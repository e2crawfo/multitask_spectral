1066 11
5 4 13 3 9 2
2 11 11
12 9 9 13 11 9 9 11 11 7 11 11 2
16 16 9 13 9 13 15 9 9 2 4 13 9 15 3 3 2
7 3 13 15 1 11 9 2
17 1 9 13 9 9 12 9 9 9 2 7 3 13 3 9 9 2
12 11 7 11 13 9 2 15 1 13 0 9 2
22 2 15 12 13 13 0 9 2 0 9 2 2 15 9 15 13 15 7 15 9 2 2
15 15 9 13 0 2 15 0 9 4 13 9 1 0 9 2
17 0 9 11 2 12 2 13 16 0 9 2 0 2 0 2 0 2
9 11 13 3 9 9 0 9 1 2
13 11 9 13 3 3 3 11 11 16 3 11 11 2
9 15 9 1 4 0 9 9 13 2
25 9 2 3 11 0 9 9 3 13 7 11 9 3 9 13 2 13 3 0 9 9 0 9 9 2
13 3 0 9 2 0 9 9 2 4 13 0 9 2
27 3 3 0 9 16 9 2 15 13 9 0 9 9 2 2 13 11 12 9 9 2 9 7 9 9 2 2
18 3 4 11 13 9 3 9 2 3 0 9 16 3 9 2 16 11 2
10 9 2 15 11 13 2 13 0 9 2
14 11 13 9 12 9 2 11 13 0 11 9 9 1 2
13 16 11 13 2 3 13 0 0 9 9 9 13 2
11 16 11 13 2 13 15 9 1 12 9 2
12 3 9 7 9 13 4 15 12 9 9 3 2
15 9 2 16 9 9 9 13 13 2 13 3 12 9 9 2
22 3 13 15 12 9 9 2 3 11 13 3 9 16 11 2 11 3 13 9 11 9 2
11 3 4 0 7 0 9 11 9 9 13 2
20 7 3 11 4 13 0 9 9 11 13 2 2 13 9 11 2 9 9 2 2
5 13 3 13 9 2
10 3 15 13 2 3 4 13 9 9 2
10 13 2 2 6 0 2 3 15 2 2
21 13 12 9 9 2 3 11 0 9 13 9 2 15 0 9 1 13 13 11 11 2
16 11 13 11 2 16 15 13 9 9 2 3 13 0 9 9 2
12 9 12 4 11 9 13 9 9 11 11 1 2
14 9 7 11 1 13 0 9 2 15 13 11 7 11 2
19 11 7 11 2 15 3 11 9 13 2 13 9 9 13 13 11 0 9 2
33 3 2 12 9 3 11 11 1 9 13 13 11 11 9 15 2 16 9 9 9 4 13 0 9 2 3 9 13 15 9 9 13 2
12 11 13 9 9 9 9 11 1 0 9 9 2
24 2 6 3 15 4 13 3 3 2 15 3 0 9 2 13 9 7 15 2 2 13 11 9 2
14 11 13 0 9 11 9 1 15 0 9 0 9 9 2
25 0 2 15 15 11 9 3 13 4 2 13 9 9 9 0 9 2 15 11 3 13 3 4 13 2
7 11 4 4 3 11 13 2
16 16 15 12 9 13 9 13 2 3 11 3 13 11 9 3 2
12 7 11 13 2 16 13 2 16 9 4 13 2
10 11 13 3 9 15 9 7 9 1 2
17 2 11 9 1 13 11 0 0 9 2 2 13 9 12 9 1 2
4 15 4 13 2
11 1 9 0 9 13 9 9 13 3 9 2
20 9 13 0 9 9 11 11 2 15 13 9 9 0 13 7 3 3 9 13 2
6 3 13 11 0 9 2
14 9 0 9 4 0 9 3 13 7 15 0 9 13 2
19 15 9 13 11 9 3 3 2 16 0 9 9 0 9 13 3 9 9 2
17 11 13 9 3 2 13 3 13 11 11 2 16 15 13 9 13 2
20 11 11 13 0 9 13 0 9 2 11 4 13 2 16 15 4 13 9 13 2
9 3 0 9 13 11 11 9 9 2
9 9 9 13 9 3 0 9 13 2
24 9 0 9 13 13 2 3 13 15 3 9 9 9 11 11 7 11 11 1 15 12 13 13 2
17 0 9 7 0 9 13 9 3 3 7 0 11 13 15 3 3 2
15 9 1 9 3 13 7 9 9 9 1 13 15 0 9 2
14 15 2 15 13 9 9 2 4 13 3 3 11 9 2
17 3 13 0 9 0 15 9 13 2 15 4 3 9 15 3 13 2
16 3 0 13 2 16 11 4 3 13 12 9 7 13 9 11 2
18 9 0 0 9 9 13 3 0 9 0 9 3 11 9 0 0 9 2
4 9 13 11 9
2 11 11
13 15 1 13 9 11 9 0 9 9 12 9 9 2
15 11 9 13 9 11 11 9 2 9 2 9 9 0 9 2
10 9 13 12 9 9 2 7 3 9 2
9 0 9 13 12 0 9 9 9 2
22 11 7 9 9 9 13 3 3 12 11 9 2 11 9 11 11 7 11 9 11 11 2
12 11 13 2 16 3 4 13 15 11 1 15 2
13 2 15 13 3 13 11 2 2 13 15 3 9 2
12 11 9 13 12 9 2 15 9 15 13 13 2
11 11 9 13 12 9 3 12 9 3 9 2
17 11 4 13 3 2 2 11 1 13 2 11 9 9 9 2 11 2
5 11 13 11 9 2
7 3 16 11 9 13 0 2
2 3 2
12 11 9 13 0 2 16 15 4 4 9 13 2
31 9 3 11 9 16 3 9 13 9 9 13 11 9 9 9 9 9 9 2 13 11 9 9 2 16 15 9 9 9 13 2
19 0 11 13 11 9 15 9 9 3 2 16 15 4 9 3 13 0 9 2
8 0 13 3 9 9 9 9 2
12 11 9 13 12 9 2 15 13 1 12 9 2
14 15 9 13 13 3 9 3 9 9 7 0 9 9 2
7 9 1 4 3 9 13 2
14 3 13 9 1 11 9 15 0 2 0 2 9 9 2
19 9 13 9 9 3 11 2 15 13 12 12 9 11 9 12 9 9 11 2
10 9 2 13 9 12 9 12 11 9 2
26 15 13 11 3 9 11 9 11 9 2 15 13 12 11 9 9 9 13 9 7 13 9 12 9 9 2
8 0 9 13 12 12 9 1 2
12 11 9 4 11 9 3 3 3 0 9 13 2
15 3 2 16 9 13 9 0 9 2 13 11 3 15 13 2
16 1 11 9 11 13 11 9 9 9 7 9 13 12 9 9 2
33 15 13 9 3 2 16 13 0 9 3 13 2 2 13 11 7 13 3 2 16 11 9 13 3 11 9 9 13 7 13 9 9 2
6 11 13 11 9 9 2
9 15 9 13 11 9 7 9 9 2
14 9 13 3 2 16 9 9 9 15 11 1 4 13 2
14 11 9 9 1 13 9 2 3 9 13 15 3 13 2
23 2 16 11 13 11 9 9 2 3 4 4 11 9 13 2 2 13 11 13 9 0 9 2
8 9 9 11 13 11 9 13 2
16 15 1 13 11 0 9 15 9 0 9 11 9 9 11 11 2
15 2 15 4 3 13 2 16 15 9 13 2 2 13 11 2
4 3 13 9 11
10 9 13 3 11 9 9 1 11 11 2
13 3 13 11 9 2 16 11 11 4 3 13 9 2
6 15 13 3 0 9 2
7 12 9 13 3 0 9 2
14 3 13 3 9 9 2 6 2 2 13 11 9 9 2
11 9 13 3 2 16 9 4 13 12 9 2
16 11 9 1 13 9 2 16 15 13 13 3 0 16 0 9 2
7 11 9 0 9 13 11 2
17 9 2 9 2 0 9 9 2 3 0 9 2 13 11 9 9 2
22 3 13 11 9 9 2 9 11 9 9 11 9 9 9 11 11 2 9 9 7 9 2
7 9 9 13 9 9 3 2
17 15 4 13 3 2 16 15 13 9 9 11 9 7 11 9 9 2
12 2 15 9 13 15 9 3 2 2 13 11 2
12 11 13 9 13 3 12 9 9 9 0 9 2
16 11 9 9 9 12 12 9 12 9 13 3 9 2 13 11 2
5 13 3 9 9 2
6 3 13 9 3 13 2
18 2 16 13 2 3 4 9 13 0 9 0 9 9 2 2 13 11 2
16 15 13 3 9 2 3 13 0 9 1 3 9 3 11 9 2
15 9 13 0 9 7 3 13 11 9 3 15 9 9 13 2
13 15 9 0 11 15 4 13 2 9 13 9 0 2
33 11 11 2 9 1 9 13 2 16 13 15 0 9 1 2 13 3 9 9 9 3 7 3 3 3 16 13 0 9 15 3 13 2
9 9 13 0 9 7 0 9 1 2
16 15 15 9 4 9 13 0 9 2 15 13 9 1 3 0 2
25 15 13 3 15 0 2 0 16 0 9 2 3 12 12 0 9 9 0 0 9 7 0 0 9 2
5 9 4 13 13 2
14 15 13 0 9 3 7 3 4 9 9 9 3 13 2
8 15 13 9 9 9 0 9 2
30 9 13 12 9 2 7 11 2 15 13 12 12 0 7 15 13 9 9 0 9 9 1 2 13 3 13 13 3 9 2
17 15 13 15 9 2 15 4 13 3 2 16 9 13 15 15 1 2
12 2 0 9 13 15 2 2 13 9 1 9 2
14 9 13 0 9 3 15 9 2 15 13 3 9 1 2
14 9 13 0 0 9 1 9 2 15 13 9 0 9 2
15 11 13 9 7 9 13 3 0 2 16 9 13 3 0 2
22 11 13 9 1 13 2 15 13 0 0 7 0 9 2 9 9 2 3 13 15 9 2
27 15 13 3 0 9 7 9 1 0 9 2 15 9 4 0 9 2 0 9 7 3 0 9 9 0 13 2
8 0 9 13 3 1 9 9 2
12 0 9 13 3 15 9 1 2 3 9 9 2
17 2 0 9 13 15 2 2 13 9 7 0 9 13 3 11 9 2
19 3 9 1 13 12 9 0 9 3 9 1 3 13 7 13 0 9 9 2
18 3 13 9 9 1 2 13 3 9 13 16 9 7 13 3 3 3 2
6 15 13 9 0 9 2
11 12 13 0 9 9 11 11 15 1 11 2
10 9 1 13 9 1 11 3 11 1 2
4 9 13 3 2
8 7 9 13 15 0 9 1 2
8 11 13 1 0 7 0 9 2
6 11 13 15 9 9 2
6 11 13 15 9 9 2
8 11 7 12 9 13 9 3 2
5 11 13 9 9 2
7 11 13 9 9 1 3 2
6 9 1 13 9 9 2
6 11 13 15 3 9 2
5 11 13 3 9 2
5 3 9 13 3 2
12 11 13 3 1 12 9 1 9 9 9 9 2
6 11 13 15 3 3 2
5 11 13 9 3 2
4 11 13 9 2
6 11 13 9 9 1 2
7 11 13 3 12 9 1 2
4 11 13 3 2
5 9 9 13 9 2
12 9 3 0 11 7 11 13 9 1 9 3 2
5 9 13 9 9 2
6 11 13 15 0 9 2
9 11 4 9 9 13 3 0 9 2
3 11 13 2
5 11 9 13 9 2
6 9 11 13 9 9 2
4 11 13 9 2
6 11 13 9 9 9 2
7 11 13 3 15 0 9 2
6 11 13 3 9 3 2
6 11 13 15 1 3 2
5 9 13 9 9 2
5 9 9 13 3 2
11 7 3 13 3 0 16 3 0 9 9 2
5 11 13 15 9 2
4 11 13 9 2
5 11 13 9 1 2
7 9 0 9 13 9 1 2
7 9 0 9 13 15 3 2
5 11 13 9 9 2
6 11 13 11 3 3 2
6 11 13 15 0 9 2
9 11 13 3 0 9 9 11 3 2
7 9 13 1 9 3 13 2
8 9 9 9 3 3 13 9 2
12 15 9 9 13 9 0 9 9 1 9 1 2
7 9 13 15 9 8 9 2
7 11 13 15 9 9 9 2
5 9 13 9 9 2
4 3 13 3 2
5 9 9 13 9 2
6 9 13 12 9 9 2
11 9 9 12 12 13 15 9 9 0 9 2
6 9 13 15 11 3 2
5 9 13 9 3 2
4 9 13 3 2
6 9 4 3 3 13 2
7 3 9 13 15 9 3 2
7 11 13 15 3 9 1 2
8 7 9 13 15 3 0 9 2
15 7 0 9 13 0 7 0 9 15 0 0 9 9 13 2
6 11 3 13 11 1 2
4 11 13 9 2
9 7 3 15 12 9 0 9 13 2
6 7 13 9 3 3 2
5 7 13 1 9 2
6 11 13 11 15 3 2
5 11 13 3 9 2
4 11 13 9 2
6 9 13 3 0 9 2
7 0 9 13 11 15 9 2
4 11 13 3 2
8 3 13 0 9 1 15 13 2
4 9 13 9 2
5 9 13 9 9 2
9 12 9 1 13 9 3 3 9 2
5 12 9 13 9 2
3 9 13 2
5 9 13 9 3 2
5 11 13 11 3 2
6 3 15 3 11 13 2
4 15 13 9 2
4 15 13 9 2
6 15 4 13 0 9 2
9 15 9 13 15 3 9 9 9 2
7 15 0 9 13 3 9 2
12 9 12 13 11 11 9 11 9 1 0 9 2
8 9 12 1 13 9 1 9 2
6 9 12 13 9 9 2
5 9 12 13 9 2
13 1 9 13 9 7 0 9 1 1 9 9 9 2
5 9 1 13 9 2
8 9 13 3 15 3 0 9 2
8 3 13 3 0 9 9 9 2
9 15 8 9 1 11 13 3 3 2
9 15 15 3 0 9 13 9 3 2
7 3 13 15 15 1 9 2
7 9 13 0 9 1 9 2
5 0 9 13 3 2
4 3 13 11 2
6 0 9 13 15 9 2
8 9 13 9 9 11 9 11 2
10 0 7 0 9 13 0 9 15 1 2
6 1 15 9 13 9 2
4 9 13 9 2
9 11 13 15 0 11 15 9 1 2
5 15 9 13 9 2
8 15 0 9 13 15 3 9 2
7 3 15 0 9 13 4 2
6 3 15 9 3 13 2
6 7 15 13 3 3 2
11 16 9 3 9 9 1 9 13 9 13 2
7 16 11 0 9 9 13 2
6 16 11 9 3 13 2
6 16 9 9 13 4 2
7 16 9 9 9 1 13 2
5 3 13 9 9 2
4 3 13 9 2
6 3 15 3 9 13 2
6 9 13 1 9 3 2
10 9 13 0 9 3 9 7 15 9 2
6 9 1 13 9 3 2
5 9 13 9 3 2
6 9 1 13 9 9 2
5 9 13 15 9 2
7 9 13 15 9 9 3 2
6 9 13 3 1 9 2
7 1 9 13 0 0 9 2
9 0 9 9 13 0 9 1 3 2
10 3 9 13 3 1 9 0 9 1 2
4 13 9 9 2
4 13 9 3 2
5 13 9 9 1 2
5 13 15 9 1 2
5 13 9 9 3 2
4 13 9 9 2
5 13 9 9 1 2
5 13 9 15 9 2
4 13 9 9 2
5 13 12 9 1 2
6 13 9 1 9 3 2
4 13 9 3 2
5 9 13 15 9 2
5 9 13 9 1 2
7 9 13 3 7 3 9 2
5 11 13 9 1 2
7 9 13 3 9 15 3 2
5 3 13 9 3 2
8 9 13 0 9 1 0 9 2
6 11 13 3 9 1 2
5 11 13 3 9 2
6 9 13 11 9 9 2
6 15 13 9 1 9 2
4 11 13 9 2
6 15 13 3 9 9 2
5 11 13 3 9 2
5 11 13 9 1 2
4 11 13 3 2
4 11 13 9 2
8 9 0 9 13 15 1 9 2
4 15 13 3 2
7 15 13 9 15 9 9 2
5 15 13 3 9 2
6 15 13 9 3 3 2
19 1 15 0 12 12 0 0 7 15 9 3 0 9 13 9 1 11 9 2
5 9 13 9 3 2
7 9 13 9 9 9 9 2
7 9 13 0 9 3 9 2
3 9 13 2
4 9 13 9 2
5 9 13 9 3 2
3 11 13 2
8 15 13 11 3 3 15 1 2
7 11 13 9 1 9 3 2
6 9 4 13 12 8 2
8 15 13 9 9 1 9 9 2
6 15 13 3 9 3 2
7 9 1 13 9 12 9 2
7 11 13 15 9 15 9 2
5 15 13 9 1 2
6 9 11 13 3 9 2
6 9 13 15 3 9 2
6 15 13 0 9 9 2
8 15 13 0 9 9 9 1 2
6 15 13 9 9 1 2
4 15 13 9 2
10 15 1 13 9 15 0 9 0 9 2
5 15 13 9 1 2
6 9 0 9 13 9 2
5 9 13 9 3 2
8 9 2 15 15 3 9 13 2
10 15 9 1 13 12 15 11 9 11 2
10 15 9 1 13 15 15 9 9 3 2
9 9 4 13 1 9 9 9 1 2
11 8 11 13 16 9 9 0 9 9 1 2
10 3 4 15 3 9 1 13 9 13 2
5 15 13 9 3 2
5 11 13 3 9 2
6 3 13 1 9 3 2
5 15 13 9 1 2
6 15 13 0 9 9 2
5 15 13 3 9 2
8 15 13 9 1 0 9 1 2
5 15 13 3 3 2
10 15 13 9 1 0 9 1 0 9 2
4 15 13 9 2
6 15 13 9 11 1 2
7 15 13 15 9 9 3 2
4 15 13 11 2
8 15 13 3 16 9 15 9 2
5 15 13 9 1 2
5 15 13 0 9 2
6 9 13 3 9 1 2
5 9 13 9 9 2
5 9 13 9 9 2
8 3 1 9 9 13 15 9 2
9 3 13 11 3 3 3 0 9 2
6 3 13 15 3 3 2
5 3 13 9 9 2
8 15 9 1 13 15 9 3 2
10 3 15 3 0 9 7 9 13 3 2
9 11 13 3 1 0 9 9 1 2
5 11 13 0 9 2
9 7 3 13 9 9 9 9 3 2
5 7 9 13 13 2
8 0 9 13 3 1 9 3 2
11 0 7 0 9 13 3 3 15 0 9 2
6 0 9 13 15 9 2
5 9 13 15 1 2
6 9 0 9 13 9 2
6 4 9 0 9 13 2
8 9 11 13 9 0 11 9 2
9 12 9 4 15 1 9 9 13 2
4 9 13 9 2
5 9 13 0 9 2
6 9 13 9 1 3 2
5 9 13 15 9 2
8 3 13 0 1 9 12 9 2
5 11 13 9 3 2
4 9 13 13 2
4 11 13 9 2
6 11 9 11 13 9 2
5 9 13 3 3 2
5 9 9 13 3 2
6 0 9 9 13 11 2
4 9 13 9 2
7 0 9 13 15 3 9 2
9 0 4 1 9 15 9 3 13 2
8 9 13 9 1 3 1 9 2
4 9 13 3 2
5 9 13 9 1 2
5 9 13 9 9 2
3 9 13 2
4 9 13 3 2
5 9 13 9 1 2
6 11 13 3 9 9 2
3 13 9 2
8 13 0 9 3 0 0 9 2
5 13 9 1 3 2
5 9 9 13 9 2
6 3 13 15 9 1 2
5 9 13 9 13 2
5 11 13 9 9 2
8 0 9 13 9 3 15 1 2
9 9 3 0 9 13 11 15 9 2
9 9 0 9 13 9 1 15 9 2
5 11 13 9 3 2
6 11 13 0 9 1 2
5 11 13 15 9 2
11 0 9 13 15 3 3 7 3 16 0 2
6 3 13 11 15 9 2
5 15 13 15 9 2
5 11 0 9 13 2
9 11 13 11 11 9 15 9 0 2
6 15 13 0 9 3 2
8 3 13 0 9 0 9 9 2
5 9 13 3 3 2
5 15 13 15 0 2
5 15 13 9 9 2
5 15 13 9 9 2
8 15 0 0 9 13 9 9 2
8 9 1 13 11 15 9 9 2
8 3 9 1 13 15 15 3 2
7 9 13 3 3 9 9 2
7 13 15 1 9 3 9 2
5 13 9 9 3 2
7 13 9 15 9 9 3 2
4 13 15 9 2
3 13 3 2
4 13 15 0 2
4 13 9 1 2
4 13 0 9 2
4 13 9 3 2
5 13 11 9 3 2
5 11 13 9 3 2
13 9 13 3 1 15 9 1 0 9 3 9 1 2
4 9 13 3 2
5 9 13 9 9 2
7 15 13 9 15 9 3 2
8 11 13 3 15 9 3 13 2
5 15 9 13 11 2
7 3 13 9 3 16 9 2
6 13 3 1 9 9 2
5 13 11 9 1 2
6 13 9 1 9 1 2
4 13 12 9 2
4 13 3 3 2
5 13 3 15 9 2
4 13 9 1 2
4 13 9 9 2
5 13 9 1 3 2
5 13 3 9 1 2
6 13 0 9 9 1 2
3 15 13 2
7 3 15 3 1 9 13 2
7 15 9 15 9 9 13 2
7 3 13 15 9 9 11 2
5 3 13 9 9 2
8 3 13 0 9 0 9 9 2
9 3 13 0 9 0 9 9 9 2
5 15 13 3 3 2
14 3 9 12 1 13 9 12 0 9 9 9 9 9 2
9 15 9 1 15 3 9 3 13 2
6 9 13 9 16 9 2
12 13 15 9 9 3 0 9 2 15 0 1 2
5 13 15 12 9 2
4 13 9 9 2
6 9 13 9 1 3 2
7 3 4 15 13 11 1 2
17 3 13 9 0 9 0 15 9 7 9 1 9 1 0 9 9 2
5 3 13 11 9 2
6 3 13 15 0 9 2
7 3 13 15 12 9 9 2
6 3 13 11 9 3 2
6 3 13 15 9 3 2
7 0 9 13 15 3 3 2
7 3 4 15 3 11 13 2
4 13 11 9 2
5 13 9 9 9 2
5 13 9 1 9 2
5 13 9 1 9 2
9 13 9 1 9 0 0 0 9 2
6 13 0 9 3 13 2
4 13 9 9 2
4 13 12 9 2
4 13 9 3 2
3 13 3 2
5 13 9 1 3 2
4 13 15 9 2
5 13 9 9 1 2
8 13 1 11 9 1 9 13 2
5 13 9 0 9 2
4 13 9 3 2
7 13 9 12 7 12 9 2
4 13 3 11 2
4 13 9 9 2
7 9 1 13 0 9 9 2
8 3 16 9 13 15 15 9 2
5 9 13 9 3 2
6 9 13 15 11 3 2
5 9 13 9 9 2
5 0 9 13 9 2
6 11 13 9 15 13 2
5 11 13 9 1 2
4 9 13 9 2
4 9 13 9 2
4 13 9 9 2
5 13 9 1 9 2
5 13 1 9 3 2
4 13 15 9 2
3 13 3 2
4 13 9 1 2
4 13 9 1 2
4 13 9 3 2
4 13 15 9 2
5 9 13 9 1 2
5 9 13 3 9 2
5 15 3 13 9 2
7 3 13 1 9 0 9 2
5 11 13 11 9 2
6 9 13 0 0 9 2
5 15 9 13 9 2
6 9 4 9 9 13 2
6 15 13 3 15 9 2
5 15 13 15 3 2
5 15 13 3 9 2
10 15 13 9 9 9 15 9 1 3 2
10 15 13 15 9 11 9 3 3 3 2
4 15 13 9 2
6 15 13 9 0 9 2
4 15 13 13 2
4 15 13 3 2
7 15 13 9 1 0 9 2
6 11 13 9 1 9 2
6 15 4 13 11 9 2
9 15 4 3 13 15 9 9 1 2
5 15 13 9 3 2
5 9 13 15 1 2
5 15 13 9 3 2
6 15 13 3 15 1 2
7 15 13 0 9 9 9 2
6 15 13 15 3 9 2
6 15 13 15 9 13 2
6 15 13 15 3 3 2
7 15 13 15 9 1 9 2
8 15 13 15 9 9 9 9 2
7 15 13 15 9 1 9 2
8 15 13 15 1 0 9 9 2
6 15 13 3 0 9 2
4 15 13 9 2
8 15 13 9 9 0 0 9 2
5 15 13 9 1 2
10 15 13 0 9 1 0 9 9 1 2
4 15 13 3 2
7 15 13 16 9 1 9 2
4 15 13 9 2
5 15 13 9 3 2
4 13 9 3 2
3 13 9 2
5 13 9 1 3 2
4 13 9 13 2
6 13 15 9 15 9 2
7 15 13 9 11 11 1 2
6 15 13 9 1 9 2
5 15 13 9 9 2
5 15 13 11 9 2
6 15 13 3 9 3 2
6 15 13 9 9 1 2
4 15 13 3 2
4 15 13 3 2
7 15 13 0 9 9 3 2
4 15 13 9 2
9 15 13 3 3 9 1 3 3 2
6 15 13 0 0 9 2
6 15 13 3 11 9 2
5 15 13 11 9 2
5 15 13 3 9 2
5 15 13 9 3 2
5 15 13 15 9 2
6 9 13 9 9 3 2
7 9 1 13 9 0 9 2
5 9 13 15 9 2
4 9 13 9 2
5 9 13 0 9 2
7 3 3 3 9 3 13 2
10 0 1 0 9 13 11 9 1 3 2
8 15 0 0 9 13 9 9 2
10 15 0 9 1 13 9 15 9 15 2
8 9 13 9 15 0 9 3 2
4 11 13 9 2
6 11 13 15 9 9 2
5 9 13 0 9 2
5 9 13 12 9 2
6 0 11 13 3 9 2
7 11 13 3 15 1 3 2
6 9 13 9 0 9 2
9 3 9 9 13 1 9 0 9 2
4 9 13 3 2
8 11 13 1 9 0 9 9 2
6 11 4 3 13 9 2
8 11 9 9 13 9 7 9 2
5 11 13 11 9 2
6 11 13 9 15 1 2
4 13 9 1 2
4 13 3 9 2
3 13 9 2
5 13 9 1 3 2
3 13 9 2
4 13 15 0 2
4 13 9 9 2
7 13 9 1 3 7 3 2
5 13 9 1 3 2
6 13 9 1 16 0 2
4 13 15 9 2
4 13 3 3 2
4 13 3 13 2
4 13 9 3 2
4 11 13 9 2
9 0 9 13 9 9 1 9 1 2
8 0 9 13 9 9 1 9 2
9 0 9 13 9 9 1 9 1 2
11 0 9 13 9 9 1 1 9 9 1 2
10 0 9 13 9 9 1 9 1 3 2
8 0 9 13 9 9 1 9 2
4 13 9 3 2
6 13 9 9 9 3 2
6 13 9 9 1 9 2
7 13 9 1 9 1 9 2
6 13 9 15 9 3 2
5 13 15 3 3 2
6 13 15 9 1 3 2
6 13 15 9 9 13 2
6 13 9 15 3 3 2
4 13 15 9 2
4 13 9 3 2
5 13 9 1 9 2
6 9 13 13 1 9 2
7 3 13 9 9 9 1 2
4 9 13 9 2
6 9 13 3 0 9 2
6 9 13 9 1 9 2
4 9 13 9 2
7 9 13 9 9 1 3 2
6 9 13 9 0 9 2
6 9 13 9 0 9 2
4 9 13 3 2
4 9 13 9 2
6 9 13 9 15 9 2
7 9 13 0 9 1 9 2
5 9 13 15 9 2
5 9 13 15 9 2
4 13 9 1 2
4 13 9 9 2
5 13 9 9 1 2
3 13 3 2
4 13 9 1 2
4 13 15 0 2
4 13 9 1 2
5 13 9 1 3 2
4 13 9 3 2
4 13 9 3 2
3 9 13 2
4 9 13 3 2
4 9 13 3 2
7 11 0 9 13 15 9 2
5 11 13 9 15 2
10 3 12 9 1 4 11 1 13 9 2
12 3 4 9 12 0 9 1 3 13 15 9 2
8 3 4 9 3 13 0 9 2
7 3 12 9 4 15 13 2
6 7 3 13 3 9 2
5 13 9 9 0 2
5 13 9 9 9 2
5 13 9 9 9 2
7 13 15 9 0 9 3 2
5 13 15 9 9 2
6 13 9 9 12 12 2
5 13 9 3 9 2
6 13 0 9 9 3 2
5 13 9 9 9 2
5 13 9 1 9 2
3 13 9 2
5 11 13 9 9 2
6 0 9 1 13 9 2
11 9 2 15 3 0 9 3 9 4 13 2
7 9 9 13 15 0 9 2
5 9 13 3 9 2
9 9 9 4 9 9 15 9 13 2
8 0 9 0 9 13 9 1 2
7 9 13 3 0 0 9 2
5 9 4 3 13 2
9 9 13 11 9 1 15 1 3 2
9 9 0 9 1 4 13 0 9 2
5 9 1 13 9 2
5 9 13 3 9 2
3 9 13 2
6 9 13 15 0 9 2
8 9 13 1 0 0 9 3 2
8 9 13 9 2 9 7 9 2
5 9 13 9 9 2
5 9 13 9 1 2
6 9 13 15 0 9 2
5 9 13 9 9 2
6 9 13 12 9 9 2
5 9 13 12 9 2
6 3 13 15 9 3 2
5 3 13 9 9 2
5 9 13 3 9 2
10 0 9 13 15 9 11 9 3 3 2
9 0 11 13 1 9 0 9 13 2
6 11 13 9 9 1 2
7 9 13 3 3 7 3 2
5 11 13 3 3 2
10 0 9 13 15 9 1 0 0 9 2
11 7 13 3 9 9 9 1 7 15 9 2
5 13 1 9 9 2
5 13 15 9 1 2
4 13 3 3 2
4 13 9 9 2
3 13 3 2
5 13 9 1 3 2
13 11 4 16 9 9 1 0 9 3 9 9 13 2
7 9 13 11 3 9 1 2
5 13 9 1 9 2
4 13 0 9 2
5 13 9 9 13 2
7 0 9 13 15 0 9 2
6 9 13 9 7 9 2
6 9 13 0 0 9 2
7 9 9 1 13 9 9 2
7 11 13 1 9 9 13 2
5 11 13 9 3 2
7 9 13 9 9 9 13 2
8 11 13 9 1 9 1 9 2
9 11 13 9 1 9 1 9 13 2
8 9 13 3 9 1 15 9 2
6 9 13 9 9 9 2
5 9 13 1 9 2
6 9 13 9 1 9 2
6 9 13 9 1 13 2
6 9 13 9 9 9 2
5 9 13 11 9 2
9 15 9 13 9 1 9 9 9 2
9 15 9 13 9 1 9 9 9 2
5 9 13 11 9 2
5 11 13 1 9 2
5 9 13 11 11 2
7 11 13 9 9 9 9 2
6 9 13 9 9 9 2
4 9 13 9 2
7 9 13 3 9 1 9 2
6 9 13 9 9 0 2
7 11 13 9 9 1 13 2
5 11 13 9 13 2
8 11 13 9 1 9 9 13 2
9 11 13 9 1 9 9 9 1 2
8 9 13 9 9 1 9 9 2
5 9 13 9 1 2
5 9 13 1 9 2
3 9 13 2
7 9 13 9 1 9 9 2
8 9 13 9 1 9 1 9 2
5 9 13 9 9 2
5 9 13 9 1 2
6 9 13 9 9 1 2
9 9 13 9 1 9 9 9 1 2
8 9 13 9 1 9 9 1 2
6 1 9 13 9 9 2
7 9 13 9 9 15 1 2
6 9 13 1 9 9 2
6 9 13 9 9 9 2
5 1 9 13 9 2
6 11 13 9 9 9 2
6 11 13 9 1 13 2
5 9 13 9 9 2
5 9 13 11 9 2
7 11 13 9 9 9 13 2
5 11 13 12 9 2
7 11 13 1 9 9 1 2
7 11 13 9 7 9 1 2
5 9 13 9 0 2
6 9 13 9 9 0 2
8 9 9 13 11 1 9 11 2
4 9 13 9 2
5 11 13 11 11 2
5 9 13 9 9 2
7 9 13 9 1 9 9 2
8 9 13 9 1 9 1 9 2
6 11 13 9 3 0 2
4 11 13 9 2
9 9 13 9 1 0 9 9 1 2
8 9 13 3 1 9 9 1 2
6 9 13 9 3 0 2
6 11 13 9 9 0 2
8 9 13 9 9 1 9 9 2
8 9 13 9 9 9 9 13 2
4 11 13 9 2
8 11 13 1 9 9 9 1 2
4 9 13 15 2
9 9 13 9 1 9 1 11 9 2
5 11 13 15 3 2
6 9 13 9 9 3 2
4 9 13 9 2
6 11 13 9 3 3 2
4 9 13 9 2
6 9 13 9 9 1 2
6 11 13 9 3 3 2
8 9 13 9 1 0 9 1 2
8 9 13 1 9 0 9 1 2
5 9 13 0 9 2
5 11 13 9 9 2
6 9 13 9 9 9 2
5 9 13 9 3 2
5 9 13 9 9 2
7 9 13 12 9 12 9 2
6 11 13 9 9 9 2
4 9 13 9 2
9 9 13 1 9 11 11 9 1 2
5 9 13 9 13 2
5 9 9 13 3 2
9 9 13 1 9 9 1 9 13 2
9 9 13 1 9 9 1 9 1 2
6 9 13 9 9 3 2
6 11 13 9 9 1 2
6 11 13 9 9 1 2
5 9 13 9 9 2
5 11 13 9 9 2
5 9 13 9 13 2
8 9 13 3 3 9 9 1 2
6 11 13 9 9 9 2
6 9 13 9 9 9 2
4 9 13 3 2
7 11 13 9 7 9 1 2
4 11 13 9 2
6 9 13 9 9 9 2
6 9 13 9 1 3 2
5 9 13 1 9 2
5 9 13 9 9 2
7 11 13 9 1 9 13 2
7 11 13 9 1 9 13 2
7 9 13 9 9 9 13 2
6 0 9 13 9 0 2
6 0 9 13 9 0 2
7 9 13 9 7 9 1 2
6 11 9 13 9 1 2
5 9 13 9 1 2
7 9 13 9 7 9 9 2
5 9 13 9 1 2
6 9 9 13 1 9 2
7 0 9 13 1 11 9 2
5 1 9 13 9 2
5 9 13 9 9 2
5 9 13 9 3 2
6 9 13 9 9 1 2
6 11 13 9 1 9 2
5 9 13 9 9 2
5 9 13 9 3 2
5 9 13 9 9 2
7 9 13 9 9 3 13 2
6 9 13 9 9 9 2
8 9 13 9 9 9 9 13 2
6 9 13 3 9 1 2
6 9 4 13 9 9 2
6 9 4 13 9 3 2
5 9 13 9 9 2
6 9 13 9 9 3 2
5 9 13 9 9 2
5 11 13 9 3 2
9 9 13 9 9 1 9 9 13 2
7 11 13 11 11 9 1 2
7 9 13 9 1 9 9 2
5 9 13 9 1 2
7 9 13 9 9 1 9 2
6 9 13 9 9 9 2
7 11 9 13 9 9 1 2
5 3 13 9 9 2
5 9 13 9 3 2
4 9 13 9 2
4 9 13 9 2
5 9 13 1 9 2
5 9 13 9 1 2
6 9 13 9 9 0 2
7 9 13 9 15 9 15 2
7 9 13 9 9 9 13 2
5 9 13 1 9 2
6 9 13 9 7 9 2
4 9 13 9 2
6 9 13 9 1 9 2
5 9 13 9 3 2
7 11 13 11 11 9 9 2
7 9 13 11 11 9 9 2
6 9 13 9 9 13 2
7 11 13 1 9 11 1 2
7 9 13 9 9 9 13 2
6 9 13 9 1 9 2
6 9 13 9 9 9 2
8 11 13 1 9 9 9 1 2
5 9 13 9 1 2
6 9 13 0 9 1 2
8 11 13 9 1 11 9 1 2
6 11 13 11 9 1 2
7 9 13 9 9 1 9 2
9 11 13 11 9 1 9 9 1 2
6 9 13 9 3 13 2
6 9 13 9 0 9 2
5 15 9 13 3 2
6 9 13 9 9 1 2
7 9 13 9 1 9 9 2
6 9 13 9 11 11 2
6 9 13 9 9 1 2
6 11 13 9 9 3 2
5 9 13 9 9 2
6 9 13 9 9 9 2
8 11 13 9 9 9 1 9 2
9 11 13 9 9 9 1 9 1 2
6 9 13 9 9 0 2
4 9 13 9 2
8 11 13 9 1 9 9 1 2
7 11 13 12 9 0 9 2
4 11 13 3 2
5 9 13 9 9 2
5 9 13 9 9 2
9 9 13 9 1 1 9 9 1 2
5 9 13 11 11 2
6 9 13 9 9 1 2
5 9 13 9 3 2
5 9 13 9 1 2
5 9 13 1 9 2
5 9 13 9 9 2
6 11 13 9 1 9 2
5 9 13 9 9 2
5 11 13 11 9 2
7 9 13 1 9 9 1 2
6 9 13 9 9 9 2
8 9 13 1 9 0 9 1 2
5 11 13 11 9 2
6 11 7 11 13 9 2
4 9 13 9 2
4 9 13 9 2
5 11 13 9 13 2
7 11 13 9 9 9 13 2
6 11 13 9 9 13 2
4 9 13 9 2
5 9 1 13 9 2
7 11 13 9 9 9 9 2
6 9 13 9 11 9 2
6 9 13 9 11 1 2
7 9 13 9 9 9 13 2
2 13 2
3 13 9 2
5 9 13 9 1 2
8 11 13 11 11 11 11 1 2
7 9 13 9 9 1 13 2
5 9 13 9 1 2
5 9 13 1 9 2
7 9 9 13 3 9 9 2
5 9 13 0 9 2
4 9 13 9 2
5 11 13 9 3 2
7 11 13 9 1 9 0 2
5 11 13 1 9 2
8 9 13 9 9 9 9 1 2
5 11 13 9 0 2
4 11 13 9 2
9 9 13 9 1 9 9 9 13 2
5 9 13 9 9 2
6 11 13 1 9 9 2
9 11 13 1 9 9 9 9 1 2
6 11 13 9 9 9 2
7 11 13 9 9 9 13 2
6 11 13 9 9 3 2
6 9 13 9 9 1 2
7 0 9 13 0 9 1 2
7 9 13 9 1 9 9 2
10 11 13 9 9 1 9 9 9 1 2
7 11 7 11 13 0 9 2
5 9 13 0 9 2
6 11 13 9 9 9 2
8 9 13 9 9 1 9 9 2
5 9 13 9 1 2
5 9 13 1 9 2
6 9 13 9 1 9 2
6 9 13 9 1 9 2
6 9 13 9 9 1 2
11 11 13 9 9 9 1 1 9 9 9 2
13 11 13 9 3 9 1 1 0 9 9 9 1 2
6 11 13 9 1 9 2
6 9 13 3 9 9 2
6 11 13 9 1 9 2
7 9 13 9 9 9 9 2
6 11 13 9 9 9 2
7 9 9 13 1 9 9 2
2 13 2
5 15 13 0 9 2
5 13 3 0 9 2
5 11 13 13 9 2
6 9 13 9 13 9 2
5 11 13 9 9 2
5 9 13 9 1 2
4 9 13 9 2
5 9 13 9 9 2
5 9 13 9 9 2
6 11 13 9 1 9 2
5 9 13 9 1 2
5 9 13 9 1 2
6 11 13 9 9 9 2
6 9 13 9 9 9 2
6 9 13 9 1 9 2
5 9 13 9 1 2
8 9 13 9 1 9 0 9 2
4 11 13 9 2
7 9 13 9 1 9 9 2
5 11 13 9 9 2
5 11 13 9 1 2
5 9 13 9 0 2
7 11 13 9 9 1 9 2
6 9 13 9 9 9 2
7 9 13 9 1 9 9 2
8 9 13 15 9 1 9 9 2
6 9 13 9 9 1 2
7 11 13 9 9 9 9 2
7 11 13 9 9 9 1 2
7 9 13 9 9 9 13 2
8 9 13 9 11 9 1 13 2
5 9 13 1 9 2
7 11 13 3 9 1 9 2
6 11 13 3 9 9 2
5 11 13 9 9 2
6 9 13 15 9 3 2
5 9 13 9 9 2
6 9 13 9 9 1 2
6 9 13 9 9 0 2
6 11 13 9 9 13 2
4 9 13 3 2
5 9 13 1 9 2
4 9 13 0 2
7 9 13 9 1 9 9 2
8 11 13 3 7 3 9 1 2
6 9 13 9 9 13 2
7 9 13 9 7 9 1 2
4 9 13 3 2
5 9 13 9 9 2
6 9 13 9 9 9 2
4 9 13 3 2
27 11 7 11 8 3 3 9 15 13 2 13 15 13 7 2 7 13 3 2 11 1 13 3 3 9 7 2
2 3 14
15 15 13 15 13 15 15 3 9 1 3 0 2 14 15 13
6 14 2 11 4 13 2
16 11 13 11 13 14 9 2 13 16 13 14 0 9 15 1 2
1 14
9 14 11 13 3 12 9 13 3 2
2 3 9
22 14 14 7 11 13 16 4 13 0 9 16 15 13 14 12 9 14 13 3 8 3 2
5 15 15 13 2 8
12 15 13 12 2 3 15 13 7 15 13 3 16
2 9 14
13 7 14 3 9 13 3 16 3 12 4 13 3 16
20 14 11 13 3 15 3 12 2 7 15 13 15 12 3 3 2 14 15 13 16
1 14
7 15 13 3 3 12 3 2
