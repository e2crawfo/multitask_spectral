1552 17
22 15 13 13 10 0 9 13 1 11 1 15 13 9 1 10 9 0 1 10 11 0 2
34 3 3 15 13 10 9 1 10 9 2 13 15 10 12 0 9 1 10 9 1 12 9 1 9 1 10 0 9 1 15 12 5 13 2
17 10 11 1 10 11 1 11 2 4 13 1 10 9 1 10 9 2
37 1 10 9 1 10 9 2 13 10 9 16 15 13 1 10 9 13 15 1 13 2 13 1 0 9 10 0 9 1 9 1 9 2 9 7 9 2
28 16 4 13 13 1 10 9 0 2 10 9 2 9 13 9 1 10 11 7 1 15 13 15 1 10 0 9 2
19 10 9 1 10 12 9 4 13 1 10 9 1 10 9 0 11 11 11 2
27 10 8 13 1 10 9 1 9 1 10 9 1 11 2 7 15 13 1 13 10 9 0 1 10 9 0 2
29 11 11 11 7 11 2 11 2 9 1 11 11 2 12 1 11 1 12 2 12 2 2 9 2 9 7 9 0 2
21 11 13 10 9 0 1 10 9 1 11 2 9 0 2 9 1 11 11 2 11 2
35 12 9 3 10 9 11 11 13 1 10 9 11 11 2 3 1 0 11 1 10 9 2 1 16 13 1 9 0 10 15 9 1 10 9 2
20 11 2 11 13 16 10 9 13 9 0 13 9 0 1 9 1 10 9 0 2
31 1 9 2 13 10 9 11 10 16 13 10 11 11 2 0 16 1 11 2 7 11 13 10 9 0 7 1 3 0 9 2
21 3 3 11 4 13 10 9 2 7 11 13 1 13 1 10 9 1 16 15 13 2
12 1 10 9 2 13 12 9 1 3 12 9 2
21 10 9 0 13 10 9 1 10 15 10 9 4 13 10 9 0 1 10 11 11 2
9 3 13 15 13 1 10 9 11 2
18 11 11 13 16 11 11 13 0 1 13 10 11 1 10 11 1 11 2
16 1 9 15 13 1 11 16 13 15 1 11 3 13 1 13 2
14 13 1 10 9 2 1 15 10 0 9 1 10 9 2
5 15 13 3 0 2
16 1 12 15 13 10 9 16 13 11 1 10 15 1 10 11 2
33 11 2 11 2 11 13 10 9 7 9 0 13 1 10 9 1 11 11 2 9 1 11 2 1 10 9 1 11 7 9 1 11 2
27 13 1 10 9 7 1 10 15 1 10 9 1 11 2 1 10 9 1 11 2 7 1 10 9 1 11 2
12 3 13 9 0 2 7 3 13 1 10 9 2
36 13 1 11 11 2 7 1 10 0 11 11 11 13 10 9 2 4 13 1 10 9 11 11 10 9 1 15 15 13 10 12 9 1 10 9 2
9 1 10 9 1 11 2 13 0 2
43 10 9 3 3 7 1 10 3 9 1 10 9 15 4 1 13 10 9 0 2 16 13 16 15 13 10 9 1 11 7 3 1 10 10 9 16 13 1 10 8 2 12 2
7 10 8 13 1 0 9 2
14 1 10 9 1 12 2 13 12 9 13 1 11 11 2
32 3 15 13 0 9 16 13 9 1 9 1 0 9 2 11 11 2 2 9 13 1 9 0 2 9 2 7 0 2 9 2 2
10 1 10 9 13 12 9 7 12 9 2
23 11 13 10 9 16 3 13 2 16 13 16 10 9 4 13 10 0 9 2 13 9 2 2
27 10 9 1 11 2 1 9 2 11 11 2 13 10 9 13 1 10 9 1 11 1 10 9 0 1 11 2
28 15 13 3 0 7 13 13 10 9 1 11 7 16 4 13 1 10 11 2 1 15 10 11 13 1 10 11 2
16 10 12 1 11 2 10 11 15 13 1 10 9 1 10 11 2
34 10 11 13 10 9 13 1 11 1 11 11 1 12 7 12 1 9 1 10 9 13 1 10 9 1 9 0 13 1 11 11 1 12 2
27 13 3 7 0 16 13 1 11 3 16 13 1 11 7 11 16 13 10 9 7 10 9 1 16 15 13 2
31 11 11 11 1 10 11 7 11 2 12 1 11 1 12 2 12 1 11 1 12 2 2 13 9 0 7 9 0 1 11 2
53 10 9 1 10 9 13 13 10 9 0 7 10 9 1 3 13 10 9 0 1 10 9 0 2 16 13 9 0 9 1 9 1 11 2 11 7 11 11 2 15 1 10 0 9 2 7 1 10 9 1 10 9 2
19 1 9 2 10 9 1 10 9 0 4 13 13 1 10 9 0 9 0 2
31 15 1 9 13 10 0 9 1 10 9 1 11 2 8 10 9 13 1 10 0 9 16 13 10 9 0 1 13 10 9 2
5 11 11 1 10 11
20 13 9 1 10 11 1 11 2 3 7 1 11 2 11 7 11 1 10 11 2
19 11 11 13 10 9 0 1 0 9 1 11 2 3 13 1 10 9 0 2
12 10 9 13 9 1 9 1 13 7 13 3 2
39 3 13 1 11 7 10 2 9 2 1 13 15 0 1 10 9 2 11 13 1 10 9 0 2 15 15 4 13 1 16 15 15 13 1 10 9 1 9 2
20 13 12 12 9 7 10 9 1 12 9 5 2 1 10 9 12 9 13 9 2
8 0 1 9 2 9 7 9 2
16 11 11 13 10 12 5 1 11 1 12 1 11 11 2 11 2
13 11 13 10 9 1 9 0 1 10 10 9 11 2
10 11 15 13 7 11 3 15 15 13 2
35 3 15 2 10 9 1 12 9 4 13 15 1 10 9 1 10 9 11 11 2 3 4 13 1 9 7 3 4 13 10 9 1 10 9 2
20 10 9 1 11 13 3 13 15 13 1 9 7 2 1 10 9 2 13 3 2
33 11 13 1 10 9 0 1 11 11 1 10 15 3 13 1 0 3 1 10 9 13 1 13 9 1 11 11 3 1 10 9 0 2
36 1 11 13 10 9 1 10 11 1 10 9 1 13 15 10 9 3 0 1 10 9 2 3 15 13 10 9 1 10 9 0 11 11 1 11 2
43 10 9 13 9 1 10 11 11 0 7 15 13 1 9 1 10 9 1 10 11 11 2 1 10 9 1 10 9 1 11 11 7 13 10 0 9 1 9 1 10 9 0 2
14 13 10 15 16 13 1 13 15 7 13 10 0 9 2
34 10 9 4 13 1 10 9 11 1 11 2 9 0 7 9 0 1 10 9 1 11 2 15 1 11 11 2 0 9 13 1 10 9 2
32 10 9 0 15 13 1 10 9 1 10 9 1 10 9 7 13 10 9 1 10 9 1 10 0 0 9 2 9 7 9 2 2
43 11 11 1 11 11 2 11 2 13 10 9 0 0 1 10 11 11 2 15 13 10 9 1 10 9 1 13 7 13 10 9 7 10 9 7 9 1 10 9 1 11 11 2
9 13 10 9 13 7 10 9 0 2
20 16 15 13 10 9 1 12 2 13 3 1 10 9 7 9 1 11 2 11 2
21 11 13 10 9 13 1 10 9 13 1 10 9 1 11 1 10 9 0 1 11 2
62 1 10 12 9 2 10 9 1 11 4 13 1 10 12 5 9 2 10 12 5 13 9 2 10 12 5 13 9 2 10 12 5 13 9 2 10 12 5 13 9 1 10 11 2 10 12 5 13 1 10 9 7 10 12 5 13 1 12 7 3 9 2
19 10 9 1 10 9 13 11 11 11 2 11 11 8 11 2 11 11 2 2
47 3 4 13 10 9 0 1 10 9 3 1 10 9 1 11 11 11 2 1 10 15 15 13 9 1 10 9 1 9 1 10 9 1 9 1 13 10 9 0 7 3 0 1 10 9 0 2
13 10 9 1 10 9 4 13 1 9 0 1 12 2
61 13 13 10 9 1 11 2 16 4 13 3 1 13 1 10 0 1 13 15 1 10 9 2 13 9 1 11 2 11 7 9 0 2 1 10 9 1 13 1 0 1 9 13 1 10 9 2 1 15 15 4 13 1 10 9 1 9 1 11 2 2
13 10 9 1 9 13 1 12 9 2 2 9 5 2
11 3 4 1 13 15 9 0 7 9 0 2
46 15 1 10 9 4 4 13 1 10 0 11 11 11 2 0 13 1 10 11 1 11 1 10 11 11 2 11 11 11 11 2 11 2 7 15 3 13 10 11 2 10 9 1 9 0 2
25 15 13 16 13 12 9 1 9 5 12 9 1 9 2 7 1 10 9 13 3 12 9 1 9 2
25 1 10 9 1 10 9 15 13 16 16 13 10 9 1 10 9 12 4 13 10 9 1 12 9 2
22 1 10 9 2 11 2 11 7 10 9 1 10 11 13 3 1 10 9 1 10 11 2
28 1 10 9 10 9 13 13 1 10 9 1 12 9 0 2 7 10 9 0 13 1 10 9 16 4 13 15 2
47 10 9 1 11 1 10 11 2 11 11 2 4 13 10 9 1 13 10 9 16 13 10 0 9 1 10 0 9 1 10 9 1 10 11 1 10 0 9 1 10 9 1 10 11 7 11 2
57 13 10 9 1 13 1 10 9 0 2 13 1 15 1 10 0 9 0 1 10 9 7 16 4 13 1 10 9 1 11 1 10 9 1 9 2 7 13 1 10 9 2 13 1 10 0 9 1 10 9 16 3 13 1 11 11 2
19 1 12 10 9 1 10 9 13 1 10 11 3 7 10 11 13 10 9 2
5 10 9 13 11 2
13 10 9 1 9 13 1 12 8 2 2 9 5 2
10 13 0 9 1 10 9 12 7 12 2
38 10 9 13 3 0 16 10 9 1 9 3 4 4 13 2 1 15 15 3 3 10 9 0 4 13 1 10 9 1 9 13 1 10 9 1 10 9 2
55 1 9 2 10 9 1 9 13 0 2 7 10 9 7 10 9 13 1 10 9 16 13 10 9 1 9 1 10 9 0 4 13 10 12 1 11 1 12 1 10 11 1 11 2 13 1 11 11 2 10 9 1 9 0 2
9 11 11 15 13 0 1 10 9 2
11 10 9 13 1 9 0 7 13 1 13 2
29 10 9 1 11 11 11 7 11 11 13 16 10 9 13 0 7 0 2 7 13 10 9 1 11 1 13 10 9 2
32 1 9 1 10 9 2 15 13 13 15 10 9 1 9 0 7 13 9 2 15 1 10 9 1 10 9 0 7 1 10 9 2
8 16 13 2 13 0 7 0 2
18 11 11 13 12 9 1 12 9 1 12 9 1 11 2 11 7 11 2
24 15 13 16 10 9 1 10 9 15 13 11 1 10 9 0 1 11 2 3 1 10 11 0 2
23 10 0 9 0 1 10 9 7 10 9 1 9 1 10 0 9 13 10 0 9 1 9 2
8 11 15 13 13 1 10 9 2
40 10 9 0 1 9 0 15 13 1 13 2 1 9 2 9 1 10 9 1 9 1 2 8 2 0 1 15 1 10 9 1 9 1 10 9 7 10 9 0 2
13 13 1 9 1 10 9 0 1 9 1 0 9 2
69 11 1 11 13 10 9 1 9 1 9 1 11 2 11 2 1 10 9 12 7 10 9 12 7 16 2 0 1 11 11 2 13 10 9 1 10 9 0 1 10 11 1 11 1 12 2 16 13 15 1 10 9 1 9 1 10 15 12 9 1 9 3 3 2 12 1 12 2 2
30 10 9 1 10 11 0 0 1 11 0 2 11 11 2 13 1 9 0 7 0 13 1 10 9 2 10 9 0 2 2
7 3 15 13 9 7 9 2
39 11 11 2 13 10 9 1 11 11 2 11 2 12 1 11 1 12 2 11 2 12 1 11 2 12 2 2 13 10 9 3 0 1 11 1 10 9 12 2
15 3 10 11 11 11 12 4 1 13 9 1 10 9 0 2
26 16 1 10 11 7 10 11 11 10 9 13 3 13 1 9 1 10 9 2 4 1 13 10 9 0 2
20 10 9 13 10 10 9 7 10 9 1 10 9 11 1 10 9 1 10 9 2
53 10 12 9 2 13 1 10 9 2 13 3 9 16 10 9 0 2 1 10 9 1 10 9 1 10 9 2 13 1 10 9 7 13 1 10 9 16 10 9 2 3 16 4 13 1 9 0 1 13 3 10 9 2
16 13 1 8 5 1 9 1 10 9 1 10 9 1 10 9 2
29 1 9 2 10 9 13 13 3 7 3 1 10 9 2 1 10 9 7 0 9 2 7 13 15 16 15 13 9 2
19 13 10 9 1 9 7 1 9 0 7 0 16 13 1 8 5 1 9 2
39 10 9 1 10 11 0 7 11 1 13 15 1 10 9 1 11 13 3 0 1 15 13 1 11 1 10 11 2 10 9 1 13 1 0 9 10 9 0 2
19 3 11 13 10 9 1 10 9 0 2 7 10 11 11 15 15 13 3 2
34 10 9 13 1 13 15 1 13 1 10 9 12 2 1 0 1 9 1 10 9 1 10 0 9 0 7 1 10 9 1 9 1 9 2
52 13 16 11 13 10 0 9 0 16 13 1 10 9 0 2 7 11 11 13 10 0 9 0 13 1 10 9 7 9 0 2 10 0 9 15 13 10 0 9 1 10 9 7 9 1 9 15 13 1 10 9 2
30 7 10 0 9 2 10 9 13 10 9 1 10 11 7 13 10 0 9 1 10 9 1 11 2 13 10 9 1 11 2
15 10 9 1 10 9 15 13 0 2 7 1 0 13 0 2
45 10 9 2 11 11 11 11 2 15 13 1 10 9 1 10 9 11 11 11 11 12 2 3 7 10 9 2 10 11 2 2 11 11 2 15 13 1 10 9 1 11 11 2 11 2
53 3 10 12 9 3 0 13 15 1 10 11 7 15 1 10 11 2 16 13 1 10 11 16 13 15 1 15 1 9 1 10 9 2 16 13 15 1 10 11 2 3 13 10 9 1 9 2 3 0 1 10 9 2
16 1 10 9 1 12 2 13 12 9 13 1 10 9 1 11 2
8 15 13 3 1 10 9 0 2
24 1 9 13 10 9 1 11 16 13 1 3 9 0 7 2 1 9 2 10 3 9 1 9 2
17 15 13 10 12 5 9 1 13 9 1 9 1 1 10 9 0 2
37 10 9 2 0 2 13 16 10 9 0 15 13 3 1 7 15 0 1 3 3 13 15 16 15 13 10 9 2 7 15 16 15 13 1 10 9 2
30 1 10 9 0 7 10 9 0 13 0 9 1 9 0 2 16 3 13 0 9 1 10 9 13 10 9 1 9 0 2
18 13 1 10 9 1 11 11 7 10 9 13 1 12 9 2 12 2 2
66 1 15 2 10 9 0 2 11 11 2 13 9 16 13 10 9 1 13 13 10 9 16 13 10 0 9 1 2 3 13 15 3 1 10 0 9 7 13 16 10 9 16 13 1 3 15 13 7 1 9 13 1 9 1 9 1 10 11 1 11 2 2 13 1 11 2
36 1 13 2 10 10 9 1 10 9 13 15 13 1 3 3 13 1 9 1 9 3 0 2 1 9 0 0 15 13 2 13 10 9 2 2 2
11 11 13 10 9 0 1 10 11 1 11 2
8 2 3 4 13 10 10 9 2
37 10 9 16 13 3 15 13 9 1 10 12 9 2 15 13 2 15 4 13 9 2 15 4 1 13 7 3 16 3 13 1 11 15 4 13 9 2
9 10 9 3 0 1 11 13 11 2
25 10 9 0 13 13 10 9 0 1 10 11 0 13 1 10 9 1 9 1 10 9 1 10 9 2
37 1 10 9 10 9 3 13 1 10 9 0 10 0 9 16 13 10 9 1 12 7 12 9 13 10 9 1 16 10 9 13 1 3 1 10 9 2
20 1 9 1 9 2 10 11 13 10 3 0 1 10 10 9 13 1 10 9 2
16 11 4 13 10 9 16 4 13 10 9 1 13 10 0 9 2
23 13 10 9 0 1 13 1 10 9 2 16 13 1 9 0 15 15 4 1 13 1 9 2
14 2 4 7 13 1 10 9 9 1 16 13 9 0 2
7 15 4 13 10 0 9 2
37 1 10 9 2 1 10 12 9 4 13 9 1 9 1 10 11 11 11 11 1 11 2 1 10 15 13 10 9 1 9 1 10 9 0 2 0 2
6 15 9 1 10 3 2
18 1 13 10 9 2 1 12 13 3 1 10 9 10 2 11 11 2 2
20 10 9 1 9 4 13 1 3 1 10 9 1 10 12 2 2 13 10 9 2
49 1 12 10 0 9 0 2 11 1 11 2 3 13 1 11 11 2 2 13 10 0 9 1 13 10 9 1 11 11 2 4 10 9 13 1 10 0 9 1 11 11 1 12 16 13 3 11 11 2
62 1 10 12 9 2 10 9 1 11 4 13 1 10 12 5 0 2 10 12 5 13 0 2 10 12 5 13 0 2 10 12 5 13 0 2 10 12 5 13 0 1 10 11 2 10 12 5 13 1 10 9 7 10 12 5 13 1 12 7 3 9 2
32 11 13 10 9 7 9 0 2 1 10 9 1 11 2 9 1 11 2 11 2 1 10 9 1 11 7 9 1 11 2 12 2
53 10 9 3 13 3 1 10 0 9 1 2 9 7 0 2 2 10 9 0 7 10 9 0 2 1 10 9 2 2 7 1 10 9 0 1 16 15 0 13 1 9 2 13 1 10 0 9 2 1 10 9 11 2
14 11 13 10 9 0 1 9 9 1 10 9 0 11 2
50 13 10 9 1 11 11 1 11 12 2 7 15 13 10 9 2 10 9 2 10 9 7 10 0 7 9 1 9 16 15 13 1 10 9 1 10 9 1 10 9 2 3 1 10 9 1 3 0 9 2
48 9 9 1 10 9 2 3 13 15 1 10 9 2 13 15 13 10 9 0 1 10 9 7 3 15 4 13 1 10 9 1 13 10 9 0 1 9 2 16 8 13 3 15 2 10 9 0 2
33 4 13 1 10 11 1 10 9 0 3 1 13 10 9 12 1 10 11 2 7 13 1 9 0 1 10 11 11 10 12 1 11 2
48 1 0 9 1 9 1 9 7 9 2 7 1 10 9 0 7 13 0 1 10 9 11 11 2 10 9 13 1 11 7 13 1 11 11 11 7 11 11 11 2 13 10 9 1 13 1 11 2
10 1 3 2 15 13 1 11 11 11 2
27 10 9 16 10 9 15 4 13 15 13 16 13 1 10 10 9 2 1 10 10 9 7 1 10 10 9 2
19 13 9 0 2 1 9 3 0 1 9 1 10 0 9 0 15 13 13 2
20 10 9 1 9 15 4 13 1 9 0 2 0 2 8 2 0 7 1 9 2
9 15 13 1 11 2 11 7 11 2
30 10 9 13 10 9 1 9 7 4 13 1 10 9 1 12 16 13 10 9 16 13 1 10 9 0 16 13 10 9 2
17 1 12 11 13 1 10 9 0 1 10 11 11 11 8 11 11 2
18 15 13 10 9 0 2 7 13 16 10 9 15 13 0 1 10 9 2
39 0 1 15 7 11 2 11 15 13 1 11 3 1 16 15 13 1 10 11 11 2 1 10 9 11 13 10 9 1 15 7 15 3 13 15 9 1 15 2
38 3 2 11 13 10 9 1 11 11 1 10 9 1 16 10 9 15 13 1 16 15 13 1 10 9 1 10 15 11 15 13 1 9 0 7 15 13 2
62 3 2 1 9 0 2 3 4 13 15 1 10 9 1 10 11 2 10 9 1 10 9 13 10 0 9 3 10 9 13 3 0 15 15 13 9 2 1 10 9 2 1 10 9 1 9 7 9 13 1 9 0 1 10 9 0 7 0 1 10 9 2
15 10 11 2 7 10 9 16 15 13 2 13 1 9 0 2
23 1 10 9 1 12 9 2 11 13 10 9 0 1 10 9 1 10 8 8 2 11 2 2
32 15 15 13 1 10 9 1 10 9 7 3 1 10 9 1 9 1 11 2 13 10 9 13 1 10 9 0 1 11 7 11 2
11 10 9 1 11 15 13 13 1 10 9 2
24 4 13 1 10 9 0 11 11 2 1 10 9 9 1 11 2 1 15 13 3 1 13 0 2
42 12 9 3 3 10 12 1 11 2 9 1 10 11 11 1 11 2 11 15 13 1 10 0 9 1 12 9 16 15 13 10 8 8 1 16 11 11 15 13 1 12 2
26 13 10 9 16 15 13 1 10 11 2 11 13 3 15 1 15 16 13 13 1 10 9 0 3 3 2
12 3 13 1 11 11 1 10 9 0 1 9 2
9 13 10 9 0 1 13 1 9 2
26 10 9 11 13 10 9 1 10 12 9 1 11 16 13 9 2 13 16 11 13 1 12 1 13 9 2
22 10 9 3 0 13 2 11 11 2 11 2 2 11 11 2 11 11 11 7 11 11 2
19 9 0 2 9 0 7 9 3 3 2 0 13 10 9 1 10 0 12 2
28 15 13 16 15 9 15 13 1 10 9 1 10 9 7 10 9 1 9 3 0 2 15 13 2 10 9 0 2
12 1 0 2 10 9 1 11 11 3 13 0 2
37 15 1 10 9 2 16 15 13 16 4 13 13 10 9 2 3 15 13 1 10 9 0 1 10 9 7 13 9 16 3 15 13 1 10 0 9 2
35 15 13 10 9 16 4 13 15 1 10 9 7 13 1 10 9 12 2 11 2 3 13 9 10 1 10 9 11 2 16 13 10 0 9 2
42 1 10 9 1 10 9 1 10 11 11 2 11 13 10 9 0 1 12 9 5 2 1 10 15 12 9 5 13 1 9 0 7 2 12 5 2 12 9 5 13 9 2
38 11 13 1 10 9 7 9 1 10 12 0 9 1 10 9 1 11 11 2 3 1 10 9 1 0 9 1 10 15 10 3 9 13 10 11 1 11 2
54 10 9 0 4 13 1 9 10 9 13 1 10 9 2 13 1 10 9 2 7 3 13 10 9 7 10 9 7 4 13 10 10 9 1 10 10 9 2 10 10 9 2 10 10 9 2 2 13 10 9 1 10 9 2
19 10 9 16 13 10 9 0 1 10 9 8 13 7 13 1 4 1 13 2
12 11 13 10 9 0 1 10 9 11 1 11 2
15 3 15 13 2 7 15 15 13 3 1 9 10 9 0 2
38 10 9 0 1 11 11 11 13 10 0 9 1 11 7 11 1 10 9 1 10 9 2 1 9 4 13 11 15 4 4 13 1 10 9 1 9 0 2
37 1 10 11 2 11 2 4 13 10 9 7 15 13 16 16 13 4 13 7 1 10 3 1 10 9 16 15 13 13 1 10 9 13 1 10 11 2
22 13 0 10 1 10 9 7 15 13 1 10 9 1 10 0 9 1 9 1 10 9 2
30 13 1 12 1 11 2 11 2 2 13 10 9 1 10 9 7 1 13 1 12 15 13 1 13 1 10 9 1 11 2
44 1 10 9 1 10 12 1 11 1 12 2 11 2 10 9 11 11 2 11 11 7 10 9 1 9 13 1 12 9 1 9 1 10 9 1 11 2 11 1 10 9 1 11 2
19 10 9 1 10 9 4 3 13 1 11 1 11 2 11 11 7 11 11 2
45 11 13 10 9 3 0 1 10 15 15 13 10 9 2 10 9 7 10 9 7 10 9 2 3 7 10 9 1 10 9 1 9 0 2 9 2 9 2 9 2 9 2 9 2 8
15 11 13 10 9 3 9 0 2 1 15 1 9 7 9 2
45 1 12 2 13 1 11 11 1 10 9 1 10 9 0 1 9 1 10 0 9 2 1 12 2 7 11 13 1 0 9 1 10 9 1 9 2 1 0 9 2 7 1 9 9 2
26 1 15 2 10 9 13 10 0 9 7 13 9 1 9 16 13 1 10 9 7 10 9 0 1 15 2
17 10 9 1 10 9 1 10 11 13 1 10 9 0 1 10 9 2
25 13 9 2 9 7 9 1 10 9 1 11 7 11 2 10 9 13 1 9 7 9 1 10 9 2
32 13 1 10 9 1 10 11 11 11 2 16 3 4 13 1 10 9 1 10 11 11 11 12 16 3 15 13 1 10 9 0 2
12 9 11 7 11 1 13 15 10 9 3 0 2
10 10 11 11 13 9 1 12 1 12 2
25 1 9 1 10 9 1 9 1 10 9 2 13 10 9 12 2 8 7 8 2 1 10 9 0 2
16 1 10 9 1 12 2 13 12 9 13 1 10 9 1 11 2
25 1 10 9 3 0 2 1 9 1 9 2 15 4 13 9 2 9 2 9 2 3 1 0 9 2
35 1 9 1 16 15 13 9 0 7 3 13 7 10 10 9 13 1 10 11 11 2 10 9 4 4 13 1 9 1 10 9 13 1 10 8
15 15 13 1 11 2 11 2 11 2 11 2 11 7 11 2
19 1 10 9 1 12 2 15 13 10 9 15 15 13 10 9 1 10 9 2
35 4 13 1 10 11 1 11 1 10 9 1 10 9 0 1 10 11 11 11 2 1 10 15 13 0 1 10 9 1 9 1 11 1 11 2
38 10 12 1 11 1 12 15 13 3 10 0 9 1 10 9 1 9 1 10 9 1 9 7 1 10 9 0 7 15 13 9 1 10 9 1 0 9 2
28 9 13 1 12 9 2 13 9 1 9 1 10 11 11 2 12 2 1 10 11 7 11 1 9 2 12 2 2
42 1 10 9 1 10 9 1 10 11 11 2 11 13 10 9 0 1 12 9 5 2 1 10 15 12 9 5 4 1 9 0 7 2 12 5 2 12 9 5 13 9 2
15 3 15 13 1 9 15 13 10 9 1 10 9 1 11 2
13 7 15 1 9 0 1 9 2 7 15 13 0 2
22 15 13 9 1 0 9 1 10 9 16 4 13 9 2 9 7 10 9 1 0 9 2
10 10 10 9 0 15 13 1 10 9 2
18 4 13 10 12 1 11 1 12 1 11 11 7 13 1 11 11 11 2
32 10 9 1 9 16 13 11 1 11 2 13 1 10 9 0 2 4 13 2 16 13 1 9 0 9 16 13 1 10 0 9 2
42 3 13 10 9 1 10 16 2 3 3 1 12 9 2 15 13 11 2 12 9 1 11 2 12 1 11 7 12 1 11 2 7 12 3 1 12 7 12 2 11 2 2
28 1 15 15 4 13 1 10 9 0 16 13 10 9 7 15 13 10 9 1 10 0 9 1 9 1 10 9 2
13 11 11 11 13 10 9 1 9 1 10 9 11 2
13 10 0 9 4 4 13 1 11 8 11 2 12 2
5 15 13 1 12 2
47 1 9 1 10 9 1 10 0 9 1 10 9 1 10 9 1 10 9 9 1 11 11 2 0 2 0 7 0 13 1 12 2 10 1 10 9 1 10 9 4 13 1 0 9 1 9 2
39 10 9 13 1 0 9 16 13 3 1 10 9 1 11 1 11 2 3 7 7 13 15 1 10 3 0 9 1 10 9 0 2 11 11 11 2 12 2 2
26 10 9 13 1 9 13 1 9 2 13 1 9 1 10 9 7 10 9 2 7 13 0 1 10 9 2
24 10 9 1 9 15 13 3 1 10 9 13 1 9 1 11 2 11 11 7 10 9 11 11 2
18 1 10 9 0 1 11 1 10 0 9 2 11 7 11 13 10 9 2
16 11 11 13 0 1 11 11 2 10 9 1 10 9 1 11 2
16 11 11 2 13 1 9 10 9 1 10 9 0 1 11 11 2
69 10 11 11 1 11 13 10 9 1 10 9 11 11 12 2 11 11 11 2 1 9 2 11 11 11 11 11 2 2 11 11 11 11 11 2 2 16 16 10 2 11 11 2 4 13 0 1 2 11 11 11 2 1 11 11 11 12 10 12 1 11 1 12 1 10 9 11 11 2
32 1 10 9 2 1 12 2 10 9 11 11 1 11 2 9 7 9 1 11 11 1 11 2 15 4 13 1 10 9 1 11 2
20 13 16 13 9 1 9 7 13 3 0 1 13 7 13 10 10 9 16 13 2
30 10 11 13 8 10 9 13 1 9 11 1 3 1 12 9 2 7 8 4 13 0 9 7 9 0 1 10 9 0 2
25 13 1 12 1 10 9 1 10 3 3 13 11 11 1 11 7 11 2 15 13 13 1 10 11 2
23 15 1 10 13 15 1 10 0 9 2 13 1 10 9 7 13 10 9 1 10 9 0 2
11 15 3 13 0 9 7 3 13 15 3 2
30 10 9 1 12 9 13 1 9 1 10 9 2 12 9 0 1 10 9 2 12 9 7 12 9 3 1 9 7 9 2
35 1 15 1 10 9 1 11 11 13 10 9 1 10 9 1 11 1 11 2 3 7 10 9 0 2 11 11 2 13 10 9 1 10 9 2
20 11 13 10 9 1 11 13 1 10 9 7 9 1 10 9 13 1 10 11 2
8 10 11 11 13 10 9 0 2
25 1 10 9 4 13 1 10 9 3 4 1 13 9 0 1 10 9 1 10 9 13 1 10 9 2
33 10 9 13 10 9 1 10 9 2 0 1 10 9 2 1 9 0 0 7 0 13 3 1 10 10 9 13 1 10 9 0 0 2
30 7 1 9 13 15 9 1 9 7 15 2 7 3 13 13 15 3 1 11 7 1 9 15 13 10 12 9 1 9 2
25 9 7 9 13 1 10 9 7 10 9 9 1 10 9 13 10 9 1 9 13 1 13 15 0 2
16 1 10 9 0 3 15 4 13 11 11 2 11 2 7 11 2
23 7 10 0 9 13 9 1 0 7 0 9 0 1 10 11 2 11 2 11 7 10 12 2
19 10 9 3 13 15 1 11 1 10 9 0 7 11 7 11 1 10 9 2
16 10 9 7 10 9 4 13 1 10 9 10 9 1 9 0 2
23 15 1 10 9 13 10 9 1 10 9 1 9 2 10 9 7 9 1 0 9 1 9 2
52 10 11 11 1 11 11 11 4 13 1 12 1 10 9 1 13 10 9 3 1 9 2 1 10 9 16 13 1 9 1 9 13 10 9 1 13 2 13 7 13 10 9 2 13 10 9 0 1 9 1 9 2
53 10 9 15 13 1 10 9 0 12 1 10 9 0 1 9 0 16 13 11 1 10 11 1 10 9 0 2 1 10 9 1 11 1 10 11 7 11 2 1 10 9 1 11 1 10 11 7 1 9 1 10 11 2
27 1 9 2 10 10 9 0 15 4 13 1 11 1 10 9 2 13 11 11 11 7 10 9 11 11 11 2
11 4 13 3 1 10 9 0 1 10 9 2
8 3 13 3 0 13 1 9 2
8 13 10 12 1 11 1 12 2
34 1 10 0 9 2 11 13 13 1 11 2 11 7 11 2 10 9 3 13 10 9 1 10 9 1 11 11 2 7 10 9 13 15 2
20 11 4 13 3 3 2 7 10 9 4 3 3 13 1 11 2 10 9 0 2
18 10 9 13 15 0 2 15 16 9 1 11 2 1 11 11 2 13 2
26 11 11 11 11 11 13 10 9 0 1 10 9 0 11 11 2 13 10 12 1 11 1 10 9 12 2
16 1 10 9 1 12 2 13 12 9 13 1 10 9 1 11 2
88 10 9 0 15 13 1 10 9 1 10 11 13 1 10 9 0 1 10 9 2 1 10 16 10 9 0 7 10 9 13 10 9 0 1 10 11 11 2 9 7 9 16 13 10 9 1 10 11 11 2 3 10 9 1 10 11 1 11 15 4 13 1 10 9 16 10 9 13 1 9 1 0 9 0 2 7 10 10 9 1 10 11 1 10 11 1 9 2
57 1 10 9 15 13 11 3 16 1 10 9 1 10 11 11 1 11 1 12 2 10 9 1 11 11 13 10 9 1 16 10 9 13 10 9 2 10 15 13 10 9 1 10 0 9 11 11 2 10 9 12 1 11 1 10 9 2
23 10 9 1 11 1 9 11 15 13 1 16 11 13 0 1 13 1 10 9 0 3 0 2
29 13 1 9 2 13 9 10 9 1 9 2 13 1 10 9 1 11 1 11 2 1 10 9 1 11 11 1 11 2
19 13 1 15 15 10 9 0 2 1 10 9 2 2 8 8 2 8 2 2
9 10 9 4 1 13 15 11 11 2
24 13 1 10 11 1 11 2 7 13 10 9 0 1 13 9 1 10 9 1 10 9 11 11 2
13 1 10 9 1 12 2 11 11 13 1 10 9 2
14 10 9 1 9 4 13 0 2 7 3 4 13 9 2
28 1 10 9 1 11 16 13 3 1 10 0 9 16 15 13 10 9 2 10 9 15 13 7 11 13 9 0 2
21 15 13 16 1 10 9 1 9 1 9 4 13 15 1 15 2 9 0 7 0 2
21 10 9 0 13 10 9 1 11 2 16 16 10 9 0 15 13 1 10 11 0 2
42 13 1 10 9 1 10 9 1 11 2 1 10 9 1 10 9 1 11 2 1 10 9 1 10 9 1 11 7 10 9 1 11 7 1 10 9 1 10 9 1 11 2
39 1 10 9 1 11 2 1 12 2 11 13 1 11 2 1 15 15 4 13 10 9 1 13 9 1 10 11 7 15 13 9 1 10 9 7 1 10 9 2
18 10 9 0 1 9 7 9 13 0 1 9 0 1 9 0 1 9 2
21 10 9 1 9 4 13 15 0 1 0 9 1 9 13 1 10 0 9 1 9 2
17 13 16 10 9 13 0 2 16 3 13 13 1 10 10 9 0 2
20 3 4 13 1 10 9 7 3 1 13 0 9 1 10 9 15 13 1 13 2
29 1 15 4 7 13 1 10 0 9 1 10 9 3 0 7 15 0 7 10 9 13 1 10 0 9 2 2 13 2
24 4 13 1 9 7 9 1 9 0 7 1 10 4 13 1 10 9 13 10 9 1 10 9 2
35 11 13 10 9 7 9 0 2 13 1 10 9 1 11 2 9 1 11 2 1 10 9 1 11 7 9 1 11 2 1 2 11 2 11 2
29 3 15 13 10 9 11 11 2 15 4 13 16 2 10 9 13 0 7 13 16 10 9 0 4 13 1 9 2 2
27 10 9 1 11 2 1 9 2 11 11 2 13 10 9 13 1 10 9 1 11 1 10 9 0 1 11 2
25 16 3 13 1 10 9 0 2 11 15 13 2 1 10 9 2 1 10 9 0 0 1 11 0 2
11 1 10 0 9 13 9 1 11 1 9 2
13 15 15 13 10 0 9 1 10 9 0 0 0 2
22 10 9 2 13 9 1 9 1 10 9 2 7 16 13 3 3 13 9 1 10 9 2
37 3 3 2 0 1 10 9 1 10 9 1 10 0 9 7 10 9 3 1 10 9 2 10 9 4 1 13 1 10 9 2 7 3 2 13 0 2
45 1 10 9 1 11 10 9 4 13 1 11 2 10 9 1 11 11 2 7 13 10 9 3 11 12 15 13 11 2 9 1 11 2 2 10 9 16 15 13 10 9 1 11 11 2
17 13 1 11 11 2 11 11 2 7 13 1 11 2 11 2 11 2
30 10 9 0 4 13 1 10 9 1 10 11 12 7 10 11 12 3 1 11 11 11 1 10 9 1 11 2 11 11 2
11 3 9 13 1 11 7 15 13 1 9 2
10 13 1 10 0 9 1 10 0 9 2
6 2 11 1 9 2 2
17 13 0 1 10 9 1 10 9 7 1 10 9 1 9 15 13 2
35 13 10 9 0 2 0 1 12 7 12 2 10 0 9 0 15 13 1 10 11 1 11 2 3 13 12 9 1 9 1 10 9 1 12 2
13 10 9 13 0 2 13 10 3 0 1 10 9 2
14 11 13 13 10 9 1 13 1 11 7 3 15 13 2
16 10 9 0 1 13 10 9 1 9 7 13 10 0 9 0 2
38 13 10 9 13 10 9 1 9 1 10 9 2 13 10 9 7 1 0 3 3 3 2 3 0 1 10 9 2 15 13 10 9 16 13 3 1 8 2
18 10 9 1 8 8 13 0 7 10 8 7 9 1 13 15 1 9 2
35 1 10 9 2 10 9 13 3 9 8 5 8 2 16 13 1 10 9 13 10 9 3 1 9 1 9 2 9 1 10 0 9 1 9 2
5 4 13 1 12 2
18 3 4 4 13 1 0 9 2 1 9 1 9 0 2 1 9 2 8
7 10 9 1 9 13 3 2
18 10 11 11 12 13 10 0 0 9 1 9 1 3 0 9 1 11 2
40 10 9 1 11 1 10 13 2 9 1 9 2 13 13 15 1 9 1 10 9 0 2 0 7 0 0 1 10 9 0 7 1 10 9 13 1 13 10 9 2
61 1 10 12 9 2 11 11 12 4 13 1 10 12 5 0 2 10 12 5 13 0 2 10 12 5 13 0 2 10 12 5 13 0 2 10 12 5 13 0 1 10 11 2 10 12 5 13 1 10 9 7 10 12 5 13 1 12 7 3 9 2
10 10 9 13 1 12 13 1 12 9 2
53 15 2 13 1 16 3 13 15 3 1 10 9 2 13 1 16 3 13 10 9 11 11 11 2 7 13 1 16 10 9 15 13 1 15 13 1 10 9 0 1 10 9 3 0 2 1 3 3 12 9 1 9 2
14 10 9 11 2 11 4 13 10 12 1 11 1 12 2
14 4 13 12 9 1 10 9 0 13 10 9 3 0 2
24 10 9 13 1 10 10 9 1 9 3 0 2 10 9 0 13 3 0 7 10 9 15 13 2
22 13 16 10 9 13 1 9 13 10 9 1 10 11 11 1 11 2 3 13 1 11 2
18 3 13 13 10 9 1 10 9 0 1 11 11 1 13 15 15 0 2
26 10 9 13 3 1 10 9 1 11 11 2 1 10 0 9 2 10 9 16 13 1 11 13 11 11 2
16 10 9 1 9 15 13 1 10 9 1 9 1 10 11 11 2
33 3 1 11 2 10 11 1 11 13 10 9 3 0 1 10 0 11 2 1 10 9 16 13 1 10 1 10 0 9 1 10 9 2
27 10 9 15 13 1 10 0 9 1 9 1 16 1 10 9 4 13 10 9 1 10 9 1 10 9 12 2
77 13 0 10 0 9 1 9 2 1 15 9 2 16 4 13 3 7 3 1 9 1 9 1 9 2 13 1 10 9 0 7 13 0 9 1 10 9 2 1 10 13 10 9 0 1 10 9 2 1 9 3 1 10 9 0 1 16 15 13 10 9 7 1 7 13 10 9 0 1 10 9 0 1 13 10 9 2
31 10 9 0 4 13 1 10 9 1 12 9 2 11 2 11 2 11 2 11 2 11 2 11 2 11 11 2 11 7 11 2
15 10 11 11 11 1 11 1 10 11 15 13 1 11 11 2
25 10 9 0 1 11 11 13 15 1 10 12 9 16 13 10 9 1 11 2 13 1 10 9 0 2
14 15 13 1 10 9 13 1 12 9 13 15 1 15 2
16 8 9 15 13 0 2 15 13 10 9 7 10 9 13 0 2
12 10 9 1 11 11 15 13 0 1 10 9 2
36 8 8 13 16 10 9 13 1 13 1 10 9 13 10 9 2 16 2 10 9 15 4 13 15 3 2 1 10 9 0 2 0 7 0 2 2
45 10 9 2 16 3 4 13 15 1 11 2 15 13 1 9 1 10 9 1 9 2 16 13 1 10 9 1 10 11 11 8 11 2 16 3 13 9 0 1 10 9 0 1 11 2
39 9 1 9 13 1 10 9 1 9 7 1 10 9 1 16 3 13 0 9 1 10 9 4 13 10 11 2 12 11 2 10 9 0 1 10 3 0 11 2
48 3 2 13 15 1 10 0 9 1 10 9 1 10 9 0 1 10 9 1 10 11 1 10 11 1 9 13 10 12 1 11 1 12 16 13 1 10 11 11 11 7 1 10 11 11 1 11 2
23 3 10 0 9 13 3 0 13 10 9 1 9 2 4 15 13 10 9 1 11 7 11 2
46 2 11 13 1 16 10 0 9 1 9 13 0 2 2 1 16 10 9 4 2 13 10 9 0 3 3 1 10 0 9 1 10 9 1 9 1 15 2 7 1 10 9 1 10 9 2
60 4 1 13 10 9 0 1 10 9 1 11 2 11 11 2 10 12 1 11 1 12 2 3 10 9 11 11 13 10 9 7 13 3 1 2 11 11 11 2 2 9 1 10 9 11 2 15 10 9 13 1 0 9 1 10 9 1 10 12 2
18 1 10 9 10 9 11 11 2 9 1 11 2 15 13 1 10 9 2
14 13 1 15 9 16 13 1 10 9 2 3 10 9 2
7 10 9 15 13 3 8 2
26 1 10 9 1 10 12 1 11 1 12 13 12 9 1 10 9 1 10 9 11 2 16 13 1 11 2
44 10 9 1 10 9 13 0 2 2 11 13 0 1 15 0 7 0 2 1 9 3 0 7 0 2 10 9 1 10 9 1 11 4 4 13 1 10 9 3 0 1 11 2 2
10 13 9 0 16 4 13 1 12 9 2
12 2 13 15 10 9 1 9 1 9 1 9 2
46 13 1 10 9 0 11 11 1 10 9 11 11 11 11 11 2 15 13 1 9 1 11 7 13 9 1 9 0 1 11 11 11 11 7 11 2 3 1 13 1 11 11 1 0 9 2
29 2 4 1 4 1 13 10 9 0 2 13 10 9 1 9 1 9 0 7 0 1 11 2 2 13 10 9 11 2
24 10 9 0 2 0 13 0 2 7 10 9 0 7 0 13 3 10 10 9 0 1 10 9 2
29 10 9 0 1 10 11 11 13 2 11 2 2 16 13 10 9 0 1 10 9 1 11 2 11 1 10 9 0 2
5 2 15 13 15 2
8 10 9 0 13 2 10 9 2
39 13 10 0 9 1 10 9 1 10 9 11 16 13 10 9 1 9 2 10 9 4 13 3 1 11 11 1 10 9 13 3 0 2 13 3 1 10 9 2
25 13 1 15 2 10 9 0 15 13 1 11 13 15 1 13 10 9 3 0 1 9 1 13 9 2
43 11 13 10 9 0 7 10 9 13 1 10 9 2 3 9 2 1 10 9 13 1 9 7 9 7 9 3 0 1 9 7 3 3 0 1 9 13 16 10 9 13 0 2
25 11 13 9 1 13 9 1 10 9 1 10 9 0 1 12 1 11 7 1 11 2 3 4 13 2
23 10 10 9 16 3 13 13 10 9 11 16 13 10 9 0 1 9 1 12 9 1 9 2
19 10 9 0 13 1 10 9 1 10 0 9 7 13 3 3 9 1 15 2
37 10 9 9 13 13 2 3 1 10 9 2 7 15 4 13 1 13 15 1 0 9 16 13 3 1 10 9 1 16 13 10 9 16 13 1 15 2
14 13 10 9 1 10 9 1 16 10 9 13 13 9 2
18 1 0 3 13 9 0 2 16 3 13 10 9 1 9 1 10 9 2
27 10 9 13 10 9 1 9 1 10 9 1 10 11 1 10 11 13 1 11 11 2 16 3 13 10 9 2
25 13 9 7 1 10 3 13 9 1 9 2 13 1 13 1 10 9 9 3 2 15 15 13 13 2
41 13 10 9 0 3 1 9 1 4 13 13 2 16 13 9 1 0 9 2 7 13 9 1 13 2 16 13 9 2 2 15 13 3 1 9 16 13 10 15 0 2
21 10 9 0 0 1 10 9 1 10 9 3 13 3 0 1 10 9 1 10 9 2
43 1 10 11 1 10 11 1 10 11 11 2 10 9 13 10 9 0 1 12 5 12 2 1 10 15 12 5 12 13 1 9 0 7 2 12 5 2 12 5 12 13 9 2
15 10 0 9 1 10 9 13 1 9 1 9 1 10 9 2
42 13 1 8 1 0 9 1 10 9 2 1 9 1 10 8 3 13 2 9 12 5 0 1 0 9 7 3 1 9 3 13 15 7 15 13 1 15 9 2 10 9 2
23 10 0 9 1 10 9 13 1 9 0 1 9 0 7 0 13 1 3 15 13 10 9 2
20 1 9 1 10 9 12 10 9 4 4 3 13 1 10 9 1 10 9 0 2
27 10 10 9 1 10 9 15 4 13 2 7 15 13 0 1 10 9 1 12 9 1 9 1 9 7 9 2
19 13 9 0 1 10 9 11 2 1 10 15 13 15 1 10 3 0 9 2
22 11 1 11 2 10 11 11 13 10 0 9 0 1 10 9 0 11 11 13 1 12 2
30 1 10 0 2 0 9 2 13 10 0 9 2 3 0 2 1 10 15 3 13 11 11 13 1 10 9 1 9 2 2
11 15 1 10 9 1 10 9 0 0 0 2
9 11 11 13 1 10 9 1 11 2
43 9 0 1 10 9 3 0 1 10 9 1 10 9 1 10 9 1 10 11 1 10 11 2 9 2 9 7 9 1 8 8 2 1 10 9 13 10 9 1 10 9 0 2
29 11 11 13 12 9 16 13 3 1 10 9 2 10 0 11 11 2 7 10 9 11 11 9 1 11 11 1 11 2
42 1 9 2 10 9 11 7 10 10 9 4 13 13 13 10 10 9 1 9 2 1 9 11 5 1 10 11 11 2 7 11 1 11 2 7 11 1 11 7 11 2 2
29 10 9 1 11 11 2 1 9 2 11 11 11 2 13 10 9 13 1 10 9 1 11 1 10 9 0 1 11 2
30 11 13 10 9 1 10 9 9 12 1 10 9 2 12 11 2 2 13 1 11 11 1 11 10 12 1 11 1 12 2
17 2 7 15 15 13 16 13 10 9 13 1 10 2 0 2 9 2
22 4 13 1 10 0 9 16 10 11 1 11 11 1 11 2 11 11 11 2 11 11 2
15 13 3 1 10 9 2 11 2 10 9 13 1 10 9 2
11 10 9 1 9 13 12 9 2 9 5 2
24 15 13 10 9 1 13 10 9 1 10 9 0 1 10 9 0 2 0 2 0 7 0 2 2
19 10 9 13 16 13 7 16 13 1 9 2 3 13 10 9 2 8 2 2
20 11 7 11 15 13 1 10 9 2 7 11 13 13 15 1 13 1 10 9 2
34 16 10 9 15 13 3 1 9 2 10 9 15 13 1 10 9 4 13 1 11 2 7 10 9 13 10 9 2 13 1 13 0 9 2
55 2 10 9 11 11 11 4 13 3 1 10 9 1 9 1 10 9 16 13 10 9 1 9 7 1 10 16 4 13 1 10 9 0 11 11 1 10 11 1 11 1 10 11 2 11 2 2 13 3 10 9 10 11 11 2
19 10 9 15 13 10 9 0 2 13 10 11 11 1 11 10 0 9 0 2
27 10 9 1 10 11 13 15 1 10 9 1 11 11 7 13 3 0 16 13 13 10 9 1 13 15 15 2
32 10 9 9 13 1 10 0 2 8 2 2 9 2 9 2 7 15 13 1 10 9 0 1 9 0 16 15 13 13 1 9 2
19 1 1 10 10 9 16 1 10 9 15 13 13 10 9 1 9 1 11 2
39 1 11 1 12 2 11 13 10 9 1 11 11 11 2 10 9 12 2 11 2 12 1 9 1 9 1 10 9 1 13 1 10 9 1 9 1 10 9 2
34 1 9 10 9 3 0 13 0 7 15 13 1 10 9 1 11 1 11 2 7 3 1 10 11 2 1 9 0 1 9 0 7 0 2
20 10 9 11 11 15 13 1 11 1 12 7 10 9 15 13 1 11 1 12 2
17 15 13 1 11 1 11 2 12 9 3 2 4 13 1 10 9 2
45 16 13 16 10 9 0 13 2 3 2 1 10 9 2 0 2 2 4 13 1 9 16 15 13 1 9 0 1 10 9 16 15 13 2 3 13 1 10 0 9 7 1 9 0 2
35 10 0 9 0 15 13 10 9 13 10 9 0 3 11 13 10 9 2 3 0 1 13 2 16 15 13 1 10 9 3 0 1 10 9 2
26 2 10 9 2 2 12 2 2 1 11 11 2 7 2 9 2 2 12 2 2 9 13 1 11 11 2
55 13 16 10 9 1 9 2 15 4 13 3 2 13 1 10 12 12 9 1 9 16 3 13 10 11 1 9 1 9 0 2 13 1 13 10 9 13 10 9 0 1 9 0 7 10 9 2 11 2 7 11 2 1 12 2
19 1 11 1 12 13 1 10 9 1 11 1 10 9 1 10 11 1 11 2
42 1 13 10 9 1 10 9 2 4 13 1 13 10 11 1 11 11 1 10 2 11 11 2 2 3 10 0 9 13 11 11 11 2 11 11 2 11 11 7 11 11 2
22 1 10 11 1 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 9 5 2
38 10 11 3 13 9 1 10 11 1 10 9 1 10 9 1 10 0 9 1 12 7 12 1 10 9 1 12 7 12 3 2 2 3 3 3 13 2 2
8 13 15 1 15 7 1 15 2
35 16 13 2 11 4 1 13 15 1 10 9 1 11 1 11 11 2 7 10 9 11 11 11 15 13 7 13 1 11 10 9 1 10 9 2
16 13 1 11 1 12 2 11 11 4 13 3 10 10 9 0 2
25 11 3 4 1 13 1 2 11 11 2 2 7 3 2 11 2 2 3 1 10 9 1 10 9 2
50 2 11 11 11 11 2 13 1 10 9 3 13 3 1 11 7 13 10 9 1 9 2 7 16 2 11 11 11 11 2 2 13 10 10 9 2 7 10 9 1 10 0 4 13 1 10 11 1 11 2
29 11 13 0 1 10 9 2 11 11 2 10 9 0 1 10 9 1 10 13 15 1 9 1 10 2 9 2 0 2
17 9 0 1 13 2 13 10 9 2 9 1 9 2 9 7 9 2
29 1 13 1 11 12 2 10 9 4 13 10 9 1 9 7 13 10 9 1 9 1 10 9 0 1 9 1 11 2
37 15 13 12 9 2 10 0 9 1 10 9 2 10 9 1 10 9 1 10 9 1 9 3 3 15 4 13 10 9 7 10 9 1 10 9 0 2
22 10 9 1 9 0 7 9 0 2 11 11 2 13 10 9 1 9 1 10 9 11 2
52 9 1 9 0 2 1 10 15 10 0 9 1 9 1 10 9 1 10 9 16 15 13 13 1 9 0 7 16 13 16 2 1 10 3 2 1 10 12 5 7 12 5 1 10 9 15 13 0 1 9 0 2
27 15 13 1 9 1 12 2 7 13 10 9 3 13 10 9 1 10 9 2 0 7 0 11 11 1 12 2
15 10 9 13 10 9 1 3 0 9 1 10 9 1 11 2
9 3 16 1 10 9 13 11 11 2
17 1 10 9 11 11 2 3 13 10 9 11 2 13 3 1 15 2
21 10 9 13 7 13 1 10 9 3 7 3 15 0 13 13 9 1 11 7 11 2
11 11 13 1 10 9 1 9 1 10 11 2
38 3 3 1 10 9 2 1 10 9 1 11 2 10 9 1 10 9 1 10 11 2 2 15 13 12 9 1 9 13 1 9 9 1 10 9 1 9 2
28 10 0 9 13 1 10 9 2 1 10 12 9 1 9 2 7 3 3 13 3 9 16 4 13 1 10 9 2
16 1 11 4 13 1 13 15 1 9 1 10 9 0 7 0 2
31 10 9 1 9 1 9 2 8 2 13 10 9 1 10 9 2 13 1 10 9 1 10 9 1 10 16 10 9 13 13 2
55 1 3 1 12 9 0 7 12 9 1 10 9 2 10 9 13 1 11 11 2 13 1 12 7 12 10 9 11 7 11 0 1 11 11 7 1 12 4 13 1 10 9 11 11 1 13 10 11 1 10 11 1 10 11 2
11 9 9 2 9 5 12 2 9 5 12 2
9 13 1 10 11 11 1 10 11 2
47 10 9 13 10 9 2 10 9 1 9 13 1 9 1 9 13 10 9 0 1 13 15 2 16 1 10 9 1 11 11 7 11 11 13 12 2 10 9 11 11 7 10 9 1 10 9 2
51 10 9 1 10 11 1 11 1 10 11 11 1 11 2 11 2 2 11 11 2 13 1 10 9 1 9 16 1 10 9 16 15 13 13 10 9 0 7 10 9 1 10 9 1 10 11 2 9 0 2 2
21 10 9 13 10 9 16 3 13 9 7 1 15 4 13 10 9 1 10 9 0 2
30 10 9 1 11 11 13 15 1 10 10 9 3 15 4 13 9 1 10 0 9 7 1 0 2 10 9 7 10 9 2
18 16 11 13 10 9 1 12 2 3 13 10 9 1 9 1 10 9 2
11 10 9 3 15 13 1 9 1 10 9 2
28 11 11 11 2 12 1 11 1 12 2 12 1 11 1 12 2 13 15 1 10 9 0 1 9 0 3 0 2
40 11 13 1 9 13 10 10 9 1 11 11 2 11 11 11 11 11 2 7 13 1 13 1 10 9 2 1 9 10 9 1 9 1 10 9 15 13 4 13 2
43 10 9 1 10 9 13 1 12 9 2 12 5 9 2 12 5 9 2 12 5 9 2 12 5 9 1 10 11 2 12 5 1 10 9 7 12 5 1 12 7 3 9 2
27 13 1 11 1 11 11 11 1 10 9 1 9 1 9 1 10 11 1 11 1 11 11 1 11 1 12 2
36 3 3 10 9 7 10 9 2 10 0 9 1 15 13 10 9 2 3 4 13 16 13 10 9 0 2 7 3 0 9 10 15 13 1 9 2
11 1 9 1 15 10 9 4 3 3 13 2
32 14 2 15 13 12 5 15 15 8 13 9 1 10 9 7 9 3 7 13 1 15 9 1 9 7 1 3 0 9 1 9 2
16 10 8 2 9 3 13 3 3 0 7 10 9 1 13 9 2
25 1 3 10 9 8 1 9 8 2 10 9 0 1 10 9 1 10 11 13 10 9 1 10 9 2
48 10 9 4 13 3 1 10 9 1 11 11 7 10 9 1 12 2 10 11 1 10 11 2 10 11 1 10 11 1 10 11 2 7 4 4 13 1 10 9 1 10 9 0 7 1 10 9 2
49 13 10 9 13 10 9 13 1 8 9 1 10 9 0 1 11 2 10 9 1 9 2 1 10 9 1 9 1 15 2 9 2 9 2 9 2 9 0 2 9 0 2 9 2 11 1 11 11 2
33 10 9 0 1 10 9 1 10 2 11 2 4 13 9 1 10 9 1 10 9 1 9 1 10 9 1 10 9 0 1 10 9 2
59 1 10 12 9 2 11 13 0 1 10 12 5 9 2 10 12 5 13 9 2 10 12 5 13 9 2 10 12 5 13 9 2 10 12 5 13 9 1 10 11 2 10 12 5 13 1 10 9 7 10 12 5 13 1 12 7 3 9 2
62 9 1 10 9 1 12 9 0 15 4 13 10 9 0 1 10 16 1 9 1 10 9 11 11 9 1 10 9 2 9 7 9 15 13 7 13 1 10 9 1 9 1 11 1 13 15 7 13 10 9 7 10 9 16 13 10 9 7 10 9 0 2
25 13 1 10 11 0 2 2 11 7 11 2 13 10 9 0 1 12 9 2 11 11 7 11 11 2
38 3 2 10 9 11 11 11 2 11 11 2 2 16 13 10 11 1 11 11 1 10 11 1 11 2 13 10 9 1 10 9 1 4 1 13 10 9 2
24 3 1 10 9 1 10 9 11 1 9 1 10 9 12 3 13 9 10 9 1 9 7 9 2
16 10 0 9 15 13 1 10 9 0 1 10 9 1 10 9 2
26 11 1 10 11 11 2 11 2 11 12 1 11 1 12 2 2 9 0 2 3 9 11 11 1 11 2
20 15 4 13 1 10 9 0 1 9 0 1 10 9 7 4 13 9 1 9 2
6 15 13 1 10 9 2
11 10 11 7 11 3 4 13 1 9 0 2
54 13 0 9 2 1 15 10 9 1 11 13 1 12 1 11 11 10 11 1 10 9 1 11 11 12 2 7 10 9 1 9 1 11 16 13 9 1 12 13 1 11 12 1 11 2 16 13 9 1 10 9 1 11 2
19 1 9 2 1 10 9 10 9 13 0 2 16 13 10 9 1 10 9 2
17 1 10 0 9 13 10 9 1 9 7 9 1 10 11 1 11 2
32 11 13 12 9 7 11 7 11 12 10 15 2 15 16 13 1 10 9 1 10 9 0 1 10 11 11 16 15 13 1 12 2
38 15 13 9 1 9 0 2 9 0 7 9 2 9 16 3 1 10 0 9 1 11 11 1 10 11 4 3 13 1 10 9 1 10 9 1 10 9 2
13 3 13 1 10 9 1 0 1 9 1 12 9 2
23 10 9 1 10 9 1 11 2 1 9 2 8 8 2 4 13 10 12 1 11 1 12 2
10 11 11 2 12 2 13 10 9 0 2
41 10 9 3 0 3 1 9 1 3 16 10 9 3 10 9 13 10 9 2 10 9 0 2 13 16 13 9 7 13 10 9 2 7 10 9 1 9 0 7 0 2
8 2 3 13 10 9 1 15 2
43 10 9 0 13 10 2 9 2 11 11 1 9 0 2 0 1 13 1 9 1 10 9 7 10 9 2 13 10 9 2 7 13 1 10 9 0 2 13 1 10 11 11 2
63 1 10 12 9 2 10 9 1 11 11 4 13 1 10 12 5 0 2 10 12 5 13 0 2 10 12 5 13 9 2 10 12 5 13 0 2 10 12 5 13 0 1 10 11 2 10 12 5 13 1 10 9 7 10 12 5 13 1 12 7 3 9 2
15 11 2 2 15 13 15 16 3 15 13 13 1 10 9 2
10 15 13 1 10 9 11 2 11 2 2
26 15 13 10 9 1 10 9 1 10 9 12 2 7 3 3 15 4 4 13 1 9 1 10 9 12 2
20 10 9 0 4 13 1 10 0 11 1 9 1 10 9 11 11 2 12 2 2
24 13 1 9 7 10 0 9 13 10 11 11 1 11 2 8 2 1 10 0 9 8 1 11 2
30 10 9 1 11 2 1 9 2 11 11 2 13 10 9 13 1 10 9 1 11 1 10 9 0 1 11 1 10 11 2
31 1 12 13 10 9 1 10 9 13 1 10 11 11 1 11 1 10 2 9 2 9 1 10 9 13 15 1 10 11 0 2
24 10 9 1 9 13 10 9 0 1 10 11 0 2 1 10 11 0 2 11 2 11 7 11 2
21 10 9 0 1 10 9 13 2 11 7 11 11 1 10 11 7 10 9 0 2 2
43 10 9 4 13 1 11 11 1 10 11 2 1 11 1 10 12 5 1 10 12 5 9 1 11 11 7 1 10 12 5 9 1 11 11 7 1 11 1 11 11 7 11 2
41 10 9 15 13 1 10 9 0 1 10 11 2 13 1 9 1 10 9 2 16 13 9 3 0 1 10 9 1 9 7 9 1 10 0 9 1 9 1 10 11 2
50 1 10 9 0 2 10 9 15 13 1 0 1 9 7 9 2 1 9 0 1 10 9 7 10 11 0 2 7 15 13 1 9 1 9 13 1 9 2 15 16 15 13 10 9 0 1 10 11 0 2
18 10 9 7 0 9 13 0 1 10 9 1 10 9 1 10 11 11 2
9 11 11 15 13 13 1 10 9 2
34 13 1 11 11 2 1 10 9 15 13 10 9 1 10 9 2 10 9 1 10 9 1 10 9 7 10 9 1 10 9 1 10 9 2
60 10 0 12 1 11 2 1 10 9 1 11 1 11 2 10 9 11 11 13 9 1 10 9 1 11 7 11 11 1 11 11 2 10 9 3 13 0 2 7 13 2 2 4 3 13 15 1 10 11 3 4 1 13 10 9 1 10 9 2 2
17 15 13 1 10 11 11 12 2 1 12 9 1 10 9 1 11 2
15 1 12 4 13 9 1 10 9 7 1 12 9 1 11 2
16 1 15 15 2 13 0 16 11 15 13 3 3 1 12 3 2
34 1 10 9 1 10 9 2 15 13 1 13 9 2 13 15 1 10 9 2 2 10 9 0 15 13 3 1 15 7 1 10 9 2 2
15 11 11 3 4 13 3 9 7 15 16 15 13 10 9 2
9 15 4 13 1 10 9 16 13 2
15 10 9 13 11 11 2 11 11 2 11 11 7 11 11 2
21 11 13 1 10 2 9 1 9 2 2 11 11 2 2 1 9 0 1 9 0 2
23 1 10 12 15 3 1 10 9 2 12 5 2 1 10 9 1 9 1 13 15 13 3 2
26 10 9 0 1 11 13 13 15 1 11 16 10 9 13 15 15 16 4 13 1 10 9 1 10 9 2
17 15 1 10 0 9 1 10 9 13 10 9 1 9 1 10 9 2
19 10 9 13 3 0 1 15 1 10 9 11 2 13 0 1 15 1 11 2
25 11 2 11 11 2 13 10 0 9 1 9 1 10 9 0 1 9 0 11 11 11 13 1 12 2
36 10 9 13 13 10 9 1 10 9 1 10 9 7 2 1 9 2 13 10 0 9 1 9 1 10 9 7 10 9 0 7 10 9 1 9 2
41 13 16 13 1 10 9 1 10 9 0 1 11 7 1 11 2 7 13 3 7 3 16 13 10 11 11 7 13 11 7 10 9 1 10 11 1 11 1 15 13 2
33 3 13 9 0 1 9 0 1 9 1 11 2 11 2 11 2 11 11 2 11 2 11 2 11 11 2 7 10 9 0 1 11 2
12 11 13 10 9 1 9 0 1 10 9 11 2
31 1 12 13 9 0 1 11 11 11 7 1 10 9 0 13 1 10 9 7 15 13 1 10 11 11 1 11 7 11 11 2
8 9 2 13 0 10 9 2 2
34 3 13 10 9 1 9 13 1 10 9 11 11 7 10 2 11 11 2 2 15 16 15 13 13 1 11 7 13 10 0 9 1 11 2
26 1 10 9 13 10 9 0 16 15 9 2 1 10 9 13 10 9 0 7 9 1 10 15 13 0 2
57 10 9 15 13 1 9 2 10 9 1 9 3 0 1 10 9 1 9 1 11 7 11 13 1 10 0 11 0 2 10 9 0 3 0 13 1 10 9 1 10 11 1 9 1 10 11 2 3 1 10 9 1 11 1 12 2 2
10 9 13 1 9 7 9 1 0 9 2
25 10 0 9 1 10 11 11 4 13 10 12 1 11 1 10 12 1 10 11 8 11 11 1 11 2
22 1 12 2 10 9 2 15 11 11 2 15 13 1 15 3 0 1 10 9 1 9 2
51 15 13 3 1 10 9 0 1 10 9 7 13 1 10 9 1 10 9 1 10 3 9 1 10 11 2 11 11 11 2 15 13 13 0 9 1 9 13 15 1 11 11 2 9 1 11 11 1 10 9 2
10 15 13 1 9 1 10 9 1 11 2
33 13 10 0 9 1 11 1 10 9 0 2 1 10 15 13 1 9 1 12 2 7 1 10 9 2 16 13 1 13 10 0 9 2
15 10 9 7 10 9 4 13 10 9 1 10 9 0 11 2
13 10 9 0 4 13 15 16 4 0 1 11 11 2
12 10 9 1 9 1 10 9 13 1 5 12 2
9 11 11 11 13 10 9 0 0 2
27 10 9 1 10 9 11 4 3 13 1 10 9 1 9 9 1 11 11 2 11 2 9 1 11 11 2 2
24 15 13 10 9 1 10 11 11 11 2 10 9 0 16 13 1 10 9 7 15 1 9 0 2
20 10 9 1 10 9 7 10 9 13 2 16 13 1 13 2 13 10 9 0 2
40 1 10 9 0 2 11 2 10 9 1 10 15 13 10 11 0 2 2 3 1 10 9 13 2 13 13 1 15 2 7 11 13 10 9 0 1 13 15 13 2
23 4 13 12 5 1 10 9 1 11 7 12 1 10 9 1 11 2 10 9 1 10 9 2
15 10 9 4 3 13 7 13 1 10 10 9 1 10 9 2
45 10 9 16 4 13 1 13 12 9 11 2 10 0 7 3 0 9 1 9 1 10 9 2 13 3 9 3 7 13 10 9 16 15 13 1 9 1 10 9 1 9 1 0 9 2
10 7 1 10 0 9 3 13 10 9 2
33 15 4 1 13 1 10 9 2 3 1 4 13 16 10 9 13 1 10 9 7 2 3 0 2 13 1 10 9 1 10 9 0 2
57 3 2 11 13 1 16 10 9 1 10 11 1 11 2 11 11 2 13 3 10 2 9 0 2 1 10 9 0 0 1 10 9 16 13 1 10 9 1 9 1 11 7 11 2 1 10 16 10 2 9 2 13 10 9 1 9 2
25 10 9 9 1 11 2 11 11 2 2 1 9 2 13 10 9 1 9 1 9 1 10 11 11 2
28 13 10 9 0 1 11 11 7 1 11 11 2 16 15 4 13 10 9 0 16 13 10 9 1 12 1 11 2
52 1 9 2 10 9 2 1 9 2 9 2 13 10 9 1 10 15 10 9 16 13 10 9 0 2 4 3 13 7 4 1 13 2 1 10 9 2 1 16 13 1 10 9 1 9 1 10 9 1 10 9 2
23 10 9 4 13 1 0 9 1 11 2 7 3 3 1 11 1 10 11 2 11 7 11 2
29 10 0 9 1 10 9 13 10 9 1 9 0 1 10 9 1 9 1 10 11 1 10 11 7 10 11 1 11 2
27 10 9 15 13 1 0 9 15 1 10 9 0 13 10 9 2 7 16 1 10 9 15 13 10 9 0 2
19 13 1 10 9 1 10 11 10 12 1 11 1 10 9 1 10 11 11 2
10 10 9 13 1 10 9 12 1 9 2
17 10 9 7 0 9 1 9 1 10 9 1 10 9 13 10 9 2
21 0 1 10 9 13 10 9 1 9 1 12 9 1 10 9 1 9 9 0 11 2
14 13 1 10 11 2 11 2 10 12 1 11 1 12 2
14 15 13 1 10 9 0 10 12 9 1 13 10 9 2
82 11 11 11 2 11 7 11 2 9 2 8 8 8 2 13 10 12 1 11 1 12 1 11 2 11 11 2 2 13 10 9 1 10 11 1 11 1 10 11 2 11 2 16 4 1 13 9 0 2 8 2 1 10 9 1 10 11 1 11 2 7 16 4 13 1 10 11 11 2 13 15 1 10 9 1 3 0 9 1 10 9 2
24 10 9 13 1 10 9 1 9 1 10 9 1 10 11 11 16 13 1 10 9 0 3 0 2
29 10 0 9 16 13 10 12 1 11 1 12 13 10 9 0 7 13 0 9 1 10 9 1 10 9 1 9 0 2
67 3 15 13 10 9 1 10 11 2 9 11 11 11 2 15 13 16 13 10 9 10 9 2 13 1 10 9 1 9 0 2 7 10 8 8 13 13 1 10 9 7 13 1 10 9 1 13 15 1 10 9 3 13 10 9 7 1 10 9 13 1 9 16 13 10 9 2
18 4 13 1 0 1 10 11 11 11 1 12 1 10 9 1 11 11 2
30 4 13 9 1 0 9 1 10 9 2 1 10 13 9 1 15 13 10 9 16 13 1 10 9 2 13 10 9 0 2
22 1 10 9 1 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 5 5 2
21 3 4 13 1 11 11 2 10 0 9 1 11 11 2 1 10 0 9 11 11 2
18 15 9 13 13 9 0 1 10 9 1 9 2 9 0 7 10 9 2
55 1 9 2 1 9 1 10 9 1 9 15 15 13 16 13 10 9 2 13 10 9 1 16 2 1 10 9 1 10 12 9 2 10 0 9 4 4 13 3 10 9 4 13 3 13 2 15 13 2 3 3 1 10 11 2
40 4 13 1 10 0 9 1 10 9 1 11 11 2 10 9 13 0 16 13 10 9 2 7 15 13 1 9 3 0 7 13 1 10 9 1 9 1 10 9 2
12 1 10 0 9 2 11 13 13 10 9 0 2
18 10 9 13 1 10 1 10 11 1 10 15 11 15 13 13 1 11 2
5 9 1 9 0 2
12 10 11 11 2 13 10 9 13 1 11 11 2
50 10 9 0 13 1 10 9 1 10 11 1 11 4 13 3 1 10 9 0 2 9 7 9 2 7 1 10 9 0 2 9 2 2 16 3 4 13 10 9 13 1 1 10 9 0 2 9 9 2 2
34 10 0 9 1 10 9 15 13 1 10 9 1 9 0 7 0 2 3 7 1 10 0 9 1 0 9 0 1 10 9 1 10 9 2
20 13 12 9 1 9 1 10 9 0 1 11 2 9 1 9 3 13 7 13 2
15 10 9 0 15 13 3 13 1 9 13 10 9 0 13 2
31 1 15 13 9 2 11 11 2 2 10 9 0 16 1 10 9 13 1 10 9 1 11 2 7 16 1 9 13 1 11 2
17 13 10 12 9 1 9 0 0 2 9 1 12 9 7 9 0 2
18 1 15 9 16 3 13 9 1 10 9 10 9 15 13 1 10 9 2
26 10 9 1 11 15 11 13 3 0 2 7 10 9 8 1 10 9 3 13 15 9 1 10 0 9 2
21 10 9 1 10 9 13 10 9 2 10 9 2 10 9 2 10 9 7 10 9 2
43 10 9 13 1 10 9 12 1 10 9 1 9 7 9 0 13 1 10 9 1 10 11 2 1 10 9 1 9 1 12 1 10 9 0 11 11 7 1 11 1 11 2 2
18 13 9 7 9 1 10 11 11 1 11 1 9 7 9 1 10 9 2
25 10 9 13 16 10 9 0 4 13 1 3 1 12 9 1 9 1 10 9 3 0 1 10 10 9
32 13 15 1 10 9 1 9 0 2 8 2 1 11 2 16 1 10 9 10 8 2 8 13 15 3 7 10 9 9 1 9 2
26 10 9 13 12 9 1 9 2 7 10 9 1 11 13 3 3 3 9 13 7 10 11 3 15 13 2
25 10 9 13 10 12 1 11 2 13 1 0 9 7 11 0 1 9 0 2 16 13 0 1 9 2
12 15 13 1 11 13 1 10 11 11 1 11 2
41 10 9 0 1 9 13 10 9 1 11 11 2 16 1 10 9 1 10 9 13 16 10 11 3 4 13 1 13 3 0 1 16 13 0 1 10 10 9 0 0 2
7 1 15 13 10 9 11 2
17 15 13 1 10 9 1 11 2 10 11 2 1 10 11 1 11 2
43 1 15 15 16 15 13 13 16 15 13 10 10 9 2 16 13 15 13 10 9 7 10 9 16 13 1 11 11 2 1 10 9 7 1 10 9 1 10 9 1 10 9 2
22 1 10 9 1 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 5 5 2
13 3 12 9 0 15 13 1 13 10 12 0 9 2
29 1 10 9 2 10 9 13 0 1 10 9 3 0 7 0 7 1 15 1 15 16 13 3 10 9 1 9 0 2
27 10 12 1 11 1 12 2 11 11 4 13 1 0 9 1 10 9 11 11 1 10 9 12 3 1 11 2
37 11 7 11 11 1 11 7 11 2 10 0 9 1 11 1 11 2 7 10 11 11 11 11 11 11 11 1 10 12 1 11 7 10 12 1 11 2
23 10 9 0 7 1 9 4 4 13 1 11 11 11 2 11 11 2 11 11 7 11 11 2
19 13 9 1 9 0 2 9 1 9 2 11 2 9 7 9 0 1 9 2
38 11 11 13 10 9 3 0 2 12 9 1 9 2 10 15 13 10 11 11 3 1 10 9 1 11 1 10 11 16 13 16 3 15 13 1 10 9 2
24 10 9 13 16 10 9 1 10 9 1 10 10 11 4 13 1 10 9 0 1 12 11 11 2
24 1 10 9 2 9 0 2 2 13 10 9 1 9 16 13 1 9 7 15 13 1 10 9 2
34 10 11 13 10 9 0 13 1 9 1 10 9 12 1 9 1 10 9 1 9 1 10 9 0 5 2 12 1 10 9 1 10 11 2
39 16 10 11 1 11 13 3 3 16 11 4 3 13 1 10 9 2 10 9 13 1 11 2 13 16 13 10 9 1 13 0 9 1 9 1 9 7 11 2
21 10 9 15 13 3 1 10 9 1 9 2 10 0 9 1 10 9 1 10 9 2
19 10 0 9 13 1 13 15 1 9 1 10 9 16 1 15 4 13 15 2
13 1 10 9 1 12 2 13 12 9 13 1 11 2
15 3 13 10 9 0 7 15 7 10 9 3 15 4 13 2
21 1 9 3 13 10 9 1 10 9 2 7 3 1 12 15 13 13 10 9 0 2
27 11 11 13 10 9 0 2 2 13 10 12 1 11 1 12 1 11 2 16 13 1 10 9 0 11 11 2
10 1 15 15 13 1 10 9 10 9 2
39 10 11 11 2 7 3 9 2 13 10 9 0 13 1 11 2 1 10 9 1 11 11 2 12 2 2 1 10 9 1 13 10 0 9 0 1 10 11 2
16 1 9 1 10 9 10 12 5 13 0 7 9 1 10 9 2
25 7 2 1 9 2 10 9 1 10 9 13 16 10 9 13 0 1 10 9 1 3 13 10 9 2
46 3 10 9 11 3 15 13 1 2 9 2 7 2 9 1 10 9 2 7 13 13 10 9 1 9 1 9 0 3 16 13 3 0 1 10 9 1 10 9 2 3 1 10 9 11 2
32 4 13 1 10 9 1 10 0 9 0 1 11 7 1 10 9 0 1 11 2 1 10 9 3 13 10 9 1 10 9 0 2
32 13 10 9 16 15 13 1 10 9 0 1 11 11 11 1 10 9 1 13 10 9 16 3 13 10 9 1 13 1 10 9 2
31 10 9 0 1 11 13 1 0 9 0 3 7 13 13 10 10 9 1 9 2 0 1 9 7 0 2 0 7 0 2 2
42 16 10 9 13 3 1 9 1 10 0 9 2 10 9 1 11 13 9 0 2 7 3 1 9 1 13 1 10 9 2 13 15 16 13 1 10 9 16 3 4 13 2
18 1 10 9 10 9 0 4 1 13 13 10 9 0 1 9 1 11 2
25 1 15 15 13 3 10 9 1 9 7 10 9 16 15 13 1 11 2 11 2 11 11 7 11 2
15 3 10 9 13 1 11 11 2 4 13 1 10 9 0 2
24 11 13 10 0 9 1 9 16 13 9 1 9 0 1 10 9 2 10 9 2 11 11 2 2
25 10 9 0 1 9 13 16 1 11 1 3 12 9 15 4 13 13 10 9 1 10 0 12 5 2
24 13 1 11 2 11 7 15 13 1 11 2 11 2 16 15 13 1 10 9 0 1 10 9 2
10 4 13 9 10 12 1 11 1 12 2
5 11 13 1 11 2
13 13 1 13 1 9 2 4 13 1 9 1 12 2
67 1 9 2 1 10 11 11 1 10 11 1 12 2 11 11 11 2 11 11 7 11 11 13 1 10 9 1 10 9 0 1 10 0 9 1 11 1 10 9 2 7 15 13 16 11 4 13 10 9 7 3 13 10 9 1 10 11 1 10 9 0 1 9 1 11 11 2
9 13 9 7 9 2 13 9 2 2
18 13 7 9 2 11 11 1 10 9 1 11 2 11 7 11 2 11 2
21 15 3 13 0 9 2 13 15 3 0 2 11 1 10 9 7 11 1 10 9 2
24 10 9 0 12 9 1 11 1 11 2 11 2 13 1 11 2 11 2 11 2 11 7 11 2
51 13 12 5 2 12 9 2 1 0 2 12 5 2 12 9 2 1 9 7 10 9 9 1 12 5 2 12 9 2 1 10 9 1 10 9 2 2 12 5 7 12 9 1 3 1 10 11 1 11 2 2
32 13 1 10 11 1 11 2 3 1 11 11 2 10 12 1 11 1 12 2 9 1 10 0 1 10 9 16 13 0 1 9 2
24 10 9 1 10 10 11 11 13 10 9 3 2 0 9 15 13 7 13 9 1 10 9 2 2
46 10 9 1 10 9 0 1 10 9 1 10 9 13 16 1 10 12 1 10 9 1 10 11 2 3 1 4 13 3 10 9 2 10 9 13 1 10 9 7 13 16 15 13 12 9 2
38 10 9 13 0 2 13 13 2 16 3 13 3 1 10 9 0 2 7 1 10 10 9 7 2 3 2 13 1 9 0 16 13 15 9 1 15 9 2
5 15 13 1 12 2
14 10 9 13 1 10 9 13 10 12 5 1 10 9 2
14 11 13 3 10 9 1 10 9 1 10 0 9 0 2
8 13 10 0 9 1 15 2 2
15 15 13 10 9 1 9 2 10 9 2 10 9 1 9 2
15 10 3 2 9 13 3 0 1 10 9 1 8 8 11 2
13 10 9 1 10 9 1 10 9 4 13 1 11 2
41 1 9 2 10 9 13 0 1 9 0 3 0 2 7 1 11 2 10 9 0 16 13 10 9 16 15 15 13 10 9 1 10 9 7 1 10 9 1 10 9 2
13 10 9 13 3 15 1 15 16 13 0 9 0 2
19 13 12 9 2 11 2 11 2 11 2 11 1 10 11 2 11 7 11 2
12 10 9 13 10 9 10 12 1 11 1 12 2
14 11 13 9 1 10 9 1 9 1 10 9 11 11 2
23 10 11 13 10 9 0 1 10 9 0 2 11 1 11 11 2 9 1 11 11 2 11 2
30 10 9 1 9 1 10 9 0 13 1 10 12 1 10 12 9 2 7 16 15 1 10 9 13 1 10 12 7 12 2
14 1 9 2 11 4 13 1 13 0 9 0 1 11 2
28 13 1 10 9 0 11 11 2 15 16 13 2 13 0 7 13 0 13 1 10 9 10 9 16 13 10 9 2
9 11 13 9 1 10 11 1 11 2
43 11 13 10 0 9 1 10 9 1 10 11 10 12 1 11 2 13 1 10 9 1 10 0 9 1 10 11 1 11 2 9 1 12 9 1 10 9 7 10 9 1 9 2
15 3 15 13 11 11 11 2 7 11 2 7 10 11 11 2
28 10 9 0 1 11 2 1 15 3 1 12 5 1 10 9 2 13 0 1 13 9 1 10 9 0 7 9 2
39 10 9 0 0 13 11 1 10 9 2 11 1 10 9 7 9 2 11 1 10 9 2 13 1 10 9 7 10 9 2 7 10 9 1 11 1 10 9 2
14 3 2 11 13 10 9 1 11 2 7 4 13 9 2
23 3 1 9 2 15 4 13 16 10 9 1 11 3 4 13 3 1 11 0 7 9 0 2
18 13 10 9 0 16 15 13 1 15 1 10 9 3 0 1 10 9 2
28 2 3 13 0 16 16 15 13 7 13 13 1 13 15 10 9 12 9 0 7 1 10 9 13 1 12 9 2
34 3 10 9 13 10 0 9 1 10 9 1 10 11 1 10 11 2 1 10 9 15 13 1 10 9 10 0 9 11 11 2 11 2 2
33 10 9 4 13 10 9 1 9 0 2 7 0 1 11 2 1 9 2 10 9 0 1 11 2 7 10 9 0 1 10 9 2 2
30 3 15 13 0 13 10 9 13 15 2 16 3 0 15 13 13 1 10 9 1 9 9 0 1 9 7 9 10 9 2
45 1 10 9 2 13 16 10 9 1 10 9 2 1 9 1 9 7 1 10 9 2 3 0 2 2 13 1 10 9 1 10 9 1 10 9 16 2 13 10 9 1 10 9 2 2
20 3 13 1 11 2 1 15 10 9 1 11 13 10 9 1 9 1 10 12 2
25 11 13 10 0 9 1 10 11 11 1 12 9 5 16 15 13 1 11 2 11 2 11 7 11 2
40 1 11 13 10 9 1 11 11 2 1 10 9 0 7 3 13 1 9 10 9 1 10 9 1 10 11 2 16 15 13 1 10 15 2 10 9 1 10 11 2
21 1 10 9 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 9 5 2
37 10 9 13 10 9 7 10 9 1 9 1 10 11 11 2 10 9 1 9 2 10 9 1 9 7 9 0 2 3 7 1 10 9 1 9 0 2
32 10 9 12 11 2 1 9 2 11 12 2 11 2 13 10 9 13 1 10 9 1 11 1 10 9 0 1 11 1 10 11 2
36 10 9 13 13 1 10 9 0 1 12 8 1 0 2 12 8 1 0 7 12 8 1 9 2 1 10 9 0 0 1 10 9 1 12 9 2
16 3 2 16 10 9 13 10 9 0 2 15 4 7 13 0 2
37 10 9 3 0 7 1 10 9 13 1 9 1 3 1 12 9 2 7 1 3 9 13 1 10 0 9 1 10 0 9 1 10 9 1 10 9 2
13 13 13 1 10 9 2 15 15 13 1 9 9 2
33 13 13 15 16 1 10 0 9 1 10 9 0 1 10 11 11 2 3 13 10 9 0 1 11 16 13 0 10 9 1 10 9 2
25 13 1 10 9 16 15 13 7 15 1 12 9 13 10 9 2 15 13 2 15 15 13 3 3 2
14 13 13 16 10 11 11 13 10 9 0 1 9 0 2
19 10 9 0 1 9 0 1 10 9 1 10 9 0 13 10 9 3 0 2
7 13 1 9 12 9 0 2
16 11 1 11 11 2 11 1 11 2 12 1 11 1 12 2 2
35 10 11 13 3 1 10 9 1 9 0 0 2 13 3 16 10 9 2 0 2 3 4 13 15 1 10 9 16 15 13 1 10 9 0 2
40 3 16 3 1 10 9 1 9 10 9 13 1 9 2 13 1 9 9 0 7 0 2 11 13 1 10 9 10 15 1 10 12 9 2 13 10 9 3 0 2
29 15 13 1 10 9 1 9 1 11 2 13 7 15 13 3 1 10 9 0 16 13 0 2 3 4 13 1 9 2
14 16 10 9 3 13 13 16 3 13 9 1 10 9 2
20 3 13 9 1 11 11 2 10 9 15 13 1 10 9 0 2 7 1 11 2
35 10 9 13 10 9 0 7 0 1 10 9 0 2 7 3 0 2 1 9 2 3 16 1 11 15 13 12 9 0 1 9 1 10 9 2
27 13 10 9 1 10 9 11 11 11 7 9 1 10 9 11 11 11 2 9 1 10 9 0 1 11 2 2
13 10 9 3 3 11 13 2 2 7 10 12 9 2
31 1 10 9 1 10 9 1 12 10 9 0 1 9 1 10 9 13 1 5 12 2 7 10 9 0 1 9 13 5 12 2
21 11 4 1 13 1 11 1 10 9 1 11 2 1 12 2 1 15 1 10 9 2
23 11 11 13 10 9 7 10 9 13 10 9 0 1 9 0 7 9 0 1 10 10 9 2
15 13 1 9 1 10 9 0 1 10 11 1 10 11 11 2
13 2 9 8 8 8 1 10 9 1 10 11 2 2
8 10 11 0 13 0 7 0 2
43 13 3 1 12 9 0 2 12 1 10 9 12 2 2 10 9 13 9 2 1 10 9 1 10 9 1 10 9 0 1 11 2 7 7 10 9 1 9 13 3 10 9 2
11 10 9 1 11 15 13 13 1 10 9 2
22 10 12 9 1 11 1 9 0 13 1 10 0 9 7 13 3 1 12 9 1 9 2
35 10 9 0 13 13 16 11 13 1 11 1 13 15 1 10 9 1 9 1 9 1 10 9 15 15 13 2 7 11 15 13 1 13 15 2
17 1 12 13 12 9 2 9 2 2 12 1 12 7 12 1 12 2
38 13 0 16 10 9 1 10 9 4 7 13 1 10 11 2 7 13 3 16 15 13 10 9 16 3 4 13 1 10 9 1 10 11 1 10 10 9 2
12 10 0 9 1 9 13 10 9 8 2 8 2
27 11 11 2 13 10 12 1 11 1 12 1 11 2 11 2 11 11 2 13 10 9 9 7 9 0 0 2
12 15 13 1 10 9 0 3 1 10 9 0 2
59 1 10 12 9 2 11 13 0 1 10 12 5 0 2 10 12 5 13 0 2 10 12 5 13 0 2 10 12 5 13 0 2 10 12 5 13 0 1 10 11 2 10 12 5 13 1 10 9 7 10 12 5 13 1 12 7 3 9 2
14 13 16 10 9 1 10 9 3 13 1 10 9 13 2
24 12 9 0 2 1 10 9 1 15 13 0 2 15 13 1 10 9 1 10 9 1 10 9 2
44 10 12 9 13 0 9 0 2 7 13 3 0 16 3 10 9 0 1 10 9 1 10 9 1 10 9 1 9 7 10 9 1 10 0 9 1 10 9 0 0 15 13 13 2
11 13 16 10 9 0 4 13 1 9 0 2
48 1 12 2 10 9 0 1 11 13 10 11 12 2 10 9 1 9 16 13 10 9 1 10 10 9 1 10 9 0 2 7 16 15 13 1 9 1 10 9 1 10 11 1 10 11 1 11 2
55 13 10 12 1 11 1 12 1 10 11 2 11 11 2 11 13 1 10 11 11 1 11 7 3 10 11 11 2 8 11 2 3 13 10 9 1 11 1 12 2 10 9 1 11 1 12 2 7 10 9 1 11 1 12 2
58 4 13 1 10 9 1 10 9 2 10 9 1 9 7 10 9 2 3 7 1 10 9 1 10 9 2 13 10 9 0 2 10 9 2 10 9 2 10 9 2 10 9 2 10 9 1 9 2 10 9 2 10 9 0 7 10 9 2
16 13 1 13 1 10 9 10 9 0 1 10 9 1 9 0 2
31 1 12 2 4 13 0 9 1 10 9 1 9 1 10 3 0 2 11 11 11 0 2 2 10 9 15 13 1 12 9 2
29 1 9 2 1 10 9 1 11 2 11 9 12 13 10 9 0 15 13 12 15 13 1 10 0 9 7 15 13 2
29 10 9 1 9 0 13 10 9 1 13 2 10 9 1 10 9 1 10 9 2 7 3 10 2 9 1 13 2 2
28 10 9 1 9 0 13 10 9 1 9 1 15 9 1 10 9 16 13 13 1 10 9 13 1 10 9 0 2
47 11 13 16 3 13 13 10 9 1 9 7 13 1 15 2 7 10 0 9 13 15 16 15 13 1 10 12 9 2 13 1 15 9 1 12 9 1 12 9 0 1 10 9 1 10 11 2
20 15 1 10 9 3 0 16 10 11 11 11 11 2 13 13 10 9 11 11 2
17 11 15 13 3 10 9 1 10 9 7 11 2 10 1 10 9 2
15 15 13 15 16 4 13 10 9 1 10 9 2 1 9 2
20 1 12 13 1 11 1 10 4 13 11 1 10 9 1 10 9 0 1 11 2
55 1 3 12 9 4 13 1 9 1 10 9 1 9 13 10 11 1 11 1 10 11 1 10 9 1 11 2 9 1 9 13 1 10 9 1 10 9 9 1 10 9 2 1 10 0 9 0 13 1 10 9 1 9 11 2
39 3 4 13 9 1 9 1 13 10 0 9 16 13 13 10 9 2 15 16 13 10 9 1 9 1 10 16 15 7 15 15 13 13 1 10 9 16 13 2
29 10 9 15 13 1 10 9 1 9 1 9 1 10 9 2 3 16 13 15 1 9 1 9 2 1 9 1 9 2
17 0 1 10 9 11 2 13 1 10 9 1 10 0 9 1 11 2
18 10 9 0 3 15 13 1 3 1 10 12 5 1 10 9 0 0 2
30 10 9 1 9 1 9 7 9 1 11 13 10 9 0 1 10 9 0 7 10 9 1 9 13 3 1 10 9 0 2
24 13 3 15 1 10 9 3 0 1 13 10 9 1 11 7 10 1 11 11 2 3 1 11 2
12 11 11 13 10 9 1 9 1 10 9 11 2
9 3 4 13 3 0 1 10 9 2
24 16 1 10 9 8 2 8 5 12 2 1 9 11 13 10 9 9 1 9 1 8 5 12 2
14 11 15 13 1 10 0 9 0 16 13 10 0 9 2
29 16 15 13 13 10 9 2 10 9 7 10 9 2 3 13 7 13 15 15 1 10 11 11 16 15 13 3 0 2
20 10 11 11 11 1 11 13 10 9 1 9 0 16 13 1 10 0 9 0 2
62 10 9 2 13 1 10 9 0 2 4 13 1 10 9 11 11 11 2 1 10 9 0 1 10 9 11 11 11 2 15 13 1 2 10 9 1 10 9 1 10 9 1 9 0 2 11 11 2 1 13 1 15 9 1 9 16 13 9 1 9 2 2
31 1 10 9 2 10 9 13 1 10 0 9 0 16 13 13 1 10 0 9 1 10 9 0 7 10 9 1 10 9 11 2
12 10 9 0 13 3 3 10 9 1 10 9 2
21 10 9 4 13 15 3 7 12 9 2 16 13 1 13 10 9 1 10 9 0 2
37 13 13 10 9 0 1 10 11 11 2 0 9 1 10 11 11 3 0 1 10 9 11 7 1 3 1 12 9 1 9 7 0 1 9 1 9 2
30 11 7 11 2 3 11 13 10 9 1 10 9 0 2 10 0 9 13 13 1 10 11 7 13 1 10 9 0 11 2
33 10 9 15 4 13 1 12 9 13 1 10 9 1 9 1 9 1 11 7 11 1 10 12 0 1 10 0 9 1 10 11 11 2
32 13 1 10 11 11 2 1 0 9 1 11 2 15 13 10 9 11 2 10 0 9 1 9 0 0 1 10 9 1 9 11 2
34 13 1 10 0 9 0 1 10 11 11 7 13 1 10 9 1 11 7 11 7 11 2 11 2 15 0 9 1 10 9 1 15 13 2
34 11 13 10 9 1 9 0 13 1 10 11 11 2 1 0 9 1 11 7 11 2 1 10 11 11 2 1 10 9 1 10 11 11 2
10 1 10 9 1 13 15 13 10 9 2
39 1 10 9 0 2 10 9 9 13 3 1 10 12 5 1 10 9 1 10 9 2 12 5 1 15 1 10 9 0 7 12 5 1 15 1 10 9 0 2
7 13 10 9 1 11 7 8
27 3 16 8 4 1 10 9 2 11 13 1 10 11 1 10 9 16 13 10 9 1 10 9 7 15 13 2
16 1 9 1 13 0 1 10 9 0 2 13 10 9 3 0 2
18 10 9 4 13 3 1 10 9 2 3 7 10 9 13 1 10 9 2
29 1 9 1 10 9 2 10 11 2 13 10 9 1 10 13 15 1 10 9 1 9 3 13 10 9 1 11 11 2
31 3 13 3 3 12 9 2 11 2 11 7 11 2 13 1 10 9 10 9 13 1 15 16 3 15 13 9 1 10 11 2
60 10 9 13 16 10 9 4 13 15 1 10 9 1 9 12 2 13 10 0 9 16 13 10 9 2 1 12 9 1 9 2 13 15 10 9 1 12 9 2 12 9 2 1 11 2 11 2 1 10 9 1 12 9 2 5 2 12 8 2 2
63 2 1 9 2 10 9 1 9 1 11 11 2 11 2 1 10 9 1 9 2 4 13 1 16 2 15 4 1 13 10 9 2 16 13 10 9 1 9 1 9 0 1 11 2 1 15 15 10 9 2 4 13 3 1 10 9 2 2 4 13 10 9 2
5 9 0 1 11 2
12 1 9 0 2 13 1 10 9 1 9 13 2
27 13 10 0 9 2 3 0 1 15 13 13 10 9 7 13 10 9 0 1 11 2 10 9 7 10 9 2
39 2 10 11 1 10 11 2 2 16 15 13 11 1 10 9 2 4 3 13 1 10 9 1 10 9 3 10 0 11 13 9 1 10 0 9 1 10 9 2
52 10 9 2 11 1 10 11 11 2 13 1 9 13 10 9 1 10 9 0 13 1 10 9 1 9 7 9 1 9 0 1 10 9 2 3 15 13 1 10 9 1 9 8 10 9 1 10 9 1 10 9 2
25 3 11 11 2 9 1 10 9 2 11 1 10 9 7 1 10 9 2 13 1 11 1 10 9 2
12 10 9 0 1 11 13 3 3 0 7 0 2
22 11 1 11 13 10 9 0 0 1 10 9 1 11 1 10 9 0 1 11 2 11 2
12 1 9 2 11 3 13 3 0 16 13 15 2
33 10 9 0 13 1 11 2 11 11 11 11 2 2 10 9 1 11 2 10 15 13 1 10 9 2 10 9 1 11 2 10 11 2
19 10 9 13 10 9 1 10 9 2 10 9 7 9 11 11 1 10 9 2
15 10 9 15 13 1 10 9 1 13 10 9 1 10 9 2
36 1 10 9 2 15 13 3 1 9 1 10 11 1 11 7 10 11 11 11 11 11 7 13 10 9 1 10 9 2 11 2 2 1 11 2 2
24 1 10 9 13 10 9 1 10 0 9 16 13 10 0 9 1 9 1 10 9 1 10 9 2
24 10 9 15 13 16 13 1 10 9 2 16 13 0 1 10 9 1 13 7 16 13 1 9 2
23 1 10 9 11 15 13 10 9 9 1 10 11 0 2 11 2 13 1 0 9 1 11 2
30 10 9 1 11 7 10 9 3 13 1 9 1 10 9 2 7 13 16 4 13 1 0 7 13 1 10 9 1 13 2
24 11 13 10 9 1 9 1 10 9 1 10 9 2 11 2 11 2 2 9 1 11 7 11 2
8 13 1 12 9 7 12 9 2
59 1 10 12 9 2 11 4 13 1 10 12 5 0 2 10 12 5 13 0 2 10 12 5 13 0 2 10 12 5 13 0 2 10 12 5 13 0 1 10 11 2 10 12 5 13 1 10 9 7 10 12 5 13 1 12 7 3 9 2
24 10 11 11 1 11 2 13 1 10 9 11 2 13 10 9 0 0 1 9 0 2 11 2 2
20 9 1 10 3 3 0 11 1 11 2 10 11 11 13 15 0 7 3 0 2
42 13 12 9 0 1 10 9 1 0 9 7 10 9 0 2 3 12 9 1 9 1 2 8 8 2 7 9 0 1 10 9 0 13 1 9 2 9 9 5 12 2 2
13 10 9 15 13 1 10 9 0 1 11 1 12 2
61 10 9 13 16 10 9 1 13 15 16 10 11 7 10 9 4 13 13 3 1 10 9 1 10 9 2 3 16 10 9 1 10 9 4 13 1 10 9 2 1 0 9 16 10 9 1 10 9 4 13 1 10 9 1 9 0 13 1 10 9 12
52 10 9 10 9 13 1 10 9 2 1 9 2 13 10 9 1 11 1 10 9 11 7 11 2 2 2 7 2 10 9 3 15 13 2 13 2 1 9 2 10 9 1 11 1 11 8 11 7 11 1 11 2
41 10 9 1 9 1 10 9 1 9 2 7 10 9 1 10 9 1 15 2 13 10 9 1 10 9 7 9 1 10 9 1 12 9 16 13 10 9 1 10 11 2
24 16 15 13 3 1 10 9 1 10 9 0 1 10 9 2 3 15 13 1 9 0 1 12 2
20 10 0 9 15 4 13 1 10 9 7 10 9 15 4 13 1 10 9 0 2
42 16 10 9 13 10 9 1 9 0 2 10 9 1 10 9 1 13 4 13 0 7 10 9 1 9 2 1 10 9 10 9 0 15 13 1 9 1 10 9 1 9 2
28 10 9 1 10 9 13 10 0 9 16 13 16 3 13 10 2 11 2 16 13 15 1 15 16 13 10 9 2
31 10 9 1 9 1 11 15 13 10 9 12 2 1 9 1 10 9 16 13 1 10 0 9 1 10 9 2 3 13 0 8
29 8 0 9 15 13 1 12 9 13 1 10 11 1 10 11 1 11 11 11 1 11 2 7 4 13 1 10 9 2
32 15 16 3 13 1 0 13 16 10 9 13 10 16 13 10 9 2 10 9 2 9 7 13 0 1 9 1 9 7 9 0 2
8 15 13 9 0 15 13 9 2
38 10 9 15 13 15 13 1 9 2 7 1 9 1 9 10 9 16 10 9 13 2 9 2 7 16 15 13 13 10 9 2 13 12 9 1 10 9 2
25 1 11 3 15 13 13 1 11 2 9 16 15 13 7 16 4 13 10 9 1 13 1 10 9 2
24 10 9 1 9 0 7 10 9 16 4 13 0 4 13 3 0 1 10 9 1 9 1 9 2
23 10 9 0 13 1 10 9 12 2 7 4 13 1 10 9 1 10 9 1 10 9 12 2
49 15 13 16 4 13 10 9 1 9 1 13 15 1 13 1 10 0 11 12 1 11 1 9 1 11 2 7 16 11 10 11 4 4 1 13 9 1 15 1 10 13 10 9 13 1 10 9 0 2
27 11 13 1 11 10 9 7 10 9 0 2 3 1 13 15 1 10 9 10 9 0 1 11 1 3 13 2
41 1 10 11 2 13 1 11 11 10 9 2 13 1 10 9 0 1 10 11 11 1 10 11 2 13 1 10 0 9 1 10 9 1 11 11 2 3 13 12 9 2
20 10 9 13 1 10 9 1 15 15 13 10 9 1 0 16 3 15 13 0 2
27 1 9 2 10 9 1 9 0 3 13 10 9 1 16 10 0 9 10 9 0 4 13 9 1 10 11 2
29 1 11 2 10 9 13 10 9 1 10 9 1 10 0 11 11 1 15 1 11 11 2 10 9 0 13 3 0 2
41 11 2 11 2 11 2 1 11 11 11 15 9 2 13 10 9 7 9 1 11 2 1 10 9 1 11 2 9 1 11 2 1 10 9 1 11 7 9 1 11 2
57 3 10 9 4 13 10 9 0 2 1 9 1 9 1 10 9 2 1 10 9 7 9 1 9 2 1 10 9 7 2 9 2 1 10 9 2 1 13 10 9 2 9 2 8 2 7 3 1 9 1 13 10 9 1 10 9 2
16 10 12 9 13 10 9 0 16 13 10 9 1 12 9 0 2
134 10 11 1 9 7 9 15 13 1 0 9 10 9 1 9 3 13 10 0 9 1 9 2 10 15 13 10 9 13 1 10 9 2 11 11 11 2 1 10 9 1 10 9 2 15 13 10 12 9 7 13 9 1 10 9 13 10 10 9 2 16 13 10 0 9 1 10 9 2 10 9 15 13 1 13 10 9 1 9 1 9 16 13 10 9 1 11 7 1 16 10 9 13 9 1 9 1 15 7 9 10 15 4 13 16 13 10 9 2 15 1 10 9 4 13 1 9 15 4 13 1 10 9 2 1 10 9 1 9 1 15 3 0 2
37 3 13 10 9 1 13 1 15 1 10 0 9 1 9 16 15 13 1 10 11 1 10 9 1 10 9 7 13 10 0 9 3 1 10 0 9 2
6 13 10 9 0 0 2
14 11 13 10 9 7 13 10 9 1 10 9 1 12 2
30 1 9 1 11 2 13 15 1 10 9 1 9 0 1 10 9 12 2 12 2 7 10 0 9 1 10 9 0 0 2
10 13 0 16 13 11 16 13 10 9 2
42 10 9 3 4 4 13 3 1 2 11 2 1 10 9 2 13 1 9 1 9 0 9 1 10 9 0 1 12 5 8 2 0 9 1 10 12 5 7 10 9 0 2
43 10 9 13 10 9 1 10 9 2 1 15 16 10 9 4 13 1 10 9 0 2 7 1 10 9 2 16 10 9 3 13 0 1 10 9 1 15 15 13 10 9 2 2
45 10 9 13 16 1 9 16 13 2 12 9 16 13 1 10 9 0 1 10 9 1 10 9 1 10 0 2 13 13 1 10 9 0 1 10 0 9 16 15 4 1 13 10 9 2
44 11 1 11 11 1 9 0 2 1 10 9 0 1 10 9 1 11 16 13 1 10 9 11 2 11 2 9 1 10 9 7 10 9 2 7 11 2 9 16 13 10 9 2 2
28 1 3 1 11 2 13 16 13 13 10 9 1 10 11 11 1 0 13 10 9 1 10 9 1 13 3 9 2
38 10 0 9 0 2 11 2 13 1 10 9 12 9 0 2 15 16 13 1 10 1 10 9 7 13 10 9 1 10 10 9 2 9 2 9 7 9 2
47 10 9 1 9 15 13 1 10 9 0 1 10 11 2 1 16 10 12 1 11 1 12 2 10 12 9 13 3 3 10 9 0 1 10 11 2 7 10 9 1 13 7 13 10 9 0 2
19 15 15 13 13 10 9 1 10 9 1 11 11 7 10 9 1 11 11 2
68 1 9 15 13 1 10 12 2 7 10 9 13 1 10 9 1 10 9 1 10 9 11 2 15 3 15 13 1 9 1 10 9 7 1 10 11 2 1 9 1 10 9 0 15 4 13 10 9 0 16 4 13 1 10 9 7 16 13 16 10 11 13 9 1 10 9 0 2
7 10 9 13 1 10 9 2
54 10 9 3 1 10 9 1 11 11 2 11 2 1 3 13 10 9 1 10 0 9 0 2 10 9 0 11 15 4 13 1 10 9 1 10 9 1 3 10 9 1 9 0 7 0 13 10 9 3 0 2 13 8 2
11 10 9 2 15 13 1 12 9 1 9 2
23 10 9 13 1 9 7 9 2 7 1 9 0 2 13 1 10 9 16 13 10 9 0 2
20 11 11 11 11 2 8 11 1 11 2 9 0 2 12 1 11 1 12 2 2
40 10 9 7 10 9 1 11 11 13 0 1 10 9 1 11 11 1 10 11 11 2 9 16 1 15 4 3 13 16 4 13 1 10 0 9 1 10 9 11 2
16 10 11 15 13 1 13 10 9 2 0 2 0 7 0 2 2
34 1 10 9 0 1 10 11 15 15 13 1 10 9 1 11 2 9 16 1 9 15 13 1 15 3 0 1 10 9 7 10 9 2 2
11 13 1 10 9 1 9 1 11 1 12 2
34 4 13 1 10 11 1 11 1 10 3 9 11 11 2 7 13 1 9 1 11 11 2 13 1 2 9 7 9 1 10 9 0 2 2
12 10 9 1 9 1 10 9 13 1 5 12 2
21 13 0 2 1 9 10 9 1 10 15 9 1 9 7 15 15 4 13 7 13 2
17 4 13 0 1 10 9 1 9 1 11 2 4 13 12 9 0 2
18 1 9 4 13 10 9 0 2 13 2 11 2 7 2 11 11 2 2
34 13 10 9 11 11 2 12 1 11 1 12 2 2 15 13 1 10 9 10 9 11 2 13 16 10 10 9 1 11 7 11 4 13 2
23 11 11 2 1 9 2 13 10 9 1 9 0 1 10 9 7 10 9 13 1 10 9 2
19 3 13 1 0 9 13 1 10 9 11 7 3 16 15 13 10 9 0 2
11 15 13 10 9 7 10 9 16 15 13 2
14 1 9 2 10 9 0 1 11 11 13 1 10 9 2
27 13 10 9 1 10 9 11 16 13 10 9 1 10 9 11 7 1 12 9 2 15 1 15 3 0 11 2
38 11 11 2 11 2 11 2 12 1 11 1 12 2 7 13 10 9 0 2 16 15 13 1 9 7 16 3 13 2 1 10 11 1 10 11 1 11 2
9 4 13 1 9 1 11 11 11 2
25 10 11 11 1 11 11 15 13 3 13 3 1 12 9 2 9 1 10 15 15 13 1 0 9 2
17 3 15 13 13 10 9 0 0 1 10 0 9 1 10 11 11 2
24 10 11 11 11 2 1 9 2 11 11 11 2 13 10 9 0 16 15 13 1 11 2 11 2
19 15 4 13 9 1 10 9 7 1 10 9 1 9 1 9 16 13 0 2
23 1 16 13 1 10 9 2 13 15 3 0 1 3 1 10 9 0 7 0 1 10 9 2
52 11 11 11 11 2 11 11 2 12 1 11 12 2 13 10 9 8 7 9 0 13 1 13 10 9 1 11 1 10 9 1 11 11 7 13 1 10 9 1 10 9 1 9 11 11 11 11 13 1 11 11 2
21 10 9 0 4 13 10 9 16 13 2 0 2 1 9 1 10 9 1 9 0 2
31 10 9 15 13 3 16 11 11 13 0 7 10 9 13 0 2 1 15 15 10 9 1 11 7 10 11 4 13 15 3 2
19 10 9 15 13 1 10 9 1 0 9 7 1 9 13 10 9 1 9 2
25 11 5 12 2 3 11 5 2 13 10 9 1 9 0 0 2 1 9 2 1 10 9 11 11 2
22 10 9 1 10 9 3 13 10 9 1 10 12 5 1 10 9 2 16 13 12 9 2
40 13 1 11 2 1 9 1 12 4 1 13 1 10 11 10 0 7 0 9 0 0 11 13 1 11 12 2 3 15 13 10 0 9 7 9 1 10 9 0 2
22 10 9 1 10 9 2 11 2 15 13 1 11 1 11 10 10 11 1 12 1 12 2
17 10 9 1 10 9 13 0 1 13 1 10 12 1 11 1 12 2
26 15 13 10 0 9 1 9 1 11 2 11 1 11 13 1 9 1 9 13 15 1 9 1 1 9 2
22 1 12 13 9 1 10 11 1 11 2 13 1 13 10 9 1 11 1 11 1 12 2
14 15 15 13 1 4 13 10 9 1 11 11 1 12 2
26 1 10 9 1 10 9 2 1 12 4 1 13 9 1 10 9 2 9 1 10 15 10 9 4 13 2
37 13 9 0 15 16 13 10 11 2 10 11 7 10 11 1 10 11 11 2 3 7 10 11 2 10 11 2 10 11 7 11 11 1 10 11 11 2
37 10 11 11 11 11 11 13 16 1 9 1 10 9 13 2 15 13 9 1 9 2 9 1 9 7 9 1 0 9 1 10 9 1 10 9 11 2
21 10 9 11 13 13 2 7 4 13 7 13 1 11 2 1 3 15 13 10 9 2
48 15 1 10 9 13 3 0 7 2 16 15 13 1 10 9 9 1 9 2 4 13 1 10 9 7 9 9 2 3 1 4 13 1 13 7 13 16 1 9 1 10 9 10 9 15 15 13 2
46 1 0 9 2 10 9 3 15 13 2 3 3 4 13 10 9 2 2 1 15 15 15 4 7 4 1 13 1 10 9 2 13 15 0 3 1 13 1 10 9 12 9 1 10 9 2
29 1 9 1 9 1 10 9 1 10 9 0 1 10 11 11 2 10 0 9 1 10 9 13 1 10 9 1 11 2
12 10 9 13 1 12 2 16 15 13 10 9 2
13 1 12 2 10 9 1 9 0 13 10 9 0 2
13 11 11 13 10 9 1 9 0 1 10 9 11 2
38 11 13 2 1 10 9 1 9 1 11 2 11 11 2 2 1 10 0 9 1 13 11 16 13 13 10 9 1 11 7 10 9 1 3 1 12 9 2
18 10 9 7 10 9 15 13 13 1 9 10 9 16 13 1 0 9 2
52 2 1 12 9 4 13 9 0 2 3 1 12 12 12 9 1 9 1 9 0 2 0 7 1 10 10 0 9 16 4 13 10 0 9 1 10 0 9 16 15 13 1 3 2 13 10 9 2 11 11 11 2
23 15 13 1 9 1 10 12 9 2 7 13 16 10 9 1 13 15 1 10 9 13 0 2
28 7 16 3 16 15 15 13 15 13 1 10 9 16 4 13 0 1 10 9 8 10 9 16 15 13 1 9 2
30 10 9 0 1 13 10 0 9 1 11 2 12 2 13 7 13 10 9 2 13 10 9 0 16 13 1 10 9 0 2
33 10 11 11 4 4 13 10 9 0 2 7 3 4 13 13 15 1 9 0 2 16 15 13 3 1 10 9 0 1 11 7 11 2
10 3 8 13 1 10 9 1 10 9 2
16 11 13 10 9 13 1 10 9 1 11 2 1 10 11 11 2
39 13 10 11 1 10 11 1 10 11 1 11 11 7 11 13 1 11 2 11 7 11 2 11 2 11 2 10 9 1 10 9 13 1 11 11 7 11 11 2
40 11 13 10 9 7 9 0 2 1 10 9 1 11 2 9 2 11 11 2 9 1 9 11 2 1 10 9 1 11 7 9 1 11 2 11 2 11 2 11 2
25 1 11 15 13 13 1 10 9 1 10 9 0 7 13 1 10 9 3 15 13 2 10 11 11 2
10 10 9 13 10 9 0 1 10 9 2
27 13 1 10 9 1 11 2 1 10 9 1 10 11 1 10 11 7 13 1 10 11 1 12 9 1 11 2
17 15 13 10 9 1 9 0 2 7 13 13 1 9 1 9 0 2
23 11 7 11 15 13 2 7 10 0 9 15 13 1 13 10 9 7 13 15 1 10 9 2
19 11 13 10 9 1 11 13 1 10 9 1 10 9 0 13 1 10 9 2
37 1 13 10 11 11 10 9 16 13 10 9 1 9 0 2 0 7 9 2 10 9 1 10 9 4 13 1 13 9 0 7 16 4 13 3 0 2
29 1 15 15 3 10 12 5 13 3 1 11 2 16 10 9 13 9 16 15 13 3 1 10 9 7 1 10 9 2
39 10 11 1 11 3 13 10 9 16 13 1 10 9 1 9 0 2 3 15 13 10 11 11 16 13 1 10 9 11 11 1 0 9 16 3 13 11 11 2
44 10 9 1 10 12 9 0 2 16 13 1 10 9 0 0 2 8 2 2 13 10 2 9 0 2 1 10 9 7 1 10 9 16 15 13 2 16 13 10 9 1 10 9 2
15 10 9 13 3 0 2 10 9 0 7 10 9 3 0 2
30 1 10 9 1 10 9 1 12 10 9 0 1 9 1 10 9 13 1 9 12 7 10 9 0 1 9 13 9 12 2
34 10 0 9 11 11 15 13 10 9 1 10 9 1 11 11 1 10 11 11 1 11 2 11 2 1 10 9 1 10 9 1 10 11 2
46 11 4 13 10 9 2 10 9 1 10 9 1 11 2 13 1 10 9 1 4 13 10 0 9 1 10 9 0 2 10 9 1 10 15 13 7 13 10 9 0 13 9 0 1 11 2
47 13 2 1 10 9 2 10 1 0 9 7 9 1 10 11 11 1 10 11 1 11 2 1 11 7 11 1 12 2 3 1 10 1 9 1 10 11 7 10 1 9 1 10 11 1 11 2
38 10 9 1 9 13 4 4 13 1 10 9 1 9 16 13 1 10 12 1 11 2 9 1 9 1 10 9 2 1 10 9 2 12 9 7 12 3 2
42 11 7 11 2 1 9 7 3 11 2 13 10 9 1 11 11 2 8 2 8 2 13 10 9 1 10 9 1 10 11 1 10 9 1 11 2 11 11 2 11 2 2
9 10 9 13 1 10 9 1 9 2
18 10 9 1 10 9 13 13 10 9 1 9 0 1 10 9 0 0 2
28 12 9 3 3 13 9 1 10 9 11 11 1 11 11 2 1 11 11 2 1 10 15 4 13 1 11 11 2
34 1 9 1 10 9 1 10 9 11 2 15 13 16 10 12 13 1 10 12 5 1 10 9 2 0 1 10 9 1 10 9 10 12 2
53 13 1 10 9 2 1 10 9 0 2 3 13 1 10 8 12 2 7 13 5 12 1 9 2 7 13 1 9 10 9 2 12 2 2 4 13 15 10 9 1 12 9 2 3 2 1 9 1 12 10 12 9 2
41 10 9 1 9 1 10 9 1 11 13 10 11 0 7 0 2 13 15 3 1 11 2 11 2 11 11 2 11 2 11 2 11 2 11 2 11 2 11 7 11 2
13 10 9 13 1 11 2 13 1 10 9 1 12 2
27 7 13 16 11 11 15 13 3 1 9 13 9 1 11 11 2 3 7 10 9 0 15 13 10 9 11 2
23 13 1 10 9 2 3 15 13 3 1 10 9 0 2 1 15 15 15 13 3 11 11 2
13 10 9 13 3 10 9 1 12 9 1 9 0 2
48 10 9 1 11 11 11 2 1 9 2 11 11 11 11 2 13 10 9 0 0 13 3 3 1 10 9 1 10 9 1 10 11 11 11 11 11 2 8 2 2 7 3 1 10 9 15 13 2
38 11 11 7 11 2 11 2 11 2 11 2 12 1 11 1 12 2 11 2 11 2 11 2 12 1 11 1 12 2 13 10 9 7 9 1 9 0 2
32 10 11 2 11 13 10 9 7 9 0 13 1 10 9 1 11 11 2 9 1 11 2 1 10 9 1 11 7 9 1 11 2
21 11 13 0 9 16 11 11 15 13 9 1 10 9 7 15 13 1 10 9 0 2
40 1 10 9 10 9 3 0 13 10 9 7 10 0 9 10 9 15 13 13 16 10 9 15 13 1 10 10 9 1 10 9 7 13 9 3 1 10 12 9 2
12 10 9 1 3 13 16 13 0 1 9 9 2
67 10 11 13 1 15 1 11 2 15 1 11 13 1 10 11 2 2 13 15 3 9 1 10 9 1 1 15 15 13 1 15 16 15 13 3 1 10 9 2 7 10 9 0 3 15 13 2 13 1 13 2 10 11 7 11 13 10 9 0 1 13 9 1 11 7 11 2
24 3 15 13 10 9 1 10 9 1 10 9 1 10 9 16 4 13 12 7 3 9 1 9 2
16 1 10 0 9 10 9 1 9 4 13 10 9 1 10 9 2
53 1 10 9 1 10 11 11 11 2 4 13 1 10 9 1 3 1 12 9 0 1 13 15 1 10 9 1 9 1 11 2 10 9 1 9 1 9 1 10 0 9 1 9 13 11 2 16 13 1 12 7 12 2
8 11 2 11 11 11 2 12 2
39 11 11 11 2 12 1 11 1 12 2 13 9 2 9 7 9 1 11 11 2 15 1 10 0 9 1 11 11 2 10 15 13 7 13 1 12 1 12 2
17 10 9 3 13 9 1 13 10 9 2 13 0 1 13 9 0 2
54 9 1 10 9 7 9 2 4 13 1 13 10 9 1 10 11 11 1 9 13 1 9 1 9 1 10 9 1 10 9 1 11 11 11 2 11 11 2 11 11 2 11 11 7 11 11 7 1 0 9 1 11 11 2
43 10 9 13 10 9 10 12 1 11 2 16 10 9 13 10 0 9 13 10 9 1 10 9 9 2 1 10 9 15 15 13 1 10 11 1 11 11 10 9 1 10 9 2
42 9 0 16 13 1 3 1 12 9 2 4 3 3 13 1 13 10 0 9 1 10 9 0 0 11 11 11 11 11 2 1 10 15 15 13 12 9 1 12 7 12 2
22 10 9 13 10 9 0 1 10 9 1 10 9 1 9 1 9 7 1 10 9 0 2
23 15 13 15 1 9 2 7 1 9 8 9 1 9 16 13 13 10 9 1 10 9 0 2
14 13 13 1 10 13 15 10 9 0 9 1 9 0 2
14 9 0 1 10 9 2 9 1 9 0 7 10 9 2
38 10 0 9 1 9 1 9 1 10 11 2 3 7 10 9 1 10 9 0 2 13 10 9 1 10 9 1 16 11 4 13 10 9 1 10 9 0 2
42 10 9 3 2 15 13 1 10 3 11 12 1 10 0 9 1 12 2 16 10 9 11 11 13 10 9 7 13 1 13 15 11 11 13 10 9 1 2 9 0 2 2
16 10 9 1 9 0 13 3 0 7 10 9 0 1 10 9 2
7 3 2 15 13 10 9 2
12 10 9 1 11 11 15 13 13 1 10 9 2
26 10 9 13 15 0 2 8 1 10 9 2 2 16 10 9 13 1 4 15 1 13 1 9 2 3 2
12 11 13 1 11 11 7 1 10 11 1 13 2
48 10 9 1 9 1 10 9 1 11 7 10 11 11 13 10 9 0 1 10 9 0 1 10 9 1 10 9 16 4 13 10 9 3 7 16 13 1 10 9 0 1 10 9 1 10 12 9 2
37 10 9 2 16 4 13 1 10 9 0 2 13 10 9 0 1 10 0 11 1 10 8 1 10 9 2 11 11 2 16 4 13 1 10 9 0 2
63 1 10 12 9 2 10 9 1 11 11 4 13 1 10 12 5 9 2 10 12 5 13 9 2 10 12 5 13 9 2 10 12 5 13 9 2 10 12 5 13 9 1 10 11 2 10 12 5 13 1 10 9 7 10 12 5 13 1 12 7 3 9 2
43 1 12 2 16 13 12 9 2 10 9 13 10 9 0 7 13 1 10 9 2 7 15 7 10 9 4 13 1 10 9 1 9 0 1 11 2 1 9 3 13 1 11 2
17 10 9 13 0 2 3 0 2 1 10 9 1 12 1 12 9 2
62 1 10 12 9 2 10 9 1 11 4 13 1 10 12 5 0 2 10 12 5 13 0 2 10 12 5 13 0 2 10 12 5 13 0 2 10 12 5 13 0 1 10 11 2 10 12 5 13 1 10 9 7 10 12 5 13 1 12 7 3 9 2
27 1 10 10 9 1 10 9 2 13 10 9 1 12 2 1 10 9 0 1 11 2 9 2 11 11 2 2
31 3 1 10 9 15 4 13 10 0 9 1 9 1 10 11 11 1 9 3 0 1 9 2 0 2 7 1 2 9 2 2
10 11 11 2 2 10 9 15 13 2 2
28 0 1 9 1 12 2 1 10 9 11 13 1 11 2 9 7 11 2 13 10 9 1 9 1 9 3 0 2
20 10 9 13 3 1 10 8 1 9 4 4 13 1 10 9 9 1 11 11 2
37 10 0 9 1 9 1 9 1 9 4 4 13 7 15 13 1 10 0 9 1 9 1 9 1 13 9 7 9 1 13 1 13 10 9 3 0 2
43 1 2 10 11 11 2 15 13 1 9 1 10 0 9 0 2 16 1 13 15 2 13 12 0 9 1 10 9 16 15 13 1 13 7 13 1 10 9 11 11 1 11 2
16 11 7 10 15 9 13 1 9 7 15 13 0 1 10 9 2
36 15 1 10 9 3 13 1 10 9 0 13 10 9 11 2 10 9 3 0 1 10 9 16 10 9 13 10 9 1 13 15 1 9 1 9 2
17 10 10 9 1 10 9 0 0 4 13 1 10 9 0 11 11 2
16 13 10 0 7 0 9 1 11 12 1 11 7 11 1 11 2
20 10 9 0 13 10 0 9 1 11 1 3 1 10 9 1 10 9 0 0 2
20 10 9 1 10 9 15 13 1 10 9 1 10 9 1 9 2 9 7 9 2
48 3 15 13 1 9 0 2 1 9 2 10 11 11 2 9 7 11 13 3 0 2 1 15 15 13 3 1 10 9 2 2 7 16 1 10 9 1 11 2 9 2 13 1 13 15 3 0 2
18 1 10 9 0 7 0 0 3 15 13 9 1 12 9 1 12 9 2
23 16 10 9 1 10 9 15 13 2 11 13 1 10 9 0 1 10 9 1 11 1 11 2
11 10 9 1 11 15 13 13 1 10 9 2
25 1 3 13 15 2 13 1 10 10 9 13 16 10 9 11 1 11 13 9 10 1 13 10 9 2
16 1 10 9 13 1 11 2 1 10 9 3 0 13 10 9 2
14 13 1 13 15 1 12 1 10 9 2 11 11 11 2
10 13 0 1 11 1 10 9 1 11 2
54 13 9 1 9 0 1 9 0 2 11 1 11 2 10 9 15 15 13 2 10 9 1 10 9 2 10 9 16 13 10 9 0 2 11 10 0 9 2 11 0 2 10 9 1 11 11 2 11 7 10 9 1 11 2
33 10 11 13 13 3 1 10 0 9 1 13 15 10 9 2 13 1 16 3 13 16 10 9 13 7 3 10 9 1 10 10 9 2
51 16 15 3 13 10 0 9 1 10 9 1 11 9 1 10 9 1 11 2 16 13 3 0 13 1 10 0 9 1 11 7 10 9 0 2 3 15 13 16 10 9 1 11 3 4 4 13 3 1 12 2
6 10 9 3 13 9 2
12 3 7 4 13 15 10 9 1 10 0 9 2
16 15 13 1 12 9 2 15 0 7 12 9 7 1 12 9 2
12 10 9 0 7 0 9 0 13 1 10 9 2
27 10 9 1 11 2 1 9 2 11 11 2 13 10 9 13 1 10 9 1 11 1 10 9 0 1 11 2
34 1 10 9 15 13 1 9 1 9 7 9 7 1 16 15 15 13 9 13 13 10 9 1 10 9 2 16 13 0 9 1 10 9 2
25 3 1 10 9 2 10 11 2 12 13 1 3 1 10 9 0 7 13 1 10 9 1 10 11 2
7 15 13 1 11 7 11 2
36 1 10 9 1 11 11 15 13 3 1 10 9 0 1 10 9 1 10 9 1 11 1 11 2 15 3 4 13 3 1 10 9 0 1 11 2
24 10 3 0 9 1 9 13 10 9 1 9 1 11 11 2 11 15 8 11 2 1 10 12 2
18 10 9 0 13 10 9 0 0 7 4 7 13 15 10 9 1 9 2
37 10 9 0 13 1 10 0 9 1 10 12 2 10 9 1 11 11 2 15 13 10 9 1 10 9 1 15 15 13 10 9 0 1 10 11 11 2
14 3 4 13 1 10 9 0 7 15 1 10 9 13 2
17 10 9 4 13 9 1 9 0 7 13 0 2 13 7 15 13 2
29 11 13 10 9 1 9 1 10 9 0 13 1 10 9 1 13 10 9 2 9 2 1 9 0 1 9 1 9 2
33 1 10 9 2 1 12 2 10 9 13 13 10 9 1 11 11 1 10 9 1 11 11 7 15 15 13 1 11 1 16 15 13 2
45 1 9 2 1 10 9 12 11 4 13 10 9 1 10 0 9 11 11 7 2 3 1 13 10 9 2 4 1 13 1 10 9 0 1 10 9 0 7 0 2 3 0 11 11 2
38 10 9 1 11 13 10 9 1 9 2 10 9 1 10 16 10 9 1 9 13 10 9 0 1 0 9 1 9 7 10 0 9 1 10 9 1 9 2
26 11 1 11 2 12 2 12 2 13 10 9 0 1 11 11 16 13 1 10 9 1 10 9 11 11 2
16 1 10 9 2 12 12 9 15 13 1 10 9 1 10 11 2
23 1 9 1 12 2 13 1 11 2 10 0 9 7 10 9 1 10 9 1 10 9 0 2
6 10 0 9 13 11 2
14 3 3 1 10 9 13 10 9 16 13 1 10 9 2
19 3 9 10 15 1 10 9 13 3 0 9 1 9 1 0 9 1 11 2
29 16 10 9 13 3 10 0 9 2 10 9 13 10 9 1 13 10 9 0 1 10 9 2 13 3 0 10 9 2
19 0 9 13 10 9 2 13 15 1 13 12 9 2 12 9 2 1 9 2
13 10 9 1 9 13 1 12 9 2 2 9 5 2
17 11 10 9 13 10 9 1 10 11 11 10 12 1 11 1 12 2
56 11 2 7 10 9 2 11 11 2 13 3 10 9 13 1 10 11 2 8 8 8 2 9 1 9 0 2 2 1 15 15 1 9 10 11 13 1 11 13 10 9 1 10 9 1 10 9 11 2 9 1 10 15 3 13 2
54 1 13 1 10 12 1 11 1 12 2 10 9 1 9 1 10 9 1 10 9 2 3 7 10 9 0 2 10 15 13 10 9 1 10 0 9 1 9 1 10 9 2 15 13 1 9 1 10 9 1 9 7 9 2
21 9 13 0 2 10 9 15 13 3 3 1 15 9 7 1 9 2 9 7 9 2
41 10 9 1 11 15 13 10 12 1 11 1 12 1 10 9 1 10 11 2 11 2 1 9 1 11 7 11 2 16 13 0 1 11 1 10 11 11 2 7 11 2
30 1 10 9 2 10 9 0 15 13 1 0 9 1 10 9 0 2 1 12 9 2 1 12 1 10 9 2 11 2 2
22 1 10 9 1 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 9 5 2
31 10 9 2 10 11 2 3 13 10 11 9 1 11 11 13 1 10 9 11 11 1 10 9 1 15 1 10 9 1 11 2
22 10 9 10 11 1 10 11 2 12 2 2 4 13 1 10 9 1 10 9 3 0 2
31 8 3 15 2 9 4 13 10 9 13 1 11 12 9 7 12 9 1 10 9 1 10 9 11 7 10 9 0 9 12 2
42 1 12 2 3 1 16 10 9 4 4 13 16 13 10 9 2 13 9 10 11 11 2 1 10 15 10 9 15 13 1 13 15 7 13 10 9 1 10 9 1 9 2
19 1 9 1 12 2 1 10 9 1 9 2 4 7 13 1 10 9 0 2
15 10 11 11 1 10 0 9 13 9 1 15 1 10 9 2
51 10 0 12 9 3 15 4 13 9 1 10 11 1 10 11 2 7 16 10 12 0 9 4 13 1 10 9 16 13 10 9 9 9 1 10 9 1 10 2 11 1 11 11 1 11 2 13 1 10 9 2
14 11 4 7 13 10 9 1 12 9 7 13 10 12 2
30 10 11 2 11 11 1 10 11 2 13 10 9 1 9 13 3 1 9 3 1 9 16 13 2 13 7 13 10 9 2
15 1 12 13 11 16 13 15 3 1 10 9 0 2 11 2
25 1 10 9 10 9 13 0 9 2 9 2 9 2 8 2 7 13 10 9 1 13 10 12 9 2
33 11 7 11 11 2 11 2 2 10 9 0 9 1 10 9 11 2 13 10 9 1 10 9 0 1 13 1 10 0 12 1 11 2
35 11 11 11 10 11 2 11 11 2 11 2 12 1 11 1 12 2 13 10 9 0 7 9 1 9 2 0 1 9 2 13 1 9 0 2
13 10 9 11 15 13 1 11 1 10 11 9 12 2
16 1 9 0 13 0 16 10 0 9 13 10 9 1 10 9 2
24 10 9 1 10 0 9 2 3 15 3 2 15 13 1 13 10 9 7 13 1 10 9 0 2
20 13 16 10 9 2 11 2 15 13 1 13 7 13 1 10 9 1 10 9 2
32 1 9 12 1 11 1 12 2 15 15 13 9 0 1 10 9 1 9 1 9 1 9 0 1 10 11 11 1 10 11 11 2
29 13 9 1 10 9 12 1 10 9 11 11 11 1 9 1 10 11 11 2 13 1 12 1 10 9 11 11 11 2
20 3 2 13 1 10 9 0 16 13 1 11 1 11 7 11 2 13 1 11 2
24 11 3 13 1 10 9 2 3 16 11 11 12 1 11 13 10 9 3 1 9 1 10 9 2
13 13 10 9 5 12 1 8 8 8 12 8 8 2
19 10 9 0 3 13 3 7 16 15 4 13 7 4 13 3 1 10 9 2
22 1 10 9 13 10 9 16 3 13 1 10 9 7 10 9 3 13 1 15 4 13 2
35 10 9 1 10 9 4 13 3 16 9 1 9 15 13 1 10 9 2 16 13 1 10 9 10 9 7 2 3 3 2 10 9 7 9 2
7 2 11 11 13 1 11 2
30 11 11 13 3 3 13 1 13 10 9 1 11 11 2 7 11 11 1 13 10 9 1 10 11 2 7 11 11 11 2
26 13 3 1 0 9 10 9 1 9 0 1 11 1 10 0 11 1 11 0 1 10 9 1 11 11 2
19 9 12 8 1 0 7 12 8 1 0 2 11 7 11 2 0 7 9 2
20 13 13 1 9 1 10 11 11 11 2 1 10 9 1 11 11 2 11 11 2
21 13 2 15 13 1 15 9 1 10 9 7 13 3 7 8 1 9 15 15 13 2
44 10 9 15 15 15 13 13 1 9 2 9 2 9 0 7 0 2 9 2 3 1 9 2 2 9 2 9 1 9 2 9 9 0 2 9 7 1 9 10 9 4 13 0 2
36 10 9 1 10 9 1 10 9 13 0 9 2 7 13 9 1 10 9 1 10 9 7 1 10 9 0 1 10 0 9 1 11 11 1 9 2
9 1 10 9 2 13 13 10 0 2
18 13 15 9 16 15 13 1 10 9 7 3 1 10 9 1 10 9 2
9 3 13 16 15 13 1 10 9 2
13 13 10 9 13 0 9 1 9 7 10 9 0 2
27 16 15 13 10 9 0 2 15 4 13 1 10 9 10 9 0 1 9 0 2 1 13 10 9 1 9 2
48 10 12 1 11 1 12 4 13 9 1 10 11 1 10 11 1 10 12 9 1 12 9 1 9 1 10 12 9 1 10 11 11 2 1 10 13 1 10 9 1 10 11 11 7 11 7 11 2
58 13 10 9 0 1 0 1 10 9 0 1 10 9 0 1 10 9 2 13 1 9 0 9 2 9 0 2 1 10 9 0 15 13 1 0 9 2 1 9 13 1 10 9 2 16 13 10 9 0 2 1 9 0 2 0 7 0 2
20 11 11 13 10 0 9 1 9 1 11 11 1 9 1 10 9 0 11 11 2
8 13 10 12 1 11 1 12 2
49 10 9 2 3 0 2 3 0 7 15 0 1 10 0 9 0 2 4 13 3 10 0 9 0 1 9 2 9 2 9 2 2 13 9 0 1 9 1 10 9 2 3 0 1 10 0 9 2 2
38 11 11 2 13 10 0 9 2 2 13 11 11 11 2 10 9 1 10 11 1 10 9 2 2 7 13 3 0 13 15 15 4 13 15 15 13 2 2
21 10 11 11 11 7 11 9 11 13 10 9 1 9 3 1 10 9 1 11 11 2
7 3 15 13 1 10 9 2
13 10 9 11 15 13 1 10 0 9 0 1 11 2
18 3 1 12 9 4 13 2 1 10 0 12 9 2 0 9 7 9 2
18 15 13 1 0 13 1 10 9 1 10 9 11 11 1 10 9 0 2
26 1 12 7 12 13 10 9 1 0 9 1 9 2 1 15 2 10 1 10 11 11 8 11 1 11 2
34 1 10 9 3 13 3 0 13 1 9 12 9 0 2 9 0 1 10 9 7 16 13 1 10 9 0 2 13 10 8 11 11 11 2
11 4 13 10 9 7 10 9 13 0 9 2
19 13 1 9 0 7 9 13 10 9 1 10 15 15 13 9 1 10 9 2
23 3 15 13 16 15 13 12 5 1 9 7 10 9 1 12 5 7 9 10 9 16 13 2
38 11 13 10 9 16 3 15 13 0 1 2 11 11 11 11 2 11 2 7 1 9 2 15 13 7 8 2 13 10 9 1 10 0 9 1 10 9 2
13 3 0 2 1 12 13 10 9 9 1 10 9 2
11 1 10 9 10 9 13 1 10 9 0 2
26 1 9 2 1 13 10 9 2 10 9 15 13 10 9 1 10 11 11 11 7 1 10 11 11 11 2
20 11 13 0 9 0 1 10 9 2 9 0 1 9 0 9 3 3 3 13 2
26 10 9 13 1 10 9 1 10 0 9 11 1 10 9 11 2 9 1 10 15 13 10 9 1 9 2
56 1 9 1 10 9 1 9 11 8 2 1 11 1 12 13 10 9 1 10 11 1 11 1 10 9 7 0 9 2 13 1 9 0 7 1 9 1 11 10 11 2 13 1 10 13 10 9 1 10 9 1 10 9 1 9 2
20 1 9 3 15 15 13 9 0 7 11 13 1 10 9 1 11 1 12 9 2
39 13 1 10 11 11 1 11 10 12 1 11 1 10 9 11 8 11 11 11 2 7 12 9 3 3 13 10 0 9 2 12 1 11 1 10 11 11 2 2
16 9 7 9 0 1 10 11 11 1 10 11 11 2 11 12 2
47 10 9 13 10 9 1 10 9 16 13 1 3 9 7 1 10 9 1 12 1 10 0 11 1 9 1 9 1 12 8 5 9 13 15 2 1 10 9 2 1 12 1 12 8 5 9 2
23 11 4 13 9 0 2 9 1 9 2 9 7 9 0 1 10 9 1 9 11 7 11 2
13 13 1 11 11 11 7 3 1 10 9 1 9 2
18 11 1 12 11 13 10 0 9 13 1 10 9 1 11 11 10 11 2
9 13 10 0 9 1 10 9 11 2
4 0 1 11 2
26 10 9 1 10 9 0 13 10 9 2 1 15 15 4 10 9 1 13 10 9 15 13 10 10 9 2
16 11 11 13 10 9 1 9 1 10 9 11 1 10 9 11 2
59 1 9 2 1 10 9 1 9 0 2 15 2 1 10 13 10 9 1 10 9 2 15 13 16 1 9 3 13 1 11 1 15 15 13 13 15 2 13 1 10 9 7 13 16 15 13 1 10 9 10 9 7 10 9 16 13 10 9 2
11 10 9 1 11 15 13 0 1 10 9 2
38 11 2 15 15 4 13 1 11 11 1 12 15 13 1 13 1 12 7 13 10 9 0 1 9 3 0 1 11 11 2 13 10 9 11 12 7 12 2
31 1 9 2 10 11 1 11 1 10 11 13 16 15 13 9 1 9 0 1 10 9 7 2 1 10 9 1 10 9 2 2
26 15 13 3 0 1 10 9 1 9 1 10 9 1 10 0 9 1 11 2 13 1 13 1 10 9 2
20 10 9 13 1 9 2 9 7 9 0 1 9 7 10 9 3 0 1 9 2
22 10 9 1 10 9 4 13 3 1 10 9 7 13 1 9 1 10 9 13 1 15 2
32 7 16 3 3 13 1 10 0 9 2 10 11 11 12 13 13 1 9 1 8 16 15 13 1 10 9 16 13 3 10 9 2
10 15 4 13 1 9 3 1 12 9 2
30 1 10 9 15 13 10 9 1 10 9 16 13 10 9 1 10 11 1 11 1 9 1 10 0 9 13 1 9 0 2
15 10 9 1 10 15 15 4 13 10 9 13 1 11 11 2
18 10 9 1 11 13 0 7 15 13 10 9 0 1 10 9 1 11 2
14 10 9 12 13 10 3 0 1 10 10 9 1 11 2
41 10 9 1 10 9 0 13 16 1 10 0 9 15 4 13 1 10 9 1 10 9 1 12 12 9 1 9 13 10 9 1 9 1 9 0 1 10 9 1 11 2
36 1 10 9 2 10 0 9 15 13 10 9 1 10 9 2 3 1 9 0 7 0 1 10 9 1 10 9 0 1 9 7 15 0 1 9 2
11 10 9 13 10 9 1 11 7 11 11 2
23 13 1 11 16 15 13 10 9 1 4 4 13 7 13 10 0 9 1 11 1 10 9 2
33 1 10 9 0 13 9 12 1 10 12 9 0 1 10 9 2 10 15 1 10 9 1 10 9 2 11 2 11 2 11 7 11 2
45 1 12 13 3 11 1 13 11 1 10 9 13 1 11 11 2 9 2 2 11 11 2 9 2 2 11 11 11 2 9 2 2 11 1 11 2 9 2 7 11 11 2 9 2 2
11 10 9 1 9 15 13 1 11 1 12 2
29 1 10 2 9 2 16 15 13 1 10 13 1 15 2 4 13 15 10 9 16 13 1 10 9 1 13 10 9 2
15 1 11 13 10 12 9 2 7 3 12 9 1 9 0 2
23 9 13 16 11 2 9 15 4 13 1 10 11 1 9 7 13 10 9 0 1 10 9 2
27 10 9 0 11 11 13 10 9 1 9 1 11 2 1 10 9 0 1 11 1 11 1 10 9 1 11 2
42 10 9 1 9 15 13 1 10 9 1 10 9 11 11 2 15 13 10 9 1 9 7 9 1 13 10 9 1 9 2 1 10 9 1 13 1 10 9 1 9 0 2
14 11 11 11 13 10 9 16 3 10 10 9 13 0 2
9 10 9 0 13 12 7 12 9 2
20 16 13 3 13 7 9 7 10 9 16 1 10 9 15 13 7 15 13 15 2
18 10 9 2 1 9 2 13 1 9 0 1 10 9 16 13 10 9 2
21 1 10 9 13 1 10 9 0 1 10 9 2 11 7 11 15 13 1 9 0 2
29 13 9 1 9 1 10 9 1 10 11 1 12 7 12 2 9 1 10 15 13 1 10 9 0 1 9 1 11 2
19 10 9 1 9 1 11 13 10 9 0 1 9 1 10 9 1 10 11 2
22 10 2 11 11 11 2 15 13 1 10 9 2 13 1 10 9 16 15 13 10 9 2
14 11 13 10 9 9 1 9 1 10 9 11 11 11 2
32 1 12 2 1 10 9 1 11 12 1 11 2 10 9 13 10 9 1 9 1 13 10 9 0 0 2 16 13 1 10 9 2
60 10 3 0 9 1 10 9 0 15 13 1 10 9 1 10 11 1 11 13 2 10 9 0 2 2 10 15 13 10 9 1 10 11 3 16 1 9 1 13 10 9 2 10 9 13 10 9 1 10 15 15 13 10 9 1 10 11 1 11 2
8 13 9 7 9 1 0 9 2
18 3 1 13 10 9 1 11 2 11 11 13 1 10 9 1 13 11 2
30 10 0 9 13 1 10 9 7 9 4 13 10 9 1 3 7 4 4 13 1 9 0 1 9 1 10 9 1 9 2
49 1 12 2 10 9 11 11 13 15 1 10 0 9 16 3 13 10 9 1 10 9 1 9 1 9 1 10 9 2 0 1 10 9 1 9 1 10 11 11 2 1 0 9 2 1 13 10 9 2
26 1 12 13 10 9 1 9 11 1 10 9 0 11 11 11 7 10 9 0 1 9 0 2 11 2 2
21 11 11 11 11 2 13 1 11 1 11 2 0 9 1 11 9 1 11 2 11 2
61 13 7 13 1 10 9 1 2 3 7 3 13 3 2 10 9 3 0 1 2 9 2 4 13 1 13 15 1 15 0 3 1 10 0 9 1 9 2 16 4 13 16 3 3 2 13 9 9 2 13 0 2 7 16 3 15 13 3 13 15 2
29 11 13 10 9 11 1 10 9 9 9 1 11 11 11 11 7 10 9 8 2 15 3 13 10 9 2 11 2 2
7 3 3 4 7 13 9 2
12 15 9 13 13 1 9 1 10 9 1 9 2
15 11 11 4 13 16 11 13 9 1 10 9 1 10 9 2
30 15 13 1 9 1 10 9 1 10 0 9 1 9 1 9 9 1 10 11 11 1 10 11 1 11 11 1 11 11 2
15 9 1 9 1 10 9 1 10 9 1 10 9 11 11 2
24 16 13 11 2 10 9 15 4 13 13 10 9 7 13 13 1 13 10 9 1 10 9 0 2
34 10 9 1 9 1 13 10 9 13 0 1 10 9 1 9 16 1 10 9 15 4 13 2 1 10 9 10 9 15 13 1 11 2 2
29 13 1 10 9 1 10 9 2 10 9 3 4 13 1 0 2 7 3 13 3 3 7 13 1 10 9 1 9 2
19 3 10 9 13 1 10 9 2 16 13 9 2 15 13 9 3 9 2 2
12 15 13 1 9 1 9 1 9 1 9 0 2
23 1 9 1 10 9 10 9 0 15 13 0 1 16 11 13 10 9 0 0 1 10 9 2
36 10 15 13 1 10 9 1 11 1 9 1 11 2 10 9 15 13 10 12 1 10 9 2 2 1 10 9 1 12 2 12 7 12 9 3 2
9 15 13 16 10 9 3 13 0 2
25 10 11 13 10 9 1 12 13 7 13 1 11 11 2 1 11 11 7 11 11 13 10 9 0 2
25 10 9 2 13 1 0 1 12 2 15 13 1 10 9 1 13 1 10 9 0 1 10 9 0 2
22 11 13 10 12 1 11 1 12 2 1 10 12 9 1 9 2 13 1 10 9 0 2
16 11 13 12 9 1 10 9 2 1 10 15 13 3 0 9 2
21 1 10 9 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 9 8 2
16 10 9 4 13 10 9 1 10 9 1 9 1 10 9 0 2
59 11 2 1 10 13 10 9 2 15 13 7 13 1 10 9 2 7 1 10 13 4 1 13 10 9 1 11 2 1 9 1 10 9 15 13 9 1 16 11 13 15 9 15 11 13 2 7 3 13 10 9 1 10 9 2 1 13 15 2
38 10 9 0 1 10 11 7 10 9 0 1 11 15 4 13 1 12 1 10 3 0 9 1 10 9 0 0 2 13 10 9 1 10 9 7 9 0 2
28 13 3 0 1 10 9 0 1 11 1 11 1 9 0 7 0 1 9 1 9 2 9 7 9 1 10 9 2
51 11 13 10 9 1 11 7 11 1 10 9 1 10 11 1 10 11 13 1 10 11 1 10 9 0 1 11 7 1 10 16 13 10 9 1 11 11 2 10 9 13 8 15 13 13 2 0 7 3 2 2
21 10 0 9 13 9 9 1 9 7 10 9 0 13 10 9 7 10 9 9 0 2
16 3 13 10 9 16 13 13 2 3 15 4 13 11 1 11 2
18 10 9 0 11 11 13 12 9 1 9 1 11 1 10 9 1 9 2
17 15 13 1 10 9 0 2 11 2 10 9 1 10 9 1 11 2
45 11 7 11 11 2 2 9 1 10 9 2 11 1 10 9 8 2 2 2 16 4 0 1 10 11 2 13 10 9 13 16 13 10 0 9 1 3 15 13 1 10 4 13 0 2
29 10 9 1 11 2 11 15 13 1 11 2 11 2 11 2 7 4 13 2 12 2 1 11 11 1 10 11 11 2
28 1 9 1 13 10 0 9 7 1 11 2 10 9 0 15 13 1 9 1 0 9 1 10 9 1 10 9 2
13 1 10 9 15 13 10 9 11 7 10 9 11 2
13 1 10 11 1 12 2 13 12 9 13 1 11 2
19 1 12 13 13 1 10 9 2 13 3 10 0 9 1 9 10 9 0 2
24 12 9 1 10 9 0 0 2 13 12 9 2 4 13 1 10 9 0 2 4 13 7 13 2
46 7 10 9 0 7 10 9 13 10 0 9 2 7 10 9 0 13 15 1 10 3 9 1 10 9 2 15 16 1 15 15 13 10 9 2 1 11 12 1 11 7 11 12 1 11 2
5 4 13 1 12 2
26 13 1 9 16 10 9 1 10 9 2 3 0 2 15 13 1 11 11 1 10 9 1 10 9 11 2
20 1 10 9 1 12 2 13 12 9 2 12 9 7 12 9 13 1 10 9 2
24 15 1 10 0 9 1 10 9 1 11 15 13 2 1 9 2 1 10 9 7 1 10 9 2
23 10 0 9 13 1 10 9 1 9 11 3 13 1 11 2 10 9 16 15 13 1 9 2
7 3 13 3 0 1 11 2
29 16 10 9 13 3 0 2 16 13 1 8 11 2 10 9 1 10 9 7 10 9 1 10 9 15 4 13 0 2
14 15 4 13 10 9 1 13 9 0 1 10 0 9 2
21 11 11 2 8 12 1 11 1 12 2 3 0 1 11 11 13 10 9 0 0 2
13 3 7 15 13 16 11 13 10 9 1 10 11 2
16 9 1 11 11 7 11 11 13 15 1 10 9 1 10 9 2
9 10 0 9 1 13 1 10 9 2
12 10 9 1 9 1 10 9 13 1 9 12 2
27 1 10 9 2 11 13 16 3 3 4 3 9 0 1 11 11 2 10 9 16 15 1 10 9 4 13 2
58 10 9 2 0 1 10 1 10 12 1 11 2 13 9 1 9 0 9 1 9 0 2 9 0 2 9 1 15 9 1 9 2 9 7 9 1 9 0 2 9 1 9 0 1 9 0 2 9 1 9 2 9 1 9 11 7 9 2
8 9 7 9 9 1 12 9 2
13 1 9 2 10 9 13 13 3 10 9 7 9 2
18 10 0 9 16 13 1 10 9 1 10 9 11 11 7 11 11 11 2
16 4 13 1 10 9 0 1 10 9 1 9 2 11 11 11 2
50 1 3 1 12 9 13 1 10 12 7 10 12 1 11 2 10 9 13 1 10 0 9 1 9 1 9 0 2 1 11 2 11 11 2 11 2 11 11 2 11 11 2 7 11 1 11 8 2 11 2
35 15 4 13 1 13 10 9 0 1 9 0 2 11 13 9 1 10 9 1 10 9 7 10 9 1 10 9 2 2 11 13 1 13 9 2
22 11 11 13 10 9 1 10 9 0 3 1 10 9 3 13 3 1 9 1 11 11 2
26 11 2 11 11 7 11 13 13 10 9 0 1 10 9 1 11 16 13 10 9 13 1 10 9 0 2
30 10 9 7 9 1 10 9 13 10 9 1 10 9 7 13 10 9 1 10 9 1 10 9 1 10 9 13 1 15 2
28 10 0 9 13 11 11 11 2 7 13 1 10 9 1 10 9 1 10 11 2 11 11 2 13 1 10 9 2
8 10 9 1 10 9 13 0 2
14 15 13 10 9 3 7 13 0 1 10 9 1 9 2
39 11 2 11 13 10 9 7 9 0 2 13 1 10 9 1 11 2 11 2 9 1 11 2 11 2 1 10 9 1 11 7 9 1 11 2 1 2 11 2
22 10 11 11 1 11 1 10 11 13 10 9 1 9 0 0 1 11 2 13 1 11 2
33 1 10 0 9 13 1 10 9 1 11 11 2 7 1 10 0 9 13 2 15 1 10 9 1 1 10 9 0 2 1 11 11 2
16 1 9 0 1 9 0 3 0 2 1 9 1 0 7 0 2
14 11 11 2 13 10 9 1 9 0 9 1 10 11 2
34 10 9 1 10 9 1 10 11 2 11 11 1 10 11 11 2 13 10 9 0 13 1 10 11 1 1 10 0 0 9 1 10 11 2
52 10 12 9 2 16 13 9 1 10 12 9 1 10 11 11 1 9 2 13 16 10 9 13 10 9 1 10 9 1 10 12 5 2 1 10 16 15 13 1 10 12 9 2 10 9 3 0 1 11 1 12 2
18 10 9 13 10 9 0 1 5 12 9 1 10 5 12 1 10 9 2
12 10 9 1 9 13 1 12 8 5 5 5 2
17 10 0 9 0 4 13 1 9 1 10 9 0 1 11 1 12 2
13 15 13 15 16 15 13 7 3 13 9 1 9 2
32 10 0 9 4 13 10 9 1 3 1 10 9 1 13 1 9 1 10 3 13 0 1 10 9 3 13 1 10 9 1 11 2
36 11 2 15 2 11 13 10 9 7 9 0 2 1 10 9 1 11 2 9 1 11 2 1 10 9 1 11 7 9 1 11 2 1 2 11 2
27 1 9 2 10 9 0 13 1 10 9 7 10 12 1 11 1 12 2 10 9 13 1 0 1 10 9 2
45 2 10 9 3 0 2 1 10 9 2 13 16 4 13 10 9 1 11 1 10 9 2 16 13 9 1 16 4 13 10 9 1 9 2 2 13 11 1 10 9 9 10 11 11 2
8 10 9 1 10 9 13 11 2
37 10 9 11 13 10 9 16 13 1 10 9 0 1 11 2 10 0 9 1 10 9 11 16 13 10 9 1 11 2 11 2 11 2 11 7 11 2
35 15 11 13 10 9 7 9 0 2 13 1 10 9 1 11 2 9 1 11 2 1 10 9 1 11 2 11 2 11 7 9 1 15 11 2
41 10 9 1 15 2 13 12 11 2 13 1 0 9 1 10 11 1 11 2 1 10 13 10 9 2 13 11 11 2 13 1 10 9 7 10 9 0 1 11 11 2
30 10 9 0 11 13 1 10 0 9 10 9 1 10 9 1 12 9 1 10 9 11 11 3 10 0 9 7 11 11 2
47 10 9 1 10 9 0 1 11 7 9 1 10 9 1 10 9 11 2 11 11 2 15 4 13 0 1 13 1 9 2 0 2 10 9 1 10 9 16 10 9 15 13 1 13 10 9 2
6 11 2 11 2 12 2
50 1 10 11 2 7 1 10 0 9 1 11 2 10 9 1 9 0 1 10 9 0 1 10 9 4 3 13 2 1 10 0 9 1 10 15 10 9 13 3 1 10 9 7 3 3 3 1 10 9 2
28 13 10 13 2 9 2 10 16 2 3 2 3 15 13 1 15 16 10 9 13 10 9 1 10 9 3 0 2
18 4 13 1 11 7 3 13 13 16 13 9 1 10 9 1 11 11 2
28 3 2 10 9 13 1 10 9 10 9 1 15 13 10 9 1 9 15 15 13 1 13 7 13 10 10 9 2
13 3 13 9 1 10 9 1 11 11 2 0 9 2
10 10 9 13 3 1 12 7 0 9 2
49 1 16 10 9 0 4 13 1 11 2 11 2 10 9 2 8 2 12 1 11 1 12 2 10 0 9 0 4 13 1 10 9 1 10 11 11 7 13 11 7 11 2 10 9 1 9 3 0 2
24 11 13 10 9 0 1 10 9 1 11 2 1 12 9 5 1 9 7 12 9 2 12 2 2
28 10 9 16 13 1 10 9 1 10 9 0 2 1 10 0 9 15 13 1 15 1 11 1 9 1 10 9 2
50 8 2 10 9 0 2 11 11 2 1 9 2 13 0 3 1 13 10 9 1 10 9 1 9 0 1 10 0 9 1 10 9 1 9 1 10 9 1 11 7 10 9 3 1 15 15 13 10 9 2
29 10 9 1 9 13 16 2 13 1 10 9 1 9 1 10 15 10 9 13 0 9 2 13 10 9 16 13 0 2
37 10 9 13 1 9 9 1 10 9 1 10 9 1 10 9 11 7 1 10 9 1 10 9 11 2 15 13 1 11 1 12 1 9 1 10 9 2
21 10 0 9 13 9 1 9 3 0 7 10 9 2 7 10 9 0 7 12 9 2
37 11 11 2 2 11 2 11 2 13 10 12 1 11 1 12 1 11 2 11 2 13 10 8 9 7 9 1 9 0 16 13 12 9 1 10 11 2
29 2 1 10 9 13 3 1 12 9 16 15 13 1 10 9 7 13 3 12 7 12 15 16 15 13 1 9 0 2
30 13 3 0 1 10 9 1 9 16 13 9 1 10 9 0 1 10 9 1 10 9 2 9 1 10 9 2 0 2 2
19 13 10 12 5 1 9 0 7 10 9 1 12 5 1 9 0 1 9 2
23 3 15 13 1 10 9 11 11 2 13 15 1 4 13 9 16 13 10 9 1 9 2 2
16 3 10 9 13 0 1 10 0 9 2 16 13 3 15 13 2
21 11 4 4 13 3 2 16 10 9 3 15 4 13 1 13 10 9 1 10 9 2
5 11 1 11 11 2
25 1 10 9 1 9 2 10 9 13 1 10 9 7 15 13 1 10 9 13 9 1 10 9 0 2
26 10 9 1 10 9 1 9 13 10 15 0 7 1 10 9 1 9 0 2 10 12 1 12 9 2 2
25 13 0 9 7 13 13 15 10 9 1 10 9 2 3 13 15 3 0 2 13 9 7 15 13 2
58 10 9 1 11 1 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 4 13 1 13 3 0 1 9 1 10 11 2 11 11 2 1 10 9 7 10 9 13 3 0 1 13 0 1 10 9 1 10 10 9 1 9 2
21 11 13 10 9 13 1 10 9 13 1 10 9 1 11 1 10 9 0 1 11 2
26 11 4 13 1 10 9 1 12 7 13 1 9 1 9 1 11 1 11 1 10 9 11 12 1 11 2
28 10 10 9 0 4 13 1 9 11 2 8 2 9 9 2 16 3 4 13 1 10 0 11 2 9 11 2 2
19 10 0 9 0 4 13 1 10 2 11 11 2 2 3 1 10 9 0 2
50 1 9 7 9 0 1 9 1 9 4 13 9 7 9 1 10 9 1 10 9 0 7 10 9 2 9 7 0 9 2 9 0 2 9 1 10 9 2 7 9 1 10 9 0 1 10 9 1 11 2
51 10 9 11 13 3 0 3 2 1 13 9 0 1 0 9 1 9 16 2 13 1 10 9 2 13 10 9 1 9 1 10 9 1 10 11 2 11 2 11 2 2 16 13 9 1 10 9 1 10 11 2
17 3 3 15 13 1 9 1 11 11 2 8 2 2 10 9 0 2
13 13 0 9 1 10 0 9 1 10 9 1 11 2
10 1 10 9 15 13 16 13 1 11 2
18 10 9 15 13 1 9 1 10 9 7 1 10 15 10 9 1 9 2
41 10 9 1 9 2 1 9 2 13 1 10 9 1 10 12 1 10 9 1 9 0 0 2 13 1 9 1 10 9 16 9 1 9 1 9 1 13 1 10 9 2
23 16 15 1 10 12 13 1 9 0 2 4 13 1 9 1 9 0 1 10 9 1 12 2
26 1 9 2 3 1 13 10 9 2 13 10 9 0 7 13 12 9 3 3 2 1 12 9 1 9 2
12 9 1 12 3 15 4 13 1 13 1 12 2
17 11 15 13 1 11 1 13 10 9 7 13 15 1 9 7 9 2
20 15 4 13 0 1 9 1 12 2 12 2 12 7 12 9 1 9 1 9 2
11 15 13 1 11 2 9 1 10 9 11 2
48 10 9 1 12 9 15 13 1 12 2 15 16 13 10 9 1 10 12 5 9 1 10 9 3 7 15 13 3 10 9 1 9 13 1 12 2 1 10 9 1 9 0 1 10 11 1 9 2
21 4 13 1 9 1 12 2 1 9 1 10 9 9 1 10 9 1 9 1 11 2
32 10 9 1 10 11 1 11 16 13 10 9 1 9 1 11 3 13 9 1 9 16 15 4 13 1 13 10 9 1 0 9 2
26 10 9 0 2 16 3 3 13 10 9 1 10 9 1 11 2 15 13 1 10 9 1 9 1 11 2
19 10 9 16 3 13 1 9 13 1 9 0 1 0 9 1 10 9 12 2
32 9 1 15 13 2 1 9 2 10 16 1 3 0 9 11 13 9 1 15 16 2 1 10 9 1 9 2 4 13 10 9 2
54 10 9 1 9 13 1 3 12 1 11 1 10 9 1 9 1 10 11 1 10 11 1 10 9 1 13 1 10 9 16 13 1 10 9 1 10 9 13 1 10 9 0 2 1 9 1 10 9 1 10 9 1 9 2
22 1 10 9 13 9 1 10 9 11 11 2 11 2 11 11 2 11 11 7 11 11 2
11 11 13 9 1 10 9 1 11 11 11 2
23 1 10 9 2 16 13 1 10 0 9 1 9 1 0 9 2 15 13 10 9 1 11 2
27 10 9 12 2 1 9 1 13 9 1 10 9 2 15 13 1 10 9 0 1 11 2 1 10 9 11 2
19 1 9 13 1 10 9 0 1 10 9 11 11 2 11 11 11 11 2 2
14 10 9 1 11 13 10 9 0 1 9 13 1 11 2
27 1 10 9 0 2 0 13 1 10 9 1 11 2 11 7 1 10 9 2 9 13 1 10 9 1 11 2
8 13 3 10 0 9 7 9 2
14 10 0 9 16 15 4 13 1 10 9 1 10 9 2
20 11 11 13 10 9 1 9 1 10 9 1 10 9 1 10 9 1 10 9 2
21 11 13 10 9 1 10 9 1 11 1 10 9 1 11 13 1 10 9 1 11 2
23 10 9 16 13 13 10 9 2 13 1 10 11 1 13 10 9 1 9 3 1 11 11 2
44 10 12 1 11 1 12 2 11 11 2 1 11 1 11 2 9 1 10 9 2 13 1 12 9 1 9 2 15 1 9 7 10 9 0 2 1 11 2 1 9 1 11 11 2
23 1 9 1 10 9 2 10 12 1 11 1 12 15 13 10 9 1 9 0 2 11 2 2
51 3 1 11 2 10 9 0 2 0 3 8 9 15 13 1 9 2 1 10 1 15 1 10 9 1 10 9 1 11 13 1 10 9 0 11 11 7 1 11 11 1 9 0 1 10 9 1 10 0 9 2
28 10 9 13 12 9 3 1 10 9 1 10 9 7 3 13 1 0 9 10 12 1 11 1 10 9 1 9 2
24 1 10 9 1 10 9 2 15 13 9 16 13 9 0 1 9 1 10 11 7 10 0 9 2
29 10 11 13 1 10 9 1 10 9 11 11 3 1 10 9 1 11 1 10 11 2 11 7 11 1 10 11 11 2
17 11 15 13 1 10 9 0 1 10 9 1 9 13 1 10 9 2
38 11 13 1 10 9 1 9 1 10 9 1 10 12 9 2 10 11 11 2 12 2 2 7 3 15 13 9 1 11 7 1 15 16 4 13 1 15 2
14 10 9 1 12 13 12 9 2 1 3 1 10 9 2
22 1 9 3 4 1 13 10 9 1 10 9 1 10 9 1 9 16 7 15 15 13 2
55 4 13 15 1 9 2 8 15 15 13 10 9 0 13 1 9 7 1 9 8 2 9 0 2 12 9 8 13 1 12 9 1 9 2 16 4 13 15 16 13 10 9 0 7 10 9 1 9 1 9 7 9 1 9 2
24 16 4 1 13 10 0 9 1 9 0 2 13 1 11 11 7 13 10 9 1 0 9 0 2
24 10 9 7 9 4 13 1 11 1 12 2 10 0 9 4 13 1 10 9 0 1 9 0 2
12 2 15 13 13 15 1 10 9 1 11 11 2
40 1 15 13 1 16 4 7 2 13 3 2 2 7 13 16 10 9 15 13 3 1 15 1 10 0 9 11 11 1 3 1 9 2 9 1 9 7 9 0 2
30 3 2 10 9 15 13 1 0 9 1 10 9 1 10 9 1 10 9 0 2 1 3 1 11 2 11 11 7 11 2
28 1 15 9 2 10 9 13 9 1 10 9 1 9 2 16 3 3 13 2 3 0 13 15 2 7 10 9 2
27 3 13 10 0 9 1 9 1 11 7 10 9 11 1 10 9 1 11 2 1 0 9 1 10 9 0 2
45 10 11 12 2 11 12 8 1 12 2 2 13 1 11 11 1 11 12 2 13 10 9 1 10 9 8 1 9 0 13 1 13 1 10 11 12 7 13 1 12 7 12 1 11 2
27 13 1 11 13 1 10 9 1 10 9 1 10 0 9 16 13 3 0 1 10 9 9 1 10 9 0 2
20 3 2 10 9 13 1 10 9 2 8 2 1 11 2 1 10 9 1 11 2
16 11 13 10 9 1 9 0 2 0 1 10 9 1 10 9 2
36 1 10 9 1 13 10 9 7 13 1 10 9 10 9 1 10 9 2 1 10 9 10 9 16 15 13 1 10 9 13 9 0 1 15 13 2
13 1 9 1 10 9 2 10 9 4 13 1 12 2
9 1 10 9 2 15 13 10 9 2
16 1 9 1 10 9 10 12 5 13 9 7 9 1 10 9 2
74 10 12 9 0 1 9 0 15 13 1 11 2 9 0 2 1 10 12 7 10 12 1 11 7 1 11 2 9 0 7 1 9 2 1 10 12 7 10 12 1 11 1 12 1 10 9 1 10 9 0 1 9 1 9 2 11 2 2 10 9 0 1 9 1 9 7 10 9 0 1 9 1 9 2
71 1 10 12 1 10 9 2 1 10 9 13 1 10 9 0 2 10 9 1 10 11 11 11 7 11 11 13 1 9 1 10 9 1 9 0 2 11 11 2 10 9 1 9 1 9 0 2 11 11 7 10 9 1 10 9 0 1 10 9 2 11 11 11 2 10 9 1 10 9 0 2
13 10 9 13 10 9 1 11 2 1 3 12 9 2
28 7 3 10 9 4 13 3 2 4 13 1 10 9 0 7 10 9 0 1 10 9 2 1 9 1 10 9 2
18 10 9 1 2 11 2 13 3 10 9 1 10 9 0 2 11 2 2
22 1 12 2 10 9 11 11 13 10 9 7 15 13 1 11 11 2 1 11 11 11 2
36 1 12 1 12 2 1 10 9 14 2 0 1 8 2 11 15 13 1 10 9 1 11 2 1 10 11 0 2 3 13 1 13 10 9 0 2
4 2 15 13 2
19 10 9 13 16 10 12 1 11 8 11 11 1 11 1 11 11 11 11 2
31 11 11 2 12 1 11 1 12 2 13 10 9 7 9 0 13 1 10 13 2 9 0 2 1 10 9 1 12 7 12 2
15 3 1 10 9 15 13 9 1 9 1 10 10 9 0 2
19 4 13 1 10 9 0 0 2 1 1 10 9 0 0 1 10 9 0 2
20 4 13 1 9 1 3 2 7 13 1 10 11 7 8 11 1 11 1 12 2
34 11 2 1 10 9 1 13 1 10 9 3 0 16 13 1 10 9 2 10 9 2 7 1 0 10 11 2 16 13 0 10 10 9 2
46 16 13 10 9 0 1 11 2 8 2 2 9 1 10 9 2 10 9 15 4 13 1 10 9 1 10 9 1 10 16 10 9 0 13 10 9 2 13 1 12 9 2 1 10 8 2
36 1 10 9 1 10 0 9 2 10 9 0 15 13 1 13 10 9 1 10 9 2 3 16 10 9 3 4 4 3 13 3 1 10 9 0 2
29 10 9 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 11 2 11 11 2 11 11 11 2
18 11 13 10 9 1 10 9 1 11 1 10 9 1 11 2 1 11 2
21 13 1 10 0 9 1 10 9 2 3 4 13 15 15 1 10 9 1 12 9 2
11 13 1 9 7 10 0 9 13 11 11 2
14 12 9 4 13 3 1 9 0 2 16 3 4 13 2
32 1 10 9 2 11 13 1 13 1 10 9 13 13 1 11 1 10 9 7 3 13 1 11 7 11 15 13 1 13 10 9 2
15 3 13 0 1 13 13 10 9 1 10 9 1 9 0 2
60 10 9 0 4 13 1 10 9 0 1 10 9 1 10 9 1 9 0 2 10 9 0 4 13 1 10 9 0 1 10 9 1 10 9 2 1 9 0 7 3 1 10 9 0 1 9 0 2 10 9 0 4 13 1 10 9 1 10 9 2
40 11 11 15 13 1 10 9 1 9 13 9 1 9 2 0 2 0 7 0 2 16 13 10 0 9 1 9 7 9 0 15 1 10 9 7 1 10 9 13 2
20 10 9 13 10 9 0 7 10 9 3 0 3 10 9 4 13 1 10 9 2
10 15 13 9 10 9 1 10 0 9 2
26 10 9 11 11 11 11 13 1 10 9 1 10 9 11 1 10 9 13 1 9 1 10 9 1 11 2
19 1 10 9 13 10 9 1 9 2 10 9 1 10 9 16 13 1 11 2
34 1 9 2 11 13 16 3 13 9 1 10 9 3 1 10 9 1 9 0 16 13 16 10 0 9 1 10 9 13 1 9 1 11 2
42 11 7 11 4 13 11 2 1 10 9 1 9 1 9 0 7 2 3 3 10 0 9 2 10 9 0 2 13 7 13 1 11 7 11 11 2 4 13 1 10 9 2
24 10 9 1 10 11 1 11 7 11 13 10 9 2 4 13 10 9 1 10 11 0 3 3 2
29 1 10 0 9 2 11 15 13 1 15 1 10 3 0 9 0 1 10 11 11 2 3 13 10 0 9 1 9 2
34 3 15 2 10 9 1 11 15 13 1 10 9 0 3 1 10 11 1 11 11 2 13 1 10 11 1 10 11 1 11 11 1 12 2
38 3 2 10 9 13 10 9 1 9 0 7 0 2 1 15 15 13 10 9 1 10 10 9 16 13 10 11 11 1 10 11 11 2 11 7 11 2 2
24 10 9 1 9 1 10 9 0 15 13 1 10 9 1 11 11 2 11 11 1 10 11 2 2
39 10 9 0 3 4 13 1 10 0 11 11 2 16 4 13 11 11 2 7 1 11 7 10 9 16 13 1 10 0 9 0 1 13 15 2 9 0 2 2
11 10 9 1 10 9 13 10 9 1 9 2
30 10 11 2 1 9 2 7 11 1 11 2 2 3 2 10 9 0 2 13 15 1 10 12 9 1 11 1 10 9 2
17 10 10 9 2 3 10 3 0 2 4 13 15 1 9 3 0 2
49 10 9 1 9 7 9 2 1 12 2 12 9 1 9 0 7 0 2 16 10 9 13 1 3 1 12 1 12 1 10 9 2 4 13 2 10 9 3 4 13 7 13 7 10 9 13 7 13 2
23 10 12 5 1 10 10 9 13 10 0 9 7 10 12 5 13 3 9 0 1 12 9 2
35 10 10 4 4 13 1 10 9 0 2 7 10 12 9 0 8 2 12 1 10 11 13 1 10 9 2 1 3 16 10 9 15 13 2 2
17 10 9 15 13 1 15 1 10 9 0 16 13 3 1 10 9 2
80 10 9 13 9 1 10 9 0 7 1 10 9 0 1 10 9 2 9 2 9 1 10 9 1 9 0 1 11 7 9 1 9 0 2 9 1 9 1 9 0 7 9 1 10 9 2 9 1 9 2 9 1 9 1 9 1 9 0 7 9 1 9 1 9 1 9 0 2 15 13 1 9 2 9 0 2 0 7 0 2
12 11 13 10 9 1 10 11 1 10 9 0 2
11 11 13 1 11 13 15 1 13 1 11 2
34 11 11 11 2 13 10 12 1 11 1 12 1 11 11 2 13 10 11 0 1 11 11 16 13 1 10 9 1 10 11 1 11 11 2
17 10 9 0 1 10 9 13 10 9 13 1 10 9 7 10 9 2
7 1 15 15 13 9 0 2
21 4 13 10 1 10 11 11 1 10 9 11 11 7 1 10 11 11 1 11 11 2
8 13 9 3 7 3 3 0 2
6 4 13 3 1 11 2
41 10 9 1 10 9 13 13 1 11 1 9 0 7 13 9 0 1 10 11 2 13 10 9 1 10 9 1 9 2 3 1 9 1 9 0 2 0 2 7 0 2
19 13 3 10 9 3 0 1 10 9 1 11 7 4 13 1 9 0 0 2
37 16 1 10 9 13 0 16 13 1 10 9 2 12 2 10 0 9 7 10 9 1 10 11 11 13 10 9 1 10 9 3 1 3 12 9 0 2
19 10 9 13 13 10 9 7 13 1 10 9 0 10 9 0 1 10 9 2
23 3 4 13 1 13 10 9 1 9 1 10 11 11 1 11 1 12 15 4 13 1 11 2
51 1 9 2 10 9 1 11 4 13 3 1 11 1 10 0 9 1 10 8 2 13 16 3 1 10 9 10 9 15 13 1 9 0 7 13 10 9 1 9 0 7 1 9 16 4 13 1 10 9 12 2
24 15 4 13 3 0 1 10 9 1 13 9 7 1 13 10 0 9 1 9 16 15 13 9 2
14 1 0 9 2 10 11 1 10 9 3 13 3 0 2
20 10 9 1 10 9 13 0 7 0 2 7 3 13 0 7 13 1 10 9 2
13 3 13 9 13 1 10 9 7 1 10 9 0 2
61 11 13 10 9 1 10 9 1 10 9 7 10 9 0 1 10 9 1 10 11 11 1 10 9 1 11 11 2 3 9 2 9 2 9 2 9 1 9 1 9 2 9 7 9 1 0 13 1 9 1 0 9 7 0 13 1 13 10 9 0 2
24 10 9 13 1 10 9 1 10 9 13 2 13 15 16 15 13 2 1 10 9 9 7 9 2
16 13 16 15 13 0 3 1 10 0 9 7 1 10 9 0 2
37 10 9 0 13 16 10 9 0 13 1 10 12 5 1 12 2 1 10 12 5 1 10 9 0 7 16 13 1 10 9 1 10 12 5 1 12 2
18 1 9 1 10 9 1 12 2 10 9 4 13 1 9 0 7 0 2
38 10 9 0 0 13 10 9 16 15 13 13 1 10 0 9 2 1 0 9 13 9 1 10 9 1 10 9 7 1 0 13 15 1 10 9 1 9 2
44 10 0 9 3 13 0 9 2 13 10 9 1 10 9 1 10 9 7 10 9 1 10 9 0 2 13 3 0 10 9 2 10 9 2 10 9 2 10 9 2 10 9 0 2
19 15 13 9 1 10 8 1 10 9 1 9 7 3 9 1 10 9 0 2
31 13 13 0 1 10 9 2 3 0 1 3 1 10 0 13 10 0 9 1 9 7 2 1 9 1 8 2 13 1 9 2
31 13 1 10 11 1 11 11 2 11 11 11 2 11 1 11 11 2 7 1 10 11 11 2 11 2 11 2 7 10 11 2
50 1 10 9 0 2 10 9 4 13 1 9 1 10 9 0 2 13 1 0 9 1 11 16 13 10 9 1 10 12 9 1 10 9 7 13 0 9 1 10 9 13 1 9 0 1 10 11 1 11 2
20 13 1 10 9 1 11 1 11 2 1 10 9 1 11 2 11 2 11 2 2
31 1 0 9 2 3 15 13 10 9 1 15 1 10 9 2 10 9 13 10 0 9 1 9 15 4 13 3 1 10 9 2
28 15 13 1 9 0 2 10 12 1 11 1 12 2 11 11 0 1 10 9 11 11 2 11 11 7 11 11 2
13 1 10 9 1 12 2 13 12 9 13 1 11 2
53 10 9 1 10 9 2 16 13 1 10 3 0 9 0 1 10 9 2 13 15 1 11 1 11 2 15 16 2 3 2 15 4 1 13 16 0 9 3 13 1 9 1 10 0 9 2 7 1 9 1 10 9 2
30 10 12 1 11 1 12 4 13 10 16 13 9 1 10 9 2 11 11 11 11 2 1 10 11 1 9 0 7 9 2
22 1 11 1 12 2 10 9 13 11 1 10 9 1 13 10 9 13 1 10 11 11 2
90 11 13 2 1 12 2 16 10 9 0 3 4 13 7 13 13 1 10 9 1 15 1 10 9 1 10 9 2 1 11 2 1 15 3 0 2 1 11 2 1 15 3 0 2 2 1 11 2 1 10 9 1 15 9 1 9 1 9 2 1 11 2 1 10 9 1 10 9 1 9 1 15 0 2 2 1 11 2 1 10 9 2 1 11 2 1 10 9 2 2
29 2 10 9 0 13 10 0 9 1 10 9 16 3 4 13 15 3 3 1 15 3 9 2 2 15 13 10 9 2
46 10 9 1 10 9 1 10 9 13 10 9 10 9 16 13 0 2 13 10 9 2 10 9 7 10 9 2 3 3 13 1 9 10 9 1 10 0 9 7 1 15 2 10 9 0 2
26 13 10 0 9 1 11 1 4 13 3 1 10 9 0 1 10 11 11 2 10 12 1 11 1 12 2
21 4 13 1 10 9 1 11 11 1 10 11 1 11 2 16 4 13 1 10 12 2
31 1 10 9 0 2 3 13 9 2 9 2 9 7 9 13 3 0 16 15 13 10 9 7 1 11 13 1 10 9 11 2
32 10 9 11 11 13 10 9 3 3 1 13 9 1 10 11 11 16 4 13 1 10 9 10 11 11 7 15 13 10 0 9 2
25 11 11 13 10 9 1 9 0 13 1 10 9 1 10 9 16 15 13 15 3 1 10 0 9 2
18 10 9 2 11 11 2 4 13 1 10 9 2 11 11 11 12 2 2
35 10 9 13 1 9 0 2 15 13 1 10 9 1 10 9 1 10 9 7 3 13 9 1 10 9 7 9 1 13 16 10 9 15 13 2
42 10 9 1 9 13 1 9 1 9 1 12 1 3 9 2 13 1 16 15 3 13 1 10 9 1 10 9 2 3 13 1 9 1 10 9 7 1 10 9 1 10 9
40 3 2 11 11 2 9 1 11 1 11 2 13 10 9 1 10 2 11 11 12 2 2 0 1 10 0 9 1 10 11 11 2 9 7 9 0 1 10 9 2
12 13 1 11 2 11 2 11 7 10 9 0 2
18 11 11 13 10 9 13 1 10 9 1 11 1 10 9 0 1 11 2
35 1 10 0 9 13 1 10 2 11 11 8 11 2 2 9 0 1 9 2 1 11 2 13 15 1 10 12 0 9 2 0 1 11 11 2
29 10 9 1 10 9 1 9 15 13 1 10 0 9 2 3 13 10 0 9 1 9 1 0 9 1 10 9 9 2
13 10 9 1 9 13 1 10 12 7 12 1 12 2
18 1 12 13 9 1 11 1 11 7 2 3 2 4 13 10 9 0 2
12 11 15 13 1 10 9 13 1 10 12 9 2
45 10 9 13 10 0 9 1 10 9 1 10 9 12 1 10 11 2 9 1 10 11 11 1 11 2 16 13 1 10 9 1 9 0 1 10 9 0 1 9 16 11 13 1 9 2
14 3 2 13 1 9 7 13 10 9 0 16 10 9 2
33 10 12 1 11 1 10 9 2 16 13 1 9 1 10 11 13 10 9 1 13 10 11 11 1 10 9 11 2 11 13 1 11 2
36 1 10 0 9 2 1 13 16 10 8 13 1 0 1 10 9 0 2 2 3 1 11 2 10 9 13 3 9 2 7 1 0 15 13 9 2
37 7 15 1 15 9 13 1 15 15 13 3 7 4 13 1 10 9 1 11 11 8 2 7 10 9 7 10 9 15 4 13 1 10 9 3 13 2
5 13 1 10 11 2
10 13 10 0 9 1 10 11 11 11 2
7 3 2 15 13 1 15 2
24 10 9 13 1 13 2 7 1 12 15 13 10 9 1 3 1 10 12 5 1 9 1 12 2
30 1 9 1 11 11 11 13 0 13 3 0 9 2 1 10 9 0 2 3 1 9 12 11 7 9 11 11 11 2 2
5 10 9 4 13 2
21 10 9 1 11 11 2 0 1 11 2 13 10 9 1 10 12 1 9 7 9 2
39 7 15 7 11 15 13 9 1 16 3 3 13 9 1 13 11 2 3 1 16 15 13 16 11 13 0 7 10 9 1 10 9 13 3 16 13 1 11 2
35 10 9 13 1 0 9 1 10 9 7 4 13 3 0 9 1 10 9 2 13 10 9 16 3 13 10 9 1 10 9 7 10 9 13 2
34 2 1 10 9 0 2 10 0 11 2 1 10 9 0 2 10 9 2 7 10 9 1 11 3 15 13 15 7 15 2 2 13 11 2
32 3 2 10 9 1 9 1 10 11 13 1 9 1 10 9 1 10 9 16 13 10 9 1 10 0 9 1 13 9 7 9 2
45 1 12 2 10 9 0 11 11 13 1 11 11 1 10 9 12 1 10 9 1 10 12 0 9 1 10 10 9 2 7 1 12 10 9 4 13 1 10 9 11 1 10 9 0 2
61 10 9 11 11 2 9 1 11 1 10 11 1 10 11 1 11 10 12 1 11 1 12 2 13 16 10 9 13 10 9 1 13 0 2 1 15 15 13 10 9 1 10 9 1 11 2 3 15 13 10 9 0 0 7 10 9 1 9 1 9 2
43 1 10 9 1 10 9 1 10 11 11 2 10 9 13 10 9 0 1 12 5 5 2 1 10 15 12 5 5 13 1 9 0 7 2 12 5 2 12 5 5 13 9 2
15 3 4 13 10 0 9 1 9 0 13 16 3 13 9 2
32 1 10 9 1 10 9 1 12 2 10 9 0 1 9 1 10 9 13 1 9 12 2 7 10 9 0 1 9 13 9 12 2
25 1 12 2 13 1 10 9 10 11 8 11 7 15 13 1 10 9 1 10 9 2 11 11 11 2
34 10 9 5 1 10 9 1 11 11 2 13 10 12 1 11 1 12 2 15 13 1 15 9 1 12 9 1 10 9 11 2 11 11 2
5 9 1 12 9 2
29 11 11 15 13 10 0 9 1 12 9 2 1 12 1 10 12 2 13 9 1 10 9 1 11 1 10 9 12 2
25 10 0 9 15 13 16 11 4 13 1 12 3 1 12 9 1 9 1 10 9 1 11 1 9 2
13 13 1 10 0 9 2 16 13 10 9 1 0 2
16 15 0 2 1 10 13 15 13 10 9 13 10 9 3 0 2
16 10 9 1 9 1 9 13 13 1 10 9 7 1 10 9 2
28 13 1 11 9 7 4 13 10 9 0 1 3 3 2 13 7 3 13 1 11 7 3 13 9 3 1 11 2
13 11 4 13 1 11 11 1 10 9 13 1 11 2
15 3 0 3 10 9 7 10 9 15 13 1 10 0 9 2
20 11 13 1 12 7 12 1 9 1 10 9 1 10 11 11 1 10 11 11 2
24 4 13 10 11 1 11 1 10 0 9 7 4 13 1 10 9 1 10 9 7 1 10 9 2
7 10 9 11 13 1 12 2
22 15 13 1 9 0 13 1 16 10 9 13 10 9 0 1 10 13 10 9 1 9 2
36 10 9 11 11 13 10 10 9 1 9 1 9 1 9 1 3 1 12 9 1 9 1 10 9 13 10 9 1 9 1 11 11 11 1 12 2
28 16 13 10 9 0 13 0 15 13 10 0 9 7 15 13 15 16 15 4 13 1 13 16 15 13 10 9 2
39 10 9 13 0 1 10 9 1 11 2 3 1 10 11 1 10 11 2 1 10 9 1 11 2 3 1 10 9 2 1 10 0 9 0 7 9 1 9 2
23 10 9 1 10 9 13 13 10 9 0 16 13 1 11 11 2 16 13 1 10 9 12 2
45 3 1 15 2 13 10 9 1 9 1 11 2 7 13 1 10 9 1 16 10 12 5 1 10 9 4 13 1 9 1 10 9 2 3 3 1 10 12 5 2 13 1 10 9 2
22 3 2 13 10 9 1 11 1 12 1 10 9 1 10 2 9 1 10 9 0 2 2
8 1 10 11 3 13 10 9 2
21 1 10 9 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 5 5 2
51 10 0 9 2 13 1 10 9 1 9 1 10 9 2 7 1 3 10 9 0 1 11 2 13 3 1 9 1 9 0 1 10 9 13 3 1 10 9 1 10 9 1 10 11 7 10 0 9 1 11 2
23 1 3 13 10 9 1 10 9 0 11 11 2 10 9 15 13 1 10 11 1 11 11 2
16 10 9 1 11 13 10 9 1 10 9 1 10 11 1 11 2
25 1 10 9 1 9 2 9 0 7 9 2 2 10 9 0 13 1 13 0 1 10 9 7 9 2
13 10 9 13 0 9 2 1 10 0 7 10 9 2
39 16 15 4 13 16 11 11 13 9 1 11 2 1 9 13 10 9 3 13 2 16 13 9 13 9 1 11 7 16 4 1 13 1 9 1 15 1 15 2
7 9 1 11 11 1 11 11
35 1 13 10 9 2 15 13 10 9 1 10 9 1 10 9 1 13 7 13 1 9 10 9 2 3 7 1 10 9 1 9 1 10 9 2
21 11 2 1 0 9 0 2 9 1 9 0 1 10 9 1 10 9 7 10 9 2
30 11 3 13 10 11 1 11 1 12 2 10 11 11 1 12 7 10 11 1 11 1 10 11 1 10 11 11 1 12 2
27 1 12 10 9 1 10 9 15 13 10 11 11 11 1 9 1 10 9 1 10 9 1 10 9 0 0 2
24 1 10 9 2 13 1 10 2 9 0 1 9 2 7 1 10 2 9 0 7 0 11 2 2
17 10 9 9 13 10 9 1 11 2 16 13 10 9 1 10 9 2
10 4 1 13 16 13 1 10 9 0 2
28 10 9 1 10 9 11 2 10 9 13 0 1 10 9 0 1 10 9 2 15 13 1 10 9 1 10 9 2
42 10 9 1 10 9 1 11 1 9 1 10 0 9 1 9 13 1 10 3 0 9 16 15 13 10 0 9 7 9 7 16 13 10 0 9 1 10 9 1 10 9 2
43 10 9 13 3 1 12 12 9 0 2 0 7 0 1 10 9 0 2 3 1 16 13 9 1 9 2 9 1 9 1 9 7 10 15 13 1 9 0 2 0 7 0 2
8 3 15 13 1 3 12 9 2
28 15 13 1 9 2 1 10 15 10 3 0 13 11 11 2 9 7 11 11 2 3 1 10 0 9 2 11 2
34 4 13 15 1 10 0 9 2 3 16 3 13 15 16 3 15 13 2 3 1 10 9 1 10 9 2 7 1 10 9 1 10 9 2
20 10 9 0 1 11 13 1 12 5 9 1 10 9 7 12 5 9 1 11 2
27 11 15 13 9 1 16 3 13 13 10 9 3 1 11 11 2 13 1 10 9 7 13 10 9 1 11 2
13 10 9 1 9 13 1 12 9 2 2 5 5 2
29 10 9 1 11 13 13 11 1 10 9 16 13 10 9 1 10 9 7 13 3 1 9 1 9 10 9 1 11 2
29 10 9 4 13 15 1 9 2 9 2 9 7 9 7 4 13 1 10 9 0 2 1 10 9 1 10 9 0 2
28 10 15 16 4 13 13 11 11 1 10 11 16 13 10 9 7 13 13 1 9 7 9 0 2 13 9 2 2
30 10 9 13 10 9 2 7 1 10 9 1 10 9 2 3 1 10 9 1 10 9 2 1 10 16 7 3 4 13 2
13 3 2 1 10 12 9 1 13 3 15 4 13 2
42 1 12 9 1 9 2 10 11 11 4 13 1 10 9 10 9 1 13 10 9 1 0 9 1 10 9 0 1 10 9 2 1 13 1 13 1 10 9 1 9 0 2
20 1 9 2 10 9 1 11 7 11 2 16 3 13 10 9 2 13 15 0 2
16 15 13 10 0 9 16 13 16 1 10 9 1 9 4 13 2
22 11 13 10 9 1 9 1 10 9 11 1 10 9 11 16 15 13 1 9 1 11 2
23 1 10 9 2 10 9 1 10 9 15 13 1 10 9 11 11 11 5 12 2 1 11 2
16 10 0 9 2 11 11 2 11 2 8 2 13 0 1 11 2
17 15 4 13 16 13 9 0 1 15 1 10 9 7 10 9 0 2
13 3 15 13 1 10 9 0 7 10 9 1 9 2
22 1 10 9 13 15 9 7 3 13 1 10 9 13 16 10 9 1 10 11 15 13 2
63 1 10 9 15 11 7 11 13 13 15 13 10 9 1 11 7 10 9 16 13 1 10 9 15 13 16 15 15 13 1 10 9 2 15 1 10 12 13 15 16 13 10 9 1 10 9 1 9 2 9 7 9 16 13 10 9 2 10 9 13 7 13 2
7 13 1 10 9 1 12 2
47 13 1 10 9 1 10 9 0 1 13 10 9 3 0 7 0 2 10 9 13 1 13 9 1 10 9 1 7 4 2 1 9 1 10 9 2 13 10 9 7 13 9 1 10 0 9 2
26 3 2 1 12 2 11 11 2 10 9 13 1 11 11 2 4 13 1 11 11 10 15 13 1 12 2
25 13 3 2 7 1 3 10 9 1 10 9 10 9 3 13 10 9 1 10 0 9 1 10 9 2
18 13 1 12 9 2 12 1 11 2 9 7 10 9 1 11 7 11 2
10 10 0 9 0 13 10 9 1 11 2
14 11 11 11 13 13 1 9 0 1 10 11 1 11 2
13 10 9 1 10 9 0 13 1 12 9 1 9 2
42 11 11 13 2 1 1 9 2 1 10 9 2 7 9 1 10 9 2 1 15 2 12 9 0 7 0 1 13 15 16 10 9 1 9 0 13 13 3 3 2 13 2
21 1 10 9 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 5 8 2
34 10 0 9 1 10 9 15 13 1 10 9 1 9 0 7 0 2 3 7 1 10 0 9 1 0 9 0 1 10 9 1 10 9 2
16 11 1 11 1 11 13 10 0 9 1 9 1 10 9 12 2
18 3 13 1 10 9 1 10 9 11 11 2 13 10 9 1 10 11 2
74 10 11 1 11 0 2 9 2 0 7 9 0 1 10 11 11 11 11 11 2 15 13 13 1 10 9 1 11 11 1 10 11 2 11 2 13 10 9 0 13 1 12 2 16 13 10 9 0 1 10 9 0 1 10 9 0 2 0 2 0 7 1 9 0 2 1 9 1 9 0 7 9 0 2
25 10 9 9 15 13 1 10 12 7 12 9 1 9 7 10 9 9 15 13 10 9 1 10 11 2
31 15 15 4 13 3 1 10 15 1 10 9 1 11 7 13 3 0 1 15 1 11 2 16 3 3 13 0 1 9 0 2
11 10 9 13 9 13 1 10 9 0 0 2
30 13 15 1 10 9 1 10 11 11 2 15 4 13 1 11 11 1 10 9 1 13 1 10 9 1 10 9 1 11 2
16 1 10 11 1 12 2 13 12 9 13 1 10 9 1 11 2
13 11 2 11 3 4 13 9 1 10 9 1 11 2
26 3 3 10 9 1 10 11 4 13 1 13 1 10 11 2 7 3 15 13 1 12 9 2 1 12 2
35 3 1 11 13 16 3 7 3 10 9 1 10 11 13 1 9 0 2 1 9 16 4 13 1 10 0 9 11 7 13 1 10 9 11 2
5 13 10 9 9 2
40 9 2 9 1 9 2 9 7 9 13 1 9 7 9 1 9 1 10 0 9 16 13 1 10 9 2 3 9 1 11 7 11 4 4 3 13 1 10 9 2
23 3 3 2 4 13 15 9 0 1 9 16 3 15 13 1 13 10 9 1 10 11 12 2
43 11 13 10 9 2 13 10 9 1 13 10 9 7 4 13 10 15 13 16 13 1 10 9 2 7 11 12 3 15 13 10 9 3 16 13 11 10 12 1 11 1 12 2
43 10 9 1 3 1 12 9 0 2 3 1 10 9 2 13 1 10 9 0 1 9 0 16 13 10 9 1 10 9 0 2 16 4 13 3 10 9 1 9 2 11 11 2
14 1 10 9 12 2 13 1 9 8 1 11 11 11 2
27 11 2 10 2 11 13 10 0 9 1 10 9 0 7 15 13 1 13 7 13 10 9 0 1 10 9 2
20 1 12 13 1 13 1 10 11 1 11 11 2 3 13 9 1 10 9 11 2
51 3 7 13 10 9 13 1 10 9 1 16 3 10 9 3 13 10 9 7 15 13 10 9 1 10 9 2 7 16 10 9 13 10 9 7 13 15 16 13 10 9 1 10 9 2 7 3 15 13 9 2
7 15 13 1 10 9 0 2
13 10 9 1 9 13 1 12 9 2 2 9 5 2
23 10 12 1 11 1 12 13 1 0 9 1 10 0 9 1 10 11 1 10 11 1 11 2
8 3 13 10 9 0 7 0 2
37 10 9 0 13 13 1 10 9 16 10 9 13 0 2 16 1 10 9 13 13 15 1 10 9 13 10 9 1 10 9 1 13 15 1 10 9 2
20 15 13 1 10 9 1 10 9 2 10 9 0 2 10 9 2 7 10 9 2
26 1 10 9 1 10 9 1 11 1 10 9 2 11 13 16 11 11 13 10 9 3 1 10 9 11 2
47 11 2 15 13 3 1 10 9 1 11 2 3 15 13 1 10 9 11 11 2 10 15 15 13 1 13 1 0 9 1 10 9 1 10 9 11 11 2 13 10 8 1 10 10 9 12 2
21 13 9 1 10 9 1 10 9 13 15 1 10 9 16 15 13 1 10 11 12 2
45 15 16 13 1 10 9 13 16 11 15 13 1 10 9 2 3 16 10 9 13 10 9 1 11 7 11 15 15 13 1 10 9 9 1 10 0 9 3 1 13 10 9 1 9 2
20 11 2 3 2 2 11 2 15 2 2 11 2 1 15 2 2 11 2 7 2
63 10 0 9 0 2 16 1 10 9 13 10 0 9 0 1 9 1 11 2 3 13 1 10 9 16 13 10 9 7 4 1 13 16 1 10 0 9 1 10 9 2 10 16 13 10 9 1 3 2 13 10 9 16 13 15 10 9 7 13 3 0 3 2
21 7 3 2 15 13 9 0 1 10 9 3 0 7 0 16 3 13 10 9 0 2
64 10 9 1 10 11 1 11 2 10 11 2 11 11 2 4 13 16 16 3 13 1 10 9 1 9 1 10 9 0 2 11 11 1 11 2 10 9 2 9 2 13 1 10 9 1 9 13 1 9 2 1 10 0 9 1 10 9 2 10 9 11 11 11 2
45 10 9 12 1 10 9 1 11 13 16 10 9 4 13 1 10 9 1 10 9 11 2 16 13 1 11 11 1 10 11 2 7 3 1 3 1 12 9 2 12 9 2 1 11 2
29 1 10 9 0 1 10 9 13 12 9 0 7 15 0 1 9 0 15 13 1 10 9 1 3 2 1 10 9 2
49 9 11 12 2 13 1 12 9 7 16 4 13 1 12 1 12 12 9 2 13 15 1 10 9 1 10 11 11 11 2 11 11 1 9 1 10 9 7 9 0 16 15 13 13 1 10 10 9 2
57 1 10 9 4 13 1 10 9 10 9 1 10 9 11 2 13 1 10 9 0 2 16 1 10 0 9 13 10 9 0 0 1 10 9 2 10 15 13 3 0 1 10 9 0 16 4 13 1 10 9 1 10 9 0 3 13 2
12 13 10 9 1 9 3 0 2 0 7 3 2
19 10 9 1 10 9 13 10 9 3 0 2 9 0 7 9 1 0 9 2
16 1 9 1 10 9 10 12 5 13 0 7 9 1 10 9 2
12 11 11 13 7 15 13 3 13 10 9 0 2
36 10 9 3 0 2 1 10 9 1 10 11 2 10 9 11 7 10 9 1 10 11 15 13 1 9 1 10 0 7 0 9 2 13 15 3 2
22 1 12 15 13 1 10 0 9 1 10 9 1 11 9 1 10 9 1 9 1 9 2
40 11 2 11 2 11 13 10 9 7 9 0 2 13 1 10 9 1 11 2 11 2 9 1 11 2 1 10 9 1 11 2 9 2 11 7 9 1 15 11 2
15 13 9 2 0 7 9 0 1 11 11 11 1 10 11 2
12 1 10 0 9 15 13 10 9 1 10 11 2
12 11 11 13 10 9 1 9 1 10 9 11 2
29 13 10 9 1 9 1 10 9 3 0 2 11 2 1 10 15 13 10 0 9 13 1 10 0 9 7 10 9 2
16 3 1 10 12 5 1 10 9 13 1 10 9 1 9 0 2
7 2 13 10 0 1 11 2
25 13 10 9 1 10 9 12 2 12 2 12 2 12 2 12 7 12 2 3 7 10 9 13 11 2
20 10 9 13 1 12 9 0 16 13 1 13 9 7 13 9 1 9 1 0 2
16 1 10 0 9 2 10 9 1 9 13 13 7 13 1 11 2
22 10 0 9 13 10 12 2 1 10 15 13 12 9 2 12 9 7 12 9 1 9 2
40 1 10 9 1 9 1 11 11 2 10 9 1 10 9 3 13 0 2 16 15 13 10 9 1 13 9 2 1 10 9 16 13 10 9 2 7 3 13 2 2
55 1 0 9 11 15 13 1 13 1 10 9 1 10 9 2 7 15 15 13 10 12 9 1 10 9 1 10 9 1 11 11 1 9 1 10 11 11 2 13 1 10 9 1 11 7 13 10 9 1 9 1 10 11 11 2
32 1 10 9 1 11 1 10 12 1 11 7 1 11 11 2 10 12 1 11 1 12 2 11 13 10 9 1 10 9 1 11 2
33 10 9 1 10 15 10 9 0 4 13 13 7 13 10 9 1 9 2 9 1 9 7 9 2 13 0 1 15 1 10 9 0 2
47 11 1 11 2 11 11 1 3 1 12 9 4 13 10 11 11 1 10 0 9 1 9 0 2 10 9 15 15 13 1 9 0 2 0 7 0 2 10 9 15 15 13 10 11 1 9 2
42 11 13 10 9 0 0 1 9 0 0 7 9 11 0 2 4 13 15 1 9 1 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 11 11 7 11 11 2
29 11 13 10 9 7 9 0 2 13 1 10 9 1 9 2 9 1 11 2 1 10 9 1 11 7 9 1 11 2
22 1 10 11 11 15 15 13 10 9 0 7 10 10 9 4 13 1 10 9 1 9 2
22 9 1 10 9 11 2 10 9 13 15 3 0 1 13 10 9 1 10 10 10 9 2
31 1 10 9 1 10 9 11 1 10 9 1 11 1 11 10 12 1 11 1 12 2 4 13 1 10 9 1 10 9 0 2
24 13 1 10 9 1 7 13 10 9 1 10 9 16 13 1 13 10 9 1 11 1 10 9 2
24 10 9 0 1 9 2 1 13 15 1 10 9 7 1 10 9 7 1 10 9 7 10 9 2
31 0 2 0 2 0 2 0 2 15 13 10 9 1 13 15 16 4 13 10 9 1 11 2 15 16 13 3 3 1 11 2
23 3 4 13 1 10 9 7 13 0 1 13 2 13 2 10 9 16 3 13 1 10 9 2
43 1 10 9 10 9 1 0 9 15 4 13 1 13 9 1 10 9 1 9 1 11 2 1 10 0 9 1 9 1 10 9 2 9 7 10 9 0 1 9 1 9 0 2
22 1 10 9 1 12 13 10 9 1 12 9 7 10 9 0 1 12 9 1 9 5 2
14 3 13 10 9 1 10 9 11 11 11 2 8 2 2
28 10 9 1 9 12 1 11 4 13 3 10 9 7 13 9 0 1 10 9 2 16 13 1 9 0 1 3 2
135 1 10 9 2 11 11 13 16 13 10 9 16 1 10 9 3 0 1 9 1 9 1 9 16 3 13 15 13 2 9 1 11 11 13 9 1 10 9 1 9 0 1 9 1 9 1 9 1 9 1 10 9 0 7 13 16 13 0 16 10 10 9 16 1 11 11 1 11 4 13 9 1 13 1 9 1 9 13 1 10 9 1 10 9 16 13 15 1 10 9 3 13 0 16 16 15 3 4 13 2 15 15 13 10 9 1 13 15 0 9 2 15 1 15 1 10 9 1 10 9 0 2 1 9 3 0 7 1 9 1 10 9 1 15 2
13 1 10 9 2 13 1 10 9 4 13 1 15 2
13 3 7 9 16 10 9 13 15 9 16 13 3 2
20 3 0 2 1 10 9 1 10 9 2 10 4 7 13 3 1 9 3 0 2
7 15 15 13 1 9 0 2
18 10 9 13 1 10 9 13 10 9 3 0 1 10 11 1 10 9 2
29 10 0 9 13 10 9 2 1 11 2 1 10 0 9 1 10 11 11 12 2 1 10 9 1 10 11 11 12 2
18 13 15 1 10 9 16 13 10 9 1 11 11 1 9 0 1 11 2
16 11 13 1 9 1 10 9 1 9 11 11 11 2 12 2 2
11 11 4 3 13 1 10 9 13 16 13 2
42 10 11 7 11 11 1 11 2 1 9 2 11 11 11 7 11 1 11 2 2 13 10 9 2 9 7 13 0 1 10 9 1 9 0 1 12 9 2 12 5 2 2
20 1 10 9 13 10 9 0 1 9 2 13 1 10 9 8 8 7 13 11 2
17 3 1 10 12 5 1 10 9 13 1 3 1 10 9 1 9 2
12 3 13 10 0 9 15 13 10 9 13 9 2
27 1 11 1 12 10 11 13 1 10 9 1 12 9 2 15 16 15 13 1 10 9 3 0 1 10 9 2
14 9 1 10 9 16 13 10 9 1 10 9 1 9 2
31 1 9 0 2 10 9 1 2 11 10 11 11 2 1 11 13 3 0 2 13 2 11 10 11 11 1 11 11 2 2 2
23 11 11 11 2 13 1 11 1 11 2 3 10 9 2 11 11 2 13 10 9 1 9 2
25 1 10 9 7 1 9 1 9 2 10 11 4 13 13 10 9 1 10 9 0 1 10 9 0 2
7 9 0 1 9 1 10 9
36 10 9 12 2 1 9 1 10 9 1 10 9 2 15 13 10 0 9 1 9 1 10 9 11 11 11 7 9 1 10 9 11 11 11 11 2
12 10 9 13 9 0 1 10 9 7 10 9 2
28 1 10 12 1 11 1 10 12 2 10 9 4 13 1 11 2 15 16 13 0 9 1 10 9 1 10 9 2
29 3 1 10 9 1 11 2 11 15 13 1 16 10 9 1 9 4 13 15 16 13 10 9 0 1 10 9 0 2
53 13 10 9 0 0 1 10 9 16 15 13 1 9 2 1 9 10 9 1 10 9 7 10 9 13 1 10 9 11 11 10 9 3 1 10 9 2 13 10 11 7 10 11 2 2 10 9 7 10 9 2 2 2
15 15 16 4 7 13 13 13 1 10 9 7 3 13 15 2
16 13 1 12 7 12 2 3 1 11 12 7 3 1 11 11 2
45 10 9 4 13 1 0 9 7 9 7 15 1 9 0 0 2 13 1 9 16 10 9 13 3 9 0 2 10 0 9 2 10 0 9 1 10 9 7 10 9 1 9 3 0 2
20 10 9 0 1 11 1 10 9 1 10 9 1 10 9 13 1 2 11 2 2
55 3 10 9 13 10 9 1 9 0 2 15 13 1 10 9 1 10 9 1 9 0 2 13 1 9 2 15 13 10 9 0 7 3 0 1 15 16 13 10 9 1 10 9 2 13 1 9 1 10 9 2 7 12 9 2
21 1 12 7 12 13 12 1 10 9 1 10 9 9 1 10 9 1 10 11 11 2
