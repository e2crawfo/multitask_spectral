504 11
19 9 13 1 10 9 2 15 13 1 10 3 0 9 2 3 0 9 13 2
8 2 15 4 13 10 9 2 2
33 15 1 10 0 9 1 9 1 9 13 1 10 0 9 1 10 9 2 16 9 13 4 10 9 2 15 13 9 7 3 0 9 2
24 2 9 1 10 9 4 3 0 2 14 13 9 1 15 15 0 13 7 13 15 7 9 2 2
12 1 10 0 9 13 9 3 1 9 0 9 2
28 1 14 13 10 0 9 1 9 7 9 4 15 13 3 9 1 9 2 3 9 3 4 4 13 10 0 9 2
46 3 9 13 10 9 7 9 4 1 9 13 10 0 9 1 9 7 9 2 2 2 9 4 3 3 10 9 1 10 9 2 7 3 1 9 1 9 4 15 13 10 9 7 9 2 2
30 15 13 3 10 9 3 9 2 3 9 2 3 1 14 13 9 9 7 9 4 13 7 13 15 1 10 9 1 9 2
20 10 0 9 13 3 14 13 9 1 10 9 7 13 9 13 9 1 9 9 2
28 3 3 15 3 4 13 10 0 9 1 9 7 9 2 4 15 13 9 1 10 3 0 9 7 9 1 9 2
15 15 13 16 3 9 3 4 4 10 3 0 14 13 9 2
46 1 10 0 9 4 9 3 0 1 0 9 7 9 1 9 9 7 2 3 0 13 2 15 4 13 0 10 9 1 7 0 16 9 4 13 15 7 13 7 13 9 1 10 0 9 2
34 3 9 4 13 1 10 15 2 7 1 15 13 15 3 10 9 2 16 15 3 13 0 9 15 13 7 13 9 1 15 1 0 9 2
38 1 0 9 4 15 13 10 9 7 9 1 9 14 3 13 3 12 7 0 9 15 3 13 3 3 1 15 2 9 2 9 7 10 0 9 1 9 2
20 3 15 13 9 9 7 9 4 15 13 3 3 9 7 3 9 10 0 9 2
10 10 9 1 9 4 0 9 1 9 2
24 7 10 0 13 3 3 13 15 2 1 3 0 7 0 9 16 15 3 13 1 9 0 9 2
23 3 3 9 13 1 9 3 1 9 4 15 4 3 13 2 9 7 9 13 3 10 9 2
27 7 1 14 4 13 1 9 4 15 13 1 9 14 13 7 13 9 2 15 13 1 9 10 9 1 9 2
64 2 15 4 13 15 0 9 2 15 4 13 15 1 10 0 9 7 1 9 14 13 9 2 15 4 13 15 1 9 14 2 13 2 10 9 2 14 13 15 7 10 9 7 15 15 13 2 15 4 13 15 10 0 9 2 15 13 9 15 13 10 9 2 2
9 9 14 13 9 2 9 13 0 2
25 10 9 13 15 2 1 9 9 2 3 9 13 13 7 13 9 3 16 15 13 15 15 13 15 2
24 10 9 1 10 0 9 4 9 2 0 9 2 2 15 15 4 13 1 14 13 9 1 9 2
19 14 4 9 1 9 4 3 10 0 7 0 9 2 1 0 9 1 9 2
17 7 3 9 4 13 10 9 2 0 9 13 4 0 3 1 9 2
22 10 0 9 1 9 9 7 9 1 9 13 15 3 3 3 15 13 9 1 0 9 2
30 9 4 13 1 9 7 9 1 9 9 2 9 1 9 13 3 14 13 7 15 13 3 3 9 15 13 15 1 15 2
34 15 13 7 16 9 3 13 10 3 0 9 1 9 1 10 3 0 7 9 1 10 3 0 9 2 15 3 3 4 13 1 0 9 2
18 10 0 9 15 4 13 9 4 3 3 3 0 10 0 1 10 9 2
8 7 1 9 9 13 15 3 2
36 3 4 3 9 1 10 9 4 3 3 13 7 0 2 3 0 7 0 3 3 15 13 3 3 0 9 7 9 1 14 13 15 10 0 9 2
24 9 4 1 0 9 0 9 2 7 15 4 3 0 16 9 13 9 9 2 10 9 14 13 2
9 15 4 13 15 3 10 9 13 2
9 15 13 10 0 9 1 9 9 2
13 13 15 15 1 15 7 1 3 9 1 10 9 2
21 1 10 0 9 13 15 9 1 14 4 0 2 0 2 0 7 0 1 10 9 2
18 15 4 3 13 3 0 2 3 0 7 3 1 9 3 0 7 0 2
19 7 1 10 0 9 13 15 3 3 10 0 9 7 13 3 9 1 9 2
41 1 14 1 10 9 4 13 15 1 9 1 9 4 15 13 15 3 1 10 0 9 7 3 13 15 1 9 2 15 13 3 1 10 0 9 0 1 9 1 9 2
35 0 9 4 13 15 2 3 9 7 9 2 15 1 9 13 10 0 9 1 14 13 9 1 9 1 9 7 1 14 13 9 1 0 9 2
25 15 15 13 9 3 0 1 9 1 10 3 9 4 9 1 10 3 9 2 15 4 13 7 9 2
20 10 9 4 3 10 9 2 15 1 15 13 9 1 3 1 9 14 13 9 2
30 1 9 13 9 3 1 9 7 13 1 15 1 0 9 2 7 1 0 4 10 0 2 0 2 7 0 9 0 9 2
32 10 0 9 15 13 1 9 7 9 4 4 13 1 9 1 9 2 0 16 10 9 15 13 4 3 0 7 0 1 0 9 2
36 9 1 10 9 1 9 15 13 7 10 9 15 13 3 2 13 1 10 0 9 11 11 11 2 15 1 0 9 13 9 7 9 1 0 9 2
15 10 0 9 13 9 1 9 1 10 0 9 1 9 9 2
40 15 4 3 13 10 0 9 15 4 13 1 9 9 14 13 1 10 0 2 0 9 1 9 7 14 13 1 0 9 1 10 0 9 2 15 4 15 9 13 2
27 1 14 13 9 1 10 9 13 11 10 9 9 1 9 1 10 9 0 9 2 1 9 1 9 1 9 2
35 1 9 1 0 0 9 4 15 13 16 9 13 3 1 1 0 9 7 7 1 9 2 9 1 9 7 9 7 1 2 0 2 9 2 12
29 12 1 10 0 9 1 9 7 9 2 13 11 11 11 2 9 7 9 1 9 1 2 0 2 9 1 10 11 2
12 0 1 0 9 1 9 2 12 2 12 12 2
19 1 10 9 4 9 3 0 2 7 3 1 10 0 9 4 9 3 0 2
6 15 13 9 3 3 2
36 2 15 13 7 16 9 1 10 9 0 9 15 15 13 1 0 9 13 14 4 10 9 1 9 7 13 10 9 2 3 15 15 13 0 9 2
34 9 13 4 3 0 7 0 7 9 2 3 1 9 1 16 15 4 3 13 1 16 9 9 4 13 3 1 0 0 0 9 2 2 12
12 12 1 11 11 11 2 9 2 9 1 9 2
10 0 1 11 12 2 9 12 2 12 2
9 13 10 9 1 9 1 0 9 2
8 4 9 9 13 10 0 9 2
26 1 14 13 10 9 13 11 1 0 9 10 9 0 9 1 0 9 7 13 7 9 10 3 0 9 2
18 9 13 1 10 9 10 3 0 9 7 1 0 9 7 1 0 9 2
31 2 15 13 1 9 1 12 7 12 9 9 2 15 13 15 14 13 1 0 9 7 3 7 13 1 10 9 15 13 2 2
15 11 9 4 3 13 15 15 13 1 9 7 3 9 13 2
26 1 15 4 15 7 4 13 10 9 1 10 9 1 9 7 0 9 1 10 9 1 12 7 12 9 2
24 9 3 0 9 13 15 3 4 13 3 1 16 15 13 0 9 1 0 9 7 0 0 9 2
42 11 13 3 3 10 9 9 2 15 1 15 13 9 9 1 9 2 9 9 1 10 0 9 2 0 9 7 9 1 9 7 9 2 0 9 7 9 1 9 7 9 2
18 9 13 3 10 9 1 10 9 2 15 4 0 7 3 3 3 0 2
21 10 9 15 13 1 4 3 0 1 9 7 10 0 9 15 13 4 3 3 0 2
20 7 1 14 13 7 13 10 1 10 0 9 7 9 4 10 9 1 9 0 2
42 11 2 7 0 9 1 15 2 13 16 9 13 9 1 16 9 3 13 9 1 10 0 9 2 16 15 3 13 0 2 0 7 3 3 0 1 9 1 10 0 9 2
18 9 1 3 2 0 2 9 4 4 3 13 3 7 1 10 0 9 2
31 7 1 14 13 10 0 9 1 0 9 1 9 7 3 1 9 9 1 9 2 3 4 9 9 3 0 14 13 9 1 2
12 3 1 10 9 13 9 3 3 7 1 9 2
12 15 13 3 1 10 0 9 1 10 0 9 2
28 9 13 3 10 0 9 14 13 16 15 13 10 9 7 10 9 1 9 15 10 0 9 7 0 0 9 13 2
4 3 4 9 2
10 13 9 1 9 3 1 9 7 9 2
10 13 10 9 14 13 1 10 0 9 2
13 10 9 13 9 1 9 2 0 9 2 1 9 2
5 0 7 3 0 2
7 15 13 9 14 4 0 2
22 0 9 13 16 10 0 9 13 3 1 10 9 15 3 13 1 9 0 9 1 9 2
38 10 0 9 1 11 2 3 15 3 7 3 13 9 1 10 9 2 13 3 9 1 16 9 4 1 9 14 13 10 0 9 1 9 1 7 1 9 2
44 3 0 4 3 16 3 10 0 0 9 2 7 15 1 10 9 7 1 0 0 9 2 13 15 2 0 2 14 13 9 1 10 0 1 9 1 14 13 9 7 9 1 9 2
30 1 9 9 4 13 16 9 1 0 9 13 3 3 1 9 9 2 3 16 15 13 1 9 1 15 9 13 10 9 2
21 15 13 3 3 10 9 16 9 13 9 1 0 7 0 9 1 7 9 7 9 2
8 15 13 3 1 12 9 9 2
14 3 13 9 0 1 12 9 9 1 10 9 7 9 2
26 7 10 0 9 13 2 3 7 15 1 10 0 9 2 3 0 3 1 16 9 13 0 3 1 9 2
20 3 0 9 7 9 4 3 13 9 16 15 3 4 13 1 0 3 1 9 2
25 10 0 9 4 3 1 9 10 9 1 9 9 1 10 9 1 3 10 0 9 0 9 1 9 2
14 9 12 2 7 3 3 2 13 10 0 9 0 9 2
8 3 4 15 13 1 9 9 2
44 15 13 0 14 13 15 1 9 16 4 3 0 10 0 9 13 1 0 9 7 0 9 3 13 1 0 9 9 4 3 9 3 3 13 0 9 7 0 9 3 15 3 13 2
15 15 4 3 13 3 3 15 13 9 0 0 7 0 9 2
11 0 7 3 3 1 0 4 10 0 9 2
34 16 15 13 1 9 9 7 9 1 9 1 9 1 10 0 9 4 10 0 9 3 13 3 7 3 13 16 9 13 0 7 0 9 2
22 1 9 0 9 13 3 12 0 9 2 3 12 9 2 7 12 9 2 3 12 9 2
13 9 0 9 1 0 9 4 3 0 2 3 0 2
21 9 13 3 3 14 13 16 15 13 10 0 9 10 9 1 9 7 1 9 13 2
29 15 3 3 4 13 16 15 13 10 0 0 9 3 12 7 16 15 3 3 3 13 12 2 13 12 9 1 9 2
18 9 9 1 9 4 3 1 10 9 3 3 0 7 1 10 0 9 2
25 3 3 1 10 7 10 9 13 9 0 2 0 9 1 10 0 9 2 0 7 0 9 7 9 2
18 3 3 1 9 1 0 9 1 10 9 4 9 3 13 9 1 9 2
7 7 15 3 13 1 9 2
25 9 12 4 1 9 13 9 7 15 13 3 1 10 9 16 0 0 9 13 3 1 9 1 9 2
22 1 0 9 13 3 0 9 15 13 9 7 9 9 1 9 15 13 0 3 0 9 2
19 0 4 16 15 1 0 0 9 3 3 13 10 9 0 0 7 0 9 2
25 15 4 3 3 13 16 1 0 9 1 9 7 9 9 13 3 10 3 0 7 3 3 0 9 2
23 15 4 3 13 10 9 3 9 7 9 13 15 3 3 1 9 1 9 2 9 7 9 2
17 3 13 10 0 9 9 1 10 3 0 7 1 10 3 0 9 2
14 9 13 3 13 10 0 9 7 10 0 7 0 9 2
13 3 0 1 0 9 4 10 9 15 9 3 13 2
19 3 0 13 9 7 9 16 7 9 7 9 4 13 10 9 1 0 9 2
8 15 13 3 1 9 1 9 2
18 9 12 13 3 12 9 1 10 0 9 9 1 12 9 1 10 0 2
16 9 12 13 15 16 9 1 10 9 7 9 4 14 13 9 2
24 7 3 3 13 9 1 3 0 9 7 9 9 15 13 3 1 10 3 0 7 3 0 9 2
12 3 1 9 1 0 0 0 9 13 9 3 2
14 3 3 3 0 4 9 1 9 3 1 10 0 9 2
8 9 13 9 1 10 0 9 2
15 1 15 13 3 3 10 3 0 9 4 10 3 0 9 2
6 9 13 9 7 9 2
23 0 9 13 1 10 9 10 0 9 3 16 0 9 1 9 1 10 9 7 9 13 3 2
8 9 13 15 1 3 0 9 2
44 15 13 9 2 9 2 9 2 9 7 9 7 9 1 10 9 2 3 1 9 1 10 3 3 0 9 2 3 1 9 1 9 7 1 9 3 9 3 0 3 13 7 9 2
13 10 0 9 1 9 9 1 9 7 9 13 0 2
28 9 0 9 1 9 4 3 3 0 16 15 15 13 3 4 10 0 9 7 10 0 9 1 9 10 9 13 2
29 15 4 3 13 3 16 0 7 3 0 9 9 7 9 13 15 1 9 1 0 9 1 9 7 3 13 3 13 2
25 1 10 10 0 9 13 10 0 9 1 9 9 7 10 0 9 13 3 1 9 0 2 0 9 2
7 3 13 15 1 10 9 2
10 12 9 4 13 15 13 7 3 13 2
8 10 0 9 7 9 7 9 2
12 0 9 7 9 1 9 1 9 7 1 9 2
111 10 0 9 16 9 13 9 7 16 9 1 10 0 9 4 3 0 1 9 2 7 0 9 2 13 10 9 1 0 9 3 3 3 16 9 13 9 7 3 2 1 10 9 16 1 10 0 9 13 15 9 1 10 9 1 3 12 2 12 9 1 10 9 1 12 2 12 9 2 3 16 9 1 3 0 9 4 3 0 1 9 7 9 2 1 10 9 16 9 1 3 0 0 9 3 7 3 2 3 1 0 9 2 13 10 0 1 9 0 9 2
27 15 15 13 1 9 3 1 10 15 15 13 13 10 9 1 9 4 10 0 9 1 10 0 9 1 9 2
33 15 13 3 3 3 1 10 9 1 10 0 9 2 3 9 13 14 13 10 0 9 7 3 15 7 9 13 0 7 0 0 9 2
32 3 3 13 15 3 3 3 10 9 15 13 0 9 0 7 3 0 7 15 15 3 13 1 0 9 7 1 9 9 13 9 2
15 1 3 0 9 13 9 4 3 0 7 9 3 3 3 2
25 9 13 3 3 3 2 3 15 4 10 7 0 7 0 9 2 16 9 4 13 15 7 3 3 2
14 15 13 3 16 10 9 4 13 15 3 3 1 9 2
14 9 13 3 1 0 9 3 1 9 1 10 0 9 2
18 15 15 4 13 4 10 3 0 9 1 9 9 2 9 1 9 9 2
11 10 9 1 9 4 0 1 9 0 9 2
11 15 4 3 13 10 3 0 9 1 9 2
37 15 4 10 9 15 3 3 13 12 7 12 9 7 9 1 3 0 0 9 2 3 9 7 3 9 9 1 0 9 4 13 1 0 9 7 9 2
19 3 1 10 9 1 9 7 9 4 9 3 7 3 4 3 13 1 9 2
25 1 0 0 9 1 10 0 9 13 15 3 1 9 3 1 9 1 9 2 9 7 9 1 9 2
5 10 9 4 13 2
9 7 15 4 0 9 16 3 13 2
20 0 1 15 3 4 16 9 13 0 1 9 1 9 1 9 1 9 1 9 2
7 3 4 15 3 10 9 2
34 3 9 0 1 10 3 0 9 4 13 16 15 4 13 9 7 3 4 10 3 3 0 9 1 16 9 4 4 13 9 7 9 13 2
31 15 4 3 13 16 2 3 3 10 0 2 3 0 9 13 15 4 13 9 9 2 9 1 9 7 9 3 13 3 0 2
16 15 13 3 9 9 14 13 1 16 9 13 3 0 7 0 2
15 1 9 13 1 10 9 0 7 0 9 15 13 9 9 2
13 9 0 9 14 13 15 1 0 9 4 10 9 2
17 1 9 13 9 14 13 9 14 13 15 1 10 3 3 0 9 2
33 0 9 13 7 15 4 14 13 1 9 3 9 13 7 9 3 3 13 9 1 10 0 7 0 9 3 3 15 13 3 1 9 2
14 1 7 1 16 9 13 3 0 9 13 15 0 9 2
16 3 13 9 1 3 0 9 15 15 3 4 13 9 1 9 2
11 0 9 4 14 13 9 0 1 0 9 2
15 10 0 13 1 9 14 13 0 7 3 0 3 7 3 2
23 15 13 7 16 9 3 3 13 13 16 3 3 4 13 1 14 13 9 0 9 7 9 2
47 16 9 13 7 3 0 9 16 9 4 13 9 14 3 7 0 13 9 7 10 9 7 10 9 1 10 9 7 10 0 2 13 3 7 0 9 7 9 1 0 3 7 15 15 4 3 2
9 7 15 13 10 0 9 14 13 2
21 9 4 13 9 14 3 3 13 7 10 9 2 3 7 10 9 0 9 1 9 2
19 15 13 1 9 9 3 0 9 1 16 9 9 7 9 1 9 4 13 2
16 15 13 10 0 9 15 13 9 1 0 9 7 3 9 9 2
39 9 4 1 0 9 10 9 1 9 9 2 9 9 14 0 13 1 10 9 7 9 2 9 7 0 2 7 10 9 13 3 7 15 1 15 1 0 9 2
10 9 9 4 13 1 9 1 9 9 2
27 10 0 9 15 1 9 13 15 13 3 0 9 14 13 9 7 9 1 10 3 0 9 0 7 0 9 2
16 9 1 9 9 13 10 0 9 1 9 9 2 9 7 9 2
18 4 15 3 2 13 15 2 4 9 9 14 13 1 2 9 9 2 2
38 7 3 10 9 15 15 0 1 9 4 13 15 2 16 15 13 3 1 0 9 7 9 7 1 9 1 10 0 2 3 0 7 3 0 7 0 9 2
11 6 2 9 4 13 3 15 7 10 9 2
52 9 13 3 16 9 4 13 10 9 1 0 9 7 9 2 16 15 4 13 0 9 1 9 7 9 2 16 15 4 13 9 14 7 13 10 9 7 13 9 7 9 2 16 15 4 4 10 0 7 0 9 2
22 7 15 13 3 1 14 13 9 0 1 10 9 7 14 13 13 0 9 1 0 9 2
20 10 0 9 4 16 9 13 3 1 1 9 7 16 15 13 9 1 0 9 2
21 15 1 13 10 0 9 2 3 7 3 3 2 10 9 0 9 1 10 0 9 2
105 15 13 1 10 9 15 15 15 13 9 1 3 1 15 2 9 15 13 0 7 0 9 1 9 1 9 2 1 16 15 4 13 15 2 2 9 15 13 10 0 9 1 14 13 9 2 15 4 13 15 3 2 2 9 15 13 3 10 0 9 1 14 1 9 13 10 9 2 15 4 3 3 0 2 2 9 15 13 9 2 1 14 13 3 3 0 2 2 9 15 13 15 7 13 9 2 1 14 4 13 9 7 9 2 2
24 15 13 3 2 16 10 15 4 1 9 1 10 0 9 2 16 0 9 3 13 1 0 9 2
17 3 13 15 1 2 16 0 9 1 9 3 4 3 9 7 9 2
47 3 1 10 9 3 15 13 16 9 4 4 0 2 3 1 9 7 9 1 0 2 0 9 2 13 15 9 1 9 1 10 9 7 9 16 9 1 9 7 9 1 3 13 7 9 9 2
13 10 0 9 7 9 14 13 9 13 3 10 9 2
20 7 16 15 1 9 13 1 9 7 4 13 3 9 3 13 15 10 0 9 2
13 1 12 9 3 13 10 9 1 10 0 0 9 2
7 9 4 9 9 1 9 2
29 10 0 9 13 3 16 9 9 13 1 9 2 7 3 12 0 1 9 13 13 10 0 9 2 1 9 0 9 2
28 3 15 3 13 10 9 1 9 9 13 10 9 16 15 1 15 4 13 14 13 0 2 1 9 1 9 9 2
9 3 10 9 1 0 9 2 3 2
31 7 15 4 0 7 0 14 13 10 9 15 2 1 14 13 10 9 0 2 9 0 7 9 0 2 13 0 9 7 9 2
26 9 13 15 3 3 1 16 9 3 4 10 0 9 9 2 10 0 9 2 6 2 0 9 13 3 2
16 15 13 3 3 15 3 0 13 13 1 10 10 0 1 9 2
6 13 15 15 3 0 2
30 6 2 1 15 13 9 1 10 0 0 9 2 15 4 13 1 9 2 13 2 13 9 2 13 9 2 13 9 9 2
9 10 9 1 9 4 13 7 13 2
8 15 13 3 15 4 13 15 2
12 15 4 13 13 9 9 1 10 9 1 9 2
39 15 4 13 1 10 9 1 9 1 9 1 9 1 0 7 0 9 7 1 10 9 1 9 1 9 1 9 1 9 7 9 2 1 9 1 9 7 9 2
41 10 0 9 15 0 9 13 1 9 1 14 3 13 15 1 2 10 0 9 2 2 2 2 4 3 3 0 7 10 0 9 2 1 15 9 1 9 4 3 0 2
28 15 4 3 3 13 2 16 9 7 9 2 9 1 10 0 0 9 3 2 4 3 0 9 7 3 3 0 2
45 15 4 0 7 0 2 14 3 0 0 9 13 2 13 9 0 9 7 9 1 9 7 9 2 13 10 0 9 7 9 2 1 14 13 10 9 9 14 1 9 13 10 0 9 2
17 15 13 1 9 9 15 13 2 16 15 4 13 3 3 3 3 2
18 3 0 9 13 13 1 10 9 7 9 15 13 9 1 9 7 9 2
4 9 4 13 2
20 7 15 13 16 15 13 1 9 1 10 0 2 0 2 3 3 13 0 9 2
17 15 13 3 1 16 9 9 13 1 9 14 13 10 9 7 9 2
16 15 13 10 9 3 3 16 15 3 4 13 14 13 10 9 2
16 16 9 4 13 10 9 7 9 2 13 15 3 15 15 13 2
28 7 15 4 13 16 15 3 13 9 2 15 4 0 1 10 0 9 2 7 15 15 7 9 4 3 0 1 2
10 15 13 9 2 15 13 9 1 9 2
3 3 9 2
8 10 0 9 0 1 0 9 2
17 15 4 1 0 9 13 16 15 3 13 0 9 1 9 7 9 2
23 11 11 2 9 1 9 7 9 2 13 16 1 10 0 9 4 9 0 7 0 1 9 2
18 15 13 3 16 9 13 2 16 10 9 13 1 0 9 14 13 9 2
20 3 0 9 13 2 13 15 1 9 7 9 2 15 13 15 9 1 3 9 2
11 10 0 9 13 1 3 0 7 0 9 2
30 3 7 3 1 11 2 3 9 1 10 0 12 9 13 7 13 1 10 9 7 9 2 13 9 3 0 7 0 9 2
20 15 4 3 10 9 16 12 9 1 9 2 9 7 9 1 11 13 1 9 2
30 3 4 10 0 9 1 0 9 13 7 10 3 0 2 7 15 15 13 15 1 0 2 0 2 9 1 9 7 9 2
45 4 3 9 14 13 1 9 13 7 10 3 0 0 9 2 15 9 4 13 9 1 2 3 15 1 10 0 9 1 10 9 13 0 9 7 4 13 3 0 9 1 10 0 9 2
21 4 15 0 2 16 9 1 14 13 10 9 4 13 15 1 9 7 13 10 9 2
17 4 15 3 1 10 9 13 1 14 13 10 9 9 1 10 0 2
12 3 13 15 3 1 9 1 14 3 13 15 2
20 4 3 9 1 9 9 1 9 1 9 9 13 10 9 2 15 13 1 9 2
52 15 4 3 3 13 10 0 7 0 1 9 1 10 0 9 2 16 9 13 10 9 14 13 3 1 2 10 2 9 2 14 4 13 1 1 10 10 3 0 1 9 2 14 13 2 13 7 13 10 0 9 2
10 10 9 4 15 9 13 1 0 9 2
29 4 15 3 13 15 1 15 1 10 3 0 9 9 7 14 13 16 15 3 4 3 0 7 9 3 15 13 9 2
9 4 15 3 13 9 1 9 3 2
15 1 9 1 14 3 13 9 9 7 9 4 15 13 9 2
21 15 4 13 16 10 0 9 13 3 3 7 10 0 9 7 3 7 13 1 11 2
15 3 3 9 3 1 4 13 1 7 13 1 9 7 9 2
4 15 4 0 2
11 15 15 13 15 4 3 3 0 7 9 2
20 7 15 9 4 3 1 10 9 4 13 1 15 10 9 14 13 1 0 9 2
15 15 13 3 0 9 2 13 15 0 3 1 3 0 9 2
18 10 0 9 1 10 9 13 3 3 1 9 1 10 0 9 1 9 2
7 7 4 15 3 13 0 2
39 10 9 2 15 4 10 0 7 3 10 3 0 2 0 1 9 7 1 10 0 7 9 2 10 9 1 9 3 9 9 13 2 10 9 4 13 3 3 2
16 15 13 10 9 1 9 10 0 9 2 10 9 9 9 3 2
6 3 13 15 1 15 2
13 4 15 13 10 0 9 7 4 15 0 0 9 2
13 3 9 13 13 1 0 9 1 9 1 0 9 2
13 13 15 9 14 13 1 10 9 3 1 10 9 2
6 4 15 13 1 15 2
13 3 13 15 9 14 13 10 9 15 13 3 1 2
23 10 9 2 15 3 13 3 1 10 3 0 2 1 9 1 15 14 13 1 3 0 9 2
13 3 13 15 9 14 13 10 9 1 10 3 9 2
20 7 3 4 15 13 10 0 2 0 7 0 9 1 15 15 4 0 1 9 2
14 9 15 13 10 9 4 3 13 3 1 10 0 9 2
24 15 13 3 3 15 14 13 2 7 15 4 13 15 1 9 2 1 9 1 10 9 15 13 2
23 9 9 14 13 1 7 4 13 7 10 0 7 0 9 1 9 1 10 0 9 7 9 2
12 15 13 3 0 9 2 15 4 13 0 9 2
9 15 4 13 3 16 9 4 0 2
6 15 4 15 1 9 2
9 3 13 15 15 15 4 3 0 2
4 15 13 9 2
7 10 15 13 15 1 15 2
8 13 1 16 15 4 3 13 2
9 3 13 9 15 14 13 15 1 2
6 9 13 3 1 9 2
13 3 15 4 9 13 15 15 0 3 15 13 15 2
12 3 3 9 13 9 1 9 4 15 3 13 2
15 7 3 13 15 14 13 9 1 12 0 9 7 12 9 2
11 7 12 9 13 10 9 1 10 0 9 2
21 15 13 9 15 13 3 1 0 9 4 4 3 0 14 13 3 7 15 15 13 2
5 13 9 2 9 2
7 13 1 15 1 0 9 2
13 15 13 10 9 2 10 9 2 6 2 0 9 2
22 14 3 0 13 9 9 7 0 9 1 9 13 1 10 0 9 1 9 15 4 0 2
10 0 9 7 10 4 13 3 1 9 2
10 15 4 3 3 0 16 15 13 15 2
21 15 13 14 13 1 10 9 1 9 7 13 16 7 9 4 15 3 13 9 3 2
16 15 13 16 15 4 13 9 3 15 4 13 15 9 0 9 2
12 15 13 9 1 9 7 3 13 15 10 9 2
33 0 9 13 3 1 9 1 9 0 9 1 0 9 2 3 0 9 2 9 2 9 2 0 9 7 7 9 1 14 13 10 9 2
30 9 15 3 13 9 1 9 2 9 3 10 0 2 0 9 3 4 13 1 10 9 1 9 2 3 0 15 3 4 2
8 7 15 3 13 1 15 0 2
13 15 4 3 13 13 15 1 9 1 9 7 15 2
15 7 16 15 13 12 9 1 9 3 15 4 13 4 0 2
27 13 3 9 1 0 9 9 1 9 1 10 10 9 2 15 4 13 1 7 13 2 4 10 15 3 13 2
31 13 10 9 13 9 1 9 1 9 1 0 9 2 0 9 2 0 9 15 4 13 1 10 3 7 3 0 9 1 9 2
15 11 13 3 12 9 10 0 9 3 9 7 9 4 0 2
9 15 13 15 1 9 3 2 3 2
6 15 4 13 1 9 2
15 0 4 15 0 1 10 9 7 13 9 1 9 1 9 2
19 3 4 15 13 1 10 9 7 15 4 13 9 1 10 3 3 0 9 2
18 0 13 15 3 10 9 1 14 13 3 1 9 3 3 9 4 0 2
19 15 13 3 3 10 0 9 9 2 0 3 2 7 15 15 13 7 0 2
24 15 4 0 14 4 9 3 9 13 3 3 16 15 13 1 9 7 9 2 3 4 15 15 2
9 7 10 9 4 15 3 9 1 2
14 7 9 13 3 0 1 9 3 1 14 13 13 1 2
17 2 15 13 3 9 14 13 15 3 15 13 15 2 2 13 15 2
12 3 15 13 1 9 13 15 10 3 0 9 2
28 10 0 9 13 0 9 1 16 15 13 0 2 0 0 9 1 9 1 9 7 1 15 15 4 0 7 0 2
19 7 10 0 9 1 9 4 3 13 9 9 7 10 0 7 3 0 9 2
7 9 4 13 3 1 9 2
6 10 0 9 13 3 2
29 3 9 13 2 13 15 3 16 15 3 4 13 9 10 9 2 7 1 9 4 15 13 10 0 9 14 13 9 2
6 7 15 13 3 3 2
46 4 13 15 4 0 2 0 7 0 2 3 13 9 7 0 2 13 10 0 2 3 16 10 9 13 9 1 9 1 9 7 9 1 0 9 9 1 10 0 9 2 3 0 1 15 2
26 15 4 4 10 0 9 1 10 0 9 2 2 4 10 1 11 0 9 3 3 0 4 13 10 9 2
7 15 13 3 0 1 9 2
9 15 13 2 15 10 4 10 2 2
14 7 3 15 13 3 1 9 13 15 3 10 9 3 2
19 3 13 15 2 3 6 3 4 10 10 10 2 3 15 0 13 15 3 2
5 15 4 3 0 2
11 7 15 4 13 1 16 9 4 13 3 2
10 3 4 15 13 9 13 16 15 13 2
11 15 4 3 0 16 15 4 13 0 9 2
12 10 0 9 13 9 3 1 16 15 13 9 2
9 1 9 9 13 15 12 9 1 2
8 9 4 3 3 3 0 3 2
14 15 13 1 10 9 7 3 3 13 15 1 9 9 2
12 15 4 9 1 0 9 14 13 1 10 9 2
18 6 2 10 9 2 15 3 4 0 1 9 2 4 14 13 3 3 2
38 1 9 4 15 14 13 3 0 9 1 9 7 15 4 13 3 0 9 7 15 3 3 4 0 7 10 9 1 3 0 9 4 3 3 0 14 13 2
7 9 13 9 1 0 9 2
8 1 10 0 9 7 0 9 2
6 1 9 13 15 9 2
16 15 4 9 15 3 4 0 1 9 7 13 15 7 15 13 2
4 15 4 0 2
4 3 1 9 2
9 15 4 0 1 14 4 13 3 2
8 0 1 14 4 13 10 9 2
8 15 13 3 3 0 15 4 2
16 15 13 3 3 0 10 3 9 4 7 3 3 15 13 13 2
40 9 4 0 1 0 9 9 2 9 1 9 2 2 0 9 2 0 9 2 7 11 11 2 9 7 9 2 11 2 11 2 12 2 0 9 2 0 9 2 2
10 10 0 13 0 9 14 13 9 0 2
13 15 1 15 4 14 13 9 3 2 4 0 9 2
15 3 15 13 9 13 15 13 10 0 9 1 9 2 9 2
15 7 16 15 3 3 2 3 3 3 2 13 15 1 9 2
31 1 0 9 9 13 15 10 0 9 3 3 2 1 14 1 10 0 9 2 9 1 2 13 3 10 0 9 1 11 9 2
16 7 13 15 10 9 1 11 11 9 1 9 1 11 13 9 2
8 15 13 3 1 9 2 9 2
5 15 13 1 9 2
5 15 13 1 9 2
11 1 10 0 9 13 0 9 1 0 9 2
17 9 15 13 1 2 7 13 2 10 9 10 0 9 1 9 13 2
25 3 16 15 13 9 14 13 3 1 14 13 3 7 13 3 2 3 1 14 13 9 7 13 9 2
17 1 10 0 9 13 9 10 9 4 0 7 10 0 9 1 9 2
9 10 9 4 10 0 9 3 13 2
30 15 13 13 10 0 10 9 1 10 9 2 3 9 1 0 9 7 9 13 3 2 3 1 9 1 10 0 9 9 2
5 15 13 1 9 2
8 10 0 9 13 3 10 9 2
38 15 2 13 9 2 2 13 1 10 0 9 2 13 1 10 0 2 0 9 2 15 3 13 1 14 13 9 0 7 0 9 1 10 9 7 9 9 2
36 16 9 13 3 1 10 9 3 16 15 3 13 13 3 7 3 1 14 13 10 0 9 2 7 1 9 10 0 9 15 4 9 1 10 9 2
5 15 13 1 9 2
18 9 4 14 13 3 2 7 13 1 10 0 9 2 3 3 9 13 2
9 3 16 10 0 9 13 1 9 2
19 15 13 9 9 7 13 7 10 0 9 3 16 10 9 4 13 3 3 2
27 15 13 7 10 0 9 15 4 13 3 1 7 13 1 9 3 15 3 13 9 7 15 4 13 1 9 2
9 15 4 0 9 15 13 9 3 2
23 15 13 9 7 10 0 9 15 1 10 9 13 9 14 13 1 0 9 2 0 1 9 2
16 15 13 15 1 10 0 7 0 9 15 13 15 0 7 0 2
7 9 9 13 3 1 9 2
21 3 15 3 13 13 15 1 10 0 9 2 0 9 7 10 9 2 15 13 15 2
15 15 4 13 3 10 9 1 10 9 2 3 3 1 9 2
14 10 0 0 9 1 9 1 9 4 13 0 9 3 2
27 0 9 10 9 4 3 10 0 9 2 7 3 0 9 3 2 7 10 1 3 10 0 9 3 0 9 2
20 9 1 10 0 9 13 10 9 1 9 2 15 1 9 13 3 1 0 9 2
30 9 7 9 1 0 9 13 3 10 9 1 10 0 9 7 9 1 9 1 9 14 13 10 9 3 16 15 13 0 2
10 7 15 13 3 15 15 4 9 1 2
44 1 0 13 15 3 3 10 9 0 1 9 1 9 7 10 9 3 9 7 7 9 13 3 7 3 14 4 9 1 9 7 9 7 9 14 13 13 10 9 1 10 0 9 2
10 9 4 13 16 9 13 0 13 15 2
16 1 15 13 9 9 7 0 1 9 3 15 3 2 13 2 2
5 9 4 3 0 2
17 1 0 9 13 9 1 10 9 16 9 1 9 4 3 3 0 2
10 15 13 1 10 9 14 13 15 9 2
35 13 15 3 10 2 0 0 2 9 13 15 3 3 15 3 15 13 3 1 9 15 7 16 10 9 3 4 3 0 7 10 0 0 9 2
16 7 1 10 9 10 0 9 13 15 13 9 9 3 1 15 2
22 9 7 9 2 10 3 0 2 13 15 1 0 7 0 9 1 14 13 3 10 9 2
11 3 4 3 9 9 7 9 13 1 9 2
38 15 4 3 13 0 7 0 7 1 10 9 0 16 10 9 13 3 1 14 2 13 10 9 7 10 9 2 3 16 2 9 2 3 13 1 10 9 2
43 16 9 13 10 0 9 7 13 14 13 1 9 2 1 16 15 3 13 15 2 2 0 9 13 3 1 9 9 2 2 3 13 15 3 3 1 0 9 2 10 0 9 2
14 15 13 10 9 7 14 13 10 9 4 3 3 0 2
11 14 13 10 2 9 2 13 15 3 3 2
25 15 13 15 1 1 9 2 3 4 9 3 7 3 13 1 1 16 15 4 4 13 9 14 13 2
6 3 13 3 9 9 2
17 6 2 14 4 13 10 0 9 3 15 4 0 4 3 10 9 2
7 15 4 3 10 0 9 2
4 7 10 9 2
12 7 3 4 3 9 1 10 9 7 10 9 2
4 4 15 0 2
5 13 15 0 9 2
10 4 15 0 1 9 2 9 2 9 2
6 13 15 10 0 9 2
2 9 2
4 9 1 9 2
8 1 10 9 4 15 13 6 2
33 7 1 10 9 4 15 3 13 3 10 0 9 7 3 0 10 9 1 0 9 15 13 10 9 15 13 2 13 3 1 2 9 2
24 9 2 13 15 2 3 13 15 9 2 10 9 13 10 9 1 9 3 15 13 3 1 9 2
29 6 2 7 10 9 15 3 13 3 7 10 9 1 10 9 13 2 3 13 15 10 9 3 7 9 13 15 3 2
2 9 2
11 6 6 13 15 9 2 12 9 1 9 2
21 15 13 15 4 13 10 9 1 12 9 1 9 10 9 15 13 0 7 3 13 2
2 9 2
10 15 13 9 1 10 9 2 13 15 2
52 7 15 13 3 1 9 1 10 9 7 1 9 1 10 9 9 3 15 13 10 9 7 16 15 3 3 4 0 1 15 3 9 13 3 13 15 10 9 3 16 15 1 3 3 0 9 4 13 10 0 9 2
16 6 2 7 10 0 9 13 15 3 1 10 9 9 2 9 2
10 15 13 15 3 7 1 9 7 9 2
23 9 1 0 9 1 9 1 9 1 9 9 13 1 10 0 9 1 9 9 10 0 9 2
18 15 13 0 9 1 16 9 4 13 10 9 1 9 1 10 0 9 2
16 1 9 9 4 10 0 9 1 3 13 3 0 9 3 4 2
12 3 4 15 1 9 13 7 15 13 7 3 2
17 7 7 0 9 15 13 1 9 7 9 1 9 7 0 13 9 2
17 3 0 0 9 4 3 10 0 15 13 10 0 7 9 1 9 2
15 10 0 9 1 9 7 3 9 1 9 7 1 9 9 2
10 15 4 13 3 1 10 0 9 9 2
6 3 3 9 0 9 2
17 9 0 9 13 1 16 9 4 0 1 14 13 3 9 1 9 2
26 9 1 0 9 1 9 1 0 9 2 9 2 9 7 0 9 9 7 9 13 9 10 3 0 9 2
38 1 15 1 9 13 15 0 9 7 9 1 9 2 15 13 10 10 9 15 13 7 3 13 9 14 13 0 9 1 10 9 2 1 0 7 0 9 2
36 3 4 3 10 0 9 0 9 0 1 10 0 9 16 9 4 9 2 3 16 9 1 9 4 13 10 9 1 9 15 4 3 0 7 9 2
18 10 9 1 9 7 9 9 1 9 13 1 9 3 3 1 9 9 2
13 15 15 1 10 9 13 1 0 9 7 0 9 2
27 13 3 3 9 1 16 15 13 0 1 9 7 3 1 16 15 3 4 14 13 10 9 1 9 1 9 2
10 7 15 4 3 10 9 0 14 13 2
19 13 15 13 3 9 1 10 0 9 2 15 13 15 0 1 9 7 9 2
14 7 13 15 1 10 9 13 10 0 9 1 0 9 2
24 3 1 0 9 7 9 1 9 1 0 9 7 9 1 9 1 9 1 9 3 9 4 0 2
10 15 13 3 10 0 9 1 10 9 2
17 15 4 10 9 1 11 11 2 2 14 13 0 9 1 9 2 2
5 2 1 0 3 2
6 9 11 9 9 2 2
23 15 4 4 13 15 1 15 15 13 15 0 1 9 9 7 15 4 13 1 14 13 1 15
36 2 10 0 9 15 1 10 0 9 13 3 1 0 9 4 3 0 9 9 7 4 3 3 10 3 0 9 1 14 13 9 1 9 0 9 2
23 3 4 9 13 16 10 9 9 13 3 3 7 13 0 0 1 16 9 13 7 13 2 2
23 15 13 16 3 3 15 3 13 10 9 2 4 15 13 13 1 10 0 9 1 10 9 2
22 3 9 4 0 7 10 0 9 3 3 0 2 13 0 9 3 0 1 9 7 9 2
13 1 9 4 1 9 10 0 9 13 10 0 9 2
17 3 13 15 3 1 9 10 9 15 4 13 9 1 9 1 9 2
18 9 1 9 7 9 13 1 10 3 0 9 1 10 9 1 0 9 2
6 10 0 9 4 13 2
15 9 15 4 13 0 9 13 10 0 9 7 10 0 9 2
34 1 15 4 9 13 3 3 0 2 9 4 13 10 7 0 9 9 16 15 13 0 7 16 10 9 7 9 13 0 9 1 10 9 2
14 3 13 3 9 1 3 7 3 0 0 7 0 9 2
17 15 4 13 1 0 9 15 1 9 13 1 14 13 7 13 9 2
26 10 0 9 2 1 9 1 3 0 9 2 4 13 10 0 9 1 10 3 0 9 14 13 3 1 2
17 1 9 1 3 13 9 3 1 3 0 9 15 13 9 3 0 2
23 10 0 9 13 3 3 1 14 13 9 1 9 2 1 0 7 9 2 1 9 7 0 2
5 10 0 9 7 9
11 15 4 13 9 1 9 1 3 10 9 2
10 1 9 1 9 13 10 9 15 13 2
13 2 1 9 4 9 9 13 7 10 0 9 2 2
12 10 0 9 1 7 9 7 9 13 10 9 2
12 1 0 9 13 15 10 9 2 0 7 0 2
10 2 15 13 3 3 1 9 15 2 2
27 10 9 13 15 3 0 1 9 2 7 3 3 4 15 3 0 1 9 2 12 9 1 12 9 1 9 2
8 2 9 4 3 3 3 2 2
23 16 15 1 9 4 10 9 15 13 13 1 16 3 0 10 0 13 10 9 1 7 1 2
35 15 4 3 13 3 9 13 15 3 16 10 0 9 1 10 9 3 13 1 9 7 10 0 1 10 9 15 1 0 9 4 13 1 9 2
10 15 4 13 9 1 9 1 12 9 2
17 1 15 4 12 0 1 16 15 4 13 3 15 14 13 1 1 2
11 1 12 9 4 0 9 9 1 9 9 2
35 9 13 3 15 3 16 9 13 1 9 1 12 9 3 3 9 13 15 1 15 16 9 4 13 9 1 12 9 3 9 13 1 10 9 2
5 11 1 12 9 2
8 9 9 2 10 9 1 9 2
18 10 0 9 13 1 0 9 2 15 13 14 13 2 15 13 14 13 2
10 10 9 13 1 9 1 3 7 0 2
26 1 10 0 9 13 15 1 0 9 9 14 13 7 13 2 9 2 9 7 9 13 14 13 15 3 2
10 10 9 1 9 4 10 9 1 9 2
18 10 0 9 13 1 9 10 9 1 9 0 1 9 2 9 7 9 2
27 9 4 10 9 1 10 9 3 15 13 2 9 4 13 1 1 9 14 13 15 7 1 9 7 1 9 2
21 10 0 13 1 9 9 1 9 0 9 1 9 1 10 0 3 1 10 0 9 2
8 9 13 9 0 9 1 9 2
43 10 0 9 13 7 10 9 0 1 0 9 2 15 13 7 13 1 0 9 1 9 7 9 2 15 13 3 3 7 13 9 3 2 15 13 15 7 13 9 1 10 9 2
26 10 0 9 4 3 15 1 9 13 2 1 10 9 10 0 9 13 10 9 1 0 9 1 0 9 2
16 9 1 9 9 13 10 9 1 3 15 13 1 10 0 9 2
22 7 15 13 0 9 15 13 1 16 0 9 3 3 7 3 13 15 1 10 0 9 2
17 0 9 1 9 13 16 10 9 3 4 13 9 1 9 7 9 2
43 0 9 13 10 9 7 9 15 13 9 1 10 9 3 9 4 9 9 7 9 13 7 0 7 0 2 9 13 1 9 7 13 9 10 9 2 9 13 1 9 7 9 2
17 9 7 9 13 15 3 3 9 1 7 3 3 1 10 0 9 2
15 1 10 9 1 0 0 7 0 0 13 3 9 7 9 2
23 15 15 13 1 9 1 0 9 13 3 9 1 9 3 15 13 1 9 1 3 0 9 2
28 10 3 0 2 0 7 0 9 15 13 9 1 10 0 9 13 3 3 1 9 0 2 0 7 3 0 9 2
2 9 2
39 13 1 9 1 0 9 9 1 3 0 9 15 1 0 9 13 9 7 9 2 3 0 9 15 13 0 9 9 2 1 10 9 0 0 13 1 9 9 2
28 1 10 9 13 15 3 10 9 14 13 9 1 2 9 2 2 14 13 1 10 9 7 2 0 2 7 15 2
19 16 15 13 10 0 9 1 2 9 7 9 2 2 15 13 15 3 1 2
33 3 3 4 15 13 1 9 1 9 1 9 1 3 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2
15 3 13 15 1 10 0 9 9 1 10 0 1 9 9 2
10 2 13 10 0 9 1 0 9 2 2
13 13 15 10 9 14 3 13 3 15 7 13 3 2
14 4 15 1 3 9 10 9 15 15 4 13 7 13 2
14 13 13 3 9 1 9 13 3 3 1 11 3 3 2
11 13 15 0 2 0 9 1 10 0 9 2
6 1 3 9 2 3 2
10 2 13 3 9 9 12 7 12 2 2
14 9 1 9 9 13 3 3 4 3 3 7 3 0 2
43 15 1 9 4 9 9 1 9 0 7 3 0 7 3 2 15 3 16 10 0 9 1 9 7 9 9 13 15 3 3 0 2 10 9 2 15 13 14 13 0 7 0 2
65 9 13 3 3 10 9 7 10 9 1 0 9 2 15 13 3 10 9 7 13 3 10 9 1 9 2 15 13 1 9 0 9 7 13 10 7 0 9 1 9 9 2 9 7 9 1 9 2 2 15 13 15 7 13 15 7 13 3 7 3 1 10 0 9 2
45 3 15 13 9 7 15 15 3 13 2 13 3 3 9 1 9 9 2 15 13 15 14 13 1 15 2 15 13 15 1 0 9 2 15 13 3 14 13 1 9 2 3 1 15 2
26 1 9 13 3 9 2 9 7 9 1 10 2 0 2 7 2 3 7 3 3 2 10 9 7 9 2
28 15 13 1 9 7 3 1 9 2 15 4 0 7 9 7 13 15 3 3 9 1 15 1 10 0 0 9 2
29 9 13 10 9 1 9 9 2 15 15 3 13 4 10 0 9 7 9 1 15 15 13 1 9 7 9 1 3 2
50 15 13 15 15 3 4 10 0 9 1 9 2 7 9 13 3 3 3 1 0 9 2 7 9 2 9 2 0 9 1 3 2 15 4 3 13 1 10 0 9 1 9 7 9 2 1 9 7 9 2
18 9 1 9 9 4 1 9 13 1 10 0 9 7 13 1 9 0 2
43 9 4 3 3 13 3 10 9 2 15 4 13 10 9 7 10 9 1 0 9 2 15 4 13 9 1 9 1 9 2 15 4 13 10 9 7 9 1 9 7 0 9 2
31 15 4 3 13 14 13 9 1 10 2 0 2 2 3 16 15 1 9 1 9 7 9 13 1 15 10 0 9 7 9 2
40 3 4 9 4 13 15 3 16 15 4 13 3 9 2 3 9 7 0 1 9 3 16 15 3 1 10 9 15 13 2 3 4 14 4 13 15 7 9 9 2
49 10 15 4 14 13 10 9 7 15 4 13 1 14 13 9 13 1 1 9 2 9 7 9 1 9 1 14 7 3 13 1 10 9 1 16 15 13 15 10 0 9 7 9 7 9 1 9 9 2
