400 17
25 11 1 11 11 11 11 2 0 2 11 9 14 9 15 9 1 9 13 4 14 9 11 13 4 2
9 15 3 2 15 9 0 9 2 2
29 9 10 11 9 13 0 9 9 13 2 0 9 1 11 9 13 14 2 3 0 11 9 13 14 0 9 9 4 2
20 3 2 11 2 11 2 11 2 11 0 11 9 13 0 9 13 4 13 4 2
15 11 14 2 9 14 11 11 11 9 13 11 13 4 4 2
30 3 2 10 9 11 1 13 4 0 11 11 11 9 9 0 9 11 9 9 11 2 11 9 11 9 0 9 13 4 2
26 0 9 3 13 0 9 9 9 9 9 9 0 9 13 15 13 13 4 14 11 9 11 9 13 4 2
7 3 15 13 0 9 2 2
15 11 9 13 9 9 9 13 4 2 0 9 13 4 4 2
13 3 2 10 9 13 3 10 9 9 14 13 4 2
31 3 0 9 2 15 9 1 13 2 11 9 1 0 9 2 9 0 11 2 11 9 9 3 0 9 9 9 13 4 4 2
19 9 1 2 11 0 11 9 14 7 9 14 0 9 14 0 9 13 4 2
19 0 9 1 2 13 0 9 9 1 12 9 1 10 9 14 13 9 4 2
11 9 0 12 11 9 1 12 9 9 9 2
41 9 9 13 11 9 0 9 15 9 0 9 9 4 14 2 0 9 14 2 9 14 2 9 9 14 13 14 10 9 1 9 9 14 2 0 9 9 14 13 4 2
20 3 13 0 9 9 9 9 13 13 4 4 2 15 13 14 9 13 4 4 2
10 10 9 3 9 9 3 13 4 4 2
16 10 0 9 11 11 13 13 4 0 9 9 0 9 13 4 2
24 9 9 9 13 2 11 9 13 13 13 1 2 9 9 13 4 0 9 14 13 9 13 4 2
11 9 10 0 9 9 11 0 9 13 4 2
25 11 9 14 11 2 11 9 9 2 9 2 9 2 9 0 9 9 3 13 13 10 9 13 4 2
26 11 0 9 14 11 0 9 14 2 11 0 9 14 11 7 11 9 1 12 7 0 9 14 4 4 2
18 11 9 2 11 2 11 2 11 0 12 9 14 0 12 9 1 4 2
17 10 9 0 12 9 0 9 2 11 2 11 2 11 2 11 9 2
17 11 0 9 14 2 11 0 9 14 2 11 0 9 14 13 4 2
17 11 9 1 0 3 9 1 9 9 1 0 11 10 9 13 4 2
29 9 2 9 9 14 14 9 14 14 0 9 13 14 0 9 14 15 0 10 9 13 13 2 2 14 9 13 4 2
17 15 1 9 1 13 10 9 13 4 14 10 9 1 13 4 4 2
27 15 14 11 2 2 10 13 0 11 9 15 2 2 14 9 9 2 11 9 11 11 9 13 14 13 4 2
11 11 3 2 12 12 11 9 13 4 4 2
30 3 13 4 11 9 1 2 9 7 9 9 1 9 0 2 12 12 3 13 9 11 11 9 0 0 9 9 13 4 2
24 3 2 11 1 9 2 12 12 1 2 12 12 1 13 13 4 14 11 0 9 9 13 4 2
5 15 9 13 4 2
16 0 9 0 0 9 9 11 9 2 12 12 1 13 13 4 2
7 15 11 0 9 9 13 2
21 11 9 1 9 9 11 11 11 2 11 11 2 11 7 0 11 9 9 1 13 2
12 3 9 0 9 13 14 11 11 3 13 4 2
14 10 9 3 2 12 12 9 13 9 9 13 4 4 2
17 11 11 11 9 11 3 11 9 14 9 9 14 14 11 13 13 2
9 3 9 11 9 14 3 13 4 2
16 15 9 9 14 9 14 11 1 13 4 0 9 13 4 4 2
11 11 0 11 9 9 9 3 11 1 13 2
6 9 3 12 9 13 2
12 9 11 9 14 3 9 12 9 9 13 4 2
6 12 9 11 9 13 2
7 12 9 11 11 9 13 2
7 15 1 0 9 9 13 2
45 9 12 9 9 1 9 9 13 9 9 12 9 1 9 9 13 4 4 2 9 12 9 9 13 2 9 13 2 9 9 9 1 2 9 0 9 9 9 2 11 9 9 13 4 2
27 11 1 9 11 11 9 9 13 14 13 4 2 15 9 9 13 4 14 11 9 0 9 11 11 9 13 2
25 0 9 9 13 4 14 0 11 2 10 9 14 9 13 13 4 15 9 10 11 13 13 4 13 2
31 11 13 0 11 11 9 3 13 9 13 2 3 13 14 0 11 2 3 10 9 9 3 13 0 9 9 1 13 13 4 2
12 11 0 9 9 0 9 11 11 9 13 4 2
22 3 11 9 1 9 9 0 14 11 9 13 4 14 10 9 9 9 9 11 11 13 2
11 11 9 1 10 9 13 4 14 15 13 2
21 11 0 9 11 9 9 3 13 1 11 11 11 9 14 11 11 9 3 9 13 2
10 11 1 11 9 15 3 9 11 13 2
11 3 11 11 1 15 15 0 9 13 13 2
28 11 11 11 9 11 14 14 0 11 2 11 3 9 11 9 1 9 4 4 0 9 9 13 4 14 13 4 2
28 11 1 9 14 12 9 9 0 0 11 9 14 9 0 11 9 11 9 14 10 9 13 4 4 14 9 13 2
26 11 11 9 9 9 14 11 12 11 9 1 13 15 1 12 9 14 13 14 10 11 9 11 11 13 2
23 11 9 14 11 11 11 1 0 0 9 1 13 1 9 13 13 14 11 9 0 14 13 2
25 9 11 9 9 9 13 0 9 0 9 13 0 14 10 11 13 14 0 9 9 9 11 11 13 2
14 11 0 12 9 13 4 4 14 11 11 9 13 4 2
32 9 0 9 11 11 9 13 0 11 11 9 9 11 9 13 0 0 9 11 11 2 11 13 11 9 11 9 9 1 13 4 2
28 10 9 11 9 13 9 13 4 4 14 14 2 15 13 0 12 9 13 4 4 14 14 11 11 9 13 4 2
21 11 9 13 4 14 0 9 9 15 9 9 13 14 11 11 11 11 9 11 13 2
13 11 9 13 4 0 12 11 9 3 9 13 4 2
18 9 9 13 14 15 9 13 4 4 14 9 0 9 15 13 4 4 2
18 3 2 12 9 0 9 9 4 4 14 11 9 9 9 11 11 13 2
19 9 9 9 0 9 9 13 0 9 3 9 14 9 13 4 14 13 13 2
25 15 0 9 14 12 0 9 13 14 3 0 9 9 1 13 4 4 14 10 9 9 11 11 13 2
18 11 9 14 12 0 9 13 14 11 9 9 11 9 9 9 13 4 2
22 9 12 12 9 14 13 14 14 2 15 3 13 4 14 14 10 9 9 13 4 4 2
25 3 11 9 14 0 9 12 9 13 14 14 2 15 3 12 9 14 13 4 14 14 15 13 4 2
19 15 9 1 9 9 0 11 2 15 1 9 1 15 3 13 4 4 13 2
19 11 9 13 0 11 9 11 9 9 4 4 14 11 11 11 9 13 4 2
35 11 11 0 11 9 3 0 9 3 9 13 4 0 11 11 9 9 11 11 2 11 11 2 11 11 9 11 11 9 0 3 3 13 4 2
10 3 15 9 13 4 4 14 13 4 2
32 10 9 2 3 9 0 11 11 9 9 11 11 2 2 9 13 0 12 9 14 11 9 13 11 11 11 9 14 13 14 4 2
12 3 11 11 9 14 0 3 13 4 2 13 2
28 3 3 15 1 11 11 9 13 4 14 13 0 15 2 9 1 9 13 14 9 9 13 4 4 14 14 13 2
13 3 15 9 4 0 9 13 14 15 3 13 4 2
9 11 9 9 11 9 11 11 13 2
19 11 1 9 0 9 1 11 0 11 2 3 9 1 11 9 9 9 13 2
20 0 9 11 11 9 14 9 11 11 9 11 2 11 11 11 9 11 9 13 2
13 3 11 9 11 9 9 11 9 9 0 9 13 2
19 3 2 11 9 11 11 9 14 2 11 9 11 11 9 14 9 13 4 2
13 3 11 2 11 2 11 0 9 14 9 13 4 2
17 11 11 9 0 11 0 9 11 2 11 9 11 2 11 9 13 2
11 3 13 0 9 9 0 9 11 13 4 2
18 11 11 9 12 9 1 13 4 0 9 9 13 4 14 11 9 13 2
15 11 9 0 9 9 1 11 9 2 9 12 2 13 4 2
14 9 9 3 0 11 13 1 2 11 10 9 13 4 2
19 11 3 13 0 9 9 7 9 9 9 15 1 14 0 3 13 4 4 2
17 0 9 9 1 13 4 15 9 13 4 2 9 11 1 13 11 2
7 0 9 11 9 9 11 2
10 11 9 14 0 15 2 0 9 13 2
16 11 2 9 2 11 2 9 0 9 13 14 2 13 14 9 2
16 11 2 9 9 11 9 0 11 2 11 9 1 9 9 13 2
12 9 9 9 14 2 9 2 15 11 9 13 2
20 0 9 9 9 14 14 2 9 7 9 9 9 7 9 9 14 14 9 13 2
8 0 9 11 11 9 14 13 2
20 0 9 9 7 9 9 9 14 14 2 0 9 9 9 9 14 14 9 13 2
12 0 9 9 9 7 9 9 9 9 14 13 2
14 0 9 1 12 9 9 7 9 9 0 9 3 13 2
8 0 9 9 9 9 9 13 2
12 0 0 9 9 9 7 9 9 3 13 4 2
9 3 2 9 9 3 9 13 4 2
10 0 11 9 11 11 9 9 3 13 2
11 15 1 0 9 9 9 14 9 11 13 2
11 12 9 0 9 9 9 3 13 11 11 2
7 3 12 9 1 9 13 2
14 11 0 9 11 9 1 15 9 9 13 4 13 4 2
9 9 0 3 9 15 13 14 2 2
11 9 0 9 11 11 9 9 13 13 4 2
18 10 9 9 15 14 13 9 9 1 15 0 9 9 3 13 13 11 2
18 9 9 9 1 9 13 14 2 11 9 9 1 11 13 4 14 13 2
13 0 9 9 11 9 13 4 14 9 11 9 13 2
12 11 9 9 14 9 13 0 11 9 9 13 2
23 9 9 9 9 13 1 11 9 13 4 2 11 9 9 9 15 13 13 14 9 13 4 2
24 11 2 9 9 14 9 11 9 9 9 7 9 9 9 14 12 0 9 14 9 13 4 4 2
14 9 9 3 11 14 2 11 11 3 11 11 14 4 2
15 9 9 0 10 12 0 9 14 9 13 4 4 13 4 2
8 11 11 9 13 0 9 13 2
13 12 11 9 0 9 13 14 11 9 9 11 13 2
16 11 11 9 1 0 9 13 9 4 2 12 12 9 4 4 2
28 11 11 9 9 9 11 9 9 0 14 2 11 9 9 1 9 9 9 3 13 0 9 13 14 9 13 4 2
13 9 0 9 11 9 3 0 9 11 9 13 4 2
29 3 11 11 9 11 9 3 0 9 2 9 11 9 13 9 11 9 9 14 11 9 1 0 9 11 9 13 4 2
15 9 1 9 9 4 4 2 0 9 13 14 11 9 13 2
6 9 13 14 11 9 2
8 15 14 0 9 14 13 4 2
15 10 9 13 4 9 9 12 12 12 9 9 9 13 4 2
6 12 12 9 9 13 2
13 3 13 0 9 12 9 14 14 14 11 13 4 2
7 9 13 0 9 3 13 2
10 11 9 9 11 9 9 14 10 9 2
9 3 2 11 9 9 1 9 13 2
14 0 0 9 11 0 9 11 9 3 13 9 4 4 2
9 11 11 9 0 9 10 9 13 2
15 10 9 9 0 9 9 13 4 14 9 13 4 4 11 2
24 11 9 13 4 9 9 13 0 11 11 0 9 14 13 14 11 9 9 9 11 11 9 13 2
17 11 13 0 11 11 2 3 9 9 13 0 11 13 9 9 13 2
7 11 1 9 15 9 13 2
9 0 9 9 2 9 13 13 4 2
25 2 15 3 15 13 15 3 4 2 3 3 13 14 9 9 1 14 9 9 0 11 15 9 4 2
18 11 1 9 1 11 11 9 0 15 3 3 9 1 11 13 13 4 2
6 11 0 9 15 13 2
13 9 11 14 9 0 11 9 12 9 9 15 13 2
13 0 11 9 2 9 11 11 9 11 1 3 13 2
19 9 0 9 13 4 0 11 13 15 11 9 14 11 11 9 14 15 13 2
10 3 11 0 9 9 1 15 9 13 2
28 11 15 0 9 3 13 1 14 9 9 0 11 14 9 9 14 9 9 13 4 1 14 9 9 1 15 13 2
14 9 9 0 11 9 11 9 13 0 14 15 9 13 2
17 9 11 14 11 9 11 11 9 9 11 11 7 11 9 14 13 2
13 3 9 13 13 4 0 11 9 0 9 15 13 2
11 11 9 0 9 11 1 12 9 13 4 2
18 11 9 0 3 11 3 13 4 14 13 2 11 9 13 4 11 9 2
17 11 11 13 3 2 9 9 11 9 14 9 9 11 14 9 13 2
18 11 0 14 9 9 11 11 7 11 9 9 1 15 9 13 14 13 2
5 11 1 9 2 2
11 9 11 9 11 7 9 9 11 11 13 2
17 11 14 11 9 7 0 9 1 11 3 12 12 12 9 13 4 2
14 3 11 9 0 12 12 11 11 9 14 11 13 4 2
18 15 1 9 2 11 9 0 12 9 12 11 9 14 3 13 4 4 2
11 9 7 9 9 1 12 9 11 13 4 2
9 3 12 12 9 9 14 11 13 2
11 11 0 9 13 10 9 9 13 4 4 2
18 3 9 7 9 9 11 1 12 12 9 13 14 14 14 11 13 4 2
12 3 2 9 9 9 0 9 9 11 13 4 2
18 9 9 13 2 9 2 11 9 2 11 9 9 0 9 11 13 4 2
20 11 0 11 11 9 9 9 1 13 11 9 0 9 9 13 14 9 13 4 2
18 11 0 11 9 12 13 13 14 11 1 12 11 0 9 9 13 4 2
14 9 9 11 1 9 0 11 9 11 11 9 13 13 2
16 9 13 0 14 15 9 1 3 13 11 9 9 13 14 13 2
8 10 9 11 11 9 13 4 2
21 11 9 1 11 9 1 9 0 9 13 14 14 15 15 13 4 4 14 13 4 2
12 3 15 1 0 9 14 10 9 9 13 4 2
37 3 12 9 9 10 11 9 15 11 9 9 13 4 4 14 14 2 11 1 14 2 11 11 9 1 14 13 15 9 13 4 14 14 10 9 13 2
17 15 10 9 14 4 0 9 0 14 15 11 9 13 14 14 13 2
18 9 9 13 2 9 9 4 4 2 9 0 14 15 11 9 13 4 2
7 15 3 11 13 14 13 2
13 9 11 9 11 1 0 0 9 11 9 12 13 2
4 12 9 13 2
27 11 9 9 9 0 10 9 9 9 0 11 11 9 9 11 11 11 9 14 13 14 9 11 9 11 13 2
11 0 9 0 11 11 0 9 10 9 13 2
12 3 11 1 0 11 9 9 3 13 9 13 2
12 11 9 9 0 9 11 9 11 9 13 4 2
18 11 13 0 9 1 2 11 9 0 12 9 9 13 14 11 3 13 2
11 11 0 9 13 4 0 9 9 9 4 2
27 11 9 13 4 0 12 9 9 4 9 0 9 9 13 4 4 14 0 9 9 13 0 9 13 4 4 2
28 15 1 2 11 7 11 9 1 0 12 9 14 2 11 9 1 9 14 2 11 9 1 12 9 14 13 4 2
12 0 12 9 13 4 4 14 9 9 13 4 2
15 10 9 3 12 9 13 4 2 11 1 11 13 4 4 2
20 3 3 12 9 13 4 4 13 10 9 0 12 9 11 9 13 4 13 4 2
17 11 11 9 9 11 11 11 13 11 9 14 9 9 11 13 4 2
9 9 9 0 9 9 15 3 13 2
10 2 11 11 9 13 4 7 13 4 2
10 11 9 15 9 14 0 9 3 13 2
15 3 9 10 0 9 14 9 14 9 14 9 14 13 4 2
16 11 9 9 3 10 0 9 14 14 13 14 14 11 13 4 2
29 11 11 9 9 11 11 9 0 9 13 13 9 9 9 1 9 13 4 14 11 9 0 9 11 11 9 13 4 2
24 9 11 9 2 11 9 7 9 2 0 9 9 9 9 1 13 14 3 9 11 11 13 4 2
32 10 9 2 9 0 9 14 11 9 0 9 14 14 11 11 2 9 9 1 9 13 4 4 14 11 11 13 4 9 13 4 2
16 15 3 2 9 9 11 11 9 9 1 13 4 14 13 13 2
9 11 9 9 0 9 11 9 4 2
24 11 2 11 2 11 2 11 2 11 2 11 0 12 9 0 0 12 9 9 12 11 9 4 2
22 11 9 11 9 9 9 3 0 11 11 11 9 9 0 9 9 9 0 9 13 4 2
22 3 3 9 0 9 11 11 2 2 11 2 11 9 9 9 9 13 4 2 14 13 2
17 11 9 9 2 12 9 14 0 9 12 9 9 15 9 9 13 2
22 11 11 9 2 12 12 9 9 9 14 9 9 11 11 2 11 11 11 11 9 13 2
12 3 2 11 0 11 9 9 12 3 13 4 2
17 9 2 11 11 2 11 11 11 9 12 12 9 9 9 9 13 2
14 3 2 9 14 12 12 9 11 11 9 9 13 4 2
27 0 3 9 13 13 4 14 0 9 3 9 13 4 14 11 9 0 9 11 11 13 4 14 9 13 4 2
16 3 13 0 11 9 9 13 13 4 0 9 11 9 13 4 2
19 9 2 9 3 0 14 2 11 0 9 13 14 11 11 9 9 13 4 2
5 2 15 15 13 2
3 13 4 2
9 15 9 9 14 9 11 1 13 2
7 3 2 15 14 3 13 2
23 15 9 9 13 14 7 0 9 9 14 13 4 14 0 9 3 15 1 14 9 13 4 2
18 2 14 9 13 0 15 9 1 11 13 14 10 11 9 13 4 4 2
15 11 11 9 9 9 13 14 9 9 9 9 11 13 4 2
11 3 15 3 13 0 9 13 4 14 2 2
25 11 11 9 9 9 9 0 9 1 11 11 9 13 4 14 13 0 9 0 9 14 9 14 13 2
29 11 11 9 1 9 9 13 0 11 11 13 13 0 11 9 9 13 3 12 9 14 0 0 11 13 14 13 4 2
15 3 9 9 9 0 0 9 0 9 3 0 9 13 4 2
48 11 14 11 9 14 9 9 13 9 1 9 9 9 13 4 14 9 1 9 0 0 9 13 0 9 2 0 9 15 3 0 9 9 9 9 4 0 9 9 0 9 9 15 14 13 14 4 2
10 0 9 10 9 9 9 9 3 13 2
12 11 0 9 3 13 4 14 14 11 1 13 2
13 11 9 0 9 9 9 13 15 14 9 13 4 2
12 3 0 9 11 9 9 0 9 9 15 13 2
17 11 0 11 9 7 9 15 11 9 0 9 9 13 4 14 13 2
7 3 11 15 9 13 4 2
16 11 9 9 9 9 13 4 14 11 11 9 11 11 13 4 2
10 3 15 3 13 0 9 4 14 2 2
19 11 9 9 13 9 0 9 2 12 9 11 1 12 11 9 9 4 4 2
7 9 9 9 9 11 13 2
18 3 2 9 9 9 13 12 11 11 0 9 14 15 9 9 4 4 2
18 9 9 1 0 9 3 13 11 9 9 4 14 13 11 9 14 9 2
19 9 0 9 2 9 2 9 2 9 9 9 14 0 9 0 11 9 4 2
14 3 2 3 11 9 13 4 3 9 9 9 13 4 2
8 3 11 11 15 9 13 4 2
29 11 11 11 9 9 1 9 9 9 13 13 0 11 9 13 3 3 9 11 1 9 13 14 9 9 11 13 4 2
11 3 15 3 13 0 9 13 4 14 2 2
11 11 2 11 9 0 11 9 9 13 4 2
20 11 13 0 2 11 2 11 9 12 9 14 0 11 9 9 9 13 13 4 2
48 11 9 9 2 11 11 11 11 9 1 0 9 9 1 9 0 9 9 9 1 13 4 9 13 14 9 3 13 4 14 14 2 3 10 0 9 9 11 9 13 4 4 14 14 9 9 13 2
39 3 9 9 9 1 9 9 13 9 9 3 13 4 14 14 2 9 13 0 9 13 14 14 2 9 9 3 13 2 9 9 13 4 14 14 9 9 13 2
20 11 11 9 9 0 9 11 9 2 15 13 13 9 0 9 11 9 13 4 2
55 11 11 11 9 9 9 1 11 9 13 13 0 11 9 13 14 2 3 15 13 13 13 14 2 11 9 2 11 9 11 1 2 12 9 9 9 12 9 9 2 11 9 9 1 11 11 9 9 11 11 9 11 9 13 2
7 3 11 15 9 13 4 2
8 11 9 9 9 12 9 13 2
17 11 9 0 11 9 9 2 9 9 0 9 12 9 0 9 13 2
8 3 2 9 9 12 9 13 2
15 11 9 11 9 9 9 0 11 12 9 0 9 1 13 2
12 3 2 10 9 13 11 9 14 12 9 13 2
13 9 0 9 7 9 9 0 9 11 3 13 4 2
17 11 2 12 9 1 9 9 1 3 3 12 14 0 9 13 4 2
10 12 9 13 4 14 11 9 13 4 2
11 11 9 11 9 1 9 13 12 9 13 2
10 9 9 11 9 0 11 9 9 13 2
8 0 11 11 9 9 13 4 2
11 3 2 11 11 13 3 9 13 4 4 2
12 3 2 9 13 14 9 9 14 13 4 4 2
13 3 2 15 13 9 9 9 9 13 13 13 13 2
11 3 2 0 9 0 9 11 1 3 13 2
9 9 2 11 9 14 12 9 13 2
6 10 9 12 9 13 2
8 15 3 9 0 9 13 4 2
8 3 2 9 9 9 3 13 2
9 9 11 9 9 11 11 9 13 2
9 10 9 9 15 9 9 9 9 2
19 9 11 9 9 13 11 13 4 3 11 11 11 11 9 9 9 13 4 2
27 11 9 9 11 2 11 9 12 0 9 9 13 4 1 15 0 0 9 12 14 0 9 9 9 13 4 2
7 3 11 9 13 4 4 2
11 9 2 9 11 11 9 9 13 4 4 2
7 3 11 9 13 14 2 2
11 9 11 9 9 9 12 9 0 11 13 2
11 15 2 11 9 9 11 3 9 4 4 2
11 3 2 15 13 0 9 12 9 13 4 2
15 9 9 3 0 14 9 13 14 11 13 14 11 9 13 2
17 10 9 9 11 1 11 11 9 11 9 11 9 9 11 13 4 2
14 11 12 11 0 12 9 13 4 14 11 9 13 4 2
12 11 0 9 9 11 0 0 9 9 13 4 2
26 9 11 9 11 9 0 11 11 9 9 1 14 11 11 9 11 9 1 14 9 9 13 14 13 4 2
24 3 12 11 0 12 9 13 14 11 11 9 9 9 2 11 1 0 9 12 0 9 13 4 2
9 3 15 11 0 11 9 13 4 2
9 11 15 13 4 14 9 13 4 2
12 11 9 9 9 9 11 9 9 4 13 4 2
13 3 12 9 9 1 11 9 0 9 9 13 4 2
8 0 9 11 9 9 13 4 2
18 11 9 9 9 9 9 0 9 9 3 13 0 11 9 1 13 4 2
6 3 11 9 13 4 2
21 11 2 11 2 11 11 9 0 9 0 0 9 14 13 10 9 9 13 13 4 2
8 9 9 12 9 14 9 13 2
13 10 12 11 11 2 11 2 11 0 12 9 13 2
7 11 9 11 9 13 4 2
16 3 12 0 11 9 14 11 2 11 2 11 0 9 13 4 2
28 0 9 9 9 11 2 11 2 11 2 11 0 9 10 0 13 14 11 9 9 14 11 9 11 11 11 13 2
15 11 9 9 9 9 13 9 9 12 12 9 9 13 4 2
7 3 11 12 9 9 9 2
9 3 0 9 9 9 11 13 4 2
22 9 9 9 0 9 3 0 11 2 11 2 11 2 11 2 11 9 9 9 13 4 2
8 3 0 9 11 0 9 13 2
15 11 9 9 9 9 13 4 4 4 14 11 3 13 4 2
23 11 9 13 12 9 2 11 2 11 2 11 2 11 2 15 9 9 13 4 14 9 13 2
11 0 9 9 0 9 9 0 9 1 13 2
18 0 9 11 0 12 9 9 9 9 9 9 9 4 4 1 13 4 2
15 3 9 4 4 1 3 13 4 14 14 3 9 13 4 2
22 11 9 9 0 14 2 11 7 9 1 9 9 13 4 14 11 9 9 11 11 13 2
4 15 10 13 2
12 3 0 9 13 9 3 13 14 15 3 13 2
21 11 9 11 11 2 11 0 9 9 9 0 14 10 9 1 3 13 4 14 13 2
14 11 9 9 9 11 11 11 9 11 11 13 4 4 2
20 9 1 11 11 9 14 11 9 9 9 9 14 14 11 11 2 10 9 13 2
10 10 9 9 3 0 9 1 11 13 2
12 9 11 9 7 9 11 9 13 9 13 4 2
7 0 9 10 9 13 4 2
7 3 12 9 9 13 4 2
12 11 11 9 9 11 11 11 0 9 9 13 2
19 11 9 11 11 0 9 3 0 11 9 11 9 11 11 9 9 9 4 2
16 11 11 2 0 9 0 11 9 11 9 11 11 9 3 13 2
9 3 2 11 0 9 14 15 13 2
9 11 11 10 9 11 0 9 13 2
8 11 9 11 9 9 9 13 2
16 11 11 9 0 11 9 1 0 9 13 4 14 14 13 4 2
13 3 11 11 9 1 11 9 2 11 9 9 13 2
11 11 11 1 0 9 14 14 14 9 13 2
9 9 11 11 15 9 9 4 4 2
18 3 15 9 2 15 9 14 2 9 14 9 9 13 14 15 13 4 2
7 9 0 13 15 13 4 2
18 15 9 15 9 14 13 4 13 0 14 3 12 9 13 4 4 13 2
14 11 11 0 0 11 11 9 1 0 9 9 13 4 2
12 15 2 11 0 9 14 11 1 9 13 4 2
17 13 0 9 13 0 14 10 9 11 9 9 11 11 9 13 4 2
10 9 13 9 1 0 9 14 13 4 2
11 2 12 12 9 13 4 14 15 13 4 2
8 0 9 15 14 9 13 4 2
5 15 9 13 4 2
16 9 9 13 4 14 13 15 13 13 4 14 14 11 11 13 2
8 11 0 11 11 9 9 13 2
15 10 9 11 0 9 3 11 0 0 11 9 13 9 13 2
11 11 9 3 0 9 9 9 11 9 13 2
18 9 0 12 9 11 9 9 14 12 9 14 2 3 12 9 14 13 2
17 9 0 9 9 9 9 3 0 9 11 9 3 9 9 3 13 2
9 9 9 13 9 9 13 13 4 2
12 11 9 11 9 9 11 11 11 11 9 13 2
8 3 0 9 9 11 11 13 2
20 0 11 12 14 9 0 11 2 0 12 11 14 12 2 12 14 9 9 13 2
11 3 12 14 11 9 11 13 11 9 13 2
5 11 9 9 13 2
15 11 13 0 9 1 11 0 11 9 9 12 3 13 4 2
9 15 1 11 9 11 0 9 13 2
9 12 11 9 0 11 0 9 13 2
23 11 9 11 11 13 9 13 11 3 9 0 11 9 9 11 0 9 14 9 9 13 4 2
20 11 3 0 11 9 9 9 0 9 3 13 13 14 11 9 11 13 4 4 2
25 15 9 9 13 11 2 9 9 2 11 9 9 2 11 11 9 1 9 11 0 9 9 13 4 2
16 11 11 11 1 11 9 11 9 0 9 11 11 9 13 4 2
13 3 2 9 0 11 0 9 14 9 9 9 4 2
23 3 11 11 9 11 11 9 7 9 9 9 9 11 9 2 11 9 2 11 9 9 13 2
6 3 15 9 9 4 2
21 9 9 13 14 0 9 9 11 9 0 14 13 4 14 11 9 11 9 9 13 2
20 9 0 12 11 9 1 9 0 14 9 9 13 4 14 9 9 11 9 13 2
17 3 9 11 1 9 13 4 4 15 13 4 14 9 9 11 13 2
16 3 11 9 1 9 9 0 9 9 13 4 9 9 13 4 2
17 11 9 13 11 1 9 9 0 9 14 9 0 9 14 13 13 2
9 11 9 0 9 0 9 13 4 2
6 3 9 9 9 4 2
17 3 11 0 9 9 9 0 9 0 9 13 14 9 9 4 13 2
15 9 0 9 14 12 9 0 9 9 9 9 12 9 13 2
26 9 13 14 11 2 11 2 11 2 11 2 11 1 11 9 0 9 9 9 14 9 0 9 13 13 2
12 0 9 9 9 14 9 0 9 9 13 13 2
17 9 9 13 0 11 9 9 13 3 11 9 0 9 3 13 4 2
24 12 9 12 11 1 11 13 4 9 13 0 9 9 0 0 11 9 10 0 9 9 13 4 2
8 3 11 9 9 3 13 4 2
14 9 9 13 9 9 14 9 10 13 14 11 9 13 2
13 3 9 7 9 9 9 2 11 9 13 4 4 2
12 3 0 9 13 0 9 15 13 14 9 4 2
22 11 11 1 13 4 9 13 0 12 9 1 9 0 9 0 9 11 9 9 13 4 2
13 11 9 13 4 14 9 7 9 9 11 9 13 2
44 11 11 11 9 9 11 9 0 9 9 2 11 11 9 9 9 11 9 1 0 9 9 9 2 11 9 7 9 9 9 2 11 9 9 9 9 13 4 9 11 13 14 2 2
15 11 11 9 9 14 15 9 11 9 1 9 13 4 4 2
7 15 0 9 1 13 4 2
12 10 9 1 13 4 0 9 1 13 4 4 2
20 11 9 9 11 9 0 9 13 4 4 14 9 0 9 3 11 9 13 4 2
19 15 13 2 11 9 9 9 14 3 0 9 13 4 14 9 15 1 13 2
35 3 2 11 9 15 13 2 15 11 9 9 14 13 4 2 10 9 3 11 9 9 9 9 13 4 0 9 15 1 0 9 1 13 4 2
41 11 0 9 9 15 11 9 1 0 9 3 3 11 9 1 13 0 9 13 14 14 2 11 9 9 13 0 9 2 10 9 3 13 4 14 0 9 13 11 14 2
6 11 9 14 9 13 2
7 3 15 12 3 13 4 2
18 3 2 10 3 10 9 13 4 3 0 12 12 12 9 13 4 4 2
15 10 9 13 4 2 15 11 9 9 9 9 13 4 4 2
6 9 9 13 3 13 2
9 3 3 9 14 9 13 3 13 2
31 10 9 14 1 0 9 2 10 9 3 0 9 0 0 9 9 15 15 14 0 9 13 14 13 10 9 15 13 13 4 2
19 10 9 11 11 9 15 13 14 10 9 13 9 13 4 2 9 13 4 2
5 9 9 13 2 2
14 9 13 4 14 9 2 9 0 11 9 15 13 4 2
