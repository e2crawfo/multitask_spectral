2077 11
7 15 16 11 13 1 11 2
23 15 16 11 13 1 15 9 2 9 2 7 3 9 2 9 1 10 3 2 0 9 9 2
9 2 1 11 11 1 11 11 11 2
25 2 7 2 1 10 9 2 13 9 0 3 10 0 9 1 10 9 3 15 13 10 0 9 2 2
31 10 11 9 13 16 11 14 9 1 9 4 13 2 10 15 4 3 13 3 2 7 15 13 3 3 2 13 1 10 9 2
7 11 13 10 0 9 9 2
8 4 9 13 15 1 9 0 2
7 15 13 11 2 3 3 2
6 13 15 10 9 9 2
8 15 4 13 3 1 10 9 2
28 15 13 10 3 0 15 3 13 15 9 4 14 13 1 15 3 2 7 15 13 15 4 13 15 3 3 3 2
22 11 11 1 11 4 13 1 10 0 9 9 16 15 4 3 13 7 13 1 1 11 2
6 13 3 14 13 15 2
12 15 13 10 0 9 1 10 0 1 10 9 2
13 12 1 10 9 13 10 9 10 4 13 1 11 2
13 1 10 0 12 9 15 13 9 1 12 9 9 2
8 13 10 9 1 10 11 9 2
11 15 13 14 13 10 9 2 15 13 0 2
24 10 11 9 4 13 1 14 13 10 3 0 9 13 1 10 11 9 1 10 9 1 10 9 2
42 13 15 13 10 9 1 9 1 11 14 0 9 2 10 2 16 13 1 10 13 9 2 13 3 3 10 9 10 0 9 4 13 2 7 13 1 10 0 0 9 3 2
12 15 13 14 0 1 10 11 2 13 2 9 9
81 2 15 4 14 13 14 13 15 9 2 15 4 13 2 1 16 13 15 9 2 15 4 14 13 14 13 9 1 9 1 10 11 9 2 7 16 2 9 1 9 2 15 13 0 16 15 4 13 9 1 9 15 4 13 10 9 1 9 15 4 3 13 15 1 10 11 9 2 15 13 3 2 3 3 0 9 1 15 9 2 2
9 3 2 10 9 13 3 0 9 2
10 1 10 0 9 2 15 13 3 0 2
12 11 13 15 4 13 0 9 16 13 0 9 2
10 10 11 11 4 14 13 10 0 9 2
7 15 4 13 10 0 9 2
6 7 15 13 10 9 2
26 15 13 10 9 1 11 11 13 10 0 9 16 13 0 14 13 10 0 9 7 15 13 1 10 9 2
18 15 4 3 13 0 1 10 11 11 11 11 1 9 1 10 9 9 2
27 10 11 4 3 13 15 4 13 14 13 11 13 1 10 9 10 15 4 14 3 13 14 13 1 0 9 2
13 7 15 4 13 16 15 13 0 9 1 0 9 2
13 0 9 13 14 13 9 1 11 1 1 0 9 2
5 7 4 9 13 2
9 7 4 9 13 0 9 1 9 2
19 12 9 13 1 16 10 11 13 10 11 1 10 9 3 15 13 15 9 2
5 15 4 13 15 2
8 15 4 14 13 14 13 15 2
7 7 15 4 14 13 15 2
16 15 4 13 16 11 3 13 9 7 3 13 1 9 1 9 2
33 0 9 13 0 9 1 10 0 9 1 11 2 9 12 2 16 10 9 9 13 1 10 0 9 9 1 11 9 4 13 1 11 2
44 11 13 16 2 0 9 1 10 9 13 10 2 9 1 10 9 1 11 2 13 10 9 1 10 9 9 7 9 2 13 12 9 1 9 2 7 13 1 10 0 9 9 2 2
25 15 13 2 2 10 9 1 11 13 10 9 10 4 13 1 11 1 9 0 1 10 9 1 11 2
34 13 0 2 0 2 9 7 9 13 16 15 13 0 16 13 10 9 14 9 7 9 2 7 13 15 14 13 15 9 1 10 9 2 2
9 10 9 13 9 1 0 11 9 2
32 11 4 3 4 13 1 0 9 1 10 11 9 3 2 16 0 11 7 13 0 1 0 9 7 4 13 0 9 7 3 9 2
22 9 0 1 11 13 0 9 1 11 7 13 10 0 9 1 10 9 14 9 7 9 2
28 15 13 16 10 0 9 13 1 15 10 9 2 7 10 9 1 10 11 7 11 2 7 15 13 14 13 3 2
2 13 8
46 10 11 11 13 15 9 9 1 11 1 11 13 1 0 9 16 11 11 13 1 1 15 9 1 10 11 11 9 7 11 11 13 10 9 1 10 12 5 12 9 10 13 12 9 0 2
8 10 0 9 13 10 0 0 2
76 13 1 15 3 2 11 11 11 13 10 9 1 10 9 1 9 1 9 12 1 12 2 12 1 12 2 9 2 12 2 12 2 9 2 12 2 7 12 2 1 10 11 2 11 2 11 2 7 11 13 2 7 10 9 1 9 1 9 12 7 12 2 9 2 12 2 1 10 11 2 11 2 7 11 13 2
16 9 13 10 13 9 2 1 10 11 2 11 2 7 11 13 2
24 11 13 10 9 13 1 0 2 1 10 11 2 11 2 7 11 13 1 1 9 12 7 12 2
13 11 13 10 13 9 2 1 10 11 7 11 13 2
36 11 13 10 13 9 2 1 10 11 13 2 7 1 10 11 13 1 1 10 7 9 12 2 12 2 9 2 12 2 7 12 2 9 2 12 2
19 11 13 10 13 9 2 1 10 11 7 11 13 1 1 9 12 1 12 2
24 15 4 13 15 10 0 9 14 13 10 0 9 2 7 15 3 13 1 10 11 11 11 9 2
14 15 4 13 9 1 10 9 7 9 3 15 13 0 2
75 0 9 0 1 11 11 14 0 9 1 15 9 9 5 0 2 9 2 15 13 14 1 9 1 10 9 2 3 1 10 9 2 3 3 3 15 9 4 14 3 4 13 1 7 4 4 3 13 2 4 13 11 3 3 1 10 0 9 2 7 10 9 9 2 7 1 1 10 11 11 7 11 11 3 2
11 15 13 14 13 1 10 11 1 10 9 2
52 15 13 0 2 15 13 2 1 15 0 2 13 2 12 9 9 2 9 9 2 16 10 0 0 2 9 0 9 1 10 9 4 3 4 13 2 16 15 11 1 11 13 0 1 15 9 9 2 1 10 9 2
5 15 13 3 0 2
27 3 0 2 3 2 13 10 9 16 10 0 9 14 13 10 9 13 10 0 0 9 3 13 14 4 13 2
24 1 10 9 2 11 11 11 11 11 13 9 4 13 14 13 10 0 9 1 11 1 12 9 2
9 12 9 3 2 7 10 9 13 2
30 10 11 11 13 3 14 1 1 10 9 16 13 10 9 2 13 12 9 1 10 9 10 4 13 12 2 13 1 9 2
22 7 0 9 4 13 3 9 1 10 9 9 10 11 13 2 13 1 10 0 11 9 2
34 3 3 15 13 2 12 9 3 2 1 10 0 11 9 12 9 3 1 11 7 11 2 7 10 9 1 10 9 1 11 13 3 0 2
20 11 11 4 13 1 12 5 1 15 9 2 3 1 10 11 7 11 11 11 2
50 15 13 10 9 10 3 13 15 2 11 14 0 9 16 13 0 1 15 9 13 16 15 4 3 13 10 9 1 15 9 1 10 3 0 9 2 3 10 9 3 4 13 3 0 9 1 10 9 3 2
39 15 13 10 0 0 14 13 2 7 1 10 9 15 0 9 13 16 10 11 13 3 0 9 2 9 2 7 15 13 15 14 13 10 9 3 3 16 0 2
17 10 3 13 16 15 13 0 16 11 7 11 4 13 14 13 3 2
26 15 13 15 0 9 13 16 15 13 0 16 11 11 3 4 14 13 3 3 14 13 15 0 9 9 2
10 15 13 14 0 3 10 9 4 13 2
32 15 4 14 13 10 9 14 0 9 2 7 16 10 9 13 2 10 9 4 4 13 1 10 0 9 16 10 9 13 3 0 2
35 1 10 0 9 2 15 13 3 10 9 16 10 9 13 0 1 10 9 15 13 15 3 2 7 13 14 13 10 0 9 1 10 0 9 2
30 6 2 6 2 10 11 9 3 13 1 0 9 7 9 2 15 13 13 3 13 10 0 9 13 16 13 1 12 9 2
12 16 10 12 9 13 1 9 4 3 13 0 2
2 8 2
35 15 4 14 13 12 5 1 2 15 4 13 10 9 1 9 10 9 10 13 1 9 1 10 9 1 12 5 10 9 2 16 0 2 2 2
12 15 13 15 9 14 9 13 10 9 1 15 2
46 15 13 3 0 16 15 4 13 16 11 7 11 13 1 10 0 9 2 3 13 10 9 9 3 13 10 0 9 2 7 11 4 3 13 0 1 15 9 1 1 11 3 15 4 13 2
38 11 3 1 10 11 11 13 10 0 9 16 3 10 11 7 10 11 2 3 10 0 9 1 11 2 4 3 13 0 9 1 0 9 1 10 0 9 2
29 1 10 0 9 11 13 1 9 1 11 7 11 2 10 0 9 11 4 13 15 4 13 1 10 13 0 0 9 2
26 1 10 9 1 11 2 15 13 0 9 1 11 16 13 10 0 0 9 1 9 1 11 14 13 9 2
20 11 4 13 14 13 1 10 9 13 3 1 11 11 12 2 10 4 3 13 2
32 11 11 2 11 11 11 4 13 15 13 9 14 2 13 11 2 16 3 4 13 1 2 10 9 1 10 9 15 4 13 2 2
22 10 9 1 3 0 9 1 0 9 9 13 10 0 9 1 10 11 11 7 10 9 2
46 3 12 9 1 12 2 10 11 11 2 1 15 9 14 13 9 16 13 9 2 3 4 14 3 13 10 9 2 9 2 2 13 1 10 9 16 16 10 9 1 0 9 13 0 9 2
26 10 9 3 13 10 9 1 9 7 0 9 2 16 10 0 9 1 11 11 1 10 11 11 11 13 2
1 5
42 10 9 14 13 10 0 14 13 10 9 14 13 9 4 14 13 9 2 7 3 13 10 0 9 16 10 9 1 11 7 11 13 10 0 9 1 10 9 7 10 9 2
35 15 4 4 13 1 10 9 1 10 0 9 3 2 3 16 10 9 7 9 13 15 13 14 13 10 9 16 11 4 13 0 16 13 11 2
4 15 13 15 2
9 15 13 10 0 9 0 7 0 2
28 15 13 10 9 10 13 15 11 9 1 12 2 13 11 9 1 10 9 7 3 15 4 4 13 10 0 9 2
17 15 13 3 10 9 14 3 13 10 11 2 7 3 3 10 11 2
31 10 11 11 11 13 1 11 11 11 2 4 13 1 10 0 0 0 9 0 14 13 2 3 16 3 3 2 1 10 11 2
13 15 4 3 13 14 13 1 1 10 11 9 9 2
34 10 11 4 3 13 10 0 9 13 0 11 14 13 1 10 9 13 1 11 2 7 4 4 13 1 10 9 1 10 11 1 11 11 2
40 16 10 11 11 11 4 3 13 13 10 11 9 13 10 9 16 16 10 0 0 11 9 1 10 9 13 1 10 9 2 3 3 13 10 9 1 10 0 9 2
22 11 2 11 2 10 11 1 11 11 13 11 14 13 1 10 9 1 11 1 10 11 2
46 1 10 9 2 10 11 13 16 16 11 14 13 9 1 2 13 9 2 1 10 9 1 10 9 2 10 9 1 10 13 0 2 0 1 11 2 4 4 13 10 3 0 1 0 9 2
32 10 0 11 13 11 2 2 15 13 3 15 13 1 9 9 1 10 9 1 11 2 7 13 16 15 13 10 0 9 1 11 2
8 13 16 10 9 13 0 2 2
23 10 0 0 11 9 13 10 9 13 10 9 1 0 9 1 10 9 1 11 2 3 3 2
70 10 9 13 2 2 15 13 10 9 1 10 9 1 10 0 9 2 16 0 9 7 9 2 10 9 1 15 13 0 2 13 1 15 14 13 16 13 10 0 9 1 10 9 1 9 10 4 14 13 15 9 7 10 9 1 0 9 2 7 15 13 15 14 13 10 9 1 0 2 2
19 15 13 10 2 9 2 10 9 16 10 9 13 3 1 0 9 1 11 2
47 10 9 1 9 1 10 3 0 0 0 9 1 11 7 10 0 11 1 10 11 9 4 4 13 3 2 0 9 1 10 0 11 9 1 11 7 1 10 11 9 1 11 11 9 1 11 2
30 0 11 2 3 2 13 3 0 14 13 0 9 14 13 10 11 1 11 2 0 1 15 4 13 11 7 15 0 9 2
13 11 11 13 10 0 9 9 1 15 9 1 9 2
5 11 2 11 2 2
35 11 0 9 13 11 11 1 11 16 13 10 13 9 14 13 1 9 9 1 10 2 9 1 0 9 2 2 13 10 9 4 13 0 9 2
28 11 9 4 13 10 9 2 13 1 11 2 14 13 1 0 9 1 10 11 13 0 1 10 9 1 11 11 2
43 2 15 13 15 13 10 3 2 13 9 7 15 13 16 15 13 0 14 13 11 7 11 1 9 2 2 13 11 11 2 0 9 1 10 11 1 11 2 11 11 9 9 2
15 10 13 3 15 4 14 13 15 13 1 9 1 0 9 2
8 15 13 1 9 1 0 9 2
23 16 13 10 9 2 0 2 1 10 9 11 4 3 14 13 11 1 9 2 3 10 9 2
25 7 16 15 4 14 13 1 3 2 10 9 1 13 9 13 3 10 11 2 11 7 11 1 15 2
7 11 11 2 12 2 11 11
8 11 11 11 2 12 2 11 11
7 11 11 2 12 2 11 11
8 11 11 11 2 12 2 11 11
7 11 11 2 12 2 11 11
8 11 11 11 2 12 2 11 11
7 11 11 2 12 2 11 11
6 11 11 2 12 2 11
7 11 11 2 12 2 11 11
8 11 11 11 2 12 2 11 11
8 11 11 11 2 12 2 11 11
8 11 11 11 2 12 2 11 11
8 11 11 11 2 12 2 11 11
7 11 11 2 12 2 11 11
12 11 11 2 12 2 2 13 11 11 2 11 11
7 11 11 2 12 2 11 11
7 11 11 2 12 2 11 11
8 11 11 11 2 12 2 11 11
33 11 11 2 12 2 11 11 16 15 13 0 1 10 9 1 10 0 9 13 1 11 10 0 9 3 2 11 11 2 12 2 11 2
9 11 11 2 12 2 11 2 11 2
7 11 11 2 12 2 11 2
7 11 11 2 12 2 11 2
8 11 11 11 2 12 2 11 2
9 11 11 2 12 2 11 2 11 2
8 11 11 11 2 12 2 11 2
7 11 11 2 12 2 11 2
8 11 11 11 2 12 2 11 2
11 11 11 11 9 11 11 2 12 2 11 2
8 11 11 11 2 12 2 11 2
11 11 11 2 12 2 1 11 11 2 11 2
29 15 4 13 10 11 2 10 12 9 10 4 14 13 15 9 2 9 2 16 15 4 13 1 10 11 11 11 11 2
16 9 2 16 15 13 0 2 7 0 2 15 13 10 0 9 2
29 7 16 15 4 14 13 14 13 0 15 4 13 9 13 10 0 9 7 13 9 9 3 0 16 15 4 3 13 2
53 1 10 9 9 1 11 7 11 11 2 11 2 11 11 11 2 11 2 2 10 9 3 13 2 2 15 13 16 10 11 7 11 11 2 15 9 7 9 2 4 13 9 1 10 9 1 10 9 11 11 11 2 2
7 10 9 13 10 0 9 2
25 11 11 11 2 11 7 15 9 4 13 14 4 13 0 9 1 11 2 11 1 10 0 9 9 2
34 12 9 1 10 11 9 1 11 13 16 11 4 14 13 11 7 11 11 14 13 9 1 11 2 11 1 10 0 9 1 10 0 9 2
30 16 10 9 13 0 2 15 13 10 0 9 16 3 10 13 0 0 9 9 4 4 2 13 3 2 1 11 2 11 2
21 10 9 13 3 10 9 1 11 14 0 9 1 11 7 1 10 9 1 10 9 2
10 15 13 10 9 1 10 9 1 9 2
26 11 2 11 1 11 13 10 9 1 3 10 0 12 2 0 11 2 15 13 0 9 1 11 11 11 2
28 15 4 3 4 13 14 13 10 12 2 0 2 11 11 2 1 10 11 9 2 16 15 13 14 10 0 9 2
33 16 11 13 0 2 15 9 13 16 15 4 3 13 1 10 9 9 1 10 0 9 1 11 10 13 1 11 14 10 12 12 9 2
36 1 12 15 4 13 1 11 1 10 11 2 11 11 2 11 9 1 11 11 2 11 2 0 1 15 13 1 11 11 2 3 11 7 9 2 2
30 1 10 9 2 11 2 11 13 10 0 9 1 10 0 9 7 10 9 11 1 11 11 2 3 10 1 15 13 0 2
27 11 13 10 11 2 7 15 11 7 11 11 9 1 11 3 13 10 0 9 1 3 0 2 0 7 0 2
14 15 3 13 10 0 9 1 10 9 1 11 7 11 2
37 15 4 3 3 13 1 10 0 9 1 0 0 9 2 10 13 10 11 2 0 9 16 13 3 1 10 0 9 1 10 0 9 1 10 11 11 2
30 2 0 11 13 14 0 7 0 2 16 15 13 14 13 3 0 2 0 1 15 9 2 1 10 9 1 11 9 2 2
31 11 7 11 11 3 4 13 10 0 9 1 11 2 3 16 10 10 9 1 10 3 2 13 11 11 11 1 0 11 13 2
33 10 0 9 13 16 0 0 0 9 13 1 10 11 9 1 11 4 13 13 11 7 11 11 2 7 13 15 0 0 7 0 9 2
16 15 4 4 13 1 0 9 1 11 11 1 11 7 1 11 2
19 3 3 15 13 9 1 11 2 11 9 1 11 3 15 4 13 9 3 2
57 10 9 1 0 0 0 0 9 1 11 2 11 4 3 4 13 1 10 9 1 10 11 9 1 9 10 13 16 10 11 11 11 11 2 13 9 15 13 1 11 12 9 11 11 2 7 3 13 1 0 0 1 10 11 9 9 2
11 10 11 11 11 4 13 15 9 1 11 2
20 15 13 12 9 1 10 10 11 13 0 9 10 4 4 13 11 11 14 9 2
11 12 1 15 13 1 11 7 12 1 11 2
32 11 13 3 9 7 13 16 16 15 4 13 15 4 13 2 15 4 4 13 10 9 14 13 15 2 7 16 3 4 13 11 2
17 10 9 13 2 1 15 9 1 0 2 9 2 3 0 9 9 2
17 3 3 11 4 4 13 14 13 12 16 15 4 13 15 4 13 2
14 10 9 13 2 2 4 15 4 13 15 4 13 2 2
8 10 9 13 2 2 6 2 2
15 15 3 13 16 11 7 15 9 13 1 9 0 1 11 2
26 11 4 13 1 9 1 11 9 9 7 13 1 9 1 11 9 3 2 3 1 11 7 11 1 12 2
52 11 13 9 9 11 11 3 10 0 13 1 10 11 2 11 9 2 13 16 10 0 9 1 9 1 10 11 13 1 11 2 7 13 15 13 11 11 14 9 9 9 16 11 13 1 10 12 11 11 11 9 2
48 16 15 13 9 9 3 16 13 1 10 9 2 15 13 10 11 2 11 9 3 13 1 1 11 2 11 11 2 11 2 10 0 9 9 13 1 11 11 2 3 15 4 13 1 10 0 9 2
14 3 1 10 9 1 11 12 2 11 4 13 1 11 2
21 11 13 1 15 7 13 16 15 13 10 12 1 12 5 9 16 11 13 1 15 2
5 2 1 10 9 2
24 10 9 13 3 11 2 11 2 7 10 0 9 1 11 2 11 7 11 4 3 4 13 2 2
24 11 3 13 10 9 1 11 2 11 9 1 11 2 13 15 13 2 10 0 9 2 1 11 2
24 2 15 1 12 11 2 11 9 10 4 13 10 12 9 7 0 9 13 1 10 11 11 2 2
29 10 11 4 14 3 13 10 9 16 13 1 11 7 11 2 11 10 15 4 13 1 10 9 2 13 1 11 11 2
10 11 4 14 13 15 9 1 10 9 2
9 7 13 11 2 11 2 7 11 2
12 15 4 13 11 11 1 11 14 0 0 9 2
31 0 9 13 10 9 16 9 1 9 1 10 11 7 0 9 3 1 10 11 9 13 3 1 11 11 7 10 9 15 13 2
11 15 4 1 10 9 13 7 14 13 1 2
22 11 13 11 11 2 1 10 3 0 7 0 1 10 11 2 11 9 2 1 15 9 2
57 11 4 3 3 13 10 0 9 1 10 9 9 2 15 13 15 2 7 15 4 14 13 15 14 13 1 9 9 1 10 9 1 12 3 11 11 14 9 13 2 1 9 2 1 10 0 9 10 11 4 13 1 1 0 11 9 2
15 1 1 10 11 9 2 13 15 13 12 9 1 15 9 2
39 11 4 13 1 10 9 1 0 11 11 11 11 1 9 1 12 10 4 4 13 10 11 14 13 10 0 9 9 3 1 11 11 1 11 2 13 1 11 2
16 15 13 15 13 10 11 9 1 9 9 16 9 9 13 0 2
7 15 3 13 0 9 9 2
10 10 9 13 3 0 7 4 4 13 2
16 7 1 9 1 12 2 11 11 11 13 10 9 1 11 11 2
22 10 0 9 13 0 1 9 0 1 10 11 2 7 10 0 0 9 13 1 10 9 2
21 11 13 11 15 4 14 13 0 9 7 9 9 14 13 10 9 3 1 11 11 2
29 13 1 10 9 7 15 13 14 13 1 3 2 1 9 1 12 2 15 4 3 13 1 10 10 9 1 0 9 2
12 3 3 2 15 4 3 13 3 1 0 9 2
18 7 1 15 1 15 13 1 10 9 2 6 13 1 11 14 11 9 2
6 15 4 4 3 13 2
7 11 13 2 7 13 3 2
10 10 9 13 14 1 15 1 10 12 2
15 15 13 3 15 13 15 14 13 1 15 1 2 10 9 2
6 15 4 14 13 3 2
4 15 13 10 9
1 6
3 13 0 2
16 13 14 13 1 9 1 15 16 15 13 15 2 11 9 2 2
6 3 13 14 3 13 15
5 15 13 2 15 2
7 15 4 13 15 13 3 2
6 15 4 15 13 9 2
3 1 15 2
7 15 4 13 1 10 0 9
4 15 13 0 2
6 15 13 14 13 12 2
5 15 13 0 9 2
5 9 9 13 0 2
11 3 4 15 13 15 4 13 12 1 15 2
8 4 14 13 15 13 0 9 2
3 0 9 2
21 15 13 0 2 15 4 14 13 14 13 15 3 2 15 3 13 14 13 10 9 2
4 15 4 14 13
13 15 4 13 9 10 13 10 9 2 1 11 14 2
9 9 10 13 1 5 12 10 9 2
10 6 2 15 4 13 9 1 11 14 2
7 15 4 13 3 0 3 2
5 15 4 15 13 2
6 15 4 13 9 0 2
3 0 9 2
2 6 2
3 15 9 2
17 15 4 4 13 15 13 1 1 10 0 9 15 13 10 9 1 2
2 9 2
12 3 2 15 13 10 9 15 15 4 13 1 2
8 15 4 4 13 1 9 0 2
14 15 4 14 3 13 11 2 15 4 14 13 1 15 2
5 11 13 11 11 2
7 15 13 15 13 10 9 2
2 6 2
6 15 13 15 9 3 2
15 15 13 14 13 1 1 10 9 11 1 10 0 9 9 2
5 15 13 1 15 2
7 15 13 10 9 10 9 2
11 4 15 13 1 1 10 0 9 11 9 2
6 6 15 4 14 13 2
6 15 13 3 0 9 2
4 4 15 13 2
6 15 13 1 1 9 2
5 15 13 1 11 2
10 15 4 13 15 9 3 15 13 3 2
6 15 13 0 15 13 2
15 11 4 14 13 3 0 16 0 1 10 9 13 9 9 2
6 9 4 13 0 3 2
7 3 15 4 14 13 15 2
8 15 4 3 13 13 0 9 2
17 15 13 16 0 4 4 13 3 1 9 1 10 0 9 7 3 2
12 9 13 15 16 11 4 13 10 9 1 9 2
11 15 13 14 0 3 0 15 13 2 3 2
11 15 4 13 14 13 16 15 4 13 9 2
2 11 11
2 12 12
2 11 2
5 6 1 11 11 2
15 15 3 13 15 9 7 15 3 13 16 11 13 10 9 2
9 15 4 13 10 0 9 1 11 2
17 15 13 10 9 10 15 13 7 15 4 13 9 1 11 13 9 2
11 15 4 14 13 3 3 15 4 13 3 2
24 11 11 7 11 11 11 4 13 10 9 3 7 15 13 0 15 4 3 13 1 15 1 15 2
13 15 13 0 3 10 9 13 0 1 10 0 9 2
25 3 15 13 15 2 15 4 13 14 13 3 1 15 9 7 9 7 10 12 9 4 13 15 0 2
19 15 4 14 13 16 15 13 9 15 4 13 7 15 13 3 0 14 13 2
3 0 9 2
1 11
8 10 9 13 10 11 11 9 2
9 3 15 13 9 1 15 9 9 2
19 11 11 11 11 11 9 9 9 7 9 9 2 12 9 2 12 9 2 8
4 0 11 11 2
34 13 1 1 15 7 11 11 14 9 1 11 11 2 15 4 13 14 13 10 13 9 2 13 1 10 1 11 11 11 11 7 11 11 2
19 11 11 11 11 11 9 9 9 7 9 9 2 12 9 2 12 9 2 8
3 14 13 3
3 6 11 2
18 15 13 15 4 4 13 0 1 10 10 9 2 3 15 4 14 13 2
6 13 15 4 4 13 2
7 13 15 16 15 13 9 2
1 11
3 6 13 3
2 11 2
13 15 13 3 12 9 1 10 9 15 13 0 9 2
6 0 9 9 9 0 9
6 11 11 5 12 5 12
5 11 5 12 5 12
1 2
5 9 5 12 5 12
11 6 13 15 13 16 15 13 10 0 9 2
1 11
13 14 0 2 7 15 13 16 10 9 9 13 15 2
5 13 15 1 9 2
6 15 4 13 14 13 2
10 15 4 13 14 13 3 1 15 3 2
2 3 2
5 15 13 10 9 2
3 6 11 2
7 13 16 15 4 13 0 2
2 0 2
1 11
6 6 2 15 13 9 2
14 4 15 13 10 9 1 10 9 9 10 15 13 9 2
54 15 13 15 13 3 10 0 9 2 13 15 9 13 1 10 3 3 0 9 1 9 2 13 15 9 1 10 9 3 0 2 7 13 11 1 1 10 11 11 9 1 10 9 14 13 11 14 0 9 2 10 0 9 2
2 6 2
8 6 2 4 14 15 13 15 2
19 15 4 14 13 9 2 7 15 13 16 15 4 13 10 9 3 1 11 2
17 15 13 14 0 2 7 15 13 16 15 13 13 9 9 2 3 2
20 15 4 13 15 1 1 9 7 1 10 9 7 13 16 15 4 13 15 1 2
5 0 9 1 11 2
4 15 13 0 2
22 15 13 14 3 13 10 9 1 11 1 11 16 15 13 10 0 9 14 13 10 9 2
22 10 9 13 3 7 3 11 13 2 10 9 9 4 13 14 13 1 10 9 1 9 2
14 3 14 13 10 9 4 13 14 4 13 1 11 9 2
15 4 14 13 1 10 0 11 9 16 15 13 10 0 9 2
41 16 9 4 13 1 9 2 15 4 13 14 13 10 9 1 10 9 16 11 4 13 1 10 11 11 2 16 11 2 11 2 11 13 1 1 10 0 12 9 2 2
24 3 2 4 14 13 9 16 15 13 10 0 9 2 10 9 15 13 13 10 11 9 0 9 2
1 8
1 8
1 8
1 8
1 8
8 15 13 0 9 16 15 13 2
7 11 1 11 3 15 13 2
14 15 13 0 15 4 4 13 15 14 13 15 10 9 2
6 3 4 11 13 1 2
8 15 4 14 13 15 14 13 2
8 15 4 3 13 14 13 3 2
10 15 13 3 0 14 13 15 10 9 2
5 11 4 13 1 2
2 11 2
29 15 4 3 13 14 13 10 9 9 9 2 3 16 10 9 9 4 13 0 14 13 10 9 1 9 1 10 9 2
18 3 1 15 9 2 15 9 1 9 4 13 10 9 1 10 9 9 2
15 15 4 3 13 12 5 13 13 1 10 12 9 13 9 2
18 9 1 9 2 9 4 13 1 10 9 1 1 12 5 7 12 5 2
18 4 12 1 15 9 9 13 10 0 12 9 9 9 1 9 2 9 2
9 3 2 15 4 13 10 0 9 2
22 1 9 2 13 15 9 15 4 13 10 9 1 11 9 7 10 9 2 9 9 9 2
25 10 9 9 4 3 13 16 15 13 10 9 7 4 3 4 0 13 10 9 9 1 10 9 3 2
10 0 1 10 9 7 9 15 4 13 2
1 11
2 11 2
12 15 13 15 1 10 9 9 0 9 1 11 2
7 15 13 15 9 3 3 2
21 15 4 13 16 15 4 13 15 10 9 13 10 9 1 9 9 1 10 9 9 2
3 13 15 2
38 11 11 11 9 11 11 11 11 7 11 11 11 11 11 2 11 2 12 2 12 0 9 12 11 11 2 11 2 12 2 12 9 11 2 11 12 8 9
2 8 8
3 12 12 9
12 15 4 13 10 11 2 11 2 11 11 9 2
11 10 9 14 13 15 2 3 13 15 9 2
20 3 2 15 13 10 9 1 11 11 7 15 13 16 11 4 13 15 5 12 2
19 11 4 13 14 13 11 2 11 2 11 7 10 9 2 0 9 7 9 2
10 15 4 3 13 10 7 10 9 9 2
20 10 9 13 16 15 14 13 1 1 15 9 7 16 15 14 13 1 3 3 2
15 15 4 13 11 11 14 13 10 9 9 13 10 10 9 2
3 6 13 2
2 8 8
3 12 12 9
17 11 2 3 13 10 9 1 9 9 13 1 15 1 9 1 12 2
8 6 13 9 1 15 0 9 2
10 13 15 1 15 9 16 13 10 9 2
10 11 7 11 2 11 2 9 12 13 12
19 11 11 11 7 11 2 11 2 9 12 2 9 12 7 9 12 13 12 2
11 11 11 11 9 9 2 11 11 12 11 12
5 15 13 1 9 2
16 16 10 9 13 3 3 2 15 4 13 15 1 2 9 9 2
4 11 11 2 8
3 12 12 9
16 4 15 13 15 3 1 11 14 13 11 13 1 9 3 3 2
17 15 4 13 15 9 1 10 9 1 9 9 1 10 9 1 11 2
20 3 2 10 9 3 13 14 2 13 2 10 9 10 4 13 3 2 6 13 2
12 15 13 1 11 14 9 13 1 15 0 9 2
8 4 14 13 10 9 10 9 2
2 2 11
8 11 2 4 15 13 9 3 2
12 15 13 1 1 10 9 16 15 13 0 9 2
15 16 13 9 14 13 10 9 4 15 14 13 13 9 0 2
2 11 2
13 13 3 4 11 11 14 9 13 10 13 11 11 2
11 15 4 13 10 9 11 11 9 9 3 2
1 11
11 9 2 0 1 10 9 16 13 15 3 2
14 6 13 3 15 4 13 14 13 9 0 1 15 9 2
2 9 2
1 11
2 11 2
32 15 13 1 11 11 2 12 2 9 2 7 12 2 9 2 2 15 13 1 15 16 10 9 13 10 13 12 5 12 13 9 2
10 6 13 10 13 9 1 9 1 15 2
2 9 2
1 11
13 15 9 11 11 13 9 2 9 9 14 13 15 2
7 15 4 13 3 1 11 2
27 11 11 11 0 9 12 11 11 2 11 12 11 2 11 12 9 2 2 12 2 12 9 2 2 12 2 12
2 9 2
1 11
2 11 2
37 3 15 13 10 0 2 9 2 1 15 9 9 10 4 13 1 15 0 9 1 2 8 2 11 0 2 2 8 2 9 9 2 2 8 2 0 2
21 15 4 13 10 9 1 10 11 0 9 12 7 13 1 15 9 1 11 11 11 2
14 10 9 13 15 2 9 2 2 3 15 4 13 0 2
1 11
2 11 2
21 16 11 4 13 9 2 4 15 6 13 10 2 0 9 9 12 2 1 10 9 2
4 3 15 0 2
12 9 2 0 1 9 9 3 16 15 13 9 2
2 9 2
1 11
6 11 11 11 2 11 2
3 6 11 2
33 15 3 13 14 13 1 16 16 15 4 13 10 9 14 13 10 9 9 9 9 2 0 1 9 1 10 9 3 13 1 11 2 2
22 15 13 15 4 14 13 9 9 3 3 3 15 4 13 10 0 9 0 1 10 9 2
4 9 7 9 2
30 11 11 11 9 9 9 9 11 11 11 2 11 9 2 2 12 2 12 9 2 2 12 2 12 9 2 8 2 8 2
2 8 8
3 12 12 9
2 11 2
29 15 4 13 16 15 4 13 0 16 15 14 13 3 1 15 12 9 14 13 10 0 9 1 15 9 1 10 9 2
20 11 4 13 15 16 15 13 16 15 4 13 15 3 13 10 9 1 10 9 2
25 15 13 10 0 0 9 4 13 9 0 2 3 3 4 14 13 10 0 9 14 13 1 15 9 2
29 7 13 15 13 16 15 4 13 10 9 2 9 2 7 3 3 10 9 3 3 1 15 3 15 13 10 0 9 2
12 15 13 15 4 13 15 3 3 1 15 9 2
2 9 2
1 11
11 10 0 13 9 9 1 11 13 9 12 2
1 11
1 11
40 15 3 13 10 9 1 10 9 1 10 9 1 12 5 9 1 9 9 12 9 2 12 1 5 12 2 4 15 13 15 7 11 11 13 15 10 9 9 13 2
1 9
2 11 2
14 15 13 16 15 3 13 12 1 9 9 1 10 9 2
1 11
4 11 12 2 12
10 11 11 12 2 11 11 2 12 2 11
7 11 11 11 11 12 2 11
4 11 12 2 12
10 11 11 12 2 11 11 2 12 2 11
7 11 11 11 11 12 2 11
4 11 12 2 12
10 11 11 12 2 11 11 2 12 2 11
7 15 4 13 3 1 15 2
4 3 1 12 2
18 15 13 10 0 9 2 3 15 4 13 14 13 15 3 10 0 3 2
6 13 15 4 13 3 2
1 11
1 2
6 13 1 10 0 9 2
1 2
9 15 1 9 13 15 1 5 12 5
1 2
1 11
5 15 4 4 13 2
2 11 2
5 9 1 10 9 2
9 13 16 10 9 13 10 0 9 2
23 15 13 15 4 14 13 2 7 15 4 13 9 14 13 15 1 10 9 9 9 1 8 2
17 16 15 13 14 13 10 9 9 9 1 1 0 9 2 13 0 2
16 16 15 13 10 9 9 1 10 9 9 2 13 15 10 9 2
2 9 2
31 11 11 2 2 8 2 9 2 11 11 12 11 11 2 11 2 11 12 2 12 2 12 2 9 2 12 2 12 9 2 8
8 2 8 8 2 8 2 9 12
2 11 11
10 6 13 15 10 9 14 13 11 9 2
2 11 11
10 13 15 0 1 9 10 9 10 9 2
20 3 2 15 13 10 0 9 1 10 11 9 1 11 15 13 15 13 14 13 2
11 10 9 13 1 12 2 11 1 11 11 2
8 4 13 16 15 14 13 15 2
10 15 4 13 12 1 15 9 1 11 2
2 11 11
9 11 3 13 10 9 9 15 13 2
9 15 4 13 15 10 9 1 9 2
1 11
21 4 12 1 15 6 13 15 10 9 1 10 0 9 15 13 1 11 9 9 9 2
22 16 15 4 13 0 7 0 1 10 9 2 15 4 13 14 13 10 9 1 0 9 2
2 9 2
27 11 11 11 11 11 11 2 11 2 0 9 8 2 12 2 12 9 2 12 2 12 9 2 12 2 12 9
5 9 13 0 12 2
4 9 13 0 2
8 15 13 0 10 9 7 11 2
8 15 3 13 1 10 11 9 2
14 15 9 13 14 4 13 1 1 9 9 2 9 9 2
4 13 15 3 2
7 13 15 0 1 9 9 2
10 15 13 14 13 1 10 9 1 9 2
8 13 15 13 16 15 13 0 2
24 11 11 0 9 11 11 2 9 9 2 2 12 2 12 9 2 2 12 2 12 9 9 2 8
10 13 15 0 1 9 10 9 10 9 2
20 3 2 15 13 10 0 9 1 10 11 9 1 11 15 13 15 13 14 13 2
11 10 9 13 1 12 2 11 1 11 11 2
8 4 13 16 15 14 13 15 2
10 15 4 13 12 1 15 9 1 11 2
2 11 11
3 6 13 15
3 3 12 2
24 11 11 0 9 11 11 2 9 9 2 2 12 2 12 9 2 2 12 2 12 9 9 2 8
5 9 13 0 12 2
4 9 13 0 2
8 15 13 0 10 9 7 11 2
8 15 3 13 1 10 11 9 2
14 15 9 13 14 4 13 1 1 9 9 2 9 9 2
4 13 15 3 2
7 13 15 0 1 9 9 2
10 15 13 14 13 1 10 9 1 9 2
8 13 15 13 16 15 13 0 2
24 11 11 0 9 11 11 2 9 9 2 2 12 2 12 9 2 2 12 2 12 9 9 2 8
1 8
3 12 12 9
5 13 1 2 8 8
10 15 13 3 0 16 15 14 13 9 2
10 15 4 13 14 13 15 1 10 9 2
6 13 15 1 15 9 2
11 10 11 13 1 1 11 1 12 1 12 2
12 1 11 1 10 9 10 11 4 13 1 12 2
14 10 11 3 13 1 10 9 1 12 1 11 1 12 2
26 1 11 1 12 10 11 4 13 1 12 2 3 14 13 1 10 3 0 9 1 12 1 11 1 12 2
11 10 11 3 13 1 12 1 11 1 12 2
22 1 11 1 12 10 11 4 13 3 1 12 2 3 14 13 1 12 1 11 1 12 2
25 10 0 9 3 13 10 11 2 0 2 1 10 0 9 1 12 1 11 1 12 2 13 9 0 2
12 7 1 11 1 12 10 11 4 13 1 12 2
21 13 15 13 0 2 1 11 1 12 10 11 4 13 1 10 9 9 9 1 12 2
27 1 10 9 2 10 9 7 9 1 11 11 4 13 10 12 11 7 0 4 13 3 1 10 9 1 9 2
7 3 3 2 15 13 10 9
17 7 15 13 10 9 10 0 9 9 1 10 11 13 15 9 3 2
27 1 0 12 9 13 0 2 15 13 0 2 15 4 13 2 1 2 15 4 13 11 11 2 0 1 0 2
9 6 2 15 13 3 16 13 15 2
2 11 11
3 12 12 9
17 15 4 14 13 3 1 12 2 7 4 13 15 3 12 1 11 2
3 0 9 2
2 11 11
2 11 11
3 12 12 9
2 3 2
15 1 10 9 2 11 14 9 9 4 4 13 1 12 9 2
3 11 11 11
3 12 12 9
24 10 9 1 10 11 9 9 9 13 1 11 4 4 13 1 10 1 15 1 10 0 12 9 2
28 16 15 4 13 2 0 11 9 2 11 4 13 10 9 1 11 14 9 7 9 9 14 13 10 11 9 9 2
16 15 13 1 11 11 2 7 15 13 16 10 13 9 13 0 2
9 13 4 10 9 10 13 10 9 2
10 10 9 1 10 13 9 13 12 9 2
15 10 9 1 10 11 9 9 13 10 13 9 1 12 9 2
46 1 9 2 15 13 10 9 1 12 9 10 13 10 9 1 10 9 9 2 0 0 2 10 11 13 1 10 11 9 9 9 7 10 2 0 2 11 9 9 10 11 11 13 1 9 2
18 14 13 2 11 14 9 9 4 3 13 12 9 2 3 1 12 9 2
11 11 14 13 9 4 4 13 1 12 9 2
8 13 15 16 15 13 10 9 2
1 3
7 6 15 4 13 1 3 2
19 15 13 14 13 15 13 14 3 0 7 11 4 14 13 10 1 10 9 2
15 15 13 15 16 1 11 7 11 15 13 15 4 3 13 2
16 3 15 13 15 15 13 15 4 13 0 14 13 11 3 3 2
6 15 13 15 13 0 2
57 4 15 13 1 3 0 9 16 15 13 10 9 2 11 13 14 13 15 13 14 13 9 2 15 13 15 15 13 0 14 13 10 9 1 10 9 2 3 13 1 9 3 15 4 14 13 10 10 9 3 7 13 14 13 3 13 1
6 2 9 9 9 9 2
11 0 2 0 9 4 4 13 1 10 9 2
34 16 15 13 14 10 9 13 1 10 9 2 7 0 1 9 1 10 9 1 0 9 2 2 15 4 14 13 7 13 10 9 1 9 2
18 1 0 9 2 15 4 13 10 9 7 3 13 10 9 1 9 9 2
20 6 13 3 16 15 7 15 9 4 14 13 1 9 9 1 9 1 10 9 2
31 9 2 9 7 0 9 1 10 9 10 4 14 13 1 10 0 9 1 15 9 4 4 13 16 7 13 7 13 1 15 2
4 9 9 2 9
4 9 9 2 9
6 9 2 11 2 11 11
6 9 2 5 12 5 12
2 9 2
26 15 9 13 10 0 9 9 10 4 13 1 10 9 14 13 15 9 13 0 9 1 10 0 9 9 2
26 15 13 10 0 9 9 13 10 0 9 2 0 9 9 2 7 0 9 16 9 14 13 1 10 9 2
1 11
2 9 2
26 15 4 13 0 14 13 15 12 5 12 9 1 9 1 0 9 14 13 15 9 14 13 1 10 9 2
2 9 2
24 11 11 2 11 12 11 11 11 2 11 12 11 9 2 8 2 8 2 9 2 12 9 2 12
1 9
29 15 4 13 1 15 10 0 9 1 10 0 0 9 2 4 14 13 14 13 1 10 3 0 9 1 15 9 9 2
15 15 4 13 10 3 0 9 1 10 9 15 13 1 11 2
12 15 13 15 13 10 9 14 13 15 0 9 2
13 15 4 13 9 7 9 3 3 1 10 9 3 2
5 15 4 13 3 2
63 15 4 13 10 9 1 11 7 11 1 9 2 9 2 10 11 2 9 2 2 9 2 11 7 11 2 1 0 9 2 13 15 0 9 10 9 3 2 7 15 0 9 13 1 11 7 13 0 9 1 0 2 16 15 13 14 0 1 10 9 9 2 2
13 13 15 10 0 9 2 7 15 4 13 1 9 2
1 11
27 15 9 13 10 9 9 1 8 0 9 9 10 13 15 3 3 0 9 3 12 12 1 10 0 12 9 2
19 14 0 3 3 3 11 4 13 14 13 3 7 15 4 13 1 15 9 2
1 11
16 16 15 13 2 3 13 10 0 9 1 10 13 9 9 9 2
34 15 13 10 1 9 9 1 10 9 1 9 13 1 10 9 9 9 7 9 2 14 0 16 15 9 0 16 15 15 10 13 1 9 2
20 6 13 15 13 10 9 15 10 13 10 9 4 14 13 7 15 4 13 3 2
1 9
2 11 12
9 13 15 3 1 12 16 15 13 15
3 11 11 11
5 13 1 2 11 11
3 12 12 9
15 6 13 10 9 13 3 13 10 0 12 9 1 15 9 2
4 6 13 0 2
3 11 11 11
5 13 1 2 11 11
3 12 12 9
8 6 13 10 13 0 9 9 2
7 13 10 13 9 1 9 2
3 13 15 2
2 11 11
3 12 12 9
8 16 11 14 9 13 1 9 2
2 6 2
6 3 0 14 13 14 13
20 10 9 4 13 16 15 13 14 13 7 10 9 13 10 12 9 14 13 15 1
10 4 14 15 13 15 13 0 9 14 13
9 3 13 16 13 3 1 9 1 11
2 0 3
3 1 15 9
2 8 8
3 12 12 9
44 13 4 0 7 13 9 1 10 11 9 14 4 13 1 9 1 11 14 9 1 10 11 11 11 11 11 11 11 2 2 11 2 2 7 11 11 11 11 2 2 11 2 2 2
49 10 9 1 10 11 4 13 1 10 11 9 9 9 1 9 1 10 9 10 4 13 1 9 1 15 11 11 11 11 2 10 9 3 3 13 1 11 2 7 10 11 9 4 13 1 10 11 9 2
54 16 15 13 0 9 2 16 10 11 9 4 13 14 13 1 10 9 10 4 0 1 15 9 9 7 9 9 2 15 13 16 15 4 13 1 10 9 10 4 13 1 15 0 9 7 10 4 13 1 11 7 10 9 2
31 15 13 14 13 10 0 0 9 1 10 11 9 10 4 4 13 1 9 1 11 1 9 1 10 9 14 9 1 10 11 2
13 15 4 13 10 9 1 10 9 1 15 3 9 2
18 6 13 0 14 13 15 10 9 16 15 13 10 9 13 10 13 9 2
3 13 15 2
3 2 8 9
3 2 8 9
4 2 8 8 9
4 2 8 8 9
1 2
2 11 11
3 12 12 9
2 11 11
3 12 12 9
20 15 4 13 14 13 10 0 0 9 16 11 11 11 13 1 11 12 2 12 2
14 15 0 9 1 10 11 9 4 13 11 12 2 12 2
13 15 13 13 1 15 7 13 15 10 0 1 9 2
26 15 0 9 4 13 2 11 11 0 0 9 11 11 11 11 11 11 11 2 11 12 2 12 2 12 8
1 11
11 3 13 10 13 9 1 10 9 9 9 2
4 9 13 9 2
42 10 9 14 9 13 16 10 9 9 1 12 5 4 4 13 1 10 11 3 3 1 9 7 10 0 9 9 9 4 13 14 13 12 12 2 3 1 10 12 3 13 2
1 11
13 16 15 13 2 3 13 10 9 1 10 9 9 2
1 9
2 11 12
6 13 15 3 1 9 12
13 9 15 4 13 14 13 3 1 9 1 10 12 9
14 3 13 0 9 1 9 9 2 3 1 9 9 2 2
8 15 13 9 1 15 1 9 2
10 4 15 13 10 0 9 1 9 9 2
1 9
2 11 12
2 11 2
15 4 15 13 14 13 0 14 13 10 9 9 9 1 11 2
1 11
2 11 2
23 15 4 3 13 1 9 2 11 11 2 7 15 13 10 0 9 14 13 3 1 10 9 2
9 15 4 15 9 14 13 10 9 2
1 11
9 11 11 2 8 2 1 12 12 9
2 11 2
19 15 3 13 14 13 1 15 13 10 9 9 15 13 10 9 1 9 3 2
42 3 2 15 4 13 1 3 10 12 7 12 9 9 3 15 13 10 9 1 10 9 1 9 10 15 13 7 13 1 11 14 13 15 0 9 7 0 9 1 0 9 2
2 9 2
1 11
25 11 11 9 1 9 11 1 11 11 11 1 11 11 2 11 12 12 2 9 2 12 2 9 2 8
2 11 2
16 4 15 13 10 9 14 13 10 9 1 10 9 15 13 15 2
10 15 13 1 10 0 9 1 15 9 2
1 11
2 11 2
3 10 9 2
16 15 13 10 0 9 3 10 9 9 1 11 11 11 1 11 2
6 10 9 1 11 11 2
6 6 2 13 15 13 2
1 12
1 11
2 8 8
3 12 12 9
5 1 15 9 9 2
3 6 11 2
24 3 1 15 9 13 4 10 9 15 13 1 10 11 11 11 11 1 11 1 10 9 1 12 2
22 15 4 13 7 13 12 1 11 11 14 3 3 7 4 13 10 9 1 1 9 9 2
13 1 10 9 2 15 9 4 13 15 10 9 9 2
1 11
2 2 9
2 11 2
4 9 10 9 2
19 10 0 9 2 15 4 14 13 15 9 1 10 0 0 9 2 9 9 2
9 6 2 13 0 16 15 4 13 2
7 11 2 11 9 13 3 2
8 15 4 13 15 10 9 9 2
1 11
9 11 11 2 8 2 1 12 12 9
8 6 13 1 11 11 2 8 2
3 11 2 11
16 1 9 15 13 0 2 15 13 10 9 1 9 9 9 9 2
2 0 2
1 11
1 5
20 11 11 9 11 11 11 12 11 9 12 12 12 9 12 12 12 9 8 9 8
1 5
2 2 8
2 11 2
11 15 4 13 1 11 11 7 15 13 0 2
27 3 16 15 4 14 13 15 3 1 11 2 15 4 13 0 14 13 15 1 9 1 0 9 9 1 9 2
13 6 2 13 15 3 7 13 15 9 1 10 9 2
4 2 12 2 12
3 0 9 2
1 11
3 11 11 11
3 12 12 9
2 11 2
14 15 4 13 11 11 7 13 10 9 1 15 9 9 2
1 11
9 11 11 2 8 2 1 12 12 9
2 11 2
15 15 9 14 13 10 9 13 1 12 1 10 11 4 13 2
15 15 13 16 15 4 13 16 15 4 13 0 1 10 9 2
20 10 9 1 10 9 7 15 0 9 4 13 0 16 3 0 10 9 4 13 2
20 11 4 13 10 0 9 1 10 1 10 9 9 1 1 9 4 4 3 13 2
16 6 3 13 9 16 15 13 0 7 13 15 1 10 9 13 2
15 15 13 0 14 13 3 1 15 9 7 3 10 13 0 2
3 0 9 2
5 11 11 12 12 12
2 11 2
3 10 9 2
7 6 2 13 11 3 3 2
1 11
28 15 13 16 16 11 13 10 9 9 2 15 4 13 0 14 13 15 13 1 9 1 11 11 1 11 3 3 2
5 4 15 13 0 2
2 9 2
1 11
13 15 4 3 13 14 13 1 10 1 10 9 9 2
13 16 15 13 10 9 1 11 15 4 13 15 13 2
1 9
1 11
2 11 2
10 13 15 10 0 9 1 10 9 9 2
25 15 3 13 10 9 7 9 10 15 13 0 9 2 7 13 14 13 16 15 13 10 9 1 15 2
20 6 13 15 13 16 15 13 10 9 16 16 10 9 4 13 1 10 0 9 2
2 9 2
1 11
2 6 2
10 15 4 13 14 13 14 13 15 9 2
10 3 2 15 4 13 1 11 10 9 2
7 15 13 15 4 13 15 2
10 15 4 13 1 1 10 9 9 9 2
13 4 15 13 3 7 13 10 0 9 15 13 0 2
5 13 1 15 3 2
1 11
3 6 9 2
25 15 4 4 13 1 15 0 9 16 15 13 14 13 10 0 9 9 16 15 4 4 13 15 9 2
23 16 15 4 13 3 0 2 4 15 3 13 15 13 1 15 9 1 10 0 9 1 9 2
16 1 15 1 15 15 3 13 15 10 9 9 3 2 6 13 2
5 9 1 15 9 2
1 11
6 11 11 4 4 13 2
9 4 15 13 10 0 9 2 9 2
20 15 13 9 1 10 11 9 3 15 13 14 0 3 15 4 14 13 15 1 2
6 10 9 4 13 3 2
1 9
8 9 9 9 9 12 2 5 12
7 9 9 9 9 12 5 12
7 9 9 9 11 12 5 12
9 9 9 9 9 5 12 5 5 12
9 9 9 9 11 2 12 2 5 12
8 9 9 9 9 12 5 5 12
7 9 9 9 9 12 5 12
8 9 9 9 9 12 2 5 12
7 9 9 9 9 12 5 12
9 9 9 9 9 2 12 2 5 12
9 9 9 9 9 2 12 2 5 12
1 9
4 16 13 3 2
20 6 13 13 10 9 9 12 9 3 1 10 9 9 12 9 14 13 1 11 2
11 10 9 13 14 4 13 14 13 9 14 2
1 9
1 11
13 4 15 3 13 15 10 0 0 9 15 13 15 2
27 16 15 13 9 1 11 7 11 9 4 13 15 13 9 14 9 1 11 2 15 4 13 15 1 9 9 2
19 6 13 10 11 9 9 9 1 15 0 9 1 15 9 1 9 1 11 2
13 15 4 13 10 0 9 9 13 1 10 12 9 2
11 10 9 7 9 9 4 13 1 5 9 2
20 13 1 11 2 15 4 13 0 14 13 10 9 2 16 13 16 13 10 9 2
2 9 2
14 11 11 9 2 9 9 0 9 9 8 2 8 2 12
2 11 2
10 13 4 10 0 0 9 1 9 9 2
17 16 15 4 13 2 10 9 9 13 3 0 14 13 1 12 9 2
14 1 9 2 15 4 3 3 13 9 1 10 9 9 2
26 11 11 4 4 13 1 10 9 1 10 9 9 9 7 4 13 0 14 13 15 1 15 9 13 3 2
1 9
1 11
2 11 2
15 3 13 10 9 1 10 9 9 10 4 13 1 10 9 2
29 1 10 9 2 15 4 3 3 13 9 1 10 9 9 2 10 9 4 13 0 14 13 15 1 10 1 15 9 2
11 15 4 3 13 3 14 13 15 16 13 2
1 9
1 11
4 3 15 13 2
1 11
2 11 2
15 15 4 13 10 9 1 9 2 9 1 15 1 12 9 2
38 1 11 2 15 4 3 3 13 9 1 10 9 2 3 16 15 4 13 15 1 8 3 16 15 4 13 9 1 10 9 14 13 1 15 4 13 15 2
10 13 15 13 16 15 4 14 13 0 2
1 9
1 11
14 6 15 13 1 11 7 15 13 14 13 1 9 12 2
5 13 0 7 0 2
5 15 13 15 9 2
1 9
1 11
4 15 13 0 2
5 15 4 13 15 2
8 9 9 1 11 7 11 13 0
8 15 13 0 2 0 1 9 12
43 10 13 2 12 2 9 0 0 9 13 11 13 10 3 0 11 9 10 9 2 10 9 9 3 1 15 2 9 1 10 11 11 1 11 11 7 15 9 2 10 11 2 2
4 11 11 11 9
2 6 2
29 15 4 13 10 0 9 1 10 0 7 0 9 1 9 7 9 7 9 1 3 13 9 2 9 9 2 9 9 2
20 15 13 3 1 15 0 9 14 13 10 9 10 0 9 9 1 0 0 9 2
1 9
1 11
36 13 15 9 2 12 2 9 2 9 1 9 2 9 2 9 12 5 9 2 7 9 9 1 10 0 0 9 2 15 4 13 10 0 9 9 2
18 0 1 0 11 9 2 10 9 4 4 13 15 13 3 0 2 9 9
5 9 3 13 0 9
7 1 11 11 2 10 11 11
2 11 11
41 3 0 9 11 11 13 16 15 13 1 10 0 9 1 11 2 15 9 1 12 9 2 12 0 9 4 13 15 2 0 2 9 1 0 9 15 13 14 13 0 2
1 2
38 13 13 0 9 8 8 8 8 2 3 1 10 9 3 3 2 9 4 13 1 10 9 2 8 8 8 8 8 2 3 13 15 1 7 13 2 6 2
1 2
4 0 9 2 2
6 13 10 0 9 2 2
1 2
1 2
3 9 7 9
1 11
1 8
1 9
3 12 12 9
26 15 3 13 13 10 3 0 9 2 15 13 3 10 9 2 1 10 0 9 13 10 10 11 1 11 2
38 10 9 13 0 9 9 2 0 9 7 9 2 10 0 9 9 2 7 15 13 15 0 1 10 0 9 1 10 9 5 13 1 8 14 13 0 1 15
7 9 2 11 11 2 8 2
9 9 2 9 2 9 2 9 2 9
5 13 2 1 2 9
43 15 4 3 13 0 9 1 2 11 11 11 8 2 0 0 9 9 9 2 7 15 7 10 11 8 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 7 0 2
1 5
3 9 2 8
54 15 13 10 9 1 10 9 1 11 11 11 2 9 3 2 11 12 5 12 2 15 4 13 1 11 9 11 11 2 11 1 7 9 7 9 1 11 7 16 15 4 14 13 14 13 9 14 9 15 13 15 3 5 11
14 1 10 9 15 3 13 10 2 9 2 1 10 9 9
1 13
8 9 2 2 11 2 2 8 2
3 9 2 9
31 15 4 13 15 9 14 13 10 9 7 9 9 7 15 4 3 13 15 9 7 13 10 0 1 2 9 9 1 10 9 2
13 6 4 13 15 7 13 0 14 13 10 9 1 8
18 9 2 15 3 13 0 9 13 3 1 9 13 15 2 9 13 2 9
3 9 16 13
4 11 2 9 8
5 0 11 9 9 13
26 9 1 10 0 9 11 13 15 4 13 10 13 9 7 9 1 0 9 14 0 9 9 1 10 9 2
23 11 9 9 11 11 11 13 10 9 1 11 11 11 2 7 13 9 4 13 1 12 9 2
27 15 13 11 11 2 12 2 4 13 1 0 2 13 11 7 13 1 10 13 11 2 11 2 11 0 9 2
3 10 11 11
41 15 13 10 9 11 11 2 1 2 11 2 15 11 2 11 7 11 2 2 3 13 10 9 1 9 9 16 13 15 1 12 1 10 9 1 10 11 11 1 11 2
44 2 9 13 1 10 0 1 10 0 1 10 0 9 16 3 10 0 9 4 13 1 10 9 1 0 9 2 7 9 7 9 4 13 9 3 16 10 9 4 13 0 14 2 2
1 11
10 15 13 10 0 9 7 10 0 9 2
17 7 10 9 1 10 9 7 9 13 13 1 10 9 1 15 9 2
41 3 13 0 14 13 15 9 14 9 1 10 9 7 16 15 13 10 9 2 9 2 13 0 15 4 13 1 15 9 16 15 4 13 10 1 10 9 1 10 9 2
2 0 2
1 11
23 2 2 15 13 10 9 3 3 0 2 3 0 2 3 0 7 3 0 1 10 9 2 2
2 2 11
7 9 2 11 11 2 8 2
10 0 9 13 10 9 1 9 1 10 9
37 2 0 9 13 0 16 13 10 9 1 9 1 10 9 2 10 13 0 9 1 10 9 1 0 9 2 13 1 10 11 11 1 11 9 1 11 2
43 10 9 13 10 0 9 13 0 16 13 3 3 10 9 2 9 7 9 1 9 1 0 0 0 9 2 7 3 10 0 9 1 9 9 2 7 2 3 2 9 9 2 2
1 2
12 13 1 11 11 1 11 11 11 1 12 12 9
10 9 2 2 11 11 11 2 2 8 2
1 2
15 2 11 13 9 4 13 3 0 9 2 0 9 1 9 2
6 2 11 2 11 2 2
49 10 0 0 7 0 9 1 11 11 13 0 9 16 0 7 0 9 13 1 10 11 11 7 0 9 4 13 14 13 1 15 9 1 10 0 9 9 2 13 1 10 9 13 9 1 10 11 11 2
28 9 1 10 11 11 7 10 9 1 9 1 15 9 4 13 10 9 1 11 11 3 0 1 10 9 1 9 2
34 13 1 0 9 2 10 0 9 1 0 9 2 12 9 11 9 9 1 10 9 7 13 9 9 2 4 4 13 10 0 9 1 11 2
3 2 2 2
1 8
6 9 2 11 2 8 2
15 11 13 10 9 1 11 11 11 7 13 15 4 13 15 2
8 2 11 13 11 1 9 9 2
21 9 9 11 4 13 10 9 1 10 11 14 13 15 14 13 15 9 4 13 1 2
3 2 8 2
5 2 11 11 11 2
19 13 10 9 7 9 9 15 13 2 3 15 13 15 2 3 1 12 0 9
3 2 8 2
3 2 9 2
29 10 11 13 14 0 1 10 9 1 10 9 2 7 9 13 1 10 9 4 14 3 13 10 11 14 9 7 9 2
16 6 13 16 7 10 9 9 7 9 1 10 9 4 4 13 2
33 16 15 4 14 13 14 13 0 9 1 10 9 7 13 14 13 0 1 10 11 14 13 10 9 9 2 6 13 15 3 13 9 2
1 8
3 2 8 2
31 16 9 13 1 1 10 0 9 1 11 2 1 10 0 9 2 2 11 11 13 0 11 11 11 7 0 0 9 1 11 2
17 10 9 1 10 9 1 10 3 0 9 9 1 11 13 11 11 2
29 11 4 13 10 0 9 16 13 11 11 1 10 9 7 11 4 13 16 1 15 9 11 4 13 10 0 0 9 2
4 11 2 11 11
19 11 11 11 11 11 13 9 1 0 11 11 11 1 10 0 9 1 11 2
18 11 13 1 11 1 10 0 11 2 11 11 11 2 11 2 9 9 2
27 3 11 11 4 13 10 9 10 4 3 3 13 13 15 0 9 2 7 4 3 13 13 10 9 1 9 2
2 11 2
1 2
11 13 1 11 11 1 11 11 1 12 12 9
6 9 2 11 2 8 2
3 9 2 9
10 15 13 10 9 14 13 1 15 9 2
13 15 13 0 11 9 2 3 15 13 0 1 9 2
15 15 13 13 9 7 9 3 14 13 1 15 9 7 9 2
13 15 13 10 9 7 13 14 13 15 1 15 9 2
14 3 15 13 10 0 9 9 7 13 15 9 1 15 2
15 1 1 10 9 1 10 9 1 15 14 13 10 9 9 2
7 15 13 1 12 9 9 2
7 15 3 13 3 12 9 2
14 15 9 7 15 4 13 16 15 14 13 7 13 15 9
5 8 15 9 1 9
19 8 16 13 0 2 15 13 10 0 9 9 2 13 7 13 7 13 15 9
9 5 13 1 8 2 0 9 9 5
11 8 2 10 9 12 9 9 1 10 9 2
10 5 3 12 9 2 12 0 9 2 5
11 13 0 9 3 2 13 1 10 9 3 2
1 12
19 13 9 0 9 0 9 13 1 9 7 9 9 2 9 7 9 14 9 2
20 9 2 9 2 9 2 9 2 9 2 9 2 15 13 15 2 15 13 15 2
14 9 13 14 13 10 0 0 0 9 1 9 7 9 2
8 15 13 3 3 13 7 0 2
6 9 9 9 7 9 2
12 15 4 13 14 13 15 0 9 1 10 9 2
35 16 15 13 10 9 9 7 13 10 0 9 15 13 1 9 2 9 2 7 9 9 7 13 0 16 13 15 9 2 6 13 15 10 9 2
1 12
17 15 13 10 0 9 9 7 0 9 9 0 14 13 1 15 9 2
5 10 0 9 9 2
16 10 9 1 7 1 5 12 10 0 12 5 1 10 0 9 2
23 15 13 2 11 2 11 2 11 2 11 14 11 2 11 11 2 7 0 9 2 9 9 2
14 8 8 8 11 11 8 12 12 11 11 11 2 11 12
4 11 14 0 9
24 11 11 2 10 13 9 1 0 9 1 11 2 3 13 10 9 1 11 2 12 1 11 11 2
7 15 4 3 13 1 11 2
9 15 9 3 13 9 7 0 9 2
16 15 4 13 1 12 1 10 13 9 2 9 9 1 0 9 2
12 15 9 4 13 7 13 1 11 11 1 12 2
33 2 11 4 13 10 9 9 1 9 7 9 2 3 13 0 0 9 1 10 0 9 2 2 13 11 11 11 2 9 1 10 9 2
20 1 10 9 1 2 11 14 0 9 2 2 10 13 14 13 3 13 7 0 2
8 10 13 0 2 10 13 0 2
40 1 11 14 9 2 10 9 4 13 0 9 2 10 9 4 13 10 9 1 12 0 9 2 10 9 9 4 13 9 2 7 11 11 4 13 12 13 0 9 2
18 2 2 14 13 1 11 14 9 13 16 13 10 13 9 1 9 2 2
15 2 10 11 1 11 1 11 11 2 11 11 11 2 12 2
3 2 8 2
4 9 1 11 11
31 11 11 11 2 10 9 1 10 11 0 9 9 2 13 11 16 9 9 11 4 13 14 13 10 1 15 9 1 9 9 2
4 2 11 11 2
16 15 13 16 10 9 1 11 7 11 4 3 13 1 10 9 2
26 11 13 12 5 12 2 15 13 1 11 2 11 11 2 11 7 11 2 7 11 4 13 15 0 9 2
18 11 4 3 13 10 9 14 13 11 11 13 11 2 15 0 9 2 2
3 0 3 2
21 7 15 13 16 11 4 14 13 15 9 1 10 9 1 10 9 16 11 11 13 2
30 2 16 15 4 14 13 9 0 14 13 9 2 11 7 10 11 11 4 3 13 0 9 14 13 8 7 15 9 2 2
19 6 11 2 16 15 4 13 15 1 9 1 0 9 1 10 9 1 12 2
30 15 4 13 0 14 13 16 7 3 11 4 3 13 10 11 9 2 15 4 13 10 0 9 7 13 14 13 10 9 2
2 11 2
1 2
11 13 1 11 11 1 11 11 1 12 12 9
8 9 2 2 11 2 2 8 2
2 6 3
18 11 11 13 10 11 9 1 9 15 4 13 9 1 9 10 13 15 2
19 15 4 13 1 9 16 15 13 15 4 13 0 1 9 13 1 9 9 2
31 15 4 13 10 9 13 1 9 1 9 2 8 2 7 10 9 13 11 11 4 3 13 1 10 9 1 9 9 1 11 2
26 15 4 13 14 13 15 1 14 13 10 9 1 10 10 9 2 10 9 3 9 4 13 9 7 9 2
35 15 4 13 0 16 10 9 1 11 15 13 10 9 4 13 3 10 0 9 1 10 9 7 10 9 1 10 9 9 1 10 11 11 9 2
30 11 11 13 3 10 0 9 14 13 9 1 9 2 7 13 14 13 3 10 9 16 15 13 14 13 9 1 15 9 2
23 15 4 13 9 15 13 1 9 1 15 0 9 2 3 3 1 1 10 2 9 2 9 2
25 15 13 0 1 0 14 13 9 1 10 9 7 13 10 9 1 11 11 2 3 13 15 10 9 2
8 3 2 13 14 13 15 3 2
2 0 9
3 11 11 8
7 11 11 4 13 10 9 2
21 1 12 9 2 15 13 10 9 16 9 4 13 15 10 9 1 10 2 9 2 2
39 12 0 9 13 3 7 13 16 2 2 16 15 0 9 15 13 0 9 4 13 1 10 9 3 10 9 13 3 7 13 15 2 15 4 13 10 9 2 2
15 2 6 2 2 11 13 2 2 15 4 13 10 9 2 2
6 10 9 13 15 9 2
24 2 16 10 9 9 13 12 9 13 1 10 9 2 13 9 0 2 15 4 13 10 9 2 2
22 2 15 13 0 14 2 2 13 11 2 2 15 13 15 15 4 13 10 0 9 2 2
12 10 9 13 0 2 9 1 10 0 9 13 2
25 2 15 2 2 13 11 2 2 13 14 15 8 9 3 15 4 13 15 10 9 1 10 9 2 2
11 3 2 10 9 1 10 9 13 15 9 2
29 1 10 0 9 2 15 13 2 2 16 10 9 13 11 11 4 13 1 1 10 9 2 10 4 13 10 9 2 2
7 2 0 2 2 11 13 2
3 2 0 2
13 7 4 15 13 15 3 15 4 13 10 9 2 2
28 2 6 2 2 13 10 9 2 2 16 15 4 14 13 10 9 2 7 15 3 4 14 13 10 0 9 2 2
3 2 8 2
3 9 1 8
3 2 8 2
28 15 13 16 10 11 11 11 2 11 4 13 10 2 9 9 2 13 1 10 11 1 11 2 7 3 3 2 2
33 2 15 0 0 9 9 13 10 0 9 10 4 13 10 9 1 10 12 2 9 9 1 10 11 7 10 11 2 2 11 13 8 2
36 2 15 9 13 13 0 9 14 13 2 13 2 9 13 2 7 13 10 11 2 11 9 1 10 9 1 10 9 7 10 9 1 15 9 2 2
23 0 9 14 13 1 10 0 9 2 11 14 9 4 13 3 0 14 13 10 9 1 15 2
8 10 9 4 13 3 0 3 2
22 10 11 11 11 2 11 2 4 3 4 13 1 12 9 9 2 11 11 7 11 11 2
28 10 1 10 9 13 3 0 1 10 0 9 1 10 9 9 2 7 10 13 3 0 1 10 9 9 13 11 2
28 15 13 14 13 11 14 13 1 11 14 9 1 9 9 2 7 13 0 16 10 11 11 4 13 1 10 9 2
48 2 15 13 3 0 16 10 11 11 7 10 0 0 9 9 9 13 10 9 14 13 10 0 9 16 13 11 13 15 9 1 10 0 9 1 9 9 2 2 13 11 11 2 11 9 7 9 2
26 1 15 9 1 10 2 11 2 11 2 9 2 15 13 16 9 9 4 13 10 9 3 16 15 13 2
2 11 2
1 2
11 13 1 11 11 1 11 11 1 12 12 9
3 2 8 2
3 2 8 2
43 11 9 4 13 1 10 9 1 0 2 0 2 9 9 9 7 10 0 0 0 2 9 9 10 9 4 13 1 0 1 10 9 2 11 7 10 11 4 13 10 11 11 2
35 0 9 7 0 9 13 1 0 9 1 10 11 4 4 13 1 0 9 3 0 1 10 11 2 9 11 11 2 10 3 0 9 3 13 2
30 15 13 16 16 11 4 13 3 1 10 9 9 2 16 1 10 9 15 4 13 14 13 3 0 16 11 4 3 13 2
42 16 10 0 9 13 3 3 0 2 15 4 13 0 14 13 1 10 3 0 9 1 15 9 9 2 16 15 4 3 3 13 0 1 10 9 7 13 10 11 3 3 2
49 2 11 4 13 9 1 10 9 9 9 13 1 9 9 0 9 9 1 10 0 0 9 1 0 9 2 2 13 10 9 2 13 1 11 9 11 11 7 10 11 14 0 9 9 2 9 11 11 2
43 2 11 3 13 14 13 10 0 12 2 0 2 9 2 9 9 9 13 1 13 9 1 10 9 9 0 9 7 0 9 9 1 0 9 1 10 11 2 2 10 9 13 2
25 11 4 13 16 13 10 0 9 14 13 10 0 9 2 16 9 9 13 10 9 3 0 1 12 2
35 10 0 9 9 4 13 3 1 15 9 2 1 10 9 16 10 9 7 9 4 13 3 1 12 0 9 10 7 13 1 1 9 3 3 2
18 13 10 9 4 3 13 0 9 2 13 0 9 16 11 13 10 9 2
1 2
11 13 1 11 11 1 11 11 1 12 12 9
3 11 7 11
1 9
3 12 12 9
2 0 9
4 13 1 10 9
2 11 5
1 2
18 15 4 3 13 10 9 9 1 16 15 13 14 13 15 9 1 11 2
3 2 11 11
13 15 13 10 9 13 1 15 7 15 13 3 0 2
27 7 15 13 14 0 14 13 10 9 1 10 9 2 2 3 0 1 10 9 2 7 0 1 10 9 2 2
3 2 11 11
1 2
7 11 11 13 10 0 9 2
7 13 9 3 3 10 9 2
3 2 11 11
1 2
7 2 1 10 9 2 13 2
25 16 15 13 10 0 9 2 15 4 13 0 2 16 15 13 10 0 9 2 15 4 13 10 9 2
2 2 11
1 2
7 15 4 13 1 10 9 2
8 15 4 4 13 1 10 9 2
3 2 11 11
1 2
10 15 9 13 10 0 9 1 15 9 2
9 3 3 7 3 15 13 14 13 2
3 2 11 11
1 2
13 15 4 3 13 10 9 3 14 13 15 9 1 2
4 2 11 11 11
1 2
22 3 0 9 13 1 10 0 9 10 12 0 9 9 2 9 2 9 2 9 7 9 2
3 2 11 11
1 2
19 9 4 14 13 15 9 2 7 15 4 13 15 10 3 0 9 1 9 2
3 2 11 11
1 2
13 16 15 13 12 2 15 13 15 9 13 13 1 2
3 2 11 11
1 2
15 9 4 13 10 0 9 16 15 13 10 0 3 1 9 2
4 2 11 11 11
1 2
6 15 4 14 13 0 2
8 15 4 14 13 9 1 9 2
8 3 15 13 9 1 15 9 2
3 2 11 11
1 2
17 4 14 13 16 13 9 2 16 15 13 0 2 15 4 13 15 2
3 2 11 11
1 2
25 3 15 13 0 16 9 13 1 12 2 7 9 0 13 14 13 1 2 13 1 2 7 13 1 2
3 2 11 11
1 2
21 1 10 9 10 9 13 0 3 14 13 15 9 2 15 13 3 0 14 13 3 2
3 2 11 11
1 5
4 4 15 13 2
4 0 1 9 2
8 11 11 13 10 0 9 9 3
1 9
3 12 12 9
7 10 9 4 13 1 11 2
1 11
1 11
6 0 9 7 0 9 2
1 0
3 0 9 2
2 0 9
5 15 13 10 11 2
7 15 13 10 9 1 11 6
9 4 9 13 10 0 9 1 11 2
4 14 15 6 2
10 4 9 13 1 10 0 9 1 11 2
4 14 15 6 2
14 10 0 9 1 15 4 9 13 10 15 0 9 5 2
1 5
9 15 13 10 0 9 9 1 11 2
8 9 2 9 2 9 9 2 9
13 4 15 13 10 0 9 9 1 11 11 12 11 2
4 10 9 9 2
2 6 2
5 3 9 1 11 2
6 11 13 10 0 9 2
8 6 2 11 13 14 1 9 2
1 6
8 10 4 15 13 9 7 9 2
11 15 13 9 2 13 2 13 2 7 13 2
1 9
1 9
11 3 0 4 15 13 14 13 11 11 11 2
6 4 14 13 10 9 3
5 13 15 1 9 3
3 9 2 8
1 11
8 15 13 9 11 11 2 13 2
1 8
2 15 9
1 8
15 3 0 4 15 13 14 13 10 11 11 9 1 15 9 2
17 3 1 11 15 13 15 13 6 5 12 7 5 12 1 10 9 2
8 11 7 11 1 10 11 9 2
25 10 9 9 4 15 13 13 3 0 1 11 7 11 7 0 1 10 11 9 1 11 11 7 11 2
8 3 14 13 9 9 1 11 2
11 10 0 9 10 15 13 1 7 15 9 2
6 11 11 2 11 11 2
8 3 13 11 11 11 1 11 2
10 4 15 13 15 13 10 11 1 11 2
9 6 15 4 13 3 3 12 11 2
17 6 2 7 15 4 13 10 11 13 1 10 9 1 11 2 11 2
17 4 15 13 10 2 13 15 9 2 9 14 13 9 0 14 9 2
21 15 4 13 15 11 9 7 9 2 16 15 13 15 3 6 15 4 13 10 11 2
13 16 13 0 9 2 15 3 4 9 13 1 11 2
18 6 2 15 13 10 9 1 9 10 15 13 1 9 2 9 2 8 2
8 6 15 13 10 11 1 15 5
5 13 11 11 0 2
9 10 11 11 15 13 13 3 0 2
14 15 13 10 9 2 7 15 13 15 9 10 10 9 2
13 15 13 1 15 0 3 15 4 13 15 9 9 2
6 9 1 11 1 11 2
5 3 15 13 0 2
14 15 4 7 4 14 13 9 2 13 1 0 9 9 2
18 1 10 9 9 9 2 15 4 3 13 9 2 13 9 1 10 9 2
15 11 13 15 0 14 13 15 9 9 7 3 13 15 13 2
5 9 1 15 9 2
25 1 1 10 0 9 2 9 4 3 13 1 10 0 9 1 9 1 9 2 9 2 9 2 8 2
5 0 9 9 5 2
25 15 4 13 1 9 1 8 8 7 8 7 9 10 13 14 3 0 7 13 10 9 1 0 9 2
11 6 13 15 9 1 9 7 9 14 13 2
3 13 15 5
1 8
12 3 4 15 13 9 7 9 1 10 9 9 2
7 13 12 1 15 13 9 2
4 13 10 9 2
2 13 2
14 13 1 9 2 3 13 10 9 7 13 10 9 1 15
11 15 13 10 9 1 0 9 7 9 9 2
12 4 15 13 9 2 9 7 9 1 15 9 2
7 1 10 9 2 9 2 5
7 3 13 9 7 3 0 9
24 1 15 9 15 13 9 7 9 3 15 13 10 0 9 1 10 0 9 1 9 7 10 9 2
13 4 9 13 10 9 9 3 16 15 4 13 1 2
13 4 9 13 10 9 9 3 16 15 4 13 1 2
12 6 15 13 14 13 15 2 15 13 10 0 9
12 6 2 15 10 13 0 9 9 2 3 1 9
2 6 2
10 11 14 11 0 0 9 1 11 11 2
20 13 11 14 11 1 12 11 9 1 11 11 3 10 0 0 9 1 10 9 2
21 16 10 1 10 9 9 15 4 13 13 3 7 15 4 13 1 11 16 15 13 0
1 6
6 9 7 9 1 11 2
29 15 13 1 12 5 7 13 1 10 0 9 14 13 15 9 3 1 9 3 15 13 9 7 15 13 10 9 9 2
10 15 13 0 16 15 13 10 0 0 2
8 10 0 9 4 3 4 13 2
2 11 11
5 11 10 0 9 2
26 1 10 9 2 3 1 11 13 15 11 2 2 3 0 0 9 2 9 13 15 7 15 13 10 9 2
5 9 1 9 2 8
10 15 4 3 13 15 1 10 9 9 2
10 15 4 3 3 13 1 10 9 3 2
13 13 9 15 13 1 10 9 10 13 1 10 9 2
2 9 9
2 9 9
2 9 9
2 9 9
15 9 1 10 9 2 9 1 0 9 9 9 1 9 2 2
4 10 1 15 5
3 9 9 2
7 10 9 4 15 13 1 2
11 15 13 15 9 9 1 10 9 1 0 2
13 3 13 10 9 13 14 13 10 9 1 10 9 2
7 15 13 1 15 3 3 2
12 16 3 0 9 4 3 3 13 1 10 9 2
6 9 13 14 13 0 2
6 15 4 3 13 3 2
19 6 2 15 4 14 13 9 3 16 15 13 10 9 15 2 11 2 13 2
8 15 4 15 13 1 11 11 2
5 15 13 11 11 2
19 15 9 13 0 2 9 7 15 3 13 10 0 0 9 13 3 1 9 2
12 15 3 13 15 9 3 0 1 0 0 9 2
8 7 15 13 1 10 0 9 2
11 15 13 1 1 15 9 14 13 11 11 2
1 0
14 15 13 10 9 1 0 7 0 9 7 0 9 2 2
31 15 4 13 14 13 10 0 9 2 13 10 9 1 9 2 2 15 13 10 3 0 9 9 2 9 2 9 2 9 2 2
11 7 13 12 0 9 10 13 10 9 0 2
9 3 4 9 13 15 10 9 13 2
1 9
16 16 15 13 10 9 1 11 4 9 0 13 15 1 1 15 2
10 15 13 5 12 9 1 1 15 3 2
43 6 15 4 14 13 0 14 10 11 4 14 13 9 1 10 9 3 10 9 4 13 3 16 13 15 7 10 9 1 9 13 14 13 15 9 7 2 7 15 9 1 10 9
9 4 9 3 13 1 11 11 11 2
19 15 4 13 13 10 9 1 11 7 13 15 13 14 13 1 10 15 9 2
17 4 13 16 9 13 10 0 9 16 3 0 15 13 1 9 7 9
14 15 4 14 3 7 15 13 10 9 1 9 15 13 2
12 11 4 13 1 15 13 10 9 1 15 9 2
6 0 9 9 1 11 2
13 15 13 10 0 9 9 15 4 13 1 11 11 2
8 15 13 9 0 7 0 0 2
8 11 11 13 10 0 9 9 2
27 15 13 15 1 15 9 7 3 13 9 1 10 0 9 1 10 9 9 3 14 13 3 0 10 9 13 2
10 13 15 10 9 7 13 15 10 9 2
1 8
7 15 13 2 0 2 9 2
32 15 4 4 13 1 10 11 11 11 12 15 4 3 13 10 11 8 9 9 2 15 4 13 15 4 13 10 0 9 1 9 2
12 15 13 9 3 0 7 1 10 9 1 9 2
17 3 15 4 13 2 13 15 0 16 10 0 10 9 13 10 0 2
1 9
4 0 7 0 2
4 11 13 14 0
7 11 9 1 11 2 11 2
9 15 4 13 11 9 0 12 9 2
11 15 4 4 13 13 11 9 9 0 9 2
9 4 15 13 14 13 9 1 11 2
8 15 13 10 9 1 15 9 2
13 3 4 13 14 13 9 16 15 13 10 9 2 2
11 15 3 13 15 13 10 9 9 1 9 2
2 6 2
8 6 2 15 4 13 9 9 2
7 12 9 0 9 3 3 2
13 6 15 13 11 11 14 2 11 11 2 11 11 2
17 7 15 9 13 3 0 1 10 1 15 2 7 15 13 3 3 2
12 15 13 3 1 10 9 7 3 1 10 9 2
3 1 15 2
14 11 2 11 11 2 11 11 2 0 9 2 0 9 2
6 11 13 10 0 9 2
7 11 14 11 11 11 2 5
13 11 2 4 15 13 15 15 4 13 14 13 1 2
8 7 4 15 13 1 0 9 2
5 15 13 3 0 2
12 11 1 11 2 13 15 3 0 3 14 13 2
1 6
3 14 0 3
5 11 11 2 7 6
3 3 11 2
18 11 11 13 3 0 13 1 15 0 9 2 16 10 9 1 15 13 2
8 6 2 15 4 3 13 11 2
7 15 4 13 15 1 10 9
10 13 1 11 1 10 0 9 1 11 2
16 4 15 4 13 14 13 9 0 9 1 15 13 9 1 11 2
16 1 15 9 9 7 4 15 13 14 13 15 1 15 13 9 2
2 6 2
6 15 4 14 13 15 13
9 15 4 13 15 1 2 9 9 2
22 6 15 4 13 15 9 0 9 2 7 9 1 15 9 16 15 13 3 10 0 9 5
6 13 1 11 2 11 2
15 16 15 13 1 10 2 0 2 9 16 9 9 1 9 2
13 13 16 15 13 10 12 9 7 15 13 10 9 2
26 4 15 13 0 14 13 3 1 9 1 10 9 9 1 10 9 14 13 10 11 14 9 1 9 9 2
5 10 9 4 13 2
2 13 15
8 15 4 13 0 14 10 9 2
9 9 4 13 15 10 9 15 13 2
13 15 4 15 13 10 9 10 13 1 15 9 9 2
7 7 3 4 15 13 15 2
4 9 9 9 2
3 7 9 9
9 13 15 1 10 0 9 9 9 2
1 9
3 9 3 2
10 0 13 15 13 10 9 1 10 9 2
1 8
3 9 9 2
24 13 10 9 7 13 9 9 9 7 13 15 1 10 9 9 2 7 13 1 9 9 9 2 2
19 1 1 11 2 11 11 2 7 11 2 9 2 10 13 10 0 7 3 2
9 15 13 11 11 1 1 10 10 2
8 15 13 3 0 14 13 3 2
17 10 0 11 11 4 13 0 2 16 15 4 14 13 1 15 3 2
5 9 1 10 0 2
15 1 10 12 2 15 13 10 9 2 9 1 11 7 11 2
14 11 13 10 9 1 10 2 1 9 1 9 7 9 2
21 4 9 13 9 9 3 13 3 16 15 4 13 1 1 10 9 10 4 13 1 2
3 15 13 2
6 15 13 10 11 11 2
4 13 1 10 9
23 16 10 9 4 3 13 1 2 10 9 9 4 14 13 9 2 3 15 4 14 13 15 9
30 0 9 13 9 7 9 3 2 10 13 10 9 14 13 1 9 9 2 7 3 13 10 9 9 14 13 9 1 9 2
10 15 13 10 0 9 1 10 0 9 2
13 2 1 11 2 9 4 13 2 13 2 7 13 2
9 13 13 3 15 13 10 9 2 2
5 10 9 1 11 2
12 3 13 10 9 10 13 10 9 1 9 9 2
10 3 0 9 13 7 3 10 13 14 2
11 15 4 13 15 0 16 13 10 0 9 2
6 10 9 1 9 2 8
5 0 9 9 2 8
3 0 9 2
6 10 0 9 2 0 2
9 10 0 9 9 4 15 13 2 2
23 15 4 13 1 10 9 10 13 3 0 9 1 10 9 7 9 2 7 0 9 9 2 9
25 15 4 13 16 13 10 0 9 9 1 11 11 2 3 6 13 10 9 2 8 2 15 4 13 2
12 3 3 0 4 0 9 9 13 1 11 11 2
15 2 7 15 4 13 15 9 7 9 1 10 9 2 11 2
6 13 10 9 1 11 11
6 15 13 0 9 9 2
24 15 13 10 0 9 16 13 10 9 13 10 9 9 1 10 0 9 1 10 0 7 0 9 2
18 10 0 9 2 9 2 13 14 13 1 10 9 7 13 1 10 9 2
42 9 13 0 2 7 0 2 3 15 13 10 9 1 15 2 15 4 13 10 9 13 2 3 10 9 2 7 3 13 3 10 9 1 9 0 9 2 13 15 13 0 2
3 13 11 2
3 9 11 2
7 15 13 10 9 1 11 2
13 4 9 13 15 3 15 15 13 7 15 13 9 2
8 15 4 14 13 10 9 1 15
24 3 10 11 13 1 11 1 10 9 1 11 11 10 11 11 13 1 9 1 10 11 11 11 2
15 15 13 10 11 1 1 10 9 2 11 2 7 13 9 2
8 13 15 15 15 4 13 1 2
24 15 13 14 13 1 10 0 11 11 2 12 5 12 2 7 10 11 11 2 12 5 12 2 2
9 4 10 9 3 13 10 9 9 2
7 7 3 9 0 7 9 2
10 15 13 15 4 13 1 10 9 9 2
15 6 2 3 15 4 14 13 10 9 9 2 15 13 0 2
14 3 2 15 3 4 14 13 16 15 13 14 13 12 2
28 10 9 9 4 13 10 9 9 10 13 10 9 9 1 10 0 9 11 1 3 3 12 5 12 9 10 9 2
20 4 14 13 14 13 10 9 9 3 10 9 2 0 9 13 0 1 9 9 2
8 9 0 0 9 9 11 11 2
10 13 1 10 9 9 14 13 15 9 2
11 10 9 4 13 0 7 3 9 3 0 2
17 15 4 13 14 13 12 1 10 3 0 3 0 9 3 2 9 2
23 6 7 10 0 10 0 2 15 4 13 14 13 9 3 2 3 2 15 4 13 0 2 9
19 3 14 13 3 10 9 1 9 2 10 9 7 13 10 9 1 11 11 2
8 0 2 0 9 2 9 3 2
7 15 13 9 1 0 9 2
2 13 8
9 15 9 9 0 9 4 14 13 2
37 1 10 0 0 9 15 4 4 13 7 4 14 13 7 15 4 13 3 15 0 9 4 14 13 7 15 13 3 1 15 9 2 15 4 15 13 2
49 3 13 1 15 7 13 14 13 15 9 7 13 10 0 9 1 10 0 9 7 13 15 1 10 9 7 16 15 13 10 0 9 13 9 1 15 9 7 9 7 16 15 4 14 13 13 15 1 9
6 13 15 1 10 9 2
6 3 13 15 1 10 9
20 3 0 4 15 13 16 15 14 13 15 7 12 9 1 11 14 9 1 9 2
29 6 2 15 4 13 14 13 15 7 15 0 9 7 15 9 9 7 10 9 15 3 13 1 1 9 1 15 9 2
29 15 3 13 14 13 1 11 14 1 15 9 7 15 4 3 13 3 0 15 4 13 16 10 12 1 15 14 13 3
14 13 10 9 10 9 1 9 15 13 7 3 15 13 2
11 3 13 1 5 12 1 9 3 3 15 2
7 7 0 16 15 13 9 2
15 15 13 9 1 11 11 9 1 0 9 7 0 9 9 2
16 15 13 9 1 9 1 11 11 1 0 9 7 0 9 9 2
15 15 13 12 0 9 12 13 1 12 7 10 13 1 12 2
16 0 9 2 9 9 2 0 2 0 2 7 0 13 10 9 2
11 3 13 10 0 9 1 0 9 1 11 11
1 8
16 6 16 15 4 14 13 15 9 2 15 13 11 11 1 0 9
8 15 13 0 7 15 13 0 2
11 11 11 13 3 0 9 7 15 13 3 0
2 13 8
9 3 0 9 1 10 9 1 11 2
4 13 1 15 2
8 9 13 9 2 9 13 9 2
16 16 15 13 0 9 2 12 2 1 13 1 10 12 1 11 2
10 10 0 9 13 0 1 10 11 9 2
8 12 0 9 1 10 9 1 11
15 16 11 2 11 13 2 15 13 3 12 1 10 0 9 2
40 13 15 3 16 15 13 10 2 0 2 9 1 10 9 1 11 15 13 1 1 13 14 13 10 0 9 1 11 1 9 2 7 15 13 15 1 0 0 9 2
9 10 9 4 14 13 0 3 3 5
6 13 9 13 0 9 2
11 15 13 10 11 7 13 15 13 1 11 2
8 15 4 13 0 9 1 15 6
23 10 9 1 10 11 13 15 4 14 13 3 0 2 15 4 13 14 13 15 13 1 11 2
24 6 16 15 13 0 2 15 13 15 13 10 9 1 11 11 2 11 11 11 11 7 11 11 2
7 15 13 15 4 13 0 2
15 15 13 15 4 13 10 0 9 1 10 2 9 2 9 2
2 2 11
9 7 15 13 9 3 0 1 15 2
15 15 4 13 0 9 1 15 10 13 1 10 11 7 11 2
11 9 14 9 9 2 3 4 15 13 12 2
21 15 4 13 1 10 9 1 11 3 2 7 15 13 14 13 10 0 2 0 9 2
13 15 4 13 7 13 2 7 4 14 13 12 3 2
10 15 4 13 10 0 2 0 0 9 2
25 15 3 13 14 13 3 0 2 10 0 12 15 13 13 15 0 1 9 0 1 0 2 0 9 2
15 15 4 13 1 1 12 5 12 1 15 16 15 13 14 2
5 13 1 10 11 9
4 1 10 11 9
6 15 13 10 0 0 9
5 3 13 10 9 2
1 8
24 15 13 10 11 9 2 12 9 2 2 11 11 11 0 9 2 3 4 15 13 15 16 13 2
24 15 13 10 11 9 2 12 9 2 2 11 11 11 0 9 2 3 4 15 13 15 16 13 2
17 15 13 14 2 15 13 10 0 9 1 2 9 2 1 0 9 2
22 15 13 1 1 10 9 10 13 10 9 16 15 13 0 14 4 13 1 10 9 9 2
23 3 15 13 10 9 14 13 13 10 9 4 13 1 10 9 1 10 9 9 2 10 9 2
19 10 15 4 13 13 13 10 9 2 0 9 2 7 13 15 3 1 9 2
7 15 13 10 11 11 9 2
45 3 11 4 13 14 13 10 9 9 4 15 13 1 10 9 1 10 9 15 13 15 9 7 15 13 15 9 16 15 9 13 15 13 15 13 15 9 2 7 15 4 14 13 9 2
27 15 13 15 13 1 10 0 9 2 7 3 2 15 13 10 9 1 10 9 2 7 16 15 14 13 15 2
26 6 2 3 2 15 4 13 10 9 1 10 0 9 2 13 1 11 2 1 10 13 3 1 11 9 2
10 4 15 13 15 13 0 1 10 9 2
6 6 2 15 13 10 2
3 10 0 2
14 11 11 4 13 14 4 13 1 11 2 3 1 11 2
18 13 15 10 0 9 14 13 10 9 2 9 9 1 1 11 11 11 2
32 3 15 13 1 11 11 11 7 15 13 14 13 16 15 13 10 0 9 14 13 10 9 2 9 9 1 0 1 11 11 14 6
7 0 9 9 2 9 2 9
12 15 13 1 11 7 15 13 11 14 9 9 2
4 15 13 0 2
20 10 1 10 0 2 0 9 13 0 9 2 9 2 13 15 14 13 15 1 2
46 10 9 9 1 11 3 3 3 16 11 11 13 10 0 0 9 9 1 10 9 15 13 1 11 1 10 0 9 13 10 9 9 7 3 13 15 15 4 13 3 3 14 13 10 9 9
8 0 9 9 1 10 11 9 2
27 10 13 10 0 9 9 1 10 11 0 9 6 1 9 11 11 11 14 11 11 10 9 4 13 10 3 2
3 11 11 2
10 9 9 13 0 7 10 9 13 0 2
3 11 14 2
3 13 15 9
2 9 2
6 4 12 13 10 9 2
14 11 14 13 10 0 9 9 10 13 1 12 9 3 2
6 15 13 3 12 9 2
1 8
13 10 0 9 1 10 0 11 14 13 11 14 11 2
1 8
16 13 15 11 7 11 13 1 10 0 9 1 11 11 1 11 2
1 8
17 1 1 10 0 9 13 10 9 1 9 9 16 15 13 1 9 2
8 3 10 0 9 4 13 0 2
1 8
16 15 9 13 13 1 0 9 1 12 9 7 4 14 13 9 2
5 15 4 15 13 2
13 15 4 13 0 0 9 7 15 4 14 13 9 2
5 15 4 15 13 2
5 4 15 13 0 2
12 13 10 9 4 13 10 0 9 1 10 0 9
3 3 0 2
9 6 13 15 9 1 10 9 3 2
65 3 16 14 13 2 16 15 4 3 13 3 7 4 13 15 14 13 3 3 2 15 4 4 13 15 13 15 0 9 7 15 13 14 13 2 16 15 13 16 15 4 13 0 9 1 12 9 2 3 15 4 4 13 8 1 9 10 13 14 4 13 1 3 3 2
16 7 4 13 10 9 1 9 7 15 3 13 14 4 13 1 2
8 3 13 15 12 9 1 11 2
25 15 13 10 9 9 1 11 7 15 13 16 15 13 12 9 1 11 2 10 9 9 7 9 9 2
18 11 13 10 9 9 7 3 4 15 13 10 16 11 4 3 13 12 2
15 3 15 13 10 0 0 2 3 13 15 12 9 1 11 2
28 0 9 2 10 11 13 1 10 9 11 1 10 0 9 9 2 10 11 13 10 13 1 9 11 1 9 7 9
9 16 15 13 13 9 1 11 2 5
43 3 2 15 4 4 4 13 7 13 2 13 13 10 9 7 13 1 10 0 9 1 10 9 2 3 0 7 0 2 13 9 10 4 4 4 13 13 10 9 1 9 3 2
8 9 1 0 11 9 1 11 2
34 15 13 10 9 3 1 11 10 9 2 7 15 4 13 14 13 10 9 1 10 0 9 9 9 15 13 16 3 3 10 9 9 3 2
17 15 13 15 13 1 10 11 11 9 7 4 14 13 15 1 15 2
32 15 2 9 2 13 16 15 13 15 9 9 2 9 1 0 9 7 13 15 1 10 9 1 10 9 13 15 9 9 1 15 2
25 12 9 1 10 0 9 0 9 13 15 9 2 7 3 15 4 13 10 9 13 15 1 15 9 2
9 10 2 15 4 2 13 9 9 2
16 15 13 3 0 16 15 13 7 4 13 14 13 15 9 3 2
3 10 9 2
5 15 13 11 11 11
13 15 13 10 0 9 14 13 10 9 1 10 9 2
22 6 2 15 13 3 14 13 1 3 1 10 9 2 7 15 4 13 14 13 0 9 2
36 7 16 1 15 9 15 13 1 9 12 9 2 7 15 13 14 13 1 10 9 2 15 4 15 13 2 4 15 13 15 1 7 1 0 9 2
15 16 15 4 13 14 13 3 2 3 1 10 9 2 13 2
14 16 15 13 14 13 2 1 1 0 9 2 3 13 2
29 15 4 3 3 13 15 1 16 15 4 13 14 13 10 9 1 10 9 16 15 13 0 10 9 4 13 14 13 2
28 9 3 4 13 3 0 3 13 0 15 13 10 9 7 3 3 0 9 14 13 15 9 7 13 10 0 9 2
5 11 11 13 13 2
28 15 11 11 13 13 1 9 16 16 10 9 9 4 13 1 2 9 2 7 10 9 4 14 13 1 10 9 2
19 10 9 3 13 14 13 3 3 15 13 1 10 9 7 13 15 3 3 2
6 4 9 13 10 9 2
10 13 15 0 14 13 3 1 9 9 2
2 9 2
6 13 0 0 1 15 2
17 15 9 4 14 13 3 2 15 13 9 2 13 11 13 1 15 2
4 15 4 13 2
12 15 13 10 11 7 4 14 13 10 10 9 2
14 15 3 13 15 13 1 9 3 13 1 9 1 11 2
37 15 13 1 10 9 9 7 10 9 13 10 9 3 16 15 13 1 10 9 2 13 10 9 1 9 1 9 7 15 4 14 4 13 1 10 9 2
2 13 11
8 0 9 9 1 11 1 11 2
26 15 4 13 1 10 9 1 10 11 1 11 12 2 7 15 4 13 1 11 2 11 2 11 11 2 2
14 10 9 4 15 13 1 7 3 4 15 13 15 9 2
14 10 3 10 3 7 15 4 3 13 1 1 10 9 2
12 13 11 7 11 7 13 15 15 13 3 1 2
25 15 9 13 1 10 11 10 12 9 7 3 7 15 4 13 16 11 11 4 13 10 0 9 3 2
13 11 1 11 2 11 1 11 7 3 11 1 11 2
14 13 13 13 2 15 13 10 9 16 13 10 0 9 2
5 13 10 9 9 2
21 1 15 0 12 9 3 1 10 11 15 13 2 11 11 2 13 1 11 2 11 2
11 15 13 10 0 9 7 9 15 4 13 2
13 15 13 10 0 9 14 13 9 1 11 11 9 2
25 15 3 13 1 10 9 2 7 15 4 13 16 15 13 10 9 15 4 13 0 9 1 9 3 2
19 15 4 14 13 14 13 14 13 1 10 9 2 10 2 9 9 1 11 2
21 15 3 13 10 0 9 14 13 10 0 9 16 10 9 15 13 2 3 15 13 2
9 10 9 4 13 3 0 2 9 2
5 15 3 13 11 2
18 15 3 13 0 9 1 11 2 11 11 2 7 10 9 1 0 9 2
12 3 15 4 3 3 13 10 9 15 13 9 2
20 0 1 10 9 13 15 13 1 12 9 2 7 10 1 10 9 13 3 0 2
24 16 15 13 14 13 3 16 13 1 10 10 0 0 9 10 9 2 11 4 13 0 1 15 2
12 3 4 15 13 1 10 0 9 2 9 2 2
15 13 1 9 1 10 0 9 7 15 13 15 14 13 0 2
37 4 13 10 9 0 2 7 2 13 10 0 9 1 10 11 9 7 10 2 11 2 9 13 10 0 9 14 13 10 9 7 9 16 13 10 9 2
35 7 3 16 13 10 11 11 11 7 13 10 9 1 9 7 13 10 9 2 15 3 13 0 0 9 15 4 13 2 9 13 3 0 3 2
11 13 1 11 4 14 13 0 1 12 9 5
10 9 9 1 10 9 2 13 1 9 2
15 15 13 0 2 15 4 14 13 14 13 9 1 9 14 13
16 14 13 9 2 15 13 0 2 3 16 9 13 3 2 15 4
15 13 2 7 16 15 13 14 13 15 2 15 3 13 6 2
4 13 14 13 2
16 15 13 14 13 10 12 9 9 2 15 4 15 13 15 1 2
5 15 4 13 9 2
13 3 10 9 9 1 10 9 1 0 9 1 3 2
7 15 4 3 13 9 3 2
19 15 13 9 13 10 9 2 4 15 13 15 10 0 9 9 1 15 3 2
16 15 4 13 10 9 10 13 10 3 16 13 1 10 10 9 5
54 3 13 10 9 1 15 12 9 9 15 13 15 1 12 1 10 9 1 1 10 9 10 12 9 1 12 9 1 9 9 9 9 9 9 9 12 12 9 9 10 9 7 12 12 9 9 9 1 12 9 9 12 0 9
16 16 15 13 1 10 9 9 15 4 13 10 9 12 9 9 2
6 13 15 1 9 5 6
16 1 10 9 10 9 15 4 13 9 7 9 10 9 0 9 2
5 3 13 10 9 9
6 0 9 2 0 9 2
6 0 9 7 0 9 2
6 11 11 13 10 0 2
6 0 0 9 0 9 9
6 15 13 3 0 2 5
6 0 9 1 10 9 5
6 10 10 0 9 13 15
7 10 9 13 14 13 1 2
7 0 13 9 1 10 9 2
7 0 7 0 9 1 9 9
7 0 9 15 4 3 13 2
8 10 0 9 1 10 11 11 2
8 15 13 0 1 11 7 11 2
8 0 0 9 2 15 13 15 2
4 9 13 0 2
5 9 13 3 0 2
9 15 13 10 9 3 0 9 1 15
9 3 0 9 1 10 9 1 0 9
4 6 6 6 2
5 10 0 9 1 11
9 0 9 7 0 9 3 0 9 2
2 11 11
7 11 11 13 10 11 11 2
1 0
9 15 13 10 0 0 0 7 0 9
7 15 13 10 9 11 13 2
2 0 9
3 0 9 2
7 9 9 2 9 16 13 2
6 0 9 2 9 11 2
4 0 9 9 2
10 0 9 10 15 4 13 3 3 2 5
5 10 3 0 9 2
6 10 9 13 3 0 2
5 10 9 13 0 2
6 7 10 9 13 0 5
9 6 15 13 10 9 15 13 3 2
2 0 2
4 3 0 9 2
5 0 3 7 3 2
3 0 9 2
7 15 13 15 0 9 9 2
4 3 13 11 11
12 3 0 9 2 3 0 9 2 3 0 9 2
10 13 15 16 13 10 9 1 15 9 2
2 9 2
12 15 13 10 0 11 14 9 15 4 3 13 1
6 13 14 13 10 9 2
7 9 13 0 7 13 9 2
3 0 9 2
7 0 1 10 9 1 9 2
3 9 3 2
4 10 9 13 0
6 0 9 2 0 9 2
3 3 13 3
6 0 9 2 0 9 2
7 13 11 7 13 0 9 2
13 13 16 15 13 1 11 2 7 9 9 13 0 2
8 0 9 7 0 9 13 0 2
6 13 14 13 1 0 9
6 3 3 0 7 0 2
7 11 11 13 15 9 3 2
13 10 0 9 1 11 11 13 9 10 10 9 13 2
4 0 0 9 2
10 15 13 1 11 3 7 13 15 9 2
11 13 10 0 9 16 13 15 9 1 11 2
3 9 11 2
9 0 0 3 13 0 9 7 9 2
3 0 9 2
3 0 9 2
4 4 14 13 2
11 15 13 0 14 13 3 10 9 4 13 2
8 10 0 0 9 7 9 9 2
7 9 7 9 13 3 3 2
4 9 13 0 2
8 15 13 13 1 10 9 9 2
4 9 13 0 2
16 0 14 13 10 10 0 9 7 0 9 7 10 9 4 13 0
1 11
8 15 4 3 13 11 1 11 2
7 0 9 9 7 0 9 2
17 15 13 10 9 9 1 9 14 13 1 7 9 13 1 10 9 2
13 13 10 10 9 3 1 10 9 2 13 1 12 2
4 15 13 15 2
17 15 13 10 0 12 9 9 9 9 1 10 9 15 4 13 1 2
11 0 9 1 15 9 7 10 9 13 0 2
7 4 13 3 1 10 9 2
3 11 1 11
3 0 9 2
10 13 1 15 9 7 13 9 1 15 2
2 9 2
3 0 9 2
14 13 0 14 13 0 9 1 15 9 14 13 15 0 2
1 6
5 15 13 10 11 14
13 15 3 13 10 9 7 15 13 10 11 14 11 2
2 9 2
5 3 0 9 13 2
4 13 15 1 2
6 2 11 11 11 11 11
18 0 1 15 9 2 15 13 10 0 9 15 4 13 1 10 0 11 2
13 9 14 7 9 9 2 1 10 9 12 9 9 2
5 9 9 2 0 11
9 15 13 10 0 9 14 13 10 9
11 15 13 14 13 10 9 3 2 15 13 0
1 0
8 0 9 9 15 4 3 13 2
11 11 13 0 2 15 4 13 15 1 9 2
6 15 9 13 9 3 2
14 15 3 4 14 13 1 3 12 9 15 4 14 13 2
6 9 1 11 11 11 9
14 10 9 1 11 13 0 2 0 7 10 9 14 13 2
7 0 2 0 2 0 9 2
14 9 4 13 10 9 0 7 15 13 10 3 3 0 9
3 0 9 2
12 15 3 13 10 0 9 1 10 11 11 9 2
6 0 2 0 7 0 2
21 9 4 13 1 10 9 2 7 3 10 0 13 2 1 9 9 1 10 11 11 2
2 13 3
3 0 9 2
3 3 0 2
13 13 9 15 13 15 3 14 13 7 4 3 13 2
2 3 13
9 15 12 9 0 9 13 10 9 2
6 10 0 9 9 3 2
4 6 1 11 2
9 10 9 13 0 2 7 3 0 2
14 3 4 15 13 10 9 2 1 10 9 1 9 2 2
2 9 9
17 10 9 9 13 0 2 15 0 0 9 13 12 7 9 12 12 2
2 13 15
10 10 9 1 11 11 11 13 3 0 2
5 7 13 0 9 2
8 15 13 3 0 1 10 9 2
22 15 13 10 0 2 0 9 7 10 0 9 7 4 3 13 11 11 11 7 11 3 2
22 15 13 15 13 11 2 11 11 11 2 15 13 15 3 2 7 10 9 15 13 0 5
2 0 9
14 15 13 10 0 9 1 11 14 11 2 9 7 9 2
7 10 0 9 13 14 0 2
1 11
8 3 0 9 13 10 0 9 2
8 13 13 9 3 3 1 9 2
8 13 15 13 1 1 10 9 2
20 0 9 3 1 10 9 9 7 10 9 3 13 10 0 9 15 4 3 13 2
4 4 14 13 3
24 9 1 9 4 13 2 9 13 0 2 9 13 3 3 0 1 11 1 9 2 0 9 13 0
3 0 7 0
10 10 9 13 9 9 12 1 10 11 2
7 15 13 3 0 1 9 2
5 4 14 13 15 2
10 0 9 2 0 9 2 7 0 9 2
16 7 10 9 4 14 13 9 1 15 16 15 13 0 7 14 2
12 12 1 10 0 0 9 15 4 13 1 11 2
13 7 1 10 9 10 13 1 0 9 9 2 3 2
11 0 9 9 2 0 9 15 4 3 13 2
14 0 9 10 13 3 13 2 0 14 13 3 1 9 2
2 11 11
23 9 2 9 2 9 7 9 2 9 9 2 9 9 2 9 2 9 9 2 9 9 9 2
1 11
9 10 0 9 9 13 1 0 9 2
10 10 0 11 13 14 13 1 0 9 2
6 9 7 9 1 9 2
5 4 3 13 3 2
5 3 0 7 0 2
17 10 9 13 1 7 1 10 9 1 10 9 1 10 0 9 13 2
2 11 9
9 15 13 10 0 9 1 10 9 2
8 15 13 3 16 15 13 12 2
8 3 15 4 13 3 0 9 2
3 11 10 11
5 0 9 1 9 2
6 0 9 7 0 9 2
13 9 3 0 9 1 11 2 9 1 10 0 9 2
10 11 7 15 9 10 13 10 0 9 2
6 3 0 7 0 9 2
11 0 9 1 15 7 10 1 15 9 9 2
5 10 10 9 13 9
21 15 13 15 9 1 9 7 9 7 13 16 15 4 13 10 0 9 1 15 9 2
10 3 0 9 13 15 9 13 1 11 2
16 0 9 16 13 15 13 1 11 11 10 4 13 1 10 0 9
11 0 9 14 13 2 15 4 13 3 3 2
18 9 13 0 2 9 1 9 14 13 1 9 2 7 0 9 1 9 2
4 0 9 1 11
9 15 4 4 13 11 11 1 9 2
12 15 4 3 13 10 0 9 1 10 0 9 2
3 3 13 2
3 3 0 2
21 0 7 10 9 13 0 7 13 1 10 9 3 15 13 3 0 9 1 10 9 2
5 15 4 14 13 2
26 10 3 0 9 2 0 9 7 3 1 15 13 0 1 15 9 2 8 9 4 3 13 7 13 2 2
13 15 13 11 11 12 9 16 15 9 13 3 0 2
15 3 2 15 4 14 13 15 3 0 7 15 9 13 0 2
3 3 0 2
7 9 7 9 1 10 9 2
12 15 9 4 14 3 13 0 9 15 13 3 2
7 3 0 1 3 3 0 9
7 10 9 7 9 13 0 2
12 15 13 1 11 11 15 13 0 9 1 15 2
11 15 13 1 3 10 3 13 9 1 11 2
29 10 9 13 0 7 15 3 13 14 13 3 16 15 13 0 2 3 15 13 3 2 3 2 7 13 3 1 15 9
3 13 9 2
15 10 0 12 2 0 9 2 11 13 9 15 4 3 13 2
11 15 3 13 2 10 9 9 1 11 11 2
4 11 13 0 2
16 11 13 0 2 3 0 9 1 10 0 9 2 0 9 9 2
6 10 9 13 3 0 2
4 7 15 13 2
4 10 10 9 2
18 16 15 13 10 0 1 15 9 2 4 14 13 16 13 10 0 9 2
9 15 13 10 3 0 1 10 11 2
4 10 10 9 2
5 10 9 13 0 2
11 10 9 13 7 10 9 13 3 3 0 2
7 15 4 13 3 7 3 2
6 3 4 14 13 3 2
2 9 9
18 11 11 13 15 1 0 9 7 13 1 10 0 9 1 9 7 9 2
10 15 9 7 9 13 1 10 0 9 2
11 9 13 3 0 3 13 10 9 10 9 2
20 3 3 3 16 14 15 13 1 1 10 0 9 1 0 0 9 1 10 9 2
2 10 9
10 15 13 10 9 1 10 9 15 13 2
11 10 9 13 0 2 0 2 0 7 0 2
9 15 3 13 0 7 13 3 0 2
5 10 9 3 13 2
16 10 1 10 9 3 13 3 0 15 13 0 1 15 1 9 2
10 10 13 10 0 9 15 4 13 1 2
3 11 11 11
11 0 9 2 3 13 1 3 15 13 15 2
17 15 4 13 0 0 9 9 1 3 2 15 4 13 1 11 11 2
3 14 0 3
17 15 13 10 0 9 2 15 13 3 10 0 0 1 10 11 9 2
13 9 0 1 15 2 3 0 9 1 10 9 9 2
2 0 9
12 2 13 15 3 3 1 10 0 9 3 13 2
7 15 13 9 1 10 9 2
13 15 9 7 9 4 4 13 1 15 1 9 2 2
6 10 9 1 11 9 2
18 15 13 15 0 9 3 3 14 13 10 9 14 13 3 1 15 9 2
6 7 10 9 13 0 2
4 3 0 9 2
3 13 11 11
5 10 9 13 0 2
6 11 7 11 13 0 2
13 15 13 3 3 14 13 10 1 15 9 7 9 2
9 10 9 14 13 1 10 9 3 2
3 0 9 9
30 11 14 11 9 13 3 3 3 3 0 9 1 10 0 9 2 13 10 9 9 1 1 12 5 7 10 0 9 9 2
17 15 4 13 14 13 15 9 9 15 13 15 9 1 11 11 9 2
13 10 0 9 2 13 10 0 9 13 10 9 0 2
4 0 9 11 2
21 10 0 0 9 15 4 3 13 1 11 2 3 0 7 3 0 9 1 0 0 2
14 10 9 13 10 3 0 0 9 1 11 2 3 13 15
4 0 7 0 2
10 3 0 2 0 2 0 7 0 9 2
21 11 13 10 0 9 1 9 2 9 7 10 9 14 13 9 1 2 1 0 9 2
2 6 2
5 0 9 2 0 9
6 10 9 13 3 0 2
13 15 9 4 14 13 3 16 13 2 10 9 2 2
12 0 1 10 9 1 9 7 10 9 1 9 2
4 0 0 9 2
22 10 9 3 13 15 9 2 15 13 3 9 15 4 13 1 9 1 9 7 9 9 2
8 3 11 11 9 9 2 4 13
3 3 0 2
4 15 10 9 2
13 15 4 14 13 10 0 9 1 15 9 1 9 2
3 0 9 2
3 3 0 2
8 10 9 13 15 15 4 13 2
4 9 14 13 2
3 0 9 9
12 13 9 13 10 9 2 15 3 13 1 9 2
21 3 15 13 14 13 15 15 13 2 3 15 13 14 13 1 10 9 7 3 0 2
18 6 2 10 9 13 3 3 7 3 16 13 15 1 15 9 9 9 2
18 15 13 10 0 9 15 13 14 13 1 13 9 14 13 1 1 15 2
2 0 9
6 3 4 14 4 13 2
14 13 12 9 16 13 14 13 16 10 9 13 1 9 2
6 13 16 15 13 9 2
7 13 3 7 15 13 9 2
3 3 0 2
15 4 14 13 15 13 1 10 0 9 1 9 1 0 9 2
22 15 9 13 3 3 0 15 13 10 0 9 14 13 3 3 0 1 10 9 15 13 2
8 0 9 9 9 1 10 1 11
11 11 11 9 1 10 11 11 11 9 9 2
16 15 13 15 9 9 1 10 1 15 9 9 9 7 9 9 9
8 3 0 7 0 9 9 9 2
12 15 13 1 0 9 2 0 2 7 9 9 2
17 10 9 13 15 15 4 13 7 13 15 1 10 9 1 15 9 2
31 10 9 9 13 3 0 2 15 13 16 10 9 13 10 0 2 10 9 13 3 0 7 10 9 2 6 10 9 1 15 2
7 6 2 15 13 3 0 2
25 15 13 0 9 2 13 10 0 9 1 10 9 2 7 10 12 9 1 10 9 13 10 9 3 2
8 15 13 10 9 1 15 9 2
6 15 4 13 3 3 2
4 1 1 9 2
10 15 13 10 9 13 3 3 1 9 2
14 16 15 13 8 2 15 4 14 13 15 1 10 9 2
12 15 4 13 14 13 12 9 1 12 1 11 2
3 0 9 9
14 11 11 13 15 13 1 0 9 1 10 9 1 9 2
16 10 9 4 13 1 12 9 2 7 9 4 13 1 1 9 2
4 3 13 9 2
2 0 0
37 10 9 9 13 12 1 10 0 3 10 9 13 0 7 0 7 10 9 9 13 10 0 2 13 15 0 9 13 7 10 0 0 9 1 10 10 9
2 13 0
21 15 3 13 14 13 15 9 16 15 13 14 3 0 1 15 0 9 15 3 13 2
15 3 15 4 13 9 15 4 13 14 13 15 15 3 13 2
3 3 13 9
22 10 9 13 10 3 13 9 15 4 3 13 15 13 3 10 0 9 15 4 3 13 2
14 15 4 14 13 10 9 1 9 7 3 9 14 13 2
3 3 3 0
5 3 0 10 9 2
5 0 7 8 0 2
13 15 13 16 16 15 13 1 10 8 0 11 11 2
12 15 4 13 14 4 13 10 0 9 14 13 2
4 7 14 3 2
11 15 4 13 11 11 1 10 0 12 9 2
11 15 13 12 9 3 7 15 13 10 0 2
5 15 13 1 9 2
14 15 9 4 4 13 9 1 7 13 1 10 0 9 2
4 0 9 0 9
18 11 13 3 5 12 14 13 15 9 7 10 9 13 15 1 5 12 2
4 13 15 9 2
15 13 15 13 1 10 0 9 2 13 14 13 10 9 2 2
2 0 9
9 10 9 13 10 0 9 7 9 2
12 15 9 13 0 1 10 0 9 1 12 9 2
19 3 3 0 7 10 9 13 14 1 10 2 13 3 8 13 15 2 9 2
17 0 9 13 15 12 9 3 7 15 3 13 15 9 12 9 3 2
22 15 9 3 13 0 7 0 9 1 10 11 11 11 15 4 13 15 9 3 3 3 2
5 10 9 1 9 2
21 15 13 3 0 3 15 13 1 11 11 2 15 13 10 9 7 10 9 13 0 2
17 15 13 14 13 1 10 9 14 13 12 0 9 2 15 10 9 2
4 13 10 9 0
21 15 4 13 11 11 7 15 9 3 3 1 15 9 7 10 9 4 13 3 0 2
17 15 4 14 13 14 13 15 3 7 13 15 1 15 9 7 9 2
9 11 11 13 10 3 0 0 9 2
14 15 13 0 16 9 13 15 1 15 1 15 0 9 2
18 15 13 10 9 9 9 7 13 10 9 1 10 9 10 11 11 13 2
6 0 9 15 4 13 1
6 13 3 1 12 9 2
8 10 9 13 3 0 7 0 2
11 10 9 13 3 0 7 10 9 13 0 2
12 0 9 7 1 9 9 13 15 9 3 0 2
10 10 9 13 0 9 1 3 0 9 2
26 15 4 13 15 12 9 16 13 9 16 13 1 10 9 1 10 9 16 13 10 9 1 15 0 11 2
6 15 4 3 4 13 2
8 4 14 13 15 9 1 10 9
32 10 9 13 10 9 7 15 13 10 0 9 1 10 9 3 15 4 13 9 15 4 14 13 2 7 15 13 1 13 1 15 2
4 3 0 9 2
3 13 11 11
22 4 3 13 3 13 10 9 13 3 10 13 15 9 13 1 10 0 9 1 10 9 2
18 10 9 2 9 13 2 8 9 2 9 7 0 9 3 1 10 0 9
1 9
19 13 12 5 9 14 13 1 11 2 9 1 9 2 9 4 14 13 9 2
15 13 10 9 1 10 9 9 9 13 1 11 7 11 11 2
10 13 1 11 11 2 12 9 5 9 2
2 0 9
7 3 0 9 7 0 9 2
17 10 9 13 0 7 3 13 10 9 9 2 9 13 0 2 5 2
14 15 13 10 0 2 0 9 14 13 9 13 7 13 2
6 15 13 16 13 3 2
3 0 9 9
18 15 13 10 9 1 10 9 13 16 15 9 4 13 3 1 9 2 5
5 15 13 3 0 2
17 11 13 10 0 9 9 15 4 3 13 7 15 4 3 13 15 2
5 0 3 2 0 3
12 10 9 3 13 0 3 2 9 13 3 0 2
10 3 0 9 10 15 3 3 13 3 2
19 10 9 1 10 9 13 0 2 4 14 13 9 3 13 15 4 13 9 2
3 0 11 9
23 15 13 1 11 7 15 13 15 9 1 11 7 15 13 0 3 15 13 15 4 13 11 2
19 15 13 1 13 3 0 9 11 9 7 15 13 0 1 10 0 11 9 2
3 11 1 11
28 15 9 9 13 3 0 7 3 13 7 10 9 9 13 3 3 0 1 15 7 4 14 13 14 13 13 9 2
11 0 9 2 3 13 2 1 9 3 3 2
3 0 9 2
3 0 9 2
4 13 10 9 2
9 13 10 9 1 10 11 11 11 2
8 9 13 0 1 11 7 11 2
13 4 14 13 1 10 9 1 11 2 15 13 0 2
3 0 9 2
5 13 1 11 11 2
4 15 13 15 2
4 0 9 3 2
6 3 0 7 0 9 2
18 15 4 13 0 9 1 15 9 2 7 11 11 13 1 3 15 0 2
19 15 3 13 1 10 9 9 0 1 12 9 7 10 9 13 0 7 0 2
8 15 13 10 0 9 14 13 2
26 15 4 13 10 0 9 1 10 9 16 15 13 2 7 13 10 9 16 10 1 10 9 13 0 9 2
14 3 10 9 15 13 10 0 9 2 15 13 3 0 2
1 0
10 11 13 10 0 9 9 1 10 9 2
3 3 13 2
15 16 15 13 0 9 2 15 4 13 1 11 14 11 11 2
5 16 15 13 0 2
8 15 13 10 9 12 5 12 2
4 12 9 3 2
3 6 6 2
8 0 9 9 7 0 9 9 2
16 10 9 13 0 14 13 7 15 13 10 9 3 1 10 9 2
15 10 9 9 7 10 9 9 13 3 0 14 13 3 1 2
9 15 3 13 11 11 1 15 9 2
2 6 2
36 6 2 15 4 14 13 10 9 2 7 3 1 10 9 4 15 13 15 9 9 10 13 10 9 11 2 13 15 9 1 10 9 1 10 9 2
10 6 15 13 3 0 1 10 9 2 6
4 0 7 0 9
15 15 13 9 9 1 3 10 10 9 7 15 13 3 0 2
8 10 9 13 3 0 7 0 2
23 15 4 13 10 9 1 10 0 9 7 3 13 15 3 15 15 13 7 15 13 3 0 2
15 15 3 13 14 13 10 9 16 15 13 3 1 10 9 2
19 3 2 15 4 13 15 10 9 1 9 1 0 9 7 13 14 13 13 2
16 10 9 4 14 3 13 14 13 15 15 4 13 7 15 13 2
3 9 9 2
25 15 13 0 1 10 9 7 15 13 0 15 4 4 13 10 9 7 10 9 7 13 14 13 3 2
16 15 13 15 9 1 1 11 7 13 1 11 1 10 0 9 2
7 4 13 9 1 15 3 2
2 0 9
45 15 1 11 11 11 13 0 1 15 9 7 10 0 9 15 13 14 13 15 9 13 3 2 15 4 13 15 0 9 16 9 13 3 7 15 4 13 15 1 0 9 1 0 9 2
8 4 14 13 10 9 1 15 9
11 1 10 9 11 13 16 15 4 13 0 2
9 15 4 14 13 3 1 10 9 2
13 10 9 13 0 2 7 10 9 4 14 4 13 2
12 10 9 13 0 2 7 15 13 10 0 9 2
3 0 9 2
15 10 9 1 11 11 11 13 3 0 7 0 14 13 1 2
20 15 13 15 1 10 10 9 0 1 10 10 9 9 16 16 15 13 10 9 2
11 15 13 15 3 0 7 4 3 13 15 2
1 9
1 11
7 10 0 9 13 1 11 2
13 3 0 7 0 2 9 13 0 9 7 3 0 2
22 15 3 13 1 15 15 13 15 4 13 14 13 2 7 15 13 3 0 1 15 9 2
7 15 4 3 13 15 9 2
2 0 9
42 15 13 14 13 15 9 3 10 10 9 2 7 9 13 9 3 3 2 10 9 4 13 0 2 7 15 3 13 14 2 13 1 2 0 9 2 10 3 4 14 13 2
6 15 4 14 13 3 3
2 0 9
18 10 9 13 3 0 10 9 7 13 9 14 13 1 15 9 7 9 2
19 15 4 3 13 1 10 9 3 3 7 15 13 3 0 2 15 13 0 2
12 10 0 9 9 15 4 13 1 1 0 9 2
4 3 0 9 2
18 11 13 10 0 9 9 2 9 15 4 3 13 1 1 15 0 9 2
8 15 13 10 9 13 15 3 2
17 15 13 3 3 0 2 3 2 10 13 10 0 9 1 15 9 2
5 15 13 10 0 2
1 9
26 10 9 13 14 13 10 9 3 3 2 3 13 14 13 10 0 1 15 9 2 14 16 15 13 15 2
18 7 3 15 4 14 13 10 0 9 16 15 13 9 1 15 9 9 2
6 10 4 13 10 0 9
9 15 13 10 9 14 13 15 9 2
14 10 9 15 13 13 0 3 15 13 6 15 13 0 2
29 16 15 13 1 15 13 10 0 9 14 13 15 9 13 2 15 13 10 10 9 1 9 7 10 9 13 3 13 2
5 9 13 9 1 11
19 3 13 15 14 13 16 11 13 3 16 13 9 7 13 15 9 1 9 2
24 15 13 14 13 3 0 15 13 16 15 14 13 0 10 0 9 4 13 3 15 13 15 9 2
3 13 15 2
4 10 0 9 2
4 15 13 0 2
6 15 3 13 0 9 2
8 15 3 13 3 13 9 9 2
6 15 9 13 3 0 2
6 15 0 9 13 0 2
19 15 4 14 13 10 9 0 9 2 7 15 3 4 14 13 15 10 9 2
3 0 9 2
7 9 9 0 15 13 14 2
12 13 3 7 15 4 14 13 15 13 1 11 2
18 10 9 13 1 10 9 9 1 11 2 0 2 0 2 7 1 9 2
10 13 0 9 2 0 9 2 7 13 2
6 0 1 11 3 3 2
4 0 0 9 2
2 3 13
15 15 13 1 10 0 9 9 7 4 13 3 1 15 9 2
8 3 10 0 9 3 1 9 2
5 0 9 7 9 2
4 0 7 0 2
6 9 1 10 0 9 2
10 4 3 13 3 3 15 13 0 9 2
3 9 1 11
17 15 4 3 13 15 11 11 0 9 13 1 10 9 1 11 11 2
29 10 9 15 13 3 13 0 2 0 7 3 0 7 4 13 15 3 3 16 15 4 1 15 9 1 9 3 9 2
3 3 13 2
4 15 0 9 2
16 15 9 7 15 13 3 3 1 10 9 1 10 9 1 11 2
12 3 3 15 13 10 0 9 1 9 1 9 2
23 6 15 9 13 1 9 0 7 15 13 1 10 8 0 9 1 10 3 0 9 1 9 2
3 10 0 9
7 0 9 2 9 7 9 2
10 13 7 13 7 0 9 7 0 9 2
21 10 9 13 0 9 1 10 9 7 13 0 16 15 13 10 0 9 7 9 9 2
14 3 10 3 0 9 4 13 3 14 13 1 11 14 2
2 0 9
19 15 4 4 13 3 16 15 13 10 0 9 7 13 10 0 7 0 9 2
10 11 11 4 3 13 3 0 7 0 2
23 15 4 13 11 11 1 9 15 13 1 9 1 10 0 9 7 4 13 1 10 0 9 2
2 9 9
34 13 15 7 14 2 7 10 9 9 4 13 3 0 1 15 9 9 10 13 7 4 14 13 3 14 13 3 15 13 16 13 9 9 2
13 15 3 13 15 9 7 15 4 13 9 15 13 2
5 9 3 2 11 2
18 11 13 13 10 9 1 15 9 14 9 7 15 4 14 4 13 0 2
30 15 13 1 12 9 14 13 10 0 9 10 4 13 15 9 1 10 9 15 13 14 7 11 7 15 9 13 15 13 2
6 15 13 0 10 9 2
6 0 9 7 3 0 9
16 15 4 13 3 0 9 7 10 9 10 9 13 0 1 0 2
22 12 9 15 3 13 16 13 1 10 9 1 12 9 7 14 4 13 1 10 9 9 2
2 0 2
10 15 4 13 10 0 0 9 1 11 2
11 15 13 1 9 1 10 0 9 1 9 2
18 0 9 15 13 3 2 15 9 13 0 7 10 9 13 0 2 0 2
27 15 13 10 0 9 9 1 9 1 10 1 15 9 2 3 15 4 13 3 0 9 14 13 13 2 13 2
5 0 0 0 9 9
26 15 4 13 0 7 3 3 13 9 9 1 10 9 7 11 11 13 0 9 2 0 9 7 3 0 2
24 16 0 4 13 0 13 1 9 1 11 11 15 13 0 1 10 9 7 9 15 13 1 11 11
4 3 0 9 2
13 10 9 13 3 3 0 2 13 15 0 7 0 2
21 10 9 13 0 7 0 2 7 15 3 4 14 13 1 1 10 0 2 0 9 2
19 15 13 12 0 9 1 9 2 15 13 3 10 0 3 15 13 1 9 2
3 10 9 2
22 15 13 1 10 9 7 10 9 13 12 1 15 9 1 10 0 2 0 7 0 9 2
16 13 1 7 13 9 0 1 10 11 11 2 10 9 13 0 2
16 0 7 0 9 2 15 13 15 9 3 15 13 1 10 9 2
7 1 9 2 0 7 3 0
11 15 13 1 10 9 1 1 13 9 9 2
7 13 9 1 12 11 9 2
8 11 13 3 1 10 13 9 2
17 15 13 3 0 2 3 0 14 13 1 7 13 10 3 0 9 2
3 3 13 2
2 9 11
3 11 11 2
10 0 9 9 13 1 9 1 9 7 9
26 11 13 0 9 9 10 4 3 13 10 9 1 15 9 7 9 7 13 9 7 9 3 1 10 9 2
20 15 13 7 13 0 16 13 2 13 7 13 10 0 9 7 13 9 14 13 2
