599 11
33 9 9 9 9 9 9 13 2 10 9 0 0 1 9 9 9 9 0 1 9 9 13 7 9 1 9 9 1 1 1 9 13 2
36 15 9 9 9 0 14 1 9 1 1 9 9 0 13 7 13 2 0 9 7 9 9 0 1 9 1 9 1 9 0 1 0 9 9 13 2
45 9 9 9 9 9 9 9 13 16 0 9 9 9 7 9 4 1 9 7 9 9 1 9 0 7 0 1 9 9 9 7 9 1 9 9 2 9 7 9 10 9 1 9 13 2
26 0 9 9 9 7 9 1 9 9 9 9 9 1 12 1 12 9 9 1 9 9 9 9 0 13 2
30 9 0 7 9 9 9 7 9 7 9 9 13 2 1 9 0 9 9 0 1 9 0 9 0 1 9 13 13 13 2
20 15 13 2 9 13 1 9 10 9 9 9 2 1 9 0 9 0 13 13 2
42 9 9 9 9 2 1 9 10 9 1 9 13 2 9 9 0 1 0 9 12 7 12 15 2 1 9 9 0 7 0 0 1 9 9 9 7 9 9 0 4 13 2
32 15 13 2 1 10 9 9 9 9 7 9 1 9 0 1 9 0 9 13 7 9 13 16 1 9 0 9 9 16 0 13 2
47 15 1 9 1 10 9 16 9 9 0 1 9 9 9 3 4 13 13 2 9 9 9 7 9 9 0 1 9 7 7 9 9 9 9 1 12 9 9 1 9 9 9 7 9 4 13 2
37 9 9 9 1 9 1 9 9 9 9 10 9 13 2 1 9 9 0 0 1 9 9 0 2 9 9 7 9 9 0 0 7 0 9 9 13 2
11 1 10 9 15 1 9 9 9 0 13 2
4 9 2 9 2
27 9 0 9 0 9 9 13 2 9 9 9 0 0 7 9 9 3 1 9 1 9 9 0 1 9 13 2
35 9 1 9 9 9 7 9 13 2 10 9 9 13 16 9 9 9 0 1 9 0 1 9 9 9 0 0 1 9 0 9 0 13 13 2
31 9 0 16 1 9 9 9 10 9 9 13 13 1 9 9 13 2 1 10 9 2 9 3 1 9 9 0 9 4 13 2
44 1 0 9 9 2 3 9 9 0 1 9 0 9 9 7 9 9 9 0 9 16 9 0 1 0 9 0 9 0 14 9 13 16 4 1 9 9 1 9 9 0 0 13 2
31 9 9 13 3 1 9 9 0 9 9 9 1 9 9 9 0 9 16 9 13 9 0 9 9 15 13 13 2 9 13 2
26 9 9 9 9 9 0 9 9 9 9 9 9 9 14 9 1 9 0 9 7 1 1 9 0 13 2
48 15 9 13 2 3 15 0 9 13 16 9 9 1 9 0 15 1 9 0 9 13 7 15 3 15 13 16 15 16 1 9 9 9 9 1 9 10 9 2 9 9 7 9 9 9 9 13 2
51 9 9 0 13 2 3 10 9 9 16 1 9 9 0 1 9 7 9 0 13 2 9 9 15 14 1 9 9 1 12 9 1 9 0 7 9 0 9 13 16 9 0 14 1 9 9 1 9 13 13 2
24 10 9 1 9 9 9 13 7 9 13 16 9 9 9 1 10 9 1 9 0 9 9 13 2
46 1 10 9 16 9 4 13 1 9 9 2 9 7 9 2 9 9 2 9 7 9 7 9 9 14 1 9 13 7 1 9 9 0 2 9 9 9 9 7 9 0 9 14 9 13 2
72 9 9 1 9 1 9 9 9 13 13 2 1 1 9 9 9 1 9 9 1 9 9 9 7 9 0 1 9 9 7 9 9 9 16 9 9 0 7 0 1 9 0 9 14 1 9 9 7 9 7 9 7 9 9 13 1 15 2 9 1 9 7 9 0 1 10 9 1 9 9 13 2
35 9 13 3 1 9 9 0 9 9 7 9 9 15 9 0 0 9 1 15 9 0 9 13 7 9 0 9 1 15 14 1 9 9 13 2
21 7 2 9 0 9 9 9 7 9 9 9 9 9 10 9 7 9 9 13 13 2
25 0 13 9 13 16 1 9 9 7 9 10 9 0 2 0 4 10 9 14 1 9 9 9 13 2
27 16 9 3 9 9 1 9 13 7 9 15 14 9 13 7 0 13 2 4 15 14 1 9 9 0 13 2
19 9 2 9 7 9 9 0 2 1 9 9 1 9 7 9 9 9 13 2
8 9 9 14 1 9 9 13 2
6 9 9 14 9 13 2
18 9 7 9 9 14 1 9 13 7 9 9 1 9 9 14 9 13 2
32 16 9 1 9 10 9 0 13 1 3 9 9 7 9 0 9 7 9 9 9 1 9 9 7 13 7 13 14 1 9 13 2
18 9 1 9 9 9 7 9 13 7 1 1 9 0 15 9 9 13 2
10 1 3 9 1 9 3 9 9 13 2
18 3 0 13 3 9 1 1 15 9 9 7 9 0 1 9 0 13 2
9 9 9 15 9 1 3 9 13 2
23 0 9 9 1 9 9 0 1 9 9 9 9 13 7 9 0 1 9 9 14 0 13 2
27 7 15 16 3 0 9 14 1 10 9 13 1 9 1 15 9 13 2 1 10 9 9 3 9 9 13 2
16 16 10 9 9 12 9 0 13 3 9 1 1 15 0 13 2
12 1 9 1 10 9 3 4 1 9 0 13 2
6 4 9 1 3 13 2
20 1 9 13 9 0 1 9 4 1 9 0 1 13 7 9 0 1 15 13 2
37 9 7 9 0 9 4 9 13 7 9 1 9 9 0 0 7 9 1 9 0 9 13 7 13 7 9 0 7 0 14 1 9 0 9 9 13 2
27 1 10 13 7 13 9 0 9 0 1 9 9 13 7 9 1 9 0 1 9 7 9 1 9 9 13 2
22 1 9 10 13 7 13 9 0 1 9 15 9 0 7 9 1 9 15 14 0 13 2
22 1 9 3 13 7 9 9 0 0 13 7 9 16 9 14 1 9 9 13 0 13 2
11 9 10 9 9 7 9 1 9 9 13 2
6 4 1 15 9 13 2
9 15 4 1 9 10 9 9 13 2
17 9 0 7 0 9 9 16 1 9 15 2 9 3 13 2 2 2
47 13 13 2 9 0 9 1 9 0 9 9 12 9 14 1 9 9 9 7 9 0 14 1 9 9 9 7 9 13 7 1 10 12 9 13 1 1 10 12 9 7 7 9 9 0 13 2
34 9 1 9 16 1 9 9 9 1 9 9 1 9 13 2 13 16 9 15 14 1 1 9 7 9 9 0 13 7 1 15 9 13 2
23 7 1 12 9 9 13 9 0 0 14 13 7 9 0 0 7 0 14 1 15 9 13 2
27 9 9 9 9 9 9 9 0 3 1 12 9 0 9 9 0 9 1 9 9 1 9 7 9 9 13 2
24 15 16 1 1 9 9 13 7 1 15 1 9 1 9 9 2 9 2 1 9 9 9 13 2
17 15 13 2 9 0 9 9 2 9 9 7 9 9 9 4 13 2
27 15 9 0 7 0 13 16 16 1 0 9 9 9 0 13 7 7 9 9 9 1 9 9 14 0 13 2
25 1 1 10 9 2 9 9 9 9 14 1 9 9 9 0 9 16 1 1 9 9 0 9 13 2
29 15 13 13 2 9 9 0 9 13 16 1 9 0 9 2 9 7 9 1 9 9 1 9 7 9 9 13 13 2
14 9 0 9 1 9 13 16 9 9 14 1 1 13 2
13 1 9 0 9 9 1 9 9 7 9 0 13 2
31 1 15 1 9 0 1 9 0 10 9 0 13 2 7 9 9 9 9 1 9 9 9 0 9 3 0 7 0 9 13 2
25 0 13 16 10 9 3 9 0 14 9 13 7 3 1 9 9 0 9 1 9 0 9 9 13 2
18 9 0 9 1 9 9 9 0 9 13 2 9 0 15 9 9 13 2
33 1 9 9 0 7 9 1 9 9 2 9 9 9 1 9 7 0 9 9 2 9 14 0 7 9 15 14 1 15 3 0 13 2
29 1 9 9 9 0 9 3 9 9 9 0 7 9 1 9 9 16 1 9 0 1 9 1 9 9 13 0 13 2
36 15 16 0 13 13 9 9 0 1 1 9 9 7 9 15 16 1 1 9 9 9 7 9 9 0 13 3 15 16 1 9 9 7 9 13 2
53 3 16 9 9 9 13 13 15 9 0 14 1 9 9 0 7 7 9 1 9 7 9 9 7 9 1 1 9 9 9 13 2 16 9 9 0 1 9 0 0 13 2 3 9 1 0 9 9 1 9 9 13 2
20 9 9 1 9 9 9 9 9 0 13 2 9 9 9 9 0 14 9 13 2
27 10 9 13 13 2 9 15 15 13 16 9 0 9 0 1 9 9 14 13 7 9 9 0 14 9 13 2
43 9 9 9 2 9 9 9 9 0 2 1 13 7 13 1 9 9 9 2 9 2 1 9 9 3 13 2 9 10 9 9 14 4 1 9 1 9 9 12 9 9 13 2
27 9 9 0 3 13 9 15 14 1 10 9 9 13 7 10 9 15 15 13 13 16 9 9 14 0 13 2
49 15 1 9 1 9 9 9 9 9 9 2 13 2 1 9 9 9 9 13 16 1 9 9 9 0 9 3 0 13 7 13 7 9 14 9 13 7 7 3 9 9 14 1 9 0 1 9 13 2
81 9 9 9 9 0 16 1 9 15 16 9 9 9 0 9 9 1 9 9 2 9 7 15 9 9 9 13 13 2 9 13 2 9 16 1 9 9 0 13 15 13 16 15 9 7 9 16 1 9 9 12 9 1 9 0 1 9 7 9 1 9 13 0 13 7 9 10 9 14 1 9 9 7 16 12 12 9 0 0 13 2
18 9 16 1 9 0 13 16 15 13 16 9 9 14 1 9 0 13 2
21 15 1 9 9 13 2 1 10 9 3 15 9 9 13 1 9 9 15 9 13 2
37 9 2 1 9 1 9 1 9 9 0 9 1 9 9 1 9 9 0 2 13 2 16 1 9 0 9 9 0 9 13 15 15 9 9 9 13 2
42 15 1 9 13 2 15 1 9 9 15 3 13 16 9 0 1 9 0 14 1 9 13 2 3 7 16 10 9 14 13 3 1 9 9 0 7 0 15 16 4 13 2
74 9 9 1 9 2 9 9 12 12 2 13 13 2 3 1 15 16 9 9 1 9 9 9 9 9 9 1 9 1 9 7 9 13 7 9 9 3 9 9 9 14 9 13 2 9 0 9 9 0 0 13 2 9 9 7 9 1 9 1 9 7 9 13 7 9 13 1 9 9 9 14 9 13 2
73 3 1 9 12 9 7 0 9 9 9 9 9 9 0 1 9 9 1 9 1 9 0 16 9 13 16 1 10 9 0 10 9 14 1 9 0 9 9 13 1 0 15 16 9 9 3 1 9 9 7 7 1 9 0 7 0 9 0 9 9 9 15 14 1 9 0 0 3 1 15 9 13 2
32 3 1 15 7 12 9 1 9 0 9 13 7 0 9 9 0 9 1 9 1 15 0 13 9 9 16 1 15 1 9 13 2
22 9 9 9 1 9 1 10 9 9 1 9 2 9 1 9 1 9 9 2 0 13 2
32 3 9 9 2 9 9 9 13 16 10 9 9 1 9 1 9 9 0 9 1 9 9 3 1 1 9 9 0 9 9 13 2
20 3 9 9 9 13 16 9 1 1 9 0 9 9 9 1 9 0 9 13 2
6 13 1 15 9 13 2
41 1 9 2 9 9 0 1 15 13 16 12 9 1 12 9 13 13 2 15 3 9 9 1 9 15 7 9 9 14 1 9 0 7 9 9 9 14 0 4 13 2
17 9 9 9 0 9 1 9 0 1 12 2 12 12 9 0 13 2
37 15 13 2 1 9 1 9 9 0 2 1 9 0 10 9 0 9 1 9 0 3 13 13 7 1 12 9 9 1 12 12 7 12 12 9 13 2
32 9 9 9 1 9 12 14 12 9 9 13 7 9 9 9 0 7 9 9 9 0 1 9 0 14 1 9 0 9 9 13 2
39 15 13 2 1 9 12 1 9 9 9 0 2 9 9 16 9 12 2 12 9 9 13 2 7 1 9 12 9 9 9 1 9 12 2 12 9 9 13 2
29 9 9 13 2 1 9 0 0 9 9 1 9 12 9 1 9 9 13 16 1 9 10 9 12 9 0 9 13 2
16 9 1 9 9 16 1 9 0 9 0 1 12 9 9 13 2
40 9 0 9 0 10 9 16 9 1 9 0 15 9 9 13 2 14 9 13 7 1 9 9 0 9 12 7 12 1 9 9 9 1 9 9 0 0 9 13 2
15 15 9 0 9 1 9 9 9 9 9 0 9 14 13 2
19 9 0 9 1 9 9 7 9 0 1 9 1 10 9 9 1 9 13 2
15 1 9 9 0 1 9 9 2 12 12 12 9 9 13 2
24 9 2 9 12 7 12 7 12 9 3 1 9 2 12 9 9 12 9 1 0 9 9 12 2
30 15 9 0 9 1 9 9 9 0 7 9 9 9 12 1 9 9 1 9 9 7 9 0 14 1 9 0 9 13 2
45 9 9 9 7 9 9 13 2 9 9 7 9 0 13 9 12 12 12 9 1 9 15 1 9 0 14 16 9 9 15 0 1 12 12 9 1 9 13 2 1 9 0 0 13 2
44 9 9 1 0 9 9 9 1 9 9 7 9 9 7 9 13 2 1 9 9 9 1 9 0 1 3 12 9 1 10 9 9 7 9 12 12 9 1 9 0 9 9 13 2
29 9 9 9 7 9 9 13 2 9 0 1 9 9 15 1 9 9 9 0 1 9 1 9 0 9 0 9 13 2
66 9 1 9 1 9 0 9 9 7 9 1 9 9 0 13 2 1 9 16 9 0 1 9 9 1 9 9 9 1 9 9 13 7 15 14 1 9 9 13 9 9 15 1 9 12 9 9 4 13 7 16 1 1 1 9 9 13 12 9 9 1 10 9 9 13 2
25 1 9 15 9 9 7 9 9 9 9 0 1 9 0 14 1 12 9 1 12 9 9 4 13 2
35 15 9 13 2 1 9 9 0 1 9 9 0 10 9 0 1 9 0 9 13 7 9 9 1 10 9 0 1 9 7 9 0 4 13 2
36 9 9 13 2 9 9 0 4 1 0 9 1 1 9 12 9 0 0 9 13 16 4 0 1 9 9 7 9 9 1 9 9 9 0 13 2
14 9 9 3 1 9 9 2 9 2 1 1 9 13 2
18 16 9 1 9 0 13 2 9 7 9 1 9 9 1 1 9 13 2
6 9 13 2 6 9 2
17 16 9 1 9 9 2 9 2 9 14 1 9 15 9 13 13 2
17 13 2 1 15 9 13 3 15 7 9 2 9 2 14 9 13 2
16 9 13 2 3 1 9 15 1 9 9 2 9 2 9 13 2
11 13 2 10 9 15 1 9 15 9 13 2
14 3 15 14 9 13 2 1 10 9 7 9 13 13 2
16 9 13 2 15 9 13 16 9 7 9 15 14 1 1 13 2
8 9 13 2 8 8 8 8 2
2 9 2
7 9 15 1 9 15 13 2
31 9 13 15 16 9 9 2 9 2 14 13 7 9 2 9 2 14 9 7 9 9 13 9 3 3 7 15 13 9 13 2
38 1 10 9 2 16 9 9 9 1 9 9 13 16 9 9 1 9 1 9 9 13 2 9 9 14 9 13 2 7 9 14 1 9 9 9 0 13 2
19 9 1 9 9 13 16 1 9 3 9 0 7 0 9 1 9 9 13 2
16 9 1 9 9 7 9 7 9 9 9 13 1 9 9 13 2
4 9 9 13 2
9 7 9 9 2 3 9 9 13 2
5 9 16 9 13 2
16 9 9 1 9 13 2 9 1 9 1 9 9 7 9 13 2
14 1 9 16 3 12 9 0 1 9 1 9 13 13 2
9 9 16 9 15 14 0 13 13 2
12 15 16 1 9 7 9 1 9 13 9 13 2
12 7 7 7 15 15 2 9 2 1 9 13 2
17 9 1 9 7 9 7 9 7 9 8 9 2 9 2 9 13 2
14 1 9 16 13 16 15 9 14 1 9 9 9 13 2
23 1 9 1 9 2 9 15 14 1 9 7 0 1 1 9 8 9 2 9 2 9 13 2
11 1 1 9 9 13 16 3 0 15 13 2
38 1 9 0 16 9 1 9 7 9 7 9 7 9 8 9 2 9 2 13 1 10 9 13 0 1 9 7 9 9 9 1 9 9 7 9 9 13 2
19 1 9 13 2 15 13 15 14 1 9 9 9 1 9 9 1 9 13 2
27 1 0 15 7 9 15 1 9 15 13 2 1 9 13 2 9 9 14 9 13 7 1 9 15 9 13 2
7 9 16 9 13 0 13 2
8 7 15 1 15 15 0 13 2
26 1 9 13 2 15 3 13 16 15 15 14 1 1 15 9 13 7 1 15 7 9 15 9 9 13 2
10 1 15 9 13 16 15 14 0 13 2
8 16 9 13 9 9 4 13 2
12 7 16 1 9 9 13 1 15 0 4 13 2
24 1 9 9 13 16 9 15 9 9 1 1 9 7 9 9 13 2 3 9 9 1 9 9 2
13 9 15 1 9 9 2 9 2 0 1 15 13 2
73 9 9 2 9 2 14 1 9 0 7 9 1 9 9 13 7 15 7 9 9 2 9 2 1 15 15 7 9 15 7 9 9 2 9 2 13 2 8 8 8 8 8 8 8 2 8 8 8 8 8 8 8 8 8 8 8 8 8 8 8 8 8 8 8 8 8 8 8 8 8 8 8 2
18 1 9 15 9 13 13 16 3 9 13 1 10 9 9 9 13 13 2
19 0 9 1 9 1 9 16 3 15 1 9 7 9 7 9 13 9 13 2
28 3 1 9 9 9 13 2 1 9 13 7 10 9 14 1 9 13 7 9 15 7 9 15 7 9 9 13 2
22 10 9 9 16 9 9 9 13 16 2 8 8 8 8 2 9 9 2 9 12 2 2
14 3 15 16 1 9 9 13 15 14 0 7 0 13 2
17 9 9 2 9 2 9 1 9 13 16 9 15 9 9 9 13 2
31 3 9 9 2 9 0 1 9 9 9 2 9 16 1 9 9 2 1 9 9 13 13 7 1 9 7 9 9 13 13 2
13 9 9 2 9 2 1 9 13 2 9 15 13 2
27 0 13 16 1 9 15 9 1 15 13 16 9 15 14 13 7 9 13 16 1 1 10 9 9 9 13 2
6 9 1 9 9 13 2
26 16 9 13 9 14 1 9 9 7 9 9 13 7 16 9 15 9 13 9 9 14 1 9 0 13 2
15 1 9 15 0 13 16 1 1 15 9 1 15 13 13 2
20 9 0 14 9 0 7 0 7 9 1 15 13 16 13 9 14 0 9 13 2
16 10 9 0 16 1 9 0 9 13 1 15 9 7 9 13 2
41 15 9 9 7 9 13 7 2 1 9 9 1 15 7 9 15 16 1 9 13 1 9 9 13 2 9 0 16 9 15 14 13 1 1 9 9 7 9 9 13 2
17 16 15 9 9 7 9 7 9 15 16 9 9 7 9 13 13 2
14 15 1 1 9 9 9 7 9 9 7 9 9 13 2
32 15 1 9 9 7 9 3 1 15 7 1 15 9 13 2 9 15 14 13 7 15 14 13 7 9 14 1 15 15 9 13 2
14 16 15 9 9 16 1 0 9 9 15 0 13 13 2
13 15 14 16 3 1 15 7 1 15 9 13 13 2
25 16 15 9 13 16 9 9 9 13 7 9 15 7 9 2 9 2 13 2 8 8 8 8 8 2
10 3 1 9 9 14 1 9 0 13 2
21 15 1 9 3 13 2 9 7 9 9 14 9 13 2 15 14 1 9 9 13 2
3 6 9 2
7 3 15 1 10 9 13 2
6 15 16 1 15 13 2
6 16 15 9 9 13 2
15 9 1 15 9 13 16 9 1 9 9 2 9 2 13 2
12 16 9 2 9 2 1 3 9 9 15 13 2
8 16 15 3 1 9 15 13 2
27 0 9 7 9 15 7 9 15 1 9 15 13 16 1 9 7 9 9 9 13 7 1 9 7 9 13 2
9 3 1 9 9 1 10 9 13 2
9 7 10 9 7 9 14 9 13 2
20 3 1 9 15 1 15 13 16 9 9 2 9 2 14 0 9 7 9 13 2
10 15 9 14 0 1 9 15 9 13 2
19 1 9 15 13 16 9 15 15 7 9 15 7 9 9 2 9 2 13 2
14 1 9 9 15 0 1 9 1 15 9 0 14 13 2
17 16 4 1 15 9 13 2 9 1 15 0 9 1 15 4 13 2
16 7 16 13 9 13 7 1 9 9 9 1 15 14 9 13 2
17 1 9 15 13 2 15 1 15 9 13 15 16 1 15 9 13 2
4 3 6 9 2
22 1 15 9 7 9 13 2 3 13 9 13 2 1 9 0 3 1 9 0 9 13 2
20 0 13 16 15 1 1 15 15 1 9 9 13 7 9 0 15 14 0 13 2
6 3 3 13 9 13 2
3 6 9 2
44 1 9 13 7 13 9 9 13 16 10 9 1 9 7 9 1 15 9 13 7 13 16 9 15 14 0 13 13 7 3 15 14 0 13 7 1 10 9 7 9 9 15 13 2
14 15 3 9 14 1 9 9 13 16 0 7 0 13 2
20 13 16 15 15 14 1 9 13 7 9 15 14 0 13 7 9 14 9 13 2
29 9 9 1 10 9 9 9 2 9 2 1 9 1 9 9 0 13 13 16 2 8 8 8 8 8 8 8 8 2
13 16 15 1 10 9 13 2 15 16 1 15 13 2
61 16 9 15 14 13 13 7 9 13 2 10 9 14 13 0 13 2 9 15 14 13 1 9 13 2 1 15 3 13 13 2 1 12 9 9 7 9 7 9 9 1 15 9 7 9 13 2 0 13 16 10 9 7 9 3 9 1 9 9 13 2
14 15 1 9 9 0 13 9 15 7 9 1 15 13 2
33 16 9 9 2 9 2 1 9 13 15 1 10 9 13 2 1 3 15 14 9 0 2 0 1 9 7 7 0 1 9 9 13 2
14 9 9 0 0 10 9 7 9 1 9 7 9 13 2
42 9 9 9 9 9 7 9 0 9 9 1 9 9 2 9 7 9 0 7 0 9 9 9 13 7 9 0 9 14 1 9 0 1 15 9 13 7 1 9 9 13 2
47 9 9 1 9 15 9 1 9 9 9 1 9 1 9 13 7 13 2 0 9 3 9 1 1 9 9 9 1 9 9 13 7 10 9 9 0 9 1 9 0 9 15 14 16 0 13 2
27 1 9 16 0 10 9 9 13 7 10 9 7 9 2 9 1 1 9 14 1 9 9 0 9 9 13 2
34 15 13 2 16 7 15 0 7 1 9 9 9 13 13 7 9 13 16 1 9 9 9 13 9 7 9 1 15 9 0 1 9 13 2
74 9 9 3 1 9 9 0 2 0 9 3 7 3 1 9 13 7 3 1 9 1 12 9 0 7 0 9 9 7 9 0 9 9 9 13 2 1 9 16 9 0 1 9 13 2 9 9 2 16 3 0 7 7 9 0 3 0 13 16 1 9 9 0 7 9 9 1 9 9 0 1 9 13 2
43 9 9 7 9 0 13 2 1 12 9 3 1 9 0 7 1 9 0 2 9 9 1 9 3 0 16 1 9 0 7 7 1 9 0 1 9 9 7 9 0 13 13 2
43 15 13 2 9 1 9 0 3 9 9 2 9 2 9 9 2 9 1 9 7 9 7 9 1 9 7 9 2 1 12 9 0 0 1 9 1 9 1 9 9 13 13 2
53 9 9 7 9 0 1 9 1 9 1 1 9 9 9 1 9 1 9 10 9 1 9 1 9 9 7 9 13 2 15 2 1 10 9 13 16 15 1 15 1 9 10 9 1 1 9 2 3 9 9 13 13 2
21 15 13 2 9 9 9 0 7 0 13 16 1 9 9 0 1 9 15 9 13 2
36 9 9 7 9 0 1 1 9 9 1 1 9 15 16 13 2 1 9 16 9 1 9 13 2 1 3 9 9 0 9 1 9 9 13 13 2
34 15 1 1 9 0 1 9 0 9 13 2 9 7 9 1 9 15 1 9 1 9 9 9 13 7 1 9 9 7 9 9 9 13 2
59 15 13 2 1 9 7 9 9 9 1 9 1 9 13 2 9 9 15 1 0 1 12 9 12 9 1 9 0 1 12 12 9 9 13 7 16 10 9 13 16 16 9 1 9 0 7 0 9 0 13 2 9 9 7 9 15 14 13 2
40 9 9 13 2 1 9 9 9 3 9 1 9 13 16 16 9 9 13 9 9 9 14 13 2 1 10 9 13 16 9 9 13 7 9 1 9 3 0 13 2
46 9 9 7 9 0 1 9 1 15 16 9 9 1 9 9 2 9 1 9 9 7 9 9 1 9 0 9 0 1 9 13 2 13 2 9 1 9 0 1 10 9 1 9 9 13 2
31 9 9 13 2 1 10 9 2 9 9 0 1 9 15 9 13 7 10 9 2 7 0 9 9 9 9 9 14 13 13 2
58 15 13 2 9 9 9 16 3 1 15 0 3 13 2 9 9 9 9 1 1 9 0 1 9 3 0 13 7 9 15 1 9 9 7 9 1 9 1 9 12 9 12 9 9 13 16 9 13 9 3 1 1 9 15 9 13 13 2
45 9 9 7 9 0 13 2 0 9 10 9 2 9 13 9 9 1 9 9 3 9 13 7 9 0 16 9 13 16 10 9 0 13 7 3 9 1 10 9 9 15 14 9 13 2
31 9 9 9 9 9 0 9 9 13 2 10 9 7 9 0 9 13 9 7 1 0 9 0 9 9 1 9 7 9 13 2
46 15 1 9 9 7 9 9 9 0 9 0 13 2 9 0 1 9 9 4 9 0 7 0 13 13 7 1 9 9 9 13 16 9 0 4 9 0 7 0 15 14 9 7 9 13 2
59 9 9 0 9 13 2 10 9 0 1 9 9 16 1 9 0 9 9 13 4 12 9 9 7 9 0 1 9 0 7 0 13 13 7 9 1 9 0 9 0 7 9 2 9 9 0 14 16 1 9 0 7 16 1 9 0 9 13 2
19 9 9 9 13 2 9 9 0 4 9 9 9 1 9 0 9 0 13 2
31 9 9 1 9 0 7 0 0 1 9 0 1 9 0 3 1 9 0 1 9 9 0 1 9 9 0 9 9 9 13 2
16 10 9 0 7 0 1 9 0 9 1 9 1 9 13 13 2
49 1 10 9 16 9 1 9 7 9 15 1 10 9 1 9 1 9 9 3 9 0 2 9 0 7 9 9 1 9 7 9 9 7 9 13 13 1 9 9 1 9 9 9 1 9 9 13 13 2
49 1 10 9 16 3 1 9 12 9 0 0 7 0 7 1 9 12 9 1 15 9 13 9 0 0 1 9 0 2 0 2 0 7 7 9 0 7 0 7 9 0 0 7 0 1 9 13 13 2
21 10 9 9 9 9 9 2 9 9 7 9 9 9 1 0 9 1 10 9 13 2
38 1 9 9 9 9 9 7 9 0 1 15 1 9 0 3 1 9 13 2 7 9 0 1 10 9 1 9 0 9 0 3 1 9 16 9 13 13 2
25 1 9 9 0 1 9 0 1 10 9 9 2 9 0 1 9 1 9 9 7 9 0 9 13 2
13 9 0 1 9 0 9 1 9 9 9 9 13 2
29 9 9 9 9 9 13 2 1 9 9 9 0 9 2 12 12 7 12 9 9 0 1 9 0 9 9 0 13 2
26 9 9 2 13 2 10 9 1 9 12 9 9 9 0 2 1 9 9 2 9 7 9 9 13 13 2
22 7 1 10 9 12 9 12 9 9 9 9 2 9 2 9 7 9 9 1 9 13 2
52 9 9 9 9 9 13 2 1 10 9 16 12 9 0 1 9 9 2 9 2 9 2 9 2 9 7 9 1 9 13 16 1 10 9 0 12 9 1 9 9 9 7 12 9 1 9 9 0 9 0 13 2
14 1 9 10 9 2 9 9 0 9 1 12 9 13 2
20 9 9 0 9 2 1 9 9 9 1 9 0 1 9 1 9 9 9 13 2
35 9 9 9 2 13 2 10 9 1 12 9 0 10 9 1 9 1 9 2 1 9 9 0 9 13 7 1 3 1 9 0 9 13 13 2
31 15 13 2 10 9 12 0 1 9 9 15 9 0 1 9 9 0 2 0 2 9 0 7 0 7 9 0 9 13 13 2
24 9 9 13 2 10 9 1 9 9 0 9 2 9 14 1 9 7 9 0 9 9 4 13 2
22 15 13 2 3 1 9 9 7 9 9 2 9 10 9 0 1 9 9 9 4 13 2
35 1 9 15 2 9 9 0 7 0 9 0 1 9 0 1 9 9 2 9 9 7 9 9 7 9 9 9 0 1 9 3 1 9 13 2
27 1 9 9 2 9 9 1 9 12 0 1 9 1 9 13 13 16 3 1 9 9 0 1 9 1 13 2
27 9 9 12 7 12 7 0 9 9 9 9 9 7 9 9 9 9 9 1 9 9 9 9 9 0 13 2
34 1 10 9 16 9 0 1 9 10 9 0 1 1 7 1 1 9 9 13 2 9 9 9 9 1 9 1 9 10 9 9 9 13 2
30 9 9 9 9 9 9 9 9 1 10 9 13 2 1 9 9 9 2 9 7 9 7 15 1 9 9 13 13 13 2
25 15 13 2 9 1 9 9 1 9 0 0 13 16 9 9 1 9 15 1 9 1 9 15 13 2
18 9 9 9 1 9 9 9 9 1 9 9 9 15 9 9 9 13 2
17 1 9 0 9 1 9 9 0 1 10 9 0 1 9 13 13 2
27 0 9 0 9 3 1 9 7 9 15 1 9 0 2 0 7 0 9 9 9 1 9 9 9 0 13 2
28 9 9 9 9 1 10 9 13 2 9 9 9 9 12 1 12 0 1 9 12 1 9 9 1 9 0 13 2
26 9 9 9 13 2 3 1 9 9 3 12 2 12 9 1 9 1 9 9 0 3 1 9 9 13 2
35 1 9 15 9 10 9 1 9 0 1 9 9 9 9 9 12 9 9 13 7 9 0 16 1 9 0 7 0 1 10 9 9 13 13 2
42 15 9 13 2 1 9 0 9 0 7 0 9 9 7 9 9 0 9 9 1 9 9 9 9 9 9 9 13 7 3 9 9 12 9 9 1 9 9 0 13 13 2
23 10 9 1 9 9 7 9 9 9 9 0 2 9 0 2 9 2 9 7 9 0 13 2
22 9 9 0 9 9 7 9 13 2 9 9 0 9 9 2 9 9 14 1 9 13 2
33 9 9 9 3 9 1 10 9 13 2 1 9 10 9 7 9 1 9 15 4 1 9 9 3 0 10 9 0 1 9 9 13 2
19 15 0 13 2 4 9 9 1 10 9 0 7 9 1 10 9 9 13 2
39 10 9 9 12 9 9 13 7 1 9 0 1 9 0 9 9 13 7 1 9 9 9 1 9 9 9 1 9 9 15 9 13 7 1 9 9 0 13 2
33 9 0 9 1 9 0 0 13 7 9 1 9 9 2 9 2 9 2 9 0 2 9 7 9 0 13 16 1 9 0 0 13 2
28 9 0 1 9 15 9 2 9 2 9 2 9 9 13 7 3 1 9 0 9 10 9 9 1 9 13 13 2
23 1 9 9 9 0 2 9 1 9 0 1 9 9 0 9 1 9 2 9 9 9 13 2
21 9 9 0 9 9 13 2 9 0 1 0 9 13 16 1 9 9 9 13 13 2
29 9 9 13 2 1 9 10 9 0 12 9 9 0 1 9 9 0 13 16 9 0 15 1 9 9 9 9 13 2
22 15 13 2 9 0 1 9 0 1 9 9 9 7 9 1 9 0 2 13 13 13 2
10 10 9 1 9 12 9 0 4 13 2
26 9 9 9 9 13 2 12 12 7 12 12 9 1 9 0 0 9 7 9 9 0 10 9 4 13 2
36 9 9 13 2 1 0 10 9 1 1 9 12 12 9 9 0 1 9 2 12 9 0 0 0 7 12 9 10 9 1 9 0 9 4 13 2
28 15 13 2 1 9 0 1 9 1 12 9 12 2 12 7 12 12 9 12 12 9 9 0 1 9 0 13 2
40 9 13 2 1 9 12 12 9 9 1 9 1 9 0 9 9 9 1 9 1 9 10 12 9 12 9 7 1 9 1 9 10 12 9 12 9 9 4 13 2
29 15 9 9 1 9 9 0 1 9 9 14 12 9 9 13 7 13 2 9 12 9 9 10 9 0 9 0 13 2
17 9 9 9 13 2 9 9 9 9 16 0 12 7 12 9 13 2
19 9 9 1 12 0 9 9 3 13 16 1 12 9 12 12 9 9 13 2
30 9 0 9 9 9 9 9 1 9 9 0 9 0 9 9 9 9 9 9 2 3 1 9 9 9 9 1 9 13 2
43 1 10 9 16 1 9 12 9 1 9 0 1 12 9 9 7 12 9 1 9 2 9 7 9 9 9 0 13 2 12 9 1 9 7 9 0 9 9 9 9 4 13 2
54 9 9 9 0 9 0 9 0 9 9 9 9 9 9 2 1 9 10 9 13 2 9 9 1 9 9 0 14 1 1 7 1 9 9 13 7 16 1 3 9 12 9 1 9 9 7 12 9 1 9 1 9 13 2
47 15 13 2 1 9 12 9 9 9 9 9 9 9 9 2 12 9 1 9 0 7 12 9 1 9 0 1 9 9 7 9 9 1 9 9 2 9 2 9 2 9 7 9 9 4 13 2
29 9 0 1 9 9 2 9 2 9 2 9 2 9 7 9 1 9 0 9 0 9 9 9 9 9 9 9 13 2
7 0 9 9 0 9 13 2
13 3 0 9 9 0 9 0 1 9 0 4 13 2
48 1 10 9 16 9 0 9 0 13 2 9 9 7 9 0 9 15 14 1 9 9 9 9 9 4 13 7 3 1 9 0 10 9 2 9 1 9 0 9 0 9 7 7 9 9 4 13 2
26 0 9 1 9 9 9 0 13 16 9 9 2 1 9 0 0 9 9 0 9 9 9 10 9 13 2
33 0 1 9 7 9 2 1 9 9 16 1 9 0 0 13 2 9 9 9 7 9 0 2 3 12 1 9 9 9 14 9 13 2
25 9 16 1 9 9 9 9 13 2 0 13 16 9 1 9 9 2 9 9 14 0 9 9 13 2
41 1 9 0 1 3 9 12 9 9 9 9 13 16 1 10 9 9 9 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 7 9 1 9 13 2
19 9 9 0 0 9 9 7 0 9 15 13 16 1 9 9 9 13 13 2
26 0 9 10 9 12 0 16 9 9 13 2 12 9 3 1 9 0 9 9 9 9 9 13 13 13 2
14 9 2 9 14 1 9 7 9 14 1 9 9 13 2
35 9 9 9 9 1 9 9 1 9 9 13 2 9 9 7 9 7 9 0 9 7 9 9 9 0 9 9 2 1 9 0 9 0 13 2
51 9 0 1 9 15 16 9 9 1 9 0 9 1 9 13 7 9 7 9 0 1 15 1 9 1 9 9 1 13 13 9 13 1 9 0 3 9 0 0 1 9 0 9 13 9 0 1 15 9 13 2
64 9 9 0 9 14 1 9 7 9 14 1 9 16 1 9 0 9 13 9 13 7 13 16 9 7 9 16 1 9 9 9 1 0 3 1 9 0 1 9 13 13 2 13 1 9 0 7 9 0 9 9 15 14 3 9 13 7 9 9 15 14 13 13 2
12 9 1 2 9 9 2 9 0 9 0 13 2
44 9 9 1 9 2 9 1 9 9 2 0 9 9 13 2 12 7 12 9 3 1 9 9 9 2 9 9 9 0 1 9 2 9 1 9 9 2 9 9 14 1 9 13 2
46 10 9 16 1 9 0 15 1 10 9 13 2 1 1 15 13 2 16 12 9 2 9 1 9 9 2 7 9 14 4 1 15 9 13 2 7 9 15 0 12 9 14 9 13 13 2
23 9 3 1 9 10 9 9 2 15 14 9 0 7 9 9 0 1 9 0 9 13 13 2
26 1 9 0 1 9 13 16 9 2 9 1 9 9 2 9 0 1 9 9 0 9 9 9 12 13 2
52 15 1 9 13 2 9 3 0 13 2 7 9 9 0 0 13 7 4 9 1 9 9 13 16 1 9 0 9 13 7 9 9 1 15 7 9 9 0 7 9 7 9 1 9 9 7 9 9 14 13 13 2
5 9 9 2 9 2
31 9 9 0 2 3 1 12 9 9 9 1 9 0 12 9 9 9 9 9 2 9 16 1 9 9 9 13 2 9 13 2
34 1 10 9 9 1 9 12 9 3 1 9 9 0 2 9 7 9 16 1 9 12 2 12 7 12 9 9 13 2 1 9 0 13 2
44 1 0 9 10 9 2 9 9 12 9 9 15 1 9 9 9 7 9 9 1 9 0 7 0 1 9 13 16 10 12 9 0 1 9 1 9 15 1 9 1 9 1 13 2
23 9 9 16 9 9 9 0 14 1 9 13 2 1 9 0 15 9 1 10 9 13 13 2
32 9 0 1 10 9 1 12 9 9 1 9 9 1 9 0 7 12 9 1 9 9 7 9 9 1 9 0 7 0 9 13 2
15 9 9 1 10 9 12 9 9 7 12 9 9 13 13 2
26 9 12 0 0 9 9 9 0 9 9 2 3 1 9 9 9 1 9 9 2 9 7 9 9 13 2
20 1 9 10 9 9 9 9 7 9 9 1 9 1 9 15 9 9 0 13 2
22 1 9 9 9 9 9 9 9 9 7 9 9 1 9 0 12 1 12 1 9 13 2
24 9 9 1 9 12 1 9 9 9 7 9 9 1 9 12 1 9 9 1 10 9 9 13 2
27 1 9 9 9 9 2 9 9 0 13 1 9 9 1 9 12 1 12 1 1 9 9 9 1 9 13 2
37 9 0 7 0 10 9 1 9 12 1 12 1 9 9 9 9 13 7 1 9 1 9 12 1 12 9 1 9 9 2 9 1 9 9 13 13 2
41 1 9 9 9 9 9 10 12 9 15 14 9 13 7 12 9 9 9 9 9 1 9 9 1 9 13 7 1 10 9 9 9 9 14 1 9 0 15 0 13 2
18 9 10 9 14 9 9 2 1 9 9 9 7 9 9 1 9 13 2
18 9 9 1 9 9 9 1 9 12 1 12 1 9 9 9 0 13 2
34 1 10 9 9 9 1 9 12 1 9 9 9 9 13 7 9 9 1 9 12 7 9 9 1 9 12 9 9 9 14 1 9 13 2
33 1 9 15 16 9 9 7 9 9 10 12 1 9 9 13 2 0 12 9 0 13 7 1 10 9 9 9 1 9 0 9 13 2
12 1 9 0 9 9 1 9 9 9 4 13 2
16 9 9 9 9 9 7 9 1 9 1 9 0 9 4 13 2
4 9 2 9 2
44 9 13 9 12 12 9 0 3 1 0 9 2 9 0 9 2 1 9 1 9 0 0 0 1 10 10 9 1 9 0 9 0 0 13 7 1 9 9 1 15 1 9 13 2
21 15 0 9 0 1 9 1 9 9 1 9 13 16 1 9 9 0 9 0 13 2
32 12 9 1 9 9 3 1 9 9 9 0 10 9 1 9 9 9 13 16 9 0 0 13 7 1 9 0 9 15 9 13 2
20 9 12 0 1 9 9 0 12 9 1 9 9 1 13 7 3 9 9 13 2
53 1 9 9 12 1 9 9 2 3 1 9 0 9 7 9 15 1 9 9 2 1 9 12 9 12 9 9 0 1 10 9 9 13 2 1 9 7 1 10 9 0 3 12 9 9 0 1 10 9 9 13 13 2
18 9 9 9 10 9 9 12 9 14 9 13 16 9 9 9 0 13 2
25 9 9 0 9 13 13 16 9 0 1 9 0 1 9 9 9 0 13 9 15 14 1 9 13 2
51 10 9 3 1 12 9 9 1 9 16 1 9 0 0 1 9 9 0 7 9 0 13 2 9 13 16 9 9 0 7 9 1 9 9 9 13 9 14 1 9 0 9 13 7 1 9 9 15 9 13 2
23 10 9 9 13 13 16 3 9 9 0 0 13 2 9 9 0 9 0 1 9 15 13 2
26 9 0 9 13 9 0 0 1 9 9 7 9 9 0 9 9 1 9 9 14 1 12 9 9 13 2
34 9 9 9 13 13 16 9 0 0 1 9 7 9 1 9 0 9 0 13 7 9 0 9 1 10 9 2 9 9 9 14 9 13 2
23 12 1 9 9 9 9 0 9 13 2 16 1 9 9 9 9 9 9 0 9 9 13 2
16 9 13 10 9 1 9 0 9 1 9 9 0 9 0 13 2
4 9 2 9 2
21 9 9 9 9 9 9 0 7 9 0 10 9 14 1 9 9 1 9 0 13 2
25 9 0 9 9 9 3 1 9 9 9 9 13 16 9 7 9 0 1 9 9 9 9 9 13 2
34 9 9 2 9 0 9 14 1 9 1 9 9 0 7 9 1 15 1 1 9 9 1 9 9 15 2 12 1 12 2 9 13 13 2
29 9 9 9 12 0 2 12 9 1 9 9 9 9 13 7 12 9 9 9 14 1 9 0 10 9 1 9 13 2
5 9 0 2 9 2
32 9 9 2 9 9 0 9 1 9 9 1 9 9 9 9 1 9 9 9 0 2 9 9 1 9 9 1 9 9 9 13 2
28 1 9 9 9 2 9 9 13 2 16 9 1 1 9 9 0 9 3 9 13 2 1 9 15 9 4 13 2
32 1 9 16 9 9 1 9 9 9 13 2 13 13 2 9 9 1 9 9 0 2 1 9 0 9 9 1 9 15 9 13 2
4 9 2 9 2
38 9 0 9 9 13 2 9 9 0 9 0 13 2 3 9 0 7 9 15 14 9 13 16 9 0 1 9 0 9 0 12 9 0 2 9 4 13 2
28 10 9 0 9 13 2 7 10 9 0 13 9 1 9 9 9 9 16 0 1 13 9 12 9 13 2 13 2
49 10 9 0 0 13 7 9 9 9 9 1 9 9 12 2 1 9 16 10 9 1 9 9 0 9 9 9 9 13 2 1 9 16 1 9 9 9 1 12 0 9 9 0 9 9 13 2 13 2
44 3 1 12 9 9 7 0 0 1 12 12 9 9 1 9 1 1 10 9 2 9 9 0 0 9 3 9 15 14 9 13 7 3 9 9 1 9 0 16 1 9 13 13 2
6 9 2 9 0 9 2
29 3 1 12 9 0 9 1 9 1 9 2 10 9 0 1 9 9 9 9 13 16 4 1 12 9 9 9 13 2
23 10 9 12 1 12 9 13 16 9 1 9 1 9 12 0 1 9 9 1 9 13 13 2
14 9 0 0 9 9 13 16 1 9 9 9 4 13 2
30 9 0 12 9 12 9 13 16 3 1 3 9 1 9 15 1 9 9 2 1 3 9 1 12 9 9 9 4 13 2
18 10 9 9 3 1 9 0 9 13 7 9 3 1 9 15 4 13 2
6 9 2 9 0 9 2
35 9 9 9 9 0 2 9 9 0 1 9 1 9 1 9 12 2 1 9 7 9 9 1 9 1 9 0 9 9 3 13 2 0 13 2
27 1 9 9 9 2 10 9 0 0 0 1 9 7 1 9 9 0 9 9 13 13 2 15 9 14 13 2
14 15 16 3 9 9 9 13 2 1 9 9 0 13 2
23 9 9 9 9 13 1 12 9 9 13 16 1 1 9 7 9 9 15 1 9 9 13 2
34 9 9 9 12 0 3 1 15 7 1 9 12 9 9 9 0 14 1 9 9 9 9 13 2 1 12 9 9 0 7 3 0 13 2
4 9 2 9 2
13 9 9 9 0 1 9 2 9 0 3 9 13 2
38 9 0 9 0 9 1 9 9 2 9 9 9 13 2 1 12 9 0 9 12 0 2 12 9 9 1 9 9 1 9 0 9 15 14 1 9 13 2
30 1 1 10 9 2 9 9 9 0 1 12 9 0 9 12 0 1 9 1 9 0 1 9 0 2 12 9 0 13 2
48 1 9 0 0 2 12 12 7 12 9 2 9 9 9 0 2 1 9 9 2 9 7 0 9 0 0 2 1 9 13 16 1 9 1 9 10 9 1 9 12 2 12 2 12 9 0 13 2
68 9 9 9 16 3 1 10 9 15 1 9 9 9 9 0 9 9 2 9 9 2 0 13 13 7 1 9 9 9 1 3 9 1 9 13 13 9 9 1 9 0 1 9 0 10 9 1 9 7 9 9 0 15 9 9 14 1 9 13 1 9 9 9 9 14 0 13 2
48 1 10 9 16 1 9 9 9 0 13 2 9 9 9 1 12 9 1 9 9 9 1 9 9 13 7 12 9 0 10 9 14 1 9 15 13 16 9 15 14 1 9 9 10 9 9 13 2
22 9 9 9 1 9 12 1 9 9 7 12 7 12 1 9 9 9 9 1 9 13 2
15 10 9 14 9 9 1 9 9 9 7 9 9 9 13 2
55 9 0 3 1 12 9 1 12 9 1 0 9 0 1 9 9 7 0 9 7 9 1 9 0 9 9 13 2 1 0 9 16 9 9 9 14 13 7 9 0 13 2 9 1 9 9 4 13 7 9 1 9 9 13 2
27 7 16 9 7 9 10 12 13 2 9 4 9 14 1 3 12 9 13 16 4 1 9 9 0 9 13 2
13 7 16 10 12 9 13 9 9 3 9 4 13 2
9 9 0 9 9 0 9 9 13 2
22 9 9 9 0 9 0 0 9 1 0 9 9 9 0 9 9 9 14 1 9 13 2
29 9 9 9 9 12 0 9 9 9 1 9 14 1 9 12 2 12 2 12 9 9 13 7 1 9 0 9 13 2
25 9 9 9 0 7 9 9 10 9 0 1 12 9 7 12 9 9 1 9 0 7 0 9 13 2
26 1 9 0 7 1 9 9 0 10 9 2 9 9 0 2 0 7 9 1 9 0 1 0 9 13 2
39 9 9 9 9 7 9 9 9 9 0 9 9 1 9 9 1 9 0 9 9 9 2 3 1 9 9 9 2 9 14 1 9 9 9 9 9 9 13 2
43 1 10 9 16 9 12 9 9 0 1 9 9 9 13 2 9 9 9 9 9 9 9 16 1 9 12 9 9 1 0 9 9 9 0 1 9 0 4 13 2 9 13 2
23 9 9 9 9 1 12 9 0 7 0 1 1 9 9 9 1 9 12 1 12 9 13 2
30 16 15 9 9 9 14 16 1 10 9 0 13 9 9 0 1 9 10 9 1 9 9 0 0 9 0 0 9 13 2
20 15 1 9 1 9 9 9 13 16 9 9 9 9 9 1 9 0 9 13 2
37 1 9 13 9 3 0 9 1 9 9 1 1 9 9 0 1 9 0 9 13 7 15 0 13 16 9 0 9 0 9 9 0 15 14 13 13 2
49 1 9 7 9 9 3 9 13 16 9 0 7 0 13 13 7 3 1 15 1 9 9 7 9 7 9 7 9 7 2 9 13 13 7 3 1 10 9 9 1 9 1 9 0 7 0 9 13 2
13 3 9 9 10 9 14 1 3 9 4 9 13 2
23 7 3 1 9 9 9 1 9 9 9 16 9 0 9 0 1 9 14 1 9 1 13 2
13 16 9 9 14 4 1 9 9 9 9 9 13 2
34 16 9 9 0 14 4 9 1 9 9 9 0 13 1 0 15 16 9 9 9 3 1 12 9 1 9 1 9 1 9 9 13 13 2
10 16 9 13 9 0 1 9 9 13 2
12 16 9 3 1 9 9 9 0 9 13 13 2
9 16 9 13 9 9 14 2 2 2
18 1 9 13 9 9 9 9 14 1 9 9 4 1 12 9 9 13 2
38 9 2 1 9 9 9 9 1 9 0 15 1 9 9 15 1 10 9 13 16 9 9 7 9 7 9 0 1 15 13 16 1 1 9 0 9 13 2
27 9 0 7 0 9 9 1 9 9 0 15 13 13 2 12 1 9 0 1 9 9 9 9 9 9 13 2
23 0 9 9 9 9 14 0 13 7 1 1 9 12 9 7 7 0 1 15 9 9 13 2
29 10 9 16 9 13 16 16 9 9 9 0 9 1 9 9 14 0 13 9 9 0 1 9 0 4 13 7 0 2
76 10 9 0 13 1 9 9 0 9 1 9 9 2 1 9 9 2 9 9 0 3 1 12 9 9 4 0 13 2 1 9 7 9 0 1 9 1 9 9 9 9 9 7 15 16 1 9 12 9 9 3 3 9 1 12 9 0 3 13 9 13 16 16 9 0 9 0 13 2 9 9 1 9 13 13 2
24 9 9 9 9 9 13 1 9 16 0 9 1 9 9 9 13 9 4 1 9 0 0 13 2
49 0 1 9 13 1 9 16 9 15 0 13 9 9 1 9 0 0 13 2 1 9 7 9 0 9 9 7 9 9 12 9 9 0 9 9 0 13 7 4 1 9 0 9 9 9 0 0 13 2
24 9 9 1 9 12 9 9 9 13 13 2 12 9 1 9 9 9 9 1 9 13 13 13 2
20 12 9 16 1 9 9 0 2 0 9 9 2 9 9 7 0 1 9 13 2
26 9 10 0 9 2 16 1 9 0 9 9 7 1 0 2 1 9 9 9 7 9 0 1 9 13 2
96 7 1 10 9 2 9 9 9 1 9 9 0 7 0 16 1 15 9 13 2 3 9 0 7 0 13 16 3 13 15 14 1 9 0 16 1 9 13 2 9 7 9 13 2 0 9 14 4 15 13 16 9 9 3 15 9 0 2 0 0 2 9 0 2 0 1 9 7 0 7 0 13 16 1 9 7 9 0 9 13 7 4 9 9 0 7 9 0 0 2 9 7 9 15 13 2
12 15 0 7 0 1 3 9 10 9 0 13 2
12 9 0 1 0 9 7 0 9 9 9 13 2
28 15 9 13 16 9 1 12 9 9 9 7 9 9 13 7 1 9 0 7 1 9 7 9 0 9 0 13 2
71 16 9 2 9 0 1 15 13 7 7 1 9 2 1 9 0 1 9 9 9 0 4 13 2 1 9 0 2 9 9 12 9 13 16 12 2 9 7 9 13 2 0 2 9 7 9 0 13 7 9 0 15 2 9 7 9 9 13 16 1 9 9 7 9 0 9 0 9 13 13 2
44 1 0 2 9 9 2 9 3 0 0 14 1 15 0 13 7 15 2 15 7 9 9 3 9 9 0 9 13 2 7 9 7 9 16 3 13 9 9 0 14 1 9 13 2
40 10 9 7 4 0 9 1 9 13 2 4 1 9 9 9 1 15 2 16 13 2 3 7 10 12 0 1 9 13 16 15 14 1 9 1 9 0 13 13 2
124 9 2 15 9 10 9 7 9 0 9 2 7 7 9 2 9 7 9 15 2 13 7 3 7 9 13 16 9 1 9 9 9 7 1 9 9 7 9 0 9 13 7 9 13 16 9 0 2 9 0 14 0 13 7 9 1 9 9 0 7 9 9 9 7 9 13 2 1 9 0 7 0 7 7 0 9 9 13 7 3 9 16 9 14 9 0 7 1 9 9 1 9 0 1 9 9 13 16 4 1 9 7 9 7 1 1 9 9 9 0 0 7 0 0 7 0 13 2 1 9 9 13 2 2
11 12 9 9 9 1 9 9 0 0 13 2
6 9 2 9 0 9 2
29 12 9 9 9 0 9 9 16 12 7 12 9 1 15 9 13 2 9 9 1 9 9 9 0 1 9 0 13 2
23 1 9 9 9 9 9 10 9 0 9 0 13 13 7 12 1 9 15 3 9 0 13 2
21 10 9 1 9 1 9 9 13 16 0 9 0 13 7 1 9 9 9 0 13 2
37 3 1 9 2 10 9 1 9 12 9 1 9 9 9 13 16 9 15 14 9 13 7 9 1 15 14 16 3 13 16 1 9 9 0 9 13 2
12 12 9 1 9 10 9 1 10 9 0 13 2
11 9 9 1 9 9 2 1 9 9 13 2
4 9 2 9 2
24 9 9 9 1 9 0 9 2 9 9 12 9 9 14 1 9 0 12 12 9 2 9 13 2
27 9 9 9 9 9 10 9 1 9 1 9 13 2 12 0 10 9 14 1 9 1 9 1 9 0 13 2
17 10 12 9 16 9 13 2 10 9 14 1 9 13 2 9 13 2
4 9 2 9 2
41 12 9 0 9 9 1 9 9 1 9 0 9 2 12 9 7 12 9 1 9 9 15 14 1 9 13 7 0 9 3 9 15 14 0 13 1 9 1 15 13 2
63 1 9 9 9 1 9 9 1 9 2 0 1 12 9 3 1 9 10 9 16 9 15 1 9 9 0 13 7 13 13 16 0 1 12 9 9 13 2 3 3 1 9 1 9 0 9 12 0 1 9 1 9 0 14 1 9 12 9 1 9 0 13 2
5 15 3 0 13 2
30 12 9 9 1 9 9 13 2 9 1 9 9 9 9 9 9 3 13 7 15 14 1 3 9 9 1 9 9 13 2
18 1 9 10 9 2 9 0 0 13 7 9 15 16 0 7 0 13 2
32 10 9 16 12 9 0 0 1 15 9 13 2 3 1 9 16 12 9 7 9 9 13 2 0 9 1 9 15 14 0 13 2
30 3 9 9 0 13 2 7 9 9 9 1 15 13 16 15 0 13 9 1 12 1 9 9 10 9 9 9 13 13 2
32 1 9 9 9 12 9 9 9 13 16 10 9 9 12 1 9 13 7 3 1 9 1 9 9 1 9 9 7 9 13 13 2
11 9 0 12 1 9 0 9 14 9 13 2
4 9 2 9 2
15 9 1 9 12 2 12 9 9 9 1 9 9 14 13 2
23 1 9 9 9 9 2 9 0 1 9 9 9 13 2 7 3 9 9 0 9 13 13 2
31 9 9 9 13 13 2 9 10 9 12 2 12 9 1 9 9 7 9 15 1 1 9 12 0 9 0 9 9 13 13 2
13 10 9 1 12 0 9 0 9 9 9 9 13 2
4 9 0 9 2
25 1 9 9 1 9 12 9 9 0 9 2 12 9 1 9 9 9 0 7 12 9 16 0 13 2
46 1 9 9 0 9 2 9 9 9 0 9 13 16 3 1 9 9 12 9 9 9 7 9 2 12 1 9 9 9 1 9 1 9 9 9 9 13 7 12 1 15 14 1 9 13 2
24 12 1 9 10 9 16 16 1 9 9 3 0 13 13 2 1 9 0 1 9 0 9 13 2
19 9 9 9 9 9 1 9 0 9 9 0 9 1 9 9 0 9 13 2
24 1 9 9 2 9 9 0 9 13 16 9 3 4 9 0 0 7 9 3 0 0 9 13 2
38 1 9 7 9 9 13 1 9 9 0 3 1 9 13 2 9 9 9 0 9 9 14 13 7 9 0 9 7 9 9 9 9 9 9 14 9 13 2
27 9 1 9 1 9 9 9 13 2 9 16 16 1 9 1 9 9 9 13 2 4 1 10 9 9 13 2
19 9 1 9 9 9 9 13 2 10 9 3 0 7 0 1 9 9 13 2
25 9 9 13 9 0 13 7 1 15 16 9 13 1 9 1 9 15 9 13 2 0 9 13 13 2
25 9 0 13 2 3 9 9 16 9 13 9 15 0 13 3 0 2 9 9 9 0 13 1 0 2
14 7 1 10 9 9 15 9 9 0 14 9 13 13 2
21 12 9 9 9 1 1 9 0 10 9 7 0 9 9 9 9 9 9 9 13 2
22 9 0 9 0 9 0 9 2 1 1 9 9 2 9 9 7 9 0 9 15 13 2
31 7 9 1 9 10 9 13 2 9 9 9 1 9 7 9 0 9 0 13 2 9 16 3 1 9 9 9 9 13 13 2
11 1 9 9 9 9 9 12 9 9 13 2
4 9 2 9 2
21 9 1 9 1 9 9 9 13 2 9 0 9 1 9 0 7 0 9 9 13 2
34 9 9 9 1 9 0 15 13 2 12 9 9 1 9 0 9 13 16 9 15 14 1 9 0 2 3 9 1 1 9 15 9 13 2
18 9 9 13 9 9 7 9 9 1 9 0 2 3 9 1 15 13 2
34 1 9 9 0 16 1 9 0 9 9 13 9 9 13 1 9 9 0 1 9 7 9 1 9 0 9 2 0 9 15 3 0 13 2
27 9 0 1 10 9 1 3 0 13 16 9 0 1 9 0 7 15 9 1 9 9 0 13 2 9 13 2
30 1 9 12 0 12 9 0 1 9 3 1 9 0 9 12 0 15 1 9 9 0 1 9 9 13 7 3 9 13 2
16 9 0 9 1 9 1 9 9 0 9 12 0 15 9 13 2
36 1 9 0 12 9 0 1 9 9 2 9 0 14 3 1 9 9 0 13 2 7 1 9 0 7 0 0 1 15 1 9 9 15 9 13 2
26 1 9 0 9 1 9 0 3 9 2 9 2 7 9 2 9 0 9 1 9 15 14 0 9 13 2
18 1 9 7 9 9 0 9 1 9 15 3 1 9 0 9 0 13 2
27 1 10 9 3 9 16 3 1 9 9 9 13 7 9 9 1 9 0 13 10 9 14 16 0 9 13 2
44 9 1 9 9 9 13 2 9 16 1 9 9 1 9 0 1 9 0 9 13 13 2 1 9 9 1 9 0 3 9 7 9 1 9 0 0 13 7 1 15 9 0 13 2
76 1 9 0 7 9 0 9 15 2 1 9 0 1 9 0 7 0 2 1 9 16 9 9 7 9 9 15 13 2 1 9 9 15 2 1 10 9 0 16 1 9 9 9 9 13 13 7 1 1 9 9 16 1 9 7 9 0 1 1 9 9 9 13 7 1 3 13 2 9 9 9 1 9 0 13 2
2 3 2
13 13 9 3 9 1 13 7 3 9 7 9 13 2
46 3 10 9 14 1 9 0 13 2 16 3 1 9 7 9 1 9 7 9 15 2 1 9 0 2 9 0 9 9 16 9 9 7 9 14 13 7 3 1 9 0 13 1 9 13 2
89 3 15 9 15 2 15 9 15 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 7 9 7 0 12 9 1 15 2 0 1 9 9 0 9 0 7 0 2 0 1 9 1 15 9 9 9 7 7 9 9 0 2 1 9 1 9 0 9 7 9 7 9 7 9 0 0 2 9 2 8 9 7 9 7 9 9 7 9 2 9 13 2
33 9 0 13 16 9 9 7 9 1 9 7 1 9 9 9 15 14 13 2 16 9 15 14 1 9 0 1 9 1 15 13 13 2
31 9 3 1 15 7 9 0 1 9 13 2 9 9 14 0 13 7 1 9 0 7 0 15 9 1 9 0 15 1 13 2
16 1 10 9 9 9 7 9 1 9 15 1 12 9 0 13 2
13 1 9 9 7 9 7 1 9 9 7 9 13 2
4 9 2 9 2
17 3 1 9 0 0 2 9 9 0 1 9 7 9 12 9 13 2
18 9 9 9 9 9 13 2 12 9 0 1 9 9 9 9 13 13 2
46 9 9 0 9 13 16 1 9 7 9 9 9 1 9 1 15 9 13 7 10 9 0 9 13 13 16 9 0 0 1 9 10 9 1 12 9 1 9 1 9 1 10 9 9 13 2
38 9 0 2 9 2 9 15 13 2 13 16 12 9 3 9 0 7 0 14 1 0 1 9 0 9 0 13 7 0 1 12 12 9 9 1 9 13 2
38 9 0 16 1 9 12 9 0 1 9 9 4 13 1 9 9 1 9 9 1 9 9 13 4 13 16 9 1 9 0 15 14 1 9 15 9 13 2
42 9 9 0 15 13 16 10 9 9 2 9 2 14 16 1 9 0 9 0 2 9 9 2 9 13 2 9 13 7 1 9 0 9 9 2 9 0 9 15 14 13 2
30 9 9 12 1 9 9 9 9 1 9 9 0 9 13 2 9 3 9 9 2 9 15 13 2 1 9 0 9 13 2
30 9 9 0 9 15 13 16 9 9 9 14 1 9 9 1 0 9 9 9 13 16 3 0 13 7 3 1 9 13 2
18 9 0 2 10 9 9 0 9 14 16 9 9 13 13 2 0 13 2
29 16 9 1 10 9 9 13 2 4 9 15 14 1 9 0 9 13 7 1 9 0 1 9 9 1 9 15 13 2
10 0 9 9 9 0 1 12 9 13 2
4 9 2 9 2
21 0 9 9 9 2 9 9 1 9 0 1 12 12 9 0 1 9 9 0 13 2
22 9 9 9 9 9 13 2 9 10 9 13 9 0 14 1 9 9 9 1 9 13 2
31 9 9 9 7 9 9 9 10 9 9 9 1 10 9 1 15 13 7 1 9 9 0 9 9 0 14 1 9 1 13 2
22 10 9 1 9 9 9 0 15 1 9 9 9 0 1 9 9 12 9 14 9 13 2
21 9 10 9 0 12 9 1 9 13 7 0 1 12 12 9 9 1 9 13 13 2
16 9 9 9 9 9 9 9 0 1 10 9 14 0 9 13 2
34 1 9 12 12 7 12 9 1 10 9 9 13 7 1 10 9 9 12 9 3 14 16 0 1 12 12 7 12 9 0 13 2 13 2
4 9 2 9 2
43 12 9 9 0 9 16 1 9 9 9 9 13 2 9 9 9 13 16 3 1 1 12 12 9 1 9 0 13 7 1 9 0 9 9 0 1 0 9 9 1 9 13 2
29 9 10 9 9 16 1 9 9 0 9 0 0 13 2 0 13 2 9 9 1 9 0 1 12 2 12 9 13 2
21 9 9 10 9 1 9 0 0 13 7 1 0 1 9 9 0 9 9 13 13 2
20 9 12 9 0 1 9 15 13 16 9 2 3 1 12 9 0 0 9 13 2
16 9 13 1 10 9 9 13 7 9 0 1 9 9 0 13 2
17 9 0 9 9 1 9 0 7 9 9 0 1 0 1 9 13 2
28 7 1 10 9 9 13 13 16 9 0 9 9 13 1 9 12 1 9 15 16 3 9 9 9 13 9 13 2
36 9 9 9 9 0 9 13 2 1 9 0 7 9 0 2 15 9 9 13 2 16 9 7 9 0 1 9 0 9 9 13 2 7 0 13 2
12 15 13 2 15 1 12 9 0 0 9 13 2
15 15 1 9 0 3 13 1 9 9 9 0 1 9 13 2
35 7 1 10 9 1 9 1 9 9 7 9 9 13 13 16 9 15 1 9 0 1 9 0 9 13 7 9 13 9 14 1 15 9 13 2
6 9 2 9 0 9 2
29 9 0 9 1 9 9 16 12 9 9 15 14 1 9 13 2 0 13 7 10 9 0 9 0 9 9 0 13 2
44 1 9 9 1 9 2 9 9 9 0 9 1 1 9 9 1 9 9 1 9 9 9 2 9 2 9 2 9 2 9 0 7 9 2 1 9 12 9 9 7 9 13 13 2
37 1 9 0 13 13 2 10 9 0 1 15 13 16 0 9 1 9 3 1 9 9 9 0 1 10 9 0 1 9 9 0 1 1 9 0 13 2
58 1 9 0 1 10 9 16 1 9 9 9 9 0 13 13 2 1 15 7 10 9 0 1 9 9 9 9 9 13 2 10 9 4 1 10 9 1 9 0 9 0 1 1 9 9 13 7 9 0 1 9 9 0 1 9 9 13 2
33 9 9 0 16 9 0 15 14 1 9 0 9 9 13 2 9 9 1 10 9 3 9 2 9 2 9 7 9 7 3 9 13 2
18 1 9 0 1 10 9 9 9 1 9 0 1 1 9 9 13 13 2
26 1 9 15 1 9 9 1 15 13 16 9 9 1 9 16 3 1 9 9 0 9 13 2 0 13 2
20 9 9 0 0 1 9 1 9 0 1 1 9 2 1 15 1 9 0 13 2
4 9 0 13 2
4 9 2 9 2
12 9 0 9 9 14 1 9 9 0 9 13 2
51 9 0 9 9 9 9 2 1 9 0 15 16 3 0 13 2 9 13 13 2 9 9 9 1 9 9 0 15 13 16 9 0 9 13 10 9 16 1 9 9 9 9 9 13 2 1 9 3 9 13 2
51 9 9 0 9 9 9 9 9 13 2 9 9 1 15 10 9 14 1 9 13 13 16 1 9 0 7 0 1 10 9 9 13 16 9 9 1 9 2 1 9 9 1 9 13 16 1 1 9 9 13 2
27 15 13 2 3 9 1 9 13 1 12 9 0 2 1 1 9 9 1 10 9 16 1 10 9 0 13 2
30 10 9 1 1 9 2 9 9 2 9 16 1 9 9 0 7 0 1 15 9 13 14 16 1 9 9 0 9 13 2
10 9 9 9 9 0 0 1 9 13 2
6 9 2 9 0 9 2
31 9 0 16 1 9 9 7 9 9 0 3 9 9 13 2 13 1 9 0 16 3 1 9 0 1 9 9 13 2 13 2
36 1 9 9 9 2 1 9 0 1 9 9 0 9 9 2 10 9 16 1 9 9 0 0 13 2 16 1 9 9 9 7 9 16 9 13 2
15 7 9 0 9 0 1 10 9 14 1 9 15 0 13 2
14 10 9 9 9 1 9 9 12 16 0 9 13 13 2
16 9 10 9 1 9 12 9 1 9 1 9 9 9 13 13 2
41 9 10 9 13 2 9 9 9 2 12 1 1 9 1 9 0 1 10 9 9 13 2 1 9 7 1 9 9 0 13 1 9 0 1 9 0 1 9 13 13 2
31 12 1 9 10 9 13 2 9 9 0 9 9 9 1 9 9 13 7 9 9 12 9 9 9 1 9 0 1 9 13 2
9 9 0 9 9 9 14 9 13 2
4 9 2 9 2
17 9 9 9 9 16 1 0 1 9 9 13 2 3 9 4 13 2
28 1 9 9 0 0 1 9 1 9 2 0 1 9 16 3 1 10 9 1 9 7 9 0 9 9 9 13 2
28 10 9 2 16 1 9 1 9 7 9 9 9 13 7 7 9 9 13 9 9 7 9 0 14 1 1 13 2
37 9 0 16 9 0 1 15 1 9 9 13 1 9 9 13 16 1 9 1 9 9 9 0 0 13 7 9 9 9 1 9 9 14 1 9 13 2
19 1 10 9 2 9 1 9 0 1 9 13 7 9 15 14 9 4 13 2
25 1 9 0 9 12 12 9 1 9 1 9 1 9 9 9 1 9 9 0 9 1 9 9 13 2
24 9 13 16 1 9 12 0 9 9 12 9 9 0 1 9 2 9 9 1 9 14 1 13 2
2 9 2
18 9 16 9 0 1 9 9 0 13 2 9 9 14 9 0 9 13 2
13 16 4 9 9 15 1 9 14 16 9 0 13 2
33 9 9 1 9 7 9 9 7 9 0 9 0 1 9 0 1 9 0 9 9 13 2 7 1 13 16 1 9 0 9 0 13 2
44 9 9 9 0 9 1 9 9 13 2 9 16 1 12 9 0 9 9 0 9 7 9 0 13 3 0 1 9 9 0 0 9 9 13 7 9 15 1 9 9 9 0 13 2
34 9 9 13 16 1 9 0 9 9 2 9 0 1 9 9 0 9 13 7 9 9 9 9 9 7 9 0 9 1 9 10 9 13 2
25 9 9 7 9 0 9 9 9 1 9 14 9 13 2 16 9 0 1 9 1 9 9 9 13 2
36 9 16 3 1 9 9 9 0 13 7 9 9 0 13 2 1 9 9 0 0 9 7 9 13 7 9 15 9 9 15 1 9 9 9 13 2
11 1 12 9 0 9 0 9 1 9 13 2
47 9 2 15 13 16 1 9 9 9 2 2 9 2 9 9 2 9 2 9 2 7 9 13 2 7 9 3 0 13 2 7 7 1 9 0 9 2 9 0 9 14 1 15 3 9 13 2
48 1 9 9 2 1 9 1 9 7 9 2 9 9 0 13 13 2 7 0 9 9 1 15 9 13 13 2 1 9 9 13 2 13 9 0 1 9 7 9 0 2 1 12 12 9 7 9 2
9 0 3 7 9 9 3 13 0 2
17 9 0 13 9 1 9 9 2 10 9 13 16 13 3 9 0 2
18 7 10 9 13 16 13 3 9 0 2 3 13 9 7 3 13 0 2
9 3 13 9 2 9 1 9 9 2
32 9 0 15 13 16 9 9 9 16 2 1 9 0 13 2 10 0 9 0 9 2 13 3 9 9 2 1 9 9 9 9 2
13 1 9 13 12 12 9 2 1 9 9 9 9 2
15 3 10 9 9 13 1 9 2 1 15 9 9 13 0 2
33 1 15 3 13 16 15 0 13 2 16 9 9 15 13 10 10 9 16 13 9 7 9 7 9 2 3 1 9 1 15 13 9 2
30 16 12 0 14 9 9 9 13 0 1 12 0 7 12 0 2 9 10 9 0 1 13 1 12 9 2 9 12 9 2
43 10 9 14 4 9 9 13 2 16 3 9 1 1 10 12 9 0 1 9 1 9 10 9 0 13 7 3 9 1 9 9 2 1 9 0 7 9 0 0 9 13 13 2
31 9 9 1 9 10 9 9 13 2 7 0 13 13 16 1 9 10 9 9 2 9 9 1 9 15 2 9 2 9 13 2
7 9 9 3 9 4 13 2
29 15 0 13 16 10 9 1 9 9 13 16 1 9 2 9 7 9 15 2 9 0 9 9 14 1 1 9 13 2
27 9 16 1 9 3 1 9 2 1 9 9 2 1 15 0 13 13 2 7 9 1 9 10 9 9 13 2
29 3 9 1 9 9 7 9 13 9 13 16 3 10 9 2 3 3 1 12 9 0 1 0 1 9 9 13 13 2
16 9 13 2 16 9 3 9 13 0 2 9 0 3 9 0 2
10 10 9 7 10 9 14 3 9 13 2
60 9 16 9 14 1 9 4 13 7 9 9 4 13 2 3 12 9 12 12 9 14 0 13 2 7 1 15 9 7 9 7 9 16 1 9 1 15 9 13 13 2 7 7 10 15 16 1 9 7 9 9 0 13 2 1 9 13 4 13 2
48 16 1 15 4 13 9 16 9 15 1 9 9 13 2 3 9 7 9 7 9 7 9 2 1 9 0 7 0 1 9 9 7 9 7 9 2 9 9 1 9 10 9 0 7 0 9 13 2
32 9 7 9 7 9 7 9 2 9 14 1 9 16 15 3 1 9 9 13 1 13 7 9 15 14 1 9 9 0 0 13 2
19 9 9 1 9 9 1 10 9 0 13 2 16 1 9 9 15 9 13 2
10 9 9 10 9 9 7 9 9 13 2
20 1 9 9 7 9 7 9 7 9 9 7 9 9 2 9 15 14 9 13 2
60 9 16 0 13 1 9 9 1 9 13 2 4 9 1 9 9 13 2 1 10 9 7 9 2 9 9 1 9 9 7 9 9 2 1 13 1 9 9 0 1 9 2 3 9 9 2 15 1 9 9 13 2 7 3 1 12 9 9 13 2
8 9 9 0 1 15 0 13 2
35 9 7 9 1 9 2 9 1 9 9 2 7 9 7 0 1 9 2 7 15 10 9 13 16 9 0 1 9 0 9 15 9 13 13 2
11 1 9 9 9 4 9 1 9 9 13 2
20 4 1 0 9 9 13 16 9 1 9 0 15 0 13 7 9 1 9 13 2
49 9 0 9 2 9 7 9 9 4 13 2 1 9 15 0 13 16 0 9 0 1 9 7 9 7 9 9 1 9 0 9 13 2 1 9 9 1 9 0 7 9 16 1 10 9 0 13 13 2
59 1 9 2 9 4 13 1 9 9 2 1 9 9 2 7 9 13 16 1 10 9 10 9 0 2 10 9 16 13 13 2 16 1 9 9 15 7 7 1 9 9 2 13 13 2 7 7 9 15 9 13 16 0 1 3 9 0 13 2
13 10 9 7 10 9 2 3 0 1 9 9 13 2
25 16 1 9 9 0 9 13 16 1 9 9 1 15 4 10 9 7 10 9 0 15 14 1 13 2
22 7 3 10 9 7 10 9 9 15 1 9 13 16 4 1 9 0 9 0 9 13 2
14 4 10 9 1 9 7 9 7 9 1 15 0 13 2
26 3 9 0 13 2 9 9 7 9 0 4 13 2 7 9 15 16 9 9 1 9 0 9 4 13 2
18 9 13 16 9 10 9 1 9 0 9 13 7 1 9 9 0 13 2
49 7 0 9 9 15 13 16 1 9 12 9 0 0 1 9 9 13 2 1 10 9 16 9 9 1 9 0 9 15 0 13 2 7 1 9 0 1 9 0 2 15 14 1 9 9 9 9 13 2
35 1 10 9 9 12 9 9 1 9 7 9 9 7 9 1 9 9 9 9 10 9 9 13 13 2 7 9 13 16 9 9 15 9 13 2
18 3 13 1 9 10 9 16 9 1 3 9 13 9 13 2 9 13 2
29 9 9 0 9 13 16 9 1 9 15 14 1 9 9 9 13 2 10 0 7 9 1 9 15 1 9 9 13 2
22 15 1 9 15 1 9 15 16 1 9 15 0 1 9 9 13 2 0 7 0 13 2
37 9 9 9 3 1 9 9 1 9 9 13 13 7 16 9 0 13 2 9 14 16 1 1 9 9 7 9 15 1 9 9 13 2 1 9 13 2
48 9 9 3 0 1 12 9 1 9 9 3 13 13 2 7 9 14 16 9 1 9 13 2 1 9 13 2 10 0 7 9 0 10 9 14 0 7 0 13 2 7 9 15 14 1 15 13 2
9 9 13 2 9 9 9 13 13 2
17 1 9 9 7 10 9 0 9 13 7 1 15 12 9 3 13 2
16 9 9 13 13 1 12 9 9 7 9 16 1 7 0 13 2
14 9 13 16 9 1 9 0 0 9 12 9 0 13 2
28 9 9 13 13 16 3 1 9 9 12 9 1 9 9 13 13 2 16 1 1 10 15 1 9 9 0 13 2
17 9 16 9 9 9 13 2 1 9 9 12 1 10 12 9 13 2
38 3 1 12 0 9 9 2 9 13 1 9 0 2 1 10 9 9 7 10 9 14 3 13 16 16 15 10 9 13 16 9 1 15 9 1 9 13 2
29 16 3 13 2 10 9 3 1 9 13 16 3 9 1 12 9 9 13 7 1 9 0 15 1 9 13 13 13 2
25 9 9 13 16 16 9 9 15 1 9 9 13 2 3 9 14 13 1 9 0 15 1 9 13 2
22 9 12 9 15 13 2 1 9 9 13 2 9 9 2 15 14 1 10 9 9 13 2
