1939 17
16 9 13 2 0 9 2 2 2 9 2 7 2 0 9 2 2
11 15 13 10 9 15 13 0 7 1 9 2
6 1 0 13 15 9 2
40 1 7 0 4 10 0 9 4 13 9 1 14 13 9 9 1 0 9 1 9 2 3 1 14 13 15 15 4 13 1 1 9 2 3 1 14 13 1 9 2
28 3 0 13 10 0 9 2 16 9 9 1 9 4 13 16 10 0 9 1 10 9 13 1 9 1 10 0 2
10 10 0 9 13 2 9 1 9 2 2
30 15 13 1 11 11 9 2 1 10 0 9 1 2 9 13 9 2 2 2 9 13 9 2 2 2 9 13 9 2 2
50 10 9 1 15 15 13 10 9 2 13 14 13 10 0 0 7 0 9 2 1 1 10 9 16 10 9 0 4 13 15 14 13 2 7 3 13 0 0 14 13 1 9 2 1 9 1 9 7 9 2
37 1 10 0 1 9 4 10 9 4 13 2 3 1 10 9 1 9 1 16 15 13 1 2 9 2 1 0 9 2 7 10 0 0 7 10 0 2
28 1 9 4 15 13 15 1 16 15 1 10 9 3 13 0 1 9 14 13 15 1 9 7 1 10 0 9 2
18 16 9 9 13 9 2 4 15 13 0 1 1 9 7 10 0 9 2
12 1 9 2 11 14 13 1 2 13 11 11 2
9 3 0 9 13 3 0 13 9 2
15 3 0 9 13 1 9 3 0 13 15 15 4 13 3 2
9 1 11 11 13 15 3 12 9 2
9 1 11 7 11 3 10 0 9 2
14 7 9 13 7 13 7 9 10 13 0 7 0 0 2
19 0 13 15 0 1 9 3 2 7 4 13 1 10 9 0 10 9 9 2
5 7 15 13 15 2
7 3 4 15 13 1 11 2
2 11 2
13 15 13 0 1 3 11 13 1 7 11 13 1 2
17 7 1 10 0 0 9 13 15 11 7 11 15 13 10 0 9 2
10 1 12 13 11 7 3 3 11 9 2
7 15 13 15 0 1 9 2
13 10 0 9 4 13 0 0 1 11 1 0 9 2
11 0 4 13 1 11 1 9 1 11 9 2
20 11 4 13 10 9 1 10 9 16 15 4 13 14 13 0 9 7 0 9 2
13 0 4 9 13 1 12 1 3 14 13 12 9 2
36 0 4 15 13 1 10 11 7 11 1 10 0 0 0 0 9 1 10 1 0 9 0 9 7 1 0 9 1 14 13 10 0 9 7 9 2
25 3 13 15 3 0 15 13 16 10 10 12 9 13 15 10 9 7 16 15 3 3 0 4 13 2
8 3 13 15 3 9 1 9 2
9 11 4 3 0 13 0 0 9 2
24 1 9 1 11 2 15 3 13 1 2 4 10 0 9 9 1 10 0 11 3 0 13 9 2
21 11 7 11 4 13 0 2 7 11 2 11 2 7 3 3 11 4 0 13 1 2
8 10 10 13 11 7 3 11 2
17 1 0 0 9 13 15 0 9 1 16 11 4 13 9 1 11 2
18 10 0 0 13 11 2 11 7 11 7 3 3 3 10 9 1 11 2
30 11 13 10 0 9 2 7 15 13 0 14 13 16 11 4 13 9 1 11 1 16 15 4 13 1 9 0 1 9 2
20 10 0 9 13 3 3 11 2 7 3 11 0 9 7 3 3 11 10 9 2
13 15 13 0 14 13 1 15 11 1 9 1 11 2
13 11 4 0 13 9 2 15 4 4 13 0 0 2
30 10 12 15 1 0 9 4 4 13 9 1 10 0 0 9 2 13 0 16 11 13 1 15 15 4 13 3 1 11 2
10 1 10 0 9 13 11 3 0 9 2
8 0 9 1 9 13 0 0 2
15 9 1 10 0 9 4 13 1 1 11 7 11 1 12 2
16 11 2 15 4 13 10 0 0 9 2 4 3 13 1 11 2
13 3 4 11 1 0 13 1 9 1 11 1 12 2
18 1 9 1 9 13 15 16 11 13 0 9 1 14 13 1 0 9 2
21 10 0 9 13 3 7 0 1 9 2 11 9 13 0 1 9 1 10 0 9 2
8 9 1 11 13 3 10 9 2
15 1 16 11 4 13 10 0 9 2 4 0 11 13 9 2
13 15 13 3 3 10 9 14 13 10 0 9 1 2
18 1 10 0 9 4 10 0 9 7 9 13 2 7 0 1 10 9 2
7 9 1 11 7 11 13 2
3 9 13 2
11 11 4 3 13 2 10 9 1 9 2 2
27 9 13 0 9 1 2 7 9 13 3 0 1 16 11 4 13 10 0 9 15 0 4 13 1 0 9 2
23 10 0 9 1 11 9 13 16 0 7 0 0 3 4 13 0 7 13 16 9 13 9 2
24 11 2 3 2 7 11 11 13 12 9 2 7 4 3 3 4 13 16 9 4 13 1 0 2
17 11 7 11 11 4 13 1 3 12 9 1 9 11 11 11 9 2
19 11 13 0 9 1 9 7 10 9 13 9 1 14 4 13 10 0 9 2
13 2 3 13 15 0 2 7 15 13 14 13 1 2
13 15 13 9 1 9 7 13 0 9 2 13 11 2
24 1 9 1 10 12 9 9 4 13 1 0 9 1 11 9 2 4 15 13 0 9 7 9 2
17 7 10 0 9 1 9 1 0 4 13 0 9 7 9 1 9 2
20 2 15 13 9 15 13 9 3 1 0 9 2 7 15 13 1 0 0 9 2
33 9 13 10 1 10 0 9 15 13 1 2 7 3 13 15 13 10 0 9 1 15 2 13 9 1 9 2 11 11 2 1 11 2
30 3 1 9 11 11 4 15 13 9 1 14 13 10 0 9 2 15 13 1 1 14 13 9 1 9 1 9 1 9 2
10 13 3 15 13 9 1 0 11 3 5
27 0 9 2 13 9 2 13 0 10 0 0 9 1 9 1 0 9 2 3 16 9 13 16 15 13 0 2
20 0 9 13 9 1 9 1 0 2 7 10 3 0 13 0 10 9 1 9 2
15 2 1 0 9 4 15 13 1 1 9 7 13 9 1 2
20 16 15 13 9 1 9 2 3 15 13 2 13 15 9 0 0 2 13 11 2
24 2 9 1 10 9 13 16 9 4 13 0 1 10 0 7 0 9 1 9 7 9 1 9 2
12 10 0 13 7 13 3 1 16 9 4 13 2
30 9 13 3 10 0 9 1 9 7 9 2 7 15 4 13 0 9 1 10 9 16 15 3 13 9 7 9 1 9 2
35 9 1 11 2 15 13 11 0 9 1 10 9 1 12 9 0 10 9 2 4 3 13 16 10 9 2 1 0 2 4 13 1 10 9 2
22 9 13 9 15 13 9 1 10 9 7 10 9 2 7 10 0 15 13 9 1 9 2
16 9 9 13 9 3 2 3 16 9 9 4 13 16 15 13 2
14 2 0 13 10 9 1 9 7 13 10 9 9 0 2
13 3 13 15 0 9 9 15 13 3 15 4 13 2
31 3 13 15 1 10 9 15 13 0 0 1 9 2 7 13 1 16 10 0 9 13 0 7 0 16 9 13 2 13 11 2
17 1 9 13 15 1 16 15 13 1 10 0 9 9 4 13 1 2
9 9 11 11 11 13 0 1 9 2
13 2 15 4 3 13 10 0 16 15 4 13 9 2
34 1 15 13 15 1 16 15 13 0 14 13 9 1 9 2 3 15 13 1 10 0 0 9 7 13 1 14 13 1 9 2 13 11 2
5 9 13 1 9 2
16 9 1 11 13 0 9 1 9 16 12 9 13 1 10 9 2
22 1 0 9 4 15 13 1 16 10 9 13 1 12 7 12 9 1 10 0 9 9 2
13 3 13 11 7 11 16 10 3 0 9 13 0 2
12 2 15 13 15 13 3 0 16 15 13 15 2
23 3 0 15 13 9 15 13 10 9 2 13 15 15 13 0 14 3 13 15 2 13 11 2
18 11 7 11 4 3 13 1 1 9 7 13 9 1 9 1 10 9 2
21 1 11 0 9 13 9 16 10 9 4 4 13 0 7 0 9 1 9 1 9 2
19 2 15 13 1 14 13 1 9 1 10 9 16 15 13 0 0 1 9 2
32 15 13 1 9 1 9 10 9 1 9 15 13 0 2 7 9 13 14 3 13 10 0 0 9 2 13 9 11 11 1 11 2
3 0 0 5
2 9 2
4 0 9 12 2
3 0 9 2
3 9 1 2
2 9 2
4 0 14 13 2
9 11 11 13 3 10 0 12 9 2
9 9 4 3 13 0 2 13 15 2
24 1 9 13 11 11 1 1 11 2 1 9 16 15 4 13 0 9 7 3 15 0 13 9 2
23 1 1 9 2 3 1 10 9 1 11 1 11 13 10 9 1 0 9 0 1 10 9 2
15 2 6 2 13 15 7 13 1 10 12 9 3 1 9 2
11 9 13 12 9 0 7 0 1 0 9 2
15 2 15 15 13 1 0 9 2 13 11 11 2 12 2 2
17 2 15 13 10 0 9 2 15 13 15 16 15 13 12 9 0 2
9 15 4 13 3 0 2 13 9 2
9 12 9 4 13 16 11 13 9 2
14 10 0 15 13 13 16 15 13 1 10 9 1 11 2
21 15 13 3 15 15 13 7 3 15 13 2 15 9 10 13 7 15 10 9 13 2
11 16 15 13 9 1 9 2 9 7 9 2
21 15 13 3 16 10 0 9 1 9 1 15 13 9 15 4 13 1 7 13 0 2
23 16 15 13 1 10 9 15 13 11 7 16 9 13 1 0 9 7 10 1 15 13 11 2
8 15 13 15 1 9 7 9 2
15 15 13 3 16 15 13 10 0 1 3 14 13 10 15 2
9 15 1 9 10 4 13 1 9 2
13 12 9 1 9 7 9 2 9 2 9 7 9 2
34 15 13 3 16 15 15 13 15 1 9 13 10 9 9 7 16 15 13 15 1 13 15 3 0 16 15 13 15 1 15 9 1 9 2
12 9 2 10 0 9 2 9 2 15 4 13 2
17 3 3 13 15 16 9 10 4 13 1 9 2 16 15 13 3 2
13 1 10 9 1 1 9 1 11 13 10 9 9 2
9 0 9 13 9 11 1 9 9 2
9 15 13 9 7 9 1 10 9 2
24 10 9 1 9 1 15 15 0 13 1 11 2 10 0 9 1 14 13 10 0 9 1 9 2
12 11 11 4 3 13 15 1 9 1 12 9 2
22 15 4 13 9 10 1 9 9 7 13 1 9 3 1 1 10 9 1 9 1 11 2
20 15 13 15 3 13 15 2 15 13 3 0 15 13 9 1 9 1 10 9 2
9 10 0 9 13 3 14 13 15 2
5 15 4 15 13 2
8 13 1 11 1 10 0 9 2
9 2 4 15 13 10 9 2 2 2
9 3 13 15 10 0 9 1 11 2
8 0 9 4 15 13 1 9 2
12 16 15 3 4 13 15 2 4 15 13 9 2
21 16 15 13 15 1 9 1 9 10 9 9 13 15 16 15 13 10 9 1 11 2
6 15 13 1 11 11 2
19 15 13 15 0 2 7 9 13 0 9 16 15 13 16 15 4 13 9 2
30 2 15 13 16 15 4 4 4 13 1 10 9 0 7 15 13 0 7 0 2 7 15 13 1 16 9 13 15 10 5
20 1 10 9 9 3 13 15 3 9 1 10 9 15 15 4 13 1 10 9 2
24 15 13 0 2 7 15 13 3 15 13 10 9 1 9 1 9 15 13 15 13 9 1 15 5
17 11 13 16 15 3 4 13 15 2 7 15 13 15 10 9 1 2
26 15 1 10 9 13 10 9 15 13 1 2 9 2 2 15 13 1 10 9 9 1 0 2 0 9 2
14 1 15 3 13 3 15 10 9 15 15 13 3 0 2
11 7 3 13 3 15 10 0 9 15 3 2
22 3 15 13 9 13 3 10 0 15 15 3 3 4 13 0 2 7 15 15 13 0 5
17 15 4 3 13 15 0 0 7 3 13 10 0 9 1 9 1 2
4 15 13 0 2
8 0 9 7 9 1 11 11 2
18 1 9 15 4 13 13 15 10 10 9 2 7 15 13 10 2 2 2
9 9 2 7 9 2 13 12 9 2
4 0 7 0 2
8 11 4 13 9 1 10 0 2
22 15 4 13 16 15 4 13 15 15 13 16 10 0 9 13 2 7 4 13 0 9 2
10 9 4 13 2 1 14 13 15 0 2
20 15 15 13 1 0 9 13 9 1 14 13 15 15 13 1 16 15 13 9 2
9 11 4 3 13 9 7 0 9 2
25 9 1 9 11 11 11 13 10 0 13 10 0 9 2 16 15 13 0 1 3 0 9 10 13 2
13 2 15 13 0 2 0 0 10 9 2 13 15 2
7 9 13 0 1 0 9 2
26 10 0 13 16 15 13 3 10 3 0 15 4 13 2 1 9 15 15 13 0 1 7 1 10 9 2
13 10 0 9 13 3 10 0 7 3 10 0 0 2
12 15 4 3 13 14 13 15 0 0 1 9 2
7 9 1 9 4 13 0 2
14 9 2 9 1 9 2 9 2 9 7 9 1 10 2
9 11 4 13 10 0 9 1 9 2
11 9 1 9 13 0 7 15 13 0 0 2
18 2 15 4 0 13 9 1 10 0 9 2 15 4 13 9 7 9 2
11 10 0 9 1 16 15 13 0 9 9 2
10 15 4 15 13 9 1 2 13 11 2
25 10 0 9 13 10 0 9 13 9 1 16 15 13 15 1 9 1 11 11 1 0 9 1 9 2
12 9 13 3 0 2 3 0 2 9 3 0 2
12 1 9 4 15 13 9 15 4 13 9 1 2
5 2 6 2 11 2
18 15 13 9 10 2 13 15 7 13 15 10 9 2 7 11 13 3 2
15 15 13 1 14 13 15 16 15 13 1 11 2 13 15 2
10 15 13 1 9 2 15 13 10 0 2
10 9 4 3 13 16 9 4 13 1 2
9 11 4 3 13 10 9 1 9 2
10 7 4 15 0 13 15 15 3 13 2
9 3 12 9 4 15 13 15 0 2
32 12 9 1 16 15 13 10 0 9 1 9 13 15 1 9 1 1 11 2 1 10 0 9 11 11 11 16 15 0 13 9 2
16 15 13 15 1 10 12 0 9 15 4 13 1 10 10 9 2
11 15 13 15 0 2 15 13 15 1 9 2
9 1 1 9 13 15 0 1 9 2
8 15 13 2 13 3 14 13 2
23 1 12 9 13 9 2 15 13 15 1 1 9 7 13 9 1 16 9 13 3 0 0 2
9 7 15 13 15 15 13 9 13 2
17 3 3 3 0 1 10 0 9 2 7 3 10 0 9 1 9 2
8 2 15 13 10 0 0 9 2
22 15 13 1 9 1 9 1 9 1 9 1 11 2 15 3 4 4 13 1 10 9 2
10 15 13 2 15 13 3 0 0 9 2
12 9 13 9 1 9 10 4 13 1 10 9 2
11 2 3 4 15 13 0 1 15 15 13 2
8 15 13 3 10 0 0 9 2
13 10 0 9 13 15 0 2 15 13 3 0 0 2
20 3 16 10 0 13 9 2 13 15 16 10 9 4 13 10 9 1 15 3 2
10 7 16 15 4 13 10 9 1 15 2
30 11 13 3 0 0 1 10 9 15 4 13 15 2 15 4 13 9 1 14 13 15 9 1 9 10 2 13 15 9 2
12 9 13 0 10 0 9 1 16 15 13 1 2
12 15 13 1 10 9 15 13 15 1 15 10 2
20 1 11 13 15 9 1 9 2 9 2 9 2 9 7 9 2 9 7 9 2
19 15 13 1 16 15 13 10 0 9 7 13 10 0 9 0 1 0 9 2
5 15 13 15 0 2
9 1 9 13 15 0 2 13 9 2
6 15 13 15 3 3 2
13 13 15 10 10 9 15 4 13 9 1 9 10 2
8 9 1 9 7 9 13 1 2
28 11 4 3 1 0 13 16 15 3 13 1 9 7 3 4 15 3 13 1 9 2 3 13 15 3 10 9 2
14 10 0 2 0 9 1 12 9 13 3 0 14 13 2
7 7 15 4 15 13 1 2
13 15 13 3 3 0 9 1 3 15 4 13 9 2
16 1 10 9 9 13 15 15 2 9 13 0 0 1 1 9 2
9 15 13 1 10 0 9 1 9 2
20 2 9 1 0 7 0 13 3 2 15 13 3 3 16 15 4 13 0 0 2
12 15 4 0 9 13 10 9 1 9 7 9 2
12 10 0 9 1 11 13 3 1 15 0 0 2
9 15 13 15 0 0 1 10 9 2
13 16 15 13 0 7 0 13 15 3 2 13 15 2
9 2 14 3 13 4 3 13 0 2
15 16 15 3 13 3 9 1 9 1 11 11 13 3 0 2
9 2 15 13 10 7 10 9 0 2
7 10 13 15 3 1 9 2
15 3 13 15 14 13 1 9 11 7 9 11 11 11 11 2
15 15 13 3 15 1 12 9 3 13 10 12 9 1 9 2
13 1 9 13 15 9 7 0 1 10 9 1 9 2
13 9 4 13 2 15 4 13 9 2 9 7 9 2
27 15 13 16 9 4 13 1 1 0 0 9 2 16 9 4 13 10 9 1 9 1 9 7 9 1 9 2
13 15 13 0 9 1 15 15 4 4 13 1 11 2
15 15 13 10 9 2 10 10 9 1 9 2 15 10 9 2
12 1 9 4 11 13 16 15 4 13 12 9 2
20 15 4 1 9 13 10 9 3 16 9 11 11 1 9 13 14 13 10 9 2
11 15 13 3 1 1 9 9 16 15 13 2
9 15 13 9 13 1 12 0 9 2
13 2 15 13 10 9 15 13 0 14 13 1 1 2
17 15 13 3 10 9 1 10 9 2 7 15 13 15 1 10 9 2
14 15 13 3 10 0 9 1 10 0 9 2 13 15 2
17 2 15 13 3 1 14 13 15 2 7 1 14 13 9 1 0 2
11 15 13 0 14 13 1 11 2 13 15 2
6 13 9 1 9 3 2
6 13 9 1 0 9 5
14 11 9 13 10 9 9 0 0 4 13 1 12 9 2
32 11 11 13 0 0 2 2 10 9 13 1 0 9 2 2 2 15 13 3 1 16 15 1 9 1 14 13 9 3 13 9 2
16 3 13 15 10 0 9 1 14 13 9 1 10 0 1 9 2
13 15 13 7 1 0 9 7 15 15 3 13 0 2
20 1 9 7 9 4 15 13 10 0 9 16 9 13 10 9 2 13 1 9 2
16 7 13 3 10 9 13 1 10 0 9 2 11 7 11 11 2
24 9 1 9 13 0 9 1 10 9 1 11 7 11 1 0 9 1 10 10 9 2 3 11 2
16 10 9 11 4 13 1 2 9 2 2 13 1 9 1 9 2
27 9 11 11 15 13 1 0 9 2 13 1 9 11 11 9 2 7 11 11 4 0 13 1 9 1 11 2
53 7 11 13 14 13 7 13 2 15 13 10 0 9 1 10 0 1 9 2 1 10 9 9 15 10 4 13 7 13 2 1 9 1 9 2 1 10 0 9 1 10 0 9 2 1 10 0 9 1 10 0 9 2
6 7 10 0 13 15 2
32 9 13 3 1 12 2 9 1 2 7 9 1 2 10 9 9 4 13 10 0 9 1 0 9 7 1 0 9 1 9 3 2
12 11 9 13 3 3 10 9 1 10 0 9 5
56 10 9 11 0 7 0 13 1 14 13 2 13 9 1 3 9 1 10 9 1 12 9 13 9 1 8 11 2 2 10 10 2 2 10 0 7 0 9 15 4 13 1 0 9 3 2 7 15 15 4 13 2 13 2 13 2
6 4 15 13 1 15 2
5 15 13 9 9 2
16 11 4 13 1 16 10 0 9 7 4 13 7 3 13 9 2
14 1 0 0 9 13 15 16 15 13 0 9 1 15 2
15 15 4 13 1 9 1 14 4 4 13 1 9 1 9 2
40 1 14 13 4 15 13 9 1 9 1 9 2 7 1 16 15 4 13 2 13 7 13 9 7 9 10 0 9 2 15 3 0 13 2 7 15 13 0 9 2
32 7 3 9 1 11 13 15 1 14 13 9 7 9 2 7 16 15 0 3 13 1 3 2 1 0 9 2 13 15 3 0 2
27 9 1 11 7 10 0 2 2 0 2 9 4 15 7 15 13 1 2 15 13 10 0 9 1 10 0 2
20 3 16 15 13 1 10 0 9 2 1 9 2 7 16 15 13 0 1 9 2
14 2 3 10 0 13 3 9 2 2 13 15 10 9 2
12 11 9 13 10 9 7 10 9 1 10 9 2
7 9 13 1 9 1 11 5
5 13 1 0 9 5
3 2 9 5
4 1 12 13 5
4 2 9 13 5
8 9 4 13 10 9 1 9 2
12 11 9 1 11 4 4 13 0 1 12 9 2
14 9 13 9 9 10 9 1 9 1 11 9 1 11 2
8 13 15 9 7 9 10 9 2
11 13 10 9 1 11 7 13 11 1 12 2
10 15 4 3 13 11 5 11 1 12 2
25 11 9 13 1 9 9 12 9 1 16 15 4 13 9 1 0 9 13 1 11 0 9 1 11 2
8 9 4 13 1 9 1 9 2
10 9 4 13 10 9 1 9 1 9 2
13 9 13 0 10 0 0 2 7 13 9 1 0 2
31 2 15 4 13 10 9 1 9 2 7 13 3 1 16 15 13 10 9 15 4 13 1 9 2 13 9 11 11 1 11 2
19 1 10 9 4 9 4 4 13 1 10 9 1 11 16 15 13 1 9 2
19 2 10 9 4 13 1 9 1 12 9 1 9 2 13 11 11 1 11 5
8 1 11 13 3 9 0 0 2
20 2 15 13 3 0 16 15 13 1 15 9 7 13 9 1 9 2 13 15 2
5 9 13 1 9 2
17 1 15 11 13 1 4 9 4 13 16 15 13 15 1 10 9 2
11 9 1 11 4 13 9 1 11 1 9 2
11 2 15 4 4 13 10 0 9 1 11 2
23 15 13 1 10 9 2 7 13 14 13 9 2 13 9 11 11 11 1 11 9 1 11 2
25 2 15 13 10 9 0 0 2 7 10 0 1 15 3 13 14 13 9 1 1 9 2 13 9 2
21 9 13 16 15 13 1 9 7 4 13 9 1 9 7 0 1 9 1 9 9 2
7 9 4 13 1 11 9 2
9 1 9 4 1 12 9 4 13 2
21 11 13 1 16 10 9 4 13 9 10 1 1 9 1 10 9 16 9 13 0 2
14 0 9 2 9 7 9 4 13 3 16 9 4 13 2
27 2 15 13 9 1 9 12 7 13 9 1 9 1 12 1 12 9 2 13 9 1 9 11 11 1 11 2
23 15 13 16 9 13 10 10 9 1 10 9 2 7 16 15 4 13 1 9 1 0 9 2
12 1 9 1 9 13 15 14 13 9 3 9 2
12 11 11 11 13 9 1 9 7 9 1 11 2
10 15 13 16 9 13 0 0 1 15 2
16 2 15 13 9 1 1 9 1 14 3 13 1 1 1 9 2
18 15 13 0 0 1 0 9 2 7 9 13 0 2 13 15 1 11 5
9 9 11 11 11 13 9 1 0 2
19 2 15 13 9 1 14 13 15 1 3 0 1 0 1 9 1 10 9 2
19 15 13 3 3 1 9 16 9 13 3 0 9 13 2 13 15 1 11 5
13 9 13 16 15 13 10 9 9 1 9 1 9 2
25 2 16 15 13 1 4 7 9 7 9 13 2 7 15 13 0 9 15 3 13 0 2 13 15 2
28 0 9 13 16 3 10 10 9 1 9 2 11 10 0 9 2 4 13 2 7 15 13 9 1 9 1 11 2
7 3 9 13 15 1 11 2
4 11 13 9 2
7 13 0 0 9 1 9 5
4 13 1 9 5
4 13 1 9 5
4 2 0 9 5
21 16 9 7 9 4 13 0 9 1 16 9 13 11 2 13 9 1 11 11 1 2
15 12 9 4 3 13 0 1 11 11 1 10 9 1 11 2
2 9 2
5 11 11 5 11 5
9 2 3 15 1 3 4 13 15 2
20 9 13 1 9 2 13 11 11 2 9 1 9 1 11 9 9 2 1 11 2
22 1 9 1 10 0 9 4 0 9 13 9 1 11 2 7 0 10 4 13 1 9 2
16 11 11 11 4 13 16 15 1 9 13 1 11 1 10 9 2
26 15 4 3 13 1 3 15 13 9 1 9 2 7 13 15 13 10 0 9 14 13 15 1 10 9 2
8 2 15 4 13 1 12 9 2
27 7 15 13 0 14 13 9 1 0 9 1 9 15 13 1 9 2 13 11 2 15 13 9 1 11 11 2
19 1 11 1 11 13 15 1 9 1 9 2 11 2 9 7 10 9 9 2
8 7 11 13 3 9 1 11 2
9 2 15 13 15 15 13 11 3 2
20 15 15 13 15 13 9 2 7 13 15 3 1 2 13 10 0 9 1 9 2
14 1 9 13 0 9 0 3 15 0 4 13 11 3 2
19 1 0 9 4 9 13 9 1 11 2 15 13 1 0 0 1 0 9 2
14 3 1 11 9 2 16 10 9 4 13 1 9 9 2
24 2 15 13 16 9 13 1 9 2 7 16 11 13 1 11 2 13 9 11 11 1 11 9 2
23 10 0 9 1 15 15 4 4 13 1 11 1 11 13 9 15 3 13 10 0 0 9 2
24 2 15 13 1 9 7 13 9 2 0 1 15 13 9 2 7 13 11 1 9 2 13 11 2
13 1 0 9 13 9 12 9 11 13 1 12 9 2
28 15 13 10 0 9 2 13 11 2 15 13 16 9 1 14 4 13 1 11 0 13 0 1 1 10 9 9 2
37 2 16 9 7 9 1 11 7 0 9 13 0 9 2 4 15 3 13 1 1 16 9 3 13 9 1 10 0 9 2 13 11 1 9 1 12 2
23 1 11 4 9 13 16 11 2 15 0 13 0 2 4 4 13 0 9 7 13 1 9 2
16 2 3 13 15 3 3 0 1 9 14 13 15 2 13 11 2
18 1 9 13 11 16 11 13 1 10 0 9 1 9 1 11 1 11 2
11 2 11 13 0 1 14 13 0 0 9 2
11 15 13 1 0 9 2 7 9 13 0 2
23 15 13 16 9 1 9 13 0 1 1 10 9 2 13 11 11 1 11 1 11 0 9 2
9 15 13 10 9 1 10 9 11 2
16 9 11 13 9 13 0 9 15 3 13 9 1 10 0 9 2
12 2 15 4 3 13 11 1 9 7 0 9 2
14 7 0 15 3 4 13 11 1 2 13 3 9 0 2
11 3 13 11 10 1 10 0 9 15 13 2
9 10 9 13 12 9 2 13 11 2
24 1 9 4 15 13 1 9 2 1 14 4 13 1 9 1 9 1 10 9 1 11 1 11 5
4 13 1 9 2
4 10 0 9 2
3 0 9 2
4 13 0 9 2
3 9 13 2
4 9 1 9 2
5 9 0 1 13 2
4 10 0 9 2
6 15 15 3 13 3 2
7 11 11 13 10 0 9 2
13 9 13 10 9 13 1 16 9 10 13 1 9 2
16 16 11 11 13 12 9 2 13 15 10 9 1 14 13 9 2
9 14 13 15 1 9 13 9 10 2
21 9 13 11 1 9 2 13 11 1 9 7 13 12 9 1 9 1 9 1 11 2
17 16 15 13 12 13 15 9 2 7 3 13 15 15 4 13 3 2
11 9 0 9 12 13 11 11 10 0 9 2
8 15 13 1 9 14 13 15 2
18 7 10 0 9 1 9 13 15 0 0 7 13 3 1 15 0 9 2
16 16 11 11 11 13 1 1 9 1 9 2 13 9 0 0 2
27 2 6 2 11 2 15 4 13 9 2 13 15 2 7 15 4 13 1 9 1 16 15 13 15 1 15 2
14 9 1 13 11 12 9 16 15 13 14 13 1 15 2
19 15 2 15 9 3 4 13 1 1 3 0 2 13 1 11 11 1 9 2
28 3 13 15 15 16 9 15 3 13 0 2 15 13 0 1 9 7 3 4 13 10 9 2 13 9 1 12 2
4 15 13 0 2
15 1 16 15 4 13 15 2 4 9 1 9 13 14 13 2
19 9 15 0 4 13 10 0 9 2 13 1 9 1 14 13 1 9 0 2
18 11 4 3 13 0 1 11 16 9 13 16 15 13 10 9 7 9 2
25 15 13 1 15 15 15 13 2 11 7 11 2 12 9 15 4 13 10 9 15 13 0 0 1 2
33 15 4 13 9 2 7 11 4 11 13 1 0 9 1 9 2 7 11 2 15 15 4 13 1 1 10 0 9 2 13 3 9 2
19 7 9 4 3 13 1 9 3 0 2 7 15 13 0 9 15 13 15 2
18 1 14 13 1 10 0 9 2 13 11 3 9 10 9 1 9 11 2
35 11 4 3 13 10 9 1 9 7 0 9 2 7 1 9 4 15 13 11 1 10 0 2 15 13 15 13 3 0 1 0 7 0 9 2
7 7 15 13 2 13 11 2
19 3 13 15 15 3 7 3 2 16 15 4 13 9 1 9 2 1 9 2
13 7 15 2 11 7 9 13 15 0 13 0 3 2
18 7 16 9 11 13 3 9 1 14 4 13 9 2 13 15 9 3 2
8 9 4 4 13 1 10 9 2
2 9 2
2 9 2
2 9 2
19 9 13 15 3 1 15 0 2 7 0 2 7 0 13 3 9 14 13 2
6 0 9 13 11 9 2
6 15 13 3 3 0 2
6 15 4 13 9 3 2
21 1 12 13 15 1 16 11 11 2 11 7 9 11 7 11 13 15 1 10 9 2
18 10 9 15 4 13 0 0 1 2 10 1 14 13 1 11 1 9 2
7 9 13 1 9 7 9 2
4 9 7 9 2
17 7 10 0 15 13 1 9 7 9 10 2 13 9 0 9 1 2
9 7 15 13 9 1 9 7 11 2
11 1 9 13 11 1 9 7 9 1 9 2
15 7 16 11 4 13 15 14 13 2 13 15 0 9 1 2
11 15 13 3 3 10 9 2 0 1 9 2
7 7 9 4 3 3 13 2
33 15 7 15 7 9 1 11 13 2 16 15 3 13 1 9 7 10 10 9 2 13 16 10 9 11 4 13 2 4 13 9 9 2
12 10 0 7 0 9 15 3 4 13 1 11 2
17 9 4 13 0 0 1 9 7 4 3 13 1 9 1 0 9 2
23 10 0 12 9 4 11 12 2 9 2 9 2 9 2 9 7 9 13 0 9 1 11 2
18 1 9 13 9 2 9 2 9 7 9 9 1 9 1 12 9 9 2
29 13 15 1 15 15 4 13 1 9 2 1 9 7 1 9 2 13 15 0 1 1 12 9 2 13 11 1 11 2
22 1 0 11 13 15 0 14 13 16 9 13 9 1 9 15 13 15 7 15 0 9 2
13 7 9 1 15 13 0 0 0 16 15 4 13 2
38 16 9 1 9 7 9 4 13 7 13 2 3 16 15 13 9 7 0 9 2 13 15 0 1 9 1 10 9 9 1 9 13 1 9 1 10 9 2
16 9 12 13 11 2 11 7 11 9 10 9 1 12 9 9 2
18 9 13 0 9 1 9 2 15 4 13 9 2 13 0 7 13 0 2
5 3 13 15 0 2
9 2 12 1 9 4 13 0 9 2
15 1 10 12 13 9 1 12 9 3 0 1 15 11 13 2
16 2 12 1 10 0 9 4 13 9 2 10 9 1 0 9 2
24 15 13 3 9 2 3 16 9 1 9 7 9 4 13 0 1 9 1 9 7 10 0 9 2
12 2 1 0 1 9 4 15 13 9 1 9 2
20 2 9 2 10 0 0 9 2 4 13 1 0 9 1 12 1 10 0 9 2
17 2 15 13 0 0 16 15 13 9 1 9 1 14 13 0 9 2
31 9 13 10 9 1 14 13 15 9 0 13 16 9 3 13 1 9 2 7 9 3 1 13 1 0 7 0 9 1 9 2
26 15 4 1 0 9 13 9 9 7 9 1 9 2 7 13 16 15 13 9 1 0 0 9 1 9 2
30 10 9 4 3 13 0 9 2 13 9 11 11 11 1 11 1 9 1 9 2 16 10 0 9 1 9 4 13 1 2
10 15 13 11 15 4 13 9 1 9 2
14 3 4 3 9 13 10 0 9 1 9 1 10 9 2
16 2 15 13 10 9 1 16 15 4 13 10 9 1 0 9 2
21 7 11 13 0 0 9 2 7 15 4 0 9 13 10 9 16 15 13 0 9 2
18 9 2 15 0 13 10 9 2 4 3 13 0 0 16 15 4 13 2
30 15 13 0 0 9 3 1 2 7 3 10 9 9 2 3 0 9 13 9 1 14 13 0 9 1 9 2 13 11 2
15 1 9 13 15 15 13 9 9 1 14 13 9 1 11 2
19 15 4 3 13 9 1 9 15 13 2 7 9 13 3 3 9 13 0 2
30 9 1 9 4 3 4 13 16 10 9 15 13 1 9 2 1 16 15 4 13 9 7 13 0 1 9 2 0 13 2
21 7 11 13 3 0 16 10 9 13 0 3 2 7 16 15 1 10 0 13 13 2
7 2 15 13 3 3 9 2
18 9 13 3 3 16 3 16 15 13 10 9 2 3 4 15 13 0 2
39 15 13 9 7 9 7 4 13 9 2 7 1 0 7 3 13 15 9 7 15 15 13 9 15 13 9 1 16 9 13 0 7 9 1 9 2 13 11 2
8 1 11 13 11 11 7 13 2
34 9 10 13 3 0 3 0 9 15 15 13 2 7 9 13 15 3 1 9 2 7 13 14 13 1 9 10 7 1 1 9 7 9 2
9 0 9 13 2 7 9 10 13 2
15 9 1 9 4 13 9 7 13 9 0 2 0 7 0 2
8 1 11 13 15 0 14 13 2
11 0 13 15 1 9 15 3 13 14 13 2
21 7 10 9 13 15 1 11 7 11 16 15 13 1 2 7 13 15 13 9 10 2
26 9 13 0 16 9 4 13 2 7 0 9 13 11 1 11 2 15 4 13 16 15 4 13 10 9 2
5 15 13 15 3 2
18 15 13 1 9 3 0 9 1 9 7 13 3 0 1 12 0 9 2
17 9 12 13 11 11 2 11 2 11 7 11 9 1 9 7 9 2
10 9 1 0 9 13 11 3 1 11 2
32 9 2 15 15 3 4 13 3 2 9 2 9 1 9 7 9 15 3 4 13 9 1 15 7 9 2 13 3 14 13 9 2
10 3 13 15 14 13 15 7 13 0 2
20 15 13 0 14 13 1 2 7 12 9 13 11 7 10 9 11 1 0 9 2
21 10 0 9 13 15 9 1 9 2 13 9 7 13 15 1 14 13 9 0 0 2
5 3 13 15 15 2
16 11 13 15 1 1 9 2 13 9 7 13 1 11 0 9 2
6 13 9 1 7 13 2
7 2 3 13 9 0 2 2
9 7 0 13 15 3 9 10 0 2
7 11 13 0 2 9 12 2
15 10 9 16 9 4 13 7 13 2 9 2 1 9 10 2
22 3 2 3 12 9 0 2 13 10 9 1 10 9 1 9 1 11 2 3 7 3 2
7 0 16 15 13 14 13 2
22 16 11 13 1 9 2 4 11 1 11 7 11 13 14 13 1 9 1 9 1 11 2
5 15 13 1 9 2
28 16 9 13 1 9 1 11 1 12 7 1 11 1 12 2 4 15 4 13 12 9 9 1 9 7 1 11 2
23 10 0 11 13 9 0 1 11 2 15 1 9 1 9 13 1 9 1 9 2 11 11 2
14 15 13 9 2 9 2 9 2 9 2 9 7 9 2
16 11 13 10 9 11 1 9 1 11 1 16 15 4 13 15 2
25 11 9 13 1 10 9 11 1 0 9 7 1 11 2 11 7 11 2 1 12 9 1 0 9 2
12 10 0 9 13 15 3 14 3 13 0 9 2
11 3 13 11 9 1 14 13 9 1 9 2
30 1 11 9 13 9 11 16 15 3 4 13 0 9 1 15 15 13 1 2 7 13 11 2 9 1 9 1 11 9 2
21 10 9 13 11 11 11 7 13 16 15 3 13 10 9 11 15 11 4 13 1 2
4 15 13 15 2
11 15 13 1 11 2 7 0 9 13 15 2
12 9 11 4 13 2 4 13 0 9 1 9 2
11 11 13 10 0 15 13 15 1 11 9 2
15 11 13 11 7 13 1 16 15 13 9 10 15 13 1 2
15 16 11 11 13 9 2 13 15 3 0 1 16 11 13 2
43 10 9 13 15 0 16 3 3 11 7 12 10 9 2 7 10 0 1 11 15 4 13 1 11 2 1 15 12 9 9 2 4 4 13 9 2 3 11 13 1 1 9 2
14 1 9 4 7 11 2 11 2 9 7 9 10 13 2
5 13 14 13 11 2
19 7 15 13 0 1 3 9 0 13 1 2 10 12 9 0 9 1 11 2
30 11 11 13 10 0 9 1 10 0 9 1 11 2 1 10 9 1 11 2 12 0 9 7 9 1 0 9 1 15 2
15 1 10 0 9 3 4 15 13 2 0 1 12 0 9 2
28 9 13 14 13 9 1 9 2 9 1 9 2 9 7 1 0 9 14 13 9 7 9 15 4 4 13 9 2
27 9 11 4 1 10 9 13 15 1 9 7 0 9 2 7 13 3 9 1 14 13 10 0 9 1 11 2
19 15 4 3 4 13 1 14 13 11 13 9 2 1 9 1 9 1 9 2
6 2 15 4 13 15 2
22 16 9 11 3 4 13 2 3 13 9 14 13 15 1 10 0 9 15 13 3 0 2
4 15 13 0 2
17 10 9 1 9 7 9 2 13 11 11 2 11 9 1 0 9 2
13 1 9 1 14 13 9 2 4 9 3 13 9 2
12 15 4 3 13 1 10 9 15 4 13 9 2
9 2 15 13 10 0 11 11 13 2
12 1 15 4 10 11 13 0 0 2 13 11 2
13 9 11 13 15 15 13 1 15 15 13 11 9 2
8 2 15 13 16 9 4 13 2
6 4 13 14 13 11 2
20 15 13 10 9 0 9 1 11 11 2 11 11 11 2 13 13 0 14 13 2
12 2 7 15 13 1 10 0 16 15 4 13 2
27 16 11 0 4 13 9 13 0 0 2 7 15 4 3 4 13 1 10 9 7 9 15 13 2 13 15 2
12 2 10 9 13 15 16 15 13 14 13 11 2
36 2 15 4 0 13 16 9 13 10 9 15 13 9 1 9 7 9 2 7 9 15 4 13 1 9 1 11 4 13 15 14 13 0 0 9 2
8 9 4 3 13 1 0 9 2
13 2 3 13 15 10 9 1 10 9 1 9 11 2
21 2 11 11 4 0 13 0 1 11 2 16 15 4 13 14 13 10 0 9 3 2
19 7 9 10 4 0 13 2 7 15 4 13 0 9 1 10 9 1 15 2
8 9 4 3 13 10 9 0 2
11 11 13 3 3 10 0 9 1 9 11 2
13 15 13 15 3 1 10 9 2 11 11 1 11 2
25 15 13 10 9 2 15 1 9 1 11 11 13 10 9 1 11 9 2 15 4 13 11 1 11 2
24 11 11 13 3 1 16 15 4 13 1 9 11 1 12 9 2 7 13 15 13 10 0 9 2
12 2 11 4 1 9 4 13 1 10 0 9 2
18 15 13 15 3 3 1 9 2 7 4 3 13 2 13 9 11 11 2
22 7 11 11 7 11 13 1 16 9 11 13 9 15 4 13 1 14 13 11 1 9 2
12 7 10 9 13 3 10 9 1 10 0 9 2
35 2 7 0 1 15 13 3 1 11 2 7 15 13 16 10 9 3 13 15 15 13 2 13 11 2 15 3 10 9 13 14 13 11 3 2
18 2 15 13 1 11 11 9 1 11 2 3 15 13 0 9 1 9 2
22 9 4 3 13 14 13 1 9 1 11 11 10 2 7 0 9 13 10 9 1 9 2
16 11 11 11 13 9 15 1 15 4 13 15 14 13 0 0 2
25 2 15 13 0 14 13 16 9 0 13 10 9 1 9 15 10 12 9 13 0 9 2 13 15 2
13 1 0 9 13 15 3 0 14 13 15 1 9 2
21 11 9 13 16 9 15 13 0 9 1 0 9 2 4 13 1 9 1 0 9 2
19 1 0 9 1 11 13 15 16 9 1 9 1 9 7 9 4 13 0 2
18 9 15 4 13 16 15 13 1 0 2 4 1 9 4 13 1 9 2
43 15 4 13 9 1 9 7 9 1 9 1 9 1 9 1 0 9 2 7 0 9 4 13 0 1 14 4 13 0 0 2 0 9 15 4 13 0 7 0 9 2 9 2
10 3 1 11 4 9 13 0 1 9 2
24 1 11 13 3 9 1 7 9 7 9 2 7 9 1 9 4 1 0 9 13 1 9 10 2
33 10 9 13 0 2 13 0 9 11 11 1 11 1 11 2 3 10 0 9 7 10 0 9 11 2 11 7 11 2 8 13 9 2
12 2 7 15 7 9 13 14 13 9 0 9 2
10 3 4 10 9 0 13 15 10 9 2
31 9 13 10 0 9 1 9 1 10 0 7 0 9 1 11 2 16 15 13 9 7 13 16 15 13 15 15 13 1 9 2
30 13 15 3 0 9 2 7 15 13 9 15 3 13 15 3 14 13 2 13 3 9 7 13 3 1 9 2 13 11 2
7 2 13 15 3 1 9 2
12 2 15 4 3 13 1 0 10 9 15 13 2
9 15 13 3 3 16 9 13 0 2
6 10 0 13 0 0 2
13 9 1 11 13 0 1 14 4 13 1 1 9 2
10 9 13 3 11 2 1 14 13 9 2
31 2 15 13 16 9 13 3 0 9 15 15 13 2 7 15 13 3 3 1 10 9 15 3 3 4 13 3 2 13 11 2
13 1 9 13 15 1 12 9 14 4 13 1 11 2
11 9 4 13 14 13 12 1 10 0 0 2
47 12 9 4 4 13 1 9 1 9 7 9 2 9 1 9 2 12 2 2 9 2 12 2 2 9 2 12 2 2 0 9 2 12 2 7 16 15 3 13 9 1 9 7 9 1 9 2
12 0 1 15 4 13 0 2 16 9 4 13 2
16 11 11 2 9 1 11 2 13 9 13 16 11 9 3 13 2
9 2 9 4 13 1 9 1 9 2
10 14 13 9 1 9 13 10 0 9 2
27 1 11 4 15 13 10 9 1 0 0 9 15 13 16 15 13 10 10 9 1 10 9 2 1 0 9 2
8 2 1 9 13 9 1 11 2
37 15 13 15 13 0 16 9 1 11 3 4 13 0 9 1 14 13 10 9 1 1 10 9 2 13 11 2 15 13 1 10 11 9 1 0 9 2
10 11 11 1 11 13 16 9 13 3 2
32 2 7 10 0 9 4 3 0 13 1 10 0 9 3 2 7 0 13 1 0 9 1 11 1 3 15 4 13 15 1 15 2
19 15 4 13 16 15 4 13 1 12 12 9 14 13 10 9 0 1 9 2
12 15 13 15 0 0 9 15 3 13 9 1 2
10 0 9 12 13 15 0 9 1 11 2
13 15 13 3 1 9 2 3 13 11 9 3 0 2
18 1 10 0 9 13 11 7 11 7 13 1 10 9 15 3 13 3 2
17 16 3 13 1 15 9 1 0 9 1 14 13 0 9 1 9 2
24 16 13 15 14 13 2 7 13 3 0 1 9 16 15 3 3 13 9 1 9 1 9 3 2
29 9 1 9 1 9 2 11 2 4 13 1 16 11 13 1 10 0 9 15 13 1 16 3 10 9 13 14 13 2
31 15 13 3 0 14 13 1 9 16 9 13 11 7 9 15 13 2 7 11 13 16 9 13 1 14 13 10 3 0 9 2
19 2 3 0 9 13 3 1 9 2 13 10 0 9 15 15 13 0 1 2
21 15 4 13 9 1 12 9 2 7 15 13 3 9 13 15 16 15 13 10 9 2
23 7 15 13 1 0 9 16 9 13 14 13 9 10 1 15 2 13 11 9 2 11 11 2
10 1 9 4 11 11 11 13 9 3 2
12 15 4 13 1 9 7 13 1 9 10 9 2
12 7 9 1 11 4 15 3 13 14 13 1 2
5 7 15 13 15 2
7 1 9 7 9 7 9 2
11 15 13 10 16 15 13 0 9 1 15 2
3 3 15 2
2 12 2
6 7 15 13 1 15 2
7 7 1 15 15 4 13 2
3 10 0 2
11 7 3 2 16 15 13 2 13 15 15 2
7 10 0 2 0 2 9 2
8 10 10 13 3 1 0 3 2
15 3 1 16 15 4 13 15 2 7 13 2 13 9 0 2
3 7 0 2
5 15 13 1 9 2
3 1 15 2
18 3 13 15 3 3 16 15 4 13 3 10 9 16 15 4 13 15 2
12 7 16 9 1 4 13 1 9 0 1 15 2
9 16 15 3 4 13 0 1 15 2
8 3 13 15 10 9 1 15 2
7 7 15 13 3 0 0 2
5 15 13 15 3 2
5 9 9 1 11 2
26 1 9 13 15 2 1 10 9 9 7 0 9 2 1 9 1 11 2 11 0 0 9 1 0 9 2
24 9 13 0 9 1 15 15 13 1 9 2 1 9 0 0 1 1 9 2 1 10 12 9 2
11 15 13 1 0 10 12 9 11 0 9 2
11 15 13 3 9 1 11 13 1 1 9 2
9 13 15 3 13 0 1 3 15 2
10 10 9 1 9 2 3 13 15 3 2
17 15 13 1 11 2 9 15 3 4 13 1 9 1 14 13 9 2
6 15 13 0 3 0 2
5 9 13 1 13 2
20 9 1 2 0 0 2 9 15 4 13 1 1 9 10 1 14 13 1 9 2
31 15 13 3 0 14 13 15 1 1 9 1 14 13 15 10 9 2 7 15 13 15 7 13 10 10 1 14 13 1 15 2
59 9 13 10 12 15 13 0 1 10 9 2 7 15 13 0 0 1 10 9 16 15 4 13 0 2 3 16 9 13 16 15 13 9 0 3 0 1 1 9 16 9 1 9 1 11 4 13 9 1 16 15 0 4 13 1 1 10 9 2
12 15 4 3 3 13 16 9 3 13 10 9 2
38 10 9 4 3 13 1 7 13 9 1 15 15 13 1 9 2 3 1 14 13 10 9 1 9 15 1 1 9 13 10 0 9 10 1 9 7 9 2
11 7 2 13 15 9 2 15 15 13 15 2
14 1 9 1 9 13 15 14 13 15 10 9 14 13 2
27 3 3 0 2 7 1 10 9 13 9 0 0 2 7 15 4 0 3 13 9 1 0 9 1 3 0 2
43 3 13 15 0 3 0 9 2 15 15 13 0 0 2 11 11 7 15 1 3 1 11 2 15 4 2 13 2 15 3 15 10 13 15 10 0 9 1 9 10 9 3 2
10 10 9 4 3 13 1 2 0 3 2
27 9 1 15 7 2 10 1 15 2 13 16 15 13 1 1 0 15 1 3 2 1 9 1 15 1 3 2
18 14 13 9 1 0 9 1 11 7 13 15 1 10 9 13 0 0 2
26 14 13 1 9 2 15 15 13 14 13 9 1 1 11 1 10 10 9 2 9 12 13 3 0 0 2
6 1 10 0 9 3 2
2 6 2
6 7 1 1 10 9 2
66 15 7 10 12 9 13 3 14 13 15 1 1 9 16 10 0 9 15 4 13 1 2 13 11 11 7 9 2 0 2 13 9 2 10 0 9 15 4 13 0 2 16 15 2 13 2 1 9 1 1 9 1 0 2 0 9 2 15 13 0 1 1 9 10 3 2
18 5 13 9 0 2 11 2 15 4 13 9 1 10 0 9 10 5 5
4 6 2 9 2
14 15 13 10 0 9 16 15 13 0 14 13 1 9 2
36 16 15 4 2 13 1 9 2 13 15 3 16 15 3 4 13 1 1 9 15 1 0 13 3 0 16 15 3 0 13 9 1 9 7 9 2
44 10 0 9 16 15 4 2 13 1 9 2 4 0 3 9 13 15 1 2 7 1 10 0 12 9 0 9 13 15 3 0 9 16 10 3 0 9 1 0 9 13 3 0 2
61 15 13 0 0 1 14 13 2 7 15 13 3 0 16 15 13 0 1 16 15 13 15 1 9 1 10 9 15 13 16 15 3 13 10 0 9 15 3 4 13 9 7 13 7 3 13 10 1 3 0 1 9 1 9 1 10 9 1 0 9 2
30 15 4 13 16 9 10 1 9 3 13 10 0 9 1 14 13 1 10 2 9 2 7 15 13 3 3 9 10 1 2
9 1 10 0 13 15 3 10 9 2
32 1 10 0 13 15 3 1 9 1 14 13 1 9 2 7 1 9 1 11 13 15 0 9 1 10 0 0 9 15 13 3 2
17 15 13 15 0 2 7 13 9 1 10 0 2 9 2 2 0 2
27 16 9 1 11 13 14 13 1 15 16 15 4 13 5 13 15 1 9 2 13 15 16 10 9 4 13 2
18 15 13 1 9 10 2 13 15 1 9 2 13 15 1 9 7 13 2
17 10 9 1 9 10 13 1 1 3 2 7 15 13 3 1 9 2
11 16 15 0 13 4 15 3 13 1 15 2
10 13 9 10 1 14 13 2 3 2 2
19 15 13 3 3 1 9 2 9 2 9 7 14 13 9 1 10 0 13 2
23 15 13 1 10 0 9 1 9 13 1 1 10 9 1 0 9 15 3 13 1 14 13 2
10 1 10 7 10 9 13 15 3 15 2
21 3 4 15 13 0 9 10 2 7 15 13 1 9 16 15 3 13 10 9 1 2
16 15 4 3 13 9 3 3 2 10 9 4 3 13 10 9 2
12 13 15 1 10 9 2 9 2 9 2 3 2
8 15 13 14 13 0 2 15 2
20 7 15 13 3 9 2 7 3 13 15 14 13 1 11 16 15 13 15 10 2
6 13 9 2 7 6 2
5 3 13 1 9 5
14 1 9 4 15 13 1 9 11 11 1 11 1 11 2
31 15 4 13 10 9 1 3 15 4 13 1 9 1 14 13 1 3 15 13 1 7 13 1 16 15 13 10 9 1 15 2
6 7 15 13 15 3 2
20 7 15 13 0 0 0 14 13 9 1 9 1 9 16 15 4 13 1 9 2
35 2 3 0 9 15 13 2 7 2 3 0 9 2 13 15 0 2 2 3 13 1 0 1 15 10 1 16 9 4 13 14 4 13 1 2
8 7 15 13 3 15 13 0 2
29 9 13 0 13 0 1 15 15 13 0 9 1 2 7 3 0 15 0 13 1 9 3 0 13 9 16 15 13 2
33 1 10 9 3 13 15 15 1 14 13 1 11 11 1 10 9 1 3 0 15 13 2 7 15 13 15 3 3 1 9 10 2 2
33 15 13 1 10 1 9 2 9 2 9 2 10 9 15 4 13 7 15 15 13 9 1 14 13 16 15 13 0 2 5 0 9 2
6 13 1 2 9 2 2
11 13 15 0 1 15 15 13 1 1 9 2
19 13 15 15 13 9 1 3 15 13 1 9 7 9 7 1 3 9 3 2
9 2 9 1 11 4 15 13 3 2
17 13 3 9 11 11 8 8 8 8 8 8 8 8 1 11 2 2
8 15 13 1 16 15 13 9 5
12 0 9 4 13 0 9 2 13 11 11 11 2
5 7 13 15 15 2
5 3 13 15 15 2
16 15 4 3 13 16 15 4 13 9 2 7 3 0 13 3 2
54 1 0 9 4 15 3 13 15 1 9 1 2 10 10 13 15 3 2 2 2 15 13 15 13 10 0 9 1 9 10 2 7 2 13 16 15 13 10 9 16 15 13 12 9 7 13 1 16 15 3 13 15 2 2
31 3 1 10 9 4 15 13 1 7 13 1 10 9 15 13 1 15 7 15 13 0 7 0 1 14 13 15 9 1 9 2
9 16 15 13 1 16 15 13 9 2
14 1 10 0 4 10 9 1 11 13 1 1 9 10 2
17 15 13 16 2 14 13 9 1 9 13 3 14 13 1 10 9 2
11 15 13 1 10 9 1 10 0 7 0 2
15 15 13 10 9 1 14 13 2 13 2 13 7 13 2 2
26 7 3 13 15 16 6 2 10 9 3 4 0 4 13 0 0 9 1 0 9 15 13 14 13 0 2
18 7 0 0 2 9 13 3 3 9 12 1 9 9 1 10 0 9 2
12 7 11 13 3 16 15 4 13 14 13 9 2
28 11 13 0 13 16 15 4 13 14 13 9 2 3 16 15 13 14 13 0 9 7 15 4 13 3 0 9 2
12 11 13 3 3 1 14 13 0 9 7 9 2
29 15 13 3 10 0 9 1 10 0 9 1 9 15 13 0 9 1 14 13 15 1 14 13 15 2 0 2 9 2
14 4 15 10 9 13 1 3 9 13 3 0 0 9 2
4 15 13 15 2
28 2 7 15 13 3 15 15 13 15 2 11 13 1 9 2 9 1 15 15 4 13 9 1 9 2 2 2 2
33 15 13 15 3 16 15 13 15 13 0 1 10 0 9 2 7 16 15 13 10 0 9 1 14 13 9 1 10 9 1 0 9 2
17 3 0 15 13 9 13 10 0 9 2 3 0 13 14 13 9 2
9 7 3 13 9 0 9 1 9 2
13 15 13 0 14 13 16 15 3 4 13 1 15 2
9 1 9 13 9 0 2 0 0 2
25 7 9 9 1 16 15 4 13 9 13 3 0 1 9 16 10 0 1 15 0 4 13 1 15 2
10 7 13 15 0 0 1 14 13 9 2
9 13 15 0 16 15 3 13 9 2
20 7 13 9 0 0 9 7 4 15 3 13 0 9 1 15 15 3 13 3 2
5 9 13 9 9 5
14 9 13 15 1 1 9 1 9 2 13 11 1 9 2
11 7 15 13 16 15 13 3 0 0 0 2
41 7 10 9 13 10 9 3 1 16 15 13 9 2 7 9 13 2 6 2 15 13 15 3 10 0 9 1 14 13 2 3 16 9 10 4 13 1 1 9 2 2
26 9 13 0 1 0 9 2 10 1 15 13 16 15 13 15 0 1 9 14 13 1 9 1 0 9 2
14 7 0 0 2 15 13 3 3 14 13 1 1 9 2
17 7 15 13 3 1 10 9 1 15 7 15 13 3 1 9 3 2
10 15 13 3 15 16 9 13 15 9 2
13 7 15 13 1 9 9 13 9 1 14 13 3 2
29 2 9 10 13 1 10 0 0 9 1 10 9 15 9 13 1 3 2 2 13 9 1 10 0 9 11 4 13 2
22 7 16 15 13 3 0 9 2 13 15 3 0 0 14 13 1 1 9 1 12 9 2
16 3 13 10 9 0 1 1 9 1 16 9 3 4 13 9 2
10 13 9 0 0 1 9 10 1 9 2
26 1 3 9 13 15 1 15 1 10 9 10 9 13 10 9 10 0 9 1 10 0 9 13 1 9 2
25 2 10 10 9 1 9 4 9 3 13 9 1 10 0 9 16 9 13 1 9 1 9 0 9 2
31 2 10 0 9 13 15 0 15 13 2 15 13 0 1 15 14 13 1 1 3 0 9 2 13 10 12 9 0 9 2 2
5 7 1 10 9 2
14 13 15 3 0 0 16 9 13 9 1 9 1 9 2
10 7 13 15 3 9 15 4 13 15 2
51 14 13 9 1 10 0 9 16 15 13 10 0 9 7 13 16 15 3 13 9 1 9 13 3 3 0 0 0 9 7 13 1 10 9 15 3 1 10 9 4 13 0 1 14 13 1 1 10 10 9 2
11 3 0 3 2 14 4 13 9 1 9 2
9 6 2 15 13 3 0 1 15 2
21 7 3 13 9 1 16 9 1 9 4 13 10 9 1 9 7 13 1 0 0 2
9 7 15 13 15 13 10 0 9 2
4 7 6 3 2
16 15 13 0 3 15 13 10 10 9 15 13 1 9 1 9 2
6 3 13 15 0 0 2
7 11 9 13 11 1 9 2
32 12 9 0 2 1 9 12 2 13 0 9 11 11 1 11 16 9 13 1 9 1 10 9 0 9 7 9 1 14 13 9 2
20 11 13 16 11 4 4 13 0 9 1 10 9 2 15 11 13 15 0 1 2
5 10 0 0 9 2
6 1 12 13 15 15 2
10 10 9 13 1 0 1 9 0 9 2
13 10 9 4 13 9 9 1 14 13 9 1 9 2
9 9 13 9 1 14 4 13 9 2
12 9 4 13 2 7 13 3 10 9 1 9 2
15 9 11 13 3 9 1 0 9 7 13 9 9 12 9 2
5 3 13 15 9 2
13 9 9 7 12 9 13 1 9 0 9 1 11 2
13 11 4 13 1 14 4 13 0 2 0 7 0 2
3 2 0 2
6 15 13 15 15 13 2
9 15 13 3 16 9 4 13 3 2
19 15 13 3 0 0 16 15 4 13 15 0 16 15 13 1 1 10 9 2
18 7 15 4 13 1 10 0 0 2 13 9 1 9 9 13 15 1 2
4 9 13 9 2
7 11 9 13 3 11 9 2
4 9 13 9 2
21 1 9 1 12 13 9 16 15 13 2 0 15 4 13 1 16 9 4 13 9 2
24 9 4 3 1 10 9 3 13 15 0 14 13 0 1 1 15 7 14 13 9 1 15 2 2
18 11 4 3 13 10 0 9 1 9 2 7 13 1 10 9 1 9 2
17 15 15 3 13 3 0 9 2 13 16 9 0 13 10 10 9 2
9 9 13 3 9 1 11 1 11 2
14 1 12 13 9 1 16 9 4 13 9 0 0 9 2
22 11 13 3 9 1 11 9 1 9 2 7 9 13 16 11 13 0 7 9 13 0 2
12 11 9 2 11 11 2 13 1 9 11 13 2
12 2 15 13 0 16 11 4 13 1 10 9 2
13 9 13 3 16 15 13 15 15 13 10 0 9 2
8 11 4 13 9 2 13 11 2
2 9 2
16 11 13 16 15 4 13 1 10 9 1 10 9 1 11 9 2
17 16 15 0 4 4 13 0 15 2 7 13 15 15 13 1 15 2
23 9 12 13 9 11 11 11 0 1 16 11 13 1 9 1 9 3 2 1 9 1 0 2
4 11 9 13 2
29 2 15 13 1 9 1 10 0 9 1 9 2 7 1 9 1 10 9 15 13 1 10 10 9 1 10 9 2 2
13 11 13 15 1 9 7 13 15 13 11 0 9 2
10 7 13 15 10 0 1 9 1 9 2
18 7 11 7 10 9 13 11 3 4 4 13 15 0 1 1 11 9 5
20 2 15 13 16 15 13 9 1 14 13 9 2 13 11 2 7 13 1 9 2
12 2 8 8 8 8 8 8 2 8 8 8 2
25 8 8 8 8 8 8 8 8 8 8 8 8 8 2 8 8 8 8 8 8 8 8 8 2 2
5 10 9 1 9 2
10 11 13 3 3 9 1 9 1 9 2
12 1 9 13 15 3 3 1 9 16 15 13 2
13 15 13 15 13 10 0 7 0 9 1 0 9 2
11 0 9 12 13 11 9 11 11 1 11 2
10 11 13 1 15 10 9 2 11 11 2
7 9 11 11 11 13 3 2
23 1 9 13 15 16 2 15 1 0 9 13 9 1 16 11 13 0 1 14 13 9 2 2
35 11 13 16 11 9 1 9 4 13 1 16 10 9 4 4 13 1 7 13 1 9 1 3 0 9 2 15 15 4 13 10 0 9 0 2
10 0 9 4 4 13 9 1 11 9 2
16 10 1 15 15 13 15 2 13 11 11 11 2 9 1 11 2
20 15 13 1 9 12 10 9 1 11 11 2 16 15 13 1 9 1 0 9 2
12 15 13 16 11 2 0 13 3 0 1 9 2
18 15 4 3 0 9 13 15 13 0 3 9 12 2 16 9 4 13 2
14 15 2 1 9 4 3 13 0 1 9 7 13 2 2
10 11 13 16 15 4 13 0 0 9 2
18 2 15 13 12 9 16 15 13 12 9 3 0 1 10 9 9 3 2
18 10 9 15 3 4 13 9 2 4 15 3 13 0 7 13 1 9 2
15 3 13 15 9 1 16 15 4 13 3 15 2 13 11 2
11 12 9 1 9 13 11 10 9 1 11 2
10 9 13 10 1 9 1 9 7 9 2
4 4 11 13 2
20 15 15 13 0 1 11 2 13 16 10 0 9 13 1 16 15 3 4 13 2
22 2 1 10 9 4 15 13 0 1 9 10 7 13 9 1 9 1 14 13 1 15 2
16 11 13 3 14 13 9 1 9 7 13 0 1 9 1 9 2
12 1 15 13 15 0 2 13 9 11 11 11 2
21 15 13 0 9 1 9 11 11 2 15 1 3 4 13 12 9 1 11 1 9 2
12 1 9 13 9 1 9 15 13 0 1 11 2
26 2 15 13 15 1 0 2 3 16 15 1 0 10 4 13 0 0 10 9 1 1 2 13 11 11 2
9 11 9 13 15 13 0 1 0 2
10 1 12 13 11 16 15 13 0 9 2
13 9 11 11 2 10 0 1 0 9 2 4 13 2
12 11 13 3 9 11 11 11 1 14 13 9 2
17 2 1 9 1 15 13 15 0 9 16 15 13 16 11 13 0 2
34 15 13 0 1 16 9 13 15 2 7 15 4 3 3 3 13 16 15 13 9 2 16 15 3 4 13 3 9 1 11 2 13 11 2
13 15 13 0 10 0 9 7 13 14 13 1 9 2
20 11 13 15 1 1 14 13 10 1 12 9 1 9 15 15 4 13 9 1 2
15 3 0 11 13 2 3 0 13 15 15 1 9 1 9 2
18 2 15 13 15 15 1 10 9 4 13 9 1 14 13 9 1 11 2
15 7 15 13 15 15 13 1 16 15 13 0 2 13 11 2
6 11 13 9 1 9 2
7 9 4 13 1 0 9 2
4 10 0 9 2
8 11 13 3 9 1 11 9 2
20 1 10 9 1 9 13 15 1 11 9 1 11 9 7 13 1 9 1 15 2
5 9 13 3 0 2
15 11 13 2 0 9 2 7 2 0 9 2 2 13 15 2
10 15 13 0 9 7 13 9 1 9 2
17 2 11 4 0 13 9 1 16 15 13 0 2 13 11 1 9 2
9 9 10 13 11 13 0 1 9 2
15 2 11 13 3 9 1 14 13 16 10 9 13 0 9 2
16 16 15 13 9 1 16 15 13 9 2 4 15 13 1 9 2
18 15 13 0 16 15 13 15 1 14 4 13 15 2 13 9 11 11 2
20 1 1 1 10 0 9 1 11 1 12 2 13 3 11 16 15 4 13 9 2
12 1 0 9 13 15 3 9 1 14 13 15 2
25 3 13 11 14 13 9 2 3 16 10 10 9 13 15 13 10 0 9 15 13 10 9 1 9 2
27 1 1 1 9 13 15 10 9 0 9 2 0 15 15 10 4 13 1 14 13 1 0 9 7 0 9 2
20 2 15 13 3 3 16 15 13 15 2 7 15 4 13 3 0 9 1 9 2
7 15 13 3 15 15 13 2
11 15 13 3 0 14 13 1 10 10 9 2
7 15 13 0 1 10 9 2
15 15 15 13 7 13 2 4 13 1 0 9 2 13 11 2
4 9 0 9 2
12 1 11 4 10 0 3 13 0 1 9 10 2
15 1 12 4 11 13 1 11 11 1 10 0 9 1 9 2
17 16 15 13 1 9 2 13 15 1 9 1 10 9 1 11 9 2
8 11 13 1 15 15 3 13 2
23 1 9 0 9 4 15 3 13 1 10 9 1 9 11 11 11 1 10 9 9 7 9 2
7 3 13 15 9 1 9 2
17 2 1 9 13 15 9 1 9 7 15 4 15 13 1 1 9 2
10 15 13 1 14 13 0 10 9 3 2
25 3 13 15 3 3 9 2 9 13 0 1 15 15 13 1 9 16 15 4 13 1 9 2 2 2
11 11 13 0 9 1 9 0 0 1 15 2
10 0 13 15 16 10 0 9 4 13 2
16 11 11 13 0 7 15 13 0 16 15 13 1 2 2 2 2
13 10 0 9 1 9 2 13 11 9 2 11 11 2
18 2 15 13 0 14 13 1 10 10 9 1 0 0 9 1 10 0 2
26 15 4 3 13 3 0 1 9 1 11 9 16 0 3 13 9 16 15 4 13 1 9 2 13 11 2
4 13 1 9 2
15 10 1 9 1 9 1 11 13 9 1 0 9 1 11 2
20 1 10 0 0 13 9 1 16 11 13 1 11 11 11 1 9 1 9 12 2
10 9 13 12 1 9 1 9 1 11 2
13 11 13 15 10 1 10 9 13 0 1 10 9 2
17 11 13 0 1 16 11 13 0 2 7 13 0 10 9 1 9 2
17 3 13 15 16 11 2 13 14 13 15 1 9 1 9 10 2 2
11 11 13 11 13 15 1 9 1 10 9 2
8 3 3 4 11 4 13 15 2
11 1 10 0 9 13 11 16 15 13 11 2
12 9 13 3 1 10 9 14 13 9 1 9 2
25 2 16 15 13 9 1 9 2 13 15 3 0 16 11 0 4 13 2 2 13 15 1 9 9 2
7 11 13 3 14 13 9 2
6 2 15 13 3 11 2
18 3 1 13 15 0 2 16 15 13 1 15 7 13 15 1 9 10 2
9 15 13 3 10 9 1 9 10 2
23 9 9 13 16 11 3 16 15 13 2 13 1 10 9 16 15 13 0 0 2 13 11 2
5 15 13 1 9 2
11 2 1 12 9 4 11 13 0 1 9 2
28 16 15 13 10 3 0 9 16 15 13 0 9 1 14 13 9 1 15 2 4 15 4 13 1 0 9 3 2
27 15 13 15 10 16 15 3 4 3 1 12 9 16 15 13 3 0 15 9 13 16 15 13 2 13 11 2
31 9 11 13 1 9 1 11 2 7 0 1 16 11 3 0 1 1 12 13 0 16 11 4 13 15 1 11 0 9 0 2
21 2 15 4 13 1 1 16 15 13 10 9 15 13 9 1 11 1 10 9 3 2
17 15 13 16 9 4 4 13 1 9 1 14 13 15 2 13 11 2
10 15 13 0 10 9 1 12 1 11 2
13 11 13 10 0 2 9 2 13 9 1 10 9 2
10 10 9 15 4 13 1 1 12 9 2
17 1 3 15 13 15 1 9 1 11 2 3 16 9 4 13 1 2
7 13 15 0 15 15 13 2
33 9 10 2 11 2 13 0 16 2 11 11 11 1 9 13 15 1 10 9 1 9 1 11 2 3 1 9 7 10 10 9 2 2
12 9 4 13 1 2 9 2 1 11 0 9 2
9 2 15 13 1 9 1 0 9 2
11 15 13 1 10 9 2 16 9 10 13 2
15 1 9 4 15 4 13 10 10 9 2 13 11 1 9 2
9 15 1 9 15 13 1 1 11 2
41 2 15 4 13 16 9 2 1 9 7 9 2 9 2 4 13 1 9 1 1 15 16 9 13 0 2 2 2 2 2 13 0 9 11 1 10 9 1 11 9 2
22 1 9 1 9 15 13 1 9 2 13 15 15 1 16 11 4 13 9 7 13 15 2
9 9 13 1 9 1 9 1 9 2
7 12 0 13 3 1 9 2
27 2 15 13 0 9 9 0 1 16 15 13 16 15 4 13 9 1 15 1 9 2 2 13 15 1 9 2
11 1 12 2 12 9 4 9 4 13 15 2
15 11 4 13 1 10 9 15 13 0 0 1 11 10 9 2
13 2 15 13 3 9 1 14 13 16 11 13 15 2
12 15 13 3 3 10 9 13 1 2 13 0 2
8 11 4 13 11 9 1 9 2
52 2 1 9 1 10 9 15 4 13 1 1 9 1 10 9 1 9 2 13 15 9 1 16 10 9 15 4 13 1 11 9 2 3 0 9 1 9 2 9 2 2 13 10 0 9 1 9 2 2 13 9 2
10 11 13 1 9 16 15 3 13 9 2
34 2 15 13 15 0 0 1 16 11 4 13 16 10 9 4 13 15 16 15 13 0 16 15 3 13 15 15 4 13 2 13 11 11 2
3 4 13 2
9 9 11 11 13 0 1 9 10 2
28 15 13 15 13 0 1 11 2 7 13 9 4 13 0 7 16 15 4 13 1 1 9 10 3 0 1 0 2
18 2 1 12 9 1 9 1 9 2 13 15 15 15 4 13 9 1 2
3 2 6 2
12 15 13 10 1 10 9 15 4 13 9 1 2
30 7 15 13 0 16 10 9 15 4 13 10 3 0 9 1 12 9 2 4 13 9 1 14 13 9 15 4 13 0 2
2 9 2
15 15 13 0 16 11 0 9 1 9 1 11 9 4 13 2
6 15 4 13 0 9 2
11 0 4 15 13 1 9 1 9 1 9 2
10 16 9 3 13 9 2 13 15 9 2
8 15 4 3 13 1 11 9 2
9 15 1 11 11 11 9 13 0 2
4 15 13 9 5
8 12 9 13 10 9 1 11 2
8 9 7 9 4 13 1 9 2
9 9 4 13 7 13 1 0 9 2
2 9 2
12 1 11 11 9 1 11 13 15 10 10 9 2
21 0 4 13 1 9 1 9 11 11 11 1 11 1 1 10 11 11 9 1 11 2
14 2 15 13 11 1 10 0 2 0 0 7 0 9 2
9 15 13 0 2 0 7 3 0 2
13 15 13 0 1 15 15 13 9 1 10 0 9 2
2 0 2
12 3 13 2 11 2 9 11 11 1 11 11 2
14 9 13 12 2 11 13 0 7 4 13 1 9 10 2
15 9 11 1 11 9 1 9 7 9 13 9 1 11 9 2
35 3 1 9 11 11 2 9 11 11 7 9 11 11 13 15 0 1 12 9 15 13 0 12 9 1 11 1 9 1 12 7 1 1 12 2
7 11 11 13 9 7 9 2
22 1 10 0 9 7 9 13 15 15 1 9 7 0 7 0 1 12 1 9 1 9 2
5 11 11 13 9 2
20 15 13 1 9 1 11 9 1 9 9 1 12 7 1 1 10 9 1 12 2
20 11 11 13 10 0 9 1 11 9 2 16 15 13 1 9 1 12 1 12 2
19 11 11 13 1 10 9 1 11 9 1 9 1 0 11 1 12 7 1 2
8 0 13 15 1 9 1 9 2
25 16 15 13 9 1 10 0 9 15 13 15 1 9 1 9 2 13 15 0 9 1 14 13 1 2
24 11 11 4 13 9 1 7 1 9 2 7 10 0 9 1 9 1 9 13 9 3 9 1 2
42 2 15 13 10 9 1 9 16 15 13 0 0 9 15 3 13 1 10 0 9 2 7 1 10 13 15 15 1 7 13 0 0 2 13 10 3 12 9 0 11 11 2
5 9 2 11 2 2
15 16 9 11 1 12 13 11 2 13 15 10 0 0 9 2
19 1 9 1 9 7 9 4 15 13 1 1 12 0 9 15 13 14 13 2
13 0 1 9 13 1 1 14 13 1 15 9 10 2
13 15 13 1 9 1 11 9 1 9 12 2 12 2
19 15 13 0 1 1 14 13 16 9 2 9 7 9 4 4 13 1 9 2
11 9 1 11 13 3 1 10 9 1 9 2
20 11 13 9 2 1 9 2 1 10 0 9 9 2 7 1 11 7 1 11 2
40 2 10 9 2 15 1 10 7 10 9 4 13 10 9 1 1 9 2 4 9 1 9 4 13 1 0 1 9 2 2 13 15 1 10 1 9 1 11 11 2
12 16 9 4 13 2 4 9 0 13 1 15 2
10 9 11 4 13 1 11 11 1 12 2
20 2 9 4 13 1 1 9 1 12 9 2 3 9 13 10 9 1 12 9 2
11 15 13 3 15 15 13 15 9 15 13 2
14 11 13 9 1 11 1 11 2 7 1 11 1 11 2
11 15 13 1 10 1 10 0 9 1 9 2
34 2 16 9 4 13 1 2 4 15 13 1 14 13 15 1 9 7 15 13 9 1 9 7 13 15 1 1 11 1 9 2 11 2 2
3 13 9 2
32 0 1 9 15 4 13 1 9 10 13 9 1 11 11 1 11 9 2 16 15 13 1 9 1 11 7 1 10 9 1 11 2
15 15 1 14 13 16 9 2 9 7 10 4 13 1 9 2
30 2 15 13 3 0 16 9 1 11 13 1 9 7 13 15 1 16 15 4 3 0 9 0 1 9 13 1 10 9 2
27 15 13 1 9 16 9 13 15 9 2 7 3 4 15 3 13 0 1 10 9 2 13 9 11 11 11 2
8 15 13 9 7 11 11 1 2
13 10 0 9 15 13 2 13 3 0 9 1 9 2
18 2 15 13 0 1 9 2 9 2 1 9 2 7 15 13 3 0 2
28 15 13 15 13 1 10 0 1 9 16 15 4 13 1 16 15 3 13 15 0 3 1 14 13 9 1 15 2
23 15 4 3 13 1 9 16 15 13 0 2 16 15 3 4 13 15 1 15 14 13 2 2
16 9 2 1 10 0 1 9 2 13 3 1 9 9 4 13 2
9 9 4 0 0 13 1 11 10 2
4 9 1 9 2
8 3 0 13 11 9 1 9 2
9 1 9 1 11 11 2 13 11 2
8 2 15 13 1 9 1 9 2
14 13 9 9 1 1 10 9 2 7 13 15 1 9 2
21 16 9 1 9 1 9 2 9 7 9 4 13 1 9 13 9 1 9 1 12 2
14 2 10 9 1 9 1 14 13 1 9 4 13 0 2
58 9 4 1 10 0 9 13 9 1 16 9 2 15 0 0 4 13 14 13 1 10 0 9 2 0 4 13 9 2 7 16 9 13 0 1 9 2 4 13 15 1 14 13 10 9 1 1 0 9 1 15 15 3 4 13 9 2 2
22 10 0 9 1 10 0 9 1 9 7 9 15 13 9 2 13 3 16 15 13 9 2
31 1 12 1 11 13 9 2 2 9 13 1 9 2 2 1 12 13 9 1 11 2 2 12 1 9 1 9 1 11 2 2
13 15 13 0 16 15 4 4 13 15 15 13 9 2
10 11 11 13 1 10 0 9 1 12 2
38 2 1 16 15 1 10 9 13 0 1 16 0 9 4 13 10 9 3 2 4 15 13 1 9 1 10 9 2 3 0 15 13 1 1 0 9 2 2
53 9 11 11 13 1 10 9 2 11 0 2 1 16 9 1 9 13 0 0 1 9 2 7 16 7 11 11 7 11 9 13 1 0 1 10 9 7 1 14 13 9 7 1 14 13 9 1 14 13 0 1 9 2
31 11 11 13 1 11 16 15 15 13 9 1 9 4 4 13 0 0 1 16 9 4 13 2 1 16 15 4 13 9 3 2
8 2 15 13 1 14 13 15 2
14 15 13 3 10 9 1 9 1 16 15 4 13 9 2
4 10 0 9 2
20 10 0 9 1 11 4 13 1 11 9 1 11 7 11 2 11 9 1 11 2
17 9 11 11 7 0 11 11 2 15 13 9 2 13 1 10 9 2
18 10 12 0 9 13 0 0 9 2 1 10 0 9 2 9 7 9 2
16 11 4 13 1 1 9 1 11 2 11 9 1 11 1 12 2
15 11 11 4 0 9 1 13 1 9 9 1 11 10 9 2
19 10 0 9 1 9 13 15 3 10 9 9 10 9 15 4 13 1 9 2
15 15 13 1 9 1 9 16 11 13 9 1 0 1 9 2
9 15 13 11 3 2 0 1 11 2
17 1 12 2 10 9 11 4 13 1 9 1 11 2 13 9 1 2
24 1 9 12 1 12 4 10 9 1 12 7 12 9 1 11 2 11 9 13 2 15 1 11 2
15 15 13 1 12 1 12 9 1 9 16 15 4 13 9 2
18 10 0 9 1 9 13 16 9 13 1 11 2 11 1 11 7 11 2
19 11 2 15 3 13 9 2 4 13 1 0 1 9 2 13 9 1 9 2
27 1 11 9 1 9 1 11 11 4 15 13 0 9 1 9 1 11 7 11 15 11 13 1 9 1 9 2
12 15 13 1 16 9 3 13 1 9 1 11 2
19 9 1 11 11 4 13 16 3 11 11 13 9 1 9 1 9 1 11 2
15 11 13 9 1 10 0 9 1 11 15 13 15 1 11 2
9 10 9 4 13 1 9 1 11 2
10 11 13 10 0 9 1 11 11 9 2
21 15 13 3 0 9 1 11 2 10 0 0 2 7 0 0 9 1 9 7 9 2
19 15 13 0 14 13 16 10 1 9 15 4 13 13 1 10 9 1 11 2
14 15 4 3 4 13 0 9 1 11 9 1 11 12 2
12 3 4 13 0 9 1 0 1 9 1 9 2
13 11 13 1 9 1 12 9 1 11 2 11 9 2
9 9 1 9 1 15 13 3 0 2
17 15 13 3 3 16 11 13 15 0 1 9 1 14 13 0 9 2
9 11 9 4 3 13 1 0 9 2
8 2 10 0 9 1 9 2 2
15 11 11 13 9 1 9 7 13 0 10 10 9 1 11 2
7 15 4 13 1 0 9 2
13 15 13 10 9 15 13 1 9 15 4 13 1 2
24 2 15 13 16 15 13 10 9 2 15 13 9 1 14 13 1 1 14 13 15 0 1 9 2
20 15 4 15 13 7 3 4 15 13 0 0 1 10 0 15 0 13 7 13 2
22 3 1 9 13 3 10 9 1 3 15 13 2 0 13 15 1 10 9 2 2 2 2
22 2 15 4 13 0 15 3 13 9 1 10 9 16 15 13 15 3 1 10 9 2 2
7 3 0 13 1 11 9 2
14 7 0 0 9 1 11 13 0 1 9 1 10 9 2
16 11 11 2 9 1 10 1 11 11 10 9 2 13 10 9 2
16 2 15 13 16 15 13 0 0 1 14 13 0 9 1 9 2
15 9 11 13 10 9 1 10 9 15 13 1 10 0 9 2
12 15 4 15 13 1 9 15 3 13 0 0 2
7 10 9 13 1 0 9 2
22 15 13 16 15 13 15 9 1 9 1 9 2 1 14 13 10 9 1 14 13 1 2
12 15 13 14 13 3 15 13 1 9 15 13 2
17 10 0 9 1 10 9 1 11 11 10 9 1 12 13 1 15 2
5 2 0 10 12 2
31 12 9 1 0 2 15 13 10 0 9 1 15 3 14 13 3 1 15 10 0 9 2 15 13 3 10 0 9 1 9 2
7 13 15 1 9 1 9 2
21 9 11 4 13 0 2 15 4 13 0 1 14 13 0 1 15 1 10 0 2 2
4 0 1 9 2
13 9 1 9 1 11 2 11 9 13 1 0 9 2
38 1 9 1 9 2 15 10 9 4 13 1 1 9 2 4 3 9 13 1 10 9 2 1 1 1 16 10 0 4 13 3 0 1 10 0 0 9 2
22 3 16 9 1 12 13 9 1 9 1 10 9 1 9 2 13 9 1 10 0 9 2
19 11 11 13 1 12 2 7 1 12 13 11 1 15 9 1 14 13 9 2
23 11 2 11 9 4 3 13 1 9 1 9 1 0 1 9 2 7 10 9 13 1 9 2
19 1 12 13 10 0 9 11 11 1 0 9 1 9 1 11 2 11 9 2
13 2 15 13 1 9 1 11 14 13 1 1 9 2
13 4 3 15 13 2 4 9 4 13 2 13 11 2
10 9 13 10 9 1 9 0 1 9 2
16 9 13 0 14 13 7 9 1 9 15 4 13 1 9 13 2
13 11 7 9 11 11 13 9 15 4 13 9 9 2
20 3 4 9 13 9 1 10 9 1 9 2 3 4 9 13 10 0 0 9 2
4 3 13 9 2
17 3 1 12 13 10 0 9 2 7 3 4 11 13 15 1 9 2
3 13 1 2
8 9 1 9 13 1 10 9 2
13 0 0 9 13 16 0 9 13 14 13 10 9 2
14 3 13 15 9 2 7 1 1 9 13 10 0 9 2
10 1 9 13 11 11 10 9 1 9 2
9 15 13 9 1 10 9 11 13 2
19 1 10 0 0 9 1 9 13 15 7 9 7 9 2 7 15 13 9 2
21 15 13 0 16 15 13 7 13 9 1 11 2 11 9 2 13 0 0 1 9 2
15 1 9 13 15 9 1 9 2 7 13 10 9 9 13 2
21 1 9 1 9 7 9 1 9 13 11 9 1 9 1 0 9 7 10 0 9 2
11 15 13 7 1 9 1 9 7 1 9 2
10 9 4 1 10 9 13 1 0 9 2
15 0 9 2 0 9 7 0 9 13 1 9 1 11 9 2
22 11 9 4 1 10 9 1 12 13 11 9 1 9 1 9 1 9 15 13 1 9 2
55 2 16 15 13 10 0 9 15 4 13 1 10 0 9 1 9 2 13 1 9 9 3 10 9 1 16 10 9 1 9 1 9 1 9 13 0 1 1 15 15 10 9 13 10 0 9 7 0 7 1 9 1 0 2 2
20 11 11 13 1 11 16 15 3 13 9 1 10 9 7 3 3 4 13 15 2
12 11 11 13 1 9 1 11 1 0 12 9 2
22 15 13 1 9 14 13 1 10 0 9 1 9 1 11 1 16 9 4 13 1 12 2
12 15 13 1 1 9 1 12 2 12 9 0 2
4 9 1 9 2
7 12 9 1 13 11 11 2
9 15 13 9 1 10 1 10 9 2
12 1 9 1 15 1 11 9 13 9 11 11 2
22 2 0 9 15 13 15 2 13 15 15 9 1 10 10 9 15 4 13 1 14 13 2
6 15 13 10 0 9 2
22 15 13 3 15 4 13 1 10 0 7 4 0 0 13 1 0 10 9 1 9 2 2
26 9 2 15 9 1 11 11 4 13 9 1 2 4 13 1 9 9 1 1 9 13 13 1 0 9 2
13 15 13 1 10 0 9 2 7 1 12 0 9 2
16 3 13 10 9 2 3 9 1 10 9 1 11 11 0 9 2
13 15 13 0 1 10 9 15 15 4 13 12 9 2
10 7 15 4 3 13 15 1 12 9 2
9 2 7 13 3 10 9 12 12 2
18 2 6 2 15 13 15 10 9 2 7 9 1 9 13 10 0 10 2
7 3 4 15 13 10 0 2
20 15 13 3 3 2 7 15 13 15 15 10 9 2 15 15 13 0 9 1 2
22 2 16 15 1 9 4 4 13 2 4 15 13 16 15 13 9 1 9 7 3 9 2
3 2 6 2
12 2 15 13 15 15 14 13 1 10 10 9 2
9 2 15 13 1 1 14 13 9 2
7 15 13 10 9 1 15 2
6 2 15 13 10 9 2
3 2 6 2
8 7 15 13 0 0 14 13 2
8 6 2 15 4 13 15 9 2
6 15 13 3 3 3 2
9 9 13 10 9 2 9 10 10 2
20 15 13 9 15 13 9 2 9 15 13 7 9 1 0 0 9 16 15 13 2
5 7 9 7 9 2
18 7 3 13 3 15 3 0 1 10 9 2 13 11 7 13 9 1 2
6 15 13 0 1 9 2
3 10 0 2
16 11 9 1 9 1 10 0 9 4 0 13 1 10 10 9 2
11 9 1 11 13 1 15 1 9 1 9 2
9 2 15 13 15 1 15 1 9 2
13 2 15 13 3 3 16 15 13 1 9 1 9 2
9 3 2 15 4 3 13 15 3 2
49 1 9 13 15 1 9 1 10 9 1 11 2 7 1 9 13 15 9 1 16 15 13 1 14 13 0 7 0 7 15 4 13 12 9 2 15 4 13 9 7 13 1 12 9 9 10 1 9 2
18 3 13 15 10 9 7 13 16 15 3 13 0 0 14 13 1 11 2
4 8 8 8 2
6 0 9 13 10 9 2
5 15 13 0 3 2
18 2 3 13 15 14 13 0 16 9 1 9 1 11 13 15 3 0 2
6 2 15 13 3 0 2
6 15 13 3 12 15 2
18 15 13 10 9 15 13 10 9 1 9 15 15 4 13 15 3 13 2
24 16 15 4 13 1 3 0 15 13 2 13 15 16 15 13 1 10 9 2 7 3 13 15 2
8 2 8 8 8 2 8 2 2
15 2 3 0 4 15 13 1 14 13 1 1 9 1 9 2
9 2 15 4 15 3 13 0 1 2
8 3 4 15 13 1 1 15 2
18 16 15 4 13 10 9 2 4 15 3 3 13 0 7 0 1 9 2
7 3 13 15 10 0 11 2
6 15 13 14 13 12 2
14 3 13 15 15 12 1 9 2 7 15 13 1 9 2
8 15 13 1 10 9 12 3 2
20 2 15 4 3 13 16 10 0 9 1 9 4 13 15 2 1 9 7 9 2
15 3 4 15 3 13 1 9 10 15 13 16 15 13 12 2
14 7 1 9 4 15 13 9 7 1 9 7 1 9 2
7 15 13 0 0 14 13 2
11 3 4 15 13 0 14 13 10 12 9 2
4 12 7 12 2
19 2 9 1 9 2 16 15 13 1 15 2 13 3 0 1 9 1 9 2
18 7 15 13 0 1 14 13 16 15 13 0 1 9 15 13 3 1 2
23 15 13 3 1 9 16 15 13 12 9 0 1 15 2 7 15 13 3 1 15 10 9 2
7 7 3 2 10 0 9 2
6 10 9 13 0 9 2
21 7 15 13 10 9 1 2 7 3 4 3 10 9 1 11 11 13 3 0 9 2
15 15 13 0 1 9 7 11 11 4 4 13 3 1 11 2
11 2 15 4 13 10 9 13 0 7 0 2
15 9 2 1 11 2 13 0 0 9 1 11 2 11 11 2
12 15 4 0 13 3 1 11 11 1 0 9 2
7 3 13 15 1 11 9 2
11 2 15 13 10 9 15 13 0 0 1 2
19 9 11 11 4 13 9 11 11 4 13 1 15 7 13 15 10 9 9 2
9 2 13 15 15 3 11 12 9 2
8 2 6 2 6 2 10 15 2
9 7 15 13 2 0 9 7 9 2
11 15 13 3 10 9 10 9 9 1 9 2
11 7 11 13 3 15 13 15 3 0 9 2
8 1 9 13 15 1 11 11 2
2 11 2
2 11 2
5 7 9 1 11 2
11 2 3 13 15 7 13 15 15 4 13 2
6 7 15 13 15 13 2
3 11 13 2
7 7 3 13 15 1 15 2
13 15 13 3 3 0 9 2 15 13 0 10 9 2
7 11 13 1 10 0 9 2
11 2 15 13 0 10 12 9 15 4 13 2
6 7 15 13 0 0 2
22 7 2 15 15 13 2 15 13 3 3 3 16 15 3 13 10 0 2 3 13 9 2
22 2 15 13 3 9 15 13 0 0 1 15 2 15 13 0 9 1 15 15 13 1 2
5 3 13 3 15 2
9 15 13 0 7 0 3 0 0 2
5 15 13 1 9 2
8 0 13 15 9 1 9 3 2
8 15 13 3 9 15 3 13 2
10 15 13 1 9 1 1 9 1 11 2
9 9 7 9 11 11 4 13 15 2
9 15 13 10 0 9 1 1 9 2
12 2 3 13 15 0 16 15 13 9 1 9 2
6 15 13 3 3 15 2
2 6 2
20 7 15 13 3 12 9 1 0 9 2 10 9 1 9 2 9 1 1 9 2
11 15 13 1 9 2 13 1 10 0 9 2
6 13 0 1 7 1 2
3 2 6 2
7 3 13 15 0 3 3 2
5 3 13 15 9 2
22 2 15 4 3 3 3 13 1 9 1 11 2 3 13 0 1 15 15 13 1 9 2
19 15 13 10 9 1 16 15 3 4 13 1 15 15 4 0 13 1 0 2
8 11 13 10 0 9 1 9 2
15 2 16 15 13 1 9 2 13 3 3 16 15 13 0 2
6 15 4 13 0 10 2
5 15 13 0 10 2
5 15 13 10 9 2
26 7 15 13 9 2 15 13 0 2 15 13 3 1 0 9 2 15 13 15 0 2 13 1 0 9 2
3 10 15 2
25 15 4 3 13 1 9 1 10 0 9 7 13 16 3 13 15 15 4 13 1 15 9 7 9 2
8 15 4 3 4 13 15 3 2
3 13 15 2
5 2 9 1 11 2
4 3 1 9 2
9 11 11 13 10 1 11 0 9 2
3 0 9 2
12 1 9 13 3 0 9 7 9 1 1 9 2
3 9 1 2
7 11 7 11 13 3 0 2
11 1 14 13 1 9 13 9 1 1 9 2
2 13 2
10 9 13 3 0 0 1 9 7 11 2
16 9 4 13 1 9 2 1 9 13 11 2 11 2 0 9 2
2 0 2
7 9 13 1 10 0 9 2
2 9 2
13 16 15 4 13 3 9 2 4 15 13 10 9 2
9 9 1 9 13 9 1 1 9 2
4 9 1 9 2
6 11 13 9 7 9 2
5 9 13 1 11 2
2 9 2
6 11 13 0 1 9 2
8 10 0 9 13 0 1 9 2
16 9 4 13 1 10 0 9 2 15 3 4 13 9 7 9 2
2 9 2
11 9 1 9 1 9 13 1 10 0 9 2
9 9 9 1 9 13 0 1 9 2
8 9 1 9 13 1 11 11 2
2 13 2
13 0 3 2 0 1 9 7 9 9 2 13 11 2
2 9 2
10 9 4 13 1 9 1 11 7 11 2
7 3 1 9 13 15 9 2
14 10 0 9 13 1 9 1 1 11 11 2 12 2 2
6 2 15 13 14 13 2
8 9 13 10 10 2 13 15 2
5 1 9 13 0 2
15 10 9 9 13 1 9 2 7 1 9 13 10 0 9 2
23 1 9 13 9 11 11 11 2 12 2 7 9 11 11 2 12 2 1 9 0 1 9 2
13 2 9 13 0 16 15 3 4 13 2 13 11 2
11 1 0 12 9 4 15 13 3 1 9 2
19 1 9 13 15 9 1 11 11 7 11 2 1 11 9 1 11 7 9 2
12 9 7 9 13 0 7 10 9 4 13 9 2
19 13 15 9 7 0 2 13 15 1 9 10 0 9 7 3 10 0 9 2
7 9 4 0 13 1 9 2
14 9 1 9 13 0 1 10 9 1 10 9 1 9 2
16 4 15 13 9 1 0 14 13 1 2 13 15 12 9 1 2
12 2 15 13 15 3 0 16 15 13 12 9 2
12 15 13 3 1 9 2 7 13 3 10 9 2
8 15 13 10 9 1 11 3 2
15 3 0 2 7 15 4 13 1 9 2 13 15 7 13 2
17 10 0 9 4 15 13 0 9 1 10 9 15 13 1 0 9 2
14 1 10 9 13 9 15 3 13 9 1 11 8 11 2
13 9 1 9 13 1 9 2 9 1 10 0 9 2
12 2 15 13 9 7 0 9 2 1 9 11 2
9 7 15 13 3 3 9 15 13 2
11 1 0 1 9 4 15 13 0 1 9 2
16 15 13 1 10 9 7 13 16 9 4 13 0 2 13 15 2
9 9 1 11 13 0 1 12 9 2
8 15 4 13 7 9 7 9 2
22 15 13 0 7 13 3 12 9 1 9 2 3 1 9 2 7 1 9 1 10 9 2
16 3 13 15 1 9 2 13 9 2 13 10 0 9 7 13 2
14 1 3 13 15 1 2 1 9 2 9 2 7 9 2
24 13 0 0 1 14 13 9 1 10 0 2 11 11 2 1 11 7 1 9 11 11 1 11 2
15 10 9 13 15 1 11 7 13 15 9 1 9 1 11 2
21 3 13 15 9 16 15 13 1 9 2 0 1 9 2 0 9 7 9 1 9 2
17 0 13 15 1 10 9 2 3 0 13 15 10 0 9 11 11 2
15 2 11 0 9 2 2 13 9 1 2 11 2 1 11 2
19 11 4 13 1 9 0 9 7 13 9 1 1 10 11 11 9 1 11 2
13 16 15 13 11 2 13 15 0 0 9 1 9 2
14 2 10 9 13 15 11 10 9 1 10 0 0 9 2
9 10 9 13 15 7 13 10 9 2
9 15 13 15 10 9 2 13 11 2
5 9 13 1 15 2
5 15 13 3 9 2
15 3 13 9 7 9 1 9 16 9 13 1 9 1 9 2
25 3 4 15 13 1 14 13 11 0 9 7 1 10 0 9 1 9 2 15 13 1 9 1 9 2
16 2 15 13 0 3 14 13 9 1 14 13 0 2 1 9 2
13 15 13 1 14 13 9 1 9 2 13 0 3 2
20 16 10 9 13 2 13 15 10 10 2 13 11 16 15 0 13 10 12 9 2
6 2 13 9 0 0 2
14 3 13 15 9 1 0 9 7 13 14 13 3 0 2
14 11 4 13 1 1 9 1 9 7 4 3 13 9 2
16 14 13 1 9 7 13 9 13 3 3 0 1 14 13 1 2
8 9 11 2 3 2 13 9 2
6 9 13 3 3 0 2
7 3 3 13 15 0 0 2
11 15 13 1 1 9 7 13 2 11 2 2
12 11 13 1 2 8 8 11 2 9 1 9 2
8 1 9 13 15 2 9 2 2
10 2 1 9 13 15 3 0 7 0 2
12 15 13 3 3 9 13 15 1 2 13 11 2
17 15 13 9 1 9 16 15 4 13 1 10 9 2 9 7 9 2
5 15 13 9 3 2
23 15 13 1 9 7 9 1 2 0 2 0 9 2 2 1 9 2 9 2 9 7 9 2
12 15 13 9 2 9 7 9 7 13 3 9 2
5 2 9 1 11 2
4 3 1 9 2
18 16 3 11 13 1 15 3 11 1 10 0 9 2 13 15 10 9 2
6 11 7 9 13 3 2
4 13 9 1 2
16 15 4 3 13 15 1 2 9 2 2 9 7 9 0 9 2
15 2 9 13 1 9 1 9 2 7 15 4 13 0 1 2
12 15 15 13 1 2 13 15 15 13 9 1 2
14 0 1 2 9 2 4 13 0 9 7 4 13 0 2
5 15 13 15 9 2
17 15 13 3 3 2 0 2 2 3 16 15 13 10 9 1 9 2
7 2 9 13 3 3 0 2
13 15 13 0 1 15 2 0 9 2 9 7 9 2
9 15 13 0 9 1 0 9 3 2
5 3 13 15 9 2
25 1 9 11 9 1 9 1 9 1 9 7 9 0 2 1 10 9 1 1 10 0 2 0 9 2
6 9 13 10 12 9 2
7 2 0 13 2 13 11 2
23 2 15 13 15 13 1 0 9 2 1 9 1 9 2 1 9 1 9 1 10 0 9 2
11 10 0 9 13 15 1 12 9 1 9 2
16 13 1 16 2 9 13 2 2 13 1 9 1 9 7 9 2
6 15 4 13 10 9 2
6 2 3 15 13 9 2
7 16 9 13 10 0 9 2
4 9 13 0 2
14 13 15 9 2 13 15 16 15 13 0 14 13 9 2
6 3 13 9 0 0 2
7 9 7 9 13 0 9 2
15 9 13 0 2 7 15 13 10 0 9 2 13 11 11 2
9 15 4 3 3 13 1 12 9 2
7 3 0 4 11 11 13 2
21 9 4 13 3 0 2 7 13 3 1 1 10 9 1 0 9 7 9 1 9 2
12 2 3 4 15 13 3 0 3 2 13 15 2
10 2 10 0 1 13 14 13 0 9 2
18 13 9 1 1 9 2 3 9 7 9 1 9 1 9 9 7 9 2
10 15 13 15 13 1 0 9 1 9 2
6 9 13 1 1 9 2
8 0 1 10 0 9 1 9 2
13 2 15 13 0 2 11 11 7 11 11 2 11 2
6 9 13 0 1 11 2
7 2 11 11 2 13 11 2
9 2 3 13 15 0 2 13 11 2
11 2 15 13 14 13 15 7 13 11 11 2
7 2 9 13 1 10 9 5
5 11 1 9 1 2
5 11 11 1 0 2
23 11 11 11 7 11 11 11 13 1 12 0 1 9 1 12 9 9 9 1 11 1 9 2
10 0 11 11 13 1 9 1 9 12 2
8 11 13 1 12 9 1 9 2
9 11 11 11 13 9 12 1 11 2
10 7 11 7 11 11 13 12 9 10 2
9 1 9 9 13 11 11 11 3 2
18 15 13 3 0 9 1 0 11 2 7 0 11 11 2 15 13 9 2
14 11 11 11 9 4 13 1 16 9 9 13 1 9 2
9 2 9 13 1 10 9 1 15 2
16 15 13 3 0 1 3 15 4 4 13 2 13 11 1 11 2
8 9 4 13 1 9 1 9 2
24 2 1 10 9 13 15 10 10 1 0 14 13 3 12 7 10 0 9 1 9 0 1 9 2
25 15 13 3 0 1 16 15 13 0 2 7 15 4 3 13 2 13 11 2 15 3 4 13 0 2
8 2 15 4 3 13 0 9 2
18 10 0 12 9 4 15 1 0 13 1 1 9 1 12 9 1 9 2
16 1 9 9 13 11 16 15 13 10 0 9 1 14 13 9 2
8 1 9 13 15 3 3 1 2
20 1 10 0 9 1 9 13 15 0 1 11 2 7 15 13 3 3 1 9 2
14 2 10 0 12 0 9 13 0 2 7 9 13 0 2
32 1 1 0 9 13 15 10 9 1 14 13 1 11 2 7 15 13 15 15 13 2 7 15 13 3 0 2 13 9 1 11 2
17 11 11 13 10 12 15 13 0 0 2 7 13 9 1 9 12 2
23 11 11 13 9 12 2 11 11 12 2 16 11 11 11 11 13 1 1 3 0 7 9 2
6 11 13 1 12 9 5
4 13 1 9 2
15 0 11 11 13 10 0 9 1 9 1 9 1 11 9 2
10 11 11 13 15 1 1 9 1 9 2
18 9 11 13 0 3 1 9 7 13 12 9 9 1 11 11 1 9 2
12 11 13 1 9 7 13 3 9 12 1 9 2
20 15 13 12 9 1 11 2 7 13 10 0 9 7 13 1 9 1 9 12 2
11 1 9 13 15 12 9 1 10 0 9 2
8 11 11 1 11 13 9 12 2
7 15 13 12 9 1 11 2
8 0 11 11 11 13 1 9 2
16 11 11 13 3 0 0 1 9 2 16 11 11 13 1 9 2
32 11 11 13 9 12 2 11 11 9 12 2 11 11 9 12 2 11 11 11 9 12 2 11 11 9 12 7 11 11 9 12 2
6 11 11 13 15 1 5
4 13 1 9 2
3 12 9 2
10 11 11 13 3 0 0 2 1 9 2
16 1 9 13 15 0 2 7 1 9 13 3 11 11 3 0 2
18 9 13 12 9 2 7 13 3 0 1 0 11 11 2 15 13 0 2
7 11 13 12 9 1 9 2
11 1 9 1 9 13 15 1 1 9 12 2
26 1 14 4 13 1 15 12 9 1 10 12 0 0 2 7 12 9 1 0 0 2 13 9 10 9 2
18 1 9 13 11 11 7 11 11 1 0 9 2 1 3 10 7 9 2
14 0 1 11 13 11 11 12 0 9 1 10 12 0 2
15 11 13 3 12 9 2 7 9 1 9 13 3 1 9 2
6 11 1 0 1 11 5
4 2 13 9 2
10 11 11 13 9 1 9 1 11 9 2
8 11 11 13 0 9 1 9 2
15 2 15 13 3 12 9 9 7 0 1 9 1 10 9 2
15 15 13 0 9 2 7 9 13 0 3 0 2 13 9 2
10 11 11 11 13 3 10 0 0 9 2
14 9 4 13 1 10 0 9 2 7 13 15 9 9 2
6 9 13 15 9 12 2
5 2 15 13 0 2
14 15 13 1 10 9 2 13 11 1 11 1 9 9 2
22 11 13 1 9 1 10 9 1 12 9 2 15 13 9 1 11 11 9 1 9 9 2
17 1 9 13 9 1 12 9 7 13 12 9 1 11 11 1 11 2
19 11 13 9 12 1 0 9 2 7 13 10 9 1 10 9 1 12 9 2
7 15 13 12 9 1 9 2
17 11 11 11 13 3 0 0 1 9 2 16 11 11 13 9 12 2
13 11 11 11 13 1 9 7 11 11 13 9 12 2
13 11 11 11 13 9 12 7 13 15 3 1 9 2
6 2 11 4 13 0 5
4 11 13 9 2
2 13 2
12 9 11 11 11 13 11 11 11 4 13 0 2
19 9 11 11 11 13 0 1 9 1 11 11 11 1 9 12 9 1 11 2
18 9 1 11 4 13 1 10 0 7 13 15 0 1 1 9 1 9 2
13 0 1 9 4 13 1 11 1 9 9 1 11 2
13 9 13 11 9 12 2 7 9 13 15 10 9 2
15 3 13 9 3 1 16 9 4 13 0 1 10 0 9 2
25 2 16 15 13 3 2 13 15 1 9 9 16 15 3 13 1 2 13 11 11 11 1 9 9 2
15 1 9 1 9 1 3 0 11 4 13 2 13 11 3 2
6 2 15 4 13 0 2
13 3 13 9 0 7 0 0 1 9 9 1 9 2
6 2 15 4 15 13 2
4 15 13 0 2
12 15 4 13 1 10 9 2 13 11 1 11 2
3 13 9 5
10 3 13 11 1 14 13 9 1 9 2
20 2 9 1 9 13 14 13 9 2 7 9 1 9 13 14 13 15 1 9 2
12 3 4 15 3 13 9 0 0 2 13 15 2
15 9 11 11 2 15 13 9 12 9 2 13 3 1 11 2
9 2 15 13 3 0 2 7 0 2
26 15 4 13 15 1 0 9 7 9 2 7 15 13 3 10 9 16 15 4 13 2 13 11 1 11 2
15 2 0 1 11 2 13 11 11 2 15 13 9 12 9 2
17 3 13 11 0 0 1 14 4 13 1 1 10 9 15 13 0 2
25 2 9 13 15 14 13 1 9 2 7 15 13 0 1 15 14 4 13 1 10 0 2 13 15 2
8 11 11 13 11 1 12 9 5
8 7 13 1 9 1 11 11 2
17 11 11 13 15 9 1 2 11 2 1 9 16 9 4 13 9 2
10 11 13 3 16 9 4 13 9 1 2
21 9 9 13 1 1 1 9 1 10 0 9 13 12 9 2 7 1 9 12 9 2
22 2 11 13 10 0 9 2 7 15 4 13 10 9 16 15 4 4 13 1 1 9 2
16 3 13 15 1 16 15 4 13 9 2 13 11 1 11 11 2
19 9 1 10 0 9 2 10 0 9 2 4 9 13 1 9 1 12 9 2
13 9 1 10 0 9 11 4 13 9 12 9 9 2
26 15 4 13 1 12 9 2 7 12 9 13 1 14 13 1 1 9 1 9 1 9 1 10 0 9 2
19 2 11 2 4 13 1 9 1 9 1 9 1 16 10 0 9 4 13 2
11 10 0 7 0 0 9 4 3 13 3 2
16 9 4 13 1 9 7 9 1 0 1 10 0 9 1 9 2
29 9 2 10 0 9 11 11 2 13 2 11 2 10 0 9 15 13 1 0 9 7 15 4 13 1 0 0 9 2
13 2 0 9 1 14 13 10 9 2 9 7 9 2
26 2 11 2 13 0 1 10 0 9 2 7 13 1 2 11 2 1 11 9 11 2 13 15 1 9 2
6 10 9 1 0 11 5
6 11 11 1 9 3 2
27 11 11 11 13 7 9 7 9 1 11 11 2 10 10 9 15 13 7 13 7 15 10 7 10 9 1 2
18 1 9 13 15 9 2 7 3 1 9 13 15 9 1 10 0 9 2
36 2 15 13 3 0 0 2 13 11 11 1 11 1 9 0 0 9 2 7 13 15 4 13 0 14 13 3 10 12 0 9 1 10 0 9 2
6 15 13 15 3 3 2
22 11 11 13 9 15 13 12 9 1 2 7 1 9 13 11 3 12 9 1 11 11 2
11 3 1 10 15 13 11 11 9 1 11 2
5 13 0 1 9 5
22 2 3 1 10 9 13 15 0 14 13 1 9 1 9 1 10 12 9 0 1 9 2
21 15 4 15 13 1 2 10 12 10 9 13 0 0 2 13 11 11 11 1 11 2
14 2 15 4 13 10 9 2 15 4 13 0 1 9 2
17 3 13 11 11 9 1 12 9 1 11 11 12 9 7 10 9 2
9 10 0 9 1 10 0 9 3 2
11 10 0 9 4 13 1 11 11 0 9 2
17 11 13 1 0 9 1 0 2 7 13 1 1 0 9 1 0 2
18 10 9 13 0 16 11 13 15 1 0 12 9 7 13 9 1 15 2
17 11 11 13 11 9 1 9 2 7 13 3 0 1 9 9 13 2
19 2 15 13 0 0 2 15 13 1 9 10 7 15 13 0 0 1 9 2
6 7 15 13 3 0 2
11 11 13 10 0 0 9 2 13 11 11 2
6 13 11 4 13 1 5
23 11 9 13 9 0 2 7 1 10 9 13 15 10 0 9 10 9 16 15 13 1 9 2
20 2 15 13 11 4 13 15 10 9 7 13 15 9 1 2 13 11 1 11 2
20 11 11 13 3 3 12 9 1 0 11 15 0 3 13 3 0 9 1 9 2
8 3 15 13 3 9 11 11 2
15 2 15 13 0 0 15 15 13 2 7 15 13 3 0 2
23 15 13 3 3 3 0 15 13 15 2 7 11 13 0 9 1 9 1 9 1 11 3 2
13 1 15 4 15 13 0 0 1 9 2 13 11 2
17 2 15 13 3 14 13 15 1 10 9 2 3 13 15 9 3 2
14 3 4 15 13 0 16 15 13 11 15 13 1 11 2
4 9 1 11 5
6 13 12 9 1 11 2
11 11 13 1 9 1 11 1 11 11 9 2
25 1 12 9 13 15 12 2 12 1 11 2 11 2 11 9 2 7 3 13 11 15 4 13 3 2
17 1 9 4 11 13 9 7 10 12 9 13 1 1 12 2 12 2
16 1 9 13 15 0 16 9 11 11 4 13 1 9 1 9 2
8 3 13 11 0 9 1 9 2
21 15 13 12 9 1 1 11 11 2 15 13 11 11 1 12 2 12 1 9 9 2
25 11 1 9 13 3 10 0 9 2 7 9 13 15 0 0 9 1 12 2 12 1 11 1 11 2
18 9 4 13 1 1 10 0 9 7 13 9 1 11 1 12 2 12 2
26 1 9 1 11 7 11 13 15 1 9 11 11 15 13 1 10 0 9 1 16 9 3 13 10 9 2
9 15 13 12 2 12 1 12 9 2
5 11 13 1 11 5
6 13 9 12 1 10 2
29 11 13 1 1 14 13 3 10 0 9 1 9 1 11 2 7 13 1 0 9 7 13 12 2 12 1 11 9 2
32 2 15 13 0 0 1 12 9 2 7 3 13 15 10 9 0 9 1 2 0 1 9 1 0 9 2 13 11 9 11 11 2
8 15 13 11 9 1 12 9 2
17 3 11 11 2 11 11 2 11 11 7 11 11 13 15 1 9 2
10 7 15 13 3 3 1 9 1 9 2
20 1 12 0 9 2 12 2 12 2 12 2 12 2 13 11 0 0 1 9 2
9 9 13 10 0 9 12 2 12 2
12 9 13 11 11 12 2 12 1 10 0 9 2
4 9 13 11 2
35 2 15 13 0 3 3 11 13 14 13 1 9 1 10 0 13 16 15 1 3 4 13 1 14 13 9 1 15 1 3 2 13 11 11 2
15 9 4 13 15 0 0 1 11 9 1 9 9 1 9 2
24 3 13 15 1 9 1 15 15 13 13 9 1 9 15 10 0 12 9 4 13 9 1 9 2
10 2 11 4 13 9 1 11 1 12 2
13 15 13 10 0 9 15 4 13 1 9 1 11 2
14 3 13 15 1 15 7 10 10 2 1 9 1 9 2
16 15 13 15 1 10 9 3 16 15 13 1 9 2 13 15 2
2 9 5
34 9 13 1 1 14 13 10 0 9 1 9 9 2 7 3 4 11 4 13 0 9 1 16 9 1 9 1 0 9 3 3 4 13 2
35 11 13 16 15 3 13 0 9 1 9 2 7 13 15 3 1 13 0 9 1 11 15 13 9 1 16 9 1 0 9 3 3 4 13 2
21 2 15 4 13 1 12 9 0 1 9 1 15 11 11 13 1 10 9 1 9 2
25 7 15 13 9 10 15 13 9 2 7 1 9 1 9 13 15 16 11 7 11 3 13 10 0 2
11 15 4 15 3 13 9 1 2 13 15 2
30 16 0 11 10 0 12 9 4 13 10 9 1 9 1 0 11 2 4 0 11 13 1 1 12 9 9 10 0 9 2
22 9 13 15 1 9 4 13 15 1 10 9 1 0 9 1 14 13 1 9 1 9 2
22 2 15 13 3 9 2 7 15 13 16 9 13 16 0 9 3 13 9 2 13 15 2
3 10 9 5
17 11 13 3 9 1 16 9 13 10 0 9 1 11 1 9 9 2
9 2 0 9 13 10 10 0 9 2
28 15 13 3 15 4 13 10 0 9 2 7 15 4 13 9 1 9 1 15 15 13 15 1 12 2 13 15 2
10 7 9 13 1 9 16 9 13 9 2
17 2 15 13 3 10 9 3 16 15 3 13 0 14 13 1 9 2
29 16 11 4 13 0 9 1 15 15 13 0 1 1 2 13 15 0 14 13 1 1 0 9 1 9 2 13 15 2
20 11 13 3 16 3 0 9 4 13 10 9 1 9 1 14 13 1 1 9 2
13 2 15 13 0 9 3 1 0 9 16 15 13 2
22 7 15 13 0 1 14 13 10 0 9 1 14 13 1 9 2 9 7 9 1 9 2
5 15 13 3 9 2
3 10 9 5
3 9 9 5
34 9 1 15 15 4 13 10 0 9 1 9 1 9 13 0 9 2 7 1 9 9 13 9 1 11 11 11 2 11 2 9 1 9 2
24 1 9 1 16 9 13 10 9 1 3 0 9 15 4 13 1 10 0 9 2 13 15 0 2
32 2 10 0 9 4 1 10 7 10 9 4 13 1 9 16 0 9 13 2 7 15 13 3 1 9 1 14 13 3 3 2 2
22 1 9 1 16 9 13 10 9 9 16 9 1 9 13 1 9 2 13 9 3 0 2
2 6 2
16 1 12 13 10 0 1 11 2 0 0 9 2 1 12 9 2
20 9 4 3 13 1 12 9 2 7 0 13 1 16 10 0 9 13 3 0 2
14 7 15 4 3 13 10 9 2 13 15 15 13 4 2
30 5 9 1 9 0 1 11 13 0 0 0 2 7 0 0 1 1 13 15 13 9 1 14 13 9 9 15 4 13 2
24 9 13 3 1 3 0 0 9 0 13 1 14 13 9 11 13 1 14 13 1 1 9 1 2
8 16 11 11 13 1 0 9 2
12 2 8 8 8 8 8 8 8 8 8 2 2
18 9 1 11 13 14 13 10 0 0 9 15 4 13 0 12 10 9 2
20 11 4 13 12 9 2 7 1 12 4 13 1 1 10 0 2 1 10 11 2
18 10 0 9 9 4 13 10 9 0 2 7 9 4 13 0 1 12 2
21 10 9 4 13 2 0 1 12 2 7 9 1 9 13 1 11 11 0 1 13 2
18 9 13 16 3 9 11 11 3 13 16 15 4 13 1 1 9 9 2
17 5 1 9 1 15 13 15 0 14 13 1 11 0 9 1 11 2
27 15 13 13 10 9 1 3 0 9 15 4 13 1 10 9 2 7 15 4 13 9 1 9 9 1 11 2
3 0 9 5
3 9 9 5
24 1 9 7 9 1 12 13 15 1 0 9 1 12 9 1 9 1 12 9 13 1 10 9 2
13 3 13 9 0 0 2 3 12 9 1 9 13 2
6 9 1 9 13 0 2
35 9 1 11 1 11 2 11 1 11 7 11 1 11 13 10 1 12 9 9 2 16 11 7 11 1 11 13 0 2 1 12 7 12 9 2
20 9 1 11 2 11 11 11 2 13 1 11 16 15 13 0 1 9 0 9 2
19 11 4 3 13 1 14 4 13 1 1 9 1 0 9 7 9 1 9 2
35 2 8 8 8 8 8 8 8 8 8 8 8 2 8 8 8 8 8 8 8 8 8 8 8 8 8 8 8 8 8 8 8 8 8 2
19 8 8 8 8 8 8 8 2 8 8 8 8 8 8 2 2 13 11 2
35 15 13 1 9 1 11 4 13 1 9 2 7 1 9 1 10 0 9 1 14 13 2 7 3 16 15 4 13 0 9 1 10 0 9 2
18 15 13 3 0 1 16 9 7 0 9 1 15 10 13 1 0 9 2
11 15 13 3 1 16 9 13 1 0 9 2
20 3 0 15 13 9 1 0 9 2 3 0 4 15 13 4 4 13 1 9 2
36 15 4 3 13 16 9 13 9 1 1 10 9 9 13 16 10 9 13 15 7 16 9 0 13 1 9 1 14 13 9 1 10 9 9 13 2
21 3 13 10 0 9 1 9 2 0 1 9 2 16 9 7 9 13 9 7 9 2
27 10 0 9 1 0 9 7 9 15 9 13 14 13 1 1 9 2 13 1 9 10 9 1 9 7 9 2
22 3 0 4 9 13 10 9 16 3 10 0 9 3 4 13 1 9 1 10 0 9 2
4 2 11 0 5
3 10 9 2
8 10 0 11 4 13 1 9 2
15 7 9 4 3 13 0 1 9 9 2 13 11 11 11 2
6 16 9 4 13 15 2
8 9 13 9 1 10 0 11 2
19 9 11 11 11 13 16 0 1 11 0 9 4 4 13 1 9 1 9 2
2 9 2
7 11 11 2 11 5 11 5
18 2 7 11 2 9 2 7 11 4 13 0 1 14 13 9 1 9 2
21 9 4 13 0 1 9 7 9 2 13 9 7 9 11 11 11 1 11 1 11 2
23 11 0 9 11 11 13 1 10 9 11 11 2 9 1 9 1 16 15 4 13 1 9 2
12 10 0 9 2 11 2 13 9 10 10 9 2
30 2 16 15 4 13 15 3 4 15 13 15 1 9 7 13 1 15 2 13 11 11 2 9 7 9 1 9 2 9 2
22 9 4 13 10 9 1 12 9 9 7 9 1 15 15 13 11 7 13 15 1 9 2
4 9 1 9 5
9 9 4 13 10 0 9 1 9 2
17 9 4 13 0 1 14 13 1 9 2 3 16 11 3 13 9 2
14 2 9 4 3 3 13 10 9 1 9 2 13 11 2
15 1 9 1 9 9 13 9 3 0 9 1 10 0 9 2
24 0 10 9 13 11 10 9 1 14 13 9 1 9 15 13 1 2 9 2 7 2 9 2 2
12 11 13 10 0 9 13 10 0 9 1 9 2
13 2 15 4 13 0 14 13 11 9 1 9 3 2
19 9 4 0 9 13 15 15 3 4 13 9 2 16 11 4 13 1 9 2
17 16 15 4 13 9 2 13 15 15 1 14 13 9 2 13 11 2
5 13 9 1 11 5
15 9 13 9 3 9 1 9 11 2 12 9 1 1 11 2
18 11 13 11 9 7 10 1 0 9 3 10 0 9 3 13 1 9 2
16 3 13 9 10 0 7 0 1 9 1 9 13 11 10 9 2
18 9 4 13 9 7 13 9 16 15 4 13 15 1 9 1 12 9 2
19 9 0 9 4 13 14 13 1 9 1 9 1 9 1 9 1 0 9 2
10 9 4 13 9 10 1 14 13 9 2
13 3 4 15 13 1 9 1 9 0 9 1 9 2
14 2 13 15 9 1 14 13 9 1 11 9 1 11 2
7 2 6 2 15 13 15 2
14 1 11 4 15 13 1 0 9 1 9 1 11 9 2
10 11 13 10 0 9 1 0 0 9 2
18 16 9 13 9 1 9 10 1 9 1 15 4 9 13 2 13 11 2
12 2 10 9 13 3 0 9 2 15 13 9 2
13 15 13 3 16 0 4 4 13 2 0 3 0 2
28 7 15 4 3 13 3 2 15 13 10 9 1 16 15 13 15 2 13 10 1 9 9 2 11 11 11 9 2
5 0 9 1 11 5
13 1 11 13 0 0 16 9 1 9 3 13 15 2
10 0 9 4 13 1 9 1 0 9 2
10 0 4 0 9 1 9 1 9 13 2
18 3 1 9 13 15 0 9 1 10 9 1 9 7 10 0 9 0 2
19 9 1 9 13 15 15 13 1 14 3 13 1 0 9 1 9 1 9 2
13 7 13 15 13 10 0 1 14 13 9 1 11 2
20 3 4 15 13 1 15 3 2 7 7 9 2 9 7 9 13 9 1 15 2
12 9 1 9 4 13 10 0 9 1 10 9 2
18 15 4 13 10 9 7 0 1 7 16 15 13 9 7 9 1 9 2
44 16 10 1 9 1 11 11 4 4 13 1 10 9 13 1 9 1 9 1 10 0 9 15 15 1 7 1 15 4 13 16 15 13 9 4 10 0 9 3 13 0 1 15 2
46 10 9 4 3 13 10 0 9 1 9 1 9 15 9 13 1 9 2 7 15 13 0 0 9 1 14 13 1 1 9 1 9 1 9 1 15 15 4 13 1 9 1 9 7 9 2
21 9 13 3 1 16 9 9 4 0 0 13 1 9 7 9 1 1 10 0 9 2
33 15 4 0 13 9 1 14 13 10 9 15 0 13 1 0 16 9 4 13 10 10 9 1 0 9 16 15 13 1 1 1 9 2
19 15 4 1 9 3 13 16 11 11 4 13 1 10 0 0 9 1 9 2
20 16 0 9 0 13 0 2 13 3 14 13 16 11 11 4 4 13 1 9 2
40 1 9 1 9 13 9 1 9 16 10 9 3 9 13 0 1 11 9 2 3 1 9 2 4 13 1 0 9 1 11 11 2 7 3 13 1 9 1 9 2
6 12 9 1 0 9 5
18 9 13 0 9 1 0 9 1 11 11 2 7 1 0 7 0 9 2
11 9 13 3 16 15 4 13 10 0 9 2
27 0 13 9 9 1 16 15 0 13 9 1 0 9 1 11 7 11 11 2 15 3 3 13 1 11 11 2
29 9 1 9 13 0 1 11 2 7 15 13 10 9 1 15 15 13 15 1 7 0 3 13 9 1 9 1 11 2
13 10 10 9 1 11 11 4 1 10 9 13 0 2
21 0 4 9 1 0 13 16 15 13 0 10 9 9 13 1 14 13 9 1 9 2
44 1 9 13 16 15 0 16 15 13 10 3 0 7 0 9 1 11 11 4 13 9 1 14 13 9 1 14 13 16 10 0 9 4 13 0 9 7 13 0 9 7 0 9 2
24 15 13 3 0 16 9 9 13 9 1 14 13 10 3 9 7 9 1 9 15 3 13 0 2
18 15 13 10 9 1 9 16 10 0 9 3 13 0 9 1 1 12 2
27 0 9 13 3 1 16 9 4 13 1 12 2 3 0 1 9 1 10 9 11 11 13 1 10 10 9 2
30 9 4 3 13 9 1 1 0 14 13 10 9 1 10 0 0 9 2 11 11 2 2 15 13 1 1 9 1 12 2
27 3 4 15 1 3 0 13 10 9 1 9 1 11 1 11 2 15 4 13 1 10 0 0 9 1 12 2
9 12 9 1 0 9 1 11 11 5
12 10 0 9 1 11 11 4 13 1 0 9 2
36 1 9 1 0 9 1 0 9 1 11 7 11 11 1 10 9 1 11 11 1 14 13 9 1 11 11 1 10 0 9 1 9 1 11 9 2
16 10 9 1 10 0 9 1 11 11 4 13 0 7 0 0 2
30 1 10 9 4 10 9 13 16 9 1 9 13 0 1 15 15 9 13 1 11 2 7 15 13 15 1 10 0 9 2
21 10 0 0 9 3 1 11 11 4 1 9 9 13 9 1 10 0 9 3 3 2
16 9 7 9 1 11 11 13 0 1 0 1 11 1 1 9 2
34 13 15 9 1 11 11 2 4 15 13 16 15 3 13 10 0 9 1 9 2 7 0 9 1 9 4 13 0 1 9 1 11 11 2
33 15 4 13 10 3 0 0 9 14 13 1 15 1 14 13 9 1 10 9 1 9 15 3 13 7 4 13 2 0 1 0 9 2
23 15 13 3 0 9 1 11 7 11 11 16 15 13 0 9 2 0 9 2 9 7 9 2
34 9 1 9 1 10 9 1 11 4 3 13 1 9 1 11 11 2 7 1 10 9 4 15 13 0 1 9 1 11 11 13 1 11 2
16 1 10 9 13 15 0 1 10 0 9 1 11 7 11 11 2
23 10 10 9 1 9 1 11 11 13 1 10 10 9 15 0 1 9 1 9 9 7 9 2
37 1 10 9 4 9 1 9 13 16 9 1 11 11 3 0 1 9 13 1 10 0 9 7 16 11 9 13 10 0 9 1 14 13 10 10 9 2
8 12 9 1 9 1 11 11 5
35 9 13 16 10 0 2 0 9 1 11 11 3 7 0 4 13 9 2 9 7 9 2 15 1 9 13 10 12 0 0 9 1 11 11 2
25 1 9 4 15 13 9 1 14 13 1 9 1 9 1 9 7 9 3 2 16 10 9 4 13 2
37 16 9 13 10 0 9 1 11 13 1 0 9 2 13 15 15 3 0 16 9 1 7 9 1 10 9 13 1 9 1 9 1 9 1 11 11 2
27 1 0 9 4 15 3 13 0 14 13 9 1 9 1 11 11 7 13 9 15 9 13 1 9 1 11 2
20 15 13 3 0 16 9 9 1 9 3 4 13 1 1 10 9 1 11 11 2
9 10 10 13 1 9 1 11 9 2
24 9 13 3 16 15 13 0 9 1 14 13 1 10 0 9 1 9 1 10 9 1 11 11 2
39 15 4 3 13 9 1 14 13 16 15 4 13 0 9 1 11 11 2 1 0 9 1 9 7 1 14 13 0 9 2 0 10 9 3 9 13 0 2 2
33 7 10 9 4 13 1 9 0 1 10 0 9 15 9 13 1 11 9 9 12 0 9 2 1 16 15 13 10 0 9 1 9 2
4 9 1 9 5
2 9 5
11 15 4 0 13 9 1 10 9 1 9 2
7 3 13 0 9 1 11 2
28 15 4 3 13 9 1 16 10 9 1 10 9 13 0 2 3 16 9 1 9 13 9 1 9 1 0 9 2
52 3 2 3 13 15 16 9 4 13 10 9 0 0 1 1 9 1 14 13 10 9 1 1 11 2 3 11 2 1 14 13 9 1 10 9 16 3 11 9 1 10 9 1 9 13 14 13 1 10 0 9 2
18 15 4 13 10 0 3 2 7 3 13 1 1 3 10 9 13 0 2
38 10 0 11 13 16 15 13 1 1 11 2 13 14 13 1 9 7 13 1 16 9 1 9 1 4 13 2 0 16 15 13 0 1 11 5 11 9 2
36 15 13 16 10 0 9 1 16 11 13 1 9 2 13 16 15 1 14 4 13 10 9 13 16 10 0 9 3 4 13 0 0 1 10 9 2
40 11 13 16 16 15 4 13 1 3 0 9 1 11 5 11 2 3 4 9 13 3 0 2 7 3 0 1 11 15 13 0 1 0 9 2 16 9 13 0 2
20 15 4 3 3 13 10 0 9 1 16 10 9 1 9 1 10 9 13 0 2
20 1 0 9 3 2 3 13 11 5 11 1 14 13 0 9 1 9 1 11 2
11 15 13 9 1 9 1 10 10 0 9 2
16 9 13 16 9 3 13 3 0 2 7 0 0 1 1 11 2
33 9 1 15 13 9 1 11 5 11 15 4 13 1 1 0 9 3 2 3 15 3 13 1 11 16 15 13 9 1 0 12 9 2
26 3 13 9 1 11 2 16 9 1 10 0 9 1 11 2 13 3 0 0 9 1 11 7 0 11 2
27 1 10 10 9 3 13 3 9 16 16 15 3 13 9 1 10 0 9 1 12 2 3 4 15 4 13 2
27 16 15 13 2 3 4 0 0 0 1 10 0 1 0 9 13 0 9 1 1 11 1 11 2 11 3 2
34 15 4 3 0 0 3 13 1 9 1 14 13 9 1 11 2 7 15 13 3 16 15 4 13 15 1 10 9 3 15 3 13 9 2
6 15 4 13 15 1 2
41 9 13 0 1 16 9 2 4 4 13 12 9 1 9 7 9 2 7 10 0 9 1 9 2 9 7 9 2 1 16 15 13 0 1 14 13 10 0 1 9 2
13 15 4 13 15 1 9 2 3 13 15 0 9 2
38 15 4 3 13 1 9 1 10 1 9 1 11 1 0 9 3 2 3 9 13 0 1 9 1 10 9 2 3 1 9 1 0 9 1 9 7 9 2
9 10 0 9 1 9 4 13 10 2
5 9 13 3 0 2
24 13 9 1 9 2 3 16 0 9 13 0 1 10 0 9 2 3 10 1 10 0 0 9 2
19 3 15 1 7 1 4 13 9 1 11 0 1 10 7 0 9 1 11 2
8 9 13 9 2 7 0 9 2
4 9 1 11 5
13 11 11 11 13 1 9 7 9 1 11 12 9 2
14 15 13 11 1 14 13 9 7 13 15 1 0 9 2
18 11 13 3 1 10 9 15 4 13 1 14 13 9 1 11 7 11 2
37 15 13 1 10 9 1 9 15 4 13 9 1 9 1 9 1 14 13 10 9 15 13 1 1 2 1 0 0 9 2 1 14 13 1 0 9 2
17 11 7 11 13 9 15 13 9 7 9 1 9 15 13 1 11 2
14 9 13 9 1 14 13 9 7 9 1 1 9 10 2
20 9 1 11 7 11 13 3 16 15 13 1 9 1 9 10 1 0 0 9 2
33 15 13 3 14 13 16 15 13 11 0 9 1 9 10 7 3 4 13 1 1 12 2 12 2 9 0 1 9 16 15 13 9 2
12 7 4 15 13 10 16 9 13 9 1 9 2
19 0 9 4 0 15 2 15 13 9 1 3 1 1 1 1 10 0 9 2
5 11 13 0 9 2
10 10 9 13 0 9 1 9 7 9 2
9 3 3 1 9 2 7 1 9 2
28 15 13 15 1 9 2 9 7 9 1 9 2 3 1 9 1 9 15 3 13 15 1 0 9 1 0 9 2
8 1 11 13 9 3 0 1 2
13 1 10 9 1 11 9 13 1 9 1 10 9 2
13 15 13 9 15 15 1 9 3 4 13 13 0 2
15 3 4 11 13 0 1 1 14 13 1 10 9 1 9 2
35 11 13 10 9 1 9 1 11 2 15 2 1 0 9 1 11 2 13 12 0 9 1 0 11 2 7 0 3 0 9 15 12 9 13 2
13 0 9 1 10 0 9 13 1 9 0 1 9 2
28 16 15 4 13 9 1 10 0 9 4 9 13 0 9 9 2 7 13 16 15 13 14 13 0 7 0 9 2
9 7 15 4 13 9 1 0 9 2
5 9 13 0 9 2
9 11 9 4 1 9 13 1 9 2
26 11 9 9 13 9 1 10 0 0 9 1 9 2 3 1 9 7 9 2 9 2 9 5 9 3 2
28 0 1 10 0 0 9 13 15 1 9 1 9 2 1 9 4 11 11 9 13 9 1 9 1 1 10 11 2
16 1 9 13 11 12 9 9 2 7 1 12 9 1 0 9 2
15 11 4 1 0 9 13 10 9 1 1 12 9 1 12 2
16 10 0 9 1 9 1 11 4 13 1 12 0 9 1 12 2
4 15 13 0 2
49 9 11 13 16 2 0 9 1 9 4 13 12 2 12 0 9 1 9 2 2 0 9 12 2 7 13 1 9 1 9 1 9 15 13 16 15 4 3 13 9 1 9 13 1 9 3 1 9 2
41 0 12 9 1 10 0 9 1 9 4 13 1 9 2 7 16 0 13 1 1 9 4 15 13 0 9 9 2 13 9 1 9 1 9 7 3 13 0 1 9 2
21 11 9 13 16 15 13 10 9 0 15 1 11 7 13 10 0 9 13 1 9 2
13 15 1 9 4 13 9 1 0 1 10 0 9 2
15 9 2 9 2 9 7 9 13 14 13 9 15 13 1 2
32 1 15 13 15 10 9 16 0 7 9 1 11 7 11 13 16 16 15 13 0 7 13 1 0 9 3 4 9 13 1 9 2
7 3 3 1 10 0 9 2
6 11 13 9 1 9 5
29 11 11 2 11 0 0 9 2 4 13 9 1 1 9 7 13 1 0 1 0 9 1 9 1 9 7 0 9 2
19 11 4 0 13 9 1 14 13 15 15 13 7 13 1 15 15 13 1 2
16 9 4 3 13 14 13 15 15 13 0 9 1 9 1 9 2
16 9 1 9 15 4 13 0 1 0 4 3 13 1 10 9 2
30 7 16 11 1 0 13 9 1 1 10 3 0 9 2 13 15 15 9 4 13 0 1 14 13 15 10 9 15 13 2
29 1 9 1 10 9 15 13 7 1 14 13 1 10 0 9 2 4 15 3 13 1 14 13 9 1 9 15 13 2
15 15 4 3 13 11 9 1 14 13 10 0 9 1 9 2
19 11 13 10 9 1 9 9 7 13 16 10 0 9 4 13 1 9 10 2
32 15 4 13 9 9 1 0 9 1 12 9 16 15 13 0 14 13 1 1 9 9 1 14 13 15 1 10 0 9 1 9 2
24 0 13 15 16 9 2 1 9 7 9 2 4 13 1 16 0 9 13 15 0 14 13 9 2
6 6 1 10 0 9 5
13 2 1 9 13 11 11 10 0 0 9 1 9 2
29 0 9 11 11 7 10 3 0 9 2 11 11 11 11 2 13 1 9 1 11 3 1 0 9 1 11 7 11 2
15 9 4 3 13 1 10 0 9 2 7 4 13 1 9 2
8 3 13 10 9 0 0 2 5
15 10 0 9 4 11 13 0 1 9 1 0 9 1 9 2
21 9 4 3 13 0 1 9 1 9 1 9 7 9 2 7 10 9 4 4 13 2
28 16 0 9 3 13 1 9 1 14 13 9 1 9 1 9 3 13 15 10 9 1 9 7 9 15 13 9 2
10 9 13 3 1 16 15 13 0 9 2
3 0 9 2
25 15 15 0 4 13 9 1 0 9 13 16 9 13 3 1 14 13 9 1 10 0 9 1 11 2
20 1 9 11 13 10 9 12 9 0 2 7 9 1 10 9 1 12 9 9 2
25 9 1 11 4 13 12 9 0 16 15 3 4 4 4 13 16 9 13 9 1 9 1 10 9 2
22 1 9 13 0 9 0 9 1 10 9 1 9 1 16 15 4 13 1 9 1 11 2
29 15 13 15 0 9 0 4 13 9 1 2 7 15 15 9 4 13 9 1 1 12 9 1 14 4 4 13 0 2
3 0 9 5
19 1 9 1 9 13 9 1 9 1 10 0 9 1 3 12 9 9 0 2
6 1 9 13 9 12 2
9 15 13 3 10 9 1 0 9 2
21 15 13 15 0 1 2 7 3 4 15 3 13 1 0 1 16 15 4 13 0 2
22 9 13 3 15 16 15 13 1 16 9 4 13 3 1 0 9 1 9 3 1 9 2
7 10 9 13 9 1 12 2
16 9 1 9 13 16 9 1 9 1 9 13 1 1 12 9 2
11 15 4 13 16 15 13 0 9 1 9 2
20 10 0 9 13 1 16 9 1 1 9 13 0 7 16 9 1 9 4 13 2
3 0 9 5
14 15 4 7 11 2 11 7 11 13 16 15 13 1 2
23 11 7 11 4 13 16 15 4 13 9 2 7 13 1 16 10 0 9 4 13 0 9 2
25 1 10 0 13 15 3 1 10 0 9 2 7 14 13 9 1 9 1 10 0 9 3 1 9 2
18 1 10 0 13 3 10 0 9 9 10 9 1 15 15 4 13 9 2
21 9 13 3 0 0 16 15 13 1 2 7 10 9 13 1 10 0 9 1 9 2
2 9 2
13 0 9 13 3 1 9 1 10 0 9 1 9 2
7 13 15 3 13 0 0 2
10 9 13 10 0 9 1 9 1 9 2
24 15 13 3 10 9 1 9 16 9 1 1 13 3 0 0 9 1 15 15 13 1 1 1 2
22 1 9 13 15 0 14 13 9 1 9 1 2 16 15 13 0 0 14 13 10 9 2
17 1 9 13 15 9 15 13 1 9 1 7 15 13 1 9 1 2
44 15 13 9 1 9 15 4 4 13 14 13 9 5 9 1 11 11 16 15 13 0 0 1 10 9 14 13 10 9 13 15 1 1 10 9 3 16 15 4 13 10 0 9 2
7 15 13 0 7 0 0 2
16 15 4 13 0 9 1 10 0 9 1 11 1 9 7 9 2
3 9 13 5
24 9 1 10 0 9 13 0 1 1 0 2 3 0 16 10 0 9 3 13 1 10 0 9 2
27 1 10 0 9 4 11 13 10 0 9 1 0 9 1 9 2 15 13 0 0 16 10 9 4 13 0 2
37 16 1 12 9 1 9 13 0 2 13 1 0 9 2 13 15 3 0 7 0 16 15 13 0 1 10 12 9 15 15 4 13 1 9 1 3 2
7 7 15 13 9 1 9 2
8 15 13 0 1 9 1 9 2
14 15 13 1 9 1 9 7 9 2 7 13 1 9 2
13 9 13 1 12 9 1 9 1 10 9 1 9 2
24 3 13 15 1 9 16 9 13 15 1 9 1 14 13 1 0 9 7 13 10 9 1 9 2
17 15 13 0 0 1 10 9 16 15 13 10 9 1 9 1 9 2
7 3 4 15 13 9 1 2
8 15 13 16 15 13 1 15 2
12 15 13 0 14 13 2 7 3 1 0 9 2
6 9 2 9 2 9 2
15 3 13 9 1 9 3 7 9 1 1 9 13 1 3 2
18 9 1 1 2 9 7 9 13 3 9 1 9 1 10 9 7 9 2
16 9 2 9 2 7 0 9 13 9 1 0 0 9 1 11 2
16 0 9 4 3 13 9 1 10 0 0 9 1 14 13 9 2
13 15 13 14 13 14 13 1 9 1 1 12 9 2
15 3 13 16 9 13 1 9 1 14 13 9 1 12 9 2
9 15 13 3 0 1 10 0 9 2
7 3 4 9 9 13 0 2
7 15 13 3 3 10 9 2
11 9 13 1 0 9 16 9 13 0 9 2
31 0 9 13 0 9 7 15 13 0 16 15 13 9 15 13 9 7 9 1 14 13 15 16 9 4 13 1 9 1 9 2
7 9 13 1 9 1 9 5
29 10 9 13 1 9 16 9 2 11 2 9 1 9 13 1 9 1 10 9 1 10 9 1 11 1 11 7 11 2
25 2 10 9 4 13 2 7 9 13 1 9 2 13 9 11 11 1 11 11 2 11 2 1 11 2
17 15 13 12 9 1 9 1 9 2 11 2 2 7 12 1 9 2
19 9 1 9 4 0 13 1 9 1 9 2 0 15 12 9 13 1 9 2
28 10 12 1 15 2 11 2 11 2 2 13 1 15 9 15 13 2 7 13 1 9 9 9 1 9 1 11 2
15 9 13 1 10 9 1 10 9 1 9 1 9 1 9 2
8 2 15 13 3 9 1 9 2
20 15 13 0 9 1 9 2 7 1 0 0 9 1 9 1 9 2 13 11 2
8 11 13 9 1 9 9 12 2
4 2 11 2 5
6 13 0 9 1 11 5
19 11 7 9 4 13 9 1 16 0 11 11 9 3 4 13 0 0 9 2
14 9 1 11 13 16 9 1 10 0 9 3 4 13 2
31 1 10 9 1 9 9 13 11 11 9 1 16 15 3 4 13 0 9 1 9 7 9 13 1 9 1 0 9 1 11 2
20 0 13 9 16 9 12 1 0 11 11 9 4 13 1 9 1 11 11 9 2
14 1 9 4 9 3 13 10 0 9 1 9 1 9 2
19 9 4 13 0 9 2 9 1 9 2 0 9 7 0 9 2 13 11 2
20 2 3 4 9 13 2 7 15 13 10 0 9 14 13 1 15 16 15 13 2
23 15 13 3 0 16 15 4 13 1 10 9 1 9 2 13 0 9 11 11 1 11 11 2
6 2 15 13 3 3 2
18 15 4 4 13 10 0 0 9 7 13 14 13 3 1 10 0 9 2
13 1 14 13 9 1 10 0 9 2 4 9 13 2
30 9 13 14 13 10 9 1 9 1 14 13 9 2 15 15 13 10 9 1 9 2 13 9 1 11 2 11 11 11 2
4 2 11 2 5
13 10 9 13 9 1 15 7 0 9 1 0 9 2
9 1 14 13 9 4 0 9 13 2
8 3 4 0 9 13 7 13 2
12 3 4 15 13 9 0 9 2 9 7 9 2
17 15 13 1 9 16 15 4 13 9 1 0 7 0 9 7 9 2
6 10 9 4 13 1 2
19 15 4 13 9 1 10 0 9 1 9 2 15 15 13 0 9 1 9 2
17 9 1 9 1 0 9 4 13 1 16 9 1 0 9 4 13 2
10 15 4 13 10 0 0 9 1 9 2
12 11 4 13 0 1 14 13 1 9 7 9 2
7 15 13 0 9 1 9 2
10 10 9 13 12 12 0 0 1 9 2
9 3 4 15 13 0 10 0 9 2
7 9 4 13 10 0 9 2
21 11 4 13 1 0 1 0 9 1 0 9 1 0 9 7 9 1 10 0 9 2
11 15 13 3 9 7 9 1 0 0 9 2
8 9 0 9 13 10 0 9 2
9 3 4 11 13 1 9 7 9 2
13 3 13 15 9 7 1 9 7 1 9 1 9 2
9 15 4 13 7 13 9 1 11 2
17 11 4 13 0 9 1 9 7 0 9 15 4 13 9 0 9 2
17 15 4 13 1 0 9 7 13 9 1 11 2 7 0 7 0 2
17 0 4 15 13 1 9 1 10 9 16 11 13 9 7 0 9 2
11 11 13 1 9 1 10 0 9 1 9 2
30 15 4 13 0 9 2 13 1 9 1 12 12 9 1 0 9 12 7 13 9 1 9 1 9 16 0 9 4 13 2
11 11 13 10 0 9 2 15 13 9 9 2
10 15 4 3 13 9 1 9 0 9 2
14 11 4 13 1 10 0 9 1 14 13 9 1 11 2
17 15 4 13 0 1 1 9 2 3 16 0 4 13 1 10 9 2
12 15 4 13 0 9 1 9 15 13 1 9 2
9 10 0 9 4 13 1 1 9 2
7 11 13 0 9 1 9 2
18 15 4 13 1 9 1 0 9 7 9 1 0 9 2 0 7 0 2
23 15 4 13 10 9 15 13 9 2 13 0 9 7 13 1 0 1 9 1 9 7 9 2
11 15 4 13 15 0 14 13 0 1 9 2
10 15 4 13 9 9 1 9 7 9 2
6 11 4 13 1 9 2
14 15 4 13 10 0 0 9 1 11 7 10 0 9 2
5 11 13 10 9 2
19 15 13 0 9 7 0 9 9 13 1 9 2 9 7 9 1 0 9 2
5 15 4 13 9 2
17 15 4 13 1 0 0 9 2 7 15 4 13 9 1 10 9 2
10 15 4 13 9 15 13 9 1 9 2
33 11 4 13 1 16 10 0 9 1 9 15 13 1 0 9 2 13 1 9 1 2 1 9 2 9 7 9 2 1 10 0 9 2
10 11 4 13 0 1 0 9 1 9 2
12 9 4 13 1 9 1 9 1 9 1 9 2
10 15 4 13 1 0 1 9 7 9 2
24 11 4 13 1 16 9 1 14 13 10 0 9 1 9 1 11 13 2 7 13 0 1 15 2
11 1 11 10 4 15 3 13 9 1 9 2
37 16 10 0 9 13 2 4 15 1 10 0 9 1 11 7 1 2 13 11 2 13 10 9 15 4 13 2 7 10 9 15 3 4 13 9 1 2
24 15 4 13 1 0 1 16 11 4 13 10 1 10 0 2 0 2 0 7 0 9 1 9 2
18 9 7 0 9 1 9 13 1 10 9 1 9 2 9 7 10 0 2
6 10 0 9 4 13 2
20 15 4 13 0 9 1 9 1 0 9 2 0 9 2 9 2 9 7 9 2
19 15 13 10 9 1 11 14 13 1 0 1 0 9 1 0 9 1 11 2
15 9 13 10 0 9 1 9 2 9 7 9 1 0 9 2
7 11 4 13 9 1 9 2
18 9 1 10 0 9 4 13 1 10 9 1 9 7 1 9 7 9 2
15 11 4 13 10 0 9 1 14 13 1 0 1 0 9 2
18 1 0 9 7 9 1 9 4 10 0 9 1 9 1 0 9 13 2
14 15 4 13 0 9 7 1 0 9 13 9 0 9 2
24 15 4 13 10 0 9 1 0 9 7 13 9 9 7 0 9 1 9 1 10 9 1 9 2
7 11 4 13 10 0 9 2
21 15 4 13 1 9 10 0 9 1 14 13 9 1 10 9 15 4 13 1 9 2
9 15 4 13 12 0 9 1 11 2
17 11 4 13 9 1 10 9 1 14 13 10 0 7 0 0 9 2
34 11 13 10 0 7 0 9 1 10 9 1 10 0 9 1 0 9 2 7 4 13 10 0 9 1 14 13 1 10 0 9 1 9 2
20 1 12 4 15 13 10 0 9 1 10 9 1 12 9 9 1 9 0 9 2
10 9 1 9 13 1 10 0 0 9 2
11 3 4 15 13 10 0 0 9 1 9 2
15 15 13 14 13 0 2 13 0 2 13 0 7 13 0 2
13 11 4 13 10 9 1 0 9 1 9 1 9 2
19 15 4 13 9 1 9 7 9 10 0 9 2 0 15 15 13 0 9 2
30 1 10 9 16 10 3 0 13 15 0 13 0 2 4 15 3 3 13 15 14 13 1 2 7 3 15 14 13 1 2
11 15 4 3 13 9 7 9 9 1 9 2
11 11 4 13 1 0 9 1 9 7 9 2
9 15 4 13 10 0 7 0 9 2
18 15 4 13 1 11 1 10 9 1 9 1 12 9 1 9 1 12 2
17 15 4 13 1 0 1 16 11 0 9 13 10 0 7 0 9 2
18 15 4 13 1 1 10 0 9 1 9 7 9 1 9 1 9 9 2
33 11 13 14 13 15 9 1 14 13 10 9 2 0 1 9 2 9 2 0 9 2 9 2 0 9 2 9 2 9 7 0 9 2
9 3 4 15 13 10 9 1 9 2
28 15 4 13 9 1 9 7 0 9 2 7 13 1 16 11 13 0 9 1 9 15 13 0 1 10 0 9 2
13 11 4 13 10 0 9 15 13 1 0 0 9 2
16 10 0 9 7 9 4 13 1 10 9 15 15 13 1 12 2
12 9 1 9 1 9 4 13 1 9 1 9 2
23 3 0 15 13 1 14 13 10 9 2 4 13 1 10 0 9 15 13 1 0 0 9 2
21 9 1 0 9 2 0 9 2 0 0 7 0 9 13 0 9 1 11 0 9 2
12 11 4 13 1 10 0 9 3 1 0 9 2
33 3 4 15 13 9 15 4 13 1 11 1 9 2 3 16 15 4 13 7 10 0 0 9 7 10 9 15 9 4 13 1 9 2
27 16 15 1 12 9 3 4 13 16 11 1 12 4 13 10 1 9 3 0 9 2 4 15 13 1 15 2
10 1 11 4 15 13 7 0 7 0 2
18 15 4 13 9 10 0 2 7 15 4 13 1 10 0 9 1 9 2
10 13 15 3 13 10 0 9 11 13 2
54 10 9 13 14 13 11 3 0 2 10 0 9 14 13 1 1 2 10 0 9 14 13 2 13 7 13 15 1 7 10 0 9 14 13 0 1 1 0 9 2 0 15 15 3 13 0 2 7 13 15 3 0 0 2
9 11 13 10 9 1 11 1 15 2
11 15 13 3 16 15 4 13 15 15 13 2
3 3 1 2
16 15 13 1 10 0 9 1 14 13 11 0 10 10 12 9 2
7 10 9 4 13 15 3 2
31 15 13 16 9 1 10 9 13 1 0 9 7 9 2 0 1 0 0 9 2 10 1 0 9 1 9 2 9 7 9 2
10 15 13 9 1 15 9 7 15 9 2
21 3 9 2 9 7 9 4 13 15 1 3 15 4 13 11 7 13 9 1 9 2
31 15 4 13 0 2 7 15 4 13 9 1 9 1 0 9 7 1 9 1 9 2 3 16 15 3 4 13 1 0 9 2
40 11 4 10 10 12 9 13 1 10 11 1 0 9 7 0 9 2 10 11 15 13 0 0 2 0 0 0 2 0 14 13 1 1 10 11 15 13 9 1 2
17 3 0 9 2 3 0 9 2 4 11 13 15 1 1 10 9 2
25 15 13 1 1 10 0 9 1 10 9 1 11 1 14 13 10 9 2 1 14 13 9 1 9 2
2 9 2
15 9 4 13 16 11 9 13 1 1 9 1 10 0 9 2
5 2 15 4 13 2
11 1 14 13 9 1 9 4 15 13 9 2
30 2 9 4 13 1 3 10 10 15 15 13 14 13 9 2 13 11 11 2 9 1 9 1 9 7 9 1 11 11 2
11 10 9 13 1 15 9 7 10 0 9 2
13 13 15 15 2 4 15 13 9 16 15 13 9 2
16 11 11 4 1 0 9 13 1 9 2 9 7 9 1 9 2
9 9 13 10 9 1 10 0 9 2
7 9 1 10 9 13 0 2
34 11 1 9 1 0 0 9 1 11 2 11 2 4 13 1 12 9 1 14 13 9 2 15 3 4 13 9 1 9 1 9 7 9 2
14 11 11 11 11 11 13 3 10 0 0 9 1 11 2
20 2 16 9 2 9 7 10 9 13 9 2 4 15 13 0 9 1 0 9 2
21 1 9 4 15 13 0 9 1 1 10 9 2 13 11 11 2 9 1 0 9 2
28 16 9 13 0 1 9 2 4 15 13 9 2 13 9 7 9 3 1 10 0 9 15 3 13 9 1 9 2
27 0 9 13 15 12 9 16 11 11 7 10 0 2 11 2 9 13 10 0 9 7 13 9 1 0 9 2
18 11 13 9 1 0 9 2 1 9 1 11 11 11 7 11 10 11 2
18 15 13 16 9 13 1 0 9 2 1 14 13 10 9 1 9 11 2
