4303 11
4 0 9 1 9
11 1 9 13 0 9 2 9 2 1 9 2
16 15 13 3 16 3 12 9 4 14 13 1 9 1 0 9 2
9 15 13 0 1 10 9 1 9 2
9 15 13 3 1 0 9 7 9 2
11 10 9 15 1 10 9 13 3 13 9 2
65 10 9 4 2 9 1 9 2 9 2 9 2 9 2 9 7 0 9 2 2 9 2 0 9 7 3 0 0 9 2 2 2 9 1 9 2 16 10 0 13 1 9 1 3 3 0 9 2 2 9 1 9 2 16 10 0 13 1 9 1 3 3 0 9 2
11 9 0 9 4 9 7 4 7 3 13 2
14 0 9 4 3 9 1 9 2 0 9 2 0 9 2
20 9 15 1 9 3 13 1 3 12 9 4 3 13 7 9 7 3 13 3 2
12 0 9 13 0 9 1 9 1 12 9 9 2
12 13 16 9 3 4 13 3 10 12 9 12 2
2 9 13
22 1 0 9 2 9 7 9 13 9 14 13 9 1 9 3 10 9 15 4 13 12 2
17 1 9 12 2 15 3 13 12 9 9 2 4 9 13 7 3 2
2 9 13
15 9 4 13 1 9 2 16 15 13 0 9 3 12 9 2
10 0 9 13 1 9 13 1 0 9 2
11 9 9 13 1 9 10 12 9 1 9 2
20 3 15 13 9 12 2 9 12 2 4 9 3 4 0 1 10 12 9 12 2
26 1 9 13 15 15 1 14 4 0 13 3 16 15 3 4 0 1 15 7 13 7 4 13 9 3 2
8 0 9 1 9 1 3 0 9
20 9 1 0 9 1 3 0 9 13 1 12 9 1 12 9 1 9 7 9 2
7 3 13 9 1 12 9 2
16 3 15 13 12 9 9 4 9 4 0 1 10 12 9 12 2
6 9 1 9 4 13 2
15 9 4 3 3 13 1 9 1 9 2 9 7 0 9 2
12 15 13 1 16 9 7 0 0 9 13 9 2
20 7 9 4 13 9 7 9 1 9 1 9 1 0 9 7 9 1 0 9 2
5 9 13 1 9 2
28 10 0 9 2 15 13 0 9 2 13 1 12 9 1 10 0 1 10 1 0 9 0 9 1 3 12 9 2
17 1 0 0 9 13 9 1 10 9 1 10 9 15 13 12 9 2
11 9 13 3 1 10 0 9 1 12 9 2
2 9 2
8 3 0 9 13 1 12 9 2
15 9 13 12 9 2 2 12 0 1 12 1 12 9 2 2
22 9 13 1 10 9 1 0 7 0 9 7 13 1 9 1 10 1 0 9 0 9 2
13 0 9 4 13 3 1 9 1 0 9 7 9 2
16 1 0 9 0 9 7 9 3 4 3 13 1 10 0 9 2
16 1 0 9 13 3 10 0 9 9 1 9 2 13 3 2 2
30 0 9 13 1 2 0 15 4 0 3 1 9 1 10 0 9 1 9 2 0 15 13 9 15 13 1 9 1 9 2
25 9 1 10 9 0 9 3 4 13 1 0 9 1 14 13 9 13 1 10 0 9 1 12 9 2
3 9 1 9
20 1 10 0 9 13 10 0 9 16 0 15 3 13 9 2 3 13 10 9 2
16 10 9 4 16 10 0 9 13 0 3 3 0 9 9 13 2
22 3 4 10 0 9 14 4 13 10 9 1 12 9 1 9 1 9 7 3 13 0 2
15 0 9 13 0 16 9 13 1 3 12 9 1 9 3 2
10 3 13 15 1 10 0 9 1 9 2
23 1 14 13 9 1 9 1 10 0 9 14 13 0 9 13 9 1 9 1 9 0 9 2
4 1 0 1 9
16 10 3 9 4 13 15 10 9 1 15 15 13 1 10 9 2
8 13 15 7 13 15 1 9 2
1 9
7 10 0 7 0 9 13 2
18 9 1 10 9 4 14 13 15 1 10 0 9 7 13 15 1 9 2
14 1 9 13 15 0 9 2 15 13 1 10 0 9 2
16 9 4 3 13 15 10 9 9 7 15 13 3 3 1 9 2
1 9
18 10 0 0 9 15 15 13 13 1 0 9 1 10 9 2 1 9 2
30 15 4 3 3 3 13 15 0 9 2 15 4 3 13 15 13 3 1 10 9 7 3 3 13 1 15 1 10 9 2
1 9
6 9 4 0 7 0 2
8 10 0 9 13 9 7 9 2
10 10 0 9 13 3 3 1 10 0 2
29 10 0 7 0 9 15 10 0 9 13 2 13 3 10 9 1 10 0 2 3 1 10 9 3 9 13 1 9 2
13 9 1 9 13 15 1 10 0 0 9 1 9 2
18 1 9 4 15 3 13 15 1 10 9 2 15 3 4 0 7 0 2
11 7 13 3 15 4 13 1 10 0 9 2
15 15 4 7 4 13 3 7 13 1 14 13 10 0 9 2
12 1 9 13 15 3 3 1 9 1 0 9 2
11 1 9 13 10 9 1 2 0 9 2 2
26 15 13 1 9 1 10 9 15 9 3 13 2 3 9 1 0 7 0 9 7 1 9 3 1 9 2
19 10 9 9 7 9 7 10 1 9 0 9 4 13 15 7 3 9 9 2
1 9
9 15 4 14 13 3 1 12 9 2
15 15 4 13 10 9 7 3 10 9 1 9 7 0 9 2
7 15 13 3 1 15 0 2
14 13 3 1 0 9 14 13 9 7 13 9 1 15 2
10 0 9 2 9 7 9 13 0 9 2
1 9
6 10 9 4 3 0 2
15 15 0 4 3 0 7 0 7 13 15 0 1 15 0 2
6 13 3 10 0 9 2
14 13 15 16 10 9 1 9 13 2 3 13 1 9 2
10 15 4 3 9 2 15 4 10 9 2
10 9 4 3 1 9 0 7 3 0 2
1 9
11 15 13 3 0 9 9 1 10 9 9 2
20 15 13 10 9 15 4 4 0 7 1 15 0 7 1 9 16 15 13 3 2
14 15 13 3 9 1 10 9 15 4 0 0 12 9 2
17 15 4 14 13 1 9 2 3 9 4 0 2 16 15 13 3 2
17 15 4 3 3 1 9 13 15 0 14 13 9 1 15 15 13 2
1 9
16 15 4 1 10 9 14 4 13 7 13 15 15 4 13 0 2
13 13 3 3 1 9 3 14 3 13 9 1 0 2
5 10 9 2 10 9
23 15 13 3 3 10 0 9 9 2 9 2 9 2 9 3 2 15 15 4 14 13 3 2
8 9 1 10 9 4 3 0 2
28 3 4 15 13 0 9 1 10 9 7 13 15 1 9 3 2 16 9 4 0 14 13 7 0 14 13 1 2
20 3 4 9 2 3 1 9 2 13 10 0 9 2 0 1 15 1 10 9 2
14 15 4 3 13 1 14 13 10 0 9 1 0 9 2
3 13 1 15
20 9 2 4 3 13 1 9 2 2 9 7 9 2 3 16 15 13 0 9 2
7 15 13 15 1 9 1 9
1 9
1 9
1 9
1 9
1 9
1 9
1 9
12 13 15 15 1 0 9 3 13 1 3 15 2
1 9
8 9 2 3 9 2 9 2 9
7 9 2 1 0 7 10 9
4 9 4 10 9
12 9 13 15 3 7 3 1 9 9 7 9 2
13 9 13 15 0 1 9 1 9 1 9 7 9 2
3 10 0 9
9 1 9 13 15 3 12 1 9 2
11 10 0 9 1 9 13 1 9 3 12 2
35 3 4 15 4 13 1 9 7 9 2 9 1 9 2 9 7 9 1 9 2 9 2 9 3 2 3 16 15 4 2 0 2 1 9 2
15 1 9 13 15 1 0 9 2 1 9 1 3 3 12 2
8 3 13 15 10 0 9 9 2
12 3 13 9 9 2 15 3 13 1 3 12 2
15 16 15 13 1 10 9 7 13 15 13 15 9 1 9 2
15 13 15 3 13 1 9 1 9 2 4 15 13 15 3 2
18 10 9 13 12 7 3 12 9 2 3 15 4 13 15 13 1 9 2
1 9
8 10 0 13 3 3 0 9 2
23 16 0 9 1 10 0 9 13 0 9 2 15 13 3 0 9 14 13 2 4 9 13 2
18 1 10 9 13 9 3 1 14 13 3 7 10 0 9 1 10 9 2
11 12 9 1 9 1 9 4 0 7 9 2
24 1 16 15 4 13 10 9 7 4 13 10 9 15 13 1 10 9 4 15 13 3 0 9 2
20 15 15 13 3 1 9 4 14 13 10 0 9 7 10 0 9 1 10 0 2
13 15 13 15 13 9 1 10 9 1 3 12 9 2
6 10 9 13 12 9 2
18 16 15 13 15 3 4 15 3 13 15 1 9 2 15 3 4 0 2
10 15 15 13 3 1 9 13 1 9 2
6 10 9 13 12 9 2
8 3 1 0 4 9 3 0 2
14 0 9 11 13 9 15 15 13 3 0 9 14 13 2
14 10 9 1 10 0 4 3 13 3 0 7 0 9 2
12 15 13 3 3 0 9 7 0 0 1 9 2
13 10 0 0 13 9 11 2 15 13 12 9 9 2
9 0 4 3 13 15 13 1 9 2
13 0 15 13 9 11 13 10 0 9 2 12 9 2
9 15 13 3 1 0 9 7 9 2
38 16 15 13 3 1 0 9 7 0 15 13 15 1 16 15 1 9 13 16 3 15 13 9 14 13 10 9 7 13 10 9 15 13 1 9 7 0 2
11 13 16 15 4 13 15 15 13 1 15 2
16 10 0 9 4 15 13 0 9 1 3 15 3 13 0 9 2
36 0 2 15 1 9 3 4 13 1 9 7 15 13 9 1 9 7 9 2 4 13 15 1 0 9 1 9 1 14 4 13 3 1 0 9 2
18 0 15 13 0 9 7 12 9 13 0 9 2 15 13 1 9 9 2
12 1 15 4 15 13 1 9 2 10 9 2 2
9 1 9 13 0 9 1 10 0 9
14 0 9 1 9 1 9 1 9 1 9 7 1 9 2
5 0 9 1 9 2
7 0 9 1 3 0 9 2
9 0 9 1 9 1 9 1 9 2
12 15 4 0 1 15 14 13 1 10 3 9 2
12 3 13 15 3 3 1 15 1 10 3 9 2
8 0 9 1 9 1 9 1 9
17 1 12 9 12 13 10 0 7 0 9 1 9 1 9 1 9 2
29 15 13 3 15 13 0 7 13 9 1 10 0 0 9 2 9 2 9 2 9 7 9 1 0 9 1 9 2 2
2 0 9
32 10 0 9 13 16 15 13 12 9 3 15 13 9 1 9 12 9 3 9 13 3 1 15 12 9 3 15 13 9 1 9 2
16 1 10 9 13 9 12 9 3 1 9 2 1 9 9 2 2
9 1 9 13 9 12 9 1 9 2
10 15 4 3 3 13 3 1 10 9 2
11 3 3 13 1 9 1 14 13 3 9 2
21 10 0 9 13 16 15 3 1 9 13 15 15 13 14 13 9 16 15 13 0 2
6 1 9 13 9 7 9
12 1 10 9 15 13 13 3 0 9 7 9 2
10 3 13 9 2 9 7 9 1 9 2
19 16 15 4 13 1 10 0 9 9 7 9 13 15 3 15 1 0 9 2
30 10 0 9 2 16 15 13 9 1 10 9 1 10 9 1 10 9 4 15 3 13 15 3 1 10 0 9 1 9 2
8 9 1 9 13 7 0 9 2
4 9 13 7 3
23 16 15 13 9 1 9 1 7 1 9 7 9 13 15 9 1 9 1 10 9 7 3 2
21 15 4 13 9 1 10 9 1 7 1 9 1 9 1 10 9 15 13 1 9 2
18 13 3 9 7 13 15 1 9 3 13 15 10 9 15 13 9 1 2
9 16 15 13 0 9 13 10 0 9
9 10 0 9 13 10 0 0 9 2
15 16 15 13 0 9 13 15 7 3 0 10 9 15 13 2
11 3 13 15 7 3 10 0 9 1 9 2
4 0 9 1 9
10 9 13 3 9 1 0 9 1 12 9
15 3 4 9 13 9 1 3 12 9 0 9 1 0 9 2
11 1 9 13 10 0 9 1 3 12 9 2
13 3 13 9 9 1 12 9 1 9 1 0 9 2
16 16 3 9 13 3 9 1 9 1 9 9 7 13 1 9 2
7 0 9 13 3 9 1 9
29 9 15 4 0 2 1 9 1 9 2 13 1 9 9 1 7 9 1 3 12 9 7 0 9 1 3 12 9 2
15 10 0 9 13 3 1 9 15 13 1 9 0 9 12 2
18 2 16 15 7 9 13 9 1 3 12 9 1 10 12 9 12 2 2
6 13 9 1 3 0 9
20 1 0 9 13 16 15 13 1 9 3 0 9 1 9 7 0 9 1 9 2
9 9 1 9 13 7 2 9 2 2
17 9 1 9 1 9 7 9 13 1 9 3 15 4 9 1 9 2
14 9 1 9 1 9 7 1 9 13 7 3 1 9 2
18 16 15 4 13 9 1 9 1 9 13 3 10 9 7 1 0 9 2
8 0 9 1 9 1 9 1 9
22 16 15 4 13 9 2 3 9 2 3 3 4 9 1 0 9 13 10 9 1 9 2
16 1 10 0 9 4 15 13 9 1 0 9 7 1 0 9 2
6 9 13 12 9 1 9
11 9 1 9 13 1 12 9 9 1 9 2
22 15 13 1 16 9 13 7 16 10 9 15 9 13 1 9 13 1 12 9 1 9 2
8 9 13 1 0 9 7 9 2
8 10 0 0 9 13 3 3 2
7 9 4 3 13 15 0 9
13 10 0 9 13 16 9 3 4 13 15 0 9 2
8 3 13 3 16 15 4 0 2
3 13 3 2
8 7 13 3 1 15 1 9 2
8 3 0 9 13 15 1 11 2
21 15 13 15 1 0 12 7 13 3 3 7 9 7 15 15 13 0 9 1 9 2
11 1 9 1 11 13 3 12 9 1 9 2
13 15 13 12 0 0 9 1 11 10 12 9 12 2
6 15 4 10 0 9 2
8 9 0 0 1 10 0 9 2
35 9 2 12 2 2 9 2 12 2 2 9 2 12 2 2 9 2 12 2 2 9 2 12 2 2 9 2 12 2 7 9 2 12 2 2
14 9 1 10 0 9 13 3 12 1 10 9 1 11 2
6 3 1 11 13 9 2
10 15 4 0 1 0 7 0 11 9 2
12 10 0 9 4 9 1 11 2 11 7 9 2
6 1 10 9 4 9 2
8 10 0 9 4 1 0 9 2
32 9 12 13 12 9 1 9 7 12 9 1 9 9 12 9 2 16 3 12 9 1 9 1 12 9 1 9 4 3 12 9 2
13 4 15 7 3 13 15 3 1 11 7 13 13 2
8 10 0 9 13 10 0 9 2
26 9 1 11 2 11 2 11 2 11 7 11 4 3 1 9 13 9 7 13 15 3 7 3 1 11 2
12 9 1 0 9 4 13 9 1 9 1 11 2
19 9 13 1 9 9 2 11 2 1 9 1 9 2 15 13 9 1 9 2
12 10 0 9 4 1 9 13 15 16 9 13 2
17 9 2 15 4 13 9 2 4 3 13 1 16 10 0 9 13 2
7 10 9 13 9 1 9 2
13 9 4 1 10 9 7 9 0 1 10 0 9 2
6 10 0 13 1 9 2
24 9 3 13 12 9 1 12 9 7 9 7 1 9 1 9 7 9 9 4 3 12 9 9 2
22 9 13 7 9 16 9 7 10 9 4 13 10 1 10 9 0 9 1 10 0 9 2
8 10 9 13 0 9 1 11 2
15 0 9 4 13 3 1 0 9 2 15 4 10 0 9 2
21 15 13 10 9 1 10 9 7 9 2 10 9 1 9 2 9 7 9 7 9 2
11 10 0 9 4 1 0 9 0 1 9 2
6 9 13 9 7 9 2
16 0 9 13 10 9 1 0 9 7 15 13 3 9 1 11 2
9 11 13 1 3 12 9 1 9 2
44 10 9 15 13 10 9 2 3 15 1 9 1 10 9 2 9 1 0 9 7 0 9 7 3 1 9 1 0 9 13 14 13 10 9 7 13 1 9 4 13 9 1 9 2
23 1 9 13 10 9 9 14 13 10 9 9 1 9 9 1 16 9 13 7 10 0 9 2
8 15 13 1 14 13 0 9 2
9 9 4 4 13 15 7 10 9 2
9 15 4 13 9 1 16 15 13 9
18 1 14 13 9 4 0 9 4 13 1 11 12 9 7 9 12 9 2
17 9 4 3 13 0 9 1 9 1 9 1 12 9 9 1 11 2
12 3 12 9 4 13 0 9 1 9 1 9 2
11 10 0 9 13 15 3 15 13 1 9 2
30 9 15 13 10 9 10 12 9 12 13 9 7 9 2 9 7 9 2 9 2 9 2 9 3 2 2 9 7 9 2
5 1 9 13 9 2
7 15 13 3 9 1 9 2
15 11 13 9 1 9 9 7 1 9 9 1 9 1 9 2
13 10 0 9 1 9 9 2 9 2 13 9 12 2
14 15 4 13 9 9 7 9 7 13 9 1 0 9 2
18 1 10 0 9 13 10 0 9 2 15 4 13 1 9 1 9 9 2
34 9 13 1 10 0 9 2 1 9 12 9 2 1 0 7 0 9 7 10 3 0 9 2 1 9 12 9 2 1 0 9 7 9 2
8 0 9 4 13 1 0 9 2
12 9 13 1 16 9 4 4 13 3 7 3 2
16 9 1 9 1 9 2 9 7 9 13 9 1 14 4 13 2
16 7 3 3 9 13 3 2 13 15 16 9 4 0 1 9 2
5 3 13 15 9 2
3 9 12 2
20 3 4 9 10 9 0 1 9 2 7 3 13 15 9 1 10 0 9 9 2
16 1 10 9 9 2 15 13 0 9 2 13 0 0 9 0 2
20 3 13 3 2 16 15 13 15 1 9 1 9 3 2 10 0 1 10 9 2
28 3 15 13 10 9 1 9 7 9 13 15 9 1 10 1 9 9 2 3 9 13 10 9 1 9 7 9 2
14 1 9 15 13 9 0 4 9 15 7 1 0 9 2
22 1 10 9 9 13 9 1 9 12 3 1 10 9 1 10 9 1 9 12 1 9 2
35 16 10 9 3 13 14 13 1 9 12 2 4 15 13 1 16 15 13 1 9 12 2 9 1 0 7 0 9 2 15 13 1 9 12 2
12 3 13 1 3 9 9 1 9 7 0 9 2
3 9 12 2
34 1 10 9 0 9 7 3 1 0 9 15 13 1 10 12 0 9 9 13 10 9 3 3 10 0 7 10 0 9 7 10 0 9 2
17 1 10 9 4 9 3 3 13 1 14 3 13 9 1 0 9 2
109 10 9 2 3 3 9 13 1 10 0 9 2 4 0 2 11 2 11 2 11 2 11 2 11 2 11 2 1 11 2 11 11 7 0 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 1 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 7 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 7 11 2
22 1 10 9 1 9 12 13 9 1 9 1 9 7 9 7 1 0 9 2 9 3 2
24 3 3 10 9 1 10 9 13 10 9 2 13 9 1 10 3 9 2 9 0 1 11 2 2
16 0 9 12 2 12 2 12 2 12 12 12 2 2 12 2 12
16 15 13 16 0 9 3 12 7 0 9 3 12 13 9 12 2
18 10 0 9 3 12 7 3 7 10 0 3 12 7 3 13 9 12 2
18 1 10 9 9 4 0 9 7 9 1 3 0 0 9 13 0 9 2
15 10 9 7 10 9 4 15 13 3 1 9 1 3 9 2
15 1 9 1 9 12 13 3 9 4 13 1 10 0 9 2
15 3 13 15 16 15 3 4 13 10 9 15 13 1 9 2
10 15 4 3 13 15 1 10 0 9 2
21 7 3 4 15 13 9 1 10 9 7 10 9 1 10 9 3 15 3 13 9 2
25 3 13 15 1 10 9 1 9 12 10 0 9 2 2 9 2 2 15 15 4 13 1 0 9 2
12 9 1 10 9 13 1 9 3 1 3 9 2
32 9 1 9 12 1 10 9 2 9 2 2 15 13 1 11 9 3 11 9 2 4 0 1 12 0 9 2 12 1 10 9 2
14 10 9 13 1 10 9 1 10 9 15 13 0 9 2
15 15 4 0 1 10 1 0 11 9 3 11 9 0 9 2
14 3 13 9 1 9 1 9 7 9 1 10 0 9 2
23 1 9 13 10 9 1 9 3 10 9 2 9 3 4 0 1 10 1 0 9 0 9 2
17 1 10 9 4 15 13 3 3 10 0 9 7 3 9 1 9 2
39 15 4 3 3 13 16 15 13 10 9 7 10 9 9 1 11 3 11 2 7 4 0 16 10 0 9 4 3 11 2 11 7 11 2 11 7 0 11 2
36 9 1 9 1 11 2 11 7 11 2 11 11 2 11 11 2 11 11 3 2 4 3 13 2 3 15 13 3 9 1 11 2 11 3 11 2
3 9 1 9
26 3 15 13 1 10 0 9 15 3 13 9 2 4 15 13 9 1 10 9 15 4 0 1 10 9 2
17 10 9 13 0 9 7 15 1 9 1 9 2 3 11 7 11 2
27 7 10 0 1 10 0 9 2 15 3 4 13 1 9 2 4 1 15 13 9 0 1 9 1 9 9 2
20 3 15 13 1 10 0 9 2 4 15 1 9 3 13 3 9 9 1 9 2
10 1 9 7 0 9 13 15 10 9 2
19 3 15 1 9 13 1 11 4 15 13 2 9 2 2 1 10 0 9 2
22 1 10 9 4 15 13 2 16 10 9 13 10 0 9 1 10 9 1 10 0 9 2
34 10 9 15 4 13 1 9 1 9 1 9 4 0 2 11 11 11 11 11 11 11 11 11 11 11 11 11 11 11 11 11 11 11 11
26 16 9 1 7 11 7 11 13 9 11 2 13 15 3 14 13 3 10 9 1 9 1 9 1 11 2
21 3 15 13 3 4 15 3 2 1 14 13 9 2 13 2 11 2 2 1 9 2
3 9 7 9
25 9 15 13 9 4 1 9 1 9 3 13 10 9 1 10 9 15 13 1 16 15 4 13 9 2
22 9 1 3 9 4 4 0 1 9 13 1 9 2 9 2 2 15 4 13 1 9 2
6 9 1 9 1 9 3
39 9 13 3 10 9 1 0 9 1 9 2 3 15 4 13 9 1 1 10 9 10 0 9 13 15 7 3 13 9 1 1 10 9 7 10 9 9 13 2
14 9 15 13 9 1 10 9 4 13 15 1 10 9 2
19 10 9 1 11 2 3 3 12 13 1 9 1 9 2 13 1 11 9 2
11 3 9 7 9 13 3 7 13 3 9 2
10 15 13 0 9 14 13 9 1 9 2
25 3 10 12 9 12 4 15 13 1 0 2 12 0 9 12 0 9 2 9 12 9 12 9 2 9
17 9 1 0 9 13 1 9 15 4 0 1 10 0 7 0 9 2
9 15 13 3 3 3 3 7 9 2
11 9 9 4 15 3 13 16 15 13 9 2
6 9 4 0 1 9 2
34 1 9 7 9 4 9 1 10 9 13 10 9 0 1 9 9 2 9 3 1 9 2 3 12 1 9 2 3 9 7 9 13 0 2
19 0 9 2 3 9 3 4 3 0 7 9 3 13 9 1 10 9 9 2
1 9
9 10 0 9 13 1 9 7 9 2
1 9
18 9 1 0 9 13 1 10 9 15 4 0 1 10 0 7 0 9 2
23 9 2 15 13 16 9 13 14 13 1 9 9 2 13 3 1 9 1 0 9 1 9 2
34 1 0 0 9 13 9 3 0 9 2 0 9 13 3 1 9 2 16 9 4 13 3 3 1 0 7 1 9 1 0 9 1 9 2
18 0 9 2 9 2 3 15 4 13 9 1 9 14 13 9 1 9 2
1 9
17 9 7 9 4 4 0 1 2 9 2 3 15 13 3 1 9 2
1 9
19 7 9 7 9 13 3 1 9 9 2 9 3 3 1 0 9 1 9 2
36 1 0 0 9 13 9 3 0 9 2 0 9 13 3 1 9 2 16 9 4 13 3 1 9 3 1 0 7 1 9 1 0 9 1 9 2
8 9 13 3 1 9 7 9 2
11 9 4 13 1 9 0 1 3 12 9 2
14 0 9 4 13 9 16 10 0 9 13 10 3 9 2
19 9 1 10 9 15 13 9 13 15 3 1 2 9 1 9 1 11 2 2
20 15 13 12 9 7 4 13 1 9 7 9 1 9 9 12 2 9 2 9 2
17 9 2 3 15 4 0 16 9 13 3 1 9 3 3 7 0 2
1 9
13 9 7 9 4 4 0 1 2 9 2 1 9 2
1 9
10 10 9 13 1 9 1 0 0 9 2
11 9 13 3 1 9 1 0 9 1 9 2
27 1 0 9 1 0 9 13 3 3 9 1 1 16 9 7 9 4 13 13 3 9 1 9 16 9 13 2
24 1 0 9 13 9 1 9 13 1 9 1 9 1 9 1 14 13 16 10 9 13 14 13 2
28 9 2 9 2 3 15 13 16 9 7 13 9 3 3 7 0 2 7 13 3 1 9 1 0 9 3 0 2
1 9
17 9 7 9 4 4 0 1 2 9 2 7 2 11 2 1 9 2
1 9
19 10 9 7 3 2 3 9 13 1 9 3 1 9 1 0 9 1 9 2
25 3 0 1 15 16 10 9 1 9 4 13 3 1 9 2 13 15 3 1 9 9 2 9 3 2
14 1 9 7 9 13 0 9 15 9 4 13 9 1 2
11 9 4 13 1 9 0 1 3 12 9 2
14 0 9 4 13 9 16 10 0 9 13 10 3 9 2
19 9 1 10 9 15 13 9 13 15 3 1 2 9 1 9 1 11 2 2
20 15 13 12 9 7 4 13 1 9 7 9 1 9 9 12 2 9 2 9 2
2 9 13
12 10 0 9 1 10 9 4 7 9 0 9 2
20 15 4 3 13 1 0 9 2 3 15 3 4 10 0 9 1 16 9 13 2
12 0 9 1 9 13 7 4 1 9 4 0 2
4 3 13 9 2
12 10 9 1 0 9 4 9 13 1 10 9 2
12 13 9 0 4 9 13 1 9 1 10 9 2
5 9 13 0 9 2
13 9 4 13 1 9 1 9 2 15 13 1 9 2
3 3 9 2
15 1 9 13 9 10 0 9 2 15 3 13 9 1 9 2
10 10 9 13 1 0 9 3 1 9 2
11 1 14 13 10 9 1 9 4 9 13 2
13 1 9 13 10 0 3 0 9 0 1 0 9 2
18 9 13 9 14 1 10 9 7 1 0 9 13 16 9 13 7 3 2
3 3 3 2
24 10 3 0 9 13 1 0 9 1 9 3 3 12 9 1 10 9 10 0 9 4 4 13 2
10 1 10 9 4 9 1 10 9 0 2
17 4 9 4 0 2 4 15 13 12 9 1 9 2 16 9 13 2
3 3 0 2
17 16 9 13 1 0 9 13 15 16 9 9 4 0 7 12 9 2
29 3 7 12 9 1 9 13 0 2 0 3 1 16 15 1 0 9 3 13 0 9 1 10 3 0 9 1 9 2
13 15 4 10 9 13 16 9 9 4 0 14 13 2
12 9 4 3 13 13 10 0 9 1 10 9 2
14 10 0 9 13 0 2 0 16 0 9 13 1 9 2
4 3 13 15 2
80 1 14 9 9 4 13 0 13 16 15 2 12 0 12 9 1 10 0 9 0 0 9 7 0 12 9 1 0 9 13 2 12 10 9 1 10 9 2 3 12 9 2 2 12 9 2 2 1 10 3 0 9 2 9 7 9 2 2 15 13 1 10 9 7 15 2 12 13 7 13 1 9 3 1 10 1 15 0 9 2
9 9 7 9 13 0 3 9 13 2
11 15 4 3 13 1 9 7 13 1 9 2
6 3 7 3 13 9 2
38 9 4 13 9 2 9 1 3 12 2 12 1 9 1 11 2 11 12 2 12 9 7 1 3 12 2 12 1 9 1 11 2 0 9 2 9 11 2
16 16 9 13 1 9 1 3 12 4 15 13 9 3 10 9 2
11 10 9 13 12 9 7 13 3 9 13 2
1 9
68 9 1 9 4 15 13 9 2 9 1 9 12 1 3 12 2 12 2 9 2 9 2 9 3 12 2 12 2 3 9 12 1 3 12 2 12 2 12 10 9 3 9 13 1 15 1 9 1 3 12 12 10 9 3 9 1 11 3 11 13 9 1 9 7 1 0 9 2
45 15 4 3 7 1 9 13 9 9 1 11 2 11 12 2 12 9 7 11 12 2 12 9 1 3 12 2 12 2 3 1 11 2 0 9 2 9 11 2 1 3 12 2 12 2
14 15 4 3 13 15 0 1 9 1 10 0 0 9 2
17 15 15 13 9 13 3 3 9 1 9 1 16 0 9 4 13 2
12 15 13 0 1 9 3 15 13 9 1 9 2
5 3 15 13 9 2
33 13 9 16 15 2 3 4 0 2 7 9 4 13 1 9 1 0 9 2 4 15 2 16 15 13 15 0 2 4 13 0 9 2
9 13 3 3 10 9 4 9 13 2
22 13 9 16 15 4 2 0 2 4 9 13 2 3 9 13 0 9 1 10 0 9 2
15 15 4 13 1 9 2 1 0 9 7 0 9 1 9 2
4 13 9 9 2
16 13 9 0 0 7 0 9 2 13 11 9 1 9 1 9 2
4 15 15 13 9
40 4 15 13 14 13 12 7 0 9 7 3 13 1 15 7 13 16 15 4 0 2 13 1 16 9 13 0 3 12 9 1 10 9 3 9 4 4 13 9 2
9 15 13 9 14 13 10 0 9 3
8 1 9 0 9 1 9 12 2
10 7 15 13 3 3 12 9 14 13 2
6 9 13 3 12 9 2
15 12 1 9 3 15 4 13 10 0 9 1 12 9 9 2
14 12 1 9 2 9 12 3 9 13 1 9 12 9 2
20 1 0 9 3 9 1 0 9 2 1 12 2 12 2 12 2 12 9 3 2
6 7 10 9 4 0 2
24 1 14 3 13 10 9 2 3 7 3 2 3 12 9 2 2 4 15 13 1 1 0 9 2
17 7 1 9 1 10 0 9 13 15 3 1 10 0 2 9 2 2
8 13 3 1 15 1 0 9 2
10 3 13 15 0 9 3 10 0 9 2
15 10 9 1 9 4 3 10 9 15 13 1 15 1 9 2
23 15 13 3 3 9 14 13 0 9 7 13 3 0 9 3 10 0 0 9 1 12 9 2
28 16 15 3 13 3 0 10 9 2 7 10 9 1 15 2 1 10 9 7 13 9 13 3 1 12 9 9 2
6 16 15 13 3 10 9
7 13 1 10 10 3 9 2
6 3 4 15 3 3 2
29 15 13 3 10 9 3 15 13 14 13 1 12 0 9 7 3 13 3 9 1 0 9 3 10 0 2 0 9 2
11 1 0 9 13 15 1 3 15 13 1 2
5 15 4 3 0 2
5 15 4 13 1 2
13 9 13 3 9 2 3 9 3 2 15 13 9 2
8 10 9 13 3 1 0 9 2
4 13 3 3 2
17 15 13 3 0 10 9 2 7 10 9 1 15 2 1 10 9 2
15 10 9 4 15 13 1 9 7 1 9 2 9 7 9 2
21 7 13 3 3 16 15 4 13 9 3 3 15 13 3 9 1 15 1 10 9 2
9 0 9 4 9 10 12 9 12 2
40 16 15 13 3 7 12 9 7 16 15 3 13 0 9 9 3 1 9 4 15 2 16 15 13 2 13 1 10 9 15 13 16 15 13 3 1 0 9 9 2
2 9 2
19 1 14 13 1 9 4 15 13 3 12 9 0 1 10 9 1 3 9 2
8 10 9 13 12 9 1 9 2
9 7 15 4 13 3 7 12 9 2
5 0 9 3 9 2
9 1 10 9 13 15 10 0 9 2
20 15 13 3 10 0 9 1 12 9 1 10 9 15 13 3 10 12 9 12 2
10 9 13 1 10 9 1 3 12 9 2
2 0 9
7 9 1 9 4 3 0 2
14 0 9 2 7 9 3 2 4 13 3 3 7 3 2
29 7 2 16 15 13 9 1 9 1 9 12 7 9 1 9 3 4 14 13 12 9 2 13 15 3 1 0 9 2
7 9 9 1 9 13 3 2
30 3 13 9 1 10 9 15 13 1 9 1 12 9 9 2 9 13 1 9 7 16 15 4 0 1 9 1 12 2 2
15 16 9 13 7 13 13 9 1 9 7 9 1 9 0 2
9 0 9 13 1 0 9 7 9 2
5 13 7 13 1 9
3 9 1 9
3 0 7 9
15 9 4 13 9 3 1 9 12 2 3 1 9 12 2 2
16 1 9 13 9 15 1 9 7 9 1 9 1 9 1 9 2
12 10 9 13 9 1 7 9 7 9 7 9 2
1 9
19 9 13 0 0 9 1 2 3 4 15 0 3 9 12 2 3 0 2 2
15 9 2 9 7 9 13 0 9 1 10 9 9 1 15 2
15 9 13 1 9 12 7 12 2 9 7 9 1 0 9 2
14 9 4 13 9 10 9 2 7 9 7 9 7 9 2
27 9 7 9 4 14 13 0 1 9 12 7 12 2 3 4 9 0 1 9 12 7 4 3 13 3 2 2
23 0 9 2 9 2 2 3 9 1 10 9 2 4 10 9 1 9 12 13 1 12 9 2
7 3 13 9 1 9 12 2
11 10 0 9 13 1 0 9 1 9 12 2
2 0 9
24 1 9 4 10 9 13 12 1 12 9 2 2 9 2 9 7 9 2 2 9 2 9 2 9
10 10 12 0 13 7 0 7 0 9 2
3 9 1 9
27 1 9 2 9 2 9 7 9 2 7 9 13 9 14 13 1 0 2 0 2 7 0 2 0 2 9 2
4 9 1 0 9
8 0 9 13 0 9 1 9 2
3 3 0 9
11 10 3 0 9 1 9 13 3 0 9 2
12 12 9 4 13 1 15 1 10 9 1 9 2
24 9 4 3 13 1 0 9 1 0 9 7 9 2 7 9 4 13 9 1 9 1 0 9 2
18 9 1 10 9 13 1 9 1 9 7 9 10 9 15 4 13 9 2
15 9 4 3 14 13 1 9 1 9 2 1 9 1 9 2
8 9 13 3 1 0 0 9 2
4 0 1 10 9
23 1 9 1 0 9 4 9 13 16 9 4 13 1 9 9 1 9 15 13 9 7 9 2
12 3 12 9 4 13 1 10 9 1 10 9 2
16 1 0 9 4 9 1 0 9 9 13 2 16 9 3 13 2
7 9 13 9 7 13 9 2
41 9 13 10 0 9 1 10 9 9 2 1 9 9 7 9 1 9 9 2 9 2 9 2 9 7 9 1 9 9 2 9 2 9 2 9 2 9 2 9 7 9
23 9 4 13 3 1 10 9 1 15 7 13 1 9 1 9 1 12 7 15 1 10 9 2
15 9 13 3 0 9 15 3 4 13 1 10 9 1 9 2
13 9 13 7 3 1 9 12 1 12 7 0 9 2
19 9 9 4 13 2 7 9 13 3 1 9 1 9 12 2 12 7 12 2
6 3 13 9 10 9 2
16 1 0 4 9 14 1 0 9 13 9 1 9 9 7 9 2
3 9 1 9
15 10 0 9 13 3 16 9 1 10 9 9 13 7 13 2
5 3 13 10 9 2
13 1 9 13 9 1 0 9 7 1 9 7 9 2
6 10 0 9 13 0 2
15 15 13 0 9 1 9 0 9 14 13 15 0 7 0 2
25 9 1 9 9 13 7 13 2 3 16 9 1 0 9 13 1 9 9 7 9 7 13 1 9 2
13 9 4 3 14 1 0 9 4 13 1 0 9 2
9 1 9 9 13 7 9 7 9 2
12 15 4 3 7 3 13 3 1 9 0 9 2
4 9 1 0 9
26 9 4 13 1 3 2 9 2 9 7 9 2 9 2 0 9 7 9 2 9 2 9 2 9 7 9
11 9 1 10 9 13 1 15 1 9 9 2
11 10 9 1 9 1 10 9 13 3 0 2
5 9 1 9 0 9
15 10 0 9 1 9 4 14 13 9 9 7 9 1 9 2
18 9 4 14 13 0 9 1 9 1 10 9 7 3 0 9 1 15 2
17 10 9 13 3 0 0 9 1 0 9 14 0 13 9 7 9 2
16 9 4 3 4 3 13 1 0 9 2 3 16 9 4 15 2
11 9 13 10 0 9 3 1 0 0 9 2
15 9 7 9 4 9 15 4 14 13 1 0 9 7 3 2
17 3 13 9 2 15 9 4 13 7 1 0 9 13 1 0 9 2
14 9 13 1 10 9 2 15 4 13 12 7 0 9 2
24 2 14 13 2 13 7 13 10 9 2 4 9 1 10 9 15 13 9 9 2 9 7 9 2
20 1 10 0 9 4 15 3 13 15 10 9 1 9 7 9 2 9 7 9 2
19 1 14 13 9 3 0 4 15 13 9 1 0 9 7 10 0 12 9 2
11 9 13 1 10 0 9 1 9 1 9 2
9 9 13 1 0 9 0 1 9 2
18 0 9 4 14 13 1 14 13 9 7 3 1 14 13 9 1 9 2
17 1 10 9 1 15 4 15 3 0 14 13 10 9 1 10 9 2
14 10 9 4 13 9 14 13 10 0 0 1 10 9 2
16 9 13 1 15 1 16 9 4 13 3 1 9 1 0 9 2
8 9 13 0 9 14 13 9 2
11 15 4 13 7 1 9 7 1 0 9 2
20 1 0 9 13 9 1 0 9 7 13 0 9 9 1 9 2 3 1 9 2
16 9 4 3 13 1 9 7 13 3 1 9 1 10 0 9 2
24 9 2 9 7 9 13 3 0 9 14 1 0 9 13 9 3 3 3 13 1 10 0 9 2
13 1 10 9 9 13 9 0 9 7 10 0 9 2
11 15 4 3 3 0 3 10 9 4 13 2
9 9 1 9 1 9 4 12 9 2
14 1 9 4 12 7 0 9 13 1 12 7 10 9 2
23 15 4 3 13 9 1 9 1 9 2 9 7 9 7 1 9 1 0 2 3 0 9 2
15 3 13 9 1 9 9 2 9 7 9 1 9 7 9 2
10 15 4 3 13 3 15 4 13 15 2
13 1 0 9 13 10 9 15 13 1 9 7 9 2
10 13 3 9 9 12 7 9 9 12 2
1 9
17 9 9 4 13 1 16 9 7 9 13 10 0 9 7 0 9 2
98 15 13 3 2 14 13 9 2 9 2 9 7 9 1 9 7 9 2 2 14 13 9 7 9 1 9 1 10 9 15 13 15 2 2 14 13 9 1 9 2 13 9 7 9 1 9 2 2 14 13 3 9 7 9 2 2 14 13 3 7 13 16 9 7 9 13 1 9 2 13 1 9 7 13 1 9 2 2 14 1 0 9 13 1 9 7 14 13 10 0 1 9 2 3 1 10 9 2
20 9 9 1 9 1 9 7 1 9 13 16 15 13 12 9 2 13 0 2 2
8 9 9 13 1 9 7 9 2
6 9 9 13 1 9 2
17 1 0 9 13 9 0 9 15 13 1 15 15 13 9 7 9 2
6 15 13 15 1 9 2
1 9
7 10 0 9 13 1 9 2
15 3 13 9 15 3 13 9 0 9 2 9 7 0 9 2
17 9 9 13 9 1 9 1 9 7 9 3 15 13 9 1 9 2
12 9 1 9 13 1 9 9 1 9 1 9 2
10 9 1 10 9 13 1 14 13 3 2
6 13 3 9 9 12 2
6 15 13 15 1 9 2
1 9
9 1 10 0 9 13 9 10 9 2
14 3 13 3 9 1 9 1 9 3 9 3 13 3 2
26 9 4 13 1 16 9 9 13 3 1 3 0 9 2 13 9 1 9 7 13 9 1 9 7 9 2
14 10 0 0 9 4 1 0 9 1 9 13 10 9 2
6 13 3 9 9 12 2
6 15 13 15 1 9 2
1 9
19 10 9 3 12 9 13 12 9 1 9 7 9 2 3 12 9 1 9 2
14 9 13 3 1 9 7 1 15 15 13 9 1 9 2
11 15 4 0 7 13 3 3 3 1 9 2
10 9 13 3 9 1 10 3 9 13 2
7 15 13 10 9 1 9 2
13 1 9 13 9 13 3 16 9 4 13 7 0 2
10 9 13 1 16 9 13 3 1 9 2
19 9 4 13 3 1 16 9 4 13 1 12 9 2 9 1 12 9 12 2
6 15 13 15 1 9 2
1 9
6 15 13 0 9 9 2
9 9 1 9 1 9 3 12 9 2
9 9 1 9 1 9 3 1 9 2
11 9 1 0 9 1 9 3 1 9 9 2
10 9 1 9 15 13 9 1 0 9 2
8 15 13 15 1 9 7 9 2
1 9
22 9 7 0 9 4 13 9 3 1 12 9 9 7 9 1 9 1 12 9 7 0 2
10 10 9 4 0 1 0 7 0 9 2
10 9 7 9 13 3 7 1 0 9 2
11 0 9 13 3 9 2 1 9 1 9 2
8 15 13 15 1 9 7 9 2
1 9
5 13 9 9 12 2
1 9
8 0 9 13 0 9 1 9 2
4 1 15 13 2
5 9 2 15 13 1
14 9 15 1 0 9 13 1 9 16 9 13 7 13 2
13 15 4 0 1 9 1 9 12 9 2 12 9 2
13 9 13 1 9 7 13 3 1 3 0 9 4 2
19 9 15 13 3 9 10 7 10 9 1 9 2 3 1 12 9 1 9 2
6 9 4 1 9 0 2
16 9 15 13 3 0 9 1 10 0 9 1 9 3 9 13 2
9 9 13 3 1 3 0 9 4 2
4 9 13 3 1
15 3 0 9 1 9 15 1 9 13 3 9 16 9 13 2
9 9 13 3 1 3 0 9 4 2
6 15 13 15 1 9 2
16 0 9 10 9 13 4 13 9 1 9 1 9 2 9 2 2
14 15 13 1 3 3 1 0 9 7 9 4 1 9 2
5 9 13 1 9 2
8 15 13 15 1 9 7 9 2
4 0 9 7 9
15 9 7 9 1 3 0 9 13 0 9 7 9 1 9 2
5 15 13 1 9 2
14 9 13 1 9 7 10 0 9 11 2 11 7 11 2
13 15 13 15 1 9 1 0 9 7 9 7 9 2
1 9
11 1 10 0 9 13 0 9 10 0 9 2
13 15 4 13 3 9 2 9 2 9 7 0 9 2
9 9 13 3 1 10 9 7 9 2
12 9 7 9 13 3 9 2 9 7 0 9 2
7 0 9 13 9 1 9 2
25 1 9 3 3 13 0 3 15 4 13 15 1 9 7 1 9 1 9 15 13 1 9 14 13 2
3 9 1 9
11 3 12 9 1 9 3 12 9 13 9 2
17 9 4 0 0 1 3 0 9 15 13 7 1 9 9 7 9 2
7 9 9 13 3 1 9 2
14 9 15 13 3 7 3 12 9 2 9 13 0 9 2
13 16 9 4 0 7 3 12 9 2 9 13 9 2
11 10 0 9 13 1 10 9 7 10 9 2
11 9 1 12 9 7 0 4 13 0 9 2
12 9 4 12 9 1 9 3 15 13 12 9 2
13 15 13 1 12 9 1 9 1 10 9 1 12 2
9 9 13 0 1 9 9 7 9 2
13 15 4 10 9 13 3 16 9 3 4 10 0 2
10 3 10 0 9 15 13 1 10 9 2
15 9 1 9 13 1 9 15 13 0 9 7 3 12 9 2
35 9 13 16 9 13 10 0 9 2 3 12 9 7 9 2 7 0 9 2 9 7 9 1 9 7 1 0 9 9 7 9 1 9 2 2
24 0 9 4 10 9 13 1 10 0 9 16 15 13 10 9 1 1 9 3 12 9 1 9 2
20 1 14 13 10 0 9 13 3 16 9 13 10 9 15 13 1 10 0 9 2
11 9 4 13 9 1 10 9 15 13 3 2
1 9
6 15 4 13 1 9 2
11 9 13 10 9 1 10 9 15 13 9 2
8 15 13 15 1 9 2 9 2
3 9 1 0
19 0 9 13 10 0 9 1 0 15 13 1 9 7 1 0 3 0 9 2
10 15 13 0 9 1 0 2 11 2 2
6 15 13 15 1 9 2
4 9 1 9 2
20 0 9 2 11 2 4 13 1 15 15 13 9 2 9 7 9 2 9 7 9
9 13 9 2 0 9 2 9 12 2
1 9
10 11 0 9 13 3 10 0 0 9 2
16 1 10 9 0 9 13 9 1 9 2 9 7 0 0 9 2
7 9 9 1 9 4 0 2
1 9
16 9 13 9 2 1 9 9 2 1 14 13 7 13 1 9 2
10 3 12 9 1 9 13 1 0 9 2
18 10 0 9 4 1 1 12 7 12 9 1 9 1 10 0 0 9 2
10 1 0 9 4 15 1 9 12 9 2
7 10 0 9 13 1 9 2
5 9 13 1 9 2
10 13 3 9 9 12 7 9 9 12 2
8 15 13 15 1 9 2 9 2
1 9
8 10 0 9 13 1 0 9 2
6 9 9 13 3 0 2
23 9 9 4 9 7 9 13 3 1 1 0 9 2 1 9 1 10 9 3 9 3 13 2
12 1 0 9 4 3 10 0 0 9 13 9 2
16 16 15 4 13 15 4 0 4 9 13 15 1 10 0 9 2
13 15 15 4 0 1 9 9 4 13 15 1 9 2
10 9 9 14 13 3 1 9 4 13 2
20 9 13 3 9 9 14 1 0 9 13 9 3 16 9 4 13 15 10 9 2
9 9 4 13 0 9 14 13 9 2
11 9 4 13 3 12 7 13 1 12 9 2
20 3 4 9 1 3 0 3 13 16 3 9 13 1 9 2 1 9 7 9 2
12 9 15 4 13 1 9 12 13 3 1 9 2
13 9 1 9 1 10 9 13 1 10 0 0 9 2
6 15 13 15 1 9 2
2 0 9
18 16 15 4 13 1 3 0 9 2 0 9 3 13 15 15 1 9 2
9 9 13 15 0 1 15 14 13 2
4 3 3 0 2
16 0 9 13 10 9 10 0 9 1 10 9 7 9 15 13 2
8 9 13 1 9 2 9 2 2
13 1 14 4 13 0 9 4 15 13 9 1 9 2
15 1 9 3 10 9 4 13 13 3 9 1 9 0 9 2
4 3 13 9 2
16 0 15 1 9 7 9 4 3 0 1 16 10 9 4 0 2
12 3 10 9 0 13 10 9 0 3 1 9 2
21 3 9 2 9 2 9 2 9 2 9 7 0 0 9 4 0 1 9 1 9 2
1 9
7 9 4 3 13 3 3 2
25 10 9 13 15 9 1 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 3 2
20 16 15 4 10 0 9 14 13 9 1 10 9 4 15 13 15 1 10 9 2
16 9 4 3 13 1 14 13 9 1 10 9 1 9 7 9 2
16 1 9 1 10 9 13 0 9 3 12 9 1 3 12 9 2
25 1 10 9 9 4 9 13 3 3 3 16 9 4 0 1 0 9 2 3 9 2 9 7 9 2
19 3 13 10 0 9 1 10 9 7 9 13 3 1 10 0 9 2 9 2
18 1 10 3 9 13 9 1 3 0 9 10 0 9 13 1 10 9 2
14 10 0 9 13 3 1 9 7 0 9 1 3 9 2
8 2 13 9 1 9 12 2 2
1 9
11 9 4 13 9 1 0 9 1 0 9 2
18 0 9 2 3 9 2 9 7 9 2 13 3 9 7 3 4 9 2
10 3 0 9 1 10 9 13 1 9 2
22 16 9 4 13 13 9 3 4 9 13 2 1 0 9 4 3 10 9 1 9 13 2
14 1 14 13 0 3 9 4 0 9 13 9 1 9 2
7 3 13 9 10 0 9 2
21 15 13 3 10 0 9 1 9 1 9 2 9 7 9 15 13 9 1 10 9 2
19 9 13 3 9 1 9 1 9 1 9 2 15 13 1 9 7 0 9 2
2 9 0
5 10 9 4 13 2
19 3 13 1 9 1 9 9 7 9 2 0 9 2 9 2 9 7 9 2
26 10 9 4 13 7 1 9 13 15 9 1 9 1 0 9 2 0 9 2 9 9 2 9 7 9 2
7 3 0 9 1 9 13 2
18 10 9 4 13 16 15 13 1 15 9 7 9 1 12 9 1 9 2
14 1 10 9 2 9 2 9 2 13 9 1 0 9 2
11 1 10 9 13 9 9 1 3 9 13 2
19 9 4 0 7 10 9 1 9 15 13 16 15 4 13 9 9 1 9 2
1 9
9 9 4 13 0 9 1 10 9 2
14 7 13 1 9 1 0 9 13 9 1 9 0 9 2
13 9 13 1 15 3 3 0 15 4 13 14 13 2
20 7 10 0 9 1 3 9 13 4 15 13 3 9 1 9 12 1 9 12 2
14 9 4 1 9 12 2 12 7 1 9 12 2 12 2
22 9 13 3 7 12 2 12 2 12 15 13 10 9 1 12 15 13 13 1 12 9 2
24 9 12 13 16 9 1 12 9 1 9 12 13 1 9 1 12 9 7 12 9 12 9 3 2
33 1 15 15 4 13 3 1 9 4 0 9 13 3 10 9 2 15 4 13 1 9 7 13 1 0 9 2 9 2 12 11 12 2
7 9 3 12 9 1 9 2
6 12 9 12 13 9 2
10 10 0 9 1 9 9 13 1 9 2
4 9 13 0 2
6 15 13 3 0 9 2
6 15 4 13 0 9 2
14 15 4 1 9 4 13 1 9 1 10 9 7 9 2
14 1 10 9 1 10 9 13 7 10 0 7 0 9 2
13 12 9 12 13 10 12 7 9 7 10 0 9 2
10 12 7 9 7 0 9 13 3 0 2
10 10 0 9 4 14 13 3 3 3 2
18 10 0 12 7 9 13 3 0 2 7 15 13 3 1 3 0 9 2
4 9 13 3 2
9 15 7 10 0 9 13 7 3 2
4 10 9 1 12
13 3 4 15 4 0 3 15 7 13 9 7 9 2
5 6 2 15 13 2
12 1 10 12 9 12 13 3 10 9 1 9 2
6 15 13 1 9 0 2
15 9 15 13 1 12 7 12 9 4 13 3 1 0 9 2
15 9 15 13 1 12 7 12 9 4 13 3 1 0 9 2
15 13 9 1 12 7 12 9 4 15 13 3 1 0 9 2
16 7 13 15 1 12 7 12 9 4 15 13 3 1 0 9 2
8 10 3 9 13 3 9 13 2
11 7 15 13 3 9 1 9 15 4 13 2
5 3 10 0 9 2
12 9 15 4 13 12 4 13 15 3 1 9 2
10 7 3 4 9 13 1 12 9 9 2
2 9 2
14 16 15 13 12 9 9 1 12 9 9 13 15 12 2
7 3 13 9 3 1 12 2
13 13 15 12 9 13 15 12 15 13 3 1 12 2
4 13 15 0 2
26 16 15 13 10 0 9 9 1 12 2 10 9 1 12 7 10 0 9 9 1 12 13 15 3 12 2
6 3 3 4 15 13 2
11 7 16 9 13 1 12 7 9 13 12 2
8 3 3 4 15 4 13 3 2
10 2 10 0 9 13 15 3 3 2 2
5 15 13 1 9 2
5 7 15 13 0 2
17 16 3 9 13 13 15 15 3 1 12 7 12 9 1 10 9 2
17 7 10 0 4 0 3 16 15 13 3 15 1 9 1 10 9 2
12 9 4 16 15 13 0 9 14 13 9 1 2
12 9 7 9 13 14 13 7 13 10 9 9 2
6 9 1 9 13 0 2
18 15 4 3 13 15 16 12 7 9 1 10 0 3 13 1 0 9 2
6 9 13 3 1 15 2
7 7 9 13 3 1 15 2
6 9 9 7 9 13 2
12 15 4 9 9 16 9 3 4 13 1 9 2
9 3 13 9 3 3 9 4 13 2
16 15 4 3 0 1 9 1 0 9 15 13 3 1 9 9 2
23 1 9 9 2 9 2 9 2 9 4 3 4 13 9 15 3 13 1 12 7 12 9 2
20 3 3 4 15 7 9 1 9 7 9 1 9 13 3 16 12 7 9 13 2
8 9 9 7 9 13 9 3 2
12 15 4 3 14 13 9 1 0 9 1 9 2
10 2 10 0 9 4 12 3 12 2 2
14 3 7 10 0 9 9 13 1 9 1 10 0 9 2
8 13 15 9 1 10 9 3 2
7 9 1 9 4 13 9 2
7 15 13 13 3 1 9 2
8 15 4 10 0 9 1 9 2
9 3 0 4 1 0 9 13 9 2
14 9 4 3 0 7 13 3 3 1 10 0 0 9 2
9 10 0 7 0 9 4 3 13 2
9 12 9 13 12 1 9 1 9 2
6 1 15 4 12 9 2
24 15 4 10 0 9 16 15 15 13 9 3 4 13 9 1 0 9 16 15 13 3 1 9 2
7 1 9 4 9 13 1 2
14 15 13 1 9 3 1 10 9 1 0 9 1 0 2
28 0 9 15 13 15 1 9 7 13 1 9 4 1 0 3 13 9 2 3 16 9 13 1 9 1 10 0 2
8 1 9 4 10 9 4 0 2
6 9 1 9 1 11 9
4 15 4 0 2
17 10 9 1 9 1 13 1 0 9 1 9 7 9 3 1 9 2
5 15 13 0 9 2
8 10 9 1 0 9 13 0 2
4 9 4 13 2
10 9 4 13 10 9 1 16 9 13 2
4 15 13 9 2
3 14 13 1
13 15 15 13 9 4 13 1 16 15 3 13 0 2
19 15 13 3 14 13 3 0 9 1 9 2 1 14 13 7 13 1 2 2
10 3 13 3 10 0 9 1 0 9 2
8 10 0 9 1 9 4 0 2
7 15 13 16 15 13 3 2
14 9 4 10 9 2 3 10 9 1 14 13 1 9 2
29 1 10 9 1 9 15 13 1 9 13 15 15 10 9 1 9 1 11 9 13 1 9 2 9 2 9 7 9 2
2 13 15
7 13 9 9 7 9 9 2
8 13 9 7 9 2 0 2 2
11 15 4 13 15 1 9 1 9 1 9 2
15 13 1 9 3 7 3 7 13 16 15 13 3 15 13 2
9 4 10 9 2 9 7 9 0 2
6 13 9 1 0 9 2
8 15 4 13 16 15 13 3 2
3 13 9 2
4 15 13 9 2
18 9 1 11 9 1 10 0 9 13 1 3 12 9 7 3 12 9 2
25 1 9 1 9 12 4 15 13 10 9 15 13 1 9 7 10 9 15 13 1 11 1 9 12 2
14 15 4 3 13 10 9 1 3 3 9 13 7 13 2
14 10 9 2 11 11 11 2 4 13 1 9 1 9 2
11 3 13 10 9 15 13 1 11 1 11 2
16 15 4 13 1 9 10 9 9 4 0 1 7 16 9 13 2
12 13 10 0 9 1 10 3 0 9 1 9 2
13 1 9 1 9 13 15 10 0 9 15 13 15 2
18 10 0 9 2 11 2 13 3 1 16 9 1 11 9 13 10 9 2
12 15 15 13 4 3 10 9 1 9 7 9 2
15 9 1 9 1 9 12 9 13 1 3 12 7 12 9 2
19 1 9 0 1 9 1 12 7 12 9 4 15 13 10 0 9 1 9 2
1 9
10 9 4 10 9 1 2 0 9 2 2
12 15 13 0 9 15 3 13 1 1 9 9 2
24 9 13 2 0 9 2 7 13 3 7 9 7 7 9 1 0 9 1 14 13 15 0 9 2
17 15 13 3 14 13 10 9 3 0 7 0 7 9 1 0 9 2
16 7 15 4 10 0 9 1 15 15 13 16 9 13 0 0 2
20 0 9 13 3 1 0 7 10 0 9 4 3 3 0 13 3 15 1 9 2
12 9 4 3 10 3 0 9 15 13 0 9 2
9 10 0 9 1 11 4 12 9 2
18 15 4 0 16 10 0 9 2 3 0 2 1 10 9 13 1 9 2
33 16 15 13 16 15 7 15 1 15 13 0 9 1 12 0 9 4 15 12 9 9 16 15 1 10 9 13 0 9 1 10 9 2
12 10 0 9 13 3 1 10 0 2 9 2 2
14 15 13 3 3 16 9 13 3 0 9 1 10 9 2
20 9 13 1 9 9 2 7 15 13 1 9 3 9 9 4 0 7 9 9 2
8 9 4 13 3 7 3 0 2
10 7 9 0 9 13 14 13 9 0 2
8 9 13 3 7 10 0 9 2
11 3 13 15 0 9 1 0 9 1 9 2
9 3 1 3 13 9 9 1 9 2
11 7 3 10 9 15 13 0 13 0 9 2
3 9 1 9
8 9 4 10 0 9 1 9 2
14 9 13 9 14 13 15 15 2 15 13 3 9 1 2
11 10 0 9 4 3 13 0 9 1 15 2
13 10 9 9 4 14 13 15 0 7 15 1 9 2
24 7 9 4 3 4 13 9 1 10 0 9 10 9 13 2 3 15 15 4 3 0 7 15 2
3 11 2 9
8 1 12 9 13 11 10 9 2
11 10 9 9 9 12 2 12 9 0 3 2
3 9 13 2
12 9 13 1 9 7 9 2 1 9 7 9 2
5 15 4 13 9 2
4 15 13 9 2
10 3 9 13 13 9 1 10 0 9 2
5 10 0 9 13 2
5 15 4 13 9 2
4 15 13 9 2
3 15 13 9
7 15 4 3 0 1 9 2
8 1 10 9 2 1 10 9 2
12 9 13 0 9 2 0 9 2 0 9 14 13
9 12 13 9 1 12 9 1 9 2
6 3 4 9 12 9 2
13 7 9 4 3 13 1 10 9 3 9 4 13 2
8 7 9 1 9 9 13 9 2
35 3 13 9 16 15 3 13 10 9 1 10 0 9 7 1 12 9 10 9 1 10 9 2 3 12 9 9 2 3 3 0 7 3 2 2
14 7 3 1 9 4 15 14 13 1 9 2 3 3 2
11 9 4 3 0 1 0 9 7 1 0 2
3 12 9 13
12 10 9 13 12 9 9 3 3 1 10 9 2
10 1 10 9 13 10 9 9 1 9 2
10 9 1 10 9 13 1 7 1 9 2
15 9 1 9 1 7 1 9 13 1 9 7 9 1 9 2
20 10 0 15 13 1 9 4 1 9 13 15 1 9 2 1 9 3 7 3 2
6 10 3 9 4 13 16
7 9 7 9 13 3 15 2
12 9 13 3 16 0 9 3 13 3 1 9 2
5 0 9 13 3 2
14 12 9 7 9 13 0 9 1 9 2 0 9 2 2
6 9 0 4 3 12 2
17 1 15 13 10 0 7 0 15 3 0 13 9 2 9 7 9 2
10 15 4 13 9 1 14 13 1 9 2
23 9 13 15 10 9 1 0 9 1 12 7 12 9 9 1 3 9 2 9 7 0 9 2
3 3 0 9
12 1 9 13 9 2 9 7 9 3 10 9 2
24 9 4 0 1 9 15 13 9 9 1 0 9 2 9 2 9 2 9 2 0 9 2 9 2
13 10 0 9 13 3 0 9 1 9 7 13 9 2
6 10 9 13 10 9 2
8 7 0 9 2 3 0 9 2
14 7 0 9 2 3 0 9 1 9 7 3 0 9 2
24 3 9 13 3 1 10 0 7 0 9 15 13 1 9 9 3 13 9 1 9 7 9 13 2
6 3 4 15 13 15 2
23 10 9 1 9 13 15 3 2 0 9 2 0 9 2 0 9 2 0 9 7 0 9 2
21 10 9 13 15 1 3 15 13 9 2 9 2 10 9 2 9 2 9 2 9 2
14 10 9 13 15 3 15 13 1 7 1 9 2 9 2
4 15 13 9 2
6 15 13 9 2 9 2
12 4 15 10 9 15 9 2 9 4 13 3 2
5 7 9 1 9 2
19 13 15 9 1 9 1 10 9 15 4 13 15 0 2 0 7 3 0 2
8 13 0 9 1 9 7 9 2
23 13 15 9 1 9 1 9 4 15 3 4 0 1 15 14 13 9 1 10 9 7 9 2
8 13 0 9 3 15 13 1 2
12 10 3 9 1 9 4 3 0 14 13 1 2
9 15 4 13 1 9 16 0 13 2
9 15 4 3 13 1 9 7 9 2
36 4 15 13 1 9 1 10 9 7 9 1 9 1 0 9 2 4 15 13 3 1 9 1 9 9 3 16 15 13 10 7 0 9 1 9 2
9 1 9 4 15 3 13 1 9 2
35 9 15 4 13 1 9 1 9 7 4 4 3 0 13 3 3 1 9 7 13 3 1 9 2 13 7 13 9 1 10 0 9 7 9 2
6 9 13 3 1 9 2
13 13 3 1 9 7 9 15 4 13 3 1 9 2
8 13 15 9 1 9 7 9 2
9 9 1 9 4 0 1 0 9 2
16 9 4 3 1 9 1 9 3 13 0 9 1 10 0 9 2
13 1 10 9 4 15 3 13 0 9 1 10 9 2
13 7 9 7 9 4 0 1 0 2 9 7 9 2
12 15 4 3 3 13 1 9 2 9 7 9 2
22 15 4 3 0 14 13 2 15 7 1 9 7 9 2 2 13 7 13 1 0 9 2
14 3 15 13 9 1 9 7 9 2 13 3 9 1 2
13 13 3 3 1 0 9 3 16 15 13 1 9 2
6 13 3 1 1 9 2
16 1 9 4 15 13 9 1 9 15 13 3 1 9 7 9 2
13 13 10 9 3 16 15 3 13 3 1 10 9 2
15 1 9 2 13 9 1 0 9 7 13 3 3 1 9 2
6 15 13 15 1 9 2
10 0 9 13 1 0 9 1 0 9 2
7 9 4 4 0 7 0 2
22 13 15 1 0 9 7 9 4 15 3 13 1 0 9 1 14 13 9 1 0 9 2
19 15 4 3 3 13 1 0 0 9 15 13 9 1 9 7 9 7 9 2
9 0 0 9 1 9 9 4 9 2
25 15 4 0 14 13 1 10 9 1 9 1 9 1 3 15 13 10 0 0 9 1 9 1 15 2
14 10 9 0 9 13 9 2 0 9 7 0 9 2 2
16 10 0 9 13 16 9 4 4 0 1 10 0 7 0 9 2
41 16 15 3 13 1 9 1 9 7 16 15 4 13 1 9 4 15 13 10 9 1 9 1 0 7 3 15 13 1 0 2 9 7 9 15 13 3 7 13 3 2
17 9 4 3 13 1 9 1 12 7 0 9 1 9 1 10 9 2
28 13 0 9 3 1 9 1 0 9 2 0 9 2 4 15 3 13 9 7 13 3 16 10 9 13 10 9 2
10 13 15 0 2 7 9 9 7 9 2
17 9 4 1 0 9 13 3 16 15 4 13 9 7 13 1 0 2
8 3 9 13 0 9 1 9 2
9 13 3 10 9 1 10 0 9 2
6 15 4 13 1 9 2
10 13 15 0 9 4 15 10 0 9 2
15 7 13 15 15 0 2 13 10 9 1 10 9 7 9 2
11 13 10 9 7 13 1 15 1 0 9 2
14 13 3 1 9 1 9 2 3 12 0 9 13 9 2
10 10 9 9 4 13 10 9 7 9 2
20 2 9 3 2 4 9 13 3 3 2 9 13 3 3 12 9 9 1 9 2
18 1 9 7 10 9 9 13 2 13 10 9 2 9 9 9 9 9 9
4 15 4 13 2
24 0 4 0 9 15 2 4 0 12 7 3 2 2 3 4 0 2 7 2 4 0 1 9 2
14 15 1 9 1 9 9 4 16 9 13 1 12 9 2
14 15 15 13 12 9 3 10 12 9 12 13 3 9 2
1 9
16 15 15 4 0 1 9 13 10 9 1 9 1 10 12 9 2
33 16 15 13 15 3 2 7 3 13 15 1 10 12 9 2 4 15 13 15 1 0 9 1 10 9 3 15 4 0 1 9 12 2
23 9 4 13 1 1 9 1 9 7 4 13 1 1 9 1 9 2 1 9 7 1 9 2
20 1 9 13 15 1 10 9 15 4 13 7 1 10 9 15 4 0 1 9 2
14 10 9 4 16 10 0 9 3 12 2 12 4 0 2
11 10 0 9 4 3 0 3 12 2 12 2
4 15 4 13 2
31 15 7 15 15 4 0 1 9 7 0 7 0 3 4 13 12 9 3 10 12 9 2 4 13 1 9 2 9 7 9 2
19 15 4 3 13 10 9 1 9 2 0 1 3 1 9 15 7 15 13 2
10 10 3 9 4 13 1 9 1 9 2
10 1 9 1 9 7 9 13 3 9 2
13 15 15 4 13 4 3 4 0 1 9 3 9 2
4 3 13 9 2
11 13 1 9 9 9 1 10 9 1 9 2
8 3 13 9 3 9 1 9 2
11 1 0 9 13 15 1 9 9 2 9 2
8 1 9 13 15 3 1 9 2
16 3 13 15 9 1 9 7 9 1 10 9 3 15 4 13 2
10 1 15 13 15 0 9 7 0 9 2
10 10 9 4 16 15 13 1 3 9 2
18 9 4 13 2 2 9 2 0 9 2 9 15 13 1 10 9 15 13
27 9 4 13 2 9 1 12 7 0 9 2 9 2 9 1 1 10 9 15 13 2 9 2 9 7 9 2
9 3 3 4 15 13 9 1 9 2
44 9 13 0 2 16 15 13 9 15 13 3 1 0 9 14 13 15 2 13 3 9 2 2 16 15 13 9 7 13 3 7 12 9 2 16 3 7 12 9 13 1 10 9 2
27 16 15 1 9 13 1 12 9 1 10 9 1 12 9 13 3 9 12 9 2 7 9 1 9 13 3 2
6 9 1 9 10 12 9
44 0 9 13 1 3 0 1 7 3 1 10 9 16 15 13 12 9 2 2 1 11 2 11 7 1 11 2 3 9 0 13 9 9 2 13 15 12 9 2 3 9 2 3 2
8 9 7 9 13 0 1 9 2
16 2 3 15 13 9 1 9 2 9 7 9 13 9 12 2 2
1 9
14 1 9 15 13 0 14 13 1 9 13 0 9 9 2
6 10 9 13 0 9 2
7 3 9 13 13 1 9 2
24 16 15 13 3 2 13 1 9 9 9 2 15 4 4 0 1 9 2 7 3 9 4 0 2
18 13 3 1 10 9 2 3 16 15 3 4 10 9 1 14 4 13 2
12 16 15 13 9 1 10 9 2 13 1 15 2
14 16 15 3 13 1 15 9 13 15 1 9 1 9 2
24 15 4 13 12 9 2 10 0 2 9 2 2 10 0 2 9 2 7 10 0 2 9 2 2
14 3 1 9 13 15 12 0 9 2 12 1 10 9 2
5 13 1 10 9 2
8 13 10 0 9 1 10 9 2
5 9 4 13 3 2
16 13 3 3 1 9 7 13 10 9 16 15 13 15 1 15 2
21 3 13 15 1 9 16 15 13 2 13 3 10 9 7 13 15 1 10 0 9 2
6 3 4 15 13 10 2
6 3 13 9 7 9 2
4 11 0 9 13
18 10 9 2 3 10 9 15 13 1 9 7 9 9 2 4 11 0 2
9 9 4 1 12 7 9 1 12 2
7 10 9 4 10 0 9 2
13 1 9 13 16 9 13 9 1 0 7 0 9 2
11 1 9 13 16 9 4 0 1 9 9 2
20 15 13 3 9 2 7 3 9 2 15 13 10 0 9 1 9 9 7 9 2
16 9 1 9 1 0 9 4 13 0 1 9 1 9 1 9 2
17 9 4 3 3 4 0 1 9 2 7 4 1 9 13 1 12 2
10 1 9 1 9 13 9 1 10 9 2
25 1 0 9 7 9 1 10 12 0 9 13 9 1 0 9 15 4 13 1 9 10 12 9 12 2
54 15 13 16 2 9 13 1 10 9 1 12 9 2 2 10 0 9 1 0 9 1 0 9 7 0 9 13 2 9 13 3 1 9 9 2 2 9 13 3 3 1 9 2 2 9 1 9 2 9 7 9 13 3 2
9 9 13 1 9 3 1 0 9 2
15 9 13 9 14 13 1 9 1 9 7 1 10 0 9 2
18 10 0 9 4 13 3 1 9 16 3 12 9 1 9 9 13 15 2
17 1 9 1 9 13 3 12 9 2 3 3 7 9 1 9 9 2
9 9 13 16 10 0 9 4 13 2
16 16 15 13 9 2 13 0 9 2 7 13 9 1 12 9 2
11 9 4 13 7 9 13 3 9 13 15 2
16 9 13 7 13 1 9 1 9 2 3 16 9 3 13 9 2
25 9 1 9 1 9 4 13 2 15 13 16 15 4 4 13 1 10 0 9 16 15 15 13 1 2
9 1 9 7 9 13 3 9 3 2
3 9 13 2
11 15 13 3 9 10 9 15 13 12 9 2
8 9 13 7 13 3 1 9 2
12 15 4 0 16 15 13 12 9 3 1 9 2
5 9 13 10 9 2
14 15 4 3 13 9 9 7 9 9 1 10 0 9 2
15 10 0 9 4 14 13 1 10 9 1 11 9 1 11 2
10 15 4 13 0 9 1 10 0 9 2
7 1 9 13 15 3 3 2
8 15 13 3 1 11 12 9 2
7 7 9 4 13 0 9 2
22 15 13 3 0 0 7 0 15 4 13 15 0 9 2 7 3 15 4 13 0 9 2
24 3 16 15 3 4 13 10 9 7 9 3 4 13 1 9 2 13 3 12 0 9 1 9 2
16 1 15 13 9 1 12 0 9 1 9 15 13 3 7 9 2
7 15 13 3 12 0 9 2
33 16 9 3 4 13 1 0 9 2 3 16 10 0 9 13 10 0 9 9 2 7 15 4 15 4 0 1 2 13 3 12 9 2
17 15 13 3 9 13 3 15 4 13 9 1 12 0 9 1 9 2
6 3 15 4 15 3 2
23 3 13 3 12 7 10 0 9 9 1 10 12 9 2 1 11 2 15 13 1 11 9 2
12 10 9 4 3 15 7 9 2 7 9 2 2
18 15 13 15 3 12 9 1 9 1 9 7 12 9 1 9 1 9 2
9 9 4 3 3 3 0 7 11 2
5 9 13 14 13 2
5 15 13 9 1 2
17 15 13 0 9 15 13 3 1 0 9 1 9 7 15 13 3 2
11 15 13 0 9 7 10 9 9 15 13 2
10 0 9 13 14 13 15 3 1 9 2
18 9 13 15 1 10 9 1 16 9 4 14 13 1 12 9 10 9 2
14 1 10 9 4 15 13 1 0 9 12 9 9 12 2
17 10 3 0 9 13 1 10 0 7 0 9 1 10 9 15 13 2
13 9 4 3 10 9 1 9 9 1 10 0 9 2
31 15 4 0 1 14 13 10 0 9 2 3 16 15 1 10 9 3 15 13 13 0 9 1 9 2 9 2 9 2 9 2
1 9
13 9 9 7 9 4 13 15 3 1 9 1 9 2
13 1 9 1 9 12 4 9 3 12 9 1 9 2
19 3 12 9 4 9 2 12 9 4 9 1 0 9 7 12 9 1 9 2
7 9 12 4 9 12 9 2
31 1 0 9 13 12 9 1 9 2 3 12 9 13 3 1 0 9 1 11 7 9 2 3 12 9 2 4 9 3 1 2
16 15 4 13 15 1 14 13 0 9 1 9 1 10 0 9 2
6 3 3 13 9 4 13
23 13 1 9 2 10 0 9 13 12 9 3 2 10 0 9 10 9 1 12 9 1 12 2
25 10 9 13 1 1 0 9 7 11 7 0 11 2 10 0 13 1 0 9 1 0 9 1 11 2
20 1 10 0 9 4 9 3 7 3 0 1 9 1 3 0 9 7 0 9 2
16 1 0 9 13 9 0 3 3 1 12 2 3 1 0 9 2
11 1 11 9 13 9 13 1 3 12 9 2
8 0 9 13 7 0 13 3 2
12 1 0 9 7 1 9 13 9 1 12 0 9
20 3 16 9 3 4 13 4 15 13 0 0 9 1 14 13 0 7 0 9 2
5 3 13 9 0 2
10 9 12 13 3 12 9 1 10 9 2
9 1 9 13 0 9 1 0 9 2
16 9 0 13 13 1 12 1 12 2 16 9 13 3 3 13 2
26 10 0 0 9 13 3 10 0 9 13 13 2 7 10 0 9 15 15 13 3 1 10 3 12 9 2
8 10 9 7 9 13 12 9 2
25 9 0 1 11 9 2 10 0 0 9 3 1 9 2 4 1 9 13 0 1 3 12 1 9 2
20 0 9 2 3 1 9 2 13 3 1 11 7 1 11 2 3 0 9 13 2
38 0 9 13 1 9 1 12 9 1 12 2 0 9 2 11 9 2 11 2 9 1 11 2 1 12 9 7 0 11 2 11 7 11 2 1 12 9 2
36 1 10 9 13 3 9 13 1 12 2 11 9 2 1 11 2 1 12 2 11 1 12 2 9 2 11 2 11 2 1 12 7 11 1 12 2
15 1 0 13 16 3 10 9 1 10 9 4 0 1 9 2
2 9 9
41 12 0 1 9 0 9 13 10 0 9 2 16 10 0 9 2 9 2 3 4 13 1 9 7 2 1 9 2 13 1 16 15 13 13 9 1 9 1 0 9 2
17 10 9 13 9 7 15 13 9 1 10 9 11 2 15 4 0 2
9 0 9 13 1 12 9 1 11 2
8 1 9 13 9 1 12 9 2
10 3 13 10 0 9 2 15 13 9 2
12 9 9 7 9 13 1 9 3 1 0 9 2
16 16 10 0 9 13 10 0 9 2 4 15 13 10 0 9 2
7 1 3 9 13 10 9 2
24 3 13 3 2 16 9 13 0 9 2 3 4 15 0 9 16 15 4 13 1 10 0 9 2
12 15 13 3 9 1 10 9 2 10 3 9 2
24 0 2 0 2 9 4 10 0 9 7 13 10 9 2 16 15 13 10 9 1 10 0 9 2
32 15 4 3 7 9 1 10 9 13 3 0 9 2 3 0 9 2 3 15 13 9 1 11 1 12 1 3 12 1 12 9 2
15 1 16 9 4 4 13 1 9 2 4 15 4 13 15 2
11 1 10 9 4 3 13 0 7 12 9 2
38 1 10 9 13 0 3 9 2 15 13 1 9 1 9 2 3 15 9 1 9 2 15 13 0 9 7 3 9 1 0 9 2 3 10 0 11 13 2
11 12 9 1 9 4 13 1 9 1 11 2
12 10 0 9 13 9 2 11 7 0 9 9 2
14 9 1 10 9 13 1 10 9 2 15 13 1 9 2
18 1 9 1 9 13 9 3 1 9 7 13 1 9 1 9 1 9 2
15 10 0 9 4 0 7 13 3 1 9 1 9 1 9 2
9 9 4 3 12 9 1 10 9 2
11 10 0 13 9 2 11 7 0 9 9 2
14 1 10 9 13 9 1 9 2 15 13 1 10 9 2
8 9 1 9 13 1 0 9 2
4 15 13 7 13
12 10 0 9 7 9 4 3 1 9 1 11 2
20 1 9 13 11 2 11 0 7 0 9 7 11 2 9 9 2 9 1 9 2
9 15 13 1 0 9 13 12 9 2
21 1 9 4 15 13 9 9 7 9 2 9 9 7 9 7 9 1 0 9 3 2
16 1 9 13 11 10 9 9 3 1 14 13 9 7 13 9 2
5 15 13 3 9 2
7 9 13 3 1 9 9 2
11 10 0 9 13 1 3 15 3 4 13 2
10 15 13 0 9 1 0 7 0 9 2
7 15 13 1 10 0 9 2
6 9 13 1 3 9 2
12 9 13 10 0 9 7 3 0 9 4 13 2
7 1 9 1 9 13 9 2
10 10 9 13 10 9 1 3 12 9 2
9 9 13 3 7 13 3 1 11 2
11 9 7 9 4 14 13 1 10 0 9 2
5 9 2 9 7 9
9 3 12 9 13 9 12 1 9 2
21 9 12 2 3 10 12 0 9 4 1 9 2 13 9 13 1 3 3 12 9 2
11 1 9 1 10 0 9 13 3 12 9 2
10 1 9 0 1 12 9 3 12 9 2
20 10 0 9 1 9 2 3 9 7 9 2 13 3 12 7 0 9 1 9 2
12 1 3 10 9 4 0 9 1 9 14 13 2
17 10 9 2 15 4 13 1 0 9 2 13 15 3 9 1 9 2
9 0 9 1 9 4 3 14 13 2
10 9 4 14 13 9 3 1 0 9 2
12 10 0 7 0 9 4 13 15 4 13 9 2
15 9 1 11 4 14 1 0 9 13 9 1 9 1 11 2
10 9 1 10 9 4 3 12 9 9 2
16 0 9 1 10 9 0 1 12 9 13 3 3 12 9 9 2
2 0 9
10 1 14 13 10 9 13 0 0 9 2
8 1 9 1 11 4 11 13 2
4 9 1 9 2
10 9 13 13 1 0 9 1 9 12 2
4 9 1 9 2
9 9 13 1 9 1 9 1 9 2
8 9 1 9 14 13 1 9 2
10 9 13 1 11 9 1 9 1 9 2
4 9 1 9 2
10 9 1 9 13 4 13 1 9 12 2
1 9
12 11 9 4 14 13 9 10 0 9 1 9 2
6 9 4 1 12 9 2
5 9 1 9 1 9
6 9 1 9 9 0 9
3 10 0 9
36 3 3 0 9 13 1 9 9 12 13 10 9 13 3 12 9 9 1 9 2 1 14 1 9 1 12 9 13 1 3 12 9 9 1 9 2
3 9 13 3
7 11 9 13 3 1 9 2
19 9 1 9 1 11 4 3 12 9 7 9 3 1 9 13 1 0 9 2
13 9 13 1 1 12 7 9 13 1 9 1 9 2
9 12 13 9 1 9 11 11 9 2
5 9 4 3 0 2
16 9 13 3 2 1 9 2 9 2 9 2 9 2 9 3 2
16 11 4 1 9 10 9 1 9 9 7 4 3 14 3 13 2
17 15 1 9 1 9 7 10 10 9 15 4 14 13 10 0 9 2
10 13 15 10 9 15 15 13 1 9 2
13 13 15 10 9 2 15 15 3 4 13 9 1 2
9 7 10 9 7 9 14 13 1 2
12 13 3 1 11 2 9 7 9 9 2 12 11
7 9 4 9 9 1 9 2
16 9 13 1 14 13 10 9 15 0 4 13 14 13 0 9 2
11 9 4 13 0 9 1 10 12 9 12 2
11 15 13 1 12 9 7 10 0 9 9 2
8 3 13 0 9 1 10 9 2
93 9 13 15 9 1 0 9 3 1 9 9 7 1 0 9 2 15 13 3 10 0 9 1 9 1 9 1 0 9 7 1 0 9 1 9 2 13 15 9 1 9 1 9 7 9 7 13 15 14 13 10 9 1 0 9 2 13 15 1 0 9 2 9 2 14 13 7 13 10 9 15 10 9 4 13 1 15 1 9 7 13 13 10 0 9 1 0 9 7 13 0 9 2
15 4 15 13 1 16 9 4 13 15 10 0 7 0 9 2
4 9 13 3 2
8 0 9 13 1 7 0 13 2
8 3 13 9 1 9 7 9 2
16 9 1 9 4 10 9 1 15 3 15 13 14 13 0 9 2
5 9 13 0 9 2
5 0 9 14 13 1
15 10 0 9 1 9 13 1 0 9 0 1 9 7 9 2
7 10 9 13 1 11 9 2
13 9 13 9 1 0 9 15 3 3 13 0 9 2
19 9 13 0 9 1 0 1 14 13 15 9 14 13 9 1 10 0 9 2
19 15 4 10 0 9 1 10 9 15 13 1 10 9 9 3 1 12 9 2
14 15 4 3 13 3 7 3 7 9 13 3 1 9 2
15 9 13 10 0 9 1 0 0 15 3 13 10 0 9 2
6 15 13 3 0 9 2
16 9 13 1 0 9 1 15 15 10 0 9 13 3 1 9 2
18 9 7 9 1 3 12 9 13 9 7 9 1 14 13 9 7 9 2
13 15 4 3 13 9 1 10 0 9 7 1 9 2
13 15 4 0 14 13 15 2 7 15 4 13 0 9
10 10 0 9 4 9 2 9 7 9 2
8 9 13 15 15 13 1 9 2
24 9 1 3 12 9 2 9 1 15 15 4 0 7 3 12 9 2 9 1 15 15 4 0 2
27 9 1 0 9 1 0 9 1 9 7 2 16 9 13 1 0 9 2 9 1 12 9 2 9 1 9 2
14 15 15 3 13 0 9 13 9 1 12 9 2 9 2
43 9 1 2 9 7 0 1 3 12 9 2 9 16 9 13 1 9 2 2 9 3 12 9 1 12 9 2 9 7 9 2 1 0 9 3 12 9 2 9 7 9 2 2
13 0 9 13 3 1 9 2 9 2 9 7 9 2
10 9 13 1 9 1 0 7 9 9 2
16 0 9 2 9 1 9 7 10 0 9 13 3 1 9 3 2
4 9 4 0 2
71 9 1 9 2 16 10 0 4 7 13 9 14 13 0 7 13 0 14 13 0 9 2 16 10 0 13 12 9 2 9 13 3 1 10 9 2 2 2 16 15 13 9 1 9 2 2 16 9 4 13 0 9 2 15 3 4 13 1 9 1 9 2 2 16 9 13 1 9 1 9 2
17 9 13 14 3 13 9 1 0 9 1 0 9 1 9 1 9 2
16 15 7 3 2 15 13 12 9 7 13 4 13 9 4 13 2
16 15 4 3 3 4 0 7 13 14 13 15 1 14 4 13 2
6 9 13 1 0 9 2
15 1 0 9 13 9 1 9 2 15 13 9 1 0 9 2
19 15 13 3 9 1 9 2 15 13 7 13 10 9 1 9 1 0 9 2
11 0 4 3 13 3 9 13 0 7 0 2
15 1 0 9 4 10 0 9 1 0 13 1 9 1 9 2
13 9 13 3 1 0 9 2 15 13 9 1 9 2
9 9 1 15 13 3 1 10 0 9
26 3 15 3 13 0 9 1 9 4 9 13 9 1 15 15 4 13 1 10 9 3 15 4 13 9 2
31 9 1 9 13 16 10 0 3 4 13 3 3 1 9 1 9 2 7 3 3 7 0 13 10 9 1 9 1 9 0 2
19 10 9 1 10 9 1 9 1 9 13 0 9 7 0 9 1 0 9 2
7 15 4 13 0 9 1 9
11 9 7 9 1 9 1 9 1 0 9 2
15 0 9 7 9 1 14 13 9 7 13 1 10 0 9 2
7 3 9 4 13 0 9 2
10 0 9 1 14 13 13 1 0 9 2
11 9 1 9 1 9 7 9 3 9 13 2
9 9 1 9 1 9 1 0 9 2
10 9 13 1 9 0 9 7 9 9 2
6 15 13 1 12 9 2
12 9 1 10 9 3 9 4 13 1 12 9 2
7 9 13 1 3 12 9 2
20 0 9 4 9 12 9 2 9 2 12 9 2 9 1 10 9 3 12 9 2
7 1 0 9 13 0 9 2
14 10 9 13 12 0 9 1 9 1 9 7 9 3 2
29 1 9 1 9 4 15 1 10 0 9 13 9 1 10 9 1 9 15 13 12 9 2 3 3 12 9 2 9 2
10 3 10 9 13 1 9 1 10 9 2
33 9 1 12 9 2 12 9 1 10 0 9 3 12 9 4 13 1 0 9 1 9 1 11 7 1 0 9 1 11 7 11 9 2
4 9 4 0 2
65 9 1 9 2 16 10 0 4 7 13 9 14 13 0 2 16 9 3 4 13 1 7 1 9 1 9 2 16 15 13 9 1 9 1 0 9 1 0 9 2 16 15 1 10 0 9 13 9 1 9 1 10 9 15 9 13 2 16 15 13 9 1 9 9 2
1 9
27 1 9 7 9 13 9 1 9 16 9 13 3 9 13 1 9 7 9 16 9 13 1 9 16 9 13 2
27 9 4 13 3 9 7 9 1 15 15 13 1 15 1 10 12 0 9 7 3 4 13 10 9 7 9 2
11 3 4 9 3 13 1 0 9 1 9 2
6 15 13 3 9 14 13
16 15 4 3 4 0 14 13 15 3 3 15 4 13 7 13 9
20 0 9 4 13 1 14 13 9 1 9 1 9 3 15 4 0 14 13 9 2
17 15 13 3 9 1 0 9 7 1 9 14 13 15 3 13 9 2
13 0 9 13 3 1 14 13 9 1 9 1 0 2
4 0 9 13 2
7 0 9 4 13 1 9 2
11 0 9 1 9 4 0 9 7 0 9 2
10 9 13 1 9 2 15 13 1 9 2
12 15 13 9 1 3 12 7 12 9 2 9 2
17 1 15 15 4 12 9 2 3 12 2 4 9 13 1 12 9 2
10 1 10 9 9 4 15 13 0 9 2
19 15 13 1 0 2 15 3 13 1 1 10 9 7 10 9 1 9 13 2
15 1 14 13 10 0 9 4 15 1 9 13 3 12 9 2
18 16 9 13 1 9 1 10 9 3 4 3 15 15 13 12 13 9 2
64 3 4 10 0 2 2 4 13 10 0 9 7 4 0 9 2 3 13 9 1 9 2 4 13 3 12 9 1 10 12 9 1 9 2 4 4 0 7 0 1 9 1 0 9 2 1 9 12 9 2 2 4 0 7 0 14 13 10 0 9 15 9 13 2
18 9 2 3 12 9 2 9 2 4 0 7 9 13 1 9 1 9 2
7 9 1 12 9 13 9 2
16 1 15 15 13 0 14 13 9 1 0 9 4 9 13 0 9
16 0 9 13 1 0 7 15 15 3 4 13 9 1 0 9 2
5 9 9 13 3 2
8 1 0 9 4 3 9 13 2
4 9 1 9 2
15 0 1 9 14 13 15 1 10 9 13 9 14 13 9 2
6 9 13 1 0 9 2
9 9 4 13 1 9 1 0 9 2
8 9 13 1 10 0 9 9 2
25 0 7 0 9 13 0 2 15 1 0 9 3 4 13 9 1 10 0 9 2 9 1 10 9 2
15 10 0 9 13 1 9 1 9 7 13 9 1 0 9 2
14 10 0 9 13 3 9 1 7 1 0 9 1 9 2
9 9 7 9 13 1 10 0 9 2
5 9 1 0 9 2
24 9 15 13 9 1 0 9 4 13 9 1 12 9 1 9 7 9 16 9 13 1 9 9 2
30 9 4 13 1 0 2 0 7 0 9 2 15 3 4 13 10 0 9 1 10 0 9 2 7 15 4 13 0 9 2
19 9 4 3 13 1 0 1 14 13 9 7 9 7 1 0 9 1 9 2
22 16 10 0 1 10 9 2 7 1 14 4 13 1 9 13 9 4 9 7 9 13 2
13 3 15 13 9 4 15 13 3 0 9 7 0 2
23 15 13 3 0 0 9 1 9 7 1 9 7 1 0 9 13 15 3 0 9 1 9 2
23 13 15 1 15 15 13 13 9 1 9 3 4 15 3 13 13 1 3 15 4 13 3 2
19 15 4 3 13 9 7 13 13 3 16 15 13 0 7 0 14 13 9 2
36 15 13 3 3 3 9 1 0 9 15 4 0 1 9 14 13 10 0 9 2 15 4 3 13 1 9 2 9 7 3 9 13 15 1 9 2
14 7 3 15 13 3 1 2 7 0 9 4 15 13 2
3 13 7 13
18 15 13 3 15 4 13 16 15 13 9 1 10 9 1 14 13 9 2
11 15 15 4 0 14 13 3 1 4 13 2
27 4 15 1 9 13 10 0 9 7 15 15 13 9 1 2 13 15 15 1 9 1 9 1 9 7 9 2
24 13 15 3 9 1 0 9 7 3 1 10 9 15 15 3 13 3 3 1 13 3 0 9 2
23 3 4 15 13 3 1 9 7 3 13 7 9 7 9 1 14 13 3 15 15 4 13 2
25 3 15 13 3 7 13 0 9 1 9 7 1 9 4 15 3 0 16 15 13 10 9 15 13 2
9 1 14 13 4 15 3 13 3 1
3 9 7 9
3 9 1 9
1 9
3 9 7 9
3 9 1 9
4 9 9 7 9
1 9
2 0 9
7 9 4 13 9 1 15 2
17 15 4 3 13 10 9 15 13 1 9 12 1 14 13 0 9 2
4 3 14 13 0
14 3 4 15 0 14 0 13 3 10 9 15 15 13 2
10 9 13 1 13 3 9 1 0 9 2
10 7 1 9 7 1 0 9 1 9 2
22 1 0 9 13 9 3 0 9 7 1 9 9 13 10 9 1 0 9 1 0 9 2
6 3 13 15 3 1 9
20 1 16 15 3 4 13 10 9 13 15 16 15 13 1 15 15 13 14 13 2
12 3 13 15 3 1 9 1 10 9 0 9 2
18 1 9 9 4 15 3 1 10 9 13 1 10 9 1 9 7 9 2
28 9 4 3 13 15 1 9 7 1 9 1 9 1 0 9 7 1 16 15 4 4 13 10 9 1 0 9 2
2 13 3
14 15 4 0 14 1 0 9 13 13 15 1 1 9 2
16 13 9 1 9 16 15 4 0 1 15 15 4 13 1 9 2
22 13 15 13 10 9 14 3 13 1 0 9 2 7 15 13 3 13 10 3 0 9 2
87 9 13 15 9 1 0 9 3 1 9 9 7 1 0 9 2 15 13 3 10 0 9 1 9 1 9 1 0 9 7 1 0 9 1 9 13 15 9 1 9 1 9 7 9 7 13 15 14 13 10 9 1 0 9 13 15 1 9 14 13 7 13 10 9 15 10 9 4 4 1 15 1 9 7 13 13 10 0 9 1 0 9 7 13 0 9 2
7 11 13 1 10 9 7 9
5 9 1 9 7 9
1 9
1 9
1 9
5 9 7 9 1 9
12 15 4 0 14 13 3 1 3 15 13 9 2
20 9 4 10 0 9 7 3 13 15 15 14 13 1 1 9 1 9 7 9 2
5 11 4 10 9 2
24 15 4 9 9 15 1 0 9 13 1 9 2 12 11 12 11 12 11 12 11 12 11 12 11
26 9 4 3 13 3 2 13 10 12 7 13 15 3 1 0 9 2 3 1 14 13 13 1 0 9 2
6 1 9 4 9 13 2
12 3 13 15 1 9 2 9 2 9 2 9 2
18 12 0 9 7 11 3 11 7 11 4 3 0 1 11 1 3 9 2
14 11 4 3 3 0 16 11 13 15 1 10 0 9 2
19 11 4 13 3 10 0 0 9 2 15 13 9 9 9 14 13 1 9 2
8 13 1 11 11 9 3 3 2
10 15 4 9 2 0 2 0 2 0 2
24 3 4 15 13 9 1 9 7 0 9 4 13 1 10 9 2 3 7 1 10 9 1 11 2
5 15 13 1 15 2
18 15 13 1 10 9 1 14 1 9 4 13 0 0 9 1 9 9 2
8 10 3 0 9 13 1 11 2
18 2 15 15 13 16 11 4 13 7 10 9 9 1 9 4 3 0 2
21 3 11 11 13 1 11 10 9 12 13 15 10 9 15 13 1 11 9 3 3 2
17 2 4 15 13 1 1 11 3 4 15 3 13 1 1 11 3 2
6 2 15 13 3 15 2
8 3 4 0 0 9 13 2 2
8 1 11 11 13 9 1 11 2
19 3 3 13 15 16 11 4 13 10 3 0 9 1 15 9 3 4 13 2
4 15 4 11 9
21 15 4 9 1 9 2 1 9 9 7 3 2 10 9 11 3 4 13 3 1 2
2 9 2
11 3 13 12 9 1 15 7 15 1 9 2
17 3 0 9 13 4 15 9 2 3 9 13 3 4 15 9 3 2
7 15 4 9 9 1 11 2
8 9 13 9 1 10 0 9 2
3 9 9 2
7 13 1 12 3 0 9 2
17 10 0 9 2 15 3 13 10 0 9 1 9 2 13 3 2 2
4 0 9 9 2
18 10 9 13 1 3 0 7 0 9 2 12 1 15 7 15 1 9 2
14 10 9 13 1 10 9 1 15 10 9 1 12 9 2
8 9 9 4 13 3 7 3 2
21 15 13 0 9 1 9 7 9 7 13 10 9 0 0 9 15 9 3 13 1 2
3 11 9 2
8 4 3 0 1 10 0 9 2
26 13 1 12 9 15 13 1 16 10 9 13 2 13 9 1 9 2 4 0 9 1 11 0 9 3 2
7 9 13 10 3 0 9 2
10 10 9 1 0 9 4 15 3 13 2
2 9 2
3 11 9 2
15 13 1 12 9 15 13 1 10 3 9 9 2 9 2 2
17 9 13 0 0 9 2 0 9 2 9 2 9 2 9 2 9 2
7 9 9 4 3 0 0 2
23 15 4 3 13 1 10 9 0 9 16 9 13 9 2 7 9 4 3 0 1 9 9 2
2 9 2
6 15 4 10 0 9 2
28 1 9 13 9 7 10 9 1 10 9 2 1 0 0 9 2 7 3 4 15 13 1 10 0 2 9 2 2
13 9 13 1 9 12 9 7 3 3 7 12 9 2
21 1 9 4 3 9 1 9 13 1 10 0 9 7 4 3 10 0 7 0 9 2
9 15 4 13 9 1 0 0 9 2
9 13 9 1 9 7 13 9 3 2
15 9 13 9 1 7 9 2 10 9 7 10 0 9 9 2
29 9 4 0 1 9 7 9 15 15 1 15 13 3 9 2 9 2 9 2 9 15 13 9 7 9 2 11 3 2
12 1 15 13 10 9 0 9 0 1 12 9 2
9 10 9 4 13 3 3 1 9 2
23 15 13 3 0 7 15 4 3 13 10 9 1 9 2 15 4 3 13 15 10 1 9 2
14 3 2 1 10 9 13 10 9 9 1 10 0 9 2
21 9 4 9 1 3 9 2 15 13 3 7 3 1 10 3 9 7 9 1 11 2
8 15 13 1 16 15 13 1 2
12 15 13 3 3 0 16 11 13 1 1 11 2
23 6 2 9 11 11 2 9 11 11 2 9 11 11 3 4 3 7 3 13 9 1 9 2
14 9 11 11 3 13 3 10 9 1 10 0 9 9 2
22 3 4 15 13 13 3 12 9 2 9 1 9 1 0 9 7 15 3 13 9 0 2
10 3 13 15 9 1 15 1 0 11 2
5 15 4 3 0 2
12 7 11 13 9 1 9 7 15 4 13 3 2
11 10 0 0 9 4 3 0 9 11 13 2
20 3 11 13 3 1 9 13 10 12 0 2 11 2 11 7 11 12 9 15 2
12 11 7 11 13 12 9 15 7 11 12 9 2
6 1 9 13 12 9 2
11 10 12 0 4 3 13 3 10 12 0 2
21 7 3 12 0 7 12 0 2 11 7 11 2 4 13 3 12 0 7 12 0 2
21 16 11 2 11 2 11 7 11 15 13 9 1 11 13 1 4 15 13 0 9 2
8 11 9 4 3 13 0 9 2
11 11 2 11 2 11 7 11 12 9 15 2
19 11 2 11 12 9 15 2 11 12 2 11 2 11 7 11 12 9 15 2
6 3 13 15 12 9 2
9 1 0 9 13 12 9 1 12 2
9 10 9 4 3 13 1 12 9 2
4 7 11 3 2
9 6 2 15 4 3 13 9 3 2
5 15 13 9 0 2
8 7 15 4 13 3 1 11 2
18 7 13 15 1 2 3 13 15 1 16 15 1 0 9 13 12 9 2
6 12 9 1 9 1 11
2 3 2
7 11 13 10 0 9 9 2
10 3 11 13 1 9 4 15 13 1 2
15 0 4 3 15 4 13 12 2 15 15 13 10 9 1 2
6 15 13 3 1 0 2
22 11 0 9 4 9 12 14 13 3 12 9 9 2 3 0 0 13 3 10 9 2 2
21 1 9 13 15 3 12 9 9 7 1 9 12 9 9 2 3 13 15 12 9 2
6 15 13 3 0 9 2
23 3 4 15 3 12 13 10 9 13 3 10 9 1 9 7 9 1 10 0 9 1 11 2
16 3 4 10 9 1 10 9 13 3 3 12 9 1 10 9 2
4 9 4 0 2
32 1 11 9 4 15 13 16 15 3 0 13 1 9 1 10 0 9 14 15 0 13 3 3 15 13 12 9 1 9 1 9 2
35 10 3 0 4 3 3 3 10 11 15 13 1 9 7 10 11 15 15 4 14 13 16 11 2 11 2 11 2 11 7 3 11 13 1 2
7 2 15 13 9 1 9 2
9 3 4 3 10 0 9 13 11 2
11 11 13 3 9 14 13 3 10 9 3 2
15 1 10 9 13 3 10 9 1 11 1 11 11 0 9 2
2 3 2
31 2 13 15 3 9 2 3 13 15 1 15 9 2 9 7 9 7 3 13 15 9 1 9 7 0 11 9 13 1 9 2
2 9 2
14 11 2 0 0 9 2 10 0 9 2 10 12 2 2
11 11 2 0 0 9 9 2 10 0 9 2
10 11 2 0 11 9 9 2 9 2 2
4 10 9 1 11
9 1 10 12 9 13 12 9 9 2
10 10 9 1 0 9 3 1 11 9 2
13 1 10 0 9 11 7 11 13 3 12 9 9 2
11 1 10 12 0 9 3 11 13 12 9 2
21 13 11 2 11 2 11 2 11 7 11 1 3 13 11 1 3 3 12 9 9 2
15 1 10 9 9 3 11 3 13 4 15 13 3 3 3 2
12 10 0 9 1 11 9 3 4 4 3 0 2
11 9 9 1 11 1 12 13 1 12 9 2
9 1 11 4 15 10 9 12 9 2
8 1 11 4 9 3 12 9 2
33 9 2 10 0 9 1 15 10 9 13 1 9 1 9 7 9 2 4 13 1 12 9 9 12 1 11 2 1 12 9 1 11 2
11 11 13 1 10 9 10 9 1 12 9 2
15 10 0 9 4 0 2 12 9 1 11 1 9 1 9 2
15 3 4 15 13 3 2 7 4 3 0 2 3 12 9 2
17 1 0 9 13 10 0 9 1 10 9 0 9 1 9 7 9 2
6 9 4 13 1 9 2
21 7 9 4 3 3 13 3 7 9 4 13 3 2 3 3 3 3 7 1 11 2
10 15 13 1 9 16 11 4 13 0 2
12 15 13 1 12 11 2 12 11 7 12 11 2
23 1 16 11 4 4 13 15 7 13 1 9 4 15 13 2 11 13 2 13 3 0 9 2
4 10 0 9 11
14 9 12 9 9 9 12 9 9 12 9 0 9 9 9
3 15 4 9
9 10 12 9 12 13 7 11 9 2
20 9 1 10 9 13 1 9 15 10 12 9 13 1 10 12 9 12 1 11 2
16 15 13 1 10 9 1 11 12 15 11 9 11 11 13 9 11
5 9 12 9 7 9
18 0 9 1 9 13 1 9 15 3 13 9 9 11 11 9 9 0 9
45 1 15 13 10 9 9 2 3 9 1 9 2 9 2 9 3 2 15 7 15 1 12 9 2 3 10 9 1 9 2 9 4 9 15 13 3 7 3 1 11 7 10 3 9 9
48 0 9 2 9 15 13 0 1 0 9 2 9 0 9 2 9 1 11 2 0 9 0 9 2 9 3 2 0 9 1 9 0 9 0 9 0 9 0 0 9 9 9 9 2 11 0 9 2
16 10 3 0 9 1 9 13 16 0 9 13 3 0 1 9 2
20 16 15 3 4 9 13 3 1 16 15 3 13 3 0 15 4 14 13 1 2
12 1 12 9 3 12 9 4 12 9 1 9 2
12 7 1 10 12 13 3 12 1 9 1 9 2
6 10 0 12 13 3 2
6 7 15 13 3 9 2
21 1 14 13 10 9 4 15 4 13 10 9 1 1 0 9 3 12 9 1 9 2
9 15 4 3 0 14 13 1 9 2
9 3 4 10 0 9 13 1 9 2
11 15 15 13 1 9 13 12 9 1 9 2
10 10 0 12 9 13 1 9 7 9 2
15 1 9 13 15 1 9 12 9 1 3 0 9 1 9 2
6 12 9 13 15 1 2
6 12 9 4 0 9 2
1 9
8 9 1 0 9 4 3 0 2
10 15 13 15 15 13 3 9 1 9 2
10 15 13 3 15 15 13 12 9 3 2
6 9 9 13 1 9 2
13 3 10 9 15 12 9 1 10 0 13 1 9 2
26 15 15 13 1 12 1 9 7 13 1 10 9 1 9 13 12 9 1 9 1 14 13 9 1 9 2
12 10 0 9 1 9 4 13 1 9 1 9 2
7 3 13 15 10 9 12 2
10 10 0 9 1 14 13 1 9 4 2
5 9 1 9 13 2
9 9 14 4 13 1 3 9 13 2
5 9 4 13 13 2
11 7 15 13 16 3 10 0 9 13 3 2
2 9 9
8 7 0 4 3 10 0 9 2
10 10 9 4 4 10 9 1 9 9 2
15 10 9 9 13 16 9 0 9 4 3 0 7 10 9 2
9 10 9 13 3 3 1 0 9 2
11 7 15 13 3 0 9 1 14 4 9 2
22 10 7 0 9 13 16 15 4 0 14 13 9 0 9 0 9 1 9 7 3 0 2
17 15 13 15 13 3 14 13 1 9 9 3 16 10 0 9 13 2
14 15 4 3 0 14 13 3 1 9 7 14 13 1 2
14 15 15 13 10 9 7 13 9 1 9 13 3 9 2
9 9 1 0 9 13 3 1 9 2
9 10 0 9 4 13 3 0 9 2
7 9 4 3 3 13 9 2
6 1 0 9 13 9 2
10 3 3 0 4 15 14 13 1 9 2
7 9 13 1 10 0 9 2
6 9 13 13 1 9 2
14 15 15 13 3 9 1 9 13 3 0 9 0 9 2
13 7 15 13 3 0 9 1 14 13 1 1 9 2
17 3 13 15 3 3 3 2 16 15 3 13 1 9 9 1 9 2
12 15 13 3 10 9 9 7 13 3 3 3 2
24 14 13 1 9 9 1 9 13 1 15 7 0 1 14 13 1 9 7 13 3 10 0 9 2
12 7 10 0 4 16 15 4 0 7 0 1 2
4 13 3 1 9
12 15 13 10 0 9 2 10 0 13 10 9 2
11 10 9 9 7 9 4 15 13 9 1 2
23 13 3 9 2 13 9 2 13 9 7 13 1 16 15 13 9 3 1 14 13 0 9 2
12 13 9 4 15 13 3 16 15 13 1 9 2
17 3 15 13 1 9 2 1 12 9 9 2 16 15 1 9 13 2
5 15 4 0 0 2
9 1 12 9 4 9 13 0 9 2
25 1 9 4 15 13 1 1 15 16 15 13 10 9 2 1 12 9 2 1 16 9 4 13 0 2
30 10 0 9 14 13 3 9 1 9 7 13 9 4 0 2 3 4 15 3 13 16 0 9 13 2 7 3 3 3 2
15 7 9 4 15 1 10 3 0 9 1 9 3 3 9 2
26 16 15 13 1 9 3 2 3 1 9 2 4 15 3 3 13 9 10 0 9 1 14 13 0 9 2
3 13 9 0
6 9 4 15 13 0 2
24 13 15 9 13 15 9 14 13 1 15 2 15 13 9 3 0 9 1 15 15 13 1 11 2
9 9 15 13 0 9 4 3 13 2
8 13 1 3 0 9 15 13 2
10 3 4 15 4 3 12 9 1 9 2
21 4 15 12 4 15 13 3 12 9 2 7 3 4 15 13 1 9 7 13 0 2
15 15 4 3 0 0 14 13 0 9 1 9 3 9 13 2
10 9 13 7 9 3 1 3 0 9 2
15 9 1 9 15 15 4 13 1 9 2 9 15 4 13 2
15 9 2 13 15 3 0 2 13 1 10 3 0 9 2 2
9 9 2 3 10 9 1 9 2 2
25 9 2 15 4 13 15 0 2 7 4 9 13 3 7 13 7 13 4 15 10 9 1 9 2 2
23 15 13 16 15 4 0 3 1 9 16 15 13 3 9 13 2 0 3 2 0 3 3 2
14 15 4 3 0 16 9 13 1 10 9 7 0 9 2
8 3 13 9 3 7 9 13 2
6 13 0 9 1 9 2
10 15 4 3 0 7 14 13 1 9 2
20 13 3 9 2 13 1 0 9 1 0 9 2 1 9 15 13 9 7 9 2
17 4 9 13 3 13 15 3 2 3 13 9 1 9 1 10 9 2
9 15 4 13 9 0 16 9 13 2
13 15 13 9 2 13 3 10 9 2 1 10 9 2
33 4 15 9 3 4 15 13 1 16 9 4 3 0 16 15 13 3 2 3 13 9 2 9 13 0 14 13 2 9 13 3 3 2
25 15 13 1 15 3 15 4 13 3 1 9 2 3 16 15 13 10 9 1 0 9 7 0 9 2
3 13 9 2
17 15 13 3 12 9 14 13 0 9 2 7 15 13 15 9 1 2
9 9 4 13 10 9 3 1 9 2
24 1 9 2 15 13 3 0 1 0 9 2 13 15 10 9 2 15 13 3 10 9 9 2 2
6 13 16 9 13 3 2
3 1 9 2
6 13 3 10 0 9 2
4 13 1 9 2
10 13 9 2 0 9 2 0 14 13 2
11 13 9 2 15 4 4 0 7 3 0 2
4 9 2 9 2
10 3 9 13 7 9 13 9 1 9 2
8 3 15 13 9 13 9 1 2
13 15 13 9 2 13 1 9 2 14 13 1 9 2
4 15 13 9 2
14 9 4 4 3 0 2 13 10 9 14 13 1 9 2
21 15 4 3 10 0 9 15 3 13 10 9 1 10 12 9 9 13 13 1 15 2
4 13 3 9 2
10 1 9 4 15 13 0 9 1 9 2
16 13 3 9 2 13 0 2 13 3 0 9 7 13 1 9 2
10 3 9 2 13 9 7 9 1 9 2
6 15 4 0 7 0 2
12 13 3 0 9 1 9 2 16 9 13 3 2
2 9 2
9 13 3 10 9 1 9 7 9 2
72 13 1 16 15 13 0 9 1 9 2 12 0 9 12 9 2 13 3 7 12 9 2 12 9 2 13 10 9 9 2 12 9 12 0 9 12 9 2 2 13 3 12 9 2 2 0 14 13 16 15 13 1 9 2 4 13 2 7 13 0 1 9 2 12 0 9 2 13 12 9 2 2
20 6 2 13 15 1 14 13 15 3 1 9 2 4 15 13 0 9 1 9 2
4 15 13 0 2
18 15 4 3 14 13 3 0 16 15 13 0 16 15 13 3 1 9 2
5 12 9 14 13 3
8 9 2 13 9 2 13 9 2
4 9 7 9 2
14 9 4 4 1 0 9 2 0 9 13 1 9 9 2
20 1 9 2 9 2 9 1 9 2 13 9 2 0 9 2 2 9 1 9 2
13 9 13 0 2 9 1 9 4 3 0 7 9 2
3 13 9 2
7 13 9 2 9 7 9 2
8 13 0 9 1 2 13 9 2
25 3 9 4 0 1 2 13 16 15 2 13 3 2 2 16 9 4 0 2 16 15 13 7 13 2
18 13 10 9 1 9 15 13 1 9 7 15 13 9 1 14 13 3 2
6 13 9 2 13 9 2
19 9 13 13 3 3 2 13 9 3 0 1 0 9 2 13 1 10 9 2
5 4 13 10 9 2
20 13 16 9 4 0 3 3 2 9 2 9 2 0 9 2 9 2 0 9 2
31 16 15 13 9 1 11 7 1 10 2 0 2 9 1 11 3 13 15 11 11 1 11 2 11 2 15 4 13 3 15 2
12 11 4 11 0 2 9 9 2 2 0 3 2
30 1 0 9 3 13 15 7 9 1 10 9 15 9 9 2 0 1 9 7 9 3 2 13 1 10 0 9 1 9 2
15 15 4 3 14 13 1 9 3 1 11 2 3 1 11 2
25 3 10 0 9 13 2 3 1 9 11 2 11 2 11 2 13 9 1 9 1 9 1 0 9 2
12 10 9 4 14 13 1 9 3 12 9 9 2
14 3 1 9 13 15 3 0 2 3 12 9 1 9 2
13 15 13 9 15 13 1 10 7 3 9 1 9 2
6 9 13 3 7 13 2
16 9 4 13 3 9 1 10 0 9 0 2 0 7 0 9 2
13 15 4 13 3 7 1 15 4 15 3 13 9 2
27 9 2 15 13 1 12 9 3 2 13 1 0 9 12 9 14 13 1 1 7 9 14 13 3 12 9 2
25 10 0 9 9 4 13 3 1 10 9 1 0 9 15 13 2 1 9 2 1 9 7 1 9 2
8 7 10 3 0 9 13 3 2
4 12 9 13 9
19 15 13 1 9 1 9 3 9 4 13 3 11 11 4 13 10 0 9 2
16 3 4 10 9 1 9 13 16 15 13 9 1 10 0 9 2
6 15 4 3 13 9 2
8 1 9 4 15 3 13 9 2
19 15 4 3 3 0 1 10 1 10 0 3 12 9 1 9 15 4 13 2
8 9 1 10 0 9 13 3 2
20 16 9 13 7 9 4 3 0 16 15 4 3 13 13 9 10 9 1 9 2
16 15 13 1 10 3 9 1 12 15 13 1 1 10 3 9 2
4 9 1 12 9
12 0 9 13 3 14 13 3 7 12 0 9 2
15 16 10 9 13 15 4 0 3 13 9 1 9 12 9 2
21 3 9 11 2 11 2 11 4 0 13 9 13 1 10 9 1 11 3 1 11 2
15 15 4 13 1 9 1 11 3 7 3 3 7 12 9 2
18 3 13 15 1 0 7 0 9 3 1 0 9 1 3 12 9 9 2
5 9 4 3 13 2
11 3 4 15 13 13 1 9 3 10 9 2
9 7 3 4 3 9 0 1 9 2
12 9 13 3 3 1 9 3 1 9 1 12 2
4 9 9 7 9
10 11 11 4 13 1 0 9 1 9 2
19 3 13 15 1 11 9 7 11 2 15 13 1 11 7 0 9 1 9 2
6 15 13 15 1 11 2
7 6 2 15 13 3 0 2
16 7 3 1 11 13 0 9 1 9 2 0 9 2 0 9 2
19 2 9 4 14 13 9 7 9 7 4 13 7 12 12 9 2 13 15 2
13 15 4 13 1 1 9 12 9 9 1 10 9 2
20 1 14 13 10 9 13 10 9 9 2 15 4 9 0 9 7 3 10 0 2
7 3 13 0 9 1 9 2
19 16 9 13 15 3 1 9 13 9 3 1 9 3 16 9 3 13 3 2
29 3 9 13 13 10 0 9 2 7 1 16 3 9 4 13 3 3 1 9 13 9 1 9 7 10 9 0 9 2
7 15 4 11 13 9 1 2
14 9 1 9 13 3 3 1 9 3 1 9 1 12 2
17 2 10 9 2 0 3 12 9 9 2 13 3 7 13 1 9 2
30 15 13 10 9 1 3 12 9 15 13 1 9 2 12 9 9 1 9 1 12 9 9 13 1 10 9 9 1 9 2
24 9 1 9 14 13 9 1 9 1 11 7 11 13 3 16 11 13 9 1 12 9 9 3 2
22 15 4 10 0 9 1 9 15 10 0 9 4 4 13 3 2 1 0 9 3 13 2
17 7 7 11 11 7 10 0 13 3 16 9 4 14 13 10 9 2
7 11 11 13 9 1 11 2
6 9 9 13 0 9 2
6 3 15 13 13 15 2
11 10 0 9 4 4 13 1 10 0 9 2
9 9 0 4 0 1 3 0 9 2
11 15 13 0 9 15 11 4 13 1 9 2
7 9 13 3 0 7 0 2
11 9 1 9 2 9 7 9 4 3 0 2
9 1 10 9 13 10 9 0 3 2
13 9 1 9 4 13 9 1 12 9 2 2 2 2
15 7 9 4 13 16 10 9 1 0 9 13 3 1 12 2
20 11 0 9 1 9 2 9 11 11 11 2 1 11 0 9 2 13 1 11 2
8 2 10 9 4 0 1 9 2
8 9 4 15 3 3 13 1 2
6 9 4 7 0 9 2
16 10 9 4 1 9 1 0 9 13 10 9 7 12 15 3 2
6 9 4 15 13 15 2
21 10 9 2 3 9 2 15 3 13 1 9 1 9 7 9 13 12 1 12 9 2
8 9 13 9 7 9 1 9 2
3 9 11 2
15 2 1 10 0 9 13 10 0 9 1 9 9 1 3 2
12 10 9 4 4 3 13 3 1 10 0 9 2
7 15 13 3 9 15 13 2
11 9 1 9 13 3 9 1 10 9 3 2
12 1 9 3 9 9 13 13 13 9 3 0 2
12 9 0 13 10 9 1 16 15 13 0 9 2
11 9 15 15 4 14 4 13 1 3 3 2
11 9 11 4 13 1 14 13 9 3 0 2
13 1 12 9 3 13 15 3 2 9 1 9 2 2
10 10 9 15 13 1 9 7 0 9 2
13 11 4 0 1 9 9 15 4 0 1 10 9 2
6 1 9 13 9 9 2
18 3 13 3 3 10 9 1 3 9 2 13 3 1 10 0 9 2 2
12 15 4 3 13 15 3 0 1 9 1 9 2
11 9 4 4 13 1 9 1 10 0 9 2
18 1 10 9 1 12 9 13 15 3 3 1 10 9 1 9 1 9 2
9 9 11 4 0 1 9 1 9 2
12 2 9 1 0 9 1 10 0 4 13 3 2
10 10 0 9 13 3 3 14 4 0 2
12 3 4 15 13 16 15 4 10 9 1 9 2
9 9 4 3 13 9 14 13 9 2
16 1 9 12 1 11 13 10 9 1 10 9 9 1 0 9 2
13 15 13 16 9 13 1 9 1 10 9 1 11 2
17 3 13 15 1 0 9 9 7 13 3 16 9 9 13 0 9 2
10 15 4 15 3 0 1 1 10 9 2
9 9 4 4 0 1 10 0 9 2
5 15 13 1 11 2
20 2 15 4 13 3 0 9 13 1 9 1 9 1 14 4 13 15 15 13 2
10 15 4 3 10 9 4 4 13 1 2
8 9 1 10 0 4 3 0 2
26 15 13 3 9 1 10 0 9 2 7 7 13 3 10 0 9 7 3 13 15 15 3 1 10 0 2
14 9 4 9 1 9 7 9 1 9 7 9 1 9 2
25 15 4 13 9 1 9 2 3 7 9 7 1 9 9 2 1 14 13 10 0 9 1 9 9 2
8 10 0 9 4 3 4 13 2
11 9 11 13 1 10 9 1 10 0 9 2
9 9 1 10 0 4 10 0 9 2
6 9 13 15 3 0 2
8 3 4 0 9 13 3 3 2
2 9 2
17 10 0 9 2 9 2 9 3 2 4 3 0 1 10 0 9 2
16 3 4 15 3 3 4 13 1 10 0 9 15 15 13 9 2
9 9 13 3 1 10 9 1 9 2
21 10 0 15 13 2 0 2 9 4 13 1 3 12 9 16 15 13 3 0 9 2
10 9 4 3 13 3 0 9 1 9 2
9 10 9 4 4 13 1 3 3 2
15 9 13 3 3 1 12 1 12 9 15 13 1 10 9 2
9 10 0 9 15 13 1 0 9 2
26 2 1 10 10 9 9 9 15 1 12 9 3 13 9 1 11 4 3 1 9 10 0 9 13 13 2
20 16 15 12 13 3 12 9 1 15 9 4 10 9 1 9 13 1 12 9 2
18 15 4 10 9 15 15 3 13 13 1 3 15 13 1 9 10 9 2
19 15 13 15 1 9 0 9 2 9 11 11 2 1 10 9 1 9 9 2
19 9 11 4 9 1 0 9 1 9 7 9 2 10 0 9 9 1 9 2
28 9 11 4 13 1 1 15 1 10 0 9 15 13 1 9 7 13 1 11 2 9 2 7 9 1 10 9 2
11 15 4 3 1 10 9 9 9 1 11 2
21 10 0 9 1 9 14 13 0 9 14 13 13 13 1 9 11 1 10 9 9 2
21 15 13 1 12 9 3 2 3 9 13 1 9 2 1 10 9 1 3 0 9 2
27 13 1 1 9 16 9 4 0 2 13 1 10 0 9 3 15 4 13 13 2 13 10 0 9 9 13 2
25 2 9 13 16 9 3 7 3 13 13 1 3 15 3 13 1 14 13 10 9 2 13 9 11 2
2 9 13
18 3 13 9 11 10 3 0 9 1 3 3 9 7 10 9 7 9 2
15 10 9 9 2 9 2 9 2 9 7 0 9 13 13 2
19 15 13 16 15 4 0 14 13 0 9 14 13 13 16 10 0 13 9 2
31 9 13 3 1 9 3 15 0 4 13 15 15 4 1 9 9 2 3 15 13 2 10 9 15 4 13 16 15 4 13 2
24 2 1 12 7 10 0 9 3 13 15 3 9 1 9 1 10 9 1 9 2 13 9 11 2
22 15 13 3 16 10 9 4 13 10 9 1 9 15 13 1 9 1 10 9 9 13 2
10 7 10 9 4 13 10 3 0 9 2
17 1 9 11 4 10 10 9 13 15 1 10 9 1 9 1 11 2
23 15 1 10 9 2 3 9 13 13 1 3 3 3 9 4 0 7 10 0 9 1 9 2
3 9 1 9
37 2 7 0 15 4 13 9 14 13 3 15 3 13 2 10 9 15 13 13 1 9 2 3 0 4 15 14 13 15 14 13 13 2 13 9 11 2
4 9 4 9 2
19 1 9 11 4 15 10 9 9 1 9 1 11 1 14 13 13 3 9 2
16 0 0 9 3 4 13 13 9 16 9 4 0 1 0 9 2
8 15 1 14 13 13 0 9 2
17 2 10 0 9 4 1 10 0 12 9 13 13 2 13 9 11 2
16 1 10 9 4 15 3 0 1 15 14 13 15 14 13 13 2
12 9 4 3 13 13 3 0 1 14 13 9 2
3 9 11 2
20 2 10 12 9 0 9 4 15 0 14 13 9 1 9 1 0 9 7 9 2
15 3 4 10 9 3 0 1 9 2 1 9 7 9 3 2
11 7 9 13 9 11 4 4 14 13 3 2
4 16 15 4 13
16 2 10 9 1 9 4 13 10 0 0 9 1 9 1 9 2
9 10 9 13 10 9 9 7 9 2
19 15 4 1 9 13 9 16 9 4 0 1 9 7 1 0 9 3 0 2
22 10 0 9 13 1 9 11 16 15 3 3 4 0 14 13 10 9 9 14 13 13 2
26 2 7 1 15 15 3 4 13 13 3 13 15 3 10 0 9 1 9 14 13 13 15 14 13 3 2
9 9 1 10 9 13 1 9 11 2
14 13 3 1 10 9 15 13 0 9 1 9 7 9 2
4 13 0 9 2
7 13 0 9 1 10 9 2
4 13 3 9 2
4 9 11 11 2
14 2 15 13 15 14 13 13 3 16 15 13 3 3 2
33 9 11 11 13 1 3 10 9 3 1 10 9 1 11 2 13 9 1 9 2 13 1 9 1 10 9 2 3 9 3 13 9 2
31 15 13 0 9 7 13 1 10 9 2 14 13 10 0 9 2 15 13 9 1 9 7 9 1 16 9 4 13 10 9 2
21 1 9 13 15 7 9 7 9 15 13 9 2 15 4 0 16 15 13 1 11 2
9 7 1 9 1 9 4 15 0 2
11 3 13 1 9 1 9 2 1 0 9 2
12 3 13 10 9 2 4 13 1 10 0 9 2
8 9 13 3 10 9 0 9 2
17 15 13 1 9 2 13 13 2 7 15 13 11 1 9 1 9 2
15 15 4 14 13 1 10 9 1 9 15 9 4 13 1 2
23 10 2 0 9 2 1 9 11 1 9 1 11 11 13 1 9 1 11 11 9 1 11 2
2 1 9
52 9 4 13 3 3 14 13 10 9 1 9 7 9 2 1 7 1 15 3 3 0 2 7 10 0 7 0 4 4 16 2 0 9 2 3 4 13 7 9 1 9 14 13 9 1 16 9 4 13 10 9 2
12 0 9 13 10 9 15 3 13 10 0 9 2
9 10 9 13 3 1 9 1 9 2
11 9 13 1 10 9 3 15 13 10 9 2
8 3 9 0 13 15 1 9 2
12 15 4 4 0 1 9 1 0 9 14 13 2
15 2 0 9 2 13 15 1 10 0 9 1 10 0 9 2
15 9 2 15 3 13 1 10 9 1 0 9 2 13 9 2
6 0 9 2 0 9 2
6 12 9 2 0 9 2
11 1 2 0 9 2 13 12 9 2 9 2
3 9 13 2
3 9 13 2
3 9 13 2
3 9 13 2
19 15 4 0 1 3 12 9 2 9 2 9 2 9 2 9 2 9 3 2
21 1 9 9 1 11 13 3 12 9 2 0 1 9 1 9 1 9 1 10 9 2
16 9 1 0 9 4 13 1 10 0 9 3 9 1 9 13 2
13 0 9 4 13 1 3 3 0 9 1 11 9 2
3 9 7 9
10 10 0 2 0 9 13 4 4 0 2
23 15 13 1 10 9 2 3 15 4 13 10 9 2 1 10 9 3 15 4 13 10 9 2
9 15 13 0 9 9 14 13 1 2
30 15 13 9 1 16 15 4 4 13 1 0 9 2 4 13 9 2 9 2 9 3 7 16 15 4 4 13 1 9 2
18 1 10 0 9 13 9 9 2 16 9 4 13 9 2 9 7 9 2
5 15 13 3 3 2
9 7 1 10 0 9 13 15 0 2
12 3 13 15 9 15 13 3 3 0 15 13 2
3 10 9 2
9 0 9 1 0 9 7 12 9 2
22 15 13 3 0 16 15 4 13 3 9 3 13 1 9 7 3 13 15 3 1 9 2
10 15 4 4 10 3 0 9 1 9 2
3 9 7 9
9 13 15 0 2 0 7 0 9 2
5 15 13 14 13 2
23 0 4 14 13 16 15 3 4 0 1 9 2 13 9 7 16 15 3 13 1 0 9 2
10 13 15 3 3 9 7 9 13 3 2
24 13 15 0 1 9 3 1 15 4 13 7 12 2 12 9 3 2 15 13 3 0 14 13 2
13 16 15 4 3 13 0 9 1 0 9 1 9 2
31 0 9 4 0 9 2 7 1 0 9 1 9 15 3 13 10 1 11 0 9 4 0 9 3 14 13 3 3 0 9 2
1 0
20 15 13 3 3 9 1 0 9 7 10 0 9 15 13 9 1 10 0 9 2
29 9 15 3 4 13 13 10 3 0 9 2 3 0 2 0 9 7 15 15 3 4 13 1 9 1 0 0 9 2
8 9 4 0 7 0 14 13 2
8 2 0 9 2 4 13 9 2
12 0 9 13 9 1 9 3 7 1 9 3 2
10 3 13 10 0 9 10 0 0 9 2
8 10 0 7 0 4 13 15 2
11 1 9 9 13 11 3 10 9 1 9 2
25 4 15 13 9 1 10 9 13 15 1 9 3 2 7 15 4 3 13 15 1 10 12 0 9 2
20 9 13 1 16 15 13 1 15 1 9 2 0 9 7 0 9 2 0 9 2
15 9 1 9 3 3 4 4 13 7 13 1 9 1 9 2
12 15 4 13 16 15 4 0 1 9 1 9 2
14 15 4 4 13 3 0 1 10 9 15 3 13 1 2
24 3 4 9 4 13 3 7 9 2 15 4 4 13 15 1 9 1 9 1 14 13 3 9 2
16 7 10 0 9 4 4 13 3 9 7 9 4 0 1 9 2
14 7 9 13 1 0 9 7 15 4 13 1 0 9 2
11 0 9 2 12 2 13 9 3 1 9 2
15 3 13 15 3 0 1 15 9 7 1 10 3 0 9 2
6 15 13 13 3 9 2
10 9 13 0 2 0 7 0 7 3 2
9 1 0 9 13 15 3 0 9 2
15 7 3 15 13 3 1 9 13 15 12 0 9 1 9 2
14 1 9 13 15 3 12 9 0 7 9 1 10 9 2
6 15 13 3 1 9 2
15 15 13 10 0 9 1 15 1 9 2 10 3 0 9 2
9 9 13 2 10 9 13 1 9 2
20 3 13 9 1 10 0 9 2 15 13 15 12 7 12 1 10 9 1 9 2
22 9 1 9 2 12 9 1 9 1 10 9 1 9 2 9 13 1 9 3 1 9 2
16 9 13 1 9 1 9 7 13 3 3 1 9 1 0 9 2
10 15 4 9 9 0 7 0 1 9 2
35 2 14 13 7 13 12 9 9 13 9 12 9 9 0 9 2 10 0 9 13 3 0 2 13 9 11 11 1 0 9 7 9 2 11 2
9 2 1 0 9 13 3 12 9 2
12 7 12 9 2 12 9 1 10 9 7 9 2
11 9 7 9 4 14 13 3 12 9 9 2
10 3 13 9 3 0 7 10 0 0 2
11 1 15 3 16 15 4 13 1 0 9 2
8 7 9 1 9 13 3 0 2
14 7 9 7 9 4 3 14 13 3 1 12 0 9 2
6 15 4 13 1 15 2
13 1 12 9 4 9 13 3 9 1 9 7 9 2
19 7 10 0 1 10 9 4 3 3 9 1 9 1 9 7 10 0 9 2
25 7 10 0 9 1 10 0 9 4 16 9 1 9 4 14 4 1 12 9 0 16 9 4 0 2
11 9 12 13 15 10 0 0 9 7 9 2
26 15 4 1 10 9 14 13 15 3 0 9 3 10 9 13 1 10 9 9 1 9 2 9 7 9 2
30 9 4 10 0 0 9 2 15 13 3 9 7 13 14 13 3 9 15 13 12 9 2 15 4 3 13 12 1 10 2
26 1 9 15 13 9 1 9 13 15 3 12 9 2 3 16 15 13 9 1 10 9 3 3 1 9 2
8 10 9 13 1 9 1 9 2
41 3 9 13 1 9 7 9 4 0 13 9 2 15 15 7 15 4 13 12 9 2 3 0 7 9 1 0 9 2 1 9 1 0 9 2 10 9 1 0 9 2
12 3 13 9 2 9 1 9 2 9 7 9 2
13 16 9 4 13 3 1 9 2 13 15 3 3 2
6 3 13 15 0 9 2
21 16 9 13 3 1 9 1 9 4 15 13 3 10 9 9 1 16 9 4 0 2
7 1 9 4 3 9 0 2
14 2 3 9 7 9 4 14 13 12 2 13 11 11 2
10 7 3 13 15 9 3 3 1 9 2
15 2 3 13 9 2 15 4 0 7 13 3 14 3 13 2
15 15 4 13 16 9 13 2 16 10 0 3 13 1 9 2
14 3 13 15 7 3 9 1 9 1 9 1 10 0 2
13 2 7 10 9 4 3 14 13 3 3 7 3 2
20 12 9 9 13 3 7 10 0 9 2 7 1 10 9 0 3 3 1 9 2
20 9 13 3 1 9 0 9 1 9 2 7 3 4 9 13 3 1 12 9 2
7 15 4 0 9 1 3 2
54 7 1 9 1 15 3 12 9 4 13 1 9 7 9 4 15 0 14 13 3 9 1 12 9 0 9 2 0 1 9 9 2 11 12 2 7 0 3 10 9 15 3 13 2 3 4 13 1 9 1 12 9 9 2
28 11 11 15 4 9 1 10 9 7 1 12 9 3 4 9 1 9 1 11 4 0 9 14 13 1 10 9 2
7 2 15 4 0 0 9 2
24 9 4 1 0 9 1 10 9 2 9 1 10 9 15 4 13 0 9 13 1 9 1 9 2
43 15 13 3 1 9 1 9 1 12 9 1 9 1 9 2 1 9 1 0 0 9 2 3 9 13 1 9 16 15 3 3 4 13 9 1 9 1 3 0 9 1 9 2
7 3 13 9 12 10 9 2
29 10 0 9 9 13 3 2 0 9 2 0 9 1 0 2 9 1 9 2 9 1 9 3 12 2 12 2 3 2
17 7 9 2 9 7 9 2 0 9 1 0 9 2 15 4 13 2
7 15 13 10 3 0 9 2
14 9 13 14 13 3 9 7 13 1 10 3 0 9 2
10 3 13 14 13 16 15 13 0 9 2
31 15 13 12 9 2 12 9 1 0 9 2 1 1 9 14 13 3 0 9 7 13 10 3 0 0 9 1 10 0 9 2
23 15 9 3 13 1 9 3 13 10 9 16 15 4 0 14 13 9 9 3 3 1 9 2
18 3 1 9 1 9 1 10 0 9 2 13 15 3 3 3 9 13 2
20 3 10 3 9 2 3 10 3 9 1 11 13 3 2 4 15 13 9 3 2
20 10 12 0 9 2 1 9 7 9 2 4 3 3 13 3 1 9 2 9 2
25 15 13 10 3 12 9 2 1 3 10 3 0 9 7 3 2 15 13 9 7 9 1 0 9 2
19 15 13 10 9 1 9 15 9 7 9 4 0 1 2 1 10 0 9 2
32 9 13 10 12 9 7 13 3 0 9 1 10 0 9 2 16 12 9 4 13 3 1 10 0 9 0 1 10 0 9 12 2
25 9 7 11 11 4 9 2 9 2 1 10 9 1 9 1 3 12 9 7 1 0 9 1 9 2
17 7 9 9 4 3 9 9 2 10 9 2 10 0 3 1 9 2
26 9 1 16 15 13 0 0 7 9 1 9 13 1 16 3 12 2 3 12 9 13 1 0 0 9 2
18 11 11 13 10 3 0 9 1 9 7 11 11 2 7 9 4 0 2
9 9 13 3 7 13 3 12 9 2
6 15 13 3 1 9 2
9 10 9 1 9 4 3 9 13 2
21 15 13 10 9 9 1 11 2 10 0 11 9 1 9 2 15 13 10 0 9 2
13 3 13 15 1 16 10 9 9 13 0 1 9 2
27 7 3 4 3 9 13 3 3 1 12 9 16 9 15 12 13 1 3 12 9 1 9 13 1 12 9 2
8 9 4 3 3 0 7 9 2
19 15 13 3 3 15 15 4 13 10 0 12 9 1 9 7 11 7 11 2
14 7 15 13 0 9 1 9 15 13 3 3 1 9 2
14 10 12 9 4 9 4 3 0 2 10 12 9 9 2
13 9 7 9 4 3 13 1 9 1 9 7 9 2
9 7 0 9 4 3 13 1 9 2
28 0 9 1 10 9 7 11 2 0 1 9 2 13 16 10 0 9 13 3 12 9 3 1 9 7 1 9 2
12 2 3 12 1 9 2 3 12 1 9 2 2
17 13 15 0 9 1 10 0 9 7 10 9 7 1 11 2 11 2
12 0 9 13 1 0 9 2 7 3 3 3 2
4 3 1 9 2
19 11 7 2 11 2 4 13 3 10 0 9 9 15 15 2 13 2 12 2
11 7 10 0 9 4 3 13 1 10 0 2
14 3 10 9 13 2 13 10 9 1 9 9 14 13 2
8 3 3 10 0 9 3 13 2
6 3 3 13 15 12 2
15 1 9 1 9 13 15 10 9 7 13 9 1 9 1 2
11 3 13 15 3 1 9 1 9 7 9 2
23 1 12 0 0 9 2 15 1 9 3 13 3 1 1 9 2 13 3 9 3 1 9 2
12 9 2 1 9 2 4 10 9 1 0 9 2
15 10 12 9 1 9 13 9 2 10 12 0 9 3 9 2
12 15 15 13 9 4 13 9 1 9 1 9 2
6 1 9 9 13 9 2
11 1 9 1 9 13 9 3 9 1 9 2
16 9 13 3 2 13 3 7 13 3 3 1 9 1 0 9 2
15 1 9 9 13 9 1 0 9 2 15 13 9 1 9 2
3 12 9 9
3 12 9 9
3 9 13 9
2 0 9
3 10 9 2
11 3 2 7 9 4 0 1 10 0 9 2
10 1 9 13 11 9 1 3 12 9 2
20 9 1 9 13 10 9 1 12 9 2 15 4 13 12 9 9 1 9 12 2
2 9 13
15 1 9 13 15 1 16 9 4 13 3 2 1 12 9 2
17 1 9 13 15 12 9 3 12 9 2 12 13 15 3 12 9 2
12 10 0 0 9 15 13 3 4 9 12 9 2
17 12 4 15 14 13 3 12 9 9 2 1 3 12 9 1 9 2
17 1 10 3 0 9 12 4 9 14 13 3 0 2 3 12 9 2
10 12 13 15 12 9 9 1 10 9 2
2 0 9
20 1 9 4 9 7 9 9 14 13 1 3 12 9 2 9 13 1 12 9 2
14 3 10 9 1 10 0 7 0 4 14 13 10 9 2
3 9 1 9
11 9 4 3 14 13 3 3 7 1 9 2
25 1 10 0 12 9 1 9 2 4 9 2 15 13 1 9 2 13 1 10 0 9 1 12 9 2
10 0 9 4 14 13 1 10 0 9 2
12 9 4 14 13 1 9 2 9 2 0 9 2
18 3 4 3 10 0 9 9 1 9 7 9 14 13 0 7 14 13 2
2 0 9
11 7 1 0 9 3 13 15 9 1 9 2
15 1 12 7 12 9 1 9 13 9 1 9 3 1 12 2
14 10 9 13 15 4 14 13 1 9 2 9 7 9 2
3 15 13 3
24 9 9 2 12 9 2 4 14 13 1 10 0 12 9 2 7 15 13 0 1 9 1 9 2
14 9 13 10 9 2 1 9 0 4 15 14 13 3 2
3 0 1 9
13 9 9 1 0 9 4 14 13 0 9 1 9 2
17 1 9 13 9 9 1 10 0 1 12 9 12 1 12 9 3 2
10 12 13 12 9 1 10 0 1 9 2
6 12 4 9 12 9 2
17 10 9 13 9 1 9 1 10 0 9 1 9 1 10 0 9 2
2 9 9
24 9 4 14 13 9 2 10 0 9 13 7 13 3 10 9 1 0 9 1 7 9 7 9 2
20 15 13 0 14 13 9 1 9 9 2 15 13 3 0 14 13 9 1 9 2
15 9 4 13 0 9 1 0 9 7 13 15 1 0 9 2
18 9 4 14 13 0 9 1 10 9 2 10 9 1 7 0 7 0 2
13 3 4 10 9 13 9 3 10 9 13 1 9 2
4 10 0 9 2
15 9 1 10 9 4 0 1 9 7 9 15 13 1 3 2
18 9 13 3 0 0 9 1 14 13 0 9 0 1 0 9 1 9 2
21 7 3 13 15 10 0 9 15 13 10 0 3 15 13 16 15 13 3 1 9 2
16 15 13 16 15 4 13 15 1 10 9 15 10 9 4 0 2
10 9 13 16 10 9 13 3 1 9 2
6 15 4 10 0 9 2
13 3 13 15 13 1 10 0 9 7 15 13 3 2
22 0 9 2 2 9 2 2 0 9 2 2 0 9 7 2 9 15 3 4 13 3 2
12 7 9 9 4 13 13 1 7 9 7 9 2
2 13 3
18 9 11 11 2 11 2 4 1 10 0 9 13 9 1 12 0 9 2
26 9 2 15 4 13 10 9 3 3 2 9 15 13 10 9 9 12 7 10 9 15 13 12 9 3 2
24 15 13 15 4 10 9 1 9 14 3 1 9 1 10 9 13 10 9 1 10 9 1 9 2
22 7 15 13 16 15 3 1 9 4 13 1 9 1 3 0 9 7 3 13 0 9 2
16 15 4 13 1 10 9 9 14 13 9 1 3 9 13 3 2
31 15 13 15 0 16 10 0 9 15 13 13 9 12 7 15 4 13 3 3 10 9 3 1 14 13 1 9 3 4 0 2
14 2 15 13 3 2 10 9 4 0 7 10 9 0 2
31 13 15 0 9 4 15 13 3 7 13 3 7 3 4 15 1 9 16 15 13 10 9 2 3 1 9 2 14 13 9 2
16 9 13 0 1 9 1 10 9 15 4 13 2 13 9 11 2
2 0 9
15 2 9 15 3 13 3 3 4 3 3 13 10 9 0 2
20 1 10 0 9 13 15 3 1 9 7 13 3 3 1 0 9 2 3 9 2
31 1 9 7 9 3 15 4 0 4 15 13 1 14 13 10 2 9 2 7 3 3 3 4 15 7 2 9 2 13 9 2
36 0 9 13 16 15 15 4 0 1 9 13 10 0 9 3 2 16 15 15 13 9 7 10 0 9 2 3 1 9 2 13 0 9 1 9 2
18 9 4 7 0 3 10 0 9 4 7 0 1 9 2 13 11 9 2
21 10 0 13 10 9 3 7 1 15 13 10 9 3 3 1 9 7 3 1 9 2
26 2 13 7 9 10 0 9 3 10 9 15 4 10 0 9 7 13 14 13 13 3 13 1 10 9 2
17 15 4 13 3 3 1 0 9 7 15 13 3 10 9 15 13 2
25 15 13 15 0 16 9 3 13 10 9 1 14 13 3 1 3 10 9 13 15 13 3 1 9 2
4 10 9 9 2
23 3 13 0 16 15 15 4 13 13 3 3 4 13 1 9 3 2 3 4 10 9 13 2
7 7 3 0 4 3 9 2
31 15 4 0 14 13 10 0 9 2 15 4 10 0 9 7 10 0 15 13 4 16 7 0 15 13 2 3 0 13 9 2
23 15 4 3 9 1 10 9 15 4 13 1 0 9 2 3 12 9 9 2 12 9 9 2
23 9 4 13 0 9 1 16 10 0 9 13 10 0 9 7 15 4 10 9 15 4 13 2
9 13 15 10 9 1 9 7 9 2
13 9 11 4 13 16 9 13 0 14 13 1 9 2
7 10 9 9 4 3 0 2
9 3 4 10 0 0 3 15 13 2
13 3 2 15 15 4 13 10 0 9 3 4 9 2
22 15 15 13 9 1 10 0 9 4 9 15 1 9 1 10 3 0 9 13 3 3 2
3 2 9 2
39 11 4 3 1 10 9 13 3 9 1 0 7 0 9 2 3 4 9 13 7 3 4 15 1 10 9 9 4 13 9 0 14 13 10 9 1 10 9 2
13 10 12 9 13 0 3 9 1 0 2 0 9 2
8 9 1 9 7 9 4 0 2
5 10 0 4 0 2
21 1 9 15 13 3 2 0 2 9 13 10 9 1 0 9 2 2 9 2 2 2
18 9 4 3 3 15 13 9 7 9 13 3 10 9 7 13 3 9 2
13 1 9 4 15 13 1 9 2 1 9 1 9 2
14 7 10 1 9 0 9 4 13 14 13 9 1 9 2
3 13 9 2
25 1 11 4 3 9 3 15 13 9 13 3 7 1 11 13 15 9 15 13 3 9 1 0 9 2
34 2 3 4 9 13 15 2 7 15 4 3 0 14 13 10 0 9 15 10 9 13 7 13 14 13 10 9 15 4 0 10 0 9 2
34 14 13 0 9 2 0 9 2 0 9 4 13 1 7 9 7 10 0 9 2 13 9 11 2 15 13 9 0 9 1 1 12 9 2
12 4 15 3 13 9 1 9 1 9 0 9 2
20 11 11 2 0 9 1 11 2 4 13 10 9 1 9 1 12 0 9 9 2
13 9 1 9 13 1 3 12 9 1 12 1 12 2
23 7 1 9 7 9 4 15 0 1 9 7 13 2 15 1 10 9 2 14 13 9 3 2
38 16 15 4 10 0 9 13 10 0 9 1 0 9 3 9 11 11 1 11 3 2 1 9 1 0 9 1 9 2 13 15 1 9 1 2 9 2 2
7 1 9 13 9 1 9 2
7 9 13 1 10 0 9 2
25 9 1 9 13 3 1 12 9 7 4 3 13 1 12 9 7 1 0 9 1 9 3 3 3 2
22 1 9 1 11 12 9 13 9 1 11 9 11 11 16 9 1 9 13 1 10 9 2
10 2 15 13 1 14 13 3 3 2 2
26 9 11 11 11 4 13 10 9 1 9 2 10 9 1 15 15 13 10 0 9 2 1 14 13 9 2
21 9 1 11 11 11 1 11 2 11 2 4 1 10 9 13 10 0 2 9 2 2
12 9 1 9 4 1 0 9 0 2 13 15 2
9 0 9 4 13 1 10 0 9 2
25 16 3 9 9 13 1 12 1 12 9 1 9 3 4 15 0 1 10 9 1 12 9 1 9 2
20 10 9 1 10 0 9 1 10 9 1 9 13 10 9 1 12 9 1 9 2
12 15 4 0 14 13 15 15 3 13 1 9 2
26 10 9 13 9 1 10 0 9 2 7 1 9 1 10 9 15 13 13 15 10 0 9 1 10 9 2
4 1 12 1 12
21 9 10 9 1 9 2 1 12 10 9 1 9 2 13 10 0 9 1 9 0 2
17 9 4 13 1 12 1 10 12 9 12 1 12 1 0 9 12 2
12 3 1 12 4 9 0 7 10 12 0 9 2
18 9 1 9 7 9 1 9 1 9 13 3 9 2 1 0 9 2 2
25 13 15 9 1 9 2 9 2 9 7 9 13 15 10 0 9 1 9 1 3 3 12 9 12 2
11 3 13 3 3 10 0 9 3 1 9 2
6 9 3 12 9 1 12
13 10 0 9 4 9 9 1 0 2 10 3 9 2
19 9 1 12 9 12 9 12 13 3 9 1 16 15 13 9 1 0 9 2
21 1 12 4 9 13 3 1 12 9 2 15 4 1 9 1 15 15 13 1 9 2
12 0 9 12 13 10 9 9 0 9 7 9 2
16 7 9 13 9 7 9 1 9 1 0 9 2 9 7 9 2
24 10 9 7 0 9 1 12 9 2 12 9 9 2 13 3 0 9 1 9 9 1 0 12 2
10 11 9 12 9 12 9 9 12 9 12
25 12 9 1 9 7 9 2 3 3 7 3 12 9 1 9 2 4 10 9 15 4 0 14 13 2
13 9 9 4 1 11 13 1 9 2 3 1 11 2
14 1 11 13 0 9 1 9 1 12 0 9 1 11 2
15 9 13 9 1 0 9 2 12 12 12 12 12 12 12 12
4 0 9 1 11
17 1 9 9 2 9 0 9 2 4 9 13 3 12 9 1 9 2
27 15 13 3 0 3 2 7 16 15 13 10 9 1 15 4 15 10 9 3 2 13 9 11 11 1 11 2
31 1 9 1 0 9 4 9 0 1 9 2 1 12 7 12 13 9 1 12 1 12 9 1 9 2 7 15 13 0 9 2
10 9 4 1 15 3 0 7 12 9 2
17 9 11 13 16 9 9 7 9 9 1 9 3 4 13 1 9 2
25 11 4 10 0 9 2 3 13 15 1 12 9 10 0 9 15 9 11 3 13 7 3 13 1 2
15 15 15 13 0 9 10 0 9 13 12 9 3 1 9 2
6 9 13 3 1 9 2
12 1 9 13 15 3 16 15 13 10 0 9 2
5 13 12 9 10 9
18 15 13 1 12 9 9 7 12 3 0 9 1 16 9 4 13 3 2
10 9 4 13 13 16 15 3 13 9 2
10 10 0 9 13 10 9 1 12 9 2
13 1 12 7 12 9 1 9 13 13 15 1 9 2
11 1 11 13 9 13 3 12 9 1 9 2
27 1 9 9 13 15 16 9 1 9 13 1 3 12 9 2 15 13 0 10 9 1 12 2 3 9 13 2
5 9 11 11 13 2
10 2 15 13 3 16 9 13 10 9 2
9 9 4 13 1 10 3 0 9 2
9 9 1 9 1 0 9 4 13 2
14 15 13 1 9 3 9 1 12 9 9 1 0 9 2
4 9 13 12 2
15 15 13 3 3 0 14 13 3 9 1 12 2 1 9 2
13 7 1 11 13 10 9 9 0 1 9 1 9 2
18 15 4 2 3 2 9 1 10 9 15 13 1 10 0 9 0 9 2
19 10 9 3 0 16 9 13 0 1 10 9 1 9 1 12 1 9 9 2
29 10 12 4 2 9 2 0 1 9 11 1 11 2 9 0 9 9 11 11 2 9 2 7 2 9 2 11 11 2
5 9 1 9 13 2
30 4 15 13 14 13 0 9 3 3 15 4 0 16 10 0 9 9 15 3 13 1 15 4 13 0 9 2 9 2 2
11 2 6 2 13 11 11 1 9 0 9 2
7 3 13 7 13 1 9 2
11 2 6 2 13 11 11 1 9 1 9 2
39 14 13 3 7 3 13 9 9 1 9 4 3 0 16 15 4 0 14 13 15 1 9 1 10 0 0 9 15 4 13 1 15 1 10 1 9 0 9 2
21 1 9 2 9 11 11 1 11 2 4 13 16 15 4 0 7 4 13 0 9 2
11 4 15 13 3 7 13 13 9 1 9 2
22 4 15 3 13 15 1 14 13 9 1 14 13 1 9 1 9 2 9 7 0 9 2
15 9 2 9 2 9 2 13 3 0 9 1 10 0 9 2
10 4 15 3 13 13 1 9 1 11 2
17 9 4 3 0 1 10 9 7 9 15 9 1 9 4 13 1 2
13 13 15 16 15 4 0 9 11 11 2 9 2 2
36 6 2 7 9 11 7 9 11 13 16 15 3 13 0 9 14 13 13 10 0 9 2 15 13 12 9 1 10 0 0 9 1 3 12 9 2
7 0 9 13 10 0 9 2
7 9 4 13 3 0 9 2
10 10 9 13 14 13 10 3 0 9 2
17 9 13 3 3 1 2 7 1 9 2 1 9 7 1 0 9 2
3 2 9 2
18 1 0 9 1 12 9 13 15 0 9 3 1 12 9 2 13 11 2
12 7 9 4 13 16 9 13 3 1 12 9 2
13 3 4 15 3 3 0 1 0 7 1 0 9 2
14 9 1 9 13 9 1 9 3 3 7 10 0 9 2
9 7 9 4 0 2 9 3 0 2
16 1 9 13 3 3 1 9 2 15 3 4 0 3 7 9 2
2 10 9
16 3 4 15 3 13 3 1 10 9 15 13 1 12 9 3 2
14 3 13 9 15 1 15 1 9 2 9 2 3 9 2
7 15 13 0 9 1 9 2
10 7 3 13 15 3 1 9 1 9 2
13 15 13 9 1 9 7 10 9 1 0 0 9 2
9 10 0 9 13 9 1 10 9 2
9 13 9 1 9 1 13 3 3 2
4 3 1 9 2
12 3 13 9 1 9 1 7 9 13 1 9 2
7 1 9 9 4 15 0 2
13 9 4 1 9 13 9 9 1 9 7 1 9 2
12 10 0 9 4 10 12 9 13 1 1 9 2
11 3 9 0 1 9 1 4 13 0 9 2
17 9 7 9 4 10 9 2 9 15 13 3 1 9 4 10 0 2
12 9 1 9 4 3 0 1 14 13 0 9 2
11 7 9 1 9 4 13 2 13 9 11 2
12 9 7 10 9 15 13 4 3 0 1 9 2
17 15 4 3 3 0 14 13 3 15 1 9 2 9 7 0 9 2
5 9 13 3 3 2
19 15 13 3 10 0 9 1 10 9 15 13 9 2 7 15 13 3 9 2
3 9 13 2
1 9
12 1 0 9 13 10 12 9 9 9 1 9 2
6 3 3 15 13 9 2
26 4 9 13 10 9 3 16 15 3 13 3 9 3 15 13 16 0 2 3 9 9 2 4 14 13 2
8 15 4 13 2 13 11 11 2
13 9 4 13 1 16 15 13 3 9 1 0 9 2
25 11 11 1 10 9 13 9 1 3 0 9 2 1 9 2 9 2 1 9 4 13 0 1 9 2
17 3 16 15 13 1 0 9 1 9 7 2 13 3 2 10 9 2
8 3 3 13 1 10 0 9 2
4 11 11 2 9
4 11 11 2 9
8 3 0 13 9 1 9 9 2
18 10 9 13 15 15 1 9 2 16 9 9 13 13 10 9 1 9 2
15 1 11 13 9 1 12 9 1 0 9 1 12 9 3 2
15 3 11 13 9 13 9 1 0 12 9 1 9 0 9 2
12 10 9 9 1 10 0 9 9 13 1 9 2
32 10 9 9 14 13 0 9 13 1 10 9 15 13 1 10 9 1 9 1 9 9 14 13 9 1 11 1 10 12 9 12 2
26 1 9 13 3 10 9 15 4 13 1 9 1 14 13 3 0 9 1 9 3 15 4 0 1 9 2
26 3 10 9 1 12 0 9 1 9 13 1 9 2 15 9 4 13 1 10 9 9 16 15 13 15 2
26 9 4 1 9 14 13 9 12 7 13 15 3 10 0 9 3 3 1 9 13 1 1 9 1 9 2
9 10 0 4 3 13 10 0 9 2
1 9
14 15 4 3 13 1 10 9 9 2 3 15 13 9 2
9 1 11 13 9 3 3 7 12 2
8 9 13 1 9 1 12 9 2
17 9 1 9 1 0 9 1 11 13 9 0 1 1 9 12 9 2
28 0 9 2 9 2 13 9 2 3 10 0 9 2 10 0 2 13 9 0 1 12 1 12 9 9 1 9 2
16 10 0 9 1 11 13 1 12 9 9 1 10 9 1 9 2
21 0 9 13 1 9 1 14 13 9 7 13 9 1 9 1 9 2 9 7 9 2
18 10 0 2 0 2 9 4 4 13 3 3 1 10 9 1 12 9 2
1 9
9 0 9 13 3 3 9 1 9 2
13 9 1 9 4 13 3 1 12 9 1 10 9 2
16 12 9 1 9 4 13 1 9 7 9 4 9 13 9 1 2
12 7 9 7 9 13 0 1 9 1 9 9 2
13 9 3 16 15 13 1 16 9 1 9 4 13 2
22 9 4 0 3 16 10 0 9 1 10 0 9 3 13 10 9 1 9 1 10 0 2
4 0 12 9 9
17 10 9 13 9 3 10 0 9 12 13 14 3 13 10 0 9 2
11 9 13 1 0 12 9 1 9 0 9 2
20 10 9 13 1 9 9 14 13 9 1 10 0 9 1 10 0 9 1 11 2
31 10 3 0 9 1 3 12 9 0 12 13 3 12 9 1 9 7 15 4 3 0 7 9 1 15 10 9 13 1 9 2
29 9 4 13 3 0 9 14 13 10 0 0 9 1 16 9 13 1 10 3 0 9 0 9 0 1 9 7 9 2
40 9 4 13 1 10 0 9 1 0 9 1 9 1 3 10 9 3 10 0 0 9 13 3 9 4 13 0 1 9 15 4 13 3 1 9 2 9 7 9 2
2 0 9
20 7 3 7 1 10 0 9 4 9 3 0 16 15 4 13 3 3 7 3 2
20 10 0 15 3 13 9 1 9 1 0 9 13 3 3 3 1 16 9 13 2
25 10 9 15 4 0 3 14 13 1 9 1 9 4 13 1 0 7 3 1 9 0 9 1 9 2
15 9 1 11 0 9 4 13 16 9 9 14 13 4 13 2
27 9 13 1 9 7 9 2 10 9 15 13 13 0 3 1 11 2 15 15 11 4 13 3 10 3 9 2
12 7 3 13 9 3 0 2 3 13 3 9 2
10 10 9 15 13 9 13 3 0 9 2
10 3 12 9 1 9 13 1 0 9 2
20 9 15 13 3 1 9 13 3 10 3 9 9 2 10 0 9 0 1 9 2
16 10 0 2 3 9 2 13 1 0 0 9 1 10 0 9 2
17 0 9 4 13 1 9 1 10 0 9 7 13 0 2 0 9 2
24 1 9 9 7 9 2 2 2 4 15 3 13 3 9 7 13 15 1 15 1 11 9 0 2
15 2 15 4 9 9 14 13 1 16 9 13 0 1 9 2
17 13 15 15 3 15 13 10 0 9 15 4 10 9 1 0 9 2
13 3 13 9 3 0 3 1 10 9 15 13 9 2
22 10 9 1 9 11 11 1 11 13 10 0 9 1 9 9 15 13 1 11 1 9 2
20 9 11 11 1 9 7 9 11 11 13 1 9 1 10 0 0 9 1 9 2
18 3 4 9 1 10 0 9 4 0 3 7 10 9 2 13 11 11 2
10 7 10 9 4 3 13 10 0 9 2
13 1 10 0 9 4 10 3 9 13 9 0 9 2
25 15 13 10 0 9 1 9 1 10 10 9 15 13 15 1 10 9 1 0 9 2 13 11 11 2
10 3 0 9 13 15 3 3 3 3 2
23 3 13 10 9 9 1 10 9 15 9 11 3 1 0 9 13 15 0 16 15 4 13 2
2 9 13
15 9 1 15 13 15 2 0 9 1 9 2 9 7 9 2
13 9 1 0 9 4 3 3 0 7 9 1 9 2
13 3 13 15 15 13 1 9 16 9 13 14 13 2
15 1 11 9 13 9 1 12 9 1 9 12 1 9 12 2
12 1 10 9 13 9 1 9 1 11 1 9 2
7 15 7 3 13 1 9 2
9 1 10 9 4 10 0 9 13 2
10 3 12 9 7 0 9 13 0 9 2
19 15 4 3 3 15 7 3 7 15 4 15 16 9 13 1 0 10 9 2
35 3 0 7 0 4 9 1 9 7 9 1 9 16 9 2 9 2 9 7 0 15 13 9 11 11 7 11 11 7 13 14 4 13 1 2
7 3 13 3 9 7 9 2
9 9 11 11 13 13 1 10 9 2
8 9 4 3 3 10 0 9 2
4 9 4 0 2
15 9 1 9 7 1 9 13 0 9 7 9 3 1 9 2
7 0 9 4 4 10 9 2
7 9 13 3 1 0 9 2
22 10 9 13 3 3 0 9 7 13 1 14 3 13 1 9 7 13 1 3 0 9 2
9 9 13 10 9 2 13 11 11 2
21 15 4 13 10 0 1 9 2 13 15 3 16 9 13 15 0 14 13 1 9 2
13 3 4 10 9 13 3 2 13 10 9 1 9 2
10 1 10 0 9 1 9 3 13 9 2
16 15 13 3 3 1 9 7 15 13 0 9 14 13 0 9 2
17 10 9 13 3 3 1 9 1 9 2 13 9 11 11 1 11 2
25 9 11 13 2 16 9 1 10 0 9 3 1 12 2 12 9 4 4 0 1 10 9 1 9 2
3 3 13 9
23 3 13 3 9 9 1 9 9 2 3 15 3 13 10 0 9 7 3 9 1 10 9 2
20 9 13 10 9 7 13 1 0 9 1 14 13 0 9 7 0 9 1 9 2
8 13 15 13 10 9 1 9 2
17 13 9 1 9 3 12 9 2 10 1 0 7 10 1 0 9 2
18 13 9 1 9 2 9 7 10 9 3 10 0 9 7 13 1 9 2
11 15 4 13 1 0 9 1 10 9 9 2
21 1 0 9 1 11 9 4 15 13 13 10 9 1 9 9 1 0 9 7 9 2
27 1 10 3 0 9 9 7 9 13 10 9 1 9 1 12 0 2 9 13 3 7 3 13 10 9 3 2
16 15 13 15 16 9 13 10 3 0 9 1 3 15 1 9 2
14 15 4 3 13 16 9 13 10 0 9 3 1 9 2
24 1 10 3 12 9 1 9 12 9 4 12 9 3 13 1 9 16 15 13 2 0 9 2 2
13 1 10 12 0 9 1 10 9 4 12 3 13 2
42 1 0 9 13 15 16 9 1 9 2 12 9 2 10 9 2 4 10 2 3 0 2 9 2 16 9 1 9 4 9 2 7 16 9 4 13 1 10 0 0 9 2
17 10 0 9 1 9 13 9 1 9 9 16 10 0 9 13 3 2
25 9 4 3 3 13 9 1 16 9 1 11 4 13 9 1 9 2 9 2 9 7 9 1 9 2
22 9 4 13 10 0 9 9 0 0 9 7 13 15 1 10 9 1 10 0 12 9 2
30 1 9 4 9 13 9 1 14 4 13 3 3 3 1 9 7 12 9 1 9 2 13 9 15 13 9 2 11 11 2
19 1 9 9 0 12 1 9 13 0 9 11 11 3 11 9 1 11 9 2
19 15 13 9 1 3 10 0 9 0 9 1 9 1 10 0 9 11 11 2
24 2 10 3 9 4 15 13 1 11 1 2 13 9 11 1 0 9 11 11 1 9 1 9 2
5 11 13 3 3 2
1 9
1 9
2 0 9
1 9
12 11 13 16 11 13 9 1 9 1 11 0 2
18 10 0 9 4 0 1 10 0 0 9 1 9 1 10 0 0 9 2
3 9 1 11
9 7 9 4 11 9 1 11 9 2
14 7 15 4 3 13 10 0 9 3 1 3 10 9 2
21 3 1 9 2 9 0 9 13 15 9 11 11 15 1 11 9 13 10 0 9 2
9 15 13 10 1 9 3 0 9 2
8 9 15 13 1 11 13 1 2
7 9 11 11 2 12 9 2
10 0 9 1 11 11 11 2 12 9 2
6 9 11 11 2 9 2
15 10 9 13 14 13 3 0 9 1 9 1 10 0 9 2
16 3 9 0 9 4 0 4 9 13 10 9 1 9 1 9 2
13 15 13 3 11 13 9 1 10 0 9 1 11 2
4 2 9 1 9
13 2 15 4 1 9 13 15 15 1 0 9 13 2
12 15 4 10 0 9 9 1 11 9 1 9 2
9 9 13 3 1 11 9 1 9 2
24 3 13 15 9 0 9 11 11 15 13 9 1 9 1 10 12 0 9 11 2 11 7 11 2
9 2 15 4 13 10 9 1 9 2
15 15 13 15 15 15 13 0 9 1 2 13 10 0 9 2
25 15 13 16 10 0 9 1 9 2 9 2 9 3 3 4 14 13 3 1 11 2 11 7 11 2
16 10 0 9 4 3 13 3 3 1 10 9 16 15 13 0 2
15 3 13 11 7 11 9 2 15 13 0 9 2 1 9 2
8 1 12 9 13 15 3 9 2
10 3 1 9 4 9 13 1 10 9 2
13 4 11 13 1 0 9 7 9 7 13 9 9 2
12 1 9 9 0 9 4 11 13 1 10 9 2
15 10 0 9 4 14 13 1 11 10 9 9 1 9 3 2
6 3 13 15 1 11 2
12 1 11 13 10 0 9 1 9 1 10 9 2
8 15 13 3 0 9 1 9 2
10 1 0 9 4 15 14 13 1 9 2
11 9 4 1 9 14 13 1 9 1 9 2
10 11 9 1 11 13 1 9 11 11 2
9 15 13 10 0 9 1 10 9 2
16 15 4 13 14 13 7 3 7 13 1 15 15 13 1 11 2
13 1 10 0 9 13 10 9 3 3 3 14 13 2
7 2 11 13 9 1 9 2
6 9 1 11 13 11 2
13 7 11 9 7 15 15 4 13 1 11 13 0 2
7 10 9 4 10 0 9 2
19 1 11 13 15 9 1 12 9 1 9 2 7 3 0 9 1 0 9 2
13 11 13 15 1 9 0 14 13 1 11 0 9 2
10 10 0 9 13 3 3 1 11 9 2
14 3 13 15 12 0 9 1 11 1 11 9 1 9 2
25 9 2 3 11 2 11 2 11 2 13 3 16 11 0 9 4 13 1 16 10 0 11 13 1 2
22 15 4 0 14 13 11 10 0 9 1 10 9 1 14 13 11 0 9 7 0 9 2
18 9 2 0 1 11 2 4 13 1 11 1 14 13 3 1 11 9 2
6 15 4 13 9 9 2
9 3 4 15 13 11 10 0 9 2
3 9 1 9
19 11 9 14 13 1 0 9 1 0 9 13 3 1 10 9 2 13 9 2
13 1 0 9 13 15 2 16 11 13 9 1 9 2
3 3 0 2
9 11 13 10 9 7 13 0 9 2
4 9 4 15 2
9 10 0 9 4 13 1 11 9 2
9 9 4 13 10 9 1 11 9 2
7 9 4 3 13 0 9 2
5 9 4 13 9 2
5 9 1 10 9 2
8 10 9 13 15 15 4 13 2
6 15 4 13 3 3 2
10 9 13 9 14 1 9 13 1 9 2
21 15 13 16 12 9 1 10 0 9 13 0 16 11 13 1 10 9 15 3 13 2
8 10 3 0 0 9 4 13 2
8 9 13 1 10 9 0 9 2
12 9 1 9 1 0 9 4 3 13 3 3 2
12 9 4 13 1 1 9 3 12 9 0 9 2
7 11 9 4 3 3 13 2
11 9 1 9 4 4 13 3 0 7 3 2
21 7 1 9 9 4 15 13 16 9 3 4 4 14 13 10 0 9 1 11 9 2
21 9 4 1 10 9 13 10 9 15 0 9 2 10 0 9 7 0 9 4 13 2
25 3 4 15 13 1 16 10 0 9 13 0 9 14 13 3 7 3 4 13 9 1 10 0 9 2
15 9 1 10 0 9 14 13 9 1 10 0 9 4 13 2
19 9 13 1 10 0 9 10 0 9 15 11 7 11 7 0 3 13 1 2
20 3 3 4 9 11 11 13 13 1 14 13 10 0 9 3 1 11 1 9 2
19 11 0 9 7 9 4 13 3 1 9 1 9 1 10 3 0 0 9 2
18 1 3 4 11 13 1 10 9 15 13 1 10 9 1 11 1 9 2
29 3 4 9 13 3 7 13 13 1 12 0 9 7 10 9 2 10 0 9 7 10 0 9 2 15 1 0 9 2
18 9 13 7 0 2 7 9 11 11 2 15 13 10 0 9 2 13 2
32 11 13 10 3 9 2 1 15 15 3 4 13 9 2 7 3 3 4 15 1 9 1 10 0 1 16 15 13 10 0 9 2
20 2 3 13 15 3 1 9 14 13 9 1 9 1 9 2 13 9 11 11 2
9 10 0 9 13 1 12 0 9 2
16 15 4 15 13 1 16 15 13 12 9 2 9 13 3 12 2
21 9 1 10 0 9 4 13 10 9 15 3 13 1 9 2 3 12 9 1 11 2
45 1 10 9 4 15 13 16 15 4 10 3 9 2 7 14 13 1 9 1 9 1 9 4 15 13 16 15 4 1 12 7 12 9 3 15 13 2 3 9 1 10 9 9 0 2
26 10 0 9 1 9 13 16 15 13 10 7 3 12 9 2 15 4 0 15 1 10 9 1 10 9 2
25 10 3 0 9 7 10 9 15 13 1 10 0 9 13 16 15 4 0 1 7 0 7 0 9 2
19 10 9 13 16 15 13 10 0 9 2 7 10 9 4 3 7 3 0 2
10 0 4 16 15 3 13 9 1 9 2
8 1 9 9 4 15 13 9 2
18 10 0 9 2 10 0 9 1 9 1 9 2 4 3 13 1 11 2
7 15 13 13 2 9 2 2
23 2 7 3 4 15 3 13 10 3 2 9 2 2 16 15 4 3 0 2 13 11 11 2
19 3 3 3 0 7 9 4 10 9 1 10 9 1 10 9 15 13 3 2
19 9 13 1 9 2 7 15 4 3 0 16 15 13 9 1 15 1 11 2
20 3 13 9 10 9 1 10 9 1 9 9 7 10 9 1 10 0 0 9 2
6 15 4 10 0 9 2
12 10 9 1 10 9 15 13 1 10 9 1 11
5 9 7 3 9 2
14 15 4 3 4 10 0 9 1 9 15 4 13 3 2
16 9 7 9 13 0 9 14 13 1 9 3 1 9 1 9 2
14 3 3 3 3 1 9 2 7 3 3 3 1 9 2
16 10 0 9 4 15 4 9 1 3 3 1 12 9 1 11 2
9 3 13 7 9 7 9 1 9 2
10 4 15 13 13 1 9 1 10 9 2
18 3 4 15 3 13 15 12 1 16 15 13 9 7 9 1 9 3 2
14 9 1 9 13 3 16 15 4 4 13 3 1 9 2
19 3 13 15 1 9 2 7 15 4 3 3 0 1 9 16 15 13 3 2
7 3 9 13 4 9 13 2
13 3 13 9 1 9 3 0 7 1 9 7 9 2
16 3 4 9 1 9 13 10 3 0 9 7 15 15 4 0 2
22 15 13 1 16 10 0 1 15 4 13 3 0 9 1 9 2 3 15 13 9 1 2
15 15 4 13 9 1 10 9 3 0 1 14 13 10 9 2
17 7 0 9 15 13 3 1 9 2 3 0 9 13 15 1 9 2
14 1 9 7 9 4 10 0 9 13 9 3 0 9 2
9 9 13 3 9 1 10 0 9 2
27 1 14 13 10 0 9 7 0 9 1 0 9 9 2 4 15 13 15 1 14 13 9 1 9 1 9 2
9 15 13 3 12 9 1 10 9 2
6 3 13 10 0 9 2
10 9 13 3 3 1 9 7 0 9 2
8 1 9 13 15 3 1 9 2
10 15 4 3 0 14 13 3 0 9 2
14 15 4 3 13 3 3 7 12 9 2 3 12 9 2
19 13 15 9 15 13 3 3 1 9 13 9 9 1 9 1 10 0 9 2
6 9 13 10 0 9 2
8 15 13 1 0 9 1 9 2
12 3 13 10 0 9 3 1 16 15 13 15 2
7 3 13 9 1 9 3 2
15 15 13 3 9 1 9 7 3 13 9 0 9 7 9 2
10 9 4 13 1 3 0 9 1 9 2
21 3 15 15 13 9 3 7 0 9 13 13 9 1 3 0 9 7 9 7 0 2
5 15 4 1 9 2
22 15 4 0 1 9 2 1 9 16 9 9 4 0 14 13 10 0 9 0 9 13 2
12 10 0 9 4 3 4 13 7 13 1 9 2
17 16 15 13 0 9 2 13 15 3 1 16 9 13 1 0 9 2
14 7 1 9 7 1 9 4 15 3 0 1 0 9 2
10 1 10 0 9 13 0 9 0 9 2
6 9 1 0 9 13 2
28 13 15 1 3 2 3 4 15 3 3 0 16 10 0 9 13 0 14 13 15 3 1 9 7 10 0 9 2
12 1 10 0 9 13 9 0 7 3 3 9 2
22 10 0 9 7 10 0 9 13 15 1 9 1 9 2 9 2 9 13 15 3 2 2
13 10 0 9 4 1 9 3 1 9 0 1 9 2
12 3 4 9 1 3 0 9 13 9 1 9 2
16 1 9 13 9 10 0 9 2 1 9 16 15 3 13 13 2
6 9 13 3 3 0 2
14 9 1 9 4 1 10 9 9 3 0 1 0 9 2
36 11 9 1 9 7 10 0 0 9 15 13 13 1 16 9 1 11 7 11 9 3 3 13 10 0 9 1 0 9 2 0 9 7 0 9 2
5 9 4 3 13 2
12 0 9 13 1 12 9 0 3 3 1 9 2
9 9 3 1 9 4 13 10 9 2
13 3 15 3 13 4 10 0 9 13 9 1 9 2
21 10 9 2 15 13 2 13 1 10 0 9 13 3 3 1 9 1 10 9 9 2
16 15 13 3 1 9 0 9 2 3 9 13 3 1 0 9 2
16 3 13 15 9 1 10 0 9 1 9 1 9 1 0 9 2
18 15 3 13 15 3 10 9 15 13 10 0 7 9 2 10 0 11 2
17 10 9 7 9 1 3 9 4 4 0 1 10 9 13 3 3 2
15 1 11 1 10 0 9 9 4 15 13 3 3 1 9 2
12 15 13 3 9 2 15 13 9 1 0 9 2
22 15 4 3 13 9 3 12 9 1 10 9 1 14 3 9 7 9 4 13 3 0 2
1 13
14 3 15 13 9 1 9 3 2 13 0 9 10 9 2
17 1 10 9 9 4 15 13 9 7 3 13 9 1 0 0 9 2
20 1 0 9 4 9 4 0 2 16 15 3 13 10 9 14 13 9 1 9 2
15 13 15 3 10 0 9 4 9 13 1 9 1 10 9 2
21 3 9 3 13 13 15 3 1 9 9 7 9 1 9 1 9 1 9 1 9 2
14 0 9 4 1 7 1 10 0 9 13 3 3 3 2
23 15 4 0 2 16 15 3 3 1 9 1 9 2 7 1 9 7 0 15 2 13 9 2
10 3 4 3 10 9 9 13 3 3 2
1 0
23 3 15 3 13 13 15 3 3 0 3 1 9 7 9 1 9 1 10 0 9 1 9 2
9 1 14 3 13 1 9 1 9 2
20 1 11 9 1 11 1 11 4 15 1 0 9 13 3 10 9 1 11 9 2
24 9 13 10 9 2 16 15 13 3 0 9 1 9 7 3 4 9 13 0 9 1 9 9 2
23 9 1 9 13 3 16 15 3 4 4 0 1 9 15 3 4 4 9 1 3 0 9 2
9 15 13 3 14 13 9 1 9 2
1 0
27 9 4 10 0 9 2 15 4 0 1 9 2 9 7 0 9 7 15 4 3 13 3 1 9 7 9 2
16 9 1 3 10 9 4 3 1 0 9 0 1 9 1 9 2
17 1 11 9 13 15 9 0 7 4 13 3 3 12 9 1 9 2
14 16 15 13 12 9 1 9 13 9 1 9 3 0 2
13 9 1 9 13 15 1 9 13 12 9 2 9 2
20 1 10 0 3 9 4 15 1 10 0 9 3 1 9 13 9 1 9 9 2
25 9 9 4 3 4 10 3 0 9 2 7 15 4 3 13 10 0 9 15 13 1 9 1 9 2
3 9 10 9
15 1 9 13 10 0 9 1 11 7 11 13 10 0 9 2
7 12 0 9 10 3 9 2
9 1 9 13 10 0 9 1 11 2
7 3 13 0 9 1 11 2
19 0 11 13 1 15 16 9 13 13 15 3 1 9 16 15 4 13 11 2
8 9 1 0 11 7 11 13 2
10 9 7 9 1 11 13 10 9 0 2
18 3 13 15 0 1 15 15 13 1 0 9 2 15 1 11 0 9 2
17 1 9 3 12 13 9 10 9 1 9 2 12 9 9 1 11 2
23 15 13 3 3 2 7 9 13 16 9 1 9 3 1 9 4 13 3 12 9 1 9 2
21 9 2 15 3 13 0 9 2 13 3 12 9 3 1 11 7 13 15 1 11 2
8 9 13 12 9 3 1 11 2
10 0 9 1 0 9 1 11 13 3 2
15 10 0 9 13 12 9 3 1 11 7 13 3 1 11 2
10 15 4 13 14 13 9 3 1 11 2
7 9 4 13 1 1 11 2
3 0 1 9
21 15 3 4 10 0 9 1 15 15 13 1 11 2 11 2 11 2 11 7 11 2
11 9 13 16 9 13 3 12 9 1 9 2
7 9 4 13 9 1 9 2
6 9 13 1 12 9 2
10 11 9 4 3 13 9 1 11 9 2
13 9 1 11 13 2 7 9 13 16 9 13 0 2
6 9 13 1 0 9 2
23 15 13 2 0 0 9 2 9 3 9 2 9 1 9 2 9 1 11 1 10 0 9 2
7 0 9 4 13 1 9 2
25 1 9 7 9 2 1 9 7 9 4 9 9 7 9 13 15 9 2 9 2 9 2 9 3 2
11 3 16 15 4 4 13 9 1 9 3 2
22 11 4 3 13 1 10 0 9 7 4 1 12 0 1 11 4 13 1 9 1 9 2
19 9 11 11 2 9 11 2 0 9 2 13 3 10 0 9 13 1 9 2
14 15 13 16 10 0 9 4 15 15 9 4 13 1 2
35 2 16 10 9 1 10 0 9 13 9 1 10 9 1 9 9 1 0 9 2 0 12 2 15 13 4 13 10 1 11 3 3 0 9 2
8 7 7 10 0 7 0 13 2
14 15 13 9 11 11 7 9 11 11 1 9 1 11 2
15 7 15 13 16 3 0 4 10 0 9 3 3 3 0 2
22 7 13 15 1 9 3 13 10 0 1 15 1 0 9 1 11 11 9 1 9 9 2
44 10 0 0 9 1 10 0 9 4 11 11 2 10 0 0 9 7 9 2 15 4 13 9 1 9 2 1 9 1 0 9 7 9 2 9 2 9 2 9 2 9 7 9 2
14 15 13 16 3 1 9 4 9 9 0 1 0 9 2
20 15 13 16 9 3 4 3 0 1 16 9 4 4 13 15 15 13 1 1 2
28 15 3 9 13 3 13 9 3 16 15 13 1 0 9 1 10 0 9 0 9 2 15 3 3 13 1 9 2
28 1 9 9 2 15 1 9 13 1 3 12 9 3 2 3 15 13 0 1 9 0 9 14 13 10 0 9 2
8 10 0 9 0 0 9 3 2
17 6 2 15 13 3 16 9 3 2 2 1 9 2 13 0 9 2
10 7 3 13 1 11 10 3 0 9 2
25 1 10 0 9 9 1 9 13 1 0 9 2 11 11 11 2 0 1 11 2 7 9 11 11 2
38 9 12 13 1 11 10 9 1 9 0 9 1 9 9 2 0 9 1 9 2 7 15 13 13 7 10 1 10 0 9 1 9 1 10 9 1 9 2
30 10 0 9 13 3 10 9 1 0 9 2 15 3 3 13 1 0 9 1 9 1 9 1 1 15 9 11 7 9 2
6 15 13 10 9 12 2
2 11 3
15 11 13 10 0 9 15 13 10 0 9 1 0 10 9 2
24 9 7 9 13 1 15 12 2 1 9 0 9 4 15 0 12 7 9 13 1 9 0 9 2
15 15 4 3 3 3 1 11 7 3 7 3 1 0 9 2
32 3 4 0 9 13 1 0 9 3 7 15 2 11 7 11 1 0 9 2 2 7 15 4 3 13 9 1 0 9 7 9 2
7 3 13 15 3 1 11 2
8 9 4 0 1 10 0 9 2
9 11 4 3 3 10 3 0 9 2
27 6 2 15 13 1 9 1 10 9 0 1 10 2 7 10 0 9 13 1 9 16 10 9 4 3 0 2
1 9
8 1 15 13 15 1 3 3 2
17 7 3 13 15 7 13 10 0 9 0 9 3 3 1 0 9 2
18 1 0 7 9 13 3 3 10 9 1 9 1 10 0 9 1 9 2
20 10 0 13 1 0 9 3 1 9 9 2 3 1 16 15 13 10 9 15 2
22 7 15 13 3 9 15 4 0 1 10 0 7 13 16 15 4 13 7 0 7 0 2
10 3 9 13 1 9 13 9 11 0 2
14 2 15 4 3 3 4 13 16 10 0 9 4 0 2
18 15 4 0 16 13 15 9 1 0 7 1 9 0 9 3 13 9 2
9 3 16 15 13 10 0 0 9 2
21 1 9 13 3 12 9 1 10 9 1 9 2 3 13 15 3 1 3 12 9 2
17 7 1 15 13 3 10 0 9 1 9 2 12 9 3 9 13 2
5 15 13 3 9 2
18 13 15 3 3 0 9 1 0 7 0 9 3 4 9 3 0 2 2
2 3 0
18 7 3 15 3 13 15 3 3 4 15 13 10 0 9 0 1 15 2
20 7 7 15 9 3 13 0 7 0 9 2 3 3 4 15 10 9 1 15 2
23 9 11 4 13 3 1 9 7 13 16 15 3 1 3 4 13 16 10 0 9 13 0 2
29 0 9 14 13 9 13 14 13 9 13 3 1 0 9 2 13 15 1 0 9 13 7 13 3 1 9 7 9 2
37 1 10 0 9 1 10 0 9 4 15 1 9 1 0 9 1 9 4 13 3 0 9 14 13 9 1 10 9 15 3 13 3 1 0 0 9 2
17 1 15 13 10 0 9 3 3 3 3 1 0 9 1 0 9 2
9 1 9 3 4 15 13 3 0 2
6 9 2 15 13 9 2
23 2 9 11 4 13 15 10 0 9 2 7 13 15 15 15 12 9 12 13 13 15 3 2
4 3 12 2 2
7 3 13 9 11 11 3 2
9 4 15 3 10 0 9 1 9 2
3 9 11 2
4 2 6 6 2
3 3 15 2
8 9 4 13 3 0 7 3 2
20 15 4 1 9 3 4 13 1 9 1 10 3 16 10 9 4 13 3 2 2
3 9 11 2
4 2 6 6 2
3 10 9 2
21 15 13 16 9 1 10 0 9 13 16 15 3 3 4 3 0 1 14 13 3 2
15 3 13 15 3 3 2 12 9 12 4 3 3 12 2 2
21 1 10 0 9 15 9 13 1 14 13 1 0 2 0 9 13 9 10 0 9 2
12 9 13 3 3 2 9 4 10 2 9 2 2
20 7 15 4 0 16 15 13 9 7 9 2 15 13 3 1 10 9 7 9 2
18 1 14 13 9 10 0 9 1 9 1 9 13 3 11 9 10 9 2
23 15 13 9 1 3 10 9 7 9 2 15 13 15 14 13 0 9 1 14 13 0 9 2
23 9 4 0 1 0 9 2 15 15 7 15 13 0 9 1 9 2 0 9 2 9 3 2
25 11 9 2 15 13 1 9 12 2 13 7 9 14 13 3 0 9 3 2 1 9 7 1 9 2
10 9 4 1 15 13 10 9 1 9 2
11 3 1 11 9 13 15 3 12 0 9 2
11 3 13 15 9 1 3 12 9 1 9 2
25 7 3 13 7 9 7 0 9 2 15 13 15 0 1 9 7 15 15 13 9 14 13 0 9 2
22 9 13 1 12 9 1 9 2 0 9 2 9 7 2 1 10 9 2 1 0 9 2
9 10 0 9 2 7 3 3 13 2
20 9 13 3 10 3 0 9 1 9 2 15 13 15 1 9 1 10 0 9 2
16 15 13 15 1 9 1 9 3 3 15 13 1 9 7 9 2
34 9 13 7 1 10 9 2 2 13 1 14 13 1 9 2 2 15 13 3 1 9 2 7 1 9 1 10 0 9 1 9 7 9 2
24 7 15 13 3 10 0 9 2 15 13 0 9 1 9 1 9 2 15 13 10 3 0 9 2
5 9 1 9 13 2
22 3 11 9 13 1 11 2 11 2 11 7 11 1 14 13 9 13 15 1 9 9 2
10 1 9 13 3 9 13 1 10 9 2
17 1 3 9 13 15 0 14 13 9 1 9 1 0 9 7 9 2
4 3 13 9 2
12 9 4 0 1 12 9 1 10 10 0 9 2
15 10 0 9 1 9 13 1 0 9 2 9 7 0 9 2
17 3 13 9 2 9 2 9 2 9 2 9 7 9 2 9 3 2
11 10 0 9 13 15 15 4 13 1 9 2
17 3 13 9 2 9 2 9 2 9 2 9 1 7 9 1 9 2
30 10 0 9 13 1 13 2 14 13 3 7 1 2 13 2 13 9 2 13 9 2 13 9 1 9 2 9 7 9 2
23 10 0 9 13 1 14 13 2 13 2 13 2 13 7 13 2 13 9 2 9 2 9 2
18 9 1 10 9 13 9 7 9 2 9 2 9 2 9 7 3 3 2
23 10 0 9 13 1 14 13 15 2 15 13 14 13 2 13 2 13 2 13 7 13 3 2
17 9 4 10 0 9 1 9 9 1 10 9 1 10 0 9 9 2
39 7 16 15 1 10 9 13 15 1 10 9 1 9 1 14 13 3 2 3 13 9 15 1 10 9 1 9 1 10 9 1 16 15 4 13 1 10 9 2
4 13 1 1 9
15 1 9 13 9 14 13 1 10 0 9 1 9 1 9 2
8 13 9 14 13 9 3 3 2
14 13 15 10 9 1 9 9 2 16 15 13 1 9 2
7 3 4 15 13 9 3 2
8 4 15 4 0 1 0 9 2
15 4 15 10 9 14 13 0 1 7 13 15 1 0 9 2
42 10 9 2 15 9 1 0 9 4 0 1 4 2 1 9 2 9 2 12 9 2 2 9 2 12 9 2 2 9 12 2 12 9 2 7 9 12 2 12 9 2 2
15 9 4 13 7 0 2 9 13 3 3 3 1 0 9 2
21 0 0 9 4 3 13 1 1 0 9 2 13 3 1 10 0 2 0 9 2 2
15 9 4 0 1 10 0 9 2 15 13 9 1 0 9 2
7 15 4 3 13 0 9 2
7 2 7 3 0 2 9 2
11 7 3 4 3 10 9 13 2 13 9 2
34 15 13 0 9 1 9 2 15 15 0 13 4 2 3 9 2 7 15 1 9 4 0 9 2 9 2 0 9 2 9 2 0 9 2
21 7 3 0 9 7 9 7 9 2 9 2 9 7 0 9 1 14 13 10 9 2
7 1 9 13 10 0 9 2
22 9 1 9 2 15 13 1 1 9 2 4 13 1 9 2 1 15 1 15 13 9 2
16 1 9 9 13 15 3 1 16 10 9 4 3 0 1 9 2
13 15 4 9 2 15 13 1 9 1 9 7 9 2
17 3 13 11 11 2 15 1 9 9 2 9 1 10 2 9 2 2
12 9 4 13 1 12 9 1 9 1 12 9 2
15 9 2 15 13 1 0 9 2 4 14 13 3 1 9 2
9 10 0 9 4 14 13 1 12 2
21 15 4 13 1 9 2 7 10 9 4 1 0 9 13 1 9 7 3 1 9 2
14 15 4 13 16 10 0 9 4 13 0 9 1 9 2
32 1 10 0 9 9 13 0 16 9 9 7 9 1 0 9 1 10 9 2 7 3 7 1 9 7 0 9 2 13 0 9 2
21 3 4 15 0 14 13 16 15 3 13 13 10 9 0 9 1 10 3 0 9 2
32 13 0 2 13 1 9 2 6 2 3 0 4 15 3 14 13 9 16 11 7 11 4 13 9 15 13 3 10 9 7 9 2
9 4 10 9 13 15 10 9 13 2
12 6 2 7 15 13 3 16 15 4 3 0 2
16 9 4 3 13 2 13 15 3 7 4 3 3 1 0 9 2
7 3 13 15 3 9 9 2
18 9 4 13 10 0 9 1 14 13 1 9 2 3 3 15 13 9 2
20 3 13 15 3 1 9 7 13 1 15 15 4 13 1 0 9 15 13 3 2
14 7 9 13 15 2 13 3 7 13 7 13 15 3 2
4 13 10 9 2
4 3 13 15 2
27 15 4 3 3 4 10 0 9 1 9 7 1 9 11 11 2 1 9 1 11 2 13 9 9 14 13 2
6 1 9 1 3 9 2
9 3 1 9 13 3 3 12 9 2
9 10 0 4 3 0 1 10 9 2
23 3 13 1 9 10 9 1 11 3 0 9 13 3 10 9 1 2 10 0 1 9 2 2
7 3 13 15 15 10 9 2
11 15 4 9 1 14 13 10 9 1 9 2
10 9 4 3 1 10 9 0 1 9 2
14 7 15 4 3 13 10 9 10 9 4 13 1 9 2
18 9 1 10 0 2 9 1 15 15 13 9 2 9 3 9 3 13 2
18 9 15 13 15 4 0 14 13 9 1 9 2 2 9 2 1 9 2
5 7 3 3 9 2
27 1 9 13 9 11 11 1 9 0 9 16 15 3 3 13 16 10 9 13 10 0 9 14 13 15 9 2
10 15 13 0 9 3 15 13 9 9 2
4 1 9 3 2
19 9 11 11 1 9 1 11 13 16 15 3 13 9 12 9 9 1 9 2
4 15 4 0 2
11 9 4 13 12 2 3 12 9 1 9 2
12 15 13 3 9 15 13 15 1 12 9 9 2
22 7 7 9 7 9 13 3 2 7 13 15 9 3 2 16 9 13 3 1 0 9 2
3 3 0 2
7 3 0 4 3 10 9 2
16 9 11 11 2 0 9 2 13 3 0 0 9 1 10 9 2
14 10 9 4 13 1 10 3 0 9 1 10 9 9 2
17 7 3 2 1 15 0 9 2 4 9 3 3 0 1 10 9 2
8 10 0 9 4 10 0 9 2
14 10 0 9 4 10 0 9 7 3 3 2 0 2 2
8 7 15 13 15 1 10 9 2
5 3 13 9 9 2
15 15 9 13 3 13 10 9 7 10 3 0 9 1 9 2
11 3 4 3 9 9 7 9 13 10 9 2
17 10 0 9 4 13 3 9 1 9 15 13 1 12 7 12 9 2
13 1 10 0 9 13 15 3 9 15 13 10 9 2
10 1 9 13 9 3 3 7 10 9 2
10 9 4 3 3 3 0 1 0 9 2
14 9 13 3 3 3 3 1 14 13 1 9 1 9 2
7 3 13 15 1 9 9 2
18 9 4 13 16 15 13 14 13 10 9 14 13 1 9 1 0 9 2
17 7 15 13 3 10 0 9 1 15 7 15 4 3 0 1 9 2
21 15 4 3 13 3 16 9 1 3 13 1 9 7 4 10 9 15 13 1 9 2
7 3 4 9 0 1 9 2
3 9 13 3
10 9 13 10 0 9 1 10 0 9 2
14 15 9 4 3 13 15 10 0 9 10 9 13 1 2
16 9 9 13 10 9 15 4 12 1 12 9 0 7 1 15 2
25 7 3 13 15 15 16 10 9 4 13 0 1 10 9 2 16 15 3 13 9 1 10 0 9 2
8 3 13 9 9 3 1 9 2
15 9 13 9 7 9 1 10 0 9 1 15 15 13 3 2
15 15 4 4 13 9 1 15 15 13 2 15 13 3 9 2
14 7 15 4 3 4 13 15 1 15 1 10 0 9 2
8 3 13 9 7 13 3 0 2
13 9 11 13 16 15 3 13 10 0 9 1 9 2
10 15 13 3 3 7 3 1 0 9 2
23 9 11 13 1 10 0 9 3 10 0 9 2 10 9 2 13 1 9 1 10 0 9 2
11 1 12 9 13 15 1 9 1 10 9 2
10 9 13 0 3 9 13 15 10 9 2
4 9 13 3 2
24 3 1 9 13 9 1 9 7 13 9 0 2 7 3 0 2 9 1 10 9 7 10 0 2
9 9 1 9 13 3 1 12 9 2
8 10 9 13 3 10 0 9 2
8 1 9 13 3 0 0 9 2
16 7 15 13 15 3 15 9 16 9 4 9 15 13 1 9 2
9 7 3 9 11 11 13 10 9 2
14 2 15 15 3 13 1 9 4 3 3 13 10 9 2
8 7 15 15 4 3 13 15 2
3 9 1 9
1 9
13 9 2 9 7 9 13 15 15 13 13 1 9 2
7 15 13 1 10 0 9 2
28 15 13 0 16 1 0 2 3 0 9 10 0 9 13 10 0 9 7 9 1 14 13 3 9 1 10 9 2
18 15 13 10 9 2 3 9 9 7 9 1 9 13 3 10 0 9 2
24 15 4 0 16 9 13 7 13 7 16 15 13 9 1 0 9 1 14 13 9 7 3 3 2
17 9 13 15 1 9 7 1 9 15 4 13 1 9 7 1 15 2
17 15 4 10 9 15 3 1 0 9 4 13 3 1 10 0 9 2
25 9 13 3 1 9 7 4 1 10 9 1 9 10 0 9 2 15 13 3 3 3 9 13 0 2
14 15 13 3 10 0 9 1 9 14 13 9 1 9 2
13 9 4 3 13 10 9 0 9 1 9 7 9 2
21 15 13 9 9 1 0 9 2 0 9 7 9 2 7 15 13 9 9 7 9 2
13 9 13 3 1 10 9 15 13 13 1 10 9 2
9 2 11 11 2 9 2 9 12 2
3 9 7 9
25 10 9 1 9 4 13 16 12 7 0 9 13 1 12 2 1 7 10 0 9 7 10 0 9 2
33 15 13 3 1 9 2 12 9 13 3 3 2 2 9 2 10 9 13 0 9 2 2 9 2 10 9 13 0 9 2 7 9 2
11 9 7 9 13 1 10 0 9 1 9 2
10 9 13 3 1 9 15 3 13 9 2
16 15 13 3 10 9 1 9 7 10 0 0 9 13 1 9 2
34 9 2 15 13 3 1 9 2 13 3 14 13 1 0 9 2 10 0 9 13 1 0 9 3 1 2 9 2 7 15 13 3 9 2
13 1 10 9 13 10 0 9 1 9 7 1 9 2
16 11 11 4 10 0 9 15 4 13 3 9 1 12 0 9 2
9 15 13 3 0 0 9 1 9 2
4 9 2 12 9
3 9 2 12
3 9 2 12
3 9 2 12
5 0 9 13 2 12
3 9 12 9
3 9 7 9
18 15 13 3 9 2 10 9 7 2 0 2 9 1 12 7 0 9 2
29 1 10 9 13 15 3 0 0 9 7 15 13 9 7 9 15 1 9 7 1 10 0 9 9 4 0 1 9 2
12 15 13 3 9 15 3 13 10 0 9 0 2
3 9 7 9
17 15 13 3 3 1 0 9 3 15 13 15 15 13 9 1 9 2
14 3 3 13 11 11 10 0 9 2 3 9 4 0 2
17 1 10 3 0 9 4 10 9 2 1 9 10 0 2 10 0 2
16 1 10 0 9 13 10 9 3 3 2 1 10 0 9 2 2
16 9 1 9 1 11 7 11 13 3 9 9 1 9 7 9 2
7 9 9 13 15 15 13 2
7 9 7 9 13 10 9 2
21 2 13 10 0 9 1 10 9 2 15 13 9 9 14 13 10 9 1 9 2 2
7 9 13 1 10 0 9 2
9 2 13 9 1 2 9 1 2 2
6 9 13 10 9 9 2
9 9 13 7 10 9 1 9 13 2
12 9 13 9 3 2 4 15 15 13 9 9 2
13 0 9 1 9 1 9 4 0 1 10 0 9 2
11 9 13 9 1 10 9 7 3 9 13 2
10 2 9 1 9 2 9 12 3 2 2
23 16 15 3 13 1 9 13 15 1 9 10 0 9 2 10 0 4 3 3 13 1 9 2
24 2 15 4 3 4 0 14 13 3 1 10 9 15 15 3 13 1 9 2 9 12 3 2 2
17 9 1 9 1 10 0 9 4 3 3 0 7 3 0 14 13 2
24 15 13 1 0 9 3 3 3 7 3 1 0 9 1 9 2 7 9 1 9 13 0 9 2
30 15 13 0 9 15 13 1 16 10 0 9 2 9 7 9 2 3 13 10 9 15 3 4 0 7 10 0 13 3 2
20 1 0 9 13 15 3 9 9 15 13 10 0 9 1 3 9 1 9 13 2
23 1 10 9 15 11 11 7 11 11 13 1 10 9 9 13 15 9 15 13 10 3 9 2
18 15 4 13 1 10 9 15 13 2 15 15 13 3 3 1 15 2 2
9 7 3 3 13 15 9 1 9 2
2 13 1
24 3 13 9 1 10 3 9 1 10 9 15 15 13 3 1 7 3 13 15 1 10 0 9 2
2 9 9
16 3 9 1 9 13 1 1 11 2 13 15 3 3 9 9 2
20 1 15 1 0 7 9 9 13 9 3 2 16 9 3 3 13 15 1 9 2
29 15 4 13 15 3 1 3 0 9 7 0 4 16 9 9 3 13 0 9 1 9 7 1 9 1 10 0 9 2
25 10 0 3 13 3 1 0 9 3 10 9 7 9 15 0 9 13 2 15 4 3 13 1 9 2
7 9 13 9 10 0 9 2
5 3 13 15 3 2
22 10 9 14 13 9 9 4 14 13 10 9 15 3 4 13 7 15 15 13 1 9 2
11 15 4 13 1 16 9 3 13 0 9 2
5 10 0 2 0 2
3 10 0 2
6 10 0 2 0 2 2
5 10 0 7 0 2
5 9 1 9 3 2
2 9 2
4 10 0 9 2
4 10 0 9 2
5 3 13 15 3 2
19 10 9 13 3 9 1 9 7 15 1 15 13 3 10 0 9 1 9 2
13 15 13 3 0 9 3 2 3 13 15 3 9 2
11 9 7 10 9 1 9 4 13 1 9 2
32 16 15 13 0 9 2 13 15 15 1 10 9 2 7 16 15 13 9 1 0 9 13 15 1 10 9 7 10 0 0 9 2
26 10 0 9 1 10 9 13 1 9 7 1 10 0 9 15 13 9 7 9 3 10 0 9 1 15 2
9 3 13 9 3 10 0 0 9 2
16 0 4 14 13 10 9 15 4 13 1 9 1 10 0 9 2
31 15 13 10 0 9 1 10 9 14 13 0 9 2 1 0 9 2 7 15 13 4 0 16 10 0 7 0 9 4 13 2
38 10 9 15 13 1 15 4 7 10 3 0 0 9 2 13 9 12 2 1 10 0 9 2 7 0 9 1 0 9 1 9 7 7 0 9 1 9 2
1 13
10 3 4 10 3 0 9 1 9 13 2
9 10 9 4 15 13 1 0 9 2
19 9 9 13 1 9 1 12 1 3 12 9 7 13 3 1 3 12 9 2
16 15 13 10 9 1 9 1 12 9 10 9 7 12 10 9 2
14 9 4 0 1 9 2 3 0 1 11 1 12 9 2
25 16 10 0 9 13 2 4 9 9 14 4 13 10 9 3 1 9 2 3 1 3 7 12 9 2
14 9 9 1 9 12 1 12 7 11 9 1 9 12 2
22 3 1 10 12 9 3 4 9 0 7 13 3 1 10 0 9 7 10 3 0 9 2
22 10 0 9 13 3 1 0 7 0 9 9 1 10 0 9 2 3 1 10 0 9 2
19 1 9 12 4 3 0 9 7 9 0 9 13 1 10 0 9 1 9 2
21 1 11 2 11 7 0 9 1 0 9 4 3 10 3 0 9 4 13 1 9 2
6 3 0 9 4 0 2
7 1 9 13 9 3 1 2
34 1 0 9 4 3 15 13 0 1 10 0 9 2 7 9 4 3 3 1 10 9 13 0 9 1 9 2 15 13 3 1 0 9 2
14 9 4 13 16 10 0 9 1 9 1 10 9 13 2
9 0 9 4 13 1 9 1 9 2
11 9 13 3 1 10 9 1 9 1 9 2
34 9 1 9 4 3 3 4 13 1 12 9 1 14 13 9 2 7 1 9 1 0 9 4 15 4 4 12 9 3 0 7 1 9 2
10 3 4 9 1 0 9 0 1 9 2
7 9 13 0 9 7 9 2
6 4 10 9 4 13 2
5 9 3 4 0 2
10 0 9 4 3 0 2 15 3 0 2
15 1 12 9 4 15 0 2 9 4 13 1 10 0 9 2
17 15 4 3 13 7 4 13 1 10 0 9 2 16 15 3 13 2
11 9 4 3 13 7 0 9 16 0 13 2
15 9 1 9 7 9 4 13 2 3 16 9 9 3 13 2
22 7 10 0 9 4 3 13 7 0 9 13 1 9 2 15 3 13 3 3 0 9 2
18 3 3 13 4 9 1 9 10 0 9 1 9 1 0 9 1 9 2
23 9 13 1 9 1 0 9 2 7 9 1 0 13 1 10 0 9 7 1 10 0 9 2
24 0 9 13 15 3 3 0 1 14 13 1 9 2 7 9 4 13 14 13 9 1 10 9 2
36 0 9 4 13 10 0 9 2 7 9 1 11 4 13 2 16 15 4 13 15 1 9 7 9 2 15 13 1 10 9 1 0 7 0 9 2
6 1 3 9 13 9 2
18 10 0 0 9 2 3 1 11 2 13 3 1 14 13 9 1 9 2
17 15 13 9 1 10 9 1 9 3 1 10 9 1 15 9 13 2
14 3 13 15 13 9 1 14 13 9 1 10 0 9 2
17 2 9 2 1 11 2 0 1 9 2 12 9 9 1 9 2 2
15 10 9 1 9 2 3 2 7 12 9 3 2 3 2 2
25 1 0 9 1 9 4 15 1 0 9 13 9 1 14 13 9 1 9 1 14 13 15 1 9 2
13 9 13 3 9 16 0 9 4 13 3 0 9 2
11 9 9 1 9 4 10 0 9 1 9 2
26 16 15 1 11 7 11 13 0 9 9 1 9 2 4 0 9 3 0 1 9 7 13 3 3 3 2
11 15 4 3 0 14 13 9 1 10 9 2
7 3 9 1 9 4 13 2
9 1 10 9 4 9 13 0 9 2
7 10 9 1 11 4 13 2
18 0 0 9 13 3 0 9 2 1 16 15 13 7 13 1 0 9 2
26 16 15 13 2 16 9 13 9 2 4 15 1 9 1 12 9 9 1 9 13 9 3 1 12 9 2
15 0 9 13 1 9 2 3 15 13 14 13 9 1 9 2
24 1 14 13 9 2 9 12 2 9 12 2 1 11 13 9 3 16 9 3 4 0 1 9 2
18 1 0 11 4 0 0 9 1 9 7 9 13 13 1 3 0 9 2
19 10 0 9 13 3 2 7 1 10 9 13 15 12 7 12 9 1 9 2
16 10 0 9 4 0 7 13 0 9 1 9 1 14 13 9 2
12 1 9 2 9 7 9 13 3 9 1 11 2
14 10 0 9 13 9 1 14 13 3 0 9 1 9 2
35 10 0 9 1 9 1 0 9 4 14 13 13 3 9 1 0 9 7 0 9 1 9 2 3 10 9 2 13 9 12 2 9 12 2 2
15 9 7 9 13 9 1 9 7 13 9 1 9 7 9 2
14 1 0 0 9 13 9 1 12 9 1 10 0 9 2
15 9 1 0 9 2 9 7 9 1 9 4 3 3 0 2
17 0 9 1 9 1 10 9 1 9 1 10 0 9 4 3 13 2
15 3 4 15 16 0 13 9 1 0 9 2 9 12 2 2
19 9 1 3 9 1 9 4 3 13 0 9 7 4 4 13 3 0 9 2
24 9 4 13 1 9 1 9 2 0 9 1 9 2 9 2 0 9 2 0 9 1 9 9 2
13 1 9 4 15 0 1 0 9 2 9 12 2 2
15 1 15 13 10 0 9 1 9 9 1 9 1 0 9 2
19 1 9 1 9 4 3 15 3 1 10 9 13 2 3 1 10 0 9 2
12 7 15 4 0 2 16 9 3 13 3 0 2
28 1 10 9 13 3 10 0 9 1 9 1 9 1 9 1 0 9 2 7 0 9 1 14 13 3 0 9 2
23 0 9 2 3 9 7 9 7 9 2 3 3 10 0 9 2 4 13 0 9 1 9 2
12 1 10 0 9 4 9 3 3 0 1 9 2
30 9 1 9 7 0 9 13 9 1 0 9 1 10 0 0 9 1 9 2 3 11 7 11 2 7 3 1 0 11 2
18 3 13 15 1 9 0 0 9 2 7 9 4 13 9 1 0 9 2
14 1 9 1 9 9 4 15 3 13 0 9 1 9 2
10 3 3 13 2 4 9 9 3 0 2
21 1 0 9 4 1 15 11 7 11 13 3 9 1 3 0 9 7 1 0 9 2
49 0 0 9 1 9 1 9 1 9 3 7 1 9 1 0 9 13 3 10 0 9 3 3 1 10 0 0 9 1 11 7 0 9 1 0 9 7 3 1 0 9 1 10 9 7 1 0 9 2
14 1 0 9 13 9 1 1 14 13 10 9 0 9 2
27 1 0 9 4 15 3 13 0 0 9 1 9 2 16 0 9 4 13 1 9 1 9 1 10 9 9 2
20 1 11 7 11 4 1 0 9 13 10 9 2 15 1 9 13 10 0 9 2
22 15 13 10 0 9 1 9 15 13 2 7 3 3 7 0 9 13 1 9 1 9 2
32 15 13 1 11 7 11 7 13 3 7 9 1 9 7 0 9 2 10 1 9 1 9 1 9 3 0 9 1 10 0 9 2
26 10 9 13 3 1 0 9 10 0 0 9 1 9 7 11 2 15 4 0 1 10 0 9 1 11 2
44 1 0 9 1 9 4 15 1 0 9 4 13 10 0 9 1 0 9 2 7 11 2 9 7 9 9 1 10 0 9 2 13 1 16 15 1 10 9 4 4 13 9 9 2
21 9 2 9 2 9 7 9 2 13 7 9 1 11 2 9 12 2 9 12 2 2
21 3 1 11 13 9 1 10 0 9 2 7 0 9 13 1 0 9 1 0 9 2
11 10 0 9 13 3 1 9 7 9 9 2
18 15 4 0 2 16 9 4 14 13 10 3 0 9 7 3 1 9 2
27 0 9 1 9 2 0 9 2 9 1 9 1 9 2 9 1 9 7 9 1 9 2 9 1 0 9 2
18 1 9 1 9 1 0 9 4 15 13 9 14 3 13 9 7 9 2
14 14 1 9 13 9 1 0 9 13 15 3 3 13 2
19 3 0 4 10 9 15 1 0 9 13 1 9 1 0 9 1 0 9 2
9 0 9 4 3 13 1 9 11 2
23 10 9 4 0 1 3 9 7 9 7 4 13 15 0 7 9 1 9 1 9 7 9 2
9 1 0 9 4 9 4 3 0 2
22 0 0 9 1 0 9 4 15 15 1 0 9 13 1 14 13 9 7 9 1 9 2
10 1 15 4 15 13 9 7 0 9 2
30 3 4 9 3 0 2 7 16 0 9 13 7 9 2 13 9 3 3 0 7 4 13 7 9 3 1 9 1 9 2
15 1 10 9 4 10 9 13 1 0 9 7 9 1 9 2
28 10 3 0 9 14 13 9 13 1 10 9 2 9 2 2 15 3 3 13 1 0 9 2 7 15 3 13 2
32 7 15 13 3 0 9 2 15 13 9 7 9 1 9 2 7 15 4 13 1 0 9 1 9 2 7 9 1 9 7 9 2
11 0 9 4 3 13 1 9 1 0 9 2
26 3 16 9 9 4 4 13 1 0 9 2 4 1 10 9 10 3 0 9 14 13 0 1 0 9 2
13 9 4 10 0 9 2 10 9 1 9 0 9 2
29 3 13 15 7 0 2 7 10 0 7 0 9 1 9 1 15 15 13 2 10 9 1 9 1 10 0 0 9 2
28 1 9 1 10 9 15 13 9 4 15 13 10 3 0 0 9 2 3 3 10 0 7 0 9 7 3 13 2
9 2 11 11 1 11 12 12 2 2
26 11 11 4 1 10 9 9 13 10 0 9 1 9 9 7 9 9 1 9 7 1 15 13 9 9 2
33 9 4 1 11 0 2 1 9 9 7 1 0 9 0 9 2 14 13 9 9 2 13 0 9 7 1 10 0 9 13 0 9 2
5 10 9 4 0 2
9 0 4 10 9 2 0 10 9 2
7 2 1 0 9 9 2 2
17 10 3 9 13 12 3 0 9 3 15 13 9 1 9 7 9 2
17 10 3 3 0 9 1 10 9 4 1 15 13 15 1 12 9 2
9 4 9 10 9 7 10 0 9 2
11 10 3 9 13 3 3 1 9 1 9 2
18 15 13 3 1 9 2 16 9 4 10 0 9 2 15 3 13 9 2
12 7 15 13 3 3 2 16 9 9 4 0 2
6 9 4 10 9 1 9
23 10 9 7 10 9 4 3 3 13 3 7 13 15 9 2 1 16 10 9 13 7 9 2
35 1 16 10 9 1 10 9 7 10 9 4 13 7 9 2 4 9 13 7 13 2 1 10 9 15 13 1 3 3 7 10 9 9 3 2
16 3 10 9 13 3 2 16 15 13 9 7 10 9 1 9 2
10 0 9 13 0 9 1 9 1 9 2
25 10 0 9 13 1 10 0 9 2 10 0 9 4 3 2 1 9 2 13 10 9 14 13 3 2
7 10 0 9 13 10 9 2
18 1 7 0 7 0 9 13 10 9 1 9 1 10 0 9 1 9 2
19 15 15 3 13 10 9 1 9 1 9 13 15 3 1 9 7 0 9 2
17 7 15 13 15 1 0 7 0 9 0 9 7 4 0 0 9 2
13 7 9 13 3 3 1 9 1 9 1 9 9 2
17 9 9 13 3 9 1 9 7 9 2 9 1 0 2 9 3 2
13 9 13 3 1 9 1 9 2 9 9 7 9 2
21 1 0 9 4 9 1 0 0 9 7 9 13 1 3 9 11 11 3 1 9 2
8 15 13 0 1 10 3 9 2
24 9 10 9 9 15 13 3 7 13 0 9 2 3 1 14 13 0 9 2 13 3 9 2 2
17 1 9 4 13 10 7 0 9 2 9 2 9 7 0 9 2 2
12 1 9 13 3 3 10 9 0 1 9 7 9
10 9 4 3 10 9 7 9 1 9 2
17 15 13 3 3 1 9 7 10 0 9 2 0 1 9 0 9 2
6 9 4 3 7 3 13
21 15 13 15 3 0 2 16 10 9 1 0 9 13 1 12 9 9 7 0 9 2
9 7 10 9 4 13 1 3 3 2
20 9 1 9 2 15 3 13 1 10 0 9 2 13 10 3 0 9 1 9 2
6 15 13 10 9 1 2
23 10 0 9 4 15 13 3 1 14 13 9 2 15 13 15 15 13 3 9 1 0 9 2
31 1 10 0 9 13 15 1 0 9 9 15 13 2 3 3 9 7 0 9 2 7 3 3 10 0 9 7 3 3 9 2
17 3 3 3 1 9 4 9 0 9 1 9 10 0 9 1 9 2
22 1 10 7 0 9 13 0 2 0 7 0 9 7 9 2 15 13 7 0 1 9 2
6 15 13 3 15 13 2
31 14 13 15 3 10 9 13 3 3 10 9 1 3 7 3 0 2 1 15 0 9 7 13 3 3 0 9 7 0 9 2
22 9 1 9 13 1 10 9 1 9 9 1 9 9 1 10 0 9 1 9 1 9 2
26 9 1 9 0 9 2 13 2 2 15 4 3 3 10 9 7 10 9 1 9 2 9 9 1 9 2
17 1 9 1 10 9 4 9 9 13 1 10 3 0 9 1 9 2
16 7 9 7 9 4 1 0 9 7 3 0 9 1 0 9 2
20 15 4 3 7 3 13 0 9 2 3 9 2 9 2 9 7 9 4 9 2
14 9 4 1 9 3 7 3 13 10 0 9 1 0 2
27 0 0 9 7 9 2 15 13 10 0 9 2 9 7 9 1 10 0 9 1 10 9 2 4 3 13 2
30 15 13 3 3 7 9 1 10 7 10 9 1 9 3 0 9 13 9 7 7 9 1 0 9 14 13 1 0 9 2
15 10 0 9 4 3 13 9 10 0 9 0 1 0 9 2
36 10 0 9 2 10 0 9 1 12 0 9 2 13 3 9 1 10 0 9 3 7 9 7 13 10 0 9 1 9 2 9 7 9 1 9 2
18 9 1 9 9 7 9 0 7 9 4 10 0 9 1 10 0 9 9
16 9 4 2 3 15 13 1 10 9 7 9 2 10 0 9 2
18 7 3 4 15 3 7 3 13 0 1 9 14 13 10 0 9 0 2
18 15 4 3 0 2 16 15 3 13 10 9 1 9 0 7 0 9 2
16 0 9 4 1 0 9 9 1 10 9 15 13 10 0 9 2
37 1 7 1 16 9 1 9 13 0 7 9 7 9 2 4 9 1 9 9 7 9 7 1 10 0 9 1 9 13 3 3 0 7 0 7 3 2
15 3 13 10 0 7 0 9 3 7 1 15 3 3 9 2
9 15 4 10 9 1 15 7 9 2
14 3 3 4 10 9 4 13 1 10 0 0 7 9 2
21 16 15 3 13 0 9 7 0 9 7 9 15 13 3 9 2 15 4 15 3 2
5 15 4 10 9 2
6 15 13 15 1 9 2
12 0 9 4 1 10 0 9 13 0 7 3 2
4 15 4 9 2
7 15 4 10 9 7 9 2
5 15 4 3 13 2
13 15 4 9 1 16 12 9 13 3 1 10 9 2
6 1 9 4 9 10 9
22 9 13 3 0 9 1 0 9 7 11 7 11 2 3 10 0 9 13 10 0 9 2
19 15 13 3 1 10 0 9 9 1 9 7 10 0 9 2 0 14 13 2
18 16 15 4 10 9 13 2 16 15 4 2 10 9 14 13 11 2 2
16 1 10 0 9 1 9 13 15 12 0 9 15 13 9 3 2
24 10 0 13 16 15 13 10 9 15 13 3 9 4 13 2 9 7 9 1 11 7 10 0 2
6 15 4 13 15 9 2
16 15 4 9 9 14 13 10 0 9 15 11 13 3 1 9 2
22 16 15 13 15 2 4 15 13 10 0 9 2 9 2 15 4 1 15 13 11 9 2
24 10 9 13 3 3 3 9 7 10 9 13 10 9 15 13 9 14 13 3 1 9 2 9 2
10 3 4 15 13 10 0 9 2 9 2
7 9 13 10 9 1 12 9
14 1 9 1 9 9 4 10 0 9 1 9 3 0 2
18 9 4 1 9 13 3 10 9 1 12 9 2 12 0 7 12 0 2
7 10 0 4 15 13 9 2
14 15 13 2 16 9 13 3 1 10 0 9 1 9 2
21 10 0 9 2 15 13 16 9 7 9 13 1 15 2 13 7 10 9 1 11 2
17 11 4 13 9 1 10 0 9 1 9 9 7 3 1 9 9 2
17 9 7 9 4 3 1 10 0 0 9 4 9 9 7 0 9 2
12 1 10 9 13 9 3 7 11 9 7 9 2
14 3 4 3 10 0 9 13 1 9 1 0 0 9 2
28 15 13 3 3 0 9 3 15 4 13 1 9 2 16 9 7 10 0 9 3 4 13 10 0 9 7 9 2
30 9 13 3 3 10 9 2 9 4 15 13 1 16 15 1 15 3 4 4 13 0 9 7 0 9 7 10 0 9 2
26 9 0 9 4 3 0 2 9 13 1 1 14 13 0 9 7 3 13 9 1 0 9 1 10 9 2
26 3 13 15 1 9 13 10 3 9 10 0 9 2 15 13 3 1 9 9 3 10 0 9 13 0 2
25 3 3 2 13 15 2 4 9 13 10 0 9 14 13 10 0 9 7 14 13 9 1 0 9 2
2 0 9
10 15 13 3 0 9 1 3 0 9 2
14 15 13 2 16 9 0 9 4 13 1 10 0 9 2
10 1 9 1 10 9 13 9 10 9 2
19 1 0 9 13 10 9 1 10 0 9 7 10 0 9 1 12 0 9 2
14 3 13 3 10 0 9 10 9 2 1 9 1 9 2
23 10 9 2 3 9 7 10 0 9 7 9 13 1 9 13 2 13 15 7 9 7 9 2
13 10 3 0 9 4 15 4 13 10 0 9 9 2
17 15 15 13 3 10 0 9 4 1 15 9 1 0 7 0 9 2
14 16 15 13 2 13 15 10 0 9 1 10 0 9 2
3 3 9 2
3 3 9 2
7 9 4 1 10 9 0 2
11 0 9 13 9 7 13 10 9 1 9 2
10 1 0 0 9 13 9 1 9 9 2
14 1 14 4 10 0 9 4 15 4 0 2 13 15 2
7 7 3 4 9 4 0 2
9 10 9 4 13 0 1 10 9 2
18 15 4 3 0 2 16 9 3 7 3 13 7 10 0 9 1 9 2
21 7 15 4 0 2 16 15 13 15 2 16 3 9 13 9 0 0 9 7 9 2
31 10 9 1 10 0 9 1 9 2 10 0 9 1 9 4 2 7 1 11 7 9 0 7 15 4 3 0 14 13 15 2
28 15 4 3 13 15 3 7 3 13 9 2 10 0 9 7 9 7 13 1 16 15 13 1 0 7 0 9 2
24 15 4 3 1 10 9 13 9 1 10 0 9 1 3 9 16 15 4 13 15 0 1 15 2
30 15 4 13 15 3 0 14 3 13 10 0 9 1 9 9 2 16 15 13 16 10 0 9 3 13 1 0 9 2 2
8 2 11 2 9 0 9 2 2
3 3 9 2
6 10 0 13 12 9 2
15 1 10 0 4 9 4 0 2 3 16 15 4 11 9 2
22 15 13 2 13 15 2 1 11 9 7 9 9 1 0 9 2 1 14 4 3 0 2
9 9 4 3 0 2 1 0 9 2
26 1 9 10 9 13 11 11 10 9 15 13 1 10 0 9 7 3 13 10 0 9 1 10 0 9 2
18 9 13 10 9 2 15 13 3 10 9 2 15 1 9 13 10 9 2
13 1 10 0 9 4 9 13 7 3 0 7 9 2
4 9 7 9 2
22 10 0 0 9 13 15 1 9 2 15 4 13 3 16 9 13 10 0 1 10 0 2
21 10 0 9 1 9 7 1 9 2 9 7 9 4 2 13 0 9 2 3 9 2
13 10 0 9 1 9 4 3 3 0 9 0 1 2
28 15 4 4 10 3 0 9 2 16 7 9 7 0 9 1 0 0 9 4 13 16 9 13 3 1 0 9 2
18 10 3 0 9 1 9 1 2 9 2 13 3 10 0 9 1 11 2
8 2 10 9 9 4 3 13 2
74 4 9 3 13 9 1 9 2 9 16 10 9 9 4 13 1 16 15 13 10 9 14 13 9 2 16 10 0 9 7 9 4 13 1 9 7 9 2 7 3 4 10 0 9 3 3 13 2 2 16 9 2 15 3 13 9 14 13 10 9 2 3 4 13 7 13 15 1 0 9 15 13 13 2
16 15 15 13 15 13 1 0 9 4 12 9 13 0 1 0 2
16 9 4 3 7 4 3 14 13 13 1 7 15 9 7 9 2
28 16 15 13 10 9 2 15 13 3 1 10 0 9 1 10 0 2 4 10 0 9 7 9 13 15 1 9 2
17 15 10 9 4 2 3 4 15 1 9 1 7 15 9 7 9 2
9 7 3 0 1 9 7 9 2 2
11 2 11 11 1 11 11 11 9 12 2 2
4 9 7 3 2
23 15 13 3 2 7 1 0 7 0 9 14 13 2 15 15 13 1 9 7 9 1 9 2
16 3 13 3 10 9 14 13 1 10 9 2 16 0 9 13 2
19 16 15 2 1 10 9 1 9 2 13 9 2 1 10 9 13 15 15 2
3 0 9 2
6 9 0 1 9 7 9
12 10 0 9 13 9 9 1 10 3 0 9 2
24 1 10 9 4 9 10 9 7 4 7 15 3 13 2 7 15 1 9 2 0 9 7 9 2
8 3 13 15 16 0 9 13 2
14 9 13 3 2 16 10 0 9 1 9 13 1 9 2
3 11 9 2
4 9 1 9 9
8 10 0 9 9 13 10 9 2
18 9 13 7 10 9 2 9 2 1 0 9 7 4 3 1 9 0 2
13 7 10 9 13 3 3 14 13 1 9 0 9 2
12 1 9 9 13 10 0 9 7 9 7 9 2
23 15 13 3 10 9 1 0 9 7 9 2 15 13 1 0 9 9 14 13 3 1 9 2
24 9 4 1 0 9 10 9 1 9 2 7 3 0 9 4 3 9 1 0 9 7 4 3 13
18 9 13 3 3 1 10 0 9 1 9 2 3 9 1 15 1 9 2
7 15 13 10 9 1 11 2
25 2 15 15 1 10 0 9 9 7 1 9 13 15 7 13 15 10 0 9 2 15 13 9 2 2
15 9 4 1 9 9 1 10 9 4 10 0 9 1 9 2
14 15 4 3 4 14 13 10 0 9 1 9 7 9 2
26 9 4 15 2 10 9 2 3 9 3 13 10 9 1 15 7 3 13 15 2 4 3 13 10 9 2
27 10 0 9 4 3 14 13 13 15 0 1 14 13 15 15 15 13 1 10 0 9 2 9 1 0 9 2
20 1 10 0 9 13 15 1 9 2 15 4 13 3 2 16 9 13 10 0 2
24 16 10 9 9 1 14 13 3 3 13 15 4 15 1 9 10 0 9 1 9 2 13 15 2
24 16 0 9 1 9 3 13 9 0 9 2 4 15 1 9 13 3 10 9 1 14 13 9 2
25 15 13 3 1 3 0 9 3 1 14 13 9 2 15 13 3 10 0 9 2 1 9 0 2 2
12 9 7 3 2 15 13 15 15 3 4 0 2
23 7 1 9 7 3 0 13 2 16 10 0 9 1 10 9 13 1 0 9 1 9 9 2
16 7 0 9 15 13 9 2 3 3 13 4 9 1 9 9 2
4 9 7 3 2
10 10 0 9 4 13 15 1 12 9 2
23 1 10 0 9 13 15 1 10 9 1 14 1 9 13 9 2 16 15 4 0 7 0 2
31 1 10 0 9 4 15 13 9 1 9 2 3 0 4 10 9 4 1 16 15 4 13 9 14 13 15 0 1 10 9 2
10 3 4 9 1 9 7 9 13 3 2
20 3 2 10 9 9 13 1 9 2 10 9 9 13 14 4 9 2 9 7 9
29 3 2 3 13 10 12 9 9 2 9 7 9 2 2 10 9 1 10 9 4 0 1 9 0 2 9 7 9 2
15 3 2 15 2 9 7 9 2 1 9 3 0 1 3 9
29 3 2 3 13 10 12 9 9 2 9 7 9 2 2 10 9 1 10 9 4 0 1 15 0 2 9 7 9 2
25 9 7 9 9 1 10 0 9 13 3 1 11 3 3 3 7 15 15 13 1 3 12 9 3 2
10 15 4 3 3 13 9 1 12 9 2
22 10 0 4 0 1 10 0 9 2 9 7 9 13 10 0 7 3 0 9 7 9 2
21 1 10 0 9 13 9 3 1 9 1 9 2 16 9 13 3 1 9 1 9 2
25 10 0 1 10 0 9 4 16 9 7 9 3 13 14 13 2 3 4 15 13 10 9 7 9 2
10 10 3 0 9 14 13 9 1 9 2
22 9 1 3 10 0 9 4 13 3 4 1 3 0 4 0 1 0 7 0 1 11 2
7 15 13 7 9 7 9 2
10 15 13 3 4 3 3 1 0 9 2
69 2 3 9 7 9 2 7 9 7 9 1 7 9 7 9 2 3 9 7 9 2 15 13 14 13 9 7 1 10 0 9 13 13 3 1 10 0 9 1 9 7 9 2 3 9 7 0 9 2 1 16 10 9 4 4 0 2 4 15 13 9 1 0 9 2 9 7 9 2
15 1 10 9 4 15 13 14 13 10 0 9 1 0 9 2
15 9 4 1 9 13 1 14 13 9 2 0 9 7 9 2
16 9 7 9 4 13 1 9 7 13 1 14 13 9 7 9 2
16 10 0 9 13 9 2 3 15 13 15 14 13 7 13 9 2
10 15 13 3 0 9 1 9 7 9 2
16 1 3 0 9 4 15 13 9 1 9 1 3 3 0 9 2
15 1 9 1 9 2 9 7 9 4 9 3 13 1 9 2
13 7 10 3 0 9 13 9 3 1 9 1 9 2
18 15 13 2 4 15 13 2 10 9 2 15 13 9 1 10 0 9 2
15 1 10 9 9 4 10 0 9 3 3 13 3 10 9 2
17 9 13 3 1 9 2 9 13 1 9 7 9 7 9 1 9 2
29 10 9 1 10 9 2 15 13 9 1 10 0 9 2 4 13 1 14 13 9 2 9 2 9 2 9 7 9 2
12 9 2 2 9 2 2 9 15 13 1 9 2
22 1 0 9 13 15 3 10 9 2 16 10 10 9 1 10 7 0 9 13 1 9 2
32 9 2 9 2 9 2 9 7 9 4 1 0 9 0 9 2 7 9 4 10 9 1 10 1 9 0 9 7 9 1 9 2
15 7 3 4 15 3 13 15 10 9 2 15 13 1 9 2
19 16 9 4 10 9 1 9 2 13 9 16 10 10 9 3 13 1 9 2
5 3 3 13 9 2
16 10 3 0 9 7 9 4 13 1 10 0 9 1 9 9 2
17 3 1 10 9 13 15 10 3 0 9 1 0 9 7 0 9 2
21 3 15 4 13 1 0 9 2 13 15 10 0 9 1 10 9 9 7 10 9 2
11 0 9 1 9 1 9 9 13 3 9 2
16 15 13 3 10 0 9 1 9 7 9 9 1 10 0 9 2
17 1 14 13 10 9 4 15 3 13 1 12 9 2 9 7 9 2
5 9 9 2 9 2
10 10 0 9 13 10 2 0 2 9 2
13 9 4 10 9 2 15 13 0 1 10 0 9 2
24 1 9 1 9 1 9 2 3 9 1 9 7 9 1 0 9 2 13 15 3 1 9 9 2
18 15 13 10 9 15 13 1 9 9 1 9 1 9 2 9 7 9 2
20 1 14 4 13 3 9 4 15 3 13 10 0 9 1 0 9 2 3 9 2
22 9 1 9 4 3 1 9 12 2 1 9 12 2 1 9 12 2 7 1 9 12 2
20 1 0 9 4 15 3 13 2 3 9 9 13 1 9 7 3 3 9 13 2
23 16 15 3 13 1 3 0 9 7 9 7 9 2 4 10 0 0 9 0 7 12 9 2
10 9 2 9 1 0 9 7 0 9 2
5 13 3 1 9 2
21 13 15 3 3 1 10 0 0 9 2 13 9 3 0 7 13 3 3 12 9 2
12 9 1 3 10 9 13 1 9 1 12 9 2
14 9 9 12 2 12 2 12 7 12 0 1 9 9 2
10 9 3 13 3 10 0 9 1 9 2
13 9 7 9 13 3 10 9 1 9 1 9 9 2
18 0 4 3 14 13 10 3 0 9 2 15 9 13 1 9 0 9 2
23 10 0 9 1 9 9 13 1 9 2 16 11 0 13 1 3 12 9 1 9 0 9 2
12 11 13 3 3 12 9 7 11 3 12 9 2
24 10 12 9 2 15 3 13 3 12 9 1 9 9 2 13 3 1 3 12 9 1 9 9 2
19 9 13 3 10 0 9 7 9 7 13 3 10 0 9 1 9 7 9 2
10 9 9 7 9 1 9 1 9 1 9
7 2 0 1 9 9 9 2
8 3 12 2 12 9 9 2 2
18 1 9 3 1 9 9 4 9 1 9 13 1 3 12 9 1 9 2
17 13 15 3 1 9 12 4 9 4 3 0 7 13 3 12 9 2
22 16 3 9 13 2 4 15 13 1 16 9 1 10 0 9 4 3 0 7 10 9 2
9 3 4 3 9 14 13 1 9 2
18 9 1 9 13 1 10 9 9 7 4 3 3 13 10 3 0 9 2
10 7 13 15 13 13 3 1 9 12 2
10 9 13 3 10 9 1 3 12 9 2
8 10 9 4 3 13 1 9 2
21 16 10 9 4 13 2 4 15 13 1 10 0 9 7 9 1 7 9 7 9 2
13 10 0 9 4 3 14 13 10 0 9 1 9 2
21 7 9 4 3 13 9 1 9 2 9 7 0 9 1 14 3 13 10 0 9 2
25 3 16 10 0 9 4 13 1 10 0 9 1 9 2 4 9 1 9 14 3 13 1 12 9 2
16 3 9 12 4 15 3 4 3 12 9 0 7 1 9 9 2
16 4 15 3 0 14 13 10 0 9 1 9 1 10 0 9 2
11 13 10 9 1 9 1 1 10 0 9 2
4 0 2 0 2
20 9 0 9 13 1 0 9 1 12 9 9 7 13 1 0 9 3 12 9 2
26 7 16 15 13 1 16 10 9 9 4 13 10 0 9 1 9 7 11 2 13 9 3 3 12 9 2
12 1 9 2 1 2 9 2 2 3 1 9 2
11 1 0 9 13 9 13 3 12 9 3 2
21 3 13 16 9 3 4 13 1 14 13 10 9 1 3 12 9 9 9 1 9 2
15 15 1 10 9 4 2 3 15 3 4 13 2 3 0 2
17 7 15 13 1 16 15 3 4 13 1 0 9 1 10 0 9 2
16 1 15 13 15 10 0 9 3 0 7 1 3 10 9 3 2
31 1 7 1 16 9 1 10 9 13 10 0 9 1 9 2 9 7 9 2 4 9 1 10 9 7 9 13 10 0 9 2
16 15 13 4 3 1 12 9 0 7 0 10 9 1 0 9 2
22 0 9 2 9 15 13 10 9 1 0 9 1 9 7 9 2 3 9 7 9 2 2
1 9
9 15 4 10 0 9 1 10 9 2
9 15 13 1 9 0 9 9 9 2
17 3 3 4 9 0 9 1 9 9 9 9 14 13 1 0 9 2
8 10 9 13 1 9 7 9 2
13 13 9 1 3 15 13 0 9 1 9 7 9 2
9 13 13 3 10 9 3 4 13 2
8 10 9 13 0 9 1 9 2
13 13 10 9 15 1 9 4 13 14 3 13 9 2
6 10 9 4 15 13 2
13 3 9 1 9 7 9 4 13 1 10 0 9 2
19 9 9 13 1 10 0 9 3 1 9 0 9 2 3 1 9 7 9 2
12 9 13 3 10 9 1 9 7 9 7 9 2
24 9 9 2 3 12 9 1 9 2 13 15 3 10 9 1 9 2 3 12 9 1 9 2 2
27 10 3 0 9 4 9 2 15 4 0 1 9 7 9 7 13 15 1 9 1 7 9 2 9 7 9 2
11 9 4 1 10 9 4 7 0 7 0 2
10 0 2 7 0 2 2 0 1 9 2
22 0 2 7 0 2 2 0 1 9 7 9 2 15 4 13 1 9 2 9 7 9 2
10 9 1 9 7 0 9 1 0 9 2
10 1 0 9 13 9 1 9 1 9 2
15 1 10 0 1 9 13 9 1 11 1 10 9 1 11 2
17 1 10 9 13 9 3 3 1 0 11 7 3 1 11 7 11 2
23 16 9 1 9 7 9 4 3 0 2 13 9 1 9 7 0 9 3 1 9 1 9 2
10 15 13 3 1 9 1 3 0 9 2
34 1 0 9 2 3 11 7 11 2 13 9 1 0 9 14 13 3 0 2 16 9 3 13 0 16 15 3 4 13 3 1 0 9 2
26 1 10 9 7 9 2 9 7 9 1 9 4 13 1 9 2 13 9 10 0 9 1 9 15 1 2
29 3 4 3 9 1 9 2 7 15 15 13 1 9 2 3 9 2 7 1 9 2 3 0 7 1 10 0 9 2
8 9 13 3 0 9 7 9 2
14 15 13 1 9 3 1 16 9 13 0 9 7 9 2
29 10 0 9 4 3 1 9 7 9 1 9 0 1 9 2 3 1 10 0 9 1 11 2 11 2 11 7 11 2
22 10 9 15 4 13 0 9 2 13 1 0 9 9 1 10 9 2 3 10 0 11 2
8 3 13 3 9 10 0 9 2
38 14 13 9 2 9 7 3 9 13 0 9 2 3 9 2 9 7 9 2 2 7 3 3 9 4 1 9 2 13 9 3 0 7 1 10 0 9 2
11 9 2 0 9 2 3 9 7 9 2 2
11 0 9 13 3 1 14 13 9 1 9 2
30 1 11 13 15 14 13 9 1 9 1 9 2 7 1 11 13 15 13 3 9 1 14 13 0 7 0 9 1 9 2
17 0 9 13 3 14 13 9 3 1 9 1 14 13 9 1 9 2
11 9 2 1 0 9 0 9 1 9 3 2
21 10 0 0 9 4 2 16 9 7 9 4 7 0 7 0 14 13 1 7 9 2
29 15 4 3 1 9 0 9 7 0 9 1 9 13 3 0 9 1 9 9 2 15 3 1 3 12 9 4 0 2
1 9
10 1 10 9 4 9 3 10 0 9 2
8 1 10 0 9 4 9 13 2
13 1 10 9 4 15 1 9 3 3 13 1 9 2
13 10 9 13 2 16 15 3 4 13 9 7 9 2
28 15 1 10 12 9 11 2 11 7 11 13 10 9 1 9 3 9 9 3 9 9 3 3 9 9 7 9 2
5 13 9 1 15 2
19 13 14 1 3 9 9 13 10 9 1 9 1 0 9 1 9 1 9 2
16 10 9 4 1 9 1 9 12 13 1 9 1 9 7 9 2
5 9 13 9 1 15
16 1 10 9 13 10 9 10 0 9 2 15 13 10 0 9 2
5 9 2 3 9 2
11 3 2 10 9 10 9 13 1 10 9 2
27 10 9 4 13 10 9 1 0 9 2 3 1 14 13 1 9 1 10 9 7 1 14 13 9 7 9 2
24 15 4 3 13 10 9 7 10 9 1 9 9 1 15 2 3 1 14 13 9 1 10 9 2
23 10 9 10 9 13 1 0 7 0 9 13 1 9 1 9 0 9 7 9 9 7 9 2
16 15 15 4 9 1 10 9 4 13 10 0 9 1 10 0 2
18 1 10 0 9 1 10 0 9 13 10 0 0 9 2 10 0 9 2
22 9 2 10 9 15 13 1 10 9 3 1 9 1 16 15 13 10 0 9 1 9 2
38 9 4 0 1 9 7 9 1 9 2 1 9 7 10 0 9 1 10 9 2 1 2 9 2 7 2 9 2 1 10 9 2 1 9 7 1 9 2
16 3 3 0 9 4 0 1 0 9 2 15 13 1 0 9 2
31 10 9 4 13 15 1 0 9 2 3 15 13 15 1 9 7 9 2 9 2 9 2 9 3 1 15 15 13 0 9 2
8 9 4 13 13 10 0 9 2
6 2 13 9 12 2 2
23 15 4 10 9 1 15 14 13 9 7 9 1 10 9 15 13 1 10 9 1 0 9 2
10 15 7 15 1 15 13 0 0 9 2
11 10 0 9 13 1 9 1 10 0 9 2
1 9
11 15 1 10 9 15 15 13 1 4 9 2
16 0 9 13 1 15 3 3 16 15 4 0 1 9 7 9 2
23 10 0 1 10 9 15 13 1 15 1 9 4 0 7 13 3 1 10 9 15 13 1 2
18 15 1 10 0 9 1 15 15 4 0 3 0 4 3 13 1 9 2
22 9 13 3 3 16 15 13 9 1 14 13 10 0 9 1 15 15 13 10 0 9 2
17 9 13 3 9 9 1 9 9 1 15 1 10 9 1 15 0 2
25 15 4 3 13 9 15 13 1 16 9 13 0 9 1 3 3 15 4 13 1 10 9 7 9 2
18 1 10 9 12 1 9 7 9 13 12 9 7 12 9 1 0 9 2
55 3 13 15 12 16 15 4 3 0 16 15 13 1 9 3 3 7 0 2 12 16 15 4 13 3 1 9 16 15 13 0 2 12 16 15 13 16 15 13 1 9 7 3 2 12 16 15 4 13 9 3 3 15 13 2
10 15 13 3 15 15 13 3 1 15 2
21 15 7 15 1 9 4 13 15 1 10 12 9 15 4 10 0 1 15 7 15 2
10 9 13 15 1 9 1 9 3 9 2
8 1 9 13 3 9 7 9 2
20 7 3 1 9 7 9 13 9 7 9 3 0 9 14 13 3 1 0 9 2
26 3 3 3 4 15 10 0 9 1 9 3 1 15 15 13 1 9 9 1 15 3 15 13 10 9 2
28 16 9 9 1 9 9 4 0 7 16 15 3 4 13 1 0 9 1 9 0 2 13 3 9 3 15 1 2
18 15 4 3 0 7 9 1 15 1 10 0 0 9 15 13 1 9 2
5 10 9 13 1 9
24 1 10 3 0 9 13 10 0 9 15 15 13 1 9 14 13 15 2 10 3 0 9 2 2
16 0 9 2 10 0 9 1 10 3 0 9 13 14 13 15 2
14 9 7 9 1 10 0 9 4 1 10 9 3 0 2
22 15 1 9 1 10 9 9 4 1 3 0 9 13 3 3 15 13 16 9 13 15 2
10 15 4 13 10 0 9 12 9 15 2
28 9 13 16 9 2 15 1 10 9 4 3 0 2 1 10 9 3 13 15 10 0 9 2 0 1 0 9 2
12 15 7 15 4 3 1 9 13 10 0 9 2
10 9 2 15 15 15 13 0 9 1 2
16 9 1 9 1 10 9 4 4 10 9 1 9 1 10 9 2
30 1 0 9 1 9 13 10 9 2 7 15 4 3 13 3 9 1 9 1 12 9 2 3 15 1 9 13 10 9 2
9 9 13 1 12 1 15 0 9 2
29 1 9 13 9 1 12 9 1 10 9 7 1 10 9 15 13 3 2 7 1 10 9 1 15 7 15 1 9 2
20 15 4 13 16 10 0 9 13 1 15 1 9 1 14 1 9 3 3 13 2
9 9 4 4 0 7 10 0 9 2
16 10 0 9 1 9 13 1 9 1 10 9 15 13 1 9 2
14 12 9 9 13 15 15 16 15 4 13 10 9 3 2
15 9 4 3 3 1 3 13 14 13 1 10 9 7 3 2
10 3 0 9 13 3 1 12 0 9 2
4 1 10 0 2
35 3 10 9 13 1 10 9 2 3 15 13 9 1 3 15 4 13 0 9 2 13 15 10 0 9 3 16 15 4 13 0 9 7 9 2
12 2 13 9 1 9 1 9 12 7 12 2 2
4 1 10 0 2
29 10 9 15 13 1 10 9 2 3 15 13 15 1 10 9 2 13 1 10 9 15 13 1 10 0 9 1 9 2
21 15 13 1 9 16 9 4 0 16 15 3 13 0 9 7 10 9 3 1 9 2
10 3 10 9 4 13 1 9 10 9 2
26 1 10 9 9 2 1 12 9 1 10 9 2 13 15 10 2 9 2 1 15 12 0 9 4 13 2
10 15 1 10 0 13 10 9 7 9 2
19 9 1 9 13 1 14 13 15 1 10 12 9 15 4 3 0 7 9 2
25 12 1 10 12 1 10 9 4 1 9 4 13 14 13 1 10 0 9 7 10 9 13 3 3 2
31 1 10 0 12 9 1 10 9 13 15 3 2 7 1 7 1 10 0 13 10 10 0 3 2 7 3 1 10 0 9 2
7 3 13 15 3 10 0 2
9 15 13 15 1 9 1 0 9 2
15 9 1 10 9 15 13 1 9 1 14 1 9 4 0 2
22 1 10 9 15 13 1 9 1 14 4 0 13 15 3 12 15 13 0 9 12 9 2
16 15 1 10 9 15 13 10 9 3 13 3 3 3 0 9 2
16 12 1 9 1 9 7 12 1 9 1 9 13 12 9 15 2
76 1 9 1 10 9 1 9 1 10 0 15 13 0 9 4 15 13 3 15 1 12 9 2 9 15 15 3 13 16 15 13 3 2 9 15 15 13 16 10 0 4 4 13 15 16 3 3 15 4 13 3 1 10 0 9 7 9 15 15 3 4 0 1 16 15 13 0 9 7 15 3 4 13 1 9 2
24 9 1 10 3 0 9 13 15 1 10 0 1 16 15 15 4 13 4 3 0 1 10 9 2
27 1 16 9 1 9 4 3 3 0 1 10 9 15 13 1 15 2 13 9 3 1 0 9 1 0 9 2
28 9 1 0 9 13 1 16 3 10 9 7 9 13 1 9 7 9 1 9 1 10 9 15 15 13 15 1 2
5 10 9 13 1 9
15 3 1 10 9 1 0 13 10 0 9 9 10 0 9 2
18 15 13 1 10 9 1 9 1 9 0 1 10 0 9 15 13 1 2
16 12 9 13 1 0 9 1 12 9 1 12 9 1 10 9 2
22 15 7 15 1 9 13 3 1 0 15 7 3 10 9 3 1 15 7 15 1 15 2
7 9 13 1 12 0 9 2
36 1 9 1 9 15 13 1 9 1 10 9 13 9 1 9 1 9 1 9 2 9 2 9 2 9 2 0 9 2 9 1 0 9 7 9 2
4 0 2 0 2
5 9 4 3 0 2
33 16 12 9 13 3 0 2 0 2 0 2 0 7 0 9 2 13 10 0 9 1 9 3 1 10 9 16 15 13 1 0 9 2
4 9 13 1 9
22 10 9 15 3 3 4 13 13 10 9 15 3 13 1 9 1 10 0 9 0 9 2
19 10 9 2 10 9 2 9 7 9 13 1 0 9 1 10 9 15 13 2
11 9 13 1 9 9 1 9 1 10 9 2
8 9 13 1 9 1 0 9 2
21 10 9 7 9 15 13 1 9 13 1 9 1 9 1 0 9 7 9 1 15 2
20 15 15 4 4 13 13 9 7 9 1 10 9 3 9 15 13 1 0 9 2
13 1 10 9 13 9 1 9 1 10 9 0 9 2
12 3 3 1 9 13 9 9 1 9 1 9 2
25 9 4 10 9 2 10 9 7 9 1 10 0 9 13 10 9 7 9 15 4 13 1 0 9 2
12 3 13 3 10 9 15 4 14 13 3 13 2
30 9 13 1 10 0 9 2 9 2 15 1 10 9 13 9 7 9 15 13 10 9 1 9 7 13 10 9 7 9 2
21 3 13 10 0 0 9 15 13 3 1 10 9 15 1 3 13 15 1 0 9 2
12 15 13 3 9 3 1 10 9 1 10 0 2
11 1 0 0 9 4 15 0 1 10 9 2
20 15 13 3 1 9 2 9 2 9 2 0 7 0 9 2 9 2 9 3 2
13 1 10 0 9 1 15 1 10 9 13 0 9 2
12 0 9 1 9 1 0 9 13 15 3 0 2
17 15 13 3 3 1 15 2 16 15 3 13 10 9 15 13 1 2
19 15 13 15 3 0 16 15 4 13 3 9 1 10 0 1 9 1 11 2
16 15 13 3 16 15 13 16 10 0 3 13 10 9 1 9 2
17 7 15 13 15 3 0 14 0 13 9 1 9 1 11 1 9 2
17 2 15 4 3 9 1 15 2 15 4 9 1 15 1 15 2 2
45 11 2 3 15 13 15 0 2 13 10 3 0 9 2 13 9 7 9 7 9 3 14 13 3 0 3 2 7 1 15 15 13 15 0 4 9 13 3 10 9 1 9 7 9 2
11 15 4 10 9 15 4 0 1 0 9 2
19 12 0 9 2 0 1 9 12 2 4 13 10 0 9 1 10 0 9 2
6 15 4 9 7 9 2
6 10 9 9 4 0 2
14 3 10 9 4 0 7 15 13 3 1 10 0 9 2
18 1 10 3 0 4 12 9 9 7 9 13 1 9 0 0 10 9 2
8 3 13 9 2 9 7 9 2
15 3 13 10 0 9 15 2 10 9 15 3 13 13 9 2
15 9 1 9 2 9 7 9 4 0 1 10 3 0 9 2
26 9 13 1 10 9 3 1 9 15 13 15 3 0 2 1 10 0 0 1 15 15 13 1 0 9 2
14 10 0 9 13 1 10 0 9 7 3 3 1 9 2
10 1 10 0 11 13 9 1 9 9 2
8 10 9 1 9 13 9 3 2
30 3 15 13 3 3 0 9 16 15 3 4 4 13 2 7 3 15 13 3 0 16 15 13 3 3 1 0 0 9 2
18 1 0 9 12 9 2 3 3 10 0 2 13 12 3 12 1 9 2
12 3 10 0 13 1 11 9 2 12 2 9 2
5 3 13 15 15 2
19 10 9 12 12 9 13 10 9 1 10 9 2 15 7 3 10 0 9 2
9 9 13 2 3 3 2 10 9 2
20 10 9 15 13 10 0 9 7 10 9 3 2 3 4 15 13 1 10 9 2
12 2 0 9 1 10 9 1 0 9 4 0 2
47 15 4 3 13 1 2 1 9 2 16 15 1 15 4 14 13 15 1 7 13 15 1 0 9 7 9 16 15 3 4 13 1 10 0 9 1 3 9 7 1 10 9 1 0 9 2 2
3 9 13 2
16 15 15 13 13 3 1 7 1 15 10 9 2 0 13 9 2
46 15 15 13 3 3 3 4 15 15 3 4 13 9 2 3 3 1 10 9 2 3 13 9 2 3 4 0 2 7 10 0 9 4 1 0 9 0 7 3 3 0 16 15 13 9 2
13 15 13 9 1 9 7 4 3 4 13 10 9 2
27 1 9 9 13 15 16 1 15 15 13 3 7 3 12 9 2 9 13 15 3 3 10 9 15 13 9 2
16 15 13 10 9 15 3 4 3 3 0 7 15 13 3 3 2
16 9 4 3 3 10 9 1 14 4 0 1 9 7 0 9 2
45 1 3 0 9 4 15 9 1 14 9 1 13 1 10 0 2 0 2 0 7 3 0 9 7 14 3 4 13 15 3 10 9 2 14 7 9 1 10 0 9 13 9 0 9 2
3 9 13 2
14 9 1 9 9 1 10 0 9 0 9 13 1 9 2
13 3 15 3 13 1 4 9 13 3 7 13 1 2
12 3 13 15 1 10 9 9 1 10 0 9 2
25 3 4 9 0 1 10 0 9 7 10 0 9 3 15 13 9 2 3 9 2 1 14 13 9 2
30 15 13 3 9 7 10 9 16 15 4 0 2 13 15 0 7 4 0 3 16 15 13 0 9 2 3 3 1 9 2
1 9
8 10 0 9 13 1 9 12 2
9 0 9 4 9 13 1 9 12 2
14 3 9 3 4 0 13 15 9 3 14 13 10 9 2
10 15 13 3 9 14 13 14 13 9 2
23 15 4 3 13 1 16 15 13 12 9 1 0 7 0 9 1 10 9 3 15 13 9 2
13 10 0 9 13 9 7 9 13 2 9 13 9 2
5 12 9 1 12 9
13 9 2 9 2 9 2 9 3 13 12 9 12 2
6 9 13 12 9 3 2
21 9 13 3 1 0 9 0 9 1 9 2 16 15 4 0 7 0 14 13 15 2
13 9 4 13 3 0 16 9 3 13 10 9 0 2
43 10 0 7 0 9 9 1 9 13 1 4 14 13 7 13 16 15 3 13 3 1 14 3 13 1 9 2 9 7 0 9 1 0 9 7 9 7 13 9 1 0 9 2
5 1 9 2 1 9
25 15 4 0 14 13 0 9 1 10 0 9 15 4 1 9 1 9 0 2 15 13 0 9 3 2
19 15 13 15 3 3 10 9 7 13 3 1 10 7 0 9 14 13 3 2
13 10 0 9 13 3 0 9 1 9 7 13 9 2
12 15 4 3 0 1 9 14 13 1 0 9 2
17 1 7 1 16 9 13 13 9 3 0 7 9 13 1 9 3 2
6 10 0 2 10 0 9
9 3 0 4 9 3 3 1 9 2
9 15 13 1 3 15 13 9 0 2
23 3 13 9 9 2 1 14 13 7 0 4 15 13 7 13 9 3 2 3 1 10 9 2
30 1 9 9 13 9 2 3 4 9 14 13 1 3 15 15 4 13 9 7 3 13 2 3 16 15 3 4 13 9 2
25 15 1 10 0 9 1 10 0 9 7 9 1 9 1 9 1 9 11 4 3 9 1 0 9 2
8 9 0 13 1 10 0 9 2
10 0 1 11 1 9 1 9 0 2 2
3 0 9 2
15 1 9 9 4 15 3 13 0 9 7 13 9 7 9 2
14 15 4 3 13 0 9 9 1 10 7 9 9 2 2
3 0 9 2
15 10 9 4 3 13 2 13 3 1 10 9 2 10 9 2
14 3 10 0 9 13 3 13 15 3 14 13 7 13 2
16 11 13 13 0 7 0 0 3 2 10 9 7 9 4 0 2
19 1 10 0 9 13 15 1 10 9 1 14 13 9 7 9 0 1 9 2
12 15 13 3 4 0 3 16 9 13 15 3 2
11 3 4 13 0 9 1 9 7 10 9 2
4 15 4 9 2
25 10 0 9 4 3 3 3 15 13 14 13 3 0 15 4 14 1 10 9 13 13 15 9 4 2
11 10 9 1 10 3 9 4 13 4 9 2
15 3 10 9 1 10 0 9 7 9 13 3 10 0 9 2
21 9 4 1 10 0 9 13 1 10 0 0 9 7 3 10 0 9 1 10 9 2
16 9 4 3 9 0 9 1 10 9 15 3 13 10 0 9 2
13 9 4 13 9 2 9 2 9 2 9 2 9 2
20 10 0 9 1 9 13 13 0 12 9 2 2 0 9 2 0 9 2 0 9
12 1 10 12 0 4 3 10 0 10 3 0 2
19 15 13 14 3 3 15 4 0 13 13 16 9 13 7 3 10 0 9 2
19 16 15 1 15 13 7 13 1 9 9 4 10 0 9 3 13 1 9 2
18 10 0 13 3 1 14 13 0 0 9 1 9 2 3 1 10 9 2
33 10 0 4 3 0 10 9 1 10 0 1 16 15 1 10 0 1 10 0 13 9 2 15 4 13 1 14 13 16 0 9 13 2
8 13 3 3 1 9 12 3 2
5 9 1 10 0 9
18 10 9 15 15 4 13 3 4 16 9 7 9 3 4 10 0 0 2
32 3 13 10 9 1 10 0 1 9 3 15 13 14 13 9 2 7 10 0 9 7 10 9 0 9 13 3 10 0 0 9 2
18 9 0 9 13 0 9 1 9 3 2 3 3 1 0 11 7 9 2
17 15 13 0 9 2 1 9 1 11 2 1 10 9 3 1 9 2
16 9 2 9 1 10 0 9 2 4 3 13 10 9 1 9 2
23 10 0 9 9 1 10 0 9 4 3 10 0 7 3 10 9 7 9 1 10 0 9 2
14 11 9 1 9 2 9 12 2 1 11 2 0 9 2
5 9 1 10 0 9
36 3 2 3 15 13 10 0 9 1 11 2 15 13 1 9 2 13 15 9 7 9 15 13 13 10 9 15 13 1 9 1 9 2 9 3 2
13 1 9 7 9 13 10 3 0 9 1 0 9 2
11 9 4 3 3 0 13 10 9 15 13 2
34 10 0 9 13 10 9 1 16 0 0 9 2 3 9 7 3 9 2 13 9 1 9 1 9 7 9 2 1 9 2 9 7 9 2
16 10 0 9 4 1 9 13 7 3 4 3 10 0 9 13 2
21 9 4 13 3 7 13 16 15 4 13 9 1 9 1 10 0 9 1 10 9 2
18 3 1 10 9 4 10 0 7 0 9 1 10 0 9 13 1 9 2
17 7 9 4 3 0 1 10 9 7 15 4 15 3 3 14 13 2
25 3 3 9 1 10 0 9 1 10 0 9 4 13 3 4 10 0 9 9 13 3 0 1 9 2
17 15 4 13 3 16 3 9 3 4 13 0 4 15 13 13 0 2
5 9 1 10 0 9
19 1 9 9 13 15 3 3 3 1 14 13 9 1 10 9 1 10 0 2
11 7 9 1 9 7 9 9 4 4 13 2
24 10 9 4 13 9 7 9 14 13 3 1 1 9 3 1 10 9 2 3 10 9 7 9 2
25 15 7 15 4 13 9 1 14 13 10 9 1 9 7 1 14 13 1 0 7 0 9 1 15 2
28 1 10 9 13 10 0 9 1 9 7 10 9 1 9 2 3 9 2 7 10 3 0 9 1 10 0 9 2
43 1 10 3 0 0 9 1 11 13 15 3 3 15 4 3 7 3 0 1 14 13 13 10 0 2 0 9 7 9 3 1 9 7 9 1 10 0 9 1 9 7 9 2
29 15 4 10 0 9 2 7 15 4 13 3 16 9 9 1 0 9 7 3 13 15 1 10 9 7 0 9 9 2
10 10 0 0 9 13 3 1 10 9 2
18 10 0 0 9 13 3 10 0 9 1 9 2 9 2 9 7 9 2
25 10 9 4 3 13 1 0 9 1 16 10 0 9 1 9 4 4 13 3 10 9 7 0 9 2
5 9 2 9 7 9
47 3 3 9 3 4 3 0 7 3 7 15 3 4 0 9 1 10 0 7 0 9 1 10 9 13 3 10 0 3 1 9 1 9 7 3 3 3 10 9 1 9 7 9 13 3 3 2
12 10 0 9 13 3 1 10 9 1 9 9 2
10 1 9 13 3 0 9 9 1 9 2
18 1 12 9 3 13 15 3 7 12 9 1 9 9 7 10 0 9 2
9 3 13 10 9 3 1 12 9 2
16 3 13 10 0 9 2 9 2 0 9 7 1 9 7 9 2
11 3 0 9 1 10 0 9 4 9 13 2
25 10 9 15 9 3 3 7 0 0 13 1 9 4 3 10 9 15 13 3 10 0 9 1 9 2
22 15 4 10 9 15 13 9 1 9 10 9 2 3 1 15 15 3 13 3 10 9 2
19 3 1 10 9 13 15 1 10 0 9 15 13 1 14 13 1 10 9 2
40 15 13 16 3 16 9 4 4 9 1 9 9 3 4 15 1 10 9 4 10 0 9 1 16 9 13 10 0 9 15 3 3 3 13 15 1 9 1 9 2
12 15 13 0 0 9 14 3 13 10 0 9 2
15 3 4 3 9 2 9 2 9 2 9 7 0 9 13 2
30 1 11 11 9 11 2 15 13 1 9 1 9 12 2 4 0 11 13 9 1 15 0 0 16 9 13 1 10 9 2
10 3 9 13 2 13 15 1 10 9 2
28 2 3 15 3 13 3 13 15 3 16 15 4 13 14 13 10 9 2 13 10 9 1 10 9 1 9 11 2
22 10 12 0 9 11 7 11 13 16 9 1 2 10 0 2 9 4 13 1 12 9 2
12 10 0 9 4 9 7 9 2 13 9 3 2
10 15 13 16 9 13 0 9 7 9 2
17 1 9 2 15 4 0 9 1 9 2 13 9 0 9 7 9 2
10 10 0 9 13 9 15 9 9 13 2
10 10 9 13 3 3 1 0 7 0 2
11 15 15 13 10 0 9 13 3 1 9 2
11 1 11 7 11 13 15 9 15 13 9 2
20 15 13 9 3 2 15 13 1 10 0 9 2 15 13 9 2 13 7 13 2
8 10 0 9 13 3 1 9 2
12 15 13 15 15 13 1 10 0 9 1 9 2
16 15 13 9 0 9 2 15 13 15 2 15 13 1 15 3 2
13 13 9 2 15 3 13 9 9 1 10 0 9 2
3 9 1 9
25 3 9 13 1 9 4 15 13 1 1 11 11 7 11 11 9 2 12 9 2 2 11 12 2 2
11 1 9 4 9 1 10 9 13 1 9 2
22 10 9 13 0 2 10 7 10 9 2 9 16 15 4 1 0 9 1 10 9 2 2
6 3 13 9 1 9 2
10 9 13 1 10 9 11 7 11 9 2
11 0 9 13 16 0 9 4 0 7 0 2
8 3 9 4 13 15 1 9 2
12 15 13 15 14 13 10 9 15 13 3 3 2
10 2 15 15 13 3 3 1 15 2 2
4 9 13 3 2
11 9 13 16 9 3 7 9 13 9 9 2
10 15 4 3 0 3 15 13 15 3 2
14 15 4 1 0 4 0 14 13 3 9 13 1 9 2
16 15 4 13 16 11 2 11 9 1 0 9 13 11 7 11 2
12 10 0 9 4 3 13 7 3 0 7 0 2
19 1 9 2 4 15 13 2 13 0 9 3 3 3 15 13 9 1 9 2
9 10 3 0 9 4 3 1 9 2
21 10 0 0 9 2 11 11 11 2 13 1 10 0 9 7 9 2 9 9 2 2
18 1 15 2 13 15 2 13 9 3 3 7 1 15 15 13 0 9 2
12 10 1 9 15 3 13 10 0 9 13 3 2
16 3 13 15 3 0 9 15 13 3 9 7 9 9 1 15 2
6 3 9 9 4 0 2
6 15 4 3 3 9 2
10 1 10 0 9 4 15 13 1 9 2
4 10 9 1 9
16 11 4 13 7 9 2 15 13 10 3 0 9 1 9 9 2
13 11 2 11 4 13 14 13 10 9 1 0 9 2
11 15 13 1 9 9 1 10 12 0 9 2
7 10 0 9 0 1 10 9
17 15 4 1 11 2 11 10 9 15 1 0 9 13 13 1 9 2
7 3 3 13 15 9 9 2
29 2 9 13 10 9 7 10 9 1 10 0 9 9 2 10 0 0 0 9 15 3 3 4 4 13 1 10 0 2
35 2 3 4 15 4 13 3 2 3 15 13 7 0 9 1 11 1 11 7 11 7 10 0 13 7 13 9 7 13 1 1 9 2 2 2
28 9 4 3 3 9 2 3 15 13 10 9 7 10 9 9 1 0 9 1 14 13 0 9 7 13 3 3 2
18 15 1 9 13 1 10 9 1 9 2 15 13 3 7 13 15 3 2
17 15 13 3 10 0 9 13 2 9 7 15 4 3 15 1 15 2
33 16 9 4 15 15 4 13 10 0 9 2 13 15 2 16 15 3 13 16 15 3 3 4 3 3 1 10 9 3 1 10 9 2
8 9 13 3 3 3 3 3 2
20 15 13 3 16 9 4 13 9 1 9 1 10 0 9 3 7 1 9 2 2
8 2 12 9 2 9 12 2 2
2 9 9
7 10 9 13 1 9 12 2
9 9 1 9 7 9 4 3 0 2
9 2 9 4 0 7 3 0 9 2
17 9 4 9 1 0 0 9 2 3 3 3 0 9 16 9 13 2
25 9 1 10 9 13 16 15 4 0 1 10 9 7 13 3 0 9 1 1 9 2 3 1 9 2
26 16 15 4 13 10 9 3 4 0 2 10 9 4 15 3 13 15 3 16 9 13 15 3 1 9 2
12 10 0 1 9 4 3 3 13 3 0 9 2
17 7 15 13 3 1 16 15 4 4 13 10 2 0 9 2 2 2
8 2 12 9 2 9 12 2 2
1 9
15 15 4 10 9 15 13 1 9 1 11 2 9 9 2 2
10 11 2 11 13 15 1 10 12 9 2
9 3 13 15 9 1 10 0 9 2
5 3 13 10 9 2
22 2 1 9 12 4 15 13 9 1 0 9 1 3 0 9 2 7 15 0 0 9 2
8 15 4 3 3 4 10 9 2
13 15 4 13 0 9 2 1 0 9 13 10 0 2
26 15 1 10 12 9 4 13 1 7 9 7 9 7 13 9 14 13 15 3 3 12 9 3 7 0 2
6 9 9 4 3 13 2
7 10 0 4 4 10 9 2
13 7 3 13 15 16 10 9 13 10 0 1 15 2
10 3 4 9 0 7 15 13 10 9 2
4 15 13 3 2
19 7 10 9 1 9 4 15 13 9 2 3 15 13 1 10 0 0 9 2
12 15 13 1 9 3 3 3 1 14 13 9 2
9 10 12 9 1 9 13 0 9 2
11 9 4 10 0 0 9 1 9 7 9 2
13 13 4 3 3 3 0 2 15 13 9 3 3 2
7 7 3 4 10 9 0 2
9 0 7 3 13 15 3 3 3 2
19 9 1 9 13 3 10 0 9 3 1 9 2 3 1 10 0 2 2 2
8 2 12 9 2 9 12 2 2
1 9
17 3 3 9 13 1 1 9 13 1 1 10 9 9 13 1 9 2
13 9 13 1 10 9 0 9 12 1 9 11 11 2
12 2 12 9 1 9 2 9 13 2 12 2 2
14 9 0 9 13 9 2 3 4 15 10 0 9 2 2
11 1 12 9 1 9 13 15 1 1 15 2
10 15 1 10 3 0 9 13 1 9 2
15 9 9 4 3 13 0 2 3 9 1 9 13 1 9 2
24 10 12 0 9 13 3 9 2 12 9 2 2 9 2 12 9 2 7 9 2 12 9 2 2
11 15 4 3 3 1 9 1 10 0 9 2
10 11 11 9 4 3 10 9 9 0 2
19 15 4 13 16 15 3 7 3 1 10 0 9 13 10 3 3 0 9 2
2 0 9
18 9 1 10 0 9 1 10 9 13 3 1 9 1 0 9 7 9 2
22 9 7 9 2 9 2 9 7 9 4 9 1 0 0 7 3 0 9 1 0 9 2
23 1 9 13 15 9 1 10 3 0 9 1 0 9 1 9 2 9 12 2 9 12 2 2
33 1 0 9 13 15 3 3 9 2 9 1 9 3 1 0 9 2 3 3 15 13 9 15 1 0 13 0 2 3 3 13 9 2
23 15 1 9 1 10 0 9 13 16 9 4 13 3 15 7 16 10 9 4 13 1 15 2
17 0 9 13 10 9 9 0 9 1 12 0 2 9 2 1 9 2
16 9 13 10 9 2 13 15 1 9 7 13 10 9 1 9 2
12 9 15 13 3 13 1 9 15 13 1 9 2
6 9 13 10 0 9 2
13 3 13 9 0 9 1 10 0 9 9 1 9 2
13 9 1 0 9 2 9 2 15 13 3 1 9 2
23 1 10 9 3 7 3 13 9 10 0 9 1 9 7 13 1 9 7 9 9 1 15 2
19 9 1 14 13 3 0 9 3 15 4 0 13 1 0 9 1 9 9 2
23 1 0 9 2 7 9 7 9 2 15 13 0 9 2 13 1 9 9 3 3 1 9 2
10 15 13 9 1 9 2 3 9 13 2
10 1 10 9 13 15 3 9 0 9 2
25 3 13 9 9 1 10 0 9 2 9 7 9 9 1 9 10 1 15 3 0 9 1 0 9 2
27 9 0 9 2 9 1 9 7 9 1 9 13 3 10 0 9 1 9 2 10 0 9 13 1 0 9 2
13 9 1 10 0 9 4 3 10 0 9 1 9 2
14 1 9 4 10 0 9 2 9 2 13 1 0 9 2
15 10 9 4 9 2 3 9 1 0 9 13 1 9 9 2
7 0 9 13 9 1 9 2
21 0 9 4 3 13 1 9 1 0 9 2 3 1 9 1 9 2 9 12 2 2
12 0 9 4 9 9 2 9 9 7 9 9 2
10 0 9 2 3 9 2 13 0 9 2
14 1 10 0 0 9 13 0 9 1 10 0 9 9 2
8 0 9 13 15 1 0 9 2
9 9 4 3 13 1 9 7 9 2
20 16 10 9 1 10 9 13 2 13 9 1 9 10 9 1 10 0 1 9 2
16 9 9 1 9 1 9 1 9 4 3 10 9 1 0 9 2
18 13 10 9 0 9 10 9 15 13 15 2 13 15 10 3 0 9 2
21 9 1 16 9 13 1 9 4 3 3 0 16 15 13 15 3 1 10 0 9 2
3 9 1 9
15 1 9 4 10 9 9 0 1 9 1 12 9 1 10 2
11 9 9 4 1 0 9 13 1 0 9 2
16 1 10 9 1 0 9 7 9 13 3 9 1 10 9 0 2
17 1 9 13 3 9 13 1 10 0 9 1 10 9 7 10 9 2
16 9 13 10 9 1 9 2 7 15 13 3 3 0 1 9 2
10 1 9 13 3 9 1 9 1 9 2
8 1 9 13 3 9 1 9 2
16 9 13 9 7 9 1 9 9 1 9 1 10 9 1 9 2
8 9 9 1 9 4 3 13 2
13 9 7 9 13 10 9 1 9 2 9 12 2 2
18 1 9 1 0 9 2 3 9 2 13 0 9 3 9 9 1 9 2
19 9 1 0 9 13 3 10 9 1 14 1 9 13 1 10 9 1 9 2
13 15 13 15 1 10 0 9 7 13 15 1 9 2
23 9 15 4 0 1 0 9 2 3 10 0 9 2 4 13 9 1 3 3 1 12 9 2
9 10 9 13 3 1 9 1 9 2
30 15 13 3 3 2 9 2 2 3 9 2 15 3 13 9 1 3 12 9 9 7 1 10 9 1 3 12 1 9 2
11 9 1 10 0 9 13 1 9 1 9 2
14 0 9 13 1 16 10 0 9 13 9 1 9 9 2
14 3 13 15 3 7 10 9 1 9 2 3 1 9 2
14 10 9 13 1 9 2 3 9 4 0 7 9 0 2
11 1 0 9 13 9 7 9 9 1 9 2
11 0 9 13 1 9 7 9 3 0 9 2
14 9 13 3 0 7 0 9 2 15 4 0 1 9 2
9 0 9 9 13 1 9 12 9 2
5 9 9 13 9 2
9 10 9 13 9 3 1 12 9 2
10 9 1 10 9 9 4 3 3 13 2
16 10 3 9 1 9 13 9 1 9 1 9 1 10 0 9 2
20 13 9 0 9 7 9 2 1 9 1 3 9 2 1 9 9 2 13 9 2
13 13 15 0 9 2 3 9 7 9 2 13 9 2
3 9 7 9
17 0 9 9 1 9 1 9 2 9 7 9 1 9 4 13 3 2
14 9 9 7 9 4 13 7 10 9 2 9 12 2 2
14 0 9 1 9 9 1 0 9 4 13 1 11 11 2
21 1 9 13 9 1 9 2 10 9 3 13 1 9 1 12 7 10 9 0 9 2
15 16 10 9 13 13 1 10 9 2 13 3 0 9 15 2
11 15 13 10 0 6 2 7 0 9 13 2
12 1 9 13 9 3 15 13 9 15 13 9 2
11 1 7 1 9 7 9 13 9 0 9 2
9 3 1 9 13 9 1 9 0 2
19 3 1 0 9 2 15 13 1 0 9 2 13 9 3 0 9 1 9 2
21 1 10 0 9 13 9 3 2 0 2 9 2 3 0 9 7 9 13 1 9 2
20 16 9 13 2 13 9 7 9 3 2 7 0 9 13 3 1 9 1 9 2
28 10 0 9 1 9 13 16 9 13 1 10 0 9 9 2 1 15 9 13 1 14 13 9 2 9 12 2 2
28 1 9 1 9 4 15 13 16 9 4 10 3 9 2 10 9 4 10 0 9 15 9 0 9 4 0 1 2
21 10 9 1 0 9 13 12 9 3 0 9 1 9 7 10 0 9 1 0 9 2
19 15 13 15 3 2 16 0 9 1 9 13 3 0 9 7 10 0 9 2
12 9 1 9 1 9 1 0 9 7 1 9 2
14 9 9 13 9 9 15 13 1 10 0 9 1 9 2
15 1 9 9 13 9 3 7 13 1 15 1 9 7 9 2
9 9 7 9 13 1 9 1 9 2
14 13 0 9 3 7 13 2 13 9 3 1 0 9 2
15 9 3 1 9 13 1 9 1 10 0 9 1 9 9 2
13 9 1 9 4 1 9 1 9 1 9 3 0 2
19 9 1 9 13 9 7 9 1 9 2 13 9 2 13 9 1 9 3 2
11 9 13 1 9 1 9 1 10 0 9 2
10 1 9 4 9 4 0 1 0 9 2
6 10 0 9 1 0 9
13 9 1 9 1 10 9 13 15 1 10 0 9 2
15 15 13 7 9 2 9 1 9 7 9 1 9 1 9 2
19 9 1 9 2 9 2 1 10 0 9 13 3 0 2 0 7 0 9 2
13 3 0 9 1 0 9 13 4 1 0 9 0 2
27 7 9 14 13 7 13 9 13 1 9 1 9 7 4 3 9 1 10 9 1 10 9 7 0 0 9 2
13 1 9 4 9 1 9 7 0 9 13 1 9 2
19 1 0 9 7 1 9 1 9 13 9 0 9 14 13 7 10 0 9 2
20 0 9 13 3 0 9 7 15 15 13 1 9 7 13 3 3 9 1 9 2
21 1 10 9 13 9 15 1 9 2 7 9 1 15 13 10 9 16 9 9 13 2
10 3 1 10 9 13 3 9 1 9 2
12 12 9 13 10 0 9 14 13 9 1 9 2
11 9 15 13 10 9 9 1 9 7 9 2
22 0 9 1 9 13 1 9 2 3 15 13 0 9 0 1 3 9 2 3 1 9 2
8 10 9 13 1 9 1 9 2
9 9 13 3 9 1 10 0 9 2
9 10 0 9 13 0 9 1 15 2
20 10 0 9 1 9 4 3 3 0 7 1 9 2 7 9 4 3 3 0 2
33 1 0 9 2 15 1 0 3 13 12 9 1 10 9 2 4 15 1 9 1 9 1 9 4 13 10 0 9 3 1 0 9 2
9 9 4 15 1 10 3 0 9 2
22 15 13 1 10 0 0 9 1 9 7 10 9 2 15 13 1 9 2 9 7 9 2
15 10 0 9 7 9 1 9 13 1 10 0 9 1 9 2
8 9 9 13 9 9 7 9 2
15 9 13 3 1 0 9 1 9 1 9 1 9 7 9 2
31 1 0 9 4 10 0 9 1 9 13 2 3 9 9 1 0 9 7 10 0 1 9 3 2 9 12 2 9 12 2 2
16 10 9 13 7 0 10 0 9 2 9 2 9 2 9 3 2
23 0 9 7 9 1 9 13 3 7 1 15 1 0 9 1 0 9 7 13 3 7 3 2
26 1 0 9 4 10 0 2 0 9 4 10 9 2 16 9 9 4 3 0 7 9 4 10 0 9 2
7 9 1 9 13 3 0 2
18 1 0 0 9 7 3 3 1 9 4 0 9 1 9 13 1 9 2
16 15 13 10 9 0 9 1 9 1 9 1 0 2 0 9 2
10 1 9 13 3 10 0 9 1 9 2
16 1 10 0 9 4 10 0 9 1 0 9 13 10 0 9 2
17 1 10 9 4 0 9 7 9 13 7 13 1 0 9 1 9 2
24 9 1 3 15 13 7 3 10 0 9 13 1 3 9 2 4 3 0 7 0 9 7 0 2
25 1 9 9 7 9 4 10 0 9 10 0 9 2 7 3 9 1 9 1 10 9 13 0 9 2
20 9 13 15 13 0 9 1 9 7 4 3 3 13 1 10 0 9 1 9 2
19 7 16 9 13 3 0 2 4 15 13 10 0 9 1 9 1 0 9 2
19 9 0 9 13 1 9 3 10 0 13 1 0 9 16 10 0 13 9 2
10 9 13 3 3 9 7 13 3 9 2
13 0 9 2 3 9 2 13 15 3 3 1 9 2
12 0 9 1 9 1 9 1 9 2 3 9 2
22 1 9 13 2 3 3 13 2 3 10 0 9 1 9 1 10 3 7 3 0 9 2
13 3 3 10 9 13 2 13 9 7 9 1 9 2
19 15 4 3 10 9 3 10 9 1 10 3 0 9 1 9 4 3 0 2
23 9 1 0 9 13 3 0 9 1 9 9 1 9 7 13 15 15 1 0 9 13 9 2
25 15 13 16 12 9 1 9 1 14 13 1 10 9 13 1 10 10 9 1 9 2 3 9 13 2
12 0 9 4 13 10 9 1 9 1 0 9 2
19 1 9 1 9 13 9 1 0 9 1 9 2 9 12 2 9 12 2 2
22 9 1 0 0 9 4 3 10 9 1 9 7 4 13 0 9 1 9 1 0 9 2
42 1 10 3 9 2 9 11 2 1 0 9 1 9 2 13 9 1 9 9 10 9 1 9 7 13 3 10 9 1 9 1 3 0 9 2 15 13 10 3 0 9 2
12 1 9 13 9 9 10 0 9 1 0 9 2
13 1 0 0 9 7 9 13 0 9 1 3 9 2
8 10 0 9 13 9 1 9 2
13 1 9 1 10 3 0 9 13 15 9 1 15 2
10 9 1 10 9 13 1 9 1 9 2
14 9 13 3 1 10 9 9 13 3 7 3 1 9 2
8 1 0 9 13 3 0 9 2
17 9 13 7 13 1 10 0 9 9 2 9 13 1 15 1 15 2
16 10 0 9 1 9 4 3 0 1 10 1 10 9 0 9 2
2 14 13
15 13 0 9 9 1 9 1 9 2 9 2 9 7 9 2
7 3 13 9 1 0 9 2
6 13 9 7 0 9 2
13 13 9 1 3 9 1 0 9 9 13 10 9 2
10 13 7 13 0 7 0 9 1 9 2
8 13 0 7 0 9 1 9 2
5 15 13 9 9 2
5 15 4 3 9 2
10 13 9 1 0 9 7 13 13 9 2
8 15 13 9 2 0 9 2 2
5 13 9 0 9 2
6 13 9 9 7 9 2
15 13 10 9 1 16 9 4 13 9 1 9 1 0 9 2
19 15 4 3 13 9 1 0 9 7 13 13 1 10 0 9 1 9 9 2
17 7 15 4 13 10 0 9 1 9 7 10 9 3 1 0 9 2
20 15 13 1 10 9 0 0 9 1 9 2 15 15 13 10 0 9 7 9 2
296 15 4 13 1 2 9 3 9 2 9 2 13 9 2 9 7 9 13 1 9 10 9 1 10 9 9 9 13 2 9 3 10 9 2 10 9 13 9 2 1 0 9 13 9 1 9 2 15 4 0 1 0 9 1 10 9 2 1 0 9 3 1 9 9 2 13 9 9 1 9 2 1 15 13 0 9 2 10 0 9 2 15 13 15 3 3 1 9 9 2 3 1 10 0 9 1 11 2 1 10 9 4 3 13 10 0 9 2 3 9 1 11 2 1 10 0 9 1 9 1 9 2 9 7 9 7 1 0 9 2 15 13 9 1 9 2 1 11 13 15 10 0 9 1 3 11 2 11 2 11 2 11 2 11 7 1 10 9 7 11 2 9 2 10 0 9 4 0 1 9 2 10 0 9 4 9 7 9 0 9 2 11 9 4 1 10 9 10 9 1 10 9 0 9 2 9 2 3 13 15 1 10 0 9 7 9 7 9 2 3 4 15 3 7 3 10 9 1 9 2 9 2 1 10 9 13 9 7 9 3 9 0 9 2 1 0 9 4 10 0 9 13 3 1 10 0 9 2 15 3 1 11 7 11 2 9 2 1 0 9 4 10 0 9 9 13 1 0 9 2 3 1 11 2 9 2 3 11 11 13 10 0 9 1 9 13 15 13 9 1 1 0 9 0 9 2
20 0 9 13 3 7 1 11 2 11 2 11 7 11 7 3 1 10 0 9 2
14 1 9 13 0 9 2 11 2 11 2 11 2 11 2
1 9
10 13 1 9 1 10 9 10 0 9 2
6 1 10 9 13 15 2
8 7 4 0 9 13 10 9 2
12 4 15 13 1 12 9 1 9 1 10 0 2
8 13 9 7 0 9 7 9 2
15 9 2 0 15 13 1 9 2 4 4 13 1 0 9 2
37 3 11 7 11 0 13 10 0 11 9 13 15 14 13 9 1 9 2 1 0 9 2 0 9 2 9 2 9 2 9 7 0 9 1 9 9 2
56 9 4 13 16 10 9 13 9 1 0 7 0 9 2 13 10 0 0 9 9 2 13 0 9 2 15 13 0 9 7 14 13 10 0 9 7 15 4 0 2 0 2 13 9 0 1 0 2 0 9 2 1 9 1 9 2
1 9
12 13 0 9 1 3 10 9 0 9 4 13 2
11 3 13 15 10 0 9 1 10 0 9 2
17 13 15 10 9 7 4 15 3 0 2 0 9 2 3 3 9 2
36 10 0 9 2 1 10 0 9 1 9 2 4 10 9 3 3 1 9 7 3 1 10 0 9 2 15 13 9 7 13 9 1 10 0 9 2
21 3 1 9 13 9 11 11 13 1 14 13 9 9 1 10 9 1 9 7 9 2
18 13 1 10 0 9 2 16 15 4 13 9 1 0 10 9 1 9 2
13 1 9 13 9 7 9 10 0 9 1 10 9 2
12 9 0 9 13 3 10 9 1 9 1 9 2
23 7 9 13 1 0 9 2 7 9 7 9 4 3 3 1 9 0 1 10 0 0 9 2
28 3 9 1 9 9 13 10 0 9 2 3 9 13 3 1 9 2 13 9 1 2 9 2 1 9 3 0 2
21 15 13 1 0 12 9 2 10 0 9 7 9 1 0 9 7 9 1 10 0 2
23 1 9 4 11 4 0 2 7 10 0 9 0 9 2 0 9 7 0 9 4 13 15 2
15 9 4 4 10 3 0 9 7 13 9 1 10 0 9 2
29 3 10 0 9 13 13 1 9 9 13 15 9 1 0 10 9 2 0 9 1 0 11 12 2 11 1 11 12 2
13 1 10 0 9 4 10 0 9 14 13 0 9 2
22 15 13 3 10 0 9 2 15 7 10 0 9 4 14 13 0 9 1 10 0 9 2
9 1 9 4 10 0 9 13 3 2
21 0 9 1 9 2 9 2 9 7 9 13 15 7 9 1 9 7 13 3 9 2
8 15 13 10 0 9 7 9 2
20 15 13 1 9 9 7 9 2 10 0 9 4 0 1 0 9 7 0 9 2
1 9
9 13 9 7 9 1 10 0 9 2
7 10 9 13 1 10 9 2
5 3 4 15 13 2
9 3 4 15 0 4 13 15 0 2
26 3 12 13 15 1 11 10 9 1 9 1 9 1 9 7 9 2 9 7 0 9 2 9 7 9 2
21 7 15 13 1 10 9 16 15 13 10 9 1 10 9 2 10 9 1 10 9 2
26 3 1 9 13 15 1 11 13 9 1 0 9 1 9 2 1 9 7 9 2 1 9 7 1 9 2
7 9 1 9 1 11 12 2
7 15 13 10 9 1 9 2
7 13 1 9 9 12 3 2
1 9
10 13 3 10 9 13 1 10 0 9 2
18 13 16 0 10 9 1 9 7 13 13 10 9 1 15 15 13 3 2
1 9
6 9 13 1 9 9 2
20 0 9 4 9 15 13 3 1 16 9 13 1 0 9 2 1 9 7 9 2
16 10 0 9 2 9 2 13 9 7 9 3 1 9 7 9 2
10 1 10 9 13 15 0 9 2 9 2
23 10 0 9 1 9 4 0 2 15 15 3 13 3 1 0 9 2 1 0 9 0 9 2
43 7 1 9 13 15 3 3 10 9 1 9 1 9 7 9 15 4 3 0 1 0 9 7 3 10 0 9 9 7 9 13 1 0 9 1 9 2 1 9 7 1 9 2
8 10 0 1 10 9 4 0 2
11 0 9 4 13 9 7 9 3 0 9 2
14 3 13 3 9 10 3 0 9 2 3 13 15 9 2
11 9 4 10 1 11 1 9 3 0 9 2
23 9 4 16 15 13 1 10 9 2 3 9 1 0 9 1 9 7 9 13 1 14 13 2
21 1 3 3 3 4 15 0 2 16 9 7 9 13 1 0 9 7 13 0 9 2
11 3 13 15 1 10 9 7 13 10 9 2
12 13 15 16 9 7 9 13 10 9 14 13 2
9 13 9 16 9 1 9 4 13 2
28 4 9 7 9 1 9 13 9 3 2 3 16 3 7 3 9 13 9 1 9 2 9 9 1 9 7 9 2
40 1 0 9 13 15 15 3 0 2 16 15 1 0 9 4 9 9 14 3 13 9 7 13 7 16 3 9 13 1 9 14 13 1 16 9 4 13 15 15 2
29 15 13 2 3 0 9 4 13 1 9 2 7 13 2 16 9 13 3 0 9 7 9 14 13 1 9 7 9 2
12 1 9 4 0 9 4 14 13 7 3 0 2
13 16 9 13 15 1 2 9 2 4 3 3 0 2
14 4 9 1 9 0 9 7 9 2 13 9 12 2 2
34 4 15 9 1 0 7 0 2 3 15 13 2 3 9 1 9 7 9 4 13 1 9 2 16 1 9 0 9 4 13 9 1 9 2
20 1 0 9 13 9 13 9 2 13 15 15 4 0 3 7 15 15 4 0 2
47 7 9 1 3 0 7 0 4 13 3 2 16 15 3 13 3 16 10 9 15 13 9 13 16 15 3 13 10 9 7 9 14 13 2 14 13 10 9 1 10 9 2 14 13 10 9 2
13 3 13 15 9 1 0 9 2 13 9 12 2 2
1 9
29 16 9 7 9 13 9 7 13 9 4 3 13 7 13 1 10 0 3 7 10 0 7 0 9 1 9 1 9 2
11 7 9 4 1 0 9 13 3 0 9 2
20 1 9 13 2 16 15 1 10 0 11 3 4 0 16 10 9 13 0 9 2
6 10 0 9 13 9 2
16 15 4 13 10 0 9 1 9 2 15 13 15 1 0 9 2
19 7 15 4 3 13 10 0 9 1 15 2 15 13 0 14 13 0 9 2
14 0 4 9 1 10 9 1 0 9 7 1 0 9 2
18 7 9 2 15 13 3 3 3 2 13 16 9 13 3 0 7 0 2
11 14 13 0 9 13 10 9 1 10 0 2
27 10 0 9 1 10 9 4 2 16 9 13 16 9 13 0 9 7 9 2 15 13 0 9 1 10 9 2
28 15 4 3 13 2 16 15 1 10 0 9 4 0 1 9 14 13 10 9 10 9 2 10 9 2 10 9 2
17 9 13 1 10 0 9 2 9 2 9 2 9 2 13 1 9 2
13 16 10 9 13 0 0 9 2 9 2 4 0 2
9 9 7 9 4 0 9 1 9 2
13 0 4 3 9 2 12 9 7 12 9 13 3 2
17 16 1 0 9 9 13 2 4 1 0 9 9 10 0 0 9 2
35 16 10 9 7 10 9 3 4 13 2 10 9 2 7 16 10 9 13 0 9 1 15 4 4 10 0 9 9 1 9 7 9 1 9 2
19 7 0 7 0 9 13 2 16 9 4 10 0 9 3 1 10 0 9 2
15 10 0 9 13 3 0 9 2 15 13 16 10 9 13 2
18 16 9 4 0 13 2 16 9 1 15 15 13 9 4 0 14 13 2
11 10 0 9 4 16 15 3 13 10 9 2
22 13 9 15 0 1 15 15 3 13 9 14 13 1 10 0 0 9 14 13 0 9 2
12 1 9 13 7 11 7 11 3 10 0 9 2
30 1 0 0 9 13 15 2 16 15 4 13 10 0 9 1 10 9 1 9 1 9 7 9 2 3 15 4 13 0 2
36 1 15 13 2 16 3 16 9 4 13 0 9 2 4 0 9 13 2 3 3 3 10 9 7 10 9 4 13 9 1 14 4 13 1 15 2
14 15 1 10 0 9 0 9 13 1 0 9 7 9 2
29 1 0 9 9 13 15 15 15 13 3 9 2 15 13 9 9 3 2 15 13 0 9 2 15 13 3 1 9 2
41 9 4 1 9 3 0 2 3 3 1 16 9 3 4 13 0 9 1 14 13 9 1 9 9 7 3 1 16 0 9 2 3 3 0 9 2 13 3 1 9 2
23 10 9 9 13 10 2 9 2 2 10 9 15 3 4 0 1 9 3 1 11 7 11 2
17 1 10 0 9 13 9 3 1 9 7 3 1 9 1 9 9 2
32 3 4 3 10 0 9 7 9 4 14 13 3 2 15 3 13 16 9 9 13 3 1 9 1 9 7 1 9 1 0 9 2
12 9 4 3 13 9 2 3 15 3 3 13 2
36 3 13 3 10 0 10 0 9 1 14 13 3 1 10 9 2 3 15 13 14 13 9 1 0 9 2 1 9 2 1 9 2 1 9 3 2
2 0 9
23 15 4 3 3 13 13 2 16 15 3 13 10 0 9 15 13 9 7 9 3 1 9 2
19 15 13 16 10 0 9 2 10 0 9 2 4 15 15 3 13 3 15 2
12 10 0 9 15 13 1 9 4 10 0 9 2
24 15 13 15 15 13 2 16 3 0 9 13 13 9 7 3 15 4 13 2 4 3 9 13 2
25 1 10 0 9 0 9 4 15 10 9 2 16 9 13 15 4 13 9 7 13 9 1 10 9 2
16 9 13 3 1 16 10 9 7 10 9 13 13 9 1 9 2
10 9 13 10 9 1 16 9 3 13 2
17 0 4 9 2 16 10 9 7 10 9 13 3 1 14 13 9 2
18 16 9 1 9 13 3 1 9 2 13 0 9 3 9 7 0 9 2
14 0 9 13 3 1 9 3 3 14 13 9 1 9 2
17 15 4 3 1 15 0 9 1 0 9 1 10 9 7 10 9 2
8 15 13 3 9 1 10 0 2
15 9 14 13 9 1 10 9 4 1 10 9 13 1 9 2
31 3 16 15 3 13 9 2 15 3 4 13 2 16 10 9 3 13 9 1 9 2 4 15 3 13 9 1 9 3 0 2
20 3 13 9 2 16 0 9 1 9 4 3 0 7 3 2 1 10 0 9 2
12 1 9 13 15 9 1 0 9 1 10 9 2
15 15 13 15 15 13 16 10 0 9 1 9 4 3 0 2
39 15 13 3 15 15 13 2 16 10 0 0 9 4 13 1 10 0 9 7 1 0 0 9 2 15 13 3 2 15 13 3 2 15 13 3 1 0 9 2
9 3 13 15 16 15 3 13 3 2
16 15 13 3 10 0 9 1 14 13 9 7 14 13 0 9 2
27 10 9 4 2 16 15 4 3 0 14 13 0 9 1 10 9 7 16 10 9 3 4 4 0 1 9 2
25 10 9 1 10 9 4 16 9 13 2 16 9 13 3 3 1 15 16 9 7 9 13 3 0 2
12 1 10 0 9 13 0 9 1 10 0 9 2
17 4 10 9 4 13 15 1 9 2 4 9 13 2 3 1 9 2
14 4 9 13 1 10 9 1 9 1 9 3 1 9 2
23 12 9 13 13 2 12 9 3 1 9 2 12 0 9 1 9 2 12 9 3 1 9 2
11 10 12 9 13 2 15 13 15 3 9 2
1 9
10 1 0 9 4 9 13 3 7 3 2
15 10 9 4 13 3 3 9 13 7 9 13 3 3 0 2
8 1 11 4 10 9 3 0 2
35 1 9 4 1 9 9 9 2 9 15 13 1 9 9 2 13 1 3 12 2 12 2 1 3 12 2 12 2 2 3 1 3 12 9 2
6 9 13 9 2 9 2
18 9 0 9 1 12 7 0 9 4 3 1 0 9 13 1 0 9 2
28 15 13 1 10 0 9 15 13 1 9 1 9 2 10 0 9 2 9 9 7 9 1 10 0 9 1 9 2
20 9 13 1 10 0 9 2 7 3 9 2 9 2 9 2 9 2 4 13 2
7 15 13 9 1 9 9 2
14 9 4 3 13 15 9 1 10 9 1 10 0 9 2
12 15 13 3 3 0 10 2 0 2 9 4 2
17 3 13 15 3 3 1 10 9 9 9 13 1 0 9 1 9 2
15 3 13 15 3 1 3 0 10 9 1 0 7 0 9 2
10 9 1 11 13 1 0 9 1 9 2
17 3 15 13 0 9 2 4 10 0 9 0 1 9 3 12 9 2
10 15 4 1 10 9 3 13 1 9 2
13 7 0 4 9 3 12 9 3 13 1 10 9 2
12 9 1 9 13 3 1 0 9 3 7 9 2
29 10 0 9 1 11 7 1 0 9 13 13 16 10 0 9 1 9 7 9 4 3 0 2 3 1 9 1 9 2
26 0 9 13 3 1 10 9 16 10 9 9 1 0 9 4 2 0 2 1 10 0 9 1 9 9 2
22 10 3 0 1 10 2 1 10 0 0 2 9 4 1 3 0 9 3 13 1 9 2
12 10 0 9 13 0 3 7 0 9 7 0 2
16 1 10 9 14 13 9 7 13 1 9 4 15 13 10 9 2
26 2 12 9 1 12 7 12 9 1 11 9 1 12 7 12 9 4 13 15 0 1 9 1 10 9 2
20 10 0 9 13 2 7 10 9 4 13 1 1 9 12 0 9 0 9 2 2
21 2 1 9 1 9 1 9 12 1 10 9 1 10 0 9 1 9 1 11 2 2
18 0 9 1 9 7 10 9 13 1 9 2 15 13 1 9 12 12 2
20 15 13 12 9 9 2 15 1 10 9 4 13 9 7 9 1 12 9 9 2
23 9 9 1 9 7 9 4 3 0 1 9 2 9 13 1 0 9 2 9 1 9 3 2
9 9 9 13 3 10 9 1 9 2
32 9 9 13 1 0 9 1 9 16 9 1 10 9 2 15 9 13 1 2 4 13 9 1 9 1 14 13 9 2 9 2 2
17 10 9 4 13 1 10 3 0 9 1 9 1 9 1 9 9 2
15 1 9 7 3 3 1 9 4 10 0 9 3 3 13 2
22 9 4 13 3 16 10 0 9 13 15 1 14 13 0 9 7 13 1 10 0 9 2
10 0 9 1 9 13 15 3 0 0 2
14 9 4 1 0 9 2 3 9 7 9 2 13 9 2
22 10 0 7 0 9 4 13 1 16 9 13 3 3 0 3 1 9 0 9 7 9 2
12 10 9 1 9 13 1 9 12 9 12 9 2
19 3 15 13 0 9 13 9 1 9 0 9 1 9 2 3 9 1 9 2
10 1 3 0 9 13 3 9 1 9 2
12 9 1 9 9 4 1 10 0 9 4 0 2
17 9 4 13 1 0 9 2 9 4 1 9 9 10 3 0 9 2
12 10 0 13 3 7 13 1 0 9 1 9 2
9 7 9 1 9 13 3 0 9 2
33 3 9 4 13 10 0 9 13 1 10 9 9 2 9 2 9 2 9 9 7 10 9 7 10 9 15 9 7 9 13 15 1 2
1 9
7 10 9 4 13 1 9 2
11 3 3 4 0 9 13 1 12 1 12 2
10 13 9 12 2 9 12 2 9 2 2
9 10 9 1 9 13 1 0 9 2
27 13 3 9 9 12 2 9 2 9 7 0 9 2 2 11 3 2 9 12 2 11 2 9 10 0 9 2
18 3 4 9 2 7 3 9 2 1 11 13 3 3 1 12 7 9 2
18 13 11 12 2 9 12 2 11 2 9 12 2 11 3 2 9 9 2
22 10 9 4 12 10 0 1 9 9 2 9 2 9 2 9 2 9 2 9 2 9 2
5 13 9 1 9 2
7 13 11 12 2 9 12 2
10 13 9 1 0 9 1 12 7 12 2
9 13 9 12 7 12 2 9 2 2
8 13 3 11 3 2 9 12 2
10 10 9 14 13 9 13 7 4 13 2
19 13 11 12 2 9 12 2 11 2 9 12 2 11 2 9 9 7 9 2
13 1 10 9 4 10 0 9 0 1 9 7 9 2
13 13 11 2 9 0 9 1 9 2 11 11 2 2
8 15 13 9 1 9 0 9 2
15 10 9 4 10 9 13 2 7 13 15 3 2 1 9 2
26 13 11 3 2 9 0 9 2 11 2 9 12 2 11 2 9 1 11 7 11 2 11 2 9 12 2
23 3 4 15 1 9 4 13 9 7 9 2 3 13 9 1 9 1 14 13 9 1 9 2
30 13 11 3 2 9 9 1 9 7 9 9 7 9 2 11 2 9 9 3 2 11 2 9 9 7 9 2 11 2 2
5 0 9 1 0 9
26 7 15 13 16 9 1 15 1 10 9 13 0 2 4 0 1 0 9 1 10 9 2 1 10 9 2
21 13 15 13 1 9 2 9 1 10 0 9 2 3 9 9 1 9 1 0 9 2
27 1 0 9 4 10 9 0 1 0 9 16 3 1 0 9 0 1 9 7 9 2 13 9 9 1 9 2
2 9 2
48 9 13 3 0 10 9 2 7 9 4 1 3 0 9 7 13 1 3 0 9 13 9 1 9 9 7 13 9 1 15 9 13 3 2 3 16 15 13 0 0 9 1 0 9 7 0 9 2
36 10 9 15 13 1 15 3 4 1 10 9 3 0 1 9 1 0 9 7 1 10 9 1 10 9 2 1 9 1 10 9 7 1 9 9 2
27 9 7 9 3 4 13 7 3 13 9 1 0 0 9 3 15 3 3 13 3 9 1 0 9 7 9 2
14 9 1 9 2 1 0 9 7 1 9 4 3 0 2
57 3 2 1 9 1 9 7 1 9 1 9 7 9 1 9 2 13 10 0 9 2 10 0 9 7 9 7 10 3 0 1 10 0 0 9 2 15 13 7 0 9 1 9 3 2 1 0 7 0 0 2 0 9 1 0 9 2
22 3 0 7 0 4 3 3 9 1 9 1 9 9 3 1 15 7 1 9 1 15 2
31 9 3 3 0 9 13 2 15 1 9 13 3 1 10 1 9 7 9 0 9 7 10 1 10 0 9 0 9 1 9 2
10 1 10 10 0 9 9 13 9 3 2
49 3 1 9 15 3 3 1 9 7 1 0 9 1 9 1 0 7 10 9 7 3 1 9 1 9 1 0 9 7 10 9 3 2 9 0 9 7 9 7 10 0 9 2 13 2 14 13 3 2
11 1 9 13 15 9 15 13 9 7 9 2
43 7 9 2 15 4 10 9 10 9 13 1 9 2 9 2 9 2 13 9 1 9 2 9 2 9 2 9 2 13 1 7 1 9 2 13 1 9 2 13 1 9 3 2
50 9 2 15 4 10 9 15 13 3 0 1 9 1 15 15 13 9 7 15 13 9 2 13 9 1 15 9 2 13 2 7 15 3 13 9 2 1 9 2 9 2 2 9 2 9 2 9 7 9 2
33 1 0 9 2 13 9 1 2 1 9 7 13 9 7 13 15 3 1 9 1 9 2 16 9 13 7 13 1 9 3 9 13 2
2 0 9
11 9 1 9 1 10 9 4 3 3 0 2
12 4 15 3 1 0 9 13 16 15 4 0 2
19 9 15 3 1 9 2 1 9 2 1 0 9 4 0 1 9 7 9 2
25 9 15 13 9 1 9 1 0 9 15 15 3 13 1 1 9 7 9 1 9 1 9 7 9 2
44 9 15 3 3 13 1 0 9 1 0 9 7 0 9 1 15 7 3 13 1 10 9 2 0 0 1 9 7 9 0 9 7 9 1 10 9 3 15 4 13 10 0 9 2
40 9 2 0 1 9 15 13 15 7 10 9 2 7 0 1 7 0 1 10 3 0 9 1 10 0 0 9 7 1 9 7 9 0 0 7 1 9 0 9 2
33 3 13 15 15 1 10 0 9 14 1 9 7 9 13 1 9 1 10 9 7 10 9 7 3 1 9 1 10 1 9 0 9 2
53 7 3 1 10 9 13 15 15 7 0 14 13 7 13 10 0 9 2 10 9 2 7 9 2 7 0 9 1 0 7 0 9 2 3 7 9 3 1 9 2 9 2 9 2 7 7 9 3 1 9 2 9 2
19 3 13 15 1 9 15 13 3 1 15 1 15 15 13 9 9 1 9 2
22 9 15 1 3 0 9 13 10 0 2 0 9 1 9 1 0 9 2 1 0 9 2
6 4 3 0 4 9 2
2 9 9
24 10 0 9 4 1 0 9 10 0 9 1 16 9 4 13 13 15 7 3 1 10 0 9 2
31 15 4 3 4 13 16 10 0 9 1 10 9 4 3 1 16 10 9 4 3 0 2 3 0 1 3 15 3 13 15 2
35 3 11 13 10 0 9 1 11 1 9 0 9 2 4 15 9 1 10 9 16 10 0 9 4 13 1 9 1 10 9 7 0 0 9 2
17 3 13 7 11 7 9 1 9 0 10 9 1 3 9 4 13 2
21 3 10 0 9 3 4 13 10 9 1 9 2 13 15 10 9 1 10 0 9 2
19 1 9 1 9 9 13 9 13 15 16 15 13 9 0 9 15 13 9 2
32 1 15 13 15 9 16 10 9 3 3 4 10 3 0 9 7 16 15 13 9 1 10 0 9 7 9 1 0 7 0 9 2
14 3 4 3 9 13 3 7 1 9 1 0 0 9 2
16 1 9 13 15 3 0 14 13 9 9 1 10 0 0 9 2
30 10 9 13 3 1 0 9 0 0 9 1 15 9 13 7 10 0 9 7 3 0 9 13 7 0 9 1 9 9 2
3 11 7 9
29 16 10 9 13 0 9 1 9 7 9 9 2 13 15 3 0 9 14 1 9 13 10 0 9 7 13 10 0 2
23 9 13 3 16 10 0 9 1 9 7 3 0 2 4 13 1 10 9 1 9 7 9 2
14 15 4 3 1 10 0 9 13 7 10 3 0 9 2
23 15 4 3 10 9 1 16 11 1 9 1 11 9 3 4 13 16 9 1 9 4 0 2
31 15 13 3 3 9 9 1 10 9 16 10 9 13 7 10 9 3 3 1 10 9 7 3 1 15 15 13 15 3 3 2
22 10 9 15 9 13 1 11 9 2 11 12 9 2 4 3 13 14 13 10 0 9 2
3 10 0 9
19 3 13 10 0 9 3 15 13 2 16 9 4 10 0 9 1 0 9 2
12 1 0 9 13 15 9 7 9 1 11 9 2
14 9 4 2 3 3 13 2 10 0 7 0 0 9 2
13 15 4 1 0 9 3 3 3 0 1 10 9 2
18 7 15 13 1 10 0 9 10 9 2 15 4 13 10 9 9 13 2
22 15 4 10 0 9 1 10 9 15 13 1 10 9 2 3 9 13 7 9 0 9 2
29 7 15 13 3 16 15 13 1 9 7 10 9 0 9 2 1 15 15 3 13 0 7 0 9 1 10 0 9 2
19 3 13 15 3 3 14 13 0 9 7 9 1 9 1 0 9 1 9 2
20 0 9 1 10 0 9 4 3 13 7 10 0 0 9 1 0 9 1 9 2
29 9 9 4 14 13 10 0 9 3 16 10 9 15 13 1 0 9 1 10 0 9 13 1 9 7 13 1 9 2
26 15 13 16 3 13 10 0 9 1 9 0 2 3 3 16 10 0 9 4 3 3 0 7 10 0 2
21 3 4 3 13 10 0 9 7 13 15 10 9 1 3 10 9 7 0 0 9 2
8 15 4 10 0 9 7 9 2
21 10 0 9 4 0 7 0 1 9 7 9 1 10 9 15 3 13 10 0 9 2
26 3 15 4 10 0 9 2 10 0 9 2 9 7 9 3 13 2 3 15 13 10 9 1 0 9 2
13 10 0 9 4 3 0 1 9 1 15 15 13 2
18 9 2 9 2 10 0 9 2 10 0 9 4 9 1 0 0 9 2
12 7 10 9 4 3 13 10 0 9 1 9 2
5 0 9 7 0 9
22 3 10 0 9 13 0 0 9 2 4 10 0 9 13 0 9 1 0 9 1 9 2
34 7 3 13 10 0 9 2 16 10 9 9 2 15 3 13 13 10 0 9 2 13 0 9 1 0 9 7 9 15 13 1 0 9 2
12 10 0 0 9 13 3 3 1 9 7 9 2
17 15 13 9 2 16 10 0 9 4 13 0 9 1 10 0 9 2
23 3 13 15 3 10 9 1 0 9 15 13 0 9 1 10 0 9 7 1 10 0 9 2
11 0 9 13 9 0 9 1 9 0 9 2
12 9 1 11 13 3 9 14 13 10 0 9 2
28 4 15 1 0 9 0 14 13 10 9 15 13 1 0 9 1 10 0 9 3 3 9 3 13 10 0 9 2
13 15 4 10 0 9 7 0 9 13 15 4 0 2
25 16 9 9 4 0 1 10 0 0 9 2 4 15 3 3 9 1 0 9 1 0 3 0 9 2
29 15 13 10 9 1 9 9 1 10 9 15 3 13 13 2 3 16 15 4 0 1 9 1 10 0 7 0 9 2
14 10 0 9 13 9 7 0 9 1 15 1 10 9 2
20 10 0 9 4 1 0 9 3 13 1 9 1 0 9 15 3 13 10 9 2
20 7 1 10 0 13 15 9 2 3 9 1 9 15 4 4 0 9 1 9 2
5 9 9 2 14 13
19 15 13 16 15 13 9 1 0 0 9 2 15 13 0 9 7 0 9 2
24 15 4 3 13 9 1 10 9 9 15 10 0 9 4 13 2 16 15 4 13 10 0 9 2
22 1 0 9 13 9 7 10 0 9 16 15 3 0 13 10 0 9 1 10 0 9 2
32 3 0 13 10 0 9 1 9 10 0 9 1 10 0 9 1 10 9 3 9 13 10 0 9 1 10 0 9 1 12 9 2
14 15 13 3 10 0 9 15 1 10 9 4 13 9 2
30 10 0 9 1 10 9 15 13 1 0 9 1 9 7 10 0 0 9 1 10 9 2 4 3 14 13 0 1 9 2
18 15 4 3 14 13 0 15 13 1 10 0 0 9 9 1 0 9 2
17 3 3 9 13 9 7 9 1 0 9 2 13 10 9 7 9 2
26 15 4 3 0 7 3 15 13 9 1 0 9 1 16 15 2 13 2 10 9 1 14 13 10 9 2
32 15 13 3 13 16 15 3 4 9 1 14 2 13 1 2 2 16 15 3 3 4 13 10 9 1 16 15 2 13 2 15 2
22 15 13 15 3 3 1 9 7 4 3 13 1 10 0 9 3 15 3 4 13 15 2
36 15 13 3 3 0 3 15 13 1 16 10 9 0 13 9 2 7 16 15 4 0 2 3 13 1 10 9 2 3 4 0 7 10 0 0 2
15 7 15 13 3 3 3 9 1 9 15 15 4 13 3 2
16 15 13 3 9 3 2 9 2 9 2 15 15 15 13 1 2
11 3 4 10 0 13 9 7 10 0 9 2
8 7 16 15 4 9 1 9 2
23 15 4 3 0 9 2 15 13 15 2 10 9 13 0 1 15 7 9 4 3 10 0 2
18 15 4 3 9 1 15 7 16 15 13 15 3 0 1 10 0 9 2
13 15 4 0 9 7 4 13 10 9 3 15 13 2
13 3 15 3 13 3 1 9 13 15 3 3 0 2
20 15 4 14 13 0 14 13 9 7 15 4 14 13 0 14 13 3 10 9 2
13 10 0 13 3 10 2 0 2 9 7 10 0 2
14 7 9 1 9 1 9 7 9 13 15 13 3 1 2
34 10 9 13 3 3 3 0 1 15 16 10 9 13 13 10 3 0 7 15 4 3 3 13 3 0 1 10 9 16 15 13 0 9 2
8 3 13 15 15 1 0 9 2
43 7 9 1 9 13 15 13 0 9 3 16 15 4 0 1 16 10 0 9 1 0 3 7 3 3 0 7 3 2 0 2 9 4 4 1 10 3 0 9 2 3 0 2
34 7 1 10 0 13 15 3 10 0 9 15 4 10 0 7 10 0 2 9 1 10 0 9 15 13 9 9 1 9 7 9 1 9 2
25 9 13 3 14 13 3 2 16 15 1 9 13 3 3 7 14 13 14 13 3 1 10 0 9 2
37 15 13 15 16 15 13 3 7 13 1 2 9 2 2 2 9 2 7 2 9 2 2 10 15 15 3 3 4 10 9 1 10 0 9 7 9 2
20 9 1 2 9 2 4 3 3 0 7 15 13 10 9 15 4 13 1 9 2
15 9 1 9 1 9 4 1 10 3 9 10 3 0 9 2
18 3 3 15 13 1 9 4 15 13 13 10 9 15 0 9 4 13 2
15 10 9 15 4 13 15 4 4 0 1 10 0 9 9 2
12 3 4 15 4 13 15 0 0 0 0 9 2
71 15 4 4 9 1 9 7 14 4 13 7 2 9 2 1 9 2 14 4 13 1 9 1 9 15 3 13 15 3 7 13 13 15 1 14 13 10 0 9 1 10 9 2 10 9 1 3 10 9 13 9 2 10 9 3 15 3 13 1 10 0 9 7 9 7 3 15 4 4 9 2
5 0 13 3 3 2
25 13 15 9 13 15 3 9 14 3 13 3 10 0 9 9 7 13 10 0 9 1 10 0 9 2
19 15 13 3 10 9 1 9 3 9 3 13 15 14 13 3 1 10 9 2
27 15 13 3 2 13 3 10 0 9 7 4 13 7 13 1 11 16 10 0 9 4 13 3 1 10 9 2
5 15 13 3 0 2
38 10 0 9 15 15 3 13 7 15 15 13 15 16 0 9 1 10 9 13 3 1 4 9 1 10 0 9 14 2 13 2 3 3 1 9 7 9 2
37 10 9 3 13 15 3 16 11 4 3 0 1 16 15 13 3 7 3 10 9 13 7 16 15 13 9 1 3 0 9 1 15 7 1 10 9 2
21 15 13 9 1 10 9 1 9 7 9 0 1 16 15 4 1 10 9 7 3 2
24 15 4 10 9 9 7 15 13 16 15 4 0 16 9 1 0 9 4 0 1 10 9 9 2
20 15 4 3 13 1 14 13 9 1 0 9 2 15 15 3 4 4 0 1 2
15 15 13 1 9 14 3 13 10 0 9 1 10 0 9 2
24 9 13 3 16 15 13 9 1 10 9 7 13 9 13 1 9 1 3 15 3 0 7 9 2
48 3 4 15 3 4 0 1 14 13 16 15 13 0 9 7 16 15 3 3 3 4 13 9 7 16 9 1 9 4 13 3 0 3 16 0 9 13 3 1 9 2 7 9 9 2 3 2 2
68 10 9 15 15 13 0 14 13 4 15 15 10 1 9 1 0 0 9 11 11 13 9 1 1 10 9 1 11 2 12 2 3 15 13 16 15 3 4 13 2 9 9 1 9 7 9 7 1 10 0 15 13 14 13 2 15 7 15 1 10 9 2 2 11 0 9 2 2
31 15 13 15 7 10 9 1 10 0 9 1 9 15 15 13 3 4 13 2 10 9 2 3 9 13 10 9 1 9 2 2
30 9 1 10 0 9 4 13 16 16 9 4 0 1 14 13 9 1 9 7 9 2 9 13 9 1 10 0 9 9 2
8 15 4 15 3 13 1 1 2
51 16 9 3 4 1 0 9 0 7 9 7 3 4 13 9 3 4 15 13 3 0 2 9 2 1 9 7 9 7 9 13 9 14 13 3 1 15 3 16 15 4 13 4 3 0 7 3 0 7 9 2
20 9 1 9 7 9 4 3 15 3 0 7 15 15 13 1 9 2 9 2 2
34 15 13 15 3 3 1 10 0 9 1 0 9 15 15 13 9 1 7 1 10 0 9 3 9 13 3 15 14 13 7 13 7 9 2
40 16 3 10 9 4 0 1 10 9 3 4 3 10 9 16 9 3 4 13 10 0 2 9 2 1 10 0 9 7 9 4 9 1 9 3 1 9 1 9 2
17 15 4 3 0 16 15 13 0 9 14 13 3 10 9 1 9 2
5 9 1 9 7 9
43 10 9 1 9 15 13 0 0 9 1 0 9 9 4 3 13 9 1 7 13 3 0 9 2 7 15 4 13 1 10 0 9 1 0 9 1 9 1 9 1 9 9 2
15 10 0 9 4 0 2 3 0 1 10 9 1 0 9 2
15 10 3 0 9 14 13 0 9 4 13 0 1 3 0 2
36 16 10 0 9 15 13 10 0 9 1 9 16 15 13 3 1 9 13 1 10 3 0 7 3 0 1 9 4 10 9 10 9 3 1 9 2
22 0 9 9 13 9 1 10 9 1 0 9 7 0 9 15 13 1 0 9 1 9 2
16 10 0 9 1 2 0 9 7 9 2 13 3 10 0 9 2
26 10 0 9 4 13 3 0 0 9 4 1 10 9 0 9 2 10 9 15 15 3 13 9 14 13 2
18 1 0 9 1 9 9 13 10 9 1 9 7 9 15 13 1 9 2
26 1 10 0 9 9 4 13 10 0 9 15 3 4 14 13 0 9 1 10 0 9 1 9 1 9 2
2 9 9
30 9 4 3 13 10 0 9 7 10 9 1 9 0 9 7 9 16 9 13 0 9 1 9 1 0 0 7 0 9 2
34 0 1 9 7 1 10 9 9 13 15 3 9 1 0 9 2 9 2 9 2 0 9 7 0 9 15 13 9 9 7 9 1 15 2
26 1 10 0 9 13 15 0 9 1 10 0 2 3 0 7 1 0 9 3 0 9 9 1 10 9 2
28 1 10 9 1 9 9 13 15 14 13 1 12 9 2 1 0 9 9 0 9 7 1 0 9 9 9 3 2
44 1 10 0 9 4 15 13 1 15 9 15 4 10 0 9 16 9 13 1 9 2 1 14 3 13 9 2 14 13 0 10 9 0 9 1 9 2 0 9 2 9 7 9 2
45 0 9 4 13 16 9 4 0 14 13 10 9 0 9 7 0 9 2 7 16 3 10 2 9 2 1 9 13 9 7 10 9 1 0 9 15 4 4 13 1 9 14 13 9 2
29 13 9 9 3 3 1 9 7 9 2 0 9 2 10 9 1 9 1 9 1 10 0 9 1 10 0 0 9 2
28 1 9 13 15 1 9 1 0 9 2 3 15 13 13 10 9 15 3 13 15 16 9 4 13 1 10 9 2
29 3 4 13 0 12 9 1 2 0 9 2 2 9 2 9 2 9 7 9 2 9 7 9 2 9 7 0 9 2
24 1 10 9 9 1 10 0 9 13 7 13 10 9 15 13 3 3 13 15 13 10 0 9 2
31 1 10 0 9 4 15 13 15 16 3 10 0 9 1 9 13 10 9 1 10 0 0 9 1 9 1 10 0 0 9 2
26 15 13 9 0 0 7 0 9 1 10 0 9 1 0 0 0 9 1 15 9 3 13 13 0 9 2
21 9 4 3 13 9 1 16 9 1 9 7 9 1 9 7 0 9 4 3 0 2
19 15 4 13 16 1 9 7 9 9 4 9 9 1 0 0 9 13 0 2
30 3 13 15 16 9 9 1 10 0 9 3 1 0 9 13 3 1 14 13 0 9 7 16 0 9 4 10 0 9 2
17 1 10 9 13 10 0 0 9 7 1 0 7 9 7 1 9 2
32 10 9 15 3 13 16 9 13 9 9 2 0 1 10 0 7 0 9 2 0 1 14 13 10 9 1 9 1 10 0 9 2
31 15 13 14 13 16 10 9 1 9 15 4 13 4 10 0 7 3 15 15 9 13 10 9 1 4 10 0 0 0 9 2
60 9 1 10 3 0 9 1 10 0 9 1 10 0 7 9 1 9 2 3 9 1 9 1 9 14 13 9 9 1 0 9 7 14 1 0 9 13 7 13 3 9 1 0 2 0 7 0 9 13 9 1 3 0 0 9 7 9 1 9 2
65 16 9 3 1 9 13 1 9 9 2 16 15 1 9 1 16 9 4 0 1 10 0 9 3 13 15 3 1 10 9 7 10 9 7 16 9 1 9 9 7 9 9 3 13 2 3 13 3 9 1 9 1 10 9 1 9 7 10 9 1 10 0 9 13 2
21 7 10 0 9 13 3 10 0 9 15 4 13 9 1 10 0 9 14 13 9 2
33 1 14 13 9 13 9 9 1 9 7 0 0 9 7 13 14 13 1 10 9 1 10 9 3 9 9 1 9 4 7 3 0 2
27 9 13 16 10 0 9 4 14 13 15 1 9 1 10 0 9 15 4 3 0 1 10 0 9 7 9 2
3 9 1 9
21 13 9 3 15 1 2 3 7 3 2 3 10 9 7 10 9 4 13 1 9 2
12 15 4 2 1 9 2 9 1 10 0 9 2
20 16 15 13 2 3 11 13 9 1 10 9 2 1 9 7 9 2 13 15 2
11 2 7 11 13 15 2 11 13 1 15 2
13 2 4 0 7 13 15 7 13 9 2 2 2 12
4 12 9 12 2
10 1 0 9 9 13 15 1 12 9 2
11 9 4 1 11 0 1 2 9 9 2 2
17 16 15 3 13 2 16 9 4 11 2 13 10 9 4 9 9 2
2 3 2
2 0 2
2 0 2
32 7 3 11 3 13 10 0 9 14 4 2 0 2 2 4 9 9 3 0 2 10 0 9 4 13 1 2 16 0 9 13 2
22 9 7 9 4 3 13 1 11 0 9 2 14 13 9 13 3 16 0 9 3 13 2
19 10 0 9 1 9 9 15 3 3 4 13 2 13 3 7 3 10 9 2
36 1 0 9 13 3 2 16 3 9 1 7 9 1 14 2 4 0 2 3 13 1 12 9 2 4 15 3 3 9 1 10 9 1 0 9 2
19 3 4 15 13 1 9 1 9 1 9 0 12 12 0 2 0 2 9 2
10 0 4 11 11 1 0 9 13 15 2
72 11 13 2 16 10 0 9 2 1 15 13 2 13 7 13 3 10 0 2 0 9 2 16 15 4 13 15 1 10 0 9 7 3 2 3 0 4 2 13 9 7 9 1 0 9 2 3 1 9 2 7 1 16 15 4 13 3 2 4 0 2 13 9 2 13 7 13 15 1 11 9 2
40 7 15 13 1 11 10 9 1 2 16 15 13 9 2 15 4 9 1 9 7 13 11 9 2 10 0 9 7 10 9 2 3 16 9 7 9 13 2 2 12
6 12 9 2 9 12 2
11 9 2 9 7 9 4 3 9 0 9 2
42 1 0 3 0 12 12 0 2 0 2 9 1 9 13 3 12 0 9 13 2 3 3 12 9 2 12 9 9 12 0 9 12 0 1 9 12 9 1 10 0 9 12
7 12 11 0 2 9 12 2
31 1 10 9 13 15 2 1 10 0 9 1 9 9 2 9 1 9 2 15 3 13 15 10 0 9 1 0 9 1 9 2
21 1 10 9 4 15 3 3 3 0 2 16 15 1 9 9 13 15 2 7 15 2
10 2 15 13 15 1 14 13 9 2 2
10 7 3 4 10 9 1 9 3 0 2
30 1 10 2 9 7 9 1 9 7 0 9 3 2 1 10 0 9 1 9 2 9 12 2 13 9 11 3 10 9 2
29 10 0 9 15 13 1 2 4 15 2 16 15 13 10 0 9 1 9 7 9 2 6 2 1 10 9 7 9 2
19 0 10 9 2 10 9 1 9 1 15 4 3 1 15 0 0 7 0 2
28 0 7 0 13 9 2 3 15 1 9 2 9 7 9 13 1 0 9 1 9 1 15 1 11 1 9 0 2
12 15 13 1 10 9 3 9 11 13 10 0 2
23 2 7 1 14 13 9 4 10 9 13 10 0 9 2 7 10 9 10 0 9 2 2 12
5 12 0 9 12 2
7 13 9 1 2 1 14 2
19 3 4 0 2 16 1 10 9 10 1 9 9 4 15 2 9 1 9 2
9 1 10 9 4 11 11 3 13 2
3 15 13 2
60 2 7 3 9 13 10 9 2 0 11 4 13 15 2 4 15 3 0 14 1 9 13 0 2 7 9 7 9 13 9 7 9 2 7 10 0 9 7 9 13 2 1 16 15 4 13 7 13 15 2 10 9 2 3 10 9 13 7 13 2
60 1 16 15 3 4 4 0 14 1 10 9 2 3 2 2 13 9 2 4 3 11 13 10 0 9 2 1 15 15 7 15 4 13 10 0 9 7 13 13 15 3 2 16 3 3 11 9 4 0 2 1 16 3 9 4 13 0 2 2 12
6 12 11 2 9 12 2
42 13 15 3 2 10 0 9 15 9 4 13 1 15 2 15 13 1 11 9 2 13 9 2 14 1 9 0 9 13 13 3 15 1 11 9 1 10 0 9 1 9 2
41 10 11 9 4 3 0 9 1 15 15 1 10 9 3 13 1 9 9 2 15 13 1 7 2 13 2 15 15 4 0 2 0 2 3 0 2 1 10 9 0 2
25 10 9 0 9 4 3 3 10 0 9 2 15 13 15 0 2 10 0 9 15 13 1 10 0 2
14 11 11 13 3 9 1 10 9 2 16 15 13 10 2
7 15 13 1 12 9 10 2
4 1 9 9 2
25 9 1 10 9 4 3 10 0 13 13 1 10 9 2 3 0 3 1 10 0 9 1 11 9 2
27 3 4 15 1 9 4 10 9 0 1 0 9 1 9 1 10 0 9 7 14 2 13 15 0 2 3 2
26 9 2 9 2 10 0 4 2 3 1 9 2 3 1 10 9 2 16 15 4 13 7 13 0 9 2
27 16 10 9 1 10 2 9 2 2 1 10 2 9 2 4 0 1 9 2 13 10 0 9 9 1 9 2
24 15 13 1 9 1 10 9 2 3 11 9 4 13 9 2 3 9 1 9 7 9 4 13 2
20 15 13 3 2 16 15 13 0 14 13 9 1 11 7 11 11 1 10 9 2
7 2 9 4 3 13 9 2
16 7 3 3 13 15 3 10 9 1 9 1 14 13 10 9 2
20 15 4 0 3 14 13 3 15 15 3 4 15 0 1 10 0 9 2 2 12
8 12 11 9 9 2 9 12 2
36 2 15 15 3 4 15 0 2 2 6 0 9 2 2 4 2 1 9 9 1 9 2 7 13 3 1 10 9 9 7 13 1 15 10 9 2
22 7 1 9 13 15 15 3 3 1 12 9 2 15 7 4 13 2 7 13 1 15 2
11 15 13 15 1 11 0 9 7 9 0 2
29 9 1 9 4 3 1 9 3 13 14 2 13 15 0 2 7 4 9 1 16 10 0 4 2 13 15 0 2 2
34 9 1 9 1 9 7 0 9 13 2 1 14 13 2 12 9 1 9 12 9 1 9 12 9 1 3 0 9 2 3 11 4 13 2
3 10 0 9
5 15 4 10 9 2
36 3 15 1 10 0 9 9 13 1 9 2 13 15 10 9 1 9 7 9 2 15 13 3 7 3 2 7 15 1 9 4 0 14 4 0 2
27 3 13 15 3 3 9 1 2 9 2 15 13 10 9 1 9 9 7 9 7 0 9 15 13 1 9 2
6 10 15 4 0 9 2
12 3 13 3 9 10 0 9 1 10 0 9 2
24 6 2 3 7 3 4 3 15 2 0 1 10 0 7 0 9 2 3 10 3 0 1 9 2
32 9 9 7 9 4 13 1 0 9 1 0 9 2 7 15 4 3 3 15 13 3 1 0 9 4 10 0 9 1 0 9 2
31 3 15 1 0 9 4 13 10 0 9 2 9 1 15 13 3 0 1 15 15 3 13 2 2 15 3 11 4 13 2 2
23 1 9 1 9 1 0 9 13 15 3 13 1 16 11 13 9 4 2 10 0 9 2 2
21 15 13 16 15 4 10 0 9 2 15 3 1 7 1 15 13 10 0 1 15 2
24 15 13 3 16 15 3 13 9 15 1 10 9 13 9 2 15 13 1 9 10 0 9 0 2
44 3 4 15 3 3 3 15 4 13 13 10 3 0 9 1 15 9 4 1 15 1 0 9 1 14 13 1 9 15 3 2 3 1 10 9 3 2 4 13 4 2 0 2 2
15 3 13 15 3 2 0 2 7 2 0 2 4 3 0 2
21 3 4 9 1 9 0 9 1 9 4 10 0 9 2 3 9 13 9 1 9 2
22 7 9 9 4 3 13 1 15 2 15 13 14 13 10 0 9 15 4 3 3 0 2
44 3 16 15 13 15 10 9 0 9 2 3 9 13 0 9 1 9 2 7 10 9 13 3 10 9 1 9 1 10 9 9 3 2 3 4 15 3 13 9 9 1 0 9 2
22 15 13 3 10 9 9 1 15 15 3 13 1 9 9 1 10 0 9 1 0 9 2
36 15 4 3 3 0 1 9 10 0 9 15 4 13 1 10 0 9 2 7 1 10 10 9 13 15 9 14 13 10 0 9 1 10 0 9 2
4 15 13 9 2
8 15 13 15 3 15 13 9 2
14 15 4 10 9 15 13 3 3 15 13 10 0 9 2
29 3 13 3 1 0 9 10 9 3 9 2 15 13 9 3 3 3 16 15 4 10 9 15 3 13 1 0 9 2
24 10 0 9 1 10 3 9 4 13 1 10 0 0 9 2 15 4 13 3 9 3 4 13 2
8 10 3 9 9 4 3 13 2
12 7 15 13 10 9 14 13 15 1 10 9 2
30 15 15 3 4 13 13 16 15 13 12 9 15 3 13 10 0 9 2 9 0 9 7 9 1 9 1 10 3 9 2
21 10 0 0 9 13 15 3 1 10 9 2 16 3 0 9 13 9 7 10 9 2
15 3 3 13 15 3 10 0 9 15 13 9 2 3 9 2
37 15 4 3 0 16 15 3 13 10 9 2 3 15 4 13 15 0 9 1 0 9 2 7 3 10 9 3 1 7 1 15 4 13 10 0 9 2
15 1 0 9 4 3 10 0 9 3 3 0 7 10 0 2
26 7 15 4 0 14 13 3 15 4 4 13 1 10 12 0 9 9 1 10 0 9 2 9 7 9 2
29 3 4 15 3 0 16 10 9 13 0 9 1 10 9 1 9 7 9 2 7 15 4 3 0 13 13 10 9 2
13 3 4 3 3 3 9 13 1 0 7 0 9 2
20 1 15 15 3 13 4 15 3 0 3 0 9 3 4 13 15 1 0 9 2
27 15 4 0 14 13 3 15 2 1 14 13 3 9 1 10 9 2 4 4 13 10 0 9 1 0 9 2
34 3 0 2 7 1 9 1 9 1 10 9 2 4 9 1 0 9 1 12 9 2 15 13 16 15 4 13 3 2 13 2 13 15 2
18 10 9 2 13 15 2 2 13 0 9 15 15 13 9 14 3 13 2
25 3 7 3 4 15 1 10 0 9 0 16 0 9 1 0 9 1 9 13 3 2 3 7 3 2
12 15 13 3 10 9 1 9 9 1 0 9 2
27 3 3 4 10 9 13 1 0 0 9 2 9 2 9 1 9 2 3 0 0 9 3 1 10 0 9 2
17 1 9 1 9 1 10 9 2 9 2 9 1 0 7 0 9 2
27 1 15 15 13 3 2 7 3 4 15 3 3 13 3 3 2 13 3 15 2 9 2 1 10 9 9 2
2 9 9
43 10 0 7 0 9 1 10 9 1 0 9 14 13 15 4 2 16 15 13 1 10 0 1 16 9 4 13 15 9 1 0 9 2 3 15 3 3 3 4 0 1 15 2
23 15 4 10 9 15 15 13 10 9 14 13 2 7 15 13 15 1 9 1 10 0 9 2
16 1 9 13 15 9 1 9 3 15 3 4 0 1 10 9 2
13 15 4 3 3 3 13 15 10 0 9 1 9 2
11 7 15 13 3 3 3 16 9 4 13 2
30 7 15 13 15 3 1 10 9 9 2 15 15 4 3 0 3 7 3 2 7 15 3 3 1 0 9 4 13 0 2
9 10 0 9 13 3 1 10 0 2
32 3 13 15 3 0 9 2 15 3 13 0 1 14 13 10 0 3 9 1 0 9 2 7 15 16 15 13 15 3 3 13 2
9 15 4 0 16 10 9 13 3 2
26 3 13 15 15 3 3 0 2 16 0 9 3 3 13 15 1 14 1 3 13 1 10 0 0 9 2
10 3 0 4 15 3 1 11 0 9 2
17 15 3 13 0 9 3 1 9 0 9 2 15 15 4 13 3 2
24 7 15 15 3 4 0 14 13 13 2 16 10 0 9 3 3 4 13 1 10 9 0 9 2
31 3 15 13 10 0 9 7 15 15 13 1 15 13 3 1 9 2 9 2 9 1 9 2 9 9 2 9 1 9 3 2
16 15 4 3 13 1 14 13 9 1 15 15 15 13 7 0 2
23 0 9 13 1 10 0 9 2 7 15 15 13 6 1 15 13 3 10 9 1 10 9 2
9 15 13 10 9 15 3 4 13 2
24 3 4 15 10 0 9 1 10 0 9 2 16 15 4 13 9 3 16 15 3 4 3 0 2
46 0 9 1 15 13 3 3 16 15 4 13 10 0 9 3 16 15 13 3 0 2 7 16 15 4 10 0 9 16 10 15 15 3 13 10 0 9 3 4 13 10 9 1 0 9 2
10 15 13 3 3 0 9 3 1 0 2
4 10 0 0 9
32 9 13 10 9 14 13 3 7 3 7 1 9 7 1 9 2 7 1 10 9 4 15 0 3 15 1 10 9 13 10 9 2
32 1 9 13 3 14 13 1 9 10 9 2 14 3 13 10 9 15 13 3 16 15 4 9 7 9 2 3 15 3 13 15 2
15 1 9 13 9 1 10 9 2 0 2 0 7 3 0 2
24 9 4 13 9 1 3 10 3 0 9 2 16 15 3 13 10 0 9 1 9 9 7 9 2
34 3 4 15 3 0 16 0 13 0 1 10 9 0 9 2 16 15 1 0 7 0 9 2 3 3 13 2 3 0 13 9 7 9 2
19 1 9 13 14 1 9 13 9 1 3 0 7 9 2 9 3 0 9 2
14 15 4 3 4 0 2 16 9 13 9 7 3 9 2
40 7 9 4 16 3 10 0 9 3 13 3 1 10 9 1 0 9 2 1 3 9 16 15 3 13 1 16 15 4 4 0 9 1 15 15 13 7 13 0 2
19 3 9 3 4 13 4 15 0 14 3 13 13 2 16 9 4 3 0 2
13 15 4 10 9 1 10 0 9 14 13 15 3 2
3 10 0 9
15 10 0 9 13 3 1 0 9 3 7 3 0 7 0 2
29 15 4 4 10 9 1 10 0 0 9 1 10 9 2 10 9 15 15 1 7 1 15 3 13 10 9 14 13 2
9 3 13 0 9 7 9 1 15 2
52 1 0 9 4 10 9 15 1 10 3 0 9 10 9 4 13 2 7 10 0 9 4 3 0 1 10 9 2 16 15 13 16 9 13 3 0 9 14 13 3 7 13 15 1 15 16 15 3 13 13 15 2
30 15 4 10 9 15 13 16 9 7 9 15 13 1 10 9 4 13 15 15 13 1 0 9 2 0 9 7 3 9 2
24 15 4 10 9 1 10 9 2 3 15 15 4 4 10 9 1 15 2 1 15 9 13 0 2
53 12 0 9 13 14 13 1 9 1 9 2 7 4 1 0 9 9 3 13 1 9 7 10 0 9 2 7 4 15 3 13 1 16 9 1 10 9 4 13 0 2 1 10 9 0 9 2 15 3 3 4 13 2
11 3 4 9 13 2 7 3 3 13 9 2
51 9 1 9 7 1 9 1 10 0 9 13 1 15 10 0 9 2 16 15 13 10 9 14 13 16 10 9 15 13 9 1 10 0 9 1 15 3 4 13 10 0 9 2 1 9 9 2 9 2 9 2
20 9 1 9 13 16 9 7 9 13 10 9 7 9 14 13 9 1 10 9 2
45 1 9 13 15 10 9 1 3 9 16 15 13 9 1 0 7 0 9 1 9 2 1 9 16 15 3 0 4 13 9 1 9 9 7 16 15 3 4 13 0 9 1 10 9 2
17 1 9 4 15 10 3 0 9 16 15 13 9 1 10 10 9 2
23 9 13 3 10 3 0 9 1 7 0 9 1 10 0 9 7 9 13 10 0 0 9 2
32 16 15 13 16 9 4 13 9 1 9 1 10 9 7 9 2 4 15 3 14 13 0 1 9 14 13 9 7 9 7 9 2
41 15 4 1 10 9 14 13 10 0 9 1 9 2 10 9 3 13 1 9 2 1 16 15 3 1 9 4 13 0 9 7 9 1 9 7 9 14 13 15 1 2
42 15 4 0 1 10 9 15 3 13 1 10 9 2 16 9 1 3 9 9 13 9 4 4 14 13 9 9 2 16 15 4 13 9 1 14 13 10 9 3 15 13 2
18 15 13 3 3 10 9 15 13 2 9 2 7 3 3 13 10 9 2
25 1 0 9 4 15 0 16 16 9 13 0 9 3 4 9 13 1 9 3 7 16 9 4 13 2
38 16 15 4 13 1 10 0 9 13 15 10 9 9 1 9 1 14 13 9 1 10 9 2 7 3 3 7 15 1 9 1 14 13 15 1 10 9 2
22 1 10 0 9 1 0 9 13 15 3 3 1 3 0 9 1 14 13 10 0 9 2
12 15 13 3 1 0 9 7 13 1 0 9 2
19 15 15 13 2 3 2 9 13 9 7 9 7 10 0 9 1 10 9 2
28 15 15 13 10 0 9 13 1 9 10 9 9 7 3 0 2 0 7 0 7 9 2 15 4 13 7 0 2
39 3 1 9 2 9 7 9 4 9 1 14 13 9 1 10 9 1 0 7 0 9 4 9 1 0 9 7 9 2 1 16 15 3 13 3 1 0 9 2
36 9 12 13 10 0 9 11 11 1 11 9 10 9 1 3 0 9 1 3 0 7 0 9 2 15 1 10 9 3 13 1 10 9 2 13 2
4 9 4 0 2
30 15 13 15 16 10 9 4 14 13 9 1 0 9 2 15 13 0 1 9 1 0 9 2 1 14 3 13 1 15 2
10 3 3 4 11 3 3 13 10 9 2
27 15 13 16 15 3 13 9 1 7 1 15 15 13 9 2 7 16 15 13 1 16 9 3 13 10 9 2
49 3 11 13 2 9 2 2 3 13 15 1 15 3 3 15 15 13 1 9 3 0 9 7 3 15 15 13 9 9 1 9 7 0 9 2 9 15 15 3 4 14 13 9 1 10 9 7 9 2
21 16 9 1 10 0 9 13 10 0 2 3 0 9 1 9 13 13 1 10 9 2
56 7 15 13 15 15 13 2 7 3 10 0 0 9 15 13 2 16 12 15 4 13 9 2 15 13 1 9 2 12 15 4 13 3 12 9 2 15 13 9 2 12 16 15 7 15 15 13 9 4 13 3 1 9 12 9 2
8 15 13 3 3 9 13 3 2
35 16 0 9 3 4 4 13 3 7 13 9 1 0 9 2 16 15 3 13 9 14 4 0 7 0 1 9 2 13 15 10 0 9 1 2
44 15 4 3 1 9 13 3 2 7 13 3 3 1 0 9 2 16 9 2 9 7 9 2 0 9 7 9 13 10 9 1 10 9 15 3 1 10 9 4 14 3 13 9 2
42 14 13 15 1 9 9 14 13 10 0 9 1 10 0 9 7 3 13 9 16 9 1 0 4 13 3 1 9 0 9 2 4 1 9 1 15 15 3 13 3 0 2
26 9 2 15 13 1 9 1 9 1 9 9 2 13 16 15 3 13 9 1 7 1 15 15 13 9 2
32 15 4 13 9 7 1 9 9 1 10 9 2 7 1 10 9 14 13 1 9 1 10 9 3 15 3 4 4 0 1 15 2
36 15 4 3 13 9 1 9 9 7 9 2 9 9 1 9 9 7 3 3 1 10 9 14 13 9 9 1 10 9 15 1 10 9 4 3 2
19 3 4 15 1 9 1 0 9 3 13 1 10 9 10 0 9 4 13 2
27 10 9 15 13 1 14 3 13 9 1 9 13 3 1 0 9 2 3 13 15 3 3 7 13 3 3 2
24 1 10 9 13 15 15 0 14 13 1 9 2 14 13 1 10 9 2 14 13 1 9 3 2
24 3 1 9 13 15 3 10 9 13 1 12 7 3 1 1 12 9 9 16 15 13 10 9 2
13 1 11 13 15 16 9 13 15 3 3 1 9 2
28 3 1 9 13 9 10 9 1 9 2 10 9 15 3 4 13 3 3 1 10 9 7 1 10 0 1 9 2
42 13 15 3 1 9 9 3 4 15 3 13 10 9 3 2 10 9 15 3 13 2 16 9 13 9 1 14 13 9 1 9 15 4 0 7 0 7 10 15 3 13 2
35 15 4 0 16 15 4 14 13 15 13 0 14 13 3 9 7 9 7 13 10 9 13 9 1 0 9 2 15 13 3 3 1 0 9 2
15 10 9 9 4 4 13 3 1 9 1 9 7 0 9 2
28 9 1 9 2 15 4 13 9 1 0 9 1 9 7 15 3 4 4 9 1 9 7 0 9 2 4 13 2
26 9 4 3 13 0 9 1 16 9 7 0 1 9 0 4 13 0 9 1 9 1 7 9 7 9 2
14 0 0 9 1 15 15 4 13 9 0 4 3 13 2
13 0 1 9 9 4 15 0 1 0 9 1 9 2
19 3 3 9 3 4 0 4 15 0 14 13 0 9 16 15 4 13 9 2
42 9 1 9 1 9 9 4 3 13 16 15 13 0 9 7 15 1 0 9 13 9 14 13 9 14 13 9 3 16 15 3 13 9 14 13 15 1 9 1 9 9 2
17 0 9 4 3 13 9 1 9 16 15 3 13 16 9 4 0 2
39 3 10 9 15 13 14 13 3 1 9 0 9 13 10 0 9 1 14 3 7 3 13 9 1 9 7 4 3 4 13 1 15 9 1 9 2 9 3 2
26 15 4 3 0 0 16 10 9 15 13 15 1 9 1 9 4 13 9 1 9 3 10 9 1 9 2
18 7 3 3 15 13 9 1 9 4 10 0 9 9 13 1 0 9 2
24 7 1 9 7 1 10 9 4 15 0 16 9 13 9 14 13 10 9 15 15 13 3 1 2
