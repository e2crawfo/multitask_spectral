2443 17
10 13 2 13 2 13 2 3 9 1 9
13 3 7 13 7 0 13 13 2 15 15 13 3 13
6 13 1 9 7 9 13
6 3 13 15 9 9 13
21 3 9 13 7 3 3 13 7 9 1 9 0 13 2 16 15 3 9 13 13 13
6 15 13 2 13 16 9
3 13 0 0
3 13 2 13
4 13 2 0 13
3 7 13 9
3 9 9 13
13 15 2 16 15 3 13 2 1 9 0 9 9 13
15 13 9 13 9 2 7 9 13 9 9 13 13 9 1 9
7 9 15 13 2 15 0 13
8 3 1 15 9 15 13 2 13
12 7 15 16 13 9 2 6 2 7 9 3 13
13 13 3 2 16 0 13 2 1 9 0 7 9 13
7 13 9 3 7 9 9 13
23 15 9 1 9 13 2 7 16 9 0 9 13 2 16 3 13 2 15 0 9 3 13 9
8 3 9 13 13 13 15 9 13
6 9 7 9 0 9 13
4 15 9 13 9
7 9 15 13 7 9 9 13
12 3 3 9 13 2 3 1 15 13 9 7 0
9 1 15 9 9 13 7 3 9 13
24 15 16 13 9 2 9 9 13 2 7 1 9 13 9 1 9 0 0 13 13 2 7 3 0
26 13 13 9 7 13 9 2 3 13 2 13 2 7 3 13 3 0 13 9 9 13 7 13 9 13 13
12 13 15 13 7 13 2 16 1 9 9 15 13
15 8 3 3 0 9 13 13 9 2 13 15 0 1 9 13
26 3 7 13 9 3 9 0 2 1 9 3 0 13 2 13 2 15 1 0 9 9 0 7 9 9 13
29 3 3 9 1 9 15 13 13 2 15 0 9 1 9 13 13 2 7 9 3 0 0 9 9 7 9 13 9 0
14 3 1 9 9 13 2 7 3 0 9 9 9 3 13
11 13 7 0 9 2 0 9 2 9 9 13
14 15 3 0 9 15 9 2 16 3 9 13 2 13 13
22 16 3 0 0 9 7 0 9 15 13 2 9 1 9 13 7 13 13 3 13 1 9
7 13 3 3 13 8 7 13
13 3 9 0 13 2 16 13 15 9 2 16 15 13
1 13
2 13 3
7 15 7 15 13 2 15 13
5 0 13 13 3 13
9 15 16 9 13 2 0 9 13 13
8 16 3 13 2 13 1 9 0
4 3 9 9 13
17 7 15 3 6 3 15 7 1 9 0 13 2 7 3 16 0 13
9 16 15 1 15 13 2 3 15 13
5 13 9 2 0 13
13 15 13 2 1 15 9 13 2 7 7 3 13 13
7 15 9 1 9 0 9 13
7 13 7 2 1 9 9 13
8 9 9 9 13 1 9 13 13
13 13 15 9 13 9 0 2 3 15 1 0 9 13
9 13 15 1 9 2 9 13 3 9
3 13 1 9
15 3 3 13 1 9 2 15 13 15 7 0 9 1 9 13
11 7 15 13 9 0 2 7 3 9 13 13
7 16 13 2 0 9 0 13
13 15 3 13 3 13 2 3 13 2 16 9 15 13
5 15 7 0 13 13
5 15 13 9 16 15
16 9 3 13 7 1 0 9 9 13 2 16 1 9 9 0 13
21 3 9 13 2 3 9 13 2 9 15 1 0 13 2 9 9 2 3 3 13 13
22 9 0 13 13 2 16 3 3 13 2 7 2 16 3 2 13 2 13 2 3 15 13
14 9 7 9 13 7 0 9 13 2 3 9 9 15 13
8 7 7 3 13 2 7 16 13
7 9 7 0 9 9 15 13
39 15 16 13 2 13 9 3 3 13 2 7 9 0 9 0 9 13 3 9 13 2 7 16 13 1 15 9 2 1 15 0 9 13 13 2 9 13 16 9
18 3 3 9 13 2 13 9 0 1 9 3 9 2 7 9 15 9 13
18 13 15 9 13 2 7 7 3 1 15 9 13 13 2 3 16 15 13
6 13 9 15 1 15 13
8 15 16 13 2 9 0 13 13
24 13 9 0 13 13 0 9 9 16 15 9 13 2 16 15 9 13 2 16 13 9 15 9 13
6 3 0 13 7 3 0
4 13 9 9 13
4 13 9 13 13
24 15 3 13 9 1 9 13 2 13 9 9 3 2 7 9 3 15 9 0 13 2 15 13 13
8 13 9 2 8 3 8 3 13
24 9 7 0 13 15 13 1 9 2 7 9 0 0 13 3 9 13 2 16 3 15 13 0 9
23 15 13 9 13 3 1 9 2 7 16 9 13 9 9 0 2 13 7 13 9 1 9 13
9 3 9 13 2 3 9 2 3 15
9 3 3 9 9 13 7 13 0 9
20 13 15 2 13 13 2 13 9 0 2 13 0 2 7 15 3 13 2 3 13
18 3 9 15 0 1 15 9 3 9 0 13 2 3 1 0 9 0 13
21 13 15 7 3 13 2 7 13 9 13 9 2 3 0 15 13 2 16 13 1 9
3 3 15 13
11 7 13 3 13 2 13 3 9 2 13 9
6 6 6 2 13 8 8
10 3 16 13 9 2 13 3 0 13 13
6 3 0 13 16 0 9
15 7 13 1 9 9 13 15 0 13 2 15 3 0 13 13
18 7 7 3 9 15 1 9 13 13 2 1 9 0 13 2 15 9 13
28 9 7 0 2 0 9 2 9 0 7 3 0 0 13 9 16 9 0 13 1 9 7 2 15 2 9 13 13
24 7 7 9 2 0 9 13 13 9 9 9 2 7 9 0 9 2 16 13 2 1 9 15 13
13 3 9 13 0 9 9 13 1 9 0 15 3 13
21 13 9 2 16 9 3 3 13 2 9 1 9 13 7 13 13 2 16 1 9 13
16 9 2 0 3 13 9 2 0 9 9 13 7 9 9 3 13
24 7 7 1 9 9 13 2 7 9 3 1 9 13 7 9 9 9 13 7 9 13 15 9 13
14 9 16 13 9 13 2 13 9 7 13 1 9 13 0
18 3 13 15 13 13 9 7 9 0 9 15 3 13 2 7 1 9 13
8 13 3 3 9 9 0 13 13
9 16 15 13 13 13 2 9 15 13
18 15 9 13 13 9 2 15 3 9 15 2 16 15 13 13 9 2 13
16 1 15 9 9 9 13 2 7 13 9 0 1 0 9 9 13
6 15 9 13 9 13 13
9 3 13 13 7 0 9 1 9 13
10 13 15 9 9 7 13 15 13 9 0
12 9 9 13 7 15 9 2 15 13 9 3 13
11 13 15 9 13 9 2 9 13 8 0 13
31 15 7 3 0 9 0 9 13 9 2 7 13 15 9 7 9 1 9 1 9 13 0 9 15 13 3 7 9 7 0 13
15 13 15 9 9 7 15 0 13 9 7 13 2 3 13 13
5 0 13 13 1 15
4 7 6 3 13
12 9 0 9 9 0 0 13 2 15 0 9 13
8 7 13 2 7 9 0 9 13
15 7 3 3 13 2 7 16 13 13 0 9 1 9 15 13
7 3 13 9 15 13 1 9
4 13 13 16 13
14 7 9 13 2 7 16 0 9 2 8 13 2 3 13
12 13 9 13 9 0 7 1 9 0 13 3 9
13 3 1 9 3 3 0 13 2 1 9 15 3 13
10 15 3 0 13 7 6 1 9 13 13
10 15 3 3 9 13 2 16 15 9 13
14 7 16 2 13 2 9 9 13 3 3 9 13 9 13
30 1 9 13 9 0 1 9 7 9 0 7 9 9 7 9 1 9 7 9 0 7 9 7 9 7 9 13 2 9 9
14 7 1 9 13 13 9 2 3 15 3 3 0 9 13
20 3 13 13 15 9 16 9 13 2 16 9 9 13 2 9 1 9 0 3 13
30 3 3 9 9 13 2 15 1 9 13 2 13 15 15 9 2 1 15 9 9 13 9 2 7 13 13 13 15 13 13
16 3 3 13 13 2 3 9 9 0 0 13 9 7 9 13 13
13 3 3 9 13 7 9 9 2 15 1 9 13 13
12 13 15 9 7 13 13 0 7 13 13 9 9
4 3 15 9 13
6 12 3 7 9 13 13
12 7 15 3 0 13 12 3 9 1 0 9 13
14 3 3 2 16 13 13 2 9 13 13 7 13 13 9
18 3 0 9 13 7 9 1 9 13 13 7 9 13 0 9 9 13 0
10 13 9 13 15 2 16 15 13 9 0
8 3 16 9 13 2 9 15 13
9 9 16 3 13 2 0 1 9 13
8 3 15 13 9 13 7 0 13
23 3 9 0 1 15 13 7 0 13 9 2 16 0 9 9 9 13 2 0 9 7 9 9
15 7 16 3 13 2 9 3 13 7 9 9 13 1 9 13
8 6 6 15 13 13 9 1 9
10 13 3 1 9 9 0 9 9 9 13
37 13 3 9 16 0 9 9 13 13 2 13 9 0 9 7 0 13 2 7 9 9 7 9 13 13 7 2 15 3 3 13 2 1 9 0 9 13
9 3 9 13 3 13 15 9 13 13
7 7 16 15 0 13 2 13
6 3 9 9 3 9 13
7 0 9 3 0 13 9 0
21 9 3 2 16 3 13 2 13 9 7 3 13 13 2 7 15 1 9 15 13 13
4 0 3 0 13
13 0 3 9 13 2 15 16 3 13 2 13 0 9
4 0 13 7 13
3 3 9 13
8 3 3 13 2 3 9 0 3
4 15 13 0 9
12 13 13 9 7 3 13 3 0 9 9 0 13
2 9 13
5 7 13 2 9 13
6 13 9 7 13 13 0
8 15 15 13 2 7 6 13 15
4 3 3 9 13
6 13 15 2 7 15 13
17 3 15 0 13 2 16 15 3 13 9 0 13 2 16 3 9 13
6 7 3 15 1 9 13
7 7 13 2 9 2 13 9
24 3 13 13 0 9 2 9 1 9 0 13 7 3 9 9 13 13 13 9 7 0 9 9 13
41 3 3 1 9 13 7 3 9 13 9 13 13 2 3 0 1 9 9 9 13 2 16 9 1 15 9 13 2 7 9 15 13 7 0 0 13 9 2 13 15 9
11 13 13 9 3 9 9 13 2 16 9 13
18 7 15 3 0 13 2 16 3 9 3 0 13 2 16 3 9 13 13
7 13 9 9 3 9 9 13
7 7 13 9 2 16 9 13
14 3 13 9 2 3 9 2 16 15 9 0 1 9 13
5 3 13 13 0 9
9 7 3 9 0 13 13 15 9 0
13 7 16 0 9 13 2 13 15 9 9 9 9 9
8 15 3 13 13 7 13 13 13
10 7 15 9 13 2 16 9 1 9 13
11 3 13 0 9 2 3 15 9 1 9 13
6 3 1 9 3 9 13
18 16 3 9 9 1 13 13 2 0 9 13 13 2 7 0 9 9 13
21 13 15 9 9 13 9 1 13 13 9 7 9 1 9 13 2 15 13 9 9 13
5 15 9 13 0 9
12 1 9 3 0 9 13 7 0 7 0 9 13
5 13 13 2 15 13
22 13 7 9 9 0 13 9 1 0 9 7 9 13 13 2 16 3 9 7 9 9 13
11 3 1 15 9 1 9 7 9 0 13 13
11 3 1 9 13 13 8 3 0 9 9 13
18 3 15 13 1 15 13 9 2 15 1 9 9 13 2 9 7 9 13
22 13 15 9 9 9 13 3 9 9 13 7 3 0 9 13 2 7 16 15 0 9 13
7 3 15 0 3 9 0 13
10 1 9 2 0 15 1 9 0 9 13
16 9 3 9 13 7 9 0 2 9 3 9 7 9 7 9 13
16 7 15 3 0 13 2 16 9 0 3 3 3 15 13 16 0
24 9 13 0 9 13 9 2 16 15 13 9 9 9 13 13 7 0 1 0 1 9 13 9 13
9 13 3 9 15 13 13 2 9 0
7 13 9 0 2 3 15 13
28 3 15 13 2 16 1 9 9 0 9 13 7 9 7 9 7 9 0 9 2 16 15 13 0 9 1 9 13
6 7 3 1 0 13 13
5 15 9 9 3 13
13 3 13 8 8 2 16 9 13 2 16 0 9 13
24 9 0 13 0 9 13 2 7 15 1 9 13 0 1 9 0 12 7 9 1 9 1 9 13
8 13 2 16 15 13 2 3 9
7 13 7 0 9 15 3 13
9 1 9 0 13 9 9 0 9 13
5 7 9 9 13 13
11 7 9 13 13 13 2 7 1 15 9 13
7 9 2 9 9 9 3 13
5 15 9 13 13 13
10 16 13 1 0 9 9 13 2 3 13
1 13
8 15 16 13 9 2 13 13 3
20 13 3 9 2 13 3 9 2 0 3 9 2 3 1 9 13 2 9 9 13
20 3 3 13 3 15 13 2 16 9 3 13 16 13 15 13 13 2 3 3 13
4 3 13 3 9
9 13 15 7 16 13 9 2 3 13
13 13 13 15 7 16 15 9 13 2 15 1 9 13
26 16 15 13 2 13 1 9 9 1 9 13 2 7 9 0 0 15 9 13 2 16 9 3 1 9 13
23 7 7 3 15 3 0 2 15 3 13 13 9 2 16 13 9 13 2 1 15 9 13 13
17 13 15 3 9 2 15 9 0 7 9 13 7 15 13 13 1 0
11 7 9 3 3 3 15 9 0 13 1 9
19 15 3 1 15 13 1 9 2 13 13 2 2 7 2 15 13 9 9 13
25 3 16 13 3 13 1 9 2 16 15 1 9 13 2 13 13 16 13 15 13 15 13 2 15 13
8 9 3 9 1 15 9 13 13
5 0 13 2 0 13
9 15 13 9 0 7 0 9 9 13
6 15 13 3 13 9 13
36 3 3 13 2 16 15 1 9 13 2 7 13 9 2 15 9 1 9 13 13 2 9 13 2 0 3 7 9 0 0 2 1 15 9 0 13
9 7 3 3 3 0 15 9 13 13
12 0 9 1 9 9 13 13 7 9 0 9 13
24 0 7 2 7 2 13 9 9 1 9 13 13 7 13 9 9 1 9 13 7 9 0 9 13
16 15 2 16 9 15 9 13 2 1 9 2 15 9 13 2 13
8 3 8 13 7 3 1 9 13
6 15 13 15 9 0 13
14 15 9 13 9 9 1 9 13 13 7 9 7 9 13
15 3 9 13 1 0 9 7 3 1 9 13 15 9 9 13
13 13 7 13 13 1 9 9 3 15 13 3 3 13
7 13 2 16 9 13 1 9
9 13 3 0 9 2 7 15 3 13
9 13 9 2 3 3 9 0 13 13
25 3 9 2 16 1 9 9 9 13 2 3 13 9 13 7 9 7 9 13 2 15 3 13 9 0
3 3 3 13
9 9 3 13 9 9 1 9 9 13
13 15 3 9 13 2 13 7 9 13 1 9 0 13
9 13 13 7 9 7 13 9 0 13
19 3 9 3 0 9 0 1 9 15 13 2 1 15 13 9 13 7 13 13
15 13 9 3 13 2 7 1 9 15 13 2 9 1 9 13
12 3 9 0 0 13 2 13 2 13 13 9 0
5 13 15 15 3 13
16 7 15 16 0 13 7 13 13 0 2 15 15 9 1 9 13
7 3 2 13 2 15 9 13
16 9 2 13 2 9 15 1 9 0 13 2 16 9 3 9 13
14 3 2 16 13 15 13 9 13 2 13 2 15 13 13
18 1 15 9 9 13 13 2 16 3 13 13 7 2 9 13 15 3 13
5 9 13 2 3 9
17 15 3 9 13 13 7 1 9 15 9 13 13 13 2 16 15 13
14 3 13 3 9 9 7 13 13 9 2 3 9 0 13
9 16 15 8 13 2 1 9 0 13
12 9 13 0 2 3 1 9 2 7 16 9 13
22 12 9 13 2 9 1 9 13 2 8 15 1 9 13 2 9 3 0 13 7 0 9
3 7 9 13
5 3 15 13 2 9
15 13 2 9 0 13 2 9 2 7 15 3 13 13 2 9
4 3 13 9 0
2 13 15
8 15 3 13 2 9 9 13 13
3 7 9 13
9 15 13 2 9 2 16 15 3 13
9 9 13 15 9 13 2 0 9 9
5 3 13 2 3 13
4 0 15 15 13
2 9 13
7 15 7 2 9 2 3 13
6 3 13 2 9 0 13
13 7 2 16 13 13 2 1 15 15 9 9 0 13
21 1 9 2 3 15 13 1 15 13 2 7 16 3 9 0 13 2 9 1 9 13
8 7 3 0 13 2 15 9 13
4 13 2 15 13
7 13 2 16 3 13 1 0
17 3 2 3 0 13 2 9 1 9 13 13 2 7 3 13 9 9
9 9 15 9 13 2 7 13 9 0
5 9 3 15 9 13
2 13 13
4 13 15 15 13
8 0 9 13 2 9 2 3 9
6 0 9 9 3 9 13
3 13 15 13
11 3 6 15 15 9 9 13 2 16 9 9
7 13 2 0 9 0 9 13
11 13 3 9 2 9 2 9 2 9 2 9
6 15 9 9 9 0 13
5 15 13 9 0 9
6 3 13 2 15 9 13
5 0 9 3 9 13
9 3 13 9 0 2 15 9 0 13
6 13 9 2 0 13 9
8 13 15 1 9 7 13 9 13
9 15 15 13 3 15 2 15 13 13
7 1 9 7 9 15 9 13
3 9 0 13
9 0 15 15 3 13 2 15 3 13
5 13 15 3 3 13
5 13 2 13 2 13
7 15 9 0 1 9 15 13
6 15 3 0 1 9 13
6 9 3 15 0 9 13
3 15 9 13
4 3 3 13 9
5 15 15 13 9 0
10 7 16 13 9 9 13 2 3 0 13
8 3 16 9 13 2 13 15 9
5 16 13 2 9 13
3 3 9 13
3 9 9 13
18 1 9 2 0 16 3 13 2 3 13 13 2 7 13 1 9 0 9
9 7 0 9 13 2 15 3 15 13
2 13 15
5 9 13 2 9 13
3 13 2 13
11 3 9 0 2 15 13 9 2 3 13 9
10 9 2 13 9 2 1 15 13 15 13
15 13 7 9 7 1 15 9 9 2 1 15 13 13 9 0
14 3 13 13 9 2 7 3 0 9 7 9 1 9 13
10 7 13 15 13 2 16 0 9 13 13
13 3 13 13 15 13 9 2 16 15 9 13 7 9
4 3 15 0 13
11 15 0 13 13 2 16 0 15 9 3 13
3 13 15 0
4 13 9 0 9
46 0 3 9 9 15 2 15 1 15 0 13 2 3 3 13 2 16 0 13 9 2 3 0 2 15 13 0 9 2 13 13 9 9 2 13 9 3 7 1 9 7 9 13 0 9 13
23 3 13 1 9 7 13 15 0 9 7 15 15 13 7 13 15 1 15 0 9 9 3 3
14 13 1 9 1 0 9 7 13 1 15 9 0 3 9
15 7 13 13 16 13 9 15 13 15 7 13 13 12 9 0
25 7 13 1 9 0 9 12 7 1 9 15 9 0 9 0 13 7 9 15 16 9 13 1 9 0
24 7 16 13 15 13 1 9 15 3 0 7 13 9 0 1 15 13 13 13 15 13 0 7 0
18 7 0 7 13 0 7 3 13 13 1 9 9 7 13 9 9 7 9
13 13 3 15 13 7 15 13 7 15 13 13 1 15
28 13 9 0 7 9 7 9 0 7 16 3 13 13 0 7 13 15 15 15 13 9 7 3 13 7 13 15 0
11 7 9 13 7 13 1 9 0 7 3 13
26 0 13 3 3 13 7 13 9 7 0 9 13 16 16 13 15 7 13 9 0 1 9 0 16 9 13
15 7 9 9 9 13 15 13 0 7 0 15 13 0 7 13
31 9 15 13 15 13 13 6 13 13 9 1 15 1 9 16 13 7 13 9 9 12 13 0 3 1 9 7 13 15 9 9
13 7 9 9 9 13 15 13 15 13 9 0 9 0
7 3 13 3 15 13 9 9
20 7 9 9 9 13 15 13 9 9 15 13 9 16 9 9 7 9 15 0 9
18 13 9 0 7 9 7 9 7 9 7 9 0 7 9 0 0 0 0
14 7 13 15 9 16 9 13 7 3 13 13 1 9 0
24 7 9 15 13 1 9 7 13 0 9 16 15 13 13 9 7 9 7 13 15 0 1 9 0
7 3 15 15 13 13 16 13
10 7 13 15 1 9 0 3 9 9 13
8 15 13 9 13 15 9 13 9
17 13 13 7 13 0 15 13 13 3 16 13 9 0 0 1 9 0
19 7 13 0 9 1 9 15 3 13 9 0 7 13 15 1 0 16 0 13
25 15 13 3 13 9 0 7 3 13 9 15 1 9 9 7 13 9 15 1 9 0 7 1 9 15
8 15 13 9 13 15 9 13 9
24 7 9 9 9 13 15 13 0 7 0 15 13 9 9 15 13 7 9 13 7 13 7 9 13
22 16 13 9 9 0 7 15 15 13 1 9 0 15 13 13 1 9 0 13 13 1 9
8 15 13 9 13 15 9 13 9
17 7 9 9 9 13 15 13 9 9 0 7 0 15 13 9 9 9
17 7 16 0 13 7 7 3 0 7 3 0 13 15 13 1 9 0
28 13 15 13 1 15 9 13 13 16 0 13 7 9 0 13 7 3 13 9 9 0 7 9 13 9 0 16 13
8 15 13 9 13 15 9 13 9
29 1 15 13 7 6 9 13 1 9 7 9 0 15 13 3 9 13 15 13 13 3 7 13 15 15 13 13 1 15
15 3 13 1 9 7 6 9 13 13 1 9 7 1 9 13
19 7 15 13 0 13 9 9 9 7 9 7 9 13 1 9 9 0 9 0
20 7 1 9 13 9 7 9 7 9 7 12 9 13 1 9 15 13 12 9 9
21 13 12 12 9 1 13 1 9 7 13 13 1 9 9 7 13 9 0 1 9 13
24 0 13 9 7 9 0 13 9 7 9 7 9 16 15 13 0 7 1 9 0 13 7 13 13
15 7 13 1 9 13 1 9 9 13 3 7 3 13 9 12
16 7 13 9 0 13 9 0 15 13 0 13 9 7 13 9 15
19 7 9 13 1 9 7 3 1 9 7 3 1 9 13 9 7 3 13 15
15 7 15 13 3 3 9 0 13 13 13 9 7 3 13 15
32 7 13 7 3 1 9 9 7 12 9 7 1 9 9 9 13 3 13 13 9 12 7 9 12 15 13 9 9 13 1 0 9
9 7 13 7 13 1 9 13 1 9
25 7 16 13 9 12 9 7 12 12 9 13 1 9 13 0 9 7 9 0 0 9 15 13 9 9
32 7 13 0 9 13 0 13 13 9 7 13 9 15 3 13 13 7 13 15 9 1 9 0 1 0 9 7 9 7 9 7 9
12 7 13 15 9 0 9 7 9 7 13 1 9
20 7 13 7 13 9 9 0 1 9 9 7 9 7 9 7 13 9 15 9 9
40 7 0 9 15 1 9 13 7 1 9 7 1 9 7 15 13 1 9 7 15 1 15 9 13 13 13 1 9 7 9 9 7 9 7 9 7 9 1 9 9
10 7 12 9 13 3 7 9 13 7 13
34 7 0 13 15 13 9 0 16 9 9 7 9 15 13 2 16 15 15 0 13 2 3 13 0 13 2 15 16 1 0 13 0 9 2
20 15 7 0 9 13 2 9 13 9 9 2 3 15 9 2 0 13 0 13 2
9 3 0 7 1 15 9 13 9 2
16 9 3 2 16 3 2 13 1 10 9 2 15 13 9 13 2
30 9 7 13 9 3 1 9 2 16 3 13 15 13 16 9 2 7 3 13 1 9 2 1 15 13 16 9 9 13 2
8 7 1 15 15 9 9 13 2
14 3 3 9 13 13 16 0 9 15 13 13 16 9 2
17 7 3 2 9 13 9 1 13 1 9 1 9 15 9 13 13 2
16 9 7 9 1 9 15 9 13 2 3 9 13 13 9 9 2
17 9 7 13 0 1 13 16 9 2 3 9 3 13 16 1 9 2
8 3 13 9 0 13 9 9 2
9 9 0 9 1 9 7 1 15 2
9 16 9 0 3 13 1 9 0 2
22 1 13 7 13 16 0 13 9 0 13 1 9 0 2 15 0 13 1 9 7 0 2
17 13 4 3 16 1 9 9 9 13 1 9 2 7 3 1 13 2
21 16 3 9 3 13 0 9 2 9 13 15 7 13 0 9 2 7 13 0 9 2
14 13 7 16 9 15 13 13 9 2 3 13 0 9 2
19 13 3 1 15 9 0 2 16 9 1 9 9 2 9 7 1 9 9 2
13 9 3 13 3 13 0 9 2 7 0 9 13 2
8 3 13 3 1 15 13 9 2
2 3 2
7 9 13 0 16 9 0 2
9 13 3 15 2 16 0 13 4 2
14 1 9 7 9 3 13 9 2 16 3 1 13 4 2
13 0 3 0 1 9 13 2 15 13 1 9 0 2
2 0 2
7 9 13 15 9 9 0 2
10 3 3 0 13 13 0 2 16 0 2
9 9 7 13 13 0 9 7 0 2
8 3 13 3 1 15 13 9 2
2 3 2
10 0 9 13 0 15 15 1 9 13 2
5 13 3 9 0 2
22 15 7 9 3 13 9 1 15 15 13 0 1 15 2 15 13 9 2 7 1 9 2
9 3 13 3 1 15 9 13 9 2
2 3 2
23 0 9 9 13 3 13 1 15 16 13 9 15 9 2 7 1 15 16 13 15 9 9 2
10 9 3 13 0 15 15 13 1 9 2
19 9 7 13 13 1 15 16 9 1 9 13 15 15 9 2 3 0 15 2
9 3 13 3 1 15 9 9 13 2
2 0 2
22 15 3 13 0 16 1 16 13 13 2 3 13 1 15 0 2 7 13 9 1 13 2
12 9 7 13 9 3 13 0 9 16 13 13 2
8 15 3 15 9 15 3 13 2
10 3 13 3 15 9 1 15 9 9 2
25 15 7 13 0 0 2 13 1 15 9 2 16 15 1 15 9 13 2 0 13 15 15 1 15 2
13 3 13 3 15 9 0 9 9 2 15 13 9 2
2 3 2
35 1 10 15 1 15 13 2 13 3 1 3 2 16 0 13 1 0 2 16 2 16 0 13 2 3 0 3 13 2 7 0 0 0 13 2
17 16 3 9 13 13 1 15 0 2 13 16 0 13 15 13 0 2
6 15 7 13 13 0 2
19 3 0 9 15 13 1 9 2 7 13 3 9 0 2 7 0 9 0 2
8 3 13 3 1 15 9 9 2
8 1 15 3 3 13 0 9 2
2 3 2
11 9 9 13 0 1 15 16 1 9 13 2
25 16 3 1 9 13 13 0 9 2 9 9 3 13 0 1 13 1 15 9 16 1 13 1 15 2
6 15 7 13 13 0 2
10 3 9 9 0 13 1 13 1 9 2
5 3 1 15 13 2
9 3 13 3 1 9 13 9 9 2
2 0 2
12 9 0 15 9 9 13 2 16 1 13 13 2
15 15 3 13 0 9 9 13 2 1 15 0 13 1 9 2
37 1 13 7 9 9 13 1 0 9 1 9 2 15 13 1 9 2 15 0 13 9 13 2 3 1 0 0 9 13 2 7 1 13 1 0 13 2
10 3 13 3 1 9 0 9 0 13 2
22 1 15 7 13 9 0 1 15 9 9 9 13 2 1 15 9 13 9 2 8 12 2
24 15 3 13 4 15 0 2 16 13 15 7 13 7 13 9 1 9 10 7 15 13 9 15 2
4 7 8 12 2
5 3 13 9 9 2
12 16 15 13 9 10 2 7 15 13 9 10 2
24 13 3 9 9 15 1 0 9 2 1 9 2 12 9 1 9 0 1 0 9 9 13 13 2
11 3 7 9 2 3 0 2 2 4 13 2
15 13 3 0 7 9 9 2 15 9 0 1 13 9 13 2
6 9 3 13 9 9 2
7 16 9 3 13 1 9 2
17 1 13 3 13 16 7 1 9 13 0 9 9 2 15 13 9 2
19 9 3 0 9 2 7 10 9 2 13 15 9 9 2 16 1 0 13 2
19 9 7 9 3 13 1 10 9 2 7 15 1 15 2 15 15 9 13 2
9 3 13 3 9 9 1 9 13 2
2 3 2
13 15 13 1 15 0 7 0 2 3 13 0 9 2
5 15 7 13 9 2
14 3 3 15 0 13 16 1 15 15 9 1 15 13 2
18 7 1 15 9 13 13 2 3 9 15 15 1 15 13 9 13 13 2
11 3 7 3 13 9 1 0 7 0 13 2
9 3 13 3 1 9 9 9 13 2
2 0 2
6 1 9 1 9 13 2
6 9 7 9 13 0 2
6 15 3 3 13 0 2
13 13 3 9 13 15 9 1 15 9 10 9 13 2
18 15 7 16 9 13 2 3 13 1 9 9 2 7 3 1 9 13 2
9 3 13 3 1 9 9 0 13 2
2 3 2
9 13 0 9 3 13 16 9 13 2
6 13 7 13 3 0 2
9 0 13 3 13 9 0 16 13 2
8 3 13 3 9 0 9 9 2
2 3 2
6 0 9 13 9 9 2
8 9 7 9 3 13 15 9 2
12 15 7 3 13 15 9 2 0 13 13 0 2
10 0 13 3 13 0 15 13 0 9 2
7 13 7 15 0 9 13 2
8 3 13 3 9 0 9 9 2
8 16 9 9 3 13 1 9 2
20 1 15 3 13 16 7 1 9 2 15 13 1 9 9 2 13 0 9 9 2
22 13 3 9 2 1 9 0 1 15 9 1 9 2 7 1 0 2 0 1 9 9 2
19 1 15 7 9 13 13 1 9 7 9 15 2 16 1 15 15 13 13 2
7 4 3 9 1 9 13 2
12 16 3 9 3 13 0 9 2 0 0 9 2
2 3 2
11 0 9 13 1 15 15 13 13 1 9 2
12 15 7 13 1 9 2 3 4 0 9 13 2
24 9 3 3 13 15 15 3 4 0 9 13 2 7 3 9 2 16 9 13 2 1 12 9 2
14 3 13 3 9 13 0 9 2 1 0 1 9 13 2
2 0 2
6 13 0 13 16 13 2
10 3 3 13 16 15 13 0 1 9 2
4 13 7 9 2
17 3 13 3 0 9 9 13 9 2 15 13 1 15 16 15 13 2
2 3 2
8 13 15 3 13 16 1 9 2
6 1 9 7 13 13 2
13 13 3 9 13 7 0 1 0 15 1 15 13 2
5 15 3 13 0 2
17 3 13 3 9 2 15 1 15 13 16 15 13 2 0 9 9 2
2 3 2
10 0 9 13 13 9 2 1 13 9 2
13 9 7 9 2 1 15 9 0 13 2 13 0 2
8 13 3 0 9 7 9 13 2
9 3 13 3 15 9 13 0 9 2
2 3 2
14 15 15 13 0 9 9 2 13 13 0 1 9 0 2
7 0 3 13 0 9 9 2
11 9 7 2 15 1 9 13 2 13 0 2
9 15 3 13 0 9 7 9 0 2
9 3 13 3 15 9 0 9 9 2
8 16 9 9 3 13 1 9 2
12 1 15 7 13 16 7 9 13 0 9 9 2
8 3 3 13 9 16 1 15 2
23 1 15 3 15 9 13 2 7 0 1 13 15 2 7 1 9 9 2 7 1 15 3 2
16 15 7 13 0 9 2 4 1 15 13 2 7 3 1 15 2
8 3 13 3 9 0 9 9 2
2 3 2
19 15 9 7 9 3 13 13 0 9 9 15 0 13 9 1 15 16 13 2
9 9 7 1 15 0 13 16 13 2
6 15 3 15 9 13 2
10 3 13 3 9 9 13 0 9 9 2
2 0 2
10 9 9 0 13 1 16 1 9 13 2
26 3 7 13 0 9 9 7 9 2 15 13 1 9 2 1 15 16 9 13 2 16 1 15 16 13 2
9 3 7 1 15 9 15 9 13 2
9 16 13 3 9 9 1 9 9 2
2 3 2
14 15 1 15 9 0 9 9 13 2 13 13 9 0 2
15 9 7 9 13 0 2 1 13 9 15 1 9 9 13 2
9 3 13 3 1 9 0 9 9 2
2 3 2
7 0 9 9 9 3 13 2
7 3 0 1 9 9 13 2
10 13 7 16 1 9 9 0 9 13 2
9 1 9 7 9 0 9 13 9 2
9 3 13 3 1 9 0 9 13 2
2 0 2
39 15 0 13 1 15 16 9 0 13 2 7 16 0 13 13 2 15 0 13 0 9 13 2 7 16 0 13 2 7 15 3 2 15 1 0 9 13 13 2
8 16 9 3 13 1 9 0 2
35 0 7 7 0 9 0 9 9 13 13 2 1 3 1 15 13 0 9 13 2 7 0 13 2 7 3 13 9 9 2 7 10 0 13 2
10 15 0 9 13 2 16 1 13 13 2
2 3 2
11 9 0 13 0 1 16 1 0 9 13 2
13 1 7 16 13 9 2 3 13 7 0 7 0 2
21 3 3 13 0 10 15 13 9 13 2 7 0 13 15 1 15 16 13 9 13 2
12 0 3 0 3 13 1 15 16 13 13 13 2
2 3 2
6 10 9 1 15 13 2
8 0 7 9 3 13 1 15 2
8 3 13 3 9 0 9 9 2
2 0 2
17 15 15 15 13 7 3 7 0 13 2 3 13 13 0 9 9 2
9 0 3 13 15 15 0 13 13 2
9 9 7 15 3 7 0 13 13 2
7 3 9 0 1 13 13 2
9 3 13 3 9 0 0 9 9 2
2 3 2
12 16 15 9 13 0 9 2 13 15 13 9 2
6 9 7 0 13 0 2
14 13 3 1 9 9 7 9 2 1 15 13 0 9 2
11 7 3 0 13 9 2 3 1 0 13 2
17 15 3 1 15 9 13 2 1 15 1 0 13 2 13 0 13 2
10 3 13 3 1 9 0 0 9 9 2
23 9 3 9 1 15 0 9 13 2 1 10 0 9 2 15 13 9 9 2 1 13 13 2
8 16 9 3 13 1 9 9 2
25 16 7 7 1 9 9 2 3 13 9 2 9 7 9 2 13 9 0 9 2 1 0 0 13 2
18 15 3 3 0 7 0 0 13 2 7 0 13 2 7 9 3 13 2
2 3 2
18 9 13 0 9 2 15 3 13 2 7 13 9 13 2 16 1 9 2
16 9 3 9 2 16 13 7 15 3 2 13 0 16 9 9 2
9 3 13 3 9 9 0 9 9 2
2 3 2
9 15 9 13 9 7 15 9 0 2
7 9 7 13 0 9 9 2
9 3 13 3 1 13 9 9 9 2
2 0 2
12 0 9 2 3 1 9 9 2 13 9 0 2
14 15 3 13 0 9 2 15 0 2 7 3 1 15 2
15 16 3 1 15 13 0 9 9 2 3 13 9 0 9 2
5 15 13 13 0 2
10 3 13 3 9 0 1 9 9 13 2
8 16 9 0 3 13 1 9 2
15 1 15 3 13 16 7 0 9 9 13 1 9 0 9 2
11 3 15 3 9 13 9 7 15 9 0 2
2 3 2
5 9 13 0 9 2
9 9 3 9 13 0 16 9 9 2
9 3 3 0 9 9 1 9 13 2
2 3 2
22 0 9 1 9 13 1 9 7 0 2 1 15 13 13 0 9 2 16 1 9 13 2
6 3 13 7 1 15 2
9 3 13 3 1 9 0 9 9 2
2 0 2
9 9 13 1 9 2 7 1 9 2
9 15 7 9 9 1 9 9 13 2
7 9 7 9 1 0 13 2
27 3 9 9 9 3 13 1 13 16 1 9 1 9 1 9 13 2 1 16 1 9 9 13 9 7 0 2
14 3 13 3 1 9 0 0 9 9 2 15 13 9 2
11 16 0 9 9 3 13 1 9 9 0 2
12 13 7 16 7 1 9 0 13 0 9 9 2
14 9 3 0 3 13 1 0 9 0 2 16 13 0 2
10 10 7 9 0 13 0 1 15 15 2
10 15 13 1 15 15 1 15 13 0 2
16 9 3 9 15 13 1 9 0 2 13 1 9 7 1 9 2
8 0 3 13 1 15 3 13 2
20 0 9 9 13 1 9 1 9 13 2 1 15 16 15 9 15 10 13 13 2
7 7 0 13 1 10 15 2
10 3 13 3 1 9 0 0 9 9 2
2 3 2
17 9 0 1 15 13 16 1 15 13 0 1 9 0 7 0 9 2
27 3 13 7 0 16 9 9 7 9 0 13 0 9 0 9 2 1 15 9 7 0 9 13 1 15 0 2
14 3 13 3 0 16 1 9 9 0 13 0 9 9 2
2 0 2
29 1 9 13 9 1 15 16 13 9 13 2 13 16 0 15 9 2 15 13 9 2 13 1 15 15 13 0 9 2
17 3 7 13 0 9 15 15 1 15 13 2 16 15 1 15 13 2
36 1 3 9 0 9 13 15 1 9 1 9 15 1 15 13 2 3 13 13 0 9 2 15 13 9 2 7 3 9 15 13 1 15 9 9 2
2 3 2
13 13 4 1 16 9 10 9 0 13 13 1 9 2
13 15 3 1 15 9 0 13 9 2 13 15 9 2
18 15 7 3 13 1 9 0 2 1 15 9 9 13 3 13 16 0 2
17 3 3 9 13 13 9 2 7 15 3 2 1 15 13 9 0 2
18 3 13 3 0 9 9 2 15 13 0 15 9 2 13 1 9 0 2
2 3 2
6 9 13 0 9 9 2
24 15 3 15 13 0 0 9 1 10 9 0 9 15 9 2 13 1 15 13 13 15 0 9 2
8 3 7 3 13 9 0 9 2
18 3 15 9 15 13 7 9 7 9 2 0 7 9 15 9 15 13 2
10 3 13 3 0 9 9 1 9 0 2
9 16 0 9 3 13 1 9 9 2
14 1 15 3 13 16 7 1 9 9 13 0 9 9 2
12 9 3 9 13 0 1 15 15 13 0 9 2
11 3 13 7 1 9 0 9 0 9 9 2
6 7 3 1 9 9 2
2 3 2
9 0 9 9 13 1 0 9 9 2
19 0 7 9 9 2 1 15 15 13 0 9 2 13 1 9 1 9 9 2
12 9 7 9 3 13 1 9 9 9 7 9 2
11 3 3 13 1 0 2 7 1 13 0 2
10 3 13 3 1 15 9 0 9 9 2
2 0 2
14 15 13 1 15 16 1 9 2 3 13 0 9 9 2
51 9 7 9 13 1 15 16 1 9 2 3 16 10 0 9 2 1 15 13 9 2 13 1 9 2 7 3 16 9 13 9 3 15 13 1 15 15 13 1 9 13 2 16 13 1 9 2 1 12 9 2
10 3 13 3 1 9 9 0 9 9 2
2 3 2
14 9 0 3 13 15 9 2 16 13 9 1 12 8 2
15 13 7 15 15 15 9 2 16 13 1 15 1 12 0 2
8 3 9 3 13 1 9 9 2
8 16 9 3 13 1 9 9 2
8 13 3 16 7 1 9 9 2
7 16 3 9 9 0 13 2
13 7 3 1 9 13 2 7 15 3 13 0 9 2
2 3 2
6 9 9 9 13 9 2
17 15 3 13 13 0 9 0 9 2 1 3 15 13 9 10 0 2
7 10 3 1 9 9 13 2
10 3 13 3 1 9 9 13 0 9 2
9 16 0 9 9 13 1 9 9 2
61 16 3 0 9 9 3 13 1 0 2 15 13 9 9 2 7 1 9 9 2 7 1 9 9 3 1 0 9 2 7 3 1 0 1 9 0 9 2 7 1 0 15 1 9 13 2 3 9 7 9 2 13 16 0 9 9 13 1 9 9 2
19 15 3 0 9 9 13 15 0 2 7 1 15 15 9 15 15 9 13 2
17 15 3 1 15 15 13 16 1 9 2 1 9 9 1 15 13 2
25 1 15 3 9 9 10 0 13 1 9 2 16 15 3 1 9 0 1 9 7 1 9 13 13 2
13 15 3 9 1 15 0 13 2 13 15 15 9 2
20 1 15 3 9 15 9 3 13 0 2 3 1 15 1 9 9 0 9 13 2
13 1 15 3 10 15 0 9 13 13 16 1 9 2
19 1 9 3 9 13 9 9 2 1 15 13 0 10 15 13 0 1 9 2
31 13 3 9 1 9 9 2 1 15 13 1 9 0 7 1 9 2 7 9 1 0 9 2 1 15 13 15 9 9 0 2
15 16 3 2 16 13 13 2 10 0 9 13 13 13 9 2
50 3 13 7 0 16 0 9 9 13 1 9 15 13 1 9 9 2 15 13 0 2 16 0 0 2 9 9 1 9 13 2 7 13 9 2 3 9 0 9 2 1 9 15 13 2 3 1 9 9 2
23 7 3 1 9 15 13 1 9 9 2 1 13 9 13 1 9 9 1 9 1 0 0 2
15 13 3 16 1 9 9 0 9 9 13 2 1 0 9 2
23 1 15 3 13 9 9 15 1 9 4 13 2 16 0 9 9 3 13 16 1 9 9 2
14 7 9 2 1 13 9 2 3 13 9 1 15 9 2
39 1 0 13 16 9 15 13 9 0 2 3 13 9 15 0 10 9 7 10 9 2 7 9 13 1 9 9 1 9 1 9 2 7 13 9 13 15 9 2
14 1 0 13 16 10 9 13 10 9 1 9 9 15 2
34 9 7 9 3 13 9 9 2 7 13 15 2 16 9 9 13 9 9 2 7 3 13 9 1 9 2 7 13 9 2 15 13 9 2
14 7 9 2 1 13 9 0 2 3 13 9 1 9 2
14 0 2 3 9 9 13 1 9 2 16 0 1 9 2
15 3 9 0 1 0 13 1 9 2 7 13 1 9 0 2
23 0 0 2 10 9 13 1 9 15 2 16 7 9 1 9 2 9 3 13 3 9 15 2
33 3 7 15 15 13 1 9 2 13 0 16 15 15 13 7 13 15 2 16 13 16 13 2 7 13 16 13 2 7 9 16 9 2
28 7 3 3 13 2 1 0 13 2 0 13 9 1 10 9 2 16 7 9 2 13 0 9 2 13 0 9 2
8 13 16 9 9 13 1 9 2
24 13 3 9 2 1 9 1 8 2 16 1 9 15 13 1 9 2 13 9 15 13 1 9 2
22 9 7 15 13 1 9 2 13 9 0 2 9 7 15 13 1 9 2 13 9 9 2
8 3 9 9 13 1 0 9 2
15 7 0 9 1 10 9 13 9 2 9 7 0 13 9 2
10 3 9 0 9 4 1 0 9 13 2
17 7 9 0 13 9 1 15 9 2 3 13 13 9 7 9 9 2
14 3 0 3 1 0 9 9 15 13 1 9 2 13 2
12 3 3 9 0 13 1 9 2 7 1 9 2
18 13 13 16 9 13 15 16 10 9 0 13 1 9 0 15 9 13 2
24 9 3 13 9 15 13 1 9 0 2 13 7 13 1 9 1 9 13 2 1 9 9 15 2
45 13 3 9 15 0 13 2 7 0 9 2 7 3 1 15 2 1 15 13 15 0 0 2 1 16 1 9 0 13 15 9 1 15 9 13 2 1 9 9 15 2 15 9 13 2
26 7 1 9 9 13 0 9 9 13 2 13 16 12 9 13 13 15 13 9 2 15 13 9 10 9 2
21 9 0 7 15 15 3 13 9 9 0 1 9 1 15 13 2 7 0 1 9 2
43 1 9 3 1 9 9 0 13 2 15 3 15 9 2 15 7 9 13 2 2 13 13 10 9 15 13 1 9 0 2 16 1 9 15 13 1 9 9 2 13 9 9 2
13 13 3 9 9 2 7 16 15 9 13 1 15 2
67 7 16 13 9 1 12 8 2 15 15 0 13 2 13 9 2 9 7 0 9 13 16 3 13 2 3 3 13 2 1 15 16 15 13 7 13 2 7 9 13 7 13 2 16 3 9 3 13 9 2 7 9 13 9 1 15 2 3 3 15 13 13 2 16 7 9 2
20 7 3 2 1 0 13 1 10 0 2 3 13 13 9 9 0 15 9 0 2
27 3 3 9 0 13 2 3 3 13 1 15 0 9 2 7 3 9 13 1 9 1 9 1 15 9 13 2
22 13 0 16 3 9 0 1 9 0 13 2 3 16 13 9 2 7 16 13 1 9 2
24 0 7 13 1 9 2 16 1 0 9 2 3 9 0 9 2 15 13 15 0 9 0 9 2
28 7 3 9 0 15 1 0 9 9 13 2 4 0 1 9 13 2 15 0 1 9 13 9 2 16 0 9 2
25 1 15 13 9 9 1 9 9 13 2 1 15 2 1 9 2 13 10 9 7 9 7 9 9 2
44 1 0 3 13 16 9 13 1 9 15 13 1 9 2 9 9 15 13 1 9 0 2 16 3 9 13 2 8 12 2 9 13 13 4 9 9 9 2 16 1 0 0 13 2
32 16 3 1 9 15 13 1 9 2 13 9 2 13 13 16 1 15 13 9 15 13 1 9 2 3 1 9 2 7 1 9 2
63 1 0 13 16 9 13 1 9 13 2 3 1 9 15 1 15 0 9 15 2 16 0 13 2 7 1 9 0 7 9 0 2 1 15 1 9 13 2 7 0 1 9 9 0 2 1 15 3 9 9 4 9 13 13 2 16 1 9 1 9 13 13 2
18 1 0 13 16 9 0 13 9 1 15 9 2 3 13 2 7 13 2
9 3 13 13 16 9 13 1 9 2
10 9 3 13 9 9 1 9 10 9 2
9 15 7 15 13 9 2 13 9 2
18 13 3 9 13 1 9 2 13 13 9 9 1 9 2 15 13 9 2
20 7 3 13 13 16 13 15 9 0 7 3 13 15 9 0 2 15 4 13 2
56 16 1 15 9 13 13 9 1 9 1 9 9 2 7 13 9 15 15 2 13 16 13 9 3 13 0 9 9 2 7 9 9 15 2 15 13 0 9 0 2 7 3 13 9 13 9 2 1 15 3 13 9 2 7 9 2
24 3 13 13 16 9 0 7 4 13 3 1 9 2 7 1 9 12 0 2 7 1 9 13 2
52 7 3 2 16 9 9 13 1 9 0 9 2 15 1 15 3 13 15 9 2 9 9 3 13 9 7 9 15 9 2 16 9 13 2 7 9 7 9 3 2 15 9 15 9 13 0 9 2 7 9 15 2
28 15 0 0 13 9 2 3 1 16 13 10 9 2 7 1 16 13 15 9 7 9 15 3 13 1 0 9 2
10 13 3 9 1 9 2 16 13 9 2
11 7 1 9 2 16 13 0 13 0 9 2
47 1 15 3 2 13 9 0 7 0 2 7 0 7 0 2 16 9 1 9 13 2 3 1 15 13 13 0 7 0 2 2 7 15 9 1 9 13 2 3 7 9 9 13 13 9 2 2
26 1 0 13 16 9 2 1 13 9 2 13 9 15 2 9 7 1 15 15 13 2 13 9 1 9 2
15 3 3 13 13 1 9 9 1 9 2 16 9 1 9 2
17 0 2 9 9 3 1 9 10 2 1 15 16 13 9 7 9 2
10 7 10 9 13 12 9 2 3 9 2
6 7 9 13 1 9 2
23 7 3 13 15 9 9 7 9 0 2 9 13 12 9 10 9 2 13 1 9 9 0 2
24 7 16 9 9 13 12 9 1 15 2 15 13 15 9 2 15 9 13 2 13 9 15 13 2
41 16 15 9 0 9 13 2 7 3 1 15 13 10 9 0 2 7 9 13 1 9 13 9 2 15 3 13 9 0 2 7 1 15 2 16 9 13 15 9 9 2
30 13 7 16 15 9 15 13 1 9 0 13 16 13 9 7 9 2 13 1 9 16 3 13 15 9 9 0 7 0 2
14 9 3 2 1 15 15 13 2 13 1 9 1 9 2
21 13 3 16 9 2 1 15 13 2 13 1 9 1 9 10 15 15 13 9 0 2
14 1 12 7 9 3 13 1 9 16 3 1 15 9 2
10 13 3 1 9 3 1 10 15 9 2
17 7 15 13 2 16 12 15 9 13 9 7 13 1 15 9 15 2
35 16 9 2 3 13 1 15 2 0 15 13 1 9 7 0 2 3 16 16 13 1 9 0 2 13 1 9 1 9 13 2 3 1 0 2
21 3 3 9 2 1 16 13 1 9 0 9 2 13 3 1 9 1 9 0 9 2
30 7 1 3 13 15 1 9 2 13 3 1 9 7 9 2 16 9 9 1 15 15 13 1 9 1 9 2 13 9 2
12 7 9 15 13 9 13 15 13 15 16 9 2
23 16 0 13 13 15 9 9 2 16 7 15 15 13 9 7 9 2 7 13 9 7 9 2
35 13 3 1 9 9 13 15 13 9 2 16 9 0 3 13 13 9 2 15 13 13 1 9 7 9 9 2 13 16 13 15 9 7 9 2
21 13 3 16 9 9 0 2 1 15 13 2 3 13 1 9 16 1 9 15 13 2
27 3 15 9 3 13 15 9 2 16 15 9 1 15 13 9 1 9 2 7 1 3 3 2 16 9 13 2
27 1 0 13 16 9 9 3 13 12 1 10 9 2 1 3 13 15 1 9 15 9 13 2 16 13 4 2
22 3 1 15 15 9 0 9 13 15 1 9 9 2 16 3 13 1 9 1 9 9 2
27 16 3 9 13 9 2 16 9 13 1 9 9 2 13 16 9 9 13 2 7 16 9 15 13 15 9 2
11 7 9 0 9 13 9 0 1 15 9 2
16 3 9 3 13 15 9 0 2 7 3 0 9 2 7 0 2
10 15 0 13 16 9 13 9 0 9 2
27 0 3 2 16 15 9 0 13 1 15 0 2 16 15 15 13 13 9 9 2 16 13 1 12 1 9 2
30 0 2 16 0 13 16 15 15 13 9 0 1 12 2 13 9 0 1 15 2 16 9 0 1 15 13 13 1 9 2
15 9 7 3 13 9 0 9 2 3 2 15 13 2 13 2
8 3 3 13 13 9 0 9 2
39 13 13 3 16 2 16 9 13 9 0 13 9 0 9 2 3 9 13 9 0 13 9 0 9 2 7 15 15 9 1 15 13 2 16 15 15 15 13 2
27 1 0 3 13 16 2 1 9 13 9 0 2 9 15 13 9 1 9 9 2 16 15 13 1 9 9 2
14 1 3 9 9 13 9 2 0 13 3 9 13 9 2
21 1 0 9 0 13 0 2 1 9 15 2 9 13 13 3 3 2 7 3 3 2
20 7 9 3 13 1 15 9 9 1 9 9 0 2 16 13 3 9 15 9 2
48 1 0 13 16 2 16 9 13 1 9 9 3 0 1 9 9 0 2 3 9 13 3 0 1 9 9 0 1 13 9 0 2 7 1 15 16 13 9 0 9 2 16 13 9 0 9 0 2
25 3 3 13 9 0 9 13 2 16 0 1 9 9 13 9 2 16 0 9 9 2 7 16 0 2
28 1 0 3 13 16 2 1 9 15 13 9 9 9 13 9 2 13 13 16 9 1 9 4 13 1 9 0 2
36 7 15 3 13 3 13 2 16 13 9 9 3 13 1 9 12 9 2 7 13 0 1 9 16 1 15 2 9 15 3 13 13 1 15 9 2
27 9 7 9 13 1 9 9 2 1 15 15 13 9 9 9 13 9 2 16 9 9 13 15 0 13 9 2
32 16 9 2 1 13 1 10 9 0 2 13 9 15 3 13 13 15 9 2 3 0 13 16 9 4 13 1 9 0 9 13 2
37 13 3 0 13 9 0 0 2 7 9 0 1 10 9 2 15 13 0 13 9 9 7 9 2 2 3 16 15 9 9 13 9 2 7 9 3 2
19 1 15 13 9 9 0 1 9 0 2 3 0 13 9 2 7 9 3 2
18 9 0 9 13 9 9 0 1 9 0 2 3 9 2 7 9 13 2
42 3 1 15 15 13 2 13 9 2 7 13 0 2 13 16 9 0 13 4 9 0 9 2 1 15 13 15 15 9 2 7 9 0 9 2 1 15 13 15 3 13 2
43 7 9 9 2 1 15 2 3 13 9 10 9 16 3 13 9 7 9 7 9 2 15 12 13 16 0 9 0 2 2 7 13 9 9 9 13 9 2 7 13 15 9 2
46 1 0 3 13 16 2 1 9 2 3 1 9 0 9 3 13 9 9 9 2 16 1 13 9 2 16 13 16 0 9 2 3 0 9 2 7 0 9 2 13 9 1 9 7 0 2
9 9 0 9 9 13 0 7 0 2
34 7 3 1 9 9 7 9 0 2 9 15 9 13 2 9 3 13 0 13 2 9 0 13 2 16 15 13 1 12 1 8 1 8 2
49 15 0 3 15 13 16 3 9 9 9 13 12 1 9 9 11 0 7 0 15 9 0 1 9 13 0 1 9 9 11 0 15 13 1 9 7 9 0 9 11 7 9 11 15 9 15 1 9 13
34 1 0 9 13 11 11 9 0 15 9 9 1 9 0 9 13 7 1 9 9 0 9 13 13 16 9 1 9 15 13 15 9 3 13
7 1 15 16 9 13 15 13
17 12 1 9 0 7 0 1 9 11 7 9 11 3 3 0 9 13
22 9 0 3 0 13 9 9 13 13 3 1 11 0 9 12 9 15 13 1 11 13 13
33 3 0 9 15 13 1 9 13 7 9 1 15 13 13 15 9 7 9 9 0 13 9 15 1 9 13 7 16 9 13 13 13 13
36 15 1 11 0 9 13 12 7 3 9 13 7 12 15 1 11 13 1 9 13 7 3 0 9 1 0 11 1 11 13 1 0 12 9 13 13
22 0 9 15 9 9 9 7 9 9 11 0 13 15 13 9 3 3 1 9 9 9 13
9 3 15 9 11 1 12 9 13 13
14 16 9 13 13 13 7 0 9 9 9 7 0 9 9
17 16 15 9 3 3 13 16 7 3 3 15 3 9 13 13 0 13
22 15 9 13 9 16 12 9 0 9 9 13 3 13 3 3 7 0 9 9 15 13 13
10 3 3 11 9 11 13 15 3 13 13
4 13 3 7 3
12 16 15 13 9 0 1 9 1 9 9 13 13
14 11 0 1 9 11 13 13 13 16 15 0 1 9 13
4 11 1 15 13
22 1 0 9 11 11 9 1 9 1 12 9 7 15 9 15 9 13 0 9 9 13 13
27 0 3 9 1 9 11 13 7 9 1 15 13 7 9 9 13 7 11 9 13 15 3 13 1 13 15 13
18 9 9 7 1 12 9 13 7 15 1 15 15 1 0 9 13 13 13
17 9 9 3 13 0 7 0 9 16 13 7 13 13 0 16 13 13
20 1 9 9 9 0 13 16 7 1 9 9 7 1 9 13 15 15 13 3 13
5 13 1 9 9 13
9 1 0 15 9 13 13 3 12 12
10 0 9 13 15 15 13 11 1 9 13
11 1 0 9 0 7 9 3 7 3 9 13
5 9 13 0 0 0
72 16 1 0 3 13 3 7 15 3 9 13 13 0 11 0 13 0 13 0 7 0 9 9 3 0 16 0 3 1 0 3 13 3 7 9 13 13 0 7 11 9 3 16 3 13 13 3 16 0 3 9 9 13 9 3 15 1 9 15 11 13 15 9 15 1 9 15 13 15 9 13 13
12 13 15 1 9 0 7 0 15 9 1 15 13
13 3 7 9 9 13 3 7 0 9 7 15 9 13
11 16 15 3 13 3 15 0 9 9 0 13
23 15 9 11 3 13 13 15 13 16 16 0 9 9 1 0 9 11 15 13 3 3 13 13
24 0 3 13 13 1 9 9 9 0 7 15 1 9 9 9 11 13 3 0 1 9 0 9 13
31 0 16 13 13 9 15 7 9 1 0 9 13 9 3 15 13 3 16 7 15 1 9 7 15 9 13 15 13 7 13 13
30 3 0 13 0 9 15 1 3 9 9 13 3 3 1 15 7 3 1 0 9 3 13 15 3 0 13 15 9 3 13
9 15 9 0 9 9 9 9 13 13
8 13 11 9 11 9 1 15 13
17 15 16 13 3 3 15 1 9 0 9 13 3 3 13 13 11 13
13 15 9 7 0 13 7 1 0 9 9 13 13 13
11 3 1 0 9 0 7 9 9 0 7 13
19 16 1 9 0 9 13 7 9 13 3 3 3 15 13 9 0 9 3 13
48 16 9 1 9 9 13 13 3 15 3 0 3 7 3 0 13 9 16 3 13 3 7 9 9 0 9 9 9 13 3 7 15 1 0 9 15 9 15 1 7 1 9 13 9 9 0 13 13
16 16 9 9 13 13 0 13 13 11 15 9 13 15 9 13 13
15 9 1 15 15 0 1 9 1 15 13 7 9 0 13 13
7 11 0 15 9 9 9 13
19 16 3 13 3 13 7 3 13 0 13 0 9 9 16 9 13 9 9 13
11 3 3 11 9 15 9 15 9 0 13 13
18 3 9 13 15 1 9 13 9 13 9 13 13 16 15 1 9 9 13
26 3 9 13 13 7 15 9 9 13 3 7 3 13 13 3 1 9 11 12 9 1 0 9 3 12 13
18 15 15 0 1 15 3 9 13 13 3 9 3 13 7 1 15 9 13
4 13 0 13 9
9 3 3 13 3 13 16 1 15 13
19 0 13 13 0 12 12 13 1 0 9 13 12 12 0 7 9 9 15 13
20 11 9 13 3 7 9 13 15 9 1 15 13 9 7 9 9 1 15 13 13
12 9 1 9 9 12 9 9 7 12 9 13 13
9 16 9 15 13 15 3 13 3 13
8 9 3 15 9 1 9 13 13
6 3 1 0 9 13 13
13 0 9 13 9 1 9 15 9 15 0 9 13 13
12 9 13 9 13 15 7 1 13 9 13 13 13
14 15 0 9 9 13 16 13 15 9 9 13 1 11 13
20 15 13 9 0 7 9 1 9 13 13 16 0 9 13 9 15 7 13 9 13
12 0 9 13 9 9 7 13 15 9 9 0 13
9 1 0 9 1 9 0 9 9 13
42 3 0 9 15 9 1 15 15 1 9 0 13 13 13 15 9 1 15 13 9 13 16 1 9 9 9 7 13 7 0 15 13 3 15 9 13 9 7 1 15 9 13
2 9 13
23 15 15 1 9 1 9 9 13 15 7 0 9 13 1 0 13 16 1 13 15 13 9 13
31 7 9 15 1 0 9 7 0 9 9 15 9 9 13 13 13 9 13 16 13 7 9 1 15 9 13 13 0 9 15 13
30 15 16 1 9 7 9 9 15 1 9 9 13 3 7 1 9 7 9 7 9 7 9 13 13 15 1 9 15 0 13
25 15 16 1 15 1 9 9 0 9 9 7 13 12 1 9 3 0 9 1 9 3 3 9 12 13
48 3 3 13 7 13 9 13 0 7 0 9 13 9 1 11 1 9 13 15 1 0 9 13 3 15 13 9 1 0 0 9 13 15 0 9 9 0 9 13 13 15 15 7 15 15 9 13 13
19 1 9 11 9 13 9 7 1 9 13 13 16 15 3 9 1 9 9 13
23 15 1 9 9 9 15 7 9 0 0 9 13 3 9 13 9 1 9 13 1 11 13 13
37 16 9 9 0 13 9 7 3 13 13 3 1 9 0 13 13 1 0 9 9 15 9 13 15 3 13 9 7 15 13 1 0 9 9 7 9 13
30 15 9 1 15 1 9 13 15 13 7 3 3 13 1 9 13 7 3 0 3 0 9 3 13 13 7 15 13 9 13
12 11 11 9 1 9 0 0 9 11 1 11 13
39 9 0 7 3 9 13 11 9 3 16 15 1 15 9 13 13 1 9 9 9 13 7 3 0 15 1 9 9 13 13 13 0 0 9 16 3 9 9 13
27 0 13 9 0 7 9 13 7 1 9 13 9 7 15 9 1 9 13 13 16 1 9 9 9 13 13 13
28 0 3 3 0 9 9 13 16 15 9 9 13 0 7 13 0 7 0 9 0 9 0 7 3 15 9 9 13
28 3 7 3 0 15 9 13 13 0 1 0 13 9 3 7 1 9 3 9 13 7 0 1 9 3 3 9 13
16 0 16 9 15 9 1 9 13 13 13 7 13 9 9 13 13
10 15 9 9 9 0 7 9 0 13 13
25 0 7 3 9 3 1 11 0 9 9 7 13 15 9 13 9 7 13 1 9 9 7 0 9 13
35 0 9 1 0 9 9 13 0 9 11 9 9 9 9 9 15 9 3 3 1 15 13 13 9 0 9 7 16 3 3 9 0 15 13 13
9 0 9 13 0 15 1 9 13 13
6 3 13 9 9 9 13
12 9 9 7 13 11 1 9 9 7 9 13 13
18 0 9 13 15 9 0 9 13 9 1 0 9 13 15 9 9 13 13
26 15 9 0 9 13 1 12 12 9 15 1 11 9 7 13 13 3 0 9 13 0 9 15 1 9 13
36 0 3 9 11 9 13 13 7 16 15 0 0 7 9 1 9 9 13 13 15 0 9 15 13 13 13 1 9 13 7 1 9 1 15 9 13
3 0 3 13
12 3 7 15 9 0 15 7 0 13 3 9 13
6 15 0 9 9 9 13
14 15 9 13 11 16 0 9 13 3 16 13 1 9 13
10 16 15 9 0 13 13 15 0 13 9
23 7 13 16 13 1 9 9 13 15 13 9 1 15 7 1 9 9 13 7 1 15 9 13
26 16 0 3 13 13 16 1 15 9 15 9 13 13 15 7 9 13 15 7 16 9 13 1 9 9 13
10 1 0 9 1 9 15 13 12 7 12
8 15 15 11 13 13 0 13 13
22 15 1 12 15 0 0 13 1 0 9 9 16 9 9 9 12 12 13 15 1 9 13
25 9 3 15 0 1 0 1 11 9 13 9 13 9 13 3 13 16 15 9 13 16 3 1 9 13
17 9 0 0 3 1 0 0 13 1 9 9 9 9 12 1 15 13
13 15 9 7 9 13 3 13 9 7 1 15 13 13
26 3 7 3 3 1 9 3 13 15 3 7 0 0 15 1 9 0 7 0 9 15 13 1 11 0 13
28 11 13 9 15 3 15 9 13 13 15 9 13 7 15 9 13 3 13 12 9 1 11 13 15 7 3 13 13
25 0 13 9 13 0 1 13 9 0 3 9 13 9 7 1 0 9 13 7 9 13 7 15 13 13
41 15 3 11 13 9 0 15 7 9 13 9 0 7 9 1 9 0 3 13 1 0 9 7 9 13 7 1 9 0 9 13 7 3 9 9 9 9 13 7 13 13
28 15 3 16 3 7 9 13 3 7 3 13 3 7 9 13 13 7 15 15 1 9 15 9 13 15 13 3 13
9 9 15 13 15 7 13 13 13 13
41 15 16 13 11 7 1 9 13 0 9 3 13 13 16 15 15 9 13 13 7 15 3 3 13 13 13 15 1 0 9 9 15 13 3 9 9 0 15 1 9 13
6 3 1 15 9 9 13
31 3 1 15 9 13 7 9 13 7 0 9 9 7 9 9 9 3 13 7 16 15 1 9 9 13 1 9 13 7 9 13
29 3 9 9 1 15 9 13 9 7 15 9 15 13 7 15 9 13 7 1 0 15 13 9 13 16 9 9 13 13
17 7 1 0 0 12 0 9 15 0 13 3 13 7 3 3 13 13
7 11 1 9 15 9 9 13
11 0 15 13 9 1 13 9 1 11 13 13
34 13 9 7 15 15 9 13 15 13 13 13 7 15 1 9 11 13 13 15 1 9 0 1 11 9 13 13 3 12 9 12 9 1 9
24 15 3 1 15 13 7 1 15 13 13 16 3 9 1 9 13 16 15 9 9 9 1 9 13
13 3 9 0 11 13 9 12 12 0 7 1 15 9
11 9 13 3 1 9 13 16 11 15 9 13
20 15 9 13 11 13 9 7 15 9 13 0 9 9 1 15 13 13 13 7 13
11 13 11 3 13 1 15 0 1 9 9 13
15 0 13 15 9 9 7 9 9 13 7 1 0 9 13 13
3 0 13 9
18 0 13 9 0 9 9 1 11 1 9 13 12 7 1 15 9 13 13
4 15 1 9 13
32 11 9 9 9 0 7 9 13 15 15 13 9 13 7 16 3 9 9 13 9 0 9 7 9 3 9 0 13 9 9 13 13
8 3 15 9 13 9 1 9 13
14 0 13 9 3 1 0 9 15 3 9 13 13 9 13
30 3 0 3 9 13 1 9 0 9 15 1 12 9 9 13 7 0 9 15 1 15 13 9 13 16 9 9 9 7 13
23 16 1 0 9 13 13 3 0 13 13 1 11 11 7 9 7 3 13 0 9 1 15 13
14 15 9 13 11 9 13 9 11 1 9 13 0 9 13
17 0 16 7 9 0 7 9 9 7 9 0 13 15 1 9 13 9
10 15 3 13 13 0 9 0 7 9 13
24 9 1 11 13 7 3 1 11 13 13 13 7 3 15 3 15 9 13 13 3 3 13 9 13
25 0 3 1 9 7 15 9 1 9 7 9 9 1 9 9 1 9 0 9 7 9 13 7 9 13
4 9 3 11 13
12 16 13 9 13 13 0 7 9 1 12 9 13
13 15 15 9 13 1 15 9 15 1 9 0 9 13
6 9 3 1 0 9 13
22 15 9 15 13 9 16 7 3 1 9 13 7 9 7 0 9 9 13 0 9 9 0
18 1 9 15 13 0 9 7 9 9 7 9 1 15 9 13 9 7 13
29 3 15 15 0 11 13 9 1 11 9 15 11 7 15 9 9 0 13 13 15 0 11 13 9 9 13 7 3 13
26 3 7 15 13 0 11 15 15 7 13 1 9 0 9 13 16 9 9 12 13 7 15 1 9 13 13
5 0 13 9 1 9
26 0 15 9 13 9 7 0 9 9 13 7 15 0 1 0 13 13 1 0 9 15 13 9 0 13 9
4 15 3 13 13
11 3 7 1 13 9 7 1 13 3 9 13
18 11 13 9 9 9 16 15 1 15 9 1 9 13 1 15 16 13 13
14 11 11 1 0 9 9 1 0 9 15 9 13 13 13
16 16 9 13 9 7 9 9 13 13 13 0 9 13 7 13 9
14 1 11 1 9 13 9 13 9 7 3 15 1 9 13
8 13 3 13 15 7 9 13 13
14 0 3 9 9 0 9 9 15 1 9 13 13 9 13
9 15 13 9 7 9 9 9 13 13
4 3 3 9 13
5 15 1 0 13 13
14 16 3 0 13 9 16 9 15 13 13 3 0 13 13
22 9 13 9 9 16 15 3 13 1 9 13 1 0 9 15 1 9 13 1 11 15 13
34 9 3 3 1 0 9 9 7 9 13 7 3 9 9 7 9 13 16 16 15 3 1 9 15 13 3 0 13 9 9 15 9 13 13
4 13 12 11 11
14 11 3 13 15 13 7 13 9 7 0 15 9 0 13
33 15 1 15 9 0 13 0 13 9 7 3 16 13 1 9 3 13 11 16 11 1 9 9 13 13 9 0 9 1 11 16 0 13
6 3 0 0 13 1 9
16 3 3 0 13 16 0 0 1 0 0 13 15 15 3 13 13
17 9 15 3 15 13 7 13 3 3 13 16 0 9 15 8 13 13
6 15 9 15 9 13 0
4 15 15 3 13
7 11 11 11 11 9 11 13
7 15 9 13 7 13 7 13
6 11 16 3 13 13 13
8 1 9 9 1 9 1 15 13
11 15 3 13 13 1 15 13 9 15 13 13
18 7 15 7 9 15 7 9 3 13 9 7 15 0 13 3 11 9 15
18 15 13 16 15 9 8 13 13 15 9 13 0 15 15 3 13 16 13
4 1 11 13 13
9 16 11 9 3 13 15 15 13 13
4 11 9 15 13
31 9 15 7 9 3 13 16 3 13 13 13 7 16 15 15 8 0 9 15 3 13 13 7 3 15 15 9 9 7 13 13
15 3 0 9 15 13 13 16 15 9 9 1 0 9 13 13
14 7 0 7 13 16 13 7 15 0 13 1 15 9 13
12 11 0 0 3 9 3 7 11 1 9 3 13
27 9 15 9 13 16 15 3 7 1 0 3 7 1 0 9 3 13 9 13 3 7 15 13 15 7 0 13
9 13 15 3 0 16 13 15 9 13
9 16 9 15 13 15 1 9 13 13
10 13 3 16 15 3 16 15 1 11 13
5 9 3 3 9 0
18 3 9 1 9 9 1 9 7 1 9 13 0 7 1 15 9 13 13
2 15 0
5 15 8 8 8 0
4 3 3 13 13
4 15 15 1 15
3 3 0 0
24 3 11 8 8 13 13 9 7 9 15 15 1 9 0 13 3 7 13 13 13 7 15 0 9
10 15 3 0 9 0 3 8 0 9 11
2 15 0
5 0 3 9 11 13
21 9 7 1 9 9 7 1 9 7 1 0 9 13 16 16 9 13 13 16 15 13
2 15 13
6 11 11 0 9 13 13
5 13 15 8 8 8
16 3 16 9 13 9 16 3 8 8 8 13 0 9 13 7 9
5 0 9 13 3 13
3 13 1 9
12 9 1 12 9 3 15 1 9 0 13 0 9
6 3 16 9 15 13 13
5 13 9 3 11 13
17 3 15 9 9 7 9 13 3 7 15 13 1 9 7 9 13 13
5 3 9 1 9 13
5 3 13 0 9 13
5 15 3 9 13 0
13 9 3 0 0 9 0 13 9 13 7 3 9 13
14 3 3 13 8 15 15 15 13 7 0 9 3 9 13
7 7 3 3 1 15 13 13
35 15 1 9 7 9 13 0 13 15 15 15 9 0 1 15 15 13 13 7 9 15 13 15 13 11 9 15 7 9 3 0 7 9 0 9
16 7 0 9 0 9 15 3 3 3 13 3 13 0 15 3 13
14 9 3 1 15 16 1 0 9 0 7 13 15 0 13
50 7 1 0 9 13 0 9 7 13 0 13 3 9 16 7 15 7 0 9 15 13 13 7 1 15 3 3 13 15 9 13 9 16 16 3 3 13 3 9 7 9 15 7 9 7 9 15 13 13 13
4 16 13 9 13
18 7 3 16 0 13 3 0 13 15 15 1 13 9 15 0 3 13 9
1 13
35 15 15 3 13 3 13 3 9 0 15 1 15 15 15 9 15 13 12 13 15 15 13 15 13 15 1 15 16 13 15 13 15 13 15 13
2 15 13
8 13 9 0 13 13 13 7 9
6 13 3 3 0 9 0
13 0 15 13 1 9 3 13 7 15 13 0 9 0
14 15 3 13 0 16 13 9 0 9 15 13 0 13 13
1 13
17 9 13 11 11 11 7 11 11 7 8 8 8 8 8 9 11 9
4 0 9 9 13
9 11 13 9 3 0 7 15 3 13
24 9 3 0 0 7 0 9 15 13 1 15 13 3 13 13 9 15 15 15 12 16 15 0 13
8 9 9 15 3 13 13 1 15
18 11 9 13 15 15 1 9 7 13 15 1 15 15 1 15 3 13 13
47 15 1 9 16 1 15 3 3 3 3 3 13 16 3 3 15 13 3 3 13 7 3 13 3 1 15 7 1 15 9 0 9 7 9 13 15 13 13 3 3 1 0 9 15 3 3 13
19 0 3 13 13 15 0 9 0 1 11 9 3 7 9 15 3 7 9 13
17 16 13 13 3 7 13 13 1 15 13 7 3 1 0 9 0 13
5 0 9 11 11 13
14 3 13 15 11 7 9 11 11 3 13 13 1 15 9
35 3 1 15 13 3 11 11 15 15 0 8 16 13 15 15 1 15 16 3 1 0 9 13 13 3 3 3 13 13 1 13 7 3 3 13
6 0 1 9 1 9 0
8 13 3 12 0 3 9 9 0
6 3 3 11 13 7 13
2 3 3
7 13 13 1 12 9 9 13
28 15 1 15 3 13 7 13 13 3 16 15 1 0 0 15 9 13 7 16 0 13 0 7 15 1 0 9 13
9 3 11 15 3 15 13 3 3 15
7 13 3 13 9 9 13 9
2 9 13
5 7 16 3 13 13
8 0 0 9 1 15 9 13 13
5 13 13 15 11 15
10 13 13 3 13 9 16 0 15 13 13
4 3 3 13 8
6 3 13 3 0 8 9
29 0 15 16 1 0 9 1 15 0 13 13 8 11 0 13 3 13 13 13 16 3 15 13 8 8 8 8 8 8
11 16 3 15 3 9 3 13 3 15 13 9
15 0 9 13 7 3 3 13 13 16 0 9 15 15 9 13
10 0 7 15 13 0 7 15 3 3 0
13 15 3 15 3 3 13 3 0 9 15 3 13 9
5 3 13 1 9 13
5 1 13 3 13 9
9 3 3 3 3 3 13 7 3 13
6 1 9 3 7 3 13
2 13 15
6 13 9 13 15 15 13
3 15 0 13
3 13 16 13
2 15 13
8 3 13 15 16 1 0 9 13
2 3 11
12 3 3 13 15 13 9 13 9 7 0 0 9
7 3 3 0 9 9 8 13
11 11 15 9 8 8 8 8 8 8 8 8
8 3 13 15 13 16 1 0 13
3 13 16 13
18 13 0 1 0 1 0 1 11 0 9 16 1 15 13 11 13 11 15
7 13 15 15 1 0 9 13
8 15 16 13 3 13 13 15 13
6 11 16 13 13 3 13
4 3 15 13 8
7 1 9 0 0 0 3 13
4 3 13 3 13
16 3 16 0 15 13 3 13 13 13 3 16 15 1 15 13 13
10 15 3 1 9 0 7 1 9 15 13
14 3 3 15 13 16 9 15 13 7 0 9 3 3 9
11 8 8 8 8 8 8 8 8 8 8 8
10 9 15 15 1 9 11 13 9 0 13
17 3 13 6 15 11 1 0 0 9 7 3 3 13 3 13 3 13
12 16 13 13 16 9 0 1 9 13 15 13 9
2 13 11
4 7 13 0 9
15 16 3 13 3 13 13 1 11 13 15 1 15 9 13 11
7 11 9 7 9 7 9 13
8 13 15 3 7 1 0 13 9
4 0 13 9 9
11 3 15 9 7 13 9 3 9 15 13 3
5 9 16 15 13 13
3 15 13 9
8 0 9 0 13 9 3 3 13
7 9 13 9 15 11 13 13
13 13 15 15 0 0 9 0 15 3 3 0 13 0
2 0 13
2 15 15
6 3 11 13 7 13 3
1 13
8 16 7 15 13 0 13 1 15
7 9 15 7 9 13 7 13
3 11 13 13
12 3 9 7 9 0 13 13 15 11 13 15 13
4 7 13 9 9
6 15 3 0 16 13 9
4 11 0 13 15
11 13 15 7 1 0 9 7 3 1 9 13
2 0 13
10 7 3 3 0 3 13 1 15 3 13
2 9 13
28 13 11 11 13 16 15 13 15 1 8 1 15 13 13 15 9 1 0 13 15 7 1 9 7 3 1 9 13
11 3 3 13 15 9 15 13 3 15 9 13
3 16 13 13
8 1 0 9 13 3 16 15 13
5 3 3 9 0 13
28 9 13 1 0 9 16 13 0 13 13 16 11 1 9 1 9 7 3 9 15 13 1 9 3 0 15 13 13
6 15 16 13 9 13 13
9 15 0 13 11 3 9 9 3 9
3 8 8 8
12 3 13 3 7 15 3 3 0 9 7 9 13
64 3 3 3 15 13 13 15 13 15 1 3 3 3 13 9 13 1 9 0 15 13 15 15 0 13 13 3 16 15 15 3 3 13 16 16 1 11 13 13 16 7 1 11 9 13 13 15 15 7 9 13 16 7 15 15 13 13 0 9 1 15 9 13 13
6 3 13 9 13 7 13
28 13 13 3 15 9 1 9 15 1 15 15 13 13 13 13 0 9 16 15 1 12 12 13 13 3 13 3 13
4 15 13 15 0
3 13 3 11
20 16 15 13 7 13 16 1 15 1 11 13 9 15 15 3 0 13 7 3 0
6 3 9 13 13 15 13
13 0 13 15 3 0 9 13 13 15 9 3 13 13
8 0 13 0 7 0 15 15 9
7 3 3 15 13 0 9 13
5 3 1 15 15 13
17 7 3 13 13 9 1 11 16 15 13 13 7 3 3 15 13 0
3 13 3 11
11 15 3 3 15 13 9 16 3 13 1 11
11 15 16 13 15 9 13 13 15 13 15 13
18 3 16 13 9 16 15 13 16 9 13 7 3 13 7 15 1 15 13
3 13 0 0
8 16 3 13 13 15 0 15 13
23 15 3 3 13 15 13 13 3 3 1 9 0 7 9 9 13 13 3 1 9 13 15 13
24 7 16 3 13 16 1 15 9 12 13 7 16 13 15 13 3 3 0 13 13 13 3 13 15
46 16 1 15 13 15 1 11 13 16 13 9 15 7 13 13 13 9 3 7 15 11 13 3 13 13 3 15 1 15 1 15 13 15 0 9 13 13 16 1 9 15 1 15 1 9 13
19 15 3 15 3 13 9 13 3 13 16 15 15 9 7 9 13 1 9 15
7 3 13 15 3 13 15 13
47 13 3 12 9 1 15 13 12 15 15 13 7 13 16 13 0 0 15 11 9 13 15 1 15 9 9 7 13 0 15 13 9 1 9 0 1 15 16 1 11 13 15 13 13 1 9 11
11 13 3 3 15 3 3 7 15 7 15 0
5 3 0 9 3 13
10 16 15 1 15 13 7 3 16 13 13
18 7 16 13 3 3 13 13 1 15 7 3 16 15 15 15 0 9 13
21 7 13 0 3 3 1 0 9 16 16 15 13 9 0 1 15 0 0 13 3 13
12 7 16 1 9 13 3 3 1 15 9 9 9
18 16 15 13 13 15 0 13 16 13 7 15 3 7 13 7 3 13 13
20 15 3 13 13 3 15 15 13 1 9 13 16 3 13 15 7 9 13 7 9
25 15 3 16 3 3 1 0 9 13 1 15 9 13 7 1 15 13 15 7 3 3 1 0 9 13
7 3 0 13 0 1 9 13
18 3 1 11 1 15 13 15 13 3 16 15 13 9 9 15 9 3 13
2 13 3
9 1 9 7 11 9 3 13 3 13
10 9 11 3 7 9 3 13 3 7 9
12 9 9 13 13 3 0 15 15 13 15 3 13
3 13 16 13
15 3 0 0 9 9 9 12 9 13 12 1 9 15 13 3
11 7 16 9 13 0 0 13 3 15 13 13
8 3 16 9 13 15 1 13 13
11 3 9 15 15 15 15 13 13 15 3 13
46 7 13 9 13 16 7 0 9 13 15 15 9 15 13 7 15 9 15 9 15 9 13 3 16 3 13 15 15 9 13 15 9 13 1 9 13 3 16 15 13 7 16 1 15 9 13
10 7 13 16 0 3 3 13 9 9 13
19 15 1 9 13 9 9 13 7 16 13 13 9 9 7 3 9 3 9 13
33 1 9 3 0 15 3 13 13 13 13 3 13 3 13 15 7 3 3 9 15 15 15 13 13 3 9 1 13 7 13 9 15 13
12 16 13 1 9 0 9 9 1 0 9 13 13
38 9 9 13 15 11 1 9 15 9 9 0 0 9 9 13 0 11 15 15 9 13 9 7 13 9 7 9 7 0 9 1 9 3 13 15 15 15 13
12 3 13 9 15 16 1 0 0 16 1 0 0
17 15 16 0 13 3 15 13 13 0 16 13 9 9 15 7 9 15
48 16 9 13 3 16 3 7 9 9 3 7 9 9 15 15 15 13 13 3 0 9 13 13 3 7 9 9 7 9 9 15 13 13 13 13 13 1 9 0 9 9 15 13 15 13 3 13 9
12 3 1 15 0 9 9 13 0 1 9 15 13
8 3 3 15 1 15 9 13 13
4 7 3 13 15
7 3 3 15 9 9 15 13
15 15 9 15 7 9 16 13 1 15 9 13 3 13 15 13
3 0 0 13
3 9 9 13
19 0 15 9 16 15 3 1 9 7 1 9 0 13 13 15 11 11 3 13
2 15 0
11 3 11 1 0 9 1 0 9 1 9 13
8 3 3 1 9 11 1 9 13
8 11 9 3 13 16 15 9 13
13 16 15 1 9 15 3 13 13 13 1 0 11 13
2 3 13
15 13 9 11 0 1 9 15 9 15 9 3 0 13 3 13
11 15 13 13 7 1 9 16 15 13 13 3
1 13
5 1 11 13 3 13
15 7 3 9 13 15 0 1 15 13 3 1 0 15 9 13
3 15 13 13
1 3
21 3 3 15 0 15 1 1 0 9 13 16 0 3 13 15 7 15 16 3 13 13
2 7 13
15 1 11 8 8 8 7 3 0 9 9 15 13 13 15 3
6 9 9 13 0 1 11
11 0 13 11 11 13 11 3 11 0 15 11
13 7 13 1 15 13 1 9 7 3 3 16 9 13
5 1 11 3 15 13
1 15
9 0 1 15 13 3 0 1 0 9
26 0 15 1 1 9 0 3 15 13 3 13 3 13 3 1 0 9 13 11 13 11 13 3 3 3 13
6 15 15 1 11 13 3
13 7 1 0 9 9 13 7 16 15 13 15 13 9
3 13 1 11
10 3 3 15 1 15 13 1 15 13 13
5 13 3 9 16 13
6 3 15 3 13 7 13
4 9 0 9 13
2 13 13
15 3 3 13 9 15 0 7 9 1 9 13 15 3 3 13
13 7 16 13 9 13 13 15 1 15 1 15 9 13
13 13 9 9 9 15 13 13 3 7 3 15 0 3
5 13 11 11 9 3
7 1 11 3 0 13 3 11
7 9 1 9 3 13 13 9
2 11 13
16 15 16 3 13 0 13 3 0 11 13 3 0 9 15 7 9
5 3 13 3 9 13
6 13 3 13 15 3 13
44 16 1 0 15 15 1 9 13 3 13 9 13 15 1 15 15 13 3 15 15 0 13 7 13 13 3 0 15 1 9 0 15 13 9 1 11 9 7 11 7 11 7 11 13
35 3 15 3 0 15 13 13 1 11 15 7 9 7 9 13 0 15 15 13 13 7 0 9 16 3 3 0 13 15 0 9 13 1 11 0
3 7 13 15
6 11 1 11 1 9 13
3 0 9 13
13 0 3 15 16 13 0 15 13 13 13 13 13 9
3 15 3 9
2 9 13
2 3 13
12 7 3 16 0 9 0 0 13 13 15 15 13
2 9 13
2 13 0
4 15 0 0 9
18 3 3 15 13 1 9 15 3 13 13 7 1 9 15 9 0 13 13
13 9 0 9 15 13 11 11 11 9 15 13 15 13
8 3 6 7 1 15 15 3 13
5 13 9 9 0 13
9 15 3 1 9 13 15 3 13 9
5 11 11 11 13 13
6 7 13 1 11 11 9
9 15 3 15 0 15 11 0 9 13
9 13 3 15 13 15 9 1 11 13
7 13 13 0 15 1 0 13
5 1 11 11 13 3
26 15 3 13 0 15 3 0 3 3 15 9 13 1 9 15 16 3 16 15 13 1 9 9 9 3 13
10 3 0 13 15 15 0 13 13 3 9
4 13 15 1 0
12 3 0 0 13 13 9 15 15 9 0 9 13
26 1 15 15 15 13 13 0 7 15 13 13 16 7 13 1 15 7 0 15 3 7 16 15 9 13 13
10 3 13 3 13 16 1 9 0 9 13
22 3 3 3 3 13 13 3 11 13 1 9 13 13 7 9 1 0 15 13 12 9 13
9 1 9 3 0 13 9 7 0 0
4 11 15 9 13
6 7 15 9 9 15 13
9 3 9 9 16 13 13 13 1 15
4 1 11 3 13
12 15 9 13 16 3 15 9 3 0 1 15 13
8 0 3 9 13 15 13 1 9
36 16 11 13 13 0 13 9 0 3 0 13 1 11 13 3 7 3 16 15 0 13 15 13 15 3 1 15 13 16 15 1 7 1 15 13 3
5 13 16 15 13 0
3 7 9 13
4 15 15 13 0
24 15 3 3 15 15 13 13 13 3 13 13 15 13 3 16 0 9 7 0 9 9 0 0 13
9 11 15 0 7 0 9 15 9 13
8 13 13 0 15 13 13 9 15
2 15 3
16 3 15 15 13 13 1 13 16 15 13 3 9 13 3 13 3
12 6 3 3 15 9 13 11 16 1 15 0 13
4 0 15 3 13
4 1 9 13 9
12 7 15 0 3 0 13 8 1 12 9 13 13
12 3 3 13 11 16 1 9 0 11 13 3 13
1 13
6 3 11 0 9 3 0
5 16 0 13 13 9
9 11 13 3 0 7 0 1 9 0
11 15 3 9 11 9 0 15 15 1 13 13
7 3 9 13 0 7 0 9
7 3 0 9 13 7 3 13
4 15 0 9 15
4 13 15 3 13
16 7 13 16 16 15 13 13 0 13 15 1 9 16 9 0 13
4 13 3 15 9
10 11 3 13 3 3 3 1 9 15 13
10 15 13 3 7 9 7 9 7 9 9
10 0 13 11 1 13 15 9 13 13 15
10 15 13 9 16 13 3 0 1 0 9
13 15 3 0 9 9 9 9 3 0 0 9 13 9
4 9 13 9 0
9 7 0 13 15 0 9 13 15 1
33 13 3 9 0 15 13 15 3 13 13 15 9 1 15 15 13 16 3 11 9 3 0 0 9 11 3 6 3 3 15 15 9 13
6 3 15 1 9 3 13
3 15 15 13
5 15 0 9 9 0
12 3 1 11 13 15 11 1 11 1 9 9 13
10 3 15 13 1 9 11 13 9 3 13
4 13 9 7 9
24 15 15 3 13 7 15 0 13 3 15 1 15 13 16 3 0 8 13 13 16 15 13 13 3
5 11 9 15 13 13
7 0 13 3 16 1 11 13
6 15 0 16 13 0 13
21 11 16 15 3 9 13 13 0 7 3 3 15 9 0 13 15 15 1 15 11 13
13 15 1 11 0 13 7 3 13 1 9 13 3 13
7 11 15 13 15 9 0 13
5 15 9 13 3 13
12 0 11 3 16 3 13 3 11 15 13 13 3
7 0 1 15 11 11 9 13
13 15 1 9 3 8 7 3 13 9 15 15 13 13
11 1 3 3 0 0 3 11 13 8 0 0
8 13 3 9 11 11 3 3 11
2 9 13
2 13 9
4 13 3 15 13
2 13 3
6 16 0 13 13 15 11
3 13 1 11
4 11 15 3 13
3 13 15 9
3 0 13 0
8 15 13 3 0 9 9 9 9
9 15 3 1 15 13 1 15 0 9
17 13 3 13 15 15 13 3 16 9 13 3 7 15 1 9 3 13
6 7 11 15 3 15 13
7 15 15 9 13 0 3 13
9 3 3 1 0 13 0 9 13 15
7 0 3 1 15 13 3 9
2 13 13
16 13 3 16 3 15 13 7 3 1 15 13 16 1 9 15 13
20 8 8 8 8 8 3 16 12 9 3 9 15 0 13 15 15 3 3 13 13
33 1 15 9 13 15 1 11 9 13 7 13 15 3 1 11 16 13 0 15 1 15 9 13 0 1 11 13 0 11 15 15 9 13
6 3 15 15 9 0 13
3 13 7 13
4 3 3 15 13
11 13 9 1 15 9 1 15 9 13 15 13
4 0 0 9 13
3 0 9 13
14 1 11 9 15 0 1 0 9 1 15 15 1 15 13
6 3 13 7 13 3 0
1 13
2 15 0
3 3 13 11
20 7 13 9 15 9 3 13 0 13 3 16 1 0 9 15 11 0 0 9 13
12 3 15 13 3 16 13 13 7 16 13 15 13
48 13 0 15 3 13 16 15 1 9 13 3 7 13 11 15 1 15 9 9 3 1 9 0 13 13 7 3 7 15 13 9 13 3 7 0 13 13 7 15 15 3 13 16 16 15 13 3 13
3 13 1 15
9 1 11 13 3 11 13 15 13 13
9 13 3 9 1 9 3 7 13 9
26 1 0 13 13 12 9 9 1 15 12 9 9 15 9 0 15 0 13 7 0 0 15 0 3 3 13
5 3 3 0 11 13
3 11 13 11
6 11 3 13 11 1 11
4 11 3 13 11
7 7 1 9 11 11 13 11
4 11 3 13 11
12 0 3 15 13 6 9 9 1 9 13 15 13
15 13 3 11 1 9 13 3 13 15 9 9 7 13 9 15
3 1 11 11
8 13 3 9 13 13 9 0 3
10 3 13 15 13 13 1 9 1 9 13
12 15 13 13 9 7 9 15 7 13 1 9 11
3 13 9 9
3 9 13 11
6 7 13 9 15 1 9
12 13 3 3 13 1 9 7 6 13 13 15 9
2 13 13
12 7 13 15 15 9 9 7 9 15 7 13 0
15 7 13 9 11 13 7 13 1 11 0 1 9 11 7 11
22 7 13 3 13 15 12 9 11 11 7 11 9 15 1 9 1 11 9 15 13 9 15
6 0 15 13 16 15 13
4 15 13 9 9
17 15 3 13 12 1 9 0 0 7 13 3 9 0 13 1 9 9
8 15 3 13 0 9 13 9 9
14 15 15 13 9 1 13 15 3 13 13 15 1 9 15
5 7 15 13 13 13
7 15 3 13 15 3 13 0
24 13 9 15 13 0 15 13 15 7 13 1 13 7 13 15 16 13 9 9 15 15 1 9 13
11 3 9 3 13 1 9 15 15 1 9 13
9 7 9 15 15 13 1 0 13 15
17 9 15 0 13 15 3 7 13 15 9 15 3 3 15 13 9 15
16 13 13 15 9 1 9 3 9 7 9 13 3 9 13 7 13
6 3 13 9 13 7 9
5 3 13 3 7 13
6 13 3 13 0 1 0
7 7 6 9 13 1 9 15
3 7 13 13
11 13 1 0 9 15 13 1 15 1 9 9
11 3 15 15 13 15 9 9 13 1 9 9
5 13 3 13 1 9
7 7 13 9 13 15 11 13
5 15 13 7 13 15
3 6 13 15
13 7 13 9 15 7 13 15 9 7 13 7 13 15
8 9 3 9 3 13 3 9 13
3 9 13 15
6 15 15 7 15 9 9
3 9 3 13
8 7 6 15 1 9 13 1 15
8 13 9 15 7 13 1 9 15
8 3 1 9 7 9 13 9 15
10 3 13 9 9 13 3 1 0 13 9
5 9 15 3 13 13
8 7 0 13 13 9 1 0 9
8 16 3 13 9 13 1 15 0
4 13 16 15 13
4 3 13 9 15
9 7 3 13 1 9 15 13 9 11
26 13 13 9 3 7 9 3 7 9 1 9 15 3 9 1 9 3 7 12 9 3 7 9 3 7 9
12 3 13 9 11 7 9 1 9 9 3 0 9
9 13 3 9 9 1 9 7 9 9
9 16 9 9 11 13 3 3 9 15
8 15 3 3 9 9 15 13 13
12 15 13 9 7 9 3 3 15 3 13 15 0
22 7 15 9 13 12 1 0 0 9 9 0 3 1 9 9 6 13 15 3 13 9 15
2 0 13
3 9 0 13
10 15 3 0 13 1 9 9 0 13 0
4 13 7 3 13
3 3 13 15
6 7 15 13 9 3 9
10 6 9 15 13 15 3 13 15 13 9
6 7 6 9 9 13 0
10 13 3 9 9 13 1 15 3 15 13
6 7 1 9 15 9 13
9 7 16 11 11 13 1 15 13 13
6 15 9 7 9 13 9
18 13 3 15 16 15 9 0 15 13 13 9 13 9 1 15 1 9 9
6 7 6 0 3 11 3
6 3 13 7 9 0 0
10 1 0 9 13 11 1 9 13 1 9
5 15 3 13 1 9
7 15 3 13 13 15 7 13
5 15 3 13 9 13
13 0 13 13 9 9 9 15 13 0 9 1 9 15
5 13 13 7 13 15
20 16 3 13 0 13 15 9 7 13 9 3 16 9 9 13 7 13 1 9 15
3 15 13 13
17 13 9 9 9 15 7 13 1 9 15 15 9 7 15 15 13 9
14 3 0 13 9 9 9 13 1 9 7 1 15 9 13
2 13 0
4 7 13 1 15
9 7 13 1 9 1 11 9 9 15
7 13 7 7 13 11 1 9
9 13 9 16 13 1 9 13 15 9
6 7 13 15 7 13 13
10 7 13 15 1 9 13 13 13 13 16
3 3 15 13
7 7 16 13 1 9 13 9
8 3 3 13 9 15 16 9 13
7 7 3 13 9 15 7 9
8 7 15 13 1 9 0 13 9
4 13 15 9 0
11 7 6 9 0 1 9 0 13 13 13 15
3 9 13 15
8 7 13 13 9 0 1 0 9
9 7 13 15 0 13 16 13 1 9
6 7 13 15 7 13 13
2 0 13
4 7 13 0 13
11 3 7 12 9 12 12 9 7 3 9 13
2 13 0
9 7 15 13 1 9 13 13 1 9
4 11 9 13 15
7 7 3 13 15 1 9 15
6 9 0 13 15 3 13
4 13 7 13 13
8 3 3 9 9 13 13 1 15
8 3 13 9 1 11 3 7 13
7 7 13 15 7 0 9 13
6 1 9 15 7 1 9
8 1 0 9 13 9 1 11 13
6 3 13 3 16 13 9
3 15 15 13
3 6 13 15
9 3 13 15 3 3 7 3 3 3
3 13 15 13
9 9 0 15 9 13 15 16 13 15
17 1 0 13 9 9 7 9 7 13 9 15 7 13 12 1 9 12
5 7 15 13 13 13
11 3 13 13 15 0 16 9 15 13 7 13
5 15 15 13 1 0
4 15 3 15 13
13 0 13 9 1 9 9 13 3 0 13 1 9 9
4 11 3 13 0
8 3 3 13 1 0 7 0 9
12 13 9 7 13 0 9 13 1 0 3 1 0
6 13 15 15 13 7 13
3 15 13 15
2 13 0
10 7 15 13 1 15 0 13 13 15 9
5 15 13 16 13 15
4 7 3 13 15
9 9 3 15 13 7 15 13 13 13
3 7 13 15
1 3
5 7 13 13 3 9
6 7 15 15 13 0 9
6 15 3 13 11 3 9
1 13
3 13 0 11
10 3 13 15 9 0 0 7 13 0 3
2 13 0
6 1 15 3 13 13 15
3 13 1 9
5 7 13 13 9 13
10 3 13 9 9 13 16 13 15 1 9
5 3 0 13 15 9
12 1 0 9 13 1 15 9 15 13 3 13 9
8 1 9 3 15 13 1 12 9
7 7 13 9 13 1 9 15
9 1 0 12 9 0 9 13 7 9
11 13 1 0 15 16 13 9 15 9 9 15
11 13 3 9 0 7 0 7 13 1 9 9
9 12 3 13 9 15 15 1 9 13
6 6 15 9 0 15 13
16 7 15 13 1 9 13 1 9 9 7 1 15 15 13 1 15
16 6 15 9 7 9 9 16 13 9 9 7 13 9 0 7 13
6 13 0 15 1 9 0
3 13 0 15
7 13 3 13 9 7 9 9
7 7 16 13 9 13 9 0
11 7 16 13 13 9 0 3 13 0 15 9
17 3 3 9 13 1 9 7 13 3 1 9 3 13 3 9 9 9
14 16 3 9 15 0 13 7 9 13 13 16 3 13 9
5 12 13 7 12 13
47 16 3 13 0 9 10 1 9 15 9 13 9 15 13 7 13 13 9 15 13 3 7 13 1 0 13 9 9 0 1 9 15 3 13 7 9 15 13 7 13 15 9 7 15 13 1 9
3 6 9 13
6 3 13 7 0 9 13
13 15 3 12 13 13 13 1 9 7 13 9 9 15
9 13 3 3 15 12 9 13 7 13
9 13 3 3 13 7 13 3 3 13
7 7 0 9 13 1 9 0
5 13 7 13 15 13
12 7 3 15 13 0 7 1 9 7 13 1 15
5 0 7 3 13 15
12 7 13 13 16 13 11 9 0 15 13 9 15
8 13 3 0 13 0 7 13 0
12 3 13 12 1 12 15 13 11 11 1 9 9
2 9 13
4 3 15 13 13
3 13 7 13
4 3 13 0 11
3 13 0 11
10 7 13 3 13 1 9 15 13 7 13
7 7 13 3 7 13 15 13
24 3 15 13 6 11 12 1 12 13 7 1 15 9 0 1 9 7 9 1 9 9 7 0 9
10 3 13 7 9 13 1 11 7 13 15
11 3 1 15 13 13 1 9 7 3 15 13
2 0 13
3 3 13 15
9 3 13 1 9 15 7 9 15 13
13 13 3 0 9 13 15 15 7 13 0 15 13 3
8 7 13 13 11 9 11 15 13
2 15 13
10 7 13 15 1 9 9 3 13 15 9
12 1 9 3 0 13 9 13 9 12 13 15 13
5 13 3 9 13 0
4 15 3 0 13
7 11 3 13 13 15 16 13
11 7 13 1 9 15 13 11 15 13 11 9
7 16 9 9 13 13 1 9
12 15 0 3 3 9 15 13 13 1 15 13 15
3 0 3 13
5 3 9 9 13 0
15 0 3 9 15 13 1 9 13 9 9 7 9 1 11 13
3 13 3 13
5 13 3 9 13 9
3 3 15 13
7 13 9 15 16 13 1 11
4 7 13 15 13
4 9 13 1 9
6 7 13 13 1 9 0
16 16 3 13 13 11 13 11 1 11 13 9 9 9 7 13 16
3 7 13 11
2 0 9
5 13 3 9 11 13
7 7 16 13 15 13 15 16
7 11 3 13 15 13 9 15
28 3 0 13 13 13 7 13 9 3 16 3 3 13 3 1 9 13 7 3 1 0 9 13 7 13 1 15 3
1 13
4 7 3 0 13
14 7 9 7 9 13 16 13 1 9 7 9 13 9 15
4 7 13 0 11
8 7 9 0 1 9 0 13 13
7 3 9 13 9 9 3 9
3 3 0 13
14 0 3 13 3 16 13 1 15 16 0 13 3 13 9
5 7 13 11 9 11
11 7 16 9 1 15 13 3 13 13 9 0
13 7 3 13 13 1 15 13 15 7 13 1 15 9
23 7 13 13 1 15 9 0 3 16 1 9 13 13 1 9 7 15 9 1 9 1 9 13
5 7 15 13 1 9
27 0 3 15 3 13 1 9 15 13 16 13 13 7 3 13 7 13 13 7 3 13 16 13 7 13 15 9
7 7 15 13 15 1 9 13
3 7 13 0
2 7 13
2 13 3
1 13
27 7 13 15 1 9 3 13 15 1 9 9 1 9 0 15 9 13 1 9 7 3 9 3 15 15 13 13
5 13 9 0 1 9
5 7 13 15 3 11
22 16 7 13 9 13 0 13 15 9 13 13 16 13 1 0 7 3 13 15 7 13 0
12 7 13 1 0 7 13 15 9 0 7 13 0
3 15 15 13
2 13 13
6 7 13 9 9 13 0
7 7 13 3 13 1 9 15
5 7 13 15 11 16
19 7 15 3 13 15 3 7 13 15 13 3 13 9 1 9 15 1 9 0
6 9 13 3 12 1 9
12 7 13 15 7 13 15 0 13 7 3 15 13
3 9 11 9
12 7 13 9 1 11 13 0 15 15 13 7 13
17 7 13 13 1 15 16 13 3 9 3 13 9 7 13 13 0 0
3 3 9 13
10 7 13 9 9 12 9 0 7 1 9
9 7 3 13 13 1 15 7 13 0
9 16 7 13 13 1 9 3 13 15
13 3 9 15 3 13 1 9 0 7 0 9 13 9
9 3 0 13 9 9 16 9 15 13
21 15 13 1 9 13 1 15 15 13 15 13 7 15 1 9 13 0 13 15 13 9
9 15 0 0 1 3 13 7 13 9
6 3 0 13 7 13 15
5 7 13 13 9 15
17 1 0 9 3 16 9 0 13 3 7 13 15 13 13 9 13 0
16 7 13 12 9 9 13 13 7 13 9 15 16 13 7 13 9
5 15 9 0 13 9
3 9 3 13
1 12
3 7 13 13
8 7 1 9 13 9 15 13 15
9 7 13 13 15 16 15 13 1 0
12 15 3 13 9 15 1 15 7 9 0 15 13
5 7 13 13 1 11
2 13 0
17 7 13 15 16 7 11 13 7 13 0 15 13 3 13 13 1 15
4 15 13 15 13
2 1 9
7 0 7 0 9 15 15 13
5 7 3 13 13 11
13 3 0 13 16 1 15 1 9 13 15 13 0 0
3 11 3 13
26 0 13 15 0 13 1 9 0 3 12 9 13 13 1 9 9 0 3 9 15 3 13 7 9 3 13
6 7 3 13 3 13 0
13 1 0 13 9 9 15 7 9 7 13 1 9 15
4 9 3 13 13
4 11 3 13 15
11 15 13 13 7 13 0 7 13 9 1 9
10 9 3 0 13 13 1 9 9 9 13
3 13 11 13
12 7 13 15 7 13 15 7 13 15 7 13 15
3 13 15 13
9 13 16 0 15 13 13 9 13 15
6 7 13 0 0 16 13
5 7 13 0 11 13
20 13 1 9 15 13 1 15 7 3 13 3 13 9 13 1 15 15 3 9 13
9 7 13 0 9 15 7 13 1 15
13 7 13 15 16 3 9 13 9 13 1 11 1 12
11 7 16 13 9 13 13 13 7 13 1 9
10 7 16 3 13 13 9 0 13 1 9
23 7 16 13 1 13 13 16 15 13 1 15 16 3 9 15 15 1 9 13 13 15 9 15
11 7 13 15 7 13 15 1 15 9 0 13
1 13
15 7 3 15 13 7 0 13 7 0 15 15 13 15 3 13
5 15 3 13 9 9
14 7 13 1 15 15 1 9 7 9 16 15 13 1 9
3 7 13 0
27 9 11 15 13 16 16 15 9 13 13 7 13 9 7 9 3 13 13 9 15 9 15 7 13 9 9 15
10 1 9 3 16 13 15 1 0 13 9
22 7 13 12 1 9 15 13 0 13 7 13 16 3 0 13 13 15 15 13 0 15 9
6 0 0 15 9 3 13
7 0 3 11 13 1 9 0
12 16 13 3 12 9 0 13 12 9 15 13 9
8 3 13 9 1 9 15 3 13
3 13 3 13
8 3 3 13 15 13 7 9 0
6 13 3 16 9 3 13
12 7 13 9 9 13 7 9 15 13 1 9 13
18 1 9 3 0 7 9 15 13 3 7 9 1 9 3 7 9 3 9
7 13 3 9 7 9 1 9
4 7 13 1 15
6 13 13 9 15 1 9
9 7 13 12 1 9 15 7 13 15
7 7 13 15 7 13 13 11
8 7 13 13 7 13 15 7 13
4 7 13 15 11
4 3 0 3 13
7 0 13 9 15 3 1 9
2 11 13
4 13 3 7 13
5 15 13 13 15 13
11 3 13 1 15 1 9 13 7 3 15 13
9 7 13 1 9 7 13 15 1 9
9 7 13 0 9 1 0 13 11 13
4 15 3 13 9
6 3 15 1 11 9 13
7 0 3 13 13 7 13 16
5 3 0 13 13 0
10 7 16 13 9 13 13 3 3 13 0
4 11 3 13 15
8 7 13 15 7 13 9 13 15
3 7 13 15
3 15 0 13
6 7 15 1 13 13 13
7 13 3 3 9 1 3 13
17 7 16 13 9 11 11 7 11 11 7 11 13 9 16 13 13 15
4 11 13 9 13
2 13 3
3 7 13 15
7 1 0 9 13 7 3 13
9 7 15 9 13 9 13 3 9 9
9 7 0 9 11 13 1 9 9 15
5 7 13 9 13 11
6 7 13 9 1 15 13
16 0 13 0 7 9 0 13 7 13 0 9 9 9 11 9 15
3 13 3 11
9 0 15 1 9 7 0 9 9 15
5 13 9 1 9 15
16 7 13 9 7 0 15 16 13 9 9 15 1 0 7 13 15
4 11 13 9 15
3 7 13 13
8 0 9 0 13 13 9 11 11
23 6 3 13 15 9 0 15 13 15 9 16 13 13 15 3 9 15 13 11 9 1 9 11
10 7 13 11 7 11 7 9 13 1 9
15 7 9 13 1 9 0 3 13 15 9 16 3 13 11 9
9 7 13 11 9 9 11 1 9 11
29 7 16 13 13 9 12 13 0 1 11 1 9 9 0 13 7 9 16 13 13 9 11 1 11 7 3 13 9 15
4 7 13 1 0
20 7 13 1 15 9 11 13 9 9 1 9 9 3 13 13 1 9 9 11 9
9 13 3 9 0 9 7 3 13 13
6 7 15 13 9 3 13
5 7 0 13 9 15
15 13 13 3 16 13 15 9 3 11 13 7 13 13 13 9
4 7 13 0 13
5 7 13 11 13 0
11 7 13 15 9 9 13 1 0 3 1 9
9 7 15 1 9 9 13 13 1 15
11 15 13 13 1 11 13 3 0 1 9 15
7 7 13 7 13 0 1 9
4 13 15 15 13
6 9 3 11 13 0 9
11 7 13 3 13 15 13 16 13 15 13 11
14 13 3 1 12 9 15 13 11 13 15 1 9 13 3
13 7 13 9 15 13 1 15 9 16 13 7 13 15
23 7 13 13 16 13 1 12 9 7 6 9 0 9 7 13 11 7 13 1 9 13 15 13
11 7 13 9 0 16 13 7 13 1 9 15
10 1 9 13 0 1 9 1 0 1 11
12 16 3 13 16 9 9 9 13 1 9 13 9
3 13 0 3
10 3 13 15 0 13 9 7 15 3 13
9 15 9 1 9 0 13 1 9 0
5 15 3 9 13 0
13 13 3 9 7 9 16 1 9 13 16 13 13 0
2 7 13
14 7 15 9 13 15 13 16 9 1 0 13 7 13 15
8 3 6 15 0 16 13 9 15
4 13 1 13 15
8 3 3 9 9 13 16 13 0
8 0 3 9 15 13 13 13 15
17 9 13 3 9 1 9 15 7 3 13 16 13 9 1 9 9 15
17 15 15 13 1 15 7 13 9 15 7 13 15 13 15 15 0 13
4 15 0 13 0
13 1 15 3 15 0 3 13 0 13 16 13 1 15
11 7 13 15 13 13 9 13 9 15 13 0
5 7 13 7 13 9
8 7 13 11 9 15 1 15 0
9 7 0 13 15 3 13 13 1 15
3 3 13 15
11 15 3 0 13 9 9 0 7 15 0 13
10 13 3 0 15 1 9 16 13 1 0
2 9 13
6 7 13 1 9 13 11
4 1 15 13 15
3 13 1 9
6 7 15 13 1 9 0
4 9 13 9 9
17 3 3 13 0 15 3 13 3 7 0 15 3 13 7 1 3 13
12 7 15 13 1 9 7 9 15 7 13 1 0
4 3 13 9 15
3 3 15 13
9 7 13 15 16 13 15 1 0 13
12 7 13 0 9 1 15 9 13 16 1 15 13
23 7 9 15 13 1 9 9 1 9 12 15 1 9 13 15 9 15 3 7 1 15 13 13
3 13 15 15
8 11 3 13 0 9 13 9 9
7 15 3 13 9 15 13 13
17 3 7 9 3 7 9 3 7 9 3 7 9 3 7 12 9 13
7 7 13 9 13 0 15 13
21 3 13 15 0 3 12 9 7 12 9 16 3 15 13 7 13 1 15 0 9 9
9 7 13 13 15 13 0 9 9 12
2 11 9
4 13 3 15 3
10 0 3 0 13 13 13 9 7 13 15
3 9 13 15
6 13 3 15 1 9 9
9 7 15 15 13 13 15 15 15 13
9 7 13 13 1 9 9 16 13 0
7 9 9 13 7 9 9 9
3 13 9 9
3 9 3 0
12 1 0 3 9 13 13 7 13 15 1 0 13
12 13 15 16 11 1 9 0 3 13 3 0 9
8 9 3 9 13 15 1 9 15
7 3 9 3 3 13 1 15
5 1 9 15 13 13
4 13 3 11 13
13 7 13 0 1 9 15 13 1 9 7 9 15 13
11 13 13 3 16 13 7 15 13 1 15 9
9 11 0 9 13 15 3 13 1 15
6 7 3 15 13 1 9
22 3 16 3 13 0 13 3 16 9 15 13 1 9 3 15 13 7 13 0 3 13 0
8 7 9 3 1 9 9 13 0
12 15 9 1 15 0 13 13 7 9 1 9 13
7 7 15 3 13 15 1 13
3 3 0 13
11 3 9 13 1 9 11 7 6 0 11 3
13 9 3 13 1 15 13 13 3 3 13 13 1 9
13 6 15 9 16 13 0 9 1 9 7 9 1 9
5 3 7 9 9 13
13 15 3 0 13 15 3 13 3 7 0 15 3 13
8 7 3 9 9 15 15 13 13
11 9 3 0 13 15 1 15 9 15 13 13
5 7 13 1 15 13
1 13
9 9 0 13 3 9 7 9 3 9
11 3 11 1 15 9 15 13 3 12 1 0
6 13 15 13 7 13 9
4 13 3 15 11
10 15 3 15 0 13 13 0 13 1 15
5 13 3 3 1 9
2 13 15
8 7 16 3 9 13 15 3 13
5 7 16 3 13 9
7 12 9 13 1 15 13 13
11 0 13 9 9 15 13 9 13 1 9 15
14 13 13 1 0 9 16 0 13 15 13 13 7 3 13
6 13 1 15 15 9 9
12 6 13 9 7 9 13 3 7 3 7 0 13
3 13 9 13
3 13 0 9
6 13 3 15 1 9 0
2 13 15
7 3 13 9 9 13 9 15
6 13 3 9 0 1 15
3 0 13 9
9 7 16 13 15 13 1 9 15 13
5 9 15 13 12 9
4 7 15 0 13
4 13 7 15 9
10 7 13 12 1 9 7 13 15 0 13
4 3 15 13 0
5 3 3 3 13 13
3 12 9 9
2 13 0
13 7 16 1 0 0 3 13 15 15 13 15 13 15
9 3 15 9 0 13 9 13 1 9
13 13 13 3 16 13 0 7 13 1 9 1 9 11
27 7 1 0 15 1 15 7 15 9 0 13 13 16 0 15 13 3 13 1 15 3 13 3 7 3 3 13
3 13 3 0
21 7 16 3 1 9 13 1 15 7 3 1 9 13 13 1 15 13 13 15 13 0
20 13 15 13 7 13 15 7 13 15 16 13 7 13 7 1 0 15 13 7 13
4 11 9 13 15
4 7 12 3 13
7 6 3 9 9 1 15 13
14 7 3 13 13 1 9 11 3 13 3 1 9 9 9
16 15 9 3 13 11 1 11 13 9 7 9 1 9 7 15 13
5 12 13 7 0 13
14 13 3 7 9 1 0 16 13 3 13 7 3 13 13
18 9 3 3 13 9 13 15 13 1 15 9 7 9 7 9 13 1 0
5 0 13 15 15 13
5 11 3 13 0 13
5 15 0 3 0 9
5 15 13 11 13 15
4 7 13 15 13
7 13 3 11 12 7 13 0
5 11 9 11 13 15
4 7 11 13 0
9 7 3 13 1 9 16 9 0 13
5 13 11 1 15 16
6 7 13 9 1 0 13
6 9 9 15 13 12 9
15 13 16 15 0 9 13 13 15 3 13 7 13 15 3 13
12 3 9 15 10 15 13 15 13 1 15 13 3
5 13 3 15 13 13
23 7 16 13 3 1 9 9 9 13 15 9 13 13 13 9 9 0 1 15 15 13 9 13
7 3 3 0 13 1 9 15
11 9 3 9 7 9 7 9 9 13 0 13
8 9 11 1 9 13 7 1 9
7 13 3 13 1 9 9 0
4 13 3 9 9
4 15 13 13 0
20 7 13 13 9 15 15 0 13 16 13 15 1 9 7 13 0 9 7 9 9
2 13 13
9 7 0 13 9 7 13 13 1 9
18 0 3 15 0 13 9 0 7 9 1 0 3 7 13 3 7 13 9
4 13 3 1 0
4 0 13 9 0
4 13 3 0 13
8 13 3 0 13 7 3 3 9
7 7 13 9 15 1 9 15
30 7 13 9 1 9 7 9 7 9 7 1 9 13 9 1 9 9 9 7 9 13 9 1 9 7 9 15 13 0 9
4 9 7 9 13
9 7 13 9 9 7 9 3 15 13
3 3 0 13
11 7 16 13 13 9 13 7 12 9 1 15
5 0 13 1 15 9
4 9 9 13 15
27 7 15 13 15 3 13 15 9 15 9 16 13 7 13 1 9 15 1 9 7 13 1 9 13 12 9 11
9 3 13 3 9 16 3 13 13 15
6 7 16 1 0 13 13
5 13 16 13 1 9
3 7 13 0
5 9 3 13 1 9
8 13 3 15 13 1 9 9 9
3 11 3 13
6 16 9 13 3 15 13
3 7 13 0
4 15 3 13 9
8 13 3 11 1 9 9 7 9
5 3 15 15 0 13
13 3 13 15 1 0 7 6 15 0 9 13 13 15
2 13 0
5 11 3 13 9 15
2 7 9
11 7 13 9 13 7 13 0 9 1 15 13
6 13 3 0 13 0 13
6 3 15 1 13 1 9
17 13 3 15 0 15 1 3 7 9 15 13 13 15 1 11 0 13
12 12 3 9 3 9 13 1 9 13 15 13 9
12 7 13 1 9 13 0 15 0 12 7 0 15
7 9 3 0 13 16 15 13
15 7 3 15 13 0 9 7 9 15 1 9 9 7 13 15
16 7 13 1 11 7 15 9 13 0 1 15 9 15 1 15 13
4 7 13 1 3
2 13 13
10 3 0 13 15 9 9 0 7 9 9
13 7 13 13 16 13 0 13 1 15 7 13 1 9
10 7 9 1 9 13 7 9 15 3 13
9 7 9 9 13 13 7 13 1 15
9 0 9 15 13 1 9 9 15 13
2 3 13
5 15 9 13 1 9
11 0 1 11 13 13 1 11 3 13 11 13
10 7 15 13 15 13 1 9 0 15 13
2 15 13
6 13 11 15 13 13 11
6 13 11 11 7 13 15
3 3 15 13
3 7 13 15
4 3 13 9 15
2 7 13
22 7 16 13 3 9 1 9 15 13 1 9 9 3 7 9 7 0 13 9 7 9 13
9 13 9 0 7 1 12 9 13 0
8 0 13 1 15 9 7 13 15
2 13 11
5 13 11 7 13 15
17 3 3 13 9 9 15 1 9 16 13 9 7 16 13 9 1 15
18 13 3 7 11 13 1 11 1 11 16 9 0 13 3 7 13 7 13
5 15 13 9 9 13
9 15 13 15 9 13 16 9 0 13
5 13 3 3 9 11
5 3 3 13 9 9
13 15 3 13 1 9 15 15 13 15 3 13 1 0
3 3 13 16
4 15 13 15 13
3 13 15 11
7 13 1 9 7 13 1 15
11 3 15 13 16 3 12 9 13 7 9 13
11 16 13 3 1 0 9 13 15 16 3 13
7 3 15 3 13 1 9 0
3 13 15 11
7 7 13 0 7 9 15 0
13 9 9 3 13 16 16 13 13 9 13 15 1 9
6 3 13 15 13 9 15
9 3 13 15 11 1 9 7 13 0
4 6 6 13 15
29 6 6 13 15 16 15 9 15 13 7 13 15 15 13 15 13 9 0 7 1 9 3 13 7 13 1 9 1 9
11 16 15 9 13 1 15 9 15 3 13 0
22 9 3 15 13 15 9 16 13 15 0 9 15 15 13 9 13 1 15 16 9 15 13
10 15 13 1 9 9 15 7 3 13 15
14 7 13 15 9 0 16 13 9 15 13 1 0 15 13
10 13 15 12 1 9 15 11 9 11 11
7 3 3 13 13 13 9 15
6 9 3 9 0 13 13
8 7 16 13 15 1 9 13 15
5 13 11 7 13 15
16 3 11 13 15 9 1 9 7 9 15 13 15 9 1 9 0
9 7 15 15 13 1 15 3 13 3
3 1 9 13
4 6 6 13 15
9 3 13 0 15 9 15 13 1 13
19 3 13 15 13 9 7 15 13 1 9 3 15 13 15 3 0 13 1 15
9 16 3 13 9 9 13 3 13 3
6 7 3 3 1 0 13
6 7 1 15 12 9 13
7 16 0 13 13 15 15 9
7 0 16 13 15 13 1 11
9 15 3 3 13 1 0 1 9 9
5 3 11 13 15 9
20 16 9 13 9 1 9 16 3 13 9 11 15 13 16 0 9 0 13 1 9
7 7 15 13 7 3 13 13
3 13 3 11
5 13 15 7 3 13
2 15 13
7 13 3 9 1 9 7 9
15 13 11 1 15 0 15 13 1 15 9 15 12 13 1 15
8 7 13 15 1 0 7 13 15
9 13 3 12 1 12 13 13 1 0
6 13 7 3 3 13 13
7 3 13 3 13 7 3 13
2 13 11
7 3 13 15 3 0 16 13
3 13 3 15
4 3 13 15 0
3 13 15 11
8 7 15 15 13 1 9 15 13
6 15 1 9 3 13 13
6 7 9 9 15 13 13
11 3 3 13 15 16 9 13 15 7 9 13
5 3 13 16 9 13
4 7 3 13 15
4 6 6 13 15
11 15 13 13 9 15 15 13 15 16 9 13
3 15 13 16
7 0 9 15 13 11 9 13
11 13 3 9 3 9 13 11 7 13 9 15
4 13 3 0 3
11 13 16 0 13 9 15 7 16 0 13 13
2 9 13
3 15 13 15
7 15 13 16 11 13 13 9
9 1 9 13 13 0 7 15 13 15
3 3 0 13
4 3 3 13 16
13 0 3 3 13 7 13 1 15 16 3 13 9 0
7 7 13 7 13 7 9 13
7 7 13 15 7 13 15 15
6 0 9 13 1 9 15
8 7 13 11 1 9 1 9 11
19 7 15 9 0 13 15 7 3 13 1 0 7 3 13 15 15 1 9 15
19 1 0 9 3 13 15 7 1 9 7 16 15 9 16 13 13 15 0 9
24 7 13 3 1 11 1 0 9 3 13 11 13 3 7 13 3 7 0 13 1 15 7 13 16
16 9 0 3 13 1 9 7 1 9 9 16 13 9 9 1 15
12 16 15 13 1 9 3 13 16 9 0 9 13
6 3 3 13 15 11 3
9 11 3 3 13 16 11 13 13 0
3 13 15 11
9 0 3 13 13 3 7 13 1 15
2 13 15
2 13 11
7 9 9 13 15 16 13 15
8 13 3 9 7 9 9 7 13
17 0 3 13 9 9 7 13 0 11 1 9 1 9 16 13 15 0
11 3 0 9 3 13 12 9 7 13 13 0
11 7 13 11 9 7 13 1 15 3 13 13
6 6 9 0 1 15 13
11 3 9 9 13 1 9 13 13 15 0 13
4 9 13 15 9
6 3 9 0 9 13 3
6 3 0 9 1 15 13
12 0 13 11 3 13 9 15 7 13 13 1 15
10 3 3 13 16 13 9 7 16 13 9
5 13 3 1 11 11
9 16 3 13 15 3 13 9 15 1
14 16 3 13 9 15 7 13 9 15 16 13 3 13 15
6 3 13 9 0 9 15
7 15 13 16 15 13 15 13
9 3 16 13 0 1 9 11 13 15
25 15 3 13 16 9 13 11 16 13 15 11 13 15 15 9 13 15 1 9 0 7 0 16 15 13
7 9 0 13 15 16 13 3
6 3 3 13 13 15 3
9 16 3 13 15 16 13 13 15 9
8 16 13 15 3 9 15 3 13
11 3 13 16 15 1 9 7 9 1 15 13
6 16 13 15 9 15 13
8 15 3 13 15 13 1 9 15
21 9 3 9 0 15 13 9 1 9 15 0 15 13 15 7 13 15 15 15 13 15
6 3 3 0 13 15 1
7 13 1 15 7 15 1 15
20 16 9 15 13 13 1 9 15 3 3 15 9 15 9 13 7 13 1 15 9
11 16 9 15 13 13 16 15 0 15 9 13
8 3 3 9 3 13 1 9 15
13 7 13 9 16 15 15 13 15 13 9 15 13 9
9 16 3 3 13 9 3 13 1 15
10 0 15 13 16 1 15 13 7 13 15
1 0
16 16 3 13 9 3 3 13 9 1 9 16 13 13 9 1 9
6 0 1 9 13 13 15
4 7 9 15 13
2 7 13
18 7 3 13 15 15 9 1 15 3 0 9 15 13 16 9 13 1 15
9 7 15 15 15 13 7 15 15 13
22 15 13 15 9 15 7 9 9 15 13 16 3 13 1 9 3 3 15 3 13 1 9
25 15 1 15 7 15 1 15 16 13 13 1 12 7 13 9 16 15 15 13 7 13 15 3 15 13
13 11 3 13 15 15 13 13 1 15 13 7 13 15
2 15 13
9 7 13 9 9 7 13 15 9 0
8 13 3 11 11 11 7 15 9
12 13 3 9 7 9 1 9 16 9 13 7 13
11 0 3 16 13 12 13 9 13 9 11 13
4 13 0 7 13
8 13 3 11 1 15 3 7 13
6 13 3 3 1 9 11
2 13 11
8 15 15 13 1 9 13 15 9
4 13 3 11 9
9 13 3 11 13 0 9 7 0 9
3 13 15 9
11 13 16 9 13 13 15 7 9 13 13 15
12 7 13 1 9 1 9 15 13 11 3 3 11
3 13 15 11
4 11 9 9 9
4 13 3 1 3
3 3 13 9
5 7 13 9 13 9
5 9 3 13 1 15
11 7 1 9 9 0 1 15 3 15 13 13
3 3 3 13
3 13 15 0
2 15 13
3 13 15 13
9 7 0 16 13 13 15 9 7 9
15 11 3 12 1 12 15 13 11 3 13 1 15 3 13 11
17 13 9 15 3 7 13 9 15 7 13 9 15 7 13 1 9 15
8 3 13 15 3 11 1 9 11
8 9 3 3 13 13 11 1 9
9 7 3 3 13 0 13 1 9 9
12 13 11 11 7 13 9 1 9 0 0 9 12
6 11 11 13 15 3 0
2 13 15
2 13 15
6 9 15 13 15 13 15
11 0 13 9 15 9 13 1 0 7 13 0
10 15 3 13 9 0 3 1 0 0 9
7 9 0 15 13 13 1 9
12 7 0 3 13 9 1 9 9 7 13 13 0
3 7 13 13
17 13 3 0 9 13 9 7 9 13 13 16 13 15 9 15 0 13
12 13 3 11 1 12 13 9 15 7 13 13 15
15 9 13 1 9 7 9 1 9 16 13 9 9 0 7 0
14 3 3 13 9 15 1 9 3 7 13 0 15 13 9
4 13 9 9 15
10 15 3 9 0 13 13 7 13 15 13
26 3 3 13 3 1 9 7 13 1 9 9 13 9 1 9 7 9 9 13 9 7 13 9 1 15 9
3 11 3 13
11 7 13 13 9 7 9 1 15 15 13 0
12 7 3 9 13 16 1 9 13 3 3 9 15
15 15 13 9 9 7 9 15 13 9 1 9 15 13 1 11
6 7 13 15 1 0 13
7 13 3 15 3 1 9 13
20 3 0 13 13 15 3 13 3 13 15 1 9 16 15 13 9 1 15 15 13
10 7 16 13 13 13 9 1 15 13 13
29 11 3 15 13 13 11 1 9 15 13 13 9 9 9 0 9 1 13 9 13 0 7 13 9 7 13 1 9 9
9 7 13 13 9 0 1 15 15 13
12 6 9 15 15 13 9 15 1 9 7 13 15
31 3 3 13 13 1 9 9 9 7 9 3 16 1 9 13 0 7 13 1 9 7 9 16 13 11 3 9 0 13 15 15
6 7 13 1 9 16 13
7 7 16 13 0 13 1 9
8 0 1 13 13 7 13 13 0
10 3 16 13 1 9 9 0 7 9 13
18 13 3 9 9 1 15 0 9 12 0 9 7 9 15 13 1 0 9
23 13 3 15 1 9 15 13 0 7 0 7 0 7 15 15 13 1 11 7 11 13 1 11
2 15 13
17 13 9 15 9 1 9 0 7 9 15 13 7 3 13 15 9 12
6 7 3 13 9 9 15
9 0 9 13 13 11 7 13 0 9
6 7 13 15 1 9 13
6 11 3 13 13 13 9
25 0 11 15 13 13 15 15 13 9 7 9 0 9 9 7 9 13 1 9 9 15 13 0 1 9
16 7 9 13 1 0 9 7 13 9 9 7 13 1 9 9 15
6 7 3 0 1 0 13
15 7 13 15 15 13 1 9 0 15 15 3 9 7 9 13
6 7 13 11 13 7 13
7 3 15 13 13 13 13 9
11 13 3 15 1 16 0 9 9 15 13 15
16 16 13 3 11 16 1 9 9 9 13 9 0 13 15 9 13
4 13 3 11 13
4 13 3 9 11
13 7 3 9 1 13 15 1 9 3 3 13 9 15
3 7 13 9
8 7 16 9 13 13 16 13 11
15 9 3 0 15 13 1 15 13 13 13 3 9 15 3 13
4 7 9 1 0
18 13 16 9 9 13 15 0 16 13 9 15 1 9 7 9 7 9 11
11 7 3 1 9 13 11 16 0 13 9 9
18 16 3 13 1 11 13 13 15 9 7 15 13 15 3 13 16 13 9
16 13 3 3 9 15 9 11 1 9 12 13 1 9 15 13 9
9 13 13 3 1 9 0 16 13 13
2 11 13
16 13 1 9 3 3 9 0 9 9 9 13 1 15 7 13 15
8 15 16 13 15 13 0 1 11
9 13 9 16 3 13 15 0 7 0
14 13 3 7 13 7 13 1 15 15 13 16 15 13 0
10 11 3 13 0 13 0 15 7 0 9
10 7 15 13 9 15 0 7 0 13 9
5 3 3 13 1 15
12 7 15 9 13 15 15 13 1 9 9 7 11
16 3 9 15 13 13 16 3 13 0 15 9 0 13 3 3 15
6 13 3 3 9 13 15
10 13 3 9 15 16 13 1 0 15 13
3 0 13 13
9 15 16 13 7 13 9 9 13 13
15 9 3 3 15 13 13 0 15 1 9 13 13 1 11 9
18 16 3 13 15 13 11 1 0 9 13 11 13 1 12 9 13 9 12
3 7 13 0
20 3 13 3 16 13 9 9 15 7 13 15 1 9 11 7 1 15 9 9 9
4 11 3 13 13
23 3 0 0 13 1 15 7 13 11 15 13 1 9 13 13 9 3 16 13 9 15 1 0
9 13 3 0 9 7 13 13 9 0
15 13 3 0 11 9 3 3 13 9 15 13 13 9 1 9
7 0 3 13 11 13 11 11
4 7 3 13 9
17 9 9 9 9 11 7 15 1 15 13 9 15 9 9 0 13 13
4 15 3 13 15
15 1 15 15 3 13 1 9 11 13 1 0 15 15 13 13
6 15 13 3 13 9 9
9 3 0 13 9 9 1 15 13 11
16 7 15 9 1 11 0 9 13 0 1 9 9 15 15 3 13
5 3 15 13 9 9
13 7 13 9 13 7 11 13 1 9 13 15 13 13
8 7 15 13 1 11 13 9 16
10 16 3 0 9 13 13 11 13 1 15
12 11 13 3 3 9 13 13 1 9 9 9 15
4 13 1 9 15
7 15 16 13 13 13 1 9
11 11 3 13 11 13 13 13 9 9 1 9
9 7 9 3 13 9 7 13 9 3
12 13 3 1 11 0 9 13 11 7 0 9 11
3 7 13 15
5 7 13 15 9 13
11 3 3 9 13 13 0 3 16 13 9 9
5 7 13 15 3 13
3 13 9 0
6 13 3 9 9 9 0
15 13 3 9 13 7 1 9 9 15 0 7 9 13 13 9
22 0 3 13 0 15 15 13 11 15 13 9 1 15 9 3 13 9 16 0 3 15 13
5 15 13 0 0 13
7 13 3 11 1 0 11 13
5 15 3 3 9 13
7 1 0 13 1 11 13 11
17 7 13 3 13 1 9 15 9 11 11 13 9 15 9 13 13 9
14 16 3 13 0 15 7 9 0 6 9 9 3 15 13
7 15 3 13 9 13 1 9
12 16 3 13 13 11 13 9 13 9 16 13 15
5 1 15 3 13 13
21 16 3 15 13 7 3 13 13 9 1 9 13 1 15 13 9 3 13 1 9 11
25 7 13 9 1 15 1 15 13 9 0 7 13 0 13 1 15 3 16 0 7 13 13 1 9 0
17 13 3 1 11 12 1 13 15 11 7 11 15 13 1 9 1 11
19 7 13 13 9 9 7 9 13 12 9 1 9 13 11 7 11 9 9 11
3 0 11 0
6 7 16 0 13 13 9
9 13 3 9 0 1 9 3 13 13
8 3 3 13 0 1 9 9 13
32 7 3 6 13 15 9 13 1 11 15 1 15 13 13 15 13 3 16 9 0 1 15 9 13 15 13 16 9 7 9 15 13
18 1 15 13 9 13 16 1 9 9 7 9 3 13 1 9 13 15 15
5 7 13 15 1 9
7 7 16 13 3 13 1 9
7 7 13 15 9 7 9 13
7 1 9 3 0 13 13 11
3 15 3 13
3 9 9 13
7 7 13 15 13 7 15 13
2 3 13
28 15 13 9 0 13 11 11 13 3 1 0 9 1 9 11 13 1 9 0 9 9 9 3 3 15 15 13 3
7 15 13 11 9 15 15 13
19 11 3 15 9 1 9 9 13 1 15 13 9 13 1 15 7 13 13 15
3 7 15 13
10 7 16 13 15 9 13 13 15 9 11
1 3
5 13 3 9 11 13
6 13 9 16 9 13 9
4 9 3 15 13
9 9 3 15 9 13 1 15 3 9
2 15 3
7 15 15 13 1 9 9 0
9 3 0 13 9 15 7 0 9 15
6 13 15 15 13 1 11
20 15 3 15 13 7 11 7 11 7 11 7 9 7 9 7 9 7 0 7 0
3 3 3 0
5 3 13 13 1 9
8 3 16 13 15 12 9 3 9
12 16 7 3 15 16 7 0 3 13 7 3 13
6 7 9 15 0 1 15
27 13 3 16 3 1 9 13 3 3 13 15 1 9 16 9 15 13 3 3 15 15 1 9 9 15 11 11
11 7 15 13 15 7 13 9 9 1 9 15
6 16 7 3 9 13 9
28 7 13 0 9 9 7 1 9 7 1 9 13 9 13 16 13 13 1 9 7 13 0 9 15 3 13 9 13
2 13 3
13 15 3 16 15 9 7 1 9 7 1 9 11 13
12 3 0 13 9 9 15 1 15 16 3 0 13
7 3 0 9 1 0 0 13
4 3 3 13 13
8 1 3 0 9 9 13 13 11
7 3 13 9 15 0 3 13
11 16 15 3 9 13 15 3 13 1 9 9
19 15 1 9 13 9 7 13 15 16 0 13 15 1 15 13 3 15 1 9
3 13 15 9
7 15 9 7 9 1 9 9
17 7 13 12 9 11 7 11 7 11 7 11 7 11 7 11 7 11
7 7 13 9 15 1 15 13
14 13 9 15 7 9 7 9 15 7 16 3 13 13 0
13 13 13 15 13 1 9 9 15 13 1 9 9 15
8 15 13 9 13 15 9 13 9
3 3 9 13
5 7 13 1 15 16
18 15 3 13 9 0 15 3 13 9 11 3 13 3 13 1 15 15 9
11 13 9 15 16 9 13 16 13 7 0 13
5 7 9 11 9 13
8 13 15 13 16 15 13 9 15
17 7 16 0 13 7 3 7 0 3 7 0 13 15 13 1 9 15
12 3 7 15 13 7 13 1 9 15 1 9 15
9 7 1 9 9 3 9 0 0 9
7 7 13 9 0 13 9 0
8 7 13 15 9 15 9 7 9
19 7 13 16 13 9 12 1 12 9 7 13 12 1 12 9 13 3 9 9
4 7 6 9 0
5 7 13 9 0 13
10 7 15 9 7 9 1 9 15 13 13
6 1 9 11 12 12 13
5 1 9 11 12 12
1 6
8 7 15 13 1 9 13 1 0
12 7 12 9 15 13 12 9 13 15 16 9 13
14 7 13 7 13 9 12 9 13 1 0 9 13 9 0
8 7 13 13 7 13 9 1 15
5 7 0 9 9 13
20 1 0 12 9 13 13 0 9 9 1 9 7 9 7 9 15 13 1 9 15
9 7 16 13 13 13 12 9 9 15
1 13
12 13 15 3 13 9 7 9 7 9 7 9 0
16 7 9 13 1 9 13 15 1 9 7 13 9 15 9 3 13
8 7 13 9 0 1 9 13 0
5 7 0 9 9 13
11 7 1 9 13 7 13 13 7 13 16 13
12 7 3 13 3 7 9 13 13 15 3 1 9
17 7 13 9 1 9 15 1 9 9 3 9 16 15 13 13 1 9
6 7 9 9 15 13 13
11 7 13 13 0 9 13 1 0 7 13 0
16 7 13 9 0 16 3 9 13 1 9 13 1 9 1 9 9
2 7 13
9 0 13 13 1 9 9 9 7 9
9 15 1 9 9 9 15 13 15 9
13 7 0 9 13 1 9 13 9 0 1 13 1 9
10 7 13 9 11 9 9 7 9 9 13
9 13 7 13 12 9 9 9 1 9
16 7 0 13 9 15 1 9 7 13 13 0 9 13 9 7 9
4 6 13 3 9
10 7 9 0 3 9 13 1 9 1 9
12 7 13 9 0 1 9 0 7 1 9 9 11
2 12 13
7 1 9 15 13 13 0 0
10 7 13 13 0 16 13 15 9 13 0
9 6 9 9 1 9 7 13 1 15
20 3 7 13 1 15 15 13 7 13 9 7 9 3 15 13 13 1 9 9 9
18 9 13 16 13 3 9 1 0 15 13 3 1 0 9 3 13 9 9
85 7 16 15 3 13 9 16 3 9 9 13 15 3 13 16 3 13 0 9 13 7 3 3 1 10 9 9 13 15 13 3 9 13 16 0 9 9 9 13 3 3 3 0 13 16 13 15 15 13 13 1 9 9 3 13 9 13 7 3 3 1 0 9 10 15 13 1 0 13 1 9 1 9 9 15 15 0 9 15 13 13 1 10 9 13
17 3 16 13 9 13 3 3 1 3 0 13 15 16 13 13 3 13
21 1 0 3 9 13 3 9 3 0 16 3 0 9 15 13 9 9 3 3 0 13
26 7 3 3 16 13 7 13 15 9 0 10 7 13 13 1 9 9 3 13 15 13 16 13 15 0 9
17 3 3 9 3 13 0 11 1 3 3 13 1 9 9 15 3 13
23 6 7 13 3 13 9 3 0 7 3 15 13 12 12 16 13 9 10 15 13 13 3 3
10 13 13 3 9 10 1 9 11 1 9
16 3 7 13 9 3 13 9 9 11 0 9 15 11 13 1 9
11 13 3 15 9 3 1 9 11 13 12 9
40 13 3 1 0 3 9 0 9 9 1 0 3 9 1 15 3 13 13 1 9 15 0 13 3 13 1 9 0 0 13 13 9 15 13 1 9 10 15 0 13
70 3 3 15 9 13 9 7 13 3 3 1 9 13 1 9 15 13 3 1 9 15 13 1 0 9 3 3 1 1 9 13 7 13 3 0 3 1 9 13 3 3 1 9 16 3 9 9 9 13 3 3 7 1 12 7 1 12 9 3 3 7 0 3 12 9 1 9 1 9 13
13 15 3 0 9 7 0 9 15 13 13 13 1 11
6 1 3 3 3 11 13
7 3 7 0 3 11 9 13
9 1 11 3 9 12 12 9 13 11
12 3 15 9 13 13 3 7 13 9 7 13 0
8 3 0 9 9 13 13 1 9
24 7 3 3 1 11 9 9 13 1 9 3 1 9 11 13 11 1 0 9 3 13 13 0 11
46 13 3 11 13 9 1 0 15 13 9 7 9 1 11 7 9 0 15 13 9 13 3 3 1 0 9 11 3 9 11 13 3 15 0 11 9 11 11 13 3 13 13 1 9 11 11
9 3 0 13 9 3 13 11 9 11
23 13 15 13 9 9 0 15 13 1 11 15 0 15 1 13 13 1 9 16 3 0 9 13
23 16 3 13 13 1 15 13 9 1 15 9 15 13 13 13 3 13 9 13 0 15 3 13
17 13 3 1 9 9 0 3 13 3 9 3 0 1 0 9 9 11
6 7 3 13 13 1 9
5 3 3 9 3 13
40 3 1 0 9 9 1 3 3 13 7 13 13 15 3 1 3 12 9 15 13 11 15 13 9 11 9 9 15 3 13 11 7 15 11 9 11 15 3 13 11
17 3 1 0 9 13 3 1 9 11 13 1 13 9 0 11 9 9
14 15 3 16 13 9 3 0 13 15 9 13 0 3 0
17 0 15 13 1 0 9 3 0 11 13 0 11 9 9 0 0 13
17 3 0 9 3 0 7 3 0 15 13 1 0 9 1 0 9 13
37 15 3 13 1 9 9 15 13 1 9 0 11 9 3 3 1 0 9 15 3 9 13 1 0 9 0 7 9 3 9 13 13 13 9 15 3 13
28 0 13 9 11 3 13 0 11 11 9 11 9 3 9 13 7 9 9 9 15 9 13 7 1 0 9 9 13
23 7 3 3 15 15 9 3 13 9 16 13 9 3 3 13 13 13 7 13 15 9 13 13
15 3 3 13 13 9 3 13 9 11 3 16 3 0 13 11
34 9 3 3 7 13 0 7 3 0 7 0 9 3 3 0 13 13 9 9 7 16 0 13 15 3 13 13 3 15 13 3 9 0 13
22 3 10 9 15 9 3 3 13 3 3 15 15 1 9 13 15 13 7 3 9 0 0
30 3 3 13 13 9 16 3 13 3 15 9 1 9 13 7 13 9 1 9 13 9 1 9 3 0 15 3 13 9 15
28 3 7 3 3 13 13 7 13 0 9 9 0 9 13 13 7 13 13 1 9 7 3 9 9 13 13 15 9
17 13 3 15 0 9 9 11 7 0 9 15 3 0 7 13 9 0
2 7 0
76 0 3 15 3 0 13 16 3 9 9 3 13 15 13 0 10 11 0 9 0 1 15 9 3 13 3 7 1 15 11 9 15 9 1 11 13 3 3 10 0 15 1 9 13 15 9 13 1 9 10 15 3 3 3 13 3 1 9 0 11 16 9 0 13 3 3 9 13 1 15 13 13 9 10 0 9
3 7 0 13
12 3 3 9 0 3 13 3 1 12 9 1 9
5 0 3 0 9 13
30 3 3 1 9 15 15 13 3 9 1 10 9 15 3 13 7 9 13 1 9 15 15 9 0 9 15 13 7 3 0
29 7 3 13 1 11 13 9 1 9 15 13 1 9 15 11 13 15 13 9 9 11 3 3 11 3 13 11 3 13
29 3 13 3 15 0 15 7 15 15 1 9 9 13 9 15 0 9 9 11 15 15 1 11 13 3 0 9 9 13
45 7 3 3 15 9 13 9 13 11 13 11 9 15 9 16 15 0 7 3 13 13 13 13 0 9 15 13 3 3 3 9 13 7 3 9 13 15 13 13 13 13 7 13 3 11
23 3 9 0 7 0 3 3 9 0 9 9 13 3 1 9 15 1 0 9 7 9 9 13
10 3 3 3 9 0 13 3 3 1 0
2 8 8
11 7 3 1 11 3 1 9 1 9 13 9
6 13 3 0 15 1 9
4 1 0 13 9
7 7 13 9 15 1 9 13
24 3 3 3 9 13 13 9 1 9 15 3 3 13 3 1 9 9 1 9 13 9 3 1 11
20 0 3 9 0 9 3 1 0 9 13 13 9 0 15 3 15 3 13 3 13
2 13 9
7 16 9 13 3 0 0 13
15 1 9 3 0 15 9 1 9 15 13 11 13 3 1 0
10 3 0 1 9 3 1 0 9 3 13
49 0 3 9 0 9 13 3 15 13 16 9 0 1 9 0 13 9 1 11 9 9 9 1 9 3 3 0 9 0 9 13 7 3 3 1 9 13 1 11 7 1 9 15 3 0 9 0 9 13
11 3 3 0 9 3 15 13 3 3 0 9
13 3 3 13 16 16 13 1 11 3 3 9 9 13
3 9 9 0
23 15 3 13 1 0 13 9 3 3 16 0 0 13 7 15 13 15 13 0 9 1 11 13
5 0 13 3 3 9
9 3 16 13 9 13 9 9 7 13
7 3 3 9 0 9 15 13
19 10 0 15 15 13 1 9 0 9 0 15 1 9 13 15 13 1 9 0
10 13 3 3 9 7 9 0 9 7 9
12 7 3 13 9 1 0 9 15 3 9 13 13
10 3 13 3 16 9 3 13 9 1 9
46 3 0 9 13 15 1 0 9 1 9 0 3 0 9 7 0 9 7 16 9 13 13 9 1 9 7 13 13 9 1 9 1 11 3 13 9 1 9 15 13 1 11 7 13 1 9
13 13 0 9 9 1 9 7 13 9 9 3 0 3
3 13 9 13
10 7 15 10 9 13 3 7 13 3 9
17 3 3 1 0 9 15 3 1 12 0 7 0 0 0 0 3 13
27 1 0 3 9 13 1 9 15 13 16 9 13 3 15 0 13 1 11 13 1 9 10 1 15 13 13 9
9 3 3 3 13 13 9 13 13 9
11 15 13 3 13 3 1 9 3 1 9 13
28 3 15 13 3 7 0 3 7 0 15 3 0 9 0 12 9 3 13 3 3 13 13 9 1 15 15 13 13
21 0 3 9 3 13 9 16 13 1 11 16 13 9 13 13 7 9 13 16 13 3
23 0 0 3 3 13 16 9 16 13 13 7 13 3 13 1 9 3 1 9 3 1 11 13
4 0 9 1 11
20 3 0 9 1 9 1 9 9 15 13 1 11 15 9 9 1 9 1 11 13
7 13 9 3 0 9 7 9
3 3 13 9
21 0 3 9 15 13 0 15 9 0 9 13 9 13 15 3 1 9 3 0 1 9
5 3 13 9 15 9
10 3 3 16 13 13 3 13 9 3 0
21 13 3 1 9 13 9 13 9 13 9 7 3 0 7 3 3 1 9 13 1 11
46 7 3 3 0 9 1 0 9 13 16 1 9 0 13 13 1 11 7 3 1 0 9 3 13 13 7 3 15 15 13 13 16 9 0 1 9 15 13 13 1 11 15 1 9 15 13
10 3 1 9 0 13 15 0 13 1 11
7 16 9 13 1 9 15 13
10 13 15 7 16 13 15 3 13 1 9
9 3 3 1 9 15 13 1 0 9
16 16 3 3 13 12 9 13 10 12 9 0 15 3 13 9 0
52 16 3 13 9 9 1 0 12 9 15 13 1 9 3 1 0 3 9 13 13 1 9 3 13 1 9 1 11 3 13 9 13 0 7 13 9 13 1 9 0 15 13 1 9 11 7 13 15 15 13 1 9
46 0 3 3 1 15 3 0 13 7 3 0 16 3 3 9 3 9 7 9 3 7 3 3 3 9 15 13 9 0 9 13 16 7 9 15 13 7 9 1 15 13 0 7 13 13 3
20 9 3 3 0 13 0 9 11 3 12 7 12 13 7 1 0 13 0 9 15
