274 17
42 10 9 1 10 9 16 10 9 13 2 13 16 10 9 0 4 13 10 9 0 13 1 9 0 2 13 1 9 10 9 0 2 13 10 9 0 13 1 10 9 0 2
17 1 13 3 3 2 1 11 11 2 13 9 10 9 1 10 9 2
36 11 12 13 10 9 11 12 13 9 1 10 9 7 10 9 3 1 13 10 0 9 1 9 13 1 11 11 2 9 1 9 0 7 8 8 2
20 13 10 9 0 1 10 9 0 2 9 16 13 15 9 1 10 0 12 9 2
15 9 0 1 9 1 11 1 10 12 2 2 15 13 9 2
32 13 3 3 13 15 16 10 9 1 11 13 1 11 11 2 3 13 1 11 16 4 13 9 1 10 9 1 9 1 10 9 2
48 1 13 1 11 7 11 2 10 12 9 4 7 13 10 9 1 10 9 7 13 10 9 1 9 7 10 9 0 1 10 9 1 13 10 9 1 10 9 1 10 9 1 10 9 1 10 9 2
26 4 1 13 3 1 13 9 7 1 13 15 2 7 4 1 13 16 13 9 0 1 9 1 9 0 2
20 1 11 15 13 9 1 15 9 1 11 1 10 11 2 9 1 0 9 0 2
21 11 11 2 9 1 10 9 13 15 9 1 10 9 0 2 2 3 13 15 0 2
34 10 9 1 11 11 13 13 16 10 9 0 4 13 10 9 1 9 1 10 9 16 15 4 13 1 10 9 1 13 7 13 10 9 2
67 9 1 10 0 9 0 1 11 1 11 2 3 7 10 9 1 10 0 9 2 13 10 9 1 10 9 2 8 2 11 11 2 1 10 9 9 0 8 11 11 9 1 11 1 10 9 16 13 2 7 16 13 10 9 1 13 10 9 1 9 1 10 15 1 10 9 2
32 10 9 0 13 1 10 9 1 10 9 1 10 9 10 11 2 3 7 10 9 0 13 15 9 1 10 9 1 10 9 11 2
16 15 13 10 9 1 10 16 15 13 10 9 12 1 10 11 2
25 1 10 9 13 10 9 16 13 1 10 11 11 7 16 4 13 1 9 7 1 9 1 10 9 2
21 3 13 10 9 0 16 13 9 3 1 10 9 16 15 13 1 10 11 11 11 2
47 15 15 13 16 3 15 13 3 7 15 13 2 16 13 13 15 13 2 2 13 1 0 9 10 9 2 13 1 10 9 1 10 9 1 10 9 1 9 1 10 9 1 9 1 10 11 2
46 3 13 1 10 11 11 1 13 0 2 7 3 3 2 10 11 11 3 15 13 10 9 1 10 9 2 9 1 0 9 16 4 13 10 9 3 1 10 9 1 10 0 9 1 11 2
21 2 3 4 13 10 9 1 9 2 9 2 9 2 9 2 8 2 1 11 11 2
120 3 2 13 1 9 16 1 1 1 10 9 3 13 2 15 13 1 10 9 0 2 7 13 1 10 9 1 10 9 2 2 13 12 9 1 9 2 12 9 0 2 15 1 10 9 7 15 1 10 9 2 7 1 10 9 15 15 13 1 10 9 1 10 9 2 10 9 3 4 13 3 15 1 10 9 0 2 13 12 9 15 13 10 9 2 7 3 15 13 10 0 9 0 2 2 10 9 3 0 2 1 9 3 0 2 1 9 7 9 16 15 13 1 10 9 1 9 0 2 2
10 9 13 1 9 0 7 1 9 0 2
16 11 11 7 11 11 13 10 3 0 1 3 1 9 15 13 2
37 2 10 10 9 16 13 3 1 10 9 13 10 0 9 1 10 9 13 15 1 9 7 9 0 1 15 2 2 13 11 11 2 9 1 11 11 2
32 10 9 13 2 10 9 1 10 9 1 10 9 0 11 2 13 13 10 9 1 9 7 13 15 1 10 9 0 1 10 9 2
52 10 9 1 11 3 13 0 2 3 7 4 13 16 15 4 4 13 3 1 9 2 9 16 15 4 13 13 10 9 7 13 16 3 11 13 13 15 12 9 1 10 11 16 15 13 0 13 10 9 1 9 2
56 15 4 13 15 1 10 0 9 1 10 9 7 16 13 1 10 9 10 15 13 0 9 7 10 9 1 9 3 15 13 2 15 13 7 3 15 13 1 10 7 11 4 13 1 10 9 2 10 1 10 0 9 1 10 9 2
15 15 13 16 15 13 15 1 10 9 16 4 13 11 11 2
14 1 15 2 15 15 13 1 10 9 0 1 10 15 2
54 10 9 1 11 13 16 3 4 13 9 1 15 3 7 12 9 1 10 9 1 11 12 2 1 15 15 1 10 9 15 13 1 13 16 11 4 13 1 9 2 1 9 1 10 9 16 13 10 9 1 10 9 0 2
28 10 9 4 13 1 15 1 11 2 7 3 15 15 13 3 16 11 13 0 1 10 9 1 15 4 13 11 2
22 10 9 3 4 13 10 9 1 9 1 10 9 2 13 1 10 9 7 1 0 9 2
8 13 3 9 1 10 9 5 5
27 16 10 9 0 3 13 3 0 2 15 13 13 1 10 9 0 1 10 9 16 13 10 12 9 1 9 2
20 15 13 16 13 10 9 0 4 13 1 10 0 9 16 15 13 10 0 11 2
36 13 1 11 11 2 10 9 7 9 8 4 13 1 11 11 11 7 11 11 1 10 9 1 10 0 9 2 11 11 11 2 2 3 1 11 2
17 10 4 13 15 1 10 9 1 10 9 2 1 12 9 1 3 2
27 10 11 13 1 11 13 16 13 7 13 1 1 10 1 11 1 12 2 12 13 10 12 9 1 9 3 2
11 2 4 10 0 9 13 10 9 1 0 2
19 10 9 2 1 10 9 2 13 10 16 4 13 10 9 7 13 10 9 2
21 2 16 4 7 13 10 11 11 2 13 1 10 11 2 1 10 3 15 15 13 2
8 2 1 15 4 13 0 9 2
9 15 15 4 13 3 13 10 9 2
24 15 9 13 16 10 9 1 9 3 4 13 1 9 7 10 9 1 9 1 9 13 3 0 2
60 11 11 3 13 10 9 0 1 9 0 2 16 13 10 9 1 11 3 13 10 9 1 10 9 7 10 9 0 13 10 9 15 3 4 13 1 10 0 9 1 11 11 3 7 10 0 9 7 9 3 13 7 9 7 0 1 13 10 9 2
32 10 12 12 1 9 1 11 11 13 1 13 1 10 9 1 10 11 7 10 0 9 1 10 9 1 10 9 2 11 11 2 2
12 7 11 3 4 13 15 1 13 10 9 0 2
32 3 3 2 13 10 9 1 10 9 7 9 1 9 0 3 7 3 1 11 11 2 13 0 1 15 15 13 1 10 10 9 2
20 13 15 1 10 0 9 2 1 15 15 13 1 10 9 16 13 1 10 9 2
31 1 11 1 12 2 9 0 1 10 11 13 1 10 9 1 10 9 1 13 1 10 9 0 7 13 10 9 1 9 0 2
7 2 13 13 3 10 9 2
42 1 10 9 1 9 7 1 9 2 10 9 4 13 15 1 10 9 11 7 11 2 3 13 9 0 2 9 0 2 9 1 9 2 9 1 9 7 10 9 1 9 2
23 2 3 4 13 10 9 1 10 9 9 16 7 3 4 13 15 9 16 13 1 10 9 2
9 7 15 13 10 9 1 0 9 2
25 11 13 2 1 10 9 2 10 9 1 9 16 13 1 9 1 11 11 11 2 13 1 11 9 2
30 10 11 11 4 13 1 15 1 10 0 9 2 1 15 1 10 11 7 1 0 4 13 1 10 0 9 2 11 11 2
29 11 13 1 10 11 1 10 3 12 9 1 13 2 10 9 0 13 1 10 11 0 2 7 3 15 13 1 11 2
70 10 9 4 13 15 2 4 13 1 9 10 9 16 13 1 10 9 10 11 11 2 1 10 9 2 13 1 10 9 1 12 2 13 1 10 0 9 1 9 1 9 1 10 9 0 2 1 10 9 1 10 9 1 10 0 9 0 2 0 2 1 9 0 2 1 0 8 8 8 2
24 13 1 11 10 9 1 11 12 7 1 10 0 9 3 13 10 0 9 7 9 1 10 9 2
38 13 15 0 2 13 15 2 3 15 4 1 13 15 2 1 15 3 13 10 9 2 13 15 2 13 15 1 15 2 13 10 9 2 3 13 15 2 2
36 4 7 11 13 10 3 3 1 10 9 1 13 15 1 9 0 2 7 15 3 4 13 9 1 16 13 10 9 1 11 1 11 3 1 9 2
13 10 9 0 13 9 0 1 10 9 1 10 9 2
30 10 0 11 2 0 7 0 9 2 15 13 10 9 13 15 1 10 2 11 7 0 9 2 2 3 10 9 0 9 2
18 10 9 0 13 10 9 1 11 1 10 11 11 16 13 1 11 11 2
28 13 1 10 9 11 2 11 2 2 11 2 9 1 9 12 9 2 9 1 9 11 7 13 9 1 9 11 2
13 15 3 15 13 1 15 2 13 10 2 9 2 2
17 10 10 9 7 9 0 16 13 1 10 9 1 10 9 13 0 2
28 10 9 1 10 12 9 13 13 10 9 0 1 10 0 9 1 10 9 7 3 13 9 1 13 15 1 3 2
12 1 11 11 13 1 9 1 9 1 12 9 2
42 2 13 13 10 9 1 10 9 16 13 10 9 1 10 11 11 2 13 1 10 9 9 1 10 9 0 1 10 9 1 10 9 1 9 9 1 15 1 10 9 0 2
26 10 0 9 3 4 1 13 15 1 11 11 12 2 10 9 16 13 0 13 1 10 9 1 11 11 2
13 10 9 1 10 9 1 9 7 9 4 13 9 2
19 10 9 2 10 9 2 9 7 13 10 9 1 2 9 2 1 10 15 2
27 3 13 1 10 0 9 2 7 10 9 1 11 4 13 10 9 1 10 9 9 1 16 3 13 11 11 2
50 10 11 11 13 10 9 16 13 13 1 9 0 1 12 9 7 9 1 9 1 9 0 16 15 13 13 1 10 9 0 11 11 11 11 1 11 2 9 11 2 1 10 9 1 13 9 1 10 9 2
25 10 9 13 3 9 1 10 9 2 7 10 9 0 3 4 13 1 10 9 13 1 10 9 0 2
11 4 13 2 11 10 9 2 2 1 11 2
39 1 15 2 3 13 10 0 9 1 10 9 1 10 0 9 1 10 9 2 4 7 13 16 10 0 9 16 15 4 13 1 2 9 3 13 13 12 9 2
32 13 16 10 9 1 10 9 13 1 11 2 10 9 4 13 9 0 1 10 10 9 1 9 1 10 9 1 9 0 7 0 2
14 10 9 1 10 9 13 2 13 10 9 1 10 9 2
43 10 9 11 7 9 1 10 0 9 0 2 13 1 10 9 1 10 9 0 2 13 10 9 3 13 1 10 9 1 10 9 1 10 9 1 10 9 2 1 10 9 2 2
14 2 1 9 13 9 1 10 9 1 10 11 1 11 2
16 10 12 13 9 2 4 13 9 7 15 1 15 13 10 9 2
48 3 3 10 9 13 10 12 12 9 1 9 2 3 1 4 13 1 12 9 3 1 12 12 9 1 9 16 15 4 13 3 13 2 16 3 13 10 0 9 16 13 10 9 0 1 10 9 2
47 10 9 1 10 9 1 9 1 10 9 1 10 9 1 11 2 11 2 9 1 11 2 13 2 1 9 0 2 1 10 9 0 7 0 1 10 9 1 9 7 10 9 0 1 10 9 2
9 10 9 13 3 10 9 1 11 2
28 10 9 13 9 0 7 0 16 13 10 9 1 13 15 2 7 13 9 2 10 9 4 3 13 16 15 13 2
47 2 16 1 10 9 15 13 10 9 16 13 10 9 2 4 13 2 2 13 10 9 2 7 13 16 1 10 9 16 13 9 15 15 13 10 0 9 1 13 1 10 9 10 9 4 13 2
31 7 10 9 1 10 9 0 2 1 10 11 11 7 1 10 9 1 9 1 10 11 10 10 9 4 13 1 10 9 0 2
20 3 9 1 9 13 1 15 3 0 1 10 9 2 9 2 9 7 3 9 2
8 10 9 13 0 1 11 11 2
55 16 15 13 1 9 10 9 13 1 10 0 9 16 13 1 10 9 1 10 9 1 10 12 2 9 1 9 7 9 1 9 1 10 9 0 4 1 13 1 10 9 2 1 10 9 2 1 13 15 0 1 10 9 13 2
19 2 1 15 13 1 9 2 1 10 9 1 11 8 10 9 1 10 9 2
21 1 10 9 1 15 16 13 1 10 9 2 10 9 3 13 1 9 1 10 9 2
62 11 11 3 13 13 1 10 9 11 7 10 12 9 16 4 13 10 9 13 10 11 11 7 3 10 11 11 16 13 15 0 13 3 7 13 16 13 13 12 9 3 1 10 11 11 7 1 0 1 11 3 13 9 1 10 9 3 10 7 10 9 2
71 10 9 1 9 0 16 15 13 16 15 15 13 10 9 2 13 16 4 7 13 10 9 7 16 2 13 0 1 15 16 13 2 2 16 15 13 1 3 10 0 9 7 1 3 9 7 13 1 15 1 10 0 9 2 1 9 0 2 2 10 9 1 9 1 10 9 8 2 0 2 2
62 16 10 9 1 9 13 15 13 1 13 9 1 10 9 2 13 3 1 10 9 11 2 11 2 8 13 9 0 1 10 9 2 10 9 1 0 9 4 1 13 15 9 16 13 13 2 13 2 13 10 9 16 13 13 1 10 9 10 9 1 9 2
30 10 11 4 13 3 16 10 9 3 13 13 15 1 11 13 7 3 13 9 1 13 1 10 9 0 3 10 9 0 2
18 11 11 13 12 9 1 12 9 1 12 9 1 11 2 11 7 11 2
47 2 13 10 9 0 2 7 15 13 0 1 13 15 1 10 10 9 16 3 15 13 1 10 9 1 11 2 2 13 2 3 1 13 16 4 13 10 0 9 7 10 9 0 3 4 13 2
36 10 9 15 13 1 10 9 1 16 9 0 13 1 9 1 9 1 12 9 1 10 0 9 1 9 1 10 9 1 9 13 1 11 11 11 2
46 10 9 2 10 9 3 4 13 2 4 13 1 10 9 0 1 10 9 1 10 9 2 3 4 13 1 10 9 13 1 10 16 2 1 10 9 2 13 10 9 1 9 1 12 9 2
103 3 2 10 9 13 16 10 9 1 10 9 1 9 7 10 9 1 10 9 1 11 2 16 13 1 9 10 9 11 12 2 13 10 9 0 2 1 15 2 15 1 10 9 1 10 9 16 4 13 1 13 1 10 9 1 10 9 0 2 1 10 9 0 2 16 3 13 3 7 10 9 1 10 9 16 15 13 1 12 2 1 10 9 1 12 9 1 9 1 10 9 1 10 2 11 2 2 9 1 9 0 2 2
86 1 9 1 10 9 1 10 9 1 10 9 0 2 15 15 13 16 10 9 2 9 1 9 1 10 9 11 7 0 2 2 13 3 1 10 9 7 1 10 9 0 2 10 9 1 10 9 1 9 0 1 9 1 10 9 2 13 7 10 9 1 9 1 9 0 7 10 0 9 1 10 9 1 9 13 16 10 9 3 4 4 13 10 9 2 2
52 11 11 13 16 4 13 0 9 13 1 10 9 1 10 9 11 11 2 1 11 11 2 11 11 2 1 11 2 11 11 2 11 2 1 11 11 2 11 1 10 11 2 11 11 2 1 11 2 11 7 11 2
27 2 13 10 9 0 1 10 9 0 3 1 10 9 1 10 11 2 2 4 13 11 1 10 9 1 9 2
28 13 10 9 1 9 0 1 10 0 9 1 10 9 2 1 13 16 2 3 0 9 4 13 1 11 2 3 2
91 1 13 1 10 9 1 9 1 10 0 9 1 10 11 1 11 2 13 1 10 9 11 11 11 2 11 11 2 13 16 2 1 15 15 13 10 9 7 10 9 16 13 10 9 1 10 9 2 13 7 3 1 15 2 15 2 13 10 9 1 10 9 2 3 3 1 10 9 2 13 1 10 9 0 1 10 9 2 1 10 0 9 1 9 7 1 10 9 0 2 2
10 3 13 16 13 2 7 16 3 2 2
27 3 13 9 16 10 9 1 10 9 0 0 7 10 9 1 10 9 0 2 13 10 0 9 1 10 9 2
25 10 0 9 13 16 10 9 1 10 9 13 1 9 7 16 15 13 10 10 9 3 1 10 12 2
24 16 15 13 16 15 4 13 9 7 3 15 13 10 9 1 10 9 2 4 13 1 10 9 2
63 9 1 10 9 1 10 9 1 9 9 2 9 2 9 7 9 7 1 10 9 1 11 2 15 13 10 9 0 1 10 9 2 16 1 10 9 13 0 13 10 12 5 1 10 9 1 9 0 2 1 7 3 10 12 9 13 1 10 9 13 15 0 2
15 1 10 9 0 13 10 2 10 9 2 1 9 1 9 2
45 10 9 0 1 11 11 12 13 1 10 9 1 10 9 3 0 16 10 0 9 1 10 9 1 10 9 13 1 10 9 2 1 10 9 7 10 9 1 10 0 9 1 10 9 2
28 15 15 13 2 7 1 3 11 7 11 13 10 9 0 1 9 0 2 1 10 9 2 9 16 3 13 9 2
34 10 9 4 13 1 16 10 9 13 1 9 1 10 0 9 2 16 10 9 13 1 9 1 9 1 10 9 1 11 1 10 9 12 2
58 9 1 10 9 1 9 0 13 1 10 9 1 12 7 12 4 4 13 1 12 7 11 13 16 2 1 15 2 15 4 1 13 10 9 1 13 10 9 10 9 1 10 12 5 1 12 7 3 13 0 13 10 9 7 13 10 9 2
19 11 11 13 1 9 0 1 10 9 0 1 11 1 9 1 10 9 12 2
33 11 11 2 9 1 10 9 0 2 13 1 10 9 1 9 16 2 1 10 9 2 10 9 15 13 1 10 9 1 9 0 0 2
29 10 9 15 13 1 10 9 12 1 10 9 1 11 2 12 8 2 12 2 12 1 9 2 7 11 2 12 2 2
37 2 10 11 2 13 1 11 11 2 11 11 7 11 11 4 13 3 1 10 0 9 11 1 11 13 9 1 10 9 1 10 9 1 10 0 9 2
38 11 11 2 11 11 13 10 0 9 16 4 13 10 12 9 2 16 1 9 1 13 1 12 9 7 3 12 3 7 10 9 3 13 10 9 1 9 2
31 10 12 0 9 0 1 9 1 10 9 0 13 0 1 10 9 1 10 0 11 11 7 1 10 9 1 9 1 10 9 2
11 7 10 9 13 2 3 1 10 9 0 2
44 10 9 15 4 13 1 9 0 16 10 9 4 13 10 9 1 16 4 13 1 10 9 1 10 9 1 11 1 13 15 1 10 9 1 10 9 2 3 10 10 9 13 9 2
103 10 9 0 1 10 11 1 11 2 11 11 2 4 13 1 10 9 0 1 10 11 2 11 11 2 16 2 15 16 4 7 13 13 3 13 3 1 10 9 7 10 9 1 9 0 1 15 16 4 13 1 9 0 2 2 1 10 9 7 4 13 16 2 15 9 16 4 13 1 10 9 13 13 9 1 10 9 7 9 1 9 1 10 9 16 3 13 9 1 10 9 1 9 7 10 0 9 1 13 10 9 2 2
18 10 0 9 1 9 1 15 13 10 9 2 13 15 7 13 10 9 2
40 10 0 9 1 9 1 10 9 13 13 15 1 9 1 10 9 1 10 11 2 1 9 10 9 0 1 10 9 1 11 13 1 3 12 9 7 12 10 9 2
18 10 0 9 1 10 9 1 9 3 13 10 9 1 10 9 1 8 2
34 10 9 13 10 9 1 9 1 9 16 3 4 13 1 10 9 11 11 1 11 11 2 7 10 1 11 2 1 12 9 1 10 9 2
27 1 10 9 2 10 9 1 10 9 13 9 1 13 10 9 1 10 9 1 10 9 1 10 9 1 9 2
39 13 16 1 12 9 1 9 0 13 1 15 7 10 15 1 10 9 16 13 2 10 9 1 9 0 2 10 9 2 0 2 2 0 7 9 1 9 0 2
20 16 15 13 1 10 9 0 2 10 0 9 13 1 12 9 1 10 12 0 2
18 3 3 2 4 7 13 16 15 13 1 10 9 0 13 1 9 0 2
22 10 9 16 13 13 13 10 9 4 8 10 9 1 9 1 11 13 1 10 9 0 2
25 10 9 0 1 10 11 13 10 9 1 10 9 1 11 1 10 9 16 13 10 11 12 1 11 2
24 13 3 1 10 9 0 1 10 9 2 12 2 2 10 9 4 13 1 10 9 1 10 9 2
60 1 10 12 1 10 9 1 10 11 4 13 10 9 1 9 0 1 10 9 1 11 2 13 1 10 9 11 11 1 10 9 2 11 11 11 2 2 13 9 0 1 10 9 0 1 10 9 0 7 9 10 9 1 10 9 0 1 10 9 2
15 2 15 15 13 12 7 12 9 1 10 9 2 2 13 2
50 13 9 1 10 9 1 9 1 10 9 0 12 7 12 2 13 1 3 1 10 9 0 7 15 4 13 10 11 12 1 15 15 3 13 3 13 10 9 1 10 9 2 10 15 13 1 13 15 0 2
18 10 9 0 13 10 9 0 16 13 1 9 0 10 9 7 9 0 2
47 10 9 1 10 9 1 10 9 11 2 11 11 2 13 16 10 9 16 13 3 11 11 13 1 10 9 0 2 16 10 9 3 13 3 0 1 10 16 13 1 10 9 1 12 7 12 2
31 15 13 3 10 9 1 10 9 2 1 9 1 9 13 1 13 4 13 1 10 9 7 10 9 2 13 9 1 10 11 2
67 13 0 13 9 2 10 9 0 7 3 0 1 9 3 0 1 13 1 9 2 1 13 1 9 10 12 5 1 10 9 0 2 13 10 9 0 3 1 12 9 0 2 7 10 9 1 10 9 0 16 2 13 1 10 9 2 4 13 10 9 1 9 1 9 7 9 2
32 15 1 10 9 1 12 9 1 9 15 13 1 10 0 9 1 9 1 11 7 3 15 13 12 1 10 9 16 13 10 9 2
26 11 11 2 16 13 10 11 11 11 1 12 13 16 10 9 0 13 1 13 1 9 1 10 9 0 2
53 1 9 1 10 9 1 9 0 1 10 9 2 11 11 7 11 2 1 12 3 15 4 13 10 9 0 1 10 9 1 10 11 2 16 15 13 10 9 1 10 9 2 7 13 10 0 9 0 15 16 15 13 2
7 7 3 3 15 4 13 2
66 1 10 9 1 10 11 3 15 4 4 13 10 9 16 10 9 2 16 15 13 1 10 9 1 9 2 13 1 10 8 8 2 8 2 7 1 10 9 16 13 10 9 2 1 0 9 7 10 9 1 9 16 3 15 13 1 10 9 1 9 1 10 9 11 2 2
62 1 9 3 13 11 11 2 11 2 2 11 11 2 10 11 2 2 11 11 2 11 2 2 11 11 11 11 2 11 2 2 11 11 2 11 11 2 2 11 11 2 11 2 2 11 11 2 11 2 2 11 11 2 11 2 7 11 11 2 11 2 2
43 10 9 1 10 11 11 2 11 11 2 4 13 10 11 10 9 1 10 9 16 13 10 9 1 9 1 10 0 9 2 10 11 16 13 1 9 1 2 9 2 7 0 2
47 1 12 10 9 11 11 11 2 12 2 2 11 11 11 2 12 2 7 11 11 11 2 12 2 1 13 1 9 0 1 9 0 2 13 10 9 1 9 0 1 13 1 9 0 10 9 2
66 1 10 9 2 13 13 10 9 1 11 11 2 9 1 10 9 0 2 15 3 13 1 13 1 10 11 1 13 10 9 0 16 13 13 1 9 0 7 13 10 9 13 16 15 13 1 10 11 1 9 1 10 12 9 0 2 2 13 11 2 9 1 10 9 0 2
42 10 11 4 13 16 1 10 9 1 10 9 1 11 11 1 11 4 13 9 0 2 7 13 1 16 10 9 16 13 1 10 9 13 16 1 10 9 3 3 13 9 2
33 10 9 11 11 11 1 10 11 13 10 9 16 13 1 10 12 1 10 9 1 10 9 0 7 13 1 10 9 1 11 11 11 2
42 11 13 1 10 9 2 1 10 9 0 1 9 1 10 9 2 16 10 9 13 2 0 2 2 1 15 1 10 9 1 11 2 3 7 10 10 9 13 2 0 2 2
29 1 0 9 1 9 2 9 7 9 1 10 9 0 4 13 3 1 10 9 1 9 1 13 10 9 7 0 9 2
15 10 9 2 1 10 16 11 13 3 2 3 13 10 9 2
33 3 13 3 13 10 9 2 16 10 9 1 11 11 2 9 1 10 9 1 2 11 2 7 11 11 2 1 10 9 13 9 0 2
38 1 11 2 9 1 11 7 11 3 13 10 9 0 2 1 10 15 10 9 13 1 10 9 10 9 0 2 13 15 10 9 1 10 9 1 9 0 2
46 10 9 1 10 9 1 10 9 1 11 2 11 11 2 4 13 10 11 16 13 10 9 1 13 10 10 9 0 0 1 13 10 9 1 10 9 0 1 10 9 1 9 1 10 11 2
28 0 9 4 13 1 11 2 11 2 11 2 11 2 11 7 11 2 16 1 11 7 11 10 9 15 13 0 2
29 1 9 2 15 13 13 10 9 16 13 10 0 9 2 9 7 8 2 9 7 10 9 1 9 16 13 1 15 2
22 3 13 0 13 15 2 1 15 15 3 13 10 9 16 13 13 7 15 13 1 11 2
19 15 13 3 1 10 9 2 7 10 9 3 3 13 13 10 9 7 13 2
55 10 9 1 11 11 2 1 12 9 2 4 13 1 12 9 1 9 3 1 10 9 1 10 11 2 1 10 9 1 10 9 1 10 9 2 3 13 10 9 1 13 1 10 9 2 16 13 0 2 13 10 9 0 0 2
88 10 9 1 11 4 13 10 9 9 1 9 1 3 15 13 10 9 7 3 15 13 1 10 0 12 9 1 10 9 1 11 7 1 10 12 9 1 10 9 9 1 10 9 11 2 1 10 12 9 2 7 13 16 4 13 3 0 1 15 16 3 15 13 1 15 7 15 1 10 15 2 16 1 10 9 1 10 11 3 4 13 15 10 9 3 2 2 2
21 13 10 0 9 1 10 16 13 7 1 10 0 9 15 13 10 15 16 4 13 2
13 13 15 10 9 13 7 15 13 10 9 13 2 2
28 1 15 1 10 9 1 10 13 1 10 9 13 3 10 9 13 10 9 1 9 1 10 9 1 9 1 9 2
27 10 9 1 11 2 16 13 10 12 1 11 2 13 12 9 1 9 2 13 1 9 0 1 9 7 9 2
46 1 10 9 2 10 9 1 10 9 4 13 16 10 9 15 13 1 13 1 9 1 10 10 9 16 15 4 13 1 9 7 10 15 13 3 0 2 1 10 9 1 10 12 1 11 2
34 11 13 1 9 1 10 9 12 9 16 4 13 1 10 9 16 1 9 2 3 4 13 0 7 3 15 13 1 10 9 16 4 13 2
50 10 9 4 13 16 2 15 9 2 13 16 10 9 2 13 2 7 2 13 1 10 9 2 2 7 2 10 9 13 15 16 13 2 7 1 15 4 7 13 1 3 1 13 10 9 2 2 4 13 2
31 10 8 1 10 9 2 16 13 10 9 1 11 1 10 11 2 13 10 9 16 4 1 13 15 1 11 1 10 0 9 2
25 3 15 13 13 10 9 1 9 1 10 9 2 15 13 16 15 13 10 9 0 2 13 10 9 2
16 3 13 10 9 0 7 16 3 4 13 13 1 10 12 9 2
32 10 9 13 2 15 13 16 10 9 1 10 9 4 1 13 10 9 1 10 9 1 11 1 10 9 13 1 10 9 1 9 2
33 10 9 1 10 9 1 10 9 0 2 3 3 1 10 9 2 13 10 9 0 2 10 9 0 16 1 10 0 9 15 4 13 2
21 10 8 1 11 2 11 7 11 13 13 1 9 0 10 9 1 10 11 1 11 2
36 10 9 15 13 10 9 7 9 1 0 9 7 2 1 10 13 1 10 15 2 10 9 4 13 1 13 15 2 15 15 13 2 3 0 2 2
24 10 9 1 9 1 0 9 1 10 9 1 9 8 1 10 0 9 13 0 1 13 10 9 2
51 1 10 9 9 0 1 10 9 0 1 9 2 13 13 10 9 11 11 1 13 1 10 9 16 10 9 1 11 11 13 1 10 9 10 9 13 1 11 2 7 13 0 9 1 9 7 9 1 11 11 2
31 10 9 16 3 13 9 2 10 11 2 15 13 1 13 11 7 10 9 0 1 13 15 1 10 9 1 10 9 1 11 2
41 10 9 0 2 13 13 2 10 0 9 1 9 16 13 2 10 13 3 13 10 9 7 10 9 1 10 0 9 1 9 2 15 13 3 1 10 2 9 0 2 2
15 13 10 9 3 13 13 15 1 10 10 9 1 9 2 2
40 10 9 13 10 11 1 11 11 11 1 10 11 11 13 1 9 0 7 15 13 10 9 0 1 0 7 0 2 10 0 9 0 1 11 15 13 11 11 11 2
13 10 9 3 13 10 0 9 16 13 1 10 9 2
51 10 9 11 11 13 10 11 10 9 1 10 16 13 0 3 10 0 9 1 9 1 9 1 9 2 10 15 13 10 9 0 1 10 9 1 10 10 9 1 9 1 13 15 1 10 12 9 7 9 0 2
54 10 9 11 2 16 13 9 1 10 0 9 2 13 12 9 1 9 15 4 4 3 13 3 1 11 11 2 9 1 10 11 2 2 7 4 13 1 10 9 1 0 9 7 9 13 1 10 9 1 10 9 11 11 2
70 10 9 0 1 11 15 13 1 12 9 1 9 2 1 10 16 13 12 9 1 9 2 1 10 9 1 9 1 12 9 1 9 2 16 7 10 9 0 1 11 1 11 15 13 1 12 9 1 9 2 1 10 16 13 12 9 1 9 2 1 10 9 1 9 1 12 9 1 9 2
44 1 10 9 1 10 9 1 13 10 9 1 11 1 9 1 10 9 2 10 9 15 13 1 13 16 13 3 2 15 16 13 2 16 11 13 1 10 9 1 10 9 1 11 2
47 2 10 9 1 10 9 4 13 3 10 9 1 10 9 1 10 11 1 13 10 9 7 4 13 10 9 1 16 11 4 13 3 10 9 16 13 1 10 10 9 1 10 9 2 2 13 2
18 10 9 16 13 11 11 10 0 9 1 11 13 10 9 1 10 9 2
45 10 9 1 9 1 9 1 8 1 1 12 9 1 9 2 13 13 2 15 16 1 9 0 4 13 15 1 10 9 8 2 13 10 9 1 10 12 5 1 10 0 9 1 11 2
33 13 16 1 10 9 0 9 12 2 10 9 13 1 10 9 0 13 11 11 2 1 10 9 0 2 3 7 13 12 9 1 9 2
29 1 9 2 10 9 0 4 13 16 10 9 16 13 10 9 0 13 1 10 9 7 15 15 13 1 9 1 9 2
43 10 11 4 1 13 10 12 0 9 1 10 9 13 1 11 2 15 15 13 1 11 2 11 2 7 15 1 10 9 8 2 12 2 1 10 9 1 10 11 2 1 11 2
76 10 9 16 3 4 13 1 0 9 2 3 4 13 12 2 7 1 10 9 3 13 1 9 2 7 16 4 13 2 7 3 1 9 7 3 1 9 2 3 1 10 9 1 3 2 10 9 13 16 3 4 13 9 1 15 2 3 4 1 13 16 4 13 1 9 2 7 1 3 7 3 0 3 4 13 2
10 9 1 9 7 9 1 10 9 0 2
15 15 13 16 13 10 0 9 2 7 16 3 13 3 0 2
19 13 10 9 7 3 15 13 10 9 2 1 3 13 7 13 1 13 9 2
37 0 13 10 9 1 15 16 15 4 13 10 9 7 9 1 9 2 15 13 10 9 1 1 9 16 15 15 13 15 1 10 9 1 10 0 9 2
10 16 13 10 9 2 15 13 10 9 2
3 15 13 2
33 13 9 1 10 0 9 1 9 7 9 1 9 2 15 16 15 13 13 10 0 9 7 13 15 1 15 10 9 13 15 16 13 2
19 13 1 0 9 2 3 9 15 8 3 3 13 8 9 7 13 15 9 2
15 3 0 16 13 10 9 1 10 9 1 0 9 7 9 2
7 15 13 16 15 13 13 2
12 9 16 13 3 0 7 1 9 3 13 9 2
15 10 9 13 3 0 2 0 7 13 13 10 10 0 9 2
26 4 13 10 9 2 7 15 3 4 13 9 1 10 9 3 0 16 13 1 9 2 10 9 1 9 2
5 3 13 10 9 2
10 4 1 13 2 0 9 7 0 9 2
12 3 15 13 10 9 7 15 13 1 10 9 2
19 10 9 13 0 2 1 12 7 12 5 1 9 2 7 10 9 13 0 2
23 10 9 13 3 0 7 3 2 1 1 10 10 9 3 15 13 15 2 4 7 13 9 2
18 10 9 10 9 2 10 9 3 0 2 1 9 3 0 7 0 9 2
4 15 15 13 3
21 14 2 10 9 0 13 10 9 1 9 8 2 7 13 3 0 7 10 1 11 2
23 10 9 0 13 1 10 9 1 9 1 10 9 1 13 10 9 7 10 9 1 10 9 2
17 1 11 11 4 13 10 9 0 3 0 2 0 7 1 0 9 2
5 13 0 10 8 2
9 1 3 9 13 1 10 9 0 2
22 4 13 1 13 10 0 9 1 9 1 13 3 1 10 9 0 16 3 13 10 11 11
46 1 9 13 1 0 9 16 3 15 13 3 9 7 15 13 1 10 12 1 13 10 9 2 16 1 11 3 13 7 3 1 13 15 7 1 13 15 10 0 9 3 15 13 10 9 2
8 3 13 15 0 9 1 9 2
19 13 1 15 3 9 16 15 4 13 3 3 1 11 13 1 10 10 9 2
19 10 9 13 10 9 1 9 0 9 0 8 8 1 13 15 7 1 10 9
9 15 3 13 16 15 13 10 9 2
18 10 9 13 0 2 7 1 15 2 3 2 10 9 15 13 3 0 2
25 10 9 13 10 9 0 2 3 13 10 9 0 1 15 1 10 9 2 1 15 9 16 13 11 2
12 10 9 0 13 16 3 16 15 13 13 0 2
13 16 4 13 10 9 1 11 2 3 15 4 13 2
6 1 10 12 15 13 2
8 15 4 13 10 9 7 9 2
12 10 9 13 3 0 1 10 9 1 10 9 2
11 1 9 10 2 15 13 1 10 12 5 2
5 10 9 13 8 2
16 10 0 9 1 10 9 16 4 13 2 10 9 1 9 0 2
17 1 9 1 13 0 2 13 10 9 7 9 1 11 1 10 9 2
27 13 9 16 10 9 13 1 8 1 11 11 13 9 0 1 0 9 16 2 1 9 0 13 9 1 11 2
14 13 10 9 0 13 1 0 11 1 11 10 9 13 12
16 16 10 9 1 10 9 15 13 10 12 5 13 3 10 9 2
9 3 10 9 7 10 9 13 0 2
12 13 10 9 1 10 9 7 1 10 9 3 0
8 13 9 1 13 13 1 3 2
21 13 13 2 16 1 10 9 15 13 10 9 1 7 3 13 9 7 13 10 9 2
9 15 9 16 10 9 3 13 0 2
22 13 3 3 0 7 3 16 15 13 10 9 2 4 13 10 9 1 13 10 9 8 2
11 3 13 13 1 13 1 9 10 10 9 2
6 10 9 15 13 0 2
5 1 9 2 9 2
19 1 9 13 10 9 1 10 9 1 10 9 16 13 13 9 1 10 9 2
6 0 9 2 9 0 2
25 10 0 8 8 16 4 13 2 13 9 1 9 2 7 10 9 0 1 13 15 1 9 0 7 0
54 15 9 0 3 13 10 9 1 9 2 13 1 10 9 2 13 3 2 2 2 16 10 11 2 16 13 1 10 10 9 1 10 9 1 9 7 9 2 13 3 0 7 15 13 13 7 10 9 4 1 13 1 13 2
19 10 9 8 8 4 13 1 12 1 12 9 1 12 9 2 10 12 5 2
17 4 13 1 9 1 11 1 12 7 4 13 10 9 0 2 13 2
4 13 3 0 2
10 10 3 0 2 7 13 3 10 9 2
21 10 9 2 10 9 2 10 9 2 9 0 7 3 0 2 0 9 2 9 1 9
21 10 9 1 11 15 4 13 1 10 8 5 12 1 10 9 11 11 2 1 11 11
17 9 1 11 2 10 8 2 1 10 9 1 16 15 13 3 3 2
10 0 9 1 13 15 7 13 10 9 5
55 13 13 10 9 7 15 2 13 10 9 9 1 12 9 2 15 3 0 2 9 7 9 2 13 10 9 1 9 2 16 3 15 13 3 10 9 2 13 10 9 1 9 1 10 9 3 2 1 9 2 3 13 7 13 2
58 10 9 13 1 10 9 1 16 10 0 9 0 1 10 9 15 13 1 9 1 9 0 7 1 9 16 2 1 10 0 9 2 13 0 1 13 1 15 7 1 10 9 2 1 0 2 1 10 9 2 1 15 13 1 10 9 11 2
15 10 9 13 1 10 9 1 10 11 7 15 13 9 1 9
15 0 9 13 10 3 0 1 15 16 13 7 3 13 0 2
6 3 4 13 10 9 2
21 15 13 10 9 1 10 9 1 10 9 2 3 13 0 2 7 15 13 10 9 2
6 3 4 13 10 9 2
11 10 9 13 3 0 7 13 13 1 9 2
13 13 1 7 15 4 4 13 1 10 9 1 9 2
