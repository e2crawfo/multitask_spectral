138 11
24 2 3 3 9 10 9 9 2 10 9 15 13 2 16 10 0 9 7 10 9 13 10 9 2
16 3 7 11 9 13 10 9 2 7 0 9 13 10 12 9 2
14 2 3 10 11 13 10 9 2 7 10 9 9 13 2
8 15 13 10 9 10 0 9 2
33 2 15 7 3 13 2 7 3 10 9 0 0 9 3 3 13 10 9 2 7 3 15 7 0 9 2 16 3 13 10 11 11 2
14 12 9 1 11 3 0 13 2 16 15 3 13 9 2
11 2 0 0 9 1 0 13 3 10 9 2
3 2 3 2
22 12 9 12 9 9 13 2 15 11 13 10 9 2 3 7 16 13 4 2 3 13 2
13 3 13 2 0 0 9 1 13 3 10 9 3 2
26 16 10 0 11 13 10 9 0 12 9 9 2 3 3 10 0 9 1 13 15 10 0 9 0 9 2
5 10 0 9 1 2
28 3 3 13 15 11 11 2 15 10 9 0 0 9 0 9 13 10 9 2 7 15 3 3 10 0 0 11 2
9 10 9 11 11 9 13 10 9 2
15 10 9 0 9 10 0 9 0 0 9 7 0 9 13 2
10 7 2 11 9 2 3 13 10 9 2
22 2 13 3 10 9 2 10 9 13 10 15 9 2 16 10 0 9 2 10 9 13 2
19 3 13 10 11 9 2 7 11 7 11 3 3 3 0 3 2 16 15 2
40 13 10 9 2 0 9 2 0 9 2 7 3 0 9 1 2 16 10 11 2 3 13 2 13 0 9 1 11 2 15 3 13 2 16 3 11 11 9 13 2
17 10 11 11 9 2 11 11 7 10 9 0 9 1 0 9 13 2
9 10 9 9 1 13 10 0 9 2
14 10 9 10 11 11 11 13 2 15 3 0 9 13 2
6 9 9 2 0 9 9
28 2 15 3 13 3 2 16 0 9 13 11 2 2 13 11 2 2 7 3 13 13 2 3 3 9 10 9 2
16 10 9 3 13 2 7 10 9 9 9 0 9 13 10 11 2
28 0 3 3 13 4 10 0 9 0 9 2 10 0 9 2 9 13 10 0 0 9 2 9 3 10 0 9 2
23 10 9 11 11 13 2 15 10 0 12 9 9 13 3 10 0 0 9 9 1 10 9 2
40 10 9 12 0 9 0 10 0 0 1 13 2 13 3 9 2 7 9 13 10 9 9 1 9 2 11 11 7 15 15 7 0 9 2 7 9 15 3 13 2
24 3 3 13 4 2 3 10 9 3 13 2 10 9 9 2 10 9 0 9 2 11 11 7 2
21 15 7 3 13 2 3 13 3 10 9 12 9 0 12 9 2 11 11 7 3 2
40 10 0 0 9 0 9 7 3 0 0 9 13 10 9 1 2 10 0 0 9 0 9 3 15 10 0 0 9 11 11 2 7 10 7 9 0 11 11 1 2
23 7 3 3 13 9 2 9 11 12 9 13 3 15 2 15 3 12 9 13 15 0 9 2
11 15 3 2 11 10 9 0 9 13 15 2
23 7 10 9 0 12 9 3 3 10 0 9 13 12 9 0 2 7 0 9 7 13 15 2
29 2 9 2 11 7 3 4 13 10 12 9 2 13 3 15 11 2 13 0 10 9 1 10 9 0 9 0 11 2
4 2 3 3 2
28 10 0 9 3 3 15 13 2 16 10 0 0 0 9 2 3 3 13 0 10 0 9 2 15 7 3 13 2
24 7 16 3 7 3 13 2 7 13 10 9 2 3 3 13 10 9 15 2 15 10 3 13 2
13 11 9 3 13 10 11 3 0 9 0 0 9 2
24 10 15 9 3 10 3 0 0 2 9 2 13 2 7 10 3 3 0 9 13 10 0 9 2
23 16 3 3 10 9 0 9 7 13 2 7 10 0 9 0 9 0 0 13 10 0 9 2
13 0 13 9 10 0 9 0 9 0 9 11 1 2
7 10 0 9 9 9 13 2
15 10 0 0 9 0 9 0 9 13 10 12 9 0 9 2
25 10 9 10 0 9 12 0 9 13 3 2 11 11 12 9 13 2 10 10 9 2 11 11 12 2
11 10 9 0 11 11 7 10 9 0 0 2
16 10 0 9 0 2 0 9 13 2 10 9 9 13 2 3 2
35 10 0 9 13 10 3 10 12 0 9 2 10 11 7 10 11 9 0 0 9 2 9 2 2 7 9 13 13 10 0 9 2 9 2 2
27 11 7 11 11 7 13 0 0 9 2 10 11 9 3 3 13 10 9 0 9 0 0 9 2 11 11 2
15 10 9 13 10 9 2 7 10 12 0 9 7 9 13 2
16 15 1 13 10 2 9 2 2 10 12 0 9 2 9 2 2
27 3 13 10 9 9 2 11 9 2 13 9 10 10 9 2 0 10 9 9 1 2 3 15 7 13 9 2
12 7 3 15 7 2 16 10 0 9 11 13 2
11 12 7 12 9 10 9 1 11 9 13 2
17 7 10 9 13 15 2 12 9 1 12 0 13 9 2 9 2 2
21 9 0 9 13 3 10 9 9 2 15 1 13 12 9 0 9 13 2 9 2 2
14 0 9 9 11 11 1 13 9 2 9 11 13 11 2
18 9 9 7 0 13 10 9 2 11 2 11 9 2 11 12 9 13 2
21 10 9 0 9 11 11 2 15 3 3 13 14 10 9 0 0 9 2 13 11 2
29 10 9 0 9 10 9 12 0 0 9 9 1 7 10 10 12 10 9 13 0 2 15 3 0 13 10 0 9 2
31 10 0 11 11 10 9 2 10 9 2 10 9 0 2 3 10 0 12 9 10 9 9 0 11 11 10 9 2 10 9 2
47 10 9 9 2 15 0 7 13 2 3 13 10 11 11 2 9 3 10 9 7 0 13 10 9 0 9 0 11 11 1 2 7 10 9 9 11 7 9 1 0 0 9 9 13 10 9 2
23 0 2 3 12 9 12 9 9 13 14 15 10 9 0 0 11 11 2 9 2 9 2 2
41 3 13 10 9 10 9 2 10 0 11 9 2 15 0 9 13 2 16 12 9 9 11 9 2 7 11 13 0 12 9 7 2 10 0 9 2 11 11 7 11 2
13 11 3 3 9 2 11 13 13 2 7 3 3 2
17 10 0 12 9 11 13 2 3 9 13 9 2 7 9 3 3 2
18 0 3 13 10 0 9 7 2 7 3 12 9 1 9 2 9 13 2
31 9 0 9 2 12 2 2 0 9 12 2 7 3 3 0 9 2 12 2 7 10 13 11 2 15 10 0 3 12 13 2
41 2 13 2 16 11 13 15 9 13 10 9 2 16 0 13 2 7 16 13 10 9 2 13 10 9 2 7 15 13 2 16 3 3 13 3 10 9 2 13 11 2
27 2 11 3 12 9 13 10 0 12 9 2 13 2 16 9 13 12 9 1 2 10 0 9 9 3 13 2
17 13 10 9 13 10 9 2 7 3 3 13 3 2 16 13 11 2
6 10 10 9 0 13 2
14 15 9 13 15 3 2 3 15 13 15 10 0 9 2
29 2 11 3 3 13 3 10 9 2 3 13 2 7 3 9 13 2 0 13 13 10 9 2 3 13 10 0 11 2
25 2 10 0 9 7 13 2 16 13 2 3 3 0 10 9 2 7 10 0 9 7 0 13 3 2
7 3 0 2 13 2 15 2
22 15 10 12 12 9 1 0 11 11 2 11 11 7 11 9 2 11 11 13 10 3 2
5 3 13 11 13 2
47 10 11 11 11 2 11 9 13 14 11 11 9 2 10 12 0 9 1 0 9 0 9 7 10 9 2 7 11 11 0 9 0 9 0 9 2 9 2 11 11 0 9 0 9 10 9 2
34 10 9 13 2 16 11 11 9 7 9 2 11 11 9 2 7 10 3 3 0 9 1 10 0 9 3 0 12 9 9 13 3 9 2
6 10 9 7 9 13 2
29 10 11 11 10 9 0 7 0 9 1 9 1 13 10 9 2 7 0 9 9 2 0 9 9 13 10 0 9 2
20 3 10 11 11 11 9 13 11 11 1 11 11 0 9 9 7 9 9 1 2
8 10 12 9 0 13 10 9 2
18 10 9 1 11 11 7 11 11 10 0 9 9 10 9 13 3 3 2
15 11 11 12 9 13 10 0 9 2 15 13 10 9 1 2
7 0 9 2 11 11 13 2
26 3 11 2 15 0 9 2 16 9 13 2 3 13 3 3 12 10 0 9 2 12 9 13 11 11 2
18 10 9 11 1 10 9 13 2 3 10 9 3 10 0 9 13 3 2
24 11 11 0 10 9 15 13 2 16 10 12 9 9 2 11 13 10 0 9 0 12 0 9 2
9 13 2 13 7 9 13 0 9 2
21 10 9 2 16 11 13 9 2 11 9 13 2 7 13 10 11 11 1 0 9 2
9 3 13 2 7 10 9 15 13 2
7 11 11 3 3 13 3 2
18 10 12 9 3 3 3 13 10 9 9 2 7 12 12 9 9 13 2
17 12 9 3 13 2 9 13 10 9 11 9 2 16 13 10 9 2
23 10 0 9 3 12 12 9 13 2 7 10 0 9 3 13 3 2 3 3 3 3 13 2
20 11 11 10 0 0 9 13 2 16 3 13 9 13 2 7 3 13 15 0 2
11 10 9 1 9 9 9 13 10 0 9 2
41 11 11 2 9 1 0 9 9 0 9 13 10 11 11 9 10 0 0 9 2 15 9 10 11 11 11 2 10 11 11 11 2 11 2 7 11 11 0 9 13 2
12 9 11 11 12 9 13 3 0 9 9 1 2
39 10 11 11 11 9 1 3 12 9 3 13 9 2 15 9 13 10 10 9 2 16 9 11 11 10 9 0 9 9 7 0 9 9 7 9 1 0 9 2
19 10 9 1 10 9 0 9 9 9 13 3 10 9 2 15 3 13 9 2
19 10 11 11 11 9 15 1 10 11 11 11 13 7 13 10 9 9 9 2
9 11 11 10 9 9 13 10 9 2
9 11 11 7 3 13 3 10 9 2
16 11 11 13 2 9 7 15 9 3 2 16 0 13 15 3 2
8 10 9 0 9 9 13 3 2
16 3 10 0 9 2 9 11 11 3 0 2 9 7 0 13 2
9 10 9 10 9 0 9 1 13 2
13 10 11 11 11 0 9 7 10 0 9 13 9 2
27 13 10 9 10 0 9 9 2 0 9 0 9 2 12 9 1 2 7 12 12 9 9 2 0 9 9 2
25 3 10 9 9 13 2 11 3 13 0 9 2 16 9 2 9 7 3 13 3 10 9 0 9 2
10 10 9 9 3 13 9 10 11 11 2
11 10 0 9 0 9 10 0 9 9 13 2
10 10 0 9 0 9 7 9 1 13 2
25 10 11 11 11 2 11 2 9 12 9 13 2 10 9 1 3 3 13 3 10 11 0 0 9 2
42 3 0 2 16 10 9 10 9 9 13 2 13 14 11 11 2 10 11 9 9 2 15 1 12 9 13 3 2 16 0 9 7 9 1 13 4 13 10 0 9 9 2
12 10 9 3 3 10 9 9 1 13 0 9 2
17 7 15 7 13 2 16 15 0 0 2 0 9 1 13 9 9 2
18 0 9 13 10 11 9 1 2 3 10 0 9 13 10 11 0 9 2
27 15 7 3 10 9 0 2 12 9 0 12 9 0 9 13 2 7 12 9 9 2 9 3 12 9 2 2
24 10 9 9 3 3 15 13 3 2 16 11 11 2 10 0 9 3 3 0 9 13 10 9 2
25 10 9 0 9 1 13 3 10 9 2 10 9 7 15 13 10 9 2 16 10 9 3 13 3 2
12 10 0 9 0 13 2 3 3 13 10 9 2
17 10 11 0 9 9 1 12 9 9 13 10 11 0 9 10 9 2
22 11 11 9 10 9 13 2 16 15 3 10 0 0 9 13 4 2 7 0 9 13 2
12 10 9 10 9 0 0 9 13 13 10 9 2
20 3 13 2 9 12 12 9 13 2 15 3 3 11 11 10 0 0 9 13 2
20 12 2 9 0 0 0 9 13 9 9 3 10 9 10 9 2 10 0 9 2
34 10 9 0 9 13 10 0 9 10 10 12 9 2 15 1 10 15 2 3 10 9 1 2 9 13 2 10 15 7 0 9 13 9 2
22 10 12 9 2 10 9 1 2 10 16 12 9 13 3 9 7 9 10 0 11 9 2
14 10 9 12 9 9 13 10 0 9 2 3 13 15 2
9 9 13 3 3 10 0 9 9 2
31 10 0 9 2 15 10 0 9 13 2 9 13 2 7 16 10 9 3 13 3 2 3 3 13 2 10 9 9 9 13 2
23 10 0 9 10 9 12 12 1 13 13 2 10 0 9 9 7 0 9 13 10 9 9 2
36 10 9 13 10 0 2 10 0 7 10 0 9 7 2 10 0 9 1 7 3 10 9 13 3 10 9 2 7 3 3 10 9 13 10 9 2
19 0 9 3 13 2 10 9 9 2 9 10 9 1 10 9 9 7 13 2
