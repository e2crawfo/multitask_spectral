150 17
32 13 9 9 13 9 8 12 15 1 9 9 10 9 0 7 13 9 9 7 9 1 9 1 8 2 9 10 11 7 9 9 2
29 13 9 1 9 14 13 9 10 9 1 2 13 1 2 1 9 0 14 13 15 7 13 15 10 9 1 9 1 2
8 13 10 9 14 13 10 9 2
6 9 9 1 9 1 2
6 14 13 15 14 0 2
27 13 9 0 13 0 12 9 14 9 1 9 0 1 9 16 3 14 13 15 9 14 13 9 1 10 9 2
25 9 1 9 9 1 8 10 9 0 7 10 11 2 9 7 9 9 2 13 9 10 9 1 9 2
6 13 15 1 1 9 2
10 13 1 10 9 16 14 13 15 9 2
12 13 15 1 9 1 9 11 1 12 1 12 2
22 13 9 0 1 10 9 0 2 13 9 10 9 1 9 7 13 10 9 0 7 0 2
56 9 0 13 0 1 14 9 1 9 1 1 14 13 3 2 2 7 16 13 9 0 10 9 7 13 9 2 16 13 15 2 14 9 0 2 14 9 0 10 9 3 2 7 14 13 9 0 1 3 0 7 14 13 15 3 2
27 13 9 9 7 9 1 2 13 10 9 1 9 2 7 13 10 9 1 9 9 10 9 1 9 10 9 2
31 1 9 13 15 3 7 13 15 2 13 9 1 14 11 2 14 13 15 1 9 1 1 12 9 10 14 13 15 9 1 2
10 2 1 9 2 13 3 2 14 9 2
36 8 1 9 10 9 0 7 2 1 9 15 2 1 10 9 1 9 0 2 13 9 9 1 9 2 1 10 9 7 10 9 9 2 1 9 2
19 16 14 13 10 9 1 9 13 9 1 9 10 9 10 16 9 0 1 2
17 2 13 10 9 10 0 14 14 13 15 1 2 2 14 13 15 2
27 13 1 10 9 10 14 0 14 13 10 9 1 9 7 13 1 10 9 10 14 0 14 13 9 10 9 2
55 2 11 14 13 1 10 9 0 14 13 1 9 14 0 1 9 9 14 9 1 1 9 10 13 1 11 16 13 9 1 9 0 0 1 9 9 11 1 12 9 3 7 16 13 9 1 3 16 13 11 10 9 1 9 2
21 1 9 10 9 13 10 9 1 10 9 0 7 13 10 11 1 9 0 7 0 2
34 3 13 3 15 9 9 14 13 1 9 1 10 9 1 10 9 10 7 13 9 1 10 9 9 0 7 10 9 13 0 1 9 12 2
30 1 10 9 10 2 13 11 1 9 1 9 7 9 1 10 8 16 13 15 1 10 9 16 3 2 3 2 14 13 2
13 13 1 9 7 9 8 15 14 0 7 14 0 2
51 13 3 2 1 15 2 1 9 1 10 9 14 13 1 10 11 14 9 1 9 1 9 9 7 9 1 9 1 9 14 13 1 10 9 10 9 9 2 1 9 1 9 2 14 9 1 9 3 0 15 2
28 16 13 10 9 1 1 9 10 9 2 7 1 9 1 10 9 1 2 13 14 13 10 9 0 3 0 1 2
12 13 9 0 1 9 10 9 1 10 9 10 2
2 13 2
38 1 9 10 9 3 2 13 9 1 9 11 3 1 9 9 0 7 1 9 1 9 1 1 9 10 11 1 9 2 13 9 0 1 1 9 10 9 2
19 16 13 0 3 1 9 13 9 1 13 9 14 13 10 9 1 10 9 2
2 13 2
3 10 9 2
47 16 13 13 1 9 9 11 11 2 10 11 0 2 14 13 10 9 2 9 14 13 14 13 1 9 11 10 9 9 14 9 1 15 1 9 1 9 7 9 10 9 1 9 1 10 9 2
14 1 15 13 9 1 9 3 1 10 9 9 1 9 2
48 9 9 14 13 9 1 9 1 9 7 9 10 1 9 2 15 9 2 1 9 9 9 1 9 7 9 2 13 15 9 0 0 14 13 9 9 0 1 2 9 14 13 3 3 1 9 9 2
35 2 9 9 14 13 3 0 15 1 2 13 9 1 9 1 1 9 1 9 0 2 7 1 9 15 13 1 9 9 14 13 1 9 2 2
29 13 1 10 9 14 13 9 1 9 10 9 14 0 14 13 1 9 3 2 16 13 10 9 0 1 10 9 0 2
69 13 10 9 14 13 1 10 9 3 2 2 10 9 2 2 10 9 14 13 11 14 11 10 9 13 0 1 9 2 1 9 3 2 9 12 9 3 1 9 1 9 9 7 9 10 11 7 9 9 1 9 11 10 11 14 13 9 11 1 14 9 1 9 1 1 10 9 0 2
3 2 9 2
11 13 9 1 14 13 9 9 1 9 1 2
2 7 2
3 2 3 2
3 15 15 2
13 15 1 9 14 9 2 14 13 15 1 10 9 2
5 3 14 13 15 2
7 9 0 0 14 13 1 2
12 13 10 9 10 9 1 9 0 1 9 0 2
3 9 12 2
36 1 11 13 1 9 1 11 15 1 9 1 10 11 1 12 9 12 2 9 14 13 15 2 16 13 9 2 14 13 1 10 9 9 1 9 2
32 13 15 13 9 1 2 9 14 13 9 9 1 1 10 9 0 14 9 2 9 14 13 9 1 9 0 1 9 10 9 10 2
44 13 0 14 13 1 9 10 9 2 9 0 7 0 14 9 7 14 9 7 9 14 9 1 2 9 14 13 10 9 7 10 9 14 9 7 14 9 7 9 3 14 9 1 2
19 13 10 9 9 1 2 13 10 9 9 2 16 9 1 9 14 9 1 2
7 13 10 9 0 1 11 2
28 16 14 13 10 9 0 3 2 13 15 1 10 11 11 11 7 1 1 9 13 15 1 11 1 9 10 9 2
11 13 10 9 1 9 1 9 7 13 9 2
6 13 15 11 10 9 2
35 13 10 9 0 1 9 1 10 9 0 7 13 15 14 0 14 13 15 1 9 14 13 15 10 9 1 7 14 13 15 9 0 1 1 2
39 13 10 9 1 11 2 9 9 9 2 9 7 9 3 7 3 10 9 7 9 1 10 9 7 13 9 10 9 3 1 9 10 9 1 9 1 14 12 2
11 13 9 0 1 9 0 14 13 9 0 2
20 13 9 3 1 9 1 9 9 14 13 15 1 10 9 1 1 10 9 0 2
5 13 15 10 9 2
22 3 2 3 2 13 3 10 9 10 14 13 9 10 9 0 1 2 7 13 3 2 2
7 2 13 10 9 14 0 2
11 13 0 1 9 7 9 0 10 12 9 2
19 13 15 3 10 9 9 1 8 7 10 9 14 13 1 9 1 9 10 2
14 1 9 10 9 9 2 13 9 0 2 9 0 3 2
38 9 13 1 9 10 10 9 10 14 9 1 7 13 0 15 2 16 15 14 9 1 9 1 9 10 1 9 1 15 14 9 1 10 9 1 9 9 2
6 9 12 2 9 9 2
11 13 10 10 9 9 1 9 1 9 9 2
36 13 0 14 13 15 9 14 9 14 0 14 13 15 0 1 9 2 9 1 10 9 14 13 9 0 2 1 14 13 15 3 12 9 9 9 2
6 13 10 9 9 9 2
20 13 11 11 2 12 9 1 9 1 12 9 1 9 9 7 9 14 13 11 2
15 13 9 9 7 9 1 12 9 9 7 12 9 14 9 2
17 1 15 1 11 2 9 14 13 9 0 1 12 9 1 9 0 2
12 13 15 1 9 1 9 10 9 2 11 0 2
24 13 9 10 9 3 7 14 13 10 9 2 7 2 9 2 10 2 16 15 0 1 10 9 2
23 13 9 9 3 1 9 10 9 7 13 9 1 9 0 1 9 9 3 1 3 10 9 2
36 13 10 9 16 14 13 1 1 9 2 16 14 13 15 9 14 13 0 7 0 2 7 16 14 13 9 0 10 9 1 10 9 7 10 9 2
42 2 13 10 9 15 14 13 1 9 3 0 15 1 9 10 9 1 9 7 14 13 1 9 1 9 1 9 9 10 9 1 9 7 9 9 10 9 7 9 1 9 2
24 1 9 2 13 9 10 1 14 13 10 9 1 9 14 13 9 10 11 1 11 2 9 9 2
13 13 9 9 1 2 9 14 13 9 1 10 9 2
5 13 15 3 15 2
6 13 9 9 9 1 2
32 9 9 9 13 15 15 10 9 9 9 2 2 8 9 2 8 9 2 8 9 2 8 9 7 9 2 8 9 2 8 9 2
37 9 16 14 13 10 9 0 1 9 1 2 3 13 9 1 9 2 13 9 16 9 1 10 9 9 1 11 11 2 7 10 9 1 9 9 0 2
10 13 11 10 9 0 1 10 9 9 2
4 13 0 0 2
66 8 13 1 9 9 14 13 10 9 7 13 1 12 9 0 14 9 15 2 16 13 9 0 7 12 9 0 14 9 1 9 2 7 14 13 15 1 9 9 1 9 7 1 9 10 10 9 1 9 1 9 1 10 9 13 1 9 0 7 12 9 0 14 13 15 2
21 16 10 9 1 11 11 2 11 2 2 13 15 1 9 15 7 13 15 10 9 2
5 13 15 1 9 2
2 9 2
23 13 10 9 0 1 11 2 7 13 0 1 14 13 15 7 10 9 9 1 9 9 1 2
14 13 15 9 3 1 9 10 9 2 1 9 11 11 2
10 9 0 2 10 9 1 14 13 1 2
50 8 1 10 9 10 14 13 14 9 1 9 9 8 2 2 8 8 13 10 11 9 1 9 1 9 8 7 10 9 13 1 14 9 1 9 1 9 14 13 7 1 9 7 1 9 2 16 9 2 2
31 13 15 9 11 11 13 9 1 9 10 9 10 1 9 2 13 1 15 2 2 9 0 0 10 9 13 0 1 10 9 2
4 13 11 0 2
8 13 15 10 9 10 10 9 2
4 9 14 9 2
61 13 0 14 13 1 9 10 9 2 1 9 0 9 2 10 9 14 9 2 14 9 2 14 9 1 9 7 14 9 7 9 14 9 1 9 0 0 2 8 2 8 2 1 9 14 9 1 9 14 9 2 9 9 14 9 1 9 7 1 9 2
7 1 12 9 13 15 3 2
46 1 9 0 13 9 1 9 1 9 10 9 11 1 10 9 1 9 11 1 10 9 7 13 9 1 0 14 13 9 0 1 9 1 10 9 10 16 14 13 1 10 9 0 14 0 2
14 2 2 15 9 14 13 10 9 10 1 9 11 9 2
35 13 9 1 12 9 9 1 9 13 1 9 1 9 1 2 10 9 0 10 1 9 2 2 0 9 1 13 0 1 11 2 15 15 15 2
17 1 9 2 1 9 2 7 15 16 13 15 14 0 1 10 9 2
16 13 10 9 0 1 9 10 9 9 2 7 1 9 10 9 2
20 14 13 11 14 11 14 13 10 9 0 1 9 1 9 1 9 10 9 10 2
40 13 15 0 14 13 10 9 1 10 9 1 9 0 7 13 0 10 9 9 1 10 9 9 1 9 1 10 9 16 13 10 9 1 9 2 2 13 10 11 2
12 11 7 10 9 14 13 1 1 9 13 3 2
22 13 15 15 7 16 14 13 10 9 1 14 13 10 9 2 13 15 15 14 9 0 2
8 9 9 7 9 13 3 1 2
17 13 15 10 9 11 7 9 10 11 11 14 13 1 10 9 10 2
46 1 9 10 9 14 13 9 1 9 1 10 9 9 1 2 13 9 14 13 1 10 9 7 10 9 2 9 9 9 14 13 1 9 7 11 2 9 9 1 9 9 2 0 7 11 2
4 13 15 3 2
26 16 14 13 15 1 9 1 10 9 10 2 13 0 14 13 9 9 9 1 9 0 1 9 10 9 2
35 13 9 10 9 1 9 1 9 0 0 2 16 13 15 15 9 14 13 1 1 10 9 0 1 9 1 9 1 15 14 13 1 9 1 2
22 13 10 9 14 13 1 10 9 9 14 0 7 14 0 10 9 15 1 9 14 9 2
7 2 13 15 15 14 9 2
9 9 14 13 1 10 9 0 10 2
6 13 10 9 0 1 2
21 2 14 13 15 1 9 3 1 3 2 13 9 1 9 1 11 2 10 9 0 2
12 13 10 9 1 9 1 10 9 2 1 9 2
6 9 2 13 8 1 2
16 13 9 10 9 2 9 0 2 1 9 9 0 14 9 1 2
27 13 15 9 10 9 14 0 0 1 9 9 2 9 9 14 9 14 0 2 9 14 9 1 10 9 2 2
27 2 3 1 1 9 0 1 10 9 14 13 1 9 2 7 10 10 9 1 1 9 14 0 1 10 9 2
16 13 11 11 3 1 7 13 1 14 13 9 1 11 14 11 2
13 3 0 1 10 9 1 9 2 13 9 9 1 2
48 1 9 15 13 9 10 9 0 1 9 1 9 1 10 9 2 9 16 14 13 15 1 9 1 9 9 9 1 10 9 1 14 13 10 9 1 2 14 13 1 9 1 9 1 9 0 2 2
12 13 1 15 10 9 14 13 10 9 1 11 2
26 13 1 9 14 12 10 9 14 13 9 7 13 15 10 9 1 9 9 2 1 16 14 13 1 9 2
7 13 0 15 14 9 3 2
18 3 1 3 1 9 0 11 16 1 9 10 9 13 9 1 9 1 2
20 2 13 9 1 2 14 9 2 2 13 11 2 2 14 13 10 9 8 0 2
3 15 9 2
61 16 14 13 0 1 9 14 13 1 10 9 7 13 0 14 13 10 9 14 13 10 9 10 9 1 9 3 2 13 9 9 0 9 14 9 1 9 1 2 11 2 7 13 0 1 11 14 9 1 9 9 1 10 9 0 14 9 1 9 9 2
29 16 13 10 9 1 9 3 1 9 2 13 9 10 9 9 7 13 9 10 9 1 9 9 0 2 10 9 2 2
5 2 15 15 15 2
55 13 15 1 9 1 10 9 2 10 9 1 9 14 14 13 1 10 9 0 2 10 9 1 9 1 10 9 2 10 9 1 9 2 10 9 1 9 2 10 9 0 0 13 1 11 14 13 15 16 14 14 13 15 15 2
4 9 10 9 2
9 14 9 11 7 14 13 15 1 2
37 13 15 0 2 13 0 2 9 1 10 9 14 9 1 9 1 9 10 2 1 9 1 9 2 9 7 14 13 10 9 9 1 9 1 1 9 2
15 11 14 13 15 1 9 1 9 1 9 10 9 1 11 2
16 13 0 14 13 10 9 9 1 2 13 1 9 3 0 10 2
19 13 14 13 1 1 9 1 2 9 0 9 2 9 0 2 9 7 9 2
13 12 13 9 9 1 9 14 13 11 11 1 11 2
30 13 9 1 9 1 9 9 1 9 1 10 9 0 2 14 13 13 0 9 9 9 14 13 3 2 1 9 10 9 2
50 12 1 9 10 12 9 12 2 8 8 12 8 12 2 9 12 2 8 1 9 10 12 9 12 1 9 9 9 14 13 9 1 9 1 9 9 7 1 9 9 3 1 9 2 8 8 12 2 12 2
33 13 10 9 1 10 9 0 3 1 9 1 9 2 1 10 9 2 2 13 15 15 2 13 13 15 9 10 9 15 7 13 15 2
7 13 0 1 9 7 9 2
