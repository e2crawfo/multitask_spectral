4868 11
23 1 9 4 11 13 1 9 1 9 1 9 1 16 9 11 11 13 3 1 10 0 9 2
19 7 3 7 3 0 7 0 1 0 7 0 9 2 15 10 0 13 15 2
12 1 9 7 9 1 9 13 9 7 9 3 2
32 0 10 3 13 9 13 1 9 2 11 11 13 15 12 2 7 9 4 3 0 1 0 9 2 16 15 13 0 9 7 9 2
16 15 4 15 1 0 9 3 0 1 10 0 9 2 11 11 2
26 1 12 4 10 9 13 9 1 11 2 7 15 13 15 3 9 1 2 7 15 13 1 0 7 0 2
7 3 3 1 9 2 13 9
1 13
32 16 9 1 0 9 13 1 9 2 13 15 2 16 10 7 9 9 4 13 0 3 1 2 16 15 4 4 13 1 0 9 2
20 10 0 9 13 1 10 0 9 1 9 1 12 10 0 9 1 9 1 11 2
26 11 11 13 2 16 11 3 4 13 3 1 0 9 2 10 0 9 2 9 7 9 1 10 0 9 2
8 15 15 13 9 1 15 15 2
19 15 4 11 11 2 15 13 1 14 13 9 3 7 13 1 9 1 9 2
22 1 14 4 10 9 1 2 9 2 4 11 11 10 9 1 15 2 15 4 13 9 2
10 1 9 13 9 9 3 1 9 9 2
10 2 15 4 3 3 0 2 13 15 2
11 15 4 13 14 13 9 1 14 13 15 2
34 7 12 9 9 4 9 2 11 11 2 2 3 15 4 13 1 0 9 1 9 2 9 2 9 2 9 2 9 2 9 7 10 9 2
27 2 15 13 2 16 15 4 13 1 10 7 10 0 2 16 15 13 3 7 13 2 16 15 4 13 2 2
13 3 1 11 4 15 13 9 1 12 9 13 9 2
11 2 13 15 3 1 10 9 2 13 15 2
20 3 2 16 9 13 10 0 9 1 10 0 9 2 7 13 1 10 0 9 2
17 15 13 15 1 12 9 7 10 9 4 13 9 1 10 0 9 2
20 14 13 1 9 1 9 4 4 9 2 16 15 3 13 10 0 9 3 1 15
22 9 1 10 9 7 9 1 10 0 12 9 13 2 16 9 13 10 0 9 2 9 2
19 2 15 4 3 3 3 10 0 9 2 16 9 4 4 13 1 13 9 2
29 9 13 14 13 1 9 1 10 9 2 7 9 13 3 0 9 2 16 9 2 15 3 1 9 13 3 2 13 8
23 3 4 15 13 10 0 9 2 15 13 9 2 7 15 4 10 0 9 3 13 15 1 2
33 9 9 1 10 13 0 9 13 3 1 9 9 7 9 2 3 1 9 9 1 15 9 2 15 4 13 1 10 0 9 1 12 2
16 11 9 9 13 3 12 9 3 7 13 1 9 9 1 11 2
23 1 9 13 15 9 1 11 2 7 15 13 15 15 1 10 9 1 10 0 9 1 9 2
3 9 4 3
32 16 3 3 4 13 10 9 1 10 9 2 13 15 3 3 9 2 3 1 15 3 4 3 0 1 9 2 16 9 13 15 2
12 9 4 3 1 12 9 0 7 13 12 9 2
12 2 15 13 2 16 15 3 13 15 3 3 2
17 1 9 1 9 3 13 15 15 1 9 7 13 15 3 1 15 2
15 11 11 11 4 13 12 0 9 1 9 7 9 1 9 2
26 15 13 15 10 2 9 2 9 2 9 2 9 7 9 2 7 15 4 15 3 3 13 3 1 9 2
19 3 13 9 1 10 12 9 2 15 4 13 1 9 1 11 2 13 11 2
5 13 10 0 9 2
14 15 1 9 13 9 1 14 13 2 2 13 11 11 2
6 15 13 13 1 15 2
35 11 0 9 2 1 9 11 11 11 2 11 2 13 9 1 1 9 2 13 9 1 10 0 1 9 1 11 9 3 1 9 10 0 9 2
48 9 1 10 12 9 13 2 13 1 10 0 2 0 9 2 3 1 9 2 9 7 0 9 2 16 11 12 13 10 0 9 1 9 2 15 4 13 3 1 9 1 13 0 12 9 1 9 2
12 7 16 15 13 13 9 2 13 15 1 9 2
31 11 11 4 10 0 0 9 1 0 9 2 7 3 13 9 1 9 1 2 16 3 10 0 9 4 13 10 9 1 3 2
22 7 3 13 0 9 2 7 1 15 13 3 10 9 15 3 4 13 10 0 9 1 2
4 9 13 3 2
15 3 10 0 0 11 2 11 2 4 13 9 7 9 0 2
17 7 13 15 3 7 13 1 10 9 2 13 15 3 3 1 9 2
29 9 1 10 9 4 3 10 9 1 0 9 2 1 10 0 9 1 10 0 9 2 3 15 3 4 13 9 3 2
24 1 14 4 13 3 1 9 7 9 13 15 15 15 1 9 1 14 13 1 10 3 0 9 2
4 9 13 0 2
4 9 1 9 2
3 0 1 11
8 3 3 13 15 1 9 9 2
19 9 13 9 1 10 12 9 0 9 1 9 1 9 2 13 1 12 9 2
4 0 9 1 11
22 15 13 3 2 16 15 13 10 0 9 1 9 1 9 1 10 9 2 2 13 9 2
15 9 13 1 2 16 9 9 3 4 4 13 1 12 9 2
1 9
14 0 9 2 10 0 9 13 1 1 9 1 11 9 2
20 1 11 13 15 10 9 1 14 13 10 9 1 10 0 12 9 13 1 0 2
15 1 9 1 9 13 10 0 9 13 1 9 3 12 9 2
13 10 9 4 10 0 9 1 15 1 10 0 9 2
20 1 10 12 9 1 9 4 2 9 2 3 10 13 7 1 0 9 0 9 2
19 11 9 13 2 16 15 3 4 13 2 16 10 9 3 3 13 1 9 2
24 15 2 15 13 9 2 4 1 3 3 1 10 0 9 2 2 13 15 1 10 0 9 11 2
24 10 10 9 2 11 11 11 11 1 11 9 1 11 12 2 11 2 4 3 13 9 1 9 2
11 9 13 3 1 15 1 0 9 1 9 2
14 15 13 3 9 1 2 16 3 3 3 13 10 9 2
8 7 15 4 3 13 1 15 2
17 1 9 1 10 3 0 9 13 3 0 0 9 1 10 0 9 2
27 9 9 1 0 9 13 1 10 9 1 10 0 9 1 9 1 0 9 2 9 2 11 11 11 11 2 2
10 11 13 2 16 15 4 0 14 13 2
23 3 3 0 9 4 0 1 14 13 1 10 9 15 4 2 15 4 3 3 13 15 3 2
21 10 0 11 12 9 1 9 1 12 9 13 3 9 1 10 9 12 9 0 9 2
35 3 0 4 11 9 13 2 7 1 10 9 1 14 13 13 9 4 11 9 2 0 11 11 1 9 13 1 10 9 1 3 12 9 9 2
28 16 9 1 9 7 9 13 13 1 3 12 7 12 9 2 7 16 9 1 9 8 13 3 12 7 12 9 2
7 3 4 3 13 1 9 2
7 3 13 9 3 3 11 2
29 11 7 11 13 3 3 1 9 10 9 0 9 2 3 15 1 10 3 0 9 4 13 9 9 1 10 0 9 2
18 9 1 9 2 7 10 3 13 9 2 10 12 9 13 1 9 9 2
19 3 4 15 3 9 2 15 13 10 0 9 2 7 15 13 10 0 9 2
12 7 15 4 15 0 1 9 7 13 0 9 2
1 8
9 7 3 4 11 11 3 10 9 2
7 0 9 2 7 9 1 9
22 9 1 9 9 7 0 9 13 10 9 1 9 1 0 9 2 13 9 1 10 9 2
25 9 4 3 13 3 1 14 13 9 3 1 9 2 7 1 0 9 13 9 3 2 7 9 13 2
3 9 1 9
4 9 1 0 9
17 15 13 2 16 15 4 1 9 14 13 11 1 14 13 9 3 2
19 2 7 15 4 15 2 15 13 11 2 13 11 7 13 7 13 1 9 2
6 9 4 4 0 3 2
6 11 13 3 1 9 2
4 3 1 15 2
9 10 0 7 0 13 1 10 9 2
9 2 9 4 1 0 0 7 0 2
32 3 4 15 10 0 9 7 9 2 15 4 13 1 9 1 11 2 2 13 11 3 1 10 9 1 10 0 0 9 1 11 2
10 10 9 13 1 9 12 9 1 9 2
35 4 0 9 3 13 2 3 1 10 9 3 13 1 14 13 2 3 13 10 12 9 1 10 0 2 16 10 0 9 1 1 0 9 13 2
7 11 11 4 11 0 9 2
7 3 13 0 9 1 9 2
32 2 15 4 3 13 2 16 15 1 10 3 0 9 1 0 0 9 13 2 6 2 3 2 2 13 10 0 11 11 1 11 2
13 3 4 10 0 9 2 11 2 13 9 1 9 2
13 7 3 10 9 4 15 10 0 9 1 13 9 2
33 2 3 13 4 15 10 0 9 1 10 9 2 9 4 3 13 1 10 0 9 7 9 2 7 15 15 13 0 9 2 9 2 2
25 15 13 3 1 14 13 1 9 1 9 7 9 2 7 10 9 4 15 3 13 2 14 13 15 2
20 7 3 13 3 3 3 3 0 3 2 16 15 4 13 0 1 10 0 9 2
7 15 13 0 3 1 9 2
11 9 13 0 9 2 3 11 7 11 9 2
18 2 0 13 3 1 9 2 3 1 3 3 3 4 13 9 1 9 2
11 15 13 3 9 1 9 1 10 9 2 2
9 2 9 2 3 15 13 15 2 2
22 3 4 15 0 14 13 10 9 1 3 14 13 15 1 14 13 9 1 9 1 9 2
11 15 4 10 0 9 2 2 13 11 11 2
19 2 15 4 10 0 9 2 15 13 15 2 7 3 13 3 3 15 3 2
40 9 1 10 9 4 12 2 12 2 7 3 1 15 13 2 16 2 10 9 4 3 15 14 13 3 1 2 2 3 4 15 12 3 3 15 2 15 13 1 2
8 10 9 4 3 0 7 0 2
23 10 0 0 9 11 11 13 2 16 15 1 9 9 4 13 9 1 10 9 7 13 9 2
22 9 7 9 13 3 9 1 14 2 13 2 12 9 1 9 2 1 0 10 9 13 2
41 2 15 4 13 1 2 16 9 13 3 0 9 1 11 2 7 15 4 13 9 12 9 2 16 3 4 13 10 13 9 1 9 1 10 0 9 1 0 9 2 2
26 16 15 13 9 1 14 13 15 1 10 0 9 3 1 14 4 13 11 1 10 9 2 15 9 13 2
41 9 13 9 3 1 9 2 3 9 3 4 13 15 1 10 0 9 7 9 1 9 1 11 2 3 9 13 0 9 1 9 10 9 1 9 2 3 15 4 9 2
17 11 11 2 9 2 13 1 9 1 10 9 9 2 9 9 2 2
19 15 4 10 0 9 1 2 3 0 9 2 15 4 13 2 2 13 11 2
30 7 9 1 10 0 2 13 11 1 11 1 10 0 7 0 9 7 11 1 10 0 0 9 13 3 10 9 9 0 2
13 2 3 4 15 4 13 3 3 2 2 13 11 2
17 7 15 4 3 3 0 1 10 0 9 1 0 7 0 9 9 2
18 3 13 12 9 2 1 9 1 9 1 9 0 9 7 1 0 9 2
8 15 13 1 15 1 10 9 2
13 15 4 13 2 16 15 4 13 1 9 1 9 2
28 10 0 9 4 3 13 9 1 14 13 15 1 10 9 1 15 15 0 9 1 0 9 7 0 9 1 9 2
15 10 9 2 15 3 4 13 15 15 2 9 7 9 9 2
20 3 13 15 3 10 9 1 9 13 9 1 3 0 9 2 1 9 1 9 2
26 2 15 13 2 16 16 9 13 3 2 3 4 10 9 3 13 10 9 7 13 3 1 12 9 9 2
29 9 4 0 1 2 16 9 11 11 4 13 1 14 13 9 1 9 7 9 2 16 15 4 9 1 9 1 12 2
18 7 10 0 9 13 9 1 14 4 13 7 13 1 0 1 15 13 2
10 10 9 13 11 11 1 10 0 9 2
12 2 15 4 10 9 2 15 4 13 1 15 2
2 3 2
15 3 4 13 9 1 9 2 7 10 0 9 4 13 3 2
20 11 11 13 2 15 15 3 13 1 11 2 2 9 13 12 1 9 1 9 2
38 15 4 3 3 3 0 1 9 1 9 2 7 1 9 13 9 10 9 1 9 2 15 15 3 4 13 15 1 9 16 15 13 9 1 14 13 3 2
26 9 1 10 9 3 0 1 10 0 9 13 3 1 11 3 1 11 2 11 2 11 2 11 7 11 2
22 2 1 9 4 9 13 15 1 10 0 9 2 7 10 0 13 10 0 9 1 9 2
23 7 16 10 9 13 9 1 14 13 9 7 9 2 4 10 9 1 10 12 9 4 0 2
20 12 9 4 4 13 1 10 0 9 2 7 3 4 4 13 10 9 1 9 2
10 0 9 13 9 3 10 0 9 12 2
18 1 9 4 15 9 13 2 16 9 4 13 10 9 2 15 4 13 2
12 9 1 11 4 3 13 1 14 13 9 3 2
14 2 15 4 9 2 15 3 13 15 2 2 13 11 2
12 2 2 6 2 15 4 11 2 15 13 15 2
26 11 9 2 11 11 2 13 1 9 10 9 1 11 1 14 13 9 1 11 2 7 1 10 0 9 2
56 1 9 9 4 15 13 10 10 7 3 3 0 13 9 2 3 10 0 2 16 1 10 0 9 2 1 15 13 15 3 1 2 4 3 3 3 10 13 9 13 1 9 2 16 9 3 13 9 3 2 13 15 0 7 0 2
12 10 9 2 3 1 0 2 7 1 0 9 2
26 15 13 9 1 10 9 1 3 14 13 10 0 9 1 9 2 16 3 4 13 10 9 1 11 9 2
33 2 9 2 13 9 1 11 11 2 9 1 0 9 1 11 7 9 1 11 9 2 15 4 13 1 12 9 7 1 9 12 9 2
24 10 9 4 0 2 15 4 13 9 1 11 7 3 11 9 1 14 13 13 9 7 3 9 2
10 9 4 3 13 9 1 10 10 9 2
13 3 13 15 14 13 3 2 14 13 10 9 2 2
10 9 4 0 7 0 7 0 1 9 2
10 3 13 3 9 7 13 9 1 9 2
13 11 11 9 2 9 1 9 2 4 10 0 9 2
9 7 15 4 9 1 0 10 9 2
10 1 11 4 9 9 10 9 1 9 2
23 11 11 13 1 11 11 2 11 11 2 11 11 2 11 11 7 10 0 2 13 11 11 2
13 3 4 10 12 0 9 1 9 1 10 0 9 2
15 9 13 9 7 9 2 1 9 3 4 7 13 13 1 2
17 3 3 10 0 9 3 4 4 13 3 2 2 13 11 11 11 2
10 2 15 13 3 1 9 2 13 11 2
20 2 15 4 3 3 13 2 16 3 4 13 10 9 2 3 16 9 4 3 2
35 15 4 9 2 9 9 2 2 11 11 2 15 13 15 9 2 16 15 13 10 9 2 10 0 9 2 3 13 9 7 9 1 0 9 2
39 15 13 3 1 9 2 7 13 10 9 3 2 16 15 13 10 0 9 3 1 15 2 7 13 10 9 1 15 2 1 14 13 15 15 4 13 15 1 2
3 3 5 12
20 15 4 3 3 9 2 16 15 4 13 3 1 9 2 15 15 13 1 9 2
10 4 15 13 2 4 15 13 1 9 2
21 15 4 3 13 1 9 1 9 1 11 9 7 4 3 13 0 1 11 7 11 2
19 3 13 15 1 9 1 10 0 9 1 2 16 15 4 13 1 10 9 2
11 2 10 9 4 15 3 13 1 9 1 2
16 3 4 15 3 13 15 13 1 14 13 15 2 1 12 9 2
8 7 15 13 3 3 3 2 2
6 3 4 13 12 9 2
22 15 4 3 13 9 0 1 9 1 9 7 9 2 11 12 2 11 11 3 0 9 2
10 7 3 13 9 3 1 14 13 15 2
7 11 13 9 3 1 9 2
20 3 4 15 3 3 16 9 4 13 12 9 7 13 3 0 9 7 8 9 2
24 15 13 2 16 9 4 4 0 1 14 13 1 9 2 7 3 4 9 13 3 13 7 0 2
10 15 4 3 13 14 13 3 1 15 2
32 0 9 3 1 10 0 9 1 9 13 3 1 9 2 15 13 3 1 11 2 1 0 9 2 7 0 9 4 10 9 3 2
18 0 4 15 3 14 13 10 9 1 10 0 9 2 15 4 13 9 2
7 11 11 9 11 9 9 2
19 3 9 7 9 4 3 13 1 9 2 15 3 13 9 7 10 0 9 2
31 15 4 13 10 9 1 0 10 9 2 15 3 13 9 14 13 10 9 2 7 15 13 3 15 2 7 15 13 15 0 2
14 3 4 10 0 9 13 3 2 16 15 4 3 13 2
13 13 2 9 4 3 3 13 15 14 13 0 9 2
26 9 13 1 0 0 9 2 7 10 9 13 15 3 0 1 15 2 16 15 3 4 13 15 1 9 2
9 10 7 0 15 9 13 13 9 9
13 10 9 2 15 3 4 13 2 4 0 1 9 2
48 15 4 0 1 9 7 9 1 3 14 13 7 13 1 14 13 10 0 9 1 10 0 9 7 13 10 9 1 10 0 9 2 7 13 0 9 1 15 15 1 9 2 16 15 3 13 9 2
14 16 15 13 3 1 15 2 4 15 3 10 0 9 2
31 3 1 9 4 13 2 13 3 3 9 1 10 0 9 2 16 11 11 11 3 13 2 16 15 4 13 15 10 0 9 2
7 9 13 3 1 0 9 2
15 10 0 9 13 2 16 9 8 8 13 9 7 9 9 2
1 9
9 3 9 9 9 4 13 10 9 2
3 9 1 9
16 10 9 2 15 4 13 1 9 2 4 3 4 3 3 0 2
18 7 16 15 13 3 2 4 3 3 13 9 1 0 9 1 10 9 2
16 10 0 0 9 2 1 15 3 4 4 0 3 14 13 1 2
5 11 13 10 9 2
11 9 1 10 12 9 13 1 10 0 9 2
4 10 0 9 13
53 2 15 4 13 2 16 15 15 4 13 1 10 0 9 7 3 15 12 4 13 3 3 2 16 15 4 13 1 2 16 10 3 0 4 13 9 2 2 13 11 11 2 15 3 13 0 1 10 3 3 0 9 2
17 4 15 13 2 16 15 13 16 9 4 0 2 4 15 13 15 2
18 10 0 0 9 1 10 9 2 15 4 13 15 1 9 2 4 9 2
4 11 4 0 2
7 11 13 9 7 13 3 2
8 7 11 11 4 10 0 9 2
15 15 4 9 1 0 9 11 11 2 9 2 9 7 9 2
30 1 10 9 13 9 1 9 10 9 1 9 7 9 2 1 15 10 9 1 9 2 1 9 13 10 9 1 1 9 2
8 15 4 0 2 1 15 13 2
4 13 15 13 15
34 2 15 4 10 0 9 2 3 10 0 9 4 13 3 1 9 9 2 9 2 1 9 7 1 9 2 2 13 9 11 11 2 11 2
6 13 1 9 1 9 2
29 3 13 11 3 1 9 2 16 3 13 12 9 2 7 1 9 4 11 1 12 9 1 9 13 10 9 1 12 2
15 2 15 4 3 13 0 2 15 15 4 13 2 1 9 2
11 2 10 9 2 10 9 2 4 13 3 2
18 10 0 9 13 9 1 11 7 11 1 2 16 0 9 4 4 13 2
26 3 0 15 3 4 13 2 4 0 14 13 2 16 15 3 13 2 3 10 0 4 4 13 1 9 2
11 15 13 2 16 9 1 3 13 1 9 2
23 10 0 9 13 2 16 12 9 4 4 0 2 7 16 12 1 15 4 4 13 1 9 2
20 16 15 13 1 10 9 9 4 13 2 3 4 15 3 13 3 1 8 11 2
13 15 13 10 9 7 10 9 2 15 3 3 13 2
30 10 12 13 9 1 0 9 9 2 9 11 11 11 7 9 11 11 2 13 1 9 9 1 11 9 1 9 1 9 2
5 9 16 15 4 13
25 10 0 9 4 3 4 13 1 9 1 12 2 3 0 9 13 14 4 15 1 9 2 13 11 2
26 15 13 15 3 3 13 7 13 15 1 2 3 15 3 3 4 15 2 15 4 13 2 2 13 15 2
8 11 13 7 13 14 13 15 2
10 3 4 9 3 2 2 13 11 11 2
24 15 13 3 12 9 3 1 15 2 13 3 0 7 4 3 1 9 1 9 13 15 12 5 2
16 9 9 11 2 9 1 0 9 2 13 3 1 9 7 9 2
21 15 4 4 13 3 1 9 2 3 1 10 2 9 2 2 15 4 4 13 3 2
2 0 9
23 11 11 9 2 9 11 11 2 15 1 9 13 12 9 2 4 10 0 9 1 0 9 2
3 9 1 9
3 9 7 9
16 3 4 15 3 4 13 0 9 2 7 15 4 3 3 0 2
4 10 9 1 11
5 9 13 1 9 2
13 11 0 9 11 11 4 3 3 13 3 1 15 2
7 7 15 4 10 0 9 2
31 8 8 10 0 9 13 9 4 9 7 10 0 0 9 13 0 9 1 9 2 16 15 13 2 10 0 2 0 9 2 2
20 7 15 4 3 3 13 15 7 13 1 2 15 11 13 2 16 15 4 0 2
19 12 9 1 11 13 1 2 16 10 0 9 1 12 9 3 13 3 1 9
20 3 13 3 3 3 0 9 1 10 0 9 1 10 9 1 12 3 7 3 2
8 13 9 7 9 3 1 3 2
7 15 1 9 4 0 3 2
35 11 2 9 1 12 9 0 11 2 11 11 7 11 11 2 11 1 11 2 4 13 1 2 16 10 9 13 10 10 9 1 10 0 9 2
39 15 3 13 10 9 4 3 4 9 2 9 4 3 13 10 3 0 9 1 10 9 15 9 13 3 2 7 4 3 13 3 1 15 15 4 13 3 1 2
8 7 15 13 11 3 9 1 2
11 3 13 3 3 9 1 10 3 0 9 2
6 15 13 1 9 2 2
32 2 15 13 1 10 9 10 9 2 1 15 4 13 3 1 1 12 9 2 7 10 9 13 1 9 2 16 15 13 1 9 2
16 1 10 13 9 4 15 4 0 14 13 9 1 10 0 9 2
13 13 9 1 10 9 1 2 15 3 13 9 9 2
15 1 9 1 9 13 11 11 15 13 1 1 9 12 9 2
13 3 7 3 13 7 13 10 0 9 1 10 9 2
10 9 4 4 10 0 2 13 15 15 2
2 10 0
26 16 3 13 3 3 9 1 10 9 1 10 0 9 2 2 13 9 11 11 1 9 7 9 1 11 2
22 11 13 3 14 13 10 9 13 1 9 2 7 0 9 13 1 9 9 1 10 9 2
20 16 2 11 2 13 3 1 9 9 2 4 15 13 3 1 10 3 0 9 2
9 2 9 4 13 10 9 1 9 2
5 15 4 3 13 2
27 9 13 2 3 3 13 3 2 7 16 9 13 9 1 9 1 9 2 4 15 13 15 1 14 13 9 2
8 15 13 3 10 0 9 2 2
16 15 15 13 2 2 3 12 9 1 9 9 13 15 10 9 2
6 3 13 15 3 1 9
9 9 1 9 4 10 3 10 9 2
24 10 0 9 1 11 9 1 11 2 11 11 11 2 13 2 9 1 9 13 0 1 9 9 2
9 3 13 15 3 9 1 11 9 2
22 15 13 1 14 13 12 9 0 9 1 10 0 9 2 2 13 11 9 2 11 11 2
15 10 9 4 13 9 11 13 10 0 9 1 9 1 9 2
35 11 11 2 11 11 2 2 11 11 2 11 11 2 2 11 11 2 11 11 2 2 11 11 2 11 11 2 2 11 11 2 11 11 2 2
19 2 9 13 3 14 13 3 1 2 15 4 10 0 9 1 9 1 13 2
11 15 13 3 0 14 13 11 7 11 1 2
45 0 1 10 3 0 9 2 15 3 3 4 13 3 2 4 9 9 2 8 2 15 1 12 4 13 1 11 7 3 7 3 3 4 3 1 11 1 9 1 11 2 11 13 9 2
50 15 13 1 11 2 15 4 13 10 0 9 3 1 10 0 9 1 10 0 9 2 1 9 2 15 1 13 9 2 10 0 9 1 9 1 9 7 15 15 3 13 3 1 9 2 3 13 1 9 2
28 1 10 9 1 3 12 9 13 10 0 8 11 11 1 12 1 10 9 1 10 9 2 2 9 1 9 2 2
37 10 9 4 1 9 4 3 1 14 13 10 0 9 2 15 13 1 15 1 9 2 3 15 1 10 9 1 15 2 15 13 1 9 13 3 13 2
14 9 4 10 0 9 2 15 13 3 0 9 1 9 2
20 9 1 9 4 3 13 2 7 3 3 2 1 12 9 9 1 12 9 9 2
17 3 13 0 9 15 13 9 1 9 2 3 9 3 13 1 9 2
26 15 4 1 12 9 1 9 13 1 10 9 1 11 1 11 1 9 2 11 2 2 15 13 1 9 2
46 10 0 9 4 13 3 1 10 0 9 2 7 1 9 2 15 4 13 2 16 9 4 10 0 9 2 13 3 9 1 9 14 13 1 10 9 2 3 10 12 9 13 3 1 15 2
23 9 3 12 9 1 9 1 9 1 11 13 12 9 1 10 0 1 9 1 9 7 9 2
6 13 10 0 9 14 13
13 11 2 3 9 13 1 2 13 3 2 9 2 2
10 9 11 11 4 3 4 13 9 3 2
9 15 4 10 9 2 15 13 9 2
6 3 4 0 15 13 2
35 10 12 9 3 0 9 13 1 9 0 9 1 9 2 11 2 1 12 2 13 0 9 1 14 13 15 2 3 1 15 3 4 13 9 2
14 7 3 3 10 0 9 13 2 15 15 4 13 3 2
3 2 6 2
24 15 13 10 0 9 13 15 2 16 2 11 4 0 11 9 2 16 15 13 9 7 9 2 2
5 3 3 7 3 2
16 15 4 12 9 2 7 15 4 0 14 13 9 1 10 9 2
6 15 4 3 0 9 2
6 13 9 3 1 9 2
7 3 13 10 3 13 9 2
25 10 9 2 3 4 3 0 2 16 15 13 10 9 7 3 4 13 10 9 1 14 13 10 0 2
15 15 13 10 0 9 1 10 9 2 15 4 15 3 13 2
10 1 11 11 7 1 11 7 11 11 2
24 15 4 4 3 0 1 2 16 9 13 1 2 16 9 4 13 15 2 2 13 9 11 11 2
5 15 4 15 3 2
8 10 9 2 15 13 15 0 2
10 10 9 4 13 10 0 9 1 15 2
17 2 15 4 3 3 10 0 2 15 13 9 7 9 2 13 15 2
31 15 4 0 1 12 9 3 2 16 9 13 9 1 14 13 10 0 9 1 11 7 1 9 13 0 9 9 1 10 9 2
3 2 12 2
1 9
24 11 11 11 13 1 11 11 0 9 12 2 3 11 11 11 13 1 0 2 9 2 1 9 2
13 11 13 10 0 9 14 13 1 2 16 15 13 2
18 15 13 1 14 13 14 13 2 16 15 4 13 1 14 13 11 3 2
23 1 11 4 9 3 0 2 16 9 1 10 0 9 11 4 13 3 3 1 10 0 11 2
13 9 1 9 1 10 0 9 13 3 14 13 11 2
14 10 9 1 12 13 7 10 0 9 1 12 9 9 2
9 9 4 3 3 3 13 9 1 2
37 3 3 1 9 2 7 0 9 1 9 2 9 7 9 2 16 9 3 13 1 14 13 3 7 4 13 10 9 9 1 9 1 9 7 1 9 2
6 9 13 3 3 13 2
12 7 9 4 3 0 1 14 13 9 1 9 2
19 3 13 15 9 1 14 13 3 1 10 0 9 2 15 3 4 0 15 2
42 3 13 1 10 0 9 2 15 1 9 13 15 1 9 0 9 2 15 15 13 1 9 2 10 0 9 2 15 3 9 0 13 15 15 3 1 9 1 0 7 0 2
15 10 9 2 15 13 3 1 9 13 10 0 7 0 9 2
29 15 13 1 9 1 10 0 2 15 3 13 2 16 9 13 9 9 2 7 13 3 1 3 14 13 15 1 9 2
5 9 4 9 9 2
9 2 7 3 13 10 9 1 0 2
18 3 11 7 11 13 1 9 2 7 10 0 9 11 13 1 9 3 2
11 13 3 16 15 13 2 13 7 3 13 2
29 9 13 14 13 9 3 2 3 4 15 3 13 0 2 7 3 13 3 9 1 9 2 2 13 9 11 11 11 2
11 3 13 15 1 10 12 9 0 13 9 2
14 15 4 13 2 16 0 9 1 9 13 15 1 15 2
1 9
13 1 1 9 9 13 9 14 13 3 1 10 0 2
16 7 15 4 3 13 1 14 13 3 0 9 14 13 9 0 2
13 9 4 13 1 15 1 9 1 9 1 10 9 2
20 3 13 9 1 2 9 2 3 1 2 16 9 13 9 1 9 1 9 12 2
13 2 12 9 9 2 13 11 7 13 3 1 9 2
6 3 9 4 13 15 2
22 3 13 13 9 0 9 3 1 10 0 9 1 2 9 2 1 11 11 9 1 11 2
34 3 1 10 0 13 15 9 1 9 1 2 16 10 9 4 13 0 2 10 9 1 10 0 9 4 13 2 16 15 4 13 10 9 2
15 11 11 2 9 2 4 4 0 9 1 11 9 1 11 2
14 9 2 15 13 9 1 10 9 2 13 2 9 2 2
24 9 2 15 3 13 9 2 9 7 0 9 2 4 13 3 2 7 15 4 3 13 15 3 2
23 1 10 9 1 9 4 11 3 13 10 13 9 1 10 9 2 15 9 7 9 4 13 2
19 1 9 13 12 9 1 9 1 11 2 7 3 13 10 0 9 1 9 2
22 10 2 13 2 9 13 1 11 2 11 7 11 2 7 9 4 3 13 1 10 9 2
5 15 4 3 13 2
28 2 15 13 0 2 16 9 4 3 2 2 13 9 9 15 2 16 15 3 13 2 16 15 13 9 3 3 2
7 1 9 1 9 4 9 2
12 1 9 13 15 1 9 1 12 9 1 9 2
12 2 9 0 1 0 2 3 0 1 9 7 9
34 15 4 13 0 9 1 9 2 7 9 4 1 0 9 4 10 9 2 15 13 0 7 0 3 2 7 9 4 3 0 14 13 3 2
13 3 13 9 1 3 9 1 9 15 1 10 0 2
10 11 11 4 3 13 9 1 0 9 2
8 15 4 3 13 14 13 15 2
19 9 13 0 9 9 1 9 1 9 1 9 2 10 0 9 7 10 9 2
16 16 15 13 1 11 9 2 4 15 10 0 9 1 10 9 2
3 13 12 9
33 15 13 9 12 1 10 9 2 13 9 2 13 9 7 9 2 13 9 1 9 7 4 3 1 14 13 10 9 2 15 4 13 2
9 7 15 15 13 1 10 0 0 2
1 9
24 9 1 9 13 3 3 11 11 1 14 13 2 16 15 3 4 13 10 3 0 1 15 3 2
22 11 11 4 13 10 0 11 2 15 3 4 1 9 1 14 13 9 0 9 1 9 2
15 2 9 1 12 9 2 13 2 15 9 13 2 9 9 2
9 15 4 3 13 9 12 9 9 2
14 9 13 1 11 2 10 0 9 1 0 2 0 9 2
3 0 9 2
14 7 1 10 9 13 15 0 9 1 14 13 10 9 2
18 16 10 0 9 4 13 13 9 1 9 4 3 0 1 9 1 11 2
3 9 13 2
13 12 9 4 13 1 10 0 0 9 1 9 9 2
4 12 9 1 9
15 3 4 9 4 0 14 13 7 13 1 3 1 0 9 2
2 9 2
26 10 12 9 2 10 1 15 9 2 13 10 9 1 9 1 10 0 9 2 1 9 1 9 1 11 2
33 3 1 9 4 3 13 10 9 1 11 7 11 1 9 1 10 0 9 2 7 11 4 3 13 11 1 9 1 10 9 1 9 2
22 15 4 3 13 3 3 2 7 3 13 3 9 1 14 13 15 2 7 9 13 13 2
1 8
27 3 3 9 11 11 9 13 0 9 1 2 16 3 1 9 9 9 3 13 10 0 0 9 2 4 13 2
1 9
5 2 15 3 3 2
12 15 13 3 1 10 9 1 0 1 12 9 2
9 3 13 10 9 1 9 7 9 2
11 1 9 13 11 9 9 7 0 0 9 2
37 1 9 7 10 13 12 9 13 11 11 11 9 0 1 11 9 12 2 7 3 4 15 9 1 10 0 0 9 2 11 9 2 3 1 9 2 2
16 1 9 13 10 0 9 1 10 9 1 9 1 14 13 9 2
14 11 13 3 7 13 2 16 15 3 4 13 3 3 2
10 16 3 3 4 10 9 3 1 15 2
41 4 15 13 1 9 2 7 15 13 15 3 2 6 3 4 15 3 16 2 15 13 15 13 1 2 16 15 4 0 1 14 13 1 9 1 11 1 10 0 9 2
17 1 9 13 12 0 9 1 9 11 7 12 0 0 0 1 9 2
9 11 11 11 2 11 12 2 12 11
15 0 9 4 3 13 9 1 14 13 0 9 1 9 9 2
15 10 0 9 13 3 3 1 10 0 9 1 9 0 9 2
24 9 13 1 10 9 3 1 2 16 15 3 1 9 4 13 2 1 15 9 9 4 13 2 2
5 2 15 13 9 2
16 15 4 3 13 10 0 9 1 9 1 9 7 4 4 9 2
15 7 3 4 13 9 1 9 2 15 3 13 10 0 9 2
35 2 16 3 13 10 0 0 9 1 3 14 13 0 7 14 13 9 1 9 2 3 4 10 9 1 9 1 11 11 4 10 0 9 2 2
23 9 2 11 11 2 4 13 9 1 9 1 14 13 0 1 13 9 1 9 7 1 9 2
38 15 4 9 1 9 1 15 13 2 15 4 13 3 0 2 16 10 0 3 15 4 13 9 1 9 7 9 1 14 13 9 2 3 1 3 0 9 2
22 15 13 2 16 15 4 0 1 15 7 13 0 9 9 1 9 2 2 13 11 11 2
16 9 7 9 1 11 13 1 9 1 11 1 9 9 7 9 2
13 2 15 13 3 1 2 16 15 4 13 9 3 2
1 9
6 2 15 13 1 15 2
20 15 4 3 0 4 0 13 13 9 2 9 2 1 10 9 0 9 7 9 2
17 0 9 13 3 3 3 3 1 11 13 9 2 9 11 1 11 2
18 7 16 15 13 3 1 2 11 7 11 13 1 14 13 9 1 15 2
5 2 0 2 3 2
11 15 0 9 1 10 9 13 1 10 9 2
11 3 4 11 0 1 2 16 11 13 9 2
16 15 13 2 15 13 9 10 0 0 9 2 16 15 13 3 2
39 9 1 9 4 11 4 13 1 9 1 9 2 15 1 10 13 9 13 2 16 3 4 15 3 13 9 3 3 1 14 13 3 2 16 9 13 1 9 2
12 13 0 9 9 2 11 11 2 1 11 11 2
9 2 13 15 3 2 2 13 9 2
35 11 11 2 0 9 1 13 1 0 9 13 1 11 11 1 12 9 3 2 4 13 0 9 3 3 1 10 0 9 1 10 9 11 11 2
35 11 9 4 10 0 7 13 9 2 15 4 13 1 0 9 2 7 1 3 4 13 15 14 4 3 0 1 9 7 1 9 1 0 9 2
8 9 7 15 15 3 13 2 2
13 15 13 3 2 10 9 4 13 1 0 0 9 2
5 9 13 0 10 9
7 13 15 3 13 1 15 2
27 7 15 4 13 1 9 2 7 15 4 3 13 2 3 0 15 3 13 2 16 9 13 1 10 0 9 2
12 15 4 13 1 9 3 2 3 3 15 13 2
22 2 15 13 2 3 1 15 3 4 9 2 15 13 15 1 9 1 2 2 13 15 2
16 3 4 15 13 2 3 15 13 3 2 16 9 13 15 3 2
15 9 4 13 1 12 9 7 12 9 1 9 7 9 1 8
22 13 15 13 15 14 13 10 0 9 2 15 3 13 2 13 15 3 1 9 1 9 2
17 0 0 9 13 12 9 1 9 7 12 9 9 12 9 12 9 2
26 9 1 9 2 12 9 1 0 9 2 15 13 3 1 9 2 4 3 13 1 10 9 12 9 3 2
11 0 4 13 2 3 10 13 9 13 15 2
20 15 4 13 10 0 0 0 9 2 15 4 10 0 9 1 10 9 1 12 2
27 3 6 1 2 16 0 11 13 11 9 1 10 9 1 10 9 2 15 4 13 2 16 10 9 4 0 2
20 9 9 13 1 10 0 9 1 14 13 0 9 7 13 0 9 1 9 9 2
3 13 10 9
7 13 9 5 12 9 5 11
19 10 10 0 9 2 11 2 13 1 9 10 0 9 1 9 0 9 12 2
19 0 1 9 7 13 1 14 13 3 7 13 9 2 15 15 13 9 1 2
9 0 9 4 3 3 0 1 9 2
13 9 4 2 3 3 9 12 13 9 1 0 9 2
2 3 2
15 0 9 4 3 13 0 9 2 16 15 3 13 1 9 2
8 2 3 13 15 1 15 15 2
15 15 13 3 1 10 9 2 16 15 13 9 1 10 9 2
12 3 13 15 3 1 9 2 7 3 13 15 2
26 9 2 15 3 13 1 9 1 9 1 9 2 13 15 9 1 2 7 15 13 3 9 3 1 9 2
7 7 11 9 13 3 13 2
19 9 13 10 9 3 1 9 2 3 15 13 9 1 14 13 9 9 3 2
2 0 9
32 15 13 3 1 10 0 9 7 13 1 10 12 9 0 9 2 3 3 4 13 10 9 2 1 1 9 4 4 11 0 9 2
33 3 1 12 13 9 11 9 1 9 2 7 1 9 0 9 13 11 3 1 12 9 2 10 0 4 11 11 2 10 0 9 9 2
20 11 13 3 1 9 1 15 1 10 0 9 1 9 7 15 15 1 10 9 2
26 16 15 13 9 3 1 9 2 13 15 10 9 1 9 1 10 9 1 0 9 1 1 10 0 9 2
5 9 13 1 9 2
7 0 2 0 2 0 9 2
8 3 13 15 1 9 1 9 2
7 15 13 0 9 1 9 2
9 9 4 13 1 9 16 9 13 2
26 10 10 0 9 4 13 1 9 1 10 0 9 2 16 10 0 9 4 13 9 13 1 9 1 9 2
6 9 2 9 1 8 2
19 9 1 9 13 2 16 9 3 4 13 9 1 9 1 9 1 9 9 2
54 2 1 14 13 0 0 9 7 3 9 1 10 0 9 2 13 15 15 3 2 3 1 10 9 2 1 14 13 1 11 2 3 16 15 13 3 2 3 16 15 13 2 16 15 13 15 2 15 13 9 1 9 2 2
12 2 3 3 15 4 13 3 2 13 15 3 2
13 13 12 9 9 7 9 3 3 1 10 0 9 2
34 15 4 3 13 0 9 2 16 15 4 13 9 7 9 3 1 9 1 10 3 0 7 0 9 2 1 15 4 13 15 3 1 9 2
8 2 3 4 15 13 10 9 2
29 3 13 0 9 1 10 13 9 9 2 7 3 9 13 3 2 15 10 9 13 1 9 2 16 9 4 13 3 2
5 2 3 3 3 2
10 15 9 13 3 3 3 0 3 3 2
5 12 2 12 9 2
2 10 9
6 15 4 15 3 13 2
35 3 1 9 1 14 4 13 1 14 13 8 7 0 13 15 15 1 10 9 2 15 4 8 2 9 3 4 13 1 2 2 13 11 11 2
8 0 9 1 12 9 4 13 2
19 10 0 9 4 15 13 10 0 9 1 10 12 10 0 9 9 1 11 2
11 16 15 13 9 7 9 4 3 10 9 2
10 9 1 10 0 9 2 11 11 2 11
2 9 12
9 9 4 9 7 10 12 9 9 2
8 15 4 0 12 0 9 3 2
24 9 3 13 15 1 10 3 0 9 2 15 13 10 10 9 14 4 3 1 2 1 15 13 2
17 3 4 15 3 13 15 3 2 16 15 3 4 13 3 1 9 2
10 11 11 4 9 7 4 3 13 3 2
14 2 13 15 3 2 11 2 6 3 13 3 3 3 2
35 3 4 15 13 3 0 9 1 10 9 1 9 1 11 2 3 3 13 3 3 0 9 1 1 11 2 7 3 3 9 1 15 4 9 2
15 15 4 3 0 2 13 3 9 3 7 13 10 9 2 2
7 3 9 4 13 10 9 2
34 2 15 13 15 3 3 13 2 7 10 0 9 4 13 10 9 2 16 0 9 3 4 4 3 3 0 1 14 13 1 0 9 2 2
27 1 11 9 1 11 13 15 3 14 13 9 1 13 9 1 14 13 9 1 14 13 15 3 1 0 9 2
10 7 15 13 15 2 7 15 13 15 2
2 9 12
23 9 13 2 7 15 4 9 9 2 15 13 9 1 10 0 9 7 10 0 9 1 9 2
21 1 9 1 9 1 9 13 3 10 9 0 9 2 15 3 4 13 1 12 9 2
32 9 13 1 10 0 0 9 1 11 2 7 3 13 15 1 10 0 2 15 13 3 3 2 2 13 11 11 2 11 1 11 2
14 10 0 13 9 2 15 13 1 9 2 13 11 0 2
28 15 13 11 1 9 0 9 1 9 2 7 3 13 3 10 9 1 10 9 2 15 13 1 10 13 9 11 2
1 9
16 16 15 13 10 9 2 13 15 3 3 15 1 1 0 9 2
5 3 10 9 1 9
3 0 11 2
25 7 15 13 2 16 15 1 0 9 1 9 13 2 4 10 9 13 1 10 9 1 10 0 9 2
7 7 15 13 3 10 9 2
20 15 1 9 1 9 4 13 2 16 15 3 13 9 1 14 13 9 1 9 2
22 3 13 3 11 1 9 11 7 11 14 13 10 3 0 9 2 1 9 9 4 13 2
13 1 10 0 9 4 15 3 3 13 10 13 9 2
14 1 0 9 0 9 14 4 2 13 15 15 3 3 2
24 3 4 15 1 10 9 4 10 9 1 9 2 16 9 3 13 3 1 14 13 1 9 2 2
25 15 4 10 9 1 9 7 9 2 9 11 11 13 2 16 15 1 9 9 13 1 9 0 9 2
13 9 1 9 4 3 13 10 0 9 1 9 9 2
29 2 9 4 10 0 9 2 3 9 4 13 9 1 9 2 2 13 11 11 2 15 13 1 11 1 11 1 9 2
8 15 4 1 12 7 1 12 2
22 1 9 13 15 1 14 13 10 9 1 11 2 13 1 0 9 1 11 9 1 11 2
4 3 0 0 9
16 11 3 0 9 13 15 3 3 1 9 0 9 10 0 9 2
27 16 9 4 10 9 2 3 15 13 14 13 15 0 2 2 13 11 11 1 15 11 11 11 13 0 9 2
5 11 11 2 0 2
19 11 11 13 1 12 9 3 1 11 9 2 3 15 13 10 9 11 11 2
15 15 4 0 1 10 0 2 16 0 8 4 10 0 9 2
16 3 13 15 10 9 1 14 13 9 2 7 15 13 9 3 2
14 2 13 9 11 11 1 15 2 13 15 1 13 9 2
7 9 5 2 3 3 13 2
21 7 15 13 10 0 0 9 1 2 15 13 9 1 9 1 11 1 9 1 9 2
26 2 15 4 3 0 2 16 15 3 13 1 14 13 2 2 13 10 9 1 12 2 15 13 1 9 2
5 9 2 12 8 2
13 15 4 15 3 13 2 7 15 4 3 13 9 2
11 15 13 15 13 2 16 15 4 10 9 2
7 13 3 1 9 1 9 2
5 3 13 15 9 2
22 1 9 13 11 11 7 9 11 11 2 16 9 13 10 1 3 9 1 9 1 9 2
3 9 1 9
25 9 4 3 2 7 1 3 13 15 2 7 15 4 13 7 13 2 15 11 11 13 15 3 3 2
44 16 3 1 15 3 4 11 11 2 15 13 9 9 7 9 3 1 10 9 2 4 15 3 15 1 10 9 2 3 9 13 3 1 9 1 10 13 2 0 9 1 9 3 2
7 3 4 15 3 13 9 2
2 3 0
19 2 15 4 10 0 0 9 2 1 9 10 9 4 1 2 2 13 11 2
9 7 15 4 3 7 3 1 9 2
8 7 15 4 3 13 10 9 2
31 13 4 15 3 3 2 16 9 1 13 0 9 1 0 0 9 2 4 13 9 3 0 9 2 1 9 3 3 13 15 2
8 15 4 3 13 8 8 8 2
2 0 9
1 9
25 15 13 0 9 15 9 1 9 12 2 3 0 9 4 0 1 14 13 2 15 3 13 1 15 2
27 9 9 4 3 13 9 1 9 3 2 7 3 1 9 2 15 4 13 1 9 2 4 3 13 7 13 2
50 3 13 11 11 3 9 1 14 13 1 9 2 16 15 3 1 16 2 3 1 9 2 13 10 0 9 1 2 13 3 2 16 15 4 13 7 0 1 11 7 3 1 12 1 3 4 13 12 9 2
8 15 4 15 3 13 9 1 2
29 15 4 0 9 2 7 3 9 4 3 13 1 9 7 9 1 9 4 10 3 13 9 1 3 2 11 3 2 2
10 1 9 4 3 11 11 11 9 0 2
26 11 11 4 3 4 9 1 9 7 9 11 2 7 4 1 10 9 1 12 9 1 0 9 1 9 2
26 15 4 13 1 10 0 9 7 13 1 0 9 2 16 15 4 13 9 3 1 11 11 7 10 9 2
23 13 1 15 13 15 3 1 10 9 2 16 15 4 0 2 7 16 15 13 10 9 2 2
6 2 13 15 1 15 2
4 2 0 2 13
7 15 4 13 9 3 13 2
11 2 3 13 11 2 2 13 11 1 15 2
24 10 13 9 13 3 14 13 9 13 1 10 9 1 9 7 13 3 1 10 0 2 0 9 2
19 15 4 3 3 13 15 16 15 4 13 10 9 1 9 7 1 0 9 2
22 3 1 10 9 1 9 13 15 14 13 3 9 7 9 7 14 13 9 1 0 9 2
40 15 4 4 13 12 9 1 10 9 9 2 7 1 10 9 9 7 9 2 3 3 1 10 9 13 0 9 1 9 2 13 9 1 9 1 0 9 1 9 2
11 15 4 15 3 13 3 1 3 1 9 2
13 2 15 4 4 13 10 10 9 2 13 11 3 2
15 15 4 10 0 0 9 0 9 2 15 13 9 1 9 2
12 1 11 11 9 13 10 0 9 1 0 9 2
14 0 9 4 13 9 1 9 2 0 9 4 13 9 2
12 15 13 7 15 4 0 2 7 10 0 9 2
9 13 15 9 2 2 13 9 11 2
24 10 10 9 4 3 3 3 3 13 2 15 13 3 1 9 2 0 2 7 13 1 12 9 2
11 9 4 3 4 0 2 7 0 7 0 2
17 7 9 4 13 2 16 11 3 13 3 1 10 0 9 1 9 2
11 9 13 3 1 2 13 3 1 9 2 2
25 9 1 12 9 7 3 1 9 4 9 1 11 7 11 2 9 8 2 9 1 11 7 0 9 2
16 15 13 10 9 13 9 2 16 15 13 10 9 1 10 9 2
9 15 13 15 3 3 7 13 15 2
17 15 13 10 9 1 9 1 11 2 7 15 13 3 3 2 6 2
18 9 2 1 15 13 9 11 11 2 13 12 9 1 9 1 11 11 2
8 2 1 9 1 10 0 9 2
13 3 13 15 9 2 1 15 13 3 1 1 9 2
11 9 7 9 13 3 12 9 1 9 9 2
36 3 4 3 3 3 13 0 9 7 0 9 1 10 0 0 9 2 11 11 12 9 9 2 15 4 4 13 1 10 0 9 1 9 1 11 2
32 16 11 11 1 3 0 9 13 1 14 13 1 10 0 9 2 4 15 3 3 1 10 0 4 13 1 9 9 7 9 9 2
11 10 9 2 10 9 2 15 13 1 9 2
5 7 15 13 15 2
12 15 13 2 15 9 10 0 9 4 13 1 2
28 15 4 3 10 9 13 14 13 9 1 9 1 10 0 9 7 10 0 9 1 11 2 3 3 4 15 13 2
5 1 9 1 9 2
15 10 9 4 15 13 10 9 1 12 9 2 2 13 9 2
10 3 4 15 3 13 3 1 12 3 2
26 2 15 13 3 3 15 2 15 13 1 2 16 15 3 4 13 1 10 12 9 2 15 4 13 1 2
42 10 0 9 13 3 9 1 2 16 9 1 11 4 13 1 14 13 2 16 10 0 9 1 9 1 11 13 3 1 2 16 10 0 7 0 9 4 13 1 0 11 2
16 15 4 3 0 1 9 2 16 15 4 13 1 9 0 9 2
20 3 13 15 3 2 15 3 4 13 10 0 9 2 1 14 13 9 1 15 2
4 3 13 9 2
14 9 4 13 9 1 10 0 9 1 9 1 11 11 2
15 1 0 9 13 11 11 2 11 1 11 9 2 1 9 2
25 15 13 10 9 0 9 2 7 15 13 3 0 9 2 15 13 1 15 15 2 2 13 11 11 2
18 1 10 9 4 10 9 9 1 10 0 9 1 0 9 1 0 9 2
14 1 9 4 9 3 13 7 13 9 0 9 1 9 2
20 10 10 9 1 9 4 9 13 1 3 0 9 1 9 7 9 1 1 9 2
44 11 13 9 3 1 11 2 7 1 9 12 4 9 13 1 0 11 1 9 1 0 9 2 15 3 3 13 15 7 13 2 16 15 13 9 1 14 4 9 1 10 0 9 2
22 15 2 16 15 9 13 0 9 1 9 7 9 2 13 9 1 10 0 9 3 3 2
15 11 11 2 9 1 9 2 4 13 9 12 9 1 11 2
18 7 15 4 3 0 2 7 16 10 0 13 9 2 13 15 1 9 2
32 11 9 4 3 3 3 1 9 1 10 0 9 2 16 10 0 0 9 4 0 1 2 16 9 13 1 9 9 1 9 12 2
17 9 4 13 9 7 9 9 1 10 9 2 15 4 0 7 0 2
12 15 4 3 10 0 1 9 2 15 11 13 2
6 15 13 15 1 9 2
14 9 1 9 4 10 0 9 1 14 13 3 1 9 2
19 3 13 3 0 9 1 2 16 15 4 13 0 1 11 1 14 13 9 2
17 7 15 13 10 10 9 2 7 15 13 15 2 2 13 11 11 2
37 2 15 13 10 1 9 7 0 9 1 15 4 2 7 15 4 0 1 2 16 15 4 13 9 1 9 9 12 2 2 13 11 11 3 1 9 2
28 2 1 3 12 9 1 10 0 9 4 15 0 2 16 15 1 9 4 13 1 9 1 11 1 9 1 9 2
43 2 16 3 13 9 1 10 0 9 1 0 9 1 2 3 4 15 3 13 9 1 9 2 7 0 9 1 9 4 3 13 1 9 2 2 13 9 11 11 2 9 9 2
15 2 1 13 4 15 3 0 2 16 15 4 3 1 9 2
9 1 10 0 2 9 13 9 3 2
19 9 4 0 1 14 13 1 9 1 10 9 1 11 2 13 9 11 11 2
15 11 11 1 11 4 10 9 1 0 9 13 1 0 9 9
28 3 13 9 10 9 1 10 0 9 9 2 16 15 4 13 2 16 15 13 10 9 7 13 9 1 10 9 2
11 2 11 13 3 1 14 13 9 1 9 2
28 13 15 2 16 16 10 9 13 15 1 14 13 0 9 2 7 1 0 0 9 2 13 9 1 14 4 0 2
22 1 10 9 13 1 9 11 1 11 13 3 3 3 0 9 9 1 10 12 0 9 2
23 2 15 4 15 1 9 9 9 0 9 2 3 3 4 0 0 9 2 1 10 13 9 2
24 2 11 13 3 3 2 0 7 0 7 13 1 9 7 9 7 13 15 2 16 15 4 3 2
14 1 9 1 9 11 11 11 7 1 9 11 11 11 2
14 15 4 3 13 16 3 13 10 9 1 9 10 9 2
21 10 0 9 13 15 3 1 10 0 9 1 12 9 2 1 9 1 9 1 9 2
9 13 9 2 7 13 15 3 13 2
4 11 13 3 2
32 4 15 10 9 13 3 3 1 10 9 1 12 9 1 14 4 13 10 9 3 1 1 9 7 1 9 1 10 3 0 9 2
15 3 4 10 0 9 0 9 2 3 9 1 9 4 0 2
20 9 1 12 9 1 9 4 0 7 9 13 15 13 13 1 9 1 0 9 2
24 15 1 9 1 10 9 4 4 2 2 4 15 3 13 15 2 16 9 13 15 3 3 2 2
3 3 5 12
7 2 15 4 0 2 0 2
24 0 1 10 3 13 0 9 4 3 10 0 9 1 9 7 9 7 3 0 9 1 0 9 2
14 3 15 1 11 9 13 1 2 15 4 13 1 11 2
1 9
13 2 15 4 3 10 9 2 16 15 13 1 9 2
9 15 13 1 10 0 9 7 13 2
31 9 13 3 1 9 1 9 1 14 13 9 1 14 13 15 1 13 9 2 16 11 9 1 9 4 13 1 10 0 9 2
6 10 9 4 3 9 2
14 10 10 0 9 4 14 13 10 0 9 13 1 11 2
29 9 1 10 9 4 13 15 13 2 16 15 13 15 1 10 13 9 2 15 13 10 9 2 15 4 9 1 9 2
40 0 2 13 9 7 9 1 9 1 0 2 0 9 13 15 1 10 0 2 11 2 2 11 11 11 11 2 12 2 3 1 14 13 15 10 9 7 10 9 2
21 15 4 13 1 9 1 10 9 2 15 3 4 13 1 9 12 1 9 11 11 2
25 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 7 9 1 0 9 2
20 9 4 13 3 2 16 15 4 13 9 1 10 9 3 1 10 9 7 9 2
20 1 9 4 11 3 13 10 10 7 3 0 9 2 11 11 12 1 12 9 2
12 15 4 3 13 1 0 9 1 11 11 9 2
3 4 13 3
14 3 2 16 15 3 13 2 16 15 4 13 15 13 2
6 1 14 13 10 9 2
19 9 4 3 13 3 3 7 7 13 10 9 3 2 1 15 13 15 1 2
12 13 9 7 9 1 10 9 1 12 9 9 2
14 10 9 3 4 13 3 1 9 1 1 12 1 9 2
15 13 10 13 9 3 10 9 7 3 1 0 9 1 3 2
25 9 1 10 0 9 9 1 9 1 10 0 9 4 13 9 1 11 9 1 14 13 9 1 9 2
31 9 13 1 10 9 2 11 10 0 0 9 4 13 1 3 0 9 1 11 2 11 7 11 2 1 14 13 10 12 9 2
1 2
27 3 4 3 1 0 9 13 9 1 9 3 1 11 9 2 3 1 9 12 9 4 4 13 1 0 9 2
4 3 13 15 2
34 11 11 2 9 1 10 0 9 1 11 2 4 1 9 13 10 12 9 9 2 7 15 13 1 3 0 9 1 9 12 0 0 9 2
23 1 0 9 9 7 0 0 9 4 12 9 13 3 1 2 16 15 4 4 3 1 9 2
20 7 9 13 0 9 1 11 11 2 15 13 9 1 9 1 9 1 13 9 2
11 3 4 15 3 3 13 10 9 3 2 2
13 15 13 9 9 2 15 4 13 10 0 9 3 2
21 11 13 0 1 0 9 2 3 13 15 15 3 1 15 15 7 13 3 1 15 2
7 10 0 9 13 1 9 2
19 11 11 9 11 11 13 3 2 16 9 4 13 1 10 9 1 12 9 2
19 2 15 13 15 2 13 15 3 2 13 9 1 10 9 7 13 15 3 2
12 16 15 4 13 2 4 15 0 14 13 9 2
15 11 10 9 2 3 11 2 13 3 11 7 11 1 9 2
10 15 4 4 13 2 13 9 3 2 2
7 0 9 4 9 15 13 2
15 3 13 11 2 11 7 10 0 10 0 9 3 1 9 2
16 16 10 9 13 1 9 10 9 2 4 0 13 3 1 11 2
2 0 9
24 7 16 15 13 2 4 15 3 3 3 2 16 15 10 9 13 7 15 4 13 1 9 9 2
4 9 4 0 2
32 7 3 13 9 10 0 9 2 13 11 2 15 13 2 16 15 1 0 9 13 15 1 10 9 2 16 15 4 13 10 9 2
4 10 0 9 2
36 15 4 4 9 1 9 9 2 9 1 9 1 0 0 9 2 1 9 1 9 1 9 2 1 9 1 0 9 7 9 1 9 1 11 9 2
38 15 4 0 2 7 9 4 3 3 3 0 2 2 13 11 11 2 16 15 13 1 2 16 9 1 9 1 9 13 1 12 1 12 1 12 1 12 2
1 9
17 3 4 15 13 15 14 13 2 7 15 4 13 1 14 13 3 2
8 10 9 1 9 4 10 9 2
9 11 8 8 8 8 8 8 8 2
25 0 10 9 1 15 2 3 4 3 0 2 3 2 1 9 1 0 10 0 2 10 9 4 13 2
10 13 1 9 4 9 0 9 1 9 2
48 9 13 2 16 10 9 9 7 9 1 9 7 9 12 13 2 16 2 11 2 1 9 1 10 0 9 2 10 0 9 7 3 9 1 11 2 7 10 9 1 11 13 9 1 9 1 11 2
4 3 13 15 2
6 3 4 15 13 15 2
4 0 9 1 9
1 9
11 9 13 3 1 13 2 0 7 0 9 2
35 0 4 15 2 15 9 15 13 2 15 13 15 0 9 2 16 9 9 13 1 9 9 2 16 10 9 7 10 9 3 3 4 4 9 2
41 7 4 15 13 3 1 9 2 4 15 13 2 16 10 9 1 9 7 9 1 14 13 9 1 15 13 1 9 1 9 2 13 9 1 9 2 9 11 11 11 2
2 12 9
23 2 15 4 3 3 14 13 1 13 9 2 2 13 11 1 9 1 10 0 9 1 12 2
26 15 4 15 1 11 7 11 9 4 3 0 2 16 15 4 13 9 1 9 1 10 12 2 9 2 2
25 11 13 15 1 10 0 9 2 16 11 3 13 9 1 10 0 9 7 9 2 15 13 1 9 2
16 2 9 7 9 4 3 13 7 13 1 9 2 2 13 15 2
15 3 1 9 9 7 9 13 10 9 9 1 9 1 9 2
16 3 13 3 9 1 2 3 0 9 9 9 13 3 1 9 2
34 1 10 0 13 15 10 0 9 9 1 10 9 2 16 15 4 13 3 1 15 2 15 13 2 8 8 8 2 2 9 1 9 2 2
28 7 3 4 15 1 3 0 9 2 15 4 13 1 0 9 2 7 3 13 3 10 9 2 3 4 3 0 2
14 3 16 9 13 14 13 7 13 3 1 9 1 9 2
4 1 9 1 9
20 7 16 15 4 13 10 0 9 4 11 11 11 3 3 13 9 1 15 2 2
19 9 1 10 0 9 2 0 11 11 1 11 2 4 13 0 0 0 9 2
15 3 13 3 10 9 9 2 1 15 10 9 7 12 9 2
29 9 13 9 1 9 3 12 1 9 2 3 1 16 9 1 12 9 7 10 0 9 1 9 13 1 11 11 9 2
8 10 0 10 2 3 14 13 2
32 0 13 3 9 1 14 13 3 14 13 10 0 7 4 3 1 0 9 2 7 0 13 13 2 16 15 13 10 0 9 0 2
2 9 3
6 9 1 10 9 13 2
14 15 13 14 13 9 1 10 0 9 1 13 1 9 12
11 3 13 10 0 9 3 3 1 10 0 2
1 9
18 7 15 13 15 3 16 10 0 9 9 3 4 13 9 7 9 0 2
25 3 13 9 1 9 2 16 10 0 9 1 11 3 3 4 13 10 9 2 15 4 13 9 0 2
19 7 15 4 13 3 1 0 9 2 7 3 4 15 4 13 3 1 9 2
25 3 1 11 9 2 3 15 1 9 1 9 1 9 13 0 9 7 9 1 9 2 9 12 9 2
24 0 9 7 0 9 13 2 16 3 3 4 13 0 9 1 10 0 9 1 9 1 10 0 2
18 15 4 0 14 13 2 16 11 9 4 4 3 0 1 11 9 2 2
13 9 13 2 16 9 13 10 0 9 1 3 9 2
20 3 1 11 0 9 1 11 0 9 13 10 0 9 9 1 10 9 1 11 2
4 13 15 15 2
10 3 13 15 2 3 3 9 4 9 2
13 2 3 13 15 2 16 10 9 4 13 15 0 2
32 7 3 1 9 3 4 10 0 2 9 2 2 15 4 13 1 2 3 4 15 10 0 9 1 9 7 10 0 9 2 11 2
14 11 13 10 9 3 2 15 9 1 9 13 1 9 2
13 11 11 11 13 2 2 15 4 3 0 1 9 2
28 1 14 13 9 3 2 3 4 3 13 10 9 1 9 7 9 1 3 12 9 2 1 10 11 3 12 9 2
41 9 1 9 1 10 0 9 4 3 4 13 1 9 1 10 13 9 2 15 4 13 9 1 15 3 1 10 0 9 1 11 2 15 4 13 9 1 11 1 9 2
1 11
21 2 15 9 15 13 9 2 13 15 13 9 2 0 9 2 13 9 7 0 9 2
24 7 15 13 3 1 9 2 15 13 3 3 9 1 14 4 0 2 11 11 13 1 10 9 2
18 3 13 3 10 9 14 13 9 3 1 2 7 15 13 1 14 13 2
4 15 13 13 2
7 9 13 10 9 9 3 2
36 1 0 9 4 15 13 13 3 7 13 10 9 13 1 9 2 7 13 10 9 9 1 14 13 2 16 10 9 13 7 13 3 1 10 9 2
12 15 4 3 13 9 2 15 4 15 13 1 2
17 9 13 9 7 9 1 9 7 13 1 9 1 9 1 0 9 2
20 15 4 13 15 3 3 0 9 14 13 2 0 4 9 2 1 10 0 9 2
22 1 9 4 3 13 0 9 10 0 9 2 7 10 0 9 4 1 12 7 12 9 2
19 11 11 2 0 9 2 4 1 11 13 1 9 1 10 0 9 11 11 2
15 3 4 9 1 9 1 9 1 10 9 1 11 7 11 2
7 2 3 13 15 1 9 2
15 2 15 13 3 0 9 2 3 1 10 8 0 9 2 2
27 10 9 1 9 11 9 13 2 16 9 1 9 13 14 2 13 13 9 1 11 11 7 13 11 9 2 2
11 15 4 13 9 0 2 12 9 1 9 2
36 9 1 10 0 9 2 11 11 2 7 10 0 9 2 11 11 2 13 1 2 13 9 13 2 2 15 13 10 11 1 0 0 9 1 12 2
9 7 15 4 3 13 10 0 9 2
15 10 9 3 4 15 2 15 3 4 13 2 3 13 3 2
11 7 1 9 12 13 9 10 0 9 12 2
7 13 9 5 9 9 5 8
4 2 12 9 2
9 7 10 9 4 10 0 9 13 2
15 15 4 13 3 3 2 16 15 1 3 13 14 13 9 2
27 15 13 3 10 0 9 0 9 2 7 15 4 3 13 3 1 9 1 14 13 1 14 13 3 1 9 2
9 3 4 9 3 13 10 0 9 2
14 2 15 9 4 15 13 15 2 2 13 15 3 3 2
25 15 13 3 2 16 9 13 1 13 1 9 9 2 7 3 1 9 13 15 10 9 1 10 9 2
10 9 4 13 0 1 0 9 1 9 2
10 2 15 4 9 2 16 15 13 3 2
11 9 11 11 13 9 1 9 1 11 9 2
21 0 9 4 3 0 1 9 2 7 1 0 9 2 3 3 12 9 13 1 9 2
22 11 2 2 15 4 3 0 7 0 9 1 9 9 2 16 15 3 13 9 1 9 2
4 10 0 9 2
8 2 6 2 3 10 0 15 2
13 15 13 15 3 1 2 3 15 4 13 9 13 2
14 3 8 3 1 9 9 2 15 3 4 13 1 15 2
8 13 13 1 14 13 1 15 2
34 11 11 11 2 1 3 4 0 1 10 0 9 2 4 13 9 1 10 0 9 1 9 2 15 13 3 1 9 1 9 10 0 9 2
18 2 9 2 4 4 10 0 9 9 7 9 1 14 4 13 1 0 2
17 7 4 9 13 3 2 4 15 3 13 15 1 0 9 1 9 2
69 9 4 10 9 2 3 10 9 2 16 16 10 0 9 13 3 1 14 13 10 0 9 1 14 4 13 1 0 9 1 9 2 4 9 3 3 1 10 9 13 1 14 4 0 2 1 13 1 9 11 11 7 1 10 3 0 9 1 11 9 2 1 4 0 1 10 0 9 2
27 16 9 3 15 13 1 9 1 14 13 10 13 9 2 4 15 1 0 9 13 9 1 0 7 0 9 2
45 2 13 2 1 16 3 3 3 3 0 1 0 9 2 2 13 15 3 1 12 9 1 11 2 11 7 11 2 11 9 7 11 1 11 2 15 0 4 13 9 1 10 9 9 2
7 2 15 4 3 13 15 2
18 9 13 2 16 11 11 3 13 10 0 9 3 1 10 9 1 11 2
13 3 13 15 10 9 9 2 15 15 13 3 3 2
44 3 13 10 0 9 2 7 3 4 9 10 9 2 3 15 10 0 9 2 7 3 13 15 3 7 13 10 0 9 2 16 3 3 3 13 9 1 9 1 10 3 0 9 2
1 9
23 10 0 1 9 13 2 16 10 3 13 9 1 8 7 9 13 10 9 3 1 9 9 2
25 1 9 1 11 4 10 0 9 13 15 1 10 0 13 1 10 0 9 1 9 1 9 7 9 2
33 11 11 4 1 10 0 9 3 13 9 1 9 1 2 16 0 9 1 9 4 13 0 9 3 1 9 2 15 15 13 1 9 2
8 0 1 15 13 9 1 9 2
14 3 13 15 1 14 13 0 10 0 9 3 1 9 2
4 12 9 1 9
31 3 13 15 3 2 1 9 9 10 0 9 9 12 2 13 1 9 9 1 12 12 12 12 1 9 10 0 9 9 12 2
22 15 4 1 10 0 9 10 0 9 2 15 13 9 2 1 3 1 3 4 13 1 2
1 9
14 16 4 15 3 7 3 4 15 3 2 13 8 11 2
83 1 3 4 15 3 13 10 9 2 15 3 4 13 8 1 11 9 2 1 1 9 14 4 3 13 0 1 9 1 9 2 7 9 1 9 9 2 9 11 11 2 3 15 1 11 11 4 3 3 2 13 2 16 3 4 9 1 9 2 13 1 9 7 9 1 9 7 9 1 9 7 9 2 13 10 9 2 15 13 9 1 9 2
11 10 9 2 15 13 9 2 9 7 9 2
13 15 13 3 0 0 9 1 15 1 9 13 1 2
15 15 4 3 14 13 3 0 1 2 16 9 4 4 0 2
13 11 13 3 9 1 11 9 2 7 9 4 13 2
9 10 9 13 0 1 10 9 13 2
13 10 9 13 2 7 4 3 0 2 1 10 9 2
47 2 9 13 0 1 10 9 1 9 9 2 7 15 4 13 11 9 11 11 11 7 11 11 14 13 10 9 2 15 13 3 3 1 10 0 9 2 7 3 4 15 13 9 3 3 2 2
21 15 13 10 9 1 2 15 15 13 2 11 11 13 2 15 4 13 3 1 9 2
12 1 15 13 9 15 14 13 1 14 13 2 2
17 2 7 3 2 3 13 15 1 15 2 15 13 1 10 10 9 2
15 1 14 4 13 3 2 4 15 3 0 1 10 0 9 2
18 15 4 3 3 13 2 3 4 15 0 9 2 15 10 9 13 11 2
3 12 9 9
46 2 4 3 0 7 3 3 0 9 13 1 9 2 4 15 3 13 2 16 10 0 9 3 4 4 0 1 14 13 3 7 13 9 1 10 9 2 2 13 15 1 10 0 9 9 2
6 11 13 3 1 9 9
2 0 9
15 15 4 3 13 10 0 9 2 15 13 0 1 10 9 2
18 2 15 4 3 13 9 1 9 1 9 2 1 9 2 9 2 2 2
23 11 9 4 0 9 9 1 10 0 1 10 9 9 2 10 0 9 11 11 13 1 11 2
27 15 1 10 12 13 0 9 4 10 3 0 9 11 2 1 3 4 3 0 3 1 9 7 10 13 9 2
13 10 9 4 15 13 9 1 10 12 9 0 8 2
33 1 9 1 10 0 9 13 11 1 12 9 2 11 11 2 11 11 7 11 11 2 1 10 9 2 15 4 13 1 9 0 9 2
9 13 15 9 2 3 13 15 3 2
13 8 13 3 1 3 3 15 2 15 4 13 9 2
8 13 7 13 15 9 3 3 2
20 2 15 13 0 9 1 2 16 10 9 13 0 2 16 15 13 12 9 2 2
28 10 0 9 13 15 2 16 9 11 13 1 14 13 1 9 2 7 9 13 3 1 9 3 7 9 4 0 2
5 6 2 13 15 2
53 0 9 13 9 7 9 2 7 10 0 1 9 13 1 9 2 15 13 3 7 3 2 15 15 13 1 9 2 9 2 9 2 9 2 15 13 10 0 9 2 15 9 3 13 9 2 7 13 0 1 14 13 2
22 9 1 2 11 11 2 4 0 7 0 2 15 13 1 9 1 9 7 1 9 9 2
9 2 15 13 9 13 0 9 3 2
49 3 4 8 13 10 9 1 9 1 10 0 9 2 15 4 13 9 1 10 9 2 15 3 4 13 9 1 10 9 1 9 2 3 3 4 0 9 7 9 1 14 13 0 9 1 14 13 9 2
9 3 9 4 13 11 0 1 9 2
31 11 4 13 1 0 9 1 10 13 9 7 4 13 0 9 7 9 3 1 15 15 7 1 10 9 1 10 12 0 9 2
13 15 1 15 13 1 3 9 2 2 13 11 11 2
25 3 13 15 11 11 1 11 9 2 7 3 1 10 0 13 15 3 1 11 9 1 10 0 9 2
13 7 3 3 9 13 1 9 2 15 13 3 9 2
12 15 13 10 3 3 0 9 1 8 7 9 2
19 7 15 13 3 1 9 9 1 9 7 9 2 11 11 13 9 1 9 2
25 3 13 1 9 1 11 7 1 10 9 1 11 2 3 15 1 10 9 4 4 13 1 0 9 2
20 15 13 1 14 13 2 11 4 13 15 1 10 9 2 7 15 4 13 15 2
21 3 13 15 1 9 9 11 11 2 3 4 0 9 7 4 13 12 1 12 9 2
5 9 4 0 0 9
7 15 13 3 3 1 11 2
7 11 13 3 15 1 13 2
12 15 4 3 3 13 2 15 15 3 3 13 2
9 9 13 1 10 9 1 8 9 2
14 15 4 12 3 13 0 9 2 15 3 13 0 9 2
22 2 7 15 13 14 13 9 13 10 9 1 9 2 2 13 9 11 11 11 1 11 2
28 7 15 13 15 9 14 13 2 15 0 9 15 4 13 1 9 3 1 10 0 9 1 9 1 9 7 9 2
9 0 9 1 9 7 10 0 9 2
2 0 9
14 9 4 9 9 2 7 9 13 9 1 14 13 10 9
8 0 7 0 9 13 15 3 2
26 1 9 12 4 11 9 3 1 12 10 0 9 13 1 14 4 3 1 10 0 9 2 11 11 11 2
11 10 12 9 13 10 9 1 0 1 9 2
18 15 4 0 3 13 15 1 10 10 9 2 16 15 13 3 12 9 2
13 9 13 1 11 1 11 7 1 9 3 1 11 2
10 10 10 9 13 10 9 2 15 13 2
29 9 13 0 9 9 7 10 9 1 15 9 9 1 8 2 9 1 3 0 9 7 9 1 9 7 8 7 9 2
17 13 16 10 9 13 7 3 4 13 3 1 3 12 9 0 9 2
11 0 4 13 0 3 1 11 9 1 11 2
11 9 12 4 13 1 8 0 9 1 12 2
47 11 11 4 3 13 3 1 9 1 9 1 11 9 2 9 11 11 2 7 3 1 9 1 11 9 4 15 13 14 13 11 1 10 0 9 9 1 9 1 9 1 10 9 1 9 9 2
25 15 13 15 3 1 14 13 1 10 9 0 9 1 12 9 9 7 10 0 2 0 9 1 9 2
34 2 7 15 4 3 10 0 9 1 11 2 7 3 4 15 3 13 15 3 7 13 15 1 15 3 13 15 15 13 15 1 14 13 2
21 9 9 2 15 3 13 10 0 9 1 11 9 2 4 3 3 13 1 0 9 2
8 2 15 4 3 0 1 15 2
22 3 1 11 11 16 15 9 13 7 13 1 10 9 1 0 13 7 9 1 11 9 2
28 7 1 0 9 13 9 15 1 15 2 7 15 13 1 10 0 9 1 9 1 9 7 9 3 1 9 9 2
46 7 15 4 3 15 1 10 0 2 3 16 15 13 1 2 16 15 4 3 1 10 9 2 15 4 14 13 1 10 0 9 3 1 14 13 1 10 0 9 2 2 13 11 11 11 2
27 16 15 13 11 9 1 10 0 7 10 0 9 1 15 2 13 15 2 13 2 16 9 4 13 10 9 2
51 15 13 15 1 3 0 2 16 10 0 11 1 10 0 9 1 10 0 1 9 9 13 15 3 1 9 1 10 9 2 9 7 9 1 8 7 9 2 15 9 13 10 3 0 7 0 9 1 9 9 2
14 11 11 13 2 16 9 2 13 15 1 9 9 2 2
9 15 4 3 0 16 9 4 13 2
24 3 3 1 10 0 9 2 15 1 10 9 13 1 14 4 13 1 0 9 7 3 13 2 2
25 3 9 3 1 10 0 2 0 9 2 1 9 2 9 2 9 7 9 13 10 0 0 0 9 2
16 7 1 9 13 2 13 9 2 7 9 13 0 7 0 9 2
17 10 0 7 0 9 4 3 13 15 9 1 14 13 0 10 9 2
1 9
19 15 13 1 9 11 2 3 10 0 0 9 13 10 9 1 10 0 9 2
12 11 13 10 9 2 1 15 13 14 13 15 2
1 0
8 3 4 9 4 10 0 9 2
34 3 4 15 13 9 3 3 1 10 9 2 14 13 13 10 3 12 9 0 9 2 15 13 9 9 1 14 13 2 1 15 4 13 2
19 1 0 9 13 3 11 3 1 3 1 9 14 4 4 13 3 1 9 2
27 9 11 11 13 0 9 1 2 16 9 3 7 3 4 13 7 13 10 0 9 2 7 3 13 13 9 2
10 15 4 9 2 15 13 0 9 0 2
16 1 3 4 15 13 1 12 7 12 0 9 1 10 9 2 2
10 7 15 13 3 0 1 10 9 2 2
3 15 13 2
22 3 1 10 3 13 9 1 9 13 15 10 9 2 15 9 0 9 13 1 0 9 2
8 2 9 13 13 1 11 9 2
5 9 4 4 0 2
6 3 13 15 10 9 2
41 15 13 2 11 2 1 9 1 0 9 2 3 15 4 13 1 15 1 9 1 10 9 1 9 2 15 1 9 4 13 3 1 9 1 11 2 11 2 1 11 2
22 9 7 9 1 9 1 0 7 3 0 9 1 15 4 13 15 14 13 10 0 9 2
25 3 3 3 4 15 3 3 13 2 7 10 13 0 9 4 3 13 2 16 3 13 15 1 9 2
31 11 4 4 9 11 7 11 0 9 1 10 0 9 1 10 0 9 2 7 3 10 0 9 1 10 9 1 15 13 0 2
10 7 15 13 9 1 9 2 1 15 2
63 9 13 1 10 9 9 3 1 9 1 8 2 8 7 9 2 3 13 9 1 9 1 9 2 16 15 13 1 12 9 1 9 1 9 1 10 13 9 2 1 10 9 3 1 9 2 4 15 3 0 2 16 10 9 4 13 3 3 1 9 1 9 2
12 3 13 15 12 9 1 10 0 0 9 3 2
27 2 15 4 10 9 2 16 0 9 9 4 13 13 1 10 0 9 7 3 13 7 13 3 1 12 9 2
24 10 0 9 12 13 11 9 1 11 11 9 2 16 9 4 13 12 9 1 9 1 11 11 2
8 9 1 12 9 1 0 9 2
24 11 11 2 15 15 13 9 9 1 11 13 11 10 9 2 16 15 13 9 7 9 1 9 2
11 7 3 1 1 12 13 15 15 1 9 2
43 10 0 9 13 1 9 2 16 15 3 4 13 14 13 2 15 15 4 13 1 2 7 16 15 4 4 10 0 9 1 15 2 7 16 15 13 1 2 16 15 4 0 2
26 10 12 9 2 11 9 7 11 9 2 4 13 10 0 9 1 11 2 15 4 13 9 1 10 9 2
7 10 9 4 0 7 0 2
22 15 4 13 14 13 1 0 9 2 7 4 3 13 15 1 2 16 15 13 15 13 2
8 2 10 9 13 9 1 9 2
16 7 15 4 3 10 13 9 2 15 1 3 13 9 1 11 2
28 0 9 13 1 2 16 15 1 10 0 9 13 3 1 9 9 1 14 13 10 9 1 2 3 0 9 13 2
10 9 4 3 3 3 13 1 11 9 2
19 1 10 0 9 2 7 11 11 3 0 9 1 9 2 4 9 10 9 2
32 7 11 11 13 3 3 15 1 9 1 9 2 16 15 15 13 1 9 2 3 1 11 11 1 0 9 13 1 3 0 9 2
11 9 1 2 3 9 4 13 2 4 0 2
22 15 13 0 10 0 9 9 7 13 1 9 2 16 9 9 7 9 4 10 0 9 2
22 15 4 9 2 3 4 0 2 9 1 10 13 9 2 3 3 4 0 7 0 2 2
26 11 2 13 10 0 9 1 11 11 7 10 9 2 11 11 11 2 15 13 10 9 1 12 9 3 2
12 2 15 4 3 3 0 2 15 4 3 0 2
12 1 10 9 13 15 3 3 1 9 7 0 2
2 13 9
19 10 12 9 4 1 9 1 9 13 1 10 9 1 10 0 9 2 11 2
8 2 4 15 3 4 3 0 2
11 10 12 9 13 1 10 9 10 0 9 2
19 11 11 9 2 11 11 2 2 10 9 4 3 10 9 1 0 11 9 2
32 7 9 1 10 0 9 2 3 1 9 13 8 2 4 3 13 1 2 16 15 1 0 9 13 1 9 1 14 13 9 9 2
10 15 13 3 1 10 9 1 13 9 2
8 15 13 3 3 9 1 9 2
22 12 9 9 12 9 1 9 2 7 1 9 4 3 1 12 9 1 9 1 15 15 2
12 15 4 13 2 16 9 13 1 9 1 9 2
7 9 2 3 2 4 12 9
34 1 9 13 15 0 7 3 7 1 10 9 2 15 4 13 10 3 0 9 1 9 9 1 9 1 9 2 1 9 1 2 11 2 2
22 1 11 4 9 13 10 0 9 1 10 0 9 2 10 9 2 9 7 9 2 9 2
21 9 13 13 9 1 9 2 16 15 4 13 15 3 7 13 9 2 15 4 13 9
14 2 16 11 13 2 13 15 3 2 15 3 4 13 2
20 15 13 15 13 2 11 11 11 2 2 13 15 2 7 13 10 12 9 0 2
2 3 13
7 3 4 11 8 9 9 2
22 3 4 10 0 0 11 11 7 9 11 11 11 13 0 1 9 2 16 15 4 13 2
25 2 15 13 3 8 13 1 9 2 16 16 15 4 13 10 9 1 9 2 3 4 9 13 13 2
10 9 0 9 13 15 3 14 4 0 2
9 15 13 3 3 3 3 9 1 2
14 9 4 10 9 2 7 15 13 3 1 9 7 9 2
33 11 11 13 10 0 7 0 9 2 15 1 10 0 7 0 9 10 9 3 3 1 9 13 1 9 1 9 2 15 4 13 9 2
13 1 9 1 9 4 11 3 13 1 10 0 9 2
22 9 7 9 2 3 0 2 9 4 4 13 1 9 2 16 10 0 4 13 9 9 2
9 3 13 12 9 1 9 1 9 2
18 10 9 13 1 9 1 10 0 9 2 15 13 10 9 1 0 9 2
23 2 15 4 13 9 2 7 3 4 15 3 13 10 9 2 7 15 13 15 3 14 13 2
29 7 9 4 10 9 1 10 0 0 9 2 10 9 9 2 1 10 0 9 7 0 9 3 2 2 13 11 11 2
29 11 4 9 1 11 2 7 4 13 7 13 1 9 7 9 1 11 7 1 11 2 3 15 13 1 3 1 12 2
12 2 15 13 9 9 1 14 13 15 1 15 2
7 7 15 3 3 13 15 2
12 10 9 4 3 13 1 0 9 1 0 9 2
5 15 13 15 3 2
14 15 4 3 13 9 1 9 1 16 15 4 13 15 2
14 11 11 13 9 1 9 2 9 7 10 0 0 9 2
25 1 11 2 3 12 9 4 4 13 7 13 3 2 4 12 0 9 4 13 3 1 0 0 9 2
27 2 15 13 0 9 1 9 2 16 15 4 13 1 2 16 15 4 13 1 14 13 3 1 2 9 2 2
8 13 1 10 9 9 1 9 2
21 2 7 0 2 3 13 15 3 1 15 2 13 15 2 7 13 13 1 0 9 2
49 1 9 13 15 15 1 10 9 0 9 1 10 0 9 2 7 3 13 3 10 9 2 15 13 9 3 1 9 2 2 13 10 0 9 2 15 4 9 1 9 7 9 1 9 2 16 9 13 2
13 3 1 11 13 9 9 1 9 7 9 1 9 2
25 16 11 11 13 10 2 11 2 11 11 11 2 1 9 12 9 3 2 13 9 3 10 10 9 2
15 7 15 13 9 1 2 10 3 0 9 1 9 9 2 2
27 9 2 13 1 9 2 7 13 9 2 4 2 1 15 9 13 2 10 0 7 3 13 9 1 11 9 2
2 9 12
29 9 2 13 9 1 9 2 13 15 3 2 13 9 3 2 13 9 7 9 2 13 3 1 9 2 13 13 9 2
10 7 9 2 11 2 4 10 0 9 2
4 10 9 0 9
20 10 9 13 15 11 1 10 9 9 14 13 3 1 9 7 13 10 0 9 2
29 10 12 9 13 3 9 1 10 0 9 1 10 0 9 2 15 1 10 9 13 3 1 0 1 10 0 0 9 2
12 7 15 4 15 3 13 2 2 13 11 11 2
20 10 9 1 10 0 9 4 13 8 3 2 15 4 13 10 9 1 15 9 2
13 15 13 8 0 1 11 11 1 11 9 9 9 2
49 15 13 1 9 2 16 10 0 9 1 9 4 10 9 9 2 10 9 2 15 3 13 2 7 3 15 3 13 10 9 3 2 15 13 3 2 1 9 1 14 13 7 13 15 1 10 0 9 2
17 3 13 2 16 3 4 13 10 0 9 1 9 1 9 1 9 2
11 11 4 13 3 3 0 11 13 1 11 2
14 1 9 13 3 10 9 1 2 16 11 11 13 15 2
3 12 4 3
5 1 11 1 0 9
24 1 9 4 10 9 0 1 14 13 9 3 1 9 2 9 2 9 2 7 11 1 11 9 2
22 1 9 1 12 13 9 0 7 3 0 1 3 2 7 8 13 1 11 1 3 3 2
21 7 3 13 15 2 16 9 4 13 1 14 13 12 9 7 13 0 9 1 9 2
37 15 13 2 16 15 1 14 13 10 9 9 0 9 7 12 9 15 9 13 10 0 9 7 0 10 10 9 1 9 2 15 4 13 9 9 3 2
17 15 4 3 0 1 2 16 15 4 4 9 2 7 3 13 13 2
17 15 13 3 1 10 0 9 1 0 9 7 10 0 2 0 9 2
2 0 9
10 9 13 3 2 2 15 13 15 3 2
2 0 2
16 2 16 3 15 13 3 2 13 15 0 9 2 2 13 11 2
19 10 9 13 2 16 15 4 13 15 1 9 2 7 3 3 13 15 3 2
22 15 4 3 13 2 16 15 4 2 0 2 9 2 16 15 3 13 9 1 11 9 2
6 2 6 2 3 3 2
13 7 15 4 15 3 13 15 2 16 15 13 2 2
21 3 4 15 3 0 16 0 0 9 4 13 1 14 13 10 9 1 10 9 13 2
8 15 4 3 3 13 7 13 2
12 7 15 7 11 4 3 13 15 14 13 1 2
12 3 7 0 1 14 13 9 1 9 7 9 2
11 15 4 3 13 1 9 11 1 3 0 2
22 1 9 13 15 1 11 11 2 12 2 15 13 11 11 10 9 1 10 9 1 9 2
39 9 2 9 2 9 2 9 2 0 9 2 7 3 3 0 9 2 13 10 9 2 1 3 4 4 3 0 2 7 1 15 3 13 0 10 9 1 11 2
71 11 13 3 9 11 11 1 9 1 11 9 2 16 15 1 10 9 1 10 0 9 2 11 2 13 2 16 2 15 4 0 2 16 11 9 2 3 4 10 9 1 10 9 2 15 1 3 0 9 13 1 0 9 2 13 14 13 10 9 2 15 4 13 10 9 2 15 9 13 2 2
3 11 4 0
9 13 15 0 2 16 15 4 0 2
9 11 11 1 15 1 10 0 9 2
11 13 15 13 15 15 8 2 9 13 3 2
12 1 15 13 1 9 4 0 13 10 9 3 2
18 10 9 9 1 11 4 3 3 13 9 3 2 16 15 13 1 9 2
26 1 10 9 13 15 2 16 9 4 13 3 1 2 9 7 9 2 3 3 7 1 9 7 9 9 2
26 3 13 15 1 14 13 9 1 10 9 1 0 9 2 16 16 9 13 2 13 3 10 9 1 9 2
38 10 9 9 2 9 1 11 2 11 11 8 11 11 2 2 9 1 11 2 11 11 11 7 9 2 2 9 1 11 2 11 7 11 7 0 9 2 2
11 0 9 2 0 9 2 0 9 7 9 2
19 7 3 4 15 0 9 13 3 3 0 3 2 3 13 3 3 10 9 2
12 3 4 10 0 13 9 7 13 9 1 9 2
20 0 9 13 1 2 16 3 13 0 9 1 13 9 2 7 3 13 10 9 2
4 9 8 12 9
20 2 3 13 15 6 2 13 9 1 9 7 13 10 0 9 1 9 1 9 2
20 7 3 13 3 3 9 1 2 16 15 4 13 3 1 9 9 1 10 9 2
6 8 5 11 9 5 11
20 16 15 13 9 2 3 4 15 3 4 15 2 15 4 13 1 0 9 3 2
59 10 0 13 9 10 9 1 9 2 10 0 9 2 10 9 1 9 2 4 9 13 9 1 14 13 10 9 2 2 2 1 9 1 12 9 1 9 9 1 9 13 9 2 16 15 3 4 4 0 1 9 14 13 10 0 9 2 2 2
14 15 13 3 1 15 1 9 2 7 15 13 3 15 2
24 10 0 9 2 15 3 3 13 1 9 1 10 0 9 2 4 3 3 0 1 10 0 9 2
50 9 2 10 0 0 9 11 11 9 1 9 1 10 13 9 1 15 2 3 3 4 11 2 4 3 13 3 1 0 9 1 9 1 0 9 2 9 1 11 2 11 9 1 10 0 2 3 13 9 2
9 13 12 9 9 7 13 15 3 2
11 9 3 13 9 3 1 10 9 2 9 2
41 2 13 3 7 13 3 2 2 2 13 1 0 9 1 11 2 3 10 3 12 9 1 1 9 4 13 1 9 12 12 12 12 7 13 9 1 10 9 0 9 2
19 9 4 9 1 0 0 9 2 7 15 4 3 13 9 2 9 7 9 2
27 9 1 9 13 1 2 16 10 9 13 1 10 0 9 2 15 13 2 16 15 13 13 1 9 1 11 2
21 9 4 3 0 1 9 1 10 3 0 9 2 7 3 3 13 9 1 0 9 2
25 1 0 11 11 13 15 1 14 13 10 9 7 13 9 1 9 2 2 16 15 4 3 3 2 2
26 15 15 13 2 13 15 3 3 1 2 7 3 13 3 9 1 9 2 15 13 9 1 10 0 9 2
8 15 13 3 7 13 10 9 2
21 15 4 13 0 2 15 15 4 13 0 9 2 3 1 15 13 15 3 3 3 2
30 9 1 10 12 9 2 13 1 9 11 11 2 15 1 12 4 13 12 9 9 7 11 11 2 9 7 9 1 11 2
17 10 9 2 1 3 3 4 1 9 1 10 3 13 9 7 9 2
2 12 9
18 10 13 7 0 9 1 9 13 2 16 10 9 1 15 4 3 0 2
17 9 4 3 13 1 9 2 7 3 13 9 14 13 3 1 15 2
30 1 0 7 0 9 4 10 0 9 13 10 0 9 9 2 15 1 10 3 13 9 4 13 10 3 0 7 0 9 2
13 15 13 3 2 16 15 13 3 2 15 13 15 2
2 10 9
12 2 15 13 1 9 2 15 13 15 3 0 2
24 3 3 1 8 7 9 2 15 13 3 8 1 9 2 4 9 13 8 1 0 9 1 9 2
22 1 9 1 11 11 1 9 13 15 2 16 9 9 1 9 1 0 9 3 4 0 2
38 9 4 3 4 0 2 7 15 4 2 3 2 3 0 9 2 15 3 13 10 0 9 1 9 1 9 7 9 7 10 0 9 2 9 13 1 9 2
13 15 13 16 3 0 13 9 1 14 13 10 9 2
12 11 13 3 1 9 2 15 13 3 1 9 2
50 3 4 15 4 10 3 0 9 2 15 13 15 11 1 0 9 7 9 1 3 10 0 9 2 15 15 13 1 10 0 9 0 9 11 11 11 7 11 11 11 7 10 0 9 11 11 7 11 11 2
57 3 13 3 9 1 0 9 1 9 2 16 9 4 13 2 1 10 3 0 9 13 9 9 3 1 9 2 3 10 3 0 9 13 2 16 9 1 10 3 0 9 13 3 3 1 9 1 9 2 3 3 3 13 3 0 9 2
10 2 15 4 3 13 1 14 4 13 2
24 15 4 3 3 3 2 16 15 13 3 1 9 2 7 1 9 4 9 1 9 3 3 0 2
44 2 16 15 3 4 13 9 1 15 1 9 2 16 15 4 3 0 1 10 0 9 2 3 4 15 0 2 16 3 4 15 3 13 10 0 9 2 16 15 4 13 14 13 2
20 3 13 10 0 9 1 2 3 10 9 13 2 3 3 3 2 7 3 3 2
14 16 15 13 10 9 2 13 15 2 16 3 13 15 2
12 13 15 10 0 9 1 2 3 15 4 13 2
21 15 4 3 0 14 13 1 13 9 1 14 13 9 7 0 1 10 3 0 9 2
6 9 13 1 12 9 2
6 15 4 12 9 3 2
6 9 13 12 1 11 2
17 9 3 4 15 9 1 11 2 7 3 4 15 13 10 9 2 2
18 7 15 4 13 9 1 10 9 1 9 1 12 0 9 15 0 9 2
33 9 13 1 11 10 9 1 9 1 9 7 1 0 9 1 14 13 2 16 15 13 10 9 2 15 13 3 12 9 3 1 9 2
34 10 0 9 13 15 2 2 10 0 13 2 7 9 13 3 2 2 10 10 9 2 2 10 0 13 1 15 2 7 13 15 15 2 2
31 0 9 13 1 9 1 12 1 9 1 9 12 1 11 2 3 15 3 1 9 7 3 13 1 9 1 0 2 0 9 2
6 2 6 6 2 3 2
22 10 0 9 2 15 13 3 1 9 7 1 9 7 13 1 14 13 1 9 1 0 2
15 9 13 1 9 1 0 0 9 2 3 10 0 9 13 2
12 2 1 9 1 16 9 3 13 3 1 9 2
6 11 13 10 9 13 2
15 11 4 15 1 10 0 2 0 9 2 15 3 4 8 2
4 10 0 13 2
26 9 1 3 13 3 1 2 16 9 9 3 13 14 13 9 1 2 16 10 0 9 4 13 1 9 2
17 15 4 4 11 7 11 2 15 3 13 2 1 2 9 9 2 2
12 13 3 10 3 0 2 15 15 13 1 9 2
25 2 1 15 13 15 15 13 9 2 9 2 9 2 9 7 9 2 7 3 9 4 13 1 9 2
12 10 9 4 13 3 7 13 3 3 3 9 2
5 2 6 2 15 2
6 2 15 4 3 0 2
38 11 9 4 3 3 3 13 10 0 9 1 2 2 2 16 15 4 13 10 0 3 7 10 0 1 10 0 9 2 7 15 4 3 13 0 3 2 2
32 3 4 15 13 3 1 9 2 16 15 13 10 0 9 2 0 2 7 3 3 13 2 16 2 9 3 13 9 1 9 2 2
46 15 13 3 1 9 2 7 1 10 9 13 15 3 2 2 13 11 11 11 2 7 11 11 11 13 10 0 9 1 2 9 2 2 10 9 2 15 9 13 3 1 14 13 9 3 2
11 9 13 0 9 1 10 0 9 0 9 2
12 7 9 4 4 3 3 0 2 13 11 11 2
9 11 11 4 10 0 7 0 9 2
18 15 2 15 13 1 11 2 13 10 9 1 11 1 11 1 12 9 2
23 11 9 13 3 2 3 1 15 4 13 3 1 9 1 10 0 9 2 7 15 3 13 2
17 2 6 2 11 13 3 10 0 9 2 7 3 4 15 3 13 2
9 9 2 0 9 3 7 9 3 2
19 15 4 3 15 15 13 15 1 1 9 0 9 2 3 11 11 13 9 2
6 9 1 12 9 9 2
15 15 4 10 9 1 9 2 7 15 13 1 10 0 9 2
4 2 12 9 2
10 7 15 13 1 0 10 3 0 9 2
12 15 13 1 0 9 2 15 13 7 13 15 2
37 15 4 3 13 15 2 16 15 4 10 0 9 14 13 13 9 2 16 11 3 13 1 9 3 1 10 9 2 2 13 8 11 11 2 11 9 2
1 9
23 9 2 15 4 13 1 9 2 13 9 12 2 4 3 13 1 9 2 16 9 9 13 2
18 2 15 4 3 13 3 1 10 9 12 9 1 2 16 15 4 13 2
25 15 13 15 1 14 13 1 9 2 7 3 9 2 7 13 10 9 1 9 1 10 10 0 9 2
26 15 13 9 7 9 1 15 7 4 3 0 1 14 4 13 3 1 9 2 3 3 13 9 1 15 2
10 2 3 4 15 13 9 1 10 9 2
10 16 15 4 9 2 13 15 10 9 2
15 2 15 13 9 1 9 2 7 3 4 15 13 9 15 2
20 2 15 4 3 0 1 10 0 0 9 2 3 1 10 9 4 10 0 9 2
14 11 9 9 13 9 2 15 13 11 11 1 10 9 2
11 3 1 9 13 15 9 1 15 14 13 2
5 13 1 2 9 2
15 13 15 3 2 13 10 0 9 2 7 3 13 15 15 2
13 3 10 9 2 15 13 10 0 9 1 10 9 2
37 16 9 1 9 7 9 1 9 7 9 13 3 9 3 2 13 3 0 9 1 9 2 16 9 1 9 1 0 9 13 14 13 9 1 0 9 2
4 9 2 11 11
24 3 13 15 9 2 7 15 15 3 13 2 1 11 9 2 15 4 13 12 0 9 1 9 2
31 0 9 13 3 3 1 9 1 2 9 2 2 16 9 13 15 1 0 2 16 9 3 7 3 4 13 1 9 1 9 2
10 15 13 3 7 13 3 1 9 3 2
7 3 0 9 13 3 13 2
11 15 2 15 13 1 9 2 4 10 9 2
6 13 1 10 0 9 2
17 3 13 15 3 1 9 1 10 0 11 2 11 11 1 12 9 2
14 1 10 9 13 15 12 9 1 0 2 13 15 2 2
10 9 13 3 3 1 14 13 0 1 2
22 10 0 9 9 4 13 10 0 9 1 2 3 0 9 1 10 0 9 3 4 13 2
53 9 4 2 12 9 9 2 12 9 9 2 12 9 9 1 8 2 12 0 9 2 10 9 9 2 12 9 9 2 12 0 9 1 9 2 12 9 0 9 2 12 9 0 9 2 12 9 9 7 9 7 9 2
17 15 13 3 1 9 7 9 2 3 9 7 9 1 9 4 13 2
31 15 13 3 1 11 11 11 9 2 16 10 0 9 3 4 13 3 7 13 0 9 7 9 2 15 4 13 1 0 9 2
21 9 13 8 7 13 1 10 12 5 9 1 9 10 9 3 1 3 3 12 9 2
11 15 13 3 1 9 2 16 3 13 9 2
6 15 13 15 3 3 2
10 9 13 3 1 9 2 9 7 9 2
4 2 3 0 2
33 1 9 1 9 1 9 1 0 9 1 11 4 11 3 13 12 9 1 11 2 7 1 15 4 10 0 9 13 13 12 1 9 2
10 2 15 13 15 1 3 14 13 15 2
5 3 13 15 3 2
50 15 13 3 3 13 2 7 11 4 3 10 9 1 0 1 10 9 2 1 10 9 13 9 15 13 1 9 2 16 3 10 9 4 13 2 16 15 3 4 4 11 13 1 3 3 1 15 1 9 2
12 3 2 16 9 3 13 3 1 0 0 9 2
9 15 4 0 14 4 0 1 0 2
26 6 2 15 13 1 9 1 11 1 10 9 1 0 9 12 2 16 10 0 3 4 13 3 1 9 2
40 15 4 10 0 9 13 1 10 0 9 7 13 15 0 2 16 11 3 4 13 1 14 13 3 12 9 3 1 11 7 3 1 11 7 10 1 11 13 9 2
9 15 4 4 9 1 10 8 9 2
10 13 3 9 3 3 2 16 9 13 2
38 10 9 11 11 2 9 1 9 2 13 2 16 11 4 3 0 2 16 15 4 13 1 14 13 3 3 1 9 2 13 10 9 9 7 3 13 3 2
30 3 4 15 13 10 0 9 9 1 10 0 0 9 1 9 7 9 1 9 11 2 0 9 2 9 7 10 0 0 2
17 15 13 10 9 3 1 9 7 13 10 13 9 1 11 1 11 2
25 2 15 4 15 2 13 15 2 7 3 4 15 3 13 2 16 15 13 3 1 10 9 1 9 2
9 3 1 9 7 9 4 9 0 2
19 2 15 13 10 0 9 1 2 16 9 4 13 1 0 2 2 13 15 2
16 0 9 13 1 12 9 1 9 2 9 1 12 9 1 9 2
46 2 16 10 0 9 2 11 7 0 9 3 3 13 9 1 10 9 2 15 4 13 1 0 2 0 0 9 2 3 13 10 12 9 15 10 0 9 1 10 9 2 2 13 11 11 2
26 7 11 13 10 3 0 9 1 13 1 9 2 7 9 13 2 16 11 7 11 1 9 13 1 9 2
6 9 1 15 4 9 2
30 9 13 10 0 2 0 9 1 11 1 14 13 2 16 2 15 13 3 13 1 10 0 9 1 1 10 0 9 2 2
15 11 11 9 13 3 9 11 11 10 0 9 2 3 9 2
36 11 13 3 1 10 0 0 9 1 0 9 2 1 3 1 15 1 9 1 0 9 1 10 9 0 7 0 9 11 11 1 10 3 13 9 2
18 2 9 13 2 16 9 4 13 10 9 0 1 15 2 2 13 15 2
12 2 7 15 13 3 14 13 3 10 0 9 2
26 16 15 13 2 16 15 13 0 3 2 13 15 3 14 13 9 3 3 3 2 16 15 3 13 3 2
30 7 9 4 3 3 3 0 1 9 1 3 2 7 15 4 0 14 13 2 3 0 3 1 9 13 15 3 1 11 2
18 1 9 2 13 15 2 4 10 13 9 0 1 10 0 9 1 9 2
11 10 0 13 7 15 15 4 0 1 9 2
21 13 15 1 9 1 0 9 2 13 10 0 9 12 9 0 9 1 1 0 9 2
7 3 13 10 9 1 9 2
35 3 13 15 14 13 9 3 1 3 10 9 2 3 1 2 16 3 1 0 9 2 3 1 12 2 13 1 9 1 8 3 12 9 9 2
21 0 9 1 9 13 13 2 7 15 13 3 1 10 9 1 14 13 0 0 9 2
81 7 9 4 3 0 2 9 4 13 9 2 15 4 13 9 2 9 2 9 2 9 2 0 9 1 10 9 13 2 7 15 4 0 9 3 13 2 7 3 4 15 3 0 16 1 10 0 9 7 9 13 3 3 10 9 1 7 1 0 9 7 0 9 2 7 3 3 13 0 9 16 9 3 13 1 16 0 9 13 9 2
20 1 9 13 15 3 2 9 7 9 4 13 3 3 3 2 16 15 13 9 2
6 7 15 13 15 3 2
45 15 13 2 16 9 0 9 7 13 9 4 13 9 1 14 13 1 10 9 2 2 7 16 9 3 13 14 13 15 9 1 0 9 2 13 10 0 10 9 14 13 1 9 2 2
23 9 1 9 13 10 0 9 2 7 15 3 13 1 2 16 15 4 0 1 14 13 9 2
6 9 7 9 2 6 2
23 9 1 9 2 11 11 2 13 0 7 13 1 9 1 10 12 9 9 0 9 1 9 2
12 9 7 9 4 4 3 3 12 9 1 9 2
33 11 11 13 10 9 1 13 9 1 12 9 2 3 13 10 9 1 9 1 15 12 13 1 0 9 1 10 0 9 1 11 9 2
46 11 11 4 13 9 1 9 11 11 2 7 1 9 1 9 11 11 2 2 15 13 12 2 12 2 7 4 3 3 1 10 9 2 3 12 7 12 2 16 15 13 10 9 1 9 2
7 11 13 9 1 9 9 2
21 13 15 1 9 1 11 13 9 1 10 0 2 0 9 3 14 4 3 3 0 2
25 10 0 13 9 4 3 13 15 2 16 11 1 9 3 13 2 16 9 1 9 4 13 1 9 2
22 2 15 2 2 13 15 1 1 10 9 2 2 13 15 3 9 2 16 15 4 9 2
11 10 0 9 1 11 13 0 9 1 9 2
7 9 13 1 10 0 9 2
5 9 1 12 9 2
3 3 0 9
10 3 1 10 9 0 9 13 11 3 2
1 9
1 9
13 15 4 3 13 0 1 10 3 0 9 1 9 2
16 3 13 9 1 10 9 2 15 13 1 9 1 9 0 9 2
21 15 13 10 0 9 3 1 10 9 2 1 15 3 13 2 15 4 13 3 1 2
21 9 4 3 13 9 11 2 1 1 0 9 4 9 1 10 9 1 10 0 11 2
12 10 9 3 10 8 9 3 4 4 8 0 2
21 10 0 13 1 16 10 9 7 15 13 1 9 1 11 2 15 1 10 9 9 2
9 3 13 3 15 14 13 1 2 2
31 3 4 9 2 9 7 9 13 16 9 4 13 3 1 9 1 14 13 13 10 9 2 15 3 13 3 1 10 13 9 2
37 3 4 3 1 10 9 13 10 9 1 14 4 13 11 1 11 7 11 2 3 16 9 1 10 9 1 0 9 13 10 0 2 0 2 0 9 2
17 11 4 13 2 15 3 13 10 12 9 1 9 2 7 1 9 2
37 3 1 10 0 9 7 9 4 13 15 3 3 1 9 2 3 4 10 0 0 9 2 1 3 4 10 9 1 9 2 13 0 9 1 0 9 2
20 15 4 13 2 16 3 1 0 9 9 13 10 9 1 10 0 9 1 9 2
17 7 1 10 9 1 11 13 15 1 2 14 13 10 9 1 9 2
17 3 4 15 13 2 1 9 11 13 2 2 15 13 15 1 15 2
17 9 4 4 13 1 9 1 0 9 7 4 13 10 9 1 9 2
8 2 6 2 13 15 1 13 2
29 11 4 13 3 3 1 10 3 0 2 0 9 2 15 3 4 3 1 14 13 15 2 7 15 13 0 15 1 2
25 11 11 2 15 13 1 9 2 9 2 1 9 2 4 13 10 9 3 4 15 3 0 1 11 2
11 9 1 9 13 3 1 9 3 1 9 2
26 15 4 3 3 0 14 13 10 3 0 9 9 2 16 0 9 4 4 13 1 9 2 16 9 13 2
31 2 9 13 3 2 16 9 4 13 3 7 2 16 0 9 3 4 13 1 9 2 2 13 9 11 11 1 9 1 11 2
14 3 0 4 15 2 16 9 1 9 4 13 0 9 2
2 9 9
15 0 14 13 2 16 15 13 1 10 8 7 10 0 9 2
10 15 13 1 14 4 13 10 0 9 2
10 10 9 3 1 9 13 10 0 9 2
26 1 9 13 3 10 0 9 1 10 9 9 2 11 2 15 3 3 1 10 9 13 1 10 0 9 2
49 3 13 9 1 0 1 15 2 7 15 13 3 10 0 9 2 3 3 1 15 13 0 11 11 2 15 4 13 2 3 1 9 2 7 3 0 2 1 15 13 9 1 10 9 1 10 0 9 2
12 7 15 4 13 1 2 16 15 4 13 15 2
35 7 3 13 15 3 10 9 2 3 11 7 11 13 9 1 14 13 0 0 8 7 9 3 1 9 1 10 0 9 2 2 13 11 11 2
35 9 4 4 9 2 3 9 13 15 1 12 3 3 0 9 1 11 2 11 7 10 0 0 9 1 9 2 10 0 9 11 11 1 11 2
44 10 0 9 13 12 9 10 0 9 7 13 15 9 1 10 9 2 3 12 13 9 2 1 15 12 2 15 9 1 9 4 13 1 9 9 2 13 1 12 1 9 12 9 2
18 2 7 15 4 3 10 0 2 15 15 4 13 9 3 1 10 9 2
19 2 15 13 2 15 4 0 2 16 11 11 13 10 0 9 1 10 9 2
11 2 15 8 2 13 8 9 7 8 9 2
16 9 4 4 3 0 2 7 3 4 15 9 3 4 4 0 2
21 15 13 2 15 4 15 3 2 11 4 13 2 15 4 13 2 15 4 0 2 2
3 0 9 2
16 1 9 4 15 3 7 13 3 1 9 1 9 1 10 9 2
10 3 3 0 7 0 4 9 3 3 2
20 1 9 13 2 16 16 10 9 13 12 9 2 4 9 13 9 1 10 9 2
15 10 9 1 9 9 13 9 4 13 1 10 0 9 12 2
25 10 0 2 13 9 4 13 2 16 15 13 10 9 3 1 15 7 13 15 3 1 10 0 9 2
25 2 3 4 15 9 2 2 13 9 1 2 9 9 7 9 2 2 16 15 13 1 10 0 9 2
25 1 9 9 13 15 9 1 0 13 9 2 7 10 0 4 13 13 10 9 1 0 9 1 9 2
40 15 4 13 10 10 9 13 10 9 7 13 2 16 3 15 13 2 16 15 13 1 10 9 2 15 4 13 1 9 3 1 9 1 9 2 2 13 11 11 2
6 3 4 3 13 9 2
3 9 1 9
8 3 13 15 10 0 12 9 2
11 7 3 4 15 1 9 13 15 1 9 2
18 3 13 0 2 0 9 1 1 10 9 2 2 13 10 0 9 13 2
20 2 15 13 3 3 1 15 1 15 2 15 13 1 9 3 2 13 15 15 2
21 0 9 1 15 1 11 9 13 10 9 14 13 9 1 9 1 9 1 9 9 2
13 1 15 4 15 13 10 0 9 1 9 1 9 2
17 15 13 2 15 4 3 0 2 16 15 3 13 1 9 1 9 2
43 2 15 13 3 9 2 15 4 0 2 15 13 15 3 3 1 9 2 3 1 15 4 0 2 16 15 13 15 2 15 13 2 3 1 15 4 10 9 1 10 9 2 2
10 15 13 9 7 9 7 13 9 3 2
16 10 0 9 1 3 12 9 4 13 10 0 9 1 10 9 2
10 2 1 3 13 10 9 2 13 15 2
19 3 11 0 0 9 1 7 1 11 11 4 13 13 1 10 3 0 9 2
23 3 1 10 8 8 9 2 11 2 12 9 2 11 2 12 9 2 7 11 2 12 9 2
46 16 9 3 13 1 9 2 4 15 10 9 1 2 16 15 4 9 7 9 2 15 13 15 2 7 9 3 4 10 9 0 2 16 15 3 4 10 9 1 15 1 10 9 1 15 2
10 2 6 2 10 9 2 2 13 15 2
44 1 11 3 4 15 9 9 3 3 1 9 2 16 15 13 2 13 1 9 2 9 13 1 9 1 9 1 10 13 9 2 7 9 13 13 1 10 3 0 1 0 2 9 2
19 2 9 3 1 0 2 2 13 10 0 9 11 11 1 9 1 9 11 2
16 9 2 15 4 13 1 9 9 2 4 10 0 9 1 9 2
10 7 3 4 15 13 10 9 13 9 2
28 1 0 9 4 0 9 1 0 9 13 1 10 9 2 7 10 0 13 0 9 13 1 11 11 7 11 11 2
47 1 9 12 4 11 0 1 10 9 2 7 4 3 13 10 9 1 9 2 7 1 10 0 9 2 1 9 1 10 9 2 13 15 3 9 1 10 0 9 1 10 7 12 9 1 9 2
11 3 1 9 1 9 13 10 9 1 9 2
18 15 13 15 3 2 7 15 13 0 9 1 15 14 13 3 14 13 2
16 7 15 4 13 2 15 4 10 9 2 15 3 4 13 1 2
9 15 13 9 1 15 7 13 9 2
31 10 0 9 13 3 1 9 2 15 4 13 12 1 12 9 9 1 10 9 1 11 7 11 12 0 9 1 10 0 9 2
13 9 2 9 2 12 8 2 12 9 1 12 8 2
18 1 9 4 9 13 9 0 9 1 9 1 9 7 1 9 1 0 9
2 13 9
31 1 10 9 4 15 13 2 16 15 1 0 9 4 9 11 11 2 15 13 3 1 9 7 13 0 9 1 10 13 9 2
22 1 12 9 7 0 4 4 13 1 9 2 13 11 2 7 9 4 3 3 4 13 2
21 2 15 13 3 2 15 4 13 10 0 9 1 2 16 9 4 13 1 10 9 2
20 15 4 4 9 1 10 15 1 3 0 9 2 9 2 0 9 7 13 9 2
8 9 7 9 4 4 13 3 2
4 9 1 9 9
7 15 4 0 9 1 9 2
10 7 15 4 0 14 13 15 1 9 2
21 0 9 13 14 13 9 1 9 7 1 14 13 15 15 9 1 14 13 1 9 2
22 15 13 2 16 3 15 4 13 10 9 1 14 4 3 1 15 2 3 4 0 0 2
8 9 9 4 15 3 3 13 2
23 15 4 3 0 2 16 11 13 9 1 9 1 9 2 15 3 13 9 1 9 0 9 2
6 15 13 15 3 3 2
15 9 11 11 11 2 0 2 4 13 2 16 9 4 13 2
12 2 6 2 15 4 3 1 2 11 11 2 2
25 2 3 13 15 12 9 3 1 9 7 13 15 2 3 1 15 4 0 7 0 2 15 15 13 2
52 15 13 15 3 1 12 9 1 3 0 1 12 9 13 1 10 12 9 9 1 1 12 0 9 2 10 9 2 10 0 9 1 0 10 9 2 15 4 3 1 1 9 2 9 7 9 2 10 3 0 9 2
6 9 4 3 10 9 2
12 2 11 4 3 0 2 16 15 4 15 13 2
11 1 8 4 3 15 2 13 3 3 9 2
21 2 15 4 13 10 9 3 1 11 2 13 11 2 16 15 4 13 3 1 9 2
16 1 9 13 11 1 9 1 0 9 9 1 9 1 12 9 2
4 4 15 0 2
13 2 10 9 13 3 1 9 1 14 13 15 0 2
30 10 0 4 1 3 14 4 0 13 10 0 9 1 9 2 7 1 3 10 3 0 9 4 3 13 10 9 1 9 2
8 9 13 3 3 3 1 9 2
18 2 15 4 11 2 15 4 13 1 11 11 2 16 13 11 1 15 2
21 9 1 0 11 2 11 1 11 2 11 2 11 2 0 11 2 11 2 9 7 9
19 15 4 10 0 2 15 13 1 2 16 11 7 10 9 4 13 10 9 2
26 10 0 9 2 11 7 0 9 3 3 13 9 1 10 9 2 15 4 13 1 0 2 0 0 9 2
23 2 6 2 11 2 13 2 9 2 15 4 3 3 13 0 9 1 9 1 10 0 9 2
14 10 9 1 3 13 3 1 11 11 2 13 11 11 2
29 13 4 15 3 4 1 11 1 16 9 3 9 4 13 1 9 1 9 1 9 9 2 16 15 4 13 1 9 2
12 15 4 3 3 13 1 2 15 3 13 9 2
13 13 0 9 2 13 3 3 12 9 1 0 9 2
2 11 12
4 9 13 2 2
5 9 4 3 0 2
4 2 0 9 2
34 13 11 14 13 15 1 9 2 13 10 0 9 3 1 14 13 10 9 1 9 1 11 7 10 9 2 15 4 1 9 1 0 9 2
38 15 13 14 13 1 11 7 13 9 1 3 11 11 11 2 3 11 11 11 2 3 11 7 11 11 2 15 9 15 13 7 13 2 7 11 11 11 2
3 9 3 2
25 10 0 9 1 10 0 9 13 1 10 0 9 2 16 3 4 4 13 0 9 1 9 1 11 2
18 0 2 9 7 11 11 2 15 13 0 15 3 1 14 13 10 9 2
11 15 4 3 0 14 13 3 1 10 9 2
2 9 0
20 2 1 10 9 3 2 13 15 13 2 1 4 15 13 10 9 1 10 9 2
5 0 9 13 3 2
38 2 15 13 2 16 0 3 13 1 15 4 13 2 13 15 2 2 3 13 15 3 1 9 2 15 3 3 4 13 10 9 4 13 3 1 9 3 2
18 2 16 3 13 9 1 12 9 7 12 9 4 3 1 3 3 0 2
12 3 13 15 12 9 1 10 9 1 12 9 2
18 15 13 2 15 13 0 13 2 2 13 10 9 1 9 2 11 11 2
17 13 9 3 0 1 10 9 2 13 10 0 7 0 3 3 0 2
11 13 3 1 9 1 10 0 11 11 9 2
3 2 3 2
22 15 13 15 14 13 2 16 15 3 13 15 1 9 2 15 13 3 10 9 1 15 2
15 11 4 0 9 2 15 15 9 13 11 3 1 10 9 2
22 15 4 3 4 2 15 3 13 12 9 2 7 3 13 1 10 9 15 3 2 12 2
6 9 13 10 0 9 2
16 15 13 2 16 9 1 11 13 3 3 2 16 15 13 9 2
15 15 13 15 3 2 16 10 0 4 10 0 1 9 9 2
13 11 11 2 0 9 2 4 13 9 9 1 9 2
18 9 1 3 9 4 15 13 1 0 9 7 3 13 2 3 9 13 2
9 10 0 9 4 3 13 1 9 2
13 0 9 4 13 3 3 1 10 0 9 1 9 2
16 2 15 4 3 13 11 11 11 9 2 16 15 4 13 9 2
2 9 2
15 15 4 3 13 10 9 7 9 3 1 9 1 0 9 2
34 10 9 4 3 4 10 0 9 1 9 0 9 11 7 11 2 7 9 13 14 13 9 1 14 13 9 1 0 9 2 10 0 9 2
18 3 1 9 1 0 10 10 9 4 15 1 10 0 9 13 11 9 2
21 15 13 15 1 10 9 2 16 0 9 13 1 9 4 4 10 0 9 1 9 2
8 4 0 1 14 4 10 0 2
18 13 9 1 9 9 13 12 9 1 9 2 7 3 4 15 3 0 2
18 1 9 4 15 0 1 2 16 15 2 9 2 9 2 4 3 0 2
28 3 4 15 3 0 1 9 2 7 15 4 3 13 2 15 4 13 2 9 2 1 15 1 9 7 1 9 2
28 9 4 9 2 2 11 11 11 11 1 9 2 11 11 7 11 11 2 2 7 15 13 15 3 1 11 11 2
8 1 10 0 13 9 1 9 2
23 15 13 15 3 1 14 4 13 2 7 15 13 3 3 3 1 0 15 13 1 9 2 2
7 13 3 9 10 9 3 2
17 15 13 11 11 1 11 2 15 4 13 9 1 10 0 12 9 2
15 11 4 0 1 9 2 7 9 1 9 4 0 1 15 2
11 2 15 4 15 13 1 9 1 0 9 2
23 3 13 1 0 9 2 7 3 13 0 9 2 15 13 1 0 9 1 11 7 1 9 2
11 15 4 13 15 1 15 3 3 1 9 2
8 10 9 13 0 9 1 9 2
32 11 9 2 10 0 9 11 2 15 13 9 1 11 12 2 4 3 0 7 4 3 3 13 9 2 7 4 3 13 0 9 2
11 10 3 3 0 9 13 0 1 0 9 2
26 15 13 15 3 3 10 9 1 0 9 2 16 15 3 10 0 9 13 10 0 9 1 9 1 9 2
7 16 15 13 15 1 9 2
22 3 13 3 3 10 0 9 1 10 0 9 2 7 3 4 9 9 3 13 10 9 2
17 3 13 3 10 9 1 12 9 1 11 0 8 10 12 9 13 2
7 3 4 13 10 9 9 2
6 15 4 13 1 9 2
28 7 10 0 9 2 15 4 13 2 3 1 11 9 2 4 13 2 16 15 13 3 1 14 13 10 0 9 2
22 10 9 1 0 9 2 1 4 10 9 2 10 13 0 9 3 4 13 15 0 1 2
32 1 10 9 1 9 1 11 1 11 2 3 3 1 9 2 4 11 11 2 11 11 2 11 11 7 11 11 3 13 9 1 11
16 10 0 9 13 2 16 10 3 0 9 4 13 12 9 3 2
23 12 9 4 1 9 1 1 9 13 3 1 11 1 14 13 9 1 0 9 1 9 12 2
9 9 1 3 3 7 9 1 9 2
7 15 4 10 3 0 9 2
17 15 4 13 2 16 9 3 4 0 2 7 16 15 3 4 0 2
16 7 15 4 13 10 9 2 15 4 13 3 13 1 15 15 2
32 16 11 11 13 9 1 9 1 10 0 9 1 9 1 9 13 15 1 10 9 2 16 9 4 13 1 0 9 1 15 13 2
11 11 13 7 13 14 13 9 1 10 9 2
25 15 4 2 3 1 9 11 11 2 13 1 9 1 10 12 13 9 2 12 9 7 12 9 2 2
60 11 11 2 15 13 9 11 7 11 1 9 13 2 2 1 10 0 9 13 9 12 9 1 0 9 2 7 3 1 15 3 13 9 3 3 3 7 13 0 1 9 2 13 15 3 1 10 12 9 9 1 0 9 1 9 1 0 9 2 2
17 0 9 13 14 13 3 1 9 2 16 15 13 1 9 1 9 2
16 10 0 9 2 1 10 0 9 4 4 9 1 1 0 9 2
5 10 9 4 13 2
22 9 4 3 9 1 2 16 9 3 3 13 2 16 15 4 13 10 0 9 1 11 2
6 1 0 7 0 9 2
21 15 13 2 16 15 3 4 13 9 1 10 9 2 3 1 15 4 3 1 9 2
18 2 9 13 13 2 7 15 4 3 9 1 10 0 9 1 15 15 2
19 15 13 9 3 1 9 2 7 15 13 15 1 14 13 10 9 1 15 2
26 9 9 1 0 9 4 3 13 0 2 16 15 1 0 4 10 0 9 2 13 9 11 11 2 11 2
10 7 12 13 9 1 9 9 12 9 2
15 3 13 15 3 7 3 3 3 2 13 9 7 13 3 2
18 15 4 3 13 10 9 1 9 1 11 2 1 15 13 15 0 1 2
35 2 1 0 9 13 15 14 13 2 16 15 4 0 2 7 1 9 3 13 15 9 1 0 9 2 7 15 13 3 2 3 3 15 13 2
8 2 11 13 15 3 1 15 2
46 9 4 15 3 3 3 13 15 1 9 1 15 12 8 2 7 3 4 15 3 2 7 15 4 13 0 1 14 13 7 13 15 2 16 10 9 1 8 3 13 2 2 13 11 11 2
33 11 13 1 9 1 0 9 1 0 9 2 7 13 3 14 13 3 1 0 9 2 15 13 9 9 1 10 9 1 1 10 9 2
5 3 0 3 0 2
68 9 13 3 1 12 9 2 3 1 9 4 3 2 16 9 4 13 13 2 7 1 0 9 4 10 0 9 1 9 3 3 2 16 11 13 3 1 10 13 9 7 10 3 0 9 1 10 9 2 7 10 0 9 3 0 2 16 15 13 11 1 10 9 1 14 13 9 2
33 7 11 4 3 3 1 10 9 2 1 15 4 0 14 13 2 16 15 1 0 9 1 12 13 0 1 9 2 7 13 1 9 2
11 2 9 2 4 10 0 2 7 0 9 2
3 3 2 2
6 15 13 15 3 2 2
3 2 6 2
8 3 13 15 0 1 11 9 2
6 15 4 3 4 9 2
20 9 13 10 0 9 1 14 13 3 2 3 1 9 2 15 3 4 13 3 2
19 2 1 15 13 15 10 0 9 7 10 0 9 3 2 3 7 0 9 2
14 2 11 8 11 2 11 11 8 8 8 8 2 2 2
7 1 3 13 1 12 9 2
14 2 9 4 10 9 2 15 1 15 10 9 4 13 2
29 10 0 1 11 2 3 12 9 2 16 9 4 13 3 9 1 1 11 7 11 1 10 0 9 1 11 0 9 2
21 9 1 10 9 13 13 1 0 9 2 7 3 13 15 16 3 3 3 4 13 2
42 1 10 0 9 13 15 12 9 14 13 10 0 9 2 7 1 9 4 15 13 1 12 9 2 16 15 13 10 9 3 7 3 13 2 16 10 9 13 10 13 9 2
13 7 15 4 3 3 13 15 1 15 2 3 2 2
27 12 9 13 1 11 11 2 10 9 1 11 4 13 1 9 1 12 9 1 9 2 15 13 9 1 12 8
14 9 13 3 8 2 7 15 4 3 13 14 4 0 2
14 2 15 4 3 9 2 16 9 4 13 1 10 11 2
26 2 10 9 2 15 13 9 1 11 2 7 3 13 15 3 3 1 10 0 9 2 13 3 9 3 2
30 0 9 3 0 2 7 3 0 2 9 2 1 11 11 13 3 11 13 9 2 7 4 3 13 9 1 10 0 9 2
66 9 4 1 15 13 3 13 9 1 9 3 4 13 1 8 7 9 3 3 1 0 9 7 13 9 1 10 0 9 1 9 9 3 4 13 3 3 1 9 7 13 1 9 7 9 2 3 13 3 9 4 13 1 0 2 0 2 0 7 0 9 7 9 7 2 9
18 9 4 0 2 16 9 1 9 3 4 10 0 9 9 1 0 9 2
4 9 13 15 2
28 9 11 13 13 9 2 16 15 1 9 13 13 9 13 7 12 9 9 1 13 1 10 9 1 9 1 9 2
41 3 3 2 3 1 16 15 4 13 12 9 7 13 10 9 2 13 9 2 3 10 0 2 7 9 1 9 4 1 9 2 7 15 4 13 2 3 0 15 13 2
2 9 9
27 13 2 3 4 15 13 15 13 2 16 9 4 13 3 13 7 13 2 16 13 15 3 13 1 10 9 2
3 0 3 13
9 3 13 9 1 12 7 12 9 2
10 13 15 2 16 15 4 13 0 9 2
13 3 1 14 13 15 2 16 3 3 13 0 9 2
29 13 3 1 2 15 15 3 13 2 15 13 1 15 7 13 13 1 14 13 1 9 2 16 9 13 3 1 15 2
12 15 12 4 3 1 10 0 9 13 13 9 2
8 2 3 9 7 9 13 15 2
13 3 4 11 11 7 12 9 13 10 9 1 9 2
8 3 4 15 3 13 1 11 2
25 15 13 10 0 9 1 9 7 9 1 9 9 12 2 7 13 1 3 10 9 1 9 1 9 2
51 15 4 3 13 2 16 9 1 9 9 3 0 9 3 4 4 3 12 1 2 9 2 2 2 9 2 1 9 2 2 13 9 2 13 9 15 2 4 3 12 9 2 16 3 13 3 10 2 9 2 2
54 9 11 4 3 3 13 9 11 11 9 1 2 16 9 1 9 1 9 12 13 3 1 10 9 1 14 13 10 3 12 0 9 2 15 4 13 1 11 1 1 12 9 2 10 9 1 11 1 11 4 4 13 13 2
35 9 13 3 0 9 2 9 2 9 3 1 9 3 2 9 2 2 7 9 9 2 9 2 9 1 9 2 9 1 9 2 9 9 3 2
18 3 13 9 1 11 3 2 16 9 1 0 9 13 9 12 1 9 2
26 2 15 13 1 11 3 0 9 2 10 0 9 2 2 13 10 0 9 11 11 2 11 2 1 11 2
23 15 4 13 1 2 16 15 3 3 4 3 2 16 10 3 13 9 3 4 10 0 2 2
8 11 13 3 1 10 0 9 2
12 3 1 0 9 13 15 10 9 8 3 2 2
14 15 4 8 13 1 14 4 12 0 9 7 13 3 8
22 10 0 9 9 4 10 9 1 2 16 11 4 13 10 3 3 0 9 1 9 9 2
9 13 9 13 13 1 3 12 9 2
13 7 15 4 3 0 2 16 15 13 3 1 9 2
26 7 9 1 2 16 15 1 3 4 9 1 10 0 2 0 9 2 15 3 13 1 10 9 1 11 2
19 3 0 9 13 1 7 13 10 0 9 13 1 2 3 0 9 13 9 2
9 10 9 13 10 9 3 1 9 2
26 2 16 15 2 3 3 7 0 15 2 3 4 4 0 1 10 9 2 15 4 13 1 10 0 9 2
18 9 4 3 13 10 2 9 2 2 15 2 9 12 2 4 13 1 2
15 15 4 3 0 7 3 0 2 7 9 4 3 0 3 2
1 0
18 0 9 0 9 1 14 13 7 3 13 0 7 0 0 9 13 3 2
21 3 4 9 1 11 13 2 16 15 3 13 9 2 1 15 13 9 2 13 15 2
16 9 4 13 3 1 12 9 1 10 9 9 2 15 4 9 2
9 15 13 15 2 16 9 4 12 2
21 15 4 0 2 16 9 7 9 13 3 2 3 3 1 9 2 7 3 1 9 2
30 0 9 13 3 7 0 1 9 7 4 1 3 10 9 2 15 13 0 1 3 2 3 15 3 13 3 0 9 9 2
9 16 9 13 3 13 9 1 9 2
51 2 9 4 13 10 0 9 1 15 2 3 4 0 1 9 1 11 2 1 16 10 0 9 9 4 13 3 2 7 16 0 9 7 13 9 1 0 9 3 4 4 13 2 2 13 11 9 2 11 11 2
32 10 0 9 13 1 0 9 1 11 1 14 13 14 13 10 9 7 13 1 2 16 3 1 9 13 1 10 0 9 1 9 2
14 3 13 15 10 0 0 9 1 0 7 0 9 3 2
25 3 1 9 3 1 9 13 10 0 9 1 9 7 13 1 10 0 9 3 3 1 10 0 9 2
29 15 13 1 9 1 14 13 2 0 7 0 7 0 2 3 13 1 10 0 9 7 1 10 9 13 3 1 9 2
13 10 9 1 10 7 10 9 4 3 13 10 9 2
7 3 13 1 9 7 9 2
6 13 15 3 1 15 2
17 2 6 2 15 13 1 10 0 9 1 9 10 9 1 10 9 2
12 3 13 9 1 9 1 13 9 1 9 3 2
18 1 9 4 15 3 0 14 13 7 13 1 9 3 2 13 15 13 2
31 2 15 13 3 3 1 9 2 7 9 13 15 2 7 15 4 3 13 2 16 15 13 3 2 2 13 11 11 1 11 2
6 11 13 1 10 9 2
24 2 1 9 4 15 13 7 13 1 2 16 9 13 9 2 16 9 13 3 1 3 12 9 2
22 11 2 3 4 10 0 9 11 11 3 0 1 14 13 9 3 1 9 1 11 9 2
21 9 1 10 9 4 3 12 9 7 12 9 2 3 13 10 0 9 1 11 11 2
18 15 4 13 3 3 3 1 9 2 16 15 4 13 9 1 0 9 2
11 7 10 9 1 9 4 0 2 13 15 2
8 7 10 0 9 13 3 9 2
9 0 2 0 7 3 1 14 13 2
4 2 3 3 2
40 1 10 0 9 13 1 11 9 7 9 9 0 9 4 9 3 13 9 1 14 13 9 10 9 1 12 9 1 9 2 15 15 13 1 14 13 3 1 9 2
21 10 0 9 1 9 4 13 1 9 2 16 9 13 3 2 7 9 3 13 3 2
10 7 15 4 9 3 13 9 9 1 2
23 9 13 14 13 9 1 11 11 9 7 9 2 11 11 11 11 2 3 3 4 11 9 2
4 9 13 0 2
12 3 4 15 13 9 1 11 2 3 1 9 2
15 15 13 10 0 9 7 4 4 13 10 0 9 1 9 2
16 3 13 10 9 1 15 2 15 9 9 13 3 1 10 9 2
11 2 15 4 3 3 0 2 13 11 3 2
27 16 9 13 2 7 9 13 2 13 11 11 11 3 1 10 9 1 9 11 11 3 12 9 3 1 11 2
42 16 15 4 13 3 2 4 15 13 3 1 15 2 16 15 14 13 10 9 3 4 10 9 2 2 13 11 11 2 15 3 3 4 13 9 3 1 12 9 1 9 2
18 2 15 4 0 2 13 9 2 2 7 0 2 15 13 10 0 9 2
19 3 4 13 9 2 3 10 0 9 4 13 7 9 2 3 15 3 13 2
19 9 13 3 2 16 9 9 13 2 16 9 1 9 4 9 1 0 9 2
21 1 0 9 13 15 3 10 9 1 10 9 1 0 2 3 10 9 1 15 15 2
13 3 13 12 9 1 9 2 3 15 12 4 0 2
10 15 4 10 9 2 15 9 13 0 2
8 15 7 9 13 1 10 9 2
33 7 15 13 1 13 9 0 9 1 9 1 11 11 2 10 0 9 11 11 2 9 11 11 2 9 11 11 7 3 9 11 11 2
18 10 0 11 9 13 3 1 9 2 15 13 1 15 10 0 9 3 2
8 15 13 2 2 3 3 2 2
34 9 2 0 7 9 2 2 9 2 9 2 9 2 0 9 2 9 2 12 8 2 12 8 7 12 8 2 2 9 2 9 7 9 2
21 10 9 2 15 13 1 9 2 4 3 13 9 1 9 2 3 16 9 4 13 2
17 1 10 9 9 13 10 9 3 2 7 15 13 15 1 10 9 2
24 11 9 1 9 1 9 9 4 3 3 3 13 1 10 0 9 2 15 3 4 13 1 9 2
28 9 0 9 13 9 2 12 9 1 12 0 9 2 3 1 9 2 7 9 13 2 16 15 13 3 1 9 2
12 15 4 1 15 15 10 0 9 1 10 0 2
9 3 4 13 12 9 9 1 9 2
29 15 4 3 0 2 7 0 2 3 10 0 9 2 4 0 1 15 2 16 15 13 1 9 2 2 13 11 11 2
7 2 0 2 13 9 7 11
41 15 4 3 4 4 0 1 11 2 14 13 0 10 9 1 9 2 7 13 4 15 3 3 2 16 9 3 4 4 13 1 10 0 9 2 3 15 13 9 8 2
36 15 4 3 10 3 0 9 14 13 10 9 2 3 15 1 10 0 9 4 13 3 1 10 0 9 2 16 10 0 9 4 13 3 3 3 2
15 1 9 12 1 12 9 2 9 1 9 12 0 9 2 2
25 0 9 2 15 13 9 1 9 1 9 2 4 13 9 2 1 9 4 13 9 1 2 13 5 12
46 4 15 3 1 10 9 13 11 11 0 9 13 1 9 7 1 9 13 15 10 9 1 10 9 2 9 7 9 2 2 15 1 0 9 13 9 1 11 9 1 11 7 9 1 11 2
7 15 4 0 1 10 9 2
3 3 5 12
2 0 9
15 2 9 13 3 0 9 1 0 9 7 1 10 9 9 2
7 9 2 12 9 1 9 2
14 15 4 13 9 2 7 15 4 3 13 9 7 9 2
2 0 9
6 15 4 3 13 9 2
38 3 1 11 13 3 14 4 0 2 3 1 9 1 0 9 7 9 13 1 9 2 7 3 13 9 1 9 1 9 2 13 10 9 1 10 0 9 2
27 15 4 3 0 1 2 16 9 3 13 15 0 2 16 3 10 9 1 2 15 15 13 2 13 1 9 2
24 1 9 13 3 0 9 1 10 9 2 7 15 13 9 1 14 13 9 2 1 14 13 9 2
2 9 2
15 10 10 9 1 9 13 3 14 13 15 1 9 1 11 2
35 1 10 9 9 13 15 3 3 2 16 10 9 4 13 3 2 16 11 13 15 0 0 9 2 2 15 4 3 3 13 1 9 7 9 2
16 9 9 13 14 13 2 16 9 4 10 9 7 10 0 9 2
34 1 9 1 10 0 9 1 9 2 13 11 11 7 11 11 3 9 1 9 2 15 3 13 15 0 1 11 11 14 13 13 10 9 2
23 2 15 13 3 10 1 10 0 9 1 14 13 9 7 13 15 3 1 10 0 9 2 2
32 3 0 9 13 15 3 1 14 13 10 9 2 7 15 7 9 4 3 13 9 1 14 13 10 0 9 2 2 13 11 11 2
35 1 10 9 13 9 9 1 10 9 9 1 10 0 0 9 7 9 7 10 0 9 1 8 7 9 2 2 7 3 0 10 1 0 9 2
13 9 11 11 2 2 15 13 3 9 1 10 9 2
1 9
29 1 9 1 9 4 9 4 13 10 3 0 9 1 9 9 1 9 1 8 1 9 2 3 9 1 9 4 13 2
8 15 13 15 2 15 3 13 2
10 15 4 4 3 1 14 13 9 10 9
7 9 4 12 9 1 9 2
7 3 3 13 11 12 9 2
30 10 0 2 0 9 1 11 13 15 1 9 7 13 12 9 3 2 9 2 9 2 16 15 4 13 9 1 11 9 2
10 15 13 3 13 2 2 13 11 11 2
10 1 0 9 13 9 1 0 1 9 2
38 2 3 1 0 10 9 2 15 4 3 3 14 4 13 1 10 9 2 2 13 9 1 9 1 2 16 11 11 1 0 9 3 4 13 1 10 9 2
9 7 15 4 3 3 15 1 9 2
35 7 15 4 3 10 3 0 9 1 10 12 9 2 15 4 13 2 7 3 13 3 10 0 9 1 2 16 9 4 3 0 1 0 9 2
13 16 9 3 13 14 13 2 4 15 3 13 9 2
40 1 10 0 12 9 4 11 11 13 1 10 3 0 2 9 2 1 11 3 1 10 0 9 11 7 10 9 11 2 15 1 9 1 0 9 4 1 9 9 2
21 16 11 11 13 10 0 9 3 1 0 9 0 9 2 13 15 3 3 1 9 2
20 9 13 1 9 2 15 3 13 9 1 10 9 2 16 9 1 9 4 13 2
29 15 4 0 1 2 16 10 0 9 1 11 4 4 13 3 1 10 0 9 1 9 1 11 3 0 9 1 9 2
34 15 4 3 3 0 1 14 13 9 1 10 9 2 13 11 11 7 13 2 2 15 4 3 10 9 2 1 0 9 3 13 0 1 2
9 15 13 9 9 7 13 9 3 2
2 13 9
13 1 8 13 9 3 1 10 9 1 9 2 9 2
10 9 13 3 1 0 9 7 1 9 2
65 10 0 2 0 2 0 9 4 1 10 0 9 1 10 9 2 15 13 1 2 7 16 10 10 9 0 9 2 11 2 4 15 2 1 0 9 2 13 10 9 2 16 15 4 12 2 16 15 4 12 2 3 1 10 9 1 11 11 1 10 0 9 1 9 2
4 9 1 11 0
12 16 15 13 2 4 15 3 13 3 7 3 2
17 3 13 9 1 0 11 9 3 3 13 2 7 9 13 1 9 2
19 1 10 9 4 9 1 9 1 10 0 9 7 11 13 1 3 0 9 2
35 9 13 10 9 2 7 15 13 3 3 2 3 3 7 3 2 16 15 3 4 13 2 16 10 0 9 1 0 9 4 13 9 1 9 2
14 13 3 9 12 1 9 7 9 12 1 9 1 9 2
24 11 11 13 1 9 9 2 16 9 4 0 1 9 1 10 0 9 1 9 7 10 0 9 2
24 11 13 12 9 1 9 1 0 9 2 7 9 4 1 3 12 9 1 9 3 1 12 9 2
10 2 13 15 3 7 13 15 13 3 2
16 1 11 4 10 0 9 1 9 13 9 1 0 1 9 1 9
17 11 4 0 1 10 0 9 2 3 1 1 10 0 2 0 9 2
24 15 4 1 9 13 0 16 10 9 2 11 11 11 2 1 9 1 8 9 2 9 11 11 2
42 15 4 3 13 2 16 9 1 11 3 0 9 1 0 11 13 1 14 13 7 13 1 2 3 1 14 13 1 10 9 1 0 9 7 3 3 1 10 9 1 9 2
9 3 13 15 9 7 13 1 15 2
35 3 1 9 1 11 13 11 1 9 3 3 1 9 2 3 9 1 3 4 13 2 16 9 3 4 15 1 10 0 7 3 0 1 9 2
30 11 4 1 9 13 1 9 1 15 1 10 10 0 2 9 2 1 9 2 15 1 9 1 10 0 13 13 9 1 2
22 15 4 1 11 9 13 2 16 15 1 14 4 12 9 1 12 4 4 12 9 1 12
11 2 15 4 0 9 13 1 3 14 13 2
9 3 13 15 9 9 1 10 9 2
47 10 9 2 15 3 4 13 1 12 9 2 12 9 2 12 0 9 2 10 9 7 12 9 1 11 2 4 13 1 9 1 10 0 9 2 1 1 11 11 9 4 2 10 9 9 2 2
10 16 9 13 13 9 1 9 7 9 2
10 9 1 0 9 4 15 3 13 2 2
9 10 0 9 4 15 13 1 15 2
16 7 15 4 3 13 1 2 16 3 13 9 1 10 9 9 2
21 1 9 13 1 15 0 9 11 11 11 7 9 11 11 7 9 11 11 2 9 2
6 10 9 13 3 10 9
4 9 1 9 2
6 2 11 2 13 15 2
11 1 9 4 9 13 1 9 1 0 9 2
10 2 13 3 3 3 2 13 15 3 2
30 11 2 15 1 12 9 3 13 10 0 9 1 9 1 13 9 2 13 3 12 9 1 10 0 9 1 12 9 9 2
25 3 13 3 12 9 9 1 15 9 2 7 15 13 0 7 0 2 3 3 3 2 15 4 13 2
8 2 10 9 4 13 1 11 2
8 7 3 13 11 3 10 9 2
9 15 13 9 1 11 1 9 12 2
19 7 0 1 15 13 3 9 1 14 13 3 1 10 9 7 13 9 3 2
21 3 13 11 11 3 1 15 13 2 16 15 4 0 1 11 9 1 10 0 9 2
72 15 13 3 1 10 13 9 11 8 2 11 8 1 9 11 11 0 9 2 3 9 11 11 2 9 15 7 9 11 11 1 9 13 15 3 1 9 1 11 2 15 13 2 3 13 9 3 4 13 1 9 1 10 3 13 9 2 3 1 15 3 4 13 16 9 1 9 13 1 11 11 2
4 15 13 9 2
20 15 13 1 10 0 9 2 15 11 3 13 14 13 2 3 1 9 9 9 2
61 7 3 1 9 1 9 1 10 0 15 2 9 4 9 7 9 2 2 4 0 9 2 3 4 3 3 10 9 0 9 2 2 15 4 13 9 1 9 7 4 13 3 1 10 0 9 2 3 15 4 4 0 2 7 15 4 4 10 9 2 2
1 9
4 3 7 3 2
25 1 16 11 4 13 13 2 16 9 3 4 3 0 1 14 13 9 2 13 9 9 14 13 9 2
23 7 1 0 9 1 9 13 15 10 0 9 2 16 15 4 13 10 9 1 14 13 11 2
4 9 13 3 3
24 15 13 9 1 10 0 9 3 3 3 2 9 13 3 3 1 11 9 1 12 2 13 9 2
30 10 0 11 11 1 11 13 1 10 0 9 1 9 1 11 2 16 15 13 9 1 14 4 10 0 9 1 0 9 2
4 9 1 9 2
1 9
13 15 4 3 3 0 2 16 9 4 12 9 0 2
6 13 9 5 12 9 5
14 7 15 13 1 14 13 2 15 13 15 15 3 1 2
27 2 15 13 0 9 10 9 3 1 9 2 16 15 13 2 16 15 3 3 4 15 2 15 13 15 1 2
19 3 16 15 4 13 15 2 7 16 10 3 2 0 2 3 4 3 3 2
6 10 9 3 13 9 2
17 9 13 1 12 12 12 5 1 9 1 10 13 9 7 10 9 2
50 15 4 13 14 13 10 9 9 2 7 0 9 4 15 13 9 2 3 2 2 2 2 13 10 0 11 11 2 15 4 8 10 0 9 1 14 13 10 9 2 16 10 12 9 4 13 7 1 9 2
40 1 9 4 9 1 0 9 3 13 2 6 3 13 1 9 1 12 1 12 1 0 9 1 9 2 7 9 4 3 13 1 12 9 9 1 3 12 9 9 2
23 10 9 13 1 0 10 9 2 15 4 13 3 2 16 15 4 9 2 16 15 13 3 2
12 15 13 3 3 3 1 0 9 7 0 9 2
27 2 9 7 9 2 2 2 11 8 11 2 2 13 1 9 1 10 0 9 2 15 13 1 10 0 9 2
23 1 15 13 9 11 11 2 2 11 9 9 1 2 16 9 4 8 9 4 3 0 2 2
18 2 6 1 9 2 13 9 2 2 7 15 4 13 15 10 0 8 2
12 9 7 10 9 13 3 1 10 0 9 11 2
38 1 0 9 2 15 4 13 9 2 15 4 13 1 9 1 9 2 9 7 9 2 7 13 9 3 2 4 9 7 9 13 3 3 2 13 5 12 2
2 5 12
26 10 0 9 4 15 13 2 15 3 3 3 4 10 9 1 2 16 9 4 13 1 9 1 10 9 2
12 3 13 12 9 2 15 13 14 4 13 9 2
1 11
24 7 15 13 1 14 13 9 2 7 15 4 3 3 10 9 1 9 2 2 13 11 11 11 2
16 10 0 9 1 9 13 3 1 9 10 9 1 10 0 9 2
13 3 4 9 13 2 16 9 3 13 1 10 9 2
11 0 9 9 4 13 9 1 9 1 9 2
21 9 13 13 0 9 1 2 16 9 7 9 13 1 14 13 9 1 1 10 9 2
2 9 11
9 2 15 13 3 10 9 2 11 2
1 9
19 15 4 4 3 1 2 16 3 4 13 9 1 10 0 9 1 15 8 2
37 10 9 4 10 0 1 15 2 16 15 4 13 10 0 1 10 0 9 2 7 9 4 3 1 3 13 13 3 1 10 9 1 9 1 9 9 2
12 13 15 2 4 15 13 15 1 15 2 11 2
14 7 15 4 3 3 9 1 9 2 15 13 1 9 2
14 15 13 11 11 11 3 1 10 9 12 9 1 9 2
23 15 13 10 9 9 1 9 2 7 16 15 13 15 1 15 2 13 15 15 7 13 0 2
8 2 15 4 13 3 9 12 2
11 7 3 13 10 0 9 1 14 4 9 2
25 10 9 2 15 13 10 9 2 10 9 2 10 9 2 10 9 7 10 9 10 0 9 1 9 2
9 10 0 9 13 3 3 1 15 2
25 10 0 0 9 4 2 16 15 13 3 1 14 13 3 1 14 13 3 2 16 15 13 10 9 2
9 2 3 13 15 11 2 13 9 2
12 2 13 15 3 2 16 15 13 10 10 9 2
37 2 7 15 13 9 13 10 0 9 2 2 13 10 0 9 2 16 9 13 1 9 7 11 0 9 2 11 11 2 13 9 1 11 9 11 11 2
19 10 0 9 13 15 2 16 15 1 9 13 1 9 7 13 3 1 9 2
22 15 4 4 9 1 10 0 9 1 0 1 12 9 2 3 4 0 9 13 1 15 2
33 3 13 9 1 10 0 9 2 7 3 1 3 3 4 13 10 0 9 0 9 1 10 0 11 2 3 13 9 3 1 4 0 2
20 2 6 2 6 2 0 2 0 4 15 3 3 2 13 9 7 13 3 3 2
53 2 10 9 13 15 3 3 1 10 0 2 2 13 11 1 9 2 2 7 3 4 15 3 3 0 1 2 16 15 4 3 3 3 1 11 7 3 3 13 9 1 11 7 13 15 1 10 0 2 15 4 2 2
10 10 0 9 4 13 3 16 1 3 2
5 9 13 15 3 2
15 15 4 13 1 10 9 2 16 3 4 15 13 3 2 2
91 2 15 13 1 9 12 9 1 9 1 11 1 9 1 1 9 12 9 2 7 15 4 0 2 16 15 3 4 13 15 1 2 16 15 1 10 9 4 4 13 1 10 0 9 2 2 13 11 11 2 9 2 11 9 2 1 16 0 11 11 1 11 13 3 1 11 7 13 2 15 3 13 1 10 9 2 15 1 10 7 10 0 9 13 1 14 13 10 0 9 2
36 11 11 13 10 13 11 7 1 9 1 9 1 11 11 9 13 11 11 2 11 11 2 11 11 11 2 11 11 2 11 11 7 11 11 11 2
32 1 9 1 9 1 11 4 8 3 4 3 1 14 13 2 16 9 11 11 3 3 13 1 9 1 11 1 14 13 10 9 2
52 9 1 9 1 9 1 11 2 9 1 0 9 3 1 10 0 9 1 11 11 7 10 0 9 2 7 9 1 0 2 1 9 11 11 2 4 3 13 0 9 1 9 7 9 2 1 1 0 2 0 9 2
20 1 10 9 4 3 3 3 13 10 9 2 15 3 0 9 4 13 1 11 2
6 3 4 9 12 9 2
35 15 4 0 2 3 0 15 4 13 1 9 2 3 0 9 1 10 0 9 2 3 15 1 14 4 9 3 4 2 13 2 10 9 9 2
15 2 15 4 3 15 2 15 4 13 1 2 2 13 15 2
20 3 3 0 9 13 15 1 11 11 2 16 15 3 4 13 1 10 9 9 2
36 9 1 9 4 13 7 13 1 10 9 2 3 4 4 0 1 9 7 13 1 10 9 9 13 1 9 2 10 9 1 3 12 9 13 2 2
11 9 4 1 3 13 15 1 0 9 9 2
12 1 10 9 9 4 10 0 1 9 4 3 2
20 7 13 3 15 2 15 4 13 2 3 13 15 14 13 1 14 13 9 3 2
12 11 11 7 9 13 0 9 14 13 10 9 2
7 7 15 13 15 3 15 2
40 7 3 4 15 1 0 13 10 9 2 15 13 2 16 3 3 13 9 7 0 1 9 1 10 9 15 13 1 9 10 9 1 11 7 11 1 10 9 13 2
21 13 15 2 4 10 9 1 9 4 0 2 7 13 15 2 4 15 3 4 0 2
14 0 10 9 13 3 2 15 15 4 13 2 13 9 2
17 10 12 13 9 4 4 10 0 9 1 11 1 3 1 12 9 2
22 1 11 13 9 2 16 3 1 9 2 3 1 9 2 13 12 9 9 1 15 9 2
9 2 6 2 7 13 9 7 11 2
2 11 2
16 10 9 2 15 13 1 9 1 11 2 4 3 10 9 0 2
21 3 0 1 15 2 13 3 3 3 15 2 15 13 9 1 14 4 2 11 2 2
48 0 10 9 4 13 1 10 13 9 9 10 0 10 2 7 1 9 11 4 13 1 10 9 7 4 13 10 0 9 9 1 9 1 9 2 4 15 3 3 9 1 10 13 9 4 4 13 2
8 3 13 11 15 3 1 9 2
15 9 1 9 13 10 0 9 1 3 14 13 15 1 9 2
66 3 4 3 3 13 1 9 1 10 9 2 16 15 4 13 2 16 9 11 11 3 13 10 9 1 10 13 9 2 9 11 11 2 7 16 10 0 11 11 4 13 3 0 9 2 16 15 13 9 2 15 3 13 15 1 2 16 9 15 1 15 9 13 0 9 2
10 0 9 2 3 7 3 2 13 1 9
12 1 10 9 2 16 15 4 13 15 1 15 2
28 9 1 11 11 13 3 1 9 2 9 7 9 7 9 7 9 2 9 1 9 1 10 9 1 10 0 9 2
27 10 3 0 9 1 9 13 11 11 3 3 1 12 2 3 15 13 10 11 1 13 1 2 0 9 2 2
39 7 3 1 10 0 9 13 2 13 15 3 1 0 9 9 2 3 9 2 9 7 0 7 0 9 1 0 9 2 0 3 1 3 3 13 9 1 9 2
22 0 9 1 0 9 13 9 11 1 14 13 2 10 0 9 2 2 15 15 13 15 2
3 9 3 0
13 2 9 1 0 9 13 1 12 3 9 1 9 2
17 9 9 13 3 3 1 2 1 15 9 10 0 2 9 2 13 2
17 2 15 4 10 0 2 15 13 10 9 3 1 14 13 15 2 2
10 9 13 10 13 9 7 10 13 9 2
19 2 15 13 3 1 14 13 2 2 13 9 11 11 1 9 1 11 11 2
33 12 9 1 12 7 12 9 4 13 3 3 2 16 15 1 9 4 13 0 9 1 0 9 7 3 13 15 13 1 3 0 9 2
8 11 13 9 4 4 13 15 2
3 9 2 11
31 9 13 3 11 1 14 2 13 7 13 2 0 9 3 1 9 7 14 2 8 1 9 1 10 0 9 1 0 9 2 2
24 9 1 9 11 11 13 0 2 7 16 9 13 1 14 13 3 2 13 9 9 11 11 9 2
11 9 0 9 13 3 3 1 10 0 9 2
9 3 13 10 0 9 1 0 9 2
46 9 7 9 2 13 2 1 10 9 2 15 4 13 1 9 2 9 1 10 0 9 2 7 13 2 16 9 3 13 9 9 1 2 16 13 4 13 9 1 14 13 10 9 1 9 2
10 7 3 13 15 1 9 2 15 13 2
7 15 13 3 3 1 11 2
37 1 10 0 9 13 9 3 1 9 1 14 4 13 9 1 10 0 9 1 10 0 9 2 16 15 13 1 11 1 9 1 9 1 9 11 9 2
1 8
19 15 13 10 0 7 0 9 7 13 3 3 1 9 3 2 2 13 9 2
45 2 7 16 15 13 3 1 15 2 16 10 9 4 13 1 10 0 9 1 9 2 13 15 14 13 10 9 2 9 7 10 9 3 4 13 9 1 1 0 9 2 2 13 15 2
53 15 4 0 14 13 2 0 9 2 1 15 2 15 15 13 1 2 0 9 2 2 2 15 11 3 13 2 2 7 9 13 3 2 1 9 0 9 13 1 10 9 2 10 0 9 9 4 4 3 3 0 1 2
25 15 13 3 1 9 2 16 10 0 9 1 9 13 2 7 9 1 9 9 13 15 1 10 0 2
32 9 4 13 10 9 1 14 13 15 1 9 2 7 10 9 13 15 3 3 1 9 2 7 3 13 15 3 1 9 2 3 2
7 1 10 9 13 15 3 2
13 10 9 13 15 3 7 3 1 10 9 9 11 2
43 0 10 0 0 9 13 1 9 11 11 1 10 0 9 1 11 2 10 0 0 9 2 7 15 13 15 3 1 0 2 16 9 9 7 9 11 11 3 4 11 0 9 2
12 2 15 13 3 7 15 4 15 3 13 3 2
13 6 2 6 2 15 13 9 3 3 1 9 1 2
23 15 4 0 7 0 2 10 9 1 10 0 9 1 15 2 0 1 0 9 7 0 9 2
10 15 4 10 9 2 15 13 1 9 2
18 2 15 4 3 0 2 16 15 3 13 10 9 2 1 9 0 9 2
46 15 4 15 2 15 3 4 13 10 3 3 0 9 3 2 7 3 13 10 9 1 10 0 9 1 9 1 14 13 3 2 15 3 4 9 2 15 3 4 9 7 15 3 4 3 2
17 9 13 10 0 9 7 10 9 2 15 4 3 1 14 13 9 2
19 9 4 0 1 10 9 2 9 13 1 13 9 7 13 1 9 1 9 2
8 7 15 4 3 10 0 9 2
21 9 7 10 0 9 13 1 11 1 9 8 2 7 15 4 0 9 2 15 13 2
5 7 15 4 13 2
6 15 13 15 4 0 2
31 3 3 13 15 1 0 9 1 9 2 3 1 0 0 9 4 4 13 3 3 3 1 3 3 1 9 1 10 0 9 2
20 15 13 3 1 10 0 9 2 16 3 13 3 9 7 9 1 9 9 1 2
8 9 4 13 1 12 9 9 2
36 2 15 4 13 10 0 1 9 1 9 11 2 7 15 4 3 13 15 3 1 9 2 2 13 11 11 1 9 11 2 15 4 13 1 9 2
14 15 13 15 3 1 9 1 10 9 2 15 13 1 2
7 9 3 13 15 1 15 2
8 11 13 3 10 9 1 9 2
3 15 1 9
10 2 11 4 3 10 0 9 1 15 2
4 8 4 3 3
13 15 4 3 0 2 7 3 10 9 9 4 13 2
31 16 15 3 13 1 11 1 12 2 4 15 1 10 0 9 3 13 1 9 2 15 13 7 13 1 15 7 13 15 9 2
23 7 1 11 11 9 2 2 16 11 13 10 9 2 4 15 13 15 1 14 4 3 2 2
5 3 13 15 3 2
11 3 9 1 0 9 2 7 1 9 9 2
16 2 15 13 3 2 15 3 4 3 2 2 13 10 0 9 2
5 11 4 12 9 2
17 9 13 3 2 16 11 9 1 9 11 4 10 0 9 1 9 2
42 0 9 4 3 13 3 2 16 9 13 10 3 0 9 2 7 0 13 1 2 16 9 4 13 1 9 2 15 9 12 9 13 10 0 9 1 2 0 9 2 9 2
14 15 13 2 16 15 13 10 9 2 15 3 4 13 2
9 7 15 13 1 15 1 10 9 2
13 3 4 15 4 13 2 16 15 13 9 1 9 2
1 9
19 9 4 12 9 3 1 10 9 13 9 1 10 0 9 3 1 9 9 2
15 9 13 1 0 0 9 2 1 9 13 3 1 1 9 2
52 1 10 9 3 9 3 7 3 13 1 9 7 1 9 2 7 3 15 9 13 1 10 0 9 2 13 15 13 7 13 1 9 14 13 13 1 10 9 1 9 2 15 4 13 8 9 1 10 0 9 9 2
13 13 3 10 2 9 2 2 15 13 3 1 12 2
8 2 15 4 9 2 13 11 2
4 15 4 9 2
31 16 9 13 15 2 13 15 15 3 1 10 9 2 11 11 2 11 2 14 13 13 9 1 15 1 10 9 1 11 9 2
22 15 13 1 10 9 9 1 9 2 7 3 3 10 9 13 15 14 13 9 1 9 2
16 2 15 4 3 4 15 2 15 4 13 15 0 10 10 9 2
32 3 4 15 3 3 9 9 2 15 13 1 15 2 16 15 1 9 1 10 9 3 13 14 13 3 1 14 13 1 9 2 2
11 9 15 1 3 3 4 13 3 1 9 2
28 2 0 15 14 13 10 9 2 15 13 10 0 1 9 2 2 13 10 0 9 7 13 1 10 9 1 9 2
10 3 13 15 9 9 1 14 13 3 2
13 0 2 13 9 1 0 9 13 1 9 1 9 2
23 3 1 9 2 3 1 9 11 3 0 9 2 13 12 0 9 9 2 16 15 13 9 2
4 15 4 0 2
17 10 9 13 1 0 9 4 13 9 2 16 15 4 13 1 9 2
12 2 0 2 3 4 15 13 1 15 1 9 2
12 2 10 9 13 10 0 9 2 2 13 11 2
10 15 4 3 3 13 15 1 12 9 2
9 3 10 9 2 7 10 0 9 2
15 13 9 1 10 0 1 2 9 2 9 12 2 12 11 11
15 3 13 15 3 3 3 1 14 13 15 3 1 10 11 2
35 7 15 4 13 2 16 9 7 9 13 1 10 9 0 9 13 2 16 15 1 9 13 9 1 10 0 9 1 10 0 9 1 0 9 2
18 11 0 9 13 1 12 9 13 1 3 12 9 2 3 12 9 9 2
15 2 15 4 3 13 2 16 15 4 13 1 9 1 9 2
41 1 9 12 13 9 11 11 3 1 9 1 10 12 0 0 9 1 11 15 8 7 8 2 15 4 13 11 1 10 0 9 1 10 3 13 9 1 9 1 9 2
5 3 0 4 15 2
73 9 7 9 11 11 2 15 13 3 1 15 1 9 2 9 1 11 2 2 13 2 16 9 3 4 13 1 9 2 2 0 11 2 0 3 2 15 13 2 15 4 4 13 10 0 9 2 2 1 9 1 10 3 9 9 2 15 3 1 9 4 13 3 2 16 9 1 10 9 3 13 3 2
27 2 15 4 3 0 14 13 1 10 0 9 2 16 15 3 13 10 9 1 14 13 15 1 9 7 9 2
47 7 11 11 9 4 13 15 1 9 1 9 1 10 0 9 2 3 1 9 1 11 11 2 11 13 10 0 9 2 7 3 1 12 9 1 11 11 7 11 2 12 9 1 10 0 9 2
33 1 10 9 2 3 4 3 0 9 2 13 11 9 2 0 11 2 7 0 9 1 11 9 9 2 11 9 7 11 8 7 9 2
20 9 13 10 3 3 0 9 2 1 10 0 9 13 1 10 9 1 9 2 2
13 7 15 13 3 2 16 9 3 13 3 1 9 2
15 11 11 4 3 3 9 2 16 15 13 9 1 0 9 2
37 10 0 9 1 13 3 9 7 9 4 13 9 9 1 14 13 10 9 3 1 9 2 1 15 4 13 1 0 9 2 2 13 11 11 11 11 2
17 1 10 9 1 11 7 11 13 3 9 1 3 0 1 0 9 2
14 6 2 3 3 9 13 9 3 3 1 15 13 15 2
35 9 11 11 11 2 11 9 2 4 3 3 13 2 3 0 9 13 2 7 3 1 3 13 0 9 1 9 2 13 9 3 9 1 0 2
20 2 7 1 10 0 9 0 9 4 15 3 13 9 14 13 9 1 10 9 2
17 2 7 15 4 3 10 0 9 2 15 13 2 15 3 4 13 2
29 7 10 0 9 1 11 7 11 4 13 10 9 2 15 1 10 9 1 9 13 1 2 16 9 13 3 1 9 2
4 4 3 13 15
23 11 11 2 1 9 9 1 11 9 2 4 13 9 1 10 0 9 1 9 1 0 9 2
16 9 11 13 3 1 10 9 3 1 11 2 3 15 4 13 2
19 10 9 12 4 0 1 10 9 1 9 2 7 0 9 13 3 1 9 2
14 15 13 3 0 3 2 15 4 3 13 13 12 9 2
7 9 7 9 2 9 8 2
14 15 13 15 1 0 9 1 10 9 1 9 1 12 2
1 9
19 2 15 4 3 0 2 16 9 1 9 4 13 10 9 1 10 13 9 2
6 2 9 4 3 9 2
19 1 10 0 9 4 13 3 12 9 9 1 11 2 11 7 11 1 9 2
24 15 4 13 2 11 2 2 16 15 3 4 3 7 13 2 13 1 9 7 13 10 3 9 2
9 13 15 1 0 9 1 0 9 2
3 8 5 9
8 0 9 1 9 13 11 9 2
31 15 13 2 16 15 4 10 0 9 1 10 9 2 15 4 1 9 1 8 3 14 13 10 9 1 9 1 3 1 9 2
17 15 4 2 3 1 10 9 2 4 13 9 11 11 7 11 11 2
15 15 13 3 2 15 3 13 8 7 9 1 14 13 9 2
3 2 6 2
31 9 11 11 13 1 10 9 1 9 7 13 0 9 1 0 9 1 9 2 15 9 12 13 9 12 7 4 13 1 12 2
10 1 10 0 9 1 10 9 3 13 2
28 10 9 11 4 3 13 14 13 2 7 3 13 9 1 12 9 3 1 0 9 10 0 9 1 9 1 11 2
1 9
32 3 13 15 14 4 13 10 9 1 14 13 10 0 3 3 2 7 10 9 9 9 3 1 10 9 1 3 0 9 1 9 2
16 13 9 1 9 7 13 9 7 9 3 3 1 10 0 9 2
31 1 9 4 0 9 13 15 10 0 9 1 9 7 10 0 9 7 9 10 9 1 9 2 15 4 13 3 1 0 9 2
11 15 13 1 11 1 12 9 2 9 9 2
8 9 13 13 7 0 1 9 2
16 15 13 3 1 14 13 2 16 11 3 13 10 9 1 9 2
65 1 9 4 13 12 9 8 2 8 7 9 2 13 1 11 1 12 8 2 12 9 9 13 1 12 9 2 15 4 3 1 9 12 1 1 14 13 9 3 1 9 1 2 12 0 9 2 0 3 1 14 4 13 10 0 9 1 9 2 7 10 9 0 9 2
12 9 1 11 4 13 1 0 9 1 0 9 2
22 15 13 15 2 7 11 13 3 1 15 2 16 15 13 10 0 9 1 10 0 9 2
6 15 4 3 13 3 2
12 13 9 1 9 3 7 13 9 13 3 3 2
27 9 13 3 3 7 13 2 16 9 13 2 4 15 3 3 13 10 9 2 16 15 4 13 1 15 3 2
14 15 2 15 13 2 13 11 7 13 10 9 1 11 2
29 7 3 1 15 13 15 1 11 11 11 9 2 15 13 10 9 1 10 9 2 2 4 15 0 1 0 1 9 2
16 7 1 3 4 9 3 13 10 0 2 13 9 1 10 0 2
29 3 11 1 9 9 4 2 0 9 1 0 9 2 2 3 13 10 0 0 9 3 1 2 0 2 0 0 2 2
19 7 9 13 3 1 9 2 16 15 13 0 9 2 16 11 3 4 3 2
43 3 13 9 9 1 11 9 3 1 9 2 16 9 1 9 1 9 0 9 13 10 0 9 1 12 9 1 3 4 13 2 16 9 13 9 1 14 13 1 10 0 9 2
27 4 15 3 1 10 9 2 3 15 13 15 2 3 13 14 13 9 1 2 15 15 13 1 1 9 9 2
35 10 9 2 3 4 9 1 11 9 2 4 13 1 12 9 3 2 16 15 13 14 13 10 0 9 1 12 9 9 2 3 9 4 13 2
54 11 11 11 2 12 2 2 15 1 3 12 9 3 13 10 0 9 2 9 2 13 0 9 1 11 2 7 11 11 13 9 1 9 1 10 1 10 9 2 3 9 1 9 7 10 9 1 10 0 9 13 1 9 2
10 10 9 4 3 9 1 11 11 13 2
12 3 4 9 7 9 3 13 1 10 0 9 2
14 1 9 12 13 9 0 9 2 1 9 9 7 9 2
21 3 13 15 3 1 2 16 15 13 15 3 2 13 3 8 7 4 0 1 9 2
18 15 13 1 10 0 9 2 15 4 13 9 1 3 10 0 12 9 2
25 15 13 3 1 9 1 10 9 2 15 4 1 9 1 9 2 16 10 0 9 3 4 3 13 2
26 3 13 12 0 9 1 11 9 1 9 1 9 1 11 11 11 2 12 2 1 9 1 11 1 11 2
30 2 7 15 4 15 3 13 1 2 7 15 4 3 3 0 1 0 10 9 2 15 13 1 9 2 2 13 11 11 2
29 9 13 3 3 12 9 0 9 2 9 7 11 2 2 7 10 9 4 13 1 9 1 9 2 2 13 11 11 2
7 3 10 0 9 13 3 3
14 2 7 3 4 15 13 9 2 3 16 15 13 3 2
5 10 9 1 9 2
1 9
8 11 13 15 15 1 14 13 2
20 1 9 4 10 0 9 3 13 15 14 13 10 9 14 13 10 0 1 9 2
9 15 4 3 13 15 3 3 3 2
27 3 13 3 1 10 0 9 11 11 1 10 0 9 7 10 0 9 1 9 1 11 2 3 9 11 13 2
4 7 1 9 2
7 2 4 15 13 15 3 2
27 3 13 10 0 9 1 9 10 11 11 3 3 1 9 2 15 4 13 3 1 9 7 13 13 1 9 2
17 1 9 4 10 9 4 0 2 2 13 11 11 11 1 11 9 2
26 7 10 9 4 13 1 14 13 2 16 10 0 9 2 11 11 2 12 2 13 1 14 13 1 9 2
33 11 13 10 0 9 2 1 16 11 4 13 14 13 2 15 15 4 13 2 13 14 13 10 0 9 1 10 3 0 2 0 9 2
22 1 9 12 4 9 13 1 10 9 2 7 3 13 9 1 14 13 10 0 9 12 2
8 15 13 1 15 3 1 9 2
8 7 15 4 3 10 0 9 2
35 2 15 13 9 3 2 15 13 9 3 2 15 13 9 1 9 2 15 4 13 0 9 2 7 3 13 15 1 2 16 15 13 9 2 2
6 3 13 9 3 11 2
17 9 11 11 4 1 12 13 15 1 9 1 9 7 9 1 9 2
34 1 9 1 3 3 2 7 3 2 13 14 13 3 13 3 2 2 15 13 3 15 1 15 2 16 3 13 15 2 15 9 3 13 2
26 15 4 3 11 2 15 9 1 9 1 0 9 13 2 2 13 9 2 7 1 9 13 15 9 2 2
8 15 3 13 2 13 7 13 2
13 13 15 3 2 4 15 13 0 7 0 9 13 2
1 11
24 9 2 15 4 13 12 9 1 0 9 4 3 0 1 0 9 2 13 12 0 2 9 2 2
18 7 15 13 3 14 13 10 9 7 10 1 10 9 2 15 4 13 2
87 15 4 13 15 1 10 13 9 7 9 7 13 15 1 10 9 2 16 15 13 10 9 1 10 13 0 9 2 3 0 16 9 3 3 13 1 9 3 2 7 15 4 3 13 7 8 15 7 13 15 9 1 3 14 13 10 1 9 2 7 1 15 2 9 2 2 1 14 13 15 13 10 9 1 15 1 10 0 2 0 7 3 0 1 10 9 2
28 2 6 2 11 7 0 15 4 3 13 2 16 15 14 13 9 4 15 2 15 3 13 3 7 13 15 1 2
43 15 4 3 1 9 13 1 10 9 9 2 15 4 13 14 13 10 9 2 7 15 4 13 11 3 1 9 1 10 9 2 15 9 10 0 11 3 13 15 14 13 1 2
45 15 13 10 0 9 1 9 1 16 9 2 16 15 4 13 9 1 10 13 9 1 9 1 9 2 3 4 13 2 16 9 3 13 1 10 9 2 15 4 13 1 9 1 9 2
8 3 13 10 0 9 7 13 2
10 15 13 3 1 10 0 9 7 9 2
20 2 10 0 9 1 9 13 2 16 9 13 0 9 2 3 3 15 13 3 2
15 15 4 13 10 3 0 9 2 10 0 9 7 0 9 2
12 1 9 13 15 3 1 9 7 13 15 3 2
8 2 11 2 13 0 1 9 2
16 10 13 12 9 4 3 13 1 12 9 9 1 9 7 9 2
30 9 1 10 0 9 13 2 16 10 9 4 13 1 9 7 4 0 1 14 13 10 9 2 15 13 10 0 9 9 2
31 7 1 10 9 4 11 11 0 9 2 11 11 2 13 15 14 13 3 3 1 15 8 8 7 0 9 1 10 0 9 2
13 2 15 13 3 3 3 2 15 13 15 3 3 2
16 15 13 13 12 9 9 1 9 0 9 2 12 9 1 9 2
28 9 11 4 13 0 9 7 13 15 3 1 10 0 9 1 9 2 9 2 9 7 10 12 0 9 1 9 2
39 3 4 9 1 2 10 11 2 2 2 13 1 9 2 7 10 0 2 9 1 11 2 13 2 16 3 13 10 0 9 2 15 13 3 1 9 13 9 2
17 15 4 13 1 10 9 2 7 1 9 4 15 3 4 0 9 2
51 16 11 11 4 13 14 13 0 9 1 9 7 1 9 1 3 14 13 15 3 1 9 2 7 16 10 0 9 4 10 9 1 9 2 15 15 4 13 9 7 9 2 4 0 15 15 13 1 15 15 2
18 2 15 13 15 15 2 16 15 13 15 1 9 7 0 10 0 0 2
17 0 9 3 13 12 13 9 2 13 9 3 7 13 9 1 9 2
20 3 4 10 8 9 13 9 0 2 0 11 8 1 9 1 11 9 1 11 2
20 15 4 3 0 7 0 14 13 1 12 9 1 1 12 2 2 13 11 11 2
2 1 9
13 3 4 9 11 11 11 13 12 9 1 11 11 2
10 13 12 9 0 7 13 15 1 9 2
14 7 15 4 9 1 14 13 9 1 9 2 13 9 2
39 15 13 2 16 10 9 2 15 3 4 13 10 9 1 3 11 7 11 2 3 1 13 1 11 11 3 4 13 14 13 1 11 7 13 10 9 13 3 2
26 10 0 13 1 0 9 1 9 2 3 9 2 3 0 9 3 4 13 3 1 9 7 9 1 9 2
13 15 4 10 9 1 15 3 14 13 10 0 9 2
48 10 12 9 13 9 3 2 15 3 4 13 2 16 3 4 4 13 10 0 9 1 9 8 7 9 2 7 16 10 9 1 11 7 11 1 9 1 9 2 1 9 13 1 9 1 9 2 2
11 15 4 3 13 15 14 13 13 1 11 2
9 0 9 4 1 3 13 15 13 2
15 10 9 1 11 9 2 15 3 13 1 11 2 4 13 2
17 15 13 0 11 11 11 1 10 3 0 2 0 7 3 0 9 2
16 15 4 13 15 3 10 9 14 13 10 9 3 1 9 2 2
11 10 0 9 1 12 9 13 1 12 9 2
13 11 11 4 2 1 0 9 9 2 12 9 0 2
22 2 15 13 10 13 9 1 9 7 13 2 16 9 4 13 1 9 1 10 0 9 2
24 10 0 8 9 11 11 13 2 16 11 3 3 3 4 13 3 1 10 0 9 9 1 11 2
5 15 13 15 3 2
42 1 11 1 9 13 2 16 9 3 13 1 9 1 14 13 15 3 1 9 9 1 9 1 9 2 16 11 9 1 12 13 3 1 9 1 9 7 10 13 9 0 2
7 3 1 10 0 9 2 2
58 9 2 13 1 9 2 2 3 0 0 7 0 9 13 2 4 13 10 9 3 0 2 16 15 13 15 15 1 2 16 15 4 13 1 7 13 1 9 9 1 0 9 2 15 15 3 13 14 13 11 1 3 14 13 15 12 8 2
22 15 13 2 16 10 0 4 13 1 9 1 10 0 11 3 16 2 10 0 9 13 2
9 15 4 15 13 1 10 0 9 2
21 15 4 1 0 9 13 3 1 10 9 1 0 9 1 11 2 15 4 13 9 2
5 15 4 13 15 2
42 16 3 10 0 9 13 13 7 13 1 10 3 13 9 1 9 7 9 2 0 7 0 9 7 0 9 2 13 10 0 1 0 9 1 0 7 3 0 9 1 9 2
21 2 3 0 3 13 2 13 3 3 10 0 9 1 2 2 13 11 11 2 9 2
21 10 9 2 15 4 13 1 9 1 12 9 2 4 15 3 13 1 10 0 9 2
2 0 9
15 3 13 0 9 1 9 1 9 2 13 9 1 9 9 2
14 0 9 1 0 9 7 9 3 1 9 2 9 7 9
1 0
19 7 15 4 3 13 15 2 16 15 3 4 13 10 9 1 10 9 2 2
22 2 16 11 11 11 11 13 10 9 1 11 2 13 0 15 1 10 2 0 9 2 2
15 7 1 9 13 3 10 9 1 12 0 1 7 1 11 2
2 0 9
5 7 15 4 0 2
12 10 3 0 9 1 10 9 4 3 13 15 2
62 1 12 9 4 15 3 1 9 1 11 13 1 9 2 15 4 3 4 13 1 14 13 15 13 3 2 16 15 4 13 1 11 2 7 9 1 11 13 16 10 9 4 13 0 2 7 16 9 13 1 9 4 3 11 7 9 13 10 9 1 11 2
2 12 2
20 2 0 2 15 13 15 1 10 9 16 15 13 9 1 14 13 10 9 2 2
49 1 10 9 4 9 1 10 0 9 13 0 1 2 16 0 1 9 1 10 9 4 13 9 2 3 4 3 3 0 1 11 2 16 15 4 13 1 9 2 16 15 4 13 2 10 0 9 2 2
6 15 4 3 10 9 2
41 9 4 0 1 2 16 11 11 1 9 13 13 10 12 9 9 9 2 10 9 7 0 9 1 9 2 16 15 13 9 1 9 1 11 11 9 1 10 0 9 2
23 1 10 0 9 1 9 4 15 13 2 11 13 2 16 0 9 4 13 10 9 0 0 2
12 11 13 3 3 2 15 4 0 14 4 0 2
2 9 12
38 10 0 12 10 9 2 15 13 1 2 13 1 9 12 2 3 15 13 9 1 9 11 2 7 3 13 11 13 2 13 10 9 7 11 7 13 9 2
8 2 15 4 15 3 13 1 2
14 15 4 3 13 2 2 13 15 0 9 3 1 15 2
7 3 0 9 13 15 3 2
6 8 5 11 9 5 0
8 3 9 7 10 9 1 9 2
31 1 9 4 11 2 11 2 11 2 11 2 11 7 11 13 1 9 2 15 11 11 3 4 13 1 15 1 9 1 9 2
7 3 1 15 4 13 9 2
2 12 2
3 3 3 2
15 15 13 2 16 9 4 4 13 1 14 13 3 1 9 2
6 7 3 13 15 3 2
17 11 4 4 10 13 9 2 15 13 3 3 1 9 7 3 3 2
15 3 1 16 15 13 9 14 13 2 13 15 10 0 9 2
37 4 15 13 15 2 3 13 15 15 10 9 2 7 4 3 13 10 9 16 9 11 13 15 1 9 1 9 1 9 2 9 7 9 3 1 9 2
14 10 9 7 15 13 3 3 1 9 1 10 9 2 2
22 7 0 10 9 4 15 13 15 15 7 15 2 7 13 15 3 2 2 13 11 11 2
29 11 4 13 9 1 9 11 11 11 2 11 2 15 1 15 13 13 2 16 11 11 4 13 1 10 9 7 9 2
14 15 13 11 10 9 1 9 7 13 12 9 1 11 2
13 2 7 3 13 3 1 9 2 2 13 11 11 2
8 12 9 13 15 1 10 9 2
16 9 13 1 10 0 9 2 7 3 4 10 9 0 1 15 2
31 1 10 3 0 8 7 9 4 15 3 13 2 16 10 0 9 1 10 0 2 0 9 4 10 9 2 7 15 4 15 2
12 13 7 13 9 1 14 13 3 14 13 15 2
13 1 10 0 12 9 4 15 13 1 9 1 9 2
17 15 7 10 9 9 4 1 9 13 1 9 2 9 7 0 15 2
34 1 14 4 13 15 3 1 10 9 2 13 11 11 3 9 1 2 16 11 1 12 9 4 13 10 3 0 9 1 0 9 1 9 2
24 10 0 9 4 10 0 9 13 13 9 3 1 0 9 2 7 3 13 9 3 3 1 9 2
2 9 12
12 9 4 13 0 1 12 9 1 10 0 9 2
6 15 13 7 13 3 2
13 15 4 3 13 15 13 1 10 9 1 12 9 2
16 2 15 13 9 4 13 3 1 0 9 7 8 8 0 9 2
21 9 13 0 2 13 7 1 9 7 13 3 3 1 9 2 9 2 9 7 9 2
7 15 4 15 3 4 13 2
7 15 13 15 0 1 2 2
24 13 9 1 9 2 4 10 13 9 13 0 1 9 2 16 11 13 10 12 9 9 1 9 2
31 15 4 0 1 10 9 7 4 3 13 1 14 13 15 1 10 9 2 3 9 13 2 7 10 0 9 13 3 1 9 2
7 1 9 4 0 9 9 2
14 13 9 7 13 9 3 1 3 7 1 9 1 3 2
20 7 3 15 13 1 11 2 3 3 1 10 0 9 13 9 11 11 1 9 2
16 2 15 4 3 13 9 7 9 1 10 9 7 13 10 9 2
14 7 3 13 10 9 1 2 16 15 3 4 13 9 2
10 3 13 3 15 3 13 15 10 0 2
16 3 13 10 9 1 2 15 3 13 3 0 9 1 0 9 2
4 15 13 11 3
6 16 3 13 9 3 2
12 7 15 4 4 0 9 2 14 13 3 1 2
25 1 10 0 9 1 10 0 9 9 1 9 13 10 9 2 15 13 15 1 9 1 11 1 13 2
12 3 3 9 4 13 1 9 13 15 1 9 2
25 10 9 2 15 1 0 9 13 0 9 1 11 1 0 9 2 13 0 9 1 10 7 10 9 2
15 3 4 15 1 0 9 2 9 2 0 1 10 0 9 2
15 2 15 4 3 0 1 15 2 13 15 1 9 1 9 2
46 10 0 9 3 13 2 16 15 0 13 10 0 9 1 2 16 9 9 4 13 1 2 16 15 13 9 1 14 13 3 1 3 0 9 2 15 3 4 13 9 1 9 7 1 9 2
15 16 15 4 13 15 3 3 2 3 15 13 1 9 9 2
8 15 13 3 3 3 1 9 2
4 2 11 11 2
81 10 12 9 2 3 4 9 1 11 2 4 1 10 9 1 9 3 13 2 15 3 13 1 1 10 9 1 12 2 2 11 9 4 0 1 14 13 11 9 2 16 9 1 0 9 4 10 0 9 3 1 10 0 9 2 15 1 9 4 4 13 1 10 0 9 2 3 4 0 1 9 3 1 10 0 9 2 2 11 2 2
14 15 4 13 3 3 3 2 16 3 13 3 0 9 2
7 15 4 12 9 1 9 2
7 0 9 4 3 0 3 2
8 15 12 4 13 3 1 12 2
40 0 11 2 3 2 15 13 9 1 9 9 2 13 1 9 7 10 0 9 1 9 2 9 11 11 2 16 15 4 13 1 9 11 2 10 0 7 0 9 2
18 3 4 15 11 11 9 2 7 15 4 0 14 13 15 14 13 1 2
16 15 2 6 9 2 15 13 15 2 13 15 3 1 10 9 2
1 9
12 15 4 9 2 15 3 4 13 1 9 9 2
32 7 15 4 0 1 2 16 9 1 11 4 10 0 1 10 0 9 1 9 9 1 9 1 11 0 2 7 3 3 0 9 2
27 2 1 0 10 9 1 1 9 13 15 3 3 2 15 15 4 13 2 15 13 3 3 1 10 9 2 2
28 11 4 13 3 3 2 7 15 4 13 13 3 2 16 15 13 10 9 1 9 2 2 13 11 11 9 11 2
26 2 9 11 11 13 1 10 9 1 9 1 0 0 9 1 9 1 9 2 10 0 9 7 10 9 2
31 7 11 13 3 13 1 14 13 1 11 2 15 1 3 13 2 15 4 13 13 14 13 2 9 1 15 3 12 1 11 2
3 3 15 2
28 7 1 13 2 10 0 9 4 3 10 9 10 9 1 3 10 9 1 11 2 3 15 3 13 15 3 2 2
21 15 13 1 9 3 1 10 9 1 13 9 7 9 2 7 10 0 9 13 3 2
7 11 9 4 1 9 13 2
2 9 2
3 9 1 9
21 15 13 3 3 1 10 13 0 9 2 7 3 10 0 2 10 0 13 9 2 2
10 15 1 9 7 9 7 9 1 9 2
9 1 0 9 4 11 10 0 9 2
26 1 10 9 4 15 13 1 14 13 10 8 9 2 7 15 13 2 16 15 3 4 13 9 1 9 2
12 3 9 1 9 13 9 1 14 13 15 3 2
23 7 1 0 9 1 10 0 9 1 11 2 15 3 4 13 1 9 1 0 2 9 2 2
9 9 1 15 4 0 7 0 9 2
12 10 0 9 4 3 3 0 1 10 9 9 2
21 15 4 13 13 1 2 16 10 0 9 1 9 9 13 0 2 2 13 11 11 2
26 3 13 9 9 2 0 9 7 10 0 9 1 14 4 13 1 14 13 9 9 1 9 1 0 9 2
11 9 13 12 9 3 7 13 1 9 12 2
15 2 9 2 3 4 15 0 2 4 15 2 15 13 3 2
14 9 4 13 12 9 7 4 3 3 10 0 0 9 2
15 1 9 13 11 11 0 9 1 14 13 10 9 14 13 2
3 9 1 9
9 3 13 9 1 1 9 12 9 2
28 3 10 9 1 9 4 13 1 2 9 2 2 16 15 13 2 3 1 15 4 10 0 0 9 1 0 9 2
66 2 15 4 15 2 2 13 15 1 10 0 9 9 0 9 2 13 2 1 10 9 15 4 2 1 9 1 10 0 9 2 9 2 15 3 13 10 0 0 9 1 9 2 10 9 8 2 8 8 8 8 2 9 15 3 4 13 1 11 2 7 10 11 1 9 2
19 2 16 15 4 13 15 2 4 15 1 10 9 13 15 1 10 0 9 2
36 16 15 1 9 1 1 9 4 13 9 1 9 2 15 1 0 9 7 0 9 1 9 13 3 3 1 9 2 4 15 3 13 13 7 13 2
24 0 9 13 3 2 16 15 3 3 4 13 15 14 13 1 9 1 10 0 9 1 0 9 2
13 15 13 15 0 3 7 13 10 9 1 9 12 2
23 2 0 9 2 0 9 2 2 13 1 12 9 2 16 9 13 9 2 16 15 13 3 2
12 15 13 3 1 9 1 14 13 10 0 9 2
14 7 15 4 10 0 9 2 16 9 3 13 10 9 2
20 13 10 9 10 12 9 2 13 10 9 1 12 5 1 9 1 10 13 9 2
9 0 9 2 12 11 1 12 8 2
4 15 13 9 2
20 0 14 13 1 9 4 9 1 12 9 2 7 15 1 12 9 13 9 3 2
19 1 9 4 10 9 1 0 9 3 3 13 2 3 13 15 13 1 9 2
20 1 9 4 15 3 0 2 16 15 1 9 1 9 1 9 13 3 1 9 2
11 15 13 1 15 7 13 9 3 1 9 2
15 11 2 12 9 13 0 9 1 11 9 1 9 1 9 2
22 11 11 13 15 15 2 16 16 9 13 2 4 15 13 3 7 13 1 15 1 11 2
36 1 12 9 4 9 1 7 1 11 13 12 9 1 14 13 7 13 9 2 12 9 7 12 9 4 13 2 7 12 9 9 4 13 1 11 2
10 15 13 15 3 3 1 10 9 9 2
15 2 1 11 4 15 3 3 3 0 1 15 10 9 13 2
8 3 13 3 9 1 0 9 2
27 15 13 2 16 15 3 3 13 9 2 7 3 13 15 3 1 14 13 9 1 9 1 10 9 1 9 2
39 1 9 9 2 15 13 9 2 4 2 1 10 9 2 0 9 13 1 10 0 9 2 16 0 9 1 9 1 9 3 4 13 15 1 10 3 13 9 2
28 9 4 0 2 10 9 13 9 1 10 9 2 15 3 13 11 3 3 1 2 16 15 13 9 1 10 9 2
17 15 13 3 14 13 1 15 2 7 15 4 3 3 13 10 9 2
44 9 2 15 4 0 2 16 9 3 4 13 0 2 0 2 9 1 15 2 7 16 10 0 9 4 0 1 9 1 9 1 9 2 4 15 3 13 1 1 0 9 1 9 2
22 15 13 3 11 2 9 1 9 11 2 15 13 15 15 13 1 14 13 9 0 9 2
18 7 16 15 4 0 2 13 15 3 1 15 2 3 15 4 13 9 2
13 3 2 15 4 3 13 2 16 15 3 4 9 2
27 9 1 11 4 1 15 13 1 11 9 2 15 1 9 11 9 4 13 15 8 7 9 1 11 9 11 2
51 16 10 0 0 9 11 11 13 15 9 9 1 9 1 10 9 1 10 9 9 3 2 7 10 0 0 9 2 11 11 11 11 11 11 2 3 4 13 1 0 9 2 13 3 3 13 10 9 1 9 2
12 11 11 2 11 11 7 11 11 13 1 9 2
8 13 15 1 15 3 7 3 2
3 9 2 11
23 15 13 3 3 1 14 13 2 16 3 13 10 9 1 9 1 14 13 9 3 1 8 2
4 7 1 11 2
1 9
17 10 9 2 15 13 1 10 9 2 3 3 1 9 4 0 9 2
28 0 1 10 9 2 15 4 13 1 9 2 4 13 9 1 14 13 9 2 15 3 3 4 4 13 1 9 2
21 11 11 4 3 1 10 0 9 13 2 16 15 13 2 16 3 13 9 1 9 2
16 10 9 2 15 13 11 2 7 10 0 9 2 15 13 11 2
25 15 4 13 1 9 1 10 9 2 16 15 1 12 9 3 13 10 9 1 11 3 1 10 9 2
13 0 10 9 1 9 1 10 9 4 13 1 11 2
9 7 1 9 1 11 9 1 11 2
9 15 13 1 11 1 0 1 12 2
6 13 15 1 10 9 2
15 7 15 13 3 9 11 2 1 4 10 0 9 0 9 2
7 10 9 4 13 1 9 2
15 15 4 3 13 1 14 13 9 7 3 13 15 15 3 2
29 15 4 4 7 13 8 11 0 9 2 15 3 3 0 3 2 13 9 2 13 1 10 0 9 1 11 3 13 2
7 3 2 9 7 9 2 2
17 9 2 7 9 1 10 0 9 2 9 1 9 2 9 2 9 2
22 7 15 13 3 2 16 15 2 0 2 13 10 0 9 1 14 13 13 10 0 9 2
17 9 1 9 9 13 2 16 0 4 0 1 9 1 10 0 9 2
12 3 10 13 9 4 3 13 0 9 1 9 2
14 7 1 14 13 9 9 13 11 10 12 9 1 9 2
31 3 1 3 1 9 9 7 9 13 10 9 9 1 9 1 9 2 4 3 3 10 0 9 3 2 15 4 13 1 9 2
9 15 13 15 14 13 15 1 9 2
6 11 9 13 1 9 2
17 9 4 9 1 10 0 9 2 15 13 1 10 0 9 1 9 2
3 2 3 2
7 6 2 15 4 3 0 2
5 15 3 1 9 2
20 15 13 3 9 1 9 2 15 13 9 7 9 1 14 13 15 3 1 9 2
15 9 4 3 1 10 9 13 3 2 13 7 13 1 9 2
34 10 9 13 15 3 14 4 13 1 9 7 1 10 9 1 15 15 2 15 15 13 1 10 12 0 9 1 9 2 11 11 7 11 2
15 2 7 9 4 3 0 2 2 13 9 2 8 11 11 2
42 10 0 9 1 0 9 4 3 3 13 2 16 9 1 2 16 15 2 1 9 1 13 9 1 12 9 2 4 13 13 9 2 4 13 2 10 9 4 4 13 15 2
15 3 0 2 15 4 11 11 1 11 2 11 2 13 1 2
26 10 0 2 1 9 1 13 9 7 9 2 4 13 1 12 9 2 1 15 16 9 13 1 0 9 2
11 15 12 8 9 4 3 13 9 1 9 2
20 15 13 2 15 4 0 1 11 7 11 14 4 0 1 11 1 3 0 9 2
11 15 4 11 9 2 16 13 3 3 2 2
14 15 4 1 10 9 3 13 15 9 1 10 0 9 2
13 0 1 10 9 1 9 9 13 3 3 1 9 2
21 3 1 11 2 15 1 9 4 13 2 4 11 13 10 9 1 1 9 12 9 2
31 3 4 15 4 9 7 9 2 0 13 9 13 2 16 9 13 9 2 7 0 4 13 2 16 15 13 1 9 0 9 2
20 11 0 9 2 9 11 11 2 13 3 7 13 15 1 9 1 12 9 9 2
34 15 13 3 2 16 10 0 9 4 13 3 3 1 14 13 9 9 2 7 16 15 3 13 9 1 9 1 10 9 1 14 13 15 2
5 7 9 4 0 2
5 9 1 0 9 2
11 15 13 3 10 9 7 13 3 10 9 2
34 9 11 0 9 1 0 9 1 9 13 3 3 10 12 9 11 7 11 2 16 15 1 10 0 9 1 11 1 12 13 2 3 2 2
12 7 3 13 11 11 3 3 1 9 1 9 2
51 9 2 15 13 1 0 9 9 7 9 2 7 1 4 13 1 3 0 9 2 13 1 0 9 1 10 12 9 0 2 13 9 1 9 11 1 11 1 11 2 16 10 0 9 1 8 13 1 13 9 2
8 2 6 2 15 4 15 3 2
15 15 13 1 9 1 10 13 9 7 13 3 1 9 3 2
34 7 1 9 1 11 7 1 10 9 3 1 9 4 9 1 11 1 9 13 12 9 1 14 13 1 9 12 9 0 9 1 0 9 2
4 9 5 0 9
46 15 13 0 0 9 2 7 1 10 9 12 9 3 4 15 13 2 16 10 0 9 4 4 13 3 10 0 9 7 10 0 9 1 10 0 9 2 2 13 9 11 11 1 11 9 2
16 11 2 11 7 11 13 14 13 15 1 0 9 8 1 12 2
22 2 15 13 15 1 9 2 2 13 9 11 11 2 7 15 13 3 15 3 13 1 2
1 11
14 16 15 3 3 4 15 2 15 15 3 4 13 2 2
21 15 13 10 0 9 2 12 1 11 11 2 7 3 4 15 13 15 1 0 9 2
20 9 11 4 13 10 9 9 1 10 13 9 2 3 12 0 9 7 10 9 2
43 3 4 10 0 9 2 7 1 9 13 15 2 16 10 0 9 2 13 1 11 11 2 13 15 0 2 16 10 9 4 13 2 7 3 3 4 13 15 1 9 1 9 2
6 10 9 4 0 9 2
21 7 15 13 10 0 9 9 2 1 9 13 1 3 2 3 16 9 4 13 9 2
14 1 9 13 9 13 9 13 7 13 3 10 0 9 2
31 12 2 3 13 15 0 9 1 9 7 9 7 13 15 3 1 15 2 15 15 13 2 9 2 2 10 3 3 13 9 2
7 2 6 2 4 15 15 2
5 0 1 9 1 9
13 1 9 13 3 10 9 2 7 15 4 9 3 2
13 13 9 4 9 1 0 9 1 9 1 10 0 2
35 11 13 15 9 13 13 15 1 10 10 9 2 13 9 3 1 10 0 1 9 7 13 2 3 9 13 0 9 1 14 13 15 7 15 2
29 0 9 1 13 9 2 9 2 15 13 0 2 7 10 9 2 15 4 0 9 0 1 0 9 1 10 0 9 2
21 1 12 9 1 11 13 15 10 0 9 2 3 1 9 2 7 9 4 3 0 2
2 0 9
17 16 9 13 3 1 9 12 13 15 3 3 3 3 1 0 9 2
16 2 13 0 2 15 4 13 7 13 15 2 9 4 3 0 2
20 9 11 11 11 13 3 3 9 1 2 16 9 3 4 13 3 1 0 9 2
24 15 13 2 16 9 1 12 9 1 9 1 11 9 13 1 9 1 11 11 12 9 0 9 2
2 0 9
18 1 10 0 0 13 11 11 1 10 0 9 1 15 2 15 13 9 2
11 9 4 9 1 10 9 2 0 0 9 2
14 3 13 3 9 1 14 13 1 9 1 9 1 9 2
8 7 10 9 4 15 3 13 2
12 9 11 11 9 13 1 9 1 9 1 9 2
13 9 13 1 15 2 7 0 9 2 7 3 9 2
13 1 3 10 9 13 9 3 3 1 9 1 9 2
10 4 11 3 0 2 1 15 4 13 2
45 2 15 13 0 1 11 2 15 4 3 3 13 2 16 3 13 3 3 0 9 0 10 9 2 2 13 9 1 10 0 9 11 2 9 11 11 11 2 15 13 9 1 9 11 2
10 10 10 9 4 3 9 7 9 9 2
16 11 11 2 11 2 13 10 9 1 9 1 9 1 10 9 2
44 0 9 13 1 9 7 9 2 7 9 1 9 1 3 9 2 15 13 1 9 2 9 2 15 3 13 1 9 7 9 13 9 2 15 3 4 13 7 13 3 3 1 9 2
10 15 13 9 3 3 1 9 0 9 2
44 10 13 9 7 9 4 9 2 15 3 13 2 3 13 9 1 9 1 11 2 3 3 13 10 9 1 0 3 14 13 9 1 14 13 10 0 1 15 2 15 13 1 9 2
3 11 1 9
41 9 0 9 2 15 1 10 0 0 9 4 13 11 11 2 4 13 9 1 0 9 1 9 11 11 2 0 2 1 14 13 1 10 9 1 10 0 9 0 9 2
3 10 9 2
10 2 3 13 10 0 3 1 9 9 2
70 11 2 15 3 13 15 3 1 10 0 9 1 9 1 10 0 9 1 9 9 2 4 13 10 9 2 11 2 11 7 11 2 16 15 4 2 13 9 2 2 7 15 4 1 9 13 1 10 9 2 16 11 13 3 1 12 7 3 4 13 9 1 3 14 13 15 1 10 9 2
25 1 9 13 15 1 14 13 12 9 2 15 13 1 12 9 9 2 13 9 11 11 2 11 11 2
23 9 13 9 7 9 1 14 13 7 13 0 9 1 9 2 1 9 7 9 2 13 15 2
20 7 9 13 2 16 10 9 3 4 9 7 9 2 7 1 10 0 9 9 2
6 15 4 3 3 0 2
9 15 4 9 2 15 13 1 9 2
20 9 13 10 0 9 1 9 3 2 7 10 9 10 9 4 3 3 13 3 2
1 0
16 15 13 15 3 1 15 7 13 13 2 2 13 15 3 15 2
38 16 10 0 4 13 1 10 0 9 1 10 9 15 4 1 9 2 4 15 0 16 15 13 10 9 7 13 2 3 15 3 13 16 13 9 4 0 2
28 11 13 1 9 10 9 1 9 7 9 1 11 9 2 3 0 9 13 1 0 9 1 9 1 10 0 9 2
5 9 9 13 0 2
4 9 2 11 11
21 12 2 13 1 9 2 9 11 11 1 2 9 0 9 2 1 11 11 2 11 2
10 11 11 15 13 3 10 9 13 9 2
17 11 11 4 12 9 2 13 1 11 7 9 1 10 0 0 9 2
8 2 15 15 2 13 11 13 2
20 10 12 9 4 11 11 11 2 10 0 11 11 7 10 0 11 11 11 11 2
10 1 0 9 4 15 3 0 1 9 2
2 9 5
32 11 4 9 1 9 2 9 7 9 2 3 4 0 1 3 9 7 9 1 9 2 7 13 1 3 3 10 9 2 15 13 2
13 15 4 13 1 11 1 0 9 1 11 0 9 2
33 15 13 4 10 0 11 11 2 11 2 7 11 11 11 2 12 2 11 2 7 11 11 9 2 11 11 11 11 2 12 2 11 2
8 1 11 11 11 2 11 2 2
24 9 4 3 0 7 0 2 7 13 1 10 12 5 9 1 9 10 9 1 3 3 12 9 2
16 9 1 10 0 9 2 15 3 13 1 9 2 13 15 9 2
8 15 13 1 14 13 3 3 2
37 15 4 3 2 16 0 10 9 2 13 3 1 9 2 7 15 4 3 9 2 11 11 4 13 3 1 2 16 10 9 4 13 1 10 0 9 2
4 15 4 0 2
22 2 1 3 0 9 4 9 13 3 1 9 7 13 9 2 7 3 4 9 4 0 2
8 2 6 2 15 13 15 3 2
31 11 9 13 3 9 1 0 12 9 2 16 15 4 13 10 12 9 1 10 12 9 0 9 9 1 10 9 1 12 8 2
12 15 13 15 16 15 13 14 13 1 10 9 2
5 13 3 1 9 2
5 2 9 4 0 2
13 3 1 9 13 10 0 9 1 10 9 1 9 2
11 15 13 1 9 7 13 15 1 0 9 2
4 15 1 9 2
9 1 9 13 9 1 9 1 9 2
57 1 10 12 9 4 11 11 13 14 13 15 1 10 0 9 2 13 1 9 8 7 0 9 2 16 11 11 3 4 13 14 13 15 0 1 14 13 0 9 1 11 11 9 2 3 7 0 1 9 1 10 9 7 9 1 9 2
18 2 15 4 0 2 16 9 13 9 1 11 2 7 13 1 11 2 2
9 16 15 13 3 13 15 1 9 2
13 9 13 3 9 1 9 2 15 13 9 1 15 2
22 6 2 3 13 15 15 3 2 7 3 13 3 15 2 3 4 4 3 14 13 3 2
36 11 9 4 3 13 10 0 9 1 10 0 9 2 7 16 15 3 1 3 4 13 15 13 1 10 9 2 4 15 3 13 2 3 15 13 2
28 15 13 3 3 1 14 13 1 2 7 13 10 9 10 0 9 2 16 3 3 13 9 2 1 1 9 2 2
4 9 4 0 2
18 5 9 4 13 10 0 9 2 15 13 0 2 9 2 3 1 9 2
49 15 4 1 9 13 10 9 1 10 0 9 1 1 10 0 9 11 11 1 11 1 11 11 2 11 11 11 7 11 11 7 1 10 10 9 11 11 1 11 1 11 11 2 11 11 7 11 11 2
14 10 0 9 13 3 2 16 0 9 13 10 0 9 2
22 9 1 11 13 2 16 9 3 13 0 9 2 7 3 13 10 0 9 1 0 9 2
17 10 12 0 9 13 1 0 9 2 3 9 2 9 7 1 9 2
29 10 10 9 1 9 2 13 15 2 4 10 9 2 0 9 13 1 11 1 14 13 13 10 9 1 10 13 9 2
12 1 1 0 10 9 4 9 4 10 0 9 2
26 13 1 10 9 1 8 9 4 10 0 9 11 11 13 12 9 3 1 9 1 14 13 10 3 0 9
15 2 6 2 15 4 13 15 1 2 16 15 13 1 9 2
17 11 11 13 2 16 9 4 8 9 2 16 9 9 4 13 3 2
24 11 13 1 14 13 10 9 0 1 9 9 0 9 2 7 3 13 9 1 0 9 1 9 2
17 7 12 9 3 13 15 1 11 1 14 4 9 1 0 9 11 2
37 9 4 3 3 13 3 2 7 11 11 4 0 1 2 16 9 4 3 3 0 1 9 1 10 0 9 2 16 3 3 13 3 3 0 13 9 2
22 15 4 3 3 3 14 13 3 1 9 2 15 13 1 14 13 10 0 9 1 9 2
21 9 13 3 3 3 9 2 7 13 3 7 0 9 1 9 7 10 0 9 2 2
13 15 4 13 3 12 9 3 2 16 9 13 15 2
4 15 13 3 2
20 10 9 2 15 13 2 3 3 15 4 13 9 1 9 2 0 9 7 9 2
10 3 0 1 10 9 4 13 4 0 2
25 1 9 1 9 4 11 11 2 3 3 4 9 1 11 2 1 10 0 9 13 10 9 0 9 2
20 10 0 0 1 9 13 2 16 15 4 13 0 9 1 10 9 1 15 15 2
24 3 13 15 15 15 1 10 0 0 9 2 15 3 13 10 9 1 10 0 9 7 10 9 2
5 15 13 1 11 2
11 2 15 13 9 1 3 0 2 0 9 2
8 9 4 13 1 10 9 9 2
7 13 3 9 2 9 2 2
18 15 13 0 9 7 4 13 1 0 10 9 2 15 9 4 4 13 2
19 3 4 15 3 4 13 15 1 14 4 13 10 9 1 14 13 15 13 2
8 0 9 4 15 3 3 0 2
20 15 4 0 7 4 4 0 14 13 9 7 13 15 2 3 16 15 13 3 2
1 13
6 7 15 4 13 3 2
26 9 1 9 4 13 9 2 15 15 3 13 3 13 1 9 2 7 1 9 1 2 3 15 4 13 2
6 8 5 8 9 5 8
8 15 13 9 1 3 12 9 2
12 15 4 13 3 2 7 15 4 13 0 9 2
8 11 11 13 7 13 9 3 2
22 9 1 11 13 15 1 10 12 0 2 1 16 9 1 9 13 1 10 9 1 11 2
22 15 13 3 16 9 3 13 10 0 2 3 16 9 4 0 2 7 16 9 4 15 2
55 13 15 1 3 11 2 3 3 10 0 9 4 3 13 1 9 2 13 3 3 0 9 2 7 3 13 9 3 10 3 0 9 1 9 2 16 9 4 0 1 14 13 9 2 15 13 0 9 7 15 13 3 0 9 2
3 10 0 9
9 3 4 15 13 15 1 9 9 2
10 15 13 10 9 2 7 1 0 9 2
9 13 15 1 14 13 9 10 9 2
2 9 2
5 13 9 7 13 2
17 9 13 14 13 1 0 9 2 9 3 0 9 4 13 1 12 2
13 2 1 9 1 0 10 9 2 7 3 3 0 2
7 11 11 4 10 0 9 2
5 2 15 13 15 2
14 15 4 3 13 15 3 2 3 13 15 13 1 9 2
21 15 4 9 1 11 7 13 1 11 0 9 2 3 15 13 1 11 11 0 9 2
8 9 13 1 9 1 10 0 2
19 11 11 2 0 9 1 11 2 4 0 9 1 0 9 9 9 1 11 2
34 10 0 9 7 9 13 1 14 13 10 0 9 1 0 9 1 9 0 9 1 9 2 7 9 13 3 0 9 1 14 13 10 9 2
19 15 13 9 1 9 11 2 15 1 9 1 9 13 9 1 9 1 9 2
41 3 2 1 16 11 11 2 3 4 10 9 0 1 10 9 11 2 3 4 13 14 13 1 10 3 0 9 2 4 15 3 13 9 3 2 16 3 4 13 9 2
16 1 9 4 15 1 15 0 9 4 13 1 9 1 10 9 2
11 9 2 9 1 10 9 2 15 4 13 2
30 10 0 9 13 2 15 11 11 11 3 4 13 15 1 2 16 9 11 11 9 1 9 13 1 9 1 10 0 9 2
10 3 3 13 9 7 11 3 1 9 2
15 16 9 13 3 2 4 15 3 3 13 3 1 11 9 2
46 7 8 8 9 13 9 2 3 13 3 3 10 9 1 2 16 15 13 10 9 1 9 2 7 3 3 13 3 0 9 1 10 9 1 1 1 9 10 9 2 2 13 11 11 11 2
13 7 1 11 4 15 3 1 9 1 10 0 9 2
12 3 13 10 9 7 9 1 9 2 3 9 2
6 10 9 13 10 9 2
45 3 15 4 15 1 10 9 2 11 11 13 1 9 2 16 15 1 9 3 13 1 9 1 11 1 12 7 13 1 2 10 9 2 15 13 10 9 1 9 1 9 7 9 2 2
11 7 9 4 1 15 13 15 14 13 9 2
22 1 10 9 2 9 13 15 2 13 9 3 9 7 13 9 1 9 1 9 1 9 2
26 9 1 9 4 13 3 3 2 16 0 9 9 3 4 13 1 10 0 9 2 15 13 3 1 9 2
8 3 4 11 11 3 3 0 2
15 2 10 9 13 1 11 1 9 12 9 7 12 1 11 2
12 3 3 1 10 0 9 7 1 11 9 9 2
27 2 1 9 13 3 12 2 15 13 2 2 13 15 7 13 3 1 9 2 15 13 1 10 0 0 9 2
9 15 4 15 13 2 7 13 3 2
27 15 4 1 0 9 13 9 1 10 0 9 1 9 2 7 3 13 9 1 14 13 0 9 1 0 9 2
35 11 11 13 9 1 13 9 1 9 2 2 10 9 1 9 7 9 1 10 9 2 15 13 9 7 9 1 9 7 9 2 9 7 9 2
14 3 4 15 3 13 3 7 13 15 3 1 10 9 2
11 15 4 0 9 1 9 13 14 13 9 2
10 1 9 13 12 9 1 9 1 9 2
8 9 4 13 2 7 9 13 2
23 1 11 13 15 9 1 14 13 9 7 9 2 2 13 10 0 9 1 8 2 11 11 2
23 7 15 13 2 16 15 13 3 3 2 2 13 11 11 2 1 4 13 9 1 11 9 2
13 9 13 2 16 3 13 10 0 1 0 10 9 2
2 3 9
10 13 9 7 9 1 0 9 1 3 2
11 2 15 4 3 13 0 9 1 10 9 2
14 15 13 2 3 1 15 4 13 9 3 1 0 9 2
12 11 13 15 3 7 3 1 9 1 10 9 2
16 9 1 10 9 2 11 12 8 2 2 11 12 2 12 9 2
13 2 15 13 14 13 9 7 9 1 9 1 9 2
21 10 3 0 9 1 0 9 13 2 3 11 9 2 10 9 2 11 11 9 13 2
37 9 4 15 3 2 7 1 9 10 9 1 0 9 9 2 16 9 4 13 11 11 3 1 9 12 9 1 2 16 15 3 4 13 1 9 9 2
14 1 3 0 15 4 15 13 1 11 16 15 13 3 2
28 2 9 2 3 13 15 15 2 15 15 4 13 2 2 13 9 7 13 10 13 9 7 10 9 3 1 9 2
42 15 13 1 12 9 2 10 13 9 1 9 2 7 9 9 1 10 9 2 7 3 10 9 2 16 1 10 9 13 9 2 9 7 13 1 10 0 9 1 9 9 2
33 11 11 4 3 13 2 16 15 3 13 1 9 1 10 10 9 2 3 1 11 7 11 1 10 0 9 2 15 11 4 1 11 2
9 0 10 9 1 9 10 0 9 2
12 11 13 3 1 9 2 15 4 13 14 13 2
7 3 13 9 7 9 13 2
6 9 1 11 1 11 9
13 10 0 2 9 2 9 4 4 10 9 1 9 2
16 1 9 4 15 13 3 1 9 2 3 3 3 13 10 9 2
36 10 0 9 11 4 3 13 1 10 9 1 11 11 11 11 2 7 16 10 0 9 4 13 1 12 9 2 13 11 15 12 9 3 1 9 2
23 2 15 13 15 3 2 9 4 2 2 13 15 2 2 16 3 10 9 9 1 15 2 2
27 15 4 10 0 9 2 15 4 13 3 1 12 9 2 16 15 4 13 1 1 9 12 9 1 12 9 2
26 12 4 3 3 2 15 4 3 3 13 2 7 15 4 3 0 7 13 1 9 2 2 13 11 11 2
21 3 3 9 13 4 13 13 10 9 1 9 1 11 11 2 11 12 2 8 11 2
41 11 13 11 1 9 2 16 9 4 13 1 11 1 9 12 7 13 15 1 10 0 9 1 11 2 15 13 10 0 9 3 1 11 3 1 3 1 10 9 3 2
18 9 13 15 1 14 8 9 2 13 9 7 13 13 13 9 1 9 2
20 11 4 3 1 10 0 9 13 9 1 14 13 10 12 9 0 9 1 11 2
9 0 2 15 13 14 13 1 9 2
42 15 13 15 1 9 3 2 16 3 13 9 1 10 9 2 15 13 12 9 3 1 9 2 7 16 15 4 10 3 0 9 1 10 9 14 13 1 9 1 10 9 2
43 3 1 9 1 0 9 9 13 11 10 9 1 11 1 10 9 2 15 9 4 13 1 9 1 9 11 13 9 1 9 7 9 13 1 9 1 10 9 1 10 0 9 2
22 2 15 4 9 3 3 4 2 3 1 12 9 3 2 16 15 4 0 1 10 9 2
18 15 13 14 13 9 9 2 2 13 11 11 2 3 4 9 1 11 2
6 9 4 3 0 2 2
20 1 15 13 15 3 3 0 9 14 13 10 9 1 9 2 3 15 13 13 2
28 15 13 2 16 9 11 11 2 0 2 3 4 13 10 12 9 0 9 1 9 1 9 1 9 1 0 9 2
27 11 11 11 2 12 9 2 9 2 11 2 2 15 13 2 16 3 0 9 4 13 15 3 3 1 11 2
13 11 11 11 13 10 11 2 16 15 4 12 9 2
15 8 10 9 1 0 9 2 3 4 4 9 1 10 0 2
28 1 9 1 11 13 9 11 9 11 11 15 3 1 10 0 9 1 10 9 7 10 2 0 7 0 9 2 2
25 1 11 13 10 0 0 9 1 9 12 0 12 9 2 12 9 1 9 7 12 9 1 11 9 2
12 9 4 0 2 15 13 3 1 10 0 9 2
16 15 4 3 0 2 15 13 12 9 3 1 0 10 9 2 2
24 11 11 13 2 16 10 9 1 10 0 9 9 3 13 3 1 10 0 9 2 13 9 2 2
7 2 0 9 2 15 13 2
25 3 4 15 3 0 1 9 2 8 15 0 14 13 9 1 9 1 9 1 9 1 10 12 9 2
12 7 8 11 13 3 9 1 3 0 9 1 9
2 9 13
7 11 4 3 13 1 15 2
24 1 9 13 15 15 1 12 9 0 9 2 15 4 13 1 11 1 9 12 7 9 1 9 2
18 0 10 9 13 3 0 9 2 1 15 13 2 7 13 9 7 9 2
14 1 10 12 9 4 3 3 13 1 10 0 0 9 2
22 11 13 15 1 10 0 9 2 16 11 4 10 0 0 7 0 9 1 10 0 9 2
14 3 4 15 13 2 15 4 15 13 10 0 9 1 2
15 10 0 9 1 11 13 1 9 1 10 9 7 10 9 2
6 3 1 11 13 9 2
26 3 4 15 3 2 3 3 1 0 9 2 13 11 11 13 0 9 2 16 15 13 10 9 3 3 2
9 9 13 3 9 9 1 0 9 2
31 3 13 15 1 2 11 2 15 11 11 9 13 1 9 2 3 3 13 10 9 1 2 16 3 13 10 9 13 1 9 2
18 3 13 15 10 9 1 11 11 2 2 13 11 7 13 3 0 3 2
7 2 9 13 8 0 9 2
19 13 3 1 2 16 9 13 9 2 7 13 15 1 2 16 9 13 9 2
17 3 13 15 0 9 1 10 0 0 9 2 3 1 11 7 11 2
8 11 11 4 9 1 12 9 2
21 11 11 11 13 15 1 14 4 0 2 16 15 4 13 1 9 1 10 0 9 2
18 11 0 13 1 12 4 3 13 1 10 0 9 1 11 10 0 9 2
17 9 11 11 13 1 9 0 9 2 16 9 13 9 9 1 9 2
16 13 15 1 0 9 1 9 1 10 9 7 1 9 1 9 2
24 11 9 2 13 1 0 9 2 13 3 12 9 2 16 0 9 11 11 9 11 13 12 9 2
12 9 13 10 0 9 1 10 9 1 0 9 2
5 3 13 15 15 2
3 16 9 13
16 9 1 9 9 13 12 9 1 9 7 9 1 9 12 9 2
13 9 9 2 11 2 4 13 0 9 1 10 9 2
6 9 7 9 2 12 8
11 9 1 14 13 3 4 3 0 14 13 2
14 0 11 1 3 9 7 9 13 12 9 1 12 9 2
4 9 4 0 2
12 7 1 9 4 9 3 3 13 9 1 9 2
11 15 4 15 13 14 13 1 2 15 3 2
19 11 8 13 10 9 1 9 1 9 7 13 10 0 9 1 9 1 9 2
17 15 13 15 1 9 2 13 9 1 15 7 13 14 13 15 3 2
24 1 12 4 9 13 1 12 9 2 2 13 11 11 1 9 11 11 7 0 1 9 1 9 2
3 12 9 8
21 11 11 11 2 9 2 13 0 9 11 9 1 14 4 13 9 1 9 13 9 2
78 1 9 1 9 9 13 3 2 1 16 9 13 1 13 1 8 7 0 9 2 1 9 3 10 0 9 1 2 15 3 13 1 9 2 2 1 10 9 2 15 4 13 2 13 0 9 2 9 2 0 9 2 3 9 2 9 2 9 2 0 9 2 9 2 9 2 9 2 9 2 8 7 9 7 0 9 2 2
6 4 3 2 15 13 2
40 1 10 9 4 15 13 3 3 1 10 9 1 10 0 9 2 15 13 1 14 4 13 3 0 2 16 3 13 15 3 1 11 1 9 2 2 13 11 11 2
39 2 10 9 13 14 13 9 3 0 2 7 3 13 15 1 14 4 10 9 9 2 15 3 13 10 9 7 13 15 13 1 10 9 2 2 13 11 11 2
9 7 1 9 4 3 13 1 9 2
29 16 15 4 13 9 1 9 2 13 15 13 10 9 1 9 7 10 13 9 1 2 9 2 9 12 2 12 11 11
15 9 4 13 1 9 2 16 9 7 9 13 1 11 9 2
14 15 13 2 15 4 4 13 1 0 8 0 9 2 2
13 7 15 4 0 1 14 13 10 0 9 1 9 2
17 3 9 1 0 9 1 9 4 13 15 2 13 15 1 9 9 2
11 15 4 10 9 2 15 4 13 1 9 2
12 9 1 9 13 1 10 0 9 1 13 9 2
28 15 1 10 9 13 3 9 1 2 16 15 4 13 10 0 7 0 9 2 16 15 13 1 9 1 11 11 2
17 1 10 0 4 3 1 9 13 10 9 1 10 9 1 12 9 2
27 2 15 13 10 9 3 2 15 13 10 9 3 2 15 13 10 9 3 2 6 3 13 15 15 3 2 2
1 13
39 15 13 1 10 13 7 0 9 2 13 3 1 11 9 7 13 9 2 2 11 2 15 13 15 4 13 9 3 3 1 0 2 2 13 15 1 0 9 2
10 1 11 4 3 3 3 12 9 3 2
15 2 15 13 15 3 1 9 7 3 13 3 0 9 2 2
18 9 1 9 2 11 11 2 13 2 16 10 9 1 9 13 1 9 2
6 9 4 0 1 9 2
15 9 4 1 9 13 1 10 0 9 2 3 1 9 12 2
4 9 7 9 2
9 7 3 13 15 3 1 10 9 2
11 11 11 4 13 10 9 7 4 13 3 2
35 15 13 3 14 4 10 0 9 2 3 1 11 11 13 13 15 15 1 10 9 2 3 1 9 2 9 1 9 2 7 3 2 11 2 2
21 15 4 15 1 2 9 2 1 0 9 2 15 3 4 13 10 0 12 9 9 2
20 3 4 15 13 10 0 9 0 9 2 15 3 3 3 13 1 3 0 9 2
2 1 9
20 15 13 1 9 7 9 2 3 3 2 7 15 13 3 15 15 1 0 9 2
19 2 9 13 10 0 9 2 9 1 9 1 9 7 9 2 9 7 9 2
17 15 13 10 9 1 1 0 9 14 13 10 0 9 1 10 0 2
19 2 9 13 1 9 3 2 16 15 4 10 9 2 15 13 3 14 13 2
12 2 15 3 4 13 1 9 2 13 15 3 2
15 2 15 4 13 9 1 10 13 9 2 2 13 11 11 2
17 15 13 9 2 15 13 9 2 15 13 9 0 9 7 10 9 2
9 16 15 13 2 13 15 3 3 2
39 9 13 1 8 7 9 2 13 9 7 9 2 7 15 4 1 9 11 11 11 2 11 9 2 13 10 0 0 9 2 3 9 3 13 15 0 9 3 2
23 9 4 3 13 1 0 9 2 15 9 1 10 0 7 0 4 13 3 1 9 1 9 2
2 9 2
6 9 4 13 12 9 2
8 9 1 9 4 0 1 9 2
39 1 0 9 1 11 4 11 0 9 1 10 0 1 9 13 0 12 9 9 2 16 15 15 4 13 10 0 2 7 3 0 9 1 9 1 10 0 9 2
23 3 9 4 13 2 13 3 10 9 2 15 13 9 1 9 2 7 15 4 3 3 0 2
8 3 13 10 12 9 3 9 2
19 3 4 15 3 13 1 0 2 15 15 13 2 1 15 7 1 15 15 2
7 15 4 10 9 1 9 2
7 15 13 15 3 10 9 2
14 7 15 13 15 1 9 7 15 9 13 10 9 3 2
7 16 3 2 4 15 0 2
6 15 13 3 1 9 2
52 1 3 0 10 9 1 10 2 11 11 2 11 11 2 11 11 2 11 11 7 11 11 2 4 15 10 9 2 16 3 13 3 0 1 10 9 2 3 15 0 4 3 2 15 3 13 9 1 10 13 9 2
18 1 9 2 3 11 7 11 4 4 9 2 4 15 13 1 12 9 2
24 0 9 1 11 1 11 13 1 9 9 1 10 9 1 11 2 3 9 1 9 1 11 13 2
13 9 4 4 15 1 9 3 9 10 0 9 12 2
29 3 3 1 10 9 1 11 2 9 7 11 4 3 0 2 13 15 9 10 9 3 3 1 15 9 7 15 9 2
11 10 0 9 3 4 9 1 9 1 9 2
21 9 4 13 1 0 9 2 3 0 7 9 2 3 10 0 7 10 9 4 9 2
11 15 4 9 0 9 7 4 1 9 9 2
10 2 15 13 3 1 9 3 1 15 2
19 15 13 15 9 1 2 1 16 9 4 4 0 3 1 0 9 1 9 2
10 1 9 4 15 13 3 3 15 13 2
7 1 9 4 11 11 0 2
5 15 13 9 3 2
23 1 11 4 9 3 13 3 1 9 1 0 9 2 16 15 13 3 7 13 10 9 9 2
12 15 4 3 13 1 11 2 16 15 13 2 2
9 15 13 3 1 11 7 15 13 2
20 9 7 9 13 3 2 7 9 13 1 9 1 14 13 9 1 9 1 9 2
59 9 4 1 10 0 9 13 10 9 1 9 1 9 11 11 2 2 11 2 7 2 11 11 2 2 2 11 11 2 2 11 11 2 2 7 11 11 2 2 13 1 9 2 2 2 11 2 2 2 15 8 13 0 9 1 9 1 9 2
2 0 9
6 13 1 9 1 9 9
3 9 1 11
2 13 15
46 2 15 13 3 10 11 11 9 1 12 9 7 3 10 11 12 9 2 11 12 9 1 0 9 7 10 9 9 9 2 11 12 1 9 7 9 3 9 2 7 11 12 11 1 9 2
12 9 13 3 3 1 12 1 15 1 11 9 2
26 11 13 1 9 2 13 1 15 15 2 2 6 2 13 15 2 2 15 13 15 3 3 2 3 3 2
19 2 3 3 4 15 0 2 7 3 13 3 10 9 2 13 10 0 9 2
5 9 13 1 9 2
20 15 1 9 13 0 1 15 3 13 9 1 2 15 4 15 3 4 3 0 2
7 9 1 9 13 1 12 2
35 3 12 9 2 1 4 3 1 10 13 9 2 16 15 13 3 1 9 11 11 11 2 16 15 4 0 9 2 15 13 3 7 13 9 2
20 15 4 3 10 9 2 16 15 13 2 0 9 2 1 9 2 16 9 13 2
22 1 9 13 10 9 2 16 11 13 3 1 1 9 14 13 9 2 16 15 13 9 2
36 1 9 1 10 0 9 9 7 0 9 9 1 11 13 3 3 3 3 1 10 0 9 2 7 9 9 1 9 1 9 9 4 13 3 3 2
15 11 7 9 4 3 13 1 14 13 0 9 9 7 9 2
23 2 6 2 15 13 2 3 0 9 1 15 2 0 9 7 9 14 13 2 15 13 15 2
13 7 15 4 13 15 2 16 15 3 13 10 9 2
25 15 13 15 2 3 15 3 4 13 1 14 13 1 11 2 16 15 3 4 10 0 9 1 9 2
12 10 9 13 13 1 0 11 1 12 9 3 2
11 10 0 13 3 0 2 0 7 0 9 2
10 2 9 13 3 2 2 13 11 11 2
27 7 10 0 9 4 3 4 13 12 9 3 0 9 1 10 0 9 7 3 13 10 0 9 1 12 9 2
4 9 4 0 2
21 1 9 4 10 12 9 1 10 0 9 3 4 3 0 2 13 15 1 0 9 2
3 3 5 12
11 2 15 4 3 3 10 0 9 14 13 2
3 9 5 8
25 7 3 0 1 15 3 13 1 2 7 15 9 13 4 3 3 15 15 13 2 3 15 15 13 2
16 1 11 11 13 10 13 9 3 3 1 9 1 14 13 9 2
9 7 6 2 15 4 3 3 0 2
6 11 13 3 1 9 2
31 15 4 3 13 3 2 7 13 3 2 7 10 9 11 2 15 3 4 13 15 2 16 11 4 13 15 2 13 15 3 2
9 11 4 3 13 10 9 1 11 2
34 15 13 15 2 16 15 13 1 11 11 11 1 11 11 7 11 11 2 3 0 9 7 9 13 3 9 1 7 13 15 1 10 9 2
11 10 9 1 15 13 2 16 15 4 13 2
37 1 0 9 13 15 3 10 9 9 1 3 11 1 1 11 2 7 15 4 3 10 9 2 16 15 4 13 10 9 2 16 10 9 4 0 2 2
17 10 9 13 15 3 13 2 16 15 4 3 16 15 13 1 9 2
28 2 15 4 3 13 9 1 10 0 9 2 7 15 4 13 0 9 1 2 16 10 9 4 0 1 10 9 2
40 15 4 3 0 14 13 3 1 10 9 7 13 1 9 1 3 10 9 2 7 3 4 15 3 3 0 14 13 3 1 14 13 2 16 15 3 4 0 3 2
23 15 13 1 2 16 9 4 13 2 16 15 4 13 9 2 2 13 9 11 11 2 9 2
18 15 13 3 14 13 1 10 0 9 2 1 10 0 7 8 8 9 2
27 15 13 0 3 1 9 1 10 12 9 2 15 4 13 3 1 0 9 1 10 0 2 0 2 0 9 2
20 7 15 4 3 4 3 0 2 16 0 9 1 11 4 3 1 0 10 9 2
16 10 0 9 1 10 9 2 15 13 1 11 2 13 1 11 2
29 9 9 1 11 11 4 13 10 3 3 0 9 1 10 0 2 0 9 2 15 9 3 13 3 1 10 0 9 2
9 11 7 11 4 0 1 10 9 2
14 12 9 1 0 9 13 1 9 7 12 9 1 9 2
24 1 11 13 10 0 9 7 1 11 10 9 1 9 2 9 1 9 9 13 15 1 14 13 2
11 9 0 13 0 9 8 7 9 1 11 2
11 3 4 15 13 2 3 15 4 13 3 2
5 15 4 1 12 2
11 1 9 13 12 9 1 12 9 1 12 2
18 7 15 4 3 10 3 0 9 2 16 9 4 0 2 2 13 15 2
2 12 2
7 15 13 10 9 1 11 2
13 15 4 3 0 2 7 13 3 1 14 13 9 2
39 15 4 3 13 1 9 2 7 3 13 11 11 7 11 11 1 10 9 1 14 4 3 3 2 3 10 3 0 9 13 2 1 14 13 9 13 1 9 2
12 15 13 3 1 2 16 15 13 1 0 9 2
25 10 9 13 10 0 9 1 9 1 2 15 15 13 1 9 2 15 13 9 7 9 3 1 9 2
28 3 13 10 0 1 9 2 0 15 2 3 4 4 0 1 14 4 13 7 13 3 1 10 0 9 1 11 2
6 2 15 4 3 13 2
5 15 13 3 1 2
27 10 9 4 11 11 13 1 11 1 12 1 10 12 9 2 15 4 13 2 16 15 13 15 1 10 9 2
29 11 11 4 15 1 11 0 9 2 7 15 4 13 15 3 1 9 1 11 3 1 11 2 13 1 9 7 9 2
30 0 9 4 3 3 0 3 4 9 4 0 7 3 13 2 3 15 13 9 1 0 9 7 15 4 3 3 3 0 2
4 11 11 13 9
35 9 4 13 15 14 13 15 1 1 10 9 1 11 2 3 3 3 4 0 1 3 9 7 10 9 1 9 2 2 13 11 11 11 11 2
5 2 16 2 6 2
19 2 11 2 13 2 13 15 1 15 2 7 15 13 13 0 1 10 9 2
16 1 10 10 9 4 15 0 1 14 13 0 1 14 13 9 2
8 15 4 3 13 10 0 9 2
27 13 15 3 0 10 9 2 3 15 1 9 13 3 1 9 7 3 3 13 14 13 3 1 10 0 9 2
15 1 0 9 4 15 10 9 16 9 4 13 1 0 9 2
14 15 4 13 9 2 3 3 4 13 9 1 0 9 2
23 9 11 10 0 9 2 13 2 16 4 15 10 9 13 1 11 9 2 4 15 13 3 2
23 0 2 9 2 1 11 9 1 15 15 1 9 9 2 9 11 2 4 0 2 9 2 2
20 0 8 1 10 0 9 2 3 0 11 11 2 11 11 11 2 1 0 9 2
15 2 15 13 3 1 10 3 0 2 9 2 1 0 9 2
12 10 9 4 4 3 1 14 13 7 13 9 2
25 1 15 0 9 7 0 9 4 3 13 9 2 16 9 4 13 3 2 16 15 13 10 0 9 2
33 15 4 3 13 1 15 2 16 9 13 10 9 2 16 9 13 7 9 1 10 0 9 4 13 3 1 10 0 9 1 10 9 2
25 15 4 0 14 13 2 3 10 0 7 9 1 0 3 4 13 10 9 1 14 13 10 0 9 2
7 2 6 2 15 4 15 2
10 2 9 9 2 4 15 3 13 2 2
8 11 7 11 11 13 1 15 2
23 15 13 13 2 16 9 9 4 4 4 3 1 9 2 7 15 13 9 3 1 0 9 2
21 1 10 0 9 4 15 13 10 9 2 15 13 2 3 9 13 9 7 13 15 2
5 15 13 15 15 2
21 10 9 2 15 13 3 1 9 7 3 13 3 14 13 1 1 9 2 13 9 2
26 1 12 9 13 3 10 0 9 11 11 2 15 3 4 13 9 2 7 1 10 0 9 9 11 11 2
21 10 0 9 13 1 3 0 11 11 11 2 3 4 9 2 9 7 9 1 9 2
4 2 11 2 2
10 16 11 4 0 2 4 10 0 9 2
19 15 13 3 1 11 3 3 1 9 2 7 15 13 3 1 15 1 9 2
28 11 11 13 9 1 10 0 9 2 15 15 4 13 15 1 1 10 9 2 15 9 11 11 13 1 10 9 2
12 7 15 13 3 14 13 10 0 7 0 9 2
5 9 2 11 11 2
25 7 0 4 15 14 13 10 0 9 2 3 9 4 13 1 10 0 9 2 15 1 9 13 3 2
29 3 3 3 13 9 2 4 3 1 9 13 9 7 13 2 15 13 10 9 2 7 9 13 3 3 1 0 9 2
20 13 13 2 16 9 4 13 10 9 2 3 16 15 13 10 0 9 1 9 2
28 15 13 3 2 16 0 9 4 0 1 14 13 0 1 9 1 9 1 8 9 2 2 13 11 11 11 11 2
16 13 15 3 3 2 3 13 15 1 9 15 3 13 1 11 2
2 0 9
13 7 15 4 3 4 0 1 15 2 3 10 9 2
2 9 2
8 3 4 15 1 15 4 9 2
54 1 10 9 13 0 3 1 0 9 15 1 11 7 13 15 1 14 13 1 10 0 9 2 1 11 4 0 7 0 1 2 7 3 4 15 9 13 1 9 2 2 13 10 0 9 1 3 9 11 7 11 1 11 2
6 7 15 13 15 0 2
32 9 2 15 13 12 9 2 8 2 8 7 9 2 13 3 1 9 1 11 2 7 3 4 12 9 1 9 13 9 1 9 2
21 2 9 4 1 9 3 0 9 2 15 4 13 10 0 9 1 9 1 10 9 2
5 3 13 9 3 2
4 1 10 9 2
11 15 4 9 2 15 3 2 3 10 9 2
22 15 4 13 15 2 15 15 4 13 2 7 15 15 4 13 1 15 2 2 13 15 2
14 2 6 2 15 4 11 3 2 13 15 15 15 13 2
7 11 11 4 9 0 9 2
14 0 2 16 15 13 1 9 7 9 13 9 1 9 2
11 3 13 10 0 10 13 9 1 10 9 2
26 1 10 9 1 11 13 9 1 9 0 9 1 10 9 1 12 0 9 1 0 9 7 9 1 9 2
43 9 4 3 13 10 0 9 1 9 1 9 2 7 13 1 14 13 2 16 3 10 9 13 1 9 7 15 2 16 0 9 1 3 4 4 9 1 0 9 2 13 11 8
9 9 1 9 4 10 9 0 9 2
18 3 4 3 1 9 13 10 9 2 1 15 1 9 1 0 9 3 2
12 1 0 15 4 11 11 13 0 9 1 9 2
6 13 12 9 9 3 2
15 15 4 0 14 13 1 7 0 14 13 0 1 9 9 2
33 10 0 9 1 9 13 1 2 16 10 0 9 1 0 9 2 3 12 9 2 3 4 13 3 13 1 14 13 10 0 1 9 2
18 15 13 1 10 9 10 3 0 9 3 2 3 3 4 13 9 9 2
2 3 2
18 2 10 0 13 3 9 1 15 2 7 3 13 3 15 1 4 0 2
6 3 4 9 9 13 2
10 7 3 1 9 1 13 9 1 11 2
21 15 4 3 13 10 9 1 2 16 9 4 13 0 9 3 12 9 1 9 9 2
15 9 11 11 7 9 11 11 4 13 10 9 14 13 9 2
31 9 13 3 1 9 2 7 1 11 7 11 13 10 0 9 1 14 13 0 1 0 9 2 3 1 10 0 9 1 9 2
13 15 4 15 3 2 15 13 15 1 9 1 15 2
51 0 9 1 10 9 4 13 3 3 1 12 2 1 9 10 9 2 15 9 4 13 10 0 9 2 3 11 9 2 1 12 2 7 1 4 13 10 9 1 10 9 7 9 2 15 4 13 1 3 2 2
11 15 9 10 9 1 11 9 3 0 9 2
27 1 9 13 15 10 9 3 1 10 9 2 7 1 9 3 1 9 13 15 3 2 16 15 3 4 3 2
13 2 10 9 7 15 13 15 2 15 4 15 13 2
28 10 9 1 9 9 4 9 12 13 9 1 9 2 3 3 1 9 9 13 9 2 10 9 9 1 11 9 2
9 7 3 13 3 15 2 15 13 2
42 2 9 4 4 3 0 1 9 3 16 10 9 13 15 2 2 13 11 11 2 3 4 9 1 10 0 9 1 11 11 11 1 11 2 3 1 10 9 1 11 11 2
10 11 11 2 11 12 2 12 11 11 2
18 9 1 9 9 2 11 12 1 11 2 13 3 10 9 1 12 9 2
6 9 4 3 3 9 2
15 2 15 13 0 2 16 9 13 10 0 9 9 1 3 2
25 15 13 10 0 9 1 9 10 12 9 1 11 1 12 9 1 14 13 10 0 9 1 0 9 2
33 3 4 15 4 0 0 9 2 16 11 13 3 13 2 16 13 15 3 10 9 1 9 2 13 15 14 13 10 9 1 10 9 2
8 1 9 9 4 15 4 3 2
20 11 11 4 4 3 1 14 13 11 9 2 7 3 4 15 13 1 9 2 2
74 15 4 10 9 2 16 3 13 7 13 10 0 9 2 16 10 0 2 9 2 4 13 2 15 4 3 10 0 9 2 16 10 3 13 9 4 0 2 13 1 10 10 9 2 15 4 3 13 1 2 16 15 3 4 13 10 9 1 10 0 9 2 7 3 13 1 2 16 15 13 1 15 15 2
27 9 7 9 1 11 9 2 11 11 11 2 4 3 3 13 9 1 14 13 2 16 10 0 9 13 9 2
22 9 4 9 9 1 14 13 0 9 1 9 2 7 3 13 3 9 1 14 13 9 2
19 10 9 9 3 2 3 1 9 12 9 2 13 10 0 9 11 11 3 2
5 11 13 1 9 2
8 11 11 2 11 12 2 12 11
5 7 15 13 3 2
41 16 10 9 4 0 2 15 4 11 11 2 2 13 15 0 9 2 16 15 8 3 1 2 16 10 9 2 15 13 1 10 0 9 2 3 1 0 9 4 0 2
41 2 9 4 13 3 1 9 1 9 9 2 7 15 4 3 13 2 16 9 3 13 2 16 9 9 4 13 10 1 3 9 1 9 1 11 2 2 13 11 11 2
25 12 9 1 9 7 12 9 1 0 9 9 13 1 9 2 16 3 12 7 12 9 13 1 9 2
1 0
6 7 13 9 13 15 2
15 16 15 3 4 13 14 13 3 1 10 0 9 1 9 2
3 3 5 12
10 15 4 3 3 15 2 15 13 9 2
29 7 15 13 3 8 14 13 1 9 7 9 2 3 15 13 1 14 4 0 2 16 9 4 0 2 2 13 15 2
10 2 4 15 3 13 3 2 13 11 2
29 15 4 4 0 2 16 15 3 13 1 8 7 9 9 1 9 2 7 0 2 16 15 3 4 13 1 9 9 2
10 1 10 9 13 10 9 1 0 9 2
15 15 4 0 1 2 16 15 3 15 13 3 0 10 9 2
7 3 4 4 3 1 9 2
7 14 13 9 7 9 3 2
25 3 3 3 13 13 10 0 9 2 3 15 1 10 0 9 2 15 4 13 1 9 2 13 9 2
28 1 9 1 10 9 4 9 3 13 1 9 2 7 15 4 0 1 14 13 2 3 0 15 13 3 1 15 2
47 10 0 9 1 11 11 3 3 1 11 4 3 4 13 1 9 2 8 2 2 16 15 4 13 0 9 7 3 13 9 1 10 0 9 1 10 9 1 9 2 15 13 13 10 3 0 2
14 15 13 12 1 9 2 15 4 3 3 0 2 3 2
21 9 0 9 1 9 13 10 3 0 0 9 10 9 0 9 2 16 9 4 3 2
16 7 3 13 15 16 1 9 1 9 2 15 13 10 0 3 2
5 12 9 4 13 2
25 2 15 4 3 4 13 2 13 15 1 9 2 2 7 15 4 3 3 4 10 0 1 15 15 2
25 2 0 13 2 15 4 0 2 16 15 4 3 1 14 13 3 1 10 9 16 15 4 12 9 2
35 15 13 3 3 2 15 4 4 13 15 13 2 16 15 1 3 0 9 2 3 3 1 10 0 2 3 4 3 0 2 2 13 11 11 2
35 1 9 13 11 11 1 11 7 13 3 10 0 9 9 1 0 9 13 2 16 15 13 1 11 1 2 11 11 2 1 3 12 9 3 2
12 3 13 15 3 1 9 7 4 13 10 9 2
32 15 13 12 9 1 9 2 11 2 1 11 11 9 1 11 2 15 4 9 2 9 2 9 2 9 2 1 9 2 7 11 2
21 2 16 15 4 3 3 0 2 15 4 13 2 7 15 13 3 13 10 9 2 2
7 13 15 10 9 1 9 2
10 15 4 4 3 1 1 9 2 9 2
40 15 13 9 1 10 9 3 1 9 1 9 2 15 1 0 9 13 10 0 9 1 9 2 15 3 1 10 0 9 4 13 2 16 9 4 13 1 10 0 2
13 16 9 1 11 13 10 0 9 13 11 11 9 2
2 0 2
10 2 15 4 3 15 2 1 4 9 2
23 3 3 4 8 13 1 10 0 9 1 3 12 8 9 2 16 9 4 13 1 13 9 2
24 15 4 1 11 11 11 4 13 1 9 1 9 12 2 3 11 13 1 10 9 1 10 9 2
15 14 13 9 1 10 0 9 7 9 1 10 9 1 9 2
9 15 13 3 0 1 12 0 9 2
5 15 4 3 0 2
34 9 1 0 9 13 10 0 9 12 2 16 11 1 9 1 10 0 9 0 13 2 2 7 3 4 15 13 9 1 14 13 9 3 2
32 1 10 9 1 12 9 13 3 11 9 10 9 0 9 1 10 9 2 15 13 1 9 1 11 11 2 11 11 7 11 12 2
31 1 9 12 13 11 11 1 11 9 7 13 0 9 9 1 11 1 11 2 11 2 3 15 13 14 13 9 1 9 3 2
20 7 15 13 3 1 14 13 10 9 1 10 9 1 2 16 15 13 1 9 2
23 9 4 10 0 9 2 1 9 4 1 14 13 0 9 1 2 16 11 9 13 1 9 2
19 11 8 8 2 8 8 8 2 8 8 8 8 8 2 8 8 8 8 2
13 3 4 10 0 0 9 3 1 9 1 9 2 2
25 16 9 1 10 2 9 2 4 13 1 13 9 2 4 8 13 1 10 0 9 1 3 8 9 2
16 3 4 15 3 2 15 3 4 13 10 9 1 14 13 3 2
2 11 2
9 2 7 2 11 2 13 2 11 2
31 9 1 14 13 10 0 9 1 2 0 9 2 13 1 0 9 1 2 9 2 2 7 13 15 3 1 9 1 9 9 2
9 9 1 9 13 1 10 13 9 2
34 0 13 2 3 0 15 4 13 14 13 3 2 7 16 15 13 10 9 9 1 10 9 7 13 1 9 1 9 2 4 9 0 3 2
44 3 1 11 4 9 3 3 0 1 11 11 0 9 2 0 9 1 11 2 2 3 15 13 1 10 9 1 9 7 9 2 7 9 1 10 9 2 1 10 0 7 0 9 2
28 9 1 9 7 9 4 1 0 9 13 1 10 0 0 9 1 10 9 2 1 15 4 3 0 14 13 1 2
18 2 15 13 15 3 3 1 1 0 9 2 3 15 13 15 3 3 2
29 10 9 13 2 16 15 13 2 15 13 3 1 10 0 9 2 7 15 13 15 15 3 1 9 7 13 1 15 2
7 1 9 1 9 13 11 2
14 7 2 6 2 7 2 15 13 3 3 1 15 3 2
41 1 11 13 15 2 16 3 10 0 9 1 9 4 0 2 7 3 13 9 14 13 1 10 0 2 9 2 7 1 10 9 14 13 3 1 10 0 9 1 9 2
18 15 13 11 11 1 10 9 1 11 2 3 15 3 13 1 9 9 2
39 2 16 15 1 0 9 9 13 1 14 13 9 9 1 2 16 9 7 9 3 4 13 15 1 10 0 9 2 4 15 13 10 0 9 2 2 13 9 2
3 2 11 2
21 15 4 3 3 13 2 16 11 11 11 1 9 9 10 0 9 4 13 9 9 2
1 5
27 7 15 4 9 2 16 11 9 3 4 13 3 1 12 9 1 9 1 2 16 0 9 13 3 1 9 2
26 13 9 9 2 4 11 13 1 10 0 9 1 1 10 9 14 13 10 9 1 14 4 13 1 12 2
54 9 1 9 9 2 9 11 11 11 2 13 1 9 2 16 10 9 2 16 9 3 13 2 4 13 10 9 1 2 16 3 1 10 0 9 13 10 9 2 15 2 3 7 3 13 2 16 0 9 3 13 15 2 2
9 13 3 10 9 1 14 13 9 2
17 14 13 7 13 3 1 10 0 9 7 10 0 9 4 3 0 2
10 1 0 9 4 9 3 13 1 9 2
22 9 9 2 11 11 2 4 3 3 3 3 1 2 16 3 4 13 9 1 0 9 2
17 0 9 4 13 10 9 1 14 13 9 1 10 0 2 0 9 2
31 2 15 13 3 1 9 2 3 15 4 13 3 1 10 9 2 7 3 15 4 13 9 1 9 2 13 13 9 1 9 2
5 11 9 2 9 2
22 1 10 0 2 9 4 13 9 1 14 13 2 16 15 13 1 10 9 1 9 9 2
33 1 9 13 9 1 14 4 15 1 10 13 9 9 2 9 13 1 9 7 9 2 9 1 9 2 9 1 9 7 9 2 3 2
10 15 13 3 1 11 2 11 0 9 2
7 15 13 1 9 12 9 2
5 9 2 13 15 2
9 3 4 15 13 0 0 9 3 2
3 9 1 9
21 15 13 2 16 10 3 0 9 9 13 3 2 1 15 13 13 2 7 15 13 2
11 2 15 4 0 2 2 13 15 0 2 2
28 15 4 13 2 16 15 3 3 4 10 9 2 7 10 1 9 0 9 2 15 4 13 9 1 9 1 9 2
6 13 3 1 11 1 12
37 7 9 4 3 4 10 9 2 9 7 3 3 9 2 16 3 1 11 4 13 9 3 1 14 13 0 9 2 10 0 9 2 0 9 7 9 2
40 7 3 1 11 11 3 1 0 9 13 1 10 0 9 3 9 1 9 1 9 2 11 11 2 1 9 2 13 15 3 3 0 9 1 10 9 2 13 9 2
20 7 10 0 9 1 12 9 1 9 1 10 0 2 12 9 3 1 15 13 2
25 15 13 3 3 1 14 13 11 9 2 7 3 4 15 4 10 0 1 13 10 0 9 1 9 2
14 10 0 9 13 1 9 1 0 9 1 9 1 11 2
10 11 4 4 0 2 16 15 13 9 2
20 7 1 3 13 9 13 9 10 0 9 2 9 2 1 10 0 2 9 2 2
20 7 15 13 15 3 1 2 7 15 4 3 3 3 13 10 2 3 12 9 2
21 3 0 2 7 10 0 1 9 4 13 3 3 1 14 13 2 16 9 4 0 2
8 3 3 4 15 3 13 15 2
26 13 12 9 9 2 12 9 9 7 12 9 3 0 9 7 13 9 1 9 2 16 0 4 3 13 2
8 15 4 10 0 9 1 9 2
32 3 9 11 11 13 9 1 11 11 1 10 0 9 1 11 11 2 15 15 3 3 13 1 9 14 13 1 10 0 9 2 2
29 1 15 1 10 9 4 15 13 10 9 1 10 0 11 11 1 9 1 9 2 9 1 9 7 10 9 1 9 2
5 2 13 15 15 2
10 15 13 2 15 3 4 10 9 2 2
24 2 6 2 15 4 3 13 15 1 15 2 7 15 4 3 0 7 13 3 1 0 10 9 2
16 9 2 15 13 1 10 9 2 4 4 13 3 2 13 15 2
36 15 13 2 16 10 12 0 9 1 11 2 15 13 1 9 1 11 1 11 1 11 1 11 1 10 9 1 9 2 4 13 3 3 1 9 2
29 1 3 3 0 15 13 15 2 13 11 0 9 1 2 16 9 2 16 15 4 0 2 13 3 3 1 3 0 2
21 15 13 1 9 1 9 1 10 0 2 1 9 3 4 13 9 1 3 0 1 2
40 10 0 9 1 15 12 13 3 2 16 11 11 1 11 11 9 1 9 12 4 13 1 10 0 9 9 2 3 1 2 16 9 0 9 9 11 11 4 13 2
11 15 13 3 13 2 7 15 13 1 15 2
24 15 13 15 1 2 3 0 2 2 16 10 9 13 10 9 2 3 4 0 1 10 0 9 2
14 0 4 9 1 11 1 11 13 3 1 2 13 11 2
33 2 15 13 15 10 9 2 2 13 15 2 7 13 3 2 16 15 3 4 0 3 2 7 16 15 3 4 13 2 0 2 9 2
9 2 15 4 13 1 11 0 9 2
15 3 1 12 9 13 15 9 2 13 7 0 0 1 9 2
12 11 13 3 2 16 15 13 10 0 9 3 2
27 11 9 13 1 0 9 1 10 0 9 1 11 2 7 9 12 4 3 12 1 10 13 12 9 4 0 2
26 1 10 0 9 3 1 9 13 15 9 1 9 2 15 1 10 0 7 15 9 4 4 13 1 9 2
16 1 9 1 9 9 2 13 0 9 3 2 3 1 12 9 2
32 1 9 1 10 0 9 1 9 13 3 11 11 12 9 12 9 0 9 2 15 15 3 4 13 1 10 9 9 1 9 9 2
26 12 0 9 1 9 9 4 13 0 9 1 9 2 16 9 1 10 9 13 10 0 0 8 7 9 2
13 2 15 13 3 0 9 1 9 2 13 11 3 2
14 9 11 13 1 9 1 11 1 15 1 9 13 9 2
13 9 13 2 16 9 4 3 3 3 0 1 9 2
13 2 15 4 13 15 2 2 13 10 0 1 9 2
18 0 2 7 0 7 0 9 1 9 1 0 9 7 0 0 0 9 2
9 11 7 11 9 4 0 9 13 8
9 7 3 4 9 3 10 0 0 2
45 16 9 9 7 9 3 4 13 2 13 15 3 2 16 10 9 9 3 3 4 10 9 1 9 2 15 9 3 13 3 3 3 1 10 9 3 7 3 1 1 3 0 10 9 2
41 3 4 15 15 11 9 2 16 15 4 3 3 13 15 15 2 15 3 13 2 2 13 11 11 2 15 13 15 3 1 9 2 16 10 2 13 9 2 13 9 2
13 3 4 15 9 2 11 11 2 15 13 1 9 2
30 1 10 13 9 2 3 4 4 10 9 2 13 15 1 11 0 9 2 16 10 0 0 9 3 4 13 1 0 9 2
8 0 9 13 1 9 7 9 2
11 15 13 10 0 9 1 11 1 9 2 2
38 13 15 13 15 2 16 10 0 9 1 9 3 4 13 10 0 9 3 1 10 9 7 10 9 13 1 13 9 13 1 14 13 9 1 0 0 9 2
21 11 11 13 3 1 9 2 7 15 13 15 3 3 2 2 13 11 11 1 11 2
22 15 13 3 1 9 7 13 3 7 13 1 10 0 2 15 4 13 15 1 9 9 2
27 9 1 9 2 1 3 4 10 0 9 2 4 15 3 13 1 11 11 0 9 2 9 1 12 9 2 2
19 10 0 13 1 9 9 1 10 9 2 10 9 3 1 9 1 1 9 2
18 0 15 2 15 3 13 3 0 9 2 16 15 4 13 1 0 9 2
27 9 13 0 9 2 16 9 7 9 2 0 9 15 13 1 9 3 2 4 13 1 10 0 9 1 11 2
30 2 13 15 1 0 0 9 2 2 13 11 11 2 15 1 11 3 13 9 2 1 10 9 1 9 11 11 11 9 2
7 7 15 13 15 3 3 2
32 15 4 3 0 2 16 0 9 4 13 1 10 9 2 16 10 0 7 0 9 1 10 0 9 13 9 1 0 9 7 9 2
18 11 13 3 1 9 2 7 11 13 9 3 13 1 0 9 1 11 2
3 2 6 2
36 15 4 3 0 2 16 9 1 11 7 3 3 11 9 1 11 13 9 1 10 0 0 9 1 10 9 1 14 13 0 9 13 10 0 9 2
8 11 11 13 10 9 1 9 2
19 16 15 4 0 2 13 15 1 9 1 0 9 7 13 15 1 9 9 2
23 10 0 9 4 12 9 2 15 4 13 10 0 9 2 15 13 10 9 1 12 9 9 2
13 15 13 1 15 1 10 0 9 1 10 0 9 2
22 7 1 15 13 3 10 0 9 1 14 13 9 7 14 4 13 15 1 10 0 9 2
15 1 9 3 1 11 13 15 1 3 14 13 1 0 9 2
5 9 13 1 9 2
22 7 3 13 15 1 2 16 9 3 13 3 7 3 13 1 3 11 11 7 11 11 2
22 9 13 3 10 0 9 1 0 9 9 1 14 13 15 1 0 9 2 2 6 9 2
10 13 0 7 13 9 7 0 9 3 2
24 7 15 13 1 10 9 1 9 9 2 3 3 0 1 15 2 3 4 3 1 14 13 9 2
18 2 16 15 13 9 2 4 3 13 1 14 13 9 2 2 13 15 2
12 15 4 3 13 1 9 2 15 13 10 9 2
12 9 8 9 13 3 10 9 1 9 1 9 2
52 11 11 13 9 1 9 3 9 1 11 11 9 1 2 16 15 1 9 12 1 9 1 9 4 4 13 2 15 15 15 13 10 2 9 2 1 2 16 9 4 13 2 7 16 15 3 4 13 10 0 9 2
47 2 13 15 15 9 10 9 9 1 10 0 9 2 13 15 0 10 9 2 15 13 1 10 0 9 2 7 10 9 9 3 2 13 9 11 11 2 3 4 9 1 11 11 9 1 11 2
19 15 13 2 15 4 3 3 0 7 3 0 14 13 9 1 11 11 11 2
2 10 9
40 9 1 10 13 9 4 3 4 0 2 16 9 4 13 2 16 15 4 13 16 3 13 9 1 10 9 1 10 0 9 7 3 4 13 15 2 1 4 0 2
5 15 13 9 3 2
11 11 11 4 3 1 14 13 0 9 9 2
21 7 9 9 13 1 9 2 2 7 10 9 1 9 2 2 7 3 13 3 9 2
19 15 9 13 1 3 10 9 2 3 15 4 0 7 13 1 10 0 9 2
20 15 4 1 0 3 2 15 4 13 14 13 15 7 13 9 1 10 0 9 2
29 11 11 9 13 1 9 1 9 9 9 1 9 1 9 2 1 15 13 4 4 15 1 10 3 13 9 1 11 2
19 9 4 1 10 9 9 1 10 9 2 15 4 13 2 1 9 0 9 2
23 9 1 9 4 13 15 2 15 4 3 3 13 2 16 15 4 4 3 3 0 1 3 2
16 2 15 4 3 0 2 7 9 4 13 12 9 1 10 9 2
4 3 13 9 2
7 9 2 9 2 12 8 2
16 15 13 10 9 1 14 13 2 16 9 3 13 10 9 3 2
68 15 4 9 3 2 7 10 11 1 0 9 1 9 1 9 9 2 7 3 3 15 0 1 2 16 15 3 3 13 3 1 10 9 1 9 1 10 0 9 8 2 4 13 10 3 0 9 3 3 1 10 9 0 0 9 2 15 4 13 10 0 9 9 1 2 11 2 2
10 11 13 1 9 3 1 10 0 9 2
3 0 1 9
5 11 4 3 13 2
16 10 9 13 3 16 9 4 13 7 3 2 3 8 10 9 2
7 15 4 15 13 11 1 2
10 3 1 15 4 13 1 9 1 15 2
12 10 0 13 3 3 13 1 9 7 9 2 2
23 10 0 9 13 3 1 10 10 9 2 9 2 3 1 9 12 9 9 1 10 0 9 2
9 9 4 13 10 0 9 1 9 2
1 9
14 15 4 13 10 0 9 13 1 9 7 13 3 15 2
7 3 4 15 3 13 15 2
3 9 7 9
17 10 9 13 1 12 7 12 9 16 15 4 4 13 10 0 9 2
8 13 9 1 9 7 13 3 2
8 9 13 0 1 9 7 9 2
13 1 11 9 13 9 1 9 1 9 10 0 9 2
8 0 1 15 0 9 13 3 2
14 10 0 9 13 1 14 13 10 9 1 10 0 9 2
29 3 4 15 13 1 14 4 13 15 10 0 9 2 13 9 14 13 1 15 13 3 1 9 1 9 3 15 13 2
9 15 4 9 1 9 7 9 2 2
6 10 0 9 4 13 2
9 2 15 4 13 3 2 1 9 2
10 10 9 1 9 3 13 1 0 9 2
24 11 4 3 13 3 2 7 14 13 3 1 0 9 2 13 14 13 1 14 4 13 1 9 2
8 11 11 4 15 1 10 0 2
20 11 4 1 10 9 3 13 10 9 3 1 9 2 16 15 13 10 9 9 2
44 3 15 4 13 1 0 9 1 9 2 2 15 4 13 3 1 9 9 2 10 9 2 9 7 9 9 1 10 9 2 7 10 9 4 13 3 1 2 16 15 13 1 9 2
37 2 9 13 3 1 14 13 3 13 0 10 0 9 2 7 15 4 3 13 9 3 1 9 2 16 15 3 13 9 1 9 2 2 13 11 11 2
11 9 4 3 0 2 16 0 4 13 3 2
24 15 4 3 3 0 2 7 1 10 9 13 3 3 0 3 2 16 15 13 3 1 9 2 2
12 15 13 10 0 9 12 2 16 11 4 13 2
10 2 0 9 13 3 3 8 1 9 2
34 11 4 1 9 3 4 13 15 1 0 9 7 9 2 7 3 11 9 2 15 0 13 13 1 9 0 9 2 4 3 13 1 13 2
39 15 4 3 3 13 2 16 3 12 0 9 13 9 9 1 11 2 10 9 2 15 13 4 10 0 1 9 2 1 14 13 15 9 0 9 1 9 1 2
40 3 3 11 4 1 9 3 0 2 7 9 1 11 13 1 9 14 13 10 9 1 11 7 11 1 0 9 2 15 15 13 15 1 9 1 10 0 9 9 2
19 11 11 13 9 9 2 7 4 3 1 9 9 10 0 0 9 1 9 2
24 3 1 14 13 15 3 1 10 0 9 2 3 1 10 7 0 9 4 3 0 7 3 0 2
34 1 0 9 1 3 10 0 1 10 0 9 4 15 3 4 0 14 13 9 0 1 14 13 1 9 2 8 8 3 13 9 1 9 2
61 3 1 11 7 11 4 3 1 10 0 9 9 13 9 1 13 12 9 9 2 7 1 0 9 4 11 2 16 10 0 9 3 13 15 2 13 10 9 1 12 9 9 1 10 0 9 11 2 1 9 1 10 12 9 13 9 1 10 0 9 2
3 13 15 2
20 15 13 3 2 7 15 4 13 1 2 16 15 3 13 3 1 9 1 9 2
28 3 3 13 15 9 1 9 2 16 9 1 9 3 4 13 1 1 12 2 7 16 9 3 1 11 4 13 2
3 1 9 2
24 0 7 0 9 13 1 9 3 14 13 2 16 11 11 9 1 9 4 3 1 14 4 3 2
9 3 1 10 9 7 1 10 9 2
12 15 4 10 0 9 9 3 2 15 4 0 2
41 16 3 1 9 3 13 3 13 2 0 9 1 11 11 2 4 15 3 9 9 14 13 2 16 10 13 9 1 9 4 0 3 1 14 13 2 16 11 4 9 2
13 3 1 10 0 9 4 15 13 9 1 9 11 2
9 9 4 1 10 9 13 3 0 2
21 1 12 10 0 9 4 10 0 9 1 9 13 0 9 2 16 9 4 10 9 2
13 3 11 11 11 2 15 13 0 9 2 4 13 2
29 11 7 11 2 15 4 13 1 10 9 3 1 9 13 1 10 0 9 7 13 3 1 10 0 9 1 0 9 2
27 10 9 3 4 15 13 3 1 10 0 9 2 2 15 4 10 3 0 9 1 15 2 10 9 1 11 2
13 2 15 13 2 15 4 4 3 1 0 9 0 2
14 9 13 10 0 9 9 1 11 2 15 4 13 3 2
10 11 13 10 0 9 1 9 1 9 2
12 7 0 9 13 1 0 9 1 10 0 9 2
1 9
22 11 2 11 2 4 4 3 13 1 9 2 16 11 7 15 2 8 8 2 4 15 2
16 2 3 4 0 1 15 4 3 1 9 1 1 12 9 3 2
17 15 4 3 13 2 16 9 4 10 9 1 10 0 9 0 9 2
18 15 13 1 0 11 11 2 3 9 4 13 1 0 9 1 10 9 2
21 9 13 3 13 7 4 3 4 3 2 7 15 4 3 13 7 1 10 9 13 2
23 15 4 3 0 1 12 9 2 7 15 4 13 2 9 4 0 7 0 2 2 13 11 2
7 3 13 15 3 1 9 2
21 13 0 9 7 8 7 9 3 7 13 3 1 12 9 9 3 2 16 9 13 2
2 9 2
2 9 2
10 3 13 15 3 16 15 4 13 0 2
18 0 9 4 13 2 7 9 4 3 13 2 3 11 13 3 0 9 2
14 9 9 11 11 13 12 9 9 7 10 9 12 9 2
12 1 9 4 15 13 9 1 9 7 9 3 2
14 1 10 12 9 1 2 11 2 4 15 13 1 9 2
23 15 13 2 16 0 9 13 9 1 9 2 16 15 1 0 4 13 15 1 14 13 9 2
12 9 13 9 1 10 0 9 9 2 10 0 2
22 10 0 9 4 3 3 0 7 13 1 15 14 13 1 2 7 15 13 15 3 0 2
13 15 4 9 7 13 12 9 1 9 1 9 9 2
18 10 9 2 1 9 2 13 1 11 2 9 2 13 9 7 13 9 2
16 10 0 9 1 11 13 1 9 2 15 13 9 0 1 9 2
18 15 13 1 0 9 1 15 2 7 15 13 1 9 7 9 1 15 2
10 11 11 11 13 15 8 9 1 11 2
35 1 10 9 1 9 3 1 15 13 11 2 7 1 9 1 15 13 10 0 0 9 2 15 3 13 3 1 14 4 10 9 1 10 9 2
33 1 11 13 1 15 8 10 9 1 10 9 1 12 8 2 10 0 7 0 9 2 15 13 2 16 11 3 3 4 13 0 9 2
7 9 4 3 3 13 3 2
17 11 4 13 1 9 1 9 7 13 3 9 1 9 1 0 9 2
30 1 9 4 15 1 10 0 13 8 9 4 13 10 0 13 9 3 2 3 1 10 9 9 2 13 3 3 13 13 2
39 9 13 10 0 9 1 14 13 2 16 15 2 15 13 9 1 7 13 3 13 9 2 13 0 3 0 9 1 14 13 10 9 1 9 1 9 7 9 2
6 8 5 8 9 5 8
24 2 15 13 1 2 16 9 7 9 1 9 3 13 1 15 7 13 15 3 2 2 13 9 2
30 9 4 3 13 2 16 9 1 9 1 9 3 7 3 4 13 1 10 0 9 2 16 3 13 9 1 9 7 9 2
23 2 15 13 1 9 2 16 3 3 4 13 10 9 1 10 9 7 15 2 2 13 9 2
4 7 3 3 2
10 2 3 13 15 1 9 1 10 9 2
39 9 4 9 2 7 15 4 0 2 16 11 4 0 2 16 15 4 3 13 1 9 2 16 15 13 10 0 9 1 0 9 1 10 3 0 2 0 9 2
18 3 9 13 9 1 2 16 10 9 3 3 4 4 10 9 1 9 2
22 7 15 13 3 0 1 9 2 15 15 4 13 14 13 1 12 9 0 9 7 9 2
16 10 0 2 9 2 13 1 14 13 1 11 7 3 1 11 2
13 3 13 15 9 1 9 2 1 4 0 1 15 2
26 10 8 9 4 0 7 4 3 13 3 2 9 2 15 4 3 4 0 14 13 10 0 3 13 9 2
25 9 1 10 0 9 4 1 10 13 9 1 0 9 1 9 13 10 9 1 10 0 9 1 11 2
18 7 15 13 1 14 13 9 3 2 1 13 15 0 13 1 0 9 2
1 9
47 9 1 9 1 10 2 0 0 9 2 4 3 13 15 1 2 16 15 4 13 1 0 9 1 10 9 2 7 16 15 3 4 0 14 13 0 0 7 0 9 1 14 13 10 0 9 2
32 1 15 4 2 10 0 2 13 3 3 2 1 15 1 10 0 9 1 15 1 10 9 0 9 2 16 15 13 15 1 9 2
25 10 0 9 9 2 11 11 2 13 3 2 16 3 3 4 4 13 0 1 10 12 9 1 11 2
13 1 10 0 9 4 9 0 14 13 1 9 9 2
25 9 13 2 16 15 3 4 9 9 14 13 10 9 7 13 0 10 0 9 2 9 9 4 13 2
15 9 13 1 9 1 10 9 1 12 9 1 10 0 9 2
18 10 0 9 2 15 13 2 16 11 4 13 9 1 10 11 11 9 2
11 10 9 4 3 3 13 1 9 0 9 2
50 9 1 10 12 0 9 2 9 7 11 2 13 10 0 9 11 2 15 13 9 3 7 3 13 1 9 7 10 9 2 15 15 13 1 2 0 9 2 2 9 2 15 10 9 13 1 9 9 1 2
15 11 13 2 1 15 13 2 7 3 13 15 3 1 15 2
22 16 15 13 3 2 13 15 2 2 15 13 3 1 10 9 2 7 15 4 3 3 2
17 9 11 11 13 3 9 3 0 2 16 15 4 13 10 0 9 2
14 1 9 13 9 3 3 2 7 10 13 9 13 9 2
20 9 13 2 15 4 13 10 0 0 9 11 11 1 9 1 9 1 12 9 2
16 3 1 15 3 4 13 9 9 2 4 15 3 13 1 9 2
7 2 9 2 4 15 13 2
16 3 3 3 1 9 1 9 13 13 7 9 13 13 1 9 2
38 7 15 13 3 1 10 12 9 2 15 3 4 13 3 1 11 1 9 1 11 2 16 15 3 13 14 4 13 1 0 9 1 13 1 9 1 11 2
10 3 13 15 2 15 4 13 15 1 2
8 15 4 3 13 3 1 9 2
11 9 1 11 11 12 11 9 2 9 9 2
7 9 1 11 13 1 9 2
10 1 9 4 15 13 15 1 12 9 2
4 4 15 13 2
31 11 9 4 13 2 16 0 9 1 0 9 12 4 4 13 1 15 13 2 16 3 3 4 13 1 10 9 1 12 8 2
32 7 3 1 15 4 10 9 2 7 11 4 10 10 9 2 7 11 10 0 2 13 15 3 1 3 4 13 10 9 10 9 2
6 15 4 3 9 1 2
9 0 9 13 12 9 1 12 9 2
8 9 4 3 10 0 1 9 2
10 1 12 9 4 11 11 3 1 11 2
7 3 4 13 0 10 9 2
10 10 12 9 13 1 9 1 12 9 2
8 1 10 9 1 10 9 9 2
25 15 2 15 13 1 9 1 9 2 13 15 3 2 7 3 13 15 3 1 9 1 3 10 9 2
11 7 15 13 3 3 0 9 1 14 13 2
6 3 13 15 1 9 2
14 2 15 4 10 9 13 1 10 0 0 7 0 9 2
5 9 2 11 11 2
22 10 9 13 3 10 9 1 12 0 9 3 1 9 1 13 0 7 0 9 2 11 2
26 3 13 15 3 1 9 7 3 1 0 9 2 3 9 12 9 1 9 12 1 12 9 13 7 13 2
24 3 4 15 1 9 4 0 1 12 9 1 10 9 9 2 11 11 2 1 10 0 9 11 2
43 7 1 10 9 2 16 15 4 4 0 14 13 8 7 9 1 10 0 9 1 9 3 1 10 9 9 7 3 1 10 9 2 16 0 9 7 9 3 4 13 1 11 2
11 1 10 9 4 15 3 13 1 12 9 2
29 11 13 1 10 0 9 1 10 9 2 10 0 9 11 2 10 0 9 1 9 2 7 3 1 9 1 12 9 2
2 9 9
8 13 0 9 1 9 1 0 2
43 3 3 3 2 3 11 3 13 11 11 9 12 9 1 9 1 1 12 9 2 9 2 2 7 3 1 9 13 3 1 14 13 0 9 1 9 2 1 1 12 0 9 2
10 2 4 15 0 2 2 13 15 3 2
9 1 9 4 15 1 0 9 0 2
10 1 9 13 13 12 9 1 12 9 2
28 11 11 2 9 1 9 1 9 2 11 11 2 9 1 11 2 11 11 2 9 1 9 2 12 9 2 0 11
45 1 10 0 12 9 4 15 13 15 3 12 9 2 10 9 9 1 9 1 9 2 7 10 0 9 1 9 1 15 2 15 3 4 13 2 1 16 10 0 9 13 10 8 9 2
23 2 15 13 15 12 9 14 13 9 1 0 9 2 16 15 13 11 11 0 9 1 12 2
12 11 4 13 1 9 1 9 11 1 11 11 2
10 9 13 9 2 7 3 4 13 9 2
9 8 1 9 1 9 13 9 9 2
6 4 15 3 3 0 2
18 7 3 10 9 2 15 15 4 13 1 9 9 2 4 11 13 1 2
13 1 9 13 0 9 10 13 9 1 1 10 9 2
6 2 9 4 4 0 2
50 10 13 0 9 2 11 11 2 12 2 15 1 9 4 13 1 10 0 9 11 2 13 1 10 9 1 9 2 16 15 3 4 13 9 1 9 1 10 9 2 15 4 13 15 3 1 10 13 9 2
40 7 1 10 9 2 15 15 4 13 1 9 2 13 3 3 3 0 1 10 9 1 2 16 11 11 4 4 13 15 0 2 2 13 9 1 11 2 11 11 2
14 9 1 12 4 13 1 9 0 0 9 3 1 9 2
15 2 13 15 3 2 11 4 10 3 0 9 2 13 15 2
35 3 13 15 2 16 9 0 9 1 0 9 1 9 13 13 1 10 9 1 9 1 9 7 9 3 1 9 1 9 1 10 0 0 9 2
19 9 1 9 1 11 2 11 9 7 9 4 0 9 9 2 11 11 11 2
20 9 13 2 16 3 12 9 4 13 1 9 1 11 1 12 9 3 1 11 2
27 9 1 9 1 11 11 2 11 9 4 1 9 1 9 13 10 0 9 1 9 1 3 11 7 11 9 2
17 9 7 9 1 9 13 2 9 13 2 7 9 4 13 9 9 2
20 1 9 4 3 13 12 9 9 1 9 2 1 9 13 12 9 1 11 9 2
26 1 9 13 15 1 9 2 7 3 4 15 9 2 16 15 3 4 13 1 9 1 9 3 1 11 2
22 15 4 10 9 9 1 12 9 2 16 11 11 13 15 1 3 0 1 12 1 9 2
15 3 9 1 0 9 7 9 2 15 13 9 1 15 13 2
21 2 7 1 10 9 4 3 13 12 0 9 2 7 3 4 15 3 3 1 9 2
20 15 4 3 0 14 13 2 16 16 15 3 4 11 11 2 15 4 9 3 2
27 9 13 14 13 9 13 1 10 0 9 2 7 15 13 9 1 9 1 2 16 9 4 13 1 10 9 2
39 13 15 15 14 13 1 9 2 3 13 0 0 9 2 11 2 10 9 9 1 10 0 2 7 3 1 10 3 0 9 1 11 2 11 2 11 7 11 2
13 15 13 1 12 1 12 9 1 10 9 1 12 2
23 2 7 15 13 3 3 1 15 15 3 2 15 4 10 0 1 15 2 15 13 9 2 2
24 13 15 8 10 0 2 0 9 2 15 15 1 15 2 3 4 0 2 4 4 0 14 13 2
5 2 8 12 2 2
17 2 15 13 15 1 13 15 2 16 9 4 0 1 1 10 9 2
27 16 3 3 3 13 10 9 1 9 9 2 4 9 7 9 4 9 1 9 7 9 2 7 9 13 3 2
22 7 15 4 13 2 16 15 4 3 0 2 16 15 7 9 11 11 1 9 4 9 2
14 10 0 9 4 3 1 9 13 3 0 9 7 9 2
15 11 2 12 9 1 11 9 1 11 4 13 1 9 12 2
7 7 3 13 15 3 3 2
28 2 9 4 0 1 0 9 7 13 3 12 9 1 10 0 9 2 7 12 9 1 10 0 2 13 11 11 2
19 1 12 9 1 9 13 1 9 1 9 1 13 9 13 15 3 9 9 2
10 10 0 9 4 3 1 14 13 15 2
16 9 13 3 2 3 15 13 10 9 2 15 3 3 4 13 2
12 2 13 3 2 11 2 15 13 3 3 3 2
11 3 13 3 16 3 4 13 1 10 9 2
44 15 1 15 2 15 13 9 2 4 11 11 2 15 3 3 13 15 9 1 10 9 1 10 12 9 2 2 15 13 9 7 13 1 14 13 2 7 3 4 15 13 15 3 2
24 15 2 15 4 13 15 2 4 9 2 7 15 2 15 13 15 2 15 4 13 2 4 9 2
45 11 2 3 4 0 1 11 9 2 13 3 10 0 7 3 0 9 2 10 0 11 9 2 15 13 1 0 9 2 1 9 1 15 9 7 3 0 14 13 1 1 0 9 9 2
7 7 13 15 3 13 15 2
20 7 16 15 13 3 3 2 4 15 4 13 1 10 3 0 7 0 0 9 2
20 1 9 9 13 11 11 2 15 1 3 13 1 11 2 11 11 9 1 9 2
8 2 15 13 1 11 1 9 2
15 9 13 12 9 1 9 1 9 1 9 1 9 1 9 2
13 2 16 3 13 0 7 8 9 7 9 1 9 2
11 3 0 10 9 4 11 11 3 3 1 2
13 15 4 0 9 2 16 9 4 13 1 0 9 2
15 2 11 4 13 9 1 9 2 7 15 4 13 9 3 2
28 13 9 3 2 16 15 4 4 0 2 16 9 13 3 1 10 0 9 2 3 13 15 15 3 1 10 9 2
10 15 13 15 4 15 3 13 1 9 2
23 3 4 9 13 12 9 2 16 15 4 13 11 10 13 9 2 11 2 16 9 11 13 2
6 3 13 3 10 9 2
26 3 13 15 3 1 9 2 13 10 9 7 13 10 0 9 1 10 9 2 15 13 11 13 3 1 2
48 2 15 13 3 1 11 1 0 10 9 2 3 15 13 1 12 9 2 13 1 15 1 3 3 14 13 1 12 9 7 13 1 15 3 2 1 14 13 15 3 1 9 2 2 13 11 11 2
43 3 7 3 3 3 3 1 9 13 11 11 11 2 0 9 1 11 2 3 15 1 10 0 9 1 9 13 10 0 13 1 9 1 14 13 1 10 0 9 3 1 11 2
33 15 13 3 1 10 0 9 1 10 9 7 13 3 2 13 9 3 2 16 0 9 4 3 2 2 4 15 3 10 9 2 2 2
29 15 13 15 13 10 9 1 9 1 15 2 3 3 3 2 7 13 3 1 9 2 15 15 13 1 10 0 9 2
2 13 9
9 3 4 9 13 2 2 13 9 2
14 1 12 9 13 15 3 10 9 1 9 1 10 9 2
20 7 1 9 13 15 1 10 9 10 9 1 9 1 3 14 13 9 1 9 2
15 15 13 3 7 3 1 11 9 13 1 10 9 1 15 2
16 7 15 13 10 13 9 3 14 13 2 16 10 0 9 13 2
13 11 2 15 13 3 3 1 11 1 10 0 9 2
48 1 9 1 9 13 11 11 11 1 9 2 11 2 1 9 1 9 8 11 1 9 1 11 11 10 9 3 1 11 2 16 15 1 9 9 3 13 2 16 3 4 13 2 9 1 9 2 2
13 15 13 2 15 15 13 2 4 13 9 1 9 2
7 2 1 9 2 13 11 2
19 1 10 9 1 10 9 9 1 10 12 9 13 15 1 10 9 1 11 2
23 3 13 9 10 0 9 2 3 15 9 13 1 12 9 2 15 1 15 4 4 10 9 2
2 12 2
25 11 2 2 6 2 7 15 13 3 3 2 3 1 9 9 15 4 13 15 3 1 10 0 9 2
21 9 1 15 1 10 0 1 15 3 4 4 0 14 13 1 9 1 8 7 9 2
27 16 3 10 9 13 10 9 1 12 9 2 3 4 9 13 9 10 9 2 15 13 1 3 12 9 9 2
15 3 13 15 3 1 12 9 2 12 9 7 10 0 9 2
11 15 4 15 13 10 9 1 2 13 11 2
13 15 13 3 9 1 10 0 9 14 13 0 9 2
20 3 1 9 13 10 0 9 2 0 2 9 2 0 9 2 1 9 1 9 2
14 1 10 9 2 11 2 4 15 3 0 9 9 2 2
24 3 13 3 10 0 2 15 4 12 0 2 7 15 4 3 3 13 2 7 9 4 3 0 2
13 1 0 9 4 15 3 4 13 10 9 1 9 2
16 9 4 13 1 11 11 11 2 7 9 13 15 13 1 9 2
23 15 4 0 9 13 1 14 13 10 0 9 2 7 15 4 15 3 13 2 2 13 15 2
22 7 9 1 0 9 13 3 3 14 13 9 3 2 13 11 11 2 9 1 11 9 2
10 7 1 11 11 9 4 9 10 9 2
12 16 9 13 1 15 2 4 15 10 0 9 2
33 11 13 10 0 9 9 1 3 11 7 11 7 4 13 0 1 9 3 2 16 15 13 10 9 1 14 13 10 0 9 1 9 2
19 10 9 1 9 13 3 9 1 15 0 9 2 15 3 4 13 1 9 2
37 0 9 4 3 13 9 1 2 7 2 15 13 9 1 9 2 1 14 13 1 12 1 12 15 9 1 12 9 7 3 13 10 0 8 7 9 2
27 16 0 1 10 2 9 2 2 15 3 1 9 13 1 10 0 9 2 13 13 2 15 4 10 10 9 2
17 8 8 1 9 13 14 13 10 9 1 9 7 13 3 1 9 2
7 15 13 3 14 13 3 2
26 10 0 9 13 3 2 16 9 3 1 9 4 13 3 12 9 9 2 12 9 9 7 12 9 9 2
27 15 13 10 0 9 1 9 1 2 16 3 4 13 3 0 10 9 1 9 2 16 15 4 13 10 9 2
11 15 1 15 13 2 3 10 9 13 3 2
15 6 2 3 13 3 10 9 2 3 3 3 3 4 9 2
15 1 9 1 9 4 9 3 12 1 11 7 12 1 11 2
26 13 1 0 9 13 3 9 1 10 0 9 2 15 13 9 1 16 9 4 13 2 16 9 4 13 2
13 3 4 9 13 10 0 9 1 11 9 1 11 2
5 9 2 9 7 9
15 15 13 1 1 9 11 11 2 11 11 7 11 11 2 2
8 13 9 1 9 7 13 3 2
25 2 15 4 3 3 13 2 15 4 0 9 2 7 15 4 4 0 14 13 9 1 10 0 9 2
8 15 1 10 0 9 4 9 2
55 3 3 1 9 9 1 10 9 13 11 1 10 9 1 9 1 0 9 1 9 7 9 2 1 15 4 13 1 2 16 3 13 9 2 1 16 15 13 1 2 9 1 9 2 2 15 3 13 15 1 10 9 1 9 2
17 3 13 3 15 2 7 3 4 15 3 3 2 7 3 10 9 2
27 11 4 13 10 3 0 9 1 14 13 10 9 1 15 1 11 2 16 15 4 13 1 14 13 0 9 2
11 1 10 0 9 1 9 2 4 9 0 2
17 2 7 13 3 1 2 16 15 3 13 3 0 14 13 1 9 2
8 15 13 2 16 9 13 3 2
1 9
9 15 13 9 2 16 15 13 9 2
11 10 12 9 4 1 0 9 4 0 9 2
42 2 0 9 4 3 10 3 13 9 2 15 0 9 13 1 14 13 15 1 10 0 9 2 7 3 13 15 14 13 15 2 15 4 13 1 9 7 13 15 10 9 2
18 0 9 4 1 9 13 1 0 9 1 9 7 2 9 7 1 9 2
35 11 11 4 1 12 4 13 1 11 2 10 9 9 11 2 1 12 9 7 9 11 11 2 11 11 7 11 11 11 11 1 10 12 9 2
41 1 11 13 10 0 9 11 11 11 7 13 15 10 2 0 2 9 2 16 15 3 4 13 1 9 1 10 9 2 16 15 4 13 2 16 11 7 11 13 9 2
26 2 15 13 3 2 16 15 3 4 13 15 3 3 2 7 15 4 3 3 15 2 15 13 15 1 2
20 16 15 4 0 2 13 15 3 13 15 1 9 2 3 3 1 10 0 9 2
9 3 10 13 9 4 15 3 4 2
9 3 1 9 4 9 1 11 9 2
27 2 0 9 13 1 0 9 1 9 10 0 9 2 16 15 4 0 3 1 2 15 9 13 14 13 15 2
26 9 11 11 13 3 1 9 2 16 15 1 9 13 2 16 11 11 3 4 13 0 9 1 10 9 2
13 10 0 9 1 9 2 13 1 12 9 1 11 2
8 11 11 13 9 1 11 11 2
8 3 13 15 3 1 0 9 2
25 9 1 2 16 10 9 3 13 10 0 9 2 15 13 15 2 4 4 13 1 0 9 1 9 2
18 15 4 3 13 15 14 13 9 1 9 2 16 3 3 13 10 9 2
15 0 11 13 2 15 3 13 11 9 1 15 3 3 0 2
18 15 13 3 15 1 14 13 3 3 3 2 3 3 4 15 3 13 2
20 3 4 9 13 3 3 1 9 2 16 15 13 1 11 9 7 1 9 9 2
9 3 4 13 9 1 9 7 9 2
3 8 5 8
8 11 4 3 13 9 1 9 2
16 2 15 13 3 9 1 10 9 2 2 13 11 11 1 11 2
29 9 2 11 8 2 13 1 14 4 3 0 7 3 3 0 1 10 0 9 2 7 0 9 13 1 10 0 9 2
23 3 3 15 13 3 1 10 0 9 2 3 4 15 0 14 4 3 1 0 10 9 2 2
13 15 4 3 10 9 1 0 9 2 15 13 3 2
18 7 3 13 3 10 9 1 10 12 9 2 0 9 1 9 12 9 2
24 9 13 3 10 9 1 9 1 10 0 9 1 14 13 9 1 3 3 0 2 7 3 0 2
5 9 4 11 11 2
23 1 1 12 0 3 1 11 9 4 9 1 9 13 1 10 0 9 1 3 13 12 9 2
21 15 13 3 0 9 1 9 2 16 3 13 9 1 14 13 0 9 1 11 9 2
18 10 0 4 15 13 1 9 1 9 7 0 2 9 2 9 7 9 2
21 11 13 1 16 13 9 4 13 1 9 7 9 1 9 2 0 9 15 0 9 2
25 1 3 0 9 13 15 11 13 15 1 10 0 9 7 0 9 2 7 15 13 3 0 3 3 2
25 15 13 15 3 1 0 2 14 13 10 9 3 1 10 0 9 2 16 10 0 9 4 13 3 2
16 10 0 9 13 3 0 13 9 2 15 13 1 9 7 9 2
7 15 4 3 3 4 11 2
8 15 13 3 3 3 1 3 2
29 10 9 1 11 1 9 1 12 13 3 9 7 9 1 14 13 3 3 2 7 3 13 15 15 3 3 1 0 2
8 15 4 3 13 15 1 3 2
12 15 13 2 3 0 2 7 2 3 0 2 2
1 9
23 11 11 2 15 13 9 2 4 13 10 9 1 12 9 1 10 0 9 1 12 9 9 2
16 7 1 11 9 13 11 10 9 2 15 13 3 1 9 3 2
5 15 13 3 3 2
8 1 9 1 10 0 0 9 2
7 13 9 1 10 0 9 2
11 7 16 15 3 13 15 10 0 1 15 2
8 10 0 9 4 10 9 0 2
36 9 11 11 13 2 16 11 13 9 1 10 0 9 2 11 11 2 7 10 0 9 2 11 11 2 3 16 11 9 13 14 13 9 1 11 2
13 9 2 0 7 0 9 7 3 0 9 7 9 2
17 10 9 1 1 10 9 13 9 1 10 9 1 12 9 9 3 2
9 15 4 1 9 12 9 7 9 2
22 15 4 0 2 7 3 0 3 1 2 16 10 0 9 4 13 10 0 2 9 2 2
12 9 13 2 16 11 3 1 9 13 0 9 2
13 2 8 4 11 9 1 9 1 11 2 13 15 2
12 15 13 1 14 4 10 9 1 9 7 9 2
48 1 11 9 11 13 10 0 9 1 11 9 2 11 2 2 11 11 11 2 1 9 1 11 9 2 16 11 13 2 16 10 0 0 9 1 10 0 9 1 11 4 13 10 0 9 1 9 2
8 9 13 10 9 1 11 9 2
27 0 1 10 13 9 13 3 10 9 1 9 2 3 15 4 4 13 13 0 9 1 14 13 9 1 9 2
43 15 4 13 1 10 9 1 8 1 2 16 9 2 15 3 4 13 1 9 1 10 0 2 0 9 2 13 9 1 14 13 15 1 15 2 15 4 13 1 10 0 9 2
2 9 13
17 7 3 4 3 13 9 1 10 0 9 2 15 4 13 1 9 2
31 3 13 3 0 9 2 7 13 15 9 2 4 15 13 1 10 0 9 2 11 2 7 0 9 1 1 9 11 7 11 2
14 9 13 3 1 9 7 13 1 12 8 10 0 9 2
44 1 3 10 0 9 1 11 4 4 13 9 9 1 0 9 1 12 2 3 1 10 0 9 11 13 12 9 1 11 2 7 0 10 9 1 11 3 4 3 0 1 10 9 2
18 0 7 0 7 3 3 0 10 0 0 10 2 3 4 0 1 15 2
24 15 13 2 16 11 9 13 1 14 13 11 1 14 13 11 2 3 3 4 4 0 2 3 2
12 15 4 3 3 2 15 3 3 13 10 9 2
11 3 13 10 0 9 1 14 13 0 9 2
6 15 4 10 0 9 2
35 9 9 4 3 3 3 0 2 7 10 0 9 2 2 1 11 4 13 1 2 2 4 1 9 3 3 0 2 1 3 1 12 9 3 2
14 11 11 2 3 4 12 9 2 4 0 1 11 9 2
7 13 3 1 9 7 9 2
7 9 7 9 13 3 9 2
11 13 1 10 9 14 13 0 9 1 9 2
33 15 4 13 0 9 1 11 7 13 10 9 1 10 13 0 9 1 12 2 15 13 15 0 9 1 3 11 7 10 13 0 9 2
15 2 7 1 9 1 9 13 15 9 1 9 1 11 9 2
12 1 0 9 2 1 9 2 13 15 3 9 2
16 3 3 1 9 3 4 13 9 1 0 9 9 1 0 9 2
1 9
10 15 4 3 3 2 15 4 13 3 2
48 9 2 10 9 2 3 10 9 2 15 1 9 7 9 13 14 13 10 9 1 10 9 7 10 9 1 9 2 7 1 13 14 13 10 9 2 13 10 13 9 1 10 0 9 1 10 9 2
10 11 2 3 10 9 1 10 0 9 2
3 0 9 2
14 3 13 15 0 1 9 1 9 7 13 3 1 9 2
7 3 3 15 13 15 3 2
2 5 12
15 7 15 13 15 2 15 13 10 0 9 9 1 9 3 2
18 7 3 4 15 10 3 0 7 0 9 1 0 9 2 15 4 13 2
9 15 13 3 3 10 9 1 15 2
30 1 14 13 10 9 1 9 1 9 1 9 2 15 4 13 3 1 10 9 2 4 9 11 13 9 1 14 13 9 2
15 15 13 9 13 1 9 2 7 16 9 1 3 4 13 2
31 15 4 3 0 2 7 16 3 13 15 2 15 4 13 10 13 9 1 15 2 3 4 15 3 13 3 2 2 13 9 2
23 3 13 10 0 0 2 16 11 11 3 13 10 9 2 10 9 1 10 9 2 11 11 2
12 15 4 13 1 0 9 1 11 11 1 11 2
11 9 13 0 1 3 2 7 11 13 9 2
26 9 9 13 1 9 7 1 9 14 13 12 9 1 10 0 7 0 9 2 1 9 13 1 1 9 2
7 2 3 4 15 0 9 2
24 11 11 2 9 1 9 2 9 2 1 11 1 11 2 4 1 10 9 13 9 1 10 0 2
11 7 3 16 15 13 3 1 10 9 9 2
24 7 1 15 2 15 4 13 12 9 2 7 1 3 13 10 9 1 9 1 10 0 7 0 2
10 3 13 15 15 1 9 1 0 9 2
22 15 4 11 11 2 9 1 9 1 9 1 11 2 15 13 10 0 9 1 11 3 2
15 1 11 13 15 12 9 1 9 2 1 11 3 10 0 2
31 10 0 1 11 9 4 1 9 13 2 16 10 0 9 3 13 2 16 15 3 3 4 13 9 1 2 16 9 13 9 2
24 2 9 9 4 13 15 3 3 10 0 9 2 16 15 3 3 13 10 9 2 2 13 15 2
10 9 4 13 9 1 9 7 9 11 2
30 11 13 2 16 10 0 2 0 9 7 0 9 1 10 0 0 7 0 9 1 9 1 9 4 13 10 9 1 9 2
49 9 13 3 1 0 9 1 9 9 9 1 9 1 11 2 7 9 9 2 11 11 2 3 4 9 1 11 2 4 1 0 9 13 15 15 9 1 9 2 16 11 11 3 13 3 1 0 9 2
2 9 3
31 9 11 4 2 0 2 7 3 13 3 2 16 11 11 7 11 11 1 9 13 2 15 15 4 13 1 0 9 1 9 2
28 11 1 9 13 12 8 2 15 1 9 9 13 0 9 2 10 3 0 9 13 1 10 0 12 8 9 2 2
16 2 15 4 3 13 2 16 15 4 13 10 0 9 1 11 2
13 1 10 9 7 10 9 1 9 13 15 1 9 2
20 1 1 3 0 10 9 13 9 9 1 0 9 7 0 9 14 13 1 9 2
19 1 9 13 12 0 9 1 12 9 9 2 12 9 9 7 12 9 9 2
28 3 4 9 2 9 2 3 3 3 10 0 1 11 11 1 8 1 1 11 2 1 10 9 3 13 1 9 2
12 3 15 1 9 2 7 3 15 1 14 13 2
27 1 10 0 9 9 4 15 3 1 9 13 9 1 10 0 0 9 2 3 1 16 9 13 3 3 13 2
12 11 13 1 8 8 10 9 1 8 1 9 2
33 15 4 3 13 15 13 1 10 9 1 9 2 15 4 3 0 2 7 10 0 9 1 9 2 15 4 4 3 0 7 3 0 2
17 3 3 2 13 9 2 8 11 11 2 9 1 9 1 11 9 2
12 9 13 10 0 9 7 0 9 1 0 9 2
8 15 9 13 1 10 11 9 2
6 16 15 13 1 9 2
13 7 15 4 9 1 2 16 9 3 13 10 9 2
34 3 4 3 3 13 10 9 2 7 3 13 3 10 3 13 9 1 11 9 2 16 15 13 0 9 1 14 13 0 9 3 1 15 2
24 10 0 9 11 13 1 9 2 15 1 10 0 9 1 9 4 13 1 9 1 9 7 9 2
8 7 15 4 15 3 3 13 2
6 15 4 13 1 15 2
2 10 9
18 1 9 4 9 13 1 2 16 15 4 0 14 13 0 9 1 9 2
20 3 4 15 3 13 1 9 1 11 2 9 11 1 11 7 1 11 11 9 2
21 9 13 15 1 0 9 1 0 9 1 11 2 15 13 2 16 9 4 3 0 2
7 3 2 3 13 10 9 2
11 10 0 9 13 3 1 10 0 9 9 2
2 0 9
10 15 4 4 13 0 9 1 9 9 2
14 1 9 4 11 11 0 1 0 9 1 11 11 11 2
26 15 13 15 1 14 13 3 1 2 3 1 9 2 13 15 3 1 9 2 16 14 13 1 0 9 2
56 16 3 13 10 9 1 10 0 9 2 4 3 8 13 10 0 9 2 15 10 9 4 13 1 2 7 3 4 3 13 1 9 9 1 10 0 11 11 2 2 13 11 11 7 13 1 2 16 9 1 11 11 3 4 13 2
14 15 4 10 0 9 1 2 3 15 4 13 10 9 2
12 15 2 15 13 15 15 2 15 13 15 15 2
24 11 11 13 2 16 3 3 13 9 1 14 13 0 9 7 9 1 3 1 12 9 1 9 2
10 1 10 0 7 0 7 0 0 9 2
15 3 13 15 9 1 14 13 3 3 2 3 15 13 13 2
12 3 13 3 3 9 1 14 13 10 0 9 2
12 9 2 9 2 9 7 9 4 13 1 9 2
19 3 0 1 10 0 9 3 13 10 0 0 9 1 9 9 1 0 9 2
7 15 13 10 9 1 9 2
37 11 9 4 10 9 2 15 13 9 2 1 11 3 4 13 3 1 2 15 9 1 3 4 13 3 1 2 7 15 2 15 1 11 9 4 13 2
7 0 4 13 3 1 9 2
6 8 5 8 9 5 8
18 15 4 3 4 4 0 1 15 14 13 3 1 10 9 1 0 9 2
30 3 11 11 7 9 11 11 1 11 9 13 2 16 9 4 13 10 9 2 16 15 4 13 9 1 10 3 0 9 2
18 7 3 13 15 0 9 1 9 2 9 1 9 7 0 9 1 9 2
9 2 11 13 15 3 1 10 9 2
4 6 7 6 2
10 3 4 15 13 15 3 3 1 9 2
29 11 11 2 9 2 4 3 1 9 11 11 1 0 9 1 11 13 9 1 10 9 1 9 1 11 11 1 11 2
12 3 4 15 3 13 15 2 2 13 11 11 2
2 12 2
32 1 3 0 2 3 3 2 9 7 9 4 9 7 9 3 13 15 0 3 2 16 15 3 13 10 3 0 9 1 11 11 2
13 15 4 3 4 13 3 3 3 1 9 1 15 2
26 3 1 9 4 15 13 10 0 9 7 10 9 13 1 9 2 16 15 4 13 9 1 9 1 11 2
6 11 11 11 2 0 2
41 3 4 3 9 16 9 4 13 11 2 7 16 15 1 9 13 15 2 15 3 13 2 11 2 2 10 3 0 9 1 10 0 9 10 7 10 9 3 1 11 2
27 15 13 3 9 7 4 1 12 10 0 9 3 13 9 1 10 1 10 0 9 7 9 1 10 0 9 2
15 1 9 13 15 1 11 3 1 12 10 0 9 1 9 2
18 15 4 13 10 9 2 15 13 10 0 9 1 9 2 3 1 9 2
14 15 4 3 13 3 1 2 15 15 4 13 15 1 2
25 9 11 11 13 12 9 1 9 1 10 0 9 2 16 11 13 9 2 16 3 4 13 0 9 2
29 10 0 9 1 10 3 13 9 9 1 9 4 3 13 11 1 14 13 2 16 3 4 13 3 1 10 0 9 2
37 15 4 10 9 2 15 4 13 3 2 7 2 1 15 4 13 1 9 2 3 4 15 13 9 1 9 10 9 2 15 13 9 1 9 1 9 2
18 9 4 13 3 1 0 9 2 3 1 9 2 15 3 4 13 3 2
24 7 1 10 13 9 13 15 1 2 16 15 3 4 13 1 15 14 13 15 1 9 1 9 2
19 9 13 9 1 14 13 1 9 2 7 9 4 3 4 13 9 1 9 2
10 2 15 13 0 9 9 3 1 9 2
2 0 9
12 9 2 11 2 9 2 9 7 9 4 9 2
18 1 9 4 1 9 0 9 2 9 7 9 1 9 9 7 2 9 2
6 2 6 2 3 3 2
27 2 15 4 13 1 0 7 4 15 3 2 3 3 11 7 11 13 1 9 1 9 2 2 13 11 11 2
25 11 9 4 13 14 13 10 9 1 11 1 11 1 11 2 16 10 0 9 1 11 13 1 11 2
9 2 15 13 9 10 9 1 9 2
16 15 13 2 16 3 13 1 10 0 7 12 9 9 1 9 2
6 9 1 10 0 11 2
5 3 14 13 3 2
3 9 7 9
23 11 2 3 0 9 9 4 13 9 2 4 1 9 1 9 13 1 0 9 2 13 9 2
21 1 10 0 7 0 9 1 9 13 9 11 11 0 9 1 2 16 9 4 13 2
14 7 15 13 3 3 2 3 1 15 13 9 1 9 2
1 9
13 2 3 4 15 0 7 0 1 14 13 10 9 2
9 9 4 13 14 13 9 1 15 2
11 1 9 1 9 2 9 2 9 7 9 2
9 9 4 0 1 14 13 15 2 2
40 1 10 9 4 15 0 14 13 1 2 16 10 13 2 0 11 9 9 9 2 9 7 0 9 1 9 9 3 3 13 3 1 10 0 9 9 1 0 9 2
3 13 1 11
10 2 10 0 13 14 4 13 8 9 2
21 9 2 9 1 7 13 1 9 1 9 1 9 1 9 7 9 1 9 1 9 2
16 15 13 10 0 1 14 4 10 9 7 9 1 10 0 9 2
11 2 15 13 3 11 2 2 13 11 11 2
25 3 7 3 13 10 0 9 3 2 3 0 2 2 15 0 9 2 13 15 1 10 0 9 2 2
32 15 4 13 1 9 1 9 2 16 3 13 9 1 9 2 13 11 11 2 15 1 9 13 3 1 9 0 9 11 1 11 2
10 7 3 4 15 3 11 9 1 9 2
17 11 11 13 10 0 2 10 13 2 0 2 7 13 15 0 9 2
6 15 4 13 0 9 2
22 15 13 7 13 9 3 3 1 9 2 10 0 9 1 10 0 9 1 9 7 9 2
12 2 15 13 11 1 10 3 0 7 0 9 2
25 2 15 4 3 13 15 7 13 2 16 10 0 9 3 4 10 0 9 2 2 13 9 11 11 2
5 9 2 0 9 12
15 16 15 13 14 13 0 9 2 4 15 13 9 15 9 2
2 6 2
6 3 4 3 13 15 2
8 3 13 0 9 3 1 9 2
21 4 15 3 3 4 10 9 2 9 2 16 15 4 0 3 7 16 15 13 9 2
21 3 4 15 3 10 0 9 1 10 9 2 0 4 13 3 1 1 9 0 9 2
11 13 9 2 9 7 9 2 9 12 2 2
15 1 9 2 1 9 2 1 9 2 1 9 2 1 9 2
31 12 13 1 10 9 1 9 2 7 10 0 13 15 0 3 3 1 3 2 13 0 9 11 11 1 10 0 9 1 9 2
1 9
8 2 3 1 9 2 15 13 2
16 10 9 13 15 3 3 1 14 13 2 16 15 13 3 13 2
11 11 13 0 0 0 9 2 3 11 9 2
27 16 15 3 4 13 10 9 9 2 4 15 0 2 7 14 4 13 3 1 9 1 15 4 3 3 9 2
3 9 13 15
11 10 12 9 4 3 13 1 10 10 9 2
12 9 4 13 10 9 1 12 9 1 9 0 2
3 2 11 2
3 9 1 11
33 9 1 9 4 11 3 3 0 9 1 9 2 7 15 4 0 9 2 16 9 13 0 9 1 0 9 1 9 1 10 0 9 2
10 10 0 1 11 12 9 4 3 0 2
15 16 9 4 0 13 9 3 12 9 1 9 2 9 9 2
48 3 4 15 3 10 0 1 11 2 15 13 9 2 7 4 15 3 13 1 10 0 9 2 8 2 11 7 11 2 6 3 4 15 3 3 13 10 9 2 16 15 4 10 0 2 0 9 2
14 15 13 3 2 16 15 3 13 10 0 9 1 9 2
40 1 9 13 11 11 3 10 9 1 10 0 9 2 1 11 7 9 2 7 0 9 1 10 9 9 2 1 10 0 9 1 9 2 3 0 1 9 9 3 2
6 10 0 9 1 11 2
20 11 2 3 4 4 10 0 9 2 13 3 3 3 0 14 13 1 11 1 2
73 11 0 9 13 1 9 1 9 1 10 0 9 1 9 2 7 15 13 2 16 3 13 3 3 0 1 11 11 2 7 3 3 4 15 3 13 15 3 2 16 10 9 3 4 13 3 3 3 1 15 1 9 11 2 7 3 3 4 13 1 11 11 8 14 13 1 9 2 3 3 13 15 2
23 1 10 0 0 9 13 15 15 2 16 9 1 9 12 4 0 1 0 9 1 1 0 2
20 2 15 13 10 3 0 9 1 9 1 9 1 9 2 9 2 9 7 9 2
21 0 9 4 3 3 0 7 0 1 9 9 2 3 4 3 0 7 13 9 3 2
15 1 12 13 15 1 14 4 13 10 0 9 1 13 9 2
20 1 9 9 13 10 0 0 9 3 1 11 7 4 13 7 13 3 1 9 2
32 1 12 13 15 10 9 1 10 8 9 2 7 16 10 0 9 1 11 3 1 9 4 13 1 10 9 2 13 9 13 0 2
17 9 13 3 14 13 2 16 15 1 10 9 15 4 13 10 9 2
2 0 2
17 15 4 1 13 9 13 2 16 15 4 13 9 1 9 3 2 2
27 9 4 13 1 10 0 9 1 10 0 9 1 10 9 9 1 0 9 2 9 7 9 1 9 1 11 2
4 3 13 9 2
7 2 3 13 15 1 15 2
3 9 1 11
9 10 0 9 4 13 1 0 9 2
4 0 9 1 9
41 2 15 13 3 15 14 13 1 2 16 11 4 13 15 1 10 0 0 9 1 10 13 9 7 13 2 16 10 10 9 3 3 4 13 10 9 2 2 13 15 2
12 0 7 3 3 0 9 15 4 13 1 11 2
20 7 1 11 2 6 2 3 13 3 9 1 10 13 9 1 10 12 0 9 2
12 9 13 0 9 1 9 1 14 13 15 1 2
26 7 15 12 4 0 1 2 16 10 9 3 3 1 0 9 4 13 1 14 13 9 7 9 0 9 2
27 10 9 1 10 0 7 0 9 4 3 3 3 0 1 9 2 2 11 11 11 11 11 11 2 13 15 2
3 9 9 12
40 9 1 9 9 2 11 11 2 11 2 2 4 13 2 16 10 0 0 9 1 11 4 4 13 1 11 2 7 15 4 10 9 2 9 11 11 2 3 13 2
21 9 11 1 9 11 1 11 4 0 9 1 10 0 9 9 9 2 3 12 13 2
18 15 13 10 0 13 1 10 9 1 9 2 3 13 15 3 1 15 2
43 10 0 11 2 3 4 15 1 10 3 0 9 2 15 4 13 2 13 3 3 10 0 9 1 9 3 3 1 14 13 9 1 2 16 10 9 1 9 3 3 4 13 2
37 11 13 2 16 15 0 9 1 9 13 10 9 1 10 9 2 11 11 2 7 10 0 9 1 14 13 9 1 12 8 2 12 9 2 1 9 2
23 1 0 9 13 9 2 7 11 9 13 9 9 2 16 11 11 13 1 14 13 1 9 2
17 2 15 4 4 0 14 13 9 2 16 15 3 4 13 1 9 2
25 9 2 10 9 7 10 9 2 15 13 1 7 13 10 9 7 10 9 1 9 2 7 1 13 2
15 3 4 13 10 0 9 15 13 2 3 2 6 1 15 2
2 11 11
4 15 4 0 2
12 3 1 9 13 15 10 9 1 14 4 3 2
15 1 9 1 9 11 11 13 15 9 2 16 15 4 9 2
13 15 4 13 10 9 3 1 10 0 0 9 9 2
10 3 4 11 13 9 13 15 1 9 2
18 2 15 13 10 0 9 1 11 9 2 2 13 9 11 11 2 9 2
12 9 1 9 7 11 1 2 10 0 9 2 2
13 9 13 3 13 1 2 15 3 13 3 1 9 2
33 2 11 13 1 9 2 13 9 3 7 13 3 9 13 1 10 9 1 9 2 3 10 0 9 4 13 3 1 9 1 0 9 2
19 15 13 15 3 3 2 7 16 3 4 13 10 0 9 2 4 0 13 2
18 15 4 13 15 13 1 8 8 11 11 2 1 11 8 8 11 11 2
13 1 9 12 1 0 9 13 10 9 1 10 9 2
9 3 13 10 9 1 0 9 9 2
10 3 4 1 12 13 12 9 1 9 2
15 16 9 1 9 13 3 2 13 3 9 1 10 0 9 2
21 0 0 9 7 9 4 13 1 10 9 1 9 1 10 0 2 0 0 9 2 2
46 4 15 4 0 1 2 16 10 9 7 9 2 15 4 13 1 14 13 10 3 0 9 1 9 3 9 1 9 3 3 13 15 1 15 2 7 3 13 14 13 9 1 10 0 9 2
36 1 10 9 15 13 3 3 0 0 0 9 7 13 15 1 15 1 9 2 16 10 0 9 13 0 9 1 14 13 1 0 9 1 10 9 2
8 7 11 13 3 10 0 9 2
30 15 13 3 1 11 9 9 7 9 2 15 13 2 16 15 13 15 1 0 2 16 10 0 9 4 13 9 1 15 2
18 0 9 4 15 13 1 9 1 9 11 11 9 1 11 11 1 11 2
23 9 13 3 1 10 0 2 3 0 9 1 10 9 1 11 0 9 2 3 15 13 9 2
14 2 15 13 3 2 16 10 0 9 4 10 0 9 2
36 15 13 10 13 11 11 2 2 13 15 3 2 0 1 9 15 2 1 9 12 2 0 2 1 9 12 2 0 2 1 9 12 2 0 2 2
19 15 4 3 13 10 0 9 1 2 3 15 4 13 9 2 15 15 13 2
18 10 0 9 4 10 13 0 9 2 3 3 4 3 0 1 10 9 2
9 15 13 0 2 16 15 4 0 2
19 2 11 2 13 15 1 9 11 2 7 9 1 9 4 13 13 10 9 2
10 15 13 3 2 16 15 4 3 0 2
24 1 10 0 0 9 13 9 3 1 8 8 1 9 13 3 9 1 0 9 1 11 7 11 2
7 10 0 9 1 0 9 2
19 9 2 15 4 13 2 7 1 10 0 9 3 13 14 13 10 13 9 2
38 2 6 2 15 13 3 0 2 7 3 4 15 3 13 15 9 1 9 2 0 2 2 15 13 3 14 13 1 14 13 2 14 2 4 13 2 2 2
7 3 13 10 9 1 9 2
37 10 12 9 2 2 2 8 8 2 9 13 1 9 5 8 2 11 2 9 9 2 8 2 9 9 2 11 2 9 9 5 8 3 5 0 0 2
44 10 9 1 11 2 3 3 1 3 11 4 15 1 11 3 0 9 1 13 2 13 16 9 4 0 7 0 2 7 4 13 1 3 0 1 9 7 9 1 0 7 0 9 2
19 15 13 1 9 9 1 9 7 13 10 0 9 1 3 15 7 10 9 2
33 9 13 3 3 1 0 10 0 9 1 14 13 9 7 9 0 7 14 13 1 8 7 9 1 0 9 2 7 3 3 13 15 2
2 12 2
6 15 4 11 13 3 1
12 1 9 1 2 11 2 13 10 9 1 9 2
13 15 13 3 2 3 0 0 9 9 4 13 1 2
28 12 9 13 2 15 15 13 2 7 1 13 1 11 7 11 13 15 3 2 15 3 4 13 9 3 1 9 2
20 10 0 9 13 13 9 1 9 1 9 2 3 1 9 1 14 13 0 9 2
10 9 13 2 16 10 9 4 4 13 2
30 15 13 1 9 13 2 16 2 9 9 1 9 2 2 15 4 3 13 1 9 2 4 4 10 0 9 1 9 9 2
54 2 0 9 1 9 2 2 1 10 9 4 13 2 2 2 4 0 9 2 1 9 1 11 11 9 13 2 10 0 0 7 0 9 2 15 4 13 12 2 13 3 14 13 9 9 1 12 1 3 11 1 11 2 2
13 3 13 3 1 0 7 0 9 1 9 1 11 2
41 9 13 1 15 2 15 4 3 13 1 9 1 12 2 7 1 10 0 9 1 13 9 1 9 1 9 3 1 9 2 4 9 3 13 3 1 10 0 9 9 2
12 15 1 9 9 9 11 11 13 1 13 9 2
4 15 4 0 2
36 1 0 9 13 0 12 9 13 15 11 11 11 1 11 1 0 12 1 9 7 13 3 10 0 9 2 15 13 1 9 1 10 0 11 11 2
23 2 1 0 9 2 3 0 2 1 0 1 0 9 9 2 3 16 15 13 1 12 9 2
11 7 4 15 3 9 1 14 13 2 13 2
23 3 2 3 1 9 7 1 9 2 13 9 1 2 10 0 9 1 9 1 0 9 2 2
13 7 15 4 3 3 13 3 2 1 9 2 13 2
2 11 13
8 3 4 15 3 3 0 3 2
9 15 13 1 10 10 9 1 8 2
55 15 4 1 10 12 9 3 1 12 9 2 7 15 9 13 15 1 9 7 13 3 1 9 1 14 13 10 0 9 3 2 13 9 7 4 3 1 14 13 3 7 13 3 10 0 9 7 0 1 9 13 7 13 9 2
14 15 4 3 3 3 13 2 16 15 1 0 13 3 2
3 9 0 9
16 10 0 9 13 0 9 2 16 15 13 9 7 9 1 9 2
3 11 2 11
7 15 13 9 3 1 15 2
9 3 13 11 10 9 1 10 9 2
14 10 12 0 0 9 13 3 1 10 9 7 13 11 2
18 15 13 3 3 1 2 16 3 3 13 10 0 9 1 10 0 9 2
21 10 9 9 3 4 10 3 0 9 2 10 0 9 11 11 11 2 4 13 13 2
47 3 4 15 0 14 2 13 2 10 0 9 1 11 2 7 13 15 0 1 9 1 10 0 9 2 3 9 7 10 0 9 2 11 2 2 2 13 11 11 11 2 9 1 11 7 11 2
11 2 15 13 10 3 0 9 2 13 11 2
26 11 13 15 7 13 1 9 2 2 6 2 15 13 3 2 13 2 11 2 6 2 15 13 3 2 2
9 15 4 15 2 15 3 13 15 2
14 10 9 1 9 1 11 11 7 9 4 3 13 9 2
32 7 1 11 11 1 10 0 9 2 9 9 2 4 15 9 1 14 13 1 9 3 1 9 2 3 4 4 0 1 11 11 2
31 1 12 4 11 11 13 1 9 1 10 0 9 2 7 15 4 10 9 2 15 3 13 1 9 1 10 0 9 1 11 2
6 1 9 1 11 9 2
9 11 13 15 1 14 13 1 3 2
23 7 15 4 3 15 1 9 1 9 2 13 9 11 11 2 15 13 9 12 9 1 9 2
23 2 15 13 3 3 13 15 3 2 13 3 7 13 3 2 15 13 15 0 10 0 9 2
26 9 4 3 13 3 1 9 1 9 1 14 13 15 3 1 9 7 3 13 3 2 16 9 4 3 2
18 11 13 9 3 7 3 1 9 2 16 15 13 3 1 10 0 9 2
9 15 4 13 1 0 9 1 9 2
13 4 9 10 0 9 1 9 1 2 7 15 0 2
20 9 1 9 13 3 9 1 14 13 3 1 9 2 16 9 4 13 1 8 2
18 15 13 0 9 1 10 9 1 11 1 12 2 7 4 3 13 3 2
11 15 4 0 1 15 2 7 3 1 15 2
10 11 11 4 13 7 13 12 9 3 2
11 8 4 0 1 14 13 15 1 10 9 2
11 15 4 3 3 1 10 0 9 1 9 2
32 10 0 0 9 4 13 15 2 7 11 7 15 1 10 12 9 2 15 3 13 3 2 13 2 16 15 4 13 15 1 15 2
12 2 6 2 13 15 1 10 0 7 13 9 2
15 16 15 13 15 3 1 9 2 13 1 10 9 3 3 2
5 13 12 9 3 2
8 9 4 13 2 3 7 3 2
3 3 5 12
18 13 3 10 9 2 15 4 13 15 9 2 15 13 9 1 9 9 2
17 2 6 2 3 4 15 3 13 1 0 9 2 2 13 11 11 2
46 9 13 2 16 15 1 14 4 13 1 15 1 10 9 1 9 7 9 2 3 4 13 1 10 9 3 1 15 14 13 9 7 9 2 16 9 1 9 7 9 3 3 4 13 3 2
12 3 13 9 10 0 9 1 0 9 1 9 2
16 10 0 9 13 1 9 1 11 11 1 9 1 11 7 11 2
15 13 9 1 9 1 9 7 13 1 9 2 15 3 13 2
9 1 0 9 4 15 13 3 3 2
25 5 9 1 14 13 10 0 9 2 15 3 13 15 13 1 9 2 4 3 10 13 9 1 9 2
3 9 1 9
17 15 4 3 3 4 10 9 2 16 9 4 13 3 1 9 9 2
16 3 4 3 13 1 12 1 9 2 3 11 3 4 4 9 2
18 10 0 9 4 1 12 2 3 10 0 9 13 12 9 1 10 9 2
12 15 4 12 0 1 1 9 1 9 1 12 2
36 9 1 10 12 9 4 3 7 0 9 1 9 2 7 3 4 9 3 0 8 9 2 7 3 4 15 0 2 16 15 3 13 10 12 9 2
26 1 10 0 9 2 9 1 10 0 12 9 1 12 2 4 9 3 1 0 9 13 1 12 9 9 2
36 15 4 15 1 10 9 2 10 0 9 13 3 3 1 1 2 11 2 2 3 3 3 3 4 10 0 7 10 15 2 8 3 7 0 3 2
40 9 1 12 4 13 1 9 1 11 11 2 8 8 8 8 8 8 2 11 8 8 8 8 8 11 11 8 11 2 2 11 11 12 2 12 2 8 2 12 2
22 15 13 11 1 15 1 2 9 2 2 7 15 13 3 12 9 3 1 9 3 3 2
29 15 13 1 12 9 2 3 12 9 2 0 1 9 2 0 0 9 2 0 9 2 0 0 9 7 3 1 9 2
14 11 11 13 1 10 9 13 10 9 1 9 1 9 2
12 10 9 4 13 1 0 11 9 11 11 9 2
11 9 4 10 0 9 1 0 9 1 11 2
15 3 1 15 13 3 1 10 0 13 15 1 15 1 3 2
54 9 1 11 2 10 9 9 2 15 4 8 0 9 11 11 7 15 9 0 7 0 9 2 16 15 13 1 9 1 9 7 9 2 4 3 13 1 9 9 7 4 8 13 2 15 10 0 9 1 9 4 13 3 2
22 15 4 13 14 13 1 15 1 15 2 7 15 13 3 2 16 9 3 3 13 15 2
25 9 4 10 9 1 15 1 9 3 0 9 2 15 13 10 0 9 1 0 9 1 11 9 1 9
20 3 4 13 12 9 2 7 0 9 13 2 16 15 10 9 13 3 0 0 2
33 2 10 0 9 4 1 9 13 14 13 11 2 7 3 4 9 11 11 13 10 0 0 9 2 16 10 9 3 4 13 9 3 2
26 1 12 8 1 11 13 11 3 1 12 8 2 10 9 2 15 13 1 10 9 1 3 12 1 9 2
4 13 15 15 2
9 9 7 9 2 8 2 12 9 2
41 7 15 4 10 9 2 16 0 0 9 13 1 14 13 10 13 9 2 3 1 0 9 3 1 9 4 4 3 3 0 14 13 7 13 7 3 3 0 14 13 2
31 7 11 4 3 9 1 11 2 15 1 10 9 2 15 13 3 3 1 8 8 2 15 3 4 13 10 9 1 0 9 2
24 2 15 13 3 3 13 12 9 9 2 7 13 7 13 8 7 9 1 9 1 14 13 3 2
12 14 13 1 11 4 3 10 9 1 11 11 2
14 2 10 0 9 1 12 4 3 0 1 10 0 9 2
11 3 10 9 4 11 11 7 11 11 3 2
7 10 0 9 1 10 9 2
10 9 4 4 0 7 0 14 13 0 2
12 7 15 13 0 9 1 9 1 10 13 9 2
35 3 13 9 9 1 10 12 9 0 9 2 7 10 0 11 13 1 14 13 1 0 10 1 9 2 15 1 0 9 4 13 9 1 9 2
15 15 13 14 13 1 9 7 4 13 1 14 13 1 9 2
65 1 9 1 9 13 15 3 2 16 3 3 4 13 9 1 10 9 1 9 2 16 10 0 9 13 1 9 1 9 2 7 16 3 3 4 13 9 1 10 11 2 8 8 8 2 2 3 16 10 0 9 3 3 4 13 10 9 1 9 2 1 15 13 1 2
11 2 16 15 13 2 13 11 10 3 0 2
3 0 7 0
2 9 2
16 7 15 4 3 13 1 11 2 16 0 10 9 13 1 11 2
5 3 13 0 9 2
17 7 9 1 9 7 9 13 9 3 1 10 9 2 1 10 9 2
44 11 11 2 9 2 4 13 2 9 1 9 2 2 10 0 9 2 11 9 13 15 9 2 16 9 1 10 0 9 1 9 4 13 15 1 10 0 1 14 13 15 3 3 2
17 10 0 9 4 3 13 1 10 13 9 1 9 1 14 13 9 2
39 1 9 4 15 9 1 11 7 11 9 2 9 1 9 1 11 9 2 8 2 9 2 11 7 9 9 8 2 11 9 2 0 9 2 9 7 0 9 2
2 12 9
15 13 9 4 3 13 3 1 9 1 14 4 13 10 9 2
17 10 9 4 13 13 9 2 3 3 9 7 15 3 13 1 11 2
3 9 4 13
18 2 1 9 1 9 12 4 0 3 13 9 1 15 14 13 10 9 2
44 7 9 11 11 4 3 10 9 13 2 16 15 13 3 7 13 2 9 12 2 2 15 1 10 9 4 4 13 10 0 9 1 9 1 14 4 13 3 1 10 9 1 9 2
12 3 4 15 13 1 10 9 8 1 9 2 2
2 9 2
7 13 15 13 3 10 9 2
23 7 3 16 15 4 13 12 9 9 1 14 13 12 9 1 10 9 1 10 9 1 11 2
10 9 4 13 1 11 11 9 2 11 2
30 3 1 11 4 15 4 0 1 13 9 2 7 15 13 14 4 3 1 9 1 9 2 9 7 9 2 2 13 9 2
54 3 13 15 14 13 15 1 9 1 15 1 9 1 9 2 2 1 9 9 13 3 1 2 16 10 9 1 9 1 9 4 13 10 9 1 9 2 7 10 9 4 13 1 2 1 15 9 10 0 9 13 0 9 2
20 2 15 4 3 3 0 2 15 3 13 2 16 10 9 13 1 10 0 9 2
9 9 4 1 10 0 13 3 3 2
21 15 13 2 16 15 3 4 13 3 1 10 9 0 9 2 14 13 7 13 15 2
36 1 9 4 10 9 13 1 10 0 9 7 13 3 0 9 1 11 2 1 3 12 9 1 11 2 1 15 10 9 3 13 9 1 2 9 2
43 9 1 10 0 8 9 2 11 2 9 13 1 0 0 9 9 1 10 9 1 9 2 15 9 1 9 4 13 1 12 7 3 12 4 9 2 16 3 13 9 1 12 2
19 11 7 11 4 10 0 1 13 9 1 11 2 15 13 1 9 1 12 2
20 2 15 13 3 3 0 3 1 3 10 0 9 1 9 1 10 0 9 2 2
16 10 0 9 13 1 9 2 7 10 0 13 3 1 1 9 2
18 15 13 2 16 11 4 13 3 0 1 9 1 14 13 15 1 9 2
10 2 9 1 11 4 13 3 12 9 2
42 9 1 11 11 0 9 1 9 13 3 2 16 15 1 0 9 3 13 1 14 13 1 9 1 10 9 3 2 16 15 3 13 15 0 1 3 14 13 9 1 9 2
19 10 0 1 10 13 9 4 10 0 9 2 11 2 1 9 11 1 11 2
12 3 4 13 15 2 13 10 9 1 11 11 2
5 15 4 3 0 2
23 15 13 2 16 15 13 3 13 1 7 3 0 1 10 9 2 15 13 1 10 0 9 2
5 3 3 11 11 2
8 3 13 3 3 10 13 9 2
21 15 4 10 9 2 10 0 9 2 2 11 11 11 11 11 11 11 2 2 13 2
6 15 13 3 9 3 2
1 9
22 15 2 15 4 13 14 13 10 9 1 9 1 0 10 9 1 10 9 2 13 9 2
8 3 13 12 9 9 1 9 2
18 16 10 0 9 13 12 9 3 2 13 9 2 15 4 13 0 9 2
20 12 9 3 4 9 0 9 0 1 13 2 7 3 13 9 1 10 0 9 2
20 9 1 0 7 0 9 9 2 15 13 1 9 2 4 13 13 3 1 9 2
17 11 11 7 11 11 11 4 4 0 1 10 0 1 9 1 9 2
11 1 10 0 9 1 11 13 11 12 9 2
8 3 13 9 15 3 1 9 2
22 3 4 13 9 1 10 9 1 9 2 16 15 13 9 1 14 13 10 9 1 9 2
5 11 13 1 9 2
19 12 9 9 1 9 4 11 13 3 1 10 9 13 1 10 0 0 9 2
6 15 13 3 1 9 2
22 15 13 3 1 9 1 14 13 1 9 1 9 1 10 9 2 3 2 3 2 3 2
17 7 16 15 3 13 14 13 9 1 15 2 13 15 9 1 15 2
6 8 5 8 9 5 8
6 9 13 3 1 9 2
20 15 4 9 1 10 9 2 15 9 4 13 1 9 1 9 1 8 7 9 2
26 3 1 9 3 3 4 13 9 2 7 3 15 3 13 3 3 2 4 9 9 10 0 9 1 9 2
23 2 1 10 9 9 3 13 10 0 1 9 2 16 15 13 10 9 2 3 4 4 0 2
52 15 13 9 7 13 15 1 10 9 3 1 0 12 9 2 3 15 13 9 1 14 13 12 9 7 10 0 9 13 15 1 10 9 2 15 13 1 9 7 9 2 1 9 2 9 2 1 9 7 1 9 2
3 9 13 2
14 9 1 9 1 9 4 1 0 9 13 9 1 11 2
20 2 7 9 4 0 2 16 9 4 13 9 9 3 1 9 2 2 13 15 2
6 2 15 13 15 3 2
30 7 16 15 3 13 3 1 9 1 9 7 9 2 4 15 13 10 0 9 1 14 13 9 1 9 1 14 13 9 2
49 10 12 9 4 1 9 9 13 10 9 9 15 1 15 2 7 1 9 9 4 3 13 10 9 2 15 3 4 13 7 3 4 13 1 0 9 1 10 9 0 9 3 1 11 7 3 1 11 2
43 7 12 9 3 13 10 9 1 11 1 10 0 9 14 13 10 0 9 2 15 4 0 14 13 10 9 1 10 0 9 2 10 13 9 11 11 2 1 10 2 9 2 2
15 7 11 4 3 9 1 0 9 2 7 4 4 10 9 2
48 9 4 2 1 15 4 4 11 11 0 2 1 0 9 13 1 8 7 9 2 7 9 4 3 13 1 9 2 15 13 2 15 9 3 4 0 1 9 1 10 9 2 15 13 1 10 9 2
11 15 4 3 3 0 14 13 6 3 2 2
17 15 4 3 4 9 1 9 2 2 13 9 1 11 2 11 11 2
1 9
15 13 9 3 1 10 0 9 2 3 12 9 8 12 9 2
9 3 4 9 2 11 11 2 13 2
10 15 4 0 7 4 13 1 0 9 2
15 3 3 4 15 0 14 13 0 9 1 9 2 13 15 2
13 1 11 13 10 0 9 9 1 12 9 1 9 2
21 9 1 9 1 9 1 10 0 9 7 9 2 13 0 9 12 1 11 11 3 2
9 10 0 9 2 15 13 1 9 2
12 2 3 2 2 13 15 2 2 4 15 4 2
40 9 2 15 13 10 12 9 1 9 1 0 9 12 7 10 9 3 2 13 3 2 15 11 11 2 11 2 1 9 1 11 9 9 4 13 9 1 14 13 2
17 15 13 15 3 2 13 9 1 9 7 13 9 1 10 0 9 2
24 9 1 10 0 9 9 13 2 16 15 4 4 13 1 0 9 7 1 15 13 9 1 9 2
9 1 11 13 15 10 9 2 11 2
22 15 13 15 1 10 9 14 13 9 1 0 9 1 0 9 13 1 9 7 13 9 2
25 15 13 3 2 16 9 1 9 7 9 3 4 13 10 13 9 2 16 9 1 11 13 1 9 2
14 7 3 4 15 13 9 2 3 9 3 13 1 9 2
29 3 4 0 9 2 3 12 9 1 10 0 9 2 7 3 9 13 16 15 1 0 9 13 10 0 9 1 15 2
34 15 4 13 1 10 9 1 11 11 11 1 9 1 2 11 11 2 15 1 10 0 9 1 0 9 2 7 3 4 9 3 3 13 2
6 12 0 9 4 13 2
7 3 4 10 9 15 4 3
26 15 13 3 2 15 4 4 13 10 9 2 16 16 15 4 0 7 0 2 4 15 13 13 10 9 2
32 15 4 3 13 9 1 9 7 4 1 12 9 13 3 1 12 1 9 2 4 13 9 3 0 9 1 9 1 10 10 9 2
4 9 1 9 9
20 0 9 13 15 1 12 9 3 3 1 9 11 11 11 2 7 9 4 13 2
18 10 0 13 9 7 9 1 0 13 2 15 3 13 1 11 0 9 2
57 7 10 0 9 2 15 13 3 1 0 7 0 9 2 7 10 9 2 15 3 4 13 10 9 2 1 4 3 0 2 13 9 3 1 9 7 13 15 1 9 10 0 9 13 1 0 9 9 2 9 2 9 7 13 9 9 2
31 9 4 3 3 3 0 9 2 7 16 9 4 13 13 15 3 3 1 10 9 2 16 10 1 10 0 9 4 13 3 2
8 9 4 0 1 0 0 9 2
18 9 3 13 15 15 2 16 15 4 13 9 13 3 1 10 0 9 2
22 15 13 1 9 11 1 10 13 9 7 10 9 11 2 15 4 13 1 0 1 15 2
7 1 15 4 15 13 9 2
5 13 10 12 9 2
5 2 0 2 9 2
37 2 15 4 13 1 0 9 1 9 2 7 15 4 13 2 16 9 13 9 1 11 9 2 2 13 9 11 11 2 3 3 4 9 1 11 11 2
8 7 3 4 3 13 0 9 2
21 10 0 9 1 9 1 10 0 9 2 10 3 0 9 2 4 3 9 1 9 2
11 7 3 3 15 9 13 2 15 4 13 2
35 9 0 9 4 15 3 3 2 13 3 1 2 2 16 9 2 15 13 15 1 9 7 1 10 9 2 13 0 9 1 10 9 9 3 2
3 0 14 13
19 3 13 3 15 1 10 9 2 15 13 2 15 13 9 1 10 0 9 2
12 1 9 13 10 0 9 1 10 0 9 11 2
9 11 11 4 0 9 7 11 9 2
30 11 11 11 13 2 16 9 2 4 13 1 9 2 7 10 0 9 4 13 2 16 15 4 13 3 1 3 3 2 2
21 15 13 10 9 8 1 10 9 1 9 2 16 15 1 0 9 13 9 1 9 2
9 2 6 2 15 4 15 3 13 2
15 8 4 8 3 13 0 3 7 1 12 13 3 12 0 8
80 11 9 12 9 12 8 12 9 12 9 12 9 12 9 12 9 12 9 12 8 12 9 12 9 11 9 12 9 12 9 12 8 12 9 12 9 12 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 8 8 2 12 9 12 2 9 2 9 2 8 8 2 9 2 9 2 9 2 12 9 12 8 12 9 12 9
3 0 9 2
18 15 4 3 3 0 1 9 2 7 3 13 3 3 0 0 9 2 2
14 0 9 4 3 3 13 2 3 1 15 8 7 9 2
5 15 13 3 3 2
16 11 11 2 15 10 0 9 13 9 1 14 13 2 4 0 2
27 9 1 9 1 2 11 11 2 7 2 0 9 2 4 1 0 3 9 1 9 0 9 2 11 11 2 2
15 15 4 13 1 7 1 9 2 7 15 4 13 1 15 2
1 9
27 10 0 0 9 1 3 3 12 9 13 1 14 13 3 12 9 13 1 12 9 2 3 3 12 9 9 2
3 13 12 9
25 9 13 0 9 1 9 7 13 3 10 9 1 12 9 1 9 1 9 7 13 15 13 1 9 2
2 1 9
33 9 4 13 1 9 9 1 0 9 2 7 11 11 13 1 7 13 14 13 10 9 1 12 9 1 11 3 1 9 9 1 12 2
9 11 11 13 0 1 10 13 11 2
34 9 9 13 14 13 9 1 0 9 1 10 11 9 13 9 2 3 1 9 2 15 1 0 9 4 2 13 2 1 14 8 3 3 2
20 15 13 1 15 3 7 13 15 2 1 15 1 10 0 9 13 3 1 9 2
18 15 4 0 2 15 3 3 4 4 13 9 3 14 13 1 0 9 2
7 2 9 2 11 11 2 2
20 5 1 9 13 15 14 13 3 1 9 2 15 4 13 9 1 14 13 3 2
9 11 13 1 10 0 10 0 9 2
19 9 4 13 1 14 13 10 9 1 10 9 0 2 9 2 1 10 9 2
25 16 15 4 12 9 1 15 4 12 13 15 3 1 0 9 3 1 12 9 2 10 9 7 9 2
23 10 9 13 9 7 9 2 16 3 13 9 1 2 16 9 4 3 13 1 14 13 9 2
4 0 9 1 9
34 13 2 16 13 10 9 9 12 9 2 7 15 13 3 1 9 2 13 15 1 10 0 12 13 9 13 10 9 1 12 5 1 9 2
23 1 16 11 4 13 9 2 13 15 3 3 1 2 16 9 3 4 13 1 9 7 9 2
24 9 11 11 11 2 15 1 9 13 12 9 2 4 1 12 9 13 0 9 1 11 7 11 2
6 13 9 2 12 9 2
12 7 10 0 7 13 9 13 3 3 1 9 2
17 15 13 2 16 15 3 4 9 7 9 2 15 4 13 9 1 2
33 3 4 15 3 13 3 1 15 2 1 9 3 13 15 1 2 10 9 9 13 2 16 15 4 13 1 9 2 15 3 4 13 2
9 9 2 15 13 9 1 0 9 2
23 10 0 9 1 11 9 4 1 0 9 13 1 10 9 1 15 1 11 11 0 0 9 2
27 7 1 3 0 9 4 15 3 13 2 16 9 2 13 2 15 1 14 13 15 1 10 9 2 15 13 2
25 11 2 9 1 9 1 9 9 1 11 9 4 13 13 3 1 10 9 1 9 1 9 9 9 2
13 11 11 0 9 11 4 3 13 1 10 0 9 2
3 9 13 2
19 16 11 3 13 15 10 9 0 9 2 13 15 1 10 9 3 1 15 2
17 10 9 13 15 1 3 1 2 16 15 13 10 0 9 0 9 2
16 2 15 4 13 10 9 1 9 1 9 3 1 0 0 9 2
39 16 1 0 10 9 1 9 7 9 13 3 1 10 3 0 9 9 1 10 0 9 2 7 9 4 3 13 1 10 9 1 14 13 9 1 10 0 9 2
23 15 4 3 3 13 3 1 9 1 9 12 0 9 2 12 0 7 3 0 2 9 2 2
35 16 15 7 11 3 13 10 0 9 1 13 0 9 2 1 9 1 10 13 11 2 13 11 7 11 2 16 15 4 10 0 9 14 13 2
6 10 0 13 11 11 2
9 3 13 3 0 1 3 0 2 2
27 15 4 0 2 16 15 4 13 3 3 7 3 3 2 13 15 2 2 13 11 11 2 12 2 13 9 2
16 11 13 15 1 10 9 2 15 15 3 3 4 13 1 15 2
6 2 11 2 13 15 2
5 3 9 13 9 2
41 15 4 3 10 0 9 1 11 11 0 9 2 3 3 10 9 1 11 11 9 2 7 3 10 3 0 8 8 9 2 15 13 1 0 11 11 7 0 11 11 2
36 7 15 13 3 1 10 0 9 7 10 0 9 2 16 9 13 9 1 15 3 2 7 16 10 9 1 11 4 13 9 9 2 9 7 9 2
15 2 15 4 15 2 15 13 11 2 13 11 15 14 13 2
29 15 4 3 1 0 13 15 3 1 0 9 1 9 7 9 2 7 15 4 3 13 14 13 10 9 1 9 3 2
16 15 4 3 4 3 2 16 9 13 9 7 9 3 1 9 2
19 10 0 9 4 15 13 2 7 0 9 4 15 13 1 9 13 3 3 2
30 15 13 10 0 9 1 9 2 3 9 4 0 7 0 13 1 10 0 9 2 15 4 13 9 3 2 13 11 11 2
23 9 2 11 12 2 4 3 1 12 7 4 3 10 0 9 2 15 4 4 13 1 0 2
38 7 4 13 10 0 9 1 0 9 2 9 1 9 1 0 9 7 9 2 0 9 1 0 9 7 3 0 9 1 0 9 2 0 9 1 9 3 2
8 3 10 9 13 15 1 0 2
67 7 13 15 9 1 9 9 2 10 0 9 9 7 9 9 2 7 13 15 9 1 10 0 9 9 2 9 9 7 9 9 2 9 9 7 9 9 2 16 13 15 1 15 2 15 13 9 9 2 15 4 13 1 14 13 2 15 15 13 2 3 3 1 10 0 9 2
23 9 2 15 13 3 1 9 2 4 3 3 3 0 7 0 2 13 10 9 8 7 9 2
18 9 4 3 13 10 0 9 1 11 2 13 9 7 13 9 1 9 2
20 11 9 2 11 11 11 2 3 15 4 0 1 9 2 4 13 10 0 9 2
19 15 4 1 0 9 13 2 16 9 4 3 0 2 7 16 15 4 0 2
8 2 15 4 15 3 13 1 2
14 7 0 4 9 2 3 16 15 4 0 1 10 9 2
6 0 13 3 1 9 2
2 0 9
16 15 13 15 3 9 7 9 1 14 13 2 2 13 11 11 2
6 15 4 3 13 9 2
17 15 4 3 10 0 9 2 15 4 13 9 9 1 9 1 9 2
4 3 10 9 2
1 9
30 7 15 4 4 13 9 1 9 2 16 9 4 13 10 0 9 7 10 0 9 2 7 3 13 15 3 0 1 15 2
10 2 15 4 11 2 15 13 1 15 2
12 13 9 3 2 16 15 13 14 13 0 9 2
10 7 3 13 9 1 9 3 1 9 2
11 7 1 0 0 4 10 0 10 3 0 2
24 10 9 13 3 1 2 16 11 11 3 12 9 1 10 13 9 1 9 13 15 1 10 9 2
29 13 3 2 3 11 11 2 9 1 9 2 9 2 2 1 11 1 9 2 2 13 15 2 2 9 4 3 0 2
13 10 0 9 4 13 1 10 13 9 9 1 9 2
2 3 2
35 15 4 9 0 2 0 9 3 2 2 13 11 9 2 11 11 2 3 1 11 1 10 0 9 1 10 9 7 10 9 0 9 1 9 2
7 2 10 9 2 13 15 2
18 2 1 9 1 9 1 11 1 3 2 13 3 3 12 9 1 11 2
32 15 9 4 13 3 1 10 9 1 14 13 15 3 0 2 2 13 9 2 3 4 9 2 15 13 9 7 9 1 15 9 2
29 3 1 9 13 9 14 13 3 1 10 0 9 1 2 16 11 9 1 9 11 3 3 4 13 9 1 9 9 2
9 9 13 1 9 1 10 0 9 2
15 7 9 13 3 1 15 12 2 13 9 7 9 1 9 2
16 9 4 0 1 11 0 13 9 2 15 13 1 11 1 11 2
31 10 9 1 12 9 1 9 9 2 3 9 1 9 1 9 3 13 10 9 1 10 0 9 2 4 3 3 13 1 0 2
36 11 13 1 10 0 9 2 15 15 13 10 9 2 7 13 1 2 16 15 4 13 1 9 7 3 13 3 1 9 2 16 15 13 1 9 2
49 9 4 3 13 15 15 1 9 2 7 1 14 13 9 1 10 9 1 9 1 10 0 9 2 2 13 11 11 2 15 4 13 9 1 9 1 10 0 9 2 3 9 1 9 4 10 0 9 2
8 15 13 3 2 15 4 0 2
34 2 1 9 2 2 13 15 2 7 0 2 1 10 9 2 2 15 4 3 3 13 15 3 1 9 3 2 13 15 15 4 9 2 2
45 2 15 4 13 1 9 2 7 4 1 15 13 2 16 15 3 4 4 13 9 1 11 2 16 15 4 4 13 10 0 9 1 11 0 9 1 11 7 11 2 2 13 11 11 2
10 7 9 4 3 13 10 0 9 3 2
8 2 15 4 0 2 13 11 2
22 9 13 3 9 2 16 15 13 9 7 4 13 1 14 13 3 1 14 13 1 11 2
29 7 10 9 13 2 16 15 4 4 3 3 0 2 16 9 3 13 2 16 15 4 13 9 2 2 13 11 11 2
26 1 9 1 9 9 1 0 11 11 4 11 0 3 1 14 13 9 3 2 11 2 1 12 1 9 2
35 11 13 3 2 16 3 3 4 13 0 9 2 16 15 13 9 2 16 0 9 4 4 13 1 14 13 9 1 13 9 1 10 0 9 2
13 3 13 15 0 9 1 10 0 9 1 0 9 2
23 15 13 3 9 1 11 7 13 2 16 15 4 13 9 1 10 0 9 1 14 13 9 2
36 7 3 13 3 10 0 9 1 2 16 15 13 1 9 1 9 2 15 4 13 3 3 14 13 1 11 9 1 12 13 9 2 2 13 11 2
24 2 9 2 9 7 0 9 4 13 1 0 9 2 9 13 3 3 13 2 7 15 4 0 2
34 15 13 3 1 11 0 9 1 0 9 2 15 13 1 9 2 7 9 9 1 12 9 1 10 0 9 11 7 11 1 3 12 9 2
18 9 13 3 1 9 1 9 7 13 9 1 11 11 1 11 1 11 2
22 10 0 13 9 1 9 1 9 4 15 2 16 9 13 15 1 9 1 10 0 9 2
8 7 15 4 15 3 3 13 2
12 3 13 3 0 13 2 15 4 13 9 2 2
3 11 11 11
14 11 1 12 13 3 1 10 12 9 7 12 13 9 2
8 2 9 1 11 4 3 0 2
34 2 15 13 14 13 2 15 15 13 1 9 7 13 2 7 4 13 2 2 13 11 11 2 15 13 0 9 9 1 9 7 1 9 2
45 11 11 11 1 0 9 2 0 9 1 0 9 2 0 9 7 0 9 1 9 2 13 3 1 10 0 9 2 0 3 15 13 13 10 0 9 9 3 1 9 2 7 9 13 2
4 0 9 1 11
19 2 15 4 3 3 10 9 2 3 3 2 13 11 7 8 10 9 3 2
32 9 13 2 16 11 3 4 13 11 7 10 10 9 1 14 13 11 1 10 9 2 3 11 13 2 16 15 13 9 1 15 2
19 10 8 9 4 1 0 9 13 1 0 9 1 11 7 9 11 1 11 2
29 15 4 3 1 9 1 14 13 9 3 1 9 7 13 3 14 13 11 2 16 11 4 13 15 10 9 1 11 2
9 4 15 13 3 3 1 11 11 2
34 9 13 1 0 9 2 3 0 0 2 1 10 9 1 9 1 9 2 7 3 4 15 3 10 9 2 11 11 3 7 0 4 13 2
59 13 1 9 2 3 15 4 13 1 10 0 9 2 13 11 11 11 1 10 3 13 3 0 9 1 9 1 10 3 0 9 2 3 9 1 14 13 13 9 0 1 9 4 3 0 2 16 3 3 13 9 1 14 13 15 1 0 9 2
22 15 4 9 1 9 9 7 4 3 0 7 0 2 16 15 0 10 9 4 13 15 2
21 3 4 15 3 0 14 13 15 3 1 9 9 2 16 15 3 13 10 0 9 2
13 15 13 3 10 9 2 7 15 13 9 3 3 2
31 10 0 9 1 9 7 9 2 15 13 14 13 10 0 9 11 11 2 4 3 13 9 3 1 10 9 1 14 13 9 2
16 3 9 7 0 13 2 7 15 4 10 9 2 15 13 9 2
32 1 10 9 2 11 7 10 0 9 2 15 1 0 9 4 13 15 0 14 13 9 1 0 9 2 13 3 0 9 1 9 2
10 2 15 13 3 15 2 2 13 11 2
21 9 4 13 0 2 7 3 13 3 9 1 9 2 16 15 13 1 11 0 9 2
19 2 7 3 13 15 3 10 9 2 3 1 15 4 9 7 13 1 9 2
22 9 13 15 3 1 9 2 15 15 3 13 9 9 14 13 1 9 2 3 1 9 2
7 10 0 9 4 3 13 2
6 1 11 11 2 9 2
27 1 10 0 9 1 10 8 9 4 10 0 11 11 11 13 0 9 1 10 9 1 14 13 9 7 9 2
37 1 9 13 10 0 9 3 10 9 3 1 11 2 11 2 11 7 11 2 0 9 1 10 0 9 1 10 0 11 2 15 13 3 9 1 9 2
15 15 13 9 7 9 7 13 1 10 9 1 10 0 9 2
19 0 2 16 9 4 13 9 1 9 2 15 3 4 13 3 3 3 3 2
26 9 13 2 16 11 11 1 10 9 4 13 10 3 13 0 9 1 10 9 2 11 7 10 0 9 2
5 3 15 4 15 2
26 10 9 2 9 7 9 1 9 7 9 2 3 10 9 1 9 1 9 2 4 9 9 1 14 13 2
31 7 0 1 10 3 12 9 2 15 4 13 1 10 9 2 3 4 9 1 2 4 16 15 13 1 10 9 1 0 9 2
11 13 9 2 9 7 9 1 1 9 12 2
36 10 0 9 13 15 2 2 9 13 10 9 2 1 9 13 9 2 2 10 10 9 2 2 16 9 4 10 9 2 3 4 0 9 0 2 2
12 13 9 4 3 13 15 1 0 9 1 9 2
33 9 13 2 15 9 1 11 9 13 2 7 15 4 2 3 13 2 3 13 1 0 9 1 15 4 13 1 9 1 9 7 9 2
9 3 3 4 10 0 9 13 3 2
9 9 3 13 15 10 9 1 11 2
35 16 15 4 13 4 0 14 13 2 7 11 11 13 15 3 1 10 3 13 9 2 3 9 1 11 11 2 11 7 11 11 13 1 9 2
74 1 10 0 15 2 15 13 15 1 9 9 4 13 9 11 11 7 11 11 2 9 11 11 7 10 9 11 11 2 11 11 1 10 0 9 2 15 4 13 3 3 1 9 1 9 1 9 8 1 2 10 9 2 2 7 11 4 1 10 9 3 3 13 10 9 2 8 11 11 7 11 11 11 2
16 1 10 9 4 10 9 3 3 13 15 3 1 10 0 9 2
5 16 15 4 0 2
19 9 13 1 9 1 9 9 2 9 9 2 9 9 7 9 9 7 9 2
14 15 4 13 1 11 9 2 7 15 4 13 1 9 2
32 15 4 15 3 13 3 1 9 2 7 15 13 9 1 10 12 0 9 7 13 2 16 15 4 13 10 10 9 2 15 4 2
27 1 9 3 4 11 13 10 0 0 9 7 13 10 0 9 1 9 1 10 0 9 1 10 0 9 2 2
36 10 0 9 1 10 12 0 9 13 15 1 9 1 14 13 9 2 16 15 13 10 9 1 10 9 9 7 15 9 3 4 13 1 0 15 2
37 2 9 2 4 10 9 1 0 10 1 9 0 9 2 3 1 9 1 11 9 1 2 16 9 13 1 15 2 1 10 9 9 13 13 9 1 2
5 12 2 11 1 11
26 2 16 9 13 2 4 15 3 13 15 2 16 15 13 1 14 4 15 1 15 2 15 13 1 9 2
35 1 11 11 2 10 0 9 1 9 1 11 2 4 12 9 7 12 9 13 2 16 10 9 1 10 0 9 13 10 9 2 13 0 9 2
20 1 0 9 13 15 15 0 2 16 12 9 1 0 9 13 0 9 3 3 2
16 1 11 4 15 3 11 11 1 11 7 15 2 15 4 13 2
8 15 4 3 3 13 9 1 2
11 7 15 13 11 11 3 13 15 3 1 2
35 3 1 11 11 4 0 9 7 0 9 0 2 7 9 4 3 10 9 7 0 9 2 3 3 13 4 10 9 1 9 12 9 0 9 2
47 15 4 13 1 0 9 2 8 12 2 1 15 1 9 7 4 3 3 13 1 9 1 0 9 1 9 2 10 9 2 15 11 3 13 9 1 14 13 1 9 1 10 0 9 1 15 2
4 9 1 0 9
2 10 9
6 11 11 2 0 1 9
16 9 13 3 3 2 7 11 13 9 1 14 13 3 1 9 2
3 3 5 12
17 3 12 9 1 9 11 11 4 10 9 2 1 11 13 3 1 2
10 11 8 2 15 0 9 13 13 9 2
16 3 1 16 15 4 4 3 1 10 9 13 15 3 14 13 2
14 7 9 13 3 1 9 1 2 16 15 4 10 9 2
23 3 4 15 13 10 9 0 2 3 4 15 13 9 2 7 15 4 3 13 9 1 3 2
21 2 7 2 15 13 10 0 9 3 1 9 2 2 13 15 7 13 10 0 9 2
21 15 13 1 9 2 16 3 13 10 0 9 9 2 15 3 13 12 9 1 9 2
10 7 15 4 15 3 2 9 4 13 2
5 9 13 1 9 2
32 15 13 15 1 2 3 10 9 13 1 2 15 13 15 1 9 1 14 13 15 3 1 9 7 13 3 1 15 1 13 9 2
5 2 3 1 0 2
28 2 6 9 2 2 13 15 2 2 15 4 3 13 9 1 12 3 1 9 15 4 4 13 15 1 9 2 2
30 15 4 13 3 2 1 16 3 1 9 1 0 9 2 7 15 4 3 3 3 2 3 0 2 2 13 9 11 11 2
14 7 15 13 15 2 15 15 4 13 9 1 1 9 2
23 9 4 3 2 3 0 15 4 13 1 10 9 2 3 4 3 1 10 9 1 13 9 2
45 2 1 9 1 12 9 4 15 13 1 12 9 1 15 2 7 9 1 9 4 10 3 0 2 13 11 11 2 16 15 13 1 9 1 9 11 2 9 11 11 11 7 9 9 2
5 13 9 9 12 2
30 2 0 2 3 4 4 3 3 1 9 2 16 15 4 4 13 9 2 13 3 1 12 9 14 13 15 9 1 9 2
12 9 13 1 9 2 15 13 1 14 4 0 2
12 2 1 10 9 4 15 3 13 9 7 9 2
13 1 9 13 10 9 9 3 2 10 9 1 9 2
9 9 13 1 10 9 15 1 15 2
9 15 13 9 2 1 9 13 9 2
27 15 4 13 1 9 0 0 9 1 12 7 13 1 10 9 13 1 0 9 7 13 1 9 1 0 9 2
8 2 6 2 11 13 1 9 2
14 13 9 7 13 9 1 0 9 2 7 3 3 0 2
26 1 9 13 9 9 9 1 9 1 11 9 9 2 7 3 4 9 3 13 2 15 9 3 4 13 2
6 15 4 13 3 2 2
15 3 16 15 3 13 9 1 15 7 13 10 9 1 9 2
27 2 11 7 11 13 9 13 0 1 15 2 2 13 11 11 2 1 4 9 1 11 9 11 11 11 9 2
21 15 4 9 13 1 3 7 3 0 0 9 2 15 3 13 15 7 3 13 9 2
27 1 10 0 13 15 9 3 0 2 7 1 9 3 1 9 1 15 13 15 3 1 10 0 2 13 11 2
27 9 1 9 4 13 9 2 7 1 10 9 13 11 9 10 9 1 14 13 0 9 13 9 3 1 9 2
58 1 9 1 10 0 2 13 9 2 4 15 3 3 13 10 2 9 2 2 3 9 2 9 7 9 3 3 13 1 0 9 1 0 9 2 7 13 10 9 1 10 9 2 15 3 3 3 13 15 1 9 7 0 9 1 10 9 2
9 10 9 13 3 1 10 0 9 2
13 15 13 1 11 2 7 15 4 9 1 0 9 2
53 9 0 9 7 9 13 1 10 0 9 2 16 15 4 13 10 9 1 2 16 9 13 10 3 0 9 1 9 1 0 9 2 15 4 4 4 13 3 1 9 1 13 9 7 1 10 9 1 9 7 9 9 2
10 2 7 15 4 3 13 9 1 9 2
14 15 4 3 14 13 9 1 15 7 15 4 3 0 2
49 9 1 11 3 0 2 7 3 3 0 9 7 9 0 9 1 10 9 1 14 13 9 4 10 0 9 2 3 3 13 1 11 7 3 1 10 0 2 11 7 11 1 1 10 0 9 7 9 2
18 7 3 13 15 3 3 1 2 16 3 4 13 9 1 9 1 9 2
18 9 1 11 11 9 13 10 9 2 3 4 0 1 15 1 10 9 2
7 2 7 0 9 1 0 2
7 3 1 15 4 13 11 2
27 3 13 12 9 2 10 12 7 10 12 11 11 2 11 0 9 1 9 2 3 9 13 1 14 13 9 2
27 7 1 10 9 4 15 3 13 9 1 10 9 9 3 1 10 9 2 15 13 3 2 15 15 4 9 2
47 2 7 15 4 3 0 2 16 15 4 13 3 0 1 9 2 16 15 13 9 1 9 2 2 13 9 8 11 11 2 15 3 3 4 13 0 9 1 14 13 9 9 2 7 3 9 2
7 15 13 15 2 13 11 2
21 9 4 3 0 2 16 15 3 4 0 1 9 2 3 1 0 9 13 7 13 2
3 9 2 2
29 12 1 10 9 2 15 3 13 9 13 1 10 9 0 9 2 16 15 1 0 9 13 9 1 9 7 13 11 2
1 9
14 4 15 13 9 2 13 15 3 3 12 9 0 3 2
13 15 13 3 3 14 13 15 3 1 9 1 15 2
19 4 15 13 9 2 4 15 13 2 16 15 13 15 2 16 3 13 9 2
15 0 11 13 2 16 11 13 9 13 14 13 3 1 9 2
36 7 3 4 15 1 9 13 15 1 9 2 13 9 1 10 0 9 9 1 9 1 9 2 16 11 9 1 9 13 10 0 9 3 1 15 2
34 16 9 0 9 3 3 13 1 10 0 0 9 2 3 13 9 9 1 15 8 9 2 16 10 0 9 1 9 13 10 3 10 9 2
19 15 13 10 9 1 10 0 9 2 2 13 11 11 0 9 2 11 11 2
2 12 2
14 15 4 3 3 13 9 1 0 9 2 15 15 13 2
21 16 0 13 1 9 2 4 12 9 13 9 12 1 10 0 9 1 11 1 11 2
32 15 4 3 13 1 14 13 10 9 7 1 9 1 10 9 13 3 1 10 9 2 3 4 0 1 9 2 7 3 13 15 2
18 2 15 13 3 1 14 13 7 13 3 3 9 1 10 9 1 9 2
1 9
24 15 15 2 15 13 15 1 0 9 2 13 2 16 9 4 13 9 16 15 3 13 1 9 2
22 10 0 9 13 3 3 1 0 11 2 7 11 4 3 13 9 1 3 0 9 2 2
20 13 9 11 11 13 2 16 3 3 13 9 7 9 1 11 7 11 1 9 2
14 2 16 15 13 14 13 15 2 4 15 3 3 0 2
10 9 4 3 13 1 8 9 7 9 2
34 1 9 9 1 11 1 9 4 9 11 11 11 3 13 15 1 12 1 10 9 2 15 4 3 1 9 1 11 1 9 1 11 9 2
31 11 11 2 9 1 10 0 0 9 2 13 2 2 1 10 9 13 15 15 3 1 10 3 13 9 1 1 10 0 9 2
10 3 1 11 9 13 11 9 1 9 2
16 1 12 4 15 3 13 3 0 1 10 9 1 11 7 11 2
20 7 1 10 9 2 3 11 11 13 2 13 15 3 7 0 1 14 13 3 2
25 15 1 9 1 16 10 9 4 4 3 0 2 4 9 13 9 1 9 1 10 0 0 9 9 2
20 0 9 4 9 0 1 12 9 9 1 9 7 3 13 3 0 9 3 3 2
41 11 9 1 11 2 3 15 13 9 2 13 9 1 10 0 7 0 9 1 9 2 3 11 11 4 13 10 0 9 0 9 1 9 2 0 9 7 12 0 9 2
15 15 4 0 7 0 2 7 9 4 0 2 0 7 0 2
10 9 1 12 9 9 13 11 1 9 2
40 2 7 3 4 9 1 14 13 9 1 14 13 3 0 2 16 15 13 9 1 14 13 10 9 15 15 13 3 1 2 7 3 13 9 1 14 13 3 2 2
18 11 11 4 3 0 1 14 13 10 9 1 9 3 1 10 0 9 2
15 3 4 9 1 9 1 10 0 9 1 11 4 10 9 2
20 2 4 15 13 10 9 1 9 12 2 4 15 10 3 0 9 14 13 9 2
47 7 16 2 0 11 9 2 4 13 11 11 0 9 2 1 16 15 3 13 14 4 10 0 2 2 13 3 3 7 0 10 3 0 9 2 3 15 13 10 9 1 9 2 9 9 13 2
6 7 16 9 4 0 2
23 15 13 3 10 9 1 9 1 10 9 2 15 13 9 2 1 15 3 13 10 9 1 2
7 11 1 11 4 13 9 2
3 0 9 2
15 1 9 13 11 11 1 9 1 14 13 15 13 1 9 2
5 15 4 10 9 2
25 2 15 4 3 13 10 9 3 2 13 9 2 2 4 15 3 0 9 2 3 13 3 15 3 2
31 1 9 9 4 3 13 2 16 13 9 4 10 9 2 15 3 13 1 9 3 13 9 1 9 2 3 10 3 13 9 2
33 0 9 2 1 3 4 9 1 11 2 13 3 2 16 3 1 9 4 13 9 1 10 9 1 9 7 3 10 0 9 1 9 2
27 7 10 0 11 2 15 4 13 1 0 9 1 0 9 9 2 9 11 2 13 3 9 1 9 0 9 2
13 10 9 13 13 1 10 9 2 7 15 13 15 2
17 1 9 13 15 2 3 1 11 11 7 11 11 2 9 11 9 2
12 15 13 3 3 1 0 2 7 9 4 0 2
9 15 4 1 0 0 0 10 9 2
15 7 0 4 15 3 2 16 11 13 10 0 9 1 9 2
12 10 9 13 15 1 15 2 15 15 4 13 2
27 11 9 1 11 4 1 10 0 9 1 10 0 9 1 10 0 9 9 1 12 13 1 10 3 0 9 2
24 9 1 9 2 3 9 1 9 2 9 7 9 2 4 4 0 7 13 1 0 7 0 9 2
25 9 1 9 4 15 3 3 13 9 1 2 3 3 10 9 4 4 13 9 2 2 13 11 11 2
20 9 4 13 11 11 1 14 13 9 1 0 9 2 7 15 4 15 13 3 2
2 10 9
24 1 0 13 11 11 1 9 2 7 1 9 13 15 1 10 9 2 3 15 13 1 12 9 2
20 16 15 4 13 3 2 13 15 3 1 9 2 2 15 13 3 0 9 2 2
17 9 13 9 1 1 9 1 0 9 1 9 1 14 13 0 9 2
3 5 12 2
11 2 11 4 0 2 7 15 4 15 3 2
9 9 9 2 2 10 0 9 2 2
6 9 13 11 0 9 2
7 15 13 3 1 0 9 2
24 7 9 11 11 13 3 3 11 13 1 9 2 16 9 3 4 4 13 2 1 0 9 2 2
25 1 12 9 9 4 15 0 1 9 7 9 14 13 2 15 3 4 9 2 7 15 3 4 9 2
26 1 9 0 9 13 15 1 9 9 2 7 15 4 9 1 2 16 15 3 4 4 3 1 9 3 2
40 3 10 0 9 1 9 1 10 2 11 2 2 9 11 4 13 1 9 2 13 3 9 1 2 16 3 1 3 0 9 1 1 11 4 13 9 1 9 9 2
51 7 15 4 3 13 15 1 9 1 10 0 9 2 2 13 15 1 9 9 0 1 11 11 2 9 1 11 0 9 2 11 2 16 15 4 10 0 9 14 13 10 9 1 10 0 0 9 1 9 9 2
39 1 9 13 11 11 3 3 1 11 11 2 15 13 1 9 2 10 0 9 2 2 2 10 0 7 10 0 2 7 2 9 1 9 2 7 10 0 9 2
7 3 4 15 3 1 9 2
4 1 9 1 9
40 16 11 12 13 10 0 9 2 15 4 13 3 0 9 7 9 2 4 9 0 2 9 4 15 0 1 9 2 7 3 4 15 13 1 10 11 9 7 8 2
21 15 4 13 1 9 1 9 2 9 2 9 7 9 2 7 0 13 14 4 0 2
10 15 13 3 9 1 15 13 8 9 2
27 2 10 3 0 13 3 3 2 16 15 15 4 3 0 2 16 15 13 1 9 1 10 0 2 13 11 2
2 12 9
23 13 15 4 15 13 14 13 3 10 9 9 1 9 2 11 7 9 1 9 1 11 9 2
34 1 10 10 9 4 11 7 11 13 11 0 9 1 10 9 1 0 9 2 9 7 9 2 16 10 0 0 9 13 1 14 13 9 2
14 1 11 9 13 9 1 10 0 9 3 1 14 13 2
17 3 13 10 0 9 1 9 3 1 12 1 12 9 1 0 9 2
8 2 7 2 15 13 3 13 2
22 1 10 0 9 13 15 0 9 3 1 9 7 13 9 13 3 2 16 9 4 0 2
34 7 3 13 3 3 10 3 0 9 1 3 10 0 9 7 10 0 9 2 16 15 4 13 2 14 13 9 3 2 2 13 11 11 2
18 1 9 4 15 10 0 9 1 9 1 11 11 0 9 1 11 9 2
10 9 1 9 7 9 13 9 1 9 2
32 10 0 9 13 3 2 16 3 4 13 0 9 2 7 3 16 10 0 2 15 3 4 13 15 1 9 2 4 13 9 3 2
33 10 0 9 2 13 1 10 0 9 1 9 9 2 4 0 9 1 11 9 7 10 0 9 3 0 1 14 13 10 9 1 9 2
12 16 15 4 10 0 9 13 3 3 0 3 2
24 10 10 8 9 1 9 1 9 4 11 11 2 3 10 0 9 13 1 10 9 1 0 9 2
4 11 13 3 2
25 16 3 15 4 3 1 10 9 1 9 7 9 2 4 15 4 13 15 2 3 1 14 13 11 2
19 15 13 3 3 1 9 0 9 9 1 10 9 1 9 1 10 0 9 2
7 0 9 4 0 1 15 2
10 1 9 13 11 11 3 15 3 0 2
12 9 7 10 9 2 9 2 4 3 13 1 2
32 2 1 9 2 11 2 11 13 1 15 2 3 13 15 15 3 1 9 2 3 3 13 10 9 2 15 3 4 0 10 9 2
23 15 4 0 9 2 15 3 1 10 0 9 4 13 3 1 9 1 11 1 10 0 9 2
7 7 2 6 2 3 3 2
24 2 15 4 0 1 10 9 1 14 13 8 7 13 2 16 10 13 9 1 9 9 4 0 2
13 10 9 1 9 4 0 2 13 1 9 7 9 2
35 15 13 10 0 12 9 1 9 2 9 2 2 7 3 2 11 11 2 7 2 11 2 1 9 2 15 4 13 1 14 13 10 0 9 2
14 1 10 9 15 4 1 9 2 13 9 1 0 9 2
5 15 13 15 3 2
3 2 6 2
41 0 9 4 1 12 2 3 15 13 2 16 15 4 13 15 3 1 11 7 4 0 1 14 13 1 10 10 9 9 1 10 9 2 7 3 13 3 8 7 11 2
21 9 13 11 11 2 4 12 9 7 13 1 11 2 3 9 13 15 1 9 3 2
33 11 11 13 2 16 15 13 13 1 10 9 1 10 9 2 7 16 15 13 13 2 13 15 2 16 9 4 13 3 9 1 9 2
18 10 9 13 3 2 16 3 13 12 13 2 15 13 1 14 4 13 2
11 15 4 4 0 9 1 13 9 1 9 2
32 15 4 10 0 9 1 10 0 9 2 16 15 3 13 13 1 10 0 9 14 13 9 7 13 10 3 0 9 1 0 9 2
46 9 13 1 10 9 1 9 7 1 0 9 2 3 15 13 1 2 16 9 4 4 3 3 1 10 0 2 2 10 9 2 0 10 9 7 2 1 13 1 9 2 10 0 0 9 2
21 11 11 11 2 1 0 13 1 9 0 7 3 0 9 2 13 2 15 3 13 2
10 15 13 3 3 15 1 9 1 9 2
3 9 3 0
22 10 13 9 4 0 1 9 9 1 9 1 9 7 9 1 9 1 9 3 1 9 2
22 10 0 9 4 3 13 1 9 3 1 11 9 2 3 3 13 1 10 3 0 9 2
31 0 9 1 10 9 2 1 9 7 9 3 7 3 1 10 0 9 2 4 3 0 1 9 1 9 1 10 9 7 9 2
10 1 10 0 9 4 15 13 1 9 2
24 15 4 1 9 3 13 1 2 3 9 4 0 2 7 4 13 0 2 3 1 9 1 9 2
17 15 13 9 7 1 10 9 10 0 9 1 10 0 9 1 9 2
16 3 13 0 9 2 15 13 14 4 10 3 0 1 0 11 2
29 9 13 3 1 10 9 2 9 4 3 1 14 13 2 2 15 4 15 3 13 2 2 7 11 13 15 1 9 2
44 11 11 13 2 16 15 4 13 9 1 10 9 1 9 1 9 9 2 9 11 11 2 7 15 4 3 13 2 15 15 4 13 2 2 15 13 1 9 9 2 2 13 15 2
20 7 1 10 0 11 11 0 9 4 15 3 13 14 13 9 1 14 13 15 2
18 3 1 11 13 3 9 2 7 15 13 15 15 3 1 14 13 2 2
8 7 9 13 3 10 0 9 2
9 2 15 4 13 3 1 0 9 2
24 2 10 9 4 8 8 11 11 15 13 1 10 9 1 9 1 2 16 9 13 3 0 9 2
3 12 9 13
19 2 3 13 15 9 2 7 10 9 4 15 13 15 14 13 3 1 11 2
6 9 1 9 13 15 2
42 3 10 12 13 9 13 3 1 9 7 13 13 9 1 10 13 9 2 15 1 9 7 9 7 9 1 9 1 9 13 10 8 0 9 1 10 0 9 1 10 9 2
6 11 11 13 0 9 2
17 10 0 9 1 3 11 7 11 13 3 3 2 3 9 13 1 2
22 10 0 9 12 0 9 4 13 1 9 1 15 1 11 3 0 9 2 11 11 11 2
19 1 10 9 13 10 0 0 9 15 1 10 0 9 2 15 3 3 4 2
8 3 10 9 13 1 15 15 2
39 3 3 13 9 3 2 16 15 4 15 8 8 2 15 13 3 1 2 15 1 10 0 1 10 0 9 4 9 1 2 3 10 0 9 13 13 15 9 2
2 9 0
20 8 7 9 13 3 1 3 0 9 7 10 9 4 1 9 13 1 12 9 2
12 15 4 10 9 2 9 13 2 15 4 13 2
29 3 13 13 15 2 16 9 4 9 1 2 16 10 0 13 1 9 1 9 1 12 9 1 9 2 2 13 15 2
10 10 0 9 4 3 9 7 3 0 2
16 11 11 2 0 9 2 4 1 10 0 13 1 9 1 11 2
5 9 4 3 10 9
19 7 15 4 0 14 13 2 3 3 15 4 13 1 14 13 9 3 2 2
9 15 4 13 15 3 0 1 15 2
14 15 4 0 9 0 2 7 9 1 0 9 13 3 2
30 3 13 0 9 1 2 16 9 3 4 13 15 9 1 14 13 12 0 9 1 12 9 2 3 1 15 13 1 12 2
35 2 15 4 10 9 2 13 9 7 13 2 7 13 16 10 0 0 9 4 4 0 1 10 0 9 2 13 15 7 13 9 3 1 10 9
15 9 13 10 0 9 1 9 1 11 9 1 9 1 12 2
25 3 4 10 9 13 1 9 2 1 9 0 1 1 10 13 0 9 2 2 16 10 0 13 15 2
36 11 9 13 3 3 1 0 9 2 2 15 13 9 10 0 9 7 13 0 0 3 1 15 3 1 9 2 16 10 10 9 1 11 13 15 2
26 9 11 13 14 13 15 3 0 2 1 15 13 1 9 1 15 1 9 9 2 9 1 0 9 12 2
27 3 9 1 10 0 9 2 11 11 11 2 13 9 2 16 3 3 13 10 9 0 9 1 9 1 9 2
14 2 3 4 15 3 13 15 1 9 2 15 4 0 2
9 3 4 15 3 3 1 15 15 2
13 3 12 1 9 12 13 13 15 1 10 0 9 2
12 15 4 3 13 1 11 9 2 7 3 3 2
2 13 3
35 3 1 3 13 1 10 3 0 9 1 11 2 4 15 10 0 9 2 7 15 4 3 13 2 16 15 4 13 3 1 15 2 15 13 2
15 15 13 0 10 9 1 10 3 0 2 0 7 0 11 2
31 1 10 9 13 15 2 16 9 2 1 4 10 9 9 1 9 2 4 0 1 0 2 0 1 10 9 2 1 10 9 2
15 15 13 15 3 2 7 15 13 14 13 15 0 1 9 2
19 15 13 3 1 9 11 11 11 2 7 10 0 9 4 15 13 12 9 2
27 10 9 4 9 3 13 14 13 2 9 2 2 15 4 0 1 2 16 9 7 9 4 13 3 3 3 2
21 10 0 13 3 1 9 2 16 15 1 10 9 13 10 0 9 1 10 0 9 2
18 11 4 4 0 1 11 1 12 7 4 13 12 9 3 3 1 9 2
12 10 0 9 1 9 13 3 12 9 1 9 2
19 15 4 3 15 14 4 0 1 2 2 13 9 1 0 9 2 11 11 2
4 9 2 8 8
15 10 0 9 1 10 9 13 15 3 3 10 0 9 1 2
6 11 13 2 3 3 2
16 3 13 10 9 1 10 0 9 2 16 9 13 1 10 0 2
2 9 13
23 16 15 13 15 1 14 13 9 2 13 15 2 16 15 3 4 13 1 14 13 15 15 2
4 13 15 9 2
11 2 0 2 2 13 15 1 9 1 9 2
34 7 15 13 3 3 1 9 2 3 3 4 15 3 1 10 13 9 3 4 9 1 9 1 9 1 0 9 2 15 13 0 9 2 2
25 15 13 2 7 9 13 1 10 9 2 16 15 10 9 3 13 14 13 0 9 2 3 0 9 2
4 2 0 13 2
25 16 11 13 11 2 13 15 10 9 1 10 9 1 3 0 9 1 0 7 15 15 13 1 9 2
13 1 10 9 2 15 4 3 3 0 14 13 1 2
10 1 10 9 4 15 3 13 10 9 2
29 9 7 9 13 15 3 1 15 2 7 1 10 0 9 2 9 1 11 2 13 15 3 3 3 14 13 13 9 2
23 3 4 15 0 1 14 4 13 1 2 0 9 2 2 1 1 9 4 0 7 4 13 2
20 15 13 10 9 1 14 13 14 13 2 16 3 13 9 1 15 1 9 2 2
14 10 0 9 4 13 1 9 1 14 13 9 1 9 2
20 15 4 0 1 2 16 15 3 13 14 13 1 9 3 2 2 13 11 11 2
18 11 11 2 9 1 11 2 4 3 13 9 7 10 9 1 11 9 2
3 3 16 2
27 1 9 12 13 11 0 2 0 9 2 1 11 2 15 1 0 9 13 9 1 9 9 2 13 11 9 2
2 10 0
22 9 1 9 1 0 9 1 12 1 9 2 9 1 0 7 3 11 11 7 11 11 2
27 15 13 9 1 9 7 9 1 1 9 11 11 2 7 15 4 8 0 7 0 1 2 16 15 4 0 2
17 7 3 13 9 1 10 0 9 1 3 0 9 3 3 1 8 2
27 10 9 13 15 3 3 1 9 2 7 11 4 3 3 13 2 16 15 1 3 4 13 15 1 14 13 2
18 10 0 9 4 13 10 0 9 1 10 9 2 7 10 0 10 0 2
14 2 6 2 15 13 15 2 3 4 15 13 1 9 2
77 1 10 9 2 15 3 13 9 3 1 10 0 11 2 4 11 11 13 1 14 13 2 15 3 9 9 13 3 1 10 9 3 2 2 16 9 11 11 2 11 2 3 3 4 13 9 1 10 0 9 2 2 7 2 16 15 3 4 13 3 3 2 16 3 10 0 9 1 13 9 4 13 9 1 9 2 2
31 11 11 2 12 2 13 1 0 7 0 9 1 9 1 11 2 7 10 9 1 2 11 2 4 3 13 1 10 9 9 2
21 15 13 3 9 1 2 16 10 9 4 4 13 3 2 1 16 15 4 13 9 2
2 9 13
20 9 9 13 10 0 0 9 1 15 15 2 3 1 9 4 13 0 1 9 2
4 2 13 9 2
11 15 13 15 9 2 16 15 13 1 11 2
36 7 10 0 0 9 2 1 9 1 9 2 13 0 9 2 16 15 13 1 9 1 10 9 7 13 1 15 2 1 16 15 13 10 0 9 2
21 3 14 13 1 11 2 3 14 13 10 0 9 1 9 7 0 9 1 0 9 2
14 3 11 11 7 11 11 4 3 13 15 1 10 9 2
23 13 3 9 1 9 2 3 13 1 2 9 2 2 9 9 2 11 12 2 12 11 11 2
22 10 0 9 13 1 15 1 9 11 11 11 2 9 11 11 7 11 0 9 11 11 2
7 2 16 9 3 13 9 2
14 10 9 1 9 4 1 9 9 13 1 9 0 9 2
38 2 16 9 13 2 16 9 2 15 13 9 1 9 1 9 12 2 13 0 1 9 2 3 4 9 13 10 9 2 16 9 4 13 2 2 13 15 2
13 15 4 3 3 3 2 15 4 3 1 0 9 2
11 16 10 9 13 2 4 13 2 13 8 2
44 10 9 2 3 15 4 13 16 9 2 15 13 3 3 3 1 14 13 10 0 9 3 1 10 9 2 3 4 13 1 2 16 10 0 9 3 0 4 13 1 10 0 9 2
12 7 15 4 13 2 16 15 4 13 10 9 2
25 15 13 3 10 9 2 15 3 7 0 13 11 13 9 1 10 9 2 15 3 13 9 1 9 2
19 3 4 15 0 2 16 9 2 15 13 9 1 10 9 2 4 13 15 2
25 11 0 9 13 3 0 9 2 7 11 11 11 13 15 9 13 1 10 13 9 0 7 0 9 2
27 9 4 15 1 9 1 10 0 2 0 9 2 7 15 13 3 3 2 3 1 9 2 9 2 9 2 2
42 15 4 0 1 10 0 9 1 10 9 1 12 9 9 7 1 9 2 1 11 11 13 15 2 2 13 15 3 1 12 9 2 1 15 13 15 1 3 1 9 2 2
22 15 13 15 7 13 14 13 10 9 10 0 9 2 16 15 13 2 2 3 6 3 2
19 0 9 4 1 9 9 13 15 1 2 16 3 15 0 9 13 1 15 2
17 1 9 13 15 15 1 12 9 2 1 0 9 9 1 12 9 2
27 10 9 13 15 1 10 0 9 3 13 1 12 9 2 0 9 7 9 2 3 10 0 0 2 9 2 2
9 15 4 13 2 15 4 13 3 2
10 1 9 4 15 10 9 7 10 9 2
9 2 15 13 10 9 3 1 11 2
14 2 15 4 3 13 10 0 2 16 3 3 13 3 2
5 3 4 15 9 2
12 15 3 8 8 13 14 13 10 0 1 9 2
14 9 9 4 0 9 1 9 9 4 2 13 3 2 2
3 15 13 2
7 1 9 13 11 11 3 2
4 11 1 11 2
11 3 11 11 13 15 3 1 10 0 9 2
21 3 13 9 1 10 9 2 7 15 1 10 0 10 2 0 9 4 1 3 13 2
15 2 7 15 13 9 1 14 13 10 3 3 0 9 2 2
42 1 0 9 1 9 7 0 9 1 11 11 7 11 11 13 11 3 10 9 3 13 1 9 9 2 3 16 9 4 3 0 2 16 15 13 2 16 15 13 3 3 2
58 11 11 4 10 12 0 9 13 0 9 1 11 11 2 7 1 9 9 13 9 2 2 11 4 13 3 1 10 0 9 2 3 1 15 4 13 15 1 0 9 2 7 10 9 4 13 9 1 1 0 9 2 3 15 13 1 9 2
29 15 4 10 0 9 1 10 13 9 2 16 15 13 2 16 9 4 13 10 9 7 10 9 2 15 10 9 13 2
12 2 15 13 15 1 15 2 13 15 1 9 2
40 0 9 13 9 1 11 11 1 10 9 1 15 10 0 9 1 2 16 9 9 13 15 15 1 10 0 9 7 1 10 9 1 9 1 9 1 9 7 9 2
22 3 4 11 2 11 2 3 1 0 9 13 11 2 16 15 1 10 9 3 13 9 2
20 11 11 13 3 1 8 12 11 11 2 3 15 4 13 1 9 0 11 11 2
11 9 2 11 11 2 7 11 11 4 13 2
29 1 9 1 0 9 13 9 1 0 9 1 9 1 0 9 1 0 9 9 1 14 13 11 9 1 9 1 11 2
45 9 4 13 1 14 13 10 0 9 2 7 15 13 10 12 0 9 9 11 11 10 9 1 2 16 15 1 9 13 10 0 9 1 10 13 9 7 13 1 11 1 12 2 12 2
4 11 11 2 12
7 2 15 4 13 1 9 2
5 7 15 13 3 2
11 7 15 4 3 9 7 3 9 1 9 2
7 7 15 4 0 13 15 2
3 9 11 2
41 7 15 13 3 3 2 16 10 9 13 1 13 9 3 1 9 7 13 2 16 9 3 13 7 3 3 13 9 7 9 3 1 9 2 16 9 13 3 1 9 2
2 12 2
6 13 9 5 12 9 5
4 11 13 15 2
21 10 0 9 1 2 3 10 0 13 15 1 9 2 16 15 13 9 1 14 13 2
19 15 4 10 3 12 9 0 2 0 9 2 15 4 13 1 11 0 9 2
16 15 13 2 16 9 13 7 4 13 0 9 1 9 7 9 2
24 9 4 0 9 2 16 11 11 13 15 1 10 9 2 11 11 2 3 1 10 9 1 9 2
13 1 9 4 9 13 3 1 10 0 9 1 9 2
22 1 0 9 1 9 13 2 9 2 2 1 1 9 4 9 2 9 1 10 0 9 2
13 9 9 13 10 0 9 3 1 10 0 9 11 2
6 7 13 3 9 2 2
9 15 13 0 9 1 14 13 15 2
14 10 9 2 4 15 15 1 9 2 15 13 1 9 2
12 2 16 15 13 4 15 13 15 3 1 9 2
15 2 3 13 15 1 10 0 9 1 15 15 2 13 15 2
7 1 15 13 15 10 9 2
27 7 15 4 0 2 16 0 9 4 13 3 1 9 2 7 15 4 3 4 10 9 2 15 15 3 13 2
11 10 9 0 9 7 9 4 15 3 13 2
6 15 4 3 10 9 2
8 7 3 12 9 1 9 9 2
11 2 15 13 9 1 15 2 13 15 3 2
13 9 1 0 9 1 10 0 1 9 13 12 9 2
16 11 11 7 11 11 13 15 1 0 9 1 9 1 11 9 2
5 15 4 3 0 2
9 11 13 15 1 9 3 1 9 2
33 9 1 9 1 11 2 11 2 11 7 11 4 3 3 0 2 16 15 13 1 2 16 15 9 3 1 0 10 9 13 12 9 2
10 2 7 16 3 3 11 4 0 3 2
14 9 13 3 3 2 1 10 0 9 1 9 1 9 2
17 15 15 13 1 9 2 13 2 13 2 0 2 0 2 3 13 2
23 1 14 4 4 13 1 9 1 9 9 13 15 1 9 7 4 3 9 2 9 7 9 2
15 9 1 0 9 4 13 1 11 9 2 13 15 1 9 2
8 3 4 15 3 1 11 2 2
22 1 9 2 15 15 13 1 10 0 9 1 9 2 13 15 14 13 1 10 9 2 2
26 7 16 15 3 13 15 2 3 4 15 3 13 15 1 2 16 3 13 10 0 9 1 9 7 15 2
24 13 10 0 9 2 15 13 3 1 9 1 2 16 15 9 9 13 10 9 13 0 1 9 2
6 11 13 15 3 3 2
16 15 13 1 9 1 12 8 15 7 3 12 9 1 15 9 2
40 10 9 13 3 3 3 1 0 9 1 10 9 2 15 13 9 1 10 0 9 1 10 9 2 15 1 9 4 13 1 0 9 1 10 10 0 9 0 9 2
25 9 1 9 13 3 1 9 7 9 1 9 7 3 13 0 9 3 1 14 13 3 1 10 9 2
34 15 4 13 0 9 1 14 13 9 2 1 15 15 4 13 0 9 3 1 0 9 2 16 15 4 13 1 9 1 9 1 0 9 2
11 15 13 2 16 15 13 15 1 10 9 2
36 9 1 11 9 4 2 1 11 15 2 3 12 9 3 0 1 1 11 9 2 3 16 10 9 1 9 4 13 10 9 13 1 12 0 9 2
12 2 15 4 13 1 14 13 0 15 1 11 2
8 7 10 9 1 9 13 9 2
19 1 9 13 11 1 3 12 9 1 9 1 11 2 3 4 10 13 9 2
21 7 16 0 15 13 2 16 0 9 13 15 2 2 13 9 1 9 2 11 11 2
22 0 9 1 7 1 11 4 13 1 10 0 9 2 7 1 9 12 9 13 1 9 2
31 1 10 9 13 13 15 1 9 1 11 2 9 2 9 2 9 1 9 2 9 7 10 0 9 1 3 14 13 10 0 2
8 2 13 15 10 0 9 2 2
28 1 9 1 9 13 9 15 10 10 7 3 0 9 2 3 1 9 1 9 1 10 0 9 2 3 13 9 2
9 10 9 13 1 10 0 9 11 2
4 13 7 13 2
43 10 0 8 7 9 13 1 9 2 7 1 8 4 12 1 10 12 9 0 2 16 15 4 0 1 10 9 2 16 11 11 2 11 11 8 10 3 0 9 11 8 11 2
13 15 13 15 1 10 9 3 1 2 2 13 9 2
12 15 4 1 9 7 6 1 15 0 1 15 2
16 3 13 10 9 1 3 3 14 13 1 10 0 9 1 9 2
18 16 9 13 9 1 14 13 2 3 3 1 9 2 7 1 10 9 2
24 9 13 9 13 2 16 11 11 13 10 0 9 1 3 14 4 13 1 9 1 9 0 9 2
43 11 11 2 9 1 10 0 9 11 11 2 13 3 1 10 9 1 10 13 9 2 2 16 9 3 4 13 16 15 3 3 4 10 9 2 15 13 0 9 7 9 2 2
23 1 11 10 9 3 9 7 9 13 9 1 3 12 9 9 2 15 13 0 1 0 9 2
14 11 13 1 9 1 9 2 1 10 0 9 3 13 2
32 13 15 13 15 2 2 13 10 0 9 2 11 11 2 16 15 13 14 13 15 1 9 1 11 2 15 3 13 10 0 9 2
15 15 9 4 9 13 10 0 9 1 10 9 1 9 9 2
5 9 13 1 15 2
12 7 6 2 11 11 4 13 0 1 10 9 2
19 2 15 4 0 2 16 11 11 4 13 15 15 1 14 13 10 9 3 2
11 15 4 3 0 2 15 10 0 3 13 2
18 3 4 9 9 1 9 3 0 9 2 16 15 13 15 1 0 9 2
29 1 0 2 0 2 0 9 7 9 1 9 4 2 11 2 1 9 0 9 1 9 12 13 13 10 13 9 9 2
1 11
40 9 1 11 13 2 16 11 13 2 16 10 9 2 15 11 4 13 1 11 1 9 1 9 1 2 16 11 13 7 13 9 2 3 3 4 13 1 11 3 2
19 13 9 3 1 9 7 9 2 13 0 1 9 1 9 7 13 9 3 2
31 1 10 13 9 13 9 1 9 7 9 1 3 11 11 11 8 11 2 11 11 11 11 2 11 11 11 7 11 11 11 2
27 3 13 3 9 1 10 0 9 2 7 9 4 3 13 14 13 10 9 1 9 1 10 9 1 0 9 2
2 3 0
20 13 3 9 1 9 2 9 7 9 1 9 7 13 9 1 0 9 10 9 2
47 2 7 1 10 0 9 13 15 0 9 1 14 13 11 3 3 0 1 9 2 2 13 11 11 2 15 13 1 9 1 9 1 12 3 1 2 16 9 13 3 1 10 0 9 1 11 2
14 4 9 7 9 3 13 2 13 9 3 3 1 9 2
7 7 13 2 15 4 9 2
18 13 3 10 9 2 15 4 13 15 9 2 15 13 9 1 9 9 2
13 7 9 4 0 9 2 7 3 4 3 13 9 2
11 15 4 0 2 16 9 7 9 13 3 2
16 9 13 3 3 2 3 1 9 2 12 9 1 10 0 9 2
12 15 4 3 1 9 13 2 16 15 4 0 2
38 1 11 13 9 9 14 13 9 0 9 1 14 13 10 9 1 10 9 1 9 1 11 2 15 13 1 14 13 9 1 9 1 10 13 9 1 11 2
23 10 9 2 10 0 9 9 4 13 2 4 1 3 0 9 13 9 1 9 1 0 9 2
13 15 13 10 0 0 9 2 15 4 13 1 9 2
26 15 13 3 10 9 1 10 9 2 11 2 15 3 13 10 9 2 2 0 11 2 2 1 10 9 2
7 9 4 4 0 7 0 2
17 15 13 1 0 9 7 13 1 9 7 13 3 0 9 1 9 2
22 2 0 0 9 2 2 13 9 2 16 9 1 14 13 0 7 1 9 13 1 9 2
8 9 12 1 10 0 11 11 2
52 2 16 15 13 9 1 2 11 2 2 4 15 3 13 15 2 16 15 4 13 9 1 9 2 7 15 13 3 3 1 2 16 15 4 0 1 14 13 9 1 0 9 2 8 14 13 3 1 9 7 9 2
8 10 0 4 3 14 13 9 2
17 3 13 3 10 1 0 0 9 2 15 13 10 0 7 0 9 2
14 7 15 13 3 2 16 15 3 13 3 3 1 9 2
24 9 13 3 1 11 1 12 2 12 7 12 2 1 11 1 9 12 7 1 11 1 9 12 2
15 7 1 10 0 9 13 15 15 3 2 3 3 1 15 2
9 13 12 9 0 2 13 9 3 2
1 8
42 15 13 3 10 0 9 2 15 13 3 3 7 13 10 9 2 7 1 10 12 9 0 9 2 3 9 4 0 1 9 2 4 15 12 0 7 0 9 2 15 13 2
19 16 9 13 13 2 4 9 3 13 0 9 7 9 3 1 9 7 9 2
18 15 13 11 3 13 10 9 1 11 7 11 7 3 13 3 1 9 2
16 1 11 1 11 13 15 12 9 2 10 0 1 9 1 11 2
12 9 4 3 3 10 0 9 1 11 11 9 2
21 16 10 9 13 1 9 1 10 9 2 16 15 4 13 10 13 9 1 10 9 2
23 3 4 3 3 4 1 12 7 12 9 3 1 9 15 2 2 13 9 11 11 1 11 2
27 9 1 9 12 2 9 11 11 11 2 13 3 2 16 10 0 9 4 13 2 16 11 9 13 1 9 2
17 9 1 9 1 10 9 13 1 10 9 2 1 15 9 4 0 2
19 1 10 0 9 1 9 4 9 1 9 3 0 1 1 0 9 1 0 2
14 9 11 1 11 4 13 1 15 7 13 1 9 9 2
27 2 1 15 13 10 0 9 14 13 3 1 10 3 0 9 7 3 13 9 3 1 9 1 10 9 9 2
20 9 4 13 10 9 1 10 13 9 1 9 7 9 1 9 2 3 9 9 2
33 9 13 2 16 15 4 4 13 1 9 1 12 9 2 7 15 1 9 4 15 15 13 1 2 10 0 9 2 2 13 11 9 2
6 9 9 13 15 9 2
16 9 13 2 16 9 3 4 3 3 0 0 2 1 3 13 2
19 16 9 13 1 9 2 4 9 13 3 7 3 3 13 9 2 13 15 2
6 15 13 3 3 3 2
20 15 4 3 13 9 3 1 9 2 16 15 1 11 4 13 10 3 0 9 2
12 13 9 1 3 1 0 9 14 13 13 9 2
32 11 2 2 7 3 4 11 13 2 16 15 3 4 13 15 3 14 13 3 1 10 0 9 2 10 0 9 7 10 0 9 2
34 13 15 3 1 2 9 9 2 1 9 12 2 3 13 15 3 9 1 10 9 13 2 9 9 2 9 12 2 7 2 11 9 2 2
5 0 9 1 11 9
49 0 15 4 11 13 2 16 15 4 0 14 13 3 0 9 13 2 7 16 9 3 4 15 15 13 1 2 16 15 13 7 3 13 10 9 2 7 3 15 3 4 13 1 15 15 4 13 1 2
12 15 13 1 10 9 1 3 10 0 9 9 2
21 9 1 12 9 13 3 1 10 9 2 15 10 9 1 12 9 3 13 1 9 2
20 9 13 3 0 9 2 7 9 13 13 2 1 12 9 9 1 12 9 9 2
14 2 13 15 3 3 7 13 11 1 9 2 13 11 2
24 11 9 13 2 16 10 0 9 11 1 10 0 11 1 9 1 9 4 13 1 10 0 9 2
14 15 9 13 1 11 1 9 13 1 2 15 15 13 2
10 3 4 4 15 1 10 0 9 3 2
14 15 4 1 9 9 13 15 13 1 10 0 9 9 2
5 9 2 12 9 2
26 15 4 3 7 1 9 13 3 1 10 9 2 7 3 13 9 1 0 9 14 13 15 3 1 9 2
16 7 9 1 9 7 9 13 13 2 16 15 3 4 4 3 2
21 10 9 2 3 4 3 1 14 13 0 9 2 16 10 9 1 9 8 13 9 2
18 9 1 10 9 1 9 2 16 15 13 10 9 1 10 0 9 3 2
16 16 9 3 4 0 1 15 2 3 4 15 3 13 15 2 2
24 5 10 9 13 14 13 15 1 9 2 15 4 13 9 3 1 9 7 3 13 15 1 9 2
15 1 9 1 3 14 13 3 1 9 16 9 4 13 3 2
11 1 10 0 9 4 9 13 1 12 9 2
3 0 3 2
2 9 12
43 15 4 1 9 11 2 10 9 13 1 9 2 8 2 9 1 9 2 9 7 9 2 2 8 2 13 9 13 1 9 7 9 2 7 8 2 9 1 8 7 9 2 2
42 1 10 9 3 9 13 2 16 3 3 1 9 4 13 9 1 10 0 9 2 13 15 3 1 11 2 15 1 10 0 9 13 1 9 1 14 13 15 1 9 9 2
10 15 13 1 12 9 1 15 0 9 2
6 9 13 1 0 9 2
37 15 4 3 16 2 15 13 11 1 9 7 13 15 3 2 15 4 13 15 2 15 4 3 10 2 0 2 9 2 15 4 13 1 9 1 9 2
10 15 4 1 0 3 1 8 2 11 11
17 10 0 7 0 10 1 9 2 2 11 11 2 2 4 3 13 2
20 15 4 3 3 0 2 3 9 3 3 13 1 14 13 3 2 2 13 11 2
11 2 15 13 2 15 13 15 0 2 3 2
39 9 11 7 11 13 15 3 2 3 16 15 4 13 3 1 9 11 9 2 7 16 15 4 13 3 1 9 2 13 3 9 11 7 11 14 13 1 15 2
5 1 9 1 9 2
7 13 9 3 7 13 3 2
9 2 13 3 12 9 3 1 9 2
25 3 1 10 9 4 15 9 2 3 4 10 0 9 2 7 1 10 3 0 9 13 0 9 9 2
2 9 12
9 15 13 2 7 13 3 1 11 2
20 12 1 10 9 4 4 13 1 9 2 7 15 13 1 9 1 10 13 9 2
10 2 15 13 3 2 15 4 13 15 2
32 15 4 4 3 0 14 13 9 7 9 1 15 1 9 9 2 11 11 2 15 4 13 10 9 1 9 1 9 9 1 9 2
3 2 3 2
23 1 9 1 11 7 11 13 15 0 9 2 7 3 3 9 2 1 3 4 10 13 9 2
26 3 13 0 0 9 1 10 13 9 2 13 1 10 0 9 11 11 11 9 9 9 3 7 11 9 2
14 10 0 4 13 10 0 9 1 2 3 15 13 15 2
34 1 11 4 3 3 3 13 15 14 13 0 1 2 13 9 7 13 10 9 2 7 9 13 3 3 0 9 1 10 7 10 0 9 2
14 16 10 9 13 1 9 2 4 9 13 10 9 3 2
20 0 9 2 7 3 3 13 1 9 1 2 15 3 13 1 3 12 9 3 2
12 3 13 9 9 7 9 10 9 1 10 9 2
26 11 11 13 15 13 1 2 16 9 1 10 0 9 4 13 9 1 10 9 1 9 1 9 0 9 2
12 7 3 13 3 15 1 9 2 15 13 3 2
5 9 13 1 9 2
34 3 1 9 1 3 13 1 0 9 1 11 2 13 3 3 3 0 9 14 13 3 1 2 15 13 10 3 0 9 1 9 1 9 2
10 2 15 13 3 2 3 15 13 15 2
7 15 4 3 4 10 0 2
9 9 1 10 9 1 3 12 9 2
13 10 0 9 1 9 1 9 4 4 10 13 9 2
27 12 9 3 2 16 15 13 1 9 2 3 1 15 1 9 1 9 4 13 9 1 14 13 9 1 12 2
13 15 13 3 3 3 3 2 16 15 13 1 9 2
16 2 15 4 1 0 9 13 0 0 1 11 2 2 13 15 2
22 3 13 10 9 1 12 9 1 11 0 9 1 9 1 10 0 11 1 9 1 11 2
11 16 10 9 13 1 0 9 7 9 13 2
6 13 9 5 12 9 5
33 15 13 3 2 16 2 11 4 13 1 10 0 9 1 10 0 9 7 1 10 9 2 15 4 13 10 0 9 1 10 0 9 2
39 2 15 4 13 1 9 2 16 15 4 13 15 1 9 9 2 7 4 0 1 14 13 3 7 13 9 1 14 13 2 16 3 13 9 2 2 13 11 2
12 2 15 13 3 3 3 10 9 2 13 9 2
40 9 13 1 9 13 2 7 3 1 0 4 3 0 2 3 13 15 3 2 16 11 11 11 7 10 0 9 4 13 9 1 14 13 10 9 1 10 0 9 2
19 15 13 15 1 2 7 4 15 13 15 1 14 13 9 1 14 13 3 2
29 15 4 10 0 9 2 16 9 1 0 9 1 10 0 9 1 9 4 13 1 9 1 9 9 7 9 1 13 2
7 3 4 11 11 9 15 2
10 15 13 2 16 9 4 4 10 9 2
13 3 13 15 9 2 7 11 4 3 1 14 13 2
29 11 11 2 15 1 12 9 3 13 1 12 9 1 0 9 1 0 9 2 4 10 9 13 3 14 13 1 9 2
29 9 1 9 9 1 9 13 2 16 3 13 3 1 2 0 9 2 1 9 1 2 0 9 2 2 7 3 0 2
11 7 16 10 9 4 13 3 1 11 9 2
20 2 15 4 3 0 1 14 13 1 11 7 4 13 10 9 1 9 12 2 2
11 9 13 0 7 0 2 16 3 0 3 2
26 9 9 13 2 16 0 9 1 0 9 4 4 3 1 14 13 10 0 9 13 9 1 9 1 9 2
15 9 2 15 13 3 1 9 2 13 1 9 1 0 9 2
33 9 1 9 1 14 13 1 9 13 2 7 15 13 9 1 0 9 3 2 2 15 13 1 10 9 1 10 0 2 16 9 13 2
26 15 1 15 4 3 4 10 0 9 2 15 4 13 10 0 9 11 11 1 14 13 10 12 0 9 2
32 9 13 3 13 2 0 4 3 13 1 9 2 3 16 15 3 4 13 1 10 9 1 10 9 11 2 1 15 13 3 1 2
33 9 13 3 3 9 1 9 1 11 2 11 7 11 2 7 11 11 13 3 1 2 16 0 11 4 4 10 0 9 1 10 9 2
23 1 10 9 4 9 13 1 9 1 10 0 9 2 15 13 10 9 1 0 9 7 9 2
49 2 10 9 13 2 16 0 9 4 13 15 13 1 9 7 13 1 15 15 2 16 10 9 4 13 1 9 2 16 15 3 13 15 2 2 13 10 9 1 0 9 2 11 11 1 9 11 11 2
31 11 4 3 13 1 0 9 2 3 2 11 12 11 7 11 11 11 8 2 0 7 0 9 1 0 9 1 0 0 9 2
28 10 9 1 9 1 9 13 2 16 0 9 8 1 12 13 12 9 2 7 9 13 1 12 9 1 0 9 2
26 10 0 2 2 15 4 3 13 15 3 2 16 16 15 13 1 9 2 3 13 15 1 9 7 13 2
5 13 9 9 12 2
19 10 0 9 13 1 9 2 9 2 9 2 9 2 9 2 9 7 9 2
14 12 9 1 2 16 9 4 13 9 2 4 15 13 2
9 1 10 9 13 11 9 12 9 2
21 9 13 3 1 2 16 15 3 3 4 13 0 9 3 1 14 4 13 10 9 2
22 1 9 9 13 11 11 3 9 2 2 4 15 3 0 14 13 1 10 0 9 2 2
30 15 1 9 1 10 9 4 0 9 1 15 1 10 0 9 2 7 1 0 9 4 15 0 14 13 10 9 1 11 2
13 7 15 13 3 1 14 13 3 2 2 13 15 2
18 2 11 2 13 2 16 15 1 10 9 3 13 15 1 10 0 9 2
24 15 13 9 11 11 2 15 4 13 1 9 1 9 1 9 1 12 2 7 3 13 1 9 2
10 3 10 9 0 9 1 11 11 9 2
15 10 0 13 15 3 0 2 7 15 4 4 0 1 9 2
24 1 9 1 11 9 12 9 9 13 0 9 10 9 2 16 15 4 13 10 9 1 12 9 2
13 15 13 10 9 1 9 1 9 1 9 9 12 2
16 15 13 2 16 9 4 13 2 7 16 3 13 0 1 11 2
24 15 13 1 9 1 9 9 2 15 4 13 2 7 3 1 16 11 4 13 1 9 1 9 2
21 0 9 4 4 10 9 1 2 16 9 1 9 4 0 1 9 1 11 7 11 2
15 15 13 1 9 2 10 0 9 11 11 13 9 1 15 2
17 11 9 4 2 1 9 11 2 1 9 11 2 2 13 10 9 2
16 7 1 10 9 2 15 4 13 9 1 9 7 13 10 9 2
34 9 4 13 1 10 0 1 0 9 2 7 16 15 3 4 13 15 2 4 15 13 10 0 1 15 14 13 9 2 2 13 11 11 2
9 15 4 13 15 7 13 1 15 2
13 3 13 3 3 10 9 3 8 13 3 1 9 2
10 2 6 2 9 2 15 13 15 3 2
22 15 13 1 0 9 2 7 15 13 3 14 13 1 9 2 16 9 4 13 0 2 2
10 15 13 1 10 0 9 7 13 3 2
18 3 4 15 13 15 3 2 7 15 13 1 14 13 3 3 1 9 2
27 2 9 4 13 15 1 9 2 7 9 2 15 3 13 1 11 2 13 1 11 11 1 10 9 9 2 2
11 15 4 13 9 1 9 1 0 0 9 2
20 7 4 9 1 11 11 11 0 9 0 1 9 2 4 15 15 3 1 9 2
8 11 2 9 13 7 9 13 2
18 10 9 4 4 15 1 10 12 0 9 1 2 9 9 7 9 2 2
30 3 13 10 0 9 3 2 0 9 2 2 15 4 13 1 10 9 2 13 10 9 1 9 1 9 1 10 10 9 2
32 15 13 15 13 7 13 2 16 15 13 1 14 13 9 1 10 11 2 3 15 4 13 3 13 10 9 1 3 10 0 9 2
24 11 2 0 0 9 4 10 0 9 13 9 1 11 1 11 2 7 3 13 12 3 1 9 2
4 9 7 9 2
49 7 1 10 0 9 1 9 4 15 13 2 16 10 0 9 1 9 3 4 13 12 9 1 9 2 7 16 9 1 9 4 0 1 3 0 9 3 13 7 16 15 13 15 1 9 7 0 9 2
12 15 4 3 4 13 1 14 13 10 0 9 2
18 3 13 3 0 9 1 14 13 10 0 7 10 0 1 9 1 9 2
15 15 13 3 15 1 9 7 9 14 13 2 7 9 3 2
17 15 13 10 9 3 2 1 15 13 11 3 4 13 1 9 1 2
30 11 13 3 1 12 2 7 1 9 13 11 3 1 12 2 7 1 0 9 13 3 9 1 10 12 9 1 9 9 2
11 3 13 15 13 3 1 15 2 13 15 2
11 10 10 9 4 15 13 3 1 9 9 2
9 11 4 13 1 12 9 1 9 2
52 2 11 11 2 13 10 0 9 1 11 1 11 0 9 12 2 7 3 1 10 9 4 11 11 11 2 9 1 9 2 13 15 0 1 9 2 16 9 4 4 0 1 14 13 1 9 0 9 2 13 9 2
10 3 1 9 4 15 1 10 9 3 2
14 9 13 3 1 14 13 3 1 9 3 1 10 9 2
9 11 11 4 3 3 0 7 0 2
13 16 15 13 13 3 1 10 9 1 10 9 9 2
54 3 4 15 13 8 8 3 3 7 13 11 2 11 11 11 11 11 11 11 2 7 2 11 11 11 11 11 11 11 2 2 1 4 3 1 2 11 11 2 2 10 0 9 15 4 13 1 10 3 12 9 1 9 2
17 1 15 1 9 1 10 0 9 7 1 9 1 11 9 1 9 2
17 0 4 3 12 0 9 1 12 9 2 12 13 9 10 9 3 2
33 15 13 9 1 10 9 7 9 7 13 15 15 9 1 0 9 1 9 2 9 7 9 2 2 13 10 0 8 11 11 1 11 2
19 2 15 13 3 14 13 10 9 1 11 2 16 11 13 2 2 13 15 2
20 4 15 1 9 2 16 15 13 1 9 2 13 16 9 1 11 4 10 9 2
3 1 11 11
20 2 16 15 3 13 1 10 9 2 13 15 3 3 2 2 13 11 11 11 2
16 2 10 0 9 2 13 15 2 4 13 15 1 10 0 9 2
3 13 15 0
17 15 4 9 2 15 13 10 0 9 1 9 2 2 13 11 11 2
11 16 9 13 2 3 2 1 9 2 3 2
11 15 4 3 15 2 15 13 0 9 2 2
29 1 9 13 3 9 1 9 1 9 2 7 3 13 9 11 11 1 10 9 9 1 9 1 14 13 10 13 9 2
4 13 3 1 9
7 0 9 2 0 9 7 9
16 13 9 1 9 2 13 15 1 13 9 1 9 1 12 9 2
5 11 13 3 9 2
14 7 15 4 3 3 3 13 15 2 16 15 13 2 2
33 15 4 13 7 13 7 13 10 9 2 9 1 9 2 7 15 13 3 1 15 3 4 3 2 15 13 14 13 2 15 15 13 2
2 9 12
27 9 13 1 15 9 1 11 7 9 2 7 0 9 13 2 16 3 13 10 9 1 9 1 9 1 9 2
16 1 9 13 15 1 9 2 3 1 9 4 10 9 13 3 2
11 10 0 13 10 9 2 10 0 13 9 2
1 8
12 7 3 13 15 3 4 2 2 13 11 11 2
3 1 9 2
10 2 15 13 9 1 0 9 1 11 2
28 1 9 4 11 9 13 1 9 11 8 2 2 7 15 4 3 13 1 10 9 1 10 0 0 9 1 9 2
11 1 9 12 13 15 1 11 1 11 11 2
23 9 1 0 7 0 9 1 9 4 13 3 1 10 0 9 3 1 9 1 10 0 9 2
20 9 4 13 15 2 16 15 4 0 2 2 13 11 11 7 13 3 1 11 2
11 10 9 13 9 1 14 13 9 7 9 2
21 3 1 9 1 9 4 11 11 2 9 13 1 10 0 2 0 9 1 0 9 2
39 10 10 12 9 0 2 9 2 1 11 4 1 0 3 0 2 16 15 2 16 9 2 15 10 9 1 9 1 9 4 4 13 11 3 3 1 0 9 2
33 1 0 9 4 11 0 9 13 2 16 9 3 13 14 13 9 1 2 15 3 13 2 16 11 13 9 1 0 9 1 0 11 2
21 9 2 15 13 14 13 10 0 9 3 3 0 1 10 9 2 4 10 0 9 2
14 3 1 15 13 15 1 2 4 15 3 10 0 9 2
22 0 9 13 15 1 0 9 7 0 9 2 7 15 4 3 13 3 1 10 0 9 2
20 2 15 4 10 0 9 2 16 15 3 13 15 3 2 2 13 9 11 11 2
12 9 7 9 9 2 7 9 2 4 3 0 2
18 1 10 9 4 15 13 9 2 7 15 4 3 0 2 16 9 13 2
15 15 4 0 3 13 16 11 11 4 13 1 11 2 8 2
38 2 11 4 13 15 1 10 9 1 11 2 2 13 11 11 1 2 10 13 9 1 9 2 2 10 9 2 15 4 13 1 14 13 13 9 1 11 2
16 7 3 4 15 3 1 9 2 9 9 4 13 3 1 9 2
34 2 9 4 1 10 9 10 9 1 2 16 15 4 13 10 9 1 0 9 2 15 4 3 1 9 2 13 9 1 10 9 1 9 2
10 11 13 9 1 14 4 0 7 0 2
29 3 1 9 13 15 9 1 14 13 3 1 11 7 3 1 11 2 15 13 3 1 10 9 3 1 10 0 9 2
12 3 10 0 9 7 9 11 13 1 10 9 2
29 11 2 10 0 9 1 11 4 13 3 1 9 2 16 10 9 1 10 9 1 9 1 10 9 1 11 4 0 2
23 3 13 9 1 11 0 9 1 0 1 14 4 10 9 1 9 7 9 2 16 15 13 2
1 9
27 9 11 11 2 11 11 2 13 3 3 10 0 9 1 2 16 11 9 3 13 13 10 0 9 1 9 2
14 3 4 15 13 3 3 2 1 14 13 3 1 9 2
9 3 10 12 9 4 10 3 0 2
16 9 4 3 3 10 0 2 15 13 10 9 1 10 0 9 2
32 15 13 2 16 11 2 3 3 4 3 0 2 2 16 15 3 4 13 0 15 2 15 3 4 13 10 9 1 9 12 12 2
32 2 1 9 1 9 13 11 2 16 15 4 13 9 1 9 2 15 4 13 2 16 3 13 0 9 7 9 3 3 1 9 2
23 11 2 3 1 0 9 13 15 2 16 9 12 13 2 15 10 0 9 1 11 4 13 2
10 13 9 1 0 9 7 9 7 9 2
10 15 4 10 0 9 2 15 13 9 2
42 10 0 9 1 3 4 0 1 0 9 2 7 3 0 1 9 1 3 11 11 7 10 0 9 11 11 2 3 3 1 10 9 11 11 13 1 9 1 10 12 9 2
7 15 13 1 9 1 9 2
7 11 13 1 10 12 9 2
41 3 4 15 13 10 12 9 13 3 1 9 2 3 11 4 13 13 2 7 3 3 4 10 0 9 13 1 13 9 2 13 9 7 13 9 2 16 11 4 13 2
14 13 2 16 15 4 13 1 9 2 15 13 3 0 2
27 10 9 4 3 3 4 10 0 2 15 4 13 9 9 2 13 15 3 1 9 7 9 9 1 9 9 2
14 10 9 1 10 0 9 13 10 9 2 15 11 13 2
17 15 4 10 3 0 7 0 9 2 16 9 13 1 9 7 11 2
27 7 10 0 9 11 11 11 7 11 11 11 2 15 3 13 12 0 9 1 10 9 2 4 3 3 0 2
12 3 13 10 0 9 0 3 7 3 0 9 2
17 2 15 1 9 13 1 9 1 2 16 3 13 10 9 1 9 2
7 9 13 3 1 11 9 2
31 3 4 15 13 0 3 2 16 15 3 3 3 4 0 1 3 9 1 9 2 15 3 3 13 14 4 0 2 3 4 2
34 8 0 9 1 10 0 9 1 10 9 11 2 11 7 11 7 9 1 9 2 3 9 2 15 4 13 10 3 3 0 9 1 9 2
24 1 0 9 13 3 9 2 3 0 0 13 0 1 9 7 9 2 15 9 4 13 1 9 2
1 9
24 3 4 9 13 3 1 11 2 1 16 9 4 13 12 9 1 9 1 0 1 10 0 9 2
23 10 0 9 2 15 13 1 2 4 12 9 11 3 10 0 9 11 11 12 9 1 9 2
15 1 11 4 15 13 12 9 1 3 14 13 10 0 9 2
51 3 13 10 9 2 16 10 13 9 2 15 3 3 13 9 1 2 16 15 1 10 0 9 13 15 15 2 4 13 1 14 13 9 2 16 9 4 0 7 9 1 10 9 0 2 1 15 13 15 1 2
9 1 9 7 9 2 9 7 9 2
33 15 4 13 9 2 3 0 9 2 15 4 13 1 11 1 10 12 9 3 2 1 13 9 1 10 0 9 1 11 7 11 3 2
20 2 4 15 13 16 10 9 13 10 9 2 0 2 0 9 1 10 0 9 2
28 2 7 2 3 13 15 2 13 11 7 15 2 15 13 7 13 9 1 15 2 3 15 3 13 3 1 9 2
3 3 0 13
41 4 15 4 13 1 11 11 1 12 9 9 2 16 15 13 1 10 0 9 2 13 0 10 9 3 14 13 2 13 9 2 13 9 7 13 9 1 10 9 9 2
21 3 1 11 13 11 0 10 0 9 2 15 9 4 13 2 3 1 11 7 11 2
14 15 4 13 7 13 10 0 9 3 7 4 3 0 2
13 0 13 15 3 0 12 9 3 1 0 9 2 2
26 12 9 4 0 9 2 7 1 9 13 9 13 15 1 9 1 14 13 3 1 11 7 13 9 9 2
35 1 10 0 9 1 0 7 0 9 13 15 1 10 9 3 3 2 2 6 11 2 15 13 15 4 0 14 13 10 0 9 1 0 2 2
8 12 9 13 2 13 11 3 2
19 11 8 8 8 8 13 1 2 16 15 13 10 9 13 9 2 11 3 2
6 1 11 1 1 9 2
2 12 2
3 3 3 2
8 3 13 15 9 1 10 0 9
18 7 16 15 3 13 1 9 3 1 10 9 2 13 15 9 0 9 2
12 0 9 13 3 10 0 9 1 15 7 9 2
28 1 9 9 13 15 1 10 9 1 9 2 9 7 0 9 13 1 10 9 1 9 2 9 2 9 7 9 2
27 15 13 3 14 13 10 10 12 9 1 11 9 2 11 2 2 11 2 11 7 11 2 16 15 13 3 2
19 2 15 4 13 10 0 9 2 2 13 15 13 1 10 0 9 2 11 2
11 10 9 13 11 11 3 10 9 1 9 2
12 9 4 13 1 10 0 9 1 9 7 9 2
16 9 4 0 1 14 13 9 2 15 13 0 9 2 9 3 2
20 15 13 3 10 9 2 7 13 15 9 10 9 1 12 9 1 9 11 11 2
15 11 11 4 0 7 13 3 2 7 11 11 13 1 9 2
15 3 4 9 13 14 13 15 0 1 9 1 9 1 9 2
19 1 9 9 7 9 13 9 1 9 1 11 1 14 13 10 9 1 9 2
41 16 10 0 9 4 13 10 9 1 0 9 2 15 4 13 0 7 0 9 2 4 0 9 4 3 0 1 10 9 2 13 9 1 11 9 1 11 2 11 11 2
23 1 9 13 0 3 7 3 7 3 3 1 9 7 13 2 2 13 0 9 2 11 11 2
18 2 11 11 11 11 11 11 2 4 13 3 10 0 9 9 9 1 2
16 10 9 4 3 13 1 16 9 13 10 9 1 10 13 9 2
22 15 13 9 3 1 10 9 2 15 13 10 0 9 1 14 13 3 1 10 0 9 2
13 11 9 4 3 1 12 13 1 9 1 9 9 2
19 16 11 13 10 9 1 14 13 9 9 2 13 15 15 3 1 15 15 2
15 15 4 10 3 0 9 1 10 9 1 1 12 9 9 2
8 9 1 9 1 10 0 9 2
21 15 4 10 3 13 9 2 3 9 13 9 2 9 2 1 14 13 10 13 9 2
24 15 4 3 0 14 13 13 9 1 10 9 1 11 2 7 0 9 13 15 3 3 1 9 2
7 10 9 13 2 9 2 2
11 15 13 15 3 3 1 2 2 13 15 2
9 2 7 10 0 11 13 3 3 2
14 1 11 4 9 13 0 1 10 1 15 0 13 9 2
3 0 9 13
15 15 13 0 1 9 1 15 7 13 7 13 9 7 9 2
12 9 4 13 15 3 2 7 9 4 13 15 2
41 15 4 13 9 1 11 2 3 11 11 13 2 2 15 4 3 13 15 10 0 9 7 4 3 13 1 14 13 10 0 9 2 7 15 13 3 15 10 9 2 2
1 9
12 1 9 13 3 12 9 9 1 9 1 9 2
23 9 1 12 9 0 9 4 3 1 10 0 9 2 1 11 2 13 1 12 9 1 9 2
45 1 10 0 9 4 15 13 8 1 14 13 7 13 9 1 14 13 7 13 2 7 1 14 4 13 10 9 1 9 2 9 2 9 7 9 13 15 1 10 9 3 14 13 9 2
29 1 10 10 9 4 15 13 9 1 9 7 9 2 16 15 13 1 3 14 13 9 1 15 2 15 13 14 13 2
24 10 9 13 1 10 3 0 7 0 9 2 7 10 0 9 4 3 10 12 9 9 7 9 2
22 9 4 0 2 9 13 2 11 13 1 9 2 3 2 7 9 9 13 10 0 9 2
43 9 4 3 13 1 10 0 9 2 16 9 4 13 3 10 9 3 2 9 12 9 1 12 1 9 1 12 2 15 13 10 9 1 9 2 15 3 13 9 1 0 9 2
36 10 12 9 4 3 3 13 15 1 15 1 10 9 2 16 15 12 15 4 13 10 9 10 2 15 3 3 13 3 1 10 9 1 10 9 2
24 7 3 4 9 3 3 13 9 1 14 13 9 11 11 1 11 0 2 0 7 3 0 9 2
10 15 13 11 3 2 7 3 3 3 2
21 11 13 3 1 0 9 2 16 15 13 3 7 9 4 13 1 10 3 0 9 2
1 9
19 3 4 9 13 15 1 9 2 9 2 9 7 0 9 2 9 12 9 2
9 5 3 9 13 3 13 1 9 2
25 11 4 13 12 0 9 2 3 16 9 1 9 7 9 2 15 4 13 15 2 13 1 12 9 2
18 10 9 4 3 13 3 7 3 2 7 1 10 9 13 15 3 3 2
15 1 9 4 3 13 0 9 7 9 7 9 1 9 3 2
42 3 16 15 13 1 9 7 9 2 7 15 15 3 3 13 2 15 15 13 14 4 13 2 16 15 13 10 9 3 2 7 1 3 13 15 14 13 15 3 1 9 2
52 1 10 0 9 2 15 4 2 4 9 11 11 12 3 13 10 9 3 2 15 13 10 0 0 9 1 10 0 9 2 7 1 13 7 0 9 2 15 1 9 4 13 10 0 0 9 3 1 9 1 9 2
30 2 15 4 10 9 2 16 15 13 2 15 13 15 1 15 2 11 2 13 11 10 9 2 16 15 4 3 1 9 2
25 15 13 3 10 0 9 1 10 0 9 2 10 0 9 2 16 9 13 11 11 3 3 1 9 2
13 3 13 13 15 2 15 15 13 1 9 1 11 2
10 13 9 3 7 13 3 10 9 9 2
10 10 9 2 3 4 10 9 1 0 2
17 1 0 9 13 15 8 7 9 3 2 3 15 13 1 0 9 2
39 9 4 15 4 0 1 2 15 4 13 15 0 9 1 0 9 7 1 3 0 15 13 2 4 15 0 1 9 14 13 15 3 1 0 9 7 0 9 2
3 2 3 2
29 15 2 15 13 15 2 13 2 16 15 3 3 13 2 16 3 0 9 7 8 7 10 9 4 13 1 10 9 2
22 1 9 9 13 9 9 1 14 13 15 9 1 14 13 0 9 2 3 9 13 3 2
12 9 4 10 9 2 10 0 9 4 9 1 2
29 3 13 3 10 9 1 10 9 1 9 11 11 1 9 9 2 3 1 9 1 10 0 9 4 4 11 11 0 2
10 10 3 0 9 4 3 3 13 15 2
21 15 13 14 13 10 0 2 9 2 7 9 2 15 13 3 1 0 3 1 15 2
21 2 15 13 1 11 9 1 14 13 9 2 9 7 9 0 9 2 13 11 11 2
40 1 0 9 4 15 3 0 2 7 10 0 9 1 9 1 9 1 10 0 9 2 12 9 0 9 1 9 1 10 0 9 7 9 13 9 13 1 11 9 2
10 15 13 15 3 7 13 15 1 9 2
27 13 1 10 0 9 4 15 13 1 10 0 9 2 0 9 2 0 9 1 10 0 9 7 10 0 9 2
8 3 13 3 9 11 1 9 2
6 7 13 9 7 9 2
21 15 4 3 4 0 14 4 9 1 10 9 2 10 3 3 0 9 1 9 4 2
32 9 4 1 3 13 1 11 1 9 2 7 11 8 8 4 1 10 9 3 13 13 3 7 1 0 13 1 9 1 9 9 2
8 15 4 13 9 1 0 9 2
16 2 15 13 14 13 1 9 1 15 7 4 3 13 1 15 2
24 15 13 13 1 9 3 3 7 0 9 1 10 9 3 13 1 9 1 9 1 9 1 9 2
17 4 10 0 9 3 0 3 2 6 3 4 9 3 0 9 3 2
12 3 10 3 3 0 9 2 12 12 9 2 2
27 11 7 10 10 9 13 13 7 13 3 1 9 2 16 15 3 1 10 9 13 15 3 1 9 7 13 2
4 9 13 3 2
10 1 14 13 3 2 13 15 1 9 2
9 3 9 1 0 9 2 11 11 2
15 0 9 1 9 1 9 2 9 7 9 7 9 13 3 2
3 3 3 9
2 15 13
3 9 9 2
5 3 4 15 0 2
5 15 13 15 3 2
17 11 13 11 1 10 9 9 1 14 13 10 0 9 7 0 9 2
44 15 4 13 3 2 16 11 9 3 13 9 2 7 10 9 1 9 2 7 3 4 10 0 9 2 9 2 7 10 9 1 11 1 11 9 3 0 1 10 9 2 11 4 2
4 2 1 9 2
12 9 13 2 3 3 2 1 11 11 9 9 2
21 2 9 13 3 2 16 0 8 0 9 3 1 10 13 9 4 13 0 9 13 2
28 13 15 10 9 1 14 13 9 7 13 9 3 1 9 2 13 15 1 10 0 9 2 3 2 11 9 2 2
1 0
3 9 2 9
34 10 9 13 8 7 0 9 8 1 8 9 2 7 3 10 2 0 2 9 13 9 1 3 2 13 10 0 9 1 9 9 1 3 2
8 10 9 13 11 9 4 9 2
38 0 9 13 3 3 2 16 15 13 9 1 9 1 14 13 2 0 9 13 3 1 9 1 15 2 15 4 13 2 16 15 13 3 1 10 9 3 2
19 15 4 3 0 3 0 1 9 3 2 13 15 1 11 9 9 1 12 2
11 13 9 1 9 7 13 9 3 1 9 2
15 9 4 9 1 0 9 1 10 9 2 15 13 1 9 2
28 2 15 1 15 4 13 10 9 2 15 13 3 1 2 16 15 13 1 9 1 14 4 0 2 13 11 11 2
21 15 13 1 0 2 7 9 1 0 9 13 2 16 3 13 9 1 12 9 9 2
9 2 13 15 9 14 13 9 3 2
13 2 10 0 9 4 13 2 16 9 4 13 13 2
8 3 13 15 13 1 3 9 2
21 15 4 13 1 14 4 13 9 10 9 1 1 12 9 9 1 0 7 0 9 2
56 10 0 9 1 2 16 15 13 10 9 2 13 10 0 9 11 11 3 3 2 16 11 3 4 13 9 1 2 16 15 13 9 4 3 13 1 11 11 11 2 7 4 13 2 16 15 13 9 1 2 9 2 9 11 11 2
35 2 15 13 10 9 1 11 7 4 1 10 9 4 3 1 14 13 9 3 2 13 11 11 2 15 13 16 11 11 3 4 9 1 11 2
18 3 13 3 10 0 9 7 12 9 2 16 15 4 1 10 9 0 2
10 9 4 13 1 10 0 9 1 11 2
13 2 15 4 13 1 15 14 13 1 10 0 9 2
38 10 0 9 4 4 0 1 9 1 14 13 1 9 1 14 13 2 7 1 9 13 9 14 13 10 9 2 15 4 13 10 9 1 0 9 1 9 2
17 11 9 9 13 1 14 4 4 10 0 9 1 11 1 0 9 2
19 9 2 15 4 13 1 9 2 7 1 0 9 1 9 4 13 1 9 2
41 15 4 3 0 2 16 2 0 11 9 2 3 1 9 4 13 10 9 1 9 1 14 13 10 0 2 1 13 1 10 0 2 1 9 1 9 1 0 0 13 2
29 10 9 13 11 11 15 3 9 1 2 15 13 3 1 9 2 7 13 2 15 1 11 13 14 13 3 0 9 2
24 10 0 9 4 13 15 1 10 9 2 7 1 10 9 13 9 3 16 15 13 1 10 9 2
37 0 9 4 13 1 9 1 11 7 11 1 12 2 16 11 8 11 1 11 1 12 2 1 11 1 12 2 1 11 1 12 7 1 11 1 12 2
3 9 13 2
14 3 4 15 0 9 1 10 9 1 9 1 0 9 2
10 0 13 1 3 3 0 9 1 9 2
19 3 4 10 0 9 13 1 9 7 0 9 9 1 9 3 1 1 9 2
13 15 13 10 9 2 16 15 13 15 3 1 9 2
32 15 1 9 9 2 11 11 11 3 13 2 4 13 1 0 9 1 10 9 1 10 0 9 2 11 11 13 3 1 10 9 2
6 7 9 13 9 3 2
21 16 2 10 0 9 13 3 13 2 7 11 4 3 3 1 9 1 14 13 9 2
25 15 4 3 3 13 2 7 3 3 0 4 15 3 1 13 2 16 11 11 3 13 10 0 9 2
27 11 2 10 9 1 11 4 3 13 2 1 16 9 9 7 9 4 13 2 16 3 3 3 13 0 9 2
11 15 13 1 9 2 10 0 9 7 15 2
20 9 13 10 7 10 0 9 1 9 1 9 1 9 1 10 9 7 10 9 2
5 9 2 12 9 2
15 2 1 15 2 15 4 13 11 11 11 2 13 9 3 2
7 3 4 10 9 13 13 2
29 10 0 1 9 1 10 9 9 13 2 16 10 0 9 13 2 3 13 10 0 3 2 1 16 10 9 13 3 2
15 15 13 15 7 13 1 9 1 10 0 9 1 9 9 2
39 15 13 3 1 14 4 10 9 1 9 2 16 10 0 9 2 15 13 9 1 9 2 13 1 14 13 0 1 9 2 15 4 13 9 1 10 0 9 2
23 9 7 9 2 1 9 1 9 2 13 15 1 0 9 3 14 13 10 0 9 1 0 2
12 3 4 15 13 3 1 9 1 0 9 9 9
38 11 9 11 11 13 15 3 3 1 11 2 2 1 10 0 12 9 1 9 4 15 15 9 13 3 1 9 2 15 3 4 13 15 14 4 3 0 2
16 10 0 4 10 0 9 1 9 7 9 1 10 0 1 9 2
29 15 4 3 13 1 2 16 9 13 10 0 9 1 14 13 9 2 16 10 9 1 9 13 9 1 9 1 9 2
14 10 0 9 7 9 4 4 3 0 2 16 15 13 2
9 15 13 10 9 1 9 1 9 2
18 15 1 15 13 2 7 3 4 0 9 13 10 0 9 3 1 9 2
13 3 4 15 3 3 13 13 10 0 1 15 3 2
14 7 10 9 4 10 0 2 0 1 11 7 11 11 2
19 15 4 10 9 2 15 13 2 16 15 3 4 4 0 9 1 10 9 2
10 15 4 3 4 0 7 9 1 9 2
14 10 0 9 9 4 9 13 13 9 1 14 13 9 2
26 10 9 0 9 13 13 2 15 4 3 0 2 3 9 1 0 9 13 1 0 9 1 9 7 9 2
21 1 9 1 9 4 11 13 12 9 2 13 0 9 7 13 1 14 13 10 0 2
32 0 9 13 10 3 12 0 9 2 7 10 13 2 14 13 2 16 15 4 13 15 13 8 2 1 9 2 1 10 9 2 2
29 1 10 9 13 15 2 15 4 1 9 14 13 10 9 1 9 1 3 14 13 9 2 16 10 9 4 4 13 2
20 10 12 0 9 4 13 7 0 1 11 7 13 2 16 15 13 1 0 9 2
43 7 10 0 1 10 9 13 2 16 15 4 13 7 13 2 2 13 11 11 2 1 3 4 1 9 1 14 13 0 1 9 9 1 10 0 9 2 15 4 13 1 11 2
11 2 15 13 3 0 9 1 15 1 9 2
8 1 9 13 9 1 0 9 2
12 13 9 4 3 1 0 9 13 1 10 9 2
10 15 13 1 9 2 2 13 11 11 2
10 9 2 10 0 9 4 4 10 9 2
23 3 13 9 11 7 9 1 9 13 3 7 3 1 10 0 0 9 1 10 0 11 9 2
27 10 0 9 4 3 3 13 9 10 0 9 1 2 3 15 4 13 10 13 9 1 10 3 0 9 9 2
41 3 1 9 2 9 2 9 2 9 2 9 2 9 3 4 3 13 0 9 1 14 13 10 3 0 9 1 9 2 7 9 3 1 9 9 13 9 1 0 9 2
4 12 0 9 13
11 10 9 4 10 9 2 9 7 0 9 2
4 11 13 3 2
12 9 7 0 13 13 1 9 7 10 0 9 2
8 7 3 4 15 12 1 9 2
9 9 4 13 1 9 7 10 0 2
14 15 13 3 2 15 13 2 15 15 13 2 3 2 2
9 9 13 1 9 3 1 9 2 2
17 3 13 10 9 1 11 11 9 2 16 15 4 13 1 10 9 2
15 9 12 4 10 0 9 1 8 3 13 3 0 12 9 2
28 9 2 15 15 3 4 13 2 7 1 3 13 15 3 1 10 9 2 3 15 13 1 9 2 9 2 9 2
13 7 15 4 0 14 13 10 9 2 2 13 15 2
14 3 13 15 8 2 8 2 1 9 1 2 8 2 2
5 11 13 1 9 2
14 1 9 13 15 1 9 2 16 15 4 13 0 9 2
8 3 3 1 10 0 0 9 2
16 12 0 9 2 15 2 15 1 10 9 2 13 10 0 11 2
21 7 15 13 2 16 10 0 9 9 13 1 10 0 9 2 16 10 9 13 9 2
13 3 4 9 9 2 1 9 2 3 0 1 9 2
13 15 4 15 13 3 13 7 13 9 2 13 15 2
14 13 10 9 1 9 2 9 7 9 2 4 15 0 2
25 15 13 1 10 3 0 9 1 10 0 9 1 11 11 11 11 1 11 2 10 0 9 11 11 2
3 3 3 2
7 11 13 1 9 1 9 2
9 11 11 11 2 11 12 2 12 11
14 2 15 13 3 10 9 1 11 11 1 9 1 11 2
40 15 4 3 4 13 9 1 9 7 9 2 16 10 0 3 13 9 1 14 4 13 3 1 0 9 1 9 1 10 0 9 2 15 3 13 9 1 0 9 2
43 2 15 13 3 3 10 9 2 7 15 4 13 3 1 10 0 9 2 2 13 11 11 11 2 15 13 0 9 1 14 13 9 1 10 9 2 15 3 3 4 13 1 2
12 15 13 3 1 15 13 14 13 3 1 11 2
19 11 11 11 2 13 9 2 13 1 9 3 1 10 0 2 0 9 2 2
24 3 1 9 13 11 10 9 2 16 15 1 9 12 9 3 13 1 10 0 9 1 8 9 2
25 15 13 2 16 15 3 4 0 9 2 1 15 13 3 1 2 7 15 13 1 0 9 10 9 2
12 15 4 9 2 15 13 1 10 0 0 9 2
3 11 2 11
8 7 15 4 3 3 3 3 2
12 9 1 11 13 1 0 9 10 0 9 12 2
29 16 11 9 11 11 4 9 9 13 15 1 0 9 2 7 13 15 1 9 2 15 13 3 1 7 13 1 15 2
12 15 4 12 9 2 0 1 0 9 7 0 2
14 3 13 15 3 1 0 7 4 3 3 3 13 0 2
28 15 13 3 14 13 15 1 2 3 10 9 7 9 4 13 3 1 9 2 7 3 15 13 15 3 1 15 2
30 2 15 4 9 13 2 7 3 13 9 3 1 0 9 1 0 9 9 1 3 9 7 11 2 2 13 11 11 11 2
21 15 13 3 3 2 16 15 3 3 4 0 14 13 0 7 0 1 10 0 9 2
21 15 1 9 0 9 1 9 9 4 9 2 8 11 11 1 9 11 11 2 11 2
5 0 9 7 0 9
26 10 3 13 9 11 4 3 13 2 16 1 12 8 4 13 3 1 10 3 13 9 3 1 10 9 2
18 4 15 13 9 1 14 13 2 4 15 13 3 2 1 15 4 3 2
16 15 13 2 15 13 10 9 2 7 10 9 4 13 3 13 2
18 10 0 9 13 10 0 9 1 10 0 9 2 15 11 11 4 13 2
11 9 1 13 3 0 9 13 3 1 9 2
12 3 4 15 13 9 1 14 13 9 1 9 2
21 0 9 1 10 9 2 15 4 13 1 5 12 2 4 3 13 1 9 1 9 12
2 9 3
12 11 11 4 13 10 0 0 9 3 1 3 2
12 11 13 9 2 7 9 13 3 3 1 9 2
2 0 9
15 10 12 9 4 0 1 0 7 0 2 16 9 4 13 2
17 10 12 9 13 3 1 9 12 3 13 2 11 11 8 8 8 2
15 15 4 13 1 11 2 16 15 13 3 1 12 1 9 2
9 10 9 2 15 15 3 3 13 2
13 2 7 1 9 4 10 0 9 1 3 0 9 2
21 2 15 13 1 9 2 2 13 15 15 7 13 3 1 9 1 14 13 1 15 2
35 15 4 3 0 2 16 15 1 9 1 15 1 2 11 2 1 9 3 4 13 15 10 0 9 1 14 13 10 2 0 2 1 10 9 2
15 15 4 15 2 16 11 3 13 11 1 10 0 0 9 2
23 3 4 10 9 11 11 2 15 13 1 10 9 1 11 2 13 9 1 9 1 12 9 2
11 3 3 3 1 9 13 11 2 12 9 2
13 7 11 13 3 1 9 2 4 15 0 1 2 2
8 2 15 4 13 1 0 9 2
8 2 6 2 0 10 9 2 2
16 3 3 0 13 9 11 11 1 0 9 3 0 9 1 9 2
1 9
18 1 9 13 1 9 4 9 13 3 1 11 2 1 11 9 1 11 2
8 3 9 7 15 13 15 3 2
22 3 13 3 15 2 15 4 13 1 14 13 2 6 10 9 4 13 1 0 9 2 2
14 13 10 9 2 15 13 9 1 2 2 13 9 9 2
29 15 4 0 2 15 9 15 4 13 3 1 2 7 3 9 13 9 2 16 15 13 14 13 3 1 10 10 9 2
33 11 9 11 11 13 3 1 9 1 11 7 11 1 14 13 10 9 1 14 13 1 14 13 9 1 11 1 9 2 13 11 9 2
6 2 0 2 13 15 2
14 3 13 15 9 1 10 0 9 1 9 0 0 9 2
8 2 13 15 15 2 13 15 2
18 11 11 13 10 9 1 10 9 2 0 0 9 13 15 1 10 9 2
13 15 4 3 0 1 10 9 2 15 13 14 13 2
11 11 2 2 15 4 3 0 7 0 2 2
10 1 9 11 4 10 0 9 13 0 2
19 1 9 1 9 4 10 13 9 13 1 12 9 2 10 9 1 12 9 2
5 13 9 1 0 9
13 15 13 3 3 1 14 13 10 9 1 9 9 2
14 13 15 3 10 13 9 2 13 15 3 1 10 9 2
7 15 13 3 1 10 9 2
9 15 4 10 0 9 1 9 9 2
34 10 9 4 13 2 16 10 12 0 0 9 4 13 10 0 9 1 9 2 9 9 2 2 7 3 4 3 13 0 9 1 0 9 2
17 11 11 4 9 2 7 1 10 9 13 15 1 9 1 9 11 2
18 2 9 1 9 4 13 2 7 9 4 13 10 0 9 1 9 8 2
8 2 4 15 13 15 2 9 2
14 3 13 10 9 2 15 13 10 9 1 10 0 2 2
24 10 0 9 2 11 11 9 2 4 13 14 13 1 9 1 9 3 1 14 13 15 3 3 2
24 3 4 15 15 1 9 0 9 2 15 13 16 9 11 11 13 10 9 1 10 0 9 9 2
8 15 13 15 13 1 10 9 2
26 15 4 15 13 15 3 1 9 1 10 0 9 7 13 11 11 13 10 0 9 13 1 8 7 9 2
7 1 3 4 9 4 12 2
30 3 13 15 15 3 1 14 13 10 9 1 9 2 7 3 13 15 3 9 1 14 13 9 7 4 0 1 9 12 2
11 15 13 1 9 3 2 2 13 10 0 2
25 12 0 9 1 10 0 1 12 9 13 15 9 2 16 9 4 13 3 1 9 2 11 11 9 2
6 15 13 3 1 9 2
7 2 11 13 10 0 9 2
10 10 9 1 10 9 13 9 9 3 2
16 1 0 9 13 15 1 10 9 14 13 9 1 10 0 9 2
13 4 15 3 0 2 16 15 4 13 7 13 9 2
9 9 1 9 13 9 1 10 9 2
48 2 15 4 13 0 9 3 2 7 1 0 9 13 15 2 16 15 13 0 9 2 1 15 1 9 13 1 9 2 2 13 11 11 2 15 4 13 1 14 13 10 9 1 11 7 13 9 2
9 2 9 2 15 4 0 3 9 2
8 3 3 13 0 2 7 0 2
15 2 7 11 13 3 10 0 9 2 2 13 11 11 11 2
35 2 15 4 13 2 16 1 14 13 10 0 9 1 10 0 9 2 4 9 13 3 2 2 13 11 9 0 9 7 13 9 2 11 11 2
26 15 13 3 1 10 0 9 1 9 1 10 0 9 11 7 11 2 0 1 12 9 1 10 0 9 2
3 15 9 2
29 16 9 13 1 9 2 4 15 3 4 13 2 16 9 13 9 1 0 9 3 2 16 9 3 13 1 10 9 2
37 15 9 2 15 13 2 4 13 0 9 2 15 16 15 4 10 3 0 9 2 15 3 4 4 13 1 9 2 7 15 4 9 0 9 7 9 2
12 1 12 9 4 3 13 8 7 9 1 11 2
25 3 11 2 9 1 0 9 2 13 9 9 1 10 0 9 1 9 1 0 9 0 9 1 11 2
14 2 0 2 15 13 9 12 1 9 10 0 9 2 2
11 9 13 1 10 9 1 0 0 9 3 2
5 10 0 13 11 2
22 1 9 13 10 0 3 10 9 1 12 2 16 9 4 4 0 1 9 1 0 9 2
16 9 13 15 1 9 1 0 1 10 12 9 1 11 9 9 2
9 3 13 12 9 3 10 0 11 2
27 15 4 1 10 9 1 0 9 4 13 2 16 2 15 1 4 9 1 9 3 4 15 15 1 9 2 2
1 9
15 9 4 3 1 9 13 1 11 2 11 9 7 11 9 2
37 7 1 15 2 15 1 10 9 0 9 1 9 0 9 13 10 9 1 10 9 0 9 2 7 1 3 13 15 2 13 2 1 3 3 13 9 2
28 9 9 13 12 9 1 9 2 13 1 9 1 9 1 9 2 12 9 1 9 2 0 13 1 9 1 12 2
29 15 4 9 2 15 13 3 1 9 1 11 2 7 1 13 2 16 9 3 4 13 10 9 7 10 9 1 9 2
7 15 4 3 3 4 0 2
32 15 13 3 2 16 10 0 9 4 4 13 1 10 9 9 9 1 9 2 3 1 9 1 0 9 1 9 1 10 0 9 2
24 10 9 4 13 1 9 1 3 10 0 9 7 1 9 11 11 2 15 4 13 1 10 9 2
19 15 13 10 0 9 1 10 0 9 2 7 9 13 15 3 1 10 9 2
23 15 2 15 13 2 13 8 2 8 2 8 2 11 11 2 3 3 13 2 7 3 8 2
12 11 13 10 0 9 3 7 13 9 1 9 2
22 9 13 1 9 2 3 0 11 11 2 11 11 2 11 11 7 11 11 13 1 11 2
12 15 4 3 3 3 2 15 15 13 14 13 2
5 9 9 4 0 2
2 3 0
5 9 13 1 9 2
13 9 4 4 0 7 0 1 9 3 3 0 9 2
28 15 4 9 1 11 9 2 15 1 9 2 1 10 1 9 0 9 2 13 10 9 2 15 4 13 9 9 2
10 7 13 2 2 15 4 0 9 2 2
40 3 4 15 12 9 1 11 11 2 15 3 13 1 10 3 10 9 1 9 1 10 0 2 3 0 2 0 7 3 0 9 2 15 9 13 2 2 13 15 2
27 3 1 9 13 15 10 13 2 0 2 9 13 1 12 9 1 11 2 3 4 10 0 9 9 1 11 2
2 0 9
14 7 3 4 15 3 3 3 13 9 3 1 10 0 2
10 9 13 3 1 10 13 9 1 9 2
6 15 4 4 4 9 2
16 7 16 15 13 15 2 4 15 13 3 7 13 15 13 3 2
3 7 3 2
16 0 2 10 9 4 0 2 7 15 4 3 3 13 1 9 2
8 15 13 10 9 9 1 9 2
20 2 15 13 3 3 3 2 3 0 9 13 1 0 9 2 2 13 11 11 2
15 15 13 3 1 9 2 16 9 13 15 0 14 13 9 2
28 1 13 9 7 9 4 1 9 9 7 9 1 10 0 9 9 1 0 9 3 13 11 9 1 11 0 9 2
29 9 4 3 1 9 12 13 3 1 9 2 10 9 2 3 3 4 13 1 12 2 7 3 4 9 4 3 0 2
9 0 9 13 15 3 1 0 9 2
29 9 13 3 1 9 1 10 0 9 1 3 1 9 2 9 2 9 7 9 2 1 8 11 11 1 9 1 9 2
39 2 15 4 11 2 15 13 15 1 9 1 9 2 7 15 13 3 1 9 2 16 11 13 9 4 10 0 9 2 15 3 4 13 2 2 13 11 11 2
30 1 9 13 11 11 15 1 10 0 9 1 1 9 14 13 9 7 0 9 1 9 1 3 7 3 0 9 9 1 2
13 1 9 13 15 3 2 16 9 4 13 3 3 2
16 7 1 10 13 9 13 8 9 3 9 1 9 7 0 9 2
8 8 7 9 4 15 3 13 2
23 7 15 13 1 14 13 2 4 9 13 9 7 13 10 0 9 1 9 2 4 9 13 2
16 11 13 15 13 2 15 4 10 0 9 2 7 11 13 9 2
14 1 9 1 2 16 15 13 3 9 1 14 13 9 2
6 11 2 15 4 3 2
12 2 13 15 3 1 10 9 2 13 15 3 2
20 15 13 10 9 1 10 9 2 15 1 9 1 9 13 10 9 0 1 9 2
33 15 4 9 2 16 15 0 9 13 9 1 9 2 7 3 13 2 16 2 1 9 2 4 13 10 15 1 3 9 3 1 9 2
20 15 13 3 3 2 15 15 13 3 1 9 2 16 15 13 3 1 9 3 2
8 13 9 5 12 9 5 5 13
15 16 15 4 10 0 9 3 2 4 15 3 13 15 3 2
8 3 13 15 10 0 9 9 2
1 13
53 11 13 15 15 3 16 15 13 9 2 3 11 3 13 1 2 9 11 2 7 13 1 9 2 7 13 1 10 13 9 1 11 3 13 9 1 10 0 11 2 13 3 3 0 14 13 1 1 2 11 11 2 2
10 3 0 2 13 11 2 7 3 0 2
25 10 0 9 1 9 4 3 13 8 7 13 1 10 9 1 9 1 9 8 11 1 10 0 9 2
27 9 11 11 4 3 1 10 9 13 15 9 1 11 2 7 10 9 1 9 11 11 4 13 1 9 9 2
38 7 9 2 3 8 1 0 9 1 12 9 2 4 3 0 2 13 9 11 11 2 11 11 7 11 11 2 15 12 0 9 1 11 13 1 9 9 2
18 2 6 2 3 15 13 15 1 10 0 9 2 2 13 15 1 11 2
16 7 3 13 15 3 8 13 2 15 3 3 13 1 10 9 2
42 2 15 13 10 3 0 9 3 1 10 9 2 15 15 4 3 1 14 13 2 2 13 15 7 13 1 15 1 9 7 9 2 1 3 9 2 9 2 9 7 9 2
1 9
12 10 9 1 9 1 11 11 2 3 1 11 2
25 9 4 1 9 9 9 2 16 15 4 3 13 15 10 9 7 12 1 14 2 13 1 2 9 2
20 10 0 9 4 3 13 10 0 9 1 3 0 2 15 11 11 4 13 1 2
3 9 7 9
33 9 7 9 4 13 15 3 2 7 3 4 15 3 7 0 13 15 1 14 13 14 13 0 9 2 16 15 13 1 10 0 9 2
14 1 9 1 9 1 9 13 3 9 1 10 0 9 2
15 16 10 13 9 7 0 1 0 9 13 14 13 7 13 2
22 9 13 1 0 10 9 10 0 2 0 9 1 9 2 15 11 13 1 11 11 9 2
2 13 9
54 2 16 15 4 0 13 15 1 14 4 9 1 9 7 9 2 7 15 4 13 1 9 1 0 9 2 2 13 11 2 15 1 9 13 11 2 11 11 2 1 11 2 3 15 3 4 13 1 9 2 9 7 9 2
12 2 15 4 13 15 3 9 9 2 13 11 2
4 13 9 5 12
6 15 4 13 0 9 2
14 2 7 15 13 3 0 9 1 9 2 15 4 13 2
15 7 13 1 2 16 15 3 13 0 2 1 15 4 13 2
21 3 4 11 2 3 13 2 2 15 15 13 2 1 14 13 10 9 1 0 9 2
18 15 4 0 2 13 11 11 2 15 13 9 1 9 2 0 9 2 2
16 9 2 3 15 1 0 9 13 0 1 12 9 9 1 9 2
11 15 13 15 1 3 9 9 1 1 12 2
9 0 15 2 15 4 13 9 1 2
17 10 0 0 9 13 1 9 1 13 9 1 0 9 9 1 9 2
14 15 4 3 0 7 13 2 7 6 3 15 4 13 2
20 1 11 4 15 13 10 0 9 2 15 13 3 0 9 13 10 9 1 9 2
19 2 15 13 10 7 10 9 1 9 1 9 1 15 3 3 4 13 13 2
23 9 13 2 9 13 9 9 1 9 3 3 3 3 1 9 7 3 3 1 9 1 9 2
19 1 0 9 4 15 10 2 9 2 2 10 9 3 13 14 13 1 9 2
13 12 13 9 4 13 10 12 9 1 9 1 9 2
7 7 15 13 15 3 0 2
10 9 13 9 7 13 9 1 0 9 2
15 15 4 3 3 13 0 9 1 11 1 14 13 10 9 2
15 1 2 0 2 9 13 0 9 3 1 0 2 11 2 2
20 11 4 13 9 7 9 2 12 9 1 9 2 7 1 9 13 10 0 3 2
11 15 4 3 13 7 13 0 7 0 9 2
12 15 4 10 9 3 0 7 0 1 10 9 2
16 2 11 2 13 15 2 7 2 15 0 2 15 13 3 16 2
16 9 4 2 3 2 16 15 3 13 1 0 9 1 1 9 2
7 10 9 4 3 13 9 2
8 9 4 13 1 10 0 9 2
12 1 10 7 10 9 4 15 3 4 13 3 2
12 1 0 9 13 15 14 13 9 9 1 9 2
8 11 11 11 4 9 1 11 2
11 2 3 4 15 13 10 0 9 1 9 2
16 16 15 3 4 13 15 2 7 16 9 4 13 15 3 0 2
53 1 10 0 12 9 4 15 3 13 7 13 0 9 1 2 3 3 1 9 2 7 2 3 7 13 2 7 10 0 9 2 9 0 9 2 2 2 0 7 0 2 7 10 0 2 16 10 9 11 4 0 2 2
26 16 15 4 12 9 13 15 1 15 1 10 10 9 1 9 1 9 2 7 15 13 15 1 10 9 2
7 2 15 13 3 1 9 2
13 15 13 15 2 7 15 13 2 3 15 4 0 2
5 3 13 10 9 2
6 15 13 3 3 3 2
26 3 0 2 15 9 13 2 4 9 3 3 1 2 7 3 1 0 9 13 9 3 12 1 9 9 2
17 10 0 9 13 1 9 1 10 0 9 1 11 2 11 7 11 2
23 15 13 13 2 16 9 13 0 9 1 9 1 13 9 2 15 3 13 15 13 1 9 2
22 1 9 1 11 13 3 3 9 2 0 2 3 1 9 3 4 13 15 1 10 9 2
20 7 13 16 15 2 15 13 9 2 4 13 9 1 12 9 1 9 1 9 2
12 9 2 3 15 1 0 9 4 13 1 9 2
21 3 13 15 9 1 10 9 1 9 1 11 2 3 15 13 9 1 9 9 12 2
17 10 0 9 1 9 11 4 15 1 9 1 10 0 9 11 11 2
4 9 1 9 2
17 1 0 9 4 10 9 13 10 9 2 15 13 9 7 0 9 2
30 7 3 3 0 13 9 1 9 1 2 16 9 9 4 13 1 9 1 15 1 11 12 9 2 11 2 11 7 11 2
24 11 9 13 1 10 9 9 3 9 2 15 4 13 2 3 0 9 1 10 9 1 12 9 2
32 7 15 4 3 3 0 3 1 1 10 0 9 2 15 1 9 4 13 9 2 16 9 13 13 9 1 10 0 16 0 9 2
29 15 13 9 1 11 11 7 13 1 10 9 1 9 11 11 1 0 9 2 3 15 13 2 16 9 4 13 3 2
11 3 3 2 16 15 4 10 9 1 9 2
16 15 13 2 16 11 11 13 0 9 1 14 13 9 1 9 2
5 9 0 12 9 12
3 9 12 2
27 3 13 3 0 9 1 14 4 13 1 10 0 0 9 2 7 10 0 9 4 1 3 3 3 0 0 2
6 11 9 13 1 9 2
10 15 4 3 13 2 16 9 4 0 2
30 0 9 13 1 2 3 15 8 13 9 1 9 1 10 0 9 2 9 1 9 2 9 1 9 7 9 1 9 3 2
9 0 1 15 4 10 9 1 9 2
26 10 0 7 0 0 9 4 3 0 1 9 2 15 4 13 1 9 1 0 9 2 9 7 13 9 2
6 0 13 0 1 0 2
19 2 7 15 4 3 3 13 1 15 2 16 15 13 2 15 4 15 15 2
36 2 13 15 13 10 9 2 2 13 15 1 9 1 10 9 2 7 10 3 0 9 2 13 3 2 2 4 15 3 3 3 13 10 9 2 2
29 1 10 13 9 4 15 3 0 2 16 10 9 4 0 2 16 10 9 4 2 13 2 10 9 1 14 13 9 2
21 9 13 1 9 2 15 3 13 10 3 12 9 2 1 12 12 12 5 1 9 2
15 7 15 4 3 3 11 9 1 9 2 15 4 13 9 2
13 10 0 1 10 0 9 4 13 1 3 0 9 2
27 2 13 15 1 15 2 16 15 3 3 13 15 1 14 13 10 10 9 2 3 4 9 2 2 13 15 2
