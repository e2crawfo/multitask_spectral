288 17
13 3 1 15 3 2 13 2 3 13 9 1 11 2
25 2 15 2 11 7 11 2 13 13 10 9 1 9 7 15 13 15 1 13 16 13 0 7 0 2
20 13 16 15 13 10 9 1 10 9 2 3 1 10 9 2 16 13 13 2 2
52 3 10 11 2 3 13 10 9 3 7 13 16 1 11 13 1 10 10 9 10 9 13 1 13 16 15 13 7 3 13 10 9 16 13 10 9 0 1 11 2 13 2 3 12 1 10 9 1 2 11 2 2
9 2 13 1 10 9 1 9 2 2
20 11 13 9 1 10 9 2 3 11 15 3 15 13 1 10 9 1 9 0 2
28 10 9 1 11 13 13 3 1 9 13 13 10 9 0 1 10 10 9 0 2 13 13 10 9 1 10 9 2
55 10 9 1 10 9 13 1 15 1 10 9 13 1 10 9 1 10 11 2 13 1 13 2 13 13 2 1 9 10 0 1 10 9 2 1 3 2 1 15 13 2 13 11 1 15 13 9 7 13 10 9 1 10 9 2
55 1 10 9 13 1 10 9 1 10 9 2 1 12 9 2 15 13 3 9 2 13 13 10 9 13 12 9 3 1 10 9 1 10 9 2 13 1 10 9 2 10 9 1 9 1 9 2 10 9 7 10 9 1 9 2
36 1 13 9 1 10 9 13 13 1 10 9 1 9 0 1 10 11 7 3 1 10 9 1 11 2 3 13 10 9 2 10 9 0 13 13 2
62 13 10 9 1 10 10 9 2 3 13 2 1 9 2 1 10 9 1 10 2 9 2 2 15 13 3 13 10 9 1 9 2 1 9 13 1 13 2 3 2 9 2 2 3 1 9 3 0 7 1 9 1 13 2 13 1 9 1 2 9 2 2
29 13 15 1 10 2 11 2 2 13 1 10 9 0 2 7 13 15 1 9 1 10 9 1 0 2 0 7 13 2
26 10 9 13 13 10 9 1 2 9 2 2 12 9 1 9 2 13 1 10 9 1 2 9 2 3 2
11 13 1 13 3 10 10 9 1 9 13 2
54 11 13 2 1 10 9 2 3 2 10 9 1 10 11 2 15 13 1 12 9 1 10 11 2 1 10 13 2 9 1 9 2 1 10 9 1 11 7 11 7 1 10 9 0 15 1 15 13 2 7 3 2 13 2
36 11 2 9 1 10 9 2 13 1 10 9 1 13 10 9 0 2 13 10 15 15 13 2 0 2 13 1 10 9 1 15 3 1 10 11 2
9 13 1 13 16 13 1 13 0 2
25 11 13 2 3 2 10 9 2 3 0 1 10 10 0 9 2 1 13 1 15 13 10 9 0 2
29 13 1 15 15 13 10 9 1 16 15 15 13 2 15 13 1 10 9 3 0 2 16 3 1 10 0 9 0 2
13 12 9 15 2 1 9 2 13 3 1 10 9 2
6 9 1 10 9 0 9
3 11 13 9
30 10 11 2 12 1 10 0 9 0 1 10 9 0 2 13 10 9 7 13 9 1 10 9 0 7 1 10 9 0 2
16 10 11 13 15 10 9 7 10 9 1 10 12 9 13 13 2
17 10 9 3 13 9 2 7 10 9 13 1 10 9 1 10 9 2
75 13 1 13 3 9 13 1 10 9 1 9 1 9 2 10 11 13 13 10 10 9 1 9 7 9 1 9 1 10 9 2 9 10 1 10 9 1 9 0 1 10 9 1 9 2 0 1 9 3 0 0 1 10 9 1 2 9 2 7 2 9 2 1 15 10 9 1 9 13 7 13 1 13 9 2
42 10 9 13 10 9 7 9 9 2 10 12 9 1 15 1 10 9 1 10 9 2 2 1 15 10 10 9 1 10 0 9 13 13 7 13 10 9 1 10 10 9 2
34 1 10 9 1 9 7 9 13 2 3 2 9 10 11 2 9 1 9 3 13 1 10 9 0 1 9 7 3 1 10 10 9 12 2
15 10 11 13 3 2 1 11 2 10 0 9 1 10 11 2
23 10 0 9 13 13 1 11 2 1 10 9 11 2 9 2 2 11 7 11 2 9 2 2
8 1 10 11 2 1 10 9 2
21 9 1 10 11 2 11 2 1 10 9 1 10 9 1 10 9 13 1 10 11 2
35 10 9 1 10 11 2 11 2 1 12 9 2 13 1 9 12 9 2 12 9 1 10 2 12 1 15 2 1 13 13 9 1 10 9 2
31 10 9 1 11 2 9 1 10 11 2 13 10 9 1 10 9 2 11 2 1 13 9 0 1 10 9 10 1 12 9 2
6 10 9 13 10 9 2
10 10 9 13 10 9 1 9 1 9 2
11 10 9 2 3 2 13 10 9 1 11 2
1 11
41 2 13 0 16 10 9 2 1 10 9 1 10 11 2 13 3 13 7 16 13 13 10 9 0 7 0 1 10 9 0 1 10 9 1 16 15 13 10 9 0 2
35 7 3 15 13 10 9 0 1 10 9 2 16 13 2 3 2 1 10 9 0 1 10 9 1 10 9 0 7 13 15 13 10 11 2 2
53 13 9 1 10 9 1 10 11 2 11 2 1 10 9 1 10 9 12 1 10 9 1 10 11 2 3 13 1 10 9 1 10 2 0 9 1 10 9 0 1 10 9 1 10 11 2 2 1 3 13 10 9 2
6 9 0 2 9 12 2
17 10 9 0 1 9 0 7 2 7 13 2 1 10 9 1 9 2
23 9 0 7 0 1 10 9 1 10 9 0 1 10 9 2 13 1 10 9 7 10 9 2
22 9 15 13 3 2 1 10 9 0 7 3 13 7 1 10 9 0 2 11 2 0 2
2 11 2
16 1 9 1 9 2 1 10 9 2 9 7 9 1 10 9 2
71 13 12 9 1 10 9 1 12 2 10 9 1 10 11 2 11 2 13 13 3 1 1 10 0 9 12 2 1 10 9 1 10 9 15 13 13 3 7 3 1 10 9 1 11 15 3 13 9 1 10 9 1 10 11 2 3 1 10 9 1 10 9 0 2 13 16 13 10 9 0 2
52 7 3 3 3 3 2 3 1 10 11 2 11 2 10 9 0 13 2 1 10 9 0 1 13 10 11 2 11 2 15 13 0 9 1 9 0 15 13 1 9 2 3 1 11 3 1 10 9 1 10 9 2
18 10 11 3 13 13 10 9 13 1 10 10 9 1 10 9 1 12 2
36 1 10 9 1 10 0 9 1 10 9 13 2 10 9 13 13 10 9 1 9 1 12 9 1 9 2 7 13 1 3 13 1 10 12 9 2
28 3 1 9 0 2 10 9 13 1 10 9 0 1 12 9 1 9 2 7 15 1 10 9 13 10 12 9 2
41 1 10 9 1 10 9 2 15 13 2 10 11 3 13 7 10 0 12 9 1 15 10 11 13 1 10 9 2 10 9 13 15 1 10 9 1 12 9 1 9 2
20 10 9 13 10 9 1 12 9 1 10 12 9 1 9 1 9 0 1 12 2
23 10 9 13 13 1 12 9 1 9 1 12 2 10 12 9 1 9 16 1 10 9 0 2
82 1 10 9 0 2 10 9 1 10 9 1 10 9 13 15 2 3 2 1 10 2 9 1 10 9 1 0 9 13 1 9 1 10 0 9 1 9 2 9 1 10 9 1 9 2 2 7 1 9 1 10 9 1 9 1 9 3 13 1 10 0 9 1 9 0 2 1 3 13 1 9 0 2 9 1 10 0 7 0 11 2 2
43 10 11 0 2 11 2 13 3 10 9 1 10 0 11 2 1 10 9 13 0 10 9 1 10 9 2 11 2 3 13 1 10 9 1 9 2 2 13 10 9 1 11 2
24 10 9 13 3 16 11 13 12 1 10 10 3 0 9 2 10 9 11 7 10 9 2 11 2
38 11 2 10 0 13 1 10 11 2 13 10 9 1 13 10 11 7 1 13 10 10 9 0 2 1 10 9 13 1 10 9 1 10 9 1 10 9 2
6 11 1 10 9 1 9
42 10 0 9 1 9 1 10 9 1 11 13 13 9 1 10 9 12 1 9 1 11 2 13 3 10 9 0 1 10 11 7 10 9 0 1 11 2 9 1 10 9 2
19 1 9 13 2 10 12 9 13 9 1 16 10 9 0 13 3 1 11 2
27 1 10 11 2 10 9 1 10 11 3 15 13 1 10 9 0 2 3 13 13 10 9 10 9 1 11 2
4 9 1 10 11
79 2 13 2 1 10 9 1 10 11 3 13 1 10 9 13 1 10 9 7 1 10 9 2 1 10 9 1 9 13 2 10 9 0 13 15 1 13 13 2 1 10 9 1 2 13 1 9 2 2 13 10 9 2 3 3 2 3 13 10 9 2 3 3 1 10 12 9 2 13 1 4 2 13 2 1 10 9 2 2
18 13 1 10 9 0 2 3 13 13 1 15 13 3 3 1 10 9 2
30 3 3 1 11 2 10 9 0 1 11 2 15 13 11 1 9 1 13 1 9 10 10 9 1 0 9 1 10 11 2
33 13 3 9 1 10 9 2 10 9 13 10 9 1 2 11 2 2 11 13 13 10 11 1 13 15 1 10 9 1 10 9 0 2
17 7 9 13 2 3 2 12 9 0 1 13 10 9 0 1 9 2
22 10 9 1 11 13 9 7 10 9 1 2 11 2 13 10 9 2 1 9 3 0 2
18 1 10 11 2 13 3 12 0 0 2 11 2 1 10 9 2 11 2
1 11
4 10 9 1 11
56 10 9 11 2 11 2 13 3 10 9 1 10 9 0 2 1 15 13 10 11 1 9 2 0 9 1 10 11 1 10 9 2 13 1 10 11 2 3 10 9 13 3 1 11 2 11 2 2 15 3 13 1 10 0 9 2
19 10 11 13 1 13 10 0 1 10 9 2 1 11 1 13 10 0 9 2
1 11
15 1 10 9 1 11 10 9 1 10 9 0 2 3 13 2
19 12 9 2 0 1 12 7 0 1 12 2 13 9 3 13 7 13 9 2
22 10 9 1 10 9 1 0 9 0 13 3 1 11 2 1 10 11 2 10 0 9 2
21 13 1 9 7 9 2 13 13 1 10 9 3 13 1 13 10 9 1 10 9 2
45 11 10 9 15 15 13 1 10 9 1 10 9 3 10 9 1 10 9 13 16 15 15 13 1 10 9 15 13 10 9 2 15 15 13 3 15 13 16 15 13 1 10 9 0 2
22 10 11 13 13 0 9 1 10 9 1 10 9 13 1 9 3 7 1 10 9 3 2
41 13 15 2 1 9 2 10 9 2 11 2 2 11 1 10 13 9 12 2 2 11 2 2 12 2 2 11 2 2 12 2 2 11 2 2 12 2 9 2 12 2
9 10 9 1 9 13 10 10 9 2
19 1 10 9 2 13 15 10 9 3 1 10 9 1 10 9 1 10 9 2
54 1 13 15 10 9 1 11 2 3 10 9 1 9 1 10 9 2 3 13 1 0 9 2 13 1 4 13 1 15 1 9 2 3 10 9 15 3 13 9 1 9 2 16 13 1 10 9 2 3 13 1 10 9 2
30 2 3 13 15 10 9 16 15 13 1 10 9 1 10 9 7 3 3 1 10 9 1 15 3 13 2 2 13 11 2
16 12 9 1 10 9 1 10 9 13 1 10 11 2 1 11 2
17 10 0 12 9 13 9 0 2 13 1 10 9 1 10 9 13 2
17 7 3 3 13 9 3 0 2 16 10 9 3 13 13 1 15 2
8 10 9 0 13 1 10 11 2
18 12 9 13 1 11 2 12 9 1 10 11 7 12 12 1 10 11 2
21 1 10 11 2 11 2 11 7 11 2 10 9 13 1 12 12 7 12 12 9 2
16 10 11 13 12 9 2 10 11 12 9 7 10 11 12 12 2
3 13 11 2
41 2 10 0 9 1 10 9 11 7 11 13 9 1 10 9 0 7 9 15 13 1 10 9 1 13 9 1 9 3 0 2 3 13 1 10 9 0 10 9 2 2
14 10 9 1 10 9 3 3 13 10 9 1 10 9 2
40 3 2 13 16 10 9 1 10 9 13 1 10 11 1 9 1 13 10 9 0 1 10 9 2 3 9 2 1 10 9 0 2 13 1 13 10 10 9 2 2
37 7 16 15 13 1 10 9 3 15 13 2 3 1 12 1 10 9 1 10 9 2 10 9 3 13 10 9 1 2 9 2 1 10 9 1 11 2
33 2 11 2 2 10 9 1 9 13 1 10 9 2 3 9 1 9 13 10 9 1 10 9 1 10 9 1 10 9 1 10 9 2
42 11 13 10 9 2 15 3 15 13 1 10 9 1 9 2 9 1 9 2 7 15 13 1 10 10 0 9 1 9 1 10 9 2 3 3 2 1 12 1 10 9 2
19 11 13 10 0 9 9 1 9 2 1 10 15 13 9 1 10 10 9 2
27 13 10 0 9 15 13 10 9 1 10 9 2 15 13 13 1 13 15 7 13 1 10 9 1 10 9 2
42 13 3 4 9 1 10 9 1 10 9 13 7 10 9 1 10 9 2 7 4 10 9 1 10 9 0 2 13 1 10 10 9 2 15 3 13 13 2 9 2 9 2
18 11 7 11 2 3 2 13 15 9 15 13 1 9 3 0 10 9 2
9 10 0 13 10 9 1 10 9 2
21 7 10 9 13 15 10 10 9 1 10 9 15 13 2 1 10 9 15 15 13 2
15 10 0 2 1 10 9 2 13 10 10 9 2 11 2 2
34 7 2 1 10 9 1 9 2 13 12 9 1 9 1 10 9 2 15 15 13 4 2 7 4 1 9 2 1 15 13 1 10 9 2
27 1 10 9 2 10 2 9 2 2 15 13 10 9 1 10 9 2 13 3 13 2 13 1 10 10 9 2
19 9 2 16 13 10 9 2 2 9 2 9 15 13 2 13 13 7 13 2
12 10 9 13 0 2 15 13 13 1 10 9 2
19 2 16 13 10 9 3 1 9 2 1 3 13 1 15 13 0 1 15 2
15 3 2 13 13 10 11 2 3 1 15 2 2 13 11 2
34 10 9 0 1 9 13 10 9 3 1 10 9 2 3 1 13 1 3 12 9 1 10 9 1 10 9 2 13 9 1 10 9 2 2
3 9 13 9
20 10 11 2 9 0 2 13 10 9 0 15 13 1 10 9 0 1 10 9 2
9 10 9 1 11 13 1 12 9 2
11 13 9 1 9 7 1 9 2 9 2 2
8 3 15 13 1 10 12 9 2
14 10 9 11 7 11 13 3 10 9 11 1 10 11 2
25 11 2 11 2 11 7 11 13 9 1 9 15 13 3 1 10 11 10 9 1 11 13 1 11 2
37 10 9 13 10 9 1 10 9 1 10 9 9 2 9 1 10 9 0 7 0 1 10 9 2 1 10 9 1 10 9 7 1 10 9 0 0 2
27 10 11 13 1 10 9 0 1 9 1 10 9 12 2 3 13 10 2 9 2 1 13 10 9 1 9 2
18 10 9 1 9 13 1 9 0 13 1 10 9 1 10 9 1 12 2
11 12 9 3 2 10 9 13 1 13 11 2
11 10 9 13 10 9 1 15 3 13 9 2
19 10 9 11 2 12 2 1 10 9 11 2 13 9 0 2 3 10 9 2
26 2 10 0 13 13 3 10 9 2 13 10 9 7 13 10 9 1 10 9 1 10 9 2 2 13 2
9 11 2 12 2 9 1 10 11 2
15 2 3 13 10 9 1 13 10 9 15 15 3 13 3 2
30 3 13 10 9 1 10 9 1 9 2 13 16 15 13 16 13 10 9 1 9 2 15 13 13 10 9 1 13 3 2
11 10 9 13 10 9 1 15 13 10 9 2
14 10 9 1 10 9 13 13 10 9 1 3 13 9 2
15 10 9 3 10 9 1 11 13 13 9 0 7 13 2 2
7 11 2 12 2 9 0 2
10 2 13 1 10 10 9 1 10 9 2
17 3 13 2 15 13 10 9 3 1 10 0 7 1 10 9 0 2
10 1 10 9 15 3 13 1 15 13 2
13 3 15 3 13 9 13 1 10 9 1 10 9 2
25 15 13 16 13 9 7 3 10 9 2 7 3 2 3 13 15 13 16 3 3 13 3 9 2 2
10 11 2 12 2 13 1 9 2 9 2
16 2 15 13 3 0 2 3 9 2 13 9 3 0 7 0 2
9 10 9 3 13 13 1 10 9 2
20 3 2 10 9 13 1 10 9 0 13 1 10 9 0 2 15 13 0 2 2
6 9 13 12 9 7 9
12 9 2 9 2 9 0 7 9 1 10 9 2
23 15 13 15 1 10 9 15 13 4 13 1 10 9 1 10 11 2 13 3 1 10 9 2
32 10 9 13 13 1 12 9 2 1 10 9 1 13 1 9 1 9 1 9 7 9 13 1 0 9 2 13 1 10 9 0 2
21 10 9 1 10 11 2 11 2 13 16 10 9 13 13 10 9 0 1 10 11 2
17 15 13 16 13 13 10 9 2 7 3 13 10 9 1 10 9 2
22 11 2 10 9 13 13 1 9 1 10 11 1 9 1 9 2 9 7 9 1 9 2
6 10 9 13 13 13 2
12 11 2 1 15 15 3 13 13 3 1 15 2
7 3 13 1 15 15 13 2
6 15 13 3 2 3 2
6 13 9 13 2 13 2
8 1 9 15 13 1 12 9 2
1 9
17 10 9 1 10 11 13 13 10 9 1 13 9 1 13 10 9 2
23 10 0 9 13 1 9 2 10 12 9 2 7 10 0 9 2 1 9 2 15 12 2 2
15 10 9 15 3 13 13 9 1 10 11 1 11 12 9 2
14 10 9 0 1 9 1 10 9 13 1 10 9 13 2
9 1 12 0 2 10 11 13 12 2
28 10 9 1 11 13 13 10 9 1 13 10 9 7 13 1 13 10 9 1 10 9 2 13 1 9 12 9 2
1 9
41 1 10 9 1 9 1 10 9 2 11 3 13 10 9 1 9 1 10 9 2 3 1 9 13 2 1 13 10 9 9 1 10 9 2 15 13 4 13 1 9 2
19 10 9 2 11 2 13 16 10 9 1 10 11 2 3 13 10 9 2 2
27 15 13 16 10 9 13 13 1 10 9 12 1 9 2 3 1 9 0 2 1 10 9 12 1 10 9 2
19 10 11 1 9 2 1 10 9 2 2 13 3 15 1 10 0 9 2 2
21 2 3 15 13 9 0 1 10 9 1 10 9 2 1 9 1 9 2 2 13 2
16 1 11 2 13 1 9 10 9 1 13 10 9 1 10 9 2
22 15 13 1 12 9 10 9 0 1 13 10 9 7 9 13 1 10 9 1 12 9 2
32 10 9 1 11 2 11 2 11 2 2 13 16 10 9 15 13 13 1 10 9 2 13 3 2 1 10 9 1 10 9 2 2
40 13 1 11 2 9 1 10 9 1 10 11 1 10 9 1 10 11 2 11 2 7 1 11 2 9 1 10 9 2 11 2 11 13 12 9 0 3 1 11 2
34 1 10 3 12 9 1 10 9 2 13 0 9 3 10 11 2 11 2 11 2 11 7 11 2 9 1 10 11 1 10 9 1 9 2
27 10 11 2 3 2 13 10 9 11 12 7 12 2 0 1 13 1 9 9 7 9 1 9 1 10 9 2
16 13 13 0 9 2 9 2 9 2 13 1 12 9 1 9 2
12 11 7 1 3 15 13 3 0 10 9 10 2
27 13 1 10 9 3 2 15 3 13 15 13 3 0 1 3 13 1 10 9 2 1 10 9 1 10 9 2
3 7 3 2
7 13 15 1 10 10 9 2
6 3 3 15 13 11 2
9 13 16 15 13 10 9 1 9 2
11 11 3 13 10 9 1 10 1 10 9 2
4 13 1 11 2
9 15 10 9 1 9 13 13 3 2
4 9 13 10 9
34 10 9 1 10 9 13 1 10 9 1 10 9 16 13 10 9 2 13 1 10 0 9 1 9 2 15 3 15 13 1 13 10 9 2
21 1 10 9 2 10 9 13 9 1 9 1 0 1 12 1 12 9 1 10 11 2
15 1 10 9 1 12 2 11 13 10 9 1 12 12 11 2
12 1 10 9 3 13 9 1 15 13 4 13 2
18 10 9 0 1 15 1 10 11 1 10 11 13 1 1 9 12 9 2
8 2 10 9 13 13 10 9 2
27 7 3 3 13 9 1 9 2 10 9 1 10 9 1 15 13 10 9 1 10 9 0 1 10 9 0 2
21 3 1 13 1 15 10 2 7 13 1 9 10 9 1 10 9 2 2 13 11 2
21 1 11 2 10 9 1 10 9 11 13 11 2 9 13 1 9 0 1 10 11 2
22 11 13 0 1 11 2 13 1 9 1 12 1 11 2 11 2 1 12 9 1 9 2
9 13 3 9 1 11 7 1 11 2
10 13 13 1 10 9 1 13 10 9 2
20 13 15 2 10 11 2 7 10 9 11 2 11 2 11 2 11 7 10 11 2
7 13 15 7 13 10 9 2
8 15 13 12 9 1 10 9 2
7 12 11 13 1 10 11 2
8 3 15 13 13 1 10 11 2
29 1 10 9 0 1 11 2 12 2 2 3 2 10 9 13 10 9 1 9 0 1 10 9 2 13 1 10 9 2
25 10 9 2 10 9 2 10 9 1 10 9 13 10 9 1 10 9 1 10 0 15 10 9 13 2
24 1 10 9 13 2 10 9 11 13 10 9 1 11 3 9 2 13 16 15 13 1 10 9 2
38 10 9 1 10 11 2 11 2 13 16 2 1 10 0 9 2 10 9 13 2 13 1 10 11 2 15 13 0 2 16 15 13 9 1 10 9 2 2
6 11 13 9 1 10 11
27 11 13 16 10 9 15 13 7 13 9 1 10 11 13 1 9 10 9 1 10 11 16 10 9 13 13 2
9 11 2 15 10 9 1 10 9 2
13 11 2 13 16 11 13 10 10 9 1 10 9 2
6 15 13 1 10 9 2
14 16 15 13 1 15 2 10 9 13 9 2 13 13 2
12 10 9 13 3 2 13 10 9 0 3 9 2
12 13 10 7 0 9 2 9 2 9 7 9 2
16 0 7 0 9 2 11 2 9 0 7 9 13 9 7 9 2
22 1 11 2 10 11 13 10 9 2 10 1 15 9 2 7 9 0 1 13 10 9 2
24 1 15 2 10 9 13 0 1 10 9 1 9 1 10 9 7 10 9 15 13 3 13 0 2
7 10 11 3 13 9 0 2
11 10 9 0 13 13 3 1 13 10 9 2
19 1 10 9 1 10 9 13 9 2 13 16 9 1 10 9 13 10 15 2
26 10 9 1 10 9 2 9 11 2 13 16 10 9 13 10 9 1 13 7 13 10 9 1 10 11 2
25 11 13 16 1 10 9 13 4 13 10 9 1 10 9 1 10 11 1 3 12 9 1 10 9 2
22 10 9 13 13 1 9 1 10 9 13 2 11 2 11 2 2 1 9 1 10 11 2
25 10 9 15 13 1 15 13 7 10 9 13 2 13 1 10 9 1 10 9 2 2 1 13 3 2
10 11 13 13 3 16 10 9 13 13 2
6 9 3 1 10 9 2
10 9 1 9 1 10 9 1 10 9 2
8 9 1 10 9 2 9 12 2
5 1 12 1 9 2
33 9 1 10 9 2 10 9 13 1 10 9 11 2 11 2 11 2 11 2 11 7 11 13 15 10 9 3 13 1 13 10 9 2
29 1 10 11 2 15 13 11 1 11 2 13 13 9 13 1 10 9 12 7 10 9 12 2 3 1 9 7 11 2
14 15 13 3 1 10 9 7 10 9 13 13 1 12 2
19 10 9 11 2 15 13 1 10 9 1 10 9 2 13 10 9 1 9 2
31 15 3 0 13 1 10 9 1 10 11 2 1 10 9 12 7 10 9 12 2 3 1 11 2 1 15 13 1 10 9 2
9 1 12 9 1 10 9 2 9 13
13 10 9 3 13 1 9 1 9 1 10 0 9 2
15 10 9 13 13 2 1 12 9 1 15 13 1 10 11 2
21 10 9 1 16 10 9 1 9 1 10 9 13 15 13 1 12 9 1 10 9 2
18 15 13 3 13 1 10 9 1 12 9 2 3 12 9 3 13 13 2
5 9 13 13 1 9
22 10 9 2 12 1 12 2 1 10 0 9 1 10 11 13 10 9 1 10 9 0 2
13 1 10 9 2 10 9 13 10 9 2 15 13 2
6 2 13 1 13 2 2
34 1 10 9 1 9 11 2 10 9 13 13 10 9 1 16 3 13 13 10 9 16 10 11 3 15 13 1 10 0 9 1 10 9 2
7 9 1 11 3 13 13 9
5 2 13 13 9 2
14 13 9 1 16 16 13 13 1 10 9 2 15 13 2
25 15 13 9 2 2 13 11 2 12 2 10 9 1 10 9 1 10 9 1 11 11 2 11 2 2
7 11 13 16 13 3 9 2
8 2 3 13 13 9 0 2 2
11 10 9 13 13 1 10 9 1 10 9 2
16 10 9 0 13 10 12 9 1 9 15 13 3 1 10 9 2
2 3 13
11 9 13 1 10 9 1 10 9 2 3 2
19 1 10 11 2 12 9 13 1 9 2 10 9 11 7 10 9 0 11 2
21 3 2 10 9 0 11 3 3 13 13 1 10 9 11 2 9 1 10 9 0 2
10 13 1 10 9 10 0 9 0 11 2
25 7 2 3 1 12 9 1 9 2 13 10 10 9 10 9 11 2 9 1 10 9 1 12 9 2
25 1 10 0 9 2 12 9 2 10 11 1 11 13 10 11 2 12 2 1 10 9 1 10 9 2
10 10 11 13 10 9 1 10 0 9 2
15 13 15 10 9 1 10 9 11 1 10 9 1 10 9 2
12 1 10 9 2 13 13 10 10 9 2 11 2
20 1 11 15 13 10 9 11 2 15 13 15 13 1 11 2 3 1 10 11 2
23 10 9 1 10 2 9 2 15 13 1 10 9 1 11 2 15 3 13 1 13 10 9 2
26 10 9 13 4 13 2 1 9 0 2 1 12 9 2 11 2 11 2 9 2 7 11 2 0 2 2
28 2 10 9 13 9 13 1 9 7 9 3 1 10 9 1 9 1 9 2 2 13 11 2 9 1 10 11 2
35 12 10 9 1 10 11 2 11 2 1 10 11 1 10 11 13 3 0 9 10 9 0 1 9 1 10 9 3 9 1 9 1 10 9 2
8 10 9 0 13 1 12 9 2
12 11 13 0 1 9 1 10 9 7 9 11 2
19 1 10 9 1 10 9 2 10 9 13 13 1 13 10 9 1 10 9 2
36 10 9 1 10 9 0 1 10 11 2 1 11 2 11 2 12 2 13 16 13 13 10 9 1 9 1 9 1 9 1 9 1 10 9 11 2
16 10 9 3 13 3 10 9 3 13 13 3 1 10 9 0 2
20 10 9 1 15 12 13 3 11 13 10 9 2 1 10 9 1 10 9 12 2
12 15 13 13 10 9 7 13 10 9 1 11 2
14 2 10 9 15 12 13 13 13 9 1 10 10 9 2
27 15 13 3 3 13 15 13 1 10 9 1 10 10 9 2 2 13 11 2 1 15 11 13 10 0 9 2
7 2 13 10 0 3 13 2
10 1 10 9 13 3 9 12 9 2 2
12 1 10 9 1 11 2 11 15 13 1 12 2
23 1 10 9 2 11 13 13 10 9 0 11 2 1 15 13 1 10 9 0 13 1 11 2
27 10 9 0 11 13 16 2 1 13 10 9 1 10 9 0 2 15 13 10 9 7 13 13 10 9 0 2
15 1 9 1 10 10 9 2 15 13 1 3 1 9 13 2
13 2 15 13 3 15 13 4 13 10 0 9 2 2
21 10 9 15 13 13 10 9 13 2 11 2 1 10 9 0 1 10 9 13 0 2
28 7 13 3 0 1 9 13 15 1 13 10 0 11 1 10 9 1 9 0 0 1 10 9 1 10 9 13 2
