1032 17
32 10 9 9 7 3 3 13 13 10 12 9 0 9 9 2 3 12 2 2 9 7 10 0 0 9 0 10 0 9 13 13 2
25 10 9 10 0 9 13 2 7 10 0 9 7 10 3 0 9 13 3 2 13 15 10 9 9 2
26 9 3 2 16 10 0 9 9 12 0 9 3 13 0 9 15 2 15 10 0 9 15 0 0 13 2
17 2 10 0 9 3 9 0 9 3 0 12 9 13 10 3 2 2
26 15 1 3 10 9 9 0 10 9 2 7 15 9 0 10 0 0 9 9 2 7 10 0 0 9 2
30 10 0 0 9 9 3 10 9 9 0 9 13 2 7 10 0 0 9 2 13 10 0 11 11 2 10 11 11 9 2
15 15 15 13 2 16 10 0 9 10 9 9 10 9 13 2
23 10 9 10 0 9 9 10 10 9 13 3 2 16 10 9 10 10 9 13 10 0 9 2
12 10 9 9 0 13 10 9 2 13 11 11 2
10 10 0 9 3 0 12 9 13 9 2
23 15 0 13 10 9 9 0 0 0 9 7 10 0 0 12 0 9 7 12 0 9 13 2
38 10 9 13 10 10 9 2 16 10 9 9 3 9 9 0 1 12 9 9 13 9 2 7 15 7 2 16 10 9 0 9 0 9 9 10 9 13 2
12 3 13 3 10 0 9 11 0 9 0 9 2
13 10 9 0 9 13 10 9 0 0 2 0 9 2
35 0 9 13 10 9 10 0 7 10 0 11 9 0 9 2 10 0 9 2 10 0 0 9 9 2 7 10 11 11 11 11 11 11 9 2
15 9 1 3 13 3 3 11 0 9 0 9 10 0 9 2
35 10 9 13 2 7 10 0 9 10 0 9 13 10 9 2 15 10 9 13 10 9 2 16 11 0 0 9 1 3 13 13 10 9 9 2
45 10 9 0 0 9 13 10 0 9 2 7 3 10 9 10 9 13 10 9 9 1 2 15 10 9 1 10 9 3 13 3 10 9 10 9 10 0 0 9 7 10 0 0 9 2
19 10 9 15 13 3 2 16 10 9 9 10 9 9 3 9 2 7 9 2
25 10 9 10 9 9 13 2 0 9 13 10 9 1 2 10 0 9 7 3 0 13 10 0 9 2
13 10 9 12 9 10 9 9 1 0 0 9 13 2
9 15 3 0 0 7 0 9 13 2
30 10 9 9 2 16 10 0 7 0 9 15 3 13 2 3 2 16 10 9 0 2 10 9 0 13 2 3 0 9 2
49 0 9 10 0 9 2 10 0 9 9 10 11 11 2 10 0 9 9 9 7 9 10 11 11 2 10 0 0 7 0 9 9 2 10 0 7 10 0 11 9 0 9 2 10 11 0 9 9 2
39 3 9 10 0 0 2 0 2 9 9 2 3 10 9 7 10 9 10 0 7 0 9 0 9 10 9 1 9 2 3 9 2 9 7 9 2 9 13 2
46 10 0 9 0 9 10 9 0 9 10 11 11 9 2 10 11 11 11 11 11 7 10 15 0 0 2 0 9 9 2 10 0 0 9 9 2 10 0 0 9 3 12 0 9 13 2
11 9 1 10 0 9 0 0 9 13 13 2
22 3 10 3 0 0 9 9 13 3 13 7 9 3 13 2 16 11 3 11 1 13 2
32 10 9 1 3 15 3 0 2 16 0 7 0 9 10 9 9 13 9 2 7 3 15 3 13 2 16 10 9 13 10 9 2
29 7 3 10 9 2 9 2 9 2 9 9 7 3 0 9 2 16 10 9 7 3 10 9 2 9 13 10 9 2
18 10 11 11 0 9 1 0 2 16 3 0 0 9 13 10 9 9 2
17 3 0 13 15 0 9 2 16 10 9 3 0 9 13 10 9 2
17 10 0 0 9 2 3 0 10 9 2 10 9 9 0 10 9 2
14 9 9 13 10 9 2 9 13 10 9 2 9 1 2
33 10 0 9 1 15 3 0 13 2 7 15 3 15 3 13 2 15 13 10 9 10 9 2 3 13 10 9 10 9 7 15 13 2
10 3 13 9 0 9 10 0 0 9 2
12 10 9 9 13 10 9 2 7 9 0 9 2
15 10 9 3 12 9 13 2 15 12 13 3 10 0 9 2
21 10 0 9 13 13 2 7 13 10 0 0 9 10 0 9 7 10 10 9 3 2
9 13 9 1 10 0 9 10 9 2
59 10 9 10 11 7 10 11 0 2 10 11 7 10 11 0 7 10 11 11 11 11 2 10 11 11 11 11 11 11 11 11 2 7 10 11 11 11 11 11 11 2 3 10 11 11 11 11 2 10 11 0 7 10 11 0 0 9 13 2
14 10 0 9 12 2 10 0 9 12 9 9 13 9 2
15 10 16 12 9 13 10 9 2 3 10 0 9 9 13 2
26 11 11 2 10 11 0 9 9 1 16 3 0 8 9 9 13 2 3 0 0 13 10 9 10 9 2
14 10 0 9 1 10 11 0 9 10 11 0 13 3 2
26 3 3 0 2 16 10 11 0 9 9 13 3 10 11 0 2 7 10 9 3 0 0 9 13 3 2
8 9 1 0 0 9 7 13 2
17 3 15 2 16 10 11 0 9 0 9 3 13 15 10 11 9 2
10 10 9 3 0 2 0 9 7 13 2
16 10 0 9 13 10 9 9 9 2 10 9 9 3 13 0 2
12 10 9 13 7 13 10 9 2 0 9 1 2
25 10 11 0 9 10 0 10 9 10 9 2 3 0 0 2 0 9 0 7 0 0 0 9 13 2
10 9 2 9 9 2 10 9 13 3 2
10 10 0 9 12 9 7 12 9 13 2
17 10 9 9 1 10 0 0 9 7 10 11 11 13 3 10 9 2
12 11 11 9 3 3 13 10 0 9 0 9 2
25 10 15 0 9 13 2 10 9 1 3 9 13 13 10 0 9 9 2 7 0 9 13 9 13 2
8 15 3 13 3 10 9 9 2
6 0 9 3 9 0 2
43 10 0 0 9 0 0 2 0 0 7 0 9 13 3 10 9 9 2 7 10 0 9 13 3 10 9 2 13 10 0 0 9 0 9 0 0 9 10 12 0 9 9 2
23 11 11 2 11 2 13 2 9 15 2 16 10 12 0 9 12 9 2 12 0 9 13 2
25 10 9 9 10 9 3 3 0 13 13 10 9 0 9 10 0 9 2 7 10 9 9 13 15 2
22 10 0 9 1 15 3 13 9 10 9 2 16 10 9 0 9 15 9 3 13 15 2
25 10 0 9 2 7 10 0 0 9 9 0 9 10 11 11 11 13 3 10 9 10 0 0 9 2
10 15 2 10 0 1 2 10 9 13 2
32 11 11 13 2 10 0 9 13 10 0 9 0 0 9 2 7 0 9 7 9 13 15 2 16 10 0 9 0 9 9 13 2
13 0 13 10 9 10 0 7 0 9 9 0 9 2
16 10 9 9 1 7 10 0 9 0 2 0 10 11 11 9 2
11 10 9 13 10 9 2 0 9 0 13 2
15 10 9 3 13 10 9 2 7 0 2 16 10 9 13 2
19 10 11 0 7 10 0 7 0 9 9 13 10 0 7 0 9 9 9 2
20 10 0 7 0 9 9 9 13 15 2 16 10 9 3 10 9 10 9 13 2
28 16 0 9 3 3 12 0 9 13 2 0 2 16 3 12 12 9 13 10 9 10 0 12 9 10 0 9 2
15 16 10 9 9 1 15 9 13 2 3 0 10 0 9 2
19 16 10 9 10 9 1 10 9 3 13 2 10 10 9 13 12 9 13 2
8 10 9 13 10 9 9 7 2
23 16 10 9 12 9 1 13 10 9 2 16 13 10 0 9 2 10 12 0 9 13 9 2
22 10 0 9 0 13 10 2 9 1 9 2 9 2 7 3 13 0 10 9 0 9 2
18 10 0 9 0 9 9 13 3 10 9 1 10 11 11 9 0 9 2
24 11 11 2 10 11 11 11 11 0 9 9 13 2 16 10 9 12 9 13 10 0 9 9 2
46 10 9 7 10 9 9 1 9 0 9 3 13 2 16 10 9 13 10 9 10 9 9 2 13 10 9 2 0 13 2 10 9 7 2 3 10 9 10 12 0 9 2 12 9 13 2
30 10 0 9 1 10 9 7 10 9 2 7 10 0 0 9 7 13 2 10 3 0 9 13 14 10 9 7 10 9 2
18 11 11 2 10 0 9 9 9 13 2 16 10 9 13 10 9 9 2
20 10 9 10 9 1 3 10 0 9 1 13 13 2 15 15 0 3 3 13 2
15 9 1 10 0 9 1 10 0 9 13 2 12 0 9 2
29 10 9 9 3 13 3 2 16 3 10 0 9 2 9 9 13 2 0 9 10 9 1 0 0 9 1 3 13 2
13 10 9 0 9 12 9 13 0 10 11 11 9 2
9 10 9 3 13 7 12 13 3 2
25 10 11 11 0 9 10 0 9 9 3 12 9 12 9 13 3 10 3 0 9 0 9 0 9 2
33 10 11 11 15 13 2 16 3 2 16 10 9 9 10 0 9 3 13 3 10 11 11 0 11 11 11 0 9 9 10 9 3 2
25 11 11 2 10 11 11 9 1 3 15 13 9 2 7 15 2 16 10 12 9 0 9 10 9 2
19 13 15 2 16 10 9 9 13 9 10 0 9 9 2 15 10 9 13 2
14 10 11 11 13 13 2 16 10 9 10 9 13 13 2
31 15 7 13 2 10 0 11 11 0 0 0 9 13 9 2 7 9 10 0 2 9 0 2 0 2 3 0 9 13 14 2
24 11 11 2 10 0 11 11 9 0 9 1 7 10 11 11 13 10 11 11 11 0 9 1 2
33 3 13 2 10 11 11 10 0 9 4 13 2 7 16 3 12 9 13 10 9 2 15 15 3 10 11 11 7 13 3 3 9 2
40 15 0 9 15 2 3 12 0 0 9 13 15 2 7 13 2 16 3 10 3 0 9 2 13 2 10 0 9 2 15 3 10 3 0 9 0 10 0 9 2
18 10 0 9 10 9 12 12 0 11 0 9 7 13 10 11 11 11 2
39 11 11 11 2 10 11 11 0 9 1 7 3 0 0 9 0 13 10 12 9 10 9 9 9 0 9 2 3 10 0 0 9 0 9 3 3 13 15 2
34 3 13 2 0 0 9 10 11 11 10 9 13 9 1 2 7 15 7 0 2 16 10 11 3 9 3 13 0 0 9 10 11 1 2
18 10 0 9 9 13 10 9 2 7 10 9 3 10 0 9 13 9 2
21 10 9 7 3 3 9 0 9 2 7 10 3 0 0 0 9 7 3 13 13 2
11 10 0 9 3 13 10 9 7 10 9 2
33 10 10 9 10 9 1 13 2 7 3 15 7 13 10 0 0 9 7 10 9 15 13 2 16 10 0 0 9 7 9 4 13 2
36 10 9 10 0 9 10 9 13 13 9 9 2 13 3 10 11 11 0 9 10 11 11 11 1 0 2 10 9 0 0 7 0 9 0 9 2
23 10 0 9 3 0 0 9 13 2 7 3 10 9 3 9 9 2 3 10 9 13 3 2
22 3 15 10 9 15 2 16 10 0 0 9 3 13 10 9 10 9 2 16 0 9 2
6 10 9 15 10 9 2
29 11 10 9 10 9 13 2 7 10 9 3 15 13 2 16 10 9 9 13 10 0 9 7 16 0 9 13 15 2
23 10 9 9 13 10 9 7 2 7 10 12 0 0 9 0 9 12 9 1 12 9 13 2
22 10 0 9 9 3 3 10 0 9 13 2 7 10 9 12 9 12 9 9 1 13 2
20 10 9 0 9 13 10 0 10 9 2 7 13 10 2 9 2 0 9 7 2
24 10 11 0 9 0 9 11 2 16 3 13 0 0 9 2 0 9 7 3 3 0 9 13 2
15 10 9 0 10 9 0 3 10 9 9 2 16 10 9 2
16 3 3 10 9 13 10 9 2 15 13 10 9 9 10 9 2
15 3 10 9 9 3 10 9 9 2 7 10 0 9 9 2
21 3 3 3 3 0 9 2 16 10 0 9 10 9 9 7 9 9 0 9 13 2
23 10 9 1 10 9 9 3 3 3 3 10 0 9 13 2 10 9 12 9 13 3 9 2
20 10 9 9 13 2 16 10 12 0 0 9 0 9 12 9 1 12 9 13 2
23 11 11 1 10 0 9 10 9 7 10 9 7 3 13 7 10 9 13 13 0 9 7 2
36 10 0 9 0 12 9 10 0 9 12 2 10 9 12 9 13 2 7 3 12 12 9 0 9 13 3 2 13 11 11 2 10 11 0 9 2
16 10 9 0 9 0 2 7 12 9 13 10 0 9 12 9 2
9 10 9 10 9 0 9 13 9 2
24 10 0 9 1 10 0 9 13 9 2 7 15 3 13 0 13 9 7 3 3 13 10 9 2
49 10 9 0 2 13 2 15 7 2 16 10 9 9 10 0 0 0 9 12 9 2 10 9 12 9 13 14 2 15 3 3 10 2 16 15 13 2 16 10 9 9 10 0 9 3 13 10 9 2
13 0 9 13 15 7 2 16 10 0 9 0 13 2
29 10 0 0 9 10 0 9 10 9 9 13 2 7 15 3 10 0 9 13 0 9 2 7 9 13 10 0 9 2
15 15 1 11 11 1 0 0 9 0 9 2 9 13 13 2
17 10 9 7 9 2 10 9 7 10 9 3 3 13 0 9 13 2
27 10 9 2 10 9 2 10 9 7 10 9 0 9 3 0 0 9 2 10 10 9 3 0 9 13 13 2
23 10 9 2 10 9 2 10 9 2 10 9 2 10 9 7 10 9 7 3 0 9 0 2
26 10 3 0 0 0 9 3 0 9 2 16 10 9 9 13 3 15 10 10 9 2 15 9 13 13 2
13 10 9 15 10 9 2 7 13 3 10 0 9 2
15 10 0 9 1 0 0 10 9 2 3 0 10 0 9 2
58 16 2 11 10 0 9 9 13 3 10 0 0 9 13 9 7 9 2 3 3 7 0 10 9 2 7 15 3 2 3 10 0 9 3 2 0 10 0 7 0 10 0 0 9 2 13 3 10 11 11 11 11 9 3 0 0 9 2
23 10 9 1 13 11 11 0 0 9 2 3 10 0 7 0 9 9 0 11 11 11 9 2
29 9 3 13 2 10 0 9 9 3 3 10 13 15 2 16 10 0 9 11 3 13 0 2 7 13 3 0 9 2
40 3 3 10 11 7 10 11 0 9 9 13 15 13 2 7 3 2 16 10 0 0 9 0 11 11 11 0 13 9 10 12 9 0 9 2 10 0 9 9 2
18 3 3 0 3 2 16 10 9 9 0 9 13 3 10 0 0 9 2
32 10 11 0 9 10 1 15 13 2 10 0 9 9 0 13 9 2 16 9 7 9 2 7 0 13 2 16 3 7 3 9 2
18 10 0 0 10 9 7 0 2 0 13 7 10 9 7 9 0 9 2
19 0 13 0 9 10 12 9 10 0 9 2 16 10 12 7 10 9 0 2
15 0 2 0 2 9 0 10 9 0 9 9 13 10 0 2
28 9 9 0 13 2 16 12 9 3 2 12 9 1 10 9 0 2 12 9 1 0 2 12 9 1 0 2 2
14 10 9 9 3 10 0 9 9 7 10 9 9 13 2
8 10 0 9 0 9 3 0 2
14 10 0 9 9 3 13 10 3 3 3 9 0 9 2
42 10 9 0 0 0 11 0 9 0 9 10 9 9 0 12 9 0 9 3 12 9 1 13 2 7 0 9 1 10 0 9 0 9 3 0 12 9 7 13 10 9 2
33 2 10 9 10 9 9 1 15 7 9 13 2 16 10 11 2 10 11 11 11 2 9 13 2 10 9 0 13 10 0 9 2 2
25 0 0 9 1 2 16 10 9 0 9 1 3 13 9 13 2 10 9 2 0 9 2 3 13 2
16 7 13 10 0 9 7 2 13 2 15 1 10 0 0 9 2
26 10 9 0 9 0 9 10 0 9 2 15 1 10 0 0 9 9 2 7 10 0 9 0 9 13 2
13 10 9 12 0 0 9 7 0 12 0 9 13 2
33 11 11 9 10 9 3 13 3 15 10 9 2 16 10 9 10 0 9 12 9 13 2 16 10 9 0 9 0 12 9 1 13 2
26 10 9 7 10 9 12 0 9 13 10 10 9 2 16 10 2 0 9 2 9 12 9 0 9 13 2
25 10 9 0 0 9 9 7 13 10 9 9 2 7 10 9 9 3 12 9 10 0 9 13 3 2
19 10 9 3 3 12 0 0 9 3 10 16 12 9 13 3 3 10 9 2
20 11 11 2 10 11 11 11 9 7 3 13 10 9 0 9 10 2 9 2 2
24 13 2 9 1 10 9 0 0 9 2 10 9 7 10 9 9 2 3 3 3 13 10 9 2
14 3 10 9 9 3 10 0 9 0 10 9 9 9 2
18 10 9 3 13 2 9 9 1 3 3 10 9 13 3 10 9 11 2
14 10 9 3 12 9 0 0 0 9 10 0 9 0 2
18 10 9 10 0 9 10 9 13 2 10 1 10 9 9 7 10 9 2
39 10 9 7 15 10 0 9 0 9 11 11 13 9 13 9 10 11 11 11 11 11 11 2 10 11 11 11 11 2 7 10 11 11 1 0 0 9 9 2
12 10 9 0 2 9 0 9 10 9 13 3 2
6 10 9 10 9 13 2
21 10 0 9 2 9 2 9 2 9 2 9 2 9 2 0 9 3 3 13 9 2
12 10 9 0 0 9 10 0 9 9 13 0 2
9 10 0 9 13 15 10 9 7 2
22 10 9 13 10 9 9 2 10 9 2 7 10 9 2 3 0 9 10 9 9 9 2
7 10 9 9 0 9 13 2
12 10 9 9 9 10 9 13 2 9 13 9 2
7 10 9 7 9 7 13 2
20 15 0 9 3 2 16 10 0 9 9 3 3 13 10 0 9 2 16 3 2
17 3 12 9 7 13 10 12 1 2 3 10 10 9 0 12 9 2
19 10 0 9 9 10 0 12 9 1 3 3 12 9 1 13 10 0 9 2
19 10 9 10 9 0 9 13 2 7 3 13 10 9 0 9 1 0 9 2
18 0 9 1 0 2 16 10 9 3 3 13 10 9 9 0 0 9 2
17 10 9 1 10 10 2 9 7 0 2 2 9 2 3 4 13 2
11 10 0 9 9 1 7 15 3 0 13 2
24 10 9 0 0 9 2 10 0 2 10 0 7 10 0 9 2 0 9 1 13 2 3 13 2
19 3 13 3 0 9 2 16 10 0 9 10 0 9 9 15 3 13 13 2
21 3 10 9 12 0 2 10 0 2 10 0 2 10 11 2 9 0 0 9 13 2
15 10 0 9 7 0 10 9 2 3 10 9 7 13 13 2
20 10 9 0 9 1 3 3 10 0 0 9 13 2 7 0 9 2 10 9 2
16 10 0 9 0 13 2 0 13 2 7 15 1 3 13 9 2
7 3 10 9 0 9 13 2
16 15 7 9 2 10 3 12 9 0 0 0 9 10 0 0 2
8 13 10 9 2 3 0 13 2
18 15 3 0 9 2 7 13 2 16 10 9 10 9 9 3 13 13 2
7 3 13 10 0 9 11 2
16 0 9 0 10 0 9 9 2 10 9 9 2 10 9 9 2
5 15 0 9 13 2
34 10 0 9 0 9 2 16 10 9 0 2 0 9 3 10 0 12 9 13 3 2 7 15 0 9 15 2 16 10 9 9 7 13 2
28 14 13 13 10 9 0 9 2 10 0 9 2 10 10 9 13 10 0 9 2 2 10 0 0 7 0 9 2
22 10 0 9 10 0 0 9 9 2 15 3 3 0 2 7 10 9 1 10 13 11 2
15 0 9 13 10 0 9 2 7 10 9 2 10 9 9 2
9 0 10 0 9 0 0 9 9 2
22 15 9 9 13 13 10 9 2 10 9 2 10 9 2 7 10 9 2 0 9 2 2
25 10 9 3 10 9 9 2 10 9 9 2 10 9 9 13 9 13 2 3 0 0 13 10 9 2
8 3 12 9 13 10 0 9 2
15 10 0 9 9 0 13 2 16 15 3 10 0 9 13 2
23 15 15 0 2 16 10 0 0 0 9 1 3 0 9 13 2 15 0 13 10 9 9 2
21 10 0 9 13 3 1 2 9 3 3 4 13 10 0 0 9 2 9 2 9 2
11 0 13 10 10 9 13 10 0 9 7 2
10 2 3 10 0 9 0 0 9 13 2
36 3 10 9 7 10 9 13 10 9 10 0 9 2 10 0 9 9 7 10 9 9 13 2 10 9 0 9 13 2 10 0 9 7 13 2 2
10 0 9 13 2 16 10 0 9 13 2
26 10 9 2 7 10 0 9 9 0 13 10 0 2 10 9 0 9 3 3 13 10 0 0 9 9 2
6 10 0 9 13 4 2
9 15 9 9 0 0 0 9 0 2
26 10 0 9 10 9 2 15 3 7 13 3 2 7 10 0 9 3 0 13 2 16 15 10 9 13 2
7 10 9 9 9 13 4 2
12 13 11 10 9 2 10 0 2 0 9 9 2
7 10 9 0 12 0 13 2
9 9 3 3 13 14 10 11 11 2
17 10 9 9 10 11 11 11 0 9 9 0 9 3 12 9 13 2
19 10 0 9 2 12 3 12 2 3 3 10 16 12 9 13 14 10 9 2
17 10 9 9 15 0 13 2 3 3 12 9 1 13 10 0 9 2
22 10 0 9 3 9 2 9 2 9 13 10 9 2 3 0 10 0 9 7 13 9 2
10 10 9 1 12 9 12 9 7 13 2
26 10 9 3 10 0 9 1 0 9 2 9 7 13 2 7 10 9 7 13 2 15 3 13 0 9 2
37 10 9 3 9 13 10 12 0 11 11 9 2 15 10 9 9 13 14 3 10 9 2 3 13 2 13 2 3 13 3 9 2 9 10 9 9 2
28 10 9 3 10 0 9 0 2 10 0 9 7 13 9 2 13 10 9 2 9 13 10 9 2 0 9 13 2
11 10 9 0 9 10 12 9 0 11 11 2
15 10 9 10 9 3 0 2 16 0 10 9 7 10 9 2
26 10 9 12 9 2 0 9 13 10 9 2 10 9 7 0 9 2 0 9 9 13 3 10 0 9 2
22 10 0 9 9 3 13 2 16 10 0 0 9 3 10 9 13 15 10 9 10 9 2
22 10 9 0 9 2 9 0 7 3 9 2 16 3 3 12 9 1 3 3 13 9 2
2 13 2
20 10 0 9 9 1 10 11 3 12 9 0 0 9 9 7 13 10 9 9 2
5 7 3 13 3 2
4 3 13 15 2
25 0 9 13 3 15 10 11 11 11 11 9 3 9 2 7 3 7 3 2 10 11 11 0 9 2
10 10 0 0 9 9 0 13 10 9 2
13 13 2 16 10 3 0 9 9 1 3 13 13 2
12 7 10 0 9 10 9 1 3 9 13 15 2
5 9 1 15 13 2
9 13 10 9 1 2 15 10 9 2
6 10 9 3 0 9 2
12 0 2 0 2 9 2 7 13 10 9 9 2
21 10 11 11 11 11 9 13 14 2 16 10 10 9 3 10 9 13 9 10 0 2
17 0 3 2 3 10 0 9 1 13 10 9 9 10 9 12 9 2
11 10 10 9 10 9 3 3 13 10 9 2
7 13 15 10 9 0 9 2
13 7 15 13 10 9 9 9 1 0 0 9 7 2
19 10 0 9 3 3 3 13 14 0 9 2 7 3 13 9 0 10 9 2
21 10 9 9 12 9 2 12 9 7 10 9 2 10 11 0 9 9 10 9 9 2
5 13 15 9 1 2
7 7 7 9 13 10 9 2
23 10 9 9 2 0 15 7 0 9 10 2 0 2 9 2 3 13 9 13 10 9 9 2
15 2 3 10 0 9 13 10 9 2 3 0 13 10 9 2
21 10 9 13 10 9 2 3 10 0 9 13 10 9 9 2 7 3 10 9 7 2
17 3 15 13 2 0 13 10 9 10 9 2 2 2 13 11 11 2
25 10 9 13 3 15 7 2 16 10 10 0 9 0 12 9 1 13 2 10 9 1 2 15 13 2
13 2 3 13 15 13 2 16 15 7 13 10 9 2
18 7 10 9 0 9 15 3 0 2 2 13 15 10 0 0 9 9 2
13 11 11 0 9 7 13 3 10 9 2 7 0 2
16 9 9 0 9 7 9 13 3 3 2 7 9 3 7 2 2
13 2 0 0 10 9 0 2 10 9 0 10 9 2
11 10 9 7 10 9 7 3 13 2 13 2
11 10 9 10 0 9 3 13 2 9 1 2
16 3 3 15 13 3 15 10 12 0 9 2 2 13 11 11 2
9 10 0 0 9 3 15 10 9 2
7 10 9 9 7 3 13 2
18 15 1 10 2 0 9 2 9 0 11 11 11 13 10 9 11 9 2
8 3 9 3 13 10 0 9 2
8 2 10 15 9 3 13 2 2
15 12 9 1 7 15 13 13 2 10 0 9 7 13 9 2
17 10 9 3 0 9 0 9 3 0 9 13 2 0 13 10 9 2
22 3 3 13 10 9 2 3 3 13 10 9 2 7 10 9 11 3 13 13 10 9 2
11 2 15 15 13 2 2 13 10 9 9 2
16 2 13 15 2 13 15 2 13 2 3 15 13 15 3 2 2
6 10 9 0 9 13 2
9 0 9 1 3 12 9 13 3 2
9 10 10 9 3 10 9 3 13 2
9 10 0 9 1 0 13 10 9 2
6 14 3 13 10 9 2
16 13 2 15 13 2 16 0 9 13 2 15 3 13 13 15 2
12 7 10 9 3 12 9 13 3 10 0 9 2
6 10 9 3 7 13 2
11 10 9 7 10 9 9 7 3 13 3 2
7 13 2 3 3 0 13 2
17 0 9 13 2 15 13 2 13 10 9 1 2 7 13 10 9 2
11 3 0 9 2 7 9 0 14 13 13 2
11 15 7 9 13 10 9 2 0 3 13 2
11 10 9 3 3 10 9 7 10 9 13 2
12 10 9 1 0 9 7 9 13 15 10 9 2
4 13 10 9 2
24 10 9 7 3 10 9 7 13 2 3 3 2 16 10 9 3 10 9 2 7 10 9 13 2
18 3 10 11 9 13 10 9 2 11 2 11 7 11 7 9 1 13 2
18 10 0 9 7 0 9 13 15 2 15 7 3 10 9 3 13 3 2
9 15 15 13 9 10 0 2 9 2
16 10 9 3 11 11 2 11 11 7 11 11 0 0 9 13 2
13 11 11 2 11 11 13 3 10 9 10 0 11 2
11 10 9 0 3 0 10 9 2 9 9 2
16 15 7 3 13 13 2 3 13 3 3 10 9 0 0 9 2
30 7 15 3 2 16 9 13 3 3 2 16 3 9 13 13 10 0 9 7 9 13 9 10 3 3 0 0 9 1 2
12 10 9 2 9 3 10 9 13 3 10 9 2
19 0 13 12 11 0 9 2 7 9 1 13 10 11 0 11 12 9 7 2
13 10 0 9 0 9 1 0 9 13 10 0 9 2
25 11 13 10 0 10 9 2 12 9 3 3 13 13 2 7 0 13 9 10 9 11 7 11 7 2
26 10 9 10 10 9 7 3 9 2 0 9 13 13 2 13 9 11 11 9 2 10 0 0 9 9 2
11 3 3 12 9 7 9 0 9 13 9 2
12 0 9 13 10 11 0 12 0 9 9 7 2
15 10 9 10 11 11 9 13 2 9 13 9 11 7 11 2
18 10 9 7 10 9 9 10 9 0 9 7 10 9 0 9 11 13 2
11 10 9 3 9 7 9 0 9 13 3 2
37 10 9 10 0 9 10 0 9 13 2 7 16 3 13 13 2 10 9 7 9 9 3 0 13 9 2 13 11 11 2 10 11 11 11 11 9 2
9 9 13 9 10 9 10 9 7 2
20 11 11 10 0 9 9 13 10 9 11 7 10 0 9 1 12 0 9 1 2
21 10 9 0 9 2 9 1 13 9 2 13 11 11 2 10 11 11 11 11 9 2
14 10 9 9 13 2 16 13 3 0 9 10 9 1 2
23 15 7 10 9 9 1 13 9 2 16 10 9 13 10 9 2 3 3 13 3 10 9 2
13 3 11 11 2 10 11 9 13 2 3 13 9 2
10 3 0 9 13 3 10 9 9 1 2
12 11 10 9 0 9 13 3 2 10 9 0 2
20 10 0 9 13 2 7 0 0 7 0 9 13 3 2 13 9 11 11 9 2
30 11 10 0 9 9 13 10 15 9 2 7 15 3 0 9 13 3 2 13 9 11 11 2 10 11 11 11 11 9 2
17 10 0 9 3 0 9 13 3 2 3 13 9 2 9 10 15 2
17 10 9 10 11 0 9 9 13 2 3 3 12 9 13 10 9 2
13 11 7 11 1 2 7 11 12 9 3 13 9 2
10 10 0 9 1 3 11 13 10 9 2
19 10 11 11 0 9 1 3 13 10 11 7 11 11 11 11 0 9 9 2
15 3 13 10 11 10 0 9 7 2 16 15 10 9 13 2
13 9 13 10 0 9 1 0 9 9 0 0 9 2
19 10 11 11 11 11 11 11 1 0 9 9 10 9 0 9 2 11 11 2
22 10 0 0 9 10 0 0 9 13 14 2 15 9 7 10 9 7 10 0 9 13 2
31 10 11 0 9 9 13 10 11 11 2 10 11 2 10 11 11 11 2 10 11 11 2 10 11 11 2 10 11 11 7 2
7 9 1 9 13 0 11 2
14 12 9 1 3 3 13 14 10 0 9 10 0 9 2
24 3 3 10 9 10 9 12 7 12 0 9 13 10 9 2 10 9 7 10 9 9 13 3 2
8 10 9 3 10 9 13 9 2
12 3 3 13 9 2 16 3 10 0 13 9 2
11 11 0 9 7 10 9 9 13 10 9 2
17 10 0 9 3 3 13 3 10 9 2 10 9 7 0 9 13 2
13 11 10 0 9 1 12 9 13 9 1 9 9 2
33 0 9 1 11 11 12 2 11 11 12 2 11 12 2 11 12 2 11 11 12 2 11 12 2 11 7 12 9 2 9 13 9 2
18 10 9 0 0 9 1 10 11 0 9 9 1 9 13 10 0 9 2
11 11 9 10 0 9 1 0 9 13 3 2
22 10 3 12 12 0 9 3 13 12 9 7 12 9 2 7 13 10 9 10 9 7 2
22 11 11 11 7 11 10 9 7 10 9 3 12 9 0 13 3 10 9 7 10 9 2
15 12 9 9 13 10 9 2 7 10 13 9 13 9 7 2
17 10 0 9 0 13 10 9 2 10 9 9 10 16 12 9 13 2
13 10 9 3 13 0 13 2 0 2 0 9 13 2
17 11 10 9 1 10 16 12 9 3 13 13 10 0 9 10 9 2
10 9 13 10 0 9 10 11 11 7 2
21 11 11 10 0 2 0 9 10 16 12 9 2 15 9 0 12 9 2 13 15 2
14 12 9 9 13 2 7 10 9 0 9 13 9 13 2
8 2 10 9 13 10 0 9 2
36 10 0 0 9 2 16 13 2 9 13 15 2 15 10 9 10 3 9 2 10 10 3 9 0 2 7 10 0 9 9 3 10 9 7 0 2
18 3 13 10 9 0 9 2 15 3 13 2 16 3 15 2 15 2 2
7 10 9 0 9 10 9 2
12 3 16 15 1 10 0 9 13 4 10 9 2
14 3 3 2 9 13 2 9 13 2 15 10 9 13 2
16 10 0 9 9 13 10 0 9 11 2 15 13 10 9 9 2
11 3 13 2 16 15 10 0 0 9 13 2
22 10 0 2 0 9 9 7 3 3 13 10 9 0 9 2 15 0 7 0 9 13 2
22 11 11 12 8 9 10 11 11 9 15 13 2 16 13 2 16 9 0 13 10 9 2
27 10 9 0 13 10 0 7 10 0 9 0 3 0 9 2 7 9 3 13 10 9 2 16 9 9 13 2
9 7 10 9 13 2 7 3 13 2
31 11 12 0 9 0 0 0 9 3 13 0 0 10 0 9 2 16 15 3 13 0 9 10 9 1 2 16 10 9 9 2
6 10 9 0 9 13 2
15 13 10 9 2 7 15 9 9 13 2 9 7 9 13 2
31 9 13 3 10 0 0 9 2 10 9 0 2 0 2 0 9 9 3 9 2 9 2 10 3 13 3 9 9 13 3 2
22 10 9 9 10 9 9 3 3 13 2 3 0 13 2 10 0 9 9 0 9 13 2
12 10 9 0 9 13 3 2 16 10 9 13 2
37 15 15 13 2 15 3 10 2 16 9 0 9 2 15 9 10 9 7 3 10 9 0 3 13 2 3 13 10 9 2 7 3 10 0 9 3 2
7 10 9 13 10 0 9 2
36 10 0 0 9 2 16 13 2 9 13 15 2 15 10 9 10 3 9 2 10 10 3 9 0 2 7 10 0 9 9 3 10 9 7 0 2
35 3 13 10 9 0 9 2 15 3 13 2 16 3 15 2 15 2 3 10 9 2 15 9 1 10 9 9 9 3 0 10 0 9 7 2
34 15 13 2 16 10 9 3 3 9 13 2 3 11 10 9 0 2 7 15 2 16 12 0 9 13 9 2 15 9 1 3 13 13 2
46 10 9 9 10 9 10 0 9 9 9 2 15 15 3 0 13 2 16 0 9 1 13 10 9 9 2 7 15 3 0 13 2 16 10 0 9 9 9 0 13 10 9 9 0 9 2
35 13 10 0 0 9 10 0 9 2 10 0 9 2 15 9 3 10 9 2 10 9 2 10 9 2 10 9 9 2 10 0 0 9 0 2
26 10 0 9 9 0 0 9 9 2 16 3 15 13 9 13 2 15 3 13 3 7 3 3 13 3 2
32 16 10 9 9 1 0 2 7 0 9 10 9 1 3 7 3 0 0 9 13 2 10 0 9 13 10 9 2 13 10 9 2
12 15 0 13 2 15 3 13 9 2 0 9 2
33 10 0 0 0 9 0 13 10 9 10 0 9 1 2 15 1 13 7 3 3 13 9 2 15 13 10 0 9 1 0 9 9 2
15 16 10 10 9 10 9 15 13 2 15 13 2 15 13 2
5 7 15 3 13 2
15 13 9 10 0 0 9 2 15 10 9 9 13 3 3 2
41 10 11 11 9 0 0 9 9 0 9 10 3 3 10 15 9 0 2 0 9 0 0 9 9 13 10 0 9 0 9 2 15 9 10 9 0 9 13 9 9 2
32 10 9 3 13 2 16 10 9 9 13 2 7 15 3 13 2 16 10 9 9 0 7 0 9 13 14 10 0 9 0 9 2
12 10 9 9 3 3 13 2 16 15 10 9 2
42 13 2 16 0 13 15 10 11 1 3 0 0 9 2 3 10 9 9 13 10 2 16 3 13 2 0 9 2 15 9 2 9 2 9 2 9 2 0 9 13 9 2
19 15 10 9 9 9 13 2 7 0 3 9 2 10 0 9 12 9 13 2
45 10 10 9 13 10 15 0 0 2 15 10 9 3 13 2 3 10 10 9 10 0 13 2 15 9 2 9 2 9 13 10 0 9 2 10 0 9 7 15 13 15 2 16 15 2
5 10 9 15 13 2
11 10 9 9 9 0 13 10 0 8 9 2
13 9 13 2 3 10 9 10 0 13 10 0 9 2
14 0 9 13 3 2 3 9 0 9 13 0 0 9 2
18 16 9 13 2 3 15 13 9 16 11 9 3 11 13 2 3 11 2
7 10 9 9 10 9 9 2
19 10 9 2 15 13 2 3 10 9 2 7 3 13 2 15 3 10 9 2
33 16 3 0 2 16 13 2 13 7 3 3 4 2 10 0 9 0 9 1 3 13 13 10 15 0 9 2 15 9 0 9 0 2
28 10 9 10 3 13 10 9 1 0 0 0 9 2 15 0 7 0 13 10 9 2 15 9 0 9 13 13 2
7 7 3 0 10 9 9 2
28 0 9 13 10 0 9 2 3 15 15 15 2 15 11 13 2 16 2 10 9 3 0 13 10 9 0 9 2
22 16 3 3 13 2 7 3 13 3 2 3 15 13 10 9 0 9 2 16 13 0 2
11 13 2 15 3 3 10 9 1 13 14 2
50 3 13 15 2 16 9 12 9 7 13 9 9 9 2 7 15 2 7 10 3 13 14 15 2 15 7 3 13 2 16 3 3 13 2 3 0 9 13 14 2 3 16 13 3 9 10 0 9 9 2
10 13 10 0 9 2 15 0 9 13 2
9 7 0 9 13 15 2 0 7 2
32 9 13 2 7 0 9 13 10 9 9 2 9 9 2 13 15 10 11 8 0 9 2 3 13 2 16 9 10 0 9 9 2
8 11 11 13 15 2 9 9 2
5 9 0 0 13 2
15 10 9 13 3 2 7 3 16 0 13 3 10 0 9 2
23 9 2 3 2 9 2 3 13 7 0 2 7 0 9 2 10 9 3 3 0 9 13 2
28 3 3 12 9 1 10 9 3 3 10 0 9 9 13 9 2 3 2 0 9 9 2 13 10 0 9 9 2
8 3 10 0 9 15 7 13 2
27 9 2 9 2 3 3 3 13 10 9 2 9 10 9 2 10 0 9 2 7 9 11 2 10 0 9 2
37 10 9 0 9 10 10 9 2 10 0 9 10 15 3 13 10 10 0 9 2 7 10 10 12 9 2 15 10 0 9 13 2 3 13 11 11 2
28 10 9 3 3 3 13 2 10 9 1 0 7 2 7 15 15 13 2 16 3 15 13 2 9 9 9 13 2
11 0 10 9 2 16 10 0 9 10 9 2
10 7 10 3 0 9 10 9 0 9 2
37 12 9 13 3 10 0 9 10 9 2 16 15 10 11 9 2 10 11 7 10 9 9 2 9 13 2 7 3 2 10 9 9 13 10 9 9 2
19 10 0 9 9 2 10 9 7 9 2 10 9 2 10 9 13 10 15 2
7 10 0 0 12 9 13 2
8 2 11 10 0 9 13 2 2
19 10 0 9 9 1 0 9 13 10 9 9 7 2 10 3 3 9 9 2
15 3 10 0 9 2 9 0 9 13 4 2 13 10 9 2
13 11 9 3 3 0 2 3 9 7 9 13 3 2
28 10 9 9 3 13 9 2 7 16 2 13 2 3 2 15 9 7 9 2 13 2 16 10 9 13 2 13 2
21 9 2 9 3 13 0 2 10 9 9 13 10 9 2 2 3 3 9 13 9 2
9 10 9 9 1 7 13 7 9 2
6 16 9 3 3 13 2
5 7 13 10 9 2
7 10 9 2 11 9 13 2
33 10 0 9 2 10 0 0 9 2 10 9 9 2 10 9 2 10 9 9 2 10 12 0 9 9 7 9 10 0 9 2 13 2
42 7 9 7 9 2 3 10 9 9 2 0 7 0 9 11 2 2 3 10 0 2 10 0 2 10 0 2 10 0 0 9 9 9 7 10 0 9 9 13 10 9 2
25 11 15 13 2 16 10 0 7 10 0 9 3 13 10 9 2 3 3 0 13 2 15 13 15 2
19 0 9 1 13 2 10 9 10 9 13 10 9 2 3 7 0 9 13 2
23 11 13 10 9 2 16 0 0 9 13 10 0 9 2 15 0 9 9 13 10 0 9 2
11 2 15 10 15 9 2 2 2 13 11 2
20 2 0 9 3 13 2 2 13 11 2 15 0 13 10 0 7 10 0 9 2
28 7 3 13 2 16 10 9 13 10 0 0 9 2 9 0 0 9 2 15 2 15 11 9 13 9 2 13 2
16 13 7 10 9 10 0 9 2 15 3 14 3 13 0 9 2
26 11 3 12 3 13 2 16 10 0 9 2 7 0 13 10 9 2 15 0 9 1 3 13 15 3 2
10 11 11 9 13 10 0 0 9 1 2
18 10 0 7 10 9 0 9 2 10 0 0 9 9 3 13 11 11 2
10 10 0 9 3 9 13 0 9 7 2
31 10 9 3 13 2 16 15 10 9 13 3 10 9 9 2 16 10 9 2 15 3 0 10 0 9 2 0 9 3 13 2
8 3 3 10 0 9 9 13 2
25 11 9 7 2 3 9 2 9 13 15 10 0 0 11 2 3 2 13 2 15 11 9 13 11 2
23 10 9 7 0 9 13 2 10 11 7 15 13 15 2 7 11 2 16 0 13 10 9 2
28 7 10 9 2 13 10 9 2 15 13 2 6 2 15 7 3 13 13 9 1 2 10 9 12 9 13 15 2
26 11 7 13 2 16 2 3 3 15 2 7 11 13 0 9 15 2 7 3 15 3 13 10 0 11 2
15 3 0 7 15 0 0 9 13 9 10 15 9 0 9 2
11 15 2 3 13 10 9 9 2 13 11 2
11 13 10 9 2 7 13 10 11 11 13 2
22 10 9 3 13 15 2 16 2 10 10 0 9 0 9 10 0 9 3 3 13 11 2
22 2 15 7 13 2 16 3 2 16 10 11 9 2 15 12 9 1 3 13 15 13 2
5 0 13 0 9 2
14 11 13 10 0 0 2 3 11 9 10 0 9 2 2
22 15 3 15 13 13 2 16 9 0 9 15 13 10 9 2 3 3 9 3 13 4 2
13 3 3 13 10 9 9 2 16 0 13 10 9 2
14 12 9 2 16 12 2 9 3 13 2 7 9 6 2
7 0 9 9 11 11 13 2
4 0 9 13 2
18 11 11 9 0 7 0 9 13 10 9 1 2 7 9 13 10 9 2
11 10 0 9 10 0 2 9 2 7 13 2
19 10 9 7 10 0 9 13 2 3 3 10 0 2 7 10 0 9 13 2
2 9 2
50 16 3 11 13 10 9 9 2 15 10 0 9 2 0 0 9 3 13 11 11 2 7 9 13 9 9 2 7 3 10 9 13 2 3 15 13 2 9 9 2 0 0 9 13 3 2 15 15 13 2
3 11 7 2
13 2 15 15 2 2 2 13 10 0 9 0 9 2
17 11 11 10 9 1 13 2 3 10 9 2 15 10 9 1 13 2
5 10 9 3 13 2
13 7 3 13 2 3 3 13 15 10 2 9 2 2
10 16 12 9 1 3 13 11 0 9 2
19 3 3 3 3 10 0 9 13 2 13 2 3 7 3 0 9 9 13 2
21 15 3 15 13 2 9 2 16 12 0 9 1 10 9 13 10 0 0 0 9 2
8 3 0 13 2 16 15 13 2
7 3 3 9 13 10 11 2
32 3 13 10 11 11 7 10 0 9 0 9 2 15 0 10 2 0 9 2 2 9 8 11 11 2 2 11 2 2 9 13 2
40 0 13 0 0 9 2 3 3 10 0 9 15 10 9 13 2 7 0 9 11 7 11 9 13 3 0 9 2 3 13 10 11 0 0 9 2 15 3 13 2
3 10 9 2
35 10 11 10 0 9 10 11 0 9 9 0 0 0 9 2 16 10 0 9 9 3 3 2 15 3 13 2 16 12 9 9 13 10 9 2
15 16 10 0 9 2 0 0 9 2 9 3 13 10 9 2
13 0 0 9 3 15 3 15 13 2 9 3 0 2
15 10 0 10 0 9 13 15 2 6 7 15 2 15 13 2
18 10 0 2 0 0 9 7 6 13 2 3 3 3 2 3 3 3 2
37 7 3 9 2 7 10 9 9 13 13 2 10 0 9 3 3 4 0 9 13 2 10 9 7 3 3 0 13 2 16 10 0 9 10 0 9 2
14 10 0 9 7 0 9 2 15 9 13 10 0 9 2
24 11 3 3 13 2 10 9 15 13 2 16 10 0 12 9 9 13 3 11 7 11 10 9 2
41 10 9 0 9 9 2 15 1 2 16 10 12 0 9 9 3 4 13 7 15 13 2 15 3 13 3 10 3 9 0 9 2 0 9 13 16 13 10 0 9 2
14 3 10 11 11 7 10 11 11 11 2 11 2 9 2
16 16 11 11 10 0 9 0 13 2 10 0 9 0 10 9 2
18 10 11 0 9 2 11 11 15 3 13 3 2 3 10 9 9 13 2
15 10 3 10 7 10 1 0 0 9 7 16 3 3 13 2
10 10 12 9 0 9 0 3 3 0 2
33 15 13 0 9 2 16 10 0 9 13 2 7 15 7 2 0 10 9 2 3 3 10 9 9 13 0 2 7 10 9 0 7 2
22 3 0 9 3 13 14 2 10 9 0 9 3 10 9 13 15 2 15 3 0 13 2
10 0 9 1 3 13 11 9 0 9 2
48 10 0 9 0 9 13 2 10 9 2 9 9 2 9 1 0 13 2 7 10 9 3 10 13 3 9 2 16 10 12 9 1 0 7 2 9 9 2 10 9 3 0 0 9 13 10 9 2
29 3 0 13 2 10 0 9 0 0 9 13 2 15 10 0 0 9 1 3 13 10 9 2 0 9 9 2 13 2
33 16 10 9 13 15 10 12 9 0 7 0 3 0 9 9 2 3 7 13 2 16 10 0 9 3 0 9 7 3 0 9 13 2
24 16 13 10 0 9 2 15 10 0 9 0 0 9 13 2 10 0 9 13 10 12 12 9 2
10 10 10 9 10 9 0 9 3 0 2
35 3 0 2 16 10 0 0 0 9 10 9 7 9 13 13 2 3 16 10 0 9 14 3 13 2 3 3 13 10 10 0 0 9 13 2
31 0 2 16 15 13 2 16 10 0 12 9 10 9 3 0 0 9 1 7 12 9 9 7 10 11 11 10 9 13 13 2
15 0 9 2 9 3 13 2 16 10 9 3 15 9 13 2
45 16 13 10 9 2 7 12 9 1 0 13 10 0 12 0 0 9 2 3 15 2 13 15 9 7 9 2 10 10 9 13 2 16 10 0 9 0 9 13 10 9 0 9 9 2
25 10 0 9 3 3 3 9 13 2 15 13 10 9 15 2 0 9 13 10 13 7 10 13 1 2
16 10 9 7 3 13 13 15 2 16 3 15 3 13 10 9 2
10 15 7 10 9 7 10 9 9 0 2
19 2 10 0 9 0 9 2 0 9 10 9 3 9 13 2 0 13 2 2
17 3 13 10 9 10 0 9 0 9 11 2 11 11 0 0 9 2
20 10 3 0 9 1 10 0 9 10 0 0 9 10 0 9 2 0 9 13 2
17 0 9 2 15 0 9 2 9 2 9 13 0 2 0 7 9 2
20 15 7 10 9 13 2 7 0 9 7 9 7 7 15 3 13 9 0 9 2
10 7 15 3 7 3 13 10 9 9 2
13 2 3 3 10 11 0 9 13 9 12 0 9 2
21 10 9 0 9 10 8 9 8 0 9 13 3 2 15 0 7 10 11 0 9 2
7 3 3 10 10 9 13 2
12 2 11 9 0 9 2 15 10 9 13 9 2
21 3 11 11 13 15 2 7 11 13 2 10 9 9 7 3 13 10 0 9 9 2
13 3 13 10 9 2 7 3 7 0 9 13 15 2
24 11 11 9 7 3 13 9 2 16 0 9 2 15 10 9 3 7 10 0 9 9 13 3 2
15 3 3 13 10 9 2 13 2 7 3 3 13 0 9 2
20 2 3 3 13 10 11 2 13 15 2 16 0 9 7 13 3 10 10 9 2
17 2 10 9 3 13 2 7 13 10 9 0 7 0 9 7 13 2
15 3 3 2 16 10 0 9 10 9 2 16 10 0 11 2
47 3 10 9 9 7 9 13 3 7 2 16 0 9 13 3 10 0 9 9 2 16 0 9 13 10 3 0 7 0 9 2 16 15 0 0 13 2 7 3 3 0 7 0 9 13 3 2
14 15 0 13 10 12 9 0 9 2 15 10 9 13 2
41 3 13 3 0 9 13 2 7 10 11 11 1 2 15 3 11 13 2 11 11 2 10 0 9 15 13 15 2 2 11 9 2 3 13 3 2 9 1 9 3 2
9 9 2 10 0 9 7 9 2 2
19 15 7 0 9 1 13 10 9 2 3 9 2 16 7 0 9 13 15 2
20 2 10 1 10 12 9 1 3 10 0 9 13 2 3 11 9 3 13 9 2
6 2 15 3 7 13 2
44 15 13 16 12 10 11 11 2 15 0 2 0 9 2 7 10 9 9 11 11 13 2 7 3 3 13 9 0 0 9 7 2 11 11 13 14 10 11 11 2 10 11 11 2
12 10 10 9 3 12 9 2 7 10 9 13 2
13 0 9 13 2 7 10 9 14 13 10 0 9 2
24 11 0 13 15 2 16 10 9 1 0 0 9 13 2 7 13 2 13 3 11 10 11 7 2
18 7 16 3 0 9 13 2 7 0 13 9 10 10 9 2 9 13 2
28 15 9 1 3 13 15 2 0 9 2 16 3 15 13 3 2 7 3 15 13 2 16 3 3 9 13 13 2
15 10 12 9 10 9 2 0 13 2 0 13 7 0 13 2
35 2 10 0 9 3 3 0 9 13 9 2 7 10 9 3 9 13 9 10 11 2 16 10 0 0 9 0 9 10 15 0 0 9 13 2
26 7 15 1 2 16 0 13 2 3 10 0 9 1 13 0 7 2 10 0 9 2 15 13 10 9 2
14 2 3 13 2 15 9 13 2 15 9 10 9 9 2
24 15 3 0 13 10 10 9 2 0 3 2 16 15 10 9 2 9 3 13 3 12 9 3 2
33 10 9 2 10 0 0 9 3 15 3 13 2 16 10 11 7 9 11 11 13 15 2 7 10 10 0 0 9 2 11 11 7 2
25 15 13 3 2 16 15 10 0 9 13 2 15 7 13 10 9 2 7 15 7 13 13 10 9 2
50 7 3 13 13 2 16 15 3 13 9 2 15 3 10 10 9 13 3 2 16 3 3 12 9 1 13 2 7 3 10 9 15 7 9 13 13 2 15 3 13 3 15 10 9 2 7 10 9 13 2
31 7 3 10 0 9 15 13 10 9 2 15 11 11 13 15 2 2 16 15 13 10 9 2 3 13 9 2 16 13 2 2
21 15 10 9 9 2 0 9 2 0 9 13 13 10 9 2 16 0 13 10 9 2
12 2 10 0 9 10 9 10 9 7 13 15 2
4 13 15 9 2
15 2 3 13 2 16 3 0 2 0 9 13 10 10 9 2
34 13 2 3 10 10 9 13 2 7 13 0 9 7 0 9 2 13 10 11 11 11 2 7 10 11 11 11 11 11 11 11 0 9 2
8 3 13 10 10 0 9 7 2
9 2 15 13 3 15 3 10 9 2
18 2 9 2 16 3 10 9 0 9 13 2 7 10 9 13 2 13 2
18 7 3 13 2 15 3 13 10 15 2 3 13 10 9 7 10 9 2
17 0 13 7 13 2 16 9 13 14 2 7 3 3 3 13 9 2
18 9 0 0 2 0 15 10 9 2 10 9 7 10 0 9 0 9 2
21 10 9 10 16 9 1 13 10 11 11 11 11 2 7 12 9 13 10 0 9 2
32 10 9 0 9 1 3 0 9 13 2 13 9 2 12 9 2 0 7 9 2 7 10 0 9 2 0 9 7 15 10 9 2
42 11 11 0 9 3 3 13 10 11 2 10 9 10 11 9 7 10 11 9 12 0 0 9 9 2 10 11 9 2 10 11 11 7 10 11 9 13 3 11 11 9 2
28 2 15 15 1 0 3 13 3 10 10 9 2 15 7 13 3 15 10 9 2 7 10 10 9 9 7 13 2
11 2 6 2 3 10 9 13 3 10 9 2
11 10 9 10 11 11 11 9 13 3 9 2
40 11 11 3 13 10 12 9 0 9 2 15 10 1 11 11 7 11 11 0 9 7 9 13 2 7 15 9 13 14 10 15 9 7 2 0 3 10 10 9 2
16 2 3 13 3 10 11 9 2 10 9 13 0 9 10 9 2
18 2 3 10 0 9 13 2 10 8 0 9 2 15 0 10 9 9 2
21 3 3 3 13 10 9 2 10 0 2 10 0 9 2 15 7 13 10 10 9 2
26 3 10 0 9 13 10 0 9 0 9 7 2 7 3 13 9 2 16 10 9 7 13 10 0 9 2
10 2 3 10 9 9 3 0 9 0 2
7 0 3 10 10 9 13 2
16 2 0 9 2 7 10 9 1 0 2 16 3 10 9 13 2
23 13 2 15 15 13 2 16 3 13 0 13 7 16 15 3 0 2 16 3 10 9 13 2
10 3 10 9 9 15 3 3 13 13 2
39 7 10 0 9 1 3 3 13 10 10 9 7 0 10 9 2 7 10 0 9 12 9 1 0 9 1 13 10 11 2 0 9 13 2 13 9 7 9 2
8 9 7 10 9 9 13 9 2
34 13 3 10 9 10 9 2 10 3 0 10 12 9 13 2 7 3 3 2 16 9 13 2 13 3 2 16 3 7 13 9 10 9 2
21 7 16 10 9 10 9 13 2 3 15 13 2 16 15 15 1 10 10 9 13 2
17 9 15 13 2 16 10 15 9 10 0 2 0 9 9 1 13 2
15 0 13 15 2 16 15 13 2 7 3 13 3 15 13 2
19 15 7 0 2 16 10 10 9 3 13 13 2 10 9 12 9 3 13 2
22 2 15 7 3 7 0 2 7 9 7 0 9 7 13 2 7 15 3 0 9 9 2
13 2 6 2 16 0 0 9 13 10 12 9 1 2
16 3 0 3 12 9 13 9 7 0 9 2 7 3 13 13 2
24 3 10 0 9 3 13 3 2 10 0 9 13 11 11 2 11 11 2 11 11 7 11 11 2
35 10 0 9 11 11 11 11 11 11 11 0 9 9 13 2 7 3 3 11 11 11 0 9 13 9 2 10 9 10 0 0 9 13 3 2
49 10 10 9 3 0 9 13 15 2 16 11 11 12 9 13 9 10 11 2 7 13 10 0 9 7 2 11 11 11 9 9 13 3 10 9 10 11 11 2 7 10 10 9 7 15 13 10 9 2
46 3 7 0 9 7 13 2 3 13 3 10 11 11 11 0 9 2 15 0 9 10 0 9 7 10 0 9 2 7 0 9 1 9 2 0 2 14 13 13 10 9 11 11 11 9 2
21 15 10 2 9 2 7 14 13 3 10 9 2 7 3 3 0 13 10 0 9 2
16 15 7 10 2 8 2 9 2 3 3 8 8 13 10 9 2
26 13 3 10 11 10 11 11 0 9 7 2 15 10 0 10 9 1 3 3 10 9 2 7 15 13 2
19 7 13 9 10 11 11 7 10 9 7 2 7 3 0 3 13 3 9 2
25 0 9 13 10 0 11 11 11 2 11 0 2 11 11 0 2 9 10 11 11 11 3 0 9 2
32 10 3 0 7 0 9 0 9 10 3 12 12 0 9 0 9 13 2 7 3 15 7 9 13 2 3 13 10 9 3 0 2
20 10 9 10 9 10 10 12 9 0 2 0 9 2 15 10 10 9 0 3 2
16 15 10 9 0 9 0 9 0 2 9 0 0 0 9 0 2
58 10 0 0 9 10 9 9 0 11 9 9 7 9 2 10 3 3 7 13 15 2 3 3 0 9 13 2 10 11 11 11 3 7 0 10 10 9 3 9 0 0 9 12 0 9 7 2 10 9 0 9 7 10 9 0 0 9 2
22 10 9 2 7 9 2 9 7 9 10 9 0 9 0 9 2 10 0 9 9 13 2
21 10 0 9 9 12 0 9 10 9 1 11 11 11 7 11 11 11 9 7 13 2
25 10 9 9 0 2 7 10 9 10 11 11 11 9 13 10 11 11 7 10 11 11 11 0 9 2
22 10 11 11 11 7 10 11 11 9 2 9 7 0 9 12 9 13 10 0 11 11 2
26 10 0 9 9 2 9 7 9 9 13 10 9 2 7 3 0 9 13 2 15 3 3 3 13 11 2
26 13 7 10 11 11 11 11 2 15 9 0 0 9 2 9 2 9 2 9 7 9 2 13 9 1 2
27 11 11 2 10 11 11 9 2 10 9 0 0 9 9 13 15 2 16 0 9 7 0 10 9 0 9 2
22 15 3 10 0 0 9 2 15 10 0 11 13 14 2 7 10 0 9 12 12 9 2
28 7 9 10 0 9 11 11 2 10 0 9 9 2 0 9 2 10 11 7 2 15 10 0 9 0 9 0 2
21 10 9 1 7 13 3 0 9 2 16 3 10 0 9 2 15 10 9 7 0 2
13 10 0 9 11 13 2 10 11 0 11 9 13 2
15 0 9 11 11 9 13 2 15 9 1 12 10 9 13 2
19 3 13 10 9 10 9 9 2 15 9 13 7 15 12 10 9 9 13 2
9 10 9 10 15 9 13 3 13 2
22 10 9 2 9 0 9 7 0 9 1 10 9 9 7 10 9 9 7 13 10 9 2
26 13 10 9 9 0 9 1 10 9 0 0 9 2 15 0 9 9 13 7 10 9 13 10 12 9 2
28 10 0 9 7 10 0 9 1 13 9 2 3 9 2 7 10 9 9 0 2 10 0 9 0 9 13 3 2
15 10 9 2 9 7 9 0 9 13 3 10 0 9 11 2
29 10 9 9 15 13 2 16 10 10 0 2 0 9 0 9 13 10 0 0 9 2 7 0 9 13 10 9 1 2
34 10 10 9 15 7 13 10 15 0 9 2 15 0 9 13 2 7 10 0 9 7 13 2 16 13 10 9 9 3 12 9 0 9 2
33 10 9 3 3 0 10 11 11 11 2 10 11 11 2 0 9 1 2 10 9 7 3 3 12 9 13 10 11 11 11 11 9 2
12 10 9 9 9 13 9 3 10 0 11 11 2
14 10 9 3 12 9 13 14 10 9 11 11 11 9 2
66 10 9 9 10 12 0 2 0 9 2 11 11 2 11 11 2 11 11 7 11 11 9 7 0 9 1 13 2 7 10 15 9 1 10 9 10 0 9 9 1 13 3 11 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 7 11 11 9 7 2
9 10 9 0 9 9 9 13 3 2
52 0 9 13 9 10 9 9 10 11 11 11 10 11 11 2 10 9 0 9 2 11 11 11 11 0 9 2 10 9 0 9 2 0 2 15 7 12 9 2 11 11 2 11 11 7 11 11 10 9 0 9 2
5 10 9 9 13 2
20 2 15 13 15 15 2 16 10 10 3 0 0 9 2 10 1 3 0 9 2
3 2 0 2
20 10 2 3 0 2 13 2 10 2 0 2 10 9 9 13 15 15 0 9 2
9 15 3 13 3 10 9 7 13 2
19 10 2 3 0 2 9 3 11 11 13 15 9 2 16 12 13 10 9 2
17 10 10 9 0 9 13 2 16 15 13 10 9 2 15 0 13 2
17 15 3 13 3 0 10 9 2 7 13 2 3 3 13 15 9 2
17 11 11 13 0 2 16 0 13 2 16 10 15 9 3 15 13 2
8 2 0 13 10 2 9 2 2
3 2 3 2
6 12 9 1 13 3 2
9 3 3 0 13 2 13 10 9 2
7 3 3 3 3 13 9 2
33 3 13 15 10 10 9 2 3 3 15 10 0 2 16 15 13 15 7 15 10 10 9 2 7 15 2 16 3 13 13 10 9 2
19 13 2 16 10 10 9 2 15 12 9 1 13 2 14 13 13 12 9 2
19 3 13 10 9 2 10 0 9 0 10 9 13 2 16 13 10 9 9 2
16 3 13 10 10 9 10 11 11 11 2 3 3 12 9 13 2
9 12 9 14 13 13 2 10 3 2
8 2 3 3 10 10 9 13 2
9 2 13 10 0 7 10 0 9 2
40 10 0 15 2 16 16 9 1 0 9 13 2 13 10 9 2 15 13 2 7 10 9 13 10 9 2 15 0 0 13 2 7 3 13 10 9 2 13 9 2
13 10 11 10 0 3 0 9 2 10 0 9 9 2
24 10 0 9 2 10 9 9 13 10 0 9 2 15 0 9 2 9 13 10 0 9 9 1 2
14 10 10 9 10 9 3 13 2 7 3 15 9 13 2
12 3 13 10 0 9 1 2 15 3 3 0 2
21 3 15 13 2 13 10 0 7 13 10 0 9 2 7 10 0 10 0 10 9 2
4 15 15 13 2
18 11 13 2 16 10 9 13 10 9 2 3 13 2 7 15 3 13 2
48 13 9 2 9 2 15 10 9 3 0 13 10 0 0 2 0 9 2 16 15 13 2 15 13 9 2 13 15 2 3 10 9 13 2 0 7 0 13 10 0 9 7 3 13 9 10 9 2
14 6 15 15 13 3 2 3 13 2 10 9 13 9 2
21 15 3 10 9 9 2 10 0 9 0 0 9 13 2 7 0 13 7 0 13 2
28 3 13 10 10 9 2 16 13 3 10 9 2 3 13 15 2 16 2 13 2 2 2 3 13 13 7 13 2
19 2 10 9 0 0 2 10 9 13 3 10 9 9 2 15 7 3 0 2
13 2 3 0 10 9 2 10 9 13 10 0 9 2
15 16 10 9 2 10 9 2 7 10 9 13 3 10 9 2
7 10 9 0 9 10 9 2
23 10 9 1 10 9 3 13 3 10 9 2 10 0 9 3 9 13 2 7 3 13 13 2
12 2 10 10 9 3 0 2 7 0 2 0 2
13 2 11 1 10 9 0 9 10 9 9 10 9 2
8 10 9 2 10 0 13 13 2
14 16 10 0 0 13 10 9 2 15 7 0 0 13 2
9 2 12 9 0 13 3 10 9 2
11 2 11 11 10 9 2 15 3 13 15 2
8 3 7 9 13 9 10 9 2
12 15 13 10 9 2 16 10 9 3 3 13 2
5 10 9 3 13 2
22 3 0 9 13 10 11 2 3 0 7 0 2 13 2 3 13 3 15 10 15 9 2
13 0 7 9 13 2 13 2 3 13 3 12 9 2
6 2 3 13 13 9 2
17 2 10 9 13 13 7 3 13 2 7 10 10 9 3 3 13 2
11 13 13 10 9 2 7 13 2 3 13 2
10 2 10 11 9 7 10 0 9 13 2
9 2 15 10 9 2 15 0 13 2
12 10 9 11 13 2 15 15 3 11 13 13 2
5 15 13 10 11 2
7 15 13 2 15 10 9 2
10 10 0 9 10 9 2 15 0 13 2
5 10 15 9 13 2
16 0 9 13 3 3 3 10 11 11 11 11 10 0 11 11 2
18 10 9 0 9 0 9 10 3 12 2 0 9 2 13 3 10 9 2
13 10 9 7 3 0 11 11 3 0 9 11 13 2
18 12 13 10 3 3 3 0 11 11 11 2 7 3 12 9 10 9 2
20 0 0 9 3 13 9 2 3 3 13 9 9 1 12 9 1 9 10 9 2
6 10 9 0 9 13 2
19 10 0 9 10 1 10 0 9 1 11 0 0 9 11 11 0 9 13 2
20 12 15 13 10 9 11 11 11 0 9 10 9 9 13 11 11 11 0 9 2
19 10 9 0 9 13 11 11 7 2 15 3 12 9 0 9 10 11 11 2
16 9 2 9 7 13 2 12 7 12 1 7 10 9 9 13 2
16 9 13 3 10 0 9 2 7 10 9 0 9 3 13 9 2
28 9 2 10 9 0 0 9 15 10 0 9 7 13 2 3 7 3 11 11 11 11 11 13 15 10 0 9 2
33 11 11 7 3 0 7 0 9 11 2 0 2 16 3 10 0 9 0 0 11 11 11 0 9 0 0 2 7 0 0 9 13 2
26 12 13 10 0 9 2 10 9 7 9 13 2 7 0 9 10 11 11 11 13 2 3 3 7 13 2
11 13 10 9 2 7 0 10 9 13 15 2
17 13 7 0 9 3 13 11 11 9 2 12 2 11 11 0 9 2
21 10 9 12 0 0 9 10 11 11 11 9 13 3 2 7 10 0 9 13 3 2
9 2 9 10 9 9 13 3 2 2
23 10 0 9 9 9 13 10 12 9 0 9 2 7 10 9 9 11 10 9 13 10 9 2
20 10 11 11 10 9 9 0 9 13 14 10 9 9 0 7 9 0 9 9 2
12 10 9 12 0 9 9 13 9 10 9 9 2
11 0 9 13 3 10 9 9 10 10 9 2
8 15 3 2 15 10 9 3 2
8 2 0 7 13 2 3 2 2
15 10 15 9 9 2 11 2 10 15 9 9 2 11 11 2
31 3 0 2 7 11 11 11 0 9 3 3 3 3 13 9 10 9 2 7 9 3 3 13 14 9 10 11 11 11 9 2
29 10 10 0 9 2 15 10 9 0 9 0 9 0 9 7 0 9 13 2 3 10 9 9 13 10 0 9 9 2
36 3 15 13 12 10 12 2 3 15 7 2 16 11 13 10 9 2 16 3 13 2 16 15 2 15 10 9 10 9 3 13 13 10 9 9 2
38 10 0 0 9 9 0 2 0 9 13 10 9 2 15 10 9 1 13 14 10 9 2 10 0 9 9 2 7 15 9 9 3 7 3 10 9 13 2
56 9 10 9 2 7 9 9 7 0 9 10 9 9 0 9 2 11 0 9 10 9 1 2 7 3 0 10 0 9 9 2 11 9 2 15 10 9 11 10 9 2 10 9 7 10 9 0 9 2 10 0 9 13 10 9 2
25 10 0 0 9 1 10 0 9 9 2 16 11 11 0 0 9 11 13 2 10 9 2 0 9 2
62 10 11 9 1 3 10 0 9 13 10 0 2 7 15 7 0 2 16 11 11 11 11 0 0 9 9 1 11 11 0 10 9 3 9 13 2 11 11 0 9 2 0 9 2 6 7 6 15 2 16 0 7 0 2 13 10 0 0 9 0 9 2
34 10 0 9 2 11 11 2 11 11 2 9 0 9 11 3 3 10 9 2 7 9 2 9 3 3 13 7 15 2 7 10 9 0 2
36 10 0 9 0 9 9 3 10 7 15 10 9 2 0 9 13 10 9 3 15 3 2 16 10 9 9 3 3 13 3 9 10 0 9 1 2
43 16 13 9 10 9 2 13 2 13 2 13 2 2 7 10 0 9 7 15 2 16 3 9 13 2 12 0 9 1 10 0 11 11 7 10 9 11 11 0 3 10 9 2
43 10 9 3 0 2 7 6 3 3 13 10 9 15 2 16 10 0 0 2 0 2 0 2 9 2 10 0 11 9 2 7 15 7 3 10 11 0 9 10 0 9 9 2
36 10 9 0 9 0 9 13 10 9 2 7 15 2 13 3 2 3 10 10 9 13 2 15 10 0 9 0 9 0 13 10 0 9 10 9 2
36 13 7 9 9 7 9 2 9 7 9 2 7 3 10 9 9 7 0 9 13 2 7 3 3 11 10 9 7 9 13 2 16 13 10 9 2
7 16 3 0 0 3 13 2
16 11 11 11 11 11 11 9 0 9 13 9 10 11 11 9 2
57 10 9 10 12 9 9 7 9 12 9 13 3 2 11 11 11 9 7 11 11 9 13 0 9 2 3 11 11 11 0 9 13 3 10 9 2 7 10 3 12 9 10 0 9 0 11 11 9 13 3 10 15 7 10 9 1 2
46 10 9 9 1 10 9 3 10 0 9 13 2 10 9 3 10 0 9 2 10 0 9 2 10 9 9 2 10 0 0 9 7 9 2 10 12 9 9 2 10 0 9 9 13 15 2
14 10 9 0 0 2 9 2 0 10 0 9 3 13 2
13 10 12 9 0 9 9 10 9 10 9 7 13 2
23 3 3 11 7 11 7 12 0 9 13 9 1 2 7 10 9 0 9 12 9 13 3 2
31 10 0 9 9 9 10 11 11 13 9 10 9 12 12 0 9 10 9 2 3 11 0 10 0 9 9 13 14 10 9 2
20 10 0 9 9 0 9 13 3 15 2 16 0 10 9 9 13 10 9 9 2
27 10 0 9 0 9 3 3 13 2 7 9 1 10 0 0 9 3 13 15 2 16 13 14 11 11 9 2
20 10 9 0 9 0 9 0 9 3 3 3 13 2 7 15 3 9 7 13 2
25 10 0 9 9 13 15 2 16 3 13 3 9 11 11 0 9 2 15 0 9 0 9 9 13 2
22 10 0 9 3 10 0 9 9 13 2 15 10 9 9 9 0 13 0 9 9 7 2
20 10 0 9 10 9 9 0 13 2 16 10 0 9 3 10 9 9 13 0 2
10 10 0 9 9 15 10 9 13 9 2
25 16 15 3 0 2 10 9 10 9 9 0 12 9 1 10 9 13 13 10 0 9 0 9 9 2
7 10 9 3 12 9 13 2
25 16 10 0 9 9 15 1 7 13 2 10 9 13 10 9 2 16 3 13 14 10 9 0 9 2
49 11 11 2 10 0 11 11 11 2 11 2 9 9 10 0 9 15 1 15 13 2 16 10 9 0 9 2 13 2 15 9 1 10 9 13 2 7 9 0 9 3 13 14 15 10 0 9 2 2
35 10 0 9 9 10 0 9 1 13 2 15 1 15 3 2 16 10 9 3 13 9 10 9 9 2 7 3 0 13 10 0 9 9 7 2
26 10 9 1 10 9 9 0 9 0 12 9 1 0 9 13 13 2 7 10 0 9 3 3 13 9 2
14 0 13 10 0 0 9 0 9 10 11 0 0 9 2
18 10 11 0 0 9 0 9 3 15 13 2 16 10 9 13 11 9 2
27 10 9 1 10 9 9 9 3 3 2 3 12 9 9 1 2 13 14 2 15 0 9 7 9 13 9 2
30 10 11 11 0 0 9 0 9 9 11 11 11 9 15 13 9 2 16 2 3 3 10 0 9 3 13 2 10 9 2
24 10 9 13 11 11 0 9 2 15 13 2 10 9 1 13 15 2 16 13 14 11 11 9 2
25 10 11 11 0 9 3 13 2 16 10 11 11 0 9 13 11 9 9 2 7 10 9 13 9 2
42 11 11 0 7 11 11 0 9 9 11 13 10 0 11 12 9 2 10 11 11 7 10 11 11 0 2 3 0 7 9 1 10 9 0 2 9 0 0 9 0 9 2
61 10 9 1 10 0 9 0 9 2 12 2 7 12 0 9 13 10 11 11 11 10 10 12 12 9 0 0 9 2 15 1 11 10 0 11 12 9 0 9 1 2 0 9 1 3 13 0 13 11 10 3 0 0 9 0 9 0 12 9 9 2
10 11 3 3 13 3 10 0 9 9 2
18 10 0 0 7 10 0 0 9 9 1 3 13 13 10 9 0 9 2
30 11 11 7 11 11 7 3 12 9 2 0 10 0 9 1 3 9 13 2 15 9 12 9 1 9 13 10 9 9 2
32 13 10 9 2 10 9 9 1 10 0 9 0 10 0 9 9 2 15 0 13 11 2 16 10 9 3 10 12 9 7 13 2
25 2 10 12 9 15 13 10 9 2 7 10 0 0 9 1 13 9 2 2 13 3 11 0 9 2
22 11 11 2 10 0 9 9 9 13 2 13 10 11 9 7 9 0 0 9 0 9 2
10 11 15 10 11 0 0 0 9 13 2
14 10 11 0 0 9 3 13 10 0 0 9 9 9 2
16 11 13 2 16 3 12 0 9 13 11 2 7 15 0 0 2
7 2 12 12 9 13 9 2
15 3 13 10 0 9 2 2 2 13 3 10 9 10 9 2
32 9 0 9 9 3 9 13 10 0 9 11 0 9 1 2 10 0 9 9 2 12 9 13 2 13 9 10 11 0 0 9 2
19 10 11 0 9 0 9 1 10 9 10 3 9 0 11 7 11 1 13 2
11 10 9 1 10 9 10 0 9 13 9 2
38 10 0 0 9 0 9 1 10 0 9 9 3 13 10 12 9 2 15 10 11 11 7 10 0 9 1 0 9 9 9 13 10 0 0 2 0 9 2
17 10 0 9 3 13 15 2 16 10 9 3 3 13 14 0 9 2
19 11 1 11 9 13 3 10 2 11 11 11 2 0 9 9 1 0 9 2
7 3 12 0 9 13 11 2
31 11 11 9 9 13 2 10 9 3 13 10 9 10 10 9 2 16 2 3 15 15 9 2 16 10 9 13 10 9 2 2
19 0 0 9 7 10 0 9 9 13 11 11 3 0 2 0 0 0 9 2
15 10 0 7 10 0 0 9 9 3 3 9 11 13 9 2
22 10 9 9 0 9 9 15 13 2 16 0 0 9 13 10 0 9 0 0 9 9 2
11 11 11 9 0 9 3 12 9 13 11 2
13 11 11 10 10 9 3 2 3 9 13 3 11 2
21 10 12 9 9 0 0 9 2 3 10 0 0 9 7 10 9 2 3 0 13 2
26 10 0 9 9 0 9 2 10 0 9 9 0 9 2 3 7 11 11 0 9 13 3 0 9 11 2
23 11 13 15 2 16 10 0 9 0 9 2 9 10 0 9 1 7 0 13 13 7 13 2
33 11 11 3 0 0 0 9 9 2 16 9 2 11 11 9 13 0 0 9 7 10 0 9 2 13 9 11 11 2 10 11 9 2
22 10 9 3 9 13 10 0 9 2 10 0 9 2 10 0 9 7 10 0 9 9 2
28 16 10 9 15 13 9 10 12 9 1 2 10 9 10 9 1 0 9 13 10 9 9 2 7 3 9 7 2
15 10 0 9 2 10 0 0 9 10 9 10 0 9 9 2
20 11 3 12 12 0 9 9 13 10 9 10 0 0 0 9 0 2 0 9 2
15 10 9 10 9 13 2 16 0 9 13 3 10 9 9 2
6 10 9 9 0 9 9
17 10 0 0 9 11 11 3 13 13 10 11 0 0 9 9 9 2
19 10 0 7 0 9 0 0 0 9 9 11 9 13 11 0 9 0 9 2
26 3 11 11 13 2 10 0 9 3 10 9 13 10 0 9 10 0 9 2 15 10 11 11 9 9 2
9 10 9 9 0 9 13 10 9 2
14 10 9 3 13 2 10 9 3 0 0 9 13 9 2
11 10 0 9 7 3 15 13 10 0 9 2
20 3 3 0 2 16 10 9 10 9 2 10 9 2 15 9 0 9 9 13 2
10 10 0 0 9 9 3 13 11 9 2
8 11 9 7 0 9 11 1 2
26 3 3 0 13 10 0 0 9 2 7 9 9 13 10 9 0 7 0 0 9 2 13 3 11 11 2
18 10 0 9 0 9 13 11 2 7 15 0 10 3 3 3 13 9 2
21 11 11 3 3 13 2 0 11 13 2 16 10 0 9 3 13 0 10 0 9 2
6 11 3 13 10 9 2
21 10 0 9 0 9 13 2 16 10 0 9 3 0 13 11 2 3 15 11 13 2
16 10 9 1 10 0 9 0 7 0 9 0 10 9 7 9 2
28 11 11 7 0 13 10 10 0 9 2 15 1 10 0 9 0 13 3 11 7 10 9 3 0 9 13 9 2
12 2 15 3 13 3 10 9 2 2 13 3 2
19 11 11 0 9 13 2 10 0 9 13 2 16 0 9 9 13 7 13 2
35 2 0 2 16 10 11 12 9 3 0 9 2 10 10 0 0 9 2 13 10 0 0 9 2 3 0 9 13 10 9 1 2 2 13 2
27 10 0 9 9 7 10 0 9 3 0 13 11 9 2 7 10 9 3 0 0 9 9 0 13 10 9 2
13 0 9 1 10 0 9 9 10 0 9 12 13 2
26 10 0 9 7 0 9 11 13 10 11 0 0 9 0 11 11 2 7 13 15 2 16 9 13 11 2
16 11 11 15 7 13 2 16 11 9 9 0 9 13 10 9 2
27 10 0 0 9 3 3 15 13 10 0 9 2 11 0 0 2 3 10 9 0 9 3 3 13 13 15 2
23 11 10 0 0 0 9 3 16 2 7 13 15 2 16 10 11 9 13 10 9 0 9 2
26 10 0 9 9 13 10 10 0 9 2 15 3 13 9 10 9 2 7 13 10 9 10 0 9 1 2
26 11 11 13 2 16 10 0 9 2 15 0 13 10 0 0 9 0 0 9 2 3 13 10 0 9 2
22 11 3 3 13 3 0 11 9 2 15 3 2 16 10 9 7 10 9 14 4 13 2
37 3 13 2 16 10 9 2 0 9 2 13 3 0 9 2 7 10 9 3 13 13 10 0 9 2 7 10 0 9 2 15 3 4 13 15 2 2
55 10 0 9 2 15 9 9 11 11 13 2 10 0 9 0 0 9 1 3 13 13 10 10 0 9 2 15 10 11 0 9 0 0 9 13 2 9 13 2 7 3 10 0 9 9 2 11 11 0 0 2 0 9 13 2
28 3 2 10 0 2 0 9 2 0 9 3 2 15 0 2 10 9 13 11 11 9 2 10 0 9 0 9 2
51 3 7 11 11 11 9 2 11 11 0 9 2 7 10 9 7 10 11 9 9 2 11 11 0 13 9 2 3 9 9 13 2 10 0 0 2 2 3 10 10 9 11 13 2 2 7 9 13 3 15 2
25 11 9 7 13 10 9 2 7 11 11 0 9 7 13 10 0 9 9 2 9 9 2 11 11 2
43 10 0 9 2 7 11 1 2 3 13 2 10 9 7 2 15 13 9 2 16 12 9 11 9 3 0 13 10 10 0 7 0 9 10 9 2 15 11 3 0 9 13 2
38 11 7 0 13 2 16 0 9 2 11 11 1 2 10 9 7 9 0 9 2 7 10 12 9 0 0 9 9 1 2 7 10 0 9 9 13 13 2
29 11 15 13 10 9 2 16 10 0 9 9 0 0 7 0 9 0 9 13 16 2 7 3 3 10 12 9 9 2
27 10 9 1 3 3 13 7 10 0 9 2 7 10 0 11 11 9 10 0 2 7 15 0 2 9 9 2
28 3 13 10 9 9 10 9 9 2 7 15 7 13 2 10 0 11 9 9 3 3 13 10 9 10 0 9 2
11 16 15 0 13 2 3 10 9 9 1 2
19 11 11 15 13 2 16 10 0 9 0 0 11 9 2 11 11 10 9 2
15 11 3 3 10 9 1 13 11 1 2 15 3 13 15 2
11 0 9 0 0 9 13 2 0 13 15 2
32 11 10 10 9 13 2 16 10 9 1 10 0 9 9 13 2 7 0 13 11 9 10 10 9 1 2 15 0 9 1 13 2
19 15 7 13 10 0 9 2 16 10 9 1 9 13 4 0 0 9 9 2
13 15 7 15 3 13 2 3 15 10 9 9 3 2
34 0 9 13 10 9 10 11 9 0 9 2 0 9 13 11 2 2 15 13 10 0 0 9 1 0 9 9 2 15 10 9 9 13 2
37 3 13 15 3 10 9 2 3 13 3 3 10 0 9 10 9 0 0 9 15 2 16 10 0 0 11 11 11 11 3 13 10 9 10 9 9 2
15 11 11 3 13 2 7 15 13 2 0 13 3 0 13 2
43 7 3 15 13 10 9 2 3 10 11 11 0 9 13 2 3 11 2 10 0 9 9 7 11 11 2 15 0 15 13 3 9 2 12 9 1 0 13 10 9 0 9 2
33 10 0 11 11 11 9 9 0 13 10 10 9 2 15 10 9 9 13 9 9 3 2 16 13 10 0 9 10 0 0 9 9 2
33 10 12 9 0 2 12 9 0 9 9 1 15 9 7 10 0 0 9 13 2 7 10 0 0 9 2 10 1 11 11 9 7 2
13 10 11 9 1 10 9 9 12 12 0 9 13 2
17 10 11 0 2 0 9 2 9 9 13 9 11 11 11 0 9 2
35 10 9 15 7 13 2 16 12 12 9 2 3 12 12 9 2 13 10 10 12 9 10 9 2 15 10 10 13 10 0 9 3 0 9 2
18 10 9 0 0 9 13 3 10 0 0 9 7 10 11 11 9 7 2
28 10 11 3 10 9 9 9 13 9 9 2 15 1 10 0 9 10 0 9 10 0 0 9 0 3 0 9 2
15 10 0 9 0 9 13 10 0 9 7 10 9 9 9 2
24 11 11 9 15 13 2 16 16 3 13 0 9 10 9 2 3 10 9 10 0 9 9 13 2
23 10 11 9 3 10 0 0 9 3 13 2 16 9 13 13 9 10 9 9 1 0 9 2
54 10 0 9 11 0 9 1 0 9 1 10 9 0 9 0 9 9 10 0 9 1 0 2 3 12 2 9 10 9 7 13 10 0 9 2 7 3 4 13 0 9 2 15 0 13 10 0 9 9 0 9 0 9 2
38 10 12 0 9 1 2 12 9 9 1 0 9 1 10 9 13 2 13 3 9 15 2 16 10 0 9 10 9 9 1 7 3 13 10 9 0 9 2
41 10 9 10 9 7 10 9 10 9 7 13 10 10 9 2 7 10 9 0 9 13 10 9 9 2 15 9 7 2 2 16 10 0 9 9 3 13 9 10 9 2
14 15 0 15 13 2 16 10 0 9 13 10 0 9 2
40 11 11 11 9 3 0 2 3 0 9 7 13 10 0 9 9 10 0 9 0 0 9 2 15 3 10 9 2 16 10 9 9 0 13 14 3 0 9 9 2
35 10 9 9 9 10 11 0 2 8 8 2 9 1 9 13 3 10 9 2 15 13 9 7 9 10 0 9 2 15 10 9 2 9 1 2
58 10 9 15 0 10 0 0 9 9 2 11 11 0 9 13 2 15 13 2 16 10 0 0 9 2 10 9 7 13 7 13 10 9 0 0 9 2 7 3 13 3 0 9 2 15 1 10 0 9 10 9 0 0 9 9 13 2 2
24 12 0 0 0 9 10 9 9 0 9 13 3 10 0 0 9 2 13 13 10 0 0 9 2
9 3 10 9 13 10 9 0 9 2
32 10 9 9 1 0 13 10 11 0 0 9 2 9 2 2 7 10 9 0 9 16 13 2 7 10 0 9 3 0 13 15 2
18 10 11 11 11 0 9 1 10 10 9 13 13 10 9 0 0 9 2
16 11 11 13 9 2 15 2 11 2 9 13 10 0 9 9 2
12 10 0 9 12 10 0 0 9 0 9 13 2
34 10 10 12 9 2 15 9 7 13 2 16 13 10 9 2 7 13 10 3 12 0 9 2 7 9 10 9 3 3 13 3 10 9 2
18 11 15 13 11 2 16 10 11 15 9 0 9 9 13 3 15 11 2
18 13 15 2 16 9 2 11 11 11 9 13 15 2 7 9 13 13 2
24 10 9 3 13 10 0 0 9 2 15 10 9 9 13 3 15 2 7 13 11 2 9 13 2
11 2 11 2 3 13 15 2 0 13 13 2
27 3 13 10 11 9 10 0 0 0 9 1 10 9 0 0 9 2 7 3 10 9 9 10 0 9 7 2
29 10 0 9 10 9 13 3 2 10 11 11 9 1 3 2 15 3 13 15 2 16 12 9 9 10 0 9 13 2
21 10 9 15 0 13 3 2 16 10 9 10 9 13 10 0 9 9 0 10 9 2
18 10 9 2 3 10 12 0 11 11 9 13 2 10 9 12 9 13 2
26 10 9 9 2 10 9 12 0 9 15 13 2 16 9 3 13 2 3 13 2 7 10 9 13 9 2
17 10 9 10 13 10 9 2 15 0 7 0 2 0 2 9 13 2
25 3 3 12 12 9 13 10 0 9 2 10 9 2 13 9 10 11 11 9 10 11 11 9 3 2
12 3 0 9 3 13 14 15 10 0 9 1 2
20 7 3 10 0 9 2 12 12 12 9 7 9 13 14 10 9 9 0 9 2
18 10 9 9 2 7 10 0 9 9 1 10 9 12 12 9 13 14 2
7 15 3 3 12 12 13 2
13 10 9 0 0 13 10 11 9 2 13 10 9 2
12 10 10 9 12 7 12 1 13 10 9 9 2
45 3 10 9 13 2 10 11 11 11 9 2 3 10 10 0 7 0 9 2 3 3 0 10 9 9 2 0 9 13 10 9 9 2 7 10 10 9 3 10 0 9 13 10 9 2
27 15 0 10 9 2 9 2 3 7 11 2 7 3 15 11 3 0 9 2 3 10 9 9 12 9 9 2
26 10 9 1 12 9 2 3 10 12 7 12 9 0 3 2 12 12 0 9 7 12 12 9 13 9 2
13 11 15 1 3 10 9 13 3 10 9 0 9 2
15 3 0 10 9 11 7 2 3 3 0 9 13 10 9 2
10 11 12 12 9 13 12 12 9 9 2
9 10 9 3 3 13 10 0 9 2
19 10 0 9 3 10 0 9 0 0 9 13 10 0 9 9 7 10 9 2
24 3 3 10 0 9 0 9 13 2 7 10 0 9 7 10 9 9 7 0 9 13 10 9 2
12 10 9 0 9 13 10 9 0 9 10 9 2
19 3 9 11 11 2 10 0 9 9 10 11 13 2 13 10 0 9 9 2
30 3 0 9 7 9 13 3 2 16 10 0 9 7 10 9 9 2 7 10 9 0 9 3 13 9 2 13 10 9 2
8 10 9 3 13 3 0 9 2
13 3 2 9 2 0 10 9 2 7 10 0 9 2
19 10 11 11 0 0 7 0 0 9 10 9 7 0 13 10 0 9 9 2
16 3 13 7 7 10 0 2 7 3 10 9 0 0 9 7 2
12 9 11 11 9 15 13 2 16 0 9 13 2
20 9 1 0 9 7 3 9 9 13 3 2 3 10 9 0 9 0 9 13 2
33 10 0 9 9 3 3 13 0 10 9 0 9 0 0 9 2 15 7 3 3 0 2 16 0 0 9 13 10 9 10 9 9 2
15 10 9 10 9 9 3 10 9 3 13 2 9 3 13 2
18 10 9 0 9 13 2 15 3 13 0 10 9 2 13 11 11 9 2
19 10 0 0 9 3 15 13 2 16 10 0 9 9 9 7 13 10 9 2
15 3 10 9 10 9 3 3 0 7 3 3 13 9 13 2
38 10 0 0 9 2 3 13 2 3 13 13 2 16 10 9 7 10 9 0 9 2 7 10 2 9 7 9 9 0 9 9 7 13 3 10 9 9 2
62 10 9 2 10 9 7 10 9 0 2 0 2 12 2 12 2 12 0 2 7 10 3 0 0 0 9 2 16 0 10 9 2 9 0 2 0 9 13 10 0 9 2 15 7 10 0 9 9 3 13 2 7 0 3 13 2 0 10 9 9 13 2
13 7 10 9 0 9 2 16 15 10 0 9 13 2
10 10 0 9 9 10 0 9 0 13 2
18 3 3 10 9 13 0 9 2 3 3 10 0 9 1 13 10 9 2
15 9 3 3 13 3 10 9 10 9 2 16 10 0 9 2
12 0 9 1 10 9 10 9 9 13 10 9 2
18 10 0 9 7 0 13 0 9 2 7 0 9 3 3 13 10 9 2
21 3 11 11 9 2 10 9 9 9 13 2 0 9 2 13 3 2 10 0 9 2
17 2 10 9 0 9 3 3 0 9 13 2 7 9 3 0 13 2
24 15 7 3 3 10 0 9 2 3 10 9 3 13 7 10 9 7 9 13 2 13 10 9 2
13 2 3 10 9 13 10 9 10 0 9 0 9 2
10 0 9 13 3 10 9 0 0 9 2
26 15 15 0 3 2 16 10 0 9 15 13 10 9 2 15 3 13 2 7 9 13 10 9 0 9 2
30 10 0 9 9 12 9 1 0 9 13 2 3 10 9 15 13 2 16 3 2 3 9 3 13 0 10 9 0 9 2
9 11 3 2 11 3 2 11 3 2
30 10 0 2 0 2 9 0 9 2 11 11 9 9 11 11 13 2 7 6 9 7 2 7 0 9 13 0 0 9 2
15 3 3 13 9 3 2 7 9 9 11 0 11 11 9 2
37 10 9 3 13 2 3 7 9 3 11 2 7 13 13 10 9 0 2 0 9 2 7 9 1 10 9 2 7 3 12 10 0 9 2 11 1 2
27 9 13 11 11 10 10 11 0 9 2 15 10 11 11 0 0 9 0 9 0 2 15 0 9 9 13 2
28 3 3 13 3 10 9 2 3 10 10 9 13 10 9 1 2 15 10 9 10 9 10 15 9 7 3 13 2
22 2 3 10 15 9 13 10 0 12 2 13 10 9 0 0 0 2 9 7 9 9 2
15 2 13 11 11 2 7 10 10 9 12 9 13 10 9 2
23 3 3 13 9 2 3 13 9 2 7 3 13 7 2 7 9 0 10 9 13 10 9 2
5 16 3 13 4 2
12 2 7 3 13 3 0 3 13 10 9 9 2
15 2 10 0 9 2 7 3 3 13 2 7 3 3 13 2
21 3 16 10 9 0 13 10 12 9 9 2 3 16 15 13 2 15 13 2 11 2
13 15 3 12 2 11 13 3 2 0 2 0 9 2
18 2 15 0 2 16 3 3 13 9 13 9 1 2 0 9 3 13 2
23 3 15 9 13 7 3 13 0 0 9 2 10 3 0 11 11 11 9 0 9 15 13 2
7 2 3 15 10 0 9 2
19 15 7 10 9 9 13 10 9 2 7 3 3 13 14 10 15 0 9 2
27 3 11 11 2 10 11 11 9 13 2 16 15 3 13 10 9 2 7 3 10 0 0 9 9 9 13 2
13 2 9 13 2 16 9 9 3 10 9 10 9 2
7 2 3 3 13 15 7 2
17 2 15 7 13 2 16 3 13 0 10 11 11 0 2 0 9 2
8 2 3 3 2 9 13 3 2
22 7 15 0 13 2 16 9 13 2 3 3 13 11 11 11 2 10 9 2 11 2 2
3 2 3 2
14 2 3 12 9 2 16 10 9 7 3 13 7 13 2
7 2 3 3 13 10 9 2
11 2 0 9 11 13 11 11 0 0 9 2
18 10 10 9 13 3 10 0 11 2 11 7 2 7 10 0 11 11 2
25 2 10 9 13 0 0 0 9 2 10 0 0 9 2 3 15 13 9 2 12 0 9 11 1 2
3 2 0 2
3 3 10 2
5 2 10 9 13 2
24 2 0 2 7 3 9 3 11 2 7 9 9 13 13 2 7 13 10 9 2 11 2 11 2
17 15 3 9 7 13 10 9 2 3 7 15 2 7 10 11 7 2
50 10 11 0 0 9 9 0 9 13 2 10 0 9 9 0 9 9 9 13 10 9 1 2 7 9 9 10 9 13 3 10 0 9 2 13 3 11 11 2 10 9 9 10 11 0 7 9 0 9 2
14 11 13 15 7 2 16 10 9 0 9 12 12 9 2
20 13 2 15 10 0 9 1 0 10 9 10 11 2 7 9 7 9 7 13 2
12 15 13 2 7 0 2 16 3 13 15 13 2
15 13 2 3 12 9 0 10 9 2 15 13 3 3 13 2
30 10 9 10 0 9 13 11 11 2 10 11 0 9 2 15 10 1 13 2 10 9 3 0 0 9 9 0 9 13 2
22 10 9 13 10 10 0 9 2 15 10 11 11 11 0 0 12 0 0 9 12 13 2
25 11 11 2 10 9 0 9 12 13 3 9 2 7 10 12 0 9 12 9 1 13 0 0 9 2
19 10 9 9 12 1 9 2 12 11 11 7 11 11 1 7 13 0 9 2
23 12 11 1 0 0 9 1 2 12 9 9 2 7 10 9 2 7 10 0 9 7 13 2
13 0 13 3 10 9 2 10 9 10 9 3 13 2
31 10 0 0 9 12 9 13 3 2 3 11 9 13 2 0 9 13 2 7 10 0 0 2 12 0 9 12 9 0 13 2
19 9 10 0 0 11 3 13 13 10 0 9 0 9 2 12 9 0 9 2
27 10 11 11 13 10 11 9 9 0 9 9 10 9 2 11 2 11 2 11 2 11 2 11 13 10 9 2
17 10 0 0 9 10 0 9 13 2 3 15 15 3 13 10 9 2
17 10 11 11 2 11 11 2 11 11 2 11 11 9 9 10 0 2
23 10 0 9 9 0 9 7 10 0 9 13 2 11 2 11 2 11 7 11 13 3 9 2
17 0 9 13 3 10 9 2 11 2 11 2 11 2 11 10 9 2
28 10 9 10 3 0 9 11 0 11 10 2 9 2 2 10 9 11 2 11 2 11 2 11 9 13 9 9 2
27 10 9 13 2 10 0 2 9 2 9 9 13 10 9 2 10 9 11 2 11 2 11 2 11 9 13 2
9 10 0 0 9 13 11 7 11 2
16 11 3 2 13 2 9 10 0 9 2 11 9 13 0 9 2
21 10 9 9 3 13 11 2 15 10 11 7 11 11 0 9 3 10 0 9 13 2
19 10 9 11 10 0 2 10 9 11 2 10 9 11 2 11 9 7 11 2
33 10 9 10 9 9 12 0 9 7 13 2 10 2 9 2 9 11 2 11 7 11 13 2 3 10 2 9 2 9 11 7 11 2
16 11 11 2 11 11 7 11 11 10 9 3 10 0 10 9 2
14 10 0 9 10 9 9 0 13 10 0 9 0 9 2
27 10 12 9 0 9 1 3 10 9 9 1 3 13 10 11 11 9 2 15 9 9 7 9 13 10 9 2
26 10 9 7 10 9 2 7 11 9 9 1 7 13 0 9 13 2 13 9 10 0 9 10 11 9 2
42 3 10 10 9 13 9 9 13 10 0 9 10 0 9 2 15 3 13 10 0 9 9 0 0 0 0 0 9 2 7 13 10 9 0 9 2 15 9 13 10 9 2
17 11 10 9 3 13 2 7 15 10 9 1 7 13 13 0 9 2
44 11 11 2 10 11 0 9 9 13 2 3 13 10 10 9 2 2 3 9 13 3 10 11 2 7 10 9 10 10 9 13 2 16 9 9 3 13 13 10 9 2 13 11 2
10 2 10 0 9 10 11 9 13 13 2
20 9 12 9 7 9 13 13 2 15 15 1 13 3 12 7 12 10 0 9 2
43 11 11 2 10 11 0 9 11 0 9 13 10 9 2 2 10 11 15 13 2 16 10 9 1 13 10 0 9 2 7 0 9 3 10 9 1 13 15 13 2 13 3 2
16 2 0 0 13 2 16 3 10 0 9 10 9 13 10 9 2
16 10 0 0 9 9 15 9 13 2 7 15 3 13 3 0 2
16 3 10 11 15 13 4 13 2 3 10 9 9 0 9 13 2
18 11 11 9 1 10 0 0 9 1 0 13 10 0 9 9 3 13 2
8 2 9 10 9 3 13 9 2
18 9 13 2 16 9 0 0 9 13 3 10 0 9 2 13 10 9 2
22 11 11 2 10 11 9 15 13 2 16 10 9 9 0 9 13 11 2 10 0 9 2
16 2 13 9 10 0 9 9 2 16 3 0 10 9 2 13 2
18 2 10 9 1 3 13 0 0 9 13 2 16 15 13 13 10 9 2
24 9 9 10 11 11 9 13 4 9 10 9 2 7 10 0 9 1 10 9 7 3 13 13 2
8 10 0 9 3 12 13 13 2
20 11 11 2 10 11 9 1 10 0 9 9 3 12 12 9 9 13 10 9 2
13 2 10 9 0 9 13 2 9 10 0 9 0 2
16 15 15 10 0 2 16 0 9 2 0 0 9 13 10 9 2
12 12 9 9 13 10 9 11 11 0 9 9 2
37 10 9 9 10 11 0 9 0 9 13 10 11 2 10 9 2 7 10 11 11 0 9 0 7 13 2 2 3 10 11 11 3 9 13 10 11 2
18 10 9 9 13 10 9 9 2 10 11 9 9 13 10 0 11 11 2
13 10 10 9 13 10 9 0 9 2 11 11 9 2
16 10 9 7 10 9 9 9 3 2 0 9 9 1 13 9 2
37 9 9 3 13 15 11 9 10 11 7 10 11 11 2 15 3 10 0 11 9 13 9 2 10 11 12 0 9 9 0 9 11 0 9 13 3 2
35 15 10 12 9 9 3 3 0 0 2 7 10 11 11 7 11 11 3 10 11 9 2 3 11 0 3 3 9 13 10 2 11 11 2 2
23 10 0 9 7 15 13 10 9 2 3 3 12 9 2 11 7 11 2 7 11 7 11 2
27 3 13 3 10 10 9 10 11 2 12 7 12 9 2 2 10 11 12 0 0 0 9 0 12 9 13 2
31 10 0 9 10 11 9 2 11 3 2 16 10 0 9 13 4 7 13 4 9 2 0 0 3 13 13 2 3 3 0 2
12 11 13 3 10 9 2 7 9 3 3 13 2
28 10 0 9 3 11 13 3 10 9 10 9 2 11 3 13 10 9 2 7 0 9 1 3 11 13 11 9 2
42 10 0 9 3 15 10 0 0 9 2 11 3 10 0 9 0 2 11 11 11 2 10 9 9 3 13 9 1 2 2 9 0 0 13 2 7 9 3 3 13 13 2
15 10 11 1 3 13 13 2 7 3 3 13 10 9 2 2
22 10 10 9 10 3 3 9 0 11 11 0 0 13 2 2 10 9 3 13 10 3 2
14 13 2 16 15 10 11 0 2 7 13 7 15 13 2
9 7 3 0 10 9 10 9 2 2
27 10 0 9 9 2 10 11 11 9 3 13 13 10 9 2 10 11 0 9 0 10 9 0 12 9 13 2
11 10 0 9 10 0 0 11 0 9 13 2
21 10 0 9 9 9 13 10 11 2 10 11 7 10 11 11 2 7 3 3 0 2
26 10 11 3 13 2 9 10 11 13 3 3 3 2 7 10 9 0 11 3 10 9 0 9 13 3 2
11 9 2 11 11 2 0 9 2 0 9 2
52 9 9 2 11 2 0 2 2 11 2 0 2 9 2 9 2 11 2 0 2 2 7 11 11 2 0 2 2 11 11 2 0 2 2 11 2 0 2 9 2 9 2 11 2 0 2 2 11 2 0 2 2
57 9 9 2 11 2 0 2 2 11 11 2 0 2 9 2 9 2 11 2 0 2 2 11 2 0 2 2 11 2 0 2 2 11 11 2 0 2 9 2 9 2 11 2 0 2 2 11 2 0 2 2 11 11 2 0 2 2
25 9 2 0 9 2 0 9 7 0 9 13 10 9 11 11 0 9 9 9 0 9 0 11 9 2
33 12 9 7 3 13 13 10 0 9 1 2 3 10 0 9 11 11 3 9 13 9 10 9 2 3 10 0 9 11 0 9 13 2
15 10 0 9 1 0 9 10 0 9 10 9 3 3 13 2
36 10 12 9 1 11 11 2 11 2 9 9 7 3 10 9 13 10 9 2 3 11 11 11 2 11 2 12 9 13 9 10 9 10 9 0 2
34 11 11 3 10 0 9 13 14 2 3 12 9 2 10 11 11 2 11 11 2 7 10 0 0 9 2 11 11 11 10 0 9 13 2
15 10 11 0 9 9 9 1 13 10 2 11 2 0 9 2
22 2 10 9 1 13 15 2 16 10 9 1 3 0 13 2 16 10 9 13 10 9 2
4 2 3 7 2
30 3 10 11 0 9 1 2 3 7 3 2 3 13 10 0 9 7 7 13 4 2 3 3 7 13 10 9 10 9 2
20 3 3 13 10 9 9 2 3 7 3 3 10 9 2 13 2 3 10 9 2
9 3 3 13 2 16 13 10 9 2
18 2 10 0 9 1 3 13 10 9 2 7 3 11 9 13 9 9 2
20 2 3 10 0 9 9 13 10 0 13 2 7 10 0 9 3 10 9 13 2
6 3 13 0 9 1 2
16 2 3 3 13 10 9 9 2 7 3 10 9 7 0 13 2
