200 11
20 9 13 16 4 0 9 1 11 3 12 9 13 9 9 2 3 16 7 9 2
11 0 9 13 4 13 9 1 11 7 11 11
32 0 0 9 1 9 4 15 15 15 4 3 0 16 9 15 0 9 14 4 0 13 4 0 1 9 2 0 9 7 3 0 2
41 15 4 9 2 9 9 2 15 4 9 9 11 1 11 2 15 4 9 1 0 9 2 11 2 2 2 2 13 4 1 12 11 11 2 9 0 9 9 0 9 2
39 11 4 1 9 2 12 9 2 13 9 1 9 9 15 9 1 11 0 0 9 11 2 11 2 1 15 9 13 16 4 1 9 4 0 1 0 3 9 2
26 3 1 0 9 15 9 2 0 0 9 11 0 9 2 11 2 11 2 13 15 9 9 9 1 11 2
23 15 13 1 9 15 15 13 9 0 9 9 1 0 7 0 11 2 2 2 13 4 11 2
13 3 7 1 9 0 9 2 0 4 0 9 9 2
16 11 2 15 4 3 9 15 9 11 1 0 9 1 9 11 2
16 0 9 13 16 4 0 9 13 12 9 9 1 0 9 1 11
30 9 4 1 9 2 12 9 2 13 9 9 16 16 4 0 9 9 11 11 11 13 0 9 1 9 11 1 15 9 2
16 9 4 1 15 15 4 0 9 3 0 1 15 9 1 11 2
14 9 1 9 9 1 11 7 11 3 4 13 4 0 2
28 9 0 9 1 11 7 11 11 11 11 13 4 12 9 16 4 15 9 9 0 9 7 9 0 9 1 9 2
35 15 15 13 9 1 11 15 4 13 13 11 7 9 9 9 2 11 4 13 9 1 9 1 9 2 15 9 13 9 7 9 1 0 9 2
44 0 4 9 13 3 12 9 2 9 1 9 9 1 0 9 7 9 1 9 2 16 7 9 1 0 9 1 0 9 0 9 7 9 9 11 1 9 9 0 7 0 0 9 2
12 13 15 9 15 4 15 9 13 9 0 9 2
13 11 4 13 0 9 11 9 11 0 1 0 9 2
43 13 15 16 4 0 9 2 15 4 15 13 1 11 3 9 16 4 13 12 9 9 0 9 2 13 0 9 1 15 15 13 2 2 0 9 2 2 9 7 15 0 9 2
35 7 2 13 14 15 9 9 9 3 13 15 3 4 0 9 9 2 9 9 7 9 7 9 9 1 12 9 15 13 13 7 9 0 9 2
36 2 2 11 4 0 2 0 9 13 2 15 4 9 1 15 15 4 0 2 9 2 13 16 13 1 9 15 11 2 7 15 4 13 13 3 2
10 9 4 13 9 7 13 9 1 9 2
8 15 13 9 11 1 0 11 2
18 9 4 1 9 2 12 9 2 13 9 1 9 9 9 11 11 11 2
29 9 9 7 9 11 11 13 16 15 9 7 9 14 13 13 16 13 0 9 2 7 13 16 4 15 9 4 0 2
11 9 0 9 0 9 13 3 4 13 9 2
32 0 9 4 4 2 1 11 2 0 1 9 0 9 0 11 0 1 9 1 9 2 16 4 13 13 0 9 1 15 9 9 2
25 9 13 1 12 9 9 2 1 15 4 12 9 13 2 11 2 1 9 15 9 11 1 0 9 2
13 9 11 7 0 9 9 11 11 4 4 0 9 2
16 13 14 11 2 11 7 11 13 0 2 2 0 9 2 2 2
35 3 1 12 9 1 0 9 13 4 9 1 0 0 9 1 0 9 11 2 3 1 11 2 16 15 9 13 1 9 11 1 0 9 11 2
12 0 9 2 13 9 2 4 15 15 4 0 2
23 2 2 16 13 1 11 2 13 13 9 1 9 9 1 9 9 2 2 2 13 4 11 2
13 14 4 3 13 15 1 0 9 2 13 0 9 2
12 2 2 15 4 11 7 11 1 11 11 11 2
15 15 1 15 4 4 0 9 2 7 13 16 4 3 13 2
41 9 9 9 0 4 1 9 12 2 16 16 4 0 0 9 2 15 4 9 0 1 9 11 1 9 0 9 2 0 1 9 9 2 3 15 4 13 0 0 9 2
16 0 9 9 13 4 11 16 1 0 9 13 9 1 9 9 2
31 0 9 13 4 16 4 11 1 12 7 12 9 13 0 9 1 15 0 9 2 7 16 15 0 9 14 4 13 9 9 2
6 4 3 13 1 9 2
26 0 9 11 2 9 2 13 4 15 9 1 11 3 16 15 0 9 4 9 2 3 9 9 0 9 2
29 3 12 9 2 3 1 11 2 13 4 0 9 1 9 2 7 12 15 13 4 1 0 9 2 9 0 9 11 2
21 12 4 1 0 9 9 0 9 1 9 9 9 15 15 9 14 13 1 0 9 2
15 11 2 0 9 15 9 14 13 0 9 1 15 0 9 2
23 0 9 1 12 9 15 13 13 0 9 9 1 0 9 7 13 15 15 9 9 7 9 2
39 13 15 16 4 15 9 1 9 9 13 13 2 16 16 4 11 0 9 4 9 11 2 16 16 4 9 11 11 13 1 9 1 11 1 9 2 9 2 2
19 9 9 11 13 4 1 9 1 9 11 7 13 9 1 0 9 9 9 2
21 1 0 9 2 12 9 4 4 12 0 9 2 12 9 12 2 7 15 9 12 2
20 15 4 13 13 15 9 2 7 15 4 4 0 9 2 2 2 13 4 11 2
5 0 9 11 13 9
19 0 9 11 11 11 7 15 0 9 11 11 13 4 16 4 13 0 9 2
28 11 7 0 11 3 15 13 9 0 9 7 9 1 9 1 0 11 2 3 16 3 9 0 9 13 1 9 2
24 9 13 9 9 2 15 13 0 9 7 9 1 0 9 0 9 1 9 2 7 9 0 9 2
27 0 1 9 4 4 9 2 2 9 7 9 2 2 0 0 9 2 0 9 1 11 2 1 9 11 11 2
22 11 13 12 9 1 0 9 15 13 13 15 9 1 11 2 12 3 16 1 0 9 2
25 11 2 12 2 3 4 13 1 0 11 9 1 0 0 0 9 1 2 11 2 9 0 1 11 2
40 2 2 11 4 2 7 2 3 4 1 9 16 2 1 9 2 3 7 3 13 9 14 3 7 14 3 2 3 0 0 9 2 2 2 13 4 0 9 11 2
52 2 2 11 4 13 9 9 0 0 9 2 11 2 7 13 7 13 9 7 9 0 0 9 2 11 2 15 4 4 1 0 9 2 2 2 13 4 0 9 11 11 8 11 11 1 11 2 2 13 2 11 2
15 1 12 9 9 2 0 9 13 9 7 9 15 3 13 2
26 0 9 13 4 0 9 11 11 2 15 4 13 16 0 0 11 4 13 2 7 2 12 9 1 9 2
20 9 9 11 11 0 4 1 9 1 11 2 0 9 7 0 0 9 0 9 2
23 2 2 9 0 9 1 11 13 9 1 0 9 0 11 1 11 2 2 2 13 4 11 2
12 1 15 15 13 0 9 11 11 8 11 11 2
15 15 4 12 1 0 9 1 9 2 7 4 0 16 0 2
22 2 2 13 16 3 4 13 2 13 2 13 7 13 15 15 13 9 9 9 2 2 2
27 9 0 9 11 11 2 12 2 0 4 1 9 0 9 2 1 3 12 1 12 9 9 3 1 9 9 2
14 11 4 4 0 1 9 1 12 2 12 7 12 9 2
18 9 2 15 15 13 0 15 4 3 13 9 2 13 4 15 3 9 2
15 11 2 9 0 9 14 13 2 16 4 9 1 15 0 2
26 0 9 14 3 13 0 9 2 9 7 0 9 9 15 15 3 13 7 13 15 13 2 13 0 9 2
22 15 4 9 14 3 0 2 7 9 1 0 9 0 9 0 1 15 9 4 3 0 2
27 12 9 13 4 9 1 9 0 9 12 9 2 7 4 15 13 1 9 0 9 7 3 4 0 1 11 2
25 9 0 9 11 11 2 3 0 9 9 1 0 9 2 13 4 16 4 9 13 13 9 9 9 2
18 9 0 0 9 2 0 9 0 9 2 13 3 0 3 7 0 9 2
40 16 4 9 0 1 3 12 9 13 16 15 3 1 12 9 11 3 3 13 14 15 0 9 1 11 2 0 9 9 11 11 11 13 4 9 16 13 9 11 2
37 2 2 13 13 14 3 1 0 9 15 9 3 3 13 15 9 7 13 9 9 2 7 14 13 9 3 2 0 2 9 2 2 2 13 4 11 2
28 3 1 0 9 0 9 13 4 1 15 9 0 9 11 1 0 9 11 11 11 2 15 4 13 1 9 11 2
8 0 4 9 1 0 0 9 2
21 1 0 9 2 11 13 16 4 15 9 13 1 0 0 9 16 4 13 15 9 2
15 9 4 13 9 1 9 2 0 9 11 7 0 0 9 2
9 0 9 4 4 0 1 9 11 2
17 1 15 9 2 9 13 13 0 0 9 15 4 13 13 1 9 2
13 11 13 16 4 11 0 1 9 9 11 1 9 9
28 2 2 0 15 4 15 9 2 16 4 0 13 9 1 15 4 15 0 13 1 9 15 15 13 1 0 9 2
15 1 0 9 1 11 1 9 2 12 9 2 13 4 12 2
16 9 1 9 13 9 0 0 9 2 9 9 7 0 9 9 2
36 1 9 12 2 12 2 0 9 11 13 4 1 9 9 0 3 0 9 11 2 13 4 0 9 1 0 7 0 9 2 7 13 9 0 9 2
12 9 13 16 9 4 0 2 16 4 9 0 2
25 15 4 0 9 1 9 15 13 1 9 1 9 2 7 0 9 3 0 9 1 9 13 0 9 2
20 9 15 13 16 4 9 9 0 9 13 1 9 0 9 0 9 11 7 11 2
45 3 16 13 9 9 15 4 13 9 9 9 11 16 16 16 4 0 2 13 2 9 2 11 4 13 16 4 15 11 13 1 0 9 1 0 9 2 15 15 13 1 9 0 9 2
43 11 4 13 16 4 2 2 0 9 9 1 0 9 2 1 9 12 9 9 2 3 13 2 7 13 4 7 0 9 2 9 2 9 1 9 1 9 9 2 9 7 9 2
22 1 9 15 9 13 9 1 9 0 1 9 9 2 9 7 9 9 1 9 7 9 2
23 9 0 0 9 3 13 16 16 4 15 9 0 9 0 3 1 3 9 7 9 1 9 2
30 1 0 9 2 11 4 4 0 3 1 12 9 1 9 9 2 11 2 15 15 13 1 9 0 9 1 9 1 9 2
11 9 4 1 15 9 13 2 3 2 9 2
4 0 9 13 9
14 3 12 9 2 1 2 12 9 0 4 3 12 9 2
20 11 2 16 15 13 9 7 13 0 9 2 15 4 4 3 0 1 9 11 2
17 0 11 11 13 1 9 11 2 11 2 11 2 11 11 7 11 2
13 9 15 9 4 13 7 0 9 16 3 0 9 2
17 13 15 16 4 0 9 0 1 9 3 9 1 15 4 0 11 2
12 9 4 9 15 15 13 1 0 9 0 9 2
25 0 9 4 3 0 1 0 9 2 16 4 4 3 15 13 16 2 9 2 7 16 2 9 2 2
27 0 9 3 15 13 1 0 9 2 7 15 13 13 7 1 0 9 2 16 1 15 9 0 9 1 9 2
25 9 11 4 13 16 0 9 12 16 16 4 9 11 11 1 9 13 13 0 9 11 7 11 11 2
7 9 13 1 9 0 9 2
13 0 9 13 15 1 9 2 0 9 7 0 9 2
6 9 9 1 9 13 2
9 11 4 13 11 12 9 12 9 2
11 1 15 2 3 15 13 1 11 7 11 2
23 0 9 13 12 9 1 11 11 2 11 2 0 9 2 16 9 2 15 4 3 13 9 2
11 1 9 0 9 13 1 11 1 9 9 2
18 13 15 13 1 9 3 9 13 9 2 16 7 3 4 0 7 0 2
28 9 1 14 0 9 0 9 13 4 1 9 15 4 1 9 13 1 9 9 9 2 9 7 9 1 12 9 2
27 9 7 9 1 9 4 15 0 9 2 15 15 13 1 9 2 0 0 9 7 9 2 15 13 9 9 2
9 3 15 13 1 11 7 0 9 2
12 13 4 1 0 0 9 1 9 9 7 9 2
18 13 15 1 9 16 15 13 9 1 9 2 9 9 7 13 0 9 2
26 0 9 4 0 0 9 1 9 15 4 0 9 13 16 4 0 9 2 7 4 15 13 2 9 2 2
12 9 15 14 13 0 9 3 15 13 1 9 2
11 0 9 0 4 0 9 0 9 0 9 2
14 16 15 14 9 3 13 2 13 4 15 13 1 9 2
5 0 9 4 11 2
11 3 1 15 15 15 13 7 9 11 11 2
16 9 9 7 9 1 9 4 3 0 2 16 9 1 9 2 2
21 11 4 12 9 13 9 2 15 4 13 12 9 9 11 2 15 15 0 11 13 2
22 1 9 0 9 9 13 1 9 2 1 9 3 15 1 0 9 1 0 7 0 9 2
26 0 9 1 0 9 4 9 12 8 12 9 11 2 7 0 4 11 11 2 3 0 16 9 11 2 2
33 1 9 13 1 11 2 1 9 1 11 2 11 7 11 7 11 11 2 1 9 1 11 7 11 7 1 9 1 11 7 9 11 2
53 0 9 15 15 13 9 9 15 9 4 1 9 0 2 7 1 0 2 0 2 9 2 1 9 15 1 0 2 15 9 13 12 1 12 2 7 0 9 16 7 0 9 9 2 9 2 15 13 1 9 1 9 2
18 1 9 9 11 2 1 9 11 13 15 0 9 11 7 11 7 11 2
10 11 3 15 9 13 2 7 15 13 2
13 9 4 0 9 1 9 1 15 9 2 3 0 2
12 9 4 0 9 1 9 16 0 9 15 9 2
20 1 15 9 4 13 9 11 7 7 15 16 13 15 4 13 7 0 0 9 2
21 9 2 1 0 9 2 9 2 4 0 9 15 13 3 0 0 9 3 0 9 2
44 3 15 13 9 1 9 13 15 9 16 16 4 2 2 0 2 7 2 0 2 2 3 0 0 9 2 0 9 1 9 2 0 9 7 3 2 2 1 0 9 0 9 9 2
10 11 11 0 4 12 9 12 1 11 2
14 15 9 13 2 16 9 13 13 3 12 9 9 9 2
18 9 13 7 0 0 9 2 3 0 2 0 9 15 13 9 1 9 2
18 7 2 3 13 16 15 15 3 3 7 14 13 7 15 13 1 11 2
26 3 9 15 3 13 0 9 1 9 0 9 3 9 9 7 9 2 7 9 4 0 1 0 9 9 2
13 9 0 9 3 4 15 13 3 9 11 13 9 2
8 9 15 4 1 9 1 11 2
16 0 9 3 15 13 16 9 0 0 9 1 0 9 1 3 2
13 0 9 13 13 1 9 1 15 4 0 15 9 2
27 1 0 0 9 13 15 16 9 9 0 15 9 2 9 2 9 2 9 2 0 9 2 0 9 7 9 2
15 11 4 9 0 9 2 3 11 11 2 2 9 9 9 2
10 0 9 9 13 0 9 0 1 9 2
22 9 0 9 4 2 1 0 9 15 9 2 13 3 4 11 13 15 12 9 1 9 2
41 9 16 9 7 9 0 0 2 0 2 0 7 0 9 1 0 9 13 0 7 0 9 1 9 9 0 9 2 7 9 0 9 16 0 2 0 9 9 0 9 2
10 9 9 13 9 9 2 9 7 9 2
18 9 15 13 13 1 3 9 9 2 3 2 2 3 1 9 0 9 2
14 11 2 0 9 2 9 11 2 0 4 9 1 11 2
20 9 13 0 9 1 9 9 3 0 0 7 0 9 2 15 4 1 0 9 2
14 0 0 9 4 11 11 2 1 12 9 12 9 2 2
27 0 0 9 2 11 2 0 11 11 11 2 11 2 0 4 9 0 9 15 13 16 0 9 0 0 9 2
27 1 9 11 12 2 0 9 0 0 7 0 9 0 4 3 12 0 9 2 1 15 4 12 1 0 12 2
33 0 9 9 13 0 9 0 7 0 9 7 0 0 9 2 15 4 0 3 7 3 1 0 9 2 7 3 7 3 1 9 9 2
18 0 9 11 4 0 2 1 9 1 11 2 1 0 0 9 9 11 2
23 9 1 15 4 12 9 0 2 7 0 0 4 3 0 1 9 1 15 15 13 0 9 2
50 1 15 2 1 9 9 15 13 13 15 0 0 0 9 2 9 9 2 15 13 9 9 16 4 13 9 2 9 7 13 9 2 7 9 9 2 15 13 9 9 16 4 13 0 9 2 9 7 9 2
5 9 13 12 9 2
23 9 9 2 11 11 2 7 9 15 4 13 2 11 11 2 0 4 0 7 3 0 9 2
26 1 9 1 9 0 9 2 9 4 0 2 15 13 14 3 9 9 2 7 13 13 1 12 9 9 2
20 1 9 9 13 9 1 9 7 9 2 0 9 2 9 0 9 7 9 9 2
8 13 15 1 0 7 0 9 2
28 3 0 9 0 4 15 13 13 9 12 9 7 4 3 0 9 13 9 0 0 0 9 16 13 11 1 9 2
15 9 4 3 2 0 9 9 9 2 15 15 13 9 9 2
35 16 16 9 13 1 9 1 0 9 9 2 3 15 3 13 9 9 15 9 2 15 4 0 9 1 9 0 7 0 9 1 9 3 0 2
22 16 9 13 12 0 9 2 3 4 0 2 7 16 4 15 9 0 13 9 1 9 2
12 9 9 13 2 9 2 9 2 9 7 9 2
20 15 12 9 13 15 13 1 9 1 0 9 9 1 9 9 2 9 7 9 2
20 11 4 4 9 0 9 15 4 4 3 0 1 9 12 9 1 9 0 11 2
30 9 13 4 0 2 1 9 2 2 0 2 1 9 9 2 2 0 2 1 9 2 7 0 2 0 2 0 9 2 2
29 9 4 0 9 0 9 2 1 9 9 2 9 9 2 9 9 0 9 1 9 2 13 16 9 9 2 9 7 3
10 0 9 9 11 4 4 9 11 11 2
18 1 9 1 0 11 13 15 0 9 11 1 15 4 15 12 7 13 2
22 3 4 15 13 7 11 11 2 11 2 0 9 2 2 11 11 2 9 2 7 11 2
9 3 4 15 0 2 0 7 0 2
21 9 11 4 4 11 2 11 2 11 2 9 4 4 11 11 2 7 9 11 11 2
20 0 9 15 13 9 1 9 3 4 1 12 9 1 12 9 2 3 1 9 2
8 9 15 4 1 11 1 11 2
20 9 4 0 9 1 9 2 9 2 1 9 0 9 7 1 9 9 1 0 2
12 0 9 11 4 13 7 13 15 16 0 9 2
21 9 15 9 15 14 13 13 3 1 9 2 1 0 1 0 9 13 13 0 9 2
21 15 1 9 7 9 0 1 9 4 9 2 0 9 2 9 2 9 7 0 9 2
14 13 4 12 1 9 9 1 9 1 0 9 11 11 2
36 9 13 15 9 16 13 3 7 3 1 9 0 9 15 4 13 1 0 9 2 3 13 15 1 9 1 9 7 15 1 15 15 13 0 9 2
20 1 9 0 0 9 13 1 9 2 11 2 1 9 3 13 0 9 7 9 2
18 1 0 9 2 0 9 4 9 0 9 0 9 2 3 1 9 9 2
12 0 9 4 9 0 0 9 1 14 15 9 2
7 1 9 15 13 9 9 2
16 1 0 9 15 9 13 9 0 9 1 11 0 2 0 9 3
19 9 4 1 0 9 9 0 1 9 9 2 15 3 2 3 2 4 9 2
6 3 4 14 0 9 2
12 9 13 7 13 9 2 9 0 7 0 9 2
14 9 15 13 1 12 9 2 0 2 0 7 0 9 2
14 0 9 1 9 9 2 2 9 2 2 4 13 11 2
