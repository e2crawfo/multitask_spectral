76 11
23 3 2 15 4 13 1 9 2 7 4 4 13 0 2 15 15 4 7 13 1 9 9 2
15 13 9 12 9 2 9 11 2 0 9 2 13 12 8 2
22 9 9 7 9 13 9 1 9 2 13 1 11 7 4 4 13 3 9 10 9 0 2
19 9 9 0 4 4 13 1 9 11 11 2 7 10 0 2 1 11 11 2
25 9 0 2 9 3 13 1 9 11 2 11 2 9 0 7 11 2 15 13 14 13 0 1 9 2
22 1 9 9 15 15 13 2 9 11 4 13 10 9 1 9 13 1 3 12 1 9 2
14 15 9 15 15 13 3 10 9 0 2 7 7 0 2
22 10 9 0 1 9 2 13 1 10 9 0 0 2 13 1 9 9 0 1 9 0 2
20 13 9 10 9 10 9 0 15 13 14 15 13 3 7 9 1 3 3 0 2
17 15 13 3 1 9 9 0 2 13 1 9 9 0 10 9 10 2
18 9 9 14 15 13 1 1 3 2 16 14 15 13 9 1 10 9 2
20 2 9 15 15 13 2 9 0 13 1 9 9 1 9 2 4 13 9 0 2
19 1 3 2 9 13 14 13 9 0 0 2 0 2 3 2 1 10 9 2
15 12 16 13 3 2 9 1 9 13 4 13 1 12 9 2
19 1 14 13 9 9 2 15 13 4 13 1 10 9 2 3 1 10 9 2
16 3 2 9 13 1 9 0 2 13 15 9 0 7 9 0 2
20 11 2 12 9 7 12 9 2 14 4 13 9 9 1 9 13 1 9 0 2
18 9 0 13 1 11 2 9 2 13 10 9 1 9 13 9 1 9 2
18 2 12 2 11 13 9 1 9 7 13 16 15 13 9 13 1 15 2
21 2 9 2 2 9 1 9 2 2 9 1 9 1 9 15 13 4 13 10 9 2
34 2 12 2 9 0 13 9 0 2 11 2 9 9 5 9 1 9 11 2 0 2 2 15 13 9 1 10 9 0 1 9 7 9 2
29 12 2 9 1 9 13 1 9 14 13 16 9 0 14 4 13 10 9 0 1 9 10 9 1 9 10 9 0 2
24 2 12 2 11 2 11 2 11 7 9 0 4 13 9 0 1 9 10 9 9 1 9 12 2
22 2 10 9 4 13 9 1 9 1 14 4 13 2 7 10 13 9 10 9 1 9 2
16 7 2 1 9 7 9 2 15 13 14 15 13 1 10 9 2
11 13 10 9 14 13 1 10 9 10 10 2
13 10 9 1 9 2 1 13 9 2 13 1 9 2
19 7 9 15 4 13 1 0 9 2 16 15 15 4 13 15 9 1 9 2
23 13 1 9 14 13 16 9 14 15 4 13 7 3 14 4 4 13 1 15 15 15 13 2
30 13 7 3 15 13 1 13 3 13 16 0 9 2 16 0 2 4 13 3 9 2 15 15 13 1 10 3 0 9 2
14 1 10 9 10 2 14 13 13 1 10 9 10 11 2
17 3 13 14 15 13 1 9 2 13 16 4 13 10 9 1 9 2
7 1 15 15 13 15 13 2
14 3 3 15 15 4 13 2 3 10 9 13 14 13 2
15 10 9 3 15 3 12 9 14 4 13 14 13 1 11 2
18 9 3 15 13 14 13 2 7 4 4 13 14 13 16 4 4 13 2
9 14 15 13 13 14 15 13 15 2
10 15 13 3 3 16 14 15 13 13 2
16 14 15 13 13 9 15 15 13 1 9 9 0 7 1 9 2
17 9 13 2 1 9 2 9 3 0 14 13 13 1 9 9 0 2
8 15 14 13 14 13 9 9 2
11 13 15 14 15 13 2 10 9 3 13 2
7 13 3 13 1 9 9 2
7 3 14 3 13 13 15 2
17 14 15 15 13 0 2 14 15 13 13 1 11 3 1 10 9 2
12 13 14 13 1 9 3 15 13 1 9 15 2
13 0 9 14 13 14 13 1 9 9 10 9 13 2
13 15 13 3 13 9 14 13 10 9 1 10 9 2
13 4 13 14 15 13 15 1 15 10 9 13 15 2
15 14 13 9 14 15 13 2 9 13 0 2 14 3 13 2
16 7 3 13 15 9 2 14 13 13 14 14 15 13 1 9 2
20 10 3 0 9 0 1 9 9 1 2 9 2 4 13 4 13 1 9 11 2
26 2 9 11 1 9 9 5 1 12 12 1 9 13 1 9 10 5 3 9 0 2 4 13 13 2 2
21 11 4 13 13 10 9 10 9 2 9 2 13 1 10 9 10 9 0 10 9 2
55 10 3 0 9 0 10 9 1 2 9 5 0 2 0 1 9 0 4 13 1 9 2 9 7 9 1 9 13 1 0 0 1 9 10 12 10 15 2 13 1 9 9 10 9 9 2 4 13 1 11 2 11 7 11 2
16 3 2 9 11 13 1 12 2 16 9 2 15 13 0 2 2
25 9 0 1 9 1 2 9 5 0 2 13 3 9 15 4 13 1 9 13 1 9 3 1 9 2
25 10 3 0 9 0 1 10 9 0 1 9 2 0 2 4 13 1 10 9 10 9 11 1 11 2
15 9 0 13 10 9 0 10 10 9 9 1 2 0 2 2
42 16 9 0 0 15 4 13 14 13 0 2 15 13 10 9 0 1 9 10 11 2 9 10 0 13 0 2 9 13 13 3 0 1 9 10 12 10 9 10 12 10 2
27 10 3 0 9 0 0 10 9 1 9 13 9 10 11 1 12 2 15 13 9 9 0 2 9 0 2 2
20 11 11 13 1 9 1 2 9 2 3 9 2 15 15 13 9 1 9 0 2
31 2 3 1 12 9 2 1 3 10 9 15 4 13 1 9 9 15 13 1 2 9 2 1 15 15 13 1 2 9 2 2
18 3 2 1 9 0 9 2 11 2 4 13 1 0 1 2 11 2 2
42 1 9 0 9 2 11 2 4 4 13 1 2 11 2 2 3 1 9 0 15 13 9 2 11 2 2 1 14 13 9 0 2 7 2 11 2 1 14 13 9 0 2
12 3 2 9 9 4 13 2 13 3 10 9 2
17 15 13 16 9 0 10 9 9 1 9 11 13 9 0 10 9 2
5 13 9 9 0 2
14 1 12 9 2 1 9 11 4 13 9 1 9 0 2
14 1 9 10 12 10 4 13 12 9 1 9 1 11 2
14 1 9 15 4 13 10 9 3 0 2 13 4 13 2
20 13 1 9 9 10 12 10 10 12 9 13 0 1 9 1 9 10 9 0 2
30 1 9 9 0 1 12 2 11 15 4 13 1 0 9 9 9 10 0 2 13 13 1 9 1 9 0 7 0 11 2
13 1 12 11 4 13 1 12 9 0 1 9 9 2
13 1 12 2 9 11 10 12 10 15 13 9 0 2
14 1 12 2 3 9 10 11 2 11 13 9 9 0 2
