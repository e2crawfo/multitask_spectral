120 17
11 11 1 0 9 9 13 0 9 13 4 2
14 0 9 3 13 4 11 1 9 13 13 4 13 11 2
16 11 9 11 9 13 15 0 9 9 13 14 15 1 9 13 2
9 3 15 9 9 13 14 9 13 2
6 3 0 9 9 13 2
13 9 9 13 1 9 0 9 0 0 3 13 4 2
11 3 11 14 11 9 13 14 9 15 4 2
9 9 11 9 1 0 9 13 4 2
16 11 0 12 9 14 13 0 9 3 13 11 0 9 13 13 2
21 11 9 0 9 11 11 0 12 9 1 12 9 1 11 11 9 9 9 13 4 2
15 12 9 11 9 13 14 0 11 9 9 1 9 11 11 2
18 15 12 9 1 12 9 9 1 9 0 14 0 9 13 14 9 13 2
25 15 3 11 11 11 9 11 9 11 11 2 11 11 11 9 11 11 9 3 13 9 9 12 13 2
34 15 2 11 11 9 14 2 11 9 13 2 9 13 9 13 2 9 9 13 9 11 11 0 9 9 1 13 9 13 14 13 4 13 2
16 15 1 2 12 9 9 13 4 14 14 10 9 13 4 4 2
13 10 9 2 11 0 11 9 13 9 11 9 13 2
67 3 2 9 9 13 4 0 9 7 9 9 1 13 2 11 9 9 12 2 12 2 12 2 12 2 14 2 2 12 2 11 2 0 9 9 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 9 1 11 0 11 9 9 9 9 13 9 13 4 2
12 0 11 9 11 11 0 9 3 13 4 4 2
15 11 9 14 11 9 11 11 11 13 4 14 13 4 4 2
16 11 0 9 0 9 11 13 4 0 9 9 11 9 13 4 2
11 15 10 9 11 13 14 3 9 13 4 2
12 3 15 12 0 9 11 13 4 14 13 4 2
13 10 9 14 15 11 13 4 14 0 9 9 13 2
25 0 9 15 11 13 14 14 2 11 9 11 11 11 11 0 14 15 13 4 14 14 10 9 13 2
24 11 0 9 14 2 11 0 9 14 14 11 9 9 1 9 13 4 13 14 15 11 9 13 2
8 12 9 14 11 9 3 13 2
12 9 7 11 9 15 13 4 14 9 9 13 2
20 9 11 9 2 9 9 9 7 11 11 9 0 9 14 11 13 9 13 4 2
58 9 11 11 11 9 12 12 12 9 14 2 9 9 11 9 12 12 12 9 14 12 0 11 13 14 2 3 2 9 11 11 9 12 9 14 2 9 11 9 12 9 14 2 11 11 9 12 9 14 12 0 11 13 14 9 13 4 2
46 15 9 1 2 9 11 9 2 9 9 9 2 11 9 0 12 9 14 1 12 12 12 9 7 9 2 12 12 12 12 12 12 12 0 9 0 11 1 13 4 14 11 9 13 4 2
25 11 9 11 11 7 11 0 9 13 14 0 0 9 2 15 11 9 3 13 4 4 14 13 4 2
24 11 9 14 11 9 0 9 9 13 4 4 14 13 1 0 9 11 9 11 11 1 9 13 2
10 15 9 3 9 13 4 4 14 13 2
17 11 0 11 9 14 11 11 9 0 9 9 13 4 4 13 15 2
21 11 11 9 9 1 9 3 12 12 9 13 14 11 9 14 11 0 9 13 4 2
15 11 11 9 11 11 9 9 12 12 9 13 14 13 4 2
16 3 11 9 9 12 12 9 1 12 12 9 13 14 13 4 2
7 12 0 9 11 9 13 2
16 10 0 11 9 14 13 12 0 9 9 14 13 14 11 13 2
12 12 1 12 12 12 9 10 9 13 4 4 2
8 9 11 14 10 0 9 13 2
8 3 3 9 12 12 9 13 2
19 3 3 11 2 11 2 11 9 10 9 13 14 11 9 9 13 4 4 2
23 9 11 2 11 2 9 13 0 12 9 11 11 9 9 9 13 9 13 4 14 9 13 2
12 11 1 11 11 9 0 12 9 1 13 4 2
15 3 9 1 9 9 0 15 9 1 9 9 9 13 4 2
15 3 9 1 13 13 9 13 4 14 11 9 11 11 13 2
10 15 9 13 0 14 9 15 13 4 2
11 15 9 2 15 9 1 9 9 13 4 2
10 9 13 4 14 9 15 15 13 4 2
8 3 13 4 14 11 11 13 2
21 9 2 9 1 3 13 14 13 2 3 9 13 9 13 4 14 11 9 9 13 2
35 11 11 1 11 9 9 11 11 9 1 9 2 9 1 13 14 14 2 11 3 15 13 15 3 9 0 14 15 13 4 14 14 9 13 2
13 11 11 9 11 11 2 11 11 0 9 9 13 2
22 9 1 0 9 1 9 9 14 3 11 9 0 9 0 0 9 9 9 9 13 4 2
18 9 15 9 13 14 14 11 9 14 15 9 14 14 0 0 11 13 2
43 11 9 3 13 14 2 9 0 9 0 9 13 14 2 9 2 11 1 14 11 9 3 13 4 4 14 0 9 2 9 1 9 0 9 12 9 9 9 14 13 4 13 2
13 12 0 9 14 9 14 9 9 14 9 13 4 2
8 12 9 14 11 9 13 4 2
12 12 9 14 9 13 13 0 9 1 13 4 2
11 12 9 13 14 0 9 3 13 4 2 2
11 15 1 15 9 2 9 14 9 13 4 2
26 10 12 14 13 0 9 9 13 15 1 3 13 14 13 9 13 15 9 13 13 4 14 9 13 13 2
19 10 9 11 13 1 15 11 14 0 9 13 14 14 14 0 14 9 13 2
17 11 13 0 9 11 9 11 9 13 4 0 9 1 3 13 4 2
17 10 9 11 3 9 13 4 14 11 9 9 1 9 13 4 4 2
16 9 9 9 9 14 9 0 9 14 9 9 9 13 3 13 2
15 10 9 12 9 13 14 11 9 0 11 9 13 4 4 2
8 15 11 9 14 3 13 4 2
14 3 11 9 1 11 9 13 4 14 10 9 13 4 2
25 11 0 9 9 9 11 11 7 0 9 9 11 11 7 9 11 11 9 3 0 9 9 13 4 2
25 11 1 14 9 9 1 14 2 10 9 12 9 1 14 9 10 9 13 14 1 14 9 13 4 2
18 12 9 1 14 9 3 13 4 3 12 9 1 14 9 3 13 4 2
25 3 11 14 2 11 14 9 9 9 11 9 13 4 0 9 3 13 4 14 14 9 13 4 4 2
15 3 11 9 0 9 9 11 9 2 11 9 1 3 13 2
24 9 9 0 9 11 0 9 14 9 13 13 4 14 14 2 15 12 9 13 14 14 13 4 2
7 15 11 9 0 13 4 2
10 3 10 9 13 11 3 9 13 4 2
32 15 13 4 12 9 1 0 10 0 9 13 4 1 2 9 9 12 9 1 0 9 13 14 9 13 14 14 9 13 4 4 2
29 9 9 11 9 9 13 0 0 9 11 9 9 14 11 13 15 11 11 9 10 0 3 13 14 14 13 4 4 2
25 11 0 9 11 11 9 10 9 9 14 11 11 2 12 9 1 14 9 9 9 13 0 9 13 2
26 11 13 4 0 9 9 11 9 2 12 9 1 14 9 9 13 0 9 13 4 14 14 15 13 4 2
7 11 9 9 9 9 13 2
15 15 13 11 14 0 9 13 14 14 13 4 14 15 13 2
12 9 9 0 14 2 3 9 9 13 4 4 2
8 11 11 9 0 9 13 4 2
14 9 0 9 9 13 13 4 4 14 14 11 13 4 2
17 11 2 11 1 9 3 13 9 4 4 14 11 9 11 11 13 2
12 11 9 9 0 9 13 4 11 13 14 2 2
10 0 9 9 0 9 9 9 9 4 2
14 10 9 11 7 11 0 9 9 9 3 13 13 4 2
16 11 2 11 1 9 9 9 2 9 9 9 3 13 13 4 2
10 15 3 11 9 14 13 15 13 4 2
12 11 3 0 9 0 15 9 14 15 13 4 2
15 11 2 11 1 9 9 12 9 14 10 9 3 13 4 2
11 3 9 13 0 9 0 9 13 4 4 2
16 3 9 9 9 9 10 9 13 4 11 9 1 13 9 13 2
11 10 9 9 3 9 9 13 13 4 4 2
10 0 9 9 0 9 13 4 13 15 2
13 3 9 9 13 13 0 9 9 15 9 13 4 2
11 0 9 0 9 1 9 0 9 13 4 2
15 10 9 9 14 13 4 9 11 9 9 4 9 13 4 2
9 11 9 11 9 11 9 13 4 2
13 10 9 11 9 9 4 14 14 15 9 13 4 2
15 9 9 9 13 14 15 0 9 13 4 14 9 13 4 2
26 11 9 9 0 9 13 13 9 13 14 0 0 9 14 2 11 9 0 9 9 14 14 11 11 13 2
8 11 9 9 15 11 13 4 2
12 11 9 0 9 13 4 4 14 11 13 4 2
11 11 9 9 13 4 14 13 12 14 13 2
10 3 15 3 9 14 15 13 4 13 2
8 3 13 0 9 9 1 13 2
25 3 2 0 9 14 2 0 9 14 0 14 0 9 15 3 13 0 9 9 13 14 14 13 4 2
30 12 0 11 9 9 14 11 9 14 14 11 11 0 9 9 14 3 0 9 14 0 14 15 10 9 10 13 4 13 2
9 15 9 13 4 14 9 9 13 2
7 3 3 15 13 13 13 2
9 3 15 9 14 13 4 13 11 2
22 12 11 9 9 1 0 11 11 2 11 0 9 9 1 11 9 13 4 14 9 13 2
8 0 9 11 9 10 9 13 2
16 3 2 9 0 0 9 9 14 9 3 12 9 13 4 4 2
14 0 9 9 9 9 14 1 9 13 4 8 14 15 2
