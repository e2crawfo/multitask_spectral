1596 11
10 11 2 10 9 1 10 9 1 11 2
14 10 9 13 12 9 7 10 9 13 3 1 10 11 2
9 7 3 13 1 10 9 3 0 2
52 10 2 9 1 9 2 2 1 10 9 15 13 10 9 0 7 10 9 0 0 2 13 0 7 0 2 10 9 15 13 10 0 9 1 9 2 1 9 2 1 9 2 1 9 1 10 9 13 1 3 0 2
12 9 1 3 0 9 13 1 10 9 9 0 2
36 11 11 2 9 0 9 1 10 9 2 7 11 11 2 9 0 9 1 10 9 0 2 1 10 9 0 2 1 10 9 7 10 9 0 2 2
11 15 13 1 13 1 10 9 1 10 9 2
12 10 9 0 1 0 9 14 13 3 10 9 2
12 15 13 3 1 10 9 13 10 9 1 9 2
40 10 9 0 4 13 3 10 9 10 9 1 0 9 3 1 10 9 0 1 10 11 1 10 9 1 10 11 0 15 13 15 0 1 10 11 11 1 12 9 2
12 7 2 10 11 14 13 3 10 9 1 9 2
19 10 11 1 10 9 1 11 11 1 10 9 1 11 1 11 2 12 2 2
24 15 13 3 10 9 3 0 7 15 1 10 9 1 13 10 9 1 10 9 3 13 10 9 2
43 11 11 2 13 10 12 9 12 1 11 7 13 10 12 9 12 1 11 2 13 10 9 0 7 9 0 1 10 9 1 10 12 9 2 15 10 9 13 10 9 1 9 2
23 15 13 1 10 9 16 15 4 13 1 12 7 1 12 2 13 3 10 9 1 10 11 2
29 1 12 2 16 10 11 4 13 10 9 1 10 9 2 11 2 15 4 4 13 1 10 9 2 4 13 10 11 2
22 13 12 9 15 10 9 13 1 7 10 9 1 9 2 15 13 10 9 0 1 9 2
38 11 15 13 1 10 0 9 1 9 2 7 10 2 9 2 1 10 9 1 11 11 4 13 0 2 11 13 16 10 9 14 13 3 7 13 3 13 2
23 10 9 1 9 4 13 1 10 12 9 1 10 9 1 9 11 1 10 9 1 11 11 2
36 10 0 9 2 1 11 11 7 11 11 2 13 10 9 1 10 9 13 1 13 10 9 1 10 0 0 9 0 7 15 10 9 15 13 0 2
19 10 0 11 2 9 1 11 11 2 2 15 13 1 10 9 0 7 0 2
17 15 4 13 9 1 9 0 1 10 9 1 10 11 7 11 11 2
25 10 9 13 1 10 11 7 10 9 0 0 13 16 10 9 4 13 1 10 9 1 10 9 0 2
21 11 13 10 9 1 10 9 11 11 11 2 15 4 13 10 0 9 11 8 11 2
49 10 9 1 9 1 9 13 1 10 9 1 11 0 1 10 11 1 11 13 10 9 1 11 13 1 10 9 7 10 9 1 12 9 1 9 1 9 15 4 13 10 9 2 10 9 7 10 9 2
24 10 9 10 3 13 13 10 9 1 10 0 9 15 13 10 9 7 10 9 1 9 1 9 2
7 15 4 13 10 12 9 2
35 10 9 13 1 10 9 1 10 9 2 11 11 7 11 2 13 1 10 9 1 10 9 2 1 10 9 2 1 10 9 7 1 10 9 2
23 15 4 13 3 1 9 2 10 9 11 11 2 11 11 2 10 9 11 11 2 11 11 2
31 11 11 2 13 11 11 10 12 9 12 1 11 2 1 10 11 2 13 10 9 7 9 0 2 1 10 0 9 0 2 2
31 1 10 9 1 9 2 11 2 2 15 13 3 0 2 15 4 15 13 1 10 3 0 9 2 0 1 15 1 10 9 2
11 10 9 13 9 12 9 1 10 9 0 2
23 3 3 0 9 1 10 9 3 0 16 0 2 10 9 13 0 7 13 1 10 0 9 2
17 15 13 10 9 1 9 1 9 1 13 11 1 9 1 9 0 2
22 10 9 13 1 10 0 9 13 1 10 9 1 9 1 9 0 1 10 9 0 13 2
35 15 4 3 13 1 12 9 2 10 9 1 11 1 10 9 2 7 10 9 1 11 1 10 9 2 10 9 15 13 1 10 9 1 11 2
16 11 7 11 4 13 1 12 1 10 9 0 7 13 1 12 2
29 10 0 9 2 15 4 13 10 9 1 10 9 11 11 1 13 13 10 9 13 1 9 1 10 9 1 10 9 2
30 10 0 9 2 3 2 2 9 1 9 2 2 13 10 9 1 9 1 10 9 3 13 1 10 9 1 10 11 0 2
16 11 2 10 9 9 2 13 1 9 1 10 9 2 10 9 2
48 10 9 0 0 2 15 13 10 9 1 10 9 1 9 7 10 9 1 9 13 1 10 9 1 10 0 9 2 13 10 0 9 2 16 10 9 0 13 1 10 9 0 13 1 12 1 12 2
11 15 14 13 0 3 1 10 12 0 9 2
19 10 9 0 1 9 1 11 13 10 9 0 0 2 1 3 12 9 2 2
14 15 13 10 9 10 3 0 1 11 13 10 9 2 2
20 3 13 1 10 9 1 11 2 15 13 9 13 1 2 11 11 2 1 12 2
21 10 0 9 0 1 10 9 13 1 10 9 1 10 0 9 4 13 9 1 12 2
25 1 10 9 1 9 2 15 13 1 10 9 1 12 9 7 14 13 3 10 0 9 1 12 13 2
17 10 9 1 10 9 13 10 9 0 1 10 9 1 10 9 0 2
25 10 9 1 11 13 10 9 0 0 2 13 1 10 9 1 10 11 7 10 9 9 1 10 11 2
32 10 9 4 13 1 12 9 0 2 10 11 11 2 1 15 13 10 11 12 2 7 10 11 2 11 11 13 1 10 11 12 2
14 10 9 0 4 15 3 13 13 10 9 1 10 9 2
25 10 9 1 9 15 13 1 9 1 10 9 15 13 7 14 13 3 10 9 1 9 1 10 9 2
17 1 10 9 1 10 9 2 10 9 13 1 13 10 9 1 12 2
20 10 12 11 2 13 1 9 1 10 12 9 12 4 4 13 1 9 1 11 2
44 15 13 3 3 10 11 2 15 13 1 10 9 1 10 10 9 2 7 3 10 0 9 11 2 3 16 10 9 1 11 2 15 13 10 3 10 9 1 9 1 10 12 9 2
10 10 9 13 3 0 16 10 9 0 2
17 10 9 0 13 0 1 10 9 1 10 9 1 9 2 7 0 2
8 15 13 0 1 10 11 0 2
54 10 9 11 13 1 10 9 11 11 2 15 12 9 13 0 2 3 10 9 1 10 9 2 11 11 2 10 9 1 10 9 2 11 11 2 10 9 1 10 9 2 11 11 2 7 10 9 1 10 9 2 11 11 2
7 10 9 13 11 11 11 2
16 15 4 13 9 9 2 1 9 2 1 10 9 1 9 11 2
15 1 10 9 2 10 9 4 13 1 10 11 1 11 11 2
29 10 11 1 11 15 13 10 9 1 9 7 1 0 9 2 1 10 0 9 0 2 1 13 3 10 9 1 11 2
24 10 9 2 13 1 10 9 1 9 13 1 10 9 11 11 2 13 16 15 14 15 13 15 2
23 15 13 10 9 1 10 11 10 11 11 11 11 11 2 7 4 4 3 13 1 10 9 2
16 10 10 9 0 1 10 9 11 15 13 1 10 9 1 11 2
15 15 15 4 13 10 12 1 10 12 9 7 3 15 14 2
11 9 7 9 13 1 10 0 9 1 9 2
12 15 15 13 10 11 1 11 3 10 9 1 2
11 15 13 7 15 13 10 9 15 4 13 2
19 10 11 13 10 9 1 10 9 0 0 1 12 9 1 10 9 1 11 2
31 10 9 1 10 9 2 11 11 2 4 13 16 15 13 16 10 9 2 13 11 1 1 9 1 10 9 0 7 0 2 2
26 1 9 3 0 2 12 9 13 0 16 15 13 10 0 9 7 10 0 9 2 7 13 10 9 0 2
48 10 9 0 1 10 9 4 13 10 12 9 1 10 11 7 10 9 11 2 10 9 1 10 9 11 2 1 10 9 1 10 11 1 11 10 12 9 13 10 9 1 9 1 9 1 10 11 2
28 10 9 1 10 11 13 1 13 10 9 1 10 9 1 9 1 9 2 7 13 10 9 1 10 11 1 3 2
10 10 9 12 13 12 9 1 9 0 2
34 15 15 13 1 10 9 0 1 10 9 0 7 0 3 13 7 9 1 10 3 0 9 1 10 9 9 1 13 10 9 1 10 9 2
28 10 9 1 10 11 11 2 9 9 1 11 10 11 2 1 11 13 10 9 0 0 13 1 11 1 10 9 2
26 1 12 7 12 2 15 4 13 1 9 2 9 7 9 1 10 9 2 8 8 2 13 1 9 12 2
22 15 13 10 9 1 10 0 9 0 0 13 1 10 11 2 13 10 9 1 10 9 2
46 9 1 10 9 12 1 10 9 1 11 11 4 3 13 1 10 9 1 10 11 11 2 15 13 1 9 1 13 10 9 11 11 2 1 10 9 1 13 1 10 9 0 1 11 11 2
21 11 13 10 9 1 9 2 1 12 9 9 12 7 9 12 2 1 12 9 12 2
18 1 9 12 2 10 0 9 0 15 13 1 10 9 2 12 15 13 2
39 16 15 15 4 13 2 15 4 13 1 10 9 1 10 9 1 10 9 7 1 15 13 13 2 15 15 4 3 13 16 15 13 16 15 13 1 10 9 2
24 1 12 2 15 15 13 1 10 9 3 1 10 9 1 10 9 7 15 13 1 13 10 9 2
74 15 15 13 1 13 11 11 2 3 13 1 10 9 1 10 9 2 11 11 2 11 11 2 13 3 1 10 9 11 11 1 10 11 7 10 9 11 11 11 1 10 11 2 3 16 11 11 2 10 9 1 11 7 0 9 2 13 1 10 9 0 7 0 1 10 9 2 15 13 3 1 10 9 2
15 15 3 13 3 1 10 9 0 7 10 9 3 13 0 2
18 1 12 2 10 9 7 9 0 11 13 10 9 0 1 10 9 0 2
23 1 9 2 15 13 10 9 0 1 10 9 1 10 9 0 0 1 12 2 1 11 11 2
21 15 3 13 10 9 1 9 2 10 9 2 10 9 2 7 10 9 1 10 9 2
7 15 4 13 1 10 9 2
13 10 9 1 10 11 13 10 9 7 13 12 9 2
27 1 10 9 2 1 10 9 1 10 9 2 12 9 0 2 10 9 7 10 9 1 9 2 13 1 9 2
13 10 9 1 11 4 13 1 10 9 1 10 9 2
16 15 15 13 3 1 10 9 1 10 9 2 15 13 10 9 2
48 11 11 13 3 11 2 10 9 1 10 9 11 15 13 10 3 0 9 0 1 10 9 1 10 0 9 2 0 1 10 9 0 2 13 9 1 10 9 1 12 9 1 9 7 9 1 9 2
10 2 11 13 3 0 1 10 9 0 2
30 10 9 1 10 9 13 0 7 2 3 1 10 9 0 2 15 4 4 13 1 9 1 10 9 7 10 9 0 0 2
16 1 13 16 12 9 4 13 1 10 9 1 10 9 1 11 2
48 10 9 13 12 9 1 10 9 1 10 0 9 1 11 1 9 1 10 9 1 9 1 10 9 2 11 2 1 10 9 11 12 7 10 11 11 1 10 9 1 11 2 8 8 2 1 11 2
41 11 11 11 2 1 10 9 0 11 11 11 1 11 2 2 13 10 12 9 12 2 1 11 1 11 2 13 10 9 0 0 2 9 1 10 9 11 2 11 11 2
36 10 9 1 9 2 15 2 14 4 13 3 16 10 9 0 15 13 3 9 7 16 15 14 4 3 13 1 10 9 10 9 7 10 9 0 2
29 10 12 9 1 9 0 1 11 11 11 2 11 12 1 12 2 4 13 1 10 9 0 1 10 9 1 10 9 2
18 10 9 1 10 9 4 3 13 7 10 9 13 10 9 1 10 9 2
62 10 9 11 0 1 10 9 2 1 2 13 10 9 1 9 3 13 1 11 11 11 2 7 15 13 10 9 1 10 10 9 0 15 13 1 10 15 7 10 0 9 0 2 7 2 3 0 2 15 13 1 10 9 0 1 10 9 1 10 9 0 2
62 16 11 12 7 11 13 10 2 9 7 10 9 2 1 11 2 15 14 13 3 10 9 1 9 1 11 7 13 10 9 1 10 9 1 10 9 1 11 7 10 13 1 10 9 1 9 1 10 9 3 0 1 15 15 13 10 9 1 11 7 11 11
15 15 15 13 1 10 9 1 10 9 7 10 9 1 9 2
19 10 9 7 10 9 1 10 9 4 4 13 1 10 12 1 10 12 9 2
26 11 13 12 9 2 7 2 1 11 2 10 0 9 13 12 9 1 9 7 12 5 1 10 9 0 2
16 1 3 2 15 14 4 13 10 9 0 1 10 9 1 11 2
12 10 9 4 13 11 0 1 10 12 9 12 2
14 15 13 1 10 9 13 11 9 2 9 7 9 2 2
15 11 11 13 10 9 0 0 13 10 12 9 12 1 11 2
19 13 15 0 2 16 0 2 1 13 10 9 0 1 10 9 1 10 9 2
19 1 3 2 10 9 0 13 3 10 9 0 1 3 1 10 9 1 9 2
29 10 9 4 13 9 1 9 1 9 0 0 10 9 1 9 2 10 9 1 9 2 10 9 1 9 7 10 9 2
22 10 9 1 11 13 15 1 10 0 9 15 10 9 1 10 11 7 10 11 13 0 2
7 12 8 13 3 1 9 2
20 10 9 13 1 10 9 10 9 13 1 10 9 1 10 9 1 15 15 13 2
21 11 11 13 10 12 9 12 1 11 13 10 9 0 2 9 1 10 11 11 0 2
15 10 9 4 13 1 10 9 1 10 9 1 11 1 12 2
28 1 12 11 11 13 1 10 9 11 11 7 11 11 2 10 9 9 13 1 10 9 1 10 9 1 9 0 2
37 10 9 4 13 1 11 2 15 15 4 13 1 11 1 12 2 7 15 15 13 12 9 1 12 9 7 10 9 1 12 9 1 9 1 1 11 2
18 10 9 9 1 10 9 2 13 10 11 11 2 13 1 10 9 0 2
16 10 9 1 10 9 7 1 10 9 0 1 9 13 3 0 2
18 15 13 1 10 9 0 1 11 11 2 13 10 9 7 13 11 11 2
22 10 9 1 10 9 13 11 11 15 4 13 10 9 1 10 9 3 16 1 10 9 2
13 10 9 10 3 0 13 10 9 2 1 10 9 2
45 11 13 13 2 1 10 9 0 7 10 9 0 2 10 10 9 1 10 9 7 15 13 3 10 9 2 10 9 7 10 0 9 1 13 1 10 9 7 1 10 9 1 10 9 2
13 10 9 0 1 10 9 3 16 10 9 4 13 2
25 10 9 13 10 9 0 2 1 10 9 2 1 13 7 13 10 9 2 7 1 9 1 9 0 2
17 9 0 2 9 0 15 15 4 3 13 13 10 9 1 13 10 9
23 11 11 4 4 13 1 12 9 0 1 10 9 1 11 7 9 1 10 11 0 1 11 2
17 11 11 13 10 9 7 13 1 11 11 1 10 9 1 10 9 2
14 10 11 11 13 10 9 1 10 9 11 2 1 11 2
24 15 13 1 10 9 1 10 0 9 1 9 1 9 7 13 10 9 1 0 9 1 10 9 2
16 1 9 12 2 11 11 11 13 1 9 1 11 2 11 2 2
38 1 10 9 1 10 9 2 13 1 10 9 1 10 11 1 9 1 10 9 0 1 10 1 12 9 2 2 10 9 13 3 10 9 1 9 1 13 2
9 15 13 3 0 2 1 11 11 2
26 13 1 11 2 15 13 16 10 9 4 13 9 2 7 11 4 13 1 11 11 15 15 13 1 9 2
10 11 11 13 10 9 1 10 9 11 2
33 1 9 2 16 15 13 10 9 15 13 10 9 0 1 15 13 1 10 9 2 15 13 10 9 15 13 10 9 1 10 9 0 2
15 10 9 13 15 1 10 9 0 2 3 1 10 9 0 2
53 10 9 4 13 2 1 10 9 1 10 9 12 2 11 11 2 9 1 10 9 2 7 11 11 13 1 13 11 1 10 9 0 15 11 15 13 1 9 1 0 9 2 7 13 10 9 7 10 9 1 10 9 2
23 9 1 10 11 2 1 15 1 10 0 9 2 13 1 9 13 13 10 9 1 10 9 2
22 1 10 9 2 15 13 3 10 9 1 9 7 10 9 1 9 2 15 10 11 11 2
29 1 9 2 10 12 9 9 13 10 9 13 10 9 1 10 9 1 10 11 15 10 9 13 0 1 12 5 9 2
22 1 15 2 2 15 13 1 10 9 0 2 15 13 3 15 13 1 10 9 0 2 2
29 15 13 1 10 9 1 10 9 15 15 13 13 2 15 13 3 10 9 1 13 2 3 0 2 7 15 13 9 2
17 11 13 10 9 0 1 10 9 1 11 1 10 11 0 1 11 2
18 10 9 1 10 9 4 4 13 1 9 1 1 12 9 10 9 0 2
18 10 0 9 13 1 10 9 1 9 0 2 1 15 13 11 7 11 2
8 11 4 13 1 9 10 9 2
35 10 9 13 10 9 0 1 10 9 13 2 1 15 10 9 1 9 4 13 2 7 10 9 13 2 15 10 9 1 9 14 4 13 2 2
27 10 9 0 13 1 10 9 1 13 10 9 0 1 13 10 9 2 9 12 7 12 1 10 11 0 2 2
23 10 9 14 4 1 3 13 10 9 1 10 9 1 10 9 1 10 9 1 10 9 0 2
22 15 4 13 1 10 9 0 7 1 10 9 1 9 1 9 0 1 10 9 1 9 2
6 10 9 4 3 13 2
31 15 15 13 1 10 9 1 10 9 1 10 11 1 10 9 1 1 10 9 1 10 11 7 1 10 9 1 1 10 11 2
30 11 12 13 10 9 1 10 9 11 1 10 9 1 10 9 1 9 1 13 10 9 1 10 11 1 10 9 1 9 2
18 11 13 10 9 0 2 13 1 10 9 1 10 11 7 10 9 11 2
13 10 9 1 10 9 0 13 1 10 9 0 0 2
14 15 13 10 9 1 0 9 2 12 1 12 9 2 2
19 10 9 1 4 13 3 1 10 9 0 14 13 3 1 9 1 15 13 2
19 11 13 16 10 9 0 15 13 13 11 1 10 9 15 13 9 1 9 2
23 1 10 9 1 10 9 2 10 0 9 2 7 10 0 9 2 15 4 13 1 10 11 2
25 1 10 9 1 10 9 13 1 10 11 2 10 9 1 9 0 1 10 11 14 13 3 10 9 2
27 15 15 13 1 13 10 11 11 7 13 1 15 13 0 2 7 15 14 13 9 1 10 9 1 10 9 2
30 13 1 9 1 10 9 13 1 10 9 0 1 11 2 15 15 13 1 15 1 10 9 0 10 3 0 1 10 9 2
17 15 15 13 1 10 0 9 1 10 9 2 10 9 7 10 9 2
37 3 16 15 13 10 0 9 2 1 10 9 1 10 11 7 4 13 1 10 9 1 11 2 9 13 10 9 1 10 9 0 1 10 11 1 11 2
17 11 11 4 3 13 10 9 9 15 4 13 1 10 9 1 11 2
9 15 15 13 10 9 2 0 2 2
18 1 12 1 12 2 15 13 10 9 1 10 9 1 9 1 10 9 2
34 1 3 2 10 9 1 10 11 1 10 9 0 13 0 13 3 1 9 1 13 10 9 1 10 9 1 10 9 1 9 1 10 9 2
48 11 11 2 13 10 12 9 12 1 11 2 9 10 12 9 12 1 11 2 13 10 9 0 2 9 7 9 2 9 7 9 1 10 9 1 11 2 15 13 12 9 2 1 13 1 10 9 2
25 9 1 10 9 2 10 9 0 1 10 9 0 2 11 11 2 15 13 1 15 13 1 10 9 2
31 10 9 4 13 1 10 9 1 10 11 15 13 10 9 3 1 11 1 10 9 1 11 1 10 9 1 10 9 1 11 2
30 11 12 9 13 10 9 1 9 3 1 11 12 2 10 9 0 1 13 1 3 1 10 11 1 10 9 1 10 11 2
26 10 9 1 10 9 13 3 1 4 13 2 3 1 10 9 0 2 3 1 12 9 7 0 3 3 2
22 10 9 13 3 0 2 0 7 0 3 16 10 3 0 2 7 15 13 11 3 2 2
7 10 9 15 13 3 0 2
11 10 9 0 13 10 9 1 10 11 0 2
25 1 10 9 15 4 4 13 1 10 12 9 1 10 9 11 1 11 2 1 10 9 1 11 11 2
46 15 15 13 1 10 9 1 9 2 7 4 13 1 10 9 1 9 11 2 9 11 11 2 15 13 16 15 4 4 13 1 15 1 10 9 2 7 1 11 2 15 15 13 10 9 2
45 11 11 2 12 9 12 2 12 9 12 2 13 10 9 0 4 13 2 1 10 9 12 2 1 10 9 1 10 9 1 10 9 0 1 10 9 0 1 10 9 1 10 11 11 2
24 1 9 10 9 10 9 0 13 1 10 9 0 11 2 11 13 10 9 15 13 1 10 9 2
15 15 13 15 15 15 13 3 10 11 2 7 2 11 2 2
23 15 13 9 1 10 11 7 9 1 9 1 10 11 0 1 11 1 10 9 1 10 9 2
10 1 13 1 12 15 13 10 9 0 2
42 10 9 0 1 9 13 10 9 2 10 9 1 9 7 15 15 15 13 10 9 1 9 1 10 9 2 8 3 2 10 9 2 9 1 10 9 1 10 9 2 2 2
46 15 4 4 13 1 10 9 1 9 1 10 9 2 2 4 13 3 1 10 9 1 10 11 12 2 11 11 2 9 0 1 10 11 0 1 9 1 10 9 7 10 9 2 11 2 2
20 15 15 13 1 12 9 1 9 13 7 13 10 15 1 10 15 1 10 9 2
29 10 9 11 0 2 13 1 10 9 0 1 11 13 1 10 9 1 11 1 13 10 9 2 11 11 2 12 2 2
12 15 4 13 10 10 9 3 1 10 9 0 2
16 3 13 12 9 7 15 13 3 1 10 0 9 13 1 11 2
29 10 9 0 13 0 1 10 9 0 7 15 13 15 15 13 11 10 2 12 9 2 0 1 10 9 1 10 9 2
43 10 9 13 0 1 10 9 2 7 15 4 3 13 1 10 9 3 0 1 16 10 11 15 13 1 10 9 15 15 4 13 1 10 9 0 7 1 10 9 1 10 9 2
7 15 4 13 10 9 12 2
24 10 9 0 13 15 1 13 10 9 4 13 10 3 1 9 7 15 13 10 9 1 10 9 2
11 15 4 3 13 1 10 9 1 9 0 2
34 3 2 11 4 13 3 10 9 1 10 9 2 13 1 9 9 2 7 4 13 9 1 10 9 0 1 10 9 1 11 7 11 11 13
18 10 9 13 1 11 11 13 0 1 10 9 1 10 9 1 10 9 2
17 1 4 13 10 11 2 11 13 7 13 10 9 0 1 10 11 2
32 10 0 9 2 10 9 13 1 12 1 11 11 4 13 2 2 12 2 11 2 1 10 9 1 11 11 7 1 10 9 11 2
19 10 11 13 1 13 10 9 0 1 10 9 0 1 9 0 1 10 9 2
16 10 9 4 13 9 1 11 2 9 13 1 10 9 0 0 2
40 15 13 1 10 9 1 10 9 1 10 11 1 13 10 9 1 9 0 16 10 9 11 8 11 2 10 9 11 2 7 1 9 1 11 11 7 11 1 11 2
14 3 2 15 3 4 13 10 0 9 7 13 3 13 2
38 10 9 1 10 9 13 3 0 3 16 15 1 10 11 4 13 1 3 12 9 2 1 3 1 10 9 1 10 9 1 10 9 2 3 12 9 2 2
29 10 9 13 3 10 9 1 10 3 0 1 11 1 10 9 9 2 1 9 1 11 7 1 11 1 10 11 2 2
15 1 10 11 2 11 11 11 2 2 15 13 3 10 9 2
33 10 9 1 10 9 4 4 13 3 1 10 9 1 10 9 1 10 11 11 2 15 13 3 1 3 3 1 10 9 1 10 9 2
24 1 3 2 1 12 2 11 13 13 10 9 1 9 1 10 9 2 7 15 1 3 0 3 2
20 15 14 13 16 1 13 10 9 2 15 4 13 1 10 9 1 10 3 0 2
21 3 3 2 15 4 4 13 16 10 9 1 10 9 4 13 10 9 0 1 8 2
18 10 9 0 4 13 1 10 9 8 7 8 1 10 9 10 9 0 2
16 10 11 4 1 10 9 13 2 3 3 2 12 12 1 9 2
43 1 9 1 10 9 1 10 9 2 9 4 4 13 1 10 10 9 1 10 9 2 13 1 10 9 1 10 9 1 10 9 0 2 1 10 9 1 10 9 10 3 0 2
28 11 13 11 10 12 9 7 10 9 11 15 13 1 10 9 1 11 1 15 13 10 9 1 10 9 1 11 2
10 10 9 13 3 12 5 1 10 9 2
8 3 2 7 3 15 13 15 2
30 3 1 10 9 1 9 7 1 9 2 11 13 3 10 9 7 4 13 7 13 10 10 9 1 10 9 1 10 9 2
34 10 9 1 10 9 0 1 9 0 4 13 10 9 1 15 13 1 12 1 12 9 0 11 12 12 12 1 10 9 11 1 9 0 2
30 1 15 15 13 10 9 0 2 15 15 13 1 11 2 11 2 11 2 11 2 11 2 11 2 11 2 7 3 11 2
32 3 1 10 9 1 9 2 10 9 13 0 2 7 10 9 2 0 2 2 15 13 1 10 9 2 4 13 1 10 9 0 2
24 15 13 10 9 1 15 13 1 11 11 2 9 1 11 0 1 10 9 1 9 7 1 9 2
62 10 9 1 10 0 9 1 9 2 9 9 1 0 9 9 2 13 10 9 0 0 13 10 9 2 1 12 2 10 9 13 14 13 3 3 3 13 1 10 9 2 1 10 9 1 9 9 9 7 9 2 11 2 2 15 13 3 10 10 0 11 2
21 11 11 13 3 10 0 9 2 1 9 0 2 13 1 3 1 15 1 10 8 2
21 2 15 13 11 15 4 13 10 9 1 10 9 2 16 1 9 2 16 1 9 2
13 13 16 11 11 7 10 0 11 11 13 10 9 2
26 10 9 1 10 9 0 13 1 3 16 10 9 0 1 10 9 13 1 10 9 10 9 2 10 9 2
14 3 13 1 10 9 7 1 10 9 1 10 9 0 2
18 10 9 0 4 13 2 10 9 4 13 1 9 15 4 13 10 9 2
57 10 9 15 13 3 10 9 2 11 2 15 13 1 10 9 1 9 0 2 1 10 10 9 13 1 11 11 11 2 1 10 11 7 10 3 0 9 2 0 2 7 1 10 9 2 9 2 13 1 10 3 0 9 1 10 9 0
17 1 12 2 10 12 11 13 10 9 2 13 1 10 9 1 9 2
40 10 0 9 1 10 9 13 13 1 10 11 0 2 1 12 11 2 1 11 2 2 10 3 9 1 10 9 0 13 10 9 1 10 9 0 1 10 9 2 2
12 3 1 12 11 14 13 3 16 3 12 9 2
30 1 10 9 2 11 2 1 10 9 1 10 0 9 2 13 1 13 10 9 1 10 9 7 13 3 3 16 3 11 2
25 15 13 3 10 11 2 12 2 7 15 13 13 10 9 1 10 12 9 1 9 13 1 11 11 2
25 15 4 13 1 12 1 10 9 1 10 9 0 11 11 2 7 4 13 1 10 9 11 1 12 2
51 10 9 1 11 11 4 13 1 10 9 1 10 9 2 1 10 9 1 10 11 2 1 10 9 0 1 10 11 2 1 1 10 9 1 11 1 11 7 1 1 10 9 1 11 2 10 9 1 10 9 2
4 15 13 12 2
13 3 2 15 15 13 10 9 7 10 9 13 2 2
19 1 11 2 10 9 0 11 14 4 3 13 2 7 10 10 9 4 13 2
30 10 9 7 10 9 1 10 11 13 10 9 0 1 9 0 1 10 9 1 11 2 13 1 10 12 9 1 10 11 2
25 10 12 9 1 9 4 13 10 12 9 12 1 11 1 10 11 12 1 3 16 9 1 10 12 2
27 15 13 3 2 1 10 0 9 2 10 9 13 10 9 2 3 16 10 9 0 0 9 13 10 9 12 2
18 15 4 3 13 1 10 9 1 10 11 11 2 10 9 0 1 11 2
43 1 12 2 10 9 1 10 9 1 10 9 4 13 2 11 11 13 9 1 10 2 11 9 1 0 9 2 2 9 13 1 10 11 1 10 11 1 10 0 9 1 9 2
31 10 9 13 10 11 2 9 2 2 10 12 9 2 9 2 2 10 0 9 2 0 9 2 7 10 9 2 0 9 2 2
29 10 0 9 4 3 4 13 1 10 9 9 1 10 9 2 10 0 9 15 13 1 9 1 10 0 9 13 11 2
8 10 9 13 0 1 10 11 2
21 10 9 13 4 13 1 10 9 1 10 9 0 2 11 2 7 1 10 9 0 2
19 15 4 13 1 10 9 0 1 10 11 2 3 1 10 9 1 10 9 2
59 10 9 4 13 1 10 9 0 12 2 1 10 9 0 12 15 13 11 1 11 2 1 9 1 10 11 2 11 2 11 2 11 2 7 1 10 9 0 12 2 3 12 15 13 11 1 11 2 1 9 1 10 9 2 11 2 11 2 2
25 15 13 1 10 5 1 12 2 15 13 10 9 11 2 13 8 2 1 9 1 10 9 0 11 2
31 10 9 15 15 13 10 12 9 12 1 10 9 11 11 13 10 9 13 1 10 9 1 10 9 1 11 10 12 9 0 2
46 1 9 12 2 15 4 2 3 1 4 13 1 10 0 9 0 2 11 11 11 2 13 10 9 1 10 9 7 9 1 10 9 11 11 11 2 15 13 10 9 0 1 10 0 9 2
10 3 2 10 9 13 0 1 1 11 2
11 9 0 13 3 3 1 9 1 10 9 2
23 1 9 2 15 3 13 10 0 9 2 10 9 0 13 1 10 0 9 13 1 10 9 2
36 15 4 13 1 10 9 1 11 11 2 9 1 10 9 1 11 2 0 9 1 10 9 0 2 3 9 2 7 3 9 1 9 1 12 0 2
30 15 13 10 9 0 1 13 16 10 9 4 13 3 1 10 9 16 10 9 1 2 13 10 0 9 0 2 2 2 2
24 10 9 13 1 11 13 3 0 16 10 11 13 10 9 16 15 4 4 13 10 12 9 0 2
25 10 12 0 9 0 13 10 15 1 10 15 1 12 9 1 10 9 2 1 9 7 1 10 9 2
32 10 12 9 12 2 10 9 13 10 9 0 1 10 9 1 11 11 2 9 1 10 9 2 7 11 11 2 9 1 10 9 2
18 15 4 13 1 10 0 9 1 10 1 10 9 11 1 9 1 9 2
36 1 10 9 1 10 9 10 9 13 1 9 2 11 15 13 15 7 15 13 15 1 10 9 0 16 10 9 13 1 10 9 15 13 1 15 2
13 1 3 10 9 13 3 0 15 15 14 13 15 2
20 15 4 13 1 10 11 0 1 10 11 1 10 11 1 10 9 12 8 12 2
10 1 12 11 11 4 13 1 10 9 2
36 3 10 9 15 15 13 1 10 9 2 3 0 7 9 3 0 2 15 4 13 12 5 10 9 1 10 9 3 16 3 15 13 12 5 2 2
41 1 10 9 1 10 11 1 12 9 0 2 3 12 1 9 13 1 10 9 0 3 16 15 14 13 3 10 9 0 15 15 13 10 9 15 13 1 13 10 9 2
16 10 9 13 10 9 1 10 9 1 10 9 13 1 10 9 2
40 9 1 10 9 1 10 9 1 9 13 1 10 9 1 10 9 7 1 10 9 0 2 11 11 13 10 0 9 2 13 1 9 10 12 9 12 1 12 9 2
16 15 9 13 3 0 7 10 9 4 13 1 9 0 1 9 2
8 11 11 13 10 9 0 0 2
46 15 13 1 10 11 2 1 10 9 2 1 15 15 13 10 0 9 10 3 1 10 9 1 10 11 12 1 11 11 2 7 1 10 11 8 2 13 10 9 1 10 9 0 7 0 2
44 9 1 10 9 11 2 15 13 1 15 13 1 8 2 12 1 10 9 1 10 9 11 7 15 4 13 9 1 10 9 2 0 0 2 1 10 9 2 11 11 7 11 11 2
27 5 2 10 9 0 2 13 10 9 7 13 9 1 10 9 1 9 1 9 0 7 0 1 10 9 0 2
48 10 9 1 11 15 13 1 10 9 13 10 9 1 11 2 12 2 2 1 10 9 0 0 2 1 10 9 1 10 0 9 1 10 9 0 1 10 9 7 10 9 9 1 10 11 11 0 2
15 3 15 13 1 13 10 9 1 11 13 0 1 10 11 2
29 10 9 0 4 4 3 13 1 10 9 1 9 13 1 10 9 0 0 7 13 1 10 9 9 9 2 11 11 2
21 1 10 9 15 4 13 10 9 0 2 13 1 12 9 13 1 10 9 1 9 2
17 12 13 10 9 0 0 15 13 1 10 9 1 11 2 11 2 2
16 13 1 10 11 7 13 1 15 2 10 9 13 10 9 11 2
51 10 9 1 9 2 13 1 12 1 11 11 2 1 10 9 1 11 2 11 1 11 2 2 13 1 10 9 10 9 1 9 4 4 13 3 1 13 10 9 1 10 9 13 1 10 9 1 9 11 8 2
11 10 9 15 13 10 0 9 1 10 9 2
27 11 13 10 9 0 2 13 1 10 9 1 11 7 10 9 11 7 1 10 9 1 10 9 1 10 11 2
21 15 4 13 10 0 9 1 10 9 2 1 15 10 9 1 11 15 4 13 13 2
12 1 15 10 9 13 10 0 9 0 1 11 2
21 10 9 0 2 15 13 9 1 10 9 9 2 4 1 3 13 1 13 10 9 2
32 1 9 2 10 9 13 10 9 1 10 9 2 3 13 10 9 1 10 9 1 9 7 1 10 9 1 9 1 10 9 13 2
49 11 2 7 11 2 13 3 10 9 2 13 1 12 2 3 13 11 2 7 11 7 11 2 1 10 9 2 2 1 12 7 12 2 7 11 2 7 11 2 11 2 11 7 3 11 2 1 12 2
13 1 12 2 15 4 13 1 13 10 12 0 9 2
21 11 11 11 2 11 2 12 9 12 2 11 2 12 9 12 2 13 10 9 0 2
6 10 9 13 10 9 2
15 1 12 2 15 13 10 9 1 10 9 7 1 10 9 2
14 10 9 0 13 0 1 10 0 9 1 10 12 9 2
7 10 11 15 13 1 3 2
10 15 13 10 9 0 1 10 9 11 2
23 11 13 10 9 15 4 3 13 1 9 0 2 3 16 10 15 4 13 3 1 9 0 2
15 15 4 3 13 9 2 3 16 9 1 10 9 1 11 2
6 15 4 3 13 11 2
43 10 9 1 10 11 13 1 12 1 10 9 13 1 12 10 9 2 11 11 7 11 11 11 11 2 2 1 9 1 10 9 1 11 11 11 7 9 1 10 9 11 12 2
17 7 10 9 13 10 9 1 10 9 1 10 9 0 13 1 12 2
22 10 9 1 10 11 4 13 1 10 9 1 3 16 10 9 13 10 9 1 10 9 2
9 9 1 11 9 12 2 12 9 2
9 15 13 10 9 1 9 1 12 2
12 10 11 13 3 1 10 10 9 7 13 0 2
36 10 12 9 13 0 1 10 9 1 10 9 0 2 7 13 10 9 0 2 3 0 2 1 1 10 9 15 11 15 13 3 1 10 0 9 2
20 10 9 4 13 1 10 9 10 9 1 9 13 1 9 10 9 1 10 9 2
20 10 9 13 10 9 0 13 2 15 10 9 1 10 9 0 13 10 9 0 2
24 10 9 4 13 1 12 1 10 9 1 10 11 2 15 13 10 9 1 12 9 1 9 0 2
31 15 13 1 13 16 3 10 9 1 10 9 1 10 11 13 1 10 9 10 9 0 1 10 9 11 2 11 11 11 2 2
15 10 9 13 3 1 9 9 13 1 10 9 0 1 11 2
26 3 2 10 9 1 10 12 0 9 1 9 13 1 9 1 15 13 1 10 9 0 1 10 9 0 2
15 11 11 11 11 13 10 9 0 1 9 0 13 1 11 2
28 11 11 11 11 2 13 10 12 9 12 1 11 8 11 7 13 10 12 9 12 1 11 2 13 10 9 0 2
35 10 9 13 3 10 0 9 1 10 9 0 1 10 11 2 10 9 1 10 9 2 15 15 15 13 10 9 1 10 9 7 1 10 9 2
19 9 1 9 2 11 13 10 9 0 1 10 9 1 10 9 1 10 9 2
38 15 13 10 15 15 13 1 4 13 10 9 0 1 10 11 7 10 11 1 13 1 2 9 0 2 1 13 1 9 1 15 13 1 2 9 0 2 2
23 10 9 13 3 10 9 2 11 11 2 10 9 1 10 9 1 10 9 7 1 10 9 2
7 15 13 15 15 4 13 2
14 10 12 9 0 4 13 10 9 1 9 1 10 9 2
3 9 0 2
21 10 11 13 3 1 10 9 2 11 13 1 13 10 9 1 13 10 9 1 9 2
46 3 10 3 3 0 2 11 15 13 16 10 9 14 15 13 3 3 2 11 15 13 2 1 13 10 9 1 10 9 2 2 7 13 10 9 0 2 7 16 1 3 15 13 9 2 2
19 1 10 9 9 1 10 0 9 13 3 1 11 2 11 11 13 1 0 2
39 10 9 15 10 9 13 1 13 10 9 0 1 10 11 0 0 2 0 13 1 13 10 9 2 3 10 9 2 10 9 7 10 9 2 1 10 0 9 2
11 11 11 13 3 10 9 1 9 8 0 2
24 1 10 9 12 2 10 9 4 13 1 11 2 3 1 11 2 9 3 13 0 1 10 9 2
23 12 13 10 0 9 1 10 9 0 11 7 10 0 9 1 10 9 0 0 2 11 2 2
25 11 13 11 1 9 1 9 2 15 3 10 9 14 13 1 1 12 3 10 9 1 9 1 11 2
10 12 9 1 2 10 9 13 10 9 2
30 10 9 0 4 1 3 4 13 1 10 9 1 11 1 12 1 13 10 12 9 1 10 9 1 10 9 13 1 12 2
31 0 9 1 11 2 10 9 9 0 1 11 13 9 1 10 9 1 13 3 2 1 1 10 9 2 10 9 7 10 9 2
8 11 2 15 13 10 9 2 2
11 10 9 7 9 13 0 1 13 3 0 2
34 10 9 0 13 0 7 10 9 1 10 9 15 13 13 1 11 1 11 1 10 9 1 13 1 10 11 11 7 10 11 1 10 9 2
32 3 1 10 9 2 1 0 10 9 0 2 15 15 13 1 10 9 0 7 1 10 9 1 10 9 1 10 9 2 9 2 2
21 10 0 9 3 0 13 10 9 1 9 2 10 9 0 2 7 10 9 1 9 2
28 10 11 11 15 4 13 3 7 1 10 9 2 10 9 13 10 9 1 10 11 2 15 4 15 15 13 2 2
32 10 9 1 9 13 1 10 11 4 13 10 9 1 10 9 12 1 10 9 7 9 12 1 10 9 1 9 9 2 10 9 2
14 1 15 15 14 4 13 16 10 9 2 13 10 9 2
21 3 2 1 3 2 10 9 4 15 13 1 10 9 2 3 16 15 13 10 9 2
9 10 9 4 13 1 12 9 3 2
12 1 11 2 11 13 10 9 13 1 10 9 2
38 1 12 2 10 0 9 13 3 10 9 1 10 9 7 9 1 10 9 0 1 10 0 9 7 10 9 1 10 9 0 1 10 9 0 7 0 0 2
9 3 2 10 9 14 4 3 13 2
9 10 9 13 10 9 0 1 11 2
16 10 9 15 13 14 13 3 10 9 1 15 13 7 13 0 2
23 1 10 11 11 2 10 9 13 1 10 11 4 13 3 1 9 7 1 9 1 10 9 2
25 1 12 2 15 13 3 10 9 10 9 0 7 11 11 13 1 10 9 1 10 0 9 2 11 2
21 10 9 1 10 9 7 15 10 9 0 13 3 10 9 10 3 0 1 10 9 2
48 1 0 9 2 10 9 13 1 10 11 1 10 9 1 10 9 0 4 4 13 1 11 1 10 9 15 4 13 1 10 9 15 4 13 10 10 9 1 9 1 11 1 10 9 1 10 11 2
26 1 10 9 2 15 13 10 9 1 9 2 16 15 13 1 10 9 0 1 10 9 1 10 9 0 2
36 10 9 1 9 2 7 1 9 1 10 9 2 4 13 1 10 9 0 2 7 10 11 11 2 15 10 9 4 13 10 9 1 10 9 0 2
51 10 9 13 12 9 1 10 9 2 15 12 0 1 11 2 11 2 11 7 11 2 2 1 11 2 1 10 11 7 1 10 11 2 3 16 10 9 0 1 11 2 1 11 2 1 11 7 1 10 11 2
19 3 1 12 12 1 9 4 13 1 10 9 1 9 8 1 9 8 9 2
17 0 9 1 10 9 7 13 1 10 9 2 15 13 10 0 9 2
34 1 9 1 9 1 10 9 2 15 14 13 3 12 9 1 10 9 1 10 9 12 2 7 10 9 1 10 9 14 13 3 1 12 2
10 10 9 14 4 3 3 13 1 9 2
19 1 10 9 2 11 1 11 4 13 10 9 2 9 2 1 10 9 0 2
14 15 4 13 10 9 1 10 9 0 1 10 9 0 2
35 10 9 1 10 9 1 10 9 1 9 3 0 14 4 1 9 3 13 1 13 10 9 1 10 9 0 7 10 9 1 10 9 3 0 2
17 11 13 10 9 0 2 13 1 10 9 1 11 7 10 9 11 2
26 9 1 11 13 10 9 0 0 1 10 9 1 10 11 13 1 10 9 1 11 1 10 9 1 11 2
56 1 10 9 0 2 3 1 12 9 10 10 11 1 11 7 1 11 15 4 13 10 9 1 10 11 1 10 9 7 1 10 9 0 0 2 7 10 9 13 10 9 1 10 9 13 16 12 9 4 13 1 10 9 1 9 2
33 15 15 13 1 10 9 10 3 0 13 1 13 2 1 10 9 0 2 16 10 9 0 0 13 1 10 9 0 7 3 3 0 2
9 1 9 2 15 13 13 10 9 2
19 1 10 9 2 15 15 13 2 2 2 2 10 9 1 10 9 2 2 2
15 3 2 15 4 13 10 0 9 1 9 9 0 1 11 2
24 15 13 10 9 1 10 9 2 11 11 2 15 13 10 9 1 9 0 1 10 9 1 9 2
11 1 15 13 0 7 13 1 3 0 9 2
20 15 13 10 9 0 7 0 3 0 1 10 0 9 13 1 9 1 10 9 2
20 15 13 3 10 0 9 1 13 1 10 0 9 1 11 11 11 11 1 12 2
39 10 9 13 10 9 2 12 9 1 10 11 2 12 9 11 2 12 9 1 11 2 12 9 11 1 13 1 12 1 1 15 13 1 12 1 10 9 0 2
13 11 13 3 3 0 2 15 4 13 1 10 9 2
23 1 10 9 1 10 9 2 10 9 11 15 13 1 10 11 1 11 1 10 9 0 12 2
15 13 3 1 9 3 2 15 4 1 9 4 13 1 12 2
17 10 9 13 1 10 9 1 10 9 7 13 10 0 9 1 9 2
31 15 13 1 10 9 1 15 13 1 10 9 0 1 9 2 1 13 1 10 9 15 13 3 3 10 9 0 1 10 9 2
43 10 9 4 13 1 10 9 6 13 10 9 13 10 9 0 1 10 9 13 1 10 9 1 10 9 0 2 1 10 9 0 2 1 10 9 0 15 15 13 1 10 9 2
17 1 10 0 9 2 10 9 13 0 2 2 15 13 10 9 0 2
27 10 9 13 1 10 9 1 15 13 3 13 1 10 9 7 3 3 0 2 13 11 11 1 10 9 11 2
16 1 10 9 2 10 9 4 13 1 10 9 1 12 7 12 2
36 10 9 0 13 10 2 9 0 2 3 10 9 1 9 1 10 9 1 10 9 1 10 9 7 3 3 1 9 1 10 9 15 15 15 13 2
21 11 1 11 4 13 3 1 10 9 1 10 9 2 9 1 10 9 1 11 11 2
19 10 9 13 9 1 13 3 2 1 13 10 9 1 10 9 0 7 0 2
30 10 0 9 4 13 10 0 9 0 1 10 11 0 2 1 10 0 9 0 15 13 10 0 9 1 10 0 9 0 2
20 10 9 1 10 9 1 11 13 10 9 1 9 0 7 10 9 1 0 9 2
33 1 9 2 15 13 15 13 1 9 7 15 13 3 1 15 4 13 3 3 2 7 16 15 13 3 1 15 13 1 13 10 9 2
10 3 3 2 10 11 11 13 10 9 2
12 10 9 13 1 10 9 0 7 1 10 9 2
27 11 11 2 3 13 2 11 0 2 2 1 10 9 3 2 13 10 9 1 9 1 10 9 1 10 11 2
32 10 9 1 10 9 0 2 1 10 9 0 1 10 9 0 2 4 13 1 10 12 9 1 13 10 9 1 9 7 1 9 2
7 10 9 4 13 1 15 2
9 10 9 0 4 13 10 9 0 2
10 11 7 11 4 3 13 7 1 9 2
15 10 9 1 9 1 10 9 1 10 9 14 13 3 0 2
28 10 11 1 11 13 10 9 1 10 9 8 11 2 11 2 1 11 2 7 11 2 11 2 1 10 11 2 2
50 15 4 4 13 1 10 9 0 1 10 9 1 12 9 2 3 13 1 4 13 10 9 1 10 9 13 12 9 1 10 11 11 7 10 9 0 2 7 1 4 4 13 1 10 9 13 1 11 11 2
36 1 10 9 0 2 10 8 13 13 10 8 0 2 8 2 15 4 3 13 1 10 9 1 10 9 0 7 4 13 1 10 9 1 10 9 2
18 10 9 4 13 1 10 9 0 1 10 11 2 1 10 9 1 11 2
16 9 1 10 12 9 2 15 4 13 12 9 1 12 7 12 2
29 15 4 13 1 12 7 12 9 2 7 10 9 9 14 4 4 13 1 10 9 1 9 0 2 11 1 9 2 2
35 3 2 1 10 11 2 1 11 7 1 10 11 2 15 14 13 3 10 9 0 2 7 10 10 9 13 3 1 9 2 13 1 9 0 2
20 10 9 1 10 9 4 13 1 10 9 0 2 9 0 1 9 7 9 0 2
10 1 10 0 9 2 11 13 10 11 2
15 9 11 13 10 9 0 13 10 11 2 11 2 1 11 2
45 1 13 15 2 10 9 1 9 1 10 11 4 13 10 9 1 9 1 10 9 1 10 11 11 1 13 1 10 9 1 10 0 9 2 14 4 15 3 13 2 10 11 11 2 2
25 11 13 4 4 13 1 10 9 2 15 13 1 15 13 1 15 13 1 10 9 0 7 0 2 2
48 0 1 10 9 1 9 0 7 0 2 15 4 13 1 11 2 1 10 11 2 13 1 10 9 0 2 10 9 1 11 11 11 2 10 9 1 11 2 10 9 1 11 11 7 1 11 11 2
21 10 11 1 11 0 13 15 1 10 9 1 9 1 10 11 1 10 11 11 0 2
40 10 9 2 10 9 11 2 15 13 10 9 1 9 12 9 3 3 2 3 16 10 9 1 9 2 11 1 11 2 12 2 2 13 1 10 0 9 1 9 2
35 1 3 1 13 10 9 15 4 13 10 9 1 12 9 2 9 2 15 1 10 9 1 9 7 10 9 2 3 0 2 1 1 10 9 2
13 15 13 9 1 10 9 1 11 1 9 1 9 2
11 15 14 13 3 3 0 16 15 15 13 2
27 12 9 1 9 1 3 13 10 0 9 1 11 11 2 13 1 10 11 11 11 2 9 11 11 1 12 2
18 15 4 13 10 11 12 2 7 10 11 0 12 1 10 8 8 8 2
12 10 11 13 10 9 0 2 9 1 10 11 2
36 1 10 9 2 11 15 13 1 10 0 9 11 2 11 11 2 15 13 10 3 0 1 13 10 0 9 13 1 10 2 9 1 10 9 2 2
34 10 12 9 12 2 10 9 11 11 11 13 1 11 1 10 9 1 10 9 16 15 13 1 11 2 3 11 7 3 11 2 1 1 2
21 15 15 13 3 1 12 9 1 10 9 1 10 9 1 10 11 2 10 12 9 2
12 2 11 15 15 15 15 13 10 9 10 9 2
27 3 3 10 0 9 4 13 1 11 11 2 13 1 11 11 2 10 12 9 12 1 10 9 15 13 3 2
15 10 9 0 0 1 10 10 9 0 13 3 10 9 0 2
16 15 4 13 1 13 12 9 1 11 1 11 1 3 12 9 2
13 10 9 1 9 4 13 1 10 9 1 9 11 2
12 10 9 0 15 4 13 1 10 11 1 12 2
44 10 9 15 13 10 9 1 10 11 11 13 1 3 1 12 9 7 4 13 10 0 9 2 16 15 13 1 10 9 1 1 10 9 2 1 13 1 10 9 0 1 10 9 2
11 10 12 9 2 10 11 13 1 10 9 2
7 10 9 1 9 13 0 2
35 10 0 9 1 9 1 3 16 0 9 13 1 10 9 1 10 9 11 11 1 11 11 2 1 10 9 1 10 0 9 1 2 11 11 2
33 1 9 1 10 10 9 13 1 10 9 0 2 15 13 2 1 13 2 10 9 7 1 10 9 1 10 9 1 9 1 10 9 2
18 11 13 10 9 0 2 13 1 10 9 1 10 11 7 10 9 11 2
20 10 9 1 10 9 0 1 10 9 12 15 13 1 10 9 0 1 10 11 11
35 15 13 9 1 10 9 0 1 10 12 7 12 9 1 10 9 1 10 9 9 1 10 11 0 15 15 4 13 1 10 11 7 1 11 2
33 15 13 1 15 16 10 9 1 10 9 14 3 4 3 1 10 9 13 2 1 2 13 14 15 2 10 3 0 9 1 10 9 2
24 10 9 4 3 0 13 1 13 10 9 1 12 9 9 1 10 9 1 10 9 1 9 0 2
18 1 10 9 1 10 9 0 2 10 9 0 4 13 1 10 9 0 2
16 11 13 10 9 2 10 9 2 1 13 10 0 9 1 9 2
51 15 4 13 13 10 9 1 10 11 11 1 10 9 1 3 1 12 9 2 9 1 9 1 9 2 1 10 9 1 9 13 1 0 9 1 10 9 1 10 11 1 16 3 13 10 9 1 10 11 11 2
35 10 9 0 13 10 9 0 1 9 7 1 9 13 1 10 9 1 9 2 1 12 7 12 3 2 1 10 9 13 1 12 7 12 9 2
26 15 15 13 2 3 2 1 10 9 1 9 13 1 10 9 1 12 9 1 10 9 0 1 10 11 2
45 10 9 1 10 9 1 10 9 1 10 11 13 3 1 10 9 0 7 10 9 1 10 9 1 10 0 9 2 3 1 13 1 12 9 1 10 9 1 10 9 0 1 10 9 2
9 14 4 4 13 10 12 9 12 2
22 7 15 14 13 3 10 9 16 15 4 4 13 15 14 1 10 9 0 1 10 0 2
17 9 1 10 9 7 1 10 9 1 9 2 15 13 3 9 0 2
27 1 12 7 12 2 15 13 10 9 3 0 2 1 10 9 1 10 9 7 9 1 11 11 7 11 11 2
9 15 13 9 1 10 9 1 11 2
13 10 9 4 13 3 1 11 1 10 9 1 11 2
32 11 13 1 11 16 16 15 15 13 1 11 2 10 9 0 2 15 15 4 13 10 0 9 0 1 13 10 9 1 10 11 2
45 1 10 0 9 2 15 13 10 9 15 13 1 10 9 0 1 15 13 1 10 0 9 7 1 10 9 0 2 7 3 0 7 0 1 13 10 9 1 9 1 9 1 10 9 2
24 3 2 10 0 9 1 10 9 1 11 13 11 1 3 1 10 9 2 1 10 3 0 9 2
19 10 9 1 9 13 10 9 11 11 2 9 1 9 13 10 9 1 9 2
15 10 9 13 10 9 11 1 10 11 2 9 12 2 12 11
23 15 13 10 9 1 10 9 7 3 3 10 9 1 10 9 1 15 10 9 13 10 9 2
36 1 10 9 2 16 10 9 1 10 11 13 10 9 1 9 2 10 9 3 14 13 3 3 10 9 15 13 3 10 9 15 10 9 15 13 2
43 3 13 10 9 1 11 11 1 13 10 9 9 1 10 9 1 11 2 3 16 1 10 9 1 10 9 1 11 1 12 2 11 1 12 7 11 1 12 15 13 10 9 2
30 1 10 9 1 12 2 15 13 10 9 1 9 1 10 9 7 14 13 3 1 13 13 10 9 0 13 1 11 11 2
23 15 13 1 10 9 1 1 12 1 10 11 1 10 9 2 1 1 13 1 10 11 11 2
13 10 0 9 1 9 14 13 3 3 0 3 3 2
23 10 9 1 10 11 13 10 9 0 13 1 10 9 1 11 2 1 10 9 0 1 11 2
11 10 2 9 2 13 10 9 1 10 9 2
33 16 10 9 15 4 13 1 12 2 10 9 15 4 13 7 15 4 13 9 1 10 9 1 9 1 10 9 11 1 10 9 2 2
17 15 13 11 11 2 11 11 2 11 11 2 11 11 7 11 11 2
25 7 10 12 9 2 11 11 2 11 11 11 2 11 11 7 11 11 2 4 13 1 13 10 9 2
55 2 9 2 14 13 10 9 1 2 9 1 13 2 3 3 3 2 1 10 9 1 10 12 9 2 1 9 2 3 2 1 10 9 1 10 9 1 9 3 16 15 14 13 3 10 9 1 10 9 9 15 13 2 9 2
17 10 11 7 10 11 15 15 4 3 13 13 10 9 3 1 3 2
47 1 12 2 10 9 1 10 10 9 13 4 13 1 9 12 9 1 9 2 10 15 1 12 7 10 9 1 12 9 0 2 3 0 1 10 10 9 7 13 1 10 9 0 1 9 0 2
37 10 0 9 1 11 7 11 2 10 9 11 2 13 3 1 13 10 3 10 9 2 15 10 9 1 9 2 1 13 10 9 1 11 2 12 2 2
16 10 0 9 14 15 13 1 10 9 1 10 0 9 1 9 2
19 15 13 3 1 10 11 1 10 11 1 3 16 9 1 10 9 1 11 2
14 3 10 13 9 7 10 9 9 1 10 9 1 9 2
32 10 9 11 11 2 0 1 10 9 2 15 13 1 10 9 0 15 2 1 10 9 1 11 11 4 3 3 13 10 9 0 2
15 10 9 1 10 9 4 13 1 13 10 9 1 10 9 2
20 10 9 1 9 11 12 15 4 13 1 11 1 10 12 1 10 12 9 12 2
15 13 16 10 9 0 13 2 10 0 9 1 9 4 13 2
12 15 4 15 13 1 10 9 1 10 9 11 2
22 1 10 9 2 10 9 4 13 10 9 0 0 2 3 13 1 10 9 0 7 0 2
38 1 10 9 0 15 0 10 9 1 9 0 13 11 2 10 9 1 10 9 0 13 1 9 1 10 9 2 3 16 15 13 10 9 1 10 9 0 2
36 10 9 1 11 9 13 10 9 1 10 9 1 10 9 1 10 9 15 4 13 1 10 9 0 1 10 12 9 1 9 1 9 7 1 9 2
13 10 9 1 9 4 13 9 2 9 1 9 2 2
23 10 11 12 4 4 13 1 10 9 9 1 10 9 2 15 15 13 1 13 1 10 9 2
22 15 13 3 1 15 13 1 10 9 1 11 15 15 4 13 0 1 10 9 1 9 2
12 10 0 9 1 10 11 1 11 13 11 11 2
23 10 9 14 4 3 13 4 13 1 10 9 1 0 9 1 13 1 13 13 10 9 0 2
11 9 2 9 1 11 12 2 10 9 9 2
27 1 10 9 2 10 9 1 10 9 1 10 9 1 9 0 13 1 10 9 1 9 1 10 9 10 0 2
27 15 13 1 10 9 11 0 1 11 2 11 2 2 10 9 1 10 9 0 0 2 15 4 13 10 9 2
19 10 9 0 1 11 2 0 9 1 11 2 2 11 13 10 9 0 0 2
16 1 10 9 10 9 4 13 1 10 9 9 1 10 9 11 2
22 3 13 3 12 9 1 10 9 2 9 2 10 9 1 10 9 7 10 9 1 9 2
28 15 13 3 16 13 3 10 9 1 10 9 0 1 10 9 1 9 1 9 2 0 1 10 9 1 10 9 2
51 10 9 0 1 10 11 2 4 13 1 10 9 1 9 1 10 9 0 2 13 3 10 9 1 9 2 1 9 1 10 9 13 1 11 7 11 11 2 3 1 10 9 1 10 9 1 10 0 11 0 2
26 11 11 2 10 9 0 2 12 2 13 10 9 1 11 2 1 13 0 2 10 9 4 4 4 13 2
19 10 9 1 12 9 7 10 9 1 12 12 1 9 1 9 4 4 13 2
31 1 9 1 10 9 1 10 11 2 15 13 10 9 6 13 10 9 13 1 9 1 10 9 2 13 10 9 1 10 11 2
21 10 9 1 11 2 7 11 2 4 13 1 11 1 9 11 1 10 9 1 11 2
51 10 11 9 1 11 4 13 10 9 1 10 9 1 10 9 1 10 9 11 7 1 10 9 9 1 10 11 9 2 1 9 1 10 9 1 10 9 0 1 10 9 1 10 11 2 4 15 13 9 9 2
25 10 11 4 13 12 9 1 9 0 1 9 1 9 7 3 1 12 9 1 9 1 9 1 9 2
25 10 9 1 11 13 0 1 10 9 1 11 2 11 11 2 11 2 11 2 11 2 11 7 11 2
24 10 9 1 10 9 1 12 2 3 3 13 1 10 11 1 11 2 14 13 3 10 9 0 2
30 11 11 4 13 10 9 1 9 1 9 1 9 7 16 15 13 0 2 15 13 0 2 12 9 1 4 13 10 9 2
24 10 9 15 13 1 9 1 10 9 0 1 13 3 12 9 1 9 1 10 9 7 1 11 2
11 15 13 10 9 1 10 9 11 11 11 2
40 10 9 1 10 9 0 13 9 1 10 9 0 1 10 9 1 11 2 13 1 10 9 1 10 11 1 10 11 1 11 1 11 7 1 10 11 0 1 11 2
38 3 16 15 13 10 3 3 10 9 0 2 15 4 13 1 2 13 2 10 9 15 13 7 13 10 9 0 7 1 13 10 9 1 10 2 10 9 2
46 10 9 13 1 9 2 13 2 15 4 13 10 9 1 10 9 15 15 13 1 10 9 10 9 1 11 2 0 9 2 15 15 4 13 2 7 13 1 9 1 10 0 9 11 11 2
17 15 4 13 1 12 9 1 9 2 10 9 11 11 7 11 11 2
30 1 10 9 1 10 9 0 2 10 11 11 4 13 1 9 10 12 9 12 2 3 1 10 9 1 9 1 10 11 2
8 10 9 13 0 1 13 0 2
11 10 9 13 1 9 0 7 1 9 0 2
15 11 11 13 10 9 1 9 0 1 10 9 1 10 11 2
21 9 0 1 11 11 1 10 9 1 11 11 7 11 11 15 4 13 1 1 9 2
18 1 10 9 2 11 2 2 3 1 0 9 2 11 11 13 10 9 2
23 3 2 15 13 12 9 10 9 0 1 10 11 7 10 9 10 9 1 9 1 11 11 2
31 10 9 13 10 9 0 1 15 1 10 11 0 15 15 15 13 1 10 9 0 0 3 13 1 10 9 1 1 10 9 2
24 1 12 2 10 9 13 1 10 0 9 1 10 9 1 10 11 2 1 10 9 0 9 0 2
30 10 9 13 1 10 11 0 1 10 9 1 10 11 1 10 11 7 13 10 9 2 13 10 0 9 1 10 9 0 2
8 1 0 9 2 13 10 9 2
14 10 9 15 4 13 1 10 9 11 2 8 12 2 2
23 15 4 13 12 9 1 11 1 10 9 7 3 15 14 15 4 3 13 10 3 0 9 2
19 9 1 10 9 2 15 13 3 10 9 0 1 9 1 15 1 10 9 2
48 10 9 4 13 1 10 9 13 7 13 2 13 10 9 1 9 0 1 10 9 2 3 16 10 9 1 10 10 9 1 10 9 0 2 10 9 0 2 10 9 1 10 9 7 10 12 9 2
26 10 11 11 11 13 10 9 1 10 9 1 10 9 1 10 9 1 10 9 1 10 9 1 10 11 2
26 1 11 2 11 15 4 13 15 15 13 10 9 7 15 4 13 16 15 13 0 1 15 13 1 9 2
27 10 9 4 13 1 10 9 0 1 12 9 1 12 9 7 1 3 12 9 1 9 2 13 1 9 0 2
28 12 9 1 10 9 1 11 13 3 1 10 9 1 10 11 2 1 10 9 1 10 9 10 11 7 10 11 2
13 15 13 10 9 1 0 9 7 10 9 1 13 2
32 15 13 0 1 13 10 9 3 2 15 14 13 3 3 16 16 15 4 13 3 1 9 2 10 9 7 10 9 1 11 2 2
18 11 13 10 9 0 2 13 1 10 9 1 10 11 7 10 9 11 2
21 9 1 10 9 2 15 14 13 3 2 10 9 0 13 1 10 9 3 0 2 2
20 1 9 2 10 11 1 10 9 14 13 3 1 15 13 1 13 1 10 9 2
27 10 9 0 13 1 10 0 9 14 15 13 3 1 9 1 10 0 9 7 1 10 0 9 1 10 9 2
51 10 11 4 13 10 9 1 10 9 0 7 13 1 9 10 9 1 10 2 9 1 9 2 1 9 0 1 10 9 3 1 13 10 9 1 10 9 7 10 9 1 10 9 7 9 1 10 9 0 0 2
8 10 9 13 1 10 9 0 2
20 10 9 1 10 9 0 13 10 9 0 7 1 10 9 0 13 1 10 9 2
33 3 2 1 10 0 9 2 11 15 13 10 11 7 10 9 1 11 1 13 10 9 0 0 1 9 1 10 10 9 0 3 13 2
17 10 9 15 13 1 13 9 1 10 9 2 7 13 1 10 9 2
77 0 9 1 11 9 2 15 15 4 13 9 0 2 2 1 11 9 2 10 9 1 15 13 9 0 1 10 9 13 0 2 13 10 9 1 10 9 2 1 13 10 9 1 11 11 2 7 3 1 10 12 0 9 15 13 1 10 9 7 10 15 15 13 2 10 9 2 10 0 9 1 9 1 10 9 0 2
48 15 4 1 9 13 1 10 0 9 1 10 11 2 3 15 13 1 10 0 9 1 9 0 1 12 7 15 1 10 0 9 1 10 9 1 9 1 9 2 10 9 12 2 1 12 1 12 2
22 7 3 6 15 13 9 1 10 9 0 1 10 9 3 13 1 10 9 1 10 11 2
22 15 4 15 13 1 11 2 0 9 2 7 3 1 8 8 2 9 1 10 9 2 2
11 10 9 13 10 9 7 11 13 10 9 2
11 7 10 9 1 3 13 10 9 1 3 2
10 10 9 1 9 13 1 10 0 9 2
50 10 9 2 1 10 9 1 10 9 1 10 11 11 11 11 2 15 4 3 13 1 10 11 1 10 9 1 10 11 7 1 10 11 2 1 4 13 10 9 6 13 10 9 1 10 9 1 10 11 2
26 10 9 7 11 11 11 13 10 9 0 2 0 1 10 9 1 10 9 13 2 13 1 10 9 0 2
12 1 3 2 10 9 13 1 10 9 1 9 2
35 11 11 13 10 9 1 13 10 9 2 15 15 13 10 9 1 10 9 2 1 9 16 10 9 1 11 13 3 10 9 1 10 9 0 2
28 10 9 0 4 3 13 1 12 9 1 9 2 0 7 0 2 2 13 1 15 2 13 10 9 1 9 0 2
25 15 4 13 9 0 1 10 9 11 1 11 11 7 9 1 10 9 9 1 10 9 9 1 11 2
10 11 1 11 0 4 4 13 1 12 2
41 1 10 9 0 2 10 9 0 15 13 1 10 9 0 13 1 10 9 1 10 9 2 10 9 7 10 9 13 10 9 1 9 7 10 9 1 10 9 1 11 2
41 15 3 4 13 1 10 9 1 9 15 15 13 2 15 15 13 1 10 11 1 11 1 11 2 1 15 13 3 2 7 1 10 9 1 10 11 7 1 10 11 2
23 10 9 1 9 1 9 7 1 0 9 4 13 1 10 9 0 1 9 13 1 11 11 2
32 15 13 1 10 9 1 9 1 10 9 1 10 9 0 1 10 11 11 11 1 13 1 12 1 12 9 1 10 11 1 11 2
14 10 9 0 13 10 0 9 7 9 1 10 9 0 2
45 10 9 1 10 11 7 0 9 1 12 9 2 11 11 2 15 13 1 10 9 0 1 12 1 3 16 10 9 3 16 10 9 11 11 15 13 9 1 10 9 1 10 0 9 2
24 1 10 9 2 13 10 11 1 11 7 10 11 1 10 11 1 11 2 1 11 7 11 2 2
12 10 9 13 0 1 10 9 1 11 1 11 2
23 1 9 2 15 14 4 3 13 1 10 9 1 11 7 1 11 2 15 4 13 3 13 2
40 3 2 11 11 2 9 0 1 9 0 1 10 9 1 11 12 2 4 13 1 2 3 1 10 9 2 2 16 11 11 4 13 10 0 9 1 11 1 11 2
25 10 9 4 4 3 13 1 9 0 2 7 1 12 15 13 1 9 0 1 10 9 1 10 11 2
16 1 9 12 2 9 1 10 0 9 1 11 11 1 10 11 2
28 1 9 12 2 15 13 9 1 10 9 9 1 10 9 1 9 1 10 11 2 1 15 15 13 10 9 11 2
10 9 2 9 2 9 0 1 10 9 2
49 11 11 2 11 2 12 9 12 2 11 2 12 9 12 2 9 7 9 0 9 2 4 13 1 10 9 1 4 13 9 1 10 9 1 10 11 0 1 11 2 3 1 15 4 13 10 11 11 2
9 10 9 1 10 9 13 3 0 2
33 15 13 3 10 0 9 1 12 9 2 9 15 15 13 3 2 12 9 1 9 1 10 9 11 1 10 9 1 9 1 12 5 2
7 15 4 13 1 15 13 2
35 10 9 1 9 0 13 10 9 0 13 10 9 0 1 10 9 1 10 9 7 2 7 1 10 9 2 1 10 9 1 9 1 10 9 2
11 15 13 1 11 7 13 10 9 1 9 2
15 10 9 13 10 0 9 1 9 1 10 9 7 10 9 2
17 15 4 13 10 0 9 1 10 9 3 0 13 1 10 0 9 2
26 1 13 10 9 1 10 10 9 1 9 10 9 2 9 2 2 15 4 13 10 0 9 1 10 9 2
50 15 13 3 10 9 1 10 9 3 1 10 9 1 11 11 2 9 1 0 1 15 1 11 11 7 12 2 10 9 1 10 9 1 11 11 1 15 1 11 11 2 13 1 3 13 11 1 11 11 2
34 10 9 0 4 13 1 10 9 1 10 9 1 10 9 1 11 2 12 9 1 12 4 13 1 10 0 9 1 9 12 2 1 11 2
11 10 9 0 13 10 9 1 10 11 0 2
15 10 9 3 4 13 16 10 9 4 13 1 10 12 9 2
31 1 10 9 1 12 9 2 15 13 1 9 1 10 9 2 9 1 0 9 2 9 1 9 0 3 1 13 1 10 9 2
12 10 9 0 15 13 1 11 2 1 10 11 2
16 10 11 11 4 13 1 10 9 0 7 10 9 1 10 9 2
17 11 13 10 13 1 10 9 0 1 11 1 9 1 11 7 11 2
24 10 11 11 2 3 13 2 11 11 2 2 13 10 9 0 15 13 1 10 11 13 1 12 2
23 11 11 1 10 9 4 13 10 9 1 10 11 1 10 11 2 15 13 3 1 10 9 2
15 1 12 10 9 13 1 10 9 7 1 12 1 10 9 2
26 15 4 13 1 11 1 11 2 10 12 9 12 2 3 13 1 11 1 10 9 1 9 1 10 11 2
11 10 0 9 1 11 13 10 9 1 11 2
15 15 13 10 9 0 0 15 13 10 9 1 10 9 0 2
37 16 10 9 1 10 11 13 3 1 10 9 0 7 16 10 15 14 15 13 3 3 9 2 10 9 7 3 1 10 11 1 0 15 4 3 13 2
35 15 13 1 10 9 0 1 10 9 1 10 9 10 0 9 1 10 9 1 11 2 10 0 9 1 10 9 13 10 0 9 1 10 9 2
18 3 10 9 1 10 9 0 4 13 10 9 15 13 3 10 9 0 2
8 11 11 13 1 15 15 13 2
36 1 9 1 10 9 13 7 13 1 9 2 10 9 4 13 3 10 9 1 10 9 0 2 1 10 9 2 1 10 9 7 1 10 9 0 2
32 1 9 2 15 13 2 1 0 9 2 12 9 0 1 12 1 12 9 2 15 12 13 3 1 13 0 1 10 9 1 9 2
12 11 11 11 13 10 9 0 1 10 9 0 2
9 13 15 15 13 1 10 0 9 2
45 10 9 4 13 1 10 9 2 10 9 7 10 9 15 13 10 9 1 11 2 15 1 10 10 9 1 10 9 0 15 13 10 9 1 9 7 1 9 1 11 7 1 10 11 2
21 10 9 0 13 10 11 11 1 12 2 3 3 10 11 11 11 1 13 1 12 2
19 10 9 4 3 15 13 1 9 1 10 0 9 1 9 2 9 0 2 2
42 1 9 1 10 9 7 10 9 1 9 0 2 15 15 13 3 10 9 1 9 1 12 7 1 10 9 1 12 2 15 13 16 1 12 7 12 15 4 13 10 9 2
38 15 13 10 9 1 12 12 1 9 1 9 0 7 9 1 12 12 1 9 15 10 9 13 1 9 10 0 9 2 10 9 11 7 10 9 11 11 2
22 1 10 9 2 10 11 13 1 13 9 7 13 13 3 10 15 15 10 9 13 0 2
11 10 9 0 14 13 0 1 10 9 12 2
16 3 9 1 12 2 11 15 13 1 14 3 13 10 0 9 2
11 15 13 10 9 1 9 1 10 9 0 2
31 10 11 4 15 13 1 9 1 12 1 10 9 0 1 9 1 10 9 0 2 13 3 10 9 1 13 9 1 10 9 2
17 11 13 10 9 0 2 13 1 10 9 1 11 7 10 9 11 2
36 10 11 1 10 9 0 1 11 13 10 9 15 13 9 1 10 9 0 1 10 9 1 11 7 15 15 13 1 10 9 1 10 9 1 11 2
20 10 9 0 7 10 9 1 9 0 1 0 4 13 1 10 9 1 0 9 2
38 15 13 12 9 3 3 2 1 10 9 1 12 9 2 2 13 2 2 4 15 13 2 2 1 10 9 1 10 15 15 15 14 4 3 4 13 2 2
11 15 4 13 1 10 9 1 10 9 11 2
21 10 9 0 4 13 10 9 7 10 9 13 1 10 9 0 7 0 1 10 9 2
17 1 11 11 2 15 13 11 15 15 13 12 1 12 1 9 0 2
27 1 9 11 1 11 4 13 10 9 1 10 9 1 11 2 9 1 10 9 1 10 9 1 10 12 9 2
14 1 12 2 11 13 11 7 11 1 10 9 1 9 2
16 3 2 10 9 1 10 9 13 10 9 1 9 7 1 9 2
47 13 1 9 10 9 15 13 1 4 13 2 10 10 9 0 13 9 1 10 0 9 2 3 1 10 9 0 1 10 9 1 9 2 3 12 14 1 10 9 0 0 15 4 13 10 9 2
12 0 9 2 13 10 9 1 9 13 3 0 2
20 15 13 9 1 10 11 1 11 2 1 0 9 1 10 0 9 11 11 11 2
19 1 15 13 1 10 9 2 11 15 13 10 9 2 1 10 9 1 11 2
22 15 13 3 1 11 1 10 9 1 10 9 11 11 11 7 13 3 10 9 1 11 2
14 10 9 4 3 13 1 10 9 11 5 11 1 11 2
33 10 9 13 16 15 14 13 3 3 10 9 0 13 1 10 9 0 1 10 9 1 10 9 2 7 2 3 2 1 10 0 9 2
16 3 1 9 7 1 0 9 2 15 13 10 9 1 10 9 2
20 4 15 13 15 4 4 13 1 9 12 7 4 13 1 9 10 12 9 12 2
27 15 13 3 16 10 9 11 13 10 9 1 10 9 2 2 3 13 11 16 15 14 15 13 3 1 11 2
21 10 9 4 13 1 10 9 0 15 15 13 2 7 1 10 9 0 15 15 13 2
33 13 9 10 12 9 12 1 10 9 1 11 2 15 13 10 9 1 10 9 1 11 15 15 13 9 7 9 1 10 9 7 9 2
18 15 4 3 13 16 1 10 9 2 15 13 10 9 15 13 10 9 2
11 10 3 3 0 9 15 15 13 1 15 2
42 9 1 10 9 1 10 9 0 2 1 9 7 1 9 2 9 1 10 9 0 7 0 9 1 10 9 2 15 13 10 9 0 1 10 9 15 13 1 15 10 9 2
23 16 15 13 9 1 13 1 10 9 15 10 9 13 1 13 2 15 15 13 3 10 9 2
31 15 13 3 2 1 10 9 1 10 9 1 11 2 1 13 10 9 1 10 9 0 7 10 9 1 10 9 0 1 11 2
10 15 4 13 1 10 9 0 11 11 2
36 3 1 10 9 1 11 11 15 13 10 9 1 0 9 1 10 9 1 10 9 1 9 1 9 2 11 11 4 4 13 9 1 10 9 0 2
5 15 4 15 13 2
29 10 9 1 11 13 10 9 0 1 9 0 13 1 10 0 9 1 9 1 10 0 9 1 11 7 10 9 11 2
9 7 15 13 10 9 1 10 9 2
19 1 9 1 9 1 12 9 2 10 0 9 1 9 13 10 9 1 9 2
31 10 9 15 13 1 10 9 1 10 9 1 11 1 15 15 13 10 9 1 11 2 11 1 10 9 7 11 1 10 9 2
71 3 13 3 10 0 9 1 10 9 1 10 11 2 3 0 1 9 0 9 1 10 11 11 2 3 16 1 10 0 9 15 10 11 7 10 11 2 2 7 13 1 10 9 15 15 13 13 1 15 13 1 10 9 0 1 3 1 12 12 1 9 2 1 10 9 1 10 9 15 13 2
32 7 3 10 9 0 13 1 10 9 2 10 11 1 9 0 2 10 11 0 7 3 10 11 1 9 1 10 9 13 10 9 2
14 3 15 13 10 9 3 0 2 12 9 1 11 2 2
21 1 9 4 15 13 10 9 2 16 15 13 1 13 10 9 1 10 9 1 11 2
33 1 10 9 1 12 9 15 13 10 9 3 1 13 7 1 13 10 3 0 9 1 10 9 2 9 2 9 2 9 2 9 2 2
18 3 16 10 9 13 0 2 7 10 9 14 15 4 3 13 13 2 2
29 15 13 1 3 16 9 1 10 9 16 15 15 13 1 10 9 1 11 1 12 2 13 10 9 1 11 1 11 2
13 10 9 13 0 2 0 7 10 9 13 3 0 2
17 11 14 4 15 3 13 10 0 9 1 13 10 9 1 10 9 2
22 10 0 9 0 1 10 9 11 4 13 1 11 1 11 1 10 9 1 10 9 12 2
9 2 15 4 13 1 13 12 9 2
28 15 4 13 9 0 1 10 9 0 9 1 9 13 1 11 11 7 11 11 2 11 11 2 11 12 2 12 2
18 10 9 1 10 9 15 13 1 10 11 1 9 7 1 9 1 11 2
18 15 13 3 13 3 10 9 9 15 13 1 10 9 1 10 9 9 2
26 15 2 3 16 10 9 13 15 1 13 11 7 13 11 1 10 9 1 16 10 9 13 1 0 0 2
16 15 13 1 9 10 0 9 1 11 1 10 9 1 10 11 2
27 1 12 2 11 11 13 10 9 1 10 0 9 11 11 10 11 2 12 9 2 2 7 15 13 10 11 2
13 10 9 1 9 1 11 4 3 13 4 3 13 2
15 15 13 15 15 13 10 9 1 11 2 10 9 11 11 2
7 10 9 3 13 3 0 2
22 9 0 16 10 9 1 9 13 10 12 9 1 10 9 12 9 1 4 13 1 9 2
42 15 13 3 10 9 1 10 9 0 2 10 9 1 10 9 1 11 2 1 10 9 11 11 2 15 15 13 10 11 1 11 11 11 2 2 11 11 7 11 11 11 2
15 10 9 0 1 9 13 10 9 0 7 0 0 1 9 2
47 1 12 2 15 13 10 9 11 11 11 1 11 2 1 10 9 1 10 9 2 1 9 1 10 9 1 10 9 1 10 9 1 10 9 0 2 1 10 9 7 1 1 10 3 10 9 2
26 10 9 1 11 13 10 9 1 9 0 1 10 10 9 2 15 13 1 10 9 1 10 9 1 9 2
31 11 13 10 9 0 1 9 1 10 9 0 2 9 13 1 10 9 7 10 9 0 7 10 0 9 0 1 10 0 9 2
10 15 4 13 1 1 9 1 9 16 3
53 3 9 0 7 9 13 1 12 2 10 9 1 9 2 11 11 2 9 9 9 9 2 13 15 3 10 9 13 1 12 2 2 10 9 4 15 13 1 10 9 7 4 13 12 9 13 1 10 9 3 1 13 2
27 15 13 10 9 1 10 9 2 3 10 9 1 9 2 7 15 13 1 15 13 16 3 15 13 1 11 2
35 1 1 15 15 15 4 13 2 15 15 13 10 9 10 0 9 3 0 7 15 13 3 3 0 1 13 1 10 9 13 1 10 11 0 2
21 10 9 0 7 11 11 13 10 9 1 9 15 15 15 13 1 10 9 1 9 2
83 11 13 3 10 0 9 0 2 11 11 11 2 12 2 2 9 1 10 9 1 11 2 12 2 2 9 0 1 11 2 12 2 2 9 1 10 9 1 11 2 12 2 2 7 3 0 2 9 1 10 9 0 1 10 9 1 9 0 1 10 9 1 11 2 12 2 2 9 1 9 2 12 2 2 9 0 2 11 2 12 2 2 2
10 10 9 4 13 1 13 10 9 0 2
23 10 9 0 4 13 1 10 11 1 11 7 1 11 15 2 3 2 13 10 9 9 0 2
9 15 15 3 13 3 10 9 1 9
20 10 11 0 7 10 11 1 11 4 13 1 10 11 0 7 11 10 12 9 2
14 15 13 10 9 3 1 13 10 9 1 9 1 9 2
21 3 2 10 9 13 10 9 1 10 11 0 15 15 13 1 9 1 10 9 0 2
29 10 9 0 1 10 8 2 9 5 13 10 9 1 8 15 2 1 0 9 2 13 1 5 10 9 1 9 1 8
17 10 9 1 10 9 5 14 13 0 1 10 9 1 9 1 9 2
23 10 0 9 1 10 9 13 3 1 10 9 1 10 9 2 15 1 10 9 0 1 9 2
42 10 9 8 11 2 12 9 2 10 3 0 1 10 9 1 10 9 11 11 2 13 10 9 1 9 1 12 5 2 1 10 9 13 9 1 10 9 1 9 0 11 2
9 15 13 10 9 1 9 1 12 2
13 15 4 13 10 11 11 7 15 15 4 13 2 2
25 15 13 10 9 0 1 11 7 1 11 1 10 11 7 13 1 10 9 10 9 1 10 9 0 2
28 10 9 1 9 1 10 9 13 3 0 1 15 1 10 9 2 12 2 7 1 15 1 10 9 2 12 2 2
12 10 9 0 13 10 9 1 9 2 13 9 2
20 10 9 7 10 9 1 10 9 1 10 9 13 10 9 0 1 10 0 9 2
25 15 13 10 15 1 10 12 0 9 1 10 11 1 10 9 1 10 9 0 1 11 7 1 11 2
24 9 7 9 0 1 9 0 2 11 11 13 1 11 10 0 9 0 1 10 9 1 11 11 2
30 15 4 13 2 10 12 9 12 2 9 1 10 11 1 11 2 1 10 9 1 10 9 1 10 9 0 2 11 11 2
19 10 0 7 0 9 7 9 15 13 2 7 14 13 3 1 13 10 9 2
14 10 9 0 15 13 3 1 10 9 7 10 0 9 2
19 15 13 0 1 13 10 15 1 9 2 7 1 13 10 9 0 7 0 2
34 1 10 9 1 12 1 11 11 2 10 9 0 4 13 1 9 0 1 1 15 16 10 9 1 10 9 4 13 1 10 11 1 12 2
8 10 9 13 3 0 7 0 2
8 15 13 10 0 9 1 9 2
23 11 2 11 1 9 2 13 10 9 0 2 13 1 10 9 1 10 11 7 10 9 11 2
16 1 12 2 11 13 10 9 11 11 2 3 1 1 11 11 2
20 15 13 3 16 15 13 10 9 1 10 9 1 15 13 3 1 10 9 0 2
35 10 9 4 3 15 13 1 1 9 2 7 3 10 3 9 1 10 9 4 13 16 15 15 4 13 3 10 9 3 0 1 9 1 9 2
13 10 9 2 9 0 7 0 13 3 0 1 11 2
45 13 9 1 12 2 15 13 9 1 11 11 1 10 9 1 12 3 9 1 10 9 11 1 10 9 10 12 9 12 1 10 9 1 9 1 10 9 1 10 0 9 1 11 11 2
18 15 15 13 3 16 10 11 7 10 9 1 10 11 14 13 3 12 2
20 10 9 4 13 1 4 13 10 9 1 9 1 10 9 1 10 9 1 11 2
30 1 12 2 15 13 12 9 1 11 13 1 9 1 9 0 2 2 9 9 2 2 1 10 9 1 9 1 10 9 2
20 15 15 13 1 10 9 2 7 11 0 15 13 3 2 13 10 9 1 11 2
20 1 9 11 4 13 10 9 1 10 9 1 10 9 10 9 1 0 11 9 2
25 3 2 1 0 1 10 9 15 13 1 10 9 2 15 15 15 13 1 13 1 10 3 0 9 2
19 13 1 10 0 9 15 15 13 3 13 1 10 9 10 0 9 1 13 2
22 15 15 13 3 10 9 1 10 9 13 10 0 7 10 9 7 10 9 1 10 9 2
17 15 4 13 13 10 9 1 9 1 9 2 7 10 9 13 0 2
18 15 4 13 10 12 9 12 1 10 9 11 11 11 15 15 13 0 2
31 10 9 13 1 10 9 1 10 9 2 10 9 1 10 9 1 0 7 10 9 0 1 10 9 0 2 4 13 10 9 2
26 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 10 9 2 3 1 9 7 1 9 2
29 10 12 9 12 2 11 11 11 4 13 11 1 10 9 1 10 9 0 2 9 15 15 13 1 10 12 9 12 2
23 15 13 1 3 10 9 3 0 1 14 3 13 0 1 11 9 1 10 11 1 10 11 2
27 1 10 9 1 9 2 15 13 3 3 10 0 9 1 10 9 1 10 9 16 15 3 13 13 10 9 2
12 10 9 0 13 0 1 9 1 10 9 11 2
32 1 10 9 11 11 2 2 10 9 1 10 9 1 10 11 2 1 11 2 1 11 7 1 11 13 10 9 1 10 9 2 2
10 10 9 4 13 1 11 11 7 11 11
14 10 9 13 3 10 9 1 9 0 1 10 9 0 2
12 10 9 15 4 13 10 9 14 4 3 13 2
34 7 10 9 15 2 3 13 10 0 9 15 13 1 10 9 2 1 10 9 0 2 15 13 10 9 1 10 9 0 1 10 9 0 2
7 3 2 10 9 13 3 2
19 13 1 12 2 10 9 4 13 1 10 9 0 1 10 9 1 10 11 2
25 15 4 13 10 9 1 10 9 8 13 1 10 11 11 11 2 3 16 1 10 9 1 11 11 2
13 15 4 13 10 12 9 1 10 9 1 11 11 2
31 10 9 4 13 1 15 7 13 10 9 15 13 10 9 7 10 9 2 1 10 9 1 13 10 9 1 10 9 1 9 2
18 3 12 9 3 3 2 10 0 9 4 13 1 1 10 9 1 11 2
21 10 9 13 1 10 12 9 7 13 0 1 10 9 1 10 11 2 1 10 9 2
24 3 2 10 9 2 0 2 2 15 4 13 1 10 9 1 10 9 0 1 12 2 13 11 2
14 11 11 13 10 9 1 9 1 10 9 1 10 11 2
16 15 14 15 13 3 1 10 9 7 1 10 9 1 9 2 2
19 10 9 4 13 1 9 1 10 9 9 2 13 1 9 1 9 1 9 2
18 13 15 3 1 10 9 1 10 9 2 10 11 2 1 12 9 12 2
24 10 9 1 9 0 13 3 1 0 10 9 1 10 9 1 0 2 13 10 9 1 9 2 2
11 10 9 11 12 15 13 10 9 1 9 2
17 10 9 13 3 12 9 0 1 11 11 2 11 11 7 11 11 2
29 10 9 1 11 4 13 3 1 9 0 1 10 9 1 11 13 1 10 11 2 1 12 7 12 12 1 9 2 2
28 1 10 0 9 0 1 11 2 11 13 10 9 7 15 13 1 10 9 15 15 13 1 10 9 1 10 9 2
34 1 10 9 1 10 9 11 1 11 2 15 13 10 9 1 9 1 10 9 1 10 9 1 10 0 9 7 13 0 9 1 10 9 2
9 15 13 10 9 7 13 10 9 2
28 1 10 9 1 10 12 9 2 10 9 0 2 4 4 13 1 10 12 9 12 9 13 1 10 0 9 0 2
32 1 9 0 1 10 12 9 12 10 9 1 9 1 11 2 1 11 2 11 7 11 4 13 1 13 10 9 1 9 1 11 2
11 10 11 13 10 0 9 0 7 9 0 2
16 3 13 1 10 9 12 2 10 9 12 9 0 1 10 11 2
19 15 15 13 3 1 10 9 0 2 1 10 9 7 1 10 9 0 0 2
13 1 9 1 12 15 13 1 10 9 1 9 0 2
23 15 4 3 13 1 13 10 9 1 10 9 9 9 11 11 2 3 0 1 10 9 12 2
42 1 9 2 10 9 9 4 2 4 13 1 10 9 1 10 9 2 15 14 13 3 1 10 9 2 0 2 1 10 9 7 14 13 3 3 1 10 9 1 10 9 2
35 15 15 13 1 11 7 3 2 13 1 10 9 13 1 10 9 1 15 13 1 10 0 9 1 10 9 15 14 13 3 1 15 15 13 2
29 13 10 9 0 2 15 13 10 9 1 10 9 13 1 10 9 11 11 1 13 7 13 3 10 15 1 10 9 2
15 12 1 12 9 13 0 1 13 10 10 9 1 10 9 2
15 10 9 4 15 13 1 13 10 9 15 10 9 4 13 2
37 10 9 0 1 10 9 1 10 9 4 13 10 9 9 1 10 9 1 10 9 0 1 11 11 2 9 1 10 9 0 1 10 9 1 10 9 2
27 10 9 0 4 13 1 11 11 2 15 4 13 1 12 9 1 10 9 11 7 13 1 10 11 1 11 2
10 9 0 2 15 3 13 3 1 9 2
16 10 9 1 10 9 13 10 9 1 10 9 15 13 10 11 2
25 11 1 11 2 9 1 10 11 1 11 2 3 13 1 10 9 10 9 1 10 9 12 3 12 2
40 1 10 12 9 1 10 9 1 11 11 2 10 11 14 4 3 13 10 9 0 7 4 13 10 9 15 13 1 9 10 9 0 0 15 10 0 9 4 13 2
12 15 13 3 9 1 10 11 1 13 10 9 2
22 11 4 13 10 9 0 1 10 9 15 4 13 10 9 2 3 1 11 7 1 11 2
31 11 15 4 13 1 13 10 9 1 10 9 1 10 0 9 1 15 13 1 10 0 9 11 1 10 9 11 12 3 13 2
21 10 9 4 13 1 10 9 1 9 9 3 13 2 13 1 9 7 13 1 9 2
26 9 1 9 0 2 10 11 1 12 9 4 3 13 1 15 13 1 10 9 1 10 9 9 11 11 2
18 1 12 2 12 5 1 10 9 13 1 9 0 7 12 5 13 0 2
55 3 2 11 11 13 10 9 0 3 0 1 13 13 10 9 7 15 13 10 9 3 1 10 9 0 2 7 1 12 10 11 11 13 1 13 10 11 2 1 0 7 0 9 1 10 9 1 10 11 7 1 10 11 2 2
9 10 9 11 15 13 1 12 9 2
19 15 15 13 1 10 0 13 1 9 2 9 13 10 3 0 1 10 11 2
13 15 4 13 12 9 1 9 1 13 10 12 9 2
15 3 10 9 0 15 13 1 9 1 11 2 1 9 12 2
20 9 13 1 10 9 1 9 1 13 10 9 3 13 7 3 13 1 10 9 2
17 10 9 15 13 1 13 1 9 1 10 0 9 2 0 7 0 2
13 10 0 9 1 13 10 9 1 9 11 1 11 2
16 10 9 9 13 10 9 13 1 10 9 1 9 7 1 9 2
9 15 13 10 9 1 9 1 12 2
15 15 4 13 0 9 0 1 10 9 12 1 10 11 11 2
19 12 0 9 0 0 13 0 1 10 9 2 1 10 9 1 10 9 0 2
22 11 15 13 1 10 9 1 10 9 1 9 7 10 9 1 13 10 0 9 1 9 2
44 11 13 3 1 9 10 9 1 9 1 10 9 1 9 2 1 13 10 0 9 1 10 9 7 10 0 9 1 9 2 13 3 1 11 11 1 13 10 9 1 11 1 11 2
11 1 12 2 15 13 1 10 9 0 0 2
29 13 3 1 13 1 10 3 12 9 1 10 9 1 10 9 1 9 7 12 9 1 10 9 1 10 9 1 9 2
15 10 0 9 13 1 10 9 4 13 10 9 1 10 9 2
32 15 15 13 3 9 16 10 9 4 13 1 10 9 7 13 3 16 10 9 4 13 1 10 9 2 1 9 1 10 9 11 2
48 1 12 10 9 11 2 9 1 9 2 2 1 10 9 1 10 9 11 11 7 11 11 11 2 4 13 10 9 1 9 0 1 9 2 11 11 2 15 13 1 10 9 1 9 1 10 9 2
29 1 10 9 9 2 10 9 14 13 1 9 16 10 9 13 7 10 0 9 1 10 9 4 13 1 10 9 0 2
10 15 15 13 1 10 9 1 12 9 2
30 10 9 11 11 2 13 10 12 9 12 1 11 7 13 1 10 9 1 11 10 12 9 12 2 13 10 9 0 0 2
15 3 1 10 9 4 3 13 1 10 0 9 1 10 9 2
18 10 9 0 4 13 10 9 1 13 10 9 1 10 11 7 10 11 2
11 15 13 10 9 15 13 9 1 10 9 2
37 11 11 11 13 10 9 1 11 11 2 9 1 10 9 1 9 1 10 11 0 2 9 1 10 11 1 11 7 1 11 2 7 1 11 11 11 2
19 10 9 4 4 13 13 10 9 1 10 9 1 10 9 1 10 9 0 2
23 10 9 9 1 10 11 1 10 9 11 13 1 9 10 11 7 10 9 1 9 1 9 2
30 15 13 1 15 13 10 9 1 9 1 10 9 0 2 13 1 10 9 2 13 13 10 9 10 9 0 1 10 9 2
17 10 9 13 10 9 0 0 1 10 11 2 4 13 10 0 9 2
39 1 9 12 2 15 13 10 9 1 9 0 1 9 2 11 2 1 10 11 1 11 2 15 15 13 10 9 1 9 0 1 2 10 9 0 1 9 2 2
93 10 0 9 13 12 9 13 3 1 10 9 1 10 9 0 1 9 1 10 12 0 9 1 9 1 10 9 2 15 12 13 1 9 2 15 1 2 9 8 2 2 2 3 16 10 0 9 13 10 9 13 3 1 10 9 1 10 9 1 12 3 12 9 15 15 4 13 1 12 2 15 12 0 1 10 9 1 10 9 0 2 13 1 0 11 2 11 15 13 1 12 9 2
10 7 15 4 3 15 13 1 10 9 2
37 10 12 4 13 1 10 9 1 9 11 2 10 9 1 11 11 13 1 11 11 7 13 10 9 15 10 9 1 9 4 13 7 13 1 10 9 2
15 10 12 9 2 11 11 7 10 9 11 11 3 4 13 2
28 10 11 15 13 3 1 10 9 1 10 9 1 13 1 9 10 9 1 12 9 7 1 13 10 9 0 0 2
34 10 9 4 3 13 1 10 9 2 3 16 10 10 9 13 1 10 0 2 9 2 9 1 9 7 9 1 1 10 9 0 1 11 2
22 11 13 10 9 1 11 1 10 9 0 1 10 9 1 11 2 1 10 9 1 11 2
22 15 13 10 9 1 10 9 1 10 9 0 0 7 13 10 9 1 9 0 7 0 2
18 15 13 1 10 9 1 10 9 1 10 9 2 3 1 13 1 12 2
9 10 9 1 10 9 1 9 13 2
9 10 9 13 10 9 1 10 9 2
36 10 9 1 10 9 4 13 1 10 9 7 10 9 2 1 10 9 2 10 11 4 13 10 9 1 9 0 7 13 10 9 7 10 9 0 2
37 1 10 9 1 15 2 11 13 16 10 0 9 13 1 13 10 9 2 1 13 10 9 1 1 15 16 10 9 4 13 1 11 7 1 10 11 2
51 10 11 1 11 4 13 1 9 9 2 5 12 5 2 2 13 10 9 1 10 12 9 2 1 10 9 13 1 10 0 9 1 11 11 2 10 9 1 10 9 0 7 10 9 0 13 9 1 10 9 2
42 1 10 9 1 10 9 2 11 11 13 10 9 1 9 1 3 12 12 1 9 3 13 1 11 2 15 13 3 12 5 1 10 9 3 16 11 13 10 12 5 0 2
19 15 13 3 16 1 12 9 2 15 13 10 3 0 9 13 1 12 9 2
30 10 9 4 13 1 11 11 2 9 0 1 10 9 12 7 12 2 15 15 13 1 10 9 1 10 9 2 11 11 2
5 9 1 11 1 9
6 3 13 7 13 15 2
38 10 9 11 11 2 12 2 2 9 1 10 9 1 11 2 4 13 1 4 13 10 0 9 1 10 9 1 11 11 2 10 2 11 1 11 2 2 2
17 1 10 0 9 2 10 9 0 13 10 0 9 7 13 10 9 2
12 15 13 2 1 15 2 10 0 9 1 11 2
28 15 13 10 9 1 9 1 10 11 1 11 1 10 9 1 10 9 2 1 10 9 1 10 9 1 11 11 2
23 10 9 12 1 10 9 1 11 1 9 13 10 12 9 1 10 9 1 0 9 1 11 2
24 13 1 11 2 1 10 9 1 10 11 2 10 12 9 12 2 13 1 10 0 9 1 12 2
14 10 9 4 4 13 1 10 9 9 1 9 1 12 2
21 16 10 9 4 13 1 11 11 2 10 9 2 1 9 0 2 4 13 1 9 2
14 11 12 15 13 1 12 1 10 9 2 11 1 11 2
50 3 16 10 9 1 10 9 15 4 13 1 10 9 1 10 9 1 10 11 10 9 13 1 4 13 7 15 15 13 3 1 10 0 9 0 13 1 10 9 1 10 11 11 1 10 9 1 10 9 2
7 10 0 9 13 11 11 2
20 10 9 1 10 11 15 13 9 7 9 1 10 0 7 0 9 1 10 9 2
8 10 9 4 13 1 9 12 2
24 10 9 1 10 9 1 3 0 9 13 3 10 9 1 10 9 0 1 10 9 1 9 0 2
18 10 9 0 1 10 11 13 9 1 11 12 9 3 1 12 7 12 2
12 1 10 0 9 15 13 11 11 7 11 11 2
19 1 10 9 1 10 9 2 10 9 15 13 1 10 9 1 10 9 0 2
21 1 9 1 9 2 10 9 0 1 10 11 11 11 1 11 11 13 9 1 9 2
22 15 13 3 10 9 1 9 0 2 0 1 13 1 10 9 10 9 7 10 9 0 2
11 15 13 3 3 1 9 1 10 9 0 2
61 1 11 11 2 10 9 1 11 13 1 10 9 0 1 9 0 1 10 9 1 9 0 2 1 10 10 1 10 0 9 7 10 9 1 10 0 9 1 11 2 7 13 1 10 9 1 11 2 10 9 15 4 13 1 9 3 12 9 3 3 2
67 3 16 3 13 1 10 9 9 3 3 0 2 3 0 3 0 7 0 2 15 13 10 9 1 9 3 0 7 10 9 3 3 13 2 3 16 10 9 1 9 7 10 9 0 1 10 9 13 2 10 9 1 9 1 10 11 15 13 1 10 9 1 10 9 9 2 2
20 15 13 10 9 1 10 9 11 11 2 10 9 0 1 10 9 1 11 11 2
46 3 15 13 15 2 13 4 15 2 10 11 2 11 1 10 11 2 15 15 4 13 1 10 9 1 4 13 9 7 9 2 1 13 10 9 2 10 9 2 10 9 13 1 10 9 2
17 10 9 1 9 15 4 13 10 9 1 10 0 9 0 1 11 2
26 10 9 1 9 9 1 10 11 13 10 9 2 11 13 3 1 12 9 1 9 7 10 11 13 12 2
16 1 10 9 9 0 13 1 12 2 15 13 10 0 9 0 2
19 9 1 14 3 13 1 9 10 9 1 9 3 0 15 4 13 10 9 2
53 3 15 13 10 9 1 10 9 1 9 2 10 9 1 9 7 1 9 2 10 9 2 10 9 2 10 9 0 0 2 10 9 1 9 2 10 9 0 0 0 7 10 9 0 2 9 2 9 2 9 0 2 2
24 10 9 11 12 13 10 9 13 1 10 9 11 2 1 10 9 1 10 11 2 1 10 11 2
45 10 9 1 12 9 13 9 9 1 10 9 1 9 1 11 2 11 1 11 2 7 13 1 10 9 11 1 11 2 13 3 1 10 2 9 0 2 10 9 2 1 10 9 0 2
15 15 15 4 13 1 15 13 1 0 11 11 1 15 13 2
17 11 11 11 2 13 10 12 9 12 2 13 10 9 0 1 9 2
25 15 13 10 0 9 1 10 9 0 1 11 2 13 11 11 11 11 2 15 13 10 9 1 12 2
24 10 9 4 13 10 9 0 1 10 11 11 2 9 1 10 9 11 11 15 13 1 10 11 2
49 10 12 9 1 10 11 11 11 2 13 1 10 11 1 10 9 7 1 10 9 1 10 9 7 13 10 9 0 13 1 10 9 1 10 9 12 2 15 4 13 10 1 10 11 11 1 11 11 2
22 15 15 13 10 9 1 10 9 1 9 7 10 9 1 10 9 1 9 9 1 9 2
45 11 13 10 9 1 10 9 0 1 11 11 2 13 1 10 9 1 11 11 7 10 9 1 11 2 10 9 1 10 9 1 11 1 10 9 0 1 11 1 10 9 1 10 9 2
17 13 1 12 1 11 11 2 11 15 13 3 10 0 9 0 0 2
11 10 9 0 13 2 4 15 3 13 9 2
28 15 15 13 1 13 10 9 1 10 11 11 2 11 11 2 1 12 9 2 12 9 2 12 9 7 12 9 2
10 10 9 13 1 12 9 2 12 2 2
12 15 13 3 3 10 9 2 10 0 11 11 2
21 15 13 1 10 9 0 0 1 9 1 9 12 2 3 0 7 3 13 1 9 2
17 10 9 13 1 10 9 0 1 10 9 2 13 1 11 7 11 2
13 9 2 11 4 13 1 9 0 10 12 9 12 2
14 12 9 13 1 10 9 2 12 0 7 12 0 2 2
32 10 0 9 0 2 13 1 9 1 11 1 10 11 2 13 1 10 0 9 10 0 9 2 10 0 9 7 10 9 1 9 2
23 3 2 10 9 0 1 9 0 4 13 1 10 9 1 11 0 2 1 13 10 9 0 2
19 15 3 4 13 1 10 9 10 9 12 9 12 2 7 15 4 4 13 2
21 10 9 13 10 9 15 13 1 12 1 12 9 0 7 4 3 15 13 1 15 2
14 10 11 1 10 11 1 11 13 10 3 0 9 0 2
41 1 10 9 0 1 10 12 9 12 2 15 15 13 1 10 15 1 10 12 9 1 10 11 1 10 9 1 11 2 7 13 3 1 9 2 16 10 0 0 9 2
22 3 2 15 13 1 13 10 0 9 3 16 10 9 14 4 3 13 7 3 1 9 2
6 10 11 4 13 9 2
21 1 10 9 0 2 10 9 15 13 0 2 2 15 15 13 3 7 3 1 9 2
36 2 10 9 1 10 9 13 1 10 9 1 0 9 7 1 3 1 9 1 10 9 2 2 4 13 2 1 10 9 2 10 9 1 9 0 2
23 1 9 7 1 15 2 15 13 10 9 1 9 15 10 9 14 13 3 1 10 0 9 2
18 15 3 13 1 13 1 9 1 10 9 1 10 9 1 10 9 11 2
10 11 7 13 10 9 1 10 10 9 2
31 10 11 12 13 10 9 1 9 0 1 0 9 3 0 13 1 10 11 2 11 11 1 10 9 1 10 11 11 11 11 11
29 10 9 0 15 13 15 3 1 10 0 9 1 10 9 1 10 9 7 10 9 0 15 13 3 10 9 1 11 2
29 1 9 2 10 9 1 10 9 0 13 16 10 9 15 4 1 13 0 7 1 10 9 1 10 9 15 15 13 2
39 10 0 9 13 1 0 9 1 10 9 1 9 2 10 0 9 2 10 0 9 1 9 13 10 12 16 15 15 13 1 10 9 13 1 10 9 1 9 2
24 1 9 2 1 10 9 1 9 2 10 9 0 13 10 15 1 10 9 1 9 1 12 9 2
11 10 9 13 10 3 0 1 10 0 9 2
24 1 10 9 1 10 9 0 2 1 12 2 10 9 1 10 9 1 11 13 3 0 1 3 2
22 10 9 2 15 4 15 13 9 9 2 15 13 10 9 1 10 0 9 9 1 9 2
53 10 9 13 15 13 1 10 9 2 9 1 10 9 1 11 1 10 9 1 11 2 11 2 11 2 11 2 11 2 11 2 11 11 1 11 2 11 2 11 2 11 2 11 2 11 11 1 11 7 11 1 11 2
20 10 9 1 10 9 15 13 1 10 12 9 1 10 9 1 10 9 1 9 2
10 15 4 3 13 9 1 10 9 0 2
16 11 1 11 13 10 9 1 11 2 1 10 9 0 1 11 2
53 1 10 9 1 10 0 9 2 10 9 15 13 1 2 11 11 11 2 2 10 9 1 11 11 2 7 15 14 13 3 1 10 9 0 9 1 11 2 13 3 1 12 9 3 1 10 9 11 1 11 11 2 2
40 10 9 1 11 15 13 1 10 9 1 10 9 1 11 2 1 10 9 1 10 11 2 1 3 12 9 1 10 9 1 11 2 12 9 1 11 7 1 11 2
29 15 15 13 1 10 9 0 13 1 10 9 1 9 2 13 3 1 13 1 9 2 13 1 10 9 1 10 9 2
38 10 9 0 1 10 9 13 1 12 2 16 10 9 1 10 11 0 11 11 4 13 9 1 10 9 1 13 1 9 10 9 0 1 13 1 9 0 2
40 3 3 10 9 1 9 1 10 9 0 1 10 11 7 0 1 10 11 2 3 16 10 0 9 0 0 15 15 13 1 9 3 3 0 2 14 4 3 13 2
19 10 9 4 13 0 3 2 7 15 13 16 15 13 0 1 10 9 0 2
40 13 10 9 1 10 9 0 0 1 12 2 15 1 10 0 9 1 10 0 11 2 15 4 13 2 3 2 1 10 9 0 2 9 0 2 1 10 0 9 2
20 1 10 12 1 10 12 9 12 2 10 0 9 1 11 4 13 1 9 9 2
31 3 1 10 9 1 10 9 2 10 9 1 9 1 9 1 10 9 4 13 10 12 9 10 9 1 9 1 10 9 0 2
25 10 9 0 1 9 0 4 3 3 13 1 10 9 0 2 7 10 9 13 3 9 6 15 13 2
16 15 13 2 13 1 9 1 9 1 10 9 2 10 9 0 2
11 15 15 13 10 9 1 9 1 10 9 2
15 10 11 13 10 9 1 10 9 1 10 11 0 1 10 11
39 11 11 2 13 10 12 9 12 1 11 2 11 2 2 13 10 0 9 0 2 15 13 1 10 9 1 9 1 9 1 10 11 11 7 1 9 1 11 2
46 10 9 9 4 13 1 10 9 1 11 11 1 11 2 11 2 2 10 9 1 10 11 4 9 1 10 11 0 1 10 11 2 11 2 2 7 10 9 1 10 11 4 9 1 11 2
9 11 13 10 9 3 1 9 1 2
24 10 0 9 2 10 11 11 13 1 10 0 9 10 9 1 10 12 5 1 10 9 0 13 2
19 1 12 2 15 13 10 9 0 15 10 9 4 4 13 1 13 10 9 2
17 9 0 2 9 0 7 0 2 10 0 9 1 15 7 10 9 2
44 3 1 9 1 9 15 13 10 9 7 3 10 9 0 3 16 1 9 15 15 13 3 1 10 0 9 3 3 0 7 15 13 10 9 0 1 9 1 9 1 10 0 9 2
26 15 4 13 10 9 1 10 2 0 2 9 9 2 15 13 3 0 2 7 15 15 4 3 3 13 2
36 10 9 11 2 3 1 9 10 0 9 2 4 13 1 9 1 12 5 1 12 9 2 1 4 10 9 13 10 3 0 9 1 10 12 9 2
11 11 4 13 1 10 11 1 10 9 0 2
37 10 9 1 10 11 11 2 13 3 1 10 9 1 9 1 10 9 1 10 9 7 0 1 10 9 0 2 4 3 15 13 1 10 11 11 12 2
20 10 9 13 10 9 1 10 9 1 10 9 2 10 9 11 11 2 12 2 2
19 10 9 1 10 9 13 0 2 15 10 9 1 10 9 13 10 9 13 2
29 10 9 1 9 13 1 10 9 1 9 1 12 9 1 12 9 13 1 10 9 13 10 9 13 1 11 12 9 2
17 10 0 9 0 13 10 11 1 11 1 10 9 1 10 9 12 2
15 10 9 0 2 10 9 1 9 1 10 9 15 4 13 2
26 11 13 10 0 9 1 10 9 0 10 12 9 12 2 1 10 9 0 9 9 11 7 9 9 11 2
33 15 4 13 10 9 2 10 9 0 2 10 9 1 9 1 9 0 2 10 9 3 16 10 9 2 3 0 1 10 9 11 2 2
29 10 0 9 1 10 11 2 10 9 1 10 11 2 13 10 9 1 10 3 0 9 1 10 9 7 13 10 9 2
36 11 11 2 10 9 1 10 9 13 9 1 11 2 7 9 1 10 11 1 11 7 10 9 1 9 2 4 13 10 9 1 10 9 11 11 2
14 1 3 9 2 10 9 1 9 13 0 7 3 0 2
39 1 9 1 10 9 2 3 0 2 15 4 13 1 10 9 1 10 9 0 13 1 10 11 1 11 7 1 10 9 1 10 9 0 1 10 9 1 11 2
12 1 12 2 15 13 10 9 1 0 9 0 2
31 11 2 1 9 0 2 2 2 1 9 10 9 2 13 10 9 13 1 10 9 1 11 1 11 2 10 9 1 10 11 2
15 11 11 13 10 9 0 13 1 11 11 2 13 1 12 2
13 1 10 9 2 13 1 10 9 0 1 10 9 2
13 10 9 1 10 9 1 10 9 4 13 1 11 2
8 10 0 9 1 9 15 13 2
36 1 10 9 7 10 9 2 10 9 4 13 10 9 1 9 0 2 7 3 2 1 10 9 2 15 4 13 10 3 0 9 1 13 10 9 2
41 10 0 11 11 11 15 4 13 1 10 12 1 10 12 9 12 1 10 9 2 1 9 0 2 9 0 2 2 11 11 2 11 11 2 11 11 2 11 11 2 2
21 12 2 10 11 13 10 9 1 10 9 1 10 11 7 1 10 9 1 10 9 2
13 10 9 1 9 13 3 1 9 0 1 11 11 2
7 10 9 13 0 1 11 2
37 15 4 13 10 9 0 1 10 9 0 7 10 9 0 7 0 3 1 13 10 9 1 3 1 3 0 2 1 10 9 1 10 2 9 0 2 2
27 1 10 0 9 1 10 9 2 10 9 13 1 9 13 2 11 11 2 7 15 13 1 13 1 10 11 2
20 10 9 13 10 11 7 15 13 1 11 1 11 2 9 1 9 1 10 9 2
10 9 1 10 9 0 2 1 9 0 2
35 10 11 11 7 10 11 11 2 13 11 11 1 10 9 0 2 4 13 2 1 10 9 11 11 2 1 10 9 11 9 1 13 1 12 2
14 15 4 3 13 10 9 1 10 9 15 15 4 13 2
5 10 9 13 0 2
31 3 0 1 10 9 2 10 9 15 13 1 10 9 0 13 7 1 10 0 9 0 9 1 10 9 1 10 9 11 11 2
23 11 11 11 13 15 1 10 9 1 10 9 1 9 0 11 13 1 11 11 7 11 11 2
12 10 9 13 7 15 13 3 9 1 10 9 2
17 13 1 11 2 15 13 12 0 9 1 10 9 7 10 9 0 2
12 10 9 13 10 9 1 11 7 10 11 0 2
22 10 9 0 0 1 10 9 15 13 3 1 10 12 5 9 7 10 9 12 5 9 2
25 15 15 13 1 11 11 1 10 3 0 9 0 1 10 9 7 12 9 1 9 11 11 1 11 2
30 15 13 10 0 9 1 9 13 1 12 1 12 9 7 10 9 13 2 1 10 9 15 15 13 12 9 1 10 13 2
10 10 9 1 9 4 13 1 10 9 2
7 11 14 13 3 1 9 2
7 13 0 2 0 7 0 2
24 15 13 1 10 11 1 10 9 12 7 13 10 9 1 10 11 11 11 1 11 2 11 11 2
17 3 2 15 13 15 1 10 0 9 1 10 9 2 15 1 3 2
40 10 9 1 10 9 0 7 1 10 9 2 1 10 9 0 2 4 13 10 0 9 1 10 9 15 2 1 10 9 1 10 9 12 2 4 13 10 9 0 2
10 15 13 1 9 12 1 10 11 11 2
39 15 4 13 1 12 1 13 10 9 1 10 9 1 10 9 1 10 9 1 12 2 7 15 14 4 13 3 1 10 11 12 2 1 9 1 9 1 9 2
20 11 13 1 13 10 9 1 11 1 10 9 15 13 1 10 9 1 10 9 2
25 11 11 14 13 3 2 15 13 1 10 10 9 1 10 9 2 15 13 1 10 9 9 7 9 2
24 10 9 11 11 4 4 13 9 1 9 1 10 9 0 15 13 1 9 10 9 1 11 12 2
50 11 13 1 10 0 9 15 4 13 10 11 4 13 1 10 9 0 7 2 3 1 10 9 2 15 4 13 10 9 1 10 12 1 11 11 15 10 9 1 9 13 9 7 13 12 9 1 10 11 2
20 15 15 13 1 10 9 2 3 1 10 9 13 3 1 10 9 1 10 9 2
42 10 9 13 10 9 1 10 9 13 2 1 10 9 1 10 9 2 11 11 2 11 11 2 11 2 11 2 11 11 2 11 2 11 11 2 11 2 11 7 11 11 2
38 3 1 10 9 2 0 11 2 7 11 2 4 13 1 11 1 13 10 9 2 3 1 4 13 1 12 1 10 0 9 15 13 10 9 1 10 9 2
4 15 4 13 2
22 3 2 1 11 11 2 10 9 11 12 14 4 3 4 13 2 7 14 15 13 3 2
36 10 9 0 13 9 1 12 1 12 7 15 15 13 3 1 10 9 0 15 15 13 12 9 1 9 2 12 9 1 9 7 12 9 1 9 2
24 11 13 10 9 1 10 9 0 1 9 1 11 1 10 11 2 13 1 10 9 0 1 11 2
33 2 11 13 16 10 9 13 0 1 15 1 10 9 0 2 2 1 15 2 11 7 11 2 1 3 16 11 2 13 15 3 11 2
16 10 9 13 16 12 9 4 4 13 1 10 9 1 10 9 2
38 15 14 4 3 13 1 13 1 10 9 12 2 10 9 13 1 13 10 9 0 1 10 11 9 1 10 9 0 1 10 9 0 1 10 9 0 2 2
12 1 10 9 0 2 10 9 13 1 10 9 2
13 1 10 9 1 15 13 10 9 7 13 10 9 2
22 1 0 9 1 10 9 1 10 9 15 13 10 0 9 1 10 9 7 10 9 13 2
40 12 0 9 0 2 10 9 11 2 11 2 11 7 10 9 11 13 10 9 1 13 10 9 1 9 0 1 10 0 9 0 2 1 1 10 9 0 13 9 2
19 15 13 9 1 10 9 0 1 10 0 9 0 2 13 11 2 1 12 2
36 10 9 13 1 12 9 1 10 9 0 15 13 1 10 0 9 0 0 7 13 10 9 1 10 11 3 1 4 13 1 10 9 1 10 11 2
37 10 9 1 11 4 3 13 1 10 11 2 15 13 3 10 9 0 1 9 13 1 10 9 0 2 10 9 2 10 9 7 10 0 9 1 9 2
22 1 3 2 10 0 9 13 1 10 9 4 13 9 1 10 9 1 10 9 1 11 2
16 10 0 9 15 10 9 13 13 10 9 1 9 1 10 9 2
41 3 1 10 9 0 1 10 9 1 10 9 1 10 9 2 11 13 3 2 3 2 1 13 10 9 0 1 10 9 0 1 9 1 10 9 0 2 0 7 0 2
18 15 13 1 10 9 0 1 10 9 1 11 11 16 15 13 1 12 2
24 1 12 2 15 13 10 9 1 10 9 1 11 1 15 13 1 12 9 1 12 9 1 9 2
21 11 2 11 2 11 2 12 2 13 10 9 0 0 1 10 9 1 10 12 9 2
34 13 1 11 11 2 10 9 1 10 11 13 3 10 11 1 11 2 3 0 9 0 2 7 10 11 1 11 2 0 9 1 10 11 2
15 15 15 13 10 9 1 3 1 12 9 1 9 1 9 2
15 0 9 7 10 9 1 9 1 10 9 4 13 3 0 2
37 14 15 13 3 10 9 2 15 15 9 1 11 11 15 2 1 9 2 13 1 13 11 7 11 1 16 11 11 15 13 1 10 9 1 10 9 2
22 11 2 13 15 1 10 9 1 9 1 10 9 0 2 11 2 1 10 11 11 0 2
17 15 13 1 0 9 15 15 13 1 10 9 15 10 9 0 13 2
30 10 9 2 1 2 12 9 1 9 2 2 1 10 9 2 7 1 2 15 1 9 2 2 13 3 1 9 1 12 2
30 15 13 1 11 1 12 1 10 11 11 15 15 13 1 10 9 12 7 12 16 12 9 2 15 12 1 12 9 2 2
28 1 13 10 9 1 10 9 1 9 2 15 13 10 11 1 11 2 15 13 1 12 5 7 12 5 1 9 2
98 11 11 2 13 10 12 9 12 1 10 9 1 11 2 1 11 2 3 1 11 2 13 10 12 9 12 2 1 10 9 1 11 2 9 1 11 11 2 12 1 11 2 12 2 11 2 13 10 9 0 2 13 1 10 9 1 4 2 1 10 11 11 0 2 13 3 1 9 0 1 10 11 0 13 1 9 1 10 9 1 10 2 11 0 2 2 1 15 15 13 0 2 2 10 9 11 11 2
53 10 9 15 4 3 13 1 15 15 15 13 3 1 10 9 2 1 10 9 7 10 9 0 13 10 9 0 1 10 9 7 1 10 9 0 1 10 0 9 7 9 0 15 4 13 10 11 0 1 10 11 11 2
48 10 9 0 1 10 9 2 10 3 0 9 1 10 11 11 11 2 4 13 10 9 1 10 9 0 2 9 0 13 1 10 9 9 2 2 15 15 13 1 0 2 9 2 1 10 9 0 2
27 15 14 13 3 15 2 10 9 0 2 1 10 9 2 15 14 13 3 1 10 9 0 7 14 15 13 2
44 10 9 15 13 1 13 1 10 9 1 11 11 2 0 9 1 9 1 10 11 7 9 0 1 10 9 1 11 13 1 10 9 1 11 1 10 11 0 1 10 9 1 11 2
41 10 0 9 0 2 0 2 0 2 7 15 13 10 3 13 1 11 2 4 13 1 15 13 10 9 0 1 10 9 1 10 9 15 15 4 13 1 10 9 0 2
11 11 13 10 9 1 10 9 0 1 11 2
13 12 9 4 13 1 10 9 7 12 1 10 9 2
6 15 13 3 10 9 2
14 1 12 1 12 9 2 10 9 4 13 10 9 0 2
42 9 1 10 9 4 13 1 10 9 1 10 9 1 10 9 1 10 11 2 1 9 10 9 1 10 9 11 10 11 6 13 10 9 1 10 11 1 10 9 1 11 2
6 10 9 4 3 13 2
19 11 13 10 9 1 10 9 1 11 1 10 11 1 10 11 1 10 11 2
12 11 11 13 10 0 9 0 0 13 1 12 2
13 11 11 13 12 9 1 10 11 7 1 10 11 2
27 13 1 10 0 9 1 10 9 1 10 9 7 10 9 2 1 16 15 13 10 0 9 1 10 0 9 2
65 10 9 11 1 10 11 13 10 9 1 10 9 2 10 9 7 10 9 0 2 0 1 10 9 1 9 11 2 2 1 13 1 10 9 2 1 10 9 1 10 9 2 1 13 10 9 0 1 10 9 1 10 9 0 7 1 13 9 1 10 9 3 0 2 2
28 3 16 15 15 13 1 9 2 15 13 0 1 13 16 10 9 1 10 9 14 15 13 3 1 10 9 1 9
16 10 9 13 10 9 13 10 9 7 13 10 9 1 11 11 2
17 10 9 2 12 5 2 13 0 1 10 9 0 2 12 5 2 2
20 1 9 2 15 4 13 1 11 7 13 1 10 9 1 11 2 3 1 11 2
19 15 14 15 13 3 10 9 2 10 9 4 13 1 12 9 10 9 0 2
26 10 9 0 13 10 0 9 0 2 3 16 10 11 13 2 0 2 2 1 9 3 1 1 9 2 2
26 1 10 9 2 15 4 13 3 1 13 13 10 9 0 1 9 0 16 11 2 11 11 2 7 11 2
13 10 9 0 11 15 4 13 10 9 1 12 9 2
12 9 11 4 1 3 13 13 15 1 10 9 2
25 10 9 4 13 1 10 9 1 9 2 3 11 2 11 7 11 11 11 2 9 0 1 10 9 2
42 13 1 11 1 1 10 11 2 11 13 2 1 9 7 1 9 2 10 9 1 10 9 0 7 0 2 10 9 0 7 10 9 2 7 10 9 1 9 1 10 9 2
12 15 4 3 13 1 10 9 1 11 1 11 2
30 15 13 16 9 1 10 9 0 2 15 13 9 16 10 9 15 13 1 13 1 15 15 15 13 2 10 9 0 2 2
32 10 9 13 10 9 13 1 10 0 9 13 3 1 9 7 13 1 10 0 9 1 10 11 11 2 10 9 1 9 1 11 2
26 10 9 1 9 13 1 10 9 1 10 0 11 1 11 13 1 9 1 9 10 9 1 9 11 11 2
45 10 12 9 15 4 3 3 13 3 1 9 3 0 2 10 12 9 12 2 12 1 10 2 11 11 1 11 2 2 3 10 12 9 12 2 10 12 9 12 7 10 12 9 12 2
20 3 1 15 1 11 11 2 15 1 11 13 10 9 4 13 10 9 1 11 2
23 15 4 13 10 9 1 9 1 9 1 10 9 0 1 10 11 11 15 15 13 10 9 2
16 1 12 2 15 4 13 9 1 10 9 11 11 1 10 11 2
12 10 9 1 10 12 0 9 13 10 0 9 2
15 10 9 14 15 13 3 12 9 3 3 1 10 9 11 2
17 10 10 9 11 2 0 9 2 4 13 3 16 12 1 10 9 2
38 10 9 13 10 9 1 10 9 10 9 1 10 9 2 7 15 4 13 10 9 0 2 1 10 9 7 10 9 2 1 9 1 10 9 1 10 9 2
21 10 9 0 2 15 4 13 1 10 11 1 10 9 1 10 11 1 3 16 9 2
16 11 13 10 9 0 2 3 0 7 0 1 15 1 13 0 2
23 3 1 3 2 10 10 9 1 10 9 1 10 11 4 13 2 3 13 10 0 9 9 2
26 10 0 9 1 10 11 2 0 9 1 10 9 1 11 2 13 10 15 1 10 3 0 1 10 11 2
31 10 9 13 3 9 1 10 9 7 10 9 0 14 4 13 3 1 10 9 2 4 13 1 10 9 0 15 13 10 9 2
9 9 11 15 13 11 11 1 9 2
20 10 9 4 1 0 13 7 10 9 13 16 11 4 13 11 16 15 15 13 2
25 11 15 13 1 4 13 10 15 1 10 12 9 1 10 2 9 12 2 2 15 13 10 11 0 2
17 1 12 2 15 13 10 9 1 10 0 9 1 10 9 1 9 2
26 15 13 10 9 1 10 9 1 10 9 11 11 2 15 13 10 9 13 1 11 11 2 3 1 11 2
17 10 9 15 13 3 1 10 9 1 10 11 1 13 10 9 0 2
27 15 4 3 13 1 13 10 9 1 9 1 10 9 1 9 1 10 11 11 7 1 10 9 0 1 11 2
13 10 9 0 2 11 11 2 13 10 0 9 0 2
31 1 13 10 9 3 0 2 15 13 9 1 10 9 0 2 1 9 2 9 2 15 13 1 10 9 0 1 9 10 9 2
37 9 11 4 13 16 10 11 4 13 1 13 10 9 1 10 11 0 1 9 1 11 7 10 9 0 1 11 2 1 16 10 9 0 4 13 2 2
11 10 9 15 13 0 1 13 1 10 9 2
11 3 13 15 2 15 14 13 3 10 9 2
27 11 13 10 9 2 7 14 13 3 10 9 2 9 1 10 9 1 10 9 1 10 9 1 10 9 12 2
7 9 1 10 9 3 0 2
33 3 2 10 9 13 0 1 10 9 1 10 9 0 13 1 10 9 2 9 7 9 2 13 1 0 9 1 10 9 1 10 9 2
15 15 13 1 15 4 13 10 9 1 10 9 1 16 0 2
51 1 14 13 3 3 10 9 1 9 1 10 11 1 9 1 10 11 0 2 10 11 7 10 11 14 15 4 3 2 1 9 2 13 1 10 9 0 1 10 9 1 10 11 1 10 9 1 10 9 0 2
18 16 15 13 2 3 10 9 2 11 13 3 1 15 13 10 0 9 2
30 10 11 13 10 9 1 0 9 1 1 10 9 1 11 2 3 16 15 15 3 13 1 15 10 9 1 10 9 11 2
13 15 13 10 9 1 15 10 9 13 1 9 0 2
32 10 9 11 15 13 1 0 9 1 10 9 0 1 10 9 1 1 15 16 10 9 1 10 9 14 15 13 1 13 10 9 2
13 15 4 13 1 0 9 1 10 9 1 10 9 2
4 9 7 9 2
12 7 2 10 9 1 11 13 0 1 10 9 2
27 11 13 3 1 13 10 9 1 10 9 1 10 9 2 7 3 15 13 1 4 13 7 13 13 10 9 2
18 10 9 7 13 2 11 2 13 1 9 10 9 1 9 1 10 9 2
16 10 11 2 1 10 9 1 10 0 9 2 13 10 9 0 2
21 10 12 9 12 2 11 11 13 10 9 1 11 11 7 11 11 1 10 9 11 2
58 2 15 13 10 9 1 10 11 1 10 9 1 10 9 1 10 9 2 3 1 10 11 16 1 10 9 1 10 11 7 3 7 15 15 13 3 0 2 2 4 13 11 11 1 10 9 1 9 13 1 10 9 1 10 11 1 11 2
12 15 4 3 13 1 12 9 2 1 12 9 2
18 1 10 9 1 10 9 15 13 10 9 11 1 9 2 0 7 0 2
16 3 1 11 11 2 15 13 10 9 1 10 9 1 10 9 2
59 11 11 2 13 10 12 9 12 1 11 7 13 1 9 12 1 11 2 13 10 9 0 2 9 1 9 1 10 11 1 11 1 12 1 12 2 9 1 10 9 1 10 9 1 12 1 12 2 9 13 1 10 11 1 10 11 1 12 2
13 10 9 1 10 9 15 13 1 10 9 1 9 2
26 1 10 9 10 9 0 4 13 1 9 1 10 9 3 3 13 7 1 10 9 15 15 4 4 13 2
15 15 13 10 9 1 12 9 7 13 10 9 1 12 9 2
17 1 10 9 1 10 0 9 2 10 11 15 13 1 11 9 9 2
62 1 10 0 9 2 15 13 1 10 9 1 11 2 15 13 1 10 9 10 9 1 9 1 9 1 10 0 9 1 10 9 1 9 2 1 15 3 13 1 13 15 15 15 13 10 2 9 2 2 1 4 13 2 2 7 13 2 10 0 9 13 2
9 10 0 9 4 13 10 9 1 12
20 13 1 10 9 0 11 12 2 15 13 10 0 9 0 1 13 10 9 0 2
31 1 12 2 1 11 2 11 11 11 13 7 13 10 10 9 9 9 1 10 9 13 1 10 9 2 10 9 11 11 11 2
18 10 9 1 10 9 13 1 10 9 12 7 15 13 1 10 9 12 2
37 10 9 0 13 1 0 9 1 10 9 2 3 16 15 13 3 1 9 2 1 3 1 11 2 15 4 13 1 12 9 2 3 13 1 11 2 2
14 10 9 13 10 9 1 9 2 9 2 9 2 9 2
13 10 9 13 1 3 12 9 1 9 7 1 9 2
20 10 9 1 9 15 13 1 15 13 1 11 11 15 15 13 1 1 10 9 2
9 15 13 16 11 11 12 4 13 2
17 10 11 0 7 10 11 4 13 1 10 11 11 1 10 11 0 2
34 10 0 9 4 4 13 1 10 11 1 12 1 10 9 15 4 13 1 12 1 10 9 15 15 13 1 15 13 1 10 9 1 11 2
19 1 12 2 15 4 13 9 1 10 11 2 9 15 15 13 1 1 12 2
21 10 9 11 11 13 3 9 1 10 9 1 10 9 3 1 15 13 1 0 9 2
13 15 13 12 9 3 0 16 10 9 14 13 3 2
20 15 4 13 1 9 1 13 10 9 1 9 0 1 13 1 10 9 1 9 2
20 10 0 9 1 11 2 11 7 11 13 3 10 9 1 10 9 1 10 11 2
22 10 9 15 4 13 10 9 7 10 9 1 9 4 13 1 9 1 1 10 9 12 2
17 10 9 1 10 9 4 13 1 10 9 7 10 9 1 10 9 2
21 10 9 1 11 1 9 1 12 12 13 10 9 1 10 9 1 10 9 1 12 2
21 15 4 3 13 1 10 9 1 10 9 11 2 11 2 2 15 13 11 1 11 2
19 10 12 9 12 2 15 13 1 10 0 9 9 1 11 11 1 11 11 2
19 10 9 13 1 13 16 15 14 13 3 10 9 3 1 13 10 9 0 2
29 1 9 11 2 10 9 1 9 11 4 2 3 13 1 10 9 0 2 2 16 15 13 10 9 0 1 10 9 2
34 3 15 13 1 10 9 0 1 10 9 0 1 10 9 0 0 16 4 13 10 0 9 1 9 1 11 11 1 10 9 1 9 0 2
17 11 11 11 11 11 4 13 10 0 9 12 1 11 2 11 2 2
31 1 10 9 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2
29 10 9 4 13 2 3 1 15 2 1 2 0 2 7 15 13 0 1 9 0 1 10 9 0 16 1 10 9 2
25 10 9 4 3 13 1 10 9 0 2 0 2 0 7 0 2 3 1 13 10 9 2 9 2 2
30 3 2 1 10 9 2 10 9 0 2 10 9 2 7 10 9 0 0 16 11 13 1 10 9 1 9 10 9 0 2
12 10 9 10 3 0 4 13 12 1 12 9 2
42 10 0 9 2 1 10 9 1 10 11 0 2 1 10 0 9 1 10 9 11 1 10 11 1 10 9 2 12 2 13 3 16 15 4 3 13 10 9 7 10 9 2
14 10 9 1 10 9 4 13 1 15 13 1 10 9 2
33 1 9 2 3 10 9 0 13 0 2 3 15 4 15 13 10 9 0 1 15 13 2 1 9 0 2 1 10 9 1 10 9 2
21 11 11 13 10 9 0 13 1 12 1 11 11 1 1 10 9 0 1 11 11 2
16 15 4 4 13 10 0 9 1 10 9 11 10 12 9 12 2
51 10 9 0 15 4 13 1 9 2 8 5 12 2 1 10 12 9 12 2 1 10 9 0 0 1 10 11 1 10 9 15 15 4 4 13 1 10 12 9 1 9 1 10 9 12 7 12 1 10 9 2
32 1 9 1 11 11 1 10 9 12 2 15 13 13 1 10 9 7 10 9 1 9 1 10 9 1 9 0 1 10 9 0 2
39 10 9 0 13 10 0 9 3 1 10 9 1 12 1 10 9 1 11 1 10 9 11 12 1 11 2 15 13 3 10 9 0 7 13 1 10 9 0 2
35 10 9 13 3 3 10 0 9 2 11 2 11 2 11 2 2 15 14 13 3 10 9 3 1 10 9 2 7 1 10 9 1 10 9 2
18 10 11 11 11 11 11 13 10 9 1 9 13 1 11 1 11 11 2
16 13 1 11 2 11 2 2 1 11 2 11 13 10 9 11 2
10 15 13 10 9 1 11 7 1 11 2
21 10 9 1 10 9 1 11 13 1 10 9 1 10 9 2 7 1 10 9 2 2
34 10 9 4 13 1 9 13 1 10 9 7 1 9 0 0 16 10 9 2 10 9 0 2 10 9 1 9 7 10 9 1 10 9 2
34 1 3 2 10 9 13 3 0 7 10 9 13 1 10 9 1 9 13 1 9 13 1 10 9 1 9 1 10 11 7 1 10 11 2
36 10 9 4 13 1 12 7 12 1 10 9 0 11 10 11 2 1 9 1 10 9 2 1 10 9 0 2 9 1 10 9 7 1 10 9 2
11 10 9 0 14 4 13 1 9 0 11 2
23 10 9 0 2 1 9 0 2 15 13 1 10 9 0 7 3 3 1 10 9 1 9 2
10 15 13 10 9 1 9 0 1 11 2
19 15 15 13 3 1 10 9 1 9 1 10 9 7 10 10 9 1 9 2
23 11 13 10 15 1 10 12 9 1 10 9 1 9 0 0 1 10 9 1 10 11 11 2
18 1 10 9 1 9 0 11 11 11 2 10 9 13 3 0 1 11 2
49 1 9 2 1 9 0 2 10 9 1 9 13 3 10 9 1 9 0 2 10 9 0 14 13 10 9 8 5 5 13 3 1 10 9 1 10 9 0 3 1 10 9 1 10 9 1 9 2 2
13 11 11 13 10 9 13 1 10 9 1 10 11 2
19 3 1 12 9 15 13 1 10 9 1 10 9 1 10 9 1 10 9 2
22 3 2 1 9 12 2 11 11 2 9 1 10 9 11 2 9 1 11 7 10 9 2
35 10 9 0 1 10 9 2 10 9 1 10 9 1 9 2 10 0 9 6 13 10 9 0 2 13 1 13 16 10 0 9 13 10 9 2
9 10 9 4 3 13 10 0 9 2
7 15 4 13 1 11 11 2
23 11 13 10 0 9 1 10 9 2 7 10 9 1 10 9 2 9 1 10 9 1 9 2
13 1 10 9 0 2 15 13 10 9 0 1 9 2
31 15 1 10 9 14 4 4 13 1 11 7 10 9 1 9 13 15 1 10 9 1 11 11 1 11 7 11 11 11 11 2
15 10 0 9 15 13 13 1 13 1 10 9 1 11 11 2
15 3 10 9 1 11 15 13 1 0 9 1 10 9 13 2
19 3 13 1 10 9 2 13 10 9 1 9 7 1 9 13 1 10 9 2
17 10 0 9 13 3 1 13 10 9 1 9 0 7 1 10 9 2
25 15 13 11 7 15 13 1 10 9 0 1 11 3 16 15 13 10 9 7 10 9 1 10 9 2
25 10 9 1 10 9 13 13 10 8 8 15 15 13 10 9 0 2 0 7 0 1 10 11 0 2
35 10 12 11 11 4 13 9 1 11 2 1 9 0 3 2 15 10 9 9 4 13 1 11 2 15 13 3 10 2 9 1 10 9 2 2
22 10 11 11 15 4 13 1 10 9 1 9 1 10 9 0 1 10 11 7 10 11 2
23 10 9 11 4 13 10 9 1 9 1 9 3 16 11 4 4 13 1 10 9 1 12 2
25 10 0 9 1 10 0 9 13 16 15 4 3 13 10 9 1 10 9 13 16 13 1 10 9 2
22 10 11 0 13 3 10 9 1 10 9 0 1 9 1 10 9 0 13 1 12 9 2
21 2 15 15 4 13 3 15 15 13 10 9 2 7 15 9 15 3 1 10 9 2
14 1 12 1 12 2 10 9 13 3 10 9 2 9 2
10 10 15 1 10 0 9 1 12 5 2
12 10 9 13 1 10 3 10 9 1 10 9 2
24 11 11 11 2 9 2 11 11 11 2 2 13 10 12 9 12 1 11 2 13 10 9 0 2
33 11 2 1 11 13 10 9 0 2 9 0 2 13 1 9 1 11 2 1 11 11 1 12 1 11 11 2 11 11 7 11 11 2
14 10 0 9 4 4 13 1 11 2 1 11 1 11 2
16 1 9 2 15 13 10 9 0 2 15 13 3 10 0 9 2
14 15 14 13 3 0 2 10 9 13 10 9 1 11 2
11 10 0 9 13 1 10 9 13 1 12 2
19 1 9 2 10 9 14 13 3 1 10 9 16 15 15 13 1 10 9 2
12 10 0 9 1 10 9 1 11 13 1 12 2
11 1 10 9 1 12 2 15 13 12 9 2
24 10 9 1 10 9 4 13 3 16 10 15 4 13 1 10 9 0 2 13 1 10 0 9 2
55 10 9 0 2 1 10 11 11 11 2 13 10 9 13 1 10 9 1 10 11 2 10 9 13 2 1 10 11 3 1 10 11 11 2 10 9 15 4 13 1 10 9 0 2 1 13 10 9 1 10 9 1 10 11 2
21 1 10 9 13 1 10 9 1 11 2 1 10 9 1 11 2 4 13 12 9 2
16 10 9 13 1 3 10 9 3 0 1 10 9 1 10 11 2
39 15 4 13 1 12 1 13 10 9 1 10 9 1 10 9 1 10 9 1 12 2 7 15 14 4 13 3 1 10 11 12 2 1 9 1 9 1 9 2
24 3 3 10 9 1 10 9 16 1 10 0 9 11 2 11 7 11 4 13 10 9 1 11 2
20 10 9 13 10 0 9 2 7 10 9 14 13 3 3 0 1 15 1 3 2
19 10 9 4 13 1 10 9 1 10 9 0 1 9 1 10 12 9 12 2
38 10 2 9 2 15 15 13 3 1 9 13 10 9 0 1 10 9 1 9 1 9 1 10 9 0 7 0 15 15 13 1 11 1 10 11 1 12 2
18 11 13 1 10 9 1 9 1 10 9 1 9 1 11 2 10 9 2
47 13 10 9 0 15 13 10 9 2 11 11 13 9 1 10 0 9 1 10 9 2 13 1 13 1 10 0 9 0 13 1 10 9 0 7 0 0 15 13 3 10 9 0 1 10 9 2
6 11 7 11 4 13 2
15 1 10 9 1 10 9 2 15 13 15 14 13 3 0 2
6 10 9 4 3 13 2
29 13 1 10 9 10 12 9 12 2 10 9 4 13 1 10 9 1 10 12 12 2 12 9 7 1 10 9 0 2
36 11 2 9 1 10 9 1 10 9 2 11 2 11 11 2 13 10 9 1 9 13 1 11 11 2 9 13 1 10 9 1 9 0 0 11 2
29 10 9 13 3 0 2 10 9 4 13 1 9 0 1 3 1 9 3 13 1 10 0 9 1 10 9 1 9 2
14 15 4 3 13 1 0 9 7 9 2 3 15 13 2
42 1 12 2 10 11 13 10 9 1 9 3 1 10 9 0 1 11 2 3 16 1 10 11 1 10 9 1 11 2 15 13 1 10 11 11 11 7 10 11 11 11 2
26 11 13 10 0 9 1 10 11 0 0 1 10 11 15 4 2 3 2 13 10 9 10 12 9 12 2
16 15 15 13 1 10 11 11 11 2 1 11 7 3 1 11 2
47 1 10 11 2 10 12 1 12 1 9 4 13 11 1 13 10 9 1 10 9 11 11 11 2 15 15 15 4 13 1 10 9 0 11 11 7 4 13 11 7 10 11 1 13 10 9 2
10 10 9 1 9 0 7 0 13 3 2
8 10 9 4 13 1 10 11 2
20 2 2 11 13 1 10 9 1 13 9 1 10 11 2 2 3 0 16 3 2
19 15 4 3 13 16 10 9 13 3 10 9 1 13 10 0 9 1 11 2
28 1 3 2 16 15 13 16 10 9 1 10 9 13 10 0 9 2 15 13 16 10 9 13 3 1 0 9 2
16 10 9 13 10 9 1 12 9 7 1 16 15 13 10 9 2
18 1 12 2 11 13 2 16 10 9 1 12 5 1 9 1 12 2 2
18 13 1 10 9 1 10 9 7 10 9 0 2 11 13 1 13 11 2
36 10 9 0 1 10 11 2 15 15 13 1 10 9 0 2 11 2 4 3 13 10 9 0 1 2 13 3 10 10 9 1 10 9 0 2 2
12 9 11 13 10 9 13 1 11 2 1 11 2
40 1 13 1 15 2 10 11 13 1 9 10 9 1 10 0 9 1 9 1 9 0 2 13 12 9 1 10 9 1 10 9 2 15 10 0 9 13 10 9 2
8 10 9 13 10 9 1 9 2
24 10 9 0 7 0 1 10 9 13 10 9 16 15 14 13 3 13 1 10 9 1 10 9 2
20 10 12 11 1 10 9 0 4 13 1 10 9 1 10 9 1 10 12 9 2
41 10 9 13 3 3 0 1 1 12 9 1 10 9 13 1 10 9 0 7 1 10 9 2 15 13 12 5 1 10 9 1 10 0 9 3 12 5 1 10 9 2
33 15 13 3 10 9 2 11 8 11 11 2 15 13 10 0 9 7 2 11 11 2 15 13 9 1 10 9 0 1 10 9 11 2
22 12 2 10 9 1 10 9 1 9 2 11 2 15 13 3 0 1 10 9 1 11 2
23 1 10 9 1 9 7 10 9 1 9 2 10 9 7 10 9 1 10 9 15 13 3 2
38 16 10 9 1 10 10 9 1 11 13 10 9 0 1 10 9 0 7 0 2 10 9 4 3 3 13 2 1 1 12 5 1 3 1 9 12 2 2
19 11 11 2 13 10 12 9 12 1 11 2 13 10 0 9 0 1 9 2
22 11 11 14 4 3 4 13 1 10 9 1 10 9 7 14 4 1 9 3 13 3 2
21 1 13 10 9 1 10 10 0 11 2 11 4 13 9 1 9 0 1 10 9 2
7 10 9 0 15 13 15 2
38 10 0 9 13 10 9 1 10 9 15 13 10 0 7 0 9 2 16 15 14 13 16 15 4 4 13 0 2 9 2 9 2 1 9 1 10 9 2
24 10 9 1 11 13 10 9 1 10 12 9 1 10 11 1 11 13 1 10 11 0 1 11 2
13 11 1 11 13 10 9 1 11 1 12 1 12 2
26 10 9 1 10 9 13 1 10 9 1 10 9 3 16 10 9 1 9 2 11 11 13 1 11 11 2
50 10 11 2 1 10 9 0 2 0 2 9 2 9 2 13 10 9 1 10 9 1 10 9 15 13 10 9 0 0 13 1 10 9 0 7 2 10 3 3 2 1 12 9 2 10 9 7 10 9 2
32 10 9 0 13 1 13 10 9 1 10 9 2 10 9 3 0 15 13 2 10 9 1 10 9 3 2 3 10 9 15 13 2
54 1 12 2 10 9 15 13 1 11 7 13 3 1 10 9 1 10 9 11 1 11 10 9 4 13 3 3 2 11 13 3 1 13 10 9 7 10 9 1 9 2 7 13 1 9 11 12 7 10 9 11 1 11 2
20 15 13 3 12 1 4 13 10 9 1 10 9 1 9 2 3 1 10 9 2
49 7 3 1 10 9 1 10 9 0 1 9 1 9 2 15 13 10 9 16 3 1 9 7 16 1 9 0 2 15 15 1 10 9 4 13 1 10 9 1 10 9 16 1 9 15 13 1 9 2
17 10 9 13 10 9 0 13 1 12 7 12 1 11 11 1 11 2
21 1 4 15 13 0 2 15 14 4 3 15 13 16 15 13 10 9 15 13 2 2
38 10 9 1 11 13 10 9 0 0 13 1 10 9 1 10 11 2 1 9 0 1 10 9 10 11 0 2 1 10 9 1 10 11 7 10 9 11 2
53 2 10 9 1 10 9 1 10 9 13 3 3 0 7 0 1 10 9 0 15 1 10 9 0 1 10 9 1 10 9 0 4 13 7 13 1 13 10 9 1 0 9 2 2 4 13 10 9 1 13 10 9 2
34 3 10 15 1 10 0 9 13 1 9 0 1 11 2 15 13 10 9 0 2 12 9 0 7 12 0 9 1 10 9 1 10 9 2
15 15 13 16 10 9 1 9 13 0 1 10 3 1 9 2
19 15 13 10 9 11 15 15 13 1 13 1 11 2 1 11 7 1 11 2
26 0 1 11 11 11 2 10 9 13 1 10 9 0 1 10 9 7 10 9 0 2 1 10 9 0 2
25 10 11 4 3 13 10 11 1 10 9 0 7 1 9 1 10 9 15 13 0 1 10 9 0 2
41 10 9 1 10 9 0 1 10 9 2 10 9 0 2 10 9 1 10 9 1 9 1 9 7 10 9 1 10 9 13 3 1 9 15 4 13 10 9 1 9 2
58 15 13 1 10 0 9 16 13 10 9 1 9 13 1 0 9 4 13 10 9 1 9 0 1 10 9 2 9 0 2 7 13 3 10 9 1 9 13 1 10 9 0 2 3 16 10 9 7 10 9 3 0 4 3 15 13 9 2
19 3 12 9 4 4 13 1 13 16 0 10 9 1 10 9 1 10 9 2
22 3 1 13 3 10 11 0 2 10 11 1 11 1 12 13 10 9 1 10 0 11 2
28 9 0 1 9 13 1 10 9 1 11 2 10 9 4 13 3 1 9 1 10 9 1 9 9 1 10 9 2
39 1 3 2 10 9 2 1 10 9 13 2 4 4 13 3 1 14 3 13 10 9 6 13 10 9 1 10 9 2 3 10 9 1 10 9 1 10 9 2
18 1 12 15 4 13 10 9 0 2 1 9 1 10 9 1 0 9 2
6 15 4 13 1 13 2
13 6 2 15 13 3 10 9 3 0 7 3 0 2
32 10 9 4 3 13 1 10 11 3 1 10 9 1 10 9 2 1 10 9 2 15 11 13 10 0 7 0 9 1 10 9 2
27 11 11 2 13 10 12 9 12 1 10 11 7 13 10 12 9 12 1 11 2 13 10 9 1 9 0 2
25 10 9 1 12 9 4 13 1 10 9 0 1 1 10 9 1 12 1 12 9 1 3 12 9 2
46 10 9 6 13 10 9 13 10 9 0 1 10 0 9 15 2 1 9 1 10 9 0 3 13 1 10 9 2 14 4 4 13 3 1 10 9 1 9 2 12 9 1 9 0 2 2
19 11 7 11 11 15 13 13 10 9 1 11 2 10 9 7 10 9 0 2
33 3 16 11 13 1 10 9 2 11 15 13 7 10 9 13 1 13 10 9 11 7 10 9 15 13 3 2 15 13 1 10 9 2
38 10 11 13 3 10 9 0 1 10 9 1 10 9 2 7 13 1 10 9 1 10 9 7 13 10 9 1 10 9 13 1 9 1 9 7 1 9 2
8 3 13 10 9 1 10 9 2
10 9 7 9 1 10 12 9 1 13 2
25 10 9 14 15 13 3 0 7 15 13 10 9 0 1 10 9 1 11 2 11 2 11 7 11 2
8 15 13 10 9 1 13 3 2
24 10 9 0 4 13 1 10 9 1 10 9 1 9 0 7 1 10 9 0 1 0 9 0 2
25 10 9 11 11 11 4 13 1 10 9 7 10 9 1 10 9 1 10 9 7 1 10 9 0 2
12 10 9 7 9 0 11 11 15 13 1 12 2
4 11 15 13 2
16 11 4 13 1 10 9 7 15 13 1 9 1 10 11 11 2
28 10 9 1 10 9 7 10 9 1 10 9 15 3 4 13 1 9 0 3 4 3 13 10 9 1 10 9 2
35 1 9 2 1 10 9 3 1 10 9 1 10 9 2 10 11 1 10 11 1 9 1 11 2 11 11 2 13 11 11 1 11 1 12 2
24 15 15 13 0 1 10 11 1 11 1 11 15 10 9 11 11 15 13 1 13 10 9 0 2
21 11 15 15 11 7 13 1 15 13 2 1 10 9 1 11 2 1 10 0 9 2
15 10 11 4 13 1 10 9 1 10 11 1 13 1 12 2
8 10 9 4 13 1 11 11 2
21 10 9 4 3 13 1 10 9 2 11 11 2 16 10 9 4 13 1 10 9 2
83 3 1 10 11 1 11 2 15 15 13 1 12 1 10 9 1 10 9 1 10 11 16 3 1 10 11 1 11 2 1 12 7 12 2 10 9 1 11 7 10 9 13 1 9 1 10 9 13 1 10 9 1 9 2 1 10 9 15 13 3 1 12 9 1 10 9 0 2 7 13 1 9 1 13 10 9 1 10 11 1 10 11 2
34 9 13 3 1 10 9 1 10 9 2 15 13 3 10 9 1 10 9 1 10 0 9 15 13 0 1 9 0 7 2 7 1 9 2
9 15 13 16 10 9 13 3 0 2
31 0 9 2 15 15 13 1 9 3 16 15 4 13 16 10 9 0 1 10 9 13 1 13 10 9 1 10 9 1 9 2
18 10 9 13 3 10 3 3 0 1 10 9 16 15 1 10 0 9 2
33 10 9 0 2 12 0 9 2 11 11 2 11 11 7 11 11 2 1 12 9 0 7 10 9 4 4 13 9 1 10 0 9 2
40 3 2 1 4 13 10 9 1 10 9 0 2 10 9 1 10 11 13 1 13 10 9 7 13 11 11 11 2 3 9 1 11 2 1 10 9 1 10 9 2
22 15 13 3 10 9 6 13 10 9 1 9 1 10 11 11 2 10 9 1 12 9 2
24 1 12 2 11 11 13 10 11 1 11 2 12 2 1 10 9 1 10 12 0 9 0 13 2
16 1 11 4 13 10 0 9 1 11 1 9 1 11 7 11 2
51 1 16 15 4 13 1 9 0 0 2 15 15 13 3 1 10 9 0 1 10 9 1 10 11 1 10 11 0 7 1 10 11 15 10 9 4 13 1 10 9 8 12 7 0 1 10 9 1 10 9 2
7 13 1 10 11 2 6 2
40 11 4 4 13 10 9 1 10 9 2 16 16 15 13 0 1 13 12 9 2 7 1 15 14 4 3 13 10 9 2 11 11 13 0 1 10 9 1 11 2
26 11 11 13 10 9 0 0 1 12 9 1 12 9 13 1 11 11 7 13 1 12 1 10 9 9 2
23 9 1 10 9 15 13 3 3 16 10 9 15 13 3 1 10 9 1 10 9 11 11 2
25 15 4 13 11 11 1 12 9 7 12 9 1 11 2 11 16 11 1 1 10 9 11 1 12 2
34 15 14 13 3 1 0 10 9 0 10 9 2 1 10 0 9 13 16 11 11 2 3 0 7 15 14 4 13 10 9 16 9 0 2
30 15 13 1 9 1 10 9 1 13 1 3 13 1 10 9 1 10 9 1 10 9 11 11 2 9 12 9 12 2 2
8 10 9 11 13 10 9 0 2
11 15 13 3 1 3 16 9 0 7 0 2
10 10 3 0 9 1 9 0 1 11 2
6 10 9 4 13 6 2
25 10 9 12 1 10 9 0 1 11 11 13 10 9 1 10 9 1 9 4 13 1 1 12 9 2
22 10 9 1 0 9 13 1 10 9 13 1 10 9 0 1 10 9 2 1 0 9 2
31 15 13 10 9 1 9 1 10 9 7 9 1 10 9 2 15 10 11 13 1 9 2 0 2 7 10 9 1 9 0 2
33 15 13 3 11 11 2 11 2 11 11 2 7 11 11 2 11 2 11 11 2 15 13 10 12 10 9 1 9 1 10 11 11 2
11 13 1 11 2 11 11 13 1 15 13 2
24 1 9 12 2 11 11 4 13 0 1 10 11 0 1 10 9 2 9 7 9 2 11 2 2
17 11 13 3 1 11 1 13 10 9 0 2 7 13 3 10 9 2
30 15 4 13 1 10 0 9 0 1 10 11 7 11 11 1 10 9 0 1 10 9 0 13 1 10 9 11 1 11 2
14 15 13 10 9 1 10 9 0 13 1 10 9 11 2
19 3 2 11 4 3 13 1 16 15 13 0 2 15 13 3 0 7 0 2
6 10 10 9 4 13 2
19 15 4 13 10 9 1 9 1 13 1 12 2 3 1 13 1 3 13 2
9 15 13 3 13 10 9 1 9 2
26 1 15 13 2 10 9 0 3 1 10 11 2 4 13 7 13 10 9 1 10 11 1 13 10 9 2
35 1 9 1 10 0 9 2 15 13 2 1 11 11 2 10 9 0 2 10 11 11 2 15 13 3 10 9 11 2 11 11 7 11 11 2
15 10 9 15 13 1 13 7 1 13 1 1 13 10 9 2
22 10 0 9 1 11 11 11 13 1 12 16 11 12 15 13 9 1 10 9 1 11 2
45 11 11 2 1 10 0 9 11 11 13 10 12 9 12 1 11 2 11 2 13 10 9 1 10 9 1 10 9 0 1 10 9 1 10 9 12 2 10 9 13 3 0 16 9 2
20 10 9 1 10 11 13 1 12 9 0 7 1 9 13 1 10 0 9 0 2
18 1 3 1 9 2 13 10 9 1 9 7 9 0 1 10 0 2 5
40 13 3 1 10 9 0 2 15 13 1 10 0 9 0 7 0 1 12 2 9 1 9 1 10 9 1 11 1 11 3 1 10 9 1 10 9 1 11 2 2
16 3 1 10 9 2 10 9 4 13 1 13 10 9 1 9 2
17 10 9 0 2 9 2 13 10 9 0 0 12 9 1 10 9 2
20 15 14 13 3 1 10 9 1 10 9 15 10 9 4 4 13 1 10 9 2
21 10 9 13 10 10 9 1 11 2 1 11 2 1 11 2 1 11 7 1 11 2
7 15 13 10 12 9 12 2
36 1 12 5 1 10 9 12 2 15 4 13 1 12 5 1 10 9 12 2 16 15 1 10 9 1 10 11 4 13 1 12 5 1 12 5 2
16 9 1 12 7 1 12 1 12 2 15 13 3 11 1 12 2
16 7 2 1 1 10 9 1 10 9 2 4 13 3 4 13 2
13 15 4 13 15 1 10 9 7 15 1 10 9 2
20 9 13 1 10 9 16 10 10 9 15 13 1 11 4 13 1 10 9 0 2
8 11 13 10 9 1 10 11 2
24 10 11 15 13 12 1 12 9 1 10 0 9 1 11 2 12 9 2 2 9 1 10 9 2
16 15 13 1 3 10 9 1 10 9 11 11 2 10 11 2 2
23 10 9 1 9 2 13 3 1 10 11 2 4 13 10 9 1 10 9 7 1 10 9 2
18 11 4 13 3 1 9 2 1 10 9 15 10 0 9 0 15 13 2
40 15 13 3 0 2 7 13 3 12 9 0 2 15 4 4 13 10 9 7 10 9 2 0 1 10 12 9 0 1 10 9 1 10 9 2 9 7 9 2 2
22 15 13 9 1 13 16 10 9 9 1 10 9 13 1 15 15 13 3 1 12 9 2
24 10 9 1 10 11 0 13 1 10 9 1 9 4 4 4 13 1 10 9 1 10 9 12 2
17 10 11 1 11 7 11 13 3 1 10 9 1 10 9 1 9 2
26 2 3 2 1 10 9 1 9 2 3 1 10 9 1 10 9 0 2 15 4 13 10 9 1 9 2
8 10 11 13 0 1 1 12 2
54 15 13 10 9 1 10 9 0 1 11 2 7 2 1 4 13 10 9 11 1 15 15 13 2 13 10 9 1 10 9 0 2 10 9 1 11 2 2 1 10 9 1 10 9 0 2 2 1 10 9 0 1 11 2
23 10 9 1 10 9 1 10 9 13 3 15 13 1 10 9 1 10 9 7 1 15 13 2
55 1 9 0 2 15 13 3 10 9 1 10 11 1 10 11 1 13 1 12 2 3 13 1 10 0 9 0 7 0 2 1 15 10 9 11 2 10 9 0 7 10 11 1 10 11 2 1 15 15 13 3 1 12 9 2
38 10 9 2 13 9 0 1 10 11 2 11 2 7 2 3 3 2 9 1 10 11 2 4 13 1 9 10 9 8 7 10 9 8 1 10 9 8 2
45 3 16 10 9 13 10 9 1 3 1 3 0 2 9 13 2 9 0 2 9 13 2 16 9 2 2 10 11 4 15 13 1 10 12 9 0 7 3 10 9 0 13 1 9 2
18 1 10 9 1 12 9 2 11 13 1 10 9 1 11 11 1 11 2
24 10 12 1 9 4 13 1 10 11 11 1 11 13 1 11 11 1 9 1 10 9 1 11 2
9 15 13 1 9 0 2 3 0 2
43 10 9 1 10 9 1 10 11 13 3 1 9 6 13 10 9 1 11 1 10 9 2 1 10 9 1 10 9 1 10 9 2 15 13 9 1 4 15 13 9 1 11 2
9 15 4 13 3 1 10 11 8 12
9 9 4 3 13 1 10 9 9 2
11 10 9 1 10 9 0 3 13 1 3 2
12 10 9 13 0 1 10 9 1 11 1 11 2
25 10 9 16 10 9 4 4 13 7 13 1 10 9 1 9 2 10 9 0 4 4 13 10 9 2
39 3 2 1 11 2 10 9 14 13 3 10 9 0 1 10 9 2 7 3 10 2 9 0 2 1 10 9 15 15 4 13 1 10 11 2 7 11 2 2
30 10 9 1 15 4 13 10 9 13 1 10 12 9 7 4 4 13 1 10 9 1 10 9 1 10 12 7 12 9 2
18 10 9 15 13 2 2 7 10 9 3 15 13 0 16 9 4 13 2
14 15 4 13 1 2 9 1 9 0 2 2 9 2 2
17 10 9 1 10 9 4 3 13 1 10 9 1 9 13 1 12 2
114 1 3 10 3 0 9 0 1 10 9 1 10 11 2 10 9 4 4 13 1 12 12 1 11 10 9 1 10 9 1 10 11 1 10 9 2 2 10 9 1 12 5 1 10 9 1 10 9 1 12 7 12 2 7 10 0 9 1 9 0 1 10 9 1 10 9 0 1 11 1 10 11 2 9 1 12 5 1 10 9 13 1 10 9 0 2 9 1 12 9 1 9 1 12 1 12 1 12 2 4 13 10 9 0 1 15 13 1 10 11 1 10 11 2
35 11 11 4 13 10 11 1 13 10 9 0 1 9 7 1 9 1 10 9 0 1 10 9 1 10 9 1 10 11 1 10 9 0 0 2
21 1 10 9 1 9 2 10 9 1 10 9 11 4 13 3 1 12 9 1 9 2
30 1 10 12 9 1 10 9 15 4 13 10 9 12 9 1 9 2 2 10 9 1 10 9 2 15 4 13 1 11 2
7 7 15 15 4 13 3 2
26 10 11 4 3 13 10 9 0 1 10 9 0 7 0 7 10 9 14 4 3 3 13 10 9 0 2
18 1 9 12 10 11 12 4 13 1 10 9 0 11 2 11 11 2 2
21 15 15 13 1 10 9 1 10 12 0 9 1 10 0 9 0 11 11 7 11 2
15 10 9 1 10 9 4 13 3 13 10 9 1 10 9 2
17 10 9 1 9 4 13 1 1 10 9 0 1 10 9 1 11 2
27 7 10 9 15 13 10 0 9 1 9 4 13 10 9 1 10 9 3 0 7 1 10 9 15 15 13 2
48 13 1 10 9 1 10 9 1 10 9 0 7 13 1 10 9 0 1 10 9 10 3 0 2 11 11 4 13 1 10 9 3 1 13 10 9 1 10 11 7 13 10 9 1 10 9 0 2
18 6 1 10 9 1 11 1 10 9 0 1 10 0 9 1 10 9 2
53 1 13 10 9 1 9 1 9 2 3 1 9 1 10 9 2 1 10 9 0 1 10 9 2 7 3 3 1 10 3 0 1 10 9 7 3 1 10 9 2 10 9 1 9 1 9 7 4 14 13 3 0 2
15 15 4 4 13 1 9 1 12 2 7 13 3 12 9 2
15 10 0 9 11 13 11 1 11 3 9 1 11 1 12 2
12 1 12 2 10 9 13 1 9 1 10 11 2
17 1 10 0 9 11 11 13 12 5 1 10 9 2 12 5 2 2
22 3 2 10 9 14 13 3 1 10 9 15 10 0 9 1 10 0 0 4 13 13 2
30 15 13 9 1 10 11 7 1 10 11 1 12 7 12 2 1 15 15 13 10 9 1 10 9 1 10 9 1 12 2
15 3 2 15 13 10 9 0 1 13 10 9 1 10 9 2
17 11 13 9 1 11 7 9 0 7 0 9 1 10 9 1 11 2
25 10 9 13 1 10 9 0 10 9 1 10 9 0 2 1 15 1 10 9 0 15 13 10 9 2
18 3 1 10 9 1 12 2 10 10 9 1 0 9 4 13 7 13 2
17 1 12 2 15 13 9 0 7 13 1 10 9 0 0 1 12 2
13 11 11 1 9 0 13 15 3 9 1 10 11 2
43 1 10 9 0 2 11 2 1 9 0 11 2 11 2 2 9 1 11 7 1 11 2 9 1 11 7 9 1 11 10 11 7 1 11 2 13 9 1 10 9 1 11 2
21 11 11 4 4 13 1 10 9 11 11 11 1 12 1 10 9 0 1 11 11 2
34 10 9 0 4 13 9 1 12 1 10 9 1 10 11 15 10 11 11 11 11 4 1 9 13 10 2 9 1 10 11 0 0 2 2
59 10 9 1 10 11 2 7 9 2 15 13 1 10 9 0 1 10 9 2 9 2 2 7 10 9 11 13 4 13 1 10 9 1 10 9 0 2 10 9 13 10 9 11 0 3 15 13 13 12 9 1 15 10 9 11 0 4 13 2
15 10 9 13 10 9 1 10 9 1 10 9 1 10 9 2
52 1 3 2 10 11 4 13 10 10 9 1 13 1 9 2 1 10 9 1 10 9 0 7 10 0 9 15 15 13 9 2 1 16 10 9 4 13 1 10 9 1 10 9 1 10 9 1 10 9 3 0 2
24 10 9 1 10 11 2 3 9 11 2 13 1 12 2 13 10 9 1 10 12 9 1 11 2
30 16 15 13 1 10 9 7 16 15 15 13 9 1 13 1 10 9 1 10 9 2 4 15 13 1 10 9 1 11 2
15 10 9 13 0 2 7 10 9 13 10 0 9 1 9 2
21 15 13 1 10 9 1 10 0 9 16 11 11 4 13 1 10 9 15 15 13 2
15 1 10 9 1 10 9 2 15 3 13 3 7 1 15 13
30 15 13 11 11 1 13 10 9 15 4 13 1 13 10 11 0 1 10 9 1 9 1 10 0 9 1 10 9 0 2
35 11 2 10 11 4 13 10 0 9 1 13 1 10 9 1 10 9 1 15 13 1 13 9 2 9 7 9 2 4 13 9 10 11 11 2
18 10 9 1 10 11 7 10 11 13 10 9 13 10 11 7 10 11 2
33 15 1 10 9 1 10 9 1 11 11 2 15 13 16 15 13 10 0 9 1 10 9 1 10 9 1 10 9 1 10 11 0 2
21 15 14 15 13 3 1 13 13 10 9 2 7 3 1 13 10 9 1 10 9 2
16 3 13 1 10 9 1 10 9 2 15 4 13 10 9 0 2
14 10 9 1 10 11 13 10 9 1 10 11 0 0 2
19 10 11 11 1 11 13 10 9 13 1 10 9 1 10 11 7 10 11 2
31 15 13 3 13 1 12 2 1 10 9 1 12 9 1 1 10 9 1 10 9 1 12 2 15 13 10 9 1 12 9 2
13 13 10 9 0 2 15 13 10 9 1 9 13 2
11 10 9 1 10 9 13 10 9 1 9 2
33 10 9 13 4 3 13 1 10 9 1 13 16 10 9 13 1 10 9 3 1 10 11 13 1 10 9 15 4 13 1 10 9 2
37 13 1 10 9 0 0 2 11 11 11 11 1 11 13 10 9 1 11 11 11 11 2 9 1 11 2 12 2 7 11 11 10 9 1 10 11 2
18 10 9 15 13 10 9 2 1 9 16 10 9 15 13 13 3 0 2
18 3 1 10 0 9 0 1 12 2 15 15 13 1 11 7 1 11 2
37 11 1 11 13 10 9 7 10 9 0 1 9 1 10 12 9 2 15 10 9 15 13 1 10 9 1 10 9 0 7 10 9 1 10 0 11 2
39 15 3 13 10 0 9 1 1 11 2 7 10 9 7 10 9 2 13 1 10 9 1 10 9 1 9 0 2 4 13 1 10 9 7 13 1 10 9 2
43 9 11 4 13 9 10 9 1 1 13 10 0 12 9 1 13 11 11 2 15 10 9 1 9 15 4 13 10 12 9 1 10 9 1 10 9 1 10 9 1 10 11 2
14 10 9 0 15 13 1 10 9 1 9 7 1 9 2
37 15 15 13 1 12 10 0 9 1 11 1 12 9 1 10 9 1 10 9 2 15 13 1 10 9 10 9 1 10 9 0 1 10 9 1 11 2
37 10 0 12 9 2 15 13 10 11 0 12 15 13 1 10 9 10 9 13 10 9 1 10 10 9 0 1 9 1 11 2 13 3 3 10 9 2
27 3 16 15 13 0 1 15 13 1 12 9 1 10 9 16 12 9 13 1 10 9 13 3 1 9 0 2
40 10 9 13 1 10 9 1 10 11 7 1 10 11 15 2 1 15 4 13 1 10 11 2 13 10 11 2 13 10 11 1 12 2 13 1 11 3 1 11 2
20 10 11 13 10 9 9 1 10 9 1 10 11 1 10 9 1 12 1 12 2
36 11 15 13 3 10 9 0 16 15 13 1 10 9 10 9 11 1 11 2 13 1 11 1 10 9 6 13 10 9 1 10 9 1 10 11 2
45 7 10 9 1 9 4 13 7 15 13 1 10 9 1 9 1 15 13 12 9 2 13 16 15 4 13 10 9 1 10 9 0 2 7 15 13 10 9 15 15 13 10 12 9 2
11 3 12 9 12 15 13 15 12 8 12 2
24 13 11 11 7 9 11 2 11 11 4 13 1 15 1 10 0 9 1 10 9 1 10 11 2
27 15 3 4 13 16 10 2 9 1 10 9 0 13 10 9 2 1 10 9 1 10 9 2 9 2 2 2
18 3 15 15 13 1 10 9 1 12 7 4 13 1 10 11 11 11 2
14 11 2 12 9 2 13 9 1 10 9 1 12 9 2
15 10 9 0 7 10 9 15 13 3 3 1 9 1 11 2
18 11 13 10 9 0 2 13 1 10 9 1 10 11 7 10 9 11 2
10 9 6 0 7 3 0 1 10 9 2
16 10 9 13 10 9 0 7 0 1 10 9 7 1 9 13 2
19 10 9 3 13 1 10 9 13 11 12 1 13 10 9 1 9 1 11 2
29 1 10 9 10 9 0 2 13 1 12 2 15 13 2 2 15 4 13 15 15 13 10 15 2 15 4 4 13 2
12 10 9 0 14 4 3 13 9 1 10 9 2
19 3 2 10 9 13 10 11 11 1 12 9 1 10 9 1 11 11 11 2
24 11 14 13 3 10 9 6 13 10 9 1 9 14 4 3 13 1 10 9 1 10 11 11 2
15 15 4 13 10 0 9 1 10 9 0 1 10 9 0 2
19 15 3 13 1 10 12 9 1 10 9 16 1 10 12 9 12 3 3 2
22 9 0 1 10 9 2 15 13 12 9 2 15 10 3 9 7 3 0 13 1 12 2
32 10 9 13 1 10 9 1 10 9 10 9 1 10 9 1 10 11 1 11 2 13 10 9 0 1 10 9 1 10 11 0 2
11 15 4 13 1 12 1 11 1 11 11 2
26 13 10 9 13 13 10 9 2 13 1 13 10 9 7 15 15 13 15 3 2 1 10 9 7 9 2
26 15 13 1 10 9 1 10 9 11 1 10 11 1 11 11 2 12 2 1 11 11 7 11 11 2 2
20 15 13 10 9 1 14 3 4 3 13 10 9 1 5 1 10 9 10 9 2
46 10 12 9 12 2 9 1 10 9 2 10 9 0 1 9 2 11 2 13 2 1 3 13 10 9 2 10 11 11 1 10 9 0 1 11 15 15 13 1 13 1 10 9 1 12 2
4 11 15 13 2
94 7 1 10 9 1 10 12 9 2 3 1 10 9 1 10 9 1 11 13 10 9 1 9 7 10 9 1 10 11 0 2 10 9 1 10 9 0 15 13 3 1 3 7 10 9 3 0 2 3 16 10 9 1 10 9 13 3 3 0 2 4 13 1 10 9 7 10 9 2 15 13 10 9 3 0 2 10 9 2 10 9 1 9 7 10 9 2 1 10 9 7 10 9 2
11 11 11 2 12 2 0 13 1 0 9 2
71 10 9 4 13 1 10 9 1 10 9 11 2 12 9 2 7 10 9 1 11 2 12 9 2 2 1 10 9 1 10 9 1 11 2 12 9 2 7 10 9 1 10 11 2 12 9 2 2 7 1 10 9 1 10 11 11 2 12 9 2 7 10 9 1 10 11 2 12 9 2 2
36 1 9 1 10 9 7 10 9 0 1 10 9 2 15 4 3 13 1 10 9 1 2 9 11 2 2 0 9 13 1 10 9 12 1 11 2
11 10 12 9 13 13 10 9 1 12 9 2
35 2 2 2 10 9 2 15 13 1 0 9 10 9 0 1 15 13 3 1 10 9 2 4 13 10 9 1 9 7 13 9 1 10 9 2
21 10 9 13 9 1 9 0 13 1 10 11 11 11 1 15 1 10 9 1 9 2
20 10 9 4 4 13 1 12 1 10 9 1 11 1 10 9 1 10 11 11 2
51 10 9 0 13 1 13 13 7 13 10 9 0 13 1 11 10 9 1 9 0 3 13 7 10 9 1 9 1 15 10 9 4 13 7 13 1 10 2 0 0 11 2 15 15 4 0 13 3 10 9 2
9 15 13 3 10 9 1 11 11 2
18 10 9 13 10 9 0 3 0 7 3 0 2 4 13 10 10 9 2
9 1 12 13 10 9 11 11 11 2
27 15 15 13 1 11 2 15 15 13 10 9 1 9 0 2 3 1 11 2 15 15 15 13 1 11 11 2
42 10 9 0 1 10 9 1 11 4 13 1 10 9 0 2 3 0 2 13 1 9 7 1 10 9 3 16 1 10 9 1 9 13 1 12 1 10 9 1 10 9 2
25 10 9 0 15 13 3 1 10 9 0 2 15 15 13 10 9 7 0 9 1 10 9 1 9 2
34 10 9 14 13 0 16 1 10 9 1 12 9 2 1 12 9 3 2 2 7 15 4 13 1 10 0 9 1 9 1 10 9 0 2
19 11 1 11 2 11 13 10 0 9 1 10 9 1 9 9 0 11 11 2
18 15 13 1 10 9 16 10 9 0 7 1 9 1 10 9 15 13 2
36 11 11 11 2 13 10 12 9 12 1 11 2 11 0 2 13 10 9 0 1 0 9 1 10 9 15 4 13 10 9 1 9 0 1 12 2
14 11 13 10 9 2 15 13 10 9 2 15 13 0 2
25 12 5 2 16 9 2 4 13 10 9 0 7 0 7 3 9 2 16 12 5 2 4 4 13 2
13 1 10 9 2 10 9 13 10 9 7 10 9 2
18 10 9 2 13 1 11 2 13 3 0 2 10 9 13 10 0 9 2
31 10 9 13 9 1 9 2 15 13 1 13 1 15 0 1 16 10 9 4 4 13 1 13 16 15 13 3 9 1 11 2
43 1 10 9 1 10 11 2 1 12 1 12 9 2 9 9 2 7 1 12 9 1 10 9 2 15 13 0 1 10 9 0 16 1 10 9 0 1 10 11 1 10 11 2
21 10 9 1 9 13 16 10 11 4 13 10 9 1 10 9 0 1 13 10 9 2
37 1 10 9 2 1 9 1 10 9 2 15 13 3 1 10 9 15 15 13 10 9 1 9 1 1 10 11 11 0 2 10 9 1 10 9 0 2
13 10 9 13 10 11 1 11 7 1 11 1 11 2
19 11 11 2 13 10 12 9 12 1 11 1 10 11 2 13 10 9 0 2
24 1 12 2 3 1 11 1 9 2 15 13 10 9 1 9 1 9 1 10 9 0 1 11 2
8 10 9 15 13 1 10 9 2
29 1 10 9 1 10 9 2 10 9 0 15 13 1 10 9 2 3 3 16 10 10 9 0 15 13 1 10 9 2
38 11 11 13 10 9 7 9 0 2 13 11 11 11 1 11 2 11 2 10 12 9 12 2 13 1 10 9 1 11 11 2 11 2 10 12 9 12 2
18 10 9 1 13 1 10 9 15 14 13 10 9 3 1 10 9 13 2
19 10 9 1 10 9 7 10 9 15 13 1 10 10 9 3 0 1 9 2
56 15 13 3 3 13 10 9 2 10 9 0 2 7 13 10 9 0 2 9 2 2 10 0 9 1 15 13 13 16 15 14 13 3 1 9 1 10 9 1 10 9 1 0 15 13 10 9 8 1 10 9 0 1 8 2 2
12 3 2 10 9 1 9 13 1 0 9 2 2
15 11 11 4 3 1 15 13 2 2 11 2 15 4 13 2
7 9 13 10 9 1 11 2
20 15 13 1 9 1 11 2 3 10 11 11 3 1 13 10 11 1 11 11 2
44 11 11 2 12 2 13 10 9 2 4 3 1 10 11 11 0 2 13 1 10 9 1 10 9 7 9 0 0 2 1 10 9 1 10 9 1 10 11 1 10 11 1 12 2
32 11 13 10 9 13 16 11 2 1 10 9 1 10 9 1 10 9 2 14 15 13 3 7 15 13 3 16 15 4 15 13 2
34 15 13 2 1 9 7 1 9 2 10 9 0 2 1 12 9 7 15 13 1 10 9 2 15 0 13 1 10 0 9 1 0 9 2
33 1 10 9 2 10 12 9 1 10 11 1 11 7 1 10 9 1 11 13 10 9 1 9 7 1 9 7 13 9 1 10 11 2
30 15 4 3 13 10 9 1 10 11 1 11 12 2 10 9 1 10 11 1 11 12 7 13 12 1 11 10 0 9 2
14 10 0 0 9 1 10 9 13 11 11 7 11 11 2
32 11 11 13 10 9 0 13 10 12 9 12 1 11 11 2 11 11 2 11 2 2 13 10 12 9 12 1 11 2 11 2 2
38 10 9 1 10 9 0 1 13 1 10 9 13 3 10 9 2 15 13 3 3 10 9 1 10 11 1 11 2 7 3 1 10 11 7 1 10 11 2
24 9 13 2 9 2 0 0 9 9 2 16 1 9 2 2 9 1 9 0 1 9 0 2 2
34 1 10 0 9 7 1 13 10 9 1 10 9 1 10 9 2 10 9 0 0 4 13 1 10 9 12 10 9 0 1 10 9 0 2
27 10 9 13 13 3 10 9 2 10 10 9 2 10 10 9 2 10 9 2 10 9 7 10 10 9 13 2
22 10 9 13 10 9 0 1 16 10 9 0 1 10 9 4 13 1 9 0 1 11 2
12 15 13 0 1 1 10 9 1 10 11 11 2
14 10 12 9 12 2 15 13 10 9 1 10 9 0 2
11 13 1 10 9 13 3 3 10 0 9 2
56 11 11 2 13 1 9 12 1 10 9 1 11 2 11 2 2 13 10 9 0 1 10 9 0 1 11 2 15 13 10 15 1 10 0 9 1 10 9 0 0 1 1 13 10 9 2 7 13 9 1 11 1 12 1 12 2
33 9 4 13 1 10 0 9 1 10 9 0 2 1 10 12 7 1 10 12 2 1 10 9 3 16 1 10 0 9 1 9 0 2
31 10 9 1 11 14 13 3 10 9 0 1 10 9 1 10 9 7 2 7 1 10 9 1 9 2 1 9 7 1 9 2
19 10 9 0 13 1 10 9 10 3 0 2 13 2 9 1 10 9 2 2
16 15 13 1 13 10 9 0 2 1 10 9 15 4 13 0 2
30 10 9 4 4 13 10 1 10 12 9 12 9 12 2 7 4 4 13 1 10 9 12 1 12 3 1 13 10 9 2
9 15 4 4 13 1 10 9 0 2
20 15 15 13 3 1 10 9 0 2 0 1 10 9 0 1 10 9 7 9 2
27 10 9 11 2 15 13 1 10 9 1 11 7 11 2 7 1 15 1 11 7 11 2 13 10 12 9 2
28 10 9 1 10 9 1 9 1 10 9 4 13 7 15 15 4 13 2 2 15 13 15 15 15 13 2 2 2
14 11 11 11 2 12 2 12 2 12 2 12 9 2 2
12 11 15 13 3 1 10 9 3 0 7 0 2
22 11 13 1 10 9 12 1 10 11 1 11 1 10 9 1 9 0 0 1 10 11 2
23 10 9 1 10 9 1 9 1 11 7 9 13 10 9 1 9 1 9 0 7 1 9 2
24 16 10 9 13 0 2 11 11 13 1 2 12 9 2 10 9 1 10 11 7 10 9 2 2
25 15 4 13 1 11 3 1 10 9 0 12 1 10 11 1 11 2 1 10 9 1 10 11 2 2
53 16 2 15 15 13 0 2 10 12 9 0 13 1 10 9 1 10 9 7 16 10 9 13 10 9 1 9 0 0 2 10 9 1 10 9 1 10 9 11 15 13 0 7 2 1 9 0 2 10 9 1 15 2
15 10 9 0 1 10 11 15 4 13 10 9 1 10 9 2
18 11 11 2 13 10 12 9 12 1 11 2 13 10 9 0 0 0 2
20 2 11 11 2 13 10 0 9 1 10 0 9 9 1 11 1 10 0 9 2
23 3 1 10 9 1 10 9 9 2 9 15 13 10 9 1 10 11 1 15 1 10 11 2
26 1 10 9 1 10 12 9 2 10 9 1 11 2 11 11 11 2 13 1 11 2 13 10 9 11 2
9 1 11 2 15 15 13 3 12 2
18 10 9 2 1 9 3 2 4 13 1 12 12 1 9 1 9 11 2
14 13 3 10 9 2 10 9 7 9 1 10 9 0 2
22 10 9 13 1 10 12 9 13 1 9 6 13 10 9 1 10 12 9 2 9 2 2
14 10 9 4 13 1 10 9 1 12 9 2 12 2 2
31 1 9 2 10 11 11 11 13 10 0 9 1 10 9 1 10 11 1 10 9 0 1 10 12 9 13 1 9 1 9 2
27 15 13 10 9 0 1 9 1 11 2 3 1 10 11 0 2 12 2 7 10 11 0 2 9 12 2 2
14 10 9 1 11 13 1 9 1 10 12 9 1 9 2
48 10 9 1 9 1 10 11 0 7 10 9 0 3 0 2 10 3 0 2 1 10 9 2 9 0 2 13 10 9 0 1 10 9 2 15 13 10 9 0 15 13 1 10 9 1 10 9 2
20 1 12 2 10 9 1 10 11 11 11 11 2 12 2 4 13 1 10 9 2
8 15 13 9 0 1 10 9 2
23 11 11 1 11 2 7 11 11 2 4 13 10 0 9 1 11 2 1 10 9 1 11 2
51 10 9 0 1 10 11 2 4 13 1 10 9 1 9 1 10 9 0 2 13 3 10 9 1 9 2 1 15 1 10 9 13 1 11 7 11 11 2 3 1 10 9 1 10 9 1 10 0 9 0 2
36 3 2 3 16 11 13 1 10 9 1 10 9 12 1 13 10 9 9 0 2 10 9 1 10 9 9 14 4 13 1 10 9 13 1 11 2
14 1 12 15 4 13 7 15 13 3 2 1 11 2 2
21 3 2 10 9 0 11 11 2 15 13 10 9 1 10 11 1 9 2 13 2 2
30 10 9 1 11 14 4 13 3 1 10 9 0 1 11 2 11 2 11 12 2 7 11 2 1 1 2 11 12 2 2
70 15 4 3 13 1 9 10 11 8 8 11 2 10 9 1 10 9 1 10 11 11 2 2 10 9 15 15 4 13 1 12 9 2 10 0 9 1 12 9 12 7 12 9 12 1 10 9 0 1 11 11 7 10 12 0 9 2 12 7 12 9 12 1 10 9 0 1 11 11 2
21 10 0 9 1 10 9 2 11 12 13 1 11 2 4 13 1 10 11 1 12 2
27 15 4 3 13 1 10 9 0 2 1 9 1 14 3 13 10 9 3 3 0 1 15 1 10 8 8 2
25 15 13 3 13 10 0 9 1 10 9 1 10 9 7 10 9 16 15 4 13 1 13 10 9 2
15 10 0 9 2 15 13 10 9 0 2 13 1 10 9 2
37 9 2 10 9 1 10 9 4 13 10 9 4 4 13 10 9 2 7 2 1 10 12 9 1 10 9 2 15 13 10 9 15 15 4 13 9 2
25 3 10 9 9 13 1 10 9 15 15 15 13 10 10 9 1 9 2 10 10 9 1 10 9 2
29 10 9 4 13 1 11 11 2 9 2 2 11 11 2 9 2 2 11 11 2 9 2 7 11 11 2 9 2 2
23 10 9 13 10 9 1 9 7 15 15 4 4 13 1 10 9 1 16 15 15 4 13 2
14 10 9 15 13 1 10 9 12 1 10 9 12 9 2
20 11 4 13 1 11 2 11 2 3 11 1 11 2 1 10 9 1 9 0 2
16 15 13 1 13 10 9 1 9 1 15 13 1 10 9 0 2
34 13 10 9 1 10 9 2 10 9 15 13 1 10 9 0 7 15 15 13 3 1 10 9 0 1 10 9 0 15 11 13 3 9 2
12 10 11 11 13 10 9 0 2 13 10 9 2
15 15 13 10 0 9 1 9 0 1 10 9 1 10 9 2
36 15 4 13 1 10 9 1 9 2 13 10 9 1 10 11 7 10 9 0 1 11 13 1 10 11 2 10 9 13 1 9 7 1 9 9 2
28 10 9 4 13 1 10 9 1 10 11 10 9 3 0 3 1 13 3 10 9 1 9 2 1 9 7 9 2
20 10 9 1 9 4 4 13 1 10 11 1 10 9 1 10 9 0 1 11 2
16 10 9 1 10 9 13 1 10 9 1 10 9 1 10 9 2
14 15 4 4 13 1 1 9 1 10 9 1 10 11 2
22 10 9 1 10 9 11 11 11 11 11 4 3 13 12 9 1 10 9 1 10 9 2
46 10 0 9 7 9 1 10 9 1 10 11 2 1 11 0 2 13 10 9 1 10 9 1 10 11 0 1 10 11 2 11 2 1 10 9 1 10 9 1 10 11 1 10 11 0 2
32 10 9 4 13 1 10 9 1 12 5 1 10 9 7 10 9 1 12 5 3 16 12 5 1 10 9 13 10 12 9 0 2
20 10 11 11 4 13 1 10 9 1 12 1 13 10 11 1 10 11 1 11 2
40 9 0 1 10 9 0 1 9 12 2 11 11 13 3 10 9 1 10 11 10 12 9 12 16 10 9 11 11 4 13 1 10 9 1 10 9 1 9 0 2
15 15 14 13 3 10 9 7 10 9 0 13 1 10 9 2
25 1 3 2 15 4 4 13 1 13 11 10 9 2 1 9 1 10 9 0 1 10 9 1 9 2
22 16 15 15 13 2 3 11 11 12 14 4 13 1 9 10 9 1 10 9 1 9 2
9 10 9 1 9 13 3 3 0 2
40 15 4 13 1 2 11 2 11 11 2 2 10 9 1 9 3 0 15 13 1 9 1 10 9 2 13 1 9 13 1 9 0 7 1 9 1 10 9 0 2
32 15 14 13 3 3 0 1 13 10 9 2 13 15 15 15 13 3 7 10 9 1 10 9 16 15 4 13 1 10 9 11 2
33 11 11 13 10 9 1 9 2 10 11 11 2 15 13 10 9 1 10 0 9 2 3 13 1 10 9 1 10 11 11 1 11 2
18 7 10 9 3 2 13 10 9 0 15 14 15 13 3 1 10 9 2
24 10 9 1 11 4 13 3 0 2 12 5 2 7 3 0 2 12 5 2 1 10 0 9 2
22 1 10 9 1 9 2 10 9 13 10 9 2 13 1 10 9 1 9 1 12 9 2
16 11 15 13 3 1 10 9 2 13 11 7 13 11 1 9 2
28 10 9 3 3 2 15 13 1 13 10 9 1 9 10 9 2 3 1 13 10 9 9 7 9 1 10 9 2
32 2 10 9 1 10 11 13 16 10 9 0 4 13 1 13 9 1 10 10 9 2 1 9 1 10 9 2 2 13 10 9 2
75 10 9 1 15 11 13 15 1 10 9 15 13 10 9 1 3 16 11 13 9 1 10 11 1 11 2 1 15 10 9 13 10 9 16 10 9 13 1 9 1 10 9 10 9 0 1 10 9 7 16 10 11 14 13 15 1 9 1 10 9 7 1 11 2 7 13 3 1 10 9 0 1 10 9 2
54 1 9 2 1 10 9 1 10 9 0 2 10 9 0 13 1 13 10 9 7 16 15 4 13 1 13 10 9 1 9 7 9 2 15 4 13 15 15 15 13 10 9 2 3 13 2 15 4 13 10 9 1 9 2
34 10 9 1 10 9 0 7 10 9 0 1 10 9 2 9 1 9 2 7 10 9 2 9 1 14 2 13 10 9 1 9 0 0 2
20 15 13 10 0 9 1 10 9 0 10 9 0 7 10 9 0 11 11 11 2
23 1 12 2 15 4 13 1 10 9 0 1 11 11 1 10 0 9 2 12 2 12 2 2
38 11 11 11 7 9 1 10 9 2 9 13 1 10 9 1 10 9 1 9 0 2 13 10 9 13 1 10 9 1 10 9 1 11 2 1 9 0 2
27 10 0 9 13 0 7 0 13 1 10 9 0 2 1 10 11 1 10 11 1 10 11 1 10 11 2 2
9 3 13 3 3 10 9 1 9 2
10 11 11 2 12 2 13 10 9 0 2
16 9 1 9 7 9 2 15 13 1 10 9 11 1 10 11 2
24 1 10 9 1 10 9 0 1 9 12 2 11 11 2 11 2 4 4 13 9 1 10 9 2
36 10 9 0 2 9 1 10 9 1 10 0 9 1 11 2 4 13 10 9 0 1 10 9 1 9 2 15 10 9 13 1 0 9 12 9 2
32 10 9 13 0 1 9 7 9 1 10 9 1 0 9 3 16 1 10 9 1 12 9 2 10 9 13 0 1 10 9 9 2
23 10 9 13 1 10 0 9 1 10 11 13 10 9 1 10 9 11 1 9 12 1 12 2
8 10 9 15 13 3 1 9 2
9 9 1 9 1 10 9 1 9 2
14 15 13 3 10 9 1 9 1 1 10 9 1 12 2
30 11 11 13 3 10 9 1 10 9 1 10 9 7 10 9 1 10 9 0 1 10 11 2 13 10 9 1 10 9 2
22 1 3 2 10 9 0 1 10 11 1 10 9 4 4 13 1 10 9 0 1 11 2
55 3 16 15 4 13 10 9 2 11 2 11 13 0 7 4 13 10 0 9 1 11 11 2 1 11 11 2 10 9 2 3 0 2 3 0 7 3 13 7 1 10 9 9 10 9 13 15 15 9 2 2 3 2 2 2
28 15 13 1 10 9 1 9 0 7 13 1 9 1 10 0 9 10 9 13 9 0 13 1 10 9 1 12 2
13 10 11 1 11 13 10 9 0 0 1 9 0 2
17 1 12 2 10 11 13 10 9 1 9 1 10 9 1 10 9 2
13 1 1 12 2 10 9 0 1 11 13 10 9 2
34 10 11 14 13 3 3 1 9 0 10 9 1 9 2 3 15 13 9 1 10 9 1 10 9 0 15 15 4 13 10 9 1 9 2
23 1 10 9 0 2 10 9 1 9 13 0 7 15 13 2 15 13 1 2 1 10 9 2
48 10 9 4 4 3 13 1 11 11 2 9 1 10 9 0 1 10 9 2 5 16 1 11 11 2 9 7 9 2 15 2 1 10 9 1 10 9 4 13 10 9 1 9 13 1 10 9 2
39 10 9 1 10 12 9 12 13 10 0 9 0 0 2 12 9 2 2 16 10 9 11 11 4 4 13 1 10 9 2 12 5 2 0 1 10 9 0 2
36 10 9 1 10 9 0 1 10 9 1 10 9 4 13 1 10 9 1 10 9 1 13 10 9 1 10 9 7 3 13 10 0 9 1 13 2
16 11 11 2 13 10 12 9 12 1 11 2 13 10 9 0 2
