735 17
9 0 0 9 4 13 14 11 11 2
3 8 8 2
6 6 2 3 13 0 2
10 3 4 15 13 2 3 4 15 13 2
27 11 0 9 0 9 4 13 2 16 4 0 9 1 0 9 0 0 9 13 0 0 9 1 9 11 11 2
19 0 0 9 13 0 2 16 13 0 9 10 9 7 9 1 3 0 9 2
14 0 9 0 9 13 3 11 2 0 9 7 13 11 2
37 11 1 11 1 11 1 0 14 4 13 14 9 2 0 9 0 9 3 1 0 9 2 9 1 9 13 14 1 0 9 1 9 3 0 0 9 2
37 1 10 9 13 0 9 11 11 7 11 11 2 9 9 0 9 2 3 1 11 13 0 7 0 9 2 16 13 12 1 12 0 0 9 10 9 2
9 13 4 9 9 7 12 12 9 2
44 9 9 11 13 9 9 1 9 7 9 2 16 15 1 9 1 9 9 9 1 9 1 9 12 13 9 1 9 9 0 9 1 9 0 9 2 16 15 4 13 9 0 9 2
15 9 13 9 9 1 9 10 9 1 3 0 9 1 9 2
19 11 11 2 11 13 3 0 9 1 9 2 16 13 0 0 7 0 9 2
12 9 13 2 16 0 9 13 9 1 0 9 2
21 13 15 15 2 16 1 11 14 13 3 13 10 9 9 2 16 13 1 0 9 2
4 16 13 9 2
21 1 11 13 1 10 9 0 9 7 9 2 4 7 15 13 3 13 0 9 9 2
11 9 7 9 0 9 13 1 15 3 0 2
10 0 9 14 13 9 7 9 0 9 2
26 9 13 9 2 1 15 4 3 13 7 3 13 9 1 0 9 7 3 0 9 7 9 9 7 9 2
19 10 9 3 13 9 14 1 12 9 2 16 15 1 0 9 14 13 13 2
12 0 9 4 13 13 0 9 7 13 10 9 2
11 1 15 13 13 9 1 0 7 0 9 2
23 9 13 13 14 0 9 2 1 9 1 0 9 2 16 4 9 1 10 9 13 0 9 2
17 1 9 2 16 15 9 13 0 9 2 13 0 0 0 9 9 2
21 9 13 0 1 0 9 13 0 7 0 9 2 1 15 15 15 13 0 0 9 2
20 9 1 0 9 4 1 9 1 11 11 1 9 9 13 9 3 13 1 11 2
11 10 0 7 0 9 4 13 9 11 11 2
16 13 4 0 9 0 9 7 9 0 9 2 1 0 0 9 2
12 0 9 13 2 16 1 10 9 13 9 9 2
13 1 0 13 9 2 16 4 1 11 13 10 9 2
12 9 13 9 9 2 7 13 13 9 0 9 2
26 1 0 9 9 0 9 1 9 1 9 13 9 9 9 7 9 2 16 4 3 13 14 9 10 9 2
43 0 13 9 14 1 0 9 2 0 9 9 2 2 1 11 2 1 11 2 11 2 1 11 2 11 2 1 11 2 0 9 2 2 0 11 7 11 2 3 0 9 2 2
18 9 13 0 14 1 0 7 0 9 2 1 9 7 9 7 1 9 2
22 9 0 9 2 16 13 0 9 2 13 0 9 0 9 2 16 15 13 1 0 9 2
22 1 0 9 13 9 3 0 2 3 13 0 9 1 9 2 16 11 13 14 1 3 2
9 7 13 9 7 9 9 9 0 2
23 3 0 9 1 12 9 13 0 13 2 4 13 11 11 2 9 1 9 1 9 1 11 2
37 9 1 9 12 2 16 15 4 13 9 9 11 2 4 13 13 14 9 12 2 16 4 1 0 9 13 0 7 0 9 0 9 1 0 12 9 2
23 9 9 1 9 12 4 13 13 2 16 4 13 0 0 0 9 2 15 13 1 9 9 2
32 0 0 9 2 16 13 9 0 9 2 13 9 1 10 0 9 9 2 13 15 4 0 9 2 16 13 9 0 2 0 9 2
31 14 1 10 9 4 13 1 9 9 0 9 2 16 0 9 3 7 3 13 2 1 0 9 9 7 9 13 0 0 9 2
23 0 9 11 2 16 4 9 9 13 9 8 1 11 2 15 4 0 0 9 13 9 12 2
32 9 1 9 2 9 7 9 2 9 1 9 2 0 9 9 7 9 1 9 1 9 4 9 1 0 9 12 13 13 9 12 2
11 0 9 15 4 13 1 3 0 0 9 2
14 0 0 9 7 9 0 9 4 13 1 0 0 9 2
11 1 15 3 13 0 9 0 9 9 11 2
15 16 15 14 4 13 2 14 4 13 14 3 0 9 9 2
26 12 15 13 9 1 0 9 7 10 9 2 0 9 1 0 9 2 10 0 2 0 0 7 0 9 2
23 9 2 16 4 13 0 1 0 9 2 14 15 13 9 7 9 7 0 9 7 0 9 2
15 9 12 9 12 4 1 9 0 9 13 0 9 9 9 2
17 3 14 3 1 0 9 13 10 9 1 0 9 0 15 0 9 2
8 7 15 13 9 2 9 2 2
16 14 13 7 13 0 1 7 1 9 2 0 2 0 9 2 2
30 13 15 2 16 14 13 1 12 2 1 10 9 0 9 9 0 9 2 16 4 13 1 0 0 9 3 0 7 0 2
12 0 13 0 9 1 9 9 1 10 9 9 2
10 9 0 9 11 13 3 0 1 9 2
19 13 4 7 15 4 1 0 9 13 1 0 9 1 9 7 1 10 9 2
47 9 1 9 9 4 13 14 9 9 1 0 0 9 11 2 16 1 0 9 2 16 15 7 10 9 13 1 9 9 7 9 0 9 2 13 3 0 9 2 7 14 9 9 7 0 9 2
22 1 10 9 9 13 0 9 9 11 7 0 9 1 11 1 0 9 1 11 9 12 2
21 13 0 9 10 9 2 1 15 4 11 7 0 9 1 11 13 1 9 9 11 2
9 14 15 1 15 14 13 13 0 2
17 1 15 9 13 9 11 7 9 9 1 11 1 9 9 9 11 2
24 9 1 9 15 1 0 9 1 9 13 2 7 15 13 14 9 2 16 15 9 13 0 9 2
18 9 15 13 13 9 7 9 14 1 3 0 9 2 16 3 13 0 2
10 1 9 0 9 13 0 13 10 9 2
19 9 13 1 9 3 9 16 9 2 7 13 9 2 16 15 13 2 3 2
37 1 0 9 7 9 15 9 3 13 1 9 0 9 7 9 2 1 9 10 9 7 1 9 2 1 9 1 0 2 9 2 9 2 9 7 9 2
8 1 9 9 0 9 13 0 2
6 9 9 1 9 13 2
16 3 16 13 9 3 0 1 0 9 7 9 2 3 4 13 2
22 1 11 13 14 0 1 15 2 16 13 13 7 13 1 15 2 16 13 14 3 0 2
12 15 13 14 0 9 1 15 2 15 14 13 2
37 3 7 13 2 16 13 0 13 2 16 13 9 3 1 9 15 2 16 15 13 14 0 9 1 0 9 2 16 15 2 16 15 13 9 0 9 2
34 7 16 13 0 9 3 0 9 2 13 13 15 14 3 0 9 9 2 7 14 13 14 2 16 4 1 10 9 13 2 14 2 0 2
40 0 9 4 1 9 2 0 2 2 2 0 2 2 0 9 11 11 7 9 1 9 0 9 13 0 9 9 2 16 15 13 1 0 9 2 1 9 0 9 2
37 0 9 2 16 15 1 10 9 1 0 9 13 1 0 9 2 1 0 9 1 9 1 0 9 9 2 16 15 13 0 9 3 2 13 3 0 2
52 0 9 2 0 9 2 3 13 1 0 9 0 9 0 0 9 1 9 0 1 9 0 9 2 16 1 0 0 9 1 0 0 9 13 1 10 9 2 16 4 1 9 2 9 7 9 9 9 13 14 0 2
35 9 4 13 1 9 0 9 2 9 0 0 9 2 16 4 13 0 9 2 15 4 3 13 0 9 2 1 9 7 0 9 0 0 9 2
16 1 15 7 1 15 4 15 3 3 13 0 3 0 9 9 2
15 7 15 13 1 0 9 9 11 2 11 2 11 2 11 2
28 16 13 14 1 15 2 16 4 13 9 2 3 1 9 0 9 2 9 1 0 9 9 2 3 4 13 3 2
30 12 9 1 12 9 2 1 15 4 13 12 9 2 4 13 0 9 11 2 16 13 1 9 14 3 2 3 1 9 2
17 7 9 13 14 1 10 0 9 1 10 9 2 16 7 4 13 2
37 3 2 16 4 15 13 1 10 10 9 1 11 2 4 13 14 9 1 9 11 2 16 4 13 3 9 2 16 15 10 9 1 9 13 12 9 2
21 13 4 10 9 7 10 9 4 13 2 16 4 13 0 9 11 2 16 15 13 2
9 1 10 9 4 15 14 14 13 2
24 9 4 13 1 9 1 0 2 1 11 7 4 13 9 2 16 4 10 0 9 13 7 13 2
42 16 3 9 13 9 9 1 0 9 2 16 4 9 13 2 16 13 10 0 9 2 7 3 9 13 0 7 3 0 9 9 9 2 16 13 0 9 1 0 0 9 2
21 16 1 10 9 13 0 9 2 15 3 13 2 3 9 3 13 14 10 0 9 2
10 7 7 13 14 0 9 7 0 9 2
21 9 11 4 3 13 0 9 2 16 4 13 2 15 13 0 1 9 9 1 9 2
11 9 14 4 13 9 0 9 7 14 9 2
8 1 15 14 4 13 0 9 2
25 1 0 9 7 9 15 3 13 2 16 4 11 13 15 1 0 0 9 7 7 4 13 14 3 2
21 7 14 1 9 15 3 11 13 1 9 7 9 1 11 13 1 9 1 0 9 2
13 7 4 13 0 0 9 9 16 0 9 0 9 2
28 16 13 9 1 9 9 2 16 15 13 2 7 9 2 16 15 13 0 9 2 0 2 13 10 9 14 0 2
12 7 7 2 3 0 9 13 7 13 9 9 2
20 11 11 7 11 11 11 2 16 14 3 13 9 0 9 2 9 3 13 3 2
12 7 10 9 13 1 3 0 9 0 0 9 2
27 0 9 13 14 2 3 15 4 11 3 13 13 0 9 2 15 4 3 13 3 13 9 9 1 0 9 2
4 9 13 0 2
17 1 0 9 4 13 0 0 9 0 0 9 2 16 13 3 0 2
15 3 7 15 4 1 10 9 9 13 9 9 1 0 9 2
10 0 4 3 1 0 9 3 3 13 2
21 3 7 13 3 0 9 0 14 1 15 2 16 4 1 9 9 13 9 1 9 2
7 9 9 9 14 13 0 2
7 9 13 3 0 9 9 2
12 0 9 15 13 7 1 15 13 0 0 9 2
13 14 3 13 7 13 2 3 4 13 10 10 9 2
15 9 4 0 13 13 1 10 0 9 2 1 11 2 11 2
13 13 4 16 9 7 4 1 9 13 3 10 9 2
22 16 4 13 2 16 15 0 9 14 13 1 9 2 4 15 3 13 10 0 0 9 2
25 1 9 9 1 0 9 4 9 12 9 13 0 9 1 8 8 2 8 8 7 8 8 1 11 2
28 1 15 4 13 7 13 12 9 9 9 2 9 9 2 12 9 9 2 12 9 9 7 0 9 1 12 9 2
22 1 8 8 7 8 8 4 13 0 9 1 9 9 0 9 0 9 7 9 1 9 2
6 1 10 0 9 13 2
13 7 9 13 10 9 2 16 3 13 1 10 9 2
15 7 15 13 9 10 9 2 16 13 2 3 13 1 15 2
4 15 13 9 2
3 4 13 2
10 13 7 15 2 16 14 13 14 0 2
8 13 7 3 10 9 1 9 2
10 14 12 7 12 4 13 1 10 9 2
17 16 16 4 9 14 13 9 13 9 7 9 10 9 1 12 9 2
50 0 11 2 1 11 15 1 0 9 13 3 12 9 2 3 9 15 7 15 13 1 9 0 2 0 9 2 16 13 1 9 9 0 0 2 0 9 0 14 1 9 0 9 7 9 9 1 9 9 2
22 1 0 0 9 9 4 9 13 2 16 4 3 13 3 0 9 14 1 0 0 9 2
19 16 13 9 1 0 9 2 13 9 10 9 3 13 7 15 13 0 9 2
47 2 3 1 15 2 16 4 1 9 7 0 9 9 0 9 3 13 2 4 13 0 9 1 9 3 0 2 2 15 4 13 9 9 2 16 4 13 1 9 13 9 1 9 0 12 9 2
20 3 4 1 15 13 9 9 1 9 9 2 1 15 4 13 9 3 1 0 9
26 11 11 1 9 1 9 15 4 13 2 16 9 13 9 9 1 11 2 13 14 1 9 1 11 11 2
17 15 10 9 13 9 2 1 15 15 3 13 9 1 0 0 9 2
21 2 9 1 9 1 9 7 15 14 13 1 0 7 0 9 2 2 4 14 13 2
31 9 0 7 3 0 9 2 16 15 11 13 1 10 9 2 3 14 13 0 0 9 2 1 15 4 13 14 0 0 9 2
30 1 10 9 13 0 0 0 9 0 7 0 9 9 2 10 9 1 0 9 1 0 0 9 7 9 0 9 0 9 2
18 14 7 13 0 0 9 1 0 9 7 9 2 16 13 3 9 9 2
21 15 13 9 0 9 7 9 9 0 9 9 7 0 9 0 9 1 15 1 9 2
22 1 11 4 3 13 11 2 16 15 4 13 15 14 0 9 1 12 2 0 9 9 2
21 0 9 3 1 9 2 16 4 3 13 9 2 4 3 13 7 0 4 13 9 2
20 2 1 15 13 12 9 0 9 7 3 13 2 16 13 3 0 9 1 0 2
18 11 4 3 14 13 12 9 2 13 7 4 14 1 0 9 1 12 2
25 9 12 4 0 9 11 3 1 11 11 2 16 14 3 13 0 0 9 2 13 0 9 0 11 2
24 1 9 4 9 13 14 1 10 9 0 7 0 9 1 0 9 2 16 4 13 14 0 9 2
19 3 3 4 15 11 13 1 0 9 1 11 7 11 7 13 0 0 9 2
23 1 9 0 9 4 13 14 0 9 11 11 2 11 7 11 11 2 11 11 7 11 11 2
20 9 0 15 13 1 15 2 16 4 0 0 9 1 0 13 1 9 7 9 2
28 11 0 9 1 0 0 9 4 0 9 13 0 9 9 7 9 2 3 1 0 9 13 3 3 3 7 3 2
21 3 13 1 9 9 9 11 2 16 13 10 14 0 0 9 1 0 1 0 9 2
21 0 9 15 13 3 3 2 13 7 4 1 9 0 13 15 7 9 1 10 9 2
39 1 0 9 9 0 7 9 2 0 0 9 2 1 9 2 0 9 7 0 9 7 0 0 7 0 9 13 9 1 10 9 13 14 10 9 16 0 9 2
40 11 11 1 11 13 2 16 4 0 9 1 0 3 3 7 3 13 9 9 1 0 9 2 10 9 7 4 13 0 11 2 16 15 13 9 9 3 1 9 2
7 1 10 9 13 9 0 2
3 2 8 2
34 3 9 3 14 13 14 9 1 9 9 2 4 15 0 9 13 13 14 9 0 9 2 9 9 1 0 9 11 7 4 13 9 9 2
15 13 4 0 0 9 11 11 1 0 9 1 0 9 11 2
21 11 4 13 9 1 10 9 1 0 9 1 10 9 2 16 4 13 1 9 11 2
24 0 9 1 9 2 12 9 0 7 0 9 13 1 9 12 9 2 15 13 1 9 7 9 2
18 12 0 9 13 2 13 7 13 1 0 9 7 1 15 13 9 9 2
8 9 13 7 15 13 1 9 2
24 1 9 3 13 0 9 2 13 12 0 9 2 12 0 9 2 9 9 7 10 9 0 9 2
14 16 15 3 13 2 13 9 7 15 13 0 12 9 2
25 0 9 13 1 9 2 1 15 13 0 9 7 13 1 9 2 16 15 3 13 1 9 7 9 2
19 0 9 0 9 1 11 4 13 0 9 12 1 9 9 1 11 1 11 2
15 9 11 11 11 4 13 9 12 1 0 0 9 10 9 2
12 9 11 11 4 13 1 10 0 9 0 9 2
24 3 4 13 1 9 9 2 15 13 0 9 7 1 9 0 9 13 9 1 9 7 1 15 2
10 0 9 14 13 1 15 12 0 9 2
22 0 0 7 0 9 7 14 15 13 0 9 1 9 9 2 16 15 13 16 0 9 2
32 0 9 11 11 4 14 9 3 1 0 9 14 13 2 3 4 15 0 9 11 3 2 1 0 0 11 2 13 1 0 9 2
17 0 9 4 14 13 1 0 9 2 7 13 1 9 1 8 11 2
20 3 4 1 9 7 0 9 3 13 9 0 9 2 9 0 9 7 0 9 2
18 1 0 9 4 3 1 0 0 9 13 11 2 16 4 13 0 9 2
16 7 15 13 14 0 9 2 1 15 4 15 13 15 15 0 2
30 1 0 9 9 9 3 13 9 9 7 10 9 1 0 2 3 0 7 0 9 2 16 13 15 0 1 9 7 9 2
11 1 15 13 0 7 3 13 14 0 9 2
16 13 9 2 16 4 13 1 9 7 4 1 15 13 1 9 2
19 1 9 15 4 13 2 15 15 13 13 7 3 1 15 3 13 2 2 2
11 7 15 4 1 10 9 13 14 1 9 2
15 1 9 9 13 9 9 2 16 13 1 10 9 0 9 2
3 9 13 2
15 11 11 13 9 2 16 15 3 13 1 9 9 7 9 2
15 0 11 13 7 9 11 11 2 12 1 0 9 1 9 2
34 16 15 0 9 13 13 9 0 9 2 13 2 16 13 3 3 0 1 0 9 0 9 9 2 16 15 1 0 9 13 1 0 9 2
13 9 3 1 9 9 13 2 16 9 13 12 0 9
28 1 9 1 0 9 15 3 13 1 0 9 2 1 9 1 9 7 9 1 9 7 9 14 15 4 3 13 2
14 16 13 2 7 13 14 1 11 14 3 9 1 9 2
20 10 10 0 9 2 9 1 12 13 14 14 3 12 9 2 13 1 15 14 2
23 1 9 2 9 7 9 3 13 9 12 9 9 2 16 15 4 13 2 16 9 3 13 2
9 0 0 9 1 10 14 0 9 2
24 9 15 0 9 4 3 13 2 16 15 14 13 2 16 13 9 1 9 9 2 9 7 9 2
28 1 9 9 2 9 9 1 9 1 0 9 7 11 11 9 13 3 14 9 0 9 9 1 0 9 7 9 2
9 3 0 7 13 9 9 1 9 2
32 1 0 7 13 0 14 9 2 16 15 9 13 7 1 15 9 13 3 13 2 15 15 3 13 7 10 9 15 15 13 0 2
17 14 13 14 9 9 2 15 9 1 9 13 2 16 13 2 2 2
30 0 7 0 13 1 9 1 15 3 0 7 0 9 7 13 9 1 0 9 1 9 2 16 4 3 11 13 0 9 2
29 11 11 2 2 0 9 11 1 9 12 2 12 15 4 3 13 2 0 13 0 9 1 9 12 2 12 2 2 2
9 2 1 9 14 4 13 9 9 2
32 0 9 2 10 9 2 16 13 9 1 0 9 2 4 3 13 2 16 4 13 0 9 9 12 3 3 0 9 1 0 9 2
47 3 1 3 1 11 4 13 1 3 0 0 9 2 0 9 1 10 0 9 7 0 9 2 7 14 1 11 15 4 1 9 9 13 2 14 2 12 0 9 2 1 15 4 13 0 9 2
20 1 0 9 3 13 9 2 1 9 0 9 1 9 9 13 13 15 0 9 2
8 0 9 13 0 9 1 9 2
33 13 14 0 9 11 3 2 16 4 13 3 3 0 2 7 1 0 0 9 2 16 4 13 1 9 9 2 4 15 15 13 13 2
29 9 0 1 9 4 3 13 9 11 11 2 11 2 2 1 15 4 1 12 0 9 13 9 9 9 1 0 9 2
20 9 4 14 1 9 13 9 1 9 11 11 2 16 14 3 13 1 9 11 2
24 16 13 9 0 2 4 13 3 3 3 13 0 9 16 7 1 9 3 1 0 13 9 1 9
17 9 3 13 1 9 0 9 2 1 15 13 0 9 14 9 9 2
7 7 15 3 1 15 13 2
3 13 3 2
26 9 13 0 1 0 9 0 9 2 0 9 7 9 9 9 2 16 4 13 1 9 1 10 16 9 2
12 9 13 2 16 15 13 0 7 7 14 0 2
28 3 13 0 2 16 3 10 9 2 16 15 13 1 0 9 2 13 1 10 0 9 2 16 16 15 13 0 2
4 15 13 9 2
9 0 7 0 9 13 10 9 0 2
10 14 3 3 9 9 13 1 9 3 2
5 2 13 10 9 2
8 15 14 13 2 15 13 9 2
11 1 9 0 0 9 4 13 14 12 9 2
22 13 15 1 9 1 9 7 9 2 1 15 4 13 9 2 13 1 0 7 0 9 2
23 3 13 0 9 12 1 0 9 2 16 13 9 7 9 10 9 7 9 2 16 15 13 2
8 14 15 13 13 0 0 9 2
13 0 13 2 16 13 12 1 12 0 9 1 9 2
16 14 13 2 16 4 3 3 13 7 14 9 3 15 4 13 2
33 9 2 9 9 1 0 9 13 1 15 2 16 4 3 1 0 9 7 0 9 13 9 3 7 15 13 2 15 15 1 9 13 2
15 7 3 3 4 13 14 15 2 15 15 3 13 7 13 2
16 16 13 3 2 16 15 15 14 4 13 2 7 3 4 13 2
33 7 16 4 15 13 13 1 9 2 16 13 0 9 9 1 9 7 0 9 1 9 1 9 2 3 13 15 0 14 13 0 9 2
8 7 15 13 1 9 1 9 2
31 2 13 0 9 1 9 2 7 16 13 10 9 14 3 0 3 2 9 2 16 4 13 1 9 2 7 13 14 3 0 2
19 9 4 14 3 13 9 1 9 7 3 4 13 1 9 2 13 15 4 2
10 0 9 4 15 13 2 9 4 13 2
22 9 13 1 10 0 7 0 9 2 9 1 0 9 2 9 2 9 7 9 0 9 2
10 13 15 14 1 10 0 9 1 9 2
10 1 10 9 13 0 14 1 0 9 2
25 1 9 0 9 14 3 13 9 1 9 11 11 2 16 4 13 1 9 1 11 0 9 11 11 2
19 2 16 4 13 12 0 9 2 4 15 3 13 13 1 11 2 2 13 2
11 0 9 2 1 9 15 13 3 13 9 2
7 14 3 13 9 13 3 2
38 16 13 3 1 10 7 15 9 2 3 13 2 3 13 1 9 15 15 2 15 4 3 13 1 0 9 9 7 9 2 16 13 15 0 1 9 9 2
14 16 13 9 12 0 9 2 3 13 9 3 14 0 2
11 1 0 9 13 3 14 0 7 0 9 2
12 13 15 12 9 2 16 4 13 1 15 0 2
24 7 15 4 13 1 9 7 3 4 1 10 9 13 1 9 2 16 13 3 15 13 13 9 2
20 15 4 1 9 13 9 7 4 13 2 3 4 13 3 2 15 13 7 13 2
8 13 4 0 9 7 15 13 2
18 13 4 3 9 2 1 3 15 14 13 13 7 3 13 3 9 13 2
8 10 9 13 2 16 15 13 2
21 3 7 13 1 15 3 13 7 14 13 2 16 15 15 13 1 9 7 0 9 2
31 16 13 3 2 15 13 14 9 2 16 14 4 13 9 2 9 2 9 2 1 15 9 3 13 7 15 3 7 3 13 2
18 11 13 0 9 1 0 9 1 11 2 16 13 1 9 9 1 15 2
20 3 13 14 3 9 3 13 9 1 15 2 16 4 13 13 9 1 0 9 2
18 10 0 9 13 2 14 13 15 15 13 7 1 9 15 10 9 13 2
17 1 0 9 2 9 2 9 2 9 7 9 13 0 1 9 9 2
23 1 0 9 9 7 9 15 13 1 3 0 2 3 13 1 10 9 13 9 1 10 9 2
15 1 9 13 14 3 0 9 2 16 9 0 14 14 13 2
6 13 15 14 1 0 2
10 1 0 9 15 13 14 3 9 9 2
14 9 0 9 2 10 9 7 9 0 0 9 1 0 9
27 9 4 1 12 9 9 13 9 9 1 9 9 7 9 9 2 16 14 4 13 0 9 8 8 0 9 2
21 0 9 1 9 9 14 4 13 9 0 0 9 7 9 10 9 1 0 0 9 2
20 1 9 1 9 9 13 9 13 9 7 13 9 1 9 9 2 0 1 9 2
36 1 9 0 9 1 9 4 1 9 0 9 11 11 13 9 10 0 9 2 1 15 9 9 1 9 9 9 1 9 0 9 14 4 13 14 2
5 2 10 9 13 2
29 0 0 9 11 11 2 16 13 1 9 9 1 0 9 2 4 1 0 9 13 12 3 0 9 1 3 12 0 2
24 16 13 9 3 2 7 13 9 1 0 0 9 2 7 11 13 10 9 1 9 12 12 9 2
18 1 9 11 13 9 9 2 0 9 9 2 9 9 7 0 0 9 2
15 9 9 13 3 0 1 9 0 9 7 14 1 9 9 2
29 12 9 1 0 9 2 16 15 13 1 9 9 1 9 2 13 9 2 16 4 10 9 3 13 1 10 9 11 2
16 7 15 14 3 14 13 2 16 1 10 9 3 11 3 13 2
32 1 11 4 13 1 10 9 14 1 9 11 2 1 15 13 14 3 3 13 0 9 2 16 4 9 10 9 13 0 0 9 2
40 9 1 9 11 0 1 15 14 13 3 0 2 7 0 9 1 9 1 10 0 9 1 10 9 2 14 2 13 9 2 1 15 4 3 3 1 9 13 11 2
38 9 13 14 15 2 16 13 9 1 10 9 3 10 9 2 1 15 13 3 13 14 14 9 0 0 2 0 9 2 16 15 3 1 0 13 3 9 2
4 9 13 0 2
41 16 1 9 13 2 16 13 0 9 1 9 0 9 0 2 16 0 14 14 13 13 2 7 13 1 9 1 9 1 9 0 9 2 9 9 7 14 13 13 3 2
20 9 1 0 0 9 15 4 14 13 9 2 7 1 3 13 10 9 1 9 2
40 3 0 9 2 16 9 9 13 1 0 9 0 9 2 1 9 1 15 2 16 13 14 9 2 0 1 9 2 7 15 15 14 14 13 14 0 1 15 0 2
45 7 3 16 4 9 13 1 0 9 9 7 0 9 2 1 15 15 4 14 3 1 9 16 9 13 9 1 0 9 2 4 15 1 9 13 15 15 2 16 4 15 13 1 11 2
10 10 0 0 9 15 4 13 1 15 2
20 11 4 13 0 9 0 9 2 1 15 13 11 13 7 2 13 2 0 9 2
7 14 11 4 1 9 13 9
9 2 11 14 4 13 14 0 9 2
12 9 13 0 9 2 9 9 9 1 0 9 2
14 1 0 9 15 13 10 9 7 1 15 13 9 9 2
12 10 0 9 1 11 0 0 9 13 1 9 2
12 9 13 1 0 9 1 0 0 9 1 9 2
20 3 13 0 9 9 9 2 3 1 0 9 9 2 16 13 0 9 0 9 2
19 1 9 4 13 10 9 16 3 3 7 14 9 0 4 13 14 3 0 2
17 9 1 9 4 13 2 13 4 3 12 9 3 1 0 0 9 2
20 7 4 13 3 0 1 9 2 7 0 0 9 4 14 13 0 1 0 9 2
17 13 15 2 16 4 15 0 0 9 1 11 13 1 9 0 9 2
16 9 4 13 0 7 0 7 11 4 13 1 0 2 0 9 2
12 7 15 1 15 15 4 13 2 16 4 13 2
7 14 0 4 13 3 0 2
35 9 9 2 16 4 13 1 9 0 12 9 2 7 15 4 3 7 3 3 13 1 9 2 16 4 13 2 0 2 2 0 7 0 9 2
6 14 3 4 15 13 2
16 15 14 13 7 15 13 14 0 13 0 7 15 13 1 0 2
6 7 4 15 3 13 2
12 3 4 3 13 1 0 9 0 9 1 15 2
12 13 4 2 16 15 4 0 9 7 3 13 2
12 13 4 7 15 13 2 3 14 13 10 9 2
33 1 11 13 15 0 2 9 9 2 0 1 9 0 9 7 9 2 0 9 2 14 1 12 9 0 0 9 13 3 14 1 3 2
11 0 0 9 1 0 9 13 1 0 9 2
11 9 2 14 16 15 13 2 13 1 9 2
13 9 9 2 16 13 1 9 0 2 13 3 0 2
15 7 16 13 0 9 0 9 2 1 15 9 13 0 9 2
10 9 0 9 14 1 9 13 0 9 2
19 1 0 11 15 4 9 13 2 16 15 13 2 15 13 0 9 0 9 2
15 11 4 13 13 2 14 13 4 9 2 16 15 4 13 2
15 11 4 13 3 0 9 2 1 15 15 15 4 13 13 2
16 13 4 15 13 7 13 15 2 15 9 1 11 14 13 13 2
5 0 9 13 0 2
8 1 11 15 4 13 1 11 2
23 11 11 13 9 1 9 0 9 1 0 9 2 16 14 4 15 13 9 0 9 11 11 2
10 9 10 9 4 13 0 9 1 0 2
31 1 10 9 4 3 11 11 13 1 0 9 1 9 1 11 7 1 9 11 1 0 9 0 9 7 1 9 1 0 9 2
28 9 9 11 11 4 13 2 16 13 9 1 9 9 2 7 13 2 16 4 9 9 1 9 7 0 9 13 2
28 9 3 13 13 1 9 1 11 7 1 10 9 4 14 13 10 9 9 7 9 2 15 1 3 4 13 3 2
16 1 3 13 9 0 9 1 9 9 9 2 13 9 1 11 2
20 9 9 13 1 10 0 9 9 2 16 13 10 9 1 9 0 2 13 9 2
3 2 8 2
14 3 4 3 11 13 3 2 16 4 9 13 14 11 2
16 7 9 0 9 11 7 11 1 11 4 13 0 9 0 9 2
19 15 3 14 4 13 2 16 4 0 0 9 13 1 14 3 0 9 9 2
23 9 9 1 0 9 3 1 9 12 9 13 1 9 2 9 2 9 2 9 7 9 9 2
9 10 0 9 13 1 10 9 9 2
9 0 0 9 13 14 9 7 9 2
11 14 9 9 13 2 10 13 10 0 9 2
22 1 0 9 4 15 13 9 10 0 9 1 0 9 7 0 9 1 0 7 0 9 2
4 13 7 13 2
10 1 15 4 13 3 14 3 0 11 2
11 13 15 14 9 0 9 7 0 0 9 2
25 7 4 13 1 15 0 2 16 15 14 4 4 9 14 3 13 2 7 16 15 3 14 13 14 2
14 0 9 0 9 13 9 1 12 0 0 9 1 9 2
45 16 0 9 11 7 11 13 3 0 0 9 2 14 4 13 9 11 2 16 15 13 3 1 12 9 3 2 16 13 9 1 9 9 11 2 9 12 1 12 9 0 16 1 9 2
18 0 1 9 0 9 7 13 9 12 9 2 16 13 1 0 0 9 2
10 9 4 13 13 1 9 1 0 9 2
19 9 2 16 13 3 0 9 2 16 13 0 7 0 9 2 13 13 3 2
4 9 13 3 2
18 1 9 1 9 7 15 13 13 2 16 9 13 7 7 15 13 0 2
17 14 3 13 1 10 9 1 9 13 14 1 0 9 0 9 9 2
25 1 9 9 9 3 0 9 13 1 12 1 12 9 1 9 12 1 12 9 7 0 9 12 9 2
30 1 9 13 3 0 2 16 0 9 13 1 0 9 2 16 9 14 13 13 9 2 7 3 0 9 13 0 1 9 2
41 11 13 1 9 0 0 9 3 0 1 9 9 1 9 11 2 7 15 3 3 13 2 16 13 14 1 0 13 9 11 2 16 1 15 3 4 13 10 0 9 2
29 14 4 15 15 1 3 13 11 11 7 11 11 2 16 3 13 1 11 2 0 9 7 14 3 3 13 1 11 2
26 1 0 9 0 9 14 4 15 1 0 9 9 8 0 9 1 11 13 13 14 1 0 9 9 12 2
33 16 13 0 9 2 13 0 9 9 8 8 9 2 0 1 9 0 0 9 7 9 1 9 2 1 15 13 0 0 9 1 9 2
21 1 10 9 7 1 9 0 9 9 13 0 9 2 16 4 13 9 1 0 9 2
16 1 9 9 13 1 9 12 9 9 2 16 13 14 0 9 2
13 1 3 9 13 0 1 0 9 9 2 9 2 2
11 9 2 16 15 13 2 4 13 0 9 2
16 0 13 3 9 11 1 0 9 2 1 15 13 15 3 3 2
14 0 0 9 15 13 1 9 7 9 7 13 0 9 2
13 0 7 0 4 3 13 9 2 16 4 15 13 2
16 2 3 7 14 13 15 2 2 15 15 4 1 9 13 11 2
19 1 9 9 11 0 9 11 11 13 0 12 0 0 9 0 9 2 2 2
12 1 12 9 7 9 9 0 9 13 0 9 2
26 9 0 9 13 1 0 9 1 0 9 2 1 0 9 7 1 9 2 16 13 1 9 9 0 9 2
20 1 10 9 13 0 9 9 0 9 1 0 9 7 9 9 9 1 10 9 2
20 1 10 9 13 9 9 1 9 2 10 0 9 13 3 0 1 0 0 9 2
11 1 0 9 1 9 13 9 1 0 9 2
29 10 10 9 2 16 13 1 12 9 12 3 0 1 11 2 13 13 14 0 9 2 16 13 3 0 9 1 0 2
22 9 9 2 16 4 13 0 1 12 9 12 2 13 3 1 9 0 9 1 0 9 2
26 1 15 2 3 13 9 2 9 7 9 2 15 3 13 7 10 9 13 0 1 9 2 4 14 13 2
17 1 0 9 4 13 1 9 9 2 9 9 7 9 9 7 9 2
18 2 3 0 1 0 9 13 9 0 9 7 9 9 7 0 9 9 2
12 7 13 0 2 16 13 9 1 0 9 9 2
21 9 1 9 13 13 0 2 7 15 13 1 9 9 7 7 9 1 9 3 13 2
37 14 7 13 2 16 4 13 15 15 2 16 4 13 10 9 2 16 15 13 9 2 0 1 0 9 7 9 2 16 15 13 3 2 16 13 9 2
15 0 9 13 0 3 3 13 2 16 3 3 13 9 9 2
22 9 4 14 3 13 0 9 1 0 9 2 0 7 13 13 9 0 9 1 0 9 2
35 2 10 0 0 9 15 4 13 13 1 0 9 2 16 15 13 11 7 16 13 3 0 7 3 0 2 2 4 13 11 11 1 9 11 2
38 16 4 13 1 0 9 1 9 2 4 11 2 16 4 13 1 10 9 14 3 2 1 9 14 1 0 12 9 1 12 9 13 0 9 0 9 9 2
19 1 10 9 2 1 15 4 3 13 2 4 3 13 1 10 9 7 9 2
13 7 13 4 0 2 1 15 7 15 4 13 9 2
6 11 4 13 3 3 2
12 13 4 15 13 9 2 16 4 13 15 0 2
15 7 4 15 14 13 1 0 9 2 14 16 4 3 13 2
9 1 9 3 13 9 1 10 9 2
16 2 16 13 0 9 2 9 2 9 2 0 9 7 0 9 2
8 9 14 13 2 7 15 13 2
7 9 15 13 1 0 9 2
26 13 7 1 9 13 9 1 9 9 2 16 4 3 13 2 15 4 3 13 2 7 13 9 14 3 2
16 9 13 3 7 13 1 9 2 16 9 1 15 14 4 13 2
19 1 9 13 0 9 1 9 2 7 7 15 13 1 0 9 7 0 9 2
4 13 12 9 2
6 0 13 1 0 9 2
23 1 0 11 13 1 9 0 1 0 9 14 9 9 2 1 9 1 9 2 9 7 9 2
6 15 1 10 9 13 2
21 13 13 2 16 15 4 13 3 15 2 15 4 13 2 16 4 15 14 13 9 2
5 9 13 0 13 2
13 13 15 0 13 7 13 2 14 13 7 3 13 2
12 13 13 2 16 15 4 13 0 7 0 9 2
20 0 4 13 1 0 9 9 3 1 0 0 9 2 0 9 7 10 9 13 2
24 9 4 13 2 16 15 4 0 9 13 1 9 1 0 9 7 3 15 4 13 13 9 9 2
12 3 15 13 16 9 2 0 1 12 0 9 2
14 1 9 15 13 9 2 16 15 13 13 7 13 0 2
18 0 9 13 0 1 0 2 0 13 15 1 9 1 12 7 12 9 2
14 16 15 13 0 2 13 9 2 16 13 14 10 9 2
14 3 3 13 10 9 9 1 10 9 1 9 10 9 2
12 1 10 9 13 9 2 9 7 0 0 9 2
25 1 10 9 7 9 2 16 15 3 13 1 9 2 9 14 13 9 1 9 2 16 13 1 9 2
18 10 0 9 3 13 2 11 13 12 9 2 0 1 10 9 7 9 2
26 9 14 13 2 3 3 13 2 16 13 1 10 9 2 7 9 2 1 9 2 1 15 15 14 13 2
16 0 9 13 0 7 0 2 9 7 1 9 13 14 10 9 2
17 9 13 14 0 7 0 9 2 13 14 0 0 9 1 9 9 2
19 16 13 2 16 13 9 10 9 0 7 0 2 13 14 12 0 0 9 2
18 1 9 13 9 2 3 15 13 7 9 13 1 9 2 9 7 9 2
27 0 9 9 13 1 0 9 7 9 13 13 12 9 2 3 7 15 13 1 9 7 9 13 1 0 9 2
10 13 2 13 0 1 15 7 10 9 2
11 1 0 9 14 13 7 9 7 9 9 2
20 14 3 13 0 9 2 15 9 13 13 2 10 9 13 1 10 9 0 9 2
25 9 9 13 9 2 1 15 13 9 7 9 7 13 1 9 2 16 3 13 15 2 15 15 13 2
21 16 4 13 9 2 4 3 13 9 1 9 2 16 13 15 0 2 0 2 0 2
14 14 0 9 3 13 1 0 9 2 9 7 9 9 2
9 1 9 13 14 9 1 0 9 2
15 3 0 9 1 9 13 9 9 2 16 15 13 1 9 2
20 13 3 9 2 16 15 13 9 2 15 7 13 0 9 9 2 9 7 9 2
24 3 15 9 9 13 1 0 9 2 16 13 0 2 0 2 0 7 3 3 14 13 1 9 2
17 9 15 3 1 0 9 2 16 15 13 2 13 14 1 0 9 2
18 9 1 9 3 13 0 2 16 7 13 9 0 2 9 15 13 9 2
6 0 9 2 13 0 2
8 14 13 9 2 16 13 9 2
4 13 0 9 2
7 13 9 9 1 0 9 2
39 13 9 13 9 1 9 9 1 9 2 15 13 2 16 13 9 9 1 9 2 3 13 9 9 7 9 9 2 16 13 14 2 15 7 9 9 3 0 2
8 9 13 2 15 13 1 9 2
26 1 0 9 13 12 1 12 9 9 7 1 15 1 0 9 13 9 2 0 9 7 1 9 0 9 2
9 2 9 13 2 13 7 15 13 2
6 14 3 13 14 9 2
16 2 0 9 15 13 0 13 14 2 16 1 0 9 13 9 2
24 9 2 16 4 13 9 2 13 7 15 14 13 14 1 0 9 2 16 15 3 13 1 9 2
8 1 10 9 13 0 13 9 2
13 14 0 9 13 2 16 9 13 2 9 7 13 2
28 1 0 9 9 2 3 0 9 0 9 7 12 7 12 9 1 0 9 7 1 0 9 0 9 9 3 13 2
26 13 9 0 9 2 16 13 9 7 9 9 1 0 9 2 1 15 13 9 0 2 0 7 0 9 2
13 16 9 13 1 0 9 2 15 13 1 0 9 2
12 0 9 9 2 0 9 7 9 2 9 9 2
26 0 9 4 13 2 16 1 10 0 9 0 9 13 3 9 9 1 9 1 9 9 7 9 1 9 2
7 3 4 15 13 7 13 2
30 0 13 2 16 4 13 15 3 0 9 2 16 4 3 13 2 16 4 15 1 10 9 13 2 1 0 9 1 11 2
5 7 10 9 13 2
3 9 0 2
55 4 7 1 9 1 9 10 9 13 1 14 0 9 2 16 4 13 1 9 9 2 16 13 0 9 9 7 16 1 9 13 9 9 10 9 1 9 2 15 13 0 9 1 0 9 2 1 15 14 4 15 10 9 13 2
4 7 13 3 2
53 15 15 4 7 3 13 7 4 3 14 3 13 2 16 4 13 1 11 2 4 13 15 2 16 15 4 0 9 13 2 16 14 13 9 2 16 13 3 9 10 9 2 16 15 9 13 1 0 9 7 1 9 2
25 14 2 14 2 15 13 0 2 15 13 0 7 14 10 9 3 3 7 0 9 15 13 1 9 2
10 3 4 15 13 2 3 15 14 13 2
4 15 14 13 2
6 0 9 2 0 9 2
19 14 10 9 4 13 1 9 2 7 13 3 0 2 16 16 4 13 9 2
16 13 13 14 15 2 16 4 1 0 0 9 13 1 0 9 2
10 1 15 4 13 13 3 9 9 12 2
10 1 10 9 13 0 13 1 0 9 2
12 0 9 4 14 13 2 16 13 9 1 9 2
35 15 9 13 3 1 12 9 9 7 14 9 0 9 7 9 9 13 2 16 4 15 10 9 13 1 0 1 12 9 1 3 12 9 9 2
10 0 9 4 14 13 10 9 1 9 2
12 1 10 9 13 0 0 9 9 1 11 11 2
3 9 9 2
8 15 4 13 13 1 10 9 2
6 3 1 15 4 13 2
5 13 14 0 9 2
5 15 13 10 9 2
10 13 4 2 16 13 14 0 12 9 2
17 13 4 2 16 4 0 0 9 1 11 13 9 7 4 13 9 2
42 16 9 10 0 9 7 16 10 9 10 9 13 2 10 0 9 4 13 1 0 9 7 0 9 2 16 4 13 10 9 1 9 2 16 4 0 9 15 10 9 13 2
19 16 13 2 13 3 1 10 9 7 4 13 1 0 9 2 16 15 13 2
6 7 3 4 13 9 2
32 13 10 9 2 3 4 13 2 3 14 4 13 9 1 10 0 9 9 7 15 3 3 7 3 13 2 3 13 10 9 0 2
23 16 7 15 14 13 2 14 15 13 10 9 10 9 2 16 13 15 9 7 16 9 13 2
15 3 4 3 15 0 13 1 9 1 0 9 2 11 2 2
17 9 1 2 14 2 0 0 9 7 0 9 7 0 9 13 0 9
4 15 15 13 2
14 16 15 13 11 7 16 13 0 2 4 1 9 13 2
19 0 9 13 2 16 4 0 9 11 13 0 9 9 2 16 13 0 9 2
29 1 12 9 13 1 11 0 9 9 9 2 11 7 4 10 9 9 13 16 0 9 1 9 9 1 9 0 9 2
38 11 2 3 16 4 0 9 1 0 9 1 0 0 0 9 1 11 0 9 9 13 9 7 9 2 4 13 0 9 9 1 11 0 14 0 0 9 2
30 1 11 11 1 11 2 0 0 9 2 15 4 1 0 9 1 9 9 11 11 1 0 9 1 9 9 13 11 11 2
28 0 0 9 15 3 13 1 9 2 16 15 14 13 13 2 9 15 1 0 7 0 9 3 13 1 0 9 2
8 7 9 9 14 13 16 9 2
24 13 1 9 2 16 13 0 9 2 1 9 15 14 4 13 1 0 9 7 3 0 0 9 2
10 3 13 1 0 9 0 9 7 9 2
10 3 13 1 9 13 9 0 9 9 2
9 7 16 13 3 2 10 9 13 2
18 0 9 1 9 7 4 3 16 1 12 9 14 3 13 9 0 9 2
53 9 9 4 14 13 3 2 16 0 0 9 14 9 9 14 4 13 0 14 1 0 2 9 2 2 16 0 9 13 0 9 9 1 11 2 7 3 1 9 2 2 15 4 3 3 13 9 11 1 9 1 9 2
41 7 0 16 1 0 0 9 1 9 2 16 15 1 9 4 13 14 1 0 9 1 10 0 9 2 7 4 14 13 9 11 2 1 0 9 14 3 4 13 15 2
27 1 11 4 3 13 9 0 9 2 16 14 4 15 13 14 1 9 0 9 2 7 4 3 13 9 9 2
16 3 4 15 13 0 9 2 16 1 0 9 13 14 3 0 2
21 1 12 9 4 11 13 9 1 0 9 1 0 0 0 7 0 9 2 11 2 2
32 7 3 1 12 9 15 4 13 2 16 11 4 13 1 0 9 2 2 0 9 2 4 13 2 9 2 1 0 9 1 11 2
46 9 9 2 16 15 14 3 3 13 0 9 0 9 2 9 9 9 7 9 1 9 2 7 10 0 9 3 13 14 3 2 16 15 4 0 9 9 1 0 14 3 13 10 0 9 2
13 11 11 4 1 0 9 13 3 16 9 0 9 2
22 1 9 0 9 4 11 1 0 12 7 12 9 13 1 9 10 9 14 12 9 9 2
10 1 15 4 13 14 0 9 11 11 2
14 16 4 3 13 1 9 2 15 4 13 10 0 9 2
16 1 0 9 13 10 9 2 16 4 13 1 15 3 0 9 2
17 14 3 3 1 0 9 13 10 9 9 1 10 9 1 0 9 2
25 10 0 9 13 1 0 0 9 1 9 3 10 16 12 9 7 13 3 12 0 9 10 0 9 2
24 15 4 3 13 9 2 1 0 9 7 9 2 16 15 4 13 2 7 4 15 15 3 13 2
44 16 14 3 13 14 1 9 9 2 4 13 2 16 14 4 13 0 2 0 0 9 2 1 15 4 15 9 13 7 14 1 12 9 13 10 9 1 0 9 2 15 9 13 2
12 1 9 4 14 13 0 9 2 0 1 9 2
14 13 4 15 1 0 9 0 9 2 16 13 3 0 2
19 9 4 1 0 13 3 1 9 1 0 9 7 0 9 1 9 0 9 2
19 0 9 4 13 3 1 9 2 9 1 9 7 13 1 0 9 3 0 2
11 1 10 9 13 3 0 14 0 9 9 2
11 9 0 9 4 14 13 1 0 9 9 2
19 9 15 4 3 13 1 0 9 2 16 0 9 15 4 13 1 0 9 2
9 1 0 9 4 9 9 13 3 2
24 16 4 3 13 10 9 1 9 2 4 3 13 1 0 9 2 7 15 3 13 9 1 9 2
21 3 4 13 10 9 2 16 15 13 2 1 12 2 12 9 7 15 3 13 9 2
15 4 15 15 1 9 9 1 0 9 9 13 1 3 7 3
19 11 1 9 1 9 14 14 13 13 10 9 2 3 14 13 7 13 15 2
45 7 4 15 3 3 13 0 9 11 2 1 10 9 0 7 0 11 11 11 2 16 4 1 0 9 13 2 16 11 13 0 9 1 9 11 2 1 15 4 9 13 1 0 9 2
10 16 4 13 2 4 15 13 16 9 2
54 9 9 2 16 13 0 0 0 2 0 9 2 4 13 14 0 2 16 4 3 13 1 3 0 11 2 11 7 15 4 14 13 2 16 4 13 1 0 9 9 1 11 2 16 4 11 3 3 13 9 11 2 11 2
48 13 4 14 2 16 4 15 13 14 0 9 1 9 11 11 7 0 9 1 9 11 11 2 7 4 13 3 0 9 2 16 4 15 13 2 16 4 13 3 1 3 0 9 0 9 1 11 2
3 2 8 2
12 11 11 13 9 2 0 9 0 0 9 11 2
17 1 10 9 11 13 2 16 3 1 12 9 15 14 13 1 9 2
20 16 4 13 9 2 4 13 14 12 9 13 1 11 7 13 0 9 1 11 2
9 10 10 9 13 1 9 11 11 2
20 9 1 11 4 3 13 0 9 2 0 9 2 13 0 9 7 9 7 9 2
31 0 9 7 0 2 0 9 2 2 16 15 13 7 4 13 1 9 14 0 2 13 1 0 9 11 1 0 9 0 9 2
14 1 11 15 4 13 0 9 7 14 3 13 7 13 2
54 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 7 0 9 3 13 0 7 0 9 2
46 1 0 0 9 2 16 13 14 3 13 0 9 7 9 14 13 1 9 11 0 9 7 13 9 2 16 1 11 13 0 9 11 2 7 13 2 16 4 3 13 0 7 3 0 11 2
9 7 15 13 13 0 9 0 9 2
13 9 2 16 15 4 13 2 14 4 13 12 9 2
22 1 9 9 4 15 1 9 11 13 1 0 9 2 16 4 13 14 3 3 0 9 2
35 11 11 4 15 9 13 16 9 7 0 9 3 2 11 11 7 13 14 2 3 15 13 13 3 2 1 15 2 16 3 13 1 9 11 2
20 14 0 3 13 2 16 13 9 1 2 3 0 2 9 7 0 9 15 0 2
12 0 9 11 4 1 9 11 3 13 14 0 9
21 9 4 9 13 9 3 2 16 4 13 14 1 9 2 7 15 4 13 10 9 2
11 9 14 4 13 2 16 4 13 3 0 2
26 7 15 4 13 3 2 16 4 9 13 1 0 0 9 9 2 1 0 9 7 4 13 9 13 9 2
16 9 15 4 3 13 1 0 9 2 9 7 4 14 13 9 2
20 10 9 13 9 9 2 16 4 0 9 13 1 11 7 3 13 13 0 9 2
15 9 10 12 9 4 13 0 0 9 11 11 7 11 11 2
24 13 15 4 14 2 16 4 10 9 13 1 0 9 2 16 4 13 10 9 1 0 9 11 2
19 0 0 7 0 9 4 15 3 13 7 1 9 9 11 13 3 1 9 2
26 0 9 4 13 0 14 1 0 9 2 16 4 13 9 10 16 12 9 7 14 4 13 9 0 9 2
15 3 1 9 1 11 4 15 0 9 13 13 1 0 9 2
28 0 9 0 9 11 11 4 13 0 9 2 0 0 9 11 11 7 4 13 2 16 4 3 13 1 0 9 2
17 0 0 9 2 1 9 2 4 3 13 1 9 9 9 1 11 2
5 9 4 13 0 2
12 9 2 9 7 9 4 13 0 1 0 9 2
13 9 4 13 2 1 0 9 4 15 13 0 9 2
13 11 4 13 1 0 9 2 7 3 4 13 11 2
15 1 0 9 1 9 7 9 9 1 11 4 13 14 12 9
14 11 11 15 14 13 1 11 2 16 13 10 9 1 11
16 1 9 4 3 13 7 13 3 0 2 16 13 9 0 9 2
6 13 4 3 1 9 2
13 1 0 9 4 11 13 2 3 0 13 1 9 2
15 1 10 9 13 9 9 9 0 14 1 15 2 3 13 2
29 10 9 15 13 13 14 1 9 1 9 2 16 15 4 13 0 9 2 16 14 13 1 0 9 2 9 9 2 2
28 1 0 9 13 0 14 0 9 3 1 0 9 0 9 2 16 9 9 13 1 9 2 0 1 9 1 9 2
9 3 0 9 3 3 13 1 9 2
12 1 0 9 3 1 9 13 14 10 0 9 2
17 9 13 3 0 14 3 2 16 15 1 0 9 7 9 14 13 2
25 10 9 9 2 3 2 13 3 13 1 9 14 1 9 9 2 7 15 14 3 13 9 0 9 2
19 0 9 13 9 1 0 9 1 0 9 2 1 15 13 0 9 0 9 2
13 10 9 13 3 3 3 1 9 7 3 1 9 2
20 0 9 15 4 3 13 1 0 7 1 9 0 9 7 1 3 0 0 9 2
23 16 13 3 0 9 2 15 13 0 13 1 0 9 1 0 9 2 16 13 10 10 9 2
24 9 1 10 0 9 3 13 10 9 2 3 7 13 15 0 2 16 9 9 13 10 0 9 2
25 16 13 0 9 0 14 1 0 9 2 13 14 3 0 9 2 16 7 15 13 3 13 1 3 2
19 9 0 9 0 0 9 13 3 0 2 1 15 7 3 13 3 0 9 2
28 10 9 13 3 7 3 7 13 0 9 0 2 3 0 7 0 9 2 16 15 3 13 1 3 0 0 9 2
28 1 0 15 9 13 3 0 1 9 0 9 2 16 3 2 16 15 14 13 2 13 9 2 8 1 0 9 2
18 0 9 13 0 1 9 9 7 1 3 0 16 14 1 3 0 9 2
11 3 15 13 7 13 1 9 0 0 9 2
17 14 13 15 7 0 7 0 9 2 10 9 7 13 13 3 0 2
10 9 13 3 13 2 16 13 0 9 2
21 3 13 9 10 9 9 2 9 7 9 1 0 9 2 16 1 15 13 0 9 2
10 10 9 4 3 1 9 13 0 9 2
20 1 9 0 9 4 9 13 9 1 0 9 9 0 9 7 0 9 0 9 2
31 0 9 9 0 9 13 1 15 2 16 9 0 9 4 13 10 0 9 7 15 4 13 1 9 2 16 15 13 1 9 2
33 9 4 3 3 13 2 16 4 0 9 1 9 13 14 9 12 7 16 4 1 9 12 1 9 9 12 13 15 1 10 0 9 2
38 16 4 9 13 10 0 9 2 4 13 1 0 9 2 3 7 4 13 9 7 10 9 2 16 1 10 9 13 2 16 4 13 0 2 3 14 13 2
33 0 9 4 13 2 16 4 9 13 1 10 9 3 12 9 2 16 1 0 9 13 2 16 4 3 13 14 1 12 1 12 9 2
21 9 4 13 2 16 10 9 2 16 15 13 9 2 1 12 9 4 13 0 13 2
18 1 15 15 13 9 2 3 4 3 9 3 13 9 7 14 13 9 2
21 9 0 9 4 1 9 13 9 1 9 9 1 9 1 0 9 7 13 0 9 2
14 3 4 13 9 1 9 7 13 0 9 9 0 9 2
26 14 3 7 3 4 13 2 16 4 9 3 13 2 1 0 9 1 9 7 4 15 13 9 2 2 2
12 1 9 4 13 2 16 13 11 3 0 9 2
29 1 0 4 13 9 2 16 4 1 9 2 16 4 13 1 11 2 16 15 3 13 2 0 9 13 12 9 9 2
19 14 1 9 7 4 13 2 16 15 4 1 11 13 14 9 8 11 11 2
11 3 10 9 13 2 16 13 9 14 9 2
38 2 10 9 13 2 16 15 13 2 16 15 4 1 0 9 3 13 2 2 13 11 11 2 0 1 9 2 9 7 9 1 9 9 11 1 11 11 2
15 0 9 15 4 3 3 13 3 1 9 13 9 1 9 2
24 16 4 13 2 15 1 10 9 13 2 16 4 1 9 12 13 9 9 0 9 1 12 9 2
11 7 14 4 13 1 9 16 1 9 9 2
6 9 4 13 9 13 2
8 14 7 13 9 13 0 9 2
14 7 9 15 4 13 9 0 1 9 0 9 1 11 2
21 2 6 2 2 4 13 2 16 4 13 11 1 9 1 9 7 15 13 1 9 2
24 16 4 15 9 13 1 10 0 9 2 4 9 14 13 2 7 1 15 3 4 13 15 13 2
6 14 9 4 13 3 2
9 7 16 15 13 12 9 1 9 2
12 9 15 4 13 1 9 1 9 7 13 13 2
7 14 14 3 13 1 9 2
7 9 14 4 13 15 0 2
36 9 1 0 13 3 13 2 16 4 1 9 1 9 2 16 13 1 15 0 7 0 2 13 14 10 9 7 9 7 10 0 0 7 0 9 2
22 14 4 1 15 3 13 2 1 15 13 2 16 4 3 15 13 2 15 9 4 13 2
15 3 1 9 0 9 4 9 3 13 9 1 0 9 9 2
44 1 12 9 9 2 16 15 4 13 3 1 9 11 11 2 4 3 13 9 2 0 0 9 2 16 3 13 2 16 4 13 11 11 7 1 9 0 9 13 14 0 0 9 2
36 7 14 3 13 2 16 4 1 9 11 3 13 1 0 9 1 0 9 2 16 15 10 0 9 1 10 0 9 2 1 0 9 2 3 13 2
34 0 9 1 9 13 0 2 0 9 1 3 0 11 11 12 11 7 14 13 2 16 13 3 10 9 1 0 9 9 3 16 1 9 2
17 10 9 13 7 1 9 1 9 0 9 2 16 15 15 13 0 2
44 10 9 1 9 2 16 13 1 15 1 9 2 13 1 10 9 3 13 10 0 9 2 16 7 13 1 9 2 1 15 15 14 13 3 2 9 13 9 2 16 13 15 0 2
16 15 3 1 9 9 13 1 9 7 13 10 0 9 7 9 2
21 9 1 9 0 9 13 14 0 9 2 16 4 15 9 13 9 2 7 0 9 2
9 9 0 9 3 13 14 1 9 2
16 1 9 4 13 14 0 9 2 16 1 9 1 9 3 13 2
21 14 9 7 9 1 9 9 1 9 13 14 9 9 2 16 10 9 13 1 0 2
35 11 10 12 9 0 9 15 4 3 13 1 10 0 0 9 1 0 9 1 9 9 2 16 4 15 1 9 13 1 0 9 1 0 9 2
14 13 4 10 9 2 7 14 4 13 9 1 15 0 2
23 7 1 10 9 4 13 9 2 7 4 15 9 9 2 1 15 4 15 13 2 13 9 2
20 11 11 7 11 11 13 9 0 0 9 1 9 1 9 1 11 0 11 11 2
33 1 10 9 4 13 2 16 4 0 9 11 11 1 0 0 9 13 1 9 7 15 4 16 9 0 9 13 1 0 9 0 9 2
24 0 9 4 3 1 9 11 11 1 9 11 13 9 2 1 15 4 13 12 9 0 0 9 2
3 2 8 2
17 14 1 10 9 4 13 13 0 9 1 9 9 1 9 7 9 2
9 15 13 9 1 0 9 0 9 2
14 7 4 3 3 3 2 16 4 13 2 13 0 9 2
18 16 13 11 11 1 11 2 4 14 1 0 0 9 11 13 0 9 2
15 15 4 7 9 0 9 1 9 0 0 9 3 14 13 2
10 1 0 9 4 0 9 13 16 0 2
17 1 15 7 4 14 11 13 2 16 15 4 13 1 0 9 9 2
12 3 13 0 9 2 16 4 3 13 3 9 2
7 9 11 4 13 1 9 2
7 13 4 12 7 12 9 2
4 9 4 13 2
23 13 15 4 13 9 1 3 14 0 0 9 2 16 7 15 4 1 9 13 1 9 9 2
7 2 9 0 9 3 13 2
14 9 9 7 9 13 14 1 0 9 7 9 3 0 2
12 1 11 13 1 14 9 10 9 12 0 9 2
13 9 13 15 2 16 4 13 1 9 3 3 3 2
31 14 16 15 4 1 0 9 13 0 9 0 9 2 16 4 9 13 3 1 9 2 4 13 2 15 4 13 3 1 15 2
10 0 9 1 11 15 13 1 0 9 9
11 1 9 7 9 0 9 13 0 0 9 2
3 13 0 2
4 15 7 13 2
8 3 13 0 2 4 15 13 2
16 4 13 3 0 1 9 2 4 14 3 13 7 3 13 9 2
36 1 9 2 3 15 4 3 14 13 1 9 13 9 2 4 13 2 16 3 9 13 14 0 9 9 7 9 2 14 13 7 13 1 0 9 2
11 15 4 3 13 14 9 1 9 0 9 2
12 15 3 13 2 16 4 9 9 13 1 9 2
40 1 12 9 4 15 9 13 10 10 9 2 3 7 4 13 0 9 2 16 4 13 3 16 10 9 14 3 3 13 2 15 15 13 1 0 9 1 0 9 2
17 1 10 0 0 9 4 9 13 1 0 9 2 9 13 0 13 2
16 15 4 13 0 9 1 3 0 9 7 9 9 1 0 9 2
29 9 10 0 9 13 9 8 11 11 2 16 15 4 13 9 12 0 9 0 9 2 16 13 3 1 0 0 9 2
10 3 15 4 1 15 13 9 2 2 2
53 13 4 3 0 9 11 11 2 16 13 9 9 13 11 11 2 9 10 0 9 1 11 2 16 15 4 1 10 9 1 0 9 13 14 1 9 0 9 11 1 11 2 2 16 13 1 0 9 13 1 11 2 2
27 10 9 7 3 0 9 2 9 7 9 10 9 4 13 11 9 2 16 0 9 13 1 9 0 9 9 2
17 11 2 1 0 9 1 11 13 3 1 12 9 9 1 9 9 2
18 1 0 9 4 9 7 9 13 9 9 2 16 4 15 13 10 9 2
32 9 9 15 4 13 1 0 7 0 9 2 9 0 9 7 15 4 1 9 9 3 13 10 0 9 7 9 7 13 0 11 2
8 1 9 4 9 13 0 9 2
11 1 9 4 13 9 9 7 0 13 9 2
20 9 14 13 2 1 15 13 14 0 9 7 12 9 1 9 7 3 0 9 2
28 16 4 13 10 9 0 1 3 0 9 1 9 2 15 4 3 1 0 9 3 13 9 14 1 9 1 9 2
30 2 1 9 1 9 13 1 9 9 12 13 0 9 9 2 13 0 9 1 9 0 9 7 15 13 1 12 1 12 2
15 3 13 3 13 2 16 13 1 3 0 0 7 0 9 2
30 1 15 13 13 2 16 9 1 0 9 14 4 13 10 9 1 0 9 11 2 2 4 13 9 9 11 11 11 11 2
27 9 0 7 0 9 4 15 7 13 2 16 4 13 0 9 7 16 1 0 0 9 14 0 9 14 13 2
28 1 9 1 9 7 9 4 15 13 2 16 0 9 2 16 13 0 1 9 2 13 10 9 1 0 9 11 2
11 11 4 1 0 9 9 13 1 0 11 2
31 9 9 11 11 7 9 11 11 4 3 1 9 1 11 1 9 13 1 11 2 16 15 4 1 3 13 9 0 9 11 2
18 0 9 2 16 13 14 12 9 2 13 0 2 16 16 4 13 12 9
13 9 10 9 2 1 9 15 10 9 4 14 13 2
35 2 3 1 15 2 16 4 9 14 3 13 3 1 9 1 9 2 15 13 2 3 4 13 0 2 16 15 14 13 3 7 13 0 9 2
16 1 9 13 0 14 12 0 9 2 16 15 4 13 11 11 2
7 9 13 0 9 1 9 2
9 9 9 1 9 13 9 0 9 2
11 1 11 4 15 9 13 1 11 7 11 2
28 1 0 9 4 9 13 1 9 10 9 2 15 0 2 1 9 0 9 2 13 7 15 15 4 3 12 9 2
41 3 15 4 13 1 9 11 2 16 4 1 0 9 1 12 9 7 1 9 0 9 1 9 9 13 9 9 1 11 2 16 0 9 14 13 1 9 9 0 9 2
13 11 9 11 11 11 4 3 13 0 9 0 9 2
32 16 13 1 0 13 0 9 1 11 2 0 9 7 11 2 15 3 9 2 16 15 4 13 1 12 9 2 13 1 12 9 2
3 2 8 2
22 11 4 1 9 13 9 11 2 16 4 1 9 12 2 12 13 1 9 9 0 9 2
18 3 14 0 9 4 13 2 16 15 3 2 9 2 3 13 3 3 2
29 1 15 4 10 9 9 13 2 7 3 16 3 2 9 7 4 13 0 2 9 2 2 15 9 4 13 0 9 2
19 9 0 9 7 10 9 13 1 15 9 0 9 1 9 9 1 0 9 2
15 0 9 13 1 9 9 1 0 9 9 2 0 1 9 2
35 0 13 2 16 1 12 7 0 0 9 0 9 13 0 2 0 9 2 16 13 9 9 1 9 10 9 7 0 9 1 9 7 9 9 2
23 0 9 1 9 1 10 0 2 9 2 13 14 0 9 9 1 9 2 7 14 10 9 2
18 9 1 9 9 7 13 10 9 7 1 0 13 9 1 3 12 9 2
20 0 9 13 1 9 0 0 9 0 9 2 1 9 7 4 13 3 0 9 2
30 1 9 9 0 9 4 13 14 15 1 9 9 1 15 2 1 15 14 4 13 0 9 2 7 14 3 0 16 9 2
14 1 9 15 4 9 14 0 13 2 15 9 13 13 2
15 15 13 2 16 4 15 13 15 15 0 13 14 1 9 2
19 15 4 13 3 0 1 11 2 7 15 13 3 15 2 16 13 1 9 2
21 1 0 9 7 14 13 13 2 16 4 13 15 0 7 7 16 4 13 15 0 2
23 10 9 13 2 16 4 15 9 13 3 13 1 9 9 2 1 15 4 13 1 9 9 2
13 9 4 15 13 13 1 9 9 1 0 0 9 2
24 9 4 3 13 3 1 15 2 16 4 11 9 13 14 16 0 9 2 7 16 0 0 9 2
21 1 0 9 15 4 9 13 3 1 0 9 2 15 15 15 13 1 10 9 0 2
29 16 9 3 13 9 3 3 2 16 15 13 2 14 16 15 1 9 9 13 9 2 15 13 2 16 9 4 13 2
16 3 16 1 9 11 11 13 14 1 0 0 9 3 0 9 2
38 1 0 9 11 4 1 9 9 1 9 1 11 11 11 10 0 9 13 0 1 9 11 11 2 16 15 4 13 15 3 0 0 9 8 12 1 9 2
11 1 0 9 4 13 0 9 12 9 9 2
14 1 15 14 13 14 9 2 16 9 14 14 13 9 2
4 3 13 0 2
20 0 9 7 14 13 2 7 9 4 1 0 9 13 14 3 12 2 0 9 2
22 11 4 1 9 13 2 16 13 1 10 9 1 12 1 12 9 0 9 1 9 9 2
26 14 13 2 1 15 15 13 15 2 16 13 2 16 15 9 3 13 1 9 2 3 7 13 10 9 2
17 14 11 11 13 14 12 9 11 2 7 13 10 9 1 11 9 2
21 11 4 13 0 9 2 16 4 15 2 16 4 13 9 2 3 13 9 1 9 2
11 0 9 9 14 4 13 1 9 0 9 2
30 9 14 4 1 10 9 13 3 1 9 2 9 1 9 7 14 4 13 1 9 3 12 2 0 9 14 3 0 9 2
13 9 14 14 4 13 3 13 9 1 0 0 9 2
35 13 9 9 9 1 9 0 9 7 9 2 9 2 9 7 9 9 9 2 16 13 3 0 0 9 1 9 1 12 1 12 9 0 9 2
25 10 9 13 9 1 9 9 2 16 15 1 9 12 13 1 9 11 7 13 1 9 1 9 11 2
31 1 0 9 2 16 15 13 1 9 11 7 13 1 9 1 9 11 1 9 1 9 12 2 15 13 0 9 2 3 2 2
38 1 0 7 0 9 2 16 13 0 1 9 1 12 1 12 2 15 1 9 1 9 11 13 9 1 0 0 9 14 1 9 0 9 0 1 10 9 2
7 0 0 9 15 14 13 2
36 9 2 16 13 9 1 9 2 13 13 0 2 1 0 9 7 0 9 9 0 8 1 9 9 0 7 1 9 1 9 0 9 1 9 9 2
20 1 0 9 3 13 1 0 7 0 9 0 9 7 9 1 0 14 0 9 2
31 0 9 1 15 13 13 7 14 13 9 2 7 13 0 2 16 4 9 13 15 7 2 13 2 0 9 1 9 7 9 2
22 14 3 13 0 0 9 0 1 9 2 16 15 13 13 1 9 1 12 7 12 9 2
11 9 13 9 9 1 9 7 9 0 9 2
13 1 9 9 7 4 14 3 13 14 9 1 11 2
13 14 13 2 3 0 9 13 1 0 9 10 9 2
16 15 13 14 9 0 9 2 16 15 9 9 13 1 0 9 2
20 13 13 14 12 2 0 9 2 7 15 4 9 1 12 9 9 13 1 9 2
27 1 9 9 7 9 9 9 10 9 0 9 7 13 10 9 2 16 4 15 13 1 9 9 12 1 9 2
27 0 9 13 3 0 9 2 1 15 15 0 3 13 9 2 7 15 13 9 1 15 9 14 13 3 13 2
14 3 15 13 1 0 9 9 2 16 13 0 9 9 2
17 1 15 4 15 3 13 9 9 2 7 3 13 14 1 0 9 2
17 0 9 4 13 3 2 0 9 9 9 13 0 9 1 0 9 2
35 15 1 9 9 1 10 9 13 9 1 9 1 0 9 1 9 2 16 13 0 9 1 9 9 2 9 7 9 9 2 16 15 13 15 2
