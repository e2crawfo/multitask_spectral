68495 11
6 11 2 9 1 9 2
1 9
2 11 11
47 16 12 1 12 0 9 1 0 11 2 9 0 9 11 11 2 1 11 13 9 1 0 9 12 0 9 7 9 10 9 3 13 16 9 0 9 2 13 15 3 1 9 13 1 0 9 2
7 9 2 13 3 0 9 2
31 7 3 2 9 7 9 3 0 2 9 12 0 9 1 0 9 1 11 2 15 13 0 9 0 9 13 7 13 1 9 2
18 1 0 0 9 1 9 11 13 13 2 16 15 15 3 13 16 13 2
47 1 15 2 16 4 13 2 16 15 1 11 2 0 1 9 9 11 2 1 0 9 9 13 3 0 2 13 9 12 9 9 2 16 4 15 3 13 2 16 14 2 7 3 15 15 13 2
24 0 2 3 0 9 2 16 4 11 1 9 13 13 14 12 9 1 9 2 13 3 1 9 2
24 1 9 11 11 2 16 4 11 7 11 13 3 13 1 9 2 9 11 13 2 11 3 13 2
26 0 13 2 16 9 1 9 9 2 16 13 11 3 1 11 13 2 13 10 0 9 2 15 13 9 2
32 9 1 15 2 16 11 13 11 1 11 9 7 9 2 3 7 0 2 7 0 2 13 1 0 9 13 0 9 12 2 9 2
11 1 10 0 9 1 11 13 2 13 9 2
21 13 0 13 9 1 9 9 2 16 4 13 0 9 1 9 0 9 1 9 9 2
11 0 9 2 0 9 2 13 3 0 9 2
2 0 9
2 11 11
9 9 0 9 15 14 13 0 9 2
8 4 15 3 13 9 0 9 2
26 15 13 9 2 13 15 2 16 9 0 13 3 9 9 2 1 15 13 2 3 13 11 11 2 0 2
13 9 0 0 9 2 1 10 0 9 13 10 9 2
9 3 13 0 9 7 9 0 9 2
7 1 0 9 13 15 9 2
33 1 15 1 0 9 15 13 1 15 2 16 9 13 9 7 9 13 3 1 15 2 16 4 9 13 7 10 9 13 1 0 9 2
10 0 9 10 9 0 9 1 15 13 2
57 0 9 13 3 1 9 0 2 13 15 10 0 0 9 1 10 0 9 7 13 9 1 10 9 2 16 9 13 0 9 2 3 13 7 13 9 2 16 0 9 13 0 1 10 0 7 0 9 2 15 4 1 9 10 9 13 2
12 9 1 9 13 0 9 7 9 15 3 13 2
21 13 0 9 13 15 2 16 12 9 0 9 13 15 0 2 16 12 9 0 9 2
66 16 7 12 9 0 9 1 9 9 0 2 15 13 12 9 0 9 2 7 0 0 9 1 9 13 2 13 15 9 9 15 12 9 0 1 9 1 10 15 0 9 7 1 10 9 15 13 9 3 15 1 15 2 1 0 0 9 2 15 13 3 0 1 0 9 2
14 14 2 16 4 13 15 15 2 15 13 13 10 9 2
12 7 9 13 3 15 2 15 15 3 3 13 2
26 10 0 0 3 7 13 13 7 3 15 13 1 9 0 9 7 15 3 10 9 13 1 10 0 9 2
13 3 15 13 9 7 10 9 7 13 3 9 0 2
11 0 9 0 4 13 3 1 9 3 13 2
26 13 15 1 0 0 9 15 13 3 3 2 16 13 9 2 16 4 9 2 1 15 15 13 2 13 2
5 0 9 7 13 2
26 13 15 1 0 0 9 0 2 0 7 0 9 2 15 13 3 7 3 10 9 13 2 3 7 13 2
23 0 9 13 3 3 0 9 0 9 7 0 9 2 15 3 1 10 9 13 0 9 0 2
14 13 15 1 9 0 3 3 2 3 3 15 13 9 2
10 13 12 12 9 13 1 15 10 9 2
13 13 1 3 0 0 9 0 9 13 14 0 9 2
4 3 2 7 3
1 9
2 11 11
25 9 9 11 11 1 9 13 2 16 3 1 1 10 9 13 10 9 13 1 9 9 2 14 9 2
12 7 16 3 10 0 9 13 13 1 0 9 2
15 1 9 0 9 15 9 13 1 0 9 3 2 7 3 2
20 0 9 9 11 11 13 14 1 9 2 3 15 1 0 9 13 3 13 9 2
18 1 15 7 2 15 13 1 0 9 0 7 0 9 3 0 9 0 2
20 0 9 13 1 0 9 1 9 2 3 1 9 13 0 9 11 2 3 3 2
18 1 9 2 9 7 9 13 9 2 0 9 2 9 9 7 0 9 2
18 3 15 9 11 13 0 2 3 13 7 1 10 9 1 9 9 13 2
6 13 2 16 9 13 2
20 7 16 1 10 9 2 14 3 1 0 9 0 0 7 0 9 2 13 13 2
18 0 9 2 15 9 3 1 9 0 9 13 2 13 1 10 9 3 2
48 9 9 0 0 9 2 9 9 9 1 0 9 7 3 9 9 1 9 0 0 9 2 13 15 2 16 11 11 3 13 13 0 0 9 9 9 9 2 7 13 13 3 0 9 3 0 9 2
31 13 2 16 0 0 9 15 13 7 1 15 2 16 1 0 9 13 9 9 9 7 13 9 1 0 9 1 9 0 9 2
9 16 4 13 14 15 3 2 2 2
2 0 9
1 9
2 11 11
13 1 9 13 9 9 9 1 9 0 0 0 9 2
83 10 9 2 1 9 2 16 15 1 15 7 13 7 9 2 13 0 0 9 3 0 9 2 9 2 9 7 9 4 13 1 9 2 15 15 15 13 2 1 9 10 9 15 13 0 9 2 13 15 10 0 9 2 4 13 7 13 0 2 0 2 0 7 0 9 2 1 0 9 13 3 13 1 9 9 7 0 9 1 0 9 9 2
14 3 0 2 1 0 9 15 13 9 1 9 0 9 2
22 1 15 3 13 9 2 1 15 10 9 1 9 13 2 0 9 9 15 13 7 9 2
12 3 3 13 9 1 9 7 9 9 10 9 2
19 1 9 1 0 9 1 9 9 1 9 9 13 12 10 9 9 0 9 2
45 11 11 3 3 13 2 16 9 9 9 13 1 0 16 10 9 7 9 2 10 9 7 13 1 9 9 1 0 7 3 3 0 9 9 7 0 9 15 1 9 7 9 0 9 2
30 0 15 7 13 13 9 2 3 9 9 13 3 9 2 15 13 0 9 0 13 1 10 7 15 9 0 3 0 9 2
26 0 0 9 15 7 13 2 1 15 0 13 1 9 10 9 16 9 9 2 3 4 13 10 0 9 2
14 9 0 9 7 13 3 9 9 9 7 9 10 9 2
15 0 9 13 9 2 16 9 9 7 10 9 15 13 3 2
47 1 10 9 13 3 0 9 9 1 9 0 9 1 0 9 0 2 9 13 9 2 10 9 13 3 1 9 2 7 14 1 9 10 9 15 3 2 13 0 9 11 1 9 12 9 2 2
23 1 15 2 16 0 9 4 13 13 9 9 9 7 0 9 0 0 9 2 13 3 15 2
17 9 10 9 3 13 9 2 1 9 9 7 10 9 13 13 3 2
8 9 15 3 4 13 1 9 2
24 1 10 9 7 13 9 9 11 2 16 4 15 3 3 9 15 1 0 9 13 1 12 9 2
5 0 9 1 0 9
4 11 2 11 2
31 9 0 0 9 0 9 1 0 9 11 3 13 2 16 0 9 1 9 15 13 3 3 2 16 3 13 13 10 0 9 2
25 9 0 9 11 1 9 13 9 2 16 7 0 9 13 0 13 9 9 0 9 7 9 12 9 2
25 11 13 0 9 11 11 2 11 11 2 16 4 11 13 0 9 2 15 4 13 9 1 0 9 2
4 11 11 3 0
2 11 2
30 0 9 0 9 0 9 11 2 0 9 2 11 2 2 13 9 11 11 2 15 1 0 0 9 13 3 3 1 9 2
17 10 0 9 13 9 0 9 11 11 3 0 3 2 3 0 2 2
21 12 1 9 13 9 1 11 2 11 1 9 2 3 9 11 13 2 13 1 11 2
17 1 9 15 7 13 10 0 9 1 11 7 10 0 9 11 11 2
22 11 2 15 15 3 13 0 9 1 0 9 2 3 13 13 1 9 9 1 0 9 2
22 11 13 9 2 16 1 12 9 13 0 9 0 9 2 16 4 13 9 1 0 9 2
5 0 9 13 1 11
2 11 2
30 0 0 9 2 0 0 9 9 11 7 0 9 9 11 2 11 2 13 3 1 11 1 9 1 0 9 11 2 11 2
23 3 13 9 1 11 1 0 11 1 9 1 11 2 11 2 9 11 11 2 0 9 11 2
10 0 9 1 0 11 10 9 3 13 2
41 13 15 1 9 11 1 0 0 9 7 13 9 2 16 15 13 1 9 0 7 0 9 3 1 9 2 3 15 13 13 3 0 2 16 11 13 9 10 0 9 2
25 11 7 0 9 1 0 9 3 13 2 16 13 0 10 9 1 0 9 2 16 11 13 0 9 2
15 9 11 11 12 2 13 3 1 9 11 1 9 0 9 2
11 9 0 12 9 13 9 0 9 0 11 2
15 11 11 12 2 1 9 13 9 9 1 10 9 1 11 2
2 9 11
3 9 0 9
5 13 13 0 11 2
4 9 1 9 2
5 3 13 9 11 2
4 13 11 9 2
16 2 10 7 15 0 9 15 10 9 13 1 0 7 0 9 2
16 9 9 15 13 9 0 11 1 11 2 9 0 0 0 9 2
17 3 0 9 1 10 0 0 9 13 3 14 9 9 1 0 9 2
16 0 9 7 13 1 3 16 12 9 0 9 9 2 11 11 2
9 2 11 2 2 11 12 2 12 2
5 11 2 0 9 9
2 11 2
22 1 11 13 3 16 12 9 1 0 9 0 9 1 9 11 1 9 11 1 9 9 2
16 13 15 3 9 0 0 0 9 1 0 9 11 2 11 2 2
44 1 9 13 3 9 2 16 15 0 9 13 13 7 9 13 9 1 0 9 0 9 2 13 9 0 2 0 9 1 9 0 9 1 11 2 15 4 13 1 0 0 9 11 2
5 9 13 9 12 11
3 0 11 2
19 0 9 1 0 0 9 1 9 12 1 11 13 9 0 9 11 0 11 2
20 13 15 0 9 2 15 13 0 9 9 2 15 13 1 0 7 0 0 9 2
11 0 9 15 13 1 3 0 9 0 9 2
17 9 3 13 13 2 3 15 13 10 9 7 3 9 13 0 9 2
20 9 11 11 13 2 16 3 10 9 3 0 9 13 0 13 16 9 1 9 2
14 13 2 16 4 10 0 9 4 1 9 13 0 9 2
18 1 0 9 15 9 13 1 0 9 9 14 1 0 11 1 0 9 2
11 10 9 7 13 7 3 0 0 0 9 2
4 11 13 9 9
4 11 2 11 2
25 11 13 1 0 9 2 16 4 13 1 0 9 2 7 13 2 16 0 11 15 13 1 10 9 2
34 1 0 9 13 0 9 0 11 10 9 11 11 11 1 9 1 9 0 0 9 7 0 12 9 2 7 10 0 9 13 1 0 9 2
20 0 0 9 3 13 2 16 9 13 1 0 0 0 9 2 9 0 0 11 2
23 0 0 9 4 3 13 9 0 11 7 10 9 0 9 1 0 2 0 9 1 9 11 2
12 13 15 0 9 2 15 15 13 1 10 9 2
2 0 9
21 1 0 9 13 0 0 9 2 15 15 13 0 9 2 12 0 7 12 0 9 2
37 3 3 13 0 9 2 9 2 16 15 0 9 2 1 10 9 0 9 7 10 9 0 9 2 13 9 0 9 9 2 13 1 9 9 1 12 2
9 16 15 13 2 13 3 1 9 2
43 1 9 9 13 2 13 0 9 2 0 11 11 7 13 2 7 1 9 4 13 2 16 11 13 0 9 7 0 9 16 15 2 16 10 9 11 13 0 7 0 16 11 2
4 11 13 9 11
2 11 2
31 11 3 13 0 9 0 9 11 11 1 9 9 1 0 9 1 12 9 1 9 9 1 9 7 9 1 11 2 11 2 2
36 9 0 9 9 13 2 16 11 13 13 14 1 0 9 7 1 9 2 16 11 13 9 1 12 0 11 7 16 4 13 9 0 9 1 9 2
20 11 1 0 11 3 13 1 0 2 0 9 1 11 1 9 0 9 11 11 2
17 0 2 0 9 15 3 13 0 9 2 1 9 9 1 0 11 2
8 0 3 13 1 0 0 9 2
5 12 9 13 1 11
2 11 2
32 1 11 4 1 0 12 9 2 3 9 1 9 0 9 1 9 2 13 1 0 9 0 7 0 9 1 12 9 0 0 9 2
31 0 9 2 15 3 13 1 11 2 1 15 7 0 9 9 11 2 11 2 4 13 13 0 9 1 11 1 9 1 9 2
15 13 7 3 9 13 9 2 16 9 4 13 1 9 9 2
38 11 4 13 1 0 7 0 9 2 11 3 13 9 1 11 2 3 1 9 0 9 9 1 9 2 7 7 1 9 13 9 1 9 0 9 1 11 2
5 0 9 9 14 9
2 11 11
14 13 2 16 4 13 0 13 15 3 2 13 11 11 2
16 11 13 0 9 1 10 9 2 13 15 0 9 9 11 11 2
16 12 10 9 15 13 3 0 9 9 9 9 0 9 11 11 2
27 12 9 13 3 1 0 9 0 2 0 2 16 9 1 0 9 2 13 16 9 11 1 0 9 0 9 2
34 0 13 10 2 0 2 9 0 9 2 15 15 3 1 9 13 2 7 9 1 15 13 2 7 13 1 15 2 15 0 2 0 9 2
12 9 1 9 13 3 3 3 7 3 13 9 2
18 12 0 13 2 3 2 0 0 9 7 3 16 4 15 3 3 13 2
40 12 13 7 3 9 9 7 3 13 3 0 10 9 13 2 0 9 13 7 1 0 9 3 0 2 16 15 13 13 0 9 7 3 15 1 10 0 9 13 2
8 15 13 7 1 9 9 9 2
35 1 0 9 12 0 9 0 15 9 10 2 15 11 1 9 13 2 7 2 0 0 9 2 0 9 7 9 1 12 9 13 0 9 3 2
13 0 9 3 4 1 0 9 13 1 9 9 3 2
26 1 0 2 7 3 3 0 9 13 2 2 9 3 3 0 0 9 2 16 0 9 1 9 0 9 2
29 2 9 0 0 9 2 15 13 0 9 0 9 2 7 16 0 2 0 9 10 9 1 9 2 3 15 9 13 2
16 2 9 0 9 0 0 9 1 3 3 0 9 2 1 9 2
8 9 0 9 1 0 9 9 2
18 2 3 0 9 1 0 9 0 7 0 9 2 15 3 13 9 9 2
16 2 9 12 9 9 1 9 1 9 0 9 0 9 9 9 2
24 1 3 0 13 0 13 9 9 2 9 7 9 2 15 13 13 9 2 3 10 9 3 13 2
30 1 10 9 4 13 2 16 3 3 13 3 1 0 9 2 7 3 3 2 7 16 0 9 3 3 3 13 9 2 2
21 1 0 9 1 0 9 9 3 11 13 2 16 13 9 9 9 1 0 0 9 2
7 13 15 15 2 7 15 2
5 3 3 1 15 2
21 10 0 9 2 10 0 9 15 0 9 3 3 13 2 13 1 0 9 1 9 2
20 1 9 10 0 2 10 0 9 15 3 3 3 13 2 15 3 13 9 9 2
11 9 3 13 2 16 15 0 13 3 3 2
25 9 2 15 15 13 13 1 9 2 7 3 3 13 1 0 9 2 15 13 3 14 0 9 9 2
23 10 9 13 1 9 0 9 2 1 0 9 15 13 0 7 0 3 3 16 1 0 9 2
27 13 15 7 13 3 0 15 2 16 7 10 9 13 3 7 1 10 9 15 4 13 13 0 9 16 3 2
6 3 7 9 13 0 2
1 3
17 1 0 9 1 11 13 3 0 9 16 9 9 9 1 12 9 2
26 1 9 12 9 15 13 9 1 9 10 9 2 15 3 13 1 9 12 2 9 12 1 9 0 9 2
36 1 9 1 9 0 9 0 9 0 11 1 11 2 0 1 0 9 9 2 13 0 9 11 2 11 0 9 2 16 4 3 13 0 9 11 2
29 0 9 9 0 0 0 9 1 11 1 9 11 2 1 15 13 12 9 2 13 9 9 2 15 15 13 13 9 2
5 13 15 0 9 2
24 1 11 13 13 1 9 12 12 7 12 7 9 9 9 0 9 9 2 15 13 0 9 9 2
12 13 15 0 9 9 1 9 1 9 9 9 2
12 9 1 9 12 9 0 9 13 3 9 11 2
16 9 15 13 1 9 12 9 1 0 9 12 9 3 1 11 2
25 0 9 11 2 11 13 3 1 9 1 11 2 15 13 10 0 9 1 0 9 1 12 0 9 2
18 11 13 0 0 9 2 15 13 1 11 1 9 0 9 1 9 12 2
26 9 0 0 9 0 0 0 9 11 2 11 4 3 1 11 13 12 0 9 2 15 13 1 10 9 2
6 1 9 1 9 13 2
16 1 9 0 9 13 1 9 0 9 9 0 0 7 0 9 2
14 9 13 1 0 9 9 0 9 1 11 1 0 9 2
28 9 7 9 1 0 0 9 3 13 12 0 9 7 13 9 7 9 1 12 9 2 15 13 13 1 0 9 2
10 1 12 9 4 13 1 9 11 11 2
15 0 9 4 13 1 9 1 9 9 11 0 1 0 9 2
22 0 9 13 0 9 2 15 13 9 11 11 1 9 12 1 0 9 9 11 2 11 2
29 9 13 9 1 3 0 9 2 15 4 13 1 9 1 11 7 13 15 9 9 12 3 0 9 7 10 12 9 2
12 11 11 2 12 2 13 1 0 9 0 9 2
22 13 16 9 1 9 0 9 11 11 9 7 9 9 2 3 13 16 0 7 0 9 2
56 1 10 9 13 13 9 11 9 2 0 9 11 7 11 2 11 2 11 7 11 2 11 2 2 9 0 9 9 2 1 11 2 11 7 11 2 11 2 2 9 0 9 7 0 9 1 0 9 9 2 1 11 2 11 2 2
9 2 11 2 2 11 12 2 12 2
6 11 2 12 12 1 11
2 11 11
16 0 0 7 0 9 13 7 0 9 1 0 9 9 15 13 2
16 0 9 12 1 12 13 1 0 0 0 9 2 11 2 9 2
7 10 9 3 13 1 9 2
6 3 7 3 0 9 2
12 7 3 1 10 9 15 4 0 9 3 13 2
9 10 9 7 1 9 0 9 13 2
16 1 9 0 9 0 11 3 13 9 2 16 4 9 13 3 2
21 9 0 9 13 11 13 2 16 9 13 1 9 2 15 1 15 13 14 3 0 2
6 0 9 13 3 0 2
20 3 2 16 4 4 13 2 16 3 13 10 0 9 0 3 1 9 0 9 2
11 1 0 9 9 13 0 7 0 0 9 2
27 0 9 2 0 1 0 9 0 9 2 11 2 7 9 0 9 0 15 1 0 9 2 13 10 0 9 2
28 1 9 9 13 13 12 9 0 3 0 9 9 3 0 11 7 13 15 14 1 9 2 7 7 1 9 9 2
12 9 1 9 9 13 7 0 0 9 0 9 2
14 3 16 0 9 1 9 15 1 0 9 13 16 9 2
16 9 13 2 16 0 2 0 0 2 9 13 9 9 1 9 2
9 13 15 7 2 16 9 13 0 2
18 3 9 10 9 13 3 9 0 9 2 15 9 13 3 1 9 12 2
22 11 11 11 2 9 11 2 15 1 9 9 13 10 9 11 11 1 11 2 13 3 2
14 1 12 9 9 0 0 9 9 13 3 12 9 11 2
8 1 9 13 9 9 3 0 2
8 1 12 9 15 11 13 12 2
12 0 9 9 13 7 13 9 15 2 15 13 2
24 3 16 0 9 15 13 2 16 13 1 9 2 0 9 13 9 2 15 15 13 9 0 9 2
17 0 9 11 11 11 13 10 9 2 16 15 15 13 0 9 13 2
15 0 9 13 2 16 1 15 9 13 7 0 9 3 0 2
15 1 10 9 13 10 9 0 9 2 0 9 13 3 13 2
39 3 7 9 13 2 10 9 13 3 10 2 16 13 13 0 9 9 2 1 15 11 11 13 1 11 11 1 11 2 11 2 1 9 12 9 9 1 12 2
13 1 9 7 13 2 16 4 0 9 4 13 3 2
17 1 9 0 9 1 9 9 15 3 0 9 2 3 3 2 13 2
24 0 1 0 9 12 0 9 2 11 11 11 1 9 0 9 2 15 1 9 9 3 13 13 2
14 0 12 9 9 2 15 1 15 13 2 13 1 9 2
22 1 9 10 9 1 0 0 9 11 2 2 3 9 9 13 11 2 13 9 0 9 2
18 16 9 3 0 13 2 3 14 3 13 3 3 2 16 1 12 9 2
8 1 10 9 15 13 15 13 2
26 16 15 9 9 0 0 9 0 9 1 9 12 3 13 2 0 9 0 9 15 3 1 12 9 13 2
21 1 9 0 9 4 15 14 0 11 11 11 13 3 3 13 7 15 15 3 13 2
7 9 1 0 9 1 11 13
2 11 11
30 11 11 2 11 2 3 0 0 9 7 3 0 0 9 2 15 1 15 3 13 0 0 9 11 11 2 11 2 11 2
18 3 16 0 9 1 0 9 1 0 9 2 13 3 11 1 0 9 2
12 13 7 15 2 16 15 13 13 9 0 9 2
15 9 0 9 13 1 9 10 9 7 13 15 1 0 9 2
10 14 13 15 13 2 16 13 3 3 2
10 15 13 1 0 9 3 2 3 0 2
19 3 1 15 13 9 11 2 15 1 10 9 13 7 13 1 15 9 11 2
18 7 3 13 0 15 11 2 15 9 7 9 15 9 3 7 3 13 2
6 13 3 1 0 9 2
11 15 15 13 7 3 2 16 13 1 9 2
27 3 15 2 16 15 1 0 9 13 3 3 9 1 0 0 9 2 13 11 0 10 9 0 9 0 9 2
10 2 3 2 13 9 1 11 0 9 2
30 9 3 1 9 0 9 3 13 2 13 1 0 9 2 7 1 0 9 3 13 0 9 2 1 9 10 0 9 2 2
9 3 13 11 0 7 3 0 9 2
15 13 15 2 16 13 0 9 7 16 10 9 13 0 9 2
26 13 7 0 2 16 15 13 9 2 1 15 15 3 13 2 9 2 3 1 9 12 13 11 11 11 2
20 7 3 15 9 3 1 11 13 13 1 9 2 15 13 1 9 1 0 9 2
47 1 0 9 2 15 13 10 0 9 2 15 1 0 9 13 9 11 11 2 11 2 9 9 7 9 2 2 11 11 2 9 7 9 9 2 7 11 11 2 11 2 9 2 9 9 2 2
7 0 11 13 9 3 0 2
18 7 3 15 13 1 10 9 2 1 0 9 13 0 9 9 2 2 2
15 1 0 9 15 13 3 0 9 2 13 1 9 10 9 2
20 13 9 0 0 9 1 9 11 11 2 7 0 9 15 14 1 15 13 9 2
5 3 3 0 9 2
11 1 0 9 13 3 9 11 2 12 2 2
17 10 0 9 13 1 9 1 9 11 2 11 2 11 9 0 9 2
10 9 13 9 2 9 13 1 0 9 2
10 1 0 9 4 13 13 9 1 9 2
15 9 11 2 3 0 16 11 2 4 3 13 1 11 11 2
17 13 15 9 2 9 1 0 9 7 9 9 2 3 1 0 9 2
12 13 9 7 10 0 0 9 13 1 0 9 2
21 1 9 0 9 13 14 15 1 15 12 3 0 2 16 4 15 13 0 9 9 2
9 7 15 13 13 0 9 0 9 2
14 13 15 7 13 9 2 16 13 0 2 3 0 9 2
12 3 0 11 11 2 7 0 11 11 2 11 2
19 11 15 11 13 15 2 16 13 0 9 2 1 15 15 13 15 0 9 2
5 13 9 0 9 2
11 7 15 13 2 16 1 10 9 15 13 2
5 3 13 9 9 2
10 11 13 0 9 9 7 0 0 9 2
24 1 9 0 9 13 1 15 9 2 13 3 1 0 9 1 9 2 7 13 15 1 0 9 2
8 3 15 13 1 9 1 9 2
6 3 3 2 13 15 2
8 1 15 1 15 15 13 9 2
20 11 0 2 13 1 0 9 2 15 16 13 10 9 2 3 13 2 15 0 2
8 11 15 1 0 9 13 11 2
10 16 13 3 15 15 0 2 13 9 2
6 7 3 2 16 0 2
7 9 1 9 7 0 0 9
8 11 11 2 9 9 1 9 9
55 1 9 1 9 11 11 2 15 15 1 9 10 9 2 11 12 2 12 2 2 13 0 9 1 9 2 16 13 1 11 9 9 1 9 2 13 13 2 16 15 15 3 13 7 13 2 16 10 9 3 13 14 1 11 2
33 16 9 3 13 9 0 7 0 15 13 3 16 15 2 16 3 13 7 9 0 9 7 9 7 0 10 9 1 9 13 7 13 2
33 9 13 13 3 0 2 9 7 9 13 15 1 15 2 16 9 1 9 9 1 9 3 7 1 15 13 3 0 16 1 0 9 2
15 13 0 3 13 2 10 9 13 0 9 9 2 0 9 2
16 7 13 3 3 0 15 9 1 0 9 7 1 0 9 13 2
23 13 3 7 13 9 7 9 7 9 13 15 3 0 0 9 2 7 7 9 0 9 9 2
24 13 3 9 2 16 15 3 13 2 16 4 13 0 13 15 9 1 9 3 7 1 0 9 2
10 13 7 13 9 0 7 3 15 0 2
23 13 10 9 2 3 13 3 0 9 1 9 13 0 9 2 7 3 9 0 9 3 13 2
8 3 15 3 3 13 3 3 2
20 16 15 3 0 13 2 13 3 7 9 11 2 15 1 9 13 7 9 9 2
52 9 2 16 9 9 1 9 7 10 9 0 9 0 13 2 13 7 9 0 9 11 1 0 11 2 15 13 1 9 10 2 9 2 1 11 11 9 0 2 7 15 15 13 0 9 0 9 1 9 7 11 2
30 9 13 1 9 1 9 9 3 0 2 0 9 2 15 1 15 13 1 0 9 15 16 0 0 9 2 9 0 9 2
33 0 9 13 7 14 12 9 9 9 2 3 15 13 7 13 9 7 3 15 9 0 9 13 3 7 1 0 9 2 1 9 3 2
23 10 9 15 13 3 15 9 2 1 15 13 9 2 16 1 15 4 9 13 1 0 9 2
34 13 15 3 7 0 0 2 9 1 9 2 0 7 0 9 2 13 15 7 3 7 3 0 7 0 9 1 9 9 2 0 9 3 2
18 0 9 15 1 10 9 3 13 9 9 0 7 0 14 1 15 9 2
19 9 2 16 15 9 13 13 2 10 9 13 1 0 9 0 9 9 9 2
8 9 13 1 9 9 15 13 2
47 3 2 16 1 12 9 12 0 9 15 3 13 14 1 10 9 0 0 9 2 1 0 9 3 13 15 9 1 12 9 3 2 1 11 15 9 13 1 9 1 12 1 12 9 1 9 2
24 16 4 0 9 13 1 10 9 7 3 2 3 13 9 9 1 10 9 2 13 4 15 0 2
32 15 13 3 0 2 16 1 9 9 13 1 10 9 14 9 2 15 15 9 13 7 13 3 7 3 7 3 1 0 9 0 2
30 16 1 9 0 9 4 3 13 0 9 7 16 9 3 13 9 9 3 13 2 16 3 15 4 13 13 10 0 9 2
14 0 1 9 9 13 13 3 2 0 13 3 3 13 2
11 13 1 15 7 13 10 0 7 0 9 2
6 9 13 7 0 7 0
4 11 11 2 9
16 13 14 0 2 16 9 13 1 9 9 2 13 0 9 9 2
27 3 7 3 4 13 2 13 2 14 9 9 9 1 0 9 2 13 11 12 2 12 2 2 1 0 9 2
20 1 9 0 9 13 9 0 9 9 9 1 0 0 9 2 15 4 3 13 2
45 9 9 15 16 3 2 16 13 1 9 0 1 0 2 2 7 1 0 9 9 9 1 9 2 13 1 9 1 9 2 14 3 3 15 13 2 15 13 7 16 0 13 1 9 2
40 1 12 9 3 1 9 13 9 9 2 3 0 9 0 16 3 0 0 9 2 13 16 6 9 2 2 7 3 13 3 10 9 1 9 1 9 2 15 13 2
36 7 1 0 12 9 3 13 9 0 0 9 1 9 0 9 2 15 13 2 16 0 9 10 9 15 13 1 10 0 9 7 1 0 9 9 2
40 3 0 0 9 2 13 0 2 13 9 1 9 2 9 0 9 9 2 3 0 2 7 9 2 9 9 9 1 0 0 9 2 1 9 9 9 3 13 2 2
5 9 13 14 12 2
15 13 15 9 1 9 9 2 1 0 9 1 10 0 9 2
11 13 1 15 9 0 9 1 0 9 9 2
48 1 9 1 15 9 1 0 9 7 9 13 3 1 0 9 0 9 2 3 1 0 9 12 0 9 2 16 4 2 3 3 7 3 2 13 0 0 9 9 3 0 2 9 3 3 0 2 2
58 9 9 2 9 1 9 2 13 16 0 9 7 13 15 2 1 9 9 9 7 9 2 13 1 9 2 16 3 1 3 0 9 0 7 7 14 3 3 0 9 9 2 9 2 0 9 13 3 9 2 7 3 3 0 9 9 2 2
47 13 3 3 13 10 9 16 9 1 10 7 15 9 9 2 7 9 2 15 4 13 1 0 9 2 2 7 16 9 1 9 9 13 13 2 13 7 1 15 2 16 3 13 1 0 9 2
14 9 2 1 9 1 9 2 4 0 0 3 13 3 2
43 16 13 13 15 0 1 9 1 9 1 9 1 0 9 2 7 13 9 7 9 15 3 0 2 15 13 13 0 9 2 16 1 9 9 2 9 7 9 2 15 13 9 2
46 15 13 7 0 1 15 0 9 13 1 0 9 2 3 7 3 2 13 13 0 9 9 3 1 9 0 9 2 0 9 2 7 0 1 9 1 3 0 0 9 2 1 0 9 2 2
17 9 4 13 3 16 9 13 0 9 2 15 7 13 9 0 9 2
28 0 9 9 2 11 2 11 2 11 0 2 2 2 15 13 1 0 9 7 13 15 2 13 15 9 3 9 2
10 0 9 1 10 9 15 13 0 9 2
29 3 2 9 0 1 9 1 0 9 13 2 9 2 9 1 9 2 0 9 2 0 9 9 1 9 1 9 3 2
21 0 9 10 0 9 3 4 2 1 9 9 2 13 4 3 13 0 9 3 0 2
30 0 9 1 0 0 9 2 0 2 1 9 9 2 13 9 1 15 2 16 13 0 1 0 2 0 2 0 2 2 2
37 16 15 13 2 16 0 9 13 13 0 2 0 7 0 9 2 3 15 13 13 2 3 15 3 1 10 9 0 9 2 3 3 0 9 2 13 2
10 1 9 1 15 13 9 0 0 9 2
62 16 0 9 13 1 9 0 9 1 9 7 3 13 0 0 9 1 9 0 9 9 9 2 14 9 0 9 2 2 7 2 9 13 3 13 3 2 3 7 1 9 2 15 15 13 1 0 9 2 3 15 13 13 2 16 13 14 12 9 2 9 2
45 16 9 0 9 3 13 0 9 1 9 9 3 0 9 1 9 9 10 9 7 0 9 1 9 9 13 1 9 1 9 0 9 7 9 0 9 2 13 1 9 0 9 10 9 2
12 14 2 10 9 3 13 1 9 12 9 9 2
4 7 3 3 2
18 1 15 3 13 0 15 3 13 2 16 4 0 9 13 10 0 9 2
13 13 15 1 9 0 9 2 7 3 7 0 9 2
23 13 9 0 2 9 0 0 9 2 9 9 1 0 9 2 15 15 1 9 0 9 13 2
15 13 15 9 9 7 3 9 0 9 3 0 1 9 0 2
6 1 9 13 0 0 9
12 11 11 2 9 9 9 0 9 1 0 9 11
28 1 9 1 0 9 0 9 0 9 13 9 11 11 3 0 9 2 1 11 12 2 12 2 2 1 10 9 2
38 13 0 2 0 9 1 0 1 0 9 9 7 1 9 2 16 2 2 2 13 0 13 9 2 9 7 0 9 10 9 1 10 7 15 9 15 13 2
19 1 15 1 0 9 13 9 9 1 10 9 0 9 0 9 9 9 9 2
26 13 3 9 1 9 9 2 9 2 15 14 13 2 16 11 2 11 3 13 1 9 7 9 9 11 2
16 13 3 1 9 1 15 2 7 1 9 2 15 9 13 9 2
19 3 2 13 1 0 9 0 9 7 9 0 9 13 9 9 1 9 12 2
14 0 9 13 10 9 13 0 9 2 13 15 7 13 2
12 13 3 2 16 0 9 13 9 1 0 9 2
25 1 9 0 9 7 9 7 9 0 7 10 0 9 13 15 13 7 13 0 9 1 9 0 9 2
9 9 9 13 1 0 9 9 9 2
16 15 1 10 9 13 0 9 2 3 16 1 9 9 0 9 2
19 13 3 9 9 2 15 7 13 13 2 16 4 13 9 1 0 0 9 2
8 13 3 10 9 1 0 9 2
21 0 9 13 0 9 2 9 0 9 7 9 0 9 9 2 0 7 0 0 9 2
12 1 9 9 13 1 12 9 1 9 0 2 2
17 9 9 15 13 3 13 14 0 9 2 9 9 14 0 9 3 2
30 9 1 10 9 13 0 7 0 13 1 0 9 2 16 4 13 0 13 9 9 0 9 1 9 7 9 9 7 9 2
10 13 3 2 16 0 9 13 0 9 2
19 1 9 2 15 13 13 0 9 9 7 15 15 13 13 2 13 13 9 2
21 10 9 13 1 9 9 9 1 9 9 1 9 14 1 9 9 9 1 0 9 2
15 15 10 9 15 7 13 14 1 9 9 2 15 13 9 2
16 13 4 13 9 2 3 2 9 0 0 9 1 9 0 9 2
22 3 1 10 9 13 1 0 9 0 9 2 9 14 1 9 0 2 0 1 15 9 2
11 3 9 10 9 13 3 13 1 9 9 2
13 3 9 13 0 9 2 13 2 14 15 9 9 2
18 1 9 13 9 1 0 9 7 9 1 9 1 0 9 3 3 0 2
28 7 16 4 15 9 3 1 9 9 0 9 13 1 9 13 11 1 9 1 9 2 9 9 10 9 13 13 2
10 13 0 0 9 13 0 0 9 9 2
9 3 13 13 0 9 13 7 9 2
25 9 13 1 15 2 16 9 0 9 13 1 0 9 3 0 7 13 15 13 14 0 7 0 9 2
18 9 1 3 0 0 9 2 3 2 11 2 13 9 10 9 3 9 2
10 7 3 13 15 1 0 0 9 9 2
42 1 0 0 9 0 9 11 11 13 12 5 0 1 0 9 9 1 9 0 0 9 2 12 5 9 13 1 3 7 3 0 1 0 9 9 0 9 2 9 7 9 2
37 3 0 13 9 12 5 9 2 16 9 4 13 13 9 2 15 4 13 0 9 7 9 13 0 9 2 16 4 15 13 4 13 9 1 0 9 2
6 10 9 9 13 9 2
17 9 13 2 16 9 13 9 2 7 4 13 1 9 1 10 9 2
5 11 11 13 3 2
12 13 1 9 1 0 9 9 2 15 13 9 2
7 0 9 11 13 1 0 9
17 0 9 13 13 9 0 9 2 13 1 9 1 11 9 9 11 11
2 11 11
36 1 0 12 9 13 0 9 3 12 1 0 9 1 0 9 2 15 13 9 9 1 15 2 1 10 0 9 4 1 0 9 13 10 0 9 2
14 14 1 10 0 9 13 0 9 3 12 0 0 9 2
21 16 4 13 9 1 9 15 0 9 3 2 13 10 9 0 9 0 0 9 11 2
22 1 0 9 4 13 0 9 0 9 2 9 7 9 9 1 9 7 0 9 11 11 2
10 3 13 0 13 3 0 9 0 9 2
17 12 1 9 13 2 16 15 10 9 9 3 13 1 10 0 9 2
23 13 1 15 13 9 1 0 9 2 15 13 3 3 0 2 16 13 1 9 12 7 12 2
39 13 15 9 0 9 2 10 0 7 3 1 15 0 0 9 9 1 0 9 13 3 0 3 2 16 4 15 13 0 9 1 0 9 7 1 9 0 9 2
13 10 0 9 13 7 0 2 7 7 13 13 2 2
29 7 15 9 13 13 3 9 1 0 9 1 15 2 16 13 1 10 9 2 7 3 1 9 1 0 0 0 9 2
10 15 13 13 0 9 0 9 0 9 2
36 10 9 15 13 3 3 16 9 1 0 9 1 9 0 9 9 2 3 7 1 9 3 0 2 0 9 2 15 4 15 13 13 0 0 9 2
13 10 9 13 0 9 0 9 9 7 9 10 9 2
15 3 4 13 0 0 9 1 0 9 1 9 9 0 9 2
11 15 10 9 3 13 0 9 0 12 9 2
32 0 9 2 15 4 13 2 13 9 10 12 9 3 7 3 0 2 3 0 9 13 9 0 2 7 2 0 9 7 9 9 2
10 15 13 1 9 0 0 9 12 9 2
34 1 10 9 9 2 12 9 13 2 16 9 13 13 15 2 15 15 13 9 13 2 7 15 15 13 13 13 15 2 15 15 9 13 2
17 13 15 3 1 9 2 3 1 0 9 2 0 3 1 9 9 2
16 1 10 9 13 3 3 9 7 9 10 0 9 13 3 0 2
20 0 9 0 0 9 13 2 16 3 13 0 7 0 9 1 0 7 0 9 2
13 1 0 9 13 0 9 9 9 7 9 0 9 2
18 1 0 9 13 3 0 13 1 9 9 0 9 2 3 10 9 13 2
13 9 10 12 9 9 4 3 13 1 9 9 0 2
13 15 15 1 0 9 0 9 13 7 9 3 0 2
12 13 13 9 0 9 2 15 4 3 3 13 2
11 13 3 2 1 0 0 9 2 9 9 2
16 15 13 3 0 1 9 0 9 2 15 10 9 13 7 13 2
23 1 9 2 16 15 13 1 0 9 2 13 9 3 14 9 2 7 7 0 9 10 9 2
9 3 15 13 3 7 1 9 0 2
13 1 15 4 13 4 1 15 13 3 0 0 9 2
23 0 0 9 0 9 1 9 13 1 12 9 9 2 1 9 0 0 0 9 2 0 9 2
15 9 9 13 3 9 0 9 16 0 0 9 10 0 9 2
26 3 1 15 13 0 7 0 9 2 9 10 9 2 15 13 1 10 9 14 0 2 7 7 3 0 2
12 3 13 12 0 9 13 1 9 12 10 9 2
18 15 13 3 0 9 2 15 13 1 9 9 1 0 0 9 3 0 2
11 3 4 15 0 9 13 1 10 9 13 2
8 10 9 3 1 0 9 13 2
16 15 2 3 9 1 9 7 0 9 7 0 9 13 0 9 2
20 3 13 1 0 2 16 4 15 9 7 9 0 9 13 9 9 0 9 3 2
22 9 9 0 9 13 13 0 9 2 13 3 1 9 0 9 2 3 13 0 9 9 2
18 0 9 9 15 3 13 3 9 2 7 10 9 9 9 13 3 0 2
11 3 4 13 0 0 9 1 9 0 9 2
11 0 0 9 13 2 15 13 3 3 0 2
20 1 9 12 15 15 2 7 3 3 13 1 15 2 16 9 9 13 7 3 2
16 16 13 0 9 9 12 13 0 9 0 9 7 13 0 9 2
29 13 15 7 0 2 13 4 15 1 0 9 1 15 0 0 9 2 13 4 13 9 0 9 7 9 4 13 13 2
12 1 0 0 9 3 10 0 9 16 9 13 2
36 7 13 3 0 9 14 0 9 2 0 9 1 9 2 15 13 13 14 9 2 7 7 0 9 2 10 9 13 3 3 0 1 9 0 9 2
10 15 13 1 0 9 0 9 1 9 2
30 1 0 9 15 13 13 9 10 0 9 2 15 13 9 0 9 7 9 0 9 2 3 3 9 9 9 15 9 9 2
22 15 13 3 0 9 2 15 4 13 2 16 0 0 9 13 3 0 7 0 10 9 2
7 10 9 9 13 0 9 2
10 3 13 1 9 9 9 0 7 0 2
12 3 13 9 9 12 10 9 9 1 0 9 2
26 3 13 3 9 9 0 2 15 13 0 9 2 16 0 9 13 3 10 9 0 9 1 9 7 9 2
35 0 10 9 9 4 13 4 3 13 2 9 9 4 15 13 3 13 14 1 0 0 9 0 9 7 9 0 9 4 13 13 9 0 9 2
18 1 9 1 9 9 0 9 13 13 3 1 0 9 0 2 0 9 2
8 15 15 13 0 0 9 13 2
11 0 9 0 9 7 3 15 1 0 9 2
15 0 9 7 10 0 9 1 0 9 13 1 10 9 0 2
14 7 13 13 2 16 1 10 9 13 12 7 12 9 2
15 3 4 13 1 9 0 9 2 15 3 13 1 9 0 2
10 13 3 4 13 1 9 0 0 9 2
15 9 0 9 13 13 7 1 9 9 1 10 0 0 9 2
12 13 3 3 1 0 9 1 9 16 1 9 2
13 3 3 13 9 0 9 1 9 1 9 0 9 2
9 14 3 2 3 2 7 3 3 2
23 0 9 13 9 2 15 13 13 3 2 3 13 9 2 10 9 7 0 9 10 0 9 2
9 1 10 9 13 3 9 3 0 2
7 13 9 9 7 10 9 2
9 10 9 3 13 9 1 0 9 2
7 9 9 13 3 0 9 2
8 13 3 1 9 10 0 9 2
24 9 7 13 4 13 10 0 9 3 2 3 15 10 9 13 13 2 3 10 0 9 13 13 2
13 9 2 15 4 13 1 0 9 2 13 3 0 2
16 15 15 15 3 13 2 7 9 7 9 13 3 10 0 9 2
18 16 10 9 0 9 3 13 2 0 2 3 2 0 9 2 15 13 2
4 9 13 3 2
5 15 13 10 9 2
21 13 7 1 15 2 16 4 9 10 9 13 14 3 2 3 1 0 9 13 13 2
25 13 9 0 9 0 9 3 9 13 10 9 9 0 9 1 9 1 10 9 1 9 1 10 9 2
7 0 4 9 13 16 9 2
12 13 3 1 0 9 15 0 9 7 10 9 2
39 15 15 13 0 9 2 15 13 9 11 2 13 15 1 0 0 9 2 7 1 0 9 0 1 9 0 9 2 15 1 10 9 13 3 7 9 0 9 2
13 13 3 1 9 0 2 0 2 0 2 0 3 2
16 13 4 3 2 16 9 9 10 0 9 3 13 1 0 9 2
19 3 2 1 9 9 13 13 9 9 1 9 9 15 10 0 9 9 11 2
10 3 13 3 10 9 0 1 9 11 2
19 1 0 0 9 7 9 1 9 1 11 13 3 0 15 1 10 9 13 2
19 1 11 13 9 2 15 15 0 0 9 13 1 9 0 9 7 9 11 2
16 7 13 9 15 1 0 9 0 9 1 0 9 1 0 9 2
30 16 3 13 1 11 11 2 4 13 1 0 9 14 12 12 10 9 2 7 14 14 1 12 2 1 15 9 13 9 2
19 3 15 7 13 1 9 2 3 1 11 4 13 11 2 13 3 15 13 2
22 3 13 13 10 0 9 2 15 13 0 1 9 0 9 2 0 1 10 9 3 3 2
10 15 7 13 2 16 15 13 9 9 2
12 13 13 0 9 1 10 9 7 13 10 9 2
10 3 1 10 9 13 9 0 9 9 2
18 3 13 1 9 15 2 15 13 9 3 7 15 13 9 1 0 9 2
15 0 9 13 0 9 9 2 1 15 15 13 9 7 13 2
23 15 1 15 13 9 2 16 13 3 9 0 9 7 16 4 10 9 9 13 3 0 9 2
15 3 15 7 13 13 2 3 13 15 0 2 0 7 0 2
24 3 15 1 0 9 9 13 9 1 9 7 9 2 16 15 7 1 10 0 9 9 13 3 2
9 0 9 15 3 1 0 9 13 2
15 13 15 7 3 9 0 16 0 7 13 1 9 0 9 2
9 9 15 1 10 9 9 13 15 2
27 15 13 1 10 9 2 13 0 9 7 13 2 3 13 0 13 3 0 2 7 14 3 0 9 1 9 2
10 15 13 3 3 2 16 15 0 13 2
7 13 3 10 9 3 0 2
6 1 0 9 13 0 2
25 9 0 9 13 3 0 2 13 3 15 2 15 13 13 1 0 9 7 9 9 16 9 7 9 2
13 15 13 0 9 2 1 15 13 0 0 0 9 2
16 3 13 0 2 16 1 9 0 9 13 13 0 9 0 9 2
22 3 13 0 13 9 10 0 0 9 2 16 15 13 3 2 1 0 9 1 0 9 2
20 15 13 13 0 9 0 9 2 1 10 9 7 9 13 2 16 13 3 0 2
8 0 9 13 0 9 0 9 2
21 3 1 9 0 9 9 2 13 15 1 10 9 3 1 9 9 0 9 1 11 2
27 0 9 13 2 16 15 0 9 13 0 9 1 9 10 9 7 13 3 15 2 15 13 1 10 9 0 2
39 13 15 7 2 16 9 13 4 13 3 0 9 10 9 2 3 4 13 10 0 9 2 13 2 10 9 0 9 1 15 13 7 15 15 13 1 9 0 2
9 15 13 1 10 9 0 9 9 2
8 13 15 0 0 9 9 3 2
11 3 3 9 10 9 9 13 13 0 9 2
12 1 10 0 9 13 3 0 9 1 9 9 2
20 7 15 1 0 9 7 3 3 13 3 0 0 9 9 2 15 13 13 0 2
10 13 1 15 9 2 14 9 7 9 2
22 9 13 10 9 1 9 0 9 1 10 9 1 9 2 16 4 13 10 0 0 9 2
5 0 2 3 0 2
27 13 15 3 2 16 1 0 9 13 0 9 9 2 15 3 1 9 0 9 13 2 15 3 13 3 13 2
24 13 15 13 7 3 3 2 0 9 0 9 13 13 1 9 7 3 13 3 13 0 0 9 2
13 3 15 3 3 13 0 9 13 0 9 0 9 2
9 13 0 1 10 9 1 9 9 2
21 9 0 0 9 2 1 15 3 13 9 2 15 1 0 9 3 13 1 0 9 2
25 13 2 16 1 9 2 16 13 3 0 2 7 13 0 2 3 0 9 1 9 0 0 9 9 2
12 0 9 13 0 9 2 15 3 2 15 3 2
13 13 7 1 9 9 2 3 15 1 10 9 13 2
12 0 13 3 3 3 9 0 9 1 9 9 2
14 1 10 9 15 13 9 0 9 7 9 1 0 9 2
21 9 9 9 1 0 9 13 9 3 1 3 0 2 9 15 3 7 1 9 13 2
6 3 0 13 0 9 2
33 9 13 2 16 0 1 9 13 7 1 0 9 9 10 9 9 13 2 7 3 15 3 3 1 10 9 13 7 9 10 9 13 2
15 7 1 9 0 9 7 13 1 10 0 9 9 15 13 2
17 3 15 13 2 16 0 9 13 2 3 13 10 9 0 9 0 2
14 9 1 9 2 15 13 1 15 9 9 1 0 9 2
31 1 9 9 13 2 16 4 15 13 9 1 9 0 0 9 7 10 3 0 9 1 9 9 2 3 0 2 3 7 0 2
5 9 13 10 9 2
20 10 9 4 13 15 2 16 9 13 9 9 2 7 2 9 2 9 7 9 2
10 13 9 1 9 0 9 7 0 9 2
21 9 13 9 2 1 15 13 13 9 9 2 15 15 13 3 1 0 9 2 9 2
33 0 9 9 13 2 16 4 15 13 3 0 10 10 9 2 16 4 13 9 3 0 9 7 16 4 13 14 3 0 9 0 9 2
9 0 9 15 13 13 0 9 1 9
40 0 9 0 9 2 15 13 9 9 3 13 2 13 1 9 0 9 3 10 9 9 1 9 9 1 0 9 1 11 2 11 2 0 11 2 11 7 3 11 2
10 1 9 15 1 9 13 3 0 9 2
17 1 11 3 13 9 9 2 15 15 1 9 0 0 9 9 13 2
52 1 11 11 1 0 9 1 0 11 2 15 13 9 9 2 15 10 3 0 9 9 13 1 10 0 9 1 0 3 3 2 16 1 0 9 3 13 9 9 9 0 9 0 9 9 7 9 0 9 1 9 2
22 0 9 2 15 15 3 13 2 4 13 1 0 0 2 0 9 0 9 9 7 9 2
22 13 9 9 13 1 9 0 9 7 0 9 7 1 0 9 2 7 3 13 10 9 2
8 0 9 13 9 9 9 9 2
39 10 9 3 13 13 7 3 2 16 3 9 9 13 1 9 7 9 9 2 15 4 9 0 9 1 9 13 13 13 2 13 11 11 11 1 9 1 9 2
6 1 9 13 0 9 2
18 13 15 1 0 9 7 16 9 9 13 1 10 9 2 13 9 13 2
14 10 9 13 0 13 7 0 9 0 9 2 13 11 2
14 0 9 9 0 9 13 0 9 1 11 1 9 12 2
24 13 15 1 12 9 2 1 15 12 13 0 3 1 9 0 9 2 13 11 11 2 2 11 2
13 9 9 7 0 9 13 9 1 0 9 1 0 11
5 9 11 11 2 11
6 11 11 7 9 1 11
18 3 13 9 9 1 9 0 9 0 9 0 9 2 11 11 2 11 2
11 13 15 1 9 12 1 11 1 0 9 2
16 1 12 9 13 13 9 1 11 2 3 15 13 1 0 9 2
12 9 9 1 9 12 13 10 9 14 1 11 2
19 16 15 1 12 9 13 1 11 2 13 15 13 0 9 1 9 0 9 2
13 1 9 12 13 1 10 9 1 11 0 0 9 2
21 13 15 1 9 10 0 9 7 16 0 9 13 1 9 15 0 0 7 0 9 2
10 9 2 11 11 2 11 12 2 12 2
4 9 13 12 9
30 0 9 1 0 0 9 2 1 15 12 2 9 13 9 0 0 9 6 11 2 13 13 1 12 9 3 9 12 9 2
12 0 13 3 9 7 9 9 7 0 0 9 2
21 1 9 9 11 2 10 9 15 9 1 11 13 2 13 9 1 11 3 12 9 2
11 10 9 7 9 13 12 0 9 0 11 2
32 0 9 13 9 9 3 1 11 11 7 9 11 11 2 15 15 3 13 3 1 9 1 11 11 7 3 1 0 9 1 11 2
1 3
14 11 11 13 1 0 9 0 9 0 0 9 0 9 2
18 9 15 4 13 1 9 9 7 9 7 13 4 13 3 1 9 9 2
21 9 15 1 9 13 0 9 11 2 3 11 3 13 3 1 11 11 7 11 11 2
5 0 11 13 1 11
19 0 9 0 11 12 2 12 13 3 1 12 9 1 0 0 9 1 9 2
16 0 9 9 1 9 1 9 4 13 13 14 1 9 1 9 2
9 1 9 15 3 13 1 12 9 2
66 1 9 1 11 2 0 9 2 11 2 11 7 11 1 11 13 3 9 11 11 7 11 2 0 9 2 9 2 11 7 11 2 11 1 11 2 11 2 9 12 2 11 11 7 3 2 9 11 2 3 13 3 2 9 9 2 11 2 11 11 7 0 2 2 11 2
5 15 2 3 2 3
28 9 11 1 11 13 3 1 12 9 1 9 1 11 7 0 0 9 1 0 9 1 0 9 9 0 2 9 2
7 9 13 9 9 0 9 2
14 9 0 0 9 13 13 1 9 11 11 1 0 9 2
5 9 1 9 0 9
2 11 11
10 3 1 0 9 13 0 9 9 9 2
23 12 3 0 9 13 14 1 0 9 9 2 15 3 13 1 9 7 1 9 0 11 3 2
39 9 13 1 0 9 0 3 0 9 2 1 12 9 2 12 2 9 12 2 4 11 11 2 10 9 11 7 11 11 7 9 11 1 11 13 0 9 9 2
11 13 7 13 1 0 9 14 1 12 9 2
11 0 9 9 9 13 0 9 1 0 9 2
23 9 9 11 11 7 11 11 13 2 16 4 1 15 13 9 0 1 9 0 9 3 3 2
11 9 7 13 1 9 0 1 0 0 9 2
26 9 13 9 3 1 12 9 0 9 2 0 2 11 2 9 2 9 2 9 15 0 7 0 9 2 2
24 12 0 9 4 13 9 2 15 15 13 13 9 2 1 15 1 11 11 13 0 9 3 3 2
24 9 9 13 13 3 3 7 9 2 13 9 11 2 0 0 9 1 9 9 13 3 3 3 2
25 0 11 1 0 9 13 0 9 2 15 4 13 4 13 14 1 0 9 2 7 7 1 0 9 2
12 3 13 9 1 0 9 0 9 2 11 11 2
9 15 3 1 9 9 0 9 13 2
25 11 2 12 2 13 9 1 0 2 11 1 11 7 1 9 12 13 16 9 1 0 9 0 9 2
20 0 9 15 1 9 13 3 2 3 16 1 9 0 9 11 11 2 12 2 2
17 9 0 9 13 0 9 9 11 11 2 9 0 0 9 1 11 2
49 9 9 0 0 9 0 9 4 13 13 3 9 0 11 2 1 11 0 11 2 11 11 3 2 2 7 13 0 0 9 2 0 0 9 2 11 0 2 15 13 0 9 2 15 15 9 13 2 2
13 0 0 11 13 7 0 0 9 0 7 0 9 2
25 9 13 12 0 9 2 1 9 13 11 11 0 9 1 0 9 7 0 9 11 13 0 0 11 2
19 0 7 0 9 1 9 4 13 0 9 0 11 7 0 0 9 1 11 2
15 9 0 9 2 15 9 13 2 13 0 0 2 0 9 2
23 15 14 13 1 9 2 9 7 0 9 2 7 1 0 9 11 11 13 0 9 0 9 2
12 1 0 9 0 9 13 3 0 9 1 9 2
36 0 9 2 15 4 15 13 13 12 2 9 2 4 13 1 9 9 7 4 1 15 3 13 0 9 11 11 2 15 13 9 1 11 1 11 2
18 9 0 9 13 9 9 7 9 15 3 4 13 13 1 10 0 9 2
2 0 11
1 9
2 11 11
24 0 2 0 9 13 3 1 9 1 11 0 0 9 2 3 15 13 9 9 7 9 11 11 2
13 11 15 13 9 12 1 0 9 1 9 1 11 2
21 1 11 2 3 15 10 9 3 13 16 0 9 2 15 13 9 0 12 9 9 2
46 0 9 0 9 2 9 9 2 0 9 1 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 7 0 11 2 7 10 9 2 0 3 1 0 9 2 13 9 3 14 3 2
18 1 11 11 13 1 9 2 13 1 0 9 9 1 0 7 0 9 2
23 1 11 13 1 0 9 1 9 10 9 1 9 2 1 15 13 1 9 13 9 7 9 2
35 7 1 11 3 3 3 13 2 15 16 16 0 9 13 1 9 0 9 7 13 10 0 9 2 10 9 2 15 13 1 0 9 2 2 2
35 3 3 7 3 0 0 9 3 13 1 0 9 9 9 2 1 1 10 9 2 0 9 9 2 7 1 1 9 10 9 13 15 0 9 2
19 1 9 3 3 13 11 2 3 9 7 9 0 9 2 9 0 1 9 2
4 3 13 14 2
17 1 15 15 0 9 16 0 9 1 0 9 9 3 3 13 13 2
21 1 15 4 14 3 3 13 9 2 15 13 0 9 7 15 13 1 10 0 9 2
9 14 2 10 15 13 1 0 11 2
13 7 3 2 1 9 13 7 10 9 2 10 9 2
30 3 1 15 2 15 1 11 13 2 1 0 9 9 13 1 9 3 2 7 13 3 0 9 1 0 9 0 9 11 2
5 3 15 3 13 2
25 16 15 13 13 0 9 0 9 0 2 0 7 0 9 1 0 9 2 3 9 0 9 3 13 2
10 0 9 2 11 12 2 12 2 12 2
36 13 15 9 11 2 16 0 9 1 9 13 2 16 0 9 13 0 2 16 1 9 1 12 9 4 0 9 13 9 1 0 9 1 0 9 2
31 13 2 14 1 0 9 2 3 1 9 2 16 9 13 2 16 15 15 9 13 2 4 13 10 9 13 14 1 9 9 2
6 1 9 11 11 2 11
4 0 2 2 2
8 2 11 12 2 12 2 12 2
16 3 0 9 15 13 1 9 2 15 1 0 9 13 14 13 2
7 3 13 3 13 1 9 2
20 16 13 15 9 15 2 16 4 15 13 1 10 9 2 7 13 3 10 9 2
11 15 3 9 3 13 7 3 2 7 3 2
18 13 7 10 9 2 7 9 1 9 10 9 1 10 9 1 0 9 2
7 13 15 1 0 0 9 2
16 9 9 15 13 2 16 9 1 0 9 15 4 13 7 13 2
11 13 15 3 2 16 1 0 9 13 9 2
25 10 9 15 0 9 13 9 7 13 15 2 16 13 9 2 16 4 15 1 15 1 9 13 3 2
6 1 9 11 11 2 11
2 9 9
23 3 0 9 11 11 1 9 0 9 15 3 13 1 9 1 9 12 1 9 9 11 11 2
20 1 3 12 9 1 15 0 9 13 3 2 3 1 0 9 9 11 11 11 2
23 0 9 11 11 15 1 9 13 3 3 2 7 15 3 13 0 7 0 9 9 11 11 2
8 2 11 2 2 11 2 12 2
5 1 9 2 2 2
8 2 11 12 2 12 2 12 2
36 16 9 11 13 2 16 15 9 13 9 7 1 9 2 15 13 1 10 0 9 7 9 15 0 2 13 15 9 9 1 9 1 0 9 9 2
14 1 15 13 9 9 15 3 0 16 0 9 10 9 2
26 1 0 9 4 13 1 15 9 7 3 13 0 2 7 15 3 13 2 16 9 0 9 13 1 15 2
57 7 16 15 9 0 9 2 3 16 9 9 11 2 13 7 13 10 9 2 13 2 3 4 13 13 1 9 7 1 9 0 15 0 9 1 10 9 2 15 15 13 1 9 9 2 1 9 9 0 9 7 1 0 9 0 9 2
13 13 15 3 2 3 14 9 13 14 12 5 9 2
6 1 9 11 11 2 11
7 13 9 14 9 1 9 2
16 9 9 3 13 1 0 9 1 9 1 9 9 0 0 9 2
11 10 9 13 1 0 9 0 1 9 12 2
26 3 1 0 9 0 9 9 7 9 11 2 11 16 12 1 0 9 4 13 0 9 2 15 13 13 2
24 3 0 9 1 15 2 15 15 3 13 2 15 3 13 2 1 0 15 3 13 13 9 9 2
13 13 15 7 9 1 9 0 9 2 3 3 0 2
23 12 1 0 9 3 13 16 9 1 0 9 0 0 9 2 1 15 15 13 1 9 13 2
8 13 15 1 9 11 7 11 2
8 10 9 7 4 3 15 13 2
26 3 1 0 9 15 13 0 9 1 9 0 9 2 9 1 0 9 13 9 7 9 1 9 0 9 2
9 9 12 7 13 15 9 1 9 2
11 3 1 9 12 15 9 3 13 1 9 2
34 1 9 9 2 15 4 13 9 11 7 9 9 2 15 3 13 1 9 0 9 2 7 13 1 10 9 3 2 3 1 15 13 9 2
17 1 0 9 13 1 9 0 9 2 15 14 13 1 11 3 0 2
25 1 0 9 15 13 0 7 0 9 1 9 9 2 7 10 9 3 13 9 0 9 1 0 9 2
19 0 9 1 0 9 0 9 13 13 0 7 0 16 10 0 3 0 9 2
16 9 9 4 13 0 9 7 13 3 13 1 9 0 9 3 2
28 13 2 16 9 9 7 9 9 4 1 9 13 0 9 1 15 9 7 3 1 9 15 2 15 15 15 13 2
6 1 9 11 11 2 11
4 15 0 9 13
28 1 11 13 12 2 12 2 12 13 9 11 2 11 2 0 1 9 11 2 11 2 11 12 2 12 2 2 2
25 1 10 0 9 13 7 14 14 3 10 9 7 9 2 0 2 16 1 9 9 13 9 7 9 2
38 9 2 11 13 0 9 11 13 12 2 12 2 12 1 0 9 2 7 1 9 9 2 3 2 9 0 9 11 2 11 2 15 13 0 7 0 9 2
57 13 15 15 0 1 0 2 0 9 1 11 1 10 9 2 13 3 1 10 9 1 9 1 0 9 2 15 13 9 2 0 3 1 10 9 0 9 7 3 3 0 9 0 9 2 15 13 1 0 9 2 7 13 0 0 9 2
29 0 9 0 9 13 9 13 9 9 12 2 12 2 12 1 0 9 2 10 9 13 0 2 16 13 1 0 9 2
21 0 2 9 3 3 13 0 11 14 1 11 2 9 15 13 1 0 9 1 11 2
18 9 0 2 9 4 13 9 11 2 11 2 7 9 0 9 1 11 2
24 9 9 1 9 2 12 3 1 11 2 16 1 11 13 0 9 2 13 1 9 0 11 3 2
32 11 2 11 13 0 9 7 9 1 9 12 1 0 9 9 1 9 12 7 9 12 2 3 9 9 13 1 0 9 1 11 2
94 11 2 11 14 3 9 13 1 9 1 0 0 2 2 0 9 1 11 1 9 2 3 3 13 9 0 9 1 11 12 1 10 9 9 2 9 9 2 11 3 3 13 1 9 9 11 1 9 9 9 12 2 12 2 12 3 1 11 2 3 1 9 1 9 12 1 11 2 11 2 11 7 11 7 3 13 10 0 7 0 9 2 7 0 9 2 15 13 1 9 11 9 11 2
70 13 0 13 1 9 0 9 2 13 3 3 9 0 9 1 12 2 12 2 12 2 7 13 0 13 10 9 2 0 10 9 1 9 1 9 0 9 11 2 11 2 3 13 9 1 9 1 0 9 2 15 4 13 0 1 9 1 12 2 12 2 12 7 7 7 1 9 0 9 2
11 1 9 9 2 9 2 11 2 11 2 11
2 0 9
26 9 13 2 9 13 1 9 2 9 15 13 1 9 0 9 7 3 15 13 15 0 9 1 0 9 2
8 3 13 9 2 3 13 9 2
6 3 10 0 9 13 2
16 3 15 13 3 2 0 9 15 13 2 9 9 13 2 13 2
5 3 9 13 9 2
12 1 9 1 9 2 3 0 9 2 13 0 2
14 9 3 13 2 15 14 2 13 15 3 2 15 13 2
23 15 13 3 1 9 2 9 7 9 2 9 7 9 2 9 2 9 2 9 2 15 13 2
6 14 9 2 9 13 2
4 15 15 13 2
18 3 15 13 2 3 1 15 4 13 0 9 1 0 9 0 1 9 2
18 1 9 3 7 0 9 0 3 2 16 13 0 9 1 9 15 0 2
33 13 2 14 3 2 13 15 9 2 13 9 1 15 2 15 13 1 15 2 15 2 15 13 3 16 15 2 9 7 9 2 9 2
21 7 9 0 3 13 3 2 16 0 9 4 13 0 9 9 1 11 2 10 9 2
9 1 9 11 11 2 12 9 2 11
18 9 11 11 15 13 1 9 0 9 1 9 10 9 1 9 11 11 11
2 9 11
4 11 1 9 13
2 11 2
19 0 9 7 9 1 9 11 11 13 1 0 9 13 10 0 0 0 9 2
9 13 15 3 1 0 9 1 11 2
2 11 13
2 11 2
21 9 9 11 11 11 13 0 0 9 1 0 9 9 9 11 11 2 11 0 11 2
6 13 15 3 9 11 2
17 13 13 2 1 10 9 15 13 2 16 3 13 0 9 0 9 2
15 10 9 13 1 9 15 2 16 0 9 13 15 9 11 2
3 11 15 13
2 11 2
16 0 9 0 0 9 11 11 4 13 1 0 9 13 9 11 2
25 3 15 15 13 9 9 9 11 11 2 15 13 2 16 11 13 9 10 9 2 16 13 11 11 2
7 9 1 11 1 9 9 11
5 11 2 11 2 2
30 9 0 9 1 0 0 9 7 9 11 13 1 9 9 11 11 11 2 15 4 0 9 13 13 1 9 11 11 11 2
24 9 0 9 2 13 1 9 9 12 2 9 13 9 11 11 11 2 7 11 1 15 9 13 2
26 9 9 2 15 13 0 0 9 7 0 0 9 11 2 13 14 9 9 11 2 11 1 11 2 11 2
19 1 15 9 11 13 9 1 9 9 2 15 9 0 9 13 1 0 9 2
39 4 15 13 13 3 2 16 4 15 13 0 10 9 7 10 9 2 15 4 3 13 4 0 9 13 2 13 11 2 11 9 9 2 15 4 1 11 13 2
20 14 1 9 10 0 9 15 13 2 16 13 1 0 9 0 9 13 7 3 2
4 11 14 11 13
16 1 9 11 1 9 9 15 1 10 9 13 10 9 11 11 2
5 3 4 13 9 2
9 13 15 0 9 14 1 9 11 2
21 1 15 15 13 9 2 15 4 13 3 1 9 9 2 16 9 1 15 3 13 2
10 3 3 2 15 13 3 0 0 9 2
8 1 15 13 13 1 0 9 2
7 14 3 0 2 7 0 2
16 13 2 14 15 0 9 2 3 13 2 16 11 13 1 9 2
10 13 13 2 13 0 0 9 1 9 2
10 13 9 2 16 9 3 13 3 0 2
10 13 1 9 13 15 1 9 1 9 2
22 16 15 13 9 9 2 13 12 9 2 7 3 1 9 9 13 2 15 3 2 2 2
7 1 10 9 13 0 9 2
3 3 0 2
27 3 4 13 3 13 2 7 3 4 15 13 13 1 0 9 16 15 13 1 0 9 1 11 7 13 15 2
30 16 13 13 1 9 2 15 13 1 0 9 12 9 2 12 9 9 2 3 15 13 9 9 7 7 0 9 1 11 2
20 1 9 15 13 9 2 16 1 9 9 1 9 9 1 9 11 13 2 2 2
10 3 4 15 15 9 9 13 2 2 2
18 15 4 15 0 9 13 1 9 2 15 13 14 9 7 1 15 13 2
17 11 13 3 0 2 7 3 15 1 15 13 13 10 0 0 9 2
16 3 15 13 9 2 3 9 7 9 2 15 4 13 0 9 2
3 2 11 2
3 1 0 9
18 11 11 1 0 11 15 3 13 13 1 11 2 7 13 1 0 9 2
20 9 12 2 9 12 2 9 0 9 2 11 15 13 3 1 9 1 12 9 2
23 11 11 2 0 0 9 1 11 13 1 9 1 11 7 3 1 0 0 9 13 13 13 2
5 2 11 2 11 2
5 11 13 1 0 9
16 9 9 13 9 2 9 3 13 9 2 13 9 11 9 11 11
4 11 11 2 11
12 0 9 13 9 0 9 11 9 11 1 9 2
28 3 4 15 3 3 13 2 13 13 1 9 2 7 15 15 13 0 9 2 15 9 9 13 1 0 9 9 2
33 1 15 4 13 13 0 9 14 1 9 0 9 9 1 9 1 9 2 16 9 15 13 13 0 9 1 0 9 1 0 0 9 2
46 15 13 3 1 9 2 3 15 9 1 0 9 11 13 2 16 1 0 9 4 13 0 0 9 16 1 15 0 2 15 3 3 1 9 1 9 13 0 9 9 2 12 2 12 2 2
14 3 3 7 9 2 15 13 1 2 13 13 1 9 2
22 16 3 1 9 9 13 9 13 2 9 15 13 2 16 15 15 13 2 15 3 13 2
66 13 4 1 10 9 3 1 9 9 7 7 16 4 3 1 12 9 13 1 0 9 0 2 13 4 1 9 3 2 16 1 9 12 2 12 2 3 4 15 13 1 0 7 0 9 2 13 9 11 11 2 9 9 7 3 1 11 2 11 7 11 12 1 9 9 2
10 13 15 1 15 1 0 9 7 0 2
12 16 13 9 2 3 13 2 1 15 4 13 2
31 1 15 2 15 13 9 2 15 1 9 13 9 2 15 15 13 2 3 3 13 1 10 9 1 15 9 12 9 2 2 2
36 9 3 13 2 16 15 0 9 13 3 2 16 13 0 9 1 9 1 0 9 2 3 1 12 9 1 9 1 0 9 14 1 12 1 0 2
21 1 9 9 11 11 9 1 9 3 1 0 9 13 9 2 16 13 0 0 9 2
21 1 9 3 13 1 9 2 16 16 15 13 13 2 13 3 1 0 9 1 11 2
25 9 11 9 11 15 7 13 2 16 15 13 1 9 3 13 0 9 0 9 2 0 3 1 9 2
26 15 15 7 13 2 7 1 9 15 13 3 12 1 12 9 9 2 0 13 1 10 9 1 9 2 2
6 13 15 3 15 13 2
7 13 4 15 13 1 9 2
12 13 4 7 15 13 1 2 13 9 11 11 2
20 3 13 2 13 15 3 9 11 2 15 15 13 1 9 13 3 1 0 9 2
7 0 7 13 13 1 15 2
13 1 9 9 13 12 9 7 15 13 13 0 9 2
5 1 0 9 13 2
14 1 12 9 13 0 9 13 1 9 0 9 1 11 2
26 1 0 9 11 3 13 9 7 3 2 3 1 9 2 13 1 0 9 9 9 11 0 9 0 11 2
23 11 15 13 13 2 9 11 2 15 15 3 13 13 1 11 1 0 9 2 13 0 3 2
29 9 13 13 2 7 1 9 0 0 9 4 13 1 11 9 10 0 9 2 13 15 13 9 0 9 11 11 11 2
19 9 0 9 3 13 1 9 2 3 13 1 9 0 9 0 9 11 9 2
12 1 15 4 13 9 13 10 9 1 0 9 2
10 13 12 0 9 9 2 13 11 11 2
17 7 15 9 13 15 2 7 13 0 9 2 7 13 1 10 9 2
19 15 3 13 2 16 9 13 1 9 2 16 4 15 13 9 1 15 13 2
24 13 15 15 3 9 2 16 3 15 13 9 1 9 2 3 3 4 15 1 15 13 13 3 2
15 15 13 2 16 16 4 15 13 2 16 1 11 13 11 2
12 9 15 13 2 3 15 13 14 1 0 9 2
14 9 10 9 13 13 9 2 3 15 15 13 3 13 2
7 10 9 13 7 1 9 2
20 9 2 3 15 13 9 14 1 15 2 16 15 9 13 9 2 3 3 13 2
11 9 13 0 9 7 9 10 9 13 9 2
10 15 13 9 7 9 15 10 9 13 2
2 0 9
12 9 9 1 11 2 9 9 2 12 9 2 2
1 9
2 9 11
12 2 9 0 9 1 9 2 3 0 9 13 2
4 9 9 11 2
3 0 9 2
19 11 11 2 11 9 12 2 12 2 12 2 12 2 2 0 9 0 9 2
10 9 2 12 2 11 2 12 2 11 2
1 9
42 0 9 2 12 2 9 2 11 11 2 11 11 12 2 12 2 12 2 12 2 12 2 12 2 12 2 12 2 2 9 2 11 12 2 11 2 11 2 11 2 11 2
1 9
5 0 9 1 11 2
5 0 11 2 12 2
3 11 11 2
4 11 2 12 2
2 11 2
4 11 2 12 2
3 11 11 2
4 11 2 12 2
2 11 2
5 11 11 2 12 2
3 0 11 2
5 11 11 2 12 2
2 11 2
5 11 9 2 12 2
2 9 2
4 15 4 13 2
43 12 2 9 2 0 12 2 1 12 2 9 12 9 12 9 2 1 12 2 13 12 9 12 9 2 1 12 2 13 12 9 12 9 7 1 12 2 13 12 9 12 9 2
39 9 2 1 12 2 7 12 2 9 13 9 2 1 12 2 13 12 9 12 9 2 1 12 2 13 12 9 12 9 7 1 12 2 13 12 9 12 9 2
4 9 0 0 9
16 11 11 13 1 9 0 11 1 9 11 12 2 12 7 13 3
7 0 9 11 1 11 11 11
19 3 1 0 11 13 11 11 0 0 9 2 15 13 1 9 0 0 9 2
15 3 1 9 9 11 11 15 0 9 11 1 11 13 3 2
24 1 0 9 3 0 13 1 0 9 11 2 0 9 2 7 1 9 12 2 12 1 0 9 2
21 3 15 13 13 2 3 13 16 11 2 13 16 9 1 9 1 9 0 9 11 2
15 10 9 15 13 10 9 1 9 7 1 0 9 13 3 2
20 9 11 13 3 1 0 9 9 3 1 9 11 2 3 13 9 13 0 9 2
11 1 0 9 15 11 13 14 1 9 11 2
9 1 0 9 13 9 16 1 9 2
32 1 12 2 9 15 0 9 1 0 9 13 13 9 11 7 1 9 3 13 9 2 15 13 2 16 4 11 13 9 9 11 2
14 16 15 11 13 13 3 9 2 16 4 13 10 9 2
24 3 15 1 0 9 13 1 12 2 9 1 0 9 11 7 10 0 0 9 13 9 1 9 2
16 11 15 3 13 1 9 11 2 15 13 1 9 1 0 9 2
12 1 9 13 9 11 2 15 13 1 12 9 2
21 11 13 1 0 0 9 0 11 7 15 1 9 1 9 9 13 0 9 11 9 2
12 9 11 13 7 15 13 2 16 4 11 13 2
25 1 0 9 13 11 1 9 13 3 0 11 7 1 12 9 13 9 1 12 2 12 1 10 9 2
33 0 9 13 1 9 9 7 13 15 13 1 12 2 9 2 3 0 11 13 9 2 11 15 13 1 0 11 2 15 0 9 13 2
22 9 3 13 11 9 7 11 3 9 13 0 0 9 7 13 0 12 9 11 1 9 2
10 15 3 12 9 3 13 1 11 11 2
24 1 1 15 2 16 0 9 13 11 12 2 12 2 13 4 1 9 13 12 9 7 15 13 2
19 15 13 1 10 9 2 16 3 1 12 2 9 13 3 11 9 1 9 2
17 1 9 9 1 12 9 15 9 13 0 9 14 1 9 1 9 2
19 3 9 11 13 9 1 9 11 2 15 13 9 0 7 4 13 1 9 2
12 0 9 13 9 3 9 11 2 12 2 12 2
9 3 13 7 9 11 7 11 13 2
29 9 2 12 2 2 12 2 11 2 12 2 11 1 9 2 12 2 11 2 12 2 11 2 12 2 11 1 9 2
12 9 2 11 2 11 2 11 2 15 11 2 2
4 9 2 11 2
4 9 2 12 2
6 9 2 12 2 12 2
3 9 1 9
15 11 11 2 9 11 2 13 13 9 2 7 3 9 9 2
20 13 4 2 16 13 9 2 16 4 13 0 9 2 7 0 9 13 3 3 2
6 3 15 13 0 11 2
22 11 11 2 9 11 11 2 13 15 15 13 3 0 9 2 15 4 13 1 9 13 2
22 9 1 9 15 13 14 9 11 2 15 13 1 0 9 7 1 9 9 13 3 13 2
13 0 9 7 0 9 4 15 13 15 0 9 2 2
28 9 11 11 2 3 1 0 9 4 15 13 9 12 9 2 1 15 15 12 13 13 3 1 0 9 1 11 2
6 12 1 15 13 11 2
11 3 3 13 1 9 2 7 4 13 9 2
24 11 11 2 9 0 9 2 1 9 10 9 4 1 9 13 9 2 7 4 3 13 0 9 2
26 1 9 15 7 15 13 7 1 9 2 3 4 13 1 0 9 2 3 4 13 2 16 15 13 9 2
5 11 13 1 9 9
6 0 11 2 11 2 2
17 1 0 11 3 12 9 3 13 11 11 2 12 2 9 11 2 2
47 7 15 3 15 2 16 1 0 9 1 11 1 9 1 11 0 0 9 3 13 2 16 9 13 10 9 13 2 16 13 10 9 1 0 0 2 12 2 12 2 2 12 2 12 2 2 2
22 13 4 9 1 9 7 13 3 1 10 9 2 16 15 9 13 2 16 4 15 13 2
18 7 15 13 13 3 2 1 9 2 7 1 12 9 2 13 3 11 2
17 3 1 9 1 11 3 9 0 0 12 3 13 2 13 4 0 2
17 13 4 15 2 16 4 15 13 2 7 13 15 7 13 15 9 2
3 9 1 9
37 9 2 12 2 9 2 9 2 12 2 9 2 12 9 2 2 11 2 11 2 11 11 2 11 2 11 1 11 2 11 2 0 2 9 2 11 2
39 9 2 12 2 11 2 11 2 11 11 2 0 9 2 11 9 2 11 2 11 9 2 11 2 12 2 11 2 0 11 2 11 2 11 2 11 2 11 2
16 9 2 0 0 9 1 11 2 12 9 2 2 11 2 11 2
44 9 2 12 2 9 2 9 2 12 2 9 2 12 9 2 2 11 2 11 2 12 2 11 2 0 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2
12 11 2 12 2 11 2 11 2 11 2 11 2
9 9 2 12 2 11 2 11 9 2
16 9 2 0 0 9 1 11 2 12 9 2 2 11 2 11 2
5 0 9 1 12 9
2 1 11
6 0 9 1 0 0 9
2 11 2
22 9 0 9 2 11 13 12 2 9 1 12 9 2 1 11 0 0 9 9 11 12 2
16 0 9 11 2 11 3 13 1 0 9 11 11 1 12 9 2
32 9 13 3 14 1 12 2 9 2 3 9 13 9 11 2 11 7 11 2 11 2 13 1 11 9 0 9 11 11 11 11 2
16 9 11 3 1 0 0 9 13 9 11 11 1 9 11 11 2
6 9 13 0 0 9 2
24 13 4 9 1 9 2 16 1 9 0 9 0 9 0 9 11 11 13 9 11 1 0 9 2
15 13 1 9 1 9 2 3 15 13 9 9 0 1 9 2
8 12 9 13 1 11 0 9 2
11 1 11 11 15 13 11 11 7 11 11 2
9 3 0 9 13 13 1 0 9 2
15 9 11 11 11 13 3 9 1 9 11 9 7 11 11 2
14 11 13 1 0 9 2 1 9 2 15 13 0 9 2
14 11 13 13 1 0 9 9 9 9 7 15 13 9 2
9 1 9 9 2 0 9 1 9 2
24 1 9 12 15 3 13 0 9 1 9 1 9 9 2 15 13 1 11 2 13 11 2 11 2
14 13 2 16 9 9 11 12 1 11 13 12 0 9 2
11 0 12 2 0 12 7 0 9 12 9 2
10 9 1 9 9 13 3 12 9 9 2
11 9 1 9 1 0 9 13 11 7 11 2
14 13 4 12 9 2 12 0 9 7 9 4 15 13 2
19 13 15 9 1 0 11 2 7 10 15 13 3 13 2 13 11 2 11 2
3 12 9 3
9 11 13 12 9 9 12 1 12 9
2 11 2
16 12 0 9 1 0 9 1 9 0 9 9 13 11 11 11 2
27 0 9 1 0 9 13 12 9 0 9 1 9 12 2 12 2 15 13 1 12 10 0 9 1 11 12 2
26 3 15 13 9 9 1 12 9 12 2 12 2 15 13 0 1 12 9 16 10 0 9 1 9 12 2
8 11 13 9 12 1 9 9 2
10 0 11 13 1 9 3 0 0 9 2
14 1 0 0 9 1 9 13 3 3 16 3 11 11 2
14 13 3 0 9 2 15 13 10 9 3 1 12 9 2
13 12 9 13 3 3 7 13 13 2 16 14 3 2
12 1 15 13 1 0 9 3 12 9 0 9 2
18 11 3 16 9 0 0 9 13 13 0 14 1 0 9 12 1 11 2
14 1 0 9 13 1 9 9 11 11 9 12 2 12 2
21 1 0 9 9 0 0 9 13 0 11 11 11 9 12 2 12 11 11 1 11 2
17 11 13 7 13 13 1 10 9 0 0 9 1 9 1 9 12 2
15 13 13 2 10 9 15 1 9 1 12 9 1 9 13 2
11 3 4 13 13 3 0 2 13 0 11 2
10 9 0 9 1 12 9 0 2 9 2
3 3 3 11
7 7 1 9 15 0 9 13
2 11 2
24 0 9 11 11 15 13 1 0 9 1 11 9 9 1 0 9 2 15 13 1 0 9 9 2
31 0 0 0 9 1 9 7 9 9 1 0 9 1 11 13 3 3 7 1 0 1 9 2 0 11 11 2 13 12 9 2
24 1 12 0 15 13 12 9 2 7 1 0 9 15 13 13 0 0 9 9 11 11 1 11 2
20 9 0 9 11 11 7 11 11 13 13 0 9 1 9 9 11 1 0 9 2
13 13 3 1 9 10 9 2 7 1 0 15 13 2
43 16 0 1 0 9 2 1 0 9 0 2 13 1 3 0 9 2 12 9 2 11 7 1 0 0 9 1 12 2 9 15 13 0 9 2 11 13 1 15 1 12 9 2
29 1 9 15 13 11 9 1 12 2 12 2 15 1 10 9 13 9 2 7 15 9 13 3 1 9 7 1 9 2
10 11 1 9 13 9 1 9 0 9 2
9 3 1 0 9 13 13 1 9 2
27 9 13 3 1 0 9 1 9 11 2 7 15 13 0 9 7 13 2 16 10 0 9 1 9 13 0 2
17 3 13 11 1 11 2 7 1 0 9 13 1 11 1 12 9 2
24 1 9 0 9 0 9 13 0 9 0 0 11 10 9 11 7 0 9 15 13 1 0 9 2
13 1 9 11 2 11 13 2 13 4 14 10 9 2
15 13 0 1 15 2 16 4 13 15 2 9 3 15 13 2
15 11 2 11 2 13 4 0 9 2 14 4 13 3 0 2
15 12 9 1 9 15 13 9 7 1 15 9 9 13 3 2
9 10 0 9 15 7 3 3 13 2
12 0 11 11 1 11 13 0 9 1 9 9 2
21 1 12 9 13 0 9 1 12 2 12 9 2 15 13 9 3 12 9 2 9 2
14 0 1 9 11 11 1 11 13 1 15 1 12 9 2
24 10 0 9 1 9 10 9 1 9 13 9 0 9 11 11 2 15 13 0 9 1 9 9 2
23 9 0 11 13 0 2 15 15 13 1 0 9 2 16 9 13 3 3 7 13 14 0 2
21 0 9 9 11 13 9 1 12 2 12 9 2 0 16 9 7 13 12 2 9 2
21 0 9 0 0 9 13 3 3 16 12 15 0 9 0 9 1 0 9 11 11 2
33 1 9 9 9 1 9 4 1 0 9 13 1 9 12 2 9 11 1 12 10 9 2 15 13 0 9 9 7 9 0 9 11 2
17 0 9 2 15 13 1 9 0 0 9 2 13 9 11 1 0 2
22 0 0 9 13 0 13 16 9 2 15 3 13 2 3 11 13 2 13 1 10 9 2
2 11 2
2 9 11
6 1 9 11 14 0 9
12 16 9 13 1 9 0 9 2 13 13 3 15
5 11 2 11 2 2
24 13 0 9 13 9 9 1 9 9 0 9 11 11 1 9 2 3 3 13 13 9 1 9 2
21 11 15 13 1 9 1 9 11 11 2 0 9 9 0 9 1 11 1 9 12 2
46 11 4 13 1 9 12 16 9 9 1 9 9 0 9 2 16 1 9 1 9 12 1 9 12 3 1 10 9 11 11 3 13 9 1 9 1 11 2 16 15 13 0 9 0 9 2
8 15 9 0 0 9 1 11 2
23 1 9 9 0 9 7 3 1 0 0 9 4 13 11 1 12 9 7 11 1 12 9 2
34 1 11 0 0 9 2 13 1 15 3 2 9 2 11 11 2 7 1 0 9 0 9 13 2 16 9 1 15 13 0 9 0 9 2
29 9 13 1 0 0 9 2 16 1 9 4 3 13 7 1 0 9 9 1 12 1 12 9 1 0 9 1 9 2
18 9 13 2 16 0 9 7 0 9 3 13 2 13 15 3 9 9 2
23 0 9 11 7 11 13 0 0 9 2 15 13 0 9 1 9 2 15 4 3 3 13 2
25 9 9 13 2 16 7 16 4 13 1 9 0 9 2 9 1 9 9 1 9 9 3 4 13 2
22 11 1 9 1 10 9 13 1 0 7 9 13 7 3 3 13 1 12 9 0 9 2
15 7 16 13 13 2 16 9 9 1 9 9 1 9 13 2
15 1 9 13 3 0 0 0 9 1 11 2 15 9 13 2
44 11 13 0 2 9 0 7 9 0 9 1 9 11 13 0 9 2 16 13 1 3 0 9 2 3 4 9 10 9 1 9 13 1 9 2 15 1 15 15 13 7 15 13 2
12 11 2 11 13 3 3 1 11 1 9 11 2
8 0 9 1 9 11 13 0 9
10 11 11 2 11 2 9 11 11 2 2
13 9 1 3 0 9 11 11 7 11 13 0 9 2
26 3 4 15 13 1 9 1 0 9 2 3 4 13 0 9 7 3 13 0 2 13 9 11 11 11 2
12 9 13 0 9 1 15 2 16 13 1 11 2
9 0 9 15 13 7 3 15 13 2
8 13 0 2 16 15 3 13 2
10 0 9 4 10 13 7 1 11 11 2
8 0 9 15 7 13 1 11 2
26 0 0 9 11 11 2 2 9 9 0 9 2 15 13 1 9 1 9 2 16 15 13 1 11 11 2
18 10 9 13 1 9 9 10 9 2 16 4 0 9 13 0 0 9 2
12 9 0 9 1 11 11 13 3 15 0 9 2
18 3 1 12 9 15 15 3 13 2 13 9 1 0 9 0 0 9 2
16 3 1 9 2 16 15 1 0 9 13 7 1 11 13 3 2
19 15 2 16 4 13 0 9 2 4 13 10 9 14 1 11 7 0 11 2
8 1 10 9 13 14 12 9 0
5 11 2 11 2 2
14 1 9 13 1 9 0 9 14 12 9 1 12 0 2
20 0 9 13 2 16 1 9 9 13 1 9 3 12 0 2 3 3 12 9 2
13 13 1 15 11 0 9 0 9 0 9 11 11 2
25 0 9 13 9 2 16 4 15 0 9 0 13 3 1 12 9 2 3 13 15 0 1 0 9 2
20 9 7 13 3 3 9 13 9 9 7 13 3 1 9 2 16 15 9 13 2
23 1 0 9 15 13 0 0 9 1 9 12 9 1 9 9 3 1 12 1 12 9 3 2
11 9 11 11 2 1 0 9 15 0 9 13
5 11 2 11 2 2
32 1 9 13 9 7 13 15 1 15 0 9 2 2 2 13 15 9 2 13 1 0 11 9 0 9 9 11 11 2 11 2 2
9 9 13 2 16 0 9 9 13 2
15 13 3 1 9 0 9 9 1 10 9 1 11 7 11 2
17 10 9 1 15 13 9 7 13 15 1 9 9 9 1 0 9 2
28 9 0 9 11 11 15 1 15 13 2 16 9 1 9 3 13 2 13 7 2 16 15 1 15 13 0 9 2
10 9 1 9 1 15 13 9 1 9 2
11 9 13 9 1 9 1 0 2 13 11 2
18 1 9 9 0 9 13 0 9 9 1 9 2 1 9 7 0 9 2
12 9 15 13 9 0 9 7 0 9 1 9 2
21 14 3 13 1 12 2 9 1 9 12 9 2 3 1 0 9 2 7 12 9 2
19 1 9 9 7 9 12 9 2 3 0 9 2 7 12 9 2 9 2 2
18 9 15 1 9 13 9 2 15 9 3 13 2 3 16 13 4 13 2
8 9 1 9 14 13 9 9 2
12 9 2 15 15 3 13 2 13 3 0 9 2
8 1 0 9 1 9 11 13 2
14 1 10 9 1 15 13 1 9 9 1 9 7 0 2
26 9 1 15 13 9 2 1 15 15 1 15 4 13 13 15 2 15 15 13 2 16 15 15 13 9 2
16 13 15 13 15 2 16 4 15 9 9 13 9 1 9 9 2
17 7 7 15 11 13 0 9 0 9 2 15 15 13 13 1 9 2
9 9 0 9 13 9 1 0 9 2
7 9 13 14 1 10 9 2
18 16 13 0 7 3 0 9 2 13 10 9 13 9 7 13 1 9 2
9 1 0 9 15 7 9 13 3 2
15 16 4 1 10 9 13 9 2 9 4 1 11 3 13 2
4 1 9 13 11
37 1 0 9 13 9 2 16 15 1 9 15 2 15 15 13 1 9 2 13 1 3 0 9 2 3 15 1 0 9 13 9 7 9 3 0 9 2
21 9 11 13 1 10 9 7 13 2 16 0 13 3 9 1 9 1 11 7 11 2
32 3 7 1 9 13 0 9 2 7 3 15 16 0 9 13 2 16 13 1 9 13 15 9 2 16 15 0 9 13 0 9 2
9 9 9 1 9 13 11 15 13 2
5 12 7 13 13 2
10 9 11 11 15 1 9 13 0 9 2
9 2 11 2 2 11 12 2 12 2
4 1 15 1 11
2 0 9
2 11 11
10 1 0 9 15 9 1 11 13 3 2
5 9 13 11 11 2
20 15 15 13 7 15 1 15 13 0 2 16 11 11 13 10 0 7 0 9 2
8 9 3 13 1 11 15 13 2
11 1 9 15 3 3 13 1 9 9 13 2
8 13 1 15 3 10 0 9 2
16 9 1 9 15 11 15 13 1 0 9 2 16 16 15 13 2
4 7 3 13 2
7 9 13 1 9 9 0 2
25 15 15 13 7 15 1 15 13 0 2 16 11 13 10 7 0 1 15 13 10 0 7 0 9 2
12 1 9 0 9 15 1 10 9 13 0 9 2
12 9 1 9 15 13 3 1 10 9 11 13 2
10 13 15 7 1 0 9 7 0 13 2
8 1 0 9 13 0 9 0 2
17 15 15 13 7 15 1 15 13 0 2 16 1 15 13 0 9 2
21 9 15 15 13 2 7 3 15 1 15 3 13 0 0 9 7 13 15 0 9 2
23 15 9 13 12 9 3 2 16 13 2 16 15 0 9 3 3 2 3 7 3 13 9 2
13 15 15 1 0 13 1 0 15 9 1 0 9 2
22 1 9 2 0 1 9 7 0 9 2 9 0 12 9 13 9 2 13 9 9 9 2
6 13 9 0 9 9 2
10 0 13 0 13 15 1 10 9 9 2
10 0 0 9 14 0 13 9 1 9 2
10 1 9 9 9 3 13 7 13 9 2
6 15 13 7 14 9 2
6 1 0 15 9 13 2
13 9 1 9 3 1 9 13 2 16 13 0 9 2
9 1 9 4 13 15 12 0 9 2
4 13 7 9 2
18 3 15 1 9 13 1 9 12 9 7 12 9 9 9 1 9 9 2
35 3 13 0 0 9 2 1 0 9 15 3 14 13 9 13 2 16 4 1 0 0 9 13 1 0 9 12 9 2 15 4 13 7 13 2
17 1 9 0 0 9 15 3 13 13 9 7 13 15 1 9 13 2
21 3 3 7 4 1 9 1 9 13 2 16 9 11 13 9 9 3 16 3 3 2
20 10 9 13 3 0 9 7 10 0 9 1 9 4 3 13 13 0 7 9 2
9 1 15 13 0 7 9 13 9 2
3 15 13 2
25 9 15 3 1 0 9 9 13 10 9 2 9 15 1 9 13 9 7 9 2 15 0 3 13 2
18 0 9 0 9 13 0 9 2 3 9 1 9 1 9 13 1 9 2
7 9 15 1 9 13 13 2
8 9 9 15 9 13 9 11 2
6 9 2 9 1 9 9
2 11 11
11 0 13 0 7 3 0 2 0 3 0 2
13 1 0 9 13 13 2 16 0 9 13 9 9 2
22 0 9 2 0 9 9 2 9 9 7 9 2 9 0 9 2 9 2 9 2 2 2
14 15 2 15 13 9 2 13 7 13 2 3 3 13 2
3 1 15 2
28 9 2 0 15 0 9 7 0 9 2 13 1 10 9 1 10 0 9 2 1 15 0 9 3 13 0 9 2
14 3 3 4 3 13 2 16 12 9 9 13 0 9 2
31 0 15 13 3 1 0 9 2 3 2 9 9 7 9 0 9 2 0 9 13 3 1 9 0 1 9 7 1 0 9 2
10 3 13 2 3 13 9 2 3 9 2
18 0 9 13 2 13 2 13 9 2 3 13 7 13 9 1 9 9 2
35 0 13 9 3 2 13 15 0 9 7 13 15 13 16 9 2 0 15 1 9 2 13 9 9 13 2 1 9 13 2 13 0 0 9 2
25 9 1 9 1 15 13 2 16 1 9 10 9 13 0 0 9 13 2 7 3 0 9 9 13 2
23 13 3 2 16 0 9 9 13 3 3 13 1 9 15 2 16 15 13 15 1 0 9 2
14 0 9 15 3 1 9 13 3 3 9 9 7 9 2
17 3 13 0 9 10 0 9 2 3 0 9 1 9 1 9 9 2
11 0 9 7 9 13 2 3 13 0 9 2
19 9 9 13 1 15 2 3 3 15 13 13 0 9 1 9 1 0 9 2
18 9 7 9 15 13 0 9 2 15 0 9 13 9 1 0 9 9 2
18 13 15 2 16 9 0 9 3 13 13 2 1 10 9 3 13 0 2
17 16 4 15 9 13 1 9 2 4 1 9 13 9 9 7 9 2
14 9 13 16 9 2 0 0 9 9 2 0 9 9 2
26 13 0 0 9 2 9 2 9 2 9 2 0 9 2 9 9 2 9 0 9 9 2 9 7 9 2
19 13 14 1 15 2 3 15 10 0 9 3 1 9 9 7 9 13 13 2
8 0 11 13 9 1 0 0 9
2 9 9
2 11 11
6 10 9 13 0 9 2
23 0 11 13 11 11 3 1 0 0 9 2 1 0 9 7 1 9 2 15 13 10 9 2
20 9 13 13 1 3 0 2 7 11 15 1 15 13 7 9 2 1 0 9 2
55 13 15 1 9 3 0 2 11 11 2 11 2 11 11 7 0 9 11 11 2 7 16 4 13 9 9 11 11 2 0 3 1 9 1 10 9 16 11 7 11 2 2 13 4 13 9 13 1 0 0 9 3 15 0 2
30 0 9 13 0 9 1 0 9 9 2 7 3 13 9 7 0 9 7 3 13 1 0 9 2 1 9 1 0 9 2
56 3 0 9 2 7 10 0 9 16 9 1 11 11 2 0 1 0 9 2 13 3 16 9 2 15 3 13 9 15 2 16 13 10 0 9 7 0 9 2 16 13 1 0 9 0 9 3 0 9 2 3 9 16 9 9 2
15 0 11 7 13 0 9 0 0 9 2 7 10 0 9 2
21 3 1 10 0 10 9 11 13 10 0 9 2 15 4 3 13 3 0 7 0 2
26 9 15 13 1 9 2 1 9 11 2 3 15 1 9 13 2 16 4 15 3 13 9 2 0 9 2
24 11 2 1 9 11 2 15 13 1 11 2 13 15 15 7 1 9 10 9 15 13 16 9 2
14 13 2 16 10 9 2 10 9 7 9 13 3 3 2
32 11 15 13 1 10 0 9 11 2 11 2 2 15 3 13 0 9 2 7 3 13 3 2 0 9 2 9 7 9 1 9 2
25 11 15 15 3 9 13 13 2 3 13 13 9 2 3 1 0 9 13 0 11 1 10 0 9 2
33 9 2 1 9 1 10 0 9 2 15 3 13 3 2 3 13 9 1 9 2 1 9 0 9 3 1 0 9 13 10 9 9 2
28 13 7 0 2 16 15 9 15 10 0 7 1 0 0 9 7 1 0 13 2 3 15 13 1 10 0 9 2
13 1 9 10 0 9 1 0 9 15 13 15 13 2
19 0 11 3 13 0 9 10 9 3 3 2 16 15 13 13 1 9 9 2
50 3 0 9 2 1 0 0 9 1 11 2 3 15 3 13 2 13 9 1 0 9 2 1 11 4 13 1 0 9 7 16 15 13 9 11 11 2 13 2 16 15 13 1 9 2 15 13 0 13 2
28 9 0 11 13 2 16 4 11 1 0 0 9 2 7 1 0 9 2 7 1 10 9 13 9 2 12 2 2
25 3 3 9 0 9 13 1 9 7 0 9 9 2 13 2 16 9 7 9 13 0 3 1 9 2
9 0 0 9 15 13 1 0 9 2
11 13 11 12 1 9 12 2 9 1 12 2
4 16 13 0 9
2 11 11
17 11 11 2 11 2 11 11 2 11 11 2 11 11 2 11 11 2
13 15 15 13 16 9 2 15 13 0 9 9 9 2
24 3 13 3 0 9 2 3 15 13 14 9 13 9 3 16 3 2 7 0 15 13 0 9 2
61 13 13 0 9 10 9 7 0 9 2 13 1 9 0 9 9 2 13 0 0 9 7 13 15 0 9 1 9 7 9 2 9 9 7 3 0 7 0 9 1 0 0 9 2 2 13 0 0 9 2 16 13 9 9 1 9 0 7 0 9 2
27 13 1 9 7 13 15 0 9 2 0 0 9 15 13 0 9 7 3 13 0 9 2 15 13 0 9 2
27 13 0 9 2 13 1 9 3 0 9 2 15 15 7 3 3 13 9 2 7 13 15 14 9 0 2 2
27 13 0 13 9 9 1 9 0 9 2 13 15 3 1 9 12 2 14 3 2 1 9 11 2 3 2 2
7 3 15 9 13 0 9 2
33 0 0 9 11 3 13 1 9 0 9 2 9 15 13 0 9 2 7 11 16 0 9 13 10 0 9 2 0 11 2 12 2 2
14 13 15 7 0 0 9 2 15 15 13 13 0 9 2
12 11 13 0 9 2 1 15 13 0 10 9 2
20 0 9 0 0 9 13 7 0 9 2 16 4 13 9 3 2 11 7 11 2
41 1 9 7 3 14 12 0 9 13 10 9 9 2 15 15 3 13 1 9 9 7 0 9 2 15 15 13 0 2 1 9 1 9 2 11 2 10 9 7 0 2
29 3 13 9 9 2 1 9 12 15 13 12 2 1 9 3 12 2 16 0 9 3 0 9 15 13 1 12 2 2
12 0 9 3 13 1 0 0 9 9 11 11 2
28 4 13 1 0 9 9 2 15 13 1 9 2 1 15 13 1 9 9 2 7 0 9 10 9 13 0 9 2
37 1 0 2 7 3 0 9 1 0 9 15 13 1 0 9 1 0 9 7 0 9 2 1 3 15 2 1 15 15 7 10 9 16 9 3 13 2
7 7 3 15 3 13 0 2
38 11 1 10 0 9 13 0 0 9 2 9 9 2 9 7 9 2 13 1 9 7 9 16 0 9 2 1 9 13 9 7 3 9 0 1 10 9 2
25 0 2 3 3 0 9 3 13 1 9 3 0 0 9 2 16 3 13 1 0 9 7 0 9 2
46 3 1 15 13 9 0 9 2 0 9 13 3 10 10 9 2 0 9 2 9 2 9 11 2 7 13 7 3 0 9 0 9 2 15 13 9 0 0 9 2 1 9 9 13 13 2
21 10 0 0 9 3 13 0 9 7 13 15 13 9 10 9 2 0 1 0 9 2
11 1 11 13 3 0 9 1 3 0 9 2
29 16 1 0 9 12 2 9 15 9 13 0 9 2 13 1 15 7 15 2 1 0 9 13 1 10 9 0 9 2
17 13 7 3 0 9 2 1 15 15 13 0 9 1 3 0 9 2
60 1 10 9 3 3 13 0 0 9 2 0 3 1 12 2 9 0 0 9 1 0 9 7 1 0 9 0 9 1 0 9 2 1 10 9 4 3 13 0 1 0 9 2 7 0 9 2 3 13 0 2 3 0 9 0 0 9 1 11 2
44 10 0 0 9 13 9 1 15 0 2 15 15 1 0 9 13 2 14 7 15 13 2 2 13 1 0 9 2 15 3 3 13 7 13 1 0 2 7 3 0 9 13 0 2
17 13 13 1 9 0 0 9 7 1 9 10 9 15 3 13 13 2
15 1 15 13 15 2 15 2 13 10 9 2 1 9 13 2
46 13 1 15 0 9 2 1 0 0 9 11 11 2 15 13 9 0 9 2 13 15 3 11 2 11 11 2 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 2 2
8 0 9 15 11 2 12 2 2
29 1 0 0 9 2 1 0 9 2 3 3 13 0 9 0 9 0 9 2 15 1 9 12 13 3 3 0 9 2
22 9 0 9 9 13 9 9 11 11 2 15 3 13 7 13 10 9 9 2 11 11 2
25 13 0 9 1 9 12 2 3 9 11 11 2 9 11 11 7 9 11 11 13 0 9 0 9 2
17 13 15 1 12 9 3 7 0 9 13 0 9 2 0 11 11 2
20 3 3 13 9 0 0 11 7 0 11 2 2 11 2 2 11 12 2 12 2
16 11 11 13 12 1 0 9 1 0 9 11 2 0 12 11 2
10 0 9 0 9 2 10 9 7 9 2
7 2 13 11 12 1 12 2
4 1 9 1 9
19 11 11 2 12 1 0 0 9 10 9 2 13 1 9 0 9 1 9 2
17 13 0 9 1 0 11 1 11 7 10 9 13 1 0 0 9 2
10 1 9 1 9 1 9 13 3 3 2
27 1 9 9 4 13 0 9 1 0 9 2 9 0 9 1 9 7 9 7 0 9 1 0 9 1 11 2
9 2 11 2 2 11 12 2 12 2
2 11 11
17 11 11 11 2 12 2 12 2 4 3 13 16 0 0 0 9 2
14 0 9 10 0 9 13 0 0 0 9 2 11 12 2
8 11 13 13 3 14 1 12 2
15 13 0 9 7 13 1 9 9 2 3 15 9 3 13 2
21 0 9 13 13 9 2 7 13 9 2 0 9 2 7 3 13 1 0 0 9 2
9 2 11 2 2 11 12 2 12 2
5 11 13 1 0 9
7 11 2 11 2 11 2 2
22 10 9 1 9 11 11 4 3 13 2 13 3 11 9 0 9 9 0 9 11 11 2
30 1 10 9 3 3 9 13 2 3 4 13 9 1 11 7 11 2 11 1 9 9 11 2 15 13 11 1 0 9 2
33 9 11 2 11 13 9 9 2 1 15 9 11 1 10 9 13 2 16 13 1 9 9 9 0 11 2 13 1 11 2 11 9 2
30 9 11 13 10 9 13 1 0 9 16 15 2 4 13 1 9 7 9 2 15 1 15 13 9 2 13 11 2 11 2
3 0 0 9
9 1 0 9 3 13 9 0 9 11
5 11 2 11 2 2
21 0 9 9 11 2 11 0 9 1 11 2 11 7 11 13 9 0 0 0 9 2
44 10 9 13 12 1 10 9 2 15 9 9 9 0 9 1 9 0 9 2 11 2 4 13 1 10 0 9 2 15 15 1 9 11 12 13 1 0 9 11 3 11 1 11 2
10 9 15 13 3 9 1 11 7 11 2
15 9 13 0 0 9 3 11 13 0 9 9 9 11 11 2
22 13 2 16 0 9 13 2 16 4 1 0 0 2 0 2 9 3 13 1 0 9 2
15 1 0 0 9 4 3 13 9 13 13 16 12 0 9 2
11 15 4 15 14 3 13 9 1 0 9 2
25 13 3 3 1 9 7 13 1 15 2 16 10 9 13 0 7 1 0 7 0 9 2 13 11 2
14 9 1 9 0 9 13 3 0 9 9 11 2 11 2
26 13 10 9 1 15 3 2 16 9 9 4 13 2 1 1 10 9 1 9 9 11 2 11 2 13 2
30 1 9 11 7 0 9 0 9 9 11 13 9 0 9 9 0 9 7 9 9 7 9 0 9 9 11 1 0 9 2
13 0 9 13 3 13 9 1 10 0 9 0 9 2
21 13 14 3 1 12 5 0 9 0 11 7 9 0 9 0 9 1 11 7 11 2
25 1 0 9 15 9 1 11 11 13 13 3 9 9 7 9 11 11 7 9 9 0 9 11 11 2
4 0 9 13 9
5 11 2 11 2 2
19 0 9 2 11 2 13 1 9 1 12 2 9 0 9 1 9 7 9 2
25 0 0 9 1 9 15 13 1 12 5 1 12 5 2 1 9 13 1 9 1 12 7 12 5 2
14 9 15 13 3 3 0 2 3 7 3 0 0 9 2
62 1 9 9 1 9 13 1 0 2 9 2 1 12 2 12 5 2 2 1 0 9 1 9 0 2 7 0 9 2 1 12 2 12 7 12 5 2 7 1 9 0 9 7 0 9 2 9 1 12 2 12 7 12 9 2 1 12 7 12 5 2 2
25 1 0 9 9 1 9 2 1 12 7 12 5 2 13 1 0 9 1 12 2 12 7 12 9 2
13 0 9 2 9 7 0 2 9 15 9 9 13 2
38 3 1 0 0 9 13 9 11 2 9 9 15 13 15 9 1 0 9 3 12 9 2 9 2 7 3 10 9 1 0 9 14 12 7 12 9 9 2
29 9 1 10 9 7 13 2 7 13 2 13 9 0 9 11 11 11 7 13 2 16 0 9 9 13 1 0 9 2
25 9 0 9 13 0 9 13 10 9 2 3 1 9 1 0 9 2 15 10 9 13 3 0 9 2
20 0 9 13 7 0 9 9 9 1 10 9 7 9 3 0 9 1 0 9 2
11 9 0 9 13 9 1 9 0 9 9 2
5 0 9 1 11 11
7 11 2 11 2 11 2 2
37 1 9 2 15 4 13 1 0 0 9 0 9 11 11 9 2 13 0 9 2 13 3 11 9 11 9 2 9 2 9 2 0 2 2 11 11 2
27 0 9 11 11 13 1 9 9 1 0 9 13 3 16 9 9 11 9 2 15 13 3 9 0 2 9 2
4 11 11 9 2
10 9 1 11 9 7 11 11 13 0 2
18 1 9 9 0 9 2 15 13 0 9 11 11 9 2 10 9 13 2
24 9 0 9 9 0 9 11 11 3 11 13 2 16 15 0 9 9 11 11 13 1 0 9 2
20 0 9 1 10 9 1 9 9 1 11 9 1 11 3 13 1 11 2 11 2
25 15 11 13 2 16 16 13 0 9 9 9 1 9 9 1 0 9 2 9 13 11 9 0 9 2
4 9 13 0 9
5 11 2 11 2 2
11 0 0 9 13 10 9 3 3 1 9 2
13 13 15 3 9 9 3 0 9 9 9 11 11 2
19 0 9 0 0 9 3 13 14 1 9 9 1 9 7 9 0 9 9 2
12 15 4 13 0 9 9 13 1 10 0 9 2
21 1 11 13 9 9 1 15 2 16 9 4 9 1 0 9 3 13 1 0 9 2
24 3 11 11 13 2 0 9 4 0 0 9 2 11 2 13 13 1 0 9 1 0 0 9 2
19 1 9 0 1 9 11 3 4 1 10 9 13 9 9 9 1 9 11 2
14 0 9 1 9 12 9 9 13 9 1 9 0 9 2
28 1 3 12 9 2 9 0 1 9 0 9 4 1 9 11 13 0 9 9 1 9 9 9 0 7 0 9 2
8 9 13 13 1 9 0 9 2
17 9 9 9 13 1 11 13 7 1 9 9 9 7 9 0 9 2
17 1 9 9 11 4 15 13 9 9 3 1 0 9 1 9 13 2
14 0 9 7 3 13 9 0 7 0 9 2 13 11 2
3 0 0 9
5 12 2 0 9 2
6 12 2 0 0 9 9
3 3 0 9
10 0 9 13 1 0 9 13 9 0 9
14 1 12 2 12 5 3 3 13 0 0 9 0 9 2
11 1 0 9 13 10 9 12 2 12 5 2
20 9 9 4 1 10 12 9 13 12 2 12 5 2 3 2 12 2 12 9 2
16 13 15 0 0 9 9 1 0 9 11 1 9 9 0 9 2
11 9 13 1 0 9 9 0 9 0 9 2
8 9 0 9 11 15 7 13 2
14 0 9 0 9 13 0 1 9 1 0 9 0 9 2
25 0 0 9 11 13 1 9 12 9 1 3 16 12 5 2 0 9 7 9 1 12 2 12 5 2
14 1 9 9 12 0 9 3 13 1 0 9 0 9 2
7 0 0 9 13 9 11 2
22 1 9 9 0 9 4 0 9 13 3 0 0 9 0 0 9 1 9 9 7 9 2
16 1 0 9 12 13 9 1 0 9 0 9 12 1 12 5 2
13 9 1 11 13 1 0 12 0 9 1 12 5 2
13 9 10 9 4 13 0 9 0 9 1 12 9 2
18 9 9 7 13 0 9 1 0 9 1 11 1 0 9 1 3 0 2
16 9 0 0 9 11 4 13 13 0 9 7 9 1 0 9 2
17 9 0 9 1 9 13 1 15 2 16 0 9 3 13 0 9 2
22 13 15 2 16 1 9 1 0 9 1 12 5 4 3 13 9 9 0 9 12 9 2
5 13 15 7 9 2
16 1 9 12 3 13 9 1 9 1 0 7 3 12 5 9 2
26 0 9 1 0 9 2 0 9 0 7 0 9 1 9 12 2 12 5 2 13 7 13 9 0 9 2
36 3 0 0 9 9 0 9 1 9 12 2 9 2 1 15 13 9 0 0 9 7 0 9 2 4 3 13 0 0 9 0 9 9 7 9 2
13 1 3 0 9 13 9 9 7 1 10 0 9 2
26 13 1 15 0 0 9 9 9 2 0 9 1 10 9 2 0 9 0 9 7 0 9 9 0 9 2
14 13 3 0 9 0 9 7 9 9 1 9 0 9 2
37 9 1 0 7 0 9 13 3 0 13 1 1 0 9 1 0 9 2 0 9 9 1 0 11 2 0 9 1 11 7 1 1 0 9 0 9 2
27 1 9 9 0 9 13 3 13 1 0 9 1 9 2 16 10 0 9 13 1 9 2 13 15 1 9 2
3 2 11 2
2 0 9
9 12 2 12 2 9 9 1 0 9
14 12 2 12 2 0 9 0 2 9 2 11 2 0 9
12 12 2 12 2 0 9 0 2 9 2 9 11
13 12 2 12 2 0 0 9 0 2 9 2 11 11
13 12 2 12 2 0 0 9 0 2 9 2 0 0
13 12 2 12 2 0 0 9 0 2 9 2 9 11
14 12 2 12 2 0 9 0 2 9 2 0 0 0 9
14 12 2 12 2 0 9 0 2 9 2 0 0 0 9
21 12 2 12 2 0 9 0 2 9 2 0 9 11 9 2 9 2 9 7 0 9
14 12 2 12 2 0 9 0 2 9 2 0 0 0 9
14 12 2 12 2 0 9 0 2 9 2 0 0 0 9
7 12 2 2 12 2 12 2
22 9 2 12 2 9 2 0 9 9 2 9 2 9 7 0 9 2 11 2 9 9 2
11 12 2 12 2 0 9 0 2 9 2 11
13 12 2 12 2 0 0 9 0 2 9 2 9 11
12 12 2 12 2 0 9 0 2 9 2 11 11
13 12 2 12 2 0 9 0 2 9 2 0 0 9
4 11 2 11 11
24 15 15 13 1 9 11 11 2 13 2 1 15 1 9 13 2 1 0 9 9 1 9 9 2
12 10 9 15 9 13 1 9 7 0 0 9 2
33 1 11 1 11 15 13 0 9 1 0 7 0 9 2 0 9 7 3 7 0 9 2 1 15 13 13 0 9 2 12 12 9 2
9 2 11 2 2 11 12 2 12 2
4 9 1 0 9
10 1 10 9 11 3 13 9 1 12 9
2 11 11
15 0 9 1 0 9 11 13 1 9 12 1 9 11 11 2
27 10 0 9 13 13 9 0 0 9 2 0 9 0 7 0 9 7 9 0 9 0 1 15 1 0 9 2
16 0 9 1 9 9 13 0 9 0 9 0 1 9 9 11 2
13 9 0 0 9 3 4 13 1 9 1 0 9 2
12 1 9 0 9 15 13 13 1 0 0 9 2
24 13 14 1 0 9 9 2 7 3 1 9 0 9 2 9 9 0 9 2 9 9 2 9 2
23 1 0 9 7 9 1 9 4 13 1 0 9 11 11 2 11 7 9 9 9 11 11 2
28 1 15 2 16 4 9 9 13 0 9 2 15 13 0 9 2 1 15 13 9 0 9 2 0 9 7 9 2
9 9 13 12 9 7 12 0 9 2
13 9 9 13 1 9 0 9 16 0 9 1 9 2
23 1 10 9 13 9 1 9 1 9 2 9 2 0 9 2 7 0 13 0 9 0 9 2
31 1 9 9 1 0 9 13 11 9 1 9 1 12 0 9 2 0 9 1 9 9 2 0 9 7 0 9 1 0 9 2
15 16 4 13 15 13 2 13 9 9 9 0 0 0 9 2
14 0 9 4 3 13 1 0 9 2 9 7 0 9 2
28 1 9 15 13 9 1 9 1 9 2 1 9 1 9 2 13 15 9 7 9 7 13 15 7 0 0 9 2
20 1 9 10 9 1 11 13 2 16 0 9 10 9 13 9 9 1 0 9 2
12 3 1 0 9 13 13 15 1 9 0 9 2
10 12 1 0 9 1 9 13 0 9 2
9 9 13 3 1 0 2 0 9 2
11 3 11 13 9 13 0 0 9 1 11 2
20 13 0 2 16 1 10 9 13 9 0 0 9 2 15 4 13 13 1 11 2
14 9 13 7 1 0 0 9 2 16 13 11 7 11 2
40 1 3 12 3 0 9 13 0 9 0 11 2 15 13 0 9 0 11 1 9 11 2 9 9 2 2 7 9 0 9 11 2 0 0 9 9 7 0 9 2
10 3 0 9 13 1 9 12 0 9 2
29 16 1 9 0 9 0 9 15 13 9 0 0 9 1 15 2 13 15 9 1 9 9 10 0 9 1 0 9 2
15 1 9 12 15 9 10 9 13 1 9 0 9 1 9 2
3 11 13 9
5 11 2 11 2 2
51 1 9 3 0 9 9 0 7 0 9 1 0 9 0 9 2 11 2 0 7 0 11 2 11 2 9 2 11 2 11 7 0 11 2 0 11 2 15 13 1 0 11 1 9 12 2 7 12 2 9 2
18 10 9 13 13 0 9 13 0 9 7 13 9 0 0 7 0 9 2
64 11 15 13 3 12 0 9 7 12 0 9 2 0 1 9 9 2 9 7 9 2 9 2 9 7 9 2 9 2 9 2 0 9 2 9 2 9 2 9 2 9 2 9 7 0 9 2 9 7 9 2 9 1 9 2 9 2 9 7 0 9 7 9 2
8 9 0 9 13 0 9 11 2
21 0 9 9 4 13 1 9 9 11 1 9 12 5 0 9 1 12 9 0 9 2
37 9 13 13 1 0 7 0 0 9 1 9 0 9 2 15 13 9 1 0 9 1 0 9 2 1 0 9 7 1 0 2 9 1 3 0 9 2
8 9 13 9 3 12 0 9 2
17 9 2 0 9 7 9 13 0 13 0 9 11 1 12 2 9 2
3 9 2 9
17 0 9 2 0 2 9 2 2 13 0 9 1 0 7 0 9 2
19 9 13 13 7 1 9 0 9 1 9 1 9 10 0 9 2 9 2 2
26 1 0 9 4 13 2 2 0 9 13 1 11 1 10 9 9 2 9 2 7 0 9 2 0 9 2
5 9 13 1 9 2
64 12 2 9 2 12 2 0 9 13 1 11 1 10 9 0 9 0 0 9 0 1 9 2 0 2 0 0 9 2 1 0 9 2 0 9 2 0 7 0 2 0 7 0 2 1 9 9 9 9 0 9 0 9 2 9 1 9 0 0 9 1 9 2 2
31 12 2 9 2 12 2 0 9 13 1 10 9 9 1 11 2 15 4 13 9 1 0 9 7 9 2 9 7 9 2 2
19 12 2 9 2 12 2 0 9 13 1 11 1 10 9 9 9 1 9 2
24 13 3 2 1 9 1 9 1 12 5 9 9 2 0 9 1 12 5 9 9 7 0 9 2
7 9 10 9 1 0 9 2
13 0 9 1 9 2 9 7 9 9 13 1 9 2
5 12 2 9 2 12
4 0 9 13 9
2 11 2
13 1 0 9 9 9 7 9 11 4 13 0 9 2
26 13 15 1 9 7 9 0 9 0 7 0 9 1 9 0 7 0 2 7 15 3 0 2 3 0 2
16 9 4 13 7 13 9 1 9 7 0 9 3 7 1 9 2
25 1 10 9 3 9 13 0 9 1 0 9 0 9 2 16 13 3 2 0 9 1 9 7 9 2
18 9 15 1 0 9 13 13 3 1 9 0 9 2 15 13 9 9 2
7 0 0 9 15 13 1 11
2 11 2
50 0 9 9 7 9 9 2 15 15 13 0 0 9 7 3 13 3 0 1 0 9 2 4 13 1 14 12 9 1 9 0 0 9 15 13 2 15 15 13 1 9 12 2 7 12 2 9 1 11 2
59 3 13 9 0 9 11 11 11 2 4 0 9 13 3 1 0 9 9 9 1 9 2 1 0 9 7 1 9 7 1 0 9 0 9 9 2 16 13 3 9 9 1 9 7 9 2 1 0 7 0 9 9 9 1 9 7 0 9 2
20 9 9 13 7 9 2 15 9 4 13 3 1 9 0 9 1 0 0 9 2
30 9 13 0 9 1 9 0 9 1 9 9 0 9 11 2 15 0 9 13 9 7 9 0 2 0 7 0 0 9 2
16 9 10 9 4 13 1 9 12 7 4 13 1 9 0 9 2
11 1 9 11 1 15 4 13 12 9 9 2
1 9
28 9 2 11 11 2 12 2 1 0 12 9 1 9 9 0 9 9 9 13 1 0 9 1 10 9 0 9 2
19 1 9 12 15 15 13 1 0 9 2 16 15 13 9 1 0 0 9 2
14 13 15 2 16 13 0 10 9 13 3 3 2 13 2
15 11 2 11 13 9 0 9 11 1 11 1 9 1 9 2
14 3 12 9 1 9 9 15 13 0 9 9 9 9 2
9 12 9 1 9 9 13 10 9 2
24 10 0 9 13 1 0 9 9 0 0 9 2 3 13 16 9 0 9 7 3 13 9 9 2
19 16 0 9 9 9 0 9 15 13 7 1 9 9 7 9 1 9 9 2
22 9 0 9 9 9 15 13 9 9 7 0 9 1 9 0 9 0 1 9 0 9 2
3 2 11 2
5 9 11 11 2 11
6 0 2 7 7 0 9
26 9 9 0 9 1 9 9 5 12 13 1 11 11 2 9 0 9 0 9 1 9 0 9 11 9 2
13 9 3 13 3 9 0 9 2 7 3 10 9 2
19 1 0 9 0 9 15 3 2 12 9 13 2 1 0 9 13 9 13 2
19 9 3 13 9 7 0 9 1 9 9 5 12 2 7 7 9 5 12 2
15 1 0 9 4 13 0 9 0 9 1 9 9 5 12 2
9 9 9 5 12 0 9 13 13 2
15 0 9 0 1 9 9 1 9 2 13 1 9 3 13 2
24 0 2 15 15 13 1 9 9 2 15 3 3 2 13 0 9 1 9 9 13 1 12 9 2
20 9 0 9 13 1 9 9 5 12 2 15 9 13 13 0 9 1 0 9 2
14 1 11 13 9 9 9 1 9 1 9 9 0 9 2
14 9 1 9 13 9 2 15 13 0 9 1 0 9 2
10 15 15 3 13 1 9 9 0 9 2
33 15 9 9 1 9 4 13 1 11 11 13 2 16 0 9 9 13 9 1 9 1 9 10 9 2 3 1 9 9 5 12 3 2
19 16 13 1 9 2 13 3 13 0 9 2 16 4 13 9 0 9 9 2
18 9 1 9 13 1 11 2 11 13 16 1 9 2 9 0 2 9 2
20 13 3 2 13 2 16 9 4 13 9 2 15 13 9 9 1 9 0 9 2
14 9 4 13 4 13 1 10 9 3 7 1 0 9 2
9 9 0 9 13 1 9 9 9 2
11 13 13 7 0 1 0 9 1 0 9 2
21 9 15 7 3 13 1 9 0 9 1 9 2 9 7 9 0 9 2 11 2 2
11 9 1 11 13 3 9 2 11 1 0 2
16 9 7 3 13 0 9 0 1 9 9 2 15 4 3 13 2
15 1 0 9 13 9 1 0 9 9 1 9 9 5 12 2
7 0 9 13 13 3 3 2
11 0 9 13 1 0 9 9 1 0 9 2
19 9 1 0 9 7 9 3 2 13 2 16 4 13 13 0 9 1 9 2
22 13 15 2 16 9 2 15 4 3 13 2 13 1 9 0 7 13 1 9 15 9 2
3 2 11 2
7 9 13 2 7 9 9 13
8 0 0 9 9 9 13 0 9
2 11 11
7 0 9 13 0 9 3 2
31 1 9 9 9 12 1 12 5 1 12 9 13 3 1 0 9 9 9 2 1 3 9 9 9 2 1 12 9 2 9 2
6 15 13 13 3 0 2
22 9 13 9 1 9 0 9 2 16 0 9 2 15 4 1 9 13 2 3 13 3 2
19 0 9 9 13 12 9 2 9 7 13 1 12 9 0 16 9 0 9 2
12 9 9 7 1 0 9 13 3 1 12 9 2
27 1 9 0 9 4 13 9 9 1 12 9 2 0 2 1 12 5 2 13 11 9 2 9 12 9 2 2
16 9 13 12 9 2 0 2 9 9 3 0 9 2 11 11 2
10 10 9 13 1 12 5 1 12 9 2
15 9 12 9 1 10 9 13 1 9 1 0 9 1 9 2
21 0 9 15 13 1 12 9 0 9 7 9 13 3 9 11 1 9 3 12 9 2
23 13 15 7 9 0 9 2 0 11 7 11 0 2 7 16 1 3 0 9 10 9 9 2
23 0 9 0 9 2 9 11 2 15 13 16 0 3 7 1 9 12 0 1 0 0 9 2
25 10 9 13 3 1 12 5 1 12 9 2 7 0 9 12 9 2 9 15 13 1 0 0 9 2
20 16 7 13 2 10 9 13 3 1 9 1 0 9 1 9 2 13 0 9 2
8 9 9 9 13 3 0 9 2
21 7 13 0 2 16 9 13 1 0 9 9 9 7 16 9 1 0 9 4 13 2
16 1 9 1 9 1 0 9 9 3 3 7 0 9 3 13 2
4 9 1 0 9
13 11 11 2 12 2 12 2 13 1 0 0 9 2
8 11 9 13 3 1 3 0 2
11 1 0 3 13 9 2 9 11 2 11 2
16 3 0 13 9 9 1 0 9 2 10 9 9 12 13 9 2
18 1 9 1 11 11 13 9 2 15 13 11 2 11 2 9 9 11 2
20 1 0 9 9 1 0 0 9 13 1 0 9 11 2 11 7 11 2 11 2
9 2 11 2 2 11 12 2 12 2
5 9 7 0 1 11
6 0 0 9 1 9 12
4 9 15 9 13
4 1 9 0 9
2 11 11
15 9 9 1 9 1 9 7 0 9 1 9 13 0 9 2
27 16 4 15 15 15 0 13 2 13 9 13 9 9 1 10 9 2 7 9 9 13 10 9 1 10 9 2
19 9 2 1 15 9 13 1 9 0 10 9 2 13 9 12 7 0 9 2
41 1 9 0 9 13 9 9 1 10 0 9 1 9 7 10 0 9 9 2 3 2 9 1 9 0 0 9 9 7 1 9 1 9 2 15 15 13 1 9 2 2
24 1 9 12 9 9 15 0 9 9 13 3 1 9 2 16 13 9 1 9 9 1 0 9 2
18 1 15 2 16 4 9 9 1 9 3 13 2 13 4 13 10 9 2
31 12 2 9 13 13 9 2 7 2 13 13 1 0 9 9 10 9 2 1 10 9 15 13 7 9 1 9 0 9 2 2
21 12 2 9 7 0 0 7 0 9 2 15 13 10 9 2 13 13 10 0 9 2
19 3 9 13 1 10 9 7 3 2 16 1 15 13 1 10 7 0 9 2
20 1 15 9 13 7 1 9 2 15 9 13 0 9 1 9 9 7 0 9 2
18 12 2 9 13 9 13 1 9 10 0 9 7 1 0 9 1 15 2
34 15 13 7 15 13 1 0 9 1 9 0 9 2 13 9 12 9 12 2 12 9 2 2 15 13 1 10 9 0 9 1 9 9 2
18 1 9 10 9 13 9 1 9 2 15 13 9 1 0 9 0 9 2
27 13 15 15 7 1 0 9 2 9 0 9 1 9 1 9 2 15 13 0 13 1 9 7 1 9 9 2
36 3 9 13 1 9 2 15 9 13 1 9 1 9 7 1 15 2 7 1 9 1 0 9 2 9 13 9 2 3 9 13 1 9 9 2 2
16 13 0 13 2 16 9 9 13 1 10 9 1 9 3 0 2
16 9 3 13 1 9 1 0 9 2 15 13 9 1 0 9 2
17 13 3 0 2 16 13 10 9 7 3 2 0 2 0 9 9 2
59 15 13 1 9 12 9 9 9 15 10 9 3 7 3 13 1 9 2 16 9 3 13 1 9 9 9 1 9 9 2 10 9 2 9 0 0 9 7 16 10 9 13 0 9 9 2 15 13 13 2 16 15 3 13 13 9 1 9 2
6 1 11 3 9 1 9
2 11 2
15 9 9 1 11 13 1 9 1 12 9 1 0 12 9 2
9 13 15 1 9 0 0 0 9 2
16 1 0 9 13 9 9 1 9 1 12 12 1 0 12 12 2
13 3 1 9 4 1 11 13 1 9 12 12 9 2
3 9 2 9
33 13 1 9 9 2 9 2 9 7 0 9 2 0 9 2 0 0 9 2 15 13 0 9 1 0 9 0 1 9 7 9 9 2
20 13 10 9 2 0 9 9 2 0 9 2 0 9 9 2 0 9 1 9 2
11 9 7 9 9 2 12 2 9 1 11 2
14 9 7 9 9 2 12 2 7 12 2 9 1 11 2
23 9 9 13 0 9 2 0 9 2 9 9 2 0 2 0 7 0 9 2 9 9 3 2
11 9 7 9 9 2 12 2 9 1 11 2
20 9 2 0 9 0 0 7 0 9 2 1 10 9 13 9 9 1 0 9 2
11 9 7 9 9 2 12 2 9 1 11 2
9 13 2 11 9 2 9 2 0 2
37 9 1 9 2 0 9 2 15 13 9 1 0 7 0 9 0 9 2 3 2 1 9 0 0 9 2 9 9 2 9 9 2 9 0 9 3 2
7 0 1 9 7 0 9 2
11 9 7 9 9 2 12 2 9 1 11 2
11 13 2 11 2 2 9 2 9 2 0 2
5 9 1 11 1 9
2 11 2
42 11 13 1 12 2 9 0 9 0 9 9 0 9 1 0 9 12 9 2 14 12 9 2 2 16 4 3 13 1 0 9 9 9 2 15 15 13 1 12 2 9 2
7 9 4 13 1 9 9 2
22 13 15 2 16 1 12 2 9 13 9 1 12 9 7 9 3 13 12 9 10 9 2
16 1 0 0 9 13 1 9 0 0 0 9 1 11 12 9 2
29 9 9 13 9 0 9 1 0 9 2 15 13 2 16 4 0 0 9 13 14 12 9 9 9 1 12 2 9 2
14 9 15 1 9 0 9 13 3 9 7 9 1 9 2
2 1 9
2 11 2
25 12 1 9 0 9 3 0 9 13 9 9 9 1 11 11 11 1 10 9 13 15 9 0 9 2
19 1 15 13 13 2 16 9 9 1 9 1 9 9 3 13 14 1 9 2
31 1 0 9 10 0 9 1 9 9 13 9 0 9 0 9 7 9 1 9 9 2 0 9 1 9 7 9 0 0 9 2
19 3 1 15 13 9 9 7 0 1 9 0 9 1 9 3 0 0 9 2
24 0 9 3 13 2 16 3 0 9 2 10 0 9 13 9 9 9 2 13 1 0 9 9 2
25 1 9 13 0 15 3 13 1 9 0 0 7 0 9 1 9 10 9 7 9 1 9 9 9 2
21 7 13 1 0 9 2 9 2 9 7 0 9 2 13 11 2 11 2 2 6 2
6 0 9 15 13 1 9
17 9 0 9 1 0 9 7 0 9 1 15 13 0 9 1 0 9
2 11 11
11 9 13 2 13 7 13 3 1 15 3 2
14 3 12 9 0 9 13 0 10 9 13 3 1 9 2
18 9 9 13 3 1 9 0 9 2 7 3 1 9 9 9 1 9 2
15 3 13 3 1 9 2 15 1 9 0 9 3 3 13 2
7 0 7 0 9 13 9 2
23 13 4 9 9 1 11 13 2 16 9 0 9 13 10 9 2 7 13 15 3 14 3 2
20 7 15 7 3 2 16 0 9 1 10 9 13 13 9 2 16 9 13 9 2
21 1 9 10 9 13 0 0 9 2 15 15 13 1 9 9 1 9 1 0 9 2
14 7 3 15 9 13 1 9 7 3 1 15 9 13 2
16 0 9 13 0 7 0 9 1 9 2 16 10 9 13 9 2
28 9 9 15 13 0 9 0 9 2 7 15 3 2 16 3 3 13 7 0 2 7 0 9 1 9 0 9 2
4 9 13 0 2
29 10 9 2 3 11 13 10 9 11 11 2 13 0 9 1 9 9 2 16 1 0 9 13 0 9 13 1 9 2
34 9 15 13 2 16 16 15 13 9 2 0 9 15 3 13 2 1 9 2 15 15 1 9 13 7 3 2 3 1 12 9 1 9 2
18 1 9 12 13 3 0 9 0 9 1 11 12 9 2 3 3 0 2
12 1 0 9 15 13 3 12 2 0 3 3 2
9 14 12 0 9 3 13 1 9 2
7 9 15 13 1 9 3 2
22 1 0 0 9 3 13 0 9 2 15 13 9 2 16 9 13 0 1 9 0 9 2
9 9 15 13 3 16 1 0 9 2
12 0 9 1 9 2 16 13 15 3 0 9 2
20 0 9 1 9 1 9 12 9 13 9 0 9 11 7 13 1 12 12 9 2
15 0 9 0 9 13 1 0 9 9 7 13 14 12 12 2
24 9 1 9 13 1 11 2 3 0 9 13 2 12 7 15 0 12 2 16 10 9 13 0 2
34 13 7 14 1 15 2 13 3 3 9 2 7 7 0 9 2 15 13 9 1 9 7 0 9 2 15 15 13 9 12 9 2 9 2
25 0 9 13 1 11 11 2 9 9 9 7 9 0 9 2 9 10 9 14 1 0 9 0 9 2
11 15 13 9 9 0 13 1 0 9 9 2
20 9 0 9 4 3 13 9 0 9 1 9 2 15 15 13 7 1 9 9 2
18 13 15 3 9 13 1 0 0 9 2 15 13 0 1 9 0 9 2
13 1 0 9 15 13 9 0 9 2 3 7 0 2
8 9 15 1 15 0 9 13 2
15 13 3 1 9 2 16 3 13 14 9 1 9 0 9 2
13 0 9 3 13 10 9 16 9 7 0 0 9 2
11 1 9 9 4 1 10 9 13 13 9 2
7 16 13 2 3 3 15 2
19 9 0 9 13 13 0 9 9 3 2 16 4 15 9 13 9 13 3 2
14 1 9 1 0 9 15 4 13 13 1 0 9 9 2
2 0 9
41 9 2 15 11 11 13 1 9 0 9 2 15 3 13 2 1 0 7 0 9 9 3 1 9 1 11 4 0 9 13 2 7 3 3 13 2 12 9 0 9 2
33 9 11 11 1 9 12 13 1 10 9 9 2 15 10 0 0 9 7 0 9 3 13 1 15 0 2 15 3 1 10 9 13 2
8 2 11 2 2 11 2 12 2
3 9 9 0
2 11 2
20 0 9 1 9 9 2 15 13 9 9 7 9 9 2 13 3 12 9 9 2
18 1 0 9 13 0 1 12 5 2 7 2 14 1 12 9 2 9 2
24 1 9 15 3 13 0 9 2 1 15 13 1 0 9 9 9 1 0 9 9 0 0 9 2
3 9 9 13
2 11 2
33 0 9 9 1 9 12 2 12 2 9 2 9 2 13 1 12 9 2 1 12 9 2 9 7 13 3 0 1 9 12 2 12 2
16 0 9 7 13 1 0 12 9 1 0 9 1 12 9 9 2
12 13 15 1 10 0 9 0 9 11 2 11 2
18 0 9 15 1 0 9 12 13 1 12 9 2 1 12 9 2 9 2
17 0 9 9 1 11 13 2 16 0 9 0 9 9 13 3 0 2
23 12 0 9 3 13 9 0 9 7 9 9 15 13 3 2 16 13 0 13 0 9 9 2
32 1 0 9 9 12 2 12 15 4 13 9 0 1 9 9 12 9 2 9 1 9 1 12 9 2 9 1 9 12 2 12 2
18 1 0 9 15 13 12 9 2 9 0 9 1 0 12 9 2 9 2
25 0 9 4 13 1 0 9 1 11 13 0 0 9 2 7 1 9 11 2 3 15 13 9 9 2
13 1 9 9 15 13 13 3 0 9 1 0 11 2
14 9 1 0 9 7 1 11 4 3 13 0 9 9 2
7 0 9 9 11 1 0 11
5 0 11 2 11 2
27 0 9 11 11 2 0 2 13 12 9 0 9 11 11 2 0 2 9 2 2 1 15 13 12 9 9 2
13 0 12 9 9 9 4 13 1 0 9 0 9 2
7 13 15 9 9 11 11 2
23 0 9 1 9 12 9 9 9 9 0 9 9 13 9 11 1 0 9 11 12 0 9 2
13 11 10 9 13 1 9 1 9 9 1 0 9 2
32 9 11 15 3 13 13 1 0 9 1 0 9 3 12 9 9 2 12 9 9 2 1 9 0 9 1 9 9 7 9 9 2
12 15 15 9 9 1 9 11 13 1 12 9 2
47 16 13 0 2 16 4 10 9 13 0 9 1 10 9 1 0 9 2 13 2 16 15 11 2 0 2 9 2 2 13 1 9 0 9 10 0 9 2 13 9 7 0 9 11 11 11 2
36 0 9 11 3 1 9 0 10 0 9 1 11 2 11 11 0 2 0 2 0 2 0 2 2 4 13 11 13 9 1 0 9 1 0 11 2
20 11 13 2 16 10 9 13 1 11 9 3 3 16 12 9 7 3 9 13 2
13 11 11 2 0 2 13 1 0 2 11 1 11 2
20 0 9 9 10 0 9 13 9 2 9 7 9 0 7 0 9 7 0 9 2
17 13 12 9 1 11 7 12 1 11 7 0 9 1 11 7 11 2
1 3
20 0 0 9 0 9 11 11 4 1 9 1 12 2 9 13 3 1 12 9 2
9 0 9 13 4 1 9 0 9 13
21 9 0 0 13 9 1 9 11 1 9 9 0 9 1 0 9 0 9 11 11 2
4 0 2 9 11
7 0 9 11 13 12 9 2
18 1 9 11 12 2 11 12 5 7 9 9 11 13 0 9 12 9 2
18 1 9 9 11 12 15 13 0 0 9 2 9 2 12 9 2 9 2
18 1 9 11 12 5 7 9 9 11 13 9 12 2 3 2 12 9 2
33 1 11 13 9 12 2 9 2 0 9 9 1 10 9 2 1 11 12 2 11 12 5 7 9 9 11 12 2 12 7 12 9 2
5 0 11 3 1 11
3 0 11 2
19 0 9 7 9 3 1 0 9 13 9 0 9 0 11 7 9 1 11 2
13 13 15 0 9 0 9 1 0 9 11 2 11 2
8 1 9 11 4 15 9 13 2
33 3 13 1 9 9 0 9 2 15 13 13 1 9 1 0 0 9 7 13 9 9 9 0 0 9 2 13 13 9 7 9 13 2
17 1 11 4 13 13 15 9 7 0 9 9 9 1 11 1 9 2
19 9 1 9 13 9 12 9 9 2 7 1 0 9 3 14 12 9 9 2
3 9 1 9
7 11 2 11 2 11 2 2
29 9 9 11 2 11 3 1 9 9 11 13 2 16 10 9 1 9 0 9 15 3 13 1 9 9 11 2 11 2
15 15 15 13 2 16 9 4 13 4 1 10 0 9 13 2
42 9 9 0 2 0 2 11 2 11 2 11 2 15 9 13 2 3 13 2 16 9 11 1 12 9 10 9 13 9 9 7 1 0 3 13 2 16 9 13 14 0 9
33 1 11 11 10 9 9 1 0 9 9 13 10 0 9 7 16 4 4 13 9 2 13 4 1 15 0 2 0 2 11 2 9 2
23 11 13 2 16 13 0 13 1 12 9 9 9 2 16 4 3 13 1 0 0 9 9 2
16 1 9 13 9 0 0 9 9 10 9 2 3 9 2 13 2
8 3 1 9 12 9 1 9 12
5 9 4 13 13 11
2 11 2
17 11 4 13 13 0 2 16 13 13 3 9 0 9 7 13 9 2
23 9 9 13 1 11 2 13 1 9 9 9 0 9 11 11 11 1 9 9 11 1 9 2
31 13 3 1 9 0 9 9 11 11 2 15 13 2 16 10 9 13 13 13 1 11 2 16 15 12 9 4 13 0 9 2
15 11 13 2 16 11 13 13 9 1 9 0 9 1 11 2
10 1 11 13 7 9 13 11 1 9 2
15 0 9 11 2 11 13 2 0 9 9 11 13 0 11 2
19 1 11 4 15 13 9 13 1 9 9 2 15 4 13 9 1 0 9 2
4 3 1 9 12
2 0 9
38 0 0 9 0 9 2 12 2 15 13 0 7 0 9 12 1 0 9 10 9 2 9 0 7 0 9 2 9 7 9 11 11 2 12 2 12 2 2
45 1 9 0 9 13 0 9 2 0 9 12 2 7 12 2 9 11 11 2 10 0 0 9 11 1 11 2 7 3 7 9 2 1 0 9 0 9 12 2 9 11 2 11 11 2
8 2 11 2 2 11 2 12 2
5 1 11 13 0 9
9 11 2 11 2 11 2 11 2 2
30 0 0 9 2 15 0 9 1 11 1 12 9 13 7 1 9 9 13 9 11 11 2 15 1 0 9 9 3 13 2
15 11 15 3 13 9 9 9 9 1 11 9 2 11 11 2
35 16 9 0 9 4 0 9 13 1 9 12 7 9 9 9 13 12 9 2 9 0 9 13 3 12 7 0 2 3 13 1 9 13 9 2
44 0 9 13 3 3 13 0 9 2 7 16 1 15 15 13 0 9 2 9 7 9 0 9 2 7 4 15 12 7 12 9 13 3 9 2 13 15 0 9 7 3 7 9 2
12 1 0 9 11 13 3 13 9 9 0 9 2
23 9 10 12 9 0 0 9 2 15 13 12 9 0 9 2 9 13 12 2 9 0 9 2
15 1 9 11 7 9 1 9 11 11 13 3 9 0 9 2
20 9 9 0 9 9 11 9 2 11 13 2 16 9 4 13 1 11 16 9 2
9 1 0 9 13 0 7 0 9 2
5 9 9 11 13 2
18 0 9 13 2 16 9 4 9 13 16 0 9 2 3 13 7 13 2
39 9 9 1 9 11 3 13 1 9 2 7 1 9 9 11 3 13 12 9 9 2 10 0 9 9 0 1 9 9 9 13 1 11 11 2 0 0 9 2
19 9 10 9 1 9 7 1 9 13 3 0 2 16 4 13 0 0 9 2
17 15 13 2 16 1 11 13 13 0 9 9 2 13 9 2 11 2
12 9 11 3 3 13 9 0 1 0 9 13 2
19 1 11 2 11 9 9 13 0 2 7 0 9 9 1 10 9 13 0 2
28 0 9 4 1 11 13 3 15 2 7 1 9 2 11 7 3 15 13 13 2 3 15 0 9 1 9 13 2
5 9 1 9 9 13
13 1 0 9 13 9 11 11 1 0 9 9 11 11
19 9 3 13 0 9 9 9 2 7 1 10 0 9 3 13 3 3 13 2
22 0 12 9 0 1 0 9 11 15 3 13 2 16 0 9 13 0 9 16 0 9 2
5 15 15 15 13 2
7 13 3 0 1 10 9 2
20 9 13 13 1 9 1 15 2 15 13 9 9 9 7 9 9 0 9 9 2
6 13 4 15 0 9 2
13 13 2 10 0 9 0 9 9 13 9 1 9 2
11 13 15 13 0 9 16 9 10 0 9 2
16 13 3 0 1 15 2 15 13 0 15 13 1 0 9 9 2
14 13 13 0 9 13 15 10 9 2 13 15 7 13 2
10 15 3 2 13 2 13 9 1 9 2
21 16 15 13 0 9 9 11 1 0 9 2 3 15 13 13 2 16 13 0 9 2
11 1 10 9 15 3 0 9 13 1 9 2
6 13 3 2 15 13 2
18 0 9 4 15 3 13 2 16 4 13 1 9 11 1 0 9 9 2
5 15 9 13 13 2
5 7 15 0 9 2
17 3 13 1 9 2 16 4 0 0 9 13 9 16 9 0 9 2
4 3 15 13 2
20 0 13 2 16 9 0 9 13 3 10 9 2 1 15 1 9 9 7 9 2
3 15 0 2
22 13 0 9 2 0 0 9 2 0 9 2 9 2 9 1 9 2 10 9 1 9 2
14 15 15 10 9 9 13 2 15 13 3 2 3 13 2
47 16 13 3 1 15 2 16 4 13 13 9 1 9 2 3 3 3 13 2 3 13 0 9 1 0 11 2 15 4 15 15 3 13 2 16 4 15 13 3 0 9 7 1 10 13 9 2
16 15 13 9 0 9 2 15 9 13 10 0 9 1 0 9 2
17 13 1 15 3 0 13 10 9 3 1 9 2 16 15 4 13 2
28 10 9 1 15 13 1 12 12 9 0 9 0 9 7 0 9 13 3 3 0 9 1 9 1 0 0 9 2
31 3 4 15 13 1 0 9 2 16 0 9 2 15 13 13 0 0 9 2 13 0 0 9 2 15 4 13 13 7 13 2
18 9 2 16 4 15 15 13 13 0 9 0 9 2 13 1 9 0 2
14 13 1 0 9 0 3 7 13 15 9 9 0 3 2
6 13 3 9 13 9 2
14 9 13 13 0 9 3 1 10 9 12 2 9 12 2
34 0 9 14 13 15 2 16 9 9 1 11 13 3 0 16 1 12 9 2 1 10 9 13 13 9 9 2 13 2 1 11 7 11 2
22 1 15 13 1 0 9 9 7 10 9 1 0 9 1 9 9 13 12 2 12 9 2
11 9 9 9 4 13 13 0 9 0 9 2
17 16 4 10 9 13 3 0 16 9 2 3 4 13 9 1 9 2
13 13 4 3 9 2 13 9 7 13 9 0 9 2
8 1 15 7 13 9 3 0 2
33 0 9 13 9 1 0 9 9 16 9 7 1 0 9 1 0 0 9 0 9 13 2 16 0 9 13 9 12 2 12 9 9 2
13 10 9 4 13 0 9 2 3 0 9 7 9 2
15 13 3 9 2 16 4 13 1 9 13 9 7 13 9 2
11 10 7 0 9 13 0 13 3 1 9 2
6 13 15 9 0 11 2
8 0 11 15 3 13 9 3 2
11 4 1 15 3 13 7 1 0 0 9 2
22 0 9 4 13 2 16 4 15 12 0 9 13 13 12 1 0 2 7 13 9 0 2
10 1 10 9 1 10 0 9 15 13 2
12 16 15 3 13 3 2 13 1 15 0 9 2
11 0 9 13 1 0 9 2 15 13 0 9
4 9 11 2 11
6 11 10 9 11 14 13
2 11 2
36 9 9 11 11 13 1 1 0 9 13 9 2 16 0 9 11 11 2 11 2 15 15 13 1 0 9 1 11 2 13 9 12 0 9 11 2
7 11 15 3 13 1 9 2
15 9 10 9 14 13 9 11 1 11 2 15 13 0 11 2
14 1 9 9 11 13 1 0 0 0 9 3 1 9 2
6 9 9 4 13 13 9
5 11 2 11 2 2
24 9 0 9 13 9 9 2 15 15 13 9 1 9 0 0 9 7 9 9 0 7 0 9 2
18 16 1 0 7 0 9 13 0 9 3 3 2 9 15 15 13 13 2
9 3 7 3 14 3 7 14 15 2
10 9 4 13 10 9 9 1 0 9 2
22 1 15 13 9 0 13 14 1 12 9 3 0 2 15 13 0 9 13 2 14 3 2
16 1 0 9 15 9 0 13 1 12 7 0 9 1 12 9 2
19 9 9 1 11 12 0 13 9 9 1 10 9 2 15 13 0 0 9 2
7 0 12 9 15 7 13 2
14 7 1 0 9 0 1 0 9 13 9 9 10 9 2
33 9 11 11 11 13 2 16 9 9 13 1 0 9 0 9 3 3 2 16 15 9 4 13 0 9 13 1 15 1 9 0 9 2
13 1 10 9 15 1 15 4 3 13 3 16 3 2
12 3 13 1 9 9 0 1 9 1 12 9 2
25 0 0 9 2 16 3 9 2 13 3 14 9 0 9 0 9 2 7 15 14 1 9 12 9 2
28 3 9 9 0 15 7 13 1 9 2 16 13 1 0 9 14 1 9 7 4 3 13 0 9 1 0 9 2
20 9 1 9 9 1 0 9 1 9 12 9 13 1 9 3 0 1 9 0 9
5 9 11 11 2 11
4 0 9 1 9
5 11 2 11 2 2
36 1 12 9 0 0 9 2 9 11 2 0 1 9 12 2 15 13 1 11 1 0 9 2 4 13 9 0 9 13 2 1 10 9 15 13 2
22 9 13 1 15 9 1 9 12 9 7 1 9 13 0 9 2 15 13 1 10 9 2
10 9 1 0 9 9 3 13 9 9 2
6 0 9 13 1 9 2
26 13 4 3 13 3 2 16 4 15 13 0 13 1 9 2 7 3 13 13 0 9 2 13 11 11 2
19 3 15 14 1 11 13 13 0 9 2 15 13 13 7 12 9 1 9 2
8 9 9 13 3 0 9 9 2
25 13 2 14 15 9 1 10 9 2 4 13 7 1 0 9 7 13 15 3 1 10 9 1 9 2
12 9 4 13 13 3 9 2 9 9 3 2 2
15 3 4 13 0 9 0 9 1 9 13 1 10 0 9 2
21 3 3 4 13 3 1 11 1 0 0 9 7 1 11 7 1 11 1 0 9 2
15 9 1 9 12 9 13 1 9 3 0 1 9 0 9 2
7 0 0 9 13 12 9 2
5 9 13 1 9 11
2 11 2
20 1 9 0 9 11 7 1 10 9 1 9 4 1 0 9 13 12 9 9 2
14 13 15 1 9 0 9 2 15 1 9 13 9 11 2
12 1 9 4 15 1 0 9 13 12 9 9 2
11 9 9 7 9 11 13 3 12 2 12 2
20 3 16 12 9 9 0 9 2 12 9 2 13 1 9 0 9 9 0 9 2
11 9 13 12 12 2 3 2 12 9 0 2
4 12 9 13 2
14 9 13 2 16 1 9 0 9 3 13 12 9 9 2
7 0 9 13 12 9 9 2
3 0 9 9
20 1 0 9 9 11 11 13 1 9 9 3 3 0 2 7 3 0 0 9 2
27 1 0 9 9 15 13 1 9 2 3 9 13 3 9 2 3 13 1 9 0 11 2 13 10 0 9 2
28 1 0 7 0 9 12 0 9 1 9 12 2 7 12 2 9 13 9 0 9 2 0 15 1 9 1 9 2
9 2 11 2 2 11 12 2 12 2
5 0 9 9 1 9
5 11 2 11 2 2
22 9 9 2 0 9 7 9 0 9 13 0 1 9 12 2 9 1 9 12 2 9 2
11 9 13 0 2 9 7 9 0 9 9 2
17 9 15 13 3 1 9 7 13 15 1 15 0 9 0 1 9 2
43 1 12 2 9 13 3 15 9 2 1 9 1 9 7 0 9 2 3 1 9 13 0 9 2 3 0 7 0 9 2 11 2 13 1 0 0 9 1 0 1 0 9 2
6 3 7 11 15 13 9
2 11 2
33 1 12 9 9 2 9 7 9 9 1 12 9 12 9 15 3 1 9 0 9 13 1 10 0 9 1 0 9 0 9 1 11 2
10 15 4 13 9 1 0 9 10 9 2
20 1 0 9 13 0 9 9 3 3 1 0 9 0 9 1 0 9 9 0 2
15 3 16 1 0 9 13 1 9 1 11 0 9 7 3 2
22 3 3 13 0 9 1 11 2 12 9 2 11 12 2 11 12 7 1 11 12 9 2
12 3 11 13 1 12 9 1 0 11 7 11 2
1 3
30 12 0 9 0 9 2 0 9 2 9 7 9 1 9 13 1 9 13 1 0 9 1 11 9 9 16 9 0 9 2
31 9 11 11 13 1 0 11 9 12 2 9 12 1 12 2 9 2 1 0 9 9 9 11 11 2 0 9 1 10 9 2
20 9 9 0 2 9 2 9 2 9 7 9 11 12 13 3 1 11 1 11 2
6 11 13 12 5 0 9
3 0 9 2
11 0 9 13 13 13 9 0 9 1 11 2
14 1 1 0 0 9 13 0 9 9 3 1 9 11 2
20 13 15 1 9 1 9 9 7 9 11 11 2 11 10 0 9 11 2 11 2
20 1 9 0 9 13 2 16 3 3 13 1 12 9 0 9 9 1 0 9 2
16 9 0 9 9 1 11 1 11 1 11 13 1 11 3 3 2
11 1 11 15 0 9 13 3 12 2 9 2
23 11 13 2 16 0 9 9 1 11 1 11 4 3 13 1 9 9 12 1 9 0 9 2
12 0 9 9 4 3 13 4 13 1 9 12 2
5 1 9 11 1 11
5 11 2 11 2 2
18 9 9 11 11 3 11 13 2 16 1 9 1 9 3 9 9 13 2
17 15 3 4 15 1 15 13 2 15 3 4 1 10 13 10 9 2
29 11 4 13 2 15 9 13 2 14 1 15 2 13 15 15 10 9 2 9 2 9 2 2 2 13 11 2 11 2
17 0 9 4 13 13 3 9 0 9 9 11 1 9 9 11 11 2
20 11 3 3 13 2 16 4 1 9 1 9 0 9 9 13 9 10 0 9 2
6 11 2 11 1 9 9
3 1 0 9
6 0 11 2 11 2 2
20 9 9 7 0 0 9 13 0 9 11 2 11 1 9 1 0 9 1 9 2
13 13 15 3 1 0 11 9 11 2 11 11 11 2
26 13 13 10 9 9 2 15 13 13 1 0 9 2 9 9 1 0 3 0 9 2 13 11 2 11 2
18 1 0 13 9 9 0 9 1 9 2 16 15 4 13 10 0 9 2
35 1 11 2 11 4 15 4 13 3 9 2 15 13 3 1 12 9 9 10 9 2 15 13 9 2 15 4 13 9 3 13 2 3 13 2
11 1 0 9 4 13 9 1 9 1 11 13
5 11 2 11 2 2
26 0 9 0 9 2 11 2 13 0 9 0 9 0 2 9 0 9 2 9 0 9 7 3 0 9 2
15 0 9 0 9 13 1 0 0 9 11 11 1 0 9 2
8 3 1 15 13 9 0 9 2
25 1 9 0 9 0 9 13 10 9 1 15 2 16 4 15 0 9 13 9 1 9 1 0 9 2
33 1 9 11 2 16 13 9 11 9 2 16 0 9 1 11 13 1 0 9 9 1 9 2 13 11 2 11 2 16 3 3 14 2
36 1 0 9 13 11 3 13 0 9 9 1 9 2 13 0 9 7 9 0 9 2 13 9 3 0 9 2 7 13 9 1 9 7 0 9 2
44 1 9 2 3 4 13 0 9 13 9 1 3 0 9 2 13 10 9 11 11 2 11 2 2 16 9 0 11 4 13 9 2 7 3 3 13 9 1 9 9 1 9 11 2
3 0 9 13
7 11 2 11 2 11 2 2
22 7 1 0 9 9 0 7 0 9 15 9 9 2 9 7 9 13 1 9 0 9 2
12 1 9 15 13 9 9 2 9 9 11 11 2
25 9 15 1 15 13 2 16 0 9 13 9 2 7 13 0 15 13 14 1 9 0 9 0 9 2
14 9 9 7 9 13 2 16 9 4 13 4 13 3 2
18 9 1 9 9 1 0 0 9 4 1 11 13 13 1 9 1 9 2
10 9 15 3 13 9 9 1 0 9 2
16 1 11 9 3 13 13 7 9 4 1 15 13 13 3 3 2
14 3 9 3 13 9 0 9 9 1 9 1 0 9 2
26 1 10 9 2 3 13 9 2 16 15 1 9 0 9 13 0 9 2 13 3 1 9 9 1 9 2
45 1 11 15 15 9 13 1 15 2 16 9 13 9 2 7 13 0 13 0 9 9 7 13 9 9 9 1 9 3 2 16 4 4 9 3 13 1 9 9 2 9 7 0 9 2
3 1 0 9
26 1 0 9 2 3 0 1 0 9 0 0 9 2 15 1 10 9 13 1 0 9 2 0 11 11 2
29 1 0 9 1 9 7 9 9 0 9 1 0 9 13 9 9 0 11 1 11 2 9 2 15 13 0 9 9 2
16 9 0 0 9 15 13 1 9 2 15 15 7 13 0 9 2
8 2 11 2 2 11 2 12 2
6 9 9 0 7 0 9
6 9 11 2 11 2 11
11 13 2 14 9 9 0 2 13 0 13 9
7 11 2 11 2 11 2 2
19 9 9 15 13 9 0 9 2 15 1 10 9 13 13 9 1 0 9 2
26 16 15 13 2 16 9 9 13 3 1 9 1 9 2 4 10 9 13 13 0 9 7 9 1 9 2
28 9 9 11 11 2 11 2 11 2 13 1 11 2 16 1 9 13 9 2 16 15 1 0 9 13 9 9 2
16 13 4 2 16 11 13 10 9 2 15 4 1 15 13 13 2
25 13 2 16 1 9 4 3 13 0 9 2 15 4 13 9 0 9 1 9 1 0 9 0 9 2
27 16 4 13 9 2 16 1 10 9 13 1 0 9 10 9 2 1 15 4 15 1 9 13 2 13 11 2
13 1 0 13 9 0 9 9 11 11 2 11 2 2
11 1 0 9 1 0 9 10 9 13 9 2
17 0 9 3 13 13 9 1 9 14 3 2 16 13 1 15 0 2
23 11 13 13 2 16 13 0 13 0 9 7 9 1 9 2 15 13 0 7 13 0 9 2
26 0 9 0 9 4 13 13 9 12 9 2 3 0 0 9 2 16 4 3 15 0 13 0 2 13 2
19 9 11 11 2 11 2 9 2 16 1 9 13 9 3 7 9 2 13 2
15 13 4 1 9 2 16 9 0 1 9 13 0 2 13 2
19 9 11 13 1 15 3 0 1 0 9 2 7 15 1 9 13 0 9 2
10 0 9 3 13 3 1 9 2 13 2
6 0 9 0 9 3 13
2 11 2
11 0 9 13 9 0 9 11 1 3 0 2
19 13 15 1 9 9 9 1 9 0 9 0 9 9 1 0 9 12 9 2
21 9 0 9 13 12 5 9 1 3 0 7 1 12 5 9 1 10 9 7 13 2
17 3 1 3 0 13 9 0 9 12 5 0 7 1 0 12 5 2
20 1 11 7 1 11 13 9 9 2 15 9 9 13 16 0 2 14 3 0 2
15 9 9 0 9 13 1 9 1 9 12 1 9 9 3 2
20 0 9 9 16 1 9 15 3 13 2 16 1 9 9 0 9 13 0 13 2
22 9 2 16 13 0 13 0 0 9 1 0 9 0 9 7 9 2 13 12 5 0 2
11 3 12 5 9 13 2 16 15 13 0 2
9 9 1 11 11 2 9 11 2 11
14 1 9 9 13 9 1 9 0 9 3 1 0 9 2
10 13 10 9 1 0 9 10 0 9 2
26 15 0 3 4 13 7 13 1 15 2 16 13 0 9 2 3 9 9 2 15 13 0 9 2 13 2
18 13 4 1 3 0 2 16 4 11 13 10 9 9 1 9 1 9 2
26 13 9 10 0 9 13 9 2 14 7 13 13 2 16 13 3 0 2 16 9 1 9 11 3 13 2
29 1 9 10 0 9 13 1 3 0 9 9 2 16 13 2 16 1 9 12 13 1 9 9 9 1 11 3 15 2
31 1 0 9 1 9 13 0 9 2 1 15 7 13 9 2 7 13 0 9 13 2 16 1 9 11 13 9 10 9 13 2
3 2 11 2
5 11 13 0 0 9
3 1 0 9
4 11 1 11 2
35 9 0 9 0 11 13 1 9 11 11 2 11 13 9 0 9 7 10 9 2 9 0 9 1 0 7 9 9 2 15 13 0 9 9 2
15 1 11 13 13 1 9 0 0 0 9 1 9 0 11 2
21 11 13 2 16 0 9 13 0 9 0 9 2 7 7 13 0 13 1 9 9 2
4 11 13 0 9
3 1 0 9
5 11 2 11 2 2
12 0 9 1 0 9 11 11 13 1 11 0 2
7 13 15 9 9 11 11 2
35 1 10 9 15 3 13 1 9 0 0 9 13 9 7 9 0 9 2 13 7 14 0 3 13 0 9 7 13 9 0 9 1 10 9 2
17 15 14 13 15 2 16 4 9 13 13 9 9 7 9 9 9 2
2 0 11
5 11 2 11 2 2
15 1 0 9 9 11 13 0 11 2 15 13 1 0 9 2
20 1 9 2 3 13 1 0 9 2 1 0 9 13 1 9 7 3 15 13 2
9 9 13 10 9 14 1 12 9 2
12 9 13 1 9 1 0 9 1 9 1 11 2
3 9 1 9
6 0 9 2 11 2 2
23 9 12 0 9 1 0 9 2 12 0 11 2 11 2 2 4 13 1 9 7 9 9 2
12 3 3 13 9 7 13 1 0 9 12 9 2
39 3 1 0 9 1 9 9 1 0 9 2 15 13 9 2 1 15 4 13 2 13 1 9 1 9 2 12 0 11 2 11 2 1 11 2 9 12 9 2
5 11 11 9 11 11
32 16 0 9 11 13 1 9 0 9 0 9 0 9 2 13 9 9 2 11 11 12 1 10 11 2 15 4 1 0 9 13 2
12 9 1 9 13 1 9 0 9 2 3 13 2
24 7 3 15 7 1 10 9 13 15 9 9 2 14 3 7 3 9 10 9 0 1 0 9 2
12 12 1 10 9 13 7 13 7 9 2 11 2
24 10 9 9 0 9 1 11 7 3 7 9 9 1 9 1 11 2 13 3 1 10 0 9 2
9 2 11 2 2 11 12 2 12 2
2 9 9
5 11 2 11 2 2
33 0 9 1 0 9 0 9 1 3 0 9 13 1 0 9 1 9 3 2 16 13 0 9 1 0 9 0 9 1 0 9 11 2
13 0 9 13 9 2 15 13 9 0 9 7 9 2
3 9 1 9
5 11 2 11 2 2
10 1 0 9 1 11 15 13 12 9 2
23 11 2 11 2 2 12 2 3 0 9 1 0 9 13 12 0 11 2 11 2 1 9 2
8 15 15 13 12 9 0 9 2
12 0 13 0 9 7 13 1 0 9 1 9 2
27 9 4 3 13 1 0 9 7 9 15 13 1 9 9 2 1 15 13 4 13 9 9 14 1 12 9 2
1 9
12 1 0 0 0 9 0 0 9 13 12 9 2
16 13 12 0 9 7 12 0 0 9 2 15 13 9 1 9 2
2 9 13
6 0 11 2 11 2 2
30 9 0 0 9 11 11 2 1 15 4 12 2 9 13 0 0 9 0 9 2 4 3 1 9 13 9 1 0 11 2
24 11 13 13 1 9 1 9 1 0 0 9 1 0 9 1 11 12 2 9 2 15 9 13 2
43 3 13 1 11 9 0 0 9 9 9 2 11 11 2 9 11 13 0 9 9 11 11 11 2 15 13 1 9 9 9 2 7 11 13 1 9 9 9 1 12 1 9 2
7 1 12 9 13 9 1 9
2 0 9
2 11 2
63 12 9 9 9 1 9 12 9 7 12 9 9 9 1 9 12 9 13 0 9 1 11 11 2 11 2 2 12 2 2 11 2 11 2 2 12 2 7 11 2 11 2 2 12 2 2 15 1 9 12 9 9 9 12 13 12 9 1 9 11 7 11 2
12 10 0 9 13 1 0 9 9 1 12 9 2
19 9 9 0 9 11 11 1 15 13 2 16 10 9 9 3 13 0 9 2
25 0 9 15 1 15 1 0 9 1 9 0 9 1 9 13 2 7 15 15 0 9 13 3 0 2
41 0 9 9 9 1 10 9 13 12 7 12 9 2 13 11 2 11 7 13 2 16 9 9 1 9 9 4 13 3 2 7 15 2 16 15 9 1 10 9 13 2
6 9 13 9 3 14 13
2 0 9
3 11 11 2
21 0 9 3 13 9 1 0 9 9 7 9 9 0 11 11 2 1 11 1 11 2
22 0 9 15 13 1 0 9 2 3 16 0 2 13 1 9 0 9 1 9 0 9 2
28 9 15 13 1 9 0 9 2 15 13 2 16 11 11 2 13 13 9 1 9 2 7 13 15 15 3 13 2
7 3 0 9 4 13 3 2
36 11 11 2 13 1 9 1 0 9 1 9 12 9 1 0 9 12 9 1 9 0 9 9 9 0 9 7 1 9 9 0 9 1 12 9 2
14 11 11 2 3 3 13 9 2 7 16 13 0 9 2
12 3 13 3 1 0 9 1 9 0 9 9 2
15 0 9 13 0 9 2 16 9 7 9 15 13 9 9 2
8 0 15 1 3 0 9 13 2
15 13 2 16 9 13 1 9 7 13 2 16 15 15 13 2
8 7 13 9 7 13 15 13 2
9 1 10 9 15 13 13 1 9 2
12 1 9 9 13 2 16 13 15 1 15 9 2
7 9 9 15 13 13 9 2
1 9
20 0 9 13 1 9 1 11 9 11 1 9 7 13 1 15 9 1 9 11 2
7 11 11 13 9 12 9 2
3 2 11 2
17 0 0 9 1 12 2 0 9 13 9 9 1 11 1 9 9 2
4 9 9 13 2
7 9 9 1 10 0 9 13
8 0 9 2 11 2 11 2 2
18 9 9 1 9 1 11 2 15 13 0 9 2 4 1 10 9 13 2
28 3 15 13 1 9 7 1 11 2 3 3 13 0 9 9 9 1 9 1 0 9 2 7 0 9 9 13 2
11 13 15 2 16 0 9 0 9 13 13 2
16 9 3 13 1 9 2 7 7 3 15 0 9 13 1 0 2
38 3 15 13 11 2 11 2 9 9 9 9 0 9 1 0 9 2 14 1 10 9 13 9 1 9 1 12 2 9 1 12 2 9 1 12 2 9 2
11 13 13 12 9 2 12 0 7 12 9 2
8 0 9 13 1 10 9 12 2
27 0 1 15 13 0 0 9 1 9 11 2 3 9 0 9 9 13 9 2 15 12 0 9 13 12 9 2
13 13 1 15 12 9 0 9 7 1 12 9 9 2
5 9 13 12 9 2
2 0 11
34 9 0 11 13 14 9 0 0 9 11 11 2 7 3 4 13 1 9 2 15 13 9 12 1 0 9 1 9 9 2 0 0 9 2
31 0 9 1 9 12 0 11 4 13 1 0 9 0 0 9 2 3 15 1 9 13 11 2 11 2 2 11 2 11 2 2
9 2 11 2 2 11 12 2 12 2
5 11 13 1 9 11
3 0 11 2
24 1 9 0 9 1 0 11 13 11 11 11 1 0 9 11 11 12 2 12 2 12 2 12 2
26 11 2 15 1 9 13 1 9 13 2 13 10 9 1 9 12 9 7 13 15 10 9 9 2 9 2
22 11 3 13 1 0 9 0 9 9 10 9 2 7 7 9 12 2 12 15 13 0 2
20 3 9 0 9 13 3 11 2 7 0 0 9 11 3 13 1 9 0 9 2
29 1 0 9 2 15 9 15 13 0 12 9 1 9 0 0 9 9 0 0 1 0 11 2 13 12 0 0 9 2
4 9 0 9 9
16 0 9 3 3 13 1 12 9 1 11 7 1 9 1 0 11
35 11 2 11 11 1 11 2 9 0 9 2 9 11 11 2 11 1 11 11 7 0 9 11 11 13 0 0 9 9 0 9 1 0 11 2
16 11 2 0 1 12 9 9 2 4 13 9 0 0 9 9 2
28 9 11 13 13 0 9 2 7 1 10 9 13 13 9 2 0 9 2 15 3 9 7 9 3 13 10 9 2
34 1 1 15 2 16 11 13 3 12 9 2 13 15 0 9 9 9 1 0 9 1 9 12 2 1 10 9 13 0 9 11 11 11 2
16 0 9 13 11 11 2 11 2 0 9 1 9 1 12 9 2
20 0 9 13 0 0 9 9 2 13 13 9 7 3 4 13 1 0 9 11 2
14 0 9 0 9 0 9 9 3 1 9 13 0 9 2
53 16 0 4 13 3 1 9 1 9 0 9 0 9 11 11 2 15 9 13 1 10 9 0 0 9 2 0 12 9 2 15 4 13 1 9 9 2 13 0 9 11 11 7 10 0 9 9 1 12 9 11 11 2
36 0 9 11 1 10 9 13 9 2 15 13 1 9 0 0 9 2 11 2 1 11 11 7 1 15 13 3 1 0 9 0 12 0 0 9 2
23 9 11 11 11 7 9 1 9 13 2 9 9 13 2 10 9 4 13 1 0 12 9 2
14 13 4 2 16 3 12 9 15 13 0 7 0 9 2
12 0 9 4 3 3 13 2 10 9 13 0 2
9 3 13 9 1 12 0 9 9 2
8 14 9 13 9 1 0 9 2
22 0 9 3 13 1 12 9 2 15 1 9 9 13 0 9 7 13 15 1 0 9 2
14 13 15 1 12 9 1 11 7 12 9 1 0 11 2
21 9 0 9 11 11 13 2 16 15 1 12 0 15 3 13 13 1 11 1 9 2
8 3 15 7 1 11 9 13 2
18 0 9 11 11 1 11 1 12 9 2 12 2 13 0 9 0 9 2
22 9 9 1 11 3 13 11 11 11 7 13 15 3 7 9 9 2 15 13 9 12 2
15 11 13 1 0 0 9 1 11 2 16 15 13 0 9 2
32 1 9 1 12 9 13 0 9 7 1 0 9 11 11 11 2 1 9 1 12 9 9 13 9 9 1 11 11 11 1 11 2
35 11 15 13 13 1 11 1 0 9 3 2 16 13 1 0 0 9 0 9 1 9 12 9 2 15 15 0 0 9 13 3 1 9 12 2
12 1 0 9 9 13 0 9 11 11 1 11 2
27 0 9 1 0 9 13 1 9 1 12 9 11 11 2 15 13 0 0 11 2 15 13 9 1 9 11 2
3 0 9 11
6 0 9 11 0 9 13
2 11 2
30 1 0 9 15 1 9 1 11 1 11 13 1 0 0 9 9 0 11 11 11 2 15 1 0 9 13 0 9 9 2
17 1 0 9 13 11 11 11 7 9 13 9 11 11 3 1 11 2
17 0 0 9 11 11 13 1 12 2 9 1 12 2 12 9 2 2
23 12 9 9 9 15 13 0 9 16 9 11 2 11 2 11 7 15 0 1 9 9 9 2
15 9 0 9 9 13 1 9 9 9 1 0 9 2 11 2
17 9 1 9 11 13 9 3 1 9 7 13 9 12 2 12 9 2
20 0 15 7 7 1 0 13 2 1 0 9 15 13 7 11 3 1 15 13 2
10 9 1 12 2 9 13 1 0 9 2
30 1 9 13 9 11 2 11 11 2 11 7 12 1 0 9 11 2 0 1 11 0 2 11 7 0 1 11 1 11 2
24 1 0 9 15 7 0 9 0 13 1 0 9 14 12 9 2 15 15 13 1 0 9 3 2
28 9 15 3 13 7 1 0 9 13 3 11 2 11 2 2 2 11 2 11 2 2 7 11 2 11 2 2 2
28 1 15 15 13 11 2 11 2 11 2 2 2 11 11 7 9 9 11 11 7 12 9 1 9 12 9 13 2
18 16 0 13 1 9 11 2 7 3 15 1 15 13 9 11 2 11 2
19 0 9 7 3 3 13 7 9 1 0 9 15 13 1 9 1 0 9 2
13 3 15 13 1 9 0 9 2 7 3 0 11 2
6 9 15 3 3 13 2
18 0 9 4 3 13 2 7 3 4 13 10 9 2 3 1 15 13 2
44 1 10 0 0 9 3 13 13 2 13 1 9 11 11 2 15 13 2 16 15 13 0 0 9 2 15 13 0 9 2 1 9 12 15 15 1 11 13 0 9 11 11 2 2
3 9 1 11
5 0 9 13 0 9
27 9 11 11 2 15 9 1 9 13 9 2 9 9 7 9 9 1 0 9 1 12 9 2 13 0 9 2
19 9 3 13 0 9 2 15 13 0 9 9 9 9 1 9 1 0 9 2
19 0 9 13 9 13 9 1 15 9 7 13 1 15 0 9 16 1 11 2
6 7 3 13 9 9 2
19 13 9 10 9 3 13 2 7 0 9 13 14 1 9 9 9 1 9 2
19 1 10 9 15 13 1 11 9 0 0 9 1 9 13 0 7 0 9 2
25 1 15 13 7 9 2 16 9 9 1 9 4 13 1 0 9 2 15 9 13 13 7 0 9 2
44 15 15 13 1 9 0 9 2 16 4 15 3 13 1 9 9 0 12 9 2 3 0 9 13 2 7 16 3 0 9 2 3 0 0 9 13 0 9 2 4 4 3 13 2
10 7 3 11 13 3 1 9 0 9 2
9 1 0 9 13 1 9 3 15 2
30 12 1 9 0 9 11 11 1 15 3 13 2 13 15 13 2 16 9 1 9 9 13 15 0 2 15 1 9 13 2
21 7 7 13 2 16 4 0 9 13 10 9 1 9 9 15 9 1 0 10 9 2
16 3 0 2 11 1 12 9 13 3 12 9 1 0 9 9 2
46 9 0 9 13 13 1 12 9 2 12 2 9 9 2 12 2 9 9 1 9 1 9 1 9 2 12 2 9 9 2 12 2 0 9 2 12 2 9 2 12 2 9 9 1 9 2
15 10 15 3 9 13 1 10 9 7 1 10 9 13 9 2
27 9 9 1 9 13 2 9 1 0 9 13 2 13 1 9 15 2 15 15 13 9 13 15 1 10 9 2
9 3 9 10 9 1 9 0 9 2
11 3 0 9 13 3 0 3 7 10 9 2
8 1 11 15 15 7 3 13 2
11 13 9 1 15 9 13 3 1 0 9 2
41 9 2 4 2 14 13 9 2 13 7 1 10 9 13 9 12 10 9 1 9 2 15 13 2 16 1 9 9 13 9 13 10 0 0 9 2 9 7 0 9 2
3 2 11 2
16 9 11 1 0 9 11 2 1 15 11 13 11 0 12 9 9
2 9 9
18 1 15 2 3 3 15 13 0 9 11 11 2 15 1 9 13 0 11
3 9 9 11
6 1 0 9 11 7 11
16 11 11 3 1 0 12 9 13 10 0 9 9 1 0 9 2
23 3 1 12 9 13 3 3 0 9 2 16 11 3 13 11 11 7 11 11 3 11 11 2
21 11 13 3 3 1 9 16 1 9 2 1 0 11 13 3 3 3 13 9 9 2
11 16 0 11 13 0 9 14 1 11 11 2
17 1 9 7 0 9 13 1 0 0 9 2 15 4 13 13 9 2
15 3 15 4 13 10 9 1 12 2 9 0 9 3 0 2
8 11 11 2 1 11 13 0 9
23 11 2 0 11 2 11 4 13 1 9 12 2 13 12 9 2 0 9 13 0 7 0 2
12 10 9 13 1 0 9 1 9 1 12 9 2
13 0 9 2 12 0 9 2 12 9 1 0 9 2
24 0 9 9 12 1 0 0 9 2 11 11 2 7 11 2 2 13 1 9 1 0 0 9 2
23 11 3 13 1 10 12 0 9 12 1 9 12 7 12 1 12 0 9 13 3 1 9 2
12 3 3 11 11 7 0 9 11 13 0 9 2
22 3 3 13 11 1 9 0 9 1 0 9 3 1 11 11 2 12 9 15 13 12 2
22 1 9 9 13 11 3 3 1 0 9 2 7 3 15 1 9 3 13 1 0 9 2
24 1 0 12 9 13 11 1 9 3 1 0 9 2 3 13 0 2 3 0 7 3 9 13 2
22 9 9 15 1 0 9 13 3 3 1 11 2 7 3 1 12 2 9 15 13 11 2
26 1 0 11 3 11 13 3 3 2 7 1 12 9 1 11 13 3 11 7 3 13 3 1 9 11 2
36 16 1 12 9 13 0 9 1 11 11 11 7 11 11 2 15 13 2 16 13 13 0 1 9 0 0 9 2 15 13 11 11 7 11 11 2
19 0 3 1 11 2 1 10 9 13 0 9 11 11 11 2 13 3 9 2
4 7 11 13 2
14 11 13 1 10 9 3 0 2 7 16 14 0 9 2
26 10 9 1 0 9 14 1 9 2 3 1 0 9 1 0 9 15 9 13 1 9 2 0 9 13 2
28 0 9 13 11 1 11 7 1 9 0 0 9 2 3 15 13 9 9 2 9 2 2 1 15 11 13 0 2
28 1 9 3 1 9 13 11 2 11 2 11 7 11 11 1 0 0 9 7 1 9 15 13 7 11 7 11 2
10 13 7 1 15 9 2 7 9 13 2
11 7 10 9 1 10 9 13 2 16 3 2
6 0 9 13 11 11 2
15 15 13 1 9 11 11 2 15 1 9 12 13 0 9 2
10 7 0 13 2 16 9 11 3 13 2
16 1 0 12 9 9 1 9 1 11 14 12 9 7 0 9 2
8 3 1 15 9 13 11 13 2
21 7 1 9 9 11 11 7 11 11 1 0 9 0 9 13 11 0 9 1 9 2
24 3 1 11 13 11 0 9 16 12 0 9 11 7 11 11 2 7 15 13 13 1 11 9 2
28 1 9 13 9 3 1 9 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2
15 9 9 13 1 0 9 2 9 9 4 13 1 9 9 2
19 1 0 9 15 13 13 9 0 9 2 15 11 1 9 11 13 7 13 2
16 11 13 3 2 12 9 2 0 9 13 7 12 0 9 11 2
20 9 11 13 12 1 11 9 1 9 7 9 13 1 0 0 9 1 12 9 2
11 1 15 1 0 0 9 13 7 11 11 2
8 11 11 2 0 9 1 9 9
22 11 11 4 13 1 9 12 2 0 9 13 0 2 1 15 4 13 7 9 0 9 2
25 9 13 1 10 9 1 9 1 11 11 1 9 12 2 1 15 12 9 0 2 0 9 12 2 2
17 0 9 2 12 7 9 2 3 13 0 9 2 9 9 7 11 2
26 0 9 11 13 1 0 9 1 9 12 7 1 10 9 13 1 0 7 0 9 1 9 9 1 0 2
27 10 0 9 13 12 9 1 9 0 9 1 9 12 1 9 0 9 2 3 13 3 0 9 7 3 11 2
40 10 9 1 0 9 11 16 9 13 3 0 9 1 0 9 14 3 2 3 13 1 11 16 0 9 0 9 2 12 2 12 1 11 0 2 15 13 9 2 2
10 0 0 9 13 1 11 0 16 9 2
12 1 9 9 13 10 9 3 3 3 1 9 2
34 3 13 1 9 12 1 11 0 2 2 12 2 12 2 2 3 1 9 12 1 11 2 12 2 12 2 7 1 0 3 1 11 0 2
25 9 1 9 12 13 0 2 1 15 13 14 0 9 2 7 16 10 9 13 13 3 1 9 12 2
31 1 9 1 9 1 9 12 13 11 3 0 11 0 1 11 2 11 2 11 2 11 2 11 2 11 2 11 7 9 11 2
13 0 9 13 1 11 12 2 12 7 13 15 13 2
22 0 9 15 13 1 11 0 2 1 0 11 7 11 13 9 11 7 11 12 2 12 2
5 0 13 9 11 2
21 1 9 11 3 11 13 11 11 12 2 12 3 1 0 9 1 9 12 2 12 2
7 12 9 15 13 1 11 2
39 1 0 9 10 9 15 1 10 0 2 0 2 9 13 9 0 9 16 3 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 3 2
33 1 11 2 11 2 11 7 11 3 13 3 3 0 9 16 11 11 2 11 11 7 3 11 11 2 15 13 3 15 0 0 9 2
41 0 9 9 2 12 0 11 11 2 13 11 1 12 9 2 13 1 11 2 1 11 2 7 11 2 1 9 1 11 13 0 9 1 11 2 15 13 1 0 9 2
26 7 16 13 9 1 11 2 13 1 9 9 1 11 1 11 2 3 13 0 9 9 7 7 0 9 2
13 1 15 13 9 11 1 9 9 9 1 0 11 2
19 10 9 13 3 3 0 7 13 13 1 9 10 9 2 1 10 9 13 2
26 9 9 10 9 1 11 13 11 11 2 15 13 9 11 2 16 11 13 1 11 2 16 13 1 11 2
10 1 11 13 10 9 13 0 0 9 2
15 3 15 13 9 2 16 9 1 11 13 0 1 9 13 2
17 11 13 1 11 3 2 3 1 11 2 3 13 1 9 0 9 2
22 1 12 9 11 11 13 9 2 15 15 15 13 13 2 16 3 10 9 13 9 9 2
12 7 0 9 1 0 9 9 9 1 9 13 2
26 9 11 15 13 0 9 2 16 13 11 0 2 15 12 9 7 3 3 2 3 3 13 12 2 12 2
8 1 12 9 9 13 11 11 2
25 11 13 9 1 3 0 0 9 2 7 3 13 3 13 16 10 9 2 16 4 15 13 1 9 2
36 1 11 13 0 9 16 11 2 11 11 2 2 11 2 11 2 2 0 11 2 11 2 2 11 2 11 2 7 3 11 2 11 2 11 2 2
83 0 9 11 13 11 11 1 11 0 2 1 12 9 2 9 2 3 13 9 11 11 1 0 11 1 12 12 9 2 0 9 11 11 2 0 9 11 11 2 7 3 9 11 11 1 11 1 12 9 2 9 2 15 13 0 9 2 1 0 9 3 13 12 9 2 1 11 1 11 2 2 9 11 11 1 11 2 11 11 1 11 11 2
14 9 9 13 3 11 2 15 9 13 9 1 0 9 2
14 13 1 11 2 11 7 11 11 2 7 12 7 13 2
16 9 11 7 11 13 11 9 2 13 1 15 9 1 0 11 2
13 1 9 1 11 2 11 4 13 11 9 1 9 2
34 13 13 12 2 13 15 12 2 0 9 11 2 9 11 2 11 2 2 11 2 11 2 2 7 3 12 11 2 11 2 11 2 11 2
21 11 4 3 11 13 1 0 9 16 9 2 16 1 0 9 11 4 13 1 9 2
13 9 9 13 0 9 11 11 2 15 13 1 11 2
4 1 9 13 9
7 11 3 13 9 0 9 2
9 13 15 0 11 11 11 1 11 2
29 9 0 9 11 11 11 11 3 13 10 9 1 15 1 9 2 7 3 1 9 1 9 15 13 13 12 0 9 2
31 3 13 1 11 1 9 2 1 11 1 9 12 2 12 1 10 0 9 12 9 13 2 3 15 13 9 7 0 9 13 2
7 7 11 13 1 10 9 2
17 11 13 9 0 9 11 1 9 12 11 2 15 13 3 9 11 2
24 1 9 15 13 1 9 0 11 7 1 9 2 16 13 2 15 13 9 1 0 11 0 11 2
10 1 10 9 1 12 9 13 12 9 2
16 3 7 11 13 15 2 15 13 1 12 9 11 2 13 11 2
17 1 0 9 13 11 1 9 0 0 9 2 16 4 15 13 9 2
22 11 2 9 2 11 11 2 11 2 11 11 2 11 2 15 10 9 15 13 11 13 2
25 11 7 13 1 0 9 2 15 3 1 10 9 13 10 0 9 2 0 9 1 9 12 9 9 2
6 15 7 3 13 3 2
17 11 13 1 9 10 9 2 3 3 11 2 1 15 13 0 9 2
24 13 15 1 11 11 2 3 13 1 9 1 0 9 11 7 11 7 11 2 11 7 3 11 2
25 15 15 13 11 16 0 9 2 15 3 13 2 3 0 0 9 2 15 11 13 9 1 0 9 2
14 11 15 13 2 16 10 0 9 1 11 4 13 11 2
23 15 1 0 9 2 9 2 9 7 9 13 3 0 2 7 3 3 0 9 1 0 9 2
10 11 13 11 1 0 0 9 1 11 2
11 7 15 4 10 9 13 2 13 11 9 2
20 3 2 16 9 1 9 11 13 3 11 2 15 1 15 3 13 12 9 9 2
13 0 9 13 1 10 9 1 11 0 11 11 11 2
11 15 15 13 1 0 9 11 0 2 11 2
12 13 15 2 16 13 3 2 13 9 11 11 2
12 13 15 0 9 7 13 15 1 15 13 3 2
6 1 11 3 13 4 2
15 9 1 11 13 1 0 9 1 0 11 0 9 1 9 2
14 7 15 13 13 9 2 3 13 1 10 0 9 9 2
10 1 10 9 13 0 13 1 0 9 2
8 1 0 2 11 13 3 12 2
6 1 15 11 7 11 2
20 7 16 13 1 11 2 13 15 2 16 3 7 3 4 13 9 10 0 9 2
6 3 0 9 15 13 2
5 13 3 0 9 2
8 13 15 12 2 10 9 13 2
4 13 9 12 2
8 0 12 9 13 11 1 9 2
16 13 15 3 3 2 16 4 13 1 9 16 13 11 7 11 2
7 13 4 10 9 1 9 2
7 7 3 4 1 15 13 2
11 7 1 10 0 9 1 9 11 13 11 2
17 9 1 15 3 13 16 1 0 11 2 16 1 0 9 0 9 2
6 7 13 14 12 11 2
21 13 4 13 0 16 15 2 16 4 9 13 3 13 2 16 3 13 14 12 11 2
3 2 11 2
1 3
9 11 11 13 0 9 1 0 11 2
15 9 9 0 0 9 11 1 0 9 15 13 9 11 11 2
16 1 0 11 13 0 9 9 11 11 11 1 9 12 2 12 2
24 0 9 9 0 9 0 0 0 9 2 11 2 11 11 11 13 1 11 1 9 11 10 9 2
22 0 9 11 11 13 1 11 3 10 9 9 9 1 0 9 0 0 9 2 11 2 2
3 11 13 9
2 11 2
24 0 0 9 7 9 9 1 9 1 12 9 9 12 0 11 11 11 13 1 9 1 0 9 2
30 0 0 9 2 15 13 10 9 1 12 9 1 9 9 2 13 3 1 9 3 1 9 7 13 15 0 16 1 9 2
14 13 4 15 15 9 13 7 13 4 1 15 0 9 2
27 3 13 1 15 16 3 7 13 15 2 16 13 13 9 1 12 9 7 13 7 9 0 9 2 13 11 2
34 11 13 0 9 12 1 9 12 7 10 9 15 13 13 14 1 12 9 3 1 9 9 0 9 1 11 10 9 11 11 2 12 2 2
14 11 13 0 9 1 9 12 1 11 7 12 1 0 11
5 9 9 9 1 11
6 9 13 0 1 10 9
2 11 2
20 0 9 11 11 15 13 9 0 0 9 9 9 2 0 9 0 9 9 9 2
39 0 9 1 11 13 3 1 10 9 11 11 1 9 12 9 0 9 9 12 9 1 11 11 11 7 12 2 12 9 2 1 0 9 11 11 2 11 11 2
29 1 0 9 9 13 7 3 1 12 9 11 7 13 1 0 9 13 0 9 9 9 2 15 3 1 10 9 13 2
13 13 15 0 9 10 9 2 13 1 9 0 9 2
8 13 10 9 13 9 0 11 2
44 9 9 1 0 9 11 11 1 11 1 9 1 0 9 13 3 1 0 9 1 9 12 2 12 9 2 2 7 1 0 9 9 15 13 0 9 7 13 3 9 1 9 9 2
50 0 9 11 11 7 11 11 13 1 0 9 1 0 9 12 2 9 1 9 12 2 12 9 2 7 10 9 1 9 11 11 11 11 7 11 11 13 1 0 9 12 2 12 9 2 1 12 2 9 2
19 1 10 9 9 12 0 9 1 9 11 11 12 11 13 0 7 0 9 2
4 9 11 1 11
9 1 11 13 3 3 1 9 1 11
2 11 2
10 0 11 11 15 0 9 13 3 13 2
16 1 0 11 2 0 9 1 9 11 2 13 1 11 11 11 2
16 12 9 15 13 1 9 1 9 9 1 9 1 12 2 9 2
11 1 9 9 11 13 9 10 9 1 9 2
12 0 11 4 13 13 3 1 0 9 1 11 2
34 3 13 1 15 9 1 9 9 7 9 1 11 3 2 0 9 13 9 0 9 2 13 1 0 9 1 9 1 0 9 0 9 11 2
11 1 15 0 13 1 0 9 9 1 9 2
25 11 13 9 1 9 2 11 0 9 2 11 15 3 13 1 9 1 9 7 1 11 15 13 9 2
13 1 9 1 9 9 11 13 2 13 9 13 13 2
15 9 1 11 15 13 2 9 13 13 9 1 9 0 9 2
2 0 9
5 0 9 0 11 2
5 11 13 9 1 11
9 11 2 11 2 11 2 11 2 2
21 9 0 9 13 1 12 2 9 0 0 9 2 1 9 9 7 1 0 0 9 2
7 3 15 10 9 13 11 2
24 11 2 15 1 0 9 13 1 11 2 13 3 1 9 11 2 16 13 1 0 9 0 9 2
13 9 9 13 9 11 1 0 9 1 9 1 11 2
14 9 2 11 2 11 2 11 2 11 2 11 2 11 2
14 9 2 11 2 11 2 11 2 11 2 9 2 11 2
3 1 0 9
13 0 11 11 13 11 11 2 15 13 1 0 11 2
9 0 9 1 15 13 12 9 9 2
14 11 13 3 0 9 0 9 2 15 4 1 11 13 2
5 11 13 1 0 11
3 0 11 2
19 0 0 9 7 9 0 0 9 11 13 1 10 9 9 1 9 1 11 2
32 0 9 0 9 15 3 13 1 0 9 2 16 10 0 0 9 7 0 9 11 11 13 0 9 7 9 4 13 3 12 9 2
36 9 9 11 11 11 13 2 16 7 1 12 11 9 1 9 13 2 3 13 2 16 1 0 9 13 9 1 9 0 9 11 11 1 11 11 2
36 9 11 13 2 15 4 13 9 13 1 9 9 2 15 13 13 14 1 12 9 2 7 13 0 2 16 11 13 0 9 1 9 12 9 9 2
13 0 0 9 7 4 13 13 3 16 1 0 11 2
22 16 4 13 13 9 1 0 0 9 2 13 4 4 13 9 14 1 9 12 9 9 2
1 3
27 9 9 0 0 9 1 11 15 1 9 1 0 9 13 1 12 9 7 1 0 9 13 0 1 12 9 2
12 0 9 9 15 0 9 1 10 9 13 12 2
18 1 9 15 9 9 0 9 13 3 1 12 9 7 3 1 12 9 2
26 1 0 12 9 10 9 13 9 0 0 9 9 12 2 15 13 1 12 9 3 16 1 0 9 3 2
14 9 9 15 9 15 7 13 1 12 9 1 12 9 2
26 9 9 0 9 11 2 11 1 11 1 0 11 13 3 0 9 16 0 9 9 9 10 9 1 11 2
12 0 9 13 3 12 9 7 14 12 0 9 2
17 9 9 0 11 13 12 0 9 7 0 9 1 0 9 7 9 2
30 9 0 9 11 2 12 9 2 15 1 0 9 13 1 0 9 2 15 3 13 10 0 9 2 16 13 9 3 9 2
18 3 16 12 9 9 13 0 0 9 1 9 9 11 2 11 11 12 2
17 13 15 7 14 12 0 9 2 1 10 9 15 13 1 0 9 2
8 9 13 13 9 1 12 9 2
13 0 11 2 3 2 13 1 11 1 0 11 0 2
7 9 9 13 12 2 12 2
2 9 11
5 0 11 13 1 9
11 1 0 9 11 13 7 0 9 2 9 11
2 11 2
15 3 12 9 1 0 9 1 11 13 0 9 9 0 9 2
19 0 9 2 1 0 11 2 13 1 12 2 9 9 3 11 12 2 12 2
13 9 13 7 9 11 2 15 1 11 1 9 13 2
20 9 9 15 13 0 9 11 2 15 1 9 12 2 7 12 2 9 13 9 2
16 9 11 12 2 15 9 13 11 7 11 2 13 3 1 11 2
15 0 9 9 13 1 12 2 9 11 2 15 9 3 13 2
21 9 1 9 11 13 9 1 12 2 9 9 1 11 2 12 2 12 2 11 11 2
32 10 12 0 9 13 1 9 1 0 11 2 11 2 1 0 9 13 1 12 2 9 7 13 9 1 0 9 11 1 0 9 2
2 11 2
21 0 9 9 11 1 0 0 9 1 11 13 14 1 12 2 9 0 9 11 0 2
11 0 9 9 13 12 9 1 9 9 11 2
31 9 2 15 15 13 1 0 9 0 9 11 2 15 1 0 12 9 13 12 9 2 13 0 9 1 9 1 12 2 9 2
10 1 9 1 9 11 7 11 13 9 2
21 1 9 9 15 13 11 0 2 15 13 11 2 7 1 0 12 9 13 12 9 2
30 13 15 7 0 9 11 11 2 0 11 2 15 13 1 9 11 12 2 12 2 16 3 1 12 9 13 12 2 12 2
15 11 13 1 0 9 14 12 9 2 7 1 12 13 3 2
2 11 2
27 0 9 9 11 2 11 11 11 11 13 7 1 12 2 9 0 9 9 2 16 13 1 11 12 2 12 2
35 1 0 9 15 13 13 0 11 0 2 11 2 15 13 1 9 0 9 11 11 11 12 2 12 7 1 12 9 15 13 1 12 2 9 2
9 11 13 11 9 12 9 1 12 9
4 3 13 12 9
7 1 9 1 9 3 14 11
2 11 2
14 1 0 0 9 13 0 0 9 0 9 12 2 9 2
19 11 15 13 12 9 1 9 1 11 2 7 1 0 9 15 3 13 9 2
28 0 15 13 1 9 9 2 7 10 9 13 13 0 0 9 11 1 11 11 2 1 12 9 1 0 9 2 2
14 3 9 13 1 0 9 9 7 16 0 9 3 13 2
15 11 13 10 0 9 9 12 2 12 1 0 9 1 11 2
15 0 14 13 1 9 3 0 0 9 3 1 0 9 9 2
11 3 0 9 11 15 13 2 7 13 11 2
6 0 9 13 11 11 2
23 11 3 13 1 11 12 2 12 2 7 12 9 1 9 12 9 13 9 3 1 9 11 2
6 11 2 11 12 2 12
18 13 15 9 9 2 16 0 11 13 9 1 9 9 7 0 13 9 2
4 7 11 13 2
15 7 3 15 13 3 1 0 9 2 7 10 9 13 9 2
6 3 0 13 9 11 2
12 1 12 2 9 9 11 1 9 13 9 11 2
21 1 12 2 9 15 1 9 11 1 9 13 11 7 3 13 11 2 12 2 12 2
10 0 7 1 10 9 13 10 9 13 2
29 1 12 2 9 15 11 3 1 0 9 13 9 2 9 11 13 3 9 0 11 2 16 11 13 2 12 2 12 2
14 1 0 9 0 13 1 11 2 7 9 9 15 13 2
14 13 15 14 1 12 2 9 2 3 1 9 11 13 2
15 0 9 0 3 13 3 7 3 11 12 1 0 9 13 2
16 11 11 2 9 11 2 3 0 0 9 4 0 1 15 13 2
11 11 11 2 9 11 2 11 13 3 3 2
14 13 4 13 0 9 2 15 7 13 1 0 9 11 2
3 2 11 2
6 11 2 11 12 2 12
16 11 13 0 2 0 7 0 2 0 3 13 14 0 9 9 2
18 1 12 2 9 13 11 9 1 0 9 2 7 9 13 1 0 9 2
15 3 15 13 1 12 9 3 11 2 16 13 0 9 11 2
20 1 9 13 0 9 1 0 9 1 12 2 9 2 7 11 1 0 9 13 2
17 12 9 1 9 13 1 9 9 11 3 11 7 13 1 15 13 2
21 3 15 9 13 1 9 2 13 11 15 9 7 0 9 1 12 9 13 0 9 2
18 11 13 9 7 0 9 2 3 13 1 9 11 2 15 7 11 13 2
26 3 9 3 13 7 9 11 15 14 13 2 16 15 1 9 11 7 1 9 7 11 13 9 1 9 2
18 1 12 2 9 3 11 13 9 7 1 9 11 15 13 12 2 12 2
13 14 1 9 15 13 0 9 0 9 1 12 9 2
18 1 12 2 9 11 13 1 0 9 0 9 2 7 13 14 1 9 2
12 3 1 9 13 11 7 11 13 9 1 9 2
4 9 2 12 2
4 11 2 12 2
4 11 2 12 2
2 9 2
4 9 2 11 2
18 9 2 11 2 11 2 11 2 9 2 11 2 11 2 11 2 11 2
4 9 2 12 2
5 11 2 11 2 2
4 9 2 12 2
6 9 2 12 2 12 2
24 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 12 2
11 11 11 2 9 11 2 9 13 12 9 2
16 16 4 13 1 12 2 13 4 0 2 9 4 13 1 9 2
18 1 9 4 15 7 13 13 2 0 9 9 13 7 15 15 13 13 2
14 11 11 2 9 11 2 13 15 0 0 9 0 9 2
20 9 16 4 13 13 3 3 16 1 9 1 9 2 3 4 13 1 0 9 2
3 2 11 2
8 0 2 11 2 11 12 2 12
14 1 9 1 0 9 1 11 0 9 11 13 1 9 2
23 1 9 15 13 11 2 1 9 0 11 7 1 9 13 11 2 15 13 1 9 1 11 2
20 0 9 13 0 1 9 2 3 9 9 13 3 1 15 1 0 9 9 11 2
19 1 0 9 13 1 9 0 11 7 3 13 9 11 2 15 7 13 11 2
9 1 12 2 9 13 11 11 9 2
9 15 13 1 3 1 9 0 15 2
19 11 2 3 0 0 9 1 9 11 2 13 9 7 3 1 9 13 11 2
24 1 12 2 9 15 0 11 13 0 9 2 11 7 10 9 1 9 13 7 0 11 13 9 2
12 11 3 7 3 1 15 13 2 0 3 13 2
4 9 2 11 2
16 11 11 2 9 11 2 9 3 13 9 2 9 9 13 0 2
21 11 11 2 9 0 2 11 2 9 13 9 1 9 2 7 1 9 15 13 9 2
11 13 4 3 9 2 13 0 9 1 9 2
9 11 13 2 16 13 1 15 9 2
3 2 11 2
6 11 2 11 12 2 12
14 0 13 1 0 9 2 0 0 9 7 9 1 9 2
19 1 12 2 9 15 15 13 2 11 3 13 9 11 2 15 3 13 11 2
21 1 9 0 9 15 0 13 2 16 11 15 13 12 9 1 9 12 9 1 9 2
28 1 12 2 9 3 13 0 0 9 7 13 2 3 1 9 1 9 15 13 0 0 9 7 0 9 13 11 2
21 1 9 9 9 13 9 1 9 13 3 9 2 13 15 12 0 9 11 7 11 2
8 1 12 9 13 3 9 11 2
10 0 15 9 9 13 1 0 9 11 2
11 12 0 9 11 7 12 11 7 11 13 2
7 9 2 12 2 7 12 2
4 11 2 12 2
2 11 2
4 9 2 11 2
16 9 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2
4 9 2 12 2
6 9 2 12 2 12 2
16 11 2 11 2 11 2 11 2 11 2 11 2 11 2 12 2
22 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 12 2
8 11 11 2 2 11 12 2 12
10 1 0 9 15 13 3 1 12 9 2
17 0 2 15 13 1 10 9 1 0 9 7 9 2 13 0 9 2
16 1 12 2 9 13 0 9 9 11 2 3 13 0 0 9 2
12 3 13 11 2 11 13 0 9 3 1 9 2
6 9 9 15 7 13 2
29 0 9 0 3 13 11 9 1 9 2 3 1 12 2 9 13 1 0 9 1 9 7 0 9 13 1 9 11 2
14 0 9 13 1 9 2 16 9 13 1 9 0 9 2
13 9 15 13 10 0 9 2 7 9 11 15 13 2
22 0 9 0 13 9 11 2 9 11 13 3 3 1 9 1 0 9 7 11 15 13 2
4 9 2 12 2
2 11 2
4 9 2 11 2
12 9 2 11 2 11 2 11 2 11 2 11 2
4 9 2 12 2
6 9 2 12 2 12 2
25 11 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 12 2
20 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 12 2
13 11 11 2 9 11 2 13 4 1 0 0 9 2
20 13 0 2 16 1 9 12 2 12 2 3 11 13 12 9 2 9 13 3 2
9 0 13 12 9 2 11 7 11 2
21 11 11 2 9 11 2 0 9 15 15 13 2 13 9 7 1 9 13 0 11 2
18 1 9 4 13 3 7 13 15 2 3 4 15 13 13 3 10 9 2
13 1 0 9 13 3 0 11 9 1 0 9 11 2
3 2 11 2
6 11 2 11 12 2 12
13 0 9 1 0 9 0 9 13 0 9 10 9 2
29 1 15 9 0 13 11 7 11 13 10 9 3 1 9 2 3 16 9 11 13 0 9 1 12 2 9 1 9 2
17 0 0 9 3 13 9 2 0 9 13 9 11 2 12 2 12 2
5 0 15 7 13 2
17 1 12 2 9 1 9 11 13 11 9 7 1 0 9 11 13 2
23 1 9 0 1 0 9 13 7 9 9 12 2 12 2 16 1 9 9 13 12 2 12 2
22 1 9 15 11 13 0 9 7 9 9 13 11 1 9 2 7 9 15 15 3 13 2
15 1 12 2 9 3 0 11 13 0 9 7 3 13 11 2
10 9 2 12 2 11 2 12 2 11 2
4 9 2 11 2
16 9 2 11 2 9 2 11 2 11 2 11 2 11 2 11 2
4 9 2 12 2
6 9 2 12 2 12 2
13 11 11 2 9 11 2 13 4 3 0 0 9 2
12 13 15 2 16 4 1 9 13 7 0 9 2
19 11 11 2 9 11 2 13 4 15 2 16 4 0 13 9 1 0 9 2
27 7 13 15 2 16 16 4 13 10 0 9 7 1 0 9 4 13 13 1 9 2 3 13 3 1 0 2
18 13 9 12 9 1 9 2 16 3 7 0 13 1 9 2 15 13 2
3 2 11 2
4 11 7 11 9
5 11 2 11 2 2
15 0 9 1 9 0 0 9 15 1 11 13 13 9 9 2
14 1 11 13 10 0 9 11 7 0 9 13 7 11 2
33 0 9 11 13 3 0 9 1 11 2 7 3 2 16 1 9 0 9 13 1 9 2 13 7 13 15 2 16 13 1 9 3 2
14 1 0 9 13 9 9 2 15 4 13 13 0 9 2
15 11 13 0 9 1 9 7 13 2 16 4 15 13 13 2
16 13 4 3 2 13 2 16 13 13 2 16 1 9 13 3 2
17 11 13 9 7 13 2 16 7 15 15 13 2 13 9 11 11 2
10 9 1 11 4 13 4 13 3 3 2
8 7 11 11 15 13 2 2 2
5 11 2 11 2 2
34 0 0 9 12 2 9 0 0 9 11 11 2 11 11 4 13 0 9 2 15 15 13 1 0 9 2 15 11 1 0 9 3 13 2
9 0 9 12 9 3 9 3 13 2
12 1 0 9 0 9 0 9 13 0 12 9 2
37 14 13 9 15 2 15 13 9 0 9 2 16 1 0 9 3 13 9 0 9 1 9 1 9 11 0 1 0 9 2 7 3 12 0 9 11 2
40 15 1 12 2 7 12 2 9 13 1 9 9 1 12 2 12 1 12 2 12 7 0 1 9 3 0 11 9 7 9 0 9 1 0 12 9 12 2 9 2
23 1 9 11 15 13 3 9 2 7 15 14 9 15 2 16 11 13 10 9 13 1 9 2
16 16 7 11 1 9 1 9 13 2 13 15 15 1 0 9 2
17 3 13 9 2 16 0 0 0 9 9 11 13 11 7 13 13 2
13 1 10 9 3 13 11 3 16 9 1 0 11 2
23 15 1 10 12 2 0 9 1 0 9 2 1 12 0 9 13 12 0 9 2 13 13 2
33 3 1 9 9 13 0 0 9 1 0 9 1 9 7 1 12 9 3 1 9 1 0 9 11 13 9 7 3 13 1 0 9 2
17 9 11 15 7 13 13 7 13 15 0 0 9 7 3 7 0 2
9 0 11 15 13 2 7 13 3 2
4 16 4 11 13
2 0 9
2 11 11
18 9 11 11 13 9 2 16 13 9 9 7 13 15 1 3 0 9 2
10 13 13 9 7 1 9 13 9 0 2
16 7 1 10 9 15 3 10 3 0 9 13 7 9 1 9 2
37 16 4 13 2 13 15 3 13 1 9 1 10 9 1 11 1 11 2 13 9 7 15 13 15 13 1 9 2 1 15 13 1 9 1 9 11 2
12 13 4 15 3 3 0 9 1 3 0 9 2
16 1 9 3 3 0 9 11 3 13 1 0 9 12 0 9 2
54 1 0 2 1 12 2 9 12 2 15 13 2 16 9 1 9 9 1 9 0 9 2 11 2 0 0 0 11 11 2 13 2 16 4 9 11 13 0 9 0 9 2 0 11 12 2 9 11 2 0 11 12 2 2
16 0 9 4 13 9 9 12 2 9 12 1 9 11 1 11 2
46 0 9 1 12 2 9 1 10 9 2 9 1 9 11 2 13 2 16 9 11 2 0 2 9 2 2 4 9 13 16 9 1 9 9 1 0 9 9 12 2 0 9 11 12 2 2
13 7 10 9 4 13 12 2 9 1 0 9 11 2
35 16 9 11 9 9 1 9 0 9 13 1 0 9 3 1 9 12 2 13 9 13 15 0 9 11 0 9 7 13 15 1 10 0 9 2
12 1 0 1 0 9 1 0 11 1 0 11 2
17 16 1 0 9 11 1 0 9 4 13 9 2 1 11 14 13 2
14 1 11 15 13 13 2 3 4 3 1 11 13 13 2
27 16 1 11 14 13 2 13 15 15 1 9 2 16 11 1 9 1 10 9 13 0 9 13 3 16 9 2
6 3 13 3 15 9 2
8 16 13 9 2 3 3 13 2
11 3 13 2 16 0 9 0 11 3 13 2
16 15 15 13 1 0 7 0 11 2 13 15 13 1 0 11 2
7 16 4 11 13 2 2 2
16 9 11 7 11 0 13 1 10 0 9 0 9 1 11 11 11
5 9 11 11 2 11
10 1 9 9 15 3 13 0 0 9 2
28 9 9 2 1 0 9 1 15 13 9 0 9 11 2 1 9 9 12 9 2 7 13 3 0 7 0 9 2
27 16 12 1 10 0 9 7 3 9 2 3 7 11 2 13 0 9 2 16 9 10 9 13 1 10 9 2
14 1 9 0 9 13 1 3 0 9 7 11 7 11 2
5 9 13 3 11 2
18 3 4 1 10 9 13 12 9 0 9 7 12 0 9 9 15 9 2
1 9
4 0 9 13 0
7 9 9 13 9 11 2 11
2 11 2
25 1 9 15 13 0 9 9 1 11 1 11 2 15 0 0 9 11 13 9 10 0 9 11 11 2
36 3 16 12 9 9 2 3 1 9 9 2 11 2 9 9 0 9 7 9 2 0 9 7 3 0 9 2 13 9 1 9 2 9 7 9 2
14 9 13 14 12 9 9 1 9 0 9 0 0 9 2
16 1 11 13 7 0 9 7 15 0 9 4 13 0 0 9 2
11 9 1 9 13 10 9 9 7 0 9 2
25 9 0 9 11 2 11 13 2 16 9 13 3 3 12 0 9 2 15 4 9 1 9 9 13 2
23 1 9 2 1 15 9 13 11 1 9 0 11 11 7 3 1 9 9 2 13 10 9 2
19 1 9 9 1 9 1 9 13 9 9 9 7 0 13 9 0 9 9 2
19 3 13 0 0 9 11 2 11 2 0 9 13 3 9 1 9 0 9 2
9 9 10 9 13 1 15 3 0 2
25 0 9 9 2 15 15 13 4 13 2 13 2 16 1 9 9 7 9 15 13 7 9 10 9 2
15 13 2 16 3 0 9 11 13 1 9 12 0 0 9 2
19 0 9 7 0 0 9 13 2 16 13 9 0 9 13 1 9 9 9 2
15 0 11 11 4 13 12 2 9 1 9 1 9 7 9 2
8 9 0 9 1 9 1 0 9
5 11 2 11 2 2
28 13 9 9 0 9 13 9 0 9 9 9 2 15 13 9 12 2 9 10 9 3 1 0 9 1 0 9 2
35 3 11 13 11 11 1 0 9 9 9 2 10 9 15 1 11 13 9 9 0 9 1 0 0 9 0 9 2 11 2 7 1 0 9 2
17 11 13 1 10 9 3 1 9 12 2 7 3 1 9 9 0 2
17 9 10 9 13 1 11 9 9 1 0 9 7 9 1 9 9 2
22 9 13 4 1 0 9 3 13 0 9 7 13 13 0 9 1 9 1 9 0 9 2
18 9 2 15 4 13 9 2 13 1 10 9 13 3 1 9 9 12 2
18 9 9 0 0 9 13 13 0 9 2 15 13 9 0 7 0 9 2
28 1 15 15 13 1 0 9 1 10 9 2 9 9 1 9 7 1 9 2 1 9 9 7 9 1 9 9 2
18 13 4 15 13 3 9 10 9 2 1 0 0 9 13 0 0 9 2
3 0 0 9
7 11 2 9 11 11 2 2
15 0 9 15 13 1 12 9 9 1 9 9 11 2 11 2
19 1 9 0 0 9 13 10 0 9 2 16 1 0 9 13 3 0 9 2
15 15 0 0 9 15 13 9 7 13 15 1 9 0 9 2
39 1 9 2 3 15 13 2 16 15 15 13 1 9 7 1 0 9 2 13 0 9 2 16 0 9 13 3 0 2 16 4 15 13 13 9 1 10 9 2
35 9 15 3 13 2 16 7 10 0 0 9 13 14 3 0 1 9 2 7 13 3 0 1 15 2 16 10 9 13 1 9 0 3 15 2
6 9 1 0 9 13 11
8 0 9 13 0 9 16 0 9
2 11 11
46 9 1 9 2 9 7 9 0 9 1 0 11 2 15 13 0 9 1 9 0 9 1 9 2 15 13 1 9 0 9 2 15 14 13 1 9 7 9 9 0 9 1 9 0 9 2
29 10 9 13 0 0 9 2 15 9 14 13 2 3 3 16 1 0 9 7 1 0 9 0 9 2 0 9 13 2
11 13 15 15 9 7 0 9 0 0 9 2
18 13 2 16 0 7 0 0 9 13 13 1 0 9 1 0 9 9 2
17 9 1 15 13 3 7 15 2 15 4 15 13 1 9 9 13 2
16 0 9 13 13 1 9 2 16 1 10 9 13 0 9 9 2
12 14 15 13 13 9 1 9 9 9 0 9 2
43 1 9 11 2 16 1 0 9 0 9 4 0 9 1 9 3 13 2 0 9 13 2 16 10 9 11 7 0 0 9 13 1 0 9 9 2 15 3 3 13 3 0 2
16 0 9 13 1 15 0 9 1 9 2 15 13 3 3 0 2
10 10 9 10 9 4 13 0 0 9 2
22 3 7 9 9 2 16 4 15 13 9 2 7 15 9 1 9 13 2 13 9 13 2
15 15 13 3 9 2 15 13 9 11 7 3 7 9 9 2
24 0 9 3 13 7 1 9 0 9 7 0 0 9 11 2 9 13 9 1 9 1 10 9 2
17 9 0 0 9 15 13 2 16 0 9 9 13 1 9 0 9 2
1 3
20 0 0 9 11 13 1 12 2 9 1 0 9 3 3 2 16 15 3 13 2
23 0 9 9 1 12 2 9 13 0 9 9 9 1 12 5 2 16 0 9 13 12 5 2
24 11 15 13 3 3 13 1 0 9 0 9 2 15 1 9 11 13 1 12 2 9 0 9 2
26 9 1 0 9 0 9 2 15 4 13 13 0 1 9 12 2 13 3 11 2 11 2 11 7 11 2
29 9 11 11 11 2 13 9 1 10 0 9 1 9 9 11 12 7 9 14 1 12 5 1 9 1 12 2 9 2
23 11 2 15 13 0 9 9 1 11 2 13 1 10 9 0 9 1 9 9 1 9 12 2
16 1 9 0 9 1 9 13 1 9 9 9 0 1 0 9 2
9 0 9 13 4 13 1 9 9 2
12 11 13 3 12 9 0 9 1 12 9 9 2
16 1 12 2 9 4 13 0 9 1 9 11 2 11 1 9 2
9 0 9 13 0 9 12 9 9 2
4 0 9 13 9
9 0 0 9 4 13 1 9 0 9
2 11 11
15 0 0 9 0 9 2 15 15 13 0 9 2 4 13 2
16 9 13 9 0 9 9 13 0 9 1 12 7 12 9 9 2
36 13 13 9 3 2 3 1 10 9 7 9 9 13 2 13 0 9 0 9 11 11 7 13 2 16 10 0 9 13 13 0 9 3 0 9 2
12 12 1 9 13 1 10 9 3 0 0 9 2
22 13 15 2 16 15 3 4 13 13 3 10 9 2 15 13 3 9 0 9 2 13 2
12 9 12 9 9 4 9 13 13 9 9 12 2
6 13 4 9 0 9 2
23 12 1 15 13 3 0 9 1 12 7 12 9 2 9 2 1 15 4 13 0 0 9 2
37 9 13 0 9 1 9 2 13 11 11 7 13 2 16 0 9 13 10 9 7 9 13 9 1 10 2 16 4 13 10 0 9 1 9 0 9 2
16 16 4 3 13 10 0 9 2 13 4 15 10 9 1 9 2
11 1 9 13 0 9 12 9 9 0 9 2
8 10 0 9 13 3 12 5 2
31 7 16 10 9 13 3 3 2 7 1 12 0 9 13 9 0 0 0 9 1 0 9 2 13 15 1 15 7 0 9 2
24 10 9 13 3 0 3 2 16 13 9 9 7 1 9 15 0 9 0 9 2 13 11 11 2
26 1 0 9 2 15 13 2 4 13 13 1 12 9 9 3 9 2 7 3 4 13 9 1 0 9 2
11 7 15 1 10 12 9 13 9 2 13 2
17 13 9 7 13 9 0 9 13 3 9 7 9 0 9 0 9 2
10 0 9 13 3 1 12 9 1 9 2
28 10 0 13 0 9 9 2 9 0 9 13 7 9 9 1 0 9 13 2 1 9 1 9 9 0 0 9 2
7 0 9 13 9 0 9 2
17 9 1 10 1 15 3 3 3 0 9 13 9 1 0 9 11 2
9 15 1 10 9 3 13 0 9 2
12 9 13 4 13 3 9 2 13 11 2 11 2
25 3 0 9 15 2 3 13 9 0 9 2 13 1 0 9 9 1 0 0 9 1 9 0 9 2
11 0 0 9 7 13 13 1 10 0 9 2
18 9 9 9 9 13 1 9 0 9 9 2 7 15 7 1 9 9 2
19 16 15 9 13 1 9 0 9 2 4 3 3 13 2 13 11 2 11 2
9 0 0 0 9 4 13 9 9 2
11 1 0 0 9 15 13 7 9 3 0 9
2 9 9
5 12 9 13 0 9
10 9 0 0 9 7 3 13 14 0 9
2 11 11
17 3 12 9 0 0 9 2 9 2 0 9 13 0 2 0 9 2
9 13 15 1 0 9 0 0 9 2
19 0 9 1 0 9 13 3 0 9 9 2 15 13 9 0 7 0 9 2
42 1 9 0 9 3 13 3 1 15 1 9 3 0 9 7 9 2 15 15 13 13 9 10 9 2 3 7 9 9 2 0 9 2 9 9 2 9 7 0 0 9 2
17 1 0 9 0 0 9 13 9 0 9 1 0 9 12 9 9 2
32 3 12 9 13 1 9 11 1 0 9 9 1 0 7 0 9 2 12 9 9 1 9 9 1 0 0 9 7 0 0 9 2
30 0 9 2 12 9 2 9 2 1 0 9 0 9 1 0 9 13 9 0 0 9 2 0 7 0 9 2 9 3 2
42 1 12 9 9 3 13 1 0 9 9 0 1 0 9 0 9 2 16 13 9 1 9 0 0 9 1 0 9 2 0 9 9 1 9 2 0 9 9 0 9 3 2
34 0 0 9 2 15 13 3 2 1 0 9 7 1 9 1 0 0 9 2 13 9 11 1 12 9 9 2 9 1 9 1 12 9 2
28 1 9 11 11 1 9 9 13 0 7 0 9 9 0 9 1 9 2 15 13 11 2 3 0 9 0 9 2
67 7 0 9 1 0 0 9 2 16 13 0 9 11 2 11 2 11 2 13 1 10 9 9 0 9 1 9 1 12 1 12 9 2 9 9 3 1 12 7 12 9 2 13 11 11 7 13 2 3 15 13 2 16 15 9 0 9 1 9 1 15 13 3 1 12 9 2
11 1 11 11 13 9 11 3 3 0 9 2
18 3 9 1 9 1 15 3 3 13 0 9 2 16 13 0 12 9 2
13 9 11 3 13 1 0 9 11 1 0 0 9 2
17 3 11 11 13 2 13 0 9 7 1 0 0 9 0 9 9 2
25 13 2 14 15 1 9 2 13 2 16 15 13 1 9 2 7 16 9 13 9 7 14 0 9 2
17 13 0 2 16 15 1 9 9 13 7 0 9 2 13 11 11 2
29 1 10 9 13 7 10 9 1 0 9 3 0 16 1 0 0 9 2 3 1 10 0 9 13 13 14 12 9 2
6 0 9 1 9 0 9
12 1 9 0 9 9 7 9 13 1 9 0 9
7 9 2 9 11 2 11 11
5 9 7 9 13 2
7 1 9 7 13 3 9 2
7 9 2 15 13 12 9 2
14 1 9 13 1 3 0 9 0 3 9 7 1 9 2
29 0 9 3 13 1 9 2 3 13 9 0 7 9 15 3 13 7 3 4 15 1 9 0 9 13 9 1 9 2
28 9 3 0 9 9 1 9 3 14 13 2 7 1 9 13 10 9 1 0 9 0 16 1 0 7 0 9 2
23 9 9 15 3 1 0 9 1 9 0 7 0 9 13 7 13 3 3 0 0 9 9 2
13 3 3 0 9 4 7 10 9 13 13 1 9 2
9 13 13 1 0 9 7 3 3 2
18 9 0 9 1 9 9 13 0 9 9 9 1 0 9 1 0 9 2
29 13 3 12 9 2 16 1 9 15 10 0 9 13 1 12 9 2 7 3 3 3 0 2 16 4 15 13 9 2
17 1 12 10 9 15 13 0 9 0 9 7 13 3 16 9 9 2
15 16 4 15 13 3 3 2 13 9 9 7 13 15 9 2
25 3 15 3 9 13 2 9 13 7 9 13 0 2 16 9 13 13 7 9 9 4 13 0 9 2
20 15 4 13 1 9 7 1 3 0 9 3 2 16 1 9 3 13 9 3 2
12 0 9 15 13 1 9 9 1 11 1 11 2
52 0 0 9 4 15 13 1 10 9 3 2 3 1 9 1 0 9 2 15 4 0 0 9 9 13 1 9 0 9 2 11 2 11 1 2 11 2 2 0 11 2 11 2 11 2 11 2 11 3 2 2 2
12 1 0 9 13 9 1 9 9 0 3 3 2
28 13 15 7 1 12 9 3 0 9 0 9 7 1 0 9 0 9 1 9 1 0 9 9 1 0 0 9 2
38 9 13 3 1 9 0 9 1 9 2 3 0 10 9 13 1 9 1 9 9 2 7 15 1 9 3 3 1 3 0 16 13 9 0 9 1 9 2
23 16 4 10 3 0 9 13 0 9 1 9 2 13 15 0 2 16 1 15 0 3 13 2
13 9 3 3 13 2 16 15 10 9 13 3 3 2
8 9 9 13 0 7 0 9 2
24 9 13 7 13 3 9 1 9 2 9 7 9 9 2 1 15 4 13 13 1 12 9 9 2
28 15 13 9 2 1 15 15 9 0 9 1 9 0 12 9 0 9 13 13 0 9 1 0 0 7 0 9 2
22 0 9 13 0 2 16 10 0 9 4 13 0 0 9 7 0 9 0 1 0 9 2
13 13 7 0 9 1 9 0 9 9 7 1 9 2
17 9 13 13 7 10 9 13 7 1 15 2 16 13 0 0 9 2
19 15 13 0 1 0 9 2 3 1 9 13 0 9 1 1 0 9 0 2
18 9 13 3 13 1 9 0 9 1 9 7 3 7 13 9 0 9 2
9 13 15 7 9 2 7 9 9 2
11 13 0 9 2 16 3 13 13 15 3 2
11 13 0 9 7 3 13 1 9 0 9 2
27 0 9 1 0 9 4 15 13 13 1 10 9 0 9 7 13 10 9 15 1 10 9 1 9 9 9 2
14 7 1 9 13 3 3 16 12 9 7 10 9 13 2
24 16 3 13 9 0 9 9 2 3 4 0 0 9 13 13 9 1 10 9 7 13 1 9 2
16 13 3 7 0 9 7 1 15 2 15 1 10 9 3 13 2
7 12 2 9 2 0 1 9
9 9 0 9 2 11 11 12 11 11
44 9 2 15 13 9 15 1 9 9 7 9 0 9 7 3 13 7 10 0 9 9 2 9 2 15 13 1 9 11 11 12 2 15 15 1 0 9 13 9 2 11 0 9 2
21 9 0 1 0 9 13 1 0 0 9 12 9 2 1 0 0 1 12 12 3 2
14 1 10 9 15 7 0 9 13 14 1 9 0 9 2
35 0 9 4 13 0 9 7 1 0 9 1 9 12 9 1 3 0 9 9 15 13 13 0 2 3 1 0 1 15 13 3 0 9 9 2
21 9 13 1 12 2 12 9 2 9 2 7 1 9 9 12 2 12 7 12 9 2
16 3 13 1 10 9 9 2 16 0 0 9 9 13 3 13 2
14 11 11 15 3 1 9 3 13 7 9 13 3 9 2
21 9 0 7 0 9 0 3 0 9 1 0 7 0 9 4 3 13 0 0 9 2
17 7 3 15 13 1 10 0 9 2 15 3 1 10 9 3 13 2
35 9 1 9 9 7 9 13 13 3 10 0 9 2 1 9 9 1 9 13 3 1 9 12 9 1 9 7 0 9 3 10 10 0 9 2
20 0 9 3 0 9 1 9 13 2 16 1 9 1 0 9 13 1 0 9 2
16 1 9 1 9 7 9 9 15 1 10 9 3 3 15 13 2
17 0 9 9 13 3 0 0 9 1 0 2 3 12 9 0 9 2
16 0 9 1 3 0 9 7 0 9 9 13 13 7 7 0 2
10 3 3 4 13 3 2 3 2 9 2
34 11 11 13 3 3 0 0 9 2 16 4 15 1 15 13 0 9 9 1 0 0 9 2 16 15 13 3 3 0 9 9 0 9 2
15 1 15 13 13 3 9 2 15 3 13 0 9 13 9 2
10 7 15 13 3 9 9 9 11 11 2
4 11 13 9 9
4 9 1 0 9
2 11 2
32 1 9 0 9 13 0 9 11 11 2 15 4 13 9 1 0 0 9 2 16 4 0 9 13 13 9 9 9 1 0 9 2
37 11 4 15 13 10 9 9 7 13 4 9 1 10 0 9 2 15 4 13 1 9 0 9 1 9 7 15 9 0 9 1 0 0 9 2 13 11
21 1 9 9 3 11 13 2 16 9 13 0 9 9 0 9 2 15 13 10 9 2
24 9 9 4 13 13 1 11 0 9 9 9 1 0 9 2 15 4 13 9 1 9 0 9 2
26 1 9 0 9 13 0 0 9 11 11 9 1 9 0 9 2 15 13 4 13 0 9 9 11 11 2
25 1 0 9 13 0 9 13 1 0 9 9 9 1 9 0 7 0 0 9 9 7 10 0 9 2
13 1 12 2 9 13 4 3 13 9 1 0 9 2
13 0 9 13 3 1 9 13 9 1 9 0 9 2
28 12 1 9 9 9 13 9 2 1 15 15 13 3 13 9 9 0 9 2 14 9 1 15 7 1 0 9 2
16 0 9 3 13 9 1 3 12 9 2 16 0 9 13 12 2
11 0 9 1 11 1 9 13 1 12 5 2
19 1 0 0 9 11 11 7 1 9 9 13 9 9 1 12 7 12 5 2
8 9 9 4 13 13 1 12 2
12 9 0 9 15 3 13 3 2 16 15 13 2
26 9 9 3 2 3 1 9 13 1 12 5 1 12 9 9 2 15 13 0 9 9 9 1 10 9 2
18 0 0 9 11 3 13 9 10 0 9 11 2 1 15 15 3 13 2
28 1 11 0 0 9 4 13 13 0 9 1 9 0 10 9 16 11 9 2 11 11 2 11 11 7 11 12 2
11 1 0 9 4 13 11 13 12 9 11 2
9 3 15 13 7 0 9 0 9 2
36 9 11 13 9 10 0 9 1 0 9 1 12 5 1 12 9 9 7 0 7 0 9 11 13 1 10 9 9 1 12 5 1 12 9 9 2
9 0 9 13 7 1 0 0 9 2
37 9 0 0 9 11 3 1 0 0 9 13 1 12 5 1 12 9 9 2 1 9 9 7 10 9 3 13 1 9 7 3 15 13 3 14 9 2
22 0 9 0 9 11 11 13 1 0 9 10 0 9 9 1 12 5 1 12 9 9 2
12 0 9 4 13 13 0 9 1 9 0 9 2
13 13 7 1 0 9 0 0 9 1 9 1 9 2
7 0 9 1 11 14 13 3
2 11 2
18 9 0 9 9 0 2 0 9 1 9 10 0 9 3 13 1 0 2
9 13 15 1 0 9 0 9 9 2
20 1 9 9 9 11 11 13 0 9 1 9 9 2 3 15 13 9 10 9 2
15 1 10 9 9 2 15 4 13 9 2 3 9 3 13 2
7 15 15 13 3 0 9 2
12 1 9 9 9 13 7 3 9 2 13 11 2
14 13 2 16 9 0 1 9 13 1 9 9 7 9 2
7 0 9 13 9 0 9 2
12 3 0 0 9 4 13 9 7 9 0 9 2
19 1 11 7 0 9 9 13 1 9 0 9 2 7 15 7 9 0 9 2
11 0 9 13 0 9 13 3 12 2 9 2
6 13 15 12 9 9 2
23 1 0 9 13 3 1 9 0 1 0 9 7 1 9 2 15 3 13 0 9 0 9 2
33 1 11 11 4 9 13 7 1 9 0 9 2 7 1 12 2 9 12 2 3 13 1 9 0 9 1 9 7 9 2 9 2 2
19 1 10 9 9 2 3 9 2 13 4 9 13 7 3 2 13 11 11 2
10 9 13 0 1 11 16 1 9 0 9
13 1 9 12 13 1 0 9 0 9 7 0 9 2
23 10 9 13 3 3 0 1 11 7 10 0 9 2 1 9 11 2 16 1 0 9 11 2
14 13 15 15 1 9 0 9 2 15 4 13 0 9 2
16 1 0 9 9 13 3 1 9 0 9 2 0 0 9 11 2
22 0 9 13 9 0 9 1 11 2 0 9 9 9 12 5 4 13 1 12 5 2 2
11 11 7 11 13 9 9 2 11 0 9 2
18 9 1 0 0 15 9 13 2 16 1 9 12 13 1 9 10 9 2
20 3 13 13 2 16 0 9 4 13 1 0 9 3 3 1 9 1 9 12 2
13 13 0 10 0 9 2 15 4 3 13 0 9 2
20 0 9 13 0 9 2 1 0 9 9 2 1 0 9 2 0 3 0 9 2
3 9 1 11
1 9
16 1 9 12 0 0 9 1 11 13 3 12 9 0 0 9 2
7 0 13 3 1 9 11 2
26 0 9 10 0 9 1 9 13 1 0 9 1 0 9 11 1 9 9 2 13 9 7 0 0 9 2
3 2 11 2
4 11 13 0 9
8 0 9 13 9 7 0 9 11
30 0 9 0 9 1 11 1 0 9 2 1 9 1 3 0 9 1 10 10 9 2 13 9 10 0 9 1 0 9 2
37 0 0 9 3 13 9 9 2 9 0 9 2 0 9 7 0 9 0 9 2 7 7 3 1 9 13 11 0 9 0 9 1 9 12 9 9 2
12 15 15 13 9 7 1 0 0 9 0 9 2
14 1 9 0 9 7 1 11 3 13 3 15 1 9 2
24 13 0 2 16 0 9 13 3 0 1 15 2 16 4 13 1 0 9 13 0 0 9 9 2
10 1 15 3 13 9 7 1 0 9 2
8 7 13 0 9 3 16 3 2
18 3 1 0 9 4 0 9 0 9 1 11 13 7 9 0 0 9 2
32 9 0 9 4 1 12 9 13 10 9 16 0 0 9 11 2 9 1 12 9 9 7 3 3 0 2 7 3 0 0 9 2
29 1 0 9 4 7 13 10 0 9 2 3 3 0 0 9 2 0 9 1 9 9 2 0 9 2 9 7 9 2
13 15 13 9 2 15 9 1 9 1 0 9 13 2
54 13 3 9 2 16 1 9 4 1 0 12 9 1 11 13 14 12 9 9 2 1 9 12 15 13 2 16 1 15 13 0 12 9 2 2 16 1 11 2 15 13 3 3 9 2 15 1 0 9 13 12 9 9 2
17 1 0 9 15 7 13 2 16 15 9 1 0 9 1 11 13 2
30 0 9 15 3 13 0 9 0 0 9 7 9 9 2 15 1 9 13 2 7 13 15 2 16 9 13 0 3 13 2
19 9 11 13 3 2 16 13 15 3 2 3 15 9 13 3 9 0 9 2
36 4 13 9 1 0 9 2 15 13 15 15 2 7 4 13 9 2 15 13 0 9 1 9 11 7 15 4 13 3 13 9 0 9 1 9 2
30 9 13 2 2 13 9 0 15 9 0 9 7 13 0 9 1 0 9 2 15 4 13 13 3 0 9 1 9 12 2
40 2 13 0 9 2 16 15 15 13 0 9 1 9 2 7 15 1 9 12 9 2 16 10 0 9 7 9 13 12 12 9 2 13 15 13 3 12 9 2 2
21 2 13 0 0 9 3 2 16 4 9 4 13 1 9 9 1 9 0 12 9 2
27 2 13 9 1 0 9 1 11 1 0 9 7 13 15 2 16 4 15 13 15 9 1 9 1 0 9 2
19 2 13 0 9 2 16 4 15 13 13 7 13 9 0 1 9 0 9 2
30 11 2 11 3 13 2 16 10 9 4 3 3 3 13 1 0 9 2 15 3 13 13 1 9 1 11 10 0 9 2
27 1 10 9 13 1 9 2 15 9 2 3 15 13 0 9 2 13 3 3 0 16 9 15 0 9 3 2
21 16 4 15 0 9 7 9 13 13 13 1 9 2 13 3 10 9 1 0 9 2
35 13 15 7 1 15 2 16 16 9 13 0 0 0 0 9 2 3 13 7 10 9 2 15 13 0 9 1 3 0 9 10 9 3 13 2
37 1 9 13 3 3 0 9 0 1 9 7 9 2 7 7 15 13 15 0 15 2 16 13 3 3 3 13 9 11 1 9 7 13 3 0 9 2
3 2 11 2
6 11 13 0 13 1 11
2 11 2
15 11 1 9 1 9 3 13 9 13 1 11 1 0 9 2
7 13 15 0 9 9 11 2
10 1 10 9 13 11 15 1 9 9 2
14 9 11 7 13 2 16 10 9 13 1 9 0 9 2
4 9 1 9 12
8 0 11 1 9 3 13 0 9
2 11 2
19 1 9 0 2 11 2 1 11 2 3 13 0 9 1 0 9 0 9 2
27 9 1 15 13 9 1 0 9 0 9 11 7 11 1 11 7 0 2 0 9 1 9 12 1 12 9 2
13 9 0 9 11 11 13 3 3 9 9 1 0 2
20 13 2 16 15 15 1 0 9 13 1 12 1 12 0 9 3 12 9 9 2
11 10 0 9 13 1 9 7 10 9 12 2
13 3 15 13 1 15 2 16 9 0 13 9 9 2
17 16 0 9 9 13 0 9 1 11 7 9 1 9 0 0 9 2
10 1 11 3 13 9 9 11 11 11 2
10 3 1 9 13 9 1 9 11 11 2
31 13 2 16 13 3 0 9 2 3 13 9 11 7 0 9 1 9 2 15 13 1 0 9 9 1 11 2 13 3 11 2
4 3 1 9 12
6 9 1 0 9 13 13
7 11 2 11 2 11 2 2
32 0 0 9 1 0 9 13 13 2 7 1 10 3 0 9 2 11 2 0 11 2 11 2 11 7 11 2 13 10 9 0 2
26 9 0 9 1 0 9 13 1 9 9 0 9 1 9 11 11 9 10 9 13 0 9 9 7 9 2
21 12 9 9 12 13 1 11 1 0 9 12 9 2 0 9 9 12 1 12 9 2
22 1 0 0 9 7 9 13 0 9 1 9 2 14 0 9 3 13 12 9 1 9 2
21 0 9 1 0 9 4 3 13 7 9 10 9 0 9 13 9 0 9 0 9 2
17 1 9 9 12 15 7 1 11 3 13 13 2 13 11 2 11 2
36 0 2 0 9 3 9 13 1 9 2 7 1 10 9 0 9 13 2 13 13 1 9 0 9 7 1 0 0 9 2 15 14 13 0 9 2
12 1 9 0 9 13 3 0 0 9 0 9 2
21 1 9 12 15 13 14 12 9 2 1 9 12 3 13 12 9 2 9 9 2 2
23 10 9 2 16 13 1 0 9 2 13 1 9 11 1 9 13 1 9 1 9 1 9 2
14 13 2 16 9 12 13 1 0 9 7 3 0 9 2
23 0 1 0 9 13 7 15 2 16 9 7 1 0 9 13 13 2 1 10 9 4 13 2
21 0 9 3 13 1 15 0 9 2 1 15 15 13 3 3 13 9 9 0 9 2
23 9 0 0 0 9 15 13 2 16 11 15 13 3 1 9 0 9 0 9 1 0 9 2
30 10 9 3 13 2 0 9 7 13 1 0 9 0 9 7 9 0 9 1 9 0 11 1 9 0 15 13 0 9 2
16 13 3 1 3 0 7 0 9 2 16 13 9 9 7 9 2
4 3 1 0 9
6 9 1 9 1 11 13
2 11 2
37 9 1 0 9 1 0 11 13 3 3 3 2 16 9 0 9 0 0 9 11 11 13 2 16 3 13 0 9 1 9 9 7 9 1 0 11 2
15 11 15 13 1 9 1 9 9 0 9 7 9 11 11 2
4 9 1 9 12
5 11 2 9 13 9
6 0 11 2 11 2 2
27 0 0 9 13 1 9 11 0 9 15 1 0 9 2 13 15 9 2 7 9 1 9 7 10 0 9 2
44 1 0 0 9 12 2 9 11 15 13 9 11 11 2 15 3 13 2 16 9 11 13 10 9 2 16 7 1 10 9 15 13 1 9 9 0 9 2 9 2 9 7 9 2
18 9 0 0 9 15 13 3 9 11 2 11 2 11 2 11 7 11 2
11 1 11 11 15 10 9 13 0 9 11 2
14 0 9 13 2 16 11 13 9 7 1 9 0 9 2
4 3 1 9 12
57 9 1 9 13 9 0 9 1 9 0 9 0 0 9 2 7 13 9 1 15 2 16 13 9 9 15 0 0 7 0 9 0 7 0 9 7 16 15 15 13 13 9 0 2 9 9 2 9 3 0 2 3 9 0 2 0 2
7 9 11 2 11 1 9 12
5 13 15 0 0 9
2 11 11
11 9 11 11 13 11 9 1 9 0 0 9
11 10 9 13 0 7 0 9 1 0 9 2
7 0 9 13 9 0 9 2
20 3 1 9 4 13 13 1 9 9 0 9 7 9 9 1 0 9 7 9 2
25 15 13 3 2 9 1 9 9 9 2 16 9 7 9 9 4 13 0 9 13 10 9 7 9 2
9 3 4 13 9 3 0 0 9 2
12 13 2 14 0 9 2 3 1 15 3 9 2
11 16 10 9 13 9 7 13 15 13 3 2
10 3 13 3 0 9 1 9 0 9 2
22 9 2 15 4 15 13 13 1 9 2 3 4 13 0 9 2 16 13 3 0 9 2
19 15 13 0 0 9 7 1 15 4 15 13 13 13 7 0 9 0 9 2
16 9 3 3 3 13 9 2 16 9 15 3 4 13 13 9 2
7 13 2 16 13 1 9 2
24 1 0 9 4 9 13 10 9 9 1 0 9 7 7 3 3 4 13 9 1 3 0 9 2
15 1 15 13 9 2 16 15 9 13 13 0 9 1 15 2
31 0 9 13 3 9 1 15 2 16 4 3 9 13 0 9 1 0 9 2 15 4 15 13 13 1 12 9 0 1 15 2
17 3 2 3 13 13 0 9 7 9 2 16 4 13 9 1 9 2
5 0 13 0 9 2
18 16 13 2 16 13 9 14 1 9 1 9 2 0 9 15 3 13 2
9 0 4 7 13 1 0 0 9 2
12 1 10 9 7 13 3 1 9 1 9 9 2
11 3 0 9 13 3 9 0 2 0 9 2
17 14 2 1 10 0 9 13 1 15 3 9 2 3 0 0 9 2
5 7 3 15 13 2
35 13 15 9 2 3 13 0 9 3 0 9 0 3 14 9 2 7 13 15 3 9 1 0 9 9 2 9 2 7 7 0 15 9 9 2
27 16 3 15 1 0 9 13 14 9 0 0 9 2 3 2 3 13 9 9 9 2 15 9 0 9 13 2
16 16 4 13 13 9 1 9 2 13 4 9 0 2 7 0 2
17 3 4 15 13 1 9 9 2 7 3 1 15 2 15 15 13 2
23 1 11 3 13 3 0 0 0 9 2 1 9 9 4 3 1 12 0 9 13 0 9 2
38 13 4 2 16 4 15 9 2 1 9 2 16 4 13 0 2 13 3 3 1 0 9 2 7 4 13 9 15 2 16 4 13 0 9 3 0 9 2
29 16 4 13 9 2 10 9 13 0 9 1 9 9 15 9 3 12 9 7 9 2 14 4 13 0 9 7 9 2
3 12 9 11
2 11 11
10 0 0 9 13 9 0 1 15 9 2
9 3 15 13 11 0 9 13 15 2
14 13 15 3 1 9 2 7 13 7 9 1 10 9 2
9 7 1 9 15 9 11 13 3 2
29 13 15 3 3 3 2 1 0 9 0 9 1 11 2 16 3 13 1 15 2 13 2 14 1 11 7 1 11 2
16 1 9 0 0 9 1 9 15 13 9 7 1 0 0 11 2
5 13 15 0 9 2
22 3 3 13 0 9 2 15 13 9 0 9 11 11 2 9 1 11 2 0 0 9 2
24 10 0 9 13 13 9 2 15 3 13 0 9 16 9 9 0 9 13 15 9 9 1 11 2
20 7 3 1 10 9 13 9 0 0 9 1 0 9 2 16 9 13 11 9 2
19 0 0 9 13 0 9 2 13 1 9 1 9 7 13 15 1 0 9 2
8 3 7 3 1 9 9 0 2
32 1 12 9 4 3 3 13 2 11 7 3 13 4 13 1 0 9 2 16 1 9 0 0 9 13 1 9 9 12 0 9 2
26 1 9 3 13 0 13 7 0 9 0 9 7 1 15 0 9 1 9 0 2 0 9 1 0 9 2
9 1 15 7 9 11 13 0 9 2
39 3 1 9 12 2 3 0 0 9 4 11 13 1 0 9 7 1 0 0 9 13 14 9 2 3 1 12 9 3 2 3 1 9 13 14 3 0 9 2
22 13 2 14 0 9 9 1 0 0 9 2 13 0 2 16 15 11 13 7 9 0 2
7 3 0 9 1 9 0 9
6 11 11 2 11 2 2
20 9 9 13 1 9 1 0 0 9 11 12 2 9 0 9 0 9 11 12 2
30 9 13 12 0 9 10 9 2 11 11 1 9 0 9 1 9 13 0 9 7 9 11 11 7 11 11 1 9 0 2
21 9 1 9 1 11 2 11 13 0 9 9 1 11 2 0 11 2 11 7 11 2
30 3 15 13 9 0 9 11 11 2 15 3 13 0 9 2 7 3 0 9 1 0 9 2 13 9 11 9 0 9 2
13 1 0 9 0 9 15 9 13 0 9 0 11 2
1 3
16 9 9 1 9 3 13 0 9 1 11 2 15 13 3 0 2
17 1 12 9 15 3 13 12 0 9 2 1 15 13 12 9 13 2
23 0 9 1 9 0 9 3 1 9 1 11 13 2 9 11 11 15 13 1 9 9 12 2
18 9 0 7 0 9 2 0 0 0 9 11 2 13 1 9 1 11 2
10 13 15 15 12 9 0 9 7 9 2
14 0 9 11 11 13 1 9 12 9 1 11 1 11 2
16 11 2 15 13 0 0 9 1 11 2 13 9 9 7 9 2
9 0 0 9 4 13 3 0 9 2
16 0 9 1 9 0 9 11 7 11 13 1 9 1 12 9 2
12 13 15 1 0 9 0 9 11 1 9 9 2
27 12 9 1 0 11 13 1 9 1 9 1 0 0 9 1 9 9 7 9 9 11 1 11 11 2 11 2
13 3 0 9 13 9 9 1 9 0 9 10 9 2
2 13 9
2 11 2
26 9 0 9 0 4 1 9 1 11 1 0 12 9 13 11 11 2 0 9 1 0 9 0 2 11 2
12 0 9 1 9 3 13 9 9 7 0 9 2
11 0 9 9 0 9 13 14 12 9 9 9
5 11 2 11 2 2
21 0 9 0 9 0 9 9 2 15 13 9 9 2 4 13 4 3 7 3 13 2
6 15 9 13 4 13 2
13 13 15 1 9 11 11 1 0 0 9 1 9 2
18 10 9 13 0 2 9 9 1 0 9 0 9 0 15 9 1 0 2
10 1 11 13 10 9 1 9 1 11 2
12 9 15 3 13 3 3 13 9 1 0 9 2
17 9 13 3 0 15 15 1 15 13 2 7 0 0 9 3 13 2
21 13 1 15 7 1 0 9 0 0 9 2 0 2 0 9 2 13 11 2 11 2
13 1 9 13 13 9 2 10 9 13 7 3 0 2
23 9 1 9 13 3 0 9 9 2 7 13 15 7 1 0 9 0 1 9 0 0 9 2
19 9 9 9 13 3 9 9 2 7 9 15 0 9 2 15 10 9 13 2
27 1 11 2 11 9 0 0 9 9 13 2 15 4 13 4 13 2 7 7 15 3 13 9 1 0 9 2
16 13 15 2 16 0 9 9 0 9 13 14 12 9 9 9 2
3 0 9 9
5 11 2 11 2 2
19 3 0 9 1 11 15 1 9 13 1 0 9 9 0 1 11 1 11 2
30 10 9 13 9 0 2 11 2 11 11 2 2 15 13 9 0 9 7 0 9 0 1 15 1 9 0 9 7 9 2
18 1 0 9 3 1 11 13 12 0 9 7 9 1 9 3 12 9 2
4 9 0 0 9
5 11 2 11 2 2
23 9 12 9 2 15 13 1 0 0 9 1 9 0 9 2 13 1 9 1 11 1 11 2
40 9 0 9 0 9 1 0 9 2 16 13 13 1 0 9 9 9 0 9 9 7 1 0 0 9 9 2 13 3 2 16 1 9 13 3 9 12 2 12 2
29 9 9 11 1 11 2 1 11 7 1 11 11 11 13 9 11 2 16 9 0 9 13 3 9 9 1 0 9 2
13 0 13 2 16 1 12 9 13 9 9 3 0 2
23 9 11 16 0 9 12 9 1 9 13 1 11 9 9 0 9 2 15 13 0 9 11 2
18 1 9 1 11 13 9 0 9 1 11 2 0 9 13 7 0 9 2
27 11 13 1 9 11 1 9 12 11 2 9 11 13 14 1 9 12 2 3 3 1 9 12 1 9 12 2
14 0 9 4 13 3 1 12 9 1 11 2 3 3 2
3 0 0 9
5 11 2 11 2 2
33 0 12 9 9 11 2 15 15 1 11 12 2 9 1 9 0 9 11 2 11 13 0 9 2 13 0 9 9 1 0 9 9 2
8 9 0 15 3 13 1 12 2
6 3 0 9 13 9 9
12 1 9 9 9 13 0 3 13 0 0 9 2
6 0 9 3 13 12 9
12 11 11 2 0 9 9 0 9 2 0 0 9
8 9 4 13 16 9 0 9 2
10 0 9 2 9 0 9 2 13 9 2
10 9 13 2 13 2 14 0 0 9 2
24 1 9 9 4 13 0 9 2 3 9 0 9 2 15 13 9 0 0 9 0 9 7 9 2
13 1 9 13 13 2 16 9 9 13 9 9 9 2
5 9 9 1 9 9
24 0 9 0 9 13 13 9 2 15 13 9 0 9 9 1 9 2 3 9 7 1 9 9 2
9 15 13 0 13 1 9 0 9 2
67 9 9 9 7 9 15 13 9 0 9 9 2 15 13 10 9 2 3 1 9 15 9 0 1 0 3 0 9 9 2 3 0 9 2 15 13 9 9 10 0 9 12 7 3 10 3 0 9 2 3 2 9 16 9 0 0 9 7 0 9 16 9 0 0 9 2 2
36 0 9 15 3 13 9 0 9 2 9 2 9 0 15 0 9 2 3 2 0 9 2 7 9 2 3 2 0 9 0 7 0 9 0 2 2
37 0 9 0 9 1 0 9 9 7 9 1 9 3 1 9 7 1 10 0 9 13 3 0 9 0 9 7 9 1 0 9 2 0 9 2 9 2
15 9 15 9 13 0 2 0 9 2 15 13 9 15 9 2
41 0 9 2 9 2 12 9 2 3 0 9 2 1 0 9 13 13 3 0 1 0 9 7 10 9 3 3 2 16 13 13 1 9 0 0 9 2 9 2 9 2
12 1 10 9 13 3 0 9 9 1 0 9 2
2 0 9
21 1 9 9 9 7 9 13 0 3 13 1 9 9 2 1 15 4 0 9 13 2
20 0 7 3 0 9 15 13 1 0 9 2 9 2 9 2 9 0 2 2 2
22 3 15 3 1 9 0 9 0 9 13 1 3 12 0 9 12 0 9 1 12 9 2
21 9 0 9 7 2 0 9 1 0 9 9 0 9 13 9 0 9 1 9 12 2
3 9 9 9
53 16 4 13 0 13 3 0 2 0 0 9 1 9 9 9 2 13 0 13 1 9 9 9 9 9 2 15 4 1 9 13 9 9 1 0 9 2 9 2 9 9 2 9 2 9 7 3 9 0 7 0 9 2
14 13 9 9 13 0 3 1 0 9 9 9 7 9 2
31 7 15 13 0 9 2 15 13 2 16 15 13 9 2 15 15 3 13 7 15 13 0 2 0 9 3 3 0 1 0 2
10 1 9 9 9 13 13 3 0 9 2
16 0 9 9 13 16 13 2 7 13 1 9 0 9 0 9 2
28 13 2 14 1 0 9 0 9 2 9 2 16 13 9 2 9 2 9 2 9 3 2 13 13 9 1 0 2
37 3 13 2 14 1 0 9 9 2 15 13 7 13 0 9 9 2 13 15 9 9 0 1 0 9 3 1 9 0 0 9 2 9 7 9 2 2
37 0 0 9 13 1 10 9 9 1 0 9 3 10 9 2 15 15 1 0 2 0 2 13 0 2 0 2 2 16 13 15 1 9 2 9 3 2
31 9 0 9 13 1 9 0 9 9 9 7 0 9 0 9 9 2 9 2 0 3 0 9 1 15 3 0 9 9 9 2
75 9 9 7 9 0 0 9 13 0 0 9 2 15 15 13 3 1 12 2 12 9 7 13 9 0 2 0 9 0 9 2 15 3 13 9 0 0 9 2 9 9 7 9 9 2 0 9 9 7 9 2 2 9 0 9 2 9 0 7 0 9 7 3 9 0 7 0 9 1 9 7 9 0 9 2
13 1 9 9 9 0 9 15 3 13 9 0 9 2
38 1 3 0 12 9 2 7 2 0 9 1 9 0 9 7 9 9 1 9 0 9 4 0 9 13 3 1 9 9 7 10 9 3 0 9 0 9 2
7 10 9 3 13 0 9 2
4 9 9 0 9
29 1 9 9 13 0 3 13 0 0 9 2 0 0 9 2 0 9 2 0 9 2 0 9 2 2 1 15 13 2
26 0 0 9 13 0 0 9 9 2 15 13 9 0 0 9 1 9 0 12 9 1 9 12 0 9 2
23 10 0 2 0 9 13 9 0 9 0 1 0 9 7 1 0 9 9 7 9 0 9 2
22 9 0 9 9 13 2 10 9 13 0 9 1 0 9 0 9 1 0 9 0 9 2
22 3 4 13 9 16 9 0 9 0 9 1 9 9 0 2 9 0 9 5 12 2 2
25 10 9 13 9 9 9 1 9 0 9 7 1 9 0 9 13 0 1 0 9 1 9 0 9 2
18 0 9 13 9 0 9 2 15 13 9 0 9 0 9 1 0 9 2
6 13 0 9 9 9 2
4 9 13 0 9
12 1 11 13 3 12 7 12 9 0 9 1 9
5 11 2 11 2 2
38 1 0 9 4 10 9 9 1 9 0 9 13 1 0 9 9 1 9 9 1 9 1 0 9 2 3 0 9 1 9 9 1 9 0 7 9 0 2
24 3 13 9 0 9 9 9 0 9 9 9 11 11 2 13 3 1 0 9 9 1 9 9 2
18 9 9 0 9 13 1 11 9 1 10 2 15 13 13 1 0 9 2
43 13 7 2 16 10 9 2 15 13 9 13 7 13 1 9 2 13 1 0 9 9 3 13 1 9 0 9 7 1 9 15 13 14 1 0 0 9 9 7 9 0 9 2
37 0 9 0 9 13 1 0 9 9 2 1 0 7 0 9 13 13 1 11 0 0 9 0 9 2 3 2 1 9 2 10 9 15 13 1 9 2
32 9 9 9 1 9 0 9 0 9 1 0 2 9 2 11 11 11 11 13 2 16 3 12 7 12 9 0 9 13 1 9 2
8 1 0 13 0 13 0 9 2
15 15 13 1 0 9 13 0 9 0 9 1 12 12 9 2
16 0 9 3 13 2 16 15 0 9 3 13 16 9 0 9 2
12 0 9 13 7 9 0 0 9 1 0 9 2
23 1 11 3 13 9 9 0 9 9 7 0 9 2 3 0 9 0 9 2 15 3 13 2
23 1 9 0 9 1 0 9 13 0 9 9 13 7 10 9 2 15 15 13 1 10 9 2
19 0 9 9 0 9 4 13 2 3 13 11 2 0 9 0 3 1 9 2
4 0 9 0 9
5 11 2 11 2 2
34 12 12 9 0 0 9 2 12 7 9 9 9 2 1 9 1 9 9 9 13 1 9 1 9 9 0 9 9 1 9 7 0 9 2
42 1 10 9 11 11 4 9 13 1 0 9 12 9 1 9 3 1 9 7 1 9 1 12 1 12 9 1 9 0 2 9 2 11 2 0 12 2 11 12 2 11 2
36 3 4 1 11 13 3 16 12 12 12 9 16 9 1 9 0 9 2 15 15 13 1 10 0 9 2 7 3 9 7 9 0 9 2 13 2
13 9 1 9 12 9 9 4 13 1 0 0 9 2
27 1 9 13 13 12 7 9 9 9 1 15 0 9 1 9 2 9 2 9 2 9 2 9 7 0 9 2
20 1 0 9 13 1 9 1 9 0 9 0 9 9 7 0 9 9 2 12 2
29 1 12 9 0 9 13 9 0 9 7 9 2 1 15 13 3 0 9 11 11 7 0 0 2 0 11 11 11 2
18 9 13 9 7 0 9 11 11 2 0 9 2 12 15 13 1 9 2
3 2 11 2
5 9 11 11 2 11
4 0 9 13 9
5 11 2 11 2 2
48 1 9 0 9 0 9 1 0 9 11 11 7 0 9 11 11 4 1 9 1 0 0 9 0 11 1 0 9 3 13 9 1 9 0 0 9 7 0 9 0 11 11 11 2 0 9 12 2
22 0 9 4 13 3 1 9 1 0 9 2 3 15 13 0 9 1 9 9 9 12 2
24 1 9 1 9 4 13 3 1 9 9 0 9 9 1 0 9 7 0 3 9 9 1 15 2
24 0 9 9 11 2 15 13 1 0 9 7 9 10 9 2 13 9 2 11 11 1 0 9 2
25 15 9 11 13 2 9 13 0 2 14 12 9 0 9 2 3 0 7 1 9 13 10 0 9 2
14 13 15 12 9 7 1 10 0 9 15 3 13 9 2
3 9 1 9
2 11 2
42 9 0 9 2 10 9 2 9 9 0 0 9 7 0 9 9 1 0 9 4 1 9 1 9 1 0 9 13 1 0 9 1 10 0 9 1 11 7 0 9 11 2
27 14 15 0 9 7 13 0 9 3 3 0 9 2 7 13 1 9 9 9 1 9 7 1 9 10 9 2
15 9 11 13 1 10 9 9 1 0 9 1 10 0 9 2
18 0 9 1 9 0 9 13 9 9 0 0 9 9 1 12 2 9 2
31 9 0 9 0 9 2 15 15 13 12 2 7 12 2 9 2 13 9 1 9 1 9 1 9 1 12 2 9 0 9 2
14 1 15 13 4 9 0 9 13 1 9 12 2 9 2
7 9 9 9 13 9 0 9
5 11 2 11 2 2
27 0 0 9 3 13 9 0 0 9 2 15 13 13 0 9 2 7 1 9 9 4 15 13 13 9 9 2
22 1 0 0 9 9 15 1 9 1 9 11 11 11 13 9 9 11 11 2 11 2 2
27 1 9 9 9 15 1 15 4 13 3 3 1 9 0 9 1 0 9 2 7 0 9 9 3 11 13 2
16 9 11 11 2 11 2 13 2 16 0 9 13 13 3 3 2
11 1 0 9 0 0 9 13 9 0 9 2
20 3 13 2 3 1 9 4 13 13 9 0 9 2 15 4 13 9 0 9 2
19 0 9 2 3 9 1 9 1 0 13 14 9 2 1 11 13 3 0 2
36 9 11 11 2 11 2 15 13 2 16 1 9 0 9 15 1 9 13 12 0 9 2 3 0 9 2 15 13 9 2 7 3 0 9 9 2
9 9 15 13 13 3 2 13 11 2
22 1 9 11 3 9 1 9 13 2 7 13 3 0 2 7 15 9 13 15 3 13 2
10 13 2 16 9 9 13 1 9 13 2
5 9 1 9 13 13
9 9 11 11 15 13 1 9 9 11
5 11 2 11 2 2
24 9 3 0 9 9 11 11 13 10 9 9 9 11 11 1 9 0 9 1 9 9 11 11 2
11 11 2 11 15 13 1 9 1 9 11 2
26 11 3 3 13 1 11 2 11 9 1 9 0 9 7 9 11 2 0 1 11 1 9 1 0 9 2
7 9 7 1 15 13 0 2
32 13 15 2 1 10 0 9 15 9 9 9 1 9 13 7 3 1 15 13 1 10 9 2 1 11 7 1 9 2 13 11 2
14 9 11 11 2 11 3 13 3 1 9 1 10 9 2
23 13 2 14 1 0 9 2 3 0 2 15 13 10 9 13 2 13 2 16 1 15 13 2
21 9 13 3 0 2 16 4 9 13 2 16 15 15 13 2 13 15 11 2 11 2
27 0 9 13 1 15 1 9 1 0 9 9 9 0 9 2 15 13 7 0 1 9 9 9 1 9 9 2
7 3 15 13 9 1 9 2
15 9 13 0 2 16 15 15 9 13 2 13 11 2 11 2
29 9 0 9 3 13 0 9 9 1 9 9 2 15 1 11 13 13 1 9 1 9 9 2 15 15 13 0 9 2
27 16 9 3 13 1 0 9 9 1 9 7 0 9 13 2 13 15 1 15 3 0 2 13 11 2 11 2
15 1 15 13 3 0 1 10 9 13 3 3 9 0 9 2
37 11 2 11 15 13 2 16 13 3 0 2 16 4 4 1 9 2 15 13 1 9 7 1 9 2 1 9 10 9 13 0 9 16 1 0 9 2
21 9 11 3 13 2 16 9 13 3 3 0 9 2 7 10 9 1 9 13 0 2
9 1 9 11 2 11 15 7 13 2
20 9 1 9 4 13 13 3 0 9 2 16 13 1 10 9 2 13 15 11 2
5 9 11 13 0 9
2 11 2
34 9 9 1 9 0 9 9 7 0 11 2 11 2 1 0 11 1 11 13 16 0 9 2 13 1 9 9 0 9 9 9 11 11 2
36 9 15 3 13 2 7 13 15 15 2 15 4 3 1 9 13 1 9 2 7 3 3 13 13 13 1 0 9 2 1 0 9 2 13 11 2
21 13 3 1 9 0 9 7 9 2 15 1 9 3 13 9 9 1 11 1 11 2
15 9 4 13 1 9 0 11 2 3 13 10 9 3 0 2
15 0 9 15 13 1 12 9 9 1 12 9 9 1 11 2
14 0 9 4 9 13 1 9 9 0 9 12 9 3 2
6 11 15 13 9 0 9
7 11 11 2 9 11 7 11
19 0 9 0 0 9 9 0 9 13 3 0 9 0 9 0 9 10 9 2
16 3 13 0 1 0 9 2 3 15 13 0 9 9 0 9 2
8 13 3 1 0 9 0 9 2
30 3 15 1 11 13 0 9 0 9 2 0 9 0 9 7 0 9 2 3 0 9 9 2 0 9 7 9 0 9 2
23 7 3 1 9 0 7 0 9 2 3 3 13 11 2 13 7 1 0 9 1 0 9 2
23 10 0 9 13 10 9 3 1 3 0 9 0 7 0 9 0 9 1 0 9 0 9 2
28 1 9 13 13 10 9 2 0 7 0 9 0 9 13 1 9 9 0 9 7 9 15 0 0 9 7 9 2
16 1 10 9 3 0 9 13 3 0 9 0 0 9 1 9 2
27 1 12 0 9 0 9 13 0 9 2 14 1 12 5 2 2 16 0 9 13 1 0 9 1 12 5 2
16 9 9 0 0 9 2 9 2 1 15 0 9 13 0 9 2
29 1 0 9 15 3 13 0 9 2 15 3 1 9 12 13 9 0 9 1 12 5 7 1 9 12 1 12 5 2
18 1 11 1 9 12 13 1 9 1 12 5 7 1 11 1 12 5 2
12 7 1 0 7 0 9 0 9 13 0 9 2
9 0 9 13 1 9 12 3 11 2
13 1 9 0 9 12 13 7 1 11 1 0 9 2
8 0 9 9 13 3 0 9 2
21 1 9 9 1 12 9 13 11 1 12 9 1 12 1 11 7 12 9 1 11 2
13 0 9 13 0 7 1 9 9 9 9 1 9 2
21 9 0 9 13 1 9 12 0 2 0 2 3 1 0 9 9 12 9 2 9 2
6 1 0 9 13 0 2
15 3 1 11 12 9 2 9 7 1 11 12 9 2 9 2
17 9 0 9 0 9 1 3 0 9 13 0 3 3 1 0 9 2
9 1 9 12 13 12 9 2 9 2
25 0 9 9 13 0 9 9 2 1 15 0 9 1 0 9 7 3 1 9 0 7 0 0 9 2
15 1 0 9 1 9 0 9 9 9 9 13 3 0 9 2
12 7 7 3 13 0 0 9 0 9 0 9 2
21 9 9 1 9 12 1 11 7 1 11 3 13 9 12 5 2 3 2 12 5 2
22 1 11 15 13 1 12 5 2 16 1 0 9 15 3 13 1 3 0 9 12 5 2
10 0 9 13 3 0 9 9 9 9 2
11 1 9 9 12 1 15 13 3 9 0 2
18 9 1 9 13 12 9 2 7 15 13 14 12 5 0 0 0 9 2
13 1 11 15 13 12 9 2 3 2 12 5 9 2
23 3 15 13 11 1 12 9 7 12 5 9 7 0 9 1 12 9 7 0 12 5 9 2
25 7 1 0 9 0 15 9 9 9 7 9 9 0 7 0 1 9 0 9 11 3 13 10 9 2
29 3 1 0 9 0 9 2 0 9 0 9 2 1 3 0 9 0 9 2 1 0 9 0 9 7 0 9 9 2
14 3 3 13 0 9 9 7 0 9 7 3 0 9 2
8 15 13 0 9 9 0 9 2
25 13 0 2 16 9 11 15 1 0 9 13 10 0 0 9 7 13 15 3 3 9 0 0 9 2
7 11 15 13 9 0 9 2
2 9 9
2 11 2
17 1 0 9 1 11 15 1 9 13 9 1 9 9 15 9 9 2
13 9 0 9 1 11 15 3 3 13 9 0 9 2
24 9 9 11 11 11 13 2 16 0 0 9 4 1 9 1 0 9 3 3 13 3 0 9 2
12 9 0 15 1 0 9 9 7 4 15 13 2
3 0 9 9
7 11 2 11 2 11 2 2
25 9 9 4 13 0 13 14 1 0 9 9 2 16 15 13 9 0 9 1 9 12 0 9 9 2
9 9 11 15 13 9 1 0 9 2
9 9 10 9 4 3 13 1 9 2
22 9 9 13 1 9 0 9 11 11 9 1 9 1 3 12 9 0 2 16 13 3 2
6 9 13 14 12 9 2
24 9 0 9 13 3 9 0 0 9 2 3 1 0 11 2 11 2 11 2 11 7 0 2 2
17 9 9 13 1 11 11 1 10 9 2 10 9 13 0 13 9 2
8 12 9 9 9 13 1 9 2
11 0 9 13 7 9 1 9 1 0 9 2
15 0 9 4 11 13 10 9 1 11 7 1 0 12 9 2
21 1 9 9 2 3 13 11 2 11 2 15 3 4 13 9 2 16 4 9 13 2
21 9 9 13 2 16 10 9 1 9 12 13 12 9 2 15 4 13 3 0 9 2
8 1 9 13 9 12 9 9 2
15 9 9 11 11 13 9 16 9 1 9 9 7 9 9 2
28 9 15 1 15 13 3 13 0 9 2 16 4 13 1 0 9 13 0 7 0 9 2 1 15 13 7 9 2
35 9 9 13 1 0 9 1 9 9 1 9 12 1 0 13 0 9 2 13 11 0 9 11 11 2 9 9 1 9 13 12 9 9 2 2
17 13 7 2 16 7 9 9 13 1 9 1 9 12 1 9 9 2
12 13 15 3 1 9 0 9 7 9 9 9 2
26 1 0 9 4 0 9 13 1 9 9 1 12 9 2 1 9 2 7 7 1 9 0 7 0 9 2
13 0 9 13 1 9 0 9 1 0 9 7 9 2
22 1 9 9 9 13 2 16 9 15 1 9 9 1 9 12 13 13 9 1 0 9 2
4 11 13 0 9
3 1 0 9
5 11 2 11 2 2
21 9 9 0 9 0 9 15 9 1 9 0 9 11 11 11 13 1 0 9 11 2
21 15 9 1 9 0 13 3 14 3 9 9 1 0 9 7 0 9 1 15 0 2
11 11 13 3 9 9 11 11 1 3 0 2
29 9 9 7 14 13 9 9 0 9 2 15 4 1 9 12 3 13 9 2 7 3 0 9 0 9 11 1 9 2
34 3 13 9 11 11 11 2 9 9 11 1 0 9 1 11 13 9 1 12 2 9 2 7 10 9 9 13 3 3 15 1 0 9 2
9 11 2 11 2 9 9 4 13 3
3 1 0 9
2 11 2
24 1 0 9 7 1 0 9 1 0 9 13 9 0 0 9 11 11 0 9 9 1 0 9 2
7 9 9 13 12 2 9 2
22 11 15 13 2 16 0 9 13 1 9 13 0 9 2 7 3 15 0 2 9 9 2
35 1 9 2 10 0 9 15 13 13 2 11 13 2 16 3 0 9 13 3 13 9 2 15 3 13 2 7 13 1 10 9 10 9 13 2
30 1 11 4 13 4 1 9 13 0 9 1 9 2 16 1 10 9 4 13 15 9 13 2 7 9 9 13 1 9 2
8 11 7 11 13 1 9 9 9
3 1 0 9
2 11 2
28 3 0 9 7 0 9 9 3 13 0 0 9 2 16 4 15 13 1 0 9 7 13 13 0 0 9 9 2
16 1 9 1 9 9 9 7 9 11 15 13 9 11 11 11 2
28 9 9 7 11 1 9 12 9 1 12 2 9 2 15 4 1 9 3 13 2 13 11 1 0 9 10 9 2
34 1 0 9 4 0 7 0 9 9 1 11 13 0 9 1 15 9 2 1 15 15 13 1 0 7 0 2 1 11 7 11 2 11 2
30 11 13 1 9 1 9 0 9 2 9 0 9 7 0 9 0 0 9 1 0 9 1 9 0 9 1 9 0 9 2
4 9 9 7 9
2 9 2
2 11 11
28 13 15 15 15 0 1 15 2 16 4 15 13 0 9 11 1 9 13 1 9 2 16 4 3 13 1 0 9
26 16 4 15 11 13 3 13 9 1 9 1 0 9 14 3 2 16 4 13 9 2 15 14 13 15 2
18 3 3 13 1 15 2 13 9 1 9 9 2 16 4 13 9 0 2
28 13 3 0 2 16 4 9 13 0 9 1 9 9 2 13 7 3 3 0 2 16 13 0 9 1 0 9 2
29 15 3 15 7 9 15 0 9 13 1 0 9 1 9 9 9 7 10 0 9 2 15 3 9 4 13 13 9 2
16 3 9 2 13 2 14 4 13 9 3 0 2 3 7 0 2
5 0 9 7 0 9
6 11 11 2 9 0 9
26 9 0 9 7 1 15 1 0 9 0 9 0 0 9 13 3 1 0 9 3 3 1 9 10 9 2
31 13 15 3 1 10 9 2 16 15 9 0 9 13 3 1 10 15 13 2 3 1 10 9 2 16 3 13 9 15 13 2
41 3 3 15 13 2 16 9 0 9 13 3 0 2 7 7 7 0 2 0 9 1 9 1 0 9 16 3 1 9 7 16 1 15 7 13 13 3 3 7 3 2
32 14 3 13 0 9 1 9 9 9 0 9 9 0 9 2 14 3 15 1 11 9 9 13 9 0 9 9 3 1 0 9 2
9 14 15 13 7 0 7 3 0 2
38 1 12 10 9 4 15 7 13 10 9 13 1 9 0 7 0 7 3 0 2 0 9 2 1 9 2 3 3 13 2 1 9 0 9 7 0 9 2
48 3 3 2 13 2 14 1 9 7 9 9 2 7 14 1 9 9 7 9 2 13 1 0 9 2 1 0 0 9 2 7 15 13 14 3 15 2 1 15 13 9 10 7 15 9 3 13 2
52 1 10 9 1 0 9 9 7 9 4 7 13 2 1 10 9 2 1 0 9 2 9 9 2 3 13 10 9 3 0 7 3 13 4 3 13 14 1 0 9 2 13 0 9 9 0 9 2 1 15 13 2
12 13 9 9 9 9 9 2 15 1 15 13 2
6 13 9 10 0 9 2
26 15 13 3 9 1 9 1 15 1 0 9 0 7 3 0 2 7 1 0 9 15 13 13 3 3 2
54 3 15 13 1 15 2 16 9 0 9 13 9 9 3 15 15 2 7 9 14 10 1 15 2 16 13 3 9 9 10 0 16 15 15 7 16 13 3 9 10 7 15 9 9 2 10 0 9 3 1 9 0 9 2
12 13 13 1 15 2 16 10 9 13 0 9 2
79 9 2 16 4 1 9 1 0 9 9 0 9 0 9 3 13 7 9 0 9 0 9 3 3 13 2 13 2 3 0 16 9 1 9 9 0 1 15 2 2 0 16 9 1 9 9 2 2 3 0 2 16 13 9 1 9 9 0 1 15 7 16 13 0 9 1 9 15 1 15 13 1 15 0 0 2 0 9 2
23 10 12 9 9 3 13 2 16 13 1 9 0 2 7 16 13 1 0 9 10 0 9 2
42 13 3 13 2 16 0 9 9 1 9 0 7 0 7 0 0 9 0 9 7 0 9 13 10 0 9 1 9 9 9 7 0 9 2 15 4 16 9 3 13 13 2
35 0 9 2 0 1 0 9 0 9 7 1 0 0 9 2 13 9 1 10 9 0 2 13 9 9 0 2 7 16 15 13 10 0 9 2
30 3 3 13 9 10 0 9 2 10 2 3 3 0 9 9 2 9 7 0 9 13 10 9 13 2 13 15 14 13 2
20 3 0 9 2 7 3 0 9 2 13 9 2 3 0 1 0 9 1 9 2
55 3 9 2 0 0 9 1 9 2 9 7 9 2 15 13 0 9 1 9 2 7 13 4 13 2 16 1 10 9 13 0 9 7 10 0 9 3 13 2 7 15 15 13 1 9 9 7 10 0 9 7 13 0 9 2
27 10 0 9 1 0 9 2 15 4 3 3 3 13 7 13 2 13 7 13 4 1 0 9 13 9 9 2
26 9 0 2 0 0 9 13 14 0 9 7 9 15 0 9 2 7 13 7 9 0 9 1 0 9 2
44 0 13 2 16 1 0 9 0 0 9 13 10 0 9 9 15 15 2 0 9 7 9 0 9 9 0 9 2 7 16 10 0 0 9 13 2 3 2 7 0 2 7 0 2
60 9 1 9 7 9 9 13 9 0 9 1 9 0 9 0 0 9 2 7 13 9 1 15 2 16 13 9 9 15 0 0 7 0 9 0 7 0 9 7 16 15 15 13 13 9 0 2 9 9 2 9 3 0 2 3 9 0 2 0 2
30 13 10 9 4 15 13 1 0 9 2 15 4 3 3 13 7 15 2 3 15 1 15 2 3 13 3 13 1 9 2
28 9 2 3 3 0 9 2 2 0 3 1 10 0 0 9 2 13 3 3 0 16 0 0 9 10 9 0 2
18 3 10 9 13 13 9 10 9 7 1 9 0 9 7 9 0 9 2
6 13 9 1 9 9 2
3 11 11 2
8 9 13 9 11 1 0 0 9
29 12 1 3 0 9 1 9 1 0 0 9 13 9 7 9 9 1 9 0 9 2 0 1 0 9 1 0 9 2
37 3 1 9 0 9 2 7 14 1 15 2 3 13 2 16 9 13 1 9 0 9 9 2 7 3 3 7 15 2 16 13 9 0 9 3 0 2
9 9 2 1 15 13 2 13 0 2
32 0 9 2 0 9 2 7 3 0 9 2 15 10 9 3 13 7 15 13 10 9 2 13 0 7 10 9 7 9 3 0 2
14 9 13 3 0 9 2 0 15 9 1 0 9 9 2
37 9 13 7 15 2 10 9 13 4 1 9 0 9 7 1 9 3 0 9 13 2 7 3 15 2 3 13 2 16 4 10 9 13 10 0 9 2
13 9 2 10 9 1 9 9 13 2 13 9 0 2
36 16 9 13 15 15 13 2 13 2 14 1 9 9 2 15 13 4 1 9 13 2 13 3 13 0 9 1 9 9 2 15 13 9 10 9 2
9 9 13 3 0 2 13 9 9 2
15 9 9 0 9 1 9 9 0 0 0 9 13 3 0 2
16 13 1 15 3 1 12 2 9 9 0 9 1 9 11 11 2
11 13 1 15 2 13 9 1 9 1 9 2
20 10 9 2 15 15 3 13 9 13 0 9 2 13 1 10 9 0 3 13 2
17 10 9 13 3 0 9 2 7 4 1 3 0 9 13 1 9 2
30 1 9 12 4 0 9 13 9 1 9 9 2 15 3 13 0 9 9 9 9 0 0 9 0 0 9 2 3 9 2
14 9 13 10 9 13 1 9 9 12 10 9 1 9 2
10 3 10 9 13 9 1 9 1 9 2
11 0 9 13 9 9 12 9 9 0 3 2
33 16 10 9 13 9 9 3 2 16 15 13 13 1 9 2 13 13 10 0 9 9 0 9 2 15 3 13 13 9 1 0 9 2
8 0 9 9 9 13 3 13 2
21 0 11 11 13 0 9 10 0 9 1 0 9 10 9 2 10 9 13 3 0 2
21 0 11 11 13 0 9 10 0 9 1 0 9 10 9 2 10 9 13 3 0 2
13 3 13 1 9 2 16 3 13 9 1 9 9 2
22 1 15 2 16 9 13 1 9 2 13 9 9 9 9 1 12 9 1 12 0 9 2
10 0 9 13 3 0 2 0 12 9 2
26 9 7 13 10 9 7 13 9 1 9 9 9 2 0 9 9 1 12 9 9 13 3 0 12 9 2
45 1 15 2 16 4 13 9 9 9 3 3 2 13 0 7 15 2 16 9 1 9 0 9 3 13 2 16 1 9 12 4 13 0 9 9 2 12 9 9 2 1 0 12 9 2
37 1 9 4 10 0 9 13 12 9 2 1 0 0 9 13 9 1 0 9 9 2 16 13 9 2 16 13 15 1 15 3 0 16 1 0 9 2
24 7 1 0 9 13 9 1 0 9 9 9 2 13 3 1 0 9 9 9 1 0 9 9 2
17 10 9 13 13 3 1 9 0 9 2 3 1 9 0 0 9 2
6 7 7 15 13 9 2
23 13 15 3 1 0 9 9 1 9 1 9 9 0 2 16 13 15 3 1 9 1 11 2
3 9 1 11
2 11 2
13 0 9 9 11 13 9 11 0 9 3 1 9 2
20 1 9 9 11 2 11 1 9 0 9 15 4 3 1 0 9 13 3 9 2
12 9 9 13 1 9 1 12 1 12 12 9 2
38 3 2 16 9 0 9 11 13 9 1 9 2 9 11 3 13 9 1 12 9 2 15 13 13 0 9 2 14 12 9 2 9 2 0 1 0 9 2
15 9 13 1 15 2 16 9 4 13 1 11 1 12 9 2
9 9 13 0 9 12 9 1 9 2
20 1 9 0 0 9 13 9 9 14 12 9 2 1 0 0 9 14 12 9 2
3 0 9 11
1 9
2 11 11
20 16 16 13 1 9 9 2 13 1 9 1 9 0 9 0 0 9 10 9 2
4 3 15 0 2
26 1 0 9 2 13 15 13 1 0 9 9 0 9 2 15 13 11 3 1 10 9 13 9 0 9 2
37 0 7 3 3 15 0 9 9 11 15 13 3 13 2 16 4 15 13 13 1 9 10 9 0 9 2 7 0 9 7 9 15 13 13 1 9 2
21 14 3 3 1 9 13 1 0 9 1 11 2 3 13 0 9 11 2 13 9 2
17 0 9 3 13 13 14 0 9 0 9 2 7 3 9 10 9 2
24 13 0 2 16 1 9 0 9 13 0 13 1 9 7 13 9 0 1 0 9 9 16 3 2
21 0 9 15 3 13 15 2 16 16 15 13 1 9 2 4 15 0 9 3 13 2
18 1 0 0 0 9 4 3 3 3 1 9 13 13 1 0 0 9 2
35 7 13 1 9 1 0 9 0 9 0 9 2 15 4 15 1 3 0 9 13 13 0 9 2 13 3 0 9 2 15 13 1 9 9 2
25 9 13 9 0 9 1 9 9 7 9 7 13 2 16 15 15 3 13 13 3 2 15 3 13 2
18 1 1 15 2 16 15 11 1 0 9 0 9 1 9 7 13 13 2
19 1 9 9 2 15 3 13 7 9 9 1 0 9 2 0 9 13 13 2
17 7 1 0 9 15 13 13 2 16 1 10 9 13 7 9 9 2
10 15 3 13 0 9 1 9 0 9 2
5 13 3 1 9 2
23 13 4 3 1 9 2 16 4 15 9 10 9 13 15 9 0 9 11 2 1 9 11 2
18 1 9 9 1 3 0 9 7 0 9 13 0 2 7 0 0 9 2
38 13 2 16 0 0 9 3 13 2 7 13 2 4 13 2 9 11 15 3 13 1 9 2 16 10 9 13 15 0 1 15 2 15 13 9 1 9 2
15 1 0 15 0 9 13 9 1 9 0 9 0 0 9 2
6 15 3 2 15 3 2
23 9 11 11 11 1 9 1 0 9 11 1 11 1 9 13 0 9 1 9 11 2 9 11
2 9 11
1 3
10 9 11 1 11 13 0 9 1 9 2
40 13 15 3 0 9 9 11 2 11 2 15 3 13 2 16 13 1 10 0 9 2 7 13 2 16 0 9 3 13 1 0 9 11 2 15 4 13 9 9 2
30 0 9 11 2 11 13 9 2 15 13 1 9 9 2 15 15 13 13 1 9 1 0 9 3 1 0 9 7 9 2
8 13 1 15 3 9 0 11 2
30 0 0 9 1 11 1 9 0 9 11 2 11 7 9 9 11 2 11 15 1 12 9 13 1 12 0 7 12 0 2
5 13 15 0 9 2
11 0 9 13 1 9 12 1 0 9 9 2
9 11 2 11 13 1 9 12 9 2
21 1 9 12 15 3 13 1 9 1 9 11 2 11 2 15 13 9 9 1 11 2
27 9 9 11 11 2 11 13 1 9 1 9 1 11 2 16 4 3 1 0 0 9 13 1 9 0 9 2
16 1 9 9 11 13 1 12 0 9 12 1 0 9 11 11 2
4 0 9 13 3
8 1 0 9 3 13 0 0 9
4 11 2 11 2
22 9 1 0 2 0 9 2 3 13 14 12 0 9 1 0 11 2 15 3 3 13 2
26 1 9 0 9 1 9 1 9 1 0 9 1 0 9 0 0 11 1 15 11 3 13 10 0 9 2
27 3 7 9 2 15 13 1 0 9 1 9 0 9 11 11 2 15 1 0 9 0 9 1 10 9 13 2
26 3 0 9 2 15 13 9 13 1 0 9 2 3 9 11 15 3 13 3 10 9 9 13 1 9 2
20 0 9 13 3 9 13 2 16 4 15 9 13 13 9 7 13 1 0 9 2
13 11 7 10 9 13 3 9 3 1 9 0 9 2
24 1 9 4 12 1 9 2 15 1 0 9 13 1 9 0 9 11 2 13 3 1 0 9 2
49 9 9 9 0 9 1 0 11 11 1 11 15 1 9 13 3 1 11 11 7 1 9 9 0 9 2 11 1 11 2 11 11 2 1 15 13 1 9 9 2 15 1 9 0 9 13 1 11 2
22 1 9 13 1 9 11 2 12 9 3 1 11 2 1 0 9 2 15 13 0 11 2
25 11 1 9 13 2 16 13 3 0 13 9 9 9 2 7 1 10 9 13 10 9 1 9 11 2
20 10 9 15 7 13 1 11 7 11 1 9 2 13 15 1 0 9 9 9 2
34 9 9 13 0 9 9 0 0 11 2 15 1 0 9 13 0 9 2 7 13 15 1 0 9 1 9 15 2 15 13 1 9 9 2
21 11 15 7 13 13 10 9 1 9 2 16 3 13 0 13 0 9 0 0 9 2
17 1 9 1 0 9 13 1 15 2 16 4 15 13 1 10 9 2
9 1 11 7 1 11 3 2 13 11
2 11 2
22 1 0 9 9 11 11 3 0 9 13 1 15 2 3 14 15 13 0 9 0 9 2
27 1 9 1 9 11 13 11 9 2 16 0 9 11 2 15 13 9 1 0 9 2 4 13 7 1 11 2
35 1 15 9 16 11 2 11 7 0 9 1 9 1 0 9 13 13 2 13 11 7 13 2 16 3 1 11 7 11 13 0 13 0 9 2
6 0 9 15 13 1 9
2 11 2
17 9 0 9 1 0 9 13 12 0 9 7 13 0 9 0 12 2
9 13 15 1 9 0 0 9 11 2
29 9 2 0 15 1 0 9 2 13 2 3 0 9 13 2 7 1 9 9 9 1 9 1 9 0 9 13 9 2
17 0 9 11 11 13 3 0 9 2 15 13 13 1 11 0 9 2
23 0 11 15 13 13 1 9 3 2 16 0 9 1 9 13 1 0 9 1 9 0 9 2
6 9 11 13 0 9 11
8 11 2 0 9 2 11 2 2
23 0 9 1 9 3 13 9 2 1 10 9 13 11 1 0 9 11 9 1 12 0 9 2
25 0 9 13 13 9 11 7 9 1 9 11 2 11 2 1 11 1 9 1 11 7 9 11 3 2
13 0 0 0 9 2 11 2 13 9 3 1 9 2
32 11 3 13 2 16 1 11 13 9 7 9 0 9 2 15 1 9 1 9 11 3 1 11 11 13 1 9 12 0 0 9 2
27 1 9 15 13 0 9 0 9 2 11 2 2 15 13 0 9 1 11 7 11 7 13 1 9 1 11 2
21 0 7 0 9 15 3 13 1 9 1 9 0 9 2 3 7 3 1 0 9 2
15 13 13 1 9 2 15 13 13 1 0 9 1 12 9 2
24 3 16 12 0 9 13 3 9 1 9 2 15 13 1 9 1 0 9 7 9 1 0 9 2
17 0 0 9 11 11 13 9 2 16 11 7 11 3 13 1 9 2
5 11 2 9 0 9
2 11 2
20 0 9 13 1 9 1 9 1 9 1 11 12 0 9 7 10 9 3 13 2
21 1 0 9 1 11 4 9 13 1 9 1 9 11 2 14 12 9 3 1 11 2
14 12 0 9 4 13 0 9 7 12 0 9 4 13 2
15 3 1 9 4 13 1 0 9 2 10 9 7 13 13 2
5 9 9 13 0 2
3 9 1 9
2 11 2
15 11 1 9 9 13 2 16 7 1 9 13 4 0 9 2
8 3 13 1 9 1 12 9 2
16 16 9 13 3 1 9 2 0 9 0 9 13 0 9 9 2
14 1 0 9 13 9 1 0 7 1 9 1 0 9 2
13 13 15 7 3 0 9 1 9 9 7 1 9 2
5 0 9 13 1 11
5 11 2 11 2 2
23 0 0 9 0 9 15 1 9 1 0 11 13 0 9 2 15 13 0 9 1 9 11 2
6 9 13 0 0 9 2
21 9 11 11 4 13 1 0 9 1 9 2 15 13 1 11 12 9 3 1 11 2
12 1 0 9 9 10 9 1 9 13 10 9 2
33 9 13 13 2 16 13 3 1 9 0 9 0 0 2 11 2 15 15 13 3 1 0 9 1 0 9 2 15 13 9 0 11 2
6 12 9 9 1 9 11
4 11 2 11 2
17 0 9 13 0 9 9 1 9 12 9 9 1 9 9 0 9 2
21 13 15 3 1 11 0 9 11 1 15 2 16 9 4 13 9 13 1 10 9 2
18 1 10 9 11 13 9 3 1 9 2 1 9 0 9 7 1 9 2
15 12 9 1 9 0 9 0 9 13 9 1 9 0 9 2
35 0 9 0 9 1 11 1 9 13 0 9 9 2 16 4 3 9 12 0 0 9 13 2 16 13 3 13 1 9 7 1 9 0 9 2
23 0 9 9 11 2 11 1 9 13 9 1 0 9 2 15 15 13 1 0 9 1 11 2
11 11 13 2 16 13 3 0 0 9 13 2
25 15 2 16 0 9 13 1 0 9 11 1 9 2 1 11 13 2 16 10 9 13 10 0 9 2
7 1 9 2 7 0 9 2
4 11 11 2 11
25 0 9 9 2 3 4 1 0 11 13 0 0 9 2 3 3 13 9 7 9 1 9 10 9 2
22 16 0 9 1 12 9 13 12 2 9 1 0 9 2 13 15 16 15 0 0 9 2
19 3 15 13 9 2 15 11 13 1 0 9 2 1 0 9 0 0 9 2
22 10 9 13 7 0 9 9 2 15 13 9 2 16 11 13 0 9 1 9 0 9 2
43 9 11 11 2 15 9 7 9 13 2 1 9 13 2 0 9 13 1 9 7 15 3 1 9 2 1 9 7 9 10 0 9 7 0 0 9 2 1 0 9 7 9 2
27 1 15 2 16 11 13 3 0 9 14 1 9 7 9 2 13 7 9 11 1 9 10 0 9 7 9 2
15 9 0 9 13 2 16 10 9 13 1 11 10 0 9 2
22 1 11 13 3 9 2 15 15 1 11 13 3 2 3 7 15 2 15 13 9 0 2
12 0 13 9 2 15 13 14 3 13 1 9 2
30 9 9 0 9 11 11 13 11 1 0 9 1 9 11 2 16 15 15 11 13 1 9 2 15 15 3 13 1 9 2
25 15 1 15 15 3 13 9 1 9 0 15 2 16 0 0 9 13 9 11 1 0 9 2 13 2
18 9 1 9 11 13 2 16 10 9 15 13 13 0 11 9 0 9 2
37 9 9 11 11 1 9 2 16 13 1 9 1 9 2 13 2 16 9 13 9 2 16 15 9 13 7 11 0 1 9 0 9 2 15 13 9 2
41 13 1 9 3 2 16 4 15 1 11 13 9 2 9 2 16 1 10 9 15 1 9 7 9 13 13 2 13 15 9 1 9 2 7 14 1 9 2 13 11 2
42 9 0 0 9 11 11 13 2 16 11 13 3 16 0 0 9 9 16 9 1 9 2 7 3 7 16 9 2 3 15 13 1 0 9 2 15 1 9 9 13 9 2
26 13 3 0 9 7 15 15 13 1 15 2 16 4 13 0 1 9 10 9 13 2 16 1 0 9 2
16 1 10 9 15 13 9 9 1 0 9 2 15 13 0 9 2
24 9 9 0 0 9 15 3 13 1 9 3 13 2 1 0 0 9 13 7 0 0 9 9 2
16 1 15 13 3 12 12 2 12 9 2 9 0 9 11 3 2
5 11 13 0 9 11
2 11 2
29 0 0 9 1 0 0 9 2 11 2 3 13 0 0 0 9 2 11 2 9 11 11 1 11 9 1 0 9 2
9 1 9 13 1 11 1 12 9 2
14 0 9 7 13 2 16 15 3 13 3 16 12 9 2
31 15 11 3 13 11 2 16 13 1 0 9 1 11 2 11 1 0 0 9 1 0 1 9 0 9 0 9 2 11 2 2
5 9 13 9 15 13
2 11 11
48 16 15 9 1 0 9 13 13 3 0 9 0 7 0 9 1 11 2 11 13 15 2 15 13 3 2 13 15 15 2 13 11 11 11 2 11 2 9 0 9 0 11 0 2 0 1 11 2
45 9 0 0 9 13 13 3 3 2 7 13 2 14 15 1 0 9 0 9 1 11 7 11 2 13 11 11 13 9 2 1 15 1 10 3 0 9 13 1 9 0 7 0 9 2
26 9 11 13 0 9 9 1 10 9 0 0 9 1 9 1 11 1 9 13 3 0 9 9 1 11 2
13 11 15 1 0 0 9 13 10 0 9 3 13 2
11 0 0 9 1 10 9 13 9 1 9 2
17 0 9 1 9 0 9 3 13 2 16 4 9 1 9 13 9 2
25 9 0 9 13 2 16 9 9 1 0 0 9 13 7 13 15 14 2 1 0 9 2 1 9 2
10 10 11 13 3 0 9 16 0 9 2
18 7 9 2 15 13 1 9 3 13 2 13 13 1 0 9 7 13 2
17 9 1 15 13 13 1 9 12 2 3 11 3 3 13 0 9 2
9 3 13 9 2 15 15 13 13 2
23 11 11 13 1 0 9 10 9 7 3 2 7 13 9 0 9 2 7 13 10 0 9 2
15 15 2 16 13 9 0 1 9 1 11 2 13 0 9 2
32 1 0 0 9 2 15 13 3 9 1 0 9 1 11 0 2 15 11 3 13 2 3 15 9 13 7 13 15 13 1 11 2
12 1 0 9 15 11 11 3 13 14 3 3 2
12 15 15 14 13 0 13 1 10 9 11 11 2
23 0 9 2 15 9 13 2 13 2 16 3 13 2 16 4 15 1 0 9 13 0 9 2
16 0 0 9 1 11 13 11 1 9 2 7 3 13 0 9 2
44 1 9 15 2 10 9 4 13 13 11 3 1 9 2 3 0 11 2 13 3 0 9 2 15 13 9 11 12 2 9 7 15 13 0 9 1 11 7 13 9 9 0 9 2
19 1 11 11 13 14 3 0 0 9 10 9 13 0 12 9 12 9 9 2
14 10 0 1 11 13 1 9 9 7 9 1 11 13 2
21 11 13 2 16 1 11 3 13 9 9 3 2 1 9 10 0 9 1 0 9 2
5 15 13 3 13 2
9 0 13 15 1 0 9 1 11 2
25 1 11 1 11 13 1 11 0 9 7 1 15 13 9 0 1 10 9 9 7 13 9 1 11 2
5 15 3 13 0 2
20 0 2 15 13 1 0 9 1 11 1 11 13 2 13 0 9 9 7 9 2
19 11 11 10 0 9 13 9 10 0 9 2 15 15 13 9 0 11 13 2
17 1 0 9 15 0 9 13 2 1 9 0 13 7 0 9 0 2
15 3 2 7 3 1 0 9 2 13 1 9 11 16 15 2
15 7 10 9 1 9 1 0 9 3 13 0 16 1 15 2
4 15 4 3 13
7 14 2 13 15 0 9 2
11 7 13 12 1 15 2 15 15 13 13 2
31 9 2 11 11 2 9 2 2 9 0 9 7 9 0 9 0 9 2 15 13 4 13 1 11 2 11 2 1 9 12 2
33 2 11 13 9 1 0 0 9 2 3 16 11 7 0 9 7 11 2 7 15 10 9 1 9 9 13 2 16 13 0 1 9 2
11 9 2 15 10 9 13 2 3 13 13 2
10 11 11 2 9 9 0 0 11 11 2
7 13 13 1 9 9 11 2
19 11 2 11 2 15 13 2 16 3 13 9 10 9 1 0 9 1 11 2
24 2 1 0 9 13 0 2 13 2 14 10 9 0 9 13 0 9 1 10 9 16 1 9 2
12 9 9 11 11 11 1 0 9 1 0 9 2
34 9 11 2 15 13 0 9 9 7 0 9 2 13 1 9 13 9 3 0 2 16 13 1 9 2 3 13 10 9 1 9 0 9 2
6 1 9 9 11 11 11
4 3 0 11 11
8 0 9 2 9 2 7 0 9
2 11 11
21 3 3 16 12 9 13 11 9 2 15 1 15 13 9 0 9 0 11 11 11 2
23 0 9 11 11 13 1 0 9 1 11 0 9 2 13 2 14 7 10 0 7 0 9 2
20 13 15 9 9 2 15 9 0 9 11 13 1 9 1 0 9 11 7 11 2
24 1 9 12 0 9 11 3 13 7 1 9 1 15 15 3 3 13 9 15 1 0 0 9 2
14 9 2 15 11 1 0 9 9 13 2 11 14 13 2
19 13 15 3 10 9 2 3 11 13 3 3 1 0 2 7 15 3 13 2
13 11 11 13 1 10 9 11 2 1 9 0 9 2
24 13 7 0 13 14 12 12 9 1 0 12 9 3 0 9 2 3 15 15 0 9 11 13 2
23 0 9 9 11 11 13 3 15 0 9 9 2 7 1 9 2 16 15 4 13 0 9 2
12 11 11 3 13 2 16 1 0 9 13 15 2
38 0 9 15 3 13 2 16 4 11 13 9 11 3 13 2 16 4 15 13 13 0 9 7 9 2 15 9 13 1 9 9 2 7 13 9 9 0 2
16 9 15 13 0 2 7 9 1 11 13 1 0 9 3 0 2
12 13 15 15 1 9 7 3 7 15 3 13 2
30 0 9 1 0 9 2 16 13 9 9 11 7 9 11 11 15 13 2 16 13 0 13 1 9 7 9 13 0 9 2
33 1 0 9 3 0 11 13 9 2 16 13 2 16 15 1 11 3 3 13 9 1 9 0 9 7 13 1 0 9 1 0 9 2
21 7 1 11 15 13 9 2 16 4 15 9 13 16 14 13 2 3 3 3 13 2
23 0 9 0 1 0 9 13 2 16 4 13 0 9 13 7 0 9 4 3 3 15 13 2
19 9 0 9 1 9 7 0 0 9 13 2 16 13 0 13 1 11 13 2
14 15 15 7 13 3 1 11 0 0 2 0 0 9 2
29 13 3 1 9 3 9 2 7 10 9 7 9 11 11 11 4 13 1 3 0 9 16 11 2 14 1 0 9 2
13 0 11 14 13 13 9 9 1 0 9 1 11 2
26 4 7 3 3 13 3 10 9 7 3 0 9 13 12 1 0 9 2 15 4 13 10 0 9 13 2
19 0 9 3 0 9 3 13 2 7 13 3 0 2 0 2 7 0 9 2
11 13 3 1 9 7 9 13 1 0 9 2
7 15 7 13 0 0 9 2
24 9 2 16 4 11 11 13 13 13 7 16 13 1 10 9 0 9 2 13 13 1 0 9 2
37 9 1 0 9 13 3 3 15 0 2 15 11 7 0 0 9 13 2 16 15 13 13 0 0 9 7 13 15 13 0 9 9 13 1 0 9 2
28 14 2 3 2 16 7 11 15 3 13 3 3 0 9 11 13 15 9 1 9 2 16 15 13 9 1 11 2
20 0 0 9 9 7 0 9 9 13 9 2 16 4 15 1 11 13 15 13 2
28 1 9 2 3 0 13 9 11 11 16 0 9 0 9 7 0 9 1 9 1 9 2 7 13 9 1 9 2
36 1 9 10 9 2 15 13 3 15 0 2 3 0 7 3 0 2 4 1 11 13 13 9 7 9 2 15 9 15 1 10 9 15 13 13 2
5 0 9 1 0 9
5 11 11 2 11 11
33 0 9 11 11 15 1 9 13 1 0 9 2 3 0 1 11 0 9 2 2 15 15 1 9 10 9 13 13 9 9 0 11 2
21 10 0 9 13 14 13 0 0 9 2 11 2 2 16 4 3 13 0 9 9 2
16 0 9 13 11 11 2 0 9 9 11 7 0 9 9 11 2
16 0 10 9 13 11 11 2 11 2 9 0 9 1 0 11 2
17 1 11 13 3 1 10 9 3 0 9 7 1 10 9 14 3 2
27 11 1 10 9 13 1 9 0 9 2 16 4 15 13 1 9 13 0 11 2 9 11 7 0 9 9 2
23 1 9 13 9 3 1 9 11 2 11 9 1 0 9 11 2 15 13 0 9 0 9 2
21 11 3 9 13 1 0 9 1 0 9 2 15 9 1 11 7 11 3 3 13 2
13 1 9 9 3 13 0 9 1 9 1 0 11 2
53 11 2 11 15 13 3 2 9 1 11 7 11 2 11 11 13 9 0 9 0 9 7 9 2 0 0 0 0 9 2 2 9 0 9 1 11 7 11 7 3 0 9 2 15 13 1 9 9 0 9 2 2 2
23 0 9 9 1 11 13 2 16 11 11 13 0 9 2 16 4 13 13 9 1 0 9 2
15 9 7 9 0 2 0 9 13 3 0 1 0 9 11 2
10 9 0 11 13 9 2 9 7 9 2
9 3 15 13 1 9 0 0 9 2
10 9 4 13 1 9 0 9 11 11 2
7 9 9 9 10 9 13 2
27 13 15 2 16 9 2 16 9 9 11 13 9 2 15 15 13 7 3 13 1 9 1 11 2 11 13 2
21 1 9 1 9 11 11 9 13 2 16 10 9 13 0 9 1 11 3 0 9 2
21 11 2 11 3 13 2 13 9 13 2 16 10 9 13 3 16 0 9 1 9 2
15 7 15 7 15 3 13 2 7 13 2 16 11 13 9 2
18 3 16 13 0 9 11 2 16 4 15 10 0 0 9 13 12 9 2
7 0 9 0 9 3 13 2
36 7 16 9 13 2 16 0 9 2 9 0 9 11 7 11 2 13 0 9 0 9 2 10 0 9 1 11 2 11 11 7 11 11 3 13 2
16 9 1 11 7 11 13 0 7 0 9 1 11 15 3 13 2
16 11 7 0 9 11 13 1 9 9 13 10 1 9 0 9 2
14 11 15 3 13 2 16 11 3 3 13 9 1 9 2
28 3 1 9 1 9 2 1 15 13 16 9 13 9 9 2 7 1 0 0 9 2 15 3 3 13 0 9 2
13 0 9 15 13 2 16 15 11 3 13 13 9 2
14 10 9 13 2 16 15 15 13 3 1 9 9 9 2
3 13 15 2
18 3 1 9 11 11 1 0 9 1 9 13 1 12 9 1 0 9 2
12 9 2 15 15 13 3 12 0 2 0 13 2
16 13 0 2 16 9 13 9 7 9 7 0 9 15 3 13 2
16 16 0 15 7 13 2 16 1 0 11 13 0 9 1 9 2
9 9 4 3 13 1 9 10 9 2
5 9 13 2 9 13
2 11 2
19 9 12 0 0 9 11 7 11 1 9 13 2 9 10 9 15 7 13 2
8 13 15 1 0 9 12 9 2
29 0 9 11 1 9 1 0 9 13 1 12 9 1 12 9 2 16 1 0 9 9 13 10 0 9 1 12 9 2
11 0 9 7 13 1 12 9 1 12 9 2
21 9 11 15 1 9 13 1 12 9 1 12 9 1 9 9 1 0 11 7 11 2
16 0 9 13 1 12 9 1 12 9 1 9 9 1 0 9 2
23 9 11 1 0 9 3 13 1 12 9 1 12 9 7 9 3 13 12 2 9 0 9 2
16 1 9 15 7 13 12 9 11 2 15 13 9 1 12 9 2
27 9 9 11 15 1 9 13 1 12 9 1 12 9 2 16 1 9 9 13 10 0 9 9 1 12 9 2
21 9 1 0 9 7 3 13 3 0 9 1 15 2 3 1 12 9 1 12 9 2
5 9 11 1 12 9
2 11 11
9 16 4 15 9 9 13 1 9 2
11 1 9 1 0 9 13 12 9 9 11 2
6 3 16 1 12 9 2
22 3 15 7 13 0 9 9 7 9 1 9 2 7 9 9 11 11 7 9 11 11 2
10 12 1 0 9 0 9 9 11 13 2
19 1 12 2 9 1 12 2 9 13 0 9 1 10 0 9 1 12 9 2
19 3 15 3 1 11 13 2 16 9 11 13 0 0 9 1 9 1 11 2
17 14 10 9 1 9 0 9 15 9 10 9 0 11 13 1 9 2
23 1 0 9 1 0 9 13 3 0 7 9 11 15 10 9 13 13 1 11 0 0 9 2
28 1 10 9 7 1 11 3 13 2 16 4 15 11 9 13 1 10 9 7 4 13 11 2 7 2 0 9 2
24 15 15 15 2 3 1 9 9 11 2 1 15 15 1 11 3 13 3 16 1 11 2 13 2
20 1 0 9 12 2 9 1 0 9 3 13 9 2 15 13 1 9 0 9 2
11 0 9 9 9 11 4 13 16 0 9 2
11 0 9 13 7 0 9 15 13 1 9 2
21 1 10 9 15 13 0 9 9 11 11 2 3 12 1 0 9 12 2 0 9 2
22 9 12 15 11 1 11 13 1 9 1 0 0 9 2 16 13 3 13 1 0 9 2
14 10 9 1 10 0 9 1 0 9 7 13 1 9 2
20 0 9 13 9 0 9 9 1 11 2 15 1 9 12 13 0 9 1 11 2
16 13 3 1 11 1 9 13 11 1 9 7 13 1 0 9 2
7 9 1 15 15 3 13 2
19 1 9 2 12 13 1 0 9 11 7 1 12 9 3 1 0 9 11 2
22 1 11 7 3 1 10 9 1 11 13 1 11 7 13 15 3 1 0 0 9 9 2
13 1 9 1 11 3 13 9 2 16 15 9 13 2
8 4 7 3 3 13 15 13 2
14 3 2 16 15 13 2 16 1 0 9 13 0 9 2
23 1 9 15 3 3 13 7 9 9 2 15 12 9 9 13 12 2 9 9 0 9 11 2
12 7 10 9 15 7 13 1 9 0 1 0 2
12 0 7 0 9 15 3 13 1 9 7 9 2
29 13 13 9 2 16 9 2 15 15 3 13 12 9 2 13 9 2 13 9 9 7 12 2 9 13 11 9 9 2
26 1 9 9 13 3 3 3 15 9 9 1 15 2 16 11 1 9 12 13 1 11 9 7 0 9 2
14 16 15 9 1 11 13 1 11 7 10 9 3 3 2
8 1 0 9 13 9 0 9 2
32 16 15 11 13 1 0 9 9 1 9 9 7 9 1 11 13 1 0 11 1 0 0 9 2 13 15 13 1 9 0 9 2
16 0 9 1 15 13 11 0 9 7 1 11 1 10 9 9 2
14 3 15 0 13 1 9 2 16 15 13 9 0 9 2
22 0 9 1 15 2 16 0 9 12 13 1 9 0 9 3 2 3 13 2 1 9 2
7 9 2 16 9 13 14 12
8 11 11 2 9 0 9 0 9
56 1 9 9 0 9 2 2 2 13 11 2 11 2 11 12 2 12 2 2 9 1 15 2 16 3 4 1 9 0 9 13 0 9 2 1 15 4 13 13 13 9 2 9 2 9 2 9 7 0 0 9 1 0 10 9 2
30 13 15 16 4 13 1 15 0 2 7 1 9 3 10 9 13 1 9 10 2 7 1 0 9 2 7 15 0 9 2
20 9 9 2 15 13 9 9 1 9 2 12 2 4 13 1 9 1 10 9 2
10 3 13 0 9 13 7 13 3 3 2
26 1 12 2 9 13 10 9 11 11 2 1 12 2 9 9 11 11 2 1 12 2 9 9 11 11 2
23 15 1 10 12 9 15 0 13 2 7 15 3 2 16 15 10 9 13 1 15 0 13 2
15 1 0 1 10 9 13 12 2 12 9 2 15 0 9 2
7 7 10 9 2 10 9 2
16 0 9 13 10 9 3 3 2 16 0 9 13 1 9 9 2
17 9 1 12 2 9 13 3 3 10 9 0 1 0 9 0 9 2
11 9 9 10 9 15 13 3 13 3 3 2
16 9 11 11 15 3 15 13 2 16 0 9 13 3 12 9 2
16 13 9 2 16 15 13 14 12 2 3 4 0 9 13 3 2
36 7 13 13 2 16 7 15 12 13 1 15 9 0 9 2 16 0 9 13 12 7 12 9 7 0 15 3 13 2 16 4 9 13 4 13 2
16 13 0 2 16 4 1 0 9 13 9 0 16 1 0 9 2
13 13 0 3 3 13 2 10 9 4 1 9 13 2
16 13 9 2 3 15 12 1 15 13 1 9 1 12 0 9 2
35 11 11 1 10 9 1 0 9 13 2 16 13 9 9 1 10 0 9 7 3 2 16 15 15 13 2 7 3 2 16 13 10 9 0 2
23 11 11 1 15 13 9 1 15 2 16 1 9 9 7 9 15 13 9 9 16 1 9 2
22 3 9 9 13 3 0 0 9 7 9 13 3 0 9 7 1 15 15 0 9 13 2
33 3 12 9 2 1 0 9 1 9 9 9 9 13 3 0 9 2 1 15 9 11 11 13 1 15 2 16 4 9 13 3 0 2
12 13 4 3 12 9 9 0 9 1 12 9 2
17 7 3 15 14 4 13 1 9 2 15 4 13 3 3 12 9 2
2 0 9
14 1 0 9 9 3 13 3 3 13 9 0 1 9 2
15 3 13 3 13 12 9 9 11 2 15 13 3 12 9 2
13 3 1 15 9 7 9 1 9 13 3 0 9 2
12 3 4 13 9 2 13 0 9 9 7 9 2
20 13 15 1 0 9 2 15 13 9 9 3 1 9 9 1 9 11 2 9 2
8 9 3 13 12 9 0 9 2
19 9 1 10 9 2 15 4 1 0 9 13 2 4 13 4 3 3 13 2
18 9 15 13 0 9 13 1 0 9 2 1 9 9 7 0 0 9 2
12 13 4 13 4 7 0 9 9 7 10 9 2
13 0 0 9 1 9 0 9 13 3 3 13 16 13
14 9 1 9 0 9 13 3 1 10 9 3 0 9 2
10 13 15 3 0 2 3 3 0 9 2
23 1 9 13 2 16 9 13 1 9 0 2 7 7 13 4 13 7 1 9 9 1 9 2
19 13 15 7 2 16 9 13 9 2 16 9 1 9 0 9 13 1 15 2
14 9 2 15 1 15 13 2 13 0 16 1 9 9 2
5 15 1 0 9 2
8 1 0 4 3 13 0 9 2
12 15 7 13 13 2 16 15 0 9 13 13 2
17 1 0 9 9 7 9 9 13 13 1 9 9 0 9 1 9 2
15 15 4 15 15 13 13 2 13 4 15 13 10 0 9 2
25 1 0 9 0 9 13 0 9 2 9 9 7 0 9 2 2 15 3 13 9 0 9 1 9 2
16 15 15 13 10 2 3 9 2 9 7 9 0 3 0 9 2
18 16 15 10 9 0 9 1 9 13 2 13 0 10 9 13 1 0 2
27 0 9 2 15 13 9 0 9 2 13 3 13 0 7 0 9 9 7 13 15 3 3 1 9 0 9 2
20 0 9 2 16 13 0 9 2 4 15 13 13 13 9 9 2 15 13 13 2
15 7 3 4 13 13 0 0 9 15 2 15 1 9 13 2
11 1 9 9 1 9 13 13 1 9 9 2
14 16 13 9 0 9 1 9 2 13 15 14 0 9 2
14 1 9 0 9 1 11 4 13 3 0 9 7 9 2
11 1 9 0 9 13 0 9 1 0 9 2
13 9 0 9 1 9 1 11 13 0 7 14 0 2
16 10 9 13 2 3 10 0 9 13 14 0 9 1 0 9 2
30 1 11 13 3 0 9 9 2 15 13 10 9 1 9 13 2 1 0 9 2 3 0 9 2 3 0 9 2 3 2
20 1 11 13 1 12 7 12 9 0 9 2 1 15 15 13 2 10 9 13 2
28 3 9 1 15 2 3 1 0 9 13 9 1 9 1 9 0 9 2 12 2 4 12 9 0 9 13 9 2
18 3 13 7 1 0 9 7 0 2 15 7 13 1 0 9 1 9 2
16 15 15 13 1 15 0 2 7 4 13 15 1 11 3 13 2
15 0 9 3 13 9 1 9 3 0 7 3 0 0 9 2
23 1 9 13 13 9 2 15 13 0 9 7 9 0 9 2 0 9 9 7 0 0 9 2
27 13 0 13 1 9 2 1 15 4 15 13 9 13 9 2 1 15 13 2 7 13 4 3 3 9 9 2
33 7 2 1 1 15 2 16 10 9 13 3 7 3 3 0 7 9 0 0 9 13 3 0 2 13 0 9 3 3 3 1 9 2
22 1 9 4 15 13 9 3 13 0 7 0 9 1 9 2 9 2 9 9 7 9 2
16 1 10 9 4 15 7 13 13 9 2 15 13 9 0 9 2
12 3 4 13 0 13 15 1 9 0 0 9 2
5 15 13 1 0 9
20 3 15 13 12 9 9 0 9 2 3 3 12 2 13 0 9 9 11 11 11
1 9
2 11 11
16 1 12 9 4 13 0 9 0 9 1 9 11 1 12 9 2
6 1 11 3 12 9 2
20 1 0 9 1 9 9 13 3 0 9 12 9 2 15 13 3 11 7 11 2
18 3 15 7 3 3 13 2 16 0 9 1 15 13 7 13 3 13 2
24 14 12 2 1 11 14 12 9 2 15 3 13 1 9 2 16 0 9 13 3 1 0 9 2
20 1 0 12 9 2 3 1 9 9 9 7 9 2 15 0 0 9 9 13 2
21 0 9 0 9 1 9 11 13 1 9 12 9 2 3 15 0 7 0 12 9 2
10 9 1 0 9 15 3 13 3 13 2
13 1 15 3 4 15 13 9 13 1 9 0 9 2
3 9 9 13
24 1 9 1 9 0 9 11 1 9 12 13 2 16 1 9 9 4 13 3 9 7 0 9 2
13 0 9 13 9 9 2 9 2 0 9 7 9 2
17 0 9 9 4 7 13 7 1 9 2 9 2 9 7 0 9 2
27 16 13 1 0 9 2 9 9 1 3 7 3 3 0 9 13 1 11 12 9 1 0 9 0 0 9 2
42 0 9 9 3 9 4 13 1 11 2 11 2 2 11 2 11 2 2 11 2 11 1 11 2 2 11 2 11 2 2 11 2 11 2 2 11 2 11 7 11 2 2
16 9 9 7 9 13 1 9 12 9 2 3 7 13 9 9 2
34 3 4 13 1 9 11 2 9 9 1 9 9 0 9 2 3 9 2 9 2 9 2 9 7 9 2 13 1 10 9 3 3 0 2
22 10 9 2 15 15 3 13 1 9 2 15 13 1 9 7 4 3 13 1 9 11 2
5 0 9 1 0 9
15 0 9 13 1 9 12 1 0 9 1 0 9 1 11 2
20 13 15 3 7 0 9 2 15 13 10 9 2 13 0 9 9 11 11 11 2
11 3 15 13 12 9 9 2 3 1 12 2
30 1 9 1 9 1 9 0 9 7 10 9 2 15 13 9 9 2 15 9 1 0 9 1 0 12 9 1 9 13 2
11 3 12 9 9 1 15 13 0 0 9 2
18 1 9 1 11 13 1 10 9 9 9 0 9 0 9 1 0 9 2
17 1 0 9 9 15 13 0 9 9 2 1 15 4 3 13 9 2
26 1 9 12 4 13 1 0 9 12 9 9 2 1 9 12 15 13 12 9 2 2 15 13 12 9 2
31 1 9 11 13 7 0 2 16 4 1 0 9 2 15 13 0 13 0 7 0 0 9 2 4 13 12 7 12 9 9 2
4 11 13 9 9
17 9 0 9 1 11 3 13 2 3 13 1 9 9 12 7 12 2
11 1 11 15 13 9 11 2 11 7 11 2
15 0 9 2 12 9 2 13 9 0 9 1 0 9 11 2
14 11 7 11 13 0 9 0 9 2 1 12 9 2 2
17 1 9 13 0 9 1 9 2 15 4 13 13 1 9 0 9 2
14 0 9 1 9 1 9 13 12 7 12 9 0 9 2
7 0 13 0 9 1 11 2
9 11 7 11 13 3 1 0 9 2
10 13 1 0 9 2 15 15 13 13 2
16 0 9 13 13 1 15 3 16 11 2 7 13 10 9 0 2
14 9 1 11 4 3 13 1 9 0 0 9 9 11 2
15 9 9 13 1 0 0 9 1 11 9 1 15 12 9 2
27 1 0 2 0 7 0 0 9 4 3 13 9 1 11 2 13 11 11 2 9 0 9 2 9 9 9 2
4 9 1 11 13
5 11 13 14 11 2
13 0 9 1 10 9 13 1 11 2 11 7 11 2
10 0 1 11 1 11 7 11 1 11 2
14 1 9 13 9 1 0 11 7 13 15 0 1 11 2
10 9 1 11 4 13 3 0 9 9 2
22 1 0 9 9 0 9 1 9 4 13 9 9 9 2 15 15 13 9 9 1 11 2
31 10 9 2 15 3 13 1 0 9 0 0 9 1 9 2 15 13 7 1 11 2 11 2 11 2 0 9 7 1 11 2
13 1 10 9 7 1 11 4 13 3 0 9 9 2
12 0 9 13 10 9 1 0 9 1 12 9 2
16 0 9 1 11 13 9 7 16 13 1 0 9 7 0 9 2
17 14 1 9 13 0 1 9 9 2 13 9 0 9 11 11 11 2
4 9 1 9 11
23 1 9 9 13 9 1 15 0 9 0 9 2 3 4 13 1 9 12 7 12 0 9 2
13 1 9 0 0 9 9 11 13 13 9 0 9 2
11 3 7 4 13 2 15 0 13 13 13 2
7 9 15 13 1 9 0 2
5 0 9 13 13 2
18 3 0 15 13 2 7 1 9 15 13 9 9 2 15 13 3 0 2
14 3 13 15 3 0 9 3 13 7 13 15 0 9 2
13 13 4 3 14 12 9 9 2 13 11 2 11 2
4 0 9 1 11
12 0 9 4 13 0 9 1 0 9 1 11 2
10 1 0 9 4 3 13 1 9 12 2
13 1 9 9 13 1 9 3 0 9 9 1 11 2
7 9 4 13 1 11 11 2
13 10 9 13 3 0 9 2 15 13 1 9 9 2
26 3 1 0 7 0 9 13 9 1 0 7 0 9 16 13 9 2 9 2 9 2 15 9 3 13 2
36 13 3 1 9 2 15 3 13 1 0 9 9 2 4 7 13 9 7 13 10 9 2 13 11 11 2 9 9 0 9 0 0 9 1 11 2
8 9 11 4 13 0 0 9 2
15 9 9 2 11 2 11 2 11 2 3 14 9 1 11 2
12 1 0 9 9 15 0 9 13 1 12 9 2
9 1 9 13 0 9 1 11 9 2
10 1 9 9 13 7 0 0 9 0 2
9 10 9 7 9 9 13 3 0 2
11 7 15 13 0 9 2 3 1 9 12 2
30 1 9 13 13 9 0 9 7 13 9 1 11 2 15 3 4 13 9 9 0 1 9 1 0 2 13 11 2 11 2
5 11 14 1 0 9
14 0 9 2 15 4 13 1 9 9 2 13 12 9 2
16 1 11 4 13 7 1 9 0 9 1 11 2 9 7 3 2
15 13 13 0 3 9 0 9 2 7 0 9 9 9 13 2
8 3 15 13 1 9 9 12 2
21 0 9 15 3 13 1 9 11 2 7 4 13 1 10 0 9 2 1 9 9 2
15 13 1 0 0 9 2 3 13 0 13 9 1 0 9 2
16 7 13 3 3 0 2 15 13 2 16 3 3 13 13 9 2
28 10 0 9 13 15 9 1 10 2 16 4 15 13 7 1 9 10 0 9 2 15 1 11 3 13 1 9 2
25 15 4 13 1 9 9 0 9 7 13 13 2 3 15 13 9 2 1 9 9 0 2 0 9 2
1 3
29 0 9 13 9 2 15 4 3 1 0 9 13 9 0 3 2 9 0 9 2 9 2 9 1 9 7 9 9 2
15 0 9 13 1 0 1 9 7 3 13 12 7 12 9 2
20 15 3 4 13 0 9 1 0 0 9 2 1 10 9 13 7 9 9 9 2
10 13 4 3 0 9 0 15 0 9 2
18 9 11 2 3 0 9 11 11 2 13 9 13 14 1 12 2 9 2
18 1 0 0 9 13 3 1 0 9 0 9 11 9 10 0 0 9 2
17 10 9 4 13 1 9 12 2 9 3 1 9 11 1 0 9 2
3 0 9 9
1 9
2 11 11
25 1 0 9 13 1 9 9 9 9 2 15 0 0 9 13 0 0 12 2 9 9 9 0 11 2
20 0 9 15 2 16 0 1 12 0 2 13 3 1 0 9 7 9 3 13 2
26 1 9 11 11 9 0 9 7 0 0 9 1 11 11 7 11 11 13 0 9 0 0 9 12 9 2
14 11 0 9 13 7 1 0 9 0 3 0 0 9 2
26 0 0 9 10 9 11 11 13 1 12 9 10 9 0 11 0 9 2 0 9 7 3 0 0 9 2
12 7 3 9 11 11 13 9 0 9 3 13 2
26 0 0 9 13 3 0 2 3 0 0 9 2 15 1 0 2 11 1 0 9 13 3 1 0 9 2
10 7 15 15 1 9 13 1 0 9 2
23 1 0 9 9 0 11 7 9 11 0 15 13 13 1 0 9 1 0 9 1 9 12 2
20 1 9 10 0 9 15 7 13 9 2 15 0 13 10 9 1 9 0 11 2
23 1 9 0 9 13 0 2 16 9 13 1 0 9 1 0 9 2 15 15 0 9 13 2
19 1 9 9 7 3 13 3 3 0 9 0 1 0 2 11 1 9 0 2
21 1 15 13 0 9 9 2 0 0 9 7 1 9 3 12 1 0 9 2 2 2
5 16 3 0 9 2
4 0 9 4 13
26 9 11 11 2 12 2 13 1 9 11 11 0 1 0 0 9 0 11 2 15 9 15 13 0 9 2
20 11 3 1 9 0 9 13 9 0 0 9 12 7 12 2 12 2 12 2 2
32 0 9 2 1 0 9 0 0 9 0 9 2 12 2 0 9 1 9 12 13 2 2 13 1 9 1 0 9 11 11 13 2
16 0 9 9 15 13 12 1 0 0 9 0 9 2 9 9 2
32 9 15 13 9 9 13 0 9 2 7 13 0 9 12 9 0 9 2 3 15 13 1 0 9 7 13 15 13 1 9 0 2
9 9 13 0 9 12 9 0 9 2
24 9 9 1 9 12 2 12 13 13 1 0 0 9 3 3 1 9 12 2 9 7 4 13 2
17 0 9 1 9 9 1 9 13 0 11 1 0 11 1 9 12 2
21 10 9 3 16 0 0 13 7 0 2 7 10 0 9 3 13 1 9 0 9 2
13 9 9 4 15 1 0 9 13 13 1 9 9 2
19 3 1 15 0 9 13 3 9 11 11 11 11 2 15 13 0 0 9 2
12 0 9 9 4 15 13 13 1 0 9 0 2
3 2 11 2
2 0 9
2 11 2
14 3 16 12 9 1 12 9 15 13 12 2 0 9 2
13 0 0 9 13 1 11 0 7 3 15 0 9 2
27 13 15 1 10 9 2 16 4 13 9 10 9 7 13 0 9 2 13 1 0 9 12 1 9 11 11 2
54 1 11 13 13 1 0 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 0 11 2 11 2 11 11 2 11 2 11 2 11 2 9 2 11 2 11 2 11 2 11 2 11 2 13 7 7 11 2 2
26 0 9 13 2 16 1 0 9 0 9 13 9 2 16 1 15 3 3 10 0 0 9 13 0 9 2
25 9 1 0 9 13 1 11 0 7 1 0 9 3 9 0 0 9 13 3 13 0 11 7 11 2
22 1 11 4 3 13 0 9 3 12 0 9 2 16 3 1 10 9 15 13 12 3 2
13 1 9 15 13 1 9 3 9 1 9 7 9 2
4 0 9 0 9
4 11 11 2 11
18 0 9 0 0 9 13 3 1 11 9 0 9 2 0 9 7 9 2
18 1 11 15 1 0 9 13 9 1 0 9 2 1 15 15 13 3 2
14 15 15 9 0 9 13 1 9 2 3 13 1 9 2
6 13 7 13 15 13 2
14 9 0 9 3 13 0 0 9 1 9 0 2 11 2
31 0 0 9 11 11 3 1 0 9 1 9 7 9 0 11 11 3 13 3 16 0 9 0 0 9 7 9 1 0 9 2
22 0 9 0 9 2 0 9 3 9 1 9 7 0 9 11 11 13 10 0 0 9 2
40 13 15 13 3 3 3 1 9 0 9 1 9 11 2 3 0 2 0 0 9 13 0 9 9 0 7 0 9 7 3 13 0 0 9 2 9 1 9 2 2
39 9 0 9 15 7 9 13 13 0 7 3 2 11 11 13 13 1 9 3 3 13 0 9 1 0 0 9 0 9 2 16 1 9 0 0 9 15 13 2
23 7 1 9 9 0 10 9 2 0 9 2 9 7 9 2 13 15 9 3 1 0 9 2
9 12 10 9 7 13 3 10 9 2
17 9 15 3 13 1 0 0 9 3 13 1 9 12 9 7 9 2
34 1 11 3 3 13 9 2 0 1 0 9 2 9 0 9 2 7 7 16 4 13 1 0 9 2 13 1 0 9 3 1 10 9 2
20 15 3 13 12 10 9 2 13 13 0 9 1 0 0 2 3 0 2 9 2
33 15 2 3 11 2 13 3 3 1 0 9 10 9 2 0 3 2 3 9 11 2 7 3 12 1 0 9 2 13 3 12 9 2
18 1 0 9 15 3 13 12 9 1 0 2 16 1 9 1 0 9 2
22 10 9 4 13 7 9 10 9 2 9 2 1 15 13 0 9 2 7 3 9 9 2
17 3 0 9 11 11 13 9 15 2 3 10 9 13 4 13 15 2
22 9 13 0 9 3 10 9 2 1 0 9 0 0 9 2 15 13 0 9 3 13 2
26 1 9 15 3 13 3 3 0 7 0 9 7 3 3 3 13 3 0 9 16 1 9 0 2 11 2
23 7 3 13 0 9 1 9 3 1 9 7 1 9 3 0 7 3 0 16 0 0 9 2
48 9 9 2 0 1 9 13 0 0 9 2 15 7 13 9 7 9 1 9 7 0 9 4 13 7 1 0 0 9 2 0 9 1 11 2 11 2 0 11 2 2 2 13 1 9 9 2 2
39 1 9 3 0 11 11 2 9 0 0 9 2 9 9 2 9 9 7 9 2 15 3 13 1 11 12 1 0 9 0 9 2 13 0 10 9 0 9 2
25 0 9 11 11 1 15 13 2 16 15 13 9 15 2 15 13 1 0 9 1 0 9 11 11 2
31 11 11 1 9 13 1 11 3 1 9 12 7 12 0 9 9 7 9 2 1 15 1 9 12 13 0 9 0 0 9 2
23 16 3 1 0 9 13 1 9 15 0 9 2 13 15 15 12 7 12 2 13 11 11 2
17 13 15 15 2 16 3 15 13 2 16 10 9 1 0 11 13 2
16 3 15 9 13 1 12 7 9 9 13 3 1 0 9 9 2
6 7 9 13 2 2 2
4 0 11 1 9
1 9
38 9 2 0 9 0 2 0 9 2 12 2 13 1 0 0 9 2 15 1 9 1 11 13 1 9 12 7 4 13 1 9 0 9 1 9 9 0 2
43 9 11 11 2 0 16 9 0 9 0 9 11 2 13 0 9 2 0 9 15 13 12 9 7 13 15 1 9 12 2 1 0 0 9 2 0 1 0 0 9 0 11 2
20 3 16 9 3 0 0 9 2 0 3 13 9 3 0 2 7 7 3 0 2
36 0 9 1 9 1 12 0 0 9 13 1 15 2 16 9 13 9 2 3 7 13 9 0 9 2 0 9 7 0 9 2 0 15 3 3 2
81 0 9 2 0 9 11 2 11 11 2 2 10 0 9 11 2 11 11 2 0 16 0 9 11 1 0 9 0 11 2 2 0 9 1 0 9 11 11 2 11 11 2 2 0 0 9 2 1 10 9 15 1 12 9 13 1 9 0 11 11 2 7 10 0 9 11 2 11 11 2 2 13 9 0 0 9 7 10 0 9 2
46 9 9 13 3 0 9 2 1 0 9 3 13 0 9 1 0 9 2 16 0 9 13 0 0 9 2 3 0 13 0 9 1 9 7 0 9 2 2 2 16 9 9 13 0 9 2
41 9 9 13 1 3 0 9 14 0 9 2 7 7 0 9 2 10 9 2 13 3 3 9 2 2 9 7 0 0 0 9 1 0 0 9 2 11 7 0 9 2
23 9 0 13 3 0 7 0 11 2 3 15 7 0 0 9 13 3 2 7 3 3 13 2
43 1 3 7 3 0 9 2 0 0 9 7 9 1 0 2 9 2 15 9 1 9 3 13 1 0 0 9 2 1 9 10 0 7 0 9 7 1 10 0 9 1 9 2
24 0 13 14 0 9 1 0 9 2 7 3 0 9 0 9 9 2 0 9 7 3 0 9 2
9 9 1 11 2 11 2 9 11 2
22 13 2 11 11 2 11 11 2 11 11 2 11 11 11 2 11 11 2 11 7 0 2
12 11 11 2 11 11 2 1 10 0 9 0 9
5 9 11 2 9 11
11 0 9 1 11 2 0 2 0 9 1 11
9 11 2 11 2 11 2 11 2 2
14 9 0 0 9 11 2 11 1 10 0 9 13 0 2
12 0 9 13 1 9 1 11 11 12 2 12 2
18 1 0 0 9 15 13 0 2 0 9 7 9 13 9 12 2 12 2
12 0 9 2 2 11 12 2 12 7 12 2 12
33 0 9 13 0 9 2 7 11 11 3 1 0 9 13 1 0 9 7 10 0 9 2 15 9 15 13 14 3 2 3 3 13 2
52 7 16 15 10 9 3 13 9 2 16 13 1 0 9 9 10 9 2 13 0 2 16 9 0 9 11 11 11 2 15 1 9 13 9 9 9 1 10 9 1 11 2 15 1 0 12 9 9 3 13 13 2
9 9 13 15 9 9 9 9 9 2
23 1 15 15 1 11 3 13 7 0 9 9 7 9 2 1 15 15 3 13 9 12 9 2
4 3 13 11 2
21 1 12 2 9 1 9 11 13 3 0 9 1 9 3 0 12 0 9 11 11 2
30 9 9 3 13 9 3 15 0 0 9 7 1 9 0 9 15 9 1 9 0 12 13 1 0 0 9 13 11 11 2
31 1 0 9 1 9 2 15 15 13 1 9 1 0 0 9 2 13 9 11 11 0 9 9 3 2 10 9 13 3 13 2
15 13 15 3 1 9 9 2 1 15 15 13 9 0 9 2
11 10 9 13 1 9 1 0 9 0 12 2
18 3 11 13 0 9 1 0 9 7 13 3 3 0 9 0 0 9 2
11 3 11 3 13 3 0 0 9 11 3 2
19 1 9 7 3 13 3 9 7 15 1 10 9 13 2 3 0 13 9 2
28 1 12 2 9 13 0 9 9 2 1 15 13 11 2 11 7 11 2 11 0 9 7 11 12 5 12 9 2
25 1 9 3 4 3 13 1 9 11 7 11 15 13 12 9 1 9 1 0 9 12 1 12 13 2
11 1 10 9 15 13 7 11 13 1 9 2
16 0 9 11 7 3 13 1 15 2 16 13 13 1 0 9 2
18 1 10 9 15 3 1 9 13 2 7 10 9 0 9 9 3 13 2
19 0 9 13 9 1 0 9 7 0 9 1 9 11 3 1 12 9 9 2
18 3 16 1 11 13 2 3 7 1 0 0 9 2 9 1 0 9 2
35 11 15 13 13 3 1 9 0 12 2 7 16 11 1 12 2 9 3 13 9 1 10 9 2 13 15 2 16 15 11 13 7 0 9 2
12 1 7 13 11 11 2 15 13 0 9 11 2
13 1 12 9 13 0 9 2 3 1 9 15 9 2
62 13 2 16 16 15 4 1 0 9 13 7 9 2 13 10 9 3 2 13 3 1 11 9 11 11 2 1 0 9 15 13 2 16 9 13 9 2 15 13 0 2 3 2 9 2 7 13 9 1 9 2 15 15 13 13 2 3 9 7 0 9 2
11 13 15 7 0 9 7 15 13 9 9 2
10 0 9 4 3 1 11 13 9 3 2
3 11 4 13
4 11 2 11 2
37 0 9 11 11 13 3 1 9 0 9 11 2 0 9 9 9 9 12 1 11 2 11 0 2 7 10 9 1 9 4 13 1 0 9 10 11 2
28 9 9 13 1 15 2 16 0 0 9 1 0 9 9 13 10 9 9 7 11 3 13 1 10 9 0 9 2
11 9 9 13 7 9 0 0 9 11 11 2
25 9 0 9 11 15 3 13 0 0 9 11 11 1 11 7 13 0 9 1 0 9 1 12 9 2
5 1 9 13 7 9
7 11 13 0 11 1 0 9
5 11 2 11 2 2
19 0 9 0 9 2 15 13 9 0 0 9 2 15 13 12 0 11 11 2
17 1 11 13 1 10 9 3 1 11 11 2 11 11 7 11 11 2
20 1 9 9 11 15 3 13 11 11 2 15 13 1 0 0 9 7 9 9 2
42 11 11 15 13 1 11 2 3 3 13 1 9 2 1 9 1 9 3 13 9 11 7 1 9 1 0 9 2 9 9 2 9 2 13 3 3 0 0 9 1 11 2
21 3 13 0 9 2 15 13 0 9 2 9 1 9 7 13 15 0 9 7 9 2
12 15 3 1 9 13 9 13 15 1 0 9 2
23 1 11 4 16 9 13 3 3 0 9 1 9 7 11 15 1 10 9 13 3 0 9 2
35 3 4 13 2 13 11 11 2 15 1 9 12 3 13 1 9 7 0 9 1 9 13 9 7 1 0 0 9 9 1 9 11 1 11 2
23 1 10 9 13 9 11 11 2 15 15 7 13 1 0 9 7 13 0 1 11 13 9 2
18 11 15 3 1 9 9 13 1 11 2 3 15 1 9 13 13 3 2
6 1 9 13 15 0 2
27 1 11 2 11 7 11 13 1 9 3 14 0 9 7 13 2 16 4 15 13 2 16 1 15 15 13 2
6 7 15 3 13 3 2
27 1 0 9 15 14 10 0 9 13 2 16 1 9 2 15 15 13 1 9 2 13 3 0 9 2 2 2
4 9 9 1 11
7 11 1 11 2 11 2 2
22 0 9 1 12 2 9 0 9 0 9 13 1 9 0 9 11 2 1 9 1 9 2
21 9 9 11 11 11 1 0 9 14 1 0 9 9 13 3 9 2 3 0 9 2
14 10 9 13 1 0 0 9 7 9 9 2 9 9 2
14 1 1 9 0 9 4 1 0 9 10 9 13 9 2
18 1 0 9 15 0 9 1 9 0 2 0 9 13 1 3 0 9 2
33 1 9 1 9 9 1 9 13 3 9 1 9 2 1 9 1 0 9 7 1 9 1 0 9 2 15 3 13 9 0 0 9 2
24 15 9 7 13 13 9 9 11 11 2 15 13 3 3 1 9 3 0 9 1 9 11 11 2
17 15 1 0 9 2 9 1 9 7 12 9 9 13 9 9 9 2
8 9 13 1 9 3 0 9 2
3 11 1 0
2 11 2
16 0 9 11 1 11 2 0 9 11 11 2 4 13 1 9 2
32 0 9 15 13 12 2 9 1 0 9 9 11 1 0 2 11 1 11 0 9 2 15 9 13 9 1 11 0 0 9 9 2
30 1 9 0 0 9 2 11 2 15 7 15 13 2 11 3 13 10 9 1 0 9 2 3 3 15 13 1 0 9 2
11 1 9 0 0 9 15 7 13 1 9 2
9 9 0 9 1 0 9 3 13 2
38 7 3 1 9 13 13 2 16 0 9 9 9 1 9 12 2 12 11 11 11 13 0 9 9 2 13 13 12 9 2 1 0 9 15 13 12 2 2
20 16 4 15 1 9 9 9 9 13 1 0 9 0 9 2 13 15 0 9 2
5 0 9 13 1 0
2 11 2
11 0 9 1 11 13 12 1 0 1 9 2
15 1 0 9 3 1 0 12 9 1 9 13 3 12 9 2
9 9 0 9 1 0 9 13 12 2
8 1 9 0 15 13 13 12 2
12 9 0 9 13 1 0 9 1 12 1 12 2
25 3 9 13 1 11 7 1 11 11 0 11 2 3 13 3 16 9 1 0 12 9 0 0 9 2
25 9 1 9 13 0 9 9 0 9 2 0 9 7 0 9 0 9 2 15 13 0 9 9 0 2
5 14 0 9 0 13
30 9 1 10 2 16 15 3 1 9 0 7 0 2 11 12 2 12 2 2 15 13 10 0 9 7 9 1 0 9 2
28 13 15 3 9 1 0 2 13 0 9 2 7 16 9 13 1 0 2 15 2 1 9 2 1 10 9 13 2
15 16 15 9 13 1 10 0 2 7 13 2 3 15 13 2
20 14 1 9 13 10 0 9 9 2 15 15 13 7 13 15 0 2 7 13 2
8 3 1 10 0 9 13 13 2
17 13 9 1 9 1 10 9 1 9 9 2 16 15 13 3 9 2
4 13 15 0 2
28 0 9 13 0 9 0 9 1 0 9 9 2 15 3 13 0 2 0 9 2 9 9 1 9 7 0 9 2
21 0 9 13 1 0 9 1 9 2 1 15 13 9 7 9 2 7 3 3 13 2
25 3 3 13 9 1 9 2 3 13 13 7 1 9 0 9 7 15 9 15 2 15 13 1 9 2
16 1 9 3 9 7 0 9 2 1 9 9 9 7 0 9 2
10 1 12 9 15 13 1 9 1 9 2
19 16 9 1 9 13 7 15 1 9 13 2 13 1 9 2 3 15 13 2
23 13 13 9 7 9 2 3 4 15 13 9 7 9 1 9 2 16 10 0 9 15 13 2
12 7 13 13 7 9 1 9 2 7 7 9 2
25 13 1 15 0 9 1 9 2 16 15 1 9 0 9 13 7 1 12 0 9 7 15 13 9 2
4 9 13 0 2
38 9 9 13 0 2 13 0 7 13 1 10 9 3 2 3 2 10 9 9 2 9 0 9 7 9 2 3 0 9 2 16 4 1 15 15 3 13 2
23 0 9 13 0 7 1 9 2 15 13 15 2 13 10 9 7 10 9 2 1 0 9 2
23 13 15 7 1 0 2 16 15 1 15 13 2 13 9 2 13 2 7 3 15 15 13 2
37 1 9 0 9 4 13 1 10 9 1 9 13 7 0 9 2 0 9 2 13 4 15 13 10 9 2 16 4 13 9 1 9 9 10 0 9 2
6 11 2 11 2 2 11
3 11 15 13
2 11 2
23 11 2 15 13 3 1 0 9 11 9 1 9 1 9 12 2 15 13 13 1 9 12 2
5 9 0 16 9 9
5 11 2 11 2 2
36 9 11 15 13 2 16 13 9 9 0 9 11 11 11 0 2 9 2 11 11 2 15 15 13 9 9 16 9 1 9 9 1 9 0 9 2
31 13 4 15 2 16 9 9 1 10 9 2 1 15 15 0 9 1 9 10 9 13 2 4 15 13 3 1 12 9 9 2
29 9 9 9 11 4 3 13 0 9 2 7 15 4 13 1 9 1 9 1 9 2 13 15 9 9 11 11 11 2
14 16 9 0 9 13 2 3 1 15 4 13 0 9 2
8 12 1 9 13 7 9 9 2
31 1 0 9 11 12 13 0 9 1 9 1 9 2 16 15 0 9 13 0 0 7 0 9 1 10 9 2 13 9 9 2
12 9 11 15 13 2 7 13 2 16 1 9 13
7 11 2 11 2 11 2 2
15 13 4 15 2 16 10 9 1 9 9 0 9 13 0 2
17 13 15 0 2 16 10 2 7 0 9 4 15 13 13 3 9 2
24 1 0 9 15 13 9 2 9 11 9 11 7 15 9 9 1 11 7 11 11 11 2 12 2
22 1 10 9 13 1 9 3 9 9 0 9 11 11 1 9 1 9 1 0 9 9 2
26 15 15 13 9 9 2 1 15 9 13 0 9 1 9 3 2 16 15 13 0 9 1 0 0 9 2
39 9 15 13 2 16 4 13 13 9 14 1 9 1 0 9 9 2 7 14 3 2 3 13 15 1 15 1 0 9 9 2 1 9 9 1 0 0 9 2
22 7 13 1 11 11 7 13 2 16 16 4 10 9 13 2 13 7 1 10 0 9 2
36 1 0 9 0 9 11 9 11 1 9 9 2 11 2 11 2 11 2 11 2 15 1 9 9 11 11 1 0 9 13 3 1 0 9 9 2
17 13 4 15 3 1 15 2 16 0 9 4 13 1 0 0 9 2
12 0 9 13 7 9 2 13 15 0 0 9 2
13 1 15 4 13 0 9 2 15 15 15 4 13 2
8 9 13 3 2 3 15 13 2
14 13 2 16 15 13 3 1 9 9 2 13 11 11 2
19 1 9 2 16 4 9 3 13 1 3 0 9 1 11 2 13 2 3 2
25 0 9 7 13 9 14 1 9 1 11 7 9 11 11 13 2 13 2 16 1 9 13 0 9 2
17 1 9 2 16 13 3 9 3 1 9 2 13 2 13 15 13 2
17 3 2 13 3 2 9 2 9 2 2 15 9 13 7 4 13 2
15 7 1 0 9 9 9 1 9 9 7 9 1 11 13 2
26 15 3 2 16 11 11 1 9 2 16 13 0 9 0 13 1 9 9 2 13 2 10 9 13 0 2
3 11 13 11
2 11 2
30 0 0 9 13 0 9 11 12 9 2 12 9 2 1 9 1 0 9 1 11 2 15 15 13 12 2 9 1 11 2
18 0 9 3 13 11 13 1 0 9 7 13 1 10 9 3 0 9 2
41 0 9 11 11 2 9 0 9 9 7 1 0 9 9 9 1 0 0 9 2 9 13 2 7 13 2 16 15 3 1 10 9 13 11 13 1 9 1 0 9 2
14 9 11 1 0 9 1 9 1 11 13 12 2 12 2
2 11 13
2 11 2
19 12 1 0 0 9 11 11 13 1 0 9 1 11 2 16 13 0 9 2
21 3 3 13 9 7 0 4 13 2 7 9 15 15 13 2 13 9 9 11 11 2
6 11 13 9 0 9 2
12 13 15 0 9 9 2 3 15 9 13 9 2
4 11 11 13 9
3 0 11 2
13 0 9 0 9 11 11 15 13 9 0 0 9 2
17 1 0 9 13 1 10 0 9 1 9 7 9 1 9 11 11 2
8 11 13 1 0 9 10 9 2
16 13 9 0 9 3 2 16 4 15 0 9 13 3 16 3 2
3 0 9 11
2 11 2
25 0 9 11 11 2 15 0 0 9 13 1 9 2 15 3 3 13 1 9 9 1 9 0 9 2
18 13 2 16 15 13 13 7 16 9 10 9 11 13 15 9 1 9 2
40 11 4 13 1 9 9 2 15 13 0 0 9 1 9 0 9 2 0 0 9 2 11 2 7 0 0 9 2 11 2 7 10 9 13 2 16 13 1 9 2
6 15 13 3 0 9 2
18 0 9 13 3 10 9 0 0 9 7 9 13 0 9 1 10 9 2
12 13 0 9 3 15 1 9 7 3 13 9 2
19 13 2 16 9 1 12 2 9 4 13 1 0 9 1 0 9 1 9 2
3 1 0 9
86 9 11 11 13 9 1 0 9 9 1 9 1 9 2 11 2 11 2 2 11 2 11 2 2 11 2 11 2 2 11 2 9 2 2 11 2 11 11 2 2 11 2 11 2 2 11 11 2 11 2 2 11 2 11 2 2 11 2 11 2 2 11 2 11 2 2 11 2 9 2 2 0 2 11 2 2 9 2 11 2 2 11 2 11 2 2
11 0 0 9 11 11 13 0 9 11 11 2
16 11 11 2 1 15 11 13 2 13 9 1 9 12 9 9 2
4 9 1 0 9
2 11 2
31 0 9 0 0 9 13 1 0 9 12 2 0 9 2 15 15 9 9 1 9 0 0 9 1 0 11 13 0 0 9 2
9 9 15 4 13 3 12 0 9 2
25 0 13 13 1 0 9 2 0 1 9 0 9 2 0 1 0 9 9 7 0 1 0 0 9 2
10 9 15 13 3 3 3 13 0 9 2
13 9 15 13 7 1 9 2 9 7 0 9 9 2
23 13 15 4 3 1 9 2 15 15 3 13 10 0 9 7 4 7 13 0 9 7 9 2
4 11 13 0 9
3 0 11 2
23 1 3 0 9 4 13 0 0 0 2 15 13 1 0 11 9 0 9 1 9 1 9 2
14 0 9 0 9 11 7 11 3 13 10 9 0 9 2
28 15 4 13 13 1 9 3 2 0 9 11 11 2 15 1 9 9 13 1 11 3 16 3 1 12 2 9 2
12 11 11 2 12 2 0 2 13 3 1 9 2
7 13 13 2 13 1 9 2
18 13 4 2 16 15 10 9 13 2 7 13 15 3 15 3 15 0 2
8 9 3 13 2 13 0 9 2
6 13 15 11 11 11 2
27 1 0 9 2 0 1 12 9 9 2 13 0 9 11 2 11 1 11 11 12 2 12 2 12 2 12 2
28 3 1 15 15 1 9 1 0 11 13 11 11 2 15 9 3 13 2 12 2 12 2 7 3 13 1 9 2
29 9 9 15 1 0 9 13 0 9 16 1 0 9 2 11 11 11 2 15 1 9 13 1 0 9 1 9 13 2
6 9 12 9 1 11 2
8 0 11 13 1 9 0 11 2
5 9 11 11 2 11
5 7 9 13 9 9
15 9 0 9 0 0 9 2 11 11 2 11 11 12 2 12
7 11 2 11 2 11 2 2
15 1 0 9 15 9 11 13 9 1 9 12 2 0 9 2
11 1 11 13 0 9 0 11 12 2 12 2
6 1 9 9 13 11 2
20 1 0 9 1 9 9 13 0 9 11 2 7 1 0 9 14 13 9 9 2
15 3 13 11 9 2 15 13 1 0 9 1 9 0 15 2
22 1 12 2 9 13 9 0 9 1 0 9 11 7 0 11 13 9 2 12 2 12 2
20 7 3 13 0 9 1 9 11 2 10 0 9 13 1 0 9 1 15 9 2
12 3 16 12 12 9 15 13 3 1 15 13 2
12 1 9 11 13 0 0 9 2 15 11 13 2
20 1 9 11 13 9 9 7 11 13 0 9 1 9 9 2 7 13 0 9 2
25 1 12 2 9 2 13 9 2 11 15 13 1 0 9 2 13 11 7 13 11 2 12 2 12 2
6 0 7 13 15 9 2
20 1 12 2 9 2 13 11 14 3 13 11 9 7 11 1 9 13 1 9 2
18 1 12 9 3 11 13 0 9 2 13 15 1 11 7 15 13 13 2
18 1 9 1 10 13 11 1 0 9 11 2 7 9 15 9 13 3 2
35 11 13 15 1 9 2 13 15 9 0 9 2 0 9 13 11 2 11 1 0 9 13 9 2 2 7 7 11 13 1 0 9 0 9 2
7 9 9 15 7 3 13 2
20 1 9 1 9 15 9 11 13 13 1 9 2 16 15 3 13 1 15 13 2
12 1 9 10 9 15 3 13 9 12 12 9 2
15 13 3 9 11 2 15 7 3 13 7 1 9 0 9 2
12 11 11 2 1 0 9 4 13 0 9 3 2
15 13 4 0 9 2 16 15 15 13 3 13 0 9 11 2
16 11 2 9 11 2 11 13 3 2 16 13 0 9 1 9 2
15 16 4 11 13 0 9 2 11 4 15 1 9 3 13 2
14 11 11 2 9 11 2 13 4 12 9 1 0 9 2
12 16 13 11 1 10 9 2 13 13 1 9 2
4 9 13 0 2
2 0 9
1 9
31 1 0 9 4 9 13 1 9 0 9 13 9 12 2 9 11 2 11 2 15 0 13 1 9 9 11 3 12 2 12 2
9 13 15 7 13 9 1 0 9 2
5 9 1 9 9 2
3 0 9 9
4 15 4 13 2
35 1 12 2 9 9 1 12 2 9 13 12 9 1 12 9 2 1 12 2 12 9 1 12 9 2 1 0 9 13 12 9 1 12 9 2
21 1 9 1 12 2 9 13 10 9 2 1 12 2 9 13 12 9 1 12 9 2
55 1 12 2 9 11 1 12 2 9 13 9 2 1 12 2 9 13 12 9 12 9 2 1 12 2 9 13 12 9 1 12 9 2 1 12 2 9 13 12 9 1 12 9 2 1 12 2 9 13 12 9 1 12 9 2
59 1 12 2 9 11 1 12 2 9 13 12 9 12 9 2 1 12 2 9 13 12 9 1 12 9 2 1 12 2 9 13 12 9 1 12 9 2 1 12 2 9 13 12 9 1 12 9 2 1 12 2 9 13 12 9 1 12 9 2
34 1 9 12 1 12 1 12 2 9 13 9 2 1 12 2 9 13 12 9 1 12 9 2 1 12 2 9 13 12 9 1 12 9 2
53 1 9 1 12 2 0 9 13 9 2 1 12 2 9 13 12 9 1 12 2 1 12 2 9 13 12 9 1 12 9 2 1 12 2 9 13 12 9 1 12 9 2 1 12 2 9 13 12 9 1 12 9 2
5 3 1 11 1 11
11 11 13 13 9 2 15 13 1 9 15 13
7 11 2 11 2 11 2 2
18 0 0 9 13 1 15 1 9 0 0 9 11 2 11 0 12 9 2
31 0 9 2 12 2 12 2 7 0 9 2 12 2 12 2 15 3 16 10 0 9 13 2 7 1 0 9 13 3 0 2
44 16 0 9 11 11 13 1 9 11 3 0 9 2 15 13 0 9 1 0 9 9 1 11 2 11 15 13 1 0 0 9 3 12 9 2 9 11 2 9 11 7 9 11 2
39 1 12 9 2 11 2 11 2 11 2 13 9 12 9 7 0 9 2 1 15 1 9 4 15 9 1 0 9 1 9 0 9 13 13 1 9 12 9 2
24 0 9 13 1 15 2 16 15 0 9 13 13 1 9 7 1 9 13 15 2 13 11 11 2
9 9 9 13 1 15 3 0 9 2
11 13 15 13 9 3 1 9 7 1 9 2
18 10 9 13 9 1 10 9 2 15 13 9 1 9 15 13 2 13 2
10 3 3 13 0 9 0 0 9 9 2
33 1 11 13 1 0 0 9 1 11 2 15 1 0 9 13 12 0 9 1 0 9 1 11 1 9 12 2 12 7 12 2 12 2
17 9 2 15 13 1 12 9 0 9 1 0 9 2 13 0 9 2
21 11 15 3 13 13 15 1 9 1 0 9 1 12 2 9 2 12 2 12 2 2
17 11 13 3 3 16 11 2 16 13 9 1 10 9 7 0 9 2
15 13 1 11 1 0 2 7 14 1 0 9 2 13 11 2
31 9 0 9 13 12 9 11 1 9 1 11 2 11 2 13 15 1 11 11 2 7 11 11 2 13 13 3 1 11 2 2
16 1 9 15 13 11 11 2 11 2 7 11 11 2 11 2 2
18 13 4 9 11 11 2 11 2 2 15 14 3 13 1 9 1 11 2
22 11 11 15 3 13 1 9 0 9 11 2 15 10 9 13 1 9 1 9 9 9 2
21 7 16 4 15 1 9 9 9 11 9 1 9 7 9 13 2 10 9 11 13 2
6 13 3 1 9 9 2
3 11 1 11
5 11 2 11 2 2
11 0 9 11 11 11 11 13 1 0 11 2
17 1 10 0 0 9 15 13 0 9 1 11 11 1 9 10 9 2
18 1 9 13 11 1 9 3 15 13 2 16 15 11 13 1 0 9 2
22 11 3 13 9 2 15 13 13 1 10 9 12 12 9 2 1 11 3 12 12 9 2
4 9 12 2 9
42 0 0 9 13 3 3 12 9 12 2 9 2 11 2 11 2 11 2 11 2 11 2 0 11 2 11 2 11 2 11 2 11 11 2 11 2 11 2 15 12 2 2
30 0 12 9 15 13 1 9 2 11 2 11 2 12 9 2 2 13 9 11 2 2 11 2 11 2 12 9 2 2 2
35 1 9 13 9 9 2 7 0 9 13 9 1 0 9 9 9 1 9 2 15 13 1 9 1 9 12 2 9 1 12 9 1 0 11 2
17 0 9 12 2 9 13 3 3 1 0 9 1 9 11 2 11 2
3 2 11 2
5 11 11 13 1 11
5 11 2 11 2 2
11 0 9 11 11 7 3 13 9 0 11 2
39 1 11 15 3 12 2 9 13 9 2 7 2 13 9 10 9 2 1 9 4 13 4 9 13 2 13 15 9 11 11 11 2 15 7 9 0 9 13 2
13 13 4 15 2 16 1 9 0 9 13 9 9 2
8 13 11 13 9 1 0 9 2
11 3 4 1 9 13 7 1 9 0 9 2
16 13 7 2 16 1 9 0 9 1 9 13 3 0 1 9 2
5 9 7 9 9 11
10 9 1 9 11 2 11 15 13 12 9
5 11 2 11 2 2
15 14 3 3 9 13 1 9 9 11 1 0 9 1 11 2
22 16 13 3 16 9 9 1 3 0 9 2 1 9 13 9 1 0 9 12 2 12 2
19 12 9 13 1 9 9 1 0 9 10 9 1 7 1 9 11 1 11 2
37 0 11 11 13 2 3 10 9 13 1 0 9 13 1 10 9 2 16 1 9 2 11 1 11 15 3 13 1 9 1 9 9 1 12 2 12 2
21 9 13 2 16 11 1 9 3 13 9 9 2 16 0 3 13 7 3 3 13 2
14 1 9 9 7 11 13 1 9 7 13 15 9 9 2
9 1 12 0 9 13 3 13 9 2
25 13 4 9 7 9 2 13 15 14 3 12 1 12 2 13 9 11 2 15 9 10 9 14 13 2
17 9 1 15 13 1 0 9 1 9 2 16 15 4 13 0 9 2
8 1 10 9 4 3 13 9 2
30 9 9 4 15 3 13 1 0 9 2 3 15 1 9 1 0 9 13 9 1 9 2 7 3 3 4 15 13 13 2
7 9 12 2 9 12 2 9
19 9 2 12 2 1 15 11 2 11 11 2 12 2 11 2 11 2 12 2
21 0 9 2 12 2 3 11 7 11 2 12 2 2 3 11 7 11 2 12 2 2
22 0 9 2 12 2 11 2 11 2 7 11 2 11 2 2 3 3 4 13 12 9 2
18 0 9 2 12 2 9 2 3 2 11 11 2 11 2 12 9 2 2
9 0 9 13 1 9 3 1 9 2
5 2 11 2 11 2
4 11 13 11 3
8 1 11 13 9 1 9 1 11
5 11 2 11 2 2
25 3 1 9 0 12 0 9 13 9 11 9 0 9 2 3 13 3 0 2 1 0 9 1 11 2
15 14 3 2 1 9 1 11 2 13 13 2 3 3 13 2
28 16 1 15 13 9 9 1 12 2 9 1 11 2 13 3 0 0 9 1 0 9 9 1 9 12 2 12 2
10 1 9 15 13 9 0 9 1 11 2
14 1 0 9 7 9 1 0 9 4 3 13 11 13 2
22 1 9 12 2 12 7 13 9 2 1 15 15 13 13 2 13 15 9 11 11 11 2
19 1 0 0 9 1 9 1 11 2 12 2 12 2 13 1 10 0 9 2
12 9 13 1 10 9 2 13 7 1 0 9 2
17 13 7 0 9 2 16 4 15 13 10 9 7 13 9 1 9 2
7 3 13 1 9 1 9 2
19 15 4 13 10 9 2 7 0 12 9 13 2 15 13 3 2 13 9 2
16 9 11 11 13 1 9 1 11 13 2 16 9 13 3 3 2
13 13 4 3 9 2 7 9 4 15 13 3 10 2
23 11 13 7 3 13 0 9 2 16 13 1 0 9 9 7 13 4 3 12 9 1 9 2
29 16 9 7 13 13 12 7 12 9 1 9 9 2 15 15 13 2 13 9 1 9 11 2 15 4 1 9 13 2
41 9 0 11 11 11 13 9 1 0 9 2 15 7 13 9 1 10 0 9 2 1 9 11 13 3 0 9 2 7 13 15 3 2 16 4 13 3 1 10 9 2
13 13 4 3 2 16 4 13 1 12 9 1 11 2
34 0 13 1 9 11 7 11 2 7 3 1 0 9 0 9 11 2 15 1 9 9 3 1 0 9 13 1 9 14 1 12 2 9 2
18 13 15 14 3 2 7 13 2 16 13 9 1 9 9 7 1 9 2
12 3 4 15 13 13 0 9 9 2 13 11 2
5 11 13 1 9 9
29 1 0 9 7 3 7 1 9 1 9 0 9 13 1 12 2 9 0 0 9 0 9 1 0 9 2 0 9 2
13 3 1 0 9 9 13 0 11 2 15 3 13 2
9 7 3 10 9 15 1 9 13 2
18 3 13 2 1 11 4 13 9 2 13 1 9 9 0 9 11 11 2
14 9 14 13 3 2 7 0 9 3 13 12 2 12 2
11 13 14 9 9 2 3 15 11 13 13 2
39 9 15 1 9 3 13 2 1 9 1 0 2 9 13 7 9 0 11 2 9 2 9 2 2 7 15 15 13 9 13 2 13 11 0 9 10 0 9 2
3 11 3 9
28 0 11 2 15 1 9 13 1 11 2 13 9 12 2 12 1 0 11 2 16 4 13 1 0 9 1 9 2
24 3 3 13 0 9 1 9 7 13 1 12 9 12 9 2 15 15 13 1 0 9 1 9 2
13 13 15 9 9 2 7 4 13 3 1 0 9 2
29 0 13 9 2 0 12 2 9 2 9 2 2 7 3 15 13 7 9 2 13 15 9 9 11 2 11 11 11 2
25 16 10 9 1 0 9 11 11 3 13 2 0 13 3 2 7 13 4 15 15 9 1 0 9 2
15 1 0 9 15 13 11 11 1 9 12 2 12 1 11 2
21 11 13 2 15 13 10 0 9 2 9 11 2 9 1 11 2 15 3 13 9 2
3 0 0 9
48 7 11 1 9 0 9 1 11 3 13 2 12 2 12 1 11 2 2 16 13 1 9 9 1 9 9 2 9 13 1 0 9 9 1 9 7 11 1 11 13 1 9 1 9 1 0 11 2
11 11 13 0 0 9 7 13 15 12 9 2
15 12 1 15 13 9 11 2 0 13 10 9 1 0 9 2
16 1 0 9 13 1 11 0 9 2 15 3 13 12 2 12 2
16 0 9 0 13 0 9 1 9 11 2 13 0 9 11 11 2
12 9 13 2 16 11 15 0 9 13 0 9 2
6 3 13 9 0 0 2
23 9 2 16 3 13 1 10 9 9 11 2 3 13 13 9 0 2 13 0 9 11 11 2
13 11 13 3 15 1 9 11 2 7 7 3 13 2
14 3 3 15 13 13 11 1 9 12 2 12 1 11 2
16 0 9 11 11 4 1 9 13 1 12 2 9 9 1 9 2
20 1 9 0 11 11 13 7 9 9 11 9 7 13 1 15 9 1 9 9 2
15 11 14 13 12 9 2 10 0 9 7 9 13 1 9 2
4 11 1 9 9
27 0 13 9 11 2 3 1 9 11 1 9 2 1 11 2 1 15 9 3 13 0 2 12 2 12 2 2
14 13 4 3 0 9 2 7 1 9 4 13 14 0 2
16 13 4 15 3 9 2 13 0 0 9 11 11 2 11 11 2
37 1 15 13 3 0 9 11 11 2 15 13 2 1 9 9 15 13 0 9 0 9 2 15 15 13 12 9 1 0 9 11 11 1 9 1 11 2
31 11 13 1 10 9 9 9 1 0 9 2 7 1 9 9 9 11 11 15 9 13 1 0 9 0 9 7 13 1 11 2
11 7 1 9 15 13 13 14 1 9 9 2
28 0 9 11 11 3 13 2 9 11 4 13 1 9 9 9 7 4 15 13 1 9 9 2 1 15 15 13 2
22 1 12 9 1 11 2 11 7 1 11 3 13 11 2 16 9 1 0 9 13 3 2
29 11 15 3 13 9 0 9 1 12 2 9 2 7 0 13 9 12 9 1 9 12 9 1 9 0 7 0 9 2
27 1 0 9 12 2 12 1 11 7 0 9 12 2 12 15 1 9 13 9 1 9 2 16 4 3 13 2
38 3 4 7 13 13 9 2 13 15 0 9 2 16 0 11 11 13 13 2 13 15 9 11 2 7 15 15 13 1 12 2 9 2 3 9 13 11 2
14 3 0 9 2 13 2 1 9 11 9 7 4 13 2
14 11 15 1 0 9 1 11 2 11 13 9 1 9 2
22 9 12 2 12 13 1 0 9 1 11 3 0 1 9 9 2 13 9 9 11 11 2
9 2 11 2 11 2 11 2 11 2
3 11 13 3
5 11 2 11 2 2
13 11 11 13 1 9 3 3 0 11 1 0 9 2
16 1 12 9 15 13 9 9 7 13 15 15 0 9 11 11 2
13 3 15 7 3 13 7 3 0 9 1 9 13 2
11 1 9 15 1 9 13 13 3 1 11 2
9 7 3 13 9 7 13 0 9 2
20 0 9 1 9 11 13 10 9 9 2 15 13 9 11 1 11 12 2 12 2
28 12 9 4 13 2 7 14 1 9 11 11 4 15 13 2 16 1 11 15 13 1 0 9 3 16 1 11 2
25 3 4 7 3 13 1 11 12 9 7 15 3 4 15 3 13 1 15 2 16 15 13 1 9 2
13 3 4 13 1 9 9 1 11 2 15 15 13 2
15 0 2 15 13 9 2 14 10 0 0 9 15 3 13 2
16 7 1 9 1 9 15 15 13 2 16 4 10 9 3 13 2
4 3 1 11 2
12 13 4 2 16 15 9 13 1 9 9 9 2
17 13 4 1 9 9 13 12 9 2 7 9 1 15 0 13 0 2
14 0 13 2 16 13 0 13 9 14 1 11 2 2 2
4 6 2 6 2
9 13 15 3 2 7 15 13 0 2
13 0 14 2 7 3 3 3 16 9 1 11 13 2
10 9 13 1 9 9 7 3 15 13 2
23 3 13 3 2 7 16 15 1 9 13 2 3 4 13 13 15 2 15 15 1 15 13 2
12 1 9 13 11 1 11 2 13 7 15 9 2
14 16 15 9 13 2 3 1 0 9 1 9 7 13 2
23 7 15 13 12 2 15 13 9 2 0 13 13 7 9 9 2 15 13 14 1 0 9 2
9 11 13 1 9 2 7 15 3 2
11 1 9 15 9 13 2 15 13 14 13 2
6 15 13 3 0 9 2
11 1 11 4 9 13 3 14 1 9 9 2
9 9 1 9 15 1 15 3 13 2
5 9 11 11 2 11
5 11 13 9 1 9
6 0 11 2 11 2 2
11 1 0 9 15 1 9 13 12 9 11 2
26 13 15 1 12 5 3 16 12 9 2 15 11 2 0 0 2 9 2 2 13 1 0 9 0 9 2
16 1 0 11 13 1 10 9 0 9 11 1 9 1 0 9 2
13 11 2 15 15 9 13 2 4 13 1 12 9 2
12 3 13 13 9 9 11 1 11 0 16 3 2
7 9 15 14 13 9 1 9
13 15 13 9 1 9 2 13 9 9 9 11 2 11
5 11 2 11 2 2
30 0 9 1 9 2 1 15 13 0 9 13 1 9 2 13 1 9 11 11 2 11 2 1 9 9 9 9 11 11 2
23 10 9 3 2 13 1 9 9 0 0 9 2 16 4 15 9 9 9 13 16 0 9 2
13 9 14 1 15 13 14 9 9 1 9 0 9 2
17 11 11 15 13 2 16 9 1 3 0 7 0 9 15 13 13 2
37 1 9 2 3 1 9 13 9 9 9 1 0 9 2 13 3 0 1 10 0 9 2 2 11 13 1 0 9 1 0 2 16 4 1 9 13 2
15 1 9 9 7 9 1 9 3 13 2 13 15 7 11 2
19 13 1 15 7 14 13 2 16 4 1 10 9 13 7 13 1 0 9 2
11 9 11 15 1 11 3 13 9 1 9 2
29 9 0 9 1 9 9 2 9 7 9 1 9 9 13 0 9 0 0 9 2 15 15 9 3 13 2 13 11 2
30 0 9 2 16 1 0 9 13 1 9 12 9 2 13 0 2 13 15 1 0 9 9 11 11 1 0 9 0 9 2
14 1 12 2 12 2 13 12 9 1 0 9 7 9 2
7 1 9 9 13 12 9 2
24 12 9 13 9 1 9 2 3 9 1 0 9 2 2 1 9 9 7 13 1 0 9 9 2
4 9 15 3 13
7 11 2 9 11 11 2 2
19 0 9 9 11 9 11 11 2 10 0 2 0 0 9 4 13 9 11 2
10 13 2 16 13 1 9 10 0 9 2
34 9 1 9 0 11 9 11 11 2 10 0 9 15 3 13 2 16 4 3 13 0 9 2 16 4 13 10 9 9 13 7 1 15 2
14 0 11 2 11 2 9 0 2 13 9 10 9 13 2
26 9 2 16 7 0 9 7 9 1 0 9 13 14 3 13 2 7 7 13 2 13 9 0 0 9 2
31 9 11 11 11 2 9 9 0 11 2 9 2 16 0 9 0 1 9 13 4 13 2 13 1 0 9 10 9 1 9 2
18 13 1 9 13 0 9 10 0 9 2 16 4 15 13 10 0 9 2
9 0 9 1 11 11 4 13 3 0
5 11 2 11 2 2
19 0 9 1 0 0 9 9 9 11 11 13 13 3 9 2 15 15 13 2
22 7 1 10 9 4 9 9 13 1 9 0 0 9 2 16 0 13 9 1 0 9 2
12 13 15 3 11 9 0 9 9 9 11 11 2
18 9 9 11 13 1 15 1 9 13 1 9 0 9 1 12 2 9 2
22 13 0 9 13 1 11 2 15 13 0 9 11 2 3 0 9 0 9 1 0 11 2
47 9 0 9 11 11 2 15 11 1 12 9 13 2 1 9 1 9 13 2 16 13 9 9 0 9 2 3 11 13 2 16 4 1 9 13 2 7 3 16 13 1 10 9 13 9 9 2
17 9 9 13 7 1 11 2 11 3 1 9 9 2 15 13 9 2
20 11 4 13 4 13 2 16 4 13 1 9 2 3 2 16 13 0 9 9 2
19 11 3 13 2 16 13 13 0 9 2 1 9 2 16 4 11 13 11 2
11 11 13 1 9 12 11 1 12 9 9 2
21 3 1 15 13 1 0 9 7 0 9 9 11 11 11 7 10 0 9 11 11 2
11 9 13 10 2 7 9 0 4 13 13 0
5 11 2 11 2 2
20 0 9 9 2 15 13 1 0 9 3 0 9 2 13 1 9 9 9 9 2
17 3 13 9 11 2 9 15 4 13 9 9 3 14 1 0 9 2
23 15 13 2 16 4 15 1 9 13 3 2 16 4 0 9 13 10 9 1 10 0 9 2
7 10 9 4 7 13 3 2
17 1 15 9 9 13 3 1 9 9 2 1 15 13 3 0 9 2
32 9 13 9 2 16 9 15 13 3 3 1 9 9 2 7 16 13 2 13 9 0 9 2 7 15 1 15 13 0 0 9 2
13 3 1 0 9 13 1 9 1 0 9 12 9 2
11 0 9 9 3 7 13 7 1 0 9 2
19 13 3 0 9 9 7 1 9 13 0 13 7 9 0 15 1 0 9 2
29 3 1 0 0 9 2 1 11 12 2 13 3 3 1 3 12 9 9 3 9 2 1 15 9 2 9 7 9 2
12 1 9 0 0 9 13 0 9 1 12 9 2
13 9 0 9 7 13 2 16 1 9 15 9 13 2
13 9 1 9 1 9 3 13 3 1 0 0 9 2
26 1 11 7 1 0 9 2 1 15 15 15 13 13 9 2 7 13 3 0 9 0 9 1 0 9 2
15 3 14 1 0 9 9 0 13 1 12 9 0 9 3 2
13 7 1 0 9 13 3 7 3 0 9 3 12 2
4 3 1 15 13
2 0 9
2 11 11
16 3 15 13 2 1 10 9 1 10 9 13 9 1 9 9 2
20 7 3 3 13 3 9 2 1 15 4 10 9 13 9 9 1 9 1 9 2
19 7 1 10 9 13 3 13 9 2 0 9 9 2 15 3 13 9 9 2
21 7 15 15 3 13 2 16 15 13 2 16 10 9 13 1 9 2 13 15 9 2
19 1 15 2 16 9 1 9 9 13 9 3 2 3 15 13 2 7 13 2
10 13 4 15 7 9 13 3 0 9 2
4 9 1 9 2
7 1 10 0 9 13 14 2
31 16 9 1 9 9 13 2 16 15 9 13 3 1 0 9 2 13 3 1 0 9 2 16 3 13 9 2 7 13 9 2
8 9 9 7 9 7 13 15 2
18 9 13 1 0 9 1 9 3 0 9 2 16 13 15 0 1 9 2
31 9 4 7 0 13 9 3 2 9 15 13 9 1 10 9 2 16 4 15 1 0 9 1 0 9 13 9 1 0 9 2
14 9 1 9 13 2 16 15 1 15 9 0 9 13 2
8 9 0 9 7 13 3 9 2
25 15 13 1 9 3 0 1 9 2 3 13 13 1 9 0 9 9 2 0 1 15 3 10 9 2
29 3 3 10 9 13 1 9 1 9 0 9 2 14 10 9 1 9 9 2 3 0 2 13 9 10 0 0 9 2
12 9 2 0 1 9 9 2 9 13 13 9 2
11 14 7 15 4 3 1 9 13 2 2 2
8 3 1 15 13 3 1 9 2
19 16 15 13 9 2 1 0 13 15 15 2 16 16 15 1 0 13 9 2
22 13 0 15 13 10 0 9 2 15 4 13 2 16 4 13 3 9 0 2 3 0 2
5 13 15 0 9 2
18 16 15 15 10 9 1 9 9 7 1 9 13 3 3 0 2 13 2
29 13 15 3 1 10 0 9 1 10 10 9 9 2 15 15 3 4 3 13 1 9 2 1 15 15 1 15 13 2
6 11 13 1 9 9 3
2 11 2
27 0 9 15 1 9 1 11 13 1 12 9 1 9 7 13 12 9 2 15 13 1 9 14 12 0 9 2
7 13 15 3 0 0 9 2
12 1 9 15 9 13 3 1 9 1 12 9 2
18 1 9 1 0 9 15 0 0 9 13 1 0 9 3 1 12 9 2
4 0 9 0 9
2 11 2
31 9 1 0 9 1 9 7 9 0 9 13 3 1 9 11 12 9 9 2 15 13 1 12 9 3 16 1 0 9 3 2
6 9 13 12 9 9 2
10 1 0 9 15 3 13 1 12 9 2
14 9 0 9 1 0 0 7 0 9 13 12 9 9 2
18 1 0 9 15 1 11 13 1 9 1 9 12 9 1 12 9 9 2
8 9 1 11 13 12 9 9 2
1 3
19 1 0 0 9 0 9 0 2 9 4 13 9 1 9 12 9 2 9 2
9 9 1 9 13 3 7 3 0 2
14 13 15 12 9 0 9 12 9 1 0 9 12 9 2
26 0 9 1 9 0 9 1 9 11 7 11 13 0 9 2 15 3 13 11 11 1 10 9 1 11 2
6 1 9 4 13 13 9
5 11 2 11 2 2
15 0 9 1 9 11 3 13 14 14 12 9 0 9 9 2
10 3 13 1 9 1 9 1 0 9 2
21 3 13 0 9 10 0 9 3 0 7 13 1 0 9 1 9 14 1 0 9 2
11 3 1 3 0 0 9 13 9 0 9 2
34 10 0 9 13 3 0 1 9 2 7 13 3 0 13 9 0 0 9 2 0 7 0 0 9 2 13 11 0 9 9 11 11 11 2
14 1 9 12 13 1 0 9 12 9 2 3 14 12 2
24 1 0 9 9 1 12 9 13 1 9 0 9 2 0 0 9 3 1 11 2 11 3 13 2
22 0 9 9 13 3 13 7 1 11 4 3 13 0 0 9 0 1 0 9 10 9 2
17 3 1 12 2 0 9 13 10 9 3 14 12 0 7 0 9 2
18 15 13 10 0 0 9 2 1 15 4 13 0 2 13 11 2 11 2
3 9 11 13
5 11 2 11 2 2
13 9 0 9 12 1 0 0 9 11 9 13 13 2
22 9 1 9 9 2 15 12 9 13 9 9 9 11 2 15 13 0 9 11 11 11 2
13 16 4 9 4 13 2 13 4 13 1 10 9 2
13 1 0 9 10 9 3 13 2 13 11 2 11 2
20 3 13 2 4 3 0 9 1 9 1 9 13 7 0 9 1 10 9 13 2
19 0 9 15 13 0 9 15 12 0 9 2 15 13 9 9 7 0 9 2
7 10 0 9 13 3 9 2
12 9 9 0 9 1 9 3 13 7 3 13 2
17 11 2 11 3 2 13 2 16 0 0 9 11 11 11 3 13 2
15 1 0 9 13 11 9 1 0 9 0 9 1 0 11 2
17 1 12 2 9 4 13 13 9 7 10 9 4 13 2 13 11 2
9 0 9 4 9 9 13 0 9 9
25 12 1 0 9 11 13 9 9 2 1 15 13 9 13 9 1 9 1 9 1 0 7 0 9 2
22 1 3 0 9 9 12 9 1 12 9 9 1 0 9 15 4 13 10 7 0 9 2
7 0 9 1 9 0 9 13
2 11 2
13 9 11 1 0 9 13 0 9 1 9 0 9 2
10 1 9 13 3 9 0 9 3 0 2
24 3 9 9 2 3 0 9 0 0 9 1 0 9 2 13 12 9 1 0 9 1 10 9 2
19 0 9 9 11 13 1 0 9 9 3 12 9 9 7 9 12 9 9 2
14 0 9 13 2 16 4 1 0 9 13 9 7 9 2
4 9 11 13 9
5 11 2 11 2 2
27 0 9 1 0 0 9 7 11 2 0 9 0 9 2 4 13 9 10 9 2 15 13 1 11 1 9 2
7 11 15 3 13 11 11 2
20 9 15 1 10 9 13 7 0 9 1 0 9 2 13 15 7 10 0 9 2
24 16 1 9 0 0 9 13 10 0 9 1 11 0 2 1 11 13 0 9 11 1 9 9 2
39 1 9 0 0 9 1 12 9 13 11 1 11 10 9 1 10 2 3 9 1 9 1 9 9 1 11 7 11 2 15 13 3 12 9 2 9 2 13 2
15 3 0 9 13 3 1 0 9 10 9 7 11 7 11 2
19 13 7 2 3 13 11 2 11 2 3 0 2 16 13 15 1 9 11 2
4 0 9 0 9
2 11 2
21 0 9 0 9 15 1 9 9 1 0 9 7 9 2 11 2 1 0 9 13 2
27 1 0 9 1 10 9 11 13 2 16 9 0 0 9 13 12 9 7 1 0 9 15 13 1 12 9 2
18 1 9 0 9 11 13 3 9 2 9 7 3 7 0 9 0 9 2
7 9 9 15 7 3 13 2
13 1 0 7 0 9 13 11 11 0 0 9 9 2
21 1 0 9 9 13 1 0 9 13 9 9 12 9 2 1 0 0 9 12 9 2
19 1 3 0 9 4 15 13 9 13 1 0 12 1 12 9 1 9 12 2
18 16 0 9 3 13 1 12 9 2 1 0 9 11 3 13 0 9 2
26 1 10 9 3 13 11 9 0 9 1 12 9 7 1 9 12 9 3 1 12 9 2 13 9 11 2
4 11 13 0 9
2 11 2
23 1 12 9 13 1 12 2 9 0 7 0 9 0 9 0 2 0 2 0 7 0 9 2
9 9 0 9 13 1 12 0 9 2
11 9 9 15 3 13 1 12 7 12 5 2
7 13 15 1 0 9 11 2
27 0 0 9 4 11 13 1 0 9 12 5 2 0 1 12 5 2 0 1 12 5 7 0 1 12 5 2
7 0 9 13 1 12 9 2
18 0 0 9 11 13 1 12 9 2 13 13 12 0 0 9 0 9 2
5 0 9 1 0 9
3 0 9 2
29 3 0 0 2 0 9 0 9 0 9 15 0 9 13 13 1 3 0 9 0 9 2 1 0 9 1 0 9 2
10 9 0 9 13 9 11 1 0 11 2
11 1 0 9 15 9 9 13 12 9 9 2
26 1 10 12 9 2 12 9 9 2 13 9 0 9 0 9 2 1 0 12 9 1 9 0 0 9 2
17 0 9 13 0 9 9 0 9 9 11 2 15 15 13 9 9 2
9 0 9 4 13 13 1 9 0 9
12 0 13 0 9 9 1 0 3 1 12 9 2
22 9 13 0 7 1 0 0 9 0 9 7 13 3 13 1 0 9 1 9 0 9 2
19 1 0 9 9 3 13 9 9 1 0 9 0 9 9 0 9 14 3 2
4 9 11 1 11
5 11 2 11 2 2
26 0 9 1 9 0 0 9 1 9 12 7 9 9 12 13 3 0 9 11 11 1 9 11 9 11 2
14 9 2 15 13 9 9 9 12 2 13 1 12 0 2
17 1 0 9 15 13 9 9 12 2 15 13 4 13 9 9 12 2
27 1 9 3 0 9 4 13 7 3 13 1 9 12 0 0 0 9 9 9 7 12 0 0 9 9 9 2
17 4 3 13 10 3 0 0 0 9 1 0 9 12 12 0 9 2
4 0 11 9 13
2 11 2
17 0 9 2 15 1 9 3 13 0 9 1 9 1 11 2 13 2
19 0 9 13 2 16 15 3 3 13 9 1 9 2 1 15 13 10 9 2
14 1 9 1 9 0 9 9 15 3 13 0 9 11 2
26 9 3 13 9 2 15 15 13 1 9 1 9 1 9 1 9 1 9 11 14 12 9 3 1 11 2
11 1 9 4 13 0 9 12 0 11 11 2
27 10 9 11 11 2 2 12 2 15 7 1 0 9 13 13 1 9 2 3 15 0 9 13 7 13 9 2
4 11 13 11 9
2 11 2
27 9 1 9 0 9 1 3 0 0 9 11 11 13 3 1 11 9 11 7 9 1 9 11 2 11 2 2
22 1 9 9 13 1 0 9 9 9 2 9 2 0 9 2 0 9 2 9 7 9 2
22 9 15 13 7 9 0 9 7 9 1 0 9 1 0 9 2 3 13 3 9 11 2
9 0 9 13 12 9 1 0 9 2
23 0 9 3 13 1 0 9 11 3 11 2 15 13 3 1 9 11 1 0 9 1 9 2
28 16 9 9 13 11 1 1 0 15 9 0 9 3 0 9 2 0 9 0 1 9 13 1 10 9 0 9 2
4 3 1 9 12
6 9 11 1 9 1 11
2 11 2
37 0 0 9 9 9 7 9 11 11 11 1 0 9 0 9 2 0 9 2 13 9 11 1 9 9 1 0 9 7 9 11 0 12 2 9 12 2
14 9 11 13 0 9 11 11 2 16 4 3 13 9 2
7 11 13 9 9 9 1 9
5 11 2 11 2 2
39 16 0 11 13 0 9 1 9 11 7 11 2 13 1 12 2 9 1 9 9 11 1 9 2 16 4 4 1 9 0 9 13 9 1 9 9 0 9 2
16 1 9 11 15 3 1 0 9 13 9 11 1 11 11 11 2
25 1 0 9 4 7 13 0 2 16 4 0 11 1 10 9 13 10 0 9 7 0 9 9 13 2
15 1 9 0 9 7 0 9 1 9 1 11 13 0 9 2
42 11 2 11 13 1 0 9 13 15 2 3 0 13 10 9 7 9 0 9 9 9 11 2 11 2 15 3 13 1 0 11 7 1 15 0 9 1 9 10 9 13 2
33 11 2 11 2 15 15 3 13 1 9 9 11 2 11 7 9 9 11 2 11 2 13 2 16 15 1 0 9 1 10 9 13 2
12 3 15 3 13 1 9 9 11 1 9 9 2
29 9 9 2 1 15 11 13 2 16 4 13 4 13 1 0 9 2 13 3 12 1 9 10 9 1 11 2 11 2
4 9 13 0 9
9 13 9 1 9 9 0 0 9 9
24 9 15 13 3 2 1 9 9 9 2 15 15 12 2 9 12 13 3 1 11 2 13 9 2
11 9 15 13 7 0 9 3 13 1 9 2
22 1 9 1 15 13 12 9 1 12 0 9 2 12 0 9 7 12 9 1 0 9 2
11 9 13 1 9 0 9 1 9 12 9 2
24 13 1 12 1 3 0 9 0 9 2 15 13 0 0 9 11 2 11 2 11 7 0 11 2
23 1 0 0 9 3 13 0 9 3 16 0 9 2 9 13 1 0 9 7 13 0 9 2
17 16 4 1 9 13 0 9 2 1 9 0 9 13 1 0 9 2
13 0 9 4 15 13 13 1 0 9 0 0 9 2
21 9 3 16 12 9 0 9 1 9 12 9 4 1 0 9 13 1 12 9 9 2
23 11 2 15 15 10 9 13 13 2 13 13 9 9 9 7 9 2 9 0 1 9 9 2
14 10 9 3 13 9 13 1 15 0 9 16 13 9 2
13 10 0 9 4 1 15 13 9 9 3 1 9 2
18 9 1 10 9 13 0 0 9 2 15 15 3 13 1 0 9 11 2
12 9 1 9 3 0 9 4 13 1 12 9 2
29 1 0 2 15 3 13 3 1 9 2 15 9 0 0 9 11 13 1 0 9 13 12 0 9 1 0 9 9 2
34 1 0 9 2 15 13 1 0 9 2 4 1 9 13 9 1 9 12 9 12 2 15 13 3 7 3 13 0 0 9 1 9 9 2
16 9 0 9 15 13 1 9 0 9 1 9 0 7 0 9 2
16 11 11 1 0 0 9 11 13 0 9 7 13 1 0 9 2
17 13 2 16 10 9 13 13 1 0 2 16 13 9 1 0 9 2
29 16 7 13 10 9 9 1 0 0 9 1 11 2 4 13 1 0 2 7 13 9 0 0 9 1 9 12 9 2
26 3 3 0 0 9 1 12 2 9 13 9 0 9 1 0 9 1 0 0 9 2 0 9 0 9 2
31 1 9 9 9 9 11 11 2 0 9 7 0 0 9 11 13 12 0 9 2 3 1 9 2 0 1 0 7 0 9 2
9 12 1 15 3 13 7 0 9 2
15 1 15 0 0 9 13 1 0 9 12 9 1 0 9 2
30 1 9 2 3 0 9 13 0 9 1 9 0 11 2 13 1 15 2 3 4 3 13 12 9 0 0 9 0 9 2
14 9 9 3 9 0 9 1 0 9 13 2 7 13 2
3 2 11 2
10 0 9 9 11 13 1 9 9 1 11
4 11 2 11 2
24 1 9 11 1 9 0 9 1 11 3 0 9 1 10 9 0 11 13 0 9 9 11 11 2
21 13 0 2 16 4 0 9 13 10 0 9 2 13 11 1 11 0 9 11 11 2
33 0 9 9 13 1 11 1 11 2 3 1 9 1 0 9 11 2 11 3 13 9 0 9 0 9 1 0 9 2 15 13 11 2
16 0 9 13 15 9 1 0 11 1 10 9 0 9 1 11 2
31 1 11 2 15 0 9 13 3 1 11 2 11 13 1 0 9 10 9 11 1 11 2 9 1 0 9 9 1 0 11 2
22 1 0 9 3 13 1 9 11 2 3 16 13 1 9 9 1 11 7 11 7 11 2
44 1 9 0 9 9 11 11 0 9 11 11 1 9 1 11 13 2 16 11 13 1 10 9 0 9 1 11 7 0 9 2 16 4 13 14 9 1 11 2 7 7 1 9 2
8 3 1 9 1 11 1 9 12
19 0 9 11 11 2 3 2 15 13 9 9 2 15 13 4 13 1 11 2
10 1 9 15 10 9 13 0 1 9 2
4 9 11 2 11
3 0 9 9
13 11 13 2 16 4 9 13 13 0 9 7 0 9
5 11 2 11 2 2
24 9 7 9 0 9 2 0 9 7 0 9 2 4 13 1 0 9 3 13 12 9 2 9 2
15 1 0 0 9 0 9 9 1 15 13 9 9 11 11 2
21 1 10 9 15 9 0 9 13 1 9 12 1 9 1 9 1 12 2 12 9 2
18 1 12 0 9 4 15 13 3 3 13 9 0 9 1 0 0 9 2
17 1 9 15 3 1 9 11 2 11 13 12 7 12 9 2 9 2
11 1 0 9 13 9 9 13 0 9 9 2
26 1 9 1 15 13 11 11 13 9 7 9 2 16 4 0 0 9 13 0 9 13 3 1 9 12 2
23 9 9 13 1 11 10 9 13 0 9 9 1 9 2 15 13 0 3 1 0 9 9 2
23 3 11 3 13 2 13 9 1 9 1 0 9 1 0 9 3 0 9 9 0 0 9 2
14 9 7 3 1 0 9 13 7 1 9 9 0 9 2
16 15 7 4 3 13 1 3 9 2 16 10 9 4 13 3 2
40 1 0 9 0 9 9 1 0 9 7 9 1 9 0 9 1 12 9 9 1 9 13 7 3 1 9 9 13 9 11 11 2 13 1 10 9 13 0 9 2
24 16 11 3 13 2 9 1 9 9 13 10 9 7 15 1 9 3 10 9 1 10 9 13 2
29 0 9 0 0 9 15 1 9 11 11 13 7 1 0 0 9 11 7 3 7 1 0 9 1 0 9 1 9 2
3 9 0 9
2 11 11
14 0 9 9 1 0 9 1 9 12 13 3 16 3 2
58 11 11 7 11 11 3 13 1 0 9 15 2 15 4 15 1 15 13 13 1 9 0 9 2 15 13 1 2 7 3 3 13 13 9 1 0 9 2 1 9 9 2 1 9 9 7 1 9 2 15 4 13 13 0 9 0 9 2
39 13 3 1 0 2 7 3 9 9 9 11 11 13 13 1 9 9 16 0 9 2 9 0 9 1 0 0 9 4 13 1 0 9 13 1 12 0 9 2
28 9 1 9 0 9 7 9 1 0 9 4 13 1 15 13 0 1 12 9 2 0 9 9 4 15 13 13 2
24 15 2 15 0 9 13 1 0 9 2 4 13 13 2 7 13 4 15 13 7 1 9 12 2
18 13 15 3 2 16 3 1 9 12 4 0 9 13 1 3 0 9 2
26 13 3 0 2 16 4 13 0 0 9 2 1 9 15 3 9 1 9 3 13 7 9 1 0 9 2
22 13 13 1 9 2 3 0 9 1 9 13 9 9 3 3 2 16 13 1 9 9 2
38 13 2 14 15 9 1 9 11 2 1 0 9 11 11 2 1 9 1 0 9 3 13 0 9 9 0 9 1 3 0 9 2 3 10 9 3 13 2
44 13 2 14 15 3 2 16 3 1 9 0 9 13 1 0 9 9 1 3 12 9 9 3 2 1 12 0 12 9 2 2 3 3 3 13 0 9 1 11 1 10 10 9 2
22 1 10 9 13 13 0 9 0 9 11 11 11 2 16 13 0 9 13 3 9 9 2
29 13 2 16 10 9 9 3 7 1 9 0 13 2 7 15 7 1 0 0 9 2 15 10 9 13 3 9 9 2
5 0 0 9 1 9
2 11 2
45 16 15 9 0 0 9 2 7 15 3 1 0 9 2 0 7 0 0 9 2 2 3 1 0 9 2 13 1 12 2 9 1 9 9 2 13 9 14 12 1 0 9 1 9 2
9 3 15 13 9 9 9 11 11 2
27 3 4 0 9 13 3 12 9 9 2 13 7 13 2 16 1 0 9 4 9 13 7 1 9 0 9 2
21 13 2 16 9 9 7 13 2 16 4 9 9 4 13 0 9 1 0 0 9 2
22 9 9 7 0 9 13 0 9 0 9 2 10 12 9 4 13 13 9 2 13 11 2
1 3
32 0 0 9 1 9 13 1 9 0 9 1 0 11 1 11 2 16 4 15 9 1 0 9 1 11 2 11 13 0 0 9 2
22 0 0 9 2 15 4 13 9 1 9 9 2 4 3 13 1 9 1 11 1 11 2
7 1 0 9 13 12 9 2
7 9 11 15 13 12 9 2
18 1 9 10 0 9 15 12 2 9 12 13 9 0 0 9 11 11 2
7 9 0 9 13 3 10 9
5 11 2 11 2 2
30 9 0 9 4 1 9 13 4 13 16 10 0 9 2 7 13 4 7 13 10 0 9 2 7 2 0 7 0 9 2
11 13 15 1 9 0 9 9 0 0 9 2
14 1 0 9 1 9 12 13 13 9 0 9 3 9 2
29 1 0 9 2 15 13 0 9 1 9 2 13 0 2 16 4 13 0 0 9 0 9 7 0 1 15 0 9 2
20 9 4 15 7 13 13 9 0 9 1 9 1 15 2 3 4 13 9 9 2
16 10 9 13 1 9 11 3 0 16 9 9 2 0 9 3 2
37 3 11 13 11 11 1 0 9 9 9 2 11 2 2 1 9 0 9 13 1 15 3 1 0 9 0 9 2 7 2 9 7 9 2 0 9 2
20 9 9 4 7 13 3 13 0 9 1 9 9 7 9 0 9 1 10 9 2
11 15 9 7 9 4 15 3 13 0 9 2
26 11 13 2 16 4 13 1 0 9 2 7 9 9 4 13 3 2 13 1 9 9 7 0 9 13 2
30 9 1 0 9 2 15 4 10 9 13 13 2 4 15 3 13 1 9 0 9 2 15 4 15 13 0 9 1 9 2
26 1 11 4 7 9 7 9 13 13 0 9 2 16 4 13 0 9 7 0 9 0 2 15 9 13 2
21 3 13 15 3 2 1 11 7 1 11 2 10 9 13 1 11 3 7 3 0 2
8 9 13 13 1 9 9 0 9
5 11 2 11 2 2
23 9 0 0 9 13 3 3 9 2 1 9 3 9 0 9 7 3 16 3 15 0 9 2
15 9 13 2 16 3 9 0 9 7 9 13 3 1 9 2
10 9 13 1 9 3 0 9 9 9 2
18 7 16 15 13 3 16 0 0 9 2 10 9 15 10 9 3 13 2
24 1 9 13 9 1 0 12 9 3 1 9 1 12 9 2 1 15 13 9 1 9 12 9 2
23 3 0 1 9 9 13 0 2 16 3 0 9 3 0 9 2 0 9 2 9 0 9 2
18 1 0 4 13 9 12 9 2 9 9 13 12 7 9 3 12 9 2
20 0 9 9 1 11 15 13 2 7 1 9 2 15 1 12 12 9 13 9 2
8 13 15 3 1 9 1 9 2
24 1 0 9 3 0 9 13 13 9 9 12 9 1 9 2 1 9 4 3 13 13 12 9 2
6 10 9 4 7 13 2
10 9 4 15 13 13 1 3 12 9 2
24 0 9 4 15 13 3 13 1 9 1 12 9 9 0 9 9 2 9 0 9 7 9 9 2
6 0 9 13 3 9 2
24 0 9 1 0 9 13 7 9 0 0 9 1 9 2 15 15 1 11 13 13 3 1 9 2
2 9 11
5 9 1 9 1 11
5 11 2 11 2 2
23 0 9 0 9 1 12 2 7 12 2 9 13 9 0 9 9 0 9 1 9 1 11 2
18 1 0 0 9 13 7 10 0 9 7 9 0 9 0 1 0 9 2
6 9 1 15 13 3 9
6 0 11 2 11 2 2
26 14 9 9 3 13 9 13 15 13 9 1 9 2 15 1 9 9 9 1 0 11 13 0 0 9 2
15 9 1 9 11 2 15 13 14 12 9 2 13 9 3 2
18 13 15 2 16 15 9 13 13 1 10 9 2 9 9 7 13 0 2
29 13 15 1 10 9 2 3 1 0 9 9 2 0 9 3 2 2 13 9 9 9 9 11 0 2 11 11 11 2
33 13 2 16 1 9 13 9 9 2 15 9 13 12 9 1 9 2 0 9 2 0 15 3 1 9 1 12 1 12 9 1 9 2
25 9 3 13 13 9 0 9 11 2 3 15 1 9 0 9 13 0 0 9 7 13 9 1 9 2
21 3 13 11 2 11 2 9 13 10 9 3 2 7 13 1 9 9 0 9 9 2
4 9 0 13 9
2 11 2
24 0 9 13 9 9 12 9 0 9 7 9 0 0 9 1 9 9 9 1 9 1 0 9 2
30 10 9 2 15 11 13 3 1 9 2 13 3 12 1 9 9 2 9 0 9 0 9 11 11 2 15 13 9 9 2
24 9 2 15 13 4 1 0 1 9 13 2 13 9 9 0 9 9 9 0 12 9 9 9 2
8 9 1 9 9 1 11 13 13
7 11 2 11 2 11 2 2
11 3 12 12 0 9 13 3 1 9 11 2
25 13 15 9 9 2 15 15 1 0 11 13 3 1 0 9 0 9 1 9 0 9 0 9 11 2
27 3 15 1 10 9 1 0 2 0 9 13 12 3 0 9 7 0 9 13 7 1 9 16 11 7 11 2
7 9 11 11 13 12 9 2
10 13 12 9 2 12 0 2 12 0 2
12 13 15 9 7 9 2 10 9 13 1 9 2
6 3 15 3 13 3 2
3 0 9 2
11 0 0 9 15 13 1 0 9 0 9 2
6 7 9 15 13 9 2
19 13 3 3 0 0 9 9 1 0 0 9 2 15 3 1 0 9 13 2
16 10 9 2 9 0 2 7 9 4 13 3 2 13 9 11 2
7 1 0 9 15 13 9 2
13 15 0 2 3 15 7 1 0 9 13 13 11 2
8 3 15 3 1 0 9 13 2
9 14 13 2 16 11 13 3 13 2
26 1 0 9 13 1 9 13 2 15 15 13 2 7 0 9 15 3 13 2 9 13 2 9 13 0 2
20 9 13 1 9 7 9 13 0 2 13 9 2 1 9 3 2 13 0 9 2
19 0 9 2 1 15 15 13 0 11 7 11 2 15 13 7 1 9 11 2
19 3 3 3 13 0 9 7 9 1 9 13 7 11 11 1 0 9 11 2
18 1 0 7 0 9 2 1 15 9 1 11 13 2 1 0 9 13 2
14 3 7 9 11 15 13 2 16 3 9 13 3 3 2
23 16 15 0 9 13 13 2 7 15 15 3 13 2 13 1 11 13 0 9 1 9 9 2
9 1 9 7 9 15 13 13 15 2
11 9 0 9 0 11 15 3 13 0 9 2
12 1 9 9 15 10 9 13 9 2 11 11 2
22 13 15 2 16 1 9 0 9 9 1 0 9 13 13 9 1 0 9 12 9 9 2
19 13 9 0 9 2 9 2 0 9 2 9 7 9 9 2 9 0 9 2
9 9 9 13 3 3 13 0 9 2
19 9 1 0 9 2 3 13 0 11 2 15 13 1 9 0 9 13 9 2
14 9 13 2 16 15 1 9 1 11 13 12 9 9 2
3 9 11 11
13 9 1 11 11 2 11 2 11 2 2 9 0 9
21 13 4 13 9 9 13 9 1 9 0 9 14 1 9 2 7 7 1 0 9 2
20 3 10 9 9 13 2 7 0 9 9 1 0 9 9 15 13 10 9 13 2
22 3 9 1 0 0 9 1 0 9 1 10 9 13 0 2 0 7 13 3 0 9 2
26 9 9 2 7 15 3 2 15 13 2 16 9 1 9 0 7 0 4 13 4 13 3 1 9 9 2
30 3 15 13 13 2 16 4 15 16 9 1 0 9 7 9 11 1 11 13 13 1 9 9 1 10 9 9 9 11 2
19 13 15 3 0 2 16 13 13 1 0 0 9 7 13 9 3 1 15 2
33 1 0 9 15 13 13 2 16 9 4 9 10 9 13 3 13 9 0 9 2 15 4 13 10 9 2 7 13 15 1 0 9 2
35 13 15 9 9 0 9 2 15 4 9 13 2 16 4 13 10 0 9 7 3 15 13 9 1 9 2 7 13 15 13 15 3 1 15 2
3 2 11 2
5 11 13 9 1 9
3 1 0 9
5 11 2 11 2 2
17 0 9 0 9 11 11 13 9 11 1 0 9 1 0 0 9 2
26 11 1 10 9 11 11 13 1 0 0 9 0 9 2 7 13 1 9 1 0 9 2 11 7 11 2
9 3 4 13 3 1 9 0 9 2
21 9 9 13 0 0 9 7 9 1 15 2 16 0 13 9 15 1 9 0 9 2
27 9 11 3 13 0 9 9 0 9 2 13 15 3 14 7 9 0 9 2 15 13 3 1 9 10 9 2
5 9 1 11 1 9
4 11 2 11 2
36 9 0 9 1 0 9 2 0 9 9 7 1 9 1 9 15 13 1 0 9 1 11 9 9 7 0 9 11 7 11 11 11 7 11 11 2
32 3 9 11 13 2 9 9 1 0 9 9 1 9 0 9 13 1 0 9 7 13 13 2 16 1 9 9 13 10 0 9 2
27 9 1 0 9 9 13 1 9 11 13 9 7 9 1 9 0 2 9 2 10 0 9 7 12 9 13 2
27 0 9 11 13 2 16 1 9 10 9 1 11 13 10 9 3 0 9 2 7 9 15 13 13 9 3 2
5 0 9 13 0 9
26 1 0 9 11 15 13 15 2 1 10 0 9 0 1 9 7 0 9 9 15 2 15 13 10 9 2
17 9 0 1 9 7 0 11 15 1 0 9 13 3 1 12 9 2
5 3 13 1 15 2
24 0 9 15 1 0 0 9 13 3 0 9 2 0 9 2 3 0 9 7 3 9 13 9 2
29 0 1 10 9 13 15 2 16 13 9 9 1 9 2 1 0 9 13 9 3 0 9 7 13 13 1 12 9 2
12 16 4 10 9 13 1 15 2 9 3 13 2
22 13 15 15 0 2 0 7 0 2 13 9 11 11 1 9 1 9 9 7 0 9 2
21 3 9 2 15 15 13 3 0 9 2 0 9 13 2 16 3 15 13 13 9 2
22 13 10 9 2 16 1 0 9 13 1 15 15 1 0 0 9 2 13 11 2 11 2
8 0 9 3 13 1 9 15 2
10 13 3 0 2 16 13 7 10 9 2
6 10 9 13 13 15 2
10 0 9 4 13 16 0 0 0 9 2
17 1 0 9 15 3 13 1 10 0 9 2 13 9 3 0 9 2
7 1 15 15 0 9 13 2
14 9 13 9 7 1 15 0 9 15 3 14 15 13 2
3 2 11 2
9 0 9 13 3 1 0 9 7 9
5 11 2 11 2 2
21 3 0 9 15 13 0 9 2 10 9 1 0 11 7 11 15 3 13 1 11 2
21 0 0 9 0 0 9 13 9 0 9 11 11 1 0 9 10 9 1 0 9 2
11 9 9 4 13 9 0 9 9 2 11 2
31 1 1 15 2 16 9 1 9 13 1 0 9 0 2 13 9 9 13 0 9 9 9 7 0 9 13 7 13 0 9 2
12 1 15 13 0 2 0 9 7 0 0 9 2
22 9 4 10 9 13 3 3 2 13 2 14 15 2 16 10 9 13 1 0 9 0 2
43 1 9 9 0 9 13 1 11 3 9 0 9 1 11 9 11 11 2 15 3 1 0 9 7 9 0 11 11 2 16 7 1 9 0 9 2 13 3 9 1 0 9 2
6 9 3 13 10 0 9
1 9
2 11 2
14 3 9 13 9 11 1 10 0 9 7 1 15 15 2
23 13 15 1 9 9 9 1 9 0 9 0 1 9 9 1 0 9 12 9 0 12 9 2
9 9 13 3 10 9 16 15 15 2
15 10 9 2 9 2 7 9 2 9 2 13 12 9 0 2
9 1 12 9 3 9 13 15 15 2
14 1 0 9 15 13 0 9 0 9 2 12 9 2 2
18 1 15 0 9 13 9 0 2 12 9 2 7 9 2 12 9 2 2
10 9 13 9 13 1 11 0 1 9 2
8 10 0 9 13 12 9 9 2
15 9 0 9 13 12 9 9 2 9 7 9 12 9 0 2
9 3 9 13 9 0 9 1 9 2
7 13 15 0 12 9 9 2
17 0 9 9 1 9 15 13 1 0 9 11 16 1 9 0 9 2
10 1 3 0 9 13 9 3 9 9 2
28 1 9 2 15 1 3 0 9 13 3 2 13 0 3 11 11 2 12 9 2 7 11 11 2 12 9 2 2
5 13 0 9 1 11
2 11 2
30 0 0 9 2 10 9 7 0 9 13 9 9 9 0 0 9 11 11 1 10 0 9 1 9 0 0 9 11 11 2
17 11 3 1 9 9 0 9 13 1 11 9 1 0 9 0 9 2
23 1 15 4 15 13 3 13 1 9 11 11 2 9 9 11 11 7 9 9 9 11 11 2
22 0 9 13 9 3 15 0 0 2 0 9 7 13 1 0 9 9 0 9 1 11 2
5 9 13 13 0 9
14 9 1 9 15 1 9 9 13 13 2 13 11 2 11
5 11 2 11 2 2
22 9 9 2 3 13 1 0 9 9 9 2 13 0 9 2 15 13 0 9 0 9 2
30 9 3 0 9 9 11 11 2 11 2 3 13 1 9 9 0 9 11 11 2 16 9 13 3 9 13 15 0 9 2
11 13 2 16 9 13 15 1 10 9 13 2
18 3 15 13 2 15 13 13 9 9 9 7 0 9 2 13 9 11 2
23 16 15 3 13 0 9 2 3 13 15 15 3 0 1 15 2 15 15 15 3 0 13 2
20 15 3 3 13 9 0 0 9 2 16 15 0 9 13 2 13 11 2 11 2
42 9 9 1 0 9 13 7 1 15 0 15 2 16 4 3 13 0 9 2 15 13 3 3 0 1 0 9 0 9 2 16 1 9 13 0 9 2 3 1 0 9 2
8 13 9 13 2 16 15 13 2
32 13 0 15 13 1 9 7 13 3 0 13 9 0 9 3 16 15 2 15 0 9 13 1 0 9 2 13 15 11 2 11 2
14 1 15 15 13 9 2 15 4 15 13 13 9 9 2
18 9 1 9 13 0 16 1 9 9 7 1 9 2 13 11 2 11 2
16 1 10 9 3 1 15 13 9 2 15 3 3 1 9 13 2
21 16 13 9 1 0 9 2 1 0 9 2 9 7 9 13 13 9 0 0 9 2
10 1 9 7 13 1 9 13 9 9 2
13 13 4 15 7 7 4 15 15 1 9 13 13 2
16 4 4 7 13 9 2 16 13 0 9 2 13 11 2 11 2
7 9 13 9 9 11 2 11
2 11 2
28 0 9 9 13 9 1 9 0 0 9 0 9 11 11 7 13 9 0 0 9 1 11 1 9 1 9 9 2
28 9 1 0 9 0 9 13 0 9 0 9 9 2 11 2 2 16 13 0 9 1 9 0 10 9 1 0 2
37 0 9 9 13 2 13 2 4 2 14 13 3 9 1 9 2 7 13 2 16 15 13 3 0 9 2 16 0 9 13 2 7 16 0 9 13 2
27 0 9 13 9 2 16 15 13 1 9 9 7 9 9 9 9 1 9 2 16 13 15 3 1 9 9 2
8 11 2 11 13 0 9 1 9
3 1 0 9
5 11 2 11 2 2
49 9 9 11 11 1 9 13 1 9 0 0 9 11 2 11 11 11 9 9 9 2 16 13 1 0 9 2 15 13 0 9 2 7 1 9 2 16 0 9 13 9 9 7 13 0 15 7 13 2
42 11 15 13 3 1 9 1 15 2 16 9 3 13 9 0 9 11 1 9 9 0 9 0 9 1 0 9 7 3 15 13 9 9 1 9 2 16 13 3 3 0 2
28 1 11 13 1 9 9 1 9 0 9 1 9 9 0 9 2 0 9 9 2 16 3 2 0 0 0 9 2
16 11 13 2 16 0 9 13 9 2 15 15 13 3 1 9 2
18 1 10 9 15 10 9 13 1 3 0 9 14 1 0 9 2 13 2
5 9 0 9 1 11
3 1 0 9
9 11 2 11 2 11 2 11 2 2
15 1 9 1 9 9 11 4 11 13 3 1 9 1 11 2
10 13 15 3 9 0 9 11 11 11 2
10 1 15 4 13 1 9 11 0 9 2
12 1 10 0 9 4 9 13 3 3 1 11 2
21 1 11 4 0 11 13 3 1 10 0 9 0 9 7 1 11 7 11 2 11 2
19 1 11 7 11 2 11 4 13 1 0 9 2 16 15 13 15 2 13 2
32 16 1 11 13 1 9 11 3 1 11 2 11 7 11 1 0 9 9 0 9 2 1 11 7 11 13 9 1 11 7 11 2
11 1 11 1 15 13 9 9 11 2 11 2
27 9 1 11 2 11 2 11 7 11 4 13 11 1 9 9 11 2 1 10 9 13 7 1 9 1 11 2
10 1 0 9 13 9 13 1 9 3 2
12 10 0 9 15 10 9 13 2 9 11 13 2
2 0 9
5 11 2 11 2 2
14 3 13 9 1 12 9 1 0 9 1 11 1 11 2
34 1 0 9 13 0 11 2 11 2 10 9 2 0 11 2 11 2 2 0 0 9 1 9 3 3 2 16 0 13 9 7 13 9 2
7 11 2 11 2 9 13 2
22 11 2 11 2 1 9 1 9 3 13 9 2 3 15 7 15 13 1 9 1 11 2
10 9 4 13 1 0 9 9 1 9 2
6 0 9 2 11 7 11
17 16 13 13 10 9 1 0 0 9 2 1 9 1 11 13 14 13
1 9
8 11 11 2 9 9 0 0 9
50 3 15 4 1 10 0 9 13 0 9 11 1 0 9 9 7 13 4 15 3 13 9 0 11 2 3 16 0 0 9 11 11 2 15 12 2 9 12 13 3 0 0 9 2 9 12 9 2 9 2
24 9 0 9 2 9 2 3 1 9 12 13 0 9 9 0 9 0 9 0 9 1 0 9 2
22 10 0 9 13 0 0 9 1 9 0 7 0 9 0 9 1 0 9 1 9 12 2
8 13 3 9 11 1 0 9 2
23 1 9 9 0 0 9 7 0 15 0 0 9 15 13 14 0 9 9 9 1 10 9 2
30 9 0 9 7 13 1 9 12 13 1 12 9 9 1 9 12 9 2 9 7 12 9 9 1 9 12 9 2 9 2
15 13 1 15 13 3 12 9 9 2 3 14 12 9 9 2
8 9 0 9 15 1 9 13 2
14 0 9 0 9 15 13 1 9 7 3 13 9 0 2
12 9 9 7 0 9 0 9 13 9 0 9 2
18 0 9 15 3 3 1 0 9 0 9 13 1 9 13 1 9 9 2
29 3 9 0 11 13 3 1 12 9 0 7 13 0 9 1 0 0 9 1 11 2 15 13 1 10 9 0 9 2
27 13 4 15 3 13 2 16 7 0 9 16 9 0 9 9 15 3 3 13 1 9 9 0 9 0 9 2
4 13 15 3 2
25 1 9 9 7 9 9 1 12 2 12 2 12 15 14 13 0 9 11 2 11 2 11 2 11 2
8 10 9 7 13 13 0 9 2
28 14 15 3 1 0 9 13 0 9 2 10 9 4 13 9 2 7 3 15 13 9 0 0 9 1 0 9 2
20 0 9 13 1 0 9 0 7 0 9 9 2 9 0 9 7 9 0 9 2
44 3 2 1 0 9 13 9 0 9 2 7 13 0 15 13 2 16 15 3 13 13 1 0 9 2 16 15 4 13 13 1 10 9 2 1 15 13 0 9 7 0 9 3 2
22 0 9 3 13 0 9 1 0 9 2 7 3 15 3 13 1 9 9 7 0 9 2
17 16 4 1 0 9 13 1 0 0 9 2 13 13 15 10 9 2
7 1 9 3 10 9 13 2
15 3 13 2 15 3 4 9 13 2 15 0 3 13 9 2
21 1 9 11 4 13 0 9 1 0 9 2 3 3 16 9 2 0 9 16 9 2
41 13 15 2 16 0 9 1 9 15 13 13 12 12 9 9 9 1 9 7 1 9 0 9 13 13 3 0 1 9 9 0 1 9 1 9 1 9 9 7 3 2
31 16 9 13 10 9 7 13 0 7 9 9 2 3 1 9 0 9 9 7 9 2 3 13 1 0 9 13 3 9 0 2
26 10 9 13 7 13 14 1 0 9 12 9 2 9 1 0 9 7 9 12 9 2 9 1 0 9 2
42 1 10 9 13 3 0 13 0 0 9 1 0 0 7 0 9 1 0 9 12 7 12 9 2 9 2 15 13 13 0 7 0 9 7 13 1 9 9 1 0 9 2
40 3 13 2 0 0 9 13 9 9 1 9 2 13 10 9 7 9 9 2 13 0 9 0 7 0 9 2 3 9 9 2 7 3 3 13 1 9 0 9 2
24 15 4 3 13 13 3 0 9 11 1 11 1 11 1 12 9 7 3 1 11 1 12 9 2
27 9 1 15 13 13 11 2 15 1 12 9 13 12 9 0 9 11 2 0 11 11 2 1 11 1 11 2
13 3 13 9 0 9 2 7 13 9 1 0 9 2
20 7 15 13 2 3 4 13 2 3 1 0 2 13 11 1 11 0 0 9 2
48 1 0 9 13 1 9 14 12 9 2 15 15 13 13 0 0 9 2 9 0 0 9 2 11 2 0 1 9 12 1 11 7 0 9 0 7 0 9 2 11 2 0 1 11 1 9 12 2
13 12 9 13 9 9 9 1 9 0 9 1 11 2
5 3 1 0 9 2
36 1 0 9 15 12 9 1 9 1 11 13 1 0 9 2 15 13 9 9 2 9 9 7 0 9 0 9 1 9 9 0 9 1 0 9 2
19 13 15 0 9 9 9 0 1 9 3 0 9 2 15 0 0 9 13 2
11 13 2 16 3 13 3 9 1 0 9 2
3 9 4 13
5 11 2 11 2 2
29 9 3 13 0 9 1 9 0 1 9 10 9 2 13 3 9 0 9 0 9 0 9 1 11 9 2 11 11 2
17 1 11 4 9 3 13 1 9 0 9 2 1 0 7 0 9 2
11 9 15 3 13 2 16 9 13 1 9 2
14 3 3 7 13 13 2 16 1 15 13 2 13 9 2
15 1 0 9 4 1 10 9 13 9 9 1 0 9 13 2
10 3 15 3 13 3 7 14 3 3 2
12 13 3 0 13 9 9 9 1 9 0 9 2
10 11 2 11 13 3 0 9 1 9 2
16 1 0 9 9 1 11 13 3 7 9 9 1 9 7 9 2
29 9 2 11 11 15 13 2 16 3 12 9 1 11 13 13 0 9 2 1 9 1 0 9 15 3 9 13 13 2
12 0 9 13 2 16 7 10 9 13 3 0 2
3 9 1 9
5 11 2 11 2 2
20 3 1 9 3 13 0 0 9 1 0 9 0 9 9 9 1 9 0 9 2
9 0 9 1 15 13 9 0 9 2
11 1 0 4 0 9 7 9 0 9 13 2
10 0 9 13 13 15 0 9 1 9 2
5 9 13 0 9 2
13 14 1 9 9 13 2 16 9 15 1 9 13 2
15 1 12 9 2 3 13 0 9 2 1 0 9 9 13 2
17 3 13 0 9 9 9 0 9 11 11 2 0 0 9 13 9 2
10 0 9 13 3 0 9 1 0 9 2
13 1 0 9 9 13 14 0 9 1 9 1 9 2
7 1 9 11 2 11 13 9
7 11 2 11 2 11 2 2
22 1 0 9 1 9 0 9 9 11 11 13 0 9 7 9 2 13 3 9 1 9 2
11 13 15 11 0 9 0 0 9 11 11 2
26 9 9 9 0 2 9 2 11 13 0 9 9 2 16 0 9 13 9 1 9 0 9 9 0 9 2
6 9 7 3 13 0 2
23 9 4 3 13 13 2 16 4 4 1 15 13 0 9 7 0 9 4 9 13 1 9 2
16 11 11 7 9 11 11 13 9 9 0 9 1 0 11 11 2
14 10 9 11 1 15 9 9 13 2 3 7 3 13 2
13 11 1 9 0 9 13 0 9 3 1 12 9 2
10 3 15 9 3 13 2 16 4 13 2
20 1 0 9 9 0 9 13 4 9 13 9 1 9 1 12 9 7 0 9 2
17 11 11 2 4 13 1 9 10 9 0 1 9 12 1 12 9 2
19 1 9 9 2 15 13 4 3 3 13 2 4 1 9 12 13 1 9 2
16 9 11 2 11 2 15 13 9 11 2 13 1 9 9 9 2
45 9 11 2 11 1 10 9 13 9 2 16 9 13 9 0 9 2 7 13 3 2 16 16 4 9 3 13 2 13 0 13 1 15 2 16 4 4 13 9 1 9 1 9 0 2
9 0 0 9 1 11 2 11 9 9
2 0 9
2 11 2
32 0 0 9 1 11 11 7 11 11 1 9 1 0 0 9 0 0 2 9 11 11 4 13 12 2 9 1 0 9 1 11 2
8 13 4 13 3 0 12 9 2
26 1 9 2 16 15 9 11 11 13 1 9 1 0 9 11 2 11 2 13 4 15 9 7 0 9 2
26 9 11 13 3 3 13 2 7 16 15 13 2 13 4 15 9 7 12 2 9 2 13 11 2 11 2
31 11 11 13 3 1 9 1 9 9 2 15 13 1 9 1 12 2 9 1 9 1 9 1 11 1 11 1 11 1 11 2
18 0 9 9 13 1 9 9 9 0 7 9 1 9 0 9 1 9 2
11 11 2 11 13 2 16 15 15 3 13 2
15 0 2 15 1 15 13 1 0 9 2 13 10 9 11 2
32 11 11 4 1 9 1 9 9 0 9 7 0 9 3 1 0 9 13 1 0 9 9 1 9 1 9 9 7 9 0 9 2
21 0 0 1 9 1 9 1 9 7 1 0 9 9 13 11 11 1 11 1 11 2
12 15 13 11 11 1 9 1 11 13 16 0 2
1 9
15 0 0 0 9 2 0 0 9 2 13 1 11 1 11 2
12 9 9 13 3 0 0 9 7 0 9 9 2
27 1 0 9 1 9 13 11 11 2 1 0 11 9 2 1 15 1 9 2 16 15 13 9 2 13 9 2
14 15 15 13 13 1 0 9 12 9 7 9 15 13 2
11 3 9 13 9 2 15 11 11 2 13 2
3 2 11 2
5 0 9 1 11 13
1 9
2 11 11
13 9 0 0 9 1 11 15 1 0 9 3 13 2
9 1 9 1 9 0 1 0 9 2
9 3 13 4 10 9 9 7 9 2
16 3 13 9 9 2 9 2 9 2 9 2 9 7 0 9 2
10 0 9 15 10 9 3 3 14 13 2
20 13 1 15 12 9 2 0 0 9 13 4 9 1 11 13 14 1 9 9 2
36 3 9 0 9 1 0 9 4 3 10 9 1 12 5 13 0 9 2 1 9 2 16 11 13 9 10 9 1 9 7 4 9 3 13 2 2
20 0 0 9 2 15 1 0 9 3 4 13 2 13 9 0 9 9 0 9 2
15 9 9 1 12 9 1 10 9 3 3 13 10 0 9 2
18 13 15 15 7 1 0 9 9 9 0 9 1 0 9 2 11 2 2
28 0 9 9 11 11 15 3 3 13 1 9 9 2 7 2 3 13 2 1 9 13 13 14 1 0 0 9 2
14 0 0 9 7 3 3 1 9 10 9 4 3 13 2
14 3 3 2 16 15 13 13 2 15 1 15 4 13 2
24 3 13 1 9 0 9 2 9 1 0 9 11 2 11 7 11 2 13 1 9 9 3 0 2
27 13 7 13 2 16 3 9 11 7 11 1 9 9 13 3 13 0 10 0 9 1 9 1 0 9 11 2
3 0 0 9
3 9 11 11
20 9 11 13 1 9 9 2 15 4 13 13 10 0 9 7 13 0 9 9 2
44 0 9 0 9 2 12 9 9 1 9 7 9 2 3 0 9 9 1 12 9 9 7 3 9 2 16 4 2 14 9 12 0 9 3 13 2 13 4 13 3 14 1 9 2
19 13 15 2 16 9 13 1 3 0 0 7 0 9 9 9 9 10 9 2
27 9 0 9 13 4 10 9 13 1 0 9 2 16 4 15 3 13 1 15 2 16 9 9 13 7 3 2
28 1 0 0 7 0 9 7 0 9 2 15 4 13 9 2 13 9 9 9 2 16 10 0 9 4 3 13 2
27 0 13 3 9 2 10 9 0 3 7 3 2 15 13 9 9 1 0 9 9 1 10 0 9 3 3 2
9 1 0 9 15 13 1 9 3 2
47 7 9 13 10 9 1 0 9 10 9 13 1 0 9 1 9 7 9 9 9 0 0 7 3 0 9 2 3 16 15 13 2 16 0 9 13 3 0 9 7 9 9 9 7 0 9 2
42 1 9 13 0 13 16 1 0 9 9 7 3 13 7 9 2 15 4 13 3 9 9 2 15 15 7 15 13 9 3 2 16 15 13 3 0 9 16 9 1 9 2
36 9 15 13 1 0 9 2 9 0 9 9 13 9 15 7 13 1 9 9 2 16 4 1 15 16 0 3 13 7 13 15 9 0 0 9 2
26 10 0 9 4 3 13 1 9 2 16 4 13 13 2 13 13 2 7 3 13 13 2 16 3 13 2
20 13 15 9 2 15 9 13 2 7 15 15 13 2 3 13 3 9 7 0 2
21 9 15 1 10 9 13 7 13 15 3 3 1 9 9 7 9 3 0 7 0 2
56 13 0 13 2 16 10 9 3 10 9 13 7 13 10 0 9 2 15 3 13 3 9 9 16 9 7 1 9 0 9 1 0 9 0 7 0 9 3 13 3 1 15 2 15 13 9 13 2 16 1 15 2 15 13 13 2
25 9 9 2 16 3 3 7 3 2 13 10 9 1 10 9 2 16 15 0 9 0 9 13 13 2
20 0 13 2 13 2 14 15 0 9 2 0 9 2 7 0 7 0 0 9 2
15 0 9 2 15 13 1 9 0 9 2 13 3 0 9 2
3 9 1 9
1 9
2 11 11
17 1 0 9 15 3 13 13 0 9 2 15 13 9 1 15 13 2
20 13 3 9 9 2 15 13 10 9 7 13 15 3 3 0 9 16 9 0 2
17 9 9 15 3 13 13 9 0 9 3 1 0 9 1 0 9 2
26 9 9 2 15 13 0 9 7 13 9 1 9 9 2 7 3 13 10 9 2 16 4 0 9 13 2
23 10 9 7 9 9 2 15 15 13 1 0 9 7 9 2 13 0 9 7 9 13 9 2
12 13 7 0 15 1 9 13 7 1 0 9 2
21 14 1 15 2 16 9 9 15 13 2 16 4 15 15 13 7 3 3 13 9 2
24 9 13 1 9 1 9 0 1 9 9 2 13 9 10 9 7 1 9 9 13 1 9 9 2
14 1 9 2 15 13 1 9 2 15 9 9 3 13 2
17 9 2 15 15 9 0 9 13 2 3 7 13 2 15 3 13 2
20 13 15 3 13 2 16 1 9 0 0 9 10 9 13 7 9 2 14 9 2
9 0 9 15 7 3 4 13 3 2
5 0 0 9 1 9
2 11 11
18 1 9 0 0 9 13 1 0 9 1 0 0 9 0 9 3 0 2
12 3 0 9 9 7 7 1 0 10 9 13 2
31 13 14 9 1 0 9 2 7 3 13 7 1 9 7 1 11 4 1 0 9 9 1 9 0 9 13 1 0 9 3 2
18 3 0 9 15 13 12 1 0 0 9 11 11 1 10 0 9 9 2
14 9 15 7 1 10 9 13 2 0 13 3 0 9 2
12 0 9 0 9 13 7 7 3 0 0 9 2
25 15 1 9 0 9 13 14 1 0 9 1 9 9 0 9 7 0 9 0 9 11 1 9 0 2
22 13 15 2 16 1 9 4 3 9 0 9 13 2 1 0 9 11 11 2 11 11 2
13 3 15 7 13 2 16 10 9 13 1 9 0 2
11 1 0 9 3 13 0 9 0 11 11 2
21 15 9 0 9 11 13 1 10 9 3 7 3 13 7 10 9 9 0 9 13 2
20 1 10 0 9 3 11 13 3 7 0 9 1 9 0 9 1 9 0 9 2
28 13 15 3 3 2 16 11 11 13 9 0 9 2 7 3 15 3 13 2 7 0 9 2 11 11 1 11 2
11 9 1 0 9 15 13 1 10 9 0 2
18 0 9 7 13 15 2 15 13 3 9 0 9 11 11 11 3 3 2
26 3 13 3 0 2 16 11 11 13 3 3 16 1 9 9 9 1 9 7 3 9 1 10 11 12 2
14 3 4 3 13 3 3 13 10 0 9 1 9 11 2
29 1 9 1 11 15 0 9 9 11 13 0 0 9 9 11 11 2 15 13 1 9 9 1 0 9 1 9 11 2
27 0 0 9 7 13 11 11 2 7 0 9 2 7 3 13 1 9 10 9 11 7 3 3 0 11 11 2
20 16 0 3 15 13 2 7 15 13 2 16 15 10 9 13 9 2 11 11 2
40 13 15 3 2 16 10 0 9 0 3 0 9 13 1 15 14 9 0 9 7 0 9 1 10 0 9 2 7 3 0 0 9 11 2 0 9 11 11 11 2
11 1 0 12 1 0 9 1 0 0 9 2
18 13 7 13 2 12 9 2 1 15 12 0 2 11 2 11 7 11 2
42 1 9 1 15 2 16 9 0 9 13 1 9 10 0 9 13 15 9 2 13 0 9 1 9 14 3 0 9 1 0 9 2 7 7 0 0 9 1 0 9 11 2
13 7 3 2 16 3 3 15 13 9 1 11 11 2
8 11 7 11 13 13 9 1 11
2 11 2
19 1 9 9 11 1 11 13 3 1 11 0 9 11 11 7 0 9 11 2
25 1 9 0 9 9 13 2 16 12 9 4 3 13 9 1 11 1 10 9 1 11 1 9 12 2
16 13 2 16 11 4 3 13 0 9 1 10 9 2 13 11 2
17 11 13 2 16 16 4 11 3 13 2 13 0 13 10 0 9 2
13 0 9 3 13 1 9 1 0 9 1 0 11 2
11 1 0 12 9 1 15 3 13 12 9 2
5 9 9 4 13 2
20 13 13 2 16 13 1 9 9 0 9 1 0 9 1 9 10 3 0 9 2
6 0 9 13 0 0 9
2 11 2
18 1 9 9 0 9 3 13 9 12 0 0 9 0 1 9 11 12 2
9 9 3 13 1 9 1 0 9 2
9 13 15 3 9 9 9 11 11 2
24 9 2 15 15 13 3 3 2 13 0 9 1 11 2 11 2 11 2 11 2 11 7 11 2
14 1 10 9 13 9 11 12 3 1 12 0 0 9 2
28 9 9 11 13 0 9 11 11 2 0 9 9 11 11 2 9 0 9 0 2 11 9 7 0 0 9 11 2
7 9 0 9 4 9 13 2
10 9 3 4 13 2 7 3 1 9 2
5 11 13 1 0 9
2 11 2
11 11 3 13 1 10 3 0 9 1 11 2
10 13 15 1 9 0 9 9 11 11 2
12 13 9 2 16 11 13 1 0 7 0 9 2
11 13 3 0 9 2 16 4 15 15 13 2
32 16 15 1 9 13 7 11 11 7 14 2 15 13 3 14 1 15 2 13 11 7 13 2 16 11 13 1 9 10 0 9 2
27 0 9 11 11 13 1 9 9 7 0 9 2 16 4 13 1 9 15 2 15 4 13 13 11 1 9 2
15 10 9 13 11 0 0 9 1 9 9 1 9 0 9 2
27 9 9 9 11 11 11 13 0 9 1 11 1 9 2 16 1 0 9 4 11 13 0 9 9 1 11 2
9 11 13 0 9 1 9 12 9 11
3 0 9 2
32 1 9 12 11 2 15 13 0 1 0 9 12 0 0 9 1 11 1 11 11 2 3 3 13 11 0 0 9 1 9 11 2
5 13 15 0 9 2
27 10 0 9 13 9 11 11 2 15 13 11 1 0 2 0 0 9 1 9 7 9 2 0 9 11 11 2
20 9 12 0 9 0 0 9 11 2 15 15 13 1 9 1 9 2 4 13 2
10 12 9 13 3 1 0 9 9 11 2
15 1 9 1 0 9 10 0 9 3 13 9 11 7 11 2
11 0 9 13 1 9 1 0 9 0 9 2
44 3 16 12 0 9 2 15 3 13 1 0 9 12 2 9 2 13 1 9 0 9 0 15 3 9 0 9 2 3 9 1 12 9 1 9 2 0 9 2 9 7 0 9 2
4 0 14 0 9
4 11 2 11 2
33 0 9 0 11 2 1 0 0 9 1 12 9 2 15 1 0 9 13 1 9 0 0 9 1 11 2 15 13 0 2 0 9 2
23 1 0 0 0 9 0 11 15 14 13 12 9 9 2 16 1 14 15 13 14 12 9 2
13 9 0 1 12 0 9 1 10 9 13 12 9 2
20 9 1 11 13 9 0 0 9 2 3 15 1 9 13 12 2 12 9 9 2
15 0 9 13 1 0 9 11 2 3 9 9 13 12 9 2
17 9 0 11 9 10 9 13 15 2 16 15 9 13 0 9 9 2
28 9 9 0 11 15 1 9 0 9 1 9 3 1 9 3 13 7 13 1 0 9 2 15 4 13 3 3 2
9 9 9 13 9 1 9 0 9 2
26 16 1 12 2 9 0 11 9 13 2 13 11 13 3 9 1 9 9 0 1 0 2 3 0 9 2
23 9 0 11 7 0 9 13 1 9 9 2 15 13 9 9 1 0 9 11 1 9 11 2
22 0 9 0 9 11 11 2 11 3 13 2 16 9 13 0 0 9 1 9 9 11 2
17 11 0 0 9 11 4 13 0 9 1 0 9 2 0 9 11 2
21 9 11 2 1 9 1 10 0 9 2 13 1 10 9 11 2 11 12 12 9 2
15 0 9 11 2 15 4 13 2 15 1 9 13 7 13 2
5 9 2 11 2 11
1 3
9 12 9 13 3 1 9 9 11 2
17 12 1 9 13 9 9 7 0 12 3 9 0 0 9 9 11 2
17 9 1 9 9 1 11 7 11 13 9 9 9 0 9 1 11 2
17 13 15 3 9 0 9 11 1 15 2 16 1 9 9 15 13 3
46 15 0 9 2 15 13 1 9 2 3 13 11 2 16 4 15 13 13 3 10 9 2 15 13 1 11 7 15 13 13 10 9 3 13 3 2 16 11 13 0 9 1 0 0 9 2
25 12 0 0 9 0 9 1 9 1 9 13 2 16 15 10 9 1 0 9 1 0 9 11 13 2
15 13 15 3 9 0 9 1 9 9 2 11 2 1 11 2
26 0 9 9 9 1 9 11 1 9 7 9 2 15 4 1 9 13 1 11 2 15 0 9 13 13 2
14 13 15 3 0 9 9 0 9 2 11 2 11 11 2
14 9 0 0 9 3 1 0 9 13 7 13 0 9 2
8 13 15 1 11 9 0 9 2
20 3 12 9 13 1 9 1 0 9 9 1 0 9 2 0 1 0 0 9 2
4 0 9 1 11
2 11 2
15 0 0 9 1 12 2 9 13 3 0 9 11 11 11 2
22 1 9 15 11 13 13 9 0 12 9 3 1 9 2 16 13 9 1 0 0 9 2
29 10 0 0 9 9 13 2 16 0 9 9 13 0 9 3 13 3 13 3 12 2 9 2 3 13 0 9 9 2
18 11 13 1 9 9 1 9 12 2 3 13 13 0 9 11 2 11 2
3 9 0 9
2 11 11
13 1 12 9 15 13 0 9 9 1 11 7 11 2
6 1 0 9 3 9 2
12 3 2 16 9 13 14 0 9 1 0 9 2
19 13 1 9 9 9 10 9 1 11 7 11 15 13 12 9 13 1 9 2
5 11 11 3 13 2
8 11 3 13 3 13 0 9 2
28 1 0 9 0 9 7 13 0 13 15 2 16 15 3 0 9 11 11 2 3 0 11 11 0 9 0 13 2
14 9 13 3 7 3 2 3 3 15 13 16 1 9 2
13 9 1 0 9 13 1 0 9 12 9 0 9 2
9 0 16 15 13 1 10 9 3 2
10 9 15 3 13 0 9 0 9 11 2
21 7 16 1 9 0 9 13 14 1 9 2 3 15 3 3 13 0 9 0 9 2
14 9 1 10 9 13 14 1 0 9 0 2 0 9 2
43 3 3 4 15 3 13 3 12 0 9 2 15 4 13 2 16 15 3 13 9 2 16 1 10 0 9 13 9 7 16 3 15 13 2 16 15 0 3 3 13 9 9 2
22 15 15 15 3 13 2 7 1 0 9 0 9 2 15 9 3 13 2 7 1 15 2
41 13 15 2 16 9 2 16 0 9 3 3 13 1 0 9 2 15 3 13 2 16 3 13 1 15 9 13 2 7 15 15 3 4 13 2 16 15 15 13 2 2
14 3 0 9 9 9 13 1 0 9 7 1 0 9 2
10 9 0 9 1 0 9 3 3 13 2
23 3 1 15 3 13 9 3 0 2 9 10 9 0 9 2 1 15 15 13 1 9 11 2
12 9 0 2 15 2 15 15 13 2 3 3 2
26 1 9 9 1 9 11 11 7 11 11 15 13 13 2 16 15 13 2 16 15 9 9 11 3 13 2
24 13 3 2 16 4 2 14 13 2 11 15 13 13 15 9 0 0 9 2 11 2 1 11 2
27 15 0 13 13 2 16 16 16 4 13 13 2 15 15 13 4 2 7 16 13 2 16 4 11 9 13 2
21 0 13 2 16 15 0 13 14 7 1 9 0 9 11 11 2 15 13 11 11 2
26 0 0 9 15 13 13 2 16 15 11 13 2 16 3 13 11 13 0 9 7 3 15 13 13 9 2
21 0 9 10 9 13 7 10 9 9 1 15 2 16 4 11 3 13 1 11 13 2
37 1 0 9 13 0 11 1 9 11 11 2 15 3 3 13 2 16 4 11 13 13 15 0 9 2 16 4 13 11 13 2 16 15 13 9 13 2
28 0 13 2 16 1 0 9 15 11 1 9 13 2 1 3 0 9 2 1 15 0 9 13 9 1 0 9 2
25 13 2 14 15 9 15 2 16 15 1 15 3 13 9 2 13 0 2 16 10 9 13 0 13 2
17 13 15 3 3 2 9 3 13 3 2 1 0 9 7 1 11 2
2 0 9
21 1 9 1 0 9 1 0 11 15 13 0 9 7 13 1 9 9 1 12 9 2
15 13 1 9 9 7 9 15 2 15 13 4 13 1 9 2
14 3 0 9 13 9 1 0 0 9 7 13 0 9 2
15 9 0 9 13 9 2 16 9 13 13 9 1 9 9 2
20 15 1 12 9 15 7 13 1 15 2 16 9 9 13 9 10 9 0 9 2
7 11 2 11 13 1 0 11
4 11 11 2 11
19 0 9 1 9 0 11 13 3 1 11 0 9 9 0 9 11 11 11 2
15 13 1 0 9 11 2 11 1 9 9 11 1 9 11 2
30 11 2 11 2 9 1 9 1 0 11 2 13 2 16 11 13 1 0 13 9 9 1 9 2 15 13 12 2 9 2
8 13 2 15 3 3 9 13 2
13 16 4 0 11 13 13 2 15 15 1 15 13 2
23 10 9 13 13 0 9 7 9 13 3 9 2 13 11 1 9 11 9 0 9 1 9 2
15 13 15 3 1 9 11 1 0 2 0 9 1 9 9 2
4 11 13 0 9
2 11 2
28 0 9 2 15 4 13 9 1 9 9 11 1 0 0 9 2 3 13 9 0 0 9 2 11 2 11 11 2
17 1 9 9 9 13 11 11 2 9 10 0 9 7 0 9 11 2
18 9 9 9 4 13 1 10 9 13 9 0 9 11 11 2 11 11 2
9 9 9 4 13 0 9 11 11 2
22 11 15 13 13 7 10 9 2 9 0 9 11 11 2 16 4 15 13 1 9 9 2
13 1 0 11 4 1 9 13 3 9 11 11 11 2
12 11 13 9 9 9 9 9 1 12 1 12 2
7 12 9 4 13 13 9 2
4 9 11 2 11
25 1 12 9 2 12 2 9 12 2 13 0 9 11 11 1 9 9 1 0 9 0 9 11 12 2
14 1 9 9 15 13 9 0 9 7 13 0 0 9 2
11 9 0 9 13 0 0 9 7 0 11 2
14 0 9 2 0 1 12 9 3 2 13 0 9 9 2
18 13 15 7 1 9 2 7 1 9 7 13 1 9 0 9 0 9 2
6 0 9 9 13 11 2
36 1 9 12 4 13 0 0 0 9 2 0 0 9 2 15 13 13 9 13 9 1 0 9 2 13 7 13 9 2 13 9 7 13 0 9 2
31 16 15 13 2 11 15 13 7 13 9 0 9 2 1 15 13 0 9 13 0 2 0 9 2 10 9 4 13 15 9 2
23 10 9 2 15 13 3 9 2 3 9 2 7 10 0 9 0 1 9 13 1 0 9 2
21 1 9 1 11 9 15 1 0 9 1 9 12 13 0 9 0 9 0 0 9 2
11 9 9 4 13 1 0 0 0 0 9 2
33 1 0 12 9 11 9 4 13 3 0 7 3 7 15 0 9 7 9 2 4 13 0 9 12 0 9 7 0 12 0 0 9 2
10 1 0 9 11 13 9 0 0 9 2
16 15 1 15 4 13 2 1 0 4 13 9 1 0 0 9 2
13 11 15 1 11 9 13 12 1 0 9 0 9 2
25 1 9 12 2 9 13 11 13 12 0 9 0 1 9 1 9 9 11 1 0 11 1 9 12 2
27 9 9 11 7 1 9 12 13 0 9 1 11 7 9 1 9 12 13 0 9 7 13 9 10 0 9 2
10 11 7 11 15 13 1 9 0 9 2
48 11 7 11 13 1 15 9 0 9 1 0 7 0 9 2 15 13 1 9 12 15 2 16 9 11 13 0 0 9 11 1 10 9 9 7 13 9 11 1 11 2 16 4 15 13 0 9 2
13 1 9 12 15 13 2 16 1 11 13 0 9 2
14 1 9 12 15 13 1 9 1 11 1 10 0 9 2
7 13 7 1 9 0 9 2
22 9 1 9 13 3 2 16 0 0 9 13 3 1 9 12 9 1 9 2 0 9 2
15 7 1 12 9 0 0 9 13 0 9 3 1 15 9 2
4 9 1 0 9
6 9 13 9 3 1 9
7 0 9 11 1 11 11 11
33 9 3 0 9 9 13 9 9 2 9 1 0 9 13 1 9 2 9 13 9 0 9 9 7 9 11 2 12 11 13 1 9 2
6 1 0 9 0 9 2
9 9 15 7 3 3 14 15 13 2
9 1 9 3 13 1 0 9 9 2
17 1 9 1 0 9 13 9 1 0 9 0 9 1 11 3 9 2
15 14 3 0 9 9 0 9 1 0 9 10 9 3 13 2
12 3 7 13 9 13 13 9 1 0 0 9 2
11 1 0 0 9 13 9 3 1 9 9 2
17 9 9 11 1 9 12 4 3 13 9 12 9 1 12 0 9 2
25 0 3 0 9 9 13 11 11 2 15 15 1 9 12 2 1 9 12 9 2 3 13 1 9 2
14 16 4 15 15 13 2 13 0 9 7 9 11 11 2
21 1 9 1 11 4 3 13 7 3 13 13 1 9 2 16 4 15 10 9 13 2
16 14 16 16 9 9 11 9 9 13 2 4 10 0 9 13 2
14 11 11 15 3 2 7 16 1 9 2 13 1 9 2
28 1 10 9 13 3 11 11 2 15 12 1 9 0 9 2 1 15 15 13 1 9 2 13 9 1 11 11 2
12 11 3 13 1 0 0 9 2 0 0 9 2
15 1 9 11 11 15 13 2 7 4 13 2 1 0 9 2
10 13 1 0 9 11 7 13 10 9 2
19 7 15 13 9 2 7 0 9 2 0 9 2 15 13 16 0 0 9 2
17 1 9 0 9 13 14 1 9 9 3 16 12 9 1 0 9 2
8 9 10 9 4 13 11 11 2
20 0 9 13 9 11 11 2 15 0 9 0 9 13 1 10 9 13 16 9 2
15 13 15 3 1 0 9 7 3 13 1 12 9 0 9 2
21 1 10 9 1 9 9 7 3 13 7 13 3 0 9 1 9 9 9 9 11 2
18 1 12 9 4 13 7 9 13 1 9 2 16 15 13 1 0 9 2
19 9 15 1 15 13 0 0 0 9 0 0 9 2 0 11 1 11 2 2
19 0 9 15 13 14 1 9 12 2 9 15 13 7 13 15 1 9 9 2
12 11 7 13 9 13 7 13 15 14 1 9 2
19 0 9 0 9 15 3 13 14 1 9 12 2 3 15 4 9 3 13 2
17 1 0 0 9 13 1 9 3 12 9 2 1 15 12 1 11 2
11 1 12 9 15 1 9 13 1 0 9 2
14 9 13 3 1 9 2 3 4 3 13 1 0 9 2
15 16 15 7 13 9 9 13 2 13 13 0 0 0 9 2
16 1 9 13 9 1 0 9 2 7 0 9 13 1 9 13 2
6 3 15 11 13 3 2
10 9 2 9 3 13 9 1 0 9 2
8 0 0 9 15 13 12 11 2
13 1 0 9 13 1 9 14 0 2 9 11 11 2
7 1 0 9 13 12 9 2
3 15 13 2
16 0 13 9 11 2 9 2 15 13 9 1 9 1 0 9 2
8 9 11 13 1 9 0 9 2
17 10 9 2 11 11 2 15 13 9 0 9 0 9 0 0 9 2
15 1 0 2 0 7 0 9 13 9 1 11 7 1 11 2
9 1 9 1 0 9 13 12 9 2
8 0 1 15 13 16 9 9 2
16 1 9 15 1 0 9 13 1 9 9 3 9 9 11 11 2
23 1 9 13 2 16 4 9 3 13 2 0 9 2 3 4 9 13 1 9 0 9 2 2
22 1 15 3 3 13 2 16 1 9 2 15 13 0 0 9 2 15 13 14 12 3 2
15 3 13 1 0 0 9 2 3 7 1 9 2 12 9 2
8 1 12 9 9 13 0 9 2
11 7 9 9 13 3 10 9 1 15 0 2
8 9 1 9 13 14 1 0 9
7 0 9 13 1 0 11 9
4 11 11 2 11
14 1 10 0 9 1 11 0 9 11 11 15 0 13 2
10 13 9 2 13 3 13 2 13 15 2
15 13 3 10 9 1 9 2 13 15 9 9 2 15 13 2
27 7 1 9 9 7 10 3 0 9 13 13 9 2 0 9 13 3 0 2 7 1 15 15 9 3 13 2
30 1 12 9 15 0 9 1 11 13 0 0 9 2 0 9 2 9 2 9 2 9 3 2 4 1 10 9 13 2 2
4 7 13 15 2
20 1 11 15 15 0 9 13 1 0 0 9 1 9 11 2 3 1 11 2 2
40 1 11 15 13 1 0 0 9 1 9 2 1 11 15 13 1 11 7 0 9 0 12 0 9 2 3 12 9 12 2 0 2 9 2 7 13 1 0 9 2
26 3 3 13 9 0 9 2 0 9 9 9 1 9 12 13 2 16 15 9 0 9 13 3 16 3 2
21 9 9 13 2 16 0 9 13 3 0 9 2 16 15 1 15 13 0 9 9 2
13 9 0 9 4 1 0 9 13 1 9 0 9 2
13 3 13 1 0 2 0 9 2 15 13 3 11 2
22 3 12 5 9 11 2 11 13 0 9 2 15 1 11 13 14 1 9 1 9 12 2
16 12 5 0 9 13 9 2 15 1 10 9 13 3 1 11 2
14 12 5 9 13 11 1 10 9 2 3 0 9 11 2
11 1 9 9 13 12 5 9 1 0 9 2
15 3 7 9 11 7 9 11 11 13 0 9 1 9 11 2
7 3 0 9 9 13 9 2
9 1 0 9 15 13 0 12 5 2
11 1 0 9 15 1 0 9 9 13 9 2
24 12 12 0 9 13 9 9 2 3 15 7 13 1 0 0 9 7 13 0 9 1 0 9 2
7 9 1 9 9 13 0 2
20 1 0 9 10 9 15 9 13 2 9 13 1 9 0 9 3 9 9 3 2
9 13 15 7 1 0 9 0 9 2
14 0 9 2 1 11 3 0 2 13 9 9 0 9 2
23 3 16 0 0 9 13 7 0 0 9 0 9 7 13 15 12 9 1 9 0 0 9 2
20 9 9 13 0 2 11 13 9 2 15 15 13 7 0 9 2 7 2 2 2
9 9 14 4 13 0 9 0 9 2
17 9 1 9 13 1 0 9 7 0 15 9 1 0 9 0 9 2
23 0 9 0 9 1 11 13 0 9 12 9 2 13 9 2 15 15 9 3 1 9 13 2
11 12 9 1 9 3 13 0 9 1 11 2
26 1 9 13 9 7 3 9 9 2 3 2 15 15 13 12 9 2 7 10 9 1 0 9 9 9 2
7 13 9 9 11 1 11 2
14 0 9 13 12 9 7 13 15 0 9 9 0 9 2
28 15 2 16 15 1 15 3 9 2 3 0 9 13 1 15 9 10 3 0 0 9 2 13 3 0 0 9 2
9 9 13 2 16 0 9 13 0 2
12 1 0 9 15 0 9 13 3 14 0 9 2
13 16 15 3 9 9 13 2 9 1 9 3 13 2
12 1 9 13 1 0 0 9 3 12 9 9 2
27 12 9 13 9 9 2 0 13 1 0 9 2 3 2 9 9 1 0 9 7 3 0 0 9 9 2 2
14 9 1 0 9 15 2 3 16 1 9 2 3 13 2
27 14 3 13 9 11 1 0 9 1 9 2 1 9 9 2 0 9 2 12 1 0 9 0 9 1 11 2
8 3 15 13 1 0 9 13 2
21 14 3 13 9 1 9 1 9 2 1 9 0 9 9 7 1 9 0 9 9 2
21 11 13 9 3 0 2 16 11 13 10 9 2 13 11 11 7 13 9 10 9 2
12 0 9 11 11 11 2 15 15 13 9 9 9
2 9 11
3 12 9 9
10 11 11 2 9 9 9 1 9 9 11
9 0 9 13 9 13 1 9 9 2
19 9 4 15 13 13 1 9 9 15 1 0 10 9 9 0 11 2 2 2
15 15 13 0 9 9 11 11 12 2 1 9 1 0 11 2
17 0 9 11 2 11 2 1 11 13 3 9 9 2 9 7 9 2
18 15 1 15 15 7 13 9 9 2 15 11 13 1 9 0 0 9 2
24 3 1 11 4 13 1 0 9 7 13 15 9 0 0 9 2 10 9 13 0 9 10 9 2
13 9 10 9 13 3 9 10 0 9 7 10 9 2
25 13 1 15 1 9 2 3 2 7 12 1 0 2 0 9 2 13 9 1 9 11 1 0 9 2
20 9 10 9 4 7 13 3 13 3 2 3 13 15 2 15 4 13 7 13 2
12 9 11 1 0 9 15 13 1 0 0 9 2
23 3 15 13 2 16 4 13 0 9 10 9 0 9 1 10 9 11 1 0 9 0 9 2
17 0 9 2 9 7 9 1 0 9 13 14 12 0 7 0 11 2
33 10 9 1 9 0 0 9 13 10 9 1 0 9 2 15 3 1 0 9 13 1 0 7 0 9 0 9 0 9 1 0 9 2
28 3 15 13 2 3 4 15 10 9 13 7 10 4 15 13 13 9 7 9 1 0 0 9 7 10 0 9 2
50 16 4 1 9 12 1 0 9 1 11 2 11 13 1 9 0 9 0 9 2 15 3 1 9 9 13 11 11 2 3 9 1 0 9 2 4 10 9 13 2 16 1 9 13 3 16 12 12 11 2
11 13 1 15 11 1 11 2 11 7 11 2
16 1 0 9 1 11 2 11 13 3 12 11 1 11 7 11 2
18 1 0 9 15 13 3 3 0 9 2 11 2 11 2 11 2 11 2
32 10 9 15 3 3 1 0 0 9 13 2 16 15 13 0 11 2 15 1 0 9 13 3 13 14 1 9 1 0 0 9 2
12 3 13 9 0 9 1 11 2 11 3 13 2
34 9 0 9 13 3 7 15 2 16 0 7 0 11 2 0 1 0 9 1 0 11 2 13 14 14 15 13 1 9 0 9 10 9 2
27 13 15 2 16 1 0 9 15 0 9 13 2 7 13 3 2 16 13 15 1 9 0 2 0 0 9 2
23 9 13 0 9 2 15 9 9 10 9 13 9 11 1 11 1 9 9 7 9 0 9 2
13 1 9 0 7 0 11 15 13 7 9 0 9 2
22 1 12 9 2 1 9 12 2 4 0 9 1 11 13 7 0 9 13 1 0 9 2
22 13 4 13 1 9 11 1 10 9 14 3 2 16 4 3 13 16 9 0 0 9 2
25 13 4 15 13 10 9 3 2 16 13 9 13 0 9 9 9 9 2 7 15 14 9 1 11 2
15 9 1 0 9 4 15 3 13 13 1 10 11 2 11 2
3 9 7 9
8 11 11 2 9 0 9 7 9
35 1 9 11 1 12 9 13 9 11 11 2 16 9 13 9 0 9 1 9 7 0 9 11 2 16 11 13 0 11 11 2 13 3 0 2
17 0 9 15 13 2 15 15 13 13 10 9 7 9 1 12 9 2
32 1 9 2 15 9 13 1 9 11 2 13 3 13 9 7 13 15 1 9 9 0 9 7 0 9 1 9 9 0 1 9 2
15 15 0 9 1 9 0 9 1 9 15 7 13 0 9 2
33 1 9 0 15 0 9 1 9 3 13 1 10 9 2 7 1 9 9 0 3 1 9 9 2 3 1 9 2 1 9 0 11 2
32 1 9 2 15 13 3 3 0 9 2 1 0 0 9 2 15 11 13 1 9 1 0 9 3 0 2 7 3 13 9 0 2
12 9 3 13 14 0 9 2 15 9 15 13 2
13 4 13 3 0 9 2 7 2 9 9 7 9 2
44 0 2 9 0 9 0 1 9 12 1 9 11 13 0 9 7 9 16 3 0 11 2 13 3 9 2 13 9 0 2 14 0 2 9 7 13 1 0 2 14 0 2 9 2
26 9 0 7 0 9 15 13 7 1 0 9 2 3 13 14 9 11 7 9 2 15 15 0 13 15 2
13 1 10 9 3 13 7 11 11 15 3 3 13 2
56 9 1 9 9 15 0 2 9 13 2 15 15 13 2 4 3 13 13 1 9 2 7 1 0 9 0 9 2 3 3 13 1 9 0 9 0 9 2 0 16 14 0 9 1 0 9 2 15 15 13 1 10 9 3 13 2
18 0 9 2 16 9 1 9 0 9 13 9 9 2 3 13 10 9 2
25 9 1 9 10 9 13 3 15 2 15 9 0 9 1 9 13 9 10 9 12 1 10 0 9 2
9 9 7 9 13 3 9 1 9 2
44 9 9 13 3 1 10 0 9 0 9 2 3 1 0 2 0 9 2 1 0 9 9 12 2 3 9 10 0 9 2 1 0 9 2 3 2 11 7 11 2 13 0 9 2
13 0 9 15 10 9 7 9 13 3 1 10 9 2
28 9 13 9 0 9 1 10 0 9 1 9 7 13 15 9 9 2 9 0 9 1 0 9 7 9 0 9 2
6 3 15 10 9 13 2
30 1 9 0 9 2 15 13 10 9 2 15 4 15 4 3 13 1 11 2 2 2 2 16 4 1 10 9 13 0 2
13 13 15 3 13 11 2 15 4 3 13 1 11 2
5 1 11 12 9 13
5 11 11 2 0 9
25 0 9 11 3 1 9 9 13 0 9 10 0 9 1 9 2 1 9 2 1 9 2 1 9 2
32 1 9 4 13 2 3 10 9 13 2 3 9 9 2 3 13 4 0 1 0 0 9 3 13 1 0 2 16 3 0 9 2
29 13 3 9 2 7 1 15 0 9 1 10 9 2 2 16 9 0 9 1 9 7 1 9 0 9 13 3 3 2
26 0 3 13 2 16 0 9 9 4 13 0 2 16 4 0 9 13 9 9 7 9 1 0 9 3 2
59 1 15 7 3 13 9 2 13 0 9 2 7 9 12 0 0 9 7 7 0 0 0 9 2 1 10 9 7 1 10 9 0 9 3 3 13 14 0 9 2 3 9 9 11 7 11 2 2 7 7 0 9 7 9 1 3 0 9 2
38 0 9 2 3 15 1 9 3 13 9 0 2 15 13 7 1 9 9 0 9 13 2 14 3 2 0 9 9 7 9 13 3 0 16 9 1 9 2
30 3 3 9 3 1 9 13 0 7 0 9 2 3 9 9 2 3 0 9 13 13 0 9 9 9 2 10 9 13 2
41 3 2 16 4 13 13 1 9 0 9 2 9 2 16 3 2 13 2 9 13 2 9 13 7 9 0 0 7 3 0 9 1 9 13 0 9 1 0 0 9 2
4 7 1 9 2
4 10 9 13 9
8 11 11 2 9 0 9 1 11
59 1 0 9 13 1 9 0 0 9 7 0 0 9 2 15 4 13 3 1 0 9 2 0 12 0 9 2 15 13 9 2 9 7 9 2 1 11 2 11 2 0 11 2 11 2 11 2 11 7 11 2 7 0 9 1 11 1 11 2
7 10 9 13 10 9 9 2
11 1 0 9 13 1 9 0 7 0 9 2
15 9 15 1 9 12 13 10 0 9 2 15 13 1 9 2
26 15 7 13 1 0 9 0 9 2 0 2 1 9 0 9 2 0 0 9 7 3 0 9 0 9 2
15 3 9 0 9 13 7 1 15 9 15 13 13 10 9 2
9 13 15 7 1 15 3 0 9 2
30 9 9 15 1 10 9 1 10 9 13 12 9 2 0 9 13 7 9 0 9 13 9 2 7 15 1 9 9 9 2
18 9 9 9 1 9 0 9 9 3 9 1 9 1 11 13 7 0 2
45 7 3 11 2 7 7 11 2 11 7 0 9 15 3 13 1 9 15 2 15 4 3 13 7 15 15 1 10 9 13 2 1 0 0 9 3 0 9 1 0 9 1 0 9 2
14 9 9 15 13 2 16 13 1 9 1 10 9 13 2
12 9 3 13 7 3 1 9 13 0 0 9 2
25 14 1 0 9 1 11 13 2 16 9 9 1 9 12 13 12 12 2 1 9 12 3 12 12 2
16 0 9 15 3 13 3 1 12 9 7 9 9 13 7 3 2
30 1 9 12 2 12 13 0 13 0 0 9 2 16 15 0 2 0 0 9 2 7 1 9 0 9 2 13 3 13 2
20 10 9 3 13 14 1 12 9 11 2 9 13 9 1 0 11 7 1 9 2
20 9 9 9 7 9 1 0 9 9 1 9 9 13 3 1 0 9 9 9 2
19 15 2 15 13 0 1 9 2 13 2 16 0 9 13 3 0 7 0 2
15 13 7 3 2 16 1 15 1 10 9 3 4 13 9 2
35 15 13 1 9 3 0 9 2 15 4 10 9 13 1 0 9 2 7 1 9 0 0 9 2 1 15 13 9 0 9 7 0 9 3 2
17 1 0 9 13 3 0 7 0 9 3 0 1 0 7 0 9 2
18 1 15 7 0 9 7 9 1 0 9 13 12 7 12 9 0 9 2
4 15 13 9 2
51 1 9 12 7 12 9 13 10 9 0 9 1 9 9 2 15 4 13 1 0 9 9 10 3 3 0 9 1 9 0 9 0 9 9 2 9 3 3 13 12 2 12 9 9 2 13 9 7 3 2 2
11 10 9 9 13 9 1 9 3 0 9 2
17 9 9 9 13 1 10 9 13 9 10 9 7 0 9 9 0 2
14 9 13 3 0 2 9 15 0 7 0 3 3 0 2
23 3 0 9 9 0 9 2 12 1 0 1 10 9 2 13 1 0 9 12 7 12 9 2
22 1 9 9 7 1 9 13 0 9 0 9 16 0 9 13 13 0 9 3 0 9 2
61 13 2 16 3 16 9 9 2 15 3 10 0 0 9 13 2 7 0 9 9 2 3 9 13 2 13 9 2 16 4 13 9 0 1 9 12 7 12 9 7 0 9 1 0 9 2 16 9 0 9 13 13 1 9 7 1 0 9 7 9 2
16 1 9 9 7 4 1 9 9 1 0 9 13 9 0 9 2
5 13 14 9 7 9
8 11 11 2 9 9 9 0 11
15 1 9 2 1 9 12 2 13 0 9 0 9 0 9 2
19 13 15 1 15 2 10 9 15 13 1 9 7 9 1 9 0 0 9 2
28 13 15 1 0 9 2 1 11 2 1 9 0 9 2 7 15 2 15 15 13 1 0 11 2 3 13 9 2
41 1 9 12 10 9 2 11 7 14 1 12 12 11 2 10 9 3 15 13 2 13 3 0 9 1 9 9 1 0 9 7 13 1 10 0 9 2 3 1 11 2
13 13 15 14 9 2 15 13 10 9 3 7 9 2
8 0 9 1 9 13 11 11 2
34 12 2 9 12 13 0 9 1 11 2 1 12 9 3 4 13 0 0 9 7 3 3 13 1 11 11 1 10 9 2 13 0 9 2
40 0 0 9 13 3 3 2 0 0 9 11 11 2 11 1 9 12 13 0 9 1 10 9 7 13 7 9 1 9 0 0 9 2 10 9 13 14 3 0 2
18 0 0 9 1 11 2 11 15 3 13 13 11 0 9 9 0 9 2
16 13 13 1 9 11 1 0 11 2 15 11 13 1 9 12 2
28 15 15 13 13 9 1 9 11 1 0 9 2 16 15 13 3 1 0 9 2 3 1 0 9 1 9 11 2
19 13 15 0 2 3 7 0 2 16 4 13 10 11 2 13 11 15 0 2
6 1 9 4 11 13 2
22 10 9 1 11 15 13 13 1 11 2 3 13 0 7 0 9 0 11 7 0 9 2
17 0 9 12 12 12 0 9 2 11 7 11 2 15 15 7 13 2
7 3 15 13 7 0 9 2
36 1 9 13 3 13 7 9 0 11 2 10 9 15 1 0 9 3 13 2 1 11 13 0 9 2 13 0 9 2 13 15 15 0 9 2 2
35 1 0 9 15 3 15 13 9 0 15 3 0 9 7 9 2 0 0 9 2 15 13 0 9 1 11 2 15 13 11 1 12 9 9 2
15 13 15 0 9 2 15 1 12 9 13 3 1 0 9 2
45 13 9 10 9 2 13 15 13 2 16 4 13 2 14 3 2 16 3 1 9 13 7 1 15 2 3 1 11 2 7 10 0 9 2 9 2 9 2 9 2 9 2 0 9 2
20 13 2 14 15 3 7 13 1 0 0 9 12 2 13 15 14 9 1 9 2
7 15 15 13 9 13 9 3
2 11 11
3 9 9 9
17 9 13 9 2 13 15 9 2 3 9 13 3 2 16 13 0 2
12 9 13 1 0 3 2 3 7 13 2 13 2
15 3 0 4 13 2 16 4 9 1 0 9 13 2 2 2
8 9 13 3 3 9 9 9 2
48 2 9 1 9 13 15 9 1 9 2 15 13 0 9 11 1 9 1 0 0 9 2 11 12 2 0 9 13 0 9 1 0 9 2 0 9 2 0 9 2 7 1 9 15 13 0 9 2
17 9 1 9 1 9 3 13 7 9 15 13 2 13 1 15 9 2
15 0 9 3 13 1 9 1 9 0 9 7 13 1 15 2
10 9 1 9 13 9 0 9 2 9 2
14 13 2 14 9 0 2 0 2 9 2 13 15 9 2
18 1 9 0 9 15 1 9 1 9 13 13 9 0 1 0 9 9 2
35 9 2 11 11 1 0 0 9 1 9 0 9 2 15 15 13 9 1 9 9 2 13 2 16 9 13 3 9 1 9 2 1 15 13 2
10 13 15 13 9 2 9 7 3 9 2
9 15 10 9 13 0 9 10 9 2
8 0 9 9 4 13 0 9 2
2 0 9
15 0 9 2 1 15 15 9 13 2 13 9 7 0 9 2
55 9 13 3 0 9 2 15 0 3 1 9 2 0 15 3 13 3 2 9 9 1 9 2 9 1 9 2 9 2 9 9 2 9 2 9 9 2 9 0 9 7 0 9 2 9 2 9 2 9 7 0 9 1 9 2
22 0 9 13 10 0 9 2 15 15 13 13 14 1 9 7 3 13 9 7 0 9 2
8 9 9 13 3 15 0 9 2
12 9 13 9 0 1 9 7 13 0 9 0 2
13 10 9 1 9 3 13 2 16 13 1 9 0 2
34 13 1 9 2 13 15 3 1 9 9 7 9 2 1 9 2 0 9 15 13 3 0 0 9 2 7 15 13 10 3 1 9 9 2
14 3 13 0 9 2 7 7 9 10 9 13 16 9 2
24 0 9 13 1 0 9 1 0 9 2 1 15 9 0 3 9 13 9 0 2 13 11 11 2
4 9 0 7 0
7 9 15 13 13 10 9 2
24 9 2 11 11 1 0 9 0 9 13 2 16 1 9 13 9 2 1 15 4 13 9 13 2
7 1 0 15 13 3 3 2
11 3 7 13 4 9 13 0 9 1 9 2
26 9 15 13 13 16 9 9 2 0 9 2 0 9 9 2 0 9 7 7 16 0 9 3 1 9 2
15 10 0 9 13 1 0 9 2 0 13 9 9 7 9 2
12 0 9 9 1 0 9 13 3 0 9 9 2
10 0 13 2 13 2 14 15 9 9 2
21 9 11 13 2 16 4 1 10 9 4 13 0 9 9 2 9 13 0 13 3 2
15 3 0 9 13 3 9 1 9 1 0 9 0 9 0 2
10 13 15 13 0 9 0 9 1 9 2
19 10 9 7 13 10 2 13 11 11 7 13 2 13 15 1 9 0 9 2
37 13 13 12 9 9 2 0 2 0 9 2 9 2 9 2 9 7 9 2 15 15 13 13 9 9 2 7 0 2 15 13 0 13 9 1 9 2
10 10 9 13 3 0 3 1 0 9 2
7 9 13 13 9 1 9 2
32 9 0 0 9 9 13 7 9 0 9 0 9 7 13 15 3 1 9 2 1 15 9 13 2 7 1 0 9 7 10 9 2
20 13 0 13 15 7 1 9 1 9 2 1 9 9 13 13 9 7 0 9 2
14 9 13 3 0 9 7 1 0 9 15 13 3 3 2
19 13 15 13 2 16 13 2 14 9 1 0 9 9 2 13 1 9 0 2
11 0 9 3 9 13 4 2 13 11 11 2
22 7 15 7 13 9 2 16 0 9 13 13 1 3 0 9 2 15 15 4 13 9 2
10 1 9 0 9 9 13 0 9 9 2
14 3 13 2 16 15 13 15 3 2 15 13 9 0 2
18 3 7 13 13 9 3 0 2 7 3 4 13 3 0 9 9 9 2
24 13 15 2 16 1 9 13 14 12 9 9 0 2 7 3 13 9 11 2 9 13 3 9 2
12 7 7 15 13 9 1 9 9 1 9 9 2
5 14 0 9 13 9
21 0 9 9 3 13 9 2 3 13 3 2 3 13 1 0 9 2 13 11 11 2
35 13 1 0 9 2 16 13 9 2 13 2 16 13 0 9 9 1 9 2 1 15 15 13 9 2 7 9 13 0 2 16 9 3 13 2
27 13 15 7 2 16 9 4 13 9 9 2 7 13 15 1 15 2 16 9 13 0 0 9 7 0 9 2
27 16 1 9 13 1 9 1 0 9 9 2 0 0 9 15 13 9 7 13 15 2 16 9 13 0 9 2
22 16 3 13 2 13 15 2 16 15 13 13 9 9 2 7 9 13 2 13 11 11 2
3 1 9 9
24 16 9 2 15 0 9 9 13 3 2 4 13 0 9 2 0 9 13 9 9 1 0 9 2
32 3 13 0 2 16 4 9 13 2 1 10 9 13 9 0 2 1 0 9 2 3 10 9 13 2 4 9 13 3 13 3 2
13 0 13 1 15 9 0 9 2 3 9 7 9 2
15 9 4 13 0 9 0 9 2 9 4 13 13 3 0 2
10 0 13 3 0 9 2 13 11 11 2
13 0 9 13 1 15 9 2 15 15 13 2 0 2
14 13 7 13 2 16 1 0 0 9 15 4 13 0 2
25 13 2 14 15 9 1 9 2 4 9 3 3 13 7 1 9 1 9 7 9 2 13 11 11 2
23 3 3 0 9 13 9 2 10 9 1 9 13 3 10 9 1 15 2 16 9 9 13 2
11 0 9 13 0 9 2 7 0 9 13 2
12 13 3 0 9 2 7 13 1 15 0 9 2
31 10 9 0 9 15 13 2 16 15 13 2 16 15 1 0 9 13 1 0 9 2 7 3 13 11 11 2 13 15 9 2
15 1 9 13 0 9 3 9 2 3 1 9 13 3 9 2
13 13 15 13 3 9 2 3 9 2 0 0 9 2
10 9 3 13 9 1 9 9 13 3 2
4 13 3 0 9
14 9 9 13 14 1 9 2 13 1 9 0 0 9 2
26 13 0 13 0 9 9 2 1 15 1 10 0 9 13 2 13 9 2 13 0 9 2 13 11 11 2
9 9 13 13 3 0 2 1 9 2
25 13 9 1 9 1 9 13 0 2 7 1 9 13 0 0 9 2 15 9 13 0 13 0 9 2
14 1 9 13 13 10 0 9 2 9 7 0 9 9 2
18 13 15 7 0 9 1 9 2 15 13 3 1 9 2 9 2 9 2
7 0 13 0 9 0 9 2
23 9 1 9 4 13 13 0 9 1 9 0 3 12 9 11 2 9 13 1 12 9 11 2
7 0 9 13 0 16 0 2
10 9 4 15 13 13 9 3 0 9 2
15 9 1 9 13 13 3 0 9 0 9 7 0 9 9 2
15 0 7 0 9 0 9 13 9 7 3 15 1 15 13 2
9 1 9 9 4 15 13 3 13 2
5 9 13 9 1 9
15 1 0 9 13 11 11 9 0 1 9 1 9 0 9 2
12 13 4 2 16 3 13 10 9 0 16 0 2
6 13 3 0 2 13 2
5 15 13 1 9 2
15 1 9 0 4 13 3 16 1 10 9 10 0 9 0 2
9 9 15 3 13 2 13 11 11 2
20 10 9 3 3 13 7 9 13 0 2 16 0 9 1 9 13 12 9 11 2
13 9 13 0 9 2 16 4 4 13 10 0 9 2
21 0 13 2 16 3 0 9 13 9 9 2 3 3 2 16 10 9 13 0 9 2
21 9 2 1 15 15 9 13 2 16 4 3 13 13 9 9 2 1 9 13 4 2
6 13 15 7 3 9 2
16 9 4 1 0 9 13 2 16 1 9 9 9 1 9 13 2
11 11 11 13 1 0 13 9 3 1 9 2
9 9 9 7 0 9 15 3 13 2
16 0 9 13 2 16 4 4 13 16 1 9 2 13 11 11 2
20 1 0 9 15 13 2 16 7 1 9 0 9 13 9 7 16 3 9 13 2
16 9 9 3 13 10 9 2 7 9 13 9 7 9 0 9 2
10 3 13 14 12 7 12 9 9 9 2
16 0 9 3 1 15 13 1 9 7 13 2 15 10 9 13 2
14 3 15 13 0 15 13 1 10 9 2 13 11 11 2
5 13 1 15 9 2
6 9 3 1 9 13 2
12 9 13 9 1 15 2 15 13 10 0 9 2
22 0 1 15 15 13 2 16 9 9 15 10 9 15 13 2 3 10 0 2 0 9 2
7 9 15 13 3 9 9 2
10 13 15 2 16 13 7 1 9 0 2
10 13 15 3 1 9 7 1 12 9 2
8 0 4 13 13 12 2 9 2
16 13 2 14 9 9 2 13 0 9 2 16 10 9 13 0 2
13 1 9 15 1 9 9 0 9 13 7 9 9 2
16 9 0 9 15 13 7 1 15 2 1 10 0 9 15 13 2
10 3 9 13 1 0 1 9 1 9 2
28 1 15 4 0 9 9 13 1 9 9 2 7 3 13 11 11 2 15 15 13 3 1 0 9 0 9 0 2
10 9 13 9 11 3 1 9 0 9 2
26 13 1 9 0 9 0 9 2 15 13 2 16 3 9 13 1 3 0 11 16 1 0 9 0 11 2
24 13 15 2 16 9 13 9 0 0 9 2 16 10 0 9 2 0 15 9 2 13 1 9 2
23 7 0 0 9 7 9 9 15 3 13 1 9 0 9 2 13 9 7 13 0 9 9 2
13 7 7 13 1 0 9 0 9 11 7 0 11 2
13 15 15 13 9 13 9 3 2 13 15 11 11 2
21 12 1 0 9 2 15 9 0 9 13 2 13 9 2 0 9 2 9 2 2 2
25 15 2 15 15 0 9 10 7 10 9 13 13 0 9 7 13 0 9 2 13 15 9 1 9 2
10 2 13 15 9 1 9 2 11 12 2
3 9 0 9
26 9 9 2 11 11 7 11 11 13 1 11 9 2 15 1 10 0 9 0 9 13 2 9 0 9 2
22 13 2 16 1 10 9 13 14 9 0 2 7 3 9 9 2 9 2 9 7 9 2
16 0 9 1 9 9 13 3 3 3 14 7 0 2 7 0 2
37 13 0 2 16 9 9 2 15 15 13 10 9 2 13 1 9 9 14 9 9 7 9 1 11 2 11 2 11 2 0 1 9 3 1 9 12 2
37 7 1 15 1 11 2 11 3 0 9 0 7 0 12 2 12 1 9 12 2 12 2 1 15 15 7 3 3 13 2 16 13 0 9 2 9 2
28 1 0 9 13 3 0 9 13 9 0 9 2 7 14 3 14 15 2 15 15 2 13 2 13 0 0 9 2
32 0 9 9 9 7 13 13 15 0 2 3 13 9 10 0 9 2 1 15 15 3 13 13 2 16 13 0 9 1 10 9 2
24 7 1 0 13 2 15 13 3 0 7 0 9 1 9 0 2 16 15 13 0 2 15 13 2
37 10 9 2 15 14 13 9 9 2 1 0 9 2 3 2 2 13 3 14 9 2 15 10 9 3 13 7 15 3 9 16 0 9 7 3 13 2
22 0 7 11 9 13 0 2 1 0 9 13 9 9 7 13 3 1 0 9 12 9 2
47 13 1 15 3 10 9 2 15 15 3 13 13 2 3 13 15 9 3 0 9 7 3 9 1 0 9 2 16 4 1 15 1 0 13 15 2 15 15 14 7 14 13 1 10 0 9 2
17 16 7 9 9 1 0 9 3 13 2 3 15 13 7 10 9 2
10 13 4 13 3 1 9 0 9 0 2
23 9 13 1 9 3 0 7 3 0 9 9 7 13 1 15 13 0 9 13 13 9 9 2
20 7 13 13 2 16 15 1 15 13 0 9 2 15 4 15 3 13 14 9 2
21 9 4 3 13 0 13 3 9 2 15 4 13 0 7 0 9 1 9 0 9 2
14 3 15 13 0 2 0 7 0 9 1 11 7 11 2
20 3 15 13 3 9 11 1 9 9 0 9 1 9 12 1 9 9 0 9 2
58 0 9 0 9 1 9 2 9 7 3 9 9 0 9 2 9 9 1 9 9 2 10 15 15 13 2 16 7 0 0 7 11 0 9 3 13 2 0 9 9 13 1 9 2 16 4 15 0 9 13 2 16 4 15 1 15 13 2
8 7 16 15 15 13 2 2 2
10 9 9 13 7 0 9 1 0 9 2
26 13 2 16 3 1 10 0 9 3 9 13 9 3 10 0 9 3 1 9 9 2 3 1 10 9 2
54 3 15 2 3 1 15 3 1 9 13 9 0 9 2 7 15 2 16 13 0 0 9 1 0 9 2 3 9 2 0 9 2 9 2 9 0 15 3 10 7 15 9 2 2 13 2 3 3 3 13 1 0 9 2
2 11 11
10 11 11 2 11 11 2 9 0 9 2
11 13 11 2 9 0 9 2 2 11 12 2
11 12 9 2 9 13 2 0 9 12 9 2
2 9 9
1 9
2 9 2
16 0 9 11 2 9 11 9 9 9 13 13 1 0 12 9 2
28 9 13 1 9 1 0 11 2 11 7 11 1 9 9 12 7 1 9 9 0 1 0 9 9 11 2 11 2
21 9 11 9 2 15 13 3 0 9 2 15 13 9 11 11 9 7 3 0 9 2
24 1 3 0 9 7 3 13 0 9 1 9 2 15 15 3 1 0 9 13 1 3 0 9 2
27 9 13 0 0 9 0 1 0 9 9 2 13 0 0 0 9 7 3 1 9 9 15 13 7 9 9 2
29 9 1 15 13 0 0 9 2 1 1 8 9 3 13 0 9 9 7 9 2 2 1 15 15 13 0 9 9 2
26 9 1 9 9 13 9 1 0 9 7 13 3 1 0 0 9 2 15 13 3 0 9 0 0 11 2
36 11 11 1 9 13 0 0 9 2 15 9 13 11 2 11 2 1 3 7 3 0 9 2 15 13 0 0 9 9 2 7 7 13 0 9 2
7 9 13 1 10 9 0 2
2 11 11
18 11 9 2 3 2 11 2 9 11 2 9 2 11 2 11 2 12 2
1 3
21 0 9 0 11 7 9 13 3 1 0 9 2 15 13 0 11 2 0 9 9 2
17 1 9 9 13 13 10 9 9 12 7 12 9 9 10 0 9 2
9 0 9 15 13 3 1 0 9 2
9 11 4 13 3 3 2 3 1 9
29 0 9 2 15 3 1 9 13 1 9 0 9 9 2 13 4 1 9 11 13 9 11 2 3 9 0 0 9 2
23 1 9 9 1 9 9 11 11 11 7 0 9 9 2 0 9 9 2 13 13 3 3 2
10 11 15 13 9 9 11 9 11 11 2
14 9 9 11 11 11 7 10 9 3 3 1 9 13 2
31 9 11 4 1 10 9 1 9 13 1 15 2 16 0 9 1 0 9 4 13 7 16 3 13 1 0 9 2 13 11 2
11 9 4 13 13 3 1 9 9 0 9 2
11 9 11 13 1 0 12 9 0 0 9 2
10 1 0 0 9 13 9 0 9 9 2
35 1 0 12 9 13 9 0 9 13 0 0 9 0 2 0 9 11 11 7 13 3 0 9 1 0 9 1 0 9 2 0 2 0 9 2
7 15 15 3 13 1 11 2
20 9 11 2 15 13 0 9 0 9 11 11 11 2 13 1 9 0 9 13 2
32 10 0 9 13 1 9 9 13 1 0 7 0 9 1 9 11 2 15 4 1 0 9 13 1 0 9 7 1 9 13 9 2
8 9 9 13 9 0 0 9 2
3 2 11 2
1 3
34 0 11 11 11 13 3 1 9 0 9 11 11 1 0 9 0 2 11 2 12 2 1 9 0 9 0 9 9 11 2 11 2 11 2
13 0 9 13 3 1 12 3 9 0 9 1 11 2
7 0 0 9 1 12 12 12
36 12 1 3 0 0 9 9 2 0 12 12 12 2 0 1 9 0 9 13 15 9 7 13 15 3 2 13 9 9 1 0 9 1 0 9 2
51 1 9 0 2 0 0 9 12 12 12 2 15 13 9 7 9 11 7 9 11 2 9 2 13 1 11 2 12 2 9 2 2 1 9 3 1 11 2 9 13 3 13 2 7 12 2 9 1 11 11 2
26 16 9 15 1 10 0 9 13 0 0 9 12 0 11 2 15 13 12 0 9 2 11 7 12 11 2
3 2 11 2
5 0 9 13 0 9
25 3 0 9 13 1 9 3 1 11 1 0 9 0 9 11 11 2 1 0 9 9 0 0 9 2
23 0 0 9 11 2 15 13 3 1 9 2 13 9 1 9 1 9 12 3 3 16 3 2
26 3 0 12 2 9 13 1 0 9 1 3 16 12 9 1 0 9 16 12 1 3 0 9 0 9 2
20 9 11 13 3 0 9 9 7 3 3 0 9 10 0 9 15 13 13 3 2
25 9 9 13 10 12 2 9 2 7 0 0 9 7 3 1 11 13 14 1 9 3 1 0 9 2
13 9 11 11 13 0 1 0 9 0 9 0 9 2
17 1 12 9 0 9 13 9 12 0 9 7 9 3 12 0 9 2
17 3 0 0 9 1 0 9 13 11 1 9 0 9 0 0 9 2
12 13 1 9 3 9 16 0 9 2 13 3 2
30 0 9 13 1 9 9 10 9 0 9 7 13 1 15 14 12 0 9 2 0 0 0 9 0 11 7 0 9 11 2
31 1 11 13 9 1 9 11 7 11 0 1 0 9 9 11 7 0 9 2 3 0 0 7 0 9 0 1 9 0 9 2
29 9 11 13 9 1 3 0 0 9 2 11 13 9 1 9 11 11 7 11 11 7 9 0 9 9 7 0 11 2
19 0 1 0 9 13 9 1 12 2 9 1 9 0 12 2 9 1 11 2
22 13 13 11 2 1 9 11 7 11 2 1 0 9 1 9 0 9 7 1 9 11 2
23 13 13 2 16 1 9 12 13 0 9 1 12 9 1 0 11 7 1 9 12 1 11 2
36 0 9 9 9 2 0 0 9 2 12 2 2 10 3 0 9 1 9 11 11 13 3 0 9 2 13 0 9 2 15 3 13 15 0 11 2
24 0 9 0 11 2 0 0 9 0 1 9 0 9 2 4 1 15 3 13 1 9 9 0 2
28 0 9 1 11 9 1 9 7 0 9 3 13 9 0 9 2 1 9 11 0 9 1 9 7 13 1 0 2
19 0 9 0 1 0 0 9 13 0 0 9 2 0 9 7 0 0 9 2
30 11 0 9 1 0 0 9 15 3 1 0 11 13 7 0 9 1 9 2 16 4 1 15 13 1 10 9 7 9 2
5 2 11 2 9 11
3 9 7 9
1 9
2 11 11
30 1 0 9 15 9 1 15 13 1 9 2 13 0 0 9 11 11 1 0 0 9 2 15 1 9 3 13 0 9 2
19 9 0 0 9 1 10 0 9 15 13 9 1 9 11 1 0 0 9 2
30 7 0 9 15 13 1 0 9 9 7 13 3 0 9 1 9 9 13 1 9 2 13 9 7 3 15 1 9 13 2
37 13 3 1 15 2 15 0 0 9 13 2 13 3 13 0 0 9 2 2 1 0 9 7 1 10 0 9 0 9 7 0 9 13 3 16 3 2
28 0 0 9 13 9 11 11 1 0 9 9 9 2 15 15 2 1 9 11 11 2 13 1 3 0 7 0 2
29 9 11 9 15 1 15 13 1 9 1 0 0 9 7 0 9 0 9 13 2 16 0 9 13 1 9 0 9 2
22 0 9 1 15 2 16 1 9 13 13 2 16 4 3 13 12 1 0 9 0 9 2
25 13 1 15 1 0 9 7 3 15 2 3 3 9 7 9 2 13 1 15 9 11 3 0 9 2
18 16 0 9 9 15 3 13 1 9 2 11 1 0 12 9 13 9 2
30 0 9 11 1 9 12 9 15 13 1 0 7 0 9 2 1 0 0 9 2 1 0 9 1 0 9 7 0 9 2
41 1 9 1 11 2 0 12 11 9 2 13 0 9 13 0 9 9 2 13 15 3 1 9 11 11 2 11 11 7 11 11 2 7 3 15 13 3 9 1 9 2
21 9 11 1 0 9 7 3 13 0 7 1 9 11 2 11 13 1 9 0 9 2
25 3 3 13 16 13 2 16 11 15 0 9 1 9 13 7 16 1 15 13 7 0 0 9 9 2
34 11 11 2 9 9 11 2 3 12 9 13 2 13 12 1 0 7 13 2 16 9 0 1 9 0 9 15 10 9 13 1 0 9 2
25 15 13 9 1 9 2 7 0 9 9 2 1 15 4 15 13 1 9 2 13 13 1 0 9 2
20 1 15 2 16 4 15 0 9 13 1 0 9 2 4 3 13 13 12 9 2
5 9 9 13 0 9
2 11 11
25 9 9 13 16 12 1 9 1 9 3 0 9 0 9 13 9 9 7 9 9 2 15 13 11 2
34 1 9 0 2 0 9 0 9 9 7 9 2 15 15 1 12 2 1 12 2 9 13 1 0 11 2 15 3 13 9 9 11 11 2
24 13 4 13 3 9 0 2 0 9 2 3 4 9 0 0 9 3 13 3 1 9 12 9 2
31 10 0 9 15 1 9 13 2 9 13 7 0 9 1 0 7 0 9 2 15 13 0 9 7 9 0 9 15 1 9 2
18 13 4 15 0 13 1 0 7 1 9 9 1 0 9 2 13 11 2
15 13 2 16 0 9 3 3 13 9 2 7 3 10 9 2
15 13 4 1 0 9 13 3 9 1 9 0 9 0 9 2
10 1 11 15 1 15 13 14 12 9 2
20 1 9 11 13 0 9 9 9 10 9 1 9 1 9 2 3 13 0 9 2
22 1 11 4 9 13 3 2 7 9 1 15 2 1 15 4 13 2 13 10 0 9 2
16 9 4 13 9 9 7 9 3 3 1 0 9 2 13 11 2
23 11 11 1 0 9 13 2 16 0 9 15 13 0 9 13 10 9 16 9 9 0 9 2
12 13 4 0 9 3 13 1 9 10 0 9 2
29 1 10 9 13 3 0 9 0 9 7 9 9 1 15 2 15 15 0 9 13 2 1 9 2 9 7 0 9 2
14 0 13 3 13 9 0 9 7 10 9 2 13 11 2
7 1 11 13 0 9 9 2
15 9 0 15 0 9 13 1 10 9 1 9 9 7 9 2
9 9 1 9 13 13 1 12 9 2
39 0 15 13 0 9 2 0 9 2 3 13 3 9 2 9 2 9 2 0 9 7 9 2 7 1 9 0 9 13 0 9 2 9 7 9 2 13 11 2
32 9 9 0 9 1 0 9 9 7 9 11 11 13 1 15 2 16 0 9 13 1 0 9 9 9 9 3 3 0 16 9 2
11 1 0 9 13 1 10 9 12 12 9 2
24 9 0 9 2 9 2 9 7 0 0 0 9 4 1 15 13 3 1 12 9 2 13 11 2
8 1 15 15 13 13 10 9 2
5 13 4 15 1 15
9 13 2 16 15 13 13 9 0 2
6 13 1 10 3 9 2
10 13 3 15 13 2 16 10 11 13 2
8 3 3 3 13 3 7 11 2
15 13 4 3 0 15 13 1 9 0 2 0 2 0 3 2
30 13 4 3 9 0 7 0 7 3 15 13 2 16 4 13 1 9 2 16 0 9 11 13 1 9 2 7 9 0 2
14 2 11 11 2 11 2 15 13 9 1 9 0 9 2
25 13 15 1 0 9 7 9 2 0 9 7 9 2 15 13 9 1 9 2 1 15 4 13 13 2
9 1 9 12 13 9 9 3 13 2
40 0 9 9 2 12 2 12 9 2 13 2 16 1 9 0 7 0 1 15 13 9 0 2 0 2 0 7 0 2 0 2 2 7 9 15 7 13 3 13 2
41 9 0 9 7 9 0 1 9 12 2 15 13 9 0 9 7 13 9 0 2 13 2 16 0 13 9 3 13 1 10 9 2 16 4 15 13 15 7 3 13 2
10 1 9 15 15 7 13 2 9 13 2
35 1 9 9 0 9 0 0 9 9 2 11 4 9 9 11 13 3 2 1 9 9 2 3 9 13 10 9 2 1 15 15 13 13 0 2
7 10 0 9 3 13 13 2
19 1 0 9 15 7 13 9 10 9 2 1 15 15 13 3 16 12 9 2
55 13 3 0 13 9 0 2 7 16 0 9 7 9 3 13 2 7 13 1 9 2 13 2 14 15 15 11 7 11 2 16 13 0 9 7 15 13 13 3 0 1 9 2 3 13 2 10 0 9 15 1 15 13 13 2
18 13 7 13 1 15 2 16 1 0 9 15 13 16 9 0 2 11 2
4 0 9 3 3
9 9 13 3 0 2 16 9 13 0
2 11 2
17 1 0 9 13 9 9 7 9 3 16 12 9 9 0 0 9 2
13 13 15 1 12 5 3 16 1 0 9 9 12 2
23 1 0 9 4 1 0 0 9 13 12 9 9 12 0 9 7 1 11 12 9 9 12 2
14 3 9 4 13 1 11 2 7 15 12 9 9 12 2
27 1 9 4 1 0 9 13 1 11 3 3 12 9 9 2 15 13 1 12 9 3 16 1 0 9 3 2
17 1 11 4 13 3 16 12 9 9 7 1 11 3 12 9 9 2
20 9 1 11 13 1 0 9 3 16 12 9 9 2 1 12 9 3 16 3 2
18 1 11 15 1 9 13 0 12 9 9 7 1 11 3 12 9 9 2
8 1 9 7 11 13 9 1 9
2 11 11
18 1 0 9 11 11 4 3 13 9 0 9 0 9 7 0 9 9 2
25 10 9 13 0 7 13 1 0 0 0 9 9 1 0 9 2 3 1 9 9 2 9 11 11 2
24 13 4 15 13 15 2 16 4 15 10 9 13 1 0 9 9 2 13 11 9 9 1 9 2
12 10 9 7 13 3 3 3 7 0 3 3 2
18 9 0 9 2 15 9 7 9 13 2 3 11 13 3 1 0 9 2
19 1 10 9 13 13 3 14 1 12 9 2 9 0 9 13 13 1 9 2
32 0 9 15 15 13 3 1 9 7 12 9 3 13 9 1 0 9 2 15 9 2 0 9 9 11 2 13 13 3 9 9 2
15 9 13 10 0 9 1 9 9 11 11 2 13 11 11 2
35 13 4 9 13 0 9 10 0 9 2 3 9 2 15 13 3 1 0 9 1 0 9 11 2 7 1 11 4 13 13 3 7 1 9 2
18 13 3 9 0 2 1 15 13 12 0 0 9 7 0 9 0 9 2
26 0 9 11 11 7 11 11 2 0 9 0 9 2 9 9 3 13 2 3 13 10 0 9 3 0 2
14 1 11 13 3 9 7 9 9 11 11 7 11 11 2
36 13 15 7 3 1 9 3 0 2 3 9 13 11 16 9 1 0 9 2 1 9 13 7 0 9 13 15 3 7 13 3 7 12 9 0 2
21 15 4 3 2 3 2 13 1 0 2 3 0 9 7 13 2 15 13 0 9 2
25 13 3 3 1 9 2 3 0 9 13 13 0 9 7 16 0 15 13 3 2 13 10 9 11 2
19 2 3 1 0 9 9 13 9 1 11 13 0 0 9 3 12 9 2 2
11 1 11 13 9 1 9 9 9 3 0 2
21 13 3 0 9 9 7 15 15 1 9 13 1 9 7 3 2 16 13 1 9 2
28 11 11 13 3 0 9 2 15 13 7 3 0 9 13 9 2 1 15 1 0 9 13 1 0 9 11 11 2
30 9 9 9 7 0 9 13 12 3 0 0 9 1 0 9 2 13 9 7 9 2 15 1 0 9 13 3 11 11 2
11 13 15 10 9 9 2 13 1 15 11 2
15 1 0 9 13 3 0 15 2 15 13 0 16 12 9 2
13 7 13 0 13 15 1 9 2 10 9 13 9 2
19 9 3 3 13 15 15 1 15 7 3 14 13 15 2 15 1 15 13 2
30 13 7 9 13 10 9 2 16 0 9 13 12 1 0 1 9 7 13 0 9 1 9 0 2 0 7 0 2 2 2
6 10 9 13 9 0 2
9 3 9 13 9 13 3 1 15 2
7 0 0 9 1 11 13 9
9 0 9 1 11 3 13 3 15 2
30 1 0 9 11 15 1 12 2 1 12 2 9 13 9 0 9 2 0 9 2 2 15 13 9 1 9 11 1 11 2
16 10 9 13 0 1 12 9 2 15 11 13 1 0 12 9 2
12 1 9 13 13 9 2 9 2 9 7 9 2
13 0 9 15 9 4 13 13 1 0 9 0 9 2
16 10 9 15 9 11 13 3 12 9 7 9 15 13 10 9 2
20 1 9 13 3 9 11 11 1 11 2 11 11 1 11 2 11 11 1 11 2
9 13 4 7 9 11 11 1 11 2
3 2 11 2
6 0 2 0 7 0 9
8 9 0 9 13 0 9 1 11
19 11 11 2 9 2 0 2 12 2 13 9 9 2 9 9 9 9 9 9
49 1 9 0 9 11 2 9 11 1 0 9 9 7 1 9 1 0 9 7 9 15 3 13 0 9 2 0 9 13 1 0 2 9 0 9 9 0 9 2 9 9 0 9 1 9 12 2 12 2
16 9 0 11 13 0 9 9 0 9 7 9 1 3 0 9 2
17 3 7 9 13 0 9 0 9 9 1 0 9 9 9 11 12 2
17 0 9 2 3 0 9 1 10 9 9 2 15 3 3 13 3 2
15 1 9 9 11 11 1 9 11 11 1 9 9 11 11 2
15 3 13 1 9 9 11 2 11 2 11 2 11 7 11 2
52 10 9 1 0 2 0 9 7 1 9 9 2 15 11 7 11 13 1 10 0 2 0 2 0 9 9 2 13 13 1 3 0 9 2 3 7 3 0 2 9 1 9 1 11 2 11 7 11 2 11 2 2
19 3 0 13 9 12 1 0 0 9 11 11 2 15 9 12 13 1 11 2
20 3 13 1 10 0 9 2 3 0 9 1 9 11 2 11 1 9 12 2 2
17 3 0 13 9 11 1 10 0 9 2 3 3 13 10 0 9 2
22 12 9 13 0 2 13 9 2 1 9 9 2 1 9 9 2 0 0 9 2 2 2
12 9 0 9 15 13 1 9 9 9 1 9 2
30 3 13 9 9 11 2 11 2 1 9 0 9 0 9 2 9 9 0 2 11 11 2 15 13 9 11 2 11 2 2
13 0 9 9 13 9 9 0 0 9 1 9 12 2
23 1 9 1 9 13 3 3 9 2 0 9 9 11 2 0 11 2 9 11 7 0 9 2
19 3 0 13 9 9 11 2 7 11 2 1 9 12 2 0 3 1 11 2
31 9 13 13 0 9 2 9 3 11 2 11 2 11 7 11 2 0 0 9 7 9 2 15 7 1 0 9 13 0 9 2
47 16 4 15 13 15 2 1 10 9 9 15 13 13 9 7 13 0 9 2 0 9 11 2 11 2 11 2 11 2 9 11 7 11 2 3 11 2 11 7 0 9 9 11 2 11 2 2
10 0 9 13 9 11 9 0 0 9 2
23 0 11 13 0 9 9 0 9 0 1 12 9 9 1 9 9 2 7 1 0 9 2 2
18 1 15 13 1 9 13 12 9 1 0 0 9 2 0 9 11 0 2
9 9 13 0 9 2 7 0 9 2
28 7 1 0 9 13 9 9 2 13 15 3 0 0 9 3 0 1 9 1 0 0 9 11 11 7 11 11 2
14 1 9 1 15 0 11 13 9 9 9 1 0 9 2
3 15 13 2
5 0 11 2 11 2
8 12 2 9 2 12 2 9 2
3 14 0 9
23 11 11 2 0 2 12 2 13 0 9 2 0 9 7 9 2 9 0 9 9 0 11 2
11 9 3 9 13 9 1 0 9 11 11 2
39 9 9 15 13 1 9 0 9 2 15 3 13 0 9 2 9 10 0 9 2 0 9 1 11 2 0 13 3 1 15 13 2 16 3 9 14 13 11 2
18 1 10 9 13 9 11 11 1 9 12 2 0 0 0 9 0 9 2
38 1 9 9 4 15 13 1 9 7 13 2 15 15 1 12 9 1 0 9 13 2 0 9 9 11 2 9 0 9 1 9 2 0 9 9 0 9 2
52 7 3 9 2 9 2 9 2 9 2 3 10 0 2 15 1 12 9 3 3 13 1 9 9 9 7 9 1 0 9 0 9 2 10 9 7 1 0 9 3 3 13 1 9 0 9 9 11 1 0 9 2
11 3 4 10 10 9 13 2 7 3 14 2
12 15 4 7 13 13 2 13 0 9 1 9 2
17 13 15 3 15 2 15 1 9 0 9 13 0 0 7 0 9 2
25 9 0 9 15 13 3 9 9 2 16 11 15 3 13 1 9 0 2 3 0 0 9 2 9 2
5 9 9 3 13 2
18 9 10 7 0 9 15 3 13 2 16 15 1 10 9 13 9 9 2
21 1 0 9 15 13 0 9 2 1 0 0 9 1 0 9 7 9 1 0 9 2
31 3 13 2 16 1 11 9 13 2 7 15 2 15 13 1 10 0 9 2 13 1 9 9 2 1 9 11 1 9 3 2
9 13 1 15 2 9 1 11 13 2
21 1 11 13 14 0 9 2 15 0 0 9 13 9 1 0 9 0 7 0 9 2
42 15 13 3 0 9 2 7 15 15 4 13 2 16 2 3 2 9 0 9 11 1 9 10 9 1 9 9 1 9 11 2 11 13 0 9 7 11 1 3 0 9 2
32 1 11 15 1 0 9 0 9 1 0 9 11 2 15 15 13 9 1 11 2 13 9 9 1 0 9 14 1 0 0 9 2
11 13 15 13 2 16 0 9 4 13 9 2
47 1 11 15 0 9 1 0 0 9 13 1 9 9 16 9 9 12 2 2 2 1 0 0 9 2 9 2 15 15 3 13 1 0 9 12 2 12 7 13 15 0 9 1 10 9 11 2
20 13 15 2 16 0 9 9 2 9 7 0 9 13 3 0 9 1 11 0 2
28 13 9 4 13 9 10 9 2 1 10 9 13 2 16 15 13 0 9 13 15 1 9 7 13 15 1 9 2
23 16 1 10 9 9 1 11 13 0 9 2 9 11 13 1 11 0 1 9 12 0 11 2
14 13 2 16 4 15 3 1 11 13 9 0 0 9 2
19 7 16 14 2 9 9 2 15 4 13 1 15 2 4 13 3 12 9 2
2 11 11
4 0 2 7 0
1 9
39 9 2 0 9 2 9 7 9 11 11 13 1 9 12 0 0 0 9 11 2 15 0 7 0 9 13 1 0 9 0 9 0 9 2 0 9 7 9 2
38 16 11 13 0 9 9 2 7 7 0 9 9 9 0 2 13 15 11 11 0 9 1 9 10 9 1 9 12 0 9 13 7 13 15 3 0 9 2
32 1 10 0 9 2 15 13 1 0 9 11 11 7 13 15 9 1 0 0 9 2 3 13 0 9 2 0 11 1 0 11 2
28 9 4 9 11 13 1 9 9 7 11 11 15 1 15 13 12 9 2 15 13 2 15 13 1 11 0 9 2
29 9 1 15 15 3 13 3 0 9 2 0 9 7 0 2 16 0 2 0 9 2 9 2 0 2 0 9 2 2
19 1 0 9 11 13 7 0 9 3 0 7 0 2 0 11 2 13 2 2
64 0 9 9 13 7 1 0 0 9 1 3 0 2 16 15 13 1 11 2 0 9 13 0 2 0 7 0 9 1 0 9 2 9 2 11 2 2 0 9 2 15 13 1 13 1 0 0 9 2 7 14 3 0 9 2 0 0 9 7 0 9 9 2 2
21 13 3 7 9 9 2 9 2 9 2 7 2 9 2 9 2 0 9 2 2 2
11 0 9 9 15 7 3 13 1 10 9 2
17 11 11 15 13 15 2 15 9 11 1 9 9 2 1 9 12 2
25 1 9 13 0 0 9 1 9 1 0 0 9 13 1 0 9 9 0 9 7 1 10 0 9 2
2 11 11
8 11 11 2 11 1 0 11 2
4 9 12 9 2
14 13 9 12 11 2 12 2 9 1 11 2 11 11 2
5 9 1 9 13 6
17 1 12 2 9 15 13 9 13 1 10 9 1 9 9 12 12 12
2 11 11
10 13 0 1 9 9 1 12 9 3 2
6 13 15 14 12 9 2
8 13 9 2 2 13 4 15 2
2 13 2
5 13 15 15 13 2
3 13 9 2
20 16 4 13 9 3 13 2 3 4 15 13 7 13 4 15 2 13 4 15 2
10 9 13 7 3 13 2 15 4 13 2
9 10 9 4 3 1 9 9 13 2
32 9 9 12 12 12 2 15 1 0 9 13 1 11 9 10 9 2 4 13 3 1 9 13 3 7 3 0 7 3 0 9 2
10 15 15 1 15 13 2 3 15 13 2
10 1 0 9 15 13 14 10 0 9 2
9 13 15 13 2 16 15 13 9 2
20 1 10 0 9 7 13 3 13 15 9 7 9 2 15 15 13 1 0 9 2
16 13 4 15 15 2 16 4 10 9 1 9 13 1 0 9 2
11 9 1 15 13 2 16 4 15 13 6 2
17 13 0 7 0 0 9 2 13 0 9 11 11 2 9 9 9 2
18 15 15 13 9 13 0 9 2 13 1 0 9 3 7 1 0 9 2
11 1 10 9 15 1 10 0 9 13 15 2
4 9 9 0 9
12 0 11 15 9 9 3 13 2 16 13 9 2
10 1 0 9 15 13 2 15 13 9 2
5 9 7 9 9 2
10 13 15 2 16 9 15 13 9 9 2
6 7 15 15 13 3 2
12 3 1 15 13 2 1 9 15 3 13 13 2
8 13 9 7 1 15 9 9 2
9 13 15 15 2 3 1 9 13 2
7 13 2 1 15 13 9 2
11 9 7 9 15 13 2 16 3 3 13 2
6 11 13 1 11 11 2
17 15 3 3 13 2 7 10 9 3 13 9 9 9 7 0 9 2
3 0 13 9
14 1 0 9 12 12 12 4 3 13 9 1 0 9 2
26 13 2 16 9 15 9 13 1 9 10 9 2 16 4 15 1 15 13 7 15 2 15 4 3 13 2
9 0 13 2 16 4 15 13 9 2
27 16 15 9 4 13 2 16 4 15 1 10 9 15 1 9 7 9 13 2 13 15 13 2 13 11 11 2
16 3 15 13 2 16 15 13 10 9 2 15 13 13 0 9 2
14 3 13 9 12 12 0 2 9 2 15 4 13 0 2
16 13 1 15 3 9 0 9 2 9 2 9 2 9 2 9 2
10 13 9 1 0 9 1 9 1 9 2
4 3 9 3 13
11 9 12 12 12 13 1 9 3 12 9 2
4 13 12 9 2
7 0 9 4 13 9 3 2
22 1 9 1 9 15 13 13 2 16 0 9 9 13 3 1 12 2 7 12 2 9 2
12 7 3 1 9 9 2 15 13 1 0 9 2
7 1 9 1 7 1 9 2
4 1 9 9 2
11 9 13 3 3 3 2 3 1 0 9 2
22 9 13 3 1 9 2 7 3 13 13 3 7 1 9 9 9 7 13 15 15 9 2
14 1 10 9 4 9 1 9 9 13 2 13 9 9 2
18 16 9 13 2 13 7 9 3 2 7 15 1 15 9 13 0 9 2
11 13 15 3 10 9 2 15 4 13 13 2
29 16 15 13 9 7 9 1 15 13 9 2 13 15 1 9 9 7 0 9 1 0 0 9 2 15 13 9 9 2
8 3 15 1 15 13 9 9 2
24 16 9 13 2 16 13 1 9 9 7 9 9 2 13 15 1 0 9 1 9 9 7 9 2
3 0 0 9
9 9 4 13 9 13 2 7 13 2
17 9 15 1 10 9 13 13 9 2 7 16 13 1 3 0 9 2
11 0 9 15 1 0 9 3 13 15 0 2
13 3 13 3 0 9 3 9 1 10 9 16 3 2
6 13 7 15 3 13 2
12 7 15 15 13 2 7 9 13 3 3 0 2
17 13 10 9 3 3 13 2 16 13 2 16 13 9 3 1 9 2
20 9 13 13 7 1 9 2 3 0 9 2 15 3 3 13 9 1 10 9 2
11 3 9 13 3 14 9 2 13 11 11 2
24 9 9 9 9 13 13 10 9 2 16 4 15 9 1 10 0 9 13 13 7 13 15 15 2
6 13 15 9 1 9 2
7 13 4 9 13 7 13 2
7 13 13 2 3 3 13 2
6 13 13 2 15 13 2
10 13 2 16 4 1 15 9 13 3 2
13 16 15 13 13 2 3 15 1 15 13 15 13 2
12 13 1 15 2 16 4 15 1 9 13 9 2
17 16 4 9 13 1 10 9 2 13 11 11 2 9 9 10 9 2
2 0 9
17 1 11 15 10 0 2 7 3 0 9 1 9 0 9 13 13 2
8 0 9 3 13 3 12 9 2
6 1 9 13 0 9 2
18 3 15 1 15 13 1 9 1 9 2 7 13 9 9 1 9 9 2
9 3 2 16 13 9 7 1 9 2
4 15 14 13 2
37 16 4 13 2 16 1 0 9 0 9 13 3 15 2 15 13 0 15 1 15 13 2 13 3 3 3 2 16 15 4 3 13 2 13 11 11 2
11 1 9 9 1 9 13 9 9 1 9 2
15 1 15 13 13 0 9 0 9 2 15 15 1 9 13 2
8 1 11 13 10 9 3 0 2
18 15 3 13 9 2 15 4 1 15 13 0 9 13 2 13 11 11 2
17 9 15 3 13 7 0 9 9 2 1 15 4 1 0 9 13 2
23 1 9 15 13 3 9 0 9 2 0 9 9 2 13 15 1 9 0 9 9 1 9 2
3 13 13 9
15 0 9 15 13 3 10 9 9 9 2 1 15 9 13 2
14 1 12 9 13 1 0 9 2 1 12 9 1 0 2
22 1 10 9 3 13 2 16 0 9 3 13 9 1 12 9 9 2 9 1 12 9 2
14 9 1 12 9 2 9 2 7 12 9 2 9 2 2
16 1 15 3 3 13 9 2 16 10 9 15 13 3 0 9 2
8 9 9 13 0 1 9 9 2
14 0 9 13 2 16 15 13 10 9 13 10 0 9 2
18 7 4 1 15 13 9 9 7 0 9 1 9 7 9 13 7 3 2
17 13 15 3 11 2 11 7 0 2 16 4 10 9 13 9 13 2
1 3
11 9 11 1 9 9 15 13 11 1 9 2
20 0 9 0 0 9 9 1 11 13 0 9 11 2 11 7 13 1 0 9 2
3 0 9 13
2 11 2
38 0 9 9 9 9 12 11 11 1 11 2 9 9 11 2 11 2 4 13 1 0 9 0 9 11 1 11 7 13 9 9 1 12 9 9 0 11 2
44 0 9 0 0 9 2 11 2 1 11 13 0 9 0 9 11 2 15 13 11 1 15 2 16 13 9 9 9 0 9 11 12 2 9 1 11 7 13 1 9 0 0 9 2
6 11 7 11 11 1 9
10 3 0 0 9 0 9 3 13 10 9
2 11 11
19 1 9 1 0 0 9 15 9 13 1 0 9 0 9 2 13 9 9 2
18 1 0 0 9 15 7 3 9 3 3 13 7 13 12 9 2 9 2
30 9 13 3 0 2 7 13 2 16 4 0 0 9 13 13 3 0 16 1 0 9 2 3 13 14 12 9 2 9 2
11 13 4 1 15 0 9 0 16 12 9 2
10 3 15 15 13 1 9 13 1 0 2
20 0 9 4 3 13 9 0 9 2 15 3 13 1 12 5 1 0 12 9 2
11 13 7 9 9 1 9 9 1 0 9 2
21 3 1 15 13 0 12 2 7 15 0 0 9 2 11 2 7 9 9 11 11 2
36 16 9 9 11 13 0 9 2 15 13 2 16 10 9 13 1 12 5 1 12 9 2 9 11 15 13 1 9 3 3 7 13 1 12 9 2
12 10 9 15 3 13 1 0 9 3 1 9 2
21 16 15 15 13 2 16 9 9 10 9 15 1 0 3 13 9 3 2 13 9 2
11 0 9 3 13 12 2 3 0 9 9 2
30 7 3 3 13 1 0 9 9 1 0 9 2 1 12 15 13 9 12 2 1 11 2 15 10 9 3 13 0 9 2
11 7 3 15 13 0 9 2 15 13 3 2
32 10 9 13 1 12 5 1 12 9 7 9 2 3 13 10 9 1 9 1 12 9 2 15 13 0 9 2 13 3 1 15 2
13 10 9 4 13 2 16 3 13 2 1 15 0 2
52 3 0 13 1 10 9 7 9 0 9 2 12 2 2 7 7 1 9 0 9 13 12 9 1 9 9 7 13 2 3 16 0 9 9 13 12 5 2 14 1 9 9 9 9 2 15 13 10 9 3 0 2
19 7 0 9 12 9 13 1 9 1 0 9 2 12 9 2 3 3 0 2
29 0 9 13 3 11 2 7 15 7 1 0 9 2 12 9 2 9 2 2 7 1 9 2 12 9 2 9 2 2
18 1 12 0 9 9 1 9 15 3 13 9 12 2 2 2 0 9 2
9 13 15 2 16 15 0 9 13 2
3 7 3 0
2 11 2
30 9 9 11 11 11 4 13 1 9 1 0 9 1 0 9 9 9 11 9 11 2 11 11 2 9 2 12 2 9 2
15 9 2 15 13 0 0 9 2 13 1 9 9 9 11 2
13 0 7 0 9 11 13 0 9 1 10 9 3 2
3 13 9 2
2 11 2
34 7 0 0 9 0 9 2 15 13 0 9 1 9 1 9 9 9 2 1 9 9 11 9 11 13 1 9 10 9 9 1 10 9 2
14 9 7 9 1 0 9 12 9 1 9 9 3 13 2
6 3 15 4 13 9 2
5 11 2 11 2 2
19 12 9 1 0 9 11 1 11 13 0 2 3 15 4 10 0 9 13 2
14 1 11 15 3 13 9 9 2 7 3 13 0 9 2
42 16 3 4 3 13 2 9 11 2 15 13 1 0 9 9 1 9 2 13 9 1 9 11 1 9 2 16 13 0 9 7 0 9 2 1 15 10 9 9 9 13 2
31 13 4 15 3 13 9 11 11 11 2 9 2 0 2 9 2 2 11 11 2 7 10 9 2 16 13 9 2 4 13 2
12 9 11 13 1 11 13 2 14 13 3 13 2
10 14 1 0 9 15 13 3 9 9 2
15 1 9 15 3 3 13 7 9 0 9 9 0 9 11 2
24 1 10 9 13 0 9 2 16 4 9 13 4 3 13 7 13 2 13 15 10 9 9 11 2
24 3 3 15 13 1 0 9 11 11 12 2 16 13 9 1 9 7 0 9 1 9 0 9 2
4 13 9 11 11
2 11 2
30 3 0 0 9 1 9 0 0 9 11 11 11 2 15 15 3 1 9 13 1 0 9 1 9 0 11 2 13 9 2
26 1 0 9 9 13 9 9 11 11 1 0 9 3 12 9 1 9 2 3 4 3 1 9 13 9 2
24 1 0 11 11 2 15 3 13 9 1 0 9 1 9 1 9 2 13 1 12 9 12 9 2
10 9 15 13 12 9 3 1 0 9 2
2 9 9
2 11 2
15 9 11 15 13 1 12 2 1 12 2 9 9 1 11 2
35 1 9 13 9 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2
3 1 0 9
16 11 13 9 11 2 11 2 1 9 9 9 1 12 2 12 2
3 9 0 9
11 0 0 11 2 11 2 0 9 12 2 12
7 11 2 11 2 11 2 2
37 3 16 1 9 1 0 9 1 11 2 12 2 12 2 13 0 9 7 1 11 1 9 0 9 0 11 10 0 9 3 3 2 3 12 2 12 2
28 16 1 0 9 9 0 9 13 2 1 0 9 13 0 9 1 12 2 9 14 11 2 11 2 11 7 11 2
21 9 13 0 9 0 9 2 7 7 15 1 0 9 9 13 1 0 9 0 9 2
24 9 0 9 0 9 3 13 0 9 2 3 3 1 9 0 9 13 0 7 1 0 9 0 2
19 0 9 9 1 0 0 9 13 3 14 9 1 9 9 0 9 11 11 2
25 1 0 9 9 13 0 9 11 14 11 10 0 9 2 15 13 1 0 9 13 9 1 0 9 2
25 1 12 2 9 3 7 9 1 9 11 2 11 2 11 2 11 13 1 0 9 2 12 2 12 2
16 1 12 9 13 1 12 2 12 11 2 15 1 9 13 11 2
31 1 11 13 1 12 2 9 13 11 2 12 2 12 2 2 7 12 9 1 9 12 13 1 0 9 1 12 2 12 11 2
13 13 15 0 9 7 1 11 13 10 9 3 0 2
11 1 0 0 9 13 3 9 1 9 9 2
20 1 0 9 13 12 9 9 1 9 7 9 15 13 9 14 1 12 2 9 2
16 15 11 3 13 0 9 1 0 0 9 7 3 13 9 11 2
13 15 13 3 1 11 0 9 7 13 15 13 11 2
10 1 10 9 4 1 9 9 3 13 2
22 7 7 0 9 0 12 13 9 11 1 9 11 2 15 0 9 11 13 12 9 9 2
20 15 13 9 9 1 9 7 1 9 7 9 1 10 9 0 0 9 15 13 2
2 11 2
8 9 2 11 2 11 2 11 2
3 9 1 9
5 11 11 2 9 11
29 2 13 4 15 1 9 16 1 9 1 11 2 7 3 16 1 3 0 9 2 3 4 10 0 9 13 13 9 2
4 14 4 13 2
20 1 9 9 4 13 2 16 13 7 13 7 9 1 0 9 1 11 1 11 2
28 11 11 2 9 0 9 2 10 9 13 1 9 1 9 1 11 0 9 1 15 2 16 4 13 1 0 9 2
15 3 15 13 2 16 0 13 13 14 0 9 0 1 9 2
4 11 13 1 11
11 11 13 3 7 13 1 12 2 9 0 0
8 0 11 2 11 2 11 2 2
33 1 0 9 11 11 2 13 1 15 1 0 9 2 13 1 12 2 9 0 0 7 0 9 11 11 2 0 16 9 2 12 2 2
10 1 0 11 0 9 13 0 11 11 2
33 3 15 3 13 11 11 2 15 1 12 2 9 13 11 11 2 3 15 1 9 13 12 2 12 2 12 2 12 2 12 2 12 2
13 13 3 0 2 13 4 3 3 2 13 0 11 2
34 0 11 13 0 9 2 1 0 0 13 12 9 1 0 9 7 1 9 13 1 0 9 12 2 12 2 15 1 9 1 10 9 13 2
39 1 0 0 9 11 11 2 12 2 9 11 2 15 15 13 0 0 9 2 12 2 12 2 12 2 12 2 12 2 12 2 12 2 12 2 12 2 12 2
8 3 4 13 0 9 10 9 2
14 3 1 0 9 4 13 13 0 9 2 13 15 9 2
24 9 1 0 9 13 0 9 11 1 10 0 9 1 0 0 2 3 15 1 12 9 13 9 2
18 11 11 13 11 11 11 12 2 12 2 12 2 12 2 12 2 12 2
30 0 9 10 0 0 9 11 11 1 11 2 12 2 13 10 9 11 11 12 2 12 2 12 2 12 2 12 2 12 2
24 3 15 13 3 0 9 11 11 2 15 3 13 1 11 11 11 12 2 12 2 12 2 12 2
25 7 9 13 1 9 1 9 2 15 15 0 9 13 2 7 13 10 12 0 9 1 0 12 9 2
14 3 3 0 9 4 15 13 0 2 16 4 3 13 2
16 1 9 4 7 13 13 7 3 15 13 15 3 2 13 11 2
4 11 13 1 11
3 0 11 2
25 9 1 9 0 12 9 9 16 9 0 9 0 9 13 3 0 9 11 11 2 7 11 11 11 2
37 9 2 0 1 0 9 9 2 13 12 9 13 9 1 9 0 9 2 9 7 0 9 1 9 9 1 9 7 1 0 9 2 13 9 12 9 2
4 11 13 1 11
5 11 13 13 1 11
2 0 11
7 11 2 11 2 11 2 2
19 0 9 0 11 13 9 11 11 2 15 13 1 9 1 9 9 1 11 2
20 11 13 1 9 9 11 2 3 13 1 11 2 7 15 15 9 13 1 11 2
10 3 15 7 13 3 1 9 2 9 2
26 11 4 15 13 1 0 9 3 13 1 0 0 9 1 11 11 2 3 7 11 13 1 0 9 11 2
10 11 13 9 11 7 1 15 14 13 2
14 1 9 13 1 0 9 13 2 13 15 0 9 11 2
30 11 11 3 13 9 1 11 2 7 1 0 9 15 13 9 2 16 1 9 1 0 2 11 13 0 9 1 9 11 2
9 10 9 15 3 3 13 1 9 2
9 11 7 3 13 13 0 9 11 2
6 1 9 9 3 13 2
3 2 11 2
4 9 13 0 9
10 11 14 13 1 11 1 9 0 2 11
9 11 2 11 2 11 2 11 2 2
27 16 4 13 0 9 9 9 1 9 1 0 0 9 1 9 2 13 15 12 2 0 9 3 3 7 3 2
25 0 13 13 2 16 11 13 0 9 7 1 9 1 0 2 11 7 16 11 1 11 13 9 9 2
13 9 13 12 0 9 11 2 11 7 11 2 11 2
5 3 13 0 9 2
31 11 4 1 11 13 0 11 7 0 11 2 1 9 9 7 9 13 11 2 15 13 0 0 9 2 7 13 4 13 0 2
21 0 2 11 4 13 3 1 9 7 0 9 11 11 2 15 15 13 9 1 11 2
15 3 7 13 0 0 9 7 13 2 16 13 1 9 13 2
11 9 11 11 15 7 13 9 10 9 13 2
24 1 11 4 13 3 3 1 9 9 13 11 2 13 13 7 9 1 11 2 3 13 9 11 2
15 1 9 15 1 9 13 11 2 13 7 4 1 9 11 2
11 0 4 13 11 2 15 13 9 1 9 2
19 9 11 11 1 11 13 0 9 11 2 15 11 13 1 11 1 0 9 2
2 0 9
2 11 2
20 11 4 13 0 9 3 1 0 9 0 11 2 15 1 0 9 13 3 11 2
19 1 11 13 1 0 0 9 0 9 2 3 7 1 11 2 3 13 11 2
15 15 4 13 0 9 11 2 15 13 9 9 11 11 11 2
7 1 9 1 11 13 11 2
8 11 13 1 11 1 0 9 2
34 3 13 0 11 2 3 1 0 9 4 1 9 13 11 2 16 15 9 11 1 9 3 13 2 16 1 10 0 9 7 0 9 13 2
16 0 9 9 13 11 7 9 13 7 11 2 15 13 1 11 2
19 0 9 11 13 9 1 9 2 11 2 11 2 11 7 11 13 0 9 2
3 0 9 9
2 11 11
9 1 14 3 0 9 15 9 13 2
28 13 15 7 9 11 2 15 15 13 0 9 1 10 9 1 0 9 1 11 3 2 16 13 1 9 9 13 2
14 15 2 15 0 9 13 2 14 13 9 12 12 9 2
15 13 15 2 16 4 4 0 9 13 9 9 2 3 3 2
27 13 15 3 0 9 1 0 9 1 9 9 2 16 9 15 15 13 9 3 15 13 7 3 15 7 13 2
6 13 15 3 14 15 2
24 3 2 13 4 1 9 15 9 0 2 16 4 1 9 9 13 3 1 11 9 9 1 9 2
4 11 13 0 9
7 11 2 11 2 11 2 2
21 1 0 9 1 11 7 11 2 12 2 12 2 15 9 13 9 14 1 0 9 2
16 12 0 9 13 0 9 7 9 3 13 13 0 9 12 9 2
26 3 0 9 12 2 9 1 11 3 13 13 9 1 9 0 9 2 15 4 13 0 9 12 2 9 2
5 13 4 3 3 2
33 14 16 4 13 1 9 9 2 7 3 15 3 3 13 2 13 9 7 9 11 11 9 2 15 13 9 12 9 7 1 0 9 2
15 9 13 14 11 9 2 1 15 13 12 9 13 9 9 2
22 1 9 13 9 11 2 15 10 0 9 13 0 9 7 13 7 1 9 12 0 9 2
23 1 0 9 13 0 2 1 0 15 9 13 2 7 11 9 3 11 13 7 13 14 11 2
35 3 1 0 9 13 11 9 9 2 9 11 1 15 13 2 9 2 15 13 1 10 9 13 11 7 11 2 13 2 15 15 13 2 2 2
28 1 9 9 3 13 2 0 9 1 0 9 4 3 13 2 0 9 4 13 3 1 9 2 16 4 13 3 2
29 9 13 1 11 0 9 2 16 4 1 9 13 9 1 11 2 16 13 4 9 11 3 13 1 9 1 9 9 2
16 16 11 9 13 2 4 7 1 9 13 11 2 13 9 11 2
19 1 9 13 3 16 12 12 9 2 13 7 9 2 10 9 13 9 13 2
29 13 0 9 1 11 2 0 9 2 1 15 15 13 0 9 9 2 14 1 0 9 1 9 3 12 9 1 9 2
16 3 7 3 2 16 4 13 15 9 7 16 10 9 4 13 2
24 1 10 9 15 3 7 13 13 9 9 2 15 15 1 9 1 9 13 15 2 16 13 9 2
14 10 9 14 10 0 9 13 1 0 9 2 2 2 2
24 1 9 12 2 9 12 2 0 9 11 2 11 2 12 2 12 2 15 0 11 13 13 0 11
2 9 11
5 9 1 9 1 9
6 9 13 9 0 0 9
5 9 2 11 2 2
22 0 9 1 12 9 7 9 15 13 1 9 9 1 0 9 9 1 0 9 1 9 2
26 1 9 12 9 13 11 11 2 0 9 0 3 1 9 2 1 9 2 2 7 0 9 0 9 11 2
13 9 1 9 13 0 1 15 2 3 4 9 13 2
15 1 10 10 9 1 9 13 7 9 9 1 9 11 9 2
10 3 4 13 1 0 9 1 9 9 2
16 0 9 9 4 13 1 11 7 3 1 15 13 9 1 9 2
18 14 7 1 0 2 15 13 10 9 7 16 13 9 2 7 15 13 2
39 0 9 1 11 2 11 2 9 11 7 11 15 9 9 13 2 3 7 16 0 9 13 9 13 7 9 3 13 2 15 15 13 1 9 2 16 15 13 2
10 1 0 9 15 15 13 1 0 9 2
8 0 9 13 0 9 3 0 2
8 9 13 1 9 9 3 3 2
14 16 4 3 13 3 9 2 7 3 13 12 3 0 2
14 3 13 9 2 16 0 9 13 0 16 10 0 0 2
6 13 15 15 12 9 2
16 13 1 9 3 0 9 7 3 14 3 13 0 9 1 9 2
15 16 13 2 11 13 9 13 1 9 7 1 9 15 13 2
20 9 11 3 13 0 16 15 2 15 13 0 0 9 2 7 9 13 3 0 2
18 3 7 9 13 1 0 9 13 9 7 1 0 9 15 13 15 9 2
17 0 9 13 1 15 2 16 3 13 0 9 3 3 9 1 9 2
5 3 13 9 0 2
9 0 9 7 13 9 3 9 11 2
4 13 1 9 2
18 0 9 3 13 1 9 7 9 4 13 13 9 1 0 9 1 9 2
8 1 10 9 3 13 10 9 2
18 1 11 2 11 7 11 13 13 3 1 9 2 11 2 11 7 11 2
16 13 3 12 9 2 1 15 12 13 9 1 9 1 0 9 2
4 11 13 1 9
9 1 9 14 13 0 9 2 7 9
6 0 11 2 11 2 2
26 15 3 13 0 9 11 11 1 9 2 3 12 2 9 11 2 2 15 3 15 15 13 1 0 11 2
18 1 9 12 13 11 1 12 2 9 0 0 2 15 13 10 0 9 2
34 1 10 9 13 10 9 1 0 11 3 0 9 2 15 13 7 0 9 2 1 0 0 9 9 15 11 11 11 13 1 12 2 9 2
9 16 3 13 2 3 15 13 13 2
13 13 2 15 15 13 2 7 3 15 15 3 13 2
27 3 15 13 2 3 3 3 13 2 13 1 9 11 2 15 1 9 13 1 9 9 2 0 1 0 9 2
14 13 4 1 15 2 16 1 15 0 3 4 14 13 2
27 0 9 0 9 13 1 0 9 1 0 9 0 9 2 0 9 1 0 9 2 15 15 1 0 0 13 2
32 13 15 1 10 9 13 2 13 2 15 13 2 13 15 11 2 1 0 9 7 10 9 13 13 2 3 13 0 9 2 2 2
16 11 13 2 16 13 0 9 2 16 1 15 15 13 0 11 2
27 13 15 0 9 2 3 15 3 13 1 9 2 3 1 0 9 2 16 3 15 13 9 2 13 0 9 2
9 0 9 3 13 9 1 10 9 2
8 3 0 9 3 13 0 9 2
29 0 9 0 11 2 12 2 9 11 2 15 3 13 3 0 9 2 1 0 9 1 10 9 14 3 13 0 9 2
11 9 9 15 1 0 9 13 9 11 11 2
5 9 11 1 9 13
2 11 2
30 0 0 9 11 0 11 13 1 10 9 1 9 1 0 9 12 9 2 15 13 1 12 9 3 16 1 0 9 12 2
5 3 13 12 9 2
17 1 9 13 1 0 9 9 9 0 9 11 1 9 1 0 9 2
20 1 10 9 4 15 9 11 2 15 15 10 9 13 2 1 12 9 3 13 2
49 9 10 9 1 11 13 0 9 9 1 0 9 1 9 2 3 2 9 9 11 11 13 1 9 12 3 12 9 2 1 9 12 9 2 2 9 11 11 11 12 9 2 3 1 9 12 9 2 2
20 1 9 12 9 1 0 9 9 11 13 7 13 1 15 1 0 9 0 9 2
25 9 11 13 2 16 7 1 0 9 13 9 9 1 9 1 0 0 9 2 3 1 11 12 2 2
5 0 9 9 13 2
7 11 2 9 11 11 2 2
21 10 9 13 2 16 1 9 1 3 0 9 0 9 13 3 9 0 2 3 0 2
21 9 9 2 9 2 1 10 0 9 2 9 2 13 0 9 9 0 0 9 9 2
15 15 13 9 1 9 1 0 9 0 0 9 2 9 2 2
14 13 15 15 13 10 9 9 2 15 13 0 0 9 2
17 1 9 0 15 13 3 13 2 9 2 7 3 0 0 9 9 2
13 3 4 1 9 13 9 9 2 9 2 16 9 2
16 13 13 7 9 9 2 9 9 4 13 9 9 2 9 2 2
29 1 0 9 13 10 9 0 9 1 9 11 11 2 11 1 0 9 12 2 12 2 15 13 1 0 9 0 9 2
4 0 9 3 0
5 11 2 11 2 2
36 9 1 9 7 9 9 11 15 13 13 9 9 9 1 9 12 2 3 3 0 9 11 11 13 1 9 9 1 11 12 9 0 9 7 11 2
24 12 1 0 9 0 9 13 9 2 10 9 3 13 0 9 9 11 1 0 9 7 0 9 2
12 9 1 9 15 13 1 9 11 12 2 9 2
16 0 12 9 3 1 3 0 9 9 13 0 9 7 1 11 2
19 11 7 0 9 4 13 2 0 4 13 1 9 7 0 3 13 7 13 2
11 3 12 2 9 4 13 0 9 0 9 2
9 13 15 12 2 1 15 12 9 2
9 1 12 1 15 13 13 9 9 2
50 0 9 9 11 1 9 11 2 11 2 11 7 0 3 3 13 1 15 2 3 4 9 13 2 13 12 9 9 2 13 2 16 4 9 13 13 9 0 2 16 4 4 1 9 3 13 10 0 9 2
28 0 9 11 13 7 1 15 2 16 4 13 9 9 2 16 4 13 0 9 2 15 4 3 13 1 9 9 2
17 9 0 9 13 13 9 0 9 1 9 2 3 13 0 0 9 2
17 3 12 2 9 4 13 9 7 12 2 9 4 0 12 0 13 2
21 13 15 14 9 9 0 3 1 0 9 7 0 9 2 15 13 13 1 12 9 2
8 11 0 9 1 9 9 3 13
5 11 2 11 2 2
31 0 0 9 1 0 0 9 2 1 15 13 9 0 9 11 11 9 7 9 9 9 1 11 11 2 4 3 13 1 9 2
33 0 9 0 13 1 9 11 11 9 1 9 2 16 4 1 15 13 10 9 1 9 11 9 11 1 9 1 11 1 10 0 9 2
25 0 9 9 0 9 1 9 12 13 9 11 3 0 9 2 1 15 9 11 13 10 9 9 0 2
23 7 15 15 2 16 13 3 9 0 9 2 1 15 13 9 11 9 11 2 0 9 9 2
6 9 13 9 0 9 2
20 11 3 1 9 13 1 9 11 2 15 15 13 9 13 7 13 15 9 12 2
9 10 9 13 1 9 1 0 9 2
25 11 1 10 9 13 9 9 11 11 2 0 9 11 2 16 4 15 13 1 0 9 1 9 9 2
17 11 13 9 9 0 9 7 1 10 9 1 11 2 7 1 11 2
39 11 1 9 11 13 1 0 2 16 4 13 10 9 0 2 16 4 1 15 13 3 2 16 15 15 3 13 9 9 2 7 1 9 4 15 9 13 3 2
18 3 2 16 9 13 9 0 0 9 2 13 0 9 11 9 1 9 2
25 0 9 13 3 2 9 0 9 11 2 15 4 15 13 1 15 2 16 9 13 9 2 7 11 2
10 11 2 1 9 0 9 15 13 3 13
5 11 2 11 2 2
23 9 0 9 1 9 1 9 1 9 9 9 9 11 9 13 3 0 9 9 11 11 11 2
16 0 9 1 0 7 0 9 13 10 9 1 9 0 9 9 2
26 16 13 9 11 1 9 11 2 1 9 0 9 4 9 13 7 15 15 15 1 10 9 13 1 9 2
12 1 10 9 15 13 3 13 2 13 3 11 2
16 1 0 9 10 9 13 11 9 9 15 1 9 0 0 9 2
33 16 15 10 9 13 2 4 15 13 16 0 9 2 15 15 13 2 3 13 0 9 7 1 10 9 13 9 0 9 2 13 11 2
12 13 15 9 9 2 7 13 0 9 0 9 2
16 10 9 13 13 14 1 9 0 9 1 0 9 2 13 11 2
5 0 9 15 13 13
10 1 9 4 15 13 13 1 9 0 9
5 11 2 11 2 2
25 9 2 15 13 0 9 0 9 0 9 2 15 3 13 13 1 0 9 9 9 9 7 9 9 2
31 1 9 11 2 11 2 11 2 11 7 10 9 11 2 11 7 11 2 11 15 9 13 7 9 0 9 9 11 2 11 2
21 9 1 0 9 13 0 9 2 3 11 2 11 13 1 9 0 9 0 9 13 2
18 0 9 13 9 1 9 0 9 0 9 1 9 9 1 9 0 9 2
18 9 0 9 13 0 9 9 7 10 9 13 13 3 1 9 0 9 2
32 1 9 0 9 15 13 11 9 1 0 9 1 9 12 9 9 7 13 12 9 1 11 2 1 0 9 0 7 9 1 9 2
27 3 10 9 15 13 12 1 9 2 1 15 15 0 0 9 13 13 9 9 7 3 7 9 9 7 9 2
29 9 9 0 2 0 2 11 2 2 15 1 0 9 9 0 9 3 13 2 15 1 10 0 9 1 9 3 13 2
32 3 13 9 9 9 11 1 10 9 1 0 0 9 2 3 13 2 16 0 9 4 15 13 13 2 16 10 9 13 3 13 2
18 11 2 11 3 13 9 2 16 4 15 13 13 9 0 9 0 9 2
19 9 0 2 0 2 11 2 13 0 9 0 9 1 10 9 1 9 9 2
50 0 2 0 2 11 2 3 3 13 9 1 9 0 9 2 15 15 13 1 9 9 9 15 9 0 0 2 9 2 9 1 9 12 2 12 2 12 2 3 0 9 13 9 1 9 0 9 0 9 2
30 1 0 9 9 0 2 0 2 11 2 9 2 3 0 9 13 7 0 9 9 2 13 9 9 2 12 1 9 12 2
22 1 15 13 13 2 16 9 13 13 1 10 9 3 0 9 2 16 13 9 3 9 2
12 1 0 9 13 9 0 9 13 9 9 3 2
48 9 0 9 13 2 16 1 9 1 0 0 9 1 10 0 9 13 9 9 1 10 0 9 7 16 4 9 13 2 13 13 1 9 0 9 13 9 9 9 1 0 12 9 14 1 12 9 2
5 9 0 9 1 11
2 0 9
2 11 11
13 13 13 1 9 0 12 0 9 2 11 7 11 2
33 1 15 15 3 3 13 9 0 9 2 16 4 1 10 0 9 13 15 3 3 0 9 7 13 1 15 0 9 0 9 0 9 2
25 1 0 9 0 9 1 0 7 3 0 9 15 11 7 11 2 0 9 0 9 2 13 3 9 2
18 3 1 15 13 9 1 9 0 0 0 9 11 2 11 7 11 11 2
39 9 10 9 13 0 1 12 9 1 0 0 9 2 1 0 9 0 2 11 7 11 9 9 7 9 0 2 13 1 12 0 0 9 9 11 7 11 9 2
12 3 7 1 11 7 11 13 11 7 11 12 2
26 1 9 12 13 0 2 14 1 9 0 9 2 16 1 0 0 9 13 3 9 3 1 12 0 9 2
23 9 15 13 2 16 15 1 10 0 9 13 12 0 0 9 2 15 13 0 9 1 11 2
14 3 0 9 9 13 1 10 9 12 9 3 0 9 2
12 15 15 13 9 0 9 2 9 2 14 9 2
31 16 15 3 12 13 2 16 0 13 1 12 9 0 9 0 9 1 9 2 13 15 9 3 13 7 13 7 0 0 9 2
29 9 15 15 3 13 13 14 9 0 1 0 9 2 15 1 15 3 13 2 14 7 1 0 9 2 15 13 12 2
12 0 9 15 3 0 9 15 15 3 13 0 2
13 16 15 0 9 13 9 2 13 11 1 0 9 2
14 13 9 15 0 0 9 2 16 13 11 9 7 9 2
26 11 2 15 15 10 9 13 13 2 13 9 2 1 15 13 2 16 15 13 9 7 16 9 13 11 2
24 11 2 15 15 0 9 13 13 2 13 0 2 3 0 9 2 1 15 13 2 16 11 13 2
32 11 2 15 15 0 9 13 13 2 1 15 13 2 16 15 13 2 7 16 11 3 13 2 7 15 14 13 2 15 3 13 2
22 16 13 9 9 2 1 15 13 9 0 9 2 13 15 13 9 1 0 9 15 0 2
22 16 13 1 9 9 2 0 3 9 0 9 2 13 15 12 9 9 0 1 0 9 2
9 9 15 13 9 1 9 0 9 2
12 13 15 0 9 2 15 13 7 1 0 9 2
14 9 15 1 9 10 9 7 1 9 9 9 3 13 2
15 12 9 13 11 7 11 0 1 15 2 12 1 9 9 2
4 13 15 3 2
20 0 9 2 15 1 9 1 0 9 0 0 9 13 0 9 2 15 13 9 2
3 0 0 9
1 11
5 11 11 2 11 0
8 9 13 2 13 15 0 9 2
12 0 9 13 2 9 15 13 13 1 0 9 2
17 3 10 9 15 7 1 11 13 9 1 0 9 7 9 0 9 2
19 3 0 9 13 1 9 1 11 1 9 3 0 9 9 1 0 9 9 2
22 9 0 9 3 13 2 16 4 13 9 0 7 1 0 9 2 3 1 0 0 9 2
5 9 3 13 9 2
22 9 9 15 13 7 9 1 9 1 11 7 0 9 2 15 13 3 0 9 11 11 2
41 9 0 9 2 9 0 9 2 15 13 1 9 0 9 1 9 2 13 2 16 0 9 15 13 14 1 9 2 16 4 13 0 9 2 3 3 1 9 0 9 2
26 9 13 3 1 9 10 0 9 2 10 9 2 3 9 9 1 0 9 2 13 9 12 0 9 3 2
9 16 9 10 9 13 14 9 11 2
19 7 0 9 15 2 16 9 7 9 13 1 9 9 2 13 0 0 9 2
20 9 9 3 13 1 15 2 16 9 13 1 9 0 9 9 0 9 10 9 2
20 1 9 1 9 9 13 9 1 0 9 9 1 9 2 13 15 0 0 9 2
9 7 3 7 13 1 9 9 9 2
13 9 10 9 13 2 3 1 10 9 2 0 9 2
23 7 1 9 0 9 1 9 9 13 1 0 9 0 13 9 9 2 15 13 1 9 3 2
6 1 9 1 9 7 3
14 0 9 3 13 2 9 2 13 13 10 7 15 9 2
40 3 1 0 3 0 0 9 1 9 12 13 0 3 13 3 0 0 9 2 1 10 9 13 12 1 0 0 9 2 0 9 2 15 1 0 9 13 9 2 2
16 1 12 9 3 2 1 0 0 9 2 9 13 3 3 3 2
17 9 13 10 2 3 9 9 0 9 2 9 9 1 9 2 2 2
25 9 14 3 13 2 16 9 9 2 3 15 13 1 9 9 2 13 1 0 7 0 9 3 0 2
9 1 15 3 13 0 0 9 9 2
8 3 0 13 0 9 1 9 2
11 9 9 4 3 1 9 13 16 9 9 2
14 9 10 9 15 9 13 16 9 0 9 1 0 9 2
3 7 3 2
13 9 15 3 13 2 16 1 9 13 9 0 11 2
10 3 3 13 9 15 1 9 9 13 2
4 9 1 0 9
7 9 7 13 1 0 9 2
13 1 0 9 2 0 7 0 2 7 4 13 15 2
7 4 3 7 3 13 9 2
12 9 13 9 1 9 9 2 7 9 15 13 2
13 13 3 0 2 16 4 15 9 13 10 9 13 2
30 16 4 15 15 7 13 2 9 1 9 0 4 15 13 12 1 0 9 0 9 11 11 1 0 9 2 7 14 15 2
19 13 2 14 15 9 1 10 9 2 4 13 13 13 9 0 9 1 9 2
37 16 15 7 9 13 13 9 9 11 2 3 15 9 13 9 0 9 1 9 9 9 7 9 1 0 0 9 13 13 1 0 0 9 9 0 9 2
15 1 10 9 15 13 14 3 13 2 16 4 9 13 0 2
16 3 15 13 7 1 9 2 15 4 1 0 9 14 3 13 2
9 7 15 13 2 16 9 13 0 2
33 9 15 13 9 2 7 13 9 1 9 2 13 3 0 9 9 11 11 2 15 13 13 9 9 7 9 1 0 9 1 0 9 2
3 9 0 9
9 9 0 9 1 11 13 3 11 11
4 11 11 2 11
32 1 11 13 3 13 9 2 16 1 0 7 0 9 13 9 3 11 11 2 15 16 0 9 1 9 12 13 9 13 0 9 2
27 1 9 12 3 13 3 9 0 9 2 11 2 1 12 12 9 2 16 3 15 1 0 9 13 3 9 2
27 1 0 9 13 0 9 12 7 12 9 1 0 9 9 11 2 3 13 15 3 12 9 2 0 9 2 2
5 11 11 9 9 13
35 1 9 1 0 9 0 9 7 1 9 9 11 11 2 11 11 7 11 11 7 13 2 16 0 9 4 15 3 16 3 13 1 0 9 2
27 16 15 11 11 10 0 9 10 0 9 1 0 11 3 13 2 7 14 2 13 0 2 16 15 15 13 2
28 13 0 2 16 16 4 9 13 0 9 1 9 11 3 1 12 7 12 9 2 13 4 0 0 9 3 0 2
15 9 11 13 7 3 0 9 7 10 9 9 1 9 13 2
25 1 9 3 13 2 16 3 1 9 12 13 9 9 11 2 16 15 1 11 4 0 9 3 13 2
11 13 15 15 9 7 0 0 7 0 9 2
31 0 9 11 13 3 1 9 2 16 1 9 9 1 11 2 11 7 0 9 13 0 9 1 9 2 9 1 9 3 13 2
21 2 0 0 9 3 13 10 9 9 9 2 16 3 12 5 13 1 9 9 2 2
4 9 1 0 9
18 9 13 0 9 1 11 3 13 9 9 9 11 1 0 7 0 9 2
13 0 0 9 13 1 9 9 10 9 9 9 13 2
19 9 13 3 0 9 2 13 15 9 9 1 9 1 0 9 1 0 9 2
7 15 7 13 13 1 9 2
16 1 0 9 13 0 2 16 1 15 13 9 2 15 13 13 2
10 14 3 13 9 13 13 1 0 9 2
6 0 9 7 13 9 2
20 0 13 7 9 2 15 1 9 9 13 10 9 9 2 15 13 1 10 9 2
43 7 3 1 0 9 2 9 2 13 1 12 12 9 1 0 12 2 1 11 2 0 9 2 0 9 2 12 1 12 12 7 1 11 2 0 9 2 12 9 1 0 12 2
21 9 3 13 2 16 1 9 1 0 9 9 1 9 4 9 1 9 0 9 13 2
12 3 1 15 13 13 0 9 7 9 13 9 2
22 9 15 13 9 13 1 10 0 9 3 9 1 9 12 9 9 1 9 9 0 9 2
11 9 0 9 13 7 3 0 16 0 9 2
3 0 9 9
22 1 9 1 0 9 13 3 7 3 0 9 9 9 16 0 2 3 0 9 1 9 2
28 0 9 3 1 12 9 13 9 9 0 9 2 9 11 2 0 9 0 0 9 7 10 0 0 9 11 11 2
26 13 15 0 9 1 9 2 3 15 11 13 7 11 13 1 9 2 10 0 9 13 3 3 9 11 2
14 15 15 13 1 9 13 1 0 9 0 1 9 9 2
11 3 15 13 15 2 16 13 3 0 9 2
21 3 15 13 13 7 15 2 16 9 2 15 11 13 1 9 2 3 14 13 11 2
18 11 3 13 7 11 15 13 9 9 11 11 13 0 9 11 2 12 2
23 11 2 3 16 11 7 11 2 13 3 9 10 9 2 7 1 9 12 13 7 12 9 2
22 13 10 9 2 16 3 13 13 15 3 2 16 3 13 9 0 9 1 9 0 11 2
23 0 9 3 13 2 16 9 1 0 9 13 1 9 9 1 0 9 2 1 9 0 11 2
27 11 13 0 9 2 10 9 13 0 9 1 0 9 7 13 0 13 9 1 0 9 1 0 7 0 9 2
17 3 13 0 13 0 9 2 16 9 11 7 9 11 10 9 13 2
19 13 15 13 9 1 11 7 13 15 3 1 0 9 2 1 9 0 2 2
3 9 0 9
30 13 0 2 16 7 1 3 0 9 0 9 2 3 9 1 9 9 3 13 2 13 9 2 16 13 1 9 1 11 2
20 11 7 11 1 9 2 3 13 13 1 9 0 9 2 13 7 15 13 3 2
10 1 0 9 7 9 0 9 3 13 2
10 10 9 3 1 9 0 9 3 13 2
1 3
30 0 9 1 0 9 11 7 0 11 1 9 13 9 13 1 9 0 9 11 0 0 9 0 0 0 1 12 9 9 2
23 0 9 9 1 9 13 1 12 5 1 1 0 9 9 7 9 0 9 1 0 15 9 2
1 9
7 1 9 1 11 15 13 13
6 11 11 2 0 0 9
22 11 13 1 0 9 1 9 12 0 9 2 15 13 2 16 0 13 7 9 13 0 2
8 15 7 13 9 1 10 9 2
19 1 9 9 13 3 0 2 16 0 0 9 13 0 13 1 9 1 9 2
14 1 9 15 13 3 7 13 1 15 13 7 0 9 2
41 3 0 9 2 3 1 9 14 12 9 2 13 0 0 9 2 9 1 9 0 9 2 9 2 0 9 2 0 9 3 2 2 7 0 0 9 15 3 3 13 2
19 9 13 1 9 12 9 2 12 0 9 2 2 7 0 9 13 3 0 2
31 3 15 10 9 13 1 14 9 9 2 7 9 9 13 3 9 2 16 15 2 15 13 13 3 16 9 2 3 9 13 2
17 13 0 15 0 9 13 1 9 9 2 7 7 13 13 1 9 2
15 1 9 0 0 9 13 0 15 13 9 0 9 7 9 2
13 10 9 13 3 12 0 9 0 9 1 12 9 2
35 15 15 13 1 9 1 12 9 2 16 0 9 13 12 9 2 12 9 7 0 12 9 2 2 7 13 15 3 0 0 9 2 3 0 2
19 1 9 9 3 13 13 2 16 15 13 15 0 2 15 3 13 9 0 2
32 9 10 12 7 0 9 13 1 0 9 2 1 0 7 3 7 1 0 9 2 3 1 10 0 0 9 7 1 0 9 11 2
28 9 0 9 0 9 7 9 2 3 0 1 0 2 7 0 9 2 13 1 10 0 12 7 0 9 0 9 2
43 3 3 13 9 1 9 2 15 1 9 0 9 2 1 0 9 7 1 0 9 13 1 0 9 13 2 0 0 9 7 9 2 16 14 1 9 2 3 3 1 0 9 2
12 1 9 0 15 9 1 0 1 15 13 9 2
13 3 0 13 9 9 9 2 15 13 3 12 9 2
16 0 0 9 13 12 9 2 7 7 0 9 3 13 12 9 2
17 10 9 13 1 15 0 16 9 1 9 3 0 9 1 0 9 2
15 7 7 9 13 9 2 7 15 13 15 1 0 13 9 2
22 13 15 2 15 3 13 2 14 16 4 15 13 9 2 0 13 13 13 1 0 9 2
5 10 9 13 0 2
21 13 3 1 9 1 9 1 9 2 0 9 15 13 9 9 2 9 7 0 9 2
17 3 1 9 9 15 0 0 9 13 9 1 9 0 9 7 9 2
55 7 3 13 9 1 9 9 2 0 9 2 0 9 2 9 1 3 0 2 0 9 2 0 9 9 2 0 9 1 0 7 0 2 9 1 0 9 7 9 2 10 9 15 1 11 13 1 3 12 12 2 7 0 9 2
16 9 1 15 13 0 13 3 0 9 2 15 14 13 10 9 2
14 9 0 1 10 9 13 1 9 0 0 9 3 0 2
26 15 2 15 13 13 1 9 2 15 13 13 3 1 9 0 9 2 3 13 3 0 9 0 9 9 2
12 9 13 2 16 0 1 10 9 13 0 9 2
22 3 13 2 16 15 2 15 13 12 9 9 2 13 13 0 2 7 16 4 15 13 2
14 10 9 4 13 3 1 0 9 2 7 7 1 9 2
25 0 9 13 0 9 9 2 16 10 9 2 7 15 14 0 7 0 9 2 13 9 1 0 9 2
45 9 10 9 13 9 12 9 9 2 12 9 9 2 2 7 3 1 9 10 2 9 2 13 3 1 9 0 9 9 12 9 9 2 12 9 9 2 2 15 4 13 1 0 9 2
53 0 9 2 15 15 13 1 9 0 9 2 1 9 12 2 12 0 13 2 3 1 9 2 1 10 9 3 0 9 2 7 9 9 1 0 9 13 1 9 14 1 12 7 12 9 1 9 9 2 1 9 12 2
33 0 9 13 7 0 9 2 16 0 9 13 1 0 9 1 9 1 10 9 2 16 4 3 13 10 9 7 13 0 9 0 9 2
8 9 13 3 0 1 15 0 2
44 3 1 9 0 9 13 9 2 15 3 13 2 13 1 9 1 9 10 12 9 2 7 16 13 9 9 0 2 16 9 9 1 12 9 7 1 9 3 0 13 10 9 13 2
32 1 9 9 13 0 9 3 0 9 2 15 13 1 9 16 12 1 10 0 9 13 0 9 2 16 4 13 3 10 0 9 2
25 1 15 13 13 1 9 0 9 0 9 2 9 1 9 7 0 9 9 2 3 9 1 0 9 2
18 3 13 15 0 2 13 0 9 2 16 15 13 1 9 11 1 11 2
9 7 3 3 13 13 9 0 9 2
17 13 2 16 15 13 9 0 1 9 2 1 9 2 1 9 9 2
24 1 0 9 13 13 2 1 9 12 13 1 9 9 12 3 0 2 1 9 12 3 14 12 2
15 1 9 12 1 9 9 13 12 7 1 9 12 3 12 2
16 9 9 13 2 16 1 9 9 9 13 14 1 9 9 9 2
19 13 0 2 16 1 9 0 11 15 3 1 11 3 13 9 9 0 9 2
33 1 11 15 9 13 12 9 2 1 11 12 2 1 11 1 12 9 1 9 12 1 9 12 15 13 0 9 1 12 1 12 9 2
17 9 13 12 9 9 0 1 9 1 12 2 12 9 16 1 9 2
14 13 15 2 9 9 1 9 9 2 0 9 7 9 2
22 1 9 12 3 13 10 9 12 9 2 1 9 12 3 12 9 7 1 0 9 12 2
13 1 0 9 11 11 13 1 0 9 12 0 9 2
17 0 9 3 13 2 16 0 9 15 3 13 1 9 16 1 9 2
20 11 13 9 0 1 0 9 0 11 2 1 15 15 3 1 9 9 13 9 2
8 0 9 13 9 1 9 9 2
22 1 9 12 15 9 9 1 9 0 9 7 9 13 0 9 13 1 12 2 12 5 2
10 0 0 9 13 0 9 3 9 9 2
8 1 9 12 9 13 12 9 2
26 9 13 15 2 15 4 13 7 1 15 2 16 15 3 15 9 13 1 0 9 2 15 0 9 13 2
21 1 0 9 4 13 9 9 7 3 9 0 9 9 9 1 0 9 9 1 9 2
58 0 9 13 2 16 1 9 2 1 15 13 0 9 2 13 0 13 1 9 0 9 2 9 0 7 0 2 1 9 0 2 1 0 9 2 1 9 1 9 7 9 2 1 9 0 9 2 0 9 7 0 9 2 1 0 9 9 2
34 1 11 13 9 9 1 9 0 7 0 9 0 16 1 10 0 0 9 2 9 15 13 0 9 7 9 9 15 13 1 0 1 11 2
23 13 13 2 16 7 1 0 9 13 0 9 13 0 9 1 9 7 15 7 9 1 9 2
25 13 0 13 9 1 9 7 0 9 2 7 9 7 9 1 0 9 9 13 9 1 9 1 9 2
17 15 13 9 2 15 13 9 7 9 2 1 15 15 13 1 9 2
22 9 13 13 1 9 9 2 9 13 9 2 13 0 9 1 9 7 13 1 9 9 2
31 16 15 1 9 0 9 0 9 13 3 2 0 9 9 15 10 9 13 7 13 15 9 9 2 13 15 7 9 1 9 2
24 7 16 15 10 9 13 13 2 13 13 1 15 2 16 4 15 1 9 10 9 4 13 9 2
30 15 2 15 3 13 1 9 2 13 0 2 0 7 3 13 1 9 1 0 9 15 0 7 0 2 15 3 15 13 2
2 11 11
3 9 1 11
27 1 9 0 9 0 9 13 0 9 11 11 9 9 2 13 11 1 9 1 10 2 15 15 15 11 13 2
8 1 9 7 13 0 9 11 2
42 9 0 9 13 1 0 0 9 9 2 16 1 11 4 0 9 13 1 9 0 1 9 9 2 7 0 9 13 1 9 12 1 0 9 9 7 13 0 11 1 9 2
23 11 7 10 0 0 9 15 13 1 9 1 9 2 15 13 1 9 10 9 7 9 9 2
11 9 15 1 9 1 9 13 1 15 13 2
14 13 7 0 9 2 16 4 9 13 3 1 10 9 2
18 15 9 7 9 2 14 1 12 2 1 0 0 9 13 12 9 0 2
20 14 1 9 0 9 7 9 15 9 13 1 3 0 2 7 16 3 0 9 2
20 9 7 3 13 9 10 9 0 1 12 9 2 3 13 4 1 9 9 13 2
23 1 11 15 1 9 0 9 1 9 9 13 15 2 16 13 1 9 9 0 9 11 0 2
10 0 0 9 11 11 13 1 10 9 2
19 1 0 9 11 0 1 9 0 9 13 11 1 9 1 9 1 0 9 2
19 0 9 2 10 9 13 13 14 1 9 2 13 9 11 11 9 0 9 2
10 11 13 9 0 9 3 1 9 9 2
23 1 0 9 11 3 2 13 9 0 0 9 9 2 9 9 2 12 7 9 0 9 11 2
23 1 11 4 13 1 9 2 7 13 15 3 12 9 2 1 9 12 4 13 1 0 9 2
17 0 9 1 11 13 2 16 4 9 11 13 11 13 9 1 11 2
19 15 13 7 9 11 11 2 16 9 9 13 2 16 4 0 9 9 13 2
8 1 12 9 9 11 13 15 2
29 13 9 4 12 9 0 9 1 9 9 11 11 7 11 11 2 0 2 16 1 9 12 13 9 0 9 11 11 2
11 9 13 2 16 13 0 9 1 9 9 2
20 9 2 15 13 1 0 1 9 9 12 9 9 2 13 1 9 1 0 9 2
33 9 12 12 9 9 15 1 10 9 3 13 9 0 0 9 11 11 2 7 10 9 11 11 2 15 1 9 1 9 13 12 9 2
3 9 1 11
22 0 9 15 13 13 1 9 0 9 1 9 12 2 16 15 4 15 13 3 0 9 2
25 1 0 9 11 12 15 13 11 1 11 3 1 9 0 9 2 9 11 7 1 9 10 9 13 2
12 0 3 0 9 3 13 0 9 3 0 9 2
9 0 9 13 13 1 9 1 9 2
20 0 0 9 4 1 11 13 3 1 9 2 16 11 13 0 9 1 9 9 2
15 13 15 0 9 9 11 11 2 9 0 9 0 9 9 2
33 9 1 0 0 9 7 0 9 13 1 11 10 9 2 16 0 9 13 1 9 10 9 7 9 13 3 13 9 7 9 0 9 2
12 9 13 10 9 2 4 7 13 13 9 11 2
12 3 15 13 2 16 9 13 12 7 12 9 2
25 0 0 9 13 9 1 12 9 1 0 9 2 16 4 13 9 9 7 13 10 9 1 0 9 2
14 0 3 0 9 13 1 0 9 9 1 9 7 9 2
20 0 0 9 1 0 9 0 9 13 12 9 2 15 2 13 2 3 12 9 2
13 13 15 1 12 5 3 16 1 0 9 0 9 2
13 9 0 9 3 1 0 9 13 14 1 12 5 2
34 11 13 0 13 1 0 9 9 0 9 7 13 15 2 16 4 13 1 11 10 0 9 2 13 1 10 0 9 11 9 9 11 11 2
12 0 0 9 1 11 13 0 13 11 0 9 2
17 1 9 7 11 13 2 16 4 11 13 9 0 9 1 10 9 2
17 9 0 9 11 13 3 12 1 12 0 0 9 13 1 11 9 2
28 11 3 13 1 11 9 1 9 9 2 15 3 13 0 9 2 15 15 11 3 13 16 9 9 15 12 9 2
22 11 11 15 1 10 9 13 1 9 0 1 0 11 2 13 0 9 11 11 9 11 2
36 0 9 9 13 7 13 2 16 15 13 3 3 2 11 14 13 11 2 16 4 15 13 1 9 0 11 7 1 9 10 9 1 9 0 9 2
23 9 0 9 3 13 9 0 9 2 1 10 9 7 13 9 2 1 15 10 0 9 13 2
25 1 9 2 16 4 15 11 13 11 2 13 9 11 11 11 11 2 3 0 9 7 9 0 9 2
21 1 11 13 11 10 9 0 1 9 11 15 11 2 7 13 1 11 9 0 9 2
10 11 11 15 13 1 0 9 0 9 2
17 13 15 15 2 16 9 9 15 13 13 3 1 9 0 1 9 2
30 9 0 9 2 0 9 0 0 9 2 3 13 7 13 1 15 2 16 1 0 0 9 13 10 9 1 9 1 9 2
15 1 0 9 13 1 0 9 0 3 15 13 1 0 9 2
15 0 3 0 9 13 1 10 9 0 9 1 9 0 9 2
11 1 9 0 9 7 4 13 10 9 13 2
34 1 0 9 0 9 13 0 9 9 9 0 9 2 15 15 1 0 9 13 1 9 1 9 13 9 0 0 9 1 10 9 1 11 2
5 9 4 3 13 2
11 9 0 9 13 9 1 0 9 1 11 2
15 9 0 0 9 4 13 1 0 9 1 11 1 0 9 2
16 9 13 10 9 2 16 9 15 13 1 0 9 1 9 11 2
13 13 7 13 2 16 15 3 13 7 1 9 11 2
20 12 1 0 9 12 2 0 9 1 0 11 13 3 9 0 9 0 1 9 2
16 9 9 3 13 0 9 2 16 4 13 9 3 1 9 11 2
19 11 11 1 10 0 9 11 11 11 13 1 0 9 11 2 3 13 9 2
4 9 0 0 9
1 11
5 11 11 2 11 0
42 3 1 0 11 1 0 11 7 1 3 0 0 9 9 2 1 0 9 1 15 3 16 0 0 0 9 15 13 1 9 9 1 0 11 0 9 2 9 0 0 9 2
45 0 9 0 9 0 9 13 3 1 0 0 9 0 9 2 9 7 9 2 16 4 0 9 0 0 9 1 9 0 11 1 11 7 11 13 10 9 1 15 2 15 15 3 9 13
7 9 1 9 13 0 9 2
28 9 0 9 11 11 7 9 0 9 11 11 2 0 1 10 9 2 7 3 3 13 2 15 15 13 1 11 2
33 11 3 13 2 16 1 9 0 9 9 13 13 2 9 7 9 15 4 13 1 9 1 9 9 2 7 1 0 9 9 13 9 2
13 15 7 13 0 2 13 0 9 9 1 9 0 2
22 7 3 0 2 13 15 9 15 2 15 15 9 13 2 7 15 2 15 15 13 13 2
36 12 9 11 1 9 9 13 0 9 2 14 2 14 0 9 2 3 1 9 1 0 9 0 9 11 2 0 9 7 3 1 0 9 1 9 2
20 0 0 9 13 15 9 9 2 15 1 10 3 0 9 0 9 13 9 11 2
19 9 7 1 15 0 0 0 9 15 3 13 2 16 9 9 13 3 3 2
27 9 1 9 4 13 3 9 9 2 3 3 9 0 9 2 7 13 4 2 16 11 13 0 9 3 3 2
12 9 4 13 7 13 15 10 2 7 15 9 2
15 9 9 7 9 1 9 13 2 7 4 15 13 3 0 2
30 13 15 2 1 9 11 2 15 2 15 0 9 2 9 9 2 9 7 9 2 15 13 0 9 1 0 9 7 9 2
22 16 13 2 13 15 0 9 10 0 3 0 9 2 1 0 0 9 4 13 0 9 2
6 11 13 7 0 9 2
25 4 13 3 9 0 0 9 2 13 7 3 2 3 15 4 0 9 9 13 1 10 0 0 9 2
21 9 2 9 9 1 12 9 13 3 0 2 3 0 2 15 15 4 3 13 13 2
42 11 2 11 7 10 0 9 11 11 13 2 16 0 9 15 13 3 1 0 9 7 16 7 0 9 13 3 2 3 13 0 0 9 2 13 3 0 9 1 0 9 2
2 9 9
12 9 9 11 13 1 9 7 1 12 9 9 2
33 11 13 9 9 2 13 12 0 9 1 9 9 9 2 7 3 13 1 9 0 9 9 1 0 9 1 12 1 15 2 1 11 2
29 0 9 0 9 13 15 7 0 7 0 9 11 1 9 13 3 15 13 2 16 4 13 9 0 0 9 0 9 2
24 0 7 0 0 9 1 11 11 11 2 3 9 0 9 1 0 9 2 13 1 0 9 9 2
40 11 13 0 9 1 0 9 2 7 7 13 1 15 0 14 1 9 3 0 2 2 0 9 13 3 1 0 9 0 2 15 3 13 1 10 9 0 0 9 2
31 11 3 3 13 2 16 0 9 13 13 0 13 1 0 7 0 9 2 15 13 1 0 9 3 0 1 9 1 0 9 2
11 15 13 3 0 9 0 9 1 0 11 2
11 13 15 3 13 2 7 14 13 0 9 2
18 9 0 9 1 11 11 11 15 13 0 2 7 3 0 2 9 11 2
38 7 9 2 7 11 0 7 0 11 1 9 13 13 2 13 15 16 9 2 16 15 2 1 15 13 10 9 2 7 14 16 9 1 15 7 0 11 2
3 9 0 9
10 0 11 15 3 3 13 1 10 9 2
17 3 0 9 1 0 9 7 1 11 13 13 10 9 1 9 9 2
16 9 11 1 9 0 9 2 15 4 13 9 0 9 0 11 2
11 13 15 1 0 11 2 7 15 3 13 2
5 2 11 2 2 2
10 9 1 0 9 0 9 13 3 3 2
12 3 13 11 11 2 7 1 11 9 13 9 2
14 16 4 15 13 9 2 9 4 15 13 9 0 9 2
10 1 11 13 9 2 14 9 2 9 2
22 9 9 7 9 2 13 3 1 11 0 0 9 11 11 1 15 2 15 11 0 13 2
8 15 15 13 2 13 0 9 2
11 13 15 15 2 1 9 9 2 13 3 2
12 0 9 0 9 15 1 15 13 9 0 9 2
14 11 3 13 2 7 13 13 0 9 2 11 2 2 2
2 9 9
11 11 13 3 1 3 0 11 3 0 9 2
18 0 0 9 2 0 0 9 7 0 0 9 13 1 15 3 0 9 2
31 3 15 7 13 15 1 11 13 3 0 9 9 7 0 9 1 0 9 2 15 13 3 3 9 0 9 3 1 0 11 2
14 13 4 15 2 16 11 4 13 10 9 1 0 9 2
42 9 7 1 9 0 2 0 7 3 7 0 9 9 13 9 2 9 13 0 0 9 7 0 9 2 7 0 9 0 0 9 7 0 11 4 13 16 9 10 0 9 2
29 9 0 0 9 13 0 9 2 9 2 9 9 2 3 3 2 0 9 11 11 11 2 3 0 9 1 11 2 2
21 13 3 9 2 16 15 1 15 11 13 3 3 16 15 1 15 7 13 13 3 2
13 0 11 13 13 0 9 2 16 9 13 1 0 2
20 7 1 0 9 15 1 15 7 0 11 3 13 15 2 1 15 3 13 9 2
9 0 9 1 9 2 7 1 9 2
1 11
2 11 11
2 11 0
19 1 9 13 9 11 0 0 9 2 9 2 0 9 0 2 0 9 11 2
16 9 15 3 3 13 1 0 9 0 11 2 15 13 1 9 2
7 0 9 11 7 9 13 2
21 9 2 0 10 9 9 2 0 1 9 9 11 11 2 13 3 16 9 12 9 2
18 13 15 12 1 0 9 9 11 11 11 7 13 15 0 9 9 9 2
13 1 9 13 9 2 0 1 0 9 9 1 9 2
14 1 9 15 13 9 11 2 15 1 9 15 9 13 2
16 9 1 9 13 1 0 9 7 3 13 1 9 1 9 11 2
17 9 13 0 9 1 0 9 2 3 13 13 1 3 0 0 9 2
4 9 1 9 13
24 9 1 9 1 9 7 9 1 9 2 15 13 1 9 1 9 12 2 3 13 9 1 9 2
6 1 9 15 7 13 2
18 9 13 9 2 13 9 1 9 9 2 13 11 11 1 9 11 11 2
27 1 10 9 13 9 2 15 13 11 11 2 3 0 9 1 9 2 13 9 0 9 0 9 11 11 11 2
21 11 13 11 11 1 0 9 1 9 9 7 9 7 1 0 9 1 9 1 9 2
12 1 9 10 9 15 3 3 9 13 1 9 2
22 13 13 2 16 13 1 10 9 3 0 9 9 2 13 11 11 1 9 9 0 9 2
7 3 4 1 10 9 13 2
9 1 10 9 15 13 1 9 13 2
18 13 9 2 7 13 1 9 0 9 2 13 9 9 0 9 11 11 2
14 11 11 13 1 0 9 9 11 1 0 9 0 9 2
18 15 15 7 1 9 1 9 2 15 15 4 3 13 2 13 13 9 2
17 1 0 0 9 13 0 9 2 15 15 13 3 2 0 9 11 2
5 11 13 9 11 2
15 0 9 1 9 1 15 13 7 9 1 9 9 9 13 2
2 0 9
43 3 13 1 11 13 2 16 15 13 9 1 9 2 7 3 15 1 10 0 9 13 13 0 9 2 16 11 11 13 9 1 9 11 2 13 15 11 11 1 9 11 11 2
11 13 1 0 9 1 0 9 9 11 11 2
16 13 1 15 3 2 13 0 9 1 9 2 0 9 7 9 2
26 15 9 9 13 2 7 16 15 13 13 2 16 1 9 3 13 9 1 9 7 1 9 2 13 11 2
13 1 0 9 15 13 1 9 9 2 13 11 11 2
14 9 1 9 1 9 7 9 13 3 7 1 11 0 2
3 9 1 11
18 0 0 9 12 2 9 7 12 2 9 15 13 12 0 9 7 9 2
21 1 12 0 9 1 0 9 0 9 15 4 13 12 9 2 1 15 12 9 2 2
7 0 9 9 13 12 9 2
19 3 9 2 12 2 13 9 1 0 11 2 3 2 14 12 2 9 9 2
17 1 0 9 0 9 0 9 13 15 1 9 13 3 12 0 9 2
7 11 13 0 9 11 11 2
10 13 1 9 11 11 7 9 11 11 2
27 1 10 9 12 9 13 0 9 2 9 1 9 0 9 2 9 1 0 9 7 9 1 9 0 0 9 2
32 9 0 9 2 0 9 0 0 9 7 0 0 0 9 13 0 9 1 0 9 0 1 0 9 0 0 9 1 9 0 9 2
31 1 9 15 13 9 0 0 9 2 0 9 2 15 15 1 9 0 0 9 13 1 9 0 9 7 9 9 11 2 11 2
26 0 9 11 13 13 2 16 9 0 9 13 1 9 9 1 0 9 2 15 13 9 9 0 0 9 2
8 9 9 13 1 0 9 11 2
22 1 10 9 3 13 3 16 12 9 2 1 15 1 12 9 1 9 1 12 9 2 2
10 0 12 9 13 9 1 0 9 11 2
17 1 9 13 9 9 9 0 1 9 0 9 1 12 1 0 9 2
36 1 0 9 11 13 9 9 11 11 11 9 9 0 11 11 2 1 15 13 3 11 1 9 0 11 1 9 12 2 12 9 1 12 9 9 2
18 1 11 2 11 0 9 3 13 9 11 0 9 9 1 9 0 11 2
34 16 13 9 0 0 9 11 1 9 9 2 13 0 9 11 11 13 1 0 2 0 9 2 15 15 4 13 1 9 10 9 1 9 2
16 1 10 9 15 13 0 9 7 0 9 15 15 13 13 15 2
21 0 9 15 13 15 2 16 1 9 10 9 4 13 9 2 7 0 9 9 11 2
24 0 9 9 7 0 9 0 9 9 13 0 9 1 11 13 9 9 1 0 9 1 9 9 2
16 3 1 9 9 4 3 1 0 9 13 12 9 0 0 9 2
12 9 9 15 7 13 1 9 1 0 0 9 2
47 9 0 0 0 0 9 9 11 11 2 0 1 9 9 12 0 9 1 11 1 12 9 9 1 9 0 9 1 9 0 9 2 3 3 13 9 9 1 0 9 2 3 13 1 9 11 2
25 16 11 13 13 9 9 1 11 2 4 1 9 9 11 11 11 0 9 13 10 9 1 15 9 2
8 1 11 13 9 3 0 9 2
15 13 15 13 1 9 9 0 0 9 9 1 9 9 9 2
33 1 9 9 4 9 1 0 9 1 9 13 1 0 7 0 9 2 1 9 0 9 1 10 9 7 9 9 9 1 9 0 9 2
19 1 0 9 4 3 13 0 9 2 13 15 10 0 9 2 9 7 9 2
3 9 1 9
1 11
28 1 9 11 13 9 2 3 0 9 1 9 1 9 2 1 0 9 0 7 0 9 7 1 9 1 9 9 2
11 13 3 7 3 13 0 9 2 13 15 2
30 15 3 2 16 9 3 13 2 3 9 1 12 2 9 1 12 7 9 1 9 12 9 2 15 13 1 0 11 0 2
28 1 9 1 0 0 9 2 1 9 11 9 9 2 12 2 15 3 13 9 9 2 12 7 9 9 2 12 2
4 9 1 9 2
1 11
27 0 0 9 1 11 2 15 15 4 1 10 0 9 13 12 2 7 12 2 9 2 13 3 0 1 9 2
8 9 9 13 13 9 0 11 2
20 9 9 13 13 3 0 9 9 11 11 11 11 2 15 13 1 10 0 9 2
9 1 9 11 2 12 13 9 3 2
25 13 15 13 1 0 9 1 0 9 2 3 9 9 9 2 12 7 9 9 2 12 1 9 11 2
3 2 11 2
4 0 9 13 11
12 9 1 0 9 11 11 2 9 0 9 1 9
5 11 11 2 0 9
18 1 11 13 9 9 0 9 1 9 0 9 3 1 9 12 2 9 2
21 0 9 13 10 9 13 9 11 11 10 0 9 9 11 2 15 13 0 9 11 2
30 11 1 10 9 0 9 13 3 7 3 1 10 9 9 9 2 15 9 7 9 13 1 15 1 15 0 9 11 0 2
9 1 11 13 1 11 15 0 9 2
34 7 16 1 11 0 13 0 9 0 9 0 0 2 0 9 2 0 9 11 3 13 9 9 9 2 16 4 9 10 0 9 3 13 2
22 15 15 13 1 15 2 16 4 15 10 9 13 2 7 15 1 10 9 13 1 0 2
9 3 3 16 11 13 11 0 9 2
7 16 13 11 10 0 9 2
21 0 13 2 16 4 1 9 11 13 3 16 1 11 2 15 3 13 9 0 9 2
6 10 9 3 3 13 2
19 1 9 4 15 13 7 3 2 16 0 9 13 13 1 9 9 0 9 2
17 9 1 3 0 0 0 9 2 0 7 3 0 9 13 0 11 2
17 1 15 4 15 9 0 9 0 9 0 11 13 1 3 0 9 2
14 7 13 2 16 1 0 9 4 4 13 7 9 0 2
7 15 11 1 9 12 13 2
11 13 3 7 1 0 9 9 9 0 9 2
24 15 15 13 1 9 0 9 1 9 2 15 13 7 9 12 2 16 3 9 9 9 7 9 2
19 15 13 2 16 0 7 0 9 13 15 0 2 15 13 2 16 13 0 2
10 13 4 15 13 3 1 9 7 9 2
11 13 4 7 9 2 1 15 13 9 13 2
30 3 0 0 9 0 0 9 11 11 2 1 15 13 3 2 16 11 13 9 1 15 2 16 13 1 11 12 0 9 2
15 16 4 15 1 10 9 13 13 1 11 3 0 7 0 2
31 13 11 7 1 9 1 0 9 2 3 15 0 9 2 0 9 2 14 0 9 3 7 13 2 15 1 9 3 13 3 2
22 1 9 13 2 16 0 9 2 15 15 13 1 0 9 2 13 1 9 11 3 0 2
19 0 9 2 15 9 11 13 1 0 2 13 1 9 11 0 2 3 3 2
24 9 0 13 1 0 9 2 16 1 9 0 9 13 3 0 13 9 16 0 9 7 0 9 2
14 9 9 0 9 13 1 9 0 11 0 3 3 3 2
11 0 9 13 3 0 2 3 3 16 0 2
47 3 13 1 11 1 9 2 1 15 1 15 9 3 13 3 2 16 15 2 15 3 11 1 9 13 1 0 0 9 7 1 0 2 0 9 2 1 15 11 13 1 0 9 2 13 9 2
41 9 3 13 12 0 9 2 12 1 15 13 11 11 2 9 0 9 2 15 13 10 9 1 9 2 3 9 0 9 2 7 1 9 4 15 7 13 3 13 2 2
17 1 3 3 0 13 9 1 12 2 9 2 13 15 10 9 2 2
15 13 15 0 9 2 7 1 9 9 13 10 9 3 0 2
7 0 9 13 1 0 9 2
8 3 0 13 9 9 1 11 2
13 0 15 13 2 16 13 1 9 3 0 9 9 2
32 0 13 2 15 15 13 1 0 0 9 2 15 3 1 0 0 0 9 13 15 13 2 16 4 15 7 13 9 0 9 2 2
8 13 10 0 9 1 0 9 2
16 14 2 9 1 9 13 9 3 1 9 1 0 2 0 9 2
23 0 9 1 11 7 1 11 13 3 3 15 2 16 1 9 13 0 9 7 0 10 9 2
10 3 4 9 9 13 1 9 14 3 2
5 15 13 0 9 2
19 13 4 1 9 9 0 9 2 1 15 4 3 1 0 9 13 9 2 2
16 0 9 4 3 13 2 16 4 15 1 15 3 13 0 9 2
11 1 10 0 9 4 15 3 13 9 9 2
7 15 13 9 1 9 11 2
8 12 9 9 0 9 13 13 2
4 13 0 9 2
31 10 0 9 13 13 0 9 1 11 2 15 3 13 2 16 4 1 9 13 2 16 4 1 15 13 1 9 9 9 9 2
27 13 4 15 3 9 2 16 4 9 13 1 9 0 2 0 2 1 0 9 0 2 7 14 0 0 9 2
6 9 13 7 0 11 2
11 7 15 13 0 2 0 9 1 10 9 2
4 9 15 3 13
13 1 0 9 13 1 0 9 9 9 7 9 0 9
5 11 11 2 11 0
21 0 0 9 1 0 9 13 1 9 7 1 0 9 9 3 3 2 16 13 13 2
7 13 9 2 9 7 9 2
11 7 3 15 9 13 7 1 9 0 9 2
15 3 0 9 15 13 9 13 0 9 7 13 1 10 9 2
11 1 0 9 9 9 7 9 13 0 9 2
18 9 0 9 7 9 0 0 9 15 13 13 1 9 14 1 12 9 2
3 9 13 3
14 16 9 13 2 9 15 13 0 9 2 9 13 9 2
4 15 15 13 2
16 3 15 13 2 2 13 15 9 1 9 1 0 9 1 11 2
8 9 9 1 9 13 10 9 2
19 0 9 13 9 1 9 0 2 13 3 12 7 12 2 7 12 12 9 2
7 15 1 9 15 3 13 2
11 9 13 3 2 13 9 9 1 0 9 2
11 0 9 1 9 9 4 13 12 9 9 2
7 3 15 13 3 12 9 2
11 13 4 15 2 16 0 9 13 1 9 2
15 7 1 0 9 9 15 9 7 9 3 13 1 0 9 2
8 0 9 13 3 2 7 13 2
16 1 0 9 1 0 9 15 13 2 16 9 7 9 13 4 2
11 0 14 13 13 15 7 13 9 0 9 2
7 0 9 3 10 9 13 2
22 1 9 11 11 1 0 9 11 2 0 9 9 0 9 2 7 9 3 13 10 9 2
18 13 2 16 13 3 1 9 0 9 2 7 13 15 3 3 2 13 2
36 13 15 9 7 9 1 0 11 7 13 15 2 13 2 14 4 1 9 0 9 13 2 3 13 13 9 1 0 9 2 15 13 1 0 9 2
3 9 1 9
33 13 2 16 9 9 13 2 7 16 15 2 1 9 13 2 3 13 2 13 11 11 1 0 9 11 0 11 2 9 7 9 2 2
20 0 9 9 4 13 9 1 9 3 10 9 2 7 9 15 1 15 13 13 2
8 0 9 1 9 13 3 13 2
17 9 13 1 9 2 16 13 15 1 9 9 1 0 9 7 9 2
20 13 0 15 13 1 9 2 16 13 9 7 13 1 15 3 12 7 12 9 2
11 16 0 9 13 9 9 3 3 16 0 2
12 3 13 1 15 9 7 1 15 3 9 13 2
4 9 7 9 2
10 0 9 9 0 9 13 9 9 9 2
15 13 15 9 3 0 2 9 13 1 0 11 14 1 12 2
6 13 15 7 3 9 2
9 1 9 9 7 13 0 0 9 2
29 1 9 11 11 1 11 2 15 1 0 9 13 9 11 2 3 13 9 9 1 9 2 15 15 1 11 3 13 2
14 11 11 13 1 10 9 1 9 1 11 1 12 9 2
8 1 9 9 4 13 0 9 2
17 1 11 13 9 0 2 15 15 3 13 9 1 12 2 12 9 2
7 9 9 15 15 13 13 2
11 13 15 1 0 9 2 3 1 9 2 2
25 13 9 7 13 13 13 1 9 7 9 1 9 1 9 10 9 2 13 9 0 9 11 11 11 2
9 7 15 1 0 1 15 3 13 2
18 9 2 15 13 13 0 0 9 7 13 1 15 9 2 15 3 13 2
15 9 13 0 9 9 0 9 2 1 10 9 13 11 11 2
18 3 13 7 1 10 9 14 10 9 9 2 13 1 15 3 0 9 2
19 9 9 9 2 9 13 9 10 0 9 9 1 9 9 9 2 11 2 2
7 15 7 3 13 10 9 2
19 11 11 13 2 16 9 13 9 1 0 9 0 9 2 9 9 7 9 2
3 3 9 9
29 1 9 2 3 9 13 13 2 4 13 12 9 2 13 0 9 2 9 1 9 0 9 2 15 15 13 4 13 2
22 10 9 15 13 13 2 3 3 13 0 0 9 2 1 0 9 7 13 9 2 13 2
8 9 1 9 13 3 1 9 2
25 16 15 13 1 0 0 9 9 9 1 0 9 0 9 2 13 4 13 1 9 9 1 10 9 2
23 9 0 9 11 2 10 9 13 9 11 2 7 0 2 9 15 1 10 9 13 3 3 2
16 0 2 9 13 0 9 1 0 9 2 9 1 12 2 9 2
4 9 2 9 11
1 3
17 0 0 9 11 15 13 13 0 9 1 0 9 1 0 0 9 2
17 0 9 2 0 0 0 11 2 0 2 2 13 13 1 0 9 2
12 0 9 4 13 13 1 0 9 3 0 0 2
6 13 15 9 10 9 2
16 11 13 7 1 0 9 0 9 0 9 9 9 1 10 9 2
23 9 15 13 1 0 1 0 9 0 9 7 1 10 3 15 0 9 1 0 7 0 9 2
8 9 11 3 13 1 12 9 2
3 9 1 9
2 11 2
22 0 9 0 0 9 13 9 9 12 9 9 2 1 15 9 0 0 9 13 12 9 2
19 9 0 0 9 13 1 9 1 12 9 2 1 9 13 10 9 12 9 2
18 9 11 15 1 9 13 1 12 9 2 1 9 15 13 9 12 9 2
15 0 9 0 9 1 0 9 13 1 9 9 12 9 9 2
11 13 15 9 1 9 9 7 9 0 9 2
26 1 9 9 15 13 1 12 2 3 2 12 9 2 1 9 9 15 13 12 2 3 2 12 9 2 2
31 3 15 13 0 0 9 2 7 15 0 1 0 12 1 12 9 2 0 1 12 1 12 9 7 0 1 12 1 12 9 2
9 1 11 15 4 1 9 0 9 13
2 11 2
26 0 9 9 0 0 9 1 11 11 1 9 13 9 0 7 0 9 2 0 1 0 9 1 10 9 2
6 3 15 13 9 11 2
21 1 15 13 11 1 10 0 9 1 9 9 1 9 1 0 9 7 3 10 9 2
16 1 0 9 0 9 4 9 0 9 1 0 9 11 11 13 2
9 9 13 3 7 13 12 5 9 2
16 1 9 0 0 9 9 15 9 13 7 13 9 0 0 9 2
38 1 1 15 2 16 0 9 1 9 7 9 13 9 2 16 0 9 13 13 0 9 9 2 13 9 11 3 1 9 9 0 9 1 9 9 1 0 2
18 0 9 15 13 2 16 9 13 3 1 9 0 0 9 2 13 11 2
6 9 0 9 13 9 9
7 11 2 11 2 11 2 2
42 9 0 9 1 10 0 9 12 2 9 3 13 2 16 13 1 0 2 16 4 4 9 9 2 10 9 4 3 1 9 0 9 13 2 13 0 9 3 1 9 9 2
8 13 15 3 9 9 11 11 2
18 1 11 2 11 13 10 9 0 9 9 7 13 3 1 9 0 9 2
15 9 10 9 3 13 1 9 2 15 13 13 3 0 9 2
10 9 13 12 1 12 0 9 0 9 2
12 10 9 13 3 9 0 9 7 0 0 9 2
25 9 7 3 13 10 9 2 15 3 3 13 2 3 1 9 9 9 9 1 0 9 7 0 9 2
5 0 9 13 1 9
9 9 9 1 0 9 13 0 7 0
5 11 2 11 2 2
20 1 0 9 1 0 9 3 12 9 13 0 9 0 7 0 9 2 9 2 2
36 9 0 9 2 1 15 15 9 13 1 0 11 2 13 1 9 0 9 9 11 11 7 9 0 9 12 9 2 15 13 3 9 9 10 9 2
10 9 9 1 12 9 4 13 0 9 2
24 0 9 13 9 0 7 0 9 2 3 13 1 9 0 9 1 15 13 12 5 9 9 9 2
21 3 13 9 9 9 2 1 15 13 1 9 12 7 12 9 2 9 1 9 9 2
16 1 1 9 12 9 2 9 13 10 9 1 11 2 11 0 2
9 9 0 9 1 0 9 13 0 2
13 3 0 9 0 9 1 9 9 13 1 12 9 2
17 9 2 15 13 9 1 0 9 2 13 0 9 1 12 12 9 2
13 3 7 9 13 1 0 9 2 0 9 13 0 2
44 1 0 11 3 13 9 10 9 2 1 15 7 13 13 9 2 1 15 15 3 13 3 1 9 1 12 9 2 9 2 2 16 1 9 13 9 1 9 1 12 9 2 9 2
27 1 0 9 0 9 1 0 9 13 3 0 0 9 13 2 7 11 2 11 15 13 2 16 13 15 3 2
33 0 9 1 9 0 1 11 2 15 13 1 9 2 9 3 2 2 13 12 7 12 9 2 9 2 12 7 12 9 2 9 2 2
8 13 3 12 9 15 13 9 2
9 15 13 1 9 15 7 0 9 2
12 13 15 9 0 9 9 2 13 11 2 11 2
21 15 0 9 2 11 2 11 3 2 2 9 13 7 13 15 3 1 9 2 13 2
15 1 10 9 13 0 9 9 1 9 0 1 0 9 11 2
19 15 4 13 13 12 0 9 2 7 0 3 12 7 12 9 1 9 9 2
11 9 13 13 0 0 9 3 1 0 9 2
14 9 1 0 9 4 13 4 13 9 9 7 0 9 2
30 1 9 0 9 0 0 9 2 15 13 0 9 1 9 2 11 2 11 13 2 16 3 10 9 13 9 1 0 9 2
15 9 9 13 7 0 10 9 13 3 2 13 15 13 9 2
24 9 2 15 13 1 9 9 2 4 1 0 9 1 9 13 7 1 0 9 9 1 0 9 2
8 0 9 13 1 10 0 9 0
6 11 11 2 0 9 11
22 9 1 0 9 13 1 15 13 0 9 9 7 3 0 9 9 13 1 0 0 9 2
14 9 3 13 3 0 7 9 13 14 1 0 0 9 2
9 9 13 13 3 1 9 0 9 2
17 0 9 1 9 0 9 3 13 9 1 0 9 9 1 0 9 2
11 0 9 13 3 9 9 9 0 0 9 2
51 16 13 9 15 2 9 4 13 13 2 16 3 13 9 2 3 13 1 9 7 0 9 10 9 13 0 9 16 1 0 9 2 7 7 16 3 14 13 3 1 0 9 2 15 3 13 13 1 0 9 2
4 0 13 12 2
12 0 9 9 1 9 9 9 3 3 15 13 2
18 0 9 3 3 13 2 16 9 2 10 9 13 2 13 9 7 3 2
18 1 9 2 3 4 9 13 1 9 2 15 13 7 9 0 0 9 2
12 9 13 1 15 0 15 1 9 13 3 3 2
13 15 2 15 3 13 9 1 9 2 13 13 0 2
17 13 15 1 9 3 1 9 7 0 9 2 15 3 10 9 13 2
7 11 9 13 13 3 0 9
2 11 2
21 1 12 0 9 1 0 9 7 1 11 13 13 0 9 11 9 1 9 1 11 2
10 1 9 0 11 13 13 1 9 12 2
18 3 13 13 1 12 0 9 2 1 15 12 1 11 7 12 1 11 2
16 1 0 9 13 9 0 9 2 7 15 9 13 9 0 9 2
33 16 13 1 0 0 9 1 11 0 9 11 9 11 11 2 1 9 9 1 9 0 9 13 9 1 0 9 0 9 9 9 11 2
10 15 9 1 0 9 9 1 11 13 2
9 1 0 9 13 9 1 0 9 2
11 0 9 4 13 13 9 1 9 0 9 2
14 11 9 3 13 1 9 9 1 9 9 1 9 11 2
14 9 1 10 9 13 7 0 9 2 1 15 9 13 2
7 0 9 4 13 9 11 2
11 0 9 11 9 13 9 0 9 1 9 2
8 0 9 13 9 0 0 9 2
12 0 0 9 7 13 10 9 14 1 0 9 2
9 3 1 15 7 4 13 0 9 2
19 1 9 13 14 9 9 2 3 11 9 13 9 0 0 9 12 2 9 2
4 11 3 13 9
16 0 0 9 11 11 11 13 9 10 9 1 0 9 10 9 2
25 9 0 9 15 1 9 1 0 9 0 9 13 1 12 5 2 1 12 9 2 9 1 12 9 2
12 13 1 0 9 2 10 9 13 3 12 5 2
22 13 15 3 9 2 7 16 3 3 2 7 15 1 12 9 2 9 1 0 12 9 2
23 10 9 13 9 2 16 15 0 9 1 11 3 13 7 13 9 2 3 1 0 9 11 2
7 9 1 0 9 3 13 2
13 0 9 11 3 3 13 13 9 0 9 1 11 2
21 1 15 0 9 9 2 1 0 7 1 9 0 7 0 11 2 15 9 11 13 2
42 0 9 9 13 1 11 2 11 7 11 2 9 1 0 9 2 2 1 0 9 1 11 2 1 9 0 9 1 11 7 1 0 0 0 9 2 15 4 13 1 11 2
13 0 13 9 1 9 9 1 9 0 0 9 9 2
12 1 11 7 11 9 13 7 0 9 7 11 2
14 9 0 9 13 9 9 11 1 0 9 9 12 12 2
19 1 10 9 13 1 10 9 2 3 3 2 7 9 13 0 9 12 9 2
3 2 11 2
5 11 15 13 1 9
3 0 9 2
15 11 0 9 13 1 0 9 9 1 0 9 12 9 9 2
11 3 1 0 9 13 9 9 12 9 9 2
8 13 15 0 9 9 11 11 2
12 1 12 2 9 0 9 13 11 3 12 9 2
14 1 0 9 13 1 0 9 9 12 9 13 12 9 2
12 0 12 9 9 4 13 9 0 9 0 9 2
8 1 0 9 15 13 0 9 2
7 0 9 4 13 0 9 2
23 12 9 9 9 13 13 1 9 9 2 12 9 1 0 9 7 12 9 13 0 9 9 2
12 9 1 12 9 13 13 1 0 2 0 9 2
27 11 2 15 13 9 0 7 0 9 2 3 3 9 7 0 9 2 13 1 0 9 0 9 12 9 9 2
9 1 9 13 14 12 9 9 9 2
29 9 1 11 7 9 0 0 9 13 3 0 16 1 9 12 2 3 1 10 9 13 11 3 9 1 12 9 9 2
11 9 1 0 9 13 11 11 1 3 0 2
20 1 1 9 1 9 7 10 0 9 13 0 0 9 9 1 9 14 12 9 2
5 1 9 3 3 9
2 11 2
20 0 9 1 9 13 0 0 9 9 1 12 9 9 1 0 9 12 9 9 2
17 1 9 12 2 12 13 0 9 9 12 9 9 2 13 9 11 2
30 0 9 4 13 3 1 9 1 0 9 0 0 9 2 15 4 13 13 3 12 9 9 9 1 0 9 12 9 9 2
25 0 9 9 11 4 13 3 13 0 9 9 1 0 9 2 3 1 0 0 9 7 0 9 11 2
15 9 9 0 9 1 0 9 4 7 13 13 1 9 9 2
29 0 9 9 0 0 9 4 13 3 13 9 9 9 16 9 1 9 2 7 9 15 4 13 13 1 0 9 9 2
12 9 9 1 0 9 3 13 14 12 0 9 2
20 0 9 9 4 1 9 13 13 1 12 9 9 1 9 1 12 9 9 3 2
12 9 15 13 1 12 9 9 1 12 9 3 2
17 0 0 9 9 15 13 1 12 9 9 1 0 9 12 9 9 2
12 1 9 12 15 0 9 13 1 12 9 9 2
20 9 0 9 13 1 0 9 9 9 1 11 2 11 2 11 2 11 7 11 2
20 0 9 9 1 0 11 2 1 11 7 1 11 13 9 1 0 9 9 13 2
6 0 9 9 1 0 9
27 0 12 9 13 1 0 9 13 3 0 9 2 7 16 0 9 13 9 9 1 11 7 1 0 0 9 2
8 13 15 1 9 0 0 9 2
21 0 9 0 9 13 1 0 9 1 0 9 1 0 9 7 9 13 13 7 3 2
35 0 9 9 15 3 13 1 12 5 1 12 9 2 9 2 16 1 9 0 9 13 9 9 12 5 7 1 9 0 7 0 11 12 5 2
33 1 9 11 4 1 10 9 13 1 0 9 3 12 12 0 9 7 1 0 0 9 1 11 1 0 12 9 14 12 12 0 9 2
7 9 15 13 16 0 9 2
16 16 9 0 9 3 13 2 13 14 14 13 0 9 1 9 2
31 1 15 13 9 2 16 9 1 9 3 13 2 3 1 0 9 2 15 15 3 1 0 9 1 9 13 3 16 12 5 2
34 15 11 13 13 1 9 9 10 9 1 12 9 2 9 7 11 7 11 13 13 1 9 9 9 9 10 9 13 1 12 9 2 9 2
3 2 11 2
4 0 9 1 9
15 1 9 7 0 9 0 9 1 11 4 13 0 0 9 2
16 9 13 10 9 13 1 0 9 3 12 2 9 1 0 9 2
13 1 12 9 4 9 0 9 13 13 1 9 9 2
15 13 15 15 1 9 0 9 2 15 9 13 1 10 9 2
24 9 0 9 10 9 1 9 12 12 9 0 13 3 2 9 1 15 9 1 10 9 7 9 2
30 9 4 3 13 13 9 9 1 9 9 7 13 9 0 9 0 9 1 9 9 1 1 15 2 16 13 1 0 9 2
10 0 9 3 13 1 9 9 0 9 2
21 9 9 13 13 1 12 9 1 9 0 9 1 12 9 2 7 15 3 1 15 2
21 1 9 0 12 9 13 9 9 1 9 12 9 9 2 1 0 3 9 1 9 2
37 0 13 13 3 9 9 1 0 9 1 9 11 7 11 2 3 13 0 0 9 1 9 0 9 11 7 3 4 1 9 13 13 0 9 0 9 2
5 2 11 2 11 2
3 9 0 9
8 0 9 13 1 0 9 13 9
3 0 11 2
14 3 3 13 9 13 0 9 0 9 0 9 0 9 2
11 1 10 9 13 9 10 9 1 12 9 2
21 13 1 15 13 7 9 9 9 0 9 3 1 9 2 15 7 4 13 0 9 2
17 1 0 9 0 9 9 13 9 9 9 1 0 9 3 1 12 2
21 1 9 0 9 11 11 3 1 0 9 1 0 0 7 0 9 3 13 0 9 2
15 0 9 0 9 13 13 9 2 15 13 3 0 7 0 2
40 1 9 9 0 9 13 12 2 9 0 9 3 2 3 13 9 9 9 9 11 7 11 2 1 15 13 1 9 1 9 0 9 3 1 0 9 9 11 11 2
26 13 1 0 9 0 9 2 15 4 1 9 12 7 12 3 13 1 10 9 9 9 7 9 11 11 2
11 9 0 9 13 1 10 9 1 0 9 2
50 0 9 0 9 3 13 12 0 9 1 0 11 2 3 15 3 2 13 3 0 9 11 11 2 3 1 11 2 11 2 11 2 11 7 11 2 12 0 9 7 0 9 0 9 1 11 1 0 11 2
33 1 0 12 9 0 9 1 12 9 9 9 15 9 0 9 3 13 0 9 2 7 7 4 13 9 2 15 15 13 1 0 9 2
5 10 9 1 0 9
5 11 2 11 2 2
13 10 9 15 13 1 0 0 9 1 0 9 11 2
42 1 0 9 7 0 9 13 9 0 0 9 1 9 9 2 0 9 12 9 2 7 9 9 2 0 9 12 9 2 2 1 0 9 4 13 3 9 9 7 9 9 2
10 0 0 9 15 4 13 12 2 9 2
7 11 9 13 0 0 0 9
2 11 2
18 0 9 7 9 11 9 13 9 1 9 10 9 1 0 9 0 9 2
10 13 15 3 0 0 9 1 0 9 2
15 1 0 9 13 9 3 0 7 9 13 4 13 1 9 2
31 11 9 4 13 14 12 9 1 0 9 2 7 15 7 1 0 9 2 7 7 1 9 10 0 7 0 9 1 10 9 2
18 1 1 0 0 9 13 1 11 0 13 3 0 9 1 11 1 11 2
8 1 9 1 9 13 0 9 2
32 9 9 13 9 9 9 0 0 13 0 0 9 1 0 9 0 11 1 9 2 11 7 11 1 11 2 7 15 1 0 9 2
18 10 9 3 13 9 1 9 10 9 1 9 0 11 1 9 2 11 2
9 0 9 4 13 4 13 1 9 2
5 13 9 15 14 13
9 9 9 7 13 13 3 16 0 11
3 0 11 2
21 16 3 0 15 7 1 0 0 9 1 9 0 9 9 9 11 11 13 9 9 2
43 16 0 0 9 13 1 10 9 9 1 12 0 9 2 0 0 9 1 12 7 12 9 7 0 0 9 13 13 3 1 9 12 0 9 11 2 13 15 9 0 0 9 2
30 9 0 9 2 15 13 14 3 10 9 2 15 3 1 11 1 0 9 13 1 9 1 9 12 7 12 9 1 9 2
32 3 0 0 9 13 3 3 0 0 9 7 0 9 2 10 0 0 9 13 11 2 3 1 9 1 9 2 13 11 2 11 2
19 9 9 13 1 0 11 13 3 1 11 2 7 13 3 1 11 7 11 2
14 1 0 9 15 9 10 9 3 13 3 0 9 11 2
24 1 12 0 9 9 13 13 12 7 12 9 3 7 1 10 9 13 13 12 7 12 0 9 2
20 15 1 11 1 12 9 13 1 9 9 2 15 1 15 13 12 7 12 9 2
12 0 9 9 1 12 9 13 3 1 12 9 2
16 9 15 13 3 12 9 2 16 10 0 9 13 3 12 9 2
20 1 0 9 13 10 9 9 1 12 9 11 7 7 3 13 0 1 0 9 2
14 1 9 11 13 1 0 0 9 3 12 9 9 9 2
9 0 0 9 13 12 9 1 9 2
3 9 2 11
4 9 11 13 13
13 9 9 13 9 7 9 13 9 9 11 16 0 9
2 11 11
20 9 7 9 9 1 9 11 1 11 13 1 9 12 1 3 16 12 9 9 2
15 1 0 9 9 12 9 1 0 9 15 13 1 0 9 2
31 16 13 11 11 2 12 1 12 9 0 9 11 2 0 9 13 1 0 9 1 9 9 1 9 7 13 9 9 1 9 2
22 0 9 13 1 9 0 9 9 9 12 9 9 2 11 11 2 11 11 7 11 11 2
16 1 9 12 9 15 15 13 13 15 0 0 9 1 9 9 2
13 1 9 11 2 11 13 9 9 0 9 0 9 2
12 1 15 13 7 9 0 9 7 0 9 9 2
14 9 13 1 9 0 1 0 9 7 1 3 0 9 2
15 13 15 3 1 0 9 2 9 1 11 2 9 1 11 2
11 0 9 13 1 11 1 0 9 0 9 2
17 1 9 15 13 1 9 9 11 16 9 2 15 13 1 9 0 2
18 1 9 11 2 11 13 3 1 10 9 10 9 2 16 3 13 13 2
12 9 13 13 9 0 0 9 3 1 12 9 2
18 16 13 1 11 11 2 11 2 9 4 3 13 13 0 0 0 9 2
14 3 15 7 13 3 0 0 9 1 9 7 0 9 2
7 10 9 13 3 1 9 2
16 9 11 13 2 16 15 3 13 9 1 9 0 7 0 9 2
7 15 13 1 15 3 0 2
11 9 13 1 0 9 2 7 0 7 9 2
19 1 0 9 13 9 11 0 9 12 9 9 2 3 13 14 12 9 9 2
28 9 9 1 0 9 13 11 2 11 16 0 1 0 9 2 7 1 15 0 9 1 9 2 0 9 7 9 2
9 9 3 13 9 2 7 13 13 2
18 14 13 9 7 13 1 9 13 9 3 1 9 2 13 11 2 11 2
6 9 11 13 12 9 2
15 1 10 0 9 13 0 9 2 9 2 9 7 0 9 2
25 1 12 9 13 9 1 9 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 7 11 2
11 3 1 12 9 1 9 9 13 1 11 2
20 1 0 9 1 9 10 9 1 0 12 9 13 1 9 11 1 0 9 9 2
14 1 9 0 0 9 13 3 1 0 9 3 3 15 2
23 9 11 4 3 3 13 7 13 1 0 9 9 7 9 11 12 0 9 0 7 0 9 2
4 9 1 0 9
12 0 9 1 11 13 12 9 9 1 12 0 9
2 11 2
27 14 12 0 9 2 7 2 12 9 2 1 9 11 13 0 9 1 11 9 1 0 9 1 9 12 9 2
32 9 2 15 13 0 9 9 2 13 0 9 14 1 9 9 1 9 7 9 9 3 0 9 0 1 9 9 0 9 0 9 2
17 0 11 2 3 9 1 9 9 9 2 4 13 1 0 0 9 2
26 13 0 9 9 9 2 1 15 4 13 9 2 15 4 1 0 9 3 13 1 9 1 0 0 9 2
12 0 9 13 9 2 1 15 13 14 12 9 2
18 1 11 11 2 9 0 9 2 13 0 9 2 15 1 10 9 13 2
32 9 1 0 9 13 14 12 9 9 0 7 13 3 9 12 9 2 16 15 1 10 9 13 1 0 9 1 9 11 1 11 2
12 1 9 9 13 1 11 3 9 0 16 11 2
8 3 0 9 13 3 0 9 2
23 3 0 0 9 13 9 9 2 7 15 13 9 2 3 15 3 0 9 1 9 9 13 2
19 1 11 11 2 11 2 13 12 9 2 9 1 9 7 9 10 12 9 2
13 3 16 12 9 9 4 13 1 9 1 9 12 2
10 0 9 12 9 13 3 12 9 9 2
23 7 1 10 9 13 0 9 3 3 16 12 9 9 2 15 4 13 9 0 9 1 9 2
21 3 11 13 1 0 9 9 1 9 12 9 2 1 12 9 3 16 1 9 12 2
11 3 15 13 2 16 9 13 3 3 9 2
22 1 0 9 13 9 11 14 12 0 0 9 9 1 9 7 3 3 16 12 1 9 2
5 11 13 9 1 11
3 0 11 2
39 0 9 11 11 11 2 11 3 13 9 1 9 9 0 9 1 11 0 9 7 1 9 1 9 1 9 11 1 0 11 13 2 16 0 9 13 13 9 2
20 11 13 2 16 0 9 13 0 2 16 9 1 11 13 13 1 10 0 9 2
40 3 1 9 13 3 1 9 1 11 12 0 0 9 2 0 9 9 9 11 11 7 0 9 9 9 11 11 2 15 13 0 9 9 1 9 1 12 0 9 2
16 3 3 13 9 9 2 15 4 15 0 9 13 13 2 12 2
6 9 1 9 9 0 9
95 11 13 9 0 9 7 13 15 1 10 9 2 2 15 13 9 1 9 9 1 10 9 2 2 1 10 9 13 0 9 2 2 1 10 9 13 0 9 2 2 1 15 15 13 13 9 2 1 9 2 7 0 9 2 2 15 13 0 9 2 9 1 9 12 2 2 2 9 9 9 7 0 9 2 2 9 9 2 15 15 13 2 7 15 15 13 2 3 2 0 9 1 10 9 2
14 11 2 0 9 2 9 9 2 11 2 9 2 11 11
19 1 11 13 1 9 1 9 9 9 2 9 13 2 13 15 0 9 9 2
6 9 0 9 13 0 2
20 0 9 13 1 0 9 2 0 0 9 7 1 9 1 0 9 1 0 9 2
19 0 13 9 1 0 9 2 1 0 9 1 0 9 7 1 0 0 9 2
46 0 9 1 11 15 13 13 1 9 1 12 1 12 9 2 9 2 0 9 1 9 7 9 1 12 9 2 7 12 9 2 9 2 0 9 1 9 1 12 7 12 9 5 9 12 2
27 1 9 0 9 15 13 1 12 9 2 9 12 1 9 2 1 9 9 1 12 9 2 9 12 1 9 2
17 10 9 15 13 9 12 7 12 9 1 9 7 13 15 9 9 2
9 1 9 13 12 7 12 0 9 2
22 0 9 10 9 13 9 7 9 0 9 1 9 11 2 9 9 0 9 1 0 9 2
14 1 9 15 10 9 13 12 7 12 9 3 1 9 2
8 11 11 2 0 9 2 11 11
20 1 1 9 9 7 1 9 9 2 0 9 2 13 9 1 9 9 3 0 2
25 10 9 13 9 1 9 1 0 9 2 7 7 13 9 14 1 0 9 2 7 7 1 0 9 2
16 0 13 7 9 7 9 2 7 1 0 9 7 1 0 9 2
18 13 9 1 0 9 2 0 9 7 1 0 9 0 3 1 0 9 2
14 9 9 2 9 7 9 13 3 0 1 9 7 9 2
37 3 2 9 9 12 5 12 1 12 1 12 9 2 9 2 9 1 12 9 2 1 12 9 2 9 2 0 9 1 12 1 12 9 5 9 12 2
13 9 9 13 1 12 1 12 9 2 9 12 3 2
11 9 1 0 9 15 13 1 9 3 3 2
15 9 9 13 0 2 13 1 9 7 9 2 15 13 9 2
6 3 7 13 12 5 2
15 3 16 9 13 7 1 0 9 13 2 13 9 10 9 2
16 10 9 4 13 1 9 2 12 7 13 0 9 1 0 9 2
14 13 9 9 0 9 11 7 3 0 9 0 9 11 2
27 13 1 9 0 9 1 10 9 2 13 1 9 1 9 1 11 2 11 2 11 2 11 2 11 7 0 2
19 0 11 2 9 2 11 2 0 7 0 9 2 0 9 2 9 2 11 11
11 9 1 9 1 9 9 10 9 13 0 2
14 1 10 9 3 13 9 9 7 9 9 13 9 9 2
42 3 1 10 9 13 12 0 0 9 2 1 15 2 7 13 15 2 16 1 0 9 7 12 1 15 2 16 4 13 7 0 9 2 13 0 15 0 9 0 9 13 2
37 3 13 3 0 9 9 2 3 1 9 9 1 0 9 0 0 9 7 10 9 2 13 1 0 9 9 9 7 3 15 13 7 13 15 1 0 2
39 0 9 13 1 9 7 9 9 7 0 9 0 3 3 9 9 2 0 9 2 0 11 2 11 1 11 2 0 9 1 11 2 11 2 11 1 11 2 2
16 3 0 13 9 1 0 0 9 7 9 1 9 1 0 9 2
38 0 9 9 12 5 12 15 13 1 12 9 2 9 2 12 5 12 1 12 9 2 9 7 0 9 0 0 9 1 12 9 2 1 12 9 2 9 2
12 9 0 9 13 9 1 9 7 9 0 9 2
11 13 15 1 12 1 12 9 2 9 12 2
26 9 9 9 7 0 9 3 13 1 9 1 9 2 13 1 9 1 12 1 12 9 2 9 12 3 2
21 10 9 15 13 1 12 1 12 9 1 9 0 9 7 1 12 5 4 13 0 2
9 10 9 13 13 1 9 9 12 2
20 1 0 0 9 13 0 9 1 9 9 1 0 9 7 13 0 9 1 9 2
5 9 0 9 3 13
5 11 2 11 2 2
42 0 9 13 13 13 0 9 1 9 0 9 1 12 0 9 3 2 3 4 3 13 2 3 3 2 13 3 9 9 11 2 11 1 9 1 10 0 9 11 2 11 2
7 1 11 13 15 0 9 2
41 13 4 15 2 16 13 9 0 9 1 11 7 0 0 9 2 16 4 13 13 1 9 12 9 3 1 11 2 7 3 1 9 13 0 9 1 11 2 13 11 2
13 11 4 13 1 9 9 13 1 9 9 12 9 2
20 3 4 15 13 3 1 15 2 16 4 15 13 0 9 2 15 0 9 13 2
27 13 4 15 1 11 13 11 2 11 2 15 4 1 10 9 13 2 16 1 15 13 15 0 2 13 11 2
7 1 0 9 1 12 9 9
2 11 2
19 1 0 9 0 9 0 9 1 0 9 13 9 9 0 9 3 12 9 2
13 13 1 0 9 2 16 3 13 9 1 0 9 2
12 1 9 13 1 12 2 9 13 3 12 9 2
33 9 13 13 9 12 9 2 10 9 13 3 12 5 9 0 1 9 0 9 2 16 9 1 0 12 9 13 3 12 5 0 9 2
9 9 11 13 13 0 9 7 13 9
2 11 2
7 4 4 13 1 9 9 2
9 3 15 13 14 3 2 7 3 2
3 13 15 2
6 10 9 13 3 0 2
5 13 3 9 9 2
29 10 9 7 9 13 3 0 9 1 11 1 9 9 2 13 9 11 1 9 2 15 4 3 13 1 0 9 11 2
5 9 9 13 9 2
14 11 13 3 1 9 9 1 0 9 1 0 9 11 2
8 1 9 1 15 13 15 13 2
27 9 9 11 11 13 2 16 15 1 11 13 2 7 13 13 9 2 15 15 9 13 2 3 1 0 9 2
22 9 13 1 9 9 1 15 2 16 15 0 9 13 1 9 1 9 11 1 9 12 2
12 13 2 16 4 1 9 9 3 13 1 11 2
6 13 9 2 13 15 2
8 13 12 1 9 0 9 9 2
7 1 10 9 15 9 13 2
16 7 14 15 13 1 15 2 16 4 13 0 9 7 13 9 2
20 1 10 9 13 2 15 13 0 9 2 16 15 7 3 0 9 13 9 9 2
4 0 9 13 9
14 12 1 0 9 1 11 2 9 9 2 12 2 13 9
5 11 2 11 2 2
21 9 9 9 11 11 13 1 0 0 9 1 11 9 0 11 3 9 0 15 9 2
11 13 15 13 1 0 9 7 9 1 11 2
48 1 0 9 4 9 9 11 11 1 9 0 9 11 13 2 16 3 10 9 2 1 11 15 13 0 11 2 13 1 9 9 1 0 0 0 9 9 2 12 2 15 13 1 11 11 2 0 2
18 15 3 2 16 15 3 13 1 9 12 0 9 9 2 12 1 11 2
11 11 7 9 13 7 11 15 1 11 13 2
24 1 0 9 9 11 7 9 9 7 9 13 2 16 13 1 9 2 3 15 11 13 1 9 2
9 11 15 13 7 9 7 0 9 2
24 14 3 2 9 1 11 13 1 12 9 9 7 1 11 15 1 9 9 13 1 3 12 9 2
15 9 7 13 0 9 7 9 13 9 11 2 16 13 11 2
33 0 1 0 9 11 7 9 9 9 13 2 16 13 4 3 1 12 9 1 0 9 9 13 9 1 9 9 1 9 9 2 12 2
20 9 11 11 11 9 1 10 9 3 13 2 13 15 1 0 9 2 0 11 2
52 1 9 0 9 11 7 13 2 16 9 11 2 1 15 2 16 13 1 0 9 0 1 11 7 13 1 0 9 0 2 13 1 9 9 0 0 11 7 11 2 15 15 1 9 1 9 9 2 12 3 13 2
31 9 13 2 16 16 4 4 3 13 0 9 0 9 11 7 9 2 15 13 1 9 12 9 2 13 4 1 9 9 11 2
28 11 13 1 15 0 13 11 7 1 9 9 12 1 0 9 1 11 2 1 15 4 9 2 12 1 9 13 2
6 3 13 9 2 3 2
21 9 9 3 13 2 16 13 9 1 9 13 9 11 2 11 1 0 9 1 11 2
18 3 7 13 13 9 2 16 9 13 3 1 9 9 0 1 0 9 2
1 9
2 11 11
31 3 0 9 1 9 0 9 11 2 0 9 2 0 9 7 9 13 0 9 1 9 0 9 2 0 0 9 13 0 11 2
20 0 9 1 15 13 1 12 9 2 1 9 12 12 9 1 9 12 2 12 2
19 9 1 9 2 9 2 9 2 9 2 0 9 0 9 14 1 0 13 2
16 1 9 9 0 9 1 0 11 13 3 0 0 9 0 9 2
39 0 9 1 10 9 4 13 1 9 9 12 2 3 11 11 3 13 13 0 9 2 3 0 9 7 1 9 0 9 13 1 9 11 0 9 12 7 12 2
19 11 13 0 11 1 0 9 2 15 3 13 1 9 9 0 0 0 9 2
33 9 11 1 9 0 9 2 11 3 13 10 0 9 3 2 16 15 15 13 13 10 0 0 9 2 13 1 9 1 9 11 9 2
15 9 0 2 0 9 1 0 9 13 9 0 7 0 11 2
16 16 13 2 13 1 11 1 9 1 0 9 9 1 0 9 2
33 13 15 13 9 1 11 1 9 12 2 13 13 0 9 0 9 1 9 12 2 3 1 9 13 4 13 0 9 1 12 9 3 2
17 11 15 13 0 2 3 0 9 1 9 9 0 11 1 9 13 2
15 1 0 9 1 9 12 15 15 13 13 1 9 0 9 2
15 13 3 9 1 9 11 1 12 9 9 7 9 0 11 2
22 9 11 9 13 2 1 0 11 4 4 3 9 0 11 13 1 9 7 9 0 9 2
16 7 11 1 0 9 10 0 9 13 1 9 0 11 0 9 2
18 10 9 1 11 15 4 1 9 9 13 2 13 13 1 15 7 3 2
17 1 9 12 13 15 3 2 0 9 0 0 9 1 11 15 13 2
6 13 3 11 7 11 2
9 10 9 2 16 0 2 7 0 2
10 13 15 9 2 0 9 15 13 15 2
6 7 10 9 13 0 2
4 0 9 0 9
5 11 2 11 2 2
24 11 13 1 9 9 1 0 9 0 9 11 11 2 15 9 13 2 13 9 0 9 1 11 2
29 11 11 9 12 1 9 12 9 9 13 13 1 0 2 3 0 9 2 3 1 9 0 9 1 9 7 0 9 2
11 1 0 9 13 10 9 3 9 1 11 2
20 16 13 11 9 0 9 1 11 9 2 11 11 2 13 0 12 9 3 13 2
23 14 3 2 16 13 13 0 9 2 7 9 13 7 3 0 9 9 1 9 2 13 9 2
6 9 1 0 9 1 11
5 11 2 11 2 2
27 0 0 0 9 0 9 2 0 2 9 2 2 11 13 1 9 1 9 0 0 9 1 9 9 9 11 2
20 1 9 7 12 9 4 13 1 9 9 12 2 9 13 7 9 9 11 11 2
10 9 1 9 9 13 9 12 9 9 2
10 0 9 13 3 16 12 9 0 9 2
13 9 9 13 13 15 9 2 15 15 13 1 0 9
5 11 2 11 2 2
22 9 9 12 12 12 13 1 12 2 9 1 9 15 9 2 15 15 13 1 0 9 2
12 13 15 9 10 9 2 10 9 13 11 11 2
10 9 13 1 0 9 0 9 7 9 2
11 1 10 9 4 13 9 1 0 0 11 2
32 13 15 0 0 9 7 9 11 11 2 15 15 3 1 11 13 9 9 3 1 9 0 9 1 9 9 2 11 2 11 11 2
23 9 11 2 15 15 13 9 10 9 2 13 2 16 1 11 3 0 11 13 12 9 9 2
12 13 1 9 12 9 2 15 13 1 9 9 2
11 15 15 13 1 9 7 15 13 2 3 2
22 9 0 0 9 2 1 15 13 2 15 13 9 2 16 4 15 15 1 10 9 13 2
11 9 2 15 9 13 2 13 3 1 9 2
40 0 9 9 9 13 3 0 9 11 11 11 11 7 9 11 2 11 2 9 9 7 0 9 13 9 0 9 2 2 11 2 11 2 11 2 11 7 11 11 2
24 9 9 13 9 9 7 13 2 16 1 9 2 15 13 9 7 9 9 2 13 0 9 0 2
10 13 15 15 13 15 9 9 0 9 2
4 3 1 9 12
8 7 0 9 13 13 10 0 9
27 1 9 0 9 7 1 9 9 9 4 10 9 13 13 0 9 1 9 7 9 0 0 9 16 0 9 2
28 0 9 2 15 10 9 13 2 13 0 9 1 9 9 1 9 9 2 15 13 9 0 7 0 0 9 2 2
24 9 13 1 9 7 9 0 1 0 7 0 9 2 9 1 9 9 2 0 9 7 0 2 2
24 1 9 9 7 9 13 1 0 9 2 3 1 0 2 0 2 0 2 0 7 0 9 2 2
18 1 9 1 0 0 9 13 9 2 0 9 2 0 9 7 9 2 2
17 13 1 9 9 0 9 2 9 2 0 9 2 1 9 9 2 2
7 13 9 1 0 9 2 2
35 13 0 9 1 9 1 9 9 1 9 7 0 1 9 2 9 2 9 1 9 2 0 9 2 9 1 9 2 9 1 9 9 2 2 2
19 13 1 9 0 9 1 0 9 1 9 2 13 0 9 2 0 9 2 2
13 3 3 3 13 9 9 7 9 1 9 1 9 2
9 2 13 9 9 1 9 0 9 2
17 0 9 13 3 1 12 2 12 2 9 0 1 9 0 0 9 2
15 16 0 9 13 0 9 2 13 15 13 1 12 2 12 2
24 9 15 13 13 16 9 9 1 0 9 2 16 10 9 13 1 12 0 9 9 12 12 9 2
27 1 9 1 9 1 9 15 13 9 9 9 1 9 7 9 2 16 13 1 9 7 1 9 9 7 9 2
18 13 2 14 9 0 9 0 1 9 2 13 15 7 9 0 9 2 2
35 1 9 13 1 0 9 3 1 9 12 9 9 1 9 0 9 2 9 1 0 9 7 9 1 0 9 9 7 9 1 0 0 9 2 2
9 13 9 0 9 0 0 9 2 2
4 13 0 9 2
16 2 16 1 0 9 13 0 9 1 9 2 13 9 13 9 2
7 2 13 9 9 7 9 2
22 2 13 9 9 2 13 0 9 0 9 2 13 0 9 9 2 9 9 7 0 9 2
3 2 11 2
2 0 9
5 11 2 11 2 2
20 9 1 9 11 11 2 15 13 13 9 3 0 9 2 13 0 9 1 11 2
16 9 0 9 3 13 1 9 7 3 13 1 10 9 7 9 2
39 0 9 13 1 11 3 12 9 7 1 10 9 3 15 15 13 13 9 0 9 9 0 9 2 13 3 0 9 2 13 1 9 11 1 9 1 9 9 2
18 1 0 9 15 13 1 9 9 2 3 13 4 1 0 9 13 9 2
20 16 13 11 9 0 0 9 11 11 2 0 9 1 9 0 9 13 0 9 2
19 1 11 13 14 14 12 9 1 9 9 2 7 13 12 9 15 0 9 2
5 12 9 13 12 9
5 11 2 11 2 2
16 0 9 9 0 9 9 11 11 15 13 3 1 9 1 11 2
10 9 15 13 12 9 2 3 0 9 2
48 9 1 9 2 0 2 11 11 2 15 15 1 9 9 13 3 9 9 7 9 2 13 1 0 9 3 16 12 9 1 11 7 9 2 13 12 9 1 9 7 1 9 13 10 9 3 13 2
13 9 1 9 0 9 15 13 1 12 2 12 9 2
11 0 9 13 1 12 7 12 9 1 9 2
32 9 13 1 9 9 7 9 3 0 16 9 2 13 0 2 13 1 9 0 7 0 9 3 13 2 13 11 9 9 11 11 2
6 9 1 0 0 9 13
5 11 2 11 2 2
24 14 1 9 13 1 9 9 2 15 3 3 13 9 0 9 1 9 0 1 9 0 0 9 2
23 16 15 13 9 1 0 9 2 13 1 9 3 13 10 9 7 13 9 9 9 0 9 2
23 16 9 0 9 4 3 13 2 1 9 11 9 13 9 2 3 4 10 0 9 13 13 2
14 1 15 13 0 9 1 9 9 9 0 0 9 11 2
18 3 15 13 9 3 13 3 9 0 9 2 7 9 1 10 9 13 2
32 9 9 11 2 15 15 3 13 9 2 7 13 14 1 0 9 2 13 1 15 0 9 2 1 15 13 10 9 1 9 9 2
20 9 13 9 12 9 9 7 13 1 0 2 15 15 1 11 1 0 9 13 2
6 9 1 0 9 0 9
5 9 11 11 2 11
5 9 0 9 1 11
2 11 2
21 1 12 9 0 9 1 0 9 13 1 9 3 1 9 11 1 9 11 1 11 2
12 1 0 9 9 13 9 0 9 7 9 13 2
15 3 1 15 13 9 0 9 9 0 9 1 11 11 11 2
27 0 9 9 0 9 2 9 2 0 2 11 13 9 9 2 1 0 9 13 1 0 9 7 13 1 9 2
11 9 15 3 13 1 9 7 13 1 9 2
16 9 1 0 9 13 9 2 15 15 13 9 1 9 12 9 2
25 7 16 0 9 9 2 15 1 9 9 13 1 12 9 2 4 0 9 13 2 9 15 13 13 2
22 0 9 1 9 4 13 1 9 1 11 11 1 9 7 3 15 13 1 9 0 9 2
13 0 9 7 13 1 9 3 12 9 2 13 11 2
1 3
15 1 0 9 9 1 11 12 3 13 9 0 9 11 11 2
10 1 9 9 4 13 1 9 0 9 2
19 0 9 0 9 1 0 9 13 1 9 0 9 1 11 1 0 9 12 2
21 9 0 9 1 9 2 9 13 9 2 15 13 1 9 1 9 1 0 9 9 2
17 13 15 15 3 12 9 1 0 9 2 15 15 4 13 3 9 2
26 9 0 9 0 1 12 2 9 1 0 9 0 9 1 9 9 13 10 9 11 11 9 1 0 9 2
13 1 9 0 9 13 9 0 9 3 12 9 9 2
13 9 4 13 1 9 9 0 9 11 1 0 9 2
10 15 4 13 1 9 13 15 9 11 2
31 0 9 13 7 3 1 9 1 11 1 11 2 7 16 11 11 2 15 4 9 13 1 9 2 13 3 1 10 0 9 2
14 3 15 9 13 1 15 2 16 4 9 13 1 9 2
11 13 7 1 9 9 1 9 12 9 9 2
4 0 9 1 11
5 11 2 11 2 2
16 3 9 9 11 11 9 13 4 1 11 13 0 0 0 9 2
24 1 10 9 15 13 3 3 3 7 1 9 2 3 4 9 13 0 2 13 0 9 7 9 2
23 1 9 2 10 9 13 12 9 9 2 13 3 0 9 2 9 1 12 9 7 0 9 2
16 9 9 13 3 3 3 2 1 9 15 7 13 14 1 9 2
18 1 10 9 15 4 12 9 0 2 0 7 0 9 13 1 0 9 2
16 9 4 13 3 9 0 11 0 1 11 7 9 1 0 11 2
30 1 9 11 2 3 13 9 3 10 2 13 9 11 11 11 2 9 13 1 12 9 7 3 13 1 9 3 0 9 2
15 13 4 2 16 3 9 10 9 4 10 9 13 0 9 2
13 3 15 13 2 16 15 13 3 14 9 0 9 2
18 12 9 4 3 1 10 9 13 9 2 9 1 15 3 15 7 13 2
11 1 0 9 9 15 3 13 13 0 9 2
6 7 7 9 13 10 2
14 0 9 4 13 16 9 1 0 9 1 9 1 10 9
5 11 2 11 2 2
22 0 9 4 13 16 9 1 0 9 2 15 4 1 9 0 9 13 13 1 9 0 2
28 3 13 7 3 0 2 7 7 13 2 14 10 0 9 3 0 9 1 9 1 0 9 2 4 1 15 13 2
11 9 0 13 3 0 16 1 9 3 0 2
16 13 15 1 10 9 2 13 15 1 9 9 7 3 7 13 2
13 3 13 9 9 1 15 2 15 0 9 3 13 2
34 1 12 9 10 9 2 3 13 1 12 9 2 13 1 11 3 12 2 16 9 13 3 0 2 13 9 0 9 1 0 9 11 11 2
15 13 1 9 14 3 3 0 9 13 1 0 9 3 0 2
8 9 3 13 9 1 9 9 2
13 7 7 1 12 9 13 1 10 9 15 13 9 2
13 1 9 0 7 0 9 15 13 10 9 1 9 2
20 13 3 3 14 3 2 13 2 14 15 13 1 9 9 2 13 11 2 11 2
25 3 1 0 9 7 9 2 15 13 1 10 9 12 7 12 9 1 9 2 13 0 0 9 9 2
7 13 3 1 12 9 3 2
35 13 2 14 9 9 7 13 0 9 10 9 2 13 15 3 1 0 9 0 9 2 3 3 9 2 15 13 13 1 9 9 1 0 9 2
7 0 9 13 7 3 0 2
9 3 9 13 1 9 3 12 9 2
7 9 13 13 0 0 9 2
8 3 10 9 13 0 0 9 2
29 1 10 9 13 2 16 9 13 1 0 9 7 9 0 9 13 0 9 3 16 1 12 9 2 13 11 2 11 2
12 0 9 2 3 13 0 9 2 1 11 13 2
5 9 13 0 9 2
15 9 1 0 9 13 1 9 9 2 15 13 0 9 0 2
17 3 13 3 1 0 0 9 1 0 9 0 2 0 7 0 9 2
13 16 15 0 9 13 2 4 13 7 1 0 9 2
7 4 15 0 9 13 11 2
2 11 2
23 9 9 1 9 9 1 0 9 1 11 11 3 13 0 0 9 11 11 9 9 11 11 2
22 9 2 16 15 9 13 2 13 9 0 9 1 11 2 15 9 13 0 9 1 9 2
5 11 15 13 3 2
30 9 1 15 13 0 2 16 0 0 9 13 9 1 0 9 2 0 9 1 9 2 1 9 2 15 13 0 1 9 2
30 9 13 9 7 1 15 2 16 9 3 13 0 9 2 16 13 2 16 11 1 9 0 9 13 0 9 2 13 11 2
14 16 9 9 13 2 4 1 15 13 0 9 1 11 2
28 15 7 9 0 9 13 2 7 9 7 10 9 13 7 0 9 13 13 2 16 4 1 9 3 13 7 13 2
10 0 9 3 13 9 13 9 0 9 2
6 0 9 13 9 0 9
7 11 2 11 2 11 2 2
20 3 1 0 2 0 9 3 13 0 9 1 9 0 9 0 10 9 11 11 2
34 16 11 13 9 0 9 9 11 11 2 11 2 2 1 0 9 4 4 13 1 9 1 0 0 9 0 15 9 0 11 1 9 12 2
19 9 1 15 13 1 3 0 7 3 0 9 7 13 15 9 0 9 9 2
28 1 9 2 16 0 9 13 9 9 0 9 2 11 13 2 16 4 4 3 13 2 16 4 15 1 15 13 2
8 10 9 7 14 9 9 13 2
27 1 10 9 13 0 9 16 0 9 2 3 4 13 10 0 9 7 13 15 13 9 2 15 13 1 0 2
13 11 15 3 3 13 1 10 0 9 11 2 11 2
24 0 7 0 9 1 15 13 0 9 0 15 9 9 9 1 9 1 9 13 1 15 0 9 2
15 13 4 15 1 0 9 9 2 14 1 0 2 13 11 2
21 3 0 0 9 1 0 9 1 9 13 14 3 0 2 16 15 13 13 10 9 2
6 11 2 11 13 0 9
7 11 2 11 2 11 2 2
13 0 9 0 9 11 2 11 15 3 13 11 11 2
16 16 9 0 9 13 1 12 9 1 11 1 0 3 0 9 2
15 1 9 11 3 1 9 13 7 1 9 13 16 0 9 2
5 9 9 9 13 0
9 0 9 13 2 16 13 11 2 11
5 11 2 11 2 2
28 0 9 0 9 11 11 3 13 10 9 1 15 2 16 4 4 13 1 9 1 10 9 1 3 0 9 9 2
29 13 15 3 13 1 9 2 1 15 0 9 9 13 1 10 9 9 7 13 9 0 0 9 1 9 1 9 9 2
28 9 1 0 9 0 9 13 0 9 0 9 9 2 11 2 2 16 13 0 9 1 9 0 10 9 1 0 2
16 9 13 11 2 11 1 9 0 9 7 1 9 1 0 9 2
18 15 15 13 13 15 2 16 9 2 15 15 13 9 13 2 13 9 2
21 9 0 9 11 9 13 2 16 4 1 0 9 13 16 1 9 0 9 7 9 2
12 9 0 9 1 0 9 4 13 13 1 9 2
22 9 4 13 3 2 16 9 9 13 0 9 0 9 9 1 9 11 7 10 0 9 2
17 9 13 9 13 3 1 9 2 16 15 9 9 13 9 0 9 2
7 0 9 0 9 9 13 2
7 9 7 13 9 0 9 2
35 16 4 15 13 2 13 4 1 9 9 0 2 16 0 9 9 1 9 13 2 13 3 1 9 11 11 11 1 9 9 7 9 9 9 2
12 9 11 2 11 1 0 9 1 15 0 13 2
20 0 9 9 1 9 9 1 9 2 16 13 0 9 2 4 13 3 16 9 2
38 9 9 3 13 3 2 16 9 4 13 9 1 9 2 15 13 1 9 0 9 2 13 3 2 16 15 13 1 0 9 9 2 13 15 11 2 11 2
3 13 11 11
2 11 2
31 0 0 9 7 9 10 9 13 9 0 9 9 11 2 11 1 0 0 9 9 11 11 2 15 13 1 0 0 9 11 2
7 13 15 0 9 11 11 2
28 1 10 9 13 14 9 9 9 1 0 11 2 1 15 13 1 15 0 9 13 3 3 7 13 3 9 9 2
28 12 9 13 2 16 9 0 9 15 0 0 0 9 13 7 13 15 1 15 9 0 9 2 13 11 2 11 2
5 0 9 1 9 11
2 11 2
33 1 0 9 1 0 9 7 11 1 9 0 9 0 9 2 11 2 15 3 13 9 0 9 11 11 3 1 0 9 9 11 11 2
9 13 15 11 11 1 9 9 9 2
27 12 9 15 3 13 1 0 9 2 9 0 9 7 1 0 9 1 0 9 1 9 12 9 1 0 9 2
26 9 11 2 15 3 13 1 0 9 0 9 2 15 3 13 1 9 11 11 7 9 0 9 11 11 2
12 13 1 0 0 9 0 9 9 1 0 11 2
4 11 2 13 9
7 11 2 11 2 11 2 2
25 13 9 13 1 9 2 15 13 2 16 13 3 0 2 16 4 9 13 1 9 9 0 0 9 2
21 1 15 2 16 4 9 10 9 13 3 13 2 13 0 9 15 10 9 13 9 2
13 13 15 11 9 0 9 9 11 11 2 11 2 2
15 16 15 10 9 13 1 0 9 2 3 15 15 3 13 2
20 13 4 15 1 10 9 9 7 13 4 15 0 13 0 0 9 2 13 11 2
8 3 7 13 10 9 11 9 2
8 0 9 1 9 0 9 13 2
35 15 0 13 2 16 1 15 13 13 0 9 2 3 9 13 0 9 1 9 9 7 10 9 1 9 9 13 1 0 9 0 9 1 9 2
7 10 9 13 9 13 3 2
15 1 9 0 9 11 13 2 16 7 10 9 1 9 13 2
24 13 9 13 3 7 13 15 3 1 0 9 2 13 9 2 15 9 13 1 9 2 13 9 2
5 15 3 3 13 2
6 13 10 9 3 9 2
5 1 9 9 13 2
13 7 13 15 9 2 15 13 13 0 9 0 9 2
11 13 4 0 2 16 4 9 9 11 13 2
19 13 7 13 15 9 2 16 0 9 13 0 9 2 7 13 15 15 13 2
9 11 13 2 16 13 9 15 13 2
19 7 1 9 0 9 9 11 0 2 11 2 13 0 9 1 0 9 9 2
7 0 9 3 13 9 11 2
18 13 7 2 16 1 0 0 9 7 7 1 11 15 1 9 13 13 2
24 1 0 0 9 13 0 2 16 9 10 9 13 0 2 7 15 13 7 1 0 11 2 13 2
11 0 13 0 9 1 0 9 0 0 9 2
22 13 15 2 16 9 13 4 3 13 9 2 15 15 3 13 16 0 9 1 0 9 2
9 0 11 4 1 11 13 3 1 9
5 11 2 11 2 2
17 9 0 11 7 9 4 13 4 1 11 3 13 1 9 9 12 2
12 1 10 0 0 9 15 13 10 9 11 11 2
26 9 1 9 9 0 0 9 2 3 15 12 0 9 13 1 11 2 3 0 11 1 9 9 11 13 2
6 13 15 3 10 9 2
27 10 9 13 2 13 11 1 9 2 16 0 11 3 13 9 1 9 10 9 2 16 15 3 3 3 13 2
31 13 4 12 9 1 11 3 1 12 2 9 12 1 15 2 3 15 4 1 9 13 0 9 7 3 4 3 13 0 9 2
21 11 11 2 15 9 13 2 13 2 16 4 0 9 1 11 13 13 3 1 9 2
12 9 0 11 4 1 0 9 13 13 0 9 2
16 0 11 3 13 13 3 0 0 9 7 13 9 0 0 9 2
21 1 11 4 15 1 15 13 13 9 7 9 2 10 0 9 4 13 3 10 9 2
17 9 1 15 14 12 0 9 4 0 11 13 1 9 0 0 9 2
22 3 13 3 3 13 1 15 2 16 4 0 10 9 13 9 1 10 9 2 13 11 2
13 3 4 13 1 12 9 1 11 13 14 12 9 2
13 9 1 15 4 1 9 11 2 11 13 13 11 2
9 9 1 11 11 2 9 11 7 11
13 9 9 0 11 7 9 9 15 4 13 1 11 2
22 3 3 1 9 0 11 2 7 14 1 0 0 9 1 11 2 1 15 15 13 9 2
12 10 9 4 3 13 2 13 4 15 7 13 2
16 9 7 14 9 0 0 0 9 4 3 13 7 10 0 9 2
18 3 15 13 13 1 9 15 7 13 13 14 15 2 15 3 3 13 2
10 9 9 9 0 9 4 13 13 0 2
6 9 13 1 0 9 2
19 9 1 11 3 14 4 1 0 9 13 7 1 10 9 1 11 13 13 2
3 2 11 2
4 11 13 9 9
3 1 0 9
2 11 2
35 9 9 9 2 0 9 9 0 9 2 9 0 0 9 1 9 9 13 1 0 9 3 0 0 9 0 9 2 15 13 13 0 9 9 2
8 3 15 13 9 11 11 11 2
48 9 3 13 1 9 9 1 0 9 1 9 13 9 2 3 0 9 7 0 0 0 9 2 0 9 1 0 9 0 9 2 3 4 9 1 10 9 7 0 0 9 13 9 1 9 0 9 2
5 11 13 9 9 11
3 1 0 9
5 11 2 11 2 2
25 0 9 9 3 0 0 9 11 2 11 2 11 2 11 2 1 0 9 0 9 13 9 0 9 2
29 1 9 0 0 9 9 0 9 11 11 11 13 9 2 16 4 13 9 7 9 0 9 2 15 15 0 9 13 2
21 15 0 9 4 13 4 1 11 13 0 9 9 2 15 13 1 9 9 0 9 2
21 10 9 4 15 13 13 9 1 9 15 2 15 13 9 1 9 7 9 9 9 2
8 0 9 13 9 1 9 0 2
25 13 7 13 2 16 0 9 7 15 13 1 9 9 1 0 7 0 11 2 13 15 1 9 11 2
7 9 13 1 9 2 9 3
5 11 2 11 2 2
26 1 9 13 0 11 11 2 2 15 3 13 13 9 9 1 9 9 1 0 9 1 0 9 1 11 2
20 9 15 13 13 10 9 2 15 15 1 9 13 3 7 15 15 13 13 9 2
23 16 9 1 0 9 3 13 1 9 2 3 13 12 9 0 0 9 2 15 15 13 13 2
20 12 1 15 15 13 3 2 16 0 9 13 1 0 9 7 13 9 1 9 2
8 0 9 1 9 9 13 9 2
14 9 12 9 13 3 0 7 4 15 13 1 0 9 2
7 9 9 1 9 15 13 2
5 0 9 13 0 9
6 0 11 2 11 2 2
34 16 9 0 9 9 9 9 1 11 1 11 2 15 15 13 12 2 9 2 13 9 1 0 11 9 9 1 9 1 12 1 12 9 2
26 15 1 0 9 12 0 9 13 1 9 0 9 7 0 9 15 13 1 9 3 2 16 13 1 9 2
26 16 3 15 0 9 13 1 0 9 7 13 15 13 9 12 9 9 2 13 15 9 0 1 9 9 2
29 7 3 2 16 9 9 1 9 3 4 13 0 9 2 15 15 13 1 9 2 9 15 13 7 1 9 9 13 2
19 1 9 0 9 13 9 12 1 9 9 2 16 4 13 1 9 1 9 2
8 0 9 4 13 3 0 9 2
2 9 13
6 0 11 2 11 2 2
22 12 11 7 12 11 13 1 9 1 0 9 12 9 7 13 15 1 9 1 9 11 2
24 12 13 0 9 1 9 2 0 13 1 9 10 9 2 3 15 13 13 0 9 1 12 9 2
7 16 9 15 13 0 11 2
13 0 9 15 13 9 11 2 10 9 15 9 13 2
6 9 15 13 1 9 2
2 0 13
6 0 11 2 11 2 2
24 1 9 1 12 9 13 1 9 2 12 0 9 9 11 2 11 2 15 13 9 0 9 11 2
9 0 9 7 3 13 3 12 9 2
9 9 15 13 1 9 9 0 9 2
3 9 1 9
5 11 2 11 2 2
15 1 0 9 9 2 11 15 13 9 0 9 9 0 9 2
10 12 1 9 9 13 9 7 0 13 2
11 9 15 13 13 12 9 7 12 9 9 2
7 0 9 11 4 13 0 9
2 11 2
15 1 11 1 11 1 11 4 13 0 0 9 0 9 11 2
58 0 9 11 11 13 2 16 9 2 15 4 13 12 9 2 4 13 12 1 15 0 9 2 0 9 1 0 9 7 1 9 0 7 0 9 2 15 13 9 11 2 7 0 0 9 11 2 15 4 13 1 0 9 1 9 10 9 2
11 0 9 4 13 7 16 0 9 9 11 2
10 12 9 4 13 0 9 1 0 9 2
10 13 3 10 9 1 9 3 12 9 2
27 10 0 9 13 9 0 9 9 11 2 15 13 1 10 9 9 3 1 9 7 9 2 13 11 2 11 2
16 11 13 10 9 9 14 1 11 2 7 7 1 11 7 11 2
11 1 15 13 0 7 16 0 7 0 9 2
4 9 13 1 11
7 11 1 11 2 11 2 2
23 1 9 4 13 1 9 0 11 2 11 2 1 11 2 9 9 12 0 9 1 0 11 2
31 12 2 9 1 0 9 0 9 2 1 9 2 3 9 13 9 11 2 13 10 0 9 1 9 2 1 15 1 15 13 2
9 9 15 13 12 9 7 12 9 2
14 13 15 3 0 9 2 7 9 3 0 9 13 0 2
39 13 1 0 9 2 16 9 13 4 13 1 9 9 9 1 9 1 12 9 1 12 9 2 13 3 9 11 0 9 0 9 9 1 11 1 11 11 11 2
14 9 1 9 0 9 13 2 16 9 13 1 9 1 0
5 11 2 11 2 2
18 0 9 13 1 12 0 9 3 0 1 9 1 0 0 9 11 11 2
24 0 11 2 11 2 15 13 0 9 9 2 13 1 0 9 1 0 9 9 1 11 2 11 2
13 1 9 13 12 2 9 3 1 11 9 1 11 2
19 11 2 0 1 9 1 0 11 2 13 9 1 9 7 13 1 9 9 2
20 1 9 1 9 13 0 9 12 9 2 15 11 2 11 13 0 9 1 9 2
25 16 13 0 9 0 9 11 2 11 2 9 3 2 13 2 16 1 9 7 9 13 10 0 9 2
14 11 4 1 9 13 1 9 2 10 9 13 1 9 2
7 1 11 13 0 9 9 2
13 1 0 0 9 13 3 0 12 0 9 1 11 2
30 0 11 11 2 15 4 1 9 15 13 1 0 0 9 2 13 12 2 12 9 0 2 0 9 7 13 0 0 9 2
20 0 11 11 13 12 2 12 9 0 2 0 9 7 13 3 0 3 0 9 2
14 1 0 9 13 13 9 9 12 9 2 15 3 13 2
17 9 4 15 13 13 1 0 9 11 1 0 0 9 9 12 12 2
13 9 13 2 16 12 1 0 13 1 9 0 9 2
17 10 9 1 0 9 13 9 13 1 0 0 9 7 1 9 12 2
5 9 15 13 1 9
2 0 9
5 11 2 11 2 2
32 1 9 0 9 1 9 0 9 2 15 15 13 13 12 2 12 2 1 9 9 11 2 15 13 9 9 0 9 13 1 9 2
22 9 9 13 2 16 4 13 1 9 13 9 9 1 10 9 7 13 1 10 9 9 2
16 10 9 13 13 3 9 15 2 15 13 13 9 0 0 9 2
16 1 15 13 9 0 11 9 1 10 9 7 9 1 9 11 2
8 9 2 3 13 2 15 13 2
15 0 9 13 9 9 2 3 3 11 2 11 13 13 0 2
1 9
19 0 9 1 11 2 3 0 1 0 9 1 11 11 2 4 1 9 13 2
20 9 4 1 9 13 2 3 15 7 13 2 16 13 3 2 7 3 3 13 2
31 1 9 13 3 12 9 2 7 13 0 2 16 15 3 13 3 13 2 13 11 1 9 9 0 9 0 9 9 11 11 2
3 2 11 2
1 9
25 9 11 13 3 0 9 1 9 1 9 9 1 9 11 0 9 2 15 9 4 13 1 12 9 2
3 2 11 2
4 9 1 0 9
1 9
2 11 11
32 9 1 9 9 0 9 1 9 9 13 10 9 15 13 2 16 4 4 13 1 10 10 9 1 9 9 0 9 1 9 12 2
12 9 15 13 1 9 1 9 9 2 15 13 2
10 9 2 11 11 2 0 9 9 11 2
7 9 2 12 2 9 12 2
6 3 0 9 0 9 2
49 1 15 2 15 11 2 11 13 2 15 13 2 1 10 9 15 9 11 13 1 10 0 7 0 9 1 0 9 2 16 15 3 1 9 0 9 13 11 7 1 15 3 15 9 13 10 0 9 2
7 3 3 9 11 3 13 2
16 3 15 13 7 13 10 9 2 16 4 0 9 13 3 0 2
9 9 1 9 11 4 7 3 13 2
38 3 1 15 13 13 9 0 0 9 2 16 3 3 13 10 0 0 9 2 7 0 7 0 9 0 9 11 7 0 0 9 11 2 15 3 15 13 2
15 9 7 4 13 1 0 9 1 10 9 2 13 1 15 2
6 9 9 11 13 13 0
1 9
2 11 11
25 9 0 0 9 13 1 0 9 12 0 9 2 0 9 9 2 11 2 2 9 9 7 9 9 2
31 9 9 0 9 4 13 3 13 15 9 0 1 9 7 0 9 12 0 0 9 2 9 1 0 9 0 7 9 1 9 2
37 10 12 9 3 9 11 11 11 2 15 13 3 9 9 9 2 13 16 9 1 9 1 9 0 9 7 12 1 15 3 1 0 9 13 0 9 2
22 10 9 1 0 9 3 13 9 1 10 9 7 9 1 9 11 13 3 10 0 9 2
19 13 1 9 2 16 9 11 15 13 3 13 9 9 9 1 0 0 9 2
23 13 15 3 9 9 9 2 15 13 9 1 9 3 0 0 9 0 9 7 3 7 9 2
28 7 15 7 3 2 16 0 9 9 2 12 1 9 12 13 3 2 16 13 9 9 2 13 3 13 15 0 2
18 1 10 9 13 16 13 2 16 9 13 0 0 9 1 0 9 9 2
26 16 13 0 13 9 9 11 2 3 3 15 13 13 0 2 16 10 0 9 13 1 10 9 3 9 2
7 9 0 9 2 9 0 9
2 11 11
22 13 14 0 9 2 3 4 9 0 9 13 3 3 16 1 9 2 3 1 0 9 2
28 3 15 0 0 9 0 1 9 13 3 10 9 2 7 0 9 4 13 1 0 9 3 14 1 12 1 15 2
16 13 0 2 16 4 15 10 0 9 1 0 9 3 3 13 2
7 9 13 10 2 15 0 2
8 1 0 9 13 0 13 9 2
21 15 15 3 3 13 1 0 9 9 2 7 13 15 3 3 2 3 13 0 9 2
15 9 0 9 2 15 13 0 9 2 15 13 3 0 9 2
18 16 13 0 9 2 13 7 0 9 13 1 9 7 9 0 9 9 2
20 3 2 0 9 9 2 15 0 9 15 0 9 13 2 15 3 13 1 9 2
9 3 3 3 9 13 2 0 13 2
10 7 1 10 0 9 4 13 13 9 2
19 13 4 3 0 13 2 7 0 3 3 13 2 2 16 9 13 9 9 2
32 7 16 9 9 0 9 4 13 1 12 1 0 2 0 2 9 9 2 13 3 1 9 0 0 9 9 13 2 13 7 13 2
17 13 2 14 3 0 15 13 2 3 14 9 0 0 9 0 9 2
9 1 9 4 13 13 1 12 9 2
17 3 15 13 2 16 0 9 15 3 13 1 0 9 9 0 9 2
13 9 15 9 9 13 3 0 9 9 9 9 11 2
44 13 15 2 10 0 9 13 0 0 9 13 2 16 15 13 9 2 9 9 13 0 9 1 12 1 12 0 9 2 9 12 9 13 9 9 0 3 2 7 13 15 9 9 2
14 3 12 9 0 9 13 7 13 1 0 2 0 9 2
7 9 13 7 13 12 9 2
7 15 13 1 11 9 9 2
34 10 9 12 9 13 3 0 9 9 1 9 2 9 9 0 9 2 9 9 7 9 1 0 9 2 9 9 1 9 9 3 2 2 2
12 0 9 9 9 1 9 1 9 7 3 13 2
15 9 9 13 13 12 9 2 15 3 3 13 9 9 11 2
19 0 9 3 3 13 2 13 1 15 0 9 9 7 12 9 13 0 9 2
11 15 3 13 12 9 13 10 0 0 9 2
26 16 15 13 1 9 9 2 14 12 7 12 9 4 3 13 2 7 2 9 13 3 7 3 0 9 2
4 13 15 15 2
5 15 13 0 13 2
4 3 0 9 2
17 13 0 15 13 2 16 4 15 13 13 3 0 2 0 7 0 2
17 0 9 15 3 13 7 0 9 15 4 13 13 2 16 3 13 2
21 3 0 9 9 0 9 13 0 7 2 3 13 0 0 9 2 3 7 0 9 2
16 0 0 9 4 3 13 0 9 2 3 1 0 9 7 9 2
25 10 0 9 1 0 9 13 1 15 2 9 12 9 9 2 3 3 9 1 0 9 1 9 2 2
17 9 2 15 13 13 9 9 9 0 1 9 2 13 9 9 9 2
8 13 15 15 1 12 9 9 2
9 9 0 1 9 0 13 0 9 2
31 13 0 2 16 0 1 15 1 0 9 1 0 9 3 4 13 13 7 3 2 16 10 0 9 13 13 1 0 12 9 2
32 9 3 3 13 1 9 9 2 0 9 2 2 7 3 4 1 0 9 13 2 3 15 13 3 2 0 9 2 9 2 2 2
6 1 9 13 0 9 2
24 16 4 7 3 1 9 13 1 0 9 9 2 13 4 15 9 9 9 9 1 0 9 13 2
26 1 0 9 4 13 3 3 13 7 13 4 15 13 15 9 1 9 0 0 9 9 2 9 7 9 2
5 9 1 9 9 13
2 11 11
14 9 2 15 13 1 11 2 3 13 9 1 10 9 2
10 0 0 9 15 13 1 9 1 9 2
10 15 7 0 0 13 9 0 9 9 2
14 7 3 1 0 9 9 7 0 9 15 13 9 11 2
14 1 9 13 3 9 12 2 9 1 11 7 10 9 2
18 9 13 9 1 9 11 2 3 15 1 9 13 7 9 1 9 9 2
10 9 13 7 1 9 2 7 1 9 2
13 10 9 13 10 9 9 2 13 9 9 11 11 2
14 9 1 9 15 13 3 1 12 7 3 1 12 9 2
18 1 9 13 13 0 9 2 15 9 1 9 13 2 7 15 15 13 2
25 9 15 13 1 9 9 13 2 7 3 13 0 13 3 9 0 1 9 2 13 1 9 3 9 2
13 0 13 0 9 1 9 2 1 12 12 9 3 2
18 0 9 2 15 9 3 13 2 13 9 1 11 1 12 12 9 3 2
25 3 13 1 12 9 10 9 9 2 3 13 10 9 1 0 9 12 2 12 2 13 11 2 11 2
14 13 9 9 2 15 13 1 10 0 9 9 1 11 2
20 9 13 1 10 9 13 9 7 1 9 2 3 13 9 9 7 9 13 0 2
27 9 15 13 2 3 0 9 2 1 10 9 11 2 1 10 9 2 1 10 9 7 1 15 15 13 13 2
22 1 9 3 13 7 9 2 15 15 1 10 9 3 13 2 7 9 1 12 0 9 2
16 15 13 2 16 9 13 3 1 0 9 11 7 13 0 3 2
23 9 13 13 9 7 3 2 7 1 0 9 15 13 3 13 1 9 9 1 9 0 9 2
33 13 0 0 9 16 0 0 9 2 15 1 9 13 2 16 1 9 9 1 9 14 12 0 9 15 1 0 9 13 15 13 9 2
27 1 10 9 4 0 9 13 13 7 9 2 16 1 0 9 13 0 13 9 2 7 4 13 0 9 13 2
9 10 0 9 9 7 9 3 13 2
16 1 10 9 15 10 9 3 13 1 9 2 13 11 2 11 2
10 1 9 9 7 9 1 9 9 13 2
27 1 9 2 16 1 11 16 9 13 9 9 1 0 9 9 2 13 10 9 9 1 9 12 9 0 9 2
20 16 9 11 13 9 1 0 9 9 9 2 13 9 1 9 12 9 0 9 2
10 9 13 3 2 16 13 15 0 9 2
13 10 9 7 13 9 9 1 0 9 7 9 9 2
15 10 9 13 1 0 9 9 0 9 2 13 11 2 11 2
5 9 1 11 2 11
5 11 2 11 2 2
14 0 9 1 0 0 9 13 9 0 9 9 7 9 2
24 1 9 12 2 9 0 0 9 13 9 11 1 9 9 9 9 11 7 0 9 9 11 11 2
18 16 0 13 11 2 15 0 9 13 1 0 7 0 9 0 1 11 2
44 1 9 11 15 3 13 2 16 11 13 9 7 10 9 1 0 9 13 12 9 2 16 1 9 12 13 2 1 10 0 9 9 9 2 9 9 9 9 1 9 9 7 9 2
8 9 13 1 9 7 0 9 2
20 10 9 11 11 13 2 16 1 9 4 13 13 9 1 9 2 7 14 9 2
5 0 9 7 1 11
2 11 2
28 9 9 13 0 9 0 9 2 15 1 9 11 2 0 9 7 0 0 11 3 13 7 3 13 15 12 9 2
12 11 3 9 13 16 12 1 12 0 0 9 2
24 1 9 15 13 1 0 13 1 0 2 0 2 0 9 0 9 7 13 3 13 0 0 9 2
20 1 12 0 9 13 0 9 13 0 9 2 7 3 13 0 0 9 1 9 2
27 0 9 4 15 13 13 0 0 0 9 7 0 9 1 0 7 0 9 2 15 13 1 9 0 0 9 2
16 12 1 9 13 3 9 0 0 9 1 0 11 1 0 11 2
5 11 13 9 0 9
2 11 2
10 0 9 13 13 3 13 1 9 9 2
28 1 0 9 4 15 13 3 0 9 2 7 13 4 15 0 9 0 9 2 13 3 0 9 11 11 9 11 2
32 3 4 13 2 16 9 4 13 3 2 13 7 13 2 16 9 9 13 13 9 12 9 7 13 0 9 1 15 7 0 11 2
13 13 3 2 16 9 9 9 1 11 15 3 13 2
6 13 15 9 1 11 2
23 11 15 13 1 9 9 1 9 9 1 10 9 2 16 10 9 4 1 11 13 1 0 2
9 13 3 0 11 9 1 0 9 2
41 1 9 9 1 12 1 12 0 9 15 13 2 16 1 9 2 15 13 13 11 1 0 2 0 9 1 11 7 0 11 3 1 9 2 15 13 3 12 9 0 2
22 1 9 13 9 9 0 9 11 1 0 11 2 9 2 1 9 9 9 1 0 9 2
9 9 13 1 9 9 1 9 9 2
9 7 13 15 14 0 9 1 11 2
20 13 1 15 13 7 9 9 0 1 0 2 9 0 9 2 11 2 1 11 2
16 11 13 0 9 2 16 9 11 11 12 2 13 0 9 11 2
13 1 9 1 9 0 11 15 13 0 9 11 11 2
20 9 4 1 11 13 13 12 2 9 2 7 13 9 1 10 9 7 0 9 2
16 9 0 11 11 11 3 13 2 16 0 9 1 11 13 13 2
19 13 15 9 15 2 15 13 9 1 9 7 9 2 13 0 0 9 11 2
16 9 15 2 15 3 13 1 15 2 15 13 11 2 13 9 2
5 0 9 13 10 9
10 9 9 11 11 11 13 0 9 1 11
2 11 11
31 0 9 13 9 2 3 13 3 0 0 9 0 11 7 13 15 3 9 1 9 0 9 1 10 9 2 9 0 0 9 2
38 0 9 13 0 9 13 0 9 0 1 9 0 9 9 0 9 7 9 0 9 2 13 0 9 9 11 11 2 15 13 1 0 9 1 0 9 11 2
37 0 9 13 9 1 3 0 9 9 1 0 9 7 11 2 13 11 2 7 13 0 9 14 0 2 7 3 0 9 7 9 1 9 9 0 9 2
19 3 1 9 0 9 2 3 10 9 1 11 15 0 1 9 0 9 13 2
22 3 13 1 0 9 9 2 15 13 1 9 1 11 0 0 9 2 9 9 11 11 2
42 1 10 9 13 9 0 9 2 16 4 16 9 1 10 2 16 0 9 3 13 11 3 3 0 9 0 9 2 13 13 1 0 9 0 9 2 13 11 1 0 9 2
11 3 1 9 11 13 0 9 2 13 0 2
21 0 9 3 13 2 16 3 4 9 0 9 1 11 13 1 0 9 1 12 9 2
31 7 13 0 9 2 16 7 3 1 9 11 11 13 1 11 0 9 1 9 2 0 9 2 9 7 9 9 0 9 0 2
16 3 13 9 2 16 0 9 13 1 10 9 1 11 3 3 2
8 1 9 9 11 11 3 14 2
27 0 9 13 3 3 9 11 2 15 15 1 0 9 1 0 9 0 9 15 1 15 3 13 1 0 9 2
6 11 11 0 9 13 2
10 10 0 9 13 3 1 9 1 9 2
15 3 3 3 13 9 0 0 9 1 9 3 12 9 9 2
31 3 15 15 13 13 9 0 2 0 9 1 0 9 2 15 4 13 1 9 3 1 9 1 9 1 0 9 9 0 9 2
21 9 1 3 3 0 0 2 0 9 4 13 13 9 7 0 9 11 11 1 11 2
21 0 9 15 1 9 13 1 0 0 9 1 11 1 10 0 9 11 11 2 11 2
29 16 3 13 1 0 9 1 12 9 1 9 2 13 0 2 16 1 11 13 0 9 0 2 0 9 1 0 9 2
19 3 1 10 9 0 9 13 9 1 0 9 2 15 4 1 11 3 13 2
18 0 9 15 15 2 1 15 2 15 1 0 0 9 13 2 13 13 2
19 0 9 10 9 13 7 13 3 2 3 0 13 13 15 10 9 1 9 2
19 15 0 13 13 0 9 10 9 1 9 0 9 2 15 13 1 11 13 2
25 1 9 15 3 13 2 16 0 9 4 13 13 1 15 2 16 10 0 9 13 1 9 9 9 2
14 16 15 15 15 13 13 2 3 11 10 9 9 13 2
24 16 14 2 13 9 1 9 0 9 0 0 9 3 1 9 0 9 7 10 9 9 11 11 2
5 0 0 9 13 11
2 11 2
24 0 14 9 0 9 3 1 9 1 11 2 11 3 13 0 9 2 15 15 3 13 1 11 2
29 0 9 0 0 9 9 13 1 12 9 1 0 9 11 1 9 0 11 2 3 9 11 13 1 0 9 11 11 2
9 0 9 13 1 11 3 3 3 2
19 0 9 11 11 2 15 13 1 0 11 2 4 1 11 13 1 0 9 2
22 10 9 13 13 9 0 2 0 9 1 11 7 9 7 3 9 11 1 9 0 9 2
28 0 9 3 13 0 9 1 15 2 15 15 13 2 16 1 9 0 9 1 11 13 11 1 9 1 11 9 2
24 3 0 9 0 9 1 0 9 4 3 13 1 9 0 9 2 13 11 1 9 1 9 11 2
13 13 2 16 1 11 7 11 13 10 0 0 9 2
19 11 7 11 3 13 9 7 9 7 1 10 9 15 13 9 2 13 9 2
10 9 9 0 9 1 11 13 0 9 2
31 9 7 9 9 0 0 9 13 2 16 0 9 15 13 1 0 9 1 11 13 1 0 9 1 11 2 3 15 15 13 2
8 13 15 3 0 9 0 11 2
16 11 13 9 10 9 1 12 9 7 11 0 9 13 12 9 2
9 7 15 9 9 9 1 12 9 2
13 15 13 0 9 2 15 13 3 9 2 13 9 2
4 0 9 13 11
2 11 2
27 0 9 1 11 3 13 9 1 9 11 2 16 13 1 9 2 4 2 14 11 1 0 9 13 0 9 2
25 9 13 0 9 9 2 11 2 2 10 9 1 9 1 9 12 13 1 11 0 9 9 7 9 2
20 11 3 3 13 10 0 9 1 11 2 16 1 10 0 9 13 9 0 9 2
24 1 0 0 9 1 11 9 9 13 0 9 1 9 9 7 3 15 3 13 0 9 1 9 2
13 0 0 9 13 2 16 0 9 1 11 3 13 2
13 9 11 4 3 13 1 0 9 2 3 4 13 2
5 9 11 13 1 9
2 11 2
21 0 9 11 11 4 3 13 9 0 9 2 15 4 13 9 9 1 0 0 9 2
8 10 9 13 1 0 9 9 2
18 13 15 1 0 0 9 1 9 9 1 9 7 0 9 1 9 9 2
17 0 0 9 11 11 11 13 9 0 1 15 1 0 9 9 9 2
25 11 13 2 16 9 0 9 1 0 9 2 15 13 1 9 10 9 0 2 4 13 1 9 9 2
11 10 9 14 4 13 1 9 9 7 9 2
16 1 9 11 13 3 0 9 9 9 2 15 13 0 0 9 2
15 1 9 13 9 1 9 9 9 12 9 1 0 0 9 2
2 9 11
22 1 0 9 1 9 15 13 12 9 3 16 9 1 9 2 13 2 9 7 0 9 2
9 16 9 10 9 13 2 13 15 2
2 9 9
13 0 9 11 13 11 7 13 1 0 9 1 11 2
28 13 15 2 16 1 1 0 9 11 1 0 0 9 9 13 1 9 9 9 11 1 11 2 15 13 9 9 2
9 1 9 9 13 9 7 1 11 2
2 9 11
1 3
49 0 9 1 9 0 9 1 9 2 6 2 2 15 13 1 9 0 11 1 0 9 2 3 13 2 16 0 9 1 9 0 0 9 2 11 2 13 9 1 9 7 16 3 13 9 1 0 9 2
10 11 3 13 1 9 12 1 0 9 2
27 13 3 1 9 0 9 2 15 9 3 13 1 9 12 1 9 0 0 9 1 11 7 13 15 1 9 2
25 9 0 9 0 9 7 9 11 11 4 3 13 10 9 1 9 2 16 13 1 10 9 1 11 2
6 1 9 15 3 13 2
9 11 3 13 9 10 9 1 11 2
29 13 15 1 9 1 9 0 2 0 9 2 15 13 9 9 1 9 0 9 2 9 9 0 9 9 9 11 11 2
29 9 0 9 1 0 0 0 9 15 3 3 13 1 9 0 9 0 0 9 2 15 4 13 1 9 0 0 9 2
11 13 15 0 9 11 1 11 11 11 11 2
17 0 9 13 1 9 11 1 11 13 9 2 15 13 10 0 9 2
20 9 15 13 1 10 9 2 15 13 1 9 2 7 13 15 1 9 7 9 2
14 16 15 9 9 13 3 2 9 3 13 1 0 9 2
18 11 11 2 9 0 9 0 9 2 15 3 13 9 0 9 1 9 2
5 9 11 11 2 11
6 0 9 0 7 1 9
14 0 9 13 1 0 0 9 1 0 9 0 0 9 2
49 1 9 9 12 9 9 2 0 1 9 9 2 15 3 3 13 0 9 0 9 2 12 9 9 2 2 0 9 11 11 2 12 9 2 7 0 9 0 2 12 9 2 2 0 7 1 10 9 2
32 1 9 13 0 9 1 11 11 1 9 0 9 2 12 9 2 7 9 0 9 2 12 9 2 2 15 1 0 9 13 3 2
32 1 0 9 15 0 9 13 0 9 9 2 3 12 9 9 2 7 9 0 9 2 15 1 0 12 9 1 9 13 12 9 2
27 1 9 13 9 0 0 9 9 2 16 4 9 13 3 9 2 7 16 15 1 9 1 10 9 13 3 2
17 0 9 13 0 9 7 9 0 9 2 16 15 0 9 3 13 2
6 9 13 7 0 9 2
33 0 9 0 13 3 3 13 3 9 1 9 2 9 0 11 7 1 0 9 13 3 10 9 0 7 0 2 15 13 7 9 0 2
24 9 0 9 1 9 0 15 3 3 13 1 9 0 9 11 2 15 1 9 13 7 9 9 2
5 2 11 2 11 2
4 12 0 0 9
13 0 0 9 12 0 9 13 10 9 9 0 9 2
30 9 1 11 11 11 1 9 11 11 7 12 9 2 11 11 2 11 11 1 9 11 11 3 13 1 3 0 0 9 2
18 4 7 3 13 2 13 0 7 0 9 2 13 9 7 13 0 9 2
16 0 9 0 9 0 1 0 9 12 9 13 13 1 12 9 2
17 3 0 9 11 11 2 12 2 9 10 13 13 0 9 10 9 2
17 13 4 3 7 10 0 9 2 7 7 0 9 1 9 11 11 2
3 2 11 2
5 12 9 7 12 9
1 9
2 11 11
12 1 0 9 9 11 15 3 13 1 0 9 2
10 1 0 9 13 0 0 9 0 9 2
21 3 0 9 15 1 10 9 13 3 9 9 10 0 9 1 0 9 1 9 12 2
14 0 9 13 0 0 9 7 0 9 3 13 0 9 2
16 1 11 1 11 13 13 0 0 9 0 0 9 9 10 9 2
25 0 9 2 15 1 0 9 13 0 9 11 11 2 9 0 11 2 2 15 3 13 13 3 3 2
18 9 9 0 9 2 0 9 3 9 2 13 13 12 3 15 0 9 2
19 0 9 0 7 0 9 13 1 15 2 16 9 10 0 9 13 1 9 2
13 9 0 7 0 9 1 0 9 15 13 0 11 2
10 3 4 3 13 13 3 12 9 3 2
21 16 7 9 9 13 0 9 3 2 13 13 9 3 0 2 15 4 13 9 15 2
16 9 2 16 4 0 9 13 9 0 7 0 2 13 3 0 2
19 1 0 9 7 3 13 9 12 0 9 2 15 4 15 7 13 3 13 2
12 2 0 9 9 13 9 9 9 7 10 9 2
13 1 9 0 2 0 15 1 9 13 3 11 2 2
17 1 9 9 1 9 0 9 15 13 0 9 2 9 1 15 0 2
17 3 15 9 13 1 9 9 2 1 15 13 10 9 0 9 9 2
20 9 2 7 9 0 9 2 7 4 3 13 7 3 4 3 13 13 9 0 2
21 16 0 9 3 10 9 13 7 13 2 1 0 9 15 4 10 9 13 0 9 2
10 9 9 4 15 13 13 1 9 9 2
24 1 1 9 9 7 13 3 0 2 16 4 15 9 12 9 1 0 9 1 9 3 14 13 2
5 0 0 9 0 11
18 1 0 0 9 15 9 1 9 1 0 9 13 7 0 9 0 11 2
33 9 0 9 15 13 2 3 1 0 0 11 7 0 11 2 1 0 9 3 3 0 0 0 9 2 15 13 7 9 0 0 9 2
17 0 0 9 11 2 12 2 15 0 11 3 13 1 0 9 9 2
22 9 3 13 3 0 9 11 11 7 14 3 0 2 3 0 9 9 9 11 7 11 2
13 15 3 13 13 0 9 9 2 3 0 0 9 2
38 0 12 3 0 9 2 0 11 3 2 12 2 7 11 1 0 11 2 12 2 2 7 3 10 9 7 9 0 9 7 13 0 9 3 3 14 13 2
17 1 15 0 9 13 1 9 3 3 3 2 16 15 1 15 13 2
29 3 15 7 0 11 13 0 9 0 11 2 15 13 3 0 0 9 1 0 0 9 9 0 7 9 9 9 0 2
24 7 16 9 0 11 13 2 1 0 11 9 13 13 0 0 9 2 9 1 9 7 9 0 2
3 2 11 2
1 3
24 12 0 9 13 13 1 11 1 12 2 7 12 2 9 1 9 12 2 9 0 9 11 12 2
21 3 1 0 9 0 9 13 0 0 9 11 0 2 3 0 0 9 11 0 9 2
5 9 13 1 12 2
21 0 9 3 13 4 7 1 0 9 3 7 13 2 13 11 9 9 11 11 11 2
25 0 9 9 2 13 1 9 0 9 2 13 3 1 9 0 9 9 2 15 1 10 9 13 9 2
12 9 9 13 7 0 9 2 15 4 9 13 2
8 1 11 4 1 9 13 9 2
3 2 11 2
6 9 9 7 9 13 0
2 11 11
16 1 9 0 2 0 15 9 2 15 13 7 0 2 0 9 2
18 15 13 9 9 9 9 1 0 9 7 13 13 0 9 1 9 9 2
20 16 3 13 9 0 9 2 3 15 13 1 9 9 2 9 2 9 7 9 2
14 0 9 12 2 9 12 13 12 9 1 15 12 9 2
12 1 9 9 13 1 3 0 9 1 12 9 2
16 1 9 0 9 15 7 9 9 13 13 1 0 12 9 3 2
20 3 12 2 9 13 12 9 2 16 9 9 9 13 12 7 9 13 12 9 2
17 15 4 13 3 9 2 15 13 9 3 0 0 9 1 0 9 2
20 7 0 9 13 1 10 9 9 12 9 2 11 12 7 0 9 3 12 9 2
18 1 9 13 9 9 12 12 9 7 0 12 9 4 13 12 2 9 2
18 1 10 9 9 9 3 13 0 9 2 12 2 7 9 13 12 9 2
16 9 2 15 13 9 1 9 0 9 2 7 3 13 3 9 2
22 3 12 2 9 13 10 0 9 9 12 9 2 7 3 1 9 13 9 9 9 0 2
19 1 9 2 16 15 12 13 2 0 15 13 2 15 3 3 13 9 9 2
23 15 15 3 13 1 9 10 12 9 2 7 13 15 7 1 0 9 9 9 13 1 9 2
14 3 3 15 13 7 9 9 2 15 13 13 0 9 2
14 9 9 15 13 3 1 12 9 7 13 3 0 9 2
5 15 2 3 2 3
28 9 9 2 9 2 9 7 9 11 11 1 9 12 2 12 4 13 3 1 0 9 7 13 1 12 2 9 2
18 11 0 13 3 1 0 9 15 0 1 12 9 1 9 9 9 9 2
16 9 9 0 9 13 13 1 0 9 1 11 1 12 2 9 2
12 3 4 13 9 9 11 11 1 9 0 9 2
7 9 13 1 12 2 9 2
31 9 11 11 11 11 12 2 13 1 9 0 1 0 9 11 1 9 0 2 11 2 0 9 2 7 13 1 12 2 9 2
5 0 9 9 1 11
24 9 1 11 15 1 10 9 1 9 12 13 1 9 9 3 12 9 0 0 9 1 0 9 2
33 9 9 2 15 13 9 9 2 1 10 9 15 0 9 13 2 15 1 9 13 3 2 16 1 9 1 9 9 13 9 11 9 2
28 9 1 11 3 1 9 13 9 1 9 0 9 2 15 0 9 2 9 2 9 2 4 13 13 7 0 9 2
18 13 4 15 3 13 9 1 9 2 7 15 7 9 2 7 0 9 2
18 0 9 9 1 11 15 3 13 11 9 2 9 12 1 0 0 9 2
17 1 9 13 9 9 1 11 11 11 2 15 13 1 9 0 9 2
5 2 11 2 11 2
5 9 0 9 13 9
15 0 9 9 9 9 3 1 0 0 9 13 9 0 9 2
20 13 15 15 7 9 11 1 9 9 9 1 11 1 11 2 15 0 9 13 2
25 13 15 1 0 9 2 9 2 9 7 9 2 1 10 9 15 13 0 9 13 3 0 0 9 2
7 0 13 3 15 9 9 2
21 9 13 1 9 2 9 7 0 0 9 2 13 11 9 0 9 1 11 11 11 2
17 9 4 13 1 12 2 9 2 3 13 1 11 7 0 0 9 2
3 2 11 2
9 1 11 3 13 0 9 1 0 9
21 0 9 0 9 9 9 11 11 13 3 3 12 2 9 0 0 9 1 0 11 2
25 9 11 4 9 12 1 0 0 9 13 1 12 2 9 2 3 9 13 9 0 9 7 0 9 2
33 1 0 9 15 13 13 3 0 9 9 7 0 9 9 11 11 0 9 11 11 2 1 0 0 9 9 9 4 13 0 9 12 2
22 1 0 9 2 15 3 13 9 9 1 11 2 4 9 0 9 13 1 10 9 0 2
27 9 0 9 13 0 9 11 11 2 0 1 10 9 3 1 9 2 9 0 9 13 1 0 9 0 9 2
25 0 9 4 3 13 0 9 11 11 2 12 2 12 2 7 13 0 9 13 10 9 0 7 0 2
3 2 11 2
4 6 11 1 15
1 9
2 11 11
38 1 0 15 9 6 11 1 11 15 1 9 0 9 0 9 13 0 9 9 2 15 9 13 15 2 15 14 3 4 1 15 1 9 1 10 9 13 2
23 0 9 1 0 0 9 1 9 13 3 12 9 2 7 15 1 10 9 3 1 15 9 2
60 1 9 11 13 0 9 2 0 9 1 9 0 9 9 0 0 11 2 9 9 3 13 0 9 1 9 9 1 11 7 3 3 3 13 0 9 2 1 9 1 9 2 2 15 4 1 9 13 3 12 0 9 0 9 2 7 7 9 2 2
16 3 3 0 7 0 13 1 9 9 2 9 3 16 0 9 2
13 0 9 15 13 7 9 11 11 9 0 6 11 2
25 10 9 13 3 3 0 9 2 7 16 12 1 10 9 13 0 9 1 9 13 7 13 10 9 2
24 1 15 13 11 10 9 2 16 13 13 7 9 9 2 15 4 9 13 1 9 9 6 11 2
50 1 1 15 2 16 11 13 1 9 1 3 0 7 3 3 0 9 0 9 2 13 10 9 3 0 2 3 0 7 0 9 2 15 1 0 12 9 9 13 7 3 0 9 1 9 9 0 6 11 2
13 0 9 13 13 9 11 2 15 9 1 15 13 2
21 10 9 3 13 1 12 9 7 0 0 9 1 10 9 13 9 9 1 9 0 2
14 13 1 15 7 3 0 9 1 0 9 0 0 11 2
32 7 3 15 0 9 1 9 9 13 13 3 0 9 2 16 15 13 1 0 7 0 9 2 15 14 3 1 10 0 9 13 2
19 9 1 9 4 15 13 2 16 4 9 13 9 0 9 1 0 9 9 2
4 15 15 13 2
6 11 9 13 2 7 13
2 11 11
20 9 11 11 2 12 2 13 1 15 2 15 13 2 7 3 1 0 9 9 2
17 7 13 7 1 0 9 0 9 0 9 9 2 15 13 3 11 2
22 3 4 13 9 0 0 9 1 10 0 9 11 1 11 2 13 1 12 2 9 2 2
10 0 9 0 9 13 9 1 9 9 2
21 9 2 9 2 9 2 9 1 9 2 9 2 9 2 9 2 0 9 7 9 2
26 9 1 9 13 13 9 2 0 9 0 9 2 0 9 2 9 10 9 2 9 2 9 0 1 9 2
12 0 9 13 1 0 16 9 9 2 13 11 2
12 9 3 13 0 9 16 10 2 1 15 13 2
12 9 13 10 9 2 16 13 4 13 10 9 2
18 9 1 9 1 10 9 13 3 1 11 2 1 10 9 3 1 11 2
27 16 15 13 2 9 1 9 13 3 1 0 9 0 9 2 10 9 13 9 0 9 2 7 0 9 9 2
12 9 0 13 3 0 9 9 9 7 10 9 2
19 9 0 9 15 3 13 2 9 13 0 9 2 0 9 3 13 0 9 2
15 9 9 3 13 2 13 15 15 13 15 9 2 13 11 2
15 9 15 1 15 13 9 2 0 9 9 13 0 16 9 2
19 1 10 0 9 15 13 3 1 9 2 3 7 2 16 15 3 3 13 2
10 9 3 13 13 1 9 2 7 0 2
14 11 13 0 2 16 4 15 13 13 1 9 0 9 2
12 9 15 13 9 16 15 1 15 2 13 11 2
16 13 15 2 16 13 0 10 9 13 2 0 13 13 0 9 2
11 3 0 13 13 1 0 0 9 0 9 2
20 0 9 7 9 15 13 2 7 15 15 1 9 13 2 14 15 13 0 9 2
12 9 1 0 9 2 15 13 14 9 1 15 2
7 9 1 9 13 9 9 2
15 9 3 13 2 16 9 13 1 15 7 15 15 15 13 2
21 11 9 13 7 9 2 13 15 13 1 0 9 2 1 9 2 15 13 0 13 2
4 13 15 13 2
4 3 1 9 9
40 0 9 1 0 9 0 9 3 13 7 12 0 0 9 2 9 1 9 0 7 9 9 2 9 7 9 2 13 15 2 13 1 9 7 9 7 3 7 9 2
16 16 4 15 13 2 9 1 9 15 13 13 7 13 9 9 2
7 7 15 3 3 13 9 2
11 3 13 9 9 2 7 15 9 3 0 2
16 9 9 13 1 0 9 3 0 2 7 9 9 3 3 0 2
8 0 13 3 2 15 2 16 2
7 3 1 15 9 9 13 2
21 1 0 9 15 3 3 0 9 13 1 9 2 0 2 9 2 9 2 9 3 2
15 10 9 13 9 2 13 15 1 0 9 3 1 9 9 2
15 1 0 9 9 13 14 1 9 0 9 1 12 2 9 2
29 3 15 3 13 2 16 0 9 9 1 9 9 0 9 13 3 0 2 16 15 15 13 2 16 4 13 3 3 2
12 15 15 14 13 3 9 1 0 9 0 9 2
7 15 4 15 13 0 9 2
14 1 0 9 15 3 13 13 1 13 2 13 1 13 2
32 13 4 15 3 13 2 16 3 13 13 1 12 2 9 12 7 12 1 0 12 7 12 7 1 9 13 3 1 9 1 9 2
13 7 3 1 15 4 13 9 9 1 9 0 13 2
25 13 4 13 1 0 9 7 0 9 0 7 0 9 7 9 0 9 2 16 10 0 9 3 13 2
12 7 15 13 3 0 9 2 0 13 13 9 2
28 13 7 3 0 2 16 4 15 2 15 13 3 0 9 9 2 13 1 9 9 2 16 15 3 13 1 9 2
10 7 16 4 0 9 10 9 9 13 2
6 1 9 11 11 2 11
8 3 9 13 9 14 1 9 2
5 13 4 15 1 15
26 10 0 9 15 13 2 16 1 12 2 12 2 15 4 13 9 1 9 2 15 13 13 1 9 9 2
5 9 15 3 13 2
9 9 15 7 4 13 1 0 9 2
5 1 15 13 13 2
21 13 1 0 9 2 15 13 13 9 9 7 13 14 13 2 16 15 15 9 13 2
6 2 11 11 2 11 2
13 13 9 2 11 11 2 9 9 9 1 9 9 2
24 9 9 13 9 2 15 13 9 14 9 2 7 7 0 9 2 10 9 13 13 9 1 9 2
17 9 15 13 7 1 9 2 3 7 10 0 9 9 1 9 13 2
22 4 3 13 7 1 0 9 2 7 1 0 9 9 2 15 13 3 1 0 0 9 2
35 13 0 9 2 16 0 9 9 0 9 1 0 9 4 1 15 2 1 9 1 9 2 0 9 13 2 7 16 7 10 9 10 9 13 2
21 1 15 9 9 13 2 7 13 15 3 15 2 15 15 13 1 9 0 9 13 2
11 0 9 13 9 1 9 14 13 7 3 2
28 13 2 14 15 7 15 9 9 1 9 2 15 13 1 9 9 13 2 3 13 13 2 16 9 4 3 13 2
16 1 9 9 3 13 1 0 9 2 7 1 9 0 0 9 2
23 1 9 15 9 1 10 9 13 3 2 13 2 14 9 1 9 13 2 9 15 13 13 2
21 1 15 15 9 13 9 0 15 0 3 3 13 2 10 9 15 13 1 9 9 2
12 13 7 1 9 0 7 0 2 15 3 13 2
16 0 9 13 9 1 9 7 0 9 2 15 3 9 15 13 2
38 3 4 13 13 9 9 7 15 0 13 2 13 14 0 0 9 2 14 15 1 9 1 9 2 2 13 15 1 9 1 15 2 15 13 3 3 3 2
6 1 0 9 9 13 9
3 9 1 0
2 11 11
21 0 1 15 15 13 13 2 16 1 10 0 2 0 7 3 0 9 15 13 3 2
13 1 10 9 13 0 13 2 10 9 15 13 13 2
15 1 0 0 9 1 9 9 0 9 9 13 9 1 9 2
15 1 9 1 0 9 9 3 13 10 9 0 9 1 9 2
19 13 1 9 0 9 2 16 9 1 9 1 9 7 10 9 13 1 9 2
48 15 13 2 16 16 9 1 9 9 9 13 2 13 9 9 2 0 2 9 2 9 3 2 2 1 10 9 2 16 15 13 13 2 7 9 9 2 0 2 9 2 9 3 2 2 9 13 2
16 15 13 9 9 0 15 3 1 9 9 9 1 9 1 9 2
38 9 9 13 1 9 2 3 13 10 9 1 0 9 2 7 2 1 9 2 3 13 0 0 9 2 16 15 1 15 13 2 7 13 1 9 0 9 2
7 9 9 9 9 13 0 2
14 9 1 9 9 15 3 13 7 1 9 3 0 9 2
9 13 3 7 9 0 2 0 9 2
11 9 9 1 9 1 9 13 7 3 13 2
8 13 13 7 0 1 9 9 2
10 1 0 13 2 16 13 13 12 9 2
15 1 0 13 1 9 2 16 9 9 1 9 4 13 9 2
13 13 7 0 13 1 10 9 2 16 15 9 13 2
6 13 7 1 9 0 2
20 15 15 13 0 9 9 2 13 13 9 0 0 9 2 9 12 0 9 2 2
9 9 0 0 9 13 3 3 0 2
19 1 9 1 9 13 9 3 1 9 12 9 2 12 2 1 15 13 3 2
18 1 0 9 15 13 1 9 2 3 9 13 9 1 9 9 1 9 2
15 1 10 9 15 13 0 9 9 12 9 2 12 0 9 2
27 1 15 13 9 0 13 9 9 1 9 1 9 1 12 9 0 2 16 13 0 9 9 1 9 0 9 2
23 1 1 0 0 9 0 9 1 0 9 15 1 9 10 9 13 9 9 1 9 9 9 2
17 9 0 1 9 13 9 9 9 2 1 10 9 13 0 9 9 2
33 16 4 0 0 9 9 1 9 9 9 13 0 9 1 9 2 15 4 13 1 10 9 2 13 1 9 13 9 1 9 9 9 2
10 10 9 13 9 9 12 9 2 12 2
5 0 9 2 2 2
8 2 11 12 2 12 2 12 2
26 13 0 7 0 9 2 3 4 7 0 15 13 7 0 9 2 7 7 10 9 0 0 9 0 9 2
22 1 0 0 9 10 9 9 15 13 14 1 0 2 7 1 0 9 9 3 1 0 2
41 0 9 4 13 13 2 16 13 13 3 9 10 9 9 2 13 2 16 9 3 0 7 0 2 0 9 2 7 3 3 13 7 13 9 7 0 9 13 3 3 2
33 16 7 13 9 3 9 15 2 16 15 13 2 10 9 13 10 0 9 3 0 9 10 9 1 0 0 9 2 13 15 13 0 2
20 13 4 15 3 13 9 0 9 0 9 7 13 0 9 1 9 9 10 9 2
22 9 4 13 13 9 0 0 9 1 9 0 9 9 1 0 9 2 3 9 0 9 2
26 3 0 12 0 0 9 7 9 1 15 0 4 13 1 0 9 10 0 9 1 10 9 1 9 9 2
6 1 9 11 11 2 11
6 11 7 9 2 15 13
2 11 2
11 0 9 13 1 0 9 0 0 9 11 2
25 1 9 15 1 9 13 11 1 11 2 11 1 11 0 2 2 11 1 11 11 7 11 1 11 2
6 9 13 2 13 15 3
5 11 2 11 2 2
33 3 9 13 9 0 9 2 15 13 13 12 9 1 9 11 11 1 11 7 1 11 2 7 15 15 13 0 9 1 0 0 9 2
29 1 9 9 11 9 11 11 11 15 9 1 9 13 2 16 1 0 9 1 0 0 9 1 11 1 0 9 13 2
11 1 0 9 4 7 1 9 9 3 13 2
3 0 9 11
7 0 9 3 1 0 9 9
5 11 2 11 2 2
24 0 0 9 3 13 1 0 9 11 11 2 11 2 12 2 12 2 0 9 0 12 2 9 2
28 10 9 15 7 3 13 9 1 0 9 2 15 3 13 11 3 1 0 9 2 7 1 9 9 13 0 9 2
29 0 9 1 0 13 13 3 14 15 2 16 15 15 1 12 2 9 13 13 0 2 11 3 0 9 1 0 9 2
25 1 0 9 15 1 0 9 13 0 11 2 15 12 9 13 9 10 9 1 9 1 11 2 11 2
15 3 0 13 0 11 2 15 13 9 1 0 9 1 11 2
14 14 0 9 13 0 9 1 10 9 0 11 1 11 2
4 9 2 11 2
2 11 2
4 9 2 11 2
4 9 2 11 2
6 11 1 0 2 9 2
4 9 2 11 2
10 9 9 11 1 12 1 11 13 9 11
5 9 11 11 2 11
6 11 15 13 7 13 11
6 9 11 15 13 1 11
6 0 9 0 11 3 9
2 11 2
33 0 0 12 9 12 2 9 0 0 9 2 11 2 11 2 12 9 2 11 2 11 2 12 9 2 3 13 9 1 9 0 9 2
24 0 11 3 13 3 3 9 1 0 11 2 15 1 9 0 9 9 13 10 0 0 0 9 2
28 0 9 1 15 13 9 12 9 11 2 15 3 1 9 1 9 11 13 1 11 7 3 15 13 3 0 9 2
11 11 13 1 9 12 9 1 9 0 9 2
18 11 11 13 3 3 14 1 9 11 2 7 7 10 9 13 9 11 2
22 1 9 9 11 13 11 12 9 2 7 13 2 7 1 15 7 10 9 2 9 11 2
17 15 1 0 9 1 9 7 3 7 0 9 13 1 12 2 9 2
30 11 15 13 1 9 1 9 7 15 15 3 13 2 13 0 9 2 15 13 10 9 1 0 9 9 1 11 1 11 2
6 11 2 11 12 2 12
13 16 0 9 13 2 3 13 2 16 15 9 13 2
22 13 15 9 1 12 2 9 2 3 11 13 0 9 1 12 9 1 9 9 9 11 2
14 11 13 9 3 2 1 9 11 13 1 9 0 11 2
11 11 13 0 0 9 2 7 15 3 13 2
14 13 15 7 11 3 1 9 2 16 13 15 1 11 2
13 3 1 12 2 9 13 0 1 11 7 9 13 2
15 7 1 0 9 0 13 2 7 9 11 13 7 0 9 2
4 9 2 11 2
23 11 2 11 2 9 11 2 13 13 9 2 13 15 3 16 9 7 13 1 9 10 9 2
12 11 2 11 2 9 11 2 12 9 13 13 2
8 15 9 13 2 13 15 3 2
9 2 11 2 11 2 11 12 2 12
12 0 3 3 13 9 1 0 7 0 9 9 2
17 3 12 9 1 9 1 9 11 13 11 2 15 13 11 0 9 2
15 11 1 10 9 13 3 1 9 2 7 10 9 13 0 2
4 9 2 11 2
22 11 2 11 2 9 11 2 1 9 11 1 0 9 13 9 2 13 4 9 1 9 2
21 11 2 11 2 9 11 2 0 9 15 13 3 3 2 16 16 4 13 12 9 2
8 11 2 0 2 11 12 2 12
11 0 0 9 13 11 14 1 12 2 9 2
14 11 13 11 2 7 15 1 9 9 3 13 1 9 2
7 9 13 9 11 7 11 2
16 3 1 9 1 9 13 11 3 3 9 1 0 9 1 9 2
5 0 9 13 9 2
22 13 15 3 12 9 2 16 11 1 0 9 13 1 9 9 9 11 2 12 2 12 2
12 1 0 12 9 13 12 9 9 1 9 9 2
11 11 13 11 7 15 13 1 12 2 12 2
19 9 11 13 11 2 15 1 0 9 13 9 11 7 13 1 12 2 12 2
15 9 0 9 0 7 1 9 9 11 13 0 9 11 3 2
26 1 12 2 9 4 1 0 0 9 13 0 11 2 7 1 12 9 15 13 11 1 9 1 0 11 2
4 9 2 11 2
24 11 2 11 2 9 0 2 11 2 3 4 13 2 16 15 1 11 13 9 7 16 13 9 2
16 11 2 11 2 9 11 2 1 0 9 9 4 15 3 13 2
13 14 15 10 9 15 13 3 2 3 4 15 13 2
9 2 11 2 11 2 11 12 2 12
9 0 9 13 0 9 14 1 9 2
12 0 15 13 1 9 2 13 15 7 9 11 2
20 0 15 7 7 1 12 0 13 2 7 7 12 9 1 9 15 13 3 11 2
4 9 2 11 2
5 11 1 0 0 2
14 11 2 11 2 11 2 11 13 3 2 7 16 3 2
16 7 16 4 13 1 12 2 13 4 14 0 9 1 9 11 2
23 11 2 11 2 11 2 13 0 2 16 4 7 1 12 13 9 2 13 9 11 7 13 2
6 11 2 11 12 2 12
18 9 3 13 12 9 11 7 11 2 7 15 13 1 0 12 9 15 2
18 1 12 2 9 13 9 1 9 0 11 2 15 13 0 9 1 11 2
17 3 1 9 0 9 0 11 13 1 9 9 9 1 12 2 12 2
19 9 13 9 7 1 12 2 9 15 15 13 9 11 13 1 12 2 12 2
13 9 13 1 12 2 9 11 2 15 13 9 11 2
16 0 7 3 13 2 7 1 0 9 9 7 11 15 11 13 2
4 9 2 11 2
16 11 2 11 2 9 11 2 0 13 1 9 7 9 15 13 2
14 11 2 11 2 9 11 2 13 13 1 12 0 11 2
6 10 0 9 13 11 2
7 11 2 11 11 12 2 12
6 0 15 13 0 9 2
14 12 1 0 9 11 13 11 9 13 1 0 9 11 2
17 9 13 7 1 3 0 9 0 11 11 14 3 13 7 13 9 2
4 9 2 11 2
5 0 9 13 3 0
12 0 2 0 2 9 7 9 3 1 9 9 12
2 11 2
22 9 1 9 9 1 0 9 13 0 9 9 0 9 0 9 12 2 0 9 1 11 2
18 13 15 9 2 15 13 2 16 4 9 13 0 9 1 9 0 9 2
13 1 0 9 4 3 13 2 16 9 13 3 0 2
28 1 0 9 4 13 13 1 15 3 16 12 0 9 2 16 0 9 4 13 9 13 0 12 9 1 10 9 2
26 13 9 2 16 0 9 13 0 2 13 9 2 3 9 2 13 11 11 2 9 0 9 0 0 9 2
14 1 9 9 13 4 1 9 11 13 9 1 9 12 2
26 9 11 11 11 11 13 2 16 4 13 4 13 3 12 9 2 7 15 9 7 0 2 0 2 9 2
9 9 13 1 9 1 0 9 1 9
2 0 9
16 13 0 7 0 9 3 9 9 2 3 9 2 9 7 9 2
11 13 9 1 10 9 13 9 9 0 11 2
18 9 10 9 4 13 1 9 0 0 9 7 3 1 9 0 0 9 2
27 1 15 9 4 13 0 9 2 3 2 0 9 2 0 9 7 9 0 9 2 3 0 9 7 0 9 2
29 1 12 9 9 1 12 9 13 9 0 9 12 9 2 7 15 3 1 9 0 9 0 9 2 0 7 0 9 2
12 12 9 13 9 1 9 7 12 0 0 9 2
18 13 9 1 0 2 0 2 0 2 0 7 0 9 7 1 11 11 2
13 1 12 9 9 1 0 9 13 1 0 9 12 2
10 9 13 0 9 9 7 0 9 9 2
15 1 9 9 7 9 15 15 9 13 16 3 0 7 0 2
26 1 12 9 9 12 13 1 12 0 9 2 12 1 12 9 1 11 7 12 1 0 9 1 0 9 2
15 1 0 9 13 1 12 0 9 12 7 1 12 0 12 2
24 1 9 13 2 16 0 9 13 0 0 9 2 7 0 9 13 0 1 0 9 9 7 9 2
20 1 12 0 15 12 13 1 9 3 0 7 0 9 2 1 12 0 3 12 2
38 0 13 9 2 16 9 0 9 7 0 9 13 1 15 9 9 2 9 7 9 3 0 2 16 13 0 9 2 7 15 1 9 0 7 0 0 9 2
3 2 11 2
1 3
19 11 7 11 1 0 9 0 9 1 0 9 1 11 13 11 12 2 12 2
4 9 1 9 13
7 9 11 2 9 13 13 9
5 11 2 11 2 2
20 16 13 0 9 1 0 9 2 9 11 3 13 9 1 0 9 1 0 9 2
27 9 9 12 9 9 1 9 4 1 9 13 1 12 2 9 2 7 1 0 0 9 13 1 9 7 9 2
19 3 1 9 14 2 9 3 13 2 13 9 1 9 1 0 9 1 11 2
41 1 10 9 4 9 9 9 13 1 9 2 1 9 15 7 13 2 16 1 9 1 0 0 9 1 11 13 9 0 9 11 1 9 11 2 15 4 13 13 9 2
26 0 13 2 16 3 0 9 1 0 9 13 9 11 2 14 9 13 13 9 2 15 13 1 15 0 2
6 1 11 4 13 3 2
15 1 10 9 13 2 7 13 9 9 2 16 4 15 13 2
7 13 13 9 7 9 9 2
4 11 13 13 9
5 11 2 11 2 2
33 11 11 2 0 9 0 9 9 1 9 0 9 2 13 13 0 9 13 10 0 9 1 11 0 9 2 0 9 11 1 0 9 2
21 0 9 11 0 9 13 1 0 9 1 11 0 9 7 13 15 13 9 1 9 2
30 12 9 1 9 9 11 13 9 9 9 11 11 13 9 2 3 13 13 1 9 2 7 3 3 13 9 1 9 3 2
4 0 9 1 11
7 11 11 13 11 1 10 9
5 11 2 11 2 2
19 0 9 12 2 9 0 11 1 0 11 13 11 11 12 2 9 1 11 2
10 3 4 13 1 0 9 13 10 9 2
24 7 1 9 15 13 0 9 11 2 7 16 15 13 1 9 9 10 9 2 13 15 0 9 2
20 13 4 13 9 1 9 2 16 1 11 13 15 0 2 13 9 11 11 11 2
21 1 11 4 9 11 13 1 3 0 2 7 7 11 13 0 9 1 0 9 9 2
20 13 4 13 14 12 9 9 1 9 2 16 10 9 4 13 9 0 12 9 2
17 1 11 9 13 2 16 15 12 12 9 13 1 9 2 13 11 2
21 1 9 13 13 1 12 9 1 9 7 11 13 1 12 7 12 9 9 1 9 2
8 1 11 4 13 0 9 9 2
19 7 16 4 15 13 14 12 9 2 0 4 13 1 0 9 2 13 11 2
23 0 9 13 9 11 1 9 1 9 11 13 0 9 7 1 9 13 0 9 0 9 11 2
6 11 4 13 1 11 2
4 1 11 9 0
8 12 9 13 12 2 9 0 9
2 11 2
15 0 0 9 3 13 12 9 2 1 15 13 1 9 9 2
22 1 11 15 1 12 9 1 0 9 9 11 13 12 3 0 9 2 0 9 7 11 2
12 12 9 13 0 2 11 13 14 3 0 9 2
21 9 11 15 3 13 2 16 9 9 11 13 1 0 9 2 7 3 14 1 9 2
23 9 11 3 1 9 3 13 9 9 2 15 15 2 3 2 13 9 9 2 9 11 11 2
7 1 9 1 11 7 13 2
27 1 9 3 2 3 1 12 9 2 13 9 1 11 2 3 13 9 1 11 2 0 3 1 0 0 9 2
21 0 13 9 2 1 10 9 13 2 1 9 13 9 11 2 11 2 11 2 11 2
8 11 3 3 13 1 0 9 2
6 1 9 3 13 11 2
10 9 11 13 1 9 1 0 2 11 2
15 9 15 3 4 13 13 1 11 2 15 15 13 1 11 2
14 9 11 7 3 13 9 11 2 0 1 9 1 11 2
6 3 0 2 0 0 9
12 1 11 13 12 2 9 9 11 1 9 12 9
7 11 2 11 2 11 2 2
34 9 0 9 2 11 2 12 2 7 11 2 11 2 12 9 2 13 3 1 9 11 11 1 11 0 9 0 0 9 9 11 2 12 2
21 10 9 13 9 12 9 2 0 1 9 12 2 0 9 13 12 7 0 12 9 2
7 0 9 3 13 12 9 2
29 0 9 13 1 11 3 1 0 9 1 0 11 1 11 7 4 13 2 16 4 15 9 9 13 9 1 12 9 2
21 1 9 3 1 10 9 13 2 7 9 11 7 11 13 11 11 10 9 9 13 2
5 13 4 3 11 2
36 3 9 13 1 15 2 10 9 15 9 13 2 13 9 11 11 7 1 0 9 13 2 1 9 15 13 9 11 2 15 13 15 3 2 2 2
18 10 0 9 2 11 2 13 3 1 11 7 3 15 13 9 1 11 2
23 16 13 9 0 3 1 9 0 9 2 3 16 15 2 2 1 10 0 9 13 0 13 2
20 7 16 1 9 13 0 9 1 0 0 9 2 9 11 11 3 1 9 13 2
24 13 7 0 0 9 11 11 1 9 11 7 11 11 2 9 0 9 11 11 7 3 0 9 2
12 0 9 1 11 13 1 9 9 11 0 9 2
19 1 9 4 0 9 10 9 13 13 1 12 9 2 9 9 13 12 2 2
14 1 3 0 0 0 2 0 9 15 3 13 0 9 2
13 0 9 15 1 0 9 4 13 13 1 12 9 2
19 0 9 11 15 1 9 13 0 9 7 11 11 13 0 9 1 11 11 2
29 11 11 2 9 11 2 0 9 11 2 13 1 11 9 0 1 9 9 2 11 2 11 2 11 2 7 10 9 2
16 0 9 1 11 7 0 9 1 0 9 9 13 0 9 9 2
23 1 9 11 13 1 0 0 9 11 2 11 2 12 2 12 2 0 9 11 1 0 9 11
2 9 11
4 0 9 0 9
10 9 9 13 0 9 7 9 9 1 9
2 11 2
25 1 0 0 9 12 2 9 9 1 0 9 1 9 11 11 3 0 9 13 0 9 7 9 9 2
11 9 13 1 9 14 1 9 12 2 9 2
12 0 9 1 9 9 13 0 11 11 1 11 2
9 0 9 11 13 1 12 0 9 2
8 13 7 2 1 15 13 11 2
17 13 3 11 2 7 16 1 10 9 13 10 0 9 2 13 11 2
13 3 1 9 9 9 13 0 0 9 2 11 2 2
7 13 12 9 1 0 9 2
32 9 2 15 13 1 0 9 14 12 9 2 4 13 0 0 9 16 9 2 15 13 1 0 9 1 12 0 2 15 13 9 2
17 7 9 2 10 9 9 11 13 2 15 4 13 1 0 9 13 2
19 3 13 13 1 12 9 7 12 9 1 9 2 16 3 13 1 0 9 2
12 0 9 4 13 7 1 9 1 9 1 9 2
30 0 9 13 1 0 9 0 9 1 9 12 9 7 12 9 2 3 12 9 2 12 0 9 7 1 9 14 12 9 2
6 9 13 13 9 0 9
2 11 2
27 13 9 9 7 9 13 9 9 0 9 2 15 1 9 9 13 9 9 9 2 11 2 1 9 1 11 2
21 1 0 9 15 13 12 0 9 2 9 9 13 9 12 9 2 15 13 0 9 2
23 1 9 11 11 11 4 15 13 9 2 15 3 13 1 11 2 3 13 1 0 0 9 2
9 1 0 7 0 9 13 3 9 2
26 9 1 0 9 7 13 11 3 1 0 0 9 2 0 9 7 1 9 7 9 9 3 1 0 9 2
14 9 2 15 4 13 1 12 9 2 4 13 1 9 2
8 0 9 4 1 10 9 13 2
10 1 9 9 0 9 13 4 9 13 2
13 3 3 13 11 2 11 2 13 0 9 12 9 2
7 0 4 13 1 0 9 2
16 9 15 13 1 9 0 9 7 9 2 0 9 7 0 9 2
15 15 13 1 11 0 9 2 15 13 0 3 1 0 9 2
28 1 0 9 13 2 16 0 9 9 1 3 12 0 13 0 1 9 7 9 9 7 9 2 3 3 1 9 2
17 0 9 15 13 2 16 1 0 9 9 15 4 10 9 9 13 2
5 9 1 9 13 0
7 0 9 11 11 1 0 9
5 11 11 2 11 11
10 13 15 15 2 3 4 13 1 11 2
7 13 15 3 0 3 13 2
23 9 4 3 13 13 2 3 4 13 3 2 7 3 4 9 13 2 16 15 13 3 0 2
38 0 9 11 11 2 15 13 1 11 1 0 9 2 13 7 0 9 0 15 11 2 16 4 13 13 2 16 13 1 11 3 2 13 4 15 3 0 2
5 11 13 16 11 2
21 7 3 13 0 13 3 2 16 4 1 15 13 3 15 3 1 10 9 7 9 2
5 4 3 13 11 2
10 15 13 0 2 11 13 3 1 9 2
15 13 1 15 7 9 2 13 9 7 13 2 7 15 13 2
4 13 1 9 2
9 13 15 0 9 9 1 0 9 2
11 13 2 16 4 13 9 2 9 1 9 2
24 3 4 13 9 1 9 1 9 2 7 9 2 15 13 9 1 9 2 16 4 15 13 9 2
37 16 4 15 15 3 13 13 9 1 9 1 9 7 1 9 2 7 15 9 1 9 13 2 13 4 9 1 0 9 14 1 9 2 7 1 9 2
19 16 4 13 1 9 2 13 4 15 2 16 13 1 9 7 4 13 9 2
5 13 13 9 11 2
6 11 13 1 0 9 2
18 3 15 13 7 3 13 1 9 2 16 4 13 12 7 3 7 0 2
8 11 13 0 9 2 1 0 2
11 9 3 13 13 3 1 9 0 0 9 2
8 11 15 13 13 0 9 9 2
11 15 13 0 9 2 3 3 13 9 13 2
10 0 9 1 11 11 13 0 9 0 12
3 13 9 9
7 11 2 9 11 11 2 2
10 9 9 0 9 13 13 0 1 11 2
22 1 9 0 9 3 13 9 0 0 9 2 15 13 14 9 9 2 7 7 0 9 2
30 9 9 13 13 9 0 9 2 13 15 9 2 9 9 13 4 13 2 7 3 7 9 9 0 9 15 9 4 13 2
26 1 9 9 9 13 13 0 9 1 9 1 9 13 2 16 9 9 13 9 3 1 9 7 9 15 2
30 16 0 9 13 9 0 9 1 9 12 9 15 13 2 15 1 9 13 0 0 9 1 9 15 13 1 11 12 9 2
17 1 9 9 7 10 0 9 13 9 1 0 9 3 4 15 13 2
21 9 9 13 4 13 1 0 9 2 9 1 9 0 9 0 9 1 0 9 9 2
8 0 9 13 9 1 9 11 11
7 11 2 11 2 11 2 2
43 0 9 1 11 3 1 0 9 13 1 0 9 9 0 9 1 11 2 1 15 4 0 0 9 11 11 13 1 9 0 9 1 0 0 9 0 11 1 12 9 9 9 2
9 0 9 13 9 0 9 1 9 2
7 13 15 9 9 11 11 2
17 0 9 15 9 13 1 0 9 1 9 0 0 9 1 9 12 2
28 15 15 13 1 15 2 16 1 0 9 12 2 9 13 7 13 9 9 9 1 9 9 0 11 1 9 9 2
13 15 15 1 0 9 13 9 1 0 9 0 9 2
28 9 2 15 0 9 1 11 1 9 9 13 2 11 13 1 15 2 16 1 9 9 15 3 13 13 0 9 2
3 9 13 9
7 9 1 9 0 9 13 0
5 11 2 11 2 2
38 9 2 15 9 9 9 11 11 13 9 9 0 11 11 11 2 2 16 13 9 0 9 1 9 9 1 9 0 11 2 13 0 9 13 9 9 9 2
42 1 0 9 0 0 9 11 13 9 2 16 0 1 9 0 9 9 2 15 13 9 1 9 9 0 15 1 0 9 2 15 13 16 9 11 2 15 9 0 11 13 2
14 10 9 4 0 9 3 13 1 9 7 9 1 11 2
8 9 15 9 13 16 0 9 2
33 1 10 9 0 9 9 9 10 9 15 13 1 0 9 0 9 1 9 9 2 15 13 1 9 9 1 0 2 9 2 7 3 2
32 0 13 7 9 9 2 16 9 9 13 7 1 9 9 1 9 9 7 16 13 0 9 13 9 2 15 9 9 13 1 9 2
26 3 2 16 13 1 9 9 2 1 15 13 0 9 1 0 9 7 9 7 0 9 2 9 9 13 2
18 0 9 2 15 1 0 9 13 2 13 1 9 11 3 3 1 9 2
38 9 0 15 0 9 15 13 2 16 10 9 1 0 9 1 0 9 13 13 1 10 9 2 7 7 1 15 2 16 13 0 9 0 9 1 0 9 2
7 4 13 9 0 9 1 0
5 11 2 11 2 2
34 9 0 9 2 15 13 1 0 9 2 7 3 1 0 9 1 9 13 1 11 3 3 1 9 3 2 1 0 11 3 0 0 9 2
18 9 13 9 1 12 9 2 13 3 0 9 7 10 9 13 3 0 2
30 11 11 2 9 9 0 9 1 9 9 7 0 9 2 11 2 15 7 13 2 16 10 9 15 4 7 1 15 13 2
20 16 0 9 13 3 13 0 9 0 9 2 0 9 4 13 13 3 0 9 2
25 11 2 11 13 1 9 9 16 0 9 2 16 9 13 3 3 3 9 1 0 9 3 1 9 2
30 1 9 1 9 13 15 2 15 15 13 9 2 1 11 13 13 0 9 14 12 9 2 16 1 9 13 3 1 9 2
13 3 1 9 1 9 7 9 13 9 9 0 9 2
31 9 1 0 2 15 13 3 0 9 16 1 9 2 13 13 9 3 15 0 9 9 9 7 0 2 15 15 13 0 9 2
30 0 4 13 2 16 4 15 9 9 12 9 13 1 0 12 9 1 12 9 3 2 3 13 15 0 1 0 0 9 2
18 9 1 15 2 16 4 10 9 1 9 12 3 13 2 4 3 13 2
22 9 9 13 2 13 15 0 9 9 0 0 9 2 3 16 15 13 9 9 15 9 2
46 1 0 9 1 9 9 0 9 11 2 15 9 13 3 1 9 2 15 13 2 16 9 9 0 9 13 13 9 9 1 3 0 9 2 16 13 9 2 9 2 9 2 9 7 9 2
23 9 9 13 13 0 9 1 0 9 1 9 7 13 9 9 2 13 15 7 13 1 9 2
8 3 0 9 13 0 16 9 2
16 1 9 1 0 9 13 9 1 9 14 3 0 16 1 9 2
2 13 3
2 0 9
2 11 11
16 13 3 2 13 1 9 9 2 13 9 7 13 1 12 9 2
12 13 3 2 1 10 9 13 1 12 9 3 2
25 13 3 3 7 3 3 2 13 9 2 16 4 13 13 1 2 1 9 0 2 0 12 9 9 2
25 13 3 2 13 1 0 9 0 9 7 0 9 0 9 15 13 1 12 9 0 16 9 1 9 2
14 1 9 1 9 9 15 9 13 1 12 9 1 12 2
27 13 3 2 13 15 13 7 9 1 9 2 7 15 13 2 16 1 0 9 13 13 1 9 9 0 12 2
33 7 16 4 13 9 2 13 1 15 9 2 7 1 16 4 15 13 2 3 15 13 2 16 1 9 7 1 9 13 1 9 9 2
22 11 2 3 13 2 13 9 2 9 13 1 9 7 13 15 13 1 0 9 1 9 2
17 9 15 7 13 3 0 9 7 13 15 13 2 3 13 1 9 2
31 13 15 7 14 15 2 1 9 3 15 13 2 3 15 13 1 0 9 10 9 2 16 9 0 9 13 3 1 0 9 2
20 10 9 13 3 15 2 7 16 10 9 4 1 10 9 3 13 2 13 9 2
34 3 1 10 9 1 15 13 13 9 7 9 2 7 14 3 2 16 13 9 0 2 13 15 1 15 3 1 9 2 15 3 13 9 2
2 3 2
11 16 3 15 1 15 2 3 15 1 15 2
20 3 15 2 16 15 2 9 7 9 2 15 13 1 15 9 7 9 3 13 2
12 15 15 15 13 7 1 10 9 4 15 13 2
11 1 9 15 13 2 7 3 3 13 13 2
30 13 15 3 2 16 13 13 15 9 2 16 4 15 1 15 13 9 2 7 13 0 9 2 16 4 15 13 3 9 2
22 10 9 2 1 15 13 2 3 3 2 7 3 13 0 2 16 1 15 15 13 9 2
29 7 15 13 2 16 9 15 4 7 3 1 9 13 9 14 3 2 16 1 15 13 7 16 9 13 1 12 9 2
18 1 10 9 15 13 2 16 4 13 2 16 4 13 3 1 0 9 2
8 13 15 13 13 16 13 9 2
8 13 13 13 16 13 1 9 2
14 7 0 9 15 1 15 15 13 2 3 15 15 13 2
5 13 15 10 9 2
18 7 13 15 13 2 14 2 15 14 2 13 15 2 0 9 1 9 2
6 13 15 16 0 9 2
11 3 4 13 1 9 9 1 12 9 3 2
13 13 15 1 9 2 3 3 13 7 9 13 13 2
20 9 15 13 1 9 2 14 2 9 2 3 2 9 2 3 15 13 2 9 2
5 9 9 7 9 2
17 9 0 9 2 7 9 2 15 15 0 13 3 7 3 13 9 2
14 1 9 0 9 13 15 2 15 15 13 1 0 9 2
21 0 9 7 0 9 2 3 14 13 2 15 13 2 7 0 13 2 15 4 13 2
4 15 2 11 2
6 3 15 1 15 13 2
4 7 13 9 2
13 9 15 13 9 1 9 2 16 4 15 13 9 2
33 13 15 9 2 16 4 15 1 15 13 9 2 1 15 15 3 13 10 9 2 15 15 13 3 14 3 2 16 15 3 13 0 2
4 9 9 9 13
5 11 2 11 2 2
25 3 12 5 1 0 12 5 4 13 1 0 9 13 1 0 9 1 9 9 1 0 9 0 9 2
9 0 12 5 13 13 9 0 9 2
21 11 15 3 13 0 9 9 9 11 11 1 15 2 16 15 3 13 1 0 9 2
19 1 10 9 13 3 9 1 9 1 0 9 1 9 12 3 1 12 5 2
15 3 0 9 13 1 11 2 11 12 1 0 9 0 9 2
41 9 3 13 2 16 4 9 1 9 1 0 9 2 15 13 0 9 2 4 13 1 9 7 0 9 1 9 12 2 12 1 9 9 2 1 0 9 12 2 12 2
10 1 0 9 13 9 9 9 10 9 2
4 11 13 0 9
5 11 2 11 2 2
17 0 9 1 12 9 9 13 1 0 9 0 0 9 2 11 2 2
12 11 15 3 13 9 9 0 9 9 11 11 2
13 1 0 9 0 9 4 9 13 4 13 1 9 2
18 16 11 11 13 2 4 9 1 0 9 1 0 2 0 9 3 13 2
29 0 9 13 1 0 9 0 9 7 0 9 2 9 13 3 0 9 2 0 7 0 9 7 0 0 7 0 9 2
12 1 0 0 9 0 9 13 0 11 7 11 2
8 0 9 12 9 13 12 9 2
21 1 9 11 11 15 9 13 1 0 9 2 0 0 9 13 12 12 5 12 9 2
22 16 11 11 13 2 13 0 0 9 3 3 1 9 0 9 2 3 1 12 9 9 2
12 0 9 12 9 13 1 10 9 9 0 9 2
1 3
9 9 0 0 9 4 13 1 11 2
9 3 13 1 11 9 0 0 9 2
12 1 9 1 11 15 1 15 13 9 12 9 2
38 2 11 2 0 9 0 9 2 15 13 9 9 1 9 9 2 9 7 9 1 0 12 9 2 15 1 9 13 1 12 9 2 1 12 9 1 9 2
9 1 9 13 10 9 3 12 9 2
7 9 13 1 9 12 9 2
5 0 9 1 9 13
11 0 9 13 0 9 0 2 0 9 13 11
2 11 2
18 0 9 0 9 3 13 12 9 9 1 12 9 2 9 1 9 12 2
7 1 12 9 7 3 13 2
17 9 1 0 9 15 13 1 12 9 9 2 3 9 9 9 12 2
21 13 15 1 0 9 1 0 9 2 15 13 9 11 1 9 7 9 2 11 2 2
22 0 9 0 0 9 13 11 2 15 15 0 9 12 9 9 13 1 0 9 1 11 2
12 1 9 12 13 11 14 12 9 9 0 9 2
22 1 11 13 7 9 9 9 1 0 9 3 13 1 12 7 12 9 11 7 0 11 2
18 0 9 1 15 13 0 12 9 9 7 10 9 1 0 9 15 13 2
22 13 15 7 9 2 1 15 4 9 0 11 13 9 2 15 4 3 13 1 0 9 2
20 9 9 1 0 11 3 13 14 12 9 9 2 15 13 1 9 9 1 11 2
24 0 9 9 1 10 9 3 13 12 9 9 7 13 14 1 9 0 16 0 0 9 1 11 2
16 1 0 9 3 3 13 0 9 9 9 11 1 12 9 9 2
17 11 13 3 0 9 0 0 9 2 16 3 13 0 12 9 9 2
18 1 11 13 3 0 9 9 0 11 2 15 13 3 0 0 0 9 2
16 3 2 14 1 12 9 2 9 2 15 13 9 9 1 11 2
7 13 15 12 9 9 12 2
9 0 9 1 9 1 9 3 1 9
5 11 2 11 2 2
15 9 9 1 9 4 13 4 9 3 13 3 14 1 9 2
13 13 15 11 11 2 9 9 9 0 9 9 9 2
16 9 0 9 9 13 0 9 2 9 7 0 9 2 1 9 2
8 10 9 13 0 0 9 9 2
16 9 11 13 2 16 9 13 13 0 9 2 15 1 9 13 2
17 9 15 3 13 2 16 1 9 13 13 9 9 9 9 1 9 2
13 13 15 2 16 15 13 13 1 9 2 13 11 2
25 1 9 9 13 7 0 2 16 4 10 9 4 3 13 1 9 3 1 9 9 1 9 0 9 2
11 13 15 0 2 16 15 15 13 0 9 2
22 1 11 1 15 2 16 4 15 0 9 4 3 13 1 9 2 13 7 9 9 9 2
12 4 13 1 9 13 10 0 9 2 13 11 2
3 11 13 9
5 11 2 11 2 2
12 0 9 13 1 9 0 9 15 1 0 9 2
15 9 9 0 9 15 1 9 11 11 13 3 9 0 9 2
8 13 3 1 9 1 10 9 2
16 1 10 9 13 1 15 7 0 9 1 9 16 3 1 11 2
28 3 2 9 9 11 15 1 15 13 3 3 16 0 9 2 15 1 0 9 1 9 0 9 7 9 13 9 2
16 9 9 7 0 9 7 9 15 1 15 9 13 1 9 3 2
22 1 9 11 11 2 11 13 2 16 9 3 4 13 1 0 0 9 9 0 0 9 2
17 15 13 4 1 0 9 13 9 1 9 1 9 9 9 2 13 2
19 9 9 1 9 11 13 3 13 2 16 11 13 0 9 1 9 0 9 2
6 11 1 9 14 1 9
5 11 2 11 2 2
19 0 9 11 1 9 11 2 11 15 4 13 0 0 9 13 14 9 9 2
17 9 0 9 11 11 3 13 2 16 15 11 13 1 9 13 3 2
19 13 2 16 0 9 4 3 13 3 3 7 9 9 13 13 3 9 9 2
27 1 9 9 11 13 11 2 11 13 2 16 9 9 9 9 0 9 4 1 0 9 13 1 12 2 9 2
21 9 9 1 0 2 0 9 13 3 1 0 11 13 14 1 9 12 9 0 9 2
7 3 13 1 0 0 9 2
14 1 0 9 13 3 1 9 3 14 12 11 7 11 2
14 9 11 13 11 2 11 13 3 3 1 9 12 9 2
6 0 9 13 9 13 2
31 0 9 9 11 15 13 13 13 9 0 9 7 0 0 0 2 9 4 13 1 9 1 9 9 1 11 1 9 9 12 2
8 9 9 13 3 9 16 9 2
17 16 15 9 3 13 2 1 9 1 0 9 9 3 13 13 9 2
8 9 15 13 3 1 0 9 2
3 9 11 11
3 9 1 9
2 11 2
11 1 9 9 1 12 0 9 13 0 9 2
9 13 15 3 9 9 11 11 11 2
15 0 9 1 10 9 15 1 0 9 13 1 12 9 9 2
11 1 0 9 4 15 13 3 12 9 9 2
21 12 1 0 9 1 11 13 9 2 16 13 3 2 9 1 9 9 1 9 9 2
11 3 13 9 1 9 3 12 9 2 9 2
13 9 13 3 0 9 0 9 7 0 9 1 9 2
1 3
21 9 0 7 0 9 11 2 11 13 3 1 0 9 1 12 9 1 12 9 9 2
20 9 15 1 10 0 9 13 1 0 2 16 9 0 0 9 13 3 3 0 2
22 9 0 9 1 0 9 0 7 0 11 13 1 0 9 1 12 9 1 12 9 9 2
19 9 1 10 9 1 11 7 1 0 9 13 1 12 9 1 12 9 9 2
3 9 1 9
14 0 0 9 9 1 9 13 0 9 1 9 0 11 2
9 1 11 7 11 13 1 9 11 2
15 11 11 0 2 4 13 7 9 9 1 11 7 1 11 2
29 1 9 12 2 2 12 2 9 15 1 11 13 12 2 0 9 9 1 0 2 0 1 9 0 9 1 0 9 2
14 9 16 9 1 0 7 0 9 13 3 3 0 9 2
34 0 9 9 11 2 15 15 13 1 0 0 9 2 13 1 9 0 1 9 9 0 9 11 0 13 1 0 0 9 1 15 0 9 2
27 9 13 13 1 15 0 9 1 9 2 9 2 9 2 9 2 7 7 1 0 9 16 9 2 9 3 2
22 0 9 9 11 13 1 9 0 9 11 0 11 1 9 12 5 12 9 0 0 9 2
18 9 13 0 9 2 3 10 9 1 11 13 3 12 12 9 1 9 2
16 0 9 1 0 9 11 11 12 1 9 11 13 10 0 9 2
16 1 15 2 16 13 0 1 11 2 13 9 9 1 0 9 2
11 1 0 7 9 13 9 0 0 9 9 2
14 12 2 9 13 9 11 12 1 10 1 0 0 9 2
19 1 9 1 0 0 9 4 13 0 9 10 0 9 2 9 11 7 11 2
4 2 2 11 2
7 11 3 3 13 0 9 9
8 0 11 2 11 2 11 2 2
26 0 9 9 13 1 0 9 9 7 9 2 13 3 11 9 0 9 9 9 1 0 9 11 2 11 2
14 9 11 11 1 15 13 9 1 0 9 1 12 9 2
10 3 3 0 0 9 7 13 0 9 2
38 11 2 11 2 9 0 2 9 2 11 11 2 15 13 12 9 0 9 1 11 2 10 9 13 7 13 2 13 1 0 9 16 0 9 0 0 9 2
19 9 13 3 16 9 1 9 1 9 9 7 0 9 2 15 13 10 9 2
7 13 3 2 7 1 9 2
16 9 15 15 13 13 2 16 15 4 9 13 7 1 10 9 2
10 1 0 9 9 9 9 13 0 13 2
11 1 11 2 11 13 1 11 3 10 9 2
28 13 15 1 15 2 16 4 13 0 3 13 9 1 15 2 0 9 4 13 9 0 9 7 3 4 13 13 2
10 0 9 15 7 3 1 15 13 13 2
17 9 13 0 0 9 2 15 13 9 9 14 3 1 0 9 9 2
17 15 15 3 13 1 9 0 9 1 9 0 0 9 7 0 9 2
15 0 9 2 13 15 2 1 10 9 13 7 9 7 9 2
4 9 1 9 11
2 11 2
16 9 1 0 0 9 11 13 0 9 11 11 9 9 11 11 2
21 11 3 2 13 2 16 1 11 13 3 0 0 9 2 1 15 13 0 13 9 2
29 11 13 3 12 9 9 0 9 2 16 3 0 9 12 9 1 9 0 9 13 1 9 9 0 9 1 10 9 2
14 0 9 13 2 16 4 4 13 7 13 9 9 11 2
28 3 13 13 9 9 1 9 11 1 0 9 0 9 2 7 3 9 9 9 11 2 15 13 11 3 1 9 2
14 11 3 13 2 16 1 10 9 13 1 0 9 11 2
26 9 9 9 4 13 4 13 11 7 9 9 11 2 16 0 9 15 1 9 1 0 9 13 0 9 2
4 0 9 0 9
9 0 9 11 13 1 0 9 0 9
3 0 11 2
21 3 12 9 9 4 13 13 0 9 0 9 11 2 0 1 9 0 7 0 9 2
26 16 13 1 9 9 9 11 11 2 12 1 9 9 2 13 15 0 9 9 1 12 5 10 0 9 2
15 9 13 1 9 3 12 9 9 2 15 13 1 12 9 2
11 11 13 12 9 1 0 9 14 12 9 2
23 3 12 5 9 9 13 1 9 2 1 9 15 13 10 9 13 14 1 12 7 12 5 2
10 1 9 13 9 12 9 1 0 9 2
14 3 12 5 9 13 9 2 0 9 9 7 3 9 2
24 0 9 11 13 7 9 7 0 9 9 2 1 15 13 11 9 1 0 9 2 0 2 9 2
19 1 9 13 0 9 9 0 9 2 15 13 12 2 12 9 10 0 9 2
20 0 0 9 13 3 9 0 0 9 7 11 2 3 15 13 0 9 1 9 2
17 11 13 1 9 3 12 7 12 9 9 9 1 9 1 9 9 2
12 9 9 13 1 11 2 11 3 16 12 9 2
29 9 0 9 13 9 1 10 0 9 9 3 12 9 9 0 0 9 2 15 3 13 1 9 7 3 16 0 9 2
18 9 11 13 1 9 12 1 9 1 9 1 9 11 0 9 11 11 2
14 13 15 3 3 9 1 9 2 9 2 9 7 9 2
6 9 3 13 0 9 2
5 11 1 9 1 9
3 0 9 2
18 0 9 12 9 9 13 1 12 2 9 0 9 0 9 11 0 9 2
8 13 15 0 9 9 11 11 2
40 0 2 9 2 11 0 9 2 3 0 2 9 2 0 9 7 9 2 15 13 9 0 0 9 2 9 7 9 0 9 2 0 9 9 7 9 1 0 9 2
9 0 9 3 13 10 0 9 9 2
11 9 1 15 13 7 11 2 13 11 11 2
14 13 2 16 0 9 1 0 9 15 0 13 7 13 2
12 0 9 9 13 1 0 9 3 12 9 9 2
10 3 12 15 1 0 9 9 13 9 2
14 0 9 13 1 11 9 0 0 9 1 0 0 9 2
20 11 2 10 0 9 13 12 9 2 9 2 4 13 1 0 9 3 0 9 2
10 11 13 12 9 9 2 9 12 9 2
4 0 9 9 11
2 11 2
22 0 9 9 11 0 2 2 0 0 9 9 7 0 9 13 1 0 9 1 12 5 2
14 0 9 13 3 1 0 9 1 9 7 0 0 9 2
21 9 13 1 10 9 9 12 9 9 2 16 1 0 9 0 9 14 12 9 9 2
18 9 13 1 12 9 1 12 9 9 1 12 9 9 1 0 9 3 2
10 11 3 13 9 3 9 10 0 9 2
19 15 13 13 12 9 9 2 15 13 1 12 9 3 2 16 13 0 9 2
13 13 2 1 9 12 9 2 9 13 0 9 9 2
17 1 0 9 13 0 9 11 12 9 9 2 9 9 12 9 9 2
20 9 11 13 2 16 9 15 13 9 3 0 9 1 10 9 1 0 9 12 2
11 1 0 9 13 9 9 1 9 12 9 2
13 11 13 2 16 1 0 9 13 1 0 12 9 2
11 0 9 4 3 13 0 2 16 15 13 2
18 0 9 0 9 2 3 0 7 0 9 2 13 13 3 0 9 9 2
5 9 13 13 11 11
4 11 1 11 2
26 9 0 9 3 13 9 1 9 3 0 9 0 0 9 1 0 9 1 0 9 9 11 11 1 11 2
19 13 3 9 2 15 15 3 13 9 12 0 9 1 0 9 2 11 2 2
17 13 15 3 9 11 11 2 9 2 9 2 0 2 2 11 11 2
15 11 13 0 9 7 0 0 9 15 3 13 2 13 9 2
19 1 9 0 9 7 9 0 9 4 9 9 7 9 11 13 3 1 9 2
16 9 11 2 1 15 4 9 13 2 13 1 9 0 9 9 2
21 1 10 0 9 7 0 9 1 11 2 11 13 13 0 9 1 0 9 0 9 2
13 9 0 9 4 1 3 0 9 13 1 9 12 2
17 1 9 2 3 13 1 9 0 9 2 0 9 10 9 3 13 2
14 10 9 0 9 1 9 11 13 7 13 9 1 9 2
7 1 9 13 13 12 12 9
2 11 2
18 1 12 12 9 4 1 9 13 9 1 9 9 1 9 1 0 9 2
10 13 1 15 9 9 7 0 0 9 2
9 3 13 0 13 3 12 9 9 2
15 14 2 11 2 13 0 9 1 9 1 9 1 0 9 2
2 9 11
9 11 15 15 0 9 13 3 3 2
16 9 11 12 11 2 9 13 3 1 11 2 7 13 3 3 2
10 1 9 13 3 13 7 9 7 9 2
11 1 9 13 7 0 9 7 0 0 9 2
11 13 13 2 16 15 9 1 11 3 13 2
2 2 11
4 0 9 13 11
2 11 2
27 0 9 9 0 0 9 3 1 9 0 9 1 9 1 9 0 1 9 7 11 1 9 13 11 7 11 2
8 13 15 1 11 0 9 9 2
21 13 3 2 16 0 9 0 3 1 11 15 13 3 1 0 9 7 1 0 9 2
39 9 9 12 0 9 1 9 1 9 1 9 1 0 9 11 13 9 1 9 0 9 2 0 9 1 11 7 11 2 7 13 11 2 16 4 10 9 13 2
3 11 13 9
2 11 2
21 0 0 9 2 11 2 3 13 2 16 13 10 0 9 1 9 0 11 1 11 2
11 0 7 15 0 9 13 1 9 1 9 2
13 0 9 11 11 13 2 16 13 10 9 3 13 2
26 0 9 13 9 11 13 9 1 0 9 7 0 9 1 9 9 7 9 9 1 9 9 1 0 11 2
16 14 10 9 1 9 9 7 13 9 1 9 9 11 0 9 2
16 0 9 1 9 11 13 0 9 7 0 9 13 1 0 11 2
10 3 1 9 12 2 0 15 3 13 9
4 9 13 0 9
5 11 2 11 2 2
18 1 0 12 1 12 5 4 15 1 0 9 13 13 9 1 0 9 2
12 3 9 1 9 1 0 9 4 13 4 13 2
14 13 15 1 9 9 9 1 9 2 15 3 13 9 2
22 16 13 9 9 11 11 2 9 10 9 13 0 9 0 9 7 9 9 15 9 11 2
18 15 13 0 9 9 1 12 7 12 9 7 0 1 12 7 12 9 2
17 9 4 15 14 13 3 13 1 0 9 2 3 3 1 0 9 2
19 1 9 0 9 15 9 13 13 0 9 1 9 9 9 9 13 10 9 2
15 9 9 1 0 9 13 3 9 1 12 9 13 0 9 2
21 1 11 15 13 1 9 9 2 7 1 9 0 0 9 13 9 0 0 9 13 2
21 9 13 3 13 0 9 2 13 4 13 4 9 0 1 0 9 7 0 0 9 2
9 3 1 9 12 2 9 4 9 13
11 11 11 13 9 9 2 13 9 9 0 9
7 11 2 11 2 11 2 2
30 9 0 2 9 2 11 2 15 13 1 0 9 0 7 0 9 2 11 2 2 13 1 9 9 9 0 9 11 11 2
5 11 13 9 11 2
23 1 9 11 13 9 11 13 2 16 1 9 9 13 13 1 0 9 0 9 11 11 11 2
47 1 10 9 13 9 9 1 9 0 0 9 9 11 11 1 11 2 11 2 1 15 15 15 9 11 13 2 16 3 10 0 9 11 2 11 13 9 9 7 13 1 9 9 11 2 11 2
31 1 12 1 9 9 11 9 11 2 11 1 9 11 2 11 3 13 1 0 9 9 1 9 9 11 1 9 9 1 11 2
26 1 9 15 1 9 11 11 11 2 15 11 13 2 13 9 2 1 15 4 11 2 11 13 1 9 2
31 1 9 11 15 9 11 1 9 2 16 10 9 13 1 9 2 13 0 9 2 9 1 11 2 3 9 0 9 9 9 2
13 11 10 9 3 13 7 13 1 0 9 10 9 2
22 0 0 9 9 9 11 11 11 13 2 16 1 10 9 15 3 0 9 13 0 9 2
13 9 9 13 0 0 9 2 10 0 9 13 11 2
10 1 10 9 13 12 0 0 9 9 2
33 1 10 9 11 2 11 1 9 13 9 9 11 2 1 15 15 13 2 16 11 2 11 3 13 9 2 15 13 13 1 10 9 2
22 9 15 3 9 13 2 16 10 9 13 1 0 7 16 11 2 11 3 13 13 9 2
16 11 11 3 11 9 2 16 4 15 13 13 9 11 2 13 2
10 13 15 9 2 15 15 13 9 11 2
25 3 4 15 1 9 1 10 3 0 13 9 11 2 16 13 9 2 16 1 9 13 1 9 9 2
20 16 15 10 9 13 2 4 15 13 1 0 9 10 9 2 13 11 2 11 2
11 1 11 13 13 9 10 9 0 9 9 2
13 1 9 2 3 9 13 2 9 13 2 13 11 2
3 9 16 9
2 11 11
8 0 11 13 2 15 3 13 2
11 1 9 13 0 9 0 9 11 7 11 2
17 1 0 9 2 0 9 0 9 7 11 2 10 9 13 12 9 2
29 7 13 0 9 13 1 9 11 11 7 10 0 9 7 13 0 9 13 3 2 16 4 3 13 9 0 0 9 2
18 0 9 2 13 0 11 2 15 3 13 12 9 9 2 1 10 9 2
28 16 1 15 10 13 2 15 13 13 2 13 15 2 13 9 0 9 1 11 11 11 2 9 0 7 0 9 2
27 0 9 13 15 2 16 0 9 1 0 9 1 9 13 9 11 1 11 7 13 9 0 9 1 0 9 2
41 16 15 7 9 2 1 11 13 1 10 9 13 2 13 13 2 16 9 1 9 9 4 13 3 2 4 0 11 3 13 2 16 15 9 1 9 13 1 10 9 2
9 1 15 13 0 9 9 1 9 2
11 1 0 9 2 13 0 0 9 3 3 2
12 15 13 1 9 13 2 16 15 15 15 13 2
21 0 13 3 15 2 16 9 13 0 11 13 7 9 3 0 9 10 9 3 13 2
33 16 0 9 13 13 9 2 4 3 13 9 2 15 4 15 15 13 13 2 14 15 15 13 13 2 13 3 12 1 0 0 9 2
35 0 11 15 10 9 2 1 10 9 11 13 13 2 13 13 9 1 9 2 16 0 9 7 11 3 13 9 2 15 1 9 1 11 13 2
7 10 9 13 7 11 11 2
21 11 13 9 13 0 9 7 13 15 9 0 9 2 15 13 9 0 2 0 11 2
12 13 1 15 13 7 1 10 0 9 1 11 2
14 1 9 0 9 9 11 13 2 13 0 9 11 0 2
8 15 3 13 9 9 9 13 2
7 9 1 0 11 13 13 2
18 13 4 7 13 1 11 11 2 7 16 10 9 1 11 13 3 3 2
7 9 1 9 9 2 12 13
14 1 11 11 13 14 9 2 16 15 9 9 13 1 9
5 11 2 11 2 2
49 0 9 9 2 12 2 15 13 1 11 11 2 9 13 1 0 9 2 1 15 13 11 7 11 3 13 2 16 3 13 1 0 9 2 9 0 9 2 9 9 12 0 9 2 7 9 0 9 2
30 9 2 15 15 1 9 2 12 13 2 13 1 0 9 2 7 7 9 9 9 1 9 9 1 9 1 9 2 12 2
39 1 9 9 13 3 1 9 1 0 9 3 1 9 7 9 13 9 9 9 11 2 11 9 9 0 11 0 2 11 2 2 15 1 11 13 0 9 11 2
14 11 15 1 11 13 7 12 0 9 11 7 0 11 2
25 9 11 11 2 11 15 13 9 1 11 2 15 15 14 1 9 9 1 9 13 13 1 0 9 2
20 1 9 2 15 11 13 2 13 2 16 11 13 0 9 1 9 1 0 11 2
11 10 9 13 0 9 2 3 11 3 13 2
20 9 9 11 2 15 15 13 13 7 0 9 9 1 11 2 1 11 13 0 2
32 1 9 11 2 1 10 9 13 7 0 7 0 9 2 13 9 2 16 10 9 2 3 15 13 1 9 0 9 2 13 11 2
18 11 7 13 9 3 1 9 9 2 12 2 15 9 11 1 11 13 2
37 1 11 13 15 2 16 10 9 13 0 1 11 2 0 13 7 1 0 9 11 2 1 0 9 13 9 12 1 0 7 0 0 9 7 1 9 2
15 1 11 13 14 9 2 16 15 9 2 12 13 1 9 2
34 1 0 9 15 7 13 13 9 2 16 1 11 4 9 13 16 1 0 9 7 14 1 0 9 2 1 15 15 13 9 9 7 9 2
9 1 9 1 0 9 2 9 13 9
5 1 0 9 1 11
10 9 0 9 13 11 7 13 1 9 2
20 13 1 0 0 9 10 9 2 1 15 13 13 12 9 1 9 7 1 9 2
19 9 2 15 4 13 10 9 3 2 4 1 0 9 13 1 0 9 9 2
9 1 9 1 9 15 13 0 9 2
17 9 13 2 16 0 9 7 9 0 9 15 9 1 10 9 13 2
58 1 15 2 15 13 12 0 9 1 9 2 16 15 13 9 9 7 13 9 9 1 9 2 10 9 13 1 0 9 9 9 9 11 2 15 13 1 9 1 0 9 2 15 13 11 3 1 12 2 7 13 15 15 7 0 0 9 2
3 2 11 2
4 10 9 13 9
5 11 2 11 2 2
19 9 2 16 1 9 3 13 10 9 2 13 13 13 9 9 1 0 9 2
14 1 0 0 9 15 13 9 12 1 15 2 11 11 2
21 1 0 9 13 1 0 9 12 7 12 0 9 2 15 15 13 3 9 0 9 2
24 9 3 13 9 2 9 7 9 13 3 3 0 9 9 16 3 2 3 7 13 7 1 9 2
11 3 3 13 0 9 0 9 1 0 9 2
16 9 9 11 7 13 2 16 4 13 13 1 9 3 1 9 2
16 9 13 9 1 0 9 2 3 15 2 15 15 13 1 9 2
12 13 3 3 14 0 9 2 15 15 9 13 2
21 16 11 13 9 0 0 9 2 9 15 13 3 9 7 3 15 9 13 1 15 2
17 0 9 9 15 3 4 13 3 1 9 2 15 13 0 0 9 2
5 0 9 1 0 9
2 11 11
34 0 9 9 0 9 1 0 9 2 15 4 9 9 13 1 0 9 1 11 2 13 0 9 0 7 3 9 3 0 9 10 9 9 2
17 3 13 7 9 10 9 1 9 2 9 2 15 9 13 3 3 2
38 0 11 13 0 9 13 15 1 9 9 0 0 9 2 1 0 9 9 2 1 9 0 9 7 0 9 7 1 0 9 7 1 0 9 9 11 11 2
27 1 0 0 9 13 1 0 9 1 9 9 0 9 2 1 9 9 10 9 13 1 11 7 3 1 11 2
30 3 13 3 1 0 9 1 9 9 1 11 1 11 2 3 15 3 13 1 9 1 11 7 0 9 0 0 0 9 2
24 1 9 15 11 13 1 11 2 3 1 15 13 9 7 0 0 9 2 0 9 10 0 9 2
17 13 7 0 9 0 9 11 2 3 13 1 9 3 0 0 9 2
25 9 0 9 2 15 9 2 11 13 2 15 3 13 2 16 3 13 0 9 0 9 2 0 11 2
14 0 0 9 9 2 11 7 10 9 13 0 9 11 2
30 13 1 15 1 9 12 2 1 0 9 4 7 11 13 2 1 1 9 1 9 9 7 1 0 9 2 14 9 12 2
9 11 13 3 0 3 1 10 9 2
20 0 9 11 15 10 9 13 3 1 0 9 2 0 9 12 2 9 9 12 2
5 15 14 13 3 2
35 4 13 1 9 0 0 9 9 12 2 3 1 9 2 3 1 9 13 3 3 0 9 12 2 9 2 0 2 7 1 9 13 9 0 2
27 1 10 9 13 10 0 9 1 0 9 9 14 12 9 2 15 15 1 0 9 13 13 14 1 9 12 2
21 9 11 9 12 13 1 11 2 13 0 9 7 0 9 2 10 10 9 15 13 2
6 15 15 9 3 13 2
40 0 0 9 0 0 9 13 9 0 9 11 12 0 3 1 11 11 2 10 9 0 9 10 9 1 9 7 12 1 3 10 0 0 0 9 1 9 0 9 2
47 1 1 0 9 9 9 13 0 13 3 14 1 0 9 2 7 7 13 16 13 1 9 9 1 11 2 11 12 2 11 12 2 7 3 7 1 9 2 11 2 11 2 11 2 11 2 2
27 1 0 9 0 3 13 9 3 0 9 11 12 2 0 1 9 9 11 2 11 1 9 12 1 11 11 2
12 13 9 11 2 11 7 0 9 1 0 9 2
11 1 0 9 9 13 14 13 0 9 9 2
20 1 15 13 7 0 0 9 0 0 9 2 3 3 0 9 9 2 11 11 2
18 0 10 0 9 13 9 9 11 2 12 2 0 1 9 12 11 11 2
41 15 13 12 1 12 9 9 0 9 2 0 13 1 11 1 11 2 11 12 2 12 1 9 11 9 11 2 2 0 1 11 2 11 1 9 9 11 2 11 2 2
36 1 9 13 2 16 15 13 3 15 9 0 9 2 15 15 13 7 13 13 2 1 9 0 9 1 0 9 14 1 9 9 0 7 0 9 2
11 1 10 9 0 7 0 9 0 9 13 2
21 1 9 9 0 7 0 9 4 13 7 0 9 11 7 11 2 0 9 9 11 2
56 11 0 13 1 0 9 14 9 0 9 2 3 0 1 9 9 10 9 2 7 16 12 1 10 3 3 3 13 2 3 0 9 13 9 7 3 0 4 13 13 1 15 2 7 3 9 3 0 9 1 9 0 7 0 9 2
32 1 9 2 15 15 13 0 9 2 13 7 13 0 9 11 2 12 2 0 9 11 2 12 2 9 1 9 0 11 2 2 2
27 1 9 9 2 15 1 3 0 9 3 10 9 3 13 9 2 3 7 13 13 1 9 0 9 0 9 2
22 9 12 9 0 7 0 0 9 1 9 13 7 3 13 9 10 9 1 0 9 9 2
31 1 0 9 2 1 9 9 9 7 9 2 3 0 9 9 13 13 2 16 13 15 2 15 3 13 9 9 11 7 0 2
14 16 15 1 10 9 13 2 4 15 13 1 15 13 2
18 9 0 9 11 11 13 3 1 9 1 0 9 1 11 0 0 9 2
19 16 9 13 9 11 11 2 15 1 9 12 13 9 1 9 0 11 11 2
5 9 11 11 2 11
12 9 0 9 4 1 9 13 13 7 9 1 9
5 11 2 11 2 2
36 1 9 0 9 1 9 1 9 0 9 9 13 2 16 0 0 9 1 0 9 13 1 0 9 0 9 3 2 1 9 1 12 9 12 9 2
27 0 9 1 9 2 9 2 9 2 0 9 2 9 2 9 2 3 0 9 13 1 0 9 9 12 9 2
7 3 15 3 13 12 9 2
32 9 0 9 1 0 0 9 9 13 3 1 0 9 13 1 12 9 2 9 0 9 0 1 0 9 0 9 13 12 9 2 2
33 9 1 0 9 9 7 0 9 2 15 9 13 2 7 13 2 16 4 1 9 0 9 4 9 1 0 9 9 13 9 1 9 2
11 15 4 13 0 9 1 0 9 7 9 2
23 10 9 13 3 1 0 9 0 9 0 9 7 10 9 1 9 9 15 4 3 3 13 2
34 9 13 15 2 16 15 9 2 15 4 15 13 1 0 9 1 0 9 2 4 13 9 1 0 9 2 15 4 13 0 9 1 9 2
20 3 13 3 12 12 9 11 1 0 9 2 0 12 1 0 7 0 1 0 2
26 1 0 7 0 9 13 1 12 5 0 9 2 14 12 5 0 7 3 1 12 5 0 7 0 9 2
27 13 15 2 16 4 9 1 0 9 13 1 0 9 2 13 3 0 2 16 10 9 1 9 13 1 9 2
4 13 11 9 2
5 11 2 11 2 2
13 9 9 9 11 13 1 0 9 0 9 1 11 2
27 10 9 13 3 9 9 0 9 2 15 4 13 9 12 9 7 0 9 1 10 9 13 12 9 2 9 2
37 9 10 9 1 9 0 13 9 7 0 12 9 2 9 11 11 2 0 0 9 9 11 11 2 15 0 9 13 2 7 0 0 9 1 0 9 2
16 9 0 9 13 13 0 9 2 9 2 9 2 9 7 9 2
17 16 15 9 13 9 2 13 11 9 13 15 1 0 1 0 9 2
3 11 1 11
5 11 2 11 2 2
29 12 9 9 4 13 0 9 2 15 13 13 9 7 0 9 1 0 9 1 11 11 2 0 9 9 0 1 9 2
18 11 13 1 10 9 12 12 9 0 9 2 0 9 13 9 1 9 2
27 0 9 13 15 0 1 9 0 11 2 10 9 4 9 13 13 1 0 9 0 9 2 3 1 0 9 2
11 7 3 4 9 1 0 9 13 0 9 2
8 1 0 9 13 1 11 9 9
5 11 2 11 2 2
27 1 9 0 9 1 0 9 2 15 4 1 9 9 1 9 9 13 1 9 2 4 3 3 13 0 9 2
27 9 13 9 1 0 9 1 9 2 3 3 13 9 1 0 9 2 13 1 15 0 9 9 11 11 11 2
23 0 9 7 13 10 9 7 3 4 13 1 15 2 16 9 13 3 1 0 9 1 9 2
41 3 2 16 15 1 9 13 7 0 9 2 0 9 3 13 13 9 1 9 2 15 4 16 9 0 0 9 13 1 11 1 12 9 7 3 13 1 3 0 9 2
29 7 16 4 9 13 13 2 13 13 2 16 10 9 0 9 13 1 10 9 1 9 3 0 2 13 11 2 11 2
7 1 9 15 4 13 1 9
5 11 2 11 2 2
29 1 9 1 11 3 13 0 0 9 2 9 1 0 9 2 1 15 15 3 10 9 13 2 4 15 7 13 13 2
21 9 3 1 9 7 9 9 1 11 3 13 13 2 16 0 9 13 0 9 9 2
12 13 1 12 9 2 3 9 7 9 1 9 2
30 10 9 9 1 11 13 15 2 16 1 12 2 9 13 9 15 9 3 1 12 9 7 13 2 16 3 13 0 9 2
29 1 9 0 9 2 3 13 9 1 10 9 13 9 2 13 9 0 9 11 11 2 9 15 4 1 15 13 13 2
12 13 9 9 9 1 0 9 2 16 4 13 2
20 9 2 9 7 9 2 15 13 9 12 9 2 15 1 9 4 13 1 9 2
9 9 15 15 4 13 13 1 9 2
16 10 9 15 13 3 2 16 1 0 9 15 13 9 9 9 2
19 9 4 13 0 7 9 9 2 15 15 1 9 13 13 2 13 11 11 2
15 1 11 15 14 3 13 13 9 2 7 4 13 3 0 9
5 11 2 11 2 2
16 1 0 9 4 15 13 13 1 11 13 9 3 1 9 12 2
21 13 15 1 9 9 11 11 2 15 7 3 13 2 16 13 1 9 1 0 9 2
10 10 9 3 0 0 0 9 3 13 2
21 3 15 1 11 13 3 14 14 12 9 7 1 0 9 15 13 3 1 0 9 2
21 9 15 13 1 0 9 13 2 7 0 9 1 0 9 13 0 9 7 1 15 2
19 4 2 14 9 13 9 2 1 15 9 13 2 4 9 0 9 13 15 2
21 13 14 9 2 13 15 9 7 13 15 2 3 1 0 0 9 2 0 0 9 2
18 9 2 15 3 13 2 4 13 3 3 0 9 2 16 13 3 9 2
20 1 0 9 15 7 13 1 15 2 16 3 0 9 9 4 13 9 1 9 2
13 9 1 0 7 0 9 4 3 13 1 9 9 2
27 16 3 15 13 9 2 15 7 3 3 13 15 0 2 3 4 13 9 13 3 1 9 2 3 1 9 2
26 1 10 0 9 3 13 12 9 1 12 9 7 3 15 13 0 13 1 9 2 16 13 15 0 9 2
27 11 11 7 13 2 16 9 0 0 9 13 1 9 9 1 12 9 2 15 4 13 4 1 0 9 13 2
6 9 1 0 9 1 9
7 11 2 11 2 11 2 2
31 1 9 9 4 15 13 0 9 13 1 15 2 10 0 0 9 4 13 1 0 9 1 10 9 7 15 4 15 13 13 2
21 13 1 15 3 0 0 9 1 0 9 2 0 9 9 11 2 11 2 11 2 2
49 0 9 13 9 9 2 1 15 13 13 10 9 3 1 9 12 9 1 11 7 1 11 2 1 9 9 11 2 11 7 11 2 7 16 15 13 1 0 9 1 0 2 0 2 0 7 0 11 2
11 9 4 15 3 13 13 1 9 0 9 2
29 9 11 11 2 11 2 13 2 16 9 13 13 1 10 9 2 15 13 1 9 0 9 2 7 2 3 12 9 2
25 9 9 13 2 16 0 9 0 9 2 1 15 9 1 0 0 9 13 9 12 9 2 9 13 2
1 9
31 9 13 9 1 9 1 9 2 9 1 9 2 7 1 9 9 13 2 10 9 3 7 3 13 9 9 0 1 9 13 2
47 0 9 2 16 13 3 2 13 13 1 9 0 9 7 0 9 15 13 1 15 2 3 0 9 13 7 3 3 13 0 0 9 13 3 2 16 4 9 9 7 9 9 13 0 2 0 2
13 9 12 5 12 9 13 3 12 9 1 0 9 2
18 0 9 13 0 3 1 12 9 2 1 10 9 15 3 13 9 11 2
21 1 9 0 9 15 1 10 9 13 0 9 2 7 3 9 0 9 15 9 13 2
19 1 0 9 15 13 0 0 9 7 13 15 0 9 2 15 13 0 9 2
16 9 13 3 0 9 9 9 1 9 1 9 0 9 2 9 2
12 0 9 13 9 9 3 1 9 9 0 9 2
10 3 9 9 9 13 13 10 0 9 2
14 9 9 0 9 13 3 12 5 0 16 1 0 9 2
11 9 7 0 0 9 13 0 9 1 9 2
10 9 13 9 2 3 1 9 13 9 2
25 13 0 2 16 9 10 9 13 4 13 1 9 0 9 9 2 9 2 9 2 9 2 9 2 2
18 0 9 7 0 9 13 1 9 0 9 13 2 7 3 13 1 9 2
42 0 9 11 2 9 2 9 3 13 13 7 9 11 13 3 1 0 9 2 15 13 12 2 12 5 0 9 9 2 9 3 13 12 9 2 9 2 13 15 9 2 2
21 10 0 9 13 9 1 9 7 1 15 15 13 9 0 3 1 15 3 0 9 2
14 15 13 13 7 9 0 2 0 3 2 1 9 11 2
14 15 3 13 9 9 9 7 10 0 9 3 13 3 2
4 2 2 11 2
5 9 11 13 1 9
10 11 11 1 9 1 9 0 9 1 11
2 11 11
28 9 9 13 9 9 11 1 0 9 1 9 0 9 2 0 0 0 11 2 9 1 9 0 9 1 0 9 2
6 9 0 0 11 13 2
7 13 3 1 9 7 9 2
9 9 11 13 3 1 9 10 9 2
21 1 9 0 9 3 13 1 9 9 1 9 0 9 2 11 2 1 11 11 11 2
23 3 15 13 13 2 16 1 3 0 0 9 4 13 9 2 15 1 9 0 9 3 13 2
7 9 9 11 4 3 13 2
18 1 9 2 3 2 16 4 15 13 2 16 13 10 0 9 1 9 2
24 9 2 15 4 13 12 2 7 12 2 9 12 1 11 2 7 13 1 9 12 7 9 12 2
7 1 10 9 3 11 13 2
18 1 9 2 1 9 9 2 4 3 3 0 9 9 0 0 9 13 2
6 3 9 9 13 3 2
8 1 9 11 4 15 7 13 2
11 13 15 10 9 2 3 1 9 10 9 2
13 10 9 0 9 2 15 13 1 9 13 2 13 2
23 9 10 9 13 1 0 9 11 7 11 2 3 9 13 2 7 13 9 1 0 0 9 2
14 9 11 15 13 10 9 2 15 13 1 9 0 9 2
10 10 9 4 1 0 9 1 9 13 2
13 1 0 9 9 15 13 3 12 0 7 0 9 2
8 1 0 9 15 13 14 11 2
4 11 1 9 11
2 11 2
18 9 11 11 2 0 9 0 9 1 9 0 9 2 13 9 9 11 2
33 10 9 1 9 13 2 16 11 15 13 1 11 7 11 13 9 7 16 10 9 13 4 1 9 12 13 1 9 9 1 0 9 2
10 11 13 1 3 0 9 2 13 11 2
11 13 2 16 10 9 13 1 9 11 9 2
20 9 1 9 9 15 11 13 1 9 1 0 9 3 13 7 13 1 0 11 2
19 3 13 11 11 13 1 0 9 0 9 1 11 12 2 3 13 0 9 2
10 9 15 13 2 16 11 13 9 0 9
8 11 2 11 2 11 2 11 2
14 9 1 9 11 13 9 0 9 3 13 0 9 11 2
52 9 0 9 2 16 4 9 9 0 9 13 0 9 1 3 0 0 9 7 9 9 13 1 0 9 9 11 1 0 9 2 13 0 9 1 9 11 1 0 9 1 9 2 3 15 15 0 9 13 0 9 2
23 9 11 11 2 9 0 2 13 2 16 4 9 11 9 9 9 13 3 1 10 0 9 2
38 11 13 2 16 9 9 11 13 3 0 9 7 3 0 13 7 9 11 2 16 3 1 9 9 7 1 9 13 9 2 15 4 3 13 9 9 9 2
25 13 2 16 4 13 0 2 16 4 15 15 13 7 13 1 0 9 7 16 4 15 13 0 9 2
25 9 11 3 13 1 9 10 0 9 2 16 4 9 9 3 1 0 9 11 13 13 9 0 9 2
23 13 2 16 13 9 2 15 13 1 3 0 9 2 9 0 9 7 9 7 0 0 9 2
7 11 11 13 1 9 9 9
5 11 2 11 2 2
15 0 9 9 7 10 9 1 9 13 9 0 9 0 9 2
18 16 15 9 9 3 13 2 13 1 9 11 11 11 12 7 12 9 2
24 1 10 9 13 14 0 9 9 9 2 15 15 1 0 13 14 1 12 9 1 9 2 13 2
22 11 3 1 9 11 11 1 0 0 9 11 13 2 16 9 9 13 14 1 12 9 2
15 9 13 1 10 9 15 1 9 2 7 0 9 13 0 2
19 10 0 9 13 14 12 9 1 9 0 9 2 16 4 13 3 15 13 2
10 0 9 13 3 9 2 13 9 9 2
15 11 13 2 16 13 7 0 9 2 15 13 7 12 9 2
22 1 10 9 13 1 10 9 9 0 2 1 9 7 9 2 13 1 15 11 2 11 2
10 0 9 10 9 13 2 14 15 13 2
15 11 13 9 9 2 16 15 3 13 13 10 9 9 9 2
32 16 4 13 3 2 0 9 9 9 2 15 4 13 0 1 9 13 2 9 4 13 2 15 3 13 2 7 13 4 9 3 2
10 3 13 15 1 11 1 9 0 11 2
9 9 0 9 4 11 1 9 13 2
11 11 2 13 4 13 4 7 0 9 1 9
5 11 2 11 2 2
32 1 0 9 1 0 7 0 1 0 9 4 15 13 13 9 9 2 15 13 4 13 0 0 9 1 9 1 9 0 0 9 2
15 13 15 3 9 0 9 9 1 9 2 11 2 11 11 2
18 9 4 1 10 9 13 1 9 2 16 4 1 0 9 9 9 13 2
25 1 9 9 2 15 13 4 13 9 1 9 2 15 9 13 1 0 0 9 7 15 9 7 9 2
29 1 0 0 9 9 13 12 9 2 9 7 9 2 10 9 4 13 7 1 0 9 13 2 3 3 12 12 9 2
29 1 9 11 2 3 4 9 13 10 3 0 9 1 0 9 2 11 13 2 16 15 1 9 9 3 13 7 13 2
10 3 9 13 7 13 0 9 0 9 2
16 1 11 13 9 3 13 9 2 7 0 9 13 13 7 11 2
17 9 9 14 9 3 13 1 15 2 16 4 10 9 1 11 13 2
7 1 0 9 11 1 11 13
5 11 2 11 2 2
27 1 0 9 11 0 1 0 9 4 3 3 13 2 16 4 4 13 1 9 1 9 0 1 0 0 9 2
14 3 4 13 1 9 2 15 13 0 9 1 0 9 2
21 9 15 3 1 11 13 0 9 9 11 11 2 15 3 13 0 0 9 0 9 2
29 0 9 13 2 16 9 10 9 2 15 15 0 11 13 2 13 13 9 0 2 7 3 9 2 15 1 9 13 2
16 0 9 13 0 7 13 13 7 15 1 9 13 2 13 11 2
7 0 9 9 13 3 0 2
18 1 15 1 10 9 13 0 9 1 10 0 9 1 11 1 0 9 2
17 1 0 9 1 9 9 0 9 11 11 4 13 2 13 0 9 2
21 11 11 3 13 1 9 11 11 2 1 9 11 11 2 1 9 0 9 11 11 2
23 1 9 3 0 9 11 11 11 7 0 9 3 13 3 13 7 1 0 9 9 12 9 2
34 1 9 0 9 13 3 15 13 2 13 0 9 11 11 1 15 2 16 0 9 13 3 2 9 13 15 1 0 9 3 1 0 9 2
14 9 11 11 15 13 2 16 10 9 13 3 3 13 2
7 0 9 1 9 1 0 9
5 11 2 11 2 2
22 1 0 9 0 9 11 1 9 0 0 9 13 3 10 9 0 9 2 0 9 0 2
18 10 9 0 3 7 3 2 1 0 0 9 9 2 13 3 0 9 2
24 9 1 15 13 3 1 9 2 16 10 9 13 1 0 9 16 1 9 2 3 10 9 13 2
14 0 9 1 10 9 13 9 2 15 13 9 3 3 2
12 1 9 9 9 13 7 0 9 3 7 3 2
22 9 11 2 11 11 11 13 2 16 4 10 0 9 13 13 7 9 0 9 1 11 2
17 13 4 15 3 1 10 9 1 0 9 2 16 4 15 13 9 2
24 13 2 16 4 13 9 3 13 7 13 16 9 9 9 2 7 3 13 0 0 9 1 9 2
16 13 4 0 0 9 1 9 2 16 13 10 9 0 0 9 2
17 13 1 9 9 3 7 3 2 7 16 13 3 1 9 0 9 2
24 0 9 13 3 0 2 16 13 13 0 7 0 9 2 3 3 9 1 0 9 0 9 13 2
20 10 9 0 9 2 15 1 10 9 3 13 9 9 2 11 2 11 13 13 2
17 10 0 9 1 9 9 13 2 10 9 13 3 1 0 9 9 2
14 11 13 2 16 0 9 4 13 9 0 7 0 9 2
22 11 2 11 4 13 2 16 4 15 1 10 9 1 9 0 9 13 7 0 0 9 2
12 9 1 11 11 2 11 2 2 9 0 9 9
25 13 0 9 9 1 0 9 3 1 0 9 1 9 12 2 7 13 0 9 2 16 3 13 3 2
18 3 13 13 0 9 11 1 11 2 16 1 0 9 9 7 13 13 2
23 10 0 9 7 3 15 13 2 0 13 13 15 3 2 16 4 1 15 13 4 3 13 2
13 13 9 7 3 12 9 13 13 1 15 0 9 2
21 1 9 2 3 13 9 2 15 3 13 16 13 2 16 15 15 1 10 9 13 2
38 7 13 2 16 13 0 13 1 9 1 11 14 1 9 2 3 4 13 9 15 13 2 16 9 13 9 2 3 13 2 13 2 14 15 1 9 12 2
24 16 13 2 0 9 9 13 0 9 10 0 9 7 1 9 15 0 9 13 9 11 1 11 2
27 16 16 9 1 9 12 13 3 2 1 0 9 13 13 2 16 1 10 0 9 1 0 9 15 15 13 2
6 13 3 0 3 13 2
3 2 11 2
8 1 11 1 11 7 0 0 9
16 3 14 15 13 2 10 15 1 10 9 13 0 0 9 11 2
26 10 9 15 13 10 9 2 10 9 7 1 9 9 13 1 12 0 9 2 7 15 13 9 10 9 2
23 15 2 15 15 13 9 1 9 9 1 11 2 1 15 13 13 15 2 15 0 14 14 2
30 1 9 0 9 7 9 3 0 9 15 13 10 9 13 1 9 0 9 7 3 15 13 1 0 9 11 7 10 9 2
16 10 9 7 13 10 7 3 10 9 7 9 9 3 3 13 2
18 11 1 9 2 9 0 9 11 2 13 0 2 15 3 3 13 9 2
20 1 12 9 2 1 9 2 13 3 0 9 7 3 9 1 9 11 1 11 2
29 13 15 14 3 13 2 13 11 2 13 1 9 15 2 15 15 13 13 2 7 1 9 15 15 9 13 1 9 2
8 3 15 13 7 1 0 9 2
26 1 11 13 9 1 9 7 13 7 13 7 9 9 13 7 9 7 9 1 11 2 9 7 11 11 2
23 9 13 13 1 3 16 12 9 0 9 11 2 11 12 7 11 12 7 11 2 9 2 2
27 11 1 9 13 9 2 15 3 13 10 0 9 2 7 10 9 2 9 9 1 11 7 11 2 13 3 2
20 1 12 9 9 13 15 3 0 2 7 1 0 9 0 9 1 9 10 9 2
3 2 11 2
7 11 14 13 1 9 1 9
3 1 0 9
5 11 2 11 2 2
43 0 9 9 2 11 2 13 0 9 1 0 9 1 9 0 11 7 11 2 11 2 2 15 15 1 11 13 2 7 1 0 0 9 2 11 2 2 15 13 1 10 9 2
10 11 15 3 13 9 11 11 2 11 2
28 13 3 9 9 0 9 11 11 2 11 2 16 14 9 0 9 1 10 9 13 2 3 3 1 11 7 11 2
23 1 9 13 0 13 2 10 9 1 9 0 15 1 11 13 2 16 3 13 9 0 9 2
18 3 13 14 12 9 2 15 13 0 9 11 7 13 9 2 13 11 2
4 9 9 13 9
2 0 9
6 11 11 2 11 2 2
39 0 11 11 1 11 11 2 15 4 1 0 0 9 1 0 9 13 0 9 1 9 0 9 9 9 2 9 7 9 2 3 9 9 2 11 11 13 9 2
41 10 0 9 15 13 11 2 11 13 1 9 12 15 2 16 13 9 2 1 15 15 13 2 16 4 9 13 0 9 2 7 10 9 13 0 3 16 9 7 9 2
24 0 9 0 9 13 9 2 16 15 9 13 9 1 10 0 9 2 15 13 13 1 10 9 2
27 9 2 11 1 9 9 13 2 16 9 9 1 0 9 2 15 4 13 16 0 9 2 1 10 9 13 2
20 1 1 15 2 16 1 0 9 13 3 12 9 2 13 9 13 7 16 9 2
12 12 9 13 9 13 3 1 9 0 2 0 2
31 13 0 2 16 15 9 13 10 9 2 16 13 9 11 2 15 9 13 14 1 9 12 9 7 1 0 9 13 13 9 2
26 3 16 0 9 15 13 9 1 0 9 2 13 1 9 9 9 0 9 9 0 9 9 2 11 11 2
4 0 9 1 9
5 11 2 11 2 2
26 1 0 9 0 9 7 9 0 7 0 9 7 9 4 1 0 9 13 0 11 2 11 2 1 11 2
11 0 0 9 13 9 1 9 0 0 9 2
18 1 9 13 13 9 1 9 9 2 9 0 1 9 9 7 0 9 2
16 9 2 15 9 3 13 2 13 4 1 9 13 1 0 9 2
6 1 0 9 12 9 9
2 0 9
5 11 2 11 2 2
28 1 0 9 1 11 15 13 0 9 1 9 0 11 11 2 2 15 3 1 9 13 1 0 11 9 12 9 2
14 9 13 1 9 0 2 7 15 15 1 0 9 13 2
36 1 9 11 11 2 0 9 3 13 1 9 10 3 0 9 2 13 15 1 9 10 9 2 15 13 9 2 7 0 9 13 7 3 0 9 2
33 0 2 15 9 4 13 1 9 1 9 1 0 9 2 1 9 13 2 16 9 13 3 7 13 13 3 9 2 15 15 13 9 2
7 3 14 3 14 13 9 2
19 13 2 16 15 1 9 13 15 3 2 7 16 13 2 16 15 15 13 2
44 12 1 9 2 15 11 2 11 2 3 3 3 13 0 9 2 13 2 16 15 0 10 9 13 7 1 0 9 7 3 1 15 13 13 2 3 0 4 15 13 1 0 9 2
18 13 15 14 16 0 9 2 15 9 13 3 1 9 2 7 1 9 2
34 9 13 1 9 2 16 15 13 1 9 0 7 3 0 2 16 1 0 9 13 2 16 11 2 11 2 13 9 9 3 0 16 9 2
14 16 13 9 2 13 9 2 16 10 9 13 13 9 2
39 15 0 11 11 2 2 15 4 13 1 9 2 7 1 9 13 0 9 2 4 13 0 1 0 9 9 1 9 7 13 1 12 9 3 1 9 1 9 2
1 9
30 9 13 9 9 2 1 15 9 9 9 2 12 13 12 2 12 2 1 12 9 2 1 0 9 2 1 11 12 9 2
13 9 13 13 1 9 12 7 0 2 9 2 12 2
7 0 9 7 9 1 0 9
2 11 11
16 3 0 9 9 1 9 0 0 9 13 1 9 12 11 9 2
14 1 9 12 13 10 9 10 9 1 11 7 0 11 2
11 1 0 9 7 13 3 10 9 0 9 2
12 13 3 1 3 3 0 0 9 1 10 9 2
27 15 1 15 13 13 15 2 16 0 9 1 9 12 13 9 9 9 12 2 0 1 9 1 0 0 9 2
14 9 13 7 1 12 9 1 9 1 0 7 0 9 2
5 14 13 0 9 2
14 9 9 13 2 13 15 7 9 2 15 9 13 3 2
12 1 0 9 15 0 2 0 2 0 9 13 2
10 13 15 15 9 2 9 1 9 3 2
4 14 11 9 2
15 15 13 1 9 10 0 9 9 1 9 10 12 0 9 2
4 9 9 13 2
33 14 0 9 2 7 9 0 0 9 2 15 1 0 9 9 7 1 15 3 9 11 7 0 11 11 2 13 1 9 0 0 9 2
19 9 7 13 9 9 2 1 15 15 3 13 2 7 1 10 9 15 13 2
13 0 9 13 9 2 9 1 9 15 13 13 13 2
17 9 3 3 0 9 13 2 16 9 15 3 13 1 9 0 9 2
3 13 9 2
35 15 7 13 9 13 9 0 9 1 0 9 7 3 3 13 9 1 9 9 1 9 2 10 9 13 1 9 2 7 1 10 9 13 0 2
9 3 13 9 9 9 13 9 9 2
8 7 15 1 15 2 0 9 2
3 9 1 9
1 9
2 11 11
15 3 3 13 1 9 1 11 0 9 1 0 0 11 11 2
9 1 10 9 13 1 9 3 3 2
9 1 9 2 11 13 9 0 11 2
17 1 9 10 9 11 11 7 3 1 10 9 9 13 0 0 9 2
25 3 15 1 9 2 15 13 0 9 0 9 2 13 2 16 15 1 0 9 4 13 0 9 9 2
25 9 3 1 9 0 0 9 2 3 15 1 9 0 9 13 9 0 1 9 0 9 2 9 13 2
11 13 15 7 9 1 0 0 9 1 11 2
4 11 15 13 2
15 13 13 9 1 9 7 13 9 1 0 9 7 0 9 2
15 3 2 13 15 14 9 9 2 16 9 3 15 3 13 2
15 3 9 13 1 9 0 9 9 2 1 9 1 0 9 2
7 9 1 10 9 15 13 2
35 3 0 9 0 9 13 3 1 9 9 2 1 15 2 16 15 9 3 13 0 0 9 2 0 15 13 13 9 7 10 9 9 1 9 2
8 13 0 13 2 15 13 0 2
12 13 9 0 9 0 9 4 7 13 3 0 2
7 0 9 15 13 1 0 9
1 9
5 11 11 2 11 11
20 0 9 13 13 13 9 1 9 0 2 0 9 1 12 0 0 9 3 3 2
27 9 0 7 0 0 9 7 0 9 15 3 3 13 13 2 16 3 7 1 3 3 15 4 0 9 13 2
31 3 13 9 2 15 9 11 13 1 9 3 1 9 1 10 0 0 9 11 2 7 13 0 13 2 16 13 15 9 0 2
43 1 9 2 3 1 9 0 9 1 15 0 1 0 9 2 13 0 9 7 9 9 0 0 9 1 9 3 2 3 13 2 2 13 0 9 9 3 0 9 13 1 9 2
23 3 13 15 1 0 7 0 9 1 9 9 9 7 0 9 2 3 1 9 16 0 0 2
32 0 9 9 15 1 11 13 3 3 2 13 2 16 9 9 13 13 0 2 16 0 9 13 4 1 9 13 7 1 0 9 2
11 13 3 9 2 1 15 15 3 3 13 2
22 9 12 9 15 3 13 9 2 1 15 15 13 3 13 2 7 13 3 10 9 13 2
40 11 11 13 7 3 14 0 16 11 11 2 3 3 15 2 3 3 4 0 9 13 1 10 9 2 13 1 9 9 13 1 15 2 3 15 9 0 9 13 2
19 9 0 7 15 9 13 7 0 7 0 9 15 1 15 9 11 3 13 2
9 9 9 4 3 13 9 0 9 2
12 9 0 9 3 7 10 9 1 11 13 4 2
26 0 0 9 10 9 2 15 3 13 13 2 3 13 9 1 9 3 1 11 2 13 7 3 1 15 2
2 3 2
5 0 9 2 0 9
7 1 9 0 9 2 12 2
2 11 11
7 9 15 3 13 1 9 2
24 1 0 9 2 3 1 9 12 2 15 16 0 9 13 9 2 15 4 1 0 9 13 9 2
39 0 9 0 9 7 9 2 0 2 3 0 0 9 2 4 1 9 9 3 13 9 11 2 7 15 1 0 9 11 2 12 2 0 1 9 1 9 12 2
13 11 11 2 12 13 0 9 7 15 9 0 9 2
38 1 12 2 9 13 7 10 0 9 3 0 9 2 15 13 1 10 9 7 0 9 2 7 3 10 0 9 1 0 9 1 9 2 9 2 9 3 2
16 1 10 9 15 13 13 9 9 2 3 3 0 1 0 9 2
13 9 1 9 15 13 12 2 7 0 9 1 9 2
10 7 15 13 9 3 0 9 16 3 2
23 3 9 3 13 2 7 1 0 9 9 15 9 1 0 9 3 3 13 0 3 3 13 2
24 9 13 11 2 1 0 0 9 13 9 11 2 11 2 1 15 3 11 2 11 7 0 11 2
17 11 13 1 9 12 9 11 2 12 2 1 9 12 3 9 12 2
8 3 13 1 9 0 9 12 2
13 0 9 7 0 0 9 9 13 9 9 1 15 2
7 10 0 9 13 0 9 2
15 9 9 13 9 9 2 9 2 1 15 15 13 0 9 2
12 1 9 13 9 14 9 0 1 0 9 9 2
30 1 9 13 3 10 9 9 2 9 1 0 9 9 9 2 9 2 9 9 2 9 9 2 0 7 0 9 2 2 2
34 0 9 9 2 15 1 15 13 13 10 0 9 2 3 9 9 2 0 9 3 2 2 13 3 1 9 9 2 7 15 3 0 9 2
8 0 9 9 9 3 3 13 2
12 13 15 2 16 4 3 13 1 0 9 0 2
5 15 13 10 9 2
12 0 9 0 9 3 13 7 3 3 13 4 2
21 16 1 12 2 7 12 2 9 13 9 1 0 9 2 3 13 10 9 3 0 2
14 1 15 4 3 13 1 9 9 2 15 13 0 9 2
30 1 10 9 9 7 9 10 9 13 0 9 2 3 2 9 2 2 7 0 9 9 1 15 2 3 10 0 0 9 2
9 1 10 0 9 15 3 7 13 2
35 1 9 1 9 15 9 13 9 1 12 9 2 0 9 2 15 4 13 3 0 7 3 0 2 16 4 15 13 13 0 9 7 3 9 2
22 0 9 13 9 12 2 9 9 11 7 11 2 11 2 15 13 0 9 0 2 9 2
8 1 10 9 3 13 0 9 2
28 10 9 7 3 13 13 3 0 2 9 4 3 13 10 0 0 9 7 10 9 13 3 9 9 0 0 9 2
6 1 0 9 0 9 2
21 0 9 9 13 14 15 2 16 13 1 0 9 0 9 2 3 9 0 1 9 2
15 13 3 1 9 1 11 2 15 13 7 13 9 0 9 2
19 1 15 1 9 13 9 1 9 0 9 2 7 1 0 7 3 0 9 2
22 1 12 2 7 12 2 9 1 15 13 3 10 0 9 0 1 9 9 11 7 11 2
26 13 1 0 9 2 10 9 0 9 2 7 3 7 0 9 2 4 13 1 9 11 1 0 0 9 2
34 3 13 1 9 9 11 12 2 3 12 7 12 2 9 11 2 9 2 7 9 11 12 2 3 7 0 9 2 9 11 2 9 2 2
5 14 1 9 9 13
1 9
2 11 11
52 0 9 2 7 3 3 1 9 0 0 9 2 15 1 15 3 13 1 15 2 16 13 0 0 7 0 9 2 16 9 13 3 9 2 7 3 9 7 13 2 14 9 3 13 9 2 7 13 3 0 9 2
10 15 15 13 2 13 15 15 2 0 2
26 3 0 13 2 16 4 9 9 2 9 9 2 16 7 9 15 15 2 4 13 3 3 7 3 3 2
13 0 9 13 10 9 2 15 13 9 9 1 9 2
8 0 13 2 9 2 9 9 2
9 0 13 2 13 15 7 15 13 2
7 13 15 7 15 15 13 2
8 13 15 15 13 7 15 13 2
18 9 2 15 15 13 9 9 2 13 3 1 9 2 10 15 15 13 2
53 13 15 14 12 9 1 10 2 15 13 2 12 9 1 10 2 15 13 2 12 9 1 9 2 1 15 13 2 12 9 1 10 2 15 3 13 7 13 2 7 12 9 1 9 7 9 2 15 15 13 13 0 2
7 9 0 9 13 3 0 2
22 15 13 2 16 3 13 9 2 15 13 1 10 9 0 2 7 16 1 15 4 13 2
26 7 3 2 16 13 9 2 16 4 15 1 10 0 9 9 3 3 13 15 2 14 1 9 0 9 2
6 13 15 3 13 0 2
13 9 13 3 7 1 9 2 13 13 7 13 0 2
20 9 11 11 3 13 0 9 0 9 11 11 2 15 13 0 9 0 0 9 2
12 11 13 1 9 2 15 15 13 0 9 9 2
22 13 1 9 1 0 2 16 13 2 3 3 16 0 0 2 16 3 0 13 0 9 2
31 10 9 7 9 13 0 9 2 3 13 2 12 1 10 12 9 2 15 15 2 1 9 1 0 12 2 13 1 0 9 2
20 9 12 9 13 2 16 15 13 9 0 9 1 9 7 13 9 1 10 9 2
31 3 15 13 2 3 15 13 2 16 14 15 2 15 13 1 0 0 9 3 9 2 13 13 0 9 7 13 15 0 9 2
16 10 9 7 9 13 15 0 9 2 7 15 15 2 15 13 2
20 13 15 2 16 1 10 9 4 15 13 1 9 0 0 9 13 7 1 15 2
19 13 3 3 9 1 9 1 15 2 15 13 7 15 13 0 9 1 9 2
3 9 13 0
4 11 11 2 9
15 15 13 2 16 9 0 9 0 3 13 3 1 12 9 2
12 0 3 2 16 1 15 13 14 1 12 9 2
35 3 0 13 7 9 15 2 15 13 3 0 9 1 0 9 7 3 15 13 15 2 16 15 3 3 13 9 1 9 7 0 9 0 9 2
40 1 9 2 15 9 1 0 9 13 16 0 9 0 9 2 15 13 2 7 13 3 0 13 7 9 0 9 1 11 2 13 2 14 0 9 15 13 3 3 2
18 3 13 13 0 9 1 10 9 1 15 2 15 0 9 13 9 9 2
12 7 13 7 15 2 7 15 3 13 1 9 2
20 15 3 13 0 15 13 2 16 9 9 1 9 12 1 15 13 9 3 3 2
16 13 15 9 15 13 16 4 2 7 13 15 1 15 3 13 2
12 15 3 13 1 9 0 9 7 0 9 9 2
26 13 2 16 15 9 3 13 2 16 9 0 9 13 14 1 9 9 7 10 0 9 13 10 0 9 2
13 3 13 0 2 16 10 9 9 13 10 0 9 2
43 13 4 15 2 7 1 10 0 0 9 13 9 0 9 7 1 9 13 9 1 0 9 10 9 2 15 15 13 13 2 7 3 13 7 1 9 13 3 2 3 13 11 2
6 0 9 0 9 13 2
8 0 9 3 3 13 7 15 2
25 10 3 0 9 13 10 9 3 3 2 3 1 9 13 0 0 9 0 9 1 9 1 9 12 2
16 16 4 15 3 1 9 15 13 2 16 15 3 13 1 9 2
41 3 7 13 0 9 2 15 13 1 9 10 9 2 7 3 4 15 13 3 0 2 16 0 9 3 13 7 10 9 13 0 15 7 13 2 14 15 1 15 13 2
25 7 13 4 13 3 0 13 10 9 1 9 1 0 9 9 2 3 1 11 7 11 13 0 9 2
17 15 3 13 13 9 13 1 9 7 1 10 9 10 0 9 13 2
10 16 4 15 13 0 9 1 9 9 2
4 7 9 2 2
30 16 13 0 9 13 1 9 10 9 2 15 1 9 13 1 11 2 15 3 4 13 13 15 2 15 13 1 9 3 2
15 16 9 9 13 0 9 2 1 15 3 0 13 9 9 2
35 9 1 0 9 3 13 0 0 9 1 9 0 9 2 15 13 0 9 11 2 7 13 15 9 11 2 9 0 9 11 7 9 9 11 2
51 13 2 3 13 0 3 0 2 7 11 15 3 3 2 13 16 13 2 16 13 3 14 1 9 2 3 9 13 1 9 2 15 15 13 16 9 3 0 2 16 1 10 9 3 13 7 13 1 0 13 2
31 3 4 1 15 3 13 3 1 10 9 2 16 4 15 15 13 0 9 2 7 3 4 15 3 3 13 9 15 0 9 2
17 3 16 9 13 0 7 1 9 1 15 0 3 3 13 1 15 2
8 9 11 13 13 11 7 11 9
2 11 2
26 0 9 11 11 13 0 13 0 9 10 9 0 11 2 16 4 0 9 13 7 1 9 11 7 11 2
12 9 10 9 4 13 13 9 9 1 0 9 2
18 11 13 0 13 1 9 11 12 9 1 11 2 11 7 0 0 9 2
6 13 15 3 0 9 2
33 0 9 0 9 11 1 0 11 11 11 13 3 0 9 0 11 2 16 9 11 11 12 2 13 13 15 0 0 9 1 9 11 2
9 0 9 15 13 13 12 2 9 2
13 9 0 9 0 1 11 13 9 10 9 1 11 2
13 9 1 0 13 9 9 0 11 2 0 1 11 2
31 9 0 9 1 9 11 1 9 11 11 11 3 13 9 9 14 12 9 1 11 1 10 9 2 15 4 13 1 9 11 2
12 9 15 1 9 13 9 11 1 11 11 11 2
5 0 9 11 2 11
4 11 11 2 11
23 0 9 9 9 11 11 3 1 9 9 1 12 9 0 11 13 0 9 11 7 11 11 2
18 1 0 9 15 1 0 13 1 9 11 11 2 9 9 7 9 9 2
36 7 16 0 9 13 0 2 1 9 4 15 13 2 16 3 13 9 2 16 0 9 13 1 15 9 0 2 13 11 2 11 1 11 9 11 2
20 9 11 11 13 9 1 10 0 9 11 11 7 13 1 9 7 9 0 9 2
27 0 9 13 9 0 9 13 1 11 0 9 2 10 0 9 4 13 9 1 0 7 0 9 1 12 9 2
13 1 0 9 0 9 11 1 11 15 7 3 13 2
7 9 1 11 2 9 7 9
10 11 11 2 9 11 14 1 9 1 11
2 11 2
17 0 9 13 0 9 9 7 10 9 15 13 13 0 9 0 9 2
24 3 13 15 9 0 9 2 13 3 1 11 1 0 9 9 0 9 1 11 0 9 11 11 2
20 13 9 0 9 1 9 0 9 7 3 13 2 3 3 13 13 0 9 11 2
18 0 9 15 13 3 13 2 16 11 3 3 4 1 0 9 13 9 2
12 1 11 13 9 11 0 1 0 2 0 9 2
12 0 9 12 9 13 4 3 13 0 0 9 2
30 1 10 9 11 13 1 9 1 9 7 9 1 11 2 11 2 2 15 13 15 0 9 2 16 4 13 9 7 9 2
15 0 0 9 11 1 11 4 13 1 10 9 13 0 9 2
20 0 9 11 11 13 2 16 9 0 9 1 11 13 0 9 1 0 9 11 2
17 1 11 13 13 1 15 2 16 11 13 12 2 9 12 0 9 2
9 11 9 11 13 0 9 0 9 2
11 3 3 13 13 2 15 11 3 13 11 2
12 1 15 15 15 13 13 3 9 2 13 9 2
22 13 7 9 11 1 9 11 7 13 2 16 11 7 11 13 3 3 1 9 0 9 2
31 13 10 10 0 9 7 9 13 7 3 13 2 7 9 7 9 11 13 4 13 1 11 2 7 14 1 0 9 1 15 2
12 9 3 13 1 0 9 9 1 9 0 9 2
20 9 11 7 9 11 13 1 0 9 9 2 16 13 13 9 0 9 1 11 2
23 13 15 1 9 9 1 0 9 12 9 7 1 9 13 2 16 3 13 9 9 1 15 2
10 13 15 1 9 0 9 0 0 9 2
19 9 0 9 11 11 11 13 2 16 11 13 0 9 1 9 9 1 11 2
4 11 3 13 11
2 11 2
32 0 9 3 13 2 16 0 0 9 7 0 0 9 4 1 9 9 1 0 11 1 9 12 13 7 16 3 4 13 0 9 2
31 0 0 9 11 11 1 10 9 13 2 16 0 9 13 9 1 11 2 7 13 15 1 3 0 9 1 9 7 1 9 2
12 0 12 0 0 9 13 3 0 7 3 0 2
14 3 13 9 2 1 15 13 9 1 11 9 0 9 2
16 0 0 9 1 9 9 9 13 7 13 2 16 4 13 9 2
4 9 11 2 11
6 0 9 13 0 11 11
2 11 2
35 9 0 0 9 1 9 15 13 2 16 13 0 13 0 9 2 15 13 1 3 16 12 9 9 1 9 9 2 3 7 1 0 9 11 2
8 11 11 15 13 1 9 9 2
16 13 4 9 3 13 2 13 3 11 11 2 9 9 11 9 2
12 13 15 13 0 2 13 1 0 9 1 11 2
33 11 7 13 2 16 4 0 9 13 10 9 1 9 2 15 13 13 1 0 9 0 9 1 9 2 1 15 0 9 13 1 9 2
22 0 9 4 13 13 9 13 0 9 2 16 4 13 10 9 1 9 2 13 0 9 2
14 12 0 0 9 0 9 1 11 15 13 1 0 9 2
11 10 9 13 0 2 9 9 9 13 9 2
7 1 0 9 15 13 12 2
7 9 13 3 3 12 9 2
15 11 9 13 1 11 0 9 9 2 7 9 13 2 15 2
11 1 9 3 3 13 9 0 9 1 9 2
11 1 0 0 9 15 4 1 9 13 12 2
18 15 1 12 11 2 15 3 13 1 9 1 11 2 15 13 13 3 2
19 10 9 13 9 0 2 0 9 1 9 2 15 13 3 13 1 0 11 2
5 10 9 13 0 2
17 13 10 9 2 13 3 0 9 11 11 1 0 9 11 1 11 2
10 11 13 9 1 0 9 9 1 11 2
5 0 0 9 1 11
3 0 11 2
22 13 0 9 1 0 9 1 11 15 13 0 0 0 0 9 11 7 11 2 2 0 2
23 0 9 2 0 0 0 0 11 2 0 2 2 11 2 13 1 10 9 13 1 0 9 2
18 13 0 9 2 0 1 0 9 2 1 15 0 9 15 3 4 13 2
14 11 7 13 0 9 2 3 15 3 13 1 0 9 2
31 1 0 9 13 13 1 9 9 11 0 11 2 15 4 13 1 11 7 15 3 9 11 13 16 12 1 0 9 1 9 2
23 1 9 1 0 0 9 2 15 13 3 1 15 0 9 2 15 11 13 3 1 0 9 2
5 9 9 1 11 13
5 11 2 11 2 2
22 3 15 3 3 1 9 0 9 1 11 13 3 9 14 2 9 2 7 1 0 9 2
10 0 0 9 15 13 13 1 12 9 2
18 1 9 12 4 13 9 7 1 0 9 2 15 13 7 1 9 9 2
24 9 2 16 0 9 13 9 0 9 7 13 15 16 0 2 0 7 0 2 15 13 16 0 2
24 9 0 9 9 1 9 9 3 13 1 12 2 12 2 12 2 13 3 11 9 9 11 11 2
4 0 9 13 9
2 11 2
28 0 9 13 1 9 0 9 0 9 11 11 11 2 11 2 0 11 7 3 9 2 7 13 1 15 0 9 2
9 0 9 13 0 9 1 9 11 2
18 0 9 13 1 0 9 1 9 1 9 2 0 9 7 1 9 9 2
30 11 13 0 1 9 12 9 2 15 13 13 1 9 0 9 11 2 0 1 9 0 0 9 1 9 11 7 9 11 2
13 9 13 2 16 9 13 9 11 1 10 12 9 2
4 11 13 9 9
2 11 2
38 11 3 13 2 16 13 9 12 9 9 2 1 15 4 1 0 12 9 13 9 1 9 9 7 9 0 9 1 9 2 15 13 0 9 1 9 12 2
38 9 13 0 7 0 9 2 0 0 9 9 0 0 9 2 9 11 2 15 13 1 11 1 11 2 7 9 11 2 15 13 1 0 9 1 9 12 2
25 9 2 15 4 13 13 0 9 0 9 1 9 2 4 13 9 9 9 1 9 9 1 0 9 2
1 3
29 9 12 9 0 9 1 0 9 7 1 9 0 1 0 9 13 11 11 3 1 9 11 11 13 0 9 0 9 2
14 9 15 3 13 1 0 9 1 0 9 9 13 0 2
28 12 9 1 9 9 13 1 0 12 9 9 1 11 2 15 13 7 1 0 11 16 0 9 9 3 0 9 2
28 9 0 9 13 9 2 16 4 13 1 9 2 16 16 9 13 9 9 2 0 0 9 9 13 13 3 0 2
27 9 0 11 13 15 3 1 11 3 13 9 0 9 11 2 11 2 13 7 2 16 11 13 0 9 13 2
21 1 11 0 11 13 16 15 3 13 1 11 2 16 4 0 9 11 13 1 11 2
23 0 9 1 9 13 3 0 0 9 0 0 9 2 15 15 3 13 13 1 0 0 9 2
22 9 11 2 11 13 2 16 12 0 9 1 0 9 13 9 9 7 1 0 9 13 2
11 11 7 11 15 13 0 9 9 9 11 2
21 0 9 0 9 11 2 15 13 1 9 9 2 15 3 13 13 1 0 9 11 2
17 9 13 2 16 12 9 13 0 9 1 11 11 14 1 9 12 2
34 0 9 1 0 9 11 13 3 0 9 9 2 15 13 9 0 0 0 9 2 11 2 2 1 0 9 7 13 0 9 2 16 13 2
5 11 13 2 7 13
2 11 11
30 9 0 9 1 0 11 7 1 11 2 15 3 13 2 13 0 9 3 16 0 0 9 1 9 1 0 9 1 9 2
16 7 1 0 12 9 4 1 11 13 12 9 9 1 0 9 2
12 14 1 0 11 4 13 12 9 7 12 9 2
23 7 0 9 13 9 2 9 1 9 1 11 13 9 1 9 7 9 1 9 9 9 9 2
17 14 15 9 7 9 9 1 0 9 13 0 9 9 12 9 9 2
14 7 1 0 9 2 7 1 9 15 7 0 9 13 2
22 13 15 3 15 2 16 9 13 3 0 7 16 15 15 13 7 0 9 1 9 11 2
19 10 9 1 9 1 11 13 0 9 15 2 3 15 11 13 0 0 9 2
14 1 11 7 3 3 1 11 13 0 13 9 0 9 2
14 3 16 4 13 1 10 9 3 3 2 1 9 9 2
18 9 0 9 0 11 7 11 13 3 14 16 9 9 13 7 13 9 2
9 0 9 13 1 0 11 0 9 2
18 1 0 9 3 13 7 0 9 0 9 1 0 9 7 1 0 9 2
21 1 0 9 3 13 11 13 14 1 9 1 0 9 7 9 9 0 0 0 9 2
12 1 10 0 9 7 13 1 9 13 0 9 2
29 9 9 1 0 9 11 2 1 11 2 1 15 1 0 9 3 13 0 9 2 13 1 0 9 3 14 0 9 2
11 1 11 13 0 0 9 3 3 10 9 2
21 0 9 1 0 11 4 13 14 1 9 12 2 0 9 1 0 11 1 9 3 2
15 14 3 7 13 10 9 1 0 9 7 3 1 0 9 2
21 1 0 11 7 1 11 13 0 9 9 9 9 2 0 9 9 7 9 0 9 2
9 14 3 13 10 9 1 0 9 2
14 1 9 0 0 0 11 13 0 9 11 3 9 3 2
16 9 0 9 13 9 1 11 2 15 13 7 1 0 0 9 2
9 1 0 9 9 15 13 0 9 2
18 0 9 13 3 1 0 11 0 1 9 0 9 7 1 9 0 9 2
17 1 11 7 1 11 15 1 0 9 11 13 7 9 2 7 9 2
15 9 9 7 3 0 0 9 10 9 7 0 9 13 9 2
24 11 3 13 1 9 0 9 2 1 9 9 1 0 9 7 11 2 7 0 9 2 0 9 2
8 0 9 13 13 3 1 11 2
10 7 16 3 15 3 13 9 0 9 2
11 9 1 15 13 0 9 0 12 2 9 2
5 0 9 13 11 2
29 3 1 9 13 0 9 1 9 0 9 0 11 7 1 9 0 9 1 9 2 16 4 15 13 13 1 0 9 2
19 10 0 9 2 15 3 13 0 9 9 2 4 7 1 0 0 9 13 2
11 0 9 11 15 13 1 9 9 1 11 2
12 14 11 7 11 15 13 13 0 9 1 11 2
16 9 9 1 0 7 0 9 11 13 9 0 9 3 14 3 2
25 16 0 9 2 16 9 0 9 7 1 9 9 13 3 3 10 9 7 10 9 16 1 9 11 2
13 3 13 9 0 9 1 9 0 9 1 0 9 2
7 14 13 1 0 9 11 2
8 9 1 15 13 9 1 9 2
14 3 13 7 0 9 9 2 16 4 15 9 3 13 2
21 10 9 13 3 0 9 11 1 0 0 9 7 3 1 0 11 1 0 9 9 2
29 9 13 7 9 2 16 11 13 14 0 7 0 9 9 7 16 14 0 9 9 7 9 15 13 13 3 0 9 2
23 7 3 13 3 14 1 15 2 16 15 3 0 9 13 13 10 9 1 0 9 0 9 2
16 7 16 13 9 3 13 7 1 0 2 7 1 0 0 9 2
6 13 11 13 0 9 2
6 11 11 2 9 9 9
38 3 7 3 15 1 0 9 0 9 2 1 11 2 13 9 2 15 4 13 0 0 9 2 16 3 13 3 2 7 2 4 2 14 9 13 7 13 2
25 1 9 9 15 3 13 9 1 0 9 9 2 15 3 0 9 13 14 9 2 7 0 0 9 2
20 0 11 1 12 9 13 9 2 15 1 9 1 9 0 9 3 13 9 9 2
33 0 11 2 15 13 1 0 0 9 2 10 9 1 9 13 2 16 10 0 0 9 3 13 0 9 9 7 1 0 2 0 9 2
12 9 11 11 7 1 9 13 7 13 9 13 2
11 15 13 1 0 9 9 1 9 7 11 2
14 16 4 0 9 13 2 13 15 1 9 11 3 13 2
10 3 7 3 3 0 2 7 0 9 2
36 1 9 2 16 15 0 9 11 13 15 12 9 2 15 13 14 9 3 0 2 16 14 3 13 0 15 2 4 15 13 1 0 9 13 12 2
20 9 1 15 2 16 15 13 13 1 11 10 9 3 2 15 1 0 9 13 2
30 0 1 9 9 13 3 13 9 0 9 0 0 9 2 16 3 15 13 2 16 1 12 9 13 13 13 1 0 9 2
21 13 3 1 12 9 9 0 9 2 12 1 9 9 7 15 0 1 0 0 9 2
18 4 2 14 1 0 9 13 12 12 9 2 4 3 13 0 0 9 2
14 15 7 13 2 16 9 4 3 1 3 13 1 9 2
2 3 2
18 13 15 2 16 4 13 9 1 9 0 9 7 16 4 13 1 9 2
28 9 1 9 9 13 1 11 0 3 3 7 3 4 15 3 13 1 15 2 16 4 15 10 9 13 9 9 2
20 1 0 9 0 9 0 12 9 2 0 9 2 9 9 2 4 7 13 0 2
29 3 0 9 7 13 2 16 11 3 14 0 9 13 2 7 11 11 3 13 2 16 7 1 10 9 13 9 13 2
11 1 0 9 13 9 9 13 1 12 9 2
20 16 3 13 2 13 1 9 1 9 7 13 4 7 13 7 13 1 0 9 2
35 16 4 7 1 15 10 13 13 2 13 15 1 15 13 0 9 0 9 2 11 7 9 2 1 9 3 12 12 2 12 2 9 0 9 2
13 15 4 13 3 2 13 3 0 1 10 9 13 2
11 1 0 9 4 13 1 11 0 0 9 2
29 13 15 2 16 9 13 9 3 3 3 2 7 13 2 16 10 0 9 13 1 0 9 9 1 3 0 9 9 2
13 9 0 9 4 13 13 2 16 13 10 9 0 2
13 9 9 13 0 9 1 0 9 9 7 0 9 2
24 1 9 13 1 11 9 11 1 9 7 0 9 2 1 15 13 0 9 9 12 1 0 9 2
26 1 9 1 9 13 2 16 15 1 11 3 13 0 9 3 0 7 0 9 2 15 0 9 9 13 2
16 11 15 13 1 9 2 10 9 13 1 11 13 10 0 9 2
25 16 4 13 13 1 9 1 0 0 9 2 3 4 15 13 0 9 13 1 9 1 0 9 9 2
11 7 1 9 15 13 0 9 1 11 13 2
34 0 9 3 13 9 3 2 16 1 0 9 13 1 9 9 9 2 13 15 9 9 7 9 9 11 2 11 2 15 13 9 0 9 2
14 13 0 13 2 10 9 0 0 9 3 1 11 13 2
3 9 13 11
2 11 11
17 9 7 9 13 3 0 9 2 1 15 15 13 1 9 1 11 2
20 1 0 9 7 10 0 0 9 13 7 3 13 15 3 0 2 12 0 9 2
29 3 0 9 11 11 1 9 1 0 9 3 13 2 16 9 2 0 7 0 9 9 2 4 13 4 13 7 13 2
32 0 9 3 3 13 2 16 10 9 13 2 7 13 0 9 1 9 10 9 2 9 0 9 7 9 9 7 4 13 1 9 2
24 9 15 13 13 1 0 9 2 16 9 13 10 9 7 9 15 3 13 1 9 0 9 9 2
35 1 0 9 13 0 9 2 13 9 1 9 2 1 0 9 0 0 9 15 1 12 9 13 9 9 7 9 2 1 0 9 1 0 9 2
23 9 15 13 13 9 2 1 15 1 12 9 13 9 11 7 3 9 9 0 7 0 9 2
44 9 9 13 1 9 2 3 16 1 0 9 11 11 2 13 7 13 9 1 15 2 15 13 1 9 0 9 3 13 0 9 7 9 9 1 9 7 15 3 13 10 0 9 2
31 11 9 1 11 15 1 9 0 9 7 0 9 9 0 9 13 0 9 1 0 9 1 0 9 7 3 7 1 0 9 2
14 0 9 13 1 9 11 9 1 9 0 9 0 9 2
20 3 0 9 1 0 0 9 9 0 9 2 3 3 0 9 2 13 0 9 2
15 9 0 0 9 4 1 0 9 0 9 3 3 4 13 2
21 9 0 9 1 9 11 3 13 1 0 0 9 2 9 2 1 15 15 3 13 2
13 9 3 1 9 1 9 13 3 9 9 3 9 2
15 1 9 15 13 0 9 2 15 4 3 13 1 10 9 2
20 1 0 9 1 9 12 13 0 9 0 11 0 12 0 9 1 0 12 9 2
29 0 9 1 11 15 13 13 13 0 9 2 3 13 13 1 9 2 16 4 13 0 2 1 9 9 0 2 9 2
18 1 11 15 1 0 9 3 13 9 1 0 9 9 1 0 0 9 2
21 0 9 1 9 12 3 13 2 16 9 13 1 9 9 2 9 2 9 7 9 2
11 1 12 9 3 4 0 9 13 1 9 2
14 1 0 9 1 9 12 13 3 9 13 16 0 9 2
17 11 11 13 3 9 2 16 1 9 0 9 13 11 1 0 9 2
49 10 0 2 3 0 0 9 3 13 2 16 9 13 1 9 9 2 16 1 0 9 13 9 9 1 9 7 13 15 13 3 1 9 3 0 7 0 9 2 15 15 13 7 0 0 7 0 9 2
15 10 0 7 0 9 13 9 9 1 9 0 9 3 3 2
14 14 3 3 13 2 3 15 2 15 15 3 7 13 2
6 11 3 1 11 13 2
21 1 9 11 7 0 0 9 13 9 9 7 13 2 16 16 13 2 13 1 9 2
11 1 11 15 13 13 2 16 10 9 13 2
16 3 3 13 0 9 2 16 16 13 3 2 9 9 13 3 2
9 1 11 7 3 3 7 3 13 2
25 15 14 12 9 1 12 9 2 15 13 9 1 11 2 13 13 9 0 9 7 0 9 1 11 2
18 12 2 9 12 13 9 1 9 11 2 11 1 0 11 0 0 9 2
14 1 10 9 15 12 0 9 13 9 9 1 0 9 2
1 9
11 1 9 15 0 9 13 1 12 9 1 9
5 9 1 0 2 9
17 12 0 9 1 9 13 1 0 9 0 2 9 1 10 0 9 2
7 10 9 13 3 10 9 2
18 9 9 1 10 9 3 3 13 0 9 2 1 0 9 7 3 13 2
19 1 0 9 13 10 9 9 2 16 15 0 9 13 1 12 9 2 9 2
21 15 13 15 2 16 4 1 10 9 13 13 9 9 0 1 9 0 9 0 9 2
14 9 9 1 0 9 0 2 9 13 3 3 16 0 2
22 1 3 0 0 0 0 9 9 9 3 13 2 7 15 1 12 1 12 9 2 9 2
10 9 9 15 7 13 1 12 9 9 2
9 13 15 12 12 0 9 12 9 2
11 0 9 0 9 13 1 12 1 12 9 2
17 9 9 12 15 1 10 9 13 1 12 5 1 12 1 12 9 2
15 12 9 13 15 0 2 3 9 1 9 1 9 0 9 2
30 3 15 13 1 9 0 0 11 2 0 0 11 2 11 0 9 2 11 0 9 2 11 11 2 0 0 7 0 11 2
22 0 13 1 12 9 0 9 2 13 9 9 0 1 9 2 9 2 0 9 7 9 2
21 1 9 1 9 15 1 0 7 0 9 13 7 1 9 9 2 15 13 1 9 2
20 9 0 0 11 2 11 11 2 11 7 11 13 3 1 0 2 9 1 0 2
23 16 3 4 13 2 13 1 0 9 9 9 1 0 9 0 2 9 0 12 9 2 9 2
11 3 0 9 13 7 12 12 0 0 9 2
21 0 9 2 1 12 1 12 9 2 13 0 9 9 2 1 15 4 13 0 9 2
19 1 9 1 0 9 13 0 9 10 9 2 9 9 9 12 2 14 3 2
23 1 0 0 9 1 12 9 13 7 0 2 16 3 13 9 1 0 9 0 16 1 0 2
21 16 0 2 9 13 12 0 9 1 9 1 0 9 2 0 9 13 14 0 9 2
20 0 9 12 3 0 9 15 13 1 12 2 9 2 3 13 0 9 3 9 2
3 2 11 2
2 9 9
13 9 2 11 11 2 9 9 1 0 0 9 1 11
1 9
10 1 0 9 9 4 15 13 13 9 2
38 3 13 3 12 9 15 7 13 15 2 16 13 15 15 3 15 0 2 7 1 0 9 15 13 15 0 2 15 15 12 3 13 2 9 1 9 3 2
20 3 7 3 13 9 1 10 9 1 0 0 9 1 10 3 0 9 1 9 2
6 13 15 1 0 9 2
6 13 13 1 0 9 2
11 13 13 9 1 0 9 2 7 0 9 2
32 9 13 15 9 1 9 9 13 1 9 3 0 9 7 13 13 7 9 9 2 3 15 12 1 9 1 10 0 9 13 13 2
26 9 15 1 0 9 1 10 9 1 9 13 1 9 9 9 1 9 0 0 9 1 9 10 0 9 2
12 3 15 15 13 0 0 9 1 0 0 9 2
25 0 9 13 9 1 0 9 0 1 0 9 2 13 15 1 9 1 9 0 9 1 10 0 9 2
14 9 0 9 9 13 7 9 1 9 9 7 9 9 2
28 0 9 0 9 13 3 1 9 7 1 9 2 7 7 1 9 1 0 0 9 7 13 0 1 9 9 9 2
29 0 9 1 9 13 13 1 0 9 1 0 0 9 9 9 7 0 9 11 9 0 9 0 0 9 1 0 9 2
14 0 0 9 13 9 9 1 9 1 9 0 0 9 2
12 3 10 9 1 11 13 1 12 9 0 11 2
19 3 13 0 9 1 9 2 0 9 13 10 9 3 0 9 10 0 9 2
27 3 7 13 0 9 1 9 9 7 9 9 0 1 9 1 9 0 9 2 7 7 13 9 1 9 9 2
32 10 9 15 1 12 9 9 13 1 0 9 1 9 0 9 2 0 9 7 9 9 1 9 13 0 9 1 3 12 9 9 2
20 10 9 13 1 9 0 7 9 2 1 15 13 0 9 2 7 3 9 9 2
16 2 9 1 9 4 9 1 9 10 0 9 13 1 0 9 2
20 1 15 13 9 0 9 1 0 9 7 9 9 7 3 13 0 9 2 9 2
24 0 9 1 9 15 13 1 9 10 9 7 13 1 9 0 9 0 9 1 0 9 9 9 2
30 0 9 13 3 1 0 0 9 2 15 13 9 3 13 1 9 0 9 7 1 9 1 9 9 13 10 0 0 9 2
29 0 9 9 15 13 13 9 1 9 2 9 9 7 9 1 0 9 9 2 0 9 9 7 0 9 9 0 9 2
24 9 4 1 10 9 3 13 1 9 0 9 1 12 1 0 9 7 3 13 1 0 9 9 2
20 9 9 9 13 3 0 7 7 1 9 13 13 2 16 9 0 9 4 13 2
20 9 9 7 9 4 13 3 7 3 13 0 9 10 9 7 9 1 9 9 2
24 13 4 15 15 13 9 7 0 9 9 1 9 2 15 13 3 13 1 9 0 9 1 9 2
8 9 0 9 13 0 0 9 2
14 1 0 11 13 9 9 1 9 1 12 7 12 9 2
5 0 9 2 9 9
20 9 2 9 2 11 11 2 9 2 2 0 9 12 2 0 9 1 11 2 11
1 9
19 1 0 9 4 1 9 13 9 16 9 9 0 9 7 9 0 0 9 2
16 9 15 13 0 9 2 7 2 9 2 15 13 1 9 9 2
20 9 13 9 1 9 0 9 1 0 9 0 9 9 2 9 2 9 7 9 2
12 13 2 14 9 0 9 2 13 3 1 9 2
30 9 0 9 13 1 0 9 9 1 9 2 9 2 9 7 9 7 9 1 15 0 2 16 13 9 2 9 7 9 2
10 1 0 9 15 13 1 12 9 9 2
14 1 15 0 13 9 0 9 2 1 15 0 13 9 2
15 1 0 9 13 3 0 9 2 0 9 2 9 2 9 2
36 1 0 9 13 9 0 9 2 9 1 9 2 9 2 9 2 9 0 9 2 9 1 9 1 9 9 2 16 13 0 9 2 9 2 9 2
12 3 1 10 9 13 10 9 2 9 2 9 2
11 1 9 13 9 3 0 9 7 0 9 2
10 9 7 9 13 1 9 3 13 9 2
37 9 9 7 0 9 1 9 13 1 0 9 2 3 4 7 9 13 1 0 0 9 1 15 9 9 2 3 9 0 9 13 3 13 7 3 0 2
30 1 0 15 9 7 1 9 0 15 0 9 9 0 9 15 13 7 0 9 9 7 9 13 13 9 7 13 0 9 2
37 0 9 13 0 9 7 0 9 15 13 0 9 2 0 9 7 0 9 2 0 9 7 0 9 2 0 9 2 9 2 9 1 9 9 7 9 2
19 13 13 7 0 9 2 7 14 15 2 15 4 3 13 7 13 3 0 2
22 9 7 3 9 0 1 0 9 13 13 1 10 9 13 0 0 9 7 0 0 9 2
20 0 0 9 1 9 13 0 9 7 13 15 1 15 3 3 7 1 10 9 2
32 16 9 0 9 1 0 9 13 10 9 2 13 9 0 9 2 15 4 13 1 0 9 7 4 3 13 7 1 9 9 9 2
19 9 9 1 3 0 9 2 15 13 0 9 2 13 9 1 9 0 9 2
5 9 2 9 7 9
2 11 11
23 1 9 13 1 9 11 9 9 2 9 7 9 1 9 0 9 1 9 0 9 1 9 2
28 10 9 9 2 9 2 11 11 7 9 2 9 2 11 11 1 12 9 13 9 1 9 9 2 15 3 13 2
14 11 2 11 15 13 9 7 11 2 11 0 9 9 2
25 11 11 2 1 9 9 1 9 0 9 15 13 9 13 10 9 2 15 15 1 9 3 3 13 2
25 9 11 7 15 4 4 13 2 16 4 15 1 10 9 13 1 15 2 16 9 13 13 0 9 2
6 3 13 7 9 13 2
23 1 0 9 15 13 1 0 9 2 13 3 13 0 2 10 9 13 15 13 7 15 13 2
7 13 3 1 9 0 9 2
23 10 9 13 1 12 9 0 9 2 1 0 9 9 14 1 0 9 7 9 9 1 9 2
14 15 14 12 0 9 13 13 3 12 2 3 12 9 2
25 11 11 2 3 10 9 13 13 1 0 9 2 7 15 3 1 9 2 15 13 1 9 1 9 2
17 1 0 9 15 13 2 16 10 9 13 3 0 1 9 7 9 2
11 15 15 3 13 7 1 0 7 0 9 2
18 7 16 3 13 9 0 2 3 15 13 2 16 13 0 7 1 9 2
9 3 14 0 9 14 1 0 9 2
21 11 11 2 16 4 15 3 13 10 9 12 9 2 3 4 15 13 3 0 9 2
10 7 13 12 7 3 15 13 7 3 2
26 13 15 2 10 13 9 2 12 12 3 1 9 2 15 13 2 3 12 9 9 13 9 10 9 13 2
32 1 10 9 13 9 2 3 13 9 9 7 3 1 15 13 2 7 9 2 3 15 13 9 13 2 16 4 15 9 9 13 2
17 7 3 13 0 0 9 2 15 13 1 10 0 9 12 9 9 2
7 10 9 15 3 3 13 2
17 9 13 0 2 0 7 13 0 15 13 2 7 3 13 3 0 2
23 9 15 13 1 9 7 4 13 3 1 0 9 1 9 2 15 15 13 9 1 9 3 2
6 7 15 9 13 13 2
13 3 7 9 7 1 10 9 13 9 15 1 15 2
12 11 11 2 13 7 9 2 1 15 15 13 2
9 7 3 9 9 7 9 0 9 2
20 3 13 14 1 9 2 7 7 1 9 2 15 13 13 2 3 15 13 13 2
16 7 9 1 9 7 10 9 1 9 7 13 15 13 3 9 2
22 13 15 13 2 16 9 1 10 9 2 15 15 0 9 13 2 13 1 9 10 0 2
9 11 11 2 14 2 15 13 0 2
15 7 3 9 1 0 0 9 13 14 1 9 7 1 9 2
9 10 9 13 10 9 2 9 3 2
28 15 7 10 9 13 13 0 9 2 7 15 2 15 13 2 13 9 7 13 15 7 3 15 9 1 9 13 2
10 7 16 13 3 2 3 7 13 13 2
12 9 2 15 3 13 1 9 2 13 0 9 2
26 11 11 2 1 9 12 2 3 4 13 1 0 0 9 0 9 1 9 9 2 15 3 13 10 9 2
18 13 4 3 9 9 7 1 12 9 4 1 9 13 3 0 9 9 2
6 7 3 0 9 9 2
18 13 4 12 9 1 9 2 15 15 13 1 0 9 7 1 10 9 2
16 15 13 10 0 9 1 9 2 3 15 9 13 2 7 13 2
25 11 11 2 13 4 9 2 15 13 1 9 1 3 0 0 7 0 9 2 15 13 13 0 9 2
11 3 3 1 9 1 9 9 13 15 0 2
12 13 15 9 2 15 13 0 9 1 0 9 2
19 1 0 9 15 13 9 2 15 15 13 1 15 1 9 0 9 7 9 2
23 11 11 2 1 15 13 0 13 2 16 1 0 9 1 11 13 9 9 1 0 0 9 2
13 15 4 10 9 13 7 13 15 14 1 12 9 2
11 13 4 15 16 0 9 9 9 7 9 2
9 13 4 2 15 15 13 1 9 2
16 15 13 9 7 13 15 15 1 15 0 9 7 1 9 3 2
18 13 9 2 3 15 9 13 3 7 13 9 1 0 9 7 1 9 2
8 10 9 13 3 0 2 0 2
15 9 15 13 1 15 7 13 0 9 2 15 3 13 9 2
18 13 15 0 9 7 15 15 13 2 3 16 9 1 0 9 7 3 2
3 11 11 2
8 10 9 4 13 1 12 9 2
30 9 2 15 15 13 1 9 9 2 15 13 0 2 15 13 0 1 10 0 0 9 2 7 3 3 2 7 9 0 2
16 7 9 2 15 13 0 9 7 13 15 13 14 16 1 9 2
17 11 11 2 10 9 2 10 0 2 13 12 9 7 13 0 9 2
32 11 11 2 12 9 2 15 3 13 2 13 13 1 0 9 9 2 15 13 3 0 7 13 9 2 7 13 1 3 0 9 2
15 12 9 13 9 2 15 3 13 9 7 13 1 0 9 2
33 1 0 9 13 15 2 15 1 0 9 13 1 0 9 2 7 9 0 9 2 7 1 0 15 2 15 15 13 1 0 0 9 2
31 3 13 9 2 15 13 1 9 0 1 3 0 9 2 3 2 0 9 2 7 3 13 9 0 2 15 13 0 2 9 2
5 13 10 0 9 2
8 11 11 2 13 15 12 9 2
8 12 13 0 2 9 0 9 2
43 3 2 16 9 13 9 7 9 15 15 13 1 10 9 2 13 15 3 7 13 0 9 2 7 15 13 13 15 2 16 7 10 9 15 1 9 4 13 1 10 9 3 2
23 3 10 3 0 9 4 13 1 9 1 9 2 15 13 1 10 9 9 0 0 9 11 2
26 9 2 15 15 13 0 9 2 16 1 9 10 9 4 13 0 9 2 1 10 9 3 13 10 9 2
24 11 11 2 3 13 9 1 0 9 2 16 13 10 9 0 2 3 13 0 9 13 7 13 2
16 11 11 2 7 1 15 4 9 13 2 3 15 13 7 13 2
16 11 11 2 10 9 13 0 0 9 7 13 1 15 9 0 2
18 14 16 4 15 13 9 7 16 4 13 15 15 2 7 13 15 9 2
8 13 15 2 16 13 0 9 2
11 11 11 2 13 13 9 2 3 15 13 2
23 7 15 13 7 1 0 9 2 3 13 9 0 2 0 2 15 13 1 15 0 1 9 2
18 11 11 2 3 13 9 2 15 1 10 9 13 1 0 2 0 9 2
2 3 2
11 13 14 1 15 13 9 2 7 7 9 2
4 15 15 13 2
11 3 15 13 13 9 2 9 2 9 3 2
8 3 15 2 15 15 13 13 2
22 11 11 2 10 9 2 15 13 10 9 0 9 2 13 0 9 7 15 13 9 9 2
4 13 15 0 2
23 13 1 15 2 13 1 0 7 10 9 15 13 2 13 0 9 7 15 15 1 15 13 2
7 15 15 13 9 0 9 2
18 1 0 9 15 13 0 7 0 7 3 7 13 2 15 13 1 9 2
11 13 15 13 3 9 9 9 2 3 9 2
17 11 11 2 16 10 9 3 13 2 3 15 3 9 0 9 13 2
4 13 15 13 2
15 13 15 1 9 2 15 13 1 9 9 1 10 0 9 2
18 11 11 2 13 15 0 2 7 13 1 15 9 10 9 7 13 9 2
30 13 9 2 3 13 0 9 14 3 0 2 15 2 3 13 0 2 14 1 15 2 15 13 1 10 9 13 1 9 2
5 13 15 13 3 2
15 3 3 13 12 9 2 3 15 13 13 15 1 0 9 2
9 16 4 3 10 9 1 9 13 2
39 11 11 2 13 15 3 2 1 15 15 13 2 7 9 1 9 13 14 2 16 15 13 9 0 2 7 13 1 9 1 9 2 15 13 1 9 3 0 2
5 13 15 0 9 2
8 7 15 13 3 3 9 9 2
16 11 11 13 1 10 10 9 0 7 0 3 1 12 9 7 9
2 9 9
2 0 9
25 9 9 2 0 0 9 0 0 9 13 0 9 2 9 11 11 2 12 2 2 0 9 0 9 2
30 9 1 9 1 0 0 9 1 9 0 9 15 13 1 9 9 1 10 9 1 0 2 0 7 0 9 9 0 9 2
30 9 2 14 0 9 7 0 9 2 13 9 0 9 11 11 2 3 3 9 11 11 1 11 7 0 9 0 0 9 2
64 11 11 15 1 15 9 13 13 9 1 0 9 0 9 2 10 0 9 14 3 13 15 9 7 9 14 1 0 9 7 0 9 10 9 2 7 7 1 0 9 9 7 9 2 0 9 2 3 13 9 2 7 0 9 2 0 3 3 3 11 16 3 11 2
40 13 15 3 13 7 0 1 0 9 9 1 12 9 9 2 9 1 0 0 9 13 1 9 9 2 16 13 2 13 2 14 15 15 0 9 3 13 2 2 2
28 13 0 0 9 7 3 0 9 9 9 7 9 2 7 3 9 9 1 0 9 13 9 9 1 3 0 9 2
25 16 1 10 10 9 11 11 13 0 9 1 15 9 2 13 3 3 14 1 9 2 9 7 9 2
5 7 1 0 9 2
45 16 9 1 0 9 13 7 9 0 7 10 9 0 2 13 2 14 3 1 9 9 11 11 1 0 9 2 13 15 3 3 1 10 9 13 15 1 0 9 7 9 10 0 9 2
10 1 0 9 15 13 9 0 1 9 2
25 2 13 7 0 9 2 15 4 3 14 3 3 13 9 7 9 13 15 3 2 3 15 13 2 2
25 0 2 9 7 9 0 11 2 7 11 2 13 14 1 9 14 9 0 2 7 0 2 0 9 2
2 11 11
13 11 11 2 0 9 2 0 9 1 11 7 11 2
7 13 0 9 2 11 12 2
4 13 11 11 2
8 12 9 2 9 7 9 13 2
22 9 2 0 11 2 11 11 2 15 3 13 9 0 9 0 9 0 11 2 11 11 2
3 9 0 9
2 0 9
1 9
27 9 2 1 12 9 13 9 11 11 0 0 9 0 9 2 15 13 1 3 0 0 0 9 0 11 3 2
42 16 9 13 10 0 9 7 13 3 14 0 9 0 9 2 0 9 7 0 9 2 15 13 3 12 0 9 11 11 7 11 11 2 13 15 0 9 1 9 7 9 2
21 9 1 0 9 13 0 9 2 11 2 11 7 11 2 11 2 7 0 9 9 2
21 9 13 1 9 9 3 0 11 2 7 7 13 14 9 9 2 3 13 0 9 2
41 0 9 12 2 11 2 9 9 12 2 13 16 0 9 0 9 11 11 1 9 2 15 13 11 11 7 11 7 11 0 2 15 12 15 13 3 1 0 9 2 2
17 9 15 14 3 13 14 1 3 0 9 0 0 9 7 0 9 2
44 2 16 1 0 9 15 11 13 13 9 0 0 9 11 2 1 15 15 13 0 0 9 2 1 0 9 13 13 15 9 2 16 4 10 9 13 1 0 9 2 3 0 2 2
36 1 0 2 16 3 3 0 0 9 9 0 0 7 0 9 11 2 15 13 0 0 9 2 13 9 9 2 16 10 9 13 1 3 0 9 2
52 0 9 4 15 13 13 1 9 12 9 7 3 13 0 7 3 14 0 9 1 9 0 0 9 2 0 9 2 9 2 0 11 2 11 2 11 2 7 0 9 2 0 0 2 9 2 0 9 2 3 2 2
29 9 13 13 9 9 0 9 2 3 2 11 2 11 11 2 12 14 11 7 11 2 7 13 9 3 0 11 11 2
25 15 14 15 13 1 9 2 16 9 9 13 3 3 0 7 10 0 9 13 13 3 14 0 9 2
2 11 11
8 0 9 12 2 11 2 12 2
7 9 1 11 2 0 9 2
20 9 2 11 11 2 9 11 11 2 11 11 2 11 11 2 9 2 11 11 2
16 13 2 11 11 2 11 11 2 11 11 2 11 11 7 0 2
4 0 9 0 9
11 0 9 13 0 9 7 13 1 11 7 9
2 11 11
25 0 9 7 9 11 11 15 1 9 12 3 13 0 9 7 1 9 0 9 3 1 11 3 13 2
15 1 10 0 9 15 3 13 12 9 9 7 9 1 9 2
33 1 9 12 15 13 9 0 9 9 7 3 13 0 2 9 11 11 2 0 1 0 9 0 0 9 2 1 9 0 9 1 9 2
20 3 11 1 10 9 2 15 13 10 9 2 13 1 0 12 0 9 1 9 2
23 11 13 1 9 0 9 0 9 16 0 9 2 14 9 3 13 0 9 3 14 3 0 2
11 3 15 13 1 0 9 1 9 0 9 2
6 13 1 9 3 0 2
19 9 9 4 3 13 2 13 3 13 3 1 10 9 10 9 1 0 9 2
12 1 0 9 2 9 10 9 13 14 3 0 2
32 3 9 11 11 13 1 9 1 12 9 9 2 9 11 11 13 1 9 3 15 7 9 10 9 1 0 9 13 13 3 0 2
9 3 13 0 2 16 3 0 9 2
15 7 14 9 9 1 10 0 9 2 1 15 13 1 15 2
24 1 12 10 0 9 2 0 2 3 0 2 0 7 0 2 13 1 11 3 0 7 0 9 2
19 16 1 15 13 9 1 10 9 1 0 9 2 3 13 9 10 0 9 2
17 3 9 7 13 7 13 2 7 13 7 13 2 7 13 3 2 2
15 13 0 0 9 0 0 9 2 15 10 9 13 1 9 2
11 3 1 0 9 13 0 9 7 1 11 2
12 1 9 9 15 13 0 7 0 9 10 9 2
40 7 3 13 3 0 9 1 9 1 0 9 2 13 2 14 9 10 0 9 1 0 9 2 3 13 2 0 2 9 0 0 9 13 1 0 0 9 10 9 2
17 0 9 1 9 0 0 9 15 13 1 9 12 9 0 9 9 2
28 1 10 0 9 13 9 11 2 11 2 11 2 11 2 11 2 11 2 9 11 2 11 7 9 11 2 11 2
26 10 9 0 9 13 3 7 3 2 7 3 13 9 1 11 14 1 11 2 7 7 1 9 2 2 2
14 9 9 2 0 9 1 0 11 2 13 3 0 9 2
16 16 13 1 0 9 2 15 15 13 13 14 1 0 0 9 2
8 0 0 9 3 13 13 9 2
15 9 1 0 9 1 9 13 2 14 2 3 9 0 9 2
22 1 0 11 13 3 0 9 0 7 3 0 9 2 0 13 0 0 9 7 0 9 2
10 3 0 9 13 3 0 0 9 11 2
15 1 10 9 15 1 15 15 13 9 9 7 0 0 9 2
15 7 16 13 0 9 0 16 10 2 14 10 9 4 13 2
14 9 15 13 0 9 7 3 14 14 9 0 0 9 2
31 1 10 0 9 15 13 2 16 0 0 9 3 13 9 1 3 0 9 9 2 7 13 7 1 10 9 2 15 3 13 2
10 15 15 13 0 7 0 9 7 9 2
22 15 13 7 9 10 9 2 7 0 0 9 7 3 7 10 0 0 0 9 2 11 2
10 13 0 9 0 9 7 3 15 11 2
7 10 13 9 1 0 9 2
7 1 9 9 13 9 0 2
23 13 3 2 7 3 3 3 2 2 3 0 11 2 13 0 2 11 7 0 10 0 9 2
8 0 11 3 13 13 1 9 2
17 3 4 15 13 3 1 9 12 2 7 3 13 14 1 9 9 2
17 9 13 3 0 9 1 9 7 9 2 15 13 1 9 7 3 2
10 14 3 1 10 9 13 0 0 9 2
20 3 4 13 9 1 9 0 0 9 2 7 11 7 11 13 1 0 9 3 2
19 13 1 10 9 9 2 15 1 0 9 0 13 2 7 3 15 13 3 2
17 0 9 1 9 13 0 9 9 12 2 9 11 7 9 0 9 2
12 3 15 1 15 11 2 7 3 9 2 13 2
10 9 13 2 13 9 2 15 3 13 2
7 9 13 1 3 0 9 2
28 9 3 3 1 9 13 9 1 0 7 0 9 1 9 7 9 7 14 15 15 13 2 15 3 2 15 3 2
10 12 9 13 14 3 0 9 1 9 2
24 0 15 3 13 2 16 13 0 0 9 2 15 15 13 13 9 11 1 11 2 11 1 9 2
30 10 0 9 2 3 0 9 11 11 0 9 2 13 3 7 3 13 1 0 9 1 0 9 7 13 15 3 10 9 2
8 3 15 7 1 0 9 13 2
15 9 15 14 13 2 16 0 9 7 13 0 2 7 0 2
8 0 9 13 3 0 1 9 2
10 3 15 1 9 1 9 13 0 9 2
12 3 15 13 2 16 1 9 3 1 9 13 2
5 13 15 3 9 2
10 3 4 3 13 13 9 7 9 9 2
7 7 0 9 3 3 13 2
5 7 1 0 9 2
16 3 11 11 2 3 13 10 3 0 9 2 0 15 13 9 2
29 10 0 9 1 0 9 9 1 9 4 1 0 2 0 9 3 13 2 3 7 15 13 0 2 7 15 7 0 2
11 3 13 1 9 11 10 9 12 0 9 2
5 1 15 13 3 2
11 1 11 4 3 13 9 0 9 1 11 2
8 13 2 16 15 3 13 9 2
9 3 2 1 9 2 13 15 0 2
3 7 0 2
7 3 15 3 13 10 9 2
7 7 9 0 9 2 2 2
6 9 13 1 0 9 9
7 9 13 9 0 0 9 9
15 0 9 0 9 13 1 0 9 9 7 0 9 9 11 2
15 0 9 13 9 0 2 7 1 10 9 3 0 0 9 2
25 10 9 9 2 9 2 9 7 9 13 0 9 1 0 2 15 13 9 1 12 9 0 12 9 2
18 16 0 9 13 1 9 9 0 9 9 9 2 15 13 12 9 0 2
19 3 15 13 0 9 2 9 1 0 9 2 1 0 9 7 1 0 9 2
15 0 3 0 9 13 9 9 2 1 15 13 12 9 9 2
13 1 0 9 13 1 0 9 11 1 12 9 9 2
16 13 15 9 0 1 0 9 2 3 15 13 9 12 9 0 2
22 1 0 9 13 9 11 2 9 7 11 2 15 13 1 10 9 3 1 12 9 9 2
8 12 9 0 13 10 9 9 2
25 1 9 3 13 0 9 11 2 15 1 0 13 12 9 0 2 1 0 0 9 3 12 9 9 2
25 0 9 13 9 11 1 12 9 9 7 0 3 0 9 13 11 2 1 15 15 13 12 9 0 2
18 15 3 16 11 13 0 9 1 9 1 12 9 2 3 13 0 9 2
29 11 13 3 0 9 9 9 2 15 13 1 0 9 2 12 5 2 7 1 9 1 0 0 9 2 12 5 2 2
11 0 9 13 1 0 12 3 0 0 9 2
15 0 9 13 16 0 12 9 0 2 11 7 11 12 9 2
9 1 9 0 9 13 9 11 11 2
29 1 0 15 13 12 9 0 2 3 9 0 12 9 2 12 5 2 7 9 1 9 1 0 9 2 12 5 2 2
17 0 3 0 9 13 11 11 2 15 13 0 0 0 0 12 9 2
16 1 0 9 13 0 11 11 2 15 16 0 13 12 9 9 2
14 3 9 2 12 5 0 2 13 10 9 9 16 0 2
35 3 1 9 15 1 0 9 13 0 9 2 7 11 1 12 9 2 1 0 9 1 0 9 11 1 12 9 7 0 13 11 1 12 9 2
18 12 9 0 13 9 11 2 1 12 9 13 9 11 2 11 7 11 2
3 2 11 2
9 9 9 13 3 13 1 9 0 9
19 9 9 15 4 1 9 0 0 9 13 1 0 9 9 0 9 11 11 2
10 11 15 3 13 9 9 9 11 11 2
32 13 1 0 9 1 9 0 9 2 11 2 11 12 2 13 15 11 1 9 9 9 2 15 13 1 0 9 13 9 0 9 2
21 11 3 13 9 11 11 2 15 12 2 9 10 9 9 11 3 13 2 0 9 2
19 9 1 9 1 11 15 3 13 1 9 2 16 9 4 13 1 0 9 2
30 16 4 13 2 13 13 3 3 2 13 11 7 13 2 16 4 9 13 13 9 9 3 1 0 9 9 12 2 9 2
3 2 11 2
1 3
11 9 11 1 11 15 1 0 0 9 13 2
22 0 0 0 11 1 9 11 11 13 1 0 9 1 0 9 3 3 7 12 2 9 2
6 0 9 3 13 10 9
15 1 9 12 2 9 13 1 10 9 1 0 9 0 9 2
41 1 9 11 12 2 15 4 1 9 9 13 13 9 13 3 0 9 9 2 15 1 0 0 9 13 3 2 0 9 11 1 9 0 0 0 0 9 0 15 9 2
22 12 9 0 9 13 0 0 9 7 0 9 4 1 15 1 9 13 13 7 0 9 2
11 3 1 15 13 0 9 0 9 11 11 2
27 1 10 9 15 13 3 1 9 2 16 4 9 13 9 9 1 9 0 9 2 1 0 9 12 9 2 2
11 1 0 9 4 15 15 13 9 0 9 2
28 11 13 7 13 2 16 9 13 1 3 0 0 9 2 15 4 13 13 9 12 7 0 9 10 0 9 9 2
12 9 1 9 0 9 15 13 7 0 0 9 2
56 1 9 13 1 11 12 0 0 9 2 15 13 9 1 0 9 1 0 1 0 9 2 4 1 15 13 3 9 9 1 9 2 0 9 2 9 12 9 2 9 2 0 9 15 13 2 3 15 13 9 2 9 10 0 2 2
68 0 9 13 1 0 9 7 0 0 9 2 3 0 11 2 0 2 9 1 11 2 9 12 2 0 9 2 9 2 9 2 7 0 7 0 9 2 13 1 9 11 2 0 9 1 9 7 0 9 0 9 0 7 0 0 0 2 9 0 11 1 9 0 9 3 2 2 2
13 0 9 13 0 9 9 9 0 0 9 11 11 2
14 0 0 9 15 1 9 1 0 9 13 1 0 9 2
41 1 9 9 15 9 13 13 3 0 0 9 0 11 2 13 0 9 2 2 0 0 9 11 3 9 7 12 9 0 9 1 9 11 11 9 11 11 1 0 11 2
29 1 9 11 2 1 10 9 13 9 1 0 9 0 9 1 9 11 2 11 11 13 2 16 9 3 3 13 13 2
13 11 15 1 0 9 13 12 9 2 11 7 11 2
11 13 1 15 3 0 2 7 3 3 0 2
8 15 3 13 0 9 3 3 2
8 3 4 13 13 1 9 9 2
3 2 11 2
6 0 9 13 2 2 2
8 2 11 12 2 12 2 12 2
22 16 13 3 0 0 9 0 9 7 10 0 9 1 10 9 13 2 10 9 15 13 2
21 13 10 9 1 9 7 1 9 3 2 7 13 15 2 16 13 15 16 9 9 2
33 15 1 15 13 2 16 1 0 9 2 3 7 1 9 2 15 13 9 13 2 16 9 3 3 3 0 13 1 12 0 9 0 2
17 1 10 9 13 3 0 1 9 13 9 0 7 0 1 12 9 2
18 16 7 1 9 13 2 13 4 2 1 10 0 9 2 13 9 0 2
23 13 2 16 0 9 0 9 2 15 13 1 15 9 2 13 1 9 2 7 3 1 9 2
37 1 9 9 9 7 1 10 9 1 0 9 15 7 13 2 16 0 9 2 3 9 0 9 9 2 13 9 14 0 2 7 3 0 1 1 9 2
19 3 15 13 2 16 0 9 3 9 13 2 7 13 13 9 3 1 9 2
21 3 15 3 13 0 9 10 9 13 2 3 16 15 15 13 10 9 13 0 9 2
12 0 9 13 9 0 0 9 1 9 7 9 2
20 9 15 13 3 0 2 7 15 1 15 4 13 1 0 9 1 9 0 9 2
17 3 13 7 3 1 9 2 16 4 15 7 15 9 13 3 13 2
22 14 16 4 3 1 10 9 1 9 1 0 15 13 10 9 7 10 9 1 10 9 2
21 15 15 3 3 13 2 7 15 15 13 2 16 0 0 9 13 10 9 3 15 2
6 1 9 11 11 2 11
4 9 2 2 2
8 2 11 12 2 12 2 12 2
26 3 1 9 2 12 4 15 13 2 16 15 13 3 0 9 2 16 4 0 9 13 10 9 1 9 2
25 7 0 9 1 15 13 3 13 7 13 2 16 4 1 0 9 13 1 9 9 0 9 7 9 2
6 1 0 9 13 4 2
22 16 15 3 13 2 16 15 3 13 2 3 15 13 2 10 9 13 7 16 15 13 2
14 3 1 9 9 4 15 13 13 2 16 13 9 9 2
14 13 9 2 16 15 1 10 9 13 9 1 0 9 2
12 3 13 9 1 9 2 15 15 13 3 13 2
11 13 15 15 2 16 15 0 9 13 9 2
23 13 2 16 15 9 13 10 9 2 0 1 0 9 2 15 3 10 0 9 1 9 13 2
6 1 9 11 11 2 11
5 0 9 2 2 2
8 2 11 12 2 12 2 12 2
12 1 9 1 0 9 3 13 7 10 0 9 2
29 3 2 16 15 13 2 16 15 1 9 13 9 7 0 2 0 7 3 0 0 9 2 13 9 10 0 0 9 2
21 13 15 1 9 12 1 9 1 9 0 9 9 11 1 9 0 9 1 9 11 2
25 11 13 0 11 7 11 7 0 9 0 9 2 0 9 2 0 0 9 7 3 0 9 2 2 2
16 16 10 9 13 15 1 9 2 13 15 3 2 7 3 13 2
16 15 7 13 0 9 9 7 13 9 2 9 7 9 1 9 2
17 9 15 2 14 2 10 9 13 1 0 7 0 9 7 0 9 2
6 1 9 11 11 2 11
4 12 9 1 9
22 1 9 0 9 15 13 12 9 3 2 11 12 2 12 2 2 2 16 13 0 9 2
41 13 2 16 15 1 10 9 13 16 0 0 7 0 9 9 0 9 2 9 2 9 9 11 2 0 0 9 2 11 11 7 9 11 2 11 7 0 3 0 9 2
18 11 7 1 15 0 9 0 9 13 12 2 9 0 9 9 1 11 2
12 3 13 11 9 10 3 0 9 1 0 11 2
6 3 13 9 9 11 2
19 15 10 0 9 13 3 9 9 2 0 11 2 7 0 9 3 0 11 2
12 9 1 9 13 10 0 9 1 15 0 9 2
9 3 4 9 13 3 0 0 9 2
13 3 11 13 7 13 15 3 2 16 15 13 3 2
21 3 2 16 1 10 9 13 12 9 7 15 2 15 15 13 2 13 3 3 9 2
13 7 15 0 7 3 13 10 9 7 9 1 11 2
20 7 15 15 13 2 16 4 15 1 15 7 11 13 0 9 2 7 7 9 2
16 3 4 15 13 1 10 9 11 1 9 1 11 7 1 11 2
10 12 9 13 13 0 9 10 0 9 2
10 11 13 1 0 9 1 9 0 9 2
20 7 3 15 13 1 9 11 2 11 7 1 9 1 9 0 9 0 9 11 2
25 1 9 13 0 9 9 9 2 15 15 1 15 1 9 1 11 13 1 9 0 9 7 9 9 2
41 13 4 15 2 16 4 10 9 13 1 10 9 9 1 9 9 7 9 0 0 9 2 9 9 0 9 7 3 3 9 1 10 2 16 4 1 9 13 9 11 2
26 13 4 15 2 16 4 0 9 9 10 9 13 3 2 7 3 1 0 9 2 13 15 15 7 9 2
11 13 15 1 9 7 13 0 9 1 11 2
20 3 15 13 1 9 9 2 3 7 1 9 2 15 4 13 13 0 10 9 2
38 13 1 15 2 16 4 15 13 1 0 9 9 0 9 2 15 13 16 9 11 1 11 2 1 9 1 11 2 1 11 2 11 2 11 7 0 11 2
6 1 9 11 11 2 11
6 9 0 9 13 3 0
47 0 9 9 0 9 7 9 0 9 2 1 15 1 10 9 9 9 3 13 2 11 12 2 12 2 2 13 11 2 11 1 0 9 9 9 2 15 1 9 0 9 0 9 13 3 0 2
20 0 9 0 9 15 1 9 1 9 12 2 14 1 10 0 9 2 3 13 2
27 3 2 1 0 9 1 12 5 9 9 2 12 2 9 12 5 2 9 1 9 9 1 12 5 7 3 2
35 16 15 1 9 10 9 13 9 10 9 2 13 0 13 2 16 1 9 0 9 4 9 9 1 0 9 13 0 0 9 1 0 0 9 2
21 1 10 9 4 10 9 13 2 1 0 9 1 0 9 2 13 10 0 9 9 2
13 10 9 13 0 2 9 0 9 13 3 9 9 2
10 3 13 0 13 1 9 12 0 9 2
29 10 9 13 0 1 9 0 9 0 9 2 15 13 1 9 9 0 2 9 2 0 9 2 15 9 3 2 2 2
35 13 0 2 16 13 1 10 9 13 2 3 3 2 10 9 9 10 9 2 15 13 1 9 1 10 9 2 16 4 10 9 10 9 13 2
24 13 0 2 16 1 9 0 9 13 10 0 9 0 9 1 0 9 0 9 7 10 0 9 2
35 1 9 12 9 13 10 9 7 1 0 9 2 14 1 0 2 7 13 7 0 2 16 9 13 13 0 9 2 7 14 9 0 9 9 2
27 1 9 3 0 0 0 9 15 13 0 0 9 2 1 15 13 3 2 9 9 9 0 9 1 0 9 2
10 0 15 13 1 9 1 0 9 11 2
29 1 9 12 4 13 9 1 9 2 15 13 15 9 9 9 7 9 0 9 1 9 1 9 12 1 9 2 12 2
19 13 3 0 0 9 9 0 9 0 9 1 9 2 0 1 11 7 11 2
6 7 3 13 9 0 2
18 15 7 13 2 16 1 0 9 15 15 0 0 9 13 1 0 9 2
20 1 10 0 9 13 0 13 3 0 0 0 9 2 3 0 9 9 0 9 2
13 1 9 9 2 11 11 2 9 2 2 9 9 11
16 1 9 0 9 4 3 13 9 9 2 9 13 7 9 0 9
1 9
17 0 9 0 2 0 9 11 11 11 13 9 0 9 2 9 11 2
5 9 11 11 2 11
12 0 11 2 3 2 1 9 1 12 1 0 9
5 9 11 11 2 11
1 3
15 1 0 11 11 13 9 11 1 9 9 1 9 11 11 2
14 0 9 9 0 2 11 0 15 3 1 0 9 13 2
7 13 15 9 11 11 11 2
15 9 0 11 0 11 15 13 0 9 11 11 7 11 11 2
12 0 9 11 11 13 9 1 9 0 0 11 2
11 13 15 3 12 9 1 9 1 0 9 2
2 11 13
3 0 11 2
12 0 9 11 13 7 3 1 0 9 0 11 2
24 11 13 13 3 1 9 2 7 10 0 9 13 0 13 9 12 9 9 2 15 0 11 13 2
5 12 9 9 1 9
7 11 2 11 2 11 2 2
27 3 0 9 7 9 12 2 12 0 9 1 11 13 3 12 9 1 0 9 9 9 11 2 12 1 11 2
13 1 0 0 9 13 11 1 9 11 12 2 12 2
13 3 13 1 9 9 11 2 11 2 12 9 2 2
6 11 2 11 12 2 12
6 9 1 15 13 3 2
25 3 1 12 9 9 4 13 11 7 9 13 1 9 2 16 0 9 1 0 13 1 0 9 11 2
25 10 9 13 1 9 0 12 3 2 16 4 13 12 9 9 12 1 12 2 13 11 2 11 2 2
11 1 0 12 9 13 0 9 12 2 12 2
45 3 2 16 15 3 3 13 1 0 9 11 2 13 0 0 9 9 11 2 13 1 0 7 13 2 16 1 0 9 9 9 1 9 13 2 7 7 15 3 13 9 1 0 9 2
11 3 0 11 15 3 1 9 13 1 9 2
14 1 0 12 9 13 11 9 7 3 3 11 13 9 2
4 9 13 9 2
30 9 15 3 13 14 11 2 15 1 12 2 9 1 9 12 1 12 13 1 9 9 7 1 3 0 9 13 11 0 2
15 1 10 9 13 7 10 9 9 7 3 13 0 9 11 2
9 1 0 9 1 9 13 7 0 2
35 1 9 2 3 15 13 2 16 9 13 9 9 1 10 9 2 13 1 9 0 9 1 0 0 9 9 11 7 13 15 14 1 0 9 2
33 1 10 9 13 0 9 11 1 9 13 10 9 7 13 15 3 3 0 9 1 0 0 9 7 0 9 9 7 9 1 12 9 2
18 1 10 9 13 3 3 2 16 3 11 11 13 1 0 9 3 3 2
23 1 9 1 9 13 1 11 14 9 7 13 15 1 9 11 2 15 15 3 13 0 9 2
21 9 12 11 2 15 13 0 0 9 1 11 2 15 1 12 2 9 13 0 9 2
30 15 4 13 3 13 1 0 9 2 11 3 13 1 11 2 2 7 1 0 9 9 4 3 1 9 13 7 0 9 2
7 0 9 2 11 2 11 2
18 11 11 2 9 11 2 13 15 3 0 9 16 0 1 11 7 11 2
24 9 9 13 1 0 9 2 15 15 3 13 2 3 16 15 2 16 15 3 13 13 1 9 2
18 11 11 2 9 11 2 9 13 3 3 2 13 4 15 16 1 9 2
30 11 11 2 9 11 2 10 9 15 3 3 13 1 9 2 13 1 15 3 12 9 2 15 1 10 9 13 13 13 2
13 13 4 9 0 9 1 9 7 9 15 3 13 2
6 11 2 11 12 2 12
6 0 9 13 9 0 2
15 11 13 3 1 12 2 9 9 1 9 2 15 13 11 2
17 0 9 0 9 13 9 2 7 7 11 13 1 9 14 0 9 2
4 9 12 2 9
4 11 9 13 4
5 11 2 11 2 2
14 11 13 9 1 0 9 1 0 9 11 1 11 11 2
48 1 9 11 2 10 9 4 0 9 13 9 11 2 11 2 9 0 9 2 11 13 2 16 9 11 1 0 9 11 3 13 2 7 16 4 11 11 1 9 13 2 16 4 13 1 9 11 2
14 3 11 1 11 13 11 9 10 0 9 9 0 9 2
10 15 15 13 1 0 9 0 2 13 2
25 1 9 9 9 4 11 13 0 9 9 1 0 9 0 9 11 2 15 15 13 7 0 15 9 2
3 9 1 11
2 11 2
16 3 1 9 13 9 9 1 11 3 1 12 7 13 12 9 2
27 9 0 0 9 13 1 9 0 0 11 1 12 9 3 16 1 9 9 12 2 15 13 9 1 12 9 2
18 1 15 15 9 9 1 0 9 11 13 1 12 2 3 1 12 9 2
3 9 1 9
5 11 2 11 2 2
23 1 0 0 9 15 1 9 12 2 9 13 0 9 9 0 9 0 0 9 7 0 9 2
30 0 9 13 9 1 9 2 15 13 10 0 9 9 1 12 9 1 3 0 9 2 15 15 13 1 11 9 1 11 2
30 0 9 9 11 13 0 9 9 9 2 12 2 12 9 2 9 1 0 9 11 12 2 2 12 2 12 2 1 11 2
3 0 0 9
5 11 2 11 2 2
29 9 9 0 9 0 9 2 12 2 12 2 9 1 12 9 2 15 13 7 13 3 0 9 9 0 9 11 11 2
27 1 11 15 13 0 9 1 0 9 11 2 11 2 15 13 1 9 0 9 3 9 0 9 9 1 11 2
18 7 7 0 9 13 9 2 16 10 9 15 13 14 1 0 0 9 2
70 1 0 9 13 15 9 11 1 9 1 11 7 0 9 11 11 2 0 1 9 11 11 2 9 0 9 1 11 11 11 2 0 11 11 2 15 3 13 0 0 9 11 2 11 2 11 11 2 10 9 11 2 15 15 3 3 13 0 9 2 0 0 9 11 7 0 0 9 11 2
36 11 11 2 15 1 9 13 3 12 9 1 11 7 3 12 1 11 2 15 0 9 1 0 9 3 13 1 0 9 2 7 9 13 3 13 2
16 3 3 13 9 0 9 2 15 7 1 10 0 9 15 13 2
9 15 0 4 1 9 10 9 13 2
25 1 3 0 9 0 9 9 13 9 1 0 9 9 2 7 13 15 3 2 16 13 1 0 9 2
21 16 13 3 13 9 1 10 9 2 13 3 1 12 7 3 1 12 9 2 2 2
16 0 9 1 10 9 13 7 0 9 13 3 0 2 13 11 2
6 11 7 11 3 1 9
10 11 1 0 11 3 16 3 13 1 9
8 0 9 11 1 0 11 11 11
53 1 12 9 2 15 13 1 12 2 9 0 0 2 13 7 12 0 9 11 11 2 13 11 11 12 2 12 2 12 2 12 2 7 11 11 2 13 1 11 11 12 2 12 2 12 2 12 2 12 2 12 2 2
42 0 9 0 0 9 11 11 11 13 1 0 9 7 3 16 3 13 1 9 2 3 1 12 2 9 1 9 12 2 12 2 12 2 12 2 12 2 12 1 11 11 2
26 3 9 1 9 13 0 0 11 2 12 2 9 9 11 2 0 2 0 9 1 11 2 12 2 2 2
23 14 15 13 7 9 2 13 15 3 0 2 13 15 11 2 15 15 1 9 9 13 13 2
7 10 0 9 13 11 11 2
14 0 9 0 9 11 2 12 2 2 15 3 3 13 2
17 3 15 7 13 2 13 1 9 1 11 2 12 2 2 0 9 2
21 7 15 1 0 9 13 2 15 15 3 1 9 10 0 9 1 0 9 9 13 2
18 3 15 1 9 13 11 11 2 1 9 0 9 12 2 9 0 9 2
15 10 9 4 15 13 14 3 1 9 7 13 4 3 0 2
25 11 15 3 13 2 1 11 15 13 9 7 3 3 15 16 11 13 1 9 2 13 1 9 11 2
37 1 0 9 13 1 10 9 12 2 12 7 12 2 12 2 3 15 15 0 9 3 13 7 13 15 7 9 0 9 12 2 12 2 3 9 13 2
35 11 13 3 14 2 9 2 7 14 3 10 9 2 13 15 12 9 2 9 2 9 2 2 2 7 15 1 9 13 9 2 13 0 11 2
32 9 1 12 2 9 13 3 10 0 9 2 1 1 15 2 16 0 10 9 13 0 9 11 2 14 3 4 10 0 9 13 2
15 14 11 2 12 2 9 11 2 13 1 0 0 0 9 2
24 3 13 3 1 9 11 11 2 3 15 1 9 13 2 7 12 2 9 3 1 9 9 13 2
36 13 15 3 1 9 0 9 9 1 11 2 12 2 2 2 3 9 13 11 0 9 2 7 15 15 14 13 1 9 2 7 13 15 0 9 2
48 13 15 2 16 9 13 14 1 0 9 9 2 15 4 13 2 14 2 7 1 10 9 13 2 2 13 1 9 9 1 9 11 2 7 16 13 2 16 9 4 15 3 13 13 7 1 9 2
24 3 0 9 13 0 9 2 1 15 13 3 12 2 12 2 7 1 12 0 9 15 3 13 2
3 11 1 11
2 11 2
38 1 0 9 11 1 9 1 11 2 12 2 9 2 13 1 9 7 11 1 11 2 1 9 9 1 12 9 13 9 11 7 11 7 0 11 2 11 2
18 1 9 9 4 13 9 11 2 16 15 1 11 13 9 9 0 9 2
6 1 9 13 7 11 2
3 9 1 11
2 11 2
26 0 9 1 0 9 12 2 9 0 0 9 15 13 1 11 2 3 0 11 13 0 11 12 2 12 2
4 0 9 1 11
6 0 11 2 11 2 2
16 16 11 15 3 1 10 9 1 0 0 13 0 9 11 11 2
19 11 3 13 1 9 0 9 1 0 11 2 15 15 14 10 9 13 13 2
19 3 15 4 13 2 7 13 1 15 9 9 7 13 15 2 16 9 13 2
20 7 3 13 15 13 2 9 3 13 0 1 9 2 16 15 4 13 13 9 2
12 13 15 1 15 0 2 16 3 13 9 1 2
28 3 13 1 9 9 0 9 2 16 15 13 2 1 9 9 13 3 0 13 1 0 11 9 2 13 9 11 2
14 1 0 9 15 4 3 13 13 7 9 0 9 11 2
5 1 9 15 13 13
5 11 2 11 2 2
13 1 9 3 15 3 13 2 1 9 13 7 9 2
34 1 15 15 13 13 2 7 16 4 13 2 16 15 13 3 3 2 13 1 0 9 1 0 2 11 2 12 2 12 2 9 11 11 2
22 0 15 1 9 1 9 11 0 9 13 2 1 0 9 13 12 9 9 12 2 12 2
19 11 3 13 9 1 9 3 9 7 1 0 9 14 0 9 1 0 9 2
34 9 13 9 1 3 0 0 9 2 15 10 9 15 3 1 9 9 13 1 10 9 1 0 9 7 9 15 10 0 9 3 13 13 2
12 16 7 11 13 9 11 2 13 1 15 9 2
9 3 15 1 9 9 13 0 11 2
19 1 12 9 15 7 13 9 1 11 2 15 15 1 0 9 3 3 13 2
43 13 2 16 1 10 9 13 3 2 1 15 13 3 9 2 13 1 9 9 11 7 1 0 9 1 9 13 2 9 0 9 13 12 9 0 9 2 15 13 1 10 9 2
4 0 0 0 9
2 11 2
15 0 0 0 0 9 13 1 9 1 11 1 11 9 11 2
22 9 9 2 0 7 0 9 13 1 12 2 9 0 9 12 9 1 9 9 2 9 2
24 1 11 15 13 2 16 9 9 1 0 9 13 0 16 3 2 7 2 3 12 9 3 2 2
6 9 9 13 9 9 2
33 3 4 15 3 13 1 0 0 9 0 1 11 1 11 2 16 1 15 10 0 9 13 1 0 9 13 2 13 9 9 11 11 2
17 1 9 9 13 1 0 0 7 0 0 9 7 9 7 9 9 2
4 0 9 1 9
5 11 2 11 2 2
20 1 0 9 13 1 9 1 9 11 2 11 2 12 2 12 2 9 12 9 2
31 13 4 15 13 1 9 7 15 15 3 13 2 16 1 9 12 2 12 2 3 4 15 13 1 9 2 13 11 1 9 2
14 9 2 16 15 9 13 9 2 13 15 0 9 11 2
24 1 0 9 13 1 9 16 9 7 13 3 2 16 15 9 11 13 3 1 10 9 1 9 2
11 16 4 15 13 2 7 4 13 1 9 2
29 7 15 13 3 2 13 0 9 7 13 2 16 9 13 13 1 15 2 16 9 13 2 7 13 13 1 9 13 2
6 7 15 9 3 13 2
16 13 2 16 15 9 3 13 2 7 13 15 1 9 13 15 2
17 12 1 9 4 13 1 0 0 9 2 3 13 4 9 13 3 2
18 9 15 3 13 9 9 2 9 3 13 1 9 7 15 13 1 9 2
16 3 13 1 9 0 0 7 15 2 9 2 13 1 9 9 2
9 13 2 15 15 1 15 13 13 2
25 0 9 0 9 4 13 2 10 9 13 1 9 9 3 1 9 7 9 15 3 13 1 9 9 2
23 7 15 3 1 10 9 2 16 1 9 1 10 9 13 0 12 9 2 16 11 0 9 2
8 0 13 12 0 9 1 9 2
22 13 9 11 7 1 9 13 1 11 2 15 10 9 13 9 0 12 9 2 9 11 2
16 15 11 13 0 2 16 4 15 13 2 3 4 9 14 13 2
24 1 9 13 1 15 0 9 2 16 3 1 15 13 3 9 2 11 2 11 2 11 2 11 2
19 1 11 15 11 3 1 9 13 2 13 1 9 9 1 9 9 11 11 2
8 11 13 1 9 3 0 9 2
14 3 13 1 9 13 9 7 13 9 1 9 7 9 2
26 3 1 9 2 0 12 9 2 9 2 9 2 2 15 10 9 13 7 13 15 13 1 9 7 9 2
19 13 7 9 2 16 1 12 0 9 13 0 0 9 1 9 2 13 11 2
27 9 1 9 13 1 0 9 11 2 1 0 9 13 1 9 1 0 9 9 9 1 11 2 14 3 0 2
47 11 13 9 1 12 0 9 2 1 15 13 12 9 2 11 2 11 2 1 12 9 13 0 9 9 2 7 11 2 15 13 0 9 3 1 15 2 16 13 1 0 0 9 1 12 9 2
6 11 12 2 3 1 11
5 11 2 11 2 2
14 0 9 15 1 9 13 12 0 9 11 11 11 11 2
18 15 1 15 13 2 16 13 9 0 0 2 9 7 3 9 11 11 2
33 13 3 0 7 0 9 2 16 13 9 1 0 9 9 2 13 0 9 2 7 16 15 13 1 10 9 2 13 3 16 0 9 2
11 7 9 1 9 12 13 1 9 11 0 2
18 3 0 2 15 15 11 1 9 1 11 13 2 13 0 9 1 9 2
15 1 9 4 13 1 9 9 2 1 15 4 13 0 9 2
20 15 13 1 9 9 2 7 3 7 7 4 15 13 1 9 14 1 12 9 2
24 9 4 3 13 13 3 1 9 1 0 11 2 7 9 15 13 9 9 7 15 0 9 13 2
7 13 9 11 1 15 9 2
3 3 3 2
7 3 1 15 13 9 3 2
8 1 15 13 1 15 11 0 2
17 13 0 9 2 13 13 1 9 7 13 15 1 9 12 1 12 2
9 1 9 7 9 13 1 15 3 2
7 3 4 15 13 1 9 2
4 16 9 3 2
13 1 9 4 13 1 11 2 1 0 9 1 11 2
22 1 15 4 13 3 2 3 1 0 9 2 3 11 13 1 11 7 15 13 1 11 2
18 1 9 13 2 1 11 15 3 13 2 3 4 3 13 1 12 9 2
8 7 3 13 2 16 3 13 2
6 9 15 1 0 9 13
11 11 2 11 2 11 2 11 2 11 2 2
50 7 1 12 2 9 2 1 0 9 7 0 12 2 2 0 0 9 2 15 15 13 1 9 7 1 9 2 13 9 1 0 11 1 0 9 7 13 2 16 4 16 0 9 13 13 1 9 0 9 2
15 1 9 1 11 2 12 2 12 2 15 13 3 9 9 2
28 0 15 3 1 12 2 9 13 3 13 7 13 3 9 9 11 2 15 13 3 1 0 9 1 12 9 9 2
10 1 0 9 3 13 7 3 9 11 2
25 3 13 12 2 12 1 9 0 9 1 11 1 11 2 15 15 3 1 9 13 3 1 0 9 2
41 15 11 2 15 4 1 9 12 1 0 9 1 9 1 0 9 13 3 1 9 9 2 1 0 9 13 2 16 10 9 1 12 2 9 1 11 13 3 14 0 2
26 3 13 1 0 9 11 2 11 12 2 12 2 16 12 9 13 11 2 15 3 13 7 1 0 9 2
24 7 3 13 0 9 11 1 9 0 9 2 0 13 3 1 9 2 1 9 15 3 13 0 2
25 10 0 0 9 2 11 2 11 2 11 2 15 13 13 1 0 9 0 1 0 0 9 0 9 2
9 3 4 3 13 3 12 0 9 2
12 13 15 3 9 2 16 0 9 2 13 11 2
21 15 10 9 11 13 7 1 9 0 9 2 13 4 0 9 7 13 4 7 9 2
14 9 12 0 9 2 16 13 1 9 2 15 13 13 2
15 0 9 10 9 13 9 11 1 11 1 11 12 2 12 2
19 11 1 10 9 13 9 14 1 0 9 1 11 7 1 9 13 0 9 2
16 1 12 9 1 9 12 2 12 1 11 4 13 3 0 9 2
14 9 10 9 13 0 9 1 9 2 13 0 9 11 2
16 11 7 13 7 9 9 2 16 9 1 9 13 11 0 9 2
28 13 15 0 9 2 15 4 13 9 13 1 9 2 3 15 15 13 2 13 0 9 1 0 9 0 9 11 2
22 11 1 0 9 3 14 13 2 3 1 11 2 7 1 9 15 13 3 1 9 9 2
33 0 9 11 13 9 10 9 7 1 0 9 2 1 15 1 10 0 2 0 7 0 9 3 13 2 13 10 9 9 1 10 9 2
26 11 2 9 11 13 9 3 1 9 10 9 2 13 4 3 12 9 2 1 15 13 10 9 1 9 2
10 3 15 13 2 16 9 13 9 9 2
4 3 11 13 0
5 11 2 11 2 2
35 9 9 11 2 0 2 11 2 12 2 12 2 15 13 12 0 9 9 11 11 2 15 13 12 9 7 1 9 1 15 4 3 13 11 2
9 1 9 15 13 1 10 9 2 2
6 3 4 13 0 9 2
12 1 0 9 4 9 13 2 16 15 3 13 2
17 1 0 9 15 9 1 11 13 1 15 7 9 4 15 3 13 2
18 1 0 9 4 3 13 3 2 7 3 15 9 7 7 13 1 9 2
3 9 11 2
22 13 4 2 16 13 1 15 2 7 4 13 7 16 15 15 13 2 3 4 15 13 2
15 7 9 15 3 13 2 3 4 3 13 1 9 2 2 2
26 13 9 2 15 4 1 9 1 0 2 11 13 1 11 7 11 2 3 4 14 13 1 9 1 9 2
16 3 14 2 10 9 15 13 3 2 3 3 13 0 7 0 2
20 9 15 1 15 13 7 15 15 13 2 13 2 14 13 2 13 1 0 9 2
9 3 4 15 13 10 9 9 9 2
11 13 15 9 9 7 15 15 3 15 13 2
17 13 9 2 16 13 1 9 0 2 3 15 13 15 13 2 2 2
19 13 2 16 9 1 11 13 9 7 3 3 4 13 11 15 2 15 3 2
13 3 15 9 3 13 2 1 3 4 13 1 9 2
13 16 9 13 1 9 1 11 2 7 3 13 3 2
3 0 13 11
5 11 2 11 2 2
20 9 11 15 1 9 3 3 13 7 10 9 2 9 11 2 14 10 9 13 2
9 3 15 15 13 13 1 9 0 2
27 3 15 0 9 13 9 0 9 11 1 0 11 2 3 15 13 1 9 9 2 9 7 9 13 1 11 2
14 3 15 9 7 1 9 13 1 0 9 1 9 11 2
13 9 13 1 9 2 16 15 13 13 10 0 9 2
34 1 9 9 13 9 0 9 11 2 7 9 1 0 11 2 9 11 3 0 9 13 11 2 13 15 0 9 11 7 9 11 11 11 2
5 9 1 0 9 2
9 11 1 11 2 9 11 11 2 2
33 13 0 9 10 0 9 13 3 9 11 0 3 0 9 2 1 15 13 9 0 9 1 0 9 2 1 15 15 13 9 0 9 2
21 13 3 0 9 1 3 0 9 1 9 9 7 0 9 1 11 2 12 5 2 2
14 3 12 5 9 11 13 10 9 1 0 9 0 9 2
15 1 9 11 13 3 0 9 9 7 9 0 2 0 9 2
25 0 9 11 13 3 13 2 16 4 15 13 13 0 9 7 1 0 9 7 0 9 1 0 9 2
20 13 2 16 3 3 0 0 9 4 13 0 13 9 1 0 9 9 0 9 2
13 1 9 1 9 11 13 3 0 9 3 3 0 2
6 9 15 2 15 13 3
11 9 0 1 9 1 9 15 13 7 1 11
9 11 2 11 2 11 2 11 2 2
34 1 9 11 0 15 1 0 0 9 11 4 3 1 9 0 9 9 11 13 0 9 2 15 3 13 3 13 1 10 0 9 9 0 2
31 1 9 13 1 9 12 2 10 9 7 4 13 2 7 1 0 9 13 1 0 9 13 3 0 9 1 12 9 0 9 2
7 0 9 13 7 0 9 2
16 0 3 13 13 7 1 9 13 7 16 13 13 12 12 9 2
16 3 1 9 0 9 13 2 16 13 0 3 0 9 1 9 2
10 0 9 9 13 13 9 1 9 9 2
36 9 11 15 13 9 7 13 9 15 0 9 1 0 9 2 13 9 9 0 9 11 11 11 7 13 2 16 9 11 13 3 0 7 0 9 2
23 16 0 9 11 11 13 0 9 7 3 15 13 2 16 15 7 3 13 13 3 16 0 2
12 0 9 13 13 1 11 7 0 9 1 0 2
9 9 1 9 4 13 1 9 9 2
17 0 9 2 7 9 0 1 9 1 0 9 15 13 7 1 11 2
18 16 7 11 13 9 9 11 11 2 9 3 13 3 14 1 12 9 2
5 3 13 1 9 2
21 1 12 9 13 9 9 1 11 2 3 15 12 9 13 0 9 1 9 1 9 2
40 9 15 13 2 7 3 3 13 9 1 9 2 13 11 2 11 7 13 2 16 9 1 9 7 1 9 13 3 3 7 11 2 11 11 2 15 13 1 11 2
17 0 9 0 9 13 7 9 9 11 1 11 2 15 13 1 9 2
18 3 3 13 1 0 9 9 1 9 2 15 13 3 0 9 0 9 2
14 11 12 13 10 9 1 9 9 2 15 7 13 3 2
10 9 11 3 13 1 9 9 1 9 9
7 11 2 11 2 11 2 2
34 9 1 9 9 1 9 9 7 0 9 1 9 13 1 0 9 3 13 1 9 9 7 9 0 9 9 11 2 0 12 9 0 9 2
10 13 15 3 9 9 9 11 2 11 2
10 9 3 9 9 9 13 7 3 13 2
6 15 13 1 0 9 2
35 9 7 1 9 0 9 13 9 3 2 16 13 9 2 16 0 9 9 9 15 13 3 2 15 4 13 2 16 3 13 13 14 1 9 2
14 3 13 1 9 9 0 9 1 0 9 1 0 9 2
19 1 9 9 9 4 9 13 13 9 3 2 16 0 3 1 0 9 13 2
14 0 9 13 9 0 0 9 2 1 15 13 9 13 2
35 10 0 0 9 9 2 3 3 15 13 0 0 9 11 2 13 3 1 9 1 9 2 9 2 0 9 7 3 2 13 9 1 9 11 2
3 9 2 9
18 13 1 9 9 2 9 2 9 7 0 9 2 0 9 2 0 9 2
11 9 7 9 9 2 12 2 9 1 11 2
36 13 2 11 2 9 2 9 2 0 2 2 0 12 2 12 12 11 12 2 9 2 12 2 12 12 12 2 12 2 9 12 2 12 12 12 2
45 9 0 0 9 9 0 2 11 9 2 0 0 9 2 15 13 13 1 9 0 9 1 9 0 0 9 2 3 1 9 0 9 1 9 7 1 15 9 2 3 13 3 0 9 2
19 9 13 9 1 9 9 0 9 0 2 11 9 7 0 9 1 12 9 2
11 9 7 9 9 2 12 2 9 1 11 2
10 13 2 11 2 9 2 9 2 0 2
15 9 9 7 0 9 2 0 9 0 1 9 9 9 9 2
38 10 9 15 13 1 9 7 9 9 11 2 1 10 9 0 9 2 9 7 9 13 1 0 9 7 9 13 13 1 9 9 2 1 9 9 7 9 2
14 9 7 9 9 2 12 2 7 12 2 9 1 11 2
35 13 2 11 2 0 2 9 2 2 11 2 11 2 11 12 2 12 12 11 12 2 9 2 12 2 12 12 12 2 9 12 2 12 12 12
4 3 7 3 2
2 0 9
2 11 11
21 0 2 7 15 0 7 0 9 13 2 3 15 13 9 9 2 1 9 0 0 2
53 9 3 16 13 1 9 9 14 3 1 11 2 9 1 0 9 7 1 9 1 0 9 2 15 13 3 2 7 3 2 9 9 7 9 2 13 1 0 7 0 9 2 1 9 2 16 4 9 12 9 13 13 2
22 13 15 15 3 13 2 9 1 0 7 0 13 0 7 1 0 9 1 15 7 0 2
13 7 2 10 9 15 13 2 13 7 3 3 13 2
17 13 3 0 7 0 2 3 1 9 2 9 1 10 9 1 11 2
30 0 9 13 3 9 2 10 9 15 3 13 2 16 1 9 3 13 2 3 3 3 4 2 9 0 7 0 2 13 2
45 1 0 9 4 1 15 13 0 9 3 15 2 15 3 13 2 3 16 9 2 3 16 9 1 9 2 7 13 4 3 1 0 9 7 13 15 14 1 0 9 2 3 15 13 2
50 1 0 0 2 7 3 14 15 2 9 2 1 9 0 11 7 0 0 9 2 1 9 2 3 15 3 13 13 0 2 0 7 0 9 0 9 2 4 15 13 0 7 9 2 7 9 2 7 9 2
4 14 3 9 2
56 1 9 0 9 2 0 9 1 9 9 11 2 7 0 0 0 9 2 13 13 1 15 0 9 1 0 7 0 9 7 9 2 7 3 15 13 10 0 9 2 0 3 1 10 0 9 2 1 15 15 13 2 3 9 10 2
26 13 4 1 10 9 3 9 9 9 9 2 7 3 3 15 15 13 2 7 13 3 0 0 15 10 2
26 9 9 2 7 15 7 1 9 1 9 2 13 3 1 10 9 7 13 3 1 10 9 7 10 9 2
35 1 0 9 2 13 2 14 1 15 3 3 3 2 13 4 3 2 16 13 3 3 1 9 2 3 1 10 9 2 2 14 3 1 11 2
32 16 15 13 13 15 2 13 9 9 2 2 13 3 2 7 3 13 4 2 9 2 16 9 13 13 0 9 1 9 3 0 2
37 15 4 15 7 13 13 2 13 2 14 15 15 3 3 1 9 0 9 7 0 11 2 13 2 16 13 2 1 9 9 1 9 2 7 10 0 2
12 13 4 15 2 13 3 2 14 0 0 9 2
17 3 2 7 3 4 15 13 2 15 13 2 16 13 1 0 9 2
18 9 0 9 15 13 7 13 15 2 16 3 2 1 0 9 0 9 2
12 3 4 3 13 3 2 15 13 3 3 11 2
8 3 0 1 10 9 0 9 2
4 9 1 0 9
2 11 2
23 9 9 0 9 3 13 1 9 0 9 2 15 9 1 9 13 7 13 1 9 1 9 2
11 13 15 1 0 9 9 9 9 11 11 2
17 9 13 1 11 13 2 16 9 13 9 9 7 9 9 13 3 2
12 1 10 9 9 3 13 9 1 0 9 9 2
38 1 9 9 1 9 1 0 9 2 9 2 2 1 15 9 1 9 13 9 2 15 13 1 0 1 0 9 13 10 0 9 1 12 5 1 12 5 2
5 11 13 1 9 9
2 11 2
17 9 1 9 0 0 9 1 12 9 13 3 0 9 9 11 11 2
13 9 13 13 0 9 1 9 0 9 13 9 12 2
16 4 13 7 9 11 11 2 15 3 13 1 0 9 0 9 2
27 9 9 11 11 13 9 9 9 2 9 7 3 0 9 2 4 2 14 3 13 1 0 9 12 2 9 2
19 1 11 9 1 9 0 9 13 7 0 0 7 0 0 9 1 0 0 2
18 0 9 4 10 9 13 13 3 1 12 9 2 1 0 0 9 9 2
8 3 9 4 13 0 9 9 2
4 0 9 13 9
7 0 9 13 0 0 9 2
4 0 9 15 13
2 11 11
8 1 0 9 13 12 0 9 2
24 10 0 9 13 0 9 9 7 0 9 0 9 2 9 2 0 9 7 1 0 9 0 9 2
11 1 0 0 9 1 11 15 13 12 9 2
15 0 9 13 1 3 12 9 0 9 7 12 9 0 9 2
20 9 13 1 0 9 0 9 9 1 12 9 2 9 13 14 12 9 2 9 2
12 3 16 12 9 9 7 1 9 0 9 13 2
12 1 9 12 7 12 0 0 9 0 9 13 2
20 3 15 1 9 9 9 0 7 0 0 9 11 11 1 10 9 0 9 13 2
5 9 3 1 0 9
9 0 9 13 0 9 9 0 9 2
10 1 10 9 4 13 3 13 3 9 2
33 1 9 1 0 3 0 9 1 0 0 9 1 9 15 3 13 1 9 7 9 0 9 7 0 9 2 7 15 3 1 0 9 2
15 0 9 0 9 1 0 9 13 0 9 7 9 0 9 2
5 9 13 9 9 2
28 9 9 1 10 9 9 13 1 0 12 9 3 0 16 1 9 2 16 9 1 9 13 0 9 1 10 9 2
12 1 9 15 3 13 9 0 9 9 7 9 2
14 1 0 9 13 10 9 10 9 1 9 9 7 9 2
7 0 9 13 9 0 9 2
11 15 9 13 1 9 1 0 9 10 9 2
9 9 13 0 9 1 9 10 9 2
20 9 0 1 0 0 9 4 15 13 3 13 1 9 0 9 1 0 0 9 2
3 9 1 9
7 0 9 13 10 9 9 2
15 3 13 15 9 1 9 1 9 12 7 12 9 1 9 2
19 4 13 1 9 9 0 1 0 9 7 1 9 9 1 9 9 0 9 2
14 3 13 15 0 9 2 9 0 9 2 0 9 3 2
9 0 9 15 13 7 1 9 9 2
10 0 9 13 1 0 12 9 0 9 2
9 3 15 13 7 0 9 10 9 2
31 0 9 0 9 13 3 1 11 2 11 0 0 9 0 3 0 0 9 2 7 16 0 9 15 1 9 1 0 9 13 2
8 11 13 0 9 1 9 0 9
2 11 2
19 0 0 9 1 10 0 9 13 9 0 0 0 9 1 9 0 0 9 2
19 1 11 7 4 13 1 9 9 9 7 9 0 9 13 3 0 9 9 2
12 13 15 3 9 11 1 9 1 9 1 9 2
11 1 0 9 9 11 13 9 11 0 9 2
12 1 10 9 9 0 0 9 3 13 9 9 2
21 11 3 13 9 3 3 7 0 0 9 1 0 9 13 1 12 9 1 12 9 2
20 1 11 4 13 0 9 7 3 13 9 7 13 13 1 9 9 1 0 9 2
30 0 9 13 3 1 10 9 9 3 0 16 11 2 7 15 7 13 1 10 9 1 0 12 1 12 9 1 0 9 2
11 9 1 9 11 7 9 15 7 3 13 2
11 3 0 9 13 12 9 1 9 0 9 2
28 9 13 2 16 9 11 3 13 3 1 10 0 9 2 16 9 15 13 2 16 9 13 3 1 0 9 9 2
13 7 13 11 0 9 9 1 11 0 16 0 9 2
16 11 13 9 0 9 11 1 0 9 1 0 12 1 12 9 2
20 1 0 9 15 13 0 9 9 13 1 12 9 7 1 0 9 1 12 9 2
17 0 9 13 1 0 9 9 1 12 7 1 0 9 1 12 9 2
5 9 1 9 13 3
6 0 11 2 11 2 2
28 16 1 9 1 0 9 13 1 0 9 0 9 0 9 1 12 9 2 1 9 0 11 15 13 1 12 9 2
26 1 9 0 0 9 0 2 11 15 13 13 9 1 9 0 9 2 7 15 7 0 9 9 0 9 2
22 16 13 1 9 9 2 1 0 0 9 13 1 9 7 0 9 2 1 12 9 2 2
23 1 0 9 9 9 2 15 13 9 7 0 9 2 15 3 9 1 9 13 1 12 9 2
4 9 9 3 13
2 11 2
14 0 0 9 9 0 9 15 1 12 2 9 3 13 2
17 13 15 1 0 9 9 0 9 9 0 0 9 1 12 2 9 2
21 1 0 0 9 1 12 2 9 13 1 0 9 1 9 2 7 15 1 12 9 2
17 1 9 1 9 1 9 0 9 3 9 1 10 9 13 12 9 2
21 3 9 0 9 2 9 7 0 9 13 0 7 0 9 13 9 9 7 0 9 2
11 3 1 0 9 13 9 0 7 0 9 2
10 9 9 13 3 0 1 0 9 11 2
34 0 9 9 3 1 0 9 0 1 9 1 9 9 12 13 1 0 9 2 7 15 12 9 2 16 1 11 13 10 9 3 12 9 2
8 0 9 1 0 9 3 13 9
2 11 11
25 13 13 2 16 13 10 0 9 2 13 3 1 9 1 11 7 0 9 0 9 0 9 11 11 2
33 13 2 16 9 9 15 13 3 0 0 9 2 15 4 3 13 16 0 9 7 15 10 9 3 13 0 9 1 0 9 9 9 2
22 1 0 9 2 3 0 9 13 1 9 10 0 0 9 2 13 11 2 11 10 9 2
23 13 2 16 0 9 3 13 2 16 9 1 0 9 13 0 2 15 15 9 9 9 13 2
36 13 4 13 1 15 2 16 9 4 15 13 1 9 2 3 4 13 13 9 1 3 0 9 2 16 15 4 4 13 13 1 0 9 2 13 2
29 11 2 11 3 13 2 16 1 0 9 13 9 0 9 3 1 9 2 7 16 9 9 14 13 0 9 16 0 2
13 0 9 1 0 9 13 13 1 12 9 9 3 2
27 9 10 0 9 3 13 2 16 10 9 13 14 3 0 2 7 13 2 16 11 13 9 7 1 0 9 2
10 10 9 13 7 3 2 16 13 0 2
16 7 15 14 3 2 16 4 10 9 13 3 0 9 2 13 2
28 11 2 11 3 13 2 16 0 0 9 13 9 0 9 2 15 1 10 0 9 13 1 9 1 9 0 9 2
11 0 9 1 15 1 10 9 3 13 13 2
13 9 7 1 10 9 13 9 0 9 1 0 9 2
23 1 9 2 3 13 14 1 9 9 2 11 2 11 13 2 16 7 10 9 13 3 0 2
5 0 9 13 1 9
2 11 11
4 1 9 0 9
18 0 9 15 9 13 1 9 2 3 1 10 0 9 13 13 0 9 2
13 1 0 1 15 13 1 9 9 13 0 0 9 2
22 9 7 13 2 16 9 9 10 9 13 9 7 13 15 2 15 13 1 0 9 9 2
13 9 13 13 0 9 3 7 12 10 9 13 9 2
35 16 13 1 0 9 0 16 12 9 2 13 0 9 14 3 2 13 2 14 1 15 9 7 16 4 0 9 1 0 9 13 7 13 9 2
15 16 9 13 0 9 0 9 2 13 10 9 0 9 9 2
9 9 7 13 7 0 9 0 3 2
46 0 9 13 3 13 2 2 9 9 2 9 2 2 1 15 4 9 13 2 2 9 9 9 2 9 2 9 7 3 0 9 2 2 2 9 9 1 9 2 10 9 13 0 9 2 2
35 10 9 13 0 1 9 9 9 1 9 7 9 9 1 0 9 7 3 3 2 16 4 15 9 13 13 2 16 4 9 13 0 0 9 2
34 9 9 13 4 13 3 2 3 2 9 1 0 9 2 7 3 2 3 2 9 2 9 2 9 3 2 2 2 15 13 1 0 9 2
15 3 0 9 9 9 13 13 9 9 2 3 1 9 9 2
21 3 3 0 9 13 9 1 9 2 7 13 15 9 7 1 9 1 0 0 9 2
18 7 13 0 2 16 4 0 9 13 7 0 9 2 7 0 9 9 2
17 3 4 13 4 9 9 13 3 2 16 15 13 1 0 0 9 2
13 2 9 3 2 9 9 9 7 9 1 0 9 2
1 3
22 0 9 1 11 15 1 9 1 9 3 13 2 1 0 9 7 13 10 9 3 0 2
24 1 0 0 9 0 9 9 13 9 1 0 12 9 9 1 9 1 0 9 3 1 12 9 2
10 0 0 9 15 13 1 9 0 9 2
22 1 0 9 0 9 9 13 1 0 9 2 1 9 0 9 2 1 3 16 12 9 2
8 11 13 0 0 9 1 11 2
15 16 10 9 13 9 0 11 2 0 9 13 3 16 12 2
10 11 13 9 0 9 1 9 9 7 9
2 11 2
27 16 0 9 13 2 16 4 11 13 9 1 11 2 13 4 13 0 9 2 15 3 1 9 1 11 13 2
7 13 15 3 0 9 9 2
48 0 9 9 11 11 2 15 13 1 0 9 1 11 1 9 13 0 9 2 7 13 2 16 0 9 0 1 0 9 9 1 9 1 0 9 11 2 11 2 11 1 9 12 0 9 13 13 2
19 1 0 9 13 0 9 0 9 7 1 9 15 3 9 1 11 1 11 2
16 9 15 1 0 13 9 0 9 7 9 0 9 1 9 9 2
13 11 13 7 13 9 9 0 0 9 1 0 9 2
2 1 9
2 11 2
19 0 9 11 2 11 1 10 0 9 13 0 9 14 1 12 3 0 9 2
33 1 9 9 9 9 9 9 11 11 11 13 1 9 2 15 13 1 0 9 9 1 12 9 1 0 0 9 2 3 13 12 9 2
26 1 9 0 9 2 15 9 3 3 13 9 9 0 0 9 2 3 1 9 1 0 9 13 0 9 2
21 9 13 0 9 2 0 9 1 9 2 3 2 9 2 2 13 0 0 9 3 2
12 3 13 9 9 12 10 0 9 12 9 9 2
28 0 12 9 1 0 0 7 0 9 13 0 9 0 9 11 1 0 9 2 15 13 1 0 9 9 1 9 2
9 4 15 3 13 0 9 0 9 2
2 11 2
19 1 9 0 9 13 0 9 9 12 9 1 9 1 9 0 7 9 9 2
17 1 11 11 1 9 9 9 7 0 9 9 13 1 0 12 9 2
10 9 9 1 0 9 13 7 0 9 2
17 13 15 9 2 3 9 1 9 1 9 9 9 13 3 0 9 2
25 1 9 2 16 13 3 9 2 9 1 9 2 9 7 9 2 13 9 3 0 9 1 0 9 2
5 3 0 9 13 9
12 9 13 9 0 7 0 9 2 13 15 15 13
2 11 11
17 1 0 9 15 10 0 9 13 3 13 2 15 13 7 15 14 2
17 3 13 1 9 0 9 9 7 0 0 9 16 1 12 2 9 2
23 3 3 13 13 1 0 9 9 2 13 11 11 1 0 0 9 11 11 2 0 2 9 2
30 0 0 9 13 3 9 2 15 1 0 0 9 13 7 9 0 7 3 13 3 0 9 7 9 1 9 0 0 9 2
16 1 9 1 9 2 15 13 9 9 2 10 9 1 9 13 2
15 16 11 2 11 13 2 13 15 10 9 13 1 0 9 2
22 1 0 9 13 0 7 1 9 7 0 9 1 9 0 9 9 0 9 1 0 9 2
14 13 3 1 0 9 2 7 13 7 9 1 9 9 2
18 1 0 15 1 9 3 13 2 3 15 13 7 13 3 0 0 9 2
17 3 0 7 0 9 0 9 13 3 9 1 9 2 13 10 9 2
33 13 15 1 9 0 9 7 13 1 15 10 9 13 1 9 2 1 9 7 1 15 7 3 1 15 3 13 2 13 11 2 11 2
30 9 9 1 9 13 7 3 1 3 0 9 2 7 7 7 9 1 9 2 1 15 4 0 9 13 2 3 13 10 2
13 7 15 15 9 13 13 9 0 9 2 3 0 2
33 1 11 2 11 7 9 13 9 7 3 0 9 2 1 10 3 1 9 0 9 13 9 9 1 0 9 7 15 13 0 9 9 2
14 3 0 9 13 1 9 9 1 0 9 0 0 9 2
22 13 3 1 9 0 9 2 9 1 9 2 1 0 9 2 15 13 13 3 2 3 2
12 3 1 15 13 1 9 10 9 0 0 9 2
28 16 15 10 9 13 7 13 2 16 13 0 15 13 2 13 15 9 3 1 9 9 7 1 9 10 0 9 2
17 13 15 3 2 16 4 10 9 13 3 0 2 13 11 2 11 2
15 9 7 0 9 9 13 3 1 9 9 7 0 0 9 2
10 3 0 9 13 7 10 9 7 9 2
18 9 0 9 15 15 3 13 7 13 9 2 3 13 0 9 10 9 2
25 7 3 9 11 2 15 15 13 3 1 9 0 9 2 1 0 9 13 3 0 9 9 7 9 2
17 15 3 13 1 9 16 0 7 10 9 13 1 0 9 0 9 2
31 7 1 15 9 13 1 0 9 11 9 3 0 9 2 1 15 15 13 13 9 0 9 2 9 2 9 9 7 9 3 2
14 0 9 15 3 13 7 1 15 9 0 7 0 9 2
22 1 9 0 0 9 7 9 2 15 1 3 0 9 9 13 2 13 10 9 0 9 2
10 13 1 15 3 7 0 9 0 9 2
15 10 9 10 9 13 9 9 2 3 11 2 11 7 11 2
17 0 9 9 15 1 10 9 7 9 1 0 0 9 13 3 3 2
19 1 0 9 9 1 11 7 9 0 9 1 9 3 13 0 9 0 9 2
23 9 13 2 16 0 9 2 15 13 13 9 1 0 9 2 1 15 13 0 7 0 9 2
15 15 7 13 13 3 14 0 9 2 7 7 9 0 9 2
17 1 10 9 13 0 9 0 9 1 0 9 0 7 3 0 9 2
4 9 9 0 9
25 11 11 1 11 15 13 1 9 13 1 9 9 1 9 2 15 1 12 9 11 13 9 1 9 2
20 1 10 9 4 13 13 9 1 15 1 9 1 9 2 3 0 9 13 9 2
18 9 1 10 9 3 3 13 2 16 3 3 13 1 10 9 1 11 2
17 13 15 14 3 3 1 12 9 2 15 1 10 9 13 0 9 2
6 1 9 15 13 9 2
26 16 15 13 1 0 0 9 2 13 15 1 9 7 9 0 9 1 11 7 3 13 13 1 0 9 2
30 9 1 9 11 15 13 13 1 9 1 11 1 0 0 9 2 15 1 9 9 1 0 9 9 13 9 1 9 9 2
13 3 0 9 13 1 0 9 7 13 9 2 9 2
19 10 9 15 15 13 2 16 13 0 9 1 9 7 15 13 1 15 9 2
18 3 1 9 9 13 1 10 9 1 11 7 13 15 9 2 15 13 2
9 9 13 2 7 13 15 1 9 2
15 1 15 2 15 15 13 2 7 9 9 13 2 13 11 2
15 1 9 2 15 1 9 13 2 13 3 12 12 1 9 2
11 9 0 9 1 9 15 7 13 1 9 2
24 1 9 2 16 0 0 9 13 1 9 1 10 0 9 9 0 9 2 13 1 10 9 9 2
15 10 9 4 13 1 11 2 3 4 13 9 1 0 9 2
11 13 9 7 13 4 15 15 13 2 13 2
27 1 9 2 3 13 10 9 2 1 0 9 13 9 12 12 9 2 2 13 2 16 15 13 0 9 13 2
13 9 9 1 9 13 3 0 1 0 7 0 9 2
17 11 15 3 3 13 2 7 7 10 0 9 13 13 3 0 9 2
18 3 13 14 9 0 9 7 1 9 1 9 15 3 3 13 0 9 2
25 16 15 15 14 13 13 9 1 15 1 0 7 0 9 2 13 1 15 2 16 15 4 13 3 2
13 3 16 15 15 1 10 9 13 7 0 10 9 2
14 15 7 4 1 0 9 13 2 16 13 0 9 9 2
21 1 11 13 7 1 10 9 0 2 16 10 9 13 9 0 9 9 7 0 9 2
15 16 13 2 1 0 9 4 13 1 9 13 1 11 9 2
14 16 13 15 3 3 12 9 2 0 9 1 11 13 2
15 1 0 0 9 1 0 9 13 9 1 9 9 10 9 2
21 15 1 15 1 10 9 1 11 14 13 2 0 3 1 0 9 13 7 10 9 2
20 15 1 15 1 15 13 1 10 9 9 9 2 16 13 2 16 7 3 13 2
16 11 11 13 1 0 9 7 13 2 16 1 15 10 3 13 2
3 2 11 2
5 9 11 11 2 11
3 3 0 11
2 11 2
20 0 9 11 2 11 9 3 13 9 9 0 9 1 12 9 1 12 9 9 2
11 7 3 7 1 10 9 13 0 0 9 2
22 1 0 9 9 11 11 4 13 4 1 15 3 13 9 9 1 9 12 12 0 9 2
17 3 13 2 16 0 9 15 1 0 9 9 13 3 1 9 12 2
34 1 0 12 9 9 11 13 12 12 0 9 2 1 10 12 9 1 11 7 12 9 9 1 0 9 2 15 13 9 0 9 0 11 2
8 11 11 13 0 9 9 11 11
2 11 2
29 11 11 2 11 13 0 13 14 12 9 9 0 9 2 15 4 13 3 1 9 0 0 9 13 0 9 11 11 2
9 13 15 3 0 9 11 11 11 2
26 13 3 2 16 9 0 1 9 9 0 0 9 2 0 1 9 0 0 9 2 13 9 12 9 9 2
16 0 9 11 11 2 11 13 0 0 9 0 7 0 0 9 2
8 10 0 9 13 12 9 9 2
18 1 0 9 13 12 9 2 16 1 9 4 15 13 10 9 3 13 2
5 9 3 4 13 2
23 1 0 9 13 12 5 9 12 0 0 9 2 15 3 12 5 9 13 0 9 11 9 2
12 0 12 5 9 4 13 1 0 9 0 9 2
8 9 9 4 13 1 0 9 2
5 0 9 1 0 9
5 11 2 11 2 2
34 9 9 12 0 2 0 7 0 9 11 2 15 13 13 1 9 9 1 0 9 0 9 1 0 9 7 9 2 13 9 1 0 9 2
8 13 15 0 9 9 11 11 2
14 16 13 2 9 9 13 9 13 9 1 9 0 9 2
13 9 9 13 3 2 9 0 11 2 11 7 11 2
28 9 0 9 1 9 0 1 11 13 12 7 12 9 1 0 9 12 7 12 9 2 16 3 13 14 12 9 2
8 11 11 13 9 1 9 11 11
2 11 2
16 9 11 11 3 13 9 0 9 11 2 11 2 1 0 11 2
23 16 0 9 4 1 0 9 11 11 13 9 12 9 9 9 0 9 1 0 9 12 9 2
23 1 9 0 9 9 2 15 13 9 12 9 9 2 4 13 1 15 13 1 9 0 9 2
21 1 9 0 9 1 9 0 9 2 15 13 12 9 2 13 11 9 3 1 9 2
26 13 3 9 7 9 9 13 9 1 0 0 9 2 15 15 13 2 16 13 1 9 0 9 1 11 2
17 1 9 9 1 0 9 4 13 11 13 3 3 12 9 2 9 2
35 0 9 11 2 15 15 1 11 3 13 1 9 9 2 13 1 10 0 12 0 0 9 1 9 0 0 9 7 1 0 9 1 10 9 2
14 15 13 2 3 3 13 11 2 13 3 0 0 9 2
25 0 9 13 2 16 15 0 9 1 9 3 13 7 1 0 9 13 3 9 0 9 12 9 9 2
8 9 0 9 11 13 3 0 2
22 9 11 11 15 7 13 2 16 1 9 0 9 0 9 13 0 0 9 1 11 13 2
26 3 16 1 11 1 9 9 12 2 12 13 0 13 9 11 0 9 2 3 13 9 7 13 9 9 2
15 1 9 1 0 9 13 1 0 0 11 9 3 0 9 2
5 0 0 9 1 9
15 11 11 13 1 9 0 9 1 9 0 9 1 9 0 9
2 11 2
17 9 0 9 4 1 11 13 0 9 1 9 0 9 1 0 9 2
8 9 13 3 1 12 9 9 2
12 13 15 3 0 9 0 9 11 11 11 11 2
15 10 9 4 11 13 1 9 1 3 0 9 16 0 9 2
23 1 0 9 0 0 9 4 13 9 13 12 9 2 9 0 9 15 4 13 1 12 9 2
13 0 9 0 9 11 11 4 13 13 12 9 9 2
12 10 9 13 11 2 11 3 1 12 9 9 2
24 11 13 3 3 12 9 9 2 1 15 12 7 12 9 13 1 0 9 7 9 13 9 0 2
18 1 0 0 9 0 9 13 11 3 12 9 1 12 9 9 0 9 2
33 12 9 9 9 13 9 2 12 9 9 4 3 13 1 9 11 2 12 9 9 13 9 9 7 0 9 4 13 9 11 7 11 2
13 11 11 13 14 12 9 2 10 9 13 3 13 2
25 0 9 1 11 2 15 13 12 9 2 4 15 13 1 11 2 11 1 9 9 13 1 12 9 2
29 9 9 1 9 1 9 9 13 14 12 9 9 2 12 7 12 9 9 1 10 9 13 9 1 0 9 1 11 2
26 3 12 9 9 13 0 9 2 15 13 0 3 1 0 9 2 9 9 2 0 9 7 0 0 9 2
23 1 11 2 11 11 1 0 9 3 13 1 11 2 3 1 9 0 0 9 1 0 9 2
14 0 0 9 13 3 9 0 0 9 2 11 7 11 2
27 0 9 9 15 13 1 9 12 9 7 13 12 0 9 2 9 9 2 9 0 9 7 9 7 9 9 2
21 0 9 9 9 2 15 11 13 2 13 1 12 2 1 15 13 3 12 9 9 2
4 0 9 3 0
9 1 9 9 13 9 9 0 9 9
2 11 2
14 14 12 12 9 9 13 3 1 9 0 9 0 9 2
19 1 0 9 0 9 11 11 13 13 1 0 9 9 1 12 12 9 9 2
16 1 9 9 9 13 0 9 2 15 13 1 11 7 0 11 2
16 1 0 9 13 9 0 9 12 9 9 2 13 7 1 9 2
10 13 15 9 9 0 9 1 0 9 2
13 3 1 0 9 9 13 0 9 9 12 9 9 2
8 3 9 0 0 9 13 0 2
18 0 9 4 13 1 9 11 16 9 1 9 9 0 9 7 0 9 2
11 12 9 13 3 13 14 12 12 9 9 2
17 0 9 13 7 0 2 1 9 3 3 13 3 12 12 9 9 2
17 0 7 13 12 9 13 7 13 15 0 9 2 3 9 7 9 2
13 1 9 0 0 9 13 1 9 7 1 0 9 2
17 3 12 9 9 9 13 2 1 9 13 0 9 7 9 9 9 2
11 1 9 12 7 12 13 1 11 9 9 2
43 1 0 0 9 2 9 2 9 2 9 2 15 1 0 9 13 3 0 9 11 2 0 9 11 2 0 9 1 0 9 12 5 12 2 0 9 11 7 0 9 1 9 2
24 0 9 2 15 13 1 9 12 0 9 7 13 12 9 2 13 0 9 1 9 12 9 9 2
34 1 0 9 0 9 13 1 12 9 9 0 9 2 12 9 13 9 0 9 2 12 9 13 1 0 9 2 9 13 1 9 0 9 2
5 0 0 9 1 9
2 11 2
23 0 9 0 2 0 2 0 2 0 2 15 13 1 12 9 9 0 9 0 9 11 11 2
29 1 9 11 11 11 11 15 1 9 9 9 1 0 9 13 9 1 9 0 9 7 0 2 0 2 0 2 0 2
11 10 9 13 7 0 0 9 2 9 11 2
19 11 11 2 15 13 0 9 0 0 9 2 13 13 1 0 9 0 9 2
9 1 15 13 13 12 9 9 9 2
23 0 12 9 9 13 0 9 2 12 9 13 0 9 2 9 13 13 1 0 2 0 9 2
16 1 12 2 9 12 2 9 13 9 11 1 9 14 12 9 2
6 9 1 12 9 1 11
5 11 2 11 2 2
24 0 9 9 11 9 9 2 0 9 1 9 12 9 2 13 0 9 9 2 11 11 1 11 2
11 9 11 13 1 9 1 0 9 1 9 2
17 16 4 15 13 13 2 16 13 2 13 15 2 16 13 1 9 2
12 13 2 16 13 9 2 15 4 13 15 9 2
13 11 13 3 2 7 7 15 13 2 16 9 13 2
24 9 1 9 11 15 3 13 13 1 9 11 2 16 4 15 13 13 3 10 12 9 1 9 2
5 9 9 1 9 12
8 9 13 9 9 1 9 0 11
5 11 2 11 2 2
24 0 9 1 11 2 11 2 11 7 11 13 1 9 12 2 9 7 12 2 9 0 9 11 2
12 11 1 15 13 9 10 9 0 9 11 11 2
10 9 0 11 13 0 0 9 0 9 2
62 1 9 12 1 9 0 9 1 10 9 13 9 7 9 2 16 3 2 0 2 0 2 0 2 0 7 0 9 2 9 2 0 7 0 9 2 9 2 9 2 0 7 0 9 2 0 9 2 9 7 9 2 0 9 2 0 9 2 0 9 3 2
37 1 0 9 15 13 3 9 2 9 2 9 2 9 2 0 9 2 9 2 0 9 2 9 2 0 9 2 0 9 2 0 9 2 9 7 0 2
27 9 0 11 13 1 11 2 11 0 13 10 0 7 0 9 1 0 9 2 10 9 7 0 9 13 3 2
28 3 15 13 13 15 2 16 4 15 9 1 10 9 13 1 10 0 9 2 9 13 1 11 2 11 1 9 2
19 1 0 9 15 13 7 0 9 0 9 2 0 9 7 9 1 0 9 2
20 9 9 9 1 9 1 9 2 15 13 9 0 9 11 2 13 12 2 9 2
10 1 9 4 13 12 9 1 0 9 2
24 3 4 15 13 2 16 0 9 0 9 13 13 2 13 9 9 1 12 9 9 2 11 11 2
5 9 11 11 2 11
6 0 11 13 9 1 9
2 11 2
21 0 7 0 9 0 0 9 2 11 2 13 1 9 1 9 1 0 11 1 9 2
23 9 0 0 9 1 0 11 13 1 9 2 3 13 9 11 9 1 9 9 2 1 9 2
13 1 0 9 13 1 9 9 9 9 1 0 9 2
17 1 9 0 0 9 1 0 0 11 13 0 9 9 1 0 9 2
4 3 1 9 12
10 13 0 2 16 4 0 9 13 10 9
16 9 11 11 13 1 0 9 1 0 9 9 0 9 11 11 2
19 13 15 2 16 15 15 13 13 0 9 1 9 13 0 9 1 0 9 2
19 1 15 13 13 3 3 2 16 13 3 1 0 9 9 7 9 10 9 2
33 13 15 3 7 9 0 2 0 7 15 13 9 2 16 0 9 13 13 1 15 0 7 16 0 9 13 13 1 3 1 9 0 2
37 7 10 9 13 0 2 13 2 16 13 1 12 1 0 9 10 9 2 7 7 4 15 13 3 13 9 7 13 15 1 10 0 9 1 0 9 2
21 13 2 16 3 2 1 0 9 2 4 15 13 2 13 2 7 15 13 0 2 2
20 13 11 16 0 9 1 0 9 0 9 2 15 4 3 13 10 9 1 9 2
17 13 15 1 10 9 1 9 2 15 3 13 1 11 7 9 11 2
7 11 3 13 10 10 9 2
18 15 4 15 13 15 2 16 13 0 2 16 4 0 9 13 10 9 2
5 1 15 15 13 2
4 9 13 12 2
60 1 9 1 9 7 9 13 1 10 9 10 9 7 10 9 2 16 13 0 9 15 1 10 9 13 1 10 0 9 2 7 7 13 12 9 10 7 15 9 4 13 1 10 9 3 0 7 13 2 16 1 15 15 13 7 1 0 0 9 2
7 0 9 13 1 0 9 2
25 13 0 9 1 0 9 2 3 9 15 12 0 13 3 3 0 2 7 3 1 9 15 9 13 2
46 13 3 13 3 0 9 1 9 0 9 2 7 7 3 15 15 15 13 3 0 2 16 0 15 13 13 0 9 7 13 15 13 2 16 4 13 1 0 11 2 11 2 11 7 11 2
6 7 10 9 13 2 2
14 13 3 9 2 16 15 11 13 13 9 1 9 11 2
35 3 4 15 13 2 16 16 4 13 1 0 9 9 13 9 2 1 15 4 15 13 2 16 13 3 10 9 0 2 7 4 15 13 11 2
19 16 9 2 16 4 13 9 2 16 4 15 15 13 2 13 1 3 0 2
16 1 15 4 3 13 2 10 0 9 11 15 10 9 13 2 2
11 10 13 9 1 9 0 9 1 0 9 2
35 11 3 13 9 2 15 13 3 7 9 10 2 16 0 9 10 0 9 13 0 9 2 7 16 9 13 0 9 15 0 13 3 3 9 2
28 9 13 10 2 0 15 2 16 1 9 0 9 13 9 14 0 9 2 7 7 0 9 2 15 13 10 9 2
6 13 0 0 0 9 2
20 13 9 10 9 7 13 3 0 2 3 3 0 9 9 2 1 15 15 13 2
10 4 15 13 2 13 10 9 3 13 2
23 15 13 10 0 9 2 7 7 3 4 13 0 9 16 0 9 0 9 1 0 0 9 2
25 1 0 9 13 2 16 1 9 0 9 13 0 0 9 2 9 13 0 9 13 7 13 10 9 2
11 15 13 2 16 4 13 1 9 0 9 2
10 1 9 0 9 13 9 1 15 13 2
31 9 11 1 9 9 9 1 9 9 9 9 1 11 3 13 9 11 11 3 0 9 0 9 11 11 1 9 14 1 9 2
8 12 7 10 9 13 1 9 2
5 9 11 11 2 11
3 9 1 11
7 11 2 11 2 11 2 2
14 9 0 11 11 11 3 13 9 9 7 13 1 9 2
10 3 13 9 10 9 7 9 0 9 2
10 11 1 9 13 0 9 9 11 11 2
25 1 11 13 11 2 15 1 11 13 0 9 1 11 2 11 2 0 1 9 11 7 3 3 0 2
8 11 15 1 0 9 13 13 2
41 11 2 11 3 11 13 2 16 9 0 2 9 2 11 2 15 13 0 9 0 7 0 9 2 11 2 7 13 11 2 13 9 1 10 9 9 1 0 9 9 2
24 9 13 1 9 10 0 9 1 0 9 9 0 2 0 9 2 15 9 11 13 2 13 11 2
18 13 13 2 16 1 9 9 13 1 0 9 0 9 11 11 2 11 2
20 13 13 1 9 1 0 9 11 2 16 1 10 9 11 3 13 2 13 11 2
16 13 2 16 0 9 1 11 15 13 1 0 9 11 2 13 2
7 11 0 9 13 1 9 2
19 9 11 13 16 9 9 13 9 1 9 9 7 13 15 3 3 0 9 2
16 13 15 9 11 11 2 11 1 15 2 16 11 13 0 9 2
15 1 9 11 7 9 11 9 11 13 3 1 12 12 9 2
38 1 9 11 2 15 1 9 11 13 9 2 9 9 11 13 2 16 1 0 9 13 3 2 9 9 9 11 11 2 11 7 9 9 9 11 2 11 2
7 1 11 13 0 9 9 2
5 9 13 9 9 9
11 1 9 9 4 9 11 13 1 9 1 9
5 11 2 11 2 2
11 9 9 1 0 9 13 3 9 9 9 2
16 1 10 0 9 1 9 9 11 11 15 13 9 9 11 11 2
18 9 11 15 1 9 13 10 9 9 9 2 15 13 9 9 13 3 2
12 11 2 11 3 13 2 16 13 12 9 9 2
39 16 3 13 11 2 9 3 13 7 1 9 9 9 7 9 0 2 0 2 0 2 2 15 0 9 1 0 9 9 13 2 1 9 0 9 0 9 11 2
21 1 15 13 9 12 0 9 9 1 9 2 15 3 9 0 16 0 0 9 13 2
10 1 9 15 13 3 3 2 13 11 2
25 1 10 9 13 9 9 13 2 16 10 9 0 9 13 0 7 1 9 1 15 13 13 3 9 2
17 9 0 2 0 2 0 2 13 1 15 2 16 9 11 13 0 2
12 3 15 13 11 11 1 0 2 0 2 0 2
26 13 3 2 16 9 13 0 9 2 15 1 15 13 0 0 0 0 0 9 1 0 9 12 9 9 2
7 0 9 13 1 11 1 11
2 11 2
25 12 12 9 2 15 13 9 9 9 1 0 9 2 13 1 0 9 1 9 1 9 1 9 11 2
14 13 1 15 3 0 9 0 9 0 9 11 11 11 2
10 13 2 16 3 13 10 9 12 0 2
15 0 9 7 13 14 3 1 9 2 3 4 13 12 0 2
7 0 12 4 13 9 9 2
12 0 9 0 9 13 1 15 13 3 0 9 2
5 9 9 13 1 9
2 11 2
35 9 0 9 9 11 11 13 13 1 0 9 9 2 15 15 13 13 15 2 16 1 0 9 13 1 9 12 0 9 3 1 12 9 9 2
7 3 1 15 13 9 11 2
15 1 9 13 0 9 2 16 11 13 2 16 9 13 0 2
5 9 13 7 1 9
12 9 9 0 9 11 13 9 1 0 9 9 11
2 11 11
15 9 9 13 1 0 7 1 15 2 10 9 13 1 9 2
23 0 0 9 15 1 10 9 3 3 13 2 16 9 0 1 9 0 9 15 15 3 13 2
21 12 1 9 2 3 13 13 0 9 1 0 9 7 1 9 2 13 0 9 11 2
16 1 9 2 15 13 9 9 2 13 11 1 10 9 11 11 2
12 10 9 13 2 16 4 9 13 1 15 3 2
23 7 15 13 9 1 0 0 7 0 9 7 13 1 15 9 7 1 11 2 7 1 9 2
8 13 15 0 9 9 2 13 2
14 3 0 15 13 0 9 2 15 0 9 3 14 13 2
23 13 15 9 9 1 0 9 0 2 11 2 0 0 11 2 2 15 13 9 11 1 11 2
18 10 9 13 13 3 0 7 0 9 1 9 0 9 1 12 9 9 2
18 0 9 1 9 15 13 9 9 2 15 13 1 9 7 9 0 9 2
24 9 1 9 13 0 2 9 1 9 13 0 7 9 1 9 13 13 3 0 9 1 9 9 2
17 0 2 11 13 0 9 2 9 15 13 13 14 1 12 9 9 2
42 1 9 1 0 9 13 9 9 0 9 1 0 9 2 15 13 9 0 1 10 9 1 0 7 0 9 2 0 9 2 0 9 7 9 9 2 9 9 0 2 2 2
8 10 9 15 13 1 0 9 2
6 1 15 13 9 3 2
21 0 9 13 0 9 2 0 1 9 9 7 9 2 15 1 9 13 1 0 9 2
14 13 13 0 9 0 9 7 3 3 0 9 10 9 2
19 0 9 7 9 1 0 9 13 3 0 9 0 9 9 7 0 9 11 2
3 0 9 9
14 0 11 2 9 7 10 9 13 10 9 1 0 9 2
7 0 9 13 9 1 9 2
10 9 7 9 13 1 9 7 0 9 2
29 0 9 2 15 13 15 13 0 9 2 13 13 0 2 11 2 9 0 13 0 9 1 0 7 0 9 1 9 2
18 9 0 9 4 1 9 2 9 7 9 1 9 13 3 1 12 9 2
18 9 2 15 3 0 9 13 2 4 15 13 13 10 9 2 0 9 2
15 13 15 13 1 9 0 0 9 11 2 11 0 1 9 2
19 1 9 9 13 1 9 9 1 3 16 12 9 9 1 3 16 12 9 2
19 9 7 13 1 0 9 13 0 9 2 15 15 13 13 9 9 1 9 2
10 11 2 11 13 7 1 0 9 9 2
19 3 13 13 0 9 0 9 11 2 15 13 9 0 9 0 9 1 9 2
15 10 9 15 13 1 9 2 1 9 11 7 1 0 11 2
6 0 9 1 9 3 13
2 11 2
30 9 13 4 1 9 13 9 11 1 11 2 15 4 1 0 9 13 9 2 16 13 9 1 9 0 2 3 0 9 2
27 0 0 9 9 9 2 15 4 13 3 1 9 2 13 1 15 2 16 13 1 9 3 0 9 1 9 2
26 9 11 11 1 15 3 13 2 16 3 15 0 9 13 7 3 0 9 9 13 1 9 9 0 9 2
33 1 9 15 3 2 13 2 16 1 12 2 9 0 9 13 4 3 0 9 13 9 1 9 12 9 7 0 9 1 9 12 9 2
6 9 1 9 13 1 9
2 11 2
18 1 0 9 1 11 1 11 4 3 1 9 0 9 13 12 0 9 2
5 13 15 9 11 2
24 9 13 3 15 2 16 9 0 9 13 1 9 11 9 1 9 9 12 9 3 1 0 9 2
8 9 15 13 3 3 0 9 2
16 1 0 9 13 0 2 16 4 9 1 9 13 14 12 9 2
25 1 9 9 9 11 11 4 9 13 1 9 13 9 1 0 9 7 0 9 13 2 3 7 3 2
18 9 9 9 9 1 9 13 1 9 0 9 2 15 4 13 4 13 2
11 9 1 9 1 9 4 13 3 12 9 2
4 9 13 4 13
5 11 2 11 2 2
18 9 13 1 12 2 9 9 0 0 9 0 9 7 10 0 0 9 2
23 9 9 2 15 15 3 13 13 2 13 3 0 9 1 9 0 9 1 0 9 7 9 2
34 1 9 4 15 13 3 13 0 0 9 2 9 2 1 9 0 1 9 1 9 1 12 9 0 9 1 12 9 1 9 12 9 3 2
17 0 9 4 13 4 13 1 9 12 9 3 2 3 12 9 2 2
15 3 13 1 9 9 10 9 13 9 2 15 13 12 9 2
10 9 4 13 13 1 12 1 12 9 2
30 1 9 13 9 9 9 9 2 16 4 1 9 1 9 9 7 0 9 13 1 9 9 9 0 9 9 9 0 9 2
21 9 3 13 9 1 9 3 9 1 9 0 9 7 9 0 1 9 12 7 12 2
31 4 13 2 16 4 15 0 2 0 2 3 0 2 1 9 9 2 0 7 0 9 13 1 12 9 7 0 9 12 9 2
13 3 1 10 9 4 13 13 0 0 9 0 9 2
23 10 9 7 4 13 1 9 2 13 15 10 9 2 16 15 1 3 3 0 12 9 13 2
14 0 9 4 13 0 9 9 13 1 10 9 0 9 2
10 0 9 1 11 13 13 9 1 0 9
5 11 2 11 2 2
24 1 0 0 9 11 4 3 13 12 1 0 7 0 9 0 7 0 9 1 0 7 0 11 2
26 13 15 9 1 0 9 2 11 9 2 9 2 0 2 2 2 15 13 0 9 0 2 0 11 11 2
16 0 9 1 15 13 11 1 11 2 1 10 9 4 9 13 2
10 9 13 1 9 9 7 9 0 9 2
8 11 13 1 9 9 1 9 2
12 9 9 13 13 9 1 9 0 9 10 9 2
39 13 3 1 0 9 0 1 0 0 9 2 15 4 13 13 9 1 0 9 7 3 9 1 9 10 3 0 9 2 13 3 1 0 9 9 9 11 11 2
11 0 9 3 0 9 13 12 9 0 9 2
25 9 3 4 13 1 9 9 0 11 7 11 2 1 9 11 2 11 2 9 7 1 10 9 11 2
5 9 9 15 13 9
5 11 2 11 2 2
22 1 9 2 7 3 1 0 0 9 13 3 3 0 9 9 0 9 16 1 12 9 2
6 3 15 13 9 9 2
22 13 15 1 9 9 9 2 15 15 13 9 2 1 15 1 10 9 13 1 9 12 2
22 9 3 13 12 9 0 9 1 0 12 7 0 0 9 13 9 9 1 3 16 9 2
11 0 9 1 9 9 0 9 13 0 9 2
16 12 9 0 9 13 1 0 9 2 12 7 9 9 1 0 2
17 1 0 0 9 13 0 0 9 3 12 9 2 1 9 12 9 2
31 1 9 9 15 3 13 9 1 9 0 0 9 2 7 13 13 15 16 0 9 2 1 15 15 9 1 0 9 13 9 2
26 9 9 13 13 7 3 13 9 1 9 0 9 7 3 13 1 0 9 2 3 4 9 4 3 13 2
11 1 0 0 9 13 9 13 10 0 9 2
18 13 15 2 16 12 1 9 13 9 9 9 7 0 9 1 9 9 2
32 9 13 7 7 13 0 9 9 2 7 2 3 13 9 9 11 11 2 7 1 9 9 13 0 3 0 9 9 16 15 0 2
12 9 9 7 13 1 3 0 9 9 1 9 2
9 3 3 13 10 9 1 9 9 2
7 9 9 2 15 13 1 9
8 11 11 2 9 9 2 9 11
30 0 9 13 9 9 11 2 7 7 15 0 9 1 10 9 13 9 9 2 15 1 0 0 9 11 13 13 0 9 2
17 11 13 9 9 2 1 15 15 13 3 2 7 14 3 7 3 2
9 9 11 2 13 1 9 1 9 2
8 13 16 9 7 9 15 13 2
11 1 9 13 1 0 9 0 12 12 9 2
12 1 9 13 10 9 3 3 3 2 1 9 2
12 0 9 1 9 15 1 15 13 9 0 9 2
7 13 4 3 1 0 9 2
12 13 4 1 9 2 13 13 2 13 4 9 2
13 9 1 0 9 2 9 7 9 13 1 15 15 2
8 14 3 0 9 0 0 9 2
10 7 13 9 2 15 13 9 0 9 2
5 13 13 1 9 2
2 3 2
8 3 3 3 16 3 2 2 2
9 9 11 2 13 0 9 10 9 2
8 1 9 9 15 13 3 9 2
14 13 1 9 1 9 1 0 2 13 15 7 13 9 2
13 3 1 9 1 9 1 15 13 0 9 0 9 2
7 13 15 3 13 3 15 2
8 1 10 9 15 10 9 13 2
16 0 9 15 13 3 0 9 7 3 15 13 3 9 0 9 2
10 3 2 1 9 2 15 9 13 15 2
20 9 11 2 15 3 13 1 0 9 2 1 15 15 10 0 9 13 0 9 2
13 9 9 11 2 13 1 9 11 3 3 1 12 2
28 16 9 2 15 13 9 1 0 9 9 9 2 13 13 9 2 11 11 1 9 0 7 0 9 11 1 11 2
8 9 1 15 13 0 9 3 2
10 11 11 13 0 9 1 9 9 0 11
5 11 2 11 2 2
29 16 13 1 9 1 0 9 0 11 2 13 9 9 11 11 1 0 9 11 9 1 9 2 15 4 13 9 13 2
20 11 15 3 13 0 9 11 1 11 11 11 2 15 10 9 13 16 0 13 2
32 9 0 9 9 0 11 2 15 13 13 1 9 1 0 9 2 13 3 7 1 9 9 9 0 9 0 1 12 0 9 11 2
19 1 9 11 13 3 3 9 9 2 1 15 4 13 10 9 1 0 9 2
22 1 9 9 15 7 13 13 9 1 9 9 11 11 7 10 9 11 11 1 9 11 2
17 0 9 13 13 9 3 3 0 9 9 2 15 13 12 2 9 2
21 10 9 4 3 13 1 9 1 9 9 2 1 0 9 13 1 9 0 0 9 2
9 15 7 10 9 9 13 1 0 2
27 11 2 11 13 9 2 16 1 9 9 13 13 1 9 2 15 4 13 9 12 7 0 9 1 0 9 2
14 1 10 9 4 13 11 2 11 13 9 0 9 11 2
8 11 13 9 9 1 0 9 9
5 11 2 11 2 2
18 0 0 9 3 13 9 1 9 9 2 15 13 1 10 0 9 9 2
21 1 10 9 11 11 13 10 0 9 11 0 9 9 9 1 0 0 9 7 9 2
24 9 1 9 13 1 9 2 16 15 9 1 9 13 1 9 3 2 16 15 13 1 9 9 2
26 16 1 10 9 3 3 1 9 11 11 11 13 9 11 2 13 4 15 3 13 1 9 11 15 9 2
32 0 9 13 7 11 2 11 1 3 0 2 3 13 13 9 1 11 7 9 2 14 13 14 1 10 9 2 7 13 13 9 2
27 3 13 1 11 0 13 9 2 16 9 9 4 13 1 15 2 16 4 15 1 15 0 9 13 9 13 2
19 1 9 1 11 13 12 0 9 1 0 9 0 9 2 0 7 0 9 2
16 14 1 10 9 4 0 9 13 9 11 7 13 1 9 11 2
15 15 0 9 4 3 1 11 13 9 3 1 9 1 9 2
3 9 1 11
2 11 2
30 0 0 9 11 2 12 2 0 1 9 0 9 1 9 7 9 0 9 1 0 9 2 15 13 1 9 9 1 11 2
12 9 9 1 0 9 13 0 0 9 11 11 2
28 11 2 15 13 1 9 0 9 11 1 9 0 9 1 0 9 2 15 13 1 9 12 3 1 10 0 9 2
8 0 9 3 13 9 0 9 2
35 0 9 0 9 15 13 9 1 0 2 0 2 0 2 0 2 0 2 0 2 0 2 0 2 0 7 0 9 7 3 3 2 9 9 2
18 9 7 9 15 13 11 13 16 0 9 7 15 13 1 9 0 9 2
13 9 15 13 13 1 9 11 11 1 12 2 9 2
4 9 9 0 9
23 0 9 2 1 0 9 2 9 12 2 9 2 13 0 9 10 9 0 0 9 0 9 2
24 1 10 9 13 1 0 0 9 0 9 2 15 3 13 1 0 9 0 2 0 0 9 11 2
27 13 15 15 10 9 1 0 9 13 1 0 9 9 0 9 2 15 4 13 1 0 12 9 1 12 9 2
30 13 2 16 10 9 13 1 9 2 7 13 13 10 9 7 9 13 1 10 0 9 2 9 2 12 2 12 12 12 2
22 13 2 14 9 1 10 9 2 13 15 15 9 1 0 9 2 16 4 13 13 9 2
9 11 2 11 2 9 11 13 0 9
7 11 2 11 2 11 2 2
26 1 0 9 1 9 13 3 9 10 0 9 11 11 2 11 2 9 11 13 3 0 0 9 0 9 2
12 16 3 13 11 2 13 1 0 2 0 9 2
11 13 15 7 9 2 7 13 9 1 9 2
19 11 1 9 13 2 16 13 3 2 3 15 13 13 1 9 1 0 9 2
23 13 9 2 16 9 1 0 9 1 15 13 9 2 7 4 15 13 13 1 9 7 9 2
10 13 4 15 13 0 9 7 10 9 2
7 0 9 3 9 0 9 13
5 11 2 11 2 2
21 0 9 3 13 0 9 2 15 13 9 9 0 9 7 14 9 1 9 0 9 2
15 3 7 13 1 0 10 9 1 0 9 2 3 13 11 2
17 3 0 0 9 4 15 9 3 13 2 13 3 9 11 11 11 2
18 0 9 11 11 13 9 11 1 0 9 2 15 13 0 9 1 9 2
11 1 15 13 1 10 9 9 3 9 13 2
17 9 3 0 0 9 7 9 1 9 9 13 1 9 1 0 9 2
23 9 0 0 9 2 11 2 11 2 15 13 9 11 1 0 0 9 13 1 9 9 9 2
22 9 11 2 11 11 11 3 13 2 16 13 0 13 9 11 1 0 9 1 10 9 2
27 9 15 1 10 9 10 9 13 2 7 2 3 13 2 15 13 13 2 16 4 1 9 1 10 9 13 2
11 9 11 11 11 7 11 11 13 1 0 9
5 9 11 11 2 11
6 1 0 9 13 10 9
3 1 0 9
7 11 2 11 2 11 2 2
12 3 12 12 9 11 1 0 0 9 13 9 2
9 13 15 3 0 9 9 11 11 2
13 9 0 9 1 9 11 1 15 13 1 9 9 2
29 1 9 2 16 15 11 13 0 9 1 9 2 13 0 9 11 2 11 2 16 9 1 0 7 0 9 15 13 2
34 13 7 2 16 1 9 0 0 9 4 15 15 12 0 9 2 15 15 9 13 2 13 13 1 15 2 15 13 0 9 1 0 9 2
18 0 9 4 1 15 13 9 1 0 9 2 15 4 15 11 13 13 2
35 1 9 9 12 5 12 5 12 13 0 0 9 1 0 11 13 11 11 2 16 15 13 1 0 9 2 15 13 4 3 3 13 9 9 2
5 11 4 13 9 9
3 1 0 9
2 11 2
26 9 11 13 9 9 9 2 16 4 13 2 16 0 9 2 15 13 10 9 1 9 11 2 13 9 2
12 1 0 0 9 11 15 13 9 9 11 11 2
33 0 9 11 11 11 1 15 13 2 16 10 9 0 0 9 0 7 0 9 13 1 11 9 1 0 7 0 9 1 10 0 9 2
12 13 2 16 13 3 3 1 9 9 11 11 2
38 9 0 9 1 10 9 13 9 2 15 9 13 13 10 9 3 1 9 2 7 1 11 15 4 2 3 13 11 2 13 9 2 15 0 9 3 13 2
8 9 13 9 9 7 1 0 9
3 1 0 9
2 11 2
46 9 7 9 1 11 2 11 13 1 9 0 9 1 0 9 9 9 9 2 16 4 12 9 1 9 1 9 1 0 9 2 0 1 0 9 2 0 9 3 2 2 13 1 0 9 2
8 13 15 3 9 9 11 11 2
25 11 2 11 13 1 15 1 15 2 16 4 9 9 0 9 4 16 3 13 1 9 9 7 9 2
15 1 9 13 0 3 13 9 1 9 0 9 7 0 9 2
27 9 1 10 9 7 9 4 13 13 13 7 13 4 15 13 9 9 1 9 9 1 0 9 2 13 11 2
6 11 2 11 1 0 9
5 11 2 11 2 2
22 9 0 9 1 11 13 1 9 9 1 0 9 11 11 7 10 9 2 0 11 11 2
9 3 3 4 13 1 0 0 9 2
21 16 4 3 13 1 11 2 12 9 13 1 9 0 9 1 0 9 1 0 9 2
26 11 11 2 11 11 7 11 11 4 13 1 0 9 9 2 15 15 13 13 1 9 7 9 10 9 2
15 1 9 9 9 15 13 9 9 9 1 12 1 12 9 2
5 0 9 1 0 9
2 11 2
44 1 9 9 0 9 11 2 0 1 9 0 2 0 7 0 0 9 2 15 1 9 12 2 2 12 2 9 13 1 11 9 1 9 9 0 9 0 9 7 9 2 9 2 2
25 9 0 4 13 3 0 0 9 2 10 9 7 3 9 10 0 9 1 0 2 0 7 0 11 2
14 1 11 15 9 13 1 3 0 9 16 1 0 9 2
14 7 3 13 0 9 10 9 1 9 7 1 0 9 2
8 1 0 9 1 9 14 1 9
5 11 2 11 2 2
21 1 9 3 16 12 9 9 15 1 0 9 1 11 13 0 9 9 2 11 11 2
23 16 13 13 1 9 2 13 1 9 9 7 1 9 9 2 3 7 1 9 0 0 9 2
11 1 9 15 1 11 13 1 9 2 12 2
7 13 15 9 0 9 11 2
7 3 15 13 1 0 9 2
5 13 15 0 9 2
6 13 13 0 9 9 2
8 3 13 1 9 3 13 9 2
15 9 2 15 13 3 13 1 9 2 15 7 13 1 9 2
27 1 9 0 9 2 11 2 11 13 9 2 0 15 0 9 3 16 12 7 12 9 9 2 1 0 9 2
13 1 9 2 3 1 9 13 2 13 9 0 9 2
11 3 4 13 14 1 12 2 12 2 12 2
18 1 10 9 4 13 16 9 7 1 15 13 11 11 2 9 3 13 2
16 0 13 2 16 15 13 0 2 16 4 15 13 0 9 9 2
16 13 2 16 13 1 10 9 1 9 2 7 3 9 0 9 2
11 9 13 3 0 9 1 9 9 1 9 2
10 15 1 15 13 0 9 7 13 15 2
13 1 0 9 4 15 13 1 3 15 0 9 13 2
29 7 0 9 2 1 15 4 13 13 2 7 0 9 15 9 13 13 2 16 13 9 2 16 15 13 1 10 9 2
14 11 1 15 3 13 13 7 9 1 0 9 1 9 2
8 13 15 9 2 13 11 11 2
9 0 9 13 1 0 9 0 9 2
8 0 9 1 9 1 11 2 11
2 0 9
5 11 2 11 2 2
26 9 13 1 9 0 9 1 0 9 2 13 11 9 9 0 9 1 11 11 11 1 9 10 0 9 2
32 10 9 13 1 0 9 9 0 9 1 11 1 11 11 2 15 4 13 1 9 12 1 0 9 0 9 1 12 9 9 9 2
19 9 13 2 16 1 9 12 7 12 13 0 9 1 0 0 9 0 11 2
24 9 9 11 2 11 13 2 16 9 1 11 2 11 4 13 2 16 13 1 9 9 0 9 2
15 9 4 13 1 12 1 12 9 0 9 9 12 0 9 2
26 1 9 9 13 13 2 0 9 9 2 15 9 13 2 3 9 9 2 3 9 7 9 10 0 9 2
19 0 9 13 2 16 15 9 13 1 15 0 9 7 9 1 9 0 9 2
7 9 11 13 1 9 12 2
15 0 15 13 2 7 13 1 15 2 16 9 13 3 13 2
35 9 9 0 0 9 11 11 2 15 9 1 11 11 13 2 13 1 9 11 9 1 9 2 16 0 0 9 13 1 9 0 9 3 13 2
5 1 15 13 13 2
8 10 9 4 13 1 9 9 2
29 16 4 0 9 1 11 13 9 2 16 0 0 9 13 13 2 13 4 0 9 2 15 15 13 2 13 11 11 2
1 9
20 1 9 11 13 3 3 0 0 9 1 11 9 1 12 9 2 15 3 13 2
19 9 13 2 16 3 1 12 9 13 9 1 9 7 9 9 0 1 9 2
3 1 9 9
1 9
2 11 11
24 0 9 13 11 3 0 9 1 15 9 1 3 0 9 1 9 0 9 9 0 0 9 9 2
28 0 9 13 9 1 9 12 9 11 2 15 11 0 0 9 13 1 12 9 11 2 3 12 9 0 9 2 2
17 10 9 13 1 9 0 0 9 2 11 2 0 9 1 0 9 2
21 1 9 13 0 9 0 9 9 3 1 0 9 12 12 11 2 7 4 3 13 2
18 9 0 9 1 12 9 3 1 0 9 13 0 9 1 9 1 9 2
12 3 0 9 13 1 0 9 3 1 9 9 2
14 13 15 3 2 16 0 9 1 9 0 9 13 0 2
43 16 1 9 12 13 0 9 1 12 5 7 9 0 9 13 11 10 9 1 0 11 1 0 12 9 2 13 0 9 13 1 9 7 1 9 1 0 9 3 12 9 9 2
16 3 1 9 13 11 0 0 9 7 13 0 9 1 9 9 2
23 16 9 9 13 13 16 0 9 2 13 9 9 0 9 9 2 15 0 9 13 3 13 2
22 11 3 13 0 0 9 7 9 1 0 9 2 15 3 7 1 0 9 13 0 9 2
23 3 13 3 0 2 16 9 1 0 9 9 13 1 9 7 0 2 0 9 4 3 13 2
17 1 11 13 1 0 9 0 3 9 1 11 1 9 9 7 9 2
18 0 9 9 0 9 0 9 13 15 0 2 16 0 9 9 3 13 2
13 0 0 9 9 12 9 11 7 3 0 9 13 2
9 0 9 0 9 4 7 3 13 2
29 1 0 9 13 3 0 2 0 9 9 1 0 9 12 2 12 7 13 15 1 0 9 2 15 9 13 1 9 2
12 1 9 9 4 13 13 9 9 11 7 11 2
8 10 9 15 3 13 0 9 2
20 16 15 3 13 3 2 0 9 0 9 7 9 0 9 13 13 3 0 9 2
25 0 9 1 11 2 7 1 9 1 9 0 9 9 2 1 0 9 0 9 1 9 9 3 13 2
10 1 15 13 1 0 9 3 15 13 2
32 1 0 9 9 0 0 9 1 11 13 0 13 3 1 9 0 9 2 15 13 0 9 1 0 9 2 11 2 7 0 9 2
5 9 0 9 13 9
8 11 11 2 9 11 7 9 9
18 1 0 2 0 9 0 9 13 3 0 0 9 1 9 7 0 9 2
23 9 4 13 13 0 9 2 10 9 13 9 2 16 3 9 13 2 7 3 9 4 13 2
17 0 9 0 9 1 9 13 3 1 9 13 9 9 7 0 9 2
22 13 1 0 9 2 1 15 4 13 0 13 3 2 7 1 9 9 9 9 9 0 2
22 13 3 0 9 1 9 9 1 0 9 2 15 2 15 9 13 13 3 2 13 9 2
6 9 7 3 13 9 2
19 9 13 3 0 9 7 0 9 2 15 13 10 9 13 0 9 7 9 2
26 3 7 9 13 13 0 9 2 0 1 15 9 7 0 13 7 1 9 0 9 2 1 9 3 0 2
21 7 3 9 0 7 0 9 10 9 2 15 13 0 9 9 7 0 9 1 9 2
26 0 2 7 16 3 0 9 0 9 1 9 15 13 3 1 0 9 2 3 3 0 9 15 1 9 2
40 9 13 15 3 1 9 0 9 2 13 0 10 3 0 9 2 9 0 1 9 2 9 2 3 9 4 13 9 2 13 3 0 7 13 0 0 7 0 9 2
26 1 9 0 9 0 9 2 10 2 15 13 0 7 1 9 3 3 7 0 9 0 2 13 7 0 2
31 9 3 0 0 9 1 9 1 9 13 3 9 2 16 15 13 12 3 0 0 9 2 10 9 13 1 9 0 0 9 2
11 0 1 15 13 1 0 0 9 1 9 2
31 0 0 9 1 9 12 13 0 9 9 1 0 7 0 9 2 0 1 0 0 9 7 0 9 2 1 10 9 15 13 2
19 3 1 10 0 9 0 9 13 0 13 0 0 9 1 10 9 7 9 2
30 1 10 9 13 7 13 15 9 2 16 1 0 9 13 0 13 0 9 9 7 9 2 7 13 3 2 1 9 9 2
6 10 9 13 3 9 2
23 9 0 13 1 9 1 15 9 1 15 15 7 13 1 0 9 7 9 13 0 0 9 2
22 9 3 0 7 0 3 13 0 2 0 9 2 3 9 2 0 1 9 7 0 9 2
35 9 1 15 2 16 9 15 1 15 15 13 2 13 1 9 9 2 15 9 13 3 3 0 9 2 0 1 9 1 9 2 0 0 9 2
41 1 10 9 13 0 9 0 9 2 0 10 9 1 0 9 10 7 10 0 9 2 14 0 0 9 2 15 15 1 10 9 1 9 0 9 7 0 9 3 13 2
16 0 9 13 1 10 9 0 9 2 15 14 13 0 9 9 2
6 1 9 7 13 13 2
14 1 9 1 3 0 9 7 0 9 13 0 0 9 2
52 9 7 9 1 9 3 0 9 2 3 0 9 7 9 13 13 7 3 13 1 10 0 9 2 10 0 9 15 3 13 2 13 1 9 3 3 0 0 9 2 15 1 10 9 13 14 1 0 7 0 9 2
48 1 9 9 13 2 16 1 9 13 0 9 2 13 10 9 9 0 9 2 16 0 9 13 3 0 0 9 2 16 15 9 2 1 15 1 9 0 9 13 2 4 13 0 9 2 0 9 2
24 10 9 0 9 13 7 3 0 7 0 9 9 2 7 3 7 0 7 0 9 1 10 9 2
28 0 13 9 2 16 15 3 13 3 13 0 9 1 9 2 9 2 9 7 9 2 1 9 0 9 0 9 2
29 0 13 9 2 16 15 9 10 9 13 13 0 9 9 9 2 16 3 0 0 9 15 13 1 0 9 0 9 2
40 1 9 0 9 2 15 15 3 13 0 0 9 2 13 13 0 9 0 7 1 0 1 10 9 3 3 0 9 10 9 1 0 9 0 9 1 12 2 9 2
74 13 15 0 2 16 14 9 1 9 2 7 3 9 7 0 0 9 2 0 1 0 9 9 7 0 9 2 13 0 9 15 2 16 10 9 3 3 2 7 3 14 13 0 7 0 9 2 0 9 2 16 9 13 0 9 2 15 1 10 9 13 10 0 9 7 13 3 1 15 7 10 0 9 2
16 13 15 7 2 16 16 9 13 2 13 13 10 0 0 9 2
42 1 10 9 1 15 2 15 1 0 9 3 13 1 9 9 2 13 15 3 13 1 9 2 7 3 13 0 9 2 7 15 2 15 3 7 3 13 7 13 9 0 2
26 13 13 2 16 0 9 9 0 1 0 9 13 0 9 1 9 9 1 9 7 0 9 1 10 9 2
36 3 0 15 15 13 7 0 0 0 9 7 9 2 15 13 9 1 9 2 15 13 9 13 15 0 9 7 3 1 9 9 13 7 10 9 2
4 9 9 1 11
2 11 11
20 0 9 15 1 10 9 13 13 1 0 2 13 3 0 2 0 9 0 9 2
30 0 9 2 3 9 11 2 4 15 13 13 1 15 3 3 2 1 15 3 15 1 15 13 9 7 9 0 0 9 2
13 13 9 2 1 15 15 9 3 13 2 13 9 2
24 15 13 0 0 9 11 9 12 2 7 0 9 9 12 7 12 2 3 13 9 10 9 0 2
20 16 15 10 0 9 13 13 9 9 1 15 7 1 11 2 13 15 3 0 2
27 3 2 16 1 9 13 9 9 3 3 9 16 1 15 2 3 1 0 9 2 2 7 13 15 3 3 2
14 9 11 9 13 9 1 0 12 9 13 1 12 9 2
11 15 13 0 7 13 15 15 1 0 9 2
33 9 3 13 1 9 2 16 3 13 1 9 2 3 4 13 9 0 9 2 1 9 2 3 9 13 3 9 16 9 1 0 9 2
11 13 4 3 4 3 13 9 9 16 9 2
37 7 15 13 2 16 3 1 10 0 9 13 3 3 9 2 9 7 9 16 0 9 7 0 0 9 15 4 13 3 1 0 2 0 7 0 9 2
9 10 9 15 3 1 0 9 13 2
9 13 15 15 3 9 1 0 9 2
11 7 1 10 9 15 3 11 1 11 13 2
24 16 3 7 10 9 9 0 9 3 13 1 9 9 7 9 2 13 15 13 1 12 9 3 2
30 13 15 2 16 4 1 9 12 9 13 3 13 7 3 4 13 12 9 9 3 16 9 1 9 0 2 0 9 9 2
16 0 9 4 3 13 0 9 9 2 1 15 4 3 13 9 2
17 9 4 13 0 9 1 9 9 1 9 2 3 1 9 0 9 2
11 9 9 9 4 13 1 9 13 2 2 2
4 1 10 9 2
4 15 3 0 2
9 9 9 4 9 13 9 1 9 2
11 15 4 13 1 9 2 9 2 0 9 2
21 13 0 15 13 2 16 4 9 10 3 0 9 3 13 7 13 15 13 0 9 2
2 3 2
25 3 2 3 3 4 13 9 9 7 9 2 4 4 3 3 13 1 9 7 1 15 7 0 9 2
12 13 7 15 2 16 10 9 4 13 3 0 2
18 12 9 4 9 13 2 16 3 13 3 13 7 9 15 7 13 13 2
10 1 9 4 15 13 9 7 9 9 2
6 1 15 0 16 3 2
20 0 9 9 13 3 3 0 2 7 3 1 9 4 13 3 0 7 3 0 2
15 0 9 13 0 9 1 0 9 7 3 14 13 3 13 2
15 10 3 0 0 9 1 0 9 13 9 7 13 10 9 2
32 9 0 0 9 1 0 9 13 1 0 9 2 1 3 0 9 13 3 1 15 0 1 9 9 3 9 16 1 9 12 2 2
16 13 15 15 1 0 0 7 0 9 2 3 4 13 9 2 2
26 15 4 1 15 13 11 2 3 15 13 2 16 1 9 1 11 4 13 13 10 9 14 12 12 9 2
13 0 9 1 0 9 13 3 2 16 4 15 13 2
23 13 15 1 12 9 0 2 16 9 13 1 0 9 3 0 9 16 0 9 1 9 12 2
23 3 1 12 9 2 3 3 4 3 13 9 11 2 4 0 9 11 13 13 3 16 3 2
12 1 9 0 9 4 9 14 13 13 0 9 2
17 7 16 0 9 13 3 0 2 9 9 3 13 1 9 9 9 2
16 3 2 15 0 9 13 1 9 3 3 0 2 16 15 0 2
5 11 13 13 0 9
5 11 2 0 11 2
17 9 0 0 9 9 11 11 13 0 9 2 15 15 13 1 11 2
11 13 15 1 11 9 9 9 11 11 11 2
28 9 9 9 0 9 11 11 13 2 16 0 9 2 15 4 13 9 1 11 13 2 4 13 3 1 9 11 2
7 11 13 1 14 12 9 2
14 13 4 15 13 1 12 9 0 9 3 1 0 9 2
12 11 1 9 0 9 13 0 9 2 16 13 2
18 0 0 9 11 11 15 1 10 0 9 13 1 0 9 1 11 3 2
8 0 9 13 9 1 0 9 2
17 10 9 14 13 9 11 2 15 15 13 9 12 2 9 9 11 2
2 9 11
4 1 0 0 9
8 11 11 2 11 2 9 9 2
16 9 0 15 9 2 9 0 11 2 11 12 2 12 9 2 2
49 9 2 15 3 13 12 1 9 0 9 1 9 2 9 2 9 2 9 7 0 9 2 1 10 9 3 13 9 0 9 2 7 0 9 13 7 9 9 2 16 9 3 13 13 0 9 0 9 2
23 11 1 15 13 7 13 9 0 9 1 9 0 7 0 9 2 7 15 1 12 0 9 2
21 1 0 13 1 0 9 0 9 2 15 13 1 9 9 0 0 0 9 7 9 2
12 1 0 1 9 1 0 7 0 1 0 9 2
22 1 0 1 0 0 2 0 9 0 9 2 15 13 3 0 0 2 0 7 0 9 2
22 1 0 13 1 0 9 9 7 9 7 10 9 1 9 2 0 9 7 9 0 9 2
15 9 9 2 9 0 9 2 13 1 11 3 9 0 9 2
8 11 11 2 9 13 1 9 2
19 9 9 1 9 7 0 2 9 0 11 2 11 12 2 12 9 2 2 2
43 9 13 13 1 0 9 2 13 1 15 0 9 7 13 3 12 9 1 15 2 16 4 15 13 7 13 0 9 9 7 13 15 1 9 3 2 16 4 1 15 13 0 2
29 0 9 3 7 3 0 9 13 13 15 13 15 0 9 7 13 15 2 15 15 13 7 15 13 13 1 0 9 2
21 13 9 1 15 2 16 9 13 13 14 15 2 15 13 0 1 9 13 0 9 2
63 9 2 9 9 7 9 1 9 9 9 7 0 9 2 9 7 0 9 2 13 2 3 10 0 9 13 3 2 16 4 15 13 9 2 3 13 0 0 9 7 13 9 0 9 2 3 13 9 7 15 13 10 0 9 7 9 2 3 15 13 1 9 2
7 11 11 2 3 13 9 2
15 9 9 2 9 0 11 2 11 12 2 12 9 2 2 2
21 0 9 4 13 10 0 9 0 12 9 2 16 0 9 13 1 10 9 3 12 2
22 7 15 13 14 9 1 15 2 16 4 15 9 1 0 9 9 13 9 0 0 9 2
24 9 2 9 9 9 0 0 9 11 0 2 1 0 9 7 0 9 13 0 9 9 0 9 2
30 9 1 9 13 9 15 13 3 9 9 7 9 9 9 9 2 9 9 1 9 9 2 9 9 9 7 9 9 9 2
38 13 1 0 9 2 15 15 9 1 9 9 13 2 13 15 7 1 9 9 1 10 9 13 0 9 2 16 15 1 0 9 9 7 1 10 9 13 2
4 9 1 9 12
22 0 9 2 15 13 1 0 9 1 11 2 15 13 13 10 9 1 0 12 0 9 2
32 0 0 7 0 9 11 1 9 13 0 7 0 9 3 0 9 2 9 2 9 7 0 9 1 9 9 7 3 0 9 9 2
12 9 15 13 7 1 0 9 7 9 1 9 2
4 9 11 13 3
4 11 11 2 11
20 1 9 9 7 9 11 11 15 3 13 1 10 0 0 9 0 9 0 9 2
21 9 9 11 2 11 13 10 0 9 2 1 15 4 13 12 9 7 12 0 9 2
25 13 2 16 7 1 15 9 2 15 15 1 10 9 13 2 13 1 10 9 3 0 9 0 9 2
26 1 10 9 13 9 9 1 9 0 9 7 0 9 0 0 9 2 12 9 2 15 13 9 0 9 2
26 13 15 1 9 2 3 1 0 9 1 9 13 0 9 2 15 13 1 9 0 9 7 9 0 9 2
29 13 9 2 16 0 9 4 13 1 9 0 9 1 9 0 9 7 13 15 13 9 7 0 9 3 1 0 9 2
7 11 15 13 13 9 1 11
2 11 2
29 9 2 16 4 12 9 0 9 13 11 1 9 9 2 13 3 1 9 1 9 0 9 0 9 9 11 11 11 2
29 1 9 9 2 15 15 13 1 0 9 1 0 9 11 2 3 15 13 9 9 2 13 11 9 1 12 2 9 2
20 13 2 16 10 9 13 13 9 11 2 15 1 0 9 1 11 13 0 9 2
14 9 0 0 9 14 11 13 7 13 15 1 12 9 2
6 0 9 1 9 1 11
2 11 2
18 1 9 1 9 11 1 0 9 2 11 2 13 1 0 9 0 9 2
7 9 13 0 9 16 0 2
12 13 15 3 9 11 1 9 1 0 0 9 2
16 9 0 9 1 0 9 10 9 3 13 7 13 10 0 9 2
28 1 9 13 1 9 14 0 9 0 9 2 15 13 9 7 0 9 2 13 9 9 1 0 9 11 2 11 2
5 9 9 15 13 2
9 0 9 4 1 11 13 4 3 13
4 11 2 11 2
17 9 1 0 0 0 9 0 1 12 2 9 4 13 4 3 13 2
10 13 15 3 1 0 9 9 11 11 2
32 1 9 9 9 9 9 1 9 9 13 2 16 11 13 9 13 1 15 2 16 4 13 9 0 9 1 3 0 0 9 11 2
11 1 10 9 4 9 13 4 13 2 13 2
43 9 2 15 15 1 0 9 1 9 0 9 13 1 0 9 13 3 1 12 2 9 2 4 1 9 1 9 1 9 9 13 3 1 12 2 9 7 3 1 12 2 9 2
19 11 7 11 3 13 2 16 15 13 1 0 9 0 9 9 9 0 9 2
20 11 4 15 3 13 1 11 0 0 9 2 15 3 13 0 9 1 0 9 2
5 9 14 1 11 13
4 11 2 11 2
18 9 11 11 12 2 3 13 2 16 4 13 0 9 3 9 13 11 2
20 13 2 16 1 0 9 13 9 9 1 9 2 15 13 1 0 0 9 13 2
11 13 15 3 0 9 11 2 11 2 11 2
16 9 15 14 13 13 1 0 11 2 1 9 9 7 0 11 2
18 3 16 12 5 0 11 15 1 9 13 1 9 1 0 9 1 11 2
14 1 11 1 11 15 3 3 13 9 0 9 11 11 2
9 9 15 13 12 9 15 0 9 2
14 1 11 4 3 13 12 9 1 0 0 9 9 11 2
9 1 9 13 3 13 1 0 9 2
6 9 15 13 10 9 2
7 13 15 9 0 9 11 2
22 12 1 0 9 1 9 9 1 11 13 13 9 9 0 9 2 3 1 11 7 11 2
12 1 11 15 3 13 0 9 9 11 2 11 2
13 10 9 13 7 9 11 11 7 9 9 11 11 2
15 16 13 2 11 13 9 9 1 0 0 9 2 11 2 2
15 13 7 2 16 4 1 9 11 1 0 11 13 0 9 2
4 11 13 0 9
5 11 2 0 11 2
25 12 11 2 15 15 13 13 1 9 0 9 11 2 4 3 13 2 16 12 1 15 13 1 9 2
8 13 15 3 9 9 1 11 2
24 1 9 11 15 13 2 16 12 11 15 13 13 0 9 2 15 13 9 1 9 1 0 9 2
12 0 9 15 7 1 9 13 1 9 1 9 2
23 16 9 9 1 11 1 0 11 13 2 13 3 1 0 11 0 2 0 9 1 9 9 2
15 0 9 13 1 15 2 16 4 15 9 13 1 9 9 2
11 11 7 13 1 9 9 7 1 0 9 2
4 9 13 1 9
8 0 0 9 0 9 9 3 13
4 11 2 11 2
23 9 2 15 13 0 0 9 2 11 2 2 13 1 0 11 1 9 3 1 12 0 9 2
14 13 15 3 12 9 3 2 16 11 10 10 9 13 2
25 1 9 9 15 1 11 9 1 9 13 1 0 9 2 1 9 2 15 13 13 1 0 9 9 2
10 1 9 3 13 0 9 1 0 9 2
31 15 15 7 3 2 16 13 9 9 1 9 0 0 9 2 13 9 0 9 0 9 2 0 1 9 0 11 1 0 9 2
23 11 11 2 9 0 9 11 11 2 0 9 11 2 13 2 16 11 13 9 1 15 9 2
29 0 0 9 3 13 2 16 13 1 9 1 9 9 2 15 4 13 14 10 9 1 15 2 16 9 13 1 9 2
18 1 9 1 9 11 15 13 0 0 0 9 0 0 9 2 11 2 2
16 9 1 11 0 9 13 1 9 1 9 1 9 1 0 9 2
29 9 0 9 1 15 2 16 11 13 1 10 0 9 0 9 16 0 2 3 13 9 2 16 9 13 3 3 0 2
28 16 13 1 11 3 9 2 13 1 9 2 15 15 3 13 1 9 2 3 13 9 2 13 3 0 9 11 2
22 1 9 0 0 11 13 9 1 0 9 7 0 9 1 0 11 0 9 9 16 9 2
22 16 9 13 12 9 2 0 9 1 9 13 13 1 9 2 16 4 13 9 1 11 2
22 11 11 7 13 1 9 13 2 16 13 0 2 16 15 9 13 9 3 2 13 9 2
2 0 9
14 12 2 12 2 0 9 0 2 9 2 9 0 9 11
14 12 2 12 2 0 0 9 0 2 9 2 11 11 11
12 12 2 12 2 9 9 13 3 2 0 9 11
15 12 2 12 2 0 9 0 2 9 2 0 0 0 9 11
11 9 13 1 0 9 1 0 11 9 0 11
2 9 11
4 9 1 11 13
2 11 2
12 11 3 13 3 0 9 9 1 0 0 9 2
29 1 9 0 0 9 0 9 7 9 9 0 9 1 0 11 7 4 1 9 3 1 9 12 13 9 12 9 9 2
20 1 9 12 13 9 9 1 12 2 15 13 1 12 9 3 16 1 9 12 2
7 9 10 9 13 9 9 2
14 1 9 15 4 13 0 9 1 0 9 7 9 9 2
23 1 9 0 9 1 9 9 1 9 12 13 3 0 9 9 1 10 9 7 3 0 9 2
51 1 0 9 1 9 9 9 13 13 9 9 9 1 9 1 9 1 12 9 2 9 9 9 1 12 9 9 9 7 1 9 12 9 1 9 1 0 9 1 9 1 12 9 2 15 3 13 1 11 0 2
24 1 9 2 3 13 9 9 2 15 1 9 13 12 9 11 1 0 0 9 7 0 9 9 2
10 3 12 9 13 1 9 9 1 9 2
22 9 0 9 7 3 0 0 9 9 9 11 13 1 9 9 0 9 9 1 0 9 2
12 3 0 9 13 1 0 9 9 13 9 9 2
16 3 4 3 13 9 1 9 9 2 15 13 13 3 3 0 2
19 0 9 9 3 13 9 0 9 2 7 3 15 13 1 9 12 2 9 2
34 9 9 1 9 9 9 15 3 13 16 0 16 3 9 0 0 9 2 16 3 1 9 7 1 0 11 1 0 9 12 2 9 2 2
13 1 0 0 9 15 9 1 9 3 13 0 9 2
17 1 9 12 15 3 13 9 9 1 12 9 7 9 1 12 9 2
37 0 9 3 1 11 13 0 0 9 2 15 13 1 9 11 1 0 11 2 1 9 0 11 1 9 7 3 3 1 9 0 11 1 9 7 9 2
5 1 9 13 1 9
12 11 2 11 7 11 15 13 2 16 3 13 13
10 0 9 1 0 9 11 11 2 11 11
33 13 15 3 2 16 15 15 10 9 13 2 14 3 4 15 13 13 9 1 0 9 0 9 9 11 11 1 0 0 9 1 11 2
31 9 11 13 9 13 9 9 11 7 13 4 15 4 2 7 3 7 13 2 9 0 0 9 1 9 1 0 9 0 9 2
16 13 7 2 16 4 15 1 10 9 13 13 7 1 0 11 2
6 15 13 0 0 9 2
5 9 11 15 13 2
13 7 2 3 13 0 0 9 2 13 15 13 15 2
21 16 1 0 9 13 3 9 9 2 16 9 9 13 3 13 15 2 7 13 15 2
17 11 1 10 0 9 13 9 1 11 2 16 4 15 13 0 9 2
17 9 0 9 9 13 0 9 2 4 15 13 0 9 1 9 11 2
26 3 13 0 9 1 11 1 9 11 1 0 2 0 2 7 0 2 9 2 16 4 13 9 10 9 2
26 0 9 15 1 0 9 13 13 12 9 2 1 0 9 2 12 2 7 3 15 13 2 16 9 13 2
4 9 15 13 2
7 3 2 13 15 13 15 2
33 13 15 3 11 11 2 13 15 2 16 3 1 15 15 13 9 9 2 2 7 13 2 16 0 9 13 0 9 1 9 1 9 2
11 13 15 3 11 11 2 15 0 9 13 2
31 1 10 9 15 14 15 0 13 2 16 2 3 13 2 13 1 3 0 9 7 13 13 9 2 16 4 1 15 13 13 2
22 3 2 9 9 0 0 9 1 11 13 14 13 9 0 9 7 3 0 2 0 9 2
17 3 2 9 9 11 14 13 13 3 1 11 9 9 1 0 9 2
18 3 16 3 3 1 9 0 9 13 7 15 13 0 9 9 11 11 2
34 1 9 1 9 13 3 11 11 7 13 15 2 16 15 13 3 2 16 13 15 14 9 9 7 15 16 4 13 9 0 7 0 9 2
24 16 4 4 11 1 9 9 11 13 3 7 1 0 9 2 15 4 15 4 4 1 9 13 2
30 11 13 2 16 0 9 9 3 13 2 7 1 15 13 10 9 2 7 16 15 9 11 13 13 15 1 11 2 13 2
4 3 14 3 2
11 15 3 15 13 0 7 0 9 1 11 2
34 13 15 2 16 15 9 13 2 0 9 4 13 2 15 3 13 1 0 9 2 1 15 3 13 2 7 11 11 0 9 1 11 13 2
18 3 3 1 9 13 14 0 9 2 15 3 9 3 13 2 16 13 2
13 15 2 16 9 0 9 13 2 14 13 9 9 2
3 9 0 9
9 0 9 9 1 0 11 1 0 9
20 9 9 9 1 11 15 3 13 1 15 9 3 12 0 2 13 4 12 9 2
9 0 9 13 0 9 1 0 9 2
21 12 2 12 2 9 0 9 2 10 9 13 7 0 0 9 2 7 0 0 9 2
22 9 12 2 1 9 0 9 13 0 9 1 0 11 0 9 2 15 13 13 0 9 2
14 9 12 2 9 0 9 13 0 9 0 11 1 11 2
8 9 13 0 9 1 0 11 2
4 0 9 13 2
15 9 12 2 13 13 0 9 0 11 2 0 1 9 12 2
10 1 0 0 0 9 13 7 0 9 2
19 9 12 2 1 0 9 0 9 1 9 9 1 0 9 13 9 0 9 2
7 13 3 0 9 1 11 2
10 9 12 2 1 0 11 13 0 9 2
13 9 12 2 0 9 13 9 1 0 9 0 11 2
24 9 12 2 9 9 0 11 7 11 11 11 7 11 11 15 13 1 9 0 2 0 0 9 2
7 0 11 1 15 13 13 2
7 13 1 0 9 0 11 2
12 9 12 2 0 9 13 9 1 0 9 9 2
9 9 12 2 13 12 0 0 9 2
14 12 9 13 11 11 2 13 15 7 1 10 9 13 2
12 1 9 1 0 9 13 9 9 7 0 9 2
5 9 9 12 13 2
31 9 12 2 9 1 0 11 7 0 9 2 15 13 9 0 11 1 0 11 7 0 9 13 0 0 9 1 9 0 11 2
7 9 13 9 9 7 9 2
30 9 12 2 9 1 9 11 1 11 1 0 0 9 7 0 0 9 1 9 7 3 0 0 9 7 9 9 1 9 2
17 9 13 2 9 13 13 9 9 1 0 9 7 9 1 0 9 2
22 9 12 2 0 11 13 0 9 9 1 0 0 9 1 0 11 1 9 13 9 9 2
7 13 1 0 9 16 0 2
24 9 12 2 0 0 9 11 11 2 3 0 7 0 9 2 7 9 11 11 11 11 13 9 2
8 1 10 9 13 3 0 9 2
16 9 12 2 11 11 13 0 9 9 1 9 9 1 0 11 2
23 9 12 2 11 11 13 2 16 13 0 9 1 9 2 16 15 9 7 9 13 1 9 2
11 13 10 9 1 11 2 16 15 13 9 2
8 13 15 1 9 0 0 9 2
23 11 11 13 2 16 9 4 13 4 13 1 9 2 16 4 4 13 10 7 0 0 9 2
26 12 2 9 12 2 0 0 9 9 1 9 11 7 0 0 9 13 9 0 0 9 1 9 0 9 2
18 12 2 9 12 2 11 11 13 9 1 11 11 2 16 11 13 9 2
15 0 9 13 13 15 9 2 1 15 4 13 13 11 11 2
40 12 2 9 12 2 0 9 11 11 7 0 9 11 11 13 1 11 9 0 9 0 9 1 0 11 2 13 9 12 9 2 16 4 13 9 9 1 0 9 2
18 12 2 9 12 2 9 1 9 11 13 2 16 4 13 1 0 9 2
34 12 2 9 12 2 0 9 13 9 11 1 12 2 9 1 9 2 16 11 13 1 9 2 13 12 0 9 1 9 11 1 11 2 2
16 12 2 9 12 2 11 11 13 0 9 1 0 9 1 9 2
12 11 11 15 13 2 16 15 9 13 9 3 2
24 12 2 9 12 2 9 11 11 13 9 11 7 0 11 1 9 0 9 9 1 9 0 9 2
29 12 2 9 12 2 11 11 2 9 11 11 2 1 9 1 9 1 11 13 2 16 1 12 9 11 13 0 9 2
18 9 9 12 2 11 13 12 2 9 9 0 9 1 11 9 0 9 2
4 0 9 1 9
11 0 9 1 9 11 1 12 9 9 9 11
2 11 2
32 3 16 1 11 15 3 1 0 0 11 13 0 9 2 10 9 13 13 9 0 1 9 0 0 9 1 0 9 0 0 9 2
37 1 0 9 13 1 10 9 2 7 1 0 9 2 15 1 0 9 13 0 0 9 11 2 16 1 9 12 1 9 1 0 11 13 9 9 11 2
29 0 9 11 13 2 16 11 13 1 0 9 14 12 9 9 2 3 9 9 2 15 13 1 0 9 1 0 11 2
19 13 3 1 9 2 16 4 15 15 13 0 9 2 15 13 1 0 9 2
23 9 15 13 1 9 0 9 11 1 0 9 0 11 2 15 13 0 9 1 9 10 9 2
28 9 1 9 9 15 13 0 9 7 9 2 15 15 3 13 2 7 16 3 14 13 0 0 9 10 0 9 2
13 0 9 15 7 13 7 9 9 13 9 1 9 2
28 15 14 13 9 0 9 2 15 15 13 1 9 1 0 9 7 13 3 2 3 1 0 0 9 0 9 13 2
27 7 15 15 7 13 13 14 0 9 1 9 0 9 7 9 2 10 9 15 7 1 9 0 9 13 13 2
11 1 0 9 13 10 9 0 7 3 0 2
27 13 15 3 2 16 0 0 9 13 10 9 1 0 0 9 1 9 2 9 7 9 11 1 9 1 9 2
23 1 15 3 13 1 9 12 7 3 15 15 1 0 9 13 2 16 4 15 15 3 13 2
27 3 13 1 9 0 9 9 0 9 2 15 13 1 0 9 0 9 1 0 9 0 9 9 0 9 13 2
11 0 9 15 3 13 1 11 7 0 9 2
45 9 1 9 13 3 3 2 3 9 9 1 11 13 1 0 0 9 0 9 7 0 0 7 0 9 2 13 0 9 7 13 2 16 1 0 9 4 3 10 9 13 9 0 9 2
8 0 9 1 0 9 4 13 9
4 11 11 2 9
44 13 3 9 2 15 3 13 9 9 0 9 1 0 9 2 9 2 15 13 2 16 10 0 9 13 3 13 2 16 9 1 9 13 13 10 9 2 16 9 9 13 3 0 2
32 13 7 15 2 16 13 15 9 3 0 2 16 3 13 11 2 13 2 16 15 0 0 9 9 0 0 9 1 9 7 13 2
14 10 9 13 9 2 15 15 13 13 3 0 12 9 2
20 15 4 15 7 13 2 16 4 0 9 1 0 9 0 9 3 14 13 4 2
17 3 13 15 2 0 0 9 13 9 2 15 4 13 4 3 13 2
51 15 1 15 13 9 2 16 0 9 0 9 2 1 9 0 7 3 0 2 0 9 13 0 9 2 0 1 10 9 7 9 12 9 0 0 9 2 3 15 2 15 15 1 10 10 9 1 0 9 13 2
38 15 1 15 13 7 9 2 16 9 0 9 3 1 0 12 9 13 9 2 15 15 13 0 9 10 9 7 1 9 11 7 11 10 9 3 3 13 2
18 1 15 3 2 13 2 14 9 0 9 2 15 0 9 13 0 9 2
18 9 0 2 7 13 15 13 2 16 3 0 2 9 7 13 9 9 2
28 9 2 16 15 0 9 0 9 1 0 0 9 2 15 0 9 13 2 13 3 1 9 1 11 7 11 11 2
42 0 2 0 2 0 9 13 0 9 2 0 0 9 2 3 9 1 9 15 2 15 15 13 2 9 9 0 9 2 0 9 0 9 2 7 3 7 0 0 9 9 2
8 7 10 0 9 1 15 13 2
8 9 13 2 16 1 15 13 2
24 1 9 0 0 9 4 15 7 15 7 0 9 13 1 0 9 3 3 16 3 9 0 15 2
49 13 2 14 15 9 0 2 15 3 0 9 2 4 0 9 13 1 9 3 0 0 9 2 4 3 1 9 13 9 0 2 4 15 15 9 13 13 9 9 2 7 3 15 4 3 7 3 13 2
8 15 15 1 9 1 0 9 2
25 13 3 2 16 0 9 1 0 9 13 0 9 1 9 0 9 2 3 15 13 7 3 13 9 2
15 13 3 9 2 16 0 0 9 13 1 15 0 9 3 2
11 10 9 7 13 0 9 9 7 9 9 2
34 13 1 9 1 9 10 9 2 15 13 9 2 16 9 9 7 10 9 13 0 9 2 1 12 1 10 9 13 1 9 13 1 0 2
4 13 9 0 2
25 0 9 9 2 0 0 0 9 2 3 13 0 9 7 13 0 9 1 9 2 16 15 13 0 2
32 0 0 9 1 11 13 0 9 2 3 13 9 2 3 10 9 2 0 9 15 15 7 1 10 9 3 1 0 9 13 13 2
29 9 13 0 9 2 15 3 13 9 12 5 9 2 15 13 3 1 11 7 9 9 2 15 13 0 0 0 9 2
11 15 13 0 0 9 2 0 9 7 9 2
11 14 9 11 13 9 1 9 7 3 13 2
30 0 9 1 0 9 4 3 3 13 1 9 13 0 9 2 7 13 1 0 9 2 2 15 4 13 9 1 0 9 2
38 13 3 0 2 16 9 4 15 13 1 0 9 2 3 3 9 2 9 2 9 0 9 2 13 1 9 2 7 15 1 0 0 9 2 13 3 13 2
13 13 3 2 16 0 9 1 0 9 13 9 0 2
14 13 4 1 9 1 9 9 9 2 9 9 0 9 2
14 9 13 10 9 16 15 2 7 13 13 1 10 9 2
10 10 9 13 0 9 2 3 9 9 2
20 13 1 15 2 16 4 13 0 9 9 7 16 4 3 13 9 1 0 9 2
4 9 7 9 9
4 11 11 2 9
37 7 0 9 15 13 0 2 0 9 15 1 15 13 0 9 2 1 15 15 13 3 13 2 16 4 15 15 13 2 16 13 1 9 9 7 9 2
29 10 9 3 13 1 9 7 0 9 2 15 3 13 9 2 7 3 13 0 9 0 9 2 0 9 7 0 9 2
40 13 15 2 16 9 15 13 13 1 9 10 9 13 7 13 9 7 10 0 9 16 15 2 15 3 13 2 0 0 9 2 1 15 15 13 14 10 9 9 2
9 9 0 9 9 13 1 0 9 2
18 13 4 13 10 0 9 2 15 4 1 9 3 0 9 13 0 9 2
48 15 15 13 9 1 0 9 2 13 2 16 0 9 13 10 9 2 0 9 1 0 9 2 9 13 9 1 0 0 9 2 0 0 9 2 0 9 2 0 9 2 15 13 3 0 9 9 2
11 0 9 2 10 9 9 2 15 9 13 2
46 0 9 2 15 15 3 13 1 0 9 2 3 3 13 1 0 9 2 1 9 2 3 15 13 13 2 16 0 9 13 9 2 13 15 1 9 1 10 9 0 9 7 13 0 9 2
46 9 15 3 13 2 16 13 1 0 0 9 2 15 13 0 0 9 9 13 1 9 2 7 1 3 0 9 2 1 10 9 13 14 0 9 2 7 7 0 9 3 3 14 9 11 2
12 1 9 2 10 0 9 13 15 1 12 9 2
24 9 2 15 9 0 13 1 9 2 16 4 3 13 9 10 9 2 13 1 9 1 9 9 2
31 9 2 1 10 0 9 2 16 4 15 13 2 16 9 9 13 13 9 0 0 9 2 13 10 9 0 9 2 0 9 2
3 9 13 2
12 0 9 13 9 2 15 13 9 2 15 9 2
7 0 9 4 13 9 0 2
9 13 9 3 2 9 1 15 3 2
17 16 9 10 9 9 13 2 13 15 9 13 0 9 2 9 9 2
10 9 15 13 3 7 13 0 2 15 2
15 15 9 13 2 13 1 0 9 2 13 2 14 15 13 2
28 15 15 3 13 9 1 9 2 16 4 3 13 15 2 15 15 3 15 13 2 13 15 3 7 13 4 0 2
18 3 9 1 9 3 13 9 0 9 2 16 4 15 15 3 3 13 2
12 7 7 4 13 0 9 13 1 10 0 9 2
12 0 9 2 15 1 15 13 9 2 15 13 2
9 0 9 1 15 15 13 13 15 2
18 13 3 1 15 2 16 9 0 9 13 1 9 9 1 9 0 9 2
11 1 9 9 13 15 0 9 1 0 9 2
7 13 15 1 3 0 9 2
19 3 14 13 9 1 9 9 2 3 13 9 2 9 9 2 3 15 13 2
7 9 0 2 9 7 0 2
6 1 9 9 13 9 2
11 7 14 3 2 0 9 13 3 0 9 2
10 13 2 16 1 0 9 15 4 13 2
5 16 1 0 9 2
16 9 15 13 2 7 15 3 13 0 9 2 16 9 10 9 2
8 3 15 13 7 10 9 0 2
10 9 13 9 2 15 13 7 15 9 2
50 0 9 13 13 13 9 0 9 7 13 15 0 0 9 7 0 9 10 0 9 1 9 2 16 13 0 7 0 0 9 2 15 1 9 2 3 9 13 13 1 9 9 2 3 13 0 16 0 9 2
3 9 0 9
4 11 11 2 9
23 1 9 9 0 9 13 1 0 9 0 9 1 9 13 0 0 9 2 0 1 9 9 2
14 15 1 9 0 13 0 9 1 9 3 0 0 9 2
13 13 9 7 13 3 1 15 2 13 14 1 9 2
17 1 10 9 15 3 13 0 0 9 2 16 4 15 13 9 15 2
29 0 9 1 0 9 1 9 12 13 3 1 9 1 12 9 0 9 2 16 1 15 1 9 13 3 9 1 9 2
23 13 15 9 2 3 3 13 3 0 9 2 7 0 3 2 16 13 1 15 3 0 9 2
51 0 0 9 2 15 3 9 13 2 13 1 9 1 9 0 9 2 9 2 1 15 13 0 15 13 2 1 15 13 0 16 0 7 0 0 9 2 10 9 4 15 3 13 2 13 9 2 10 9 13 2
23 9 0 9 13 12 0 9 2 15 4 13 4 3 13 2 15 13 1 0 9 0 9 2
14 9 12 9 0 9 3 13 2 0 13 9 0 9 2
43 0 9 3 13 12 0 9 2 9 2 9 0 9 7 9 2 0 9 0 1 10 9 2 3 3 2 3 15 9 1 9 0 9 3 13 2 7 0 9 0 0 9 2
30 1 0 9 13 9 0 9 2 15 0 9 13 3 9 0 9 2 3 2 3 15 13 2 14 13 9 0 0 9 2
30 11 3 13 9 13 9 0 0 9 0 9 2 16 15 13 13 1 9 9 9 0 7 9 0 13 0 9 3 13 2
20 1 0 9 3 13 9 3 0 2 1 9 0 9 1 9 3 0 0 9 2
18 13 3 9 9 9 1 9 11 7 13 15 1 0 9 1 9 9 2
13 13 15 9 16 0 9 2 1 15 13 15 9 2
27 16 15 9 0 9 13 1 9 9 0 9 2 13 9 9 13 2 13 10 10 9 2 13 7 13 9 2
15 9 2 15 1 9 0 0 9 3 13 2 13 9 9 2
11 13 1 10 0 9 1 9 13 0 9 2
5 1 9 3 13 2
22 1 9 9 4 13 3 1 15 2 16 4 15 0 0 0 9 13 3 13 1 9 2
22 13 3 0 9 0 0 9 1 9 3 0 0 9 15 7 13 9 0 9 1 9 2
8 0 9 13 9 9 2 12 2
1 9
4 9 2 11 11
25 1 0 9 9 0 1 0 9 15 4 13 9 0 9 1 0 9 7 3 0 9 9 0 9 2
55 0 9 0 9 0 1 0 9 13 10 9 1 0 9 1 9 12 2 12 0 9 2 15 15 13 1 0 9 0 10 9 2 7 2 3 1 0 0 9 0 1 9 1 10 0 9 7 1 10 0 9 0 1 9 2
14 0 9 13 0 1 0 9 0 9 2 0 0 9 2
40 0 0 9 13 9 9 2 9 13 0 9 2 1 15 13 9 13 1 10 9 1 0 9 9 0 9 7 1 15 3 9 13 9 9 3 9 1 9 2 2
36 13 15 15 2 16 9 10 9 2 7 2 9 2 15 9 13 2 13 1 9 9 0 0 9 13 13 0 9 1 9 2 0 2 9 2 2
27 4 2 14 9 0 1 9 3 7 3 13 2 13 10 9 9 0 9 13 7 1 9 9 13 10 9 2
23 3 16 1 0 9 13 7 1 10 9 1 9 0 9 1 9 0 10 9 1 9 9 2
31 1 9 9 2 12 2 12 9 2 1 9 13 1 15 0 0 9 13 3 9 2 7 15 14 1 9 9 9 9 11 2
20 0 0 9 2 7 3 7 9 1 15 0 2 13 4 3 13 1 0 9 2
13 9 1 9 0 0 9 13 9 1 9 0 9 2
21 0 9 1 9 12 13 3 9 0 15 10 0 9 0 1 9 1 10 0 9 2
36 0 9 3 2 13 2 16 0 9 13 1 9 10 0 9 13 1 0 9 0 9 7 0 9 2 15 13 1 15 7 1 15 13 13 13 2
29 13 7 1 0 9 3 13 9 2 7 2 9 9 2 7 9 2 7 2 9 2 10 9 13 0 9 13 2 2
17 13 2 14 15 0 9 2 13 0 9 13 9 7 0 0 9 2
30 3 0 9 9 0 9 13 1 0 9 0 1 15 2 16 13 13 9 15 2 16 4 10 9 13 3 13 1 9 2
35 15 13 9 1 0 9 0 9 0 1 0 9 2 7 1 15 15 9 13 9 10 9 1 9 13 3 1 9 2 15 3 15 9 13 2
43 7 0 9 1 0 9 2 15 4 15 3 0 9 13 2 13 7 1 10 9 12 9 15 13 1 10 9 1 0 9 2 16 15 9 7 9 1 10 9 13 0 9 2
14 3 3 13 0 15 1 9 9 13 3 0 0 9 2
13 1 0 9 4 3 13 4 3 13 9 9 9 2
28 0 13 2 16 9 13 9 2 16 4 15 9 1 9 9 13 9 2 15 13 1 9 9 1 9 0 9 2
53 1 10 9 13 0 13 1 0 10 9 9 9 2 15 13 13 9 9 9 2 1 15 4 15 1 9 3 13 9 13 2 1 10 9 4 4 3 9 13 1 9 9 2 1 10 4 13 1 9 0 9 9 2
3 9 1 9
9 1 9 7 1 9 15 13 0 0
2 11 11
15 7 16 1 9 13 7 3 0 11 3 0 0 0 9 2
5 0 15 7 13 2
10 1 9 11 1 9 7 9 13 9 2
13 0 0 9 3 13 1 0 9 0 2 0 9 2
18 9 9 1 9 13 0 9 7 11 2 7 11 13 1 9 1 9 2
10 0 9 13 13 1 0 9 0 9 2
26 10 9 13 7 13 9 2 16 3 16 0 9 13 0 11 2 10 9 15 3 13 9 1 0 9 2
7 9 1 9 13 9 0 2
10 13 15 2 16 15 15 13 2 2 2
27 3 15 13 9 2 3 13 15 0 9 2 13 9 2 11 1 11 12 7 13 2 3 15 13 9 9 2
16 3 13 0 7 13 4 13 9 2 3 9 13 16 1 9 2
11 7 10 9 15 1 15 13 3 7 9 2
16 3 3 15 0 9 13 1 0 9 7 3 15 13 7 9 2
13 9 15 3 14 3 13 15 2 1 15 13 13 2
3 13 0 9
28 1 0 9 1 9 9 2 3 10 9 13 9 1 9 9 2 15 1 0 9 9 1 9 7 9 13 13 2
10 3 13 1 15 3 0 7 0 9 2
12 10 9 13 0 7 7 13 3 0 9 9 2
7 15 15 13 7 11 12 2
27 15 3 3 13 9 7 1 11 12 2 15 13 1 0 9 13 0 0 9 1 0 9 3 12 9 9 2
31 0 9 2 15 13 0 9 2 13 0 9 0 9 2 10 9 1 9 15 13 0 9 7 3 13 0 9 2 9 3 2
12 0 9 1 15 13 12 9 7 3 0 9 2
11 10 9 13 1 0 9 9 1 0 9 2
17 3 13 9 1 9 2 3 1 12 2 3 3 1 9 7 9 2
15 3 9 1 0 9 2 15 9 13 1 15 2 13 0 2
18 15 3 4 13 13 1 0 9 9 2 16 4 15 1 15 13 13 2
14 3 15 7 9 15 3 13 1 9 2 13 9 11 2
3 9 16 9
12 9 1 0 11 2 15 13 9 15 1 15 2
14 9 9 9 7 0 9 13 3 0 9 13 3 0 2
9 3 9 13 0 0 9 1 9 2
16 16 0 9 13 2 1 9 13 15 15 0 2 1 9 3 2
6 9 9 13 3 15 2
19 16 4 9 13 3 16 1 12 0 9 2 13 13 9 12 7 12 0 2
12 15 13 3 9 1 9 9 2 9 2 2 2
8 0 9 3 1 0 9 13 2
26 13 0 2 7 16 1 11 0 2 16 1 0 9 13 0 9 1 0 11 13 0 9 9 16 9 2
11 9 13 2 3 1 10 9 13 0 9 2
14 15 7 3 4 9 13 1 9 2 13 3 0 9 2
5 15 2 3 2 3
17 0 0 9 13 3 1 12 1 9 0 9 1 9 9 9 9 2
43 11 11 2 11 11 2 11 11 2 11 11 7 0 15 13 1 9 9 1 0 9 2 15 13 1 0 9 13 1 0 9 9 1 0 9 2 7 13 1 12 2 9 2
18 9 2 9 7 9 11 11 13 1 9 13 1 0 9 11 1 11 2
28 9 0 2 0 9 0 9 2 12 2 9 0 9 1 0 9 2 13 3 1 11 7 13 1 12 2 9 2
5 9 1 9 11 11
29 0 9 9 11 11 2 12 2 9 12 2 12 2 9 12 2 13 9 2 15 4 3 13 1 0 9 1 11 2
25 1 0 9 10 0 9 0 0 9 0 9 0 9 13 7 9 0 0 0 9 2 15 11 13 2
11 13 0 2 15 11 11 1 10 9 13 2
24 10 0 9 7 13 7 9 9 7 9 2 15 13 13 1 0 9 2 13 9 9 11 11 2
19 9 9 13 3 0 9 2 15 9 1 15 11 13 9 0 9 9 13 2
14 9 2 3 0 9 1 9 2 13 14 1 9 9 2
29 9 11 13 0 9 2 15 4 3 13 1 0 9 11 2 13 0 9 0 9 0 9 0 1 11 1 9 12 2
51 0 9 1 0 9 2 9 2 9 2 9 2 9 7 3 9 13 1 0 0 9 2 10 9 15 13 13 3 1 9 10 9 7 13 15 1 0 9 11 1 9 12 2 3 13 9 10 0 9 13 2
22 1 0 9 2 11 11 2 11 11 2 11 11 0 2 2 3 13 0 9 0 9 2
16 9 13 0 9 1 9 0 0 9 1 11 11 1 9 12 2
28 1 9 9 13 0 9 12 9 2 15 15 4 13 0 9 2 1 12 2 9 2 1 12 9 1 9 11 2
3 2 11 2
2 9 9
9 0 9 11 11 4 3 13 0 9
34 9 9 3 13 1 9 9 0 9 7 9 3 0 9 0 0 11 2 11 2 0 11 7 0 0 11 11 11 2 12 2 12 2 2
25 0 9 1 0 9 13 4 3 13 14 1 0 9 1 9 1 0 9 1 0 9 7 0 9 2
30 9 9 1 0 11 13 3 16 9 0 9 0 2 0 9 2 10 9 13 1 0 9 7 1 9 0 14 2 9 2
30 0 0 9 13 9 9 11 2 12 2 3 12 7 12 2 2 15 3 13 1 0 9 1 9 0 9 2 12 2 2
24 9 3 1 9 9 1 0 9 1 9 12 2 12 9 0 9 3 13 0 9 0 0 9 2
13 9 3 13 1 9 1 0 0 9 7 9 9 2
40 1 0 0 9 3 13 9 9 11 2 12 2 2 9 2 12 2 2 11 2 9 0 9 2 12 2 3 12 7 12 2 7 9 0 0 9 2 12 2 2
32 1 0 9 15 9 0 9 13 1 0 0 9 1 0 7 0 9 2 1 15 13 0 9 1 10 9 1 9 9 7 9 2
29 12 0 9 13 9 11 2 9 1 0 9 7 0 9 2 12 2 7 0 9 2 9 7 0 9 2 12 2 2
27 12 1 0 13 9 9 1 0 9 2 12 2 2 10 0 9 9 9 2 15 15 13 9 1 0 9 2
3 2 11 2
3 0 9 9
1 9
36 9 2 0 0 9 0 9 2 11 2 12 2 13 0 9 9 11 1 11 2 0 9 0 0 9 2 11 11 2 11 11 2 11 11 2 2
20 10 9 1 0 9 3 14 3 0 9 0 9 13 1 0 9 1 0 9 2
36 1 0 9 13 2 16 9 0 9 13 13 9 14 9 0 9 2 7 7 0 9 2 0 1 9 13 15 3 1 9 3 0 9 3 13 2
30 0 9 0 0 9 11 11 2 3 0 11 11 2 1 0 9 11 2 0 11 11 2 13 0 9 1 9 7 9 2
17 15 13 1 0 9 0 9 0 9 0 9 1 9 7 1 9 2
8 7 11 1 11 9 9 13 2
17 0 9 0 9 13 9 13 9 16 3 0 9 3 0 0 9 2
44 3 0 0 9 13 12 9 2 16 11 0 9 13 9 13 1 9 9 0 0 9 2 13 9 9 1 0 0 9 7 13 9 1 9 0 9 2 0 15 1 9 0 9 2
19 12 0 0 9 13 9 0 9 2 15 15 9 13 1 9 7 1 9 2
33 0 0 9 2 1 9 0 9 0 0 3 2 3 13 2 15 9 0 9 11 2 0 2 16 15 13 2 13 1 0 9 9 2
26 1 0 15 9 2 3 0 1 9 2 13 13 0 9 14 9 2 15 3 13 9 2 9 7 9 2
17 0 11 13 14 9 0 11 2 3 0 1 0 9 1 0 9 2
26 0 9 9 3 0 9 9 2 9 7 9 1 0 9 13 1 15 2 15 15 13 7 15 4 13 2
18 1 0 0 9 3 3 9 9 1 9 0 9 13 3 15 0 9 2
2 11 11
7 0 9 2 11 2 12 2
9 9 1 11 2 11 2 9 9 2
16 9 2 11 1 11 2 9 2 11 11 2 9 2 11 11 2
13 13 2 11 11 2 11 11 2 11 11 7 0 2
4 0 9 1 11
1 9
31 9 2 1 9 9 1 9 0 9 15 9 1 0 9 9 13 13 3 12 9 0 9 11 7 11 2 15 13 11 11 2
16 1 0 9 9 15 3 4 0 9 13 3 1 12 2 9 2
37 11 2 11 2 11 2 11 7 0 9 0 9 13 1 0 9 3 3 9 2 3 16 1 0 11 9 2 7 9 10 9 15 13 14 1 9 2
20 9 11 1 11 7 13 16 9 2 10 0 9 15 13 13 0 1 12 9 2
25 3 0 13 7 11 11 11 2 15 10 0 3 3 13 3 1 9 9 2 3 15 3 7 13 2
14 1 10 9 15 13 1 9 2 1 9 7 3 3 2
33 0 9 0 9 7 0 9 1 9 9 13 3 1 15 0 2 1 15 0 9 1 15 13 1 10 0 9 7 3 14 0 9 2
38 0 9 1 9 13 3 11 11 1 9 3 0 11 2 11 11 16 3 0 11 7 10 0 2 3 0 9 2 10 0 9 13 0 9 9 7 9 2
29 1 9 1 15 13 3 0 0 9 7 3 0 2 14 0 9 3 0 9 0 9 2 15 13 1 9 3 0 2
40 10 9 13 2 1 0 9 11 11 1 9 11 2 7 9 1 9 2 15 4 15 3 1 9 9 13 13 7 15 4 15 0 7 0 9 9 11 11 13 2
27 9 2 15 13 0 9 2 15 13 7 1 0 9 7 13 3 3 0 2 7 14 3 3 0 9 9 2
49 9 1 3 0 9 11 11 2 11 2 15 1 9 1 3 0 0 9 13 1 0 9 9 7 3 16 9 1 9 1 11 13 9 9 7 13 0 9 0 9 0 9 2 1 15 3 13 3 2
2 11 11
14 9 11 2 11 7 0 2 0 2 0 2 0 2 2
7 11 11 2 11 7 11 2
4 9 11 11 2
28 9 11 11 2 9 11 11 2 9 11 11 2 9 11 11 2 9 11 11 2 9 11 11 2 9 11 11 2
12 9 0 9 2 12 2 9 2 12 2 9 2
4 16 4 15 13
1 9
2 11 11
19 16 0 9 3 13 10 0 9 0 9 2 9 9 10 9 13 3 0 2
18 0 9 15 13 3 12 9 2 16 1 9 3 13 0 0 0 9 2
27 7 3 1 9 9 2 3 10 0 9 2 9 0 2 15 4 13 10 9 13 1 9 0 0 0 9 2
37 1 9 0 9 13 1 11 0 9 0 11 2 9 2 2 15 3 7 3 2 1 12 2 13 1 11 1 9 1 11 2 16 4 15 13 2 2
23 3 15 9 0 0 0 9 13 1 0 11 1 9 12 1 0 9 0 0 9 1 11 2
37 9 11 13 9 3 2 16 15 13 1 15 2 16 4 0 9 2 7 1 9 0 2 11 0 11 2 9 9 2 2 13 1 9 12 1 15 2
24 13 15 3 2 16 14 9 9 1 0 9 2 7 3 15 9 13 1 10 9 0 7 0 2
40 1 12 9 9 13 9 12 9 2 15 15 10 0 9 7 9 9 1 0 9 0 9 13 9 9 7 0 9 2 15 13 3 11 11 2 0 9 11 11 2
32 9 13 11 0 11 2 9 0 9 1 9 1 11 2 1 2 11 2 3 3 0 11 13 2 1 0 9 3 13 3 2 2
21 9 1 9 1 12 1 12 9 15 13 1 9 1 0 11 13 1 0 0 9 2
32 13 1 0 9 2 7 3 13 0 2 3 0 9 1 9 2 1 15 13 2 1 15 15 13 9 9 2 0 7 0 9 2
18 1 9 2 1 15 1 15 13 3 2 15 11 13 1 9 0 9 2
32 1 3 3 0 9 2 9 9 7 0 9 2 13 14 12 9 9 2 0 1 9 9 11 2 0 11 2 11 7 11 11 2
16 9 0 7 0 0 9 13 13 7 16 0 9 0 0 9 2
4 11 13 0 9
12 3 0 9 13 1 9 9 12 9 9 11 2
22 1 9 9 12 9 15 13 0 9 2 7 15 1 0 9 13 13 9 0 0 9 2
9 0 9 11 13 12 2 9 12 2
22 10 9 13 1 9 12 2 9 2 3 15 9 10 9 1 9 13 3 1 0 9 2
33 0 9 9 13 12 5 9 1 0 9 2 12 5 13 9 0 9 1 0 9 9 0 2 9 2 11 2 0 12 9 13 11 2
32 11 13 16 0 2 0 7 3 0 9 2 7 15 3 1 9 0 9 7 9 1 9 2 9 7 9 0 9 1 10 9 2
14 1 10 0 9 13 11 2 0 0 9 7 11 11 2
17 9 15 13 1 12 9 2 16 3 16 9 9 11 13 9 9 2
22 3 13 15 9 9 2 0 9 2 9 2 9 9 3 0 9 2 0 7 9 9 2
26 1 9 10 9 2 7 2 1 9 12 2 10 9 13 7 13 12 9 0 9 1 0 9 0 9 2
8 13 15 7 1 9 0 9 2
21 1 9 9 12 13 9 3 13 1 9 7 9 9 9 9 1 9 9 11 12 2
9 0 9 13 13 1 0 9 9 2
17 1 9 12 4 13 0 9 9 7 1 9 3 13 9 0 9 2
15 0 9 0 9 9 13 1 9 9 12 1 12 9 9 2
7 9 0 9 13 0 9 2
17 1 0 9 13 9 9 11 0 9 12 9 2 0 3 12 9 2
10 1 0 9 15 13 1 9 12 9 2
15 0 9 13 1 9 9 11 1 10 0 2 9 12 9 2
3 2 11 2
14 0 9 9 0 0 11 13 9 11 11 7 9 11 11
3 9 11 11
8 11 13 0 9 9 0 0 11
33 1 1 9 0 0 9 15 13 0 2 3 3 0 9 0 0 11 1 0 0 9 2 15 1 9 13 1 0 9 11 1 11 2
36 7 13 0 0 11 1 0 0 9 0 9 0 0 11 2 1 15 15 1 0 11 1 15 13 7 0 9 0 11 7 0 9 7 9 11 2
11 11 1 11 3 13 1 0 9 0 9 2
34 1 3 0 9 13 12 0 9 2 15 13 9 9 2 9 7 0 0 9 3 3 16 0 0 9 2 0 9 0 9 7 0 9 2
30 16 4 15 13 1 0 9 13 2 16 15 13 1 0 9 0 9 2 9 9 0 0 11 13 3 2 3 7 3 2
3 2 11 2
16 11 11 2 11 11 2 0 9 1 11 1 11 2 11 2 12
2 9 9
5 3 13 1 9 2
2 11 11
17 9 2 0 2 12 2 13 9 9 2 13 1 9 9 9 9 9
28 9 0 9 0 1 0 9 1 0 0 9 15 13 13 9 0 3 1 9 2 9 7 9 16 1 9 9 2
27 1 9 0 9 2 0 9 1 11 1 11 1 0 0 9 1 11 15 7 3 13 1 15 15 3 0 2
16 13 15 3 9 11 11 11 2 11 11 11 7 11 11 11 2
16 1 0 9 7 0 11 9 13 0 9 0 9 1 0 9 2
24 1 9 12 13 11 14 12 9 2 10 9 13 1 9 0 9 0 9 1 11 7 1 9 2
16 0 13 9 9 2 9 2 7 0 9 2 12 9 0 2 2
8 9 9 7 9 13 1 9 2
60 16 4 15 9 3 13 0 9 0 9 2 9 2 9 2 9 2 2 16 4 15 3 13 0 0 9 1 9 1 10 0 9 2 7 16 4 15 9 10 9 13 3 13 1 9 2 9 7 1 0 9 2 1 15 15 3 13 0 9 2
26 1 0 9 7 1 0 0 2 0 9 9 11 2 13 15 1 9 9 2 15 1 15 13 15 0 2
19 12 9 15 1 9 13 0 9 2 12 3 0 9 1 9 7 0 9 2
23 13 0 0 9 1 10 0 0 9 2 0 9 1 0 9 7 9 7 1 9 0 9 2
11 0 9 9 3 13 1 9 3 11 11 2
13 0 9 0 9 15 1 15 13 1 0 0 9 2
26 11 11 7 3 3 0 11 11 15 1 3 0 9 10 9 13 0 0 0 9 1 9 9 1 11 2
28 1 9 13 10 9 1 0 11 3 14 3 0 2 7 1 0 9 15 3 16 9 13 1 9 9 11 12 2
18 1 10 0 9 16 9 11 2 11 13 9 1 10 9 11 11 11 2
16 9 0 9 1 0 9 13 9 0 9 11 11 7 11 11 2
21 10 0 0 9 1 9 9 3 13 2 7 1 15 13 0 9 1 0 9 9 2
10 0 9 2 0 9 1 11 1 11 2
14 0 0 9 1 11 2 12 2 9 2 12 2 9 2
2 11 11
2 9 9
4 9 7 9 9
2 11 11
16 9 2 0 2 12 2 13 0 9 7 9 2 13 1 0 9
3 9 11 11
26 9 16 1 0 9 2 9 9 2 9 2 9 2 0 9 2 9 3 1 9 0 2 3 1 0 2
49 7 3 10 12 9 13 1 15 9 11 11 15 0 1 9 0 9 0 9 2 9 0 15 1 0 9 1 0 9 9 2 7 0 3 13 3 3 0 9 2 16 1 15 13 10 0 9 13 2
11 9 1 9 1 9 2 9 1 10 9 2
32 15 15 2 3 1 3 0 9 1 9 9 7 9 2 11 11 13 1 0 9 9 15 13 2 15 0 9 13 1 9 11 2
28 0 9 2 3 0 1 10 9 0 7 0 2 7 3 13 3 0 9 0 9 2 0 9 10 9 1 9 2
31 13 15 15 2 1 11 9 1 9 7 9 2 9 7 0 9 2 15 15 3 13 0 9 2 7 3 7 9 0 9 2
34 11 11 15 13 12 2 9 12 1 11 2 15 13 3 11 2 3 2 16 15 15 13 2 15 13 10 9 7 15 2 2 2 2 2
18 13 1 0 9 1 11 2 3 13 3 9 10 0 9 1 9 2 2
14 3 13 0 9 1 11 7 0 11 2 9 12 2 2
27 1 9 12 2 12 13 9 0 9 0 9 2 1 9 12 13 0 9 1 11 16 9 9 11 2 11 2
32 0 9 15 13 3 1 9 12 2 11 1 15 13 0 9 2 2 2 3 13 1 11 1 11 7 13 16 9 1 0 9 2
19 1 9 11 15 13 1 11 2 3 15 1 11 13 1 0 9 1 11 2
17 1 9 12 13 1 0 9 13 1 0 9 7 13 15 9 11 2
8 1 9 12 13 1 9 9 2
37 1 9 12 13 1 11 2 13 4 13 2 16 9 13 9 2 15 13 13 7 1 0 9 9 2 2 2 2 7 0 9 3 13 16 0 9 2
9 9 12 15 13 1 9 1 11 2
10 13 16 0 9 2 9 7 16 9 2
20 1 9 12 2 12 13 9 1 0 0 0 11 1 11 2 0 9 3 13 2
20 3 2 16 15 9 12 13 1 11 2 13 16 9 0 9 14 1 9 12 2
20 10 0 9 13 3 1 11 2 11 7 0 9 2 1 9 12 3 7 3 2
16 9 11 2 9 12 9 2 15 13 0 9 3 7 3 3 2
30 3 1 9 10 9 2 9 2 12 2 2 3 1 9 12 2 1 9 1 11 2 3 2 3 13 2 13 0 9 2
22 7 3 1 9 12 2 9 9 7 9 2 2 3 15 3 13 0 9 1 0 9 2
24 0 9 1 0 9 3 3 9 13 2 9 11 7 0 9 9 4 1 9 0 9 13 2 2
42 3 1 9 12 2 1 10 0 9 2 13 0 9 1 0 9 15 0 2 0 9 2 1 15 4 13 10 9 2 9 2 9 2 9 1 9 7 9 7 9 9 2
53 16 3 9 13 3 0 9 15 2 15 1 0 9 13 2 15 13 14 10 9 2 15 13 0 15 13 2 7 15 9 13 1 15 0 9 7 13 15 1 9 3 16 9 0 2 0 1 9 10 9 2 0 2
9 11 11 15 13 9 0 7 0 2
26 0 3 0 7 0 9 10 9 2 15 13 9 13 1 15 2 16 4 15 13 1 10 0 0 9 2
16 7 0 3 1 15 2 15 15 10 9 13 2 13 3 3 2
19 0 9 2 3 1 10 0 9 2 13 9 0 9 7 3 0 9 9 2
59 1 10 9 7 9 13 7 0 9 2 1 9 2 3 13 13 1 0 2 3 0 9 2 16 7 1 0 9 2 10 10 9 15 13 0 9 2 2 13 14 9 1 9 9 2 9 2 15 15 13 0 9 7 9 2 9 7 9 2
34 9 13 3 2 3 3 15 13 13 1 10 9 2 1 15 2 15 3 13 1 15 0 2 9 9 2 10 0 0 9 0 1 15 2
12 7 11 13 13 7 10 0 9 0 7 0 2
28 0 13 2 16 1 0 9 13 1 9 11 11 2 3 1 9 0 0 2 13 2 0 10 0 9 1 15 2
23 9 3 13 2 16 13 4 11 13 1 9 9 0 2 16 13 3 11 11 7 11 11 2
13 9 0 9 13 3 9 16 9 3 7 3 0 2
34 9 14 2 7 16 9 2 15 15 13 0 13 3 3 2 1 0 7 0 9 9 2 3 9 0 1 0 9 9 3 0 10 9 2
35 7 14 10 9 13 15 0 10 9 1 9 2 15 13 13 9 0 9 7 0 9 2 1 9 9 2 9 2 9 7 9 1 10 9 2
13 7 1 15 13 11 3 9 9 0 16 10 0 2
34 1 0 0 9 13 13 9 0 0 9 2 0 9 9 2 2 2 15 13 7 0 9 7 10 0 9 2 0 0 9 2 9 2 2
65 9 0 9 2 15 3 13 0 0 9 2 0 9 2 2 16 7 0 9 2 15 9 2 15 4 13 2 2 1 9 9 13 2 2 7 0 9 1 0 9 9 2 3 1 9 7 9 2 9 9 7 9 13 1 11 1 15 0 2 15 13 11 7 11 2
20 1 0 9 13 9 7 10 9 2 9 2 15 3 13 10 9 2 0 15 2
16 3 9 2 2 9 2 1 15 9 7 9 3 3 12 13 2
13 9 9 16 3 0 9 13 11 1 9 1 9 2
27 7 15 2 9 2 0 0 9 2 15 13 9 15 9 7 9 15 9 7 9 2 2 15 9 0 9 2
35 1 0 9 9 2 15 15 3 3 13 15 2 3 2 1 0 9 2 15 13 13 11 2 11 2 11 7 10 9 0 9 0 1 9 2
38 11 13 2 3 1 3 0 11 2 11 11 2 11 11 7 11 11 0 9 2 1 9 0 0 9 2 7 15 3 9 10 9 2 7 7 9 9 2
27 9 1 15 13 3 9 15 0 2 9 7 9 1 10 7 15 2 7 14 14 9 2 3 0 7 0 2
26 7 3 10 9 2 14 2 0 2 16 0 2 13 0 7 0 9 15 2 15 13 1 0 9 9 2
10 15 9 0 7 0 13 16 0 9 2
1 9
30 1 9 11 11 1 9 9 13 9 0 9 11 2 9 0 9 2 11 2 7 9 9 11 2 11 2 11 2 11 2
29 13 1 9 1 9 9 2 3 15 1 9 9 9 9 7 9 3 7 3 3 1 11 13 0 0 13 0 9 2
29 9 9 1 12 2 7 0 0 9 13 1 12 2 9 1 9 1 9 11 7 1 0 9 11 1 0 0 9 2
4 0 9 9 3
18 0 9 0 7 0 1 11 13 1 10 9 3 0 0 0 9 9 2
29 1 12 2 9 1 12 2 9 3 13 9 7 0 9 1 0 9 9 7 13 9 0 15 9 0 9 9 11 2
33 1 9 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 13 3 13 9 2 3 11 11 2 11 11 2 11 11 2
12 9 4 13 9 9 2 15 13 12 2 9 2
9 1 9 0 9 4 3 13 9 2
3 2 11 2
3 1 0 9
18 9 9 12 2 12 2 9 11 11 2 12 9 2 9 12 9 2 2
19 9 0 9 9 9 2 13 3 3 2 13 0 9 9 0 1 0 9 2
14 1 9 9 13 9 0 9 11 11 2 9 0 9 2
15 1 9 13 9 11 11 2 15 3 13 3 1 0 9 2
12 1 11 11 2 9 0 9 2 13 11 11 2
21 1 0 9 9 13 1 0 9 1 15 2 1 10 0 9 15 13 1 10 9 2
8 13 7 9 1 9 0 9 2
3 2 11 2
18 0 9 1 11 13 1 0 9 9 2 9 7 9 0 7 0 9 2
24 3 3 0 9 13 10 0 9 2 1 15 3 13 7 0 9 9 11 11 2 1 9 2 2
26 1 10 9 0 13 3 11 7 11 0 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2
10 9 13 13 3 1 12 1 12 9 2
3 2 11 2
5 9 11 11 2 11
5 9 9 1 12 9
2 11 11
13 1 9 0 0 9 9 9 13 12 0 0 9 2
22 15 0 4 3 3 13 1 9 2 15 13 1 0 11 1 9 12 1 9 11 12 2
12 1 0 0 0 9 13 9 9 3 3 3 2
50 13 0 2 16 0 0 7 0 9 11 0 2 11 0 7 0 11 11 15 1 9 9 11 11 3 13 1 9 0 15 0 9 0 9 0 9 2 1 9 0 9 3 13 0 9 0 9 1 15 2
40 9 0 3 7 3 0 11 13 3 10 0 0 9 2 3 0 1 9 0 9 2 16 3 0 0 9 2 0 15 1 3 3 0 9 3 0 9 0 9 2
22 1 9 0 9 11 0 7 12 0 9 7 0 9 13 7 9 3 0 9 11 11 2
16 0 9 13 3 0 9 0 0 9 11 0 1 9 0 9 2
31 0 9 13 13 1 3 0 9 0 2 7 3 2 9 9 1 9 1 10 0 9 7 0 0 9 13 3 3 7 3 2
27 0 13 1 0 9 3 9 9 2 7 15 3 3 2 3 15 9 9 13 1 0 0 9 1 0 9 2
24 0 9 0 9 2 15 13 14 1 9 2 13 1 0 2 0 9 7 10 9 0 0 9 2
12 9 9 2 11 0 2 11 0 2 11 11 2
10 9 15 0 2 11 2 12 2 9 2
6 9 9 2 11 0 2
10 9 15 0 2 11 2 12 2 9 2
1 9
3 1 0 9
19 3 0 9 11 7 10 9 11 15 13 2 16 3 4 13 1 9 9 2
30 12 13 0 9 1 9 9 2 15 1 15 13 9 0 9 7 9 2 15 13 9 2 16 13 10 9 1 0 9 2
17 1 15 15 13 10 9 14 1 9 2 16 11 13 3 3 13 2
23 1 10 9 4 1 0 9 0 9 7 9 9 7 9 3 13 3 0 9 11 2 2 2
25 0 2 3 0 9 13 1 9 11 11 7 13 2 7 1 3 0 9 2 1 0 9 10 9 2
30 13 3 3 0 9 9 2 9 7 9 2 9 13 13 1 3 0 9 2 0 1 0 9 1 11 2 7 0 9 2
22 16 1 9 13 3 0 9 2 0 9 13 3 1 10 3 0 2 0 7 0 9 2
33 15 3 13 0 0 9 2 15 13 0 2 0 9 0 9 11 7 0 9 1 0 9 11 2 1 3 0 7 0 0 9 2 2
3 2 11 2
7 0 11 2 11 2 12 2
8 9 1 11 2 0 0 11 2
5 9 2 11 11 2
13 13 2 11 11 2 11 11 2 11 11 7 0 2
3 0 11 3
3 1 0 9
36 1 0 0 11 4 0 0 9 0 11 2 10 9 9 0 13 0 15 2 3 3 13 2 14 15 2 15 13 1 0 9 0 9 0 9 2
13 7 0 9 1 10 0 9 1 0 11 13 3 2
31 9 1 12 0 9 13 3 1 9 2 15 15 1 0 9 13 3 16 3 0 9 0 12 2 11 11 2 11 7 11 2
22 0 2 0 0 9 1 15 13 9 0 0 12 2 7 7 3 0 9 7 0 9 2
28 9 3 0 9 13 0 2 0 2 0 9 2 0 0 9 0 9 11 11 2 11 2 14 0 7 11 2 2
39 10 0 9 15 13 1 0 9 11 11 2 11 2 0 2 2 0 9 11 11 1 11 2 15 15 13 2 7 9 11 11 1 0 11 2 0 3 2 2
26 9 9 9 13 3 0 2 0 11 2 15 1 0 9 7 1 10 9 1 9 13 16 0 15 9 2
17 9 1 0 11 13 0 9 2 3 13 0 9 13 3 0 9 2
3 2 11 2
6 0 11 3 2 12 2
6 9 1 11 2 11 2
1 3
30 9 9 11 11 2 0 9 0 9 2 1 0 9 0 9 1 0 0 9 2 12 2 12 15 13 1 12 2 9 2
17 9 0 9 11 2 2 2 4 3 3 13 1 0 9 0 9 2
21 13 2 1 12 2 9 2 0 9 11 11 2 9 2 7 11 11 2 9 2 2
15 9 9 7 0 9 13 3 0 9 1 9 9 11 3 2
22 15 15 13 14 15 13 2 7 15 13 2 2 2 13 3 1 0 9 9 11 11 2
6 0 9 3 1 12 9
29 9 1 0 9 12 2 10 9 13 0 9 2 13 13 9 11 9 2 15 13 0 9 0 9 9 2 9 9 2
21 1 1 15 2 16 1 0 9 4 13 0 9 2 13 9 1 9 9 1 11 2
19 15 1 0 9 13 1 0 9 2 16 1 9 1 9 13 12 9 9 2
26 10 9 2 15 13 4 13 1 9 0 9 2 13 9 1 11 13 1 9 9 9 3 1 9 9 2
31 1 9 4 1 9 13 4 13 0 9 2 0 1 9 0 0 9 7 9 2 0 9 15 3 13 13 9 0 0 9 2
23 1 0 9 9 1 11 4 3 13 13 9 1 11 2 11 2 11 2 11 2 11 3 2
25 1 9 9 11 11 13 0 9 1 15 2 16 9 9 7 0 9 4 13 4 13 1 12 9 2
15 1 10 9 13 9 10 9 0 1 10 9 9 0 11 2
28 1 10 9 15 1 11 1 9 9 7 9 3 13 0 9 11 1 9 9 0 9 11 11 11 7 0 9 2
3 2 11 2
3 11 3 13
5 11 2 11 2 2
40 0 9 3 13 2 16 13 0 9 2 16 4 15 13 13 0 9 9 1 0 9 7 1 0 0 9 2 15 4 13 1 9 12 2 12 2 1 0 9 2
12 0 9 4 1 0 9 13 1 12 2 12 2
32 0 2 15 15 15 13 2 7 4 3 13 2 16 13 1 0 9 13 9 15 7 13 15 3 9 7 1 9 1 12 9 2
6 2 3 1 9 9 2
2 9 9
24 13 15 10 10 9 2 15 1 9 12 2 12 2 1 9 7 16 9 13 0 9 0 9 2
18 10 9 1 9 7 9 4 13 9 1 9 9 1 0 9 0 9 2
28 1 9 2 16 4 9 0 9 13 1 10 9 2 7 13 2 14 15 0 2 13 15 13 1 9 1 15 2
15 9 13 2 16 4 9 0 11 13 1 10 0 9 11 2
26 1 9 2 16 13 2 13 15 1 0 9 9 2 2 12 2 12 12 12 2 3 13 13 15 13 2
3 13 1 9
7 1 9 9 2 12 4 13
7 11 2 11 2 11 2 2
18 9 9 2 9 2 9 9 7 9 11 11 15 3 13 1 9 9 2
9 13 15 1 9 9 9 2 12 2
24 9 11 11 11 11 13 2 16 9 9 2 12 16 0 9 13 1 9 0 9 1 9 9 2
19 9 7 13 9 1 9 9 2 15 13 13 9 1 9 13 9 9 9 2
9 3 1 9 12 2 0 9 13 0
13 9 0 0 9 11 11 11 11 1 0 0 9 2
27 3 2 16 4 1 0 11 13 9 0 9 2 13 11 0 0 9 2 16 4 13 9 11 7 13 9 2
2 9 11
6 0 9 13 1 0 9
5 11 2 11 2 2
23 9 0 9 0 9 1 9 0 9 13 1 9 9 0 9 2 11 2 11 11 3 0 2
9 0 9 1 9 0 9 4 13 2
27 0 9 0 9 1 0 9 2 15 7 13 3 9 1 9 12 9 1 15 2 10 9 4 0 9 13 2
22 1 0 9 13 13 10 9 2 16 4 15 10 9 3 13 2 13 3 11 1 11 2
13 3 13 2 16 0 9 4 13 12 7 12 9 2
5 11 1 9 4 13
2 11 2
20 0 0 9 2 11 2 13 1 9 2 15 4 13 13 0 9 1 0 11 2
15 1 0 9 1 11 15 3 13 9 9 11 11 11 11 2
19 9 0 9 11 13 1 9 9 9 2 1 15 13 1 9 3 1 11 2
12 1 9 15 13 0 0 9 9 1 9 11 2
12 11 3 13 9 0 9 1 0 9 1 11 2
10 11 4 1 15 13 3 13 9 9 2
18 1 9 1 11 13 3 3 0 9 11 11 1 0 9 9 11 11 2
14 11 1 9 13 2 16 11 0 9 1 0 11 13 2
6 0 9 13 1 9 11
2 11 2
15 0 0 9 11 9 2 12 15 3 13 1 0 9 11 2
33 13 1 0 9 1 12 0 2 15 13 0 0 9 2 16 11 9 2 12 13 1 0 9 3 0 9 7 9 1 0 0 9 2
24 1 9 1 0 9 15 3 0 9 13 1 0 9 2 7 13 15 9 9 9 11 11 11 2
27 9 1 0 9 13 1 9 1 9 0 9 2 16 12 0 9 1 9 13 9 9 0 9 1 0 9 2
16 9 11 13 1 0 9 3 0 9 7 3 3 13 1 9 2
15 3 1 9 12 2 11 9 2 12 2 3 7 1 0 9
8 11 2 11 2 11 13 9 11
4 11 11 2 11
24 0 9 9 9 11 2 11 3 13 9 0 9 11 11 10 0 9 1 12 9 0 0 9 2
27 1 10 9 13 10 9 16 1 9 9 7 9 9 2 7 7 1 9 9 0 9 1 0 9 10 9 2
13 1 11 15 11 2 11 13 1 0 9 11 11 2
18 9 15 1 9 9 0 9 7 0 9 13 3 0 0 2 0 9 2
15 13 0 9 11 2 15 13 1 9 0 9 2 13 11 2
13 13 2 16 11 13 9 11 1 9 1 0 9 2
27 9 11 11 1 9 1 0 9 13 2 16 9 0 9 13 11 3 7 3 13 11 7 13 9 10 9 2
32 1 9 11 2 16 15 13 9 0 9 1 10 9 2 13 2 16 13 9 1 11 7 13 15 13 9 11 2 10 9 13 2
3 1 0 9
5 11 11 2 11 11
25 10 9 13 13 9 2 16 9 13 0 9 3 2 3 4 15 13 13 2 15 13 1 0 9 2
17 3 3 13 3 2 16 3 1 10 9 9 9 3 13 0 9 2
17 9 15 13 2 16 15 13 0 9 10 9 7 13 9 11 11 2
18 13 9 1 15 2 16 15 2 15 9 13 2 13 1 10 9 9 2
20 9 9 13 7 12 9 2 1 9 1 0 0 9 13 0 9 10 9 9 2
7 9 3 13 0 9 11 2
9 10 0 9 13 0 7 0 9 2
10 1 15 13 0 0 9 3 0 9 2
23 1 0 9 9 13 9 9 9 9 11 11 11 2 9 9 9 11 11 7 0 0 9 2
30 16 13 9 1 0 9 3 3 3 0 1 0 9 2 3 1 11 2 2 13 15 3 13 10 10 9 1 0 9 2
14 9 9 13 9 1 9 7 10 9 1 0 9 13 2
12 0 9 1 0 9 9 1 0 9 13 0 2
13 0 9 4 13 2 16 10 9 9 9 13 13 2
21 13 15 3 9 2 16 3 4 13 13 9 9 0 9 2 16 15 13 14 3 2
5 7 13 7 3 2
13 9 9 1 0 9 9 0 9 9 3 13 13 2
7 0 9 13 0 9 9 2
43 3 3 15 13 9 2 16 0 9 4 13 9 2 10 9 13 0 0 9 1 0 0 9 7 10 0 9 13 0 9 1 11 11 7 3 0 9 1 10 9 1 11 2
13 1 0 9 3 1 10 9 13 9 1 10 9 2
25 11 4 3 13 2 16 15 1 0 9 7 0 9 10 9 11 11 3 13 2 16 11 13 9 2
9 0 9 7 13 3 1 10 9 2
19 13 3 3 2 16 0 9 1 0 7 0 9 13 9 9 1 10 9 2
14 16 4 13 1 9 0 2 1 15 0 4 13 13 2
11 9 0 9 3 13 1 3 0 9 9 2
7 1 15 10 11 3 13 2
5 9 1 9 11 13
5 11 2 11 2 2
20 9 9 0 9 1 11 13 1 9 0 9 2 13 3 1 9 11 9 11 2
15 0 9 13 1 9 0 9 0 9 1 9 1 0 11 2
35 1 9 9 0 9 1 9 9 1 9 9 11 13 2 16 7 16 1 11 13 9 1 9 1 9 0 9 2 9 9 1 0 9 13 2
11 15 13 1 9 12 9 9 2 0 9 2
5 11 13 11 1 9
5 11 2 11 2 2
22 1 3 0 0 9 1 9 0 9 1 0 0 9 13 9 11 11 9 11 11 11 2
24 1 0 0 9 13 0 9 7 9 9 0 9 11 2 1 15 1 9 13 1 0 9 11 2
32 11 11 15 13 1 0 9 0 2 16 9 11 11 15 13 9 1 10 0 9 3 15 7 16 15 13 2 3 13 1 9 2
28 13 9 2 3 4 0 9 11 11 3 2 16 13 11 7 11 1 9 2 16 4 1 15 3 13 2 13 2
32 1 0 9 15 3 13 2 16 9 1 12 9 1 9 1 9 13 2 7 13 2 16 4 4 0 9 1 9 1 15 13 2
21 9 11 13 3 1 9 2 10 0 9 7 11 0 9 10 9 1 9 3 13 2
1 3
20 0 9 1 11 1 11 2 1 15 13 9 0 9 11 2 4 3 13 9 2
17 0 9 9 4 13 1 15 9 1 12 2 12 1 12 2 12 2
38 16 9 9 11 7 11 1 11 13 1 0 9 1 11 9 1 9 0 0 9 2 15 1 0 9 1 10 9 4 12 2 12 2 13 13 1 9 2
8 13 15 9 9 11 2 11 2
19 13 15 9 9 11 2 16 12 2 12 2 4 1 9 13 12 0 9 2
5 0 9 13 9 9
5 11 2 11 2 2
17 9 9 9 9 1 12 9 13 9 9 1 12 2 9 0 9 2
9 3 1 0 9 15 13 3 12 2
30 9 9 7 0 9 11 11 3 3 13 2 16 1 9 0 9 1 9 13 1 10 9 3 1 12 2 9 12 9 2
24 9 4 3 13 1 9 7 13 2 14 13 2 7 4 9 1 15 13 2 13 9 11 11 2
26 13 2 16 1 9 9 10 0 9 1 12 2 9 0 9 13 9 1 10 9 3 1 12 9 9 2
4 0 9 1 9
2 11 2
41 0 9 1 9 1 11 13 2 16 4 1 0 9 0 0 9 9 0 9 1 9 7 9 13 7 9 2 16 9 4 1 10 9 13 4 13 16 9 0 9 2
15 0 0 9 2 11 2 9 10 9 11 11 13 0 9 2
22 1 9 1 0 9 7 9 0 9 7 9 0 1 11 13 16 0 9 0 9 9 2
12 13 1 9 0 9 11 7 1 10 0 9 2
25 0 13 1 0 9 7 9 9 0 9 2 7 1 9 13 1 10 9 13 0 9 2 13 11 2
24 3 4 1 9 11 1 0 9 13 1 12 12 0 9 2 7 15 13 9 1 0 10 9 2
4 9 13 3 9
5 11 2 11 2 2
17 12 9 13 0 2 16 13 1 11 12 9 7 13 3 9 9 2
13 13 15 3 9 9 0 2 9 2 11 9 11 2
21 9 0 9 13 12 9 9 9 2 3 1 9 9 13 9 7 13 12 12 9 2
20 0 9 13 9 0 9 7 13 2 16 0 13 12 9 1 0 0 0 9 2
15 12 7 4 1 9 1 9 9 3 1 9 13 1 9 2
4 0 9 4 13
5 11 2 11 2 2
28 16 9 0 0 9 9 0 9 9 11 11 2 13 2 16 4 15 13 0 9 2 10 9 13 0 9 9 2
29 11 11 1 9 9 9 3 13 11 2 16 10 9 1 9 13 9 9 7 11 11 2 4 13 1 9 1 9 2
29 9 0 9 0 9 11 2 11 2 1 9 3 13 2 16 15 13 13 3 12 7 9 9 9 1 12 0 9 2
15 1 9 11 13 9 0 7 0 13 1 9 13 1 9 2
29 11 11 2 1 9 13 2 16 15 10 0 9 13 7 13 9 10 0 9 1 11 3 1 0 9 9 9 9 2
23 11 2 11 11 13 2 16 10 9 3 13 9 2 15 9 3 3 13 1 0 0 9 2
25 11 11 2 13 1 9 2 16 13 1 15 2 16 9 13 0 2 10 9 15 14 9 13 9 2
5 0 9 13 0 9
5 11 2 11 2 2
10 0 9 1 9 4 13 3 12 9 2
15 9 1 9 0 9 13 9 9 10 9 1 15 9 9 2
28 9 2 15 3 13 2 13 3 0 9 1 10 9 2 7 9 9 13 3 13 9 7 9 9 13 7 13 2
16 1 9 4 13 3 0 13 1 0 9 1 9 16 1 9 2
28 1 0 9 15 3 13 1 9 0 9 2 3 1 0 9 2 15 15 13 13 1 0 9 13 1 9 11 2
23 9 4 13 0 9 1 15 2 7 1 9 10 9 1 9 9 7 9 0 0 9 9 2
21 1 9 15 13 7 1 0 9 11 2 7 15 1 9 1 0 9 7 0 9 2
17 0 9 9 1 10 9 0 0 0 9 13 0 9 1 0 9 2
19 9 1 9 0 9 4 14 13 9 11 2 7 13 4 3 13 9 9 2
14 16 4 13 15 2 3 4 13 0 2 13 9 0 9
5 11 2 11 2 2
25 9 0 0 9 11 11 13 13 9 1 9 1 15 2 15 13 9 1 3 0 9 10 0 9 2
26 16 4 13 10 7 15 9 2 1 0 9 4 15 13 3 13 2 16 4 1 15 13 3 0 9 2
38 3 3 2 16 4 15 0 9 13 2 13 9 0 9 1 10 9 0 9 2 15 1 0 12 9 13 1 12 9 12 7 3 13 9 7 10 9 2
28 16 3 3 2 16 13 1 3 0 9 2 13 15 1 9 9 0 9 9 15 2 15 13 7 13 15 13 2
23 15 13 9 2 3 3 4 13 9 1 9 2 7 3 9 0 9 3 0 9 0 9 2
18 9 11 11 13 1 9 9 2 16 9 4 13 1 9 12 2 9 2
26 16 13 13 3 0 9 2 1 10 9 13 0 2 16 15 9 3 13 13 0 9 3 1 0 9 2
21 16 9 3 13 9 7 13 10 9 2 13 15 13 9 2 13 1 15 9 11 2
12 15 13 15 1 0 9 2 15 13 0 9 2
20 13 3 13 2 16 9 9 2 3 2 3 4 13 2 13 1 9 0 9 2
15 1 9 0 9 13 9 0 13 2 10 9 13 3 0 2
29 11 2 11 15 3 13 2 16 4 15 1 9 2 15 13 14 1 0 9 2 13 13 0 9 1 9 0 9 2
13 1 9 15 13 1 10 9 1 3 0 9 0 2
16 1 0 9 0 9 0 11 4 3 13 3 3 12 12 9 2
10 1 9 13 9 1 9 1 0 9 2
26 9 0 11 2 11 2 15 0 9 9 13 2 3 13 2 16 9 1 0 9 4 13 14 1 9 2
5 9 11 11 2 11
5 9 11 13 1 11
3 1 0 9
5 11 2 11 2 2
27 1 10 0 9 13 0 9 11 1 9 9 11 11 2 3 11 2 3 3 11 2 11 2 1 10 9 2
9 13 15 3 0 9 11 11 11 2
15 11 2 11 4 13 1 0 9 13 7 1 9 1 11 2
26 9 11 1 0 9 11 13 1 0 9 9 9 10 9 2 7 15 9 10 9 13 1 0 9 12 2
10 1 0 9 0 9 13 10 9 10 9
5 11 2 11 2 2
22 9 1 0 9 1 9 1 11 3 10 9 13 1 0 9 0 9 0 11 1 11 2
28 16 0 9 1 11 13 1 0 9 9 7 13 15 7 0 9 2 4 0 9 13 1 11 2 3 1 11 2
14 1 0 9 15 0 9 13 14 10 9 1 0 9 2
14 0 9 13 1 9 3 0 2 13 3 0 9 9 2
12 3 13 1 15 0 13 12 2 12 9 9 2
11 9 0 9 13 0 1 9 13 12 9 2
18 3 2 3 13 2 15 13 9 13 10 0 9 7 1 9 3 13 2
14 3 15 1 9 13 0 9 2 3 9 13 0 9 2
9 3 12 2 12 9 9 13 0 2
17 3 13 0 9 2 14 12 5 2 2 16 9 9 0 9 13 2
8 0 0 9 15 13 1 9 2
11 1 0 9 13 0 13 1 9 3 9 2
9 0 9 7 13 3 12 12 9 2
6 7 13 9 3 0 2
19 16 9 9 13 1 9 1 0 9 1 9 0 0 9 2 13 15 3 2
23 9 1 9 0 9 7 10 9 3 13 15 9 0 9 2 15 4 3 15 13 1 9 2
7 9 9 15 11 13 13 2
22 10 9 13 12 2 12 2 12 2 13 4 7 9 0 12 2 12 2 12 2 12 2
6 11 2 0 9 11 11
3 1 0 9
5 11 2 11 2 2
16 9 9 9 11 11 4 3 3 13 9 11 1 0 0 9 2
18 0 9 4 1 11 13 13 14 0 9 9 2 7 3 9 9 11 2
40 11 7 4 1 9 0 9 13 0 9 1 9 2 9 3 0 9 1 9 1 0 0 9 2 9 9 9 1 9 7 9 0 9 9 7 0 9 1 11 2
19 1 11 13 11 1 10 0 9 2 15 4 15 13 3 13 1 9 9 2
27 1 9 1 0 9 2 3 15 13 1 9 1 0 9 2 4 11 1 11 13 3 1 0 9 9 9 2
2 9 9
1 9
2 11 11
10 11 13 1 0 9 0 9 1 11 2
9 9 11 13 1 0 9 0 9 2
6 11 4 13 1 11 2
18 11 13 0 9 2 10 9 13 1 9 9 1 9 13 12 9 9 2
12 11 13 13 1 9 7 9 15 2 0 9 2
19 1 9 9 15 3 13 9 2 7 0 13 1 0 9 9 9 7 9 2
18 9 1 15 13 0 9 7 13 10 0 9 1 9 1 9 1 9 2
14 15 9 13 2 7 3 13 2 3 1 0 0 9 2
8 9 15 1 0 9 3 13 2
4 3 3 13 2
9 3 15 9 13 3 2 7 3 2
9 15 2 7 3 2 3 7 13 2
10 9 13 9 2 0 9 15 3 13 2
9 9 15 15 13 1 10 0 9 2
18 13 0 13 15 1 0 9 1 0 9 9 1 9 9 1 9 9 2
12 9 1 9 0 9 1 9 9 15 13 15 2
9 9 15 13 7 9 2 2 2 2
13 3 2 16 1 10 9 9 13 0 3 0 9 2
15 9 2 15 4 13 2 1 0 9 2 13 9 0 9 2
1 9
1 9
2 11 11
11 0 0 0 9 13 2 0 9 13 9 2
17 15 13 9 1 0 0 7 0 0 9 1 3 3 0 11 11 2
15 13 3 7 3 12 9 2 1 15 9 11 11 14 13 2
7 13 3 13 7 0 9 2
27 10 0 9 7 9 15 1 9 13 13 2 16 3 1 11 13 9 12 9 9 0 7 13 15 1 9 2
16 1 0 11 15 13 10 12 9 2 13 4 3 1 9 11 2
12 3 15 13 2 16 3 1 11 15 15 13 2
21 13 2 14 3 1 9 2 13 10 9 1 10 9 9 2 3 15 3 9 13 2
13 13 2 14 3 1 9 2 13 9 1 0 9 2
10 13 9 7 1 11 15 13 1 9 2
19 13 15 0 9 2 0 2 0 2 0 2 0 7 2 3 2 7 0 2
11 11 11 3 13 2 16 0 9 13 15 2
16 15 3 13 9 2 1 0 0 2 0 9 2 14 13 11 2
20 16 9 13 11 14 0 0 9 2 7 7 3 0 9 11 1 0 0 9 2
15 15 14 13 0 9 3 2 16 0 0 9 13 16 9 2
14 13 0 13 15 15 2 16 1 0 0 9 0 9 2
6 15 7 13 10 9 2
21 13 15 13 1 0 9 2 13 7 7 3 13 9 2 3 15 3 13 0 9 2
24 4 11 13 2 16 0 9 13 9 0 16 9 9 0 11 2 15 0 9 15 3 11 13 2
16 4 13 0 9 2 15 13 9 9 0 9 3 1 12 9 2
24 4 13 9 9 0 9 1 0 0 7 0 9 11 2 11 7 0 7 0 9 0 9 0 2
25 4 13 2 16 11 13 1 0 9 13 11 16 9 7 3 1 10 9 15 13 1 0 0 9 2
19 4 13 0 9 1 9 1 0 2 0 7 0 9 9 7 1 9 9 2
4 13 2 13 2
9 15 14 15 13 1 15 11 13 2
3 9 1 9
4 11 11 2 9
53 13 15 15 16 3 2 1 9 0 9 11 13 9 0 0 9 2 11 2 11 7 1 0 9 13 2 16 0 9 13 0 9 1 11 2 7 1 9 10 9 15 3 13 2 13 2 7 1 11 2 7 3 2
12 15 15 13 3 11 2 15 13 11 15 13 2
31 11 15 7 1 9 12 2 9 13 1 0 9 7 11 3 10 9 1 9 12 1 0 9 2 15 13 1 10 9 9 2
26 9 13 12 9 7 16 3 13 2 13 1 9 1 11 0 9 2 7 16 13 1 10 9 7 9 2
13 3 4 11 13 0 9 7 10 9 15 13 3 2
20 1 9 1 9 15 15 12 2 9 11 13 0 9 13 10 0 2 0 9 2
18 11 15 13 1 0 9 7 9 7 13 1 15 9 0 9 1 9 2
14 13 15 2 16 9 0 9 15 0 9 11 13 13 2
10 1 16 4 15 3 13 2 13 15 2
13 13 15 3 0 9 7 9 11 11 2 9 11 2
53 13 13 0 9 1 9 1 9 9 2 15 4 9 13 1 0 9 2 13 13 9 0 9 2 0 1 11 2 10 9 13 13 1 11 2 7 10 9 2 0 2 15 13 1 0 9 9 2 15 13 9 11 2
7 1 15 13 11 9 11 2
8 0 9 0 13 16 0 9 2
29 11 13 1 9 3 7 9 0 9 2 9 2 9 0 9 7 0 9 2 3 9 0 9 2 0 9 13 0 2
31 11 7 3 13 0 9 0 9 2 13 15 1 0 9 11 7 11 2 15 11 13 1 9 1 0 9 2 1 0 9 2
36 13 7 2 16 1 11 13 9 0 9 2 0 15 1 9 0 0 9 2 15 1 0 11 13 9 11 11 2 16 1 9 13 3 10 9 2
16 15 3 0 0 11 3 13 4 2 7 7 10 9 7 9 2
8 13 7 1 15 0 2 0 2
48 1 9 2 3 15 11 13 3 13 2 13 15 1 9 0 11 2 9 0 9 2 9 9 7 9 0 9 13 9 2 16 11 13 9 1 9 2 10 9 13 13 15 0 2 16 9 9 2
11 7 15 3 9 11 1 9 7 11 13 2
41 10 9 3 3 13 7 1 11 2 15 15 11 13 14 3 2 7 3 3 2 3 0 9 0 9 11 7 11 2 0 11 11 0 2 11 7 9 2 11 11 2
25 16 0 9 11 13 1 0 9 10 9 7 9 2 13 4 3 1 11 13 0 9 1 9 9 2
4 11 13 1 9
4 11 11 2 11
47 0 9 7 9 9 1 0 11 2 11 2 11 11 1 0 0 0 9 10 0 9 13 2 16 10 9 13 1 0 9 3 12 5 9 7 16 15 1 0 9 4 13 1 9 0 9 2
23 9 0 9 11 13 9 0 9 2 3 9 9 2 15 9 4 13 4 1 11 13 9 2
6 1 11 13 14 1 11
4 11 11 2 11
24 0 2 0 7 0 9 11 7 0 9 13 10 9 0 9 0 9 0 0 9 1 0 11 2
23 9 11 11 2 11 15 3 1 10 9 13 1 0 1 0 9 1 0 9 9 11 11 2
30 4 13 1 9 0 9 1 10 9 7 1 10 9 4 11 13 7 9 0 9 0 9 1 0 9 13 11 0 9 2
6 0 2 0 9 1 9
3 0 11 2
17 1 0 9 13 1 9 9 0 9 1 11 1 9 1 0 9 2
19 9 13 9 1 0 2 0 2 0 7 0 2 7 13 13 10 0 9 2
26 9 0 9 13 2 16 9 11 1 9 13 10 9 7 16 3 15 1 9 13 9 11 1 0 9 2
39 9 9 0 9 12 9 13 1 15 2 16 11 13 13 1 15 0 16 1 0 9 7 1 0 9 0 9 11 1 11 2 16 0 9 13 0 0 9 2
11 11 4 13 1 9 12 9 2 13 11 11
2 11 2
26 1 9 9 1 0 9 1 11 7 0 0 9 13 3 1 11 0 9 0 0 0 9 2 11 2 2
37 1 9 12 2 9 4 9 13 0 9 1 0 0 9 7 12 2 9 3 3 1 11 9 11 11 1 9 1 0 9 9 0 0 9 1 11 2
17 1 9 13 9 11 7 0 9 9 11 11 12 0 0 9 9 2
18 11 1 15 13 13 15 1 15 2 16 4 11 11 13 9 0 9 2
28 3 13 13 11 3 1 0 11 3 0 2 16 4 15 1 15 13 1 11 1 0 0 9 13 2 13 11 2
14 9 0 0 9 2 11 2 11 11 3 13 9 10 9
2 9 11
5 9 1 9 9 13
10 0 9 13 9 9 11 1 9 0 9
4 11 2 11 2
42 0 9 13 3 1 9 0 11 2 16 13 0 9 1 11 2 9 0 9 11 2 16 4 1 9 9 9 7 9 1 10 9 13 7 9 2 13 2 14 15 3 2
20 11 13 9 1 9 9 1 9 9 2 13 3 9 0 2 0 9 11 11 2
28 9 9 0 9 11 1 9 3 13 2 16 4 13 13 9 9 9 2 16 4 11 11 9 0 9 3 13 2
19 0 0 9 13 3 1 0 9 11 0 2 3 0 9 1 9 0 11 2
14 13 15 9 0 9 0 9 11 2 9 2 1 11 2
23 1 9 11 2 11 11 13 9 1 0 11 7 9 0 9 3 1 9 1 9 0 9 2
31 13 15 7 1 9 9 2 3 9 9 13 11 1 9 0 11 2 11 2 2 0 3 14 1 12 9 11 1 9 12 2
19 9 9 13 7 15 2 16 9 11 1 9 1 9 13 3 16 9 9 2
11 0 11 13 3 9 9 9 1 9 9 2
18 9 4 13 9 1 9 2 3 15 14 12 9 9 11 15 13 13 2
36 0 9 9 3 13 2 16 3 13 9 1 0 9 0 9 2 0 1 0 9 1 9 0 9 2 16 3 11 13 12 9 9 9 2 12 2
5 0 9 13 1 9
2 11 2
44 0 9 11 11 3 13 9 1 9 1 9 9 0 9 1 9 11 11 2 15 13 1 0 9 9 9 13 0 9 0 9 7 9 2 13 2 14 0 9 9 2 13 9 2
8 9 11 11 13 1 9 9 2
4 13 0 9 2
7 13 15 0 9 2 2 2
17 14 15 9 13 1 15 9 2 13 11 1 10 0 9 0 11 2
4 11 13 11 3
3 0 11 2
32 11 1 9 13 2 16 3 13 9 0 11 2 15 1 9 13 1 15 2 16 11 13 1 0 9 13 9 9 1 0 9 2
14 0 9 9 13 2 16 0 9 9 13 9 0 9 2
3 9 9 14
5 11 2 11 2 2
28 9 0 9 2 11 2 11 11 3 13 2 16 9 1 9 9 2 15 13 0 9 9 2 13 13 1 9 2
23 13 13 2 16 0 0 9 9 2 15 4 13 9 0 9 2 3 3 7 3 13 13 2
17 3 4 7 0 9 1 0 9 13 4 3 13 16 0 0 9 2
4 0 9 13 3
2 11 2
28 0 9 3 13 2 16 13 9 9 1 9 9 2 15 13 13 9 0 9 1 0 9 11 1 9 7 9 2
26 1 9 12 9 9 2 15 15 13 1 9 12 2 7 12 2 9 2 13 1 11 13 1 12 9 2
19 0 9 9 0 1 9 2 15 9 13 3 1 12 2 9 2 4 13 2
20 0 9 11 11 3 13 0 9 2 16 13 15 15 2 4 2 14 9 13 2
27 9 2 15 15 13 13 3 16 12 9 2 3 13 0 11 2 11 7 11 2 9 13 9 11 7 11 2
5 9 1 11 3 0
2 11 2
22 9 0 11 15 3 13 13 9 9 11 11 1 9 0 9 0 0 9 0 9 9 2
17 1 9 0 9 13 12 9 2 1 13 12 7 12 15 13 9 2
18 1 9 0 9 13 1 0 9 0 0 9 2 15 3 13 12 9 2
15 9 9 13 2 16 1 11 13 7 3 9 3 3 0 2
10 11 9 2 12 2 3 7 1 0 9
12 1 0 9 0 9 11 13 1 9 9 0 9
7 11 11 2 11 11 2 11
10 9 0 0 9 13 1 9 0 9 2
12 13 15 0 9 9 12 2 0 9 11 11 2
8 3 13 0 9 0 0 9 2
29 3 2 3 1 12 9 0 9 2 15 3 1 10 9 13 3 1 9 0 9 11 1 0 9 11 9 2 12 2
23 11 11 13 9 1 0 9 11 11 2 12 2 15 4 1 10 9 3 13 1 9 11 2
15 1 0 9 15 9 13 3 3 2 1 9 7 1 9 2
8 0 9 7 3 9 11 13 2
14 9 2 3 15 9 1 0 9 13 2 13 3 0 2
4 0 9 13 2
8 1 0 9 4 9 13 3 2
24 9 13 2 16 15 9 1 9 9 13 1 9 9 9 11 11 2 15 13 3 1 9 3 2
24 7 10 9 2 0 0 9 11 11 7 9 2 9 9 11 11 13 1 9 1 9 10 9 2
20 9 13 1 15 2 16 9 1 3 0 9 13 0 9 2 3 13 0 9 2
44 9 0 0 9 3 13 9 13 0 9 11 2 15 13 1 9 11 13 14 12 9 9 2 9 9 2 0 9 2 1 15 9 13 0 7 0 9 2 7 3 0 9 9 2
18 16 4 15 13 0 9 13 9 9 11 2 13 4 4 9 3 13 2
7 7 13 14 1 10 9 2
20 1 9 9 4 4 13 7 0 2 3 3 0 0 9 0 1 0 12 9 2
10 0 1 0 9 15 13 13 0 9 2
6 1 9 3 13 15 2
34 7 16 0 0 9 13 1 0 9 15 0 2 0 0 9 2 3 15 3 13 1 9 0 2 1 9 3 0 9 2 13 3 0 2
20 16 13 0 9 2 13 14 1 9 0 0 0 9 2 7 7 1 9 9 2
18 3 11 4 13 13 1 9 9 9 0 9 2 15 15 1 9 13 2
21 13 15 7 9 2 16 13 9 1 0 9 16 15 2 15 4 13 0 0 9 2
11 9 11 3 13 9 13 9 1 0 9 2
11 3 13 3 1 0 9 3 3 3 13 2
26 3 4 3 3 13 9 0 9 2 0 9 0 0 9 2 1 15 4 13 7 3 0 3 12 9 2
12 1 10 9 15 9 11 11 13 3 0 9 2
10 0 9 3 0 9 13 14 12 9 2
23 9 15 13 3 1 0 9 2 0 9 13 0 9 9 7 0 9 4 3 13 4 13 2
10 9 7 1 0 9 4 13 3 13 2
29 9 1 0 9 13 0 9 7 13 15 13 1 9 0 2 3 12 2 0 9 2 15 13 12 2 9 10 9 2
15 1 0 9 15 15 13 13 7 9 0 0 9 11 11 2
6 11 1 10 9 1 11
2 11 2
40 0 9 0 0 9 11 11 0 9 9 11 2 15 4 1 0 0 9 13 1 9 9 2 13 0 9 0 9 0 9 2 15 15 3 13 1 9 0 9 2
11 10 9 13 9 1 9 0 9 11 11 2
39 3 0 9 7 9 13 1 12 9 0 7 0 9 0 11 1 9 2 15 13 1 10 0 7 0 9 1 0 7 0 9 0 0 9 1 9 1 11 2
20 11 13 1 9 9 14 1 9 12 2 3 3 9 0 9 13 13 3 0 2
32 1 0 9 11 11 15 11 14 13 13 9 3 2 16 4 3 13 0 1 10 9 1 9 0 9 2 7 13 3 0 9 2
12 11 13 2 16 11 13 3 10 9 13 15 2
1 3
16 0 9 13 9 1 11 13 3 7 13 1 15 0 10 9 2
14 13 15 3 1 0 11 0 9 11 11 11 2 11 2
20 1 9 1 11 11 2 11 13 2 16 11 13 1 10 9 9 9 9 11 2
22 1 9 9 2 12 13 3 1 0 9 0 9 0 0 0 2 0 9 1 0 9 2
22 9 15 13 12 9 12 2 9 0 9 7 0 9 9 12 2 0 9 0 0 9 2
15 0 9 9 11 2 11 15 1 10 0 9 13 13 9 2
17 9 3 13 9 0 9 2 16 13 0 9 7 1 9 13 9 2
18 0 9 9 11 2 11 15 1 9 13 9 9 9 0 9 1 11 2
20 9 9 13 13 9 0 9 2 11 2 11 7 11 0 1 9 15 1 11 2
15 0 9 11 11 2 11 3 13 1 11 1 0 0 9 2
16 13 1 0 9 0 0 9 1 9 0 0 9 1 9 12 2
17 3 13 1 11 10 9 1 9 11 2 11 7 9 11 2 11 2
38 9 0 9 11 2 11 1 11 15 13 9 9 2 3 1 9 9 0 9 2 11 2 2 15 15 13 13 12 2 9 1 11 2 7 3 1 15 2
11 13 15 3 1 11 0 9 11 2 11 2
7 9 11 11 1 9 11 11
5 9 11 11 2 11
3 9 1 9
22 3 0 9 0 0 9 1 0 9 4 3 1 9 9 7 9 13 1 11 1 11 2
24 9 13 0 9 11 2 0 0 9 9 2 0 12 2 12 12 11 2 2 15 13 11 11 2
15 1 9 9 3 13 9 9 2 15 3 13 1 0 9 2
17 1 12 9 13 3 16 9 0 1 12 9 2 15 13 3 0 2
29 9 3 13 0 9 11 11 2 15 3 13 0 9 1 9 2 1 0 9 2 15 15 13 0 9 9 3 9 2
24 0 9 1 10 9 7 9 0 7 0 9 1 0 9 15 10 9 13 7 1 0 0 9 2
6 1 9 11 11 2 11
3 9 0 9
20 16 15 10 0 9 13 3 13 0 9 10 9 2 13 15 1 9 10 9 2
10 13 15 3 2 16 13 0 9 9 2
60 13 15 3 13 13 0 0 9 2 16 9 0 9 2 1 15 13 0 9 1 9 2 9 10 9 7 9 2 4 13 13 0 9 9 14 1 10 9 2 7 7 1 10 7 0 9 2 7 16 10 9 1 0 9 13 1 9 10 9 2
23 10 9 7 9 10 0 9 13 7 15 2 16 15 10 9 13 13 1 10 0 0 9 2
16 1 9 1 9 15 7 10 0 0 9 13 1 9 0 9 2
4 11 11 2 11
3 9 1 9
5 11 2 11 2 2
18 9 0 9 2 11 2 4 3 13 1 9 9 1 9 1 0 9 2
19 1 9 9 9 1 15 3 13 9 11 2 11 7 9 11 11 2 11 2
32 1 0 9 0 9 9 2 12 9 2 9 2 7 0 9 9 13 2 16 1 0 9 13 9 13 7 1 9 7 0 9 2
4 4 13 3 2
7 1 9 4 13 12 9 2
5 15 15 13 12 2
14 1 0 9 9 4 0 9 0 9 11 13 11 11 2
5 0 9 13 9 13
40 1 9 13 2 16 15 9 9 13 13 1 0 9 1 9 2 16 16 13 1 0 7 0 9 2 13 15 1 9 0 9 2 11 12 2 12 2 12 2 2
43 16 15 13 9 2 13 9 11 2 3 1 12 2 9 13 1 0 9 2 7 14 1 12 2 9 15 13 10 9 1 9 9 9 7 9 15 13 1 10 9 3 13 2
29 13 15 9 15 2 16 0 9 13 1 0 9 3 3 2 7 3 3 15 9 13 13 1 9 7 13 15 13 2
12 13 9 2 16 0 9 10 9 3 13 9 2
25 3 3 13 0 13 9 1 9 2 16 15 13 9 2 13 9 1 9 2 16 15 3 3 13 2
12 13 3 0 13 9 2 9 7 9 1 9 2
31 1 15 2 16 4 0 9 13 13 7 1 10 9 2 13 9 13 0 2 0 9 2 3 1 0 9 7 0 9 9 2
7 0 9 2 15 9 13 2
5 9 2 15 13 2
8 0 9 2 15 1 15 13 2
16 7 1 0 9 9 9 2 0 1 10 9 2 1 9 9 2
14 10 9 15 13 2 3 7 16 13 1 9 0 9 2
7 7 4 15 13 1 9 2
7 7 1 10 9 13 9 2
6 13 3 1 0 9 2
14 13 9 2 16 0 9 13 9 9 9 1 0 9 2
22 3 13 2 16 4 9 10 9 3 13 7 16 4 10 9 7 0 9 13 10 9 2
17 13 15 13 2 3 3 4 0 9 7 9 9 13 1 9 9 2
9 9 3 13 9 0 2 7 0 2
25 3 2 15 16 9 0 9 13 13 3 3 3 3 2 16 4 13 0 0 9 7 13 0 9 2
72 7 16 13 13 3 7 13 3 3 2 16 15 4 13 9 0 9 7 0 9 2 16 4 13 1 9 2 7 14 1 9 2 16 4 3 3 13 0 9 2 3 4 13 9 2 16 4 15 15 13 2 0 9 2 9 3 0 9 2 0 9 1 0 9 9 2 9 9 1 9 3 2
13 7 16 15 9 13 2 13 1 15 9 16 9 2
22 13 9 2 16 0 9 3 13 2 16 9 9 2 9 7 9 13 1 10 9 0 2
18 1 9 15 9 1 15 15 13 7 9 7 9 13 9 1 15 13 2
19 7 3 9 9 2 9 7 9 1 0 0 9 13 1 10 9 3 0 2
16 13 3 9 2 15 15 0 9 9 13 1 0 9 0 9 2
6 1 9 11 11 2 11
14 11 2 9 7 1 9 2 11 12 2 12 2 12 2
19 13 9 2 16 11 13 14 12 9 7 16 3 3 13 10 9 7 9 2
14 15 7 3 13 2 16 11 13 9 9 7 9 9 2
26 9 11 13 14 9 9 2 7 13 3 9 0 9 2 15 13 9 0 1 0 9 2 9 7 9 2
13 9 13 1 10 0 1 0 9 2 13 9 9 2
20 13 3 1 9 2 1 10 9 13 0 9 9 2 15 13 1 9 9 11 2
21 9 9 0 1 11 1 10 9 15 13 9 9 2 7 14 0 9 9 13 9 2
19 13 2 16 9 9 13 7 13 13 1 0 9 2 1 9 2 10 9 2
18 13 15 9 0 3 2 0 9 2 0 9 2 9 2 0 9 3 2
13 13 3 13 1 15 2 16 4 13 9 0 9 2
7 15 13 9 7 0 9 2
8 13 13 1 9 7 9 0 2
15 13 13 1 9 2 0 9 10 9 16 3 0 7 0 2
18 16 3 13 2 13 1 9 1 0 9 2 10 9 7 0 9 9 2
21 10 0 9 13 1 10 9 0 2 16 3 13 9 11 12 2 7 11 11 12 2
18 9 4 3 13 9 0 9 7 13 1 10 9 9 2 0 9 9 2
29 13 15 9 0 2 9 9 7 9 2 14 2 1 15 3 3 3 0 2 3 0 2 7 7 3 1 9 0 2
6 1 9 11 11 2 11
3 12 1 11
2 11 2
29 0 9 11 13 0 9 11 11 1 11 11 9 9 1 12 9 0 9 1 9 9 1 9 9 11 1 11 11 2
20 3 0 9 13 11 11 1 0 9 1 12 9 1 0 9 1 9 1 11 2
4 11 4 13 0
6 0 11 2 11 2 2
28 16 15 0 9 11 11 13 1 9 1 3 16 12 9 9 2 10 9 12 2 9 1 0 0 3 13 3 2
26 1 12 9 1 9 1 11 15 15 13 9 7 0 9 13 1 15 14 1 9 2 7 7 1 9 2
18 13 4 15 0 9 7 13 4 3 2 16 4 15 15 13 10 9 2
8 3 15 13 13 15 1 9 2
13 13 4 3 7 13 2 2 13 15 0 9 2 2
10 13 15 11 11 2 15 13 0 3 2
19 13 4 15 7 13 3 1 9 2 16 4 15 13 2 13 0 9 11 2
16 16 15 14 3 1 0 9 13 16 9 2 9 1 9 13 2
2 0 9
4 9 1 9 2
2 11 2
41 1 9 12 2 0 9 1 11 13 9 0 0 9 2 11 2 7 9 0 0 9 11 11 2 16 4 9 9 1 9 12 1 0 11 13 13 12 9 1 9 2
8 1 15 13 7 0 9 9 2
3 9 1 9
2 11 2
19 9 0 9 11 2 11 7 11 15 1 9 13 1 11 9 9 9 9 2
32 1 9 12 9 13 10 9 1 12 0 9 2 15 13 9 1 9 10 9 2 15 15 13 12 2 9 1 11 1 11 2 2
3 1 0 9
13 11 11 7 11 13 0 9 1 0 9 11 11 2
7 12 13 1 0 11 11 2
12 11 11 3 13 9 1 12 0 9 0 11 2
14 1 9 1 0 9 11 1 11 11 11 2 3 2 2
5 9 11 11 2 11
8 14 1 9 2 7 7 1 9
11 11 1 9 1 0 9 9 1 11 13 11
9 11 2 11 2 11 2 11 2 2
38 0 9 15 1 9 13 7 0 10 9 3 4 13 1 11 2 3 1 9 13 0 0 9 9 11 11 1 0 9 1 9 1 9 11 1 9 12 2
9 12 9 13 1 11 1 0 9 2
13 10 9 15 3 13 13 3 3 2 11 13 3 2
22 0 15 3 3 13 1 9 11 1 11 1 11 2 9 13 0 9 11 1 9 11 2
25 9 1 11 15 3 13 1 11 1 11 2 3 15 13 1 11 2 3 15 1 15 13 0 9 2
10 9 13 3 1 9 0 9 1 11 2
19 13 7 1 15 0 9 11 2 15 1 0 9 1 11 1 11 3 13 2
19 10 9 13 11 1 11 2 15 1 9 11 1 12 9 13 11 1 11 2
36 3 15 1 12 9 13 1 11 0 9 9 11 1 0 11 1 12 5 12 9 2 1 9 4 0 9 13 1 9 9 11 11 11 1 11 2
20 9 1 9 15 12 9 13 9 1 11 2 9 11 1 12 7 15 1 12 2
32 0 9 13 1 9 1 12 7 13 9 13 13 14 0 9 9 11 2 0 9 13 3 12 10 9 2 2 7 3 0 9 2
40 1 0 9 15 13 9 1 12 9 2 1 0 9 1 9 1 12 9 7 0 1 9 2 9 7 9 1 12 9 2 9 1 12 9 7 9 13 9 3 2
15 9 9 11 11 13 9 12 9 2 1 15 13 1 9 2
20 1 9 2 15 1 12 9 13 1 11 0 9 1 11 2 13 14 9 11 2
22 15 9 13 1 0 9 2 0 9 11 11 15 3 1 0 11 13 3 1 0 11 2
5 0 9 1 11 2
5 11 2 11 2 2
16 0 0 9 2 0 3 0 9 2 13 1 0 9 10 9 2
24 0 9 7 13 13 3 7 1 9 2 3 13 10 9 0 0 1 0 0 9 1 12 9 2
19 0 9 13 12 9 2 15 13 9 9 9 0 9 11 11 7 11 11 2
21 3 0 9 1 11 15 13 3 9 1 11 7 3 1 9 1 9 13 0 9 2
9 12 9 13 1 11 1 12 9 2
6 0 9 1 11 2 11
2 11 2
18 9 1 11 13 3 9 9 0 9 11 11 1 9 9 10 0 9 2
16 0 9 1 9 0 9 1 9 9 0 9 13 12 2 9 2
41 0 0 9 11 13 1 9 1 9 1 0 9 1 9 2 16 10 9 11 2 11 13 2 16 13 3 9 2 16 4 3 13 15 9 1 0 9 1 0 9 2
8 11 13 13 1 9 12 9 2
23 1 9 13 13 12 9 10 9 1 11 1 9 1 11 2 11 7 11 7 9 1 11 2
13 0 9 4 1 9 10 9 3 13 1 10 9 2
38 1 0 9 13 11 13 9 1 9 12 0 9 2 12 9 2 1 9 11 11 1 9 1 9 7 9 0 9 7 13 15 13 9 1 0 9 11 2
18 3 1 9 3 13 11 11 13 11 0 12 0 9 2 12 9 2 2
26 11 4 3 3 13 7 13 1 9 14 1 9 9 12 0 9 2 12 9 2 7 0 9 10 9 2
4 0 9 13 11
2 11 2
24 0 0 9 13 9 1 9 0 0 9 1 9 0 0 9 2 0 1 0 9 11 11 11 2
14 0 9 1 10 9 13 0 0 9 9 2 11 11 2
11 9 1 12 0 9 3 13 1 0 9 2
27 9 11 11 11 15 3 1 9 11 0 0 13 3 3 1 0 9 7 13 9 1 3 0 1 0 9 2
24 11 15 13 10 9 13 7 10 9 13 2 16 13 11 13 1 9 9 1 9 12 9 9 2
3 9 7 9
2 11 2
18 11 7 11 13 1 0 9 1 0 9 0 9 1 0 9 1 11 2
31 0 9 0 9 3 0 9 13 1 0 9 11 2 11 12 2 12 2 7 1 0 9 13 11 11 7 11 12 2 12 2
3 0 9 11
4 11 1 11 2
15 9 0 0 9 11 11 11 13 1 9 10 9 12 9 2
19 9 13 10 9 9 0 9 1 9 9 11 2 11 2 12 2 12 2 2
25 11 2 15 13 1 9 11 1 9 12 2 13 11 11 1 9 7 10 9 13 0 9 9 11 2
10 1 0 9 13 11 9 3 16 9 2
24 1 9 12 15 3 13 1 9 1 9 11 7 0 11 2 1 15 15 13 9 1 12 9 2
7 9 12 2 9 12 2 9
4 9 2 12 2
19 11 2 11 2 7 11 13 2 11 2 11 2 7 11 2 11 2 13 2
3 2 11 2
4 1 11 13 11
7 12 9 13 1 10 0 9
5 11 2 11 2 2
24 0 9 15 0 9 1 11 13 1 9 0 9 2 7 1 9 10 9 13 0 12 9 9 2
28 1 0 9 12 2 9 15 3 13 7 9 2 16 9 13 1 0 0 9 3 0 9 11 2 11 2 2 2
15 11 13 1 9 1 0 9 1 11 1 12 9 1 9 2
16 1 9 13 11 7 3 9 9 13 3 3 7 1 9 11 2
10 1 9 1 15 13 11 11 7 11 2
26 3 1 9 1 11 4 13 2 16 9 2 15 13 2 13 9 2 13 0 9 11 3 1 9 11 2
20 11 13 3 1 0 9 11 1 11 2 15 15 13 1 9 3 7 3 13 2
13 9 11 2 1 11 1 9 13 2 7 3 13 2
19 1 11 15 7 13 3 9 1 9 7 13 4 0 2 16 4 3 13 2
14 13 4 15 13 1 9 2 7 10 9 15 15 13 2
40 1 0 0 9 13 3 12 9 1 10 0 9 2 0 11 1 11 2 11 1 11 1 11 2 0 11 1 11 7 3 11 13 3 10 9 1 11 1 11 2
9 9 1 0 9 9 11 13 9 2
27 1 9 1 9 3 13 1 0 9 7 7 1 11 13 2 16 13 0 9 2 13 11 1 10 0 9 2
7 0 9 0 11 13 1 9
7 11 2 11 2 11 2 2
18 0 9 11 11 7 10 9 11 11 13 1 9 11 1 9 9 11 2
26 0 9 1 10 9 13 0 9 0 9 11 11 2 1 0 9 15 13 9 12 3 0 9 0 11 2
18 13 1 15 0 9 2 15 13 0 9 0 9 1 9 1 11 11 2
26 9 11 7 9 11 3 15 13 1 9 1 0 9 3 2 3 15 10 9 13 0 0 9 1 9 2
13 1 0 9 9 13 15 1 0 9 9 1 11 2
14 9 13 1 9 0 9 0 9 0 9 11 2 11 2
15 9 13 3 12 9 2 1 15 12 13 0 2 0 9 2
21 1 11 2 11 4 9 13 1 10 9 2 16 15 1 12 9 0 11 13 12 2
22 11 2 11 13 2 16 15 3 13 13 0 12 9 2 12 1 9 7 0 1 9 2
25 1 9 11 2 3 4 13 9 2 16 4 13 9 2 11 2 11 13 2 16 1 15 4 13 2
16 9 9 1 9 11 2 11 2 1 9 9 11 2 11 7 11
5 9 11 11 2 11
4 13 7 0 9
9 16 4 11 13 9 2 13 4 9
5 11 2 11 2 2
39 1 9 0 9 13 1 11 12 9 2 7 2 9 13 9 1 11 2 11 13 1 9 1 11 7 1 9 7 11 1 9 1 9 1 9 1 9 11 2
22 11 10 9 2 3 1 0 9 2 13 1 12 0 9 7 3 1 9 1 0 9 2
26 13 4 9 13 1 0 9 2 7 3 4 15 13 1 0 9 2 13 10 9 12 0 11 11 2 2
14 13 10 9 2 16 15 1 11 13 1 9 1 11 2
3 3 14 2
17 1 11 4 13 12 9 1 9 2 7 15 1 9 10 9 13 2
15 9 13 2 16 4 13 9 2 16 0 9 13 0 9 2
7 13 4 13 3 14 3 2
10 1 11 15 3 16 3 13 0 9 2
2 3 2
11 13 15 13 13 9 2 3 12 1 15 2
12 3 15 13 3 1 12 9 2 15 13 0 2
21 14 15 15 13 0 9 2 3 15 1 9 13 12 9 2 7 1 9 14 12 2
5 13 15 11 9 2
7 3 4 1 15 13 3 2
21 1 15 13 15 1 10 9 14 3 2 3 7 3 13 9 9 2 9 2 9 2
14 3 15 13 13 9 0 9 11 7 9 9 1 11 2
13 3 3 2 13 15 1 9 7 9 13 10 9 2
13 3 15 14 13 7 13 2 16 13 15 1 9 2
5 3 13 9 9 2
11 9 11 11 2 3 4 9 13 0 9 2
5 11 2 11 2 2
7 13 4 12 1 0 9 2
40 1 9 4 15 13 2 16 4 13 3 2 7 3 4 9 13 0 9 2 13 15 1 9 12 2 9 0 9 11 2 11 2 12 2 12 2 9 9 11 2
19 0 9 13 1 9 0 9 2 15 13 9 0 9 1 9 1 0 9 2
18 9 1 9 0 0 9 7 0 9 0 11 13 1 0 9 0 9 2
25 11 15 13 9 2 16 0 9 9 13 13 3 7 3 7 1 9 0 9 13 9 1 0 9 2
6 10 0 9 9 13 2
25 16 11 13 1 9 9 7 3 13 3 13 1 10 9 2 7 1 9 15 3 13 16 10 9 2
29 1 0 9 13 3 3 3 1 9 2 12 15 9 1 9 13 2 2 7 1 12 9 14 3 13 3 1 9 2
6 15 13 9 0 9 2
13 0 9 9 13 0 9 1 0 9 1 11 11 2
29 16 9 3 13 1 9 2 13 9 1 0 9 2 13 15 15 2 16 4 15 1 9 13 9 7 9 1 9 2
9 0 7 13 2 3 0 13 9 2
23 9 2 15 13 1 9 2 11 2 11 2 13 2 7 7 0 16 4 13 9 7 9 2
26 3 3 15 1 9 13 2 16 3 0 9 11 11 13 1 0 9 3 3 1 0 9 16 1 9 2
16 13 3 9 2 16 10 9 15 13 9 1 0 9 0 9 2
9 9 1 0 9 15 9 13 3 2
25 3 3 1 9 13 9 9 1 0 9 1 11 2 15 13 1 10 9 2 7 9 15 3 13 2
6 11 4 13 1 15 13
19 9 10 9 3 13 9 14 16 0 9 2 13 9 0 9 11 11 2 11
18 1 9 9 1 11 1 15 13 10 9 7 13 15 16 0 9 9 2
21 13 15 2 16 13 15 1 15 2 16 4 4 13 1 9 1 9 9 0 9 2
11 13 15 2 16 15 13 11 2 7 11 2
7 13 2 9 15 3 13 2
50 3 13 11 11 2 3 1 11 7 11 2 9 0 0 9 0 11 7 1 9 12 9 11 2 1 15 3 1 11 13 9 9 9 2 3 3 1 9 1 9 1 11 13 9 1 9 0 9 2 2
5 15 13 10 9 2
7 13 15 0 7 0 9 2
24 3 4 1 15 15 13 2 7 13 4 2 16 13 1 0 0 9 0 9 14 1 9 12 2
22 9 1 0 9 7 11 13 13 3 0 9 2 3 13 0 9 0 11 1 0 11 2
6 13 4 15 10 9 2
4 9 13 9 2
15 13 2 16 15 4 0 2 15 13 0 2 7 14 0 2
14 13 13 1 9 0 9 7 13 9 2 15 15 13 2
14 3 1 9 15 3 13 15 15 13 1 9 0 9 2
10 9 13 3 0 7 15 15 13 13 2
11 9 10 7 15 0 9 13 1 10 9 2
9 3 4 15 13 13 1 0 9 2
6 3 2 3 14 2 2
16 1 9 9 1 11 4 13 1 9 0 9 1 9 0 9 2
6 15 13 9 1 11 2
8 1 9 4 15 0 9 13 2
20 1 9 1 0 9 4 15 7 14 13 10 0 0 9 2 15 13 0 9 2
18 15 2 1 15 2 13 1 9 0 2 7 10 9 15 1 15 13 2
16 7 1 9 4 1 9 9 0 0 9 13 10 9 11 11 2
11 13 15 11 11 2 9 10 9 11 11 2
6 13 4 15 1 9 2
4 13 0 9 2
15 13 15 14 1 10 9 2 1 10 13 9 1 9 12 2
5 0 9 15 13 2
17 13 14 15 2 16 3 13 9 11 7 11 13 0 9 1 9 2
15 16 4 7 0 9 13 1 9 0 9 2 15 4 13 2
11 1 9 13 7 10 0 9 1 0 11 2
18 3 4 1 9 1 0 0 9 13 9 13 13 1 12 0 0 9 2
20 3 4 1 9 13 7 11 2 1 15 13 3 9 2 15 13 9 0 9 2
11 13 15 1 10 9 13 2 7 3 13 2
10 1 10 9 3 13 1 15 3 13 2
18 13 0 2 16 15 13 3 13 2 9 11 2 3 4 13 9 2 2
7 13 15 7 13 16 9 2
12 3 3 15 13 9 0 9 0 9 1 9 2
7 1 15 15 3 13 13 2
21 10 9 13 13 9 1 0 9 1 9 1 15 2 1 10 9 7 3 3 13 2
13 13 3 15 2 15 13 13 9 1 9 3 0 2
12 13 0 9 7 13 15 2 15 13 3 0 2
10 3 7 3 13 9 9 1 0 11 2
26 7 1 9 4 15 13 13 2 16 4 0 7 0 9 13 2 16 4 9 13 1 9 1 0 9 2
20 11 13 0 0 9 2 1 15 13 1 15 2 7 7 1 15 3 3 3 2
19 16 0 9 4 1 9 11 7 11 13 0 0 9 2 15 15 9 13 2
5 15 13 10 9 2
7 3 13 9 13 0 9 2
13 11 7 11 13 0 9 7 13 9 1 0 9 2
13 7 16 4 13 0 9 2 0 9 4 3 13 2
19 16 4 15 1 15 13 2 13 15 3 0 9 2 15 15 13 1 9 2
11 9 13 15 13 2 15 15 13 13 9 2
7 1 15 13 15 3 9 2
11 10 9 7 3 13 9 3 16 0 9 2
7 3 15 15 13 9 11 2
7 1 10 9 10 9 13 2
15 13 15 0 9 13 2 10 0 9 15 1 9 13 3 2
30 13 7 0 2 16 15 3 15 4 13 9 9 9 2 13 1 15 2 7 3 7 1 0 9 9 1 0 9 13 2
3 13 15 2
12 9 11 13 13 9 9 1 0 9 2 2 2
3 0 9 2
8 9 13 2 10 15 13 9 2
19 13 4 3 9 0 9 7 9 9 2 3 3 9 13 7 9 1 9 2
6 9 1 9 13 0 2
7 1 9 13 13 9 11 2
21 1 11 13 0 7 1 9 9 1 11 3 1 10 9 13 0 9 2 11 11 2
5 15 13 1 15 2
9 13 13 9 0 1 9 13 3 9
7 11 2 11 2 11 2 2
21 9 0 9 2 1 15 15 1 0 9 13 0 9 9 11 2 13 3 3 9 2
10 13 15 9 9 11 1 0 9 9 2
16 1 11 15 3 13 3 14 3 2 7 15 3 1 9 12 2
6 3 13 1 0 9 2
17 1 9 9 0 9 9 11 15 7 7 3 13 1 9 3 3 2
8 1 9 9 4 13 0 9 2
7 3 4 7 9 13 9 2
9 1 11 13 3 14 10 0 9 2
16 1 0 9 15 7 4 3 13 0 9 2 15 13 0 9 2
7 1 0 11 15 3 13 2
17 0 9 0 9 15 7 13 1 9 13 0 9 9 1 0 9 2
19 1 0 9 1 11 13 9 1 0 0 9 2 10 9 3 13 9 9 2
10 16 7 13 9 2 13 12 9 9 2
14 3 13 9 1 9 0 2 1 9 15 7 3 13 2
16 3 0 9 2 15 13 1 0 9 1 11 2 13 12 9 2
20 0 9 13 0 0 9 1 9 2 3 15 9 13 1 0 9 1 9 9 2
22 16 7 13 1 9 0 9 2 15 4 13 9 0 9 2 4 9 13 14 0 9 2
4 9 9 1 9
7 11 2 9 11 11 2 2
39 0 9 2 15 3 9 13 0 0 9 0 9 7 10 0 9 2 13 9 9 2 1 15 4 1 11 13 16 9 3 0 9 9 2 11 1 0 9 2
10 9 13 0 7 3 4 13 0 9 2
11 9 1 9 4 13 14 1 9 1 9 2
25 9 13 2 16 10 9 15 13 9 7 9 9 2 15 15 1 9 9 13 3 3 13 0 9 2
10 1 10 9 13 13 1 9 7 9 2
8 9 9 1 0 9 13 14 3
7 11 2 11 2 11 2 2
26 0 9 0 9 1 11 11 11 13 13 13 1 9 0 0 9 2 11 2 11 11 1 9 0 9 2
48 9 11 11 7 11 11 3 1 10 0 9 1 11 13 1 0 9 9 9 1 12 0 9 1 9 11 2 7 0 9 1 0 9 9 1 0 9 12 9 13 1 0 9 1 9 10 9 2
14 13 0 2 16 9 13 9 1 0 2 9 0 9 2
13 10 9 13 1 15 0 2 13 11 3 1 11 2
13 11 11 13 3 3 1 9 9 1 10 9 0 2
40 13 3 0 9 2 7 1 10 9 13 3 13 1 15 2 16 4 9 0 9 13 13 9 2 0 9 10 0 9 2 3 1 0 9 2 13 15 1 9 2
19 9 0 9 11 11 2 15 13 0 9 9 2 13 1 10 9 1 9 2
7 9 1 9 13 13 9 11
13 0 9 4 1 9 13 7 11 15 13 1 10 9
5 11 2 11 2 2
43 9 1 9 7 9 9 11 2 11 2 15 13 13 2 1 10 9 11 13 7 13 0 9 1 11 2 10 12 9 13 1 9 12 1 9 11 12 9 0 9 7 11 2
13 0 9 13 10 9 16 9 0 9 0 0 9 2
13 9 15 13 9 1 9 1 0 9 7 0 9 2
21 9 11 3 0 9 1 9 13 2 10 9 9 13 9 13 7 13 1 0 9 2
17 3 4 1 9 1 9 13 12 9 2 1 15 12 1 9 9 2
25 9 2 16 15 9 9 11 11 2 0 0 9 1 9 2 4 13 11 2 15 3 13 13 9 2
35 11 15 13 13 9 1 9 1 0 9 9 2 9 11 0 9 2 15 1 15 13 0 0 9 7 1 15 13 9 2 16 13 1 11 2
9 13 0 2 16 10 9 3 13 2
23 1 11 11 1 11 15 13 13 9 2 15 13 2 16 11 1 9 0 9 13 7 13 2
21 13 3 2 1 10 9 15 11 13 2 13 2 7 3 13 7 13 15 15 13 2
31 1 10 9 15 13 2 16 9 13 0 9 7 9 1 9 11 7 9 2 7 9 11 13 2 16 4 0 9 4 13 2
24 3 15 7 3 1 10 9 9 13 11 1 9 7 12 3 15 0 9 13 9 1 0 9 2
11 11 2 11 7 13 10 9 1 3 0 2
16 15 11 2 15 9 13 2 16 13 0 9 2 15 13 3 2
19 0 9 3 13 2 16 15 13 7 16 15 13 2 14 16 15 13 9 2
10 3 0 13 1 11 3 9 0 9 2
14 0 9 1 12 0 9 13 3 0 9 1 10 9 2
17 7 15 13 13 2 16 0 9 13 13 0 7 0 9 1 9 2
4 9 1 9 13
10 9 9 3 7 3 7 0 9 3 13
9 11 2 11 2 11 2 11 2 2
30 0 9 9 1 9 11 2 11 0 3 7 3 0 9 12 0 0 9 9 13 7 0 9 0 9 9 11 1 11 2
18 9 11 11 2 11 2 15 13 2 16 0 9 4 13 1 0 9 2
17 9 4 3 13 15 9 9 7 0 9 4 15 7 13 10 9 2
14 13 15 9 13 9 1 9 2 15 13 2 13 9 2
31 11 11 2 9 0 2 15 13 0 2 16 13 9 3 7 3 0 2 7 1 3 0 13 9 9 16 9 2 7 9 2
12 1 9 4 13 9 7 11 11 2 11 2 2
21 13 15 0 9 2 13 2 7 13 4 13 2 15 15 13 1 9 9 1 9 2
28 11 11 2 11 2 13 2 16 3 0 9 4 13 1 9 3 3 2 16 1 15 9 4 3 13 10 9 2
24 9 11 13 11 11 11 2 9 11 2 11 13 1 9 7 15 11 13 1 3 0 7 0 2
9 15 13 9 1 9 7 0 9 2
7 7 9 9 3 13 4 2
21 11 11 2 11 2 15 13 0 2 16 13 3 0 9 2 16 3 13 9 0 2
19 16 7 3 13 0 9 2 13 11 1 0 2 16 4 4 13 3 3 2
21 9 4 13 13 9 15 13 1 9 1 9 10 12 9 2 16 13 13 0 9 2
12 1 0 9 15 15 13 10 9 2 13 11 2
28 0 0 9 11 11 2 11 2 11 2 13 13 2 16 9 13 0 9 2 1 15 15 9 13 2 16 13 2
13 3 15 10 9 13 1 15 3 2 16 13 9 2
14 13 7 2 16 9 9 9 13 0 16 9 9 9 2
29 9 9 1 0 9 13 3 1 11 1 11 10 9 1 9 11 11 2 12 2 9 9 1 9 0 9 1 9 2
13 1 0 9 13 1 11 13 1 12 3 0 9 2
5 9 11 11 2 11
8 0 9 4 13 1 11 0 9
5 11 2 11 2 2
29 0 12 9 0 9 15 13 1 0 9 9 2 3 13 10 9 2 13 3 9 9 9 7 9 9 9 11 11 2
29 0 9 13 1 15 10 0 9 2 9 13 9 1 0 9 9 2 13 0 9 0 9 7 13 9 9 0 9 2
19 9 2 10 9 3 11 13 2 4 13 1 9 13 0 9 16 0 9 2
18 9 0 9 1 0 9 4 7 13 0 9 2 3 1 0 9 2 2
19 1 9 9 13 9 11 13 9 9 2 10 9 7 9 13 9 9 9 2
21 1 0 9 13 12 9 9 2 0 12 9 13 13 1 0 9 0 7 0 9 2
20 13 1 15 12 9 9 2 15 13 3 1 0 0 9 2 13 11 2 11 2
13 3 3 1 10 9 13 9 0 9 1 9 11 2
10 9 11 4 13 9 9 1 9 9 2
15 1 9 9 13 9 0 1 9 0 9 7 1 9 9 2
8 9 0 9 4 13 9 9 2
4 9 3 0 9
6 9 13 15 0 16 15
2 11 11
9 15 13 3 13 2 1 9 13 2
10 13 7 3 9 2 3 15 9 13 2
23 1 12 1 0 9 0 0 9 3 3 13 2 16 12 9 4 13 1 9 1 3 0 2
5 7 13 0 9 2
9 9 13 1 11 1 9 9 12 2
10 3 15 13 1 0 9 9 9 12 2
24 2 2 2 9 13 9 3 16 9 13 15 9 2 13 15 7 13 3 0 9 1 0 9 2
11 9 13 13 1 9 9 2 3 7 9 2
20 13 15 1 10 9 2 16 13 9 2 0 9 2 3 0 9 2 0 9 2
24 9 9 13 1 9 13 1 0 9 2 16 3 12 9 15 9 13 1 9 9 12 2 12 2
14 9 0 9 2 7 15 16 0 9 2 13 9 12 2
23 9 9 1 0 2 9 12 2 13 3 0 9 2 15 13 3 0 2 3 7 0 9 2
10 9 12 13 3 0 9 0 1 9 2
39 9 1 9 1 11 2 0 9 0 9 1 0 9 2 2 9 12 2 13 3 0 9 2 3 3 9 12 13 0 9 16 9 12 2 7 1 0 9 2
41 9 1 9 1 12 15 13 1 12 9 2 15 1 9 12 13 1 15 3 2 13 3 7 15 2 15 10 9 13 0 2 7 13 15 3 9 9 7 9 2 2
16 9 1 9 1 12 2 7 1 12 2 13 3 14 12 9 2
4 1 0 0 9
27 9 2 15 13 0 9 3 0 9 2 13 3 0 1 9 2 1 15 4 0 2 0 9 13 9 0 2
7 3 4 15 1 15 13 2
10 3 2 16 4 15 13 10 0 9 2
30 15 4 15 13 1 0 9 2 9 4 13 3 3 2 7 10 0 9 9 4 15 1 9 3 13 1 9 9 0 2
5 0 1 0 9 2
21 1 10 9 10 0 9 4 10 9 13 9 2 16 4 7 15 15 13 3 13 2
14 3 1 0 9 13 3 0 9 16 0 7 0 9 2
20 16 10 9 3 3 13 7 0 9 2 9 1 15 3 13 0 9 10 9 2
14 1 15 15 13 2 16 1 0 9 13 3 10 9 2
17 1 9 15 13 2 13 2 1 9 15 1 10 9 13 0 9 2
14 3 1 0 2 0 9 9 1 15 3 13 9 9 2
5 13 0 7 0 2
10 9 1 15 13 0 9 1 0 9 2
5 0 9 13 1 9
34 3 13 3 3 9 0 7 0 2 15 3 2 1 10 0 9 2 13 1 9 7 9 3 2 16 15 3 13 3 13 7 3 13 2
29 10 9 15 1 9 15 13 2 13 0 9 1 0 9 7 9 1 9 7 3 3 1 0 9 13 1 15 0 2
15 3 1 15 13 0 9 1 3 0 9 1 9 0 9 2
14 13 0 13 2 16 7 1 9 13 9 2 15 13 2
10 16 13 15 3 0 2 3 15 13 2
7 3 7 3 13 0 9 2
16 1 12 15 13 7 12 0 2 15 0 0 9 13 1 9 2
3 0 0 9
8 0 9 3 13 3 0 9 2
15 13 1 15 0 2 3 0 9 13 0 14 1 0 9 2
18 15 1 15 3 13 9 0 1 0 9 2 16 13 3 3 0 9 2
11 3 13 0 9 2 7 3 13 1 9 2
3 7 3 2
8 9 1 15 13 9 0 9 2
30 0 13 9 2 3 13 1 0 9 3 13 1 9 1 9 2 7 16 1 9 1 9 2 9 7 9 1 0 9 2
25 13 9 2 15 15 10 0 9 13 0 13 2 3 16 10 0 9 13 0 3 13 9 3 0 2
5 11 15 0 9 13
19 16 9 1 0 9 13 0 2 0 9 1 15 3 0 1 15 3 13 2
9 1 11 15 3 13 1 9 11 2
6 13 15 9 0 9 2
7 9 13 15 0 16 15 2
39 11 0 9 15 3 13 13 1 15 0 0 9 1 3 0 9 2 7 16 1 15 13 0 9 2 13 1 9 9 12 3 0 9 11 1 0 12 9 2
15 3 9 1 11 4 13 15 0 2 1 0 9 7 13 2
14 3 13 13 9 7 10 9 2 1 9 13 3 13 2
16 13 1 0 9 9 1 9 1 11 13 1 0 9 3 0 2
24 9 0 9 11 2 15 10 0 9 13 2 3 11 1 0 9 2 0 9 1 0 9 13 2
10 3 4 13 13 7 0 7 0 9 2
13 1 0 9 13 9 9 13 9 2 9 7 9 2
16 3 10 0 9 15 13 1 9 9 3 9 10 9 16 9 2
6 11 15 0 9 13 2
20 10 9 1 15 3 13 2 7 7 10 0 9 13 1 0 9 7 0 9 2
2 3 13
33 16 4 0 1 9 2 15 15 3 3 13 1 9 0 9 2 10 0 9 1 12 9 13 2 13 4 9 1 9 1 0 9 2
8 13 0 3 13 13 0 9 2
35 7 10 9 1 0 9 13 1 15 2 1 10 9 13 0 13 2 13 2 14 15 3 1 9 3 16 1 0 9 2 16 1 0 9 2
22 10 0 9 13 3 0 9 1 9 9 9 2 0 7 0 9 7 0 9 1 9 2
9 1 9 9 0 9 13 7 9 2
3 11 1 11
17 9 11 11 13 1 9 1 11 0 0 9 7 0 0 11 1 11
2 11 11
4 0 0 9 2
19 1 12 0 9 9 2 15 13 13 9 0 9 0 9 1 9 0 9 2
14 1 9 10 9 3 2 7 3 1 0 9 2 13 2
16 13 15 3 2 12 9 1 0 9 2 0 9 0 0 9 2
9 1 9 9 2 9 7 9 3 2
21 12 1 9 2 3 0 9 13 9 0 9 2 13 13 9 0 1 10 0 9 2
6 15 15 3 13 3 2
11 7 1 9 9 13 13 0 9 9 9 2
9 10 9 1 12 9 15 13 13 2
54 13 13 10 0 9 9 1 0 2 0 0 9 12 7 9 9 9 3 2 15 13 12 12 12 9 12 9 3 2 13 11 11 2 9 0 0 11 1 11 2 0 0 0 9 2 15 3 13 10 0 0 0 9 2
5 1 0 9 3 9
12 9 3 12 12 3 15 13 0 9 0 9 2
13 10 9 15 13 13 13 10 9 1 9 0 9 2
12 13 15 1 0 9 3 9 2 13 9 11 2
16 7 1 9 10 0 9 15 15 13 14 12 2 15 15 13 2
4 15 15 0 2
12 1 0 12 4 13 9 0 9 2 13 11 2
6 1 10 0 0 9 2
35 15 4 13 9 12 12 3 2 15 14 12 7 15 2 15 7 13 0 9 1 0 9 1 0 9 2 3 14 9 12 9 12 9 3 2
22 1 9 0 11 2 0 1 11 7 0 0 7 0 9 7 9 2 13 0 9 13 2
14 3 15 13 9 2 10 9 15 7 0 9 13 13 2
17 3 1 15 13 0 9 2 1 9 0 1 0 2 16 10 9 2
12 0 13 13 15 2 10 9 15 0 9 13 2
15 0 9 1 9 12 9 0 11 13 14 12 9 9 3 2
23 3 13 0 13 2 13 2 14 9 9 13 1 9 2 1 15 4 9 0 9 13 9 2
16 7 7 4 13 9 3 9 0 1 0 9 2 10 0 9 2
19 13 15 2 16 9 2 16 13 3 1 9 0 0 9 2 13 0 9 2
19 1 0 9 15 1 11 13 14 9 0 9 2 7 1 15 0 9 9 2
4 13 0 9 2
13 4 13 9 3 1 3 0 9 2 13 9 11 2
16 1 11 13 9 1 9 3 12 9 12 9 2 13 11 11 2
28 1 15 15 13 1 0 0 9 1 11 0 1 9 2 15 1 10 9 13 9 1 10 9 2 16 4 13 2
3 9 3 0
13 3 15 1 11 13 9 1 9 0 9 1 11 2
21 1 11 13 15 0 9 9 2 15 13 9 13 15 0 2 16 13 0 0 9 2
27 9 9 13 0 0 9 2 9 7 9 9 11 1 11 2 13 3 16 0 9 0 9 1 9 12 2 2
19 16 0 9 13 1 9 1 9 0 9 2 15 0 0 9 13 3 0 2
19 9 7 9 2 15 4 13 1 9 2 13 1 0 0 9 7 0 9 2
21 1 10 9 12 9 1 9 9 13 1 0 9 2 3 0 11 13 2 3 9 2
50 3 3 7 9 0 9 13 15 16 3 1 9 2 3 15 9 11 1 10 9 11 7 9 11 11 13 1 0 9 1 0 0 9 7 13 9 1 9 7 10 9 2 16 1 0 9 15 13 0 2
9 10 9 4 1 0 11 3 13 2
27 1 0 0 9 13 12 12 0 2 1 12 9 2 2 12 12 0 2 1 12 9 2 7 12 0 9 2
4 3 10 9 2
22 0 4 13 9 12 9 1 9 13 1 3 0 9 11 2 11 11 1 0 11 2 2
28 1 0 12 9 4 13 13 9 2 11 11 2 2 0 9 2 3 1 0 9 7 0 3 1 15 9 9 2
18 12 9 15 13 1 9 2 15 13 1 15 9 1 0 11 0 9 2
24 0 15 1 12 9 13 1 0 9 0 3 1 11 2 15 13 2 16 15 15 4 13 13 2
11 0 15 4 13 1 0 9 0 1 11 2
5 15 15 4 13 2
19 1 9 9 0 9 15 13 2 16 10 9 11 11 3 9 1 9 13 2
21 3 1 9 13 12 9 2 15 1 9 13 13 1 0 9 2 7 12 0 9 2
5 13 0 2 9 2
13 15 0 9 2 15 15 4 13 3 2 4 13 2
12 10 9 4 13 3 0 9 2 13 11 11 2
15 3 9 0 9 13 1 0 11 2 3 13 1 0 9 2
11 9 4 13 10 0 9 1 11 1 11 2
23 9 7 9 4 13 1 9 9 1 11 2 15 13 9 1 9 1 11 7 13 3 3 2
8 13 1 11 1 10 0 9 2
14 9 13 15 9 1 10 9 7 15 13 3 3 3 2
24 15 15 13 7 0 9 2 15 13 1 15 2 15 4 13 1 0 9 7 3 13 0 9 2
6 9 2 0 2 7 0
12 0 9 1 0 0 9 4 13 14 0 0 2
25 7 15 9 11 13 2 15 15 13 13 1 9 2 16 15 13 12 9 1 0 0 11 1 11 2
10 13 15 15 2 15 15 13 1 11 2
4 9 13 0 2
31 16 4 13 2 16 13 1 9 2 13 15 1 15 9 0 11 1 15 2 16 13 15 0 2 15 4 13 9 1 11 2
4 3 13 3 2
19 1 10 9 1 9 11 11 13 0 9 2 1 15 4 9 10 9 13 2
7 13 0 2 7 3 0 2
18 11 11 13 2 16 15 15 13 2 2 13 0 9 1 9 1 9 2
13 2 13 15 9 13 0 9 1 15 0 0 9 2
19 2 13 1 15 0 9 1 9 2 0 9 7 13 15 9 9 7 9 2
7 3 13 9 9 2 2 2
12 1 9 11 11 2 5 12 2 12 2 12 2
1 11
5 9 11 13 0 2
11 13 3 13 0 9 3 1 12 2 9 2
19 7 3 3 1 10 9 4 13 9 15 0 2 15 15 13 1 10 9 2
22 9 15 13 1 9 11 11 11 2 15 13 11 7 13 1 9 10 9 7 9 9 2
20 11 4 13 1 0 9 2 7 3 2 7 10 9 15 9 3 7 13 13 2
48 13 15 0 9 1 9 9 2 3 0 7 3 0 2 0 0 0 9 2 7 1 9 7 9 3 13 1 9 9 3 0 9 11 2 11 2 11 2 9 9 12 7 1 15 9 0 9 2
7 15 3 13 1 9 12 2
34 9 15 13 15 2 16 13 15 14 9 2 16 15 0 9 13 2 7 9 3 1 10 9 13 3 12 9 7 0 9 4 13 3 2
5 3 13 9 9 2
7 3 13 9 9 2 2 2
8 15 3 13 3 7 1 11 2
5 0 9 12 2 12
27 13 2 16 1 9 9 11 12 2 9 12 1 10 9 4 15 13 2 13 15 1 0 9 2 1 11 2
16 7 7 3 4 15 3 13 1 11 2 7 4 13 1 11 2
19 9 15 3 13 14 1 9 12 2 3 13 13 13 9 10 9 1 9 2
19 1 9 12 1 0 9 13 0 9 1 10 9 0 9 3 1 0 9 2
45 13 14 9 1 9 2 0 9 10 9 13 2 10 9 2 3 15 2 16 13 1 11 2 13 15 1 15 0 9 7 9 1 10 9 2 7 3 3 7 1 0 2 13 0 2
46 13 1 0 0 9 3 0 7 1 3 0 9 0 7 15 0 7 0 9 3 1 9 12 2 3 3 9 1 9 2 3 4 13 9 1 9 1 0 11 1 11 11 7 11 11 2
38 1 10 9 1 11 2 3 1 11 2 4 15 13 0 0 9 2 15 15 1 15 13 2 3 0 9 2 0 2 0 7 9 0 7 0 9 0 2
25 10 9 3 15 13 2 13 15 2 16 13 1 11 2 13 4 2 13 9 7 13 4 13 3 2
23 7 3 11 2 11 13 7 13 9 2 13 3 3 1 10 9 2 2 16 4 13 9 2
9 16 15 2 15 13 2 13 13 2
10 7 3 9 3 3 15 13 9 13 2
13 1 9 13 10 9 2 0 0 9 7 10 9 2
8 13 1 15 0 9 7 9 2
24 9 15 13 2 14 15 10 9 3 13 2 2 2 7 9 14 15 1 15 3 13 2 2 2
30 1 9 4 1 9 13 1 11 7 3 4 15 13 1 9 1 0 0 9 1 0 9 7 3 15 3 13 2 2 2
13 14 3 2 1 0 9 0 9 4 13 1 11 2
37 1 12 9 15 3 13 10 0 9 9 11 11 7 1 9 12 0 2 9 9 1 0 9 1 9 11 7 3 1 9 11 2 11 2 11 11 2
10 1 10 9 0 4 13 3 0 9 2
61 3 3 1 11 3 1 9 13 9 13 15 1 9 9 11 2 1 15 4 15 3 13 2 7 15 15 14 2 3 1 0 9 10 9 2 7 3 15 13 0 0 9 7 9 11 11 2 15 15 13 13 2 16 15 13 9 1 10 0 9 2
17 7 1 15 4 15 3 13 2 16 4 1 15 16 9 3 13 2
25 13 15 0 7 3 0 9 2 14 0 9 2 1 15 4 13 3 0 2 7 3 4 15 13 2
14 10 9 1 11 13 1 11 11 2 0 9 0 9 2
19 13 4 15 1 11 1 9 12 2 3 3 13 1 0 9 1 0 11 2
16 13 1 11 2 1 9 13 1 9 11 7 13 7 3 3 2
17 13 1 11 1 11 2 1 9 15 13 12 9 7 13 3 9 2
28 1 9 7 9 1 11 13 9 3 2 16 15 13 1 0 9 2 9 15 13 1 9 7 1 9 13 9 2
30 1 9 13 9 0 2 9 2 9 2 9 7 0 9 10 9 7 3 4 13 1 10 9 2 15 4 1 9 13 2
7 7 3 9 13 9 9 2
8 13 15 9 7 0 9 0 2
4 13 15 0 2
12 1 0 9 13 1 9 0 9 1 15 3 2
8 13 0 9 7 13 15 3 2
6 9 1 9 9 13 2
28 2 2 2 1 11 13 9 7 9 1 0 9 2 3 2 1 9 2 4 15 13 7 13 0 0 9 11 2
10 7 3 4 15 13 13 1 11 12 2
17 9 11 12 2 0 15 13 1 9 0 9 0 9 9 3 0 2
35 13 9 2 0 9 11 11 2 15 15 13 13 3 0 9 11 3 0 1 9 7 9 1 9 7 13 15 1 0 9 7 1 9 9 2
29 0 15 3 13 2 13 3 3 16 1 9 1 11 2 13 3 10 0 9 7 0 0 9 7 13 15 0 9 2
33 13 15 1 9 7 1 15 1 0 0 9 7 9 1 9 7 9 7 1 9 7 9 1 15 1 9 13 2 16 15 3 13 2
15 13 1 10 9 0 2 7 3 7 3 2 16 13 9 2
28 9 9 0 9 2 10 10 3 7 3 0 9 7 9 1 0 9 13 13 7 0 9 0 0 7 1 9 2
10 3 9 15 13 1 11 1 9 0 2
27 0 9 15 13 9 9 11 11 2 9 11 2 0 9 3 16 10 0 9 2 7 15 13 11 3 0 2
15 0 9 0 13 7 0 9 13 1 15 13 1 9 0 2
19 0 9 15 3 13 1 0 9 2 13 10 9 2 0 9 13 1 9 2
6 13 7 10 9 0 2
10 13 15 0 9 2 15 13 3 0 2
13 7 7 4 1 11 13 0 9 9 1 0 9 2
16 13 1 9 0 9 2 16 4 13 11 13 7 13 10 9 2
18 9 11 11 7 10 9 1 0 9 13 1 11 1 0 9 10 9 2
11 0 15 13 1 0 9 10 9 7 9 2
7 13 15 0 7 0 9 2
18 3 15 3 13 3 2 16 15 13 10 0 9 7 3 7 0 9 2
15 11 15 3 3 13 2 13 15 1 15 7 13 1 9 2
29 3 15 13 1 0 9 2 15 9 13 1 9 2 7 1 15 15 9 12 7 1 10 9 11 12 2 0 13 2
5 13 15 12 9 2
6 1 9 13 16 9 2
8 10 0 7 0 9 13 13 2
26 1 9 0 9 1 9 9 4 13 9 1 0 9 9 2 9 7 9 2 1 9 7 0 0 9 2
12 9 4 3 13 7 1 9 3 13 2 2 2
22 3 4 15 13 1 11 2 11 1 11 1 10 9 11 11 2 15 13 1 0 9 2
10 13 4 0 9 1 0 9 1 9 2
15 7 3 4 15 13 2 16 0 3 0 9 1 11 13 2
19 3 15 3 13 13 2 7 15 15 2 7 15 15 13 7 1 10 9 2
5 13 13 15 0 2
17 3 4 13 11 7 15 13 2 13 4 13 1 0 0 9 11 2
21 10 0 9 2 3 15 13 1 0 9 7 0 9 15 13 1 0 9 1 9 2
46 0 9 13 0 1 0 9 7 9 2 13 15 13 9 2 3 13 1 15 15 2 9 2 9 2 9 7 9 9 7 0 9 3 2 1 15 13 0 9 7 9 7 9 7 9 2
6 1 9 15 13 0 2
13 7 13 3 7 0 7 0 9 2 9 7 9 2
11 15 13 9 0 9 1 0 7 0 9 2
57 9 3 13 3 0 2 3 0 9 2 0 9 1 9 2 0 9 2 9 2 0 9 2 9 2 9 2 2 7 3 15 3 13 9 2 9 1 0 2 3 16 15 13 2 16 13 0 7 3 0 2 7 3 13 7 0 2
10 3 13 2 3 15 13 2 1 11 2
25 16 4 13 0 0 9 1 11 2 13 4 15 9 13 3 7 3 13 7 9 2 15 13 9 2
52 13 15 12 9 2 13 15 9 1 9 2 1 15 15 13 1 11 2 2 7 13 0 13 9 9 9 2 13 15 1 0 9 2 13 2 7 16 15 9 3 13 2 15 15 13 7 13 15 15 12 9 2
6 13 15 15 1 9 2
42 3 15 13 12 0 9 2 13 15 9 2 15 13 9 2 1 11 15 0 7 3 0 9 2 2 3 15 15 13 9 2 13 14 3 2 7 13 15 7 0 9 2
30 1 9 2 3 0 2 15 13 9 9 2 7 15 3 1 9 13 7 13 2 16 15 13 0 7 13 15 15 13 2
8 9 13 13 3 9 0 9 2
11 9 13 0 1 9 2 13 3 7 13 2
7 13 15 3 13 1 9 2
8 13 15 13 3 0 7 0 2
23 15 1 15 13 2 3 9 7 10 0 9 2 9 2 9 2 9 7 3 2 15 13 2
6 13 15 9 0 9 2
13 3 4 1 10 0 9 13 2 13 4 0 9 2
15 3 4 3 13 2 1 10 9 15 1 10 0 9 13 2
4 0 13 15 2
4 9 1 11 12
63 3 10 9 1 11 13 0 7 0 9 2 3 1 9 0 10 9 1 11 1 0 9 0 0 9 2 1 15 13 7 9 1 9 0 9 7 9 2 13 9 2 9 9 9 7 10 9 13 1 15 3 3 2 7 7 16 3 3 3 2 7 3 2
18 0 9 1 0 9 15 3 13 2 7 9 0 9 15 1 9 13 2
26 13 15 0 9 2 7 9 2 2 9 10 9 2 3 9 2 11 2 11 1 11 7 9 1 11 2
7 3 1 9 1 9 13 2
40 13 15 9 2 3 15 3 13 0 9 0 9 7 9 9 11 11 2 11 2 9 15 7 1 9 1 10 9 1 11 13 7 1 9 13 1 10 9 9 2
30 3 4 13 1 11 1 11 2 1 9 1 9 1 11 2 1 9 1 11 7 1 9 2 10 9 15 7 9 13 2
17 9 15 13 1 9 1 0 9 9 2 7 14 1 9 0 9 2
10 13 15 3 2 16 13 0 2 0 2
28 1 9 4 9 2 15 15 15 13 2 13 2 16 13 2 15 13 7 15 13 9 2 16 13 1 9 9 2
17 16 15 1 11 1 15 13 7 1 9 1 15 13 1 15 13 2
66 7 1 0 9 2 7 13 4 15 2 4 13 2 16 13 1 0 9 2 13 15 2 15 15 14 13 2 1 9 13 1 9 2 13 13 9 7 1 9 15 13 9 1 0 11 2 1 9 1 15 13 2 16 15 13 2 7 13 15 3 3 1 3 0 9 2
18 3 15 15 13 2 0 13 0 9 1 3 0 7 3 0 2 2 2
31 7 13 4 3 15 2 7 3 13 2 9 7 9 2 7 10 0 9 2 15 15 13 0 9 7 15 0 9 2 2 2
6 9 13 1 15 13 2
46 0 9 13 3 1 10 10 9 7 9 2 3 3 3 13 10 0 9 7 3 4 13 2 16 15 15 15 13 1 0 9 1 9 2 16 9 13 3 7 1 10 9 15 13 9 2
50 10 9 0 9 2 15 1 15 13 2 3 13 7 13 2 13 3 1 10 0 9 2 2 2 2 15 13 1 9 10 9 13 7 13 15 1 10 9 2 14 3 2 16 4 13 7 1 10 9 2
27 15 15 13 2 13 3 2 3 4 13 1 0 9 2 7 1 15 15 13 3 14 7 14 13 2 2 2
39 13 4 3 2 3 10 9 13 13 2 13 15 1 9 2 7 3 15 13 13 2 9 13 2 2 13 13 14 3 2 7 1 9 15 13 3 2 2 2
19 16 13 2 12 9 2 12 9 7 12 9 2 3 13 7 13 1 9 2
10 13 4 7 9 2 3 3 3 2 2
23 16 4 10 9 13 1 0 9 1 9 9 2 9 3 2 15 15 13 2 13 2 2 2
35 16 1 9 12 13 1 9 0 9 11 11 9 12 9 2 9 11 11 7 9 0 9 2 2 15 13 3 1 0 9 2 13 0 9 2
5 13 15 3 13 2
36 3 1 10 9 9 11 11 2 1 15 15 3 13 3 9 9 7 15 13 1 9 16 10 9 7 9 2 13 1 9 13 13 1 0 9 2
23 3 13 13 16 9 1 9 2 10 9 9 7 11 2 11 13 7 13 13 3 0 9 2
32 11 2 11 1 9 13 2 16 13 1 3 0 9 7 16 15 9 2 3 1 10 9 3 3 13 2 10 9 13 1 9 2
21 11 2 11 15 3 13 9 10 9 2 9 13 13 14 9 2 2 7 13 0 2
20 13 9 1 9 2 9 1 9 2 13 9 9 7 9 2 0 13 0 9 2
20 1 0 9 7 9 15 11 1 10 9 13 0 9 2 0 3 14 1 9 2
21 9 2 12 9 2 13 0 9 7 13 0 0 9 2 12 2 12 2 12 2 2
32 0 12 9 10 9 11 2 11 3 13 7 13 1 9 0 9 10 9 2 1 0 9 13 9 7 1 9 0 0 9 2 2
6 10 9 13 2 13 2
14 13 15 0 2 10 9 1 15 2 1 15 2 13 2
13 1 9 9 11 11 13 9 1 9 1 9 11 2
4 9 13 11 11
3 9 11 11
30 0 9 2 3 13 0 9 11 11 1 11 2 9 2 13 1 12 2 9 3 0 2 16 3 4 13 0 0 9 2
15 1 9 12 3 13 9 11 2 11 13 0 7 0 9 2
12 9 2 12 9 12 2 13 1 12 9 9 2
1 9
10 9 13 7 11 2 0 9 0 9 2
11 1 9 15 13 1 0 9 7 0 9 2
16 1 0 9 13 9 0 7 0 9 2 1 15 7 9 9 2
12 9 1 9 7 10 9 1 0 9 2 13 2
1 9
6 11 2 0 9 0 9
16 9 1 9 13 0 2 13 15 1 0 9 2 13 11 11 2
4 11 11 2 11
1 9
39 9 3 2 16 1 9 12 13 0 9 2 1 9 2 3 13 1 9 9 1 0 9 2 15 1 0 11 3 13 9 2 15 15 1 0 9 13 9 2
15 9 13 3 3 2 13 9 2 7 13 1 15 0 9 2
7 9 1 0 9 7 9 2
29 1 0 9 1 0 9 2 3 1 0 11 1 0 9 13 0 11 2 0 9 13 2 16 15 10 9 3 13 2
18 15 2 15 1 11 13 9 2 7 10 0 9 2 13 13 0 9 2
30 16 11 2 11 0 15 3 3 1 11 3 0 9 2 7 3 2 13 9 9 2 15 10 9 1 12 9 13 0 2
14 16 0 0 9 13 1 0 3 14 1 9 1 9 2
37 16 13 15 1 9 3 2 16 13 7 15 13 2 13 3 3 14 9 2 15 1 0 9 1 9 12 13 1 10 9 9 1 11 9 11 11 2
7 1 11 15 13 7 13 2
52 16 0 11 15 0 9 13 3 1 0 12 9 1 3 0 9 0 0 9 2 16 9 2 9 7 9 2 15 3 13 3 9 0 9 2 13 3 0 1 0 9 7 13 9 2 1 11 15 13 7 13 2
9 9 7 9 1 0 9 13 9 2
6 6 2 6 2 6 2
25 13 0 9 7 9 2 16 4 13 0 0 0 9 13 1 9 0 2 0 2 0 7 0 9 2
22 9 9 1 9 0 9 7 9 2 15 13 1 0 9 13 1 9 9 2 13 0 2
13 9 0 11 13 1 9 9 1 0 9 12 9 2
22 9 11 11 13 10 9 9 9 0 0 9 2 3 9 7 3 3 3 9 0 9 2
14 11 13 1 10 0 7 0 9 3 10 11 1 0 2
29 3 16 3 3 13 9 9 2 7 7 9 1 0 7 3 15 0 9 2 13 3 0 9 10 3 14 0 9 2
17 9 9 13 1 0 9 2 3 15 0 13 13 9 9 7 9 2
17 16 4 13 2 3 14 1 0 9 2 7 3 7 3 3 0 2
7 1 11 15 13 7 13 2
10 13 15 0 0 9 7 13 15 0 2
20 16 13 11 3 9 0 9 2 13 15 2 16 15 11 13 1 0 9 13 2
4 16 3 11 2
4 11 13 7 13
12 0 0 9 2 11 11 11 2 3 13 0 2
16 16 0 9 0 9 13 1 0 9 1 9 0 9 1 11 2
27 13 3 3 1 9 0 9 2 16 15 1 9 9 3 13 9 7 13 1 0 9 0 0 9 1 11 2
14 1 12 9 11 13 9 2 15 13 9 13 0 9 2
14 0 9 15 3 13 1 9 9 1 0 7 0 11 2
8 13 13 7 1 0 0 9 2
23 4 13 0 11 2 0 9 2 15 13 9 7 15 14 13 1 12 2 9 0 9 11 2
11 11 13 0 2 16 15 13 3 0 9 2
8 9 13 3 3 0 2 13 2
31 1 15 15 7 3 13 2 13 9 2 16 16 11 13 3 1 12 9 2 3 3 1 9 3 16 9 1 0 9 9 2
19 15 13 1 15 9 2 16 9 3 13 3 0 2 13 1 0 9 9 2
12 0 13 15 7 1 9 9 7 11 2 11 2
16 15 2 15 13 9 1 0 9 2 13 12 9 9 0 9 2
7 15 3 13 9 2 16 2
11 9 13 1 0 0 9 1 0 9 0 2
11 9 9 0 9 1 0 9 13 0 9 2
10 11 13 2 16 3 13 9 15 13 2
21 13 15 3 1 0 9 9 0 11 2 1 15 13 0 9 1 0 9 1 9 2
21 3 1 9 15 12 9 13 1 0 9 7 13 11 2 15 13 3 14 1 9 2
3 9 1 9
27 1 11 2 0 1 0 9 2 3 13 1 11 11 12 0 0 9 2 13 1 15 3 12 9 2 2 2
50 16 13 3 9 0 9 0 9 11 11 2 15 1 0 9 0 11 1 9 1 0 9 13 2 16 11 13 9 1 9 11 2 9 0 9 2 2 3 13 3 0 2 16 9 13 3 1 9 11 2
26 9 0 11 15 1 0 9 1 11 13 12 5 2 1 0 11 12 5 2 7 1 11 3 12 5 2
39 7 16 10 9 13 13 0 9 2 16 9 9 13 0 16 1 9 1 0 9 2 13 1 9 11 11 11 0 2 16 9 0 11 1 0 9 11 13 2
30 3 15 11 13 13 0 9 2 3 15 13 7 0 9 2 0 0 9 2 7 0 9 2 0 15 1 0 9 9 2
17 1 0 9 13 9 9 0 9 2 0 9 9 2 0 9 9 2
14 15 15 13 9 9 11 11 11 2 0 2 0 9 2
4 11 13 7 13
22 0 9 12 0 0 9 11 11 2 12 9 2 11 14 13 2 7 3 1 15 13 2
15 13 15 15 3 12 1 10 9 2 1 15 13 1 9 2
23 11 13 9 3 15 2 1 9 1 0 9 2 15 9 14 3 0 1 0 9 11 13 2
29 13 15 9 7 13 15 1 0 0 9 2 3 2 15 3 15 9 16 15 7 3 0 2 3 13 2 13 11 2
19 3 15 13 3 0 2 3 0 2 16 3 2 2 2 9 2 9 13 2
8 14 2 13 0 9 0 11 2
21 13 0 2 16 10 9 13 9 1 0 11 7 9 2 0 9 2 3 13 3 2
12 13 3 9 2 16 10 9 13 10 0 9 2
8 9 2 1 15 13 2 13 2
23 13 2 16 10 9 2 15 13 1 0 0 2 0 9 0 2 13 1 0 9 3 0 2
10 15 2 15 13 9 2 15 13 9 2
15 15 2 15 15 13 2 15 13 9 7 9 9 2 13 2
20 3 3 13 13 2 16 13 10 9 7 15 3 15 13 2 13 15 14 3 2
29 13 15 3 1 9 2 15 13 1 9 9 7 1 9 3 3 0 9 15 3 13 2 3 15 13 1 9 11 2
4 13 2 15 13
11 13 15 3 3 0 7 9 13 14 9 2
17 1 12 9 0 9 13 0 13 0 9 2 13 9 11 11 11 2
10 9 13 16 9 0 3 1 9 12 2
22 9 2 0 9 1 9 12 15 0 0 0 11 2 13 0 2 0 7 3 0 9 2
11 13 2 16 9 3 7 13 2 15 13 2
29 13 9 2 13 1 9 13 0 9 2 13 0 9 2 7 16 4 15 13 2 15 15 4 13 2 13 9 11 2
45 1 9 11 2 9 2 15 13 9 0 0 9 11 7 3 13 9 9 1 0 0 9 2 15 15 3 13 1 0 9 3 0 2 15 13 3 16 0 9 0 1 0 0 9 2
16 1 0 12 9 0 9 11 15 1 9 0 9 13 12 9 2
9 12 1 9 13 1 9 0 9 2
19 13 3 1 0 9 7 13 1 15 16 1 0 9 2 15 13 0 13 2
6 15 15 3 6 13 2
34 10 9 13 2 16 9 1 10 9 13 1 9 3 0 2 7 14 1 9 4 13 9 2 15 15 1 9 13 1 9 9 1 9 2
15 9 3 13 7 9 1 0 2 0 9 12 2 12 9 2
6 9 1 11 13 3 3
21 1 15 2 15 13 9 1 9 2 13 3 11 2 0 9 2 15 13 10 9 2
21 9 1 11 1 0 9 13 16 0 0 9 7 13 1 15 0 2 13 9 11 2
18 13 15 1 0 9 0 9 2 1 9 9 2 1 9 9 7 9 2
8 3 13 7 9 1 9 9 2
4 13 3 3 2
11 9 11 13 2 16 4 15 13 9 9 2
7 7 15 13 3 9 9 2
11 1 15 2 3 13 9 2 13 0 9 2
12 11 2 16 0 0 9 2 13 13 14 9 2
7 13 4 15 1 9 9 2
13 13 1 15 0 7 13 1 10 9 2 16 0 2
11 14 2 15 14 2 13 0 2 3 0 2
22 3 3 15 13 9 2 15 0 11 3 13 2 7 15 15 3 13 2 13 15 9 2
4 14 2 9 2
2 0 9
12 0 9 13 12 1 0 9 0 9 0 11 2
27 13 15 7 3 0 9 0 9 11 11 2 15 3 13 10 9 1 11 7 13 0 9 7 9 0 9 2
24 2 3 3 3 2 16 9 15 3 13 1 0 9 1 0 11 2 16 0 11 13 1 9 2
20 3 4 3 13 7 11 7 11 2 16 4 3 9 10 9 13 1 9 2 2
15 10 9 15 13 9 9 11 2 0 1 9 9 0 11 2
24 1 15 15 12 9 0 11 13 2 16 9 13 0 9 2 14 14 1 9 11 13 0 9 2
14 16 9 0 1 9 15 9 13 12 9 2 12 13 2
20 13 15 0 9 2 13 11 11 1 9 2 3 15 1 15 13 13 1 9 2
24 4 15 13 3 3 2 7 9 1 0 9 15 13 2 16 13 9 0 1 0 9 7 9 2
2 0 9
12 0 0 9 13 1 0 0 9 3 10 9 2
26 9 1 9 9 2 11 11 11 13 1 9 16 0 9 2 9 1 9 2 0 15 1 0 9 9 2
9 9 10 9 9 13 1 11 11 2
25 1 0 9 15 11 11 13 16 9 2 3 15 3 13 1 9 3 2 16 1 0 9 13 9 2
28 7 16 4 13 9 2 13 0 2 16 13 0 9 3 1 15 16 0 9 2 13 15 11 11 1 10 9 2
22 0 0 2 0 9 13 16 0 9 2 15 13 10 9 1 9 3 1 0 0 9 2
14 0 9 2 15 13 15 0 2 15 9 13 1 9 2
14 13 7 0 2 16 9 0 2 0 9 13 9 9 2
20 1 0 9 13 3 0 2 16 4 15 0 9 1 9 13 2 13 11 11 2
17 13 15 2 16 13 3 3 3 13 2 3 7 3 15 9 13 2
8 9 9 1 15 13 0 9 2
15 13 3 0 2 3 15 9 0 1 9 13 1 0 9 2
18 16 15 4 13 2 16 3 1 0 9 2 7 16 15 9 3 13 2
11 13 0 9 2 15 15 16 0 9 13 2
34 13 7 7 15 2 15 15 9 0 2 9 3 13 2 13 9 11 2 15 15 1 0 9 13 13 9 2 7 0 9 1 0 9 2
3 9 13 3
39 3 16 13 0 11 1 10 0 9 2 9 2 7 0 9 11 3 16 0 0 9 0 11 2 13 7 0 11 2 16 9 9 1 0 9 2 0 9 2
18 9 11 11 2 12 9 2 13 2 16 15 0 9 13 1 11 0 2
15 7 16 9 1 0 13 9 2 13 4 15 0 11 0 2
18 0 11 15 13 9 1 0 9 2 1 9 1 11 2 3 15 13 2
6 13 0 9 7 9 2
26 1 9 9 15 3 13 2 7 14 0 15 3 13 3 13 1 10 9 2 1 9 13 0 9 9 2
17 10 9 3 0 13 2 16 1 0 9 13 3 12 9 2 9 2
10 11 11 2 0 9 2 13 0 11 2
21 1 9 2 16 13 9 7 1 3 12 9 1 9 9 16 0 2 13 2 3 2
3 13 15 3
17 1 0 9 13 14 1 15 2 16 3 9 13 1 9 10 9 2
13 13 0 9 2 15 1 9 1 9 9 13 9 2
8 13 15 16 9 1 0 9 2
14 9 1 9 15 3 13 0 2 7 14 15 13 3 2
12 3 15 13 2 1 9 2 9 2 1 9 2
7 7 3 13 3 1 9 2
10 3 15 13 7 13 2 15 15 13 2
9 13 15 2 16 15 9 3 13 2
12 3 4 13 2 16 15 12 9 13 0 9 2
12 13 12 9 7 13 1 0 9 0 2 0 2
15 15 1 15 7 3 13 7 13 15 2 3 3 13 9 2
12 15 3 13 10 9 2 7 15 15 3 13 2
6 1 9 13 3 9 2
29 13 15 2 16 15 13 1 0 11 0 2 7 16 13 2 16 4 13 1 0 9 7 16 15 1 15 0 13 2
18 13 2 16 0 0 9 13 1 0 11 0 9 2 15 13 14 0 2
10 1 10 0 9 13 9 11 3 3 2
23 1 9 3 13 2 16 4 13 3 0 2 16 4 9 2 15 13 2 13 9 0 9 2
4 9 15 3 13
24 11 2 12 0 9 1 12 0 0 9 2 13 9 1 0 9 0 2 13 15 13 0 9 2
8 3 0 9 9 13 3 13 2
25 0 9 2 0 0 9 2 13 15 15 3 7 0 9 1 0 9 1 11 2 7 13 14 0 2
24 7 14 2 13 4 3 2 13 2 7 9 13 3 0 2 13 3 0 2 7 3 13 9 2
7 2 7 1 15 0 9 2
16 7 3 1 15 13 15 0 2 9 2 3 9 9 2 2 2
8 15 3 9 14 13 2 2 2
25 13 9 1 0 9 3 3 2 14 16 9 11 2 15 13 2 16 1 15 3 9 1 11 13 2
5 9 9 15 13 13
16 9 11 13 3 9 2 16 15 13 2 16 11 13 0 9 2
18 13 15 9 9 0 1 12 0 9 2 15 15 3 13 1 12 9 2
39 1 10 9 13 1 0 15 9 0 9 0 9 9 11 2 1 15 15 0 11 13 13 3 14 12 5 0 9 0 0 9 2 1 12 5 1 9 12 2
15 15 13 1 12 9 0 9 2 16 9 9 13 9 0 2
41 13 2 14 7 9 2 16 15 13 0 9 2 0 9 2 15 13 13 1 9 1 0 0 9 2 3 13 2 14 3 2 3 2 16 13 11 0 1 10 9 2
21 3 2 16 15 3 3 4 13 0 0 9 11 1 3 0 0 2 0 2 11 2
14 13 14 9 7 9 0 9 2 7 3 10 0 9 2
2 9 9
7 11 11 13 3 0 0 9
5 11 2 11 2 2
29 3 0 7 3 0 1 9 16 1 0 9 13 3 1 9 0 9 11 11 2 11 2 9 9 9 1 9 12 2
11 9 9 1 0 9 7 9 9 3 13 2
26 1 11 4 9 13 2 16 4 1 9 1 0 9 9 0 9 0 9 13 1 9 3 16 9 9 2
13 9 1 0 9 4 3 13 13 0 9 0 9 2
22 0 9 4 13 9 13 9 10 0 7 0 9 2 1 15 15 1 11 13 10 9 2
47 0 14 3 13 2 16 4 9 9 13 0 0 9 9 2 1 0 9 13 9 3 2 13 0 9 0 9 0 9 2 16 4 3 13 12 9 1 9 9 2 15 4 1 9 3 13 2
32 11 1 11 13 9 0 14 1 0 9 2 7 3 1 9 0 2 9 13 1 15 10 9 7 9 13 2 16 13 1 9 2
19 10 9 13 2 13 9 1 0 9 11 2 1 10 0 9 15 3 13 2
21 1 9 2 0 0 9 0 2 0 2 11 2 15 3 3 13 13 10 0 9 2
1 9
1 9
9 15 15 13 2 16 15 13 11 11
27 0 0 9 13 0 9 0 2 7 3 0 9 2 3 13 9 2 9 2 2 16 11 13 7 11 13 2
13 1 15 15 13 13 3 2 16 0 9 2 3 2
19 9 7 9 13 3 9 0 2 1 9 15 1 10 9 10 9 13 13 2
20 1 0 0 9 0 9 0 9 13 9 0 9 2 16 1 9 0 9 11 2
10 7 3 3 13 9 2 3 15 13 2
23 13 1 9 1 9 2 3 15 0 9 13 9 9 9 7 13 0 9 2 15 13 15 2
10 15 9 13 2 13 15 9 0 9 2
8 16 15 13 9 2 13 0 2
7 0 13 0 7 0 9 2
7 1 0 13 0 7 0 2
14 15 7 9 10 9 13 7 0 2 3 13 9 0 2
15 9 0 15 13 13 3 2 1 9 9 2 1 0 9 2
9 10 9 13 9 2 4 13 9 2
14 7 15 13 0 9 2 13 0 7 9 2 3 3 2
17 7 13 9 7 9 2 0 0 9 7 0 9 13 1 9 9 2
16 3 3 13 9 2 0 7 3 2 15 13 0 9 2 0 2
11 0 9 1 9 10 9 13 9 1 9 2
17 7 3 2 16 13 3 13 7 13 3 3 2 16 15 9 13 2
19 1 10 9 13 9 2 3 0 9 9 0 2 0 0 9 16 10 9 2
21 9 13 9 1 9 3 3 2 16 15 13 0 9 1 9 0 9 2 1 9 2
19 3 15 9 13 9 1 9 1 0 9 7 13 1 9 2 0 0 9 2
7 7 13 1 11 0 9 2
16 3 15 3 13 2 7 13 3 0 9 0 2 0 9 0 2
10 0 9 1 10 9 13 1 9 0 2
18 0 9 15 3 3 13 13 1 9 2 7 15 13 1 0 9 0 2
13 9 9 1 10 9 13 3 1 10 0 0 9 2
11 13 1 9 3 0 11 2 3 3 0 2
17 16 4 15 13 9 1 0 7 0 9 2 4 13 12 0 9 2
18 1 9 12 1 9 1 9 0 2 1 9 12 1 9 1 9 0 2
14 15 15 13 13 9 2 13 13 3 12 9 9 0 2
16 7 15 13 0 9 1 9 2 13 12 9 13 1 9 0 2
10 3 3 15 13 13 1 9 1 9 2
25 1 9 0 0 9 15 9 0 9 13 1 0 9 1 11 7 3 13 2 16 13 3 3 0 2
6 9 13 1 9 12 2
13 9 3 14 1 0 0 9 0 9 3 13 9 2
41 1 9 0 9 1 0 0 9 1 0 12 0 9 15 0 9 13 1 12 9 2 1 0 1 9 1 9 11 11 2 11 7 1 9 0 2 15 13 1 11 2
21 1 9 9 1 9 2 3 2 1 9 2 0 9 9 9 1 0 9 13 3 2
8 3 15 13 1 0 0 9 2
12 12 2 9 12 4 9 1 0 9 9 13 2
2 0 9
5 0 9 1 9 9
2 11 11
5 10 9 3 2 2
5 9 9 3 0 2
9 15 2 15 13 2 15 3 13 2
7 3 13 2 1 15 13 2
30 3 3 15 13 7 9 9 1 9 7 9 9 3 0 14 15 2 16 13 1 15 2 7 7 15 2 15 9 13 2
30 10 0 9 0 9 2 15 15 3 3 13 1 9 9 9 2 15 13 9 9 7 14 15 13 0 9 1 0 9 2
6 16 4 13 3 13 2
10 7 14 2 15 3 13 15 2 2 2
9 9 9 12 2 9 13 1 9 2
7 9 13 2 15 14 9 2
20 7 15 9 3 13 2 16 13 13 1 10 9 2 7 15 3 13 1 9 2
3 3 9 2
31 9 0 9 15 1 9 3 13 7 15 15 13 13 3 0 2 16 16 4 13 1 9 2 13 4 1 9 1 0 9 2
23 13 3 16 15 3 13 7 14 1 9 9 13 9 3 1 9 2 16 9 3 13 13 2
6 3 0 11 2 2 2
4 14 2 9 2
20 9 1 15 2 16 9 1 9 13 3 9 3 0 2 3 9 0 9 13 2
10 13 3 3 2 3 0 11 2 2 2
14 13 2 13 0 9 2 13 1 9 7 1 15 3 2
11 15 15 7 0 0 15 9 1 9 13 2
31 1 0 9 7 13 2 16 11 3 7 1 9 13 9 0 9 0 9 2 9 9 2 2 15 15 13 3 1 9 11 2
20 0 0 9 7 9 11 13 1 0 9 10 9 3 1 0 7 0 9 9 2
18 1 9 0 9 2 3 15 13 3 2 15 7 13 13 1 0 9 2
25 9 2 15 15 11 1 9 0 11 13 2 13 9 0 9 7 10 9 0 11 13 3 16 11 2
29 16 0 11 13 1 9 9 0 9 1 10 9 2 3 15 13 1 9 2 11 1 9 11 13 9 1 0 9 2
17 9 9 9 2 9 0 2 13 7 13 9 2 15 15 13 3 2
19 9 9 13 1 9 9 9 7 1 9 9 13 9 2 1 15 9 13 2
9 0 0 0 9 3 13 2 13 2
7 3 0 9 13 0 9 2
3 13 15 9
14 0 9 1 9 9 13 0 9 11 11 1 11 11 2
33 3 2 16 4 1 9 12 16 9 13 7 1 12 9 13 1 11 2 13 15 1 0 11 1 0 9 2 13 3 9 1 11 2
10 1 15 13 7 3 9 2 9 9 2
21 12 1 0 9 1 9 13 1 10 9 9 2 15 13 3 7 13 15 1 9 2
37 3 16 0 11 2 7 11 11 13 7 3 13 9 9 0 9 2 14 1 0 9 9 2 2 7 3 15 13 9 13 15 1 9 13 9 9 2
20 3 1 10 9 13 9 0 11 1 9 11 11 2 9 7 3 9 15 9 2
11 12 15 3 13 1 9 7 9 13 0 2
20 11 11 13 9 2 3 15 13 1 0 11 13 0 9 2 7 11 0 9 2
25 14 9 15 11 7 10 0 9 13 2 9 13 2 13 2 13 9 0 9 7 13 1 0 9 2
5 15 1 0 9 2
26 16 14 1 9 10 9 13 2 13 15 11 2 16 15 2 15 15 1 9 3 13 2 13 1 9 2
11 13 15 9 12 7 1 9 13 0 9 2
31 11 11 13 1 0 9 1 9 11 7 0 9 7 3 1 15 3 13 7 0 9 2 15 13 1 0 9 1 12 9 2
9 1 10 9 15 11 13 9 9 2
20 13 15 3 2 16 11 11 9 1 9 13 9 9 2 13 1 9 7 13 2
11 13 15 7 9 2 15 15 3 9 13 2
15 13 15 9 9 0 11 2 15 9 14 10 0 9 13 2
7 3 15 13 0 0 9 2
3 12 9 9
20 11 15 13 3 7 3 10 9 13 1 10 12 9 12 9 0 9 0 9 2
23 0 9 15 13 1 10 9 9 1 11 11 1 15 2 16 4 15 13 13 1 9 9 2
15 13 2 0 9 15 1 9 12 9 1 9 13 1 9 2
24 0 9 13 3 10 15 9 2 1 10 9 12 2 1 0 12 9 2 7 13 15 0 9 2
25 16 1 12 9 3 13 1 9 9 0 9 11 11 2 13 3 9 0 9 2 1 15 11 2 2
22 3 7 4 9 1 9 13 3 2 9 9 13 3 3 14 3 0 7 0 9 9 2
22 11 13 0 9 1 9 9 2 15 13 16 9 9 1 9 2 7 13 15 1 9 2
26 9 2 15 13 0 9 0 11 2 15 13 3 2 11 13 9 7 1 0 9 15 13 1 0 9 2
3 9 1 9
15 0 9 13 1 9 12 0 9 11 11 2 11 1 11 2
3 14 15 2
11 16 0 13 3 14 9 9 1 0 9 2
17 10 0 0 9 13 1 0 9 2 15 13 9 7 15 15 13 2
13 3 0 9 9 9 13 1 9 0 9 1 9 2
21 10 9 15 7 3 13 14 1 9 2 3 13 9 9 1 9 0 0 0 9 2
10 1 15 15 13 12 1 0 9 11 2
10 3 13 1 0 9 1 0 0 9 2
26 11 11 2 11 2 9 1 9 2 13 9 2 3 1 9 13 0 9 7 3 3 15 1 15 13 2
20 13 2 16 15 9 3 13 1 0 9 2 15 13 0 13 3 10 0 9 2
12 0 2 15 15 15 13 1 9 2 13 0 2
17 1 9 0 9 13 3 0 9 0 9 12 9 10 9 9 11 2
16 3 15 15 3 13 2 16 1 15 3 1 9 15 3 13 2
15 10 9 15 1 0 9 0 11 13 9 1 9 11 12 2
13 7 9 13 10 9 9 7 9 7 3 0 9 2
15 3 2 16 0 9 1 9 1 9 9 13 9 1 9 2
22 7 16 0 11 10 9 13 2 9 15 3 13 7 11 15 1 9 13 9 1 11 2
3 9 7 9
11 3 12 9 15 13 9 2 9 0 9 2
21 13 15 1 9 12 2 3 11 11 11 13 0 0 0 9 2 15 13 13 9 2
3 13 14 2
7 15 7 13 2 13 9 2
17 9 3 3 13 7 9 13 3 0 2 1 0 9 13 3 3 2
14 13 15 14 1 9 12 2 16 15 10 9 13 13 2
32 0 9 1 0 9 11 11 2 13 10 9 2 13 1 0 9 9 1 0 9 9 9 7 9 2 10 9 9 13 0 2 2
17 13 15 12 9 2 16 10 9 13 13 3 2 16 13 3 0 2
18 1 9 2 3 10 9 13 9 9 2 13 1 9 3 0 0 9 2
9 16 3 0 0 9 13 0 9 2
4 9 7 9 2
24 9 9 12 4 3 13 15 9 0 0 0 9 2 0 9 3 13 14 15 1 0 9 9 2
12 3 15 2 1 15 4 9 13 16 0 9 2
12 15 0 9 1 10 9 13 3 14 0 9 2
5 0 13 9 0 2
18 9 9 9 2 15 13 16 9 1 0 0 9 2 13 3 3 0 2
12 13 3 1 0 2 7 0 2 9 1 9 2
9 10 9 13 3 9 9 9 11 2
15 3 3 13 0 9 9 2 1 9 10 9 13 9 15 2
16 0 0 9 0 9 13 7 9 9 0 2 15 13 0 9 2
15 13 9 1 9 2 10 9 2 9 9 3 13 0 9 2
12 1 0 9 9 1 9 3 3 9 3 13 2
28 1 9 0 1 9 9 15 9 9 13 2 16 1 0 9 13 9 0 9 2 7 7 13 10 9 3 0 2
18 13 1 15 2 3 3 13 1 0 9 9 2 7 3 1 9 9 2
10 7 3 15 13 3 1 9 10 9 2
29 13 4 15 3 2 16 0 9 0 9 2 15 1 9 1 9 3 0 13 1 9 2 13 9 9 0 1 9 2
12 9 3 9 13 13 2 9 7 14 2 2 2
2 9 9
6 0 9 2 9 7 9
3 9 11 11
2 11 11
5 13 0 0 9 2
3 3 13 2
13 1 9 9 0 9 3 13 12 9 2 3 0 2
19 9 4 13 9 11 7 9 13 9 11 2 13 9 9 7 13 15 3 2
14 1 0 9 15 10 9 13 9 1 9 1 0 9 2
7 13 15 1 11 11 0 2
16 9 2 9 2 9 7 9 9 7 9 9 11 11 13 9 2
5 7 13 3 13 2
28 11 11 13 9 7 2 3 2 13 1 9 9 9 1 9 2 12 1 12 1 9 0 7 0 9 10 9 2
20 3 13 15 13 7 9 2 0 9 1 9 2 15 1 11 13 9 9 11 2
14 9 11 11 2 13 12 1 11 2 15 13 9 9 2
17 1 11 2 11 7 11 13 1 9 9 12 9 10 9 1 11 2
5 11 11 13 9 2
28 0 9 0 9 7 3 10 0 9 2 0 9 11 2 11 2 11 2 11 11 2 11 11 2 7 11 11 2
8 13 4 15 1 9 1 9 2
4 13 4 15 2
17 7 10 9 13 16 9 1 9 2 15 1 10 9 13 7 3 2
13 3 2 3 2 1 0 9 2 7 1 9 9 2
7 7 4 3 9 9 13 2
8 13 14 9 10 9 7 9 2
5 3 13 2 2 2
2 1 11
6 11 13 9 0 9 2
35 3 4 13 1 9 0 9 1 9 2 1 15 4 0 9 13 2 1 11 2 11 2 11 2 11 2 7 13 3 2 16 11 15 13 2
17 13 16 11 0 9 15 1 15 2 14 15 2 15 13 10 9 2
39 9 2 16 15 13 16 9 10 9 13 9 10 0 0 9 2 13 1 9 2 1 0 9 2 7 13 2 16 11 4 3 3 3 1 15 13 2 2 2
3 1 0 9
15 10 9 13 9 9 9 11 2 9 2 15 13 0 9 2
13 0 9 0 1 9 11 15 13 3 1 10 9 2
19 7 13 15 3 0 9 2 7 0 9 10 9 16 11 11 7 11 11 2
14 11 11 3 13 2 3 1 10 9 15 13 2 2 2
17 13 2 16 12 15 13 1 0 9 7 13 15 13 7 0 9 2
14 10 9 13 9 0 9 7 0 0 9 3 3 13 2
15 13 15 0 2 16 11 11 4 3 13 7 9 2 2 2
16 1 9 12 13 1 9 7 1 0 9 13 9 9 0 9 2
15 13 2 16 1 0 0 9 7 9 13 1 9 7 9 2
27 3 15 9 13 1 9 9 9 11 2 7 15 4 3 3 13 2 7 16 4 3 3 15 13 2 2 2
3 1 0 9
21 11 15 1 10 9 13 9 9 9 2 15 9 7 9 1 9 7 3 10 9 2
12 3 13 9 1 9 14 12 7 12 9 9 2
13 13 15 10 0 0 9 2 16 3 13 0 9 2
44 1 12 0 9 1 0 15 13 10 9 2 0 9 7 1 9 10 9 0 9 2 9 1 9 2 15 4 3 7 3 13 2 10 0 9 1 11 9 12 2 2 2 3 2
9 15 13 9 9 2 10 0 9 2
3 1 0 9
7 13 12 0 0 2 9 2
10 12 1 9 12 7 0 1 9 12 2
10 3 4 15 15 13 0 2 0 9 2
9 7 1 0 9 13 14 10 9 2
13 10 9 13 9 2 14 3 15 13 3 1 9 2
9 13 9 1 9 15 13 3 0 2
7 9 13 0 9 13 9 2
9 9 9 13 15 0 16 9 9 2
8 1 9 9 13 0 0 9 2
8 0 9 7 9 13 0 9 2
16 9 2 15 13 9 1 9 2 13 1 15 0 9 0 9 2
11 14 13 9 1 0 2 9 0 2 0 2
9 7 0 9 13 0 9 2 2 2
2 1 9
5 3 15 13 9 2
6 9 13 0 9 9 2
22 13 1 15 0 9 9 2 16 13 16 9 2 3 13 1 0 9 9 2 3 9 2
19 9 9 13 1 15 2 16 13 2 15 13 9 2 16 13 0 9 9 2
29 3 13 0 9 7 9 1 9 2 1 9 2 1 9 2 1 9 7 9 2 1 0 9 2 1 9 0 9 2
13 1 15 9 13 13 2 15 3 13 2 0 9 2
8 7 3 13 7 0 9 9 2
27 1 15 3 13 0 9 0 0 9 2 7 3 9 10 11 11 7 11 11 11 13 0 9 16 0 9 2
37 13 2 14 13 1 15 2 7 15 4 15 13 1 10 12 9 13 0 9 2 16 4 13 0 9 2 0 2 16 13 0 9 7 9 0 9 2
10 13 4 15 13 0 9 0 0 9 2
9 13 9 2 15 4 9 13 3 2
5 1 9 7 0 9
17 1 15 4 9 13 13 15 0 2 3 3 1 9 2 16 9 2
8 1 9 9 13 9 15 0 2
29 3 9 2 15 13 1 10 0 9 2 15 13 1 9 1 0 9 7 13 15 13 1 10 9 3 1 10 9 2
19 3 2 3 13 9 2 13 15 1 9 10 0 0 9 3 1 9 9 2
17 3 13 0 0 9 2 7 15 13 3 0 2 0 9 10 9 2
25 14 16 1 9 2 0 7 0 9 13 15 2 3 4 13 1 9 2 3 4 13 1 0 9 2
16 9 1 9 2 9 1 9 7 9 9 0 9 7 0 9 2
17 9 2 3 4 13 1 9 1 9 2 13 15 9 9 2 2 2
12 15 0 1 10 9 13 3 9 2 9 9 2
8 3 1 10 0 9 13 9 2
17 1 9 9 2 2 2 1 9 7 1 0 9 9 7 0 9 2
26 11 2 1 3 0 9 2 0 9 2 11 11 11 2 12 2 12 2 2 0 9 2 9 7 9 2
19 1 9 9 1 9 12 2 12 13 0 9 7 3 0 9 0 0 9 2
22 10 9 11 11 15 13 1 10 9 7 0 9 9 11 7 9 2 15 13 9 9 2
6 13 1 12 9 2 2
11 1 9 2 9 11 11 4 13 9 9 2
21 13 4 1 9 2 15 15 3 13 2 3 1 10 0 9 9 2 3 13 9 2
9 13 15 0 2 0 2 0 9 2
13 1 0 9 2 15 15 4 13 2 13 12 9 2
17 9 2 9 2 9 9 7 9 7 3 9 1 0 9 1 9 2
27 10 9 13 7 13 0 9 13 14 0 9 2 7 3 0 2 1 15 0 2 7 3 0 0 10 9 2
29 13 12 9 3 2 3 13 1 9 1 9 7 15 12 9 13 1 9 1 9 1 12 9 1 9 7 0 9 2
24 15 15 13 2 16 4 15 13 0 9 2 0 13 9 2 9 1 9 2 15 15 13 13 2
21 11 3 13 2 16 9 10 9 13 1 9 7 0 9 9 13 1 9 0 9 2
8 7 15 3 13 1 9 9 2
9 15 13 1 0 11 15 3 0 2
22 3 15 15 13 13 0 9 9 1 0 9 2 3 1 15 13 1 11 7 1 11 2
21 3 13 9 2 13 1 15 2 16 4 9 7 1 0 7 0 9 13 10 9 2
16 7 15 15 16 9 3 13 2 13 15 9 3 0 7 0 2
21 1 10 9 15 3 13 13 0 9 1 9 9 10 0 9 7 9 10 9 0 2
2 1 9
33 9 7 9 9 15 13 3 2 7 15 13 2 16 0 9 13 1 9 2 13 0 2 13 9 9 9 2 0 9 7 0 9 2
31 14 2 13 15 2 16 13 1 9 9 2 10 9 3 3 13 2 13 0 7 13 14 1 0 9 2 1 15 3 13 2
27 7 1 10 9 9 7 9 9 16 9 0 9 9 2 9 7 9 4 13 1 10 9 0 9 7 9 2
3 1 9 9
27 13 15 2 16 1 15 2 16 4 15 9 13 9 2 13 13 0 9 16 9 2 15 15 13 13 9 2
15 3 0 9 9 2 0 9 2 9 13 15 14 3 0 2
9 0 9 2 3 0 2 15 13 2
29 9 13 13 3 0 2 0 2 7 1 10 9 7 3 3 9 0 9 2 13 13 15 0 2 15 3 4 13 2
11 7 13 0 9 0 9 2 9 2 9 2
20 13 9 7 9 2 9 7 9 2 13 0 7 0 2 0 7 0 2 2 2
29 16 9 13 3 3 9 0 9 2 3 15 0 2 15 9 13 13 2 13 13 1 15 15 10 10 9 7 9 2
12 16 15 13 2 13 13 9 7 9 10 9 2
7 1 15 13 0 9 11 2
19 11 13 0 9 1 0 9 13 9 2 7 3 0 9 0 9 7 9 2
5 11 15 13 13 2
4 1 9 7 11
42 1 12 1 10 0 0 9 2 1 11 2 3 9 10 0 9 2 13 1 15 0 0 9 1 9 2 0 0 9 2 9 2 9 16 9 9 2 0 9 2 2 2
23 13 4 15 13 2 7 3 4 13 2 16 15 13 1 11 2 1 11 11 2 1 11 2
48 6 2 11 3 7 13 1 0 9 13 2 13 15 10 9 2 15 3 13 1 0 0 9 2 7 15 15 13 2 16 9 13 0 0 9 2 0 0 9 2 9 2 15 13 3 16 9 2
3 9 7 9
8 3 4 13 13 9 1 9 2
12 3 2 7 3 2 16 15 10 9 13 0 2
14 0 9 4 15 13 16 9 2 16 4 13 0 9 2
20 15 12 9 0 9 15 13 13 9 9 2 9 0 9 7 3 0 9 9 2
7 0 9 13 14 0 9 2
9 3 13 2 13 15 16 1 9 2
7 15 13 9 0 10 9 2
14 10 9 13 9 14 3 2 16 15 13 1 10 9 2
30 9 13 1 15 0 9 2 7 16 0 16 10 9 0 2 7 3 15 13 2 16 13 9 1 9 13 0 2 2 2
6 9 3 13 9 9 2
32 13 13 7 10 9 2 1 15 1 9 13 2 13 7 10 9 2 16 15 15 13 3 2 13 13 15 2 15 15 13 9 2
41 9 13 3 0 9 2 7 3 1 9 3 0 2 3 3 2 3 13 1 9 9 9 7 9 9 1 0 9 13 1 9 0 9 3 0 2 16 4 15 13 2
6 13 0 0 0 9 2
3 3 13 2
13 1 9 9 0 9 15 3 13 12 9 2 2 2
31 11 11 13 3 1 9 0 9 7 11 7 11 0 9 11 1 0 0 9 2 1 9 13 9 1 9 0 9 7 9 2
25 13 3 1 0 9 11 9 0 9 1 0 9 2 9 11 11 7 9 7 9 9 3 2 2 2
1 9
7 9 0 9 2 12 2 2
2 11 11
21 9 1 12 9 2 15 13 9 9 2 1 15 4 1 0 9 10 9 9 13 2
23 3 4 13 1 9 9 2 15 13 0 3 1 0 9 9 7 9 1 9 7 1 9 2
15 1 10 9 9 15 10 9 3 13 11 2 11 7 11 2
7 3 13 9 1 11 9 2
13 1 9 9 13 1 9 3 12 2 9 12 2 2
19 1 12 2 9 12 7 12 2 9 12 4 13 0 7 15 15 13 3 2
17 16 4 3 13 0 12 2 9 12 2 13 0 9 12 2 2 2
11 1 9 9 0 13 7 13 15 0 9 2
19 1 0 9 13 2 16 13 1 0 9 2 1 9 7 9 13 0 9 2
20 11 13 10 9 1 9 12 2 7 0 9 13 1 9 12 1 1 9 12 2
20 1 9 1 9 12 13 7 9 0 7 1 9 12 15 13 0 9 11 11 2
16 3 0 13 1 0 9 1 9 1 9 12 2 13 3 0 2
11 0 9 13 3 12 0 9 9 1 9 2
12 2 12 9 13 3 13 2 9 13 3 0 2
13 1 12 0 0 0 9 13 9 13 1 0 9 2
28 0 9 13 9 0 2 15 13 10 0 9 2 0 2 9 12 9 12 2 0 2 9 12 9 12 9 12 2
14 0 13 0 9 1 9 9 7 13 15 9 1 9 2
4 9 13 15 2
11 7 1 0 9 9 13 13 9 1 9 2
25 1 9 11 2 11 2 0 1 0 11 1 9 12 2 13 0 9 9 1 0 9 1 10 9 2
10 0 13 1 9 7 13 12 2 2 2
6 4 0 13 3 13 2
12 0 9 12 2 9 12 4 13 3 1 9 2
19 1 0 9 15 13 0 1 9 11 2 11 2 0 1 11 1 9 12 2
4 3 15 13 2
9 15 0 13 9 9 7 9 2 2
6 0 4 13 9 12 2
7 2 3 13 9 0 9 2
10 1 0 9 13 13 3 12 2 2 2
8 2 0 9 13 9 0 9 2
18 0 15 13 13 7 9 9 7 9 9 1 9 12 1 10 9 2 2
2 13 9
12 13 9 9 2 7 7 13 9 9 12 0 2
12 13 1 15 7 9 14 1 12 2 9 12 2
5 13 15 0 9 2
5 9 1 0 9 2
7 9 0 9 3 13 3 2
5 1 11 4 9 13
2 0 9
2 11 11
16 13 4 3 3 0 9 7 13 4 15 13 10 3 0 11 2
13 7 11 13 1 9 9 9 2 7 15 15 13 2
57 1 11 13 14 9 2 3 9 2 9 2 9 7 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 7 14 15 3 2
37 16 4 15 15 13 9 7 13 12 9 0 0 9 3 1 9 0 9 2 13 4 9 10 9 13 1 9 2 16 0 9 13 0 9 3 0 2
15 15 15 7 1 0 9 13 1 15 0 2 3 3 0 2
5 13 4 3 11 2
7 3 15 15 13 10 9 2
28 13 2 14 15 15 1 15 2 16 15 13 0 9 2 3 13 3 2 16 15 3 13 1 0 9 9 0 2
9 0 9 4 15 13 13 1 9 2
14 9 15 1 15 13 1 9 2 7 13 9 1 11 2
25 9 13 7 1 9 7 1 9 2 9 1 9 2 9 13 9 11 1 0 9 9 2 9 2 2
34 9 15 1 15 13 1 9 1 11 2 3 4 9 13 2 2 9 13 0 9 2 9 7 9 1 9 2 9 1 0 9 2 9 2
11 9 13 1 9 2 3 16 9 7 9 2
11 9 13 3 0 9 2 15 13 0 9 2
24 9 13 1 0 9 9 2 16 9 13 3 0 2 3 7 11 15 15 13 7 13 3 9 2
21 1 11 15 0 11 3 13 7 9 9 2 9 2 7 1 15 11 16 9 2 2
25 1 0 9 9 13 11 9 2 3 9 1 9 2 7 15 0 13 1 11 2 3 3 1 11 2
12 7 3 0 2 3 4 15 13 15 1 11 2
19 9 13 1 9 2 9 1 0 9 2 9 1 0 9 2 9 1 9 2
27 9 13 1 9 2 9 1 9 2 9 1 9 2 9 1 9 2 9 1 9 2 7 9 13 1 9 2
11 10 9 10 9 13 0 2 0 3 0 2
13 3 14 13 1 0 11 2 3 15 3 13 9 2
14 9 13 13 1 9 0 0 2 15 15 13 11 11 2
10 7 9 13 3 0 9 11 11 11 2
14 9 13 14 9 0 9 2 10 9 15 13 16 9 2
7 3 3 7 9 9 13 2
20 9 13 16 9 13 3 12 1 11 2 16 9 13 14 9 2 7 3 2 2
10 9 13 1 0 9 7 13 3 9 2
60 1 9 15 13 11 2 1 9 12 15 15 13 1 0 11 1 11 7 1 10 9 1 9 0 9 11 2 7 9 15 1 15 13 1 10 9 1 0 11 7 11 2 3 16 15 15 3 13 2 14 4 1 15 11 15 13 3 0 2 2
28 9 9 13 1 9 2 7 3 13 1 9 1 11 2 10 9 13 12 9 0 9 9 7 1 15 13 9 2
22 9 15 13 3 12 1 11 2 16 0 2 11 9 3 13 2 7 16 1 15 13 2
16 9 9 15 13 11 2 3 9 2 13 15 3 1 9 3 2
24 9 0 15 13 11 2 9 13 11 1 9 2 9 13 1 11 2 9 13 9 1 0 11 2
58 1 10 9 2 16 13 9 7 9 2 13 0 7 0 3 15 2 9 2 9 2 9 2 9 2 9 2 13 13 15 0 9 2 3 16 9 2 9 2 9 2 9 2 9 2 9 2 14 3 7 9 2 3 1 0 9 2 2
27 0 9 15 13 13 2 16 1 0 9 13 1 15 3 2 7 1 15 13 9 3 0 9 3 3 0 2
18 13 2 14 7 3 13 9 1 9 9 2 13 13 9 1 0 9 2
6 15 15 3 3 13 2
5 9 1 9 7 9
2 11 11
20 1 11 15 12 2 9 13 0 9 9 11 11 2 3 3 0 9 0 9 2
32 0 9 9 15 13 1 9 9 9 1 9 7 9 2 1 15 15 10 9 2 9 7 9 0 7 0 13 1 0 0 9 2
56 1 12 9 2 3 13 9 15 3 13 1 0 9 2 15 13 3 16 13 2 16 10 9 13 0 9 7 16 15 10 9 13 14 3 1 9 10 9 2 7 7 3 1 9 2 1 15 13 9 12 9 2 9 7 9 2
22 11 11 2 3 0 9 9 7 9 0 9 1 0 9 1 11 2 13 1 0 9 2
22 13 15 0 9 3 15 2 3 15 1 9 9 13 2 3 1 15 15 0 9 13 2
14 1 0 9 13 7 1 9 1 9 15 9 0 9 2
29 13 1 9 1 9 11 14 1 9 9 12 2 3 4 3 13 2 16 10 9 7 9 11 11 2 0 9 9 2
15 13 15 12 2 9 12 1 11 1 9 0 9 11 11 2
17 1 9 9 0 0 9 15 13 1 0 9 1 9 9 7 9 2
35 1 9 15 7 3 13 2 16 1 9 9 12 4 1 9 13 0 2 0 9 1 15 0 0 9 2 3 1 10 0 7 0 0 9 2
13 1 0 9 0 9 3 13 3 0 0 0 9 2
12 0 9 13 1 0 0 9 1 0 9 9 2
18 11 15 13 11 2 7 14 15 2 0 9 0 13 1 10 0 9 2
23 9 1 9 3 14 3 13 9 2 3 9 10 0 9 2 15 13 9 1 0 0 9 2
23 9 1 0 0 9 0 11 7 9 11 15 10 9 13 14 3 9 9 2 7 7 3 2
13 0 9 11 11 13 7 13 3 13 14 3 0 2
30 15 13 9 2 15 13 10 9 10 9 2 0 1 15 1 0 9 2 0 9 9 1 0 9 13 2 11 2 12 2
6 11 0 2 11 12 2
18 0 9 0 11 2 12 2 7 12 2 9 2 11 12 7 12 2 2
19 13 3 0 13 1 0 9 2 7 13 0 13 1 0 9 9 0 9 2
31 9 2 7 3 9 1 9 2 2 0 9 3 3 11 2 11 3 13 0 9 0 9 0 10 9 1 0 7 0 9 2
28 0 9 1 12 2 9 9 11 11 9 1 9 7 9 13 1 0 9 9 0 9 7 0 0 7 0 9 2
15 0 9 13 9 11 11 2 9 11 11 7 9 11 11 2
10 13 15 3 0 9 7 0 0 9 2
19 2 2 2 9 15 13 2 3 13 15 2 1 9 2 15 13 0 9 2
7 1 9 11 11 0 11 11
11 9 13 3 13 9 2 13 1 9 11 9
7 11 2 11 2 11 2 2
51 13 15 0 2 7 16 3 14 0 2 13 3 9 9 11 11 2 11 2 1 9 11 2 16 13 0 2 16 4 9 0 0 7 0 9 13 9 10 0 0 9 9 0 11 2 15 15 13 1 0 2
14 15 13 3 0 2 16 9 13 9 13 9 2 13 2
31 9 9 1 10 0 9 4 7 1 11 13 13 3 3 13 2 16 1 9 0 9 3 0 0 9 13 13 0 9 9 2
26 1 9 9 11 11 11 13 9 2 16 4 9 13 13 10 9 2 15 15 13 1 0 2 3 0 2
48 1 9 11 2 15 0 9 11 11 13 2 16 15 9 11 13 1 0 9 9 0 9 0 9 11 11 11 2 11 13 2 16 16 1 11 13 1 10 9 2 7 13 1 0 9 15 9 2
17 9 9 13 3 0 9 7 15 3 13 13 9 9 11 1 0 2
20 0 9 4 1 15 13 2 16 4 15 9 13 13 0 9 7 3 15 13 2
38 3 3 1 9 11 2 11 7 11 2 11 2 11 2 3 13 1 9 9 11 9 9 11 2 11 2 11 2 7 9 9 11 2 11 2 11 2 2
13 9 3 13 9 2 16 13 1 9 9 13 9 2
6 0 9 13 9 13 0
14 13 11 7 11 2 16 4 3 13 13 2 13 11 11
6 11 11 2 11 11 2
24 3 1 11 13 10 9 2 13 1 9 0 9 2 7 1 0 9 2 1 9 1 9 9 2
10 3 13 1 15 0 7 0 9 9 2
15 0 9 7 9 15 1 15 13 16 0 9 7 0 9 2
23 0 9 13 9 3 0 2 7 9 3 1 9 3 13 10 2 16 4 15 13 1 15 2
20 9 7 9 13 7 9 2 15 9 13 1 9 10 9 2 3 15 13 3 2
11 13 13 10 9 2 16 4 15 13 13 2
16 9 9 13 1 9 1 9 7 9 2 7 15 13 0 9 2
8 1 11 13 1 9 7 9 2
13 9 13 9 2 15 4 3 13 2 16 4 13 2
21 9 13 15 2 15 4 13 3 3 2 16 4 13 13 3 9 15 7 10 0 2
45 13 4 10 9 1 9 2 3 4 13 2 16 15 13 9 1 9 2 3 4 15 15 13 15 7 15 13 1 9 2 7 3 4 13 1 9 2 16 4 15 15 15 13 13 2
19 1 15 0 2 1 9 9 2 9 2 0 9 2 13 0 0 9 13 2
7 2 9 0 9 2 2 2
15 9 13 9 2 15 4 1 0 9 3 3 13 2 2 2
15 13 4 2 16 9 0 9 13 12 1 0 9 1 9 2
23 15 2 16 13 0 9 7 9 2 13 9 2 7 3 4 15 13 0 13 1 0 9 2
11 13 1 0 9 2 3 1 9 7 9 2
13 1 10 9 3 13 9 1 0 2 9 1 9 2
31 13 9 2 16 4 11 13 13 10 9 2 7 15 1 10 9 2 16 13 1 9 9 2 15 13 9 7 13 3 13 2
23 2 11 11 3 13 2 16 4 15 0 13 1 9 9 11 2 7 15 4 0 9 13 2
13 13 3 9 9 2 16 4 15 13 10 0 9 2
8 13 3 0 13 15 1 9 2
7 3 15 3 13 13 9 2
18 13 15 9 2 16 4 15 13 9 1 10 9 2 13 4 1 15 2
16 16 4 7 15 13 11 11 1 15 2 13 4 16 1 9 2
19 16 9 3 13 2 16 15 9 13 1 0 9 2 3 9 13 13 9 2
13 7 15 13 9 9 1 10 9 2 16 15 13 2
7 2 3 4 13 9 9 2
2 9 2
6 2 3 4 13 11 2
18 13 15 9 2 15 15 13 9 2 9 7 9 2 7 13 10 9 2
16 2 1 9 13 0 10 0 9 10 9 2 15 13 10 9 2
15 1 10 9 0 11 15 3 13 2 16 4 15 13 13 2
7 13 4 13 9 1 9 2
16 10 9 4 13 7 10 0 9 2 7 1 15 15 3 13 2
17 11 11 3 13 1 0 9 1 11 2 16 15 13 0 9 11 2
19 1 15 9 13 10 0 9 2 16 13 1 3 3 0 9 9 3 0 2
3 13 9 2
10 1 15 2 16 4 3 13 3 13 2
10 9 15 13 2 15 1 15 13 0 2
4 13 13 13 2
15 2 1 10 9 13 0 13 9 1 9 1 11 7 11 2
15 1 10 9 13 13 16 1 0 9 1 0 7 0 9 2
9 13 15 9 2 9 1 12 0 2
13 11 13 3 0 9 1 15 2 16 13 3 13 2
7 11 13 13 1 0 9 2
12 15 2 15 13 0 13 2 4 13 0 9 2
13 13 15 2 16 4 12 0 9 13 1 0 9 2
25 16 13 15 9 0 2 13 15 13 2 15 13 10 9 2 3 15 4 13 1 9 7 1 9 2
6 3 3 13 13 9 2
19 3 15 13 0 9 2 7 15 13 13 9 2 3 2 13 4 13 12 2
4 12 0 9 2
13 2 1 9 0 9 4 13 0 0 9 11 0 2
19 13 15 1 0 9 9 11 2 3 4 15 13 13 1 0 9 10 9 2
31 13 15 13 1 15 2 16 0 9 13 9 1 0 9 0 9 2 7 1 15 2 16 14 0 0 9 13 13 3 0 2
9 13 15 3 3 7 9 1 11 2
24 13 15 3 0 9 1 2 9 1 9 2 15 13 0 9 13 3 2 7 3 13 15 0 2
7 13 15 9 1 0 9 2
17 11 13 13 0 9 1 9 9 2 9 2 9 2 9 7 9 2
15 3 13 15 1 12 9 2 15 3 13 12 0 10 15 2
19 13 15 16 9 0 9 2 16 9 15 2 16 0 9 13 9 13 0 2
18 2 1 0 9 9 13 9 0 9 11 16 9 0 2 0 0 9 2
7 13 10 9 9 1 9 2
19 13 9 7 13 7 3 9 1 9 2 16 15 1 0 0 9 13 13 2
12 0 9 13 3 9 1 9 7 1 0 9 2
14 0 13 1 0 9 9 2 14 15 0 0 2 15 2
26 0 9 11 13 3 0 9 2 16 15 1 9 9 13 0 9 9 2 1 15 13 9 7 9 9 2
12 15 13 2 7 10 9 13 1 0 9 9 2
11 2 7 1 9 9 13 9 9 13 0 2
19 9 13 1 0 1 15 7 13 15 9 2 3 7 16 13 1 0 9 2
15 13 4 9 2 15 4 15 13 3 2 16 4 13 9 2
16 13 9 2 15 15 3 13 1 15 2 16 13 0 9 9 2
16 9 13 0 9 7 16 13 15 9 2 13 15 9 0 9 2
14 2 0 9 4 13 1 10 0 9 0 9 2 2 2
14 13 15 9 1 0 9 2 15 13 0 13 15 0 2
30 13 9 2 15 15 13 13 0 9 2 7 16 13 3 14 9 1 9 2 13 0 9 9 2 16 4 10 9 13 2
22 10 0 9 1 0 9 13 9 13 15 1 9 2 15 1 10 9 13 9 1 9 2
22 1 10 9 13 3 0 2 9 13 0 9 1 9 2 16 4 15 3 13 1 9 2
17 10 9 4 15 3 13 3 3 2 16 4 15 0 9 13 0 2
30 2 10 0 9 1 0 3 1 9 0 9 2 15 15 1 15 3 13 0 9 2 13 1 0 9 1 0 0 9 2
7 13 1 0 11 9 0 2
10 11 13 3 3 0 9 2 9 13 2
25 13 4 2 16 0 9 2 1 11 0 3 3 12 12 9 2 13 1 15 0 9 16 0 3 2
9 13 15 13 0 9 2 0 9 2
20 16 13 10 0 9 13 16 9 1 10 0 0 0 9 2 3 13 0 9 2
2 11 11
2 15 15
2 15 2
2 15 2
3 13 9 2
6 13 9 2 0 13 2
3 13 9 2
6 9 9 2 15 14 2
2 13 2
6 15 9 2 9 9 2
8 9 13 15 9 1 9 9 2
2 15 2
3 13 13 2
3 9 9 2
9 1 9 11 1 11 2 11 12 2
7 9 9 1 9 2 12 2
6 6 2 10 0 9 2
4 15 13 11 11
12 9 2 0 2 12 2 13 0 9 7 9 2
31 13 1 9 9 2 1 9 3 1 0 9 2 1 0 9 0 9 1 11 2 2 13 0 9 1 9 0 9 7 9 2
11 13 1 0 9 2 11 2 11 2 2 2
10 1 11 11 13 3 0 9 0 9 2
23 13 9 2 3 9 13 10 9 7 0 9 2 15 2 1 0 9 9 7 9 2 2 2
20 13 15 15 0 9 2 7 15 13 0 2 16 10 9 13 14 15 1 15 2
34 3 13 9 2 15 0 9 13 1 9 2 7 0 9 15 13 2 15 2 0 2 13 2 13 15 2 13 2 1 9 13 2 2 2
28 3 0 9 15 7 3 13 2 1 9 15 13 0 9 2 1 15 3 13 0 2 15 7 1 15 15 13 2
8 3 3 13 15 7 1 15 2
22 10 9 4 15 3 13 2 16 10 0 9 1 0 9 4 13 0 13 1 10 9 2
45 16 3 13 3 3 0 13 1 0 9 2 0 1 10 0 9 2 13 4 3 2 3 4 15 3 13 2 16 2 2 2 2 7 16 15 0 15 4 10 9 3 13 1 9 2
24 13 4 3 13 0 9 10 9 15 2 15 15 15 3 13 2 7 3 15 13 1 10 9 2
17 13 15 2 16 4 1 15 13 2 7 13 15 3 3 15 0 2
16 9 1 9 2 16 7 1 0 9 2 3 13 1 0 9 2
10 3 7 3 13 3 0 9 2 15 2
6 15 13 9 3 0 2
13 13 15 3 3 7 1 0 15 15 13 3 13 2
13 14 0 15 13 3 9 13 3 7 3 1 15 2
13 16 0 9 0 15 13 3 14 1 12 0 9 2
36 7 0 15 7 9 0 15 13 10 9 3 13 7 9 7 9 13 15 1 10 9 15 3 13 15 0 15 2 15 13 15 3 0 2 2 2
36 11 13 2 16 0 13 2 13 2 14 15 3 3 2 7 13 15 13 2 16 13 0 9 2 16 13 0 15 2 15 13 14 15 1 15 2
27 7 6 3 2 13 2 14 15 3 10 0 15 2 3 15 7 13 2 16 4 15 15 13 3 1 9 2
14 7 7 3 13 9 14 9 0 9 1 15 7 15 2
27 1 0 15 2 0 15 1 9 7 0 15 0 9 2 1 15 13 14 2 14 9 2 3 3 0 9 2
6 0 9 11 7 0 9
2 11 11
15 9 2 0 2 12 2 13 9 2 9 2 13 1 0 9
10 9 9 10 0 9 13 9 1 9 2
34 3 3 13 2 16 13 9 2 15 13 16 9 0 9 7 15 15 3 13 13 1 9 1 9 2 9 9 7 9 0 9 2 9 2
8 3 1 9 7 1 10 9 2
11 9 13 1 10 9 9 9 1 0 9 2
15 9 15 3 13 3 13 2 7 3 13 3 13 9 9 2
6 7 15 13 1 9 2
39 15 13 3 9 2 15 9 12 13 0 9 7 0 0 9 11 11 11 2 12 2 1 9 11 7 10 0 9 2 15 0 9 13 1 0 11 9 11 2
41 9 2 16 4 13 1 10 9 13 3 3 2 7 1 0 9 13 10 0 9 0 2 0 9 4 3 3 1 9 10 0 9 13 9 1 9 7 4 13 3 2
33 0 9 13 1 15 2 16 14 0 13 3 0 2 16 4 15 13 13 0 9 0 9 2 9 9 11 2 0 9 7 0 9 2
27 7 16 9 13 13 10 0 9 14 1 9 2 13 15 13 7 1 9 1 0 9 13 1 3 0 9 2
27 15 13 7 1 0 9 0 15 1 0 0 9 2 1 15 15 11 11 3 13 1 9 0 9 0 9 2
26 13 7 0 7 0 9 2 16 11 11 13 0 9 1 0 9 1 11 7 16 0 9 1 9 13 2
23 13 15 3 3 9 2 3 10 0 9 10 0 0 9 1 0 9 0 11 13 0 9 2
16 13 3 0 9 2 7 0 0 9 3 13 13 1 0 9 2
7 7 1 9 3 3 14 2
5 9 13 3 0 2
24 9 9 13 13 0 9 10 9 1 0 7 0 9 1 9 9 2 9 2 9 9 7 9 2
14 0 9 13 13 2 7 0 9 7 0 9 11 13 2
16 9 1 9 0 13 3 2 13 0 9 1 9 9 0 9 2
9 3 15 13 2 14 7 3 13 2
27 7 13 9 9 2 16 13 1 9 9 7 16 13 0 9 13 9 0 9 7 9 2 15 9 3 0 2
26 14 13 3 13 2 7 3 15 9 13 2 3 2 3 2 15 1 15 2 3 3 7 3 3 2 2
21 7 16 15 3 3 13 7 16 15 1 15 13 0 0 9 2 13 1 9 13 2
16 7 9 1 0 9 7 1 11 2 3 13 15 1 15 13 2
25 9 15 13 2 15 15 13 2 0 9 3 13 15 1 9 2 13 7 16 3 13 1 0 9 2
17 9 13 12 2 0 0 9 13 1 9 1 0 9 2 7 0 2
5 11 15 14 13 2
28 0 9 3 13 1 0 9 11 11 2 3 13 9 9 7 9 2 0 9 7 9 1 9 9 2 9 0 2
31 7 13 3 3 0 2 15 13 7 1 9 9 11 7 0 9 2 3 9 2 9 2 3 15 13 9 1 0 9 9 2
20 1 0 9 13 1 9 0 9 7 0 0 9 2 15 14 13 10 0 9 2
13 16 1 9 15 4 0 0 9 13 1 0 9 2
24 3 16 1 9 0 9 2 9 2 9 2 3 7 13 4 1 9 12 9 9 11 11 13 2
10 11 11 11 2 11 7 10 0 9 2
14 13 11 2 11 12 2 16 12 2 9 9 0 9 2
4 13 11 11 2
10 12 9 2 9 13 2 9 12 9 2
3 1 0 9
6 11 11 2 11 12 2
3 13 15 2
27 0 9 0 9 2 0 9 1 9 11 2 2 15 13 16 9 2 9 7 9 3 2 13 0 9 9 2
3 13 9 2
6 11 11 2 10 9 2
27 1 0 9 3 0 9 1 9 11 13 0 9 1 9 2 3 13 1 9 1 0 9 0 9 11 11 2
12 13 11 1 9 11 11 7 11 11 2 11 2
9 11 11 2 0 9 1 0 9 2
9 9 13 9 0 9 9 1 9 2
8 13 0 9 11 11 1 11 2
9 11 11 11 2 9 1 0 9 2
19 9 9 0 9 13 1 9 1 9 11 1 9 2 9 7 9 10 9 2
7 13 11 11 7 11 11 2
6 11 11 2 0 9 2
3 9 9 2
3 9 9 2
2 9 2
3 6 3 2
26 0 2 0 9 12 9 9 2 12 2 12 2 0 9 1 11 7 11 13 0 9 1 9 11 11 2
3 0 0 9
1 9
2 11 11
9 0 9 15 3 13 11 0 9 2
23 1 0 9 2 0 11 11 2 13 1 3 0 9 1 9 0 9 9 7 0 0 9 2
44 9 2 15 9 9 13 11 11 1 0 9 0 0 11 1 0 9 2 13 9 9 0 9 1 0 9 2 7 1 0 9 2 16 3 13 1 11 9 2 13 13 9 9 2
11 1 0 9 13 11 2 7 9 11 11 2
27 1 15 0 9 0 9 15 13 3 3 0 2 7 13 7 11 9 1 9 9 2 0 11 1 11 2 2
24 13 15 1 15 3 9 9 0 9 11 2 11 2 11 2 11 9 9 2 11 1 11 2 2
39 9 11 2 15 0 9 3 14 1 9 13 2 15 1 10 0 9 13 7 3 3 13 2 16 0 0 9 13 13 9 0 9 2 16 15 9 3 13 2
37 16 2 16 11 13 2 1 10 9 13 0 9 11 11 1 9 16 0 2 7 0 9 2 13 4 3 0 2 16 4 15 9 13 0 9 9 2
6 1 15 13 3 13 2
25 9 7 13 9 0 2 3 10 0 9 9 11 9 2 15 13 2 9 9 2 0 0 11 2 2
37 13 4 15 15 3 2 13 11 3 2 16 13 2 16 11 9 13 2 1 3 0 9 13 9 0 9 2 10 9 13 13 2 2 2 9 11 2
39 16 13 13 2 13 15 0 9 10 9 2 15 0 9 12 1 0 11 9 3 9 13 2 16 3 15 13 1 9 9 7 9 2 7 1 0 0 9 2
17 13 4 1 9 1 12 9 2 13 3 1 9 10 9 11 11 2
54 0 9 2 16 15 1 9 13 2 3 13 9 2 16 9 10 0 2 16 3 0 0 9 13 0 9 7 16 0 0 9 1 15 9 4 13 1 0 9 7 9 9 15 0 2 16 1 15 13 7 13 9 0 2
5 0 9 13 0 9
2 11 11
13 9 2 0 2 12 2 13 9 2 13 1 0 9
18 11 11 11 2 12 2 13 1 10 9 0 9 9 1 9 0 9 2
15 1 10 3 3 0 0 9 4 13 10 3 0 0 9 2
23 9 0 9 7 10 9 0 0 9 2 10 0 9 13 9 11 2 13 3 13 0 9 2
15 7 16 0 9 1 9 9 9 2 7 16 0 9 9 2
19 1 0 9 0 9 15 13 9 9 7 9 0 9 1 0 9 0 9 2
33 1 11 13 0 13 9 3 16 9 9 2 9 2 1 15 13 2 15 3 13 2 15 13 1 9 11 2 16 13 1 9 9 2
10 14 16 0 9 9 13 9 0 9 2
24 0 9 13 11 1 9 9 16 9 9 2 10 0 9 13 13 1 9 15 2 15 3 13 2
30 15 2 15 13 9 9 1 10 9 2 13 7 13 1 9 0 9 16 1 0 9 15 2 15 13 0 2 13 11 2
19 15 0 13 7 1 9 1 9 10 0 9 2 13 2 14 15 16 0 2
27 0 0 9 13 13 1 0 9 1 0 9 7 0 9 2 15 9 3 13 0 7 9 3 3 13 9 2
18 0 9 13 9 3 0 0 9 7 11 13 1 15 9 0 0 9 2
54 13 3 2 16 0 9 13 4 13 3 0 9 1 0 0 7 0 9 3 1 12 0 9 2 3 9 2 16 13 3 3 0 9 1 9 15 2 15 13 10 9 2 7 9 2 16 13 13 0 9 1 10 9 2
16 11 13 13 1 9 0 7 1 15 0 9 2 15 3 13 2
13 3 13 13 0 2 0 2 7 1 15 0 9 2
12 3 3 13 9 0 9 2 9 0 9 9 2
20 10 9 13 2 3 16 3 11 2 3 15 0 16 13 9 1 10 9 0 2
53 13 0 9 16 11 2 15 13 2 15 13 1 9 2 13 9 7 9 2 1 15 9 13 2 13 15 7 1 15 0 2 3 16 13 10 9 13 7 13 9 9 2 16 15 15 15 13 13 3 1 0 9 2
15 1 0 9 13 0 3 9 9 0 9 13 3 0 9 2
25 10 9 0 7 0 9 13 13 16 9 1 9 0 9 0 9 1 9 7 9 0 9 0 9 2
33 1 9 9 0 9 13 7 10 9 13 3 1 9 0 9 1 0 7 0 9 1 10 0 9 2 7 3 7 1 10 0 9 2
23 1 10 9 15 13 13 2 16 1 9 0 9 15 13 0 9 0 9 9 0 7 0 2
11 11 11 11 2 0 9 7 10 9 12 2
6 13 11 2 11 12 2
4 13 11 11 2
10 12 9 2 9 13 2 9 12 9 2
6 0 9 1 9 0 15
2 11 11
15 9 2 0 2 12 2 13 9 7 9 2 9 9 0 9
46 1 9 2 3 15 1 10 9 13 9 0 2 0 9 2 13 15 1 15 1 0 9 12 1 0 9 10 9 2 9 9 2 11 2 0 9 7 9 11 11 2 12 2 12 2 2
32 0 9 2 15 1 0 11 13 15 16 9 0 9 2 13 1 9 0 15 0 9 2 1 11 1 11 1 11 11 2 2 2
20 3 15 1 10 9 0 0 9 13 2 13 13 2 16 13 0 9 0 9 2
42 16 11 1 10 9 3 16 11 1 9 0 9 7 10 9 7 11 1 9 1 15 13 1 0 9 0 9 2 0 9 9 13 9 9 0 9 1 9 3 3 0 2
26 13 1 15 15 9 0 15 2 13 1 15 0 7 0 9 7 0 0 9 13 3 1 0 0 9 2
29 0 3 13 2 16 15 2 15 13 3 3 1 15 7 14 1 15 2 13 1 10 9 3 0 9 1 0 9 2
11 11 13 7 1 10 9 0 9 2 9 2
17 10 0 0 9 3 13 1 9 1 0 0 9 0 9 0 9 2
6 13 1 0 9 9 2
13 1 9 1 10 0 9 15 13 1 0 0 9 2
35 3 1 0 11 11 7 0 11 11 13 1 9 12 0 0 9 2 11 1 11 2 2 15 15 13 0 9 3 1 9 9 1 10 9 2
16 1 9 1 0 9 9 3 13 11 7 11 0 9 1 9 2
34 0 0 9 4 7 9 13 3 16 9 0 2 1 9 1 11 3 13 9 2 15 4 13 1 3 0 2 7 3 13 10 0 9 2
21 16 7 13 11 11 1 9 2 0 9 1 0 0 9 15 11 13 9 0 9 2
17 3 9 9 2 0 1 11 9 12 2 13 0 9 1 10 9 2
14 1 3 0 2 14 3 0 9 13 0 9 0 9 2
32 9 9 2 1 15 9 13 1 15 15 2 13 0 2 0 9 2 1 15 0 2 16 13 3 9 0 0 9 16 0 9 2
34 9 2 1 15 9 13 2 13 9 11 2 9 2 9 2 2 11 2 0 9 2 7 11 2 9 0 7 3 0 9 0 9 2 2
45 1 0 9 9 7 1 9 0 9 2 1 9 9 7 1 3 0 9 0 9 15 13 0 9 1 0 0 9 2 10 9 1 9 7 9 1 9 1 9 13 0 9 0 9 2
19 1 0 9 9 13 11 0 9 1 10 0 9 2 0 9 0 9 9 2
22 1 15 3 13 14 15 9 2 9 15 15 2 2 7 7 9 9 2 3 9 2 2
36 9 1 15 15 7 1 0 9 9 7 9 13 1 10 0 9 0 0 9 2 1 2 2 2 9 15 2 15 4 13 3 9 7 9 9 2
7 13 13 0 9 1 9 2
32 1 0 0 9 13 15 15 15 13 13 9 9 9 3 15 13 7 15 15 1 15 13 2 1 15 13 1 0 9 3 0 2
28 3 4 13 10 9 13 1 9 7 13 15 1 15 2 3 1 0 9 11 11 2 16 1 3 0 0 9 2
30 9 10 9 13 3 12 1 0 9 0 0 9 2 3 13 1 0 9 13 9 2 15 3 3 13 1 0 9 9 2
6 11 11 2 9 9 2
17 13 11 2 11 12 2 1 9 0 9 9 7 0 9 1 11 2
8 13 11 11 2 9 11 11 2
11 12 9 2 9 12 9 2 9 12 9 2
6 9 9 13 9 1 9
9 11 2 11 2 11 2 11 2 2
21 1 0 9 9 1 11 12 13 0 0 9 0 9 0 9 0 9 9 0 11 2
43 1 9 11 2 16 9 9 13 2 13 11 11 2 9 9 0 11 2 15 13 9 9 2 1 9 9 2 15 13 1 0 9 2 4 13 9 2 3 4 10 9 13 2
33 14 3 3 2 16 4 13 9 1 15 2 16 9 13 1 9 2 7 13 4 15 2 16 9 2 0 9 2 4 13 0 9 2
8 3 4 13 0 9 1 9 2
28 1 11 13 0 9 1 9 9 9 11 13 1 0 9 11 9 2 10 9 7 4 9 13 1 0 9 9 2
37 0 9 3 13 0 9 2 16 15 3 13 2 13 4 9 9 4 3 13 2 11 7 1 10 9 14 13 14 14 13 2 16 15 3 3 13 2
21 9 11 2 11 2 11 2 13 2 16 3 13 9 2 15 4 4 9 13 11 2
14 11 7 1 9 10 9 11 2 11 10 0 9 13 2
14 9 9 4 14 13 2 7 16 4 9 13 0 9 2
24 1 11 2 11 2 11 2 4 1 0 9 13 14 9 9 11 2 7 3 4 13 3 1 2
20 9 11 2 11 2 11 2 13 2 16 10 9 13 2 16 4 4 9 13 2
8 13 7 2 16 15 11 13 2
4 9 9 13 3
11 10 9 13 1 11 9 7 3 13 1 11
7 11 2 11 2 11 2 2
15 0 9 15 13 1 11 9 0 9 9 9 11 2 12 2
21 1 0 9 15 1 9 2 0 9 12 9 13 3 0 9 1 11 12 2 12 2
27 1 9 3 13 10 9 1 0 0 9 9 1 11 0 9 2 0 9 12 2 12 7 12 2 12 2 2
27 11 3 1 9 1 9 13 3 9 2 7 3 1 9 1 11 2 12 2 12 2 13 1 9 14 0 2
5 0 9 13 11 2
6 11 2 11 12 2 12
22 12 1 12 9 13 0 9 1 11 11 7 11 1 9 1 9 3 3 0 9 11 2
22 11 2 15 13 12 9 7 12 9 2 13 2 16 15 13 14 10 0 9 1 9 2
6 1 9 15 3 13 2
29 11 11 13 1 11 2 15 12 1 11 2 7 9 7 9 2 15 1 12 9 13 1 0 9 9 2 13 13 2
8 1 9 15 13 2 13 11 2
29 1 9 0 9 1 0 9 1 0 0 9 1 12 2 9 3 13 1 9 15 0 7 9 4 1 9 9 13 2
10 1 9 9 1 9 4 13 11 11 2
24 1 12 9 13 9 11 7 16 1 12 2 9 13 11 0 9 2 4 1 9 9 3 13 2
26 1 0 0 9 1 12 2 9 15 13 1 0 9 13 11 2 15 15 13 0 9 0 2 0 9 2
12 7 12 1 12 0 0 9 3 13 1 9 2
8 7 1 0 12 15 11 13 2
21 13 15 3 15 7 16 3 15 13 1 0 9 2 13 15 15 0 9 9 11 2
27 9 1 9 13 1 12 2 9 11 2 10 9 1 0 9 0 0 9 1 9 13 9 9 1 12 9 2
25 3 10 0 9 13 11 1 0 9 9 1 0 9 9 2 15 15 13 14 0 0 9 11 11 2
6 11 2 11 12 2 12
10 0 9 7 0 9 15 13 9 9 2
33 1 15 13 0 9 11 2 15 11 1 12 2 9 13 1 9 3 2 16 13 4 13 1 9 2 13 1 15 1 0 9 2 2
14 11 4 3 1 0 9 9 13 1 12 9 1 9 2
8 3 3 7 13 13 9 9 2
28 15 11 1 12 2 9 13 0 9 1 0 0 9 7 3 16 13 0 9 11 13 2 13 11 9 1 9 2
19 9 9 3 13 13 9 11 2 15 13 1 11 1 12 0 9 1 11 2
7 9 11 7 13 0 9 2
16 9 13 2 16 0 9 11 1 12 2 9 13 1 9 0 2
29 0 9 15 3 13 1 0 9 1 12 2 9 2 3 11 13 11 2 15 9 9 3 13 0 11 2 9 2 2
23 9 15 13 13 2 7 1 12 2 9 13 1 0 9 11 11 7 13 1 9 0 9 2
23 11 13 1 9 12 9 7 15 2 15 1 9 12 2 12 13 2 13 15 0 16 11 2
21 10 0 9 13 1 9 1 0 9 3 0 2 7 4 13 1 0 9 12 9 2
21 13 0 2 16 4 13 13 9 1 9 2 15 13 1 15 3 3 2 13 11 2
4 11 13 12 9
8 1 9 0 0 13 7 11 11
8 0 9 11 1 0 11 11 11
57 0 9 11 2 12 2 9 11 2 13 1 0 9 9 1 11 11 2 12 2 2 12 9 7 1 9 12 2 12 2 12 2 12 2 12 2 12 2 12 2 2 12 2 12 2 12 2 12 2 12 2 13 1 9 0 0 2
36 1 0 12 9 13 1 0 11 7 0 0 11 11 2 15 1 11 11 2 12 2 9 11 2 13 10 9 2 12 2 12 2 12 2 12 2
35 1 0 9 0 9 13 11 2 11 7 11 2 1 15 4 9 9 13 3 2 7 1 0 9 11 2 0 0 9 11 7 0 9 11 2
11 0 9 15 13 0 9 11 7 9 11 2
27 10 9 1 11 13 11 16 0 2 1 9 1 11 15 13 1 9 0 9 2 15 0 9 13 0 9 2
28 0 12 9 7 0 9 13 1 9 7 3 13 9 2 16 15 15 13 2 0 9 3 1 15 13 0 9 2
24 13 4 9 2 16 4 13 12 0 9 1 12 2 12 3 1 9 9 2 3 15 15 13 2
37 3 4 7 13 1 9 2 16 4 15 15 13 3 2 13 1 9 11 2 15 13 0 9 0 9 9 7 3 13 12 2 12 7 12 2 12 2
25 1 10 9 4 15 13 9 1 9 2 13 15 9 7 13 9 2 13 15 1 12 0 9 11 2
13 0 9 13 0 9 2 7 1 0 9 15 13 2
21 3 15 13 0 9 0 2 15 11 3 13 2 16 13 10 9 1 12 2 12 2
30 3 4 15 3 13 7 0 9 9 13 2 13 11 2 15 1 12 9 7 12 9 13 3 10 0 9 1 0 9 2
30 1 12 9 4 1 0 9 9 12 13 1 11 2 1 15 4 13 12 2 12 1 9 7 12 2 12 1 0 9 2
20 7 7 1 9 13 13 2 3 1 11 4 13 12 1 11 2 13 15 11 2
23 10 9 13 1 9 2 15 13 3 2 3 15 0 9 3 13 2 9 11 2 12 2 2
15 1 9 1 11 15 11 1 9 1 11 13 9 1 9 2
12 3 4 1 15 3 13 2 7 4 15 13 2
20 13 15 15 13 0 9 2 1 9 15 13 11 2 13 7 14 0 9 11 2
13 1 9 1 11 11 2 12 2 2 15 13 3 2
20 15 3 1 10 9 12 2 9 1 0 9 11 13 11 11 2 12 2 2 2
28 1 10 9 9 13 2 16 4 15 13 9 2 16 4 15 13 2 7 3 4 15 13 2 13 15 13 2 2
19 3 13 1 10 9 0 2 13 1 9 12 2 12 2 12 2 12 11 2
19 7 16 1 0 9 13 12 2 12 2 7 1 10 9 14 1 9 13 2
45 16 11 13 0 9 3 9 2 11 11 2 12 2 2 15 15 1 0 9 9 11 1 12 2 9 13 7 13 1 9 7 12 9 12 2 12 2 12 2 12 2 12 2 12 2
25 9 9 1 9 0 9 2 3 4 13 12 2 12 1 0 9 7 13 4 13 1 12 2 12 2
17 7 11 3 13 7 1 0 9 13 9 9 2 13 1 9 11 2
21 16 3 14 1 9 1 11 13 3 2 3 3 13 9 2 7 9 15 9 13 2
39 11 3 13 0 9 3 1 0 9 1 11 11 2 12 2 2 2 1 15 13 14 1 9 12 2 12 2 12 2 12 2 12 2 12 2 12 2 12 2
46 11 11 2 12 2 2 15 13 9 1 9 1 11 2 12 2 2 2 12 2 12 2 12 2 12 2 12 2 12 2 16 1 0 0 9 13 12 2 12 7 13 9 12 10 9 2
14 1 11 13 9 1 9 2 15 13 2 15 15 13 2
26 1 11 4 13 3 13 7 1 15 13 9 2 7 1 0 9 4 1 15 13 3 2 13 9 11 2
13 3 4 3 13 1 15 2 16 4 13 11 13 2
38 16 4 15 3 1 9 1 0 0 9 13 9 12 0 9 2 16 13 1 12 9 2 13 15 0 11 11 2 12 2 2 3 2 16 13 0 9 2
50 3 1 9 15 7 13 11 13 1 9 2 16 1 0 9 15 1 0 11 13 7 1 9 2 1 12 2 9 3 13 1 0 11 11 2 12 2 2 12 2 12 2 12 2 12 2 12 2 12 2
13 11 11 13 9 9 1 0 0 2 16 13 11 11
2 9 11
7 9 7 9 1 9 1 11
2 11 2
16 9 9 0 9 1 9 12 1 11 13 9 1 9 7 9 2
15 13 1 15 1 10 0 9 1 11 0 9 0 0 9 2
10 9 0 9 7 3 13 9 9 11 2
25 9 4 13 1 11 9 3 3 0 0 9 2 12 9 9 2 12 9 9 2 12 9 9 2 2
24 9 2 0 9 0 0 9 2 13 3 13 1 3 16 9 9 7 3 1 11 13 0 9 2
19 12 0 9 13 13 14 1 9 9 1 11 2 13 15 0 9 0 9 2
9 1 9 13 9 3 0 12 9 2
26 1 0 9 9 7 0 9 11 13 14 1 15 2 3 15 10 9 13 1 9 1 11 1 9 12 2
24 9 11 11 2 11 2 11 13 2 16 10 9 13 13 3 0 9 11 1 9 12 1 11 2
9 11 2 3 2 13 10 0 9 11
2 9 11
6 0 9 13 1 9 9
13 11 2 9 13 10 9 2 9 13 1 9 13 9
5 11 11 2 0 11
10 0 9 1 0 0 15 13 0 9 2
22 0 0 9 11 1 9 13 2 16 10 0 9 4 13 10 3 0 9 1 0 11 2
44 14 16 4 11 13 1 9 13 1 9 1 10 9 0 9 11 2 7 10 9 13 13 3 1 9 11 11 1 0 0 11 2 7 1 0 0 0 11 2 9 0 0 11 2
28 0 0 9 0 9 15 7 13 9 1 9 2 7 7 13 3 9 7 0 0 9 13 1 9 3 0 9 2
34 15 0 13 1 15 0 2 15 9 13 2 3 15 9 13 1 9 9 2 13 9 0 9 11 11 2 15 0 9 13 1 10 9 2
27 1 9 1 9 1 11 13 1 9 10 9 7 1 0 9 9 15 13 2 2 3 15 2 11 2 2 2
23 3 1 9 13 13 2 16 3 13 1 9 10 9 2 15 9 1 0 9 11 11 13 2
8 14 2 1 15 13 0 9 2
9 15 15 3 13 2 3 13 13 2
16 3 15 13 2 16 4 13 3 1 9 2 7 15 15 13 2
9 9 15 15 13 2 9 4 13 2
29 0 9 4 7 13 1 10 9 7 9 4 13 2 13 15 11 2 16 15 13 9 2 7 16 15 13 1 9 2
27 7 9 9 1 15 2 16 9 13 1 10 9 10 9 2 15 1 15 7 3 1 10 9 3 13 9 2
20 3 15 1 11 9 13 1 0 9 0 9 7 3 10 0 9 13 0 9 2
64 13 4 11 2 16 4 0 13 15 2 15 15 4 13 14 0 9 2 7 1 15 4 13 9 1 11 1 9 2 13 11 1 9 10 0 9 9 2 0 0 9 13 1 9 1 9 9 0 7 1 9 1 9 16 9 13 9 2 16 11 13 1 9 2
15 7 1 0 9 9 11 11 15 13 1 0 9 9 11 2
22 11 3 3 13 13 1 9 2 7 12 9 15 3 13 2 16 15 13 0 0 9 2
24 3 1 9 0 9 2 9 1 9 1 9 7 0 9 9 1 9 1 9 2 1 15 13 2
11 3 1 9 13 0 15 9 3 0 9 2
27 15 13 13 1 9 7 13 2 16 16 0 9 13 13 7 13 9 2 3 4 15 13 13 7 0 9 2
23 13 2 16 9 15 13 1 0 9 2 9 2 16 9 13 9 2 15 13 1 0 9 2
19 7 16 13 1 9 2 9 15 13 13 1 9 2 14 15 13 10 9 2
9 13 15 2 16 15 13 10 9 2
24 9 13 13 9 7 1 15 2 16 4 1 9 13 0 9 1 9 0 9 2 13 15 11 2
18 3 13 0 9 3 9 2 7 1 10 9 3 3 13 10 0 9 2
21 9 3 13 9 1 0 9 1 0 11 1 9 2 0 9 7 3 0 9 9 2
21 11 11 2 15 13 13 2 16 1 9 13 0 9 2 15 3 1 12 9 13 2
13 1 9 11 15 0 2 7 1 9 13 7 11 2
18 7 15 9 2 16 4 15 13 9 1 9 2 13 9 9 1 15 2
36 11 15 3 13 10 0 9 11 11 2 11 11 15 13 1 0 1 11 7 11 11 3 0 9 0 9 13 13 1 9 0 11 1 0 11 2
25 9 1 9 3 13 11 11 2 15 15 13 1 15 13 0 11 1 11 7 13 3 12 2 12 2
14 13 15 3 13 2 16 1 9 9 3 9 3 13 2
42 7 15 15 13 7 13 2 15 4 15 13 2 16 4 9 9 13 1 10 0 9 2 13 9 13 2 10 9 7 9 9 13 2 7 3 15 15 1 9 13 13 2
4 9 13 0 9
7 11 13 2 16 13 10 9
13 16 15 9 13 7 13 2 3 15 11 11 13 2
13 1 9 9 2 15 15 13 9 7 13 1 9 2
15 1 9 0 9 1 9 11 11 2 11 2 15 3 13 2
18 0 11 3 14 3 3 9 13 2 7 10 9 1 9 13 1 0 2
27 1 0 11 15 13 9 2 9 1 9 15 13 1 0 9 9 11 7 1 9 0 9 13 1 0 9 2
9 7 1 9 15 13 9 0 9 2
13 2 3 4 15 13 2 16 4 1 15 9 13 2
16 3 16 4 3 15 13 1 11 11 2 9 13 13 11 11 2
15 0 13 1 15 0 2 13 15 15 2 16 4 13 9 2
10 3 4 1 15 13 2 15 1 15 2
9 13 10 9 2 16 4 15 13 2
9 13 13 9 2 16 4 13 0 2
11 3 14 15 1 15 13 2 16 13 9 2
10 2 13 0 13 9 1 9 10 9 2
9 15 4 3 13 2 3 3 3 2
27 3 9 13 7 3 15 3 13 2 16 9 2 9 2 13 0 9 2 16 0 9 9 2 13 15 2 2
12 7 16 4 15 13 0 9 2 3 13 0 2
10 13 3 13 2 16 4 13 9 9 2
18 2 16 15 13 3 2 3 13 13 2 16 4 1 9 13 1 9 2
6 13 15 7 0 9 2
24 3 2 1 15 15 13 0 9 2 3 15 13 14 9 2 7 3 15 3 13 1 0 9 2
15 9 15 0 15 13 1 9 2 7 15 4 15 3 13 2
12 7 14 15 1 15 1 9 15 1 9 13 2
18 3 14 2 0 9 13 1 10 9 2 7 13 9 1 0 0 9 2
12 2 13 15 2 16 15 3 9 3 13 9 2
8 14 2 3 1 15 1 9 2
23 13 13 9 1 9 2 7 1 9 2 15 15 3 13 1 9 2 4 13 4 9 13 2
15 10 9 13 2 16 9 13 10 9 7 9 13 9 9 2
12 2 3 15 4 13 2 16 13 1 0 9 2
14 7 16 4 13 0 9 2 13 4 1 9 1 9 2
20 3 16 4 1 0 13 1 9 1 11 2 13 4 2 16 13 13 0 9 2
8 2 3 0 13 1 9 9 2
11 11 13 0 9 2 15 4 13 1 9 2
11 15 13 0 9 2 15 4 1 9 13 2
9 9 15 13 9 2 16 4 13 2
22 13 4 0 9 1 9 7 13 15 2 15 13 2 7 1 9 4 13 12 1 10 2
14 9 15 13 1 9 2 13 4 2 16 13 10 9 2
31 3 13 13 7 3 13 10 9 2 13 10 9 2 15 9 2 15 15 3 3 13 1 9 2 13 7 3 15 3 13 2
6 2 15 10 11 11 2
13 0 9 2 3 15 9 13 1 9 1 0 9 2
25 3 15 13 2 16 13 1 10 9 15 0 2 7 15 13 0 9 1 0 9 2 13 1 9 2
9 9 15 13 1 9 1 9 9 2
22 13 15 1 9 2 7 13 15 15 2 16 15 1 15 13 2 16 1 12 13 9 2
12 13 0 2 16 9 13 7 1 15 15 13 2
11 2 13 13 9 0 9 2 16 9 13 2
18 13 15 1 15 13 2 7 3 15 13 13 14 1 15 7 10 9 2
12 7 4 13 12 9 1 0 9 13 1 9 2
30 1 11 9 13 9 2 3 13 0 9 2 15 15 13 13 1 0 9 2 3 13 3 10 9 2 15 10 9 13 2
9 2 13 15 13 0 9 1 0 2
11 9 13 0 9 2 9 13 3 0 9 2
18 14 3 4 15 13 2 16 1 9 4 15 13 3 2 3 4 13 2
12 13 2 16 4 15 15 15 13 16 9 9 2
8 15 13 3 9 1 10 9 2
14 13 3 3 9 2 13 0 0 9 2 7 13 9 2
6 9 13 0 7 0 2
10 13 1 9 7 13 9 13 0 9 2
8 2 15 15 13 9 1 9 2
10 16 15 13 13 14 7 14 1 15 2
17 13 15 3 0 9 2 13 15 9 2 7 3 4 13 9 13 2
12 9 13 0 9 2 7 1 9 13 9 0 2
5 2 11 2 0 11
6 11 1 11 9 11 11
4 11 11 2 11
52 3 12 3 0 9 10 0 0 9 1 9 11 2 12 1 11 2 1 11 2 12 2 12 2 7 11 2 12 2 12 2 9 9 1 11 4 1 9 9 10 9 13 2 2 13 9 1 0 9 11 11 2
19 15 2 16 0 2 13 1 9 3 1 9 2 3 1 9 13 11 11 2
23 12 1 10 9 2 15 13 9 0 9 1 11 7 13 7 0 9 2 13 9 11 11 2
4 13 3 13 2
32 0 9 13 1 15 2 16 9 1 10 9 3 13 0 9 2 7 11 13 2 16 3 1 15 13 13 9 9 1 9 9 2
7 1 11 4 9 13 3 2
11 1 0 9 3 3 13 9 1 0 9 2
31 13 2 16 13 9 1 9 3 0 2 16 15 1 9 15 13 13 1 0 9 7 1 9 1 0 9 2 13 11 11 2
10 12 12 14 13 1 9 3 0 9 2
13 0 9 1 0 9 13 7 1 11 0 16 0 2
9 13 15 0 2 3 1 1 9 2
12 11 3 13 14 11 7 3 3 13 1 9 2
8 11 15 13 1 15 3 3 2
15 15 7 15 13 1 15 2 16 11 13 16 9 9 0 2
13 12 0 9 1 9 9 7 1 0 9 13 9 2
28 15 15 13 14 1 0 9 2 3 13 1 9 1 11 7 3 1 9 1 11 3 3 13 1 9 1 11 2
11 9 12 9 1 9 1 9 13 14 0 2
8 0 9 13 11 1 9 9 2
20 16 1 11 7 11 4 1 9 13 3 2 3 14 13 7 13 15 1 9 2
16 3 2 13 15 13 2 7 13 14 1 15 2 13 0 9 2
6 3 4 13 3 0 2
9 3 1 9 4 1 11 13 9 2
5 3 15 15 13 2
9 3 4 9 1 11 13 16 9 2
8 13 0 9 7 15 4 13 2
9 11 11 13 1 11 11 0 9 2
8 1 15 3 13 1 9 9 2
15 1 0 9 3 13 0 9 2 7 16 15 15 3 13 2
10 3 13 1 0 9 1 9 3 15 2
24 11 3 13 3 13 2 15 15 1 9 13 2 7 15 0 3 1 9 9 13 9 7 9 2
23 11 11 13 1 9 3 3 1 15 2 16 4 15 10 9 1 11 11 13 13 1 0 2
20 13 9 2 3 3 7 1 9 2 15 15 13 14 1 9 2 13 11 11 2
5 3 15 15 13 2
12 9 15 7 3 13 2 14 16 15 9 13 2
4 0 11 13 9
6 0 11 2 11 2 2
24 1 9 2 12 9 1 9 2 13 9 1 0 9 9 9 1 0 11 2 9 12 9 2 2
24 3 15 15 13 2 13 15 0 9 11 11 2 15 13 1 0 0 0 1 9 3 0 9 2
24 10 9 15 15 13 2 15 13 1 9 2 16 13 1 9 7 13 2 16 15 13 13 9 2
25 3 13 0 2 16 1 9 13 13 3 9 3 2 16 4 15 13 13 1 0 9 2 13 11 2
3 11 1 11
5 11 2 11 2 2
16 1 11 11 7 11 11 13 9 0 9 0 9 0 0 9 2
9 13 15 15 12 0 9 11 11 2
35 9 9 1 11 12 3 1 11 0 9 13 2 7 3 15 1 11 1 9 9 11 13 0 9 0 11 11 2 3 1 0 9 13 9 2
18 11 13 3 9 1 11 11 2 15 1 0 9 13 0 9 1 11 2
24 1 9 1 11 15 13 1 11 13 3 1 12 9 2 7 3 13 0 2 13 1 15 11 2
9 0 9 11 13 11 3 1 11 2
7 13 15 2 3 13 11 2
2 9 13
5 11 2 11 2 2
38 9 9 0 0 9 0 11 13 1 0 0 0 9 2 9 11 11 2 0 9 1 12 9 2 10 9 9 9 11 13 7 13 16 0 9 14 0 2
29 0 9 15 3 1 0 9 1 0 9 3 13 9 9 2 11 11 2 1 10 9 13 3 0 9 0 11 11 2
18 0 13 0 11 11 2 16 12 1 9 11 13 13 10 9 7 13 2
1 3
21 9 0 9 13 1 9 9 1 11 0 9 2 15 13 0 9 1 9 10 9 2
11 9 0 9 4 10 0 9 13 1 9 2
14 0 9 9 13 11 2 11 2 11 2 11 7 11 2
12 15 13 0 9 1 9 0 1 9 7 9 2
2 9 13
2 11 2
34 9 12 2 9 0 9 1 9 11 11 1 11 11 9 11 13 1 1 15 2 16 0 11 11 13 0 9 12 2 0 12 12 9 2
8 0 13 11 2 0 11 11 2
34 9 9 1 0 9 13 9 9 2 15 13 13 1 9 1 0 9 2 13 9 7 9 1 9 2 7 7 15 9 1 9 13 2 2
10 1 9 13 11 1 9 9 1 11 2
20 1 3 0 0 9 10 9 3 13 2 1 10 9 13 3 0 9 1 9 2
12 1 9 9 11 3 14 13 9 7 3 13 2
36 1 0 9 13 3 11 2 11 7 13 1 0 9 9 1 11 13 3 16 12 9 1 11 2 7 13 15 3 0 9 1 9 12 12 9 2
10 13 15 3 12 0 9 1 12 9 2
19 1 0 9 0 9 13 1 11 2 11 0 11 9 0 11 12 2 12 2
18 0 9 7 13 9 2 14 1 9 10 0 9 9 2 9 9 2 2
6 9 4 13 9 11 2
5 9 11 11 2 11
4 0 9 13 9
7 9 11 11 15 13 1 11
2 11 11
17 0 9 1 9 0 13 1 9 12 9 12 9 0 11 11 11 2
11 10 9 15 13 7 0 0 9 1 9 2
33 3 0 9 15 13 1 9 1 0 9 0 9 1 11 1 9 0 9 2 13 9 2 12 2 7 13 0 1 9 2 12 2 2
9 2 3 4 15 13 1 0 9 2
38 1 11 11 2 9 7 9 1 12 9 2 15 13 1 9 12 0 9 11 1 9 2 13 1 11 9 7 9 15 1 15 13 1 9 1 9 9 2
7 2 1 15 13 10 9 2
10 13 10 0 9 2 14 9 1 9 2
6 3 13 3 1 9 2
8 9 1 15 3 3 3 13 2
9 2 3 4 15 13 13 1 11 2
12 16 13 3 1 11 3 9 7 13 3 9 2
17 1 15 13 0 0 9 2 9 3 13 7 9 13 0 7 0 2
8 2 3 3 13 1 11 13 2
24 1 15 4 3 13 2 3 15 15 3 13 2 13 15 3 2 16 4 13 13 3 1 11 2
22 2 10 0 9 13 3 0 15 2 16 4 13 1 11 7 13 1 0 9 2 2 2
18 13 4 10 0 9 9 7 1 9 15 3 13 13 10 9 16 3 2
24 16 3 13 2 13 15 9 2 7 16 4 13 13 15 1 0 9 2 13 15 9 1 15 2
16 2 15 13 9 1 11 11 2 16 13 0 9 2 7 3 2
27 1 9 2 3 15 13 7 13 1 9 2 4 13 1 2 0 9 2 3 1 9 0 9 7 0 9 2
14 3 13 0 9 2 15 13 13 3 7 13 1 9 2
12 0 9 9 0 2 0 2 0 2 0 11 13
9 11 2 11 2 11 2 11 2 2
11 0 0 9 1 9 13 9 12 2 9 2
48 9 0 2 0 2 0 2 0 11 3 1 11 3 1 0 9 13 2 1 9 7 11 13 13 7 3 1 0 9 0 9 11 13 1 15 2 16 0 2 11 13 9 3 1 9 0 9 2
11 1 0 9 15 0 11 3 13 1 11 2
25 3 12 9 1 9 15 13 2 16 0 13 0 0 9 2 9 15 7 13 12 0 9 0 11 2
21 11 13 3 1 15 1 0 9 7 3 3 13 2 3 1 9 1 11 1 11 2
18 11 13 13 1 11 7 3 2 16 13 1 12 2 9 1 0 11 2
24 1 11 13 0 9 2 3 3 0 0 9 1 0 9 1 11 2 13 1 0 9 11 2 11
17 11 2 0 11 12 2 12 2 12 2 12 2 2 9 2 12 2
12 9 0 9 2 11 2 11 2 11 2 12 2
2 11 11
22 1 9 1 10 9 1 0 9 11 11 2 9 0 9 1 9 2 13 2 10 11 2
4 13 15 3 2
19 0 2 9 9 2 0 9 2 15 1 10 0 9 13 3 12 0 9 2
15 0 9 1 11 2 0 9 0 9 2 9 9 0 9 2
7 0 9 7 9 0 9 2
4 9 0 9 2
14 0 9 0 9 0 9 7 1 0 9 9 0 9 2
17 11 13 9 2 16 0 9 4 13 0 9 3 1 9 0 9 2
22 11 11 2 11 2 12 2 12 2 15 13 1 11 1 11 2 1 0 9 16 11 2
9 1 0 15 10 12 9 13 0 2
22 0 9 2 0 9 2 9 13 0 9 2 7 16 0 9 1 0 9 13 3 0 2
36 9 9 0 9 7 0 9 9 1 0 7 1 9 0 0 9 2 13 1 0 9 3 16 9 0 9 11 0 0 11 2 9 0 9 2 2
11 1 10 3 0 9 13 0 9 0 9 2
23 13 1 0 9 0 9 2 11 13 3 1 0 9 15 9 2 7 13 15 16 3 0 2
18 1 9 15 10 9 13 15 2 16 15 0 9 13 0 7 0 9 2
16 9 0 9 13 3 15 2 16 15 12 1 9 13 13 3 2
30 10 9 13 9 2 9 2 15 15 13 1 9 2 7 7 3 13 13 1 9 9 2 15 13 7 9 2 7 9 2
26 10 9 15 1 9 13 15 2 16 13 0 9 0 9 2 7 9 15 14 3 13 1 9 0 9 2
19 9 13 3 16 9 7 1 0 9 9 2 15 15 10 9 13 1 9 2
19 0 9 2 9 2 13 7 10 9 3 1 9 2 7 1 9 0 9 2
15 4 13 9 1 9 7 9 7 13 0 9 0 1 9 2
40 13 10 9 3 1 9 0 0 9 0 0 0 9 2 16 15 13 9 2 7 1 9 9 0 9 2 9 0 9 2 9 0 9 9 2 7 9 0 9 2
13 10 9 0 9 13 3 0 9 7 13 0 9 2
14 3 7 3 15 15 13 9 7 0 0 9 3 13 2
22 1 9 10 0 9 15 9 13 1 0 9 2 1 15 13 3 7 9 2 7 9 2
24 0 0 9 4 13 2 7 0 9 1 10 9 13 13 9 1 9 0 9 7 3 0 9 2
14 10 0 9 9 7 9 15 3 13 1 9 0 9 2
19 1 15 13 9 1 15 15 2 16 15 13 0 9 2 7 16 15 13 2
8 0 9 13 7 9 0 9 2
25 15 2 16 11 13 0 9 0 9 7 13 0 9 2 13 3 0 9 7 11 16 11 7 11 2
19 13 2 16 9 9 15 3 13 12 9 2 9 0 9 7 9 9 9 2
24 0 4 13 0 9 0 9 2 1 15 0 9 13 9 9 7 0 9 15 13 9 0 9 2
30 1 0 13 0 9 0 7 0 9 2 0 9 4 13 3 9 7 9 15 13 3 10 0 9 16 0 9 0 9 2
33 15 13 11 9 2 13 9 2 10 9 15 13 1 10 0 0 9 11 2 11 7 11 2 15 13 0 9 1 0 2 0 9 2
24 3 2 16 15 0 9 13 1 0 9 0 9 2 13 9 9 7 9 2 9 3 10 9 2
20 9 15 3 13 15 3 15 3 9 9 7 9 2 14 2 14 14 0 9 2
8 15 13 7 1 11 0 9 2
30 0 9 2 15 13 9 0 0 9 15 2 16 13 0 9 2 13 9 3 13 7 1 15 7 10 0 7 0 9 2
28 3 13 0 0 9 7 0 9 7 3 7 9 0 15 13 0 9 7 1 0 9 2 7 7 1 9 9 2
19 15 13 9 1 0 9 7 13 15 9 1 9 0 9 0 1 0 9 2
21 11 15 1 10 0 9 13 2 10 9 2 9 2 7 9 2 4 13 9 9 2
16 1 9 2 9 7 9 9 10 9 13 3 2 13 15 9 2
17 1 10 0 9 0 9 13 11 2 9 7 11 2 9 0 9 2
8 3 7 13 10 9 1 0 2
8 9 13 9 2 15 11 13 2
10 13 10 9 9 2 10 0 0 9 2
25 13 2 16 16 13 1 0 9 2 13 11 9 2 0 9 15 3 13 1 3 3 0 9 0 2
7 9 4 13 10 0 9 2
20 15 13 10 0 9 2 0 3 1 9 2 15 4 3 13 1 9 0 9 2
7 10 15 1 15 13 9 2
25 1 0 2 13 2 3 9 9 13 9 9 7 13 9 9 2 15 9 13 2 7 15 0 9 2
11 9 0 9 7 9 4 3 13 0 9 2
10 0 9 13 0 7 13 1 9 0 2
9 13 1 15 2 16 9 13 9 2
20 13 1 12 12 9 15 2 16 13 9 2 9 2 9 7 9 9 1 9 2
9 13 15 2 16 13 0 0 9 2
22 11 15 13 2 16 0 9 13 0 0 9 2 15 13 3 13 1 10 9 7 9 2
14 13 2 16 0 9 13 0 2 7 0 2 0 9 2
15 13 14 15 2 16 15 13 9 7 13 0 7 0 9 2
22 1 9 2 13 11 2 15 13 7 9 2 7 9 15 13 2 15 10 9 3 13 2
22 7 16 15 3 13 2 13 3 14 0 9 2 16 1 0 9 15 10 9 3 13 2
28 3 16 9 1 0 9 9 0 9 2 9 7 9 4 3 13 1 0 0 9 2 15 4 13 9 0 9 2
16 13 9 1 10 9 1 9 2 15 13 9 9 3 1 9 2
12 13 15 2 16 13 9 1 9 2 15 13 2
17 10 9 13 1 9 12 2 3 0 9 9 13 1 15 12 9 2
33 11 13 1 0 0 9 7 16 4 3 13 2 14 4 13 2 16 15 13 3 3 0 9 2 16 4 13 0 13 15 1 9 2
32 9 9 4 13 7 1 15 2 16 15 13 0 2 7 3 2 1 1 9 1 0 0 9 1 9 0 2 9 9 12 9 2
21 9 4 15 13 1 0 2 0 7 3 0 9 2 7 3 4 13 1 9 9 2
7 11 15 13 7 13 9 2
32 1 0 9 9 13 15 9 2 3 4 13 4 0 9 13 7 13 2 16 4 15 13 0 9 7 0 9 0 9 7 9 2
25 16 15 9 13 1 0 9 2 13 3 9 0 9 2 15 13 10 9 1 15 1 0 0 9 2
24 0 9 2 15 1 9 13 2 13 2 9 15 13 1 9 9 2 3 4 0 9 13 13 2
23 7 3 2 16 15 13 2 16 13 9 1 9 2 16 13 4 2 1 0 9 0 9 2
24 1 10 0 11 2 0 9 2 13 0 9 0 0 9 2 15 13 10 9 15 0 16 0 2
43 13 7 9 9 13 9 2 16 0 9 15 13 9 0 9 7 16 13 12 9 10 9 2 9 1 0 9 12 9 2 9 0 9 9 7 9 0 1 12 1 12 9 2
30 15 2 15 11 13 2 7 13 1 15 9 16 11 2 11 2 11 2 15 13 1 15 2 16 15 13 3 0 9 2
39 1 11 2 3 10 0 9 13 1 0 0 9 14 1 10 9 2 13 0 9 2 13 4 13 0 9 1 9 2 0 9 1 9 7 0 9 1 9 2
9 1 1 0 9 0 9 3 13 2
40 11 13 2 16 13 0 9 2 10 9 7 9 13 9 2 0 9 0 0 9 2 1 15 9 13 9 15 9 1 0 9 2 7 9 1 3 15 9 9 2
12 1 0 13 1 11 0 9 9 2 1 9 2
32 7 16 13 1 0 9 0 9 7 0 9 13 7 13 2 13 15 13 1 3 0 0 9 2 15 13 11 2 11 7 11 2
7 11 11 13 7 1 0 9
2 11 2
23 9 11 11 13 0 9 1 9 2 13 15 12 0 9 2 13 12 9 7 13 14 0 2
7 3 9 11 3 13 9 2
25 12 9 3 2 16 13 1 12 9 9 0 9 11 11 1 11 2 13 9 1 11 11 1 11 2
10 10 9 13 0 9 1 12 9 9 2
5 11 3 3 13 11
2 11 2
28 0 0 9 11 11 2 15 1 12 9 13 12 9 2 15 3 13 10 0 9 11 0 14 1 9 0 9 2
22 10 0 9 3 13 14 1 12 9 2 7 9 9 3 13 13 10 9 1 0 9 2
19 15 11 13 2 16 13 1 11 3 0 7 13 1 15 13 3 3 3 2
14 11 0 13 13 1 11 11 7 3 2 13 9 11 2
3 1 0 9
20 11 11 2 12 2 2 12 1 0 0 9 15 9 2 13 1 11 1 9 2
4 11 3 1 0
10 1 9 15 13 7 11 2 11 13 9
6 11 2 11 2 11 2
15 0 0 9 11 11 15 13 9 0 9 0 9 1 11 2
19 1 12 9 9 13 3 1 0 7 13 3 1 9 1 11 12 2 12 2
25 11 2 10 9 13 3 11 11 2 13 1 12 9 0 9 9 12 9 2 3 16 0 12 9 2
13 16 9 0 9 9 15 7 3 13 9 1 9 2
10 1 0 9 15 13 7 0 0 9 2
32 12 9 13 11 11 1 9 11 2 11 11 13 10 9 9 1 9 11 1 11 7 10 0 9 1 9 0 9 13 11 11 2
12 10 9 13 1 9 11 1 11 12 2 12 2
32 3 1 0 9 15 1 9 9 13 0 9 2 11 11 9 1 0 9 13 1 9 11 1 3 0 11 2 12 2 12 2 2
14 3 3 1 12 2 9 11 11 13 1 0 9 11 2
21 11 13 1 11 1 11 12 12 2 12 2 11 13 0 9 2 11 14 0 9 2
26 9 9 11 11 15 3 1 9 13 1 9 1 0 9 2 12 9 13 1 11 2 12 2 12 2 2
21 9 13 11 11 2 7 3 0 11 15 13 0 9 2 12 2 12 2 1 11 2
9 3 13 1 0 9 0 11 11 2
48 9 0 9 11 11 13 1 11 11 1 10 9 12 2 12 2 16 12 9 2 0 3 1 12 9 9 2 13 11 11 2 15 13 11 1 9 13 2 7 1 12 9 1 15 13 7 9 2
18 1 9 13 7 11 7 11 1 9 2 3 11 11 11 0 9 13 2
21 0 11 2 3 2 7 11 2 11 2 1 9 1 9 1 9 12 2 9 9 2
14 1 12 9 15 13 11 2 16 13 3 12 2 12 2
2 9 11
5 1 9 13 0 9
7 11 2 11 2 11 2 2
20 1 0 9 13 1 11 1 11 13 3 1 9 9 0 9 11 1 12 9 2
18 9 9 13 1 9 1 0 7 13 3 0 9 1 9 12 1 11 2
24 11 4 3 13 13 2 7 1 10 9 13 15 0 1 9 2 13 15 1 9 7 13 9 2
12 13 13 3 0 2 13 9 0 9 11 11 2
18 11 15 13 7 1 0 9 2 3 3 15 9 13 9 9 1 9 2
11 15 4 1 9 13 2 13 11 9 11 2
12 9 13 1 12 9 7 13 15 0 9 11 2
32 0 9 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 2 11 2 11 2 11 2 11 11 2 11 2 11 2
4 0 9 1 9
9 11 15 9 1 11 0 13 1 9
4 11 11 2 11
39 9 9 7 10 9 1 9 13 9 11 11 1 15 2 16 4 3 13 0 0 9 11 2 11 2 11 2 11 2 11 9 1 11 7 13 3 0 9 2
35 1 9 1 12 9 3 15 1 0 9 13 9 9 0 9 7 14 1 12 9 12 15 13 11 2 11 7 11 2 9 2 9 2 2 2
21 3 4 13 1 9 7 15 0 9 13 2 16 4 15 13 0 9 2 13 11 2
12 0 9 1 0 9 13 3 1 9 11 11 2
14 3 16 1 9 15 1 9 1 11 13 1 0 9 2
11 9 9 4 13 2 16 4 15 13 13 2
25 3 4 3 9 1 11 3 13 2 16 4 15 13 2 7 9 13 2 16 4 13 9 1 9 2
12 2 1 9 15 7 1 9 13 9 2 2 2
9 1 9 1 11 4 13 12 9 2
33 3 13 1 9 2 16 4 15 13 2 1 12 9 1 11 4 13 9 2 3 9 13 3 1 9 2 7 3 9 13 1 9 2
26 13 2 16 15 15 13 13 12 9 1 0 9 2 7 3 15 13 2 16 15 1 9 9 13 3 2
26 9 15 15 13 10 0 9 2 13 4 3 1 12 9 1 12 2 7 3 4 13 1 9 0 9 2
10 2 3 15 1 9 0 9 13 11 2
6 3 15 13 16 9 2
7 11 13 3 1 15 3 2
18 1 9 11 4 3 13 7 12 13 0 9 2 16 0 9 15 13 2
10 3 0 15 13 1 9 7 13 15 2
4 9 9 3 13
4 9 1 0 9
10 1 0 9 9 1 0 9 3 13 2
9 0 9 1 11 13 1 9 9 2
10 7 1 0 9 13 9 0 9 0 2
19 9 13 1 9 0 9 11 7 3 1 0 9 1 9 1 11 1 9 2
8 9 13 9 9 1 0 9 2
19 1 9 9 13 1 12 9 2 15 13 0 9 1 9 1 9 0 9 2
13 1 9 9 0 9 3 1 9 13 1 0 9 2
16 9 13 0 9 9 1 0 9 10 9 1 9 0 9 11 2
11 15 13 1 9 9 0 9 1 12 9 2
10 9 13 1 9 1 9 9 12 9 2
14 1 9 1 9 1 9 1 9 1 11 9 3 13 2
24 13 1 15 9 1 15 2 16 4 13 3 0 9 9 0 9 1 0 9 13 1 0 9 2
12 9 9 1 0 9 1 0 9 3 3 13 2
10 9 13 1 9 3 0 1 0 9 2
14 0 0 9 0 9 13 14 9 1 0 9 1 11 2
9 1 9 7 1 9 9 9 13 2
25 0 9 1 0 11 3 1 11 13 9 1 0 9 0 9 14 1 0 9 12 9 1 0 9 2
14 15 7 13 3 0 1 15 2 16 4 13 4 13 2
23 1 9 4 9 9 13 9 9 2 15 0 9 13 1 9 14 1 12 9 1 0 9 2
20 9 9 1 0 9 3 3 13 1 12 1 12 9 1 9 2 12 9 2 2
7 0 0 9 2 11 7 11
2 11 11
28 16 9 0 9 2 3 16 0 2 13 1 9 1 9 12 3 1 9 2 9 1 9 1 11 13 3 3 2
16 9 13 3 1 9 0 11 2 16 3 13 11 12 2 12 2
9 1 9 15 13 3 0 0 9 2
25 1 0 9 9 7 13 9 2 3 3 3 9 1 0 9 3 1 9 9 7 9 1 9 13 2
27 9 1 10 9 13 11 2 0 11 2 7 11 2 15 15 13 3 1 12 9 2 3 1 12 0 9 2
2 9 12
12 11 2 11 2 11 2 11 2 11 2 11 2
21 1 11 7 11 13 15 0 9 3 2 11 3 1 0 9 13 1 9 1 9 2
25 7 7 12 0 9 9 10 3 15 13 2 7 16 13 7 1 9 9 2 7 9 1 9 9 2
27 11 13 3 1 9 15 2 11 14 11 2 7 15 3 3 14 11 2 1 15 13 1 9 1 9 12 2
11 9 1 11 15 3 13 1 9 1 11 2
12 1 11 15 9 9 0 9 13 1 9 12 2
6 11 7 11 13 9 2
19 11 13 11 1 9 1 11 7 9 15 3 13 2 16 15 13 7 9 2
26 11 13 1 11 3 1 0 9 2 9 12 2 9 12 2 9 12 2 2 1 11 14 1 9 12 2
15 15 10 12 9 13 11 2 7 13 1 15 3 7 9 2
15 11 3 13 11 3 1 9 12 7 1 0 9 9 12 2
13 0 9 3 13 0 9 1 9 2 11 7 11 2
15 1 9 1 11 12 13 3 1 0 13 14 0 0 9 2
5 3 15 13 11 2
15 11 0 13 1 9 1 9 12 2 3 1 15 13 11 2
10 11 13 1 9 1 9 12 7 11 2
20 7 3 1 12 0 9 2 9 12 7 9 12 2 13 11 7 3 13 11 2
9 1 11 7 11 11 3 3 13 2
23 1 12 9 1 10 9 13 1 0 9 2 3 15 13 14 11 1 11 2 9 12 2 2
7 1 10 9 13 0 9 2
21 3 15 3 13 11 1 11 2 15 15 3 1 9 9 12 2 9 9 2 13 2
23 0 9 13 3 9 1 11 1 9 1 9 12 2 7 1 0 9 15 13 7 1 9 2
18 1 11 4 13 3 14 1 0 9 2 9 12 2 9 12 7 12 2
11 11 7 11 3 13 1 9 1 9 12 2
14 13 3 12 9 2 7 11 1 0 9 13 12 9 2
4 11 13 9 2
10 11 2 11 2 11 2 11 2 11 2
27 1 9 12 15 12 0 9 13 3 3 1 9 2 1 0 9 13 7 1 9 1 9 1 12 0 9 2
14 1 9 1 9 12 1 15 13 1 9 3 7 11 2
20 0 2 11 13 1 0 9 1 9 1 11 2 1 11 3 3 1 12 9 2
12 3 11 13 10 9 1 11 14 1 0 9 2
15 9 11 1 11 13 1 9 12 2 3 11 13 1 9 2
8 11 7 11 13 1 9 3 2
17 11 0 13 1 0 9 1 9 1 11 7 4 15 13 1 9 2
12 13 7 13 7 1 11 7 13 9 1 11 2
18 11 13 3 9 13 2 7 7 11 2 7 11 13 3 1 10 9 2
24 11 13 1 11 1 9 1 9 1 11 7 3 16 9 0 9 3 1 9 1 9 7 9 2
27 11 3 13 1 0 9 9 7 9 14 3 2 7 3 1 9 1 11 7 11 2 7 3 13 9 9 2
20 11 1 11 13 14 1 11 7 1 9 1 11 2 3 11 2 3 11 2 2
20 11 13 10 12 9 3 2 7 3 13 9 2 3 16 0 9 7 0 11 2
14 9 11 2 3 2 13 1 0 11 1 0 9 1 11
2 9 11
4 0 9 16 9
6 11 13 13 1 11 2
6 9 10 9 13 12 9
7 11 2 11 2 11 2 2
16 3 14 9 13 0 0 9 1 0 9 1 9 1 9 12 2
9 3 1 12 13 1 11 1 11 2
38 0 9 15 1 9 1 0 9 13 11 1 9 3 2 0 11 13 12 2 12 2 12 2 12 2 9 11 2 11 2 11 2 1 9 2 7 11 2
22 13 1 0 9 2 9 11 13 1 9 13 9 7 13 3 2 16 15 14 13 11 2
10 13 15 1 9 2 13 9 11 11 2
21 1 9 15 13 11 1 9 2 1 15 15 13 2 15 1 11 3 13 0 11 2
6 0 9 13 0 9 2
19 13 1 12 9 0 16 1 9 1 11 2 13 11 10 9 1 0 9 2
19 3 15 9 13 1 9 11 1 11 1 11 2 3 4 14 1 9 13 2
24 1 9 1 9 13 9 1 11 0 9 2 15 13 1 9 9 12 2 7 12 2 0 9 2
15 3 15 3 13 2 1 3 0 11 2 1 11 1 11 2
23 9 3 13 1 12 2 2 2 9 7 1 9 9 12 2 9 9 15 13 7 0 9 2
17 10 9 1 9 4 1 15 3 13 2 13 9 9 11 9 11 2
9 9 11 13 1 10 9 0 9 2
13 13 15 3 13 13 0 9 7 13 1 0 9 2
16 13 9 1 0 2 16 4 15 1 9 13 9 2 13 11 2
9 3 13 1 9 9 0 9 9 2
24 13 15 9 11 2 11 2 3 15 11 3 13 9 9 7 13 15 14 1 9 12 2 12 2
19 3 13 0 9 10 9 1 11 2 9 9 15 15 3 13 2 13 11 2
14 1 11 13 3 3 11 2 7 10 9 13 0 9 2
27 9 15 3 13 2 16 15 13 1 11 2 3 1 9 3 13 2 7 1 9 11 15 13 14 1 9 2
10 7 11 13 10 9 2 3 15 13 2
15 3 11 13 1 0 9 1 9 1 9 1 0 9 11 2
7 11 13 13 13 3 12 9
5 11 2 11 2 2
23 0 12 1 12 0 9 2 15 3 13 1 0 9 2 13 1 0 9 0 9 13 13 2
27 9 9 7 0 9 0 9 11 11 15 13 1 9 9 11 11 11 2 16 4 3 13 10 9 1 11 2
14 10 0 11 13 3 0 1 9 2 15 13 10 9 2
20 1 0 9 4 1 12 9 13 0 9 12 0 0 9 1 9 1 12 9 2
27 9 11 13 2 16 1 11 15 13 0 9 14 1 12 9 2 10 9 13 3 13 2 7 7 0 12 2
27 0 9 13 9 0 9 11 2 16 4 13 0 9 0 9 7 13 13 0 9 2 15 4 13 10 9 2
7 10 9 4 13 10 9 2
22 10 0 0 9 2 15 13 1 10 9 2 3 4 3 13 1 0 9 1 0 9 2
25 4 13 1 0 9 1 15 2 16 4 1 9 1 9 10 9 13 1 9 2 1 15 15 13 2
16 1 10 9 13 13 1 0 9 15 0 9 2 13 11 11 2
4 0 9 1 9
7 11 2 9 11 11 2 2
25 0 9 2 15 4 1 0 9 13 1 10 0 9 2 15 3 13 7 1 9 11 1 0 9 2
5 13 9 0 9 2
17 9 3 14 13 2 16 1 15 3 0 9 13 16 0 3 3 2
22 9 0 0 9 2 15 9 13 2 15 7 13 2 16 9 13 9 9 10 9 3 2
26 9 2 15 3 9 13 2 13 2 16 15 13 2 16 4 10 9 3 1 9 13 1 9 10 0 2
20 16 13 12 1 9 9 2 4 7 3 13 1 9 1 9 0 9 7 9 2
5 9 1 9 11 11
10 9 1 9 2 9 7 9 1 0 9
2 11 2
16 3 9 15 1 0 9 1 11 13 0 9 9 0 11 11 2
20 9 0 1 9 2 9 7 9 15 14 1 0 0 9 1 9 13 1 9 2
12 0 9 15 1 9 9 13 12 7 12 9 2
14 9 13 9 9 1 0 9 7 0 9 14 1 11 2
11 1 9 9 0 15 13 12 7 12 9 2
40 9 15 3 13 9 1 0 9 2 3 1 9 0 11 13 9 2 1 15 1 9 11 2 11 13 0 0 9 9 2 0 11 11 0 1 11 9 9 9 2
46 1 9 15 3 2 13 2 1 9 0 9 1 9 13 3 7 3 10 9 2 15 3 3 13 1 9 2 13 0 9 7 13 15 1 10 2 16 4 12 9 13 9 1 10 9 2
23 13 15 1 9 3 0 0 9 2 9 1 9 2 0 9 11 2 13 9 1 10 9 2
12 9 1 9 9 13 1 9 0 9 1 9 2
25 3 9 15 1 9 13 9 1 9 2 3 1 9 9 0 13 9 0 9 0 11 9 11 2 11
5 9 11 11 2 11
3 9 0 9
5 9 11 11 2 11
4 11 13 1 11
5 11 2 11 2 2
38 9 0 9 7 0 9 0 0 11 2 11 2 11 11 2 11 13 2 16 9 13 1 11 9 1 9 0 9 7 9 1 0 9 12 9 2 9 2
33 1 0 9 13 9 2 16 9 13 1 11 3 0 16 0 9 12 0 9 2 16 1 9 1 0 9 15 9 13 0 12 9 2
27 1 9 0 9 4 13 12 12 9 9 7 0 9 1 9 3 16 12 9 2 9 1 9 1 9 11 2
15 1 9 0 12 9 11 13 9 0 0 9 1 12 9 2
13 9 9 4 13 9 9 0 9 1 9 1 11 2
3 9 1 11
18 9 1 0 9 1 9 11 11 2 0 0 9 1 15 13 0 9 2
16 13 15 1 9 1 11 13 9 9 1 9 7 9 1 11 2
24 10 9 13 3 1 9 0 9 9 7 3 13 10 9 2 13 10 9 2 9 10 0 9 2
19 3 15 13 13 1 9 9 0 9 9 9 2 13 12 2 9 9 11 2
21 3 15 13 13 16 0 9 9 0 9 11 2 3 15 4 3 13 1 10 9 2
13 3 4 13 1 9 12 2 9 9 0 0 9 2
34 7 15 15 3 3 13 0 9 9 10 9 2 9 2 9 2 3 15 3 13 2 7 3 0 9 2 1 15 4 15 15 13 13 2
23 13 9 2 16 10 9 15 3 7 3 13 1 10 9 7 15 15 3 1 10 9 13 2
13 13 4 1 10 9 7 0 9 1 10 9 9 2
22 1 10 9 4 13 13 1 9 7 13 0 0 9 2 9 2 9 2 9 7 3 2
31 13 4 14 13 2 16 10 9 2 3 0 2 3 0 2 3 15 0 0 9 10 9 2 13 16 9 0 1 0 9 2
35 13 4 15 15 3 13 1 9 1 0 2 13 1 15 0 9 7 3 13 10 9 1 0 10 9 9 7 1 10 9 1 10 0 9 2
16 13 0 2 16 9 9 1 10 0 9 13 3 3 0 9 2
47 13 3 3 11 2 11 16 0 9 1 0 0 9 2 15 3 13 1 9 11 2 7 13 0 9 9 2 0 9 2 15 1 9 13 1 0 9 13 2 13 3 14 0 9 0 9 2
10 13 4 1 15 3 7 1 11 11 2
23 0 9 15 13 2 16 11 7 11 16 12 3 0 2 3 0 9 4 13 13 0 9 2
26 15 15 3 13 2 16 4 3 13 13 3 11 2 0 9 2 3 0 2 7 11 3 16 9 0 2
5 15 13 12 9 2
6 7 13 7 0 9 2
5 0 9 9 9 2
32 7 3 0 9 2 9 9 9 2 9 2 15 13 2 9 7 9 2 15 13 0 3 7 3 13 9 2 13 0 9 9 2
31 15 4 3 1 9 11 13 7 1 9 0 9 9 10 0 9 11 2 15 4 3 13 1 10 9 1 9 9 9 13 2
11 0 9 13 2 16 11 13 13 3 15 2
11 9 0 9 13 0 13 7 1 0 9 2
48 15 15 13 0 7 13 0 2 16 15 15 3 13 13 2 3 13 13 9 2 14 9 9 2 7 3 9 9 11 2 13 15 7 9 9 2 3 15 13 3 1 9 9 2 1 9 0 2
19 13 2 14 0 9 13 9 1 0 0 0 9 2 3 15 13 7 9 2
22 13 2 14 9 2 13 9 7 13 15 15 3 2 3 0 7 13 9 10 0 11 2
5 9 1 11 1 11
2 11 2
18 10 12 9 13 1 9 0 9 0 9 9 1 0 9 11 0 11 2
19 13 15 3 11 11 2 9 9 11 11 1 11 2 15 9 1 9 13 2
17 0 9 11 2 15 13 9 11 11 2 13 0 9 9 1 11 2
7 10 9 15 9 3 13 2
18 7 1 10 9 2 16 9 0 9 13 1 9 1 0 9 3 0 2
12 1 11 2 11 13 11 9 1 11 3 9 2
20 9 11 2 15 13 9 0 9 9 11 2 13 3 0 9 9 1 12 9 2
14 1 9 12 4 15 13 4 3 1 12 7 12 9 2
3 0 9 9
5 11 2 11 2 2
16 1 0 9 15 3 3 11 13 3 16 1 0 9 0 9 2
23 1 9 9 9 7 9 11 11 13 1 0 0 9 0 9 12 9 9 7 9 12 9 2
17 0 0 9 11 13 11 2 12 5 0 9 7 12 5 9 2 2
22 0 1 9 13 11 2 12 7 12 5 2 7 11 2 12 2 3 2 12 5 2 2
39 9 0 9 13 0 16 3 2 15 13 2 16 12 5 15 1 15 13 9 1 9 2 9 2 9 7 9 3 1 9 9 7 9 2 3 12 5 2 2
25 9 0 7 0 9 15 1 0 9 13 12 5 1 0 12 5 7 0 9 12 5 1 12 5 2
5 13 15 9 9 9
25 1 9 0 0 9 0 2 0 2 7 0 2 11 13 9 0 9 9 1 9 11 0 16 3 2
15 3 4 15 7 10 9 3 1 0 9 0 9 13 13 2
19 3 3 15 13 0 9 1 9 11 7 11 2 15 4 13 1 9 9 2
27 10 9 9 3 3 13 0 9 9 1 11 7 1 0 9 11 2 1 0 12 9 2 9 3 12 9 2
17 9 13 2 16 11 15 4 13 0 9 13 14 12 9 2 9 2
27 9 0 9 13 13 7 0 9 2 16 1 1 9 0 9 3 4 9 1 9 0 9 13 1 12 5 2
27 0 9 0 9 1 9 12 2 12 13 9 12 9 2 9 2 16 0 9 13 3 1 12 9 2 9 2
17 1 9 11 2 3 4 3 13 3 0 9 2 13 3 9 0 2
13 9 0 9 13 3 0 14 1 12 7 12 5 2
5 1 9 9 0 9
14 0 9 9 9 13 12 12 9 7 12 9 1 12 9
2 11 11
27 9 9 7 9 1 9 2 9 7 9 1 0 9 9 9 13 1 0 0 9 1 0 0 9 1 9 2
13 9 2 9 7 9 10 9 3 13 1 9 9 2
13 1 15 15 7 13 7 0 9 9 7 0 9 2
29 1 9 13 3 13 15 2 16 9 9 13 7 0 2 7 7 0 9 1 0 9 2 9 7 1 0 0 9 2
20 13 15 1 9 1 9 15 0 9 2 10 0 9 7 9 13 7 3 0 2
13 16 1 9 15 9 13 2 13 1 15 10 9 2
11 13 1 15 7 9 2 7 13 0 9 2
9 10 9 13 3 1 12 5 0 2
33 13 15 3 0 9 2 7 15 13 1 0 9 9 11 1 0 9 2 15 15 9 7 13 0 9 2 13 9 9 11 11 11 2
18 1 15 13 1 9 9 9 9 3 1 0 9 2 3 13 15 3 2
12 9 1 9 13 1 9 3 16 1 0 9 2
22 3 9 0 9 11 13 13 13 0 9 2 15 13 0 9 2 9 1 0 9 3 2
11 13 15 3 0 9 2 7 3 15 13 2
14 1 9 13 15 3 0 9 2 10 9 13 1 0 2
23 3 9 1 15 15 13 3 0 9 1 9 7 1 0 9 13 9 10 9 1 9 9 2
28 1 9 1 9 13 10 9 3 0 2 16 3 0 9 13 1 9 0 1 10 9 1 9 2 13 11 11 2
26 1 9 11 11 13 11 11 11 2 16 1 10 9 9 2 0 0 9 3 2 13 9 3 0 9 2
13 1 10 9 15 13 0 2 7 9 13 10 9 2
17 13 2 16 9 2 15 1 10 9 13 2 15 15 13 2 13 2
12 9 9 1 9 9 7 13 1 10 0 9 2
13 9 1 11 11 1 11 15 1 9 13 3 3 2
10 1 15 4 15 7 13 13 10 9 2
22 1 1 15 2 16 3 15 9 13 15 9 0 9 2 3 3 1 15 13 3 0 2
13 13 4 9 2 9 2 7 13 13 1 0 0 2
15 1 0 9 1 9 13 9 0 7 15 15 1 15 13 2
17 13 4 15 3 13 9 1 9 7 9 2 15 13 0 9 9 2
18 1 0 9 1 15 4 2 4 7 4 9 3 13 2 13 11 11 2
9 3 13 1 9 7 9 11 11 2
29 1 9 1 12 1 0 9 2 10 9 13 3 1 12 9 9 2 13 2 16 10 9 1 10 9 13 1 9 2
7 0 9 7 13 12 9 2
12 7 3 10 9 13 12 1 9 9 9 9 2
1 3
13 0 9 3 13 1 0 9 0 9 12 9 9 2
10 10 9 13 0 9 2 7 0 9 2
21 3 0 0 9 9 13 9 1 9 9 9 10 9 2 15 13 12 9 2 9 2
17 9 13 9 1 9 9 12 9 2 9 15 7 13 1 12 9 2
27 0 9 11 7 11 13 1 9 12 9 2 15 4 13 1 0 2 0 9 2 15 15 13 13 9 9 2
28 4 13 9 3 0 9 1 0 9 2 9 0 9 2 9 1 9 9 7 9 2 1 9 0 7 0 9 2
20 9 4 13 1 0 9 1 0 9 2 1 9 1 0 9 2 1 9 9 2
4 9 1 0 9
12 12 1 9 0 15 0 0 9 13 9 9 2
12 0 0 9 13 9 9 0 9 7 9 9 2
31 1 9 1 9 13 3 9 2 9 2 9 7 0 9 9 13 2 16 10 9 1 0 9 13 0 2 9 3 0 9 2
19 1 9 11 11 1 9 0 9 11 13 1 9 3 1 0 9 1 9 2
10 10 0 9 13 1 0 0 9 0 2
13 1 11 13 3 9 13 3 9 0 9 1 9 2
23 13 13 7 1 15 2 16 15 10 9 1 9 13 1 12 2 12 2 12 7 3 9 2
22 13 2 14 15 9 1 9 0 9 1 9 2 13 10 9 13 3 7 1 0 9 2
23 1 9 1 9 0 9 13 3 1 0 9 9 9 13 10 9 2 7 15 1 0 9 2
15 13 15 3 2 16 0 9 4 13 0 9 16 0 9 2
27 13 3 3 1 9 9 0 9 13 3 1 9 2 16 9 9 2 15 13 9 0 9 2 13 1 9 2
3 2 11 2
5 9 13 3 0 9
2 9 11
3 11 13 9
39 9 9 1 11 7 9 1 9 11 4 13 9 9 0 0 9 7 9 13 9 9 1 9 2 1 15 4 1 0 9 11 7 1 11 13 0 0 9 2
8 13 15 7 13 1 9 9 2
16 12 9 13 7 9 7 9 7 0 3 9 9 9 1 9 2
35 13 3 0 9 1 9 9 7 0 9 1 9 0 11 2 7 10 9 1 9 13 3 3 0 2 3 15 15 13 11 7 0 0 9 2
10 0 9 13 2 7 13 15 15 13 2
15 9 2 3 15 9 9 1 0 9 3 13 2 13 10 2
23 1 9 3 13 9 1 15 2 16 13 11 14 14 13 1 15 0 9 9 7 0 9 2
43 0 9 1 11 7 1 0 9 11 14 13 3 1 9 9 2 15 13 2 16 9 1 11 7 11 1 9 9 13 3 0 7 16 1 9 11 15 13 0 9 0 9 2
28 9 9 7 9 1 9 0 11 13 3 1 3 0 9 2 16 10 9 7 9 0 9 15 13 3 0 9 2
16 1 9 1 0 9 13 3 0 9 0 7 0 9 15 9 2
47 13 3 9 2 16 11 0 1 9 12 1 11 15 3 13 13 0 9 2 7 10 9 3 13 3 0 9 1 0 0 9 7 3 1 9 7 1 0 9 13 0 13 15 3 14 13 2
26 1 9 1 0 9 13 3 0 9 0 7 0 9 2 15 13 9 2 15 0 0 9 3 3 13 2
29 11 13 0 9 2 7 16 13 0 2 13 9 0 0 9 2 15 13 0 9 11 1 10 9 11 1 9 12 2
29 10 9 7 4 1 9 13 16 3 0 1 0 9 2 7 15 13 3 12 5 9 1 0 9 7 13 9 9 2
15 3 3 13 0 2 10 9 9 4 1 0 9 13 9 2
45 11 7 0 9 3 13 9 13 0 9 2 7 1 0 9 13 3 3 9 2 15 13 2 16 4 9 13 10 9 2 3 2 9 2 7 1 9 15 15 3 3 13 7 13 2
18 9 3 0 0 9 7 9 13 7 9 0 0 2 0 7 0 9 2
28 1 0 9 15 0 9 13 15 2 16 0 9 15 0 9 4 15 13 3 13 1 9 9 2 9 7 9 2
3 2 11 2
4 11 12 13 9
5 11 2 11 2 2
30 0 9 11 2 0 9 0 9 1 9 2 13 9 1 0 9 0 0 9 1 0 12 9 2 15 13 1 9 12 2
34 13 1 15 2 16 1 0 9 13 1 9 1 9 0 0 9 7 0 12 9 13 3 0 9 1 9 0 9 1 9 7 1 9 2
10 0 0 9 13 0 9 0 11 12 2
20 1 12 9 10 9 2 15 13 3 1 9 2 13 12 12 15 9 0 9 2
27 1 9 4 9 0 0 9 1 9 12 7 12 13 9 12 5 3 2 16 15 10 9 9 0 9 13 2
33 9 0 0 9 13 0 9 1 0 9 2 7 11 7 13 2 16 1 0 12 9 15 13 3 12 2 7 15 3 1 0 9 2
17 1 0 9 4 3 0 11 13 3 1 0 9 7 9 0 9 2
17 13 1 15 7 0 9 11 2 15 4 3 13 10 0 0 9 2
1 3
14 9 9 9 1 11 13 3 1 9 0 9 15 9 2
10 0 9 0 9 13 12 9 2 9 2
20 0 0 9 4 13 1 9 9 12 2 3 11 3 13 1 12 9 2 9 2
7 0 9 9 13 11 7 11
12 0 9 13 1 11 3 7 3 12 9 9 2
4 11 11 2 11
9 1 0 9 15 15 3 13 9 2
23 13 1 0 0 9 2 15 13 3 3 3 12 7 15 13 1 12 0 9 1 15 9 2
18 3 13 9 1 3 12 9 9 2 15 13 3 3 16 1 12 9 2
25 3 3 3 13 13 10 9 1 3 15 9 2 7 12 12 9 13 9 9 1 12 3 0 9 2
19 0 9 9 0 9 13 12 9 9 2 1 15 3 9 15 13 1 9 2
8 10 0 9 13 12 9 9 2
15 16 4 0 9 9 13 2 13 4 15 13 0 11 3 2
10 9 13 9 1 12 0 9 7 9 2
55 10 9 13 9 7 9 0 9 2 13 9 1 0 9 12 2 15 12 2 9 13 0 9 9 0 9 1 9 7 9 2 11 2 2 7 15 13 9 7 9 2 16 4 13 0 9 1 0 0 9 2 15 13 9 2
29 9 9 3 13 13 1 15 2 16 0 9 4 3 3 13 7 16 1 10 9 13 0 9 0 9 2 13 11 2
22 9 13 0 9 1 15 2 16 1 0 12 9 0 9 13 3 3 16 0 0 9 2
14 9 10 0 0 9 3 13 12 0 9 9 7 9 2
22 10 0 0 9 13 0 9 0 0 9 2 15 1 9 12 13 0 9 12 9 9 2
15 3 7 13 9 0 3 0 0 9 0 7 0 0 9 2
10 1 9 12 13 0 9 12 9 9 2
22 1 0 9 12 9 9 2 15 0 9 3 13 1 9 2 13 3 16 12 1 11 2
20 9 11 13 2 16 0 9 9 13 3 0 9 2 3 3 13 12 9 9 2
36 1 0 9 13 11 1 12 9 9 2 15 15 13 1 10 0 9 15 2 16 9 3 13 1 9 0 12 0 9 1 0 9 12 9 9 2
19 3 12 9 9 13 1 14 9 3 15 0 9 1 0 11 7 0 11 2
14 1 11 3 13 12 0 9 2 11 2 11 7 11 2
15 16 9 15 3 13 11 15 2 16 15 3 13 0 9 2
33 0 9 11 2 11 2 0 2 11 7 11 13 9 1 0 0 9 2 16 13 10 9 7 13 15 1 9 9 1 3 0 9 2
19 1 0 11 13 1 9 0 2 3 0 9 11 7 1 0 9 3 11 2
30 1 11 2 3 15 13 3 15 0 9 2 13 14 9 2 14 12 9 9 3 2 15 13 3 2 16 13 3 11 2
25 0 7 0 11 13 3 0 9 2 1 15 3 13 3 12 9 9 2 7 3 15 16 1 11 2
19 0 9 0 9 1 10 9 1 9 9 15 13 1 9 14 12 9 9 2
7 0 12 9 13 3 13 2
14 11 2 11 7 11 13 3 3 16 12 12 15 9 2
33 9 11 13 2 16 10 0 9 13 0 7 0 0 9 7 0 0 9 2 15 4 13 13 0 9 2 16 4 3 13 10 9 2
33 13 15 7 2 16 13 1 0 9 10 9 1 0 11 2 7 3 14 1 0 9 9 9 0 9 1 9 13 9 1 0 9 2
24 0 9 13 12 1 0 0 9 2 7 3 13 12 9 9 2 15 13 12 9 15 0 9 2
7 7 15 13 14 9 9 2
39 9 13 9 10 9 9 2 0 9 2 15 13 13 9 7 13 15 9 1 9 1 9 2 16 13 0 13 15 1 9 7 15 13 2 15 1 15 13 2
25 3 0 0 9 11 13 1 10 0 9 14 12 9 2 16 1 0 9 1 15 13 12 0 9 2
20 1 9 1 10 0 9 13 13 2 16 0 9 3 13 9 3 12 9 9 2
6 9 0 9 0 9 13
15 0 9 4 13 4 1 9 9 13 9 0 9 1 11 2
33 13 15 0 9 2 15 3 13 2 16 0 9 13 1 0 9 12 9 9 2 12 9 2 9 2 2 15 3 0 9 3 13 2
20 0 9 13 0 9 1 9 0 9 1 0 9 9 9 0 9 9 11 11 2
29 1 0 0 9 13 2 16 4 0 9 2 1 15 4 13 9 0 9 2 4 13 1 9 0 9 1 0 9 2
15 13 13 2 16 4 1 0 9 13 15 0 9 0 9 2
9 0 9 13 0 9 1 0 9 2
5 3 15 7 13 2
28 0 9 2 15 9 13 0 7 0 0 0 9 2 4 13 0 9 1 0 9 2 0 0 9 7 9 3 2
26 13 15 2 16 0 9 2 16 15 4 13 9 7 4 13 9 1 10 9 2 3 13 0 0 9 2
27 11 11 2 9 9 9 7 9 0 0 9 2 9 10 9 13 7 1 0 9 15 13 1 0 9 9 2
13 1 1 0 9 9 15 9 13 3 13 0 9 2
19 0 0 0 9 7 13 9 1 0 9 0 9 0 9 0 7 0 9 2
19 0 9 15 7 13 2 16 0 9 0 9 15 13 7 3 13 0 9 2
18 1 12 1 0 9 3 9 13 0 9 7 13 13 1 9 0 9 2
15 13 3 2 2 16 4 9 13 1 10 9 13 3 3 2
9 9 13 1 9 0 9 3 0 2
14 10 9 15 13 13 9 15 2 16 13 9 9 9 2
38 13 3 2 16 10 0 9 2 15 13 1 9 9 1 3 7 3 0 9 2 13 1 0 9 13 0 9 2 15 4 13 0 13 10 9 0 9 2
3 2 11 2
9 11 13 13 9 1 0 7 0 9
9 11 13 13 0 0 9 10 9 2
21 13 15 1 9 0 0 9 11 11 2 15 3 13 3 1 9 1 0 9 9 2
17 9 1 0 0 9 0 9 7 0 9 1 0 9 15 3 13 2
24 11 15 1 10 9 13 0 0 9 2 0 1 9 0 0 9 2 9 9 9 7 9 9 2
12 9 13 2 3 4 13 1 9 0 9 13 2
20 0 11 13 10 9 1 0 0 9 0 0 9 1 9 13 9 1 0 9 2
20 9 7 13 1 9 1 0 0 9 0 0 3 0 9 0 9 2 1 0 2
21 13 3 2 3 4 0 0 9 9 13 2 13 7 9 2 16 15 3 3 13 2
18 0 0 9 13 1 0 9 2 16 9 13 9 1 9 0 0 9 2
12 13 2 16 9 9 13 1 9 9 3 0 2
12 0 9 13 1 10 9 13 15 0 0 9 2
22 9 4 13 1 15 9 1 9 0 9 0 9 2 0 1 9 3 0 9 0 9 2
28 0 0 9 13 13 10 0 9 1 0 9 1 9 0 9 2 16 13 1 9 0 9 2 0 1 9 11 2
24 1 0 11 13 11 2 15 13 3 1 9 10 9 9 1 9 0 9 2 3 13 9 11 2
22 15 3 1 11 13 0 9 2 1 15 13 13 9 0 9 1 9 12 9 2 9 2
35 9 13 0 9 1 9 0 9 2 15 11 13 9 12 0 9 2 0 12 2 1 9 1 0 9 2 15 15 13 3 1 9 1 11 2
27 9 0 9 13 0 9 1 3 0 2 16 0 9 0 9 13 1 0 9 1 0 9 7 0 9 9 2
14 9 2 15 13 1 9 12 0 9 2 13 0 9 2
37 1 0 9 13 0 13 1 0 9 1 9 3 12 9 2 1 0 0 9 2 0 0 9 7 3 0 9 2 13 7 10 9 12 9 1 9 2
28 16 0 9 0 9 13 10 9 2 13 12 1 0 9 9 0 9 1 15 16 9 2 15 13 10 0 9 2
21 3 1 0 9 2 3 15 4 11 13 3 0 9 2 16 0 0 9 3 13 2
31 3 0 9 9 13 9 9 9 1 3 0 9 2 15 13 9 3 13 1 0 0 9 2 7 15 1 12 1 12 5 2
21 15 13 1 0 9 2 10 9 4 13 1 12 9 2 9 3 7 9 0 9 2
3 2 11 2
5 11 15 13 1 11
2 11 2
20 11 13 1 9 12 12 0 9 1 11 7 11 2 15 1 9 11 13 9 2
9 13 15 3 0 9 9 11 11 2
22 1 11 4 13 12 9 2 1 11 2 1 9 9 7 1 0 9 1 9 1 11 2
14 1 11 13 12 9 2 1 0 9 7 1 0 9 2
6 9 13 13 13 1 11
2 11 2
17 9 11 11 12 2 1 9 3 3 13 2 16 10 0 9 13 2
32 0 9 11 11 3 3 1 11 13 2 16 3 13 13 9 9 11 11 12 2 1 11 2 15 4 13 1 9 12 2 9 2
20 1 9 3 9 0 11 0 9 13 2 16 15 13 13 2 16 1 15 13 2
20 13 2 16 13 13 1 9 9 2 15 4 15 3 9 13 13 1 0 11 2
18 9 1 0 9 11 13 3 0 7 13 15 9 0 9 3 1 9 2
10 13 15 9 9 1 11 11 2 11 2
37 1 9 13 11 11 12 2 1 9 0 1 0 9 13 0 0 11 3 2 0 9 2 3 13 9 1 10 12 0 9 9 13 9 1 12 9 2
8 9 15 13 13 9 2 14 9
11 0 9 9 11 11 13 1 0 9 0 9
4 11 11 2 11
12 0 9 4 15 13 13 1 0 9 0 9 2
25 1 9 0 0 9 7 9 1 0 11 1 10 9 13 9 11 11 11 1 0 9 9 11 11 2
9 0 9 1 10 9 13 11 9 2
16 2 10 9 13 1 10 9 0 9 1 9 0 9 1 11 2
15 9 1 0 7 0 9 13 3 1 0 9 1 0 9 2
24 13 2 16 15 0 2 3 16 0 2 9 13 0 9 1 11 2 3 9 0 9 4 13 2
14 2 13 3 1 12 9 10 0 9 1 9 1 9 2
2 3 2
14 13 1 15 14 10 9 2 7 7 9 7 9 0 2
9 2 1 0 9 13 11 0 9 2
14 1 9 9 7 9 4 1 0 9 13 9 0 9 2
10 3 4 13 10 9 1 0 0 9 2
8 1 11 13 0 9 3 0 2
40 13 4 12 0 9 2 0 0 9 1 9 1 9 11 2 13 9 1 11 2 0 9 1 11 1 0 9 0 9 7 1 10 9 4 15 13 7 1 11 2
5 13 15 0 9 2
4 3 16 9 2
4 13 15 9 2
10 9 1 11 13 12 1 0 1 9 2
6 3 16 9 1 11 2
4 13 3 0 2
16 2 1 9 1 0 0 9 1 0 9 13 0 9 1 11 2
8 13 2 16 15 9 13 13 2
7 13 15 1 15 3 13 2
18 13 7 0 13 9 1 9 16 15 7 9 2 15 15 13 2 9 2
9 9 15 13 13 1 9 1 9 2
10 13 0 13 3 2 13 15 13 9 2
8 9 15 13 13 3 14 9 2
7 13 15 13 9 0 9 2
12 13 13 9 2 15 9 13 2 0 7 0 2
5 11 1 11 1 11
2 11 2
17 1 0 9 13 3 1 0 9 9 0 9 11 11 1 9 11 2
13 1 3 0 9 15 12 9 13 3 10 0 9 2
17 9 7 9 15 3 13 1 9 0 0 9 7 1 9 9 0 2
33 11 2 11 11 2 11 13 1 9 9 9 9 1 0 11 7 3 1 10 9 1 11 1 9 9 11 2 15 15 13 0 9 2
14 11 9 13 1 0 9 1 11 2 1 15 15 13 2
24 9 4 1 11 2 11 13 9 9 13 1 11 7 3 3 13 9 11 2 11 7 0 11 2
36 13 4 9 3 7 3 2 13 11 7 13 2 16 15 9 13 10 0 9 2 16 13 9 0 9 7 9 11 1 9 0 9 1 0 9 2
8 10 9 13 7 11 2 11 2
21 1 0 9 13 9 9 1 9 0 1 12 2 9 2 3 13 1 9 9 11 2
16 13 15 3 3 2 16 15 13 7 13 2 13 1 9 9 2
5 9 0 9 1 11
10 0 9 7 9 13 1 0 11 1 9
4 11 11 2 11
39 9 1 9 0 9 0 9 1 15 2 3 4 1 9 13 9 1 11 7 1 10 9 2 15 1 9 13 0 9 9 0 0 9 7 9 1 0 11 2
36 9 0 9 15 13 1 9 0 2 16 4 0 9 13 3 7 1 10 9 2 16 13 1 9 7 3 13 9 0 9 15 9 1 9 3 2
16 13 3 0 9 1 9 9 0 9 1 9 0 11 1 11 2
19 0 9 13 9 9 1 11 13 1 9 2 13 1 9 9 11 11 11 2
15 13 2 16 11 13 9 1 9 1 0 9 1 9 12 2
10 13 2 3 4 11 13 13 1 9 2
18 3 15 13 3 13 15 9 2 13 1 15 11 9 11 11 1 11 2
13 13 2 16 0 13 9 0 9 11 1 9 12 2
14 1 10 9 15 3 13 13 2 15 15 13 2 13 2
12 9 0 9 9 1 11 13 3 1 0 9 2
14 13 1 9 0 0 9 7 1 0 9 9 11 11 2
11 11 1 0 9 13 0 9 9 0 9 2
9 9 4 15 13 13 7 0 9 2
13 13 7 7 1 9 10 9 2 13 11 2 11 2
22 1 9 1 11 7 11 2 1 1 10 0 9 2 9 13 1 0 9 9 11 11 2
6 13 13 9 0 9 2
20 1 15 13 9 1 0 9 11 2 11 1 11 9 9 12 2 13 0 9 2
16 11 0 9 13 10 9 9 11 1 9 0 9 1 9 11 2
17 15 2 16 11 0 0 9 1 9 12 13 2 15 1 15 13 2
1 12
2 11 11
7 9 13 9 2 7 9 2
14 13 3 0 9 9 7 9 2 0 7 10 9 13 2
13 7 13 9 1 0 9 0 9 13 1 9 9 2
15 9 3 13 3 3 9 9 2 7 0 9 2 0 9 2
11 9 9 13 2 16 15 1 0 9 13 2
16 1 9 1 0 9 2 1 0 9 2 13 9 1 0 9 2
11 15 0 9 13 3 9 1 9 1 9 2
24 9 13 1 9 0 9 2 7 13 1 9 2 16 0 9 10 9 3 13 9 0 9 13 2
9 1 10 9 15 7 9 9 13 2
5 3 13 13 0 2
13 13 9 2 16 1 9 0 9 13 1 0 9 2
18 7 3 1 9 2 16 13 13 2 16 1 15 13 14 1 0 9 2
6 10 9 13 7 0 2
20 9 1 0 0 9 7 0 0 9 11 14 3 13 9 0 9 7 0 9 2
18 0 9 7 0 9 15 9 12 9 13 9 1 0 9 1 9 9 2
37 13 2 14 11 11 9 9 11 1 9 1 0 9 0 2 13 9 0 9 7 9 2 16 3 1 15 3 13 13 2 16 13 3 11 11 1 2
10 9 13 0 9 0 9 7 0 9 2
7 15 7 4 10 9 13 2
10 7 12 1 12 9 2 7 15 9 2
11 3 7 3 15 3 13 0 9 1 9 2
21 4 2 14 9 0 9 1 11 7 11 13 2 13 15 9 16 9 9 0 9 2
16 9 9 11 2 16 0 11 11 3 13 0 9 2 13 0 2
26 3 4 13 1 12 9 0 9 1 9 9 2 15 4 13 12 9 1 0 9 1 0 9 0 9 2
17 0 9 13 13 3 0 3 2 15 0 9 10 9 3 0 13 2
3 9 14 13
2 11 2
32 1 1 9 0 9 11 7 11 13 0 9 0 13 15 1 9 0 9 2 1 15 13 9 9 1 11 7 11 1 0 9 2
10 11 15 3 13 0 9 9 11 11 2
12 1 12 2 9 4 13 9 13 1 0 9 2
2 0 9
2 11 2
7 9 13 9 1 9 9 2
17 13 15 9 0 9 0 9 1 0 0 9 0 1 9 9 9 2
13 13 4 12 9 7 1 15 9 9 3 13 9 2
9 12 13 9 3 1 12 9 9 2
5 0 9 1 0 11
2 11 2
27 0 9 4 12 2 9 1 9 0 9 0 11 13 14 1 12 2 3 1 12 2 3 13 13 1 9 2
21 0 9 11 3 13 2 16 9 9 9 2 0 3 1 12 2 9 2 13 13 2
29 9 1 9 2 15 13 1 0 9 2 13 9 13 1 0 9 1 0 9 2 0 9 7 1 0 9 1 11 2
13 0 9 1 9 13 0 9 7 13 10 0 9 2
44 1 11 0 9 4 12 2 12 2 3 13 0 9 1 0 11 2 9 12 2 2 15 13 1 11 1 11 2 11 2 11 1 11 2 11 2 11 2 11 7 11 1 11 2
8 0 9 4 13 3 1 9 2
4 9 9 1 11
5 11 2 11 2 2
18 9 9 2 15 13 11 1 9 1 9 2 13 0 9 0 0 9 2
12 1 12 9 13 1 0 0 9 12 9 9 2
27 3 0 13 9 9 0 9 1 11 9 3 7 3 9 1 9 0 9 2 1 0 11 4 13 9 9 2
21 15 0 13 1 9 2 12 2 13 9 11 11 2 11 1 9 11 1 0 11 2
11 1 0 9 13 3 7 1 9 0 9 2
26 1 1 15 2 16 0 9 1 11 1 11 15 13 0 15 9 14 1 10 9 2 13 9 9 9 2
5 0 9 1 0 9
5 11 2 11 2 2
28 1 0 0 9 9 9 1 11 0 1 3 0 9 3 13 12 9 1 0 11 1 9 1 12 1 12 9 2
23 1 9 2 3 3 13 9 0 9 2 1 15 9 11 13 9 9 9 2 11 2 11 2
9 1 9 13 7 12 9 1 11 2
8 1 12 9 9 3 13 9 2
12 3 1 9 9 4 1 0 9 13 12 9 2
29 1 11 15 0 9 7 9 1 0 0 9 3 13 2 7 0 9 13 1 9 9 2 13 7 9 9 7 9 2
48 1 9 9 13 3 0 9 0 9 7 0 9 2 7 1 9 9 2 15 13 3 12 2 13 1 9 9 0 9 2 3 1 9 1 11 2 16 0 9 13 9 1 0 9 2 13 11 2
20 1 9 0 9 7 0 0 0 9 13 9 0 9 13 1 9 1 9 11 2
10 9 15 7 13 7 1 0 0 9 2
12 0 9 0 9 13 4 3 3 13 3 1 15
5 11 2 11 2 2
16 0 9 16 0 9 0 9 4 3 3 3 13 7 1 15 2
7 1 9 15 3 3 13 2
23 13 13 9 2 15 4 3 3 13 2 16 1 9 0 9 4 13 13 15 1 10 9 2
14 16 15 7 15 0 9 13 2 13 15 1 15 13 2
13 13 1 9 7 13 1 9 2 1 15 13 0 2
15 3 13 9 2 16 0 9 10 9 13 0 7 0 13 2
9 1 10 9 9 13 3 0 9 2
12 13 13 0 2 7 13 3 13 12 9 3 2
40 13 4 15 1 0 9 1 3 0 9 2 16 3 13 9 1 9 10 9 1 0 9 0 9 7 0 0 9 2 13 11 9 9 9 7 0 9 11 11 2
10 3 7 1 0 9 15 1 9 13 2
20 3 15 3 13 9 13 1 15 9 2 15 13 1 0 9 2 13 11 11 2
26 1 9 9 9 1 0 9 4 13 2 16 4 0 9 13 1 9 2 15 13 9 1 0 9 13 2
21 9 9 7 0 9 13 10 0 9 7 0 9 16 0 9 0 9 1 15 13 2
11 9 1 0 9 4 13 4 13 3 3 2
17 13 15 2 16 1 9 0 9 4 13 0 9 13 10 9 13 2
17 1 10 9 4 9 10 9 13 2 13 0 9 1 9 0 9 2
6 1 9 13 14 13 9
2 11 2
25 0 9 4 13 10 0 9 13 1 15 2 16 4 9 13 10 9 9 2 15 13 0 3 13 2
34 1 10 9 1 0 9 1 9 11 1 11 2 15 15 13 12 2 7 12 2 9 2 15 13 9 0 9 9 7 0 9 11 11 2
14 1 12 9 15 15 13 7 0 9 1 9 11 11 2
11 1 11 7 0 9 13 13 0 9 9 2
28 9 13 2 16 13 0 9 16 9 0 9 7 13 2 16 15 13 9 13 1 15 2 16 4 15 13 3 2
27 3 13 2 16 1 9 7 0 9 2 15 7 13 1 10 9 13 1 0 0 9 2 4 13 13 9 2
14 1 9 1 11 15 13 9 7 9 9 1 0 9 2
36 4 15 13 14 9 9 2 7 3 9 9 7 9 9 2 9 9 2 10 9 1 9 2 0 0 9 2 9 7 9 0 9 1 0 9 2
4 9 9 9 2
5 11 2 11 2 2
11 9 0 9 9 11 11 13 13 3 0 2
8 13 15 0 0 9 11 11 2
30 13 2 16 16 13 9 0 1 9 2 15 1 9 0 9 13 0 9 7 3 4 13 2 3 13 1 3 0 9 2
48 9 0 1 0 9 4 1 10 9 13 13 2 16 9 9 9 2 15 15 13 1 15 0 2 13 1 10 9 2 3 2 1 0 9 2 7 16 4 3 3 13 0 9 1 9 1 9 2
23 0 9 11 11 2 2 12 2 4 3 13 1 15 2 16 9 0 13 0 9 0 9 2
4 9 0 9 13
5 11 2 11 2 2
19 0 9 11 11 13 1 9 3 1 0 9 0 0 9 1 0 0 9 2
23 0 0 9 13 10 9 3 1 9 9 2 7 15 1 12 9 2 15 13 9 0 9 2
18 9 13 9 9 0 0 9 11 11 7 0 9 0 1 11 11 11 2
7 9 13 0 9 0 11 2
10 0 9 3 13 13 1 9 9 12 2
6 0 9 4 15 13 13
4 11 1 11 2
26 0 9 13 1 0 0 9 11 11 9 0 9 9 2 15 15 13 12 2 9 1 0 9 1 11 2
11 9 3 13 9 11 2 11 7 9 13 2
54 11 4 15 1 9 9 9 13 13 14 15 0 2 7 7 10 9 2 15 13 10 9 0 9 10 9 13 1 0 9 2 3 0 15 9 2 7 1 0 9 7 11 2 10 9 4 0 0 9 1 9 9 13 2
18 4 2 14 3 13 0 9 11 13 2 13 9 9 15 9 1 9 2
21 9 9 0 9 1 9 12 7 12 13 1 9 1 9 9 11 1 0 9 11 2
23 9 13 3 0 9 9 2 0 0 9 2 7 9 2 15 13 9 11 11 1 11 11 2
21 1 0 9 1 11 7 0 9 13 13 12 9 9 11 2 15 13 1 0 9 2
11 9 9 15 13 7 11 11 7 11 11 2
9 1 9 11 11 1 9 0 9 2
5 9 11 2 11 11
1 3
23 9 12 9 2 0 3 12 9 9 2 13 3 3 1 9 1 11 1 0 9 0 11 2
12 9 11 15 13 9 9 0 9 11 2 11 2
24 0 9 3 13 12 2 9 2 3 3 1 9 2 3 0 0 0 9 13 9 1 0 9 2
14 3 4 15 1 10 9 13 0 9 13 1 12 9 2
35 9 12 9 2 15 12 2 12 2 12 13 1 9 1 0 0 9 11 1 11 1 11 2 13 1 9 1 11 0 7 9 1 0 9 2
4 0 9 1 9
3 0 11 2
33 1 9 15 13 0 9 9 1 11 1 9 0 9 1 11 7 11 1 0 9 2 15 13 0 9 0 9 11 7 11 1 11 2
24 9 9 0 11 11 11 3 13 9 1 9 9 2 7 1 15 13 1 0 9 7 0 9 2
14 10 9 13 9 16 15 2 3 13 9 1 0 9 2
13 3 12 9 9 9 13 0 9 1 9 1 9 2
15 1 0 9 1 0 9 3 1 9 13 9 0 9 0 2
18 9 15 13 7 0 9 0 0 9 1 9 11 11 11 11 2 11 2
5 11 1 11 13 11
2 11 2
24 9 1 9 11 11 2 11 11 7 0 0 9 0 0 11 13 3 9 1 9 9 11 11 2
10 15 10 9 1 11 3 13 0 9 2
12 9 6 11 4 13 16 9 11 3 1 9 2
31 9 1 0 2 3 0 11 11 13 0 0 9 9 13 2 16 3 13 1 12 9 2 3 13 1 9 0 9 0 11 2
38 0 9 11 2 15 3 1 9 11 1 9 13 2 13 2 16 9 13 0 2 1 9 9 13 3 3 0 9 11 1 10 9 11 7 9 0 11 2
4 0 9 1 11
2 11 2
36 9 0 7 0 0 9 1 9 1 0 9 0 9 11 13 0 9 9 9 0 9 1 0 9 11 11 1 11 11 2 9 0 9 0 9 2
10 11 13 1 11 1 9 1 0 9 2
19 1 9 9 13 12 9 9 1 9 9 7 9 1 9 9 1 0 9 2
10 1 9 13 11 1 9 0 9 11 2
8 0 9 14 2 7 2 2 2
11 9 1 0 9 9 11 13 14 1 9 9
5 11 2 11 2 2
24 3 3 16 9 15 9 0 0 9 13 1 9 0 9 11 1 9 0 9 0 9 0 9 2
14 1 10 9 13 3 9 9 7 9 1 0 9 9 2
20 9 11 13 1 0 9 10 9 9 9 11 11 7 9 0 9 9 11 11 2
23 9 11 3 13 15 2 16 9 13 9 13 1 15 2 16 9 4 3 13 9 10 9 2
16 3 1 0 9 14 10 0 9 13 1 9 9 7 9 9 2
20 0 9 1 9 11 13 1 11 0 9 9 2 15 13 2 1 15 13 9 2
17 1 9 11 10 0 9 10 9 13 13 2 9 9 15 13 11 2
20 1 9 0 9 11 11 2 11 2 13 0 9 3 0 9 1 3 0 9 2
12 0 9 4 3 3 13 4 13 7 9 9 2
25 1 0 9 9 13 7 14 9 2 0 9 15 3 13 13 13 2 1 15 15 7 9 13 3 2
16 9 9 9 11 11 11 13 9 13 3 0 9 9 0 9 2
20 7 0 9 7 1 15 13 2 16 9 13 0 9 2 7 13 7 13 9 2
16 0 9 0 9 16 0 9 13 1 10 9 0 9 1 9 2
17 9 11 13 14 0 9 2 15 13 13 11 1 9 1 0 9 2
11 7 0 9 0 9 15 1 9 11 13 2
12 1 11 11 15 1 0 9 13 3 3 13 2
18 7 1 9 9 4 14 13 0 3 1 9 12 3 0 9 0 9 2
9 1 11 11 13 0 9 9 9 2
15 0 9 4 13 9 13 1 9 0 9 7 9 9 9 2
3 11 13 9
2 11 2
15 1 11 1 11 13 1 0 9 12 2 9 9 0 9 2
26 0 9 15 1 10 9 13 3 12 2 9 7 9 13 7 1 9 1 9 0 9 1 11 11 11 2
11 13 15 3 9 9 11 11 2 11 2 2
12 10 9 4 13 0 9 13 9 9 11 11 2
36 9 2 3 15 1 11 13 13 0 9 2 13 0 9 1 9 9 2 9 0 9 13 1 9 3 9 0 7 0 13 1 9 1 0 9 2
18 9 13 2 16 9 3 13 15 9 2 3 0 9 1 0 9 13 2
17 0 9 13 1 9 1 12 9 1 11 2 11 7 11 2 11 2
18 9 13 9 13 0 7 3 15 9 1 9 10 9 13 2 13 9 2
5 0 9 9 9 11
2 11 2
27 3 10 9 7 9 9 13 9 13 1 0 9 9 11 2 15 15 13 12 2 9 1 9 10 0 9 2
24 1 9 0 9 4 15 1 9 13 13 3 2 9 11 2 9 11 7 11 7 9 0 9 2
33 1 0 9 13 13 12 9 2 9 1 12 9 7 1 12 9 2 9 2 1 15 15 13 7 9 2 7 3 0 7 0 9 2
14 9 9 9 13 1 0 11 12 2 3 0 1 9 2
6 1 9 13 0 9 2
1 9
4 0 9 3 14
10 9 0 9 15 13 3 1 9 0 9
7 11 2 11 2 11 2 2
12 11 1 10 9 11 11 13 9 13 0 9 2
30 1 9 0 9 15 14 13 7 1 9 2 7 13 1 9 9 0 2 9 1 3 13 2 16 9 9 9 0 13 2
19 7 0 9 9 14 13 0 2 9 9 1 0 9 4 13 13 3 0 2
10 9 13 9 13 2 10 0 9 13 2
16 0 9 13 2 16 9 4 13 13 9 13 1 9 10 9 2
20 1 9 2 10 9 13 11 0 2 11 13 2 16 13 15 9 0 9 9 2
13 13 9 2 15 4 15 3 13 2 7 3 13 2
10 3 10 9 13 1 15 3 3 13 2
10 3 15 13 3 1 6 9 7 11 2
10 9 0 9 13 1 0 9 3 0 2
29 13 15 9 1 15 2 16 0 9 9 1 0 9 3 13 2 3 16 9 2 15 15 13 1 9 13 1 9 2
16 11 13 14 9 9 3 13 2 7 3 13 1 11 3 0 2
12 13 13 9 2 15 14 1 0 9 3 13 2
25 13 1 9 13 2 16 1 10 9 13 0 9 2 15 13 1 0 9 1 0 9 2 13 11 2
10 9 0 9 1 10 9 13 11 11 2
20 13 15 2 16 1 0 9 15 13 13 7 0 9 2 16 13 7 3 0 2
31 13 3 1 0 9 2 15 15 13 9 0 0 9 1 0 9 13 2 7 15 13 10 9 13 2 13 13 11 2 11 2
9 1 9 13 9 0 9 9 0 9
2 11 2
35 1 0 9 1 9 0 0 9 0 9 2 15 9 13 2 13 9 0 9 3 9 9 11 2 15 13 2 16 15 9 13 0 0 9 2
29 9 9 2 10 9 9 9 11 13 2 4 1 0 9 9 0 9 11 11 13 4 1 10 9 13 1 9 9 2
17 1 10 9 4 13 4 13 7 1 12 9 9 13 3 0 9 2
22 9 11 2 11 9 13 2 16 3 13 9 2 15 13 7 3 2 7 13 2 3 2
22 9 9 1 15 3 13 0 9 7 1 9 9 7 9 9 1 9 0 9 1 9 2
15 3 1 0 9 13 9 9 0 9 9 2 15 13 9 2
24 13 2 16 15 1 9 0 9 0 9 4 13 0 9 13 13 9 2 15 13 13 10 9 2
37 9 0 9 15 1 10 9 13 9 2 16 13 1 10 0 9 2 16 13 13 1 9 7 9 0 9 2 15 15 13 10 0 9 3 12 9 2
6 11 15 13 1 9 9
5 11 2 11 2 2
22 9 9 2 0 9 7 9 0 9 9 1 9 13 0 9 0 1 0 9 0 9 2
25 13 7 1 0 15 9 0 9 1 9 7 0 9 9 0 1 9 2 3 1 0 2 9 9 2
13 1 12 9 13 0 9 13 9 9 9 1 9 2
33 4 13 2 16 4 15 0 9 11 2 15 0 9 13 2 3 9 1 9 9 9 7 9 1 9 9 2 13 9 0 0 9 2
13 13 15 3 13 1 9 0 9 1 9 7 9 2
13 1 0 9 4 13 13 9 9 1 9 7 9 2
4 11 1 9 9
3 1 0 9
5 11 2 11 2 2
21 11 13 1 9 11 11 13 3 13 1 9 9 7 13 1 10 9 1 9 9 2
16 1 9 0 9 13 11 9 0 9 0 9 1 0 0 9 2
20 1 0 9 4 9 3 13 1 15 0 0 9 7 14 1 12 9 0 9 2
20 1 9 0 0 9 11 1 11 1 11 13 11 9 9 1 0 9 7 9 2
7 11 2 1 9 13 13 11
3 1 0 9
2 11 2
32 3 11 2 7 3 0 9 13 13 1 9 7 13 15 1 3 0 9 0 9 2 9 13 9 11 1 9 9 13 0 9 2
15 9 9 11 11 11 15 13 1 9 1 0 0 9 9 2
9 1 0 9 13 11 13 0 9 2
26 11 3 13 2 16 9 4 3 13 9 0 9 0 9 2 0 9 10 9 7 0 9 0 0 9 2
7 11 2 1 0 11 12 9
3 1 0 9
4 11 1 11 2
17 3 12 9 1 0 9 13 13 11 1 12 9 7 9 0 9 2
10 13 15 9 0 0 9 9 11 11 2
14 12 12 1 15 13 9 11 2 0 13 1 0 9 2
9 13 1 15 7 12 0 9 11 2
11 1 11 7 15 1 15 13 10 0 9 2
17 15 9 2 15 15 1 9 11 1 0 11 13 2 4 3 13 2
24 1 9 13 11 1 11 1 11 1 11 2 11 2 11 7 11 2 16 11 4 13 0 9 2
5 0 9 7 9 9
3 13 13 2
4 9 2 11 11
38 9 15 13 2 13 2 14 0 9 2 16 4 13 9 0 9 1 9 1 9 1 9 1 9 2 3 0 9 13 1 0 9 3 9 7 3 9 2
27 16 1 0 9 13 9 13 9 0 2 13 15 15 2 16 13 13 9 2 15 13 3 9 16 0 9 2
10 9 13 1 9 9 9 2 7 13 2
23 10 9 13 0 7 13 1 15 2 16 1 11 0 0 0 9 15 13 3 0 9 9 2
24 13 7 1 15 2 16 0 9 13 0 9 2 3 3 7 9 1 9 9 0 9 7 9 2
21 16 4 15 9 13 14 3 1 9 1 10 9 2 13 4 15 14 1 0 9 2
16 13 7 3 2 16 7 1 15 9 9 13 2 16 4 13 2
18 9 12 9 2 12 9 13 0 9 1 0 9 9 7 9 1 15 2
35 9 12 9 2 12 9 13 2 16 0 13 9 1 9 7 9 2 12 10 9 13 2 16 9 13 9 1 0 9 1 0 7 0 9 2
23 7 3 9 2 12 9 2 12 9 3 2 13 2 16 0 9 15 13 15 1 9 9 2
6 9 13 10 0 9 2
39 0 13 9 2 16 16 9 13 1 0 9 0 9 16 0 9 2 4 15 13 12 1 0 9 2 2 4 1 9 13 3 7 14 3 2 16 13 9 2
22 13 0 2 16 1 0 9 4 0 9 3 13 15 1 3 0 9 9 0 0 9 2
4 3 15 13 2
51 9 9 1 0 0 9 2 15 3 13 9 2 1 15 13 13 9 13 15 2 16 4 9 0 9 4 13 9 2 13 7 9 9 9 2 16 7 9 0 9 1 9 1 9 9 1 9 1 0 9 2
42 13 15 1 0 9 2 13 15 2 13 2 16 9 2 12 9 2 12 9 13 2 16 1 9 9 13 4 13 9 9 9 0 9 0 15 0 9 7 9 0 9 2
16 9 0 9 9 1 0 0 9 13 1 10 9 3 16 0 2
46 1 9 12 9 2 12 9 2 9 2 9 1 0 9 13 13 13 0 9 3 2 0 9 2 16 13 2 16 0 9 9 0 9 4 13 10 3 0 0 9 2 1 12 9 2 2
26 1 15 7 13 13 15 0 0 9 0 9 1 9 10 9 2 7 2 1 0 9 9 1 0 9 2
20 16 4 3 0 9 13 2 16 1 9 3 0 9 13 2 13 4 0 9 2
10 0 9 13 9 0 9 1 0 9 2
45 13 1 15 2 16 1 9 3 13 2 16 13 1 0 0 9 13 13 9 0 2 15 3 13 0 0 9 2 0 16 9 1 0 9 2 7 9 3 0 0 9 1 0 9 2
17 0 9 2 9 9 1 9 0 9 0 9 13 1 9 1 9 2
44 1 9 13 3 3 13 2 16 9 13 9 13 0 9 0 0 9 3 2 16 4 13 3 0 9 0 10 9 13 3 9 10 10 9 13 1 9 0 9 2 7 2 3 2
10 7 15 9 13 13 1 0 0 9 2
26 16 4 15 1 9 0 9 1 0 9 13 7 13 0 9 1 0 9 1 9 2 15 13 13 15 2
26 13 1 9 2 1 15 13 2 16 10 9 13 9 0 0 9 2 7 9 1 0 9 0 0 9 2
27 9 13 0 0 7 0 9 2 7 13 1 15 9 2 1 0 0 9 2 3 7 3 0 9 0 9 2
15 1 10 9 15 10 9 13 0 0 2 14 0 0 9 2
22 1 11 2 16 13 0 0 9 3 13 3 2 13 0 9 1 9 1 0 9 9 2
20 11 15 3 13 3 2 7 13 0 9 2 3 16 4 9 13 13 0 9 2
3 9 1 9
1 9
2 11 11
17 9 1 10 0 9 13 0 9 13 1 0 9 9 9 7 9 2
32 7 16 13 1 9 11 11 1 11 11 13 10 9 2 3 3 0 9 12 10 9 2 0 0 9 2 13 3 14 0 9 2
14 13 15 2 16 0 9 0 9 13 7 1 9 13 2
24 9 0 2 0 2 0 2 2 15 1 0 9 9 3 10 9 13 2 13 3 0 0 9 2
39 13 15 13 2 16 0 9 1 0 0 9 2 16 15 13 0 9 0 9 2 13 0 9 2 15 13 13 0 9 1 0 0 9 9 1 9 0 9 2
16 10 0 9 13 3 9 9 2 15 3 1 9 13 10 9 2
16 3 0 9 7 1 0 9 13 3 9 0 9 9 11 11 2
23 15 3 13 1 9 1 9 0 9 2 16 4 13 1 9 0 0 9 1 10 0 9 2
16 13 7 1 0 9 13 0 9 1 9 0 9 1 9 12 2
44 1 10 9 13 9 0 2 0 2 0 2 1 9 9 2 16 4 13 15 9 1 9 0 9 11 2 15 10 0 9 13 1 0 12 2 9 2 3 4 13 9 0 9 2
30 16 9 0 2 0 2 0 2 13 2 16 15 1 10 9 1 9 9 11 11 13 1 10 9 2 13 13 3 13 2
27 9 9 3 13 9 10 9 7 13 2 16 10 0 9 15 0 2 0 2 0 2 7 9 9 13 3 2
40 9 9 1 15 2 16 0 9 7 9 1 10 9 3 0 13 13 0 9 14 3 2 16 15 13 9 2 3 7 3 1 9 9 13 0 9 3 15 13 2
7 0 9 7 13 13 9 2
23 9 10 9 3 13 3 3 9 2 16 13 2 16 0 9 13 13 3 15 16 10 9 2
18 16 4 3 13 1 9 0 9 2 1 15 1 0 9 0 9 13 2
5 0 9 11 13 9
12 0 11 15 13 1 11 2 1 15 9 1 9
4 11 11 2 11
19 0 11 13 1 0 2 7 3 3 0 9 9 1 11 1 0 9 11 2
16 1 0 9 15 0 9 13 1 11 7 0 9 13 1 15 2
29 1 9 13 0 2 16 0 11 13 1 0 9 2 15 15 1 9 12 7 12 13 12 9 9 2 14 9 0 2
4 7 14 3 2
11 0 9 11 13 2 0 9 1 9 2 2
17 7 9 0 3 1 0 9 2 1 9 1 0 9 7 1 9 2
29 3 1 0 9 7 9 9 1 9 1 0 0 9 0 2 11 4 15 7 13 2 16 9 13 3 3 0 9 2
21 14 3 13 11 0 9 11 11 2 7 7 15 3 13 9 2 0 9 11 2 2
25 0 9 12 9 13 1 9 9 9 0 2 16 15 11 4 3 3 13 1 9 7 1 10 9 2
23 10 0 9 4 15 13 13 11 11 2 11 11 2 7 1 0 9 7 3 0 0 11 2
29 9 9 11 11 3 3 13 2 16 15 1 9 1 0 9 13 1 9 9 7 9 0 9 4 13 13 12 9 2
33 9 11 13 2 16 11 13 3 0 9 16 0 11 7 11 7 1 9 1 0 9 1 0 9 1 11 4 15 13 13 1 9 2
26 1 9 4 11 13 1 12 9 1 9 12 2 12 7 12 9 1 9 12 2 12 2 3 12 9 2
10 0 9 13 1 0 9 1 0 9 2
10 9 13 3 9 1 0 2 0 9 2
23 0 9 13 3 9 1 12 1 12 9 2 9 2 12 9 2 7 16 15 13 0 9 2
25 9 0 9 2 12 2 12 9 2 9 2 2 9 2 13 12 2 12 7 12 9 1 12 9 2
19 3 0 13 7 9 7 1 0 9 7 9 10 9 3 13 9 0 9 2
8 1 15 13 7 0 0 9 2
7 11 13 7 3 0 9 2
19 1 9 13 9 0 9 1 9 9 7 9 7 1 0 9 13 7 9 2
14 11 3 13 7 13 1 0 9 9 9 12 11 11 2
10 9 0 9 13 1 9 11 3 0 2
13 0 9 15 3 1 15 13 1 11 11 7 11 2
15 3 0 0 9 0 9 15 13 1 0 9 1 9 9 2
17 9 9 3 13 0 0 9 2 1 0 9 13 7 3 0 9 2
16 1 9 1 9 12 9 13 0 13 7 0 2 7 0 9 2
8 11 13 1 15 3 0 9 2
14 7 3 1 9 1 9 14 0 9 13 1 12 9 2
6 7 15 13 1 0 2
5 9 7 0 0 9
5 11 11 2 9 9
6 3 3 13 0 9 2
12 3 13 0 9 7 3 15 13 1 0 9 2
14 12 9 9 3 13 1 9 9 2 3 1 9 9 2
8 13 0 9 2 13 15 13 2
10 13 0 9 0 9 2 13 15 13 2
9 13 0 0 9 2 13 15 13 2
22 13 0 0 9 16 9 0 9 2 13 4 10 9 1 9 1 11 13 1 0 9 2
20 13 0 9 2 13 1 11 2 13 7 9 13 0 9 0 9 10 0 9 2
8 13 9 2 13 13 9 9 2
11 13 4 13 2 7 15 4 15 3 13 2
51 0 9 15 13 2 16 13 0 9 2 16 13 0 7 0 2 1 12 9 0 2 9 2 16 13 0 9 1 0 9 2 1 9 2 1 9 0 9 2 1 0 9 2 1 10 7 15 3 0 9 2
12 15 15 9 3 13 2 13 15 7 9 0 2
15 1 9 3 13 15 1 15 7 3 15 13 13 1 12 2
29 3 16 1 9 9 2 9 2 0 9 7 0 9 2 7 1 9 9 13 2 16 13 13 3 2 16 15 13 2
5 13 15 3 13 2
30 7 3 3 13 12 0 9 2 15 2 15 9 13 7 4 13 1 9 2 13 3 9 15 2 1 15 13 3 13 2
7 1 9 13 15 7 3 2
19 9 13 13 3 2 16 13 2 3 7 1 9 2 9 9 9 3 13 2
30 10 9 15 2 9 2 3 13 2 7 13 2 16 3 10 9 15 9 7 10 9 4 0 9 13 1 9 0 9 2
38 0 9 9 13 1 9 9 13 0 0 9 2 9 0 9 2 10 0 9 2 7 3 10 0 9 1 9 2 15 4 1 9 9 1 9 3 13 2
12 13 4 3 13 2 16 15 14 3 13 15 2
38 9 1 9 7 9 13 7 1 15 2 7 3 3 1 15 2 16 16 9 13 1 15 15 2 1 9 9 13 9 9 7 10 9 3 13 7 13 2
56 12 0 9 13 15 0 2 12 9 0 2 7 7 13 10 0 9 13 0 9 1 9 2 3 1 9 9 2 9 2 9 2 10 9 2 16 4 9 4 9 13 2 16 4 13 0 9 0 9 9 0 2 7 14 0 2
10 0 9 10 0 9 13 9 0 9 2
20 9 13 3 3 3 13 1 9 7 13 3 3 1 15 2 7 15 3 3 2
18 15 15 13 0 9 7 0 9 1 9 0 9 13 14 12 1 15 2
43 9 1 9 13 3 7 3 3 3 7 3 1 0 9 9 13 9 10 9 3 3 13 3 0 0 9 2 7 15 3 13 9 1 9 9 13 1 9 1 0 0 9 2
53 14 3 13 1 10 9 3 7 15 2 1 9 2 3 15 3 13 13 0 0 9 3 15 13 0 9 2 13 0 9 0 9 7 3 15 13 13 7 3 15 1 10 9 15 13 13 2 16 9 3 13 3 2
26 7 13 9 9 9 1 0 0 9 2 7 15 3 9 0 0 9 16 3 0 9 1 0 0 9 2
15 0 9 13 2 13 7 4 3 13 1 9 3 0 9 2
50 3 10 9 1 10 9 0 11 2 0 11 2 11 2 12 2 13 0 0 9 2 0 9 9 2 9 1 9 9 12 2 12 11 11 2 1 10 0 9 13 15 0 7 3 4 15 15 13 0 2
53 3 1 9 12 4 12 9 10 9 13 0 0 9 2 11 2 11 2 12 2 13 0 9 9 7 13 4 2 16 4 1 10 9 9 1 11 11 13 2 16 1 9 9 13 1 0 9 2 7 1 0 9 2
42 11 11 7 13 1 0 11 13 14 1 0 9 0 9 2 7 7 1 0 9 9 0 9 2 15 13 15 2 15 1 15 13 1 0 9 7 15 13 10 0 9 2
7 3 3 13 12 0 9 2
31 3 3 4 1 0 9 2 13 1 9 0 9 2 13 9 0 0 9 1 9 15 2 16 13 3 9 1 15 7 15 2
33 9 0 9 3 13 7 13 13 9 9 9 2 16 9 15 9 13 2 3 15 13 2 1 9 10 9 2 1 0 9 1 9 2
42 9 0 9 4 10 9 13 1 0 2 9 0 9 2 3 1 9 2 3 9 3 13 2 7 13 3 7 0 2 7 0 2 9 13 3 9 10 9 13 1 9 2
9 13 13 2 16 15 13 10 9 2
18 0 9 10 9 13 9 9 2 7 16 15 15 3 3 3 15 13 2
4 9 0 9 13
2 11 11
18 9 0 9 4 1 9 11 11 13 9 9 1 9 9 1 0 9 2
8 11 13 1 9 3 12 9 2
9 3 12 9 13 3 9 1 9 2
26 13 15 0 13 1 9 1 9 1 0 0 9 9 1 0 9 2 15 15 3 13 1 9 0 9 2
3 7 0 2
12 13 2 16 9 9 13 0 1 9 9 13 2
9 0 16 9 9 13 3 9 9 2
20 16 4 11 1 9 13 2 14 4 13 0 2 0 9 1 12 1 12 9 2
9 0 9 13 1 9 9 3 13 2
13 0 9 2 16 0 9 2 13 0 1 9 9 2
10 15 0 9 2 15 0 9 1 9 2
25 13 7 9 2 16 1 0 9 0 9 4 15 13 2 7 7 13 7 9 2 15 1 9 13 2
16 13 15 15 9 9 2 16 3 13 3 0 9 7 3 9 2
21 10 9 1 9 2 16 15 11 13 1 9 9 2 13 7 15 9 7 9 9 2
12 7 15 0 9 1 9 9 9 13 9 9 2
9 1 9 0 11 7 10 0 9 2
23 9 1 9 0 9 0 9 13 3 3 1 9 9 2 16 1 15 0 9 3 3 13 2
39 0 11 15 13 1 9 9 2 16 3 16 1 9 9 9 2 3 15 13 9 2 15 3 16 0 9 13 3 1 9 1 9 7 9 1 3 0 9 2
8 9 1 9 9 13 3 9 2
12 9 1 9 4 3 1 11 13 13 14 9 2
21 3 0 9 9 4 15 13 7 10 9 2 1 15 9 1 0 9 13 14 13 2
21 3 0 13 7 9 2 16 1 0 9 9 7 9 1 9 9 13 0 0 9 2
20 13 0 2 3 9 7 9 13 13 0 9 9 2 7 15 7 0 9 9 2
11 0 9 9 1 15 15 13 1 12 9 2
9 3 12 1 15 13 1 0 9 2
19 9 2 15 13 0 9 1 0 9 2 13 0 1 0 9 0 0 9 2
12 11 15 3 1 9 9 13 13 2 15 13 2
20 15 3 13 9 0 0 9 2 7 0 9 9 15 10 9 13 0 1 9 2
40 7 13 0 2 16 9 9 2 3 9 2 15 1 9 13 9 1 0 9 9 2 13 1 15 1 9 1 0 9 3 0 2 16 13 0 9 10 0 9 2
29 0 9 2 15 2 16 13 1 0 9 2 7 13 15 3 13 1 0 9 2 13 9 9 7 1 15 0 9 2
17 13 1 9 2 0 9 13 1 9 9 0 9 1 9 0 9 2
13 9 2 13 7 10 9 2 3 0 9 9 13 2
2 7 2
11 1 15 1 15 15 13 9 13 9 9 2
13 1 10 9 4 9 0 9 13 7 0 9 9 2
13 1 10 9 0 9 13 13 9 3 1 0 9 2
22 13 15 3 14 0 9 2 7 7 1 0 11 13 9 9 9 0 7 3 15 0 2
15 3 1 15 10 9 13 9 1 0 9 14 9 0 9 2
10 11 2 0 0 9 9 2 9 13 2
13 1 11 9 0 9 1 9 0 0 9 3 13 2
17 10 9 2 3 11 13 9 15 0 1 15 9 2 13 3 0 2
23 3 15 13 9 2 16 11 13 13 3 15 2 16 13 13 0 9 0 9 16 9 0 2
7 15 13 7 9 3 0 2
17 0 9 0 9 3 13 13 2 16 0 9 9 4 3 13 9 2
8 3 0 0 9 11 3 13 2
11 13 9 1 3 3 0 0 9 1 0 2
10 9 1 9 13 11 1 9 10 9 2
17 0 9 1 9 13 7 0 9 9 2 15 13 1 0 0 9 2
24 9 3 0 0 9 3 11 13 1 0 7 3 0 9 2 3 13 3 3 9 16 9 0 2
18 9 9 4 14 13 0 9 11 7 0 9 4 4 13 1 9 0 2
7 9 15 10 9 3 13 2
5 11 2 9 7 15
1 9
2 11 11
18 0 9 9 9 11 11 11 13 0 9 11 2 11 2 11 7 11 2
22 3 0 9 9 13 12 2 13 0 2 3 0 9 7 13 15 1 9 9 0 9 2
6 15 15 3 13 13 2
14 0 9 9 7 13 1 9 0 1 9 7 1 9 2
15 15 15 13 1 11 13 1 9 0 9 7 1 9 9 2
16 13 4 15 7 13 9 3 0 7 0 9 11 1 10 9 2
9 10 9 13 1 0 9 3 0 2
18 13 9 9 11 1 9 13 9 0 9 14 1 0 2 0 0 9 2
19 13 0 9 9 7 9 9 13 0 2 9 0 9 13 3 0 9 9 2
18 13 13 2 16 15 4 1 0 9 13 1 10 0 9 3 3 13 2
24 1 10 9 13 3 0 0 9 1 11 7 9 1 9 9 11 11 2 9 11 7 0 9 2
32 0 0 9 2 3 7 0 9 0 9 7 0 9 2 13 0 9 3 13 1 9 2 15 13 15 1 11 7 15 3 13 2
9 0 9 9 1 11 13 3 0 2
16 14 12 13 3 0 2 1 0 0 9 0 9 13 9 3 2
35 9 15 13 3 1 15 2 10 9 4 13 2 10 9 1 15 4 13 12 9 0 1 0 2 0 9 7 13 2 14 15 1 0 9 2
25 1 0 11 15 3 13 14 1 9 10 9 2 1 9 13 7 9 0 2 0 9 11 7 9 2
28 13 4 3 3 2 16 4 0 9 3 10 9 2 9 7 9 2 1 15 15 13 2 10 9 3 3 13 2
4 0 9 1 11
1 9
2 11 11
25 3 0 0 11 15 13 1 0 0 9 13 9 1 9 9 1 9 9 11 7 9 1 0 9 2
50 0 9 9 13 9 3 0 9 9 0 1 9 0 9 11 2 15 4 13 1 12 9 0 2 0 9 2 12 9 0 0 9 7 9 9 9 11 11 2 11 2 15 13 16 9 0 9 0 9 2
29 9 4 13 3 1 15 2 16 0 9 1 15 13 9 9 0 9 11 2 0 9 7 9 0 0 9 11 11 2
35 10 9 2 16 13 3 1 9 1 9 11 11 2 13 9 0 7 1 9 15 13 7 1 15 2 16 4 13 0 9 1 9 0 9 2
9 15 15 7 0 9 13 16 0 2
24 3 16 11 2 11 2 7 0 9 1 0 9 0 9 11 13 1 0 9 10 7 15 9 2
15 13 3 0 2 16 1 9 13 1 9 9 9 10 9 2
23 1 9 3 0 0 9 2 15 13 0 3 0 9 9 11 11 2 13 13 1 0 9 2
17 0 9 7 0 9 2 9 11 11 2 9 11 2 13 0 9 2
30 3 0 9 13 9 9 1 9 11 2 3 7 9 3 2 15 15 1 9 9 13 3 1 10 9 11 11 13 9 2
16 13 7 13 2 16 15 12 13 1 0 9 13 1 0 9 2
25 0 9 15 13 3 1 9 13 1 0 11 0 9 3 2 16 4 3 1 12 9 13 1 9 2
17 13 15 3 14 1 0 9 9 1 0 9 2 0 1 10 9 2
22 12 1 0 9 13 3 0 9 3 0 9 0 11 2 15 13 1 9 9 0 9 2
21 1 10 9 15 13 0 9 13 9 1 10 9 0 9 7 13 9 1 10 9 2
6 11 13 9 9 1 11
5 11 2 0 11 2
30 0 9 9 11 11 13 2 16 10 9 13 10 9 1 0 9 11 1 11 2 16 4 13 9 1 9 9 0 9 2
32 10 9 13 1 9 2 15 4 13 1 10 9 1 9 1 11 7 11 2 15 15 13 9 0 9 2 7 13 4 14 3 2
12 11 13 1 0 11 0 9 1 9 12 9 2
29 9 11 4 13 2 16 11 13 1 0 9 9 1 9 9 7 1 0 9 13 2 3 3 16 3 2 13 11 2
36 11 3 13 11 2 16 13 1 9 0 9 1 0 9 2 7 3 13 3 3 2 16 13 11 2 15 13 9 0 9 10 0 9 1 11 2
45 16 3 13 9 0 0 11 1 9 1 0 9 1 0 9 2 0 9 11 13 0 9 1 11 7 11 1 9 2 10 0 9 13 1 9 0 9 2 16 4 4 13 9 9 2
43 0 9 11 11 7 9 0 0 9 1 0 11 11 11 7 11 11 13 3 1 11 0 9 9 1 0 0 9 2 11 2 1 0 9 0 9 1 9 1 11 7 11 2
3 11 13 9
5 11 2 11 2 2
16 0 0 9 0 9 13 9 9 9 16 9 1 9 0 9 2
8 9 13 1 9 0 9 11 2
18 13 3 2 16 0 9 11 11 1 10 9 3 13 0 9 11 11 2
9 13 15 3 2 3 11 13 9 2
7 11 15 3 13 9 1 9
4 11 2 11 2
25 0 0 9 2 11 2 15 13 15 10 9 2 16 4 13 9 0 0 9 1 9 0 9 9 2
12 13 15 3 1 9 11 0 3 0 9 11 2
28 1 0 0 9 11 13 14 12 9 9 7 9 2 1 15 9 1 0 9 9 13 1 0 9 1 0 9 2
18 0 9 13 3 9 11 2 0 0 9 11 2 11 2 7 0 11 2
23 0 3 0 9 2 11 2 2 15 9 13 1 9 11 1 11 2 4 3 13 13 9 2
12 1 9 1 0 9 1 11 15 13 9 11 2
15 9 1 9 0 9 13 11 3 9 10 9 2 13 9 2
20 11 15 1 9 12 13 1 11 7 4 13 1 0 0 9 0 1 0 11 2
13 1 9 9 13 0 9 1 11 0 9 11 11 2
13 3 13 2 16 0 9 13 10 0 9 1 11 2
27 11 15 1 9 1 0 11 13 13 0 9 2 16 9 11 13 2 16 4 11 13 1 9 11 1 11 2
30 3 13 2 16 0 9 13 13 9 2 16 9 11 13 0 2 16 4 13 13 9 1 9 11 11 2 0 9 11 2
30 0 9 11 11 13 2 16 10 9 13 1 0 9 1 0 9 1 9 13 15 2 16 4 13 11 7 13 0 9 2
22 13 1 0 0 9 2 7 1 9 1 9 2 7 15 1 12 9 2 9 7 9 2
19 1 9 1 0 9 11 11 13 2 16 0 9 1 0 9 13 3 11 2
18 0 9 13 2 16 15 0 9 13 1 11 11 2 9 9 11 11 2
28 9 11 11 11 15 13 10 9 13 1 11 1 9 11 2 11 2 16 4 1 15 13 1 0 9 1 11 2
3 11 13 11
2 11 2
19 9 1 11 13 3 9 10 9 1 0 9 2 13 3 0 9 11 11 2
17 13 3 9 11 2 16 0 9 1 11 13 14 9 9 11 11 2
20 11 13 3 9 0 9 11 7 13 0 9 2 16 4 13 0 9 1 11 2
23 0 9 7 11 13 1 9 9 2 0 13 3 12 0 9 1 0 0 9 1 0 9 2
11 0 12 9 13 4 1 11 13 3 3 2
20 0 9 15 3 13 13 10 0 9 11 1 11 2 3 4 9 9 3 13 2
9 1 0 9 15 9 9 3 13 2
13 11 11 15 7 13 7 1 0 9 2 0 9 2
1 9
9 11 15 13 9 1 9 1 9 9
4 9 11 2 11
5 11 2 9 13 9
4 11 2 11 2
25 0 9 11 2 11 1 11 3 13 1 9 0 9 2 11 2 2 15 13 9 0 0 0 9 2
23 9 13 15 0 16 9 0 1 9 2 13 11 7 13 2 16 10 9 13 7 13 0 2
33 9 0 9 2 11 2 11 11 3 1 0 0 9 9 1 11 13 9 1 15 2 16 11 13 1 9 13 0 9 1 9 11 2
29 13 9 1 9 9 1 0 0 9 2 15 13 0 9 9 0 0 9 2 11 2 2 15 15 3 13 1 11 2
14 9 13 1 0 0 9 1 0 9 3 13 1 15 2
19 9 9 11 11 13 1 10 9 2 16 11 13 3 11 2 11 7 11 2
17 1 0 9 11 4 15 10 9 13 13 9 0 9 1 9 12 2
25 1 9 0 9 0 0 9 15 13 9 0 0 0 9 2 11 2 2 15 1 9 13 1 11 2
17 1 9 9 13 9 9 0 9 2 1 15 15 13 1 0 9 2
4 12 11 9 0
39 12 0 11 1 9 11 2 0 1 0 9 11 2 4 0 9 0 13 1 9 1 12 9 9 1 0 9 1 9 2 1 12 1 9 1 0 9 11 2
15 9 13 9 1 9 9 13 1 0 9 0 9 9 11 2
41 12 0 9 2 0 1 9 2 9 7 9 9 0 9 2 13 1 15 1 9 3 0 12 9 7 9 1 9 0 9 2 0 9 7 9 9 1 0 10 9 2
5 1 11 0 9 11
2 11 2
19 11 13 1 11 0 9 2 15 4 13 13 0 9 1 10 0 9 0 2
15 13 15 3 9 0 9 7 9 0 9 9 9 11 11 2
49 1 9 13 11 3 3 0 9 1 11 2 3 7 13 13 1 0 0 9 7 3 1 0 9 9 9 2 11 2 16 9 0 9 2 13 11 7 13 2 16 3 4 13 9 9 1 0 9 2
16 9 9 11 11 11 13 10 9 1 11 2 0 1 0 9 2
19 9 9 9 13 9 2 16 11 13 13 9 0 1 9 1 11 7 11 2
17 0 9 0 9 1 11 13 9 9 7 9 1 15 13 3 3 2
17 15 13 1 9 0 0 0 11 0 9 0 9 9 9 7 9 2
8 0 9 15 13 0 9 1 11
2 9 11
4 9 1 0 9
9 0 0 9 15 13 1 11 1 11
7 11 11 2 11 11 2 11
24 1 12 9 15 0 9 1 9 11 13 3 9 2 3 11 13 9 2 15 15 13 1 11 2
17 1 9 3 2 12 2 9 12 2 3 13 0 0 9 1 11 2
11 0 12 9 9 0 9 9 15 13 3 2
25 1 9 11 11 2 15 9 1 0 9 9 15 3 13 2 1 9 1 9 13 0 9 11 11 2
30 1 9 9 9 11 15 13 14 9 0 9 11 2 11 7 1 0 9 11 13 10 9 13 14 12 7 9 9 9 2
28 1 15 14 12 9 13 15 13 2 7 13 10 9 1 9 0 9 7 13 9 0 9 9 9 2 13 15 2
18 7 9 11 13 2 9 0 9 9 1 11 13 0 0 7 0 9 2
19 13 9 2 16 9 13 15 1 10 2 16 4 3 13 0 9 1 9 2
12 11 1 12 7 9 9 13 1 11 12 9 2
17 1 15 13 12 9 2 9 13 9 9 1 12 9 7 0 9 2
13 1 9 13 0 9 0 9 0 9 9 9 11 2
15 13 2 16 9 0 9 13 13 9 0 9 1 0 9 2
23 9 0 9 11 11 13 9 9 1 9 9 0 7 0 9 2 1 15 11 13 9 9 2
12 13 15 9 2 7 0 9 0 9 2 13 2
28 1 3 0 9 13 0 9 0 9 11 2 11 9 11 2 13 4 0 9 9 2 15 3 13 9 1 9 2
9 10 9 13 9 9 2 13 11 2
27 1 15 13 11 11 2 15 13 9 1 11 2 13 1 9 9 2 16 1 15 9 4 13 1 11 9 2
10 0 9 15 13 14 9 0 1 11 2
18 1 9 12 15 1 11 13 1 9 3 16 12 9 7 10 0 9 2
17 1 0 9 4 1 15 13 3 12 9 2 12 9 7 12 9 2
18 11 3 13 12 9 9 1 9 9 2 1 9 9 7 1 9 9 2
14 3 13 1 10 9 12 9 0 9 1 9 1 9 2
25 9 9 11 11 11 3 13 2 16 1 9 0 9 4 13 12 0 0 9 1 9 11 7 11 2
15 1 0 9 4 3 13 0 9 1 11 7 1 0 11 2
26 12 1 9 0 9 9 11 11 13 9 0 9 1 11 9 2 13 1 9 2 7 1 0 0 9 2
21 11 2 15 15 13 1 0 0 9 2 13 10 0 9 1 10 0 7 0 9 2
18 0 9 9 13 1 10 9 0 1 12 9 13 9 11 7 0 9 2
10 3 10 3 0 9 13 9 1 9 2
9 7 13 15 2 16 13 15 13 2
22 3 1 11 1 0 9 2 15 15 11 3 13 2 13 10 9 3 16 9 9 9 2
15 14 16 15 13 10 10 9 1 0 9 3 1 10 9 2
1 3
35 11 11 2 0 9 9 2 13 3 9 3 2 16 4 3 0 9 13 1 9 1 9 1 9 9 0 9 11 11 1 0 15 0 9 2
35 11 11 2 0 9 0 9 2 13 1 9 0 9 2 16 13 0 9 2 15 15 1 9 0 9 13 1 9 1 9 0 9 11 11 2
15 9 1 9 11 1 9 7 9 11 15 3 13 12 0 2
32 9 1 0 9 11 13 9 0 9 1 0 9 11 2 13 3 1 11 1 12 2 9 9 9 9 9 9 0 9 11 11 2
21 1 0 9 11 1 0 9 2 15 0 9 13 1 9 12 2 13 12 9 11 2
16 12 12 9 13 1 0 9 7 12 9 13 1 10 0 9 2
18 1 9 2 15 13 9 1 11 1 9 12 9 2 13 3 0 9 2
35 9 0 9 1 0 11 9 9 0 11 13 1 9 9 0 0 9 13 1 0 9 0 9 1 9 12 9 0 0 9 1 11 7 11 2
38 9 11 13 1 9 9 0 2 16 0 9 15 1 9 1 9 11 13 9 2 16 9 0 1 0 0 9 1 9 12 2 12 13 4 13 0 9 2
18 13 15 9 1 9 11 11 2 16 11 3 1 9 12 13 9 11 2
5 9 9 1 9 9
10 1 11 3 13 0 9 1 9 7 9
2 11 11
1 9
12 3 9 13 2 16 9 15 13 1 0 9 2
50 9 1 0 9 13 0 9 11 11 9 9 2 15 1 0 9 13 7 13 9 9 9 11 2 9 7 9 2 0 13 9 1 9 0 9 1 9 7 9 2 11 12 2 2 15 3 13 1 11 2
50 13 2 14 10 9 1 0 9 0 9 7 13 15 1 9 1 15 0 9 7 9 2 3 13 3 3 2 13 9 0 9 3 13 2 10 9 13 13 1 9 2 1 10 0 9 1 9 3 13 2
4 7 13 9 2
17 16 10 9 3 3 13 2 9 3 15 13 13 3 0 7 0 2
26 1 9 13 2 16 4 13 9 1 9 9 9 0 9 2 7 15 13 13 9 9 9 1 0 9 2
14 3 13 2 16 4 13 9 1 9 9 7 0 9 2
18 13 15 13 9 9 12 9 1 9 3 2 16 4 0 9 13 12 2
22 3 1 12 9 13 1 12 9 12 9 2 3 3 3 16 12 2 3 3 12 2 2
10 13 15 15 16 0 9 0 0 9 2
22 7 3 0 9 2 12 9 1 12 9 2 13 0 9 3 3 3 0 2 1 11 2
12 9 13 2 3 13 15 9 9 9 12 9 2
49 16 15 13 0 9 9 2 3 0 9 2 16 13 9 0 2 4 13 1 15 12 9 9 2 7 1 9 9 2 1 9 12 2 14 3 3 16 9 12 2 1 12 9 2 16 14 3 3 2
42 1 10 9 15 13 9 2 16 0 9 13 3 2 10 9 13 3 0 2 12 5 9 11 13 0 12 9 2 7 0 0 2 12 5 9 11 13 1 12 9 2 2
46 14 12 5 1 0 9 9 15 1 9 12 9 13 1 0 9 9 2 1 11 2 11 2 0 11 2 11 2 16 1 0 9 9 13 2 7 3 13 2 11 2 11 2 11 2 2
39 13 3 13 2 16 9 2 15 3 13 1 9 1 0 9 2 13 1 9 10 9 12 2 12 7 3 9 2 9 3 2 2 16 10 9 1 0 9 2
31 9 13 10 9 1 15 10 0 9 15 13 2 1 0 9 2 1 0 9 1 11 1 9 12 7 11 11 1 9 12 2
7 1 0 9 13 1 9 2
10 0 9 1 11 7 0 9 1 11 2
18 1 9 0 9 9 1 0 9 13 0 9 9 2 0 9 13 9 2
32 1 12 9 9 9 2 3 9 7 0 9 1 0 9 13 1 9 7 9 3 9 13 9 2 15 13 13 9 1 0 9 2
33 0 9 4 13 3 3 2 1 0 9 3 1 0 9 2 13 15 0 1 9 7 9 2 1 0 9 7 3 0 7 0 9 2
2 9 2
12 9 15 13 7 3 15 13 0 9 12 9 2
30 1 11 15 13 9 2 13 15 4 1 12 7 12 9 2 1 9 9 9 2 7 9 2 7 0 2 9 7 9 2
27 1 9 9 13 0 9 11 12 1 0 9 2 3 13 0 7 0 9 7 13 0 9 1 9 0 9 2
52 0 9 9 13 13 0 9 1 9 12 2 12 1 9 1 12 0 3 0 9 2 2 9 2 12 5 1 12 9 0 9 13 9 7 1 12 9 9 2 15 13 0 9 2 13 12 5 1 9 2 2 2
43 2 9 9 9 2 9 7 9 2 3 9 9 9 2 1 15 12 5 1 0 9 2 13 3 1 9 9 2 0 9 7 9 2 16 3 15 10 9 4 15 13 13 2
18 9 9 13 1 0 9 14 12 7 0 16 1 9 0 9 2 2 2
11 2 9 0 9 1 9 1 9 0 9 2
27 0 9 9 2 7 16 15 10 9 1 9 12 2 9 3 13 2 13 3 3 0 3 1 12 9 9 2
34 0 9 13 0 2 0 2 0 2 7 0 2 9 1 10 9 15 13 13 9 1 12 9 9 1 9 12 1 12 9 1 9 12 2
31 14 7 0 9 9 2 0 11 7 11 13 2 3 14 15 13 13 2 16 9 13 3 3 7 9 3 0 16 9 9 2
16 1 0 2 0 9 11 11 15 3 1 9 13 9 1 9 2
13 1 15 15 1 9 13 0 9 7 0 0 9 2
13 1 0 0 9 3 13 13 7 13 3 1 9 2
2 9 9
4 11 1 0 9
2 11 2
18 1 12 9 0 9 1 11 7 11 13 3 11 13 1 11 0 9 2
16 13 15 0 0 9 9 11 11 2 15 15 9 13 0 9 2
36 1 9 1 9 0 9 0 9 13 0 9 2 16 4 13 13 9 1 11 1 9 1 9 9 11 1 0 9 1 9 0 9 1 9 12 2
35 11 13 7 13 10 9 0 15 9 2 3 0 2 15 13 3 1 0 9 0 3 1 9 1 11 9 11 2 11 7 11 2 13 11 2
22 9 1 10 9 13 2 16 13 0 13 0 9 0 9 2 16 4 10 9 3 13 2
22 11 3 13 2 16 11 13 13 15 1 9 9 1 11 2 3 7 1 9 0 9 2
26 13 3 2 16 9 9 1 11 4 1 10 9 13 13 1 9 9 9 1 0 2 0 7 0 11 2
3 9 11 0
6 9 11 0 9 1 11
7 0 9 11 1 11 11 11
26 7 4 0 9 1 11 13 2 7 3 13 9 2 13 1 0 9 9 9 0 9 10 9 11 11 2
13 9 0 9 9 0 9 11 13 10 9 13 3 2
11 7 9 2 1 15 13 2 13 3 0 2
21 9 1 11 15 13 0 9 9 11 3 2 16 13 3 0 9 11 2 11 11 2
11 9 0 9 7 10 0 9 13 11 11 2
18 3 15 11 3 1 9 3 3 13 0 7 0 9 13 9 1 9 2
18 9 9 9 11 11 11 9 0 9 2 16 4 3 13 9 2 13 2
23 16 13 1 9 0 9 0 9 2 4 9 11 7 10 9 13 7 13 1 9 0 9 2
14 9 11 13 2 16 1 9 9 13 9 13 0 9 2
17 1 0 9 4 13 9 9 3 1 9 0 0 9 7 0 9 2
14 9 13 2 16 1 10 9 13 0 13 12 12 9 2
18 14 0 9 13 13 0 9 1 0 9 7 0 9 2 7 0 9 2
7 9 0 9 13 3 0 2
7 12 0 9 13 12 9 2
11 1 9 9 15 7 13 3 3 12 9 2
15 9 9 9 7 0 9 15 0 9 13 0 0 0 9 2
15 7 11 11 2 7 11 11 15 1 0 9 9 13 13 2
20 13 15 7 13 2 16 7 3 13 0 9 1 11 2 1 2 11 1 9 2
4 15 4 3 13
31 13 9 2 15 4 1 10 9 3 13 2 13 0 9 2 15 9 3 3 13 2 3 9 2 15 13 4 13 0 9 2
10 11 11 1 9 1 0 9 0 11 2
13 9 13 11 1 11 10 9 2 11 3 1 11 2
4 15 13 15 2
4 11 11 3 2
17 13 9 2 16 11 13 1 0 9 1 0 9 2 3 15 13 2
10 10 0 9 13 11 3 16 15 0 2
9 0 9 11 11 1 9 0 11 2
14 2 15 1 15 15 13 13 0 2 3 13 9 11 2
28 15 13 2 16 15 13 0 2 7 0 9 9 0 9 2 1 0 15 13 0 9 0 1 9 1 10 9 2
49 0 9 2 7 0 9 16 10 9 2 4 13 13 3 7 3 13 1 9 1 0 11 7 1 10 9 2 16 4 9 13 1 10 9 2 16 4 15 13 13 9 2 15 4 13 9 10 9 2
17 11 11 2 0 9 9 0 9 2 1 9 1 9 11 0 11 2
16 9 13 2 0 9 13 2 7 7 13 0 9 16 15 15 2
45 1 10 9 2 16 9 13 9 7 9 0 10 9 13 15 16 0 9 2 16 9 1 0 9 2 7 15 13 1 9 2 13 15 0 1 0 9 2 1 15 15 13 9 9 2
11 11 2 11 11 2 9 0 9 14 2 11
7 0 9 0 9 1 0 9
9 11 11 2 9 2 0 9 0 9
18 13 1 0 2 16 9 0 9 3 3 13 13 10 9 1 0 9 2
28 9 13 0 0 9 1 9 12 7 3 0 0 9 9 1 0 9 1 9 12 7 0 9 11 1 9 12 2
35 7 1 12 9 2 15 13 1 9 10 0 9 2 7 1 12 9 1 9 11 2 2 13 0 2 7 3 7 0 2 13 10 0 9 2
22 9 9 13 1 0 0 7 0 9 3 2 16 13 9 1 9 2 15 15 13 9 2
20 15 15 3 3 1 15 13 2 3 3 15 0 9 9 13 1 15 0 9 2
54 15 2 16 9 3 15 0 9 13 1 9 2 15 3 13 2 1 10 9 13 15 15 2 16 11 2 11 2 11 7 11 3 13 2 3 13 0 9 13 2 7 13 3 0 9 2 16 4 15 13 1 11 13 2
25 9 16 9 13 0 9 9 1 11 7 0 0 0 9 2 1 10 9 15 13 2 1 10 9 2
24 10 9 2 9 2 3 13 0 9 2 7 15 15 3 13 2 9 15 7 7 13 15 13 2
21 1 0 9 4 15 9 9 1 9 9 13 1 9 0 9 11 11 7 10 9 2
21 9 0 9 3 10 9 13 1 9 0 0 9 2 15 13 1 0 9 14 13 2
12 13 7 0 2 16 3 3 9 10 9 13 2
29 13 15 14 1 0 9 0 0 9 2 7 3 1 15 2 16 1 9 9 13 7 0 9 1 9 0 9 9 2
28 4 13 0 9 3 0 9 2 0 9 7 9 1 9 0 0 9 2 0 1 0 2 3 0 9 0 9 2
19 1 9 2 9 7 9 9 10 9 4 3 13 0 2 3 3 0 9 2
25 13 7 9 2 16 9 2 0 1 9 9 12 2 9 12 2 13 3 0 7 16 9 3 0 2
45 1 9 0 9 13 3 0 9 2 3 2 1 9 12 2 12 13 9 0 9 0 1 9 11 2 7 13 9 9 10 9 2 14 3 3 0 2 9 0 9 0 0 9 2 2
47 3 0 9 0 9 1 9 9 1 0 9 13 9 13 13 0 9 2 15 10 9 9 9 3 13 2 13 15 15 3 9 11 2 9 0 9 2 9 0 9 7 9 9 1 0 9 2
29 16 10 9 13 9 1 10 0 9 2 13 13 0 16 0 2 7 3 2 1 0 9 2 0 2 7 3 0 2
17 0 9 11 11 1 9 0 9 11 11 11 1 9 1 0 9 2
2 9 9
1 3
15 9 9 11 11 4 3 13 1 0 9 9 1 0 9 2
16 9 2 15 13 9 9 11 11 11 11 2 13 1 9 9 2
24 0 0 9 9 13 9 9 10 0 9 1 9 9 11 11 2 15 13 1 9 0 9 9 2
8 13 15 0 9 0 0 11 2
16 9 9 13 13 9 1 0 9 1 0 9 11 1 9 12 2
40 12 9 1 9 9 12 2 12 7 12 9 2 1 15 7 12 9 0 9 2 13 9 9 11 11 2 12 2 12 2 2 15 4 3 13 1 9 9 11 2
13 9 12 1 9 0 9 12 13 1 12 2 9 2
22 1 10 9 3 1 12 9 13 9 3 11 2 15 9 13 0 2 0 7 0 9 2
15 1 9 9 13 9 0 0 9 1 9 11 11 1 11 2
12 0 0 9 13 3 1 11 0 9 11 11 2
12 1 0 9 4 1 10 9 13 9 10 9 2
2 0 9
1 9
27 9 2 0 2 0 9 9 9 9 13 15 9 1 15 2 16 4 11 0 1 0 9 13 10 0 9 2
48 0 0 0 9 2 15 1 11 13 0 9 11 11 2 3 3 1 9 0 9 13 9 0 0 9 2 9 0 1 11 10 0 9 1 9 0 9 7 9 0 9 2 3 9 7 9 2 2
31 7 16 9 13 3 2 15 0 4 1 10 9 3 3 13 2 2 9 13 0 9 1 9 2 13 15 1 0 12 9 2
12 9 2 1 15 14 9 1 9 0 9 13 2
22 11 7 1 0 9 9 3 13 2 7 1 9 3 3 13 1 9 1 0 9 0 2
6 15 15 11 3 13 2
7 9 13 9 7 0 9 2
33 11 11 1 9 13 3 7 9 7 9 15 1 10 9 13 9 0 9 2 13 4 2 13 2 16 15 15 13 1 9 3 13 2
40 10 9 1 9 13 3 0 1 9 0 9 2 9 2 7 3 7 9 2 11 11 15 13 1 9 3 0 9 2 7 13 2 13 15 9 7 3 7 9 2
56 13 2 14 1 15 0 9 11 11 2 0 9 0 9 7 10 9 13 9 9 2 15 13 3 3 0 7 0 9 2 13 15 2 16 9 13 3 3 9 1 9 16 3 7 13 1 0 11 7 11 1 9 1 0 9 2
27 11 11 15 1 9 13 2 13 15 1 15 2 16 4 9 9 7 9 13 1 0 9 3 0 16 3 2
16 7 7 3 15 9 1 10 9 13 2 13 2 13 7 13 2
11 13 2 16 4 15 15 1 10 9 13 2
9 9 11 1 15 7 13 0 9 2
22 13 2 16 4 9 13 0 7 3 0 2 7 16 1 9 13 3 0 9 1 11 2
33 1 0 9 13 0 9 0 9 2 13 9 11 1 11 7 9 9 2 9 11 2 11 2 11 2 7 9 0 1 9 0 9 2
8 0 9 3 13 0 9 9 2
16 0 9 13 2 13 15 2 0 2 3 15 3 13 1 9 2
21 1 15 15 9 3 13 7 13 1 9 7 9 2 3 2 3 15 1 15 13 2
9 3 15 3 3 13 3 12 9 2
7 11 11 2 11 9 9 2
5 11 11 2 9 2
7 9 2 11 12 2 9 2
6 9 9 2 0 11 2
8 9 0 9 2 12 2 9 2
4 1 9 1 11
1 9
2 11 11
11 9 0 0 9 1 11 15 13 1 9 2
43 0 0 9 2 1 0 9 0 9 7 9 2 1 15 7 9 9 13 9 0 2 9 7 9 2 2 0 9 9 1 9 2 13 1 9 0 0 9 16 9 1 0 2
46 16 4 15 7 13 2 1 0 14 3 2 16 13 9 1 9 3 0 2 7 3 3 2 16 15 1 15 1 12 0 9 0 9 13 10 0 7 3 0 0 9 1 9 0 9 2
36 0 9 13 3 0 7 16 13 1 9 14 0 2 15 4 3 2 1 0 9 15 3 13 1 11 7 1 11 0 9 13 9 2 13 13 2
18 0 9 9 1 9 13 3 2 9 3 13 9 7 9 1 0 9 2
4 13 15 15 2
8 0 9 3 9 1 11 13 2
34 13 2 16 11 15 2 15 13 1 9 9 2 7 15 2 10 13 0 9 0 9 2 4 13 2 13 15 1 9 12 9 11 11 2
9 15 3 7 0 13 9 2 2 2
22 13 15 1 9 9 7 9 0 9 7 13 3 1 12 0 9 2 12 7 12 2 2
20 1 9 1 9 0 13 14 0 9 2 7 9 15 13 7 1 0 9 13 2
30 3 13 3 9 3 0 2 7 15 14 1 9 0 9 2 7 7 1 0 9 7 1 10 9 2 2 3 3 13 2
24 9 13 11 2 9 1 9 7 9 7 1 9 11 2 12 13 13 2 0 9 1 0 9 2
19 13 2 11 3 2 13 10 0 2 16 0 9 2 3 13 1 10 9 2
23 16 15 0 2 12 7 12 2 13 9 15 13 3 1 0 9 2 15 0 3 13 3 2
25 3 3 13 0 9 9 3 0 2 7 0 9 7 1 15 1 10 9 13 2 13 3 1 11 2
19 1 11 7 3 13 1 0 9 7 7 3 1 15 13 1 9 0 9 2
7 13 14 1 9 9 9 2
26 13 2 14 7 10 9 0 9 9 2 15 15 3 13 14 1 9 2 7 15 13 3 7 3 2 2
3 9 1 9
5 11 11 11 12 11
3 9 0 9
2 11 11
20 11 11 13 3 13 0 9 1 3 9 2 15 13 1 0 0 9 0 9 2
23 7 3 15 2 15 0 13 7 13 13 3 14 9 2 7 7 9 0 9 7 0 9 2
17 9 11 0 9 15 1 0 9 13 9 1 0 9 1 9 11 2
12 3 4 1 9 13 2 15 13 9 3 13 2
28 3 15 4 13 0 9 1 9 2 0 9 1 3 9 2 1 0 2 16 15 13 2 3 13 0 12 9 2
27 1 9 10 0 9 0 12 0 9 2 9 1 9 1 9 7 1 0 9 3 3 1 12 12 9 3 2
16 13 15 7 3 0 9 2 7 9 1 15 3 13 1 15 2
15 7 3 13 2 13 2 14 0 1 0 2 3 0 9 2
40 16 9 1 9 12 9 13 9 2 14 2 12 9 2 12 9 2 2 13 9 3 12 7 9 9 0 9 1 12 1 12 9 2 9 2 12 9 3 0 2
24 0 9 0 9 13 0 0 9 14 3 0 9 9 1 12 0 9 2 7 7 3 0 9 2
42 9 13 1 12 2 12 9 2 9 2 7 1 9 9 12 2 12 2 3 12 9 9 1 12 9 7 9 0 9 12 9 15 13 2 16 4 13 1 0 9 3 2
7 11 13 3 3 0 9 2
18 1 0 13 0 9 1 9 1 9 0 9 7 12 9 1 9 9 2
29 1 10 9 3 13 3 0 9 2 7 15 13 13 9 2 16 4 13 1 9 2 15 13 13 7 0 12 9 2
16 9 9 13 9 2 7 7 15 9 13 3 16 1 0 9 2
27 3 1 9 15 9 13 13 13 1 9 3 0 9 2 10 9 13 1 12 9 1 15 13 14 1 12 2
7 0 9 13 9 0 9 2
16 13 2 14 3 0 9 1 12 9 2 13 15 0 0 9 2
18 0 0 9 13 0 9 2 15 13 0 9 12 9 7 0 12 9 2
7 13 2 16 13 15 13 2
24 1 9 9 13 7 3 0 0 9 1 3 0 9 2 16 7 1 0 0 9 15 13 9 2
5 9 1 11 1 9
4 11 11 2 11
30 0 9 9 1 0 11 1 9 9 2 9 13 1 0 9 2 3 9 12 1 15 13 9 0 0 9 9 1 11 2
13 13 9 1 9 2 15 13 13 1 9 0 11 2
42 1 0 9 15 10 9 13 1 0 9 2 13 3 0 9 16 0 2 2 1 9 0 9 11 11 7 9 9 2 1 15 11 2 0 2 0 2 0 7 0 9 2
30 1 9 9 13 9 12 9 2 9 0 9 9 1 9 14 1 9 7 9 0 9 1 0 9 1 9 9 1 9 2
10 9 0 9 13 1 0 9 11 11 2
15 9 15 9 13 1 0 9 2 3 3 9 13 2 9 2
20 1 9 13 9 1 0 9 2 1 9 1 0 0 9 7 9 12 0 9 2
26 1 0 9 13 0 9 7 9 11 11 2 16 4 13 1 12 1 9 10 0 9 2 9 11 11 2
12 15 13 7 16 0 9 10 0 9 1 9 2
6 9 1 11 13 10 9
5 11 11 2 11 11
27 0 9 3 0 0 9 0 11 11 14 13 0 0 9 9 2 7 13 1 0 0 9 1 11 0 9 2
15 11 11 15 3 9 0 9 0 9 0 0 9 3 13 2
41 3 7 0 9 3 13 10 9 9 2 13 1 9 11 11 1 9 0 9 2 10 9 13 1 9 0 1 2 1 9 2 3 11 1 9 0 9 13 0 9 2
26 11 11 2 0 9 11 2 15 13 12 2 9 12 1 9 9 2 12 1 0 9 1 0 0 9 2
20 1 9 13 10 0 9 0 9 2 15 3 13 0 0 9 2 9 11 11 2
22 9 7 9 11 11 1 0 9 13 9 0 9 0 9 2 1 9 9 1 0 9 2
34 10 9 3 13 3 1 0 0 9 11 0 2 3 1 11 13 9 11 11 2 0 9 11 11 11 7 11 11 7 0 9 11 11 2
8 15 13 1 0 9 0 9 2
14 0 11 11 13 0 9 14 1 0 12 2 9 12 2
12 1 1 0 0 9 13 9 13 10 0 9 2
21 0 9 11 11 7 9 11 11 15 1 9 11 11 7 11 11 3 13 12 9 2
17 9 9 2 9 9 2 0 9 7 0 9 13 1 9 0 9 2
12 0 9 15 7 3 13 9 0 9 0 9 2
34 0 9 0 9 7 9 2 7 13 0 9 2 12 2 9 12 11 13 1 9 9 2 15 15 13 9 1 0 9 1 0 0 9 2
10 0 9 7 9 15 3 13 1 9 2
18 1 9 2 15 13 13 13 2 13 13 10 0 0 9 0 0 9 2
11 3 0 9 13 13 9 0 9 7 9 2
27 0 9 9 0 9 2 10 9 4 13 0 9 2 3 9 0 0 9 2 2 13 3 9 12 0 9 2
5 0 9 4 13 2
13 0 9 9 13 11 11 2 11 11 7 11 11 2
19 0 9 13 9 9 7 1 0 9 13 3 1 9 0 9 0 9 9 2
47 1 0 9 9 2 13 15 9 9 7 9 11 11 2 9 11 0 7 9 9 9 9 2 14 3 13 9 0 9 9 0 0 9 11 11 2 15 1 9 0 2 11 13 9 0 9 2
29 1 9 9 12 9 1 0 0 9 10 9 2 15 4 13 16 0 0 9 2 13 3 9 0 9 7 0 9 2
13 1 0 9 13 10 9 11 11 2 9 0 9 2
8 11 11 13 16 11 13 11 2
33 16 3 13 11 11 11 2 9 10 0 9 1 0 9 2 0 9 14 13 9 1 9 9 9 13 2 2 3 4 11 11 13 2
9 9 7 13 1 0 9 0 9 2
28 15 13 3 0 9 16 0 0 9 2 13 15 2 13 2 14 2 13 2 16 13 2 0 9 7 0 9 2
4 11 9 0 9
15 9 9 11 11 13 11 11 9 9 0 0 9 0 9 2
43 1 9 11 11 15 10 0 9 13 9 0 9 1 11 7 0 0 0 9 7 9 11 11 13 1 10 9 3 0 9 0 9 2 13 11 11 2 11 2 9 0 9 2
23 11 2 15 13 3 9 9 9 2 15 3 3 13 1 10 0 9 1 0 9 10 9 2
3 2 11 2
4 1 9 1 9
2 11 2
22 0 9 11 11 7 0 0 9 1 9 11 11 2 11 15 13 9 0 9 0 11 2
23 1 0 0 9 1 11 13 1 10 9 3 9 7 15 12 13 0 9 1 9 12 9 2
9 1 11 9 3 1 9 13 9 2
22 0 9 1 9 1 12 9 3 13 9 7 0 9 7 3 13 2 16 1 11 13 2
10 3 15 1 9 9 9 13 7 13 2
22 10 0 9 1 0 9 13 1 9 1 0 9 1 12 9 2 15 13 1 11 11 2
10 9 1 9 11 13 7 0 0 9 2
20 0 9 11 11 13 10 9 1 12 9 7 13 15 3 12 2 9 1 9 2
8 3 13 3 1 9 1 11 2
20 9 9 1 11 11 11 13 1 0 9 9 12 2 15 13 0 0 9 9 2
13 1 0 0 9 1 12 9 13 11 11 9 12 2
4 11 11 3 13
8 11 13 1 9 2 11 15 13
7 11 2 11 2 11 2 2
31 1 12 2 9 0 9 0 9 9 11 11 2 11 2 12 2 12 2 0 9 2 0 1 3 0 9 11 11 2 13 2
15 1 9 1 11 13 1 0 9 3 13 12 0 11 11 2
26 13 4 0 9 1 9 7 1 12 9 3 13 0 1 15 2 13 15 9 2 11 1 0 0 9 2
8 9 13 9 0 9 0 9 2
7 13 4 9 1 0 9 2
17 11 13 3 1 10 9 0 9 7 1 0 9 9 13 0 9 2
6 3 13 0 7 9 2
14 1 9 9 13 0 13 2 9 7 9 9 13 4 2
19 1 0 9 4 13 4 11 13 1 11 1 11 9 7 3 3 1 11 2
24 0 2 15 4 15 3 13 1 9 2 13 13 9 2 11 4 13 2 9 2 9 2 2 2
14 13 15 15 2 7 1 10 9 9 13 0 1 11 2
15 1 10 9 9 13 9 9 3 3 2 13 1 9 11 2
23 15 0 9 11 11 13 1 9 3 9 2 15 13 0 9 1 0 9 1 12 2 12 2
9 13 15 0 9 1 3 0 9 2
11 16 9 4 15 15 13 13 2 13 11 2
14 11 11 13 2 16 4 11 13 1 9 1 9 13 2
17 10 9 4 13 2 7 3 1 15 1 15 13 2 13 10 9 2
4 0 9 1 9
2 11 2
13 3 0 0 9 0 9 9 13 0 9 0 9 2
24 15 3 13 2 16 4 13 13 9 1 11 2 7 3 10 0 9 3 1 9 9 9 13 2
19 16 0 11 11 13 1 9 1 0 9 2 13 15 9 0 13 0 9 2
14 11 3 1 10 9 13 3 9 7 15 15 3 13 2
28 0 9 13 9 0 9 1 9 9 1 9 0 9 1 11 7 13 9 9 2 15 1 9 10 9 13 9 2
37 11 2 15 1 11 13 0 9 1 11 2 13 1 11 12 2 12 7 9 10 9 13 9 2 16 15 9 1 9 9 13 13 0 9 1 9 2
3 0 9 13
7 9 9 15 1 9 9 13
5 11 2 11 2 2
42 0 0 9 13 0 9 9 11 11 11 11 2 11 2 11 2 15 1 9 3 13 9 2 16 1 0 9 1 0 9 9 13 1 9 1 0 9 1 0 0 9 2
30 3 1 15 15 13 9 13 1 9 2 1 10 9 3 13 1 12 9 1 9 0 11 2 12 1 11 7 1 11 2
9 1 9 3 13 0 9 1 11 2
14 1 9 7 13 9 2 15 15 13 1 9 1 9 2
21 0 9 9 13 9 9 7 13 15 13 1 10 9 2 16 9 9 13 10 9 2
21 0 9 13 11 11 2 15 15 7 1 9 13 3 3 2 16 4 13 0 9 2
9 1 9 15 1 15 3 13 0 2
13 3 3 15 3 13 13 2 13 9 9 11 11 2
11 10 0 9 1 9 0 9 7 13 13 2
10 3 3 13 9 11 11 11 11 11 2
9 9 15 13 15 9 2 13 3 2
8 1 9 9 3 13 3 13 2
5 12 13 7 0 2
22 16 11 11 7 0 0 9 0 9 11 11 3 13 0 9 2 9 3 13 0 9 2
3 9 1 9
2 11 2
18 0 9 11 11 13 1 0 9 11 1 0 9 0 9 1 0 9 2
21 1 9 2 15 15 13 1 11 2 3 13 1 9 10 9 2 15 13 0 9 2
7 13 15 7 0 0 9 2
12 11 13 0 7 11 0 9 2 3 16 11 2
21 11 11 11 2 12 2 12 2 15 13 1 11 1 11 2 1 0 9 16 11 2
9 1 0 15 10 12 9 13 0 2
11 0 9 2 0 9 2 9 13 0 9 2
40 11 13 2 16 13 0 9 2 10 9 7 9 13 9 2 0 9 0 0 9 2 1 15 9 13 9 15 9 1 0 9 2 7 9 1 3 15 9 9 2
23 3 16 10 0 9 13 0 9 2 13 10 0 2 0 9 0 9 9 0 9 0 9 2
12 1 10 0 9 15 13 12 1 0 0 9 2
1 9
2 0 9
9 11 1 11 2 9 0 11 2 2
19 0 0 9 13 9 11 2 16 13 9 1 9 9 1 9 7 0 9 2
35 16 9 11 13 1 12 12 9 9 0 0 9 2 9 11 1 12 12 9 9 0 2 9 11 15 13 1 0 7 0 9 1 0 9 2
12 0 3 13 2 16 9 11 13 3 9 9 2
17 10 9 13 7 13 15 2 16 15 1 9 13 3 0 9 11 2
19 11 13 13 2 16 3 0 9 13 10 9 1 0 9 1 0 0 9 2
4 9 1 3 0
5 11 2 11 2 2
17 10 0 9 15 3 1 0 9 13 13 1 15 2 16 13 9 2
19 0 9 1 3 0 9 3 13 2 13 0 9 11 11 2 9 0 11 2
17 1 9 12 15 1 15 13 3 13 0 7 0 9 1 10 9 2
21 11 1 9 3 13 0 9 1 0 0 0 9 0 9 0 0 9 1 3 0 2
12 1 9 1 0 1 11 4 3 3 13 9 2
13 10 9 11 11 13 2 16 13 10 9 1 9 2
9 1 11 0 9 0 9 14 13 2
27 1 11 11 1 9 9 2 15 15 13 1 9 9 2 13 0 9 1 0 1 9 0 16 1 0 9 2
19 3 0 13 13 1 0 0 9 9 2 3 15 9 13 1 0 0 9 2
20 10 9 7 9 7 13 3 0 9 3 0 15 2 15 13 1 0 0 9 2
35 9 9 7 9 3 0 2 15 13 1 9 0 9 0 9 13 2 13 7 13 2 16 13 1 11 3 0 9 0 9 7 9 1 9 2
15 1 9 9 11 11 13 1 11 14 12 12 3 0 9 2
8 9 15 15 13 13 0 9 2
11 13 3 3 2 9 0 0 9 1 0 2
16 9 4 3 1 9 9 1 0 11 11 13 13 0 1 0 2
13 13 0 13 3 0 9 7 13 0 9 0 9 2
15 9 15 1 9 1 0 3 13 1 15 2 16 13 0 2
14 1 10 9 3 13 9 0 9 3 13 2 13 11 2
10 9 15 1 0 9 13 1 9 0 2
15 13 13 2 16 15 1 9 13 10 9 2 7 10 9 2
11 3 4 1 15 13 1 0 9 0 9 2
10 13 3 15 2 3 15 14 13 9 2
24 3 15 13 12 9 7 1 0 9 15 13 15 2 15 4 13 1 10 9 13 2 13 11 2
8 0 9 13 9 0 9 1 11
5 11 2 11 2 2
20 0 9 9 11 13 9 0 9 1 11 2 15 15 0 0 9 13 0 9 2
25 9 0 9 11 13 2 16 9 13 1 9 9 0 9 9 0 2 15 13 2 16 9 15 13 2
32 16 4 3 13 2 11 12 2 12 2 2 2 0 13 3 13 1 10 0 9 9 3 2 16 10 9 1 0 9 4 13 2
28 3 2 16 9 13 1 0 9 1 9 9 2 0 9 3 1 9 13 2 16 9 13 1 9 9 0 9 2
15 1 12 9 9 13 9 7 13 9 0 9 0 0 9 2
29 0 10 9 13 1 15 3 0 2 7 7 4 1 9 9 0 2 16 9 13 15 2 13 2 13 11 2 11 2
9 1 9 15 14 13 1 0 9 2
38 1 9 2 15 12 9 13 1 9 0 9 7 13 1 15 3 13 2 13 10 9 3 16 0 2 13 15 9 0 0 9 2 15 15 13 4 13 2
10 16 4 13 2 10 10 9 13 0 2
4 0 9 9 9
10 0 9 14 13 1 9 1 9 15 0
5 11 2 11 2 2
32 9 14 12 9 9 1 9 9 1 9 7 9 13 1 9 1 9 9 1 9 0 9 7 1 9 9 7 9 9 15 13 2
38 1 9 2 3 9 1 9 1 9 13 9 0 9 2 13 11 10 9 11 11 2 0 9 13 1 9 1 9 15 0 2 7 15 13 1 10 9 2
11 10 9 13 3 0 9 1 9 1 9 2
18 14 1 0 9 13 1 9 13 0 9 2 15 13 1 9 0 9 2
8 10 9 13 11 16 3 0 2
23 1 9 0 9 11 11 13 9 1 9 9 0 9 9 2 0 9 15 3 13 0 9 2
14 9 13 1 10 9 0 2 7 7 1 9 13 9 2
16 0 9 13 3 3 0 9 2 15 1 10 9 13 10 9 2
23 9 2 16 9 13 1 9 9 7 13 15 1 10 9 3 2 13 11 16 9 0 9 2
22 1 9 0 9 13 13 3 3 2 13 2 14 3 13 9 7 9 7 0 9 9 2
22 9 0 13 1 15 3 13 3 16 9 1 0 9 2 3 0 1 9 10 9 9 2
15 9 9 9 14 7 13 13 2 7 15 9 13 3 13 2
19 16 11 3 13 11 2 11 2 1 0 9 13 1 9 3 1 0 9 2
15 0 9 1 0 9 12 9 13 15 0 0 0 9 13 2
16 13 3 3 9 9 2 10 9 7 3 10 0 7 0 9 2
13 1 0 9 7 13 3 1 9 1 0 9 9 2
10 3 14 7 9 0 9 1 9 13 2
19 0 9 15 3 1 0 9 13 14 1 9 2 3 9 3 13 1 9 2
9 9 0 9 15 14 7 13 13 2
14 3 11 13 2 16 4 0 9 13 13 9 0 9 2
20 16 4 14 13 0 3 15 13 2 10 0 9 7 0 9 0 9 13 0 2
33 11 11 3 9 9 11 13 9 0 9 1 11 1 11 12 12 0 9 2 15 13 0 7 3 0 9 1 9 1 9 1 9 2
5 9 11 11 2 11
9 9 9 13 13 3 12 7 12 9
5 11 2 11 2 2
18 3 10 0 9 2 9 2 4 1 12 2 9 12 1 0 9 13 2
7 13 15 1 9 9 9 2
15 1 0 9 10 0 9 13 9 9 13 12 7 12 9 2
19 1 9 12 2 3 13 13 9 1 9 2 4 13 12 9 1 9 9 2
14 1 10 9 4 1 12 2 9 12 13 12 0 9 2
23 1 9 1 0 9 13 1 0 9 3 0 9 2 3 0 0 9 7 9 1 9 0 2
7 0 9 13 14 0 9 2
23 9 9 0 9 11 11 3 1 9 13 2 16 0 9 9 3 13 9 9 7 9 9 2
10 9 0 0 9 7 10 9 3 13 2
20 1 15 13 0 9 0 9 1 9 7 9 2 15 9 3 13 1 3 0 2
29 1 0 9 3 0 9 13 13 1 0 0 9 2 16 9 1 9 13 10 0 0 9 2 15 4 9 9 13 2
10 9 9 0 9 13 7 0 0 9 2
30 1 10 9 13 1 9 9 0 9 2 3 13 9 0 9 2 13 0 9 1 9 7 9 7 3 13 10 0 9 2
2 10 9
2 11 11
20 15 13 2 0 1 15 13 10 9 2 13 9 9 2 15 13 1 10 9 2
24 1 15 1 0 9 15 13 2 16 3 13 9 2 16 3 0 2 7 15 1 9 7 9 2
11 3 15 10 15 14 3 9 13 1 9 2
29 1 10 9 15 13 2 16 16 3 13 0 9 10 0 9 1 15 1 9 2 13 3 7 1 9 9 13 9 2
11 9 13 2 15 0 2 9 1 0 9 2
27 0 9 1 9 13 1 9 7 3 15 3 13 3 2 13 13 1 9 9 7 13 3 10 9 1 9 2
17 9 3 3 13 3 2 3 13 2 16 13 9 2 10 0 9 2
6 13 3 9 7 9 2
30 16 3 1 9 13 1 10 9 1 9 9 1 0 9 7 3 13 9 10 2 13 4 15 1 9 1 0 9 9 2
18 15 15 10 0 9 3 3 13 2 16 1 9 15 1 9 13 9 2
15 13 15 2 16 0 9 1 15 13 0 9 2 0 9 2
4 13 15 3 2
20 7 15 4 1 15 13 2 16 15 1 9 1 9 13 2 2 2 7 13 2
9 16 13 9 2 0 13 10 9 2
9 7 1 10 9 13 1 9 9 2
35 16 13 1 9 2 15 13 1 9 2 7 1 9 13 9 2 3 15 13 2 13 3 0 2 16 3 13 2 16 4 15 0 9 13 2
3 3 9 2
13 3 2 16 11 13 11 2 15 15 3 13 13 2
37 1 9 9 13 13 9 9 1 9 9 2 15 1 12 9 3 9 13 9 9 13 2 1 9 0 15 1 9 4 13 2 16 4 13 0 9 2
13 13 2 3 13 10 9 2 9 13 13 10 9 2
4 7 0 9 2
28 13 15 2 16 13 3 9 9 2 3 15 15 13 15 2 15 9 1 0 9 13 0 9 7 15 10 9 2
28 7 15 1 15 13 13 2 16 13 3 0 9 2 16 1 15 13 9 7 1 9 13 9 2 3 15 13 2
9 3 3 13 2 16 4 15 13 2
4 0 9 1 9
2 11 2
18 0 9 0 0 9 1 9 11 15 13 1 9 1 0 9 0 9 2
12 1 15 13 0 9 9 0 9 1 9 11 2
43 1 9 2 15 4 3 13 1 9 11 7 1 0 9 11 2 15 13 2 16 10 9 13 1 9 0 2 0 9 7 1 9 9 7 9 2 16 4 11 13 1 9 2
34 1 9 0 9 15 9 2 15 1 0 9 1 11 1 0 9 9 13 9 7 12 0 13 2 13 1 9 3 1 9 1 9 11 2
29 9 9 11 11 11 2 15 13 1 11 2 7 1 9 1 0 9 13 2 16 0 9 1 0 9 11 9 13 2
4 9 1 9 13
2 11 2
23 1 0 0 9 3 13 1 11 0 9 11 1 9 7 9 2 15 13 1 12 2 9 2
9 9 15 13 1 12 9 0 9 2
11 9 11 13 9 0 9 9 9 11 11 2
16 3 1 9 13 9 0 9 2 15 15 1 11 13 1 12 2
7 9 9 13 1 12 9 2
38 9 13 10 0 9 11 11 7 3 13 0 9 10 9 2 0 9 11 11 2 15 13 2 16 9 13 9 1 0 9 7 9 2 15 13 0 13 2
31 0 9 11 11 11 2 11 13 9 1 0 9 1 15 0 9 7 13 2 14 15 9 13 0 9 2 13 0 9 3 2
28 0 9 11 11 1 10 9 13 2 16 11 4 1 9 13 1 15 2 16 4 15 1 9 13 9 9 9 2
18 0 9 11 11 13 9 2 16 4 13 9 2 15 13 13 0 9 2
10 9 13 9 2 13 9 9 2 13 2
26 9 13 9 0 9 11 11 11 2 1 15 15 13 1 9 9 9 1 9 16 9 1 9 9 9 2
4 3 1 9 12
7 1 9 11 2 12 15 13
7 11 2 11 2 11 2 2
24 0 9 0 9 11 2 12 2 16 1 0 9 2 13 4 1 9 9 13 1 9 1 11 2
30 1 0 9 4 13 3 0 13 0 9 0 2 7 0 12 9 11 2 12 16 13 1 9 12 9 0 11 2 12 2
39 9 0 9 11 11 15 7 13 2 16 9 0 9 11 2 12 13 3 0 2 3 1 15 9 13 2 1 9 1 11 2 12 2 9 0 9 7 9 2
19 1 9 13 14 0 13 7 0 0 9 1 11 2 15 11 2 12 13 2
27 11 2 12 4 1 9 13 13 0 9 0 9 11 2 12 7 1 10 9 7 3 0 9 11 2 12 2
19 11 13 2 16 1 9 2 1 15 13 9 7 0 9 2 13 3 13 2
6 0 9 1 11 13 0
2 11 2
9 11 3 3 13 10 9 1 11 2
11 3 3 3 13 1 9 9 13 10 9 2
11 13 15 3 11 11 1 0 9 0 9 2
13 13 3 2 16 0 9 3 13 7 9 13 9 2
31 11 13 1 0 9 1 9 2 3 11 11 12 2 13 2 13 2 16 13 1 11 2 4 2 14 13 9 0 0 9 2
26 3 13 9 2 13 11 2 15 13 11 11 2 11 2 15 13 1 9 11 1 9 7 9 1 11 2
5 0 9 1 12 9
14 0 0 9 13 1 12 9 1 9 11 1 9 10 9
2 11 11
2 11 2
30 0 9 0 0 9 2 0 2 9 2 11 2 12 2 12 2 12 13 1 10 15 0 9 1 9 10 9 11 11 2
33 14 2 13 4 0 9 2 13 3 1 11 11 2 11 1 9 12 9 0 2 9 2 11 1 9 11 1 0 9 12 9 9 2
10 10 0 9 15 13 1 12 9 9 2
21 1 11 13 1 0 9 9 0 9 0 9 1 0 9 1 9 9 9 7 11 2
12 9 9 13 3 0 0 9 11 2 0 9 2
25 0 9 1 10 9 13 0 9 11 11 11 7 0 9 0 2 9 2 11 2 3 9 11 11 2
35 15 15 3 1 9 12 13 9 0 9 1 9 0 2 9 2 11 2 7 9 12 9 9 2 15 1 9 13 2 1 0 9 3 13 2
7 1 11 13 7 0 9 2
26 1 9 12 12 9 0 2 9 2 11 2 15 9 13 1 12 0 9 2 13 1 9 1 0 9 2
18 0 9 1 11 7 0 2 9 2 11 13 13 0 9 1 15 0 2
40 7 9 3 2 16 11 13 0 9 1 9 0 2 9 2 11 2 13 9 10 9 11 2 11 9 1 0 9 2 1 15 11 13 2 2 15 0 9 13 2
8 10 9 13 3 11 1 11 2
8 15 11 1 10 0 9 13 2
18 9 3 13 0 2 9 2 11 2 7 12 9 3 10 9 13 11 2
9 15 0 9 13 1 9 3 13 2
24 16 0 2 9 2 11 10 9 13 13 2 11 13 0 9 1 11 2 16 4 9 13 13 2
15 3 11 9 13 0 9 11 2 0 9 1 12 9 9 2
16 15 1 9 9 0 2 9 2 11 11 2 11 7 9 9 2
34 9 10 9 9 13 9 1 9 1 0 9 2 15 3 13 9 9 0 9 1 9 9 2 7 13 13 10 0 9 2 13 9 11 2
3 13 13 2
17 9 15 7 3 13 2 13 3 0 9 9 9 9 9 11 11 2
13 9 0 9 13 9 2 1 11 4 13 1 9 2
8 9 11 14 13 9 1 9 11
5 11 2 11 2 2
41 0 9 1 9 9 9 9 11 2 11 9 9 0 11 11 11 2 2 16 4 1 9 9 1 9 9 2 12 13 0 9 11 2 13 0 9 1 11 7 11 2
8 11 15 13 9 0 0 9 2
21 11 11 13 9 0 11 9 9 2 12 2 13 13 9 0 9 11 2 1 11 2
15 11 13 3 0 9 2 7 1 9 0 9 15 13 9 2
45 1 9 11 13 0 9 9 9 2 15 13 9 9 1 9 9 1 9 2 12 2 9 9 11 2 11 9 9 11 2 11 7 9 11 11 2 11 2 16 4 13 0 9 9 2
6 15 9 13 1 0 2
12 11 2 15 13 0 9 2 15 9 3 13 2
18 9 13 2 16 13 9 2 12 1 9 9 9 13 2 15 11 13 2
13 13 2 16 13 9 1 9 11 1 9 2 12 2
35 1 9 9 13 1 9 11 3 1 0 9 2 15 15 1 0 9 1 0 9 9 11 1 9 11 1 0 9 13 9 1 11 1 9 2
3 9 1 9
2 11 11
10 9 9 9 13 3 3 0 0 9 2
10 13 0 9 2 15 4 13 1 9 2
2 3 2
20 1 0 9 0 9 2 1 10 9 3 14 3 0 2 7 9 0 11 13 2
19 1 0 9 2 15 15 13 1 9 1 9 0 2 4 10 9 3 13 2
21 7 9 7 0 9 15 1 15 9 9 0 9 13 3 1 0 9 0 9 9 2
11 13 9 7 0 9 15 13 13 1 9 2
9 9 1 0 9 4 13 1 9 2
4 9 3 13 2
29 3 0 9 1 9 9 13 3 2 13 15 2 9 3 2 7 16 3 15 4 3 1 9 13 3 7 3 13 2
8 9 13 7 9 0 7 0 2
23 13 2 14 15 2 4 13 1 0 9 9 2 15 13 2 1 9 9 2 3 1 9 2
7 9 1 9 9 3 13 2
14 13 15 9 0 2 16 0 9 15 1 9 13 3 2
9 9 3 0 2 0 2 16 0 2
20 13 1 15 7 7 0 9 0 2 0 1 15 2 16 1 9 13 0 9 2
7 0 9 13 11 2 11 2
17 13 0 9 9 1 15 2 16 1 0 0 9 4 3 13 9 2
23 14 9 13 3 0 0 9 1 9 1 9 2 15 10 9 2 1 15 0 2 3 13 2
13 13 15 7 2 16 4 0 9 13 0 9 13 2
11 13 1 15 2 16 13 1 9 0 9 2
11 9 13 3 0 2 3 3 0 1 9 2
14 13 15 2 16 13 1 9 13 13 9 1 9 9 2
10 13 15 2 16 9 9 9 3 13 2
12 13 2 1 15 4 3 0 9 13 0 9 2
9 0 9 13 0 1 10 9 0 2
17 1 0 9 9 1 9 0 9 13 9 2 16 13 0 16 9 2
7 9 9 9 4 13 13 2
23 13 2 14 15 9 9 3 7 3 2 14 13 1 9 2 15 4 13 1 10 0 9 2
8 0 9 1 9 13 9 0 2
5 13 7 3 0 2
5 16 0 2 13 2
17 13 7 0 9 16 0 9 1 15 2 15 4 3 13 9 9 2
6 0 0 9 13 1 11
3 1 0 9
2 11 2
20 0 9 9 9 9 11 11 11 13 1 11 1 9 1 9 9 11 11 11 2
17 1 9 9 11 13 1 15 3 0 9 9 7 0 0 9 11 2
17 11 0 9 13 2 16 4 13 1 0 9 9 11 11 2 11 2
34 13 9 2 13 3 11 2 16 9 9 13 9 13 1 0 9 9 2 7 3 13 2 16 13 9 1 0 9 13 9 1 15 9 2
16 0 9 15 11 13 13 1 9 9 7 1 11 2 7 3 2
4 9 13 3 9
2 11 2
9 0 9 0 9 7 9 13 9 2
25 9 9 1 12 9 9 13 1 0 9 12 7 3 2 16 0 9 13 3 12 9 1 12 9 2
9 13 15 9 9 11 11 11 11 2
15 11 13 9 7 0 9 9 1 9 2 9 7 0 9 2
23 9 9 13 2 16 13 13 9 9 1 12 9 2 16 9 0 9 1 12 2 12 9 2
22 1 12 2 9 0 9 9 13 12 9 0 9 9 2 15 13 14 12 9 9 3 2
15 1 9 11 13 1 9 1 0 0 9 3 0 0 9 2
26 16 4 0 9 13 7 3 2 13 4 1 0 9 1 0 0 9 13 0 16 1 15 1 0 9 2
16 15 13 3 1 9 0 0 9 2 3 9 2 13 11 11 2
19 0 9 13 12 1 9 2 3 9 1 0 0 9 13 3 13 0 9 2
32 0 0 9 1 11 13 3 12 9 9 2 7 7 13 9 9 13 3 3 0 9 2 16 13 0 15 9 0 9 3 13 2
5 11 13 9 0 9
2 11 2
16 11 13 13 0 9 9 1 9 0 0 9 7 10 0 9 2
11 3 15 13 9 9 1 10 9 11 11 2
14 0 9 9 2 15 13 12 0 9 2 13 1 0 2
22 1 11 4 11 13 9 1 9 0 9 11 2 12 9 2 7 11 2 12 9 2 2
27 11 13 1 9 1 9 1 15 2 16 9 1 9 0 0 9 4 15 13 13 3 1 9 1 10 9 2
17 11 13 2 16 11 13 0 13 9 3 3 1 0 9 10 9 2
30 9 11 13 15 1 10 2 16 4 4 9 13 10 9 2 15 13 13 2 7 13 15 3 15 13 1 9 2 13 2
10 11 2 11 13 2 16 9 13 9 11
5 11 2 11 2 2
20 0 0 2 9 2 13 9 0 0 9 10 9 7 13 0 9 1 10 9 2
20 10 9 13 9 11 11 11 1 0 9 9 1 9 10 9 1 0 9 9 2
28 3 11 13 9 9 9 11 2 4 2 14 1 10 9 13 9 7 9 2 13 9 2 15 4 9 11 13 2
28 9 11 0 9 13 2 16 7 9 2 15 4 1 9 9 13 3 3 2 4 13 9 10 9 1 0 9 2
9 13 15 15 14 3 9 1 11 2
20 1 0 9 15 11 13 3 13 1 9 0 9 2 15 15 13 9 9 13 2
11 13 0 9 2 16 13 9 2 13 0 2
18 16 4 15 10 9 13 2 13 4 15 13 13 9 1 11 2 13 2
19 1 0 9 1 9 11 15 4 0 9 13 3 1 9 7 9 1 11 2
13 9 7 9 13 2 16 9 12 13 13 9 1 11
9 11 2 11 2 11 2 11 2 2
24 9 12 13 1 3 0 9 1 9 9 1 0 9 9 0 9 0 9 11 11 2 11 2 2
22 13 3 1 9 9 11 11 2 1 15 3 1 0 9 13 9 1 0 9 0 9 2
8 3 4 15 13 2 13 11 2
44 3 1 9 7 11 13 2 16 1 9 9 13 0 13 1 0 9 7 16 13 0 13 1 0 9 12 2 7 15 0 0 9 13 1 0 0 9 11 0 1 9 1 11 2
24 3 9 0 9 11 11 2 11 2 13 2 16 9 9 1 9 12 13 3 3 1 0 9 2
12 13 7 2 16 1 9 9 9 3 3 13 2
8 1 11 13 3 1 9 11 2
28 9 0 9 11 11 2 11 2 13 2 16 11 0 9 12 13 1 15 0 9 7 16 3 0 9 3 13 2
17 13 15 9 0 2 16 4 15 3 13 7 16 4 13 2 13 2
5 0 9 1 0 9
7 11 2 11 2 11 2 2
37 1 0 13 1 0 9 1 9 11 11 9 0 0 2 0 9 0 9 0 0 0 0 9 11 11 2 11 2 15 13 1 10 9 1 9 11 2
23 1 11 13 1 9 0 9 13 10 0 9 1 11 2 1 15 15 4 13 9 10 9 2
30 4 13 0 9 1 11 2 7 4 13 0 9 2 13 3 1 9 1 0 9 9 0 9 9 11 11 2 11 2 2
11 9 0 9 1 11 11 13 16 0 9 2
19 1 9 14 9 9 0 9 13 2 7 0 9 1 11 10 9 13 3 2
33 1 9 12 9 13 0 9 2 15 11 13 15 2 16 13 3 0 13 10 9 2 3 3 13 7 0 1 15 13 0 9 11 2
23 9 11 2 11 3 13 1 9 0 0 9 11 11 2 11 1 0 9 9 0 2 0 9
5 9 11 11 2 11
8 11 2 11 1 9 9 1 9
5 11 2 11 2 2
36 13 2 3 11 13 9 9 1 9 2 13 1 9 9 9 11 2 11 12 1 9 10 0 9 1 9 9 0 9 2 11 2 11 2 11 2
20 11 3 2 13 9 2 16 4 15 0 9 13 1 0 9 11 1 0 9 2
14 11 13 7 1 9 9 11 2 11 7 9 9 9 2
5 0 9 7 9 9
9 1 10 9 13 0 9 1 9 9
7 11 2 11 2 11 2 2
17 9 0 9 13 1 0 2 16 4 9 0 9 0 9 13 9 2
19 13 1 15 7 0 9 9 1 9 0 9 2 15 13 9 13 10 9 2
38 9 0 9 11 11 2 11 2 11 13 2 16 13 0 13 10 9 9 0 9 2 1 15 13 3 9 2 1 9 0 2 3 1 0 9 13 9 2
20 10 9 13 9 3 1 0 9 2 16 1 11 9 9 13 1 0 9 3 2
30 13 2 14 3 10 9 9 3 13 1 9 2 15 15 9 13 1 0 9 2 13 1 11 13 15 7 1 9 9 2
14 9 13 3 13 3 9 0 0 9 7 0 9 9 2
26 1 9 2 16 4 9 0 9 1 10 9 13 9 9 0 9 1 9 9 2 11 13 2 16 3 2
16 13 2 16 13 9 3 0 2 16 4 13 0 10 9 13 2
11 1 10 9 15 1 15 0 9 13 3 2
13 1 9 0 9 9 13 2 16 15 13 14 3 2
7 7 1 15 13 0 9 2
14 11 14 3 13 2 16 9 15 1 10 9 3 13 2
19 3 15 13 13 9 10 9 2 16 16 4 1 15 13 0 9 2 13 2
23 13 2 16 13 9 9 2 16 4 13 10 9 1 10 9 2 15 13 9 0 0 9 2
31 9 9 11 11 2 11 2 13 1 0 2 16 9 13 9 0 9 9 9 0 9 0 0 9 2 1 15 10 9 13 2
14 1 9 9 11 11 11 13 2 16 4 9 13 9 2
12 1 11 4 13 9 9 13 7 0 0 9 2
13 13 15 13 2 16 4 15 13 9 9 2 13 2
22 11 15 13 2 16 0 9 4 1 9 9 0 9 13 1 9 13 7 0 0 9 2
5 4 0 9 13 2
5 11 2 11 2 2
17 0 0 9 11 11 13 13 1 0 9 9 0 9 1 11 12 2
18 13 15 1 9 2 15 11 13 9 0 9 1 11 12 11 2 11 2
19 1 15 13 0 9 0 9 0 2 7 11 7 13 13 1 10 0 9 2
22 15 7 13 2 16 15 9 11 1 9 11 1 11 12 1 10 9 13 2 13 11 2
5 0 9 13 13 9
23 9 10 9 1 9 1 9 13 9 3 2 16 15 0 9 13 0 9 13 3 0 9 2
30 9 7 9 0 9 7 3 1 0 9 13 9 0 9 10 9 13 1 9 1 0 0 9 1 10 9 1 0 9 2
10 3 3 15 3 13 13 9 0 9 2
32 3 1 9 12 0 9 7 12 9 9 1 9 0 0 9 13 9 0 0 9 2 16 1 12 9 13 9 9 1 0 9 2
9 10 9 13 0 3 1 0 9 2
19 0 9 2 15 13 0 9 7 9 1 10 9 2 0 9 0 9 13 2
19 9 13 9 1 9 1 0 9 13 12 9 2 15 13 12 9 0 9 2
27 1 0 9 1 9 3 16 9 9 2 15 13 9 9 1 0 9 2 13 9 9 0 9 1 9 9 2
12 9 0 9 1 0 9 13 1 10 9 0 2
19 10 9 13 1 9 2 0 9 7 3 7 1 15 2 16 9 13 0 2
17 15 7 3 13 2 16 13 13 3 0 2 0 9 7 9 9 2
9 7 13 9 1 9 3 0 9 2
28 16 15 13 9 13 9 1 9 7 13 13 9 2 16 9 15 1 9 13 2 13 15 0 9 13 1 9 2
23 9 13 3 0 15 13 2 7 15 3 1 9 2 15 9 4 13 13 0 9 7 9 2
3 2 11 2
5 0 9 1 9 11
3 1 0 9
5 11 2 11 2 2
16 1 0 9 1 0 9 13 11 1 0 11 0 9 1 11 2
12 9 11 15 13 7 0 0 9 9 11 11 2
10 13 15 3 9 0 9 11 11 11 2
17 0 9 4 1 12 9 0 1 9 0 9 13 1 9 12 9 2
14 1 11 4 11 13 1 0 0 9 3 1 9 0 2
3 13 7 9
6 0 11 2 11 2 2
28 16 9 9 9 13 9 2 13 1 10 9 0 9 7 13 12 9 2 9 7 9 1 12 9 7 0 9 2
3 9 9 9
5 11 2 11 2 2
27 0 9 13 1 9 1 9 1 9 0 11 2 11 2 1 9 9 1 0 9 10 1 12 9 0 9 2
8 11 15 13 9 0 9 9 2
13 9 9 2 15 9 15 13 2 13 0 0 9 2
29 0 9 2 15 15 1 9 9 3 1 9 13 2 13 11 2 11 2 2 0 1 9 0 9 2 1 9 9 2
17 9 2 15 15 0 0 9 0 9 13 15 2 4 13 1 9 2
23 9 1 0 9 9 4 13 3 2 16 13 11 2 11 2 0 9 1 0 9 7 9 2
4 0 13 1 9
5 11 2 11 2 2
23 16 3 13 0 9 2 13 1 0 12 0 9 12 0 9 1 9 1 1 9 1 9 2
9 13 1 9 2 1 15 12 13 2
4 15 9 13 2
5 3 13 0 9 2
30 15 15 12 1 9 13 3 3 2 16 13 9 2 9 1 9 7 9 15 13 0 9 2 13 11 0 9 11 11 2
16 0 15 13 9 1 9 2 7 9 13 4 1 10 9 13 2
4 1 9 13 9
5 11 2 11 2 2
33 9 13 1 0 9 9 0 9 11 2 11 2 7 1 9 13 12 9 1 9 12 9 9 2 15 13 9 11 11 1 11 13 2
16 9 15 13 1 9 13 3 1 0 0 9 1 0 0 9 2
11 1 12 9 0 9 13 1 9 0 9 2
26 13 9 9 2 15 15 13 1 10 9 2 1 9 1 9 2 13 9 11 2 11 1 0 9 9 2
16 9 15 13 2 16 10 9 13 9 1 9 1 0 0 9 2
3 0 11 13
5 11 2 11 2 2
30 0 11 11 2 15 12 2 12 2 1 11 9 13 12 9 0 9 1 9 2 3 13 1 0 9 1 11 2 11 2
13 11 15 13 9 0 9 9 2 15 15 9 13 2
20 16 3 4 1 11 13 2 11 2 11 13 9 1 9 7 13 1 9 9 2
15 3 1 9 1 9 9 13 12 9 2 15 11 3 13 2
21 1 0 0 9 13 3 0 12 0 9 1 11 2 0 11 11 7 0 11 11 2
7 1 12 9 9 3 13 2
5 3 1 9 0 11
10 1 0 9 4 13 1 9 9 0 9
2 11 2
19 0 0 9 1 9 1 0 9 0 0 0 9 0 11 13 0 0 9 2
14 1 0 9 4 13 1 12 7 12 9 3 16 3 2
8 3 0 9 13 1 12 3 2
9 3 9 1 9 13 1 9 9 2
14 0 9 13 1 9 9 0 9 7 13 10 0 9 2
42 1 0 0 9 4 13 0 9 1 11 2 9 1 12 9 2 2 2 15 13 1 0 9 1 11 2 11 2 11 2 11 2 11 1 11 2 11 1 11 7 11 2
35 0 0 9 2 9 1 12 9 2 2 1 0 11 13 1 11 1 11 2 11 2 11 1 11 2 11 2 11 2 11 7 11 1 11 2
32 1 0 9 4 13 0 0 9 11 2 11 2 9 1 12 9 2 2 7 11 2 11 2 11 2 9 1 12 9 2 2 2
54 1 0 9 9 13 0 9 12 2 9 1 12 9 2 1 11 2 11 0 9 1 11 2 11 2 11 2 11 1 11 2 0 11 2 11 1 11 2 11 2 11 1 11 2 11 2 11 2 11 2 11 7 11 2
40 0 0 9 13 1 12 9 2 1 0 0 9 9 1 11 2 11 11 2 11 2 0 11 2 11 1 11 2 11 7 11 2 3 9 0 9 1 11 2 2
14 0 0 9 11 2 11 13 1 0 9 1 12 9 2
41 1 10 9 4 1 12 9 2 13 0 9 1 0 11 2 0 1 11 2 11 2 11 1 11 2 11 2 11 2 11 2 11 1 11 7 11 1 11 2 11 2
14 1 11 2 11 1 11 13 0 0 9 1 12 9 2
15 0 9 1 11 13 1 0 0 9 1 12 2 12 9 2
43 13 1 11 2 11 2 11 1 11 2 11 1 11 2 11 1 11 2 11 2 11 2 11 1 11 2 11 1 11 2 11 2 11 1 11 7 0 9 1 11 1 11 2
23 1 0 11 13 1 0 0 9 1 12 9 2 1 11 2 11 2 11 7 11 0 9 2
22 1 12 9 2 13 1 11 0 9 1 9 1 11 2 11 1 11 7 11 1 11 2
9 9 2 15 13 1 9 2 1 9
2 0 9
5 11 2 11 2 2
31 1 0 9 9 2 9 0 9 2 9 7 0 9 0 9 13 3 1 0 9 1 11 0 11 11 2 1 11 1 11 2
16 4 13 1 15 2 16 13 1 9 0 11 11 2 1 11 2
9 13 15 9 1 9 1 12 9 2
9 1 9 9 15 7 13 3 3 2
8 11 11 2 3 13 3 9 2
16 9 2 15 15 13 1 9 7 9 2 0 1 10 9 13 2
14 0 15 3 1 9 13 3 9 1 10 11 7 13 2
8 1 9 0 1 9 9 13 2
17 13 15 3 14 13 10 9 2 15 15 1 11 11 2 3 13 2
6 15 3 15 7 13 2
25 1 9 1 0 9 11 11 2 1 9 3 13 9 2 16 15 9 9 13 2 13 7 3 13 2
6 7 1 15 13 9 2
9 3 15 1 15 13 14 1 9 2
18 0 9 13 9 9 9 1 9 1 12 1 12 9 2 3 7 0 2
7 3 13 0 9 9 9 2
19 1 0 9 0 1 0 9 15 13 0 0 9 16 1 9 0 1 9 2
14 9 3 1 10 9 3 13 1 9 7 9 0 9 2
3 9 11 11
1 9
29 3 1 9 9 13 1 9 1 12 9 1 0 11 9 1 11 2 11 2 2 12 2 7 1 12 9 0 9 2
15 9 15 3 13 7 9 13 9 1 0 11 2 3 13 2
13 9 4 13 1 0 9 9 1 9 1 9 9 2
15 0 9 0 15 1 0 9 13 1 9 3 0 9 9 2
12 9 1 9 9 11 11 2 11 13 12 9 2
3 2 11 2
15 3 13 9 1 0 9 1 9 11 1 9 11 1 11 2
11 1 9 13 9 0 9 12 0 9 9 2
12 1 9 1 9 4 13 1 0 9 1 11 2
3 2 11 2
1 9
1 9
2 11 11
14 0 9 0 9 11 13 9 9 0 9 13 9 9 2
17 1 13 2 16 15 13 2 7 10 9 9 2 1 15 9 13 2
18 3 4 15 7 15 2 15 13 3 1 9 2 13 13 9 0 2 2
15 9 13 2 9 13 3 2 13 0 9 3 0 0 9 2
21 1 0 9 13 15 14 0 9 2 13 9 9 11 2 3 13 1 9 0 9 2
9 3 1 10 9 0 9 2 2 2
13 15 13 9 13 2 15 13 9 2 13 10 9 2
29 3 13 15 3 0 9 10 9 11 1 15 9 2 1 9 2 1 0 9 2 15 13 0 9 0 9 10 9 2
8 13 12 9 7 9 3 13 2
31 11 16 4 13 13 2 15 10 9 0 9 3 10 9 13 2 16 3 15 15 13 3 10 0 9 2 15 15 13 13 2
15 13 4 14 0 2 16 4 0 9 13 3 0 0 9 2
26 14 3 1 15 15 2 16 1 0 7 0 9 2 15 13 9 7 15 10 9 3 13 3 1 9 2
32 13 2 14 4 10 9 13 3 3 2 16 15 10 9 13 1 9 7 3 13 9 9 0 9 2 13 13 9 0 0 9 2
11 1 0 9 11 15 3 13 1 9 9 11
5 9 11 11 2 11
4 9 14 1 9
1 9
2 11 11
15 9 9 9 1 9 1 9 3 13 0 9 1 0 9 2
21 3 16 1 9 15 15 3 13 1 15 2 3 0 7 3 0 13 13 0 9 2
21 3 13 13 2 16 15 9 3 13 1 9 0 2 3 1 0 9 10 0 9 2
17 15 0 4 13 4 13 1 0 9 2 3 0 0 9 7 9 2
17 0 9 1 9 0 9 4 15 7 10 0 9 13 3 3 13 2
27 1 9 11 13 3 0 2 16 9 1 9 3 2 13 2 10 0 9 9 13 0 9 1 9 1 9 2
11 7 9 0 9 7 13 10 9 1 9 2
21 9 12 0 0 9 13 2 16 13 10 9 13 7 13 15 2 15 13 1 9 2
18 1 9 9 10 9 11 11 13 7 15 9 7 9 9 7 9 0 2
46 13 2 14 15 3 2 13 3 1 9 2 16 10 9 13 3 3 13 9 1 15 2 16 13 3 2 10 10 9 0 13 9 1 9 9 1 0 2 3 1 9 3 15 15 13 2
26 3 4 1 9 0 9 1 10 9 0 9 1 9 13 2 16 9 9 1 9 13 14 1 10 9 2
14 9 1 0 9 7 3 0 9 9 13 7 13 9 2
29 1 9 1 9 1 0 9 13 9 3 13 2 1 0 9 4 14 7 13 13 0 9 9 9 13 9 1 15 2
14 15 15 13 3 1 9 2 15 15 13 0 9 9 2
3 9 0 9
2 11 11
14 0 9 0 9 13 10 9 13 0 9 1 0 9 2
12 9 1 15 13 3 1 9 0 9 0 11 2
28 0 7 0 9 2 15 13 1 9 9 12 0 9 2 3 1 12 9 13 3 16 0 9 1 11 11 11 2
21 13 15 7 2 16 9 0 9 0 9 1 0 9 3 13 9 0 3 0 9 2
16 9 0 9 3 13 13 0 9 0 0 9 1 0 0 9 2
7 1 11 3 13 12 9 2
11 3 12 1 15 7 13 3 1 9 12 2
6 0 13 1 0 9 2
24 1 9 2 1 0 9 2 1 0 9 7 3 1 9 2 15 4 15 13 3 0 0 9 2
28 16 4 0 0 9 3 13 13 2 4 13 13 3 0 0 9 1 9 7 13 1 9 9 1 9 0 9 2
12 9 9 1 0 7 0 9 15 7 3 13 2
23 1 0 0 9 2 1 15 13 13 0 9 15 0 9 2 3 13 3 0 9 0 9 2
6 9 0 9 7 13 2
16 3 3 0 9 1 9 13 10 0 9 13 7 3 0 9 2
35 13 2 14 1 9 0 9 2 16 1 0 0 9 13 1 9 9 0 13 3 0 9 2 13 1 9 2 16 0 9 13 15 0 9 2
11 0 9 15 3 3 13 0 16 0 9 2
12 16 4 13 9 13 0 9 2 13 0 9 2
29 7 3 15 13 3 1 9 9 7 1 0 0 9 9 9 2 15 1 9 9 13 7 0 9 0 0 0 9 2
13 7 15 13 13 9 1 0 9 1 0 0 9 2
48 13 2 14 4 1 0 0 9 13 9 2 15 13 0 1 9 7 9 2 7 7 0 9 2 13 0 2 16 4 13 9 0 9 2 15 4 13 9 0 9 7 13 3 10 0 0 9 2
21 0 9 10 9 4 7 3 13 13 9 0 9 2 7 15 3 1 9 0 9 2
20 13 1 0 9 0 9 7 0 7 0 9 13 3 3 1 9 0 9 0 2
20 10 9 2 15 13 9 0 0 9 3 13 2 13 7 1 0 9 3 0 2
16 1 0 9 2 15 13 3 1 9 12 2 14 13 0 9 2
17 16 12 0 9 2 15 15 13 2 3 10 9 1 0 9 13 2
14 3 16 12 1 15 13 0 2 16 13 3 0 9 2
3 11 1 9
2 11 11
9 0 0 9 3 13 0 0 9 2
23 10 0 9 13 7 3 1 9 15 2 16 13 3 9 1 9 0 0 0 9 16 15 2
10 0 9 13 9 1 0 0 0 9 2
19 1 0 0 9 13 0 9 10 0 9 2 15 3 1 9 13 1 9 2
21 1 0 0 9 3 13 9 1 9 16 0 0 9 7 0 9 4 13 1 9 2
11 1 0 0 9 13 10 9 3 0 9 2
17 9 0 0 9 3 13 13 9 2 10 9 13 1 9 11 11 2
12 13 9 2 16 9 13 9 0 9 1 11 2
28 3 0 0 9 4 13 13 3 9 1 9 9 7 10 9 2 15 13 3 7 1 3 0 9 15 1 9 2
13 3 7 7 13 3 9 1 9 0 9 3 0 2
12 3 0 9 11 13 0 9 9 7 9 9 2
13 1 9 13 12 0 9 2 1 15 13 0 9 2
32 3 13 15 0 9 2 0 1 9 9 7 9 11 2 3 0 9 7 3 0 9 2 0 1 9 2 15 13 0 9 9 2
14 0 9 1 9 10 0 9 13 3 13 9 0 9 2
29 7 11 11 13 9 3 16 9 1 9 10 0 9 2 7 7 13 15 3 13 1 9 0 9 7 1 0 9 2
20 7 3 9 9 2 15 13 13 0 9 1 9 9 2 13 1 11 3 13 2
27 1 10 0 9 13 3 9 11 2 15 13 2 1 10 9 3 13 7 13 2 0 9 1 9 0 9 2
19 0 9 0 9 9 13 9 2 16 3 13 2 9 11 11 2 1 9 2
19 3 13 2 9 15 13 2 14 16 13 2 7 4 0 9 13 1 9 2
14 0 9 0 9 7 13 0 9 11 2 1 9 9 2
12 1 9 4 10 9 13 16 9 11 1 11 2
19 13 7 1 0 0 9 2 7 1 9 2 1 15 15 13 0 0 9 2
17 9 13 3 1 9 1 0 9 2 3 9 9 13 13 9 11 2
15 1 12 2 9 3 13 1 9 1 9 0 7 0 9 2
13 15 0 13 13 10 9 0 9 11 1 9 12 2
19 0 9 4 3 13 13 9 1 9 1 9 2 15 13 3 9 9 11 2
33 9 15 0 3 13 7 16 3 2 13 0 9 2 13 3 10 9 1 9 13 1 0 9 2 9 2 9 2 9 1 11 2 2
14 9 13 2 3 3 3 13 9 0 9 1 9 0 2
18 0 9 1 12 9 3 13 1 0 1 0 9 0 9 1 0 9 2
15 3 3 7 15 1 0 0 9 3 13 1 9 9 11 2
8 1 0 0 9 3 3 13 2
24 16 15 0 0 9 3 13 0 7 10 9 13 9 1 0 0 9 1 9 2 13 3 13 2
4 3 9 7 9
1 9
2 11 11
19 13 13 2 16 9 2 3 0 9 2 13 0 9 9 16 15 0 9 2
16 9 9 15 3 3 13 7 9 0 2 10 13 3 0 9 2
18 9 13 0 9 2 13 0 9 2 13 9 7 13 15 13 0 9 2
24 1 9 9 15 3 3 13 9 2 16 1 0 9 15 9 3 13 1 0 9 0 0 9 2
25 16 4 13 9 10 9 7 15 15 13 13 1 9 9 2 13 4 15 3 1 9 10 0 9 2
10 13 2 14 0 9 2 13 7 0 2
15 13 3 2 16 0 9 0 9 1 0 9 13 0 9 2
29 9 16 0 9 7 0 0 9 2 3 11 7 11 2 13 9 0 0 9 7 9 13 3 3 10 3 0 9 2
33 9 2 0 1 0 9 9 0 9 2 13 3 15 9 7 13 2 10 9 13 3 3 0 1 10 9 2 15 13 9 7 9 2
29 1 9 13 9 3 0 16 9 2 16 13 2 16 4 1 0 9 9 13 1 15 2 16 13 2 15 15 13 2
34 12 2 9 13 11 3 9 2 16 0 9 13 3 12 9 10 9 9 2 1 15 13 13 10 9 14 1 9 12 9 1 0 9 2
9 9 13 0 9 2 7 13 0 2
22 11 15 13 14 15 2 16 9 13 13 2 15 3 13 2 15 13 9 3 0 9 2
25 13 4 10 9 13 2 16 0 9 13 3 9 0 0 9 2 15 9 0 9 1 9 0 13 2
20 7 15 9 13 2 7 9 15 2 3 7 9 2 15 15 14 13 3 13 2
23 13 15 2 16 4 3 3 1 9 13 10 9 2 16 9 13 0 2 7 10 9 13 2
25 15 15 13 1 15 0 2 14 3 2 16 15 9 13 2 7 3 2 16 15 13 1 9 9 2
42 13 4 12 2 12 2 9 1 15 2 16 3 1 0 9 11 3 13 9 0 9 2 10 0 9 3 13 0 0 9 2 13 2 14 15 0 9 3 13 0 9 2
16 13 0 2 16 15 10 0 9 13 7 16 1 10 9 13 2
42 0 13 7 15 2 13 15 3 13 13 1 15 2 16 0 9 13 0 2 3 7 3 0 0 9 2 3 15 0 1 0 9 2 1 15 10 9 13 13 0 9 2
20 13 15 2 16 4 9 2 15 15 13 2 3 13 2 16 15 1 9 13 2
22 13 4 15 7 13 9 9 1 15 15 13 13 15 2 1 15 1 11 13 15 3 2
12 13 15 0 9 2 15 13 3 0 9 9 2
32 13 13 2 16 4 13 13 3 0 9 2 16 4 9 1 15 2 16 10 0 9 13 0 9 2 13 1 9 9 0 11 2
6 3 3 13 3 1 0
10 1 9 1 0 9 13 3 14 12 9
7 0 9 11 1 11 11 11
17 12 9 3 13 0 9 1 9 1 0 9 2 12 2 9 2 2
7 0 9 13 1 0 9 2
41 9 11 13 1 0 9 9 10 9 2 11 2 11 2 7 9 0 9 1 9 9 11 11 13 2 3 16 0 9 10 9 4 3 13 2 9 3 10 0 9 2
34 11 15 13 13 1 10 9 2 7 9 2 3 9 0 9 9 13 9 2 0 9 10 9 2 7 15 7 0 9 7 9 0 9 2
11 0 9 15 13 3 3 1 9 11 11 2
13 0 0 9 13 9 11 11 2 0 1 0 9 2
9 1 9 2 9 13 15 0 9 2
25 11 7 10 9 13 2 16 13 1 11 0 9 0 2 16 1 9 1 9 1 9 2 4 13 2
10 7 13 1 9 2 0 9 0 9 2
31 3 0 9 2 9 11 2 0 0 9 11 11 7 10 0 9 11 11 2 12 0 0 9 0 9 2 4 13 13 9 2
8 0 9 13 7 3 1 9 2
16 1 0 2 15 13 0 2 1 9 9 2 15 13 1 9 2
28 1 0 1 9 9 2 16 13 0 2 16 11 13 13 15 0 9 7 4 13 13 1 9 2 16 3 10 2
17 7 1 15 3 7 9 4 13 10 7 15 9 2 1 15 0 2
14 0 9 13 7 3 0 2 13 15 9 9 0 9 2
27 16 1 12 9 11 16 9 1 9 13 3 1 11 7 11 13 3 9 16 11 2 13 9 3 3 0 2
26 15 3 13 3 0 1 0 9 9 2 13 15 7 9 2 15 15 12 9 1 9 14 3 3 13 2
13 11 13 0 9 1 9 2 15 13 9 0 9 2
14 1 0 9 2 0 9 2 4 15 7 13 0 9 2
16 15 9 1 10 0 9 13 2 16 13 13 13 9 3 13 2
12 15 13 0 9 2 15 13 13 0 9 9 2
7 1 15 13 7 0 9 2
15 13 3 0 2 16 0 9 9 13 9 3 0 7 0 2
15 7 1 15 2 1 3 3 3 0 9 2 13 13 9 2
30 13 2 14 3 9 1 9 9 2 15 15 13 2 1 10 9 13 3 15 13 2 13 15 1 1 0 9 3 0 2
19 7 16 0 9 0 9 15 13 3 0 2 0 9 1 9 9 3 13 2
41 0 0 9 2 9 9 9 7 3 9 1 9 2 9 1 9 7 9 2 0 9 7 9 9 1 9 2 15 13 9 2 15 11 13 1 0 1 9 10 9 2
42 0 9 1 9 1 0 9 13 10 9 1 0 9 2 1 0 0 9 2 0 0 9 7 0 1 9 11 2 10 9 13 15 0 9 2 0 0 9 2 3 13 2
50 9 11 11 3 3 13 2 16 0 9 16 1 11 2 11 2 0 0 9 2 0 1 9 11 2 1 11 13 1 9 2 7 9 0 9 2 1 9 1 11 11 2 7 10 9 3 3 3 13 2
16 9 13 0 9 2 1 0 9 9 11 13 3 16 1 0 2
17 12 9 1 0 9 11 7 13 3 2 16 12 9 1 0 11 2
13 0 9 2 11 2 1 0 9 13 3 0 9 2
19 0 9 13 2 13 3 0 2 9 11 11 13 9 9 2 3 0 9 2
43 9 15 13 15 2 16 13 0 1 0 9 9 11 2 11 2 15 13 2 16 1 11 10 9 13 13 1 9 2 14 1 0 9 2 7 15 13 0 9 10 0 9 2
58 13 2 14 7 3 1 0 9 3 12 0 9 2 11 2 11 2 11 2 11 2 0 7 11 2 13 9 0 2 0 2 0 2 0 2 0 2 9 2 11 2 11 7 0 2 0 0 9 7 1 11 2 11 7 11 1 9 2
9 15 15 3 1 10 9 3 13 2
23 1 0 9 7 13 7 1 9 11 2 7 11 2 16 0 9 1 1 0 9 0 9 2
16 12 9 3 13 1 9 7 0 9 13 0 9 10 0 9 2
7 13 15 13 3 0 9 2
16 3 0 9 13 2 16 0 9 1 15 9 13 14 0 9 2
15 4 2 14 0 9 13 2 13 3 1 0 9 0 9 2
24 7 1 9 13 0 2 16 16 3 9 13 3 2 11 13 0 9 1 11 2 0 7 0 2
5 11 2 0 9 9
7 0 9 11 1 11 11 11
19 3 16 12 9 15 1 11 3 13 9 9 15 9 1 9 0 2 11 2
12 0 9 15 3 3 13 1 9 1 0 11 2
17 1 9 12 2 9 13 10 9 3 0 2 7 10 9 4 13 2
11 1 12 9 9 7 9 13 11 9 9 2
8 15 3 13 11 1 0 9 2
6 13 15 3 0 9 2
16 11 15 13 1 10 9 10 9 7 1 15 13 0 9 9 2
13 13 15 3 2 16 0 13 0 9 0 0 9 2
18 9 7 9 11 11 15 13 1 9 10 9 7 9 0 11 15 13 2
47 16 4 11 13 3 13 1 9 2 16 4 15 1 15 15 13 2 13 4 15 3 12 2 15 13 7 13 0 9 2 13 15 0 9 11 11 2 1 12 9 3 7 3 3 3 13 2
25 15 9 9 9 13 1 0 9 1 0 11 7 13 0 7 0 9 7 3 9 3 13 16 0 2
11 11 13 10 9 1 0 9 16 0 9 2
27 12 12 9 0 9 14 3 13 0 9 1 9 2 13 3 9 11 2 16 3 13 0 13 1 0 9 2
10 9 13 2 16 9 11 15 13 0 2
14 0 13 13 0 2 16 0 9 3 10 0 9 13 2
17 11 15 3 13 15 3 15 0 9 2 1 0 9 3 0 9 2
9 3 3 3 13 9 1 10 9 2
21 9 11 11 2 0 9 11 2 13 3 0 10 9 1 9 7 15 15 13 9 2
35 3 15 9 1 9 3 13 9 2 16 16 4 15 13 16 3 11 11 1 0 11 2 7 0 9 1 11 2 13 4 15 1 15 13 2
34 9 11 11 2 0 9 1 0 11 3 3 13 2 16 11 3 13 10 0 9 1 0 11 2 10 0 7 0 9 15 1 15 13 2
10 3 13 9 2 15 11 11 3 13 2
9 9 9 1 12 7 9 9 9 2
10 15 13 9 3 0 1 0 0 9 2
15 11 3 13 0 9 2 16 7 13 0 9 1 0 9 2
29 1 15 15 11 13 9 2 16 4 13 0 9 2 16 1 12 9 9 9 4 9 11 11 13 13 1 0 9 2
33 9 11 13 1 9 11 1 9 1 9 11 7 10 9 13 3 3 0 2 1 9 11 0 0 9 16 11 7 11 1 0 9 2
9 4 12 9 9 9 1 9 13 2
21 0 9 9 11 11 13 3 1 9 1 0 9 2 16 4 13 0 9 0 9 2
19 7 11 3 13 0 9 9 7 9 2 3 4 11 11 13 4 13 3 2
14 0 9 13 2 16 7 0 9 15 3 13 10 9 2
15 0 9 3 13 2 3 15 9 13 2 10 9 13 0 2
22 9 4 9 9 13 7 13 9 11 2 0 9 13 12 9 7 1 15 15 15 13 2
7 9 11 13 3 9 9 2
19 3 15 13 2 15 15 15 1 9 13 2 3 2 3 2 1 0 9 2
19 9 15 0 9 2 16 15 1 0 9 3 3 13 11 11 1 11 11 2
6 9 7 9 0 9 2
8 15 15 13 1 15 9 11 2
20 15 15 13 1 9 2 15 1 0 9 13 9 1 9 7 3 13 1 9 2
9 1 0 9 3 13 9 0 9 2
18 9 1 0 11 13 9 1 0 9 2 15 15 3 13 13 0 9 2
32 13 7 7 0 0 9 2 16 0 9 11 11 2 15 13 1 9 7 13 0 9 2 16 4 13 9 11 7 3 13 9 2
6 14 15 9 3 13 2
13 9 9 15 7 13 3 12 9 2 16 13 9 2
11 16 13 1 9 12 9 9 1 10 9 2
12 15 15 7 12 9 2 0 7 0 3 13 2
16 9 11 3 15 13 1 11 2 16 4 15 1 15 3 13 2
8 0 9 13 7 10 0 9 2
14 1 12 9 15 9 0 9 13 1 12 1 12 9 2
7 9 3 13 3 0 9 2
33 1 12 9 15 3 13 0 9 2 16 9 13 3 3 9 7 15 11 13 9 7 9 2 0 9 9 1 9 13 13 1 9 2
4 11 11 1 11
18 0 9 11 11 13 1 10 9 11 11 11 1 9 1 0 9 11 2
7 9 13 1 0 9 11 2
6 3 15 13 0 9 2
9 0 9 9 13 1 11 9 9 2
9 1 11 13 9 1 0 9 11 2
13 11 9 13 3 3 2 13 3 3 16 0 9 2
27 9 0 9 2 15 15 1 10 9 1 9 12 13 1 0 0 9 2 13 2 16 15 13 1 0 9 2
11 9 15 3 13 9 1 11 1 0 9 2
12 13 7 2 16 0 9 3 13 10 0 9 2
6 9 9 13 0 16 9
10 11 11 1 0 9 0 11 13 0 9
2 11 2
53 3 12 9 1 9 11 13 9 1 0 9 0 2 16 4 0 9 9 13 10 9 1 0 9 3 13 1 0 9 2 13 4 15 0 0 9 1 11 2 11 7 0 11 2 13 11 11 1 0 9 0 11 2
21 1 9 10 0 9 13 0 9 9 9 9 2 15 3 13 0 9 7 0 9 2
11 11 3 13 13 0 0 9 0 0 9 2
15 9 0 9 7 9 0 9 1 9 13 3 0 16 9 2
28 16 4 1 9 12 1 0 9 13 14 12 9 2 1 9 0 9 1 0 9 4 1 11 13 7 0 9 2
12 1 0 9 13 0 9 0 9 2 13 11 2
13 11 4 3 13 0 0 0 9 3 1 11 11 2
26 11 2 11 2 11 2 11 7 3 11 13 3 2 16 1 11 13 0 16 9 1 9 1 0 11 2
24 11 13 3 13 2 16 1 11 13 13 0 9 1 11 2 7 16 15 11 13 1 0 9 2
3 9 9 11
7 11 11 2 0 9 1 11
30 11 11 13 9 12 0 11 0 9 11 2 11 1 9 1 11 1 9 9 2 9 9 2 11 12 2 12 2 2 2
47 13 2 16 15 9 13 1 9 9 11 2 16 9 2 0 0 9 2 7 15 7 1 0 9 9 2 0 1 9 2 3 13 13 3 9 2 13 9 9 1 10 0 7 10 0 9 2
57 16 9 16 0 9 0 15 15 2 15 1 11 13 1 11 2 13 3 13 1 9 2 16 11 13 1 9 2 0 7 0 11 2 3 9 0 9 2 9 9 3 0 7 0 2 9 1 0 9 1 11 2 1 15 13 9 2
16 15 9 11 1 0 9 13 2 3 9 15 2 7 3 9 2
32 9 11 3 13 7 9 2 16 1 0 9 4 3 13 0 9 2 15 3 13 2 16 7 1 11 15 13 9 0 9 2 2
27 1 10 9 7 0 0 9 13 9 1 0 0 9 2 7 1 9 11 13 1 9 9 0 2 3 0 2
14 13 4 7 0 9 2 16 1 9 13 3 2 11 2
10 1 0 9 9 11 1 10 9 13 2
42 9 1 0 9 13 1 9 1 9 9 2 16 11 2 11 1 10 9 13 2 16 1 0 13 9 2 1 11 3 13 0 9 2 3 3 13 0 0 9 7 9 2
17 13 0 15 13 15 1 0 9 7 9 2 15 1 9 3 13 2
22 9 0 13 9 1 9 1 9 7 9 2 0 9 7 9 13 9 7 9 1 9 2
9 3 9 1 9 10 0 9 13 2
49 3 3 2 16 4 13 0 9 7 16 4 3 13 2 7 3 2 16 4 9 13 2 1 9 9 2 1 0 7 0 9 0 9 10 9 2 4 0 9 3 12 3 0 9 3 13 1 9 2
28 9 4 13 3 3 3 2 16 15 13 2 16 1 9 9 2 9 2 1 15 13 2 13 7 3 0 9 2
12 9 11 7 13 15 0 16 9 9 16 15 2
23 10 9 1 15 9 2 3 0 0 9 2 15 1 0 9 13 1 0 9 16 1 0 2
31 15 3 9 13 7 3 13 2 16 4 4 13 1 0 2 7 13 15 13 2 16 13 15 3 10 9 16 9 0 9 2
31 1 9 1 11 2 11 15 7 13 2 16 9 11 3 13 1 11 0 2 7 1 10 9 13 2 15 13 0 1 9 2
44 7 16 11 2 11 1 10 9 13 7 0 9 0 11 2 16 15 7 15 2 15 15 13 2 13 3 1 11 0 2 13 13 2 16 3 15 13 15 2 15 13 3 13 2
6 15 13 1 0 9 2
30 15 9 13 7 3 3 13 13 1 10 9 7 9 2 7 3 13 13 2 13 1 0 9 2 1 9 1 0 9 2
25 14 2 3 9 13 0 9 1 9 2 3 15 1 10 9 13 2 16 10 9 4 0 9 13 2
16 13 4 2 16 9 11 10 9 1 0 9 3 0 9 13 2
15 14 2 3 3 2 16 13 1 11 2 7 1 0 11 2
5 1 9 13 14 9
4 11 11 2 9
43 1 10 9 2 0 0 0 9 2 11 12 2 12 2 12 2 2 15 10 0 9 11 11 13 1 15 2 16 4 15 1 9 13 15 2 1 9 2 7 15 9 13 2
13 9 2 15 15 13 1 9 2 13 1 0 9 2
15 13 2 1 15 4 10 9 3 13 2 13 15 7 0 2
26 13 15 13 2 16 15 13 2 16 15 0 9 1 12 9 13 3 1 9 2 1 15 15 15 13 2
10 13 15 9 1 15 3 14 3 0 2
9 9 13 13 3 1 10 0 9 2
22 3 11 11 11 2 9 0 9 2 13 1 0 9 1 3 0 9 1 9 0 9 2
41 9 9 15 1 10 9 1 9 13 3 1 9 1 9 0 9 2 7 3 9 0 9 2 11 11 15 9 0 9 13 1 15 2 15 4 13 13 9 9 9 2
21 0 9 1 9 1 9 9 1 9 1 9 7 9 15 13 1 9 9 0 9 2
18 13 0 2 16 0 9 15 1 9 0 9 13 3 16 9 9 9 2
21 15 13 1 9 9 0 9 2 3 15 7 13 15 9 13 9 9 9 7 9 2
31 9 11 2 11 13 13 9 0 9 2 16 4 15 13 13 2 3 15 3 1 9 13 15 2 1 9 1 10 0 9 2
11 13 2 16 4 15 13 9 1 0 9 2
14 1 10 9 13 15 3 3 3 2 16 9 13 9 2
39 3 15 13 3 0 9 1 9 0 9 2 1 9 0 0 9 2 1 15 2 16 15 1 15 13 0 0 9 2 1 15 2 16 4 13 9 2 2 2
25 0 1 15 13 13 2 16 1 9 13 3 15 1 9 7 16 9 1 15 13 3 3 1 9 2
21 3 13 2 16 16 15 13 13 3 12 9 3 0 9 2 13 4 13 3 3 2
8 3 7 15 1 9 13 15 2
7 3 15 13 9 1 9 2
6 13 15 0 9 9 2
14 13 2 16 13 15 1 9 2 7 9 15 3 13 2
5 9 9 0 9 2
13 9 2 11 11 2 9 2 2 9 9 7 9 11
19 9 0 9 4 13 1 9 0 9 9 1 0 9 7 1 9 0 9 2
40 10 0 9 9 13 10 0 9 2 15 13 3 13 1 9 0 9 2 3 15 13 1 10 0 9 7 9 0 1 0 0 9 2 3 3 1 0 9 2 2
32 13 7 1 0 13 1 10 9 0 9 2 15 4 13 4 3 13 7 13 3 2 16 4 9 13 1 9 0 9 1 9 2
58 9 0 9 13 1 15 2 16 15 0 9 0 0 9 2 0 2 0 2 3 2 0 2 13 13 2 16 0 9 2 15 1 9 0 9 13 2 7 13 2 2 4 13 3 0 0 9 2 7 16 10 9 4 13 1 0 9 2
22 9 9 13 4 13 1 9 1 9 7 1 0 0 9 2 0 0 9 0 9 2 2
11 0 9 9 15 3 13 7 1 9 0 2
30 9 0 9 13 9 0 9 15 2 16 13 13 10 9 0 2 0 2 1 0 9 0 2 7 0 9 0 9 9 2
13 9 9 0 9 1 0 9 13 3 13 0 9 2
13 0 9 0 9 13 10 0 9 1 9 2 9 2
14 10 9 0 9 4 13 13 1 0 9 1 0 9 2
57 1 9 0 9 13 3 9 0 0 9 1 0 0 9 2 9 2 9 2 12 2 12 9 2 2 1 0 9 1 0 0 9 7 9 0 9 2 9 12 7 12 9 9 2 12 2 12 9 2 2 1 0 9 1 9 2 2
21 0 0 9 13 7 13 0 9 2 15 4 10 9 13 1 0 0 7 0 9 2
36 10 0 9 13 1 9 10 9 1 0 0 7 0 9 0 9 9 2 15 13 0 1 10 9 16 0 9 2 15 13 3 13 9 1 9 2
53 13 0 3 13 2 16 0 9 1 11 15 10 0 7 0 0 9 13 0 9 1 9 7 3 2 15 15 13 7 1 3 0 9 0 9 2 1 15 9 13 10 0 9 1 9 9 2 15 1 15 13 13 2
25 9 0 9 1 15 4 14 3 13 1 9 9 1 9 1 0 9 2 0 0 7 0 9 2 2
29 13 0 13 2 16 0 9 1 9 1 0 9 0 1 0 9 13 9 0 9 1 9 7 1 9 1 9 0 2
25 1 10 9 9 0 9 13 0 9 0 9 2 15 13 0 9 9 1 0 9 7 9 0 9 2
29 0 9 9 13 7 1 0 9 10 9 2 15 13 1 9 1 9 0 9 7 15 15 13 1 9 0 0 9 2
34 13 3 3 1 9 2 1 15 13 9 9 9 9 2 13 1 15 2 15 1 10 9 13 4 13 2 3 15 1 10 9 4 13 2
12 9 13 7 0 9 2 16 13 1 9 13 2
27 3 15 9 1 10 9 1 9 9 13 0 9 2 13 9 2 9 12 2 12 7 12 0 9 9 2 2
38 13 7 13 1 15 2 16 1 9 9 13 4 13 3 0 9 0 9 7 15 2 15 13 0 9 2 9 12 9 2 12 0 2 9 9 2 2 2
66 15 10 0 9 2 15 4 13 13 0 9 0 1 0 0 9 9 1 0 9 2 13 0 9 7 13 15 13 3 14 3 2 16 15 13 1 9 1 9 9 0 9 0 9 1 0 9 0 9 11 2 7 7 3 2 16 15 13 1 9 1 15 9 0 9 2
21 13 0 13 3 1 9 2 16 13 3 0 9 1 11 2 15 13 9 0 9 2
29 0 0 9 2 0 9 13 9 1 10 9 7 9 0 2 13 9 0 0 9 7 9 2 15 4 7 4 13 2
26 7 16 9 0 9 1 11 4 1 0 0 9 13 2 10 10 9 15 15 1 10 9 0 9 13 2
55 0 0 9 9 1 0 9 13 0 13 1 9 1 0 9 9 1 9 0 0 7 0 9 1 0 9 2 1 15 15 1 9 1 3 0 9 9 12 9 2 9 2 12 2 12 9 2 3 13 9 0 9 1 11 2
24 0 9 9 0 9 15 3 3 13 7 1 9 10 9 2 15 4 1 9 3 13 1 0 2
48 3 9 13 13 7 0 2 0 9 9 12 0 0 9 9 2 1 15 9 12 7 12 13 9 3 3 9 9 2 7 2 9 1 15 2 15 13 13 9 7 1 9 9 0 9 9 2 2
11 9 10 9 4 9 0 0 9 4 13 2
18 9 2 16 3 0 7 0 2 15 4 15 13 2 4 13 3 0 2
12 9 9 2 16 0 2 15 13 3 14 3 2
4 13 1 9 2
5 15 2 10 9 2
2 11 11
6 3 2 3 2 11 2
6 1 9 2 0 11 2
8 1 9 2 15 2 10 9 2
11 13 15 3 12 7 3 4 3 13 9 2
11 0 11 2 15 4 7 9 11 3 13 2
10 1 9 0 9 1 11 13 3 3 2
15 0 9 15 13 0 9 2 7 3 9 1 9 0 9 2
13 0 15 9 2 16 13 9 0 9 2 13 3 2
6 13 3 0 9 9 2
10 12 0 9 13 9 0 9 0 11 2
7 15 13 2 16 4 13 2
6 7 4 10 9 13 2
12 13 4 1 15 9 7 1 9 9 7 9 2
3 0 9 2
6 11 13 10 0 9 2
10 11 11 9 10 2 3 16 10 9 2
19 9 13 9 2 13 9 7 16 13 9 2 13 15 13 3 3 1 9 2
7 10 9 13 7 12 9 2
6 13 1 0 9 9 2
16 12 9 4 13 1 9 2 16 9 13 2 16 13 1 9 2
25 0 0 9 2 1 9 15 10 0 9 1 10 9 13 2 13 9 1 10 9 2 1 0 11 2
15 0 9 1 9 12 13 9 2 13 0 9 1 0 9 2
11 9 7 10 9 9 1 15 13 1 9 2
15 1 9 15 13 0 0 11 7 3 0 9 13 1 9 2
11 9 13 9 9 7 3 13 1 0 9 2
4 13 13 9 2
10 1 0 9 3 13 2 3 15 13 2
14 1 0 9 13 2 10 9 15 1 9 13 0 11 2
11 0 9 2 3 9 15 1 15 13 13 2
6 9 13 1 0 0 2
11 13 4 11 1 9 2 13 4 9 9 2
16 4 13 0 2 16 13 11 7 16 10 9 13 3 9 11 2
5 14 14 12 9 2
7 1 9 15 13 1 9 2
12 0 9 15 13 9 2 9 7 9 1 9 2
15 13 15 15 0 16 0 9 0 0 9 11 1 0 9 2
9 13 4 15 13 1 9 1 9 2
4 3 4 13 2
6 13 4 15 3 3 2
4 9 15 13 2
20 13 4 15 2 13 4 15 2 13 4 9 2 13 15 7 13 1 15 9 2
7 13 15 1 15 0 9 2
6 9 9 4 13 9 2
4 3 15 13 2
10 11 13 7 0 7 9 15 3 13 2
10 13 15 9 2 7 3 13 13 9 2
5 9 9 2 13 2
13 13 4 15 1 11 2 7 11 13 3 10 9 2
10 13 3 3 0 2 3 10 9 13 2
13 13 3 3 12 9 2 7 3 13 9 0 9 2
6 7 13 11 1 11 2
3 9 1 9
9 9 13 1 9 7 9 1 9 2
15 3 1 15 13 2 14 14 11 2 15 13 0 0 9 2
7 9 11 2 9 0 11 2
8 13 1 12 9 1 0 11 2
11 1 12 9 13 1 9 1 9 0 9 2
3 13 13 2
10 1 12 9 1 15 13 9 1 9 2
13 16 15 1 9 13 15 13 2 13 15 1 11 2
14 3 15 13 9 2 13 0 9 15 2 9 7 9 2
5 13 11 16 9 2
22 9 13 0 9 0 2 13 7 13 9 9 7 13 4 0 9 2 16 9 7 9 2
3 15 14 2
11 1 9 13 11 7 9 12 9 0 9 2
4 11 13 3 2
7 0 9 13 2 9 13 2
5 13 1 15 9 2
8 13 12 9 7 13 15 13 2
3 13 9 2
8 12 9 1 15 7 13 9 2
5 13 1 15 9 2
20 12 9 1 9 1 15 13 9 2 16 13 1 0 9 7 1 9 1 9 2
23 0 0 9 9 9 3 13 1 9 0 9 2 1 9 2 1 9 7 9 9 0 9 2
30 15 4 15 13 2 15 4 13 9 2 16 15 15 1 9 13 2 3 15 13 2 7 3 13 2 15 1 15 13 2
4 13 1 15 2
8 1 0 9 15 3 13 9 2
10 3 15 13 2 13 2 13 2 13 2
14 13 12 9 3 7 7 3 13 9 1 9 0 9 2
5 3 1 11 13 2
3 3 1 11
5 9 15 13 11 2
2 11 2
7 0 9 15 3 13 11 2
4 1 9 9 2
7 11 13 0 7 0 9 2
8 13 15 7 13 3 1 15 2
5 0 11 1 11 2
4 9 13 9 2
11 1 9 0 9 15 13 1 11 1 11 2
8 13 11 0 9 1 0 11 2
11 13 15 1 9 12 7 13 15 1 11 2
11 15 4 13 1 9 1 9 9 0 9 2
15 1 11 15 10 15 13 2 1 12 9 15 11 13 13 2
12 14 13 3 10 9 7 3 13 3 1 11 2
5 13 4 1 11 2
11 1 9 11 13 11 13 1 12 9 9 2
10 9 13 3 9 15 1 0 11 13 2
31 15 15 13 2 3 4 3 3 13 7 7 1 9 4 15 13 2 16 15 0 9 9 0 9 13 2 16 13 0 9 2
14 9 11 2 9 11 2 15 1 12 9 13 16 11 2
14 3 15 13 13 0 9 2 3 15 10 9 3 13 2
2 0 9
7 9 13 0 9 1 9 2
6 7 13 13 1 9 2
16 15 3 13 2 16 1 9 9 4 13 9 0 16 0 9 2
13 16 4 13 2 13 9 7 3 1 11 15 13 2
13 15 3 13 2 14 15 4 15 13 1 9 3 2
13 9 13 9 1 9 1 0 1 11 3 1 11 2
11 13 1 0 9 7 10 9 15 3 13 2
6 9 4 13 1 9 2
6 11 15 3 13 9 2
9 15 13 3 10 0 9 1 15 2
14 3 3 0 2 16 16 13 2 13 3 9 0 9 2
3 0 0 9
8 11 13 0 2 16 13 9 2
4 13 15 15 2
4 13 2 13 2
7 14 12 9 1 15 13 2
5 13 15 7 11 2
16 16 13 0 9 9 2 3 13 3 11 2 3 15 3 13 2
12 7 15 13 14 0 2 15 15 1 11 13 2
11 1 12 9 13 1 9 12 9 1 11 2
17 13 14 0 9 7 9 2 4 15 1 15 13 1 9 1 9 2
14 16 13 1 0 9 2 13 3 0 16 0 9 3 2
26 13 15 7 9 11 1 0 9 9 2 0 9 3 13 1 11 7 0 9 0 9 7 13 1 9 2
25 13 11 2 16 15 0 13 2 16 10 9 3 13 2 16 13 9 9 2 15 1 10 9 13 2
7 9 9 4 11 3 13 2
5 9 3 15 13 2
11 9 13 0 7 13 10 9 1 9 9 2
8 11 15 3 13 13 0 9 2
10 0 9 13 1 9 9 9 0 9 2
18 1 11 1 11 15 4 13 0 9 1 9 9 16 1 9 0 9 2
22 9 1 9 9 7 13 7 10 9 2 15 13 2 16 13 0 9 1 0 0 9 2
20 1 9 2 15 15 13 1 12 2 9 12 2 13 1 9 9 0 9 9 2
12 0 15 3 13 3 3 2 13 7 3 13 2
18 1 9 0 1 12 2 9 12 13 9 9 9 2 7 0 9 9 2
19 3 3 13 14 12 9 2 15 13 9 0 0 9 7 13 13 0 9 2
29 1 12 2 9 4 10 9 13 1 9 9 9 2 13 9 1 0 9 1 9 7 13 4 16 9 13 1 11 2
8 9 11 13 1 9 0 9 2
11 13 15 1 11 2 7 9 9 13 0 9
1 9
3 9 7 9
1 9
29 9 2 12 0 9 0 9 2 15 15 3 1 12 9 13 1 10 0 0 9 2 13 0 0 11 1 0 9 2
35 9 2 9 7 9 3 0 0 9 11 0 11 2 3 0 9 0 9 2 15 15 13 11 2 7 0 0 9 2 0 0 9 0 11 2
24 9 13 0 9 11 0 11 2 15 15 1 9 13 1 0 9 1 0 9 1 9 7 9 2
45 0 9 9 2 9 2 9 7 9 11 11 2 0 1 0 0 9 1 0 9 1 9 2 1 3 0 9 3 0 9 2 3 11 7 0 11 1 9 11 2 13 3 0 9 2
24 7 1 0 9 11 13 3 0 7 3 3 0 9 3 9 12 1 0 7 0 0 9 9 2
23 16 11 13 1 9 2 0 0 2 0 9 0 9 11 4 1 0 9 1 0 9 13 2
21 0 9 11 1 9 0 9 13 1 0 2 3 0 2 0 9 7 0 0 9 2
21 14 3 11 13 1 10 9 7 0 9 2 15 15 15 13 13 1 13 0 2 2
13 11 9 13 1 9 2 16 0 9 9 13 0 2
30 16 1 9 9 13 1 0 9 7 13 15 3 1 9 9 2 3 9 13 1 9 7 1 9 15 13 0 9 9 2
14 11 0 9 7 13 1 0 12 3 0 9 7 9 2
25 1 0 9 15 13 9 0 11 2 15 3 1 0 9 0 9 15 13 15 13 7 13 0 9 2
64 0 0 9 9 2 0 0 9 2 7 0 9 11 11 13 1 0 0 9 2 1 15 13 14 9 1 0 9 11 0 2 11 1 0 11 7 11 12 2 2 7 7 9 0 9 1 9 0 2 15 13 1 0 11 2 11 2 15 13 3 15 13 2 2
28 0 7 3 0 0 9 2 15 3 13 0 2 3 0 9 2 13 12 1 0 9 9 2 0 0 15 3 2
25 1 0 9 15 9 13 1 9 14 12 0 9 0 11 2 15 15 9 1 15 13 1 0 9 2
2 11 11
9 11 0 11 2 11 2 0 11 2
11 12 2 9 12 2 9 2 9 2 11 2
9 13 9 0 2 11 7 11 11 2
25 1 9 11 2 15 1 9 0 9 13 1 11 1 10 0 0 9 2 4 15 13 13 9 9 11
2 9 9
20 1 10 9 13 9 9 9 2 13 2 13 9 2 2 2 9 2 3 13 2
6 0 9 13 1 9 2
10 0 9 0 9 0 9 2 9 15 2
9 9 9 13 13 15 1 10 9 2
6 9 11 11 7 11 11
7 15 15 13 3 2 2 2
1 9
19 9 2 0 9 2 0 9 1 10 0 9 2 0 0 9 7 0 9 2
26 3 15 13 13 0 9 11 11 2 12 2 7 11 11 2 12 2 1 0 11 1 0 9 0 9 2
24 9 2 15 13 3 1 9 12 7 13 3 3 1 9 12 2 13 9 9 2 9 2 9 2
49 1 9 9 7 9 15 13 7 10 0 9 1 11 11 2 0 3 10 9 1 9 2 13 1 15 9 9 13 9 0 2 13 2 16 9 3 13 10 9 7 3 13 3 3 2 16 15 13 2
15 9 0 2 0 9 13 1 0 0 9 0 1 0 9 2
18 9 13 0 0 9 15 2 15 13 2 7 15 2 15 4 9 13 2
24 9 15 13 16 0 9 9 7 13 9 2 15 7 13 9 2 3 0 7 3 0 2 13 2
9 9 13 0 9 10 9 0 9 2
18 9 15 13 9 9 2 7 16 15 13 2 16 13 1 9 9 9 2
13 13 2 14 0 7 11 9 2 3 15 3 13 2
2 11 11
6 9 2 9 2 9 2
6 11 11 2 11 11 2
9 0 11 2 0 0 11 2 11 2
7 12 2 2 12 2 9 2
5 9 13 1 9 9
9 9 11 13 0 9 14 1 9 9
2 11 11
13 0 9 3 1 9 1 3 12 9 9 13 9 2
30 3 15 3 13 7 0 9 2 0 0 9 1 0 9 1 0 9 2 15 3 1 9 12 13 0 0 9 11 11 2
42 9 0 9 11 11 11 2 1 0 9 0 9 0 9 7 0 9 2 10 9 1 11 13 2 7 1 9 1 11 13 7 9 9 13 1 9 9 9 0 9 11 2
4 9 9 13 9
16 0 4 13 1 15 0 2 15 3 13 2 1 9 1 9 2
11 3 4 13 0 9 1 0 9 2 13 2
14 13 3 11 11 2 11 11 2 11 11 2 0 9 2
12 0 9 13 1 11 13 0 9 1 0 9 2
6 1 9 7 3 13 2
33 0 9 13 1 9 0 9 9 2 15 9 1 9 1 9 0 9 7 0 0 9 1 0 9 0 7 1 9 13 0 0 9 2
19 0 9 9 13 13 9 9 9 2 15 4 15 13 13 1 9 0 9 2
9 15 13 2 9 13 2 13 11 2
16 3 4 3 13 2 16 4 9 13 1 0 9 7 1 9 2
14 13 15 3 14 1 9 1 9 2 16 4 9 13 2
25 16 4 1 15 13 2 1 9 2 3 3 4 13 1 9 2 16 4 13 2 16 13 3 13 2
15 9 9 15 13 13 2 16 1 15 10 9 13 10 9 2
15 3 9 9 13 3 3 9 7 1 9 2 3 13 0 2
17 0 9 2 7 1 11 13 15 9 3 2 13 1 9 9 9 2
17 15 4 9 13 7 16 9 13 0 9 9 12 9 1 0 9 2
15 9 9 11 15 13 9 0 0 9 2 13 7 9 0 2
32 9 13 1 9 7 9 0 9 2 15 1 0 9 7 1 9 11 13 1 9 7 1 0 0 9 4 13 0 7 0 9 2
17 13 4 1 9 1 9 2 16 1 9 13 7 9 2 13 11 2
14 0 9 1 11 3 10 9 13 2 0 13 3 0 2
25 0 0 9 13 1 9 11 9 1 9 0 9 2 10 0 9 0 0 9 9 7 0 9 13 2
5 0 9 13 9 9
34 9 11 15 13 13 1 10 9 2 15 1 11 13 9 1 9 2 1 15 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2
9 13 2 13 2 13 7 9 9 2
17 9 13 13 1 9 1 0 9 0 2 12 9 9 1 9 2 2
12 13 15 0 2 7 7 0 9 2 13 11 2
17 13 4 3 1 11 9 2 16 15 13 3 2 15 15 9 13 2
15 1 12 9 13 10 9 3 7 1 9 1 12 9 9 2
22 9 4 1 9 1 11 13 13 9 2 9 0 9 4 14 13 13 9 2 13 11 2
21 13 3 0 0 9 0 9 2 3 12 9 13 3 13 9 1 0 7 0 11 2
7 9 14 2 7 1 9 2
11 0 9 13 9 9 15 1 15 2 13 2
18 1 3 0 0 0 9 4 9 11 0 13 9 1 9 0 0 9 2
30 15 13 9 13 3 2 16 4 13 0 9 2 15 1 0 9 3 13 14 1 0 9 2 7 3 7 3 1 9 2
27 9 0 9 11 11 2 15 15 1 0 9 13 9 13 0 9 2 13 13 9 11 3 1 0 0 9 2
32 3 16 1 9 0 9 13 11 11 11 1 0 9 1 11 7 1 11 7 1 9 1 15 2 15 3 3 1 0 9 13 2
14 13 3 9 13 0 9 1 3 0 0 9 2 13 2
9 9 4 13 1 11 13 1 9 2
12 3 3 13 13 3 1 9 9 2 13 11 2
15 13 7 13 2 16 15 9 1 15 7 9 13 10 9 2
11 11 11 7 11 11 1 9 9 9 1 9
5 9 11 11 2 11
7 9 2 15 13 9 7 9
11 0 9 11 2 11 7 11 4 13 9 3
2 11 11
30 9 1 9 2 0 11 2 13 9 0 9 2 15 1 12 0 9 13 11 11 11 2 11 11 11 7 11 11 11 2
33 13 15 1 9 0 9 0 0 11 1 11 7 10 0 9 4 1 11 2 3 13 9 3 1 9 9 2 13 13 7 1 11 2
36 9 15 13 1 12 9 2 0 2 0 11 2 13 11 11 1 0 9 11 7 11 0 2 0 9 0 9 2 0 2 7 0 9 11 11 2
29 0 9 9 13 9 0 11 2 0 9 2 7 1 9 11 11 2 0 9 1 9 0 9 2 15 13 11 11 2
11 0 9 13 0 9 11 11 0 0 9 2
16 9 10 9 2 15 13 9 11 2 13 11 11 7 11 11 2
20 9 0 9 15 13 3 9 2 0 9 11 11 11 2 11 11 7 11 11 2
41 1 11 11 2 15 13 9 7 0 9 0 9 2 13 10 9 13 0 9 0 9 2 1 15 15 13 9 9 1 9 0 1 0 9 9 7 0 9 1 9 2
34 9 0 9 7 9 4 3 13 1 9 13 7 9 2 15 3 3 1 0 9 13 2 7 13 15 1 0 0 9 2 9 7 9 2
19 13 15 9 1 0 9 2 3 1 0 9 9 13 3 9 0 11 11 2
26 10 9 13 11 1 3 0 16 9 15 2 16 4 13 1 0 9 2 16 1 15 13 10 9 0 2
25 9 9 13 9 9 9 2 9 0 9 2 0 9 9 0 2 9 0 9 7 0 9 7 9 2
20 1 12 2 9 15 9 1 9 4 13 1 9 2 1 10 0 9 15 13 2
5 15 2 3 2 3
23 11 11 2 0 11 13 9 9 2 15 13 1 0 0 9 9 2 12 13 1 12 2 9
27 9 9 13 1 9 9 0 9 7 9 11 11 2 11 11 2 11 11 2 11 11 2 11 11 7 0 2
7 9 13 1 12 2 9 2
7 1 0 11 15 13 9 11
2 11 2
31 3 1 9 13 0 9 11 1 11 14 1 0 9 3 12 12 9 9 7 9 1 9 11 2 13 0 9 9 11 11 2
23 1 9 13 1 10 9 9 14 12 9 2 7 10 9 4 13 13 1 9 14 1 12 2
17 0 0 9 9 13 1 9 10 0 9 11 11 3 9 9 9 2
23 0 9 13 14 12 9 0 9 2 12 9 13 9 1 9 7 12 9 9 13 0 9 2
27 10 9 3 9 13 2 3 1 0 9 1 9 9 7 1 9 0 0 9 2 1 15 13 15 10 9 2
23 0 9 9 1 11 13 1 9 0 9 2 15 13 1 9 3 12 7 13 3 0 9 2
12 1 9 9 13 9 1 11 2 11 0 9 2
19 1 9 13 9 3 12 9 2 15 13 1 0 9 0 9 12 9 9 2
10 1 0 9 15 13 3 1 12 9 2
23 9 9 13 12 12 9 9 1 9 2 1 9 9 13 15 12 7 12 12 9 1 9 2
21 1 9 11 2 11 4 1 9 0 9 13 9 3 13 12 7 12 9 9 9 2
18 9 0 9 13 9 11 1 11 2 11 2 11 7 9 12 11 9 2
24 0 9 9 13 12 9 9 7 1 11 2 11 10 9 13 1 9 0 9 1 9 10 9 2
7 1 9 9 3 13 13 2
15 9 1 9 1 9 9 15 13 1 9 1 12 9 9 2
8 0 0 9 4 3 13 1 9
39 1 9 1 9 7 0 9 1 0 2 0 7 0 9 4 3 1 9 13 0 9 0 0 9 2 0 9 0 9 9 1 11 2 11 1 0 11 2 2
39 0 9 13 3 0 1 0 0 9 11 11 2 12 2 2 0 9 7 13 1 9 7 4 13 14 1 9 9 2 9 1 9 1 15 13 11 11 2 2
31 9 1 11 1 9 11 11 13 1 0 9 9 11 2 15 3 13 13 1 10 0 9 9 9 2 0 0 9 0 9 2
26 9 10 0 0 0 0 9 13 1 9 11 11 1 9 12 2 0 9 15 7 13 3 1 9 12 2
35 9 13 9 9 2 3 0 9 0 9 1 9 2 7 10 9 13 0 9 9 11 11 1 11 2 0 0 11 0 2 9 7 9 2 2
18 11 13 1 9 0 9 11 2 13 1 10 9 7 13 15 9 11 2
34 11 9 0 9 1 12 9 1 12 12 9 2 15 4 13 0 0 9 2 13 9 0 9 1 10 0 0 2 9 1 9 0 9 2
3 2 11 2
10 9 1 0 9 4 13 2 9 15 13
20 9 0 9 1 11 7 11 7 0 9 13 1 9 1 11 1 9 0 9 2
20 9 0 9 4 13 7 9 4 13 3 3 2 13 9 9 0 9 11 11 2
19 9 13 1 3 0 9 2 15 13 9 9 2 7 13 7 9 9 15 2
46 0 9 9 11 11 9 0 0 9 2 11 2 1 11 11 11 7 11 11 1 10 9 1 9 9 11 11 12 2 9 1 11 13 2 16 4 13 0 9 1 9 0 9 1 11 2
13 1 0 9 4 13 12 9 9 2 15 4 13 2
18 0 9 9 0 9 13 3 12 2 7 12 2 9 1 9 1 11 2
14 4 13 0 9 2 15 13 9 0 9 2 13 11 2
29 9 13 1 10 9 9 1 15 2 16 0 9 4 15 13 7 15 13 7 7 12 4 1 15 13 0 2 13 2
10 13 7 9 13 1 9 1 9 9 2
13 11 3 13 2 16 0 9 13 1 9 9 13 2
22 1 9 9 2 1 0 7 0 9 0 9 2 3 13 4 13 2 13 12 9 9 2
17 9 13 0 9 3 2 16 4 13 0 9 0 9 16 1 11 2
10 9 13 0 9 12 9 7 0 9 2
3 11 1 9
1 9
12 9 2 9 11 13 1 0 0 9 0 9 2
42 11 11 13 1 10 9 0 9 16 11 11 1 11 2 10 9 2 9 11 11 2 13 0 0 9 7 9 2 9 11 11 2 13 9 0 0 9 2 0 0 9 2
20 9 9 9 9 13 1 0 9 0 9 1 0 9 11 1 9 0 7 0 2
13 9 13 0 9 9 9 0 9 0 9 11 11 2
15 0 0 9 0 9 4 7 13 2 3 0 9 1 9 2
18 0 9 4 3 13 1 0 9 2 15 13 13 3 0 16 0 9 2
33 1 0 0 9 1 9 7 9 7 9 9 9 3 13 15 1 9 2 14 1 12 2 13 15 11 0 2 7 3 0 7 0 2
21 11 11 0 2 7 0 2 13 1 10 0 7 0 9 3 0 7 3 3 13 2
26 1 0 9 11 4 13 3 0 13 9 7 1 0 0 9 2 16 13 10 9 7 11 9 0 9 2
32 1 0 9 0 0 9 9 9 13 3 0 9 1 0 9 9 2 7 4 13 3 3 2 1 0 9 2 0 9 7 9 2
2 11 11
7 9 9 2 0 0 9 2
8 9 0 9 2 12 2 9 2
11 1 0 11 1 9 2 9 2 9 7 9
23 9 9 2 0 1 0 0 9 9 2 7 2 1 0 9 0 11 2 13 1 11 13 2
21 16 11 13 9 0 9 0 11 11 11 2 13 3 14 13 0 9 7 0 9 2
24 1 0 9 4 13 1 9 12 9 2 7 1 9 9 13 3 3 0 9 1 9 12 9 2
35 9 0 9 15 3 13 14 1 12 9 2 3 1 12 9 3 2 16 16 13 13 1 9 2 7 9 4 1 10 9 13 12 0 9 2
24 9 1 12 9 13 9 1 9 2 15 0 9 15 13 1 12 9 2 13 3 1 9 9 2
17 1 9 9 1 15 13 9 13 10 9 2 9 7 3 7 9 2
20 3 13 3 13 3 9 2 9 2 9 7 0 9 1 9 0 7 0 9 2
13 1 9 9 3 13 0 9 13 7 13 0 9 2
3 2 11 2
11 9 1 9 1 9 0 11 2 9 2 12
14 11 11 2 3 2 1 9 10 0 9 1 11 11 11
5 9 11 11 2 11
2 11 13
1 9
30 9 2 10 9 2 9 9 7 0 9 2 9 9 7 9 7 1 0 9 7 9 11 13 9 0 9 9 9 9 2
25 0 9 3 0 9 13 10 9 0 11 2 15 13 1 11 7 1 0 11 2 7 9 11 11 2
29 0 9 9 2 9 1 9 9 11 11 2 11 2 11 2 13 11 3 3 2 9 13 0 9 2 9 7 9 2
17 0 0 0 9 9 9 13 3 0 9 11 2 7 7 0 9 2
13 13 3 3 3 0 9 13 1 0 9 0 9 2
22 0 0 9 11 11 13 11 1 3 0 9 2 16 13 0 2 3 9 7 3 9 2
10 3 13 10 3 0 9 7 0 9 2
12 3 7 9 13 10 0 9 7 9 10 9 2
15 9 15 13 3 0 9 2 7 1 9 10 0 9 9 2
16 0 9 9 15 7 13 9 12 2 9 9 9 11 1 11 2
20 9 1 15 13 3 0 9 2 3 0 7 0 2 1 0 9 7 0 9 2
33 16 0 9 0 0 9 0 9 13 0 0 7 0 9 10 0 9 2 3 0 2 2 13 0 9 1 9 0 9 3 16 0 2
2 11 11
16 9 9 2 0 11 2 11 11 2 9 2 11 11 2 9 2
9 0 9 0 9 2 12 2 9 2
7 11 14 13 1 0 2 11
5 11 2 11 2 2
16 9 0 0 9 11 11 15 3 3 13 1 9 1 0 11 2
12 9 4 13 4 13 1 12 9 1 0 9 2
32 1 9 4 13 3 1 12 2 9 2 3 4 1 9 9 10 0 9 11 11 11 11 1 11 13 4 0 9 13 1 9 2
3 1 11 2
2 11 2
14 1 0 9 9 0 9 1 11 4 11 3 13 11 2
12 1 0 9 15 3 13 13 10 9 11 11 2
21 15 9 7 9 11 1 9 13 2 16 15 13 3 1 9 7 13 1 9 13 2
18 0 0 9 7 13 1 11 2 11 7 0 0 9 9 1 10 9 2
18 9 1 11 13 9 2 16 15 13 13 9 2 16 4 4 11 13 2
4 9 1 9 13
4 11 1 11 2
21 1 9 0 9 0 9 13 1 9 0 9 9 1 0 7 0 9 2 11 2 2
14 1 0 9 3 13 1 9 9 7 0 9 1 9 2
18 1 0 0 9 4 1 9 0 9 12 13 0 9 1 9 0 9 2
17 0 0 9 9 0 9 1 11 3 13 1 3 16 12 12 9 2
12 0 9 1 0 9 15 13 1 12 9 9 2
15 3 1 0 9 13 1 9 0 9 12 9 0 0 9 2
20 10 9 13 3 2 0 9 2 1 15 13 3 0 9 9 1 9 0 9 2
10 11 13 3 0 13 3 0 9 9 2
23 9 0 9 2 15 9 13 9 9 2 15 13 0 0 9 2 15 13 9 13 7 13 2
36 10 9 9 0 11 15 13 1 3 0 9 1 9 0 0 9 2 15 13 1 11 2 11 1 3 15 0 0 7 0 9 7 0 9 9 2
15 3 12 9 0 9 13 0 9 0 9 2 3 1 11 2
8 13 15 3 1 0 0 9 2
2 14 9
2 11 2
21 9 0 9 9 1 0 9 9 2 11 11 15 3 13 1 9 0 9 9 11 2
15 15 4 13 1 9 1 9 0 9 1 11 0 9 9 2
15 1 9 15 13 2 16 10 9 13 1 9 13 3 9 2
24 9 2 11 1 15 13 2 9 13 0 9 2 0 9 0 9 2 7 7 13 1 9 9 2
12 10 9 13 1 0 7 13 15 3 9 9 2
23 9 11 11 1 0 0 9 9 9 13 2 16 15 13 1 9 3 3 13 9 16 9 2
2 0 11
2 11 2
26 1 9 1 12 9 0 9 9 1 9 1 0 9 1 11 13 11 11 2 11 0 0 9 9 12 2
18 13 3 0 9 11 11 11 1 12 2 9 12 2 15 9 13 12 2
27 0 9 11 1 9 0 9 1 12 9 13 0 9 1 12 2 12 2 14 1 12 9 1 10 0 9 2
26 1 3 0 9 1 9 2 3 13 0 2 15 1 0 9 13 1 0 9 7 15 13 14 1 9 2
7 13 11 11 11 2 11 2
2 0 9
2 11 2
36 0 0 9 13 1 10 12 2 9 1 11 9 1 9 2 1 15 4 1 15 9 13 1 0 0 0 9 0 9 7 1 0 0 9 9 2
17 13 15 2 16 1 3 0 9 4 3 13 1 9 1 15 9 2
12 0 9 11 3 4 13 11 1 11 1 11 2
5 0 9 1 9 11
18 9 9 9 1 12 9 2 11 2 11 12 2 12 2 12 2 12 2
5 11 2 11 2 2
26 0 0 9 1 3 0 9 10 9 1 0 9 9 9 9 1 12 9 13 10 0 9 9 1 9 2
12 1 3 0 9 11 15 10 9 14 3 13 2
41 1 12 2 9 13 1 0 9 2 3 1 9 1 11 1 0 9 13 9 1 9 9 7 10 9 1 9 14 0 9 2 7 11 15 1 9 13 3 1 9 2
19 9 1 0 15 3 13 2 7 7 1 0 9 13 9 13 3 9 9 2
16 0 9 13 9 11 1 15 2 11 13 11 2 7 15 13 2
14 3 1 9 9 3 1 9 9 3 13 11 1 9 2
15 1 9 1 11 13 11 9 1 9 0 9 3 1 9 2
3 9 1 11
2 11 2
23 12 0 9 1 9 0 15 13 9 2 15 15 13 1 12 2 1 12 2 9 1 11 2
28 1 9 13 1 12 9 11 2 1 12 9 11 2 1 12 9 11 2 1 12 9 11 7 1 12 9 11 2
3 1 0 9
20 11 11 11 2 11 1 11 11 13 1 9 9 0 0 9 0 9 9 9 2
1 3
14 0 9 11 11 4 13 0 9 9 1 0 0 9 2
13 0 9 9 4 7 1 0 9 13 1 9 9 2
36 11 7 11 13 1 9 0 9 1 0 9 1 11 1 12 2 2 12 2 9 2 16 1 0 9 13 1 0 9 11 2 11 12 2 12 2
9 9 13 0 11 11 7 1 11 2
10 9 9 2 1 11 2 7 1 15 2
21 11 7 11 13 1 0 9 3 9 2 7 13 15 13 3 1 12 1 11 1 11
7 11 2 11 2 11 2 2
34 1 11 2 7 1 15 2 15 13 0 9 9 0 0 9 11 11 2 15 13 13 1 0 0 9 9 9 1 12 1 11 1 11 2
47 9 11 13 13 12 9 9 2 1 11 3 9 9 7 1 11 1 9 2 1 11 7 11 2 13 4 9 11 2 7 1 9 14 1 9 9 2 7 1 11 2 2 16 0 0 9 2
20 1 0 9 13 0 2 16 11 13 9 9 2 3 1 10 9 13 3 11 2
6 13 2 16 4 13 2
26 7 3 13 2 1 11 4 15 13 1 9 7 1 9 10 9 13 1 9 9 0 9 2 13 11 2
26 7 9 11 15 13 0 2 16 11 13 1 10 0 9 3 3 3 2 3 13 13 9 10 0 9 2
13 1 0 0 9 1 11 4 13 12 9 9 9 2
16 13 15 3 9 2 16 15 13 1 9 9 13 2 13 11 2
19 1 9 1 0 9 15 1 9 13 9 1 9 2 13 9 11 2 11 2
20 11 3 13 2 16 7 12 1 15 13 1 0 9 9 1 0 9 10 9 2
15 11 9 13 2 7 9 13 2 11 15 13 2 13 11 2
11 12 9 13 1 9 9 3 1 0 9 2
31 0 7 13 13 15 12 9 1 9 2 13 12 2 12 2 13 11 2 15 3 1 0 0 9 3 13 9 9 1 9 2
29 11 15 13 0 2 16 9 9 9 15 3 3 2 3 15 13 1 9 1 9 10 9 14 1 9 12 2 13 2
12 9 13 3 7 3 12 12 9 4 13 13 2
19 15 7 3 3 13 3 1 9 2 13 9 7 3 15 15 13 1 9 2
28 15 13 0 2 16 15 0 16 9 2 1 15 0 1 9 13 9 12 12 9 2 4 4 13 1 0 9 2
30 11 7 0 9 13 9 2 3 3 2 13 11 12 2 12 2 11 12 2 12 7 13 1 11 1 11 12 2 12 2
43 1 0 9 13 12 9 9 9 12 2 3 0 2 9 1 10 9 13 9 1 0 9 2 9 11 7 3 3 0 9 11 2 13 1 0 11 2 7 13 15 3 2 2
35 15 13 9 9 7 13 15 12 2 1 10 9 13 2 13 11 2 15 1 0 9 13 10 9 9 15 11 2 16 4 15 10 9 13 2
11 13 1 15 7 11 2 15 13 9 9 2
11 13 0 9 2 7 13 15 13 0 9 2
7 13 3 9 4 13 9 2
22 1 0 9 15 13 13 9 3 1 11 2 11 7 11 2 13 9 11 11 11 11 2
16 9 13 1 12 9 1 9 0 9 11 2 13 15 9 11 2
29 0 9 11 2 11 2 11 2 11 2 11 2 11 2 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2
35 1 9 13 9 12 2 0 9 9 2 9 2 9 2 9 7 0 9 9 13 15 1 9 7 9 1 9 2 3 15 15 1 0 9 13
3 2 11 2
5 9 11 11 2 11
19 0 9 11 11 13 1 9 1 9 9 2 3 13 3 1 11 9 1 9
2 9 9
4 11 1 9 0
14 1 9 0 0 1 0 11 13 0 9 0 0 11 11
8 0 9 11 1 0 11 11 11
20 1 12 9 13 0 9 11 11 2 12 2 0 2 3 1 9 9 0 0 2
22 11 11 11 2 12 2 2 13 1 12 9 1 0 9 12 2 12 2 12 2 12 2
29 1 0 9 1 11 11 11 2 12 2 2 13 1 15 2 15 1 9 15 3 1 9 13 1 0 11 1 9 2
13 1 0 12 9 13 0 9 11 11 2 11 11 2
33 0 0 9 13 9 11 2 11 12 2 12 2 12 2 12 2 12 2 12 2 12 2 2 16 1 0 0 9 13 12 2 12 2
11 1 0 9 13 11 11 3 3 1 9 2
22 3 1 11 13 3 3 3 1 0 9 9 11 2 11 12 2 12 2 12 2 12 2
18 0 9 9 2 0 9 2 3 13 11 9 9 1 0 1 9 0 2
11 14 15 13 10 9 13 0 9 1 9 2
18 11 13 0 12 9 2 1 15 13 12 2 12 2 7 15 15 13 2
10 3 13 2 16 15 15 13 0 9 2
22 7 1 0 9 4 15 13 9 1 12 2 12 7 3 13 13 15 3 2 13 11 2
21 1 9 12 2 12 7 12 2 12 13 12 9 7 9 13 14 1 12 9 3 2
16 13 4 2 14 11 2 3 0 2 3 13 2 13 15 11 2
18 1 11 13 13 3 2 7 16 4 13 1 15 2 15 15 11 13 2
20 16 4 13 10 9 2 7 13 0 2 16 10 10 9 3 3 13 7 13 2
18 7 11 13 7 0 9 2 7 1 11 13 3 13 2 13 15 11 2
18 11 13 0 9 7 9 9 12 11 11 2 12 2 2 0 12 9 2
13 0 9 9 13 10 9 9 11 1 11 2 11 2
21 1 10 0 0 9 15 1 0 11 13 9 11 0 0 11 11 2 12 2 2 2
49 3 2 16 12 2 9 13 0 1 11 11 2 12 2 2 2 15 13 1 9 11 2 12 2 2 1 12 9 12 2 12 2 12 2 12 2 12 2 12 2 13 1 9 0 0 9 11 11 2
46 9 9 15 13 1 12 2 9 13 0 9 1 11 2 12 2 2 2 7 11 11 2 12 2 2 0 9 13 1 12 9 2 16 0 12 13 2 7 13 15 15 1 0 9 15 2
21 11 15 13 13 15 2 16 16 0 13 11 1 0 0 2 7 15 1 9 12 2
42 1 9 11 7 11 13 1 0 11 11 11 11 2 12 2 2 2 15 15 9 1 10 0 0 9 13 1 11 2 11 2 12 2 2 7 3 11 2 12 2 2 2
28 11 2 15 15 13 1 0 9 1 9 2 13 12 2 12 2 12 2 12 2 12 2 12 2 12 2 12 2
19 13 3 0 2 16 16 15 13 9 7 13 1 0 9 2 13 0 9 2
18 1 11 7 11 13 2 3 13 9 2 13 11 0 9 1 10 9 2
2 0 9
4 15 4 13 2
12 9 2 1 12 2 7 12 2 9 13 9 2
49 9 2 12 2 9 2 1 12 2 9 13 9 2 1 12 2 13 12 9 12 9 2 1 12 2 13 12 9 12 9 2 1 12 2 13 12 9 12 9 7 1 12 2 13 12 9 12 9 2
41 12 2 9 2 1 12 2 7 12 2 9 13 9 2 1 12 2 9 12 9 12 9 2 1 12 2 13 12 9 12 9 7 1 12 2 13 12 9 12 9 2
33 9 12 1 12 2 1 12 2 9 13 12 9 12 9 2 1 12 2 13 12 9 12 9 7 1 12 2 13 12 9 12 9 2
30 9 2 1 12 2 9 13 12 9 12 9 2 1 12 2 13 12 9 12 9 7 1 12 2 13 12 9 12 9 2
45 9 2 1 12 2 9 13 9 2 1 12 2 13 12 9 12 9 2 1 12 2 13 12 9 12 9 2 1 12 2 13 12 9 12 9 7 1 12 2 13 12 9 12 9 2
4 0 13 1 0
7 11 13 9 2 13 14 11
5 11 2 11 2 2
18 1 0 9 9 1 11 13 13 0 9 1 0 9 9 9 11 11 2
22 1 9 11 3 13 0 9 2 9 11 11 11 2 9 11 11 11 7 9 11 11 2
7 3 0 9 15 7 13 2
15 9 11 1 9 13 1 0 9 7 9 1 11 3 13 2
43 3 15 13 13 15 1 0 9 0 9 1 9 2 7 13 15 1 10 9 2 16 15 3 13 2 16 9 11 13 12 9 13 2 13 15 9 11 2 11 11 2 11 2
11 0 9 4 13 14 3 1 9 1 11 2
23 9 4 13 1 0 9 2 7 9 11 13 7 7 15 1 10 0 9 13 2 3 13 2
44 1 9 1 12 4 15 13 13 3 2 13 15 9 11 7 0 9 11 13 2 13 15 9 2 16 9 13 9 9 2 11 2 3 13 9 9 9 2 7 15 13 15 13 2
4 9 13 0 2
8 1 11 4 13 13 0 9 2
38 11 11 15 3 13 1 15 2 16 9 2 15 3 13 9 1 9 2 13 0 3 13 9 9 2 7 3 13 2 16 13 13 3 13 1 0 9 2
15 1 11 3 13 3 9 9 1 9 11 2 15 13 13 2
19 13 13 9 1 9 2 7 3 3 0 9 13 9 9 1 0 0 9 2
3 11 13 9
5 11 2 11 2 2
32 0 9 13 1 12 2 9 3 0 0 9 2 15 4 13 1 0 0 11 13 9 9 11 11 7 9 11 3 12 9 9 2
22 3 10 9 4 13 13 1 11 12 9 0 9 2 13 9 11 9 0 9 11 11 2
17 3 7 13 9 2 16 4 15 9 1 11 15 13 15 0 9 2
25 1 0 9 4 15 3 13 2 16 11 13 3 13 1 9 2 3 0 9 13 0 9 9 9 2
23 11 13 0 9 2 12 1 10 2 3 13 0 9 1 9 9 2 9 7 3 7 9 2
10 10 9 7 3 13 13 11 7 11 2
17 9 0 9 4 13 11 13 13 15 1 11 3 0 9 0 9 2
25 13 1 15 1 0 9 0 9 1 9 7 9 0 1 9 3 1 0 9 2 13 11 2 11 2
2 0 11
4 11 2 11 2
17 11 11 0 2 1 9 11 11 13 11 11 0 9 9 9 11 2
12 0 13 0 9 1 9 11 1 11 11 11 2
13 11 13 0 9 1 9 7 3 3 13 12 9 2
33 9 9 7 9 9 9 12 1 9 12 11 11 11 13 0 9 1 12 2 1 12 2 9 2 3 7 13 13 1 9 1 9 2
26 15 13 14 1 0 9 7 1 9 13 15 1 0 9 1 0 9 1 11 11 13 1 9 10 9 2
9 11 4 3 13 0 7 11 0 2
8 9 16 11 13 13 10 9 2
12 13 15 9 2 16 1 0 9 13 16 9 2
21 3 13 10 9 1 10 9 7 9 2 13 9 0 11 2 1 15 7 11 13 2
19 13 4 1 15 7 15 13 3 12 9 2 13 15 13 7 7 13 9 2
4 13 0 9 2
11 0 9 1 11 12 13 1 9 11 9 2
20 1 10 0 9 15 13 0 9 9 11 11 13 1 10 9 1 0 0 9 2
18 11 3 13 1 9 11 11 3 0 10 9 7 13 0 9 1 11 2
19 1 9 1 0 9 7 10 9 1 9 11 15 13 9 1 0 0 9 2
8 11 7 13 9 1 0 9 2
15 0 13 2 16 3 9 11 7 11 13 1 11 0 9 2
7 9 12 2 9 12 2 9
18 9 2 12 2 1 15 3 13 11 2 11 2 7 11 2 11 2 2
3 2 11 2
7 1 0 9 3 15 1 0
11 3 9 1 0 9 1 9 1 11 1 11
11 11 2 11 2 11 2 11 2 11 2 2
21 1 12 2 9 0 0 9 2 15 15 13 1 10 9 2 13 15 3 1 0 2
26 9 0 11 3 13 7 13 1 9 9 1 9 9 2 3 0 3 13 7 1 0 9 13 3 0 2
28 3 7 11 1 0 9 3 13 1 0 9 12 1 9 0 9 11 2 16 1 12 2 9 1 15 13 3 2
18 0 0 2 13 1 11 2 7 3 13 9 1 0 9 12 9 11 2
16 3 4 13 1 9 10 9 2 7 16 10 9 4 15 13 2
19 13 0 9 2 16 15 15 1 9 13 13 11 2 13 9 0 9 11 2
16 0 11 9 1 9 13 2 13 0 2 16 13 9 1 15 2
22 13 4 1 15 7 9 9 2 16 11 2 15 3 13 1 10 9 2 4 13 13 2
32 0 11 13 1 11 2 7 16 1 9 9 13 2 3 1 0 9 2 2 9 9 1 0 9 11 7 11 13 10 0 9 2
15 0 9 11 13 9 2 13 4 1 9 13 2 16 13 2
16 1 9 12 2 12 4 7 13 10 0 9 7 3 4 13 2
15 16 4 3 13 3 1 9 0 9 2 13 4 13 3 2
5 7 15 15 13 2
6 11 13 9 14 3 2
17 9 0 2 11 11 13 3 0 2 11 13 1 0 12 9 3 2
20 0 9 3 1 9 4 15 7 13 1 9 7 1 9 4 13 3 15 13 2
34 11 3 3 1 10 9 13 2 3 3 1 9 1 11 7 7 16 3 3 1 0 11 16 0 13 2 13 1 9 14 1 0 9 2
12 9 15 3 13 9 11 2 15 9 3 13 2
19 12 9 13 1 9 2 16 3 15 0 2 0 1 9 2 13 0 9 2
19 0 9 11 13 0 3 1 9 2 13 15 12 9 9 7 9 13 9 2
4 15 13 0 2
26 3 1 9 4 11 13 1 9 2 1 15 13 2 9 4 13 2 14 4 13 2 14 15 13 2 2
10 13 15 10 9 2 13 15 0 9 2
22 15 0 9 11 13 0 9 3 3 2 15 15 1 9 13 16 0 9 1 0 9 2
20 1 9 13 1 0 9 2 3 15 13 0 9 11 2 11 7 11 2 0 2
26 0 9 13 3 1 0 9 9 9 11 2 15 13 1 10 9 1 9 1 0 12 9 1 0 9 2
9 1 11 13 1 9 13 3 9 2
7 1 0 9 4 13 0 2
4 9 0 9 2
15 1 9 15 3 9 1 15 0 13 2 13 0 9 11 2
13 0 9 12 2 9 13 12 0 7 12 0 9 2
28 9 13 1 0 9 9 2 9 2 9 3 3 1 15 2 15 13 2 16 1 0 9 15 13 3 3 3 2
6 1 9 15 13 3 3
12 9 1 9 4 15 13 13 13 9 1 0 9
5 11 11 2 0 11
20 1 9 7 0 9 15 13 9 2 7 3 7 9 9 2 3 13 0 9 2
18 3 2 16 4 15 13 16 0 3 2 16 1 15 13 10 0 9 2
14 14 0 7 13 2 15 7 3 15 13 1 9 13 2
16 13 3 7 9 1 3 0 9 2 0 2 0 7 0 9 2
31 10 9 13 15 0 2 16 13 7 13 9 1 0 0 9 7 10 9 3 13 10 9 2 15 3 13 10 9 7 9 2
17 0 9 13 9 0 9 7 0 9 2 7 16 15 3 3 13 2
14 0 7 0 9 3 13 13 0 1 10 9 7 9 2
23 13 10 9 13 10 9 2 15 1 15 13 0 2 7 14 15 2 1 15 13 0 9 2
23 1 15 4 3 9 13 7 14 3 3 2 9 0 9 13 0 1 9 0 9 7 9 2
9 9 7 0 9 13 9 3 0 2
12 3 7 9 13 2 16 15 10 9 13 3 2
22 10 9 13 1 9 3 3 2 16 10 9 13 3 13 9 2 16 13 3 1 9 2
25 9 3 13 13 15 9 2 3 13 0 13 3 3 7 14 3 2 3 13 15 3 3 0 9 2
13 9 7 13 13 1 9 2 13 15 15 14 9 2
8 9 9 13 1 10 0 9 2
9 9 7 9 15 13 3 3 13 2
9 3 4 15 13 13 10 0 9 2
23 13 3 7 12 9 2 0 9 13 9 10 9 2 16 1 10 9 15 10 14 15 13 2
20 3 3 15 13 13 0 9 7 9 3 1 10 0 9 7 0 9 1 15 2
10 0 9 3 3 13 9 1 0 9 2
22 3 15 13 1 0 9 2 9 7 9 7 3 3 15 15 13 13 9 0 1 9 2
17 1 0 9 15 13 13 3 2 16 4 15 13 1 10 9 3 2
20 0 9 2 3 15 13 1 3 0 9 2 13 9 1 9 9 1 0 9 2
6 2 9 13 9 9 2
12 0 11 2 3 11 11 2 11 11 7 11 11
2 9 9
5 0 11 1 9 11
9 0 9 9 12 1 0 0 9 9
30 11 11 3 13 0 9 1 9 9 1 0 9 7 0 11 15 3 13 1 0 9 1 0 9 1 9 9 1 9 2
23 3 3 13 3 11 11 1 0 9 11 13 11 11 2 11 11 2 11 11 7 11 11 2
7 10 9 3 13 10 9 2
12 12 2 12 2 1 9 2 11 9 9 12 2
25 9 11 11 2 12 2 2 9 11 11 2 12 2 7 9 11 11 2 12 2 13 9 11 12 2
40 1 15 1 3 0 9 2 0 11 2 0 11 2 0 11 2 0 11 7 9 2 11 2 13 3 11 11 2 9 2 2 11 11 7 11 11 2 9 2 2
15 9 12 2 11 13 1 9 10 9 1 0 9 11 11 2
16 15 13 1 9 0 9 0 0 0 11 7 13 15 0 9 2
27 12 2 9 12 2 0 11 13 3 1 0 9 11 1 9 0 11 2 1 15 15 13 0 9 7 9 2
20 12 2 9 12 2 0 11 13 1 9 9 11 11 7 9 7 0 0 9 2
6 9 3 13 1 11 2
20 12 2 2 12 2 9 12 2 0 11 13 9 1 0 9 1 9 0 11 2
11 1 0 9 13 0 11 10 9 2 11 2
12 12 2 9 12 2 0 11 13 1 9 9 2
10 11 15 1 9 1 9 1 9 13 2
18 12 2 9 12 2 13 0 9 0 11 0 9 1 0 9 1 9 2
18 12 2 9 12 2 0 9 1 0 11 13 0 0 9 1 11 11 2
14 12 2 9 12 2 11 11 3 13 0 1 9 13 2
11 11 7 13 0 9 11 11 2 12 2 2
11 12 2 9 12 2 11 11 13 3 9 2
15 12 2 9 12 2 13 0 9 0 11 0 9 1 9 2
8 0 0 9 15 13 11 11 2
5 13 9 1 11 2
17 12 2 9 12 2 0 11 13 1 11 0 9 1 9 0 9 2
12 9 1 10 9 15 3 13 1 0 0 9 2
15 12 2 9 12 2 0 11 13 9 1 9 11 11 11 2
13 13 15 0 9 2 1 15 15 0 11 3 13 2
13 11 3 13 10 9 1 9 11 2 9 1 9 2
19 3 9 13 3 1 9 11 2 12 2 0 9 2 0 11 7 0 11 2
9 12 2 9 12 2 13 9 9 2
5 9 15 13 9 2
15 16 4 13 11 2 13 4 1 0 11 2 13 0 11 2
19 12 2 2 12 2 9 12 2 9 13 9 1 0 9 11 11 0 11 2
10 12 2 12 2 1 0 0 9 1 9
14 12 2 9 12 2 13 0 9 11 11 0 0 9 2
11 11 7 11 15 13 9 7 9 3 13 2
23 12 2 9 12 2 0 11 13 1 0 11 1 11 11 2 15 13 12 9 1 10 9 2
22 12 2 9 12 2 1 9 0 0 9 13 9 0 2 7 9 15 13 1 9 9 2
24 12 2 9 12 2 13 0 9 1 11 2 11 2 11 2 11 2 11 2 0 11 7 11 2
14 12 2 9 12 2 0 11 13 9 10 0 9 9 2
20 12 2 9 12 2 0 11 13 9 9 2 15 15 12 9 13 1 0 9 2
11 12 2 9 12 2 13 9 0 1 9 2
11 13 15 1 9 1 0 0 9 0 11 2
19 12 2 9 12 2 1 0 9 1 11 4 13 9 0 11 3 1 11 2
16 9 12 2 0 9 0 9 0 0 9 1 0 9 1 11 2
5 13 9 0 9 2
20 14 1 0 9 9 2 12 2 15 13 1 12 9 0 9 0 9 1 9 2
30 12 2 9 12 2 13 9 0 0 9 2 15 13 3 9 0 9 0 9 1 0 9 1 9 7 0 9 1 9 2
22 12 2 9 12 2 13 15 9 13 15 13 3 2 15 13 9 0 9 1 0 9 2
16 12 2 9 12 2 0 9 0 9 1 0 9 13 9 9 2
13 9 12 2 0 11 13 13 0 9 1 0 9 2
21 9 12 2 9 0 9 1 0 9 2 9 12 13 0 9 9 1 11 7 11 2
13 12 2 9 12 2 1 9 15 13 9 0 9 2
7 12 2 12 2 9 7 9
23 12 2 9 12 2 0 9 0 11 1 9 0 9 1 0 11 2 15 13 0 9 9 2
14 1 0 9 0 9 1 11 13 0 11 9 1 9 2
14 9 13 0 9 1 9 2 7 7 13 9 7 9 2
6 11 11 1 15 13 2
19 0 11 13 9 9 2 13 9 1 0 9 7 13 9 1 9 7 9 2
16 12 2 9 12 2 13 15 0 9 0 9 1 0 0 9 2
24 12 2 9 12 2 1 0 0 11 15 13 9 9 0 9 11 11 1 11 11 1 9 11 2
7 1 9 3 13 11 11 2
12 9 1 9 9 15 3 13 3 1 0 9 2
16 1 0 9 9 13 14 1 9 9 7 11 11 3 13 9 2
23 9 9 12 2 11 13 0 0 9 1 0 9 0 0 9 2 15 13 12 2 9 12 2
11 9 15 13 0 9 1 9 9 0 11 2
21 9 12 2 11 11 13 9 1 9 7 1 10 9 3 15 13 7 11 1 11 2
12 9 12 7 12 13 1 9 0 9 0 9 2
23 12 2 9 12 2 1 9 15 13 9 1 9 9 0 11 1 9 11 2 11 7 11 2
13 0 9 13 9 2 16 0 0 11 13 0 9 2
12 11 11 13 10 0 9 1 9 9 0 11 2
5 1 9 3 13 2
19 12 2 9 12 2 1 9 13 1 9 3 0 9 0 0 9 1 9 2
6 0 11 0 9 13 2
13 12 2 9 12 2 1 11 13 0 11 0 9 2
21 0 9 9 0 0 9 1 9 15 1 9 12 13 1 9 0 0 9 1 9 2
19 9 12 2 1 11 13 0 11 0 9 2 9 1 0 9 1 11 0 2
9 13 15 1 15 13 12 12 9 2
8 12 2 12 2 0 9 9 2
28 12 2 9 12 2 11 11 13 1 0 9 1 9 2 3 13 0 9 2 0 9 2 0 0 9 0 9 2
19 1 0 15 13 3 2 11 11 2 11 11 2 11 11 2 11 7 11 2
14 9 12 2 11 2 11 7 11 13 13 1 0 9 2
17 12 2 9 12 2 0 11 13 0 9 1 11 11 0 0 9 2
11 9 1 0 9 13 12 2 9 1 11 2
15 12 2 9 12 2 1 9 9 13 0 11 1 0 11 2
5 2 11 2 11 2
3 9 0 11
3 0 9 11
23 0 9 13 1 3 0 0 0 9 1 11 0 9 11 11 9 7 0 9 9 11 11 2
6 0 9 3 13 9 2
14 9 9 13 11 11 1 0 9 0 0 9 11 11 2
13 13 4 0 9 13 2 13 1 9 1 11 11 2
12 13 4 10 9 1 9 2 7 13 15 0 2
14 13 4 1 15 9 1 9 2 15 13 15 1 9 2
10 1 0 9 11 13 0 9 0 9 2
13 11 13 9 2 13 15 9 9 2 15 13 9 2
18 0 9 9 0 15 1 0 9 1 11 13 0 2 7 13 15 9 2
14 13 15 7 9 1 0 9 2 15 4 13 3 0 2
11 13 1 0 9 2 15 4 3 13 9 2
18 9 1 9 2 15 15 13 13 3 2 1 11 2 1 11 2 2 2
10 3 13 9 2 15 15 13 9 9 2
28 16 4 9 15 1 15 13 1 0 11 2 11 15 14 13 2 13 4 1 0 9 2 7 13 15 13 15 2
19 3 1 11 11 4 13 13 9 2 7 3 4 1 9 13 13 0 9 2
16 1 10 9 4 13 10 0 2 0 2 0 9 9 1 9 2
3 2 11 2
7 9 2 1 15 15 9 13
4 11 11 2 11
26 0 0 9 9 0 0 9 7 9 0 9 13 1 0 9 0 9 0 9 2 9 1 11 1 11 2
26 3 15 9 12 13 0 0 9 2 3 1 15 1 9 1 0 0 9 3 1 0 9 13 9 0 2
18 0 9 2 15 4 13 1 11 2 15 13 12 9 1 0 9 9 2
14 1 11 13 9 13 15 1 0 9 1 9 10 9 2
22 1 0 9 1 0 0 9 7 9 13 15 3 0 9 13 2 3 9 13 15 15 2
12 9 9 3 13 3 0 0 9 11 0 9 2
15 1 10 0 9 13 9 11 11 7 11 11 1 0 9 2
29 11 3 1 11 13 0 9 0 9 2 9 11 11 2 11 11 2 11 11 2 7 7 11 11 7 11 11 2 2
32 0 9 11 11 13 0 9 0 9 10 9 2 3 15 13 9 2 9 2 9 1 9 2 9 1 9 2 9 7 9 2 2
15 13 3 3 0 9 10 9 2 16 4 9 13 15 15 2
7 1 0 9 15 3 13 2
17 0 9 15 13 9 0 9 7 0 0 9 9 7 9 0 9 2
17 1 10 9 15 0 9 13 9 9 13 9 9 10 9 1 9 2
18 3 13 1 9 0 9 9 0 9 7 10 9 1 9 0 0 9 2
19 11 11 1 9 1 9 2 15 9 13 1 10 0 9 7 1 9 0 9
2 9 11
3 9 1 11
1 9
28 9 2 0 9 11 11 15 1 9 3 13 0 1 0 9 2 1 10 9 13 0 15 11 2 0 9 11 2
26 1 0 9 7 9 11 11 13 0 9 1 0 9 12 0 9 2 15 13 9 7 9 9 0 9 2
18 9 13 1 0 9 7 13 15 2 16 15 3 3 13 7 1 9 2
18 15 1 3 0 9 3 0 0 11 9 13 14 12 7 12 9 9 2
15 13 3 3 2 16 9 13 2 7 3 3 13 0 9 2
34 9 7 13 1 9 9 3 0 2 7 16 0 9 3 13 1 10 9 3 2 16 15 15 13 7 3 1 10 9 13 3 3 13 2
15 11 1 9 13 2 16 15 1 10 9 14 13 2 2 2
11 13 3 3 2 16 4 15 9 13 3 2
24 0 9 0 9 13 3 1 9 2 1 10 9 0 2 9 11 1 0 9 7 9 1 9 2
29 3 1 11 13 3 0 2 16 3 0 9 13 1 9 15 9 0 9 0 9 2 11 3 3 13 0 0 9 2
24 10 0 9 3 13 0 9 2 9 2 9 2 7 16 7 3 13 3 9 1 10 9 9 2
16 9 11 7 3 3 9 3 0 9 1 11 11 3 13 3 2
19 15 13 3 9 2 15 13 1 9 13 2 7 13 15 3 3 7 3 2
13 0 9 9 13 0 2 11 7 0 7 0 9 2
28 1 15 1 9 11 1 9 13 7 9 10 0 0 9 7 1 0 11 2 0 3 3 2 0 9 7 9 2
18 3 3 9 2 0 1 0 9 3 3 3 2 3 3 13 10 9 2
12 1 10 9 7 1 9 15 13 3 0 9 2
14 3 3 1 0 0 9 2 15 13 11 3 0 9 2
11 7 3 7 1 3 3 0 9 2 2 2
25 15 2 16 1 11 1 9 0 9 9 13 2 13 0 13 1 9 2 9 15 13 14 1 11 2
42 9 2 11 2 6 9 15 2 3 13 7 3 1 15 14 13 9 1 0 9 11 11 2 11 10 0 9 13 2 7 13 7 1 10 9 2 7 15 15 3 13 2
7 11 11 0 9 11 11 2
7 0 9 2 9 11 11 2
9 9 9 2 11 2 12 2 9 2
3 1 0 9
1 9
2 11 11
19 16 15 13 9 3 3 2 16 3 1 11 2 3 13 7 10 0 9 2
16 13 3 1 9 2 7 7 1 9 9 2 3 13 0 9 2
27 12 10 9 15 13 0 7 0 9 2 0 9 7 9 0 9 2 1 11 3 11 2 1 9 1 9 2
32 1 9 9 12 2 15 13 0 7 3 13 4 13 2 13 12 9 9 0 9 7 13 3 0 9 1 0 9 7 0 9 2
19 1 9 13 3 13 7 0 9 13 9 9 2 14 1 12 2 9 2 2
20 9 1 9 9 2 9 2 9 2 0 9 2 9 7 9 15 13 3 3 2
35 11 11 13 0 9 1 9 9 0 9 2 3 15 9 1 9 13 0 9 0 9 2 9 7 9 2 7 3 9 0 9 1 0 9 2
34 11 11 13 0 9 1 0 9 1 9 12 9 2 1 15 13 13 9 1 0 9 2 13 2 14 13 1 0 9 2 14 3 0 2
12 1 9 7 13 2 16 9 0 9 13 13 2
15 11 11 13 0 9 7 10 9 1 0 9 7 1 9 2
31 0 9 7 9 1 0 9 13 11 11 9 12 9 2 12 13 1 0 0 9 2 12 13 13 3 2 12 13 0 3 2
9 11 11 15 1 12 9 13 9 2
16 1 0 7 0 9 13 3 9 9 1 9 7 3 1 9 2
9 11 11 13 1 9 0 9 3 2
18 1 10 9 13 9 0 15 3 3 2 1 9 2 1 9 7 9 2
12 1 0 9 13 9 1 9 1 10 0 9 2
18 13 15 3 2 7 3 13 0 9 9 2 15 13 1 9 1 9 2
9 9 9 13 1 9 0 0 9 2
19 9 11 13 13 3 9 1 0 9 2 11 13 9 9 3 1 0 9 2
17 0 9 3 13 2 0 9 2 0 9 2 0 9 3 2 2 2
31 3 4 3 0 9 2 15 0 0 9 13 2 13 1 15 13 15 2 16 0 9 10 9 13 1 9 7 9 0 9 2
4 0 9 0 9
16 0 9 11 2 15 13 1 0 9 11 11 2 13 11 11 2
17 9 9 13 1 9 12 2 1 9 0 9 15 13 7 9 9 2
19 16 4 13 1 9 2 3 4 13 10 0 7 0 9 2 13 11 11 2
24 10 9 13 13 9 2 15 13 9 2 16 15 4 13 9 9 2 13 9 9 1 0 9 2
18 7 13 1 9 0 2 0 9 13 3 13 2 13 15 15 3 13 2
23 11 11 2 9 9 1 9 7 9 1 0 9 0 9 2 12 2 2 13 0 0 9 2
31 3 1 9 9 13 0 9 7 0 9 1 0 0 0 9 1 0 11 2 1 12 9 3 15 13 9 0 9 1 11 2
25 13 9 0 9 0 2 9 1 11 2 12 2 12 2 2 3 14 1 9 12 13 0 0 9 2
19 1 9 12 15 13 9 0 9 1 11 2 3 1 10 9 13 16 9 2
16 0 9 0 9 2 15 3 13 2 13 1 10 9 3 0 2
17 13 1 15 10 0 9 7 7 3 0 9 2 16 13 9 11 2
24 13 7 3 0 2 3 0 7 3 3 0 2 16 3 13 9 2 15 13 15 9 0 9 2
16 3 3 1 0 9 13 12 0 9 2 11 2 0 7 11 2
15 9 0 9 9 13 1 11 11 9 0 9 1 0 9 2
19 1 9 3 1 10 9 13 10 0 9 3 1 11 2 7 3 1 11 2
31 0 3 13 7 9 0 9 0 9 9 9 2 9 2 11 11 11 7 10 9 0 9 11 11 1 9 9 9 11 11 2
8 0 9 13 10 9 1 9 2
12 9 9 0 9 4 13 4 13 1 0 9 2
17 9 13 16 0 9 0 7 0 12 2 9 7 0 9 10 9 2
7 13 3 0 0 9 0 2
23 9 13 0 0 9 1 10 0 9 2 7 9 9 4 13 9 1 9 7 1 10 9 2
3 2 11 2
4 9 13 7 11
15 9 9 9 1 0 9 15 13 12 2 9 7 13 3 0
2 11 11
13 13 1 0 9 1 9 10 9 4 3 13 0 2
18 13 3 3 1 0 9 9 9 2 7 15 14 1 12 9 2 9 2
18 9 13 7 3 3 0 0 9 2 16 1 9 13 0 13 1 9 2
29 9 9 9 2 1 9 1 0 9 1 3 12 9 2 4 13 7 9 0 9 9 12 1 12 5 1 12 9 2
37 1 9 0 9 3 13 9 1 0 9 2 7 9 9 13 3 3 0 2 16 15 13 9 12 9 2 15 1 9 0 9 13 14 0 12 5 2
22 12 9 1 0 9 3 13 13 9 9 3 2 3 3 2 16 1 15 13 9 11 2
16 1 0 9 15 13 0 9 2 9 0 0 9 2 11 2 2
17 13 3 1 9 9 1 12 5 1 12 9 1 3 0 0 12 2
23 10 9 15 13 3 12 5 9 10 9 0 9 7 1 9 9 7 9 12 7 12 5 2
25 13 15 15 3 3 2 1 0 2 9 2 11 7 11 2 10 9 3 13 14 1 9 12 9 2
23 9 0 9 3 3 13 4 2 16 13 0 9 2 3 13 1 9 9 1 0 0 9 2
16 3 13 0 2 3 15 1 9 13 7 15 10 0 9 13 2
24 0 9 2 10 9 13 9 13 16 9 2 1 10 9 15 13 13 2 15 13 1 12 9 2
21 3 3 13 0 9 9 2 13 3 9 3 0 7 0 9 13 3 9 9 9 2
22 9 13 9 0 9 0 1 12 9 7 13 15 3 7 11 1 9 12 9 2 9 2
11 1 9 13 0 9 11 1 9 12 9 2
7 12 9 15 3 13 1 0
2 11 11
19 0 9 0 9 0 2 11 2 15 9 0 9 13 11 11 2 12 2 2
21 1 9 1 9 0 9 13 1 11 11 7 1 0 9 11 2 0 11 11 2 2
8 1 10 9 4 13 1 9 2
11 10 9 13 3 0 9 10 9 11 11 2
13 0 9 13 1 0 9 9 0 9 1 0 9 2
26 9 4 1 9 15 13 1 3 0 0 9 2 3 1 9 0 9 2 0 1 9 0 1 0 11 2
9 1 0 9 13 3 7 0 9 2
5 2 15 13 9 2
4 13 0 9 2
15 9 0 9 13 13 0 9 2 15 0 4 13 13 9 2
13 1 15 3 13 0 9 2 15 4 15 13 13 2
25 1 0 9 4 15 1 9 13 13 12 0 9 2 7 14 0 12 7 12 9 16 1 0 9 2
23 0 9 4 15 9 13 13 7 0 9 2 13 0 9 2 3 13 7 1 9 7 3 2
15 2 9 9 11 4 7 13 13 7 1 15 0 2 2 2
11 15 13 3 15 2 15 3 15 3 13 2
26 13 3 3 2 15 15 13 2 7 13 13 15 2 15 15 13 2 1 0 9 7 9 2 0 9 2
25 4 13 0 0 9 2 7 15 7 1 9 2 16 1 0 9 13 0 9 10 12 9 3 0 2
26 3 3 13 4 15 13 13 0 9 2 13 15 7 13 1 15 2 15 10 9 1 0 1 15 13 2
9 13 15 9 1 0 9 7 9 2
43 13 4 15 1 15 13 7 3 0 9 11 2 15 13 10 0 9 2 7 13 4 15 13 2 3 16 1 0 9 2 0 9 2 1 0 9 0 0 9 0 9 2 2
10 1 10 9 4 13 9 1 0 9 2
37 15 9 15 13 13 0 9 1 0 9 2 1 15 2 16 4 13 13 0 9 2 15 15 4 1 0 9 13 7 15 4 15 3 14 13 13 2
12 13 3 1 0 9 2 15 7 13 0 9 2
23 3 15 3 13 0 0 9 2 16 1 3 0 7 0 9 1 9 13 9 1 9 2 2
18 11 13 3 3 1 0 9 0 9 2 15 13 1 9 12 2 2 2
23 13 15 2 16 1 9 12 3 3 13 0 9 7 16 15 3 9 9 13 13 3 3 2
23 15 2 16 1 10 9 13 9 2 4 13 13 14 16 9 9 2 7 16 9 9 2 2
16 0 9 11 15 14 13 13 9 1 9 12 11 11 2 2 2
22 1 9 9 4 13 0 9 2 3 4 15 1 15 13 2 7 15 4 15 13 3 2
20 9 11 13 9 9 2 15 4 13 9 2 9 4 13 3 1 9 9 9 2
9 10 0 9 1 15 7 3 13 2
3 11 0 9
8 0 9 1 9 0 9 2 12
7 11 1 11 2 11 2 2
25 3 0 9 1 9 0 9 2 12 13 0 9 11 11 1 15 2 16 15 13 9 9 11 12 2
25 15 4 13 16 9 1 9 9 2 15 15 3 3 13 1 0 9 7 0 0 9 1 0 9 2
23 11 15 3 0 9 2 12 9 2 13 9 7 3 10 9 4 13 1 0 0 9 9 2
37 9 2 16 1 0 9 0 1 12 9 1 12 2 13 11 11 2 11 11 2 11 11 7 11 11 2 2 7 0 9 7 9 9 13 1 9 2
12 7 7 13 1 9 12 9 0 9 1 11 2
17 1 0 9 15 13 11 11 1 12 7 1 0 11 11 1 12 2
20 11 11 13 3 12 0 9 1 12 9 7 1 0 9 13 9 1 0 12 2
22 3 1 9 13 2 13 2 16 15 15 13 10 0 9 2 13 0 16 1 0 9 2
28 1 0 9 3 1 9 1 9 1 0 9 13 2 13 15 10 0 0 9 7 3 1 9 4 15 0 13 2
13 1 0 9 13 13 7 3 7 3 3 3 13 2
8 11 1 9 2 1 9 7 9
2 11 2
38 0 9 11 1 11 15 3 2 16 1 9 9 1 12 9 0 9 1 9 1 11 13 14 1 0 9 9 11 2 13 1 0 9 7 13 0 9 2
14 9 12 2 12 13 1 12 12 9 0 9 9 11 2
33 1 11 2 15 1 9 13 14 0 7 1 9 15 7 3 13 2 13 1 9 10 9 11 2 1 9 0 2 2 15 9 13 2
23 0 9 13 1 0 9 1 12 9 2 3 11 11 9 12 2 12 13 0 9 11 11 2
3 11 13 9
2 11 2
11 0 0 9 0 9 11 11 11 13 9 2
30 10 9 11 15 13 1 9 1 11 1 0 9 11 7 11 11 2 15 4 13 1 0 0 9 11 2 13 9 0 2
5 9 13 12 9 2
7 9 13 3 0 9 11 2
3 1 0 9
13 9 0 0 9 11 11 13 9 0 9 11 11 2
5 9 13 0 9 2
29 11 11 2 9 0 0 9 11 2 13 1 9 1 0 0 9 2 1 15 10 9 13 1 11 11 12 2 12 2
4 9 13 1 9
7 11 2 11 2 11 2 2
14 1 0 0 9 15 3 1 11 1 0 9 13 9 2
18 1 9 15 9 13 13 15 9 1 9 1 9 7 13 1 15 9 2
19 1 0 2 15 13 9 1 9 2 13 11 2 15 13 1 12 9 11 2
20 13 15 2 7 13 9 2 13 4 15 1 9 2 13 2 13 14 1 9 2
21 1 9 13 2 0 9 4 3 13 2 7 9 4 13 3 2 3 4 13 9 2
11 3 13 0 2 16 15 13 1 0 9 2
7 1 9 11 13 9 11 2
14 9 15 13 2 16 4 16 0 9 13 1 0 9 2
13 1 9 4 12 9 13 2 1 9 3 1 9 2
9 3 15 11 13 1 9 2 2 2
12 3 3 4 13 3 10 9 2 13 9 11 2
14 1 9 4 13 13 2 16 1 9 13 9 1 9 2
11 13 15 3 3 2 3 15 15 13 13 2
15 3 2 16 15 9 13 1 9 2 9 13 1 0 9 2
11 1 9 4 13 2 16 4 13 10 9 2
4 9 13 0 2
12 13 7 3 9 13 1 9 2 13 15 11 2
28 10 0 9 11 14 13 2 13 15 9 1 12 9 2 11 13 0 9 1 15 9 2 13 15 15 15 9 2
8 1 9 13 7 9 11 11 2
18 3 13 1 9 11 2 11 2 3 13 13 9 11 9 11 7 11 2
10 3 15 15 4 13 1 9 10 9 2
8 11 2 3 2 13 11 2 11
2 9 11
6 11 13 2 11 13 9
19 0 9 1 0 9 9 2 0 9 2 11 12 2 12 2 12 2 12 2
9 11 2 11 2 11 2 11 2 2
22 7 1 9 15 9 0 0 9 13 1 15 2 3 3 13 10 9 1 9 9 11 2
12 1 0 9 13 1 0 11 11 12 2 12 2
24 3 13 0 9 15 13 3 1 12 2 9 11 2 13 15 1 9 2 3 15 9 13 11 2
10 1 9 15 11 13 2 12 2 12 2
16 0 9 2 15 3 13 1 11 2 15 13 9 13 1 9 2
18 9 15 13 14 1 0 9 9 2 16 15 13 14 1 12 9 9 2
13 1 12 2 9 13 11 2 16 15 13 0 9 2
13 3 13 9 1 9 7 0 11 15 1 9 13 2
11 9 15 13 1 0 9 14 1 12 9 2
13 1 9 13 11 2 13 7 11 13 9 3 3 2
8 7 15 7 13 9 0 9 2
23 3 15 9 13 9 1 12 2 9 2 7 13 2 16 1 0 9 15 13 14 0 9 2
23 15 3 13 11 1 9 9 2 13 15 3 9 9 7 0 9 15 13 1 3 0 9 2
36 1 0 9 9 15 13 7 10 0 9 7 1 12 2 9 3 1 15 13 9 2 0 9 14 3 13 2 3 9 1 0 9 13 1 9 2
17 1 9 7 0 9 13 9 7 1 0 0 0 9 2 1 9 2
14 13 15 11 7 11 13 10 0 9 2 12 2 12 2
10 7 1 0 9 13 0 9 1 9 2
9 11 13 9 11 2 15 9 13 2
11 3 15 0 9 13 7 15 1 0 9 2
26 1 12 2 9 13 1 0 9 11 2 3 11 13 9 9 16 0 9 2 7 0 9 9 11 13 2
12 9 9 3 13 1 9 2 16 1 15 13 2
11 1 10 9 1 12 2 9 3 13 11 2
16 0 9 13 3 1 9 13 11 2 16 4 10 9 13 11 2
16 7 3 11 3 13 9 2 10 0 0 9 13 11 1 9 2
17 11 3 13 1 0 9 0 9 2 7 9 3 10 9 3 13 2
22 11 15 13 1 0 0 9 2 13 7 3 3 0 11 2 15 15 13 0 0 9 2
14 0 9 13 0 11 1 12 9 9 1 9 0 9 2
4 11 13 0 9
15 0 0 9 2 11 2 13 3 0 9 0 9 1 11 2
19 0 9 1 0 9 12 5 4 13 12 2 9 1 0 9 12 9 9 2
13 9 13 1 9 7 10 0 9 13 12 12 9 2
29 3 4 13 1 9 0 9 11 2 12 2 9 1 9 0 0 9 2 7 9 9 4 15 13 13 1 0 9 2
19 11 3 13 3 0 9 0 9 2 15 15 1 0 9 13 12 2 9 2
18 13 15 0 0 9 0 9 12 5 1 0 9 12 7 12 12 9 2
12 1 9 13 1 12 2 9 1 15 9 11 2
12 11 13 0 9 10 9 9 3 1 9 9 2
7 13 0 7 13 1 9 2
23 0 9 4 13 3 2 15 13 2 16 10 0 9 13 1 0 9 0 16 0 9 9 2
8 9 4 13 1 9 12 5 2
14 0 9 12 9 13 13 0 9 11 7 10 0 9 2
28 1 12 2 9 12 11 13 0 9 9 2 15 15 13 9 9 1 12 9 2 9 9 0 9 1 12 9 2
28 9 0 9 13 1 9 0 9 1 9 1 9 0 9 1 12 7 12 5 0 7 3 13 12 9 2 9 2
16 9 1 0 9 13 1 3 16 12 5 7 13 12 9 9 2
34 9 1 0 9 13 9 10 9 1 9 1 3 0 9 2 3 1 0 9 2 1 15 13 0 9 1 0 0 9 1 9 1 9 2
11 1 0 9 13 14 1 9 1 0 9 2
37 3 13 1 9 9 7 9 0 9 2 1 0 9 0 9 2 15 13 9 1 0 9 2 15 9 13 9 1 9 9 0 9 2 7 0 9 2
14 0 9 1 0 9 9 13 9 1 0 7 0 9 2
24 10 9 1 9 1 0 9 13 1 12 5 1 0 0 9 1 12 5 1 12 2 9 12 2
3 2 11 2
6 11 13 1 9 0 0
13 1 9 1 0 11 3 13 0 9 0 0 11 11
8 0 9 11 1 0 11 11 11
14 0 9 11 11 2 12 2 2 13 1 9 0 0 2
40 0 9 1 11 13 1 12 2 9 11 11 2 12 2 2 1 12 9 7 12 9 12 2 12 2 12 2 12 2 12 2 12 2 12 2 2 12 2 12 2
23 1 12 0 9 15 11 13 1 0 9 0 7 1 0 13 12 0 9 1 12 2 12 2
11 11 10 9 13 7 3 3 13 9 11 2
33 0 9 7 13 1 10 0 0 9 2 0 1 0 11 2 3 1 0 0 12 7 12 2 7 13 1 15 9 9 11 2 11 2
26 1 9 3 13 0 9 0 0 9 2 7 15 11 2 11 2 12 2 2 2 11 2 12 2 2 2
52 9 9 13 1 0 11 1 9 3 2 3 13 1 0 9 0 0 11 11 2 12 2 2 2 15 13 1 12 2 9 1 11 11 2 12 2 2 12 2 12 2 12 2 12 2 12 2 2 12 2 12 2
46 3 0 0 9 13 11 2 11 2 12 2 2 7 11 2 12 2 2 2 11 2 12 2 2 2 0 2 12 2 2 9 13 1 9 11 2 12 2 2 2 11 2 12 2 2 2
25 1 9 0 9 1 15 13 0 2 0 9 11 2 11 7 0 2 0 9 11 2 11 2 11 2
14 1 12 0 9 15 11 1 11 12 13 1 0 9 2
39 16 9 1 0 9 15 13 13 7 1 0 9 2 9 1 0 9 2 2 3 0 11 15 3 9 13 2 7 1 0 0 9 13 10 0 9 3 13 2
10 1 0 0 15 7 3 13 1 9 2
24 7 4 1 10 9 13 3 16 1 9 2 16 13 0 2 13 11 3 2 16 13 0 9 2
30 1 9 1 10 9 11 13 1 9 2 13 1 15 13 1 9 2 7 1 9 2 3 1 15 13 9 12 2 12 2
17 3 4 3 13 2 16 15 13 12 7 13 1 15 1 12 9 2
19 11 3 1 15 13 7 13 2 2 13 4 12 1 0 9 9 2 2 2
11 13 4 15 7 6 2 3 4 15 13 2
17 1 0 9 15 13 7 9 0 11 1 0 11 2 12 2 2 2
16 3 4 15 13 2 15 15 13 12 7 11 13 1 15 3 2
66 3 15 3 13 9 2 13 0 1 3 7 1 9 13 9 2 7 9 13 3 16 9 2 13 15 11 2 15 9 1 0 11 12 2 12 2 12 2 12 2 12 2 12 2 12 2 12 2 12 2 12 13 1 0 9 2 9 13 3 2 16 15 15 13 9 2
37 14 1 15 13 2 16 3 3 13 0 9 2 13 15 0 9 9 0 0 12 2 7 1 9 13 1 15 0 9 0 7 4 7 13 0 9 2
23 11 15 1 0 0 0 13 13 10 0 9 2 9 11 11 2 16 13 0 16 10 9 2
25 11 11 13 1 9 0 9 3 3 1 0 11 1 9 12 2 11 15 15 13 1 12 9 3 2
34 1 12 9 15 9 13 13 2 13 11 2 12 2 2 3 2 16 13 1 0 0 9 9 11 1 9 12 2 12 2 12 2 12 2
19 13 15 1 3 0 9 2 7 12 9 13 1 9 1 9 9 0 9 2
31 1 9 9 15 1 9 13 0 9 0 9 2 13 2 15 15 13 2 7 13 13 9 2 3 13 0 9 2 0 11 2
23 11 2 11 15 1 11 13 9 1 0 0 0 2 1 0 9 13 0 9 12 2 12 2
22 15 3 1 0 11 1 12 9 13 2 7 3 13 7 0 12 9 13 3 1 9 2
40 9 1 0 0 9 2 0 11 11 2 12 2 2 13 3 2 0 9 13 9 14 1 0 9 2 7 15 0 9 2 3 13 12 2 12 2 12 2 12 2
23 11 2 11 3 13 1 11 11 2 12 2 2 9 9 2 12 2 12 2 12 2 12 2
2 0 9
7 10 9 3 13 1 9 2
4 13 11 3 2
5 11 2 11 2 2
17 3 10 9 15 1 11 13 12 2 9 0 9 11 1 0 9 2
25 1 12 9 15 13 9 13 1 0 9 9 2 16 1 9 4 13 9 1 9 9 0 9 9 2
41 0 9 11 11 13 1 11 3 1 12 0 9 2 11 11 11 2 12 11 13 0 9 0 11 2 13 0 9 0 9 7 11 11 11 13 3 0 9 0 9 2
18 7 0 9 13 9 9 2 11 11 7 11 2 11 11 7 0 11 11
31 1 0 9 4 13 15 11 2 15 10 9 13 0 9 2 7 0 9 9 11 11 1 11 2 15 13 9 3 1 11 2
40 1 0 9 13 0 9 1 0 11 2 15 3 4 13 1 11 1 9 1 11 2 7 1 9 0 11 15 13 1 10 0 9 2 7 9 15 13 3 13 2
16 13 7 0 11 7 11 2 15 13 1 0 9 9 1 11 2
11 0 0 9 11 13 1 9 0 9 9 2
6 9 13 13 9 1 9
7 11 2 11 2 11 2 2
14 1 12 12 9 3 13 0 0 9 9 1 9 9 2
30 15 4 1 9 12 1 9 1 0 12 9 13 0 0 9 13 9 1 12 9 7 13 9 0 9 2 9 7 9 2
28 9 1 9 2 1 10 9 15 10 9 13 2 15 4 13 3 2 3 2 11 7 11 15 13 9 1 9 2
25 9 11 1 0 11 11 11 3 13 2 16 1 9 11 4 9 1 10 9 13 0 0 9 9 2
9 0 1 15 13 3 9 1 11 2
7 0 9 4 9 13 3 2
19 9 10 9 13 13 9 1 9 7 1 9 2 13 0 9 11 11 11 2
10 11 13 2 11 1 15 13 3 0 9
5 11 2 11 2 2
19 0 0 9 11 2 11 15 1 0 9 13 3 1 3 0 9 1 11 2
8 11 3 0 9 13 9 9 2
33 0 9 0 9 11 12 3 3 1 0 0 9 13 3 0 9 7 13 3 9 0 9 11 11 2 15 3 13 1 0 9 9 2
23 9 0 11 15 3 13 1 9 0 0 9 1 9 1 9 2 1 15 9 9 9 13 2
14 13 3 14 9 0 9 11 2 15 15 9 13 3 2
47 1 9 1 12 9 9 9 2 3 1 12 9 13 1 0 3 0 0 0 9 2 15 3 3 3 3 13 7 3 15 13 14 1 0 9 2 7 3 3 0 9 3 3 13 9 9 2
15 0 9 13 3 1 12 9 3 2 13 15 12 1 9 2
16 3 13 2 16 11 13 3 1 9 2 13 9 0 11 11 2
14 9 13 0 9 1 9 12 9 9 1 9 0 9 2
17 9 9 11 11 15 13 13 2 16 1 10 9 13 9 7 0 2
25 9 14 13 2 16 7 0 9 11 13 13 2 13 11 2 15 1 0 9 13 3 10 9 13 2
13 13 4 16 9 0 9 7 10 9 13 1 9 2
17 16 0 2 9 1 0 11 7 9 1 9 0 9 11 3 13 2
35 9 0 9 11 11 12 9 2 11 13 2 16 1 9 12 0 9 2 9 9 3 2 2 3 15 13 9 0 0 9 7 9 1 9 2
10 15 15 1 0 9 4 13 0 9 2
11 1 9 9 13 13 0 9 2 13 11 2
17 0 9 11 13 2 16 0 9 0 9 15 4 13 3 1 9 2
6 10 9 13 11 9 2
12 10 0 9 11 11 15 13 1 9 0 9 11
16 1 9 10 0 9 11 11 13 1 0 11 0 9 11 11 2
26 11 3 13 0 0 1 9 1 11 11 2 11 7 1 9 1 11 11 2 15 15 3 13 1 9 2
25 1 10 9 3 13 1 0 9 11 1 0 9 9 1 9 2 9 1 9 7 9 1 0 9 2
19 13 4 1 9 13 15 9 7 16 11 13 0 11 2 13 4 15 3 2
17 3 15 15 1 15 9 13 2 16 13 0 2 13 0 9 11 2
10 9 1 9 0 9 3 13 0 9 2
30 7 16 1 0 11 3 13 0 9 0 9 11 7 11 2 0 9 1 11 11 11 15 13 1 9 13 0 9 11 2
8 1 9 10 9 13 0 9 2
32 9 9 11 11 2 11 11 3 10 9 2 9 11 11 2 13 9 9 10 9 2 0 9 9 11 11 7 0 9 0 11 2
28 0 11 15 3 13 1 9 0 9 2 0 0 13 1 11 11 2 2 15 13 9 2 16 9 10 9 13 2
21 0 0 3 2 13 1 9 0 9 7 9 2 14 9 1 9 15 0 9 13 2
9 13 15 9 1 9 13 1 11 2
52 16 4 15 1 9 15 13 2 16 4 1 9 13 2 13 4 15 2 13 11 2 15 1 9 11 3 13 2 3 2 9 1 0 9 3 13 1 10 9 1 9 2 2 7 16 3 13 10 9 3 0 2
13 9 1 0 11 13 7 11 11 2 10 0 9 2
18 14 16 4 3 13 2 16 15 13 1 9 2 7 15 15 9 13 2
18 11 13 9 2 15 3 13 9 1 10 9 2 16 3 0 7 0 2
15 3 15 13 9 2 3 13 10 0 9 2 14 3 15 2
12 0 9 15 1 10 9 7 13 7 11 11 2
31 3 2 16 15 3 13 2 13 1 9 1 9 10 9 7 13 15 1 0 9 2 15 3 11 13 2 7 11 13 9 2
27 1 9 2 16 1 15 13 1 11 2 11 10 0 9 1 9 0 0 11 13 7 3 13 1 9 11 2
13 13 15 2 13 7 10 9 15 15 13 1 9 2
22 1 0 0 15 13 14 3 2 16 15 11 11 1 9 13 2 16 15 13 1 11 2
23 15 15 15 13 2 13 7 13 15 3 16 3 2 13 0 11 1 9 11 10 0 9 2
22 1 0 0 0 9 13 1 12 9 0 2 3 15 7 1 11 13 9 0 0 9 2
26 12 3 1 0 9 13 9 1 9 2 11 13 9 0 0 12 7 9 12 2 11 0 0 12 2 2
33 0 9 13 1 12 0 9 2 15 2 15 1 15 13 2 15 4 13 13 1 9 1 9 12 9 2 9 15 13 3 1 9 2
15 1 9 15 13 11 1 9 13 9 0 0 9 1 11 2
15 16 4 1 9 13 9 9 7 0 2 15 13 0 9 2
3 2 11 2
2 0 11
3 3 1 9
9 9 11 4 13 13 1 9 0 9
4 9 9 0 9
5 11 2 11 2 2
33 10 0 9 13 0 2 13 15 1 9 7 13 1 12 2 9 3 15 0 9 2 13 11 11 2 9 9 0 9 9 11 11 2
39 1 9 2 15 13 3 9 12 2 11 2 13 0 0 2 9 11 2 12 2 0 9 2 7 3 1 9 15 13 11 2 11 2 7 11 2 11 2 2
14 9 11 7 11 13 3 2 3 15 1 10 9 13 2
21 12 9 15 3 13 1 15 9 7 1 0 9 13 10 9 1 0 9 7 13 2
16 15 9 15 13 2 16 15 15 1 15 13 2 13 9 11 2
35 9 0 9 4 13 13 9 11 11 2 1 9 2 2 15 1 9 1 11 13 11 3 3 1 0 9 7 13 9 1 12 5 12 9 2
28 9 13 11 11 2 11 2 2 11 11 2 11 2 2 11 2 0 2 11 2 7 11 2 0 2 11 2 2
24 1 15 11 11 2 13 4 3 1 10 0 9 2 7 13 13 1 9 15 14 1 10 9 2
9 3 4 13 9 1 10 0 9 2
31 1 0 9 13 0 14 12 9 2 7 9 11 15 13 2 16 4 13 1 9 1 9 9 16 3 11 11 7 0 11 2
16 1 0 9 3 4 15 3 13 3 13 2 16 3 13 13 2
10 10 9 4 13 13 7 0 0 9 2
17 7 13 9 9 12 9 7 12 9 1 9 3 4 13 12 9 2
18 0 9 13 9 11 2 7 13 1 15 2 16 9 13 13 10 9 2
17 0 3 13 1 9 1 9 9 11 1 0 9 2 0 9 9 2
8 1 0 9 9 15 13 13 2
27 1 0 9 4 3 13 1 9 13 9 10 9 2 16 15 13 0 2 15 13 3 9 2 13 11 11 2
10 9 9 9 0 9 11 2 11 7 11
16 1 0 9 13 13 1 12 12 9 1 9 1 9 0 9 2
9 1 15 13 1 9 0 14 12 2
23 0 0 9 13 9 0 9 11 2 11 7 11 2 11 11 2 2 15 13 3 12 9 2
48 9 13 1 10 9 0 9 2 16 13 9 7 0 9 2 0 9 1 0 9 7 10 9 2 3 2 0 9 9 13 12 2 12 9 1 0 9 2 2 7 3 9 9 7 9 0 9 2
10 13 0 9 9 2 15 15 9 13 2
13 0 9 11 13 7 13 9 9 1 12 2 9 2
4 0 9 15 13
12 3 0 0 9 1 9 1 0 9 12 1 11
2 11 2
16 1 12 9 15 3 13 9 1 0 9 1 11 1 0 9 2
20 9 9 13 1 9 1 9 9 3 13 7 11 13 1 9 0 9 1 11 2
22 7 1 0 9 4 15 13 13 7 0 9 0 9 7 1 0 9 9 11 11 11 2
18 1 9 0 9 4 0 9 13 1 0 9 0 9 1 11 7 11 2
26 0 9 11 13 1 9 1 11 1 9 9 1 9 2 1 15 7 3 13 9 11 2 15 13 9 2
25 1 0 9 0 9 13 2 1 0 9 15 13 14 9 1 9 0 9 11 1 0 9 11 11 2
22 3 1 12 9 4 3 1 10 9 1 11 13 11 11 2 15 13 1 9 16 9 2
40 1 0 9 11 15 1 9 13 0 9 2 11 2 11 2 11 7 11 2 11 13 1 9 9 2 1 9 13 14 3 0 1 11 2 7 7 11 7 11 2
12 3 4 1 9 9 11 13 13 11 0 9 2
31 11 4 1 9 1 11 1 11 13 9 9 11 2 15 13 3 0 9 2 7 13 13 7 9 11 2 15 13 9 9 2
19 10 9 9 13 9 1 11 2 15 15 1 12 9 13 0 9 1 11 2
21 9 1 11 13 9 1 9 11 2 7 7 15 0 11 13 1 9 1 9 11 2
12 0 9 4 13 7 11 1 0 9 1 11 2
22 1 9 11 13 9 1 11 0 9 2 3 13 7 11 2 15 4 10 9 13 13 2
8 1 12 9 13 3 9 11 2
17 9 9 0 11 15 3 13 13 7 10 9 1 9 3 3 13 2
28 1 0 9 1 9 7 4 1 0 11 13 14 0 9 11 2 15 9 4 13 13 0 9 1 11 11 11 2
7 7 11 13 1 11 0 2
20 9 1 9 11 15 1 0 0 9 13 9 7 1 9 4 13 11 1 11 2
17 0 9 9 1 9 2 9 12 2 11 2 11 2 11 2 11 2
15 9 12 2 11 2 11 2 11 2 11 2 11 2 11 2
11 9 12 2 11 2 11 2 11 2 11 2
11 9 12 2 11 2 11 2 11 2 11 2
11 9 12 2 11 2 11 2 11 2 11 2
12 11 11 2 3 2 13 1 0 9 2 2 2
14 9 0 9 0 11 13 1 11 3 3 9 1 11 2
8 13 13 1 12 9 9 11 2
17 1 0 9 15 3 13 1 9 1 0 9 11 9 11 2 11 2
10 0 0 9 0 11 13 1 9 13 2
17 9 12 12 9 15 3 4 13 3 1 12 9 2 3 1 9 2
5 9 11 11 2 11
5 0 9 13 3 9
5 11 2 11 2 2
28 0 9 13 9 9 0 3 0 9 3 13 1 0 9 9 1 10 9 9 9 0 0 7 0 9 11 11 2
31 13 3 3 1 9 11 1 9 9 10 9 1 9 9 9 11 11 2 9 9 11 11 2 9 0 9 7 0 0 9 2
58 9 0 9 11 11 1 9 13 2 16 1 9 9 2 10 0 9 13 2 0 9 3 13 13 9 3 0 0 0 9 2 7 13 3 1 15 2 16 4 10 9 1 9 13 13 9 0 9 7 3 13 1 9 0 7 0 9 2
12 10 9 10 9 15 13 10 9 2 13 11 2
21 9 2 16 0 9 9 4 13 1 9 0 9 9 2 13 9 0 9 10 9 2
13 9 9 11 11 2 11 2 13 0 9 1 0 2
7 0 9 9 13 9 1 9
5 11 2 11 2 2
21 9 2 15 0 0 9 2 0 2 9 2 11 2 13 1 10 9 2 13 0 2
29 0 9 9 11 2 11 7 9 11 2 11 13 9 1 9 1 0 9 2 15 13 13 9 0 9 1 9 9 2
22 9 0 2 9 2 11 13 1 9 1 0 9 2 15 9 13 1 12 0 2 9 2
18 0 9 1 11 7 0 2 9 2 11 13 13 0 9 1 15 0 2
15 11 2 11 7 13 9 1 0 9 2 15 10 9 13 2
19 9 13 3 11 1 11 2 16 15 15 13 2 16 9 9 1 9 13 2
25 15 11 1 0 9 13 2 9 7 3 13 0 2 9 2 11 2 7 12 9 2 3 13 11 2
11 15 13 2 16 4 9 0 9 3 13 2
22 16 0 2 9 2 11 9 13 2 11 13 0 9 1 11 2 16 4 9 13 13 2
22 3 9 13 0 2 9 2 11 2 0 9 2 3 13 9 2 1 12 9 2 9 2
14 9 1 9 13 1 9 2 16 9 13 13 1 9 2
16 9 9 7 13 0 9 1 15 2 16 9 3 4 13 13 2
34 13 3 2 16 15 15 13 1 9 0 2 9 2 11 2 2 16 9 13 1 9 13 0 9 1 15 2 15 15 13 0 9 13 2
17 9 11 1 9 9 0 2 9 2 11 13 11 2 11 1 0 2
5 9 1 9 14 13
16 1 9 1 9 11 15 13 12 9 2 1 9 9 11 12 9
5 11 2 11 2 2
32 14 9 9 1 9 0 9 0 9 13 1 12 2 9 12 2 3 1 12 7 9 9 1 9 11 2 3 0 9 9 9 2
7 13 15 10 9 11 11 2
22 9 1 15 13 15 1 9 9 1 0 9 2 3 0 0 9 1 11 7 0 9 2
8 1 0 9 15 13 0 9 2
25 16 11 13 0 9 2 1 12 2 9 15 3 13 9 1 9 1 9 11 1 12 9 1 9 2
20 1 9 2 16 0 9 13 1 11 10 9 7 9 2 13 9 13 0 9 2
24 1 9 11 11 0 9 2 3 11 2 13 9 13 7 9 15 14 13 1 0 9 1 11 2
15 1 9 1 9 9 7 13 9 1 0 9 1 9 9 2
13 9 1 9 0 9 13 7 1 0 9 12 9 2
31 0 7 0 9 1 9 9 0 9 13 9 0 9 7 9 2 11 2 1 9 0 0 9 2 15 13 9 1 0 9 2
12 1 3 0 11 1 11 13 1 9 9 9 2
12 0 15 1 11 11 1 11 13 1 0 9 2
26 0 15 2 16 13 0 9 7 9 9 2 9 7 9 2 15 1 11 9 13 7 4 13 1 9 2
23 0 9 2 3 11 2 13 1 11 1 10 9 2 13 9 7 13 0 9 16 0 9 2
13 1 0 9 1 11 7 13 13 1 0 0 9 2
15 1 10 9 13 0 2 16 13 9 0 9 11 7 11 2
7 1 15 0 9 3 13 2
22 9 1 11 13 2 16 4 1 9 13 3 1 0 11 2 7 16 4 13 3 3 2
8 11 13 0 9 9 11 1 11
2 11 2
27 9 0 9 0 9 1 9 1 11 4 13 1 0 9 9 9 11 11 13 9 9 2 7 14 9 9 2
23 11 15 13 1 0 0 9 2 1 10 9 1 0 9 9 9 9 9 0 9 1 11 2
40 9 0 9 11 2 11 2 11 7 11 1 11 13 2 13 11 7 13 2 16 15 13 3 9 2 3 9 9 13 2 16 4 15 9 13 9 9 11 11 2
13 3 1 0 9 9 9 1 11 13 1 11 11 2
8 11 15 1 9 13 3 3 2
7 11 1 15 13 9 0 2
3 0 9 11
9 11 1 11 2 9 0 11 2 2
23 0 9 13 9 11 2 0 0 2 0 9 2 2 16 13 9 1 0 9 7 0 9 2
18 16 0 9 9 11 13 12 9 2 0 9 9 11 13 3 12 9 2
23 9 11 3 13 1 9 12 9 2 3 13 3 9 10 0 9 9 11 2 12 9 2 2
39 0 3 13 2 16 15 13 0 9 11 2 16 0 1 0 2 9 0 11 2 12 9 2 13 2 16 14 13 9 10 9 2 7 1 9 13 3 13 2
28 13 3 13 2 16 16 9 0 9 4 13 11 7 11 2 9 0 9 11 2 9 0 9 1 9 3 13 2
5 11 13 1 11 9
12 9 11 9 2 9 2 0 2 13 0 9 11
5 11 2 11 2 2
15 9 1 9 9 0 9 11 11 7 11 13 9 11 11 2
34 1 11 13 13 3 2 16 13 1 9 1 9 12 9 9 1 9 16 1 0 9 7 3 16 1 9 9 11 2 9 1 9 0 2
7 11 13 7 10 0 9 2
7 11 3 13 0 9 11 2
11 3 13 9 7 9 9 12 9 2 9 2
27 10 0 9 2 15 13 1 9 12 9 2 9 2 1 9 13 1 12 9 2 9 1 12 9 2 9 2
20 1 9 13 9 0 9 0 9 1 12 9 2 9 1 0 12 9 2 9 2
16 9 1 12 9 2 15 3 11 13 1 0 9 2 13 9 2
9 1 9 4 3 13 1 12 9 2
13 11 15 3 1 11 13 7 1 10 0 0 9 2
38 1 9 9 1 11 11 11 2 1 15 13 9 12 5 9 7 15 0 11 11 1 0 9 9 11 11 11 11 2 13 2 16 15 11 0 9 13 2
10 9 1 11 11 4 13 4 13 9 2
13 9 1 12 9 13 1 9 9 1 9 11 11 2
28 9 9 3 13 2 16 9 13 1 15 2 16 4 9 11 9 2 9 2 0 2 13 15 9 0 9 11 2
18 9 15 7 1 10 9 1 0 9 13 1 9 10 9 1 0 9 2
26 0 9 3 9 13 0 9 1 10 9 9 11 9 2 9 2 0 2 2 16 4 1 15 13 13 2
2 9 13
11 0 9 13 3 1 9 12 9 9 9 2
11 1 0 9 3 15 13 9 1 12 5 2
7 9 13 0 1 12 5 2
19 3 1 12 5 1 12 9 15 13 1 10 9 1 9 12 9 0 9 2
4 0 9 1 11
2 11 2
38 0 9 1 0 9 7 0 9 0 11 7 0 11 13 3 1 12 9 7 1 0 9 13 0 3 16 12 9 2 9 2 14 12 9 2 9 2 2
15 0 9 15 7 13 1 0 12 9 1 0 12 9 9 2
18 0 9 1 11 13 12 9 9 7 9 0 9 1 11 12 9 9 2
9 13 15 1 9 0 0 0 9 2
30 0 9 0 9 1 11 13 3 0 9 11 2 15 15 1 11 13 1 12 9 1 12 12 1 3 12 9 2 9 2
23 0 11 13 1 0 9 1 0 9 1 9 11 1 3 0 9 1 11 2 11 7 11 2
14 0 9 13 1 0 9 12 9 15 9 0 1 9 2
12 11 13 3 1 0 9 0 9 9 0 9 2
7 1 11 15 13 1 0 9
5 11 2 11 2 2
25 1 9 12 2 9 13 1 11 0 9 0 9 1 0 9 2 11 2 1 9 0 9 0 9 2
11 13 15 15 1 12 9 1 12 9 9 2
13 13 0 9 2 9 7 10 9 1 9 0 9 2
20 13 3 1 9 0 9 2 9 9 9 1 0 9 7 1 0 9 0 9 2
25 9 11 13 2 16 1 9 12 13 1 9 12 0 9 2 15 13 12 5 0 9 1 0 9 2
5 1 0 11 13 9
5 11 2 11 2 2
48 0 9 1 0 11 13 1 9 9 0 0 9 9 2 11 11 9 9 9 13 1 12 2 12 2 0 9 0 9 1 12 9 7 9 1 9 1 9 9 0 9 2 16 15 13 0 9 2
33 1 11 2 11 0 0 9 12 9 3 13 1 12 9 7 9 9 13 9 1 9 0 9 2 15 4 13 7 9 9 0 9 2
4 9 15 13 2
26 3 16 12 1 0 9 12 9 13 9 9 2 11 11 9 1 9 0 9 7 13 0 9 10 9 2
13 9 9 3 13 2 16 0 4 1 10 9 13 2
30 1 9 11 4 0 9 9 9 1 9 13 1 12 9 2 0 9 2 9 13 9 1 9 0 9 2 7 3 13 2
24 9 13 2 16 0 15 9 9 2 0 1 0 9 3 0 9 2 4 13 3 1 10 9 2
5 1 9 0 3 13
5 11 2 11 2 2
11 13 13 3 0 1 9 9 0 9 11 2
27 0 9 0 7 0 9 7 13 1 15 2 16 15 1 10 9 13 3 13 2 13 3 9 9 11 11 2
18 3 13 3 3 0 2 16 15 15 13 7 4 13 0 3 0 9 2
30 1 11 7 1 0 9 9 9 11 1 0 11 13 2 16 15 13 9 11 2 9 13 0 7 1 11 7 1 11 2
8 3 14 1 11 13 9 3 2
11 11 13 9 2 16 10 9 13 0 13 2
25 13 1 15 13 9 3 9 9 9 9 2 13 1 15 13 9 9 0 9 1 9 9 7 9 2
24 9 13 13 2 13 11 2 7 9 2 16 1 3 0 9 13 10 9 2 13 3 1 9 2
17 13 2 16 9 1 10 9 1 15 15 3 13 7 13 10 9 2
1 3
22 9 9 1 11 15 1 9 11 3 1 9 1 0 9 3 13 1 12 1 12 5 2
32 0 0 9 13 1 0 9 0 0 9 1 3 0 9 1 9 1 12 9 2 1 9 1 0 9 3 13 0 1 12 5 2
5 0 9 9 1 9
10 0 9 4 13 13 0 7 0 9 9
5 11 2 11 2 2
46 9 1 0 9 1 9 2 15 4 13 13 0 9 1 10 0 7 0 9 2 13 1 0 9 0 9 0 0 9 1 0 0 2 0 9 1 0 0 9 0 9 9 11 11 11 2
10 1 11 4 13 0 0 9 0 9 2
19 9 12 9 9 1 9 9 15 13 1 0 9 1 11 1 11 7 11 2
19 3 13 7 0 13 15 1 0 9 0 9 9 2 1 0 9 0 9 2
45 11 11 13 2 16 1 11 13 9 9 9 1 9 1 12 12 9 2 1 9 12 15 13 3 9 9 2 7 16 14 12 9 0 9 0 9 9 13 1 0 9 9 1 9 2
26 1 10 9 13 9 0 9 2 3 0 9 11 2 15 13 1 9 9 9 9 1 0 9 10 9 2
14 0 9 1 10 9 13 1 0 9 12 9 2 9 2
11 1 9 12 15 13 0 9 0 9 11 2
32 9 9 7 0 9 4 13 1 9 11 7 1 0 9 0 9 1 9 9 2 15 13 9 12 9 2 2 4 12 9 13 2
24 1 9 9 4 12 9 0 9 13 12 12 9 9 2 3 16 12 9 13 12 12 9 9 2
9 1 0 0 9 4 13 12 5 2
25 9 15 1 11 13 1 9 9 0 9 2 9 9 0 9 2 9 0 9 7 9 9 9 9 2
18 9 9 1 9 2 15 4 3 3 13 13 9 11 2 13 3 13 2
8 1 0 9 13 1 9 9 2
27 13 1 15 2 16 4 9 13 0 9 7 10 9 2 7 3 3 13 9 9 1 0 9 2 13 11 2
23 10 9 13 13 0 7 0 0 9 0 9 2 3 9 9 9 9 2 13 13 1 9 2
27 0 9 13 13 9 14 12 0 9 2 0 9 9 2 0 9 0 9 2 0 9 0 9 1 12 9 2
26 1 15 1 9 9 0 9 4 13 13 9 2 16 4 13 1 9 0 13 3 3 0 9 7 9 2
30 1 9 0 9 13 1 11 9 1 15 2 16 9 4 3 13 0 9 9 1 9 7 9 9 0 9 1 0 9 2
17 9 7 9 13 13 9 0 9 7 1 15 15 1 15 4 13 2
36 0 0 9 1 0 9 11 15 13 1 11 1 9 12 2 9 9 0 9 0 2 0 0 9 1 0 11 2 0 1 9 0 7 0 9 2
19 13 15 15 9 1 11 2 11 2 11 2 11 2 11 2 11 7 11 2
6 9 11 13 1 0 9
9 1 0 9 13 16 9 0 9 2
9 3 1 0 13 10 9 11 7 11
1 9
21 0 9 13 1 9 9 1 12 2 9 0 9 2 3 1 0 9 7 1 11 2
14 11 13 1 12 9 3 7 11 14 1 12 2 9 2
20 13 15 15 1 9 1 0 9 12 2 15 13 7 3 13 12 0 0 9 2
24 9 13 1 9 12 0 9 1 9 9 7 0 0 9 2 15 13 7 13 1 0 9 9 2
10 0 9 13 12 9 0 1 0 9 2
24 10 9 2 0 9 2 4 13 16 9 9 7 9 13 3 3 9 16 10 9 1 0 9 2
13 1 0 9 3 13 11 2 15 13 3 0 11 2
9 15 13 14 1 0 9 1 11 2
16 7 16 0 9 13 15 9 2 10 9 1 0 9 13 0 2
23 0 9 3 13 0 9 7 11 15 13 3 1 15 2 16 11 13 1 9 7 0 9 2
13 11 3 13 0 9 1 12 0 9 2 13 9 2
19 9 0 9 13 13 1 9 12 0 9 2 15 15 13 1 10 0 9 2
23 3 13 1 0 0 9 2 9 2 9 2 9 2 9 2 9 2 9 7 9 7 9 2
14 1 11 9 13 2 16 9 7 9 13 10 0 9 2
31 0 9 7 1 9 13 2 16 11 15 13 10 9 13 2 3 16 13 1 9 10 9 7 9 0 9 1 0 9 9 2
42 11 13 7 10 0 9 1 9 2 3 9 7 9 7 9 2 9 9 1 0 9 7 9 2 2 15 13 1 0 9 3 3 2 16 13 0 9 9 2 13 9 2
16 3 16 0 9 0 9 4 1 9 0 1 9 13 0 9 2
19 1 0 9 1 9 0 9 13 3 9 2 15 13 9 7 9 0 9 2
3 2 11 2
6 1 11 3 13 0 9
2 11 2
35 0 9 0 9 2 9 9 0 9 2 9 7 9 9 15 1 0 11 13 13 9 0 9 9 0 0 9 1 0 9 9 1 9 12 2
12 13 15 1 9 9 1 0 0 9 1 11 2
10 9 13 9 0 9 0 0 9 11 2
31 3 1 15 4 13 7 1 0 9 3 13 0 9 2 9 7 9 9 11 2 7 9 9 11 2 13 9 9 11 11 2
36 0 0 9 11 2 15 13 0 9 2 15 1 9 12 13 1 0 9 7 9 1 9 13 0 9 0 9 2 15 1 9 3 1 9 13 2
19 9 0 7 0 9 10 9 1 11 15 13 1 0 9 9 1 9 12 2
12 9 13 1 9 12 9 9 9 12 9 9 2
19 11 11 13 1 9 2 9 7 9 0 9 1 9 0 9 7 0 9 2
19 1 0 9 13 3 9 0 9 0 9 1 9 1 11 11 7 11 11 2
19 3 13 0 9 1 9 11 2 11 7 11 2 0 9 13 7 11 11 2
11 1 0 9 15 3 13 9 1 0 9 2
4 0 9 1 11
2 11 2
40 1 12 9 0 12 0 9 1 3 0 9 2 0 10 9 1 11 2 7 3 0 12 0 9 15 13 13 1 0 11 12 1 0 0 0 9 0 0 11 2
11 1 9 1 9 9 9 15 13 9 11 2
12 9 1 12 9 9 4 13 0 9 1 9 2
8 13 15 4 0 7 0 9 2
7 9 4 13 1 12 9 2
19 0 4 13 4 13 9 1 12 9 9 1 9 3 16 12 12 9 0 2
14 3 4 13 4 13 1 9 12 12 9 0 0 9 2
15 9 0 9 13 1 11 12 0 9 2 1 15 12 0 2
13 9 11 13 1 0 9 12 9 2 3 1 11 2
6 11 13 1 9 1 9
2 11 2
45 11 13 1 9 9 2 1 10 0 9 0 9 4 1 0 9 9 11 3 0 0 9 13 0 9 12 9 9 2 16 9 0 9 13 1 0 9 0 9 9 2 13 9 11 2
24 0 0 9 4 13 9 0 0 11 11 2 1 9 9 1 0 12 12 1 12 12 9 3 2
18 9 13 9 11 0 9 11 2 15 4 1 11 13 1 0 16 9 2
22 1 0 9 15 13 11 13 1 0 0 9 9 2 1 15 13 9 11 13 0 9 2
32 12 0 0 9 0 9 2 9 0 0 11 2 7 0 0 11 2 2 12 1 9 1 11 2 13 1 0 9 0 9 9 2
17 11 13 14 12 9 0 0 9 7 11 3 12 9 0 0 9 2
5 9 7 9 0 9
10 9 15 13 0 9 13 0 9 0 9
2 11 11
12 1 9 9 13 3 0 0 9 7 0 9 2
8 0 9 13 7 0 0 9 2
15 14 0 9 9 13 10 9 13 15 2 16 0 9 13 2
12 0 13 16 0 9 13 7 13 0 0 9 2
24 16 9 13 3 0 9 2 9 7 0 9 1 0 7 0 9 2 13 9 0 9 0 9 2
19 9 13 3 1 0 9 9 2 7 3 1 0 9 1 9 7 0 9 2
23 9 1 0 9 4 13 9 9 2 12 2 12 9 2 2 1 0 9 9 1 0 9 2
44 7 10 9 1 9 9 12 9 2 12 13 13 0 9 1 9 2 16 9 0 9 2 9 2 13 9 7 9 2 3 13 3 0 9 16 0 2 3 13 13 9 1 9 2
18 1 9 10 9 7 9 4 9 13 13 1 9 9 7 1 9 9 2
21 9 9 10 9 13 2 7 15 3 3 2 16 15 13 1 9 9 9 1 9 2
12 0 3 13 16 0 7 3 0 0 10 9 2
17 9 1 0 9 0 9 7 0 9 9 1 9 7 4 13 3 2
12 14 3 13 3 9 1 0 9 1 9 9 2
14 0 9 3 13 3 0 9 7 13 3 1 9 9 2
28 10 9 2 15 13 9 9 2 15 10 9 3 13 1 9 0 9 2 7 3 7 0 9 0 9 7 9 2
21 3 3 3 0 9 2 15 15 13 9 13 0 9 2 13 0 2 0 0 9 2
21 9 15 1 9 13 9 9 1 12 9 12 2 7 15 7 0 9 1 9 9 2
17 1 0 9 3 13 0 9 2 0 14 9 2 7 7 0 9 2
10 9 0 9 0 9 13 3 3 13 2
12 4 3 13 2 16 9 4 13 9 0 9 2
18 1 9 9 3 0 9 0 9 13 9 0 9 7 0 9 0 9 2
19 16 15 9 2 15 9 13 2 3 13 9 1 9 9 2 13 3 9 2
21 1 9 3 0 0 9 13 7 0 13 1 9 9 2 1 15 15 0 9 13 2
28 0 9 13 9 0 9 3 1 0 9 2 7 1 9 2 9 2 2 3 1 10 9 2 12 2 9 2 2
28 10 9 9 13 7 13 3 1 9 2 16 13 1 0 9 7 16 10 9 13 3 13 1 0 9 1 9 2
29 16 9 1 10 9 9 13 2 13 3 13 1 0 9 9 12 2 12 9 2 2 3 2 9 12 2 12 9 2
22 0 9 15 3 13 9 12 7 0 0 9 7 9 12 2 12 9 2 2 1 9 2
7 9 9 15 4 15 13 2
17 10 9 13 9 13 0 9 2 16 4 15 13 13 10 0 9 2
34 9 0 0 9 1 9 15 3 13 3 13 9 0 0 9 2 9 12 0 9 2 2 9 1 0 9 2 9 12 0 9 2 3 2
15 16 7 1 0 9 13 2 13 9 1 9 10 9 0 2
14 1 9 0 9 10 9 13 7 1 9 9 0 9 2
27 13 0 15 1 9 9 13 9 9 1 9 9 12 2 12 9 2 7 1 15 3 13 0 9 0 9 2
20 1 9 0 9 13 16 1 9 13 2 16 15 1 9 2 9 13 3 0 2
3 0 9 13
2 11 2
23 0 9 1 0 9 13 9 9 2 16 1 9 13 1 0 0 9 9 7 0 9 9 2
22 1 9 4 9 13 3 12 7 12 9 7 13 4 13 15 2 15 15 15 3 13 2
7 0 0 9 15 7 13 2
5 0 9 13 13 9
5 11 2 11 2 2
16 3 12 12 9 0 9 13 1 0 9 0 9 11 0 9 2
31 16 3 13 9 9 11 11 1 9 9 1 0 9 1 0 9 0 9 1 11 2 13 9 0 9 1 0 9 0 9 2
27 1 9 9 7 9 0 9 15 12 1 0 0 9 13 9 9 2 9 0 7 0 9 7 9 9 0 2
12 1 11 15 13 3 12 2 12 12 9 3 2
18 1 9 9 2 15 13 1 12 2 9 2 13 9 1 0 0 9 2
32 9 13 9 1 11 2 0 1 9 1 9 0 11 11 2 13 7 1 0 9 2 0 9 2 9 1 0 9 7 0 9 2
5 0 11 13 1 9
2 11 2
13 0 9 13 9 0 0 9 11 0 1 9 11 2
30 10 9 9 15 1 11 13 13 3 1 9 2 1 9 9 10 9 13 3 1 12 9 9 2 13 0 9 11 11 2
21 13 2 16 0 9 13 9 1 0 9 9 0 11 2 16 13 3 3 1 9 2
23 9 10 9 1 9 11 13 1 15 2 16 0 9 9 9 11 15 13 0 9 11 11 2
7 10 9 13 3 12 9 2
4 0 2 9 11
18 1 9 11 12 2 11 12 5 7 9 9 11 13 0 9 12 9 2
18 1 9 9 11 12 15 13 0 0 9 2 9 2 12 9 2 9 2
18 1 9 11 12 5 7 9 9 11 13 9 12 2 3 2 12 9 2
25 1 11 13 9 12 2 9 1 11 12 2 11 12 5 7 9 9 11 12 2 12 7 12 9 2
2 0 9
6 0 11 2 11 2 2
15 0 9 9 2 15 13 1 0 11 2 13 9 3 3 2
18 3 1 9 1 0 9 0 9 11 1 0 11 15 13 9 11 11 2
9 1 9 15 3 13 0 9 11 2
28 1 9 2 16 13 1 9 9 0 11 2 1 15 15 1 9 13 2 9 13 2 16 1 0 9 15 13 2
34 1 9 1 9 9 1 0 9 3 2 13 2 16 1 3 0 13 2 16 9 9 9 0 9 7 9 13 9 1 9 1 9 11 2
13 9 15 3 1 11 13 7 1 0 0 0 9 2
16 9 1 9 9 13 0 7 11 11 15 13 0 9 10 9 2
6 12 9 1 9 1 11
7 11 2 11 2 11 2 2
25 0 0 9 13 1 10 0 0 9 1 9 1 9 11 12 11 12 2 12 2 12 2 12 2 2
8 12 9 10 9 13 11 11 2
17 9 13 11 2 0 9 11 7 9 13 1 0 9 1 9 11 2
4 3 1 9 12
7 13 15 0 9 1 9 9
4 11 11 13 11
5 11 2 11 2 2
25 13 13 1 9 2 15 13 1 9 9 2 13 11 0 9 9 11 11 11 1 10 9 1 11 2
19 1 15 13 11 3 3 0 9 1 0 9 2 15 13 9 0 0 9 2
18 11 13 2 16 11 13 0 9 2 16 15 1 10 9 13 1 9 2
25 11 1 10 9 13 2 15 13 1 10 0 9 2 13 11 2 11 1 9 11 1 9 10 9 2
8 9 1 11 2 11 1 9 12
3 9 1 9
27 9 0 9 1 0 9 1 3 12 0 9 1 9 9 0 9 2 7 3 9 9 0 11 13 0 9 2
16 1 9 0 9 11 11 4 10 9 13 13 1 9 7 12 2
9 9 13 0 9 1 9 1 9 2
23 1 0 9 4 0 9 13 1 9 9 10 9 7 0 9 4 13 9 1 9 0 9 2
13 0 9 13 1 9 9 13 9 0 15 0 11 2
17 1 0 9 9 0 11 15 4 9 13 9 0 9 1 0 9 2
20 4 15 1 0 9 13 0 9 2 15 13 11 10 7 4 13 1 0 9 2
18 0 9 4 3 13 9 0 9 7 9 1 0 9 1 11 2 11 2
25 1 10 9 13 0 9 12 9 12 9 1 12 9 2 9 12 2 0 9 13 9 1 0 9 2
5 2 11 2 11 2
15 0 9 0 9 9 0 9 1 0 11 13 3 9 11 11
5 9 11 11 2 11
6 9 13 13 0 9 11
5 11 2 11 2 2
23 9 4 13 0 9 2 11 2 13 13 0 9 0 1 10 9 7 9 0 2 0 9 2
10 1 0 9 15 1 15 13 0 9 2
32 16 13 9 9 11 2 11 2 9 15 3 13 1 15 2 16 4 9 9 11 13 0 7 4 3 13 1 9 9 10 9 2
17 9 9 9 11 11 13 13 1 9 9 2 15 4 0 9 13 2
9 3 3 13 4 13 1 0 9 2
12 9 0 0 9 1 0 11 0 15 9 13 2
13 9 0 9 13 3 9 9 7 9 9 0 9 2
20 9 13 2 16 4 9 4 1 9 13 1 9 9 2 7 3 1 9 9 2
26 9 4 1 11 2 11 13 13 1 15 2 16 4 15 13 0 9 1 0 9 7 9 0 0 9 2
13 16 13 1 9 9 0 9 2 4 13 10 9 2
20 9 9 7 0 9 11 2 11 9 13 2 16 4 15 9 3 13 1 9 2
9 0 9 9 9 11 2 11 11 11
5 9 11 11 2 11
5 9 1 9 9 13
2 11 2
30 0 9 1 11 13 1 9 0 9 1 9 9 1 11 11 1 0 11 7 11 11 1 11 2 0 1 9 0 9 2
16 1 9 12 13 1 10 9 9 1 11 3 16 12 9 9 2
13 1 9 13 9 0 9 0 1 11 9 1 11 2
8 0 15 3 13 11 1 11 2
22 11 15 14 13 2 16 13 9 2 11 13 2 16 15 1 0 9 13 14 1 9 2
4 9 9 1 9
5 11 2 11 2 2
33 11 11 1 0 9 1 11 2 11 13 9 9 0 2 9 9 0 1 9 0 9 0 9 2 15 4 13 13 1 9 0 9 2
12 9 4 1 9 0 9 13 1 9 0 9 2
22 11 11 13 2 16 13 9 1 9 2 9 7 1 9 1 9 0 2 3 7 0 2
9 1 15 13 9 9 13 0 9 2
23 13 7 2 16 1 10 2 15 3 13 9 1 10 9 2 9 9 3 0 9 13 4 2
5 0 0 9 13 9
5 11 2 11 2 2
30 9 2 9 0 9 7 0 7 0 9 13 9 0 9 0 0 0 9 2 11 2 2 15 1 9 3 13 10 9 2
15 10 9 11 11 13 2 16 9 13 10 9 9 0 9 2
8 3 1 9 15 13 0 9 2
24 1 11 11 1 11 13 9 1 10 9 15 9 2 7 15 1 0 9 13 3 0 0 9 2
11 3 3 9 0 9 13 1 0 9 13 2
13 0 9 13 2 16 4 10 9 0 9 3 13 2
28 11 13 0 2 9 2 7 13 1 10 9 2 16 4 15 15 13 1 9 1 9 0 9 1 9 10 9 2
25 11 13 1 9 0 9 7 13 1 12 9 1 9 2 3 13 0 9 7 3 13 0 2 9 2
20 0 0 9 13 13 9 15 9 7 0 9 2 9 1 15 13 0 3 13 2
25 9 4 13 9 1 0 9 2 15 4 1 9 1 9 13 9 3 1 9 13 9 1 0 9 2
17 11 15 13 1 9 9 9 11 11 1 0 9 7 15 0 9 2
24 10 9 13 15 1 9 0 7 13 0 0 9 0 1 0 9 2 15 13 9 9 2 13 2
5 9 13 13 0 9
5 11 2 11 2 2
29 1 0 0 9 9 11 11 12 2 1 11 4 0 9 13 1 9 0 9 2 15 13 9 1 9 7 9 13 2
21 3 15 13 9 10 9 2 0 9 7 13 9 2 13 9 9 9 2 11 11 2
16 11 11 12 2 0 9 13 1 9 1 9 0 9 11 11 2
19 12 1 0 9 0 9 13 13 7 9 0 9 1 0 9 1 9 11 2
17 3 10 9 13 1 0 9 9 2 7 10 9 3 4 3 13 2
13 0 9 13 13 0 9 11 11 11 1 0 9 2
15 9 13 1 0 0 9 12 9 1 0 9 12 9 9 2
12 0 9 13 9 9 1 0 9 1 0 9 2
25 16 10 9 11 13 1 9 9 2 4 1 9 11 15 13 15 2 16 4 13 0 9 0 9 2
17 1 0 9 13 12 9 1 12 9 2 1 15 13 13 0 9 2
12 9 3 13 3 12 9 2 0 13 9 9 2
27 1 9 9 2 0 1 9 12 2 15 13 1 15 2 16 0 7 0 9 9 9 4 13 1 0 9 2
18 9 11 11 13 11 13 0 9 1 9 0 9 0 9 1 9 0 2
17 9 13 3 3 1 9 0 9 2 15 15 4 13 12 2 9 2
6 0 9 13 1 9 3
2 11 2
15 9 9 7 9 13 1 3 0 9 0 9 1 0 9 2
30 13 15 1 0 7 0 9 9 9 7 9 9 9 2 9 7 9 2 15 13 1 12 9 1 9 12 7 12 9 2
14 1 9 3 13 12 9 0 9 2 1 9 12 9 2
25 1 15 3 3 3 13 9 12 9 9 1 10 9 2 1 9 15 3 3 13 12 0 1 9 2
36 3 1 15 0 9 13 1 9 9 1 9 1 12 1 12 9 2 3 9 1 9 1 12 1 12 9 1 9 13 3 3 16 3 0 9 2
16 9 9 13 3 9 2 0 9 2 0 7 0 9 7 9 2
18 9 13 1 12 9 9 0 9 2 9 7 9 15 13 1 9 9 2
5 0 9 1 0 9
2 11 2
20 0 9 1 0 3 0 9 1 0 9 13 3 1 10 0 9 13 0 9 2
28 9 11 11 13 2 16 1 0 9 13 1 3 16 0 9 1 9 9 2 12 0 1 9 11 9 1 11 2
25 13 15 1 9 0 0 9 1 12 9 12 0 9 7 1 0 0 9 12 9 0 1 0 9 2
23 9 0 9 2 15 13 13 9 1 0 9 9 2 4 13 0 9 13 1 12 2 9 2
5 0 9 13 9 11
2 11 2
24 9 0 9 11 2 11 2 11 1 9 1 9 0 0 0 9 3 13 0 9 1 11 12 2
33 9 13 0 2 0 7 0 9 0 9 2 15 1 9 9 0 0 7 0 9 0 1 9 12 13 2 13 7 13 9 0 11 2
17 9 13 3 9 0 9 1 9 0 9 0 9 13 1 9 11 2
25 9 11 11 13 2 16 13 0 9 2 1 10 9 4 9 13 13 9 1 9 1 9 0 11 2
21 9 0 1 9 12 10 9 13 1 15 2 16 15 1 12 9 13 0 9 11 2
16 9 13 1 15 2 16 9 0 0 9 13 13 16 3 0 2
7 9 1 11 15 14 13 9
2 11 2
24 9 9 13 1 10 9 1 9 1 11 1 9 11 2 15 1 0 9 13 1 0 9 11 2
32 0 9 9 0 9 9 9 1 9 13 2 16 0 0 9 13 1 9 11 1 9 9 1 9 2 15 15 1 9 13 9 2
15 9 1 9 11 7 9 3 13 0 9 7 13 9 9 2
20 13 15 2 16 9 9 13 0 9 2 7 16 9 10 9 13 3 9 9 2
15 9 13 9 9 7 13 15 9 9 11 7 1 0 9 2
8 11 11 2 3 2 7 11 11
4 9 11 2 11
5 13 13 0 0 9
2 11 2
24 0 9 16 9 0 9 0 9 2 0 2 9 2 2 13 9 9 9 1 9 7 9 9 2
8 13 12 9 9 1 0 9 2
22 1 0 13 9 3 1 12 9 9 9 7 1 9 2 16 9 13 9 3 12 9 2
15 0 9 1 0 9 9 15 13 1 12 9 3 0 9 2
10 3 9 13 0 9 1 12 9 9 2
8 1 9 13 13 7 0 9 2
11 1 15 13 9 1 12 9 1 9 9 2
14 9 13 0 13 1 15 0 9 0 9 1 9 9 2
4 9 9 1 9
9 0 9 1 11 3 13 15 9 9
5 11 2 11 2 2
30 16 4 1 9 11 1 11 1 12 2 9 13 0 9 9 2 15 9 13 13 0 9 0 9 2 9 15 3 13 2
9 3 15 13 9 9 9 11 11 2
12 9 9 4 3 13 1 11 13 0 9 9 2
25 9 11 11 11 2 11 2 3 3 13 2 16 16 4 1 9 13 9 2 13 15 3 0 9 2
32 1 9 9 13 11 3 1 9 7 3 3 1 9 1 0 9 1 11 9 1 9 12 9 2 1 9 11 15 7 4 13 2
23 16 0 9 13 9 11 2 9 9 3 0 9 3 13 9 9 0 9 1 11 11 11 2
25 15 13 3 9 2 15 4 1 9 11 13 13 0 9 1 9 9 7 9 9 1 9 0 9 2
17 1 15 4 9 13 4 13 1 9 9 9 14 1 12 9 3 2
20 0 9 15 13 7 1 9 2 16 4 16 0 9 13 9 0 1 10 9 2
10 13 7 1 9 2 3 13 10 9 2
15 11 10 9 3 13 1 3 0 9 9 2 13 9 11 2
32 16 4 15 1 11 0 9 1 0 9 13 2 3 4 3 1 9 13 9 7 9 0 9 4 4 3 13 0 9 1 11 2
17 1 9 11 13 0 9 1 9 2 3 0 9 9 13 9 9 2
19 1 0 9 13 7 0 13 2 16 9 0 9 7 10 9 13 9 9 2
1 3
25 0 9 1 9 9 1 9 0 9 13 9 0 9 1 9 1 0 7 0 9 1 0 9 11 2
11 9 15 13 13 1 9 9 1 9 9 2
21 9 0 9 0 11 15 4 13 1 12 2 1 12 2 9 1 9 9 1 11 2
12 9 3 4 13 13 0 9 9 7 0 9 2
22 12 11 0 1 9 9 0 1 11 1 11 2 11 7 11 13 1 0 9 0 9 2
11 4 15 13 9 1 11 1 9 12 9 2
12 1 0 9 13 3 9 2 1 9 7 13 9
5 11 2 11 2 2
16 1 9 1 0 9 15 3 13 12 9 2 1 15 12 9 2
10 13 4 12 9 2 1 15 12 9 2
15 11 15 13 1 10 9 1 9 1 9 0 9 1 9 2
32 9 3 3 13 1 9 2 16 10 0 9 2 7 3 15 13 3 9 2 13 0 9 1 9 7 0 2 0 2 1 9 2
11 9 0 9 1 11 11 2 11 15 13 2
7 13 9 9 7 9 3 2
14 16 13 13 12 9 2 3 13 12 9 7 12 9 2
18 16 4 13 1 9 3 7 13 14 9 9 2 13 4 3 0 9 2
14 3 15 9 13 2 16 4 15 3 13 3 1 9 2
10 9 15 3 13 3 3 7 3 3 2
11 13 2 16 15 15 13 13 10 0 9 2
24 1 9 2 15 13 1 9 9 1 9 1 9 2 15 3 1 0 9 13 3 9 16 9 2
25 3 13 9 1 0 0 9 0 0 9 12 5 2 1 0 0 9 3 12 5 1 0 9 9 2
7 9 0 13 7 3 0 2
7 13 15 9 1 0 9 2
21 3 3 15 13 1 0 0 9 12 5 9 2 1 0 15 3 13 14 12 5 2
15 3 9 0 9 13 1 10 0 9 3 2 3 12 5 2
6 0 9 13 3 0 2
14 3 15 15 13 13 9 3 1 0 9 11 1 11 2
24 1 9 13 12 5 9 2 1 0 2 9 13 14 0 7 3 0 2 13 15 0 12 9 2
1 3
23 0 9 11 3 1 9 13 9 11 2 11 1 0 9 0 9 13 9 9 1 0 9 2
9 11 15 13 9 9 11 2 11 2
10 13 14 10 9 2 15 4 9 13 2
20 13 2 13 11 1 9 2 16 4 15 1 9 11 13 13 3 1 9 9 2
3 2 11 2
6 13 15 9 1 0 9
2 11 2
18 1 9 0 9 11 11 15 13 0 9 2 15 13 9 0 0 9 2
31 10 9 4 13 0 9 1 9 0 9 2 7 3 13 1 15 2 16 15 9 2 15 13 1 11 13 2 13 0 9 2
15 13 4 3 13 1 9 10 9 1 9 1 9 7 9 2
25 1 11 3 4 13 10 0 9 7 1 9 3 13 1 15 2 16 15 10 9 10 9 3 13 2
17 9 0 9 4 13 13 0 9 16 9 0 9 7 16 0 9 2
7 11 2 11 13 1 0 9
2 11 2
25 0 9 9 9 1 0 9 4 13 13 1 9 11 11 11 9 1 9 9 2 15 13 0 9 2
33 11 13 2 16 9 0 9 13 0 7 16 0 9 15 13 3 16 3 0 2 16 15 13 0 9 1 15 2 16 4 3 13 2
7 0 9 13 1 0 9 2
12 13 3 2 16 9 0 9 3 13 0 9 2
16 1 12 1 0 7 0 0 9 13 11 9 0 9 0 9 2
14 9 4 13 13 10 0 9 7 13 0 9 2 13 2
24 0 9 13 14 3 9 0 9 9 1 0 9 2 7 1 10 9 4 9 9 13 7 13 2
5 9 9 13 13 9
5 11 2 11 2 2
22 0 9 9 4 13 1 9 11 11 13 9 0 9 2 10 9 3 13 0 9 9 2
18 9 13 0 9 0 9 2 15 13 0 9 2 0 1 0 0 9 2
22 1 0 1 15 13 3 0 0 0 9 2 1 0 9 13 3 12 1 0 9 9 2
14 1 9 9 9 0 9 13 13 7 13 9 0 9 2
28 1 0 9 4 3 0 0 9 13 0 9 13 1 15 2 7 15 3 13 1 15 2 15 1 0 9 13 2
32 1 11 15 3 0 9 10 9 13 3 13 9 1 9 0 0 9 1 0 2 16 0 9 13 3 9 9 2 7 10 9 2
10 0 9 9 13 1 9 9 1 9 9
7 11 2 11 2 11 2 2
19 9 1 0 9 2 15 15 13 1 10 9 1 0 9 2 0 9 13 2
19 13 15 3 2 16 1 0 9 15 4 0 9 15 9 13 1 0 9 2
9 13 4 3 9 13 10 0 9 2
27 9 9 7 0 9 11 11 2 11 2 15 13 2 16 0 9 9 13 13 0 2 0 1 9 9 9 2
16 9 4 13 1 15 3 13 0 9 0 15 0 9 7 9 2
34 3 2 16 4 9 13 3 13 9 3 2 7 2 13 9 9 9 7 0 0 9 2 13 4 3 1 11 3 13 7 1 0 9 2
18 13 7 13 9 0 9 9 2 15 4 13 1 0 9 9 2 13 2
18 9 0 9 15 14 13 2 16 0 9 1 10 9 13 1 9 0 2
17 11 7 13 2 16 3 15 13 9 7 13 1 15 13 10 9 2
13 10 9 3 13 1 12 9 0 9 2 13 9 2
24 3 16 1 0 0 9 13 9 11 11 11 9 9 1 15 2 16 13 9 9 1 0 9 2
10 0 9 13 13 9 13 9 1 9 2
18 0 0 9 1 9 9 7 9 15 1 15 1 10 9 4 3 13 2
21 3 13 0 9 7 9 2 13 2 14 9 3 13 2 13 2 14 9 9 3 2
25 16 13 9 0 9 1 0 9 2 7 13 10 0 9 2 16 4 3 9 13 9 2 13 11 2
12 9 1 9 9 1 3 9 13 13 0 9 2
12 10 9 11 11 13 10 9 9 1 3 0 2
33 1 9 0 9 13 11 9 0 9 9 1 3 9 2 15 13 1 9 9 3 7 13 7 0 0 9 0 13 1 9 1 9 2
8 13 4 3 9 0 0 9 2
6 0 9 15 13 1 9
5 11 2 11 2 2
18 0 9 3 0 7 9 9 2 9 7 9 13 3 9 1 0 9 2
10 13 15 9 9 11 11 7 11 11 2
11 9 15 13 13 3 0 9 1 0 9 2
7 12 9 7 3 13 13 2
9 13 3 13 0 7 0 0 9 2
9 9 13 9 1 9 11 0 9 2
11 10 9 13 13 12 9 9 1 0 9 2
26 1 9 11 2 16 4 9 13 0 9 1 9 9 9 2 11 13 2 16 9 13 1 9 0 9 2
13 3 7 13 9 0 9 11 13 1 9 0 9 2
15 9 11 1 9 0 9 13 1 11 9 9 1 9 9 2
10 11 13 9 0 9 1 9 1 9 2
11 12 9 15 13 1 0 9 1 0 9 2
4 9 1 9 12
4 11 2 9 13
5 11 2 11 2 2
14 16 4 15 13 9 3 0 2 1 9 3 9 13 2
11 15 0 4 10 0 9 3 7 13 13 2
37 13 15 3 9 9 11 11 1 9 1 9 0 9 1 11 12 1 9 0 9 0 9 7 0 9 9 9 11 11 2 16 10 9 13 0 9 2
17 1 11 13 13 1 9 3 1 10 9 2 15 13 0 0 9 2
14 10 9 4 13 7 10 9 13 3 14 0 0 9 2
38 9 13 1 9 0 9 12 9 2 13 15 1 15 2 13 1 9 10 9 7 15 13 1 9 2 16 4 13 9 0 9 7 0 9 2 13 11 2
9 1 0 9 9 13 14 9 13 2
3 9 13 9
2 11 2
21 1 9 9 9 11 11 1 11 13 1 9 0 0 9 11 11 9 9 11 11 2
20 16 4 1 9 0 9 11 9 13 3 2 3 15 13 9 2 13 11 13 2
10 11 15 13 1 0 0 9 1 11 2
41 1 11 3 11 10 9 13 1 9 9 2 15 12 2 9 13 1 11 1 11 0 9 1 0 9 7 13 9 12 11 2 13 1 0 9 9 1 9 10 9 2
11 0 9 13 0 9 1 0 9 2 13 11
2 11 11
15 0 9 9 9 9 11 11 11 13 1 0 9 1 11 2
13 16 9 13 9 1 9 0 9 1 9 9 11 2
13 11 2 11 1 10 9 13 11 1 10 9 2 2
16 13 1 15 9 0 9 3 0 2 16 4 13 13 1 11 2
16 13 15 13 0 9 2 16 1 9 9 11 13 11 10 9 2
13 9 15 3 13 7 15 4 15 15 3 0 13 2
19 7 16 4 7 1 15 3 13 2 3 7 1 15 13 1 0 9 11 2
5 7 15 3 3 2
14 13 13 1 9 2 15 10 9 13 1 9 9 2 2
14 13 1 15 9 11 1 9 9 0 9 1 10 9 2
12 3 3 15 15 13 10 0 9 1 9 11 2
19 13 9 2 16 1 0 9 1 9 9 1 9 12 15 0 9 13 0 2
25 9 2 15 13 15 3 3 2 13 1 15 7 13 15 13 3 2 16 16 15 10 9 3 13 2
18 1 0 9 15 9 11 13 16 0 9 9 0 9 13 15 0 9 2
8 9 9 1 15 3 13 2 2
8 1 15 13 0 9 10 9 2
41 3 3 16 13 9 0 9 1 9 7 1 10 9 1 15 13 1 9 0 9 2 3 15 13 2 16 0 9 13 0 9 1 15 2 15 4 13 0 0 9 2
22 15 13 9 2 15 15 3 13 1 0 12 9 7 13 15 1 15 9 0 0 9 2
23 1 15 13 10 9 0 9 7 11 13 0 9 2 16 15 1 10 9 13 1 0 9 2
31 13 3 0 2 16 13 1 9 0 9 2 15 4 13 0 9 9 1 0 9 1 3 0 7 1 9 0 0 9 2 2
17 13 15 2 16 9 11 1 0 9 13 0 9 0 9 1 11 2
8 11 1 0 9 0 9 13 2
11 13 15 2 16 15 13 1 10 0 9 2
14 9 1 11 11 2 9 9 9 2 9 7 9 11 2
18 0 9 1 9 1 11 13 0 9 10 9 1 9 1 0 0 9 2
15 1 15 13 9 1 11 2 1 15 15 13 1 0 9 2
15 1 11 4 13 13 3 1 9 2 7 15 16 0 9 2
9 13 4 3 7 0 9 1 9 2
24 3 7 11 13 10 0 9 2 1 0 9 3 13 9 7 13 15 13 1 10 9 0 9 2
14 13 10 9 2 7 13 15 13 14 10 9 1 9 2
19 0 9 1 15 1 15 13 0 9 1 9 2 0 1 11 1 0 9 2
12 13 15 2 16 3 13 11 7 3 1 9 2
3 2 11 2
5 3 3 1 0 9
4 11 11 2 9
33 9 9 0 9 9 9 11 2 11 12 2 12 2 2 1 10 9 2 11 12 2 12 2 2 15 13 3 13 7 13 10 9 2
30 9 2 16 13 15 0 0 9 13 7 13 2 15 13 9 9 2 9 7 9 2 13 0 7 13 16 1 15 13 2
16 0 7 13 2 16 0 9 9 13 1 10 9 1 0 9 2
41 13 9 2 16 9 9 2 12 2 12 9 2 13 1 9 12 9 13 9 0 9 1 9 0 0 9 7 9 0 1 9 2 3 9 0 13 0 16 9 0 2
14 9 12 13 9 9 1 9 9 2 7 3 9 0 2
9 3 13 3 13 9 13 0 9 2
14 9 0 9 13 9 12 7 7 15 10 10 9 13 2
32 13 9 2 16 9 10 9 13 13 0 9 1 0 7 0 1 0 9 0 15 9 7 16 10 9 4 13 4 13 0 9 2
94 15 9 9 0 1 10 9 2 9 2 11 2 3 1 9 1 9 12 0 2 9 2 11 2 11 2 12 2 1 9 1 10 9 13 2 16 9 0 9 15 3 13 1 0 9 7 9 9 2 12 2 12 9 2 13 9 0 2 1 9 9 9 1 9 9 13 7 9 9 9 0 1 9 9 2 12 2 12 9 2 7 13 1 10 9 0 9 0 9 7 9 0 9 2
46 1 9 0 9 9 2 9 0 1 0 9 1 9 10 9 2 13 2 16 0 9 13 1 15 2 15 13 9 9 2 7 13 10 9 1 0 2 16 4 1 15 13 10 0 9 2
26 13 9 16 9 2 13 15 12 2 1 15 15 13 2 7 13 2 16 9 9 13 13 14 3 0 2
28 1 9 2 3 1 9 2 12 9 0 9 7 9 13 13 9 14 1 9 9 2 13 10 0 9 3 0 2
18 13 0 2 16 1 9 13 7 9 9 2 15 4 13 10 0 9 2
35 7 13 9 9 3 12 1 10 9 0 9 2 13 1 9 12 1 9 1 9 9 9 2 12 2 12 9 2 2 1 9 2 0 9 2
22 16 14 2 3 13 0 2 16 4 9 1 9 0 7 9 0 13 9 1 0 9 2
5 11 4 13 1 9
3 1 0 9
2 11 2
21 9 0 9 0 9 11 11 13 1 9 9 9 11 11 9 9 1 9 0 9 2
19 11 13 1 11 3 0 9 0 0 9 2 15 11 13 1 0 0 9 2
11 11 15 1 0 9 13 3 1 0 9 2
15 1 0 11 13 9 1 9 0 7 1 11 1 0 9 2
7 11 13 1 11 12 9 2
5 0 9 13 1 11
5 11 2 11 2 2
34 9 0 9 7 9 9 9 2 11 11 2 15 12 2 9 13 1 9 11 11 2 13 11 2 16 9 13 1 9 9 12 0 9 2
17 9 1 15 13 2 16 9 13 1 9 7 9 2 11 3 13 2
13 1 10 9 13 2 13 1 9 2 11 3 13 2
7 12 7 4 13 1 11 2
21 13 13 2 16 15 13 1 9 0 1 9 9 1 0 9 7 3 1 0 9 2
15 13 15 14 1 9 11 2 7 3 1 9 11 2 9 2
25 13 4 2 16 10 9 1 0 9 4 13 2 7 13 15 7 3 1 15 2 13 9 2 11 2
4 9 13 9 2
9 1 0 9 4 13 1 0 9 2
8 9 14 13 1 9 15 0 2
18 0 9 15 7 1 0 13 15 2 16 10 9 13 1 0 9 0 2
11 13 15 3 3 9 9 9 7 0 9 2
9 1 10 9 13 15 9 3 0 2
15 13 0 9 2 3 4 13 9 10 9 7 15 13 0 2
14 13 2 14 9 3 13 1 9 2 13 13 9 9 2
8 0 9 1 9 13 10 9 2
24 16 4 15 3 13 13 9 0 9 1 9 2 13 1 15 9 9 2 13 11 9 2 11 2
5 1 9 13 1 9
5 11 2 11 2 2
39 0 9 2 1 15 15 4 13 9 2 15 1 9 13 9 9 0 9 13 0 9 1 11 12 11 2 12 2 12 9 2 2 15 13 7 13 1 11 2
28 1 10 9 15 0 9 13 1 9 2 13 1 15 9 7 13 15 1 9 0 9 7 3 16 12 12 9 2
11 16 13 1 9 2 12 11 15 9 13 2
11 1 10 9 4 1 10 9 1 11 13 2
4 3 1 0 9
7 9 0 11 13 9 1 9
2 11 2
21 1 9 9 9 1 0 9 0 0 9 0 11 13 0 9 0 9 11 0 9 2
35 0 0 9 9 12 4 13 1 9 0 2 11 2 11 2 1 12 1 12 9 7 1 12 1 12 9 2 1 9 11 2 9 9 0 2
11 13 13 0 1 9 11 7 1 9 11 2
15 0 9 9 12 7 12 4 13 1 9 11 7 9 11 2
23 1 9 4 1 12 9 13 1 9 1 0 9 1 11 7 1 9 1 11 9 9 11 2
20 0 0 9 9 12 13 1 12 1 12 9 2 1 9 1 0 2 9 11 2
18 1 12 1 12 9 2 13 10 9 1 9 1 11 7 9 9 11 2
14 0 9 12 2 12 7 12 1 9 9 1 11 13 2
7 9 9 4 13 1 9 2
10 9 0 7 11 4 13 3 16 0 2
17 1 9 11 7 11 13 13 1 9 9 1 9 11 7 9 11 2
10 0 9 1 11 9 13 1 12 9 2
14 1 0 9 13 12 2 9 9 11 13 1 0 9 2
4 9 3 13 13
5 11 2 11 2 2
18 9 13 1 0 9 1 12 0 9 3 1 9 1 0 9 9 0 2
21 0 9 0 9 1 0 9 3 13 2 7 15 1 12 9 9 2 12 5 2 2
19 16 9 9 1 0 9 13 1 12 5 2 9 0 3 13 1 12 5 2
10 0 12 1 15 13 9 1 12 9 2
13 9 9 13 1 9 9 11 2 11 13 10 9 2
9 1 0 13 0 9 0 9 9 2
7 9 9 13 3 1 9 2
19 13 15 0 9 1 9 0 9 7 9 15 3 13 1 0 9 0 9 2
4 9 9 13 9
5 11 2 11 2 2
23 0 9 15 13 13 9 0 11 11 2 1 11 2 15 1 9 13 1 9 1 0 9 2
28 16 3 13 0 9 11 11 2 1 0 9 15 13 7 12 9 9 9 2 15 15 1 10 9 1 11 13 2
25 9 13 14 12 9 0 0 9 2 16 0 15 13 13 14 12 9 1 9 2 3 1 9 13 2
28 1 0 9 13 1 9 3 2 3 15 11 11 2 13 13 9 2 3 15 7 13 9 9 7 13 15 13 2
24 1 9 15 13 12 9 1 9 2 0 11 11 2 1 11 7 0 11 11 2 1 0 11 2
16 9 1 9 15 7 13 2 16 12 9 13 1 9 13 0 2
13 11 11 2 4 13 1 9 1 0 9 1 11 2
17 16 13 11 2 11 2 1 11 11 2 13 3 1 9 13 9 2
27 9 9 13 0 13 14 1 9 9 9 1 12 9 2 7 1 9 9 13 9 9 12 9 0 1 9 2
22 1 9 1 9 13 3 1 9 1 0 9 2 1 0 9 15 12 9 13 9 9 2
7 1 9 11 2 11 3 9
2 0 9
5 11 2 11 2 2
31 9 1 11 11 2 0 1 0 9 9 11 11 4 3 13 9 0 9 1 11 2 16 15 1 9 13 12 9 1 12 2
29 16 0 1 10 9 1 9 2 3 13 0 9 2 13 2 16 13 1 0 9 2 9 13 9 2 15 15 13 2
21 9 13 14 12 9 1 9 0 1 9 9 2 15 15 11 11 2 13 0 9 2
24 9 13 1 9 0 9 0 1 11 11 2 2 15 4 3 13 1 0 9 9 1 0 9 2
40 11 11 2 0 9 0 9 0 11 2 1 15 11 11 2 13 2 9 13 2 16 0 13 1 0 9 9 7 16 9 9 13 13 0 9 7 9 2 9 2
20 11 11 2 1 9 1 9 0 9 3 13 2 16 4 13 9 1 0 9 2
24 12 3 0 9 13 0 9 9 1 9 1 12 2 1 12 2 9 0 9 1 9 9 0 2
37 12 1 15 3 3 1 9 1 0 9 13 2 16 1 9 1 0 13 1 0 2 16 14 15 13 10 9 1 9 7 13 15 1 15 3 9 2
15 9 13 12 9 0 9 2 16 11 11 2 9 9 13 2
22 0 15 13 7 13 15 15 2 16 13 1 9 2 16 0 15 9 13 9 1 9 2
12 1 9 1 9 13 7 3 15 13 1 9 2
1 9
21 9 9 11 1 11 9 2 11 11 13 1 12 2 9 1 9 0 9 0 9 2
9 13 15 15 9 2 11 2 11 2
5 0 9 13 1 9
24 0 9 11 12 13 0 9 1 9 0 9 1 9 0 9 2 15 13 13 1 0 0 9 2
21 9 13 10 9 13 9 9 1 0 9 1 11 12 1 12 2 9 1 0 9 2
11 1 0 9 4 9 13 13 1 9 9 2
16 9 9 7 9 7 9 9 13 13 2 13 15 13 15 0 2
16 9 9 4 3 13 3 13 9 9 1 0 9 7 9 9 2
17 0 9 13 1 9 9 13 1 9 9 3 0 2 3 0 9 2
27 1 9 0 9 13 0 14 9 9 1 9 9 2 9 0 7 0 9 2 7 7 9 1 9 0 9 2
12 9 15 3 13 9 13 3 1 9 0 9 2
32 1 9 9 0 1 9 13 0 9 13 1 9 0 0 9 7 9 1 9 1 0 7 0 9 2 1 9 9 7 9 11 2
3 2 11 2
2 0 9
1 9
2 11 11
20 13 9 0 9 1 10 0 9 1 9 9 9 2 9 0 9 7 10 9 2
15 9 2 10 0 9 1 9 0 9 13 1 9 9 13 2
6 9 2 2 9 13 2
15 15 4 15 13 2 16 4 15 1 0 9 13 10 9 2
36 9 4 13 9 3 7 9 9 0 9 4 3 1 10 9 1 9 13 2 16 9 7 9 2 15 3 13 9 2 15 9 13 9 0 9 2
24 13 15 9 12 9 0 0 9 1 9 11 2 10 0 9 15 13 1 9 1 12 9 9 2
28 0 9 2 0 0 9 2 15 1 0 9 13 0 9 0 0 9 11 11 2 15 15 13 1 12 10 9 2
13 11 7 13 1 0 9 13 9 0 9 12 9 2
14 13 15 9 2 15 1 0 9 1 0 0 9 13 2
7 9 10 9 3 3 13 2
14 11 13 7 0 2 16 10 9 3 13 12 9 9 2
8 15 2 15 1 9 13 9 2
30 0 9 13 3 3 13 2 13 1 15 12 9 2 1 9 9 9 7 0 9 2 15 0 9 3 1 10 9 13 2
7 15 1 10 9 13 9 2
3 14 15 2
20 0 0 9 2 7 3 13 2 15 2 15 1 15 13 2 3 13 1 9 2
20 9 9 2 9 9 2 7 13 2 16 10 9 13 7 9 13 13 0 9 2
36 9 13 7 15 2 16 9 3 4 13 13 1 9 0 9 7 0 9 2 15 1 9 1 9 1 0 9 12 9 0 9 13 1 0 9 2
21 1 9 9 13 0 7 9 9 2 7 9 0 9 2 3 0 9 1 0 9 2
19 10 9 3 13 9 9 0 9 1 9 9 2 7 13 13 10 0 9 2
9 1 10 9 13 9 1 10 9 2
20 9 0 2 9 0 9 11 2 11 2 3 2 7 11 2 11 1 0 0 9
5 9 11 11 2 11
5 0 9 1 0 9
1 9
2 11 11
26 1 9 1 0 9 0 9 13 13 0 9 3 13 0 9 3 0 7 9 9 2 9 7 9 11 2
38 9 9 11 2 11 13 1 15 2 16 1 9 1 0 9 11 2 15 1 10 9 13 3 9 16 9 2 15 1 0 9 1 0 9 9 9 13 2
20 13 7 2 16 10 2 15 13 1 9 3 10 9 2 13 13 0 12 9 2
15 1 9 1 9 1 10 0 9 13 3 9 1 0 11 2
12 10 0 9 1 9 13 3 9 2 7 13 2
14 9 13 3 1 9 9 0 9 2 10 9 9 13 2
8 13 1 9 7 9 0 9 2
12 15 3 9 2 3 1 0 9 2 13 13 2
4 15 13 13 2
24 9 9 11 11 11 2 15 13 9 1 0 9 7 15 0 9 4 1 0 9 13 1 9 2
35 13 14 2 16 9 9 0 9 13 1 11 3 11 11 2 11 2 15 13 1 15 0 9 9 1 0 9 2 1 0 9 1 9 9 2
12 13 15 2 16 3 15 13 1 9 10 9 2
17 11 1 0 9 9 13 2 16 15 12 9 13 13 0 0 9 2
28 13 2 14 15 15 15 2 13 15 1 15 13 2 13 10 9 7 13 0 9 1 12 9 0 9 1 0 2
16 9 9 13 7 13 2 16 3 15 13 10 0 0 9 0 2
5 0 9 13 1 9
2 11 11
28 9 1 9 9 1 0 0 9 7 0 0 9 1 0 9 13 9 9 7 3 9 1 10 0 7 0 9 2
14 9 2 9 4 13 1 9 2 7 16 14 14 3 2
9 9 3 13 10 0 7 0 9 2
21 0 0 9 0 9 2 1 15 9 3 13 0 9 2 3 4 3 3 3 13 2
5 15 15 3 13 2
33 1 9 12 2 12 2 3 13 15 9 1 9 0 9 10 0 0 9 2 3 9 1 9 2 13 10 0 0 9 1 0 9 2
13 13 15 0 9 1 0 0 9 7 0 0 9 2
30 3 2 1 10 9 9 0 9 2 13 3 15 0 7 13 2 16 0 9 13 9 2 15 13 9 13 0 0 9 2
10 10 9 15 3 13 14 1 12 9 2
9 1 15 15 0 9 13 3 13 2
12 9 2 15 13 9 2 13 3 13 7 13 2
19 9 1 9 2 15 13 13 10 9 2 13 0 9 16 1 9 0 9 2
19 16 0 9 13 9 2 16 1 0 9 13 1 0 9 1 0 9 13 2
23 16 15 9 13 3 12 7 12 9 2 15 13 10 9 2 1 0 9 13 2 7 3 2
17 13 15 0 9 12 9 1 9 7 9 0 9 1 3 0 9 2
15 0 9 7 13 1 9 9 1 15 3 2 16 13 0 2
20 9 10 9 13 9 2 16 9 13 13 1 0 9 9 2 16 4 4 13 2
14 15 3 13 1 3 0 9 1 9 13 1 0 9 2
15 0 9 13 0 9 9 2 1 10 9 3 3 0 0 2
7 3 15 13 1 0 9 2
36 1 9 15 13 2 16 9 0 15 1 0 9 9 13 1 10 9 1 0 0 9 2 7 14 1 9 9 9 2 3 15 3 13 0 9 2
20 1 9 13 9 1 9 11 1 0 9 15 1 0 9 3 15 13 7 13 2
24 13 7 1 0 9 2 1 15 15 13 2 7 9 15 13 2 16 4 13 9 1 12 9 2
23 9 11 13 7 3 1 9 3 13 9 2 3 1 0 9 1 0 0 9 13 0 9 2
16 1 15 15 3 13 2 7 16 7 10 9 3 13 0 9 2
28 9 9 13 9 3 3 2 13 2 16 13 15 0 9 1 0 0 9 7 0 9 1 9 1 12 2 9 2
24 11 13 0 3 3 0 9 2 7 15 13 10 9 7 10 9 2 15 15 13 1 9 9 2
22 13 2 16 3 12 2 9 9 9 13 2 10 9 4 13 1 9 9 1 11 7 9
36 9 13 1 15 2 16 0 9 15 3 13 9 1 0 9 2 15 13 2 7 1 15 13 13 2 1 9 1 0 9 2 1 9 0 9 2
14 13 3 9 2 16 3 0 9 13 1 0 9 0 2
35 0 7 0 9 9 11 13 0 9 1 0 0 9 0 1 0 0 9 9 0 7 0 0 9 1 9 7 10 9 9 13 1 9 9 2
15 13 13 3 16 12 12 9 1 0 9 1 12 9 9 2
12 1 9 11 7 9 0 9 13 1 0 9 2
5 9 13 7 0 2
16 9 1 0 9 13 3 13 15 1 15 7 1 10 0 9 2
8 0 9 1 0 9 13 9 2
29 0 0 9 3 13 0 9 0 9 2 7 1 0 9 1 11 7 10 9 7 0 9 3 0 9 16 15 0 2
6 9 2 7 0 9 2
2 11 11
16 9 0 9 11 1 9 0 9 13 1 0 9 3 15 9 2
13 1 9 1 0 9 0 9 13 0 1 0 9 2
25 3 1 15 9 9 0 9 13 0 7 0 0 7 0 9 2 16 4 15 13 0 9 0 9 2
25 3 15 7 1 10 9 13 7 9 1 0 7 0 0 9 2 15 4 9 0 9 13 13 0 2
27 9 0 0 9 2 15 4 3 13 2 16 9 0 9 13 4 13 9 10 9 2 15 13 1 9 9 2
15 0 9 1 10 9 15 13 1 12 2 9 1 0 9 2
36 3 13 0 9 9 1 9 2 15 4 13 2 16 2 1 9 0 9 2 13 4 9 13 16 0 7 9 1 0 9 13 13 9 0 9 2
46 10 9 2 3 0 9 3 1 9 2 3 10 9 1 10 9 13 0 9 0 9 1 9 0 9 2 4 13 0 9 3 3 2 16 13 0 9 2 15 13 9 0 9 1 9 2
27 9 0 9 2 0 1 11 2 3 13 0 9 0 9 2 13 3 9 13 2 16 0 9 4 3 13 2
13 13 9 1 9 1 0 0 9 13 3 3 0 2
35 9 2 16 4 0 9 13 0 9 13 9 0 9 2 7 2 16 9 0 0 9 13 0 7 0 9 9 0 9 2 2 13 3 0 2
15 3 9 15 2 3 0 9 13 0 0 9 2 13 11 2
34 16 0 0 9 0 9 13 4 1 9 13 3 0 9 2 13 0 0 9 3 9 12 2 9 9 9 2 16 0 9 13 12 9 2
20 1 1 0 9 9 1 3 2 13 9 0 9 1 9 2 15 3 9 13 2
22 1 0 9 13 3 3 0 2 16 15 9 13 3 2 7 16 3 13 9 0 9 2
40 1 15 13 10 9 3 2 9 9 0 9 2 15 13 14 9 1 0 9 2 7 3 9 1 11 7 9 0 9 2 2 7 0 0 0 9 7 0 9 2
27 1 1 15 2 16 15 3 13 9 2 3 10 9 13 1 10 9 2 13 0 0 9 9 0 0 9 2
15 0 9 13 3 9 9 1 9 2 1 15 13 0 9 2
16 1 10 9 15 3 9 13 9 13 2 16 4 3 13 9 2
22 0 9 2 15 10 0 9 3 7 3 13 2 7 13 13 1 9 1 0 0 9 2
11 3 3 15 7 13 13 1 9 1 9 2
16 9 0 9 3 1 0 9 9 9 1 9 0 9 3 13 2
22 1 9 1 0 7 1 10 9 3 0 9 1 0 0 9 13 1 9 0 0 9 2
42 15 4 7 13 9 9 2 10 9 13 0 0 9 2 16 7 3 13 0 9 0 0 9 2 2 3 4 7 13 9 9 1 9 7 9 0 9 1 9 0 9 2
23 3 2 12 1 0 0 9 1 10 9 2 0 9 12 2 15 13 3 1 0 9 9 2
12 0 9 1 9 9 13 13 0 9 0 9 2
10 9 0 9 15 1 15 13 0 9 2
22 0 9 9 7 9 0 9 2 16 4 13 3 3 2 13 3 13 0 9 0 9 2
17 1 0 7 0 9 0 9 13 0 9 14 3 0 7 0 9 2
13 3 7 3 9 1 0 9 13 1 0 0 9 2
31 16 7 9 0 0 9 13 13 0 9 0 15 0 9 2 13 4 13 9 0 0 9 7 13 10 9 1 9 0 9 2
19 13 7 2 16 4 1 0 9 13 13 0 9 10 0 9 1 0 9 2
1 9
3 9 11 11
22 9 11 11 11 11 15 1 12 9 13 0 9 2 13 0 9 7 3 1 15 13 2
44 1 9 2 3 15 1 9 13 10 9 9 0 9 2 15 0 0 9 13 15 13 7 0 9 1 9 0 9 7 10 9 0 9 15 13 2 15 11 13 1 0 9 11 2
19 15 11 13 9 9 2 0 9 2 0 9 2 3 7 9 1 0 9 2
40 1 9 2 16 11 3 13 0 0 9 2 7 13 1 15 0 2 11 11 13 9 2 0 0 9 9 2 12 13 12 9 9 7 15 15 11 13 1 12 2
23 1 0 9 14 11 13 3 16 1 10 9 1 9 2 16 3 13 1 11 2 7 11 2
33 16 3 3 13 9 12 9 9 2 12 1 9 11 1 11 3 2 13 11 2 15 15 1 9 0 9 13 1 9 2 1 0 2
14 9 15 13 16 0 9 2 15 11 13 1 9 9 2
34 11 2 15 13 0 0 0 9 2 14 3 13 9 2 13 15 1 9 2 15 13 0 0 9 0 0 9 7 3 1 15 3 13 2
15 0 13 3 10 9 13 15 1 0 0 9 9 2 12 2
23 1 10 13 9 0 9 7 0 9 2 15 15 0 9 13 13 2 7 7 10 0 9 2
9 0 9 13 3 9 7 1 11 2
33 1 10 9 13 1 11 1 9 1 0 9 13 1 0 9 9 9 9 11 11 9 9 0 11 2 15 1 11 13 9 0 9 2
19 3 15 13 1 9 9 2 15 15 0 11 7 0 9 1 0 9 13 2
23 1 9 3 0 9 14 1 9 13 0 9 2 16 1 9 9 0 9 15 13 14 13 2
18 1 9 11 15 13 3 9 2 15 3 13 9 11 7 9 0 9 2
28 13 2 14 15 9 1 9 9 11 2 15 9 1 9 13 9 9 9 1 0 9 2 13 4 15 1 9 2
43 0 9 2 9 1 11 0 11 2 0 11 7 11 15 13 1 9 2 15 14 3 3 13 2 16 9 9 2 12 13 1 0 9 1 11 2 1 15 13 7 15 13 2
22 15 3 13 1 15 2 16 15 0 2 0 2 0 7 0 9 10 9 13 7 9 2
4 13 9 0 9
2 11 2
18 0 9 13 3 1 9 11 12 0 9 2 0 1 9 1 0 9 2
17 0 11 13 1 0 9 0 0 9 1 9 11 2 0 9 2 2
18 1 0 9 13 9 1 15 2 15 15 1 9 13 2 0 9 9 2
24 0 9 1 0 13 9 9 9 11 11 2 12 2 7 0 9 9 11 11 11 2 12 2 2
22 12 13 1 15 2 15 13 1 3 16 12 9 2 15 11 1 9 12 13 1 11 2
16 0 9 15 13 1 0 9 1 0 9 2 1 15 12 13 2
4 11 11 11 13
2 11 2
20 11 3 13 0 9 9 11 1 9 7 9 2 15 15 13 1 9 1 11 2
13 13 15 3 9 11 11 11 1 9 1 0 9 2
19 11 13 10 9 1 3 0 2 13 7 2 16 3 12 9 13 3 0 2
29 0 9 0 0 9 2 11 2 11 11 3 13 2 16 4 13 0 9 13 9 1 0 9 9 1 9 1 9 2
18 9 11 3 13 2 16 0 9 4 13 13 13 0 9 9 0 9 2
19 0 9 9 11 1 9 7 9 4 13 9 2 16 9 13 9 0 9 2
8 13 15 1 15 3 9 9 2
6 9 13 14 9 11 2
6 0 9 13 1 9 11
4 11 2 11 2
28 0 0 9 13 9 0 0 9 2 11 2 2 16 4 13 0 0 9 1 9 11 2 0 11 1 9 9 2
33 9 11 3 13 9 11 2 11 7 11 1 9 2 15 0 9 13 12 2 9 7 3 1 0 9 13 3 16 12 9 0 9 2
36 0 9 13 9 1 9 11 2 1 10 9 13 1 12 0 9 2 16 4 13 0 9 0 9 1 11 2 15 4 13 9 1 9 1 9 2
6 11 13 0 9 1 11
2 11 2
27 9 0 0 9 1 11 3 3 13 9 11 1 11 11 11 2 15 1 11 13 1 0 9 9 11 11 2
31 1 9 11 2 11 13 2 16 16 11 4 13 0 9 0 9 2 13 15 11 0 13 9 1 0 9 1 9 0 11 2
12 9 0 9 1 11 13 11 1 0 9 9 2
25 13 14 1 0 2 7 7 1 0 9 2 7 1 9 0 9 1 9 13 0 0 0 9 11 2
4 3 9 13 9
9 9 9 11 7 11 13 1 0 9
7 0 9 11 1 11 11 11
10 9 10 9 9 1 0 9 13 9 2
8 3 16 13 7 10 0 9 2
38 0 9 9 0 9 1 11 7 13 15 0 16 0 9 2 1 15 12 9 13 3 3 0 2 13 15 3 1 0 9 0 9 2 7 15 13 15 2
10 7 12 0 9 2 7 12 0 9 2
13 3 15 7 13 9 1 11 7 1 11 3 0 2
22 11 11 9 1 10 9 1 0 9 1 0 9 11 13 9 9 10 9 1 0 9 2
36 11 13 3 15 3 2 16 13 1 9 9 0 9 7 16 15 13 13 1 0 9 11 7 0 9 2 3 16 11 2 11 2 11 7 11 2
28 0 9 7 13 11 3 1 9 15 16 11 2 16 13 1 9 10 0 9 2 1 9 1 11 13 13 9 2
30 13 9 2 16 3 3 15 15 13 2 7 0 9 0 11 7 9 9 0 9 0 9 13 1 0 11 16 0 9 2
18 7 15 13 7 0 9 0 9 11 11 1 11 2 15 3 13 9 2
12 7 7 3 0 9 11 1 10 9 1 11 2
21 11 11 13 9 1 11 2 16 9 9 0 2 0 0 9 13 1 12 9 0 2
14 13 13 9 9 9 7 9 0 9 1 11 2 13 2
10 3 0 9 2 3 16 1 9 11 2
5 14 1 12 9 2
42 9 11 11 3 13 2 16 11 13 0 3 3 1 10 9 3 7 3 13 9 9 9 2 13 15 7 9 2 16 11 0 1 11 4 13 9 13 15 3 16 3 2
29 0 0 9 2 9 0 3 1 9 0 9 7 1 15 0 9 13 3 9 15 2 16 15 11 1 11 13 13 2
23 1 15 13 9 0 9 2 1 15 13 0 0 9 2 9 13 7 3 15 1 15 13 2
8 3 0 9 1 11 15 13 2
32 1 9 0 9 1 9 0 9 9 15 1 12 9 1 15 13 9 12 9 1 0 9 2 11 7 11 3 13 1 0 9 2
15 16 1 10 9 2 15 13 3 9 7 0 9 0 9 2
5 0 9 13 0 9
3 0 11 2
22 9 0 1 0 0 9 13 1 0 9 1 9 12 7 12 9 0 1 9 0 9 2
22 13 15 15 1 9 0 9 11 11 7 11 11 11 2 15 15 3 13 1 0 9 2
19 9 9 11 15 13 13 2 16 15 1 9 9 1 0 9 13 9 9 2
9 9 9 13 9 2 7 0 9 2
16 1 10 9 9 13 9 7 13 15 15 1 9 9 1 9 2
18 0 2 15 15 13 9 9 1 9 9 9 2 13 0 9 0 9 2
20 3 13 2 16 1 15 13 7 13 2 0 2 16 0 2 13 15 1 9 2
17 0 9 9 1 9 2 15 13 1 9 1 0 0 9 2 13 2
4 9 1 9 11
4 11 2 11 2
42 1 9 9 0 9 2 11 2 1 0 9 0 9 2 11 2 2 15 15 13 9 1 9 12 2 3 13 9 0 9 11 9 11 11 11 1 0 9 0 0 11 2
14 0 9 1 9 0 0 9 3 13 13 2 13 9 2
21 1 11 13 13 9 1 9 0 9 1 9 3 10 9 1 0 9 7 1 11 2
9 13 13 3 1 0 9 0 9 2
25 0 9 11 11 13 9 0 0 9 2 11 2 1 0 9 10 9 11 2 0 1 0 9 11 2
27 9 0 9 1 9 1 9 13 2 16 9 13 10 9 1 9 0 9 1 9 0 9 7 9 0 9 2
23 9 0 11 13 1 15 2 16 15 11 2 11 2 11 2 11 7 11 13 9 0 9 2
28 0 9 0 9 3 13 9 0 9 2 1 15 13 12 1 12 0 9 11 1 9 9 13 1 9 10 9 2
16 9 0 9 1 9 11 13 1 9 11 10 9 1 9 11 2
28 9 0 0 9 9 3 1 11 13 2 16 10 9 13 9 1 9 0 9 1 9 0 9 1 9 0 9 2
19 9 3 13 1 11 16 1 9 0 9 7 16 1 0 9 9 9 9 2
4 9 11 2 11
9 9 1 0 9 1 11 1 0 9
4 11 2 11 2
5 13 1 0 9 2
43 13 15 9 2 16 15 15 13 13 0 11 2 16 0 9 13 3 0 2 13 3 11 11 1 0 9 1 11 0 1 9 0 9 9 9 12 9 0 9 7 9 11 2
20 13 2 16 13 3 0 2 16 4 13 0 9 0 7 16 4 3 13 9 2
26 1 0 9 13 1 11 9 9 0 9 1 11 2 1 15 13 11 2 11 2 11 2 11 7 11 2
21 9 9 13 9 0 9 9 11 11 1 10 9 1 11 2 11 7 11 0 9 2
8 3 15 9 4 13 9 9 2
30 13 13 2 16 9 9 0 0 9 1 9 0 0 11 13 1 15 2 16 4 4 0 9 1 0 2 0 11 13 2
17 0 11 3 13 3 1 9 2 0 1 9 1 0 9 1 11 2
5 13 15 9 11 2
23 12 9 0 11 13 3 1 0 9 11 12 9 7 0 12 13 2 1 15 7 10 9 2
36 0 9 13 0 13 9 0 9 11 2 9 2 1 10 9 1 9 2 16 10 0 9 4 13 7 4 13 3 9 11 1 9 9 0 11 2
24 13 15 1 11 9 9 7 9 11 11 7 11 11 1 9 1 0 9 0 9 11 11 11 2
23 9 9 1 9 9 1 11 4 13 9 1 0 7 0 9 2 13 0 9 9 11 11 2
23 10 9 4 1 11 7 11 13 2 16 13 10 9 0 9 7 13 15 0 9 2 13 2
16 0 9 0 9 11 11 13 1 9 13 9 0 9 0 9 2
15 11 13 1 9 0 9 11 2 15 13 9 10 9 9 2
4 11 13 14 0
4 11 2 11 2
30 1 9 1 9 0 9 0 9 13 1 0 9 9 11 0 9 9 1 9 11 2 11 2 11 11 0 9 11 11 2
13 1 9 3 13 2 16 1 15 7 11 13 9 2
42 0 9 2 15 14 11 11 13 2 13 1 15 2 16 15 13 13 15 2 15 15 13 1 9 2 7 16 13 9 2 15 4 15 13 13 0 0 9 1 9 9 2
8 1 0 9 13 0 0 9 2
16 16 4 7 13 1 11 2 13 4 1 15 9 2 13 11 2
8 16 9 13 0 9 11 11 2
29 3 13 11 1 9 11 7 0 9 1 15 2 16 13 1 11 2 15 13 1 0 9 1 9 1 9 0 9 2
8 1 9 1 9 9 13 1 9
9 11 11 2 0 9 0 9 11 11
61 9 11 11 2 9 0 9 0 9 2 15 1 11 1 12 2 12 2 13 2 16 9 9 1 0 0 9 4 13 9 9 3 12 9 2 7 15 3 2 16 9 0 0 0 9 13 9 3 0 2 3 7 0 1 9 1 9 0 9 12 2
20 13 13 2 16 9 11 0 0 9 4 13 3 10 9 1 9 0 0 9 2
17 3 13 0 0 9 0 9 9 0 9 13 3 1 9 1 0 2
51 1 0 9 7 13 0 9 2 7 15 3 13 9 7 9 0 2 0 2 0 7 3 2 0 9 1 9 9 12 2 12 2 1 0 9 9 1 9 2 12 7 1 9 0 9 1 9 7 9 12 2
24 9 4 13 13 9 1 0 9 1 9 7 9 9 0 9 1 0 9 7 1 9 0 9 2
24 13 4 13 1 0 0 9 0 7 0 9 2 16 4 4 1 0 9 13 0 9 7 9 2
54 7 3 4 15 13 13 9 1 9 7 0 0 9 1 0 9 2 0 9 9 0 9 4 1 0 9 3 13 2 2 7 1 9 9 1 3 0 9 2 9 2 0 9 2 9 2 1 9 2 9 2 9 0 2
41 16 13 1 9 1 0 9 2 1 9 13 1 9 2 16 1 0 9 15 0 9 13 2 0 13 15 7 1 9 10 9 1 9 9 12 2 7 1 0 2 2
35 3 0 0 9 0 1 9 1 9 0 16 11 2 11 2 11 2 11 2 11 2 7 3 0 9 11 2 11 2 11 0 2 3 13 2
26 1 9 12 13 16 2 3 0 2 9 11 2 7 11 2 2 11 7 0 9 0 15 1 0 9 2
7 13 4 13 0 0 9 2
21 13 2 3 0 0 9 11 7 11 7 0 0 11 2 7 11 3 2 2 13 2
25 3 15 13 9 2 3 13 13 7 11 2 16 15 13 14 11 7 1 0 9 3 3 14 11 2
6 13 7 1 9 11 2
24 3 7 9 12 13 9 2 9 2 1 0 9 9 0 9 9 2 12 1 9 2 9 2 2
21 3 3 2 16 4 9 9 9 2 9 2 9 2 9 2 13 3 0 2 0 2
60 3 15 1 0 9 2 15 9 11 13 16 0 9 2 7 7 1 0 9 14 13 2 16 0 3 0 9 4 3 13 1 0 9 2 13 2 9 9 16 0 9 9 2 9 2 9 2 9 2 0 2 7 14 0 2 7 15 2 0 2
17 0 4 13 2 16 9 1 0 9 13 15 7 0 2 7 0 2
15 13 15 14 9 9 0 7 0 0 9 1 0 0 9 2
34 9 7 9 15 13 3 15 2 13 14 1 15 2 16 15 13 13 2 16 15 13 1 9 7 1 0 9 2 7 1 9 7 9 2
19 0 9 1 0 9 0 0 9 4 13 0 2 16 4 4 13 9 0 2
24 7 16 0 2 1 9 1 9 0 15 1 9 2 12 1 9 0 9 13 13 7 1 9 2
34 7 7 3 0 0 9 13 3 0 9 0 9 2 9 2 0 9 1 9 7 0 0 9 1 0 9 7 0 9 1 9 0 9 2
9 9 9 2 9 0 2 7 0 2
9 11 11 2 9 2 0 9 7 9
24 3 16 13 0 9 2 4 15 13 2 16 12 1 0 9 1 10 0 9 13 2 0 9 2
13 1 9 9 15 0 9 9 9 13 3 15 13 2
10 1 15 1 9 0 15 3 3 13 2
12 1 9 9 9 3 14 0 9 7 0 9 2
15 0 15 0 9 9 2 16 3 15 13 2 1 15 13 2
28 13 15 3 0 9 9 1 9 1 9 7 16 15 13 9 1 9 2 15 13 1 9 7 1 15 15 0 2
28 0 9 13 9 1 9 1 10 9 2 16 15 13 1 10 0 9 7 13 1 15 9 1 9 1 0 9 2
14 13 1 15 2 16 4 15 3 3 15 1 9 13 2
19 9 13 9 2 13 15 16 0 3 0 9 7 9 1 15 1 0 9 2
8 3 1 15 13 2 3 13 2
41 9 1 0 9 0 9 2 11 12 2 12 2 2 1 9 9 1 0 9 13 1 9 1 9 9 9 2 3 13 14 0 9 2 16 15 13 1 9 0 2 2
24 16 1 9 0 11 13 3 13 9 0 2 9 13 10 9 0 9 9 9 1 9 1 9 2
17 10 0 9 3 13 0 0 9 2 3 13 2 14 1 9 0 2
41 13 15 0 16 13 1 9 2 1 9 9 1 15 9 2 16 13 3 0 2 10 0 9 15 13 2 9 1 0 9 2 0 9 0 9 7 9 0 0 9 2
14 1 0 9 15 13 1 12 3 0 9 1 9 9 2
20 0 2 9 9 2 15 13 9 0 2 0 2 9 9 2 9 0 2 0 2
22 0 13 9 0 2 0 7 15 2 2 0 13 0 7 13 9 3 2 1 0 9 2
9 0 9 9 13 2 0 13 9 2
41 0 13 9 2 0 13 0 2 1 9 0 9 2 0 9 7 9 13 1 9 13 15 1 10 0 9 1 0 9 2 3 2 9 9 9 1 9 0 9 2 2
28 9 2 0 9 7 9 1 0 0 7 0 9 9 2 0 3 7 3 2 13 13 1 0 9 1 0 9 2
27 9 9 2 9 7 9 15 13 1 0 9 1 0 2 0 7 0 9 7 13 13 9 3 0 1 9 2
59 16 15 13 3 1 9 0 15 9 1 9 9 9 2 3 0 9 2 2 2 13 4 9 0 2 0 7 0 2 16 3 1 9 2 0 2 0 9 1 0 9 7 9 16 0 9 9 1 15 2 15 4 1 9 3 7 3 13 2
8 7 1 15 0 9 3 13 2
9 0 9 1 0 9 13 13 1 9
9 11 11 2 9 9 2 9 7 9
22 1 9 0 9 1 10 9 0 3 13 9 1 0 0 9 2 15 15 4 3 13 2
14 1 0 9 4 0 9 13 9 9 7 13 0 9 2
25 13 7 0 2 16 12 1 9 9 12 2 1 15 0 9 13 3 0 9 2 13 9 0 9 2
35 9 1 15 7 15 7 1 0 9 0 9 4 3 1 9 9 12 13 1 0 0 9 2 1 12 1 0 0 9 2 15 4 3 13 2
18 9 9 1 0 9 4 13 7 0 9 10 9 13 1 9 0 9 2
39 9 0 12 9 13 9 7 9 15 0 9 7 3 13 1 9 3 13 9 9 7 9 0 9 2 10 0 0 9 7 9 1 9 7 9 10 0 9 2
34 1 9 9 13 13 2 16 15 13 13 1 9 2 3 9 13 3 10 0 9 2 9 9 2 7 9 15 3 13 1 10 0 9 2
19 0 9 9 1 10 9 13 9 13 0 9 0 9 7 3 13 0 9 2
12 12 1 0 9 13 3 9 1 9 7 9 2
17 0 9 2 3 15 9 0 9 9 13 2 13 9 9 0 9 2
44 16 4 3 13 1 9 0 9 2 0 4 15 13 2 16 0 9 13 1 0 9 7 9 0 9 0 3 0 3 0 0 0 9 1 0 9 7 13 1 15 9 0 9 2
14 1 15 13 9 13 9 0 9 7 1 0 0 9 2
15 3 1 9 0 9 4 13 13 3 1 0 7 0 9 2
12 0 9 7 0 9 13 0 0 9 0 9 2
9 3 15 13 13 9 13 0 9 2
16 0 0 9 4 13 13 0 9 3 1 9 1 10 0 9 2
27 9 10 0 9 13 13 9 9 2 13 9 1 0 9 2 7 13 3 10 9 1 9 9 1 9 9 2
32 16 3 4 13 2 1 9 1 0 9 15 1 9 0 9 13 2 16 4 9 0 9 13 14 9 2 7 7 0 0 9 2
19 3 15 1 9 9 13 12 9 2 7 0 9 9 2 7 10 9 9 2
14 13 0 3 13 1 0 9 9 0 7 9 9 0 2
14 0 9 4 13 0 9 9 9 9 2 0 9 9 2
27 1 0 9 4 3 0 9 13 9 9 2 9 0 9 4 13 13 0 9 0 9 7 0 0 0 9 2
10 9 13 1 9 13 0 9 0 9 2
15 3 13 13 9 0 9 9 3 0 9 1 9 9 9 2
21 13 15 3 13 3 0 9 7 13 15 9 7 9 14 0 2 7 9 3 0 2
15 1 9 7 9 9 0 9 4 13 0 0 9 0 9 2
20 3 15 13 0 9 2 15 15 3 1 0 9 13 1 0 9 1 0 9 2
30 9 0 9 2 0 1 0 9 1 0 0 9 2 13 0 9 1 9 0 9 0 9 7 0 0 9 0 0 9 2
17 9 4 13 3 9 0 9 7 9 13 9 9 7 0 9 9 2
17 0 0 9 0 9 13 9 9 7 0 9 2 9 9 0 9 2
13 9 9 13 9 0 9 7 9 0 9 0 9 2
12 0 0 9 13 7 1 0 0 9 0 9 2
10 13 9 9 2 13 15 10 0 9 2
18 1 0 9 13 9 9 9 2 7 3 0 9 2 16 15 13 3 2
10 0 9 9 13 9 9 9 1 9 2
10 1 0 9 13 9 9 9 9 13 2
15 9 3 13 9 9 7 1 9 9 2 9 7 9 9 2
26 13 3 0 9 13 9 9 9 16 9 2 16 4 13 1 9 0 9 0 9 7 0 0 9 9 2
11 9 13 9 9 1 9 0 9 0 9 2
11 3 15 3 13 9 0 9 7 0 9 2
40 1 0 9 15 13 9 9 9 7 9 2 9 9 15 13 1 3 12 2 12 9 2 16 15 13 9 1 0 9 7 9 1 9 9 1 0 9 1 15 2
26 3 9 9 1 9 9 15 13 1 9 10 9 1 9 2 15 13 13 9 1 0 9 3 12 9 2
9 3 15 13 7 9 7 9 9 2
39 9 9 1 9 0 9 15 13 1 9 9 13 7 13 9 1 10 9 2 15 4 3 13 13 1 9 9 1 0 9 7 1 10 0 9 1 10 9 2
16 9 9 15 13 7 9 0 9 2 15 7 13 9 10 9 2
39 0 9 4 13 4 13 1 0 9 7 13 4 13 0 9 9 1 10 9 7 9 2 1 15 1 0 9 13 7 9 7 9 9 7 0 9 9 9 2
10 13 9 0 9 1 12 0 9 13 0
3 9 11 11
10 9 15 13 2 9 15 13 2 2 2
3 9 11 11
4 9 13 10 9
16 1 9 0 9 7 0 9 13 1 9 0 9 1 12 0 9
2 11 11
32 16 15 9 0 9 13 0 9 0 9 1 0 9 1 11 2 15 1 9 14 13 2 16 3 1 12 9 13 10 9 0 2
13 9 4 3 13 1 9 0 9 0 0 0 9 2
39 10 9 15 1 9 12 13 3 1 9 2 13 15 2 15 15 15 13 2 7 3 15 3 13 1 10 9 2 3 15 13 9 0 9 7 0 9 9 2
33 3 0 0 9 7 10 0 9 13 3 1 9 3 2 0 9 3 13 7 3 3 15 1 0 9 1 0 9 13 7 0 9 2
17 1 9 12 15 9 13 0 9 7 9 1 10 9 3 15 13 2
33 1 9 3 0 0 9 9 9 9 11 13 1 9 2 7 1 9 12 15 13 14 15 2 0 9 3 13 1 9 0 0 9 2
13 9 15 13 14 1 9 0 0 9 1 9 12 2
25 0 9 13 7 9 0 0 9 9 11 13 2 16 15 1 3 0 0 9 1 0 9 13 4 2
3 13 3 13
7 15 15 7 3 13 9 2
33 1 9 1 3 0 11 3 15 1 3 12 9 9 1 9 7 9 9 7 9 10 9 13 10 9 2 0 9 2 9 7 9 2
46 16 3 3 13 1 10 9 1 0 9 2 13 9 13 13 7 1 10 9 2 15 13 0 9 1 3 12 9 2 3 3 2 9 11 13 12 9 2 2 7 13 7 13 1 9 2
22 13 15 3 7 13 2 16 9 9 13 0 9 7 13 13 1 0 9 0 0 9 2
23 1 9 2 1 0 9 2 15 3 13 9 0 9 2 3 0 0 9 2 7 9 9 2
56 9 9 11 2 11 2 11 2 7 11 2 11 2 11 2 11 2 3 13 2 16 15 2 15 13 1 9 3 13 12 0 9 10 0 9 2 7 3 7 10 9 2 13 1 15 1 9 0 3 14 0 0 9 7 9 2
2 0 9
21 3 15 3 13 9 0 9 0 9 9 1 0 9 2 15 7 9 0 9 13 2
49 7 9 3 1 9 7 12 13 2 16 1 10 9 3 13 9 0 9 7 9 1 0 9 7 0 9 2 15 1 9 9 11 2 11 2 1 9 12 2 12 2 3 13 0 0 9 9 0 2
19 9 10 9 13 3 2 7 0 0 9 1 9 7 0 9 1 9 12 2
64 0 9 15 7 9 9 3 13 2 16 3 0 9 9 12 13 0 9 7 15 7 0 0 9 2 9 0 7 11 2 9 2 0 2 12 7 12 2 7 12 9 9 1 0 9 2 9 2 0 2 12 7 12 2 15 13 9 9 7 0 9 0 9 2
20 15 15 3 2 3 16 0 9 2 13 13 7 10 9 15 13 16 0 9 2
12 7 15 3 13 1 9 0 2 11 10 9 2
2 9 13
36 3 3 9 13 7 9 11 13 1 9 12 0 9 1 0 9 1 9 0 9 1 9 9 7 0 9 2 11 2 13 7 9 0 9 2 2
37 13 4 13 4 1 12 2 9 12 2 7 15 7 1 0 9 0 0 9 9 1 9 9 2 12 7 12 1 0 9 1 9 11 1 10 9 2
31 9 2 1 15 9 13 1 12 9 9 9 2 3 13 3 2 16 13 0 9 2 13 15 0 9 7 13 9 7 9 2
24 0 9 0 9 0 9 3 13 9 7 1 0 9 9 13 3 9 0 9 9 7 0 9 2
34 1 9 9 2 12 2 3 13 9 11 0 9 2 13 7 10 9 9 2 11 11 2 1 15 4 15 13 1 9 0 9 0 9 2
3 9 13 9
13 0 9 9 13 13 12 0 9 1 9 0 9 2
42 0 1 9 4 13 1 15 1 3 12 12 9 13 10 9 2 9 2 9 2 9 2 15 3 3 10 9 2 9 1 9 2 0 9 7 9 2 13 9 2 11 2
12 1 10 0 9 7 1 15 9 13 3 4 2
24 16 15 15 1 0 9 13 2 9 0 0 7 0 9 1 0 2 3 0 9 13 10 9 2
18 1 15 2 16 4 1 11 7 1 9 11 13 10 9 2 13 9 2
31 9 7 4 13 10 0 9 2 7 1 9 1 9 9 4 13 1 12 7 1 3 2 3 14 7 1 9 1 0 9 2
24 16 10 9 13 3 16 1 12 2 9 0 2 4 15 10 9 3 13 16 1 0 0 9 2
31 0 9 0 9 13 7 3 14 12 9 2 9 0 1 9 2 3 1 0 9 2 2 16 13 0 1 9 1 0 9 2
12 15 13 1 9 0 9 2 15 7 3 13 2
21 1 9 13 1 0 9 10 0 9 2 0 9 7 0 9 1 0 9 7 9 2
37 1 10 9 4 15 1 9 2 11 13 13 2 10 9 4 13 9 9 2 3 3 13 7 14 0 2 16 13 3 0 2 0 7 0 1 9 2
4 1 9 13 9
11 10 0 0 9 7 9 1 0 9 13 2
20 3 1 0 0 9 1 9 9 0 1 11 9 15 13 0 2 0 2 9 2
38 10 0 9 4 13 13 0 9 1 0 0 9 2 16 3 0 9 13 0 9 1 0 9 2 1 9 13 1 11 7 9 15 3 13 1 0 9 2
10 7 1 0 0 9 7 9 15 13 2
25 9 4 13 13 3 2 16 9 13 3 3 7 9 1 3 0 9 1 9 4 9 9 3 13 2
10 16 3 13 9 2 13 9 2 11 2
10 7 1 0 9 13 1 0 9 9 2
21 3 12 12 9 15 3 13 2 0 3 9 12 12 13 1 9 0 9 1 11 2
22 13 9 1 3 0 9 2 16 13 15 1 0 9 1 11 2 14 1 0 9 13 2
4 1 0 9 9
20 16 4 15 0 9 1 9 9 3 3 13 2 4 0 0 9 13 14 9 2
17 0 9 13 9 9 1 9 12 0 9 2 15 13 1 0 9 2
37 1 9 9 11 4 13 4 13 3 9 1 9 2 3 4 1 1 0 0 9 13 13 7 0 9 16 1 9 2 3 9 1 9 3 1 12 2
20 9 13 1 15 3 0 2 13 7 9 2 11 0 9 0 9 9 1 9 2
10 3 3 0 9 13 14 9 0 9 2
12 3 15 4 3 1 9 9 13 9 0 9 2
25 9 0 7 0 7 13 3 13 2 7 3 1 0 9 9 13 9 1 9 0 9 7 13 15 2
26 7 1 9 15 13 13 15 2 3 14 13 0 9 7 9 15 4 13 3 13 2 13 9 2 11 2
5 9 2 7 9 2
19 16 9 13 0 9 0 9 9 1 0 9 2 13 1 9 1 11 9 2
7 10 9 15 7 13 0 2
20 0 0 9 4 3 0 9 13 3 3 1 9 2 16 4 15 3 15 13 2
26 16 0 0 9 1 9 12 3 3 13 2 7 13 1 0 9 2 13 15 13 13 1 0 9 11 2
28 9 15 7 1 9 1 0 9 0 9 13 3 2 7 13 9 9 2 15 13 2 16 13 3 0 9 13 2
17 16 15 13 2 16 14 2 13 15 0 9 2 13 9 2 11 2
20 0 9 15 3 13 1 9 12 2 12 2 13 15 1 9 7 13 9 9 2
12 13 2 14 0 2 9 13 7 1 9 13 2
25 9 3 14 1 9 9 13 2 9 15 13 1 0 9 2 7 13 15 7 0 0 9 2 2 2
3 0 0 9
20 1 9 0 9 13 1 0 9 3 12 12 9 0 0 0 9 1 9 9 2
9 15 15 13 2 13 9 2 11 2
18 1 0 0 9 15 9 13 13 14 0 9 7 13 15 1 15 9 2
16 0 9 13 0 1 9 2 7 4 15 3 13 2 2 2 2
12 9 0 9 9 13 0 9 1 9 11 11 2
17 7 15 1 0 9 1 9 9 13 1 0 9 7 0 0 9 2
30 0 13 2 16 3 13 1 9 9 10 9 2 16 9 13 3 3 2 16 15 13 7 0 9 13 9 1 0 9 2
20 9 3 4 3 13 2 13 7 13 1 9 2 3 4 9 12 9 9 13 2
21 1 9 9 13 4 3 13 2 7 3 3 16 0 9 0 1 0 9 1 9 2
21 1 9 2 3 15 0 9 13 2 14 4 3 13 7 13 15 13 1 10 9 2
22 1 9 2 11 15 3 1 9 0 9 13 2 3 13 3 2 16 9 3 13 9 2
44 12 9 2 15 13 13 9 9 1 9 0 9 11 2 15 13 2 16 1 9 9 4 1 0 9 13 0 9 1 9 2 15 4 13 3 2 9 4 13 7 13 9 9 2
22 3 15 15 14 15 13 2 15 13 0 9 0 0 9 2 15 2 15 15 13 13 2
21 16 15 1 15 15 13 13 1 9 9 2 13 0 2 16 13 13 13 2 13 2
62 1 9 9 0 9 15 13 13 0 2 7 0 9 1 9 9 9 12 2 9 7 3 2 16 9 0 9 4 13 16 0 7 13 14 0 9 2 9 11 13 13 9 15 12 9 14 13 2 7 3 3 13 2 16 4 0 9 0 9 9 13 2
5 9 9 13 1 9
27 0 0 9 3 1 15 15 3 13 9 2 16 3 13 10 9 0 7 0 0 9 7 13 9 1 9 2
15 0 9 1 11 12 13 10 9 1 9 9 9 0 9 2
46 9 0 9 1 11 2 1 0 9 7 1 11 15 7 3 13 2 7 3 0 9 13 1 9 7 13 15 1 9 13 0 9 1 12 0 9 2 12 9 5 12 9 12 9 2 2
25 1 15 7 13 2 16 13 2 14 15 1 9 9 0 9 0 9 2 13 15 12 9 0 9 2
15 3 13 0 9 0 2 0 0 9 2 13 9 2 11 2
34 10 9 13 0 2 1 10 9 13 1 0 9 2 1 9 13 9 2 9 9 3 13 1 9 2 3 15 13 1 15 1 0 9 2
12 3 3 15 9 13 2 16 1 15 13 13 2
21 9 0 9 1 12 9 13 0 2 9 9 9 1 9 12 9 7 9 12 9 2
11 3 3 9 2 7 1 0 9 0 9 2
20 13 10 9 1 0 7 0 9 1 9 13 2 13 3 3 0 9 2 2 2
3 9 1 9
27 3 16 0 9 9 1 0 0 9 13 1 9 2 3 1 9 0 9 0 11 1 11 2 0 9 9 2
30 13 3 9 3 0 2 3 0 2 16 15 1 9 0 2 9 9 13 13 9 2 3 0 9 13 3 1 9 0 2
25 3 13 2 16 13 3 15 1 10 2 16 4 0 9 1 0 9 13 1 9 9 3 0 0 2
25 13 2 14 15 0 9 3 1 0 9 12 2 0 9 0 1 9 12 15 15 13 14 0 9 2
17 0 0 9 3 13 3 1 9 0 1 9 12 7 1 0 9 2
3 0 9 9
1 9
18 9 2 9 11 11 2 12 2 12 2 13 1 0 1 0 0 9 2
20 1 0 7 0 9 7 1 11 3 13 2 10 0 9 15 13 3 1 9 2
16 0 0 0 0 9 13 0 9 0 9 1 0 9 1 11 2
7 11 11 13 9 0 9 2
8 0 2 0 2 0 7 0 2
18 3 9 0 2 13 1 9 15 2 0 9 2 7 2 0 9 2 2
8 13 0 7 0 1 9 9 2
14 1 0 9 13 1 0 9 9 7 9 13 3 13 2
16 1 9 13 1 11 7 13 15 9 11 11 1 0 9 0 2
15 3 15 13 1 9 2 1 15 1 9 12 13 9 9 2
19 9 13 0 3 1 0 0 9 2 10 9 7 13 9 7 9 0 9 2
11 10 9 1 0 9 13 0 9 0 9 2
8 0 9 9 13 0 0 9 2
64 9 0 9 0 15 10 9 7 9 10 9 2 9 0 0 0 9 0 7 0 2 15 13 0 9 2 13 15 13 15 1 15 2 13 15 3 7 13 1 9 0 0 9 7 15 13 9 2 1 9 2 16 7 16 4 13 15 2 13 0 13 3 15 2
7 9 13 9 0 0 9 2
23 13 10 9 1 9 2 10 9 1 9 2 9 9 2 2 9 2 1 15 15 3 13 2
9 11 15 3 13 1 3 0 9 2
15 13 1 0 9 9 2 13 3 0 2 16 16 4 13 2
11 1 0 9 7 10 9 13 0 0 9 2
23 13 15 1 9 9 1 0 9 7 1 0 7 0 9 1 9 0 2 9 9 3 0 2
22 7 1 9 9 11 13 9 0 9 2 1 10 0 9 13 0 9 9 7 0 9 2
5 13 9 0 9 2
14 1 15 13 0 9 0 9 7 9 0 9 0 9 2
34 1 0 9 1 9 2 15 15 13 1 0 9 2 13 9 1 0 9 7 9 9 2 9 1 9 2 9 2 9 1 0 9 2 2
17 11 11 13 1 9 12 2 3 1 9 0 2 1 9 0 9 2
9 10 9 13 9 1 0 0 9 2
2 11 11
3 11 11 2
11 9 2 9 2 9 2 9 12 2 12 2
4 9 11 11 2
6 0 9 2 0 9 2
8 12 2 9 2 12 2 9 2
2 11 11
2 9 11
4 9 13 0 9
2 11 2
27 1 9 13 1 0 9 2 11 2 9 0 9 7 9 2 10 0 9 13 9 2 9 7 9 0 9 2
14 13 15 7 0 0 9 11 1 0 9 1 0 9 2
18 1 10 0 9 11 11 15 3 3 13 7 13 9 0 1 0 9 2
29 1 9 9 3 2 13 0 9 1 9 7 9 0 0 9 11 2 11 7 1 9 7 9 0 9 1 0 11 2
36 13 15 7 0 2 0 9 1 9 0 9 1 9 11 2 0 9 7 11 2 0 9 2 15 4 13 1 9 1 0 9 7 0 0 9 2
17 1 0 9 13 3 13 3 12 9 9 1 0 9 11 2 11 2
9 13 13 3 9 9 11 2 11 2
12 13 15 7 1 9 0 0 9 1 10 9 2
20 0 9 3 13 13 2 7 15 3 12 9 2 3 0 9 1 0 0 9 2
14 9 4 15 13 13 15 2 7 15 3 13 0 9 2
21 11 13 9 2 1 15 13 3 13 0 9 9 1 0 9 1 9 1 10 9 2
13 1 10 9 13 1 11 2 11 9 10 0 9 2
13 1 9 9 11 13 0 9 0 9 0 0 9 2
20 13 3 1 0 7 0 9 2 7 3 3 1 0 9 0 7 1 0 9 2
3 0 0 9
1 9
19 9 2 9 7 9 9 11 11 2 12 2 12 2 13 3 0 7 0 2
20 3 13 15 7 1 9 0 9 11 11 2 10 0 0 9 13 3 1 9 2
15 13 1 9 2 15 1 15 3 13 1 9 0 0 9 2
9 15 13 9 0 9 1 12 9 2
21 3 15 13 9 13 9 1 0 9 0 0 9 2 9 7 9 0 9 0 11 2
11 3 7 3 0 9 13 1 9 0 9 2
16 9 11 11 13 2 1 0 9 2 1 11 3 9 16 9 2
30 1 3 0 9 1 0 0 9 2 1 9 9 7 9 15 13 1 9 0 9 10 12 9 2 7 7 9 0 9 2
8 10 0 9 13 1 9 9 2
12 3 0 9 13 3 0 9 1 10 0 9 2
31 13 15 9 2 15 15 1 9 12 1 9 13 0 9 16 9 0 0 9 2 16 3 0 9 7 3 7 3 0 9 2
26 0 13 14 0 0 9 2 7 7 0 0 0 9 2 3 16 3 0 9 7 3 0 9 0 9 2
22 15 15 1 0 9 3 3 13 3 9 11 11 11 2 9 11 11 7 9 11 11 2
15 3 1 0 9 4 13 0 9 0 2 0 9 11 11 2
14 11 11 9 11 13 1 0 9 0 9 3 0 9 2
20 9 13 7 1 9 12 9 13 1 0 0 9 7 1 0 0 7 0 9 2
7 7 13 1 9 3 0 2
8 11 11 11 11 2 11 11 2
10 9 7 9 0 11 2 9 11 11 2
8 12 9 2 13 11 2 12 2
2 9 9
1 9
45 9 2 13 0 13 15 11 11 2 12 2 12 2 13 2 10 9 15 10 9 3 13 2 3 15 13 2 7 13 0 9 0 9 2 15 13 11 12 1 9 9 0 9 9 2
17 3 13 10 9 10 0 9 1 15 2 15 3 13 10 9 9 2
19 13 15 7 0 9 1 0 9 0 9 2 9 2 9 2 9 11 2 2
24 9 13 0 9 1 11 1 11 0 9 9 2 9 15 13 9 7 9 11 2 9 2 9 2
18 16 9 0 2 13 1 3 0 11 13 0 2 3 3 7 15 0 2
17 3 10 9 2 15 13 10 0 7 3 7 0 9 3 0 9 2
16 9 9 13 9 2 0 9 3 0 7 3 0 9 0 9 2
21 11 15 13 1 9 9 7 0 9 2 9 2 15 15 13 3 1 9 9 2 2
23 9 16 9 1 0 9 1 12 9 13 15 0 16 9 2 9 2 9 1 9 7 9 2
22 1 0 9 7 2 1 11 2 3 9 2 15 13 9 2 0 9 2 15 15 13 2
27 13 15 3 9 0 2 7 13 15 9 13 9 9 2 1 1 15 13 0 13 7 13 0 7 0 9 2
19 9 13 3 9 9 2 1 15 4 9 3 3 3 13 2 13 2 13 2
17 7 13 2 14 11 1 9 16 3 0 2 13 2 3 2 9 2
27 13 1 9 7 9 2 15 13 3 9 1 9 0 0 9 2 15 2 15 10 9 3 13 16 10 9 2
14 0 9 13 13 0 9 7 9 2 15 13 9 9 2
18 10 0 9 13 1 15 2 16 15 13 3 2 3 4 15 3 13 2
30 3 13 2 14 9 9 1 0 9 2 7 2 16 13 15 1 9 15 13 9 2 16 13 9 16 3 0 9 9 2
21 3 13 3 0 7 0 9 0 9 2 15 13 0 7 3 1 9 13 10 9 2
22 9 15 13 7 0 9 9 2 1 15 11 3 1 0 9 13 2 15 13 9 9 2
45 13 2 14 9 9 2 0 9 2 13 15 14 3 13 15 2 15 15 13 2 0 9 9 2 15 13 9 1 10 9 2 10 9 2 2 2 2 2 2 3 16 1 10 9 2
12 7 15 15 13 9 2 13 2 14 10 9 2
10 9 15 2 16 9 10 0 9 13 2
4 11 11 9 2
9 11 11 2 9 2 9 2 9 2
12 13 9 11 2 9 9 7 9 2 11 12 2
7 13 7 9 13 11 11 2
8 12 9 2 9 7 9 13 2
5 9 1 11 11 13
21 9 0 9 11 11 11 13 2 16 4 13 1 10 9 1 0 9 1 11 11 2
14 0 9 10 9 13 1 9 12 3 1 10 0 9 2
37 1 9 0 0 9 0 1 9 2 15 15 13 4 13 2 13 11 3 13 1 9 0 9 1 11 7 3 13 1 9 10 9 1 0 9 3 2
22 0 0 9 2 15 13 1 9 0 9 2 13 9 9 13 3 2 13 3 11 11 2
31 1 11 1 9 2 12 13 3 9 11 7 10 9 2 12 2 2 9 2 12 2 7 9 9 7 0 9 2 12 2 2
17 9 9 13 3 13 1 9 9 12 2 1 11 1 11 9 12 2
3 2 11 2
8 0 0 9 13 7 0 0 9
13 0 0 0 9 4 3 3 13 1 0 9 9 2
47 9 7 0 9 1 0 7 0 9 15 13 1 9 13 1 0 9 0 9 7 9 2 0 7 0 9 2 0 9 7 9 1 0 9 7 9 9 7 1 0 9 7 1 9 0 9 2
14 1 12 9 0 1 12 9 0 9 13 7 0 11 2
27 10 9 10 9 13 1 9 0 9 9 11 11 1 0 9 10 0 9 2 3 0 9 1 0 0 9 2
20 3 1 0 9 13 1 9 0 9 0 9 11 7 0 0 0 9 9 11 2
36 13 13 7 0 0 9 0 0 7 0 0 2 0 7 0 9 7 9 1 9 2 1 9 1 0 9 2 9 9 2 9 7 9 0 9 2
16 0 9 9 13 3 0 0 9 0 0 9 0 1 0 9 2
9 10 9 13 11 11 1 0 11 2
6 11 13 9 0 0 9
32 0 0 9 11 11 7 0 9 11 11 15 13 13 9 9 9 0 2 11 2 15 12 2 9 13 9 0 0 9 1 11 2
18 1 9 2 15 13 1 12 2 9 2 13 9 9 9 11 7 11 2
20 10 9 15 13 9 0 9 11 11 2 15 15 7 1 9 11 1 9 13 2
8 9 0 9 13 1 9 10 2
29 13 4 2 16 4 15 15 10 13 9 7 13 1 9 0 9 0 9 1 11 2 13 0 9 0 9 11 11 2
18 13 2 16 13 1 0 9 2 9 1 0 9 13 13 0 12 9 2
1 3
22 0 0 9 11 11 4 1 9 13 1 9 0 0 9 1 0 9 1 0 0 9 2
20 9 2 1 15 15 9 13 10 9 2 9 7 9 2 13 1 12 2 9 2
25 9 9 9 9 11 11 13 3 1 12 9 1 0 0 9 1 0 9 12 9 7 9 11 11 2
16 9 1 9 13 3 3 0 9 0 9 2 0 9 11 11 2
4 9 1 9 2
1 9
2 11 11
28 0 12 2 0 0 9 10 9 2 0 7 0 9 7 10 0 9 2 15 0 9 1 0 9 13 0 9 2
22 10 9 15 13 0 3 0 9 2 0 3 0 7 1 9 3 0 0 9 1 11 2
23 15 2 3 16 10 0 0 9 1 9 2 13 10 9 1 9 2 0 9 7 0 9 2
24 0 12 15 13 13 11 16 9 1 0 9 0 0 9 2 15 15 3 1 0 9 3 13 2
22 15 13 7 9 9 9 1 0 9 11 2 11 2 7 11 2 2 0 1 0 9 2
37 1 9 0 9 11 11 13 13 0 12 1 11 0 7 15 2 16 3 10 0 0 9 13 2 3 14 1 10 9 7 9 2 15 13 0 12 2
24 9 0 9 2 10 0 9 13 1 9 9 9 0 9 2 13 13 3 1 9 7 0 9 2
39 10 9 13 3 3 1 9 13 0 9 2 7 13 3 9 9 2 16 0 7 0 9 0 9 0 12 15 3 13 13 0 16 10 0 0 9 2 9 2
42 1 9 2 3 15 1 9 0 12 13 3 0 9 9 9 2 3 2 9 2 9 7 9 2 15 0 9 10 9 7 9 3 13 7 9 15 13 3 1 0 9 2
52 1 9 7 9 2 3 15 13 3 9 9 9 2 7 9 0 9 7 0 9 1 9 0 9 15 3 0 9 0 9 13 3 1 0 0 7 0 0 9 2 0 0 9 7 3 9 1 9 1 11 2 2
26 1 10 9 13 3 0 13 2 15 15 4 13 1 0 0 9 0 12 2 15 13 1 11 1 11 2
29 1 0 9 13 4 13 3 3 1 9 2 7 1 9 2 15 0 12 13 2 3 13 9 3 14 0 9 11 2
8 0 9 13 1 9 1 0 11
29 0 9 13 0 0 0 9 2 15 1 0 11 1 11 13 1 9 12 2 9 7 13 14 1 9 12 2 9 2
22 9 4 13 13 1 0 9 9 0 0 9 2 11 12 2 11 0 0 7 9 11 2
13 11 11 13 1 10 0 0 9 1 0 9 11 2
12 12 1 10 9 13 7 0 9 1 0 11 2
24 1 9 12 2 1 10 12 12 9 2 13 1 9 9 11 1 11 7 13 15 9 10 9 2
19 1 0 0 0 9 1 0 11 13 10 0 9 2 15 4 13 16 0 2
23 3 1 10 9 13 9 1 0 0 0 9 2 15 3 1 9 0 11 0 0 9 13 2
14 9 13 3 12 1 0 9 1 15 2 7 16 0 2
12 1 9 12 13 9 0 9 0 9 11 11 2
27 9 1 0 9 9 1 0 9 12 2 7 12 2 9 13 9 9 1 9 0 9 1 0 0 0 9 2
16 0 9 0 9 15 13 9 9 9 7 9 9 0 0 9 2
19 9 9 1 9 9 1 0 9 3 3 13 1 9 3 0 9 0 9 2
3 2 11 2
23 9 9 0 2 9 2 11 11 4 13 1 0 9 11 1 0 0 9 1 11 0 9 2
2 9 11
11 11 11 7 11 11 1 0 9 9 13 9
2 9 11
9 11 11 13 1 9 1 9 3 9
5 9 11 11 2 11
8 9 2 9 7 9 1 9 9
2 11 11
34 3 3 2 12 9 2 2 13 1 0 9 9 0 9 0 0 9 9 1 9 2 10 9 1 9 12 13 10 9 0 9 1 9 2
27 0 9 13 11 11 2 12 2 2 15 3 13 16 9 12 1 0 9 11 2 0 1 0 0 9 2 2
13 3 4 15 13 13 7 13 9 0 3 12 9 2
18 9 1 9 4 3 3 16 1 12 9 13 13 16 9 1 0 9 2
20 3 3 13 10 9 1 11 11 7 1 9 4 15 3 13 7 1 9 11 2
14 3 3 4 14 3 13 7 13 9 13 9 16 9 2
27 3 3 4 7 13 2 16 15 3 13 2 7 13 15 1 0 9 0 9 2 0 1 9 1 0 9 2
15 13 4 15 3 3 13 1 9 9 7 9 1 0 9 2
21 9 11 11 15 13 0 0 9 1 0 9 7 9 2 3 13 7 9 7 9 2
10 3 4 14 13 13 7 9 0 9 2
18 13 15 3 0 2 9 13 1 9 0 9 1 0 9 1 9 2 2
27 0 9 15 13 3 9 9 2 1 10 9 3 13 7 0 9 0 1 0 9 1 11 1 11 2 2 2
25 1 11 11 7 11 11 4 15 1 0 9 13 3 0 7 9 0 0 9 11 11 15 13 3 2
21 1 9 3 4 7 13 3 3 3 2 9 0 9 13 0 7 0 9 13 0 2
22 9 1 9 4 15 3 0 13 3 13 3 1 9 2 3 3 1 9 2 2 2 2
15 13 15 1 9 9 2 16 9 10 9 13 3 0 9 2
6 15 15 3 3 13 2
23 10 9 13 1 15 0 9 3 2 1 10 9 7 9 2 1 10 0 9 1 9 9 2
21 3 1 9 4 15 13 2 16 13 0 9 3 10 9 3 0 2 0 7 0 2
27 13 9 1 0 9 0 9 2 0 9 2 0 9 7 0 10 10 0 9 7 13 15 15 9 2 2 2
12 10 9 13 0 2 3 16 13 0 10 9 2
14 3 10 9 9 7 0 9 3 13 1 0 9 3 2
13 7 1 10 3 0 9 4 1 9 13 0 9 2
8 9 9 13 13 3 0 9 3
7 11 2 11 2 11 2 2
28 9 9 3 13 9 2 15 4 13 2 16 13 0 7 3 13 9 1 9 12 9 0 0 9 2 11 2 2
13 10 9 13 1 10 15 0 9 1 9 9 11 2
51 9 2 10 0 9 15 13 1 12 9 2 9 2 1 12 9 2 13 0 9 0 2 9 2 11 2 0 9 2 15 1 0 9 13 11 2 11 2 9 0 9 2 0 9 2 1 9 0 9 11 2
14 9 1 9 1 11 13 9 11 11 2 11 1 0 2
25 9 11 3 13 2 16 4 9 16 9 11 13 9 13 2 16 1 10 9 4 13 0 9 9 2
40 11 2 11 2 9 9 11 11 12 2 1 15 13 0 9 1 9 2 3 13 2 16 11 15 13 0 9 7 13 9 9 1 11 3 3 7 3 13 1 2
9 10 9 13 11 2 11 1 0 2
22 9 15 13 2 16 1 9 13 0 9 2 16 9 9 13 2 16 9 4 13 13 2
8 9 1 9 15 13 14 1 9
5 11 2 11 2 2
30 1 0 9 9 2 7 13 3 0 2 13 9 9 1 9 9 9 0 9 2 15 15 1 0 11 13 1 0 9 2
8 11 15 13 0 9 10 9 2
15 9 3 13 0 9 2 9 15 13 3 7 9 9 9 2
25 10 0 9 0 11 2 15 0 9 11 11 13 2 13 3 1 0 9 9 1 9 0 9 9 2
19 1 10 9 7 9 3 13 7 13 4 3 3 2 16 4 1 9 13 2
21 9 9 13 9 3 2 0 9 3 13 1 9 9 2 16 1 0 9 0 9 2
22 0 9 15 13 7 1 9 0 9 2 16 15 1 15 13 9 0 9 1 0 9 2
28 0 9 13 1 9 11 9 2 15 1 9 9 13 9 7 9 1 11 2 9 1 11 7 0 9 1 9 2
30 0 9 13 0 0 9 2 15 15 13 3 1 9 13 9 1 9 0 9 2 16 4 1 15 13 10 0 0 9 2
8 10 9 3 1 15 13 9 2
12 0 9 15 3 1 9 13 13 9 1 9 2
22 1 9 11 2 16 15 10 9 15 13 2 9 9 9 13 2 16 15 13 0 9 2
3 3 3 2
5 9 1 9 7 9
13 11 15 13 13 2 7 0 9 13 1 0 9 3
7 11 2 11 2 11 2 2
9 11 13 1 9 9 11 7 11 2
6 3 13 3 3 3 2
13 9 13 3 3 2 9 13 12 9 7 12 9 2
15 10 9 13 9 9 2 16 9 13 2 16 13 0 9 2
42 1 9 4 13 1 9 1 9 12 9 12 9 1 9 9 2 13 9 11 11 2 4 13 7 3 4 15 13 2 16 0 11 13 12 9 9 1 9 9 1 9 2
9 15 15 13 3 2 16 2 2 2
7 1 9 3 9 3 13 2
24 9 9 15 13 2 7 16 3 14 15 2 1 9 7 13 3 7 9 13 13 1 0 9 2
22 3 13 15 1 9 2 1 9 13 12 9 2 15 1 0 9 13 0 14 1 9 2
8 16 13 2 13 15 13 3 2
10 3 9 13 1 0 9 0 9 11 2
27 3 15 13 0 9 7 9 13 0 9 13 2 15 15 13 2 13 1 9 7 13 1 12 9 0 11 2
8 15 2 16 13 0 0 9 2
13 9 0 9 11 11 11 9 9 13 3 1 9 2
27 13 2 16 9 13 7 0 9 2 3 9 13 2 1 1 15 2 16 0 9 1 9 13 14 0 9 2
15 7 15 7 13 2 16 9 9 9 1 9 0 9 13 2
15 9 9 1 0 9 2 15 13 2 15 3 13 9 9 2
14 10 9 2 12 1 12 9 9 2 15 13 0 9 2
9 9 13 1 9 9 11 3 3 2
5 11 13 7 0 2
19 9 0 9 13 2 9 13 2 16 15 9 14 13 2 16 4 3 13 2
7 1 0 9 13 3 9 2
12 3 13 0 2 3 15 13 2 3 0 9 2
7 9 1 0 9 13 0 9
5 11 2 11 2 2
23 0 12 9 9 9 0 0 0 9 2 11 2 1 0 12 9 0 9 13 1 0 9 2
6 3 15 13 12 9 2
22 1 9 12 13 11 1 12 12 9 2 3 1 9 1 9 9 3 3 16 12 9 2
22 9 11 11 11 3 13 2 16 0 9 13 0 0 9 15 0 9 0 1 0 9 2
7 9 9 13 1 12 9 2
16 1 11 13 12 0 9 2 3 1 11 2 3 15 13 12 2
23 9 0 9 4 13 4 3 13 7 1 9 1 9 9 2 7 1 0 9 2 13 11 2
19 0 1 0 7 0 9 13 1 3 0 9 9 2 15 3 13 0 9 2
20 1 9 13 11 9 0 9 2 15 13 13 1 0 9 0 0 7 0 9 2
15 0 9 13 1 0 11 2 3 15 13 1 15 9 11 2
23 1 12 9 13 1 0 9 0 9 1 11 11 7 0 9 2 15 13 3 0 9 9 2
4 0 9 1 11
7 11 2 9 0 11 2 2
9 1 11 11 15 4 3 13 15 2
13 16 4 15 15 15 13 2 13 4 15 3 15 2
1 3
30 0 9 9 7 0 9 13 1 9 7 9 0 9 1 0 9 3 1 12 1 12 9 2 9 2 3 1 12 9 2
9 9 13 9 9 1 9 0 9 2
37 9 1 9 9 11 11 13 9 0 9 9 0 9 11 11 2 15 13 9 1 9 0 9 1 0 9 2 0 11 0 11 7 0 0 0 11 2
14 0 9 4 13 0 9 1 9 0 9 7 0 9 2
3 2 11 2
20 9 13 1 9 1 0 9 9 0 9 12 9 1 9 2 13 9 0 11 2
14 9 1 9 0 0 9 13 1 9 1 0 9 9 2
18 9 13 9 3 1 9 2 1 10 9 15 13 1 3 16 12 9 2
4 9 2 15 13
2 11 11
4 13 0 9 2
3 10 9 2
5 9 2 15 13 2
21 9 2 1 15 15 13 2 9 2 15 13 2 9 2 15 15 3 13 1 9 2
8 7 14 1 15 15 13 13 2
18 16 15 9 1 9 13 2 13 15 7 13 2 13 4 15 0 9 2
26 16 1 15 1 9 13 9 2 13 15 1 9 7 13 15 9 2 13 4 1 15 2 15 13 11 2
8 15 4 15 3 9 13 13 2
13 16 4 15 2 0 9 2 3 3 13 1 9 2
17 1 0 9 2 15 4 1 9 13 2 15 15 15 13 14 6 2
6 10 0 9 13 15 2
14 7 9 1 9 2 3 15 0 2 1 9 2 0 2
6 15 15 13 14 3 2
21 9 15 3 3 13 2 15 4 1 15 3 1 9 13 2 16 4 15 13 13 2
16 1 0 9 1 0 0 11 15 1 10 9 13 0 9 9 2
15 1 9 15 1 10 9 13 9 2 15 9 13 0 9 2
12 9 2 3 15 13 9 2 13 9 0 9 2
16 9 2 13 15 1 15 9 0 15 9 2 13 1 9 9 2
7 16 4 14 9 2 9 2
10 3 15 13 9 9 2 3 1 9 2
14 9 9 2 16 1 0 9 3 13 9 2 3 13 2
10 16 15 1 9 13 0 2 13 9 2
6 15 13 7 13 9 2
5 9 13 3 0 2
5 9 13 10 9 2
5 3 4 15 13 2
5 13 15 1 9 2
3 1 9 2
7 15 10 9 2 13 15 2
7 3 15 13 2 13 9 2
7 3 14 4 13 1 9 2
5 15 13 1 9 2
2 13 2
4 7 15 9 2
5 15 15 13 13 2
15 0 9 13 15 2 15 13 3 2 13 3 9 0 9 2
26 10 9 9 3 13 7 13 15 15 1 0 9 2 0 9 13 15 2 15 13 13 2 15 15 13 2
7 7 9 1 9 1 9 2
10 1 9 3 2 16 4 9 9 13 2
4 9 1 9 11
2 11 2
29 9 1 0 9 11 2 15 13 9 12 9 9 2 1 0 9 7 0 9 4 13 9 9 13 9 9 7 9 2
11 13 15 3 9 1 9 11 11 11 11 2
22 1 15 9 13 9 1 0 9 1 9 10 0 9 2 16 1 0 9 13 10 9 2
30 9 7 1 0 9 0 9 9 9 2 9 7 9 11 11 4 13 1 9 1 11 11 7 0 11 1 0 9 11 2
20 9 1 15 13 3 1 9 9 9 12 9 2 16 13 9 1 0 9 9 2
6 9 1 9 3 3 3
5 11 2 11 2 2
38 16 4 15 13 1 0 9 0 9 0 9 3 13 9 3 12 0 9 2 13 9 0 9 9 0 9 11 11 2 16 4 4 10 9 13 0 9 2
23 13 2 14 15 7 14 9 9 2 13 4 4 1 15 9 10 9 13 14 1 0 9 2
25 11 2 11 3 1 9 1 11 3 3 13 10 9 2 1 15 13 0 9 1 0 7 0 9 2
21 1 10 9 13 3 3 0 9 10 2 16 9 10 9 0 9 4 13 3 0 2
15 1 0 9 13 2 16 1 0 9 4 3 13 12 9 2
14 9 1 9 9 0 9 13 9 9 1 9 9 9 2
24 1 0 9 13 3 0 13 0 0 9 2 15 9 13 3 0 16 0 9 1 9 0 9 2
21 14 15 0 9 15 1 11 2 11 3 13 1 9 9 2 16 15 15 9 13 2
14 13 2 14 15 1 0 9 2 13 4 13 0 9 2
10 3 1 0 9 13 9 1 0 9 2
14 9 9 7 3 13 3 0 9 16 1 3 0 9 2
15 9 9 1 11 2 11 2 7 11 2 1 9 2 9 2
4 11 13 1 11
5 11 2 11 2 2
14 0 12 2 0 0 9 11 12 4 3 13 1 11 2
22 10 9 13 3 9 0 9 7 9 2 15 13 3 13 9 1 0 0 9 1 11 2
32 1 12 9 9 1 11 2 11 7 0 12 9 13 3 11 11 2 15 1 10 9 13 9 1 12 9 1 11 14 1 11 2
30 13 1 9 0 9 2 16 13 15 2 7 13 0 9 1 0 9 1 11 2 16 13 15 2 13 1 9 9 9 2
9 13 15 7 9 11 11 1 11 2
5 0 0 9 13 9
5 11 2 11 2 2
19 1 0 0 0 2 9 2 13 0 2 16 4 13 0 9 1 3 9 2
39 1 0 9 15 13 12 9 9 11 2 9 13 1 0 0 7 0 9 7 3 16 12 9 9 13 12 1 12 0 0 9 3 1 9 11 11 2 11 2
21 1 9 13 10 9 1 11 1 11 1 9 0 9 1 11 7 1 11 0 9 2
26 1 10 9 15 13 9 13 1 9 9 0 9 1 11 2 9 11 2 7 1 0 11 2 11 2 2
28 16 13 11 0 9 11 11 2 11 2 10 9 13 1 11 0 2 15 1 15 13 1 9 1 0 0 9 2
16 3 11 13 1 11 12 9 9 1 11 7 0 9 1 11 2
26 13 1 15 16 0 9 11 2 7 3 9 1 9 0 9 1 11 1 11 2 15 13 1 9 11 2
5 9 0 9 13 13
2 11 2
32 9 9 9 0 9 0 9 11 2 11 2 7 0 0 9 2 11 2 2 0 3 1 9 2 13 1 9 11 11 11 13 2
31 3 9 2 16 15 9 0 9 12 9 13 1 9 10 9 2 3 13 2 16 13 10 9 3 0 2 13 3 9 11 2
15 16 9 0 9 11 13 0 9 0 15 9 12 0 9 2
20 13 9 2 16 4 1 0 9 9 9 13 9 0 15 0 9 1 0 9 2
34 9 11 3 13 2 16 4 9 1 0 9 1 11 7 11 2 10 9 3 13 1 9 11 2 13 9 1 0 9 9 12 0 9 2
38 1 9 2 3 4 9 0 9 13 0 0 9 0 9 1 11 7 11 7 0 0 9 2 9 11 13 2 16 1 0 9 4 15 13 1 9 0 2
31 1 1 15 2 16 0 9 3 13 0 9 12 9 9 1 0 9 2 4 15 15 3 13 7 1 9 0 9 2 13 2
7 11 13 9 1 9 1 11
2 11 11
36 16 9 10 0 9 1 0 9 10 9 13 1 0 9 9 0 9 1 12 5 2 13 11 3 1 11 7 11 1 9 1 0 9 10 9 2
11 9 9 1 11 3 13 1 0 12 5 2
36 10 9 13 3 1 9 0 9 0 0 0 0 9 11 11 2 11 2 16 15 1 10 9 1 9 11 11 13 1 0 9 9 1 12 9 2
15 11 13 0 9 1 9 2 10 9 3 7 3 13 13 2
14 10 9 1 9 1 15 13 13 7 1 15 3 0 2
6 3 7 0 9 13 2
28 9 1 11 15 1 10 9 13 1 9 9 1 9 0 9 2 3 3 3 13 11 2 11 2 11 7 11 2
42 3 13 11 1 10 9 9 1 0 12 9 9 9 1 9 12 9 2 9 7 10 9 1 10 9 1 0 9 13 1 12 5 2 16 9 1 15 13 1 12 12 2
19 3 3 15 10 9 13 15 13 2 7 1 0 9 1 10 9 9 13 2
11 3 13 1 15 3 0 9 2 0 9 2
19 1 9 15 3 13 11 2 3 4 13 0 0 9 2 9 7 0 9 2
40 9 1 0 9 1 10 9 3 11 13 2 16 10 9 1 0 9 9 2 0 2 11 2 11 2 0 11 2 11 7 11 2 13 1 10 9 1 12 5 2
53 1 11 11 2 9 9 11 2 1 9 0 9 9 9 7 9 13 9 1 15 2 16 9 9 2 15 1 11 13 2 10 9 13 13 9 1 11 2 10 0 9 13 0 9 11 7 1 0 2 7 0 9 2
16 0 9 2 9 7 9 2 15 3 13 2 13 3 0 9 2
18 3 1 9 1 9 1 0 0 9 13 9 0 0 7 9 3 0 2
19 1 9 0 9 7 9 0 9 4 1 15 11 0 13 0 9 7 9 2
17 9 9 10 9 0 9 13 2 16 14 0 2 7 3 3 0 2
17 3 15 13 1 9 12 9 1 12 9 1 9 1 11 2 11 2
24 3 2 16 15 13 13 1 12 2 9 2 3 15 11 0 9 13 1 9 0 9 7 9 2
17 1 15 4 1 9 1 11 13 9 10 9 2 15 13 11 11 2
3 0 9 11
4 11 1 11 2
10 13 10 0 9 13 11 11 1 11 2
29 16 3 13 0 9 11 11 2 1 9 0 9 13 13 12 9 9 1 0 9 11 7 12 9 1 0 9 11 2
9 11 13 12 0 0 9 0 9 2
21 1 0 9 1 15 13 9 1 9 0 9 2 16 9 1 0 0 9 13 0 2
26 3 13 1 9 9 1 9 12 9 9 2 0 12 9 9 2 15 13 1 9 9 2 13 1 9 2
14 9 11 7 11 13 9 11 9 9 9 1 10 9 2
10 15 0 9 4 13 0 9 0 9 2
16 4 13 7 9 9 9 2 15 13 13 9 12 9 1 9 2
5 0 9 1 0 9
13 1 9 0 9 7 9 13 3 9 3 12 9 9
2 11 11
20 0 9 13 0 9 0 7 0 0 7 0 9 0 0 0 9 1 9 9 2
21 9 13 13 13 0 7 0 9 0 9 7 0 9 2 15 10 9 1 9 13 2
19 9 13 13 3 1 9 1 0 9 2 9 2 9 2 9 2 9 2 2
10 9 9 4 13 9 9 9 1 9 2
18 16 13 9 9 11 11 2 9 13 1 0 9 12 0 9 1 9 2
16 9 1 10 9 2 1 9 1 0 2 13 1 9 10 9 2
40 11 13 2 16 0 9 9 0 9 13 7 3 0 9 1 15 2 16 4 15 0 9 13 13 1 0 9 0 9 2 3 2 9 1 0 9 0 9 2 2
20 1 0 9 4 3 13 0 0 9 9 9 7 9 0 9 0 9 1 9 2
31 9 13 13 9 2 15 13 0 1 9 13 1 9 7 9 0 9 9 2 0 9 2 1 9 0 9 9 7 10 9 2
19 9 1 9 10 9 4 13 7 1 9 9 2 7 1 0 9 0 9 2
32 9 9 4 0 9 13 9 0 0 0 9 2 3 15 13 1 9 7 9 0 1 9 1 9 9 12 1 9 9 12 2 2
10 0 9 9 4 13 12 9 1 9 2
10 9 13 13 1 9 0 16 12 9 2
31 9 9 13 10 9 0 9 1 9 0 9 13 3 1 12 2 9 0 9 2 3 7 1 9 0 2 0 9 9 9 2
30 0 9 4 3 3 13 9 1 9 9 7 9 1 0 9 2 3 0 0 9 9 1 9 0 13 0 16 12 9 2
11 9 9 1 10 9 13 12 9 1 9 2
9 0 9 13 13 0 16 12 9 2
14 9 13 9 2 9 7 9 2 2 15 13 9 9 2
13 9 1 9 15 1 10 9 13 1 12 2 9 2
15 9 9 1 0 9 1 12 0 9 13 9 12 9 9 2
28 13 15 2 16 0 9 4 13 1 11 3 1 12 9 9 7 9 2 3 1 0 11 2 12 9 9 2 2
37 9 0 9 4 1 9 10 9 13 9 0 9 3 7 3 0 9 2 9 0 9 2 9 0 7 3 0 9 7 9 2 9 0 0 9 3 2
14 1 10 9 4 13 14 12 9 9 0 1 0 9 2
9 11 11 13 1 9 13 1 9 11
2 11 2
43 0 9 1 9 2 9 2 9 7 9 0 9 1 9 0 0 9 13 9 9 1 0 9 2 15 1 9 13 0 9 11 11 1 0 9 0 11 9 1 9 1 11 2
21 3 1 9 13 0 9 11 11 11 2 9 9 15 13 0 9 9 9 0 9 2
20 1 0 9 7 9 13 7 1 9 2 1 9 9 7 1 0 7 0 9 2
21 1 0 9 4 13 3 0 0 9 11 11 7 11 0 11 2 9 0 11 2 2
20 1 0 9 13 1 11 12 9 0 9 11 2 11 1 0 0 7 0 9 2
10 1 0 13 3 1 0 9 0 9 2
23 0 9 4 13 3 1 0 9 2 1 11 7 1 0 9 0 9 2 13 0 9 11 2
23 11 13 9 9 0 9 10 7 0 9 1 0 9 7 10 9 13 1 9 9 7 9 2
12 9 11 13 0 9 7 9 0 9 1 11 2
3 0 0 9
2 11 2
29 9 1 9 12 9 9 15 13 9 0 0 9 1 9 9 2 15 4 1 9 13 1 9 1 0 9 1 11 2
18 0 9 15 13 7 0 9 9 9 11 11 7 9 0 9 11 11 2
26 10 9 13 1 0 1 9 7 10 9 4 13 0 9 0 7 0 9 2 13 0 9 9 11 11 2
22 0 9 9 15 13 9 9 12 9 1 9 1 0 0 9 7 0 9 2 13 11 2
37 3 16 12 9 9 9 4 13 1 0 9 2 16 1 0 0 9 13 11 2 9 13 12 12 9 2 2 11 2 11 2 11 2 11 7 11 2
26 1 0 9 13 0 9 0 9 2 0 11 2 11 7 0 2 16 0 9 13 1 12 9 0 9 2
5 11 13 9 1 11
4 11 1 11 2
29 1 0 9 0 9 11 1 9 11 11 1 11 4 1 9 2 15 4 13 3 10 9 2 13 13 9 12 9 2
37 1 9 11 11 11 3 0 9 9 9 11 11 2 15 13 1 9 11 1 9 9 11 0 9 1 11 2 13 0 9 1 9 0 9 1 11 2
30 9 9 1 11 4 1 11 13 13 9 0 9 1 9 0 9 2 7 0 13 7 9 9 9 1 0 9 1 11 2
36 0 9 13 1 15 1 9 13 1 11 1 11 10 9 0 9 1 9 11 7 11 2 16 9 9 7 0 0 7 0 9 13 13 0 9 2
13 11 13 0 9 9 0 0 9 1 11 1 11 2
35 13 3 0 9 7 9 1 9 2 9 1 9 9 2 9 1 0 9 2 0 9 7 0 9 1 9 9 2 9 2 9 2 9 2 2
13 0 9 9 1 9 12 13 9 9 12 9 9 2
15 9 0 9 9 13 7 1 9 12 9 9 13 0 9 2
6 11 11 2 9 1 9
8 0 0 9 7 9 13 9 9
5 11 2 11 2 2
25 16 1 9 12 13 0 9 11 12 9 2 13 3 0 0 9 13 3 12 9 0 7 0 9 2
32 13 4 1 9 9 7 0 0 9 2 13 1 0 0 9 11 11 2 15 13 9 7 0 9 0 9 11 11 1 9 12 2
20 1 9 0 0 9 2 1 0 9 7 1 0 9 13 9 9 0 0 9 2
14 1 9 1 9 9 1 0 9 13 0 2 0 9 2
45 9 0 9 0 12 9 0 1 0 9 1 0 9 13 1 0 9 13 1 0 9 2 3 13 3 12 5 9 2 14 9 7 9 2 7 3 9 0 9 2 9 7 0 9 2
16 9 1 9 0 9 0 9 1 9 0 9 3 13 12 9 2
31 0 0 9 13 7 0 9 2 16 3 0 0 9 2 0 0 0 9 2 9 1 9 7 9 7 0 9 1 0 9 2
9 3 1 0 9 13 0 9 11 2
12 13 1 0 9 15 11 13 3 9 0 9 2
27 1 9 1 0 9 13 9 9 11 11 2 13 15 9 9 1 11 2 3 4 13 9 1 9 9 11 2
10 1 15 9 13 7 3 9 11 0 2
19 0 9 13 13 1 12 5 7 9 9 13 9 0 9 14 1 9 12 2
4 11 0 9 11
2 11 2
20 11 11 1 9 9 13 9 9 0 11 2 1 15 13 9 9 0 0 9 2
17 12 1 9 9 11 11 11 13 2 16 9 13 15 0 9 11 2
14 9 9 13 1 11 2 11 10 9 1 9 0 9 2
18 9 13 1 9 9 7 9 9 1 0 9 7 9 1 0 0 9 2
21 3 9 13 9 12 9 9 11 2 15 9 4 1 9 13 1 0 9 1 11 2
7 0 9 11 13 0 9 2
10 11 13 9 13 0 9 15 9 9 2
16 3 13 1 9 2 3 13 11 2 11 2 3 13 0 9 2
34 1 10 9 13 3 1 9 2 16 13 11 2 11 2 11 7 0 2 1 0 9 2 7 3 1 9 13 10 9 1 0 0 9 2
20 1 0 9 13 3 9 0 2 15 15 13 9 1 9 2 9 7 0 9 2
15 1 11 13 12 9 7 0 9 2 12 9 13 1 11 2
12 9 0 9 4 3 13 13 14 12 9 9 2
15 1 9 9 1 11 4 13 9 13 3 12 7 12 9 2
11 13 4 9 0 9 1 3 12 9 9 2
3 9 1 9
29 9 11 13 12 2 9 1 11 1 9 0 9 2 9 7 9 0 9 0 0 0 9 2 9 7 9 0 9 2
12 9 13 9 0 9 11 1 9 2 9 9 2
21 12 2 9 0 9 13 9 3 0 0 9 2 9 0 9 9 2 9 2 0 2
8 13 1 0 0 0 0 9 2
10 9 15 13 1 11 12 1 11 9 2
21 1 10 9 3 13 1 0 9 11 2 0 2 11 7 11 2 11 2 0 9 2
28 1 0 9 13 0 9 2 9 7 9 2 2 9 9 2 2 0 9 2 0 9 2 7 3 9 7 9 2
9 9 13 13 9 7 9 0 9 2
17 9 13 9 16 9 0 9 2 9 2 2 16 9 7 0 9 2
34 13 2 15 13 2 3 4 15 13 13 0 9 9 0 9 11 2 11 0 11 7 0 0 0 9 1 9 0 0 9 0 9 11 2
21 1 9 9 2 9 7 9 13 1 9 9 14 1 12 0 16 9 0 9 11 2
11 15 3 13 7 3 1 9 1 0 9 2
2 11 2
27 11 13 1 0 9 13 1 9 9 0 9 2 1 15 0 2 0 7 0 2 9 11 13 13 12 5 2
13 15 9 13 13 0 9 7 11 13 9 12 9 2
12 0 9 13 9 1 9 7 9 1 0 11 2
27 11 13 0 9 0 7 0 9 2 1 9 1 0 9 13 9 3 0 0 9 1 9 0 1 9 11 2
9 13 15 15 3 1 12 9 9 2
30 11 15 13 0 9 0 9 1 0 9 0 11 2 15 15 13 1 9 1 9 7 0 9 9 1 9 0 1 9 2
20 9 13 2 16 9 0 1 9 12 9 13 13 7 1 9 1 0 0 9 2
25 11 11 13 1 10 9 0 0 9 2 9 9 1 0 0 9 2 7 2 12 11 2 9 2 2
6 10 9 13 9 11 2
10 9 13 9 12 11 11 2 12 9 2
9 13 13 0 9 1 9 12 9 2
8 1 9 13 7 1 0 9 2
5 0 11 13 0 9
2 11 2
32 0 9 0 11 3 1 11 13 0 9 1 0 9 2 15 4 13 0 0 9 2 15 7 1 10 9 13 0 9 1 11 2
20 1 9 11 11 2 11 4 1 0 12 9 9 13 1 9 3 16 12 9 2
5 11 13 1 0 9
2 11 2
13 1 9 0 0 9 15 3 13 0 9 11 11 2
20 13 3 1 9 0 7 0 9 1 9 9 0 9 11 1 9 11 2 11 2
23 1 11 13 1 9 2 16 15 10 9 7 9 9 13 1 0 9 1 0 9 16 0 2
8 15 7 13 13 9 15 13 2
8 13 15 1 9 13 12 9 2
10 15 0 7 13 13 9 15 13 13 2
28 13 4 15 3 1 0 9 2 15 13 3 13 2 13 9 7 13 2 16 13 7 3 13 13 0 0 9 2
9 0 9 3 13 9 9 3 13 2
5 1 11 15 13 9
8 0 0 9 13 0 9 0 11
7 11 2 11 2 11 2 2
29 12 9 1 0 13 3 1 11 0 0 9 2 15 3 10 9 13 2 3 0 0 7 0 9 0 9 0 11 2
35 9 12 12 0 9 15 3 1 9 13 0 9 2 9 1 15 0 9 1 9 13 15 13 3 2 12 1 0 2 15 3 0 9 13 2
19 0 11 13 9 2 3 0 3 1 0 9 2 1 9 9 10 0 9 2
12 3 0 7 1 0 0 9 13 0 9 9 2
17 1 9 0 9 9 15 1 12 9 9 13 0 9 1 0 9 2
25 0 9 13 3 1 0 9 12 1 0 9 9 2 10 0 9 7 9 13 13 3 9 0 9 2
27 9 0 9 15 1 9 9 2 1 15 0 13 1 0 9 2 3 11 7 11 2 2 13 3 1 0 2
16 16 4 9 3 1 9 13 16 0 2 10 9 13 1 9 2
12 9 1 15 3 13 1 9 1 9 9 9 2
13 1 15 15 13 2 13 13 9 3 1 0 9 2
29 9 13 1 0 9 0 9 0 11 2 3 11 11 2 11 11 7 11 11 2 3 4 3 13 14 1 12 9 2
8 0 11 13 1 11 14 3 2
12 1 10 9 15 0 9 13 3 13 0 9 2
7 0 9 11 1 11 11 13
5 11 2 11 2 2
28 9 0 2 9 2 11 11 13 1 0 0 9 2 16 0 9 11 2 11 13 1 10 9 7 16 9 9 2
22 1 9 9 7 9 9 13 3 11 11 7 11 11 2 15 1 9 1 12 2 9 2
29 9 9 11 11 13 2 16 9 11 13 1 11 13 2 12 9 9 13 2 7 9 2 15 15 13 2 4 13 2
16 9 13 0 2 10 9 4 13 7 3 2 13 7 3 9 2
10 9 11 13 13 1 11 1 9 12 2
22 0 9 0 9 13 9 12 9 12 9 9 2 0 9 4 13 1 9 12 9 9 2
11 11 13 10 9 13 7 13 12 0 9 2
27 0 9 13 3 0 9 1 9 12 2 15 13 0 9 0 0 9 2 0 9 9 7 9 9 1 9 2
11 13 15 7 1 9 9 9 1 10 9 2
21 1 0 9 1 9 7 9 2 11 2 13 11 1 0 9 1 9 12 9 9 2
13 13 13 9 0 9 1 9 7 9 11 1 11 2
6 11 11 13 9 1 11
2 11 2
19 0 9 11 11 3 1 0 11 13 0 9 0 7 0 9 1 0 11 2
21 13 2 16 0 9 13 13 10 0 9 1 0 9 7 0 11 1 9 9 9 2
12 1 0 9 13 10 9 13 3 12 9 9 2
34 0 9 13 3 0 9 1 9 9 1 9 2 16 9 1 0 11 3 13 2 16 1 9 0 9 4 13 9 0 9 7 0 9 2
11 9 9 13 12 1 0 9 9 11 11 2
11 0 9 13 9 0 7 0 9 1 9 2
23 13 2 16 0 9 13 9 0 0 0 0 9 1 0 7 16 4 13 9 11 0 9 2
5 0 9 11 2 11
2 11 2
34 9 9 0 0 9 11 1 0 1 11 2 11 13 1 9 11 11 0 9 0 9 0 9 2 15 13 10 9 1 0 7 0 9 2
28 1 0 9 9 0 9 1 9 13 3 9 2 16 11 13 13 1 9 1 0 9 0 9 7 1 0 9 2
10 9 11 11 11 3 13 0 9 11 2
16 1 9 13 9 9 2 16 9 0 9 1 0 9 13 0 2
27 13 15 15 1 9 2 3 0 9 13 12 9 9 7 0 9 12 9 2 13 13 9 9 2 13 11 2
10 9 11 13 9 3 3 0 9 6 11
2 9 11
6 0 9 13 1 9 9
5 11 2 11 2 2
13 3 0 9 11 11 15 13 13 1 9 0 9 2
37 1 9 15 3 13 0 9 0 0 9 11 2 0 1 11 2 11 2 11 7 11 2 2 0 2 9 2 11 7 9 2 9 2 0 2 11 2
30 11 11 13 3 9 12 0 9 2 3 2 11 2 11 7 0 2 7 9 2 15 13 1 9 0 0 2 0 9 2
14 13 15 9 11 2 11 2 15 9 0 9 13 11 2
18 1 15 1 10 9 13 11 11 1 11 7 11 13 9 12 9 9 2
21 9 11 11 13 0 9 9 2 16 4 0 9 16 0 9 13 1 9 0 9 2
27 1 9 2 16 9 1 10 0 9 3 13 1 15 2 15 13 13 7 3 13 2 11 13 2 16 14 2
12 10 9 7 13 3 2 16 1 9 13 11 2
13 13 13 2 16 11 13 9 10 9 2 13 11 2
32 1 9 11 1 9 9 13 2 16 13 0 9 1 11 2 3 3 13 0 9 9 1 11 7 1 0 9 13 7 1 11 2
11 9 13 1 9 9 9 13 12 2 9 2
34 13 4 15 13 2 16 16 9 0 9 3 13 1 10 9 9 2 10 9 2 13 2 3 15 1 9 13 2 2 14 15 15 13 2
36 16 3 9 0 7 3 0 0 9 13 7 3 0 2 9 9 3 13 0 9 14 1 15 2 16 4 15 13 2 15 15 3 13 1 9 2
22 7 3 4 1 0 9 13 9 1 9 1 9 13 3 2 16 15 10 9 13 13 2
35 10 9 9 13 3 0 2 7 15 7 1 9 1 0 9 9 11 2 2 7 1 0 9 13 0 0 9 0 9 1 9 9 1 9 2
21 7 16 15 3 13 9 2 13 3 1 15 2 3 13 0 7 0 9 10 9 2
28 1 15 1 0 9 3 13 10 9 1 9 2 9 2 10 9 13 0 9 12 3 2 7 3 3 0 9 2
3 2 11 2
3 0 0 9
2 11 11
17 3 4 13 2 3 15 13 2 1 9 0 15 13 9 1 11 2
13 15 15 13 1 15 2 1 15 13 13 14 9 2
11 15 3 13 2 15 7 10 9 15 13 2
7 13 15 3 10 0 9 2
11 13 2 16 4 15 15 13 9 0 9 2
12 13 1 0 9 2 15 3 13 2 13 0 2
29 13 15 3 3 2 16 1 9 0 11 3 9 9 13 1 15 2 16 15 13 3 3 16 1 11 7 3 3 2
12 9 0 9 13 14 1 0 9 9 9 0 2
17 14 3 2 16 4 10 9 0 9 13 13 9 0 9 1 11 2
13 3 4 13 0 0 9 13 0 9 2 3 13 2
17 16 2 7 15 13 0 9 2 2 16 1 15 13 0 0 9 2
44 3 13 9 2 16 10 9 1 11 13 2 7 16 13 2 13 1 15 2 16 4 15 15 1 15 13 2 7 16 4 15 3 1 15 15 13 2 1 10 9 4 15 13 2
12 15 4 15 0 0 9 13 1 0 9 13 2
15 9 0 7 0 2 16 0 9 15 1 0 9 3 13 2
31 0 9 7 9 1 15 2 16 1 9 13 9 9 0 1 9 0 2 13 0 0 9 14 16 9 9 11 1 9 0 2
10 1 9 1 11 13 9 3 0 9 2
12 3 16 3 7 16 3 3 13 13 9 0 2
34 16 13 9 9 11 1 0 9 0 9 1 0 9 3 9 1 0 9 2 3 13 0 9 11 11 2 7 16 13 15 0 0 9 2
13 16 13 0 13 0 0 9 0 9 1 0 9 2
32 7 3 13 9 3 12 9 2 3 13 9 2 16 0 9 3 13 2 7 3 13 9 1 9 9 1 9 1 9 7 3 2
18 1 9 11 11 1 3 0 2 3 0 11 0 9 1 15 15 13 2
7 0 0 9 15 3 13 2
9 7 13 0 9 3 1 10 9 2
11 16 3 10 9 4 13 1 11 13 9 2
4 0 9 1 11
2 11 2
22 0 9 7 0 9 13 0 0 9 2 16 4 13 9 9 1 9 9 7 0 9 2
12 11 15 3 13 9 0 9 1 11 11 11 2
21 12 1 9 1 9 10 9 13 0 9 2 1 15 9 9 13 7 3 15 13 2
30 3 0 13 9 2 15 0 9 1 11 13 1 9 1 9 11 2 11 1 9 7 9 10 0 9 0 9 1 9 2
18 1 9 0 9 13 2 16 13 9 1 9 7 13 9 9 11 11 2
25 1 1 15 2 16 10 9 13 13 2 0 0 9 3 13 0 9 7 13 0 9 1 0 9 2
24 1 9 1 0 9 10 9 1 9 1 0 9 13 1 9 7 9 0 9 0 9 7 9 2
16 0 9 4 13 9 2 15 13 13 1 0 9 1 0 9 2
20 0 9 15 13 3 15 2 16 9 0 9 3 1 9 13 13 7 0 9 2
4 9 13 0 9
2 11 2
29 9 0 9 13 1 9 12 9 9 2 9 0 9 13 12 9 9 7 3 9 13 13 12 9 9 1 0 9 2
13 13 15 1 9 9 2 15 1 9 13 9 11 2
7 9 11 11 2 11 1 9
2 11 2
21 9 0 11 11 11 4 1 9 11 13 7 9 15 1 9 0 9 13 1 9 2
10 9 3 11 13 1 9 9 10 9 2
19 11 13 4 3 13 1 9 1 11 2 16 13 13 1 9 10 9 11 2
27 1 9 1 10 9 4 13 7 10 0 9 7 13 13 2 16 13 1 15 7 9 11 11 2 13 11 2
17 0 9 4 13 1 0 9 3 1 9 1 0 9 1 9 11 2
5 11 13 0 0 2
16 12 0 9 2 15 15 15 1 9 3 13 2 9 3 13 2
5 0 9 13 7 9
5 11 2 11 2 2
27 9 1 9 1 11 2 1 9 9 7 0 9 2 0 9 7 0 9 13 9 1 9 3 12 0 9 2
14 1 9 0 9 9 15 13 9 9 0 9 11 11 2
21 0 9 15 13 3 1 0 0 7 0 9 7 3 15 13 1 0 9 0 9 2
19 13 13 1 0 9 0 9 2 7 7 1 11 2 11 2 11 7 11 2
18 1 11 4 13 9 13 1 9 9 2 3 16 1 0 11 7 11 2
12 1 0 9 13 11 2 3 11 7 0 11 2
23 1 12 2 9 9 13 9 0 9 2 15 13 1 9 0 9 7 3 13 1 0 9 2
13 9 9 13 1 9 0 9 7 9 9 1 9 2
14 1 9 0 9 1 9 4 15 13 3 13 0 9 2
19 11 13 2 16 4 9 13 0 9 13 9 1 9 0 9 1 0 9 2
10 1 12 9 15 1 15 13 0 9 2
13 1 0 9 7 13 1 9 12 9 9 1 9 2
6 1 15 13 9 9 2
17 16 7 13 9 11 11 2 1 9 10 9 1 12 9 13 9 2
6 11 13 9 1 9 3
5 11 2 11 2 2
19 16 9 9 0 9 1 0 12 9 3 13 2 9 9 1 11 3 13 2
15 16 1 9 12 13 12 9 9 2 3 15 13 14 12 2
21 9 11 11 15 3 3 13 1 10 9 2 16 3 0 9 0 0 9 13 0 2
7 1 9 13 11 12 9 2
21 0 13 1 9 13 9 0 9 2 15 0 9 13 0 9 2 1 0 9 13 2
21 12 0 9 0 1 9 9 13 7 9 13 9 7 1 9 11 2 3 1 11 2
20 9 13 1 11 2 3 13 1 10 0 9 2 0 9 13 3 1 12 9 2
15 1 9 12 15 13 9 9 13 7 1 9 9 0 9 2
10 1 12 0 9 13 13 3 12 0 2
36 9 13 9 1 9 0 9 2 3 15 1 15 0 13 3 1 9 2 13 0 2 0 9 2 15 3 13 13 0 9 0 9 1 0 9 2
8 9 7 13 1 9 0 9 2
9 3 3 13 1 0 0 9 9 2
35 9 0 9 9 7 9 11 11 13 2 16 16 15 9 13 2 13 0 9 10 0 9 2 7 1 9 9 0 9 13 9 10 9 0 2
11 1 15 9 9 13 3 3 16 9 9 2
10 13 15 3 3 3 13 3 1 9 2
3 9 16 3
2 11 2
26 1 9 4 13 11 7 9 11 9 13 15 9 2 3 4 14 13 0 9 2 16 4 13 9 0 2
18 3 15 3 13 13 0 9 2 15 4 13 9 1 9 1 9 12 2
5 12 9 1 0 9
5 11 2 11 2 2
20 0 9 11 13 1 12 2 9 10 9 1 0 9 9 9 9 1 0 9 2
21 1 9 15 1 11 13 13 0 12 9 9 7 9 2 9 11 11 7 9 11 2
7 9 11 15 7 9 13 2
15 13 1 12 9 0 9 2 3 9 2 9 2 9 0 2
15 0 9 13 3 9 9 2 9 9 9 12 9 1 11 2
11 9 13 0 9 1 12 7 1 12 9 2
7 9 1 12 1 12 9 2
5 13 2 7 13 2
2 11 11
16 0 9 13 3 1 10 9 2 0 9 2 14 3 15 0 2
37 13 14 9 2 16 9 9 15 3 16 0 9 13 2 7 13 3 9 2 16 13 14 9 9 2 3 15 9 1 0 9 0 9 0 9 13 2
18 1 10 9 7 9 0 0 9 15 3 3 13 9 9 0 9 9 2
16 13 15 9 2 15 4 3 3 3 13 2 13 2 7 13 2
15 13 15 13 2 16 0 9 0 9 9 13 3 1 9 2
18 0 9 3 13 1 9 1 0 9 3 3 9 2 9 7 9 9 2
12 15 3 13 15 0 2 15 9 1 9 13 2
7 9 15 13 7 3 3 2
34 1 0 9 9 2 9 9 7 9 1 9 2 9 9 7 9 3 2 13 3 0 9 1 15 9 2 9 7 0 9 1 0 9 2
31 3 1 9 9 1 3 0 9 15 14 13 9 2 7 3 13 15 0 9 2 9 2 9 2 9 9 13 3 2 2 2
47 9 13 1 9 9 9 1 9 9 2 9 1 9 2 9 2 9 7 9 2 15 15 13 0 9 9 9 2 7 2 9 0 7 0 9 2 9 9 2 9 2 9 7 9 9 3 2
18 1 15 9 13 1 9 9 9 0 0 9 2 3 1 9 15 9 2
24 13 7 3 13 0 9 7 9 0 9 9 1 9 7 11 1 2 2 2 2 1 9 2 2
18 9 9 0 9 13 2 16 15 1 15 2 15 13 2 13 13 3 2
24 13 3 0 13 15 9 2 16 13 3 9 2 15 13 13 2 2 3 13 13 3 1 9 2
11 13 15 9 2 9 2 9 1 10 9 2
21 13 15 3 1 9 1 9 0 2 16 15 3 13 2 13 15 1 0 9 3 2
21 3 9 2 1 15 15 13 1 10 9 2 13 2 14 2 1 15 3 3 0 2
20 13 4 3 12 9 2 13 1 11 2 13 9 13 1 9 7 3 15 13 2
17 13 3 9 3 2 16 13 9 9 7 13 2 16 13 7 13 2
15 0 13 3 0 9 14 3 2 16 13 13 0 0 9 2
23 10 3 0 9 13 1 9 13 10 9 0 9 2 15 4 13 1 9 2 0 9 9 2
39 1 0 0 9 13 9 2 9 1 10 9 0 9 2 15 13 9 9 1 9 15 0 2 7 9 2 9 1 9 0 9 2 3 0 9 1 0 9 2
22 3 13 2 3 4 12 0 9 13 7 13 3 2 16 1 0 9 15 3 3 13 2
24 9 2 13 9 9 2 13 0 9 1 9 1 3 0 9 7 16 9 13 2 13 1 15 2
29 16 13 9 2 13 1 0 2 0 7 0 9 9 2 1 0 9 0 9 0 9 2 1 9 9 1 9 3 2
12 3 13 9 16 9 2 7 3 14 1 9 2
18 9 3 13 14 9 2 7 7 9 9 0 2 0 2 0 7 0 2
18 1 9 4 3 10 9 0 9 2 15 13 13 9 9 2 13 9 2
43 1 0 9 13 9 7 13 9 2 0 9 2 13 1 0 9 10 9 2 1 0 9 2 9 10 9 7 0 9 2 0 9 2 3 2 10 9 1 0 9 2 3 2
8 15 0 3 3 3 1 9 2
26 9 13 3 1 12 9 2 7 1 0 2 3 9 9 13 7 13 9 7 15 2 7 1 9 9 2
15 16 13 9 1 9 2 13 15 13 1 0 2 0 9 2
13 9 3 13 1 9 16 0 9 2 7 7 0 2
13 1 0 9 15 9 13 3 13 1 15 10 9 2
11 16 9 13 0 9 2 13 15 3 3 2
17 9 0 9 4 13 13 9 2 1 15 15 13 10 9 0 9 2
15 13 2 14 9 1 0 9 2 3 10 9 13 16 9 2
24 1 9 4 13 13 16 2 13 2 14 1 9 2 7 9 2 13 2 14 1 3 0 9 2
6 13 0 9 13 0 2
8 0 9 13 9 0 16 9 2
20 1 9 13 9 13 9 1 9 9 7 13 2 16 13 13 16 9 1 13 2
37 16 15 1 15 0 9 13 2 10 9 9 13 7 3 15 13 1 15 2 16 15 9 13 1 15 2 16 1 13 13 1 9 3 2 13 9 2
52 13 15 13 0 15 2 16 16 0 9 2 0 9 2 0 9 3 2 3 13 13 2 16 13 1 15 2 16 4 15 0 9 13 2 0 9 1 0 9 4 13 13 3 16 10 2 3 14 0 2 9 2
20 14 15 2 15 13 2 13 3 7 3 2 14 15 2 15 13 2 13 3 2
26 3 4 13 0 2 16 4 15 9 3 13 9 0 9 0 9 13 0 1 0 9 0 9 13 0 2
11 14 1 9 0 1 15 3 15 13 13 2
12 16 13 9 3 0 9 2 0 9 15 13 2
20 9 15 13 9 13 2 3 15 9 13 13 3 2 16 13 13 3 0 9 2
15 13 9 9 2 15 13 0 2 7 1 0 9 15 13 2
11 13 1 15 9 9 2 9 2 9 3 2
14 15 15 13 3 9 1 15 2 10 9 13 7 13 2
14 13 1 15 9 9 3 1 9 7 3 7 1 15 2
44 1 9 9 16 0 9 9 13 7 1 2 0 2 9 13 1 15 2 16 13 1 9 9 2 15 10 0 2 3 0 7 3 0 0 9 13 1 9 0 0 9 1 9 2
15 1 9 1 0 9 9 13 0 9 0 9 1 9 9 2
20 16 1 10 9 4 3 13 2 13 4 13 1 0 9 1 9 7 0 9 2
4 9 13 1 9
8 0 9 0 9 7 1 9 13
7 11 2 11 2 11 2 2
34 0 9 3 0 9 4 13 13 1 0 9 9 9 9 1 9 1 9 2 9 7 0 9 0 9 0 9 0 1 9 1 0 9 2
27 0 9 1 0 9 7 9 2 15 3 1 9 9 13 9 2 7 9 0 15 0 9 3 0 9 13 2
11 9 13 1 10 9 9 0 7 0 9 2
28 1 9 4 13 4 13 13 7 13 0 9 9 0 12 9 7 13 4 4 13 7 9 0 9 1 0 9 2
11 0 9 13 9 0 9 9 0 12 9 2
29 9 3 13 2 16 4 4 13 13 3 1 0 9 2 9 7 9 0 1 0 9 2 1 9 9 0 1 9 2
19 9 13 2 16 4 9 0 9 3 13 0 9 1 9 3 12 9 9 2
18 1 9 4 13 0 13 9 2 9 7 9 0 9 1 9 0 9 2
26 1 9 0 9 0 7 0 1 0 9 4 13 9 0 13 0 9 1 9 9 2 9 7 9 0 2
26 9 9 13 0 7 9 9 9 0 9 11 11 2 15 13 2 16 0 13 3 9 9 2 7 9 2
12 1 9 9 13 1 10 9 0 9 3 13 2
9 1 10 9 3 0 0 9 13 2
6 9 9 9 1 0 9
2 11 2
16 9 9 0 0 9 13 9 0 9 2 0 0 9 9 9 2
11 9 13 1 9 11 7 1 9 1 15 2
7 9 4 13 3 1 11 2
51 3 13 1 11 2 3 1 11 2 12 2 12 2 2 2 0 11 2 12 2 12 2 2 2 11 2 12 2 12 2 2 2 11 2 12 2 12 2 2 7 1 9 1 11 2 12 2 12 2 2 2
2 9 13
2 11 2
8 0 9 1 9 0 3 13 2
7 13 7 13 7 9 0 2
10 13 15 11 2 11 1 0 0 9 2
11 1 9 11 7 11 15 3 13 9 0 2
15 3 1 11 7 1 0 0 9 4 3 9 10 9 13 2
14 3 0 13 0 9 2 15 13 3 0 3 1 9 2
1 3
10 0 9 13 1 9 0 9 11 9 2
22 0 9 15 1 9 13 2 16 15 3 13 1 9 1 0 0 9 1 9 0 9 2
18 13 2 16 13 3 1 0 9 2 13 1 15 9 9 11 11 11 2
32 3 12 9 2 9 2 9 7 9 12 3 0 9 1 11 13 0 9 1 9 9 9 2 15 4 3 13 1 0 0 9 2
7 9 13 1 12 2 9 2
6 15 13 1 9 11 2
3 1 0 9
4 11 2 11 2
27 0 9 9 3 1 10 9 13 11 11 2 16 4 13 9 2 15 7 3 15 1 15 13 1 9 11 2
17 9 13 1 11 1 9 1 11 13 1 0 9 0 1 9 11 2
21 13 9 9 2 16 4 13 10 0 9 7 15 2 10 9 15 1 9 11 13 2
7 3 4 15 13 9 13 2
24 1 0 9 15 15 13 7 15 4 15 13 13 1 9 0 9 0 9 2 13 15 1 9 2
7 9 1 9 13 9 1 9
5 11 2 11 2 2
26 9 1 15 9 9 13 3 1 9 10 9 13 0 9 1 9 2 15 9 1 10 0 9 13 9 2
22 16 1 10 9 13 9 9 11 11 2 1 0 9 4 1 9 13 13 7 0 9 2
32 9 13 12 9 0 9 2 9 1 9 2 7 2 9 7 9 9 2 2 9 0 9 7 9 9 2 15 13 9 7 9 2
35 1 0 9 9 7 9 1 11 13 9 0 9 7 13 13 10 0 9 2 1 15 4 15 13 14 12 9 13 7 9 13 1 10 9 2
14 0 9 4 15 1 9 9 13 13 1 0 9 9 2
13 9 4 1 11 13 4 13 9 0 2 3 0 2
13 1 0 9 4 10 9 13 9 1 9 1 9 2
25 9 3 3 13 9 1 0 9 0 0 9 2 15 13 0 9 2 15 9 13 9 15 0 9 2
49 9 3 13 9 1 9 12 2 0 9 9 0 9 9 11 0 1 9 0 0 9 2 15 15 4 13 9 9 1 11 2 7 13 9 9 9 1 9 2 15 9 13 9 11 11 2 11 2 2
15 11 4 3 13 0 9 1 10 9 1 9 1 0 9 2
25 13 15 3 1 11 9 0 0 9 2 0 9 9 2 11 11 1 9 1 9 0 9 11 11 2
19 11 7 11 15 13 9 1 9 1 11 7 11 1 9 10 9 1 11 2
12 13 3 1 0 9 0 1 9 1 10 9 2
5 9 11 11 2 11
8 11 2 11 13 1 9 9 11
5 11 2 11 2 2
21 9 9 1 0 9 13 0 2 7 1 9 4 13 0 9 2 15 4 15 13 2
15 11 15 13 9 0 9 1 0 9 11 11 2 11 2 2
22 10 9 13 1 9 2 16 11 10 0 9 0 1 9 9 3 13 9 9 0 9 2
20 1 11 13 10 9 13 0 9 2 7 9 1 0 9 13 2 7 15 13 2
22 1 0 9 13 2 16 4 14 13 4 13 0 0 9 7 9 9 1 9 0 9 2
17 0 9 2 0 3 2 7 1 11 2 3 13 0 9 0 9 2
16 11 13 1 9 9 11 11 2 1 15 4 11 9 13 13 2
29 11 13 3 9 1 9 14 3 2 16 15 13 3 1 9 10 0 9 2 15 13 0 9 16 9 11 2 13 2
1 9
16 9 2 9 2 14 13 2 16 1 0 9 13 9 13 3 2
14 0 9 13 1 9 13 14 9 2 7 10 0 9 2
8 3 15 13 9 9 2 9 2
25 9 9 13 12 9 2 0 9 7 0 9 2 7 12 9 2 9 0 9 7 3 0 0 9 2
7 15 15 13 1 0 9 2
8 1 9 15 13 0 9 9 2
19 0 9 15 9 13 7 16 0 9 1 0 9 7 3 1 9 0 9 2
22 9 2 0 9 15 3 13 7 13 2 16 9 1 9 13 9 1 9 10 0 9 2
26 16 4 15 15 13 2 9 15 13 2 16 3 13 3 0 11 12 2 7 3 13 1 9 12 2 2
31 13 9 2 16 9 0 9 13 1 9 0 9 3 3 13 2 3 15 13 7 3 2 2 3 10 0 9 15 13 9 2
5 9 11 1 9 9
5 11 2 11 2 2
35 9 9 11 2 11 2 11 2 1 9 9 0 9 9 9 0 9 9 1 9 12 2 15 9 13 0 9 11 2 4 13 13 9 9 2
11 11 15 3 13 9 0 9 11 11 11 2
22 10 9 4 13 4 10 9 13 2 7 15 13 9 9 9 13 2 7 14 2 13 2
32 16 9 11 13 9 9 1 9 9 9 7 4 1 15 13 2 14 3 13 2 3 7 13 2 16 9 9 0 9 9 13 2
8 11 13 9 11 13 1 9 0
6 0 11 2 11 2 2
23 0 0 0 9 11 11 15 13 0 9 0 11 1 0 9 7 3 13 1 9 0 11 2
18 9 0 9 4 13 2 16 13 15 3 0 2 13 11 11 2 11 2
18 1 0 9 3 3 13 1 0 0 9 2 15 1 15 13 0 9 2
26 13 4 0 0 9 1 9 7 1 9 7 1 0 9 4 3 3 13 1 0 9 9 2 13 11 2
15 16 0 9 10 9 1 0 9 13 9 13 1 9 0 2
10 11 2 11 13 1 9 11 16 0 2
12 1 10 9 15 1 15 13 3 9 1 9 2
27 16 4 13 2 16 10 9 13 3 1 10 9 2 13 0 9 2 13 9 9 2 13 1 9 1 11 2
21 0 9 0 9 13 11 1 0 9 2 3 1 0 9 2 1 15 13 9 9 2
5 0 0 9 15 13
5 11 2 11 2 2
12 9 9 1 0 9 3 9 13 13 0 9 2
27 1 9 9 11 11 2 11 2 13 9 9 9 0 0 9 1 12 2 9 12 2 16 0 9 3 13 2
17 11 3 13 2 16 0 9 9 13 4 13 1 9 1 0 9 2
28 9 9 3 13 9 9 1 0 9 2 7 13 9 9 11 11 2 11 2 13 9 1 0 9 9 7 9 2
23 16 3 4 9 9 1 9 0 9 13 3 2 1 9 4 15 13 1 11 13 3 9 2
29 1 11 11 2 11 2 4 15 7 13 4 13 9 2 1 10 9 13 10 0 9 7 15 13 1 0 9 13 2
15 9 1 9 13 3 2 9 2 9 2 0 9 7 0 9
5 11 2 11 2 2
15 3 9 0 9 13 1 9 0 0 9 9 9 0 9 2
24 3 3 1 9 15 9 13 1 0 9 2 3 13 13 12 9 9 1 9 7 9 1 9 2
41 9 9 11 11 11 3 11 13 2 16 1 0 9 0 9 3 1 9 13 9 1 0 9 2 1 9 1 9 2 1 9 7 9 0 0 9 7 9 0 9 2
26 3 1 0 0 9 9 1 0 0 9 4 9 13 13 12 9 9 0 0 9 0 9 9 2 9 2
50 13 1 9 9 0 9 2 15 1 9 13 1 9 0 0 9 2 9 11 11 2 11 2 11 2 2 15 9 4 3 3 3 13 2 7 9 0 9 1 9 9 2 15 13 11 11 2 11 2 2
21 7 1 9 9 10 1 0 12 9 4 15 3 0 9 1 9 13 13 3 3 2
30 9 15 1 9 9 11 11 11 13 13 1 9 0 9 7 9 11 11 2 11 2 13 0 9 11 3 1 9 9 2
17 9 4 15 13 1 9 13 7 0 9 0 9 1 9 0 9 2
50 7 1 1 15 2 16 9 9 9 11 11 2 11 2 1 10 9 3 13 9 0 9 7 1 12 2 9 13 9 9 13 1 10 9 0 9 2 9 9 2 3 1 11 2 13 1 0 9 0 2
19 1 9 9 7 9 4 13 9 13 9 9 1 0 9 11 1 9 12 2
42 1 0 9 9 13 1 9 9 9 3 2 13 9 9 1 9 1 9 0 9 2 1 0 9 2 1 0 2 0 2 0 7 0 9 7 1 9 9 7 0 9 2
18 1 9 0 9 11 4 9 9 13 13 9 0 9 1 0 0 9 2
23 16 0 9 9 13 0 2 0 9 9 13 14 3 13 2 7 13 1 0 9 9 9 2
13 9 1 11 11 2 11 2 2 9 0 9 9 2
21 9 9 9 11 11 13 9 2 16 0 9 13 9 1 9 0 7 0 0 9 2
12 13 7 13 9 1 9 0 9 3 1 9 2
8 13 9 1 9 3 3 0 2
21 13 4 15 9 11 13 2 13 0 9 9 7 13 0 2 16 15 9 3 13 2
12 13 7 9 2 16 0 9 13 9 1 9 2
23 13 15 0 9 2 1 10 9 13 9 13 10 0 9 7 13 15 0 0 7 0 9 2
12 9 4 13 1 0 9 13 9 11 16 9 2
20 7 15 13 13 0 1 0 9 0 9 2 16 13 15 9 2 9 7 9 2
9 1 9 10 9 13 7 9 9 2
16 7 7 15 13 9 2 15 13 13 3 1 9 0 0 9 2
20 13 2 16 10 0 9 13 0 2 7 13 13 1 9 7 0 9 0 9 2
18 3 2 16 1 9 1 9 0 9 4 13 2 16 13 0 15 13 2
8 13 7 13 9 1 0 9 2
3 2 11 2
5 11 1 9 3 3
3 1 0 9
10 11 2 11 11 2 11 2 11 2 2
25 1 0 9 1 0 9 1 0 11 13 11 3 1 11 2 11 2 11 1 11 2 11 7 11 2
19 3 1 11 13 11 9 1 11 7 9 0 7 1 0 11 1 0 9 2
11 13 15 3 9 0 0 9 11 11 11 2
16 1 11 13 11 0 9 1 0 9 7 1 12 0 0 9 2
15 1 0 9 11 13 9 1 11 2 11 2 11 7 11 2
25 1 11 13 0 9 12 0 9 1 0 11 9 1 11 7 13 9 0 0 9 1 9 0 9 2
15 1 12 9 7 9 0 11 13 11 0 9 1 0 9 2
13 1 0 12 9 4 13 3 1 9 1 0 9 2
18 1 0 0 9 0 0 9 11 1 11 11 15 13 10 9 11 11 2
6 11 13 13 2 7 13
3 1 0 9
5 11 2 11 2 2
28 11 11 2 0 9 9 1 9 9 7 9 3 0 1 11 2 4 13 1 0 9 2 11 2 1 0 9 2
28 1 0 9 9 11 13 9 0 9 0 11 11 11 2 3 15 3 13 7 0 9 11 11 11 7 11 11 2
20 16 3 13 11 2 11 2 9 0 9 1 10 0 9 13 13 2 7 13 2
11 11 13 13 9 11 16 0 9 3 11 2
1 9
10 3 1 9 12 15 3 13 0 9 2
26 9 13 1 0 9 1 0 0 9 1 12 5 2 9 15 13 1 12 5 2 16 3 13 12 5 2
15 9 13 9 0 9 0 9 1 0 9 0 7 0 9 2
2 9 11
8 0 9 2 1 9 1 0 11
7 1 9 0 9 2 12 2
2 11 11
14 9 1 9 13 1 11 3 13 1 9 12 2 9 2
24 9 15 13 9 1 12 9 2 9 3 0 7 0 2 16 4 15 15 13 13 7 13 9 2
10 0 9 13 9 0 9 2 9 2 2
26 0 9 11 13 16 0 9 9 12 9 1 9 2 0 1 9 0 2 9 2 3 0 0 9 9 2
6 13 15 3 9 12 2
29 0 9 11 13 3 3 9 2 15 15 1 3 0 9 0 7 0 9 13 1 9 12 13 0 11 2 0 9 2
23 9 12 15 1 11 13 12 9 1 0 9 2 0 11 11 7 1 12 9 0 11 11 2
17 12 13 0 9 1 9 7 9 13 9 10 9 2 0 0 9 2
15 13 1 9 12 9 2 11 13 0 9 7 11 0 9 2
8 0 9 13 1 9 0 9 2
18 9 11 0 2 15 15 1 15 3 3 13 13 2 15 3 13 9 2
19 12 9 15 15 13 15 2 16 1 15 13 10 0 9 1 9 0 9 2
10 13 1 15 0 12 9 9 11 12 2
23 2 9 11 2 9 2 13 11 2 15 15 3 13 1 11 7 3 13 1 9 9 9 2
19 9 13 9 9 7 1 15 2 3 13 11 2 15 15 0 3 13 2 2
9 9 0 11 3 13 1 0 9 2
21 7 1 0 11 2 3 1 10 9 13 9 3 9 2 13 10 9 9 3 0 2
25 9 11 12 2 15 13 1 9 9 12 2 13 1 0 9 15 2 15 11 9 9 1 9 0 2
8 13 11 7 3 13 1 11 2
13 0 3 0 9 13 3 9 9 1 9 0 9 2
10 9 0 9 7 4 13 3 0 9 2
18 11 9 12 13 0 0 9 2 9 12 7 2 1 9 3 2 12 2
30 10 0 9 1 12 9 7 3 0 0 9 9 0 9 1 9 0 15 13 0 9 1 0 0 9 3 2 1 11 2
18 9 12 13 9 10 0 0 9 2 0 3 11 11 2 0 9 2 2
5 3 13 9 9 2
22 11 15 1 15 9 13 1 0 9 2 15 13 16 9 11 11 2 7 9 10 9 2
21 9 1 9 15 13 13 3 0 16 9 3 2 3 15 9 10 9 13 1 11 2
27 11 11 13 0 9 2 7 3 1 15 13 0 9 11 2 11 2 12 2 7 11 2 11 2 12 2 2
14 11 11 2 11 4 13 1 0 9 11 2 9 12 2
9 3 1 9 15 3 13 0 9 2
23 1 0 9 2 1 15 0 9 13 0 0 9 2 11 3 3 13 9 0 9 9 11 2
14 1 15 13 0 9 13 1 9 1 0 2 0 9 2
6 0 13 15 16 0 2
17 9 0 1 11 15 13 13 3 7 1 15 9 3 16 0 9 2
26 3 13 1 15 13 2 16 15 9 2 15 13 13 1 11 11 2 13 3 13 7 1 11 0 9 2
23 0 9 3 2 15 13 9 0 9 2 13 9 11 2 9 13 1 9 9 7 9 2 2
18 9 9 15 7 13 13 3 0 2 16 3 15 9 11 13 1 9 2
25 9 9 11 13 1 3 0 9 7 9 0 11 2 0 0 9 2 15 13 7 13 1 0 9 2
31 1 9 12 2 13 2 14 13 9 2 15 9 9 0 9 11 7 11 13 14 1 12 5 1 11 7 12 5 1 11 2
19 11 13 3 3 3 0 0 9 0 9 2 0 11 3 0 10 0 9 2
4 0 9 0 9
5 11 2 11 2 2
24 1 0 9 0 9 4 13 0 11 11 11 2 2 7 1 9 11 3 13 10 0 9 11 2
7 9 9 13 1 9 11 2
22 1 9 9 9 13 11 11 2 9 9 9 14 1 12 9 2 9 9 7 0 9 2
6 0 9 13 1 9 9
2 11 2
42 9 1 0 9 0 9 9 1 0 11 0 9 2 11 11 2 1 0 9 0 9 9 2 9 0 9 7 0 9 0 9 13 3 0 0 9 1 0 9 1 11 2
25 0 9 0 9 9 2 11 11 2 13 1 9 0 9 1 0 9 13 9 14 12 9 1 11 2
21 13 3 13 2 16 0 9 2 15 1 0 11 13 1 9 2 13 13 7 3 2
20 9 13 9 2 11 11 2 13 1 0 9 2 1 9 7 9 9 0 9 2
10 9 4 13 9 12 2 9 0 9 2
16 1 9 13 13 1 15 0 7 0 9 1 9 1 12 9 2
5 9 9 13 1 9
5 11 2 11 2 2
41 0 0 9 11 2 11 2 1 11 2 15 1 9 1 9 11 1 0 9 1 9 10 9 13 12 9 1 3 0 9 10 9 2 13 0 9 3 1 0 9 2
11 13 13 1 0 9 9 7 9 0 9 2
5 9 13 1 9 2
7 9 10 9 13 0 9 2
13 9 13 1 9 7 9 2 16 4 13 3 13 2
21 3 9 13 7 13 2 13 1 9 11 9 0 9 9 11 9 2 11 2 11 2
4 1 9 9 13
5 11 2 11 2 2
12 3 13 9 0 9 1 0 9 0 11 11 2
14 9 0 1 9 13 0 9 7 3 3 0 0 9 2
19 1 9 15 13 0 9 2 15 1 11 11 2 13 0 9 0 1 9 2
28 11 11 2 13 13 1 0 9 9 1 0 9 2 9 1 9 9 7 9 7 0 9 1 9 1 0 9 2
25 9 10 9 3 13 1 0 9 1 9 9 2 15 0 13 1 12 9 7 15 4 13 16 0 2
8 9 13 2 16 9 13 1 9
2 0 9
5 11 2 11 2 2
32 9 0 9 13 1 9 1 0 9 9 1 9 9 2 11 11 2 2 15 13 16 0 9 13 1 9 3 16 12 9 9 2
12 10 9 15 13 1 11 13 0 9 0 9 2
22 9 9 2 11 2 11 3 16 10 9 7 13 2 16 0 9 0 0 9 4 13 2
17 9 2 11 11 2 13 1 9 2 15 15 13 1 0 9 11 2
21 9 7 1 15 13 1 9 9 2 1 15 13 9 3 13 2 3 1 0 9 2
10 9 13 1 0 9 13 12 0 9 2
4 13 15 3 2
12 1 0 9 1 11 3 13 0 9 0 9 2
20 12 1 9 9 13 2 16 13 9 1 9 7 9 9 2 3 1 9 9 2
14 9 13 9 1 0 9 1 0 7 0 9 15 13 2
21 1 9 0 13 0 9 7 9 1 0 9 1 0 9 2 15 1 9 12 13 2
15 13 15 1 9 2 3 3 9 2 11 11 2 9 13 2
14 1 9 2 11 2 11 1 9 10 9 13 0 9 2
8 15 4 13 9 1 9 13 2
8 7 9 4 9 0 9 13 2
9 9 4 13 0 9 13 10 9 2
6 1 12 9 12 9 9
1 9
2 11 11
34 9 2 15 15 3 3 13 1 3 0 9 2 16 1 15 0 13 9 2 16 1 11 13 12 9 2 4 13 1 12 9 9 9 2
15 9 13 1 10 9 1 0 9 1 11 7 13 3 0 2
8 13 15 9 0 2 7 0 2
20 1 9 9 13 11 2 11 2 0 9 2 15 15 9 3 13 13 1 9 2
27 14 0 9 13 2 16 4 15 0 9 13 9 0 9 1 9 9 0 9 2 9 2 15 9 3 13 2
22 1 9 9 13 9 1 0 9 2 7 3 10 9 2 3 0 9 0 0 9 2 2
10 9 1 11 13 1 10 9 0 9 2
10 9 7 9 3 14 13 7 13 9 2
23 11 2 11 2 13 12 9 2 16 9 13 1 9 9 0 9 2 13 3 1 9 9 2
42 0 9 1 0 9 0 9 9 1 9 13 2 15 0 1 9 13 0 9 1 9 7 9 2 4 13 9 9 14 1 12 9 2 16 13 0 9 0 1 10 9 2
15 1 10 9 0 13 0 9 2 15 13 9 1 0 9 2
16 13 14 12 9 2 16 0 9 13 9 1 0 9 12 9 2
32 15 2 15 15 1 10 9 9 13 3 0 2 13 3 9 2 16 15 0 9 4 13 3 3 2 16 9 13 9 3 0 2
8 13 2 16 0 13 1 9 2
12 10 9 3 13 1 9 2 16 15 15 13 2
7 9 1 9 7 14 13 2
1 11
5 9 11 11 2 11
3 0 9 2
1 9
4 11 11 2 11
31 13 3 3 9 1 15 2 16 13 7 13 13 0 9 13 1 9 2 7 13 15 2 15 13 9 0 9 9 7 9 2
24 13 0 13 2 16 9 9 1 0 9 1 0 12 0 9 1 12 9 9 1 9 3 13 2
31 9 2 3 15 0 2 15 4 3 3 3 13 0 9 1 9 7 0 9 2 7 10 0 9 9 13 1 10 9 13 2
39 3 1 9 2 15 13 13 0 9 2 3 2 9 2 9 2 10 0 9 2 2 13 3 3 1 9 9 9 3 2 16 9 1 15 13 9 0 9 2
10 10 0 9 4 7 13 13 3 0 2
7 3 0 9 13 1 9 2
11 1 0 9 4 0 9 13 0 9 9 2
34 0 9 13 2 16 4 3 12 9 13 13 7 9 2 15 4 13 1 9 10 9 2 7 3 15 13 1 12 0 9 1 0 9 2
7 9 3 13 1 0 9 2
9 7 9 9 13 10 0 9 13 2
9 1 9 15 7 4 13 9 9 2
26 3 3 0 9 0 9 9 1 0 9 13 0 9 1 10 9 9 2 15 15 13 13 0 9 9 2
14 13 0 9 2 16 10 0 9 13 1 0 1 9 2
20 9 9 13 0 9 13 1 9 2 16 1 12 9 13 2 1 0 13 13 2
29 13 9 2 16 4 9 13 13 9 1 9 0 9 3 1 9 0 9 9 1 9 2 7 1 0 9 0 9 2
7 15 13 3 9 0 9 2
24 1 15 7 13 3 9 0 9 1 0 9 1 9 1 0 9 2 15 13 3 0 16 3 2
5 0 9 1 0 9
2 11 2
13 0 0 9 0 9 0 2 11 13 12 9 9 2
27 9 1 9 13 12 9 9 2 16 1 0 9 0 9 3 12 9 9 2 3 13 9 0 9 11 11 2
26 0 9 0 9 2 3 12 5 13 0 0 9 0 2 11 2 13 0 0 9 2 3 12 5 2 2
11 0 9 13 9 9 2 14 12 5 2 2
16 0 9 9 13 9 1 11 2 11 2 11 2 11 7 11 2
18 0 2 11 13 9 9 1 0 9 2 3 2 0 2 11 7 11 2
18 1 9 13 0 9 1 9 0 0 9 11 1 11 1 9 12 9 2
7 0 9 13 3 12 9 2
13 3 13 9 10 9 1 11 3 16 12 12 9 2
5 9 9 9 1 11
4 11 11 2 9
32 1 9 15 13 2 16 1 9 9 9 1 0 9 11 4 3 13 9 9 9 9 2 15 13 1 9 1 9 9 10 9 2
26 9 9 11 1 0 9 3 1 9 13 3 0 2 13 0 9 1 9 10 9 7 13 15 0 9 2
24 0 0 0 9 10 9 13 7 3 12 1 9 9 1 0 9 9 9 7 9 1 15 0 2
42 13 2 14 3 2 1 9 1 0 9 1 9 0 11 2 1 9 0 9 1 11 2 3 4 4 10 3 16 0 9 13 3 3 7 13 4 9 0 9 9 9 2
16 13 4 3 0 9 9 0 9 1 0 9 9 0 0 9 2
21 1 0 9 13 0 15 13 2 16 0 9 9 9 13 1 10 9 0 7 3 2
40 16 13 9 1 9 1 11 1 12 9 2 13 15 3 3 0 9 10 0 9 3 2 7 4 3 13 9 2 1 10 9 1 0 9 15 13 13 0 9 2
21 9 13 2 9 15 3 13 2 1 9 10 9 13 9 0 9 1 0 9 11 2
20 3 13 9 1 9 7 3 7 9 2 16 3 15 3 4 9 13 16 9 2
9 9 13 3 2 9 15 3 13 2
32 16 4 13 10 9 13 1 0 9 9 2 13 0 2 16 9 11 4 13 1 9 9 2 16 4 15 9 3 1 9 13 2
49 15 13 10 9 2 15 9 13 0 9 2 9 9 13 1 9 10 0 9 2 7 15 1 9 0 9 2 9 9 1 9 9 9 2 1 10 10 9 2 7 14 1 15 2 16 4 3 13 2
32 13 2 14 15 9 3 2 16 13 9 10 7 16 4 3 3 13 2 15 3 13 2 13 1 9 7 13 15 1 9 9 2
30 0 9 2 15 13 10 9 0 9 9 9 2 13 9 13 1 0 9 0 9 2 7 13 0 13 15 9 1 9 2
23 13 15 7 2 7 2 7 10 0 9 0 9 1 15 0 9 1 9 11 2 7 13 2
19 13 1 15 9 2 15 10 9 13 2 1 9 0 0 9 1 9 11 2
24 9 11 2 3 1 11 2 7 4 13 9 2 3 1 10 9 13 2 3 3 13 1 11 2
35 7 3 15 3 13 2 13 15 3 3 0 9 2 0 9 0 0 9 1 9 7 10 9 1 11 2 7 7 9 9 11 1 0 9 2
26 16 9 0 2 3 3 0 9 0 9 4 13 13 9 9 2 7 14 9 9 2 16 15 13 0 2
2 9 0
1 9
2 11 11
16 9 13 0 9 9 2 0 0 9 1 9 2 3 0 9 2
9 15 13 3 0 9 1 9 9 2
17 0 13 2 16 15 15 1 9 10 9 13 3 3 16 15 9 2
25 0 9 9 2 0 9 7 0 9 2 15 15 3 13 1 9 7 0 9 2 10 9 14 13 2
6 13 7 0 9 9 2
9 3 13 3 3 0 1 0 9 2
9 13 3 0 7 0 2 7 13 2
16 13 3 1 15 2 16 9 3 13 3 13 9 14 0 9 2
38 13 2 14 9 9 3 9 0 2 3 13 9 9 1 9 2 7 13 9 9 1 10 9 2 13 1 3 16 12 9 11 11 7 13 1 0 9 2
13 16 13 3 9 0 9 9 2 15 13 9 15 2
12 3 16 3 1 9 4 9 3 13 0 9 2
18 15 0 13 9 13 1 9 9 9 7 13 14 15 2 15 9 13 2
23 13 3 3 0 9 0 9 2 15 13 0 9 2 16 4 1 10 9 3 3 3 13 2
9 7 15 1 9 3 0 0 9 2
12 12 9 3 13 0 9 7 1 15 15 13 2
8 1 0 0 9 13 0 9 2
18 3 3 13 0 9 2 15 1 0 9 3 9 13 1 0 0 9 2
14 9 15 1 15 13 3 9 7 10 9 1 9 9 2
28 1 9 1 3 0 0 9 1 12 0 9 13 3 0 13 9 12 9 7 12 0 9 2 15 13 3 0 2
21 13 1 9 2 16 12 1 9 3 1 10 0 9 3 3 3 13 9 2 2 2
10 13 13 9 0 15 0 16 10 9 2
12 14 2 3 0 9 0 7 9 1 0 9 2
18 3 13 2 0 9 7 9 4 13 3 13 14 9 2 7 7 9 2
19 9 0 10 0 9 1 9 3 0 3 13 15 1 9 9 1 0 9 2
10 15 13 7 9 1 9 9 7 9 2
14 3 14 15 2 16 9 13 13 9 9 7 13 9 2
11 9 13 15 2 7 13 3 3 0 9 2
3 9 0 2
4 11 13 0 9
2 11 2
44 3 12 9 0 1 0 9 0 9 2 11 2 3 13 1 11 1 9 0 9 2 15 4 13 13 0 0 7 0 9 2 15 15 3 13 1 9 9 0 9 9 11 11 2
35 11 11 2 9 11 2 0 0 0 9 1 0 2 0 0 2 9 2 13 2 16 16 11 1 9 13 2 4 1 9 9 13 0 9 2
14 0 9 11 13 9 9 7 13 9 1 9 2 13 2
19 15 9 1 9 13 9 11 1 9 2 15 4 4 13 1 9 0 9 2
4 11 13 0 9
2 11 2
44 9 0 9 11 11 3 13 2 16 11 13 13 0 9 2 3 0 9 0 9 1 11 13 9 10 0 9 2 1 10 9 4 1 9 13 9 0 7 0 9 1 0 11 2
9 0 9 13 9 0 9 1 11 2
17 13 15 2 16 10 9 4 13 0 7 3 7 0 2 13 11 2
12 3 13 2 16 11 13 1 0 9 0 9 2
5 9 1 0 0 9
20 0 9 3 0 9 0 9 9 11 13 3 1 0 9 0 0 9 11 11 2
18 16 9 4 13 1 3 0 9 2 13 0 2 16 9 13 0 9 2
8 0 9 2 0 9 2 2 2
11 7 9 9 2 15 3 2 3 13 13 2
18 0 9 2 13 9 9 7 13 2 16 13 1 0 0 9 0 11 2
26 1 9 4 9 9 2 15 13 1 15 3 0 0 9 3 0 1 9 2 13 1 9 1 0 11 2
9 11 11 13 11 0 9 1 0 9
2 11 2
23 0 0 9 0 9 1 11 4 13 1 0 9 11 11 13 0 9 0 9 1 0 9 2
26 9 1 9 1 0 9 3 13 2 16 13 9 1 9 1 0 9 2 15 13 1 15 13 0 9 2
22 11 14 9 13 0 9 2 15 13 1 9 0 9 1 11 2 0 11 1 9 12 2
9 9 13 4 13 1 9 10 9 2
7 0 9 7 9 13 13 2
21 1 0 0 9 4 15 1 11 11 7 11 13 9 2 13 4 0 9 7 9 2
24 13 3 9 1 9 1 11 2 15 16 0 0 9 3 1 9 12 13 1 0 9 0 9 2
20 0 9 11 11 13 10 9 9 1 11 2 16 1 0 9 11 13 0 9 2
16 13 15 3 7 3 13 2 10 9 9 13 1 9 9 9 2
37 9 0 9 11 11 13 3 1 11 9 9 2 16 11 13 1 11 9 2 10 9 13 13 9 1 0 9 9 1 9 9 11 1 9 11 11 2
23 0 9 0 0 9 13 11 11 3 0 1 0 9 0 1 9 0 9 9 9 11 1 11
2 9 11
6 9 1 11 13 3 0
2 11 2
13 0 9 3 13 9 1 9 10 0 9 1 11 2
31 1 9 1 0 0 9 11 13 0 9 11 2 16 9 13 4 13 3 3 2 16 13 1 9 9 9 1 0 0 9 2
21 15 3 1 9 11 13 7 9 0 9 1 0 9 11 2 1 2 11 11 11 2
33 15 3 13 9 0 0 9 9 11 11 7 10 9 2 16 0 9 4 1 11 13 1 0 9 2 16 3 9 9 7 0 9 2
4 9 1 11 13
8 9 9 1 9 15 13 0 9
2 11 2
29 0 9 1 9 9 1 9 15 3 1 9 11 1 9 7 9 1 11 13 2 7 12 0 9 13 1 9 11 2
12 0 9 3 13 9 0 9 0 9 1 0 2
27 0 9 11 1 9 13 0 9 2 16 4 13 11 2 11 7 11 2 0 1 9 11 2 13 9 9 2
34 16 15 3 3 9 13 2 9 11 2 11 2 11 2 11 2 11 2 11 2 11 7 11 13 2 16 13 11 2 7 7 9 13 2
16 1 0 9 11 11 3 13 0 9 9 1 9 14 12 9 2
22 0 9 9 13 1 9 9 7 1 11 2 11 7 0 9 2 15 13 3 0 9 2
19 16 4 13 9 2 9 15 13 1 0 9 2 16 4 13 1 0 9 2
29 9 0 9 2 15 15 13 9 2 13 2 16 7 16 13 9 9 3 0 2 0 9 13 1 9 0 9 9 2
21 3 12 9 9 13 1 9 2 15 1 9 9 13 2 13 9 1 9 11 11 2
9 11 1 0 9 1 9 13 9 2
18 0 9 2 0 0 9 2 9 0 9 7 11 13 9 1 9 9 2
18 3 1 0 9 13 9 9 15 15 13 2 16 13 13 2 13 9 2
14 11 4 3 13 2 16 13 9 9 1 9 7 9 2
22 14 12 9 9 1 9 13 1 9 2 10 9 13 0 9 9 3 1 9 0 9 2
17 13 3 1 9 11 2 0 9 11 2 0 7 0 11 7 11 2
19 0 9 13 3 3 2 7 9 13 1 15 3 0 2 16 3 13 9 2
18 11 2 11 7 11 13 1 9 1 9 0 0 9 7 0 0 9 2
19 3 13 15 1 11 2 3 15 0 9 13 1 12 9 1 9 1 9 2
7 0 9 13 9 9 1 11
2 11 2
21 0 9 1 11 13 9 9 11 2 16 4 13 9 9 0 1 0 2 0 11 2
22 13 15 1 11 0 9 0 9 1 0 11 11 11 2 15 15 13 9 1 0 9 2
26 9 1 11 15 13 0 9 9 9 12 0 9 2 0 9 0 2 11 2 11 2 11 7 11 2 2
21 1 0 9 9 0 9 13 13 9 2 3 13 0 11 1 9 0 9 0 9 2
23 0 9 9 11 11 3 13 1 9 9 1 9 9 0 9 2 15 13 0 7 0 9 2
19 11 7 13 2 16 13 11 13 13 0 9 1 9 9 1 9 9 11 2
24 13 2 16 16 9 13 2 0 9 13 12 9 2 15 13 1 11 7 11 1 0 9 11 2
26 0 9 11 11 13 2 16 11 7 11 1 9 9 0 9 1 0 9 13 10 9 1 11 7 11 2
17 16 3 13 9 1 11 2 10 9 4 3 13 9 9 10 9 2
22 0 9 13 2 16 4 2 14 9 1 9 9 1 11 13 2 13 15 1 9 9 2
5 9 11 15 13 2
6 13 10 9 2 13 2
33 1 9 0 9 1 11 7 11 13 9 9 11 13 0 9 11 11 1 9 2 16 0 11 1 12 2 9 13 0 0 0 9 2
5 11 2 9 1 0
13 9 11 13 1 0 11 2 9 11 11 13 1 11
4 11 11 2 11
38 11 11 2 9 11 11 2 0 9 0 0 9 2 4 12 2 9 3 1 9 10 9 13 1 11 1 9 9 0 9 11 11 16 9 7 0 9 2
18 9 11 11 2 9 0 0 9 2 4 3 10 9 13 1 0 11 2
8 0 9 3 15 13 2 2 2
22 11 4 3 13 9 14 3 2 2 2 13 15 1 9 15 13 2 2 2 13 11 2
11 13 2 16 15 11 13 7 13 15 9 2
9 0 9 9 1 0 9 3 13 2
19 0 9 1 10 9 13 1 9 2 1 15 9 1 9 13 1 15 9 2
8 11 11 15 13 0 9 13 2
24 3 1 9 15 11 13 2 16 13 16 0 9 0 9 9 2 16 10 0 9 1 11 13 2
6 9 11 15 9 13 2
21 13 9 13 9 1 0 9 2 11 3 7 3 13 2 16 11 13 9 0 9 2
24 10 9 4 3 13 7 11 15 13 1 9 9 2 1 15 3 13 11 1 9 11 0 9 2
33 9 9 3 13 0 9 7 16 15 11 13 2 16 0 9 9 13 2 11 13 1 9 7 13 2 1 10 9 0 9 13 9 2
21 13 13 10 9 7 13 15 2 16 4 13 13 2 16 13 2 7 16 13 9 2
10 3 15 15 13 1 11 9 7 13 2
25 16 0 11 13 1 9 7 13 9 15 9 2 9 11 11 11 11 15 13 1 11 1 0 9 2
36 9 7 7 10 0 9 1 11 13 0 0 9 16 0 9 2 7 9 13 0 3 9 2 0 9 11 13 2 16 9 13 0 13 1 9 2
23 1 0 9 13 11 2 16 4 13 0 7 0 9 1 0 7 0 9 1 9 0 9 2
20 0 9 15 3 13 1 15 2 16 11 13 10 9 16 0 2 7 14 0 2
12 11 3 13 11 2 16 15 13 0 9 3 2
10 11 3 13 0 9 1 0 9 9 2
20 11 13 2 16 13 15 3 15 2 15 13 9 1 9 7 9 1 0 11 2
10 11 13 0 7 0 9 3 16 9 2
24 0 9 13 7 10 9 2 16 15 3 7 15 3 13 11 1 0 9 2 15 3 1 15 2
14 11 7 15 0 13 0 9 0 9 11 16 0 9 2
21 3 2 1 11 9 1 9 0 9 2 15 13 1 0 9 1 11 1 0 9 2
14 12 9 4 13 1 0 0 9 1 0 9 0 11 2
15 12 1 15 13 4 13 1 9 1 9 7 9 1 9 2
23 13 15 9 0 9 0 9 1 0 9 2 15 13 12 9 7 13 10 9 1 0 9 2
2 9 11
4 11 3 13 11
2 11 2
18 1 9 1 9 10 0 9 1 0 9 3 13 11 0 9 11 11 2
16 11 1 9 13 11 3 7 9 2 16 4 11 10 9 13 2
44 9 9 0 9 1 0 9 1 9 0 9 1 0 12 1 12 9 4 1 9 11 13 1 9 2 3 4 1 9 11 13 12 9 0 9 2 16 1 0 14 0 12 9 2
23 9 0 9 1 12 0 9 13 1 0 0 9 1 0 9 0 2 11 7 10 9 13 2
13 0 9 3 13 2 16 13 1 9 10 9 13 2
7 13 15 7 1 15 9 2
5 11 13 9 0 9
2 11 2
10 11 13 3 13 9 9 1 0 9 2
27 13 15 1 9 0 9 9 11 11 1 10 0 9 1 0 9 11 11 2 15 13 1 11 1 0 9 2
18 1 0 9 13 11 1 0 9 1 0 9 13 3 12 9 9 9 2
21 1 0 9 15 13 1 12 9 9 7 1 9 12 11 13 12 9 9 0 9 2
38 11 1 9 4 13 14 10 9 2 15 15 9 13 2 7 3 9 0 1 9 0 9 2 3 13 10 9 1 0 9 0 16 9 1 0 9 11 2
6 9 0 9 11 3 13
3 9 11 11
5 7 9 2 7 9
6 11 11 2 11 2 11
22 1 0 9 1 0 9 13 0 2 0 0 9 1 9 11 13 7 13 13 0 9 2
12 1 0 0 9 13 1 0 9 9 9 9 2
20 1 9 15 15 15 13 2 13 9 11 7 13 9 9 1 9 1 0 9 2
29 3 1 10 9 13 9 1 12 9 0 9 1 0 9 0 9 2 9 15 13 1 0 9 7 9 15 15 13 2
7 13 15 7 14 0 9 2
21 3 13 11 0 0 9 1 9 2 3 13 1 15 3 14 0 9 2 13 3 2
24 7 1 0 9 9 1 0 0 9 11 7 11 14 9 1 10 9 13 1 0 9 0 9 2
11 1 15 13 15 3 3 3 0 16 3 2
18 1 9 2 3 4 13 2 16 15 13 0 9 2 13 9 1 9 2
17 14 3 9 13 0 10 9 0 9 7 9 9 2 13 0 9 2
22 0 9 1 9 9 13 13 9 2 15 15 13 1 9 1 9 2 9 7 0 9 2
24 14 9 1 9 1 9 0 9 13 12 2 9 2 3 3 0 0 9 13 3 16 12 9 2
16 1 3 12 9 0 0 9 0 11 13 3 16 12 12 9 2
17 1 0 9 7 0 9 11 13 11 10 0 9 7 0 9 13 2
9 1 9 9 15 3 13 13 9 2
8 9 7 0 9 9 7 13 2
18 0 9 13 2 16 13 9 7 9 13 3 1 9 0 13 3 9 2
4 9 3 13 2
40 9 4 7 13 1 0 9 0 2 16 11 2 0 9 11 1 9 2 3 3 13 9 1 9 7 3 15 13 2 13 9 0 9 1 0 9 1 9 11 2
17 9 1 9 1 9 3 15 1 0 9 13 9 9 1 0 9 2
11 9 9 1 9 13 10 9 0 9 11 2
4 15 13 9 2
17 10 9 13 1 12 9 2 1 0 0 9 3 3 15 13 9 2
21 15 13 9 2 16 13 1 9 3 3 9 7 3 13 1 10 9 9 3 13 2
7 9 9 13 1 15 3 2
22 13 15 13 3 7 3 2 16 4 15 1 15 15 13 2 13 9 2 0 1 11 2
19 1 11 3 3 13 3 10 9 2 0 9 15 13 1 9 1 12 9 2
9 9 1 9 13 3 10 9 3 2
13 3 1 9 9 0 9 0 9 3 13 9 9 2
9 1 11 3 13 0 9 9 13 2
24 15 2 15 3 13 11 2 13 14 9 2 9 13 9 2 15 3 2 13 12 1 9 11 2
26 0 9 1 10 9 13 9 15 9 1 0 11 16 9 1 10 0 9 0 0 9 0 2 0 9 2
17 0 9 1 9 13 9 1 9 9 1 9 9 1 11 7 11 2
11 1 9 9 15 1 0 11 13 13 15 2
24 12 1 3 0 9 13 7 0 2 0 9 2 3 1 9 0 0 0 9 2 13 0 9 2
7 11 3 13 11 1 9 2
11 9 11 15 13 7 1 15 15 13 11 2
7 13 0 9 1 0 9 2
14 9 15 13 2 16 3 2 14 3 2 13 9 11 2
17 13 1 0 9 1 9 0 11 2 3 12 1 0 9 1 9 2
12 9 9 1 9 1 0 9 0 9 15 13 2
7 0 9 9 13 9 9 2
15 14 0 9 13 1 0 9 0 9 7 13 1 15 9 2
22 14 10 9 9 1 15 2 1 0 9 1 9 11 2 1 12 1 9 13 0 9 2
4 3 16 3 2
4 11 13 1 9
9 1 9 13 1 0 0 0 9 9
21 0 9 13 0 12 9 0 0 9 13 1 12 9 0 12 9 10 0 0 9 2
23 11 2 0 0 0 9 2 15 13 1 0 9 1 9 7 9 0 2 11 1 9 11 2
16 3 12 9 10 9 13 1 11 7 1 12 9 13 0 9 2
21 1 0 9 13 11 9 1 9 0 2 0 2 0 2 0 7 1 9 0 9 2
11 0 9 13 0 0 9 1 0 0 9 2
16 9 9 2 15 13 1 9 2 15 13 9 7 13 0 9 2
12 9 4 13 0 9 2 0 9 13 0 9 2
5 9 13 0 9 2
13 9 13 0 7 0 2 9 1 11 13 0 9 2
10 0 9 13 12 9 0 0 9 11 2
22 13 15 1 9 9 2 9 2 9 2 9 2 9 0 2 2 2 9 7 0 9 2
25 9 3 3 13 1 9 0 9 2 1 15 15 15 13 1 0 9 3 13 0 9 9 1 0 2
29 1 0 0 9 7 10 0 0 9 13 3 0 9 11 1 9 0 9 1 9 12 9 0 2 0 7 0 9 2
21 1 9 12 2 9 13 0 2 0 9 2 10 9 13 13 9 9 1 9 11 2
11 0 9 13 3 1 9 12 0 0 9 2
14 1 9 1 9 12 15 7 9 11 13 1 0 9 2
28 1 12 9 3 11 13 13 0 9 2 16 1 15 4 3 13 9 0 9 9 7 3 7 9 10 0 9 2
25 9 1 9 1 10 9 2 0 1 0 11 1 0 9 7 15 12 9 2 15 7 3 13 13 2
9 9 11 7 11 15 1 9 13 2
28 1 9 12 0 9 9 11 13 9 1 9 2 15 13 9 11 16 0 9 7 13 9 12 9 1 0 9 2
17 9 13 0 9 12 1 12 9 9 2 16 0 9 13 3 13 2
14 1 0 0 9 1 0 9 15 0 9 9 3 13 2
28 0 9 2 9 0 1 9 9 7 9 10 9 2 15 9 13 1 0 9 2 13 0 12 12 9 0 9 2
5 0 9 1 0 9
10 9 1 11 3 13 9 0 2 0 9
6 11 11 2 9 9 11
17 0 9 3 3 13 0 9 1 0 9 1 0 9 7 0 9 2
22 3 1 15 2 13 1 9 2 3 1 0 9 13 0 0 9 2 3 10 0 9 2
49 9 1 0 9 2 9 7 9 9 11 11 2 11 2 13 1 0 9 2 15 13 3 9 2 15 3 13 9 9 2 1 15 15 0 9 13 1 9 2 1 0 9 7 3 13 7 0 9 2
12 1 9 1 0 0 9 13 0 7 0 11 2
49 11 11 2 11 15 13 1 9 13 3 3 16 3 2 3 15 0 9 11 13 1 9 9 2 9 0 9 2 0 9 11 2 4 1 10 0 9 13 14 1 0 9 2 7 3 1 0 9 2
33 0 9 2 15 15 11 13 2 13 3 13 3 1 11 2 13 7 10 0 9 13 2 16 9 0 2 0 9 13 3 1 9 2
17 1 9 12 9 13 0 9 3 1 0 0 9 13 3 0 9 2
36 15 0 2 0 9 2 0 11 7 9 11 11 2 13 2 16 9 2 15 15 1 12 2 9 13 1 0 0 9 2 15 3 13 0 9 2
10 9 9 13 9 13 0 9 16 0 2
29 0 9 13 1 11 7 3 7 1 9 0 9 2 13 3 2 16 0 9 4 13 3 16 1 9 0 0 9 2
23 16 7 1 9 0 0 2 0 9 13 9 2 9 1 0 9 13 9 10 9 2 2 2
34 0 9 3 13 9 2 16 9 13 13 0 9 2 7 13 0 9 1 15 2 16 4 1 10 9 13 9 2 15 4 13 9 9 2
27 0 9 1 11 3 13 0 9 1 9 0 9 2 1 9 13 1 15 2 10 0 9 13 13 0 9 2
22 10 3 0 9 13 0 2 0 9 13 14 1 9 2 3 4 1 0 9 13 9 2
18 9 11 1 11 13 1 9 9 2 15 11 7 11 1 0 9 13 2
30 12 9 15 13 1 9 2 7 11 2 15 15 15 3 13 13 2 3 13 1 3 0 9 2 15 9 13 0 9 2
23 0 9 7 1 9 1 11 13 12 0 9 2 13 1 12 9 10 0 9 1 10 9 2
5 1 15 15 13 2
14 13 2 16 9 0 9 1 0 9 13 3 0 9 2
15 1 12 9 13 9 11 11 1 11 1 9 0 0 9 2
21 0 9 1 11 13 14 14 13 1 11 9 2 15 13 1 15 0 16 1 9 2
24 13 2 4 13 15 2 15 4 13 11 2 13 2 3 15 14 13 11 1 10 9 0 9 2
9 13 12 0 9 2 3 15 13 2
12 1 0 2 0 9 13 7 13 1 0 9 2
6 7 15 0 13 0 2
13 13 4 3 13 2 16 15 13 9 7 9 9 2
16 7 1 0 2 0 9 15 13 2 16 1 15 13 0 9 2
16 13 3 1 15 2 16 15 9 11 4 1 10 0 9 13 2
4 11 11 0 9
2 11 11
46 1 0 9 11 11 13 2 15 13 1 12 0 0 9 9 12 1 9 9 1 11 2 0 9 13 3 3 7 1 0 9 15 2 15 15 13 10 9 2 3 10 0 9 2 2 2
20 13 0 13 0 9 2 13 15 1 9 1 9 2 10 9 15 13 2 2 2
24 9 0 9 1 9 13 9 1 15 2 16 16 16 4 13 9 9 2 13 15 10 0 9 2
29 9 0 9 13 1 10 9 3 0 9 1 9 12 7 9 2 9 13 13 9 0 9 0 15 10 0 9 0 2
8 1 12 9 13 0 9 0 2
36 10 0 9 15 1 9 3 13 9 13 9 0 9 1 9 3 2 16 9 0 15 13 10 0 9 2 1 15 3 13 9 2 15 15 13 2
11 9 13 14 12 1 10 9 2 3 0 2
67 9 1 11 15 3 2 13 15 2 13 9 11 11 1 9 7 1 0 9 1 9 12 13 15 0 9 0 9 7 13 15 9 1 9 2 3 9 7 9 2 9 1 9 7 9 2 0 0 9 2 9 9 2 0 9 2 0 2 14 0 9 2 0 9 2 9 2
7 0 9 15 15 3 13 2
37 1 9 0 9 2 0 2 9 9 2 12 2 11 2 11 13 2 1 15 13 10 0 9 2 15 13 9 2 15 13 9 0 15 1 10 9 2
28 13 15 15 9 2 15 1 9 13 1 9 3 2 4 13 9 0 1 9 7 9 7 4 1 9 3 13 2
23 13 15 1 9 1 15 2 16 13 0 9 9 2 15 15 1 15 1 9 7 9 13 2
30 10 9 13 0 9 1 9 9 13 7 16 3 0 9 0 9 1 9 2 1 15 11 3 3 13 9 1 9 12 2
36 11 11 13 2 9 3 13 12 9 2 9 0 9 13 14 15 2 16 9 1 0 9 15 13 13 9 10 9 2 7 7 15 2 16 13 2
21 16 15 13 0 9 2 15 13 9 7 13 15 15 2 16 10 9 13 1 0 2
19 9 2 9 2 9 7 9 2 15 13 0 9 9 2 0 1 0 9 2
22 11 1 10 9 13 9 2 15 13 2 16 4 15 13 1 0 9 16 0 2 9 2
5 7 15 3 9 2
22 13 3 0 9 10 9 1 9 13 9 13 10 9 1 0 9 2 7 3 15 13 2
35 16 3 13 10 9 10 9 1 0 9 2 16 15 13 0 9 7 9 1 0 9 2 13 15 9 2 15 4 14 3 11 11 13 9 2
15 16 4 14 2 3 4 14 13 1 9 1 9 0 9 2
7 7 13 3 1 10 9 2
37 7 10 9 13 13 3 9 9 9 2 0 15 1 0 9 2 15 15 13 10 0 9 9 1 9 2 7 3 13 15 2 15 1 9 9 13 2
23 13 4 15 13 3 9 1 9 2 15 10 9 13 0 9 2 16 15 10 9 3 13 2
7 7 13 3 7 0 9 2
18 10 9 4 13 10 9 13 2 13 15 3 13 10 9 2 10 9 2
51 1 0 9 11 13 2 3 4 13 1 9 2 16 4 13 0 9 11 2 0 9 4 1 9 1 9 13 15 9 7 9 1 9 2 15 4 3 4 13 1 9 2 3 13 7 13 1 9 7 9 2
19 1 9 4 15 13 3 2 16 10 9 4 3 1 9 0 9 15 13 2
16 3 15 1 15 1 9 13 2 16 4 0 9 11 3 13 2
20 1 0 9 15 13 2 16 1 10 0 9 9 0 2 9 13 1 0 9 2
25 13 1 15 3 13 7 15 2 16 9 13 13 1 11 9 1 0 9 2 16 13 9 0 9 2
10 13 9 9 2 15 15 1 15 13 2
19 7 15 3 9 2 3 9 2 15 13 13 7 4 1 15 13 0 9 2
4 13 15 9 2
15 13 2 16 7 0 0 9 4 15 13 13 1 12 9 2
13 1 0 9 13 0 13 9 2 16 4 15 13 2
25 15 13 0 9 15 0 9 2 3 3 13 9 2 15 13 0 9 7 3 12 1 0 13 9 2
32 0 9 13 7 1 9 2 15 14 1 9 13 9 0 9 2 9 2 16 13 10 9 2 4 13 9 0 9 3 14 13 2
21 10 9 15 13 2 16 4 13 1 9 11 1 10 9 2 16 4 15 13 3 2
25 7 1 15 2 16 1 0 0 9 14 3 9 13 9 0 9 2 13 3 13 11 3 1 9 2
5 13 15 0 9 2
24 9 10 9 13 13 2 3 3 2 16 10 9 4 13 1 0 9 7 4 15 13 9 9 2
22 13 2 16 15 3 3 7 3 13 10 0 9 3 13 1 9 3 7 3 0 9 2
37 13 2 14 0 9 9 2 0 9 13 15 2 7 15 13 13 2 16 4 15 3 13 2 16 10 7 15 9 13 0 13 7 3 13 1 9 2
11 15 13 7 9 0 9 2 9 1 9 2
9 9 0 9 9 13 1 15 0 2
17 1 9 13 12 0 0 7 0 9 1 0 2 0 7 0 9 2
22 10 9 13 0 2 1 0 13 10 9 2 7 15 3 13 9 9 2 13 3 0 2
34 0 13 0 9 2 3 9 2 1 15 9 13 13 0 2 0 9 15 2 15 13 1 15 0 2 3 13 7 13 3 1 9 13 2
31 1 10 9 13 9 0 9 9 0 2 16 10 9 2 15 4 15 3 13 2 13 3 13 9 2 1 15 15 9 13 2
14 13 7 0 0 9 13 15 9 9 9 1 0 9 2
15 0 13 13 1 15 2 16 4 0 9 9 13 3 0 2
64 0 0 9 15 13 1 15 2 15 15 4 13 2 16 13 1 11 2 15 4 3 13 13 11 2 1 9 13 3 3 14 12 9 2 9 9 13 2 9 1 9 15 13 1 9 2 7 16 9 13 2 15 13 9 0 9 2 4 13 7 9 2 2 2
16 7 0 9 15 3 13 2 16 7 15 13 1 9 0 9 2
47 13 15 1 15 2 16 9 9 13 2 13 1 15 0 2 16 13 15 9 2 0 9 7 9 9 3 2 16 4 3 1 9 13 2 16 4 11 15 13 13 0 9 7 10 9 13 2
35 0 9 15 3 13 13 3 2 16 4 10 9 13 13 0 9 2 13 13 1 9 9 1 12 9 7 13 1 9 9 9 1 9 0 2
18 7 7 1 10 9 7 9 13 15 3 2 3 15 0 9 3 13 2
22 3 0 9 13 9 9 2 15 15 13 9 9 2 9 2 9 0 9 2 9 3 2
52 10 9 2 1 9 16 13 0 2 15 13 1 9 7 9 9 2 15 13 11 11 1 15 2 16 4 9 10 9 13 1 9 0 9 2 13 3 0 9 7 15 15 13 13 1 10 0 9 7 0 9 2
13 10 9 7 13 1 9 9 7 9 1 10 9 2
19 3 2 15 2 16 15 13 1 15 2 16 4 15 13 2 9 3 13 2
15 13 4 0 9 2 7 15 15 13 2 16 4 15 13 2
4 1 15 13 2
8 1 0 9 7 1 10 9 2
10 1 15 9 13 11 10 0 9 13 2
3 13 13 2
27 13 9 9 10 2 15 15 13 13 9 2 15 4 13 2 13 15 13 14 3 2 16 15 1 9 13 2
17 11 3 13 2 15 13 2 7 15 2 15 13 2 3 13 9 2
15 13 13 10 9 2 13 10 9 7 13 3 13 1 11 2
25 3 13 15 3 2 15 13 9 9 2 15 13 13 7 15 15 15 13 13 2 16 4 15 13 2
10 16 10 9 3 13 1 9 0 9 2
16 15 1 15 2 7 15 1 15 2 7 3 15 1 9 15 2
35 3 9 9 13 14 1 0 9 1 10 9 2 13 15 9 3 15 0 9 2 15 7 13 0 13 1 9 2 16 4 15 13 1 9 2
14 15 3 13 2 16 4 15 9 13 2 15 13 13 2
19 1 11 11 15 13 2 15 13 7 9 0 9 16 10 9 7 0 9 2
40 0 0 9 13 1 10 9 2 7 16 15 9 7 9 0 15 1 0 9 4 13 10 9 2 13 15 3 2 13 2 14 1 15 3 13 7 9 0 9 2
6 13 3 2 16 13 2
10 1 0 9 13 9 0 9 3 0 2
33 13 4 3 1 0 9 1 11 1 0 9 7 0 9 15 1 15 3 13 1 10 9 2 15 3 13 9 2 7 3 15 13 2
19 0 15 3 13 2 16 9 15 13 1 0 9 7 10 0 7 0 9 2
25 13 15 1 0 9 2 0 9 2 13 3 2 16 15 13 1 15 2 15 13 15 0 16 15 2
29 9 13 1 0 9 7 13 15 13 1 15 0 16 13 9 2 9 2 9 1 9 2 9 9 7 9 1 9 2
15 13 0 0 9 7 13 1 9 2 16 13 1 10 9 2
9 0 9 13 0 7 0 9 9 2
41 13 14 13 2 16 1 9 3 0 1 9 3 13 10 0 9 2 3 4 15 13 1 9 2 1 15 13 2 13 4 3 15 15 0 15 2 1 15 15 13 2
9 1 9 2 9 2 9 7 0 9
7 11 11 2 0 9 0 9
23 10 0 9 13 12 2 12 2 9 2 16 0 9 13 13 9 1 0 9 1 12 9 2
5 10 9 13 0 2
22 9 10 9 1 9 0 13 2 13 7 13 2 3 15 13 13 7 7 1 9 13 2
14 13 4 15 14 9 7 0 9 2 7 7 10 9 2
16 9 1 9 1 9 0 13 1 0 9 7 13 15 3 13 2
36 9 1 0 0 9 2 16 13 0 9 2 3 2 1 11 0 2 9 2 9 2 2 13 0 9 2 1 15 15 13 0 9 1 9 9 2
34 10 0 7 0 9 15 13 1 9 0 7 9 15 13 13 3 1 9 0 9 1 0 0 0 9 0 1 10 9 2 3 7 3 2
21 13 13 1 0 9 1 0 9 9 9 2 3 1 9 0 2 0 7 0 3 2
21 3 13 9 13 10 9 7 1 0 9 9 3 0 2 1 10 9 1 9 0 2
17 13 2 14 9 0 9 0 3 3 2 13 15 13 7 10 9 2
19 0 9 0 9 13 9 1 0 0 9 2 3 9 13 9 0 0 9 2
16 13 0 2 16 10 9 0 9 13 7 13 13 9 3 0 2
17 0 9 0 1 0 9 2 7 15 14 0 9 2 13 1 9 2
20 9 15 3 13 12 9 9 3 0 2 1 15 1 12 9 13 9 9 0 2
23 1 0 9 15 9 13 1 9 9 9 2 13 3 1 9 3 0 7 1 9 9 0 2
6 1 9 9 3 13 2
21 1 0 9 15 9 13 1 0 9 9 0 9 1 9 2 15 9 13 3 13 2
31 13 1 15 0 9 2 4 13 0 9 2 3 0 9 2 1 0 9 2 9 3 13 7 13 13 15 3 13 7 13 2
26 10 9 15 13 13 2 16 13 1 9 9 1 9 0 2 16 1 10 9 13 13 9 9 10 9 2
13 13 0 2 16 7 9 1 9 0 13 13 3 2
19 10 9 2 9 7 0 9 15 9 13 1 12 2 0 7 12 9 0 2
20 10 9 2 16 1 15 13 15 0 9 2 15 13 1 9 2 15 13 9 2
39 7 3 10 9 13 15 2 15 9 3 13 2 9 1 9 1 0 9 1 12 9 7 1 0 0 9 2 16 4 15 15 13 9 0 9 1 9 0 2
21 9 3 13 2 1 15 9 2 3 0 9 3 0 0 9 1 0 0 9 13 2
21 13 13 9 9 2 7 3 1 10 9 10 9 9 13 2 16 4 9 9 13 2
31 1 0 9 3 10 9 13 2 16 0 9 15 13 9 9 9 1 9 0 2 15 3 13 7 13 3 1 0 9 9 2
14 13 15 2 16 3 13 9 15 2 16 13 9 0 2
47 15 2 16 9 13 9 1 10 9 2 16 13 13 10 9 1 0 9 2 10 9 4 3 13 2 7 15 13 9 9 2 15 9 13 9 1 9 0 2 13 16 10 9 0 0 9 2
27 13 2 16 9 0 9 9 1 9 9 13 0 9 0 0 9 1 9 1 0 9 2 3 13 9 0 2
16 10 9 9 7 9 13 10 9 2 7 0 9 15 0 9 2
29 9 2 15 9 9 13 2 13 1 15 2 16 13 0 13 10 0 0 9 7 3 2 3 3 15 13 0 9 2
22 13 15 16 9 1 9 0 15 9 2 7 1 15 9 2 3 1 9 1 9 9 2
47 9 2 15 15 13 0 9 1 0 0 9 1 9 12 7 12 7 13 9 1 0 9 1 0 9 1 0 9 10 9 10 2 16 15 9 3 13 1 0 9 2 15 3 10 9 13 2
44 3 3 2 9 2 15 15 1 9 9 1 12 13 2 16 15 0 9 3 13 10 9 2 13 9 12 2 12 2 12 1 0 0 9 1 0 0 9 12 5 9 9 12 2
9 9 9 13 12 2 12 2 12 2
17 9 15 13 1 0 9 1 0 0 9 1 0 0 9 12 5 2
24 9 13 0 9 1 0 9 9 12 2 12 2 12 2 9 4 13 1 12 2 12 2 12 2
15 0 9 1 9 1 0 9 7 1 0 4 13 9 12 2
59 13 2 14 0 9 3 1 0 9 1 0 9 9 1 0 9 2 7 1 0 9 2 10 2 9 2 9 12 5 2 2 13 1 12 2 12 2 12 1 12 2 12 2 12 3 3 9 12 2 3 9 3 12 7 12 5 0 9 2
72 1 10 9 15 2 15 13 12 9 9 13 2 14 13 2 9 2 15 13 3 4 13 2 7 15 13 9 13 15 1 9 1 10 9 0 2 3 2 1 9 1 0 9 1 0 9 2 2 15 2 15 13 13 10 9 10 0 9 2 13 2 16 9 9 2 9 7 0 9 3 13 2
14 11 2 9 12 9 2 2 3 0 9 3 1 11 2
9 1 9 0 9 2 3 0 9 2
1 9
8 11 2 13 12 2 7 3 12
5 11 11 2 11 11
13 1 9 1 11 13 0 7 3 0 9 2 11 2
12 9 2 15 13 1 0 9 3 9 0 9 2
22 3 15 7 13 2 16 11 13 3 14 0 11 2 7 3 0 9 2 9 0 9 2
18 7 16 15 2 15 15 13 1 9 9 2 13 10 9 3 7 3 2
12 0 9 13 14 1 9 0 16 11 1 11 2
13 13 3 0 0 9 7 0 9 0 0 0 9 2
12 7 0 0 9 13 1 9 9 3 16 11 2
19 9 15 3 13 14 3 3 2 7 15 3 14 1 9 9 1 0 9 2
13 1 15 0 13 9 2 15 13 14 12 9 9 2
22 9 15 13 7 13 3 16 9 1 9 2 16 9 2 7 3 16 0 9 1 9 2
20 0 9 9 13 1 9 1 9 13 7 7 1 0 9 15 14 3 13 9 2
12 0 9 13 0 9 7 13 13 1 0 9 2
18 1 9 3 13 3 3 2 1 9 3 3 1 0 9 13 0 9 2
11 11 2 3 16 11 2 13 0 9 9 2
22 1 15 3 13 3 15 2 15 3 13 0 0 9 2 14 3 0 7 14 3 0 2
9 2 13 15 0 2 7 0 2 2
10 3 9 9 9 3 13 3 0 9 2
2 0 9
13 1 9 13 11 2 3 16 10 9 2 0 9 2
17 9 10 9 13 3 0 3 1 9 2 7 3 1 0 0 9 2
8 0 9 13 7 9 0 9 2
14 0 7 3 12 1 0 9 11 15 13 1 9 9 2
11 1 0 12 9 0 9 15 13 14 12 2
16 1 0 7 0 9 1 9 15 13 1 0 9 3 9 9 2
15 3 0 0 9 2 15 9 13 2 15 0 9 3 13 2
26 13 2 16 9 13 0 9 2 7 7 13 1 9 10 9 0 9 3 9 9 2 7 3 15 13 2
19 9 11 13 1 0 9 3 1 9 2 15 15 1 0 9 3 3 13 2
7 7 3 13 10 10 9 2
10 9 13 3 0 9 1 9 0 9 2
4 9 0 7 0
26 9 2 15 3 13 3 1 9 12 1 11 2 15 1 0 9 0 9 1 11 13 3 10 9 9 2
16 7 15 14 9 1 0 9 11 12 2 2 7 1 11 3 2
24 11 15 10 0 9 1 0 9 13 7 3 2 3 15 1 15 13 12 12 9 9 0 9 2
12 1 9 9 15 13 3 0 11 2 0 9 2
17 9 1 11 13 10 9 11 9 12 7 10 9 13 3 16 0 2
15 16 1 9 12 13 2 4 9 13 7 13 7 0 9 2
8 10 9 13 0 7 0 9 2
20 13 9 7 9 2 15 15 3 13 0 7 0 9 9 2 1 15 13 9 2
25 3 13 1 0 9 9 0 9 7 9 0 9 2 15 15 13 3 1 9 1 9 9 7 9 2
17 0 9 10 9 13 0 0 9 2 9 2 9 7 0 0 9 2
13 1 12 2 1 12 2 9 13 0 9 0 9 2
8 1 9 13 15 0 7 0 2
15 1 9 1 9 15 3 9 3 13 9 9 0 7 0 2
23 11 15 13 14 1 9 1 0 9 2 7 1 9 0 9 13 0 9 0 9 0 11 2
14 1 9 1 15 13 1 0 7 3 0 9 0 9 2
13 9 0 9 13 3 3 0 9 11 2 0 9 2
19 1 9 15 0 2 11 13 10 9 13 0 9 2 15 15 7 13 13 2
20 7 7 11 13 1 9 9 7 9 2 13 12 2 7 3 12 2 13 9 2
12 9 15 1 9 13 1 9 9 7 0 9 2
7 7 7 3 10 9 13 2
25 13 9 2 9 2 9 7 0 9 2 3 15 2 15 4 13 1 11 2 13 1 15 0 9 2
11 3 15 3 9 9 13 3 1 9 9 2
2 9 11
25 0 0 9 13 3 1 9 12 1 9 9 0 9 2 15 13 1 10 9 3 0 1 0 9 2
12 0 9 11 12 2 13 0 9 7 0 9 2
12 1 0 9 15 7 11 13 13 0 9 9 2
17 11 2 15 15 13 1 9 7 1 9 2 1 15 13 0 9 2
9 3 13 11 14 0 9 1 11 2
16 0 9 13 13 9 2 7 7 15 15 13 11 2 9 2 2
12 9 12 11 13 7 3 3 13 9 0 9 2
11 13 0 9 9 2 15 4 13 0 9 2
7 13 7 1 0 0 9 2
6 11 13 9 0 11 2
10 7 1 10 9 11 13 10 9 13 2
13 13 9 0 9 2 9 9 9 7 3 7 9 2
12 0 9 13 7 1 9 0 7 0 9 11 2
8 11 3 13 0 9 7 9 2
11 9 12 2 9 3 13 3 15 9 9 2
6 9 1 9 2 9 9
27 1 9 0 9 13 1 9 12 11 1 0 11 2 9 0 11 2 1 9 13 0 9 7 0 9 9 2
5 3 7 4 13 2
17 1 9 12 1 9 0 2 9 1 9 4 11 13 1 0 11 2
14 9 0 9 13 1 0 9 0 9 2 13 0 13 2
24 1 0 9 12 2 9 13 0 0 9 0 11 2 0 9 2 1 9 9 11 11 2 11 2
6 13 9 9 1 9 2
14 3 0 9 0 9 1 9 9 13 10 9 1 9 2
13 9 1 9 11 13 1 0 12 9 3 0 9 2
18 0 0 11 2 9 9 2 13 10 0 9 1 9 1 0 9 11 2
15 3 13 1 3 0 9 1 0 9 2 15 13 9 13 2
39 1 9 1 0 9 9 13 0 9 0 11 2 0 9 2 2 1 10 9 13 1 9 12 9 11 0 2 15 15 2 2 0 9 7 9 0 0 9 2
13 9 13 7 1 9 2 9 9 13 9 0 9 2
15 1 9 12 0 9 13 0 9 7 13 9 1 0 9 2
19 0 9 7 13 1 0 9 2 3 13 9 1 0 0 9 13 1 9 2
18 10 9 7 3 13 1 0 9 7 3 0 9 0 9 11 0 9 2
16 9 13 0 9 1 9 12 2 1 15 11 13 0 0 9 2
15 1 0 9 1 0 9 13 9 13 7 12 10 9 13 2
9 1 0 9 13 11 0 0 9 2
18 0 9 7 13 13 1 11 2 13 15 1 0 9 7 13 0 9 2
6 3 3 13 11 9 2
15 13 0 0 9 2 11 2 2 15 13 0 9 1 11 2
18 15 3 1 0 9 13 0 9 2 15 1 11 13 1 9 1 9 2
17 1 9 12 13 11 10 0 9 2 11 13 9 2 9 13 11 2
10 13 3 0 9 0 11 7 0 11 2
8 9 11 13 11 1 0 9 2
13 0 9 1 0 11 4 3 13 14 1 9 12 2
6 11 3 2 11 1 9
25 1 0 2 0 9 1 9 12 2 3 9 9 13 0 9 2 13 1 11 12 7 9 9 9 2
20 9 0 0 9 7 1 9 9 13 1 9 12 1 12 9 3 12 9 11 2
14 3 13 1 9 2 3 15 13 1 9 11 7 11 2
18 16 15 15 13 0 2 13 3 1 9 1 12 9 9 1 0 9 2
16 1 0 9 15 13 3 7 0 9 11 11 2 11 7 11 2
9 0 11 13 3 3 12 0 9 2
10 1 0 9 13 13 9 7 0 9 2
12 13 1 15 3 3 16 12 7 12 12 9 2
19 7 15 13 9 0 0 9 9 2 3 3 0 9 13 13 7 0 9 2
8 9 3 13 9 9 10 9 2
24 9 13 14 10 3 0 9 2 16 3 2 0 0 9 2 0 9 9 9 11 1 9 11 2
20 9 13 0 0 0 9 1 0 9 7 9 2 9 13 0 9 7 0 9 2
6 11 2 9 9 7 9
11 1 9 1 11 13 11 9 9 7 9 2
14 9 2 13 15 3 1 12 9 2 15 13 1 9 2
42 16 1 0 13 1 9 3 11 2 0 9 7 0 9 2 1 15 0 13 9 11 11 2 11 11 11 2 11 11 11 2 11 11 2 11 11 7 0 0 0 9 2
13 10 0 9 15 13 13 12 9 0 9 1 9 2
10 11 7 11 3 13 1 10 9 0 2
31 13 15 14 0 9 10 9 2 7 3 9 2 9 2 9 2 9 1 9 7 9 2 7 3 7 9 9 0 10 9 2
9 0 0 9 11 13 3 11 11 2
19 1 11 13 10 11 2 0 12 9 9 12 11 2 0 9 0 9 3 2
18 0 9 4 1 15 2 16 13 3 1 9 2 3 9 13 1 11 2
27 9 2 0 1 0 0 9 2 3 13 7 3 1 9 3 3 0 2 7 16 0 9 7 9 13 0 2
11 10 9 13 2 16 1 9 15 3 13 2
12 3 11 15 13 11 7 11 13 11 1 11 2
9 0 9 15 1 0 3 3 13 2
4 13 0 9 2
14 3 9 13 3 0 9 2 3 15 13 1 15 9 2
8 9 9 1 9 13 3 0 2
40 1 9 0 0 9 13 1 10 9 9 2 16 13 11 0 10 0 9 11 2 11 13 9 3 0 2 0 7 0 9 2 0 9 7 3 7 0 0 9 2
8 10 9 13 9 3 12 9 2
12 13 15 1 9 1 9 7 13 1 15 9 2
14 1 0 0 9 4 13 13 7 0 0 9 7 9 2
16 3 15 13 1 0 9 7 9 2 3 15 13 7 0 9 2
25 1 0 9 15 11 13 3 7 1 0 9 2 13 13 0 9 0 12 7 9 11 11 2 11 2
8 7 11 13 14 9 7 9 2
13 0 9 9 13 3 16 10 0 9 13 0 9 2
18 0 13 3 0 0 9 2 15 9 2 15 0 9 7 3 0 9 2
8 1 0 9 13 12 0 9 2
21 0 0 11 7 0 0 2 11 11 2 3 13 16 9 11 11 2 9 0 9 2
16 0 9 0 11 13 3 0 9 11 12 2 3 1 9 9 2
23 16 9 13 13 2 16 9 2 1 15 13 0 9 2 13 1 9 9 1 9 0 9 2
4 9 1 0 9
13 0 9 13 1 11 1 12 9 1 9 0 9 2
29 1 10 9 13 1 0 9 2 16 1 9 9 2 7 1 9 9 7 11 2 15 15 13 3 10 12 0 9 2
17 1 0 9 1 0 11 15 13 2 16 4 13 3 13 1 9 2
10 0 9 13 1 0 9 9 1 9 2
2 9 9
13 11 2 11 11 13 3 0 9 0 9 0 9 11
1 9
3 9 1 9
1 9
35 9 2 1 9 2 3 1 15 9 13 3 1 12 9 2 13 13 9 9 11 11 9 16 0 9 2 13 0 9 2 9 2 3 3 2
5 13 15 7 13 2
11 9 9 11 13 3 3 3 1 0 9 2
40 16 15 1 0 9 2 3 9 13 9 2 13 1 10 0 9 2 3 3 16 12 9 3 0 9 13 14 13 2 15 15 13 13 9 1 9 9 7 9 2
15 7 3 0 15 0 9 13 0 9 1 0 9 0 9 2
40 15 2 15 13 1 9 0 9 0 9 9 7 9 1 9 9 2 13 1 9 9 9 0 9 2 9 9 7 9 2 0 9 2 0 9 9 2 0 9 2
12 13 3 1 9 2 15 13 0 9 0 9 2
8 9 15 7 13 1 0 9 2
22 3 16 13 3 2 13 9 0 7 13 9 15 2 15 13 9 1 9 10 0 9 2
13 11 13 1 9 16 1 0 2 0 7 0 9 2
19 13 9 1 9 10 9 7 1 9 2 15 15 0 9 13 10 9 13 2
37 9 13 9 1 0 9 13 1 15 0 2 16 0 0 9 1 9 2 3 0 7 0 0 9 2 13 1 0 9 3 1 0 9 3 3 13 2
10 11 11 11 11 2 9 16 0 9 2
18 13 9 9 2 11 12 2 12 9 2 9 13 2 0 9 12 9 2
10 13 9 16 9 2 9 13 1 9 0
11 1 0 9 0 9 11 11 1 9 0 9
35 1 9 12 9 9 2 0 1 9 7 0 9 1 9 12 7 12 2 15 1 0 12 9 13 3 9 2 0 9 9 7 0 9 9 2
66 0 9 2 15 15 1 9 12 2 9 13 1 0 9 0 9 3 7 15 13 9 12 0 9 9 1 9 1 9 0 1 0 0 9 7 1 0 0 9 1 10 0 9 15 0 9 1 0 9 2 13 9 14 1 9 10 9 2 7 1 0 9 1 0 9 2
51 9 0 7 1 9 0 15 3 1 0 9 14 7 0 2 9 2 9 2 9 7 9 2 15 13 9 1 10 1 9 9 0 9 2 15 13 13 1 11 11 2 0 9 11 0 1 9 0 9 2 2
29 9 4 1 0 9 1 9 1 9 12 9 9 13 9 2 16 13 0 7 0 9 2 7 9 0 9 1 15 2
25 0 9 13 2 16 3 13 7 13 1 9 13 0 9 2 16 3 1 0 2 7 0 0 9 2
12 1 15 13 10 0 9 1 9 0 7 0 2
34 0 9 13 15 2 16 1 9 1 10 9 13 3 3 13 9 2 1 15 9 4 9 13 7 9 15 15 4 13 1 9 7 13 2
24 3 13 15 9 12 2 12 2 12 2 12 7 12 9 2 7 13 4 13 7 0 7 0 2
9 10 9 15 9 13 7 4 13 2
33 9 13 10 0 9 9 2 16 1 3 0 9 13 1 0 9 13 2 13 13 0 9 2 2 9 10 9 9 13 9 0 9 2
24 1 9 9 1 9 15 13 2 16 3 9 0 9 13 9 2 16 1 15 13 10 0 9 2
25 1 9 0 9 13 15 9 0 9 2 1 15 4 3 13 9 10 9 2 3 2 0 9 2 2
11 15 13 9 1 9 10 12 0 9 9 2
39 3 9 0 9 13 1 9 1 9 7 1 9 0 15 0 9 1 9 1 0 9 13 15 2 16 9 9 1 10 9 2 3 4 13 0 2 13 0 2
11 9 9 0 9 13 3 0 9 0 9 2
25 1 10 9 9 13 15 10 9 2 7 16 4 15 3 2 3 1 9 0 0 9 2 13 0 2
8 9 13 9 13 10 0 9 2
17 9 13 13 0 9 0 11 1 9 12 1 12 5 0 0 9 2
28 1 9 10 9 3 13 0 9 9 7 9 1 15 7 0 0 9 9 13 2 9 9 7 9 13 10 9 2
15 1 15 9 0 13 10 9 9 0 9 1 9 7 9 2
32 9 10 9 13 0 7 9 12 9 2 7 9 12 9 2 3 9 1 9 2 16 4 10 9 9 0 9 1 9 13 2 2
20 9 0 1 10 9 0 9 15 3 13 3 9 2 15 4 13 1 9 0 2
27 14 2 13 3 1 12 0 9 9 0 1 9 12 7 12 1 9 0 1 0 0 9 7 0 0 9 2
14 9 9 13 0 1 9 2 3 4 9 1 9 13 2
20 10 9 4 3 13 1 15 2 16 4 15 1 15 13 13 9 1 0 9 2
17 9 15 7 13 13 7 1 9 9 1 0 9 7 1 0 9 2
12 3 15 13 9 2 3 9 13 9 0 9 2
8 9 3 1 10 10 9 13 2
27 13 3 1 9 13 1 9 2 1 9 0 0 9 2 3 0 9 2 16 15 4 13 0 9 0 9 2
19 15 7 4 13 9 10 9 0 1 10 12 9 9 2 0 9 0 9 2
28 15 13 3 9 0 9 1 9 9 7 9 15 1 15 2 3 16 15 13 0 9 0 1 0 0 9 2 2
11 3 13 9 0 0 9 7 0 0 9 2
6 13 13 9 1 15 2
28 16 4 9 13 1 0 0 9 2 13 15 2 16 1 0 9 10 9 13 9 0 9 0 7 9 3 0 2
12 1 3 1 9 9 2 9 13 3 0 9 2
26 10 9 0 9 13 11 3 1 0 9 10 9 2 3 13 2 3 16 0 9 2 1 0 0 9 2
10 10 9 4 13 1 0 2 0 9 2
29 0 7 13 2 16 0 0 9 15 13 1 9 1 0 9 2 13 3 9 10 9 7 1 9 1 15 15 13 2
31 1 15 4 0 13 2 16 1 0 9 13 0 9 10 0 9 3 3 2 7 15 1 12 2 9 7 1 12 2 9 2
26 10 9 13 0 9 1 9 9 1 9 1 0 9 2 15 13 9 9 0 10 9 1 3 0 9 2
15 9 0 9 1 9 3 13 7 9 0 9 1 9 2 2
11 13 15 3 1 9 9 1 9 0 9 2
10 1 9 1 15 13 1 9 0 9 2
27 3 7 3 2 16 0 9 1 9 9 9 13 0 1 9 2 15 13 13 1 9 2 16 9 13 9 2
26 1 10 9 1 9 1 0 0 9 7 0 0 9 4 9 0 9 1 9 0 9 13 3 1 9 2
21 0 9 13 2 16 9 15 13 13 9 3 1 9 12 9 3 2 16 13 9 2
17 16 4 15 10 9 13 1 9 0 9 2 4 4 15 13 9 2
25 9 9 3 13 9 1 10 0 9 13 0 2 3 15 13 9 2 15 13 0 7 13 15 13 2
12 0 0 9 1 9 0 9 1 9 13 4 2
20 13 3 1 0 9 2 16 3 2 16 13 15 3 1 9 13 2 13 9 2
21 3 9 9 1 9 4 15 4 13 0 9 2 15 15 3 13 7 15 15 13 2
36 1 9 7 3 7 1 0 13 13 15 2 16 10 9 9 4 13 1 9 0 9 1 9 0 9 2 3 1 0 9 9 7 0 9 2 2
28 9 12 0 9 2 1 15 15 11 13 2 7 13 1 9 9 0 1 9 0 3 0 0 9 0 9 9 2
33 1 9 13 3 3 0 2 16 9 13 9 2 7 15 0 0 9 4 13 1 0 9 2 7 2 3 12 2 7 3 12 9 2
32 16 9 1 0 9 3 13 7 3 1 9 9 13 9 0 9 2 13 1 15 9 9 1 9 0 9 1 0 9 10 9 2
24 13 15 2 16 10 9 1 0 9 4 13 0 0 9 3 0 12 9 1 9 9 10 9 2
38 10 9 9 2 15 3 13 2 7 7 15 13 0 0 9 1 9 9 2 11 10 9 13 7 3 2 7 1 12 2 9 12 15 3 4 13 2 2
18 13 15 1 9 2 3 0 9 13 7 0 9 1 9 7 9 13 2
5 15 4 13 3 2
21 9 13 9 3 1 9 7 9 4 13 10 0 9 2 3 1 10 9 13 2 2
12 13 9 9 10 0 9 9 9 1 0 9 2
21 14 2 9 1 9 0 0 9 2 3 9 2 3 13 13 9 2 13 10 2 2
10 13 15 7 1 9 9 3 0 9 2
7 10 0 9 15 9 13 2
42 13 0 2 16 0 9 1 9 12 7 12 5 13 3 2 13 14 1 0 9 2 7 7 1 10 0 9 2 9 2 3 16 13 7 9 0 0 9 1 10 9 2
50 11 13 9 2 15 4 0 13 3 0 0 9 2 13 7 0 0 9 1 9 2 0 9 2 9 2 1 0 0 9 2 7 9 0 1 11 3 1 12 9 2 15 13 13 1 9 3 0 9 2
11 1 10 9 13 9 14 12 0 9 3 2
12 9 1 10 0 9 13 7 0 9 9 9 2
24 10 9 9 15 3 13 1 15 2 15 13 10 9 13 3 2 7 13 15 3 1 0 9 2
27 1 10 9 2 15 13 0 0 9 2 13 1 9 1 9 0 9 9 0 1 9 0 1 0 0 9 2
18 15 4 7 13 0 0 9 2 15 1 9 13 12 7 12 5 3 2
3 2 11 2
8 9 3 1 11 13 12 9 9
4 0 9 15 13
8 11 3 13 0 0 9 11 2
39 3 16 12 0 7 0 9 3 0 9 2 15 13 11 2 11 9 2 11 12 7 11 11 2 13 0 9 7 0 9 1 0 1 2 11 9 11 11 2
17 1 9 11 4 1 0 9 13 9 0 9 2 15 0 9 13 2
18 9 15 1 15 4 13 13 3 3 3 1 9 9 0 9 9 12 2
25 11 13 3 13 0 9 10 0 9 1 1 2 11 9 3 9 10 9 2 7 9 9 15 13 2
22 9 11 13 13 9 9 1 0 9 1 0 9 7 0 9 14 1 9 1 0 9 2
19 4 13 7 0 9 2 9 1 0 0 9 9 7 9 13 9 1 9 2
22 13 3 4 13 9 1 9 9 11 11 2 9 11 2 1 9 1 9 1 9 9 2
1 3
23 9 13 1 11 1 0 9 9 12 9 9 2 15 13 1 12 9 3 16 1 0 9 2
6 9 13 14 1 9 12
11 15 13 1 0 9 1 9 2 13 15 13
2 11 2
34 9 12 9 9 2 15 13 13 9 9 2 15 13 10 9 2 16 13 0 0 9 2 13 0 9 1 10 9 13 1 9 9 12 2
21 13 15 3 9 10 0 9 3 1 9 2 16 10 9 13 0 9 1 0 9 2
39 0 9 1 0 9 2 15 9 1 10 9 13 1 9 0 9 2 13 1 15 2 16 9 13 13 13 15 10 0 9 1 9 0 9 0 9 9 9 2
14 15 15 13 3 9 9 0 9 9 2 3 0 9 2
20 1 0 9 13 9 1 0 2 0 2 9 3 0 9 1 9 12 9 3 2
17 9 1 9 9 13 9 1 0 9 14 3 1 0 9 1 9 2
37 9 9 12 13 9 1 0 9 2 3 4 15 10 9 13 4 13 1 0 0 9 2 15 9 1 0 9 7 9 10 9 4 13 1 0 9 2
31 1 9 1 9 3 1 9 4 3 13 13 9 9 1 9 1 10 9 3 3 3 3 2 16 1 9 13 1 10 9 2
35 9 9 0 7 0 9 11 11 2 11 3 11 13 2 16 9 2 15 1 0 9 13 2 15 13 13 2 16 15 13 9 1 9 9 2
24 3 3 4 11 13 0 9 2 11 2 11 13 1 15 2 16 1 10 9 15 3 3 13 2
26 9 0 9 13 9 15 2 16 0 9 10 9 13 3 0 9 1 9 7 0 9 13 1 15 13 2
20 1 9 15 13 9 9 2 7 9 4 13 1 9 7 9 1 15 13 9 2
31 1 0 9 13 0 9 2 15 13 3 12 9 2 0 9 2 1 12 12 0 9 2 1 15 12 12 4 13 0 9 2
5 9 9 11 15 13
2 11 2
28 1 9 9 0 9 0 11 11 15 12 2 9 4 13 1 9 9 2 9 1 11 2 2 15 13 9 9 2
12 9 4 13 1 12 9 7 13 1 12 9 2
29 9 9 13 13 9 0 9 9 2 13 0 7 3 13 0 9 2 13 15 9 7 9 7 1 15 15 3 13 2
31 1 9 9 13 0 9 2 9 1 9 7 1 9 0 9 2 0 9 2 0 9 2 0 9 2 9 9 7 3 9 2
4 0 9 13 9
4 11 2 11 2
40 9 9 1 9 2 9 2 9 2 0 0 9 11 9 2 0 9 0 0 2 7 11 2 13 9 0 9 2 13 11 11 2 11 11 1 0 9 0 9 2
10 13 2 16 10 9 3 13 0 9 2
40 1 9 1 0 9 0 9 13 2 16 9 9 2 9 2 9 2 4 3 13 2 7 3 1 9 0 9 1 0 9 1 0 9 9 2 15 13 0 9 2
22 9 1 0 0 9 15 13 2 16 9 1 0 9 4 13 13 10 0 9 10 9 2
20 16 13 2 0 2 11 11 13 3 1 0 9 2 15 3 13 1 0 9 2
22 3 15 13 2 16 0 9 4 13 9 9 1 9 9 0 0 9 0 0 2 11 2
3 9 14 13
2 11 2
15 9 0 0 9 13 0 9 13 9 7 0 0 9 13 2
8 11 15 13 9 9 11 9 2
10 1 0 9 13 11 12 9 9 9 2
10 11 2 11 13 10 9 1 3 0 2
13 0 9 9 11 13 2 16 13 2 0 9 9 2
4 0 9 13 9
2 11 2
26 1 9 9 9 0 9 7 0 9 13 13 0 9 2 15 3 13 9 10 9 0 9 1 0 9 2
14 16 13 10 9 2 1 0 0 9 13 14 12 9 2
8 3 13 7 9 3 0 9 2
18 9 2 15 1 9 13 9 2 13 13 0 2 7 13 7 1 9 2
16 10 0 9 13 13 9 9 9 9 7 0 9 1 10 9 2
17 1 0 9 13 2 16 9 0 9 13 0 0 9 1 15 9 2
6 9 9 13 3 9 9
22 0 9 9 15 14 13 0 9 2 1 15 0 9 13 9 9 2 7 3 15 3 13
17 9 9 1 0 9 13 1 9 9 2 9 1 0 0 9 2 2
31 0 9 1 9 13 7 9 9 9 2 1 0 9 2 2 1 15 13 3 11 9 11 7 11 9 11 2 11 2 11 2
12 7 9 1 9 15 13 1 9 13 0 9 2
11 7 1 9 15 2 16 13 1 0 9 2
38 12 1 10 9 3 2 1 15 3 9 4 13 2 16 13 1 0 9 7 1 0 9 2 13 9 9 2 3 0 0 9 2 3 0 0 9 2 2
7 9 0 9 13 11 11 2
25 13 0 9 2 15 13 1 9 2 3 0 2 9 9 9 1 0 9 9 11 2 11 7 11 2
11 0 0 9 3 13 7 9 11 7 11 2
15 9 13 9 9 1 3 0 9 9 2 7 15 0 9 2
12 7 15 3 13 13 2 15 13 10 9 13 2
84 1 10 2 3 3 4 9 13 2 13 1 9 9 12 9 2 9 9 1 9 2 15 3 2 15 3 10 9 13 2 2 0 9 9 1 12 9 2 9 13 0 9 9 9 7 13 9 0 1 9 0 2 3 0 9 2 12 9 15 3 13 1 10 10 9 2 7 3 9 9 12 9 7 0 9 2 0 3 1 9 2 9 2 2
11 12 0 9 13 1 0 9 9 12 9 2
10 10 0 9 13 9 0 1 9 9 2
18 13 9 3 13 13 15 1 0 12 9 2 7 7 3 1 15 3 2
15 3 0 13 13 9 1 3 0 0 9 2 0 9 2 2
6 15 15 3 3 13 2
32 13 7 1 0 9 9 2 15 3 3 13 1 9 0 0 9 2 9 1 9 2 1 0 9 9 9 1 9 3 2 2 2
9 9 15 3 7 13 1 0 9 2
13 1 12 2 9 13 13 9 13 9 9 1 9 2
26 13 15 15 3 2 16 15 9 13 13 1 9 3 0 9 7 13 15 3 0 9 2 0 2 9 2
34 10 9 13 9 9 2 0 0 0 9 2 3 0 0 9 2 7 13 3 1 9 9 9 0 9 9 2 1 0 0 9 1 11 2
33 3 9 12 2 9 7 0 9 13 2 16 9 9 13 10 9 9 2 7 7 13 2 3 1 9 2 3 3 1 9 2 9 2
16 15 13 9 1 0 0 0 9 2 7 9 1 0 9 9 2
40 1 0 9 2 16 4 9 2 13 3 3 2 2 13 9 1 0 9 2 16 4 15 9 2 13 15 2 7 3 2 7 0 9 16 4 13 9 0 9 2
31 15 3 13 0 9 9 1 9 2 0 9 2 2 7 13 0 9 0 9 1 9 2 0 9 2 2 15 13 3 0 2
8 0 9 9 13 9 0 9 2
14 13 15 3 9 0 2 3 4 15 15 13 14 3 2
18 1 0 9 3 13 13 12 7 3 9 3 2 7 15 3 13 9 2
25 16 7 9 13 0 9 12 9 2 13 15 3 13 2 16 9 0 1 15 3 13 1 9 0 2
8 1 0 9 4 9 13 3 2
17 3 14 0 9 9 13 9 9 1 9 1 9 2 3 1 9 2
32 0 9 13 3 0 2 13 9 1 0 0 9 2 16 13 9 7 9 2 7 13 15 9 2 15 13 9 1 9 9 9 2
28 3 13 0 0 9 2 15 13 0 9 2 13 1 15 9 2 15 1 15 3 13 2 7 13 15 1 9 2
13 3 1 0 0 9 9 4 0 9 13 12 9 2
17 10 9 13 3 10 3 0 0 9 2 1 15 15 0 9 13 2
17 1 9 3 9 13 7 13 9 1 9 2 7 3 12 9 3 2
13 13 7 10 0 9 2 15 3 1 15 13 9 2
22 9 13 1 15 2 16 3 0 9 15 3 1 9 0 1 0 9 9 13 9 0 2
17 9 9 4 13 13 13 0 9 9 9 9 1 9 0 12 9 2
54 13 7 10 0 9 2 15 13 1 9 9 13 2 1 3 0 2 0 9 1 3 0 9 2 14 1 0 2 9 13 9 0 14 1 9 9 2 15 9 13 13 2 10 9 13 3 1 3 0 9 3 0 2 2
28 13 0 2 16 3 16 0 9 15 9 13 0 9 2 1 15 0 9 13 9 9 2 7 3 15 3 13 2
38 7 2 7 1 15 13 3 10 9 1 0 2 13 15 2 3 0 9 2 9 0 9 13 3 3 15 2 16 15 13 13 13 7 0 9 0 9 2
2 0 9
10 16 9 13 4 9 9 12 1 11 2
20 1 9 2 15 15 9 13 2 13 7 9 1 9 12 2 9 9 1 9 2
13 0 9 0 9 2 9 0 1 9 0 0 9 2
20 1 9 4 15 7 3 13 2 13 1 9 2 1 9 9 15 13 0 9 2
8 13 2 3 13 9 11 11 2
4 13 12 9 2
11 1 9 9 13 0 9 7 13 11 9 2
3 9 13 2
6 15 4 13 1 11 2
12 1 9 0 9 13 1 9 9 1 0 9 2
22 2 14 2 3 13 2 16 0 9 13 0 9 2 2 13 0 9 9 1 0 9 2
11 1 0 9 15 15 3 1 11 13 3 2
27 1 9 13 9 2 0 9 1 9 1 9 9 15 13 3 1 15 2 2 9 2 13 13 2 2 2 2
13 1 9 0 9 1 11 3 13 0 9 11 11 2
14 16 0 9 0 9 4 13 3 9 3 15 13 11 2
19 3 2 7 1 11 10 9 4 13 10 9 1 0 9 0 9 1 11 2
8 7 11 11 3 13 10 9 2
20 16 13 1 9 2 9 0 9 1 0 9 15 4 3 13 1 9 10 9 2
10 13 13 9 1 0 9 10 0 9 2
19 9 9 0 1 9 0 9 7 1 9 15 13 2 16 1 9 13 9 2
21 3 16 15 13 13 2 16 4 1 11 13 12 9 0 9 0 0 7 0 9 2
12 1 15 13 7 0 0 9 1 9 1 11 2
12 9 2 0 9 9 2 15 3 13 1 9 2
6 0 13 7 3 0 2
27 0 9 0 9 11 2 9 15 3 13 10 9 1 9 11 2 9 1 0 0 9 2 0 9 11 2 2
21 3 4 12 2 9 12 0 9 10 0 0 9 9 9 1 0 9 11 11 13 2
40 9 11 11 2 3 2 2 11 11 7 11 11 13 9 9 2 1 9 0 0 9 2 7 9 0 11 2 9 11 11 2 3 2 13 10 9 1 0 9 2
4 0 1 9 11
2 11 2
14 0 9 11 11 11 7 10 9 13 9 9 11 11 2
15 11 13 3 0 9 2 10 9 11 13 1 0 9 9 2
19 9 13 11 3 1 0 9 9 9 1 9 11 1 10 0 9 9 11 2
20 9 13 1 15 2 16 11 13 12 12 9 10 9 2 3 9 9 2 3 2
5 11 10 9 13 2
16 0 9 3 16 11 3 13 9 12 0 9 0 2 0 9 2
5 11 13 9 0 9
4 11 2 11 2
30 0 9 11 11 2 13 1 15 3 2 0 2 0 7 0 2 0 9 2 13 1 10 9 9 9 9 9 2 12 2
9 13 15 15 3 9 1 0 9 2
27 1 9 13 13 9 2 1 9 12 12 9 2 7 9 2 13 4 13 12 9 9 1 9 2 0 9 2
21 9 9 11 11 11 13 0 9 1 0 9 1 9 12 1 0 0 9 1 11 2
22 1 0 9 0 9 11 11 2 15 4 1 9 2 12 13 2 13 11 7 0 9 2
19 9 9 9 2 12 13 1 11 2 11 0 3 14 1 9 11 2 11 2
29 9 11 11 9 15 7 3 13 15 2 16 0 9 1 11 13 0 11 2 1 15 15 9 13 13 1 0 9 2
48 1 9 11 2 16 0 9 9 2 12 13 13 13 9 1 11 7 0 9 2 1 9 1 0 9 13 2 2 9 9 11 11 2 11 13 2 16 9 3 3 0 0 9 4 13 3 0 2
10 9 1 9 0 9 13 7 1 0 2
15 2 3 13 1 15 0 9 1 0 9 2 2 13 11 2
11 11 11 13 12 1 0 9 9 7 9 2
8 3 15 13 7 1 9 9 2
15 1 0 9 15 11 13 14 1 9 1 9 9 2 12 2
23 11 3 4 1 9 9 2 12 2 9 2 12 7 9 2 12 13 1 0 9 0 9 2
23 9 1 15 13 9 1 9 9 2 1 15 2 10 9 13 1 9 2 3 11 13 13 2
28 16 1 11 13 11 2 3 3 2 1 11 13 1 10 0 9 2 11 2 11 7 11 2 7 7 1 11 2
21 1 12 9 9 2 1 15 1 9 12 11 13 9 2 13 12 9 1 11 11 2
7 9 0 11 13 3 9 0
2 11 2
18 0 9 2 1 15 4 13 9 0 11 2 15 13 9 9 10 9 2
14 1 9 11 15 3 13 9 0 9 9 9 11 11 2
20 13 2 16 9 9 1 0 7 9 9 13 7 3 13 9 0 9 1 9 2
17 0 2 0 9 2 7 2 9 3 2 2 13 0 9 9 9 2
52 1 15 2 16 15 0 9 1 9 9 13 2 1 11 13 2 16 0 9 13 13 7 3 13 0 9 1 9 7 10 9 2 16 13 1 9 13 3 2 3 1 10 9 2 3 0 9 13 1 0 9 2
15 0 9 1 9 13 9 9 9 9 9 1 11 11 11 2
32 1 15 1 9 13 0 2 16 15 0 9 2 15 4 13 9 0 11 2 13 3 1 9 2 3 7 1 9 9 0 11 2
5 11 1 9 3 2
1 13
2 11 2
20 14 1 9 0 0 9 15 11 11 2 0 9 11 2 4 1 10 9 13 2
13 13 15 3 1 9 1 11 10 0 9 11 11 2
22 13 3 9 2 16 11 11 13 1 15 2 16 4 13 1 9 11 11 1 9 3 2
21 2 3 3 2 16 10 9 1 9 9 11 13 2 4 10 9 13 2 2 13 2
33 11 11 13 9 2 16 1 0 9 11 9 4 9 13 0 9 2 15 4 13 9 0 9 1 9 11 7 9 2 9 2 9 2
5 16 4 0 9 13
4 11 11 2 11
4 0 9 1 11
10 0 9 13 1 9 9 11 12 2 12
2 11 2
31 0 9 9 9 11 2 15 13 0 9 2 13 3 1 11 1 9 11 11 14 1 9 2 7 3 1 9 9 9 9 2
28 0 9 3 13 0 9 11 12 2 12 2 12 2 12 2 7 1 12 2 9 0 9 11 15 13 0 9 2
27 11 13 1 12 9 9 9 2 11 3 1 10 9 13 9 7 3 1 12 2 9 9 1 0 9 13 2
28 3 12 0 9 15 1 10 9 1 12 2 9 13 0 9 11 2 1 0 9 12 0 9 2 3 12 2 2
33 2 11 3 13 2 11 13 0 2 2 3 13 1 9 11 2 7 16 3 10 9 15 0 9 9 13 0 9 14 3 1 9 2
25 3 0 9 11 2 12 2 9 2 12 2 12 2 13 9 9 2 15 3 13 9 9 16 9 2
33 1 12 2 9 13 11 3 1 12 9 2 12 2 12 2 2 7 13 15 15 9 7 11 12 9 11 13 2 12 2 12 2 2
37 14 12 9 1 9 11 13 9 2 16 11 12 9 1 15 2 12 2 12 2 13 0 9 2 9 15 3 13 1 9 2 1 9 7 9 2 2
24 2 11 13 16 11 2 16 15 13 1 9 2 13 7 13 10 9 2 2 13 0 9 11 2
21 11 9 13 2 12 2 12 2 2 11 13 9 2 7 3 3 14 0 9 13 2
38 2 3 15 13 9 9 2 2 13 15 9 11 2 11 1 9 2 3 12 9 1 9 10 9 13 12 2 12 2 13 9 7 0 9 13 1 9 2
9 7 1 9 15 13 3 9 11 2
21 2 11 13 0 9 2 15 4 15 9 1 15 13 1 0 9 3 1 9 3 2
16 12 0 9 4 13 3 9 2 2 13 1 9 9 11 11 2
2 11 13
2 11 2
16 0 0 0 9 11 11 15 13 0 9 1 9 9 1 11 2
24 11 13 9 0 2 11 7 11 2 7 15 9 13 0 9 12 7 12 9 0 0 0 9 2
29 11 3 13 2 16 13 0 13 1 15 0 9 9 0 0 9 2 7 1 10 0 9 13 0 13 1 9 9 2
3 1 0 9
26 11 11 2 12 2 2 0 9 9 11 0 7 11 11 2 15 13 0 9 9 0 0 9 0 11 2
13 13 15 3 0 12 9 3 2 3 13 11 11 2
1 3
24 11 11 2 9 0 9 1 11 2 13 1 9 1 11 2 15 13 1 9 2 0 11 11 2
4 9 1 0 9
10 9 11 13 1 9 0 11 12 2 12
2 11 2
26 14 1 0 9 1 0 9 13 0 9 0 9 1 0 9 1 11 0 0 9 11 11 12 2 12 2
21 1 0 9 1 0 9 13 3 3 11 2 15 15 1 9 9 13 7 12 9 2
26 1 0 9 3 13 1 9 9 9 13 11 2 7 13 9 2 3 16 1 9 3 11 1 0 9 2
25 12 9 1 9 15 9 13 9 12 2 12 9 11 2 15 1 0 9 13 9 7 13 9 11 2
18 3 1 15 15 1 0 9 13 0 9 2 7 7 10 9 13 9 2
14 9 13 1 0 9 0 9 2 7 3 1 0 9 2
13 11 13 9 9 7 9 9 1 9 13 1 9 2
17 11 7 1 10 9 9 13 13 2 15 15 15 13 3 9 9 2
12 9 7 11 13 13 9 7 0 9 13 9 2
21 9 13 9 9 2 15 13 0 9 2 9 15 13 7 13 0 9 12 2 12 2
2 11 2
4 9 2 11 2
6 9 2 11 2 11 2
6 9 2 12 2 12 2
19 9 11 11 11 2 2 9 13 10 9 2 7 16 15 13 1 0 9 2
8 15 15 13 13 7 1 9 2
13 9 13 14 3 0 2 10 9 7 9 13 9 2
20 3 13 0 16 15 2 1 0 9 7 13 10 9 1 9 7 9 3 2 2
3 9 13 11
2 11 2
16 9 0 11 11 11 9 13 1 0 0 9 0 9 11 11 2
17 2 0 4 15 1 9 13 1 10 9 2 2 13 9 2 9 2
19 11 1 9 13 9 1 0 11 7 3 3 13 2 16 15 13 13 3 2
29 2 3 16 15 7 9 11 4 13 2 16 1 9 13 3 3 9 7 16 15 13 3 15 13 2 2 13 11 2
3 3 1 11
6 0 9 1 11 7 11
2 11 2
17 9 0 9 11 11 13 1 9 1 9 1 9 9 9 10 9 2
45 10 9 1 15 2 16 15 13 13 15 0 9 1 11 2 7 9 0 9 13 14 1 9 1 11 2 12 2 12 2 2 7 11 2 12 2 12 2 2 13 3 9 0 9 2
15 2 13 1 15 1 9 2 10 9 13 1 0 9 9 2
45 10 9 1 9 9 0 13 3 0 2 9 9 13 3 3 9 2 2 13 15 11 0 9 1 10 9 1 9 11 2 7 3 13 2 16 10 9 13 13 3 0 9 1 11 2
32 3 15 13 7 9 9 2 7 9 0 9 9 2 9 11 2 11 11 15 7 1 9 1 9 1 11 13 1 11 3 3 2
46 13 1 15 2 16 11 13 0 9 9 1 9 2 13 14 0 7 1 0 0 9 2 7 1 9 13 1 9 1 9 9 11 11 11 2 10 0 9 13 1 10 9 1 9 0 2
38 9 0 9 9 11 3 13 2 16 7 1 11 2 15 13 16 0 9 1 9 2 15 13 0 9 1 0 9 2 3 2 1 11 1 9 12 2 2
17 2 13 2 16 1 0 9 13 0 13 7 11 2 2 13 11 2
20 9 1 11 7 3 4 13 2 11 15 3 3 13 1 9 11 16 0 9 2
25 0 4 1 11 13 2 16 4 11 10 9 1 9 9 9 13 7 15 4 9 1 10 9 13 2
6 1 0 9 14 10 9
2 11 2
26 0 9 11 4 3 13 9 0 9 11 9 7 11 11 1 9 9 0 9 0 1 9 12 1 9 2
23 9 13 3 3 13 2 1 9 13 4 9 1 9 13 1 0 9 2 13 0 11 2 2
17 9 0 9 11 11 3 13 12 9 2 3 16 0 9 11 11 2
16 13 15 9 13 10 9 2 15 1 9 1 9 12 13 13 2
29 9 15 13 3 1 9 0 9 11 11 2 15 9 3 1 9 9 3 13 2 13 1 15 7 1 0 9 2 2
11 0 9 13 1 0 9 1 9 0 9 2
18 1 9 11 13 0 9 1 9 9 2 1 15 13 13 10 0 9 2
13 9 3 1 11 13 9 7 13 3 1 0 11 2
3 1 11 13
2 11 2
14 0 9 13 0 9 0 9 1 11 1 11 7 11 2
30 1 0 9 2 3 15 0 9 13 1 12 2 9 9 9 1 9 11 2 13 0 9 1 11 1 0 9 9 9 2
11 13 13 9 7 10 9 13 1 0 9 2
12 13 13 9 7 3 0 9 9 9 3 13 2
13 1 0 9 4 3 9 13 7 9 9 9 13 2
25 11 2 11 2 12 2 12 2 2 11 11 2 9 11 2 2 1 9 7 1 9 9 13 0 2
18 12 1 9 0 9 11 15 13 2 16 13 0 9 1 9 11 2 2
12 11 11 2 9 11 2 2 13 4 9 9 2
20 1 0 9 0 4 13 3 2 0 13 9 0 9 12 1 12 1 9 2 2
9 11 2 11 2 12 2 12 2 2
25 11 11 2 9 11 2 2 13 4 1 9 9 0 2 3 15 15 9 13 7 3 4 9 13 2
19 10 9 1 0 9 9 7 13 1 9 9 2 7 1 9 4 13 0 2
8 0 9 15 13 1 9 2 2
28 11 0 2 9 11 2 2 1 11 13 3 0 9 2 3 4 13 12 2 12 2 7 9 1 9 13 9 2
20 1 0 9 13 2 16 4 1 9 12 2 12 1 9 13 1 12 2 12 2
6 3 15 9 13 2 2
26 11 2 11 2 12 2 12 2 2 11 11 2 9 11 2 2 13 4 3 7 1 11 0 1 9 2
12 13 7 13 2 16 11 13 0 9 0 9 2
9 10 0 9 15 13 14 13 2 2
20 11 11 2 9 11 2 2 16 13 15 13 2 3 9 11 7 11 1 9 2
11 9 3 14 0 12 9 1 9 9 2 2
36 11 2 0 2 11 2 12 2 12 2 2 11 11 2 9 11 2 2 1 9 4 13 1 0 9 7 1 10 9 13 0 9 1 9 2 2
29 11 11 2 9 0 2 11 2 2 0 9 1 9 9 13 2 16 4 13 1 0 12 0 9 1 10 9 2 2
34 11 2 11 2 12 2 12 2 2 11 11 2 9 11 2 2 13 4 3 2 7 16 4 1 12 9 13 13 14 1 0 9 9 2
17 13 9 9 2 15 3 1 12 9 1 0 0 9 13 13 2 2
19 11 11 2 9 11 2 2 1 12 9 4 3 13 7 9 15 3 13 2
10 3 4 3 13 9 14 0 0 9 2
17 13 9 1 10 9 13 9 1 9 9 2 7 9 13 0 2 2
4 9 9 1 11
8 12 1 9 13 1 9 1 9
5 0 9 11 7 11
26 11 2 0 9 11 11 13 1 0 9 1 11 0 0 9 1 9 1 12 9 9 12 2 12 9 2
15 0 0 0 9 12 2 12 13 10 9 11 1 9 12 2
21 16 0 15 1 0 9 13 1 0 0 9 1 9 1 12 9 9 11 11 11 2
9 9 12 13 0 9 1 12 9 2
18 3 0 1 0 9 11 0 9 11 15 9 12 13 1 9 0 9 2
15 1 9 1 9 13 0 11 11 11 9 12 9 14 0 2
17 9 11 11 13 9 1 9 12 9 2 15 13 0 0 0 9 2
3 11 1 9
3 0 11 2
30 0 9 0 9 9 9 12 11 11 11 2 12 9 2 1 11 15 13 7 1 10 0 9 11 11 13 1 9 9 2
12 11 13 9 9 7 3 3 15 13 13 9 2
9 9 1 15 13 9 13 15 0 9
2 9 2
25 0 9 3 13 7 1 0 9 7 3 1 0 9 0 7 0 9 13 9 7 10 9 1 9 2
27 3 16 13 13 1 10 9 2 15 3 0 9 13 1 10 9 1 9 7 3 13 9 1 9 0 9 2
42 1 9 0 9 2 3 9 3 13 9 1 9 1 9 2 16 1 9 13 3 3 14 12 7 16 13 9 13 15 9 2 4 13 10 0 9 7 13 15 1 9 2
22 1 9 13 2 2 13 2 13 2 2 7 1 15 0 9 2 3 13 1 9 2 2
21 9 15 13 7 3 13 2 16 15 15 15 13 2 7 16 9 9 13 3 3 2
18 13 4 2 16 16 13 0 2 13 4 13 0 9 0 3 10 9 2
11 3 15 13 1 9 2 13 9 7 13 2
12 3 3 4 15 13 10 9 2 13 2 13 2
5 3 13 1 9 2
7 9 13 9 1 9 9 2
11 0 9 13 2 9 1 10 0 9 3 2
16 9 13 9 2 9 2 1 0 9 9 2 2 9 7 9 2
11 9 0 12 10 9 13 7 1 9 9 2
10 15 13 9 2 15 15 16 9 13 2
14 15 15 13 1 9 1 0 2 3 15 16 9 13 2
11 15 13 9 2 13 9 1 15 0 9 2
8 15 13 9 2 13 15 13 2
11 13 3 13 3 13 2 3 3 0 9 2
15 13 7 9 2 16 9 3 13 9 2 3 15 9 13 2
15 0 9 3 0 0 9 13 9 2 16 13 1 0 9 2
17 10 9 7 13 1 15 2 16 9 13 0 9 1 10 0 9 2
29 10 9 13 13 3 1 10 0 9 2 1 15 15 13 1 10 9 3 13 2 7 1 15 4 3 10 9 13 2
11 3 13 0 0 9 2 13 15 3 13 2
9 13 15 3 10 0 9 0 9 2
21 9 1 9 2 1 9 2 1 9 9 2 1 0 9 2 7 3 1 0 9 2
9 0 9 1 10 9 13 0 9 2
11 9 1 15 15 13 14 15 0 1 0 2
16 9 1 9 2 1 10 9 15 13 9 13 15 1 10 9 2
20 1 9 2 3 13 15 3 13 9 9 2 7 7 0 9 2 9 2 3 2
12 9 1 9 2 15 13 3 13 9 0 9 2
25 1 10 9 9 2 3 15 9 13 16 9 2 13 9 1 9 7 0 9 14 9 10 9 13 2
20 7 16 13 3 0 9 3 0 2 1 15 0 13 0 9 16 0 0 9 2
7 7 15 1 15 13 3 2
22 15 2 15 1 9 2 15 15 13 2 13 2 7 15 2 15 15 15 3 13 13 2
57 3 0 9 2 0 9 2 1 15 15 13 9 1 9 1 0 9 10 3 7 3 0 9 2 15 13 9 1 9 9 7 9 9 7 10 0 9 13 9 15 1 9 2 16 13 2 1 0 9 9 2 2 3 1 0 9 2
4 13 2 13 2
10 16 15 2 15 3 13 1 9 9 2
24 9 15 13 2 13 9 9 2 0 9 2 16 4 15 1 9 13 13 15 0 2 7 13 2
11 1 9 15 0 9 3 13 1 10 9 2
15 1 15 10 0 9 7 9 2 1 15 4 13 1 0 2
12 9 15 13 1 9 7 1 0 9 3 13 2
7 9 1 11 2 9 7 9
36 16 0 9 9 9 9 11 11 2 13 13 2 16 13 9 0 9 0 9 1 11 2 0 9 1 2 2 2 2 11 12 2 12 2 2 2
16 3 15 13 13 0 9 2 7 3 13 13 9 1 0 9 2
25 13 4 3 1 9 12 2 12 9 9 9 0 9 1 11 2 7 15 16 9 1 0 0 9 2
12 13 15 0 3 0 9 1 0 9 1 0 2
27 4 13 1 12 1 12 9 1 9 0 9 2 16 13 0 2 16 4 15 1 12 9 13 9 1 9 2
25 15 4 13 0 7 0 9 2 1 15 4 13 9 2 15 15 3 13 3 3 13 1 0 9 2
12 14 2 0 2 7 1 11 4 13 0 9 2
27 0 13 1 9 13 9 7 13 1 0 9 9 2 3 0 1 9 9 2 9 2 1 9 7 9 2 2
27 13 3 0 0 9 2 13 15 1 0 9 2 3 15 3 2 13 9 1 9 2 3 15 13 9 9 2
12 13 9 13 2 16 9 4 13 1 9 9 2
7 1 9 9 13 0 9 2
6 3 9 15 13 3 2
29 13 1 9 0 9 1 9 1 9 2 1 9 1 9 7 16 9 1 9 3 2 3 1 0 9 12 9 0 2
10 13 15 3 0 9 0 2 0 9 2
11 0 10 9 13 0 9 7 13 0 9 2
8 3 15 13 1 9 9 9 2
24 16 11 11 2 3 13 9 7 3 15 13 9 2 13 3 0 2 16 4 9 7 9 13 2
33 7 13 3 11 11 2 2 15 1 9 13 2 16 4 1 9 13 2 16 13 0 9 2 7 13 15 3 1 2 0 11 2 2
11 1 9 0 7 0 9 13 9 0 9 2
17 3 7 13 1 9 0 9 2 9 2 9 2 0 9 7 9 2
15 1 11 13 0 7 0 9 13 0 9 1 0 0 9 2
26 1 12 9 10 9 15 11 13 9 1 9 2 13 14 13 1 9 7 13 15 2 10 0 9 13 2
12 13 4 1 0 2 1 9 1 9 0 9 2
30 1 9 13 1 9 0 9 1 9 9 2 0 9 13 0 9 11 1 11 2 15 15 3 13 1 0 9 10 9 2
28 9 13 1 9 13 7 3 2 13 15 1 0 9 2 0 9 2 1 0 9 1 9 9 2 9 2 9 2
15 0 13 0 9 9 7 11 1 9 1 0 11 7 9 2
30 3 2 7 1 12 9 2 15 3 2 13 0 9 2 15 15 1 10 9 13 1 0 9 7 1 9 13 0 9 2
13 15 2 15 13 0 9 2 4 15 13 3 13 2
6 13 4 7 0 9 2
32 16 9 13 12 9 2 13 15 2 16 1 0 9 15 13 1 0 9 2 7 13 15 2 3 16 0 2 15 1 11 13 2
8 14 2 9 13 9 3 0 2
30 1 11 15 9 9 13 2 16 4 15 0 9 13 1 9 3 0 7 3 0 2 16 4 13 13 1 10 0 9 2
25 15 15 13 9 9 0 2 7 3 13 1 9 0 1 9 2 16 13 1 9 0 9 1 11 2
18 15 13 0 9 1 9 2 7 7 13 9 9 1 9 1 9 13 2
5 0 9 1 0 9
36 1 0 0 9 15 1 3 0 0 9 2 0 0 9 0 1 9 2 13 1 0 0 9 0 9 3 16 0 0 9 2 11 11 2 2 2
10 1 0 0 9 9 11 13 9 0 2
36 3 4 1 9 1 11 13 3 3 2 0 0 9 2 0 1 10 0 9 2 13 0 13 1 11 9 16 14 0 2 3 9 1 0 9 2
17 9 11 4 3 13 12 2 16 4 1 9 13 2 0 9 2 2
18 3 9 11 4 14 1 9 13 9 11 13 0 9 1 11 13 9 2
15 13 4 1 15 7 13 15 2 15 13 3 9 0 9 2
22 16 10 9 13 11 2 13 4 15 13 3 9 2 15 13 9 13 9 0 0 9 2
10 4 3 13 9 2 7 15 13 9 2
13 3 9 9 13 15 1 10 9 1 9 15 0 2
55 16 13 1 9 7 0 0 9 1 0 9 2 0 9 2 9 2 9 2 7 7 15 0 9 1 9 7 1 9 9 2 13 3 13 0 9 9 2 1 11 15 13 9 2 2 15 15 1 9 3 7 3 3 13 2
39 9 13 3 15 9 9 2 15 2 13 2 3 15 2 15 1 9 9 9 7 10 9 9 13 1 10 9 7 4 13 3 0 9 13 9 0 10 9 2
28 3 0 13 10 9 1 0 9 0 9 2 10 0 9 13 13 2 3 1 9 0 9 7 0 9 1 9 2
18 1 9 3 7 3 0 9 10 9 13 1 0 9 9 9 3 0 2
15 9 9 9 9 15 3 3 13 2 3 7 1 0 9 2
32 0 13 9 2 15 13 9 9 1 0 9 1 9 13 10 9 2 1 9 15 3 13 13 7 13 15 13 9 1 0 9 2
13 3 0 2 9 13 9 7 3 9 7 9 9 2
32 16 13 15 1 10 9 1 9 2 13 3 2 16 15 1 9 1 10 9 13 1 0 9 9 3 9 7 9 1 9 9 2
5 9 15 3 13 2
23 9 7 1 9 9 13 3 1 9 2 16 4 15 13 13 0 9 7 9 1 9 13 2
45 1 10 0 9 1 9 0 9 1 9 7 1 10 9 15 3 9 9 13 7 3 1 9 13 1 9 10 9 0 9 2 16 4 13 1 9 0 9 2 15 15 10 9 13 2
28 9 10 0 9 2 15 13 3 1 9 9 0 9 7 0 9 4 3 13 2 4 15 13 1 0 9 11 2
16 1 3 0 0 9 13 9 0 2 7 14 1 9 9 9 2
10 3 16 1 15 13 9 1 9 9 2
11 0 13 7 9 9 9 1 9 0 9 2
40 16 13 1 0 9 3 9 2 3 7 1 12 9 2 3 2 13 15 1 9 1 0 9 0 9 2 15 3 0 9 13 2 7 14 1 9 7 1 9 2
36 10 9 0 9 1 9 2 1 15 13 15 1 9 9 3 3 2 4 3 13 1 0 9 2 7 2 1 0 9 9 7 9 1 9 9 2
35 13 15 2 16 15 13 0 9 1 9 7 0 9 1 0 9 2 7 13 3 9 2 16 15 15 13 2 7 13 12 1 0 9 9 2
4 9 9 13 9
13 9 0 0 9 4 13 3 13 9 1 9 12 9
27 0 0 9 2 15 13 3 0 9 1 9 9 2 13 3 1 9 14 12 9 9 0 9 12 9 9 2
14 9 9 13 1 9 9 1 9 14 12 9 1 9 2
29 1 11 11 1 0 0 9 1 0 9 1 15 1 0 9 13 9 9 9 9 0 2 11 1 0 9 1 11 2
29 9 3 13 0 9 0 9 0 9 7 13 1 9 9 0 9 1 9 11 2 15 4 13 4 13 9 0 9 2
34 1 0 9 1 0 9 4 2 1 0 9 1 9 9 2 13 9 9 9 2 12 1 0 9 1 11 1 0 9 0 11 2 11 2
20 9 2 15 10 9 13 2 13 1 11 2 11 14 3 0 2 7 7 0 2
14 1 15 15 3 13 13 1 15 0 9 0 0 9 2
31 0 0 9 15 7 3 13 13 3 1 9 3 0 9 7 0 9 2 16 13 3 9 9 0 9 2 11 3 0 9 2
18 1 14 12 9 2 15 9 1 9 3 13 2 13 9 15 0 9 2
40 11 3 13 9 0 9 2 16 13 9 2 9 2 9 2 9 7 0 9 2 15 15 0 9 13 1 9 0 9 1 9 0 9 11 2 13 11 2 11 2
27 0 9 9 13 0 12 9 9 2 16 0 0 9 13 3 9 1 9 11 7 0 9 2 11 11 11 2
21 1 0 9 13 11 11 2 1 12 9 1 15 3 13 0 7 0 9 7 11 2
24 1 0 9 0 9 4 9 10 9 13 1 12 9 7 1 9 13 9 9 1 12 9 0 2
2 0 9
2 9 2
27 9 11 11 9 9 13 9 0 9 7 13 1 15 2 15 13 1 10 9 7 10 9 0 9 13 0 2
30 0 9 15 13 1 9 12 7 1 0 9 1 0 9 9 3 13 1 0 9 9 2 0 9 13 1 9 0 9 2
12 9 9 9 15 13 13 10 9 1 9 9 2
17 13 15 1 9 11 11 7 1 0 9 9 1 15 13 2 13 2
24 9 9 9 3 13 0 0 9 2 0 9 11 7 11 2 15 15 3 10 9 13 7 13 2
18 7 0 9 13 9 1 9 0 9 3 3 3 0 7 0 0 9 2
30 0 9 9 7 9 0 15 1 9 1 0 9 2 1 9 0 9 7 0 9 2 13 9 0 9 1 9 7 9 2
15 13 3 0 9 2 15 13 0 9 2 3 13 1 9 2
23 0 9 9 13 0 9 2 3 1 9 13 13 2 16 7 0 9 11 4 1 9 13 2
29 0 9 10 9 13 7 3 0 9 1 0 9 9 2 11 2 2 9 1 9 2 2 13 3 1 0 9 2 2
55 0 9 11 11 4 13 9 9 7 1 9 2 3 15 0 9 3 13 1 9 2 9 3 13 9 0 9 7 9 2 15 7 13 0 0 9 2 3 9 2 3 11 13 11 2 7 0 9 12 9 1 0 9 2 2
17 0 9 11 11 13 0 0 9 7 0 0 9 16 9 0 9 2
14 0 9 13 3 3 2 1 10 9 13 13 3 15 2
9 9 0 9 3 13 0 9 9 2
15 0 9 13 7 0 9 0 7 0 9 2 11 11 2 2
19 1 9 0 10 0 9 2 0 3 9 9 2 13 10 0 9 11 11 2
33 11 0 1 9 11 3 13 13 10 3 0 9 0 9 1 0 7 0 9 2 7 1 0 9 16 0 9 13 13 9 10 9 2
21 0 9 11 11 13 13 0 9 2 7 16 0 9 9 15 13 1 9 0 9 2
28 11 11 2 2 9 2 11 2 7 11 11 2 0 9 11 2 13 10 0 9 1 9 0 9 7 0 9 2
15 9 2 11 2 11 11 2 11 2 9 1 15 13 13 2
5 9 12 2 9 2
4 9 16 0 9
10 9 0 9 1 9 12 11 13 0 9
28 0 9 1 9 0 9 0 9 12 11 1 0 9 1 11 1 0 9 3 0 9 4 13 12 2 9 12 2
13 9 13 12 9 2 12 13 0 7 12 0 9 2
33 1 9 13 15 1 15 2 9 0 9 2 15 13 1 9 9 1 0 9 0 9 1 11 2 3 13 2 16 15 0 9 13 2
5 13 15 0 9 2
6 11 2 12 11 2 11
21 9 13 11 13 9 9 1 12 1 12 9 2 15 1 9 9 13 7 0 9 2
8 15 7 1 0 9 4 13 2
14 7 10 0 9 15 1 3 0 9 1 0 9 13 2
16 1 9 12 13 1 10 9 0 9 0 9 0 7 0 9 2
30 9 2 0 9 0 9 2 7 13 3 1 0 9 9 1 12 2 9 7 3 1 9 9 11 11 1 12 2 9 2
38 13 2 14 2 16 9 12 11 3 14 13 9 11 7 16 15 10 9 4 3 13 1 9 11 1 9 9 2 13 15 1 9 0 9 11 13 13 2
49 0 9 15 13 13 1 0 0 9 0 9 9 2 12 1 0 9 3 2 16 4 13 3 0 9 0 9 2 9 2 9 2 12 7 0 9 9 2 12 2 1 15 13 3 13 1 0 9 2
19 9 0 9 15 13 9 9 13 1 12 7 3 9 7 3 15 3 13 2
11 0 1 15 1 15 13 9 10 0 9 2
22 9 10 9 15 1 9 13 0 9 2 9 2 9 7 10 0 3 7 3 0 9 2
18 9 10 0 9 3 13 9 0 0 9 1 9 0 9 1 9 12 2
22 9 0 9 13 1 0 9 2 7 1 15 2 16 4 15 13 1 9 0 0 9 2
27 0 9 9 1 12 11 13 3 2 14 15 13 13 0 9 2 3 3 13 13 9 3 0 9 1 9 2
15 15 0 3 13 2 16 0 0 9 3 13 0 0 9 2
22 10 0 9 10 0 9 1 9 13 1 9 9 12 11 14 10 0 9 1 0 9 2
42 13 1 15 0 7 3 14 0 9 9 2 12 1 9 11 2 11 1 0 11 2 15 0 9 3 7 3 13 0 9 2 0 7 9 2 0 9 0 1 0 9 2
25 16 4 13 11 13 1 0 9 2 3 15 15 3 13 9 11 11 2 13 4 0 9 0 9 2
15 0 9 7 13 3 1 15 2 15 3 13 1 11 13 2
7 9 0 9 12 11 9 2
15 9 9 0 9 2 11 2 12 2 9 2 12 2 9 2
2 0 9
18 9 2 9 11 11 13 2 16 10 11 13 2 9 1 12 9 2 2
21 3 3 13 0 9 2 13 0 7 3 0 9 7 13 1 10 0 2 9 2 2
12 7 3 15 13 1 0 9 2 9 0 9 2
11 9 3 0 9 9 13 11 11 2 11 2
24 9 15 13 3 1 9 10 9 2 15 13 2 16 9 12 15 13 9 14 1 9 10 9 2
12 9 4 13 13 0 9 0 9 1 0 9 2
25 11 2 11 15 1 9 9 13 0 9 2 7 3 9 3 13 2 16 3 1 0 7 0 9 2
18 1 11 15 1 9 13 3 12 9 2 7 15 0 9 9 1 9 2
32 11 11 2 12 2 13 0 9 1 0 9 2 9 0 9 13 7 13 7 1 0 9 13 0 0 9 13 3 0 0 9 2
6 3 0 2 3 0 2
19 11 11 2 12 2 13 10 0 9 1 9 2 15 3 13 1 0 9 2
7 13 15 9 7 0 9 2
10 13 15 0 9 2 9 2 0 9 2
13 0 9 13 9 1 9 16 9 0 7 0 9 2
6 9 13 0 9 9 2
11 0 9 9 3 0 0 9 13 15 0 2
8 13 14 0 9 0 0 9 2
9 9 12 2 9 11 11 2 11 2
5 9 11 2 11 2
7 12 2 2 12 2 9 2
3 0 0 9
29 0 9 9 7 0 9 11 13 13 3 9 9 11 11 2 15 15 13 1 0 9 1 11 7 13 1 0 9 2
25 1 9 0 7 0 2 9 1 9 11 11 2 11 11 7 11 11 13 3 1 9 7 11 11 2
17 3 12 9 13 1 9 1 0 0 9 7 1 15 9 13 9 2
11 0 9 15 1 0 9 13 1 9 9 2
14 16 15 0 13 13 0 9 9 2 9 7 0 9 2
34 0 0 9 16 9 9 7 0 9 15 13 3 1 15 10 9 2 15 1 9 1 9 7 9 9 13 3 0 2 2 0 2 9 2
22 0 9 3 13 0 9 0 9 2 0 9 11 2 11 2 11 11 11 7 9 9 2
11 3 13 1 9 3 0 9 14 13 9 2
39 1 9 9 13 9 13 9 2 0 9 1 11 11 2 9 0 9 0 9 1 11 11 7 11 11 2 7 0 9 0 9 0 9 1 11 7 11 11 2
25 9 1 9 11 11 13 9 0 9 1 9 0 9 7 9 15 9 9 2 0 1 9 0 9 2
14 1 9 12 13 11 11 16 0 9 1 9 0 9 2
21 1 10 9 15 13 1 2 0 9 9 2 15 1 15 13 1 9 14 9 2 2
11 9 7 0 9 13 3 1 10 9 0 2
15 1 10 9 3 0 9 9 7 10 0 9 13 1 0 2
3 9 0 9
17 9 2 0 9 11 11 13 1 0 0 9 9 9 9 1 11 2
9 10 9 4 13 1 9 0 9 2
8 9 0 9 15 13 1 15 2
20 13 15 1 9 2 9 2 11 11 2 15 13 1 0 9 1 9 0 9 2
29 13 9 11 11 11 2 9 12 2 9 9 2 2 15 3 13 1 9 9 9 7 9 7 13 0 9 0 9 2
31 1 11 11 2 9 9 9 2 9 2 12 2 12 2 13 9 2 0 2 9 2 15 1 0 9 13 1 9 0 9 2
11 0 9 13 0 9 9 9 2 9 12 2
16 0 9 3 13 0 0 9 7 13 15 1 0 9 0 9 2
11 11 11 13 1 9 0 9 1 0 9 2
14 1 9 1 10 9 13 1 0 2 7 1 0 9 2
27 7 15 13 0 13 3 1 15 2 7 3 13 1 9 16 1 10 2 0 9 2 2 15 13 7 0 2
15 13 0 13 9 0 9 2 15 15 13 1 0 0 9 2
8 13 13 0 2 0 9 9 2
18 9 0 9 13 0 2 13 2 2 16 15 1 9 13 0 0 9 2
8 15 15 15 0 0 9 13 2
15 10 9 13 2 0 2 9 2 13 3 2 1 0 9 2
16 1 9 10 0 9 13 9 2 16 4 15 13 1 0 9 2
19 13 1 9 0 9 9 2 15 1 9 13 0 0 9 1 9 0 9 2
2 11 11
4 9 9 9 2
8 12 2 0 9 9 0 9 2
10 9 0 9 2 11 2 12 2 9 2
37 9 9 7 0 9 1 0 0 9 1 11 4 3 13 1 0 9 1 9 0 9 9 11 11 11 2 9 0 7 0 9 2 0 3 1 9 2
30 9 9 13 9 0 2 0 7 0 9 1 0 7 0 9 2 15 13 1 9 0 9 2 9 9 9 7 0 9 2
8 9 13 0 1 12 2 9 2
8 11 11 16 9 1 9 0 9
2 0 11
26 9 11 11 11 1 9 15 4 13 9 3 0 0 9 1 9 11 2 11 2 11 2 9 7 9 2
19 13 15 1 12 2 1 12 2 9 1 0 9 11 1 0 9 1 11 2
20 1 12 0 9 3 13 1 9 9 7 0 9 2 3 0 9 0 0 9 2
28 9 13 3 9 11 2 9 9 2 15 13 9 9 10 9 2 7 9 2 0 0 9 1 9 7 1 9 2
8 9 9 13 0 7 0 9 2
5 1 9 3 1 9
35 9 1 9 12 2 15 9 0 9 13 1 9 0 9 0 1 9 11 9 11 11 2 13 3 1 10 9 13 15 0 9 1 9 9 2
25 1 9 9 13 13 1 9 9 2 15 4 0 9 13 0 9 7 9 9 3 0 1 10 9 2
8 2 0 9 4 13 0 9 2
21 13 4 9 12 9 12 9 1 0 9 12 9 2 15 15 4 13 16 0 9 2
13 0 9 3 13 4 2 2 13 9 9 11 11 2
26 1 11 11 2 9 0 9 2 15 9 1 9 12 13 2 13 9 9 0 9 1 9 9 10 9 2
18 2 1 0 9 2 16 15 1 9 13 2 3 13 2 2 13 11 2
25 9 1 9 12 2 15 13 9 0 9 9 9 7 15 13 11 11 2 4 1 9 0 9 13 2
18 9 1 9 11 11 13 9 1 9 12 2 15 13 9 1 0 9 2
19 15 11 11 7 9 11 11 3 9 9 13 2 7 16 1 15 3 13 2
38 9 11 1 10 9 3 13 9 0 9 2 15 1 9 9 13 1 2 0 9 0 9 2 16 4 3 13 10 9 7 13 9 1 9 13 7 13 2
15 2 1 9 0 9 13 9 0 9 2 2 13 1 9 2
10 2 9 0 9 13 0 9 0 9 2
25 4 13 9 2 15 3 1 9 12 9 1 9 0 9 13 0 9 9 2 2 13 1 15 11 2
1 3
25 0 2 0 9 9 1 9 2 15 13 0 0 9 11 11 2 13 3 1 10 9 1 0 9 2
12 0 9 9 15 13 12 2 9 1 9 11 2
39 0 7 0 9 1 11 7 0 0 9 13 1 10 9 0 9 0 9 0 2 15 1 0 9 13 0 9 15 9 7 9 1 9 0 9 1 9 12 2
7 9 1 9 7 1 9 9
22 0 9 9 0 9 13 9 0 7 0 9 1 0 9 12 1 0 9 1 10 9 2
14 13 1 15 3 9 0 9 7 3 7 3 0 9 2
19 1 15 0 14 13 7 9 0 9 11 11 2 12 2 2 0 9 9 2
16 9 3 13 0 0 2 0 9 2 15 13 7 0 9 9 2
39 13 2 14 15 0 9 1 0 9 11 1 9 7 9 0 9 0 9 2 13 13 2 16 0 9 13 0 2 3 0 1 9 9 2 16 15 13 11 2
26 0 13 3 9 1 9 1 0 9 2 15 13 11 11 9 12 2 3 14 1 9 12 1 9 9 2
51 16 4 15 11 13 15 1 9 0 9 1 11 2 13 4 2 16 10 9 2 9 11 12 2 11 12 2 11 2 13 0 9 16 10 9 2 13 15 7 1 9 13 1 9 0 9 1 0 0 9 2
19 1 0 9 4 3 13 9 11 14 1 9 9 9 7 15 13 3 3 2
27 13 2 1 10 9 13 9 9 2 16 1 9 9 1 9 2 15 13 3 3 9 2 13 11 1 11 2
29 16 13 3 0 2 9 2 15 11 12 2 13 2 4 13 1 9 0 9 1 0 9 7 1 0 9 0 9 2
33 1 0 9 0 0 9 4 15 11 13 2 16 0 9 13 0 9 0 2 7 10 0 0 2 2 9 0 2 9 2 9 2 2
36 9 11 11 1 9 0 9 1 0 9 4 1 9 3 13 7 1 0 9 15 13 2 16 9 13 9 11 2 3 11 2 16 15 3 13 2
31 1 9 9 11 13 2 16 11 12 2 7 10 9 13 13 3 1 0 2 0 2 9 0 0 9 2 7 1 9 3 2
32 3 15 9 13 1 15 2 16 9 13 0 9 2 10 9 7 1 0 2 11 13 2 13 1 0 9 2 15 13 9 9 2
20 3 3 7 11 13 0 9 11 11 2 15 13 1 9 11 11 7 11 11 2
20 1 9 12 4 3 1 10 9 13 3 0 9 2 3 9 0 7 0 2 2
32 9 1 9 2 0 2 11 11 2 9 1 9 0 1 11 11 2 2 2 2 2 0 14 1 9 9 1 11 2 13 0 2
42 1 9 4 1 11 12 2 9 12 13 9 9 0 9 11 11 7 11 0 9 4 2 3 3 2 3 3 2 16 15 13 1 10 9 2 13 1 11 3 9 12 2
40 1 0 9 11 3 13 9 1 12 9 1 9 9 0 2 15 13 0 9 1 0 9 2 1 9 15 13 9 1 9 2 3 0 1 9 0 9 1 11 2
21 0 13 7 0 9 9 1 0 9 2 13 9 2 3 9 1 9 10 9 13 2
23 16 13 3 11 11 1 9 2 9 11 11 4 13 9 12 1 9 2 7 1 0 9 2
33 9 11 11 1 11 4 3 13 1 9 0 9 7 1 9 1 0 2 11 11 3 1 9 9 2 7 12 2 9 12 1 11 2
14 9 13 3 13 0 9 9 2 7 3 13 0 9 2
26 0 2 11 13 13 1 9 0 2 11 2 3 1 9 2 1 9 0 2 11 13 3 9 9 2 2
22 1 0 9 13 13 13 0 0 9 2 3 9 0 2 16 11 11 13 3 0 9 2
10 3 13 13 11 11 2 13 12 2 9
3 1 0 9
12 11 11 2 11 11 2 16 13 0 9 9 2
21 0 0 9 7 0 9 2 15 13 9 1 0 9 2 13 1 9 9 0 9 2
7 3 0 9 13 9 11 2
6 11 11 2 9 9 2
41 0 0 0 9 0 9 2 12 2 12 2 2 1 15 15 1 0 9 11 7 11 13 3 9 11 11 2 11 7 9 1 11 2 13 3 9 0 10 0 9 2
21 1 9 11 11 7 1 9 11 11 10 0 0 9 13 1 10 0 9 0 9 2
5 11 11 2 9 2
23 0 9 0 2 12 2 12 2 0 3 9 9 1 0 9 13 9 9 1 9 0 9 2
17 9 0 0 9 9 11 12 2 1 0 9 2 15 13 12 0 9
3 9 9 9
26 9 0 0 9 9 11 1 11 2 15 13 3 0 9 0 0 9 2 13 1 0 0 9 9 0 2
23 0 9 1 0 9 1 9 11 13 13 9 12 2 13 2 14 0 0 9 1 9 12 2
25 9 3 13 9 11 11 9 0 2 15 1 9 9 9 1 9 1 9 0 9 13 0 9 11 2
33 3 1 10 9 9 0 9 0 9 4 0 9 13 1 0 9 11 2 3 1 9 9 2 9 11 2 7 10 9 2 9 11 2
15 15 13 1 10 9 3 13 2 9 0 13 9 9 2 2
27 9 1 0 9 7 3 13 9 1 0 9 11 11 12 2 2 10 2 9 2 0 9 13 9 9 9 2
19 9 13 7 9 0 9 2 10 9 7 0 9 0 9 1 9 10 9 2
26 1 9 9 0 9 15 9 13 3 1 9 0 9 2 7 16 4 13 0 3 9 1 9 0 9 2
28 13 15 15 7 9 9 2 3 3 9 9 9 0 1 0 9 2 12 2 11 2 11 13 9 0 7 0 2
20 1 0 9 13 9 0 9 2 0 9 11 2 11 1 9 9 2 14 13 2
18 9 9 13 7 9 2 15 11 13 9 9 1 0 9 9 0 9 2
18 1 9 2 1 15 15 10 9 13 2 15 9 13 10 0 0 9 2
11 3 9 9 0 13 13 3 1 0 9 2
27 9 11 11 12 2 15 13 11 2 7 14 11 2 7 3 15 13 9 1 11 2 16 15 1 15 13 2
8 11 11 13 11 2 7 11 2
16 9 11 13 7 0 9 2 9 1 10 9 13 13 16 9 2
19 1 10 9 13 9 9 9 9 0 9 2 15 13 9 0 7 0 9 2
10 13 13 2 16 0 9 4 3 13 2
5 0 9 1 0 9
34 9 9 9 1 0 9 1 9 13 0 9 0 9 9 7 9 9 10 9 1 10 9 1 9 2 15 13 1 10 9 3 0 9 2
31 9 9 2 0 1 9 0 0 9 9 9 1 11 2 13 11 2 11 2 11 2 11 2 11 2 11 7 11 2 11 2
44 9 3 13 0 9 1 9 9 1 11 7 1 11 2 13 10 0 9 2 0 2 11 1 11 2 2 13 0 9 1 0 9 7 10 0 9 7 13 0 9 1 0 9 2
25 3 13 9 0 9 0 9 2 11 2 11 2 11 2 11 2 7 10 9 2 11 2 11 2 2
24 13 13 3 9 9 0 9 0 9 11 13 2 15 15 9 0 9 13 3 3 16 9 9 2
23 13 0 9 2 1 15 10 9 1 9 0 9 13 1 0 9 13 3 0 9 0 9 2
16 9 13 13 0 9 7 9 0 9 2 0 0 9 0 9 2
7 9 13 0 9 1 9 2
27 9 9 13 1 9 12 2 3 9 9 13 1 0 9 1 11 1 11 2 15 15 3 13 0 9 9 2
36 9 12 3 1 9 0 12 9 13 0 9 11 2 15 15 1 3 0 9 1 11 2 1 15 9 1 0 9 13 2 4 13 11 1 11 2
35 10 0 9 13 0 9 14 0 9 2 7 0 0 9 2 15 3 4 13 9 0 2 9 2 10 9 1 0 0 9 13 13 3 13 2
36 1 0 9 0 9 13 2 16 13 10 9 2 9 0 9 2 9 9 9 9 7 0 9 3 0 11 2 3 9 2 9 2 7 0 9 2
23 1 10 9 13 1 0 11 10 9 9 0 9 2 0 1 10 0 9 0 9 1 0 2
23 1 15 13 3 0 0 9 2 0 9 0 9 7 9 0 9 9 10 2 0 2 9 2
17 7 3 0 0 9 2 0 15 1 0 9 15 0 9 9 11 2
13 0 13 9 1 0 9 7 0 0 9 0 9 2
25 0 13 9 0 15 14 1 0 9 9 2 7 3 1 0 9 0 15 9 0 9 7 10 9 2
19 1 9 9 0 9 15 13 3 0 0 9 0 9 2 15 15 13 9 2
41 1 11 7 1 11 13 0 9 0 9 1 9 0 0 9 2 3 0 1 9 2 9 2 2 16 15 3 13 3 9 0 0 9 16 9 1 9 0 9 9 2
86 0 2 3 2 0 2 0 9 7 0 9 1 15 13 14 1 9 0 7 1 9 0 9 2 3 15 0 9 13 3 1 9 0 9 9 2 15 13 0 9 7 0 9 9 1 0 11 2 0 0 9 0 9 9 1 0 9 2 1 0 9 0 9 1 11 2 3 0 11 1 9 0 9 2 7 0 9 1 0 9 3 0 9 0 9 2
15 15 10 9 13 1 0 0 9 0 9 1 0 0 9 2
27 1 15 0 12 1 15 13 3 3 3 3 0 9 1 0 11 2 0 3 1 9 11 1 11 9 10 9
10 11 2 15 1 15 1 12 9 13 2
9 13 9 1 9 7 13 0 3 2
8 15 1 9 15 2 1 9 2
6 0 0 9 13 1 9
10 3 0 0 9 15 13 1 9 0 9
8 3 3 13 9 12 9 12 9
10 3 1 9 11 15 13 9 0 9 2
31 13 1 0 9 13 9 2 1 15 15 13 11 11 2 11 11 2 1 9 11 11 2 0 9 7 9 3 14 0 9 2
19 6 2 3 2 3 2 13 0 9 2 10 0 9 13 9 9 1 9 2
18 0 9 1 0 9 2 9 2 15 3 13 1 0 9 9 0 9 2
21 9 15 3 13 9 2 7 9 9 13 1 11 1 9 1 10 9 1 0 9 2
21 16 15 13 0 2 7 0 9 1 9 0 9 9 2 10 9 13 0 9 9 2
15 3 13 0 9 7 9 7 3 13 1 9 9 0 9 2
9 9 2 3 9 2 13 1 9 2
13 3 16 0 1 9 2 15 9 13 9 1 9 2
17 13 15 9 12 7 1 0 9 2 0 11 13 10 9 9 9 2
6 15 11 7 12 11 2
9 1 9 15 13 12 9 9 9 2
17 6 2 3 2 3 2 13 0 9 2 10 0 9 13 9 9 2
28 1 9 0 9 2 15 13 3 9 7 13 15 1 10 9 2 13 9 7 13 1 0 9 1 9 7 9 2
11 3 0 2 3 0 2 3 13 0 9 2
16 13 3 9 9 2 7 10 9 11 7 11 4 13 3 9 2
4 15 13 0 2
42 0 9 2 11 7 11 2 0 9 2 9 11 9 2 9 9 2 1 9 15 13 14 12 2 2 11 0 9 2 13 3 9 7 13 14 0 9 2 7 0 9 2
18 13 15 9 12 7 1 11 2 0 0 9 13 10 9 9 12 9 2
6 15 11 2 12 11 2
8 1 9 15 13 7 12 9 2
18 9 1 9 0 9 13 12 1 0 9 2 15 13 1 9 12 9 2
12 13 15 1 12 9 0 11 3 1 9 12 2
7 9 1 9 13 7 0 2
21 9 13 1 0 9 9 13 1 0 9 2 16 10 9 13 9 3 0 16 9 2
22 9 7 9 13 9 13 0 9 11 11 1 9 2 16 4 4 13 9 0 0 9 2
10 1 11 13 0 9 3 1 9 12 2
29 1 9 13 7 13 9 7 9 9 13 9 15 9 9 3 0 1 0 11 2 12 9 1 9 2 13 3 13 2
8 4 13 9 9 2 13 9 2
10 4 13 0 0 9 7 3 0 9 2
11 1 9 0 9 13 9 9 1 0 9 2
28 10 9 1 9 2 2 10 0 9 2 15 13 10 9 2 15 13 0 9 2 0 9 2 2 13 9 9 2
19 9 13 1 9 0 9 9 7 3 15 9 13 9 0 9 2 0 9 2
28 9 3 0 2 0 9 2 16 0 9 13 1 0 9 9 2 13 9 1 9 2 3 15 0 1 0 9 2
24 0 1 15 7 3 13 2 15 13 9 1 0 9 2 15 3 7 13 2 3 10 9 13 2
28 9 3 13 0 9 9 7 13 15 7 13 2 16 15 3 13 1 3 0 9 9 2 1 15 15 3 13 2
20 9 1 0 9 13 13 13 1 9 9 1 0 0 9 7 13 0 9 9 2
12 13 3 9 2 16 13 0 15 13 0 9 2
25 9 9 12 9 12 9 2 15 1 9 13 0 9 1 0 0 11 2 13 15 2 14 3 13 2
41 9 3 13 15 3 13 0 9 9 10 9 7 9 2 0 9 2 1 9 7 9 2 12 9 9 13 1 9 2 7 9 1 9 9 2 10 9 7 9 3 2
18 13 3 0 0 9 0 9 2 15 13 9 1 10 9 7 9 0 2
2 9 3
16 0 2 0 9 0 9 0 9 13 14 1 9 1 10 9 2
15 1 0 9 13 0 9 9 0 2 3 0 9 7 9 2
11 1 0 9 13 9 0 9 1 0 9 2
26 0 9 7 0 9 9 13 9 9 3 2 16 1 9 10 9 9 2 0 0 9 2 13 1 9 2
9 9 1 15 7 13 9 0 9 2
16 0 15 0 9 1 9 10 9 2 13 13 1 0 9 9 2
12 1 9 13 0 0 0 9 1 9 7 9 2
15 13 1 9 7 9 7 9 9 10 9 2 11 0 9 2
24 13 9 1 9 7 9 2 3 15 3 13 7 13 0 0 9 11 11 1 10 9 1 11 2
14 1 9 13 9 0 0 9 7 9 2 15 9 13 2
7 11 3 1 0 9 13 2
28 1 10 9 0 1 0 9 15 13 2 16 1 0 9 13 11 11 2 9 0 9 11 11 7 9 11 11 2
18 0 9 13 1 9 12 9 9 7 0 9 0 9 2 9 7 9 2
10 0 9 3 4 1 9 12 9 13 2
16 9 13 13 1 9 15 2 15 15 1 0 9 13 7 13 2
13 0 9 15 1 9 13 1 0 9 2 15 0 2
11 0 9 15 3 13 14 1 9 0 9 2
10 1 9 9 9 1 11 4 13 9 2
19 9 0 2 11 13 3 1 0 9 13 1 9 7 0 9 13 1 11 2
18 0 9 9 13 9 12 12 9 7 9 2 0 1 9 1 9 0 2
9 0 9 9 13 9 1 0 9 2
16 9 9 1 9 15 13 14 3 2 16 9 0 9 1 9 2
15 3 15 3 0 0 9 13 1 9 0 9 7 0 9 2
26 13 15 9 2 15 13 0 14 1 9 9 2 15 15 3 13 2 15 1 15 13 2 13 10 9 2
8 9 0 9 9 7 0 9 2
19 9 0 9 2 1 9 7 1 9 13 0 9 9 9 1 0 0 9 2
13 9 1 0 0 11 13 13 0 9 10 9 9 2
11 1 3 0 9 13 1 9 9 0 9 2
21 13 7 0 9 7 0 9 2 16 9 1 0 9 0 9 11 13 13 12 9 2
9 15 15 13 1 9 2 10 9 2
24 1 9 1 0 7 0 9 2 3 13 0 9 13 1 9 2 13 0 9 1 0 0 9 2
5 13 9 7 9 2
60 9 1 9 0 3 0 9 2 0 1 9 3 0 9 7 1 9 7 9 9 13 9 1 0 9 1 9 0 9 2 3 1 9 11 2 1 0 9 0 0 9 7 0 9 1 9 2 1 9 0 1 15 9 9 2 3 0 0 9 2
15 0 9 13 3 3 13 16 14 9 0 9 2 0 9 2
9 9 3 13 1 9 9 0 9 2
30 9 9 7 9 9 9 7 9 15 7 13 2 16 4 9 9 12 9 12 9 4 13 9 1 9 9 1 0 9 2
21 9 7 9 1 9 4 3 13 2 13 9 1 10 9 1 9 2 9 7 9 2
26 1 10 0 9 9 9 3 13 9 7 9 2 16 4 0 7 0 0 9 13 7 13 9 0 9 2
1 9
7 9 9 13 0 0 9 2
17 1 9 0 9 2 9 7 9 0 9 2 0 1 0 0 9 2
11 11 11 2 0 9 2 13 1 0 9 2
17 0 9 2 12 12 9 0 0 9 2 3 13 9 9 1 9 2
5 13 14 9 0 2
12 9 11 13 9 12 7 12 9 1 9 9 2
9 9 13 1 9 9 1 0 9 2
11 1 9 13 9 0 12 9 1 0 9 2
15 0 9 15 9 7 9 13 1 3 0 9 3 0 9 2
8 0 9 1 15 3 15 13 2
14 9 3 13 1 11 2 7 3 9 13 1 9 9 2
17 2 1 9 7 0 9 15 13 13 9 2 2 13 9 11 9 2
4 2 13 13 2
7 13 0 9 1 0 9 2
9 10 9 13 7 1 10 9 2 2
11 9 13 0 9 7 13 13 9 0 9 2
27 13 13 1 0 0 9 0 9 2 1 9 13 3 13 0 9 2 7 13 0 9 0 0 9 0 9 2
22 0 9 2 15 13 3 0 9 0 9 2 15 4 13 1 9 3 0 0 9 9 2
8 3 3 13 0 9 12 9 2
14 9 13 1 9 0 9 13 3 0 12 7 9 9 2
18 0 9 2 15 13 9 7 13 1 9 2 13 1 0 9 3 0 2
21 13 0 2 16 0 9 15 1 9 13 1 0 9 2 15 13 0 0 11 11 2
12 15 1 0 9 3 13 9 1 9 2 9 2
11 1 0 9 13 9 13 0 0 0 9 2
6 1 9 0 7 0 2
12 13 15 3 9 2 0 10 9 1 0 9 2
5 0 9 9 13 2
16 1 9 9 2 0 3 16 11 2 4 3 9 13 3 0 2
7 0 9 9 15 3 13 2
7 0 9 13 10 0 9 2
15 1 0 9 15 3 3 13 0 9 0 0 2 0 9 2
5 0 9 0 9 2
24 9 7 9 13 15 2 1 15 15 9 3 13 2 3 13 2 15 15 15 13 16 0 9 2
8 16 9 4 3 13 4 13 2
2 9 9
39 9 2 9 9 13 2 13 11 11 2 11 10 9 1 9 0 9 11 11 2 0 9 1 9 1 9 2 9 0 9 2 11 12 2 12 2 12 2 2
25 9 13 3 2 7 13 1 0 0 9 15 1 10 9 1 15 13 7 3 14 3 3 1 9 2
68 3 0 9 10 0 9 13 3 13 1 9 7 9 2 13 4 3 7 1 9 2 13 15 2 16 1 9 0 9 0 9 15 3 3 1 0 9 13 9 2 7 0 9 2 3 10 0 9 2 13 7 0 1 0 9 13 3 2 16 15 1 15 1 9 13 0 9 2
56 1 11 2 11 2 11 15 11 11 0 9 2 13 14 3 1 0 9 2 2 14 3 2 3 2 2 10 9 15 13 2 14 0 9 1 0 9 2 7 2 4 3 1 15 13 13 10 3 0 9 2 2 9 0 2 2
26 13 3 3 0 9 2 15 1 9 0 13 2 9 2 7 15 0 9 2 7 13 15 3 1 9 2
42 16 4 1 9 1 9 2 1 15 13 9 2 13 7 13 15 9 0 2 0 9 1 11 11 2 13 13 2 16 7 12 1 0 0 9 9 11 15 13 1 9 2
19 0 9 15 13 3 3 7 2 16 9 0 13 4 13 1 9 0 9 2
32 1 9 2 0 9 2 2 7 1 2 9 2 13 13 1 9 11 11 2 14 1 9 9 3 0 7 0 2 3 7 9 2
21 16 15 9 11 1 0 0 9 13 2 13 15 0 2 3 9 1 10 9 13 2
97 16 13 9 2 16 3 1 0 9 2 13 15 2 16 13 13 3 14 1 0 9 9 11 2 11 1 0 11 2 9 1 0 11 2 12 2 12 2 2 15 4 15 7 3 2 12 2 12 2 13 16 0 9 0 0 9 13 1 0 9 15 2 16 4 13 0 9 1 9 0 9 1 9 1 9 7 1 0 9 1 15 2 1 10 10 9 15 13 13 7 0 9 1 9 9 11 2
11 1 0 3 0 9 13 3 0 12 9 2
46 3 9 9 11 13 0 9 1 9 2 1 10 0 7 0 9 13 2 16 15 13 1 10 9 3 15 13 2 7 15 7 1 9 2 3 15 15 13 13 9 2 3 3 7 9 2
25 3 3 16 0 13 2 16 0 7 0 9 1 9 13 0 9 2 7 0 9 0 7 0 9 2
57 11 11 1 9 9 0 9 2 2 11 12 2 12 2 2 13 1 0 2 16 0 9 1 11 2 11 2 13 1 0 9 1 0 9 1 10 0 9 1 10 9 2 0 9 2 13 2 14 7 1 9 10 3 0 9 2 2
24 9 9 15 1 9 13 13 2 3 16 16 0 9 0 9 2 16 4 0 9 13 3 2 2
37 2 3 2 2 13 11 2 2 16 9 11 13 1 15 2 16 9 1 9 1 0 9 2 3 3 0 0 9 2 15 1 10 9 3 13 2 2
29 13 0 0 9 10 0 0 9 2 9 1 9 3 13 1 0 9 1 10 9 2 15 3 13 13 1 9 2 2
20 13 3 3 0 9 13 7 13 0 9 7 1 9 2 16 15 15 13 13 2
23 0 9 13 2 13 3 3 1 9 0 0 11 1 0 0 11 2 16 15 13 9 11 2
11 9 2 16 3 15 13 2 13 3 0 2
15 7 13 10 0 9 2 13 4 11 1 12 9 7 13 2
22 1 10 9 3 13 2 13 7 13 0 0 9 14 0 7 0 9 2 7 3 9 2
24 1 9 9 0 9 9 2 15 9 13 2 13 1 9 10 9 0 9 7 0 9 9 11 2
27 1 0 9 13 9 7 15 2 16 13 11 2 13 4 3 1 10 9 9 15 13 7 1 15 15 13 2
24 13 15 14 2 16 4 1 9 0 2 11 1 9 0 9 9 12 13 9 2 7 0 9 2
34 7 16 4 0 9 13 1 0 0 9 0 0 9 0 2 9 2 7 2 16 15 13 1 9 2 0 0 9 1 11 7 0 9 2
23 16 13 1 0 9 2 13 15 1 11 3 1 9 12 1 9 1 9 9 1 9 11 2
12 3 2 1 0 9 3 13 7 0 0 9 2
24 1 9 13 9 0 9 1 0 2 0 7 0 2 3 0 2 9 9 2 16 4 9 13 2
42 1 10 9 13 13 0 9 11 2 0 9 7 0 9 11 11 2 15 1 9 13 7 1 0 9 13 10 9 2 15 4 3 13 9 7 13 4 15 9 1 9 2
30 13 7 12 9 1 9 9 7 13 0 9 2 3 1 0 9 0 9 1 15 2 15 13 13 1 9 2 9 13 2
14 13 2 10 0 9 4 13 1 9 7 13 1 9 2
18 0 9 2 3 13 4 9 3 3 13 1 9 2 13 0 0 9 2
23 13 3 7 3 13 9 11 2 11 13 1 11 0 9 2 10 0 2 7 3 0 9 2
18 0 9 9 9 7 10 9 1 12 7 9 1 0 9 3 13 15 2
18 9 13 1 9 0 9 1 9 7 9 3 10 9 0 3 0 9 2
26 3 7 13 2 7 3 14 3 2 9 0 9 2 15 4 1 0 9 13 9 2 3 3 0 9 2
14 0 0 9 13 2 16 15 11 13 13 2 1 9 2
9 9 13 3 0 9 0 0 9 2
38 15 13 9 1 0 0 9 2 3 3 9 9 13 7 13 1 15 0 9 2 1 0 9 15 7 3 13 9 2 15 13 14 1 9 9 1 9 2
15 0 9 15 13 3 14 10 0 2 7 16 3 0 9 2
22 0 9 15 3 3 13 9 10 9 2 16 13 0 11 2 0 11 2 0 9 9 2
13 7 0 9 0 9 3 13 1 0 9 10 9 2
24 3 0 13 2 16 10 3 0 9 10 9 12 2 9 4 1 9 1 9 13 0 0 9 2
12 0 0 9 4 13 0 9 9 7 9 9 2
14 9 10 0 9 4 13 9 7 9 2 0 7 0 2
35 15 13 0 9 2 3 15 11 13 9 9 1 10 0 9 2 15 13 1 0 0 0 9 7 3 13 0 7 0 9 13 1 0 9 2
26 1 15 2 16 9 11 7 9 13 0 7 16 0 0 9 9 1 11 3 13 2 13 3 0 9 2
13 11 13 3 0 9 1 9 0 2 0 7 0 2
11 3 13 1 9 0 7 0 9 1 11 2
19 1 3 0 13 13 9 1 9 0 1 9 0 0 9 9 1 0 11 2
8 0 9 13 3 13 0 9 2
13 3 15 13 0 9 2 16 3 13 11 2 11 2
26 9 9 7 11 13 0 2 3 1 9 1 9 0 9 2 15 9 15 13 3 13 1 0 9 9 2
24 0 9 3 13 13 3 9 11 2 9 9 2 3 13 2 14 10 9 3 0 11 2 11 2
29 13 9 1 10 9 1 10 9 0 2 0 7 3 0 9 4 13 14 0 2 7 3 0 2 3 1 9 15 2
18 13 3 0 13 2 16 15 9 11 4 15 1 3 0 9 3 13 2
29 2 11 11 7 11 11 13 1 0 9 1 11 2 11 11 13 1 9 1 9 9 11 11 7 1 0 9 11 2
7 0 9 7 9 13 1 15
3 3 0 9
3 1 9 9
28 9 11 2 9 9 2 3 0 14 9 2 15 3 2 0 9 13 2 11 12 2 12 2 2 13 1 9 2
52 0 9 2 2 15 15 3 13 1 9 2 2 15 3 13 7 4 13 1 0 9 2 2 3 0 2 2 7 0 2 2 3 3 0 2 2 2 16 3 1 15 2 13 15 2 9 9 7 9 9 2 2
23 10 0 9 2 3 10 9 13 2 15 15 13 2 7 3 3 15 13 9 7 3 9 2
9 9 13 9 2 7 7 14 15 2
23 9 1 12 0 9 2 3 16 9 1 0 9 7 10 9 2 13 3 9 10 0 9 2
5 13 3 1 9 2
50 7 7 16 4 13 7 15 13 1 9 15 10 9 7 15 3 13 1 9 2 15 11 13 2 16 4 15 2 15 13 1 10 9 2 13 2 16 13 1 9 2 13 15 3 0 9 1 10 9 2
20 3 1 9 2 1 15 15 10 9 13 2 13 3 0 9 0 1 9 11 2
48 13 1 15 2 7 15 3 2 9 15 2 15 15 1 9 13 2 15 13 0 1 10 9 1 9 0 7 15 2 15 13 9 11 2 15 13 1 9 9 7 9 7 3 15 1 15 13 2
8 13 3 10 9 1 0 9 2
7 16 9 2 3 0 9 2
11 16 9 2 14 2 1 9 2 0 9 2
24 10 0 9 2 3 13 9 11 9 2 16 1 9 10 9 7 9 4 1 0 9 13 9 2
36 15 2 16 1 0 15 13 0 1 15 2 15 13 9 0 2 7 3 0 2 15 13 1 15 2 15 1 0 9 13 7 13 1 0 9 2
14 11 13 9 2 15 13 1 9 10 9 0 9 9 2
10 15 13 9 9 2 15 13 10 9 2
12 11 0 0 9 11 13 9 9 0 9 13 2
15 1 15 13 9 7 1 0 9 1 9 10 9 13 9 2
14 10 9 15 3 13 0 9 2 15 13 1 0 9 2
7 3 11 13 9 0 9 2
12 13 1 0 9 3 2 16 15 13 1 9 2
22 12 13 9 15 2 16 9 13 3 16 15 2 15 3 13 2 15 13 0 7 0 2
25 1 9 13 7 9 15 2 1 15 13 2 9 1 9 10 9 2 9 15 2 15 13 0 9 2
21 7 13 13 13 1 15 2 15 13 1 15 2 14 3 7 3 1 0 9 9 2
7 7 7 15 13 1 9 2
43 14 2 9 0 9 2 2 15 3 13 1 9 2 2 13 15 1 9 7 9 2 15 13 1 9 11 3 13 2 13 16 0 9 2 0 3 1 9 1 9 0 9 2
32 4 15 7 13 1 15 13 9 9 2 3 15 13 11 10 9 2 7 15 13 1 9 2 9 2 2 3 15 13 15 15 2
30 3 2 16 15 13 9 2 15 15 2 3 3 16 0 1 10 0 9 2 13 0 13 0 0 7 0 9 7 9 2
13 14 3 13 3 0 13 1 11 0 9 3 9 2
21 14 3 15 13 13 1 9 7 1 10 9 7 9 2 15 13 9 10 0 9 2
19 0 9 15 15 2 15 13 0 9 2 13 13 1 9 9 7 0 9 2
28 1 0 9 0 9 2 1 15 4 13 12 0 9 7 12 0 9 2 13 9 1 9 9 1 15 3 13 2
19 1 10 9 2 1 15 9 9 9 7 9 3 13 2 13 10 0 9 2
9 13 15 13 1 0 9 7 9 2
31 7 10 9 13 13 1 9 2 7 1 9 2 16 1 15 2 3 0 9 2 13 9 1 9 2 15 13 3 16 9 2
2 9 9
22 13 15 2 16 1 12 9 15 14 1 12 0 9 9 13 1 15 2 15 15 13 2
11 1 0 12 0 9 13 3 9 9 9 2
19 15 13 1 0 9 0 2 13 1 9 9 0 9 7 9 3 0 9 2
8 1 9 9 13 3 0 9 2
15 1 0 9 15 1 10 9 13 15 0 2 9 1 9 2
5 9 13 0 9 2
12 3 0 9 1 15 3 13 0 9 0 9 2
4 9 13 0 2
22 0 9 2 16 4 13 9 2 13 13 2 0 2 9 2 7 3 0 9 13 9 2
38 0 9 9 2 1 9 9 13 10 7 15 0 9 7 9 15 2 2 15 9 13 14 0 9 9 2 14 10 9 2 7 3 0 9 9 0 9 2
27 1 0 9 15 9 2 13 3 1 0 9 2 7 14 1 15 2 13 14 3 1 9 2 7 1 9 2
27 3 13 7 13 2 13 9 1 9 2 13 9 1 9 10 7 15 9 2 1 9 1 10 7 15 9 2
9 0 9 1 9 3 13 15 9 2
7 9 9 9 15 3 13 2
24 9 3 13 0 13 15 1 10 9 1 9 2 7 14 3 13 1 10 9 9 0 1 9 2
9 13 15 1 9 0 2 7 0 2
33 3 13 2 13 1 9 9 2 3 15 1 9 9 13 2 7 15 2 16 13 0 2 13 13 9 9 16 0 2 9 9 2 2
26 9 1 9 9 9 13 13 7 3 2 16 13 1 9 2 3 13 15 9 0 9 7 13 9 9 2
10 10 9 13 13 1 9 7 3 13 2
35 0 9 9 13 1 15 2 16 15 13 1 9 0 9 9 2 7 3 1 9 0 9 0 9 2 16 3 0 9 1 9 13 7 13 2
10 7 9 13 9 2 15 10 9 13 2
10 3 13 9 1 2 0 9 2 0 2
25 3 15 15 13 9 13 1 0 15 9 9 2 13 3 0 7 0 9 2 15 13 0 9 9 2
15 7 3 2 9 9 13 9 1 0 9 2 15 9 13 2
42 1 1 0 9 9 13 0 14 9 0 9 2 3 0 13 7 9 2 3 15 0 9 13 1 10 0 9 1 9 7 13 15 1 9 2 16 4 13 15 7 15 2
4 0 9 13 13
19 9 9 13 9 2 16 15 15 1 15 13 0 9 3 1 9 9 7 9
25 1 0 9 13 3 0 3 0 9 9 1 9 9 7 15 2 16 13 3 1 9 0 9 9 2
18 9 13 2 7 13 13 2 16 0 0 9 13 9 15 9 0 9 2
24 1 15 9 9 7 0 9 13 9 1 0 9 0 0 9 7 0 9 16 11 11 7 9 2
24 9 9 13 0 9 9 1 9 1 0 9 7 9 2 16 9 0 9 9 0 9 13 3 2
20 13 7 1 15 2 16 9 9 13 1 15 0 1 0 2 14 1 0 9 2
8 9 9 13 3 9 0 9 2
19 10 9 9 4 10 9 13 9 9 7 0 0 9 2 13 0 15 13 2
26 1 15 3 15 3 4 9 1 0 9 13 2 16 3 15 15 4 13 13 3 9 7 9 1 9 2
20 0 9 1 9 9 7 9 0 9 2 7 3 0 9 9 2 13 0 9 2
18 15 13 7 0 0 9 1 9 9 2 0 0 9 7 0 0 9 2
8 15 9 9 7 0 9 13 2
21 9 9 3 13 9 2 16 15 15 1 15 13 0 9 3 1 9 9 7 9 2
10 12 1 10 0 15 9 13 9 9 2
16 13 0 2 7 3 0 13 2 16 4 15 0 9 15 13 2
12 7 10 0 9 2 15 13 2 9 3 13 2
19 3 2 9 9 9 9 4 1 10 9 13 0 13 1 9 9 7 9 2
6 13 15 3 9 9 2
40 0 9 3 13 2 16 9 2 3 13 9 0 9 13 2 13 1 9 0 9 9 7 16 13 3 3 0 0 9 1 9 1 9 2 3 13 9 9 13 2
33 13 15 3 7 1 15 2 16 9 9 9 7 0 9 1 11 13 1 9 9 0 9 1 12 9 1 12 5 1 0 12 9 2
21 13 15 7 1 0 0 9 9 1 9 2 15 13 1 9 0 2 7 1 9 2
15 13 2 16 10 7 15 9 13 13 1 9 2 13 0 2
26 0 9 9 13 7 3 0 9 7 0 9 2 13 9 2 15 0 9 1 0 9 1 9 3 13 2
22 13 3 0 2 16 9 9 13 3 3 1 0 9 7 16 15 0 9 1 9 13 2
23 13 15 3 9 2 3 9 13 3 10 9 9 2 3 15 0 9 13 2 7 9 0 2
13 3 2 16 13 3 9 1 9 9 11 1 15 2
24 13 1 15 13 9 0 9 2 3 2 3 9 9 1 0 9 13 3 12 9 1 9 9 2
37 13 4 3 0 13 2 16 9 0 9 7 0 9 2 13 2 0 9 7 15 2 7 16 9 0 9 1 0 9 13 1 15 0 16 9 9 2
24 15 2 16 4 9 1 9 13 9 1 11 2 15 1 10 9 13 0 9 2 3 15 13 2
7 3 15 7 13 0 9 2
25 9 2 15 13 0 0 9 1 0 7 10 0 9 2 15 3 13 1 15 2 15 13 0 9 2
19 3 13 9 7 9 0 9 3 2 7 16 15 13 9 2 3 15 13 2
22 3 15 13 0 9 2 15 15 7 9 0 9 4 1 0 9 9 3 7 3 13 2
7 9 13 0 7 0 9 2
24 13 9 1 15 2 16 9 7 9 0 9 1 0 9 13 9 9 1 0 9 1 0 9 2
4 11 11 1 9
24 0 9 9 13 0 0 9 9 1 9 0 2 0 9 7 3 15 1 15 13 0 9 9 2
42 1 9 9 2 3 13 1 9 0 9 2 15 0 9 1 10 9 13 9 3 15 2 10 9 13 1 12 9 2 9 1 11 7 0 9 11 1 9 9 1 9 2
17 0 9 2 9 7 11 13 1 9 3 0 2 1 9 1 9 2
18 9 11 15 0 9 13 2 16 13 9 1 12 9 0 11 7 11 2
30 1 0 2 7 0 2 9 13 9 1 11 2 11 2 11 2 11 7 11 2 13 1 9 7 9 1 9 9 2 2
27 11 15 7 1 9 1 0 9 0 11 13 13 9 9 16 15 2 15 3 13 2 9 9 1 0 9 2
17 2 0 15 9 9 13 0 9 2 15 9 13 1 9 0 9 2
10 9 9 4 13 9 13 2 2 13 2
10 13 9 9 7 13 2 15 15 13 2
12 13 15 3 7 9 15 1 0 9 3 13 2
17 1 9 9 11 15 9 0 9 1 0 9 13 7 3 15 13 2
10 3 2 16 4 15 13 7 0 9 2
21 13 15 3 9 3 10 9 2 15 15 10 9 13 3 2 11 2 11 7 11 2
20 1 9 0 9 0 9 16 2 3 0 2 15 13 13 7 0 9 10 9 2
4 9 1 11 2
23 1 0 2 0 7 0 9 14 0 2 0 2 9 13 13 9 0 9 1 10 0 9 2
17 9 0 9 13 1 9 9 2 0 0 9 7 13 14 15 2 2
7 9 13 1 9 3 3 2
31 13 2 16 15 13 9 9 0 9 11 11 11 2 11 2 15 1 0 9 13 1 2 9 9 11 2 0 9 1 9 2
26 1 9 0 0 9 9 11 11 13 2 0 0 9 2 11 1 0 0 9 7 2 9 9 12 2 2
16 2 11 13 0 0 9 1 0 0 9 2 2 13 10 9 2
17 1 10 0 9 13 2 16 3 3 3 13 2 3 0 13 9 2
9 11 11 15 15 10 0 9 13 2
5 13 3 0 9 2
15 9 13 15 13 9 0 9 15 13 0 9 1 0 9 2
27 2 0 0 2 15 15 1 7 1 2 15 15 10 9 13 13 2 13 13 3 2 16 11 1 9 13 2
7 13 15 2 16 3 13 2
14 3 2 3 4 3 13 0 0 13 2 13 3 3 2
8 0 9 13 0 9 1 0 9
26 9 13 0 2 3 13 3 2 15 13 2 13 4 15 13 9 11 11 2 15 13 0 9 0 11 2
16 9 11 2 15 10 9 3 13 2 15 15 13 13 3 9 2
20 9 9 1 0 9 7 3 13 1 9 1 2 9 2 2 15 13 9 11 2
8 2 9 13 0 2 3 0 2
20 13 4 15 1 9 2 2 13 9 9 0 11 2 15 3 3 3 13 11 2
15 1 9 13 9 3 13 11 7 10 0 9 1 9 11 2
22 13 13 2 0 9 2 2 9 9 9 11 1 9 7 0 9 0 9 11 1 9 2
35 9 2 9 2 9 7 3 7 9 2 15 0 9 0 11 1 11 13 2 13 9 2 16 15 13 0 9 0 9 1 9 11 7 11 2
25 0 0 11 2 15 13 1 10 12 9 9 0 0 9 1 11 0 11 2 13 1 11 0 9 2
16 0 11 2 3 14 0 2 15 3 13 1 9 0 0 9 2
22 3 1 9 0 11 13 3 9 0 0 9 2 11 2 15 9 13 1 9 0 9 2
16 1 11 15 3 13 9 9 15 11 2 3 0 1 10 9 2
19 11 13 1 11 14 0 2 7 3 0 2 1 10 9 13 9 9 9 2
17 1 9 11 15 13 1 0 9 3 0 9 9 11 7 0 11 2
17 2 7 16 15 11 13 3 1 11 2 13 2 16 1 15 13 2
21 13 4 1 15 9 9 7 13 2 16 13 13 2 2 13 1 9 9 9 9 2
13 1 10 9 11 13 11 9 2 15 13 1 11 2
15 11 3 11 13 2 16 4 15 10 9 13 1 0 9 2
13 1 0 9 9 11 1 0 9 3 13 9 9 2
32 16 1 15 3 0 0 9 13 7 1 11 11 0 0 9 2 15 15 13 2 13 15 13 9 9 2 1 9 1 0 9 2
19 0 9 7 0 9 11 14 13 9 2 16 9 12 9 13 3 9 9 2
10 1 0 9 13 9 1 11 7 9 2
18 0 1 15 2 11 2 13 0 9 0 11 2 15 9 12 15 13 2
14 11 3 13 9 11 2 3 7 0 13 9 0 9 2
18 0 11 15 1 9 0 9 3 7 1 0 11 3 13 9 11 11 2
30 3 15 4 11 7 11 13 13 1 0 9 0 9 2 7 0 9 0 9 2 1 15 4 13 10 9 7 10 9 2
7 3 3 0 13 9 11 2
9 11 3 13 0 9 2 0 11 2
8 3 14 13 9 11 2 2 2
14 3 0 9 9 15 13 13 9 11 1 11 11 11 2
23 1 10 9 4 13 9 11 1 12 2 9 13 9 9 2 0 9 9 7 0 9 9 2
11 9 4 15 13 13 1 9 1 10 9 2
19 9 9 11 13 9 9 1 9 9 7 15 2 16 3 13 0 9 11 2
34 11 9 15 1 9 1 0 9 1 0 9 13 1 0 9 2 2 11 13 9 2 16 9 11 13 3 0 9 1 0 0 9 2 2
9 0 9 13 0 2 15 0 9 2
17 0 2 15 15 1 9 13 2 13 9 2 9 2 9 7 9 2
29 9 11 2 16 2 16 13 9 2 13 1 0 9 9 2 0 9 2 7 13 15 1 9 2 2 3 13 13 2
6 2 0 11 2 1 11
33 11 13 1 0 0 9 1 0 9 2 15 13 10 9 2 13 15 9 11 2 15 3 3 13 3 3 1 11 1 11 7 3 2
23 11 13 1 12 9 0 9 1 9 11 7 11 13 7 1 11 0 0 9 1 0 9 2
35 9 11 1 9 11 2 3 1 9 9 13 12 9 9 1 9 2 15 3 1 15 13 0 9 11 2 3 15 13 0 0 9 0 9 2
24 11 13 3 0 0 9 9 2 1 15 13 9 3 0 2 16 13 1 9 1 0 0 9 2
33 10 9 15 13 13 15 1 0 9 1 0 9 1 0 9 2 7 9 16 0 2 7 0 9 15 3 13 1 12 2 9 13 2
21 11 13 10 9 2 16 3 0 11 4 13 13 3 7 13 15 1 9 0 9 2
26 15 15 7 3 13 2 16 13 2 16 0 0 9 13 1 10 9 0 9 1 9 7 9 15 9 2
36 11 7 13 1 0 0 9 1 0 9 2 15 13 10 9 2 13 15 9 0 9 11 2 15 3 3 13 3 3 1 11 1 11 7 3 2
24 11 13 1 12 9 0 9 1 0 9 11 7 11 13 7 1 11 0 0 9 1 0 9 2
20 13 7 9 2 16 11 13 9 9 2 16 4 15 13 13 1 9 0 9 2
7 7 3 15 7 13 0 2
31 1 11 13 1 10 0 9 13 7 9 2 16 0 9 13 13 9 7 9 9 13 1 9 9 2 15 13 13 0 9 2
18 3 1 9 0 9 13 1 11 3 12 11 3 7 13 1 0 9 2
19 3 15 13 1 11 1 12 9 7 0 1 15 13 1 15 0 0 9 2
28 13 1 15 0 9 2 10 0 9 13 1 11 7 9 15 1 15 13 7 13 2 16 0 9 13 10 9 2
13 3 9 9 13 0 9 12 11 3 1 0 9 2
15 13 1 15 9 9 2 15 1 10 9 3 13 1 11 2
16 0 0 3 1 9 7 9 13 9 2 15 15 1 9 13 2
12 0 0 9 13 1 10 0 9 9 9 9 2
10 3 7 13 13 1 9 11 0 9 2
16 15 9 1 9 15 13 1 9 1 9 0 9 1 9 12 2
24 0 9 0 9 15 7 13 2 16 11 13 3 0 9 7 13 15 13 15 3 9 0 9 2
5 11 15 7 13 2
31 1 9 1 9 0 9 13 1 10 0 9 2 16 16 4 15 13 2 7 4 13 2 13 15 1 11 0 9 3 9 2
12 1 15 15 13 1 9 7 9 9 11 11 2
13 15 9 13 9 7 1 0 9 4 13 3 0 2
27 0 1 15 13 1 11 1 0 9 7 3 10 9 15 13 1 9 2 16 1 15 13 13 9 3 0 2
12 15 15 3 13 13 9 1 0 9 1 11 2
26 0 13 0 9 2 15 4 13 1 9 1 0 9 2 0 1 9 1 9 2 9 1 15 1 0 2
16 15 13 13 3 1 9 9 2 15 15 13 7 13 1 9 2
26 11 11 13 1 15 2 16 1 9 2 1 15 13 11 1 0 9 2 15 0 7 0 9 3 13 2
9 13 15 15 3 13 9 1 9 2
47 11 11 1 9 1 0 9 1 9 0 9 13 7 1 9 10 9 4 13 2 16 0 9 13 0 9 10 2 0 11 2 1 9 11 2 7 0 9 13 1 9 7 13 3 1 11 2
44 13 2 16 4 13 1 9 0 0 9 9 1 9 10 0 0 9 2 7 15 2 13 2 13 3 1 0 9 2 3 1 9 9 13 7 0 9 0 9 9 1 0 9 2
5 11 7 11 13 9
32 16 1 0 9 1 9 0 9 13 3 3 3 9 2 9 1 0 9 1 0 9 13 3 3 2 3 1 9 9 2 0 2
10 0 9 13 13 10 9 1 0 9 2
37 13 15 3 9 2 16 9 11 4 13 3 2 16 4 15 0 9 13 2 7 15 15 13 2 16 0 9 13 9 2 15 13 13 7 0 9 2
11 3 13 1 10 9 1 0 9 0 9 2
10 9 9 15 7 13 3 1 9 9 2
25 1 0 9 1 0 9 1 9 15 9 13 0 9 2 16 4 1 9 12 13 13 7 0 9 2
9 15 13 1 0 9 1 0 9 2
26 15 15 13 13 2 7 3 15 13 1 9 2 12 7 12 9 9 2 15 3 0 9 1 11 13 2
26 9 0 9 1 9 2 0 9 9 0 0 9 2 11 11 4 13 16 0 9 1 9 3 0 9 2
9 3 13 10 0 9 9 11 11 2
12 1 10 9 15 13 2 16 11 3 3 13 2
17 1 9 15 13 2 16 0 0 9 4 13 13 3 1 10 9 2
9 9 9 15 1 0 9 3 13 2
30 0 9 4 13 2 16 15 13 9 0 9 11 11 2 0 9 9 2 15 4 13 11 11 1 0 9 1 9 12 2
12 0 9 13 0 9 11 11 2 0 0 9 2
20 13 3 1 15 0 9 2 7 0 9 13 1 15 3 3 14 3 0 9 2
18 3 9 15 13 0 9 9 11 11 7 10 9 1 9 9 11 9 2
13 12 7 3 3 13 2 16 15 1 9 13 4 2
13 1 3 0 9 4 15 13 13 13 3 10 9 2
39 0 9 15 4 13 1 9 2 16 3 1 9 3 3 13 9 13 9 7 9 9 2 16 0 9 1 0 9 1 9 13 3 13 11 11 7 11 11 2
25 1 10 9 15 13 1 9 11 11 2 11 2 2 11 11 2 11 2 7 11 11 2 11 2 2
14 1 9 4 13 11 7 11 13 11 11 7 11 11 2
13 13 13 7 1 0 0 9 7 9 9 9 11 2
28 1 9 1 0 9 2 15 13 4 13 2 9 1 9 9 15 13 0 9 1 9 2 14 1 9 0 9 2
37 13 15 9 2 16 0 9 0 9 4 13 13 9 2 9 9 0 11 11 11 11 2 15 1 15 13 0 7 0 9 1 0 9 1 9 9 2
21 10 9 4 0 9 11 11 2 16 3 15 13 15 2 3 13 1 9 1 9 2
22 9 13 13 0 9 11 7 10 0 0 9 2 15 15 1 9 7 10 9 3 13 2
13 7 1 10 9 13 3 1 0 9 3 3 3 2
12 11 11 11 2 11 1 10 12 9 0 9 2
19 10 9 13 15 1 0 9 9 15 13 12 9 9 7 12 9 0 9 2
4 9 1 0 9
22 1 0 0 9 4 1 0 9 13 0 9 11 11 11 1 9 0 9 2 11 2 2
13 11 2 11 15 13 12 2 9 12 1 0 9 2
7 13 9 0 9 1 11 2
23 1 9 12 13 9 0 0 0 0 9 2 11 2 7 13 15 16 9 9 0 0 9 2
31 1 9 15 13 3 9 9 11 1 0 9 1 9 7 9 7 3 13 1 9 12 7 12 9 9 9 11 1 0 9 2
29 1 9 12 1 9 12 13 0 0 9 11 7 1 9 12 2 12 13 1 0 0 9 1 0 0 9 1 9 2
13 1 9 12 15 13 0 9 11 1 9 11 11 2
20 1 9 1 0 0 9 11 11 13 11 3 9 9 16 9 1 9 1 9 2
20 13 3 9 1 0 0 0 9 7 9 13 7 1 0 0 9 1 9 12 2
25 1 0 3 0 11 15 13 11 9 0 9 9 0 9 2 11 2 7 9 9 1 0 0 9 2
15 1 9 1 9 12 15 16 9 0 0 9 13 9 11 2
9 11 13 0 7 13 9 7 9 2
4 11 13 9 11
39 9 0 9 0 9 11 11 2 15 13 0 9 1 9 1 11 2 13 2 16 11 13 0 13 1 0 9 0 9 1 9 9 1 10 9 1 0 9 2
36 13 2 14 1 9 0 9 0 9 1 9 7 0 9 1 0 9 7 1 9 2 13 10 9 3 1 9 2 13 0 9 0 0 11 11 2
21 0 9 13 9 9 2 15 1 0 9 2 3 13 1 9 2 13 1 9 11 2
36 13 14 0 9 13 15 3 1 9 2 7 3 3 13 14 14 13 0 9 1 9 7 13 3 9 2 15 4 15 13 3 13 1 9 9 2
21 0 9 9 13 1 15 2 16 9 0 9 13 9 9 2 15 4 13 1 9 2
16 0 9 13 1 9 9 0 9 0 15 9 2 11 11 11 2
31 13 9 13 9 9 0 9 0 9 2 15 13 14 1 9 7 15 4 13 14 7 2 16 4 15 9 13 9 0 9 2
7 0 9 13 1 0 9 2
33 0 9 13 13 14 1 0 9 2 7 15 3 14 1 9 2 16 0 11 4 3 13 0 9 7 9 15 13 9 7 0 9 2
1 3
11 0 9 0 11 3 13 0 9 11 11 2
14 1 9 13 9 1 0 9 11 9 7 1 0 9 2
7 13 15 3 9 11 12 2
32 0 9 0 9 11 11 2 11 13 1 0 9 2 16 10 9 13 1 0 9 0 15 0 9 1 9 0 0 9 1 11 2
25 13 13 1 9 0 9 11 1 11 2 16 4 0 9 1 9 10 9 13 7 1 12 2 9 2
14 9 0 0 9 1 11 9 3 13 0 9 11 11 2
11 3 13 1 9 0 0 9 1 0 9 2
20 0 0 0 9 11 3 13 2 16 10 9 1 0 0 9 13 11 2 11 2
21 10 9 4 13 9 9 13 0 9 11 2 11 2 12 2 2 15 13 0 9 2
30 0 9 9 2 15 4 13 13 3 9 0 9 0 9 0 9 2 11 2 2 4 3 13 1 0 9 9 0 9 2
9 0 9 3 1 11 13 0 9 2
32 0 0 9 2 11 2 2 15 15 13 1 3 0 0 0 9 9 0 9 7 13 3 1 9 2 3 13 7 9 1 9 2
20 0 9 3 13 9 11 2 11 2 16 4 13 9 9 10 9 11 2 11 2
22 9 13 11 1 9 9 7 13 3 3 3 9 2 15 3 0 9 13 1 0 9 2
18 9 9 0 0 9 1 0 2 11 15 13 1 12 2 3 13 9 2
25 9 2 15 3 13 0 0 9 1 9 0 2 11 2 13 0 9 1 0 2 11 1 9 9 2
9 1 12 9 13 9 9 3 9 2
5 11 1 9 0 9
2 11 2
33 0 9 15 1 0 12 9 4 13 3 1 15 2 16 4 4 13 15 2 15 3 4 1 11 13 2 7 13 10 0 0 9 2
28 13 15 1 9 9 0 9 9 11 11 2 15 3 1 11 9 0 9 13 0 9 0 9 1 9 12 9 2
17 1 9 11 13 3 0 9 11 7 9 0 9 11 1 9 12 2
4 9 13 0 9
2 11 2
18 2 1 0 9 2 13 3 9 11 11 9 0 9 0 9 11 11 2
16 1 0 9 1 11 3 3 13 9 3 0 9 11 11 11 2
21 1 11 2 0 9 2 3 11 2 11 13 1 9 2 13 0 7 0 9 2 2
18 2 16 9 13 0 3 13 2 13 0 13 0 0 9 2 2 13 2
5 11 2 9 0 9
2 11 2
37 0 9 1 9 0 11 4 13 4 13 2 3 3 2 3 1 9 2 2 13 0 9 9 11 11 1 0 9 1 0 9 1 0 11 11 11 2
29 3 3 11 13 2 13 4 15 3 3 1 10 0 9 13 3 1 9 9 2 16 4 13 0 9 9 0 9 2
15 15 4 13 4 13 9 1 11 7 1 11 1 0 9 2
24 1 10 9 4 1 9 1 0 9 11 13 9 2 15 1 0 0 9 13 0 9 12 9 2
26 11 2 11 3 13 2 16 13 1 9 9 1 9 0 9 13 1 9 1 9 0 9 1 0 11 2
25 9 0 9 0 9 11 2 11 3 13 11 2 16 13 3 0 2 16 13 1 9 0 0 9 2
6 11 13 14 0 0 9
2 11 2
27 11 13 1 9 0 9 0 0 9 2 13 1 9 1 0 9 0 9 11 0 0 9 0 9 11 11 2
18 13 2 16 11 13 9 9 2 15 4 3 13 10 9 1 10 9 2
20 2 13 15 9 2 1 15 15 13 7 15 15 13 10 0 9 2 2 13 2
21 9 0 9 13 2 16 9 13 13 13 9 2 16 1 15 11 13 2 9 2 2
24 11 13 13 0 9 1 9 0 9 2 11 2 2 10 9 13 1 9 2 16 9 13 11 2
40 0 9 2 15 4 3 13 2 16 13 12 7 12 0 9 7 9 0 7 0 9 2 15 1 10 9 3 13 2 7 15 13 2 16 9 1 0 9 13 2
4 1 11 13 9
10 0 9 13 0 9 1 11 7 13 11
4 11 2 11 2
22 9 0 7 0 9 15 1 9 0 0 9 9 3 13 1 9 9 1 0 9 11 2
24 16 13 0 0 0 9 11 11 2 9 10 9 13 13 9 0 2 9 0 7 9 0 9 2
16 11 1 9 9 9 3 13 2 16 12 0 9 13 0 9 2
14 1 0 9 9 15 0 9 13 1 11 3 1 9 2
32 0 9 2 0 9 0 9 2 3 13 0 9 9 0 9 1 11 7 9 0 0 9 1 9 0 9 7 1 9 0 9 2
26 1 0 9 2 1 15 15 13 0 9 9 2 9 3 13 9 3 15 13 1 0 9 9 0 9 2
32 9 0 9 3 3 13 0 9 0 0 0 9 1 9 9 0 9 1 9 7 13 15 1 0 9 7 9 1 0 9 11 2
22 11 15 13 0 0 9 2 10 9 3 13 1 0 9 0 9 2 13 1 9 9 2
16 0 9 1 0 9 13 2 0 9 11 1 9 0 9 2 2
16 13 9 1 15 2 16 4 1 0 0 9 0 9 3 13 2
5 11 2 9 1 9
2 11 2
24 1 0 0 9 11 3 1 0 0 9 13 0 0 9 1 9 3 12 9 9 1 0 11 2
27 13 15 15 9 11 3 0 9 11 1 9 11 11 2 0 9 9 0 9 11 11 11 7 0 0 9 2
24 0 9 11 11 11 2 11 13 9 2 16 4 15 13 1 9 0 9 7 9 1 0 11 2
50 1 9 2 15 4 13 9 9 2 11 2 11 13 2 16 13 0 13 1 9 9 1 9 7 13 9 0 9 1 11 7 11 2 3 3 4 13 10 9 12 9 7 9 4 13 1 9 1 9 2
25 11 7 11 1 10 9 13 9 9 9 3 16 12 9 0 7 0 9 1 11 2 11 7 11 2
5 9 1 11 1 9
5 11 2 0 11 2
25 0 9 11 2 15 3 3 13 1 0 11 2 15 3 13 7 1 0 0 9 13 1 0 9 2
22 9 13 12 9 9 7 12 9 9 0 9 11 1 9 1 9 7 9 1 0 9 2
17 0 9 13 9 9 1 11 3 11 1 9 9 2 0 0 9 2
11 9 15 7 3 3 13 1 10 9 13 2
13 1 0 13 9 11 9 1 9 0 3 1 11 2
7 3 13 7 3 0 9 2
26 0 9 11 11 1 9 13 9 13 11 0 9 0 9 2 16 11 13 11 7 0 0 9 0 11 2
15 1 11 15 13 0 9 0 9 2 15 15 13 4 13 2
7 9 13 0 2 0 9 2
10 9 13 13 3 0 0 9 1 11 2
15 1 10 9 13 0 3 13 0 9 2 1 15 13 9 2
11 1 11 15 3 13 0 9 11 2 11 2
11 9 0 9 11 2 11 1 9 13 0 2
4 11 13 0 9
2 11 2
24 9 11 11 13 1 0 9 1 9 0 9 9 2 16 10 0 9 15 1 15 3 3 13 2
9 13 15 1 12 0 9 0 9 2
19 1 10 9 11 1 9 13 1 9 9 12 9 2 16 11 15 3 13 2
23 12 1 9 3 13 2 16 11 4 13 1 0 9 0 9 13 3 9 16 10 0 9 2
23 1 9 11 4 13 11 13 1 0 9 1 12 9 9 2 16 11 4 13 1 12 9 2
27 9 1 0 0 9 3 13 2 16 1 9 0 9 0 9 10 9 15 13 0 9 0 9 11 2 11 2
21 12 1 0 0 9 1 0 9 11 2 15 13 3 1 10 9 1 9 0 9 2
19 1 0 9 15 9 9 13 12 0 2 12 9 13 13 2 12 4 13 2
11 3 16 12 9 13 3 13 1 0 9 2
6 11 13 9 9 7 9
2 11 2
25 9 11 3 13 11 2 3 12 1 0 0 9 2 1 9 9 7 9 2 3 9 3 13 9 2
26 1 10 9 9 11 1 0 9 13 0 9 9 11 2 16 4 13 10 9 7 13 1 9 9 9 2
27 9 1 11 1 15 13 2 0 2 0 7 0 9 7 9 0 0 9 7 9 2 15 1 15 13 2 2
7 0 9 13 10 9 0 9
29 9 2 15 13 1 15 2 16 0 13 10 7 15 9 1 9 2 7 7 1 0 9 13 2 15 13 13 0 9
29 0 9 13 10 9 0 9 2 15 2 15 13 10 9 2 13 13 3 1 3 0 0 9 2 7 7 0 9 2
17 10 2 9 2 3 9 1 0 0 9 9 13 1 12 9 9 2
11 13 1 0 9 0 9 3 13 10 9 2
21 13 15 15 13 7 0 9 2 15 7 13 13 0 9 2 15 1 9 3 13 2
15 3 3 13 2 16 4 9 1 9 13 1 9 12 3 2
4 13 15 13 2
20 15 2 16 15 3 9 7 10 0 9 13 2 3 9 3 13 9 15 13 2
14 9 1 9 13 3 3 3 2 3 1 3 0 9 2
13 1 0 9 1 9 13 9 7 9 1 0 9 2
13 16 0 9 13 3 1 0 9 2 3 9 13 2
23 15 13 13 2 16 9 13 13 3 1 9 1 9 2 7 15 13 13 13 1 10 9 2
16 13 7 3 0 2 16 7 3 9 3 3 9 1 9 13 2
16 7 13 3 0 2 16 1 9 0 13 3 3 7 3 9 2
5 13 3 1 9 2
37 13 15 3 7 9 2 3 9 9 13 1 9 9 0 9 3 2 15 10 9 2 1 10 0 9 13 7 0 9 2 3 3 16 13 2 2 2
22 1 0 9 13 9 7 3 9 13 1 9 10 0 9 1 9 9 7 9 1 9 2
15 10 9 15 1 9 9 7 9 13 13 2 14 0 13 2
23 16 0 9 2 3 9 2 0 9 13 0 2 13 15 9 1 10 9 13 3 0 9 2
16 9 1 9 7 13 2 16 7 10 9 10 0 9 3 13 2
8 9 13 13 2 7 15 9 2
20 9 2 15 13 0 13 13 9 7 9 1 9 1 9 2 0 9 3 13 2
13 3 0 9 13 9 2 15 13 0 7 0 9 2
9 0 9 15 1 10 9 3 13 2
6 13 15 15 3 13 2
16 10 9 9 13 1 9 3 1 9 3 3 0 7 3 0 2
25 3 15 13 1 0 0 9 2 15 13 13 1 0 9 2 7 3 15 15 13 13 3 0 9 2
9 0 7 0 9 13 12 1 15 2
9 13 4 0 2 16 4 13 0 2
10 3 15 9 0 9 9 4 13 13 2
15 9 15 3 3 2 3 1 9 0 9 2 13 1 9 2
27 0 0 9 4 1 0 9 13 1 9 9 12 2 3 1 9 0 9 1 0 2 0 7 0 0 9 2
3 0 9 2
33 3 1 0 9 13 0 9 2 12 2 9 10 2 9 2 2 9 2 10 9 13 2 2 0 9 9 3 13 3 3 0 9 2
13 0 9 7 9 3 13 2 7 2 2 2 2 2
34 9 2 7 2 1 12 9 3 16 9 9 0 9 2 2 13 1 9 2 15 15 9 3 13 15 2 2 13 2 15 13 1 9 2
20 15 1 9 0 9 1 12 9 9 2 15 9 9 13 1 9 9 1 11 2
22 9 15 3 2 1 0 2 13 13 0 9 9 1 0 7 0 2 0 7 0 9 2
30 1 0 9 3 13 9 0 0 9 2 15 13 3 0 9 7 9 9 2 7 15 3 13 9 9 9 1 0 9 2
5 10 9 13 0 2
15 16 15 1 15 13 2 13 15 2 16 15 15 3 13 2
26 15 15 15 3 13 2 13 15 3 0 13 2 7 15 15 3 13 1 9 2 16 15 3 3 13 2
34 1 10 0 9 2 15 13 2 16 13 9 0 7 0 2 7 13 2 16 4 15 13 15 2 13 1 9 2 16 13 3 15 0 2
8 1 0 9 13 15 15 0 2
22 9 0 9 3 3 13 2 16 7 9 9 2 15 13 9 9 2 13 1 15 0 2
55 3 3 13 2 2 16 9 9 15 1 0 9 13 1 9 9 2 2 9 15 3 13 2 3 1 9 0 9 0 9 2 2 3 13 2 16 2 9 9 2 15 15 13 13 9 0 9 2 13 13 9 1 10 9 2
12 9 15 3 9 1 10 9 13 2 2 2 2
8 2 7 2 1 12 9 13 2
27 1 9 2 9 2 13 15 13 3 2 2 9 3 13 2 16 4 10 9 1 9 13 2 2 14 13 2
11 9 15 9 1 9 2 3 13 15 2 2
14 3 16 15 15 13 9 13 1 3 0 9 1 9 2
8 13 9 2 13 15 1 9 2
6 0 9 4 3 13 2
23 10 9 2 3 0 9 2 15 3 13 2 16 15 13 9 9 9 1 0 9 10 9 2
16 12 1 10 9 13 9 0 9 9 0 1 3 0 9 9 2
23 9 9 0 9 13 1 0 9 13 10 9 2 16 13 0 2 16 13 9 7 9 0 2
36 13 2 16 15 13 13 1 9 2 15 0 9 13 1 9 0 9 2 3 16 1 9 10 9 2 7 0 9 1 0 9 10 9 13 0 2
16 13 0 9 2 15 13 7 1 0 9 2 7 1 0 9 2
8 15 13 9 10 9 2 13 2
14 3 14 0 9 2 3 7 9 2 15 1 9 13 2
22 9 9 0 9 13 1 0 9 13 10 9 2 16 13 0 2 16 13 9 7 9 0
3 15 13 9
13 3 1 9 0 9 4 13 13 0 9 0 9 2
23 0 9 1 9 7 0 0 9 1 9 9 1 9 15 1 0 9 13 13 14 0 9 2
14 1 0 9 7 0 9 10 9 15 13 0 9 9 2
21 15 13 9 9 1 9 9 9 1 9 12 9 2 0 14 9 1 0 0 9 2
39 16 3 15 1 15 13 15 2 3 0 9 9 7 0 9 2 15 15 3 1 9 13 10 0 0 9 2 13 1 12 2 9 9 3 13 0 3 13 2
25 0 9 7 0 0 9 13 9 3 9 13 15 9 0 1 9 0 0 9 1 9 0 0 9 2
30 15 15 13 13 9 1 0 0 9 2 13 10 9 13 3 1 0 9 0 9 7 13 13 1 9 1 0 0 9 2
12 15 1 9 0 9 7 0 0 9 0 13 2
32 0 0 9 2 7 16 3 3 0 2 13 1 0 0 9 13 3 9 1 9 1 9 7 9 0 0 9 1 0 0 9 2
26 0 0 9 2 15 9 9 4 13 1 9 2 3 3 13 9 9 7 9 1 10 9 9 1 9 2
23 1 9 9 0 9 1 9 7 1 9 1 0 0 9 15 3 4 13 3 10 9 13 2
17 3 14 1 9 2 16 15 9 13 3 13 1 9 0 0 9 2
12 7 15 7 3 9 1 0 9 1 9 13 2
7 10 9 7 1 10 9 2
20 1 9 1 9 13 14 1 9 1 9 7 1 0 9 13 14 9 0 9 2
11 13 4 3 2 16 4 4 13 3 3 2
4 9 1 9 2
18 0 9 13 9 7 9 1 0 9 9 13 1 11 1 9 14 9 2
16 13 7 9 2 3 4 10 0 9 13 13 3 1 9 9 2
16 9 13 3 0 2 7 7 0 2 9 1 0 9 0 9 2
12 10 9 4 15 1 10 0 9 13 13 0 2
16 7 13 3 9 1 15 9 9 4 1 0 9 13 13 0 2
11 13 9 1 10 0 9 13 3 9 0 2
25 0 9 13 3 1 9 9 0 9 9 0 9 1 9 11 2 1 15 9 9 13 7 13 9 2
30 7 3 1 9 2 3 4 9 7 9 9 4 13 3 7 9 9 4 13 0 9 2 7 4 10 9 13 0 9 2
17 9 9 4 10 9 13 2 4 3 13 1 2 9 0 9 2 2
29 1 0 9 13 9 0 0 9 2 15 4 13 11 13 3 13 0 9 9 9 11 2 0 15 9 9 7 9 2
11 3 3 1 15 13 0 10 9 3 13 2
7 9 13 3 9 0 9 2
12 1 9 9 9 14 1 10 9 9 13 9 2
15 1 0 9 9 9 13 7 0 13 1 9 2 3 9 2
23 3 15 13 3 7 1 15 2 7 3 1 9 0 9 2 1 10 9 13 9 3 9 2
5 15 7 3 13 2
7 9 13 3 0 1 9 2
5 13 15 12 9 2
21 1 0 4 9 1 9 9 4 13 13 9 7 9 4 15 13 3 1 0 9 2
14 9 4 7 13 1 9 2 1 15 4 3 9 13 2
23 0 9 4 13 1 0 9 9 3 13 9 2 3 4 15 0 9 13 13 1 12 9 2
22 3 4 13 7 0 13 7 13 0 9 2 15 13 13 9 1 9 15 1 0 9 2
15 12 9 13 2 0 2 2 7 12 7 0 13 1 9 2
11 1 9 10 9 4 9 13 0 9 9 2
12 9 15 3 13 13 2 16 9 9 9 13 2
9 13 15 3 1 9 13 0 9 2
18 7 9 13 1 1 9 2 15 13 10 9 2 1 0 9 3 0 2
11 10 9 1 15 4 3 13 1 0 9 2
17 16 3 13 1 9 13 9 2 13 3 0 9 7 13 0 9 2
2 0 9
21 0 9 0 9 11 11 9 13 1 0 9 2 15 13 1 9 11 1 0 9 2
31 10 9 4 13 3 0 2 16 4 11 9 13 0 9 2 15 13 13 9 1 0 0 9 1 10 0 9 1 0 9 2
25 16 4 9 9 11 0 11 2 11 2 13 2 16 0 9 9 13 3 3 3 0 7 0 9 2
54 16 4 9 1 9 7 11 13 1 9 7 16 4 9 9 9 9 1 9 11 2 0 1 9 11 2 11 2 9 7 11 2 1 9 2 13 4 13 9 9 2 4 13 3 0 0 9 11 9 1 10 0 9 2
20 16 4 13 3 3 9 9 0 9 0 9 1 9 1 9 2 0 9 11 2
25 16 4 1 0 9 11 2 3 15 11 9 3 13 2 4 13 0 9 10 9 2 0 9 11 2
33 16 4 13 2 16 16 15 9 13 1 9 9 2 3 1 9 9 9 0 9 2 2 9 13 13 1 9 7 1 3 0 9 2
47 16 4 13 2 16 3 1 10 9 13 0 9 0 9 12 9 3 2 16 4 0 9 13 1 9 1 9 0 9 2 13 1 0 9 7 13 9 1 11 7 1 10 0 2 0 9 2
1 9
16 3 0 0 9 13 1 9 1 9 1 11 2 9 0 9 2
21 9 9 13 9 1 9 7 1 9 10 9 15 13 1 0 9 2 3 15 13 2
5 0 13 0 9 2
8 9 15 13 3 13 12 9 2
6 12 9 13 12 0 9
2 11 2
21 0 9 2 15 15 13 1 0 9 12 0 9 11 2 13 1 0 9 1 9 2
13 11 15 13 9 0 9 9 1 11 11 2 11 2
12 0 0 9 15 3 13 3 3 1 12 9 2
34 1 11 2 11 13 1 9 1 0 9 3 1 9 1 9 9 12 0 7 12 0 9 9 2 15 15 13 13 9 1 12 12 9 2
4 9 3 13 2
23 2 0 9 2 3 15 0 9 13 14 9 2 4 3 3 13 2 2 13 11 2 11 2
10 12 0 9 13 9 1 0 9 9 2
5 11 11 1 0 9
12 9 9 9 12 2 0 9 2 11 7 0 9
4 11 2 11 2
24 11 11 2 15 1 9 13 9 7 9 13 1 9 2 13 1 9 1 9 1 9 1 11 2
28 1 9 0 9 11 11 11 13 2 16 13 1 9 9 1 9 2 15 15 13 1 9 2 9 7 12 9 2
14 4 7 13 9 1 0 9 2 3 9 13 0 9 2
22 0 9 13 11 1 0 9 1 11 2 3 15 13 9 7 9 7 9 13 9 9 2
10 9 13 0 9 1 0 9 1 11 2
25 11 13 2 16 1 0 9 9 13 1 0 9 0 9 2 0 9 1 9 7 9 1 12 9 2
5 9 9 9 13 2
40 11 11 4 1 9 12 13 1 9 1 0 9 2 15 15 13 13 15 2 16 13 9 2 15 1 9 12 13 10 9 2 7 15 1 9 1 12 9 13 2
24 16 15 1 9 11 0 9 13 2 9 15 1 9 13 7 0 9 1 11 1 15 13 9 2
20 1 9 11 11 13 3 0 9 9 9 12 2 0 9 2 11 7 0 9 2
9 13 1 15 1 0 9 1 11 2
32 1 9 3 2 13 2 16 9 9 12 2 1 10 9 4 11 13 7 15 13 1 9 0 9 2 13 1 15 1 0 9 2
33 0 9 1 9 9 13 2 1 9 1 0 0 9 2 16 9 1 9 11 1 9 4 1 9 9 13 0 9 9 11 11 2 2
6 11 13 9 1 0 9
2 11 2
15 9 0 9 11 11 3 13 9 1 0 9 11 2 9 2
21 0 9 1 11 12 13 2 16 9 1 9 2 15 9 1 11 13 2 13 0 2
21 0 9 13 1 9 0 1 11 1 9 12 7 11 13 13 15 9 1 9 12 2
23 1 10 9 15 13 9 3 0 12 9 9 2 15 13 16 9 1 9 1 10 9 13 2
17 0 0 9 15 13 2 16 0 9 1 9 13 1 9 9 9 2
16 9 3 13 1 9 2 16 9 1 9 13 0 7 3 0 2
4 11 13 1 9
2 11 2
12 0 9 13 1 9 10 0 9 7 0 9 2
22 3 1 9 9 15 9 9 11 13 1 12 9 9 11 12 2 12 1 9 12 0 2
11 0 9 4 1 11 13 7 1 0 9 2
8 0 1 15 4 13 1 9 2
28 1 9 0 0 9 12 0 9 2 12 0 9 7 12 0 9 13 1 9 3 1 9 0 9 1 0 9 2
6 9 9 1 11 3 13
2 9 2
31 0 9 9 1 9 12 13 1 12 9 9 1 9 12 9 9 1 9 1 12 9 9 2 12 9 9 2 1 9 12 2
20 1 9 9 13 3 0 9 11 7 11 2 15 13 1 9 0 9 0 9 2
23 14 1 10 9 1 9 12 13 0 9 0 9 0 9 1 0 9 3 16 12 9 9 2
6 11 13 9 1 0 9
2 11 2
18 9 1 9 12 9 1 0 9 1 9 12 9 9 13 0 9 11 2
9 13 15 3 9 11 11 11 11 2
23 0 9 2 1 15 0 4 13 1 0 9 9 9 12 2 13 0 1 12 9 0 9 2
15 0 9 13 13 0 2 0 2 3 0 7 13 3 9 2
26 1 15 13 0 9 9 3 0 2 9 1 12 9 4 10 9 13 9 9 1 12 9 0 0 9 2
11 15 13 13 1 0 9 1 9 7 9 2
21 11 11 13 12 12 9 1 0 9 1 9 1 12 9 9 2 1 9 12 2 2
1 3
22 11 11 11 15 13 1 9 0 9 1 11 11 1 0 9 2 15 4 13 10 9 2
10 1 0 9 13 9 13 7 7 0 2
22 0 9 11 2 9 13 1 0 9 1 11 9 12 0 9 1 0 9 12 9 9 2
14 0 11 9 13 0 3 1 0 9 9 16 0 9 2
16 10 0 9 1 0 9 2 1 0 9 2 13 12 9 9 2
1 3
19 9 11 11 7 9 1 10 9 1 9 9 13 9 0 9 11 1 11 2
8 11 13 1 11 14 12 9 2
8 9 13 13 9 9 1 0 9
2 11 2
17 1 9 13 9 2 16 9 9 1 9 0 9 4 13 13 13 2
23 9 9 11 11 2 11 2 13 11 2 16 15 10 9 13 1 0 9 9 9 1 9 2
15 3 1 9 9 9 13 0 9 7 15 3 13 10 9 2
27 9 15 7 3 13 1 9 2 16 4 9 13 13 9 9 7 16 9 4 13 1 9 9 13 9 9 2
33 2 9 0 9 1 0 9 4 13 4 13 9 2 16 4 0 9 13 9 2 16 15 4 13 9 9 0 9 2 2 13 9 2
29 9 15 1 9 1 9 9 13 2 16 4 9 13 13 9 9 2 16 4 13 1 0 9 13 1 9 1 9 2
20 9 11 13 2 16 15 13 15 2 16 4 9 9 13 1 9 1 9 9 2
23 0 9 9 13 9 9 9 2 16 4 1 9 2 15 13 10 9 2 13 13 0 9 2
9 9 3 9 9 13 1 9 9 2
8 11 13 1 0 9 3 1 11
2 11 2
21 9 11 1 0 9 13 1 0 0 9 11 2 1 0 9 0 9 7 3 13 2
18 1 9 0 9 11 1 0 11 11 11 13 9 1 9 0 9 0 2
19 2 7 16 13 9 0 9 0 2 3 3 1 15 13 11 2 2 13 2
19 13 7 1 9 3 2 3 16 9 1 0 9 2 13 1 10 9 0 2
25 9 9 0 9 1 0 11 1 11 11 11 13 9 1 9 11 1 0 0 9 1 9 1 0 2
17 2 13 15 9 0 9 2 15 13 3 7 3 13 2 2 13 2
26 7 16 9 11 13 9 2 16 4 9 10 9 1 0 9 13 2 13 1 11 10 9 1 9 9 2
10 0 0 9 15 3 13 1 0 11 2
19 2 1 9 13 3 13 2 16 15 13 16 0 9 7 14 16 9 2 2
27 9 0 9 11 2 11 11 11 15 13 2 16 10 9 1 0 9 1 0 0 9 13 13 0 9 11 2
17 2 9 2 16 4 15 13 13 1 0 9 2 13 2 2 13 2
15 1 9 9 7 1 0 9 9 7 13 13 1 0 9 2
8 2 15 15 9 1 9 13 2
10 0 13 9 1 0 9 2 2 13 2
4 9 13 1 11
2 11 2
19 0 9 0 9 13 0 9 2 16 15 1 12 9 13 0 9 1 9 2
19 3 13 9 9 11 11 9 0 9 9 9 7 9 13 11 7 13 3 2
19 11 15 13 2 16 9 9 13 1 9 0 9 2 7 3 1 10 9 2
13 0 9 1 10 9 13 13 0 3 13 9 9 2
17 0 9 13 10 9 3 0 0 9 2 15 9 13 1 9 9 2
6 9 9 13 1 0 2
9 13 7 0 9 9 1 0 9 2
28 1 9 9 11 11 4 13 9 13 10 9 3 1 9 7 9 1 9 2 3 3 4 13 13 1 0 9 2
5 11 15 13 1 9
2 11 2
27 1 9 11 11 13 0 9 0 9 2 7 13 9 9 1 9 7 9 12 11 1 9 9 1 0 9 2
39 1 9 1 0 9 3 9 11 2 11 2 11 11 11 13 2 2 1 15 2 16 3 9 13 10 9 9 2 13 3 2 16 13 9 1 0 9 9 2
19 9 0 9 13 11 1 9 0 2 7 7 13 9 13 1 15 3 0 2
12 16 16 4 9 13 1 0 9 2 13 9 2
25 13 13 0 9 2 16 9 13 2 7 9 2 15 9 9 13 7 15 15 13 15 0 9 2 2
8 11 11 2 11 2 2 9 9
24 9 0 9 11 12 13 1 0 9 9 2 16 0 9 9 0 7 0 13 9 9 1 11 2
5 15 13 10 9 2
10 10 9 13 3 0 1 9 9 9 2
25 13 15 3 0 9 10 9 0 2 0 9 2 15 15 13 1 10 9 3 0 9 16 0 9 2
32 9 9 9 13 2 16 4 13 10 0 0 9 2 15 4 13 1 9 7 15 4 13 3 15 9 2 15 13 3 9 9 2
14 15 13 9 9 16 15 2 13 3 9 0 0 9 2
9 7 15 1 9 13 9 1 9 2
28 14 7 2 16 4 13 9 9 2 7 7 1 9 2 3 10 0 0 9 13 9 2 13 10 9 3 0 2
11 13 15 1 9 16 11 2 11 7 11 2
18 7 1 11 15 1 0 9 3 13 1 15 2 16 13 10 9 0 2
5 11 11 1 9 11
2 11 2
11 2 0 9 15 4 13 9 9 10 9 2
45 13 15 2 16 3 13 9 2 15 15 4 13 9 1 11 2 7 13 2 16 4 1 11 13 2 2 13 11 0 9 9 11 11 1 9 2 15 13 1 10 9 1 0 9 2
34 9 15 13 1 0 9 1 9 9 0 9 2 1 9 11 1 10 9 7 1 9 2 15 9 1 9 1 11 13 9 9 1 9 2
5 0 9 1 9 12
4 0 9 1 11
5 11 2 11 2 2
29 0 7 0 0 9 15 3 13 1 0 12 0 9 2 15 13 1 9 3 1 9 0 9 2 1 12 9 2 2
8 13 4 15 13 15 9 9 2
39 9 1 0 9 13 9 0 9 1 11 9 11 11 7 9 9 0 0 9 9 11 11 2 15 15 3 1 0 9 11 13 1 0 9 9 0 0 9 2
19 1 0 9 9 4 1 9 3 13 9 2 15 15 13 3 1 0 9 2
12 1 9 1 9 7 4 9 9 1 9 13 2
4 3 1 9 12
15 3 13 1 9 9 11 2 11 2 11 9 0 16 3 2
28 9 0 9 15 7 13 2 16 15 13 3 9 0 9 9 2 15 13 11 2 16 4 15 13 0 9 13 2
6 1 10 9 13 9 2
2 0 9
11 9 2 11 11 4 15 3 13 12 9 2
13 10 0 9 12 2 9 13 0 2 15 15 13 2
5 13 0 0 9 2
24 16 13 1 9 12 1 15 2 13 9 1 9 7 9 0 0 9 2 13 1 10 0 9 2
14 13 15 0 9 0 9 2 1 15 15 13 9 12 2
18 3 1 9 12 13 10 9 7 9 9 0 0 9 9 9 0 9 2
14 13 13 10 9 9 7 16 0 0 13 9 9 9 2
18 7 2 9 2 10 9 4 13 2 7 16 13 1 0 9 0 9 2
15 1 9 13 9 2 1 15 13 9 1 0 2 0 9 2
28 1 10 9 9 0 9 15 3 13 13 0 9 0 0 9 2 15 13 9 0 9 2 0 9 7 0 9 2
42 1 11 15 13 9 9 12 7 1 10 0 9 13 0 9 2 1 10 0 9 13 13 1 9 2 3 0 2 13 9 9 7 0 0 9 2 13 9 16 9 0 2
6 13 15 9 1 0 9
2 11 2
21 3 9 13 0 9 7 0 0 9 1 9 2 16 13 0 13 7 13 0 9 2
13 10 0 9 7 9 0 9 15 3 13 1 15 2
24 9 11 11 1 9 3 0 13 2 16 15 13 9 2 3 0 9 9 13 3 0 0 9 2
14 1 9 11 1 11 1 9 10 9 13 9 12 9 2
9 1 11 13 3 1 9 0 9 2
8 7 15 9 1 0 9 13 2
29 1 0 11 2 1 11 7 11 2 11 2 7 7 1 11 9 13 9 1 0 9 9 1 3 3 0 1 9 2
27 2 9 1 0 9 1 11 2 15 3 13 1 9 1 9 1 11 2 13 9 7 1 9 1 0 9 2
8 15 4 13 13 14 12 9 2
14 1 9 15 1 9 13 0 9 2 2 13 11 11 2
21 9 9 3 0 13 2 16 4 0 9 1 9 1 0 9 13 1 0 9 9 2
7 3 15 14 13 0 9 2
14 9 3 13 9 14 9 9 3 0 9 1 3 0 2
27 1 9 9 1 0 9 15 13 2 16 0 9 3 13 0 0 9 7 13 1 9 0 9 1 0 9 2
15 9 1 9 9 1 11 11 11 13 3 9 0 0 9 2
19 1 10 9 15 3 13 9 7 9 2 15 4 1 0 9 3 13 9 2
18 1 9 9 9 7 0 9 0 9 1 11 1 10 9 13 9 9 2
12 1 9 9 4 9 13 13 1 12 2 9 2
4 9 3 3 13
2 11 2
27 9 1 0 9 9 7 7 9 4 3 13 3 1 0 9 2 11 2 11 2 11 2 11 7 0 9 2
26 9 11 11 1 0 0 0 9 7 0 9 13 2 16 1 15 15 3 1 0 9 13 13 0 9 2
8 9 3 3 13 9 0 9 2
19 0 9 13 7 0 9 2 15 15 13 13 1 9 9 3 3 9 9 2
15 3 1 15 9 13 2 13 9 7 2 7 9 13 0 2
7 3 4 9 7 13 3 2
23 2 13 0 2 16 9 2 15 10 9 3 13 2 13 1 15 0 2 2 13 11 11 2
12 3 7 13 2 16 1 9 15 13 3 13 2
16 1 15 13 3 1 11 9 2 7 9 15 13 13 1 9 2
22 9 7 13 2 16 16 3 1 9 9 13 9 2 9 13 1 9 3 3 16 3 2
4 9 13 0 9
2 11 2
19 9 12 1 0 9 0 9 2 11 2 11 2 11 2 13 1 9 13 2
10 3 14 1 9 15 3 4 13 9 2
15 1 12 0 9 13 13 1 0 9 1 9 3 14 12 2
9 1 3 0 9 13 9 9 0 2
18 1 9 13 9 1 9 9 0 2 10 11 15 7 13 1 3 0 2
20 14 13 9 9 3 3 0 2 16 13 1 15 0 12 9 2 13 15 9 2
11 9 2 11 1 11 9 13 2 16 13 2
14 13 14 14 1 9 9 2 7 3 1 0 0 9 2
10 1 0 12 9 9 3 3 13 12 2
26 7 0 9 11 11 11 15 13 2 16 13 9 3 0 2 2 13 0 2 16 15 4 13 1 9 2
19 3 15 3 13 9 2 16 1 9 9 15 0 9 13 14 3 3 2 2
9 1 11 2 11 13 0 9 3 2
18 2 1 10 0 9 15 9 0 9 13 2 16 9 13 0 16 3 2
17 13 4 0 2 16 4 9 3 13 7 0 9 1 10 9 2 2
22 1 9 13 3 1 9 3 12 0 9 1 0 2 15 13 3 1 9 1 0 9 2
11 0 9 15 13 2 16 4 15 13 13 2
17 2 16 4 9 13 13 1 9 2 13 13 0 9 2 2 13 2
15 12 1 15 13 9 9 1 15 2 16 4 13 14 9 2
8 9 0 9 13 14 0 9 2
7 9 13 1 11 14 14 3
15 9 15 13 2 16 1 11 13 1 9 9 3 7 13 4
2 11 2
27 9 0 9 2 15 13 1 0 9 1 11 2 13 1 10 0 9 1 11 1 0 11 0 9 11 11 2
10 3 1 0 9 3 13 12 0 9 2
15 9 13 13 0 9 1 15 2 16 9 4 13 0 9 2
25 2 16 0 9 4 15 1 9 1 0 0 9 13 1 9 2 15 13 1 9 9 1 0 9 2
34 13 15 2 16 1 11 13 9 9 0 9 2 3 4 15 9 13 13 2 2 13 11 11 2 0 9 9 2 3 9 1 0 9 2
27 9 9 0 9 7 0 0 9 11 2 9 2 2 1 10 9 15 9 13 2 7 13 1 9 9 9 2
18 2 9 11 13 9 2 16 13 0 9 7 9 1 9 1 9 9 2
31 3 13 9 1 9 0 9 2 15 13 9 11 16 0 9 0 0 9 2 2 13 11 11 1 9 9 9 1 0 11 2
25 15 11 2 11 2 15 2 16 13 2 13 1 9 9 9 2 13 9 1 11 3 1 0 9 2
35 2 13 4 15 2 16 9 1 0 9 7 0 9 1 9 7 9 0 9 13 3 0 7 16 0 9 4 13 1 9 3 2 2 13 2
11 16 13 2 13 1 9 9 13 0 9 2
15 13 3 1 9 9 1 0 9 2 0 7 1 9 9 2
33 15 2 16 15 13 2 13 0 13 9 1 0 9 14 3 2 15 13 1 9 1 9 11 2 11 2 16 1 0 9 9 13 2
7 9 11 7 11 2 9 11
2 11 2
19 12 0 0 9 15 1 0 9 3 13 2 11 13 0 9 12 10 9 2
13 13 15 1 9 9 9 0 9 1 0 0 9 2
28 11 4 1 9 13 12 9 9 1 0 12 9 2 11 4 13 10 9 12 9 2 1 9 12 9 2 9 2
47 1 0 9 4 9 1 0 9 13 3 3 14 11 2 1 15 15 13 12 9 9 2 1 9 12 2 2 11 1 12 9 2 12 2 7 11 2 11 1 12 9 2 1 9 12 2 2
62 16 4 15 1 9 13 0 9 2 13 4 1 15 0 9 1 10 9 2 11 4 13 12 9 2 3 15 13 12 2 2 11 12 2 3 12 2 2 11 12 2 12 2 2 11 12 2 12 2 7 11 2 11 12 2 3 2 16 13 3 2 2
4 3 1 9 12
5 0 9 1 0 9
14 0 9 11 4 13 1 9 13 1 12 2 9 0 9
2 11 2
26 0 9 1 9 12 9 9 13 9 9 1 15 2 16 4 1 12 9 13 1 9 0 9 1 11 2
49 16 9 11 13 2 1 0 0 9 9 13 12 9 9 1 9 9 7 12 9 9 1 9 0 9 1 9 12 2 1 0 0 9 3 12 9 9 0 9 1 9 0 9 2 0 1 0 9 2
18 0 9 4 15 1 11 13 9 1 12 7 12 9 1 12 9 13 2
19 0 0 9 2 15 13 1 9 12 2 13 0 9 1 9 12 7 12 2
32 16 15 9 9 13 1 9 1 12 9 7 1 0 9 4 13 1 0 9 3 12 9 9 2 3 13 13 3 3 9 9 2
22 9 11 13 2 16 9 13 0 13 3 3 2 7 9 0 9 13 3 12 9 9 2
11 16 0 9 9 13 12 2 9 10 9 2
24 9 9 13 9 3 10 9 1 0 9 9 1 9 1 9 0 9 2 15 13 0 0 9 2
25 1 10 9 15 1 9 9 9 1 9 3 13 1 12 9 9 7 0 3 12 9 13 3 13 2
14 11 13 2 16 9 9 13 7 13 1 15 13 9 2
11 9 3 3 13 9 9 1 0 9 9 2
17 10 9 13 9 3 0 9 11 1 0 9 1 12 2 9 12 2
17 9 11 13 1 12 9 1 0 9 11 7 12 9 1 9 11 2
27 9 9 15 13 0 9 1 0 9 1 9 14 12 9 9 2 9 0 9 4 13 3 1 12 9 9 2
5 16 4 0 9 13
2 11 2
21 0 9 9 0 9 11 13 12 2 9 9 9 7 9 1 9 0 9 9 9 2
23 10 9 15 13 2 9 0 9 2 7 1 0 0 9 13 1 15 13 9 11 7 11 2
20 2 13 15 7 2 16 4 0 9 13 2 2 13 9 1 9 11 9 9 2
7 1 0 9 9 15 13 2
9 11 1 15 2 1 15 15 3 13
5 14 2 0 9 2
31 0 9 2 9 7 9 11 11 2 12 2 12 2 2 15 13 1 9 7 1 9 1 10 9 2 4 1 9 3 13 2
25 1 0 9 9 1 0 9 2 3 15 13 0 9 0 9 0 9 2 4 10 9 13 0 9 2
38 0 9 2 10 9 3 0 0 9 1 9 11 11 2 9 9 1 11 2 2 13 2 0 9 1 9 0 9 0 9 10 9 3 13 0 13 9 2
26 11 10 0 9 13 0 9 12 2 15 7 13 1 9 2 3 4 13 1 12 9 1 3 0 9 2
18 10 9 4 13 1 9 7 1 12 9 3 13 1 11 1 9 9 2
32 0 9 11 11 1 0 0 9 1 0 13 2 16 2 1 9 13 1 10 0 9 2 7 13 15 13 0 9 10 9 2 2
15 1 9 13 9 11 11 7 11 11 9 1 2 9 2 2
20 0 9 0 9 9 11 11 13 0 9 7 13 0 9 1 0 9 11 11 2
25 2 3 0 2 9 0 7 0 3 1 9 10 9 3 13 2 7 0 9 13 1 9 3 13 2
27 2 0 9 1 11 2 15 11 3 13 2 13 3 0 9 2 2 13 1 9 1 10 9 0 0 9 2
22 0 9 11 11 2 10 9 15 13 9 2 13 2 16 4 13 9 9 0 9 13 2
38 2 9 10 9 4 15 7 3 13 1 15 2 16 3 15 2 15 15 3 3 1 0 9 13 2 4 13 4 3 13 1 15 2 2 13 1 11 2
43 11 2 15 15 3 13 2 16 2 13 13 15 1 9 2 2 4 13 3 13 7 9 2 15 15 4 1 9 9 13 2 3 1 11 11 11 2 9 9 9 9 11 2
21 1 0 9 13 1 15 3 0 9 1 0 9 0 9 7 0 9 9 11 11 2
34 10 9 3 13 0 0 7 0 9 9 10 9 9 11 11 2 0 9 2 12 2 7 9 0 9 7 0 9 2 9 2 12 2 2
7 2 11 2 11 2 11 2
7 0 11 2 0 9 1 9
5 14 2 0 9 2
28 0 9 11 11 11 2 15 13 1 10 9 3 1 9 2 13 13 10 9 7 9 2 0 12 9 0 9 2
8 13 15 3 0 9 0 11 2
23 1 9 15 3 11 13 13 9 9 1 11 2 3 13 4 13 12 9 0 7 0 9 2
5 9 15 13 0 2
22 0 1 10 0 9 11 2 10 9 4 3 3 13 2 15 1 9 3 10 9 13 2
27 3 13 3 9 2 16 3 13 9 1 9 7 9 2 7 15 7 1 9 11 1 9 7 9 0 9 2
42 3 16 9 3 1 11 13 9 7 9 15 13 1 9 9 1 9 12 9 0 7 1 15 2 16 13 10 9 2 15 13 9 2 1 10 9 7 1 9 0 9 2
21 1 0 9 11 11 13 2 16 15 10 9 13 9 7 4 15 13 13 9 9 2
15 9 9 3 13 1 9 0 9 2 16 4 15 13 13 2
18 1 0 9 1 9 9 12 2 9 7 9 13 13 15 1 0 9 2
10 9 2 9 2 1 0 9 3 13 2
32 15 3 3 13 0 0 9 1 11 7 13 1 10 9 2 16 4 9 13 1 9 0 9 1 11 7 1 9 9 0 9 2
37 16 0 11 3 13 2 0 9 13 10 9 3 2 16 11 2 15 15 13 9 0 9 0 9 2 13 1 9 0 9 0 15 0 9 1 9 2
27 10 9 4 13 13 13 9 0 0 9 2 11 2 2 15 13 9 7 0 9 9 0 9 3 12 9 2
26 13 15 3 2 16 15 0 9 13 1 9 3 1 15 15 7 2 10 2 0 9 2 13 0 9 2
6 0 9 1 9 1 9
5 14 2 0 9 2
3 0 11 2
22 14 0 9 9 13 1 9 1 9 0 11 11 2 1 9 0 0 9 1 0 11 2
20 9 0 9 15 0 1 9 13 1 9 2 3 15 1 9 13 3 1 9 2
26 11 11 2 15 13 1 9 3 13 1 9 9 9 1 0 11 2 7 10 9 15 13 12 1 9 2
20 16 13 1 9 2 13 11 11 2 1 9 1 9 7 13 2 16 15 13 2
19 13 1 15 13 9 0 9 0 9 0 9 7 3 15 9 13 1 9 2
5 0 9 3 1 9
5 14 2 0 9 2
2 11 2
27 9 12 9 7 9 0 9 13 3 1 0 9 1 11 9 2 1 15 9 13 3 0 0 9 1 15 2
22 1 9 9 11 11 13 13 0 11 11 2 15 15 13 1 12 9 13 9 11 11 2
18 1 9 11 11 13 0 9 1 10 9 1 11 7 10 9 3 13 2
7 11 15 1 9 9 13 2
12 3 1 11 7 9 13 13 3 12 0 9 2
15 12 1 15 13 9 1 15 2 16 9 13 7 13 9 2
22 0 0 13 13 1 9 2 16 16 9 13 1 9 0 0 2 1 0 9 13 9 2
10 0 9 4 13 1 0 9 1 9 2
6 9 13 9 1 0 9
5 14 2 0 9 2
2 11 2
33 13 13 2 16 1 0 7 0 0 9 15 1 9 13 0 0 9 1 9 9 2 15 13 9 0 9 1 9 9 1 0 9 2
22 9 11 11 11 11 13 2 16 0 9 4 13 1 0 9 9 2 15 9 13 9 2
15 1 9 9 4 13 9 11 2 16 4 1 9 9 13 2
23 9 9 2 1 15 9 13 10 9 1 9 0 9 2 13 3 1 11 7 3 1 11 2
12 13 4 0 9 1 0 9 1 11 1 11 2
22 1 11 13 9 1 9 9 2 16 4 15 1 0 9 13 2 7 1 9 9 13 2
11 9 13 3 0 9 0 9 1 0 9 2
6 10 9 7 9 13 2
5 9 0 9 9 13
5 14 2 0 9 2
2 11 2
24 9 0 0 9 11 11 13 3 1 0 9 1 11 10 9 2 16 13 1 10 9 1 11 2
10 13 3 9 1 9 9 1 9 11 2
35 9 0 9 11 11 4 13 1 11 7 1 10 9 4 1 9 12 16 12 1 12 9 13 1 0 9 11 11 7 0 9 1 0 9 2
31 11 13 9 11 1 9 2 1 15 9 13 2 16 1 10 9 13 1 0 11 2 16 4 1 11 13 7 13 1 11 2
10 9 9 11 9 13 9 3 1 9 2
15 11 13 10 9 1 0 2 13 9 9 7 9 9 9 2
23 9 15 13 13 9 10 0 9 1 9 1 0 9 2 3 13 3 1 9 1 9 13 2
10 11 1 0 9 13 9 7 9 11 2
18 1 11 4 13 1 12 9 9 1 9 9 2 16 13 13 1 9 2
17 9 13 10 9 1 15 2 16 0 9 13 14 1 0 9 0 2
16 13 3 1 9 2 15 9 13 9 1 9 7 9 9 9 2
11 15 4 16 0 13 1 9 1 9 9 2
23 13 1 15 2 16 1 9 12 9 0 13 1 9 13 1 11 2 7 4 1 15 13 2
6 11 13 13 16 9 2
8 9 0 1 11 13 7 11 2
17 9 3 13 2 16 9 9 13 2 16 4 11 4 13 1 9 2
17 13 13 2 16 0 9 9 1 11 7 11 15 7 13 2 13 2
5 9 13 3 0 2
17 0 15 13 1 11 1 9 12 7 16 0 9 13 0 0 9 2
22 11 4 13 1 9 12 7 13 2 16 1 9 12 7 12 13 0 9 11 0 9 2
5 1 15 13 9 9
5 14 2 0 9 2
2 11 2
25 0 9 9 11 1 0 9 9 9 13 9 9 11 11 16 9 9 9 1 0 9 1 0 9 2
13 2 10 0 9 13 3 1 11 2 2 13 11 2
20 3 13 15 1 15 9 9 0 9 2 15 14 13 1 9 11 7 0 9 2
12 9 9 11 11 13 2 16 11 0 9 13 2
14 2 10 9 7 13 1 9 9 7 3 1 9 9 2
16 9 1 9 4 13 7 2 16 4 13 10 9 2 2 13 2
19 11 13 2 16 15 11 13 0 0 9 2 15 1 9 9 1 9 13 2
18 9 9 2 15 1 9 13 2 15 11 1 11 13 13 10 0 9 2
14 1 0 0 9 9 4 14 13 4 13 0 0 9 2
18 2 11 15 4 13 1 0 0 9 2 15 13 9 2 2 13 11 2
33 9 0 9 11 9 1 9 9 11 13 2 16 1 9 11 11 9 15 9 13 1 9 13 3 0 9 1 0 9 1 9 12 2
18 9 1 15 1 9 13 2 16 15 11 13 0 9 2 15 9 13 2
19 2 13 15 0 9 1 11 7 9 15 3 7 13 13 2 2 13 9 2
15 13 2 16 1 0 9 4 11 13 1 9 13 12 5 2
20 0 9 11 11 11 15 13 2 16 15 1 9 9 13 0 9 1 0 9 2
22 2 13 4 2 16 15 9 2 15 13 11 2 13 1 9 3 3 2 2 13 11 2
19 1 9 7 1 15 13 2 16 9 9 13 1 11 1 0 9 7 11 2
7 0 9 13 1 9 11 9
5 14 2 0 9 2
2 11 2
14 1 0 0 9 15 1 0 7 0 9 0 9 13 2
24 9 13 9 0 7 0 9 2 3 11 2 2 15 1 9 9 12 7 12 13 9 3 3 2
15 11 15 13 11 11 2 9 0 0 0 9 2 11 2 2
26 0 0 9 15 1 9 12 1 9 9 0 0 9 2 3 1 0 9 0 7 0 9 2 3 13 2
9 1 12 2 9 12 13 1 9 2
37 9 13 2 16 1 9 3 16 0 9 0 9 9 2 0 1 12 7 15 9 1 10 12 9 7 3 9 0 1 9 2 13 0 13 9 11 2
22 1 0 9 2 12 2 12 2 12 2 13 0 9 3 9 13 9 9 0 1 9 2
38 2 9 0 9 13 0 9 9 4 13 1 10 0 9 2 0 0 9 2 0 9 2 3 7 0 9 2 15 15 1 15 11 13 2 2 13 11 2
23 7 16 3 0 9 1 9 13 2 16 0 9 13 11 2 13 15 10 9 3 3 13 2
10 13 15 9 2 7 1 9 2 13 2
21 0 9 0 9 1 10 9 13 9 13 9 9 2 0 9 7 0 9 9 9 2
20 0 9 15 1 9 7 0 9 13 7 0 1 9 0 7 0 9 11 11 2
16 1 0 9 13 0 9 1 9 12 1 10 0 9 0 9 2
9 11 13 1 9 12 1 0 9 2
4 0 9 0 9
5 14 2 0 9 2
22 0 9 9 0 9 2 9 2 13 0 0 9 0 9 11 7 0 9 9 9 11 2
20 1 9 13 9 9 11 1 3 16 12 0 9 2 0 9 3 1 12 13 2
15 11 13 1 0 9 0 9 2 10 9 13 7 3 0 2
11 11 2 11 7 11 13 3 0 0 9 2
5 2 11 2 9 9
4 9 1 0 9
2 11 2
23 9 9 0 9 2 11 2 3 13 0 9 1 0 9 9 2 9 2 9 7 10 9 2
23 16 1 0 0 9 9 1 11 13 10 0 9 11 11 2 0 9 4 13 1 9 0 2
31 2 9 0 9 4 13 13 15 9 9 11 2 11 2 0 9 0 7 0 11 1 9 0 11 1 11 2 2 13 11 2
33 1 9 1 0 0 9 11 1 9 9 2 15 15 13 12 2 2 12 2 9 2 13 11 13 11 9 1 0 9 3 0 9 2
4 13 9 9 9
5 14 2 0 9 2
2 11 2
17 9 0 0 9 2 3 9 0 9 2 16 13 9 1 0 9 2
32 0 9 11 9 10 9 13 1 0 9 1 9 1 0 11 2 16 15 15 13 13 0 9 12 9 9 9 2 13 9 2 2
14 0 0 9 13 1 9 9 13 12 9 0 0 9 2
9 10 0 9 13 12 5 12 9 2
27 13 13 9 12 0 9 2 12 9 9 2 3 1 9 0 1 0 9 2 7 12 9 9 1 9 9 2
14 0 9 9 13 9 0 12 9 2 3 12 12 9 2
29 1 0 9 9 11 11 2 11 15 0 9 9 13 3 1 0 9 0 1 0 9 7 1 0 9 9 9 9 2
23 1 0 9 9 2 3 1 9 0 9 2 15 7 9 0 9 4 13 13 1 9 12 2
13 9 11 4 1 10 9 13 13 1 12 9 9 2
19 16 13 9 11 2 0 9 15 1 9 13 13 3 0 9 11 7 11 2
12 3 14 11 13 13 9 9 1 9 12 9 9
2 9 11
6 9 13 3 1 9 2
12 1 0 9 13 13 0 9 3 1 9 1 9
5 14 2 0 9 2
2 11 2
14 3 16 12 0 9 1 0 9 1 9 13 0 9 2
12 1 9 13 9 7 13 7 9 9 0 9 2
13 11 15 13 9 0 0 9 2 11 2 11 11 2
28 1 15 15 9 0 9 2 0 9 7 0 9 9 10 9 13 13 1 9 7 9 1 9 7 0 0 9 2
9 9 9 15 7 3 1 9 13 2
14 11 3 13 1 10 9 3 9 1 9 7 0 9 2
14 0 9 9 13 9 2 0 9 2 1 10 9 9 2
16 15 15 3 13 1 0 9 1 0 9 2 3 12 9 2 2
19 3 15 7 13 9 2 15 15 13 9 3 1 9 3 1 9 1 9 2
31 1 3 0 9 13 3 0 9 2 0 9 12 2 11 1 9 2 0 9 2 0 9 2 9 7 3 10 0 0 9 2
16 9 15 13 1 9 3 1 11 7 1 0 0 9 1 11 2
15 1 0 9 0 9 13 0 0 9 1 9 3 0 11 2
12 3 15 14 3 13 9 0 9 1 0 9 2
18 13 15 3 3 11 7 1 9 11 7 9 1 10 9 13 1 11 2
24 9 15 13 1 11 7 2 16 1 11 2 3 16 1 0 0 9 2 13 0 9 0 9 2
12 1 11 13 1 0 0 0 9 10 12 9 2
22 1 11 13 10 0 9 3 11 2 16 1 10 9 13 9 0 9 0 0 0 9 2
19 3 1 10 9 0 9 3 13 7 13 2 3 15 1 9 13 0 9 2
28 0 9 13 1 10 9 1 9 0 9 2 7 13 1 15 3 16 3 2 11 2 3 9 13 12 12 9 2
10 9 1 9 9 13 1 9 1 9 9
5 14 2 0 9 2
2 11 2
30 0 9 9 11 11 2 11 2 7 11 11 2 11 2 11 2 3 13 0 9 0 0 9 1 9 0 7 0 9 2
42 9 13 9 3 2 16 13 10 9 2 16 4 15 1 9 1 0 9 1 9 9 2 9 9 1 9 7 0 2 0 0 9 2 13 14 3 2 3 3 3 3 2
22 9 9 11 11 2 13 2 7 1 10 9 9 13 2 16 13 15 4 3 14 3 2
22 2 9 9 10 9 1 9 1 15 13 3 0 9 2 2 13 11 0 7 0 9 2
10 9 13 13 2 13 7 9 0 9 2
22 9 15 3 13 13 7 1 9 0 9 11 1 9 1 9 2 15 4 13 0 9 2
21 2 9 9 9 13 1 9 1 9 2 16 1 15 13 3 13 2 2 13 11 2
34 9 11 13 2 16 1 0 9 9 9 13 9 2 16 4 15 13 0 9 0 13 9 9 1 0 9 7 9 9 1 0 9 9 2
5 9 7 9 13 2
13 11 15 9 13 2 1 9 1 9 13 0 9 2
7 1 9 13 12 9 9 2
5 14 2 0 9 2
3 0 11 2
24 0 9 13 11 0 11 2 15 13 0 9 0 9 2 1 0 9 1 9 14 12 9 9 2
22 1 0 0 9 2 1 15 13 0 9 11 2 11 2 13 9 1 9 12 9 9 2
21 16 13 2 4 9 9 13 9 9 9 1 9 12 1 0 9 3 12 9 9 2
10 0 9 13 9 9 7 1 0 9 2
21 1 9 12 13 9 1 12 9 1 9 12 9 7 10 0 9 13 12 9 9 2
13 9 9 13 3 12 9 9 7 9 12 9 9 2
12 9 13 12 9 9 7 9 9 12 9 9 2
23 3 2 3 16 9 2 15 1 15 13 0 9 2 13 9 2 9 2 9 7 0 9 2
15 3 12 9 9 13 9 2 1 15 13 12 9 1 11 2
16 0 9 15 1 9 12 13 1 12 9 7 13 3 12 9 2
30 1 9 0 9 1 12 9 9 15 1 11 13 3 9 2 16 1 9 12 11 13 0 9 9 1 0 9 0 9 2
10 9 0 1 0 0 9 13 12 9 2
8 3 13 0 9 9 0 9 2
20 9 11 10 9 13 7 3 15 13 11 1 12 9 7 9 11 1 12 9 2
24 0 9 13 1 12 9 11 2 16 9 0 9 2 15 13 12 9 9 2 3 12 9 13 2
7 9 13 13 12 9 9 2
14 7 9 9 15 3 13 2 16 15 10 9 3 3 13
7 9 9 3 3 13 3 0
8 3 3 0 9 13 1 0 9
6 0 9 1 0 9 13
3 9 3 13
26 9 9 1 0 2 15 15 10 0 9 13 1 0 9 13 9 0 9 2 3 3 13 2 15 13 2
15 9 7 9 3 13 0 9 2 9 7 3 3 0 9 2
18 3 16 0 9 9 13 9 9 10 9 7 0 9 9 7 2 9 2
23 1 9 13 0 9 1 9 0 9 2 1 0 9 3 2 14 1 9 12 7 12 9 2
12 9 3 0 9 3 13 1 12 7 12 9 2
18 1 0 9 3 0 9 2 3 15 3 2 1 9 2 0 9 13 2
31 16 1 9 0 9 4 13 14 12 9 9 1 9 7 14 12 9 1 0 9 2 3 3 13 10 9 3 12 1 12 2
15 2 13 2 10 9 13 2 16 9 9 15 13 12 9 2
27 1 9 14 1 9 13 7 9 13 14 1 9 2 2 13 1 0 9 12 1 0 9 2 15 4 13 2
7 13 9 7 13 4 13 2
6 9 3 2 13 2 2
19 13 2 16 15 13 10 9 7 9 9 1 2 9 2 16 3 15 13 2
18 2 9 2 9 2 9 2 9 2 13 15 3 7 13 15 1 9 2
17 15 15 13 2 15 15 15 13 2 7 7 0 9 15 13 2 2
27 1 0 0 9 3 1 10 9 13 1 0 9 12 0 9 1 0 7 1 10 9 13 7 0 0 9 2
13 2 13 15 3 13 7 1 0 9 2 2 13 2
18 0 9 9 1 0 9 4 1 0 9 13 1 3 16 12 9 9 2
24 1 15 1 9 4 13 4 13 3 12 9 9 2 1 0 9 12 9 7 9 13 0 9 2
15 1 9 4 15 3 1 9 9 13 13 14 12 9 9 2
42 9 3 13 1 12 2 7 16 15 9 9 1 0 3 3 13 1 9 7 1 10 0 9 3 13 0 9 9 2 9 1 3 0 9 15 13 3 16 1 0 9 2
12 9 0 9 13 3 3 0 16 9 0 9 2
12 1 0 9 7 7 15 3 2 7 3 13 2
29 1 9 0 9 4 1 0 9 13 3 12 9 0 0 9 2 15 13 1 12 9 3 16 1 0 9 9 12 2
15 1 0 9 3 13 13 1 11 2 9 9 7 11 9 2
19 16 15 13 3 3 2 13 3 0 9 9 3 9 3 12 9 0 9 2
34 1 0 9 1 9 15 3 3 1 9 7 1 9 1 9 13 1 12 1 12 9 1 9 2 1 0 9 12 7 12 9 1 9 2
23 0 9 0 9 15 1 0 9 1 9 1 9 12 3 13 7 3 15 3 13 7 3 2
17 0 7 0 9 14 13 1 0 3 0 9 9 16 0 0 9 2
14 0 9 13 1 9 2 16 15 1 15 13 3 13 2
16 7 16 15 14 15 13 2 16 1 12 9 13 3 1 9 2
9 1 9 15 3 13 0 9 9 2
26 15 13 9 9 7 9 2 13 3 3 9 1 15 2 15 3 15 7 10 9 13 9 13 1 0 2
9 9 0 9 9 7 9 3 13 2
12 1 0 9 15 14 3 13 9 9 0 9 2
6 11 13 13 0 0 9
2 11 2
18 9 0 9 1 0 9 7 9 1 0 9 7 1 9 0 9 13 2
23 10 9 13 1 3 0 0 9 0 9 1 11 11 11 2 11 1 12 0 0 9 11 2
19 9 0 0 9 13 0 9 0 9 7 0 9 0 9 13 1 0 9 2
14 1 0 9 13 1 0 9 0 9 0 0 9 0 2
15 11 3 13 0 9 2 15 4 3 13 13 7 10 9 2
23 9 13 1 9 3 12 0 0 9 2 15 4 13 4 13 0 9 2 13 11 2 11 2
17 0 9 1 0 9 13 3 3 12 9 9 7 9 12 9 9 2
16 1 9 0 9 1 11 15 3 12 9 13 9 7 0 9 2
16 0 9 1 0 9 7 9 1 0 9 13 1 9 0 9 2
19 1 0 0 9 11 1 11 11 11 2 11 13 3 9 0 9 12 9 9
5 9 7 9 13 0
10 3 0 9 4 1 9 0 9 13 3
28 11 11 1 0 9 13 9 0 9 2 16 13 3 1 9 9 1 9 0 7 0 9 3 9 9 1 9 2
19 3 1 9 9 13 1 9 0 9 2 0 0 9 7 1 9 0 9 2
19 1 9 1 9 11 11 11 11 13 0 9 1 9 0 9 12 9 9 2
34 0 9 9 1 0 9 7 13 1 12 9 1 12 9 7 9 1 0 9 15 13 1 12 9 1 0 7 1 12 9 1 0 9 2
19 0 9 0 9 1 12 9 1 0 9 15 3 13 1 12 1 12 9 2
25 1 0 9 13 1 0 9 9 0 9 1 12 1 12 9 7 9 9 1 9 0 9 0 3 2
17 1 9 1 0 9 13 0 9 12 9 7 1 0 9 12 9 2
18 3 7 4 13 0 9 0 7 0 9 3 1 9 0 1 0 9 2
38 9 1 9 9 9 1 9 15 13 1 0 12 9 1 9 7 12 9 1 9 1 0 12 9 7 0 9 1 9 9 1 0 12 9 1 12 9 2
19 1 3 0 9 13 1 9 9 1 9 0 9 7 4 13 1 0 9 2
35 1 9 11 4 11 11 7 3 13 1 9 10 0 9 0 9 1 15 0 9 0 1 9 0 12 0 9 1 9 12 9 1 12 9 2
21 9 0 9 15 13 1 9 1 12 9 1 0 7 1 12 7 12 9 1 0 2
26 3 1 0 0 9 13 1 9 9 9 3 1 12 9 2 3 1 9 0 11 2 11 2 7 11 2
6 0 9 13 1 11 9
2 11 2
25 0 9 1 11 3 13 2 16 0 9 13 1 9 12 7 12 0 9 1 0 9 12 9 9 2
12 13 15 1 9 0 0 0 9 2 11 2 2
33 1 0 9 4 9 13 12 9 9 2 1 0 9 12 9 9 2 1 9 12 15 13 12 9 9 7 1 9 12 12 9 9 2
12 13 15 4 3 9 9 7 9 9 7 9 2
4 11 13 0 9
2 11 2
9 0 0 9 13 9 7 0 9 2
17 9 1 15 13 9 0 0 9 2 1 15 13 13 3 1 9 2
8 13 15 3 0 9 1 11 2
21 0 9 9 2 15 4 13 1 9 0 9 1 0 9 2 15 13 13 3 3 2
8 3 15 3 13 1 10 9 2
32 9 2 15 13 13 7 0 2 4 13 13 3 12 7 12 9 9 2 7 1 9 10 0 9 15 4 13 13 7 0 9 2
9 10 9 7 4 13 1 9 9 2
29 1 0 0 9 13 1 0 9 12 9 2 15 13 12 9 0 0 9 7 13 0 9 1 9 14 12 9 9 2
10 12 12 0 0 9 13 1 0 9 2
11 0 9 15 1 0 0 9 11 13 12 9
6 1 9 14 1 11 2
8 11 2 11 2 11 11 2 2
28 9 11 7 11 13 0 9 0 9 1 11 1 0 11 2 3 15 13 13 1 11 1 9 9 1 0 9 2
26 1 11 4 13 1 9 1 11 2 3 15 13 1 9 11 2 15 15 1 12 9 13 1 9 11 2
10 11 13 0 0 9 7 11 0 9 2
18 9 15 14 13 1 9 7 13 15 4 1 9 2 15 13 1 15 2
15 13 14 12 9 1 9 2 12 0 9 7 12 0 9 2
13 11 13 7 9 9 2 16 11 13 9 9 9 2
19 1 9 11 13 4 2 13 3 1 0 9 11 1 11 2 3 13 9 2
7 1 9 13 0 0 9 2
23 13 15 1 0 0 9 7 10 9 2 15 13 13 7 9 11 11 11 2 7 9 11 2
23 12 9 13 9 11 1 9 10 9 2 7 3 13 15 14 3 7 15 0 15 7 13 2
17 13 2 16 9 4 13 13 7 9 11 7 9 10 0 9 11 2
16 2 15 3 15 1 11 13 2 2 13 1 9 1 11 11 2
7 0 9 11 13 14 9 9
5 14 2 0 9 2
2 11 2
23 0 0 9 0 9 0 0 9 2 0 2 9 2 11 2 11 11 13 1 10 9 13 2
7 13 1 15 3 0 9 2
22 1 9 9 3 4 3 13 2 16 9 13 9 7 9 2 7 13 15 3 0 9 2
36 11 4 3 1 0 9 11 11 13 1 9 1 9 12 9 9 2 15 13 1 9 1 0 9 7 9 15 13 1 9 1 9 12 9 9 2
10 0 9 9 15 13 1 12 9 9 2
19 9 13 9 1 11 11 2 15 13 9 0 9 9 0 2 9 2 11 2
34 1 9 0 9 15 7 1 11 13 2 16 3 2 16 1 9 1 11 13 15 0 9 0 2 9 2 11 2 1 9 9 9 13 2
15 9 9 11 11 7 9 11 11 11 13 9 11 1 0 2
7 11 13 9 9 1 9 2
26 9 3 7 3 13 0 2 9 2 11 2 7 12 9 3 9 13 11 2 15 13 0 9 10 9 2
25 16 0 2 9 2 11 9 13 2 13 11 1 11 0 9 1 9 9 1 9 9 9 11 11 2
20 9 3 11 3 13 0 2 9 2 11 2 0 9 2 1 15 13 0 9 2
42 9 9 2 10 13 9 0 2 9 2 11 2 12 2 9 12 13 1 0 9 0 2 9 2 11 2 0 9 9 1 9 9 1 9 9 9 2 15 13 13 3 2
20 9 9 9 9 11 11 11 3 13 2 16 9 1 9 9 3 13 10 9 2
8 15 13 1 0 9 2 2 2
10 9 1 9 1 9 9 0 12 2 2
22 3 15 13 9 1 10 9 3 3 1 12 9 2 3 3 4 13 2 9 0 2 2
54 1 10 9 15 2 3 2 15 13 2 9 9 13 7 1 0 9 2 9 9 15 13 3 3 9 2 13 9 2 15 13 1 15 2 16 4 9 15 2 15 13 9 9 9 7 3 15 13 2 4 1 15 13 2
11 1 9 10 9 15 15 13 3 3 3 2
9 3 4 13 9 2 15 13 0 2
14 9 9 1 9 13 9 2 15 15 15 13 1 9 2
12 9 2 13 1 10 9 2 15 13 1 9 2
18 9 1 0 9 15 15 13 13 2 7 16 15 13 2 13 15 9 2
12 9 13 7 13 15 1 9 1 9 9 10 2
39 13 3 2 13 9 9 2 7 0 9 2 9 3 3 9 13 2 13 9 9 1 9 2 3 15 3 1 12 9 13 13 1 10 3 3 0 9 2 2
7 10 9 1 9 13 9 2
16 13 15 7 9 2 1 15 15 13 10 9 1 10 0 9 2
8 9 13 9 2 16 13 3 2
20 16 4 9 13 2 13 13 1 0 9 1 9 2 1 0 15 13 3 13 2
11 16 4 15 9 1 9 13 2 15 13 2
3 0 9 2
5 16 4 4 13 2
6 9 14 1 9 0 2
10 1 0 9 9 3 13 1 9 9 2
7 9 13 2 16 13 9 2
34 3 15 13 0 9 2 16 15 15 13 1 0 9 2 13 9 7 9 7 13 0 9 2 15 3 13 1 9 0 2 15 9 13 2
29 15 15 13 1 0 2 15 13 2 9 1 12 11 2 13 2 16 0 13 9 2 16 4 4 13 2 14 13 2
11 4 2 14 3 13 2 3 15 15 13 2
19 15 2 15 15 13 2 15 3 15 13 2 16 15 3 13 7 9 13 2
29 3 0 15 13 13 1 9 7 3 13 1 15 2 16 4 13 9 2 16 15 13 9 14 13 2 7 3 13 2
47 13 1 9 9 1 15 2 15 13 1 0 9 2 7 1 15 2 15 1 9 15 15 2 15 3 13 2 15 13 9 9 1 10 9 7 1 10 9 3 13 2 1 15 4 9 13 2
12 13 7 0 9 2 16 9 7 9 3 13 2
37 4 2 14 10 9 9 1 10 9 13 2 4 2 14 13 3 9 1 9 1 9 16 1 9 0 9 2 13 15 3 0 9 13 0 16 13 2
25 2 1 12 12 9 13 9 2 9 2 9 1 9 2 2 13 9 9 9 11 11 2 12 2 2
29 10 0 9 1 9 0 9 7 0 9 13 1 9 1 12 2 9 9 1 9 9 1 0 9 9 1 0 9 2
8 11 0 1 9 9 4 13 9
3 11 11 2
28 11 11 11 2 12 2 2 0 3 2 1 9 12 0 9 9 11 2 13 3 0 9 1 9 0 9 9 2
22 1 0 9 4 13 1 9 9 9 1 12 9 2 7 10 9 3 3 13 1 9 2
22 1 9 12 4 1 0 9 1 11 13 1 9 9 2 16 12 1 15 4 3 13 2
11 11 15 1 9 13 2 3 7 9 13 2
15 13 2 16 15 9 13 9 10 9 2 7 7 13 9 2
12 0 9 4 13 12 2 9 16 9 1 0 2
10 11 4 1 0 0 9 13 1 9 2
15 3 1 9 4 1 15 13 9 2 7 13 15 15 13 2
18 1 9 0 9 4 13 10 9 2 16 1 9 13 0 9 10 9 2
30 9 13 2 16 3 9 11 4 4 0 1 10 9 2 15 0 9 13 2 13 1 9 2 13 1 9 9 7 13 2
13 10 9 3 13 2 16 1 9 13 3 0 9 2
6 9 4 3 3 13 2
8 9 9 0 11 13 2 13 11
2 11 2
27 9 9 7 9 3 13 2 16 4 9 11 11 11 4 13 9 1 9 0 0 9 11 2 3 11 2 2
12 13 15 9 11 11 1 0 0 9 1 11 2
51 2 0 9 2 15 4 1 10 9 13 2 13 15 2 16 4 9 4 13 3 3 2 2 13 9 11 1 9 11 1 9 0 1 12 9 2 16 1 15 13 4 13 9 11 2 15 13 0 0 9 2
36 1 9 11 2 16 13 4 11 13 11 1 0 9 1 9 9 9 2 9 13 2 16 15 3 13 1 9 9 9 2 15 13 9 9 11 2
23 1 15 13 13 1 9 2 16 4 15 9 11 11 13 1 9 9 9 7 9 0 9 2
17 11 13 2 16 15 3 13 2 3 4 11 13 1 12 9 9 2
39 2 13 15 9 2 7 13 4 1 9 2 16 15 13 1 9 11 2 7 13 9 2 15 13 13 13 9 9 11 7 3 1 10 0 9 13 7 9 2
24 16 4 15 3 13 2 13 4 0 9 7 11 4 13 3 3 16 3 2 2 13 9 11 2
22 9 9 3 13 11 9 2 1 15 15 13 1 0 9 0 9 2 9 13 9 2 2
7 9 14 3 10 9 13 2
36 1 9 4 9 0 9 1 9 2 3 0 9 9 13 1 9 2 13 1 9 9 0 9 9 9 2 9 9 7 9 0 9 7 0 9 2
29 2 9 9 1 10 9 13 7 0 7 0 9 1 9 9 11 1 0 16 3 0 9 2 2 13 15 1 9 2
7 0 9 11 13 14 9 9
11 2 9 2 1 0 11 3 13 3 12 9
10 0 9 2 1 9 0 9 1 9 2
12 1 12 9 0 9 0 9 2 1 0 9 2
15 9 2 9 7 9 2 0 3 1 15 2 13 15 9 2
13 0 9 13 9 9 2 3 9 13 9 1 9 2
12 14 1 9 13 9 11 1 9 1 0 9 2
19 2 3 13 15 0 2 7 16 13 2 13 4 1 9 2 2 13 15 2
2 9 2
21 9 2 15 13 9 7 9 13 13 9 9 2 13 1 0 11 1 9 0 9 2
9 9 0 9 13 9 9 9 9 2
28 9 12 0 2 9 2 0 3 0 9 7 0 9 2 0 0 9 1 9 2 9 1 9 2 13 1 9 2
42 2 12 9 13 3 9 2 2 13 3 3 3 0 9 11 11 7 13 15 2 16 3 1 9 15 1 2 9 2 2 3 15 9 1 0 9 13 2 13 0 9 2
23 0 9 13 9 0 9 11 11 2 2 9 13 13 3 12 2 7 3 9 1 9 2 2
20 2 13 3 3 15 2 2 13 11 11 7 13 15 1 9 9 1 0 9 2
14 0 9 13 1 9 2 9 13 9 7 13 10 9 2
28 2 9 1 9 13 1 9 1 9 2 13 3 13 2 2 3 13 9 2 2 1 12 9 13 15 6 0 2
23 15 4 3 13 7 15 15 13 2 16 1 9 9 13 9 2 7 13 15 2 2 13 2
16 10 9 13 7 9 11 2 2 9 3 13 2 13 7 0 2
4 9 13 2 2
21 7 3 13 2 2 3 2 15 13 9 13 9 1 15 2 16 15 3 13 2 2
2 0 9
12 11 11 0 9 13 14 0 14 3 1 9 2
11 1 0 9 11 11 1 11 9 13 3 2
41 1 9 0 9 1 9 7 0 9 9 13 1 0 9 2 16 1 3 16 0 9 2 1 9 2 7 7 3 13 9 2 15 13 10 0 0 9 1 9 12 2
42 0 0 9 2 1 15 13 11 9 1 9 1 11 2 15 15 13 14 0 9 2 7 13 15 15 3 2 16 9 1 9 3 13 1 9 9 2 3 13 14 15 2
7 9 9 7 3 15 13 2
30 12 9 1 15 13 14 9 2 1 15 10 9 13 7 13 2 16 2 2 2 2 1 9 13 13 10 0 9 2 2
17 15 3 13 9 0 9 2 16 4 9 0 9 13 9 0 9 2
23 13 4 15 13 2 16 9 1 9 9 9 7 2 9 2 13 1 9 3 3 13 9 2
13 9 13 3 3 0 9 7 13 7 1 9 9 2
34 0 9 3 1 0 9 4 3 3 13 9 2 1 0 9 15 13 10 0 9 13 9 7 12 9 3 9 13 2 10 3 13 9 2
6 0 9 15 13 0 9
15 11 15 1 9 1 11 13 9 9 11 12 1 9 0 11
4 11 2 11 2
37 0 7 0 0 9 13 3 9 9 2 15 9 0 0 0 9 2 14 12 1 12 9 9 2 13 1 9 3 9 0 0 0 9 11 2 11 2
31 1 12 9 4 13 7 1 9 13 12 0 2 9 2 2 15 13 9 7 9 7 13 15 13 1 0 9 1 0 9 2
22 12 9 13 1 9 1 9 2 16 13 1 9 2 7 10 9 3 13 1 9 9 2
26 9 9 11 11 11 2 15 15 3 13 9 13 7 14 1 9 13 9 2 9 13 2 2 13 13 2
17 1 15 2 15 15 13 1 11 2 15 1 12 9 11 13 9 2
12 3 13 3 3 2 3 4 13 2 2 2 2
19 9 0 9 13 3 0 9 1 0 9 0 9 1 9 11 12 1 11 2
16 2 16 4 1 9 9 13 13 2 13 4 15 9 1 9 2
38 13 3 0 2 1 9 0 9 7 9 15 0 9 2 15 15 1 15 3 1 0 9 13 2 9 13 2 2 13 11 11 2 0 9 0 0 9 2
10 0 9 9 11 11 13 14 0 9 2
11 2 1 0 9 1 11 13 0 9 2 2
14 9 9 13 0 9 9 11 11 7 13 7 0 9 2
7 3 1 9 13 0 9 2
6 2 9 2 3 9 2
18 1 9 11 13 0 9 0 9 15 13 0 9 2 2 13 0 11 2
42 2 16 4 0 0 9 13 1 9 2 16 11 13 0 9 1 9 9 1 9 1 0 9 2 3 3 4 13 15 2 1 15 15 1 11 13 2 2 13 0 9 2
26 0 9 2 2 0 9 15 13 0 9 2 16 13 1 9 0 9 2 16 4 13 7 10 0 9 2
28 1 9 11 4 0 0 9 13 11 0 9 2 16 4 13 10 9 1 9 11 2 15 15 11 3 13 13 2
14 0 9 13 1 10 9 13 15 1 0 9 0 9 2
13 2 0 9 13 10 0 9 9 1 9 0 9 2
9 10 9 1 9 10 0 9 13 2
15 9 1 0 9 13 15 13 2 13 15 9 7 13 9 2
14 13 7 0 9 11 7 10 9 2 2 13 11 9 2
20 0 0 9 2 11 2 13 0 9 1 9 16 1 0 2 7 7 0 9 2
14 2 13 15 0 9 11 7 0 9 9 12 1 11 2
22 3 16 15 12 9 13 2 13 11 0 9 1 9 0 9 2 2 13 0 9 11 2
12 9 1 11 13 7 0 0 9 2 11 2 2
12 10 9 11 11 7 13 1 9 9 9 12 2
17 2 0 9 11 12 4 13 13 1 11 7 1 9 0 1 11 2
7 15 15 13 13 9 2 2
3 1 0 9
24 11 11 13 1 0 9 1 9 11 11 1 9 9 11 11 2 15 3 13 14 0 12 9 2
5 9 1 9 3 13
13 0 9 9 11 2 9 1 11 0 1 12 2 9
2 11 2
6 10 9 4 13 3 2
39 1 10 9 13 7 9 0 9 0 9 2 9 2 11 1 9 0 9 11 11 7 11 9 1 9 7 0 9 9 0 9 0 12 2 9 12 1 9 2
6 9 4 1 9 13 2
17 13 15 3 9 11 2 16 9 1 9 13 4 13 1 0 9 2
16 0 9 0 9 13 3 1 15 0 9 2 13 0 11 2 2
38 12 9 13 14 0 9 2 1 15 3 2 13 2 16 2 2 2 2 1 9 13 13 10 0 9 2 7 1 9 15 3 16 0 9 11 11 13 2
33 16 0 9 0 9 11 11 11 13 2 16 9 1 9 13 9 2 7 1 9 9 13 13 3 0 9 2 9 9 15 13 13 2
37 2 1 1 9 9 7 1 9 1 9 11 1 9 9 9 9 7 11 1 15 9 0 9 11 9 9 13 2 2 13 1 9 9 9 11 11 2
18 1 10 9 4 13 0 9 1 9 9 9 14 1 9 9 0 9 2
17 0 9 13 0 2 9 9 1 11 13 14 12 2 9 1 9 2
22 9 7 3 1 9 13 9 2 13 3 1 0 11 7 0 9 3 1 0 9 13 2
4 9 13 1 9
8 11 11 0 9 9 1 12 9
2 11 2
34 0 11 11 11 13 0 9 1 9 7 1 9 13 1 12 9 3 16 11 11 2 15 15 13 9 1 9 1 12 9 1 9 9 2
12 0 9 1 11 13 11 2 15 3 13 3 2
5 15 15 13 9 2
7 11 11 13 13 3 0 2
23 12 9 9 15 13 14 1 0 9 2 16 16 0 13 12 9 9 1 9 1 12 9 2
16 0 1 0 9 13 1 9 11 11 2 15 13 12 2 9 2
21 1 12 0 0 0 9 13 1 12 0 7 1 9 3 13 13 1 9 11 11 2
22 3 0 0 9 15 13 11 11 2 7 12 9 1 9 15 13 14 1 12 2 9 2
22 16 11 13 9 1 0 9 3 7 0 9 3 2 13 11 1 12 9 3 0 9 2
10 9 9 1 12 9 13 11 11 11 2
16 1 9 9 11 7 0 9 1 9 1 11 13 0 0 9 2
17 9 9 11 11 1 11 13 1 12 9 1 9 14 1 0 9 2
14 0 9 0 9 13 10 0 9 0 2 12 2 2 2
3 9 9 11
2 11 2
19 9 11 11 15 13 13 0 0 9 1 11 2 0 1 0 9 1 11 2
14 1 10 9 11 11 13 9 3 0 9 1 0 9 2
4 9 1 12 9
2 11 2
23 9 0 9 0 9 2 0 0 12 15 1 11 13 1 0 9 11 0 7 10 9 11 2
27 1 0 0 9 4 13 11 7 11 2 1 9 13 1 0 9 9 1 9 1 11 11 2 11 7 11 2
2 0 9
4 11 2 11 2
12 0 0 9 9 13 10 0 9 1 0 9 2
29 9 9 11 13 1 9 9 11 0 9 11 11 12 2 12 2 7 1 1 9 12 2 12 1 0 9 4 13 2
34 9 9 11 11 13 1 9 9 11 7 1 0 9 1 0 9 11 11 12 2 12 2 0 9 12 2 12 2 2 1 0 9 13 2
2 0 9
2 11 2
24 0 9 4 13 1 0 0 9 2 11 2 11 2 11 2 11 2 7 9 0 11 7 11 2
6 9 1 11 3 13 2
6 0 9 13 3 13 2
3 11 1 11
8 9 7 12 9 11 11 1 11
5 11 2 0 11 2
18 9 0 11 11 11 13 10 0 9 11 11 1 11 11 1 11 11 2
16 0 9 4 1 11 13 7 0 9 9 1 0 9 11 11 2
17 0 0 9 11 1 12 9 0 9 13 12 9 7 13 12 9 2
10 1 11 13 1 9 12 1 11 11 2
10 1 0 9 13 1 12 9 12 9 2
20 3 13 0 9 1 11 7 1 0 12 9 13 12 9 7 1 0 12 13 2
16 11 1 10 12 9 11 3 13 3 12 9 7 1 12 13 2
20 3 0 0 9 13 9 11 11 2 15 13 1 0 9 11 11 12 2 12 2
12 0 9 1 10 9 13 11 11 7 11 11 2
30 11 13 9 11 11 3 2 16 1 0 12 9 15 13 9 11 2 15 15 1 12 2 9 13 0 9 9 10 9 2
14 11 11 13 1 0 9 1 0 11 11 12 2 12 2
15 0 9 11 11 13 0 9 14 1 12 2 9 0 9 2
17 3 13 11 7 12 9 1 0 9 13 1 9 9 0 9 11 2
14 3 1 9 0 11 2 11 12 2 12 13 0 9 2
30 0 9 13 1 12 2 9 11 11 2 3 15 13 3 2 2 13 7 14 1 9 9 1 12 2 12 1 9 11 2
11 3 1 0 12 13 0 9 11 11 11 2
3 11 1 9
3 0 11 2
12 11 11 11 13 0 9 9 9 1 9 11 2
27 0 9 13 1 12 9 1 0 9 1 0 0 11 1 11 11 11 2 15 1 0 9 13 0 12 9 2
11 9 9 11 2 11 13 12 2 12 9 2
7 11 13 0 9 0 9 2
19 9 0 9 1 11 11 1 11 7 9 11 11 13 3 12 2 12 9 2
8 0 9 4 1 12 9 13 2
3 11 1 11
2 11 2
18 0 9 7 9 9 11 11 11 15 3 1 9 0 9 0 9 13 2
16 3 3 13 1 11 2 3 13 1 9 1 9 0 9 11 2
17 13 1 9 2 16 3 1 10 9 4 13 3 1 0 11 11 2
5 11 13 1 0 9
9 9 9 1 0 9 13 9 3 13
10 9 9 0 9 13 9 1 9 0 2
40 0 9 3 13 1 15 2 16 0 9 13 0 13 9 14 1 12 9 0 9 2 7 3 15 3 1 0 9 13 9 0 9 1 9 1 9 1 9 11 2
21 1 9 0 9 13 9 7 15 7 0 9 2 7 0 9 1 9 13 3 0 2
30 0 9 2 13 2 14 13 2 16 1 9 9 13 9 10 9 1 3 0 9 2 13 3 3 13 9 1 0 9 2
34 15 3 11 2 0 1 10 0 9 2 13 1 15 3 2 16 3 13 0 9 3 1 9 7 9 1 0 9 3 13 1 9 0 2
17 1 0 9 15 3 13 13 13 1 11 7 0 9 3 1 11 2
11 9 9 4 7 7 1 10 9 3 13 2
15 9 1 0 9 13 0 9 3 3 1 9 1 0 9 2
18 9 13 1 0 9 1 0 11 11 3 11 2 15 9 13 12 9 2
41 1 0 13 1 0 9 0 0 9 1 10 11 13 2 3 1 11 2 1 0 9 2 7 3 1 9 13 13 15 1 11 13 3 7 12 9 3 1 9 13 2
18 9 0 9 9 11 11 13 13 12 2 9 1 11 1 9 1 11 2
19 3 13 1 11 2 11 7 11 2 1 0 9 11 7 11 13 13 9 2
28 9 11 2 11 2 11 2 11 4 13 1 9 1 10 9 2 11 4 1 9 0 9 13 7 13 3 0 2
14 9 0 9 13 16 0 9 0 9 9 0 9 9 2
24 1 0 9 1 11 2 12 2 12 2 1 11 2 3 13 15 1 9 11 2 11 2 11 2
35 16 15 13 15 0 2 13 1 9 9 11 7 1 15 15 4 13 12 9 2 15 1 0 9 13 1 9 11 2 11 2 9 2 11 2
22 11 15 7 1 10 9 3 13 2 16 1 11 4 1 9 9 13 9 3 0 9 2
26 1 9 9 2 9 2 7 11 2 0 9 2 13 11 1 9 1 11 13 14 9 9 11 2 11 2
8 2 3 13 9 14 1 11 2
27 11 1 11 13 3 3 7 13 1 15 3 13 2 2 13 11 2 15 9 9 13 1 9 0 9 9 2
9 1 10 9 13 3 1 0 9 2
14 1 11 13 3 3 11 11 7 11 2 9 13 11 2
23 2 11 3 13 2 13 3 2 1 9 7 1 9 3 13 2 2 13 0 9 9 9 2
13 1 9 0 9 11 0 13 1 9 10 9 13 2
27 2 11 1 11 13 9 9 2 1 15 13 9 2 7 16 13 1 11 7 0 9 2 15 13 1 9 2
24 13 7 9 2 16 4 13 9 1 0 9 2 16 4 13 1 0 9 13 2 2 13 11 2
11 16 9 13 9 11 3 1 9 9 11 2
16 3 15 9 13 1 10 9 2 3 15 13 1 9 1 11 2
29 3 4 13 9 0 9 1 9 2 11 1 11 2 7 11 2 11 2 2 1 9 13 9 11 2 11 1 11 2
5 9 1 9 1 11
7 9 11 13 9 9 1 11
27 1 0 9 4 13 1 9 9 0 9 7 0 9 2 15 13 9 0 9 1 9 2 12 7 10 9 2
35 13 9 9 9 7 9 2 1 10 9 15 9 13 13 1 9 1 0 9 1 0 9 1 11 7 10 9 7 1 0 9 1 0 9 2
59 9 9 2 12 1 9 2 12 13 9 2 15 13 13 9 1 9 0 9 2 9 13 9 1 10 9 2 3 9 13 13 10 9 7 13 15 13 1 0 9 2 16 13 9 1 9 10 9 0 1 9 0 9 7 0 9 0 9 2
25 9 13 0 2 15 4 9 13 0 1 0 9 2 9 13 13 9 1 9 7 9 9 0 9 2
32 9 13 1 3 0 0 9 7 13 2 14 15 1 0 9 0 9 2 7 1 9 2 1 15 13 1 9 0 1 0 9 2
59 4 2 14 0 9 1 0 9 3 13 7 4 2 14 13 0 9 2 16 0 7 3 0 9 13 2 16 13 1 0 9 2 13 4 0 9 13 1 9 7 9 0 9 2 16 15 13 2 16 1 0 9 0 9 13 9 10 9 2
38 9 3 13 2 16 15 13 4 13 7 1 0 9 1 10 9 13 1 0 9 2 1 15 4 3 1 9 3 13 9 7 13 0 2 0 2 9 2
26 15 7 13 13 0 9 9 2 16 0 7 3 0 9 7 0 9 0 9 13 13 0 9 1 9 2
10 1 3 0 9 13 0 9 9 13 2
29 3 9 13 0 9 9 1 9 9 2 1 10 9 7 1 9 2 7 15 1 15 3 7 1 9 1 10 9 2
17 13 7 0 2 16 4 9 13 9 2 15 13 0 1 9 9 2
31 10 9 4 13 3 9 7 1 9 2 10 9 1 11 13 13 7 10 9 0 9 9 0 9 0 9 13 7 13 13 2
44 0 9 7 0 9 1 0 9 13 2 3 15 3 13 2 10 0 0 2 0 9 2 1 9 2 3 13 15 1 10 9 13 1 0 7 0 9 0 1 0 9 9 11 2
53 9 0 1 9 13 3 0 9 7 9 2 15 13 9 9 7 10 9 7 13 15 13 1 9 9 0 3 0 9 0 9 2 15 7 1 9 0 9 13 13 0 2 7 7 1 9 0 9 2 15 9 13 2
54 0 9 1 9 0 9 7 0 9 13 1 0 11 1 9 1 12 2 12 2 12 3 0 9 7 9 9 2 12 7 12 2 9 9 2 12 9 12 2 12 2 12 7 9 9 2 12 9 12 2 12 2 12 2
36 9 11 13 9 11 2 16 11 15 4 13 13 0 9 3 1 10 9 9 12 2 12 2 12 2 1 10 9 4 13 1 9 1 9 11 2
12 11 15 13 0 9 1 12 2 12 2 12 2
6 9 7 9 1 0 9
5 11 2 11 2 2
18 1 9 15 3 13 2 16 13 15 3 9 0 2 3 9 1 9 2
16 9 11 15 1 12 9 1 10 2 9 1 9 2 13 9 2
21 9 11 15 13 3 13 1 10 0 9 2 1 15 13 1 9 13 1 0 9 2
17 15 2 15 15 10 9 3 13 2 15 3 13 2 15 13 9 2
6 0 9 1 9 2 2
10 7 1 0 9 13 9 3 0 9 2
14 13 9 2 13 10 9 2 7 3 13 15 3 13 2
17 3 3 1 12 9 2 13 9 11 13 1 9 9 1 10 9 2
6 0 0 9 13 0 9
19 9 11 11 2 15 13 9 9 2 7 14 15 2 2 13 3 0 9 2
22 9 15 3 13 7 0 9 9 9 2 0 9 11 2 11 12 2 12 2 12 2 2
15 15 2 1 0 9 2 13 9 0 0 9 11 2 11 2
8 3 3 15 13 13 0 9 2
32 16 15 9 13 9 15 13 2 15 7 1 10 9 13 11 2 11 2 3 13 2 16 15 13 1 15 0 16 9 9 9 2
10 9 9 13 2 9 0 0 9 2 2
16 9 11 3 13 2 15 1 15 7 10 9 1 10 9 13 2
16 16 4 13 2 13 4 0 9 3 1 0 9 2 9 2 2
18 9 13 0 9 3 1 9 9 1 15 13 14 9 9 1 9 9 2
15 10 9 2 15 9 9 9 13 7 13 13 2 3 13 2
12 13 15 3 0 9 2 14 1 9 11 11 2
41 9 11 13 2 16 2 13 0 13 0 9 2 0 0 9 2 13 2 14 1 9 0 2 7 0 9 2 13 2 14 1 9 0 2 7 13 1 10 9 2 2
27 16 13 1 10 9 2 13 3 13 1 15 2 16 15 13 2 15 7 1 10 9 15 1 15 13 13 2
19 1 9 2 16 13 15 9 15 2 13 13 2 7 3 13 15 1 15 2
38 13 0 15 13 2 15 13 2 16 4 13 16 3 2 15 1 15 13 13 2 7 3 15 3 13 1 9 3 10 0 9 7 9 1 9 10 9 2
28 9 2 16 4 0 13 14 1 0 9 7 13 9 9 2 13 2 14 13 9 9 7 9 2 0 9 13 2
10 9 3 1 9 9 9 9 1 9 2
36 0 9 2 7 15 1 9 2 16 13 1 3 0 9 2 9 7 9 2 3 2 1 9 1 15 3 0 7 0 2 13 1 9 7 9 2
13 7 3 3 13 9 1 9 15 0 7 0 9 2
30 0 9 2 16 13 7 13 15 9 2 13 7 3 13 9 7 9 9 1 2 0 0 2 7 3 1 15 0 9 2
8 9 1 15 13 3 15 0 2
36 7 3 3 13 1 11 2 11 2 16 3 3 13 0 13 2 16 15 15 13 2 16 4 1 9 9 13 10 9 13 1 0 9 0 9 2
3 0 9 9
2 9 2
27 3 0 9 9 0 9 9 11 11 7 9 10 9 13 9 0 9 2 15 0 9 13 1 12 9 9 2
34 9 9 2 11 11 2 13 3 7 9 2 7 9 2 3 9 2 15 1 0 9 13 0 9 7 13 3 10 0 9 9 0 9 2
28 9 4 1 15 13 1 0 9 2 1 0 9 7 1 0 9 7 1 9 0 9 13 3 0 9 0 9 2
46 0 2 0 7 0 9 9 1 0 9 13 3 9 7 9 9 7 13 15 9 1 0 9 2 1 15 4 13 0 7 0 9 0 9 2 16 13 1 0 2 0 7 7 0 9 2
39 1 15 13 9 0 7 15 2 16 15 1 11 13 9 0 9 2 15 13 10 0 9 1 0 9 7 13 15 10 9 2 16 9 13 16 15 3 0 2
22 0 9 9 2 0 9 0 0 9 7 0 1 0 9 7 9 2 10 9 14 13 2
16 3 2 11 11 3 13 1 9 10 0 9 7 1 0 9 2
44 1 0 9 2 3 1 11 13 0 9 2 13 4 10 9 13 1 12 0 2 3 0 9 2 1 9 13 0 9 16 0 9 0 9 2 0 7 3 0 10 9 7 9 2
18 1 10 9 13 9 0 7 0 16 1 9 2 7 7 1 0 9 2
11 9 11 11 7 10 9 1 9 11 11 2
13 0 0 9 1 11 2 12 2 2 12 2 9 2
6 9 2 15 13 10 9
9 0 9 15 9 11 13 1 0 9
13 9 13 9 9 7 15 0 2 15 1 15 13 2
6 9 13 0 9 9 2
7 0 9 11 13 0 9 2
31 10 9 9 2 15 13 9 3 1 9 0 7 9 0 9 2 13 3 3 1 0 9 9 9 0 9 0 1 0 9 2
23 11 13 1 9 12 9 7 2 0 0 9 2 11 11 7 9 3 13 1 0 1 11 2
13 1 0 0 9 1 9 12 7 0 9 11 13 2
25 1 0 9 3 9 13 0 9 2 7 3 15 13 14 3 0 9 1 0 9 7 3 0 9 2
23 9 11 11 2 12 2 2 9 9 2 13 3 11 16 2 9 2 15 13 10 9 2 2
8 10 9 1 9 13 11 11 2
13 15 11 13 7 13 15 2 9 11 2 13 9 2
7 1 11 4 13 0 9 2
18 11 15 13 9 1 0 9 7 15 4 13 2 16 13 15 0 9 2
6 15 4 1 15 13 2
9 1 12 9 9 2 9 7 9 2
25 1 9 0 9 2 1 15 13 1 0 0 9 2 9 1 9 2 9 2 9 2 9 2 2 2
7 15 13 0 9 1 9 2
10 10 9 0 9 7 0 9 13 0 2
7 11 11 7 0 9 13 2
14 9 1 15 3 13 2 16 4 15 13 1 0 9 2
4 15 13 0 2
5 15 13 11 3 2
17 11 3 13 9 11 2 7 3 4 15 13 1 0 9 11 11 2
8 1 15 13 1 10 9 9 2
24 7 9 15 13 0 9 1 0 9 2 16 13 10 9 2 0 9 9 2 3 3 7 3 2
9 14 1 0 9 3 13 9 3 2
6 9 2 1 0 9 2
24 13 4 2 16 16 13 1 11 2 13 4 13 9 1 0 9 2 16 4 15 13 1 11 2
6 13 15 3 1 9 2
20 0 9 9 0 9 2 15 15 13 13 2 13 9 1 0 0 9 7 9 2
11 15 13 3 9 2 9 2 1 0 9 2
19 7 0 0 0 9 13 1 10 0 9 3 12 9 2 15 13 1 9 2
9 13 9 2 16 9 15 13 0 2
40 3 10 9 13 13 3 2 7 3 1 9 3 13 0 9 2 7 16 15 13 9 2 15 13 1 0 9 1 9 1 9 2 3 15 1 15 3 15 13 2
5 9 13 0 9 2
7 7 13 15 1 15 9 2
18 13 1 11 2 3 16 3 9 7 9 9 9 11 11 2 1 9 2
12 13 4 1 11 3 3 1 11 1 9 9 2
8 13 15 1 2 0 9 2 2
4 14 3 14 2
32 15 15 3 13 1 10 9 9 0 7 13 15 3 13 2 7 13 15 2 16 16 15 13 1 0 9 2 13 15 16 9 2
14 7 3 2 0 9 3 1 9 13 7 13 0 9 2
3 13 15 2
22 11 11 2 1 9 2 13 1 0 9 1 0 9 0 2 2 0 9 2 9 9 2
14 0 9 13 1 11 2 3 7 1 9 9 7 11 2
2 0 9
17 1 9 13 3 12 9 1 9 2 3 9 9 13 9 11 11 2
28 1 0 9 13 0 9 1 9 11 10 2 0 9 0 9 2 2 3 15 13 9 11 11 2 3 12 9 2
31 1 9 0 9 11 11 3 13 9 1 9 2 15 13 1 12 9 2 15 13 3 9 1 11 11 2 9 1 12 2 2
21 9 15 3 13 1 0 0 9 2 7 3 13 9 1 9 10 0 7 0 9 2
31 9 0 9 15 1 0 9 13 3 1 9 2 13 1 0 0 9 2 7 3 13 1 9 1 11 2 11 2 0 11 2
20 3 13 1 0 0 9 2 1 9 0 2 0 7 13 9 1 9 11 11 2
29 1 9 12 13 10 0 9 9 0 9 2 3 3 1 9 11 11 13 1 0 7 0 9 3 13 10 0 9 2
8 0 9 13 11 1 0 9 2
15 10 9 11 15 13 16 3 0 9 2 0 7 3 0 2
17 1 9 11 1 9 9 11 13 9 7 0 9 0 3 0 9 2
36 9 15 13 3 0 7 0 9 1 0 9 11 11 7 0 9 1 9 1 9 7 1 11 2 3 15 13 3 0 9 1 9 0 9 0 2
18 13 7 9 0 9 1 0 9 2 1 15 15 11 11 13 3 0 2
29 0 9 2 9 11 1 0 9 1 9 2 13 1 9 2 1 9 7 1 9 2 9 11 11 1 9 12 2 2
36 0 0 0 9 2 15 9 13 3 7 13 2 7 13 9 7 9 1 9 2 13 1 0 0 9 2 9 1 0 0 9 3 10 0 9 2
20 15 4 15 13 1 3 0 9 7 1 0 0 2 0 13 2 2 2 2 2
1 3
16 9 0 9 9 11 11 2 12 2 4 3 3 13 1 11 2
26 9 0 0 0 9 13 9 1 9 12 7 12 2 3 4 9 11 13 9 7 13 9 11 11 12 2
21 9 9 13 0 0 9 1 9 2 0 13 9 2 15 11 13 1 0 0 9 2
9 1 9 1 0 9 13 0 9 12
21 0 9 12 9 1 0 0 9 0 9 13 0 0 2 9 9 12 9 11 11 2
63 16 13 1 9 0 9 2 1 15 13 9 9 9 2 9 1 0 0 9 2 9 2 9 11 7 9 7 0 9 9 11 11 2 2 4 9 12 13 1 9 2 9 2 9 2 9 2 9 2 0 9 2 9 7 0 0 9 1 0 7 0 9 2
11 9 13 0 9 11 3 3 1 0 9 2
18 12 9 15 13 0 9 11 7 0 9 9 7 0 9 9 11 11 2
33 3 13 0 12 9 2 0 9 11 9 11 11 2 9 9 11 11 2 9 11 11 9 1 0 0 9 7 0 0 2 9 9 2
23 1 9 0 9 13 0 9 2 15 1 0 0 9 13 1 12 0 9 1 0 0 9 2
28 9 1 0 9 13 0 9 12 2 9 1 0 9 2 9 0 0 9 4 13 13 0 9 7 9 11 11 2
41 7 3 15 1 9 9 1 0 9 13 12 0 0 9 2 0 9 2 9 2 9 1 9 11 2 3 0 2 9 16 4 13 2 9 7 13 4 15 1 9 2
15 3 12 1 15 4 3 13 1 0 9 7 13 0 9 2
4 3 13 11 2
2 9 2
26 1 9 0 0 9 1 0 9 0 9 11 11 11 2 12 2 13 9 11 11 11 9 11 1 11 2
17 1 10 9 9 2 11 11 15 13 11 11 2 15 9 7 13 2
35 11 2 15 1 10 11 3 13 9 1 0 9 2 13 10 9 0 9 2 9 7 9 2 1 15 0 9 11 12 2 7 3 1 9 2
19 1 0 0 9 13 11 0 7 0 9 0 9 0 9 10 9 1 15 2
19 1 9 1 0 9 13 9 0 9 7 13 7 1 0 9 1 0 9 2
17 13 3 10 0 0 9 2 3 1 0 0 9 1 9 0 9 2
14 0 9 13 1 0 1 10 9 10 3 3 0 9 2
42 0 13 3 0 9 2 11 11 11 2 0 1 9 11 2 9 9 2 16 9 11 11 7 11 11 2 0 16 0 11 2 1 9 0 9 2 7 7 0 0 9 2
39 0 11 16 0 9 15 7 13 1 9 10 0 0 9 2 7 9 15 3 13 2 3 16 0 7 3 0 13 1 10 0 9 2 1 9 1 0 9 2
29 10 0 9 2 7 9 2 13 2 13 7 13 9 2 15 13 3 1 9 2 7 1 0 9 14 7 14 13 2
10 9 0 9 9 13 2 0 9 13 2
31 15 13 13 3 0 2 16 13 13 9 1 9 2 1 9 1 0 9 9 1 9 2 3 0 9 3 13 0 9 2 2
24 9 3 13 0 9 9 1 9 2 3 15 9 12 13 13 10 9 11 2 0 9 9 11 2
23 15 13 10 9 9 0 11 7 10 9 13 16 9 0 9 2 15 15 1 9 13 3 2
23 13 0 11 2 16 4 10 9 7 9 2 0 11 11 2 3 13 3 0 9 3 0 2
32 1 0 9 0 11 15 10 13 2 3 1 9 1 0 9 1 9 12 1 11 11 2 7 9 1 15 9 1 9 13 4 2
17 9 13 14 9 2 16 11 1 11 15 1 10 9 3 3 13 2
8 15 3 14 13 2 2 2 2
13 11 2 11 11 2 9 11 2 11 2 12 2 2
6 9 1 11 2 11 2
23 9 2 11 11 2 9 2 11 11 2 9 2 11 11 2 11 11 2 9 2 11 11 2
14 13 2 11 1 11 2 11 11 2 11 11 7 0 2
5 9 12 2 9 2
6 9 11 13 1 0 11
16 1 9 0 9 7 0 9 15 7 1 0 9 13 0 9 2
20 3 1 0 9 11 11 1 11 13 9 11 7 2 0 9 2 1 0 11 2
13 1 9 12 0 9 13 9 0 7 0 9 11 2
9 1 0 12 9 1 11 13 11 2
26 7 10 9 13 9 11 1 9 1 0 0 9 11 7 0 11 2 15 3 3 13 1 0 9 9 2
12 0 9 0 9 0 0 9 13 9 0 9 2
12 1 9 9 3 13 9 0 1 9 0 9 2
6 0 13 7 0 9 2
31 15 0 0 9 2 9 11 2 11 9 7 11 2 4 13 1 0 0 9 2 16 4 15 10 9 13 13 0 9 9 2
13 15 15 7 3 13 9 13 1 9 9 2 2 2
24 0 9 13 3 3 0 9 9 2 15 15 13 3 14 3 2 16 9 2 13 1 9 2 2
38 1 9 9 3 0 9 11 11 9 9 11 11 9 13 2 2 3 12 9 13 0 0 0 9 11 7 13 2 16 9 0 11 13 12 1 9 9 2
15 13 15 3 1 9 2 15 13 0 2 7 7 0 9 2
18 13 15 3 9 9 0 11 2 7 7 9 2 15 13 3 11 2 2
11 14 12 0 9 11 7 0 11 13 9 2
14 11 9 13 1 0 7 1 0 11 7 9 9 11 2
2 3 2
29 2 9 13 0 9 2 16 13 9 9 1 9 7 11 2 15 13 3 7 13 3 10 9 2 2 13 11 9 2
13 9 9 11 13 1 11 13 0 7 0 0 9 2
11 0 9 13 13 12 12 0 9 1 9 2
28 0 1 15 4 15 13 13 9 2 3 15 3 13 1 0 9 0 11 2 15 13 1 11 1 9 12 2 2
41 9 13 1 0 0 9 7 1 0 9 13 9 7 1 11 2 9 9 9 13 1 9 11 7 3 0 7 15 9 10 9 15 1 10 9 13 3 1 9 2 2
47 11 9 15 3 3 13 13 1 9 9 11 2 7 3 1 0 2 9 2 0 9 1 11 7 1 11 2 3 15 2 1 9 1 11 2 13 1 9 0 0 9 0 9 0 0 9 2
15 2 11 13 3 1 12 1 0 0 9 2 2 13 9 2
18 2 13 0 9 2 0 9 7 9 9 15 1 15 13 3 13 2 2
5 1 0 9 11 11
13 3 4 1 9 1 11 13 9 7 9 11 11 2
25 0 9 3 0 9 0 0 9 2 9 7 9 9 2 12 2 12 2 13 13 1 12 2 9 2
17 13 3 12 9 1 9 12 2 12 2 3 1 0 9 0 9 2
16 1 0 9 0 7 1 0 9 13 11 9 0 9 0 9 2
22 13 15 1 0 9 9 11 2 15 15 13 0 9 3 10 9 10 0 7 0 9 2
8 9 13 0 0 9 7 9 2
23 1 0 13 3 1 9 0 9 2 7 13 7 0 9 9 7 0 9 1 0 0 9 2
9 0 11 13 1 9 9 1 0 9
36 0 9 11 2 9 9 0 11 2 11 2 11 2 0 11 7 0 9 1 9 9 1 9 13 1 9 13 0 9 10 0 0 9 9 9 2
19 1 10 0 9 9 13 3 0 11 7 0 0 9 2 9 7 0 9 2
47 1 0 9 9 0 11 2 15 13 1 9 3 1 0 9 11 2 9 2 1 10 9 2 0 9 11 2 4 3 1 12 9 0 9 10 9 13 2 1 10 9 13 10 9 11 11 2
17 9 7 9 9 0 9 11 1 11 1 11 2 13 15 9 2 2
9 11 3 13 0 9 9 9 11 2
18 10 0 9 15 13 13 1 9 9 1 0 9 7 0 9 1 9 2
16 13 3 9 9 1 0 9 1 9 7 9 9 1 0 9 2
42 0 0 9 0 1 9 7 9 11 2 9 2 15 13 10 0 0 9 1 10 9 2 13 0 9 11 1 12 2 9 3 0 9 1 12 9 14 1 12 2 9 2
5 15 2 3 2 3
21 0 9 9 1 9 13 3 1 12 9 9 11 7 11 0 11 1 9 11 11 2
26 9 9 11 13 9 9 2 9 7 9 11 11 2 0 7 11 0 0 1 0 9 1 12 2 9 2
14 0 9 1 9 13 1 9 9 9 7 9 11 11 2
16 0 9 13 9 9 1 9 11 9 1 0 0 9 1 11 2
14 0 9 11 13 3 3 1 0 9 9 1 0 9 2
7 9 13 0 9 11 11 2
4 9 11 1 11
9 9 0 9 1 11 13 0 9 9
13 1 0 0 9 3 1 11 13 0 9 11 11 2
13 1 10 9 13 13 12 0 2 0 3 0 9 2
24 9 13 3 13 3 3 1 9 2 7 1 9 1 0 9 1 0 9 11 9 1 9 13 2
24 16 13 1 0 9 2 10 9 4 3 0 2 9 2 3 1 15 13 2 13 7 13 9 2
21 16 1 11 2 7 1 11 13 13 3 0 9 1 10 0 9 16 1 10 9 2
28 11 2 11 3 13 1 11 1 9 2 3 9 11 11 13 1 9 7 0 9 0 9 11 11 15 3 13 2
19 7 16 1 0 9 9 11 13 13 2 9 10 9 1 0 9 13 0 2
15 3 9 1 11 13 1 0 9 0 9 1 9 0 9 2
20 3 3 13 2 16 10 0 9 0 9 1 11 13 1 9 10 9 0 9 2
39 7 13 11 3 3 3 13 2 16 9 2 16 10 1 11 2 3 13 10 0 9 2 7 15 7 3 2 16 9 11 13 1 11 9 9 11 1 9 2
31 1 9 9 1 7 1 4 13 13 2 9 7 13 2 16 9 1 3 13 7 16 15 13 9 16 0 2 7 0 9 2
31 3 0 9 3 13 9 9 1 9 1 9 11 1 11 2 15 9 13 13 1 0 9 2 13 2 14 15 13 0 9 2
11 1 12 9 0 9 13 12 9 1 11 2
12 9 1 0 9 15 13 1 12 9 2 9 2
13 11 13 1 9 9 7 0 9 3 13 1 9 2
18 1 9 12 4 11 9 13 1 0 11 12 9 2 9 12 9 3 2
11 11 13 3 13 12 9 2 9 12 3 2
33 1 0 9 1 9 9 7 0 9 13 9 14 11 2 0 9 11 7 0 9 0 0 7 0 9 1 0 9 2 7 7 11 2
18 1 0 0 9 2 15 13 4 13 2 13 9 1 0 9 0 9 2
19 12 9 13 12 9 7 13 1 0 2 0 9 2 3 9 4 3 13 2
8 9 13 13 9 1 0 9 2
31 15 15 1 0 9 3 3 13 1 9 9 12 2 12 2 7 0 9 13 3 1 12 5 7 13 9 12 9 2 9 2
20 11 13 3 1 0 9 1 12 2 9 7 13 4 15 13 1 10 9 3 2
19 9 15 3 13 1 0 9 0 7 0 0 9 2 15 13 4 3 13 2
5 2 13 0 9 2
17 13 9 0 9 7 9 2 2 13 1 15 0 9 9 11 11 2
35 9 4 13 13 0 9 2 7 10 0 0 9 15 13 2 7 1 10 9 13 1 0 9 11 1 9 1 11 2 15 9 13 0 9 2
4 11 13 9 9
2 11 2
24 0 9 2 11 2 13 1 9 0 9 9 1 9 0 9 1 0 9 0 9 1 0 9 2
36 16 13 9 11 11 11 2 9 1 10 9 13 0 9 2 16 3 1 0 9 13 1 9 1 9 11 0 9 2 1 15 13 9 1 9 2
15 11 7 13 16 0 9 9 9 1 0 9 9 11 11 2
23 11 15 3 13 1 9 9 0 9 1 11 2 15 1 15 13 0 9 1 0 9 11 2
30 0 9 13 3 1 9 0 9 9 0 9 2 15 13 13 9 1 0 9 0 9 11 2 1 15 13 9 0 9 2
5 0 9 1 9 11
2 11 2
34 0 0 9 0 9 0 9 11 11 13 1 9 10 0 9 1 11 1 0 9 1 9 0 9 11 2 9 2 1 11 1 9 11 2
21 9 15 1 11 13 1 9 2 9 7 9 9 7 1 9 0 9 1 10 9 2
40 0 9 1 11 11 11 2 15 9 1 11 13 2 1 9 9 13 2 16 0 9 7 9 0 9 15 13 9 0 9 7 16 9 11 4 13 10 9 13 2
4 9 13 0 9
2 11 2
38 0 9 1 0 11 15 3 13 1 0 9 2 16 0 0 9 13 9 11 9 1 15 2 16 1 9 1 9 9 13 2 0 0 9 2 0 9 2
31 1 9 2 15 9 13 9 7 15 4 3 13 1 11 2 13 1 2 3 0 2 0 9 1 0 9 1 9 0 11 2
28 9 3 13 2 16 13 1 9 1 0 9 2 9 7 13 13 13 1 0 7 0 9 9 1 0 0 9 2
5 11 2 13 0 9
8 11 11 13 9 0 9 1 11
30 0 9 11 11 1 10 0 9 1 12 9 9 13 0 0 9 2 16 13 9 11 13 11 16 0 9 1 0 9 2
22 13 2 16 0 0 9 13 0 13 1 2 0 9 11 2 2 16 10 10 9 13 2
13 9 15 11 11 3 13 1 9 1 9 1 11 2
16 13 0 9 0 1 11 1 15 2 16 3 13 10 0 9 2
24 2 14 0 9 2 7 11 13 13 1 9 9 7 9 2 15 13 16 0 9 2 2 13 2
21 9 0 9 0 9 11 11 13 9 1 15 2 16 11 13 13 0 9 0 9 2
11 9 9 11 11 3 13 9 1 9 9 2
15 2 9 13 1 9 1 11 1 15 13 2 2 13 11 2
40 11 11 2 9 0 9 2 13 9 9 2 16 0 7 0 9 15 1 11 13 1 9 2 9 2 2 3 3 13 1 10 9 0 9 2 16 10 9 2 2
22 2 13 15 9 1 15 2 2 13 3 1 9 1 0 9 9 0 9 11 2 11 2
17 1 12 9 13 3 9 0 9 2 15 4 9 13 1 0 9 2
9 10 0 9 15 13 3 0 9 2
15 11 2 11 13 9 9 1 12 1 0 9 1 9 12 2
9 13 9 0 9 9 7 0 9 2
26 0 9 13 1 9 9 2 16 13 1 0 9 2 2 9 9 13 0 9 2 7 9 13 0 2 2
14 13 2 16 9 13 13 9 1 9 7 9 1 9 2
1 3
49 9 0 9 15 3 13 1 9 0 11 1 11 1 0 9 11 2 16 4 15 13 12 2 9 9 9 11 11 2 0 3 1 9 1 0 9 3 3 2 16 3 13 1 9 3 12 9 9 2
38 0 9 0 9 7 9 11 2 0 9 7 9 2 11 2 2 15 15 13 13 3 7 1 9 1 11 2 4 1 9 3 2 9 2 13 1 9 2
24 11 13 12 9 7 0 9 1 9 11 2 16 4 13 12 1 0 9 2 15 3 13 11 2
34 3 1 9 0 9 0 9 11 11 2 11 2 10 9 11 11 2 11 2 3 13 1 0 9 12 2 9 2 7 1 9 15 13 2
16 9 9 13 12 9 0 0 9 1 9 1 11 7 0 11 2
8 13 15 3 0 9 1 11 2
8 9 1 0 9 13 3 0 2
18 1 9 1 0 0 9 11 15 13 9 9 11 11 1 0 0 9 2
10 11 13 13 9 9 0 9 1 9 2
11 13 15 0 9 0 2 11 0 2 11 2
20 9 0 9 11 11 13 1 9 9 15 12 9 2 16 4 0 13 12 9 2
23 11 3 3 13 11 1 9 9 2 16 4 15 13 13 10 9 13 11 13 1 0 9 2
15 0 9 3 13 9 1 9 1 0 9 9 1 0 9 2
28 9 1 9 1 15 9 0 9 1 0 9 2 11 2 2 15 13 9 2 13 1 9 9 0 9 11 11 2
9 0 9 15 13 9 9 0 11 2
4 11 2 11 2
36 0 9 3 13 11 2 16 4 15 1 10 9 13 13 9 0 9 1 9 2 16 4 13 9 0 9 9 0 9 2 9 2 1 0 11 2
10 11 3 3 13 9 0 9 1 11 2
16 9 0 9 15 13 1 0 9 9 1 9 9 9 1 11 2
12 11 1 15 13 2 7 15 3 1 9 9 2
29 1 0 9 1 11 3 0 9 15 9 1 11 9 11 11 13 1 15 2 16 4 9 1 0 9 4 3 13 2
26 0 9 9 2 15 14 11 3 13 2 15 13 13 0 9 9 11 1 11 7 3 0 9 0 9 2
39 11 13 13 13 1 9 0 9 1 11 2 0 11 2 11 2 11 2 11 7 11 2 1 9 0 9 1 11 9 1 9 11 7 11 1 10 0 9 2
12 13 15 1 0 11 0 9 1 11 11 11 2
39 3 1 9 11 13 9 0 9 0 9 0 2 0 11 2 2 9 9 2 1 9 9 1 9 7 9 1 11 7 9 15 12 9 0 11 16 0 9 2
26 1 0 9 11 13 4 3 13 0 9 2 15 1 9 3 13 0 9 9 7 9 0 9 1 9 2
19 0 9 11 13 2 16 9 13 9 2 15 4 13 3 0 9 1 9 2
5 0 9 1 11 11
2 11 2
28 0 9 3 1 11 13 0 9 1 9 7 9 2 11 2 2 16 4 13 9 1 9 0 9 1 0 11 2
23 9 2 15 1 9 1 9 9 13 3 1 0 9 2 4 13 15 0 9 16 0 9 2
32 0 9 3 13 0 9 7 11 2 16 4 13 15 9 0 15 0 9 9 9 2 16 7 9 10 9 7 9 1 0 9 2
4 11 13 0 9
4 11 2 11 2
27 0 9 11 11 2 11 3 13 2 16 10 9 13 9 0 9 1 9 12 9 0 9 1 11 7 11 2
13 13 3 0 9 11 11 2 16 4 9 3 13 2
39 9 13 11 2 11 2 11 7 0 9 16 0 9 0 9 2 15 4 1 9 12 13 0 0 9 1 11 7 11 2 1 15 11 13 3 1 9 9 2
29 1 0 9 13 1 0 9 1 12 9 7 3 9 2 7 15 3 9 2 15 1 9 13 11 7 15 11 13 2
4 9 4 13 9
16 9 10 9 3 13 9 1 9 7 9 0 9 7 10 9 2
7 3 3 3 13 9 10 9
23 13 4 15 3 13 9 0 9 1 9 2 16 13 15 1 9 3 7 16 15 9 13 2
3 14 3 2
8 3 1 9 15 0 9 13 2
22 9 0 9 13 0 2 7 7 13 14 0 13 9 9 2 0 1 0 9 0 9 2
34 3 2 16 7 10 9 9 15 1 9 0 9 9 13 2 1 9 15 7 13 13 2 7 1 0 9 13 9 2 3 10 9 13 2
13 1 9 0 7 0 9 2 13 15 2 9 13 2
13 13 9 1 9 2 1 10 9 1 9 15 13 2
23 16 4 9 9 0 1 9 4 13 0 9 0 9 7 0 9 2 0 9 4 3 13 2
16 16 15 7 1 9 13 0 9 9 2 13 0 9 3 13 2
5 13 15 12 9 2
9 0 1 15 2 9 2 4 13 2
4 9 13 10 2
22 9 4 1 10 9 13 10 9 2 7 3 9 13 15 1 0 9 2 9 3 0 2
12 1 10 9 4 13 13 9 9 1 9 9 2
21 7 13 7 0 2 15 4 9 13 2 7 9 1 0 9 3 13 13 9 9 2
23 13 15 3 9 0 2 0 9 9 7 10 9 0 9 2 1 10 9 9 0 0 9 2
14 16 13 9 1 9 2 13 15 3 3 1 0 9 2
7 13 15 15 0 9 13 2
21 3 13 9 2 16 4 3 9 13 13 9 1 9 9 2 1 9 9 0 9 2
15 3 9 9 13 3 3 13 3 2 3 15 13 13 3 2
20 1 9 9 9 0 9 1 0 7 0 9 13 0 13 9 1 9 0 9 2
12 1 15 0 9 9 15 9 13 3 3 13 2
19 10 9 7 1 9 13 2 7 7 3 3 2 7 3 14 9 9 13 2
15 9 1 0 9 7 10 9 9 1 0 9 3 13 3 2
26 1 9 9 9 9 9 0 9 13 13 0 9 3 2 16 4 9 9 3 1 11 13 3 1 12 2
14 7 15 3 15 2 16 7 3 13 10 9 3 0 2
16 9 9 11 13 0 9 9 15 2 16 14 15 9 13 0 2
20 12 9 7 13 13 1 0 9 3 0 9 2 10 9 13 13 3 3 0 2
10 3 9 13 13 15 9 7 3 9 2
16 3 13 13 2 16 0 0 9 13 13 3 13 1 9 9 2
15 14 0 9 13 9 13 15 1 9 2 15 13 1 9 2
18 3 4 15 3 1 9 13 2 16 13 9 3 0 9 1 0 9 2
26 1 15 9 3 10 9 0 9 13 7 13 3 10 9 2 16 13 1 9 3 0 13 9 9 9 2
17 9 15 15 13 9 1 10 9 1 15 2 3 7 15 4 13 2
24 11 3 13 10 3 0 9 2 16 13 0 13 0 9 0 9 2 16 4 15 0 13 13 2
8 7 15 13 2 15 13 0 2
11 9 15 0 13 1 9 9 3 13 3 2
15 3 4 15 0 0 9 14 13 0 0 9 1 0 9 2
16 9 10 9 3 13 9 1 9 7 9 0 9 7 10 9 2
8 3 3 3 13 9 10 9 2
10 15 3 9 2 15 0 9 10 9 2
16 0 9 13 2 3 16 9 2 15 15 13 13 1 10 9 2
22 10 9 15 13 13 2 16 3 15 13 13 1 9 0 11 15 2 15 13 1 9 2
4 11 13 0 9
15 0 9 0 9 9 9 13 2 16 0 0 9 15 13 2
19 1 0 9 0 9 3 13 9 9 0 9 7 11 2 3 13 9 11 2
32 0 12 9 2 15 13 0 9 1 9 1 0 9 2 11 2 11 7 11 2 13 0 0 9 7 9 10 9 15 3 13 2
17 0 0 9 2 0 11 13 7 1 0 9 0 2 0 9 9 2
13 1 15 0 0 9 13 9 10 9 1 3 0 2
6 3 13 1 15 9 2
19 7 16 10 0 9 15 9 7 0 9 1 9 11 13 2 13 3 0 2
12 3 1 15 9 0 9 13 1 15 0 11 2
18 0 9 13 14 0 9 9 2 15 13 9 1 0 9 3 0 9 2
10 0 9 0 9 1 0 9 13 11 2
17 7 16 9 10 9 13 3 1 0 0 9 2 0 9 13 0 2
23 11 13 1 0 9 12 10 9 2 1 9 4 15 13 12 7 1 9 3 12 9 9 2
33 0 9 0 9 1 0 9 2 0 0 9 1 0 9 2 9 0 7 0 2 9 2 13 9 14 11 2 7 7 0 0 9 2
17 1 9 4 1 2 0 9 2 13 1 12 9 9 3 16 9 2
36 15 13 13 2 16 11 13 10 9 3 0 9 2 15 15 1 9 9 13 1 0 0 9 2 7 13 9 13 15 10 9 7 13 1 11 2
26 1 10 9 13 9 11 1 0 9 0 2 7 3 14 13 13 7 10 9 2 15 4 3 9 13 2
11 10 9 13 3 1 0 9 9 0 9 2
28 1 1 15 2 16 9 15 13 12 9 1 9 0 9 2 13 0 2 16 7 0 9 9 10 9 13 0 2
11 10 9 11 3 1 10 9 13 7 3 2
12 3 15 13 13 1 9 1 0 9 10 9 2
27 0 0 9 13 1 9 7 0 0 9 9 11 2 15 13 1 0 2 0 2 9 1 10 9 3 9 2
15 1 9 10 9 1 9 0 9 13 1 0 9 1 11 2
17 7 15 2 15 13 1 9 1 10 9 2 13 3 1 15 9 2
20 0 9 13 3 2 16 13 0 9 1 0 9 16 1 0 9 1 10 9 2
11 0 9 9 13 1 0 9 14 0 9 2
13 1 0 9 1 0 9 9 15 9 10 9 13 2
30 0 9 11 7 3 0 9 0 9 2 3 15 3 0 1 0 9 2 13 2 16 15 0 9 13 0 9 0 9 2
19 13 15 2 16 1 3 0 9 15 13 0 9 2 1 15 13 0 13 2
8 13 15 1 9 9 0 9 2
11 9 3 3 13 10 9 1 3 0 9 2
26 0 9 9 0 0 9 7 3 0 9 11 13 13 2 16 0 9 4 1 15 13 3 10 12 9 2
35 0 9 0 9 7 3 7 9 13 2 13 15 2 9 9 1 9 2 3 15 13 10 9 11 2 7 9 1 9 1 0 9 7 9 2
7 9 15 1 0 2 9 13
29 0 9 1 0 9 9 3 0 9 1 0 9 1 9 13 1 9 9 13 9 0 2 11 10 9 9 0 9 2
17 2 0 9 13 9 2 3 0 9 9 2 15 4 3 13 2 2
29 9 13 3 0 2 16 0 0 9 2 15 13 13 0 9 0 9 2 13 13 1 9 9 1 0 9 0 9 2
19 0 9 13 9 9 0 2 13 9 9 2 9 9 1 0 9 1 0 2
28 13 3 9 2 16 4 15 13 10 0 9 9 13 13 9 0 9 0 9 1 9 10 2 3 1 0 9 2
21 15 4 15 13 2 16 4 15 10 0 9 1 9 7 1 0 2 11 3 13 2
27 13 1 9 9 11 7 13 2 16 1 9 4 13 1 9 12 1 9 7 1 0 2 11 1 12 9 2
20 1 9 4 9 11 3 13 2 16 13 2 16 3 3 1 10 9 13 3 2
18 13 3 0 9 9 2 9 15 13 7 9 11 4 3 7 3 13 2
19 1 0 2 11 3 10 9 9 13 9 9 3 2 16 4 13 9 13 2
17 15 4 3 1 0 2 11 13 2 16 1 9 13 9 3 0 2
15 1 0 9 15 9 9 11 1 12 9 13 1 0 9 2
21 13 3 0 2 16 0 9 0 9 3 3 0 9 4 13 13 1 0 9 9 2
24 3 0 9 1 9 7 1 0 2 11 13 0 9 0 9 9 7 13 0 9 1 0 9 2
2 0 9
20 1 12 2 9 12 13 3 1 0 12 9 1 0 9 3 12 2 0 11 2
21 13 3 1 0 9 1 9 9 2 15 13 1 9 12 9 9 1 0 9 9 2
16 9 3 13 1 9 10 0 9 7 1 9 13 9 0 9 2
7 0 9 3 13 1 9 2
19 0 9 13 1 12 9 0 3 1 9 11 7 9 0 9 1 9 11 2
14 9 11 4 1 10 12 9 9 13 1 0 1 9 2
25 9 10 9 13 3 3 1 9 9 9 2 3 1 9 0 0 9 0 9 3 13 14 12 9 2
18 0 9 13 12 1 9 2 15 9 1 10 9 13 14 3 1 9 2
27 9 1 9 0 9 2 15 9 9 13 2 1 9 7 1 9 9 2 1 0 9 2 13 1 12 9 2
20 9 10 9 13 3 0 2 1 3 0 9 14 1 0 9 7 3 7 9 2
6 0 9 9 3 13 2
17 1 10 9 13 3 12 9 7 3 4 13 0 7 3 0 9 2
19 9 2 15 15 13 9 9 1 0 9 1 12 9 2 4 13 3 13 2
15 1 15 3 13 2 16 15 9 13 3 13 3 0 9 2
12 3 1 9 9 13 2 16 9 9 13 0 2
26 9 3 13 2 16 13 9 13 0 9 9 1 9 10 10 9 2 7 9 9 13 3 1 12 9 2
9 14 2 15 9 13 1 9 9 2
13 9 2 15 13 9 9 2 4 3 13 3 9 2
26 9 9 9 13 13 9 1 0 9 1 0 9 2 15 4 9 0 9 7 9 0 0 9 3 13 2
38 15 2 16 9 13 3 0 9 2 13 15 7 0 9 0 9 7 9 2 0 9 2 0 13 3 3 2 13 1 9 0 9 7 15 2 10 2 2
11 3 13 2 16 13 10 9 1 9 9 2
11 1 10 9 15 3 13 9 1 9 1 9
5 14 2 0 9 2
2 11 2
19 0 9 13 1 9 3 1 9 9 1 0 7 0 9 1 12 9 9 2
24 1 0 9 2 15 13 9 0 9 1 0 9 9 1 0 9 2 13 0 12 9 9 9 2
13 0 9 0 9 10 9 13 2 3 16 13 9 2
15 13 15 1 0 1 9 9 2 15 1 0 9 13 9 2
7 2 10 9 15 13 9 2
36 1 0 9 9 15 3 13 9 1 0 0 3 1 12 9 1 9 2 16 4 15 9 15 13 2 2 13 9 2 11 1 0 9 0 9 2
11 3 1 15 13 9 1 9 1 0 9 2
15 16 13 1 9 0 9 2 13 9 1 0 7 0 9 2
10 13 15 2 0 9 13 7 9 13 2
12 3 1 9 13 9 0 2 16 15 9 13 2
29 1 0 9 9 1 9 9 0 1 0 0 9 13 9 0 9 9 11 2 11 3 9 9 1 3 0 0 9 2
10 15 1 9 9 13 14 12 12 9 2
6 0 9 7 13 13 2
15 2 7 16 4 13 3 12 12 2 3 4 15 3 13 2
12 13 13 1 9 2 2 13 11 12 1 9 2
23 0 9 3 1 0 9 9 15 13 7 0 9 2 7 9 7 9 0 9 1 10 9 2
20 16 7 9 3 13 9 0 0 9 2 13 1 11 2 11 13 1 9 9 2
8 15 7 13 7 0 0 9 2
10 9 13 3 9 15 1 9 9 13 2
8 1 0 9 9 13 13 3 2
15 13 0 13 15 0 9 7 13 9 0 9 3 1 9 2
11 15 13 7 13 14 9 2 15 9 13 2
17 9 2 16 9 9 4 13 3 2 10 2 9 2 13 7 0 2
6 0 9 0 9 3 13
2 11 2
18 9 15 3 10 9 13 13 0 9 2 15 3 13 9 9 11 11 2
28 16 1 9 9 13 0 9 7 9 11 11 2 15 13 11 1 9 13 2 13 9 9 9 0 9 3 13 2
19 3 4 3 3 13 1 0 11 2 9 11 3 13 10 0 9 11 11 2
16 15 3 9 10 9 13 9 0 9 1 11 1 9 1 9 2
9 9 9 7 3 1 10 9 13 2
2 9 9
3 0 11 2
27 1 9 1 9 13 12 3 0 9 0 9 1 9 14 12 9 1 9 0 9 1 0 9 1 0 11 2
12 9 9 7 0 9 13 2 16 4 15 13 2
15 16 12 13 9 1 0 9 2 12 9 13 1 0 9 2
4 13 12 9 2
5 9 11 11 13 0
5 11 2 11 2 2
20 0 9 1 11 3 13 1 9 9 1 11 11 2 15 13 13 12 0 9 2
5 9 13 0 9 2
20 11 4 13 1 12 9 9 9 2 7 0 9 9 13 7 13 9 1 9 2
10 9 3 13 12 1 0 9 11 11 2
14 15 13 2 1 12 9 2 9 9 13 1 9 9 2
17 3 15 14 13 1 0 9 7 13 1 15 9 2 15 0 13 2
15 9 3 1 9 12 7 12 9 13 2 16 11 13 9 2
22 3 1 9 7 13 2 16 15 2 13 2 11 13 16 9 2 15 13 1 9 9 2
8 11 7 11 13 9 9 9 9
5 14 2 0 9 2
2 11 2
40 9 0 9 1 9 9 11 11 2 11 2 7 11 11 2 11 2 11 2 3 13 9 1 9 2 15 9 13 1 9 11 2 16 9 13 9 1 9 9 2
30 11 13 2 16 0 9 13 1 0 9 1 10 0 9 2 3 1 0 9 9 1 9 7 1 9 0 2 0 9 2
27 11 2 15 0 9 3 13 2 13 13 2 16 4 9 13 9 2 1 15 4 13 9 1 0 9 9 2
20 13 3 13 2 16 9 13 2 16 4 13 2 7 13 14 0 7 9 0 2
27 13 15 2 16 3 1 12 9 1 0 2 0 9 13 13 2 16 9 1 15 13 1 0 7 0 9 2
14 9 7 1 11 10 9 13 1 9 7 13 0 9 2
9 11 7 11 13 1 0 9 9 2
17 11 9 9 13 1 0 7 1 10 9 2 16 1 15 13 9 2
29 2 1 15 2 16 15 13 9 9 2 9 1 9 13 7 9 10 9 3 15 13 0 1 9 2 2 13 11 2
22 11 13 2 16 0 9 4 13 13 7 0 9 9 11 11 2 15 1 15 15 13 2
14 0 9 13 9 2 15 13 0 3 13 1 15 9 2
15 13 3 13 0 9 2 16 4 1 9 13 10 0 9 2
5 0 9 15 15 13
24 9 0 9 9 0 9 2 9 1 9 7 0 2 0 9 13 9 0 9 1 9 11 11 2
6 11 13 1 9 11 11
2 11 2
24 13 0 2 16 4 4 15 12 9 1 9 13 1 9 1 0 9 1 9 9 0 0 9 2
13 3 15 13 9 11 11 11 1 9 9 11 11 2
20 1 10 9 13 1 0 9 1 11 2 2 3 0 9 16 9 1 9 2 2
19 1 11 13 9 2 16 1 0 9 13 9 7 16 4 9 3 3 13 2
26 11 13 9 10 9 1 9 9 1 9 0 9 9 2 7 13 14 1 9 0 2 0 7 3 0 2
25 11 13 2 16 15 13 13 2 16 4 13 0 13 2 15 13 9 1 9 7 15 1 9 9 2
18 2 13 15 14 9 1 9 2 15 15 15 13 10 9 2 2 13 2
1 3
32 9 0 9 11 11 11 1 0 0 9 13 9 9 0 0 9 11 11 2 16 15 1 15 0 9 13 1 0 0 0 9 2
20 2 10 9 1 11 11 13 3 1 9 0 9 16 9 2 2 13 11 11 2
10 0 9 14 4 13 1 0 9 0 9
2 11 2
24 1 0 9 0 9 2 15 13 11 2 13 0 0 9 0 9 1 9 1 9 14 12 9 2
23 11 15 13 2 3 1 10 9 13 0 9 2 15 9 1 0 9 1 9 3 9 13 2
10 9 11 11 11 3 13 10 0 9 2
6 16 0 9 13 11 2
17 11 15 13 2 16 4 9 11 1 9 13 9 0 9 1 11 2
19 0 9 1 11 13 2 16 13 12 9 2 7 13 7 13 1 0 9 2
26 9 0 9 0 9 11 11 13 13 2 16 10 9 13 13 0 9 9 2 16 15 13 1 0 9 2
10 2 10 9 3 13 13 2 2 13 2
16 1 0 0 0 9 0 9 15 13 1 11 13 14 9 9 2
16 9 9 0 11 2 11 13 9 1 9 1 0 9 1 0 2
20 0 1 10 9 13 1 9 7 9 7 13 0 13 1 0 2 9 7 13 2
12 11 3 0 9 13 1 9 1 0 0 9 2
10 1 0 9 13 9 11 11 0 11 2
12 11 3 13 1 0 9 1 0 9 7 11 2
14 1 9 11 2 11 15 13 9 1 0 9 1 11 2
8 11 11 13 1 9 9 11 12
2 11 2
26 11 2 11 4 13 2 16 4 0 0 9 0 9 4 13 2 7 16 4 13 1 9 10 0 9 2
8 13 15 3 9 9 11 11 2
17 0 9 2 15 11 12 13 2 4 1 15 13 1 0 9 13 2
47 1 3 0 9 1 0 9 9 11 12 4 9 0 9 13 1 15 2 16 4 2 0 9 13 10 9 16 10 0 0 1 9 7 1 0 9 2 15 13 1 0 9 2 2 13 11 2
5 9 9 1 9 13
2 11 2
20 9 9 1 0 9 1 0 0 9 1 9 1 9 0 9 2 11 2 13 2
7 13 15 1 10 0 9 2
17 9 13 9 3 12 9 0 2 16 3 1 9 15 13 12 9 2
13 9 13 12 9 9 2 16 3 15 13 12 9 2
12 1 9 0 15 13 9 1 11 7 1 11 2
21 0 9 15 13 1 0 7 0 9 1 12 9 2 3 0 9 13 12 9 0 2
9 9 13 0 9 1 0 9 0 2
26 0 9 1 9 1 9 0 9 13 3 0 9 2 16 0 2 1 9 12 7 12 9 13 3 0 2
8 9 9 11 11 1 0 0 9
5 9 11 1 9 9
11 1 0 9 15 3 9 13 1 12 9 9
2 11 2
19 3 12 9 15 9 0 0 9 11 3 13 9 2 1 9 13 0 9 2
17 13 1 15 3 9 9 11 11 2 1 10 9 3 10 9 13 2
11 9 9 10 9 9 13 9 11 1 0 2
12 1 9 1 15 3 13 2 13 14 7 0 2
32 1 9 1 9 9 0 11 2 15 1 12 9 13 9 2 13 2 16 11 1 9 12 13 7 13 9 1 9 12 9 9 2
27 1 9 9 2 15 13 3 1 0 9 2 7 1 9 9 13 1 0 9 9 1 0 9 12 9 9 2
28 9 9 11 4 1 9 11 13 9 3 1 9 12 2 7 2 3 1 9 0 9 1 9 9 0 11 9 2
11 9 1 0 9 4 3 13 1 0 9 2
13 1 9 9 9 13 12 0 9 7 12 0 9 2
9 9 1 15 13 7 3 4 13 2
18 0 15 13 13 3 12 0 9 7 9 9 1 0 9 12 9 9 2
19 16 11 13 9 9 11 11 2 9 15 12 0 9 13 13 1 0 9 2
15 9 1 9 9 4 13 4 13 1 9 0 9 0 9 2
8 0 9 14 13 1 0 9 2
15 1 9 13 7 1 9 2 16 4 11 9 0 9 13 2
9 1 9 15 13 7 1 9 9 2
37 1 9 0 0 9 11 4 1 9 11 3 9 13 9 9 0 0 9 9 1 9 12 9 9 7 0 9 0 0 9 11 1 9 12 9 9 2
9 1 10 9 15 3 13 0 9 2
23 9 9 11 11 13 2 16 10 9 13 15 0 1 0 0 9 0 11 7 10 0 9 2
15 9 13 2 16 0 9 13 9 2 7 7 9 9 1 15
5 14 2 0 9 2
2 11 2
12 1 0 9 4 15 13 13 9 9 16 9 2
19 1 0 9 0 0 9 7 0 0 9 15 13 11 11 1 9 0 9 2
29 9 7 9 3 13 1 0 1 15 2 16 0 9 1 9 4 13 10 0 9 7 13 15 7 1 9 9 9 2
6 0 13 2 16 14 2
27 9 13 1 9 2 16 15 9 4 13 1 12 7 12 9 3 16 1 0 9 7 4 13 3 7 9 2
8 0 9 15 13 1 0 9 2
15 9 4 13 13 7 0 7 9 0 2 7 16 14 0 2
10 9 7 3 13 1 9 0 9 9 2
18 1 9 11 11 13 9 0 9 1 9 3 1 11 3 1 9 12 2
29 7 7 1 0 9 3 0 9 0 1 9 13 2 16 2 15 13 13 9 2 7 0 2 16 13 15 10 2 2
10 0 9 3 13 3 0 9 1 9 2
22 1 9 13 1 10 9 7 3 0 2 15 15 9 13 2 7 3 15 15 4 13 2
14 9 9 15 13 9 2 16 13 4 0 9 15 13 2
26 9 13 2 16 3 4 13 0 9 2 1 11 3 13 12 9 2 7 0 9 4 13 9 3 13 2
22 1 15 9 9 0 9 1 11 13 2 16 1 9 3 13 0 0 9 7 10 9 2
10 12 12 0 13 2 16 13 0 9 2
26 11 9 1 0 9 9 7 0 9 13 1 9 2 16 3 0 1 0 9 13 9 0 9 7 9 2
22 10 9 1 15 13 1 0 9 9 1 0 9 7 0 9 13 15 1 9 0 9 2
8 9 9 9 13 1 9 9 11
5 14 2 0 9 2
2 11 2
22 9 1 9 1 2 0 9 2 9 0 9 13 3 1 10 9 10 9 0 9 9 2
24 1 15 15 9 13 1 9 11 11 2 9 2 15 16 2 16 4 9 13 2 13 15 2 2
17 9 15 13 2 3 3 15 0 9 1 9 0 9 7 11 2 2
30 13 1 9 9 2 15 1 15 13 9 9 2 16 13 11 11 1 9 9 0 9 9 9 7 13 1 9 10 9 2
30 0 9 11 9 3 13 2 16 2 9 13 1 0 13 10 9 1 9 0 9 3 7 2 16 9 9 9 13 0 2
8 1 9 9 15 3 13 2 2
26 1 0 9 9 13 2 2 4 13 2 16 16 0 9 13 13 0 9 1 9 0 9 9 9 2 2
18 9 9 9 1 10 9 1 9 9 0 9 3 13 9 9 11 11 2
13 10 9 13 1 15 12 1 0 9 9 1 9 2
7 9 0 2 11 13 0 9
2 11 2
28 9 0 11 13 12 12 9 11 1 0 9 7 9 1 15 15 13 2 16 4 13 13 1 9 0 0 9 2
17 1 9 1 0 9 1 9 7 9 9 15 1 11 13 9 11 2
9 1 9 13 12 9 0 12 9 2
24 9 0 2 11 13 1 9 0 9 3 0 9 2 9 1 0 9 7 15 2 15 13 0 2
15 0 11 7 9 15 13 2 16 4 9 13 13 9 9 2
38 3 0 0 9 11 13 1 15 2 16 4 9 9 13 13 0 0 9 2 0 4 9 0 2 11 13 1 9 9 7 0 0 4 10 9 13 9 2
17 1 9 9 9 13 3 9 2 9 2 9 7 9 1 0 9 2
16 16 4 9 13 9 2 13 3 9 2 9 0 9 7 0 2
5 9 11 3 1 9
2 11 2
19 9 9 11 11 3 13 9 1 9 9 1 0 9 0 0 9 11 11 2
10 13 1 15 0 9 9 9 11 11 2
38 9 11 11 1 15 13 0 9 1 11 2 15 1 9 4 13 2 16 4 13 2 16 9 0 9 4 13 9 1 9 0 7 16 4 10 9 13 2
17 9 15 3 13 2 16 13 0 1 10 9 13 0 9 2 13 2
13 9 11 11 4 13 1 9 0 9 0 0 9 2
30 13 15 15 13 15 2 16 1 9 12 7 12 13 7 13 0 9 9 9 1 9 0 9 9 0 11 1 9 9 2
18 0 9 1 11 15 1 9 9 13 1 9 12 1 0 9 9 9 2
22 11 11 15 13 7 1 9 9 0 9 0 0 9 1 11 0 9 3 1 9 13 2
13 1 0 9 9 1 9 13 9 9 1 0 9 2
6 11 13 13 9 1 9
2 11 2
40 9 9 0 1 9 9 9 2 11 11 7 11 11 7 10 9 11 11 2 4 1 9 13 1 0 9 9 0 9 2 16 10 0 9 13 0 9 1 9 2
11 9 15 13 9 0 0 9 9 11 11 2
20 1 15 13 9 9 2 3 11 7 10 9 13 2 16 4 9 1 9 13 2
14 16 7 9 13 10 9 2 13 15 14 12 9 9 2
26 11 15 13 2 16 4 15 9 13 13 3 9 9 1 9 2 15 7 1 15 13 2 3 4 13 2
10 11 13 1 10 9 3 0 12 9 2
21 9 15 13 2 16 1 9 13 7 15 2 15 13 0 0 9 13 3 1 9 2
19 9 15 13 9 13 3 2 16 3 13 9 9 9 2 0 9 0 9 2
13 3 13 3 2 16 9 9 10 9 13 1 9 2
18 1 11 9 1 11 7 11 13 12 0 9 9 0 9 9 9 9 2
24 9 15 1 9 13 1 9 1 9 9 11 11 2 15 15 1 9 9 13 1 0 9 9 2
18 1 9 9 4 13 1 9 9 1 11 1 11 1 0 9 1 11 2
11 1 10 9 13 10 9 9 1 0 9 2
7 9 9 11 3 13 9 2
11 1 9 11 13 1 9 13 0 9 9 2
6 0 9 1 11 14 13
2 11 2
15 9 9 2 15 13 1 11 2 13 1 0 9 13 9 2
9 13 15 0 9 0 9 11 11 2
10 2 10 9 13 3 13 2 2 13 2
24 11 11 1 9 0 9 3 11 13 2 16 1 10 9 13 4 0 0 1 9 3 13 3 2
31 1 9 15 13 1 0 9 3 1 9 12 2 7 3 0 9 13 3 0 7 0 15 13 9 3 1 12 9 1 9 2
19 9 15 1 9 9 0 11 13 3 1 0 9 0 9 1 11 7 11 2
13 0 1 15 15 13 7 13 10 9 13 0 9 2
9 1 13 13 7 9 9 1 9 2
19 13 14 0 2 16 4 11 13 0 9 1 11 7 16 4 15 13 13 2
13 3 15 2 15 15 3 13 2 4 13 0 9 2
5 9 9 11 1 9
2 11 2
23 0 0 9 9 11 4 12 2 9 13 1 0 0 9 1 0 9 9 9 9 7 11 2
21 0 9 4 13 1 9 12 2 9 9 0 9 9 11 2 15 15 13 1 11 2
24 9 0 9 11 11 11 2 11 4 13 12 0 9 0 0 9 2 0 9 2 9 7 9 2
21 9 4 3 13 12 9 2 15 13 13 1 9 2 0 9 7 1 0 0 9 2
15 9 4 13 1 9 7 0 9 1 12 9 7 0 9 2
7 0 9 4 13 13 12 9
2 11 2
29 3 12 9 4 13 13 1 9 0 9 1 11 7 11 1 0 0 9 2 7 1 10 9 15 13 10 9 13 2
20 13 15 3 9 0 9 0 9 11 11 1 9 0 7 0 9 9 1 11 2
13 9 4 13 1 9 9 13 9 7 9 12 9 2
21 9 9 0 0 9 15 1 9 12 9 13 1 11 2 11 7 11 2 13 11 2
28 9 13 1 11 1 9 0 7 0 9 9 3 16 12 0 9 2 15 13 3 13 1 0 0 2 0 9 2
20 13 13 0 9 2 1 0 9 13 9 2 9 2 2 1 0 2 9 2 2
13 1 12 0 9 1 11 7 1 11 13 9 13 2
12 0 0 9 4 13 12 2 12 2 1 11 2
4 0 9 9 13
7 0 9 13 9 0 12 9
2 11 2
20 3 13 9 13 1 0 9 1 10 0 9 2 15 15 13 2 13 15 9 2
12 3 13 0 9 3 7 3 13 0 9 9 2
23 2 0 9 15 3 1 9 12 13 14 0 0 9 2 2 13 11 11 11 1 9 9 2
21 1 0 0 9 2 1 15 13 0 0 9 13 2 4 13 1 15 13 0 9 2
18 9 9 1 9 13 2 16 4 0 9 0 1 9 10 9 13 9 2
17 0 9 9 9 11 11 15 7 13 2 16 4 15 13 3 0 2
17 2 16 4 13 9 1 9 2 13 0 2 16 4 15 3 13 2
14 1 9 15 4 15 13 1 0 9 9 13 0 9 2
24 13 7 0 3 13 0 9 1 0 9 0 9 2 16 3 1 15 13 0 9 0 9 2 2
34 0 9 13 13 9 0 9 2 7 3 4 15 14 13 13 0 9 3 1 9 1 0 9 7 15 2 15 13 1 9 1 0 9 2
7 13 3 13 0 9 9 2
13 0 9 13 0 9 7 9 2 1 9 3 9 2
11 10 9 4 3 16 0 0 9 13 9 2
10 9 13 3 0 9 1 9 1 9 2
10 2 15 13 3 15 2 15 15 13 2
26 13 15 13 9 2 15 13 9 1 0 9 7 3 9 2 15 13 9 1 15 2 2 13 11 11 2
25 1 9 0 9 0 0 9 11 11 13 0 9 9 12 9 2 15 13 3 1 11 12 9 2 2
9 3 13 9 13 1 0 0 9 2
27 10 9 7 10 13 7 7 9 13 14 14 12 9 0 9 2 15 3 13 3 9 9 7 10 0 9 2
5 0 9 13 1 9
2 11 2
30 1 11 2 1 9 0 9 2 1 10 9 13 12 12 9 9 7 0 9 1 12 9 9 2 13 9 1 9 0 2
22 13 3 1 11 2 3 13 3 3 2 0 9 1 9 13 7 1 0 7 0 9 2
17 3 1 9 9 7 1 11 9 13 7 13 15 7 1 0 9 2
10 1 9 13 0 9 1 9 7 11 2
5 1 11 13 0 9
2 11 2
46 7 3 15 13 9 0 9 7 9 0 0 9 1 9 9 11 11 13 9 1 9 11 2 11 1 9 0 2 0 9 2 9 2 9 7 9 2 10 9 4 13 1 9 1 9 2
19 9 13 1 10 9 1 9 9 7 9 2 15 13 11 11 7 11 11 2
21 9 7 9 15 13 3 1 15 2 16 9 9 4 13 13 0 9 9 11 11 2
29 16 9 4 13 13 1 9 9 2 13 15 9 2 16 15 13 14 1 0 9 7 0 9 2 13 3 11 11 2
3 1 9 11
2 11 2
14 1 9 11 1 9 1 11 13 0 9 11 11 11 2
26 9 11 1 9 1 11 4 1 11 14 13 9 0 9 1 11 7 13 4 0 9 9 1 0 9 2
3 3 9 2
15 0 9 13 10 0 0 9 1 9 2 13 3 0 9 2
52 13 1 15 2 16 9 9 13 12 9 9 0 9 1 0 7 0 9 2 10 9 2 15 15 3 13 0 0 9 2 9 2 7 15 0 0 0 9 13 3 16 0 9 2 14 1 9 9 0 9 2 2
21 3 13 13 1 0 9 2 15 4 13 15 9 0 1 9 11 7 9 15 13 2
27 0 16 2 9 2 15 13 9 2 16 15 3 13 1 9 2 10 12 9 1 0 9 0 9 3 13 2
15 13 15 3 2 16 9 7 0 0 9 13 1 0 9 2
16 0 9 15 3 13 0 2 16 4 15 13 1 0 9 13 2
34 13 15 2 16 0 9 2 15 13 9 10 9 13 2 13 9 2 15 13 13 2 16 7 1 11 15 13 3 0 9 1 9 9 2
26 3 0 2 0 2 9 15 3 3 13 2 0 7 13 2 16 4 9 9 13 3 1 9 9 9 2
24 1 10 9 9 15 3 13 9 3 0 9 2 0 9 13 3 0 7 3 1 0 9 13 2
15 9 0 9 13 3 0 7 0 2 9 1 0 9 2 2
25 3 3 15 13 13 2 16 1 9 2 3 4 0 9 9 13 2 13 3 0 7 0 0 9 2
30 0 9 1 9 13 1 10 9 9 2 16 0 9 12 9 13 7 0 1 0 9 2 15 15 13 1 0 0 9 2
10 2 3 3 7 3 0 0 9 2 2
22 9 0 9 13 0 0 9 0 9 10 9 7 0 9 9 1 7 1 15 3 13 2
30 1 9 0 9 1 15 2 16 0 9 13 0 9 0 9 2 13 0 0 9 13 15 0 16 9 3 13 1 9 2
24 3 3 15 7 7 13 1 9 2 15 2 15 13 9 9 9 2 4 15 3 3 13 13 2
18 0 9 3 13 13 0 9 2 15 0 0 9 1 10 9 9 13 2
20 7 16 15 0 9 13 3 0 9 11 11 2 0 7 0 9 13 3 13 2
5 11 1 9 1 9
2 11 2
10 9 13 15 1 9 9 1 0 9 2
17 13 15 1 9 11 11 1 0 9 9 0 9 7 0 0 9 2
18 9 15 3 13 1 0 9 15 0 9 2 15 13 9 0 0 9 2
17 11 11 13 2 16 0 9 13 1 0 9 13 0 9 0 9 2
13 13 7 9 2 16 4 11 13 9 9 0 9 2
13 1 9 9 11 2 11 9 13 7 9 0 9 2
17 16 9 13 2 9 4 0 9 13 0 9 0 9 1 0 9 2
5 3 9 2 9 12
4 9 11 1 9
2 11 2
20 3 9 7 9 1 11 15 13 1 0 9 1 12 9 9 0 9 11 11 2
15 9 12 13 3 3 7 1 0 9 9 0 13 0 9 2
9 0 9 3 13 9 9 1 11 2
19 13 2 16 13 0 13 9 0 0 9 2 15 13 9 0 9 11 11 2
19 2 3 15 13 0 9 1 9 11 2 2 13 0 9 1 11 11 11 2
19 13 2 16 9 13 3 13 1 9 0 9 7 16 13 0 15 3 13 2
14 2 13 3 13 3 0 9 1 0 9 2 2 13 2
8 3 3 3 13 9 9 11 2
13 1 15 4 10 9 13 9 3 1 12 2 9 2
4 3 1 9 12
6 12 9 1 9 9 12
2 11 2
24 0 0 2 9 9 12 9 11 11 13 12 1 12 0 9 1 0 0 9 2 0 9 11 2
16 9 1 0 9 3 13 0 9 11 9 11 1 0 9 9 2
38 9 12 15 7 13 1 9 9 2 0 1 9 0 9 2 9 9 2 9 1 0 0 9 2 9 2 9 11 7 9 7 0 9 9 11 11 2 2
13 0 12 0 9 13 1 0 9 3 1 12 9 2
10 9 9 0 9 15 4 13 9 9 2
4 3 1 9 12
17 11 11 2 11 11 7 9 0 9 0 9 11 11 1 0 9 9
4 9 1 9 13
8 11 13 9 0 9 1 0 2
2 11 2
14 0 9 1 9 9 3 13 9 0 11 1 9 9 2
8 9 3 13 10 3 0 9 2
20 3 7 13 13 0 9 2 3 2 15 2 15 13 1 11 11 7 11 11 2
63 0 9 9 9 12 2 11 11 2 13 2 11 11 2 11 2 11 11 2 11 2 11 11 2 11 2 11 11 2 11 2 1 12 2 11 11 2 11 7 11 11 2 11 2 11 2 13 2 16 13 10 9 0 1 15 2 16 9 13 9 0 9 2
24 9 15 3 13 2 16 13 15 2 15 4 13 0 9 9 1 9 1 9 13 0 9 9 2
50 9 13 3 1 9 9 9 9 11 11 2 16 15 1 9 0 9 7 1 9 0 1 10 9 13 1 9 1 9 0 7 0 9 11 11 7 9 9 11 11 11 1 9 10 0 9 1 0 9 2
51 1 0 9 9 11 2 3 0 9 9 1 0 9 2 15 9 9 13 3 1 9 7 15 3 2 16 1 9 1 9 12 13 1 9 9 1 9 9 1 0 9 0 9 2 15 13 13 1 9 9 2
11 0 0 9 11 11 7 10 9 13 13 2
19 9 11 11 13 9 9 1 9 11 2 7 1 9 9 0 9 1 11 2
39 1 9 11 2 16 13 1 9 13 2 11 13 2 16 16 4 3 13 13 2 3 3 1 9 9 2 7 1 9 2 16 13 3 1 9 0 15 13 2
26 9 11 7 9 9 11 11 3 13 2 16 9 0 9 13 3 0 2 3 15 9 1 10 9 13 2
22 13 2 16 1 9 1 9 2 15 11 13 2 13 13 9 0 9 9 1 12 12 2
31 1 9 2 16 1 0 9 13 0 9 7 13 1 9 9 11 2 13 2 2 13 15 2 16 1 15 4 13 3 3 2
10 7 10 0 9 10 9 13 3 9 2
5 2 3 1 9 12
1 3
13 11 2 11 9 13 13 0 9 9 11 11 9 2
19 0 9 9 13 2 16 1 15 13 1 9 0 9 9 1 0 9 9 2
27 9 1 9 13 0 9 11 1 9 9 2 15 13 2 16 11 15 4 13 1 12 5 0 9 1 9 2
5 0 9 13 11 9
2 9 2
35 0 9 1 3 16 12 9 9 2 15 13 9 0 0 9 9 1 0 0 9 2 13 1 9 0 2 0 9 1 0 9 1 9 9 2
10 9 13 13 1 0 9 0 0 9 2
20 1 9 9 9 11 11 15 1 10 9 13 9 3 12 9 3 0 0 9 2
15 15 13 9 13 9 9 1 9 9 1 9 12 9 9 2
9 0 9 9 13 12 9 1 9 2
11 9 0 0 9 11 13 1 3 12 9 2
19 3 13 2 0 0 9 13 0 13 3 9 1 3 0 0 9 1 11 2
19 9 9 13 12 0 9 1 9 1 12 9 2 15 13 14 12 9 9 2
4 1 11 13 9
3 0 11 2
21 1 0 9 11 0 11 1 11 2 15 4 13 1 0 9 2 13 3 15 9 2
22 1 0 9 9 4 13 12 9 10 9 1 0 9 12 9 9 1 0 9 12 9 2
8 1 9 0 9 11 3 13 2
8 0 9 13 11 1 0 9 2
31 9 0 9 1 0 9 2 1 9 9 7 1 0 9 9 2 12 0 0 9 7 0 0 9 13 3 3 12 9 9 2
15 3 13 0 9 1 0 9 12 9 9 9 1 0 9 2
2 9 13
2 11 2
20 9 0 9 1 0 9 7 0 9 15 3 13 1 0 9 1 0 12 9 2
20 1 0 0 9 15 9 3 3 1 9 13 1 12 0 9 7 12 0 9 2
18 9 3 13 1 0 9 12 9 7 1 9 4 10 9 13 7 3 2
18 0 9 0 9 9 13 1 9 0 9 1 9 1 11 7 9 9 2
7 11 1 9 2 7 9 13
2 11 2
21 1 0 9 13 0 9 9 11 11 9 12 7 12 9 9 1 9 12 9 9 2
32 1 9 11 11 15 1 0 9 13 3 0 0 9 1 9 0 1 0 9 7 3 0 9 1 0 11 1 9 12 9 9 2
35 9 9 0 9 0 11 11 2 3 11 13 3 12 5 1 0 9 1 0 9 9 13 9 1 9 9 7 9 9 7 13 3 9 9 2
18 11 13 0 7 0 9 7 10 9 15 1 9 3 13 1 12 9 2
4 11 13 0 9
2 11 2
42 0 9 11 2 0 1 0 9 0 9 2 13 1 9 1 9 10 9 1 0 0 9 1 11 1 11 1 3 16 12 9 1 12 9 2 15 13 3 16 0 9 2
24 9 11 13 3 13 9 9 7 13 9 9 1 0 12 9 1 12 9 3 1 9 0 9 2
22 1 9 10 9 4 15 13 13 7 3 13 9 10 9 7 10 0 9 1 0 9 2
27 9 9 15 1 0 9 3 13 1 12 9 2 10 0 9 1 0 9 13 12 7 0 12 9 1 9 2
5 0 2 11 9 13
7 1 9 11 1 12 9 9
4 3 12 0 9
4 11 1 11 2
28 0 9 0 9 0 2 11 11 4 13 1 0 9 13 12 9 9 2 15 1 9 12 13 9 1 12 9 2
19 3 9 13 1 9 9 1 9 9 12 2 3 4 13 12 9 1 9 2
25 9 1 0 9 7 9 13 12 9 9 2 15 13 1 9 9 1 12 9 3 16 1 9 12 2
25 9 9 4 1 15 13 9 9 1 11 1 12 9 2 9 9 1 11 7 9 9 1 0 9 2
22 3 1 0 9 9 13 0 9 9 1 9 9 2 15 13 9 9 1 12 9 9 2
22 9 0 9 1 9 1 0 9 13 12 9 9 2 1 11 13 9 1 12 9 9 2
12 9 1 0 2 3 0 9 13 12 9 9 2
15 0 0 9 2 3 9 2 15 1 9 13 12 9 9 2
20 0 2 11 1 0 9 13 1 9 11 1 12 9 9 1 9 9 7 9 2
16 1 9 1 9 13 7 0 9 1 0 9 2 0 9 0 2
19 9 9 4 13 3 1 0 9 7 9 0 1 9 11 7 10 0 9 2
17 16 13 1 0 0 9 2 9 9 1 15 3 13 0 9 9 2
19 9 9 13 1 9 2 16 3 4 1 9 13 12 0 7 3 0 9 2
23 9 15 7 1 10 9 13 0 0 9 14 1 0 9 2 7 3 1 9 9 7 9 2
14 1 0 9 4 15 13 10 9 13 1 9 9 9 2
11 3 15 3 13 1 9 9 1 12 9 2
21 0 9 9 4 1 0 9 3 13 9 9 1 9 12 9 9 1 12 9 9 2
9 1 0 9 9 13 3 12 9 2
11 0 2 11 4 13 1 0 9 0 9 2
24 0 9 13 12 9 9 2 16 1 12 9 13 0 0 9 2 9 0 0 7 11 0 9 2
8 0 9 13 3 12 9 9 2
11 9 9 13 9 1 9 9 7 0 9 2
15 9 0 2 11 11 4 1 9 0 9 13 1 0 9 2
18 1 9 3 13 12 9 2 9 1 0 9 13 12 7 9 12 9 2
8 0 9 11 13 1 9 9 9
2 11 2
24 1 9 9 15 13 9 13 3 12 9 0 9 0 9 11 2 15 13 9 0 9 9 9 2
16 0 0 9 0 9 13 1 9 10 0 9 1 12 9 9 2
10 0 9 13 14 14 12 1 12 9 2
18 9 9 2 10 0 9 13 12 9 2 4 1 9 13 1 12 9 2
26 9 9 15 1 9 9 13 2 9 1 9 0 9 2 15 3 13 13 0 9 9 1 0 9 2 2
21 9 9 13 0 1 9 0 9 2 0 0 9 0 11 7 1 0 9 9 11 2
11 0 9 9 1 9 4 13 12 9 9 2
16 0 9 9 9 13 9 1 0 9 2 15 13 12 9 9 2
20 0 9 0 9 2 15 13 9 9 1 9 11 2 4 13 1 9 9 12 2
17 9 11 1 9 13 9 9 12 2 16 10 9 13 9 1 9 2
22 1 12 9 9 15 3 13 0 9 7 10 9 15 1 9 0 9 11 11 13 13 2
3 9 0 9
5 14 2 0 9 2
2 11 2
18 0 0 9 13 1 0 9 9 7 1 9 13 0 9 9 1 9 2
11 9 11 15 13 0 9 11 2 11 11 2
22 13 13 3 1 0 9 1 9 2 7 9 11 15 13 1 9 9 7 0 9 9 2
17 0 9 4 9 9 13 9 15 9 2 0 1 11 1 9 9 2
13 1 0 9 13 9 9 13 9 1 0 9 9 2
24 2 0 9 1 10 9 13 0 9 11 11 1 9 2 15 13 0 9 7 13 10 0 9 2
17 13 15 7 3 3 13 1 9 7 10 9 13 2 2 13 11 2
36 1 9 2 16 11 13 1 11 1 0 9 1 9 9 9 12 2 12 9 11 13 2 16 15 1 15 3 13 13 2 16 0 9 4 13 2
12 9 13 1 11 1 9 9 9 2 11 1 11
11 0 9 13 1 9 2 9 9 13 9 2
7 0 12 9 13 13 9 2
5 14 2 0 9 2
2 11 2
11 0 9 13 1 0 9 9 12 9 9 2
10 0 9 9 13 3 16 12 9 9 2
22 3 0 9 1 9 1 9 13 1 0 9 11 11 13 0 3 0 9 9 1 9 2
26 1 9 1 9 9 11 9 2 15 13 9 12 9 9 2 4 1 0 12 9 13 0 9 9 9 2
17 0 9 9 2 15 4 13 1 0 9 0 9 2 13 3 9 2
14 1 0 9 12 9 9 13 3 3 12 1 9 9 2
16 9 11 13 2 16 13 3 12 9 2 16 13 1 9 9 2
9 0 9 0 9 13 12 9 9 2
9 9 9 13 1 0 12 1 12 2
16 9 13 12 0 9 1 0 9 7 13 0 0 9 1 9 2
20 1 0 0 9 15 13 12 9 7 1 9 9 13 1 11 1 12 2 9 2
21 0 9 13 1 12 2 9 1 0 9 11 7 0 0 0 9 1 9 9 9 2
11 1 0 9 9 13 3 14 1 9 9 2
30 1 9 12 13 15 9 1 0 9 1 9 2 9 9 1 12 9 1 12 9 2 7 9 15 13 13 1 0 9 2
16 1 15 13 7 9 9 2 15 13 0 9 3 12 9 9 2
25 9 0 9 7 9 9 0 9 7 9 15 3 13 9 7 9 13 13 0 7 3 13 10 9 2
25 16 9 9 15 1 9 9 11 13 7 0 9 1 0 9 9 7 1 9 13 3 1 0 9 2
22 0 9 15 13 13 7 1 0 9 7 10 9 13 3 1 0 9 7 1 0 9 2
34 1 0 9 15 13 3 1 0 9 1 9 0 9 2 0 9 2 9 9 11 2 7 0 9 2 9 0 9 1 11 0 11 2 2
19 0 9 15 13 13 7 0 9 1 9 0 9 2 9 11 7 0 9 2
7 13 4 7 9 0 9 2
12 1 9 13 0 7 9 0 9 7 9 9 2
3 0 9 13
8 0 9 4 13 3 1 0 9
4 0 9 15 13
24 1 0 9 4 1 0 9 13 3 12 9 1 9 2 15 13 12 7 3 16 1 9 0 2
22 1 0 0 9 13 9 9 2 16 9 4 3 13 7 4 15 13 7 9 10 9 2
22 1 9 9 9 2 15 10 9 13 9 0 9 2 4 1 9 12 13 3 12 9 2
10 1 9 12 15 10 9 13 3 3 2
18 9 1 9 15 7 13 1 9 9 0 2 7 13 3 0 0 9 2
27 14 12 9 0 9 3 13 0 9 7 9 1 9 0 2 16 15 3 13 9 0 0 9 7 0 9 2
16 16 1 9 12 13 10 9 12 9 2 3 3 3 12 9 2
20 1 9 13 15 9 0 9 0 9 2 10 0 9 15 13 13 0 9 9 2
11 0 9 13 0 9 9 2 3 0 9 2
9 0 9 4 13 3 1 0 9 2
22 1 0 13 3 9 11 2 11 11 2 11 11 2 9 11 2 11 2 0 9 11 2
8 9 9 13 3 9 9 9 2
18 3 13 9 0 9 1 9 9 1 15 3 0 7 13 0 12 9 2
22 1 3 12 0 9 1 9 13 1 9 1 9 0 9 13 12 9 2 3 12 9 2
37 7 13 1 9 9 0 3 13 9 0 9 7 13 9 12 2 12 9 2 1 9 7 9 1 9 13 9 0 9 1 9 7 13 0 9 9 2
8 9 1 9 4 3 13 12 2
18 0 9 4 13 12 9 2 1 15 13 1 0 7 0 7 0 9 2
14 1 3 0 9 13 3 13 10 9 1 9 1 9 2
21 0 9 9 4 1 9 9 13 1 0 0 9 2 3 1 11 2 11 7 11 2
17 9 13 9 15 9 1 9 9 7 0 9 2 9 7 0 9 2
6 9 13 3 16 0 9
13 9 1 9 1 0 7 0 9 15 1 9 12 13
34 0 0 0 9 15 1 9 12 13 1 9 12 1 12 0 9 1 9 9 2 1 12 9 1 9 9 7 1 12 9 1 9 9 2
25 9 9 9 13 0 16 9 9 0 9 2 16 0 9 0 0 0 9 15 13 1 15 9 9 2
13 13 15 9 1 9 1 0 9 7 9 1 9 2
12 3 13 0 9 2 15 15 3 13 0 9 2
13 9 9 0 9 13 3 0 7 10 0 9 13 2
19 1 9 3 0 15 3 13 9 0 9 7 13 15 9 9 9 9 0 2
26 0 0 9 9 13 1 9 7 0 0 9 9 2 0 9 9 0 9 13 9 9 9 2 3 9 2
66 0 0 9 0 1 0 9 13 1 9 12 1 9 12 1 12 0 9 1 9 9 2 1 12 9 1 9 9 2 1 12 9 1 9 9 2 1 9 1 9 7 0 9 1 12 9 2 1 9 1 9 3 1 12 9 7 1 9 9 1 0 9 1 12 9 2
10 9 13 3 13 9 1 9 7 9 2
29 1 9 9 7 9 15 9 9 1 9 7 9 1 9 12 1 9 12 13 7 13 12 5 2 3 2 12 5 2
16 1 9 9 1 9 12 13 1 12 0 9 7 13 12 5 2
23 1 9 9 1 9 9 3 0 9 13 3 9 10 9 2 15 13 13 7 13 0 9 2
17 9 13 9 15 9 1 9 9 7 0 9 2 9 7 0 9 2
10 9 9 13 9 9 1 0 9 9 2
11 15 9 3 3 13 9 0 9 7 9 2
41 0 9 1 9 13 1 9 9 1 9 12 1 9 12 1 12 0 9 2 1 9 9 1 12 9 3 1 9 0 9 1 9 7 9 2 0 0 9 7 9 2
11 1 9 9 13 10 9 3 1 12 9 2
34 9 9 2 15 15 9 1 9 12 13 1 0 0 9 10 9 2 15 13 1 9 1 9 7 9 7 3 1 9 2 9 7 9 2
12 10 9 1 0 0 9 13 1 15 9 9 2
6 0 9 15 13 1 11
2 11 2
32 1 12 2 1 12 2 9 15 1 11 13 0 9 0 9 1 9 3 12 9 0 9 7 0 9 1 11 7 0 9 0 2
20 9 10 9 13 0 9 9 7 9 1 0 9 2 9 2 9 7 0 9 2
56 1 0 9 13 1 10 9 9 9 11 11 2 9 9 11 11 2 9 0 0 9 11 11 2 9 9 7 9 11 11 2 9 9 7 0 9 11 11 2 9 1 9 11 11 2 9 9 11 11 7 9 0 9 11 11 2
4 0 9 13 9
2 11 2
23 0 9 0 0 9 15 3 13 1 12 9 1 12 7 10 0 9 7 9 9 15 13 2
10 13 15 0 9 0 9 1 0 9 2
24 9 0 9 13 1 12 1 9 12 1 12 3 7 1 9 1 15 13 7 9 1 12 9 2
23 0 9 9 15 7 13 2 16 0 9 13 1 3 12 0 9 9 2 13 15 1 9 2
27 1 0 9 9 13 1 0 9 2 3 15 9 9 3 16 13 2 16 0 9 1 9 13 9 0 9 2
29 3 3 15 3 9 9 13 1 0 12 9 2 16 15 1 0 9 1 9 13 0 9 2 7 9 13 3 3 2
25 1 0 9 0 9 15 7 3 13 0 9 0 9 0 9 2 16 10 9 1 0 9 3 13 2
7 0 9 1 0 2 11 2
18 0 9 13 9 10 0 9 1 12 0 0 9 2 0 11 7 11 2
27 9 0 9 13 12 9 9 7 9 1 9 10 9 13 3 16 12 9 9 0 11 2 7 12 9 9 2
6 13 15 0 0 11 2
25 0 9 4 9 0 9 13 13 1 9 12 9 1 9 7 0 9 4 13 13 1 12 0 9 2
5 13 15 14 3 0
29 0 9 9 2 15 4 3 13 16 9 0 9 2 13 3 3 13 1 9 10 9 2 9 2 3 9 3 0 2
18 1 15 13 15 0 2 10 0 9 4 7 3 13 7 1 0 9 2
8 15 13 1 10 9 3 0 2
12 1 0 9 9 13 15 3 9 14 3 3 2
7 3 15 15 15 3 13 2
20 13 2 14 15 14 2 9 13 9 2 1 15 13 0 2 13 15 3 0 2
16 13 7 12 9 2 1 9 14 7 1 15 2 3 0 9 2
19 7 13 3 9 2 1 15 13 9 14 16 15 0 2 1 9 0 0 2
12 13 3 10 9 2 16 4 1 10 9 13 2
19 3 13 13 2 16 9 13 15 14 3 0 13 16 0 9 1 0 9 2
28 1 0 9 13 0 9 13 3 3 1 10 9 7 9 7 3 3 13 7 1 0 9 2 7 15 3 0 2
20 13 1 15 7 9 9 0 9 2 1 15 15 1 9 10 0 9 9 13 2
18 13 10 9 2 15 15 13 9 2 9 10 9 13 3 14 3 0 2
9 13 14 3 0 9 1 10 9 2
18 9 1 0 9 13 3 1 15 0 2 7 15 15 14 3 3 13 2
9 13 15 1 9 13 14 10 9 2
11 1 15 10 9 4 13 0 9 14 13 2
18 13 15 2 16 4 3 13 9 9 9 7 3 9 9 10 9 13 2
17 1 9 15 13 14 3 0 13 9 9 13 3 1 0 9 3 2
24 9 14 13 3 9 2 7 1 9 1 9 3 13 9 9 1 0 9 2 1 9 0 9 2
21 3 13 9 14 1 9 1 0 9 2 15 15 1 15 13 0 0 7 0 9 2
26 9 14 7 15 13 9 9 2 13 9 9 14 1 9 2 13 14 1 9 2 13 15 14 1 9 2
9 13 15 1 9 1 9 14 3 2
23 9 10 9 0 9 1 15 4 3 13 15 2 16 15 9 14 3 1 0 9 3 13 2
8 7 9 12 9 10 9 13 2
21 16 13 2 16 0 9 14 3 13 13 15 3 2 3 4 13 9 1 15 13 2
25 1 15 9 2 15 4 1 9 14 3 13 2 13 14 1 9 9 2 7 7 1 10 0 9 2
9 7 13 13 10 9 1 9 0 2
19 7 16 4 15 3 13 2 13 9 2 3 4 13 14 3 1 9 13 2
18 10 9 0 9 13 0 9 2 16 9 14 3 13 1 9 1 9 2
13 13 15 3 0 2 16 15 1 0 9 13 3 2
35 1 9 0 9 2 12 2 12 2 7 13 13 7 1 15 13 13 2 16 7 1 9 13 3 3 1 0 9 9 2 15 15 3 13 2
12 13 2 16 4 13 13 1 9 3 3 0 2
19 1 10 9 12 9 15 0 9 3 13 1 0 9 2 16 15 3 13 2
20 3 4 13 13 1 0 9 2 16 14 13 1 9 1 9 0 9 2 9 2
9 7 13 15 9 1 0 0 9 2
10 14 9 4 13 13 1 9 12 9 2
26 7 3 9 10 9 1 9 14 3 13 3 3 0 2 10 9 4 15 13 13 1 10 9 1 9 2
10 1 0 9 13 13 1 0 9 9 2
3 16 13 9
20 0 9 9 9 2 16 13 16 3 0 9 0 9 2 13 1 0 9 9 2
35 3 0 9 0 9 1 9 0 9 7 9 2 3 15 0 9 0 2 0 0 9 7 0 0 9 7 13 1 9 1 15 0 9 2 2
25 3 1 9 0 11 2 3 1 10 0 9 2 13 10 12 9 0 9 3 9 1 9 0 9 2
14 1 0 9 3 13 13 0 9 9 9 1 0 9 2
23 9 2 15 15 13 1 0 9 13 0 9 1 12 9 9 2 15 13 13 10 0 9 2
18 1 9 13 9 9 2 1 0 9 0 2 1 0 9 0 9 9 2
12 0 9 9 13 13 1 0 9 2 9 2 2
15 9 9 15 13 1 11 1 11 1 11 7 3 1 9 2
20 0 9 2 3 9 2 13 13 15 9 2 13 1 9 12 1 11 1 11 2
17 13 15 12 12 9 9 7 10 3 0 9 3 13 1 10 0 2
15 9 13 1 0 9 2 13 3 7 14 1 12 9 13 2
16 13 3 0 3 2 7 1 15 0 9 4 13 13 3 3 2
11 9 13 0 2 1 9 13 13 9 9 2
13 1 0 9 13 9 1 9 12 1 12 0 9 2
7 3 13 3 0 9 9 2
21 14 1 0 9 1 9 0 9 0 13 0 9 2 9 13 13 14 9 2 2 2
29 0 9 9 2 15 13 1 9 9 2 9 2 9 2 9 9 7 0 9 7 9 2 13 1 0 9 0 9 2
24 9 15 1 9 3 13 3 16 9 15 2 9 9 9 1 9 9 13 3 9 3 1 9 2
14 9 0 9 9 9 2 7 9 2 13 3 7 3 2
8 9 3 3 13 2 3 13 2
28 16 4 1 15 15 13 2 3 13 9 9 7 9 2 13 15 9 2 9 15 13 1 9 2 13 3 0 2
19 9 2 16 13 9 2 9 7 0 9 2 3 13 1 9 1 0 9 2
45 13 4 15 2 16 9 13 0 2 3 13 3 9 7 10 9 1 0 9 2 13 1 9 13 2 16 15 13 1 0 9 2 9 9 2 9 0 9 2 0 9 3 2 2 2
15 13 7 4 13 1 9 9 2 16 13 3 0 15 13 2
13 13 9 13 3 7 1 0 9 0 9 1 9 2
9 9 3 13 1 12 7 12 9 2
21 9 15 13 14 3 2 3 1 9 0 2 9 2 0 9 2 0 9 0 2 2
12 9 13 3 1 9 1 9 2 1 9 9 2
13 0 13 0 9 2 9 0 2 9 2 9 2 2
31 9 9 2 11 2 13 3 13 1 0 9 2 1 12 9 2 0 2 0 9 1 0 9 2 7 15 13 9 7 11 2
9 0 13 0 9 7 9 0 9 2
15 7 0 9 9 3 13 1 9 9 7 9 1 9 9 2
28 16 9 1 0 9 13 13 9 9 2 13 3 0 2 16 9 13 3 9 1 9 7 13 1 10 9 3 2
13 9 1 9 4 13 0 9 2 3 1 9 0 2
16 3 13 14 1 9 2 1 9 0 2 0 9 1 10 9 2
10 0 9 3 14 13 15 15 0 9 2
11 9 13 0 9 2 7 9 9 2 9 2
3 9 1 9
15 1 9 1 0 9 7 9 13 3 12 9 13 9 1 9
38 3 1 10 9 2 3 13 1 0 0 9 0 11 9 1 9 11 11 0 9 0 11 2 13 1 9 7 0 9 1 11 9 9 10 9 11 11 2
9 9 1 0 11 9 4 3 13 2
5 16 3 3 15 2
14 1 9 10 1 15 3 12 9 0 9 13 0 9 2
15 1 12 9 4 13 11 7 11 1 9 7 9 0 9 2
34 13 15 2 16 13 2 16 10 9 13 7 9 9 2 16 3 9 0 11 7 9 9 9 2 3 13 9 2 2 13 15 9 11 2
10 15 15 13 2 13 1 9 11 11 2
23 3 2 13 15 2 16 3 13 9 2 3 13 0 13 3 1 9 7 1 9 10 9 2
14 1 9 13 0 13 9 1 12 9 3 1 0 9 2
27 13 15 0 2 16 15 2 15 13 3 13 9 1 9 0 3 0 9 2 10 9 1 0 9 3 13 2
17 0 9 11 2 1 15 13 0 9 2 13 9 0 9 1 9 2
24 13 15 1 10 9 15 1 9 0 0 9 2 15 13 1 12 9 9 1 11 7 1 9 2
21 11 3 13 7 3 13 9 1 0 2 0 9 3 0 0 2 1 9 0 9 2
12 10 0 9 1 3 16 9 9 13 0 9 2
30 1 0 9 9 11 11 3 2 13 2 16 9 13 13 14 15 2 15 9 13 13 2 7 3 15 2 15 4 13 2
15 0 14 13 9 2 16 4 13 2 15 13 13 7 13 2
45 15 1 0 3 7 3 0 11 2 3 3 2 9 9 11 13 2 16 0 0 9 4 13 3 7 2 16 15 15 9 13 2 7 3 15 15 13 13 13 9 2 13 3 3 2
13 1 0 0 9 4 7 11 13 1 3 0 9 2
24 3 7 2 16 4 3 13 1 0 9 2 7 3 7 2 16 0 9 1 0 11 13 0 2
14 10 9 3 13 7 15 0 9 1 9 2 9 0 2
17 9 11 15 3 13 13 9 7 9 2 15 3 3 13 0 9 2
15 13 13 3 9 2 15 1 11 13 13 16 9 1 9 2
21 0 9 1 9 2 3 2 9 9 2 13 11 9 1 9 1 9 0 9 11 2
37 13 9 3 3 16 9 0 9 2 1 15 15 3 13 0 0 9 7 9 2 11 2 0 11 2 0 0 2 0 11 2 0 11 2 0 11 2
6 15 10 9 13 0 9
20 1 9 7 9 13 3 1 9 2 1 9 1 0 11 9 2 3 0 9 2
44 3 3 1 9 11 11 2 11 2 9 2 1 15 9 2 0 1 9 12 1 0 11 2 9 2 9 7 9 2 1 9 0 1 9 7 10 0 9 13 9 1 0 9 2
32 1 9 15 13 0 9 11 11 2 15 1 9 12 13 1 11 2 1 0 9 1 9 11 11 2 15 10 9 13 0 9 2
40 0 2 3 1 3 0 9 3 0 0 9 13 12 2 9 2 0 0 9 11 2 11 11 13 9 1 10 3 0 9 1 0 9 1 9 12 0 9 9 2
5 3 13 10 9 2
3 9 1 9
38 0 9 1 12 9 3 13 11 9 9 2 1 9 1 9 9 11 2 11 2 11 2 11 2 11 7 11 2 11 13 3 0 9 1 9 11 11 2
32 1 9 9 1 9 9 3 1 9 0 7 0 13 0 9 7 0 9 1 9 3 0 7 0 2 0 9 7 9 1 9 2
5 11 7 9 1 11
29 0 9 9 13 9 1 9 9 2 9 2 9 1 9 2 0 9 1 0 9 9 7 9 1 0 9 1 11 2
18 1 0 9 13 13 9 0 9 1 0 7 0 9 2 1 9 9 2
15 1 9 3 13 13 1 0 0 11 7 13 9 1 11 2
10 1 9 0 9 13 13 3 0 9 2
3 9 2 9
17 1 9 2 9 2 13 2 14 2 15 13 13 1 0 0 9 2
10 15 15 4 13 3 2 15 15 3 2
28 9 9 0 0 2 0 9 1 0 9 13 3 12 2 9 1 12 1 12 9 7 1 0 9 12 2 9 2
9 1 12 9 1 11 9 1 11 2
16 1 9 13 1 9 1 12 12 9 2 9 2 9 7 9 2
9 1 9 9 12 9 9 7 9 2
3 9 3 2
17 9 0 0 9 2 15 13 9 0 11 9 11 11 2 13 0 2
16 7 0 9 13 3 1 9 9 2 0 9 7 0 0 9 2
23 1 9 0 9 11 13 9 1 9 1 0 9 2 9 2 9 13 1 9 1 12 9 2
17 0 9 13 3 0 2 7 1 9 10 9 4 13 13 7 3 2
8 9 1 9 1 11 13 13 2
19 7 10 9 13 13 9 1 0 9 2 1 15 13 0 9 1 9 0 2
1 9
3 15 13 9
22 9 9 11 3 13 0 9 16 9 9 1 9 0 9 1 9 2 3 7 3 13 2
54 13 2 0 2 0 2 16 4 13 2 16 3 9 2 1 9 1 12 9 2 0 0 9 2 0 2 0 2 0 9 1 0 9 2 1 9 0 9 0 1 0 9 7 9 7 2 3 4 3 13 13 3 2 2
13 13 1 9 0 9 2 2 2 7 13 15 9 2
15 1 11 1 11 13 9 1 9 1 10 0 7 0 9 2
53 16 1 0 9 15 9 13 2 3 3 13 1 9 2 13 2 14 3 15 9 1 9 13 2 16 0 9 13 3 1 0 9 1 0 9 2 9 1 11 13 1 9 0 9 7 1 10 9 0 7 0 9 2
4 13 15 3 2
2 3 2
6 9 9 2 9 9 2
18 0 9 13 1 15 2 16 16 3 9 0 9 13 2 13 15 3 2
4 9 3 13 2
69 12 9 2 7 3 3 13 2 3 2 16 1 9 2 9 2 13 7 12 0 9 2 3 0 2 7 0 2 2 3 12 9 1 0 9 13 1 9 7 1 10 0 9 2 3 1 9 1 9 0 7 0 2 1 9 0 1 0 2 0 9 13 0 2 0 9 13 9 2
20 9 1 9 1 9 1 12 9 7 9 7 9 1 9 0 3 3 13 0 2
13 9 15 13 12 1 0 3 1 0 0 9 9 2
42 10 0 9 1 10 9 13 3 0 9 1 9 2 13 15 9 1 9 7 3 13 9 1 9 1 9 7 0 9 2 2 3 3 15 3 13 2 13 3 9 2 2
12 7 3 2 1 9 15 13 0 2 0 9 2
13 9 9 0 10 0 0 9 15 13 1 0 9 2
3 13 9 2
66 3 4 13 1 0 9 7 1 10 0 9 13 9 10 9 0 0 9 2 2 1 15 13 2 15 13 2 15 13 2 9 2 1 15 2 1 15 15 15 13 2 13 14 9 2 13 9 2 13 2 9 2 15 13 13 2 6 15 13 2 13 15 2 9 2 2
31 0 9 13 9 2 7 14 0 2 6 2 7 9 2 15 13 9 7 9 2 13 15 9 9 2 2 0 2 0 2 2
10 9 1 0 9 0 9 4 3 13 2
10 13 15 9 2 12 9 1 12 9 2
19 15 13 13 7 0 9 2 9 1 9 3 1 0 9 2 3 3 13 2
10 3 15 15 15 3 3 0 3 13 2
5 3 13 0 9 2
15 2 9 2 2 15 3 13 0 0 0 2 13 1 9 2
8 11 1 11 13 3 3 9 2
8 1 9 15 13 1 9 11 2
5 0 16 0 9 2
10 0 0 9 1 9 9 9 13 3 2
9 6 2 16 9 13 1 10 9 2
8 6 2 16 13 11 1 9 2
9 1 9 13 7 9 2 7 9 2
17 15 15 7 3 13 1 0 9 2 16 15 13 2 1 15 2 2
8 7 9 13 2 2 1 15 2
3 2 11 11
6 0 9 9 9 7 9
44 2 9 7 9 2 2 13 9 11 10 9 11 1 0 0 9 2 2 9 7 9 4 15 13 9 15 2 3 4 15 13 3 13 0 9 2 7 13 2 16 13 15 0 2
13 13 15 2 0 9 4 15 13 7 1 0 9 2
9 13 15 2 13 15 3 13 9 2
6 13 15 3 13 9 2
10 13 4 1 0 9 13 10 9 2 2
17 7 9 2 13 9 2 7 9 4 15 13 13 9 1 0 9 2
19 3 14 7 14 2 16 0 9 13 13 1 15 2 7 3 1 10 9 2
10 0 11 15 13 1 0 2 16 3 2
16 13 3 1 0 9 0 9 2 14 7 3 1 10 0 9 2
20 0 0 9 13 1 0 9 3 0 16 0 2 7 9 15 1 15 13 3 2
37 9 3 13 0 9 0 7 0 9 2 11 2 2 15 13 0 2 9 2 15 13 0 2 9 2 2 7 3 1 9 13 1 10 9 0 9 2
22 9 15 3 13 1 9 12 2 9 2 3 15 9 13 9 0 9 1 9 0 9 2
37 0 9 0 9 2 0 0 9 2 13 0 9 9 0 9 1 0 9 2 9 2 1 15 2 0 9 2 13 1 9 2 15 13 1 10 9 2
5 9 0 7 0 9
34 3 7 3 3 0 9 13 0 9 13 1 9 9 10 0 9 0 9 1 0 9 2 9 7 0 0 9 2 9 13 9 9 2 2
18 0 9 13 1 9 16 12 1 10 0 0 9 9 0 7 0 9 2
20 9 12 10 9 15 1 9 1 0 9 13 3 0 9 2 3 3 3 9 2
18 0 9 9 13 3 0 9 1 9 9 7 9 9 7 0 0 9 2
30 9 2 0 1 9 16 9 1 9 2 13 1 0 9 3 2 3 1 15 15 7 13 0 9 0 9 9 7 9 2
27 1 10 9 13 9 1 9 9 3 1 15 9 9 2 16 1 0 11 2 7 7 1 0 0 0 9 2
33 9 12 15 0 9 11 13 1 9 10 0 0 9 2 1 15 3 9 13 9 2 13 9 7 13 9 0 1 9 1 0 9 2
24 0 9 9 11 2 0 9 2 12 1 0 9 1 11 2 13 0 9 9 7 0 0 9 2
19 9 9 0 9 1 9 13 10 9 2 7 4 3 13 14 1 0 9 2
2 0 9
20 0 9 3 13 9 2 0 9 2 12 1 9 11 12 2 11 7 9 11 2
26 0 15 1 10 9 13 0 9 1 9 2 13 3 2 3 0 9 2 7 0 9 13 3 13 9 2
12 1 9 15 7 0 9 13 3 16 9 9 2
41 9 0 7 0 9 13 7 0 9 1 0 11 2 9 0 9 15 13 1 9 9 7 0 9 13 0 1 15 2 15 4 3 3 13 16 2 0 0 9 2 2
21 9 9 11 1 15 2 16 0 9 13 1 9 16 1 10 9 2 13 3 0 2
13 3 0 0 9 15 13 1 9 3 0 16 0 2
27 0 9 13 3 9 11 12 2 9 2 12 7 2 16 4 13 9 7 15 7 9 10 9 2 9 11 2
9 3 15 13 9 1 0 0 9 2
9 0 9 13 7 3 0 0 9 2
3 0 9 9
12 9 9 0 7 0 9 1 15 13 3 0 0
16 9 0 7 0 9 1 0 9 13 10 3 0 9 0 9 2
14 9 9 0 9 1 0 9 15 3 13 1 0 9 2
31 0 9 0 9 7 0 9 2 15 13 0 9 1 10 0 9 2 4 3 3 13 9 0 9 9 7 10 9 1 9 2
27 11 12 2 13 3 9 12 2 16 0 9 9 1 9 13 3 13 9 2 0 9 13 3 1 0 9 2
7 3 4 13 9 0 9 2
12 9 3 13 9 13 15 0 9 1 9 0 2
6 9 13 7 13 9 2
32 9 0 9 16 0 13 3 9 0 2 7 0 2 0 2 15 15 2 13 1 9 1 9 2 2 15 1 0 9 13 9 2
22 9 1 0 9 1 9 13 0 9 1 9 2 16 15 1 9 11 12 2 3 13 2
20 13 0 13 2 16 0 10 9 13 9 2 7 3 13 9 9 7 9 9 2
2 0 9
24 0 9 1 0 9 7 1 9 0 9 13 0 0 9 0 9 7 9 9 1 15 9 9 2
10 3 7 10 9 13 9 1 0 9 2
9 0 9 7 13 10 9 3 3 2
39 2 0 9 3 13 9 9 7 13 9 9 2 1 15 15 13 13 14 9 0 9 2 2 13 3 11 11 12 2 1 0 9 1 12 2 12 2 12 2
24 9 3 3 13 1 9 9 2 1 15 2 0 9 9 9 13 13 7 3 13 9 0 2 2
25 0 9 0 7 0 0 9 15 1 9 0 9 13 16 0 9 2 7 3 16 0 9 0 9 2
17 0 9 2 0 15 1 9 0 9 2 3 13 0 9 0 9 2
17 9 9 13 1 10 9 0 3 2 16 1 9 2 7 1 9 2
15 9 15 3 13 1 9 0 9 2 0 1 9 15 9 2
22 7 15 9 15 3 13 3 0 2 16 13 1 15 10 2 0 2 9 0 7 3 2
11 1 10 0 9 3 13 7 9 0 9 2
48 3 9 12 4 1 0 9 9 13 0 9 9 7 9 2 15 15 0 9 13 0 2 1 0 9 0 9 0 9 2 3 13 2 3 3 4 9 13 3 1 9 10 2 0 9 2 2 2
20 9 11 2 11 1 0 9 11 12 2 7 12 2 0 9 10 9 3 13 2
25 0 9 3 13 1 0 9 3 0 0 9 2 15 7 1 9 13 15 9 1 9 9 1 9 2
16 10 0 9 15 1 10 9 3 2 7 3 3 3 13 3 2
6 0 9 9 7 9 9
21 9 7 9 2 12 3 0 9 2 15 15 3 13 1 0 7 3 1 0 9 2
16 9 2 15 13 10 9 2 15 13 13 0 9 1 0 9 2
31 1 9 9 2 9 1 2 0 9 2 2 1 9 10 9 2 13 1 9 2 3 15 10 0 9 1 0 0 9 13 2
11 3 14 0 9 3 13 1 9 9 9 2
29 9 0 9 11 11 2 12 2 12 2 1 9 12 2 15 13 9 11 2 13 0 9 1 3 0 9 9 9 2
16 10 9 13 1 9 1 0 9 9 7 9 15 1 9 9 2
16 13 1 9 9 13 3 1 11 0 3 1 9 9 9 9 2
12 0 9 10 9 13 11 9 0 9 0 9 2
25 1 0 9 13 1 15 9 9 2 7 9 0 9 1 11 13 13 9 0 9 2 0 0 9 2
6 9 9 9 13 9 2
24 9 1 0 9 9 13 0 9 2 9 0 15 13 1 3 0 9 2 15 13 1 9 0 2
7 9 13 0 9 11 9 2
28 9 2 15 13 13 1 0 9 2 15 13 13 1 0 9 9 2 7 7 0 9 13 1 15 9 7 9 2
10 0 9 15 3 3 13 1 9 0 2
10 9 13 1 11 0 9 1 9 9 2
30 3 1 10 9 15 7 11 13 1 9 9 9 2 3 11 2 2 15 0 9 0 9 7 1 15 0 0 9 13 2
13 9 1 0 0 7 0 0 9 11 14 3 13 2
63 1 0 9 15 3 3 13 12 0 9 2 15 11 13 2 12 2 9 2 15 13 2 16 0 9 0 4 13 1 0 9 7 9 0 9 2 7 12 2 9 2 15 13 1 9 11 1 11 2 1 15 13 4 9 0 9 13 0 9 1 0 9 2
13 3 7 1 9 1 15 13 12 0 9 1 9 2
21 0 9 13 2 16 15 9 13 1 0 9 2 3 3 2 16 9 13 0 9 2
18 1 15 15 13 7 3 0 9 2 1 15 9 13 14 1 9 9 2
9 0 9 9 0 9 13 11 3 2
33 1 9 0 0 9 15 1 9 9 13 3 13 0 9 2 16 1 0 9 9 13 14 1 9 2 15 9 9 13 9 0 9 2
9 0 9 1 0 9 13 9 9 2
26 15 3 15 0 9 13 9 0 9 7 0 9 2 0 9 7 13 7 13 1 15 3 0 9 9 2
18 9 1 9 1 9 4 7 13 9 1 9 2 1 3 0 9 9 2
8 12 9 15 7 11 13 13 2
14 0 9 9 9 13 1 0 9 7 9 9 16 15 2
29 3 0 9 0 9 0 9 13 2 16 9 9 15 1 9 3 13 2 3 7 7 2 16 9 10 0 9 13 2
15 0 9 0 1 0 3 13 9 2 15 15 9 9 13 2
7 3 7 13 9 9 0 2
21 0 0 9 1 11 13 2 15 13 9 9 2 15 13 9 10 0 9 7 9 2
17 0 9 13 1 9 1 9 0 0 9 1 9 9 0 9 13 2
6 12 0 0 9 1 9
17 3 1 0 9 15 3 13 1 0 9 9 11 11 2 12 2 2
31 7 1 10 9 13 3 9 14 9 2 1 9 13 0 0 9 2 7 7 15 1 10 9 0 13 15 0 14 9 12 2
35 9 15 7 1 0 9 13 9 3 13 2 3 12 9 2 9 0 14 1 9 2 0 9 2 12 9 2 7 9 0 9 2 11 2 2
8 3 1 12 9 12 9 9 2
9 1 10 9 13 13 7 3 9 2
24 13 15 3 1 15 2 1 15 15 1 0 9 13 2 16 13 2 0 2 2 1 0 9 2
18 7 7 2 16 15 3 3 13 9 7 9 1 9 2 9 2 9 2
26 16 15 13 3 9 0 2 14 15 3 13 2 0 2 9 2 13 0 9 0 1 2 0 2 9 2
24 2 0 2 2 0 9 0 9 15 13 1 10 0 2 0 9 3 2 7 3 3 16 3 2
52 1 0 9 0 9 15 1 15 13 2 13 7 13 0 7 0 9 1 0 9 2 9 9 0 9 2 3 16 9 1 0 9 7 9 1 9 2 16 4 4 1 10 9 15 3 2 3 2 13 7 13 2
18 13 15 3 9 2 0 9 2 7 2 9 2 7 10 2 9 2 2
25 14 3 0 9 9 2 15 13 9 14 1 9 0 0 9 7 10 2 9 13 0 1 9 2 2
15 9 13 9 1 9 2 2 15 1 9 13 0 9 2 2
19 9 1 0 9 0 9 13 0 2 7 9 10 9 15 13 14 0 9 2
6 13 7 1 15 0 2
44 1 0 9 3 0 9 2 13 4 1 9 2 3 15 1 10 0 9 13 9 0 0 0 2 0 9 1 10 9 2 3 0 9 7 1 9 9 2 2 13 13 0 9 2
16 9 1 0 2 9 2 9 3 0 9 2 7 10 0 9 2
22 1 0 9 1 0 9 3 0 2 9 2 1 0 9 9 15 13 13 1 10 9 2
15 16 7 3 13 2 9 0 9 2 2 13 3 15 13 2
9 9 9 13 9 2 10 0 9 2
29 1 10 9 15 13 1 2 9 9 2 13 7 1 0 9 2 1 9 2 1 2 9 0 9 2 2 1 9 2
8 15 9 15 13 9 1 9 2
16 7 9 13 7 1 9 2 13 15 1 9 2 13 7 0 2
33 13 0 9 9 0 9 2 0 1 9 12 1 11 2 7 3 0 11 2 1 15 11 3 13 0 9 7 3 1 9 12 13 2
25 1 0 2 3 0 2 7 7 3 0 9 9 13 9 10 9 3 0 9 0 7 1 0 9 2
51 10 9 3 13 1 3 0 2 3 3 0 2 9 9 2 9 9 13 2 9 9 1 9 2 14 1 3 0 9 2 2 13 2 14 9 9 2 0 9 2 7 9 13 9 9 2 1 15 13 2 2
33 7 9 2 3 0 7 3 2 0 2 9 2 15 3 13 13 7 10 0 9 2 2 9 1 0 9 1 9 15 13 9 2 2
18 15 13 7 9 2 0 13 3 0 9 2 0 2 7 2 0 2 2
19 16 16 2 9 1 9 13 10 9 16 9 2 1 9 1 0 9 2 2
13 13 15 3 7 9 1 9 2 1 9 1 15 2
15 1 9 2 1 15 13 2 15 13 3 13 16 15 2 2
30 11 11 3 13 2 16 1 12 1 9 13 0 2 0 9 2 1 2 0 9 0 2 0 2 0 7 3 0 2 2
21 13 3 10 9 13 3 2 7 1 11 15 13 13 7 9 2 1 15 11 13 3
4 3 1 11 11
1 9
38 0 9 1 3 0 9 0 9 11 11 2 12 2 13 9 11 11 2 15 13 0 9 11 0 1 11 3 1 0 9 11 2 0 9 7 0 9 2
17 3 0 9 2 0 12 9 2 13 0 9 3 1 10 9 13 2
27 0 9 9 13 0 9 1 9 7 9 9 2 10 2 9 13 7 13 1 0 9 9 9 7 9 2 2
11 1 0 9 3 7 13 7 9 0 9 2
17 3 0 9 13 0 9 1 9 0 9 2 0 1 11 0 9 2
14 9 1 11 13 0 9 1 0 9 1 10 0 9 2
27 16 4 3 13 10 9 7 9 2 13 0 3 3 13 11 0 9 7 3 15 13 1 9 9 0 9 2
22 13 2 3 7 3 13 0 2 0 9 2 1 15 4 15 13 0 9 0 0 9 2
13 15 13 1 9 13 0 9 1 0 9 10 9 2
26 7 0 9 9 13 0 3 13 1 9 2 0 1 0 9 9 2 15 13 11 0 3 1 0 9 2
25 9 0 1 0 9 0 9 2 1 0 9 10 9 7 1 0 9 13 0 9 7 0 9 9 2
8 1 0 9 13 1 9 0 2
22 0 0 9 3 0 9 13 9 2 15 4 13 10 0 9 9 1 9 2 12 2 2
22 13 0 9 2 9 0 2 0 7 0 2 15 13 1 11 7 1 0 9 0 9 2
16 11 9 7 10 0 0 7 0 9 4 1 9 15 3 13 2
22 9 13 9 9 2 9 2 9 2 9 2 15 15 10 9 13 1 9 9 10 9 2
3 1 0 9
16 11 11 2 0 9 2 9 13 1 9 2 0 9 2 13 2
19 0 0 9 2 0 9 0 1 0 9 9 0 9 2 13 3 3 3 2
38 9 11 11 2 15 15 13 1 9 0 9 1 0 0 9 2 9 13 1 9 0 0 9 2 9 12 2 12 2 2 15 13 9 13 9 1 9 2
8 11 11 2 0 9 7 9 2
31 0 2 0 9 0 9 13 9 9 9 1 9 3 1 9 0 9 16 2 9 9 7 9 1 9 9 7 0 9 2 2
7 1 0 9 13 0 9 2
6 11 11 2 0 9 2
23 0 9 0 9 13 1 9 11 11 7 9 11 11 16 0 2 9 2 0 0 9 9 2
8 11 11 2 11 2 12 9 2
17 0 9 1 0 9 9 11 11 13 0 9 1 9 9 7 9 2
14 9 11 11 2 0 1 9 12 9 2 13 9 9 2
7 11 11 2 9 0 11 2
24 0 9 0 9 11 2 11 1 9 9 11 1 0 9 13 9 0 1 9 1 9 9 9 2
8 13 11 11 2 13 0 9 2
4 9 13 13 0
10 9 3 13 0 2 3 2 13 11 11
23 9 9 1 0 9 0 13 1 10 9 3 3 3 0 9 11 11 9 9 7 0 9 2
15 11 11 10 9 13 7 13 1 15 7 0 9 11 11 2
9 15 15 13 16 0 9 1 9 2
8 13 15 13 3 9 0 9 2
31 3 3 3 9 0 0 0 9 7 1 0 9 0 9 9 10 0 9 11 11 2 1 15 4 13 0 9 1 11 11 2
36 7 1 9 12 15 9 1 11 11 7 11 7 11 0 13 1 9 2 16 9 13 3 0 2 0 9 7 16 13 3 0 15 1 15 13 2
12 13 15 10 9 1 9 1 0 9 10 9 2
2 9 2
5 9 9 9 9 2
14 15 2 16 9 13 0 9 2 2 15 13 9 2 2
29 9 0 1 0 9 2 1 0 9 2 3 15 13 9 0 2 9 0 2 9 7 9 0 7 9 1 0 9 2
13 9 9 13 3 0 2 7 3 10 0 9 9 2
14 13 1 0 9 1 9 2 9 1 9 10 0 9 2
5 13 9 1 9 2
11 9 13 9 0 13 9 2 13 3 0 2
13 10 9 13 3 3 0 9 0 7 0 2 2 2
12 1 11 2 3 9 13 2 13 9 0 9 2
9 7 9 13 0 9 0 0 9 2
7 3 3 1 15 3 13 2
21 9 0 9 15 13 2 16 15 13 9 0 7 16 1 9 0 0 9 9 13 2
23 7 15 2 15 13 9 1 0 7 0 9 2 7 15 13 9 0 2 2 9 3 13 2
36 1 11 2 15 13 9 9 7 3 15 13 0 9 2 13 3 9 9 2 0 9 2 0 9 2 0 9 2 15 15 3 0 9 3 13 2
8 7 9 13 0 3 0 9 2
8 1 0 9 13 9 0 9 2
34 3 13 1 9 3 2 0 2 2 16 15 9 13 1 12 9 1 0 9 2 7 13 1 15 3 3 0 9 16 1 0 2 9 2
11 10 0 9 4 3 13 1 0 9 9 2
8 3 4 15 1 10 9 13 2
23 13 1 15 2 1 0 9 2 9 12 1 9 2 1 0 12 9 2 15 13 3 0 2
19 9 0 9 4 15 13 11 13 1 9 11 2 3 4 3 13 16 9 2
13 3 3 4 13 1 9 10 0 9 1 0 9 2
26 13 3 9 9 2 15 9 3 13 2 0 9 2 7 0 9 9 13 0 10 9 2 7 3 0 2
11 15 13 2 16 13 1 10 0 0 9 2
39 9 0 9 1 0 9 9 2 15 2 16 2 7 3 7 2 16 13 0 2 3 3 13 9 2 9 2 9 7 9 0 9 2 3 1 10 0 9 2
13 13 3 0 13 9 2 9 2 1 9 1 9 2
13 3 13 9 13 1 0 2 0 9 2 2 2 2
17 7 0 9 13 13 0 2 16 13 2 14 0 2 13 1 15 2
10 0 9 13 0 9 7 13 1 9 2
22 16 13 3 11 2 9 13 13 1 9 2 3 9 2 7 13 3 9 2 3 9 2
7 9 13 3 3 9 9 2
11 0 9 9 13 3 0 2 3 13 0 2
12 0 9 7 9 3 13 1 0 9 0 9 2
12 1 15 13 7 0 9 9 2 10 0 9 2
17 13 0 9 3 10 0 9 16 10 2 15 13 1 0 9 9 2
2 3 2
21 1 15 15 13 2 16 9 13 7 3 14 9 2 7 16 13 3 0 9 9 2
12 15 13 3 3 13 1 9 2 15 9 13 2
26 15 11 13 9 9 2 13 15 9 2 9 2 7 13 0 9 0 9 2 15 13 3 1 9 13 2
12 10 9 2 0 15 0 9 9 2 14 13 2
14 3 13 15 3 0 2 16 13 9 1 9 0 9 2
26 13 2 16 1 15 9 13 1 0 9 9 7 9 15 2 1 15 13 9 9 7 1 15 15 13 2
13 13 1 15 3 13 2 16 1 9 10 9 13 2
17 1 0 0 9 0 9 9 13 13 7 13 15 3 3 1 9 2
11 13 3 1 9 7 9 0 9 0 9 2
30 1 15 13 7 9 0 2 0 2 9 0 2 9 3 0 2 9 2 9 7 9 1 9 2 15 13 11 1 11 2
18 9 13 3 13 1 9 2 3 7 0 2 1 9 2 3 1 9 2
18 7 15 1 15 3 3 13 0 9 2 7 3 3 14 14 1 11 2
10 15 13 1 0 9 0 9 1 9 2
12 1 11 11 11 11 2 10 9 13 3 0 2
30 13 15 0 2 3 0 9 7 10 9 16 0 9 9 7 9 7 9 13 15 0 2 15 1 15 4 1 9 13 2
30 11 2 3 15 13 7 13 2 16 13 1 0 9 9 2 13 0 9 16 11 2 13 1 9 9 2 1 9 9 2
18 1 10 9 13 0 0 9 2 10 9 13 14 1 10 9 9 12 2
34 13 3 7 0 0 9 2 9 11 2 11 2 11 2 9 11 2 9 11 7 11 2 3 11 11 2 11 11 2 11 7 11 0 2
19 9 0 9 3 13 2 3 13 9 0 2 10 0 9 3 13 1 9 2
35 13 9 0 2 1 11 7 11 15 13 3 15 2 3 13 13 11 11 2 15 13 1 0 9 1 11 1 11 2 3 13 0 9 11 2
6 13 0 9 1 11 2
24 13 7 0 9 2 7 11 12 2 7 0 14 1 12 10 9 2 15 13 13 1 0 9 2
7 10 9 15 15 3 13 2
17 13 15 10 9 2 15 13 1 0 9 1 9 7 13 0 9 2
16 13 15 13 15 2 16 3 0 9 13 13 13 0 9 9 2
11 14 1 0 9 2 16 0 9 3 13 2
7 9 15 13 13 9 11 2
6 9 3 3 13 0 2
29 15 13 10 0 9 2 16 13 1 9 7 16 9 13 0 2 16 3 13 9 11 2 15 15 7 1 15 13 2
7 13 9 1 9 1 9 2
4 9 13 0 2
14 9 1 0 9 9 13 1 15 2 16 13 0 9 2
19 1 0 9 13 9 0 0 1 9 0 2 7 15 3 1 0 7 0 2
43 7 15 15 13 9 1 0 9 2 1 9 2 9 7 9 2 3 13 11 2 2 9 0 2 1 9 9 2 1 1 15 13 15 2 15 13 0 7 0 9 2 0 2
12 13 7 1 10 9 7 1 9 7 9 9 2
8 9 7 9 7 3 13 9 2
18 9 13 14 0 9 2 2 9 7 9 2 2 3 13 3 11 11 2
9 9 13 0 2 7 3 15 13 2
5 3 13 10 9 2
16 15 4 13 1 0 9 2 16 15 3 15 3 1 9 13 2
11 3 13 0 9 1 0 9 9 11 11 2
30 9 9 2 9 9 2 9 9 15 15 9 9 2 3 1 15 15 13 1 10 9 2 15 15 1 15 13 1 9 2
19 13 3 1 9 0 9 16 1 11 9 2 15 13 1 10 9 3 0 2
17 1 9 13 3 11 11 2 12 1 0 0 9 1 9 0 9 2
19 1 15 15 2 15 13 0 9 11 2 15 13 0 9 2 0 2 0 2
23 3 9 13 9 0 9 2 16 13 11 11 2 15 1 11 1 11 13 0 9 7 9 2
27 1 0 9 15 13 3 1 9 11 1 0 2 11 0 1 11 2 0 9 10 9 1 11 2 16 13 2
7 13 4 10 9 1 11 2
8 13 4 1 15 1 0 9 2
25 16 13 3 11 11 2 13 4 3 9 2 16 4 15 13 2 7 3 4 13 1 10 9 11 2
11 1 10 9 13 14 1 10 9 9 11 2
20 13 1 0 9 11 1 11 0 2 15 13 1 0 9 7 1 0 9 0 2
14 13 4 15 1 0 9 2 0 9 2 9 2 9 2
25 10 9 3 4 14 13 0 9 2 7 4 13 3 2 16 13 1 15 0 9 2 13 0 9 2
8 7 15 13 9 3 3 0 2
16 15 10 9 2 15 13 15 0 1 9 2 15 3 13 9 2
40 16 15 9 3 13 9 2 1 15 13 14 9 9 2 7 13 15 2 16 15 13 1 9 2 7 3 13 10 0 9 2 0 9 2 15 3 13 3 13 2
10 15 13 0 9 9 2 7 3 0 2
10 13 3 13 2 1 15 3 15 13 2
12 13 15 1 9 13 2 16 13 0 9 9 2
10 3 14 2 3 3 3 0 9 9 2
39 11 11 2 12 2 2 9 0 9 7 2 0 2 9 15 13 1 11 1 11 2 7 16 13 3 9 9 0 1 11 2 11 13 1 15 3 3 0 2
12 1 11 9 13 9 7 9 0 9 0 9 2
33 1 9 12 15 13 9 0 9 1 11 2 1 0 9 15 0 9 13 1 11 2 3 15 13 3 13 1 15 0 9 0 9 2
10 9 0 9 13 16 9 1 9 11 2
86 1 0 9 3 13 10 0 7 0 9 2 13 9 2 9 2 9 2 11 2 0 2 11 12 2 0 9 1 0 9 2 2 13 1 9 2 13 9 11 2 13 2 13 2 7 13 0 9 1 10 9 2 3 13 0 9 2 0 9 11 13 1 0 9 1 11 2 3 15 13 1 12 9 7 2 13 2 1 9 2 0 9 1 0 9 2
9 3 15 13 0 2 16 0 9 2
2 9 11
12 13 15 2 16 4 13 4 13 9 0 9 2
5 13 0 9 11 2
18 9 2 0 13 1 15 0 9 2 16 9 13 15 3 0 2 0 2
4 9 3 13 2
10 15 13 1 15 2 16 13 13 0 2
12 13 2 16 16 13 1 9 2 3 0 13 2
4 9 2 14 2
6 15 4 1 15 13 2
5 13 4 15 15 2
4 9 2 14 2
10 9 13 9 10 2 16 15 13 0 2
4 9 2 3 2
9 3 14 7 2 16 12 9 13 2
5 9 9 13 0 2
20 13 2 16 4 10 9 13 13 15 16 3 2 7 3 13 15 0 1 9 2
12 9 2 15 9 13 2 13 4 15 14 13 2
5 9 2 14 3 2
6 3 14 9 7 9 2
6 15 4 1 15 13 2
9 9 2 13 9 2 15 13 15 2
9 9 9 13 3 0 9 9 0 2
8 9 2 14 2 14 2 14 2
5 3 13 13 3 2
7 9 2 13 2 16 14 2
10 3 15 13 7 1 10 9 15 13 2
14 13 2 3 4 15 13 4 13 2 13 1 15 9 2
4 0 9 1 9
9 9 0 9 13 1 9 1 9 9
27 12 1 9 11 2 0 9 2 13 1 0 9 0 0 9 1 9 15 2 16 15 0 9 13 1 9 2
7 7 3 15 13 12 9 2
12 9 9 1 9 9 9 11 4 13 9 12 2
26 1 9 0 13 9 2 7 10 9 4 3 13 7 1 9 9 15 13 12 1 0 0 9 0 11 2
27 1 0 9 4 9 13 7 1 0 9 1 12 2 9 2 7 3 1 9 2 3 9 16 15 13 13 2
41 0 9 0 2 0 9 7 9 2 7 9 1 11 13 12 1 0 9 0 9 1 0 9 2 13 11 11 1 10 9 11 9 1 9 2 9 1 9 12 2 2
22 15 2 16 13 1 9 0 9 2 16 13 1 9 7 0 0 9 2 13 14 13 2
7 9 13 13 1 9 12 2
13 1 12 9 3 13 1 10 9 13 9 0 9 2
43 10 9 4 3 13 0 9 1 9 9 2 7 1 10 9 15 13 0 2 0 7 3 0 9 9 0 9 9 2 9 2 9 7 0 9 0 9 1 9 11 7 11 2
12 0 9 1 10 0 9 1 15 13 0 9 2
16 1 10 12 9 9 15 9 13 12 1 0 0 9 1 11 2
28 3 13 3 0 9 2 12 9 2 7 9 0 9 2 15 13 1 12 0 9 2 9 2 9 7 0 9 2
23 10 9 9 13 1 9 0 9 2 13 9 7 9 1 9 7 9 7 13 15 0 9 2
3 9 1 9
8 1 9 12 4 9 13 9 2
14 3 14 3 2 16 9 15 13 1 9 1 9 13 2
23 13 4 15 2 16 10 9 13 13 3 3 3 1 9 9 1 9 3 0 1 9 9 2
18 3 4 7 9 9 13 2 16 1 10 9 1 15 13 14 0 9 2
11 9 1 10 9 13 1 9 9 3 0 2
17 9 2 16 4 15 9 7 10 9 13 13 2 13 3 3 0 2
15 9 3 13 0 9 2 1 15 4 13 13 1 15 3 2
2 13 2
15 7 9 3 13 2 3 4 13 1 9 9 13 0 9 2
7 9 3 13 9 9 13 2
22 9 4 13 2 1 10 9 2 1 3 3 0 9 2 13 9 9 9 2 11 11 2
27 0 9 0 9 2 15 4 13 13 0 9 9 0 2 4 13 3 1 9 0 2 7 3 0 7 0 2
14 1 9 13 9 14 0 9 1 0 12 12 9 0 2
14 13 4 15 10 9 3 2 16 4 4 13 15 0 2
9 0 9 4 13 9 3 1 9 2
12 3 15 9 13 9 0 9 0 12 9 9 2
10 0 9 9 13 1 9 1 9 9 2
8 0 9 9 4 13 1 11 2
15 13 15 3 0 9 9 2 15 13 9 16 0 9 13 2
5 13 10 9 13 2
12 9 1 0 9 13 3 3 0 2 13 9 2
8 4 1 10 9 9 13 9 2
8 11 11 15 13 2 16 3 2
14 15 2 15 9 13 1 9 1 9 2 13 14 9 2
12 3 13 9 9 13 2 16 15 0 9 13 2
8 1 0 9 4 13 7 9 2
19 9 15 13 13 3 1 0 9 1 11 2 9 3 13 7 3 3 13 2
2 0 9
7 1 9 1 9 13 9 2
7 13 9 1 9 0 9 2
8 7 9 9 13 0 7 0 2
14 1 9 2 3 13 9 9 2 13 9 1 0 9 2
3 3 0 2
17 1 0 9 3 13 12 12 9 2 3 1 9 15 13 12 12 2
8 9 3 13 1 9 16 9 2
9 3 1 11 13 15 9 7 9 2
9 3 4 13 12 0 2 3 12 2
17 16 15 13 0 9 3 2 6 13 2 13 15 9 11 11 0 2
6 3 15 3 3 13 2
9 9 13 0 2 13 0 0 9 2
7 1 0 13 13 12 9 2
17 1 9 1 9 1 9 13 3 3 2 13 1 9 7 9 3 2
10 13 4 2 16 4 13 0 10 9 2
12 16 13 0 9 0 9 2 4 13 0 9 2
10 3 16 4 13 12 9 13 1 9 2
15 16 15 9 1 9 1 9 12 13 2 13 15 1 9 2
13 3 15 13 9 7 9 2 3 13 3 0 9 2
21 0 12 9 13 1 9 9 13 7 3 13 2 16 15 13 7 13 9 0 9 2
7 3 3 13 15 1 9 2
13 9 1 15 3 13 1 9 2 9 13 3 3 2
12 15 4 15 3 13 9 2 7 3 3 9 2
16 13 4 2 16 13 9 2 0 9 9 2 1 15 4 13 2
19 7 16 9 13 9 2 13 3 9 2 9 9 2 15 13 1 0 9 2
11 13 1 9 16 9 2 15 13 3 13 2
6 7 13 4 15 3 2
7 3 15 14 13 3 13 2
12 13 15 13 15 0 16 13 3 1 12 9 2
7 13 3 1 9 2 9 2
9 9 13 0 9 7 0 0 9 2
12 0 1 9 2 0 2 13 9 3 1 15 2
10 1 9 1 15 13 0 12 9 9 2
4 13 4 9 2
24 1 9 2 15 4 9 13 2 15 13 0 0 9 2 9 9 11 11 7 0 3 0 9 2
9 10 9 13 1 9 9 0 9 2
19 1 9 13 9 1 9 2 3 4 13 0 0 9 0 3 1 0 9 2
10 13 1 15 0 9 0 14 16 9 2
4 9 9 1 9
12 11 4 13 13 9 3 0 2 9 1 9 2
20 13 4 2 16 4 3 13 13 9 0 0 9 7 9 9 3 13 1 9 2
18 4 3 13 10 9 2 7 3 4 13 13 13 7 1 9 0 9 2
15 7 11 13 3 9 2 1 15 15 13 10 0 0 9 2
17 1 9 9 13 9 9 11 2 9 13 13 2 16 13 1 9 2
9 0 9 15 13 0 9 0 9 2
17 13 2 16 1 9 13 9 1 9 2 7 13 0 13 0 9 2
14 13 3 9 2 16 13 10 9 13 0 9 1 9 2
9 9 13 9 9 2 13 10 9 2
7 13 7 1 0 9 9 2
3 9 0 2
11 1 9 0 13 9 9 9 12 9 3 2
19 7 16 9 13 1 9 12 1 9 2 0 9 13 1 1 9 9 0 2
22 13 2 16 4 15 1 9 3 13 1 9 0 1 12 9 2 13 15 9 11 11 2
11 3 4 15 9 13 1 15 3 3 13 2
16 0 0 9 13 1 9 12 7 9 9 9 0 9 13 9 2
15 3 16 9 15 13 1 10 9 1 9 0 9 1 11 2
13 15 13 1 15 2 16 15 13 9 1 0 9 2
25 9 4 1 0 9 13 13 3 0 2 7 7 4 13 13 3 9 3 1 9 7 9 0 9 2
6 13 10 9 3 3 2
10 0 13 13 15 13 3 1 0 9 2
20 14 4 15 13 13 3 16 10 0 9 2 7 15 13 3 3 2 13 9 2
18 1 9 15 3 2 16 13 15 9 2 13 13 7 9 4 3 13 2
4 13 1 9 2
5 9 11 11 2 11
1 9
2 0 9
43 0 9 13 3 0 9 9 7 9 9 2 7 12 9 3 13 3 1 9 2 0 0 9 15 3 1 9 13 1 10 0 9 2 16 9 10 9 13 9 1 0 9 2
28 13 3 3 2 9 0 15 13 13 7 13 3 2 9 0 13 7 13 1 9 1 15 2 16 15 9 13 2
33 0 9 2 10 9 9 7 10 9 1 10 9 13 0 7 0 2 13 13 2 7 15 3 7 2 16 1 9 15 13 15 0 2
28 1 15 3 13 0 0 9 2 0 9 15 1 0 9 13 1 9 13 15 1 9 2 15 13 15 3 0 2
21 13 0 2 13 0 9 9 2 13 1 9 2 15 15 3 16 3 13 0 9 2
32 13 0 2 13 9 0 2 13 15 3 13 7 13 7 3 13 13 3 9 2 16 9 9 13 3 13 1 9 2 13 2 2
23 3 3 13 2 9 9 3 15 13 2 7 3 3 13 1 10 9 9 7 9 3 0 2
12 13 14 13 2 15 1 15 9 1 9 13 2
28 13 15 2 16 9 0 13 3 9 7 10 9 13 9 9 2 3 7 1 9 15 2 16 15 13 0 11 2
31 3 9 0 13 1 10 0 9 7 3 2 13 2 14 15 1 15 9 7 9 2 3 13 7 13 3 2 13 10 9 2
23 13 15 7 7 10 9 2 15 13 1 0 9 0 9 7 13 3 9 2 15 15 13 2
20 9 9 10 0 9 13 0 7 13 15 3 2 16 3 10 9 13 9 9 2
24 9 13 14 1 15 2 16 10 9 13 1 9 2 7 1 9 2 7 3 3 13 9 9 2
9 13 3 1 9 9 13 1 9 2
13 15 7 15 1 3 0 9 13 1 0 0 9 2
17 13 15 2 13 9 2 9 2 7 14 13 2 13 1 15 3 2
18 1 3 0 9 13 1 0 9 9 2 16 13 9 15 2 15 13 2
12 13 1 15 7 13 1 15 13 10 0 9 2
11 15 0 3 0 9 13 2 16 13 3 2
2 9 9
5 11 1 15 13 2
4 7 15 11 2
16 9 11 11 2 11 2 1 9 1 9 2 16 9 11 13 0
14 9 13 9 2 15 13 9 1 9 2 9 7 9 2
13 0 9 13 7 3 1 9 9 9 7 0 9 2
10 15 13 13 3 3 9 0 0 9 2
18 9 9 1 9 7 0 9 11 11 1 0 9 9 1 9 7 0 9
13 1 11 13 9 2 16 4 4 13 13 1 9 2
21 9 11 11 11 2 16 13 2 16 1 11 13 1 0 9 1 0 11 1 0 11
28 15 2 16 7 3 0 4 13 2 3 4 15 4 3 13 16 10 10 9 1 15 2 15 1 15 3 13 2
14 9 11 9 2 11 2 1 10 9 1 0 7 0 9
11 13 2 16 1 0 9 4 15 13 15 2
18 13 4 9 2 16 15 13 2 16 15 4 13 1 9 14 1 9 2
10 0 9 11 11 1 10 9 1 0 9
15 13 15 7 13 0 2 16 1 10 9 2 13 2 9 2
24 9 11 11 11 1 9 9 2 16 13 10 9 2 15 13 2 16 1 9 1 9 13 3 9
4 11 3 13 11
10 0 9 13 1 9 9 1 0 0 9
5 0 11 2 11 2
35 9 1 11 13 1 0 9 7 1 9 1 11 7 1 9 12 2 12 3 13 1 9 9 0 0 0 9 2 15 13 11 1 9 12 2
20 9 1 11 3 13 9 1 12 9 1 9 7 11 3 15 13 1 9 12 2
22 9 9 13 11 11 2 15 13 3 0 9 10 9 7 1 15 13 3 12 9 3 2
34 1 0 9 7 13 11 11 2 15 15 1 15 10 9 13 9 7 13 15 9 1 0 9 2 1 15 13 3 12 9 7 12 9 2
20 9 13 2 16 13 1 9 1 12 1 12 9 2 15 9 1 10 9 13 2
24 9 1 15 3 13 11 2 15 13 1 11 12 2 12 7 13 1 9 12 9 7 0 9 2
11 1 12 0 9 3 13 0 9 1 11 2
14 0 9 7 3 13 9 11 2 15 13 12 9 0 2
18 9 1 9 11 13 12 9 1 0 12 11 2 0 13 11 7 11 2
32 0 11 3 3 1 10 9 13 13 9 2 1 15 13 1 0 12 2 7 1 9 1 11 15 13 13 1 9 12 2 12 2
9 9 13 12 9 7 12 15 13 2
23 9 11 13 12 9 7 9 11 2 15 3 1 9 13 1 11 1 11 2 13 0 9 2
19 1 11 13 0 1 9 1 11 11 11 11 12 9 1 9 1 9 9 2
22 9 2 15 1 10 9 1 11 1 9 12 13 3 14 12 9 2 13 3 0 9 2
24 9 13 1 9 9 11 7 3 1 9 2 7 13 15 9 2 7 7 9 13 12 2 12 2
14 0 9 11 11 15 1 3 16 0 9 13 1 11 2
11 1 9 4 13 13 9 1 9 11 11 2
21 11 13 1 9 3 12 9 1 9 11 11 2 0 9 7 13 0 9 1 11 2
5 9 15 1 9 13
5 9 3 0 9 13
4 11 2 11 2
20 9 11 7 11 15 1 0 9 13 9 2 7 7 13 9 10 0 0 9 2
28 11 4 1 9 12 2 12 1 0 11 13 1 11 2 11 13 1 0 11 12 2 12 7 13 1 9 11 2
16 1 9 11 13 3 0 9 2 15 13 11 3 12 2 12 2
6 0 9 3 11 13 2
18 3 9 13 2 13 1 0 9 7 3 1 9 9 3 1 9 13 2
19 2 9 13 3 3 2 1 15 7 3 13 9 7 9 7 3 4 13 2
7 13 15 0 7 0 9 2
23 16 9 1 9 3 13 1 0 9 2 13 9 1 10 9 2 2 13 0 9 11 0 2
11 13 9 12 2 12 15 13 7 0 11 2
18 9 13 3 12 9 0 9 1 9 2 3 13 11 0 12 2 9 2
18 2 1 15 9 13 3 7 3 7 1 0 9 4 15 13 0 9 2
19 10 9 15 13 3 1 0 9 1 11 2 2 13 15 9 11 11 11 2
5 0 7 11 1 11
8 11 1 0 0 9 13 12 9
2 11 2
16 0 7 0 9 13 1 9 1 11 0 11 1 0 0 9 2
28 1 10 0 9 2 1 15 13 3 3 9 9 2 13 1 0 9 11 7 9 9 11 11 0 7 11 11 2
23 9 9 1 9 12 0 13 1 0 9 11 1 12 9 0 2 0 11 13 3 12 9 2
16 1 9 1 0 11 7 1 0 9 13 0 13 1 0 9 2
19 0 9 11 1 12 9 1 11 4 13 9 12 0 11 2 11 7 11 2
17 11 13 1 0 12 2 9 9 2 1 15 13 1 0 0 9 2
9 11 7 13 1 9 1 0 9 2
7 0 9 15 13 9 9 2
22 12 0 9 11 1 9 1 11 13 4 2 7 10 0 9 13 9 1 9 0 9 2
15 2 0 7 11 13 0 9 2 7 15 13 3 0 9 2
35 3 3 13 0 1 0 9 7 3 13 0 9 2 2 13 1 9 1 11 9 9 1 0 0 9 1 9 12 7 0 0 9 11 9 2
6 0 9 1 9 9 2
10 1 0 9 15 13 7 0 9 9 12
5 0 9 9 0 9
2 11 2
11 1 0 9 0 9 13 0 9 0 9 2
42 1 3 12 9 13 0 9 3 0 11 11 2 9 9 9 9 7 9 2 7 9 9 9 12 9 2 2 1 0 9 15 7 3 13 1 15 7 0 9 0 9 2
77 15 13 1 11 12 9 0 9 0 9 0 7 0 9 2 15 13 0 9 11 12 11 2 0 11 9 11 2 9 9 11 2 0 9 9 1 9 11 2 2 11 11 2 11 11 12 0 11 2 9 2 11 0 9 2 12 2 9 11 12 7 0 9 9 11 12 2 1 15 15 3 3 13 0 11 11 2
57 0 0 9 10 0 0 9 13 0 9 11 2 12 2 2 12 2 12 2 2 2 3 3 1 9 11 9 2 0 7 0 9 2 13 0 9 11 2 12 2 2 12 2 12 2 2 7 9 9 13 12 2 2 12 2 12 2
4 0 9 11 2
31 0 9 15 0 9 13 9 1 0 9 9 2 9 2 15 4 16 9 1 9 1 9 0 9 13 1 9 12 2 12 2
43 0 9 13 9 11 1 0 0 9 2 12 2 2 12 2 12 2 2 2 9 12 2 2 12 2 12 2 13 3 13 0 9 0 9 11 2 7 0 0 0 11 12 2
27 1 9 9 2 15 1 0 9 1 11 7 11 13 0 9 1 9 9 9 12 2 13 7 3 3 13 2
46 7 16 1 0 0 11 11 3 13 2 0 7 1 15 0 9 13 0 9 0 9 2 15 12 2 12 2 2 12 2 12 2 13 1 11 0 9 0 0 11 9 0 0 11 11 2
69 10 9 13 9 9 9 12 2 0 1 9 12 2 12 2 0 0 9 13 9 0 9 16 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 0 1 9 10 0 9 11 2 11 2 11 2 11 7 0 0 9 2
24 1 0 9 13 11 7 0 9 9 0 11 0 11 1 0 0 0 9 0 0 9 11 11 2
37 0 9 13 1 11 7 11 0 11 2 12 2 2 12 2 12 2 2 1 12 9 9 11 12 7 9 12 2 0 1 0 7 0 9 10 9 2
65 1 0 0 9 1 0 9 13 1 0 11 11 2 12 2 2 12 2 12 2 2 1 9 9 11 2 12 2 2 12 2 12 2 2 7 12 9 9 0 0 2 0 9 11 9 12 2 12 9 2 9 7 9 2 0 3 9 0 11 11 7 11 12 11 2
51 3 15 13 12 2 2 12 2 12 2 2 12 2 2 12 2 12 2 2 12 2 2 12 2 12 2 7 12 2 2 12 2 12 2 2 1 9 0 9 13 9 3 12 9 0 0 9 1 2 9 2
3 11 1 11
2 11 2
17 1 10 0 9 11 13 3 0 9 12 2 9 1 11 1 11 2
15 13 1 15 9 9 0 0 9 11 11 1 9 11 11 2
9 9 13 0 3 0 9 1 9 2
9 10 9 13 9 9 11 0 11 2
5 9 13 13 1 11
2 11 2
22 0 0 9 13 0 9 1 9 1 9 1 11 2 12 2 12 2 2 1 9 11 2
26 1 0 9 15 1 15 3 13 9 0 9 11 11 11 2 9 11 11 11 7 10 0 9 11 11 2
21 0 13 3 0 9 1 9 2 9 4 13 9 1 9 3 1 9 12 2 9 2
27 11 11 1 9 9 1 9 12 13 1 0 9 11 2 15 4 15 13 13 1 0 9 1 9 9 7 9
4 0 9 13 9
8 0 9 1 0 9 7 11 11
4 11 1 11 2
31 0 9 1 10 0 9 3 9 9 13 1 0 1 0 9 7 10 9 13 1 0 9 9 0 9 1 0 7 0 9 2
25 11 11 13 3 3 9 1 9 9 1 9 2 11 11 13 9 0 9 0 9 1 9 1 11 2
21 9 2 15 13 1 12 9 9 11 2 3 13 9 9 1 9 11 1 0 9 2
22 1 0 9 0 9 13 1 0 9 0 9 9 11 2 15 13 7 0 0 0 9 2
33 9 4 13 11 11 2 11 11 2 11 11 2 0 9 3 11 9 2 11 11 7 0 9 11 11 2 15 13 1 9 9 11 2
29 1 9 3 13 9 11 11 2 11 11 7 3 0 0 9 11 11 2 15 1 9 12 13 9 11 9 1 9 2
10 9 9 13 0 9 1 0 0 9 2
49 11 11 4 1 0 9 13 3 13 9 9 9 1 9 2 0 9 11 11 13 9 1 9 11 1 9 2 15 15 13 1 9 2 7 0 9 4 13 3 13 1 9 0 9 7 1 0 9 2
3 1 0 9
22 11 11 2 12 2 2 9 11 11 2 13 3 0 11 2 15 13 9 1 0 9 2
17 0 9 1 15 13 9 11 7 14 13 13 13 11 12 9 9 2
26 3 9 15 4 13 11 11 13 1 11 11 11 2 12 2 2 9 13 1 9 0 9 1 0 9 2
7 11 1 0 0 9 1 11
2 11 2
14 9 0 9 11 1 11 1 0 9 3 13 3 13 2
20 1 9 9 0 9 0 0 9 11 11 13 3 0 9 9 9 13 0 9 2
11 2 13 4 1 15 1 0 9 3 3 2
15 1 9 15 3 7 13 9 2 9 15 0 9 13 3 2
13 3 15 13 1 9 9 0 15 2 1 9 2 2
13 9 4 15 13 13 7 14 13 2 2 13 11 2
2 9 9
3 0 11 2
15 12 9 7 12 9 4 13 1 11 1 9 1 0 9 2
22 13 15 1 3 0 9 0 1 10 9 2 15 13 3 1 9 9 0 9 11 11 2
21 3 15 9 13 14 0 9 2 9 13 1 9 9 11 11 1 9 1 9 9 2
4 11 3 1 9
4 11 1 11 2
28 1 11 1 11 3 13 0 9 0 0 9 1 9 11 11 2 15 15 13 3 0 9 11 11 7 11 11 2
12 9 15 3 13 1 0 9 1 9 1 9 2
25 9 13 13 0 9 9 1 0 9 2 15 15 13 2 7 3 9 9 1 7 1 9 1 9 2
12 3 13 1 0 9 9 1 9 0 9 9 2
54 1 0 9 3 13 1 12 9 2 9 12 2 9 12 2 9 11 2 11 15 4 13 12 2 9 1 12 2 12 9 1 1 9 9 1 0 9 7 9 12 2 9 12 2 9 0 11 2 11 3 12 2 9 2
5 11 1 9 1 11
5 0 13 0 0 9
2 11 2
34 2 13 9 0 2 2 13 0 0 9 11 11 3 2 16 1 9 0 0 11 13 0 0 9 11 11 12 2 12 2 12 2 12 2
24 0 11 0 1 11 13 1 11 9 1 0 0 7 0 9 11 2 12 2 9 9 11 2 2
23 1 0 9 11 2 12 2 2 15 7 13 2 7 16 15 1 0 9 0 9 13 9 2
10 2 13 4 2 16 4 13 3 3 2
13 13 15 2 3 10 0 9 7 0 9 1 9 2
20 13 3 13 9 7 13 9 2 3 3 13 7 0 9 2 2 13 9 11 2
22 1 10 9 13 2 16 15 1 0 9 13 0 9 2 7 3 16 3 15 15 13 2
39 2 13 15 1 11 1 9 7 1 15 13 1 9 2 15 13 9 2 2 13 11 2 12 2 2 2 15 15 1 9 1 9 1 0 9 3 13 13 2
11 2 15 15 13 2 13 3 3 7 3 2
28 1 0 9 7 15 0 13 0 9 2 2 13 11 2 15 4 1 9 9 7 9 13 1 0 9 0 11 2
3 11 13 9
3 0 11 2
21 1 15 2 15 13 9 11 11 11 1 9 0 9 9 11 2 3 3 13 13 2
17 1 0 9 0 9 13 9 9 11 11 11 1 11 11 1 11 2
17 1 9 0 9 7 11 13 7 13 3 10 9 1 12 2 12 2
14 1 9 1 9 15 3 13 3 14 9 9 1 9 2
5 11 7 11 13 9
2 11 2
27 11 7 11 3 1 11 13 9 1 9 7 3 3 13 12 9 0 0 9 2 15 15 13 10 9 9 2
11 13 15 9 0 9 9 11 1 11 11 2
34 9 2 15 13 9 9 9 11 7 11 11 11 1 11 7 11 11 2 13 9 2 15 9 9 3 13 11 7 15 11 1 9 13 2
13 11 7 1 9 1 9 13 11 2 16 9 13 2
19 1 0 0 9 0 9 3 13 1 0 9 0 1 0 9 1 12 9 2
9 11 4 13 1 9 0 9 1 9
2 11 2
34 11 1 9 9 0 9 1 9 2 11 2 1 9 0 2 0 7 0 9 13 7 1 9 2 16 13 9 3 0 9 2 11 2 2
19 13 15 3 1 11 0 9 9 11 11 1 0 0 9 0 9 1 11 2
30 11 13 1 9 11 0 9 2 7 7 13 9 10 9 13 9 0 9 2 15 3 13 0 9 7 13 15 0 9 2
20 11 13 2 16 0 2 0 9 1 9 0 9 12 0 9 13 1 9 9 2
30 1 11 13 0 2 16 4 11 1 9 2 3 13 9 9 0 7 0 11 1 0 0 9 2 13 9 0 9 9 2
33 9 11 14 1 9 1 0 12 9 0 0 9 9 2 14 12 9 9 2 13 1 9 2 15 13 11 13 15 0 9 1 9 2
10 1 12 0 9 13 9 11 14 12 2
13 11 3 13 1 9 0 9 16 1 9 0 9 2
31 1 0 0 9 2 15 13 13 1 0 14 9 0 9 2 13 9 9 1 9 11 1 0 9 11 7 9 0 0 9 2
28 11 13 2 16 16 11 2 15 13 0 1 2 13 1 9 11 2 13 7 9 1 0 9 1 10 0 9 2
16 0 9 15 13 0 9 2 7 3 13 1 9 2 13 11 2
19 3 11 13 9 0 9 3 2 16 4 13 10 9 2 3 0 9 11 2
26 0 9 7 9 1 9 9 11 11 13 10 9 1 9 9 1 9 1 0 9 11 2 1 2 11 2
19 9 7 13 1 3 9 9 2 15 9 7 9 13 3 9 1 9 9 2
5 9 9 13 1 9
2 11 2
21 9 0 0 9 11 11 15 4 13 1 9 1 9 1 9 10 9 13 1 9 2
8 13 1 15 0 9 1 11 2
16 1 0 9 13 9 1 11 7 0 9 9 11 11 1 9 2
18 9 3 12 2 9 13 9 9 2 1 15 13 1 9 1 0 9 2
19 12 0 15 3 16 9 9 3 13 1 0 9 9 9 0 9 1 11 2
4 11 13 0 9
2 11 2
35 1 2 3 0 7 3 0 2 13 1 9 1 9 1 11 9 0 9 9 11 11 9 9 0 9 0 0 9 2 15 4 13 1 11 2
18 1 9 13 1 0 9 9 7 9 0 9 13 1 0 9 0 11 2
15 9 0 9 1 11 13 0 9 0 9 0 9 11 11 2
31 10 9 1 0 13 2 16 4 13 4 13 9 1 0 9 15 2 15 4 1 11 13 9 2 15 4 1 9 13 11 2
22 13 4 3 9 1 0 9 10 9 2 15 13 1 11 0 9 7 13 15 1 11 2
5 9 11 11 4 13
2 11 2
16 0 9 13 1 9 1 0 9 11 0 9 9 11 11 11 2
28 13 15 1 0 9 0 9 11 2 11 1 9 1 9 1 9 0 9 0 9 11 11 2 15 13 0 9 2
7 0 9 10 9 3 13 2
11 0 11 11 13 16 9 0 9 1 11 2
22 3 2 16 15 10 9 11 13 1 10 0 9 9 2 15 13 10 9 7 0 9 2
18 4 13 1 2 0 9 2 1 0 9 7 13 15 0 9 1 9 2
23 0 9 3 13 1 9 0 9 1 11 2 15 4 13 13 0 9 1 0 9 12 9 2
17 13 15 3 9 9 0 9 11 11 2 15 15 13 9 1 11 2
6 2 9 13 10 9 2
30 13 15 9 2 15 15 13 7 14 15 15 13 13 2 2 13 11 2 15 13 1 9 0 9 1 11 9 11 11 2
29 0 7 0 9 15 3 13 1 9 0 12 0 9 2 15 13 13 3 1 9 0 9 2 1 9 12 0 9 2
27 13 15 0 0 0 9 11 11 2 15 15 13 0 0 9 0 2 0 9 1 0 11 2 0 0 9 2
22 0 9 12 9 15 13 1 9 0 9 7 0 2 15 15 13 13 1 11 3 3 2
3 11 13 9
8 0 0 9 13 0 9 9 9
13 9 9 11 15 3 3 1 11 13 1 0 9 2
18 3 0 9 0 9 1 9 0 0 9 11 13 0 9 1 9 9 2
16 9 0 9 1 9 13 1 12 9 9 1 0 9 11 11 2
10 1 0 9 15 13 3 1 0 9 2
28 2 0 9 1 0 9 2 2 3 15 0 0 9 1 9 13 2 15 13 0 7 3 3 14 0 0 9 2
9 9 0 9 13 1 10 9 9 2
28 4 2 14 11 13 2 13 15 3 10 9 2 9 9 7 3 1 15 7 1 0 9 3 0 9 11 11 2
14 15 3 1 0 9 9 13 15 0 2 16 13 9 2
38 1 9 0 9 13 0 0 9 11 11 9 0 0 9 11 2 15 1 9 12 3 13 12 9 0 1 9 1 0 9 11 2 11 7 10 9 2 2
26 3 1 9 9 13 11 1 0 2 13 12 9 11 0 13 2 0 9 11 11 7 0 9 11 11 2
23 16 12 3 13 2 9 11 14 13 1 0 9 0 9 7 3 4 13 1 9 9 9 2
27 1 9 9 13 1 9 12 2 12 9 0 9 9 3 0 11 12 9 9 7 1 9 12 0 12 9 2
38 16 9 1 15 9 0 9 3 13 7 0 11 1 10 9 1 9 10 9 9 11 13 1 0 9 1 9 7 13 10 9 2 9 13 1 0 9 2
12 9 0 9 9 0 9 13 1 9 0 9 2
29 16 7 0 0 9 0 9 9 13 2 16 13 0 0 9 9 13 3 2 16 15 13 3 2 13 11 0 9 2
22 11 15 1 9 3 3 13 7 1 12 9 9 4 15 11 13 1 0 9 3 13 2
28 3 1 0 0 9 1 9 12 13 9 10 0 9 1 9 7 3 13 14 1 9 1 0 9 9 7 9 2
23 0 9 1 0 0 9 11 11 11 1 9 4 3 1 9 13 0 9 1 9 1 9 2
13 1 15 3 7 1 0 9 7 9 0 9 13 2
9 9 11 15 1 15 13 0 9 2
20 16 0 9 0 9 13 9 9 9 2 15 0 4 3 13 14 1 9 12 2
10 11 7 3 13 2 16 4 9 13 2
9 10 9 4 13 14 3 3 13 2
22 1 0 0 9 0 9 7 0 9 9 13 3 1 9 9 11 15 7 9 13 9 2
4 0 9 13 9
2 11 2
20 9 11 11 1 0 9 13 9 2 9 9 2 1 12 9 9 0 0 9 2
16 0 9 13 2 16 15 15 1 9 9 13 9 1 9 13 2
13 13 13 2 16 1 9 13 1 9 9 10 9 2
6 3 9 13 9 9 2
11 1 10 9 13 13 2 16 13 0 9 2
7 9 13 0 9 0 9 2
3 11 1 9
1 11
16 12 1 12 9 0 0 9 15 3 3 13 1 9 9 11 2
25 9 9 9 11 11 1 9 1 9 9 13 2 16 1 11 7 1 9 11 4 3 13 9 0 2
40 9 0 0 9 11 11 3 13 2 16 9 0 9 11 1 11 13 0 7 16 4 15 11 2 1 1 10 9 1 9 9 2 9 2 13 13 1 9 9 2
26 2 1 11 4 13 13 10 9 2 13 2 15 15 1 15 13 2 1 15 13 0 2 2 13 11 2
2 11 9
2 11 2
29 9 1 9 11 7 0 9 1 9 0 9 11 11 1 9 0 2 0 9 13 0 2 13 3 0 9 11 11 2
8 2 9 1 9 4 13 0 2
14 9 13 2 13 15 3 9 9 2 2 13 0 9 2
14 13 2 16 13 13 15 2 3 3 9 0 9 13 2
2 9 9
1 9
16 1 0 9 2 3 0 9 2 15 3 10 9 13 0 9 2
20 3 0 9 2 0 9 7 0 9 13 11 2 11 2 0 1 0 9 13 2
7 3 13 10 9 0 9 2
5 9 13 0 9 2
7 13 15 3 1 9 12 2
14 9 0 9 3 13 13 0 9 0 15 0 2 9 2
25 3 15 3 13 2 16 0 9 15 13 3 13 1 9 9 7 9 1 9 15 13 13 14 3 2
10 9 9 0 15 3 13 9 9 11 2
22 16 1 0 9 13 0 2 0 9 2 3 15 13 1 9 12 2 1 9 9 11 2
23 3 0 11 4 2 3 3 2 13 9 2 9 2 9 2 10 1 15 13 0 9 13 2
10 9 11 15 3 13 1 9 9 9 2
7 9 2 1 10 9 13 2
13 9 3 13 0 7 3 0 9 15 11 1 9 2
18 1 9 2 3 9 9 13 3 3 2 15 13 1 9 11 9 0 2
27 3 15 13 2 16 10 9 13 3 1 9 1 0 0 9 0 9 9 11 2 15 3 13 1 0 9 2
10 0 9 1 9 13 1 0 9 11 2
12 7 7 13 3 0 9 9 1 0 0 9 2
22 9 7 9 0 15 1 0 9 13 0 10 9 13 1 9 2 15 4 13 10 9 2
20 10 9 15 1 15 9 13 7 10 9 1 15 0 9 11 2 11 2 13 2
5 9 13 9 9 2
7 11 3 14 13 1 9 2
21 13 3 1 0 9 2 15 1 0 9 2 1 9 12 2 13 3 13 1 9 2
28 2 13 4 9 0 9 2 15 15 13 2 7 7 15 13 2 2 0 9 0 9 15 13 0 14 3 13 2
17 1 9 13 3 0 9 2 15 0 9 1 11 13 1 15 9 2
4 9 3 13 2
15 0 0 0 9 0 9 1 11 15 14 13 9 11 13 2
11 9 13 2 16 9 0 9 13 3 0 2
4 9 1 0 9
1 9
16 9 1 0 11 3 13 9 0 0 9 7 3 15 9 13 2
20 3 2 16 1 3 0 9 15 0 13 13 9 1 9 0 9 2 9 13 2
11 9 13 9 2 3 13 1 9 0 9 2
12 16 9 13 13 0 2 0 9 13 13 0 2
13 1 0 11 4 12 2 9 13 0 9 11 11 2
11 13 15 0 0 9 2 10 9 15 13 2
6 3 1 0 9 13 2
23 13 0 9 7 13 15 1 9 15 1 15 3 3 13 14 1 0 9 7 3 1 9 2
12 13 15 7 13 2 9 13 14 1 0 9 2
36 16 7 9 2 9 2 9 7 0 9 13 2 1 9 9 0 9 7 1 1 9 9 2 9 0 9 3 13 2 1 9 0 9 15 13 2
27 9 1 9 1 9 7 9 7 0 9 13 3 0 2 16 7 9 0 1 9 1 9 9 1 9 13 2
28 9 1 9 1 11 3 13 2 16 9 9 0 9 13 1 0 9 2 16 1 9 9 15 13 1 0 9 2
16 13 0 13 9 2 15 13 10 9 1 9 7 13 10 9 2
11 7 9 4 3 13 3 3 16 0 9 2
15 13 0 2 16 7 9 9 4 1 9 3 13 13 3 2
6 0 11 13 15 9 2
10 7 7 1 11 15 1 15 13 0 2
4 0 9 7 9
24 3 4 13 1 0 9 2 15 13 0 1 3 0 9 13 9 1 9 10 9 7 12 9 2
11 13 10 9 13 16 9 1 0 0 9 2
13 1 3 0 9 13 0 9 0 9 1 0 9 2
26 0 13 9 2 16 3 3 15 13 13 1 0 9 1 0 9 9 7 15 16 13 1 0 9 0 2
19 2 3 0 13 10 9 1 0 9 2 15 0 9 13 1 0 9 2 2
22 10 9 15 13 3 0 1 0 1 9 0 11 2 3 3 9 0 9 13 0 9 2
22 12 1 0 9 9 2 3 2 0 2 9 11 2 3 1 9 0 9 13 10 9 2
6 9 13 7 3 0 2
4 9 13 10 2
22 3 2 16 15 13 1 10 3 15 0 9 2 13 15 13 3 0 2 16 13 0 2
21 9 13 0 9 2 15 13 3 10 9 2 16 9 13 2 7 3 13 1 9 2
17 1 15 15 13 14 3 3 7 3 13 13 9 2 16 13 3 2
27 3 7 16 13 1 9 3 0 9 2 1 10 9 13 13 9 2 3 2 13 0 2 16 13 10 9 2
21 13 15 9 0 3 0 9 9 9 2 15 12 9 13 3 1 0 9 1 9 2
11 2 3 13 2 3 13 10 0 0 9 2
18 13 1 12 3 0 9 2 1 15 4 3 13 0 9 0 0 9 2
5 13 13 3 2 2
21 1 10 9 15 13 2 16 10 0 0 9 13 9 9 3 0 9 1 0 9 2
16 9 0 3 0 9 13 3 0 9 1 0 9 1 10 9 2
12 0 0 9 13 9 2 16 9 13 1 9 2
7 13 7 0 9 9 9 2
23 3 1 9 12 13 11 11 11 13 0 9 1 0 9 1 0 9 1 0 9 1 11 2
16 11 13 3 9 1 0 9 1 12 12 9 3 16 0 9 2
14 9 2 15 15 13 2 13 3 9 0 9 7 9 2
24 13 15 1 0 9 2 1 0 9 1 0 9 2 1 0 9 2 15 1 15 7 13 13 2
28 9 9 12 0 9 1 9 13 9 0 9 0 9 9 11 11 11 1 10 0 9 11 11 1 0 9 11 2
13 9 13 2 16 12 9 13 9 7 13 10 9 2
33 16 9 13 1 0 9 2 13 0 9 11 11 2 2 14 2 2 2 2 2 7 0 2 0 7 0 9 15 13 3 1 9 2
10 15 9 13 3 2 15 13 0 9 2
15 1 9 0 9 7 9 13 3 3 0 13 1 9 9 2
17 1 9 15 13 7 0 9 2 7 9 9 2 15 13 1 9 2
8 9 13 0 7 13 15 3 2
14 13 0 3 0 7 0 15 13 13 2 3 3 13 2
9 13 3 13 13 9 2 7 9 2
30 9 3 13 9 7 9 9 2 15 13 3 1 0 9 2 2 7 10 0 9 2 9 7 9 2 15 13 3 2 2
18 13 15 3 2 16 9 1 9 13 9 9 2 7 10 9 7 9 2
10 3 7 3 0 9 13 13 0 9 2
10 13 3 9 2 3 0 16 0 9 2
25 0 11 3 1 9 0 9 13 2 16 15 1 0 9 3 3 13 9 0 9 12 0 0 9 2
9 10 9 13 1 9 0 0 9 2
17 10 9 1 9 0 9 13 9 2 15 13 9 9 1 0 9 2
18 11 15 1 10 9 13 1 0 7 0 9 2 13 14 3 13 9 2
8 9 11 3 1 9 1 9 13
5 14 2 0 9 2
2 11 2
23 9 13 13 13 1 12 2 9 1 11 9 1 9 10 9 1 0 9 9 1 0 9 2
10 1 0 9 9 11 15 13 11 11 2
18 0 9 9 9 13 3 13 2 13 7 0 2 16 10 13 0 9 2
13 9 9 7 0 9 11 11 15 3 9 9 13 2
16 10 0 9 13 1 9 2 0 1 9 9 9 2 13 0 2
32 1 9 2 15 3 11 13 9 2 13 0 13 3 13 0 9 2 1 15 13 0 13 9 0 9 2 9 9 7 0 9 2
10 7 9 15 13 9 15 1 9 13 2
19 16 4 13 9 3 0 9 13 9 1 9 2 15 15 1 15 4 13 2
30 11 7 13 2 16 3 9 13 0 9 3 1 2 16 10 0 9 2 0 1 0 9 2 15 13 14 1 9 12 2
21 9 1 0 9 9 9 1 0 9 15 1 10 9 1 9 9 7 0 9 13 2
16 1 9 11 11 11 13 9 13 1 9 2 7 1 9 9 2
18 11 13 2 16 4 13 0 7 0 9 2 1 0 9 1 9 9 2
22 9 9 1 0 11 1 0 9 13 9 9 1 9 2 16 9 9 1 9 9 13 2
5 9 13 13 9 9
3 1 0 9
9 0 0 2 9 11 2 11 2 2
31 1 9 9 0 9 11 13 11 9 9 2 16 13 1 2 0 9 2 9 1 15 2 16 4 13 13 1 9 9 11 2
15 13 7 2 16 13 9 13 9 0 15 9 9 0 9 2
15 1 10 9 4 1 9 1 9 13 13 9 0 1 9 2
17 9 9 11 11 15 3 1 9 0 9 9 0 9 13 9 13 2
10 2 13 0 13 1 10 0 0 9 2
9 1 15 13 13 7 13 15 0 2
26 3 13 13 9 3 0 9 9 0 9 2 13 9 1 9 2 9 2 9 9 9 2 2 13 11 2
8 9 11 3 1 9 1 9 13
5 11 2 11 2 2
23 9 13 13 13 1 12 2 9 1 11 9 1 9 10 9 1 0 9 9 1 0 9 2
19 11 11 13 2 16 4 13 0 7 0 9 2 1 0 9 1 9 9 2
4 9 13 13 0
5 14 2 0 9 2
2 11 2
16 9 15 3 13 1 10 0 9 2 7 15 1 0 9 13 2
15 1 9 1 9 10 0 9 15 3 13 9 11 11 11 2
17 13 2 16 9 13 13 9 0 9 2 7 3 2 3 0 9 2
13 1 9 12 13 9 9 9 2 15 13 10 9 2
12 3 3 13 1 11 9 1 11 7 0 9 2
29 1 1 15 2 16 9 0 9 15 1 0 9 13 1 9 1 9 2 13 14 0 2 16 15 13 9 1 15 2
27 11 13 2 16 9 13 9 13 1 9 0 9 1 9 9 12 9 2 15 4 3 2 13 0 9 2 2
12 9 13 1 15 9 2 3 7 1 0 9 2
17 15 15 13 9 1 9 2 7 1 9 2 16 15 13 9 11 2
16 10 9 11 13 2 7 15 13 1 0 9 0 9 0 9 2
10 7 1 9 9 11 4 13 0 9 2
8 11 13 13 0 9 1 0 9
6 11 11 1 9 1 11
10 1 11 15 1 9 13 9 0 9 2
20 9 2 15 1 9 0 9 13 9 1 9 12 7 3 13 1 12 9 9 2
18 10 9 11 11 15 7 3 13 12 1 0 9 1 9 9 0 9 2
11 0 9 3 0 9 13 15 1 9 13 2
12 4 1 9 13 1 0 9 1 0 0 9 2
14 0 9 13 1 15 2 15 4 15 13 1 9 11 2
37 13 1 15 3 3 3 2 1 9 4 13 12 9 2 0 9 3 12 2 7 16 15 4 13 10 9 2 13 4 15 1 9 13 1 12 9 2
12 13 4 15 9 9 1 9 0 9 11 11 2
8 1 0 9 4 15 7 13 2
2 3 2
11 13 4 15 7 2 16 4 15 13 13 2
19 3 16 4 13 3 1 9 1 11 11 2 3 4 15 13 1 11 11 2
23 13 4 1 9 1 0 7 0 9 10 9 7 1 15 2 3 13 9 0 9 1 15 2
8 10 9 0 0 9 13 15 2
30 13 13 2 16 16 4 15 13 1 9 3 12 9 2 3 1 15 13 0 9 0 9 2 3 13 13 12 0 9 2
13 15 3 13 1 15 2 3 15 4 0 9 13 2
18 3 10 9 13 1 11 2 7 13 3 2 16 13 2 9 3 12 2
22 9 13 3 2 15 15 3 13 1 0 9 2 16 4 13 3 3 9 13 0 9 2
15 13 7 2 15 15 4 13 1 11 2 15 13 10 9 2
17 10 10 9 2 16 9 11 2 15 13 7 13 15 13 9 0 2
9 16 15 15 15 13 2 13 9 2
11 16 0 9 13 0 9 1 9 0 9 2
9 16 4 13 1 9 2 13 4 2
2 3 2
10 7 15 10 9 13 3 3 3 0 2
22 7 15 13 2 16 11 13 9 13 1 9 2 0 1 9 7 1 9 0 0 9 2
20 13 15 9 9 2 15 13 0 1 9 13 1 10 9 2 15 13 9 3 2
31 3 13 15 9 9 2 7 15 13 0 2 9 13 13 2 3 13 1 9 10 9 2 1 10 9 1 11 7 1 9 2
37 9 0 9 4 15 13 3 13 16 9 2 7 16 9 2 15 13 3 3 0 9 7 15 15 13 1 10 9 13 9 2 3 3 13 0 9 2
6 1 0 9 13 9 9
2 11 2
41 1 9 9 11 11 11 13 9 9 0 9 0 2 0 7 0 9 1 11 9 1 9 0 1 0 9 7 3 13 9 1 9 9 2 16 15 4 13 10 9 2
30 9 9 9 13 3 1 15 9 9 7 10 9 1 9 2 16 15 13 0 2 16 13 1 9 2 3 3 0 2 2
39 11 2 11 13 2 16 4 0 0 9 2 15 13 1 11 0 1 9 0 9 2 13 9 10 9 2 16 2 13 3 13 2 16 15 1 9 13 2 2
36 1 9 0 0 9 11 11 11 13 9 9 2 0 9 2 15 13 13 9 2 2 7 0 9 1 9 4 13 9 1 10 9 1 0 9 2
53 9 2 16 9 2 13 1 0 9 9 9 2 15 13 1 9 9 3 0 7 13 2 9 7 0 9 2 2 16 4 15 13 2 10 9 9 7 9 1 9 0 0 2 0 2 0 2 0 7 0 9 2 2
35 9 0 0 9 11 11 1 0 0 9 13 2 16 2 16 15 15 13 2 16 9 13 13 7 1 11 2 3 13 2 1 15 13 2 2
6 11 13 15 9 13 2
9 11 11 7 11 11 1 0 9 11
7 11 13 1 0 9 1 9
3 1 0 9
2 11 2
24 11 13 9 0 0 9 2 13 7 2 16 9 1 9 1 0 9 2 3 4 13 2 13 2
8 13 15 3 9 9 11 11 2
17 0 0 9 11 3 13 0 9 1 9 2 0 15 0 0 9 2
18 1 11 4 11 13 9 9 1 9 0 9 2 3 0 1 0 9 2
10 10 9 4 7 13 4 13 0 9 2
16 1 9 4 14 13 0 9 9 13 1 9 3 2 0 9 2
20 1 0 9 4 13 9 13 3 10 9 2 10 0 9 13 12 9 0 9 2
5 9 13 13 9 9
1 3
32 0 9 11 13 9 9 7 0 0 9 0 9 0 11 11 1 9 7 13 9 2 16 15 11 13 0 0 9 0 15 9 2
13 15 1 10 9 13 1 11 9 0 9 1 9 2
3 9 3 13
1 3
17 9 9 1 11 2 15 13 0 9 1 11 2 15 13 1 11 2
11 13 15 15 13 1 12 9 0 0 9 2
11 9 0 9 15 1 0 11 3 16 13 2
12 12 0 9 4 13 12 9 1 0 12 9 2
20 0 9 1 11 7 10 0 9 13 1 9 9 11 11 13 9 0 0 9 2
4 11 9 9 13
11 11 2 1 0 9 9 1 9 13 0 9
2 11 2
24 9 11 3 13 9 9 0 9 1 9 0 0 9 2 15 1 9 13 9 0 9 1 0 2
21 1 9 9 11 11 13 1 0 9 0 9 1 15 2 16 4 4 9 3 13 2
24 0 0 9 1 11 13 9 2 16 3 13 10 0 9 2 15 15 9 13 1 9 10 9 2
23 9 13 14 3 0 2 9 13 2 16 13 15 1 9 2 7 13 3 1 9 3 13 2
19 13 14 1 9 0 9 9 2 3 13 1 9 7 3 15 3 13 2 2
15 11 3 13 2 16 13 1 0 9 11 3 13 10 9 2
15 0 9 1 9 9 13 1 15 0 16 0 9 9 11 2
31 2 13 2 14 15 7 2 16 0 9 13 3 9 1 0 9 9 16 9 1 10 9 2 0 1 9 13 2 2 13 2
25 1 10 9 4 9 13 10 9 9 2 13 3 0 0 9 2 16 13 0 9 3 1 9 2 2
39 1 9 11 2 16 4 13 11 0 13 2 16 15 1 10 9 13 2 11 13 2 2 11 15 13 7 0 9 13 0 7 9 9 0 9 9 13 2 2
17 13 2 16 11 13 7 3 13 13 1 0 9 1 9 0 9 2
29 9 0 9 11 7 9 0 9 11 11 13 2 16 12 9 9 4 13 3 7 1 15 13 9 3 1 15 9 2
23 13 2 16 15 9 1 9 4 13 7 3 7 4 13 1 9 15 9 2 15 11 13 2
37 9 9 2 15 4 15 13 13 9 9 9 2 4 1 11 13 13 0 2 2 13 2 14 15 3 2 13 7 3 13 15 2 15 13 13 2 2
8 0 9 13 9 7 1 0 9
2 11 2
15 0 9 1 9 4 14 3 0 13 10 9 3 0 9 2
18 1 12 1 15 2 11 11 1 0 0 9 2 7 9 3 9 13 2
6 2 10 9 13 0 2
9 3 9 1 9 13 1 9 0 2
21 13 15 7 9 13 3 0 9 2 16 1 15 13 0 2 2 13 11 2 11 2
22 1 0 9 15 10 9 13 2 16 1 0 9 16 4 3 15 13 1 9 0 9 2
25 13 15 3 0 7 3 3 0 9 2 3 0 9 7 9 2 3 13 9 7 3 9 7 9 2
8 9 3 13 3 9 3 0 2
14 3 15 13 3 1 0 9 1 11 7 1 0 9 2
15 1 0 0 9 13 9 1 10 9 9 2 9 7 9 2
18 0 9 11 13 2 16 9 1 10 9 13 0 3 1 10 0 9 2
11 9 13 1 9 0 0 9 7 7 9 2
15 3 15 2 15 15 13 3 13 2 3 13 9 1 9 2
18 1 9 12 13 9 9 1 9 7 9 13 2 3 13 9 3 13 2
12 9 9 7 13 14 0 9 2 7 3 9 2
13 1 9 12 9 13 9 3 12 7 12 9 3 2
10 7 3 13 9 3 14 9 7 9 2
19 0 9 1 0 9 11 11 13 2 16 15 13 13 3 9 7 0 9 2
10 3 16 9 13 9 9 9 7 9 2
20 11 11 3 13 2 16 3 9 1 9 7 9 13 13 9 0 9 7 9 2
11 13 1 9 2 16 0 9 0 9 13 2
14 1 15 3 13 0 9 0 9 7 13 9 1 9 2
12 10 9 14 13 3 9 0 1 9 1 9 2
6 0 9 11 11 2 11
2 11 2
23 0 9 0 9 13 3 0 9 9 0 11 11 2 9 9 2 9 7 9 1 0 9 2
18 9 11 15 13 1 9 12 1 0 11 7 13 1 0 9 1 11 2
26 1 9 13 1 9 1 11 7 1 9 12 4 13 1 0 9 2 3 13 13 16 9 0 0 9 2
9 1 10 9 3 13 1 0 9 2
24 1 0 9 11 11 11 15 9 11 3 13 1 9 0 0 0 9 1 11 7 1 11 11 2
6 9 14 13 1 9 13
2 11 2
25 0 9 0 0 9 0 0 9 1 0 9 1 11 13 9 1 9 1 9 7 9 0 9 9 2
7 13 15 10 9 11 11 2
22 9 4 1 15 13 13 9 0 9 1 9 2 16 3 1 15 9 13 4 7 14 2
22 11 13 2 16 9 3 1 9 13 1 0 9 2 7 9 12 9 15 3 13 9 2
10 9 4 13 3 1 9 9 1 9 2
11 9 9 11 11 4 13 1 9 13 3 2
7 1 9 13 0 9 9 2
17 1 9 9 0 9 11 11 4 13 4 13 16 0 9 7 9 2
22 11 13 2 16 16 15 9 13 2 0 9 13 10 9 2 9 7 13 13 0 9 2
16 2 13 15 1 15 2 16 4 0 9 9 3 3 13 2 2
25 9 1 9 13 14 0 3 13 2 13 4 7 13 0 2 3 0 9 2 16 3 15 13 3 2
8 1 12 9 13 13 0 9 9
2 11 2
26 0 9 9 2 15 13 13 9 9 0 9 14 1 0 9 2 4 13 4 13 1 9 1 9 12 2
27 1 9 0 9 9 2 15 15 1 10 9 13 2 1 9 0 9 15 13 9 9 9 0 9 11 11 2
25 1 10 9 13 10 9 3 0 2 10 9 13 0 3 1 15 2 16 13 1 9 9 0 9 2
13 0 9 9 9 13 12 9 7 4 13 12 9 2
15 13 13 3 9 11 2 11 2 11 2 11 7 0 9 2
27 1 0 9 15 13 1 9 12 2 1 9 9 1 0 9 7 1 0 9 13 4 9 13 1 9 3 2
24 1 9 9 12 15 7 9 3 13 2 7 0 9 4 3 13 1 9 9 9 9 1 11 2
10 9 15 13 1 9 0 9 14 3 2
15 0 9 13 3 12 9 1 12 9 1 0 9 12 9 2
6 3 13 12 9 0 2
5 9 13 9 7 9
2 11 2
19 1 0 9 9 9 4 13 0 0 9 11 11 2 1 11 1 0 11 2
19 1 0 9 0 9 13 9 0 0 9 1 0 11 0 9 1 0 9 2
17 12 9 2 15 3 4 0 13 15 1 9 2 13 1 9 13 2
15 1 9 13 9 3 12 9 2 1 15 12 3 13 0 2
20 9 13 1 9 1 9 9 9 7 13 15 0 9 3 0 3 7 0 9 2
24 3 13 9 1 9 2 1 9 3 13 1 9 7 3 9 3 7 9 13 1 9 7 9 2
8 1 0 9 13 14 7 9 2
8 1 9 13 0 9 0 11 2
22 3 13 11 9 11 9 2 11 11 2 13 1 0 9 1 9 3 3 9 12 9 2
8 11 7 11 1 9 1 0 9
8 9 9 9 11 11 1 0 9
29 10 9 2 9 7 9 2 0 0 2 10 9 13 1 9 2 15 4 3 3 13 16 9 0 0 9 7 9 2
47 3 1 9 2 3 15 3 13 0 0 9 2 3 10 9 3 13 10 9 2 10 9 7 10 0 9 2 3 4 13 15 0 9 9 9 2 9 2 9 7 0 0 9 1 10 9 2
13 13 13 2 16 15 13 9 0 9 7 0 9 2
17 13 15 3 7 9 0 9 2 1 9 0 2 7 9 0 9 2
37 13 14 1 15 2 16 0 15 0 9 9 0 0 9 13 1 9 1 15 2 15 13 3 2 1 9 9 2 0 1 10 0 9 0 9 13 2
38 13 14 1 15 2 16 0 9 9 0 9 2 9 0 9 7 0 9 9 13 1 9 2 15 10 0 9 13 2 15 13 7 1 10 9 15 13 2
29 13 1 3 2 13 15 10 9 13 1 0 7 0 0 9 7 13 15 9 10 9 13 1 9 10 0 9 2 2
29 13 0 2 16 3 13 13 1 9 2 15 3 16 15 0 13 0 0 9 11 7 11 2 1 0 9 9 0 2
20 9 1 11 7 1 11 13 1 15 15 3 16 14 12 1 10 9 10 9 2
11 13 15 9 10 9 2 14 3 10 9 2
8 11 13 10 9 7 10 9 2
18 9 0 9 7 10 9 7 9 2 16 7 9 2 1 15 15 13 2
14 15 13 11 16 10 0 9 2 0 16 10 0 9 2
42 13 13 2 16 9 1 11 7 1 11 15 11 14 3 2 7 7 3 13 7 16 9 10 9 13 14 10 9 1 0 9 2 7 3 15 9 10 0 7 0 9 2
39 1 11 3 9 1 11 13 10 0 9 2 7 13 1 15 3 0 9 2 16 15 15 1 15 14 13 2 13 3 12 1 9 2 15 13 7 10 9 2
16 7 9 11 1 15 13 3 3 9 10 9 1 11 16 15 2
26 10 9 3 13 3 3 2 3 7 3 0 11 13 10 0 9 7 10 0 9 1 11 7 1 9 2
6 15 15 1 15 13 2
35 15 3 7 15 3 2 16 16 4 13 1 0 2 0 9 13 3 2 3 2 3 7 1 0 9 2 16 13 1 15 2 13 1 15 2
4 9 1 9 12
5 13 15 0 0 9
2 11 2
20 0 0 9 1 0 0 9 12 4 13 1 9 1 9 11 2 9 11 2 2
24 0 9 2 3 0 1 0 11 2 4 13 0 9 1 11 1 11 2 7 1 0 9 12 2
11 3 15 13 0 9 9 0 9 11 11 2
21 1 11 13 9 9 9 1 0 9 2 1 11 13 9 9 9 11 1 9 9 2
22 1 0 9 4 1 0 11 13 12 0 9 9 1 0 9 12 2 15 13 3 9 2
16 0 9 13 3 12 2 9 0 9 7 1 10 9 1 11 2
21 0 9 13 12 2 9 0 11 1 0 11 1 9 9 0 9 1 10 0 9 2
9 11 7 11 1 9 1 0 9 11
2 11 2
33 9 9 0 9 11 11 7 9 9 9 9 11 11 15 1 9 1 9 3 13 1 9 9 2 15 1 9 13 9 9 0 9 2
19 9 13 9 0 9 1 0 9 11 7 13 0 9 11 1 12 0 9 2
11 1 11 15 1 9 0 9 3 13 9 2
8 9 11 11 13 9 1 0 2
18 13 2 16 16 15 13 9 2 13 3 15 2 15 15 11 13 13 2
11 4 13 3 0 9 11 1 0 0 9 2
21 9 11 13 3 3 3 2 16 9 1 9 2 3 15 3 13 9 2 4 13 2
6 9 9 1 11 7 11
2 11 2
19 0 9 1 0 9 13 9 11 11 1 9 2 15 3 13 1 0 9 2
31 2 1 9 13 13 0 9 2 3 15 7 13 13 1 10 0 9 7 13 15 1 15 9 2 15 15 13 2 2 13 2
8 1 0 13 9 13 9 9 2
8 9 9 4 13 1 15 13 2
12 9 3 13 0 9 9 1 9 9 1 9 2
28 1 9 9 2 15 13 9 0 7 0 0 9 2 13 9 0 9 7 9 2 9 2 9 7 9 0 9 2
22 1 0 9 15 13 9 0 9 11 11 2 0 0 9 11 11 2 10 9 7 9 2
5 0 9 1 9 12
3 13 9 9
22 12 1 0 9 1 0 9 9 11 11 1 9 0 9 13 2 2 13 9 9 2 2
21 13 4 14 10 9 2 16 4 13 0 9 9 2 2 13 9 0 9 9 2 2
28 1 0 2 0 9 13 3 9 12 2 15 10 7 15 10 2 7 13 3 9 13 9 9 1 12 9 0 2
7 15 13 0 14 0 9 2
28 9 11 13 10 9 1 9 2 3 0 11 2 1 1 0 9 9 9 2 13 9 7 13 15 9 1 9 2
10 16 9 10 9 4 13 4 9 13 2
25 14 1 9 11 2 7 3 2 7 3 3 2 11 4 0 9 13 0 9 1 10 9 1 11 2
9 11 11 15 1 10 9 13 3 2
8 9 1 0 9 13 3 0 2
15 3 15 1 0 9 1 11 7 1 11 13 13 0 9 2
7 0 9 13 1 0 9 2
40 13 2 14 0 9 2 16 3 13 1 9 1 0 9 10 9 2 15 13 3 13 1 9 15 3 0 9 2 0 7 0 2 13 4 9 1 0 9 0 2
7 13 2 16 15 3 13 2
26 9 0 9 13 0 7 0 9 2 15 15 13 1 9 13 15 1 0 0 9 1 9 9 12 9 2
6 9 9 13 13 9 2
18 1 9 7 9 9 7 13 0 7 0 9 1 9 2 13 9 11 2
17 15 9 13 2 13 9 2 7 13 15 1 15 9 13 10 9 2
9 1 15 14 13 7 15 15 13 2
10 12 9 9 7 9 9 13 13 3 2
22 13 7 1 15 3 12 9 9 9 7 3 1 9 0 2 0 9 15 13 3 3 2
10 9 1 15 13 16 9 2 7 9 2
32 10 9 7 9 0 9 7 9 1 0 9 13 3 10 0 9 7 9 2 15 15 3 9 0 1 11 13 1 9 0 9 2
16 3 15 13 1 0 9 2 1 15 10 9 1 9 9 13 2
12 9 7 9 13 10 9 3 7 3 13 3 2
22 15 3 4 0 9 13 10 2 0 9 9 2 2 15 3 15 13 13 3 1 11 2
1 3
6 9 9 13 7 11 2
19 0 9 3 13 14 12 9 9 9 1 9 1 12 9 9 1 9 12 2
21 1 12 9 9 3 9 1 11 13 12 9 2 16 1 9 15 13 14 12 9 2
30 9 1 9 9 1 0 9 7 11 1 12 9 1 9 12 2 12 7 1 12 9 1 9 12 2 12 13 0 9 2
10 11 13 11 7 13 0 0 9 9 2
14 1 9 12 2 12 13 0 12 9 2 9 0 9 2
22 9 9 1 11 13 3 12 9 2 15 13 2 16 3 1 9 12 4 13 10 9 2
21 9 9 13 3 3 1 12 9 0 16 1 9 12 2 15 13 14 1 12 9 2
18 0 9 0 0 13 1 9 12 9 1 9 1 9 12 9 2 9 2
23 9 7 13 13 9 1 9 12 9 14 1 12 9 2 7 2 12 9 1 12 0 9 2
19 11 2 15 13 10 9 3 16 9 9 2 13 0 9 0 9 0 9 2
27 0 0 9 0 0 9 11 2 11 13 10 0 9 1 12 5 1 9 13 3 9 0 9 9 7 9 2
17 9 11 2 11 1 9 3 13 1 9 9 1 9 9 1 9 2
4 0 9 9 2
47 0 9 9 1 9 9 0 9 2 15 1 9 13 9 11 7 11 2 11 11 7 11 2 15 13 3 3 1 0 9 0 0 9 2 9 2 1 9 11 1 11 2 10 9 15 13 2
17 2 13 4 2 16 13 1 9 9 1 11 2 2 13 9 11 2
9 11 7 13 1 10 9 1 11 2
3 0 9 2
19 1 9 13 14 9 9 9 2 9 2 15 15 9 13 1 9 9 11 2
7 1 9 13 3 11 12 2
25 0 9 2 15 9 3 3 13 9 9 12 2 12 2 13 3 0 2 16 10 9 13 7 9 2
17 11 7 11 13 1 2 3 1 0 9 11 1 9 11 1 11 2
14 1 9 15 13 2 16 9 11 13 9 0 9 9 2
14 10 9 13 3 0 2 16 1 15 13 7 11 11 2
27 15 13 9 1 9 2 9 2 9 2 2 9 2 0 9 2 9 2 7 9 2 9 2 13 3 0 2
7 9 9 15 15 3 13 2
3 0 0 9
3 0 2 9
31 1 0 9 13 0 2 9 13 9 1 9 1 9 1 0 9 0 9 2 1 15 15 0 9 9 13 9 1 0 9 2
16 0 9 9 13 7 0 0 9 9 1 0 9 0 2 11 2
17 3 15 10 9 13 3 12 12 0 9 1 3 16 12 9 9 2
22 7 16 15 0 0 9 13 13 2 0 9 9 15 10 9 13 3 1 9 12 9 2
17 3 15 13 1 9 2 3 13 9 9 1 9 3 12 9 9 2
20 3 15 13 7 0 9 2 15 13 1 0 2 11 1 9 1 9 3 9 2
24 0 13 3 9 2 3 15 13 0 9 1 3 12 12 9 2 15 13 0 1 0 0 9 2
18 3 0 9 1 0 9 2 15 13 0 2 11 2 13 1 0 9 2
14 0 9 15 13 1 0 12 1 3 16 12 9 9 2
25 16 9 1 9 0 0 9 13 13 1 0 9 3 0 2 9 0 9 11 12 1 0 9 13 2
32 1 9 3 9 12 13 1 9 1 9 0 9 7 13 1 12 5 1 12 9 2 7 15 13 3 2 16 15 10 9 13 2
27 1 9 13 1 3 0 9 2 1 15 15 9 3 13 2 3 9 13 7 1 9 3 13 1 12 9 2
7 3 13 1 9 12 9 2
13 9 1 0 9 0 2 11 3 13 9 0 9 2
10 3 15 13 1 9 1 12 9 9 2
6 9 11 3 3 13 2
22 3 9 15 13 1 12 9 2 1 9 13 10 9 12 7 1 9 13 1 12 9 2
8 3 13 0 9 1 12 9 2
9 1 0 9 15 13 7 11 0 2
16 1 9 15 13 1 12 9 7 1 9 13 14 1 12 9 2
5 3 13 12 9 2
12 3 0 1 0 9 2 11 0 13 0 9 2
10 13 16 0 0 9 1 9 12 9 2
14 3 7 10 9 13 7 1 9 15 13 1 12 9 2
9 1 9 13 10 0 9 12 9 2
13 9 0 9 11 13 1 0 12 9 1 0 12 2
12 1 9 9 15 3 13 13 3 1 0 9 2
10 1 9 15 9 11 13 1 12 9 2
6 9 13 1 12 9 2
24 3 3 15 1 0 2 11 13 9 0 0 0 11 2 7 15 1 12 7 12 9 1 9 2
4 9 1 0 9
1 9
11 0 9 0 9 13 1 15 3 0 9 2
9 1 10 9 15 13 3 14 3 2
26 9 1 12 9 13 1 0 12 9 2 9 1 0 9 15 9 7 9 15 3 13 13 1 0 9 2
10 15 15 13 2 16 3 13 10 9 2
26 3 12 0 9 1 0 9 0 9 4 12 2 9 13 1 0 9 7 0 9 7 1 0 2 11 2
18 10 0 9 15 9 13 3 13 2 7 15 3 13 10 0 0 9 2
21 1 0 9 9 9 1 0 9 13 2 16 4 9 1 9 0 13 13 9 0 2
14 0 9 2 0 1 9 9 2 15 1 0 9 13 2
9 3 13 0 1 0 0 0 9 2
7 3 13 9 9 0 9 2
34 9 3 15 3 0 9 2 3 7 2 16 13 3 3 0 2 13 3 13 2 16 9 4 13 13 0 9 16 0 2 7 3 0 2
38 9 1 0 11 2 15 15 13 1 0 12 9 2 3 11 0 9 13 1 0 9 1 10 9 9 12 12 9 2 13 3 1 9 12 2 9 12 2
25 1 10 0 9 15 3 13 9 1 9 9 2 15 3 13 0 9 2 15 3 4 13 3 13 2
13 1 9 0 0 9 15 13 13 7 1 0 9 2
9 15 13 9 1 10 0 0 9 2
10 0 9 2 0 9 2 0 0 9 2
4 9 9 13 13
2 11 2
25 1 9 1 9 0 9 2 0 9 7 11 13 3 0 9 10 9 9 9 7 9 11 2 11 2
28 13 1 15 13 7 0 9 2 15 4 13 13 1 9 10 0 9 11 7 0 9 7 1 9 0 0 9 2
17 10 9 4 13 1 9 9 7 9 7 3 7 1 0 0 9 2
17 9 9 13 7 9 2 15 4 13 13 0 9 3 1 0 9 2
27 1 11 2 11 13 9 0 9 3 0 1 9 11 11 1 10 9 2 16 0 9 13 1 0 0 9 2
4 0 9 13 9
3 0 11 2
18 9 0 9 1 9 9 9 1 12 9 13 0 0 9 0 0 9 2
15 0 9 1 0 9 13 0 9 2 13 9 11 2 11 2
14 12 12 9 13 1 9 12 0 9 0 9 7 11 2
15 0 12 1 9 12 9 9 13 9 1 0 9 0 9 2
17 3 11 2 3 2 9 11 9 2 13 9 0 9 1 12 12 2
23 0 9 9 2 15 13 1 12 9 2 15 1 0 12 9 13 1 12 7 12 9 9 2
6 11 15 3 1 9 13
4 11 13 9 2
4 9 9 4 13
46 0 9 11 11 3 13 1 0 0 9 1 0 11 9 1 9 2 16 11 13 9 2 1 15 15 1 9 1 11 13 9 0 9 11 11 2 11 7 11 9 2 0 9 11 9 2
25 9 12 9 0 9 15 13 1 9 0 9 2 16 15 0 9 13 1 9 1 9 0 0 9 2
12 11 3 13 13 9 13 9 0 1 9 11 2
33 10 9 1 11 2 11 2 11 13 11 1 10 9 2 16 4 13 1 12 7 12 5 0 9 2 16 1 15 13 3 0 9 2
18 11 15 13 1 9 12 1 0 9 12 9 0 9 1 12 9 9 2
13 1 9 9 13 9 14 1 12 7 12 9 9 2
19 11 2 11 3 13 2 16 1 9 1 0 9 13 3 3 13 0 9 2
21 1 15 14 0 9 3 13 0 9 2 3 13 7 13 9 11 3 1 0 9 2
33 1 9 0 0 9 0 9 1 11 15 12 9 13 2 16 11 9 1 12 2 9 13 15 9 2 15 9 11 13 1 9 12 2
18 13 15 15 12 9 0 9 2 15 4 13 1 2 3 0 9 2 2
25 1 9 10 9 11 13 1 0 0 9 7 13 0 9 1 3 0 9 1 14 12 9 0 9 2
11 9 11 9 15 13 13 3 12 0 9 2
19 10 12 9 1 12 2 9 13 0 9 11 3 12 9 9 1 0 9 2
21 12 9 15 13 13 9 2 15 13 11 9 3 13 7 0 9 1 0 9 13 2
20 1 0 9 16 9 1 0 9 2 7 1 0 9 13 1 11 11 3 3 2
19 0 9 13 2 16 0 9 1 9 15 0 1 9 13 1 10 0 9 2
8 11 1 9 9 9 1 9 9
2 11 2
41 9 9 0 9 2 11 2 4 13 2 16 4 1 9 0 9 3 13 9 0 9 2 7 15 1 9 1 15 2 3 0 9 11 2 3 9 2 1 9 13 2
28 13 15 9 9 7 9 9 11 11 11 1 9 1 9 9 11 2 15 4 13 1 9 1 12 2 9 12 2
22 9 11 13 0 9 1 9 9 2 15 13 0 9 1 9 0 9 9 1 0 9 2
47 9 9 1 11 13 1 15 2 16 9 9 4 1 9 7 1 0 9 9 2 1 15 13 11 0 16 0 9 2 13 1 9 0 0 9 7 16 1 0 9 3 13 9 1 9 11 2
15 0 9 11 13 3 0 13 9 1 15 2 3 9 13 2
24 9 9 13 3 0 13 9 2 15 13 3 1 0 7 0 9 9 7 9 1 9 9 9 2
9 9 1 9 9 1 2 0 9 2
2 11 2
16 9 1 0 7 0 9 13 13 9 9 1 0 9 9 9 2
8 11 15 13 9 9 11 11 2
26 1 0 9 1 0 7 0 9 2 15 13 1 10 9 0 9 2 13 13 9 0 1 9 0 9 2
32 9 9 1 11 3 1 15 13 7 1 0 9 2 15 4 0 7 0 9 13 13 9 0 9 1 9 0 9 1 0 9 2
30 9 9 11 9 1 9 0 9 3 13 2 16 1 0 9 15 13 12 0 0 9 7 16 3 4 13 10 0 9 2
19 10 0 9 7 13 13 1 9 2 16 15 1 15 13 2 0 9 2 2
12 9 0 9 4 1 10 9 13 1 12 9 2
37 1 9 11 13 1 12 9 9 0 0 11 2 11 2 2 15 4 1 0 9 13 0 9 11 2 7 0 7 0 9 9 11 11 2 11 2 2
9 9 0 12 15 9 3 13 13 2
50 1 9 9 1 9 9 9 0 9 13 13 10 9 9 1 0 7 0 9 2 15 13 1 9 9 13 2 16 9 0 9 13 9 9 2 16 13 9 0 9 7 15 13 9 9 1 9 0 9 2
24 1 9 11 13 2 16 0 9 1 9 9 13 3 9 11 2 15 3 11 13 12 9 9 2
18 11 15 13 3 1 0 9 1 0 11 7 3 1 11 13 9 11 2
15 9 0 9 1 11 15 1 0 9 13 9 9 0 1 9
5 13 3 9 1 11
2 11 2
14 0 0 9 1 11 11 13 3 1 0 9 1 11 2
37 9 15 13 1 15 2 16 13 0 9 2 3 1 9 1 0 9 0 9 1 11 7 1 9 9 1 11 1 11 1 0 9 14 12 9 9 2
26 9 4 3 13 7 9 11 1 0 3 0 9 1 0 9 1 11 1 0 11 1 9 14 12 9 2
13 1 9 13 9 13 13 1 12 9 12 12 9 2
24 0 9 3 13 3 1 9 2 13 15 7 13 2 16 12 1 0 4 3 13 1 10 9 2
28 11 1 9 9 13 2 16 13 0 7 16 9 2 15 13 10 9 1 3 0 9 1 0 9 2 13 0 2
19 9 13 7 9 2 15 15 1 0 9 13 13 7 15 10 9 3 13 2
16 0 11 13 0 9 1 10 9 1 0 9 1 11 2 11 0
6 1 11 15 13 1 11
15 9 11 9 2 13 9 2 16 1 0 9 13 12 0 9
2 11 2
16 2 9 1 9 13 12 9 2 15 15 1 11 13 16 9 2
26 3 4 13 1 0 0 9 2 11 2 15 13 1 0 9 2 2 13 15 0 9 9 11 11 0 2
22 15 1 9 13 14 1 0 9 2 16 3 1 9 0 0 9 13 10 9 1 11 2
19 0 9 3 3 13 13 11 11 7 11 0 9 13 2 3 15 3 13 2
14 2 15 15 7 13 2 16 3 3 0 9 11 13 2
21 13 15 13 7 3 2 7 1 9 1 0 9 15 13 13 0 9 1 9 2 2
17 3 3 9 13 0 9 9 7 12 9 15 9 13 1 0 9 2
24 0 9 7 13 2 16 10 9 15 13 2 2 3 4 9 15 13 7 3 4 3 13 2 2
20 0 9 2 15 15 13 1 0 9 2 13 11 2 15 15 0 13 1 11 2
12 2 9 13 3 0 2 13 4 1 12 9 2
22 3 4 9 13 7 12 3 0 9 4 13 1 9 2 16 4 13 7 13 1 9 2
10 11 13 1 15 0 9 14 3 9 2
59 14 15 13 7 1 10 9 3 13 2 7 15 3 9 9 13 0 9 2 2 13 9 2 15 1 9 13 1 9 7 9 0 9 2 1 15 0 13 1 10 9 1 11 2 11 2 11 2 11 7 11 2 11 3 7 1 11 2 2
27 1 0 9 1 9 15 0 9 13 9 13 15 9 1 9 2 7 16 9 14 13 7 9 1 12 9 2
31 2 11 2 11 7 11 4 13 13 3 0 9 9 2 16 4 15 1 0 9 13 2 7 0 9 13 1 0 0 9 2
13 11 13 3 3 0 7 1 15 13 7 10 9 2
17 13 9 2 16 1 0 9 1 9 9 4 13 12 0 9 2 2
6 1 11 13 1 0 9
4 11 2 11 2
16 1 0 9 1 0 9 0 0 9 13 9 11 11 11 0 2
35 2 14 9 13 13 1 9 3 2 16 0 9 9 13 9 1 0 9 2 2 13 9 2 15 3 13 0 9 1 11 2 11 7 11 2
22 0 9 13 1 11 16 0 9 2 7 1 9 11 11 1 11 13 3 1 0 9 2
11 1 0 9 9 13 10 9 1 0 9 2
13 1 11 11 13 11 2 3 15 1 9 13 11 2
15 16 13 11 1 0 9 9 2 9 13 1 9 1 9 2
11 2 13 3 0 9 2 15 13 0 9 2
24 3 3 13 2 3 15 1 15 13 2 1 0 9 11 7 11 2 9 1 9 13 3 0 2
20 0 12 0 9 15 13 2 16 13 1 11 2 1 11 1 11 7 1 11 2
14 13 15 1 0 9 7 13 2 16 15 13 0 9 2
8 1 0 9 15 13 13 2 2
8 0 9 9 13 3 0 9 2
37 1 0 9 13 9 0 9 14 1 0 9 2 3 0 2 1 11 2 12 2 12 2 7 0 14 1 0 9 1 0 9 1 9 1 0 9 2
30 2 10 9 4 13 9 12 9 1 9 1 9 9 7 1 9 13 10 9 3 13 2 2 13 0 9 0 11 11 2
5 9 1 11 13 9
7 0 9 3 13 0 9 11
18 0 0 9 13 3 10 9 7 9 1 0 9 13 14 1 0 9 2
26 1 11 15 9 0 9 13 9 12 2 7 12 2 9 7 9 10 9 13 3 9 0 7 0 9 2
14 1 9 3 15 9 9 9 11 11 11 13 12 9 2
31 13 13 11 2 1 9 13 1 9 9 2 7 11 2 0 9 2 0 9 2 2 0 9 3 13 11 2 15 13 9 2
31 16 13 9 2 16 15 13 9 2 13 13 0 9 2 11 13 9 2 7 1 9 13 0 9 1 9 9 11 1 9 2
18 9 13 1 9 1 9 2 3 7 3 9 13 12 9 1 12 9 2
34 2 0 1 9 13 12 7 12 9 9 2 7 13 13 15 2 2 13 11 7 13 15 7 12 9 2 1 15 15 0 9 13 13 2
19 12 1 9 3 13 2 2 15 13 1 9 13 9 9 1 0 9 2 2
28 1 9 9 13 0 9 3 1 9 2 7 14 1 0 9 2 16 15 1 9 1 3 0 9 13 13 0 2
15 2 9 9 15 7 13 9 2 9 1 9 7 0 9 2
16 13 4 3 13 2 16 9 9 13 2 2 13 9 0 9 2
26 1 9 1 9 15 9 13 13 10 9 2 1 15 9 4 13 1 9 2 0 9 7 13 0 9 2
26 12 9 1 12 9 2 12 9 1 12 9 7 1 0 9 2 0 2 0 9 2 13 3 12 9 2
11 2 12 9 15 13 3 2 0 9 3 2
18 15 13 9 3 14 1 0 9 2 13 13 0 9 3 1 0 9 2
14 9 13 3 1 9 7 9 15 15 13 1 0 9 2
17 16 3 13 2 13 15 1 15 13 2 2 13 0 9 11 11 2
23 1 0 9 1 0 9 13 9 0 11 2 15 3 13 1 12 9 9 7 13 0 9 2
23 9 9 13 3 0 9 2 12 0 11 2 15 15 1 0 9 13 14 1 9 12 9 2
20 3 0 9 9 2 0 2 13 1 9 1 9 2 7 9 13 14 1 9 2
22 1 0 9 13 9 1 9 7 1 9 1 0 0 9 13 10 3 7 3 0 9 2
22 3 16 1 0 9 7 1 9 15 3 13 9 0 9 2 0 9 7 9 1 9 2
15 2 13 1 9 7 0 9 2 15 13 9 9 0 9 2
18 13 15 3 1 9 0 9 7 3 3 3 0 9 2 2 13 11 2
16 0 9 13 9 0 7 0 9 3 1 9 3 1 9 9 2
19 1 9 3 13 3 3 1 0 9 2 16 9 4 13 13 10 9 3 2
14 2 0 9 13 1 15 3 3 2 16 4 13 15 2
23 1 15 13 9 14 3 3 7 3 4 13 1 9 2 2 13 11 11 2 0 0 9 2
16 9 15 9 15 9 13 1 0 9 3 1 9 1 0 9 2
13 1 9 13 9 11 1 0 9 7 11 1 0 2
4 11 15 13 11
26 12 9 13 0 9 11 11 2 12 2 2 16 4 15 13 11 7 13 15 13 1 9 0 9 3 2
24 0 0 9 7 9 12 2 11 11 1 11 1 9 10 0 9 13 12 1 9 9 1 11 2
30 10 0 9 15 3 13 9 11 2 15 3 1 0 9 13 0 9 1 0 2 0 2 9 9 1 3 0 0 9 2
13 1 9 13 0 9 2 3 9 9 13 2 9 2
20 1 9 0 9 13 0 9 2 1 15 13 9 2 13 11 0 9 11 11 2
30 0 9 1 11 13 3 9 2 1 9 13 9 7 10 9 11 7 11 2 15 3 13 1 9 1 11 1 2 11 2
10 2 10 9 13 1 15 1 0 9 2
24 13 1 10 9 2 16 15 13 7 10 9 2 2 13 11 11 1 12 1 0 0 2 9 2
7 0 9 7 11 9 13 2
19 1 1 3 0 9 15 3 9 13 1 9 1 0 9 7 13 14 9 2
11 13 7 13 1 0 9 7 13 0 9 2
5 1 11 2 3 2
11 2 3 13 10 9 2 2 13 0 11 2
4 11 13 13 9
2 11 2
26 0 9 9 11 0 11 11 13 2 16 13 13 13 0 9 1 11 0 9 2 16 15 9 13 9 2
15 2 13 10 9 3 0 2 7 13 9 13 9 10 9 2
13 1 9 13 4 13 9 1 9 2 9 7 9 2
25 9 13 13 2 16 15 13 1 9 13 2 2 13 11 1 0 9 1 9 11 1 11 1 11 2
4 9 11 11 13
2 11 2
27 0 9 0 0 9 2 11 2 13 9 11 1 9 1 0 9 9 1 0 9 9 9 1 11 1 11 2
17 1 9 9 3 13 0 9 0 12 9 1 0 9 1 0 9 2
9 1 9 1 11 13 12 2 12 2
3 1 0 9
15 11 13 1 9 9 12 2 9 11 2 11 9 0 9 2
7 16 0 4 13 11 11 2
23 11 11 13 2 16 1 9 9 3 13 11 11 7 1 9 0 9 15 14 13 1 11 2
18 15 1 15 1 9 9 13 12 9 9 3 2 16 15 13 12 9 2
5 11 7 0 13 9
2 11 2
10 0 0 0 9 13 1 9 0 9 2
2 11 2
23 0 9 13 1 9 1 0 9 9 12 2 9 2 1 15 15 13 7 0 9 11 11 2
18 15 3 13 9 1 12 2 9 1 0 9 9 1 11 12 2 12 2
13 0 13 9 2 7 7 0 9 13 9 1 9 2
20 11 13 12 9 3 1 0 9 2 1 0 0 9 15 13 7 11 7 11 2
20 1 11 15 13 13 9 11 11 2 15 13 1 0 9 9 1 0 0 11 2
21 11 13 9 9 1 11 1 12 2 9 7 12 9 1 9 13 0 9 0 11 2
20 11 2 15 13 1 0 9 9 2 13 3 14 13 1 12 2 9 9 11 2
2 11 2
21 1 11 13 1 9 12 2 9 9 2 7 7 15 13 14 12 9 12 2 9 2
17 0 11 11 13 1 9 0 11 3 1 12 9 11 1 0 9 2
8 1 9 3 14 13 0 11 2
18 11 15 1 0 9 13 1 0 11 2 15 1 9 13 14 0 9 2
2 11 2
20 1 9 9 1 0 9 11 15 3 13 0 11 2 15 13 11 12 2 12 2
9 9 9 11 15 13 3 9 9 2
18 3 1 12 2 9 13 11 7 7 9 11 7 11 13 1 0 9 2
2 11 2
30 1 12 2 9 0 9 13 11 0 9 1 12 2 9 1 0 9 11 1 11 11 2 15 10 9 13 1 9 9 2
16 9 13 0 9 9 9 11 11 1 9 0 11 12 2 12 2
19 10 9 3 0 13 1 9 1 9 9 2 7 1 0 9 13 12 9 2
12 9 9 13 9 11 2 9 9 1 0 9 2
25 9 13 1 11 12 2 12 7 1 9 11 1 9 1 11 13 10 9 1 9 9 1 12 9 2
4 11 13 0 9
2 11 2
30 0 0 9 11 2 11 2 15 13 4 0 9 1 12 9 9 13 1 9 9 2 15 4 3 13 1 11 0 9 2
11 1 10 9 13 16 0 0 9 11 11 2
17 9 4 15 13 13 7 1 0 9 2 7 14 1 9 0 9 2
16 0 9 11 11 1 9 1 9 11 11 13 1 9 0 9 11
1 3
17 0 9 11 13 9 9 2 10 9 4 13 9 9 1 0 11 2
21 9 2 15 15 13 12 2 9 1 11 2 15 13 11 11 7 11 7 11 11 2
22 0 9 0 9 11 4 13 9 9 1 12 9 7 12 9 1 9 1 9 0 9 2
18 0 9 11 13 1 9 1 0 11 0 9 1 0 9 1 12 9 2
17 1 9 13 3 1 9 12 9 11 11 2 0 9 0 0 9 2
5 9 1 9 1 9
2 11 2
30 9 15 11 9 0 11 2 0 2 9 1 9 2 15 13 7 1 0 9 2 7 15 9 9 1 9 0 9 9 2
17 9 9 0 9 11 13 1 9 9 2 15 13 0 9 12 9 2
41 0 9 4 9 13 1 11 2 0 11 2 11 2 11 2 11 7 11 2 9 4 13 1 0 9 2 11 2 9 7 11 2 7 3 1 11 7 11 1 11 2
19 9 0 0 9 4 1 9 11 3 13 9 1 9 9 7 9 1 9 2
31 9 1 0 9 2 9 2 12 9 2 12 9 2 13 0 13 1 11 11 2 0 9 12 2 12 12 11 12 2 11 2
7 11 1 9 1 9 13 3
21 2 16 13 1 0 12 9 2 13 15 1 15 13 2 2 13 9 11 0 0 9
58 9 0 0 9 11 11 1 9 1 0 9 13 2 16 1 9 9 14 0 9 2 15 13 1 9 2 4 1 1 0 15 9 9 13 9 11 2 11 2 2 11 2 11 2 2 11 2 11 2 7 0 9 9 11 11 1 11 2
24 15 13 1 0 9 0 9 0 7 3 7 0 9 2 7 3 15 3 1 10 0 9 13 2
13 2 1 9 11 4 13 3 1 9 1 0 9 2
12 13 15 2 16 13 13 9 3 1 0 9 2
17 1 9 4 15 13 3 2 3 3 1 9 1 9 3 3 13 2
24 15 13 3 0 9 2 2 13 11 11 7 3 13 2 16 15 10 9 13 1 3 0 9 2
21 2 9 11 13 1 1 0 9 0 9 2 15 13 2 1 9 0 9 0 9 2
19 14 16 4 3 1 15 13 10 9 2 7 13 15 3 9 0 0 9 2
31 7 1 10 9 15 13 10 0 9 13 1 9 1 11 2 13 4 15 1 15 9 1 10 9 2 15 15 13 3 0 2
23 1 0 9 15 15 1 9 3 13 7 3 4 13 13 2 3 15 11 13 1 9 2 2
8 11 13 2 9 13 2 2 2
20 11 11 13 1 9 12 1 0 9 0 11 7 3 3 0 9 13 1 11 2
19 1 9 9 0 9 9 13 0 1 0 9 12 1 9 7 12 0 9 2
28 13 15 7 11 2 15 1 9 14 13 1 0 9 7 1 12 2 9 3 13 1 11 12 2 12 1 9 2
5 2 3 13 3 2
27 1 9 15 13 12 9 9 2 1 15 7 11 11 2 15 13 3 0 9 9 7 13 7 1 0 9 2
9 1 11 15 3 13 1 0 9 2
15 0 9 1 10 9 13 12 9 2 1 11 3 12 9 2
11 13 3 1 0 9 2 7 13 3 13 2
23 10 0 9 2 15 13 1 9 2 13 1 9 1 12 9 7 13 13 9 10 0 9 2
29 1 9 4 13 1 9 11 13 1 12 9 11 11 2 15 15 13 1 12 9 2 7 0 9 15 15 13 2 2
23 0 9 4 1 9 13 1 12 1 12 9 7 1 9 0 11 15 13 2 16 15 13 2
20 1 0 9 15 1 9 13 7 1 0 9 2 15 4 13 0 9 12 9 2
20 2 0 9 1 9 0 9 13 9 13 9 1 0 9 7 13 0 9 9 2
20 7 3 13 3 0 0 9 2 16 4 13 13 9 7 1 15 9 9 13 2
16 16 3 13 1 15 1 0 12 9 2 13 15 1 15 13 2
47 1 11 13 0 9 9 7 3 15 13 0 2 7 16 1 9 1 11 13 0 9 2 2 13 11 11 7 13 2 16 15 3 1 9 13 7 0 9 2 15 15 1 9 9 0 13 2
16 2 9 9 11 11 1 9 9 13 7 13 7 9 1 9 2
24 1 11 13 3 1 12 9 3 16 3 2 0 13 15 1 15 2 1 11 7 1 11 2 2
26 1 9 1 15 15 13 9 9 2 15 0 9 13 2 7 7 1 0 9 13 9 1 9 0 9 2
22 2 15 13 9 9 9 1 12 2 0 9 9 7 9 9 13 1 9 0 0 9 2
29 1 9 13 15 9 1 9 9 11 2 0 9 13 3 10 9 2 7 9 11 11 2 1 15 13 0 9 2 2
4 0 9 0 9
4 0 9 3 13
6 12 9 13 1 0 9
2 11 2
31 10 9 2 1 15 4 13 0 0 9 11 2 11 2 12 2 12 2 2 4 15 3 13 13 0 9 1 10 0 9 2
23 14 1 9 0 0 9 2 12 9 2 13 1 9 9 9 0 2 0 7 3 0 9 2
33 1 9 9 2 15 13 0 9 1 9 1 9 1 9 14 7 0 1 9 9 1 11 13 2 15 13 1 0 9 1 0 9 2
20 1 15 9 13 3 0 11 2 7 1 0 9 1 9 9 3 0 9 13 2
17 0 9 9 13 9 0 12 0 9 1 12 9 7 1 9 9 2
16 9 11 13 1 9 11 3 1 0 9 0 9 1 0 9 2
20 10 9 1 0 9 0 1 9 1 9 0 9 13 7 13 14 1 0 9 2
13 9 9 11 1 9 13 2 16 13 1 0 9 2
39 7 2 16 15 0 13 1 9 2 13 3 3 2 7 16 15 15 9 13 3 1 15 2 16 4 11 1 0 9 3 13 2 13 15 1 9 0 9 2
39 11 11 13 1 9 1 9 10 9 0 2 7 13 9 1 9 2 15 13 1 9 0 9 3 3 13 1 9 2 2 15 2 15 13 2 13 0 9 2
27 13 10 9 1 15 2 3 15 13 1 12 1 15 2 16 9 11 13 9 1 9 2 15 4 13 9 2
14 9 1 15 13 2 16 4 13 12 9 1 9 2 2
58 1 9 11 11 13 2 16 15 7 11 11 2 15 3 1 0 9 1 9 12 2 12 1 11 13 0 9 1 9 9 2 13 9 3 2 2 11 13 1 11 13 2 16 13 3 0 9 2 13 7 1 0 9 0 9 7 13 2
16 9 3 13 1 9 9 11 2 15 1 0 12 3 13 2 2
32 0 9 15 3 13 1 9 1 0 9 9 1 0 1 9 0 9 1 0 0 9 2 2 13 1 9 0 3 1 15 13 2
22 1 10 9 1 11 7 1 11 4 15 1 15 0 2 15 13 9 11 2 13 2 2
6 3 14 7 3 1 9
11 0 9 11 11 13 0 9 3 1 12 9
39 2 13 4 3 2 14 16 4 15 13 2 2 13 1 9 9 11 11 1 0 9 2 12 9 2 2 15 13 1 0 0 0 9 1 11 0 0 9 2
16 2 13 15 2 16 13 3 13 1 12 9 7 13 1 9 2
22 3 15 13 0 2 16 3 13 13 7 13 0 0 9 1 0 9 1 12 9 2 2
22 1 9 15 1 11 13 9 11 7 3 4 13 13 0 0 0 9 13 13 0 9 2
45 16 4 15 7 9 13 2 13 4 7 3 1 0 0 9 9 1 11 2 2 1 9 13 13 2 7 16 4 3 15 13 1 9 2 3 15 1 9 13 9 13 9 7 9 2
13 0 9 13 13 3 3 2 13 15 9 9 2 2
22 13 9 2 13 11 11 1 0 9 0 2 2 13 4 15 1 11 11 0 1 11 2
23 13 15 10 9 2 1 9 4 15 13 1 9 0 9 7 13 2 16 15 15 13 2 2
19 1 0 9 13 0 0 9 1 9 0 0 9 1 9 9 12 1 11 2
27 0 9 4 3 13 13 1 0 11 7 1 0 11 1 0 9 9 0 11 2 10 9 13 3 0 9 2
19 3 1 9 15 1 9 11 11 1 0 9 11 11 13 0 9 11 11 2
22 1 11 13 1 11 0 0 9 2 15 4 15 13 1 12 9 3 13 1 0 9 2
20 1 9 7 3 13 0 9 7 3 1 9 15 1 9 0 9 13 0 9 2
14 2 9 9 7 9 15 13 2 7 9 15 3 13 2
19 1 9 4 13 12 9 7 12 9 13 14 1 9 0 16 10 0 9 2
21 1 10 9 12 9 4 15 13 7 1 9 0 2 7 3 4 13 1 12 2 2
19 9 2 15 13 0 7 0 9 2 13 1 9 10 0 9 3 3 3 2
28 0 9 2 15 1 9 1 12 9 1 9 13 7 13 16 9 2 3 3 7 13 2 10 9 13 3 9 2
24 2 9 1 9 15 3 13 2 7 16 4 13 2 3 15 3 13 2 2 13 11 2 11 2
2 9 9
5 0 9 1 0 9
11 1 9 15 1 0 9 13 11 11 7 11
2 11 2
19 1 3 0 0 9 4 13 0 0 9 9 1 0 11 7 13 1 9 2
23 9 0 9 3 13 12 1 0 9 12 9 2 16 9 9 1 0 9 7 9 3 13 2
26 0 13 1 10 9 11 1 11 9 12 2 12 9 2 2 0 11 11 13 9 1 12 12 9 0 2
32 11 13 7 1 0 9 0 9 2 7 1 0 15 13 11 11 2 1 15 15 13 0 9 1 9 2 7 11 7 11 11 2
6 9 12 0 9 1 15
26 11 15 0 9 13 16 9 1 9 2 3 13 1 0 9 0 9 2 16 9 1 11 15 3 13 2
2 11 2
17 3 13 9 9 11 11 2 0 1 0 0 9 1 0 9 11 2
15 1 9 12 12 9 13 0 11 11 2 0 13 11 11 2
8 11 13 1 11 3 1 9 9
2 11 2
36 1 0 9 1 12 9 1 0 9 1 11 13 1 15 11 11 11 2 9 9 7 11 1 0 0 9 2 7 0 9 11 11 1 11 11 2
22 1 9 13 1 10 9 2 7 11 13 1 0 9 9 12 0 9 1 9 12 12 2
26 2 1 11 15 3 13 2 7 1 9 12 4 1 15 13 1 2 9 2 1 0 9 11 1 11 2
20 15 15 3 3 13 2 7 13 4 3 2 16 4 15 15 13 1 0 9 2
27 0 9 15 3 13 7 9 15 14 13 13 2 7 1 9 1 11 4 15 13 2 2 13 1 9 11 2
36 10 0 9 13 10 9 2 2 16 0 9 9 13 9 9 9 9 1 9 2 7 7 3 7 13 0 2 16 4 13 1 0 9 1 11 2
18 0 9 4 15 13 1 9 1 0 9 16 9 1 0 9 1 11 2
9 13 0 1 9 2 14 1 9 2
26 2 3 3 13 13 11 0 1 0 2 1 11 13 9 12 0 0 0 9 1 12 9 1 0 12 2
23 1 9 12 9 15 3 3 13 0 0 9 12 2 15 13 0 9 11 11 2 12 2 2
3 11 13 9
2 11 2
28 1 9 0 9 1 11 2 9 12 9 2 13 11 11 1 11 11 12 2 12 2 12 2 12 1 12 9 2
18 0 11 13 10 12 2 9 9 7 3 1 12 9 13 10 0 9 2
25 1 0 9 0 9 13 1 0 9 11 2 11 2 15 13 1 9 11 1 0 0 7 1 11 2
7 2 13 15 15 3 3 2
48 13 4 2 16 1 0 0 9 13 3 10 0 9 2 3 1 9 1 9 11 11 2 2 13 0 11 2 15 0 12 0 9 1 11 13 2 7 15 3 3 3 1 11 1 9 0 0 2
10 1 11 11 13 14 0 9 0 9 2
21 1 9 1 0 9 12 2 12 2 12 2 12 15 13 3 0 9 1 10 9 2
11 15 3 13 11 0 1 0 12 0 9 2
22 9 13 12 9 7 11 15 13 9 2 2 11 13 3 16 1 9 10 0 9 2 2
2 11 2
34 1 9 0 9 1 11 13 11 11 1 11 11 12 2 12 2 12 2 12 2 2 12 2 12 2 12 2 12 2 2 12 2 12 2
19 11 13 1 11 1 0 9 3 12 2 12 2 3 15 13 1 0 11 2
29 1 0 9 9 2 15 13 12 9 7 12 9 2 13 11 1 10 9 12 9 2 16 11 0 9 7 12 9 2
12 2 1 9 1 11 13 9 13 1 9 9 2
16 1 10 9 4 13 9 2 7 11 13 3 2 2 13 11 2
26 1 9 3 11 13 1 11 11 2 15 1 12 9 7 12 9 13 12 2 12 2 12 2 12 2 2
2 11 2
27 1 9 9 1 11 13 0 9 0 9 11 11 1 9 11 12 2 12 2 12 2 12 2 12 2 12 2
20 7 15 11 1 9 0 9 13 1 0 11 12 2 12 7 13 15 12 9 2
9 11 9 13 1 0 9 1 11 2
2 0 9
2 11 2
16 12 0 9 13 9 0 9 1 9 1 12 0 9 1 11 2
24 11 11 13 12 9 9 1 0 12 9 7 13 1 0 9 11 11 2 12 2 1 0 9 2
26 0 0 9 13 11 11 2 15 13 1 12 9 9 1 12 7 13 3 12 9 0 9 11 11 12 2
56 0 9 15 13 1 0 9 2 9 0 9 13 11 11 9 12 2 12 1 12 9 9 2 13 11 11 2 12 2 12 2 2 11 11 1 12 9 9 9 12 2 13 11 11 12 2 7 11 11 1 12 9 9 9 12 2
29 0 9 11 11 13 0 9 1 12 9 0 9 9 12 2 12 7 1 0 9 13 3 0 2 12 2 12 2 2
21 1 0 9 13 11 0 9 2 12 2 12 2 7 11 0 2 12 2 12 2 2
15 11 3 13 1 9 1 12 9 9 0 1 12 2 12 2
5 9 11 13 12 9
2 11 2
19 1 0 0 0 9 9 1 0 11 13 11 11 0 0 9 9 12 9 2
5 0 9 1 0 9
16 11 11 2 12 2 13 12 1 12 0 9 9 9 1 9 2
10 9 10 3 0 9 13 0 9 9 2
12 1 9 13 9 10 9 0 9 11 9 11 2
16 1 11 4 15 13 3 3 2 1 10 9 1 11 2 2 2
12 10 10 9 1 11 4 15 13 3 3 0 2
18 13 4 3 1 9 13 0 9 2 16 4 10 10 9 13 3 13 2
5 15 15 13 11 2
9 3 13 9 1 0 9 3 0 2
4 13 15 13 2
23 1 10 9 13 14 12 9 2 7 1 9 15 7 13 3 11 2 9 2 11 7 11 2
6 0 9 15 13 3 2
17 13 9 2 13 15 2 2 7 13 9 2 11 15 13 2 2 2
23 13 15 10 0 9 0 9 2 15 4 3 13 7 3 15 13 2 3 1 15 3 13 2
8 15 13 1 9 12 15 1 12
17 13 2 16 15 9 13 3 1 9 2 13 3 0 7 14 0 2
12 3 4 1 15 13 0 9 1 11 2 2 2
10 2 3 4 15 1 9 1 9 13 2
7 13 4 13 15 3 0 2
11 1 11 11 4 3 13 1 0 0 9 2
16 1 15 13 13 0 9 9 7 9 2 0 9 7 9 9 2
18 10 9 15 14 13 3 1 9 7 15 15 1 10 9 13 1 11 2
16 3 4 15 13 1 15 2 16 9 9 11 13 0 0 9 2
13 13 15 9 13 11 16 9 2 16 10 0 11 2
11 10 9 9 13 14 3 1 15 3 0 2
6 3 15 3 3 13 2
12 15 7 13 11 1 0 9 2 1 0 9 2
7 1 9 13 0 0 9 2
14 13 14 13 9 0 9 1 15 2 3 15 13 13 2
26 11 11 1 9 9 1 9 13 3 11 9 9 2 11 9 9 7 10 0 9 0 9 7 9 7 9
6 15 15 13 1 11 2
1 9
16 1 10 9 1 0 0 9 9 12 13 11 11 1 0 9 2
23 3 3 3 15 13 2 10 0 2 7 0 2 9 15 1 10 9 0 9 9 11 13 2
21 0 7 13 2 16 1 9 1 0 9 15 13 9 0 0 9 7 1 11 9 2
18 9 15 15 9 7 9 13 14 0 9 2 7 7 9 10 9 9 2
34 0 0 9 9 2 0 13 7 7 0 9 7 9 2 15 1 9 13 11 2 11 2 11 2 13 10 2 9 2 1 9 0 9 2
21 15 15 13 1 0 0 9 1 9 1 9 7 9 7 0 9 1 9 3 11 2
9 11 7 0 9 3 13 7 13 2
20 3 0 13 9 2 16 3 15 13 1 11 2 11 7 1 9 7 1 11 2
11 9 3 0 9 13 9 14 10 0 9 2
15 9 3 13 3 0 9 9 2 15 13 3 0 9 9 2
16 1 0 9 11 1 0 9 9 1 9 15 3 13 0 9 2
27 7 16 10 9 7 9 0 9 10 9 13 13 3 0 9 11 11 13 2 15 0 15 13 9 0 9 2
29 9 1 0 0 9 2 10 0 9 13 7 1 9 0 9 0 7 13 15 3 3 2 13 9 1 9 0 9 2
26 9 0 0 0 0 9 13 1 0 9 0 9 2 11 11 2 2 15 7 9 0 9 3 3 13 2
11 9 9 9 3 13 1 9 15 0 9 2
23 0 11 3 13 2 13 7 13 2 3 2 2 16 15 1 15 13 3 3 0 7 0 2
16 9 10 0 0 9 3 13 9 14 0 0 7 3 0 9 2
33 11 3 1 0 9 13 9 9 2 15 16 4 15 1 0 9 7 9 1 9 7 9 1 0 9 9 0 9 13 1 10 9 2
5 0 9 15 3 13
24 0 9 13 1 11 0 2 9 9 9 7 9 7 9 9 10 9 2 9 0 7 0 9 2
15 13 15 1 10 9 1 0 9 2 15 10 9 3 13 2
9 2 10 0 9 2 2 13 0 2
15 2 3 15 13 15 2 15 13 1 0 9 2 2 13 2
32 13 15 1 9 3 3 0 9 9 9 2 15 13 14 1 12 9 2 1 9 13 0 2 2 7 1 9 2 13 9 2 2
25 9 13 0 9 2 3 2 9 2 0 9 2 2 3 13 9 9 0 16 1 9 1 9 12 2
32 9 9 1 0 9 15 13 14 12 2 9 1 0 9 1 9 9 9 7 9 2 7 3 3 13 0 9 1 15 12 9 2
15 16 9 9 4 13 9 1 11 7 9 2 7 0 9 2
13 9 4 13 11 11 1 11 11 7 11 11 11 2
28 0 12 9 1 9 9 9 13 0 9 2 9 2 2 0 9 2 0 9 2 7 0 9 2 14 11 2 2
24 1 9 9 4 13 9 11 2 11 7 11 2 1 9 9 2 9 11 11 7 9 14 3 2
14 9 15 13 9 0 9 2 9 1 11 7 0 9 2
12 1 9 9 13 1 12 9 12 9 0 9 2
7 0 9 16 9 0 0 9
38 0 9 0 9 2 15 1 9 12 13 9 11 11 1 0 9 11 11 2 13 9 9 0 9 1 0 9 0 2 0 7 3 0 0 9 1 11 2
22 0 0 9 2 15 13 11 2 13 3 9 0 0 0 9 11 11 9 9 11 11 2
29 9 13 0 9 11 11 11 1 9 9 12 2 9 9 2 0 9 15 1 9 12 9 1 12 9 13 16 0 2
27 0 9 0 9 13 9 1 9 1 9 11 11 2 12 2 7 9 0 9 11 7 11 0 2 12 2 2
32 1 0 0 9 11 11 11 13 9 0 9 0 9 0 0 0 9 7 0 0 9 2 15 4 13 1 12 1 0 1 9 2
5 9 11 7 9 0
41 9 0 11 16 4 13 9 9 2 1 0 9 2 0 9 1 11 11 2 13 7 13 2 7 1 0 9 1 9 9 9 2 13 0 9 9 3 10 0 9 2
36 1 2 3 0 2 0 9 13 3 9 11 11 2 15 13 9 1 9 10 1 12 9 0 0 9 1 11 7 13 15 0 9 1 0 9 2
37 1 0 9 13 3 0 15 9 16 9 0 9 7 0 9 2 1 9 13 1 9 7 1 9 0 1 9 13 1 9 7 3 15 7 13 9 2
34 3 3 0 9 13 0 9 1 9 1 9 11 11 2 9 11 11 7 11 11 2 10 9 9 2 9 2 15 13 3 0 0 9 2
32 10 3 0 9 15 13 1 11 9 12 2 15 9 13 9 9 7 9 2 1 15 15 13 7 13 0 0 0 9 7 9 2
39 1 9 3 0 2 9 9 2 13 9 11 11 2 9 1 11 2 1 15 13 10 9 0 9 2 0 9 9 9 2 15 13 1 0 9 7 0 9 2
21 0 9 2 0 0 9 2 0 9 7 3 7 9 11 11 13 9 9 11 11 2
23 11 15 3 3 13 1 0 0 9 0 1 9 2 0 1 0 9 2 2 0 1 9 2
19 15 9 13 10 0 9 9 1 3 0 2 0 9 2 2 0 9 2 2
21 13 15 3 7 14 1 9 1 10 9 1 0 0 9 9 9 2 11 11 2 2
24 1 11 2 15 13 9 0 9 2 7 12 0 0 9 15 3 13 7 11 1 9 9 9 2
16 0 11 15 13 13 7 12 3 0 9 0 0 9 11 11 2
27 10 0 0 9 0 9 2 0 9 2 13 0 9 0 0 9 2 15 1 0 9 0 11 13 0 9 2
31 0 0 9 13 14 0 9 2 7 7 0 0 9 0 0 9 9 7 0 9 2 0 9 2 0 9 7 3 0 9 2
29 3 3 13 0 9 0 9 2 9 0 0 9 11 11 2 11 2 0 9 2 7 0 9 11 11 2 9 2 2
26 11 11 11 2 3 2 9 0 9 9 11 2 3 13 1 10 0 9 2 0 9 2 0 9 9 2
30 13 1 14 3 0 9 2 1 15 15 1 9 1 0 9 9 13 9 0 9 2 0 9 7 9 9 1 10 9 2
15 1 9 3 15 1 9 9 0 9 13 7 0 0 9 2
12 0 9 9 9 11 11 13 9 3 16 0 2
14 3 15 1 15 13 7 3 3 1 0 9 0 9 2
5 9 3 13 15 0
32 1 0 9 15 9 13 1 9 2 13 9 1 9 11 3 4 13 0 9 9 1 0 9 1 9 12 0 9 9 0 9 2
10 13 0 9 9 2 7 3 10 9 2
18 11 15 13 1 9 9 9 2 9 2 2 15 13 12 2 9 12 2
31 11 11 2 11 7 11 2 16 15 1 10 9 13 13 12 2 9 2 13 15 0 9 0 1 10 9 13 2 3 13 2
8 15 13 2 16 4 13 9 2
29 10 9 2 3 1 0 0 9 10 9 2 3 13 1 0 9 9 10 9 2 16 11 11 2 9 2 9 3 2
13 1 0 9 15 13 3 13 9 9 7 0 9 2
24 0 9 13 13 7 1 9 1 12 2 9 2 1 3 0 9 2 11 2 11 0 2 2 2
34 11 11 2 0 7 0 9 2 9 2 12 2 13 15 2 16 4 0 9 9 13 0 9 1 0 9 9 7 9 9 1 0 9 2
17 9 2 13 0 9 2 4 13 13 10 9 3 7 1 0 9 2
22 11 11 2 0 11 2 0 9 1 9 1 9 9 1 0 9 15 13 14 3 13 2
10 3 0 13 0 9 2 15 9 13 2
20 3 3 13 0 2 16 15 4 1 0 9 0 2 11 3 13 2 13 0 2
22 1 9 0 9 4 9 13 7 3 0 9 2 7 10 9 7 9 9 3 0 9 2
28 9 0 9 15 14 0 9 1 0 9 13 7 16 14 2 3 1 9 9 2 9 12 2 1 9 9 9 2
9 0 9 9 13 1 10 9 13 2
25 11 11 2 0 11 2 13 2 16 0 9 13 1 9 9 7 0 9 3 0 2 16 9 0 2
13 11 9 2 11 9 2 0 9 13 0 9 9 2
15 11 11 2 0 11 2 9 1 0 9 4 13 0 9 2
25 13 15 13 2 16 9 1 15 15 13 1 0 9 9 7 9 2 7 7 15 4 13 3 10 2
10 13 10 9 2 16 4 13 0 9 2
25 11 11 2 0 9 2 0 9 13 1 9 9 0 9 7 0 9 1 9 0 1 9 0 9 2
14 13 9 9 1 14 12 9 2 9 2 9 7 9 2
16 11 11 2 0 11 2 3 0 9 9 1 9 1 0 9 2
8 0 0 9 1 9 0 9 2
42 11 11 2 0 11 2 9 1 9 1 0 9 4 1 0 9 13 9 0 9 0 9 1 0 9 12 5 1 12 9 2 7 15 14 1 0 9 7 9 0 9 2
22 3 15 13 0 9 9 2 7 1 9 2 15 4 13 9 1 0 9 2 3 13 2
15 11 11 2 11 11 2 15 4 13 1 9 9 0 9 2
27 1 0 9 15 7 13 2 16 3 0 0 9 13 3 3 0 9 7 13 15 14 1 9 0 0 9 2
30 11 11 2 11 9 11 2 13 15 13 2 16 3 0 9 15 9 13 1 0 0 9 2 15 13 1 9 10 9 2
10 1 9 13 7 9 2 15 4 13 2
14 1 9 9 7 9 13 2 7 15 13 9 1 9 2
3 0 11 2
22 9 15 1 0 9 1 0 0 9 13 1 12 0 9 2 15 13 3 1 9 12 2
15 9 9 1 9 15 1 10 9 13 3 1 0 0 9 2
18 9 13 2 16 9 0 9 13 0 9 2 15 13 0 9 0 9 2
7 9 13 3 2 13 9 2
7 0 9 13 1 0 11 2
23 13 13 2 16 9 9 13 1 9 2 16 0 9 13 0 13 9 9 1 0 0 9 2
1 3
21 0 0 9 7 0 9 3 13 0 0 9 1 0 9 0 9 11 1 0 9 2
18 9 13 3 0 9 7 1 9 13 0 9 2 13 9 0 9 11 2
19 1 9 1 0 9 7 0 9 1 0 11 13 1 9 1 9 12 9 2
21 13 15 3 0 9 1 15 2 16 13 1 0 9 1 12 9 0 9 1 9 2
33 12 9 2 15 15 13 13 0 9 1 0 9 3 0 9 11 2 3 13 0 2 0 9 9 2 0 9 3 12 9 1 9 2
8 9 3 9 13 7 13 13 2
18 9 9 9 13 1 3 16 12 9 2 1 15 9 7 9 13 9 2
23 12 0 7 3 12 0 15 13 9 2 1 15 13 1 0 9 1 9 11 1 9 11 2
27 1 9 9 13 0 0 0 9 2 11 2 2 15 13 2 16 9 9 1 10 0 9 0 1 11 13 2
39 9 11 11 11 13 9 0 9 11 11 2 16 4 15 1 15 13 12 2 9 1 11 1 9 1 12 2 9 9 0 9 1 0 11 1 0 0 9 2
12 1 9 11 15 1 9 13 0 0 0 9 2
19 10 0 9 13 2 16 0 9 7 1 0 0 0 2 0 9 3 13 2
8 11 7 11 15 3 13 9 9
6 11 2 11 2 11 2
31 11 2 0 9 9 1 9 11 2 13 0 9 1 11 2 16 13 1 0 9 2 16 13 1 9 1 9 0 0 9 2
33 13 3 1 0 9 11 2 15 13 2 16 4 2 14 0 9 1 0 9 13 0 9 0 9 2 3 10 9 1 0 9 13 2
21 9 11 11 11 15 1 11 13 1 0 9 9 11 11 1 9 1 9 0 9 2
18 11 15 13 1 9 1 9 1 15 2 16 2 4 13 0 9 2 2
21 1 3 16 12 9 7 3 11 13 14 12 11 1 9 11 13 1 9 1 11 2
23 0 9 3 3 13 9 0 9 1 9 11 13 9 10 9 9 1 0 9 11 1 11 2
18 0 9 7 9 3 3 13 1 10 9 9 0 9 11 1 9 11 2
10 1 9 4 12 9 13 7 15 13 2
21 1 9 0 11 3 13 14 12 9 2 15 13 1 9 12 0 9 7 12 9 2
18 9 13 9 1 0 9 11 2 1 15 4 13 9 11 7 12 9 2
5 0 9 0 0 9
15 9 11 11 1 9 15 13 9 0 9 1 9 1 0 9
13 9 1 9 13 10 0 9 0 9 11 11 11 2
11 1 0 9 0 0 9 13 1 0 9 2
29 16 10 9 13 12 9 3 2 13 10 0 9 0 9 7 0 9 0 9 1 0 0 9 13 1 12 9 3 2
40 0 12 9 0 2 1 11 3 0 2 9 11 11 2 15 15 13 1 9 13 2 16 4 13 1 9 0 9 13 1 9 9 2 13 1 0 9 0 9 2
12 10 9 15 13 3 1 9 1 9 0 9 2
47 1 12 9 15 1 9 3 13 2 16 10 9 13 9 0 9 11 11 11 11 2 12 2 0 0 9 9 2 7 9 9 11 11 2 12 2 2 15 13 0 11 7 0 9 0 9 2
9 0 9 9 3 1 9 13 11 2
19 1 0 9 12 0 9 13 14 3 13 2 15 1 15 4 9 13 3 2
26 2 4 2 14 13 2 13 4 13 1 9 2 15 13 11 2 2 13 15 11 1 9 0 9 9 2
10 11 1 15 13 0 9 7 9 9 2
11 1 11 13 0 9 2 1 11 9 9 2
13 3 15 4 4 13 13 1 9 1 11 9 0 2
37 9 3 13 14 0 0 9 2 7 7 9 0 9 1 9 9 1 9 2 15 4 2 16 4 13 14 1 9 2 13 4 13 3 3 1 9 2
26 9 9 13 0 9 0 9 0 7 0 9 11 11 1 9 2 16 9 0 0 9 13 9 0 9 2
28 9 13 1 15 2 16 0 0 9 4 1 9 0 13 0 9 7 13 0 2 0 9 2 1 10 0 9 2
26 3 4 15 13 3 13 2 16 1 12 0 9 2 3 0 9 11 13 0 9 2 13 0 9 9 2
32 10 9 13 7 0 9 0 9 2 1 15 15 12 9 9 13 3 1 9 2 16 1 0 9 4 3 13 0 12 9 9 2
23 10 9 3 13 13 7 9 2 16 15 11 13 13 1 0 9 9 1 0 0 0 9 2
32 9 11 11 2 15 9 13 1 9 12 2 12 9 3 2 16 13 1 0 9 2 13 9 2 3 11 13 0 7 0 9 2
29 7 12 1 9 1 9 2 0 9 11 11 7 0 9 11 11 2 13 0 9 9 2 1 15 15 13 13 11 2
32 10 9 4 1 11 13 1 0 2 9 2 7 1 9 9 2 15 13 1 2 9 9 2 1 9 12 2 15 13 0 9 2
26 16 15 1 0 9 13 0 9 9 15 1 12 0 2 1 9 1 3 0 11 13 0 9 16 0 2
6 11 2 9 1 9 9
2 11 2
21 3 13 1 11 13 0 9 1 9 9 9 9 0 9 9 2 15 13 9 9 2
23 0 13 9 7 9 3 3 13 0 9 2 9 0 9 0 10 0 9 13 3 1 11 2
31 9 0 11 2 11 11 13 9 1 9 12 9 1 10 2 16 10 9 4 1 9 12 13 0 9 1 9 1 0 9 2
14 1 12 9 9 0 1 11 13 12 9 1 12 9 2
6 1 11 13 13 1 11
2 11 2
25 0 9 9 11 1 11 3 13 9 0 9 1 0 0 9 1 0 0 9 2 11 2 11 11 2
31 13 3 1 9 9 11 11 1 0 9 11 1 9 9 1 11 2 0 9 9 11 7 0 0 0 9 1 9 1 11 2
41 1 1 0 9 15 9 0 11 2 1 15 13 3 9 2 13 1 0 9 0 9 7 1 9 11 15 13 1 0 0 9 7 13 15 1 9 1 9 0 9 2
10 13 3 10 9 9 0 9 7 9 2
4 9 15 13 11
2 11 2
16 0 0 9 11 13 3 9 1 0 0 9 11 3 1 11 2
23 1 11 13 9 9 2 1 10 9 13 9 0 11 9 11 11 2 3 0 16 0 9 2
15 1 0 9 13 3 9 1 9 3 12 1 12 0 9 2
17 0 9 9 13 11 2 0 9 0 0 0 9 0 9 11 11 2
13 9 13 3 1 0 9 14 12 9 1 0 9 2
10 10 9 3 13 1 2 12 9 2 2
45 11 2 15 15 13 3 1 12 9 1 0 9 11 7 3 13 0 9 1 2 15 0 9 0 9 2 2 13 9 0 1 9 2 1 15 11 13 1 9 0 9 1 9 12 2
19 13 9 2 16 11 4 13 1 0 11 2 1 11 2 7 7 1 11 2
16 1 12 9 13 1 9 11 2 1 0 13 1 15 3 11 2
21 11 13 2 16 13 9 13 1 15 9 2 15 13 14 0 7 13 15 1 9 2
23 11 7 9 11 11 2 12 0 9 0 11 2 1 9 13 0 9 1 9 0 9 11 2
10 13 3 9 1 0 9 9 1 9 2
18 11 13 9 15 12 0 9 1 0 9 2 15 1 9 13 9 11 2
16 1 0 9 13 13 1 10 9 2 0 9 2 7 0 9 2
11 0 9 13 9 0 0 9 1 15 11 2
30 12 1 9 9 13 9 11 2 16 0 0 9 4 3 13 13 13 1 9 9 2 16 15 14 13 0 9 0 9 2
22 15 15 3 13 0 9 2 15 1 0 9 13 7 13 15 3 9 1 0 12 11 2
23 1 0 9 3 13 1 9 9 9 1 9 2 3 11 9 11 7 11 11 11 13 11 2
7 11 13 2 16 15 13 9
2 11 2
40 1 9 2 16 4 13 0 15 13 9 2 13 9 11 0 0 9 11 11 2 2 13 1 0 9 7 15 13 3 0 2 16 1 15 13 0 7 0 9 2
13 13 7 9 2 16 1 15 4 12 9 9 13 2
6 7 13 15 15 2 2
19 13 2 16 16 4 1 15 13 2 13 4 15 3 3 2 0 9 2 2
21 2 13 1 15 3 16 10 9 9 7 13 4 1 9 2 16 9 15 13 2 2
10 1 0 11 13 1 15 0 10 9 2
18 2 3 0 9 2 2 13 2 16 2 9 3 13 1 0 9 2 2
13 1 10 9 13 9 9 13 2 3 0 9 2 2
27 11 2 9 9 0 9 2 0 9 1 0 9 1 0 9 2 4 3 13 1 12 1 9 1 0 9 2
31 16 3 13 9 1 11 7 9 9 9 1 9 11 11 2 13 9 2 16 4 15 13 9 12 2 9 0 1 0 11 2
5 11 13 1 9 9
2 11 2
23 0 9 11 11 3 13 2 16 13 0 9 1 9 0 9 2 16 4 3 13 0 9 2
26 1 0 9 11 9 13 2 16 2 4 2 14 10 9 1 9 13 2 4 3 13 13 0 9 2 2
20 13 3 2 2 16 15 13 9 11 0 2 4 13 3 13 7 15 13 2 2
25 11 13 15 2 16 9 13 13 2 16 15 1 9 13 1 0 9 1 9 9 2 9 7 9 2
10 10 9 4 13 1 9 9 1 9 2
12 11 3 13 0 9 1 9 9 9 7 9 2
15 15 15 1 9 13 10 9 2 1 15 15 7 9 13 2
22 13 15 2 16 0 9 2 3 13 0 9 0 9 2 13 11 0 9 12 2 9 2
5 11 2 11 7 11
25 0 9 9 9 1 9 4 1 9 9 3 13 16 10 0 0 0 9 1 9 1 9 0 9 2
41 16 1 11 13 0 9 2 16 11 15 1 15 13 1 9 10 0 9 2 13 3 9 3 0 0 9 16 0 0 9 14 16 9 11 2 7 3 9 0 9 2
60 9 2 15 0 9 9 0 0 9 13 11 7 3 0 10 9 2 13 0 2 13 3 3 3 2 3 7 3 2 1 0 9 7 0 9 2 15 14 3 3 3 13 0 10 9 2 13 10 9 2 15 1 9 9 13 0 9 7 9 2
23 13 10 9 1 11 7 1 9 2 15 3 3 13 9 7 9 3 1 10 3 0 9 2
33 13 15 9 0 3 3 2 16 2 1 15 15 3 15 13 2 0 0 9 3 13 1 12 2 7 1 12 9 2 1 9 12 2
29 9 9 7 10 0 9 13 0 9 2 7 1 9 15 13 3 0 2 9 11 7 2 9 2 0 9 1 11 2
16 0 13 9 9 0 0 9 2 7 12 7 3 13 0 9 2
20 11 10 0 9 0 9 3 13 2 3 16 10 9 7 9 13 9 0 11 2
24 7 11 7 9 15 1 10 0 9 13 3 13 2 3 7 3 9 9 2 16 10 0 9 2
20 1 10 2 3 16 3 2 0 9 13 13 15 3 2 13 1 15 14 13 2
9 10 0 9 13 13 7 13 15 2
28 9 9 15 13 1 9 1 11 2 1 10 9 2 1 15 15 0 9 7 0 9 1 10 0 9 3 13 2
18 13 15 3 2 3 7 3 2 9 2 15 3 13 9 7 0 9 2
46 13 3 15 2 15 3 3 13 15 0 9 1 11 2 9 13 9 7 2 16 13 2 7 3 13 15 7 13 15 15 13 0 2 3 0 7 3 7 0 4 13 13 9 15 13 2
16 0 0 9 3 13 13 15 0 16 2 9 2 9 9 0 2
36 3 13 3 3 0 3 3 13 9 1 12 9 2 0 7 0 2 3 14 13 13 2 16 15 13 11 2 15 13 9 9 7 9 1 9 2
74 15 2 16 4 15 3 1 9 10 9 13 3 2 3 1 9 1 9 0 9 10 9 2 15 15 13 9 3 0 10 0 9 2 15 1 15 13 2 13 0 9 0 9 2 15 4 13 10 9 1 0 14 0 2 0 9 2 2 15 13 2 9 9 1 0 9 9 2 2 11 2 11 2 2
39 7 15 2 9 7 10 3 1 9 0 7 3 7 0 9 2 3 7 9 9 0 9 2 13 9 2 15 13 2 3 3 1 0 9 2 13 7 13 2
19 15 1 15 7 13 13 7 3 3 13 2 16 4 15 13 13 15 0 2
10 15 13 0 9 7 1 0 0 9 2
9 1 15 15 13 9 2 7 9 2
34 13 4 15 13 1 9 16 1 15 0 7 1 11 3 0 9 11 2 7 7 0 0 9 2 0 3 9 15 1 10 9 9 13 2
34 15 15 13 0 13 1 15 2 16 4 15 13 2 15 13 2 7 1 10 0 9 2 16 4 15 7 15 13 2 15 13 0 9 2
35 13 7 14 1 0 9 2 13 1 10 9 1 0 10 9 2 15 15 3 2 1 0 9 0 0 9 2 0 9 0 9 2 3 13 2
14 0 2 0 9 13 12 1 0 9 1 9 0 11 2
19 4 2 14 10 9 13 2 13 4 3 4 13 2 16 4 13 0 9 2
18 13 3 15 9 1 15 2 16 4 1 10 0 9 11 13 0 9 2
42 13 4 14 3 2 7 1 9 2 13 2 16 13 13 0 2 7 15 15 2 16 13 2 16 4 15 0 7 0 9 0 2 1 15 0 0 9 13 0 0 9 2
77 9 11 15 13 3 3 2 13 15 15 7 13 9 10 2 13 3 7 3 13 1 9 9 1 0 2 9 0 1 15 2 15 1 15 13 2 2 3 14 9 11 2 11 2 2 1 9 0 9 0 15 10 0 9 0 1 9 2 7 1 9 2 7 0 3 1 15 15 2 1 0 9 7 9 2 13 2
32 1 2 0 2 11 9 7 9 15 13 13 11 2 9 10 0 9 2 14 3 15 2 16 15 11 13 2 7 0 0 9 2
19 13 15 15 0 7 13 1 15 1 15 0 9 10 9 7 10 0 9 2
14 16 15 15 13 2 13 1 15 9 1 0 9 3 2
2 0 9
25 10 0 9 15 3 13 13 12 0 9 2 7 16 2 7 15 13 2 9 0 2 0 2 9 2
29 13 13 12 9 9 1 0 9 2 1 0 9 9 2 10 13 11 11 2 7 1 9 2 15 15 3 13 13 2
26 9 13 2 15 4 15 3 13 2 7 16 13 15 1 15 1 9 2 13 0 2 16 15 13 15 2
23 1 0 9 15 15 13 12 7 0 9 1 15 13 2 13 2 14 15 3 2 7 3 2
21 13 2 14 9 2 1 15 15 1 15 13 1 15 9 2 3 13 15 3 3 2
34 7 16 0 0 9 2 15 15 13 2 13 3 7 16 1 15 3 13 9 2 1 15 15 9 13 2 13 0 9 3 14 3 10 2
14 0 0 9 1 9 13 9 2 13 1 9 9 2 2
26 13 3 1 9 9 2 7 16 9 2 9 9 2 3 13 2 7 3 13 2 16 15 10 9 13 2
41 13 9 7 9 0 9 2 10 9 13 9 9 3 0 2 9 3 0 2 9 1 0 9 2 3 14 3 9 0 2 0 2 2 7 3 9 2 15 13 0 2
11 7 15 3 3 2 7 7 3 1 9 2
23 13 15 10 3 0 9 13 0 7 13 0 9 1 15 1 15 2 13 13 9 9 0 2
22 15 15 9 0 13 2 7 13 15 0 2 16 15 15 13 3 3 0 7 10 9 2
35 9 13 10 9 13 9 2 7 15 14 1 9 1 9 2 2 7 13 15 13 3 16 1 9 1 9 15 2 15 1 10 9 3 13 2
11 13 15 13 3 2 16 15 13 1 9 2
31 3 2 0 9 9 1 12 2 9 12 7 3 9 0 9 1 12 2 9 12 10 9 15 2 15 15 13 13 2 13 2
8 3 13 1 9 13 12 9 2
14 0 1 15 13 2 0 9 3 12 5 0 9 2 2
23 13 15 0 2 16 13 15 2 15 9 13 7 13 2 1 15 13 2 3 2 15 13 2
53 13 3 15 2 15 4 13 0 9 3 12 5 9 2 7 2 3 13 9 2 12 5 1 9 2 2 16 15 1 0 9 4 13 1 0 9 9 1 9 12 5 0 9 2 16 15 1 0 9 3 12 5 2
16 3 15 13 0 2 3 1 15 4 13 2 13 9 2 9 2
10 13 15 0 2 7 3 0 9 9 2
6 0 9 13 3 15 2
36 16 15 13 12 5 7 12 5 1 9 7 1 0 9 13 9 0 9 2 15 13 1 0 9 7 15 15 13 1 9 1 0 9 3 13 2
24 0 9 13 2 13 9 0 9 9 1 9 1 12 9 2 2 16 9 12 4 3 15 13 2
32 1 0 4 13 13 15 2 16 13 13 9 0 9 0 2 16 13 13 1 9 7 16 1 15 13 13 3 14 1 9 12 2
10 13 3 9 0 9 1 15 1 15 2
63 15 14 15 1 0 9 13 2 7 15 4 15 7 13 13 0 12 0 9 7 3 2 12 0 9 2 16 13 15 1 15 3 3 3 0 9 2 16 4 15 1 15 13 0 9 2 7 3 0 9 2 3 2 9 9 2 15 1 15 4 13 2 2
14 1 0 4 13 13 2 16 13 1 12 9 13 0 2
21 9 13 1 12 9 1 9 2 1 12 1 12 9 2 7 1 12 9 1 9 2
36 1 9 0 13 1 9 1 9 9 2 3 1 12 9 2 1 9 1 9 1 12 2 1 12 9 2 14 1 12 9 2 1 12 9 2 2
43 1 0 13 13 2 16 15 0 9 7 1 10 9 13 2 7 13 15 13 2 16 1 0 9 1 15 13 13 10 9 3 3 9 13 7 3 9 13 13 1 0 9 2
31 14 4 1 10 9 1 9 13 0 9 2 7 14 15 4 3 13 16 0 9 9 7 16 0 9 9 1 10 0 9 2
19 0 9 13 2 2 16 4 9 0 1 0 9 4 13 1 0 9 2 2
33 13 2 16 15 15 1 15 13 1 9 7 16 9 13 3 1 15 2 1 3 0 2 7 0 2 0 9 15 13 1 9 13 2
13 13 0 9 2 16 13 0 0 9 12 0 9 2
66 7 13 3 0 9 15 2 15 15 2 1 0 9 0 9 2 13 2 7 15 15 3 13 0 9 9 2 15 13 3 0 9 2 1 9 13 2 7 13 0 9 0 9 9 9 2 1 0 9 2 7 1 15 9 9 1 0 9 2 3 7 3 2 13 13 2
19 15 3 13 9 0 7 13 9 2 16 10 9 0 9 10 9 13 3 2
24 3 2 13 1 9 9 2 7 1 9 1 0 9 2 1 15 2 13 2 13 9 0 9 2
18 3 10 0 9 13 0 9 2 7 7 15 13 2 16 13 10 9 2
4 9 13 3 0
1 9
16 1 0 0 9 9 13 0 9 10 9 7 0 9 1 9 2
30 0 9 9 7 0 9 3 10 9 13 7 1 9 9 1 9 2 3 3 13 7 13 0 9 2 13 1 0 9 2
13 13 1 15 9 11 9 0 9 1 9 0 9 2
21 0 9 2 16 0 9 13 3 0 9 1 9 2 13 2 13 15 2 3 0 2
30 1 0 13 9 9 2 15 13 0 9 0 9 9 2 0 9 1 9 2 9 1 9 2 0 9 7 9 1 9 2
18 3 3 9 13 9 0 9 7 9 2 3 9 2 9 7 9 9 2
19 3 15 3 13 1 0 7 0 9 2 3 15 3 13 0 9 1 9 2
11 0 9 1 0 15 13 0 9 1 9 2
15 15 13 3 3 7 3 13 13 9 2 9 9 7 9 2
11 9 13 3 3 0 9 1 9 7 9 2
19 1 0 9 1 9 13 9 2 9 2 0 9 7 9 1 9 7 9 2
17 0 9 9 13 0 9 1 0 9 2 10 9 4 9 3 13 2
15 9 3 1 0 9 13 9 2 3 9 9 7 9 9 2
13 0 13 2 15 1 0 9 3 13 9 0 9 2
17 1 9 13 1 12 9 2 1 0 9 7 1 0 9 1 9 2
6 3 9 13 1 9 2
21 15 13 0 2 15 0 13 9 14 1 9 1 9 2 7 7 1 9 1 9 2
14 9 7 13 2 16 7 3 13 9 13 0 0 9 2
9 1 0 2 7 0 9 13 9 2
9 12 0 13 9 1 12 9 9 2
29 9 3 1 0 12 9 9 9 0 9 13 7 3 2 3 13 9 2 0 0 9 4 15 13 1 9 3 13 2
17 7 0 9 7 3 13 9 2 15 13 1 9 0 1 0 9 2
14 0 9 4 1 9 13 3 2 9 4 3 13 9 2
10 12 1 0 9 13 0 15 0 9 2
21 16 1 11 13 9 9 7 9 1 9 12 2 11 1 10 9 13 3 0 9 2
19 0 9 0 13 7 1 15 7 9 13 2 16 15 13 9 9 0 9 2
32 0 9 1 0 9 13 2 0 2 9 9 2 0 9 1 9 7 3 0 9 2 15 3 10 9 0 9 13 1 9 9 2
16 13 7 9 2 16 1 9 0 0 9 13 1 0 0 9 2
23 9 2 3 15 4 13 9 13 3 9 7 9 2 15 3 13 1 9 16 1 0 9 2
18 0 15 13 2 16 9 13 3 13 2 9 15 13 13 0 0 9 2
13 3 14 3 3 13 10 9 7 13 7 1 9 2
2 10 9
1 9
19 9 0 9 11 11 15 13 13 2 16 9 13 1 9 0 9 0 9 2
15 16 9 13 2 16 0 9 11 12 4 13 1 9 13 2
37 1 9 2 15 13 9 9 0 9 1 0 9 2 4 15 13 13 2 16 13 9 7 13 15 1 3 0 9 2 16 1 9 9 13 10 9 2
21 9 2 9 2 4 3 13 9 2 3 15 0 9 13 1 9 0 1 9 0 2
24 15 9 0 9 7 9 7 13 7 7 3 13 1 0 9 2 0 9 1 15 13 7 9 2
12 9 9 13 3 9 13 10 9 1 0 9 2
4 13 1 9 2
21 9 9 2 3 3 3 1 0 9 2 13 13 0 9 2 1 15 13 0 9 2
23 0 0 9 13 2 16 1 9 9 9 9 11 4 9 3 13 13 1 9 9 11 12 2
29 9 4 13 9 12 0 9 1 3 0 9 2 9 0 2 9 2 1 9 0 9 0 9 9 1 9 0 9 2
18 9 9 11 13 7 13 1 3 0 0 9 2 15 15 13 10 9 2
41 0 9 9 3 1 0 9 9 1 9 11 13 3 1 15 2 16 0 9 15 1 9 13 16 0 2 10 0 9 15 13 1 9 2 15 13 14 0 9 9 2
9 0 9 3 4 13 1 9 0 2
27 16 4 11 13 9 14 12 2 3 15 2 15 13 3 0 9 2 13 4 10 2 9 2 3 1 15 2
17 0 0 9 0 9 4 3 3 15 13 13 7 1 9 0 9 2
9 3 2 13 15 12 1 0 9 2
17 13 7 0 7 7 13 2 16 0 9 3 13 13 0 0 9 2
23 3 11 1 10 0 9 14 3 3 3 13 2 16 15 13 3 0 3 1 9 0 9 2
15 0 0 9 3 1 9 9 9 1 9 13 3 12 9 2
9 16 1 9 4 13 13 3 3 2
5 9 7 3 13 2
3 9 1 15
3 13 10 9
5 14 2 0 9 2
2 11 2
28 9 0 1 0 9 13 1 9 3 1 12 1 0 9 11 1 11 12 0 11 13 10 12 0 9 1 11 2
18 9 2 15 4 13 1 0 9 1 9 3 0 9 2 1 9 13 2
12 9 1 9 1 9 12 9 13 0 0 9 2
22 9 1 9 1 9 9 9 13 7 3 13 13 1 0 9 9 1 9 1 9 9 2
5 0 9 13 0 9
4 11 1 11 2
35 0 9 3 13 1 9 1 9 0 9 0 9 3 11 1 11 1 9 9 9 9 11 11 0 9 2 3 0 2 15 13 1 0 9 2
9 0 9 13 9 9 0 9 11 2
11 1 9 9 4 1 9 13 9 0 9 2
10 0 9 13 2 16 9 13 0 9 2
38 9 15 13 1 15 9 2 15 15 1 9 1 12 1 12 9 12 2 9 13 1 9 1 0 9 11 1 9 11 7 0 9 2 16 4 13 9 2
6 1 0 9 13 9 9
5 14 2 0 9 2
2 11 2
41 1 9 9 11 11 11 13 9 9 0 9 0 2 0 7 0 9 1 11 9 1 9 0 1 0 9 7 3 13 9 1 9 9 2 16 15 4 13 10 9 2
30 9 9 9 13 3 1 15 9 9 7 10 9 1 9 2 16 15 13 0 2 16 13 1 9 2 3 3 0 2 2
37 11 13 2 16 4 0 0 9 2 15 13 1 11 0 1 9 0 9 2 13 9 10 9 2 16 2 13 3 13 2 16 15 1 9 13 2 2
33 1 9 0 0 9 11 11 11 13 9 9 2 0 9 2 15 13 13 9 2 7 0 9 4 13 9 1 10 9 1 0 9 2
35 9 0 0 9 11 11 1 0 0 9 13 2 16 2 16 15 15 13 2 16 9 13 13 7 1 11 2 3 13 2 1 15 13 2 2
8 0 9 11 13 1 9 9 9
2 11 2
20 0 0 9 13 2 1 0 9 2 1 9 9 1 9 9 7 9 0 9 2
11 3 13 9 0 9 2 15 13 1 0 2
25 13 15 15 1 9 0 9 11 2 0 1 9 1 11 1 9 0 9 11 0 9 1 9 9 2
28 9 11 11 11 13 2 16 2 0 9 13 1 0 7 0 15 3 1 9 0 9 1 9 3 3 13 2 2
20 13 2 16 1 1 0 9 11 13 0 9 11 0 9 1 9 9 1 0 2
5 11 13 0 0 9
3 1 0 9
3 0 11 2
31 0 9 0 9 0 0 9 2 15 13 10 9 11 11 2 13 1 9 0 9 11 1 9 1 0 11 1 0 2 11 2
29 3 13 9 9 11 11 2 0 9 9 4 13 4 13 1 0 9 11 3 2 16 13 2 0 9 2 9 9 2
14 0 0 9 9 13 0 9 13 1 9 12 2 9 2
9 9 13 1 11 3 16 10 0 9
3 0 11 2
16 1 0 9 0 0 9 13 11 9 0 0 9 1 0 9 2
12 13 15 1 9 0 9 9 10 9 11 11 2
21 3 13 2 1 9 1 0 0 9 2 9 2 1 10 9 1 0 9 13 9 2
44 0 9 11 13 9 9 0 7 0 9 2 15 13 9 9 11 11 11 1 15 2 16 9 3 13 0 9 2 7 13 0 9 1 0 2 13 0 9 9 0 9 11 11 2
16 11 13 2 16 9 0 9 13 1 11 3 16 10 0 9 2
25 2 14 2 9 13 1 15 0 9 2 13 7 0 2 15 15 13 7 15 15 13 2 2 13 2
31 1 10 0 9 0 9 13 3 1 9 9 2 9 0 9 9 2 9 0 9 2 9 0 9 7 9 9 1 0 9 2
7 0 9 13 1 3 0 9
2 11 2
41 16 9 9 1 0 9 1 9 2 9 2 0 9 7 9 2 13 3 0 9 0 9 2 11 2 11 11 12 2 0 9 10 9 2 15 3 13 1 0 11 2
27 12 9 9 1 12 0 9 13 3 9 2 15 15 13 11 11 2 7 0 9 9 2 15 13 11 11 2
10 1 0 0 9 13 3 13 0 9 2
21 9 15 1 10 9 1 11 13 7 11 11 2 13 3 4 11 11 7 11 11 2
11 15 1 9 13 2 16 13 1 0 9 2
12 0 0 9 13 9 1 9 3 0 9 9 2
27 10 9 15 1 0 9 13 14 0 9 2 7 13 7 9 0 0 9 2 0 0 9 2 9 7 9 2
27 1 10 0 9 1 9 11 13 2 16 1 0 9 13 0 9 3 2 2 3 13 16 0 0 9 2 2
18 9 9 1 9 1 9 7 13 2 13 15 3 1 0 0 9 2 2
24 0 9 13 2 16 1 9 9 15 10 0 9 13 1 0 12 9 2 3 1 12 9 2 2
27 2 16 15 15 15 13 2 3 13 13 0 9 1 3 0 9 16 15 0 2 2 13 11 1 0 9 2
7 11 2 9 1 9 15 13
3 1 0 9
2 11 2
14 1 0 13 9 9 1 9 0 9 9 11 11 11 2
12 13 2 16 0 9 13 9 1 9 0 9 2
31 2 3 15 13 7 9 0 9 9 1 9 11 2 16 1 0 0 9 4 13 9 1 0 9 0 9 2 2 13 9 2
16 9 11 11 13 2 16 11 10 0 9 13 1 0 9 9 2
17 2 13 7 1 9 15 7 9 2 16 4 13 1 0 0 9 2
11 1 9 0 9 15 15 13 2 2 13 2
24 2 13 4 0 2 16 4 1 10 9 13 0 2 7 1 0 9 0 9 2 2 13 11 2
7 11 15 13 1 9 0 9
2 11 2
24 1 0 0 9 11 1 9 1 9 1 11 13 1 9 9 9 11 9 11 11 2 11 2 2
27 13 2 16 9 3 13 9 9 1 0 9 2 16 13 1 9 0 7 0 2 3 7 3 1 9 0 2
32 9 13 1 9 9 13 2 1 10 9 4 1 9 1 9 1 0 9 13 1 9 0 9 2 15 1 0 9 13 9 9 2
39 3 13 13 2 10 9 13 9 1 0 0 9 9 11 1 10 9 7 1 10 9 9 1 9 1 9 13 1 9 0 9 7 3 1 0 9 0 9 2
43 11 4 0 13 9 7 1 9 2 16 10 9 13 1 9 9 0 9 11 2 15 4 1 1 10 9 1 11 13 13 1 0 9 10 9 2 15 4 13 13 9 11 2
5 9 1 9 9 9
11 9 2 9 7 9 0 9 13 1 0 9
2 11 2
23 1 9 9 1 12 9 2 15 13 0 9 9 1 0 9 2 9 0 0 9 15 13 2
28 13 7 13 2 16 9 13 9 1 15 2 16 4 3 9 1 9 2 0 9 7 9 13 14 9 3 0 2
21 9 9 15 7 13 9 2 0 15 9 2 9 2 0 9 7 3 9 1 9 2
28 9 7 0 9 1 9 1 9 1 12 9 4 1 9 9 13 13 14 9 2 10 9 13 12 9 0 9 2
15 2 0 9 1 12 0 9 1 0 9 13 12 9 2 2
24 0 9 13 13 1 9 1 9 2 15 4 13 4 13 3 9 1 9 1 12 9 0 9 2
20 1 9 9 7 0 9 4 13 4 10 12 9 13 15 1 9 1 9 9 2
18 10 9 13 0 9 2 9 1 0 0 9 7 0 9 9 1 9 2
33 2 16 15 13 15 2 16 15 0 9 13 1 9 0 9 9 2 3 15 15 4 13 3 0 9 16 9 1 0 7 0 9 2
29 9 1 0 7 0 15 13 3 3 15 3 0 2 2 13 9 11 11 11 7 13 1 9 0 1 9 9 9 2
18 9 1 9 0 9 15 13 0 9 9 9 9 7 0 9 11 11 2
15 9 9 2 0 1 0 9 9 2 13 9 1 0 9 2
38 11 13 2 16 1 9 4 15 7 1 9 1 9 13 10 9 13 0 2 9 2 3 0 9 9 1 0 9 2 3 10 0 9 1 9 0 9 2
32 9 11 13 2 16 0 9 13 1 9 0 9 2 7 13 4 15 13 0 9 2 15 4 13 0 9 2 7 13 10 9 2
14 1 0 9 9 1 9 13 7 11 7 11 2 11 2
26 10 9 13 1 15 2 16 9 13 13 9 9 9 1 9 2 15 13 0 9 2 3 9 1 9 2
31 1 9 1 9 9 9 1 9 3 13 9 2 16 9 13 14 0 2 7 7 15 2 15 15 0 9 13 1 3 0 2
8 9 14 3 1 11 16 1 9
2 11 2
29 9 9 9 12 12 9 1 9 15 9 9 9 1 0 9 1 9 0 9 1 11 13 9 13 15 0 9 9 2
16 13 15 3 1 9 9 11 12 7 12 9 9 11 11 11 2
17 9 1 15 13 13 9 9 9 2 16 4 15 10 9 9 13 2
20 1 9 2 16 15 13 1 0 9 1 9 2 11 13 2 16 3 1 9 2
26 9 11 11 11 13 2 16 9 4 13 13 3 14 10 9 2 1 10 9 4 13 13 10 0 9 2
19 2 13 2 16 13 9 10 0 9 2 15 9 13 10 9 2 2 13 2
12 1 11 1 15 13 1 9 0 9 0 9 2
9 9 0 0 9 13 3 1 0 9
2 11 2
35 9 1 0 9 1 9 0 9 1 0 9 1 11 2 15 13 9 9 2 13 14 9 9 11 2 7 2 3 13 11 2 7 9 9 2
22 0 9 0 9 13 1 9 11 0 1 9 9 7 1 9 1 9 12 9 13 9 2
15 9 9 13 13 1 0 2 0 2 7 0 9 1 9 2
38 13 3 1 9 2 3 15 13 2 16 2 0 7 0 0 9 1 0 9 7 0 9 2 15 4 11 13 2 13 3 0 7 13 9 1 9 2 2
6 3 13 7 9 9 2
35 1 9 2 3 13 0 0 9 2 9 9 9 11 0 0 9 13 2 16 10 9 13 0 0 9 13 3 2 16 13 9 11 7 11 2
39 0 9 4 3 13 2 16 4 15 12 9 13 1 15 2 16 13 0 13 1 0 9 0 9 16 1 11 2 7 1 11 2 7 16 15 0 9 13 2
30 11 11 3 13 9 9 11 2 16 15 0 9 2 15 13 13 9 7 13 12 9 2 13 9 0 9 1 0 9 2
6 9 13 1 15 9 2
41 2 9 0 0 9 1 0 9 1 0 9 7 3 2 1 9 9 11 2 0 9 1 0 9 1 0 9 4 9 0 9 1 9 13 3 3 2 2 13 11 2
26 1 0 9 0 9 7 1 9 9 9 13 3 14 12 0 9 1 12 9 0 1 9 1 0 9 2
19 0 14 12 9 9 13 3 0 7 13 14 0 9 13 15 1 0 9 2
6 1 11 15 13 1 9
14 9 11 13 2 16 4 15 1 9 0 9 13 1 9
2 11 2
27 7 16 4 3 1 9 0 9 11 2 9 2 13 3 12 12 9 12 9 2 13 13 1 3 0 9 2
22 1 9 1 9 9 9 0 2 9 11 9 15 13 9 0 9 11 11 2 11 2 2
23 0 9 1 11 13 7 9 15 2 15 4 15 1 11 13 2 16 4 0 9 4 13 2
8 0 9 3 13 14 12 9 2
32 11 1 9 1 0 9 1 9 9 13 2 16 0 9 0 9 1 0 9 13 0 2 9 13 7 0 0 9 7 0 9 2
39 16 15 0 9 1 12 7 12 9 13 2 13 9 3 13 1 12 12 9 12 3 2 16 1 0 9 9 2 3 12 9 2 4 10 0 9 3 13 2
20 12 0 9 9 4 13 1 0 9 2 3 13 4 13 0 2 9 0 9 2
14 9 11 13 2 16 9 13 9 9 1 3 0 9 2
23 1 9 0 0 9 14 13 9 9 9 7 9 1 9 2 1 9 0 9 2 13 0 2
18 12 9 0 9 15 1 11 13 0 0 9 2 9 4 13 1 9 2
7 9 9 13 3 12 9 2
24 15 9 0 9 14 9 13 1 9 9 2 9 7 9 0 9 2 0 9 7 9 0 9 2
39 1 0 9 2 16 15 9 9 13 9 9 1 0 9 2 11 13 2 16 9 3 13 9 9 9 9 12 9 9 7 12 9 13 1 0 7 0 9 2
17 3 0 9 1 0 0 9 9 9 0 9 11 13 1 9 0 2
12 0 9 9 13 13 3 9 1 9 9 9 2
27 0 9 1 9 2 9 7 0 9 13 1 9 3 1 11 1 0 11 2 0 9 9 7 9 11 11 2
11 9 15 13 1 12 9 1 9 0 9 2
5 0 9 13 7 9
2 11 2
27 9 1 0 15 9 0 9 0 9 1 11 13 1 9 0 0 9 0 2 11 2 0 9 9 0 0 2
22 13 3 1 9 2 1 15 15 1 9 13 7 13 2 7 3 1 2 9 2 9 2
7 0 9 0 9 13 11 2
17 9 9 1 9 11 11 13 2 16 4 9 4 13 0 0 9 2
16 1 9 9 11 13 9 7 9 2 16 4 1 0 9 13 2
26 2 13 7 3 0 15 13 2 16 9 7 9 10 9 13 3 0 7 11 15 13 1 10 0 9 2
26 13 15 3 13 1 0 9 2 7 16 7 15 13 13 1 0 0 9 2 2 13 9 0 9 9 2
23 9 11 13 3 1 9 2 16 0 9 13 9 0 0 9 7 1 0 9 13 14 3 2
11 0 9 13 0 0 9 0 16 0 9 2
19 3 15 7 13 1 9 1 0 9 9 7 1 0 9 1 9 0 9 2
5 0 9 13 1 9
2 11 2
15 1 0 9 0 9 0 9 15 3 1 9 9 13 9 2
18 7 16 15 9 9 3 13 2 1 10 9 15 1 10 9 13 3 2
34 9 9 0 9 11 11 1 15 13 2 16 16 0 9 9 13 2 9 15 13 1 0 9 13 9 2 15 13 9 9 9 0 9 2
6 9 3 13 0 9 2
15 0 9 9 13 0 9 2 1 15 13 10 9 9 13 2
9 0 9 13 13 0 9 0 9 2
21 3 15 7 13 13 2 16 13 9 13 0 9 7 9 9 1 9 7 1 9 2
11 1 11 9 0 9 9 3 13 7 13 2
3 0 9 9
2 11 2
18 0 0 9 2 9 9 15 13 1 11 1 0 9 9 11 1 11 2
22 0 0 9 1 11 7 13 0 0 9 7 13 0 9 1 0 9 7 1 0 9 2
11 0 9 1 9 9 9 13 13 0 9 2
9 9 13 9 7 9 1 0 9 2
10 9 4 13 9 9 7 13 0 9 2
16 9 13 1 10 9 12 9 2 3 3 4 9 13 1 0 2
12 9 13 0 9 0 9 2 0 9 9 0 2
7 9 13 0 3 1 9 2
16 0 13 3 9 9 2 1 15 13 9 0 7 0 0 9 2
6 2 9 9 2 1 9
3 11 11 2
25 3 16 12 9 9 9 9 7 0 9 0 11 13 1 9 1 11 11 1 2 9 0 9 2 2
21 1 9 1 9 15 13 9 14 12 9 13 9 9 2 1 15 13 7 9 9 2
9 0 0 9 7 9 12 9 13 2
28 9 2 15 13 1 9 9 0 0 9 7 13 9 1 9 0 1 9 9 2 1 12 9 1 9 9 13 2
21 0 9 11 1 9 12 15 1 9 1 11 13 12 0 11 11 2 9 9 1 11
3 11 13 9
15 9 11 1 9 13 2 16 1 0 9 13 0 9 9 2
28 1 12 1 12 7 12 9 1 9 1 9 9 0 7 1 12 1 12 7 12 9 1 9 1 9 9 0 2
22 9 15 1 15 13 1 9 9 2 16 9 9 3 1 0 9 9 3 13 0 9 2
8 0 9 9 13 9 3 0 2
16 3 10 9 2 7 3 9 9 2 13 0 1 9 0 9 2
15 1 9 7 13 9 2 3 1 0 9 9 13 3 3 2
17 7 3 0 9 15 1 9 2 13 2 3 1 9 9 0 11 2
13 3 1 9 0 0 9 13 3 1 12 0 9 2
13 1 1 10 0 9 13 7 3 14 1 0 9 2
38 11 13 2 16 9 4 3 3 13 2 16 10 9 13 0 0 9 0 9 7 16 13 15 1 9 9 3 13 1 15 3 0 2 16 13 9 0 2
24 0 9 1 0 9 9 9 2 7 15 7 9 0 9 2 13 9 3 0 9 1 9 9 2
21 13 0 2 16 13 0 9 2 15 4 13 1 0 9 7 13 1 9 0 9 2
23 1 9 9 0 9 2 3 1 0 9 0 9 2 7 0 0 9 3 3 13 0 9 2
14 9 15 13 13 13 2 4 3 9 13 14 1 9 2
16 13 3 10 2 0 9 15 0 2 9 9 0 0 0 9 2
21 13 15 1 15 9 9 1 9 2 0 0 0 9 2 0 9 9 1 0 9 2
4 15 3 14 2
7 7 7 15 13 9 0 2
31 9 3 1 9 0 0 0 9 13 1 10 9 0 9 7 2 16 4 15 3 13 1 9 2 15 9 13 1 9 0 2
2 3 2
6 1 9 12 13 9 2
39 9 11 2 11 2 3 13 2 16 0 0 9 4 15 13 0 0 9 2 7 7 15 1 9 13 2 16 4 2 9 2 1 0 9 9 13 0 9 2
19 9 7 13 2 16 9 0 0 9 9 4 13 1 9 0 0 0 9 2
6 9 11 13 1 11 9
2 11 2
13 0 9 13 1 9 1 11 0 9 9 11 11 2
28 9 0 9 1 11 2 15 0 0 9 1 9 13 9 1 10 9 9 2 13 1 0 7 0 9 1 9 2
35 0 9 9 9 9 13 9 2 15 9 11 13 3 1 12 9 2 1 15 13 7 0 0 9 11 11 7 0 9 7 0 9 11 11 2
16 0 13 7 10 9 7 9 2 3 0 2 7 0 0 9 2
20 9 0 11 1 11 4 13 9 11 1 9 10 9 11 1 9 0 2 9 2
11 15 13 0 11 1 11 9 12 1 11 2
6 11 1 11 13 1 9
2 11 2
23 3 0 9 0 9 1 9 1 0 11 7 9 0 9 13 1 11 0 9 9 0 9 2
21 0 9 9 11 11 13 9 12 9 1 12 10 0 9 11 11 3 1 0 9 2
26 9 9 13 7 11 11 2 15 13 3 0 9 11 7 3 13 9 9 11 0 15 1 0 11 11 2
17 0 9 11 15 13 11 11 2 11 11 2 11 11 7 11 11 2
25 9 13 0 9 1 0 7 0 9 2 15 4 7 1 12 9 13 13 9 9 7 0 9 11 2
14 1 0 9 0 9 13 11 9 0 0 9 1 11 2
23 11 13 2 16 1 0 9 13 11 0 9 2 3 4 13 1 0 9 13 9 0 9 2
14 0 9 0 9 13 1 9 1 9 0 1 9 9 2
16 13 15 3 1 9 2 7 3 3 14 4 13 13 10 9 2
24 2 9 13 0 2 13 0 15 0 13 2 2 13 9 0 9 11 11 2 1 9 3 2 2
20 0 9 2 15 1 9 1 11 13 0 9 2 13 0 0 9 1 9 9 2
6 1 9 0 9 1 11
5 9 15 13 1 9
11 13 7 9 10 9 2 3 14 13 1 9
2 11 2
26 0 0 9 13 3 13 1 9 9 7 10 9 4 13 13 3 10 9 1 0 9 1 9 9 9 2
19 1 9 0 9 1 9 11 3 13 0 0 9 9 1 0 9 1 11 2
23 9 15 13 3 2 16 9 9 9 13 9 0 9 9 3 1 9 9 9 7 9 9 2
15 9 7 3 13 1 0 9 1 9 9 2 9 7 9 2
16 9 3 13 13 3 9 1 0 9 9 2 3 1 9 9 2
28 1 9 9 15 13 1 9 2 15 15 13 2 16 4 13 10 9 0 9 7 3 15 13 9 1 9 9 2
11 0 9 4 13 1 0 2 3 3 0 2
26 2 10 9 13 13 0 9 2 7 3 15 13 13 7 1 0 9 2 2 13 9 9 9 11 11 2
38 15 15 13 9 2 16 1 9 1 9 4 13 3 2 16 3 1 9 9 4 1 9 1 9 13 0 9 1 2 9 0 9 9 7 9 9 2 2
15 9 1 0 13 9 9 2 0 9 9 7 9 9 9 2
12 3 9 9 13 9 7 15 13 1 0 9 2
13 11 13 2 16 9 9 4 15 13 13 7 9 2
21 10 9 0 9 13 1 9 3 0 7 13 2 16 4 1 9 4 13 7 9 2
5 15 7 11 13 2
10 2 13 9 2 7 9 2 2 13 2
7 1 9 13 3 9 11 2
11 13 2 16 10 9 13 0 0 9 11 2
21 13 3 2 2 4 15 13 13 9 9 1 15 9 3 2 3 3 4 13 2 2
5 9 1 9 13 9
6 2 9 1 0 9 2
5 14 2 0 9 2
30 0 9 1 9 4 13 1 0 9 13 1 12 9 9 3 1 12 9 9 3 7 1 9 12 1 0 12 9 9 2
19 9 13 1 12 9 1 9 1 9 9 12 1 12 9 1 9 9 12 2
16 13 15 1 9 9 1 0 9 11 2 15 4 13 0 9 2
16 1 15 1 0 9 9 1 9 13 14 1 12 12 9 3 2
26 9 9 9 1 0 12 9 13 9 9 1 9 1 0 15 0 9 7 0 9 1 9 0 0 9 2
24 9 9 1 0 0 9 7 0 11 3 7 1 0 9 1 0 9 13 1 12 12 9 3 2
16 9 1 9 11 15 13 1 12 12 9 3 1 12 0 9 2
36 0 9 13 1 0 9 0 0 9 9 0 9 1 0 9 7 0 9 0 9 7 9 1 10 2 16 4 15 13 13 1 0 9 0 9 2
18 2 1 9 0 7 0 11 10 9 3 13 2 2 13 15 1 9 2
22 9 4 13 2 16 4 9 13 13 9 0 9 0 1 9 9 9 0 11 1 11 2
9 9 1 9 3 13 11 7 11 2
9 0 9 4 13 9 1 9 12 2
13 3 4 13 1 0 9 13 9 3 11 7 11 2
16 0 9 3 7 13 0 9 9 9 7 9 1 9 10 9 2
23 0 9 15 13 1 9 2 16 4 13 13 1 9 9 9 11 1 0 11 1 9 9 2
4 0 9 0 9
13 3 0 2 14 2 0 2 9 13 9 10 0 9
27 11 2 11 2 11 2 11 1 11 2 11 2 0 9 2 0 9 2 0 9 2 15 13 10 9 0 2
9 9 9 2 9 9 7 0 9 2
18 13 1 0 9 2 15 4 15 13 0 9 1 0 9 2 3 13 2
16 9 13 3 0 9 7 13 15 1 0 9 13 1 0 9 2
21 10 9 2 15 13 9 2 13 7 3 15 0 1 11 2 11 2 11 7 11 2
21 3 1 9 2 15 13 3 0 9 9 2 0 9 7 1 9 11 9 9 13 2
30 15 10 12 9 9 13 2 13 15 2 15 15 13 14 2 0 9 2 7 0 9 2 3 15 1 9 10 9 13 2
30 0 9 13 1 3 0 9 2 3 1 9 3 0 7 3 0 9 9 1 0 9 2 7 13 15 3 1 9 0 2
41 1 0 9 13 7 13 0 9 2 9 2 9 9 2 9 7 0 9 2 3 15 9 2 15 13 3 9 0 9 0 9 2 9 2 7 13 0 1 0 9 2
13 0 0 9 13 13 1 0 9 1 9 9 9 2
12 13 0 9 2 0 9 13 13 1 9 9 2
17 0 9 4 3 3 13 0 9 7 13 4 3 9 1 0 9 2
32 3 15 13 3 2 12 9 1 9 0 9 15 1 10 0 9 13 2 9 2 9 2 15 13 2 7 13 13 1 0 9 2
14 13 7 9 1 9 7 15 0 15 13 9 0 9 2
36 0 9 9 10 9 13 9 2 16 0 9 15 13 9 9 7 14 0 9 9 7 9 1 15 2 16 9 10 9 13 13 3 3 9 9 2
36 3 7 3 14 9 13 9 1 9 9 2 0 7 0 9 0 9 13 9 9 1 9 9 2 15 1 10 9 13 3 9 2 3 11 2 2
37 0 9 9 0 9 13 3 0 9 10 9 2 15 15 3 9 1 9 13 2 7 3 13 3 0 16 1 0 9 2 1 10 9 1 0 9 2
26 0 9 15 13 3 3 13 1 0 9 2 7 13 0 15 13 2 16 10 0 9 13 13 15 0 2
18 10 9 2 1 9 13 0 9 2 13 9 7 1 0 9 0 9 2
53 1 0 9 2 3 1 0 9 2 9 0 9 0 9 13 0 9 0 1 0 9 2 16 10 9 13 9 3 13 2 16 4 4 13 10 2 9 2 16 9 10 9 2 7 9 9 1 10 9 1 0 9 2
19 10 9 2 3 1 9 0 0 9 2 3 13 1 9 1 9 0 9 2
26 1 0 9 0 9 1 11 13 13 13 9 9 7 1 9 1 9 1 9 1 9 1 15 13 9 2
30 15 2 13 2 14 3 9 9 13 7 16 9 0 9 2 0 9 2 16 9 0 9 3 3 3 10 9 13 2 2
13 9 0 9 7 13 9 0 9 1 3 0 9 2
16 1 0 9 13 15 0 1 9 2 15 15 1 10 9 13 2
38 15 0 2 3 10 0 9 2 13 9 1 9 1 10 9 2 7 16 10 9 13 13 3 0 2 1 1 15 2 16 1 9 0 9 13 13 15 2
10 3 7 13 0 13 9 1 0 9 2
6 3 14 3 13 13 2
49 1 0 9 2 9 15 3 13 1 0 9 2 16 1 9 13 13 3 10 9 2 0 9 2 9 9 2 9 1 9 2 1 9 9 7 3 2 15 13 1 0 9 9 1 9 13 0 9 2
18 0 9 15 1 9 9 13 1 0 9 2 1 10 9 1 0 9 2
11 13 15 15 2 15 9 1 9 9 13 2
9 0 9 13 3 0 9 0 9 2
30 9 9 13 1 0 9 13 1 9 2 3 13 0 0 9 2 3 13 13 9 1 9 7 3 13 3 3 0 13 2
23 9 9 0 9 13 3 0 2 13 15 9 9 1 9 0 2 15 9 9 0 9 13 2
12 9 9 4 13 10 0 9 7 13 9 11 2
11 9 10 9 13 4 3 13 1 9 9 2
25 1 9 0 9 13 9 9 9 2 15 13 0 9 0 9 7 15 13 9 9 1 10 0 9 2
14 9 10 9 15 13 0 0 0 9 2 15 13 9 2
32 10 0 9 13 3 1 10 9 13 10 0 9 2 0 7 0 0 9 2 2 1 15 15 9 13 7 15 0 9 3 13 2
20 9 1 9 9 2 3 1 11 2 13 12 0 9 2 15 13 14 12 9 2
15 10 9 1 0 9 15 1 15 3 13 2 13 3 0 2
36 3 13 9 9 14 2 0 9 3 0 2 7 1 10 9 1 15 13 0 9 2 15 13 2 1 15 7 3 15 13 7 13 15 0 9 2
42 1 11 13 9 3 16 12 12 0 9 2 3 3 0 9 16 11 2 0 0 2 9 11 2 12 9 2 1 15 3 7 9 0 1 11 2 7 7 12 0 9 2
20 1 0 9 13 1 11 0 9 7 10 11 2 7 13 3 1 0 9 0 2
10 9 9 0 9 13 1 9 3 0 2
13 14 1 0 9 0 9 4 13 9 9 10 9 2
3 0 0 9
17 1 9 12 15 11 13 9 1 0 9 0 9 1 9 1 9 2
10 13 15 0 11 0 11 2 11 2 2
19 1 10 9 3 4 13 0 12 0 9 2 0 15 3 1 9 0 9 2
10 3 7 2 16 0 9 13 15 0 2
15 1 0 9 13 13 12 0 9 2 12 0 7 12 0 2
16 1 9 13 3 13 12 0 9 2 10 9 13 12 9 9 2
21 1 15 13 3 13 3 16 12 12 9 2 1 15 12 5 13 1 9 0 0 2
23 1 9 9 7 9 2 15 13 9 9 0 9 2 15 3 15 2 11 2 13 15 13 2
25 15 2 15 15 13 2 13 13 2 16 1 0 9 2 0 0 9 2 3 13 7 3 0 9 2
8 12 1 10 9 13 7 11 2
4 0 11 1 11
5 14 2 0 9 2
8 9 0 9 1 11 13 0 2
11 0 13 0 9 1 0 9 1 3 0 2
15 13 1 15 7 11 2 11 2 15 13 9 0 0 9 2
24 0 9 13 1 9 0 2 0 2 11 9 9 2 7 1 0 9 15 13 1 10 0 9 2
22 13 4 13 13 0 9 9 2 9 7 9 0 9 2 0 9 4 13 1 9 9 2
30 9 4 13 13 0 0 2 0 9 7 1 9 13 14 12 9 3 2 16 9 0 9 4 15 13 13 1 12 9 2
24 1 0 9 13 3 9 7 1 0 0 9 2 16 13 3 0 9 7 0 9 1 12 9 2
11 13 15 7 0 9 0 9 11 1 11 2
16 9 9 13 14 1 9 12 2 3 13 9 1 9 0 9 2
23 1 0 9 13 11 7 1 9 12 2 7 9 9 13 12 9 0 1 9 12 1 11 2
26 1 0 9 15 13 1 9 11 1 9 12 7 3 1 12 9 3 13 9 1 9 9 0 0 9 2
30 13 0 3 0 9 2 16 3 1 9 12 13 0 9 9 1 11 7 1 9 12 4 13 9 11 2 11 11 0 2
19 1 9 12 7 12 13 12 0 9 1 9 0 9 12 11 0 9 12 2
20 3 4 13 9 1 11 7 0 9 11 1 0 9 0 9 1 9 0 11 2
5 0 9 3 13 2
36 11 2 11 13 14 1 9 12 12 0 7 12 0 9 1 11 7 1 0 9 9 7 0 9 13 12 0 9 1 9 2 9 7 9 11 2
18 3 15 1 11 13 1 9 0 9 1 0 9 10 9 3 1 11 2
14 1 0 0 9 4 15 15 13 13 9 7 0 9 2
6 9 1 0 9 7 9
13 9 0 9 0 0 9 13 0 1 15 9 11 2
16 10 0 9 15 13 13 15 12 9 9 11 0 1 10 9 2
13 1 0 0 9 4 15 13 9 13 1 0 9 2
17 3 0 0 9 13 0 9 3 1 0 9 9 7 9 1 9 2
15 9 13 9 2 7 10 0 9 2 9 7 0 9 9 2
5 13 13 9 9 2
23 13 4 9 1 9 13 12 0 9 7 13 15 2 3 3 4 13 1 9 1 10 9 2
22 3 15 1 0 9 13 7 3 9 7 1 15 15 1 9 1 3 0 9 15 13 2
7 3 0 9 13 3 13 2
19 0 13 7 3 0 0 9 1 9 0 9 7 3 13 1 9 0 9 2
8 0 13 7 9 10 0 9 2
15 1 9 13 15 7 0 9 1 0 9 7 9 1 9 2
20 3 16 0 13 9 2 0 12 9 7 15 15 13 3 13 9 9 0 9 2
26 1 0 9 13 9 9 2 0 9 9 2 0 9 0 9 2 9 0 9 7 0 9 1 9 9 2
24 1 9 11 13 0 15 13 1 0 9 9 7 9 9 2 15 7 15 13 3 16 0 9 2
14 0 9 1 0 9 7 0 1 0 9 15 15 13 2
32 0 9 13 9 1 0 9 12 2 12 9 2 7 0 9 1 12 9 1 9 9 2 1 0 9 12 9 2 0 0 9 2
28 15 13 7 1 0 9 2 16 1 0 9 9 9 13 3 3 2 7 16 13 9 3 0 9 1 9 9 2
32 9 15 3 13 13 10 9 16 0 0 9 2 7 15 15 13 0 9 7 0 7 0 9 7 1 9 1 12 9 2 9 2
25 1 9 7 0 9 7 1 10 9 13 1 9 0 9 2 15 7 13 10 9 1 0 9 9 2
16 11 11 13 3 0 0 9 2 15 13 7 7 0 0 9 2
18 10 0 9 7 3 0 9 13 16 1 0 9 2 7 1 0 9 2
1 3
21 0 0 9 11 13 2 16 1 0 9 3 16 13 10 9 1 0 9 0 9 2
12 0 9 15 1 0 9 13 1 12 9 9 2
26 0 0 9 11 13 1 0 9 1 0 9 1 0 9 0 9 12 9 0 9 2 12 9 9 2 2
20 1 0 9 15 13 12 9 11 2 15 13 1 12 9 3 16 1 9 12 2
11 0 9 13 0 2 9 2 3 1 11 2
30 9 2 15 13 0 9 1 9 1 12 9 7 1 9 1 12 9 1 9 2 13 4 1 10 9 3 13 0 9 2
26 13 2 14 15 9 10 9 3 2 4 15 0 9 13 1 12 9 2 1 0 9 3 1 12 9 2
7 9 13 1 9 9 3 2
10 11 15 13 3 13 0 9 0 9 2
22 7 7 1 9 9 11 11 13 3 14 9 2 0 9 2 2 15 13 9 11 11 2
14 10 9 4 13 13 3 0 15 9 1 0 9 9 2
23 9 1 9 11 9 0 9 13 0 9 1 9 12 9 0 9 12 9 2 12 9 2 2
4 9 13 3 9
8 0 9 13 9 13 1 0 9
28 1 9 0 9 2 3 1 12 2 9 12 2 4 13 9 3 0 9 1 0 9 9 0 9 1 0 9 2
12 9 0 9 13 3 1 9 1 0 0 9 2
14 15 0 9 7 13 0 3 1 9 9 1 0 9 2
16 2 10 9 15 13 9 9 1 0 9 0 9 1 0 9 2
40 1 9 15 13 1 9 7 9 0 9 9 2 15 13 0 1 9 9 7 1 9 9 2 2 13 9 2 11 11 2 9 9 11 1 9 0 7 0 9 2
7 7 9 10 9 3 13 2
21 2 1 9 13 4 9 9 13 0 9 2 2 13 9 2 11 1 9 1 9 2
27 1 0 9 13 1 9 10 9 12 9 0 9 2 11 2 2 15 13 0 9 1 9 12 2 12 2 2
10 2 3 0 9 13 3 12 0 11 2
8 0 0 9 13 12 9 9 2
26 0 11 2 15 4 3 3 13 1 0 9 1 11 2 13 1 12 9 13 12 0 7 12 0 9 2
15 16 13 9 2 13 0 13 0 9 7 3 13 7 9 2
14 3 4 13 2 16 4 9 13 0 9 1 0 9 2
12 1 9 7 1 9 13 13 3 0 9 2 2
28 9 0 9 13 0 13 10 9 1 0 1 0 0 9 1 9 9 1 12 9 1 12 9 1 9 9 9 2
7 10 9 13 7 3 0 2
25 16 15 13 7 13 1 9 12 0 9 0 3 1 9 12 2 3 15 13 3 13 1 0 9 2
21 2 13 9 1 0 9 2 13 3 1 9 9 12 9 2 2 13 9 2 11 2
10 1 9 0 9 3 13 7 9 9 2
8 0 9 4 3 12 9 13 2
12 9 9 10 9 13 9 2 11 11 1 11 2
22 2 1 9 11 15 13 1 0 9 0 9 9 7 1 2 9 2 15 13 10 9 2
12 1 9 9 15 3 7 13 2 3 13 9 2
8 15 13 0 9 10 9 2 2
11 1 11 4 13 9 13 9 1 9 9 2
13 15 13 13 0 9 1 12 9 2 13 0 9 2
9 2 0 9 4 15 9 13 13 2
9 3 0 9 1 15 13 13 9 2
16 1 11 3 13 13 1 2 9 2 2 3 15 1 9 13 2
7 3 14 9 13 9 9 2
18 16 13 15 1 9 2 1 0 9 1 9 15 13 3 14 0 9 2
11 13 7 7 0 2 2 13 9 2 11 2
7 9 11 4 0 9 13 2
19 9 15 13 1 12 1 12 9 2 7 9 11 13 3 1 10 12 9 2
22 9 9 2 3 1 1 3 16 9 9 4 13 9 9 2 13 9 12 7 12 9 2
14 2 13 15 1 9 2 16 9 13 3 7 3 0 2
9 13 7 13 0 9 1 0 9 2
17 16 13 1 9 0 9 0 13 9 2 3 3 9 13 3 3 2
16 7 15 13 1 9 2 7 1 9 2 2 13 9 2 11 2
20 15 13 11 2 13 4 13 0 9 7 9 1 0 7 3 7 0 0 9 2
18 16 7 13 0 9 0 1 9 2 4 15 13 3 14 9 1 9 2
14 0 9 13 3 0 9 2 1 15 4 13 0 9 2
4 11 13 9 9
18 0 9 1 0 9 13 3 0 9 2 0 3 0 9 1 0 9 2
41 1 9 11 7 1 15 0 9 2 10 9 4 3 3 13 2 13 9 2 3 0 7 9 0 2 15 13 0 9 0 2 0 2 0 2 3 2 7 0 9 2
10 10 9 13 1 9 12 7 12 9 2
10 13 10 9 1 15 0 9 1 9 2
33 15 15 3 13 1 9 9 0 9 1 0 9 2 1 9 1 9 1 10 9 2 1 0 9 2 9 2 2 1 9 13 3 2
6 1 11 0 9 13 2
19 3 3 1 9 0 0 9 7 9 9 7 9 13 3 16 12 12 9 2
17 13 15 3 0 7 0 9 3 1 0 9 7 1 9 0 9 2
58 10 9 1 9 13 3 0 9 1 0 9 13 1 0 9 1 9 9 7 9 11 11 15 2 16 1 9 9 0 0 9 2 15 13 0 9 9 9 2 13 1 12 2 9 12 0 9 11 1 0 9 2 13 0 9 0 9 2
48 3 13 11 9 9 0 0 9 11 11 2 11 15 13 1 12 0 9 9 2 1 0 1 9 1 9 7 9 0 9 2 0 9 1 9 7 9 7 0 9 7 1 0 1 0 0 9 2
21 15 13 0 0 9 1 0 9 7 0 9 1 0 0 9 7 1 0 0 9 2
60 3 2 1 9 1 9 0 2 3 2 0 9 9 0 0 9 1 9 0 9 7 1 0 9 0 1 9 2 11 1 15 13 1 9 9 12 2 12 2 12 2 2 1 15 13 0 7 3 0 9 1 0 9 1 0 9 1 0 9 2
33 3 13 11 9 9 1 12 9 9 0 9 1 0 9 2 1 0 9 4 10 9 1 0 9 13 1 9 9 2 9 2 9 2
10 3 13 0 9 0 1 0 9 9 2
7 3 0 13 0 9 11 2
21 10 9 3 13 1 9 12 7 12 0 9 7 13 1 3 0 9 9 7 9 2
21 1 10 0 7 0 9 13 11 0 7 0 9 10 0 9 2 9 0 0 9 2
36 9 2 3 11 2 15 3 13 9 2 9 2 9 7 9 9 1 9 0 9 2 0 9 2 0 9 0 0 9 11 7 3 0 0 9 2
23 10 9 9 13 3 1 0 9 2 16 11 1 10 9 3 13 3 0 9 1 0 9 2
23 1 10 9 9 7 10 12 9 2 0 7 0 7 11 2 13 9 10 9 1 9 12 2
16 1 10 9 4 0 9 7 9 13 1 0 9 7 0 9 2
4 11 13 13 9
12 9 1 9 7 9 13 9 1 0 9 7 9
4 11 2 11 2
16 2 0 2 9 13 0 9 9 2 1 0 14 1 15 0 2
9 9 13 1 10 9 3 1 9 2
15 13 3 3 7 3 1 0 9 2 16 3 1 9 13 2
16 9 10 9 13 9 9 2 7 9 2 3 0 2 13 9 2
29 7 15 10 9 13 1 0 2 9 2 2 15 7 3 13 1 9 9 1 9 7 10 9 13 0 1 10 9 2
19 13 7 7 3 0 7 0 9 2 3 0 11 2 0 3 1 9 9 2
16 10 9 13 1 9 0 0 9 7 3 13 1 12 0 9 2
16 0 9 15 10 9 13 1 0 9 2 13 9 11 11 11 2
23 3 13 1 10 9 9 9 2 15 4 3 13 1 0 2 1 0 9 3 12 9 9 2
13 11 15 13 3 3 0 7 0 9 3 0 9 2
18 13 9 2 3 1 15 13 9 12 9 7 15 13 3 9 0 9 2
30 3 1 11 13 11 2 11 2 13 15 9 1 9 11 2 1 0 13 12 9 2 7 13 15 2 16 13 15 9 2
13 2 0 13 1 11 2 15 13 3 3 3 9 2
30 1 12 7 12 9 4 3 13 9 1 9 1 12 9 9 7 9 1 12 9 3 13 13 2 2 13 11 2 11 2
11 10 9 13 0 1 12 7 12 9 9 2
15 11 13 1 3 0 0 9 2 15 13 12 9 0 9 2
14 9 13 0 3 1 9 2 3 9 13 10 9 3 2
16 16 15 13 13 9 9 2 13 11 1 10 9 9 10 9 2
19 1 9 0 1 0 9 15 9 3 13 2 16 4 13 1 9 1 9 2
24 1 15 4 13 13 10 9 3 3 2 16 1 11 2 11 13 9 1 15 0 9 0 9 2
24 3 0 9 2 3 13 9 3 1 9 9 7 10 9 13 2 13 1 9 11 14 12 9 2
24 1 15 9 15 9 9 13 9 13 2 13 0 9 7 15 0 9 13 1 9 1 0 9 2
13 9 13 2 1 0 9 13 3 3 2 13 11 2
13 1 15 0 13 0 13 3 9 1 0 9 3 2
28 0 9 2 15 9 9 13 1 9 9 2 13 0 9 1 9 2 9 2 9 2 0 9 7 3 1 9 2
23 0 13 3 9 9 1 9 7 9 1 9 1 0 9 2 9 2 15 13 0 9 11 2
7 15 15 13 1 9 9 2
28 9 0 9 13 1 15 1 9 9 9 11 11 0 9 2 7 13 1 10 9 0 1 12 7 12 9 9 2
23 11 15 13 0 0 9 1 0 9 2 2 13 1 9 9 2 1 9 12 7 12 9 2
21 15 0 9 9 1 10 9 13 2 15 13 9 0 2 1 12 9 15 13 15 2
29 1 0 9 9 13 11 7 9 9 0 1 9 0 9 2 15 15 13 13 10 9 3 1 12 9 1 9 9 2
5 9 13 0 9 9
3 11 11 2
35 9 0 9 7 9 2 15 4 13 0 7 0 9 1 9 2 9 2 9 7 0 9 2 13 12 2 9 1 11 11 9 0 0 9 2
24 10 9 1 9 4 13 1 12 0 9 2 9 0 9 2 0 9 7 9 1 0 0 9 2
20 9 4 13 1 9 1 9 11 11 2 15 13 12 1 9 0 9 1 9 2
12 3 1 9 9 9 4 13 7 0 9 9 2
16 0 9 3 13 2 10 0 9 13 1 9 14 1 9 9 2
5 14 2 0 9 2
2 11 2
17 9 1 9 1 0 9 3 7 1 0 9 9 9 1 9 13 2
19 1 9 9 0 9 9 7 9 11 15 13 1 11 7 1 0 0 9 2
20 0 0 9 1 9 0 9 7 13 7 9 13 7 3 9 1 0 9 13 2
14 9 9 1 0 9 13 1 0 9 14 1 9 9 2
15 1 9 15 1 0 9 9 10 0 0 9 3 3 13 2
25 9 11 3 13 0 9 1 9 3 0 9 1 9 14 1 9 9 7 1 9 9 1 12 9 2
14 1 9 1 9 7 1 9 1 9 9 13 12 9 2
19 1 9 0 9 13 9 1 9 1 10 0 0 9 1 11 1 12 9 2
24 11 13 0 9 1 9 11 2 9 7 11 3 12 9 2 15 13 3 3 16 1 0 9 2
29 1 0 9 9 1 0 9 11 2 15 15 13 1 9 2 13 3 9 1 0 9 1 12 9 2 0 12 9 2
21 0 9 11 1 11 11 13 1 9 9 1 0 9 0 9 1 9 1 12 9 2
11 0 9 13 1 0 9 13 3 12 9 2
26 7 16 15 1 9 0 9 0 2 11 11 11 13 9 1 9 2 9 15 13 2 7 3 3 13 2
25 1 10 9 3 9 13 1 11 16 9 1 9 2 7 3 13 13 2 16 15 0 13 3 3 2
46 0 0 9 2 3 13 3 9 2 13 1 0 9 1 11 2 3 12 9 13 1 9 3 12 9 2 1 0 11 12 9 2 11 12 9 7 1 11 12 9 7 1 11 12 9 2
19 16 15 9 0 9 1 0 9 13 3 2 9 0 9 13 1 9 0 2
23 1 0 9 1 15 13 12 9 9 2 1 15 13 9 14 14 12 9 13 1 0 9 2
8 3 9 0 9 13 3 0 2
8 3 9 15 3 13 1 11 2
10 9 1 9 13 1 10 9 3 0 2
16 14 1 0 12 9 3 13 7 1 0 9 13 12 9 9 2
4 0 9 3 13
3 9 1 11
2 11 2
43 0 9 1 0 9 9 1 0 9 7 9 3 1 9 11 13 1 9 1 12 5 2 15 13 10 0 9 1 9 12 2 3 1 9 3 15 1 15 13 9 9 13 2
5 9 11 11 13 2
9 10 0 9 9 3 13 12 5 2
3 9 9 13
2 11 2
22 0 9 9 13 1 0 9 12 9 9 2 15 13 1 12 9 3 16 1 0 9 2
8 13 15 1 9 0 0 9 2
44 0 9 1 10 9 13 11 2 3 9 9 13 1 12 9 7 13 12 9 9 2 7 11 2 3 15 3 13 12 9 9 9 2 15 13 1 12 9 3 16 1 9 12 2
12 9 9 15 13 7 1 11 2 11 7 11 2
16 9 9 1 11 3 13 1 12 9 7 13 9 12 9 9 2
17 11 15 3 1 9 9 13 1 0 9 1 0 11 7 0 9 2
14 3 13 11 2 11 2 11 2 11 2 11 7 11 2
6 0 9 15 1 11 13
2 11 2
15 0 9 1 0 9 13 1 0 9 1 11 11 2 11 2
21 9 12 0 0 0 9 1 0 9 1 0 0 9 1 9 12 13 9 0 9 2
22 0 9 13 0 0 9 0 9 2 15 15 13 3 2 16 0 9 15 13 9 12 2
6 1 11 13 3 3 9
2 11 2
16 0 0 9 11 1 0 9 13 1 11 7 1 11 12 9 2
16 13 15 0 9 1 12 0 9 0 9 11 1 0 9 11 2
14 1 9 1 9 12 15 13 9 9 0 3 1 9 2
11 0 9 13 11 11 3 7 1 0 9 2
27 1 0 9 9 2 1 11 2 11 7 11 11 13 12 9 2 9 2 1 12 5 3 16 1 9 12 2
18 3 1 9 12 0 9 11 1 9 12 13 9 0 9 1 0 9 2
17 3 13 1 12 11 12 2 12 7 12 9 11 9 12 2 12 2
17 1 11 11 3 13 12 9 3 2 15 13 3 1 15 0 9 2
12 9 1 0 9 1 9 11 11 2 0 0 9
29 15 15 3 0 9 13 9 13 1 10 0 9 1 0 2 0 9 2 16 15 15 13 2 16 9 1 15 13 2
25 0 9 15 15 15 13 1 0 9 2 3 16 1 11 13 10 9 7 4 3 13 15 1 15 2
37 13 9 1 0 9 7 13 15 2 16 3 2 16 15 9 13 2 13 0 9 15 13 1 9 9 10 9 2 1 0 9 2 10 0 7 0 2
37 15 4 1 15 13 1 0 10 0 9 7 1 0 9 2 3 1 9 11 2 7 13 4 15 1 15 2 16 10 9 4 15 3 15 13 13 2
51 9 7 9 13 13 10 9 2 15 13 0 2 16 4 4 13 16 9 1 10 9 7 9 0 9 10 0 9 2 7 3 16 10 9 2 15 4 13 0 9 0 9 7 1 10 9 3 13 3 13 2
15 15 15 13 2 16 3 0 9 1 9 13 13 3 13 2
8 10 9 15 15 1 15 13 2
23 1 9 13 10 9 2 15 2 16 15 9 11 7 11 13 2 3 1 15 13 3 3 2
12 7 2 15 13 1 15 2 16 4 15 13 2
21 3 4 13 9 7 3 15 13 10 0 0 9 10 9 2 15 4 13 1 9 2
7 10 9 0 9 7 3 2
34 3 15 13 2 16 15 2 15 9 11 7 11 13 2 15 13 2 10 0 9 2 7 10 9 7 9 2 15 3 13 2 3 13 2
5 3 15 13 13 2
51 3 15 15 13 7 15 4 13 2 16 15 15 3 13 7 7 15 13 2 7 3 15 15 13 2 16 12 1 0 9 13 3 2 7 15 13 7 13 15 1 15 0 9 2 7 16 15 4 13 3 2
8 7 15 15 3 3 3 13 2
77 13 15 9 0 2 13 15 9 9 0 9 2 0 9 2 0 9 7 15 3 13 2 16 13 0 9 9 0 0 9 2 3 3 15 13 2 0 15 0 2 3 1 12 0 9 3 13 0 16 9 7 0 16 0 2 16 13 10 9 0 2 7 3 15 9 13 16 9 0 9 7 14 16 10 0 9 2
10 13 15 2 16 13 1 15 3 13 2
18 7 1 0 9 15 13 2 16 15 14 13 1 9 2 9 13 3 2
3 1 0 9
5 2 9 0 9 2
5 14 2 0 9 2
57 9 2 11 13 9 0 9 2 2 2 9 9 7 9 2 2 2 11 11 13 9 9 2 2 2 9 1 9 2 7 2 11 2 9 15 13 13 9 2 13 9 7 9 0 0 0 9 1 9 11 11 1 0 2 0 9 2
14 11 11 13 0 9 1 9 0 9 2 13 0 11 2
27 11 15 13 1 15 2 15 15 13 9 1 12 9 2 13 4 13 1 9 2 16 4 15 13 9 9 2
28 1 9 0 2 11 0 9 13 1 11 7 11 2 16 4 3 13 1 9 7 16 4 13 3 9 7 9 2
34 0 0 11 15 13 2 16 11 3 13 3 7 3 16 3 15 9 13 1 9 9 7 9 2 15 1 9 13 9 0 9 1 11 2
22 9 12 4 15 13 1 9 11 7 11 13 9 0 9 7 0 9 2 13 0 11 2
17 11 11 1 15 13 0 0 9 2 16 13 1 0 9 12 9 2
23 13 3 3 2 16 13 9 2 16 13 10 9 2 7 14 14 0 9 2 13 0 9 2
34 11 15 13 13 1 9 2 15 13 0 9 2 9 11 11 1 9 9 1 10 9 1 0 0 9 2 13 9 0 0 0 9 11 2
37 1 0 9 7 9 1 12 2 9 9 9 7 15 9 0 9 13 11 3 0 0 9 2 7 15 13 3 0 2 0 7 0 2 13 9 11 2
4 15 4 3 13
5 14 2 0 9 2
10 4 4 13 2 7 13 4 15 0 2
48 11 11 2 9 9 1 0 9 9 2 1 12 2 9 9 11 0 9 2 13 15 15 2 7 1 9 13 3 12 2 9 2 2 9 2 9 2 2 9 2 9 2 7 9 2 9 2 2
24 0 9 9 11 2 12 9 2 2 11 2 10 0 9 2 13 10 0 9 1 9 2 2 2
25 0 9 11 1 9 0 9 1 11 2 11 13 0 2 14 3 0 9 7 1 0 9 1 9 2
21 9 0 9 11 11 1 12 2 9 2 2 11 2 3 13 2 2 13 3 13 2
20 0 9 0 11 2 10 0 9 13 9 0 9 7 9 11 1 10 0 9 2
35 9 0 0 0 9 2 11 2 11 11 2 13 1 9 1 9 7 15 2 15 13 1 9 0 9 7 9 9 2 15 1 15 13 13 2
27 9 0 9 11 11 1 9 2 16 10 11 13 9 11 11 2 15 1 9 13 12 9 9 1 0 9 2
20 13 4 0 9 7 13 4 15 1 0 9 2 15 13 0 1 15 0 9 2
22 0 0 9 11 11 1 9 0 9 1 9 1 11 2 13 15 1 9 15 13 0 2
56 11 11 2 0 9 7 0 2 9 2 0 9 1 9 1 11 2 1 10 9 7 1 9 9 2 16 1 11 7 0 9 13 3 13 12 0 9 2 15 10 9 1 0 9 7 11 13 3 0 2 16 15 13 1 9 2
24 0 0 9 11 1 9 0 9 2 16 11 7 11 13 0 9 9 16 9 1 0 0 9 2
4 11 13 0 2
24 3 15 13 16 0 9 2 3 16 0 11 2 9 9 2 7 16 9 0 1 9 10 9 2
21 1 0 9 15 13 13 0 9 1 12 7 13 3 0 9 9 7 0 9 9 2
3 0 9 11
7 0 11 2 0 9 0 2
5 14 2 0 9 2
12 0 9 11 11 1 10 0 9 13 0 9 2
34 16 13 1 0 9 9 2 9 1 10 9 13 3 9 0 2 9 0 2 1 11 7 0 9 2 13 0 9 0 0 9 0 11 2
40 2 0 9 2 0 9 2 3 3 13 1 9 2 3 7 13 13 2 16 0 0 9 9 4 1 3 0 0 2 0 9 13 16 0 9 2 2 13 9 2
25 2 1 0 9 15 13 9 2 16 0 9 11 13 13 12 2 9 9 9 16 9 1 0 9 2
17 11 7 3 13 2 16 1 11 13 3 0 9 9 13 1 9 2
17 0 0 9 7 1 15 13 1 9 0 9 2 2 13 0 11 2
27 1 12 9 13 11 9 1 9 2 10 0 9 4 7 1 0 2 0 9 13 13 9 9 2 13 9 2
1 3
22 0 0 9 11 7 0 9 11 13 1 9 9 9 1 9 7 9 1 12 2 9 2
23 9 11 1 0 0 9 13 3 12 9 9 2 15 13 1 12 9 3 16 1 9 12 2
8 9 0 9 13 12 9 9 2
13 9 9 13 1 12 1 12 11 1 9 0 9 2
15 9 1 15 13 3 13 13 1 9 10 0 9 1 9 2
22 0 9 1 11 1 9 1 12 9 1 9 12 15 1 0 0 9 13 1 12 5 2
23 0 0 9 2 9 2 11 2 11 7 0 9 2 15 3 9 11 1 9 12 13 13 2
15 0 9 13 3 9 1 12 5 2 0 9 1 12 5 2
4 9 9 13 9
8 1 0 9 13 1 0 9 9
2 11 2
15 0 9 0 9 3 13 2 16 15 1 9 13 0 9 2
10 11 15 13 11 11 1 0 9 11 2
15 9 9 7 0 9 9 13 1 10 9 1 9 0 9 2
43 0 2 7 16 3 0 9 2 10 9 15 4 13 9 9 1 0 9 0 9 7 9 3 0 9 2 13 13 9 0 9 2 3 9 0 9 2 15 13 1 0 9 2
14 10 9 13 9 1 9 1 0 7 1 9 0 9 2
27 0 9 13 0 0 9 1 9 9 12 2 15 15 13 1 9 7 0 9 2 3 13 0 7 0 9 2
15 1 9 12 15 3 13 7 0 9 7 9 1 0 9 2
22 1 9 9 12 10 9 13 1 0 9 1 12 9 7 1 9 13 9 12 9 9 2
20 9 15 13 1 9 2 16 9 9 13 15 1 9 1 0 9 13 3 0 2
14 0 9 2 16 3 0 9 2 3 13 1 9 9 2
26 10 9 1 0 9 13 3 0 0 9 1 9 2 15 13 9 13 1 9 2 1 9 1 0 9 2
12 1 3 12 9 9 13 10 9 9 12 9 2
12 0 9 13 12 9 9 7 0 9 12 9 2
15 3 0 9 15 1 11 2 11 4 3 13 1 9 9 2
24 2 16 13 13 10 9 2 15 9 13 2 16 0 9 13 0 9 1 0 9 2 2 13 2
18 3 13 2 1 9 1 0 9 13 3 13 9 1 9 3 0 9 2
25 10 0 0 9 15 13 1 15 2 16 9 9 1 0 9 1 0 9 13 0 9 3 3 3 2
27 9 2 3 9 7 9 9 13 0 9 2 15 3 13 2 7 13 1 0 9 7 2 0 2 0 9 2
13 3 9 0 9 13 1 10 9 3 9 9 9 2
4 0 11 7 9
2 11 2
50 1 9 13 1 0 9 0 9 13 1 11 9 11 9 1 9 1 0 9 0 11 2 12 9 2 2 10 9 1 1 0 0 9 3 13 3 0 0 9 9 2 15 13 0 9 11 0 11 11 2
49 0 9 9 1 0 9 13 0 9 7 9 9 9 13 1 10 9 2 16 9 0 9 2 3 9 11 2 13 9 1 9 0 9 0 0 9 1 11 7 0 9 2 16 0 9 13 1 9 2
36 0 9 9 1 10 9 13 2 16 1 0 9 1 10 9 13 7 16 0 12 5 0 9 13 1 0 9 1 0 9 0 9 1 0 9 2
13 1 0 9 9 13 1 9 0 9 13 0 9 2
5 0 9 13 1 11
11 0 9 13 14 12 7 3 16 10 0 9
2 11 2
23 0 9 0 0 9 12 9 3 13 1 9 3 3 15 16 0 9 1 0 9 7 11 2
12 13 15 3 1 9 1 9 0 9 0 11 2
26 16 15 0 9 13 0 9 1 9 0 9 2 13 3 9 2 4 13 3 12 7 3 16 1 11 2
22 1 0 9 1 0 9 1 11 7 0 9 9 13 9 9 2 0 0 9 9 9 2
33 3 15 1 15 13 2 0 9 9 13 0 2 7 1 0 9 13 0 0 9 7 9 0 7 0 9 2 7 13 0 0 9 2
32 9 3 13 2 16 1 9 1 0 9 0 9 13 9 1 0 9 2 16 3 2 3 13 0 9 9 2 13 9 3 0 2
34 0 9 3 13 9 0 9 12 0 9 9 2 9 12 2 1 0 9 1 11 2 15 15 13 13 0 7 0 9 0 2 0 9 2
24 0 9 1 0 9 11 11 13 2 2 13 13 3 0 0 9 2 16 4 0 9 13 2 2
21 11 13 1 9 0 9 1 9 1 9 7 3 1 15 13 11 2 11 7 11 2
13 3 13 1 15 0 9 0 11 2 13 0 9 2
3 9 3 13
1 9
2 11 2
13 3 15 13 0 0 9 1 0 9 1 12 9 2
9 13 15 1 0 9 0 0 9 2
25 1 9 1 12 7 3 9 13 9 9 1 0 9 3 12 9 9 7 1 9 0 12 9 9 2
18 1 0 9 1 12 2 9 12 15 1 12 9 13 0 12 9 9 2
21 0 0 9 9 15 1 0 9 1 9 12 13 1 12 0 9 7 13 12 9 2
20 9 13 3 12 9 2 15 1 9 1 0 9 9 12 13 9 1 12 9 2
6 9 15 13 1 0 9
2 11 2
17 0 9 2 0 9 1 0 9 2 4 3 13 1 0 9 11 2
29 0 9 9 2 15 13 0 0 9 0 0 11 2 13 9 2 0 9 1 0 9 2 9 7 9 7 9 9 2
17 1 9 9 15 0 9 1 0 9 0 9 13 12 9 0 9 2
19 1 9 7 1 15 3 13 9 9 11 11 7 9 0 0 9 11 11 2
6 0 9 13 12 9 2
4 0 9 1 11
2 11 2
27 0 12 0 0 9 1 9 13 1 0 9 9 1 11 0 0 9 1 9 9 9 1 0 2 0 9 2
30 0 9 9 2 0 3 12 9 2 9 0 0 9 2 13 3 13 14 12 9 2 0 12 9 11 3 1 12 9 2
24 3 3 13 9 9 0 9 9 9 11 11 2 0 9 10 9 13 0 16 1 0 9 11 2
16 0 9 13 1 9 1 12 9 2 15 13 0 1 9 9 2
16 9 9 7 9 13 9 9 1 0 9 2 15 13 13 0 2
26 9 9 13 9 9 3 0 0 9 2 7 7 0 1 0 9 2 15 15 13 13 1 0 9 9 2
4 11 13 0 9
2 11 2
21 0 9 1 9 7 9 13 1 0 9 13 9 11 1 0 9 0 7 0 9 2
7 3 15 13 0 9 11 2
21 0 9 9 13 1 9 0 9 1 0 7 0 0 9 7 9 1 9 10 9 2
4 10 9 1 11
9 0 0 9 15 3 0 0 9 13
2 11 2
31 0 9 9 11 11 13 9 9 0 2 16 15 3 13 12 0 9 2 9 7 9 1 9 9 2 2 1 15 13 13 2
19 11 15 3 13 11 11 2 9 0 9 1 11 2 15 13 9 1 9 2
17 9 11 13 1 15 2 16 0 9 4 13 13 13 1 0 9 2
16 2 1 9 15 2 15 13 2 15 13 13 2 2 13 11 2
27 0 9 1 11 7 12 2 9 13 2 16 9 13 0 0 0 9 2 15 4 13 13 1 0 9 9 2
17 0 0 9 1 11 11 11 3 11 13 2 16 0 9 3 13 2
17 13 7 2 16 1 15 9 9 0 9 1 11 9 3 13 13 2
24 2 3 1 9 9 13 9 7 0 9 13 2 16 9 13 1 9 1 9 2 2 13 11 2
11 0 9 1 11 4 13 3 12 2 9 2
14 9 3 13 12 9 1 9 2 16 4 13 9 9 2
26 1 9 13 11 13 10 9 9 1 0 7 0 9 2 16 15 3 3 13 9 2 15 13 10 9 2
7 13 3 1 12 9 9 2
12 3 15 3 13 13 9 10 9 1 0 9 2
10 15 4 15 13 13 9 0 9 9 2
10 15 0 9 4 1 9 0 9 13 2
5 2 15 13 9 2
19 13 13 7 9 2 7 3 7 15 13 2 2 13 11 3 11 2 11 2
6 1 9 9 15 13 2
22 0 9 11 11 1 9 2 3 13 10 0 9 1 9 2 13 1 0 9 0 9 2
17 9 13 0 9 2 7 0 9 9 13 1 9 9 0 1 11 2
23 1 9 2 15 1 11 13 2 13 7 9 11 2 15 13 9 1 9 9 1 9 9 2
20 15 11 3 1 9 10 9 13 2 13 7 2 3 1 9 2 0 0 9 2
4 10 10 9 0
2 0 9
19 3 13 15 3 16 12 9 2 7 1 0 9 1 9 0 9 3 13 2
46 13 4 3 10 9 1 9 2 7 7 4 15 9 3 9 1 9 14 1 9 13 3 1 9 0 9 7 3 13 1 9 7 9 2 7 9 13 9 13 14 3 7 9 3 3 2
19 15 13 3 1 9 2 13 3 9 7 13 15 1 9 13 1 0 9 2
39 1 10 9 15 3 13 1 15 2 16 4 9 13 16 9 1 9 2 7 1 0 9 15 15 13 9 0 2 14 2 9 2 7 15 3 7 1 9 2
50 0 0 9 13 9 2 10 9 1 0 9 13 13 9 7 9 2 9 0 0 9 2 2 15 9 2 0 0 9 2 2 15 9 2 0 7 0 9 2 7 15 0 0 9 2 0 1 9 2 2
26 1 9 4 15 3 13 13 7 0 9 0 0 9 7 9 11 11 2 15 4 13 1 9 0 9 2
30 4 4 15 15 15 13 2 13 15 2 16 10 9 7 9 3 13 2 16 4 9 13 0 9 0 9 1 0 9 2
24 13 4 15 2 16 4 9 13 2 16 0 9 15 13 13 3 16 12 2 7 3 12 9 2
6 13 15 3 0 9 2
21 3 13 15 3 2 3 7 9 9 15 13 3 3 16 9 9 1 9 0 9 2
7 7 15 9 0 0 9 2
4 7 0 9 2
5 7 3 7 9 2
6 15 13 1 0 9 2
22 1 9 4 3 13 0 9 2 0 9 2 15 3 13 1 10 9 0 9 7 9 2
25 16 4 15 15 13 2 15 13 0 9 1 9 0 9 0 9 1 9 2 3 15 13 1 9 2
3 0 9 2
5 9 9 7 9 2
5 3 14 2 2 2
16 7 2 13 2 1 10 9 4 0 9 13 13 14 3 3 2
16 13 9 9 13 3 14 15 0 2 16 13 9 7 13 9 2
15 0 9 2 3 14 2 7 14 16 13 1 15 9 0 2
8 3 16 1 15 13 1 9 2
27 3 4 15 13 13 15 2 13 4 15 2 16 4 10 9 13 14 7 2 16 4 1 15 9 13 9 2
27 13 15 13 2 3 4 15 9 13 9 2 16 4 13 1 9 14 7 2 16 13 9 7 13 10 9 2
7 15 4 15 10 9 13 2
4 15 3 14 2
7 3 3 9 9 7 9 2
11 9 15 1 15 13 9 3 7 9 3 2
14 13 15 9 2 13 7 13 15 1 10 10 10 9 2
51 3 4 15 7 13 13 2 16 14 15 2 7 7 0 0 9 13 2 16 4 10 9 13 1 9 1 9 1 9 2 2 2 3 7 1 10 9 2 16 15 13 1 9 0 2 1 1 9 0 9 2
5 11 13 1 0 9
2 11 2
21 11 11 2 0 11 13 1 9 1 0 9 1 9 12 1 9 0 9 0 9 2
12 11 15 13 9 0 9 9 0 9 11 11 2
36 1 9 2 15 9 13 9 9 2 15 11 2 11 2 0 1 11 2 13 1 0 1 9 0 9 2 15 4 13 9 0 9 9 1 11 2
25 9 9 1 0 9 13 1 15 2 16 0 2 3 0 9 2 15 13 1 0 0 9 2 13 2
6 9 13 1 0 9 2
26 1 9 0 9 3 4 13 9 2 1 15 13 0 9 13 9 9 9 0 15 1 9 9 9 9 2
18 1 15 2 3 0 9 1 9 11 13 2 15 9 2 11 13 13 2
22 11 11 15 3 0 9 13 9 0 9 0 9 11 2 1 10 13 9 1 9 12 2
29 3 2 3 0 9 1 11 13 0 9 0 9 1 0 11 13 9 2 13 15 11 2 11 1 9 1 0 9 2
4 9 13 11 9
2 11 2
17 9 11 11 13 3 9 11 11 7 1 0 9 13 10 0 9 2
8 13 15 3 0 9 11 9 2
23 1 9 9 13 2 16 0 9 1 11 11 13 1 9 2 15 13 0 9 1 9 9 2
9 9 1 9 9 13 7 9 13 2
18 11 11 13 9 11 11 2 0 9 2 15 13 1 9 1 9 12 2
44 11 2 11 13 3 1 9 13 1 0 9 9 1 0 9 2 16 3 13 16 1 9 2 7 3 9 7 0 9 1 11 2 15 15 13 0 9 2 1 15 10 9 13 2
20 0 9 1 11 13 0 9 1 11 9 7 15 10 9 1 9 13 0 9 2
23 1 0 9 15 11 2 11 1 9 13 7 12 1 15 13 7 13 7 9 1 0 9 2
24 10 0 9 2 1 0 9 12 7 0 9 2 1 9 13 9 2 16 4 0 9 11 13 2
40 9 0 9 11 11 1 10 0 9 13 2 16 11 11 4 13 1 9 7 2 16 10 9 1 9 12 1 9 12 13 3 3 2 16 15 13 0 9 13 2
5 9 13 9 1 9
7 11 11 4 0 13 9 11
2 11 2
20 3 13 9 3 1 0 9 1 11 2 13 9 7 13 15 14 11 13 9 2
20 3 15 0 9 11 9 13 0 0 9 9 11 11 2 1 9 0 9 9 2
17 2 16 15 3 13 2 13 4 15 7 3 13 2 2 13 3 2
18 0 9 0 9 7 11 15 3 9 1 0 0 9 1 15 9 13 2
19 2 13 4 9 2 16 4 15 13 2 7 15 3 15 15 7 13 13 2
11 13 4 15 9 2 2 13 3 0 9 2
36 3 3 3 13 0 9 2 16 13 2 2 13 13 1 15 2 16 1 9 13 13 9 9 14 11 7 0 0 9 9 4 13 14 9 11 2
9 0 4 15 3 9 11 13 2 2
20 0 9 7 11 13 1 9 11 2 3 15 1 9 12 2 9 13 0 11 2
10 2 9 1 0 9 4 15 0 13 2
19 3 0 9 15 13 3 1 0 9 2 3 4 15 13 13 12 9 2 2
10 1 0 0 9 13 9 1 9 0 2
33 2 3 13 3 1 9 9 2 1 0 13 0 0 9 7 1 9 2 15 4 0 13 2 13 0 13 9 9 2 2 13 9 2
20 1 9 3 9 11 11 13 12 9 2 1 15 3 3 11 13 1 0 9 2
14 9 11 1 11 15 3 13 2 1 9 11 7 13 2
9 1 9 13 1 11 13 0 9 2
48 16 13 9 11 1 0 9 9 3 1 9 2 2 16 4 13 0 9 3 3 2 1 9 4 13 11 2 2 13 9 2 15 0 9 13 2 16 4 15 15 13 1 0 9 0 9 11 2
22 2 13 1 9 2 2 13 1 9 9 2 15 1 9 1 12 0 9 13 12 9 2
25 0 9 11 2 12 2 9 2 12 9 2 12 9 2 12 9 2 9 12 2 12 2 12 9 2
18 13 2 11 2 0 11 2 2 11 2 9 1 11 13 1 9 2 2
30 13 2 11 2 11 2 12 9 1 11 2 2 11 2 9 1 11 2 2 11 2 1 9 2 2 9 2 11 2 2
3 9 0 9
9 1 11 13 1 9 9 3 14 11
2 11 2
24 1 9 2 16 1 9 9 13 1 9 3 14 9 11 2 13 1 0 0 9 11 9 11 2
15 11 2 15 13 12 1 12 0 9 11 2 13 0 9 2
22 9 3 13 0 0 9 9 11 2 11 2 7 9 11 2 3 11 2 3 11 2 2
18 2 3 15 15 13 13 9 1 9 2 3 13 3 0 9 14 11 2
15 0 15 13 1 9 0 9 13 2 2 13 9 11 11 2
17 1 0 9 13 11 12 9 2 11 12 2 11 12 7 11 12 2
23 3 0 9 13 3 3 1 9 2 3 13 0 9 9 9 11 2 13 15 1 11 2 2
6 10 9 15 3 13 2
20 11 15 7 1 10 9 3 13 1 0 11 2 15 15 9 11 13 1 11 2
15 11 13 1 0 9 12 9 2 15 1 0 9 13 3 2
10 2 3 13 3 0 9 3 1 11 2
14 16 4 13 2 13 4 14 3 2 2 13 9 11 2
25 0 9 11 2 12 2 9 2 12 9 2 12 9 2 12 9 2 9 12 2 12 2 12 9 2
29 13 2 11 2 9 1 11 2 2 11 2 11 2 2 11 2 11 2 9 1 11 11 2 2 11 2 11 2 2
23 13 2 11 2 11 2 2 9 2 11 2 9 1 11 2 2 11 2 9 1 11 2 2
5 0 9 1 11 2
6 11 11 13 9 0 9
2 11 2
27 2 13 1 0 9 13 3 3 7 13 15 13 1 0 9 2 2 13 1 0 9 9 11 11 11 11 2
23 10 9 7 9 11 1 12 9 11 11 7 13 1 0 9 7 13 2 2 13 15 3 2
23 1 0 9 4 13 2 16 16 4 13 13 1 11 2 13 4 13 9 2 15 13 9 2
18 9 0 9 3 13 2 16 10 0 9 13 2 13 1 0 9 2 2
34 9 1 9 13 3 9 9 11 1 0 11 1 0 9 2 1 15 15 0 9 3 3 13 12 9 2 7 3 13 9 1 9 9 2
22 13 0 0 9 11 2 3 1 0 11 13 1 9 12 9 2 4 13 11 1 11 2
48 2 3 9 13 3 1 0 0 9 2 2 13 0 9 11 2 7 3 13 2 16 1 11 4 13 9 0 9 2 2 11 13 0 9 2 11 9 9 13 7 13 10 0 9 3 0 9 2
15 13 7 9 9 2 1 9 15 4 13 1 0 9 2 2
7 11 13 1 0 9 0 2
32 1 0 0 9 1 0 9 2 15 9 11 13 3 1 2 0 0 9 2 13 9 1 9 0 9 1 0 9 0 11 11 2
20 0 9 9 2 15 10 0 9 4 3 13 1 0 9 2 7 13 14 9 2
25 0 9 11 2 12 2 9 2 12 9 2 12 9 2 12 9 2 9 12 2 12 2 12 9 2
7 13 2 11 2 11 2 2
30 13 2 11 2 9 1 11 2 2 11 2 11 2 12 1 9 9 1 11 2 2 11 2 1 9 9 1 11 2 2
21 0 9 9 11 2 3 2 15 13 1 9 11 11 11 13 9 1 9 1 0 9
9 11 1 11 13 2 7 3 3 13
3 0 11 2
23 14 9 11 11 12 9 1 9 9 0 0 0 9 13 1 9 12 2 12 11 1 11 2
27 9 2 1 10 9 3 13 0 9 11 11 2 13 1 12 12 12 2 12 2 7 0 3 13 3 13 2
19 11 13 1 10 9 12 9 2 0 1 15 13 10 12 2 9 1 9 2
16 1 9 13 3 0 11 11 2 15 1 9 13 3 9 9 2
11 11 13 1 11 13 1 12 9 1 15 2
24 11 2 15 1 12 9 0 9 13 12 9 2 13 13 1 0 12 9 3 9 1 10 9 2
7 3 13 12 9 0 9 2
26 1 9 9 0 9 13 11 9 11 2 15 13 1 11 12 2 12 7 13 0 9 1 0 12 9 2
7 12 9 9 13 11 11 2
25 11 11 13 12 9 11 1 10 0 9 1 11 7 13 10 9 1 9 1 0 9 9 0 9 2
22 9 13 11 2 12 2 12 2 3 3 3 7 1 0 12 0 9 13 3 3 13 2
12 0 9 9 13 9 11 11 2 0 9 11 2
23 0 9 0 2 11 9 7 10 0 0 9 1 0 12 9 11 11 1 0 9 9 13 2
12 9 13 0 9 9 11 11 15 2 13 2 2
15 11 3 13 9 1 10 9 1 11 9 1 9 1 11 2
18 11 7 13 0 9 2 7 3 15 1 9 13 1 10 9 11 11 2
14 11 13 2 16 16 15 15 15 13 13 2 4 13 2
15 11 13 3 0 9 9 2 15 15 13 13 0 0 9 2
37 11 13 3 3 1 0 2 11 1 9 2 16 4 13 11 1 11 11 2 7 1 0 9 11 13 7 13 3 11 11 2 11 11 7 11 11 2
24 15 11 13 9 13 7 1 11 2 11 2 0 11 2 0 11 11 2 0 11 11 7 11 2
13 3 15 3 13 11 11 2 16 13 9 11 11 2
5 11 1 11 1 11
2 11 2
37 11 1 11 2 11 3 1 11 7 11 1 11 2 15 13 0 9 0 12 2 9 0 9 2 1 15 15 4 13 1 0 9 9 1 9 14 2
21 9 13 13 7 11 2 15 3 3 13 9 1 9 7 13 9 9 0 9 11 2
31 11 4 13 9 1 9 2 16 9 11 7 11 13 9 1 9 2 11 13 1 9 1 11 0 0 9 7 9 13 9 2
15 11 4 13 9 11 1 9 7 11 1 0 9 1 9 2
13 9 11 3 3 13 2 7 10 0 9 13 0 2
25 1 11 13 1 0 11 2 11 7 11 7 9 11 2 15 13 0 0 9 2 9 13 9 9 2
39 11 13 1 0 9 1 11 1 0 9 7 9 9 7 0 9 9 11 11 1 15 13 2 2 11 13 3 1 9 7 13 10 9 2 7 9 3 13 2
25 3 10 9 15 3 13 14 1 9 2 7 7 13 13 1 0 9 7 13 15 1 0 9 2 2
12 11 15 13 9 3 3 13 9 1 9 14 2
22 2 13 15 1 15 3 0 9 2 13 3 1 12 9 2 2 13 0 9 11 11 2
30 9 4 1 11 1 3 0 11 13 0 9 11 2 15 4 1 0 9 1 12 9 2 5 1 9 9 12 9 13 2
13 3 1 9 1 0 9 13 0 9 0 9 11 2
5 1 0 9 0 9
8 9 9 13 1 9 9 1 9
2 11 2
27 9 1 0 9 0 9 15 13 9 11 11 9 9 9 1 9 9 7 3 13 16 3 0 1 9 14 2
48 1 0 9 9 15 13 15 9 1 9 12 9 12 2 11 2 11 2 11 2 11 2 7 9 0 1 12 9 12 2 11 11 2 0 2 11 2 7 12 9 12 2 9 11 2 11 2 2
15 10 9 4 0 9 1 12 0 9 13 1 9 9 11 2
27 0 9 13 0 9 11 2 11 2 0 9 13 2 11 2 11 2 11 2 9 7 11 2 0 2 11 2
26 0 12 9 0 9 4 13 1 9 1 0 9 7 3 1 9 13 15 1 9 12 9 1 0 9 2
5 12 0 9 1 11
2 11 2
42 1 12 0 9 0 9 2 15 9 11 11 13 1 0 9 1 9 1 11 12 2 9 1 11 2 13 14 12 9 2 11 1 11 2 11 1 11 7 11 1 11 2
23 0 9 0 1 9 4 13 0 9 2 16 13 3 13 1 10 9 1 0 9 1 11 2
22 1 9 11 2 11 2 11 7 11 15 1 1 9 10 9 1 0 9 13 3 3 2
22 1 9 11 1 9 0 9 13 7 11 7 1 11 13 13 9 9 9 1 0 9 2
11 0 9 9 11 13 1 12 2 0 9 2
3 11 1 9
2 11 2
23 0 9 7 9 9 1 9 11 11 11 13 13 3 0 9 7 13 1 0 9 1 11 2
37 0 9 0 9 1 11 15 13 10 9 7 9 9 9 2 3 7 13 13 0 0 9 2 11 2 1 9 7 13 15 0 9 3 1 9 12 2
4 11 0 9 11
2 11 2
12 0 9 11 11 13 0 9 0 0 0 9 2
18 9 9 15 1 10 9 13 9 9 1 0 9 1 9 12 1 11 2
24 11 16 0 9 13 11 2 11 7 11 7 1 0 9 13 3 7 0 9 11 7 0 11 2
2 11 9
2 11 2
29 0 0 0 9 2 0 9 2 13 1 9 3 1 9 7 1 12 0 9 4 13 1 11 11 9 7 0 9 2
35 11 15 3 3 13 3 1 12 9 7 9 1 11 11 12 2 12 13 1 9 9 11 0 9 1 9 2 15 1 0 9 13 1 9 2
5 11 13 3 9 9
15 0 9 9 11 11 2 2 9 13 1 0 9 16 9 2
2 11 2
33 0 9 1 12 5 12 9 15 13 16 12 1 0 0 9 0 9 9 9 2 15 15 13 12 2 2 12 2 12 2 1 11 2
35 1 0 0 9 1 11 0 9 1 9 11 2 11 2 11 7 11 13 7 9 12 2 12 13 0 9 1 3 0 9 12 5 12 9 2
51 1 10 9 15 7 0 9 1 11 13 2 16 1 0 9 4 13 3 11 11 2 15 1 11 13 9 1 9 1 12 9 2 7 11 11 2 15 15 15 1 9 1 11 13 1 0 9 1 9 3 2
17 3 15 13 16 0 2 16 1 0 11 13 1 11 0 12 9 2
14 2 15 9 15 13 0 9 2 16 0 9 3 13 2
26 11 11 13 9 3 1 9 9 7 13 2 16 15 15 3 13 2 2 13 11 11 2 0 9 9 2
9 2 9 13 2 16 13 12 9 2
24 13 15 9 0 9 0 9 2 15 13 1 10 0 9 16 9 2 15 15 13 7 1 9 2
31 3 15 1 15 13 13 2 16 13 9 2 7 0 13 0 9 13 15 1 0 9 2 16 1 0 9 3 3 13 2 2
20 11 11 1 0 9 13 2 2 1 0 0 0 9 1 11 13 0 9 0 2
14 13 2 16 15 9 2 3 10 11 2 1 9 13 2
23 13 2 16 1 0 9 7 9 13 15 1 9 2 15 15 1 11 3 13 2 3 13 2
22 3 13 3 0 13 9 2 16 4 15 15 1 9 13 2 16 9 13 3 0 2 2
39 9 9 15 13 1 9 13 2 7 11 11 4 15 13 1 0 2 2 0 9 3 3 13 2 7 1 9 9 13 0 13 2 16 9 13 3 0 9 2
11 13 2 16 1 9 13 0 13 10 9 2
36 11 11 13 0 9 1 9 2 11 11 13 3 0 13 1 0 9 2 11 11 0 9 3 13 7 1 11 11 13 0 2 16 13 13 2 2
38 1 11 2 11 15 3 4 13 13 0 9 1 0 9 2 2 0 9 13 2 16 4 11 13 1 9 1 12 9 2 16 9 9 13 1 12 9 2
20 1 15 15 7 13 1 9 9 2 16 15 13 3 14 0 9 1 9 2 2
19 11 11 15 13 0 9 0 2 2 13 2 16 1 11 12 9 9 13 2
13 13 15 9 2 7 1 9 13 15 9 1 9 2
10 1 9 4 13 1 9 11 11 9 2
14 15 4 15 3 13 2 7 15 15 1 9 3 13 2
37 1 10 9 3 16 11 11 13 10 9 9 2 1 0 9 15 1 9 13 9 1 0 9 7 1 15 15 9 13 13 2 9 2 9 2 2 2
16 1 10 9 4 13 3 0 2 7 13 2 16 15 3 13 2
15 16 15 3 9 13 1 9 2 13 9 2 16 13 2 2
1 3
23 11 11 13 0 9 0 9 1 9 1 9 1 0 11 2 11 2 9 12 7 12 9 2
21 0 13 0 9 11 2 12 7 12 9 2 7 0 11 2 12 7 12 9 2 2
12 11 11 13 13 10 9 1 0 9 1 11 2
8 1 9 9 13 10 0 9 2
3 1 0 9
22 9 11 11 4 9 0 9 11 11 13 0 9 0 9 3 2 16 15 13 11 11 2
9 11 15 1 11 13 16 1 0 9
30 16 13 0 9 11 11 2 12 9 2 1 9 12 1 9 0 11 11 11 2 13 9 9 10 0 9 1 11 9 2
28 13 3 1 15 9 2 16 4 3 13 13 9 9 9 11 11 2 15 15 1 0 12 9 13 1 0 9 2
21 3 13 3 11 0 9 11 2 7 3 13 9 2 16 4 3 10 0 9 13 2
5 2 15 3 14 2
17 13 10 9 16 11 2 7 16 3 13 13 0 9 9 16 15 2
25 3 1 0 9 2 16 4 1 11 13 12 2 12 2 4 13 1 0 12 1 9 14 12 9 2
19 3 13 3 3 7 3 15 13 7 15 2 16 15 11 13 0 9 13 2
20 13 15 1 15 3 0 9 2 7 1 0 9 3 13 3 9 3 7 3 2
30 15 13 13 9 7 15 3 13 1 15 2 16 11 13 1 9 2 13 12 9 7 9 13 3 2 2 13 11 11 2
28 1 0 9 13 11 0 9 7 13 15 2 16 13 9 11 11 1 9 12 2 3 11 9 13 0 12 9 2
18 9 9 15 7 1 9 13 1 9 12 2 12 1 11 1 9 12 2
20 2 15 15 13 13 0 2 16 4 13 3 1 11 2 15 13 1 0 9 2
16 15 7 13 3 0 9 7 13 15 15 13 15 10 9 2 2
25 0 9 0 9 11 2 15 4 1 1 0 9 13 1 12 9 1 12 2 13 11 1 0 9 2
13 2 15 13 3 3 2 16 15 15 13 13 13 2
14 0 9 13 0 9 2 1 9 4 13 0 0 9 2
30 3 15 15 1 0 12 9 13 16 1 0 9 2 3 15 1 15 13 12 9 7 0 9 1 15 13 3 3 2 2
28 1 9 10 9 11 13 2 16 10 9 13 13 15 9 2 1 15 4 13 13 2 16 13 0 9 1 9 2
21 2 3 9 1 11 13 2 16 3 15 15 15 13 2 7 15 10 9 3 13 2
10 13 4 15 15 1 15 3 13 9 2
21 13 2 16 16 4 12 12 9 3 13 7 13 1 0 9 2 13 13 9 0 2
3 7 3 2
19 15 14 3 14 2 2 13 3 11 2 15 3 13 12 9 7 12 9 2
15 13 15 0 9 11 7 11 7 3 0 9 11 7 11 2
7 2 10 9 13 3 0 2
16 3 3 15 13 1 11 3 3 16 3 1 12 7 12 9 2
17 13 3 11 2 15 15 1 15 13 2 9 13 0 7 9 0 2
14 1 10 9 15 13 11 2 15 13 12 9 2 0 2
16 13 15 3 14 12 9 7 1 0 9 15 3 13 14 9 2
9 7 1 12 2 9 15 13 9 2
24 13 15 3 1 15 2 15 13 7 13 1 9 12 9 2 1 15 15 15 13 13 3 13 2
11 1 11 15 3 13 13 2 2 13 11 2
40 13 15 7 1 9 2 16 15 9 2 3 3 13 2 11 2 11 2 11 2 2 13 10 9 2 2 13 2 13 2 15 13 14 14 10 9 2 2 2 2
19 0 9 11 11 11 2 11 2 1 9 0 9 9 11 11 2 11 2 13
4 11 13 11 11
8 9 13 1 0 7 0 9 9
3 0 11 2
27 0 0 9 11 11 11 13 10 9 1 9 0 9 1 11 2 12 2 9 2 12 2 9 1 11 2 2
8 13 15 3 0 9 11 11 2
6 2 13 15 15 9 2
34 1 12 2 9 4 13 13 1 12 0 9 1 9 1 0 0 2 7 3 3 15 15 1 11 11 1 11 13 13 2 2 13 11 2
15 0 9 9 0 9 13 0 9 0 9 11 2 0 9 2
17 1 9 0 0 0 4 0 11 11 3 13 7 9 13 0 9 2
27 11 3 3 13 9 1 11 1 9 3 2 16 1 15 12 1 9 13 2 16 4 13 3 1 10 9 2
8 2 11 15 13 9 0 9 2
13 10 9 13 3 3 7 3 15 3 13 3 13 2
13 7 15 13 13 9 10 9 2 2 13 0 9 2
2 0 9
2 11 2
33 3 0 9 0 0 9 3 13 9 12 2 9 0 9 9 9 12 9 1 11 0 9 7 11 11 11 12 2 12 1 9 0 2
11 9 0 9 15 1 9 12 2 9 13 2
5 11 3 13 0 9
2 11 2
19 11 11 2 0 0 9 7 9 11 0 2 13 1 10 9 3 0 9 2
27 1 0 9 1 9 13 1 0 9 1 9 1 9 2 1 9 15 3 4 13 1 0 9 0 0 9 2
35 9 13 0 9 1 0 9 1 0 11 9 9 2 3 0 0 9 13 9 9 3 2 16 1 9 13 1 9 7 13 15 9 0 9 2
5 1 11 13 0 9
4 11 1 11 2
17 12 0 0 9 4 13 1 9 1 9 1 9 1 11 1 11 2
6 3 15 13 0 9 2
27 12 9 1 9 12 7 12 12 9 4 13 1 9 0 9 2 15 13 1 0 9 1 9 1 9 11 2
18 12 1 0 13 3 7 0 13 1 0 9 2 16 15 9 3 13 2
17 1 9 3 0 12 9 13 13 0 9 3 2 16 4 13 9 2
17 0 9 13 1 9 1 11 1 11 7 11 1 9 11 1 11 2
11 12 1 15 13 1 15 9 11 1 11 2
11 3 12 9 13 1 0 9 1 0 9 2
14 9 3 13 2 16 15 1 9 13 13 16 0 9 2
6 0 9 3 13 0 9
5 9 9 1 0 9
10 2 9 3 13 0 9 2 2 13 11
12 1 0 0 9 13 1 0 9 0 0 9 2
12 16 9 13 10 9 2 3 3 14 1 9 2
14 2 9 1 9 3 13 2 2 13 0 9 11 11 2
31 2 15 13 13 9 1 0 11 11 2 3 15 1 9 13 0 9 2 7 13 15 15 3 2 2 13 9 11 9 11 2
27 11 11 2 9 9 7 9 0 9 11 2 13 1 10 9 3 0 2 2 9 9 3 13 0 9 0 9
17 16 3 1 11 13 3 14 12 12 9 2 13 15 3 0 2 2
19 11 11 2 9 11 11 2 3 13 0 9 9 1 9 0 0 9 9 2
19 2 13 15 9 1 0 0 9 2 13 2 14 9 2 15 3 13 2 2
17 1 9 1 0 9 9 7 9 13 3 3 9 9 7 9 9 2
15 2 10 9 15 13 3 1 0 9 7 3 10 9 13 2
10 1 9 15 7 13 2 2 13 11 2
17 0 9 1 9 9 2 1 12 12 9 2 13 14 14 0 9 2
17 2 9 13 0 2 3 16 15 13 9 7 13 0 3 13 9 2
10 13 7 0 9 2 2 13 0 9 2
36 3 3 1 15 13 3 11 2 15 3 1 0 0 9 13 1 0 9 10 9 2 7 1 9 9 4 13 1 9 13 0 2 15 3 13 2
41 0 9 1 0 9 13 7 11 2 16 0 9 3 13 2 3 13 1 0 9 2 16 3 9 0 9 9 1 0 9 9 2 3 13 11 12 2 12 2 2 2
15 0 0 9 2 16 3 0 2 13 1 0 9 0 11 2
18 16 15 9 1 11 11 3 14 13 2 13 1 0 9 12 12 9 2
39 2 13 15 15 13 1 11 1 9 9 2 3 13 0 9 2 0 2 9 2 9 2 2 7 3 4 13 10 9 1 9 9 2 2 13 15 9 11 2
13 3 15 7 0 9 0 9 1 9 1 9 13 2
13 2 16 1 15 13 15 13 2 0 9 15 13 2
11 13 15 3 12 9 2 2 13 11 11 2
23 9 13 14 12 2 1 9 9 13 9 9 13 0 9 16 3 7 13 1 0 0 9 2
10 2 7 15 9 13 2 7 13 3 2
21 16 7 9 13 3 15 2 1 9 13 9 0 2 16 13 9 2 2 13 11 2
10 1 0 9 9 13 9 9 1 9 2
15 2 9 15 4 13 3 13 2 7 0 9 13 3 3 2
9 3 15 3 13 1 9 0 9 2
25 3 3 13 3 12 9 2 15 15 4 13 13 7 1 15 0 0 13 2 7 0 2 2 2 2
15 0 9 11 11 13 1 0 9 0 2 3 3 0 9 2
17 0 9 11 11 2 3 2 1 15 13 13 3 14 1 0 9 2
5 0 9 12 2 9
3 0 0 9
5 11 3 13 0 9
14 0 9 0 9 13 1 9 9 11 9 11 7 9 11
18 9 11 13 0 9 1 9 0 9 2 7 7 11 3 13 0 9 2
15 1 10 9 13 1 9 11 9 9 7 0 9 0 9 2
24 1 9 9 14 15 13 3 0 11 2 0 9 9 13 9 3 1 11 1 11 7 9 11 2
10 11 11 2 9 11 11 7 9 11 2
14 12 2 11 15 13 3 0 2 7 13 4 9 11 2
7 1 0 9 13 0 15 2
9 12 2 0 13 2 16 14 15 2
4 12 2 15 2
2 12 2
3 10 11 2
6 11 0 2 9 11 2
11 12 2 3 15 1 9 11 1 11 13 2
17 11 3 13 1 3 0 9 16 11 2 7 1 9 13 0 9 2
8 16 15 13 11 2 13 9 2
4 12 2 13 2
21 11 7 11 15 13 2 0 9 9 9 1 11 13 2 16 7 15 14 2 2 2
13 12 2 16 15 9 3 13 0 2 7 0 9 2
17 15 15 3 13 1 0 9 2 3 15 9 3 2 13 16 13 2
2 12 2
2 11 2
7 11 11 2 9 9 9 2
15 12 2 9 4 13 11 2 16 14 3 2 3 1 9 2
19 16 4 13 1 3 0 9 11 2 13 4 15 0 9 7 1 0 9 2
20 11 13 0 9 2 3 3 13 1 9 1 9 11 2 13 0 9 1 11 2
14 12 2 9 15 13 2 7 16 1 15 13 3 13 2
5 0 9 13 11 2
16 12 2 15 13 1 9 2 3 9 9 13 0 1 0 9 2
4 15 3 13 2
20 12 2 0 9 4 13 13 3 11 2 0 13 11 7 9 4 13 7 11 2
9 11 11 2 9 11 1 12 9 2
10 12 2 13 15 1 11 7 11 11 2
12 11 4 13 13 2 16 15 3 13 15 9 2
9 11 13 3 13 2 16 15 13 2
8 11 13 1 9 3 0 9 2
14 12 2 13 12 9 2 11 2 11 2 11 7 11 2
8 9 13 11 2 15 3 14 2
15 11 13 3 1 9 7 1 15 0 9 7 13 9 13 2
11 3 16 11 13 0 9 2 13 1 9 2
23 3 13 9 11 2 1 0 9 2 16 13 9 2 13 9 9 7 15 4 1 11 13 2
21 12 2 1 10 9 13 0 9 2 11 13 0 0 9 2 9 13 1 9 9 2
14 12 2 11 1 9 2 16 15 9 11 4 13 3 2
7 11 11 2 9 11 11 2
11 12 2 11 2 16 13 9 0 15 9 2
7 12 3 13 14 1 9 2
9 12 2 3 13 2 16 14 15 2
10 13 15 14 1 11 2 11 7 11 2
10 12 2 9 9 1 15 9 1 11 2
12 3 15 13 9 1 10 9 2 15 15 13 2
9 13 15 15 9 7 9 1 9 2
13 12 2 13 4 15 13 10 11 2 3 7 11 2
7 11 11 2 9 11 11 2
11 12 2 1 10 13 9 14 0 12 9 2
16 3 15 13 3 0 11 2 7 1 12 9 15 13 13 3 2
17 11 13 1 9 13 14 1 9 2 16 13 1 11 7 1 15 2
13 12 2 12 9 3 4 13 2 7 15 15 13 2
19 12 2 16 9 13 14 16 9 1 9 7 7 3 2 13 15 1 0 2
11 12 2 0 13 2 16 4 15 10 9 2
7 11 11 2 9 9 11 2
17 12 2 7 15 15 4 13 2 7 13 11 2 16 13 0 9 2
11 12 2 13 15 1 11 2 11 7 11 2
17 3 3 13 1 15 7 11 2 7 1 10 9 13 3 13 3 2
2 12 2
2 15 2
2 12 2
13 11 2 15 4 13 13 3 0 9 1 0 9 2
7 11 11 2 9 11 11 2
4 12 2 11 2
9 13 0 9 7 14 7 0 9 2
4 12 2 13 2
8 12 2 13 15 9 1 9 2
20 15 15 1 15 13 2 15 1 15 13 7 15 4 13 1 9 13 2 2 2
16 12 2 13 4 15 15 10 12 9 2 15 4 1 9 13 2
8 11 11 2 0 9 11 11 2
13 12 2 11 2 13 0 0 9 7 13 0 9 2
2 12 2
2 11 2
16 1 0 9 13 9 2 10 9 2 15 13 3 1 9 9 2
11 11 15 13 3 2 7 14 1 0 9 2
6 12 2 9 13 0 2
13 12 2 11 13 2 16 13 1 10 9 0 9 2
16 11 11 2 9 9 11 2 9 2 9 2 9 2 0 2 2
2 12 2
5 9 13 15 0 2
8 3 3 4 15 15 3 13 2
2 12 2
4 13 15 0 2
11 0 4 15 13 2 15 4 13 0 9 2
2 12 2
13 9 0 9 2 9 1 9 1 9 13 0 9 2
2 12 2
3 3 9 2
10 0 9 10 9 11 7 4 15 13 2
7 11 11 2 9 11 11 2
14 12 2 13 15 1 11 7 11 2 7 13 0 9 2
2 12 2
13 3 13 2 9 2 3 2 9 1 9 13 0 2
7 4 13 1 0 12 9 2
2 12 2
2 15 2
2 12 2
5 9 1 15 13 2
11 3 9 11 4 15 1 0 9 13 13 2
7 11 11 2 9 11 11 2
23 12 2 13 2 16 11 2 7 1 0 9 13 11 2 15 13 0 9 16 1 12 9 2
2 12 2
7 1 9 9 13 15 0 2
17 9 15 13 13 1 12 2 9 7 13 2 15 1 9 13 9 2
2 12 2
28 16 15 0 9 13 9 11 2 9 11 2 9 2 9 2 2 9 11 7 16 15 13 13 10 9 1 9 2
2 12 2
3 3 11 2
8 11 11 2 0 9 9 11 2
10 12 2 13 15 1 11 7 11 11 2
18 11 13 0 9 2 11 3 0 9 2 16 13 1 11 7 11 3 2
16 3 1 15 13 2 3 15 11 7 11 13 1 9 1 11 2
2 12 2
10 1 9 3 9 13 9 9 12 11 2
8 1 11 13 2 3 13 9 2
7 0 0 13 7 3 11 2
7 9 1 0 9 0 9 2
5 0 11 7 11 2
21 11 13 1 9 7 9 9 9 2 15 13 0 9 2 11 3 16 0 9 3 2
7 11 11 2 9 11 11 2
15 0 0 9 13 11 2 7 7 11 3 13 10 0 9 2
2 12 2
14 9 15 13 2 3 0 9 13 11 2 11 7 11 2
2 12 2
10 13 15 9 1 0 9 7 0 9 2
2 12 2
15 13 0 9 2 7 13 0 2 16 10 13 15 1 15 2
7 11 11 2 9 11 11 2
7 12 2 11 13 0 9 2
14 1 9 15 3 13 2 9 9 13 3 0 9 3 2
14 13 15 2 16 1 9 13 15 7 1 9 15 13 2
2 12 2
4 0 3 13 2
2 12 2
8 9 9 13 9 11 1 11 2
2 12 2
9 10 0 9 13 3 10 9 11 2
7 11 11 2 9 9 9 2
20 12 2 13 15 1 11 7 11 2 1 9 13 7 11 7 14 1 0 11 2
2 12 2
3 12 0 2
2 12 2
5 9 1 0 9 2
2 12 2
7 9 11 7 11 1 11 2
9 16 15 14 0 9 13 1 9 2
7 11 11 2 9 11 11 2
8 12 2 3 13 2 16 15 2
2 12 2
6 13 2 9 13 0 2
2 12 2
11 3 10 9 1 9 7 1 9 3 13 2
2 12 2
6 11 2 11 2 11 2
7 11 11 2 9 11 11 2
11 12 2 0 13 2 16 9 13 1 11 2
14 0 9 13 11 7 11 2 7 1 9 13 7 11 2
9 11 13 9 2 15 15 4 13 2
9 13 9 7 13 0 9 15 13 2
2 12 2
11 13 13 3 9 2 15 13 1 9 9 2
13 13 15 13 15 2 7 13 2 16 15 13 0 2
2 12 2
10 15 9 1 9 7 9 1 0 9 2
2 12 2
15 1 10 9 4 13 0 2 16 4 10 9 13 3 3 2
22 1 10 9 13 9 2 16 15 9 13 1 9 2 13 2 16 15 13 1 0 9 2
8 11 11 2 9 11 0 11 2
16 12 2 15 13 0 2 13 15 1 9 11 2 11 2 11 2
17 11 7 11 1 15 13 9 1 9 2 7 11 3 13 0 9 2
2 12 2
3 0 13 2
14 7 15 3 13 13 7 13 4 3 15 1 9 13 2
2 12 2
5 9 11 1 11 2
2 12 2
14 15 15 13 9 1 11 2 15 13 9 1 0 9 2
6 11 11 2 9 11 2
21 12 2 11 13 0 0 9 7 0 9 2 16 16 15 13 9 2 13 4 13 2
2 12 2
5 13 0 9 9 2
2 12 2
6 0 9 1 9 9 2
2 12 2
11 11 2 15 15 3 13 7 1 0 9 2
7 11 11 2 9 9 11 2
11 12 2 12 1 9 11 2 11 2 11 2
2 12 2
4 15 15 13 2
2 12 2
2 15 2
2 12 2
12 10 9 13 2 16 4 15 13 11 1 9 2
8 11 11 2 9 0 9 11 2
17 12 2 13 4 15 13 11 2 16 16 0 13 13 1 9 9 2
4 13 7 11 2
2 12 2
14 13 2 15 13 2 1 10 9 13 9 1 0 9 2
2 12 2
2 15 2
2 12 2
18 1 0 11 15 3 3 2 13 16 3 13 2 16 4 15 13 13 2
5 15 13 3 9 2
4 11 13 0 9
17 0 9 11 13 1 9 11 2 15 15 13 13 1 9 0 9 2
31 1 0 9 1 9 0 2 9 1 0 9 2 13 9 0 9 9 9 2 13 1 9 1 9 9 7 3 15 13 9 2
23 9 11 15 1 11 13 0 0 9 1 12 9 2 1 9 12 3 13 0 9 11 2 2
14 1 9 15 13 14 12 9 2 15 13 3 12 9 2
23 0 9 1 9 13 10 9 2 9 7 9 9 1 9 2 1 15 13 14 1 10 9 2
29 0 9 3 13 9 2 0 2 9 9 14 3 2 1 15 13 3 0 9 10 9 2 16 13 11 7 11 11 2
2 9 9
1 9
16 9 2 3 0 13 9 0 1 0 9 0 9 2 0 9 2
22 3 1 9 10 9 13 9 0 0 0 9 2 15 9 13 3 9 0 0 0 9 2
25 0 13 7 7 15 2 3 1 0 9 9 3 13 0 9 0 9 11 11 2 15 9 13 11 2
20 0 0 0 9 0 0 9 13 0 0 0 9 0 2 3 0 7 0 9 2
20 3 0 9 13 1 11 9 3 3 13 3 0 9 1 9 2 0 1 11 2
31 7 3 15 0 9 1 15 13 1 9 9 0 9 2 15 0 2 7 1 0 7 0 9 0 9 1 0 9 13 3 2
13 3 15 13 2 16 0 9 0 13 0 0 9 2
10 0 9 13 1 9 0 12 0 9 2
27 15 13 3 0 7 16 13 3 13 2 3 2 13 2 7 1 0 9 13 2 10 0 9 13 0 9 2
31 9 1 9 1 9 9 10 0 9 1 9 2 9 7 2 0 9 0 9 2 3 13 0 7 0 0 9 7 10 9 2
41 9 2 9 2 0 9 7 0 9 1 0 9 1 0 0 3 0 9 9 12 2 2 13 9 9 7 9 2 2 3 13 14 3 0 0 9 1 0 0 9 2
16 11 11 0 9 2 0 0 9 2 11 9 2 9 11 12 2
5 0 9 9 0 9
23 9 1 9 7 9 11 11 2 12 2 12 2 13 0 9 11 2 11 2 11 1 11 2
16 13 3 9 9 1 9 10 0 0 9 2 9 7 0 9 2
18 10 9 2 13 1 12 2 9 2 4 13 1 9 0 0 9 11 2
42 9 11 11 13 13 1 9 7 0 9 0 9 1 11 1 11 2 1 9 1 0 9 2 1 9 0 2 7 1 9 9 3 0 2 9 0 1 0 7 0 9 2
14 1 9 0 9 13 2 3 13 1 11 7 1 11 2
20 0 9 11 2 11 2 11 13 3 1 12 9 0 9 1 0 9 7 9 2
23 13 1 10 9 3 9 2 7 15 1 0 1 9 1 9 11 11 7 11 11 1 11 2
33 10 9 3 1 9 9 13 0 9 0 9 1 9 11 2 9 9 0 9 0 0 9 1 0 2 11 1 11 2 11 2 11 2
13 13 1 9 9 1 0 0 9 9 2 12 2 2
9 3 3 9 13 3 2 12 2 2
19 0 9 1 11 11 4 13 12 2 9 7 9 1 15 13 9 11 11 2
3 11 13 9
14 0 9 9 9 13 3 12 2 9 0 0 9 11 2
23 12 1 0 9 4 13 0 9 7 9 11 11 1 0 9 9 2 15 13 9 0 9 2
36 0 9 1 0 0 9 13 0 9 9 2 0 2 9 2 9 11 11 2 0 9 1 0 0 9 2 15 15 1 9 10 9 13 13 9 2
39 0 9 9 2 0 9 2 7 0 9 11 2 4 2 1 9 1 0 9 11 11 2 13 0 9 9 2 9 2 2 15 1 11 13 0 9 11 11 2
28 0 9 1 0 9 13 11 11 1 0 2 16 3 3 0 9 1 9 9 2 1 9 2 11 2 11 2 2
32 0 9 1 0 0 9 13 11 11 2 1 9 1 0 9 10 9 2 7 0 9 11 11 2 1 9 1 9 0 9 2 2
28 1 0 0 9 15 13 0 2 0 9 2 9 2 11 11 2 7 0 9 1 9 2 9 2 11 11 2 2
16 9 9 2 15 3 13 11 9 11 1 11 2 13 3 3 2
21 1 9 1 0 0 9 13 0 9 9 2 3 1 9 0 9 7 9 1 9 2
7 9 0 9 15 13 9 9
23 1 9 9 7 9 13 1 11 2 7 3 3 7 1 11 2 0 9 9 9 0 9 2
28 9 9 13 13 9 1 0 0 9 2 15 13 3 3 9 1 9 1 0 9 2 0 3 9 0 7 0 2
35 1 0 9 1 9 2 1 12 2 1 12 2 9 2 7 1 9 0 0 9 2 1 12 2 1 12 2 9 2 4 13 12 0 9 2
34 1 9 15 13 3 9 9 2 14 9 0 9 11 2 11 2 9 0 9 0 9 11 2 11 7 9 1 9 0 9 11 2 11 2
25 10 9 4 1 9 13 0 9 9 11 2 0 0 9 9 2 9 9 11 11 7 0 9 11 2
4 9 13 1 11
25 1 0 9 7 0 0 9 13 0 0 9 0 0 0 0 9 2 15 1 0 12 9 13 11 2
26 1 9 1 9 15 13 3 3 1 0 0 9 7 0 7 15 0 9 2 11 11 2 11 11 2 2
40 9 13 1 12 9 2 12 1 15 13 0 2 1 0 9 1 11 7 11 1 11 2 11 7 11 14 1 9 0 2 0 2 11 2 11 11 7 11 11 2
29 1 9 1 11 15 3 0 0 9 13 3 9 1 0 11 2 1 11 2 11 2 11 2 11 2 11 7 11 2
5 15 2 3 2 3
21 9 9 11 11 4 3 13 1 9 9 9 1 11 2 13 1 12 2 9 2 2
29 10 9 0 9 2 0 11 2 13 9 7 9 11 9 3 1 12 9 1 9 0 11 2 0 12 2 11 12 2
7 9 9 13 9 11 11 2
21 9 9 7 9 11 11 4 3 2 12 2 13 1 9 9 1 0 9 1 11 2
19 9 9 15 13 9 2 15 13 1 9 1 0 0 9 1 12 2 9 2
2 0 9
1 9
26 9 2 1 0 9 9 13 15 0 9 9 0 9 11 1 0 9 0 9 9 11 11 2 12 2 2
17 13 15 1 15 3 2 16 1 0 9 13 9 0 7 0 9 2
11 15 9 13 10 9 2 0 3 1 9 2
14 9 13 3 1 9 2 13 1 9 7 13 1 9 2
5 13 9 10 9 2
8 11 11 13 1 15 0 9 2
34 16 13 1 3 16 12 9 1 9 2 3 13 1 11 2 2 13 4 9 13 10 9 1 0 9 7 1 0 10 9 7 1 11 2
12 3 13 10 9 9 2 15 7 13 13 9 2
16 11 13 1 9 0 7 0 9 2 13 15 3 7 0 9 2
16 9 7 9 10 0 2 7 3 0 2 9 13 9 0 9 2
19 0 9 2 7 15 13 9 7 9 2 15 13 0 9 2 7 0 9 2
13 13 1 0 9 2 1 9 0 9 1 0 9 2
32 1 0 2 9 2 2 2 9 2 2 2 9 2 7 2 9 2 15 13 0 9 2 15 15 13 1 0 9 1 0 9 2
16 9 13 13 9 2 3 16 9 15 2 1 9 1 10 9 2
8 1 10 9 15 13 3 13 2
17 9 13 3 13 15 2 7 16 4 15 13 10 9 13 1 9 2
9 11 15 15 1 15 9 13 3 2
19 10 9 13 0 9 2 7 7 9 2 15 4 15 13 0 9 10 9 2
26 13 1 2 9 2 0 9 2 1 10 9 7 9 2 7 3 1 9 2 15 13 1 15 3 0 2
22 9 0 0 9 13 14 9 9 10 9 2 7 3 9 9 2 9 9 1 0 9 2
18 0 0 9 2 0 1 0 9 2 13 3 2 7 3 10 9 13 2
8 0 9 9 13 1 9 9 2
18 9 2 9 2 9 1 9 2 1 9 9 2 2 15 13 0 9 2
6 0 9 9 7 9 2
4 9 15 13 2
12 14 1 9 9 2 7 1 9 1 9 9 2
11 13 1 9 2 3 10 9 7 13 0 2
34 3 0 9 2 16 4 9 1 9 0 9 13 2 0 9 2 9 7 3 9 2 13 9 9 2 9 2 9 2 3 9 3 13 2
6 13 9 0 0 9 2
12 0 9 13 10 9 2 0 9 13 10 9 2
18 1 11 11 4 13 3 1 11 2 1 10 9 0 9 7 0 9 2
13 1 9 2 15 15 13 1 0 9 9 1 9 2
26 2 1 15 13 9 3 3 15 2 15 13 1 9 0 9 2 2 13 9 1 9 1 11 2 11 2
26 1 0 9 9 2 1 15 9 13 3 15 2 15 13 1 10 9 2 13 0 0 9 3 16 0 2
17 13 9 3 15 13 9 0 7 13 2 16 13 15 16 0 9 2
5 11 11 11 11 2
10 9 0 2 9 2 11 2 0 9 2
8 12 2 9 2 12 2 9 2
20 9 2 15 13 9 2 7 15 10 9 2 9 2 13 1 0 9 15 0 2
20 4 2 14 7 15 13 1 15 13 2 13 15 9 7 13 7 9 0 9 2
7 13 15 3 13 2 2 2
17 2 11 12 2 12 2 12 2 11 11 1 10 9 3 13 9 2
16 13 15 3 7 2 16 9 13 2 0 2 1 9 0 9 2
12 15 9 9 4 13 7 13 1 0 0 9 2
27 13 1 0 0 9 2 15 7 13 0 9 1 9 12 2 3 4 9 9 1 15 15 13 1 9 9 2
29 9 13 1 0 9 1 9 1 9 0 9 2 1 15 15 3 13 13 1 9 1 9 7 13 1 15 0 9 2
6 9 1 9 13 9 2
23 3 9 2 15 13 1 0 9 1 9 2 0 0 9 2 2 4 13 0 9 7 9 2
18 0 9 2 9 2 7 1 9 13 13 2 15 13 1 9 9 9 2
11 13 15 3 13 0 9 9 9 9 9 2
14 9 2 9 2 9 13 13 2 13 9 1 0 9 2
27 16 3 9 9 1 0 9 13 0 2 0 9 2 2 3 9 2 3 13 15 3 14 9 2 3 9 2
25 9 13 10 0 9 2 9 13 3 1 0 9 2 1 15 13 9 9 9 2 7 3 0 9 2
48 9 3 13 10 2 0 9 2 2 16 13 0 9 0 2 1 9 2 2 9 9 9 7 9 2 9 1 9 9 1 0 9 1 9 2 9 9 1 0 7 0 1 9 1 9 9 9 2
19 1 9 12 13 0 9 0 0 9 0 9 2 1 15 13 9 0 9 2
8 3 13 15 1 9 0 9 2
6 9 13 9 1 0 9
40 1 9 9 9 1 0 9 4 9 7 9 13 13 1 9 2 16 7 15 13 0 7 16 15 3 13 1 9 2 1 15 15 3 13 15 7 9 10 9 2
12 16 4 13 2 13 4 1 10 9 9 9 2
10 3 3 7 13 10 9 9 1 15 2
34 9 10 0 9 15 13 1 15 2 1 10 0 7 0 0 9 15 15 13 13 2 7 1 15 2 16 15 13 1 0 1 10 0 2
34 1 0 9 13 13 2 16 13 14 3 9 2 16 4 4 9 2 15 0 9 3 13 7 13 9 7 9 2 13 1 0 0 9 2
29 1 15 15 13 3 2 0 2 16 15 2 16 9 13 9 2 13 1 15 2 16 4 4 3 3 7 3 13 2
9 0 9 13 0 9 10 0 9 2
34 1 9 2 3 13 2 16 10 9 3 1 9 13 13 2 3 13 3 0 9 1 9 2 4 15 13 9 2 16 9 15 15 13 2
19 3 2 16 15 2 15 13 1 0 9 7 13 0 9 2 13 3 3 2
31 13 7 2 16 9 13 13 2 16 12 9 2 3 9 0 16 0 9 2 4 13 9 2 15 4 13 1 0 9 9 2
17 3 15 15 4 13 13 12 9 3 2 1 9 9 7 0 9 2
14 10 9 13 1 15 2 16 3 0 9 13 1 9 2
35 16 0 7 0 9 10 9 13 3 9 3 2 1 15 2 16 9 10 0 9 1 10 3 0 9 3 13 1 0 0 9 1 0 9 2
21 16 3 13 2 16 1 9 3 12 9 13 9 7 9 2 13 15 1 15 3 2
13 3 13 0 2 16 3 15 13 3 1 9 13 2
42 13 2 16 16 10 9 7 9 13 1 0 0 9 1 0 9 2 13 0 2 16 0 9 7 9 13 3 10 0 9 1 0 9 1 0 9 2 0 9 7 9 2
11 7 3 3 15 7 15 13 3 3 12 2
18 3 4 13 13 1 10 9 2 15 4 15 13 3 13 7 3 13 2
9 3 3 15 1 10 9 13 13 2
19 13 2 16 4 9 13 7 3 10 9 2 7 15 15 13 1 9 9 2
7 9 1 9 13 0 9 2
6 1 15 13 0 9 2
32 16 9 1 3 0 9 2 0 0 9 1 0 9 1 9 9 13 2 3 15 13 9 1 9 2 11 12 2 12 2 2 2
13 0 9 1 11 15 13 1 9 1 9 9 9 2
20 3 14 7 2 16 13 9 13 1 9 2 3 4 10 9 13 9 7 9 2
12 1 10 9 0 9 11 13 0 9 1 9 2
12 10 9 2 15 13 9 2 3 1 9 13 2
8 3 15 7 13 10 0 9 2
12 9 0 9 2 15 2 13 9 1 10 9 2
15 13 3 3 3 1 9 2 16 13 10 0 9 3 0 2
20 13 2 16 13 0 2 16 4 9 3 13 9 9 2 15 13 7 10 9 2
9 9 9 9 9 13 1 3 0 2
12 13 15 2 16 13 0 9 9 13 9 9 2
10 13 2 16 4 0 9 13 13 0 2
10 0 9 9 11 15 1 10 9 13 2
8 11 13 1 9 1 9 9 2
27 1 15 2 10 9 2 11 13 3 15 2 16 15 1 9 9 0 0 9 3 13 3 13 1 10 9 2
16 10 10 0 9 13 0 0 0 9 2 16 3 0 7 0 2
61 1 11 13 0 9 2 0 1 15 2 9 1 9 7 9 9 2 3 14 0 2 1 9 9 3 14 9 9 2 16 9 9 1 0 9 2 7 1 9 0 9 1 9 7 0 9 1 9 2 16 4 0 9 1 0 9 13 1 11 9 2
5 1 3 9 3 9
36 1 9 0 9 0 9 9 9 4 15 13 13 1 0 9 0 2 0 9 0 9 2 13 2 13 2 7 13 2 11 12 2 12 2 2 2
67 3 1 0 9 13 3 10 9 0 9 2 10 9 2 0 2 0 2 9 2 15 3 13 7 3 13 0 0 9 2 4 14 13 0 2 9 2 2 7 13 3 0 9 0 9 2 15 13 13 1 9 9 1 9 14 12 5 0 9 1 12 5 1 9 2 2 2
36 3 13 9 1 9 9 2 1 9 0 9 2 2 15 3 13 3 16 10 2 0 2 9 2 7 15 14 7 2 16 13 1 9 0 9 2
9 1 9 13 13 1 9 7 3 9
12 0 9 9 7 9 0 9 13 1 0 9 2
15 9 15 7 3 3 3 13 2 16 7 13 1 0 11 2
17 13 15 3 3 3 2 1 11 1 0 9 11 0 12 9 9 2
4 3 1 11 2
17 13 15 1 0 9 3 0 9 11 1 11 13 0 3 1 9 2
13 7 9 3 2 1 9 11 2 3 1 0 9 2
4 1 9 3 14
14 0 9 11 13 1 0 0 9 2 0 9 0 9 2
6 13 0 9 1 9 2
16 1 11 13 9 1 0 0 9 14 1 9 12 9 1 9 2
21 3 15 0 0 9 13 1 0 0 9 1 12 9 3 2 14 1 9 0 9 2
23 1 9 12 9 15 1 9 13 12 1 0 0 9 7 13 13 1 11 7 1 0 9 2
8 9 15 7 16 0 9 13 2
8 1 9 4 15 13 3 13 2
5 3 3 1 11 2
11 11 13 1 9 0 0 9 1 9 12 2
15 13 3 2 7 15 13 9 0 9 1 0 7 0 9 2
19 3 15 3 13 9 0 9 7 1 9 12 15 3 13 9 1 9 9 2
8 0 9 13 0 9 3 0 2
14 3 2 0 0 9 15 1 11 13 3 1 9 9 2
18 1 0 0 9 13 11 14 12 1 15 12 11 2 15 13 1 11 2
2 9 2
7 9 3 13 1 0 9 2
13 9 1 0 9 2 9 1 0 0 9 2 2 2
13 1 11 13 7 0 0 9 7 0 9 16 9 2
25 9 7 3 13 0 9 9 7 9 2 15 14 1 11 13 1 9 13 1 12 9 3 0 9 2
16 1 10 9 3 13 3 16 1 0 9 1 11 2 3 3 2
8 3 1 11 13 3 0 9 2
20 1 0 9 1 0 9 13 12 9 1 9 1 12 9 2 9 0 13 0 2
35 9 0 9 2 0 0 0 9 2 13 2 12 9 1 9 2 0 9 2 9 0 9 7 9 1 0 9 2 15 15 1 0 12 9 2
20 13 15 3 3 2 13 2 14 2 16 14 0 0 9 13 1 9 12 9 2
18 13 9 7 1 9 7 1 9 9 2 0 1 9 9 1 0 9 2
3 9 3 13
27 1 0 2 0 2 9 15 0 0 9 13 13 0 9 2 15 13 0 1 0 9 7 1 0 9 9 2
23 9 13 0 9 7 9 9 2 13 9 2 13 15 1 9 9 2 3 0 7 0 9 2
11 13 0 9 7 9 9 2 0 0 9 2
10 0 9 13 1 0 9 9 7 9 2
10 9 1 10 9 15 13 1 9 9 2
18 1 11 3 13 1 12 9 9 0 0 9 1 9 12 9 1 9 2
25 3 2 1 9 12 2 3 3 4 13 1 9 0 0 9 2 15 1 0 9 13 0 0 9 2
10 1 9 9 13 7 3 14 3 13 2
29 12 7 0 0 0 9 13 3 0 9 9 1 9 2 3 10 0 9 2 7 9 0 9 1 9 9 0 9 2
7 7 0 9 3 13 0 2
15 10 9 13 10 9 2 3 9 2 0 9 2 3 9 2
25 1 11 3 13 7 3 9 2 12 2 9 2 3 1 0 2 11 2 13 0 9 11 1 9 2
15 0 9 1 9 1 11 13 0 9 0 0 9 0 11 2
3 9 9 11
10 13 9 13 2 15 13 15 2 2 2
21 0 9 4 15 13 13 3 0 9 2 13 11 11 2 15 1 9 13 1 0 11
14 1 9 12 3 4 7 1 9 1 10 9 13 3 2
8 3 4 0 9 13 15 3 2
23 12 2 9 4 1 9 1 9 13 1 0 9 14 1 9 2 3 15 3 13 0 9 2
19 13 4 7 3 2 3 1 0 9 1 11 14 1 9 10 9 1 11 2
23 0 9 9 4 13 2 3 2 2 16 15 2 9 2 11 2 11 7 0 2 3 13 2
29 1 9 12 2 1 9 2 3 1 9 0 9 13 11 2 4 3 4 0 9 1 9 3 2 13 2 1 9 2
14 3 4 15 3 1 9 13 1 0 9 14 3 3 2
5 13 15 2 9 2
9 13 4 15 1 0 9 2 2 2
16 13 10 9 2 16 13 1 9 9 15 16 2 9 9 2 2
7 7 15 13 0 2 2 2
18 7 13 15 0 2 16 9 15 9 13 7 13 1 0 9 2 2 2
7 15 15 13 1 9 9 2
36 9 1 9 0 9 2 15 10 9 13 3 2 16 4 13 11 11 2 9 13 15 1 0 9 7 13 15 13 10 9 1 9 3 3 0 2
14 13 1 15 9 0 9 7 15 15 3 13 3 3 2
21 9 13 3 9 2 16 1 10 9 4 12 0 0 9 1 9 13 1 9 9 2
12 0 9 13 14 0 2 0 2 3 0 9 2
6 13 15 1 15 9 2
5 14 15 15 13 2
17 1 9 15 3 13 9 1 9 9 2 9 2 1 9 7 9 2
10 1 0 9 13 9 2 9 7 9 2
5 15 1 15 13 2
16 3 1 9 11 7 1 11 12 10 0 9 0 9 3 13 2
18 13 15 1 9 13 1 10 9 12 1 3 0 9 9 1 10 9 2
11 7 0 9 4 15 13 13 3 0 9 2
27 13 4 15 1 10 9 1 11 2 10 9 13 1 9 9 0 9 9 7 9 7 13 15 15 3 0 2
22 3 4 13 3 13 10 0 0 9 2 9 7 9 13 1 9 7 9 2 2 14 2
8 3 15 3 13 1 11 11 2
8 13 15 3 2 3 12 9 2
9 1 9 4 15 15 12 3 13 2
8 11 13 9 0 7 0 9 2
17 3 7 13 2 3 4 13 3 1 15 2 16 13 11 1 9 2
27 13 15 13 1 9 2 13 9 7 15 15 13 10 9 2 0 15 1 15 13 2 3 15 1 15 13 2
23 16 4 15 13 2 15 15 13 1 15 2 3 7 3 13 2 15 13 0 9 2 2 2
3 7 15 2
5 13 1 15 13 2
9 13 15 9 0 2 0 2 0 2
19 13 15 9 9 11 11 2 3 13 15 2 12 1 0 0 10 9 2 2
12 3 15 13 2 16 15 15 3 13 2 2 2
5 7 15 0 11 2
6 15 13 1 15 9 2
26 0 9 15 13 7 3 4 15 3 13 1 15 13 2 16 15 13 1 0 0 2 0 9 1 11 2
24 3 1 10 9 1 9 15 13 1 0 11 2 16 15 15 3 1 0 9 13 10 0 9 2
16 1 0 9 2 3 1 10 9 1 9 2 4 13 1 9 2
9 16 15 3 13 14 1 9 9 2
12 15 13 1 10 0 9 1 0 1 9 9 2
11 3 9 2 1 15 2 15 1 15 13 2
14 3 15 1 0 9 13 9 3 10 9 0 0 9 2
15 3 13 13 7 9 0 2 13 0 9 2 0 9 9 2
21 7 3 3 13 3 10 9 13 0 2 0 9 2 16 14 1 9 7 1 9 2
17 0 0 9 9 9 13 13 3 0 9 2 13 10 9 7 9 2
16 3 13 15 3 0 2 13 4 10 9 1 0 2 0 9 2
30 16 3 1 0 11 13 10 0 9 1 15 2 16 15 2 3 16 1 0 2 13 3 13 1 15 2 15 3 13 2
9 15 1 15 13 10 0 0 9 2
22 1 9 7 9 1 15 0 2 15 3 13 2 4 13 0 9 2 13 1 0 9 2
24 15 3 4 15 13 2 10 0 9 2 15 13 9 0 2 3 7 0 9 1 0 9 9 2
6 7 15 15 3 13 2
10 7 3 3 3 13 2 3 3 13 2
7 13 10 0 9 1 9 2
42 1 0 9 1 9 9 12 2 12 15 15 13 0 9 13 1 9 0 9 7 10 0 9 15 15 13 0 7 3 2 16 4 13 7 13 2 15 13 15 2 2 2
18 7 16 15 15 15 3 0 9 3 13 2 1 15 13 10 0 9 2
39 13 2 15 2 11 11 2 4 13 10 9 13 1 0 11 1 11 1 11 9 2 16 11 11 13 4 13 9 1 0 9 7 16 4 13 16 0 9 2
46 9 9 9 0 11 3 1 12 3 3 1 9 1 9 13 0 9 11 11 2 12 2 2 15 15 15 1 0 9 2 3 1 10 0 9 7 9 2 3 13 1 9 1 0 9 2
19 3 1 9 9 12 13 9 7 9 13 9 7 1 9 7 3 0 9 2
23 13 1 11 2 13 1 0 9 16 9 2 1 9 12 15 13 9 10 0 9 7 9 2
15 15 13 1 9 2 3 10 9 13 1 9 0 9 9 2
24 1 0 9 7 3 1 9 9 4 14 10 9 2 7 3 7 9 10 12 9 2 3 13 2
21 13 1 9 16 9 2 13 9 1 9 2 13 0 9 2 13 1 11 2 2 2
25 3 13 1 0 11 1 9 0 9 7 9 2 9 2 7 1 9 4 13 1 0 9 11 12 2
15 1 0 9 0 9 2 9 11 11 3 13 9 10 9 2
3 9 0 9
19 1 0 0 9 13 11 1 11 11 1 9 12 1 12 9 2 11 12 2
24 9 11 1 9 9 11 11 13 12 5 9 2 9 11 2 0 9 11 11 2 14 12 5 2
5 15 15 13 0 2
9 1 0 9 9 7 13 15 3 2
30 9 13 11 2 11 2 11 2 2 1 12 9 15 13 11 2 11 7 11 2 1 11 1 0 9 13 3 12 9 2
38 3 1 9 7 1 15 2 15 9 13 1 2 0 7 0 11 2 2 13 0 13 2 16 11 15 1 11 13 12 9 1 9 2 9 7 12 9 2
11 3 3 2 16 1 15 15 13 9 9 2
45 13 7 13 2 15 2 15 13 9 0 9 2 13 3 2 7 1 9 13 2 3 1 15 13 15 2 15 15 1 9 1 10 9 13 1 9 1 3 0 16 0 9 0 9 2
13 3 3 13 9 2 7 3 9 2 0 0 9 2
17 1 9 11 1 9 13 0 9 9 11 2 11 7 10 0 9 2
21 15 1 15 2 15 3 1 0 9 13 2 4 13 1 9 1 9 12 9 11 2
33 12 9 1 9 12 15 3 1 0 9 0 9 1 9 11 3 13 1 9 2 3 1 15 2 15 13 1 9 2 3 13 9 2
12 13 7 2 16 15 13 3 7 9 13 0 2
13 9 1 9 9 13 0 9 2 3 14 0 2 2
19 0 9 9 1 0 9 7 13 9 2 1 15 9 1 9 13 3 3 2
18 0 9 9 11 7 11 1 0 9 15 3 3 14 3 13 0 9 2
27 16 11 3 13 0 0 0 9 1 0 9 2 13 2 3 3 13 3 2 1 9 0 11 9 3 0 2
18 9 3 2 0 2 7 1 9 9 2 15 13 15 7 15 15 2 2
9 1 9 3 7 13 0 15 13 2
32 13 15 2 16 9 11 1 9 0 9 1 9 11 3 13 0 9 2 16 13 9 11 1 9 11 2 11 2 11 7 11 2
11 1 10 9 13 7 13 11 3 3 3 2
18 9 0 9 0 1 0 9 1 9 12 1 0 9 7 13 0 9 2
28 0 9 2 15 11 10 3 2 0 9 1 10 0 9 13 2 7 1 15 13 13 7 9 10 0 9 0 2
49 3 15 3 13 2 16 12 0 0 0 9 2 1 0 9 2 2 2 0 13 15 1 0 0 9 2 13 1 9 0 9 0 9 16 0 9 1 9 1 9 0 2 1 15 7 0 0 9 2
2 0 9
30 0 2 0 7 0 9 9 11 2 0 3 3 1 9 9 0 9 2 3 13 9 9 1 0 9 7 10 0 9 2
17 10 9 13 13 3 9 9 7 1 10 0 9 3 11 2 11 2
15 1 12 9 9 0 9 9 0 7 0 9 13 3 3 2
23 10 9 7 13 0 9 2 3 13 2 14 15 10 0 9 1 9 2 9 7 10 9 2
15 2 13 0 13 2 16 9 2 9 9 2 10 9 13 2
9 9 9 14 3 13 9 9 9 2
13 1 9 13 10 9 7 13 15 1 0 15 9 2
24 3 3 0 9 1 9 1 0 9 13 15 0 9 7 9 0 9 2 2 13 3 11 9 2
20 0 9 1 9 2 3 9 9 1 9 2 15 3 15 15 1 0 9 13 2
46 1 9 10 9 1 12 9 7 9 0 0 9 7 9 1 9 0 2 15 15 0 0 9 13 1 9 2 15 13 1 9 10 9 0 12 9 7 1 9 0 2 7 1 9 0 2
29 0 9 9 11 10 9 9 9 1 9 7 1 9 0 3 3 13 7 0 7 0 9 13 9 2 15 15 13 2
23 9 0 9 7 10 9 1 9 1 0 9 7 1 9 3 1 0 9 13 9 0 9 2
19 9 1 15 13 9 1 9 9 2 9 2 9 7 9 0 7 0 9 2
34 9 10 9 1 0 9 9 10 0 9 7 9 2 15 9 1 10 0 9 13 2 10 9 3 13 13 9 0 9 2 9 7 9 2
14 1 9 11 15 3 2 13 7 9 2 0 11 2 2
32 9 0 0 9 7 9 2 1 15 15 13 2 16 13 9 7 9 10 9 2 1 0 12 9 16 4 15 3 3 13 3 2
10 0 9 9 11 13 3 3 10 9 2
57 0 9 1 2 0 2 0 9 7 9 13 1 15 0 9 2 13 3 9 0 9 2 10 0 9 7 9 9 9 1 9 9 2 9 3 0 2 7 2 1 9 2 2 9 2 15 0 9 13 1 9 7 10 9 1 9 2
29 0 0 9 13 9 1 0 9 0 9 2 9 9 3 1 0 0 9 1 10 0 0 9 11 2 11 2 11 2
4 11 1 11 13
1 9
53 0 0 0 9 13 1 0 9 11 11 7 0 0 9 9 0 9 2 11 2 2 9 2 15 15 1 9 1 0 9 13 1 0 9 9 12 13 9 1 10 9 7 13 15 1 0 9 9 1 0 0 9 2
36 1 9 11 11 15 13 1 0 11 1 9 1 9 12 0 0 0 9 1 11 2 15 4 1 9 0 0 9 3 13 9 1 9 7 9 2
17 9 11 2 9 1 0 0 9 2 15 3 13 1 0 0 9 2
27 0 9 2 9 1 0 9 0 9 2 9 1 15 7 3 0 0 9 7 13 1 12 9 9 0 9 2
20 1 0 0 9 15 11 13 1 9 14 1 0 9 2 1 0 12 12 9 2
19 9 7 13 1 0 9 9 2 15 15 13 1 9 1 11 2 9 9 2
8 3 1 9 13 9 9 0 2
27 1 9 9 1 9 9 15 13 9 1 0 9 11 7 3 9 9 1 0 0 9 2 9 1 0 11 2
32 0 9 0 9 13 0 9 9 1 0 0 9 7 13 15 9 1 9 9 0 9 9 1 9 9 11 11 2 3 9 11 2
27 9 10 9 0 9 13 7 1 9 9 1 9 0 0 9 2 3 3 9 1 0 9 13 9 1 11 2
15 9 11 1 11 15 7 13 1 0 9 0 0 9 9 2
10 1 10 9 15 13 7 9 0 9 2
21 1 9 9 13 16 0 9 11 11 11 11 2 15 15 13 9 0 9 1 11 2
18 0 9 1 9 9 13 11 11 2 15 9 13 16 0 2 9 2 2
20 1 0 0 9 15 15 13 13 9 9 2 9 9 13 9 14 1 0 9 2
19 9 13 0 9 2 1 0 9 7 9 12 1 12 13 0 9 11 11 2
20 3 13 7 9 0 9 2 15 4 2 1 11 11 2 15 13 1 0 9 2
18 9 9 9 1 9 9 11 7 11 15 13 7 1 9 9 1 9 2
44 0 9 0 9 9 9 11 11 2 15 13 0 10 3 0 9 1 0 9 9 0 9 0 2 4 3 13 0 9 0 9 9 11 2 15 4 3 1 9 13 1 0 11 2
11 9 12 0 9 15 13 7 1 0 9 2
12 1 11 13 3 0 9 2 0 0 0 9 2
13 13 4 0 9 0 0 9 13 11 1 0 9 2
21 16 13 9 9 1 0 9 0 2 13 15 3 1 10 9 9 1 0 9 11 2
22 1 0 9 15 11 13 0 9 9 7 0 9 13 2 3 13 1 9 9 0 9 2
24 13 15 13 2 16 9 0 9 4 13 10 9 2 15 3 1 9 13 1 11 1 9 9 2
28 16 0 0 9 13 9 1 9 9 2 13 3 0 2 16 15 11 13 2 0 13 7 9 1 9 0 9 2
21 12 1 0 9 0 9 11 13 7 11 11 2 15 4 15 9 9 13 10 9 2
28 1 0 9 15 13 1 9 9 11 2 15 9 4 13 13 7 9 9 0 9 2 9 9 7 9 0 9 2
5 9 11 2 9 9
3 1 0 9
13 9 9 13 1 9 0 9 1 12 1 12 11 2
15 9 1 15 13 3 0 13 1 9 10 0 9 1 9 2
18 13 15 1 9 9 0 9 2 15 13 0 0 9 11 2 0 11 2
21 1 9 13 12 9 9 13 1 10 0 9 2 12 9 15 3 13 1 3 0 2
21 7 13 2 14 15 0 2 12 9 0 9 13 13 13 10 0 9 9 1 9 2
22 12 9 0 15 13 2 16 0 9 0 9 9 13 0 9 7 0 9 9 9 9 2
31 1 0 9 1 9 0 0 9 13 12 9 0 11 9 0 0 9 1 3 9 2 16 4 15 15 7 13 9 0 9 2
21 1 9 0 9 4 1 9 12 2 7 12 2 9 13 9 12 9 0 12 9 2
4 1 11 3 13
6 0 9 15 3 13 2
35 9 11 11 13 1 9 1 9 1 9 1 0 0 9 10 9 0 11 2 16 4 15 1 9 13 13 1 0 9 11 11 1 9 9 2
9 0 15 9 13 3 0 0 9 2
21 13 0 7 0 9 2 15 13 1 9 0 9 2 1 15 15 13 9 10 9 2
13 9 1 9 7 0 0 9 13 3 3 1 9 2
16 10 9 13 2 16 0 0 9 13 0 9 1 9 7 9 2
24 0 9 13 9 0 9 0 9 2 11 2 11 11 1 12 0 9 9 1 11 1 0 9 2
10 1 0 15 0 9 3 13 13 9 2
43 0 9 13 1 15 2 16 12 9 0 0 9 2 7 2 11 7 0 0 9 2 11 2 2 15 13 1 9 9 2 16 15 0 9 15 3 13 7 4 13 0 9 2
28 0 9 13 2 16 0 9 9 13 2 9 15 0 9 13 2 7 9 15 1 0 9 4 13 13 7 13 2
25 9 3 1 9 11 13 9 1 9 7 4 13 2 16 4 15 1 10 9 13 1 0 0 9 2
21 1 0 9 0 0 9 2 13 9 9 10 9 2 15 16 0 13 13 9 0 2
29 0 9 3 13 9 9 0 9 2 1 15 3 13 7 0 0 9 11 11 2 7 13 15 1 9 9 1 11 2
29 15 13 9 0 9 2 15 3 13 1 10 9 3 13 1 9 0 9 2 7 13 15 7 1 10 9 3 3 2
49 3 3 2 16 15 3 13 0 9 14 1 9 9 2 7 7 9 9 2 9 2 0 9 9 2 1 11 0 1 12 2 12 2 2 2 15 11 3 13 2 16 13 3 0 9 11 2 11 2
42 9 13 1 9 3 11 9 3 15 13 1 9 1 9 12 0 2 0 0 9 2 0 9 2 9 2 0 9 2 1 15 13 9 9 1 0 2 0 9 15 13 2
22 11 15 3 13 1 9 13 14 1 9 9 2 1 15 9 4 13 13 0 9 11 2
12 1 12 0 9 3 13 0 9 1 10 9 2
26 9 2 1 15 3 13 1 0 0 9 2 15 4 13 3 9 10 9 9 1 0 9 1 9 9 2
24 9 2 15 13 1 9 9 2 13 1 9 9 0 9 9 1 0 2 0 9 1 9 9 2
24 15 15 1 0 9 1 9 9 13 15 2 16 15 3 13 7 1 0 9 2 15 9 13 2
31 13 2 14 3 0 9 0 9 7 13 2 14 9 2 9 9 13 3 3 0 2 7 9 14 13 7 13 1 15 9 2
38 13 15 15 7 1 12 0 0 9 2 7 1 0 9 9 13 9 3 9 13 15 1 0 9 0 9 2 7 9 13 0 15 0 0 0 9 13 2
10 0 9 3 13 0 9 0 9 9 2
38 1 11 11 2 15 13 1 0 9 0 0 0 9 2 4 2 14 9 13 1 9 12 0 9 2 3 13 9 2 7 16 4 13 1 9 0 9 2
13 13 0 2 16 9 4 13 10 9 9 7 3 2
18 11 11 13 9 2 15 3 13 9 1 9 9 9 0 9 11 11 2
21 10 9 13 1 0 9 0 0 9 16 9 9 10 9 0 1 9 0 0 9 2
5 2 10 0 11 2
13 9 0 1 0 0 9 9 15 13 1 9 9 2
24 0 9 11 11 15 13 1 9 2 3 1 10 9 13 9 2 2 11 2 3 1 11 2 2
9 13 9 7 3 13 1 0 9 2
12 9 1 15 13 2 2 3 1 0 9 2 2
11 10 9 3 13 0 9 11 11 1 11 2
14 13 15 0 9 7 1 9 9 3 13 1 15 0 2
15 1 0 9 1 9 15 1 11 13 7 1 3 0 9 2
20 9 0 0 9 1 0 7 0 11 1 11 15 13 0 9 15 9 0 9 2
10 0 9 11 11 13 10 9 3 3 2
15 1 9 1 9 11 0 9 13 2 2 11 13 0 9 2
13 4 15 11 13 2 16 13 3 13 7 14 2 2
45 16 1 9 0 9 13 11 11 1 9 2 1 9 9 7 1 9 2 16 4 10 9 13 3 2 13 2 2 3 13 13 2 3 10 0 9 13 3 3 3 3 13 1 11 2
10 14 15 13 13 3 7 3 11 13 2
11 3 15 11 13 2 16 11 13 10 9 2
6 7 1 15 13 13 2
4 1 11 2 2
28 1 10 0 9 9 9 3 15 13 7 9 13 0 9 10 9 2 11 13 9 1 9 11 1 9 0 9 2
37 0 9 0 9 11 13 9 1 12 9 0 9 2 15 15 13 1 9 13 14 1 0 9 7 1 3 0 9 15 13 13 9 0 9 1 11 2
9 10 9 3 13 0 13 1 0 2
8 4 13 2 0 9 7 13 2
36 3 3 13 13 15 2 16 0 9 13 2 10 9 13 9 9 1 11 15 2 15 15 1 0 11 13 3 3 13 7 13 15 0 9 11 2
21 15 15 3 13 2 16 4 0 9 3 13 0 9 7 3 15 15 13 1 11 2
20 1 0 9 15 13 3 13 2 10 9 15 4 13 1 0 9 0 0 9 2
23 11 13 0 9 15 2 16 9 1 0 9 13 0 7 16 13 0 15 13 1 15 9 2
18 3 13 7 1 9 0 0 9 13 3 16 9 1 0 9 0 9 2
18 9 2 9 2 7 2 9 2 15 13 9 9 9 0 9 1 11 2
31 1 15 15 3 3 13 2 0 9 2 2 0 9 9 11 11 2 15 0 9 13 0 9 1 9 2 3 2 11 2 2
7 13 2 2 11 13 9 2
11 3 4 13 9 1 9 13 9 7 9 2
6 13 15 13 15 2 2
18 0 10 9 15 3 13 0 0 9 11 11 2 14 9 13 3 0 2
17 1 0 9 13 1 0 9 9 2 10 0 11 2 13 3 3 2
24 13 15 3 3 16 9 9 11 2 7 9 2 3 3 2 13 2 14 9 0 9 1 11 2
8 3 13 9 0 9 13 3 2
16 7 11 15 13 1 10 9 1 0 7 1 0 1 0 9 2
16 15 15 3 1 9 3 15 0 9 13 13 2 3 9 13 2
9 3 13 3 3 0 9 9 0 2
13 0 15 3 13 2 13 10 9 7 9 7 9 2
12 9 1 15 13 1 2 0 11 2 10 9 2
31 1 0 9 0 0 9 13 1 9 9 11 2 12 1 0 9 9 9 1 9 12 2 10 9 2 2 10 0 0 9 2
9 14 15 13 3 1 9 0 9 2
15 7 3 15 2 11 2 13 7 13 9 11 2 2 2 2
10 3 2 16 13 0 9 11 11 9 2
31 1 10 9 1 9 9 1 9 13 2 16 15 2 15 13 3 1 11 2 15 13 2 16 4 15 13 10 0 9 11 2
8 1 9 11 10 10 9 13 2
10 3 2 16 15 15 10 0 9 13 2
14 7 3 12 2 9 13 2 2 0 9 0 9 13 2
15 11 15 13 13 15 0 9 7 2 16 15 13 9 9 2
11 16 10 9 13 1 11 2 13 0 11 2
11 13 10 9 2 16 15 15 15 13 2 2
12 3 1 12 9 3 13 9 1 9 0 9 2
20 13 0 11 13 2 16 11 13 10 0 9 7 16 15 1 12 9 4 13 2
27 11 13 3 3 0 9 7 13 0 2 15 7 1 10 9 4 13 1 9 10 3 3 0 9 0 11 2
13 9 3 11 11 13 7 1 9 1 11 13 9 2
14 11 11 13 3 9 2 16 0 0 9 13 1 9 2
14 7 13 2 14 1 11 9 7 14 2 13 15 0 2
16 7 9 0 9 1 11 4 13 2 16 0 9 4 9 13 2
9 11 15 13 10 9 3 3 0 2
19 9 11 15 13 3 3 2 2 13 15 13 0 2 7 13 15 15 13 2
8 3 15 15 4 3 13 2 2
20 3 13 1 15 2 16 15 4 3 13 0 9 1 9 11 2 7 11 15 2
6 13 7 3 12 9 2
22 16 9 0 9 13 13 9 0 9 16 9 0 9 7 4 15 13 15 10 9 13 2
12 1 9 7 0 9 1 2 10 0 11 2 2
23 10 9 2 15 3 13 0 9 2 13 1 11 1 10 9 1 2 0 9 2 0 9 2
5 11 2 9 1 9
4 11 2 11 2
34 1 9 9 2 15 13 1 9 3 2 15 1 11 1 0 9 7 1 3 0 9 3 13 9 2 16 3 0 16 1 9 9 9 2
19 9 1 0 9 7 0 9 9 13 1 0 9 13 3 1 0 9 11 2
14 1 9 9 9 15 3 3 3 13 0 7 0 9 2
28 10 0 9 15 7 3 3 13 3 13 9 7 13 9 1 0 9 2 10 0 9 15 13 1 9 1 11 2
8 3 7 13 1 10 9 9 2
28 3 13 1 0 0 9 1 11 9 0 9 9 11 11 2 0 9 14 13 1 0 9 2 16 4 3 13 2
12 13 3 2 16 10 9 13 0 3 1 11 2
16 15 11 3 3 13 9 11 11 1 0 9 1 9 0 9 2
12 13 2 16 9 1 0 9 13 13 10 9 2
13 3 13 0 0 9 2 15 13 13 9 2 13 2
44 0 9 11 11 3 13 2 16 1 9 15 1 0 9 11 0 14 12 9 3 1 11 13 9 0 7 0 0 9 2 1 15 15 13 9 12 9 1 9 0 9 1 11 2
10 12 9 15 1 11 13 1 12 9 2
12 11 7 3 1 9 13 1 12 9 0 9 2
22 9 11 1 0 9 3 13 2 16 0 9 15 1 0 9 9 1 11 13 9 9 2
21 13 7 2 16 0 9 1 15 13 0 9 2 15 13 9 0 9 1 0 9 2
11 1 9 3 1 11 13 14 12 0 9 2
30 11 3 13 2 16 9 2 15 13 2 13 1 9 1 9 0 9 1 11 1 12 9 7 9 7 12 9 4 13 2
4 9 1 0 9
9 11 2 11 13 1 11 1 0 9
4 11 2 11 2
15 0 9 1 0 9 15 13 1 0 9 2 7 13 3 2
31 13 15 3 1 11 9 9 1 9 11 2 11 2 11 11 1 0 9 1 9 9 11 11 7 0 9 1 9 11 11 2
9 2 13 13 1 0 9 2 2 2
12 13 4 15 7 1 0 9 2 2 13 11 2
12 13 9 2 16 11 4 13 13 9 1 9 2
18 13 2 16 0 9 11 1 10 0 9 1 11 13 7 13 0 9 2
7 11 13 9 1 3 0 2
23 1 10 9 13 0 0 9 13 7 13 0 9 2 16 13 15 4 13 9 1 0 9 2
28 0 9 11 2 3 13 2 13 1 9 1 11 2 16 2 3 13 10 0 9 2 7 4 13 0 9 9 2
19 13 15 1 0 9 0 9 0 2 11 2 15 13 1 10 9 1 11 2
29 9 13 2 16 10 9 13 0 2 16 15 11 2 0 0 9 2 13 13 2 1 9 2 15 15 4 13 2 2
30 9 0 9 15 3 13 1 0 9 1 0 9 1 0 2 0 9 1 0 11 2 7 15 13 1 0 0 9 13 2
8 13 15 0 9 1 0 11 2
17 15 3 13 2 16 0 9 3 13 1 0 9 1 9 0 9 2
7 9 11 7 11 1 11 13
2 11 2
15 1 0 9 9 4 3 3 13 0 9 0 9 7 11 2
36 9 15 13 9 9 9 11 11 11 2 9 0 9 9 9 11 11 11 2 0 9 9 11 1 11 11 11 7 0 9 0 9 0 1 11 2
15 9 13 0 9 9 11 7 11 1 12 2 9 9 11 2
33 9 13 1 9 0 9 9 7 0 11 1 9 12 2 3 15 0 9 13 13 1 0 9 11 11 1 9 0 9 12 2 9 2
20 9 13 1 3 0 9 9 7 4 3 13 1 9 7 0 9 1 0 9 2
4 9 9 15 13
5 11 2 11 2 2
32 12 9 1 9 11 1 0 9 15 1 9 13 0 9 9 1 9 11 1 9 0 11 2 7 3 3 13 9 1 9 12 2
14 0 1 9 13 12 9 1 9 1 3 12 0 9 2
11 13 15 1 9 2 9 7 9 0 9 2
15 3 9 1 9 13 12 0 9 0 9 1 9 11 11 2
16 2 10 9 13 3 15 2 15 10 9 3 13 1 10 9 2
39 15 2 15 3 13 2 15 13 11 0 2 15 2 15 13 2 15 4 13 2 16 4 13 0 2 2 13 11 2 15 4 1 0 0 9 13 1 9 2
1 3
8 9 1 9 0 9 13 0 2
32 16 7 13 0 13 0 9 2 13 9 9 9 9 1 9 2 13 3 1 9 1 9 9 11 7 9 1 9 9 11 11 2
30 0 9 11 11 2 11 13 9 9 13 9 0 9 1 0 9 11 2 15 2 16 9 13 2 3 13 10 0 9 2
27 9 9 13 1 0 9 9 9 2 15 13 2 16 16 15 1 0 9 13 0 9 2 0 9 11 13 2
21 0 9 15 13 1 9 1 0 9 2 16 4 13 9 11 1 0 9 1 11 2
14 0 9 9 9 1 9 13 4 13 0 9 1 11 2
17 12 9 15 13 9 1 9 7 9 2 1 15 13 1 9 11 2
11 12 9 4 13 7 1 12 9 4 13 2
18 9 13 2 16 9 9 13 10 9 2 16 4 15 13 1 0 9 2
24 1 9 1 2 0 2 9 13 11 13 7 0 0 9 9 2 15 13 3 16 12 9 9 2
22 16 13 0 9 9 7 9 11 11 2 11 13 1 9 9 9 13 0 0 9 11 2
12 0 0 9 1 0 9 11 3 13 0 9 2
12 13 15 0 0 9 0 15 11 1 9 9 2
14 9 13 9 1 9 9 2 7 3 3 13 10 9 2
26 9 1 11 1 9 12 9 9 13 1 0 9 0 9 11 2 11 2 15 13 1 0 9 1 9 2
14 3 13 2 16 10 9 4 3 13 9 9 1 9 2
16 9 1 0 9 10 0 9 2 11 2 13 3 9 10 9 2
12 11 15 13 1 0 0 0 9 2 11 2 2
34 1 9 13 9 0 1 11 1 10 9 1 11 1 9 12 13 3 1 11 0 9 9 9 11 11 11 11 1 0 9 9 11 11 2
8 11 13 9 1 12 0 9 2
15 1 0 9 1 9 9 11 11 13 9 0 9 1 11 2
19 0 9 3 13 1 10 9 0 9 1 9 1 9 12 11 0 1 11 2
9 13 15 9 0 9 9 1 11 2
21 1 0 9 13 10 9 0 9 1 0 9 9 1 0 0 9 10 9 0 11 2
43 1 12 9 9 13 3 9 1 9 11 1 9 11 12 0 11 2 15 15 0 9 13 9 1 9 7 9 0 9 2 1 15 12 9 13 1 9 7 12 9 4 13 2
21 1 9 13 3 2 16 14 12 11 13 9 9 2 15 13 9 3 0 0 9 2
20 9 9 11 13 11 10 0 9 11 2 16 4 15 13 13 0 7 0 9 2
17 1 9 1 0 9 11 11 15 3 13 0 9 1 9 11 11 2
11 12 2 9 3 13 11 11 1 0 11 2
27 13 15 1 11 9 11 2 15 2 13 0 7 13 9 2 2 7 1 9 0 9 7 13 3 15 9 2
30 2 1 9 4 13 14 12 9 7 1 15 15 13 2 2 13 2 16 3 13 2 3 13 7 13 15 1 0 9 2
4 0 9 13 9
2 11 2
21 0 9 1 11 7 1 15 0 9 15 9 4 13 13 1 0 9 0 0 9 2
20 9 11 1 9 12 13 1 9 1 9 7 1 15 7 10 9 13 0 9 2
21 0 9 1 9 0 9 13 1 11 1 0 9 0 9 1 9 9 9 9 9 2
24 3 13 9 9 3 1 12 9 2 13 15 9 9 1 9 7 13 9 13 9 7 0 9 2
30 2 9 9 1 11 13 2 16 13 15 9 3 2 2 13 11 11 1 0 0 11 1 9 1 0 15 0 0 9 2
9 9 9 14 3 13 1 10 9 2
5 0 9 13 10 9
2 11 2
26 0 9 1 0 9 11 1 9 13 9 1 9 2 16 0 9 13 9 2 15 13 1 9 1 15 2
18 1 9 13 2 16 16 9 1 10 9 13 2 13 0 9 1 9 2
14 9 3 1 9 0 9 1 0 9 2 11 2 13 2
42 9 4 13 3 2 16 13 0 11 1 9 11 9 9 1 9 7 9 0 9 11 11 2 15 15 13 1 9 1 9 7 11 7 15 10 9 13 1 9 1 9 2
5 9 15 1 9 13
11 1 9 1 0 9 1 11 13 13 15 0
20 1 11 15 9 13 7 9 13 0 2 16 13 2 16 13 0 2 13 15 2
44 0 9 0 9 2 12 9 9 1 12 9 2 15 13 1 0 9 1 9 12 2 1 0 7 9 2 12 2 12 9 2 1 12 9 3 16 1 12 9 2 13 1 9 2
13 0 9 16 1 9 12 9 2 3 12 2 13 2
19 9 15 3 13 1 0 0 9 0 9 16 1 0 9 2 12 9 2 2
18 1 3 0 13 1 9 2 1 15 15 15 1 0 9 13 14 13 2
25 9 13 3 1 9 9 1 9 2 3 15 7 11 13 14 1 2 0 2 0 9 9 0 11 2
31 7 16 0 9 13 1 11 1 9 14 1 12 9 2 12 1 9 13 7 13 15 0 9 2 2 0 9 9 15 13 2
40 9 11 7 9 9 11 11 3 13 3 9 7 9 1 9 1 11 7 13 15 13 1 2 0 9 2 1 0 9 2 0 11 2 11 2 11 7 11 2 2
22 2 13 15 2 16 3 13 1 0 3 7 16 15 1 15 13 13 2 2 13 9 2
14 0 9 1 9 0 9 13 14 0 9 2 7 9 2
22 10 0 9 13 14 0 9 1 0 0 9 0 11 2 11 2 3 13 12 9 11 2
13 3 15 4 13 1 0 9 16 1 9 1 11 2
24 1 12 0 9 4 13 3 0 2 7 0 9 2 1 12 15 4 13 9 1 0 0 9 2
14 1 10 9 13 0 9 11 1 11 13 3 0 9 2
41 16 4 0 9 9 11 11 1 9 9 11 2 11 13 2 13 4 15 9 13 0 9 9 2 7 15 13 1 0 0 9 2 3 0 1 0 9 2 3 0 2
37 1 0 11 2 11 1 9 9 4 0 9 2 3 16 1 11 2 13 10 9 1 0 9 9 2 0 9 2 3 13 13 0 9 1 0 9 2
21 3 9 1 9 13 1 0 9 9 0 9 13 0 0 9 13 9 1 9 9 2
10 9 15 1 0 9 13 1 9 13 2
28 1 0 2 16 0 9 11 11 2 15 13 3 13 0 0 9 3 3 3 0 2 15 1 11 13 0 9 2
10 0 0 9 15 7 1 9 3 13 2
24 9 1 0 11 2 11 13 0 9 2 15 13 7 15 2 15 13 2 16 11 1 11 13 2
20 1 9 3 13 2 16 9 2 10 9 13 0 7 0 9 11 2 13 13 2
17 13 3 3 2 0 9 9 11 3 13 9 13 0 9 1 11 2
23 9 0 15 1 9 2 0 9 10 9 2 13 3 3 3 0 7 3 3 13 1 9 2
5 9 11 1 9 12
5 0 9 9 12 2
24 1 0 9 9 1 9 1 0 9 13 12 9 0 0 9 0 9 1 9 9 11 9 11 2
11 0 9 13 0 9 0 9 10 9 13 2
23 16 15 13 10 0 9 9 9 13 9 7 1 0 9 2 13 15 0 9 9 3 13 2
8 13 15 7 9 3 13 9 2
29 9 2 15 13 0 11 1 12 2 9 12 13 0 7 0 9 2 15 13 1 9 1 9 9 12 2 4 13 2
12 9 1 0 9 15 7 13 2 13 3 3 2
24 16 10 9 1 9 0 9 7 1 9 9 0 9 1 11 3 13 2 13 3 1 0 9 2
23 3 13 3 13 0 9 9 2 7 13 7 0 9 1 9 0 9 2 15 1 0 9 2
11 9 9 11 4 3 1 9 13 7 9 2
46 9 9 2 9 9 7 9 2 13 3 0 2 13 2 14 12 1 0 3 1 9 3 1 9 3 2 13 14 1 3 3 3 0 9 1 10 2 10 9 13 10 9 0 9 2 2
17 0 9 4 0 9 3 13 16 9 13 9 7 16 0 0 9 2
24 3 9 9 1 10 9 9 13 0 9 2 15 15 1 0 9 13 9 0 9 7 0 9 2
20 9 1 0 9 10 9 13 11 0 9 7 13 9 0 9 1 15 7 9 2
13 9 9 9 3 13 9 3 1 9 0 0 9 2
21 1 0 9 0 9 9 13 7 13 11 1 9 9 12 9 14 1 12 9 9 2
16 1 15 13 13 7 12 9 2 15 9 1 9 11 3 13 2
29 3 3 15 13 9 2 7 15 14 0 9 2 2 16 11 0 9 9 13 7 16 13 10 0 9 14 15 0 2
20 3 16 1 9 9 0 11 13 14 1 0 9 1 9 11 3 1 9 12 2
13 9 10 0 9 3 0 9 13 3 7 14 15 2
36 1 9 2 15 1 9 0 9 13 1 0 9 2 13 3 0 9 0 9 2 9 0 0 9 9 2 7 0 9 2 9 0 9 11 2 2
12 13 13 13 10 9 1 9 3 1 0 9 2
26 1 9 1 0 9 12 9 9 15 3 10 9 1 0 9 13 2 13 3 1 9 0 11 11 2 2
16 0 9 2 9 7 0 9 9 2 13 3 1 9 9 9 2
23 1 12 0 9 7 12 0 9 2 1 9 9 3 0 2 15 9 13 16 0 0 9 2
8 13 12 0 9 7 9 9 2
24 1 15 15 13 1 0 9 2 10 9 4 1 0 12 9 13 13 9 1 9 9 0 9 2
34 1 9 9 11 11 2 16 0 9 0 0 9 2 15 7 3 13 9 2 1 0 9 9 0 9 2 1 9 9 15 0 9 3 2
31 13 13 1 15 2 16 0 9 1 9 9 3 13 3 0 9 2 16 4 13 9 9 9 7 16 4 3 0 9 13 2
28 7 9 3 13 9 2 16 4 1 0 9 13 2 16 16 4 15 13 1 0 9 0 9 3 2 9 11 2
34 0 9 9 11 11 3 13 2 16 1 9 9 12 3 13 1 9 11 0 9 2 10 0 9 11 7 13 2 16 15 0 3 13 2
22 1 0 7 0 9 13 7 0 2 16 4 11 9 13 7 4 3 1 0 9 13 2
24 3 7 3 13 10 9 1 0 2 16 1 9 1 0 0 9 13 2 3 2 1 9 9 2
22 1 9 9 0 9 1 9 9 9 13 2 16 1 9 10 9 4 13 13 0 9 2
24 9 13 0 2 1 15 2 15 13 2 15 13 15 9 0 9 1 9 7 0 9 14 13 2
4 3 3 7 15
5 0 9 0 9 2
11 3 13 3 13 0 9 0 9 1 11 2
31 13 3 0 9 9 2 9 7 9 0 9 2 3 13 1 9 0 0 9 2 9 1 0 9 7 1 9 1 9 9 2
11 1 11 13 3 0 9 9 7 0 9 2
11 3 0 0 9 13 0 9 1 0 9 2
21 3 3 7 13 3 1 9 9 2 16 1 9 12 15 9 13 3 3 7 3 2
25 13 15 2 16 10 9 13 3 13 9 1 9 16 0 9 2 15 1 9 14 3 13 10 9 2
20 9 13 9 0 9 1 9 7 3 9 9 9 2 11 2 11 2 11 2 2
27 1 10 9 13 0 9 9 3 13 2 13 2 13 2 16 13 0 9 16 13 9 9 7 9 9 9 2
15 13 0 9 13 1 0 9 14 9 0 2 7 7 0 2
17 0 0 9 2 0 9 7 9 1 9 13 1 3 16 0 9 2
23 0 12 9 1 9 4 3 13 0 0 0 9 1 0 0 9 7 3 0 9 1 9 2
9 1 0 9 4 13 9 13 9 2
4 3 7 3 2
17 3 3 9 11 11 1 9 15 3 13 9 1 9 1 9 9 2
15 9 0 9 2 15 3 13 9 2 13 9 9 0 9 2
11 1 9 0 9 13 0 9 0 9 9 2
15 9 2 0 16 0 9 2 9 9 2 9 7 0 9 2
15 13 15 1 0 2 9 0 9 3 13 0 9 0 9 2
24 1 15 15 3 13 0 9 2 2 13 0 7 0 9 9 2 7 13 15 0 9 1 9 2
12 1 0 9 4 13 3 0 7 3 15 13 2
19 7 3 13 0 9 2 7 13 15 13 2 3 4 15 9 13 13 2 2
4 1 9 9 2
27 1 9 0 9 13 2 3 13 1 0 0 9 0 9 9 2 10 9 2 15 15 13 1 0 0 9 2
21 1 9 1 11 13 11 0 9 2 9 15 1 11 2 15 15 13 1 11 11 2
13 13 3 0 9 2 9 1 9 7 3 0 9 2
19 13 15 2 16 1 9 15 3 13 1 0 9 2 10 0 9 13 13 2
7 1 10 9 15 4 13 2
8 7 3 3 2 10 0 9 2
22 0 11 13 0 9 2 15 13 9 7 13 4 15 13 2 16 13 0 9 4 13 2
3 9 9 2
10 9 15 13 7 15 15 15 13 13 2
18 3 14 0 9 9 9 2 16 9 9 13 15 7 0 9 15 0 2
8 0 9 15 3 13 3 3 2
4 0 9 1 9
1 9
21 9 1 0 9 2 15 1 9 13 0 9 11 2 13 3 9 7 9 11 11 2
41 3 3 2 3 9 9 11 13 1 9 2 9 0 9 2 2 9 1 9 1 15 7 11 11 13 2 16 9 0 1 9 9 13 1 0 7 10 9 1 0 2
59 16 0 9 9 9 13 13 2 16 9 1 0 9 13 3 7 2 16 4 9 13 9 1 10 9 1 0 9 2 13 15 9 13 2 16 2 16 15 0 9 13 2 13 15 3 9 1 0 9 2 16 15 13 3 2 3 13 2 2
20 9 11 3 13 9 13 15 2 16 9 9 13 1 0 9 3 1 10 9 2
47 10 9 7 13 1 15 2 16 11 11 1 0 9 1 11 13 2 16 1 15 2 16 4 9 9 4 3 13 2 13 15 7 13 15 1 15 9 9 0 9 7 9 2 15 15 13 2
24 13 15 1 15 0 9 2 15 10 0 9 2 16 3 1 0 9 15 13 2 13 1 9 2
9 9 11 3 9 9 1 15 13 2
29 13 10 0 9 1 15 0 2 13 2 14 15 1 0 9 1 10 9 2 13 15 2 16 3 13 1 10 9 2
47 10 0 9 3 13 9 2 16 9 9 15 1 15 13 9 2 3 15 13 1 9 0 9 1 11 7 3 1 10 9 11 11 2 1 15 15 3 9 13 1 9 1 9 10 0 9 2
8 9 9 15 13 13 1 9 2
30 16 0 2 7 0 9 9 11 1 9 13 7 13 1 15 2 7 3 1 0 11 2 3 15 1 0 9 3 13 2
17 15 3 13 11 2 16 4 3 13 10 9 0 9 1 0 9 2
18 3 2 16 13 3 7 9 1 9 1 0 9 1 11 2 14 15 2
1 9
37 12 9 1 11 1 9 1 12 1 12 9 7 12 12 0 1 11 1 9 1 9 1 9 11 13 12 0 9 1 11 7 1 9 0 1 11 2
10 0 9 1 9 7 9 13 13 9 2
18 9 3 13 7 2 16 12 1 12 0 13 3 3 13 0 1 15 2
10 9 4 13 1 0 9 9 1 9 2
10 9 9 13 1 0 9 12 0 9 2
16 1 9 15 2 1 9 0 2 9 2 11 11 13 0 9 2
17 9 2 15 14 13 1 9 2 16 15 13 2 13 3 1 9 2
26 1 9 0 1 0 11 1 11 13 1 9 1 9 11 2 11 1 9 1 12 0 0 9 12 9 2
15 12 1 15 15 13 1 9 9 7 0 12 15 13 9 2
9 13 15 12 9 7 1 9 13 2
6 0 9 1 9 11 11
2 0 9
2 11 2
12 9 11 11 13 3 3 13 0 9 1 11 2
16 0 9 15 13 2 16 12 1 0 4 3 13 1 10 9 2
21 9 9 11 11 13 2 16 9 15 4 1 0 9 13 3 12 9 1 0 9 2
18 15 15 13 9 0 9 1 9 1 9 9 1 11 12 1 0 9 2
17 10 9 15 13 9 13 3 1 9 2 3 7 11 2 11 13 2
15 1 0 9 13 1 10 9 16 9 13 9 11 2 11 2
34 0 9 13 9 2 15 13 11 1 9 0 9 7 1 9 2 15 9 13 13 9 1 11 7 1 11 1 0 9 14 12 9 9 2
26 11 13 3 13 1 9 9 0 9 2 16 13 9 9 1 9 9 1 0 0 9 7 3 15 13 2
18 3 13 3 13 0 9 1 9 1 11 1 11 1 9 1 12 9 2
20 9 15 13 1 0 9 2 1 15 13 4 9 13 9 1 12 7 12 9 2
28 0 3 13 2 16 15 13 13 0 7 13 3 2 16 4 13 15 0 1 0 9 0 1 9 1 0 9 2
16 16 13 13 2 9 13 10 9 1 9 7 1 0 0 9 2
9 9 4 13 13 1 12 2 9 2
12 0 9 13 0 0 9 3 14 9 2 13 9
2 11 2
23 9 9 2 15 13 1 9 0 7 0 9 7 4 13 1 9 2 15 13 9 0 9 2
24 3 15 3 13 2 13 2 3 7 3 0 0 2 9 2 2 15 15 13 1 11 7 9 2
12 11 15 13 11 11 1 0 9 0 0 9 2
19 1 15 14 1 0 9 9 13 9 0 9 9 9 2 7 15 15 13 2
16 0 9 1 9 1 2 0 9 2 1 15 13 0 0 9 2
25 0 1 0 9 13 1 9 0 9 2 1 0 9 2 13 15 1 9 7 1 9 1 9 9 2
18 3 13 10 0 9 1 9 2 3 3 1 2 9 1 9 9 2 2
28 1 3 0 9 15 7 3 13 0 9 1 0 2 0 2 9 2 3 9 1 0 11 2 3 3 1 11 2
17 9 15 1 15 9 13 1 9 1 10 9 9 1 10 12 9 2
15 0 1 15 2 15 13 1 0 9 2 13 1 9 9 2
15 1 12 9 9 13 3 13 2 1 0 9 7 9 13 2
6 9 15 15 3 13 2
22 14 15 1 9 2 15 15 13 13 3 1 11 2 13 3 1 9 0 1 9 13 2
15 9 7 1 10 9 13 9 2 3 4 15 9 3 13 2
16 3 2 3 13 9 0 13 2 13 3 2 9 2 1 9 2
18 9 9 2 1 10 13 9 9 2 15 13 3 1 12 7 12 9 2
7 2 14 3 13 0 9 2
11 16 15 15 15 13 2 13 15 3 9 2
19 13 9 2 16 1 10 9 15 3 13 0 9 2 2 13 11 2 11 2
14 14 1 0 9 13 0 9 12 9 0 3 1 9 2
7 1 9 12 15 13 12 2
3 13 0 9
2 11 2
27 9 9 13 13 9 2 15 15 0 9 1 9 1 9 1 9 13 1 9 9 0 0 9 1 11 12 2
31 1 9 0 9 13 9 0 2 12 9 0 2 0 1 0 9 7 0 0 9 1 9 2 0 9 9 12 5 12 2 2
19 9 13 15 2 15 15 1 15 15 13 2 16 4 15 13 1 9 12 2
6 1 0 9 15 14 13
6 11 11 1 9 1 11
14 9 0 7 0 0 9 13 9 9 1 3 0 9 2
12 15 4 13 13 9 1 9 0 2 0 9 2
9 1 9 11 13 9 11 11 11 2
7 13 16 9 9 0 9 2
19 13 4 7 1 9 0 9 9 1 9 0 9 9 7 0 9 0 9 2
12 9 1 9 13 15 2 15 15 1 15 13 2
9 13 7 3 0 13 9 0 9 2
12 13 2 16 9 10 9 13 3 7 9 11 2
21 7 1 9 1 0 9 3 3 13 2 16 9 0 9 13 1 9 9 2 9 2
6 13 3 13 0 9 2
9 15 3 7 13 9 0 9 13 2
17 3 0 13 9 13 3 1 9 7 9 13 1 0 9 1 9 2
20 9 9 13 1 0 9 13 9 10 9 9 9 1 9 9 0 9 1 9 2
6 15 13 1 15 3 2
11 9 7 13 1 9 0 0 9 0 9 2
18 13 1 15 13 9 2 15 4 10 9 13 3 1 9 7 0 9 2
17 13 2 16 1 0 9 4 15 13 13 9 9 3 0 0 9 2
7 15 4 10 9 13 13 2
18 13 1 9 0 9 2 3 15 9 13 13 3 0 9 9 1 9 2
35 1 9 2 3 9 1 0 9 9 7 9 13 1 9 0 9 2 4 13 9 9 2 15 4 13 0 9 1 9 2 16 13 12 9 2
9 0 9 4 1 15 13 13 9 2
12 15 4 1 0 9 13 3 9 1 9 9 2
33 15 2 15 1 0 9 13 13 12 9 0 9 2 1 15 4 15 13 9 3 0 9 2 13 1 0 9 3 3 9 7 3 2
15 3 15 13 9 9 9 2 15 4 1 0 9 13 9 2
10 13 4 15 13 1 9 1 0 9 2
19 3 1 11 15 3 13 10 9 13 0 0 9 1 9 12 9 0 9 2
8 0 7 0 9 13 13 9 2
10 13 7 2 16 15 13 13 3 3 2
6 13 15 9 0 9 2
5 11 11 1 9 13
3 1 0 9
2 11 2
35 1 9 1 11 11 2 15 15 1 0 9 0 9 1 11 13 1 9 13 1 9 2 13 0 0 9 11 11 13 1 9 1 9 13 2
9 1 9 3 13 9 1 9 11 2
19 1 9 1 11 13 2 16 1 15 13 1 10 9 9 15 1 0 9 2
8 11 2 11 7 11 13 1 9
3 1 0 9
4 11 2 11 2
27 0 9 1 0 9 13 0 9 9 9 11 11 1 0 2 0 9 9 0 0 9 11 2 11 11 11 2
15 13 2 16 2 13 15 9 2 1 15 15 13 13 2 2
9 2 11 15 15 3 4 3 13 2
20 7 13 2 16 13 13 2 16 4 3 13 2 16 13 0 2 2 13 11 2
10 1 9 9 15 13 7 0 9 9 2
12 2 13 15 7 2 16 13 4 9 13 3 2
31 15 4 13 1 15 2 16 15 0 0 9 1 9 1 9 0 11 10 0 9 13 1 15 2 2 13 9 11 11 11 2
10 1 11 4 15 0 9 13 13 10 9
2 11 2
22 9 4 1 9 11 11 11 13 13 10 9 2 16 4 1 0 9 13 3 10 9 2
12 13 2 16 15 13 0 9 11 1 0 9 2
27 9 11 1 9 13 1 9 1 0 9 10 9 11 2 2 15 13 1 9 9 11 13 3 1 9 2 2
20 1 10 9 3 13 9 0 9 11 11 11 2 15 15 13 13 1 9 9 2
24 2 1 9 2 16 15 11 1 9 13 13 1 11 2 4 3 13 2 2 13 11 9 11 2
19 9 11 3 1 11 13 1 0 9 2 15 4 15 13 13 1 0 9 2
25 11 13 2 16 4 10 9 1 9 9 0 9 13 1 9 1 0 9 11 13 1 0 9 3 2
31 2 9 13 3 4 13 3 3 2 16 1 9 7 12 0 9 13 10 9 0 9 16 9 0 0 9 2 2 13 11 2
15 9 11 11 11 14 3 13 2 16 0 9 4 13 3 2
18 16 3 13 9 11 2 13 15 2 16 9 0 9 11 13 1 11 2
31 2 13 4 7 1 0 2 16 4 1 9 2 16 15 11 13 10 0 9 2 13 0 9 10 9 2 2 13 11 11 2
8 9 4 13 3 13 7 0 9
2 11 2
25 13 9 9 1 0 9 1 9 4 13 9 1 0 0 9 2 15 9 13 1 10 9 9 9 2
12 3 13 9 9 13 3 0 7 0 0 9 2
32 9 15 7 13 2 16 13 0 13 9 7 1 9 9 10 9 2 3 0 7 0 9 2 1 9 0 9 7 9 0 9 2
72 1 0 9 0 9 13 2 16 4 0 0 9 13 3 1 0 0 9 7 0 9 9 1 0 9 2 9 0 9 2 0 9 2 0 9 0 9 2 0 9 2 0 9 2 9 9 2 9 0 9 1 0 15 9 2 9 10 9 2 9 9 2 9 9 2 9 7 9 0 9 3 2
24 0 9 2 15 1 0 9 13 1 9 2 13 13 9 9 2 7 15 7 1 9 0 9 2
12 1 9 9 13 9 9 14 1 12 12 9 2
11 9 13 2 16 1 0 9 3 13 12 9
2 11 2
22 1 12 9 15 3 13 9 0 9 15 3 0 0 9 2 1 9 7 9 0 9 2
16 1 9 1 9 9 11 11 2 11 2 15 13 9 11 11 2
8 9 7 13 1 0 7 0 2
22 4 14 13 0 9 0 9 1 9 15 3 0 0 9 2 3 13 9 7 9 9 2
45 11 3 13 2 16 13 0 15 3 13 2 16 1 9 0 7 0 9 13 0 13 0 9 0 9 7 10 9 3 13 2 3 3 0 9 2 0 9 2 9 9 7 0 9 2
18 1 9 9 9 13 0 9 9 2 15 0 9 7 9 13 7 13 2
32 3 2 1 12 0 9 13 9 9 7 1 0 12 0 0 9 7 0 9 0 2 16 1 9 9 15 10 9 13 1 12 2
45 3 9 2 7 15 1 12 2 13 9 9 9 0 0 9 7 0 9 2 12 9 15 13 0 9 2 12 9 9 2 1 0 12 9 15 13 1 12 10 0 0 9 7 9 2
21 13 15 2 16 1 0 9 4 3 13 12 12 9 2 3 1 12 3 16 3 2
41 1 0 9 2 10 9 9 15 13 0 9 9 0 9 9 1 9 2 11 13 2 16 1 0 0 9 13 9 12 9 1 9 2 16 15 4 13 1 12 3 2
34 1 1 9 1 9 1 0 9 1 9 0 9 7 1 0 9 15 13 2 13 11 2 16 3 15 9 9 1 9 13 1 12 9 2
23 1 9 0 9 9 11 4 7 1 0 12 2 9 13 4 1 9 12 12 9 1 9 2
7 9 13 13 9 0 0 9
2 11 2
22 3 13 7 13 4 15 1 12 2 9 12 13 15 0 7 0 0 0 9 7 9 2
15 13 15 15 1 0 9 9 0 9 2 15 13 9 9 2
25 9 0 9 13 13 0 9 0 9 1 9 2 16 4 1 10 9 7 0 0 9 13 0 9 2
21 9 4 13 1 9 9 9 2 15 4 0 9 7 9 0 13 9 1 0 9 2
18 1 9 9 4 13 13 7 9 0 9 0 9 9 7 9 9 9 2
50 9 15 13 13 3 2 9 2 9 2 9 2 9 7 0 2 0 2 0 2 3 0 7 0 9 2 1 15 15 3 13 0 9 2 9 2 9 2 9 2 9 2 9 2 0 7 0 9 2 2
31 9 1 9 13 13 9 9 9 13 9 0 9 7 0 7 0 9 2 16 1 15 13 7 16 15 13 1 9 0 9 2
11 1 9 15 7 13 9 0 15 9 9 2
13 9 1 9 9 13 13 1 9 7 9 0 9 2
21 1 0 9 7 9 13 13 9 14 12 9 9 2 1 9 0 9 14 12 9 2
5 11 1 9 0 9
2 11 2
21 1 9 0 2 0 9 1 9 9 1 0 9 11 15 3 13 0 9 11 11 2
60 2 16 4 13 1 15 1 15 13 2 3 13 15 3 1 9 9 9 1 0 9 9 7 9 9 1 11 2 1 9 9 11 2 1 9 2 15 3 13 2 2 13 11 1 9 1 0 7 0 9 1 0 9 0 9 11 11 1 11 2
20 11 13 9 0 9 0 7 0 9 2 15 4 1 15 13 1 9 1 11 2
10 3 7 13 1 9 0 9 7 9 2
28 2 13 9 2 16 1 9 1 10 9 13 0 9 1 11 3 0 9 16 0 9 1 11 2 2 13 11 2
4 11 13 9 9
2 11 2
22 9 0 9 11 11 13 2 16 1 0 9 13 0 9 9 1 9 1 0 9 9 2
37 11 2 15 4 1 9 9 13 1 0 7 0 9 1 11 11 7 9 11 11 11 2 3 13 2 16 4 15 13 13 0 9 9 1 10 9 2
13 13 7 11 2 16 15 9 13 1 9 10 9 2
61 2 1 9 11 4 13 7 13 2 16 1 0 9 9 13 1 9 2 3 4 15 13 1 9 10 9 16 3 1 0 7 0 9 2 16 1 15 13 9 3 0 2 7 3 3 0 2 7 16 4 13 10 9 3 2 2 13 11 1 11 2
1 3
11 9 4 1 9 13 13 1 9 0 9 2
36 3 4 13 9 2 15 4 13 13 3 3 1 9 9 2 3 4 13 13 0 9 9 2 15 4 13 3 2 7 3 4 13 13 0 9 2
12 1 0 9 9 9 15 13 10 9 11 11 2
8 0 9 4 13 1 12 9 2
14 9 15 4 13 0 9 7 1 10 9 7 9 0 2
24 1 11 3 9 9 13 1 2 0 9 2 16 14 15 0 9 13 9 9 15 12 9 2 2
6 9 13 3 13 9 11
2 11 2
33 3 3 13 13 9 9 9 1 0 9 9 0 9 9 0 9 2 11 2 11 11 1 9 1 9 9 0 0 9 1 11 12 2
5 9 15 13 3 2
21 0 9 11 11 11 4 13 1 9 9 2 1 15 15 13 14 0 9 9 9 2
16 1 9 15 11 11 3 1 10 9 11 11 13 1 9 9 2
24 9 11 11 3 13 9 1 9 0 9 2 7 13 13 2 16 9 10 9 10 0 9 13 2
14 9 7 13 2 16 9 13 9 9 0 1 0 9 2
8 9 13 1 9 11 14 1 9
2 11 2
26 13 9 1 0 9 3 1 0 9 13 1 9 9 11 11 3 3 0 2 7 13 15 9 0 9 2
14 11 2 11 13 3 0 9 9 11 11 1 9 9 2
17 9 9 13 9 0 0 9 2 15 4 13 1 0 9 13 9 2
8 12 1 10 9 13 9 9 2
18 1 0 9 7 11 2 11 9 13 2 16 3 1 9 9 3 13 2
21 1 10 9 13 2 16 15 9 3 13 9 1 0 9 0 9 9 2 11 2 2
34 16 9 10 9 15 13 2 16 4 11 13 13 13 1 9 16 0 9 2 7 7 7 0 9 1 0 9 2 9 15 15 3 13 2
12 13 9 11 1 9 0 9 7 0 9 9 2
18 11 15 3 13 3 1 9 9 2 7 10 9 1 10 9 13 0 2
8 0 0 9 13 0 13 0 9
2 11 2
21 9 0 9 1 11 12 13 3 1 0 9 1 0 9 9 9 1 9 12 9 2
25 10 9 1 10 12 9 13 0 9 9 7 1 9 12 9 2 15 13 13 1 9 2 9 13 2
7 13 3 3 13 0 9 2
24 7 0 9 9 13 2 13 7 0 9 2 0 1 9 0 9 2 12 9 2 2 13 9 2
8 13 9 7 13 1 10 9 2
35 9 9 0 9 1 11 12 11 11 13 2 16 1 0 9 13 9 3 0 9 7 0 9 2 10 9 13 12 9 0 9 12 0 9 2
24 2 1 9 0 1 9 9 13 3 9 2 16 15 15 13 0 9 9 2 15 15 3 13 2
25 7 0 9 1 12 9 9 13 1 10 9 0 2 7 1 10 9 13 2 2 13 11 2 11 2
24 1 15 9 0 9 13 3 0 9 14 12 9 2 3 9 1 0 9 7 3 3 3 0 2
15 11 11 13 13 2 16 1 9 0 9 3 13 0 9 2
22 1 0 0 9 2 15 13 0 9 1 9 2 15 3 9 9 13 1 0 9 3 2
37 16 9 3 13 9 1 9 1 9 9 2 13 9 12 9 2 3 7 4 1 9 13 9 7 9 2 16 13 3 0 0 9 2 4 9 13 2
21 7 14 1 9 2 16 1 0 9 0 9 13 2 16 13 3 9 1 12 9 2
27 2 0 9 10 9 13 2 13 1 9 9 2 7 13 15 2 16 13 1 9 2 2 13 11 2 11 2
17 3 1 0 9 13 9 0 9 13 0 9 7 9 13 9 9 2
34 14 1 9 2 3 9 1 9 2 13 2 7 3 16 9 9 2 15 1 9 14 1 9 7 9 13 1 11 12 1 12 12 9 2
28 9 9 9 11 11 1 15 11 13 2 16 7 1 9 13 10 9 2 16 15 13 13 0 9 1 0 9 2
7 7 13 14 0 13 9 2
11 9 1 9 7 9 14 13 1 9 3 9
2 11 2
30 0 9 9 7 9 2 9 9 0 9 9 0 7 0 9 0 9 1 9 4 13 13 0 2 0 2 9 9 9 2
8 13 15 3 0 9 11 11 2
18 3 1 9 1 9 9 9 13 2 16 3 13 0 13 10 0 9 2
14 9 0 9 9 13 9 1 0 9 0 7 0 9 2
23 0 9 9 1 15 13 1 9 9 1 9 1 3 0 9 2 16 13 3 9 7 9 2
30 9 2 1 9 2 13 13 1 15 2 16 3 1 9 4 13 1 9 12 9 3 1 0 9 2 9 2 9 2 2
8 1 11 13 15 1 9 0 2
14 9 4 13 13 3 9 3 1 0 9 1 0 9 2
17 15 9 13 3 1 9 7 0 9 13 13 3 9 0 9 9 2
11 9 13 3 3 13 9 9 0 0 9 2
23 11 13 2 16 14 12 5 9 1 0 7 12 5 1 0 9 4 13 4 13 1 0 2
16 11 1 9 13 2 16 1 15 4 3 13 13 9 0 9 2
12 0 9 4 15 7 13 13 9 9 2 13 2
32 9 2 15 3 13 9 0 9 2 3 4 1 9 13 1 0 15 9 9 9 3 3 9 2 13 14 9 1 0 9 9 2
20 11 3 13 9 2 16 15 13 0 0 9 0 9 9 2 15 3 13 9 2
11 3 15 7 13 2 16 3 13 1 9 2
14 15 1 15 13 3 13 9 2 1 15 4 9 13 2
14 13 7 14 13 0 9 15 2 15 13 13 1 9 2
20 16 9 9 13 2 16 3 4 1 9 9 13 13 9 2 7 9 0 9 2
25 3 1 9 12 13 3 9 0 3 1 15 2 10 13 9 2 7 4 13 3 1 9 10 9 2
4 9 13 0 9
2 11 2
38 9 0 9 1 11 3 13 9 0 9 11 11 7 13 3 9 0 9 1 0 11 2 15 15 3 13 1 0 9 9 9 0 9 1 12 9 9 2
23 1 9 9 11 11 13 7 13 10 9 15 2 16 1 0 9 13 1 9 9 0 9 2
42 0 9 3 1 9 13 2 16 9 11 13 13 15 1 0 0 9 2 7 1 10 9 13 13 15 2 15 4 13 1 10 0 9 1 9 7 13 9 1 15 13 2
30 2 1 10 9 15 13 1 0 9 2 16 15 4 13 0 1 9 7 15 1 10 9 4 13 2 2 13 11 9 2
8 1 9 0 9 13 0 9 2
7 9 1 9 1 9 1 9
2 11 2
33 1 9 1 9 1 9 1 9 9 1 9 11 15 1 9 2 0 7 0 9 7 0 9 13 0 9 0 9 10 9 7 9 2
20 9 13 1 9 0 0 9 2 0 9 11 2 0 0 9 7 0 0 9 2
49 2 13 4 15 1 0 9 9 9 1 10 9 0 11 2 15 1 9 0 9 13 9 9 2 1 15 13 2 7 4 1 10 9 13 9 9 2 10 9 13 1 9 2 2 13 9 1 9 2
22 1 12 9 4 1 10 9 3 13 0 7 0 9 7 9 15 13 1 10 9 0 2
16 13 15 1 0 9 1 0 9 7 1 9 0 7 0 9 2
26 2 3 4 10 9 15 2 16 13 13 2 13 1 0 7 0 9 1 10 9 2 2 13 0 9 2
4 3 9 1 9
3 11 11 2
15 9 1 9 13 1 12 9 1 0 9 0 0 0 9 2
6 13 15 10 9 11 2
15 1 15 4 9 13 12 2 9 1 9 9 11 1 11 2
15 9 2 15 15 13 2 4 13 1 0 9 0 0 9 2
17 1 1 15 2 16 13 0 9 1 9 1 9 2 13 4 13 2
10 1 0 9 13 9 0 9 0 9 2
22 13 4 0 9 9 1 9 2 0 9 9 7 9 0 0 9 9 0 1 0 9 2
4 9 13 0 9
2 11 2
50 9 0 1 0 9 13 9 9 1 12 9 9 2 15 13 13 0 9 0 9 1 9 0 0 2 0 2 11 2 0 9 7 9 9 13 2 16 9 9 7 9 10 0 9 1 9 13 13 0 2
7 13 1 15 3 0 9 2
27 11 11 16 9 9 0 2 0 2 11 2 13 3 12 2 9 1 12 9 9 9 0 1 12 9 9 2
29 9 13 0 12 2 9 7 9 13 13 0 9 1 9 0 2 15 15 7 1 9 1 0 9 13 2 13 9 2
27 1 1 15 13 9 0 2 0 2 11 2 1 9 9 10 9 2 0 9 7 0 0 0 9 11 11 2
21 9 7 13 2 16 9 13 1 9 7 16 13 0 9 1 15 2 16 3 13 2
33 1 0 9 0 9 15 1 0 9 13 2 16 1 10 9 2 1 15 13 10 9 13 16 9 2 13 0 9 1 9 0 9 2
5 9 13 9 0 9
4 11 2 11 2
40 0 9 0 9 7 9 1 11 2 15 13 0 9 11 13 1 0 9 1 12 2 9 9 9 2 1 9 9 11 11 7 0 9 9 7 9 0 9 13 2
28 1 9 0 0 9 15 9 0 9 7 0 9 13 1 0 9 7 3 1 0 9 2 9 7 0 9 9 2
13 2 13 0 9 7 9 1 9 9 9 15 9 2
29 13 0 9 1 9 9 9 9 10 9 1 9 7 9 2 2 13 15 9 9 2 1 15 13 10 9 3 0 2
1 9
30 9 11 9 2 3 3 9 11 2 1 9 3 12 9 2 11 7 11 2 15 13 1 9 0 9 7 13 15 9 2
28 0 0 9 15 7 13 2 16 9 0 1 9 13 1 9 14 9 9 9 2 1 15 15 1 10 9 13 2
15 1 9 1 9 13 9 0 9 0 2 0 7 3 0 2
15 13 11 1 0 9 1 0 9 7 11 1 0 0 9 2
17 1 9 12 15 0 13 2 16 9 9 15 11 13 1 0 9 2
18 0 9 2 13 1 11 7 11 2 10 9 4 13 7 1 10 9 2
20 13 10 9 2 16 13 9 2 13 2 16 10 1 9 0 9 13 0 9 2
41 9 13 9 2 15 15 0 13 0 9 2 15 15 13 2 16 9 13 7 3 13 13 1 12 0 9 0 9 7 16 15 2 0 0 9 13 3 1 0 9 2
50 13 4 9 1 9 0 9 2 13 3 1 9 9 2 13 15 7 13 15 1 2 0 9 2 2 15 3 1 2 0 9 9 2 13 2 0 9 2 1 15 13 0 13 1 9 9 0 9 2 2
9 11 9 13 3 0 9 0 9 2
2 3 2
5 1 11 7 11 2
4 3 3 3 2
18 6 7 2 16 13 15 14 9 1 9 2 1 0 9 7 1 9 2
14 1 12 1 15 2 15 0 2 15 3 11 9 13 2
38 15 3 13 1 0 9 1 9 7 9 2 13 3 1 9 16 0 9 9 2 7 13 7 7 1 9 0 9 2 1 15 13 0 9 2 0 9 2
21 15 15 13 7 3 2 13 2 3 16 3 2 9 16 9 9 2 7 0 9 2
44 13 2 16 0 9 1 0 9 3 1 9 10 0 9 13 2 0 9 13 7 13 15 16 0 7 13 2 3 7 1 0 7 0 9 2 16 15 1 15 13 15 9 9 2
16 13 2 16 9 9 13 7 9 2 7 9 2 7 0 9 2
34 15 15 13 9 2 13 15 2 16 4 16 15 1 9 1 0 9 10 9 13 1 9 0 9 7 3 13 2 3 1 15 9 13 2
23 9 13 0 9 0 9 2 9 1 11 3 9 1 9 15 2 15 13 1 9 9 13 2
4 9 13 0 9
9 9 0 9 3 13 3 0 12 9
2 11 2
20 0 9 2 15 13 14 1 0 9 9 1 0 9 9 2 15 13 13 9 2
20 0 9 1 9 0 9 9 9 13 1 9 0 9 1 9 11 7 0 9 2
17 0 7 0 9 2 11 2 13 9 0 9 13 1 9 9 12 2
20 1 9 15 13 14 12 9 2 16 3 13 1 0 9 9 14 12 0 9 2
27 1 9 1 0 9 7 11 3 13 9 2 3 9 13 1 0 9 9 1 9 2 7 3 9 0 9 2
9 15 13 9 9 11 11 13 3 2
29 3 9 1 9 13 2 16 9 4 13 1 9 2 1 15 15 13 9 2 13 15 15 1 12 9 9 1 9 2
37 1 0 9 13 9 0 0 9 1 9 2 9 1 9 9 7 9 1 0 9 2 1 0 9 2 9 2 9 2 9 9 3 2 3 9 11 2
13 3 7 3 1 9 11 2 0 0 9 7 11 2
16 9 1 9 11 7 11 15 3 13 13 9 0 9 10 9 2
32 16 4 15 1 9 13 13 0 9 2 13 9 9 1 9 3 2 7 13 9 0 9 2 1 10 9 13 9 3 13 9 2
15 11 13 0 9 9 1 15 10 0 9 1 9 0 9 2
17 7 9 10 9 15 13 9 4 13 1 15 1 3 12 0 9 2
18 3 16 1 0 12 0 9 13 9 13 0 9 0 11 7 0 11 2
9 7 10 9 13 1 0 9 9 2
35 0 9 13 0 9 1 0 9 1 9 0 9 1 9 0 9 2 11 3 13 0 9 1 0 9 7 0 9 10 9 13 1 0 9 2
9 0 11 13 3 1 9 12 9 9
2 11 2
16 0 0 9 11 9 13 1 9 1 9 12 9 12 9 9 2
14 10 9 11 9 10 9 3 13 7 13 15 1 9 2
14 1 10 0 0 9 9 13 1 9 3 16 12 9 2
14 13 2 16 11 13 3 0 9 1 9 12 9 9 2
19 0 9 3 13 1 12 9 1 0 9 2 15 13 14 1 12 9 9 2
19 1 9 11 3 9 14 1 9 1 10 9 13 3 12 7 12 9 9 2
33 9 3 13 9 2 1 15 10 9 13 0 9 1 11 2 11 2 12 9 9 1 9 9 2 15 9 13 0 9 11 11 11 2
11 9 11 13 9 1 9 1 12 9 9 2
16 15 9 1 9 11 9 4 13 13 1 9 1 9 3 13 2
16 9 11 3 13 1 9 9 2 15 13 0 9 11 2 11 2
22 13 1 15 2 16 13 13 9 9 11 9 1 0 9 2 16 13 1 9 0 9 2
19 0 9 3 13 9 2 16 4 11 9 13 1 10 9 13 16 0 9 2
9 0 9 7 9 13 9 1 9 9
2 11 2
27 0 9 0 1 9 0 7 0 9 13 3 0 0 9 0 9 0 9 7 0 9 11 11 7 11 11 2
26 9 2 10 9 13 13 0 9 9 9 2 13 13 9 9 2 3 13 9 9 1 0 7 0 9 2
38 11 7 11 3 13 2 16 9 9 9 13 9 0 0 9 2 12 9 3 1 0 7 12 9 1 0 9 2 4 3 13 9 7 3 0 9 9 2
19 2 9 15 3 13 13 2 16 13 9 1 15 9 2 2 13 9 11 2
20 1 15 13 9 13 16 9 0 9 9 2 7 16 0 9 13 0 9 9 2
30 2 13 15 16 9 1 9 2 3 15 13 15 13 2 16 15 13 13 0 9 2 16 3 13 9 2 2 13 11 2
11 9 4 1 15 3 13 13 9 12 9 2
9 3 3 4 0 9 13 1 9 2
18 15 1 9 9 13 1 12 12 9 1 0 9 7 12 12 1 9 2
12 1 11 13 9 9 13 3 1 12 9 9 2
8 15 13 1 11 3 12 9 2
38 2 1 0 9 13 7 9 3 0 2 1 0 0 9 3 16 12 9 9 0 9 2 0 9 2 15 9 13 14 12 12 2 2 13 15 9 11 2
20 12 9 13 2 16 9 13 1 9 9 2 10 0 9 1 9 1 9 2 2
8 13 15 3 13 3 9 9 2
5 0 9 13 1 11
3 0 11 2
25 0 9 0 0 9 0 11 7 0 9 0 9 13 3 1 12 1 9 2 0 9 1 12 9 2
27 11 13 1 9 1 0 9 9 2 12 11 0 9 2 11 3 13 9 9 11 2 12 7 9 0 9 2
15 2 13 4 3 13 2 2 13 11 1 9 9 11 11 2
16 2 13 15 3 10 0 9 7 3 15 9 13 15 1 11 2
6 3 15 15 13 15 2
13 16 15 15 3 13 2 13 4 3 16 9 9 2
13 1 9 0 9 13 1 3 0 9 10 9 2 2
14 7 1 15 7 13 2 16 12 1 11 13 0 9 2
13 13 16 9 2 0 9 15 13 12 9 1 9 2
4 0 9 11 13
2 11 2
37 13 3 0 1 15 2 15 11 11 13 1 9 12 9 7 1 9 2 13 1 9 1 0 9 0 9 1 0 2 0 9 9 0 9 11 11 2
5 2 13 0 9 2
9 13 9 7 3 9 2 2 13 2
21 16 13 1 0 9 0 9 2 4 1 11 1 11 2 3 13 3 0 9 2 2
15 1 9 9 0 9 9 11 3 13 2 10 0 9 2 2
17 2 0 9 13 2 16 13 13 1 0 9 2 7 15 3 13 2
18 13 15 1 15 3 13 7 13 15 3 1 9 9 2 2 13 11 2
4 0 9 1 11
2 11 2
20 0 0 9 9 13 3 1 0 0 9 11 0 9 1 9 1 9 0 9 2
28 9 0 9 1 9 0 9 13 9 7 9 11 11 2 10 0 9 9 2 9 2 9 4 3 13 1 11 2
33 0 9 1 0 0 9 13 9 9 0 9 9 2 9 2 11 11 2 2 0 9 1 0 9 13 11 11 7 0 9 11 11 2
4 3 1 9 12
6 11 15 13 13 0 9
2 11 2
15 0 9 11 11 11 11 13 3 0 9 0 9 0 11 2
20 2 3 9 13 2 16 3 13 0 9 1 9 2 7 15 10 9 3 13 2
17 13 2 16 16 4 12 12 9 3 13 2 13 15 15 15 13 2
3 7 3 2
20 15 14 3 14 2 2 13 3 11 2 15 1 0 9 3 13 7 0 11 2
8 9 1 11 2 11 1 9 12
5 1 11 13 0 9
2 11 2
21 1 0 11 2 9 11 2 11 2 4 1 9 13 1 0 9 0 9 1 11 2
22 1 0 9 4 13 12 9 9 2 13 11 2 11 11 2 9 9 0 9 11 9 2
20 9 9 2 15 13 4 13 1 0 9 1 9 2 13 12 12 9 9 3 2
23 16 9 15 4 13 3 0 9 1 9 1 12 9 2 15 3 13 1 12 12 9 9 2
14 1 10 9 9 13 0 9 1 9 1 12 12 9 2
6 11 2 11 1 0 9
2 11 2
14 9 0 0 9 11 2 11 13 13 10 9 1 11 2
21 16 3 13 9 0 11 2 9 13 13 2 0 9 9 0 9 7 0 9 2 2
18 0 9 10 9 13 9 11 11 7 10 10 9 1 9 9 10 9 2
11 0 9 4 13 0 0 9 12 2 9 2
25 1 9 10 9 3 13 1 9 9 0 9 1 10 0 0 9 2 15 15 9 11 2 11 13 2
4 0 9 11 13
2 11 2
18 0 0 9 0 9 11 4 1 0 9 9 13 14 1 12 2 9 2
8 0 0 9 13 9 7 9 2
13 0 9 1 0 9 4 13 14 1 0 0 9 2
11 1 9 12 13 9 11 9 12 9 9 2
17 9 13 1 9 9 9 1 9 1 9 9 1 9 12 9 9 2
23 9 9 11 2 15 13 1 9 12 1 12 9 0 1 11 7 9 2 13 12 9 9 2
4 0 11 13 9
2 11 2
23 1 0 9 12 9 9 13 0 9 0 0 9 11 2 16 3 3 13 9 12 9 9 2
9 3 15 13 9 9 11 11 11 2
24 9 13 11 1 9 12 1 12 9 1 12 9 2 9 1 9 1 12 9 2 1 9 12 2
10 11 13 1 10 9 0 9 12 9 2
6 1 12 5 9 13 2
17 0 9 11 13 0 13 1 9 2 9 2 9 9 7 0 9 2
3 0 9 13
2 11 2
26 0 9 2 9 0 11 9 2 3 1 0 9 2 11 1 11 2 13 1 9 14 12 9 0 9 2
14 13 15 15 3 9 1 9 9 2 9 1 9 3 2
15 9 1 3 0 9 7 3 0 9 13 1 9 12 9 2
1 3
31 9 0 9 1 11 15 1 9 3 13 1 12 9 2 16 13 1 9 3 16 12 0 9 1 9 2 12 9 0 9 2
4 9 9 3 13
4 11 2 11 2
23 9 9 2 15 1 0 12 9 13 1 0 9 1 9 12 2 15 3 3 1 9 13 2
18 3 15 7 13 0 9 2 3 16 15 3 1 0 9 13 0 9 2
12 3 1 9 15 9 1 11 13 1 12 9 2
10 1 0 9 15 3 13 9 12 9 2
11 1 9 3 9 1 11 13 1 12 9 2
24 1 9 0 9 13 3 9 3 0 0 9 7 1 9 0 9 11 1 11 0 9 15 13 2
23 16 3 11 13 12 1 9 2 13 15 2 16 3 3 15 9 3 13 14 9 12 9 2
4 9 1 9 11
2 11 2
21 0 0 9 9 11 2 0 1 9 0 9 12 9 9 2 15 3 13 1 11 2
15 9 13 9 9 9 2 13 0 0 9 7 13 9 9 2
14 1 0 9 13 1 9 9 0 9 3 1 0 9 2
12 0 9 13 13 9 9 0 9 1 9 9 2
25 0 9 1 9 0 9 13 10 9 9 2 11 11 2 0 9 9 11 2 15 13 0 0 9 2
12 9 13 9 0 9 9 11 9 2 11 11 2
13 1 10 9 1 9 7 13 14 1 10 0 9 2
17 16 13 11 0 9 11 2 9 9 9 11 13 1 0 9 13 2
11 9 0 9 11 13 13 3 0 9 9 9
7 0 2 11 15 13 9 11
2 11 2
19 9 0 2 11 15 13 9 1 0 9 9 12 9 9 11 11 2 11 2
17 9 1 15 13 1 9 1 9 0 9 2 15 9 14 3 13 2
9 3 15 13 0 9 11 11 11 2
36 13 1 10 9 2 16 9 0 2 11 3 13 1 9 9 9 3 1 0 0 9 2 0 9 11 11 11 7 3 1 9 11 1 0 9 2
10 9 13 1 10 9 13 16 0 9 2
17 11 4 13 1 0 0 9 1 9 12 1 0 9 12 9 9 2
19 0 9 13 3 13 1 9 7 9 1 0 2 0 2 0 7 0 9 2
6 0 9 1 9 0 9
32 3 1 9 13 10 9 3 7 1 9 15 2 16 15 0 9 9 0 7 0 11 13 1 0 9 1 9 0 7 0 9 2
28 9 2 11 15 13 2 1 9 1 10 0 9 0 9 2 3 1 9 12 13 9 0 0 9 2 9 2 2
21 7 3 11 13 3 16 0 9 9 0 9 10 9 1 9 0 7 9 0 9 2
38 7 3 13 0 9 15 13 2 7 0 0 0 9 1 9 13 1 9 12 3 1 9 0 1 9 1 0 9 7 1 3 16 12 1 9 1 0 2
17 13 15 3 1 0 9 12 0 0 9 2 0 1 0 12 9 2
44 3 1 0 9 13 0 2 16 9 12 13 9 2 0 0 9 9 2 13 3 9 0 11 7 9 2 0 1 9 0 0 9 2 10 9 15 13 3 3 1 0 9 2 2
34 1 0 9 13 9 2 0 0 2 2 0 2 2 9 0 9 1 0 9 2 15 2 13 2 9 2 9 2 9 9 7 0 9 2
40 0 9 0 9 9 15 13 1 15 2 16 0 9 13 13 3 1 9 9 0 7 0 9 2 0 0 9 2 0 0 9 2 3 3 10 0 0 9 2 2
17 7 3 1 10 9 13 0 9 2 16 13 9 2 1 9 9 2
33 15 13 3 12 1 9 2 3 10 0 9 1 9 13 1 0 9 3 0 9 9 0 9 2 16 9 1 0 9 13 3 0 2
37 13 3 2 16 0 0 9 2 0 1 11 1 9 0 9 9 7 1 11 1 9 9 0 9 2 0 3 1 0 0 9 2 13 1 9 9 2
15 11 13 1 0 9 0 9 2 16 15 1 0 9 13 2
17 13 15 3 1 0 9 1 9 9 9 1 0 9 1 9 9 2
31 0 9 1 9 2 13 2 14 15 13 0 9 1 0 9 2 7 0 9 0 9 7 13 10 9 1 9 0 0 9 2
23 0 9 1 9 0 9 13 3 1 9 2 16 10 0 9 4 13 3 1 9 9 9 2
28 0 9 13 9 9 9 7 9 9 0 15 9 2 16 7 0 9 2 15 13 3 0 1 9 9 7 9 2
30 3 13 13 9 1 9 1 0 9 3 2 13 2 14 1 9 0 9 2 16 13 15 1 13 7 3 9 10 9 2
41 13 2 14 1 9 0 9 0 9 2 3 13 1 9 0 2 3 3 0 9 2 15 4 1 0 9 13 2 9 2 16 7 3 3 13 13 0 9 0 9 2
14 3 2 9 0 7 0 13 0 9 1 9 10 9 2
30 13 7 9 2 16 3 9 1 9 9 13 3 0 2 7 16 3 3 13 7 4 13 7 1 9 0 9 2 0 2
42 1 10 0 9 13 9 2 0 10 0 9 9 2 16 0 9 9 13 0 1 9 9 1 0 9 2 7 16 7 13 13 3 7 0 3 2 0 9 1 9 9 2
21 13 1 15 2 16 10 9 13 14 1 0 9 2 7 16 7 3 13 3 13 2
10 0 13 2 16 0 9 3 3 13 2
16 10 0 9 15 13 2 9 9 15 13 2 7 13 3 0 2
35 0 9 15 3 13 2 7 9 2 9 0 9 2 9 0 9 2 9 9 1 0 9 2 0 9 9 3 2 2 15 13 14 3 3 2
28 0 9 2 9 9 2 9 1 9 7 9 2 15 13 9 2 3 3 13 13 9 2 0 1 0 0 9 2
15 0 9 2 15 0 9 13 1 9 0 9 2 13 0 2
14 13 1 9 9 13 7 14 9 2 7 3 7 9 2
21 13 1 15 2 13 9 1 9 3 0 0 9 2 16 4 0 9 13 7 13 2
9 9 0 9 2 11 11 2 12 2
10 11 11 11 13 12 1 0 9 9 2
9 0 9 1 9 13 1 9 12 2
17 4 15 13 1 2 9 0 7 0 9 9 0 7 0 9 2 2
25 10 9 15 11 2 11 13 0 10 9 7 0 9 1 15 13 9 7 0 9 1 0 9 9 2
15 15 4 3 3 13 16 9 0 9 7 3 0 0 9 2
12 11 11 15 13 12 2 9 12 1 9 11 2
25 1 9 0 0 0 11 1 9 2 12 13 1 9 1 9 1 11 2 3 9 12 13 9 9 2
12 9 9 13 1 9 2 12 1 9 1 11 2
9 1 9 0 9 15 13 0 9 2
15 3 13 1 9 1 11 2 3 3 1 9 1 0 11 2
16 1 0 12 9 15 3 1 11 13 2 3 7 1 0 9 2
26 1 0 9 13 0 9 11 1 11 1 0 11 7 9 11 11 2 11 11 11 1 11 2 9 11 2
37 0 9 7 9 1 9 7 1 9 13 11 2 11 0 9 14 1 0 0 9 2 7 7 1 0 9 2 15 13 1 9 7 9 10 0 9 2
32 1 9 10 9 1 9 0 9 13 11 2 11 13 0 0 9 11 2 11 2 15 0 9 2 16 13 2 3 13 10 9 2
29 13 2 16 0 1 10 9 2 3 1 0 9 7 0 9 2 13 0 13 16 0 9 2 9 7 9 0 9 2
29 13 15 3 3 11 2 11 2 15 1 9 10 9 13 2 16 11 2 11 15 9 0 9 13 1 10 0 9 2
11 11 2 11 10 9 0 9 13 10 9 2
34 0 10 9 1 9 0 9 2 15 13 3 1 0 9 0 2 13 9 7 9 0 0 9 1 9 0 9 2 0 9 7 0 9 2
27 0 9 9 0 9 1 10 9 2 3 0 0 0 9 2 13 9 13 2 3 3 13 0 9 0 9 2
15 2 1 9 1 0 9 2 0 2 3 4 13 13 2 2
46 0 9 2 15 16 9 9 7 9 13 3 1 10 0 9 7 13 15 13 10 9 7 9 2 13 3 9 0 9 7 13 13 1 15 2 16 4 3 10 9 13 1 9 0 9 2
22 9 9 0 9 13 0 9 9 1 0 0 9 2 15 13 15 0 9 0 0 9 2
21 0 9 0 9 13 9 9 2 15 13 9 0 0 7 0 9 1 9 10 9 2
65 0 9 9 0 9 2 15 16 0 9 13 9 1 9 9 1 9 2 9 7 0 9 0 9 2 13 0 9 9 0 9 2 3 2 9 0 0 9 2 3 15 0 9 13 0 9 2 16 9 9 13 9 0 2 10 9 3 13 0 9 7 13 1 9 2
39 0 9 10 9 9 13 2 16 9 1 9 0 0 9 7 2 9 9 2 0 7 0 9 4 13 1 15 13 1 0 7 3 3 0 2 0 9 2 2
22 0 9 9 0 9 2 1 15 11 2 11 13 3 2 15 13 9 0 7 0 9 2
18 3 1 9 2 12 13 13 9 9 0 9 7 0 9 1 9 9 2
20 9 0 9 1 12 9 13 4 13 7 13 1 0 9 2 1 15 15 13 2
44 10 0 9 1 9 9 9 3 11 2 11 13 1 0 0 9 2 1 15 0 0 9 13 13 9 0 0 9 9 1 9 2 15 0 9 13 2 16 15 9 1 9 13 2
45 0 9 13 9 0 9 7 9 9 9 2 15 4 13 9 1 9 2 15 13 0 1 9 9 1 0 7 0 9 7 9 2 7 9 2 16 0 9 9 4 13 0 0 9 2
16 10 9 13 11 2 11 1 0 9 9 9 0 9 7 9 2
26 0 9 10 9 13 0 9 2 15 14 16 13 0 7 0 9 2 7 13 3 0 9 0 9 9 2
28 1 9 10 9 13 11 2 11 0 9 0 9 2 1 15 13 9 0 9 10 0 9 1 9 9 0 9 2
33 10 9 1 9 0 9 4 3 13 0 9 11 11 2 12 2 2 9 0 9 9 1 11 7 11 7 0 9 1 0 0 9 2
12 11 11 15 13 12 2 9 12 1 9 11 2
9 10 11 13 12 1 0 9 9 2
9 0 9 1 9 13 1 9 12 2
6 0 9 13 10 9 2
36 0 10 9 1 0 2 9 0 9 2 15 13 3 1 0 9 0 2 13 9 7 9 0 0 9 1 9 0 9 2 0 9 7 0 9 2
27 0 9 9 0 9 1 10 9 2 3 0 0 0 9 2 13 9 13 2 3 3 13 0 9 0 9 2
14 2 1 9 1 0 9 0 2 3 4 13 13 2 2
47 0 9 2 15 16 9 9 7 9 13 3 1 10 0 9 7 13 15 13 10 9 7 9 2 13 3 9 0 9 7 13 13 1 15 2 16 4 3 3 10 9 13 1 9 9 0 2
5 11 1 9 0 9
2 11 2
28 11 13 0 9 9 1 9 9 0 9 0 9 3 1 9 2 16 9 9 9 0 9 7 9 1 9 13 2
16 16 4 9 10 9 13 2 13 0 9 1 0 9 0 9 2
7 13 15 3 0 9 11 2
37 0 9 1 9 13 2 16 9 0 1 0 9 13 9 9 1 12 9 9 2 15 4 13 13 0 9 0 9 1 9 0 11 2 11 2 11 2
21 0 9 7 9 9 13 2 16 9 9 7 9 10 0 9 1 9 13 13 0 2
16 1 9 11 0 9 13 14 1 9 2 3 13 9 9 13 2
8 1 0 9 13 10 9 13 2
22 0 9 13 9 13 1 0 0 9 0 9 7 1 9 1 9 7 10 9 2 13 2
8 9 0 9 15 3 13 1 9
1 9
2 11 2
10 9 0 9 15 3 13 1 12 9 2
15 9 13 1 0 0 9 1 12 9 7 9 1 12 9 2
14 9 0 9 0 9 13 1 0 9 0 12 9 9 2
14 9 12 9 9 4 13 1 9 1 9 0 0 9 2
26 9 1 9 11 2 0 9 0 9 2 13 10 9 1 12 9 9 7 1 0 9 1 12 9 9 2
21 3 0 9 12 9 9 13 10 9 1 9 1 11 7 12 9 9 1 0 9 2
22 1 12 9 9 13 0 0 9 3 1 0 9 1 0 9 2 1 9 9 0 11 2
13 0 0 9 0 9 13 1 9 12 3 3 11 2
4 9 9 13 4
2 11 2
23 16 0 9 1 9 1 11 13 9 1 0 9 1 9 12 2 9 9 0 9 15 13 2
28 13 15 3 1 10 0 9 0 0 9 0 9 2 7 1 9 3 13 15 0 9 1 0 9 0 0 9 2
31 0 9 9 15 1 9 13 1 12 9 7 1 0 9 3 13 1 9 1 0 9 1 12 9 2 15 13 0 9 9 2
9 9 7 13 1 0 9 0 9 2
15 13 15 3 9 9 9 7 0 9 2 0 0 0 9 2
16 3 0 9 0 9 15 13 13 0 9 1 9 10 0 9 2
31 9 9 3 1 0 9 9 13 9 0 9 2 1 15 3 1 10 0 9 9 9 13 4 7 0 9 9 13 9 3 2
3 0 9 9
2 0 9
18 9 9 0 9 11 11 1 9 1 9 12 15 3 3 13 1 9 2
15 9 7 0 9 0 9 15 13 3 1 10 9 0 9 2
21 9 9 11 11 13 0 9 10 9 2 0 9 7 0 9 2 15 13 9 9 2
12 13 1 15 0 9 1 0 9 13 0 9 2
39 15 15 1 15 13 2 13 7 13 13 2 16 13 13 1 0 9 2 3 0 2 15 15 13 2 3 2 3 7 3 7 3 2 3 2 2 7 3 2
34 13 9 3 13 13 9 1 9 0 9 2 16 4 15 13 1 9 2 16 4 13 3 9 7 10 9 2 7 13 13 1 0 9 2
40 1 0 9 9 1 0 9 13 9 11 2 9 1 3 0 9 2 0 9 2 16 15 13 3 15 13 10 9 2 13 3 1 0 9 7 15 0 15 13 2
25 16 10 9 13 3 3 7 3 0 9 0 9 1 9 15 3 13 7 1 9 2 15 13 13 2
20 7 3 13 0 2 13 1 9 9 9 2 1 15 7 13 13 9 0 9 2
29 7 7 1 9 13 1 15 3 9 7 0 9 2 16 4 1 0 9 2 7 3 1 9 2 13 1 0 9 2
10 15 4 15 3 13 1 10 9 13 2
15 0 9 11 11 13 9 0 9 7 3 3 9 11 13 2
8 15 13 1 9 9 11 11 2
12 13 13 1 0 9 0 9 9 7 9 13 2
11 9 9 13 3 0 9 7 9 11 13 2
18 11 11 13 15 0 16 15 13 9 0 9 2 7 15 9 13 9 2
8 1 9 15 14 13 1 9 2
40 7 0 9 2 9 2 11 2 3 7 3 13 1 10 9 0 9 9 13 10 9 9 1 11 11 1 9 2 16 3 15 3 13 15 9 1 9 10 9 2
6 13 15 0 0 9 2
12 0 9 9 9 11 11 13 7 10 9 13 2
4 9 9 13 11
16 1 9 13 1 0 9 9 2 13 9 9 11 11 2 11 2
64 16 10 9 1 0 9 13 2 16 0 9 3 13 1 9 9 1 9 0 9 1 0 9 2 12 1 0 9 0 0 9 11 11 2 11 2 7 9 1 0 15 9 11 11 13 2 16 0 9 13 9 3 1 12 9 1 0 9 2 7 15 11 11 2
38 1 11 2 11 15 11 2 13 2 1 0 0 0 9 2 15 0 9 1 9 0 0 9 1 11 7 1 9 1 9 0 0 9 1 11 3 13 2
38 15 15 13 11 2 0 9 13 1 11 11 1 9 9 2 3 0 9 1 9 0 0 9 2 7 15 1 9 1 9 1 12 1 12 9 1 9 2
42 3 2 1 9 9 0 0 15 9 0 9 2 0 9 10 9 7 3 0 0 9 9 13 13 0 9 0 7 10 9 1 0 9 1 11 13 1 12 7 12 9 2
12 0 9 1 9 9 11 13 11 0 11 11 2
31 9 0 9 13 1 10 9 0 9 14 1 9 10 9 7 10 9 4 15 13 3 13 1 9 1 12 7 1 12 9 2
12 9 7 9 13 9 14 1 12 9 1 9 2
28 11 11 15 3 16 9 0 13 1 9 2 16 1 9 9 1 0 9 1 9 13 9 0 9 0 9 3 2
29 0 9 4 1 10 9 13 7 1 9 9 1 9 2 16 0 9 13 1 0 0 9 1 9 3 1 0 9 2
51 2 7 16 13 1 9 2 16 0 9 13 3 0 9 7 16 11 13 0 7 0 9 2 3 13 9 0 9 1 9 1 9 3 3 13 2 2 13 11 11 7 13 2 16 3 15 15 13 9 9 2
13 2 9 1 0 0 9 3 3 13 10 9 2 2
9 0 9 15 3 3 3 13 1 11
2 11 2
16 0 0 9 0 9 1 0 11 15 13 1 9 9 7 9 2
23 1 9 1 9 9 0 0 9 1 11 15 13 9 0 9 0 9 0 9 11 11 11 2
19 1 9 9 15 0 9 13 13 1 0 9 9 7 9 7 1 9 9 2
14 9 9 0 9 1 11 13 3 1 11 2 11 0 2
21 11 3 13 13 9 1 0 7 0 11 2 7 13 3 10 9 3 1 0 11 2
16 1 9 4 15 13 3 9 1 0 9 1 9 0 9 13 2
26 9 0 2 0 9 1 0 12 9 0 9 13 0 12 9 9 7 1 0 9 12 13 12 9 9 2
20 0 0 9 11 2 15 13 0 0 9 2 13 10 9 1 9 7 1 11 2
11 10 9 13 13 9 1 11 7 0 9 2
11 3 13 1 11 9 12 9 1 12 9 2
12 9 0 9 13 2 7 9 10 9 3 13 2
14 3 13 13 1 9 3 3 16 1 9 7 1 9 2
9 13 2 14 9 2 13 13 7 9
15 0 9 4 13 9 13 13 0 9 7 13 0 9 0 9
15 3 0 1 15 15 3 3 13 1 0 9 1 0 9 2
13 16 4 9 13 9 9 2 13 13 13 10 9 2
19 1 15 0 9 13 0 9 9 2 1 0 9 14 1 0 9 1 9 2
28 1 9 4 15 13 2 3 3 13 0 13 1 0 9 1 9 12 12 9 2 0 1 9 1 9 0 9 2
18 1 9 0 9 0 1 9 15 9 9 13 2 1 15 4 9 13 2
28 1 9 2 15 13 1 0 9 2 13 9 1 0 9 1 9 7 9 1 9 0 9 3 9 1 0 9 2
33 13 1 15 9 1 9 9 14 0 16 12 9 2 9 1 9 9 9 2 0 7 0 9 2 7 9 0 9 0 3 12 9 2
17 16 0 9 13 9 13 0 9 1 0 9 7 9 1 9 9 2
16 0 9 4 9 13 1 9 9 1 0 9 7 1 0 9 2
28 15 7 13 3 13 0 9 2 0 9 1 9 1 9 9 2 3 0 9 2 0 9 7 9 1 0 9 2
12 0 9 15 13 7 1 10 0 9 9 9 2
13 16 9 13 9 1 12 9 2 13 9 12 9 2
15 1 9 1 12 1 12 9 13 9 3 1 9 12 9 2
13 1 9 1 12 9 3 4 0 9 13 12 9 2
21 1 0 9 9 13 1 9 3 12 9 2 9 1 12 9 9 13 3 12 9 2
29 1 9 1 9 13 9 13 1 0 9 1 0 9 2 15 7 13 13 3 1 9 2 9 2 9 7 9 9 2
30 7 16 13 9 10 9 13 7 13 15 13 1 0 0 9 2 0 9 13 1 15 0 16 1 9 1 9 1 9 2
30 3 9 1 0 9 0 1 12 9 13 9 0 9 1 9 12 9 2 1 12 9 12 9 7 1 12 9 12 9 2
48 1 9 9 9 9 13 1 0 9 1 9 7 0 0 9 2 15 15 13 3 13 2 3 9 9 7 9 0 1 9 2 9 0 9 2 0 9 1 9 0 2 9 9 7 9 0 9 2
36 0 9 2 0 0 0 9 2 1 9 12 2 12 7 12 9 7 1 0 9 12 9 13 9 13 1 0 9 0 9 3 1 9 0 9 2
18 10 9 13 1 9 0 7 0 9 2 9 1 0 9 7 0 9 2
22 1 9 0 9 13 13 9 1 9 12 12 7 12 9 9 3 1 10 9 7 9 2
18 1 9 9 13 3 0 9 9 7 9 9 2 15 15 13 1 9 2
9 9 13 13 12 9 9 0 9 2
29 9 2 15 13 1 0 9 1 9 9 2 13 13 3 13 2 16 13 1 9 0 1 9 7 16 13 10 9 2
14 9 1 9 1 9 1 9 13 0 16 1 0 9 2
30 0 13 9 1 9 9 2 15 13 13 0 16 12 9 2 3 9 9 7 9 7 9 1 9 9 1 0 12 9 2
20 9 9 2 3 9 13 1 9 9 2 13 1 9 0 9 12 0 9 0 2
14 3 15 9 13 1 0 9 0 1 9 7 0 9 2
22 3 13 13 0 9 2 1 0 9 13 0 13 0 9 7 2 1 9 2 13 9 2
17 0 9 7 9 0 9 13 14 0 9 2 16 13 15 0 9 2
12 1 9 0 9 13 13 0 9 0 9 9 2
9 9 0 9 13 9 9 1 9 2
16 13 13 0 0 0 9 0 0 9 7 13 0 9 0 9 2
13 1 9 15 15 13 0 9 7 9 9 0 9 2
13 0 9 9 13 9 0 9 13 1 0 0 9 2
22 16 4 0 9 9 13 2 4 9 3 15 13 1 9 0 0 9 1 0 0 9 2
4 11 13 11 9
8 1 11 13 3 11 2 3 11
3 0 11 2
16 3 1 12 0 9 0 11 13 10 9 0 9 1 0 9 2
28 11 15 13 9 1 12 9 0 11 1 11 2 11 1 0 11 11 1 11 7 3 3 11 1 11 1 11 2
22 9 0 11 11 11 13 12 9 0 9 11 7 3 1 10 9 13 1 9 0 9 2
21 3 15 10 9 13 11 11 1 0 2 11 1 9 10 9 12 2 12 1 11 2
28 9 0 9 0 11 11 13 1 11 1 11 12 2 12 7 1 0 9 0 2 15 13 11 2 13 11 11 2
6 1 11 13 14 9 2
18 0 13 0 12 1 11 12 2 12 2 9 7 9 11 7 11 13 2
22 9 2 0 12 9 2 13 1 0 9 9 9 11 11 7 13 10 0 1 0 9 2
26 3 1 12 2 13 1 9 9 9 11 11 11 7 13 15 15 1 10 0 9 1 11 1 0 9 2
18 10 9 13 1 11 12 2 12 7 11 13 7 3 1 9 0 9 2
18 9 15 13 12 9 1 0 9 11 11 2 15 13 10 0 9 9 2
21 1 9 0 9 13 9 1 11 2 3 0 9 0 9 0 11 13 12 2 12 2
30 12 1 9 9 0 13 11 11 2 15 15 3 1 0 9 13 2 7 1 12 9 13 2 12 9 13 7 11 11 2
8 1 9 9 0 11 12 9 3
2 11 2
28 9 9 9 1 9 12 9 1 0 9 12 9 13 3 0 9 1 11 12 11 11 2 0 0 9 9 11 2
8 15 13 9 0 0 9 9 2
29 11 11 4 13 0 1 9 0 9 9 7 9 2 15 15 13 13 1 9 12 2 1 9 10 9 1 9 11 2
24 1 9 9 9 13 9 11 0 9 1 9 12 12 9 7 9 13 3 16 12 12 9 11 2
14 1 0 9 15 9 13 1 1 0 9 0 0 9 2
20 0 9 1 11 2 11 13 11 11 2 15 15 1 9 12 1 9 11 13 2
31 9 3 13 10 9 2 16 11 3 13 1 9 9 9 1 0 9 7 13 9 1 0 2 7 3 0 2 9 0 9 2
28 15 15 3 13 3 1 12 12 9 2 0 12 12 15 11 13 1 0 9 2 13 15 7 1 0 9 11 2
18 0 9 11 7 3 10 9 13 7 13 2 16 15 13 3 0 9 2
16 11 4 3 3 13 1 9 11 2 10 0 9 13 3 11 2
10 11 13 1 15 3 9 11 15 0 2
20 2 1 10 9 4 11 1 0 9 10 9 13 1 9 2 2 13 11 3 2
11 3 15 7 13 2 16 15 1 9 13 2
8 2 9 2 13 1 9 9 9
10 11 11 15 13 1 0 9 1 9 11
2 11 2
17 3 9 0 9 13 2 16 13 11 11 11 0 9 1 0 9 2
29 2 9 2 3 13 0 9 1 0 1 9 11 11 2 3 0 9 1 11 7 0 9 9 13 9 1 0 11 2
19 2 16 13 12 9 2 13 1 12 9 0 2 2 13 9 9 11 11 2
21 0 15 3 13 1 0 9 1 11 2 3 3 13 3 12 2 9 1 11 11 2
21 3 15 1 0 9 9 13 1 3 12 9 0 11 7 13 15 3 0 0 9 2
35 2 7 10 0 9 13 1 11 7 3 1 9 13 9 15 13 2 2 13 0 9 0 9 11 11 2 9 0 9 7 9 9 11 11 2
30 0 9 15 9 1 0 9 13 1 0 9 1 11 2 1 12 9 2 2 7 14 1 9 2 16 4 13 9 9 2
18 11 13 1 12 0 9 14 12 9 2 15 13 3 1 15 0 9 2
16 7 15 3 13 1 9 10 9 11 2 15 3 13 1 11 2
11 1 9 15 15 13 2 3 9 1 11 2
20 1 0 0 9 2 11 2 11 2 11 2 11 2 15 13 14 1 3 0 2
32 16 13 9 2 16 1 0 12 9 13 9 9 11 2 15 15 13 9 9 9 7 13 15 1 9 10 9 1 11 2 11 2
12 2 9 1 15 3 13 2 2 13 9 11 2
25 0 9 11 2 12 2 9 2 12 9 2 12 9 2 12 9 2 9 12 2 12 2 12 9 2
23 13 2 11 2 11 11 2 2 11 2 11 2 2 11 2 11 2 2 11 2 11 2 2
46 13 2 11 2 11 2 2 11 2 11 2 2 11 2 11 2 12 9 1 11 2 2 11 2 9 1 11 11 2 2 11 2 9 1 11 2 2 11 2 13 9 1 11 11 2 2
40 9 11 11 2 15 13 0 9 1 9 9 11 1 11 0 1 9 9 11 1 10 0 9 11 2 13 1 9 9 0 0 9 9 0 0 9 2 11 2 2
16 9 10 9 13 1 9 13 1 0 9 0 9 1 9 9 2
4 11 16 0 9
11 9 11 11 2 1 9 7 9 13 0 9
3 0 11 2
20 1 0 9 2 15 4 13 7 10 0 9 2 13 0 9 2 9 0 9 2
18 11 15 1 0 0 2 0 0 9 13 9 0 0 9 9 11 11 2
28 9 0 0 9 13 13 2 16 7 3 0 9 2 1 15 13 9 10 9 2 13 1 9 1 9 0 9 2
23 2 9 13 2 9 15 7 0 9 13 1 10 9 7 15 13 13 13 15 2 2 13 2
16 0 9 13 2 15 3 0 9 13 2 15 3 15 15 13 2
14 3 15 7 13 9 2 15 1 10 9 13 0 9 2
28 2 13 15 3 2 3 0 1 15 13 1 9 3 2 16 4 13 13 2 13 7 13 2 2 13 9 11 2
17 2 13 15 1 15 7 3 2 13 15 0 9 7 0 9 2 2
20 2 0 0 9 13 0 9 2 15 9 13 9 9 2 2 13 9 11 11 2
13 13 7 2 16 9 1 9 7 9 13 3 0 2
11 11 15 15 7 1 9 13 7 13 9 2
12 2 13 0 2 2 13 0 9 9 11 11 2
23 2 1 9 1 9 13 7 9 2 3 15 3 13 1 9 7 3 7 1 9 9 2 2
19 1 0 9 15 1 9 0 9 11 1 15 13 2 13 7 1 9 9 2
23 3 15 15 13 1 9 0 9 2 1 15 11 13 16 3 0 9 0 1 0 0 9 2
16 2 13 15 9 2 15 3 13 10 9 2 2 13 9 11 2
12 12 0 9 13 3 7 1 0 9 0 9 2
4 9 1 9 12
3 9 11 13
2 11 2
22 1 9 9 10 0 9 2 15 13 1 0 9 0 9 2 13 11 11 0 0 9 2
13 0 9 13 9 2 15 15 13 1 3 0 9 2
27 0 9 2 0 0 9 9 2 3 13 9 0 9 2 15 13 13 0 9 2 15 13 0 9 9 9 2
10 2 13 15 2 2 13 3 11 11 2
15 3 9 15 13 3 0 9 1 9 1 0 2 0 9 2
32 3 0 13 0 9 2 7 3 15 1 11 13 1 0 9 9 2 2 1 11 3 13 15 2 10 0 9 15 3 13 2 2
25 1 9 10 0 9 0 9 13 2 2 15 13 0 9 10 0 9 2 3 0 9 13 1 9 2
6 10 9 13 3 0 2
7 15 13 1 0 9 2 2
9 0 9 13 3 9 1 9 9 11
2 11 2
41 2 11 13 9 0 9 2 11 2 2 13 1 9 7 13 1 9 1 0 9 2 2 13 11 11 2 9 0 9 0 1 9 0 9 12 0 11 11 11 11 2
21 11 3 13 1 9 11 2 3 9 9 9 13 2 15 3 15 11 1 11 13 2
19 11 3 13 2 16 15 13 2 16 13 2 16 11 13 9 0 9 9 2
14 1 9 1 0 9 1 11 13 11 0 13 0 9 2
25 3 1 9 11 11 9 1 10 1 9 12 3 0 0 9 0 9 13 1 9 12 1 9 9 2
9 10 9 13 9 7 9 9 9 2
21 11 13 1 9 9 9 9 11 2 15 1 9 13 9 11 1 11 1 0 9 2
14 1 9 7 0 9 13 2 7 14 13 1 9 0 2
25 0 0 9 11 9 2 11 11 11 13 2 2 13 9 1 15 2 16 13 1 9 10 9 9 2
19 15 2 15 13 3 9 2 13 0 9 9 2 3 9 3 3 13 2 2
5 9 13 9 1 11
2 11 2
11 1 0 9 15 13 0 0 9 11 11 2
25 9 13 2 16 12 1 0 9 1 9 1 9 11 2 11 0 9 1 11 13 9 3 1 11 2
30 11 11 2 12 1 12 9 2 15 0 9 1 9 13 1 9 2 13 2 16 9 1 15 7 10 9 13 1 11 2
24 2 3 4 15 13 1 9 1 11 2 7 13 4 13 2 16 13 1 9 2 2 13 9 2
7 1 9 15 13 11 1 11
15 1 9 15 13 13 9 0 11 2 11 7 9 0 9 11
8 9 15 13 1 10 9 16 9
2 11 2
23 0 0 9 1 9 13 3 1 9 12 9 2 15 13 1 12 9 3 16 1 9 3 2
6 13 15 0 0 9 2
30 3 15 13 9 1 9 2 12 9 2 2 1 15 13 9 2 12 9 2 7 3 9 1 0 11 2 12 9 2 2
26 9 1 0 9 13 1 9 1 15 9 3 2 12 9 2 16 10 9 1 0 9 2 12 9 2 2
19 3 0 0 0 9 1 9 13 3 1 9 12 9 7 1 9 12 9 2
17 1 0 9 13 1 0 9 1 12 9 7 1 0 1 12 9 2
21 16 4 13 1 9 9 2 9 9 1 9 13 9 2 9 7 9 2 0 9 2
24 1 0 9 15 1 9 12 13 9 1 9 1 0 9 1 12 9 7 1 9 1 12 9 2
11 1 0 0 9 3 9 13 1 12 9 2
20 15 7 13 2 16 0 9 13 1 9 9 9 7 9 9 13 9 10 9 2
30 0 0 9 1 0 9 7 9 15 1 9 0 0 9 3 13 1 12 9 2 16 1 9 1 12 7 3 9 13 2
10 1 9 13 0 9 12 7 12 9 2
4 11 1 11 13
3 0 11 2
9 0 9 13 9 9 11 11 11 2
20 0 9 13 1 11 12 2 12 2 1 9 3 3 13 9 11 12 2 12 2
24 13 15 0 9 2 15 3 10 9 13 2 3 13 12 2 12 1 12 2 9 12 1 11 2
18 12 9 13 1 10 9 11 11 2 11 2 1 12 3 13 11 11 2
21 3 0 15 13 1 10 9 0 9 2 12 2 9 12 13 1 11 12 2 12 2
4 11 13 0 9
16 9 9 13 12 9 16 9 2 1 0 9 13 3 13 15 15
24 0 9 1 9 1 9 11 2 0 9 0 9 9 2 13 3 1 9 11 1 9 11 11 2
26 9 1 0 0 9 11 11 2 12 2 9 11 2 7 11 11 2 12 2 2 15 13 1 0 9 2
17 2 13 2 1 10 9 15 13 9 2 15 15 13 13 1 3 2
43 3 15 13 13 9 2 16 15 9 4 13 2 7 16 15 4 13 2 1 9 0 9 4 0 13 3 2 2 13 10 9 1 9 0 11 2 15 1 9 13 11 11 2
28 0 9 1 0 9 13 9 1 0 9 1 12 2 1 12 2 9 2 3 13 9 0 2 0 9 11 11 2
21 0 9 2 1 15 15 0 9 13 13 1 0 9 1 0 9 2 13 12 9 2
26 2 13 13 0 9 13 15 3 1 0 9 7 9 13 15 1 15 0 2 7 16 15 13 14 3 2
15 7 3 1 11 13 11 7 7 9 11 13 1 9 0 2
12 0 13 7 11 1 11 7 11 1 11 2 2
36 1 11 7 11 13 1 0 9 1 9 11 2 11 7 11 2 1 10 9 15 11 11 13 14 1 10 0 9 2 9 9 13 12 2 9 2
21 2 1 15 4 13 7 13 15 1 11 2 0 0 9 13 0 11 7 11 2 2
24 9 13 1 0 9 1 9 11 2 3 14 3 1 11 2 15 1 9 13 0 9 16 11 2
26 16 9 2 16 13 0 9 11 11 2 13 9 2 7 4 15 13 13 1 15 2 13 11 11 13 2
22 2 13 2 16 13 0 9 2 15 4 13 14 9 7 9 2 7 13 3 7 3 2
31 11 11 4 3 13 0 2 13 4 15 1 10 9 2 15 15 3 13 1 9 9 2 3 15 9 13 3 1 15 2 2
31 0 0 2 9 3 1 0 9 13 1 9 9 0 9 2 12 2 12 2 2 1 15 11 13 9 2 12 2 12 2 2
21 1 0 9 13 12 7 2 1 9 13 9 12 2 12 2 1 9 12 2 12 2
37 10 0 9 13 9 11 11 2 11 11 7 11 11 2 1 10 0 9 7 11 11 15 13 13 2 2 13 15 13 0 2 13 13 15 15 2 2
7 11 4 15 1 9 11 13
2 11 2
9 2 11 11 4 13 13 10 9 2
3 3 14 2
40 13 4 15 0 9 2 2 13 9 0 0 9 11 11 1 9 9 11 2 16 4 13 1 15 2 16 4 15 11 13 1 9 9 11 1 9 1 9 12 2
26 2 9 11 13 10 9 2 13 15 14 0 9 2 7 13 15 7 16 9 7 9 2 2 13 11 2
8 9 1 9 11 1 9 1 9
13 11 11 7 11 11 13 10 9 1 0 9 0 9
18 0 9 0 0 9 2 11 2 13 12 2 9 12 9 0 0 9 2
12 0 9 1 0 9 13 9 2 3 12 9 2
17 12 1 15 4 15 13 2 1 15 13 1 0 0 9 1 11 2
23 9 11 11 11 7 0 9 11 11 15 13 1 15 2 16 15 3 3 13 9 1 9 2
23 12 4 13 1 9 0 9 16 9 0 9 2 12 13 13 1 0 9 9 13 10 9 2
31 2 3 13 13 2 15 1 9 13 2 13 16 9 7 3 3 3 13 2 15 9 1 0 9 13 2 2 13 11 11 2
10 2 3 13 9 2 15 15 4 13 2
13 13 1 0 9 13 1 10 9 2 13 15 0 2
30 1 10 9 13 13 0 9 2 2 13 11 11 2 15 1 9 2 16 13 15 9 2 13 2 2 3 3 14 2 2
30 1 9 10 2 9 2 1 0 9 13 11 7 11 3 1 9 1 9 2 2 0 9 13 7 1 0 9 0 9 2
16 13 0 13 9 9 0 9 1 9 1 9 9 1 0 9 2
23 13 4 15 13 9 1 9 2 16 15 13 9 2 15 13 0 0 9 7 13 7 9 2
16 7 11 13 9 0 9 7 0 9 13 0 9 1 9 11 2
10 3 15 13 13 11 2 11 7 11 2
9 9 1 9 13 7 9 1 9 2
13 13 0 13 9 2 16 13 14 1 0 9 2 2
22 11 13 0 9 9 1 9 2 0 13 0 11 2 2 15 9 4 13 13 1 9 2
8 0 13 7 9 0 0 9 2
23 13 0 13 9 1 9 9 2 16 4 0 9 3 13 2 16 13 1 0 9 9 2 2
38 9 11 11 11 15 13 9 0 9 2 2 1 9 15 4 13 0 9 2 1 9 0 9 7 9 9 0 9 15 4 9 13 9 0 9 9 2 2
47 9 1 0 9 9 13 3 0 2 0 9 11 4 3 0 9 13 7 16 9 9 2 3 9 0 9 2 2 0 9 13 1 9 7 1 11 13 3 13 2 10 9 13 4 9 13 2
24 1 0 0 9 13 12 9 2 11 2 13 9 1 9 2 0 2 11 2 13 0 1 9 2
19 0 9 9 13 1 9 9 2 9 2 9 0 9 7 9 9 7 9 2
1 3
16 11 15 1 9 9 9 13 11 7 11 1 0 9 11 11 2
14 1 9 12 9 13 11 11 2 9 11 1 0 9 2
18 1 9 12 7 12 13 1 11 11 0 9 1 9 1 11 7 11 2
9 9 15 13 12 2 9 1 11 2
36 9 9 1 12 9 7 9 12 9 13 0 9 0 9 0 9 9 11 1 0 9 9 7 9 9 1 9 12 2 9 1 9 1 0 11 2
17 9 2 1 15 15 9 13 2 13 9 13 3 12 9 1 11 2
8 9 3 13 0 9 11 9 2
25 1 0 9 2 1 15 13 9 0 0 9 11 11 1 11 1 11 2 15 3 14 12 9 13 2
13 1 9 11 2 11 13 11 11 9 1 12 9 2
2 0 9
21 3 12 9 13 0 0 9 9 1 10 2 16 4 15 1 9 10 9 13 13 2
5 13 3 0 9 2
19 0 9 1 11 7 11 11 2 12 2 12 2 13 7 9 11 11 11 2
26 2 13 4 15 1 0 9 11 13 2 16 4 15 13 1 9 11 1 11 2 2 13 11 10 9 2
15 3 15 13 2 13 7 1 11 9 11 1 11 11 11 2
23 2 11 1 11 1 15 13 1 9 7 3 15 13 13 2 16 15 15 13 1 9 2 2
21 0 9 13 0 11 1 0 9 3 2 2 13 2 3 4 15 1 15 13 2 2
4 0 9 0 9
2 11 2
19 11 1 0 12 2 9 0 9 13 11 7 3 13 10 9 1 9 14 2
15 11 13 1 0 12 9 0 0 9 1 0 9 1 11 2
27 9 2 15 13 7 1 11 3 9 2 15 3 13 1 15 2 16 4 1 9 13 9 1 11 7 11 2
16 15 12 9 1 0 2 0 0 9 1 9 14 13 12 9 2
8 11 2 0 2 11 12 2 12
14 0 13 3 2 3 1 12 2 9 1 9 11 13 2
12 0 1 0 11 7 3 13 9 0 9 11 2
12 1 12 2 9 9 9 13 7 15 13 11 2
11 9 15 13 1 12 2 9 1 9 11 2
7 9 0 12 13 3 9 2
18 1 12 2 9 13 1 9 9 11 11 2 1 12 9 3 13 11 2
20 3 11 13 9 1 0 12 2 7 9 3 13 0 9 11 1 12 2 9 2
8 9 2 11 2 11 2 11 2
6 11 2 11 12 2 12
18 11 1 11 7 11 13 3 0 2 7 11 1 12 2 9 13 9 2
18 1 0 9 0 9 11 13 3 13 2 7 1 9 11 13 3 0 2
19 0 9 13 1 12 2 9 2 3 11 15 13 0 9 3 13 9 9 2
9 1 9 15 13 0 0 9 11 2
23 12 10 0 9 3 11 13 2 7 1 10 0 9 1 9 12 9 1 9 9 13 0 2
8 9 2 11 2 11 2 11 2
6 11 2 11 12 2 12
23 0 15 1 9 9 13 13 0 9 0 7 12 9 15 14 13 2 7 13 15 9 11 2
21 15 3 13 1 12 2 9 2 3 13 9 7 0 9 11 1 9 13 0 9 2
16 1 12 2 12 13 0 1 12 2 9 2 11 9 13 11 2
14 10 15 9 1 12 9 3 13 11 9 0 12 9 2
8 9 2 11 2 11 2 11 2
6 11 2 11 12 2 12
17 0 11 13 1 12 2 9 9 1 11 7 13 15 12 2 12 2
18 1 12 9 3 7 1 9 11 13 13 1 15 9 11 7 11 13 2
21 1 12 2 9 11 13 9 2 11 13 1 0 9 0 7 13 9 1 9 0 2
13 3 9 11 1 11 11 13 7 11 15 13 9 2
20 16 1 0 0 9 11 13 11 0 9 2 13 3 0 0 13 1 12 9 2
8 9 2 11 2 11 2 11 2
6 11 2 11 12 2 12
18 0 9 2 3 15 13 14 1 9 9 2 3 7 13 12 9 13 2
9 14 1 9 9 15 13 0 9 2
23 0 15 13 1 12 2 9 2 16 13 1 12 9 12 9 2 7 15 13 1 9 9 2
27 9 0 12 13 1 12 2 9 10 0 9 11 2 15 15 3 13 0 0 9 3 12 9 1 9 9 2
8 9 2 11 2 11 2 11 2
18 1 12 2 9 2 12 9 1 9 0 11 2 13 0 0 9 11 2
18 11 15 3 15 13 1 3 0 9 2 7 3 0 1 9 3 13 2
21 9 13 1 9 0 12 9 11 7 1 0 12 9 15 13 9 3 1 0 9 2
12 9 9 7 3 1 9 0 9 1 9 13 2
34 1 9 11 13 11 0 9 11 7 9 1 11 3 3 16 9 1 9 13 0 0 9 1 0 9 2 3 15 3 13 1 9 14 2
9 1 0 9 13 14 1 0 9 2
40 3 3 11 13 0 9 2 7 3 1 0 12 9 0 0 9 3 13 11 2 15 1 0 12 13 0 11 2 11 2 3 1 0 9 12 9 1 9 2 2
21 9 2 7 16 1 15 13 0 12 9 9 0 9 12 1 12 2 9 3 13 2
19 9 0 9 11 11 2 3 2 7 9 9 11 11 7 11 9 2 3 2
2 11 13
2 11 2
27 0 9 11 0 11 11 4 3 0 9 13 1 9 1 9 1 9 11 0 1 9 11 11 12 2 9 2
8 0 9 3 13 1 0 9 2
15 11 4 13 1 9 7 12 2 9 15 13 13 1 9 2
11 13 4 13 3 0 9 7 9 12 9 2
4 11 1 11 13
2 11 2
30 3 12 12 9 15 13 0 9 1 9 1 0 0 0 9 2 12 2 12 9 2 2 0 11 11 1 0 11 11 2
27 2 13 2 16 13 0 0 9 7 1 9 13 3 0 9 1 12 12 9 2 2 13 0 9 11 11 2
13 1 9 13 2 16 3 11 1 11 3 3 13 2
43 1 9 9 1 0 9 1 3 12 9 13 12 2 9 12 1 0 0 9 1 11 2 3 2 12 9 2 7 3 12 1 0 9 9 13 2 16 4 13 3 12 9 2
9 10 0 9 13 3 0 9 11 2
3 1 0 9
19 11 11 4 13 1 9 9 0 9 11 1 0 9 7 0 9 1 9 2
16 1 9 12 2 3 15 11 13 9 2 13 11 3 1 9 2
7 0 9 15 13 11 11 2
18 11 13 1 12 7 12 9 9 11 11 2 1 10 9 13 12 9 2
17 0 9 13 9 2 16 11 13 0 1 9 0 9 1 9 9 2
3 0 9 13
1 9
25 11 11 2 11 11 2 11 11 2 1 10 0 9 9 9 1 9 13 1 0 9 0 0 9 2
34 13 2 14 1 3 0 9 9 0 0 9 2 13 2 16 13 3 13 1 9 0 9 1 9 9 7 13 0 0 9 2 0 2 2
35 9 1 0 9 1 9 15 13 13 3 1 9 0 2 0 9 2 9 1 11 11 2 1 0 9 9 11 11 7 1 0 9 11 11 2
14 9 16 9 1 9 7 0 9 9 13 9 7 9 2
41 9 1 0 7 0 9 9 2 9 7 0 9 0 9 3 13 13 1 0 9 1 9 11 11 2 0 9 11 11 7 1 9 9 2 9 2 9 9 11 11 2
12 1 9 1 0 9 15 13 0 9 11 11 2
29 1 0 9 9 15 13 10 9 2 9 9 1 9 2 0 9 2 13 3 1 9 7 3 16 12 9 7 9 2
11 9 3 13 3 13 7 13 1 0 9 2
41 0 9 2 1 15 4 9 13 2 7 13 7 1 9 0 2 1 0 9 2 2 7 1 9 0 9 2 0 9 2 11 7 11 2 7 9 2 3 11 2 2
19 9 13 16 3 0 9 0 9 1 9 2 15 0 9 13 1 12 9 2
26 0 9 15 13 9 1 9 2 0 9 3 3 13 0 9 2 0 9 9 2 9 9 2 9 3 2
7 9 13 3 13 1 9 2
24 9 0 0 9 13 7 9 1 9 2 1 11 2 11 11 2 0 0 9 2 7 1 9 2
15 1 15 15 1 15 13 13 9 9 7 0 9 0 9 2
8 11 13 0 9 2 15 13 15
22 0 9 11 11 2 12 2 15 3 3 2 1 12 9 2 13 1 0 0 9 11 2
28 9 10 2 0 2 9 2 0 9 11 2 2 15 11 13 1 9 0 0 9 2 10 9 7 9 3 13 2
29 1 12 9 0 0 7 0 9 13 1 15 0 14 9 9 1 9 2 13 9 12 1 9 11 11 1 11 2 2
31 0 0 9 7 9 10 9 2 15 1 10 9 2 0 9 7 9 4 13 3 2 13 13 0 0 9 7 9 0 11 2
31 11 15 13 13 1 11 2 13 9 11 2 9 12 2 12 13 1 11 2 13 1 11 7 1 9 0 9 13 1 11 2
11 9 1 9 1 9 0 9 11 3 13 2
15 3 0 15 13 3 0 9 9 2 15 0 9 3 13 2
11 7 4 0 0 9 13 13 7 10 9 2
28 1 10 9 2 1 10 9 0 2 13 3 11 13 16 9 9 2 15 14 13 15 2 9 2 11 7 11 2
5 0 9 1 0 9
24 3 12 9 13 9 9 0 9 0 9 2 11 2 12 2 15 13 1 9 1 0 9 11 2
11 1 9 13 0 9 11 7 0 0 11 2
28 1 0 1 9 2 13 15 0 9 14 1 12 2 9 2 13 12 1 12 12 9 2 15 13 0 0 9 2
19 1 11 13 9 1 0 11 2 11 2 11 2 0 9 7 1 0 9 2
8 9 13 13 1 12 2 9 2
13 3 3 15 1 11 13 7 0 9 0 9 11 2
15 9 13 12 2 2 12 2 7 12 2 9 1 9 11 2
11 0 9 15 13 1 0 9 12 2 9 2
6 0 0 11 13 1 11
14 0 0 0 9 0 11 15 3 13 7 1 0 9 2
48 3 1 0 0 9 2 15 15 13 11 2 7 1 0 0 2 0 9 0 11 2 3 13 7 0 9 0 11 11 11 2 15 13 1 9 9 12 2 12 11 3 1 0 0 9 1 9 2
19 9 15 3 13 1 15 13 2 3 0 9 12 0 9 3 13 0 9 2
38 0 11 2 1 9 11 11 2 11 11 7 11 11 2 13 3 1 9 12 1 0 11 2 7 1 0 0 9 13 3 3 2 13 3 16 9 0 2
15 13 7 3 7 13 9 2 7 1 15 7 10 0 9 2
27 1 9 9 7 12 0 2 9 13 1 9 12 3 0 9 0 14 0 2 0 1 0 9 0 9 2 2
8 15 13 3 0 0 0 9 2
30 0 9 1 9 11 2 9 9 1 9 12 15 3 3 13 2 0 9 4 9 3 13 7 15 3 2 9 3 13 2
26 3 1 9 9 15 0 11 13 14 1 9 12 1 9 13 15 11 2 0 3 1 0 9 0 0 2
36 0 9 1 9 0 9 7 13 0 9 2 3 15 3 13 9 0 9 7 0 9 1 9 15 0 9 7 1 10 9 3 0 9 0 9 2
20 0 9 9 2 13 15 9 0 0 9 1 0 9 2 15 13 9 1 11 2
16 3 4 1 9 10 0 9 13 1 10 9 1 0 0 9 2
23 13 2 14 1 9 2 10 9 15 0 9 13 2 10 9 1 0 9 13 3 16 0 2
14 9 13 14 1 0 11 2 7 13 7 1 9 0 2
18 7 3 13 1 0 9 2 13 9 0 11 3 7 3 1 0 9 2
23 1 9 2 15 11 13 9 12 2 12 11 2 13 1 0 9 1 9 3 3 12 9 2
7 0 9 11 13 1 0 9
17 9 1 0 9 0 9 13 1 9 0 0 9 11 2 11 11 2
25 1 11 15 13 9 1 9 0 9 11 11 2 0 9 11 7 9 1 11 7 9 9 12 2 2
27 11 2 12 2 13 3 1 12 9 0 9 1 0 0 9 1 11 7 13 0 1 0 7 0 0 9 2
25 0 9 13 1 0 9 1 0 0 11 1 9 12 2 13 1 9 0 9 2 1 11 7 11 2
25 1 10 9 1 9 0 9 1 11 13 12 9 16 9 0 0 9 7 13 0 9 0 0 9 2
13 11 13 3 0 9 7 0 9 1 10 0 9 2
13 3 13 0 9 0 0 9 7 9 0 0 9 2
6 1 11 13 0 15 13
11 11 13 9 2 7 1 9 3 14 3 13
2 11 2
14 1 12 9 0 15 14 12 13 3 13 1 9 11 2
10 13 15 3 13 0 3 9 0 9 2
25 1 9 11 13 1 0 11 0 9 3 1 11 7 11 2 16 3 16 11 13 9 1 0 9 2
31 9 9 11 2 9 11 2 11 11 2 1 15 15 11 13 3 13 2 13 9 1 0 9 1 0 0 9 1 3 0 2
25 0 0 9 7 3 3 1 9 13 2 16 4 15 1 9 9 13 13 7 0 9 16 0 11 2
44 9 3 13 9 0 9 9 2 15 15 14 13 13 15 9 1 9 1 9 9 12 2 7 3 13 2 16 10 9 2 15 1 0 9 4 13 0 9 2 13 12 12 9 2
21 9 9 7 3 11 1 12 9 2 3 15 1 9 13 13 7 0 9 2 13 2
10 3 1 9 15 0 13 1 9 11 2
19 15 13 1 9 9 2 9 11 7 9 9 9 2 15 15 13 1 9 2
11 1 11 9 11 13 9 0 9 9 9 2
27 16 9 0 9 9 11 3 13 2 0 9 13 9 9 2 16 4 3 13 9 9 0 9 1 9 11 2
26 1 10 9 15 13 3 2 16 11 13 2 16 1 9 11 2 9 11 2 13 3 9 0 0 9 2
14 2 13 7 2 16 4 13 0 9 2 2 13 11 2
12 9 0 9 11 11 2 11 9 1 11 13 2
13 13 7 2 16 0 9 4 13 1 9 0 9 2
26 1 9 11 2 3 15 1 9 11 13 13 0 9 2 13 2 16 11 1 9 3 13 0 0 9 2
5 15 2 3 2 3
36 9 11 0 0 9 11 11 2 15 1 11 13 3 12 9 1 3 0 0 9 2 13 3 1 12 1 0 0 9 1 11 2 0 12 2 2
21 11 11 1 11 13 9 9 2 15 3 1 12 9 13 9 1 0 9 1 11 2
14 9 11 11 13 3 1 12 9 1 0 11 9 9 2
6 1 11 3 1 0 9
18 1 0 0 9 4 1 0 9 2 0 9 2 13 12 0 0 9 2
19 0 9 13 1 12 2 1 12 2 9 2 9 9 13 13 3 11 11 2
32 9 15 13 12 1 0 9 9 12 2 9 9 11 2 1 10 9 13 3 0 9 12 9 9 7 9 0 11 1 0 9 2
19 1 9 15 13 7 1 9 0 9 3 0 9 7 1 9 11 9 11 2
2 0 9
1 9
14 9 2 0 9 0 0 9 13 12 9 9 11 11 2
37 13 15 9 1 9 2 15 15 1 9 13 14 10 9 7 9 2 7 7 0 9 0 0 9 2 11 11 2 11 11 2 11 11 7 11 11 2
41 9 0 9 11 13 1 11 11 7 1 9 0 9 2 11 2 11 11 2 11 2 11 11 11 2 11 2 11 11 2 11 2 11 11 2 11 2 11 11 2 2
16 7 3 10 9 13 15 1 15 3 0 2 15 13 7 13 2
27 9 13 3 1 0 9 2 3 0 9 11 11 2 1 3 0 7 0 9 9 2 1 9 7 9 9 2
15 15 15 13 3 9 11 2 3 0 2 7 3 3 0 2
10 7 3 13 15 9 9 0 0 9 2
41 1 0 9 15 3 3 13 0 11 11 11 2 3 3 0 2 3 3 0 11 11 2 0 9 1 10 9 13 3 1 15 2 7 9 0 9 2 0 11 11 2
25 9 11 11 13 9 0 9 9 2 3 3 3 2 16 13 13 1 0 2 14 0 9 11 11 2
47 13 2 14 13 9 1 9 9 9 2 7 0 0 9 15 13 2 2 13 0 2 16 0 9 11 11 15 1 1 12 0 9 7 12 9 2 2 2 13 1 0 12 9 3 1 12 2
31 9 0 9 1 11 13 9 9 9 9 2 15 4 3 13 1 0 9 0 0 11 2 15 3 13 10 9 0 7 0 2
25 9 0 9 11 11 13 10 9 1 9 9 9 1 3 0 9 2 15 3 13 9 7 3 9 2
11 1 9 9 13 0 9 1 9 0 9 2
5 0 9 7 13 2
19 0 13 9 9 2 16 15 4 13 9 11 11 1 0 9 1 9 12 2
17 9 9 13 1 9 3 0 2 9 2 12 9 1 0 0 9 2
12 0 13 7 9 11 11 1 0 0 0 11 2
18 13 10 10 0 9 7 1 15 13 0 9 2 7 9 13 9 2 2
17 3 2 3 10 9 13 9 1 9 9 2 13 11 9 9 9 2
24 0 9 13 11 11 7 1 0 9 13 15 1 9 2 15 13 3 1 11 9 0 0 9 2
27 0 9 7 1 9 10 0 9 13 7 9 7 3 13 3 7 3 3 0 2 7 3 0 9 11 11 2
20 1 3 0 9 11 11 2 9 2 7 1 0 9 11 11 7 13 0 9 2
11 7 7 1 9 13 3 14 11 11 11 2
11 10 0 9 13 7 0 9 9 0 9 2
2 11 11
15 9 0 0 9 2 0 9 11 2 11 11 2 11 11 2
9 13 1 0 0 9 12 2 9 2
5 9 0 0 9 2
11 0 9 11 2 11 11 2 9 9 9 2
9 13 1 0 0 9 12 2 9 2
4 0 9 9 9
10 0 9 11 11 13 10 9 1 9 11
28 1 0 9 0 9 1 11 13 13 0 9 11 11 2 12 2 12 2 2 12 1 0 9 0 9 0 9 2
20 3 15 13 1 11 7 13 0 9 10 0 9 2 9 7 0 9 9 9 2
19 3 1 10 9 1 9 0 9 13 0 9 13 0 9 3 1 10 9 2
24 3 3 7 13 9 13 0 9 2 9 2 9 7 9 2 15 13 9 10 0 7 0 9 2
26 11 11 3 13 2 13 1 11 2 11 2 11 7 11 2 7 3 13 0 9 2 0 10 0 9 2
14 13 15 1 0 1 0 9 7 0 9 13 10 9 2
6 0 0 9 13 9 2
23 0 9 9 7 9 2 9 1 0 9 9 7 0 9 7 9 9 13 10 9 11 11 2
22 9 1 9 0 9 1 10 9 7 3 9 0 9 0 9 15 13 10 9 11 11 2
23 11 11 15 13 3 1 9 2 9 7 9 2 13 0 9 2 15 13 1 0 9 9 2
30 1 0 9 15 3 13 10 0 9 7 9 2 0 3 0 9 2 9 0 1 9 7 0 9 0 9 7 0 9 2
12 0 9 15 1 0 9 1 0 9 3 13 2
24 9 0 9 15 13 1 0 9 2 0 7 9 1 0 9 7 0 9 1 9 0 0 9 2
13 0 9 3 13 7 13 15 9 9 0 0 9 2
19 3 3 13 0 0 7 3 3 0 0 9 2 10 9 13 0 0 9 2
15 9 13 0 9 1 0 9 2 0 0 9 7 0 9 2
20 9 15 3 13 9 2 13 3 9 3 1 0 2 3 0 9 0 0 9 2
6 11 11 2 0 9 2
8 9 11 2 0 9 1 11 2
8 12 2 9 2 12 2 9 2
4 11 1 0 9
1 9
13 9 2 11 11 16 9 13 0 0 9 0 9 2
36 16 13 0 9 9 2 9 9 0 0 9 7 0 0 9 1 0 9 1 0 0 9 1 11 2 13 9 1 14 0 9 3 0 9 9 2
16 0 9 13 12 1 10 0 0 9 2 10 9 13 0 9 2
20 0 0 9 13 3 7 3 2 1 0 9 7 1 9 3 0 9 0 9 2
13 9 13 1 9 2 15 16 4 13 3 1 9 2
28 3 3 16 1 0 9 9 2 9 15 13 1 0 9 2 15 7 14 0 9 3 13 2 14 14 1 9 2
14 3 0 9 7 0 0 9 13 1 0 9 3 3 2
16 1 12 9 3 11 13 0 9 0 1 10 9 1 11 11 2
14 1 9 12 13 11 15 1 10 9 1 0 0 9 2
7 11 15 15 13 1 9 2
5 0 2 9 11 2
3 1 0 9
33 16 9 0 9 2 11 2 13 13 9 9 1 11 2 9 11 11 4 13 3 13 2 2 13 4 15 13 11 2 11 13 2 2
32 13 15 3 9 9 1 9 1 2 9 2 2 15 13 9 9 12 9 11 1 3 3 0 9 11 11 1 0 9 1 11 2
25 11 2 14 1 0 9 2 13 7 1 9 0 9 0 9 1 9 2 9 7 0 9 11 11 2
23 9 2 0 9 2 1 12 0 9 7 13 1 0 9 2 15 13 0 9 2 13 9 2
23 10 9 13 9 2 16 9 11 1 0 0 9 9 9 11 13 13 9 7 9 0 9 2
25 0 9 11 13 2 16 0 9 12 9 11 13 1 9 7 0 9 0 9 1 9 9 11 11 2
33 16 0 2 3 1 9 11 13 1 9 9 11 11 7 9 9 11 11 9 1 9 2 15 0 9 13 1 10 9 9 7 9 2
24 1 9 9 2 7 3 1 9 9 11 2 11 1 15 2 13 9 0 9 1 0 9 9 2
28 1 0 9 9 11 13 2 16 1 10 9 13 13 13 1 11 0 9 0 9 11 2 9 11 7 11 0 2
8 2 13 4 2 16 4 13 2
49 1 9 1 9 11 2 2 2 4 13 2 16 15 2 15 1 15 13 2 13 1 9 10 9 7 0 9 3 0 2 2 13 9 11 0 9 11 2 15 3 1 9 13 1 9 0 9 9 2
5 0 9 1 9 2
41 0 9 1 11 3 13 1 15 2 16 0 9 1 0 9 11 11 11 2 12 2 4 13 7 13 0 9 2 1 15 4 4 13 1 12 9 9 1 0 12 2
32 0 9 7 0 9 11 13 13 2 16 13 10 9 1 15 2 16 4 1 9 11 0 1 9 1 9 13 16 9 10 9 2
11 13 15 15 1 9 3 9 7 0 9 2
24 9 13 9 0 9 7 13 15 3 1 9 0 9 2 1 15 13 4 9 13 1 0 9 2
32 1 0 9 4 4 1 11 13 7 0 9 0 0 9 2 11 2 11 11 2 12 2 2 15 13 1 9 9 1 12 9 2
16 9 13 1 9 0 9 7 13 1 10 9 13 9 0 9 2
14 0 9 13 11 11 2 15 10 9 13 7 11 11 2
37 1 12 0 9 11 16 9 0 9 1 0 0 9 13 9 1 9 1 0 0 9 2 16 4 15 3 13 10 9 2 15 3 13 9 0 9 2
14 1 9 12 2 12 13 3 1 0 9 9 0 9 2
13 1 10 9 13 3 1 0 9 9 12 9 9 2
16 1 0 9 13 1 9 12 0 11 7 4 13 12 0 9 2
3 9 0 9
24 16 4 15 9 0 9 13 13 9 9 0 9 1 9 2 13 4 3 3 9 1 0 9 2
9 13 4 3 1 9 1 9 9 2
7 10 9 4 3 13 9 2
44 0 9 9 9 2 15 13 9 0 9 2 13 12 9 1 0 9 2 9 0 9 2 0 9 0 9 1 10 0 0 9 7 0 9 9 9 9 7 9 0 9 11 11 2
44 2 13 15 2 16 9 1 10 9 7 10 9 15 3 13 9 2 2 13 15 1 0 9 3 2 16 9 9 13 1 9 10 9 7 15 15 3 13 1 0 9 0 9 2
61 9 1 9 9 9 7 9 1 11 1 0 9 0 9 13 1 0 9 2 3 13 9 1 0 9 0 0 9 0 1 10 9 9 2 3 3 2 9 13 1 15 2 16 4 9 13 1 0 9 0 9 3 11 0 9 1 9 7 1 9 2
21 10 9 13 0 9 2 0 9 13 13 1 0 12 9 2 0 1 0 12 9 2
33 0 9 9 13 0 0 9 3 1 9 2 16 12 0 0 9 11 2 12 7 11 13 2 16 0 9 1 9 7 9 13 4 2
24 1 9 9 13 9 9 7 9 1 9 1 9 11 1 3 0 9 7 9 13 13 0 9 2
13 9 1 9 7 9 9 3 13 9 9 1 9 2
35 3 15 9 13 13 1 10 9 9 1 11 2 13 15 1 0 9 9 9 2 15 3 13 0 9 7 13 0 9 2 16 4 15 13 2
11 0 9 15 13 9 11 2 11 7 11 2
16 16 0 9 13 0 9 2 9 13 0 9 1 9 1 11 2
11 1 9 1 9 13 1 9 9 11 11 2
11 1 9 1 0 9 15 13 1 12 9 2
27 1 0 9 2 0 9 7 0 9 15 13 11 11 2 15 11 13 1 2 11 1 11 2 0 9 9 2
20 9 1 9 9 15 9 9 13 1 0 9 7 9 1 0 9 0 9 11 2
12 9 1 9 9 13 1 9 1 9 1 9 2
13 1 0 0 9 13 1 9 9 9 1 9 9 2
20 2 13 15 1 9 10 0 9 2 2 13 3 10 9 0 9 9 11 11 2
4 9 7 0 9
3 1 0 9
21 0 0 9 1 11 1 11 13 10 0 9 2 15 7 3 13 3 13 3 0 2
14 0 9 9 3 10 0 9 13 2 7 10 9 13 2
28 9 0 9 3 13 9 0 9 1 9 11 2 7 3 0 9 9 0 1 11 2 13 3 0 9 0 11 2
22 9 9 2 16 11 13 11 3 1 0 9 0 9 2 13 13 10 9 2 13 9 2
24 9 9 11 11 1 0 9 13 2 16 2 15 2 11 2 13 10 9 2 14 15 15 2 2
27 1 0 11 15 3 3 13 13 2 16 0 9 9 1 11 13 1 11 1 9 2 7 1 0 0 9 2
11 9 13 2 16 0 9 3 13 0 9 2
26 7 3 12 1 0 9 1 0 9 13 1 9 2 16 9 0 9 3 3 13 13 7 9 10 9 2
11 9 0 0 9 3 13 3 13 16 3 2
22 9 2 16 3 3 1 10 9 13 16 0 9 2 3 0 9 13 2 13 0 11 2
1 3
24 9 0 9 11 2 11 7 10 0 9 11 2 11 1 0 9 0 11 13 3 9 0 9 2
13 9 15 13 1 0 9 9 9 0 0 0 9 2
35 12 0 9 0 0 9 13 9 1 0 9 7 0 9 2 13 3 0 9 9 11 11 1 9 1 0 9 7 0 9 0 9 0 9 2
23 9 1 9 9 13 0 0 9 1 9 7 0 9 11 2 1 15 13 1 0 9 11 2
41 0 9 3 1 2 0 2 9 7 2 1 10 9 9 2 13 0 9 2 13 0 9 11 1 11 11 1 0 11 1 9 2 15 4 3 13 1 0 9 11 2
38 3 13 13 2 3 4 13 0 0 9 2 13 1 9 9 0 0 9 2 0 0 9 7 9 0 9 0 9 1 9 9 2 9 11 11 2 11 2
29 0 9 11 2 11 1 0 9 11 13 2 16 0 9 11 2 11 13 3 1 11 1 9 1 0 9 0 9 2
5 9 0 9 13 2
13 13 14 2 16 3 4 13 1 9 9 2 12 2
18 9 0 11 11 11 13 2 16 10 9 11 13 0 9 9 0 9 2
8 1 0 13 1 10 0 9 2
16 0 9 9 0 9 3 1 12 9 3 13 0 9 1 11 2
9 9 1 9 13 3 0 0 9 2
18 0 3 13 9 0 1 9 9 1 9 1 9 7 1 9 0 9 2
5 11 13 1 0 9
10 1 0 9 13 9 11 7 0 9 11
22 16 0 9 9 13 3 9 0 9 1 9 9 9 1 9 9 0 9 11 1 11 2
10 1 9 7 0 9 1 1 11 13 2
35 9 15 1 9 1 0 9 13 13 7 0 1 3 0 0 9 2 0 9 11 11 11 2 15 1 11 3 13 9 9 9 7 0 9 2
26 3 0 0 2 9 11 2 2 1 10 9 1 11 13 12 9 0 0 0 9 2 3 13 16 9 2
12 7 3 13 7 1 3 2 0 2 9 0 2
10 12 1 0 0 9 13 9 0 9 2
30 12 9 9 2 9 0 0 0 9 2 13 1 9 12 1 0 9 11 9 2 1 10 9 0 9 13 12 0 9 2
43 9 0 9 11 11 2 9 9 10 9 11 11 7 0 0 9 11 11 4 1 9 12 1 9 13 1 15 2 16 1 9 9 13 1 11 9 1 9 12 9 0 9 2
10 15 3 13 1 9 0 9 10 9 2
16 15 12 0 1 10 0 9 2 1 9 1 10 9 2 13 2
9 13 15 2 16 15 13 15 13 2
9 3 7 13 1 9 0 0 9 2
13 0 9 13 0 9 7 1 9 9 13 3 0 2
5 0 9 9 13 2
12 13 3 14 1 9 2 0 9 13 9 9 2
41 0 9 13 3 3 2 12 1 0 9 2 15 13 0 9 9 1 0 7 9 11 2 4 1 9 13 13 0 0 9 9 11 11 2 0 1 9 0 0 9 2
9 13 4 13 2 16 4 3 13 2
13 1 3 0 9 4 10 9 1 9 9 12 13 2
18 0 9 1 0 9 9 9 3 0 9 1 0 9 9 13 2 11 2
15 11 15 1 0 9 13 3 1 10 9 0 9 13 9 2
12 1 0 0 9 9 13 9 1 0 0 9 2
5 14 1 0 9 2
26 15 4 1 9 13 0 1 11 2 0 9 11 1 0 9 2 11 11 7 9 0 0 9 11 11 2
29 10 9 13 9 3 14 1 9 11 2 0 9 11 2 7 1 11 2 9 11 7 1 9 9 12 9 0 9 2
14 0 9 1 15 1 0 9 13 2 14 2 0 9 2
32 16 3 1 11 7 11 10 9 1 11 3 13 2 0 9 9 1 11 13 2 16 3 4 13 13 13 9 2 0 9 2 2
16 0 9 4 13 1 12 0 0 9 1 9 9 7 0 9 2
14 9 13 9 11 2 11 11 13 1 9 0 0 9 2
6 11 13 14 0 9 11
2 11 2
33 1 0 9 9 11 13 4 13 9 1 9 9 0 0 9 11 11 11 2 1 15 2 16 1 10 9 13 0 9 13 11 11 2
14 13 15 1 3 0 9 11 2 15 15 13 4 13 2
20 9 9 3 9 1 0 9 3 13 2 7 7 3 1 10 0 9 3 13 2
29 1 0 9 9 13 9 9 11 11 2 16 1 10 9 4 1 10 9 13 2 3 15 13 7 9 9 11 11 2
39 1 9 11 3 13 9 9 15 13 7 1 9 2 3 3 13 9 11 7 9 9 11 2 15 9 0 9 11 13 9 13 7 13 15 0 9 10 9 2
4 0 9 4 13
2 11 2
32 0 9 7 0 9 1 0 9 1 9 11 11 13 9 0 9 0 9 2 1 15 15 3 1 0 9 13 15 9 0 9 2
13 13 15 1 9 9 2 15 3 13 0 9 11 2
30 1 0 9 4 1 9 13 0 9 11 11 2 1 15 15 13 12 5 9 2 3 1 12 9 3 16 1 0 9 2
19 13 15 3 0 9 1 11 11 11 2 15 13 12 5 2 3 16 11 2
4 11 13 9 9
2 11 2
42 0 9 9 1 9 11 2 11 2 3 13 2 16 0 9 13 9 13 0 9 1 11 7 13 1 15 0 9 2 15 4 3 13 13 1 9 0 9 1 0 9 2
52 2 13 2 16 0 9 4 13 4 3 7 3 13 7 13 4 13 1 0 7 0 9 2 2 13 9 0 9 11 11 11 11 1 11 1 9 9 9 0 0 9 1 0 0 2 0 9 1 9 0 9 2
26 0 9 9 13 2 16 0 9 9 13 12 1 9 2 1 15 4 0 9 1 0 9 1 11 13 2
28 13 2 16 0 0 9 1 9 0 9 2 3 13 1 9 9 0 2 0 9 0 9 11 7 9 11 2 2
31 2 0 9 11 13 0 9 0 9 13 1 15 2 16 13 1 0 9 2 2 13 11 11 2 1 15 13 16 9 13 2
27 1 9 2 15 4 3 4 13 1 0 9 2 11 11 13 11 2 11 2 11 2 9 0 9 7 11 2
15 9 13 9 11 11 11 2 15 1 0 9 13 3 3 2
13 1 11 3 0 9 13 0 2 0 9 1 9 2
15 12 9 15 3 13 1 9 0 9 1 9 1 0 9 2
5 1 9 0 9 9
26 9 1 9 0 11 4 1 0 9 13 1 0 9 7 1 0 9 1 15 4 13 0 0 9 9 2
15 3 3 13 11 11 1 0 0 9 9 9 10 0 9 2
13 1 10 9 13 1 3 0 9 1 9 7 9 2
10 0 9 0 9 13 3 10 0 9 2
15 0 9 1 9 13 0 9 7 9 10 9 13 3 0 2
32 13 7 0 0 9 3 13 2 16 1 9 0 1 15 2 15 13 1 9 0 14 13 2 15 13 3 3 13 2 13 11 2
11 1 11 15 1 10 9 13 9 1 9 2
17 12 1 9 13 7 9 1 0 9 7 9 2 13 3 3 2 2
5 0 9 2 12 0
10 9 11 11 13 11 1 2 0 9 2
23 1 12 12 9 13 1 12 2 9 12 1 12 2 9 12 1 0 9 11 7 10 9 2
16 10 9 3 1 11 13 0 9 11 11 2 9 1 0 9 2
28 15 11 2 11 13 2 16 1 9 9 4 13 0 9 7 16 0 9 15 13 1 9 13 3 1 12 9 2
42 1 9 2 15 9 13 2 15 13 2 16 3 0 9 1 9 3 0 9 11 13 0 13 3 1 9 9 1 11 1 0 0 9 2 3 0 9 3 13 0 9 2
28 9 13 2 16 1 11 3 13 12 9 1 9 1 12 9 2 12 9 0 12 9 2 12 9 0 12 9 2
13 13 3 12 12 9 1 9 1 12 7 12 9 2
14 1 10 9 13 12 9 0 7 14 12 9 1 9 2
15 3 13 7 4 13 1 10 9 1 9 14 12 12 9 2
15 11 15 3 13 1 9 9 9 1 0 9 11 1 11 2
11 13 2 16 9 13 9 2 0 9 2 2
35 2 9 9 13 2 16 15 1 11 13 7 13 2 2 13 11 2 15 15 1 10 9 1 11 13 1 11 7 3 15 3 13 1 11 2
16 9 1 0 9 11 3 13 9 2 15 4 13 9 1 11 2
9 9 7 9 1 0 9 3 13 2
25 3 13 3 15 9 0 12 9 1 9 1 11 10 9 3 2 16 13 9 1 0 15 0 9 2
24 1 0 15 9 9 11 2 15 13 12 2 9 12 2 13 9 1 0 9 0 1 0 9 2
13 9 9 0 0 9 13 3 9 0 9 1 11 2
30 1 0 9 0 9 2 9 2 13 7 1 9 9 0 9 2 16 4 13 13 3 0 9 2 14 12 12 9 12 2
16 9 0 9 13 1 9 11 9 1 9 11 1 9 1 11 2
14 1 0 9 11 15 9 13 10 0 9 1 0 9 2
11 9 2 9 9 7 9 2 7 0 9 2
11 9 1 9 1 9 13 9 1 0 9 2
22 13 15 2 16 16 13 9 9 2 13 0 2 16 3 13 1 9 1 9 12 9 2
31 0 13 0 9 0 9 2 9 13 1 9 0 7 0 9 0 9 7 0 9 1 15 13 9 2 3 2 0 9 2 2
37 10 9 13 13 9 2 9 13 15 15 2 13 9 1 9 0 7 0 9 2 7 13 15 9 2 7 13 0 9 1 9 7 1 0 9 2 2
23 0 9 0 9 2 9 13 0 9 2 1 15 13 1 0 9 13 9 0 9 0 9 2
37 1 0 9 2 1 15 13 9 9 2 13 9 9 9 2 0 9 7 0 9 7 13 15 1 15 3 13 9 7 9 2 9 7 0 0 9 2
68 1 0 9 9 2 15 15 13 13 7 9 1 0 9 2 3 13 0 9 0 9 1 2 9 15 9 2 7 9 13 0 9 2 2 13 2 16 15 15 9 9 2 0 1 9 0 9 1 9 9 2 13 7 14 2 0 9 1 2 9 2 2 13 2 9 2 9 2
119 1 0 9 13 0 9 2 3 0 2 7 3 0 9 9 2 11 2 0 9 9 11 2 0 9 1 9 2 9 11 2 15 1 11 3 13 9 2 15 9 2 2 13 15 2 16 13 2 14 10 9 1 10 9 1 9 16 2 9 2 0 9 2 13 4 10 0 0 9 13 1 15 2 2 7 0 9 10 9 2 0 9 2 16 1 2 9 2 13 0 9 9 7 13 4 13 1 9 2 3 13 2 16 1 9 13 1 9 7 3 14 1 0 9 2 2 2 2 2
46 1 9 9 13 3 13 14 3 0 9 9 11 7 9 0 9 2 9 1 0 9 9 2 15 13 2 3 3 13 1 9 1 0 9 2 15 15 13 13 0 9 9 7 0 9 2
22 1 9 9 15 13 13 3 0 7 3 0 9 9 1 15 15 2 13 2 15 13 2
18 1 2 9 9 2 13 1 9 13 2 16 13 0 1 9 10 9 2
32 9 13 13 0 2 7 3 15 3 15 2 1 9 2 13 13 3 1 12 9 1 0 9 2 1 0 9 13 15 2 9 2
6 9 1 9 11 7 11
2 9 9
15 0 9 0 9 0 15 9 0 9 13 1 11 12 9 2
22 9 0 9 2 11 2 13 0 9 2 15 13 3 1 9 9 7 4 10 9 13 2
23 0 9 13 9 1 9 0 9 2 11 2 0 1 0 0 9 2 15 9 4 13 9 2
9 9 12 9 15 1 10 9 13 2
12 9 1 0 9 13 1 9 13 1 12 9 2
23 3 13 13 2 16 1 9 9 11 13 1 15 15 0 9 1 15 3 16 1 9 11 2
22 13 15 0 3 1 0 9 2 9 7 1 0 9 15 1 10 9 13 3 7 11 2
11 9 13 13 3 9 9 1 3 0 9 2
39 13 2 14 0 9 9 1 11 2 16 13 2 7 13 13 2 16 15 9 13 2 3 15 1 9 13 1 10 9 7 1 10 9 15 3 9 3 13 2
16 9 11 7 3 13 13 2 3 4 13 2 16 4 13 13 2
9 10 9 13 9 9 3 15 9 2
26 1 9 9 12 9 13 13 2 10 0 9 13 0 9 13 1 10 9 0 7 3 0 13 10 9 2
17 0 9 9 13 2 16 0 9 13 11 2 11 7 11 2 11 2
12 9 9 0 9 7 11 13 1 15 3 0 2
15 7 15 1 9 1 9 2 16 0 9 13 7 0 13 2
11 0 9 1 9 12 9 13 3 13 0 2
20 0 0 9 11 13 0 9 9 11 7 9 9 0 9 1 3 16 12 9 2
21 9 11 1 0 9 9 9 9 3 13 7 11 3 13 1 12 9 1 12 9 2
10 10 9 13 13 13 0 9 9 0 2
32 9 9 11 13 3 1 12 0 2 7 10 9 13 3 0 1 0 9 3 13 9 1 9 9 16 11 7 3 13 9 9 2
18 9 12 9 15 3 1 10 9 13 2 7 13 1 9 0 7 0 2
7 13 1 0 9 12 9 2
25 1 1 15 2 16 11 13 0 9 0 3 1 9 10 9 2 13 10 9 3 0 7 3 0 2
3 9 0 9
14 0 9 0 9 13 1 3 0 7 0 9 1 11 2
20 0 9 15 13 3 0 9 2 7 7 0 9 2 16 3 1 9 13 9 2
16 0 2 3 0 9 13 0 9 2 0 0 9 1 0 9 2
18 1 9 9 13 9 2 16 2 10 9 13 1 10 9 1 15 2 2
13 0 9 15 9 13 16 0 9 1 10 0 9 2
41 1 2 0 9 2 1 0 2 9 3 13 7 0 9 0 9 2 9 1 9 7 0 9 2 0 7 0 9 2 7 7 0 9 9 0 9 7 9 1 9 2
33 0 9 0 0 9 13 3 3 0 9 2 15 1 9 13 0 9 13 3 9 13 1 9 0 9 7 9 3 13 0 9 9 2
24 1 9 2 16 15 13 3 0 9 1 11 2 15 7 13 7 9 9 7 9 0 0 9 2
16 10 0 9 4 9 2 15 13 1 0 9 2 13 1 9 2
11 3 15 13 1 9 2 16 9 9 13 2
23 9 9 7 9 15 1 15 3 13 13 1 9 2 16 4 15 9 13 1 9 0 9 2
12 1 0 9 13 9 3 3 2 16 13 0 2
17 0 9 14 1 9 13 2 16 0 9 15 1 0 9 9 13 2
14 0 1 15 13 9 9 2 9 7 9 9 1 9 2
11 0 9 14 13 9 0 9 13 3 9 2
17 0 15 3 13 13 9 0 9 7 0 9 2 15 1 9 13 2
13 13 7 15 2 15 13 0 0 2 9 3 0 2
30 3 13 3 1 0 9 0 7 9 2 9 2 3 10 1 9 0 9 2 13 3 15 13 9 0 9 1 0 9 2
8 3 15 1 15 13 7 9 2
1 9
27 0 9 13 13 1 9 9 2 15 15 13 1 9 16 9 1 9 9 2 9 10 9 2 16 4 13 2
21 9 3 1 9 9 1 11 7 1 11 1 11 12 13 7 1 15 9 1 11 2
29 9 9 11 1 9 11 13 1 9 12 0 11 2 15 13 1 0 9 1 9 9 2 7 13 1 12 9 3 2
22 9 1 9 11 1 11 12 2 0 9 13 9 3 1 12 11 11 2 2 12 2 2
13 0 9 13 2 16 9 13 3 13 9 1 9 2
22 9 9 11 12 9 12 2 12 0 9 15 1 9 13 12 0 11 11 2 1 11 2
11 1 9 15 9 13 1 0 9 0 9 2
7 0 9 1 9 1 11 11
2 0 9
2 11 2
10 1 9 1 11 11 15 13 0 9 2
22 9 9 12 11 11 2 15 3 13 16 9 2 13 1 0 9 1 11 1 12 9 2
21 15 13 1 11 1 9 12 2 3 3 13 1 9 9 1 9 1 9 9 11 2
9 9 13 14 1 9 3 10 9 2
17 9 13 9 9 2 15 11 13 9 10 0 9 2 7 9 11 2
23 1 9 11 13 2 16 0 9 2 15 13 2 4 15 13 13 1 0 9 7 0 9 2
16 13 1 15 2 16 9 1 10 9 13 2 7 1 9 13 2
21 3 13 2 16 9 7 9 13 0 2 16 4 9 9 13 9 2 15 15 13 2
23 1 9 15 9 13 7 1 9 0 9 9 9 11 11 2 15 1 9 13 16 0 9 2
17 11 2 11 13 2 16 11 13 1 9 9 11 1 0 9 11 2
34 11 13 13 3 2 1 9 0 9 7 0 9 1 0 9 0 9 1 0 7 1 9 9 1 11 1 11 1 9 3 12 9 9 2
6 9 1 9 11 11 13
2 0 9
2 11 2
21 0 9 1 11 13 3 0 9 1 9 11 11 2 15 4 13 1 0 0 9 2
22 11 13 1 9 12 1 11 12 13 3 1 0 9 12 9 7 1 9 12 15 0 2
10 9 9 13 3 1 9 12 12 9 2
28 11 10 9 3 3 13 1 12 9 9 9 2 7 0 9 9 13 1 9 1 9 9 7 13 9 1 9 2
24 1 0 9 15 13 2 16 12 1 9 2 15 16 0 11 13 2 15 13 1 9 10 9 2
14 9 3 3 13 1 9 9 2 1 15 4 0 13 2
16 9 9 7 0 13 3 2 1 0 9 7 1 9 1 9 2
6 9 13 7 12 9 2
12 9 13 2 16 9 9 13 7 3 13 0 2
27 0 9 13 0 1 9 1 9 9 7 9 15 15 7 13 1 9 13 2 16 2 1 15 13 9 2 2
13 0 9 3 13 2 3 9 13 1 9 0 9 2
19 10 9 0 9 13 1 12 9 2 16 9 0 1 9 12 9 13 0 2
14 9 0 9 15 13 1 10 0 9 2 16 11 13 2
20 9 0 9 13 12 1 0 9 0 9 2 9 2 15 13 3 1 9 9 2
14 15 13 2 1 12 9 2 9 9 13 1 9 9 2
12 3 15 13 1 0 9 7 13 1 15 9 2
18 10 9 3 1 9 13 2 16 11 13 9 2 7 3 15 13 0 2
5 13 9 1 9 9
2 11 2
27 9 1 3 16 9 9 13 0 9 0 9 12 9 2 15 15 1 9 9 13 0 0 9 1 0 9 2
11 13 1 15 3 0 9 0 9 11 11 2
21 9 1 9 12 7 12 9 13 0 9 13 1 12 2 9 7 13 15 0 9 2
9 13 15 9 0 9 7 13 9 2
5 13 9 1 0 9
2 11 2
20 9 13 1 9 12 0 11 11 2 1 11 1 11 7 13 15 7 0 9 2
25 9 13 1 9 2 0 3 1 9 12 1 0 9 7 0 1 9 9 9 1 9 0 0 9 2
30 1 9 9 13 11 11 2 1 0 9 0 9 7 9 0 7 0 9 7 9 2 9 9 7 9 15 9 0 9 2
33 0 0 9 15 13 0 13 15 2 16 3 2 16 12 2 9 12 13 0 9 1 9 7 9 9 1 11 2 1 9 9 13 2
13 0 13 9 9 9 14 1 12 9 7 9 0 2
6 9 3 13 1 0 9
2 11 2
26 3 0 9 9 1 9 7 9 13 1 9 0 9 9 0 9 9 9 9 2 1 15 9 3 13 2
15 12 12 0 13 2 16 0 9 13 13 10 9 1 9 2
14 0 1 9 9 13 9 7 9 2 3 0 13 9 2
12 11 11 4 16 9 3 13 3 15 9 9 2
14 13 15 12 12 9 7 9 2 9 0 9 7 9 2
13 13 13 7 1 9 3 0 9 1 9 7 0 2
22 13 9 14 1 9 0 9 2 7 7 1 9 0 15 1 0 9 7 3 1 9 2
10 0 13 10 9 7 1 9 7 9 2
13 9 11 4 13 16 9 9 0 9 2 3 11 2
18 13 15 9 0 7 0 2 10 9 13 1 9 7 9 1 0 9 2
12 3 9 13 1 9 2 15 15 13 0 9 2
11 7 12 1 10 12 9 13 12 9 0 2
18 1 9 9 15 13 1 0 2 9 2 0 9 7 9 1 0 9 2
20 0 9 13 11 2 15 13 1 0 9 2 7 3 15 13 10 9 1 9 2
17 1 10 9 13 9 9 7 9 2 7 7 9 9 13 3 0 2
9 11 15 13 16 9 9 0 9 2
11 13 1 0 9 1 0 9 7 1 9 2
13 13 15 10 2 0 9 2 7 10 9 1 11 2
11 3 0 0 9 11 1 9 3 13 0 2
22 11 2 11 2 0 1 9 0 9 9 0 7 9 2 13 9 7 1 0 0 9 2
10 9 9 7 9 1 10 9 15 13 2
15 9 13 9 1 9 1 0 9 7 3 15 13 1 11 2
7 0 11 13 9 0 9 2
14 9 9 1 10 9 15 7 1 0 9 13 14 3 2
13 3 15 3 13 9 10 0 9 1 9 7 9 2
5 11 13 0 9 0
3 1 0 9
2 11 2
27 9 0 1 0 9 9 11 11 13 2 3 0 2 9 0 9 2 11 2 2 15 15 13 3 1 9 2
13 13 15 1 9 9 9 11 11 1 0 0 9 2
22 2 3 0 2 13 11 0 0 9 1 9 9 7 1 0 2 0 9 2 13 11 2
12 2 13 3 0 9 0 0 9 2 2 13 2
23 11 13 2 16 9 1 0 9 13 9 2 16 9 11 7 9 0 9 7 9 4 13 2
20 11 1 11 3 3 16 1 9 13 1 15 2 16 0 9 13 0 9 9 2
12 11 13 1 0 9 2 9 9 15 7 3 13
2 11 2
36 9 9 11 11 2 11 2 13 13 2 16 15 0 9 12 0 9 1 0 9 1 9 13 9 14 1 9 0 9 2 7 7 1 0 9 2
31 16 3 13 11 2 13 1 9 9 9 2 15 4 3 16 3 13 9 13 1 9 1 15 2 16 13 1 9 7 3 2
19 11 13 2 16 15 13 1 9 0 0 9 2 3 1 2 9 2 3 2
34 1 9 1 9 2 15 4 15 13 13 15 9 1 9 2 13 9 13 9 3 12 1 12 12 0 9 7 10 9 1 9 0 9 2
17 1 9 1 9 15 13 13 3 0 12 9 2 3 3 12 9 2
14 9 13 2 16 0 9 13 1 9 3 1 0 9 2
15 13 15 1 9 9 1 9 2 15 4 13 13 0 9 2
22 1 0 9 0 9 11 13 11 9 11 11 9 2 1 15 10 2 0 2 9 13 2
18 1 9 3 0 9 11 13 0 9 0 9 0 11 11 7 13 11 2
22 11 3 11 13 2 16 16 4 13 0 9 9 0 9 2 2 15 1 15 13 2 2
29 9 0 9 1 9 11 11 2 11 2 11 2 15 13 2 16 9 13 3 0 2 16 4 9 0 11 13 13 2
25 2 13 15 2 16 9 1 9 13 10 9 7 16 9 1 9 0 9 13 0 13 2 2 13 2
13 11 11 2 11 2 13 0 9 1 9 1 0 2
20 13 15 7 2 16 15 2 15 11 13 2 3 13 3 13 7 13 1 9 2
26 2 13 0 0 9 2 7 13 13 0 9 2 2 13 0 9 2 16 4 9 13 1 9 1 9 2
29 11 13 3 0 9 0 9 7 9 9 1 9 2 3 7 7 9 2 15 4 15 13 9 1 3 0 9 9 2
11 13 3 9 2 16 0 9 13 0 9 2
7 9 0 0 9 11 13 0
2 11 2
24 1 9 0 0 9 11 11 11 4 9 1 0 9 13 1 0 0 9 13 3 9 0 9 2
10 15 4 15 13 13 1 0 0 9 2
35 9 0 9 1 9 2 0 0 9 2 2 15 9 3 9 0 9 13 9 0 0 9 11 2 13 11 1 10 9 1 2 3 0 2 2
15 1 3 0 9 4 15 1 15 13 13 14 9 0 9 2
20 2 13 15 2 16 4 9 3 13 13 0 9 2 15 4 3 13 0 9 2
16 3 4 15 13 13 1 9 1 0 0 9 2 2 13 11 2
10 9 0 9 3 3 13 1 0 9 2
33 2 10 9 15 4 1 10 9 13 7 10 9 3 1 9 0 9 13 1 9 2 2 13 15 9 0 9 0 9 11 11 11 2
21 2 13 2 16 9 0 0 9 4 1 9 13 13 0 9 2 2 13 9 11 2
13 1 9 0 9 4 13 9 13 1 10 0 9 2
25 11 13 2 16 1 9 9 9 2 0 9 2 1 9 9 13 10 9 1 0 9 9 1 11 2
29 0 9 0 9 11 13 1 11 1 9 2 15 13 1 0 9 0 9 2 15 4 15 13 13 0 9 1 9 2
9 9 7 3 13 1 9 1 0 9
2 11 2
17 16 9 13 9 9 1 0 9 2 13 15 9 9 1 10 9 2
9 0 9 13 1 9 1 0 9 2
33 13 15 1 9 9 11 11 11 1 0 14 3 0 9 1 0 9 1 11 1 11 2 1 15 13 13 1 9 0 1 0 11 2
19 0 9 15 13 13 7 9 2 15 9 13 1 12 2 9 1 0 9 2
34 9 9 15 13 13 13 9 9 0 9 2 1 10 9 15 12 9 0 13 2 16 13 0 2 16 4 15 9 13 1 9 0 9 2
17 9 13 3 1 9 1 0 9 2 13 15 15 7 7 9 11 2
29 3 7 9 0 2 12 9 2 13 1 0 9 1 9 0 9 9 1 9 2 15 13 12 1 9 9 3 0 2
17 1 9 9 1 9 0 9 13 3 11 11 7 9 1 0 9 2
4 0 9 13 13
2 11 2
29 9 0 9 9 9 11 15 1 9 1 9 0 9 13 13 9 9 1 9 11 2 11 2 11 7 9 0 9 2
30 9 1 0 9 15 13 1 9 11 2 11 2 11 2 2 15 13 1 9 9 0 9 2 3 3 13 0 0 9 2
21 11 1 9 13 3 2 16 12 9 0 9 1 0 9 13 1 10 9 9 9 2
24 1 10 9 4 1 9 9 13 7 9 13 3 0 9 2 7 15 11 11 2 0 1 11 2
43 9 11 2 11 2 11 7 9 0 9 2 15 13 1 0 9 9 2 13 1 9 11 2 11 15 3 0 9 9 2 16 4 15 9 13 7 15 15 13 13 0 9 2
26 10 9 7 4 13 7 11 2 11 4 1 0 9 9 11 2 11 2 11 12 2 11 7 11 13 2
9 9 1 0 9 11 7 11 13 0
2 11 2
37 9 0 9 1 9 0 9 9 0 9 2 11 2 7 9 1 9 0 9 2 11 2 13 1 10 9 3 0 2 16 4 15 13 0 3 13 2
24 9 11 11 11 15 13 2 16 0 9 10 9 1 9 12 9 13 3 0 16 10 0 9 2
17 9 1 10 9 13 13 1 10 9 13 0 9 9 3 1 9 2
19 2 15 2 1 9 1 11 2 13 0 9 13 10 9 0 2 2 13 2
13 9 13 1 10 9 13 7 1 0 9 9 0 2
29 3 9 11 11 11 15 13 2 16 0 9 2 15 15 13 0 9 3 15 9 1 9 11 2 13 13 9 9 2
13 2 3 13 9 0 15 7 3 11 2 2 13 2
19 13 2 16 9 13 13 13 7 0 9 0 2 15 1 10 9 13 11 2
23 1 11 7 9 1 0 9 13 0 7 1 9 13 0 13 2 15 1 15 13 3 9 2
4 9 1 9 12
7 11 1 9 9 1 9 9
3 1 0 9
2 11 2
28 9 9 1 9 9 4 13 13 7 9 0 9 0 0 9 13 15 1 9 12 9 1 9 9 9 0 9 2
15 1 9 11 11 2 11 2 15 13 13 0 9 10 9 2
10 16 9 13 9 1 9 0 0 9 2
15 0 9 15 7 1 11 13 13 2 9 2 1 0 9 2
34 16 9 9 9 1 9 3 2 9 1 9 0 9 13 13 1 9 10 0 9 2 9 0 9 15 4 3 1 9 13 2 13 9 2
13 9 0 9 13 1 15 7 9 2 7 0 9 2
20 13 7 2 16 13 1 15 2 15 1 9 1 9 9 4 13 13 1 9 2
9 9 13 1 12 2 9 9 13 9
2 11 2
44 0 9 13 1 0 9 0 9 0 9 9 12 2 9 9 0 0 9 2 15 13 1 0 9 7 0 9 3 12 2 9 1 9 9 9 2 9 0 0 9 7 0 9 2
9 13 15 3 9 9 11 11 11 2
20 1 9 1 9 0 9 13 2 16 9 1 10 9 4 13 13 12 9 9 2
50 0 9 4 13 10 9 2 15 13 9 9 11 11 2 11 2 2 9 9 11 11 2 11 2 7 9 9 11 11 2 11 2 2 13 1 0 9 1 9 9 9 11 11 7 9 0 9 11 11 2
33 0 9 15 1 11 13 1 15 2 16 4 15 15 0 0 9 13 1 9 9 7 16 4 4 13 12 9 1 9 9 7 9 2
26 1 10 9 4 15 13 9 0 9 12 2 9 2 10 9 11 13 0 9 1 12 9 2 13 11 2
19 9 1 15 13 9 2 9 0 9 1 9 2 1 9 12 2 9 9 2
4 9 13 1 9
2 11 2
25 3 9 9 13 9 3 3 13 9 0 9 0 12 9 1 0 9 0 2 9 2 9 9 9 2
6 9 1 9 13 0 2
32 13 13 1 15 7 1 9 0 9 15 1 0 9 9 7 13 15 2 16 15 1 9 3 1 9 13 9 1 9 9 9 2
16 2 0 9 13 9 9 1 9 9 15 1 12 9 0 9 2
17 3 1 0 9 15 13 9 7 9 1 9 1 12 3 1 9 2
22 0 9 1 0 9 7 9 13 9 9 0 9 2 3 7 9 2 15 13 0 9 2
28 16 9 7 9 9 2 13 15 13 7 0 9 2 4 13 1 15 0 9 1 3 0 0 9 2 13 9 2
8 1 9 3 9 15 9 13 2
21 1 0 9 13 9 9 9 2 9 9 2 2 13 9 9 11 11 0 9 9 2
18 15 13 0 0 9 2 12 2 9 2 7 3 4 13 1 12 9 2
29 2 1 0 9 9 9 7 10 0 9 1 9 13 9 0 9 0 2 9 2 9 2 2 13 9 9 11 11 2
11 9 3 13 2 10 9 15 14 13 1 0
2 11 2
7 9 0 9 13 0 13 2
11 1 15 15 13 9 9 2 9 7 9 2
16 12 1 9 2 3 15 13 2 13 7 9 0 0 9 9 2
8 9 4 13 13 3 12 9 2
20 13 15 0 9 9 9 1 9 2 15 4 10 9 13 0 7 0 9 9 2
20 9 9 11 11 1 9 13 2 16 10 9 13 16 0 0 9 3 12 9 2
24 0 9 9 9 4 13 1 0 7 15 2 16 0 0 9 13 1 1 9 9 3 0 9 2
24 9 13 2 16 4 15 13 13 14 12 9 9 2 16 4 9 13 10 0 9 1 9 0 2
11 15 1 15 13 14 12 9 1 10 9 2
13 9 15 3 13 2 16 13 3 7 10 0 9 2
19 9 15 3 13 2 16 9 13 3 10 9 7 3 14 3 13 0 9 2
16 0 9 0 1 0 9 0 1 0 12 9 3 13 0 13 2
8 9 4 1 15 13 13 9 2
14 9 9 2 15 13 10 9 2 15 3 13 1 0 2
10 9 15 9 13 7 1 10 0 9 2
24 15 13 9 10 9 2 7 3 0 9 11 11 13 1 0 2 16 4 13 15 13 1 0 2
11 0 9 4 3 13 13 3 9 1 9 2
15 1 10 9 10 9 13 2 16 4 15 14 13 0 9 2
19 3 13 3 3 3 13 2 1 10 9 9 13 2 16 15 9 3 13 2
9 1 0 9 9 13 3 1 0 9
2 11 2
22 9 15 2 15 13 2 16 9 13 1 10 9 10 9 2 13 9 1 9 1 9 2
26 1 10 9 15 1 0 11 13 9 3 1 12 9 9 2 1 0 9 2 1 9 7 1 0 9 2
14 1 0 9 0 9 13 9 12 9 1 0 0 9 2
16 1 9 15 13 3 0 9 2 15 7 13 15 0 1 9 2
9 13 1 9 1 0 0 0 9 2
5 13 3 12 9 2
22 13 15 3 2 0 9 2 2 15 13 3 1 9 0 9 2 7 3 9 1 9 2
14 1 9 7 9 13 13 7 0 9 3 7 3 13 2
15 11 13 1 0 9 9 1 9 1 10 0 7 0 9 2
33 13 1 15 2 16 16 3 1 11 13 9 1 0 9 3 0 7 1 11 15 3 3 13 9 2 1 11 7 1 11 9 13 2
25 9 7 13 3 0 2 1 0 9 1 9 12 7 12 9 3 2 7 13 3 3 9 0 9 2
20 0 9 1 0 9 1 0 0 9 13 3 3 12 9 2 1 0 1 12 2
23 1 11 13 9 1 0 0 9 0 2 9 7 13 13 9 1 0 2 0 7 0 9 2
18 9 13 2 16 10 9 13 9 9 0 1 0 9 7 13 0 9 2
11 1 0 0 9 15 7 13 0 9 9 2
23 3 1 0 0 9 9 7 9 13 14 9 12 0 9 7 1 0 9 15 13 12 9 2
10 0 9 1 9 9 13 1 9 1 9
2 11 2
20 0 9 11 1 0 0 9 0 2 0 9 13 3 9 9 9 7 9 9 2
16 13 1 9 0 9 2 3 13 9 2 1 9 9 12 2 2
8 13 15 3 16 12 12 9 2
16 9 13 0 9 9 2 9 2 9 7 9 9 0 0 9 2
32 9 13 9 1 9 1 9 12 0 9 2 15 7 1 9 9 0 9 3 13 1 0 9 7 0 7 0 9 1 9 9 2
18 9 7 13 0 9 0 9 2 15 4 13 9 13 1 10 0 9 2
20 7 7 15 13 1 9 9 9 11 11 1 9 2 16 13 0 9 9 9 2
28 11 11 1 9 0 9 11 3 13 2 16 0 9 0 9 3 13 1 0 9 7 13 0 9 3 0 9 2
33 13 3 9 0 9 9 0 9 2 1 11 15 7 13 14 1 9 0 2 0 9 9 2 3 1 9 2 0 9 7 9 2 2
27 3 9 0 7 0 9 1 11 11 2 15 15 13 9 9 0 9 2 11 11 13 0 0 9 1 0 2
5 0 9 13 13 3
2 11 2
14 0 0 9 13 3 10 0 9 13 3 1 10 9 2
22 16 0 9 9 9 9 7 13 2 16 4 9 1 9 0 9 4 13 1 0 9 2
12 0 9 3 13 13 9 1 0 9 7 9 2
13 3 15 13 3 1 11 2 15 10 9 9 13 2
10 9 0 3 13 0 9 13 1 15 2
23 9 0 9 2 0 1 0 9 9 1 11 2 13 9 9 7 9 9 0 9 9 1 9
5 9 13 9 1 9
2 11 2
18 14 1 12 9 13 3 9 9 1 9 11 9 0 1 0 9 11 2
20 13 15 0 9 1 9 9 2 9 7 0 9 2 1 15 3 13 12 9 2
27 1 0 9 13 0 9 9 2 15 13 1 9 9 2 9 9 9 1 0 9 3 1 9 1 0 9 2
26 3 3 3 2 13 9 9 11 2 15 4 13 3 1 0 9 2 7 13 1 9 1 9 7 9 2
14 9 2 15 13 3 1 12 2 13 1 9 1 12 2
7 9 13 9 1 9 1 9
2 11 2
30 9 9 2 12 0 9 0 9 7 9 2 15 9 13 2 15 13 3 3 7 3 1 9 1 9 1 0 9 9 2
11 3 3 9 13 3 9 1 10 0 9 2
35 13 15 3 9 1 0 9 1 9 9 7 9 2 15 4 13 3 1 0 9 2 7 3 0 0 7 0 9 2 15 13 0 9 9 2
9 10 10 9 13 1 9 1 9 2
22 1 9 13 7 9 0 13 9 9 3 3 2 7 3 15 9 13 1 0 0 9 2
18 3 9 9 11 13 7 1 12 12 9 2 13 15 7 13 1 9 2
14 9 2 15 13 0 0 9 2 13 3 1 9 7 9
10 1 0 9 7 13 3 9 15 13 2
29 9 1 12 0 9 13 1 9 3 12 9 2 9 1 9 12 9 7 1 9 1 0 9 13 0 13 12 9 2
2 0 9
19 1 12 2 9 10 9 1 0 9 13 12 9 9 1 0 9 0 9 2
28 3 1 15 3 12 9 2 1 15 3 9 13 2 7 10 9 14 3 1 0 9 13 1 9 9 0 9 2
12 0 9 0 9 3 1 9 13 0 9 12 2
12 0 9 3 3 13 2 10 0 9 9 13 2
18 9 3 13 9 9 0 1 0 9 2 1 15 15 3 1 9 13 2
23 1 15 13 0 9 2 0 2 0 9 2 13 1 9 0 1 0 9 1 12 2 9 2
7 13 3 1 0 0 9 2
40 1 9 9 0 9 0 9 15 9 13 1 9 2 15 13 1 9 9 9 7 9 1 0 9 2 3 0 9 10 10 0 9 2 7 3 0 9 1 9 2
22 0 9 13 13 10 0 9 2 7 13 2 1 9 9 9 2 13 3 1 9 9 2
13 13 15 2 16 0 9 4 13 1 3 0 9 2
18 14 1 0 0 9 13 3 0 3 13 9 14 1 12 9 12 9 2
21 1 9 9 15 3 9 4 3 3 13 7 1 9 9 3 9 13 3 3 3 2
19 3 1 9 9 2 0 9 2 15 9 0 0 9 13 1 0 12 9 2
18 0 13 0 9 1 9 2 3 15 13 0 2 9 7 15 13 9 2
20 3 10 0 9 13 9 0 0 9 2 3 9 3 0 9 0 10 0 9 2
29 16 1 0 2 9 0 9 15 0 9 13 12 9 9 2 1 9 13 10 9 12 9 2 13 3 3 3 0 2
29 0 9 1 9 0 9 1 9 7 0 2 9 13 1 9 2 16 0 1 10 12 0 9 13 1 0 9 9 2
37 7 1 10 12 9 7 3 3 13 1 0 0 9 2 7 3 9 2 9 2 16 0 9 3 15 13 2 7 7 13 2 1 12 3 0 9 2
13 0 9 15 3 13 12 1 0 9 10 0 9 2
7 15 13 15 2 16 3 2
6 9 0 16 0 2 11
15 15 13 13 0 9 1 9 1 0 9 2 13 4 15 13
2 11 2
21 3 3 16 0 2 9 13 9 0 9 0 9 3 0 9 1 0 9 0 9 2
25 9 2 15 13 13 0 9 1 12 9 2 13 3 3 13 0 9 1 0 2 11 7 13 9 2
18 1 9 15 13 13 1 9 12 7 12 7 0 16 1 0 2 11 2
7 13 15 1 9 12 9 2
26 16 0 9 1 0 2 11 9 11 15 4 0 9 13 1 12 9 2 1 9 13 10 9 12 9 2
18 9 9 4 1 0 2 11 13 1 12 9 7 1 9 1 12 9 2
18 0 9 0 11 13 1 9 12 9 7 1 0 2 11 13 12 9 2
16 15 1 0 9 13 1 9 1 9 0 16 12 9 1 9 2
17 0 9 1 0 2 11 13 0 0 9 1 9 12 9 1 9 2
9 1 9 15 13 13 1 12 9 2
21 13 7 13 9 1 0 9 0 9 13 0 0 9 2 15 15 13 1 0 9 2
31 14 7 3 16 1 9 12 2 9 2 3 9 0 9 13 10 0 9 2 1 15 13 1 9 9 3 9 1 0 9 2
24 0 9 13 13 10 9 3 1 9 11 2 1 0 9 0 2 9 7 9 0 9 1 9 2
19 1 9 13 0 2 11 9 1 9 7 9 0 9 1 9 1 0 9 2
10 0 9 15 13 12 2 9 1 9 2
16 1 9 15 3 13 13 3 10 9 2 7 3 1 0 9 2
14 2 15 7 13 3 0 2 2 13 9 9 11 11 2
15 1 9 1 9 13 0 13 0 2 0 9 1 0 9 2
17 15 3 13 9 0 9 1 11 7 1 9 9 15 13 1 9 2
11 0 9 0 9 1 9 13 3 1 9 9
6 9 9 13 1 9 0
2 11 2
16 0 0 9 1 9 4 3 13 0 12 7 3 3 12 9 2
14 13 15 1 0 9 2 15 3 9 13 9 9 9 2
14 1 10 9 15 13 13 9 1 0 9 9 0 9 2
29 9 13 1 0 9 12 9 3 7 13 2 16 15 9 1 9 13 9 10 9 2 16 0 15 13 1 0 9 2
17 9 13 13 12 9 1 9 0 9 7 4 15 13 3 12 9 2
21 13 15 1 12 5 9 2 12 5 0 9 9 7 12 5 9 1 9 1 9 2
23 3 1 0 9 1 0 9 12 2 0 9 1 0 9 9 7 12 2 9 1 0 9 2
29 1 0 9 13 0 0 9 12 9 2 15 4 13 13 12 5 9 1 0 9 9 7 12 5 9 1 0 9 2
25 13 1 0 9 9 0 9 0 9 15 13 0 0 9 12 9 1 9 9 7 12 9 1 9 2
5 0 9 1 9 12
10 9 9 1 9 13 2 1 9 3 13
2 11 2
21 9 11 11 15 13 9 12 9 9 2 16 9 1 9 11 11 13 1 12 9 2
10 1 9 13 12 9 3 0 0 9 2
18 9 0 9 2 11 2 13 1 10 9 1 9 0 9 1 12 9 2
21 1 9 9 11 13 9 3 1 9 7 10 9 1 9 0 9 2 3 0 9 2
21 0 9 11 3 13 2 16 3 2 16 13 9 1 9 2 13 7 9 1 9 2
25 3 13 3 1 15 3 16 9 0 9 13 1 0 9 9 7 14 12 9 9 13 3 9 9 2
21 11 1 10 9 13 1 0 9 0 9 9 1 0 9 2 16 0 9 13 9 2
4 3 1 9 12
3 11 13 11
2 11 2
21 9 9 0 0 9 11 13 0 0 9 13 1 9 2 0 9 2 14 1 9 2
9 11 15 13 9 11 11 2 11 2
20 9 9 9 9 7 9 2 11 7 0 11 1 9 4 13 4 13 1 9 2
22 11 13 9 11 11 2 11 1 10 9 9 3 2 16 13 4 13 1 9 0 9 2
7 9 1 11 14 1 12 9
2 11 2
27 9 0 9 11 11 11 13 3 1 9 1 9 9 1 0 9 9 9 9 0 9 1 11 12 11 11 2
14 15 13 2 16 1 0 9 13 1 12 7 12 9 2
19 9 13 9 0 9 1 9 7 13 2 16 9 9 1 0 9 13 9 2
13 16 13 9 11 0 2 13 15 14 12 9 9 2
5 11 2 11 3 13
2 11 2
15 0 9 0 9 1 0 9 13 3 14 1 12 9 3 2
10 0 9 13 1 9 7 9 7 9 2
16 9 4 13 1 0 9 9 1 9 1 0 9 0 9 11 2
17 1 9 0 9 9 11 11 15 0 9 3 13 13 0 9 9 2
25 1 11 13 3 3 13 9 1 0 7 0 0 9 2 7 0 9 3 0 9 0 0 9 13 2
23 0 9 0 9 13 0 9 0 9 2 15 15 13 3 3 3 3 2 16 11 13 9 2
14 9 13 1 9 9 11 7 1 9 1 9 1 11 2
4 3 1 9 12
5 11 1 0 9 11
2 11 2
24 11 13 1 9 13 11 0 0 9 2 15 4 13 10 9 1 9 11 13 15 1 0 11 2
7 13 15 1 11 9 9 2
30 9 14 3 1 9 13 0 9 11 7 13 13 13 1 9 11 11 2 15 13 3 13 0 0 9 9 9 9 11 2
19 1 0 9 9 3 13 9 1 9 0 0 9 1 9 1 11 7 9 2
25 0 9 13 13 13 11 9 2 1 15 13 1 9 2 3 11 13 9 13 9 1 9 1 9 2
39 1 9 11 9 11 13 9 13 3 0 0 9 2 7 13 13 9 1 15 2 16 4 11 13 9 9 1 11 2 15 13 3 13 1 10 9 9 9 2
5 9 13 0 0 9
2 11 2
32 9 0 0 9 2 15 4 13 13 12 1 0 9 9 1 9 1 9 7 9 0 9 0 0 9 2 13 9 0 0 12 2
23 13 15 1 9 9 9 2 0 9 0 9 0 11 11 11 2 1 12 2 9 0 9 2
35 1 9 7 9 9 9 13 1 0 2 3 0 9 1 9 9 0 9 2 0 9 2 9 0 9 2 1 0 9 7 9 3 1 9 2
29 13 3 1 11 2 9 9 7 9 11 2 9 9 0 2 0 2 11 2 2 0 9 11 7 10 0 0 9 2
12 9 13 3 0 1 9 0 1 0 0 9 2
19 9 13 1 11 0 9 1 9 9 7 15 13 10 9 7 9 3 13 2
13 1 9 15 1 15 13 13 10 0 9 7 9 2
25 1 9 9 1 0 9 13 9 9 12 2 1 9 9 1 9 12 13 1 9 0 9 0 9 2
23 1 9 9 0 0 12 13 1 11 3 13 2 9 1 9 7 1 9 9 13 1 9 2
5 0 9 13 9 9
10 0 9 0 9 4 13 14 1 9 12
2 11 2
20 0 9 0 2 0 9 2 15 13 0 9 11 2 13 1 0 9 3 13 2
15 1 9 11 9 2 11 11 9 13 0 9 1 12 9 2
8 0 9 13 12 9 9 9 2
15 3 0 9 13 9 0 9 2 0 9 13 14 12 9 2
28 1 0 0 9 2 15 7 3 9 13 2 4 1 9 12 9 9 13 3 12 9 9 2 3 12 9 9 2
8 9 9 13 1 0 9 9 2
30 9 9 7 9 11 11 0 9 1 11 13 2 16 0 9 2 15 0 9 13 1 0 9 9 2 13 1 9 12 2
20 1 15 4 1 10 9 13 4 13 1 9 9 2 3 1 9 1 9 9 2
17 0 2 9 2 11 4 13 4 9 9 13 9 14 12 9 9 2
10 3 3 4 13 3 16 12 9 9 2
10 13 13 4 0 9 9 11 7 11 2
11 9 9 12 9 9 11 1 11 4 13 2
19 1 9 13 9 1 9 1 9 9 11 1 9 12 7 9 1 9 12 2
18 1 9 11 15 3 13 0 9 9 1 9 9 0 9 7 0 9 2
13 1 15 13 11 0 9 2 9 11 7 11 11 2
11 13 13 7 9 3 13 9 1 0 9 2
27 0 0 9 1 11 3 1 0 9 7 0 9 9 9 1 11 13 9 9 2 15 9 13 1 0 9 2
15 3 0 4 1 11 13 13 7 0 9 9 2 0 9 2
3 9 9 13
8 9 13 7 0 11 1 0 11
2 11 2
20 0 0 9 0 9 1 9 13 1 12 9 9 2 1 12 9 1 0 9 2
11 13 15 1 9 0 9 1 9 7 9 2
27 1 0 11 16 9 13 9 9 1 12 9 1 12 9 9 7 1 0 9 1 12 9 1 12 9 9 2
22 1 9 1 9 9 12 13 9 9 1 11 3 1 12 9 0 7 13 12 9 9 2
54 1 0 11 1 0 11 13 0 9 0 9 12 9 9 2 1 12 9 3 16 1 9 2 16 0 9 1 0 9 11 13 1 12 9 9 2 1 12 9 1 0 9 2 7 13 1 12 9 0 16 1 9 12 2
5 1 11 13 0 9
2 11 2
19 1 0 9 15 3 13 0 9 7 9 0 9 15 13 1 0 9 9 2
27 9 9 0 9 1 9 13 2 16 0 9 3 1 2 0 0 7 0 9 2 13 3 0 9 0 9 2
23 9 9 1 0 9 0 9 13 1 12 1 12 9 7 1 0 9 15 13 10 0 9 2
18 1 0 9 0 9 13 3 11 2 15 15 13 14 0 12 9 9 2
24 1 12 0 0 9 1 11 13 3 11 12 2 11 11 2 11 12 2 11 11 7 11 11 2
9 3 1 0 9 13 0 11 12 2
23 9 13 1 0 9 1 0 9 0 11 2 3 13 3 3 1 9 12 11 7 12 11 2
5 13 9 1 12 9
2 11 2
17 3 1 12 9 1 11 7 1 11 13 9 0 9 0 9 11 2
24 10 9 1 0 9 13 1 0 9 3 12 9 9 2 9 1 9 4 13 1 12 9 9 2
20 3 4 15 13 9 13 1 12 9 9 7 9 4 13 13 1 9 9 12 2
4 11 13 0 9
2 11 2
18 11 1 9 9 9 0 9 13 1 9 12 0 0 9 1 0 9 2
18 13 15 1 0 9 9 2 0 9 2 2 15 1 9 13 0 9 2
30 1 10 9 4 9 1 9 12 13 9 0 0 0 9 1 0 9 2 10 2 0 9 2 3 4 13 1 9 12 2
16 9 3 13 9 0 9 2 16 13 9 2 9 7 0 9 2
22 4 3 13 1 9 1 9 0 0 9 2 15 9 4 13 9 9 1 9 0 9 2
3 9 13 0
2 11 2
20 1 0 9 13 9 1 0 0 9 0 7 1 10 0 9 1 0 0 9 2
11 0 9 13 0 9 9 1 9 0 9 2
32 3 1 9 15 9 13 1 12 9 2 3 1 0 0 9 12 9 7 3 1 9 12 9 2 1 15 1 9 13 1 11 2
21 9 0 9 15 1 9 3 9 13 1 9 0 0 9 2 0 9 7 0 9 2
8 15 15 13 1 9 0 9 2
22 9 13 1 9 1 0 9 12 9 7 0 9 13 1 12 0 9 12 9 1 9 2
9 1 0 9 15 4 7 3 13 9
2 11 2
21 1 12 9 2 15 13 14 12 9 2 13 3 13 0 0 9 9 0 9 11 2
18 0 0 9 1 0 9 13 1 9 9 12 1 9 0 9 12 7 2
7 15 13 9 1 12 9 2
17 1 15 1 9 12 13 0 0 9 9 1 0 9 14 12 9 2
10 0 0 9 9 0 9 13 12 9 2
13 9 9 1 0 9 11 13 1 0 1 0 0 9
6 0 9 13 12 9 2
8 0 9 9 13 12 9 9 2
14 0 9 13 12 9 9 7 9 13 12 9 15 9 2
9 0 9 0 9 13 12 9 9 2
8 0 9 9 13 1 12 0 9
5 10 9 15 13 2
12 13 2 14 3 9 2 13 13 9 0 9 2
5 9 4 13 12 0
2 11 2
27 9 1 9 0 9 4 1 9 0 0 9 13 3 12 1 3 12 12 9 7 1 9 0 9 3 12 2
26 3 12 0 9 1 0 9 13 1 0 9 0 16 12 9 7 12 0 4 13 1 9 1 12 9 2
21 0 9 1 12 7 12 9 4 13 12 0 2 0 9 13 0 3 1 12 9 2
24 0 0 9 4 13 12 9 0 2 0 9 12 9 7 3 9 0 9 13 12 9 9 9 2
17 1 9 0 0 9 16 0 7 0 9 13 9 3 16 9 0 2
16 0 9 9 1 15 4 15 13 12 9 2 0 12 9 0 2
6 0 9 11 13 1 9
2 11 2
28 0 9 1 11 13 1 9 12 2 9 13 0 9 11 2 15 13 0 9 11 11 2 7 13 3 0 9 2
18 0 7 3 0 9 9 1 9 7 9 13 13 1 12 9 2 9 2
12 9 9 1 9 13 9 0 9 1 0 9 2
33 0 9 1 9 0 9 13 9 12 9 2 9 1 12 9 2 12 9 1 12 9 2 9 1 12 9 7 0 9 1 0 9 2
11 4 13 1 12 9 7 9 13 9 9 2
8 1 9 1 11 15 13 7 11
2 11 2
14 11 15 3 1 9 13 0 9 9 11 1 0 11 2
12 9 0 9 15 1 9 4 13 1 0 9 2
14 1 9 0 9 13 9 10 9 13 1 9 0 9 2
12 0 9 9 11 15 13 1 11 1 9 12 2
13 3 15 1 9 13 3 16 12 9 1 12 9 2
12 0 9 15 13 1 12 2 1 12 2 9 2
6 1 0 9 13 3 9
14 1 3 0 0 9 1 11 15 4 0 9 13 1 9
22 9 0 0 9 2 3 1 9 9 2 15 3 13 14 1 11 2 7 7 1 11 2
15 0 0 9 1 0 9 13 1 0 7 0 9 7 9 2
17 1 9 3 13 7 0 9 2 15 13 0 1 9 7 0 9 2
21 13 10 9 1 0 9 13 9 11 2 11 9 9 2 2 15 9 13 9 11 2
35 9 11 13 9 12 12 9 0 0 0 7 0 9 1 0 9 2 0 9 1 9 7 12 0 9 1 12 9 0 9 3 1 9 11 2
11 9 13 13 1 9 9 2 9 7 9 2
16 9 9 4 13 3 3 1 9 7 13 13 4 3 1 9 2
18 0 9 9 4 13 9 1 9 9 12 7 9 9 3 1 9 3 2
16 9 9 11 13 2 16 0 9 13 1 12 9 3 3 13 2
15 9 9 1 9 13 2 16 9 13 9 9 7 9 3 2
17 0 9 13 9 9 13 3 1 9 2 7 9 0 9 13 0 2
34 9 9 13 0 1 0 14 1 0 2 0 9 1 9 0 9 2 0 9 0 9 2 0 11 2 9 2 0 9 2 9 7 9 2
13 0 9 4 13 9 2 3 15 13 10 0 9 2
18 4 13 1 9 0 9 0 0 9 7 9 1 0 9 1 0 9 2
23 9 9 11 13 13 3 2 16 4 9 13 0 9 1 0 9 1 3 0 9 1 11 2
15 1 9 0 9 13 9 9 11 1 0 9 11 7 11 2
16 9 9 11 13 1 15 9 0 9 1 9 1 11 7 11 2
13 1 9 0 9 13 9 9 9 9 1 10 9 2
15 11 7 13 9 1 11 1 9 9 1 12 7 12 9 2
23 1 9 9 9 15 13 1 9 0 0 9 12 12 9 2 0 9 12 7 0 12 9 2
16 1 9 9 13 9 11 0 9 1 9 0 1 9 11 12 2
22 3 9 13 12 7 12 9 2 7 2 14 12 9 7 12 9 1 9 0 7 9 2
31 1 0 0 9 15 9 9 1 12 9 0 13 1 12 1 12 9 3 2 15 1 9 13 12 9 7 12 9 1 9 2
28 1 0 9 9 13 0 0 9 9 1 9 9 12 9 3 1 9 1 12 12 1 12 12 9 1 9 0 2
13 9 0 9 13 1 11 1 9 3 16 1 11 2
30 3 0 0 9 2 0 1 9 11 2 13 9 0 9 0 9 1 12 9 3 2 3 12 9 1 9 7 9 0 2
18 1 15 0 0 9 1 0 9 4 13 1 12 12 9 1 9 0 2
19 1 9 9 11 13 0 9 9 1 0 11 3 3 0 16 0 1 11 2
17 0 9 15 13 9 13 3 2 16 4 13 9 9 1 0 9 2
38 0 9 2 15 3 13 1 9 9 7 3 0 9 2 13 2 16 13 3 16 9 2 7 2 9 2 7 3 0 9 9 7 15 15 13 7 9 2
45 1 9 9 15 13 9 2 15 13 0 9 13 9 2 7 7 13 1 9 9 16 1 0 9 2 7 1 9 9 2 9 2 9 2 0 7 0 9 2 9 2 9 7 9 2
5 0 9 13 9 2
2 11 2
30 0 9 1 0 2 0 9 13 0 9 3 1 9 0 12 9 9 2 7 16 1 9 0 1 12 1 12 9 9 2
24 0 9 9 13 14 1 9 0 9 9 2 7 7 1 9 0 9 2 15 9 9 3 13 2
37 9 9 15 13 1 12 1 12 1 12 9 9 2 9 1 9 13 1 12 1 12 9 9 7 9 0 9 15 13 1 12 5 1 12 9 9 2
1 3
15 11 4 15 1 9 0 9 13 13 9 0 9 0 9 2
12 9 1 11 13 1 10 9 9 1 0 9 2
18 0 9 1 11 3 13 1 9 9 9 0 9 11 11 12 9 9 2
15 1 9 12 10 9 13 12 9 7 1 9 12 12 9 2
21 9 0 9 13 9 1 12 9 9 2 15 4 3 13 0 9 1 9 0 9 2
11 0 9 13 1 0 9 1 0 9 9 2
11 0 0 9 1 10 9 13 1 12 9 2
9 1 0 9 9 13 1 12 9 2
13 9 11 1 9 12 9 9 13 9 9 0 9 2
19 9 10 9 13 9 9 1 0 2 0 2 14 2 9 1 0 0 9 2
5 0 9 13 0 9
7 9 0 9 13 0 0 9
10 11 2 11 13 12 2 12 5 9 9
2 11 2
24 0 9 13 1 15 9 0 9 2 15 4 1 0 9 13 13 0 16 1 0 9 0 11 2
24 13 15 1 9 10 9 1 0 9 1 0 9 1 0 9 2 15 3 13 1 0 9 11 2
22 1 9 9 7 9 11 11 13 0 9 7 3 9 1 0 9 9 7 0 9 9 2
17 9 1 10 9 13 10 9 7 13 0 9 1 0 9 1 11 2
25 0 9 4 1 11 2 11 13 1 9 9 10 0 9 13 3 1 0 7 0 9 14 0 9 2
26 11 2 11 13 2 16 9 13 1 0 9 0 9 1 9 12 9 9 0 9 2 0 9 7 11 2
48 1 9 1 11 0 9 1 9 13 3 1 10 0 9 9 11 11 2 16 13 2 16 0 9 9 15 3 12 9 13 1 0 9 7 1 10 9 1 9 7 9 13 1 10 0 0 9 2
24 1 0 9 4 9 13 1 9 13 1 0 0 9 2 3 13 0 9 13 1 0 9 9 2
22 1 9 9 9 0 0 9 11 11 13 0 0 9 1 11 1 0 9 12 9 9 2
26 16 1 9 1 0 9 13 9 9 9 11 11 2 9 4 13 0 0 9 9 9 7 9 1 9 2
29 0 9 7 13 1 15 2 16 9 13 1 15 2 3 15 3 13 0 9 2 15 4 13 9 1 0 9 13 2
21 11 11 0 9 13 2 16 0 0 9 3 1 0 9 13 1 12 2 12 9 2
31 9 2 15 3 13 12 9 2 4 1 10 9 13 3 13 1 12 7 12 0 9 3 14 1 12 9 1 9 0 9 2
13 9 9 4 1 12 9 13 13 12 7 12 9 2
22 0 9 9 2 1 15 3 13 0 9 1 0 9 2 3 13 0 9 9 12 9 2
20 9 9 1 12 7 12 9 13 1 9 11 1 10 0 9 3 0 0 9 2
20 0 9 13 9 3 1 0 9 2 15 13 9 3 1 9 9 3 13 9 2
30 0 9 1 9 1 12 7 3 9 13 1 9 11 2 11 13 3 3 16 0 9 0 1 9 9 7 0 9 9 2
17 9 2 15 3 13 9 0 9 2 13 13 9 14 1 12 9 2
17 2 15 4 13 13 0 1 0 9 2 15 13 9 2 2 13 2
31 1 9 15 9 1 0 9 13 9 9 2 9 7 9 2 9 0 0 9 7 1 10 0 9 3 7 9 9 0 9 2
10 9 1 9 0 9 2 13 2 9 9
2 11 2
17 0 9 9 0 0 9 2 13 2 9 0 0 9 2 3 9 2
31 1 9 15 13 1 0 9 9 2 15 14 3 13 1 9 0 0 0 9 7 0 9 0 9 1 9 9 11 1 11 2
22 9 1 9 1 9 13 1 0 9 9 0 9 0 0 9 2 1 15 11 3 13 2
17 1 9 9 15 13 1 0 9 9 12 2 3 7 1 9 12 2
18 9 13 2 16 1 0 9 4 9 1 0 9 13 3 1 9 12 2
30 1 9 0 9 0 0 0 9 2 0 9 7 11 13 9 3 2 13 0 9 9 0 1 2 9 2 1 9 9 2
22 0 9 3 0 9 3 1 9 2 16 3 15 1 9 13 3 1 10 3 0 9 2
20 15 0 9 4 1 9 0 9 13 1 0 0 9 7 0 0 9 0 9 2
5 0 0 9 1 9
2 11 2
28 0 9 3 3 13 1 9 11 13 1 9 9 1 9 10 9 1 2 9 2 7 13 15 9 3 13 9 2
41 9 0 9 13 2 16 9 13 10 9 1 0 9 0 9 1 9 2 9 2 9 7 0 9 7 16 13 10 9 2 15 13 1 9 0 0 9 1 0 9 2
48 11 13 13 0 9 1 12 2 9 1 9 1 15 2 16 13 1 11 9 2 15 15 3 16 0 9 1 0 0 9 13 3 2 16 15 1 9 11 13 1 2 9 2 1 2 9 2 2
13 9 0 9 13 9 11 1 9 2 7 10 9 2
5 0 9 11 13 9
2 11 2
25 0 0 9 11 2 15 1 9 13 9 9 9 2 13 13 0 9 1 0 9 1 12 2 9 2
28 9 13 9 0 2 0 2 0 2 15 1 9 0 7 0 2 2 0 9 1 9 0 2 9 7 0 9 2
18 9 2 15 13 13 1 9 0 0 9 2 13 0 1 15 9 9 2
28 0 9 9 2 15 9 13 1 0 0 9 11 11 2 13 12 9 9 2 16 0 9 13 0 12 9 9 2
4 0 0 13 9
2 11 2
16 0 9 0 0 9 1 9 12 13 1 0 9 12 9 9 2
15 0 9 13 3 12 9 1 12 9 1 0 9 12 9 2
16 1 9 12 13 0 0 9 9 12 9 9 7 9 13 4 2
27 9 9 1 12 2 9 12 13 12 9 9 2 15 13 1 9 1 9 1 9 9 9 3 1 12 9 2
15 9 7 3 2 13 1 9 9 0 9 2 13 3 3 2
11 11 13 1 11 9 2 11 15 13 0 9
2 11 2
9 9 0 9 13 13 1 0 9 2
26 13 1 15 9 0 9 2 15 15 1 11 11 1 0 9 7 11 11 1 9 11 13 1 0 9 2
19 1 10 9 13 9 11 11 1 9 9 0 15 9 2 15 13 9 11 2
20 1 11 11 3 2 13 2 16 11 13 9 9 2 7 16 1 15 13 3 2
19 1 9 9 11 13 3 1 11 2 11 13 2 16 9 0 9 11 13 2
15 11 13 2 16 11 1 9 12 13 3 16 1 9 12 2
14 1 9 3 13 13 13 9 1 2 0 9 2 11 2
8 11 15 13 2 16 9 13 2
21 2 9 11 13 3 12 9 2 9 2 15 13 0 9 9 9 11 2 2 13 2
20 1 9 13 9 13 11 1 11 11 13 2 16 0 9 13 12 5 9 11 2
8 15 14 7 13 0 12 5 2
16 2 13 15 13 0 9 3 16 16 0 9 2 2 13 11 2
8 3 1 9 13 9 9 11 2
24 2 1 9 13 9 4 3 7 1 9 13 9 1 9 2 3 1 9 0 9 4 13 9 2
10 9 9 3 13 9 2 2 13 11 2
19 15 9 4 13 1 0 9 11 7 0 0 9 11 2 13 9 9 11 2
24 9 1 9 9 11 4 1 11 7 1 12 9 13 3 2 3 4 13 1 9 11 2 11 2
12 2 11 3 13 9 1 9 0 9 7 9 2
13 13 7 0 0 9 0 9 2 2 13 9 11 2
12 11 15 3 13 1 9 9 11 7 9 11 2
21 1 0 9 1 11 13 2 16 9 9 11 13 14 3 1 12 7 12 9 11 2
3 9 0 9
2 0 9
22 13 15 13 1 9 2 1 15 15 1 0 9 11 11 3 13 1 0 3 9 12 2
6 3 13 13 9 0 2
22 7 15 15 3 13 1 10 9 2 15 10 9 13 1 9 9 2 0 1 0 9 2
22 7 4 3 13 9 15 2 15 1 9 13 0 2 7 4 3 13 7 10 0 9 2
25 1 9 9 12 4 1 10 9 13 15 3 1 9 12 2 3 3 1 10 9 0 0 9 13 2
14 13 4 1 15 7 1 9 2 3 3 1 9 12 2
22 3 15 3 10 9 2 0 1 0 9 10 0 9 2 13 13 0 9 1 0 9 2
23 3 3 2 3 9 3 0 1 9 0 7 0 9 0 9 2 15 9 9 12 3 13 2
50 1 9 9 13 10 2 0 2 9 2 2 9 13 13 0 9 2 13 3 1 15 9 0 2 15 3 13 9 1 9 9 7 0 9 2 16 7 0 9 2 16 3 13 9 0 7 0 9 2 2
8 9 7 9 0 9 13 4 2
11 2 2 3 13 0 3 13 9 9 2 2
25 0 9 7 13 0 9 2 1 0 9 2 16 13 9 1 0 9 7 1 0 7 0 9 2 2
27 2 2 1 10 9 13 9 1 0 9 7 3 0 9 10 9 13 2 7 15 15 3 13 9 9 2 2
17 3 15 13 0 9 13 12 9 2 15 13 0 1 9 9 9 2
14 15 0 1 9 2 13 4 3 1 0 9 0 9 2
29 7 15 13 1 9 9 12 1 9 12 12 9 11 2 15 15 3 13 1 0 7 3 3 15 1 0 7 11 2
40 3 15 15 1 9 13 0 7 0 9 2 15 15 7 3 13 2 0 9 2 2 1 15 4 1 2 9 9 1 9 9 14 1 0 9 3 13 9 2 2
28 1 0 13 0 2 16 9 0 9 13 9 7 9 9 12 3 3 2 7 13 7 10 9 15 15 3 13 2
33 16 3 3 4 10 9 2 9 2 1 9 3 0 13 10 9 2 13 1 9 2 16 0 0 9 11 12 1 15 13 15 0 2
29 3 4 3 13 3 0 16 11 2 16 4 1 10 9 13 15 0 13 2 7 9 13 9 2 15 15 13 13 2
32 9 0 9 1 9 0 9 11 11 13 12 1 9 9 0 0 9 0 9 2 15 15 1 0 9 13 1 0 11 1 11 2
15 9 13 7 13 0 9 2 13 9 7 13 0 9 9 2
4 9 15 13 9
2 11 2
29 9 1 9 1 9 0 0 9 1 0 9 3 13 3 1 0 9 11 2 11 1 11 9 9 1 12 0 9 2
8 1 9 13 3 0 9 12 2
17 10 9 13 13 16 0 9 11 2 11 1 9 1 9 7 9 2
26 0 9 9 9 9 4 1 9 9 9 11 13 1 9 13 3 0 9 1 0 9 2 9 7 9 2
10 0 9 15 1 9 9 13 2 13 11
2 11 2
21 9 9 9 9 11 11 13 13 2 16 2 0 9 15 1 9 9 13 13 2 2
10 13 15 1 9 1 9 3 9 11 2
18 2 13 1 15 2 16 0 9 9 11 13 0 2 2 13 3 11 2
19 9 1 9 9 1 0 9 7 13 2 13 7 0 9 1 9 0 9 2
26 9 9 11 11 3 11 13 2 16 9 9 9 4 13 14 3 2 16 15 13 1 9 10 0 9 2
15 1 0 9 13 1 11 14 12 9 2 9 9 13 12 2
13 9 0 12 13 9 11 13 1 2 0 9 2 2
8 3 15 13 12 0 9 9 2
21 0 2 9 2 1 9 9 13 3 16 12 9 2 13 0 9 7 13 0 9 2
28 1 9 9 13 9 1 15 2 16 9 13 0 9 2 9 0 9 13 1 0 9 7 13 9 1 9 9 2
24 9 0 0 9 11 11 15 13 1 0 11 1 9 9 11 1 9 10 9 11 11 7 11 11
5 9 13 9 1 9
2 11 2
30 1 0 9 12 2 12 1 11 15 3 13 0 9 11 11 2 15 1 0 0 9 1 9 13 13 9 1 9 14 2
14 2 13 15 9 1 9 2 0 9 9 13 1 15 2
14 16 4 13 9 2 7 13 2 3 15 15 15 13 2
15 13 4 0 9 16 1 12 9 2 3 4 3 13 3 2
9 13 4 1 9 7 9 15 13 2
43 13 4 15 2 16 13 9 2 7 16 15 1 15 13 2 16 15 15 4 13 13 1 9 2 2 13 11 11 7 3 13 2 16 10 9 3 13 0 9 1 0 9 2
7 2 13 4 15 13 3 2
20 1 9 1 15 13 11 11 2 13 15 12 9 7 9 11 7 13 0 9 2
7 3 4 15 13 3 3 2
21 1 9 4 15 13 9 1 11 2 13 11 7 11 7 0 9 13 3 3 2 2
10 0 13 1 9 2 14 16 13 1 11
4 11 2 11 2
24 14 0 9 1 15 9 2 15 13 1 9 1 0 9 0 9 1 9 14 2 13 9 11 2
13 1 0 12 0 9 15 13 12 9 1 9 9 2
21 1 9 13 12 2 12 1 11 7 9 15 13 7 0 9 12 2 12 1 11 2
23 14 1 15 2 16 11 13 1 11 7 11 13 1 11 14 9 2 13 7 3 1 9 2
20 2 1 12 9 1 9 2 15 4 13 13 3 2 4 13 1 9 12 9 2
7 15 3 15 15 14 13 2
41 1 9 13 1 11 7 9 13 3 0 2 9 1 9 14 13 14 1 9 2 2 13 0 9 9 7 9 11 11 2 15 13 1 9 10 9 1 11 3 0 2
18 2 1 0 12 12 13 11 3 0 7 15 4 15 13 13 1 9 2
16 1 0 9 3 15 13 0 2 7 13 4 15 10 9 2 2
19 0 9 1 9 14 13 3 7 0 11 2 15 13 12 2 12 1 11 2
28 1 9 9 2 11 2 11 2 11 2 13 3 0 9 2 7 1 9 9 1 9 14 13 13 3 12 9 2
12 0 9 9 2 15 13 1 9 1 9 14 2
12 12 2 9 2 11 2 11 2 11 2 11 2
5 11 13 14 1 9
15 0 9 7 0 9 0 9 13 1 0 9 9 0 11 2
16 1 3 0 9 9 13 9 14 1 0 0 2 3 0 9 2
15 9 7 0 9 13 13 7 0 9 11 11 7 11 11 2
22 2 13 3 3 0 9 1 15 2 16 4 15 1 9 13 7 13 13 10 0 9 2
17 7 1 15 0 9 13 0 9 1 11 2 3 4 13 3 3 2
35 3 13 9 0 9 7 9 15 3 13 2 2 13 11 7 11 15 13 2 2 10 0 9 4 3 13 7 0 9 2 16 15 11 13 2
19 3 15 1 10 9 3 13 0 11 11 2 15 13 3 9 1 9 13 2
11 13 15 7 15 15 15 13 1 9 2 2
10 3 15 13 7 9 13 9 9 9 2
9 2 1 9 13 3 3 0 9 2
21 11 11 13 3 0 9 2 16 0 11 11 2 1 15 13 3 0 9 3 0 2
12 7 0 9 4 13 1 9 2 2 13 11 2
22 0 9 9 9 3 0 9 13 2 7 16 13 2 16 3 10 9 1 9 9 13 2
15 2 3 14 13 9 7 13 1 15 9 2 2 13 11 2
8 9 11 13 11 1 0 2 11
33 0 0 9 1 9 0 11 15 3 13 0 0 9 11 11 2 12 9 2 2 15 1 0 9 13 1 9 0 11 11 1 11 2
39 1 9 13 1 9 12 2 1 12 9 15 1 0 9 13 1 11 9 11 2 3 4 1 9 12 13 1 11 7 3 3 1 9 16 0 9 13 11 2
8 9 9 7 13 1 0 9 2
42 1 11 13 14 12 9 1 11 1 9 11 11 2 15 3 13 1 0 2 11 7 16 15 3 13 2 0 4 1 10 9 3 13 11 2 15 13 3 0 9 11 2
9 10 9 11 3 13 1 9 9 2
3 0 0 9
3 0 11 2
26 0 9 11 11 13 10 0 9 10 9 11 7 13 15 1 9 9 11 2 11 2 12 2 12 2 2
38 0 12 13 3 0 2 13 1 15 12 9 2 16 0 9 13 3 11 2 15 13 9 0 12 9 3 2 16 11 1 11 13 9 1 12 2 12 2
14 1 0 9 0 9 13 7 11 11 7 13 12 9 2
12 1 11 13 11 9 0 11 11 12 2 12 2
25 1 9 12 2 12 1 0 12 13 0 9 11 2 16 9 1 10 9 13 1 9 1 0 9 2
10 1 0 9 9 12 2 12 13 11 2
1 9
28 11 2 11 2 12 2 12 2 2 11 11 2 9 11 2 2 1 0 9 12 12 9 13 9 9 14 0 2
8 9 11 13 1 15 0 2 2
27 11 11 2 9 11 2 2 3 13 1 9 11 7 11 7 3 15 4 13 1 0 9 1 9 14 2 2
46 11 2 11 2 12 2 12 2 2 11 11 2 9 11 2 2 11 1 0 9 13 1 0 12 3 2 7 3 4 15 13 1 10 9 2 16 15 13 2 16 4 3 9 13 2 2
22 11 11 2 9 11 2 2 13 4 10 9 2 0 14 2 16 15 13 16 0 9 2
11 1 9 12 2 12 4 3 13 9 2 2
12 9 11 15 1 0 9 11 7 11 2 11 13
6 1 9 1 12 9 2
8 11 11 15 13 13 1 0 9
2 11 2
13 1 0 9 13 9 11 11 1 0 9 0 9 2
22 1 9 13 1 0 9 2 9 11 11 7 13 2 16 13 0 1 9 1 0 9 2
12 2 9 1 0 9 13 7 13 3 1 9 2
18 16 4 13 2 10 4 13 13 1 9 9 2 3 15 13 0 9 2
9 9 13 7 0 2 2 13 11 2
20 0 0 9 1 0 9 13 9 11 2 15 15 13 1 3 0 9 1 11 2
16 9 0 9 15 1 9 0 9 1 0 11 13 1 0 9 2
14 1 3 0 9 1 11 13 2 7 13 9 0 9 2
17 1 9 13 11 12 9 1 9 12 9 2 12 9 7 12 9 2
27 1 0 9 1 11 13 9 1 9 0 9 11 2 9 2 2 11 2 9 2 7 11 2 0 9 2 2
25 0 9 11 2 12 2 9 2 12 9 2 12 9 2 12 9 2 9 12 2 12 2 12 9 2
22 13 2 11 2 11 11 2 2 11 2 1 9 2 2 11 2 1 9 1 11 2 2
28 13 2 11 2 11 2 11 2 12 9 1 11 2 2 11 2 11 2 11 2 7 11 2 11 2 9 2 2
2 9 9
2 11 2
24 9 0 0 1 9 0 9 15 3 13 0 9 11 11 2 15 13 1 0 0 9 11 11 2
9 0 0 9 13 1 9 10 9 2
5 9 1 9 1 11
2 11 2
21 9 0 9 12 1 9 1 9 1 11 15 1 9 7 1 9 13 12 9 11 2
31 1 0 9 9 2 12 13 1 12 0 9 1 9 1 9 0 9 9 1 10 9 11 2 11 2 11 2 11 7 11 2
18 11 2 15 15 3 13 1 0 9 2 4 3 13 1 0 9 9 2
29 2 11 13 1 15 0 2 16 3 15 13 2 15 4 0 9 13 1 9 1 0 11 2 2 13 9 11 11 2
1 3
21 0 9 11 13 13 9 12 2 9 9 1 11 1 11 11 1 0 9 0 9 2
11 3 13 2 16 15 13 1 11 9 9 2
4 9 13 1 9
9 0 9 11 11 4 13 13 9 9
2 11 2
18 0 9 0 0 9 2 11 2 15 3 13 1 0 9 1 0 9 2
23 1 9 9 1 0 9 13 9 0 9 1 11 1 0 9 0 9 1 9 1 0 9 2
54 2 11 15 13 16 9 9 2 15 15 13 10 9 3 1 9 12 2 7 1 10 0 9 13 10 9 2 2 13 9 11 11 0 7 1 9 9 1 9 0 9 13 2 2 10 9 13 13 9 3 1 15 9 2
18 9 13 16 9 2 7 1 0 9 4 1 0 9 13 0 9 2 2
23 15 9 11 13 1 9 0 0 2 9 2 13 0 9 1 11 7 11 7 13 0 9 2
24 0 9 11 11 3 13 9 1 9 10 9 7 3 13 1 9 9 9 2 9 7 0 9 2
14 1 0 9 2 9 7 0 9 13 0 9 11 11 2
19 11 11 2 9 9 2 12 2 1 9 0 9 13 1 0 7 0 9 2
24 0 9 1 0 9 15 4 13 11 11 2 1 9 3 11 11 1 11 7 11 11 1 11 2
15 11 11 13 1 9 0 9 7 9 9 11 1 0 9 2
10 1 0 9 7 0 9 13 11 11 2
23 11 11 15 4 13 9 9 1 9 7 11 11 4 3 16 1 0 0 9 13 1 9 2
10 0 9 11 3 13 0 9 10 9 2
17 3 9 0 2 9 7 9 13 2 16 4 13 9 0 9 9 2
34 1 9 9 7 9 9 13 13 0 9 11 2 7 14 3 0 9 1 9 0 9 1 0 0 9 2 11 11 16 9 9 11 11 2
26 1 9 2 1 9 9 3 0 9 13 0 0 9 11 11 0 2 0 9 13 0 0 9 11 11 2
28 9 9 9 1 11 15 4 1 0 9 13 12 2 9 1 11 1 11 2 9 15 13 1 9 3 1 11 2
24 1 11 4 12 2 7 12 2 9 13 9 7 9 1 11 1 15 2 16 9 4 13 3 2
16 1 0 9 4 11 13 9 11 1 12 9 2 9 7 9 2
18 9 9 0 9 15 0 9 9 13 2 13 12 0 9 1 12 9 2
8 13 15 7 1 9 9 9 2
14 0 9 11 11 9 13 10 9 2 7 11 15 13 2
17 2 13 9 2 15 4 13 10 9 13 2 2 13 9 0 9 2
18 11 13 2 16 13 9 1 10 9 1 9 2 7 13 1 10 9 2
29 2 13 0 0 9 13 2 2 13 0 9 2 15 13 13 9 0 9 1 9 9 9 7 9 0 0 9 11 2
4 9 9 3 9
2 11 2
20 3 3 1 15 13 9 1 9 9 9 2 9 1 0 9 9 9 0 11 2
17 1 11 11 2 12 2 7 11 11 2 12 2 13 9 11 11 2
8 2 3 13 2 15 15 13 2
12 15 4 13 3 0 2 2 13 0 0 9 2
15 9 9 12 4 1 9 0 9 13 11 11 1 11 11 2
19 7 15 7 13 9 1 9 11 11 2 16 4 10 9 13 1 0 9 2
6 9 13 0 0 9 2
28 11 11 2 1 9 2 15 1 12 2 9 1 9 1 9 1 9 13 1 11 11 12 2 12 2 12 2 12
5 0 15 1 11 13
2 11 2
37 1 9 9 15 1 9 9 0 11 11 11 3 13 9 13 9 9 0 0 9 1 9 9 0 9 2 15 13 13 9 0 0 9 11 1 11 2
45 1 12 9 15 1 9 9 11 13 13 9 11 2 11 2 11 2 1 9 11 2 11 2 11 7 0 2 1 9 0 13 9 11 1 9 11 2 11 2 11 2 11 7 9 2
33 9 12 9 2 15 3 13 0 9 1 9 2 13 9 1 9 0 9 1 0 9 1 0 9 11 2 2 15 7 1 9 13 2
14 2 13 0 9 7 15 13 1 9 1 9 1 11 2
20 9 15 13 7 0 9 1 0 9 2 2 13 3 3 3 9 11 11 0 2
21 3 7 13 10 0 9 0 9 9 11 11 2 16 4 13 0 9 9 1 9 2
20 1 9 0 9 7 1 9 3 13 9 2 16 0 9 13 2 15 13 0 2
17 9 9 1 11 9 3 0 9 9 13 1 10 9 9 0 9 2
3 1 0 9
16 0 9 11 11 13 9 1 11 11 1 12 2 12 2 12 2
15 11 13 1 11 1 9 12 1 12 9 9 1 11 11 2
4 11 13 1 9
2 11 2
12 0 9 1 0 0 9 11 11 13 3 9 2
13 9 3 13 0 9 1 9 1 9 12 12 9 2
15 2 13 9 2 16 4 15 13 13 9 1 9 0 9 2
29 15 13 1 9 2 3 15 13 13 12 12 1 9 2 15 13 1 9 13 2 2 13 11 9 0 9 11 11 2
20 0 9 13 1 11 9 1 11 2 16 4 9 1 9 13 9 1 9 11 2
26 9 9 13 3 2 7 9 0 9 11 1 0 9 1 9 11 11 2 15 13 9 0 9 11 11 2
27 15 13 0 9 9 9 0 9 2 15 1 0 0 9 3 13 9 7 13 9 9 0 9 1 0 9 2
25 1 9 1 9 9 13 9 9 11 2 1 9 11 15 3 12 9 9 13 1 9 1 0 11 2
6 0 9 0 9 9 9
2 11 2
11 1 9 1 0 9 13 9 0 9 9 2
26 9 13 9 9 1 11 1 9 9 1 0 9 2 0 9 4 13 0 0 9 9 1 11 0 11 2
33 1 0 9 9 1 15 13 13 9 1 0 9 2 0 11 2 15 15 1 0 9 13 3 16 12 12 9 1 12 9 1 11 2
5 9 1 11 0 9
2 11 2
39 9 9 0 9 11 11 1 0 9 2 11 11 11 2 12 2 9 11 2 7 0 11 0 9 11 11 2 12 2 2 2 15 13 13 9 0 0 11 2
20 13 15 0 9 9 0 9 12 9 2 15 15 0 9 13 1 9 9 11 2
16 9 0 9 13 12 9 2 16 0 9 1 9 13 12 9 2
17 0 9 13 11 11 2 12 2 2 2 9 0 2 12 2 2 2
23 10 9 13 11 11 2 9 15 13 15 2 16 10 9 15 13 0 9 11 2 11 13 2
4 11 13 9 11
2 11 2
25 9 1 15 2 16 13 9 9 0 0 9 2 15 0 9 11 11 11 13 14 1 0 0 9 2
30 13 15 7 3 1 0 9 0 9 11 2 16 13 13 9 2 16 16 9 9 0 9 4 1 9 9 13 1 9 2
26 2 13 15 0 9 2 9 9 4 13 16 9 1 9 9 2 7 13 2 16 15 3 0 14 13 2
24 1 9 7 13 9 9 9 7 4 13 9 9 9 9 11 2 0 9 11 2 2 13 11 2
19 10 9 13 7 3 1 0 9 1 11 2 16 1 9 9 1 0 9 2
5 9 13 1 0 9
3 11 11 2
28 9 1 9 9 7 9 1 0 0 9 11 15 13 1 12 0 9 11 7 11 0 2 1 15 0 9 13 2
20 1 10 9 13 1 9 9 2 7 1 0 9 11 15 12 9 13 1 11 2
20 11 13 1 9 0 11 1 9 12 2 12 2 11 1 9 12 1 9 12 2
2 9 9
2 11 2
29 0 9 13 9 9 11 11 11 11 2 15 4 13 1 9 1 9 9 11 11 11 1 9 12 9 12 2 9 2
23 0 9 0 0 9 13 1 0 11 9 11 11 9 7 12 9 1 11 11 2 3 2 2
3 11 7 11
1 9
2 9 2
29 0 0 9 9 11 11 4 13 13 7 3 2 1 12 1 12 0 9 11 2 11 2 11 2 15 13 9 9 2
9 1 9 4 3 15 13 7 13 2
38 3 2 16 15 3 11 13 1 10 0 9 2 15 13 0 7 0 9 2 16 1 11 13 9 3 3 10 9 13 7 16 9 10 9 13 1 9 2
9 13 2 16 0 9 13 10 9 2
18 16 13 1 9 2 16 0 9 9 13 3 0 2 9 13 3 0 2
31 3 0 9 13 3 0 7 13 4 3 0 9 16 3 9 11 1 9 9 2 11 7 11 2 0 1 0 7 0 9 2
17 15 3 15 13 1 10 0 9 2 0 1 0 9 1 9 3 2
16 0 9 2 9 7 9 1 15 13 13 13 1 0 0 9 2
9 12 1 0 7 0 13 13 3 2
33 11 11 15 1 10 12 9 13 13 3 0 9 2 15 15 1 3 0 9 2 3 1 10 0 9 2 3 2 13 2 10 9 2
40 3 3 13 9 3 13 2 13 2 14 0 9 7 0 9 2 2 13 1 15 0 9 0 9 1 9 0 9 9 7 0 2 3 16 0 9 9 2 9 2
22 3 3 13 0 0 9 2 7 13 3 7 3 13 0 9 1 0 9 1 0 9 2
30 15 13 2 10 9 13 3 1 15 2 7 3 1 0 9 2 7 10 0 9 2 13 2 3 0 9 11 11 13 2
28 0 9 1 0 0 0 9 3 3 13 2 3 16 1 0 0 9 11 11 2 0 0 9 2 0 11 11 2
9 11 11 11 11 2 13 7 3 2
6 2 9 1 9 2 2
7 9 13 2 11 2 12 2
2 9 9
1 9
33 10 0 9 2 15 13 1 0 0 9 7 3 15 3 13 2 13 1 0 0 9 0 0 9 7 1 9 1 15 7 0 9 2
22 0 1 15 13 9 2 13 15 3 7 0 9 2 10 9 3 13 2 0 2 9 2
17 13 1 15 3 9 9 0 11 7 9 11 2 3 13 0 9 2
27 1 3 0 9 13 3 0 9 2 1 15 13 7 11 11 2 12 2 2 9 0 1 0 9 7 9 2
7 13 3 0 7 3 0 2
25 10 9 2 1 15 3 13 13 1 0 9 9 2 13 0 9 2 9 2 9 2 9 7 9 2
11 1 0 9 13 1 0 9 1 9 0 2
26 3 13 0 9 0 7 0 2 1 0 9 2 13 9 2 15 15 13 2 9 2 9 2 0 9 2
14 13 15 9 2 9 2 9 2 9 2 0 0 9 2
16 16 4 15 13 0 9 13 2 13 4 11 16 10 0 9 2
11 13 0 1 0 2 13 0 7 0 9 2
16 14 9 0 9 2 1 15 15 9 13 2 15 13 3 0 2
16 16 4 13 3 0 14 12 2 0 9 2 3 3 15 0 2
7 11 13 13 1 10 9 2
13 3 14 1 0 0 9 1 9 13 9 15 15 2
23 3 7 13 10 9 2 15 16 4 13 1 15 2 0 9 10 9 4 13 3 0 9 2
17 9 13 1 9 0 9 2 1 15 4 15 7 3 3 3 13 2
15 3 13 3 9 9 2 3 16 3 0 11 11 1 11 2
38 16 4 11 13 0 9 0 7 0 2 1 10 9 13 10 9 1 0 9 13 2 2 13 4 1 15 13 9 2 9 2 15 15 3 13 1 9 2
6 9 1 9 1 0 9
26 0 0 9 11 11 7 11 11 2 12 2 15 13 1 11 16 9 0 2 0 0 9 9 1 9 2
19 9 13 0 0 9 0 0 9 11 7 0 0 9 11 12 7 0 11 2
10 10 9 15 13 3 1 0 9 11 2
15 11 11 13 1 11 2 3 13 0 9 2 9 9 2 2
22 1 0 9 13 1 11 2 3 13 1 9 1 0 11 2 1 11 15 3 13 3 2
13 9 1 9 13 2 3 13 2 10 9 10 9 2
26 13 9 0 11 2 15 13 9 1 0 9 11 0 9 2 1 9 2 15 2 13 9 7 9 2 2
20 9 0 9 3 13 9 2 9 7 0 9 1 9 2 0 7 10 0 9 2
11 13 0 0 9 9 9 0 9 2 2 2
14 2 9 10 9 4 1 15 13 3 2 2 13 9 2
19 10 9 4 1 12 9 3 13 9 0 11 2 15 3 13 10 12 9 2
9 3 13 9 7 0 9 11 12 2
15 15 7 1 9 13 2 1 9 13 0 13 3 9 9 2
21 15 15 3 13 1 9 0 9 11 2 15 1 9 9 13 1 12 12 9 9 2
16 10 3 0 9 13 9 11 15 2 16 15 15 9 3 13 2
17 3 15 1 15 13 1 9 2 3 15 13 13 1 0 0 9 2
31 9 15 13 1 12 9 1 11 7 9 7 10 0 9 13 0 0 9 2 11 11 2 11 11 2 11 11 7 11 11 2
24 2 0 9 15 15 14 13 13 14 1 0 9 2 16 15 10 9 3 13 2 2 13 11 2
29 2 13 2 16 7 1 9 13 9 2 1 15 15 10 0 9 2 16 13 3 0 2 13 13 2 2 13 9 2
14 9 1 9 13 1 10 9 1 0 9 1 0 9 2
13 2 13 2 16 9 4 9 13 2 2 13 9 2
16 2 9 2 15 13 10 9 0 13 2 3 13 0 9 13 2
22 13 2 16 9 15 13 3 2 16 15 13 1 9 7 13 15 15 13 7 13 2 2
12 1 9 9 1 0 0 9 15 3 13 9 2
15 15 7 0 9 2 15 7 1 0 9 10 0 9 13 2
13 1 11 4 13 9 0 1 9 9 13 0 9 2
16 2 13 15 1 9 2 9 9 7 0 9 2 2 13 9 2
1 3
32 0 9 0 9 11 11 2 12 2 12 2 13 10 0 9 0 1 9 2 16 9 13 1 15 2 16 9 13 4 3 13 2
23 9 11 1 11 15 3 13 13 2 16 4 11 2 12 2 13 3 1 9 16 1 9 2
5 15 2 3 2 3
16 9 9 1 11 13 3 9 0 0 9 0 9 12 2 9 2
17 0 1 9 11 0 13 3 2 12 2 1 0 9 9 11 11 2
26 9 0 9 1 9 1 11 11 7 11 11 15 13 3 2 12 2 1 9 11 11 1 0 9 9 2
11 9 1 9 12 13 1 9 12 7 9 9
20 12 9 9 0 9 13 1 0 9 9 9 9 9 0 2 0 7 0 9 2
22 0 9 1 10 9 13 3 12 9 9 2 9 9 13 1 9 9 2 9 7 9 2
20 1 9 9 11 11 13 0 9 1 9 9 1 9 0 7 0 9 0 9 2
18 0 9 13 3 0 0 9 2 15 13 2 9 0 9 1 9 2 2
25 0 9 9 1 0 9 13 1 11 12 9 2 16 4 2 13 9 10 0 9 9 7 9 2 2
26 1 9 0 4 3 13 12 9 9 1 9 9 1 9 12 7 12 9 9 1 9 9 9 7 9 2
31 0 9 11 0 12 2 7 11 13 1 12 9 2 9 0 9 12 12 9 2 9 3 0 9 7 9 9 9 9 9 2
7 9 0 13 9 0 9 2
43 2 16 1 0 9 13 9 1 12 9 0 16 3 2 13 4 13 3 12 9 2 2 13 11 2 15 13 1 0 0 9 0 9 2 15 4 13 13 9 1 0 9 2
4 9 9 1 9
1 9
2 9 2
21 0 0 9 9 9 3 13 1 9 9 11 11 2 9 11 11 7 9 11 11 2
9 3 9 9 7 9 13 0 9 2
12 13 7 0 9 2 15 13 9 12 0 9 2
19 1 9 9 13 15 12 9 1 0 0 9 11 9 0 11 1 11 11 2
23 13 0 0 9 9 7 9 9 2 15 3 13 1 9 0 0 9 10 9 0 0 9 2
11 9 1 0 9 9 15 13 3 16 0 2
15 0 0 9 9 13 9 0 1 9 7 9 1 11 11 2
24 12 1 10 3 0 0 9 13 11 11 7 11 11 3 2 7 3 13 9 2 3 3 3 2
14 3 13 9 9 9 2 10 9 2 9 9 7 9 2
18 0 9 0 9 15 13 0 9 6 2 9 15 9 0 9 11 11 2
19 9 13 2 16 10 9 13 15 3 0 10 0 9 2 0 9 7 9 2
15 1 11 7 11 15 13 0 0 9 1 9 9 7 9 2
15 0 0 9 11 11 13 0 9 1 0 9 9 7 9 2
21 0 0 12 9 1 9 2 9 7 9 13 9 2 7 9 1 0 0 9 9 2
15 0 2 0 9 0 0 9 13 0 9 1 3 0 9 2
12 9 14 2 16 9 13 1 3 0 0 9 2
9 0 9 9 9 11 11 3 13 2
19 11 11 12 2 0 9 9 9 3 2 11 11 2 11 11 2 11 11 2
9 0 9 11 2 12 2 9 12 2
31 9 0 9 9 9 2 9 1 0 9 2 1 9 9 9 11 11 1 9 9 11 7 9 11 13 1 0 9 9 9 2
38 11 11 1 0 9 13 0 9 3 15 2 16 1 15 13 9 2 0 9 15 13 1 0 9 2 7 16 13 1 15 3 3 9 2 9 7 9 2
12 3 7 9 4 1 15 13 16 3 0 9 2
23 1 0 9 11 11 9 13 1 0 11 11 16 9 2 3 2 7 11 11 1 9 9 2
9 11 11 1 11 3 13 9 0 9
29 9 0 9 11 11 3 13 12 2 9 1 0 9 11 9 9 11 11 9 1 9 2 0 1 0 9 11 11 2
21 0 9 1 10 0 9 15 13 1 12 12 9 2 9 9 13 12 9 9 2 2
18 11 15 15 13 13 9 9 9 2 15 13 13 9 0 9 1 11 2
50 0 11 11 2 0 9 13 0 3 1 9 0 9 2 0 9 2 13 12 2 9 7 9 0 9 2 4 1 11 1 9 9 14 1 12 2 9 13 9 0 9 9 11 1 11 1 9 9 0 2
19 12 1 10 9 4 13 13 7 11 11 2 0 3 1 0 9 0 9 2
17 9 13 13 1 11 2 1 11 7 3 1 9 1 9 0 11 2
1 3
21 1 9 0 9 9 11 11 15 4 13 0 9 13 1 0 11 3 1 9 12 2
46 1 1 15 2 16 9 1 11 13 10 0 9 1 9 11 2 7 13 9 9 0 9 1 11 13 2 13 9 7 13 2 16 1 0 9 11 4 13 2 1 0 9 2 1 11 2
33 9 9 0 9 2 0 1 0 9 0 0 9 2 13 1 11 9 9 2 15 13 9 11 13 1 0 0 9 0 9 1 9 2
23 0 9 11 11 11 13 9 2 16 4 1 9 9 10 9 1 0 9 0 9 11 13 2
32 11 3 13 10 9 2 7 13 2 16 15 13 9 9 0 0 9 1 9 12 2 1 15 13 9 1 0 9 1 9 11 2
10 0 9 9 1 15 3 10 9 13 2
9 0 9 1 0 9 13 3 13 2
20 1 9 0 9 0 11 15 1 15 1 3 16 12 0 9 13 12 9 9 2
4 0 9 1 11
4 0 9 13 9
4 11 2 11 2
26 11 15 13 1 9 9 2 16 0 9 13 0 9 2 13 0 9 9 11 11 1 9 1 9 11 2
27 13 2 16 9 9 11 11 13 13 15 0 2 16 13 10 9 7 9 2 16 4 15 13 1 9 9 2
30 11 2 0 11 7 11 3 13 0 0 9 1 0 11 2 1 15 0 9 13 0 9 11 11 0 9 9 11 11 2
6 13 15 0 9 9 2
34 10 0 9 2 1 10 9 15 13 0 12 9 0 9 2 11 7 11 2 14 13 1 9 0 9 0 0 9 7 1 10 0 9 2
28 9 3 3 3 13 2 16 4 15 0 2 0 9 1 11 13 13 1 11 7 0 11 1 0 2 0 11 2
5 11 13 9 9 11
2 11 2
20 0 9 9 11 11 13 0 9 0 9 2 16 4 13 1 11 12 0 9 2
25 16 13 9 0 11 2 15 0 9 1 12 9 0 9 11 1 11 3 13 1 0 9 0 9 2
28 1 10 9 0 9 13 2 16 13 1 9 0 0 0 9 2 11 2 2 15 15 13 13 10 9 0 9 2
24 16 13 9 11 2 9 0 9 1 9 13 2 16 0 9 1 9 0 9 3 13 0 9 2
5 11 2 9 9 13
2 11 2
21 0 9 1 9 1 0 9 13 0 9 0 9 2 15 15 13 13 1 10 9 2
33 9 3 13 1 0 9 9 0 9 2 1 9 13 7 0 9 1 9 13 9 2 15 13 13 10 9 2 9 9 0 9 9 2
13 13 15 3 1 9 0 9 2 9 7 0 9 2
15 16 15 10 9 13 2 9 13 13 9 14 1 12 9 2
24 9 0 9 11 11 11 15 1 0 9 13 1 10 9 2 16 2 13 9 0 9 9 2 2
5 11 13 9 1 11
2 11 2
27 11 15 3 1 9 10 9 0 2 11 0 13 1 9 9 11 11 2 9 0 9 0 11 1 0 11 2
18 9 11 13 1 0 9 1 9 16 0 9 9 9 1 0 9 11 2
26 1 0 9 1 9 1 0 11 9 13 2 16 2 14 12 9 9 1 9 9 13 9 0 1 9 2
14 11 7 9 15 7 13 1 9 9 7 10 9 2 2
18 0 9 1 0 11 2 1 15 13 10 9 2 3 3 13 0 9 2
22 11 13 1 2 9 2 7 13 15 0 9 1 0 0 9 1 0 9 2 11 2 2
9 9 13 2 16 4 13 9 9 2
6 11 1 9 9 1 11
28 0 9 11 3 1 10 0 9 13 1 9 13 9 1 11 2 3 15 7 13 1 7 13 15 13 1 9 2
28 3 1 9 0 9 7 11 13 13 0 0 9 2 16 4 13 9 2 16 13 15 11 2 15 13 0 9 2
19 1 9 15 15 13 13 9 0 0 9 1 0 9 1 9 9 0 9 2
42 11 13 3 13 10 9 1 0 9 2 9 0 9 2 11 2 11 7 11 2 16 4 3 13 0 9 7 13 1 9 0 2 0 9 1 9 12 1 9 0 9 2
29 1 9 0 9 11 11 11 15 3 13 9 0 9 1 0 0 9 2 1 10 9 13 0 9 9 11 11 11 2
12 10 9 3 13 9 0 9 2 0 9 2 2
13 9 15 13 1 0 9 7 1 0 13 9 11 2
28 2 13 15 0 0 9 1 10 0 9 2 2 13 11 2 15 13 1 12 9 1 9 0 9 1 9 12 2
15 1 0 2 0 9 1 0 9 4 3 1 11 13 9 2
34 11 13 9 1 0 9 2 16 4 1 9 7 9 9 13 9 12 0 9 7 12 0 9 2 1 15 9 4 13 9 1 0 9 2
11 9 12 9 13 0 9 1 2 0 2 2
9 3 1 11 13 10 2 9 2 2
13 9 3 13 1 0 9 9 9 7 0 9 11 11
4 11 14 13 9
2 11 2
16 0 9 9 7 0 9 11 11 13 1 9 9 11 10 9 2
12 11 0 9 1 9 13 2 7 3 14 3 2
17 13 15 3 0 0 9 0 11 0 2 15 9 13 3 3 0 2
24 11 2 15 13 1 0 9 0 9 1 0 9 2 15 1 9 13 9 9 13 0 0 9 2
35 1 9 3 9 13 10 0 9 1 9 9 0 9 11 2 11 2 15 15 3 13 10 3 0 0 9 2 7 3 13 9 9 1 0 2
36 2 11 2 11 2 13 3 1 9 16 1 0 9 2 2 13 9 1 9 1 0 9 2 16 1 9 0 0 9 13 15 1 9 9 9 2
24 11 15 3 13 9 0 9 11 11 2 16 13 3 0 2 16 15 4 15 13 1 0 9 2
27 9 13 0 1 9 9 7 15 2 16 15 1 11 11 2 15 1 9 9 13 2 13 3 0 0 9 2
5 11 15 13 13 9
2 11 2
25 0 9 15 1 9 1 9 13 1 9 7 1 9 13 0 9 11 2 7 0 9 10 9 13 2
19 13 15 0 9 11 2 11 1 9 1 9 1 9 0 9 1 0 11 2
38 9 0 9 1 11 3 13 9 13 9 1 9 9 11 11 2 7 3 1 9 2 16 0 9 3 13 3 3 0 0 9 2 1 0 1 9 11 2
5 9 11 1 9 11
4 11 2 11 2
31 9 14 12 0 9 13 1 9 1 9 9 1 9 9 11 2 10 9 13 13 12 9 11 2 15 1 10 0 9 13 2
17 9 0 9 4 13 9 2 15 13 0 9 1 9 1 0 9 2
34 1 0 9 1 12 9 13 1 9 2 3 1 9 9 13 0 9 9 2 15 13 13 1 9 0 9 0 1 11 7 11 0 9 2
4 9 9 9 2
18 9 9 0 9 13 1 0 9 12 9 1 12 9 9 7 12 9 2
36 3 3 13 9 11 11 11 2 13 15 9 0 9 9 11 2 11 2 15 7 1 0 9 9 1 10 9 13 1 0 9 0 9 1 11 2
22 11 3 13 10 9 1 0 9 2 15 9 4 13 1 0 9 13 0 9 0 9 2
20 11 3 3 13 2 16 9 13 9 9 0 9 11 11 11 1 9 1 9 2
10 1 15 13 7 9 0 9 7 9 2
27 9 13 0 11 13 14 3 2 16 15 9 13 9 0 9 2 15 4 15 1 0 9 13 13 11 11 2
5 11 0 1 0 9
2 11 2
24 9 9 0 11 1 0 11 1 9 9 11 11 13 1 10 9 11 11 1 2 0 9 2 2
36 1 9 1 0 9 0 11 13 11 0 0 9 1 0 2 0 9 1 2 9 3 2 1 9 1 0 9 1 9 12 7 1 0 0 9 2
26 11 13 2 16 15 0 11 13 1 9 0 9 9 2 7 3 13 9 1 2 0 9 0 9 2 2
22 13 1 15 0 2 1 10 2 9 2 11 13 9 0 9 2 16 3 13 9 11 2
5 11 1 9 1 11
2 11 2
35 1 0 9 0 7 0 11 7 1 9 0 9 11 2 9 2 1 11 13 1 9 1 11 1 0 9 9 11 11 0 9 9 11 11 2
13 0 9 15 3 13 1 0 9 0 9 11 11 2
38 3 13 2 16 9 1 9 1 11 7 0 9 13 0 2 9 7 1 11 2 7 1 11 15 13 9 7 9 13 1 9 9 2 13 9 11 11 2
9 13 2 16 4 0 9 13 0 2
22 0 9 1 0 9 13 0 7 13 15 9 2 15 13 1 15 0 2 13 0 9 2
2 9 9
1 9
7 10 0 9 13 9 9 2
16 13 15 9 0 2 9 9 13 0 9 2 3 9 9 13 2
39 13 3 1 10 0 9 2 13 9 7 9 0 7 0 9 2 13 0 9 9 7 13 7 9 13 9 0 7 0 9 1 9 0 9 7 13 9 9 2
25 1 0 9 15 13 13 10 9 3 0 2 3 2 15 4 13 13 0 1 9 9 9 0 9 2
23 3 9 1 0 9 1 11 12 13 0 9 9 0 7 0 1 12 1 0 9 9 9 2
7 9 10 9 7 13 0 2
34 9 0 9 11 2 15 13 1 10 9 12 1 12 9 0 9 2 15 3 13 1 15 2 16 9 0 9 13 12 1 10 0 9 2
20 1 9 10 9 9 2 11 11 13 0 0 9 1 10 9 9 7 1 9 2
13 3 0 9 13 0 9 2 15 13 7 9 11 2
32 9 9 3 1 10 9 9 1 0 0 9 3 13 2 16 13 2 16 13 1 9 3 10 9 9 2 14 2 14 14 12 2
33 13 3 0 2 16 1 9 0 9 9 2 7 3 7 9 15 9 2 15 15 13 0 9 2 13 0 13 10 9 9 0 9 2
17 7 1 0 9 15 13 13 0 2 3 0 9 9 1 9 9 2
30 3 9 9 13 9 1 9 2 10 2 0 9 7 4 13 1 9 9 0 9 2 16 4 9 13 3 3 0 9 2
24 7 4 13 1 0 9 1 15 2 16 4 15 0 9 13 2 15 7 4 3 13 9 9 2
12 1 9 9 7 13 0 13 9 2 7 9 2
19 0 9 1 9 9 2 12 1 9 0 9 2 15 9 9 1 9 13 2
19 7 15 13 13 0 2 16 9 1 0 9 9 13 0 7 0 9 0 2
4 0 2 0 9
1 9
12 9 9 13 13 2 13 15 13 2 13 0 2
10 3 15 15 0 9 9 11 11 13 2
12 9 1 10 9 1 0 9 1 10 9 13 2
23 0 9 13 13 0 2 3 7 13 9 2 15 15 13 2 3 2 9 9 9 1 9 2
16 13 15 1 0 9 7 9 9 7 13 0 9 13 9 0 2
24 0 9 7 13 3 0 2 16 4 13 9 0 0 9 1 0 0 9 0 1 0 0 9 2
16 9 7 13 3 13 1 9 9 2 0 15 9 10 0 9 2
13 14 3 2 16 4 10 9 13 3 3 0 9 2
17 13 7 0 9 2 3 15 13 13 2 1 9 7 1 0 9 2
5 9 13 12 9 2
14 13 2 14 7 9 2 16 13 3 13 2 13 3 2
9 9 7 9 13 10 0 0 9 2
20 13 2 14 1 15 3 1 9 2 13 3 13 2 16 13 0 7 0 9 2
25 13 3 9 2 16 15 1 10 9 13 1 9 0 7 16 15 15 15 13 1 9 1 9 0 2
21 9 1 9 9 13 9 13 15 2 16 13 10 10 9 1 9 1 9 0 9 2
6 9 15 13 0 9 2
16 7 9 2 16 15 15 15 1 9 3 13 2 13 3 0 2
26 3 11 2 11 2 15 9 9 1 10 9 13 2 4 13 3 3 9 2 16 4 15 1 9 13 2
6 13 3 9 0 9 2
10 11 11 15 7 13 9 9 1 11 2
9 15 15 11 11 1 0 9 13 2
15 10 9 4 3 1 9 9 13 1 9 9 1 0 9 2
7 0 9 4 13 1 15 2
13 9 4 15 13 13 1 9 2 15 13 1 9 2
22 9 14 13 13 3 2 3 13 10 9 2 1 0 9 13 13 10 9 2 15 13 2
25 1 1 0 0 9 9 7 1 15 0 9 0 0 9 13 7 14 3 13 0 9 10 0 9 2
24 16 11 1 0 9 13 2 16 11 13 1 10 9 0 9 2 13 15 3 9 0 1 9 2
3 0 9 13
1 9
35 9 11 11 1 0 9 15 1 9 2 11 15 13 0 9 2 1 10 9 13 2 16 4 14 1 0 9 0 9 13 9 1 11 11 2
5 9 13 3 0 2
22 3 1 9 0 9 9 4 1 15 13 1 9 2 13 15 1 9 10 9 1 9 2
14 3 13 1 12 1 9 7 13 15 2 16 4 13 2
35 1 9 13 9 11 7 3 15 15 13 2 16 4 13 13 9 3 2 3 2 3 4 15 3 13 2 2 16 15 13 13 1 10 9 2
10 3 15 1 15 13 7 9 1 11 2
15 13 4 2 16 9 1 11 11 13 7 1 0 0 9 2
19 9 9 11 2 16 4 13 3 13 9 1 0 9 2 13 0 0 9 2
15 13 3 14 10 9 2 16 4 15 3 13 1 9 9 2
25 10 9 3 13 2 16 4 13 9 2 16 4 1 9 13 0 9 2 9 11 1 9 1 11 2
23 1 15 1 15 13 0 2 3 3 13 2 16 4 1 10 9 13 0 15 1 0 9 2
1 9
14 9 0 9 13 1 9 0 2 0 9 12 0 9 2
10 9 15 4 13 1 9 1 0 9 2
11 9 13 2 16 9 1 9 13 1 9 2
8 7 1 12 9 15 7 13 2
9 1 11 13 12 12 9 9 9 0
2 11 2
35 3 12 9 9 9 0 1 9 3 12 9 13 1 3 0 9 1 9 1 9 1 9 1 9 9 1 9 0 0 9 1 11 1 11 2
14 9 9 9 15 13 9 3 1 9 7 9 0 9 2
3 0 9 13
2 11 2
23 9 0 9 1 11 13 3 1 9 0 9 12 0 9 7 1 15 13 1 9 12 9 2
12 1 9 12 15 13 9 0 9 1 12 12 2
19 9 13 9 2 15 13 9 9 2 9 7 9 1 9 7 13 0 9 2
17 13 3 0 9 1 9 0 9 2 3 4 13 4 13 0 9 2
9 1 9 0 9 13 9 11 11 9
2 11 2
17 9 1 9 2 15 13 11 11 3 0 9 1 11 2 13 0 2
13 3 15 13 0 9 11 11 2 9 1 0 9 2
21 1 9 4 13 7 9 1 0 9 7 0 9 2 15 15 13 1 10 0 9 2
14 9 13 1 9 12 15 9 2 15 0 13 10 9 2
36 11 11 4 13 1 0 9 1 11 3 1 9 0 9 7 0 9 2 15 13 13 9 1 9 1 11 7 15 15 13 13 9 0 9 9 2
7 0 0 9 13 10 9 2
34 0 9 3 13 2 16 1 0 9 1 0 9 13 7 15 2 3 13 1 9 12 9 9 13 11 11 2 0 9 11 2 11 2 2
9 3 13 1 10 9 13 11 11 2
25 11 15 7 13 2 16 10 9 13 1 9 2 16 0 9 0 9 13 2 13 2 13 7 13 2
28 9 3 13 10 9 9 1 0 9 9 3 0 9 7 13 1 9 2 15 13 7 15 13 2 16 13 0 2
24 9 3 13 9 2 13 0 9 3 0 9 9 2 13 0 9 9 7 13 15 10 0 9 2
14 3 1 0 9 1 12 2 7 12 2 9 13 9 2
20 0 9 3 1 9 12 4 13 1 0 9 2 15 4 13 1 12 9 3 2
27 9 9 0 9 2 15 4 13 1 0 9 2 13 3 0 2 7 3 13 1 9 2 3 9 13 13 2
15 1 11 2 11 13 1 9 13 10 9 10 9 11 11 2
21 13 15 3 13 9 0 0 9 2 15 1 11 10 9 13 1 9 1 9 12 2
23 10 9 1 9 1 0 9 15 13 11 13 1 9 12 1 15 1 0 9 1 0 9 2
23 3 2 16 13 9 2 16 13 9 7 1 9 9 2 13 1 15 1 9 12 0 9 2
8 0 9 13 0 9 10 0 9
2 11 2
18 9 0 9 2 0 9 7 9 0 9 13 0 9 9 0 0 9 2
25 13 15 15 1 9 0 9 1 9 2 9 9 2 9 7 9 2 2 15 13 13 0 9 11 2
16 9 1 0 9 13 1 9 11 13 1 9 0 9 1 9 2
18 2 0 13 13 9 13 9 1 3 0 9 2 2 13 15 1 9 2
11 9 0 9 4 13 13 13 1 9 9 2
21 0 9 4 7 13 13 1 0 9 0 0 9 2 0 2 3 0 9 9 2 2
11 1 10 9 13 11 13 0 2 0 9 2
26 13 4 15 13 9 0 9 2 15 4 13 9 1 0 9 7 13 0 9 7 0 9 1 0 9 2
14 1 0 9 13 0 9 0 9 0 9 1 0 9 2
18 1 0 9 9 13 0 9 2 15 13 2 0 9 1 0 9 2 2
12 0 9 0 9 11 13 13 9 7 9 9 2
11 0 9 13 9 9 1 9 0 9 9 2
24 2 13 1 9 2 16 9 1 9 13 0 0 9 0 9 2 2 13 11 1 9 0 9 2
18 0 9 13 13 0 0 2 0 2 0 2 0 2 0 7 0 9 2
22 0 9 13 13 3 0 9 2 0 9 9 9 9 1 0 3 0 9 7 9 2 2
13 11 13 0 9 3 2 3 9 13 9 9 9 2
17 9 13 0 13 10 2 0 9 2 15 9 2 13 15 1 9 2
22 16 3 11 13 9 11 11 11 2 0 9 9 4 13 13 0 9 9 9 0 9 2
5 0 9 13 14 0
9 10 9 13 9 0 9 9 1 0
2 11 2
32 16 9 9 13 9 11 11 2 16 9 0 0 9 11 4 1 0 9 13 12 7 12 9 2 9 9 15 13 1 0 9 2
19 9 0 9 11 11 2 11 2 9 11 13 2 16 10 9 13 3 0 2
13 2 3 4 15 7 10 10 9 13 2 2 13 2
23 15 1 15 13 15 2 16 9 4 3 13 7 0 11 4 13 3 2 12 0 9 2 2
28 1 0 9 13 1 9 9 9 1 9 12 9 11 13 2 16 13 1 9 0 7 12 9 4 13 0 9 2
9 2 0 15 3 13 2 2 13 2
15 13 2 16 3 9 13 12 9 7 3 13 13 1 12 2
19 3 9 11 11 2 11 2 13 2 16 11 0 9 9 9 13 3 13 2
10 13 15 2 16 13 0 13 9 0 2
20 2 13 2 14 10 9 13 9 1 9 1 10 9 2 4 13 2 2 13 2
26 11 13 1 15 1 10 9 0 1 9 1 0 9 0 11 2 16 0 9 1 9 13 3 0 9 2
18 1 9 9 13 2 16 15 13 1 10 0 9 2 3 2 7 0 2
12 11 11 2 11 2 0 0 9 9 3 13 2
15 13 14 0 3 1 9 2 16 15 13 9 9 10 9 2
10 9 1 0 9 3 13 4 2 13 2
11 13 3 9 9 0 9 1 3 12 9 2
19 15 1 15 13 1 0 9 3 2 16 15 13 3 1 2 0 9 2 2
19 11 13 2 16 1 0 9 13 9 2 16 13 3 9 7 13 0 9 2
8 0 9 13 13 0 9 0 9
2 11 2
38 0 9 9 3 9 9 12 2 12 2 12 15 13 2 13 13 1 9 9 9 9 1 0 9 2 15 13 9 11 11 7 11 11 2 12 11 2 2
14 9 13 4 13 0 9 0 9 2 0 3 1 9 2
33 9 0 9 9 1 0 9 1 12 12 9 13 3 15 2 16 13 0 9 3 13 7 3 16 4 15 13 2 13 1 10 9 2
27 11 11 2 11 2 13 2 16 13 1 0 9 2 13 7 2 16 3 13 0 9 2 3 0 9 13 2
48 9 11 3 13 2 16 9 11 1 0 0 9 13 1 0 9 13 1 9 2 3 1 10 9 4 13 1 0 9 9 7 0 9 2 16 4 7 13 0 13 9 10 0 9 1 0 9 2
17 2 13 15 9 2 2 13 11 7 13 9 0 9 3 0 9 2
31 2 15 4 13 10 9 2 15 13 1 2 16 15 15 9 9 13 2 2 13 1 9 9 9 9 11 11 2 11 2 2
17 13 1 9 9 2 16 1 9 0 9 15 13 7 10 0 9 2
39 0 9 3 3 13 9 1 9 9 9 11 11 7 11 11 2 12 11 2 2 15 4 13 3 13 2 0 2 9 2 0 3 3 16 12 12 9 9 2
13 9 3 3 13 9 9 2 15 9 0 9 13 2
8 9 0 9 13 13 9 0 9
2 11 2
16 0 9 11 4 7 3 13 13 12 2 9 7 12 2 9 2
38 10 9 13 0 9 0 9 2 15 3 13 9 9 9 1 0 9 0 12 9 9 1 9 1 11 2 11 2 11 2 7 11 2 11 2 11 2 2
31 9 13 1 9 0 9 12 2 9 2 9 0 9 2 7 12 2 9 2 9 9 11 2 2 7 1 9 12 2 9 2
10 12 0 9 4 13 13 9 0 9 2
66 0 7 0 9 9 13 2 16 4 1 0 9 9 1 9 2 7 2 3 9 0 9 2 3 13 0 9 2 9 0 2 12 2 9 2 12 2 7 12 2 9 2 12 2 7 12 2 9 2 15 0 7 9 0 2 7 12 2 2 12 2 7 12 2 9 2
18 3 0 2 0 2 9 13 13 3 2 9 1 9 1 9 15 9 2
88 0 9 10 9 4 1 9 0 9 9 1 9 13 13 2 12 2 9 2 12 9 2 2 12 2 9 2 9 11 2 2 12 2 9 2 9 11 2 11 2 11 2 2 12 2 9 2 9 9 0 2 2 12 2 9 2 9 1 9 12 2 2 12 2 9 2 9 11 11 2 2 12 2 9 2 0 2 11 2 7 12 2 9 2 9 9 2 2
4 9 1 9 9
2 11 2
15 9 9 2 12 9 2 13 1 9 0 9 9 1 9 2
15 13 15 1 9 2 15 9 0 9 13 0 9 0 9 2
29 1 9 12 9 9 3 13 2 16 12 9 0 1 9 9 11 15 13 2 16 15 9 13 13 1 9 0 9 2
6 9 1 9 13 1 9
3 9 0 9
23 9 4 13 0 0 9 2 15 13 13 9 1 9 7 9 9 1 9 1 9 7 9 2
5 3 10 9 13 2
20 11 11 2 11 2 2 9 0 9 2 9 9 1 9 9 1 9 13 0 2
19 9 4 13 14 0 9 2 16 9 13 0 9 2 7 3 13 0 9 2
10 13 0 2 16 4 9 13 3 15 2
17 11 11 2 11 2 2 9 0 9 2 13 15 3 9 0 9 2
7 3 15 11 13 0 9 2
24 15 13 2 16 4 13 9 2 7 15 4 13 1 9 10 2 15 15 13 2 15 13 9 2
20 11 11 2 11 2 2 9 2 10 9 13 1 0 9 13 9 0 0 9 2
19 1 10 9 13 2 16 15 13 2 16 13 3 9 0 9 7 0 9 2
14 0 0 9 13 7 9 7 9 1 9 9 13 3 2
22 11 11 2 11 2 2 9 2 1 10 0 9 13 0 13 0 9 1 9 0 9 2
16 15 13 2 16 1 0 9 4 9 9 13 1 10 9 13 2
24 13 0 2 16 4 15 1 15 2 15 13 3 2 3 13 2 7 10 9 13 3 13 9 2
31 11 11 0 2 2 11 2 2 9 2 9 13 1 15 2 16 9 4 3 13 9 2 7 13 15 9 9 1 0 9 2
6 1 15 13 16 13 2
8 11 2 11 2 13 1 9 11
2 11 2
44 2 7 15 2 3 16 0 9 7 0 9 0 9 2 13 9 1 15 2 16 4 15 11 13 1 9 2 2 13 3 11 0 9 9 9 11 11 1 9 1 0 9 11 2
21 9 11 13 11 0 0 9 2 15 13 13 9 11 1 0 9 11 1 0 9 2
27 9 9 13 13 13 1 9 9 11 11 11 11 2 15 3 13 0 0 9 9 9 9 11 11 2 11 2
23 2 9 13 3 9 1 0 9 1 11 2 15 3 13 9 9 1 9 2 2 13 11 2
24 1 10 9 13 11 1 0 9 1 9 1 9 7 11 10 9 1 9 13 1 10 9 13 2
5 9 13 1 9 9
2 11 2
32 0 9 0 9 4 13 13 1 9 0 9 0 9 9 2 15 4 13 0 9 9 1 9 9 1 9 12 9 0 0 9 2
9 9 13 9 11 2 11 7 9 2
23 13 15 1 15 3 0 9 0 2 1 0 9 7 9 3 2 16 13 9 0 0 9 2
26 1 0 9 4 15 9 9 13 13 3 0 9 2 1 9 11 7 11 7 10 0 9 7 0 0 2
10 0 9 3 13 1 0 9 9 9 2
8 9 13 0 9 9 9 1 9
2 11 2
16 9 3 13 12 9 9 9 1 9 9 11 2 11 7 11 2
16 9 13 9 11 2 11 15 2 16 9 13 1 9 1 9 2
14 13 4 9 9 0 9 1 11 7 10 9 0 9 2
11 9 4 1 10 9 13 0 3 13 9 2
25 9 13 2 16 9 2 15 4 15 13 0 9 2 13 1 9 13 2 7 7 13 0 9 0 2
28 9 3 13 12 0 9 9 9 1 0 9 2 15 13 1 9 9 9 1 0 12 1 12 2 3 2 12 2
25 1 11 4 0 9 9 13 13 0 2 3 4 15 14 7 13 13 13 11 15 0 16 9 9 2
18 9 13 7 9 1 9 0 9 1 0 9 1 11 1 9 10 9 2
17 1 9 9 9 11 13 2 16 13 1 9 9 2 3 0 9 2
7 0 9 15 13 1 0 9
2 11 2
29 1 9 0 9 1 11 7 9 9 3 0 1 0 9 1 9 13 1 9 9 12 0 0 9 9 1 3 0 2
13 1 10 9 9 13 9 2 0 9 7 9 9 2
36 9 0 9 9 9 2 13 1 15 13 3 12 5 9 1 0 0 9 2 4 1 11 3 13 7 3 0 13 1 0 9 9 2 13 9 2
17 9 9 9 13 0 9 2 1 15 9 13 2 9 7 9 9 2
19 1 0 9 2 13 15 1 9 2 13 9 0 3 0 3 3 0 9 2
8 1 11 15 3 10 9 13 2
8 9 3 13 7 3 0 9 2
13 1 0 15 3 13 0 9 7 1 9 13 9 2
17 9 13 9 2 16 0 9 9 13 13 0 2 16 4 15 13 2
15 9 13 3 14 1 0 9 2 15 13 3 9 10 9 2
9 11 13 1 0 9 12 3 0 2
25 0 1 15 13 3 1 12 9 2 13 0 9 7 9 1 9 13 1 0 9 0 9 1 9 2
15 13 7 3 1 9 2 16 3 1 9 0 13 1 9 2
16 0 9 15 1 0 9 1 0 9 13 12 7 12 9 3 2
19 11 13 1 15 2 16 1 9 9 13 9 1 9 0 9 1 0 9 2
23 9 9 9 1 11 12 11 11 3 13 2 16 9 11 13 3 3 0 2 16 13 9 2
15 15 13 3 13 3 0 1 0 9 14 1 12 12 9 2
18 9 2 3 15 9 3 13 2 13 0 9 1 9 1 0 0 9 2
13 9 13 3 1 9 9 7 0 9 1 10 9 2
10 11 13 0 0 9 7 1 0 9 2
14 3 14 9 13 14 15 2 16 13 9 1 10 9 2
8 13 9 13 0 2 13 9 11
2 11 2
21 9 2 15 1 9 13 9 9 7 15 3 13 2 4 1 10 9 3 3 13 2
15 0 9 3 13 2 16 4 13 2 16 9 13 9 0 2
6 15 13 7 3 0 2
12 11 15 3 13 9 9 11 11 2 11 2 2
17 1 0 9 7 13 9 13 9 1 9 9 0 9 1 0 9 2
31 11 13 0 0 9 13 2 16 4 9 2 9 1 9 7 9 2 13 9 13 1 9 10 9 3 2 3 13 1 0 2
25 1 10 0 9 4 15 13 13 9 7 15 4 7 13 13 9 13 2 3 13 3 2 3 13 2
34 2 16 1 15 1 9 13 12 9 1 9 7 9 2 4 15 13 2 16 15 13 3 2 7 16 13 2 16 15 13 13 7 13 2
21 16 1 10 9 13 9 7 15 4 1 9 13 2 3 3 13 2 2 13 11 2
6 2 13 9 13 15 2
18 1 15 2 16 9 13 7 13 2 4 13 13 10 9 2 2 13 2
6 0 9 4 1 11 13
2 11 2
24 13 0 9 3 12 9 0 9 1 0 0 9 15 13 9 0 0 9 1 9 1 12 9 2
8 13 15 3 10 9 11 11 2
16 13 2 16 0 9 1 10 9 13 9 9 9 7 0 9 2
38 15 3 13 9 2 16 0 9 13 13 1 0 0 9 1 11 2 9 11 11 7 13 1 9 1 9 10 9 1 9 3 0 9 7 9 0 9 2
22 0 0 9 1 0 9 2 15 4 13 1 0 9 13 0 9 2 13 0 0 9 2
5 0 9 1 9 9
2 11 2
27 1 0 9 1 11 2 15 13 1 0 0 9 1 9 2 4 13 9 12 9 0 0 9 0 0 9 2
12 13 15 9 0 2 9 2 9 11 11 11 2
18 9 4 1 11 13 1 9 1 0 9 9 7 13 3 1 0 9 2
11 0 0 9 4 13 1 9 12 7 12 2
10 1 0 9 9 13 0 9 12 9 2
16 9 13 13 1 9 9 7 9 2 13 3 16 9 0 9 2
8 13 15 7 1 9 9 11 2
8 9 13 0 9 1 12 9 2
19 15 0 2 15 4 13 0 7 0 9 2 13 13 1 0 9 0 9 2
3 9 4 13
2 11 2
24 1 0 9 11 1 0 9 1 11 15 13 1 12 2 12 2 12 13 10 0 9 2 9 2
17 13 1 15 9 9 2 0 9 7 9 9 2 9 0 11 11 2
19 1 0 9 11 11 1 9 0 11 13 9 0 9 13 11 16 0 9 2
11 13 13 0 9 9 7 9 1 10 9 2
8 15 9 3 16 9 11 13 2
15 0 9 9 14 1 15 13 9 12 2 9 9 9 11 2
21 1 11 7 13 9 3 0 2 7 7 9 9 13 9 1 9 1 9 0 9 2
9 15 13 13 1 11 9 0 9 2
10 9 13 1 9 9 0 11 3 0 2
36 11 11 1 9 0 9 11 13 2 16 9 13 3 1 15 2 16 4 9 0 9 13 1 9 3 7 16 4 9 13 1 9 1 10 9 2
6 11 13 3 0 9 2
27 9 13 2 16 15 1 9 13 12 2 9 12 1 9 14 3 13 2 7 13 3 3 0 3 0 9 2
18 1 10 9 13 1 11 9 9 1 9 9 7 1 9 0 9 9 2
3 0 9 13
2 11 2
16 0 9 0 9 1 11 1 0 9 15 13 1 0 9 9 2
28 9 10 0 9 13 10 0 9 11 11 9 2 2 0 9 9 11 13 1 3 0 9 2 9 13 0 2 2
23 16 15 11 13 1 11 2 3 4 14 13 9 1 0 9 2 16 13 1 15 0 9 2
19 2 13 3 3 2 16 10 9 13 13 15 0 9 11 1 12 9 2 2
16 0 0 9 13 1 11 11 0 9 13 1 12 9 0 11 2
17 13 3 1 0 9 2 9 2 9 2 7 3 0 9 7 9 2
24 1 0 9 2 0 9 7 3 0 2 13 0 9 3 3 0 7 3 0 1 9 7 9 2
7 11 15 13 9 9 1 11
2 11 2
17 11 11 2 11 11 7 0 9 0 9 4 1 9 13 1 11 2
25 11 11 7 0 9 11 2 11 13 1 11 7 1 0 9 13 9 0 9 2 9 2 0 2 2
13 13 1 0 9 2 15 4 13 3 13 0 9 2
9 9 7 3 13 0 9 0 9 2
34 11 11 1 9 11 11 2 15 13 0 9 0 9 2 3 13 2 16 15 13 1 0 9 1 15 2 15 15 4 13 3 0 9 2
23 3 13 2 16 15 9 4 1 0 12 7 12 9 13 9 7 0 0 9 2 7 9 2
22 4 14 13 7 0 9 7 13 15 1 9 9 2 16 4 1 15 13 0 9 9 2
33 9 0 9 11 12 11 11 2 15 1 9 1 9 13 13 2 3 13 11 13 2 10 0 9 4 0 9 13 1 9 0 9 2
28 13 7 2 16 9 13 9 2 3 0 9 13 3 1 0 9 1 0 9 2 3 0 9 13 9 3 3 2
21 1 3 0 9 13 9 0 2 7 15 13 3 1 0 9 0 9 7 0 9 2
16 1 9 2 9 2 0 2 15 7 3 13 1 9 10 9 2
31 11 2 11 13 2 16 9 13 13 1 0 12 7 12 9 1 9 15 9 2 15 4 13 9 0 2 3 7 0 9 2
4 9 13 9 9
2 11 2
19 3 3 13 1 0 9 0 0 9 1 11 13 15 3 0 9 7 9 2
19 1 10 9 7 13 9 2 15 13 0 9 13 2 16 13 9 0 9 2
26 9 13 10 9 2 7 13 3 9 0 7 0 9 2 3 13 12 7 12 0 9 7 0 9 3 2
18 9 9 9 2 11 11 13 2 16 9 9 13 13 14 1 0 9 2
16 3 7 10 9 13 2 16 4 4 0 10 9 13 0 9 2
6 0 9 13 9 9 2
6 15 7 13 0 9 2
14 1 10 9 4 13 2 16 9 13 0 13 9 0 2
10 9 1 10 9 4 13 3 1 11 2
16 2 13 7 12 7 15 15 9 13 13 2 2 13 11 11 2
18 9 15 7 13 13 1 9 1 0 9 2 15 13 11 11 11 11 2
22 9 9 13 9 7 10 9 13 9 2 15 13 13 10 0 9 2 1 0 9 2 2
17 13 0 9 2 15 15 1 11 13 0 9 7 13 15 10 9 2
14 1 0 9 4 13 3 10 9 1 0 9 7 9 2
16 3 15 9 13 1 12 12 0 9 7 13 1 15 0 9 2
12 9 1 0 9 1 11 2 13 2 12 9 2
28 2 3 1 15 13 12 10 9 2 2 13 11 11 11 2 15 13 2 16 0 7 0 9 13 3 1 9 2
12 2 13 15 2 16 13 15 0 16 9 2 2
5 9 15 13 9 9
2 11 2
25 9 15 3 13 0 9 2 9 9 2 2 15 13 1 9 9 9 9 2 0 9 11 2 0 2
21 3 1 9 15 13 0 9 1 9 1 0 9 7 1 11 1 11 13 0 9 2
14 1 9 3 10 9 13 0 9 9 0 9 1 11 2
21 0 0 9 1 15 2 9 2 13 12 12 9 2 1 15 12 12 0 12 9 2
3 9 0 9
2 11 2
21 1 0 9 13 9 1 0 0 9 11 11 2 11 2 7 11 11 2 11 2 2
20 11 13 1 0 9 11 9 2 1 15 13 9 9 0 1 10 9 9 11 2
10 9 15 13 9 9 7 9 0 9 2
34 9 9 11 13 3 9 0 9 1 0 9 11 2 11 2 9 9 11 1 0 7 0 9 11 2 11 7 3 15 13 1 9 9 2
7 11 3 9 11 11 13 2
26 13 2 16 13 0 0 9 9 2 3 16 4 13 9 0 0 9 1 9 9 0 9 1 11 2 2
4 3 1 0 9
3 9 0 9
9 9 3 13 9 9 0 0 9 2
16 0 9 13 0 9 2 15 10 9 13 1 0 9 0 9 2
18 1 9 0 9 1 9 12 13 1 0 2 0 9 2 1 0 9 2
8 15 0 15 3 3 4 13 2
28 1 0 12 9 3 3 3 13 1 0 9 2 10 9 15 7 4 3 13 0 9 7 0 9 15 3 13 2
10 0 0 9 3 4 13 3 0 9 2
29 16 15 0 13 2 15 13 13 2 3 3 13 3 1 0 2 7 3 3 15 0 2 9 15 2 15 13 13 2
5 13 4 3 0 2
41 13 2 14 9 13 7 13 0 9 3 1 9 2 3 1 0 9 9 0 9 4 13 14 3 0 9 9 0 9 2 1 0 7 0 9 2 1 9 1 9 2
3 3 15 2
16 3 10 9 4 7 1 10 0 9 13 14 1 9 0 9 2
21 16 1 9 12 4 13 0 0 9 2 13 15 9 9 9 7 9 1 0 9 2
12 9 0 9 2 9 0 9 2 9 0 9 2
26 1 0 9 13 9 0 2 16 1 0 9 3 1 9 9 2 1 9 2 0 9 7 9 0 9 2
15 0 9 7 3 13 9 3 0 7 1 9 0 4 13 2
7 1 15 13 3 3 9 2
25 0 9 3 14 16 13 0 1 0 9 1 9 2 7 3 4 13 0 9 0 9 1 0 9 2
23 13 0 0 9 2 15 13 9 1 9 2 7 7 3 13 0 3 3 13 0 15 9 2
10 13 3 9 2 16 1 9 9 13 2
3 3 14 2
12 1 0 9 15 13 13 16 1 15 3 0 2
28 0 9 9 13 1 9 7 0 9 15 13 12 9 9 2 15 1 1 9 10 0 9 13 9 9 0 9 2
7 9 3 3 7 13 3 2
19 3 16 15 9 13 13 2 7 16 15 3 13 13 2 9 2 15 13 2
4 9 11 13 9
10 15 13 0 9 2 13 1 9 9 13
2 11 2
22 3 12 0 9 13 13 9 0 9 2 11 2 15 2 15 13 0 9 1 9 9 2
7 0 1 15 13 9 9 2
11 11 13 9 3 1 9 9 1 12 9 2
14 1 15 12 9 13 9 1 9 9 7 12 9 9 2
14 2 0 9 13 2 2 13 15 9 9 11 11 11 2
10 1 9 12 13 9 3 12 9 9 2
13 3 13 0 9 2 15 4 13 9 9 9 13 2
15 9 4 13 13 9 9 1 0 9 2 15 13 9 9 2
20 1 9 0 9 11 13 9 15 2 16 15 13 9 1 9 9 1 0 9 2
19 1 9 9 13 3 1 9 0 1 9 9 2 0 9 7 9 1 9 2
17 9 9 13 3 9 2 15 13 0 9 7 13 15 9 1 9 2
20 0 0 9 2 15 11 13 9 2 13 13 9 2 15 9 13 13 1 9 2
31 15 13 9 2 13 13 7 1 15 2 16 1 15 4 11 13 1 10 0 9 2 15 13 9 3 1 0 9 1 9 2
19 16 9 9 1 11 13 0 9 2 13 1 0 0 9 1 9 9 13 2
22 13 2 16 9 1 9 9 2 9 9 2 13 14 3 1 9 1 9 1 9 11 2
12 1 0 9 13 1 9 11 14 12 9 3 2
12 9 3 13 1 9 9 7 13 9 0 9 2
12 2 15 13 0 9 2 2 13 11 2 11 2
16 1 15 13 0 9 7 9 1 9 13 3 7 9 0 9 2
15 1 9 1 11 13 0 2 16 4 9 13 0 9 9 2
24 9 9 13 9 9 2 16 3 2 9 9 2 15 13 1 9 0 9 3 2 15 13 13 2
11 3 9 15 3 13 0 9 12 9 1 9
2 11 2
24 9 12 9 3 1 0 12 9 9 1 9 13 0 13 7 1 15 2 15 1 10 9 13 2
10 11 15 13 9 9 9 11 2 11 2
11 9 15 13 1 9 9 13 13 1 9 2
19 1 10 9 13 0 9 1 9 9 2 9 7 9 13 3 1 9 9 2
15 3 13 0 14 15 2 16 13 15 4 14 1 9 9 2
11 9 1 11 13 2 16 9 3 13 9 2
15 9 15 14 3 4 3 13 1 15 2 16 9 3 13 2
19 9 13 2 16 0 4 7 1 9 10 9 1 9 3 13 3 2 9 2
25 0 3 4 13 1 15 9 2 9 7 0 9 0 1 9 2 1 15 13 12 9 13 2 13 2
21 3 0 2 1 15 13 9 1 10 9 2 4 14 13 13 9 9 7 0 9 2
26 9 2 15 9 13 4 2 7 3 3 3 13 13 2 13 4 1 9 13 2 16 15 13 10 9 2
19 11 13 2 16 9 13 9 0 9 2 15 13 9 7 15 9 13 9 2
15 2 15 4 13 1 9 3 16 12 9 2 2 13 11 2
15 9 9 3 13 2 16 9 4 13 14 0 12 9 3 2
22 4 2 14 7 15 13 1 9 1 9 15 2 3 13 14 0 12 9 1 0 9 2
9 15 4 13 3 9 0 12 9 2
8 9 13 3 7 9 1 9 2
16 11 13 2 16 0 9 9 1 9 13 1 0 9 12 9 2
4 0 9 1 11
2 11 2
28 0 9 0 7 0 9 0 9 1 0 9 0 11 13 3 1 11 0 9 11 11 7 10 0 9 11 11 2
29 12 9 1 15 13 10 9 13 9 9 1 9 9 9 7 3 7 9 0 9 11 7 11 1 9 1 9 9 2
25 9 3 13 9 0 9 2 1 15 4 13 13 16 9 9 1 11 2 7 9 9 9 1 11 2
15 12 9 13 9 1 0 9 2 15 4 13 0 9 9 2
13 9 13 10 0 9 1 11 1 9 1 9 11 2
4 3 1 9 12
4 9 0 9 13
2 11 2
20 9 3 13 9 1 9 0 0 9 2 15 0 9 13 0 9 1 0 9 2
11 1 0 9 9 1 15 13 9 11 11 2
14 9 13 2 16 9 4 13 3 1 0 9 0 9 2
27 9 1 0 9 4 15 1 0 9 13 13 3 2 7 15 1 9 0 9 3 1 9 12 7 12 9 2
35 0 9 2 15 9 13 9 9 1 0 9 0 9 2 13 1 9 0 0 9 10 0 9 7 9 2 15 4 3 1 9 0 9 13 2
5 0 9 1 0 9
13 1 0 9 7 1 11 13 9 1 9 9 9 9
2 11 2
15 0 9 9 12 2 9 9 0 0 9 13 3 0 9 2
15 9 15 13 3 9 9 11 11 7 9 0 9 11 11 2
20 1 9 4 13 9 0 9 7 9 0 12 0 9 15 13 7 9 15 0 2
31 0 9 9 13 0 9 0 9 12 2 9 1 11 1 0 9 1 9 0 9 2 9 0 9 7 9 12 2 0 9 2
10 1 9 13 9 1 9 12 9 9 2
25 9 11 1 9 1 9 9 13 2 16 1 9 13 9 2 16 4 1 9 4 13 7 9 11 2
19 9 11 11 7 1 9 9 11 13 2 16 9 1 10 9 3 3 13 2
18 13 7 1 15 2 16 4 15 1 9 9 9 1 9 13 0 9 2
23 1 11 1 0 15 9 13 9 1 15 2 16 12 2 9 12 13 9 2 7 9 11 2
25 0 9 11 15 13 1 9 0 9 11 1 11 1 9 12 2 2 12 2 9 13 9 9 2 2
15 9 11 11 13 9 13 1 9 9 11 1 10 0 9 2
19 13 4 15 13 9 9 9 12 2 9 1 11 7 1 9 3 1 11 2
20 11 15 3 13 0 12 2 9 9 9 0 9 0 9 1 11 12 2 9 2
23 9 9 4 13 13 9 0 9 11 11 16 9 9 11 2 15 4 9 1 9 3 13 2
8 1 12 9 3 13 3 13 2
6 0 9 1 11 7 11
2 11 2
24 1 0 9 15 9 0 2 11 13 1 0 9 13 0 12 9 9 0 11 7 0 9 11 2
12 1 0 9 9 11 13 1 3 16 12 5 2
17 0 13 1 9 12 1 0 11 2 3 15 9 13 1 12 9 2
11 11 15 3 13 0 0 0 9 1 9 2
16 9 11 13 3 1 11 7 1 0 9 0 9 1 12 9 2
25 3 15 9 0 2 11 13 1 9 12 13 1 3 16 12 9 9 10 9 3 16 1 0 9 2
4 11 11 13 0
2 11 2
23 9 11 11 2 15 13 1 9 0 9 3 9 2 13 1 0 9 9 1 12 9 9 2
18 9 9 2 15 13 16 0 2 7 7 0 9 2 13 3 14 12 2
31 0 9 9 9 13 9 7 9 9 7 9 1 15 0 2 3 9 0 9 2 0 9 7 9 1 0 9 1 9 9 2
16 9 13 9 0 9 2 7 15 13 3 1 0 7 0 9 2
13 1 9 9 13 0 9 1 9 12 9 2 9 2
23 9 13 10 0 9 0 9 2 7 9 15 13 3 1 0 9 0 12 5 0 9 9 2
4 9 13 1 11
2 11 2
31 1 9 11 2 11 9 13 4 1 12 2 9 13 0 9 9 1 9 11 2 11 2 11 9 0 9 0 7 0 11 2
27 13 13 0 0 9 1 11 7 11 1 0 0 9 1 9 9 12 9 1 9 9 7 12 9 1 9 2
21 11 2 11 9 11 4 13 0 9 1 9 0 9 14 1 9 9 9 1 9 2
30 11 13 1 10 9 13 2 16 10 0 0 9 13 9 0 9 9 1 0 9 1 9 0 0 9 3 1 9 11 2
8 11 11 15 13 1 9 9 9
2 11 2
16 0 9 9 9 1 0 9 13 9 1 0 9 7 11 11 2
28 16 9 3 13 9 9 10 9 1 0 9 2 3 13 0 15 13 1 12 9 2 7 15 3 1 0 9 2
27 1 9 12 15 13 1 9 9 3 12 7 12 9 2 1 9 12 13 15 3 12 9 7 9 3 13 2
13 11 13 1 9 9 3 1 0 9 0 0 9 2
13 1 10 9 7 13 3 0 9 1 10 9 13 2
8 9 9 3 9 13 1 11 2
15 15 7 13 1 9 0 9 2 15 15 3 13 3 0 2
11 11 13 0 9 13 15 7 13 0 9 2
23 7 9 13 10 9 9 12 9 1 9 0 9 2 15 13 14 12 0 9 1 0 9 2
22 0 9 0 11 13 1 9 12 3 9 9 7 13 15 9 9 10 9 1 15 9 2
11 9 15 7 13 7 9 9 3 3 13 2
17 3 2 7 11 2 15 13 1 9 1 9 9 0 2 15 13 2
12 11 11 13 0 0 9 9 2 9 7 9 2
10 1 9 12 13 12 9 0 9 9 2
8 4 13 1 0 9 0 9 2
7 0 9 9 13 12 9 2
5 0 9 13 1 9
12 3 4 13 4 13 14 12 9 1 9 1 9
30 0 9 13 3 1 9 16 0 9 9 9 2 3 3 2 16 13 0 13 9 0 9 7 13 9 0 9 1 9 2
24 1 0 9 4 13 13 2 16 4 9 13 13 9 7 9 9 2 3 13 0 9 1 9 2
14 1 9 0 9 13 10 9 9 0 0 9 1 9 2
14 1 10 9 13 1 9 7 9 2 0 7 0 9 2
17 3 9 13 9 1 0 2 0 2 0 7 0 9 0 1 9 2
11 9 9 9 13 7 9 9 7 10 9 2
26 1 9 0 9 11 11 15 1 9 13 10 9 9 0 9 2 15 13 1 9 9 9 0 0 9 2
16 13 15 1 9 0 9 1 9 9 7 9 1 9 0 9 2
15 0 9 13 9 0 9 0 0 9 7 0 0 0 9 2
15 10 9 13 13 1 0 9 7 1 0 9 13 12 9 2
16 1 9 9 9 9 13 1 9 0 12 9 2 13 9 11 2
30 1 10 9 4 13 9 1 9 0 9 13 1 9 9 9 2 12 2 12 1 9 14 12 0 9 7 9 1 9 2
17 1 10 9 11 2 11 13 9 2 16 1 9 9 13 0 9 2
32 13 15 3 3 2 16 1 9 13 1 1 10 9 13 3 0 9 0 9 7 1 9 9 0 9 9 13 3 4 0 13 2
31 0 9 4 3 13 0 9 1 9 9 1 0 9 7 9 2 15 13 10 9 2 7 9 0 15 1 9 9 1 9 2
16 9 1 10 9 13 0 9 7 13 15 13 0 3 1 9 2
5 11 13 0 9 11
2 11 2
12 1 0 9 0 9 11 13 0 0 9 11 2
20 9 3 12 2 2 12 2 9 3 13 0 9 0 0 9 1 9 12 9 2
16 0 9 2 10 9 3 4 13 2 13 9 9 1 12 9 2
13 1 9 0 9 13 9 1 0 9 0 9 9 2
23 11 13 0 9 2 13 13 9 0 9 7 10 9 13 12 9 2 0 9 13 12 9 2
17 1 11 4 9 11 3 13 9 7 9 0 9 1 9 7 9 2
9 13 9 11 4 13 0 0 9 2
19 9 1 12 9 1 9 12 9 2 9 13 1 9 9 12 9 9 0 2
5 9 13 1 9 9
2 11 2
26 9 1 9 3 3 1 11 13 2 16 9 1 0 9 9 0 9 11 11 11 13 1 9 0 9 2
15 0 9 1 0 9 9 4 13 13 0 9 0 0 9 2
31 3 1 9 9 13 1 0 9 1 0 12 0 9 1 12 9 1 12 9 7 1 0 9 1 11 15 10 9 3 13 2
14 9 3 13 1 0 0 9 2 0 9 7 0 9 2
13 9 15 3 1 9 13 3 1 12 9 1 9 2
13 3 3 15 7 13 3 1 9 12 9 1 9 2
5 9 13 9 1 11
2 11 2
17 0 9 9 11 13 1 0 12 9 3 9 9 1 9 0 11 2
17 3 1 9 12 13 9 1 11 12 9 10 9 12 9 9 9 2
11 1 9 12 13 10 9 1 0 12 9 2
10 3 15 10 9 13 1 0 12 9 2
15 1 0 9 9 11 11 4 15 9 1 11 13 3 13 2
20 2 11 7 9 11 13 3 0 3 0 9 1 9 2 2 13 11 2 11 2
32 9 9 0 0 0 9 13 1 11 3 13 3 0 9 1 11 2 3 9 13 1 9 0 0 9 9 1 9 12 9 9 2
12 3 0 9 13 0 12 9 1 10 0 9 2
29 9 0 9 10 9 15 9 13 1 0 9 7 10 9 4 13 0 9 1 9 0 9 1 0 9 7 0 9 2
27 1 12 0 9 2 15 9 13 1 9 12 2 13 3 9 1 9 12 9 9 9 1 9 12 9 9 2
12 9 12 4 1 11 13 13 9 0 9 9 2
20 9 9 13 1 9 0 9 2 15 4 13 9 0 12 9 1 0 0 9 2
13 0 9 9 13 7 1 11 0 1 9 0 9 2
18 12 9 9 9 13 0 7 0 9 2 0 0 0 9 7 11 11 2
17 0 9 13 1 0 9 0 9 1 0 12 9 9 0 12 9 2
33 9 3 13 12 9 9 9 2 1 15 9 13 9 1 0 9 2 12 9 4 13 1 9 0 9 7 12 9 1 9 0 11 2
4 13 12 9 2
6 9 9 3 13 3 9
14 11 13 0 9 9 14 1 12 12 9 1 9 12 9
5 11 2 11 2 2
27 0 9 1 9 2 15 13 1 0 9 16 9 0 9 2 13 10 9 3 1 0 0 9 3 0 9 2
26 13 1 0 0 2 9 2 3 0 9 1 0 9 2 9 2 15 9 13 1 0 9 12 9 9 2
6 9 4 13 12 5 2
23 9 9 13 1 9 9 0 9 11 11 11 0 3 16 9 9 2 15 9 13 3 3 2
6 10 9 13 3 13 2
26 9 15 7 9 13 1 0 0 9 2 7 2 3 2 1 9 1 9 7 1 9 0 9 1 9 2
12 1 9 0 2 9 13 11 7 9 0 9 2
25 9 13 13 10 9 14 1 9 0 0 9 2 3 7 1 9 12 9 7 1 9 0 9 9 2
28 0 9 4 13 12 5 3 2 0 9 1 9 1 9 7 0 2 3 0 9 1 0 9 13 12 5 3 2
12 9 1 9 7 11 13 3 0 9 0 9 2
82 9 0 0 9 2 1 15 13 0 13 0 9 9 9 2 3 9 2 9 1 9 9 7 9 2 0 9 2 9 1 9 2 9 3 2 13 1 12 0 0 9 2 0 9 2 0 9 2 0 7 0 9 2 7 9 0 7 0 9 2 3 9 11 2 0 9 2 0 9 11 2 11 2 0 9 2 0 9 2 11 0 2
11 9 15 13 1 9 1 12 1 12 5 2
7 9 9 13 13 1 0 9
2 11 2
15 0 9 13 1 12 2 9 0 0 9 1 9 0 9 2
19 13 1 0 9 1 12 2 12 2 12 7 12 9 0 12 7 12 5 2
7 0 9 13 12 12 9 2
12 0 9 1 0 9 9 13 3 7 0 9 2
48 16 11 13 9 0 9 9 11 11 2 0 9 1 9 9 13 2 16 13 13 9 1 10 9 14 1 9 10 0 9 7 1 0 9 10 9 2 3 1 12 2 12 2 12 7 12 9 2
33 2 16 13 9 1 0 0 9 3 12 9 12 9 2 13 10 9 13 14 1 10 9 7 1 9 12 9 2 2 13 11 11 2
6 9 13 12 5 3 2
15 9 13 2 16 4 13 9 9 3 13 7 9 1 9 2
36 2 0 2 9 9 2 15 0 9 1 9 13 2 13 10 9 13 9 1 3 12 12 9 2 16 0 9 13 0 13 1 10 9 0 9 2
35 9 13 2 3 7 1 0 9 2 13 7 9 2 16 9 0 0 9 2 15 15 9 15 13 2 4 1 0 9 13 1 0 9 3 2
28 1 10 9 13 9 9 2 15 13 13 1 3 0 0 9 2 13 3 15 2 7 15 1 3 0 0 9 2
6 11 15 13 1 11 11
2 11 2
23 9 11 2 15 13 9 11 11 7 0 11 2 15 4 13 1 12 0 9 1 11 11 2
10 13 15 3 9 11 1 11 11 11 2
18 0 9 1 3 0 9 4 13 0 0 9 7 0 9 4 13 11 2
12 11 13 1 0 9 13 0 9 11 2 11 2
22 0 9 13 0 9 1 0 2 0 7 0 9 3 9 0 9 1 9 11 7 11 2
13 9 11 13 0 9 2 15 13 1 11 0 9 2
17 0 11 13 9 0 9 2 16 10 0 9 13 3 12 9 9 2
5 12 9 1 0 9
2 11 2
14 3 3 12 9 13 9 9 2 15 13 9 0 9 2
9 13 15 3 9 9 9 11 11 2
31 1 10 9 13 13 13 0 2 15 15 13 13 9 0 9 0 9 2 15 13 9 9 7 13 1 10 9 10 10 9 2
17 2 4 15 13 10 9 13 7 9 9 2 15 1 15 13 9 2
28 0 9 13 13 9 1 9 7 9 2 16 4 13 9 2 15 1 0 9 9 13 0 9 2 2 13 11 2
17 1 10 9 13 9 9 3 0 2 16 9 9 15 9 0 13 2
27 9 0 9 2 15 13 3 1 9 2 13 13 3 0 0 9 2 7 15 13 7 9 2 7 10 9 2
10 13 1 10 9 0 0 9 0 9 2
20 16 11 13 11 11 2 3 13 9 12 9 2 0 12 9 13 1 9 9 2
5 11 13 1 9 9
2 11 2
18 0 9 13 1 9 9 0 9 9 1 0 9 7 1 9 9 11 2
19 1 9 9 9 11 7 0 9 11 15 13 0 0 9 11 11 2 11 2
20 1 9 9 2 15 0 9 13 13 9 9 2 4 13 9 0 3 1 11 2
20 1 9 15 15 7 1 9 13 14 10 10 9 2 15 13 1 0 9 13 2
26 9 11 2 10 9 13 3 13 1 9 0 9 2 13 12 2 7 12 2 9 1 11 9 0 9 2
16 13 15 3 9 9 13 1 9 2 15 13 1 9 9 0 2
5 9 1 0 9 13
2 11 2
31 0 9 13 1 0 9 12 2 9 9 9 11 2 9 7 0 9 1 9 1 12 9 2 15 13 3 12 9 1 9 2
11 13 1 15 3 9 11 11 1 0 9 2
23 0 9 9 13 1 10 9 9 0 9 15 9 2 15 0 9 13 2 3 1 12 9 2
26 9 11 13 3 3 0 9 7 1 9 0 0 9 7 9 10 9 9 13 3 1 12 9 1 9 2
1 3
29 11 4 13 9 1 9 12 9 2 9 2 15 4 13 0 9 1 9 10 9 1 9 9 1 0 0 2 9 2
6 9 9 1 9 13 3
11 11 3 3 13 1 0 9 12 9 9 2
5 9 11 4 13 2
5 11 7 11 13 15
1 9
33 1 9 9 9 13 1 9 0 9 9 11 1 0 9 3 12 9 9 2 1 15 12 9 2 9 4 1 9 13 1 0 9 2
30 16 13 1 9 0 0 9 2 1 9 11 7 11 9 9 0 9 2 15 4 13 1 10 9 3 0 9 2 13 2
7 0 9 11 13 0 9 2
53 1 10 9 1 11 2 15 13 3 12 9 2 9 7 13 3 9 0 9 1 9 12 7 12 1 0 9 12 9 2 9 2 13 0 0 9 2 15 11 13 1 9 12 2 3 1 0 9 12 9 2 9 2
41 1 9 1 9 9 1 11 7 0 9 1 9 0 9 13 11 0 9 13 1 9 12 7 0 9 2 3 12 9 2 9 2 1 9 12 7 12 1 9 12 2
46 1 0 9 11 13 11 0 12 9 9 1 0 2 0 9 2 15 13 1 9 9 9 0 9 9 0 9 1 9 12 2 7 3 0 9 12 9 9 2 1 15 3 13 12 9 2
50 9 0 9 1 9 0 7 0 9 2 15 1 9 1 9 9 11 13 13 14 1 9 12 2 7 0 2 0 9 2 15 13 0 3 1 9 12 2 13 1 0 9 13 1 2 0 2 0 9 2
24 9 2 15 13 1 0 2 0 9 1 9 0 9 2 11 1 9 12 1 9 13 9 9 2
28 0 9 9 9 2 15 9 11 3 13 1 12 7 12 9 9 3 2 4 13 3 2 0 13 1 9 12 2
27 16 13 1 9 9 9 7 11 2 9 9 0 9 1 9 13 9 0 0 9 2 3 13 9 0 9 2
37 15 13 9 10 0 9 2 15 4 1 9 12 3 13 16 9 0 0 9 2 7 0 9 1 9 11 2 7 3 0 0 0 9 11 1 9 2
19 1 9 11 0 2 3 2 0 0 9 3 1 9 12 0 0 9 13 2
14 1 0 9 10 9 13 0 9 9 0 1 9 12 2
13 10 9 3 11 13 3 1 11 12 9 2 9 2
16 9 1 9 0 9 11 4 1 9 9 9 1 0 9 13 2
28 1 9 2 15 13 11 1 9 2 15 1 0 9 2 15 4 1 9 13 1 0 9 2 3 13 0 9 2
18 3 1 10 0 9 13 12 9 2 9 11 2 3 13 10 9 11 2
15 1 9 1 9 11 9 1 9 9 3 13 11 7 11 2
35 9 11 2 15 13 9 1 9 1 0 9 11 2 13 2 16 9 10 9 13 1 0 0 9 0 9 7 10 0 0 9 13 3 0 2
25 1 9 11 13 3 0 9 1 11 12 9 9 2 1 11 12 9 9 7 1 11 12 9 9 2
33 1 9 2 15 13 0 11 1 0 9 2 13 12 9 9 9 11 2 12 9 11 2 12 9 11 7 12 9 9 11 7 11 2
25 0 9 1 0 9 2 15 13 1 9 0 0 9 2 13 1 0 9 3 0 16 0 0 9 2
30 16 13 1 9 9 9 7 0 0 9 2 13 9 0 0 9 1 9 14 3 3 2 15 1 15 13 3 3 13 2
18 9 11 11 1 0 9 11 2 12 2 3 1 9 13 9 9 11 11
5 9 9 13 13 9
13 9 13 9 1 9 7 4 9 13 7 1 0 9
27 0 9 9 9 2 9 9 2 2 15 13 13 1 0 9 1 0 0 9 2 13 3 13 9 0 9 2
17 11 15 13 11 11 1 9 9 9 11 2 15 15 13 9 9 2
19 9 0 9 13 0 9 2 1 15 4 0 9 1 9 0 9 13 9 2
12 15 2 16 13 9 9 2 13 13 9 9 2
20 9 7 9 9 2 15 15 4 0 9 13 2 4 13 9 7 13 1 9 2
25 11 15 13 2 16 16 15 9 13 1 0 9 9 2 13 9 9 1 9 13 0 7 0 9 2
26 3 13 2 16 1 9 0 9 1 0 9 2 15 9 9 13 2 13 0 9 0 0 7 0 9 2
8 10 9 13 3 9 9 9 2
6 9 13 3 0 9 2
19 1 9 9 2 12 1 0 9 13 3 13 9 2 15 13 9 13 9 2
17 2 13 10 9 2 16 9 9 1 15 13 13 2 2 13 11 2
21 9 9 9 11 11 0 9 13 2 16 9 9 4 13 1 9 9 1 0 9 2
15 1 9 14 13 1 0 9 2 15 13 1 0 9 13 2
15 2 7 3 4 13 0 9 1 10 9 7 9 1 9 2
12 3 15 13 0 1 9 9 2 2 13 11 2
35 1 10 9 13 13 1 9 9 9 2 16 15 4 13 1 9 1 9 2 1 9 1 0 9 2 9 7 3 7 1 0 7 0 9 2
44 1 9 2 16 15 13 2 16 4 15 15 13 9 9 0 9 13 1 9 9 2 11 13 2 16 9 1 9 2 9 9 2 13 0 2 13 12 12 9 7 13 14 0 2
5 0 9 0 9 2
2 11 2
14 0 9 9 13 3 0 9 0 9 7 1 0 9 2
17 16 0 9 1 15 10 13 2 13 15 9 3 12 12 12 9 2
29 0 9 4 1 0 9 13 3 2 16 13 3 3 16 9 12 9 2 7 16 9 15 2 15 13 2 13 0 2
12 9 2 15 4 13 0 0 9 2 15 13 2
17 12 10 0 9 2 1 15 15 9 13 2 15 1 9 9 13 2
6 0 9 13 1 11 9
2 11 2
12 0 9 4 1 9 1 0 9 13 11 11 2
22 1 0 9 9 11 11 11 3 0 9 13 1 9 9 1 9 9 1 9 11 11 2
29 0 9 11 11 11 1 0 9 13 9 9 10 9 2 15 15 13 12 2 9 1 9 9 11 1 0 9 11 2
14 11 3 9 1 9 13 7 13 9 13 1 0 9 2
29 16 4 3 13 2 9 11 13 9 1 9 2 15 15 13 9 2 9 2 0 9 7 9 0 9 1 9 11 2
36 11 1 9 13 9 2 16 1 9 9 13 13 7 0 0 9 0 9 2 3 16 9 0 0 9 1 9 9 9 0 1 0 9 3 13 2
19 11 13 2 16 15 9 4 13 7 1 0 9 2 7 0 0 9 11 2
4 9 13 1 9
4 11 1 9 2
27 1 12 9 2 15 15 9 1 9 11 11 13 1 0 9 2 15 3 9 0 9 11 11 13 1 9 2
18 0 9 9 9 11 13 1 9 10 9 9 0 9 1 11 1 9 2
19 3 9 0 9 11 13 2 16 13 13 1 0 0 9 1 9 0 9 2
14 11 11 13 2 16 13 9 0 9 9 9 7 9 2
18 13 3 9 9 9 2 3 2 9 9 1 9 7 0 9 0 9 2
18 9 13 1 9 9 0 1 9 0 9 2 9 7 1 3 0 9 2
12 2 13 15 7 9 1 0 9 15 1 9 2
19 3 0 13 9 1 9 1 9 2 1 15 15 9 13 2 2 13 9 2
4 9 13 0 11
2 11 2
19 13 0 9 2 9 2 3 0 0 9 0 11 13 7 3 9 0 9 2
9 13 1 15 1 10 0 0 9 2
21 1 3 16 0 9 9 13 9 2 1 15 15 13 1 9 9 1 12 2 9 2
23 15 3 13 0 0 9 9 0 9 2 11 2 13 9 0 11 1 0 11 1 0 11 2
24 9 3 13 2 16 4 15 9 13 3 1 9 1 0 11 1 11 7 13 0 9 0 11 2
18 0 9 13 0 9 11 11 2 0 15 1 9 9 1 9 12 9 2
32 11 13 2 16 4 15 1 11 13 3 12 0 9 2 0 0 9 15 3 13 0 9 7 0 11 1 11 13 14 1 9 2
4 13 15 0 9
13 0 0 9 13 3 1 12 9 11 11 2 11 11
4 11 2 11 2
20 0 9 15 13 1 0 12 9 0 9 7 3 1 9 13 9 1 9 0 2
21 0 9 9 11 11 13 1 0 0 9 12 2 9 1 12 0 9 2 0 11 2
20 3 0 9 15 1 9 1 11 13 0 9 2 15 4 13 9 0 0 9 2
25 1 10 9 13 0 9 16 0 9 2 12 0 9 3 2 15 4 13 9 2 2 7 0 9 2
37 12 9 13 9 0 9 2 11 11 2 11 7 11 2 11 11 2 11 2 0 9 14 13 7 11 1 11 2 1 0 9 3 13 13 9 11 2
23 9 11 11 1 15 13 2 16 13 0 9 7 1 10 9 13 11 0 9 2 16 13 2
36 1 0 9 10 9 13 7 3 13 10 9 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2
17 13 15 2 16 13 12 9 2 14 1 9 13 12 1 0 9 2
22 2 11 13 0 2 14 13 2 16 13 1 0 9 0 13 0 9 2 2 13 11 2
16 2 13 14 9 2 16 4 15 9 13 14 1 3 0 9 2
16 11 13 9 1 9 0 11 7 1 9 13 0 13 7 11 2
38 3 15 3 3 1 10 9 13 2 0 1 9 4 13 3 2 16 4 3 13 2 2 13 12 0 9 11 2 15 13 3 7 9 0 9 11 11 2
14 7 9 11 13 2 16 0 9 13 0 9 1 9 2
21 2 13 4 15 2 16 4 10 9 13 9 2 15 13 0 2 16 4 13 9 2
19 13 13 2 10 9 15 13 2 15 15 13 1 9 9 2 2 13 11 2
4 0 9 13 0
3 12 9 11
2 11 2
10 1 9 13 1 11 9 14 0 9 2
31 1 9 1 11 2 12 2 12 2 3 13 0 0 9 11 11 2 15 1 12 2 1 12 2 9 13 9 11 12 9 2
23 11 15 1 10 0 9 2 15 13 9 0 0 9 2 13 2 2 13 15 3 12 9 2
11 13 3 3 15 2 15 3 13 13 2 2
4 11 13 3 9
8 11 11 15 13 9 1 0 9
2 11 2
30 2 1 9 1 11 13 13 0 9 2 13 3 9 7 14 9 2 2 13 15 0 0 9 0 11 10 9 11 11 2
15 0 13 1 0 9 3 1 9 14 1 12 2 9 9 2
18 3 15 13 2 16 9 13 0 9 11 2 11 2 7 3 12 13 2
39 2 9 13 0 13 7 13 0 2 16 4 13 0 9 11 7 0 9 11 2 2 13 10 9 9 11 11 7 13 1 9 9 2 2 13 4 12 9 2
8 3 9 4 13 1 9 9 2
12 13 13 1 9 7 3 13 0 0 9 2 2
20 11 13 1 0 11 11 2 3 9 13 9 11 2 15 4 1 9 9 13 2
16 0 9 11 15 13 13 0 9 2 15 13 9 1 0 11 2
41 2 1 10 9 15 13 0 7 0 9 2 2 13 1 9 11 7 13 2 2 15 0 4 13 13 9 2 7 11 13 3 7 3 11 13 9 1 9 9 2 2
25 13 2 11 2 0 2 11 2 2 11 2 0 2 11 2 2 11 2 1 9 1 11 11 2 2
37 13 2 11 2 11 2 2 11 2 0 2 11 2 2 11 2 9 1 11 2 2 9 2 9 1 11 2 2 11 2 11 2 9 1 11 2 2
3 9 9 9
10 13 2 14 1 11 9 2 13 0 9
2 11 2
20 13 15 0 9 13 9 11 11 1 0 9 2 3 9 13 12 2 9 9 2
25 2 9 13 13 9 7 9 2 15 15 15 9 11 2 11 7 11 13 2 2 13 9 11 11 2
18 10 9 13 1 9 2 3 13 2 9 2 13 1 0 9 12 9 2
9 2 9 13 9 7 9 9 9 2
14 16 15 15 13 2 13 9 10 9 13 3 1 9 2
22 13 4 1 15 7 9 2 16 10 9 13 1 9 14 1 9 2 3 13 0 9 2
14 3 4 1 11 13 0 9 2 2 13 9 11 11 2
22 3 9 13 1 0 9 2 1 9 2 12 9 9 2 16 12 9 9 13 9 11 2
9 3 15 13 1 9 11 1 11 2
17 2 13 9 2 16 4 15 13 1 15 2 16 1 15 13 11 2
19 16 13 1 15 2 1 9 15 13 2 3 15 15 13 2 2 13 11 2
25 2 9 2 14 13 11 1 2 9 2 13 2 4 15 3 7 13 7 10 9 13 1 9 13 2
24 13 2 11 2 9 1 11 2 2 11 2 9 1 11 2 2 11 2 9 1 11 11 2 2
32 13 2 11 2 11 11 2 2 11 2 11 2 11 2 9 1 11 11 2 2 11 2 11 2 2 11 2 9 1 11 2 2
6 1 0 9 13 3 9
7 0 11 13 0 9 1 9
3 0 11 2
17 1 0 9 9 0 2 11 13 2 3 13 1 0 9 1 9 2
23 9 3 15 13 2 9 11 2 11 7 11 13 2 16 1 9 9 15 13 3 0 9 2
16 9 13 11 3 2 9 13 1 12 9 1 11 7 1 11 2
31 0 9 13 3 0 2 0 2 11 13 1 9 0 2 11 11 1 11 7 3 1 0 0 9 1 9 13 1 11 11 2
9 3 15 9 11 13 1 9 3 2
10 0 13 1 9 11 7 3 13 9 2
16 9 1 9 13 13 15 9 1 9 7 13 1 9 1 9 2
12 2 1 9 9 13 3 13 2 15 13 0 2
10 0 9 15 7 13 1 9 1 9 2
16 0 9 13 9 11 9 2 1 9 9 15 13 9 7 9 2
11 13 15 0 9 2 2 13 9 9 11 2
27 0 9 0 2 11 2 12 2 9 2 12 9 2 12 9 2 12 9 2 9 12 2 12 2 12 9 2
61 13 2 11 2 0 2 11 2 2 11 2 11 11 2 2 11 7 11 2 1 9 9 2 2 11 2 11 2 2 11 2 9 1 11 13 1 9 2 2 11 2 11 2 1 9 2 2 11 2 1 9 2 2 11 2 13 9 1 11 2 2
26 13 2 11 2 11 2 11 2 11 2 2 11 2 11 2 9 2 2 11 2 9 9 1 11 2 2
4 9 1 11 13
8 1 0 9 15 1 11 3 13
2 11 2
18 1 0 0 9 3 0 0 9 13 9 9 11 11 11 9 0 9 2
24 0 9 0 9 13 11 7 11 2 3 3 13 11 2 15 13 1 11 16 0 9 0 9 2
26 1 9 15 3 13 9 11 2 15 4 1 9 11 13 11 9 2 7 12 0 9 1 9 2 9 2
26 9 11 1 9 13 0 1 10 0 9 1 9 2 13 15 1 0 9 9 7 13 1 12 9 9 2
12 1 0 0 9 9 7 15 10 9 3 13 2
8 2 16 13 10 9 9 9 2
12 15 13 14 9 2 2 13 3 3 9 11 2
15 1 0 9 9 7 9 13 2 2 10 9 13 14 0 2
18 7 15 13 9 2 15 15 13 0 9 2 13 9 13 7 13 2 2
23 9 1 11 13 1 0 9 2 1 12 1 12 9 2 2 14 1 0 9 13 0 9 2
30 16 1 9 11 13 11 16 0 9 2 13 9 9 11 11 1 15 2 16 4 0 0 9 13 13 9 1 9 9 2
17 3 13 15 13 1 0 9 2 2 9 14 15 1 11 15 13 2
13 13 1 9 2 13 4 2 16 15 13 0 9 2
8 13 15 1 0 9 11 2 2
25 0 9 11 2 12 2 9 2 12 9 2 12 9 2 12 9 2 9 12 2 12 2 12 9 2
30 13 2 11 2 1 9 1 0 2 11 2 2 11 2 11 2 2 11 2 11 2 11 2 13 1 9 2 9 2 2
37 13 2 11 2 1 9 9 1 11 2 2 11 2 13 9 1 11 2 2 11 2 1 9 9 3 1 11 2 2 11 2 1 9 1 11 2 2
3 0 9 9
7 1 0 9 3 7 0 9
2 11 2
25 3 13 4 13 9 1 0 15 9 1 0 9 1 0 11 2 12 2 2 12 2 12 2 2 2
21 1 9 0 9 7 13 1 0 9 0 9 7 13 15 16 3 4 1 0 9 2
24 0 9 9 1 0 9 9 3 9 13 2 7 0 0 9 0 9 15 3 14 15 13 13 2
22 11 11 13 1 0 9 1 0 9 9 11 2 11 2 11 2 11 2 11 7 11 2
27 9 11 11 13 9 13 1 15 9 1 9 1 9 9 2 3 12 9 7 12 9 2 7 3 13 9 2
15 10 0 9 15 1 1 0 0 9 9 13 13 14 3 2
9 0 9 11 1 0 9 13 13 2
9 11 13 13 1 9 7 12 9 2
13 13 15 4 3 1 9 9 11 1 9 1 11 2
31 16 4 15 9 1 0 9 13 1 12 2 9 2 13 4 15 0 9 1 12 9 7 9 1 9 1 9 12 1 11 2
14 1 0 9 11 13 2 2 11 15 13 3 0 9 2
20 16 13 1 9 2 1 15 4 3 13 2 7 1 9 9 4 15 15 13 2
8 1 9 13 15 0 0 2 2
11 14 16 7 11 13 9 1 9 1 9 2
15 2 9 13 12 9 7 9 0 2 2 13 0 9 11 2
24 11 11 4 13 1 0 9 9 10 9 1 0 9 1 12 2 9 2 1 9 3 1 0 2
17 1 9 11 2 11 2 11 2 11 2 11 2 11 12 9 13 2
10 3 15 13 15 1 12 3 0 9 2
16 9 0 9 4 13 0 11 2 11 2 11 2 11 7 11 2
15 0 9 13 11 1 11 2 9 4 0 13 0 0 9 2
4 0 9 1 11
2 11 2
13 0 0 9 1 0 9 9 13 0 0 9 11 2
28 15 15 10 0 9 12 9 7 0 9 12 9 12 13 1 9 9 11 11 1 0 9 11 0 0 0 9 2
8 0 9 13 1 0 9 9 2
39 15 3 1 0 9 0 9 9 1 9 2 0 12 9 1 9 2 9 7 9 1 9 2 13 3 1 0 9 1 0 9 2 16 13 0 1 0 9 2
21 1 9 3 0 9 3 3 13 12 9 2 9 7 9 2 1 15 13 15 9 2
4 0 9 1 9
12 9 12 2 9 0 9 13 9 0 9 1 11
2 11 2
45 16 0 12 9 9 0 9 2 11 2 13 1 0 9 12 2 9 13 3 1 9 9 1 9 1 9 14 7 0 11 1 0 11 3 14 1 9 2 3 12 9 13 1 3 2
13 9 11 2 11 13 0 7 9 4 3 13 9 2
18 11 15 1 9 13 9 9 1 11 7 1 11 1 9 9 13 13 2
28 7 11 4 13 13 0 11 2 3 1 11 7 11 2 2 16 9 9 4 15 15 1 0 9 9 13 13 2
14 11 13 1 0 9 1 11 0 9 11 7 9 11 2
15 12 1 0 9 13 7 1 0 9 15 13 14 1 9 2
11 1 9 9 1 12 9 15 13 9 11 2
25 11 13 1 0 9 9 1 0 9 16 1 9 1 11 2 13 4 9 11 2 15 13 0 9 2
7 11 4 13 9 1 9 2
15 11 13 9 1 9 2 11 13 9 9 7 11 3 9 2
23 9 11 11 11 1 9 13 2 2 9 1 0 11 13 0 1 9 1 9 1 9 14 2
23 11 4 13 9 0 9 2 7 16 13 13 1 9 1 0 9 2 13 13 3 9 2 2
8 0 9 1 9 11 9 9 9
2 11 2
19 0 9 1 9 2 0 0 9 11 11 2 13 9 7 13 9 9 9 2
37 0 9 2 15 0 1 9 13 15 0 9 10 9 1 12 0 9 1 15 7 3 15 13 3 9 9 2 4 13 1 0 9 1 9 15 9 2
11 1 12 9 13 0 9 7 13 15 9 2
17 1 10 9 13 13 9 1 0 9 9 11 2 12 2 12 2 2
13 9 1 0 9 13 1 9 9 11 11 2 11 2
27 3 3 1 9 1 0 9 9 1 0 11 11 13 2 15 15 3 3 13 2 16 13 1 10 9 9 2
12 0 9 15 1 11 13 13 3 1 0 9 2
21 1 12 9 15 4 3 13 2 16 15 13 1 9 2 15 15 3 3 3 13 2
21 1 0 9 11 13 2 16 1 10 0 9 15 13 12 9 1 9 12 1 11 2
14 1 0 9 3 13 0 9 9 1 9 7 13 15 2
8 1 9 15 1 9 13 9 2
14 1 10 9 7 13 9 0 0 9 2 15 15 13 2
12 13 15 14 2 16 9 0 1 9 9 13 2
28 2 13 4 7 0 9 2 1 9 9 4 15 3 14 13 2 16 4 15 15 1 15 13 2 2 13 11 2
31 0 0 9 2 9 11 11 2 7 3 9 13 2 16 9 9 15 3 10 9 13 2 16 1 0 9 15 15 13 13 2
19 11 11 15 13 12 2 9 12 9 2 1 15 0 13 3 3 12 9 2
13 9 13 1 9 11 1 0 9 2 9 13 11 2
15 9 4 1 12 9 13 7 13 1 9 0 11 1 11 2
22 1 0 9 9 13 10 9 1 10 9 2 3 13 9 2 15 15 13 9 1 9 2
21 3 15 13 9 2 9 7 9 2 0 9 1 9 15 7 13 1 10 9 13 2
32 3 1 9 9 11 11 2 0 0 9 2 15 13 11 1 9 0 9 2 1 11 13 9 2 12 10 0 0 9 2 0 2
6 3 15 13 12 9 2
22 1 0 11 13 0 1 9 9 12 9 1 9 1 12 0 9 2 13 3 12 9 2
1 3
25 0 0 0 9 11 2 11 13 0 9 2 3 0 1 0 9 1 0 0 9 1 11 1 11 2
5 9 11 15 13 9
2 11 2
16 9 0 9 11 11 11 11 15 13 10 9 1 0 9 11 2
40 2 13 1 0 9 2 16 4 1 0 9 13 1 9 0 9 1 11 7 9 0 9 9 11 10 9 3 13 1 9 2 2 13 11 1 9 1 10 9 2
54 11 13 13 1 9 12 2 9 1 11 2 1 9 7 9 13 12 10 9 1 0 9 1 0 9 1 11 2 2 9 2 2 3 2 11 2 9 1 12 9 2 7 3 1 9 13 0 1 9 0 9 1 11 2
7 15 13 11 13 1 9 2
21 2 11 13 10 9 2 1 0 9 1 11 4 13 3 7 3 15 1 15 13 2
15 13 3 1 0 9 7 13 15 15 13 2 2 13 11 2
18 13 1 10 9 2 16 0 9 9 15 13 11 11 2 3 9 11 2
4 0 9 1 9
7 0 9 13 12 9 1 11
2 11 2
30 0 9 0 9 0 9 13 0 9 11 7 13 10 9 1 9 9 1 9 1 0 11 2 15 15 13 12 2 9 2
22 0 9 9 1 12 0 9 3 13 1 0 9 1 12 9 1 12 2 9 0 9 2
15 1 0 9 9 0 9 15 13 9 0 0 9 1 11 2
12 2 3 13 9 2 2 13 9 9 11 11 2
14 0 13 9 9 2 9 7 0 9 0 9 2 9 2
7 15 13 1 0 9 0 2
24 13 15 13 9 0 1 0 3 2 1 0 9 4 15 3 13 9 1 0 9 9 1 0 2
17 13 4 9 14 2 1 10 12 2 9 4 13 0 12 9 9 2
16 0 9 9 14 15 13 1 12 2 15 0 1 12 0 9 2
15 9 2 15 13 0 9 1 9 2 3 13 3 12 9 2
3 1 0 9
29 9 11 1 11 15 13 1 0 9 1 0 11 2 15 13 12 2 12 2 9 7 10 9 1 0 9 13 13 2
16 0 9 11 15 1 9 9 13 9 9 11 1 11 1 11 2
17 15 1 0 9 3 4 13 0 9 2 7 9 15 13 1 9 2
28 0 9 13 9 11 11 11 2 11 2 15 4 13 1 9 1 9 9 11 11 2 11 1 9 12 2 12 2
5 11 3 1 9 2
2 11 2
25 1 9 1 0 9 0 9 9 1 9 1 11 13 1 12 2 9 11 11 9 9 9 12 9 2
20 0 9 15 13 2 11 15 3 13 9 2 16 13 12 2 7 12 2 9 2
11 1 12 2 9 13 11 0 9 1 11 2
9 1 9 9 13 3 14 10 0 9
7 1 9 11 11 2 0 9
33 1 0 9 15 1 9 0 9 7 9 2 15 13 0 9 1 9 2 13 3 0 9 16 9 9 2 11 2 9 9 7 0 2
23 15 3 3 3 13 2 16 0 0 9 13 1 15 2 15 15 1 15 13 1 9 9 2
20 1 9 3 13 0 9 1 9 0 9 2 15 15 13 1 11 1 9 12 2
16 1 10 9 13 9 1 0 9 1 3 0 9 0 0 9 2
14 9 0 9 15 1 0 0 9 13 0 9 1 9 2
39 1 15 4 13 3 0 0 9 11 11 2 15 9 9 1 12 9 1 0 9 13 0 9 2 0 9 2 7 3 7 9 1 3 0 7 0 0 9 2
17 15 2 16 3 15 13 9 2 13 1 0 9 9 1 0 9 2
12 9 9 1 9 0 9 13 7 13 15 0 2
23 3 15 3 15 13 1 0 9 10 9 0 0 9 1 0 9 11 2 15 13 1 9 2
11 12 1 15 4 1 10 9 13 1 9 2
11 13 2 16 4 15 1 15 13 3 3 2
34 1 9 9 9 9 11 4 15 13 2 16 0 9 15 1 9 9 13 3 2 16 1 10 9 13 1 9 9 2 14 7 1 9 2
10 7 9 1 15 2 15 1 9 13 2
14 3 3 2 9 13 9 3 0 9 13 3 1 9 2
17 9 9 9 4 1 9 9 13 13 7 9 0 9 1 10 0 2
12 13 4 13 0 7 0 1 9 1 0 9 2
12 9 0 15 13 9 9 0 9 13 3 0 2
12 3 15 13 3 0 9 1 0 9 1 9 2
15 3 15 2 15 13 14 0 9 2 7 7 0 0 9 2
8 7 13 15 7 0 0 9 2
51 15 1 15 15 1 9 9 13 2 16 4 15 13 13 3 3 3 2 7 10 9 2 14 9 7 0 9 1 15 2 15 13 0 0 9 2 15 3 13 2 16 13 0 9 2 13 7 13 0 9 2
8 3 15 3 13 1 9 9 2
6 0 0 9 2 2 2
8 2 11 12 2 12 2 12 2
12 13 0 13 2 16 13 0 9 3 9 0 2
13 3 13 9 1 15 0 9 2 15 13 9 0 2
16 13 9 2 16 9 9 1 9 13 1 9 1 0 0 9 2
14 0 9 3 13 0 9 0 0 9 7 3 9 0 2
21 16 0 9 13 1 9 0 9 2 13 0 2 16 4 15 13 1 9 10 9 2
18 0 9 13 0 0 9 7 1 10 9 4 13 7 9 9 0 9 2
17 13 1 0 13 9 9 0 9 2 15 13 9 1 0 7 0 2
29 13 15 3 9 2 15 0 9 2 9 2 0 9 7 9 13 0 0 9 0 1 9 2 15 9 0 9 13 2
14 0 9 13 10 0 9 2 15 4 13 13 1 9 2
6 9 1 0 9 13 2
15 7 4 9 13 3 10 9 0 9 13 16 9 1 9 2
32 7 16 9 13 9 2 1 10 9 3 0 0 9 2 9 9 1 0 9 7 0 9 0 1 9 9 9 2 15 13 0 2
20 13 9 3 0 2 16 4 13 13 9 7 0 9 0 9 16 9 9 9 2
18 13 3 3 9 9 9 1 9 2 15 15 13 0 9 1 9 9 2
21 3 15 3 13 7 1 10 9 2 16 13 0 0 9 2 15 13 16 0 9 2
1 3
20 0 9 7 9 11 11 13 1 9 0 9 12 2 12 2 1 0 9 11 2
5 9 1 12 9 2
18 0 9 0 0 11 15 13 1 9 12 2 9 1 0 0 9 9 2
7 16 9 15 13 9 11 2
5 9 0 9 12 2
8 1 10 9 13 9 2 11 11
25 3 15 13 1 15 2 15 13 9 9 0 9 1 0 9 1 0 9 9 0 9 1 0 9 2
7 15 9 9 1 9 13 2
26 13 15 0 0 9 2 15 13 0 13 1 9 0 0 9 9 11 2 7 1 9 0 7 0 2 2
25 1 9 9 15 0 7 0 9 13 0 9 9 11 1 9 9 9 2 15 1 10 9 3 13 2
8 9 13 4 13 9 0 9 2
15 13 3 1 0 9 9 11 2 15 15 3 13 9 9 2
34 9 15 13 13 15 2 16 4 4 13 9 9 0 9 7 0 9 13 13 13 15 9 9 1 15 9 2 1 15 13 9 1 9 2
46 13 2 14 9 2 16 9 9 7 9 13 1 9 1 9 7 16 0 9 13 3 0 9 9 10 9 2 9 3 1 9 13 13 0 9 0 9 2 1 0 9 0 0 9 2 2
57 9 12 0 9 13 2 16 9 9 0 15 1 0 1 9 9 9 0 9 13 13 9 9 0 9 1 0 9 3 14 1 9 15 0 0 9 9 1 3 0 9 0 9 7 1 9 12 9 1 9 2 3 4 13 0 9 2
29 3 9 12 9 2 12 13 0 9 1 0 9 13 0 9 1 0 3 2 13 2 14 15 1 0 1 9 12 2
16 9 12 13 3 12 0 9 2 15 13 9 0 9 3 13 2
17 3 13 13 15 0 0 9 9 2 15 13 13 0 7 0 2 2
20 1 15 2 10 0 9 9 13 0 1 0 9 3 13 2 13 13 0 9 2
7 0 13 14 9 0 9 2
27 3 13 13 2 16 13 13 13 15 1 9 1 9 0 0 9 2 0 3 16 9 2 9 3 2 2 2
27 9 1 9 12 13 2 16 1 9 2 16 13 1 9 12 9 9 9 2 13 4 13 14 1 0 9 2
31 13 2 14 0 9 1 9 3 0 0 9 9 2 13 13 3 15 1 15 2 1 15 15 13 3 13 2 16 13 0 2
32 9 12 13 3 1 10 9 0 13 3 2 16 4 13 0 0 9 9 10 9 1 9 13 15 0 9 9 7 9 0 9 2
18 9 0 9 7 13 13 2 3 13 3 0 0 9 7 1 10 9 2
37 1 1 15 2 16 0 9 7 9 13 1 15 1 9 0 9 2 13 3 0 13 7 0 9 1 9 12 9 2 12 9 2 9 2 9 11 2
24 3 7 3 13 0 13 2 16 13 0 1 9 9 0 9 1 0 9 13 3 3 0 9 2
4 9 2 0 9
18 9 9 11 13 2 2 0 2 13 9 7 13 15 9 1 10 9 2
18 13 4 15 16 9 2 13 9 7 0 9 2 16 4 15 13 9 2
31 3 10 9 13 0 13 1 10 9 2 3 15 13 9 2 15 15 9 13 2 13 13 9 7 13 15 9 2 2 2 2
8 9 13 9 0 9 0 9 2
19 16 15 13 1 9 9 2 13 15 0 9 1 0 9 0 1 0 9 2
33 1 9 9 2 15 13 3 3 1 12 2 15 1 0 4 13 3 10 9 3 13 7 16 15 9 1 10 9 13 13 0 9 2
23 1 9 2 10 1 10 9 13 9 2 11 11 1 0 9 1 11 2 13 9 0 11 2
3 9 7 9
1 9
31 0 9 7 9 11 11 2 12 2 15 1 0 9 13 16 0 9 3 15 2 13 15 2 0 9 2 3 7 3 2 2
13 1 10 9 13 0 9 9 10 9 1 0 9 2
26 1 0 9 2 13 15 9 11 1 12 9 2 2 15 9 13 9 2 1 10 9 3 0 2 9 2
15 1 0 2 9 2 15 13 3 12 9 2 9 7 9 2
26 0 9 13 0 2 9 13 13 9 10 2 9 2 1 9 9 7 13 15 13 10 2 0 9 2 2
18 0 7 0 9 13 1 9 7 9 7 1 0 7 0 9 10 9 2
18 1 0 7 3 0 9 15 9 9 13 7 3 15 13 10 0 9 2
27 1 3 0 11 2 15 1 10 9 13 9 14 9 2 15 13 9 0 9 2 15 15 1 9 13 11 2
20 3 2 16 15 9 9 13 1 0 0 9 2 13 7 1 0 9 0 9 2
37 10 0 9 1 9 9 13 9 2 16 9 2 7 9 9 7 9 1 10 9 2 13 7 10 9 13 14 3 2 2 16 4 15 3 13 2 2
19 15 13 1 10 9 2 0 15 1 9 9 7 9 2 9 7 15 9 2
14 1 9 7 1 9 3 13 0 9 0 9 2 2 2
16 1 9 13 13 14 0 0 9 9 2 7 7 9 10 9 2
42 11 11 13 10 9 1 9 14 1 0 9 2 7 13 1 9 1 0 9 3 10 9 2 10 0 9 1 9 11 3 13 9 7 0 9 2 15 9 9 3 13 2
9 9 1 12 0 9 13 9 9 2
19 11 11 15 13 1 3 0 2 3 0 0 9 1 0 9 9 7 9 2
21 11 11 13 0 2 9 0 9 2 7 1 10 9 3 13 1 9 7 0 9 2
23 1 9 9 0 9 7 0 9 13 0 9 9 2 16 1 10 0 9 15 13 3 0 2
27 0 9 1 0 9 13 0 2 7 0 9 9 2 1 15 13 9 1 0 9 7 1 9 9 7 9 2
7 0 2 0 9 13 9 11
20 9 0 2 11 2 0 9 0 0 9 2 13 0 9 1 9 0 9 11 2
23 1 0 9 9 9 11 11 15 13 11 11 2 0 0 7 0 9 3 1 9 0 9 2
28 9 13 0 0 9 11 11 2 1 0 9 9 0 11 0 1 11 2 3 1 9 7 9 11 2 11 11 2
20 13 1 15 10 9 7 0 9 1 0 9 2 15 1 9 0 0 9 13 2
54 0 9 13 11 11 0 2 2 11 2 2 11 11 2 11 2 7 11 11 2 11 2 2 1 0 9 15 13 11 11 2 9 2 2 11 11 2 9 1 11 2 7 11 11 1 9 1 11 11 2 9 11 2 2
21 9 11 12 2 13 11 11 2 9 11 11 11 2 0 0 2 11 11 11 0 2
52 1 9 13 0 7 0 9 9 9 11 2 1 11 11 2 15 3 13 1 0 9 1 9 0 11 11 2 1 15 13 3 11 11 2 1 0 9 1 11 11 2 7 11 11 2 1 0 9 1 11 2 2
19 1 9 13 1 0 2 11 7 9 9 2 9 2 9 7 0 9 9 2
19 9 7 9 13 1 9 11 11 2 15 9 0 9 9 1 9 3 13 2
24 9 9 13 0 9 7 13 1 15 0 2 0 9 7 10 9 1 9 1 0 9 1 9 2
26 3 13 0 9 1 11 1 9 0 9 9 2 0 2 0 9 7 9 2 7 0 9 1 0 9 2
27 9 2 3 16 0 9 2 13 13 1 0 9 7 9 2 7 13 7 0 9 1 9 0 9 7 9 2
32 0 2 11 13 9 11 1 9 11 11 7 1 9 10 0 9 11 11 2 15 0 9 1 0 9 13 3 3 1 0 9 2
17 12 1 10 0 9 13 9 12 3 0 9 2 15 7 11 13 2
16 9 11 11 7 13 9 3 3 2 7 15 14 1 9 9 2
13 10 9 15 7 1 9 0 2 11 9 4 13 2
14 11 11 13 9 0 2 11 3 1 0 9 9 11 11
5 15 2 3 2 3
21 9 9 9 0 9 11 11 13 3 7 3 2 12 2 1 9 0 9 1 11 2
21 0 9 1 11 13 3 2 12 2 9 0 9 11 11 9 9 1 9 11 11 2
22 0 9 1 11 13 1 3 9 9 9 11 11 1 9 12 0 9 1 9 11 11 2
11 9 0 9 1 9 13 1 9 11 11 11
22 0 9 11 11 11 13 12 2 9 1 0 9 1 11 0 9 0 0 9 1 9 2
33 0 9 13 9 2 0 7 0 9 7 9 2 15 15 13 3 1 0 11 2 1 0 2 11 7 1 9 0 2 11 7 11 2
22 1 0 9 15 3 1 9 13 11 2 11 2 11 2 11 2 11 2 11 7 11 2
20 1 0 9 15 1 11 13 3 0 9 2 0 0 9 7 0 9 1 11 2
27 3 13 7 0 9 2 0 9 0 9 2 0 0 9 2 0 0 9 7 9 0 11 7 9 1 11 2
18 1 9 9 13 0 9 11 2 9 1 11 7 9 0 9 1 11 2
31 1 9 9 15 4 13 0 0 0 9 0 11 1 11 2 9 0 2 2 9 0 9 7 9 0 9 0 9 0 9 2
17 0 9 13 0 0 9 2 9 0 9 2 0 9 7 0 9 2
4 0 0 0 9
29 9 9 11 11 2 12 2 12 2 2 9 0 0 0 9 2 4 13 0 9 1 0 0 9 2 0 0 9 2
22 1 10 9 15 3 0 0 9 3 1 9 0 9 1 0 11 13 0 9 0 9 2
31 0 0 9 1 10 9 2 3 9 12 1 11 13 10 9 2 0 2 15 13 7 1 9 10 9 11 2 9 7 9 2
17 15 3 13 1 11 1 11 11 7 3 3 13 16 9 0 9 2
29 1 10 0 9 13 9 0 0 9 2 13 4 9 9 2 1 15 15 13 1 15 13 9 3 1 9 0 9 2
13 9 15 1 0 0 9 3 13 9 1 0 9 2
17 10 3 0 0 9 15 13 2 16 13 10 9 1 9 0 9 2
30 0 9 3 1 9 0 2 3 0 2 9 2 0 0 9 7 0 9 1 0 0 9 13 7 0 9 3 3 0 2
38 15 13 11 11 2 15 1 0 7 0 9 11 11 13 3 3 0 0 9 2 12 2 2 0 9 2 1 0 0 9 7 1 0 9 3 0 9 2
19 3 0 9 15 13 0 9 9 2 12 1 9 0 9 2 9 11 11 2
17 15 13 3 0 9 9 7 9 0 9 16 9 7 9 10 9 2
35 9 0 0 9 13 0 0 9 9 2 12 2 3 0 0 9 2 15 0 9 13 0 9 2 7 3 3 0 9 1 9 1 0 9 2
21 0 9 13 3 10 9 7 13 15 9 3 3 7 1 0 2 16 3 0 9 2
1 3
17 0 0 9 9 0 9 11 11 2 12 2 12 2 4 3 13 2
19 0 9 11 2 9 15 3 13 1 0 9 2 15 13 10 9 0 9 2
24 9 13 0 0 9 2 10 9 9 1 0 9 7 12 1 0 9 10 0 9 9 1 15 2
5 11 2 11 15 13
20 0 9 11 11 2 12 7 12 2 15 13 1 11 1 10 0 9 0 11 2
23 0 9 0 9 0 9 15 4 3 13 1 0 0 0 9 7 3 1 9 1 0 11 2
12 1 9 9 11 11 13 1 0 9 0 9 2
5 9 0 9 1 11
15 9 9 1 11 3 13 9 0 9 0 9 1 0 9 2
16 9 13 9 0 9 1 12 12 9 0 1 9 12 7 12 2
16 0 9 9 13 0 0 1 15 7 13 14 12 12 0 9 2
28 9 9 13 9 1 9 9 0 0 9 2 3 11 2 11 2 11 2 11 2 11 2 11 7 11 2 11 2
17 13 7 7 1 9 0 9 2 3 11 2 11 7 11 2 11 2
20 0 9 9 13 9 0 9 2 1 0 1 9 11 2 11 7 11 2 11 2
22 9 9 12 2 7 12 2 9 2 3 2 11 2 11 7 11 2 11 2 9 13 2
3 16 13 9
1 9
2 9 2
28 9 0 9 11 11 1 9 15 13 3 13 0 9 7 3 3 13 0 9 9 2 1 15 3 13 3 13 2
35 9 10 9 15 10 9 13 1 9 13 0 0 9 2 13 1 9 11 11 0 9 7 1 9 11 11 0 9 2 12 1 9 12 2 2
11 0 9 7 1 0 9 9 0 9 13 2
31 11 15 3 13 1 10 0 9 2 13 0 9 11 7 13 1 11 2 7 13 3 0 0 9 0 9 2 0 0 9 2
49 9 2 15 3 13 2 15 13 3 1 9 0 9 1 9 0 0 9 7 9 9 2 13 7 0 0 9 2 9 9 9 7 9 13 9 3 3 0 9 2 1 15 13 9 0 13 0 9 2
21 9 15 3 13 1 9 1 9 7 3 3 9 9 13 9 2 3 13 11 11 2
6 3 11 13 0 9 2
6 3 11 13 11 2 2
51 0 9 0 9 4 7 3 1 10 9 13 3 0 7 0 2 9 13 2 16 9 13 3 0 11 2 7 7 3 2 1 0 9 10 9 2 0 9 2 1 0 9 3 0 9 10 9 7 0 9 2
14 1 10 9 4 3 3 13 9 1 0 9 0 9 2
47 15 1 9 0 9 13 15 0 16 13 9 0 7 0 11 2 1 9 2 2 13 0 0 9 1 9 11 2 9 13 1 9 3 11 2 7 1 0 9 13 2 0 9 2 1 11 2
25 11 10 9 3 13 1 0 9 1 9 0 7 0 11 7 2 3 3 2 1 15 13 0 9 2
23 3 7 3 13 12 1 0 9 9 2 3 10 9 2 3 10 9 2 15 13 3 13 2
65 7 3 3 10 9 0 9 2 3 1 9 9 11 2 15 9 13 3 1 9 12 13 12 9 9 1 9 2 7 9 2 15 4 1 10 9 9 13 14 1 0 9 2 13 1 0 9 9 0 9 7 0 9 1 0 0 9 2 3 16 15 13 0 9 2
14 9 3 0 9 15 1 10 9 13 1 9 0 9 2
18 0 9 9 2 9 1 0 9 0 9 0 9 2 7 3 13 13 2
30 11 15 13 1 15 2 15 3 1 9 13 1 9 9 7 3 0 9 0 9 9 2 7 15 14 1 3 0 9 2
38 0 13 7 10 9 1 15 2 10 9 0 9 7 0 9 4 3 13 0 9 0 9 2 15 4 13 16 3 0 7 0 15 13 1 9 2 2 2
27 13 0 15 13 0 9 3 2 1 0 9 9 0 11 2 7 13 15 1 15 2 15 1 15 9 13 2
15 11 11 11 11 2 15 13 3 7 15 13 0 0 9 2
16 13 10 9 2 11 12 2 16 12 2 9 9 9 7 9 2
7 13 11 11 7 11 11 2
4 9 16 0 9
15 9 11 2 0 9 11 11 2 1 0 9 11 7 0 11
5 0 9 1 0 9
7 0 9 13 9 0 0 9
20 2 11 4 3 9 13 1 9 9 2 3 15 3 13 3 1 0 9 2 2
26 10 9 13 9 11 11 0 9 11 1 9 2 15 3 2 1 12 2 9 2 13 1 0 0 9 2
31 9 9 15 7 13 3 11 2 7 1 0 9 7 0 9 2 13 15 3 13 1 9 1 9 15 12 0 9 7 9 2
22 15 7 13 13 0 9 9 2 1 0 9 0 9 1 2 0 2 2 3 0 9 2
29 9 9 2 1 0 9 1 0 9 0 9 2 13 11 15 2 16 13 3 0 9 2 16 4 13 16 0 15 2
18 9 0 9 3 13 0 9 0 0 9 2 12 11 2 12 0 9 2
13 1 10 9 13 0 9 2 7 7 0 9 9 2
12 1 12 9 13 0 3 13 2 13 2 13 2
34 1 0 9 15 7 0 9 13 10 9 1 9 9 1 0 9 11 1 9 1 9 9 2 7 15 7 1 0 0 9 0 0 9 2
20 1 11 7 11 13 1 0 9 9 2 15 4 15 13 13 9 3 14 9 2
13 1 9 15 3 1 11 13 9 0 9 0 9 2
30 1 15 0 7 0 9 13 11 15 9 3 2 9 0 9 11 13 3 14 1 15 10 9 2 15 13 1 0 9 2
26 0 9 15 13 3 11 11 2 0 9 0 0 9 2 7 3 3 11 11 2 15 13 0 0 9 2
23 9 0 9 3 13 2 16 0 9 13 9 0 9 0 9 7 13 4 1 15 13 0 2
14 9 2 9 1 11 2 3 13 0 7 3 0 9 2
6 3 13 9 1 9 2
59 1 10 9 13 9 0 9 7 0 9 9 2 10 9 2 9 14 13 9 9 7 13 0 9 2 7 2 9 9 4 3 1 15 0 9 2 15 1 15 13 1 9 0 9 2 13 2 7 2 0 0 13 1 11 2 13 9 9 2
14 13 9 2 15 15 13 1 9 1 0 9 9 9 2
22 1 10 9 10 9 1 10 9 13 0 0 9 2 15 3 13 0 9 7 13 9 2
7 1 9 13 9 7 9 2
22 9 13 4 13 1 0 9 10 0 9 2 13 2 1 10 9 1 0 9 0 9 2
13 15 13 10 0 0 9 7 15 1 10 9 13 2
12 15 7 3 15 3 13 7 15 1 15 13 2
1 13
16 9 1 2 9 2 0 9 1 10 9 0 9 15 13 0 2
33 1 9 11 1 11 3 9 7 13 2 7 0 3 13 3 9 2 2 15 9 9 0 9 11 13 1 9 9 1 0 0 9 2
16 13 2 16 1 10 9 13 3 0 9 7 3 13 1 0 2
27 16 9 9 13 9 1 9 10 0 9 1 10 9 2 4 13 10 9 1 9 1 9 9 1 10 9 2
22 13 2 16 15 15 13 1 0 9 1 10 9 2 2 2 2 7 3 12 9 9 2
17 1 11 3 13 9 9 9 2 15 15 1 15 9 0 9 13 2
22 0 9 3 7 13 13 7 12 9 7 0 9 0 9 10 9 1 9 3 3 13 2
8 2 1 11 10 9 13 13 2
20 15 3 13 3 0 9 7 15 16 4 15 13 1 11 2 15 4 13 9 2
28 13 4 2 16 15 13 9 2 15 1 9 9 13 13 3 1 11 2 2 2 2 13 9 9 7 9 9 2
20 9 1 2 9 2 0 11 13 1 0 11 2 3 1 15 13 3 0 9 2
8 3 4 13 1 9 0 9 2
9 1 9 0 13 3 0 7 0 2
41 13 0 9 1 0 9 2 2 1 15 2 16 13 9 0 9 2 13 3 0 2 13 15 1 15 0 9 2 7 3 15 13 1 9 9 2 2 13 0 9 2
28 16 15 9 0 9 13 2 10 9 1 15 13 2 0 9 13 7 0 9 15 13 7 1 9 1 9 13 2
25 15 15 13 1 11 2 0 13 1 9 1 0 11 7 13 15 1 9 2 15 3 4 3 13 2
13 0 9 16 1 11 13 7 9 1 11 9 11 2
18 12 3 15 14 9 2 15 13 4 13 1 9 2 13 9 7 9 2
19 0 9 2 3 4 9 9 9 13 2 13 0 9 9 7 9 1 11 2
23 3 9 1 0 9 15 13 1 9 2 9 2 9 7 9 9 2 15 15 1 9 13 2
10 1 9 10 1 15 13 1 0 9 2
14 13 15 7 0 2 16 9 15 13 2 13 7 13 2
5 15 15 3 13 2
6 0 9 4 3 13 2
16 11 13 0 9 2 3 4 3 1 10 9 13 3 1 11 2
10 13 4 3 3 0 9 2 9 11 2
32 0 9 1 9 12 7 12 9 4 1 15 13 1 9 0 9 2 9 1 9 2 1 9 1 0 0 9 1 11 1 11 2
11 1 9 11 13 1 10 9 7 0 9 2
13 13 15 9 1 9 2 1 15 13 13 0 9 2
24 13 15 7 13 1 0 0 9 10 9 0 9 1 0 9 2 3 1 11 2 11 2 11 2
13 0 9 10 9 13 9 9 1 9 1 0 9 2
10 9 1 0 9 15 1 10 9 13 2
16 7 15 15 13 1 9 1 9 2 7 7 15 13 9 9 2
15 9 13 9 7 9 2 3 13 9 2 1 15 13 13 2
6 9 13 3 10 9 2
13 9 9 9 1 11 7 1 0 9 4 3 13 2
20 3 9 11 13 9 0 9 1 10 9 14 1 0 9 16 2 1 9 2 2
23 13 15 2 16 13 0 9 13 2 7 0 9 4 1 9 1 15 14 1 9 3 13 2
2 0 9
28 15 2 15 1 9 0 9 1 0 9 13 2 13 9 9 9 2 9 2 0 2 2 15 15 13 0 9 2
13 10 9 9 2 11 7 15 9 1 0 9 13 2
23 1 15 15 0 9 13 1 15 3 16 3 0 11 7 1 15 15 9 3 7 3 13 2
36 3 9 9 11 11 11 13 1 9 9 3 2 0 9 9 9 11 2 0 9 2 2 15 15 13 1 9 11 1 9 1 9 9 9 9 2
15 9 9 7 13 2 16 13 0 10 0 9 1 10 9 2
14 0 0 9 13 15 2 16 0 9 3 13 16 9 2
15 0 12 9 7 13 13 1 9 1 9 7 3 15 13 2
3 9 1 11
15 15 13 3 9 9 0 0 9 9 1 9 1 0 9 2
22 13 15 3 9 2 16 13 9 10 9 2 16 0 9 1 0 2 0 9 13 0 2
16 0 9 2 0 9 9 1 9 7 0 9 3 13 3 9 2
28 13 7 9 0 9 3 3 0 2 16 4 15 1 15 13 13 16 1 0 9 7 0 9 13 9 7 9 2
30 1 15 15 1 10 9 7 0 9 13 3 9 9 2 15 3 13 9 1 10 9 7 1 15 2 15 13 9 9 2
18 13 3 9 0 9 7 0 9 2 16 13 1 0 1 11 0 9 2
29 13 2 16 1 3 0 9 2 15 13 0 9 4 3 3 13 0 9 1 10 11 1 0 9 16 1 0 9 2
33 9 11 11 11 2 2 16 13 2 13 15 2 16 4 15 13 3 2 16 4 15 13 9 9 1 9 7 16 0 9 13 9 2
19 14 13 3 13 2 16 15 11 3 13 0 1 9 1 11 2 2 2 2
2 0 9
14 11 11 2 2 9 9 13 3 1 0 7 0 9 2
18 1 9 15 16 13 2 13 15 2 15 13 1 10 0 9 0 9 2
12 9 2 9 2 9 2 9 2 9 7 0 2
9 10 9 13 2 7 13 15 13 2
6 15 13 0 9 2 2
25 10 9 13 11 11 2 9 1 0 9 9 2 15 13 9 1 11 1 0 0 9 11 2 11 2
15 9 13 1 0 9 16 0 0 9 9 2 9 2 9 2
51 1 9 12 4 1 0 9 9 11 13 2 1 9 0 9 1 0 9 1 11 2 13 1 0 11 2 3 16 7 1 0 9 2 1 11 2 11 2 11 2 11 2 2 0 9 1 0 9 7 9 2
15 9 3 13 1 10 9 13 7 3 15 13 3 1 11 2
8 3 4 9 13 3 1 15 2
35 2 9 11 13 1 15 0 9 2 13 1 15 1 9 9 9 0 9 2 2 13 15 11 11 2 9 0 1 9 0 9 1 0 9 2
16 2 13 15 1 9 2 15 15 14 0 9 13 1 0 9 2
9 7 7 15 13 1 15 0 9 2
19 13 15 9 2 9 2 10 9 13 1 9 2 9 9 2 9 1 9 2
7 1 10 9 15 13 9 2
20 13 9 9 2 10 2 9 2 2 3 2 9 2 2 2 13 11 2 11 2
20 1 0 9 9 15 13 9 2 16 0 9 1 10 0 9 13 13 10 9 2
12 1 9 13 9 2 9 9 2 9 2 9 2
6 9 13 1 0 9 2
10 13 3 13 9 2 9 7 0 9 2
5 13 15 10 9 2
10 3 15 9 15 13 7 15 15 13 2
6 13 15 3 3 0 2
12 0 9 15 3 3 13 1 0 2 9 2 2
13 0 9 1 9 13 3 0 9 16 1 0 11 2
16 3 0 9 11 1 15 13 1 0 12 9 9 9 0 9 2
12 9 1 0 9 2 9 7 9 1 0 9 2
11 12 9 12 10 9 13 10 9 1 9 2
10 9 4 13 1 9 2 0 2 0 2
12 0 3 13 9 1 9 9 9 9 1 11 2
32 9 11 11 3 1 0 9 13 2 16 9 13 9 1 9 2 2 7 9 1 11 13 2 7 4 13 10 9 1 9 2 2
13 9 0 0 9 11 11 13 12 1 9 0 9 2
19 0 9 1 0 9 13 2 16 0 7 0 9 15 9 1 11 3 13 2
4 13 1 15 2
24 9 2 15 15 1 10 9 13 2 13 14 1 0 9 7 1 9 2 15 15 13 1 9 2
12 2 14 2 15 4 10 9 1 10 9 13 2
11 15 15 13 3 3 2 16 15 3 13 2
15 3 4 1 9 1 9 13 0 9 16 9 0 9 2 2
10 10 9 0 9 13 1 11 3 0 2
10 9 11 11 13 1 9 0 0 9 2
25 16 13 11 2 3 1 15 15 13 2 0 9 1 9 2 9 1 9 9 2 9 1 9 2 2
7 11 11 3 15 3 13 2
6 13 15 3 1 11 2
16 13 15 1 0 9 9 7 1 9 2 16 9 15 13 13 2
2 3 2
10 2 16 13 11 2 2 13 11 11 2
6 15 0 13 1 11 2
13 0 9 9 11 1 9 13 9 1 0 9 3 2
5 13 4 15 3 9
24 13 2 16 13 15 1 15 2 9 1 0 9 2 3 0 2 13 15 1 9 1 0 9 2
14 7 3 13 15 13 1 9 10 9 2 15 3 13 2
50 13 1 9 1 15 2 16 9 2 3 9 9 2 3 2 3 15 13 3 2 4 1 0 9 13 10 2 9 9 2 2 9 9 0 1 15 9 7 3 0 9 2 16 3 13 0 2 7 0 2
44 13 2 14 1 0 9 1 9 16 1 9 3 3 0 7 3 3 0 2 0 9 2 13 15 3 13 15 2 15 15 13 1 0 9 2 15 4 13 14 3 0 9 9 2
29 13 15 10 2 3 0 9 13 3 16 9 2 7 1 9 7 1 9 9 3 2 13 10 9 9 3 16 0 2
63 15 3 13 0 9 1 9 0 9 9 2 11 2 11 2 11 2 1 10 0 0 2 1 15 9 0 9 9 2 11 11 2 1 0 0 0 2 0 7 1 9 1 9 0 9 7 11 11 1 3 0 2 14 0 2 3 1 0 9 0 0 9 2
12 3 13 1 9 10 9 3 1 0 9 0 2
30 1 10 9 15 13 9 2 13 1 9 9 2 7 3 7 1 9 9 10 3 0 9 2 3 0 1 9 0 9 2
24 13 10 9 0 0 7 0 9 1 9 10 0 9 1 9 1 15 2 16 3 13 0 9 2
37 13 2 14 15 3 2 3 10 9 1 9 2 7 14 3 2 13 9 2 7 3 3 10 2 9 2 0 9 2 15 10 9 13 9 15 0 2
44 16 3 13 1 15 2 16 9 7 9 13 0 9 9 7 16 10 9 10 9 13 2 13 3 3 0 13 1 15 9 2 16 9 10 3 0 9 4 14 3 13 10 9 2
9 15 3 13 3 9 9 10 9 2
17 13 15 15 0 2 16 4 0 9 13 15 3 0 16 15 0 2
14 13 15 15 3 2 16 0 9 13 9 1 9 0 2
22 16 4 2 9 9 2 7 1 15 0 7 0 9 9 0 13 13 2 3 4 13 2
24 13 2 14 3 1 15 2 16 13 10 9 9 2 3 13 10 10 9 3 13 10 0 9 2
51 3 4 15 13 13 13 0 9 10 1 0 9 3 3 2 7 3 6 3 2 2 0 9 2 3 13 10 9 2 13 2 3 4 13 2 7 3 3 13 2 7 13 15 13 2 15 13 14 10 9 2
20 1 0 0 9 4 15 13 3 9 2 3 10 0 9 2 0 15 1 9 2
3 9 0 9
23 1 9 10 0 9 13 3 9 2 16 4 15 3 13 1 3 0 9 0 9 0 9 2
19 10 0 9 0 9 7 13 0 9 2 16 0 9 7 9 13 3 3 2
22 16 3 0 9 13 13 9 11 11 2 10 9 9 2 2 11 12 2 12 2 12 2
15 0 9 9 1 9 13 2 13 1 9 2 0 7 0 2
27 13 15 2 3 4 3 1 0 9 13 2 1 12 0 9 2 7 13 3 3 1 9 13 9 3 0 2
28 9 15 1 9 13 1 9 2 15 1 15 12 13 9 9 2 0 9 7 9 1 9 1 0 9 0 9 2
30 9 15 13 1 3 0 9 9 14 3 2 13 2 14 0 9 0 0 9 2 7 3 15 0 9 1 9 0 9 2
23 15 3 13 10 9 1 2 0 9 9 7 9 2 7 3 9 2 7 3 3 3 13 2
8 3 13 0 0 9 0 9 2
12 13 3 3 0 2 16 1 9 9 13 9 2
27 11 7 13 2 16 4 15 10 10 9 13 2 7 16 13 1 15 13 7 1 0 9 1 9 1 11 2
46 11 0 9 3 13 2 16 9 0 9 0 2 9 0 9 2 2 3 13 9 1 9 7 1 0 9 2 15 4 15 1 10 0 9 3 3 13 9 0 9 1 15 7 1 15 2
12 3 13 2 15 13 1 9 1 9 0 11 2
23 10 0 9 13 14 3 0 9 9 0 9 2 15 13 11 2 11 7 10 0 9 11 2
39 13 15 2 16 3 0 13 0 9 9 0 9 2 3 15 1 9 13 0 9 7 0 9 11 11 1 3 0 9 7 0 0 9 0 9 2 11 11 2
19 1 9 11 13 15 9 3 0 7 1 0 9 0 2 16 3 3 0 2
36 16 4 15 10 9 13 0 9 7 10 9 3 2 16 13 3 2 0 9 13 3 9 0 0 9 2 2 10 9 4 3 13 1 9 3 2
43 13 4 7 13 2 16 11 13 7 0 9 2 7 0 0 9 2 7 3 3 0 9 9 0 9 2 15 13 1 0 9 0 9 7 1 15 15 3 1 0 9 13 2
13 1 9 9 2 9 7 9 11 7 13 0 9 2
29 13 3 0 9 0 9 2 3 15 3 2 3 1 0 0 9 2 13 10 9 2 3 16 0 0 9 0 9 2
31 1 15 13 11 3 1 10 9 9 1 0 9 2 15 10 0 9 9 3 13 2 9 1 9 9 0 9 1 9 9 2
13 3 13 0 0 9 0 9 7 1 15 0 9 2
16 0 9 0 9 13 16 10 0 9 2 3 0 9 7 9 2
20 11 7 13 7 3 0 2 7 3 0 9 2 14 9 0 9 2 9 11 2
22 0 9 13 2 13 2 1 0 0 9 9 11 2 16 14 15 13 7 3 3 13 2
7 13 15 3 1 3 3 2
34 3 1 0 9 2 15 13 0 0 9 2 1 0 9 7 9 1 15 2 15 0 9 7 9 13 7 13 15 0 2 16 0 9 2
10 0 0 9 0 9 3 3 4 13 2
14 7 16 2 3 1 0 0 9 2 1 9 2 2 2
4 3 13 1 0
7 7 11 13 9 0 0 9
20 9 2 1 10 0 9 13 9 0 0 9 2 13 0 9 1 0 0 9 2
20 3 7 13 0 9 1 15 10 10 0 9 2 3 15 3 13 1 0 9 2
33 16 13 11 11 3 10 9 2 15 1 0 9 0 9 1 10 10 9 13 2 13 15 3 1 10 9 13 7 1 10 0 9 2
11 3 1 10 3 0 9 1 11 7 11 2
6 11 9 11 13 0 2
45 13 15 10 0 9 7 10 9 2 15 3 13 11 3 2 2 9 13 1 11 0 9 2 16 11 15 13 13 10 9 1 9 0 9 1 0 9 2 1 0 7 0 9 2 2
31 13 11 16 9 0 0 9 2 13 10 11 2 15 13 1 0 9 9 7 4 13 2 13 1 9 7 13 1 0 9 2
32 13 1 9 2 16 1 0 0 9 9 12 13 0 11 12 9 9 2 13 0 9 2 15 0 0 9 13 1 9 1 11 2
30 13 2 15 1 10 9 13 7 3 0 7 15 3 13 10 9 1 9 10 11 2 15 13 7 0 9 1 0 9 2
35 1 9 12 0 9 13 1 11 16 1 9 0 9 1 9 2 7 13 1 15 0 9 2 9 2 16 0 9 4 13 3 2 15 13 2
14 9 2 15 0 9 13 9 2 1 0 9 3 13 2
42 9 1 9 0 9 3 13 13 1 10 9 1 9 7 1 3 2 3 0 2 9 10 9 15 13 3 3 10 9 11 2 15 15 13 0 9 13 2 13 7 13 2
17 13 15 7 2 16 4 15 3 3 13 1 11 9 0 0 9 2
19 9 15 13 2 16 1 0 9 13 13 7 3 2 16 15 13 11 11 2
61 3 16 0 9 11 11 1 9 12 2 2 1 9 1 15 2 1 9 1 15 7 1 9 1 9 2 16 15 9 13 9 13 2 15 13 1 15 2 1 15 4 15 13 13 2 13 0 9 1 9 7 13 1 9 9 7 10 9 7 9 2
21 13 15 1 15 2 16 4 4 13 0 7 0 9 1 15 7 1 15 9 2 2
21 15 0 9 13 13 1 9 1 15 2 3 13 9 2 15 15 13 1 12 9 2
30 3 1 15 13 1 12 9 9 0 0 9 9 9 0 9 2 1 0 9 9 0 1 9 13 9 7 0 11 3 2
48 3 15 7 3 13 1 9 0 9 1 11 2 16 1 9 1 9 11 7 1 9 1 0 9 11 2 11 2 3 13 1 0 9 11 7 1 9 1 9 0 9 11 7 1 11 0 11 2
38 0 1 15 2 15 11 13 11 2 4 13 0 13 7 1 11 2 1 0 9 1 11 11 2 15 4 1 0 9 13 10 9 7 1 9 0 9 2
31 7 11 13 9 0 9 2 13 1 9 12 11 1 11 1 9 1 0 9 7 13 1 9 12 9 3 0 9 1 11 2
24 7 1 11 13 9 0 2 0 9 2 2 11 2 0 9 1 9 9 9 1 0 0 9 2
23 3 2 16 4 4 7 11 13 3 2 16 4 13 9 2 15 1 11 13 0 0 9 2
27 7 15 13 14 9 0 9 10 2 15 15 3 13 2 3 2 16 15 9 0 9 9 1 0 9 13 2
39 3 9 1 0 9 13 0 9 3 9 2 3 13 0 3 7 3 13 1 9 2 0 15 0 9 1 0 9 0 9 2 3 0 13 13 7 3 13 2
44 16 11 13 2 13 15 13 9 9 7 13 1 0 2 15 13 14 0 2 13 13 15 0 9 2 2 13 1 12 1 0 9 2 1 15 15 1 0 0 9 3 15 13 2
37 1 15 15 13 7 9 0 2 3 2 9 13 9 9 1 10 9 2 13 0 9 9 0 9 9 1 0 2 0 9 7 13 9 1 9 9 2
40 7 3 10 9 15 13 2 16 4 1 12 9 13 7 11 3 16 14 16 9 0 9 7 9 9 2 15 4 3 1 11 14 1 9 0 9 13 0 9 2
20 11 15 13 13 10 0 9 1 0 9 7 7 15 1 15 14 1 9 13 2
21 3 1 9 10 0 0 9 15 13 1 9 2 15 1 15 13 0 9 1 9 2
57 9 1 2 0 9 2 7 9 13 10 0 9 13 3 1 0 9 9 2 7 3 1 0 9 15 9 13 3 13 2 3 0 13 0 2 0 9 2 1 15 15 3 13 9 7 9 1 0 2 0 9 0 2 0 0 9 2
20 0 9 7 9 10 11 15 13 9 1 15 9 7 9 0 15 0 0 9 2
14 13 4 7 0 2 16 4 15 15 13 3 3 13 2
41 11 4 13 2 13 7 9 9 3 13 0 9 11 13 2 13 15 13 16 0 9 9 1 0 9 0 9 7 13 0 9 2 3 15 1 0 9 13 11 11 2
35 16 13 11 16 2 9 0 9 1 9 1 11 2 2 3 15 13 11 2 2 3 4 15 13 13 7 1 9 7 9 0 7 0 9 2
5 0 0 2 0 9
23 0 2 0 9 13 10 9 0 9 2 13 15 3 13 2 9 7 9 15 1 9 13 2
13 10 9 9 15 7 1 9 0 9 13 13 0 2
28 0 9 2 12 2 12 2 2 13 2 16 0 9 1 2 9 2 0 9 2 0 9 2 13 3 0 9 2
21 14 10 9 1 15 3 13 7 13 1 0 0 9 1 9 3 7 1 15 15 2
11 1 9 15 9 13 13 7 1 0 9 2
29 0 2 0 9 13 9 12 0 2 7 0 9 2 15 13 0 9 9 7 13 1 15 14 3 1 12 9 9 2
15 9 13 1 9 2 7 1 9 7 0 9 1 12 9 2
35 7 16 1 9 12 4 1 11 7 0 11 13 0 9 2 16 1 11 2 2 13 14 9 13 15 2 16 0 9 13 3 1 0 9 2
24 13 3 3 0 2 7 0 2 2 0 2 9 1 9 1 0 9 13 1 15 9 0 9 2
11 3 1 9 9 13 13 9 1 10 9 2
18 11 13 1 0 0 9 10 9 2 13 10 0 7 2 0 2 9 2
40 3 0 9 1 12 2 9 15 7 3 13 1 9 7 1 9 1 2 15 0 2 1 9 2 15 7 15 13 7 13 13 7 1 0 2 7 1 0 9 2
19 9 12 13 13 1 9 12 2 12 7 12 2 3 3 13 11 2 11 2
47 9 9 13 15 1 0 9 11 2 11 7 11 2 1 0 0 9 2 13 15 14 0 9 2 3 1 9 0 9 2 7 13 15 0 9 11 7 11 2 2 3 13 0 15 2 2 2
27 0 11 13 13 2 16 0 9 13 9 0 9 2 15 11 13 7 15 3 13 3 15 0 1 0 9 2
5 15 15 3 13 2
16 16 15 3 3 13 0 9 2 3 13 1 0 2 0 9 2
15 3 11 13 2 16 1 9 9 11 13 9 1 0 9 2
13 0 11 3 13 2 16 13 1 11 10 0 9 2
15 1 10 9 13 10 9 9 2 13 1 9 1 0 9 2
6 15 3 13 13 15 2
42 12 16 9 10 9 0 9 1 11 3 7 3 13 2 7 1 15 3 9 2 0 2 2 0 2 0 2 0 2 9 13 9 1 9 2 15 13 13 0 9 11 2
19 1 10 9 13 0 13 0 9 2 9 2 1 9 12 16 9 0 9 2
15 9 9 13 9 9 2 15 3 13 9 1 0 0 9 2
13 10 9 14 13 2 16 0 9 7 9 9 13 2
17 11 7 11 13 3 1 0 9 2 13 10 0 2 0 2 9 2
35 13 1 15 13 9 10 9 1 0 0 9 2 1 15 13 3 2 9 2 9 2 7 7 0 9 2 0 9 2 0 9 2 0 11 2
8 10 9 4 13 13 9 9 2
26 13 4 15 3 16 3 15 0 2 0 9 2 7 16 9 9 0 9 2 7 16 0 9 7 9 2
56 13 15 13 12 0 2 9 2 2 12 5 12 2 2 1 0 9 9 9 2 1 0 2 2 0 9 7 0 9 2 7 14 16 0 0 2 0 9 2 1 2 9 2 2 2 1 9 0 0 2 0 7 0 9 0 2
15 9 9 2 0 9 2 9 1 0 9 1 9 0 9 2
7 9 13 9 10 9 1 11
2 0 9
1 9
19 9 1 9 1 11 13 3 0 9 9 11 2 0 9 1 9 0 9 2
23 11 2 15 1 12 9 13 12 0 9 2 13 1 9 13 0 9 7 13 15 0 9 2
28 9 0 9 2 13 9 11 1 9 0 9 2 2 13 10 9 1 9 1 11 0 9 11 1 11 11 11 2
26 13 2 16 4 13 1 9 0 9 1 9 0 9 2 15 13 13 15 9 9 2 0 9 1 9 2
25 11 3 15 13 9 9 11 2 0 11 2 16 4 15 13 1 9 2 15 13 1 9 0 11 2
8 11 9 13 13 0 0 9 2
11 2 1 10 9 4 13 0 9 1 11 2
11 3 15 15 13 2 2 13 3 9 11 2
9 2 13 1 0 7 0 9 11 2
17 4 13 1 0 2 15 1 15 13 2 2 13 12 1 9 11 2
7 0 9 11 13 3 0 2
22 13 13 1 11 2 13 15 13 1 9 7 13 9 1 0 0 9 2 7 13 13 2
10 0 12 9 15 3 13 1 9 9 2
13 9 13 9 7 10 9 2 1 9 7 1 9 2
28 11 3 3 13 12 9 2 9 2 16 13 9 11 2 15 1 0 9 1 9 12 3 13 1 0 9 9 2
23 1 9 0 9 13 0 9 11 11 1 0 9 10 0 9 9 9 1 11 1 0 11 2
27 13 1 9 2 0 9 2 1 15 2 3 4 1 0 9 13 9 2 9 2 9 7 0 9 0 9 2
13 1 10 9 15 3 13 14 11 2 11 7 11 2
13 11 13 3 1 9 1 11 1 10 0 9 13 2
16 15 2 15 13 11 1 9 1 11 2 7 13 1 10 9 2
9 13 1 15 9 0 9 15 11 2
9 7 15 13 7 1 0 9 11 2
10 9 1 9 11 13 7 10 0 9 2
14 2 1 9 9 13 9 2 16 10 9 13 16 9 2
16 13 15 7 13 1 9 3 2 2 13 15 12 1 9 11 2
34 1 2 0 9 2 2 15 11 3 13 1 11 2 13 7 9 9 7 9 2 9 9 1 9 7 9 9 9 1 9 1 9 9 2
18 3 15 3 10 0 9 13 2 16 3 13 0 9 7 3 15 13 2
11 9 9 11 1 11 3 13 13 1 9 2
11 13 14 9 0 9 2 0 0 9 2 2
6 1 0 13 10 9 2
6 9 1 9 3 13 2
23 16 1 15 13 7 9 11 2 4 13 11 3 14 12 0 9 2 9 2 9 7 9 2
4 15 13 11 2
3 1 0 9
75 1 9 2 3 0 11 3 3 13 0 9 9 1 9 2 0 0 9 2 2 11 2 12 2 2 7 16 15 13 3 15 10 9 2 13 12 9 10 9 2 15 13 7 11 7 11 2 3 3 2 13 15 2 9 2 1 3 0 9 2 15 4 3 13 13 9 9 2 13 9 0 9 0 11 2
13 9 0 0 9 7 9 13 1 9 3 3 9 2
27 3 12 11 2 9 7 0 0 9 2 15 11 1 9 12 13 1 2 9 2 2 13 0 9 10 9 2
29 11 15 3 2 3 13 0 9 16 0 9 2 2 13 11 11 1 0 0 0 9 7 0 2 0 9 15 13 2
18 1 11 15 9 1 11 13 14 2 0 2 9 2 9 2 3 9 2
12 15 13 3 13 9 9 7 9 1 0 11 2
30 13 13 2 16 1 3 0 2 0 9 2 0 9 2 3 1 0 0 9 2 15 3 10 0 9 13 1 9 9 2
11 2 11 1 10 9 3 13 0 9 2 2
23 15 0 9 1 11 3 13 9 2 16 4 0 9 4 13 2 7 13 2 13 0 11 2
40 3 13 0 13 2 16 9 2 15 11 9 12 2 9 13 1 9 1 0 0 9 2 1 15 11 13 2 13 9 1 10 2 16 4 3 13 9 0 9 2
13 16 4 12 9 13 9 2 13 11 1 0 9 2
18 3 15 13 2 3 0 9 15 13 1 9 2 7 3 1 0 9 2
16 13 0 13 0 9 2 15 15 13 13 14 1 0 0 9 2
20 15 15 4 13 13 9 2 0 9 2 2 11 11 2 7 3 7 0 9 2
30 3 3 15 11 11 13 1 11 13 16 2 0 11 2 2 9 0 0 9 1 9 12 2 12 2 9 9 11 2 2
16 11 4 13 0 0 9 2 15 10 9 3 13 7 3 13 2
8 11 13 1 11 2 11 1 11
30 3 2 1 9 11 2 13 0 2 16 9 11 13 3 3 0 1 11 7 1 15 1 0 9 7 9 11 1 11 2
21 15 13 9 0 9 1 12 9 0 0 9 7 15 13 9 0 7 0 0 9 2
10 13 15 3 1 9 11 9 11 11 2
8 3 15 13 0 13 2 13 2
24 15 13 9 1 0 11 2 9 9 11 7 0 0 9 2 13 11 2 7 10 9 13 9 2
18 1 0 2 0 9 4 13 3 0 9 9 9 11 11 1 0 9 2
25 9 0 9 2 9 0 9 1 9 2 0 9 2 4 13 9 1 9 11 1 0 7 0 9 2
18 11 11 1 11 3 3 13 2 16 9 1 11 13 11 13 3 11 2
18 0 0 7 0 9 1 11 2 9 2 9 11 7 9 9 13 0 2
20 3 10 9 13 13 0 9 0 9 2 15 4 1 15 13 13 0 0 9 2
25 14 3 0 9 2 1 0 9 2 13 0 9 9 1 3 0 9 0 1 9 9 2 13 9 2
12 11 15 0 9 2 1 0 9 2 13 13 2
23 13 2 16 0 9 15 1 15 13 1 9 2 7 15 13 13 10 0 9 2 13 9 2
1 3
37 11 7 11 15 1 0 9 0 9 9 11 11 1 11 13 1 9 1 9 0 9 2 11 2 7 11 15 13 13 3 1 9 1 9 11 11 2
23 9 0 9 13 2 16 1 10 9 0 15 11 2 4 13 1 9 2 1 0 14 2 2
10 13 2 16 1 0 9 15 4 13 2
31 0 9 11 11 3 13 11 11 9 9 2 11 11 9 1 9 2 15 4 13 1 9 2 7 11 11 9 0 0 9 2
9 9 1 10 9 13 9 11 11 2
47 9 0 9 2 11 2 11 11 13 3 9 7 9 0 0 0 9 2 11 2 2 16 4 15 13 1 0 9 2 1 15 13 1 9 1 11 1 9 12 1 9 1 9 1 11 11 2
27 1 9 0 9 2 15 4 13 0 9 1 11 2 0 11 2 2 13 3 1 11 1 12 9 0 9 2
22 9 9 13 2 16 4 15 1 0 9 1 11 13 3 1 0 9 2 15 13 9 2
39 0 9 1 11 11 11 13 1 0 9 10 0 9 9 9 2 1 15 7 0 9 2 16 4 15 13 2 16 13 1 9 13 9 9 1 9 9 11 2
15 9 1 9 11 1 11 15 13 1 0 0 9 9 9 2
7 13 15 3 3 0 9 2
20 13 2 16 1 0 9 2 15 1 9 13 9 7 9 2 4 13 12 9 2
15 1 15 13 12 0 9 0 1 9 1 2 0 2 9 2
8 12 15 13 9 1 0 9 2
30 9 0 0 9 0 0 9 7 9 0 9 15 3 3 13 1 9 0 9 2 1 10 9 13 13 9 11 11 11 2
19 11 1 9 13 2 16 0 13 3 0 9 9 2 13 7 13 0 9 2
15 9 11 13 3 1 9 0 0 9 13 9 11 2 11 2
4 0 9 1 11
4 11 2 11 2
26 9 1 9 0 9 1 12 9 0 9 7 10 0 9 1 0 11 13 3 3 3 0 9 0 9 2
7 13 1 15 0 0 9 2
31 1 10 9 15 9 0 9 13 1 0 9 0 9 7 0 9 2 11 2 1 0 9 3 1 11 1 0 9 9 13 2
28 9 0 9 4 13 7 1 0 9 11 14 2 11 0 15 3 1 0 9 1 0 2 0 9 0 0 9 2
15 0 9 13 9 0 11 16 9 1 9 1 0 0 9 2
32 11 13 1 11 1 0 9 0 9 2 1 15 1 0 9 3 13 2 16 10 9 13 1 9 0 9 7 10 9 1 11 2
10 1 9 3 1 9 13 9 12 9 2
16 10 9 3 3 13 0 9 11 11 1 9 10 9 10 9 2
16 11 13 2 16 0 9 1 12 9 13 4 13 1 12 9 2
16 3 1 12 9 13 3 1 0 11 2 3 13 9 9 11 2
18 1 11 15 13 0 9 13 13 1 2 9 9 2 2 16 13 11 2
13 9 1 11 7 11 13 3 0 9 1 0 9 2
29 11 13 1 15 2 16 4 15 11 3 13 1 0 11 2 16 0 9 13 2 16 4 0 9 13 1 0 9 2
17 0 9 13 13 11 2 16 4 15 13 1 9 9 1 0 11 2
15 11 3 13 0 9 1 9 1 0 11 1 0 9 11 2
27 1 0 9 13 12 11 1 9 9 1 11 2 1 2 11 9 0 1 9 1 0 9 0 0 9 11 2
10 11 11 3 1 11 13 10 0 9 2
6 11 11 13 1 0 9
2 11 2
29 10 9 1 0 9 2 0 15 9 9 1 0 9 11 1 0 9 1 9 12 2 3 13 0 9 11 11 11 2
11 3 3 13 2 16 1 9 13 15 0 2
26 0 0 9 9 1 0 9 11 11 14 1 9 13 2 16 1 0 9 10 9 3 1 9 11 13 2
43 1 0 9 0 11 0 7 1 9 13 2 16 3 9 15 7 3 0 9 0 0 9 11 11 7 9 9 11 11 13 2 16 9 11 4 13 13 0 9 2 9 2 2
10 15 12 10 9 3 13 2 13 11 2
5 11 7 11 13 9
4 11 2 11 2
24 1 9 9 1 0 0 9 2 15 4 13 1 12 9 2 15 3 3 13 9 11 7 11 2
14 0 9 3 1 0 9 13 2 16 11 13 0 9 2
17 1 0 9 9 11 11 13 0 9 0 11 2 3 0 9 2 2
8 10 0 9 7 13 1 9 2
21 0 9 11 2 11 13 2 16 4 9 13 10 9 2 7 13 1 0 9 11 2
5 9 0 9 1 11
2 11 2
24 0 0 9 1 9 11 13 13 13 0 9 11 1 9 7 13 14 14 13 10 9 0 9 2
29 13 15 9 9 9 11 11 2 15 13 9 12 0 9 2 12 9 7 12 9 7 9 2 1 15 9 13 11 2
20 13 2 16 1 9 1 0 9 0 9 13 9 13 1 2 9 7 9 2 2
15 11 7 13 2 16 1 10 9 4 0 9 13 0 9 2
5 9 1 9 1 11
2 11 2
22 12 9 7 12 0 15 1 0 9 13 0 9 0 9 1 9 1 0 0 9 11 2
23 1 9 13 9 0 0 9 2 3 9 2 0 1 11 1 9 0 9 9 9 0 9 2
20 9 0 0 9 1 11 9 11 2 11 13 2 16 9 4 13 0 0 9 2
16 2 9 13 13 3 1 9 2 7 1 11 2 2 13 11 2
12 1 15 13 1 9 0 1 9 9 9 9 2
6 0 9 13 9 1 9
21 0 0 0 9 1 11 13 4 13 3 2 16 0 9 13 12 1 15 0 9 2
15 1 9 1 0 0 9 11 15 3 1 11 13 9 11 2
37 2 1 10 9 4 1 0 13 2 13 7 13 12 9 2 12 0 9 2 12 9 0 7 12 9 2 2 13 15 9 9 2 12 0 11 11 2
9 0 9 13 9 7 0 0 9 2
5 0 9 1 0 9
2 11 2
16 0 9 1 0 9 1 9 11 7 11 13 1 9 1 9 2
22 0 0 9 13 2 16 15 9 13 3 1 9 0 11 2 3 13 0 9 11 11 2
18 1 9 15 9 1 0 9 3 13 1 9 0 11 13 9 0 9 2
18 1 10 9 13 3 1 9 0 0 9 1 0 9 0 0 9 11 2
25 1 9 0 9 2 15 13 1 9 9 2 15 3 13 9 0 2 3 0 2 9 7 0 11 2
28 1 9 9 11 13 12 9 1 9 1 0 9 7 1 9 0 9 1 9 9 0 9 1 9 9 1 9 2
10 0 9 2 0 9 7 2 10 9 2
9 13 1 9 13 15 3 0 9 2
36 13 4 15 3 2 13 1 15 2 15 13 10 0 9 2 2 13 1 9 9 9 11 11 2 0 0 9 1 0 9 9 1 10 9 2 2
30 0 9 0 9 1 0 9 4 3 14 13 13 1 15 2 16 9 4 2 13 9 0 9 10 9 7 10 9 2 2
11 13 1 9 11 11 2 13 4 15 13 2
19 1 9 13 7 0 13 2 16 3 3 4 15 13 13 2 0 2 9 2
34 12 9 15 3 13 2 16 9 13 10 0 9 2 1 15 15 0 9 1 10 9 13 9 9 2 16 4 15 15 13 1 0 9 2
24 15 1 15 13 2 9 3 3 13 2 9 13 3 1 15 2 16 13 15 3 0 16 9 2
12 13 15 3 0 9 0 9 2 9 7 9 2
21 13 3 3 16 0 9 0 9 2 16 13 3 0 9 13 1 12 3 0 9 2
24 0 11 13 13 16 9 2 15 2 13 13 15 7 0 2 1 9 1 9 2 7 9 9 2
19 13 9 2 1 0 9 2 10 9 1 10 3 0 0 9 13 3 0 2
39 3 16 13 2 16 9 2 9 9 2 7 9 3 3 13 9 2 7 3 3 2 16 7 2 9 0 2 9 13 10 9 0 2 7 16 2 3 2 2
23 13 2 14 3 13 10 9 2 13 15 1 15 0 13 1 9 2 15 13 1 0 9 2
21 16 15 13 0 9 2 13 15 9 0 7 0 2 3 7 13 2 3 0 2 2
16 13 15 9 1 9 9 2 13 15 3 9 0 9 10 9 2
22 13 2 14 15 3 2 13 2 1 0 9 0 0 9 2 13 9 3 0 9 9 2
32 13 1 15 13 15 0 1 9 7 13 15 1 9 11 11 1 9 0 9 2 13 15 1 10 2 0 9 0 9 2 2 2
20 1 15 3 13 2 13 3 9 9 1 10 0 0 9 1 9 11 7 11 2
38 13 1 9 2 14 7 1 0 2 10 9 0 9 9 2 2 9 0 1 15 2 15 1 15 13 2 2 7 1 9 0 2 0 2 9 0 9 2
37 1 0 2 2 0 2 9 15 13 2 15 15 15 13 7 3 1 15 13 9 0 9 2 1 0 9 13 7 10 0 9 3 13 10 0 9 2
22 1 15 0 13 0 9 0 9 2 1 15 0 13 1 15 2 1 10 9 0 9 2
27 1 0 9 13 1 9 1 9 7 13 9 0 15 0 2 1 0 3 7 3 13 2 13 7 3 13 2
14 0 13 3 10 9 2 13 15 15 2 15 13 9 2
32 11 11 13 2 11 1 12 2 9 2 1 9 0 9 2 16 10 9 3 13 9 2 15 11 13 0 2 9 1 0 9 2
37 9 1 0 9 4 7 13 13 9 9 3 0 2 10 9 2 3 0 9 0 9 2 4 3 13 13 1 15 2 15 13 7 3 15 13 13 2
4 9 2 9 2
13 9 0 9 13 9 0 2 3 14 3 0 9 2
11 13 15 1 9 10 0 0 9 1 11 2
28 13 2 16 15 15 9 9 13 2 16 15 10 9 3 13 1 0 9 2 1 15 13 0 9 9 10 9 2
16 9 2 15 9 0 11 15 13 1 0 0 9 13 1 9 2
47 16 1 0 0 9 13 1 0 9 10 9 1 9 12 11 11 2 13 1 15 3 9 11 11 11 1 15 2 16 0 9 13 3 0 7 13 3 0 13 7 0 2 3 2 0 9 2
24 10 9 7 13 7 10 9 13 2 16 0 9 2 3 0 9 2 15 1 9 9 14 13 2
14 11 10 9 1 0 9 13 9 10 0 9 1 9 2
26 0 9 15 7 3 13 2 7 7 3 11 13 1 9 11 7 10 9 0 9 13 1 0 0 9 2
14 0 9 13 9 9 0 9 13 0 9 3 0 9 2
13 1 9 15 13 9 2 15 3 0 9 3 13 2
12 7 7 13 10 0 2 9 2 9 0 9 2
8 15 0 13 14 12 1 0 2
27 0 9 13 1 0 9 10 9 11 1 0 0 9 9 0 9 0 9 9 12 1 9 11 1 0 9 2
37 1 0 9 4 13 0 13 2 16 15 2 15 13 13 13 1 9 0 9 0 9 2 1 9 1 10 9 13 7 13 15 13 10 9 3 3 2
20 0 0 9 15 7 13 10 9 9 11 13 7 13 9 11 1 9 7 9 2
6 1 9 3 13 9 2
35 0 9 11 1 0 9 0 15 1 9 13 14 9 0 9 1 9 0 9 2 7 3 9 9 2 1 15 4 9 11 1 0 9 13 2
27 1 3 0 0 9 15 1 10 9 13 13 2 7 13 0 9 10 9 1 9 1 9 1 0 0 9 2
9 16 0 3 0 9 4 15 13 2
20 9 7 9 1 11 11 2 1 11 2 15 2 13 7 13 0 9 11 2 2
30 7 16 11 15 3 3 13 13 10 0 9 0 9 7 0 9 2 13 15 9 10 0 9 1 9 7 1 10 9 2
22 3 15 3 13 0 2 7 9 2 9 9 7 9 1 0 0 9 3 13 0 9 2
38 1 15 15 7 9 0 9 2 7 15 14 1 9 0 9 2 13 9 2 16 10 0 9 15 1 11 15 13 3 1 9 2 1 15 15 3 13 2
70 1 9 1 2 0 0 9 2 2 1 15 13 3 3 9 14 1 9 11 2 7 3 7 1 15 2 16 4 15 13 1 9 2 2 13 0 9 2 9 9 0 1 9 9 7 9 1 0 7 0 9 2 1 9 9 1 0 9 2 7 2 9 0 3 1 0 9 9 2 2
7 9 13 15 7 3 0 2
16 9 3 13 14 9 1 9 9 0 2 0 2 0 3 9 2
15 9 13 0 9 9 2 15 13 13 13 9 0 7 0 2
4 3 7 0 2
27 0 9 15 13 10 0 9 1 9 7 9 9 2 7 3 10 9 2 15 0 9 13 1 0 9 3 2
16 13 13 9 9 2 0 9 1 9 2 7 9 13 0 9 2
36 15 7 13 2 16 9 1 9 9 13 1 0 9 9 2 16 0 9 9 13 1 9 0 9 2 16 0 9 13 1 9 0 7 0 9 2
27 10 9 13 13 3 1 9 2 16 9 15 13 2 16 13 13 9 7 16 10 0 9 15 13 4 13 2
15 0 9 2 3 0 9 9 2 13 9 10 0 9 9 2
10 15 4 3 13 4 3 13 0 9 2
26 9 10 9 4 13 14 9 1 9 2 7 9 1 0 9 4 13 3 10 9 2 15 13 11 0 2
7 9 15 1 15 3 13 2
6 9 14 2 7 15 3
1 9
27 1 0 9 4 15 13 15 9 9 1 9 9 13 0 12 9 9 12 9 3 3 13 1 9 7 9 2
9 13 0 13 2 13 7 3 13 2
15 0 9 13 3 14 9 9 2 15 9 1 9 3 13 2
8 15 15 13 1 12 9 9 2
8 1 9 13 9 3 12 9 2
18 9 9 15 7 1 9 1 9 13 3 1 0 9 0 9 1 9 2
20 0 9 7 3 13 2 16 0 9 15 13 13 2 16 13 10 9 3 0 2
17 9 7 3 3 13 0 1 15 2 16 4 15 15 9 3 13 2
30 9 9 3 13 2 16 13 13 0 9 9 2 1 0 9 13 15 1 15 7 0 2 16 13 13 3 0 9 9 2
26 12 12 9 2 15 15 9 13 2 4 13 13 3 12 9 2 9 15 3 13 13 1 3 0 9 2
8 9 15 3 13 3 1 9 2
21 10 9 13 1 9 2 16 9 4 13 9 9 1 9 12 0 9 3 3 13 2
9 13 1 15 7 3 0 0 9 2
21 1 15 4 9 13 1 9 15 3 9 1 9 2 15 3 4 1 15 9 13 2
16 9 13 2 16 1 0 9 13 9 9 3 0 2 3 3 2
22 13 7 13 2 16 1 10 0 9 1 0 0 9 13 9 0 9 7 3 0 9 2
9 9 9 13 3 13 9 13 0 2
7 9 4 7 13 13 15 2
10 13 13 9 1 9 7 13 9 9 2
27 13 0 13 9 2 16 4 13 0 7 3 14 0 9 1 9 2 15 4 15 13 13 1 2 0 2 2
27 15 4 10 9 13 3 0 1 9 0 9 7 13 4 15 13 15 2 15 3 3 13 1 0 0 9 2
7 3 3 15 3 3 13 2
1 9
1 9
12 11 11 13 11 11 9 2 7 15 13 3 2
23 9 2 15 1 0 9 13 10 0 9 2 13 0 2 16 0 9 0 9 10 9 13 2
24 11 11 15 3 13 9 1 0 9 2 3 15 13 0 9 7 0 9 1 15 1 15 13 2
29 0 9 9 7 0 9 2 15 1 9 13 10 9 1 9 2 1 15 13 2 13 0 2 12 9 13 9 9 2
9 10 9 7 13 0 2 13 0 2
22 0 9 3 13 2 16 7 1 9 2 15 13 13 9 9 7 9 2 13 0 9 2
9 0 9 7 13 0 7 0 9 2
35 11 11 1 9 0 9 13 2 16 7 9 2 7 0 9 13 10 9 9 1 9 15 0 2 7 7 15 1 9 1 0 9 13 13 2
5 15 13 3 9 2
33 1 0 9 9 13 1 9 0 3 0 9 2 3 2 0 9 9 2 15 15 13 2 13 13 0 0 9 7 13 15 0 9 2
14 1 0 0 9 13 4 9 1 9 9 9 7 13 2
8 3 13 13 3 9 0 9 2
14 1 0 9 9 13 3 2 9 0 9 7 0 9 2
33 15 2 15 9 13 13 9 1 9 7 0 9 2 4 15 13 1 0 9 11 11 13 1 15 2 16 13 12 9 0 7 3 2
31 1 0 9 3 7 1 15 2 13 2 14 0 13 15 1 0 9 1 9 9 9 7 1 9 10 0 9 13 10 9 2
17 1 10 0 9 3 13 9 2 10 9 13 1 10 9 3 0 2
3 3 0 9
1 9
30 11 11 13 10 9 1 0 0 9 1 0 9 2 16 9 13 1 9 12 2 9 1 0 12 1 14 12 9 3 2
11 13 4 0 2 16 4 15 3 3 13 2
31 13 7 9 9 2 16 4 15 9 1 0 9 1 10 2 15 7 3 13 2 13 7 13 2 13 3 3 0 0 9 2
6 0 9 9 13 0 2
30 13 1 15 0 9 9 2 0 9 10 9 7 9 0 9 13 3 0 9 9 9 2 3 2 9 0 9 0 9 2
30 3 7 3 13 2 16 9 9 2 9 2 9 2 0 9 2 9 7 9 0 9 1 0 9 1 9 9 3 13 2
13 0 9 1 9 0 9 7 13 1 0 9 9 2
20 10 9 13 1 0 0 9 0 9 2 15 3 13 0 13 1 9 7 12 2
36 3 13 3 0 3 13 3 0 9 0 15 1 0 0 9 2 13 9 2 7 13 3 9 9 1 9 2 15 4 15 13 13 1 9 9 2
20 1 0 9 0 9 13 12 3 0 2 1 0 9 13 7 9 2 7 9 2
14 15 3 13 2 7 3 1 9 2 15 4 13 13 2
31 9 0 1 9 13 3 7 0 9 9 1 0 9 7 0 9 1 9 13 3 3 0 2 16 9 9 9 7 3 13 2
15 1 0 9 2 15 3 13 3 2 3 3 13 3 13 2
56 0 9 9 1 0 9 9 7 9 13 1 0 0 9 7 0 9 9 2 15 15 13 9 2 15 1 15 13 0 9 0 3 7 3 3 10 0 9 1 10 0 9 2 7 16 1 0 0 2 7 3 7 0 2 9 2
44 13 15 3 2 16 16 4 3 13 11 11 11 1 0 9 1 9 1 9 1 9 10 2 9 2 15 13 9 2 2 13 4 1 9 2 16 4 13 9 0 9 16 9 2
18 13 3 2 16 1 15 12 12 9 4 1 10 9 3 15 13 13 2
15 9 1 0 9 9 15 7 1 10 9 13 13 3 0 2
26 3 0 9 0 9 2 15 13 3 3 1 11 2 13 9 0 9 2 7 3 0 9 7 0 9 2
7 7 15 3 13 10 9 2
6 13 15 1 0 0 9
2 0 9
2 11 2
11 1 9 1 11 11 3 13 9 11 11 2
29 13 2 16 0 1 9 12 13 10 0 0 9 2 15 3 1 9 13 3 0 3 2 16 15 1 15 13 13 2
25 2 13 2 16 9 13 11 2 11 2 2 13 7 13 2 16 9 1 10 9 13 7 10 9 2
19 1 0 0 9 4 1 9 0 9 13 12 9 9 2 15 0 13 9 2
20 9 13 2 16 11 2 11 13 0 9 9 1 10 9 2 16 13 1 9 2
19 3 2 16 9 13 0 2 13 10 9 9 9 2 15 13 1 9 11 2
27 11 3 13 0 13 2 16 13 3 1 10 9 2 7 16 15 9 2 15 9 13 2 4 1 9 13 2
10 0 15 15 13 9 7 9 0 9 2
37 1 10 9 13 0 2 16 1 9 9 13 1 9 2 7 15 16 9 1 9 13 1 9 11 2 3 13 1 11 9 7 13 15 14 12 9 2
16 11 4 13 1 9 0 9 7 0 9 1 0 9 0 9 2
22 1 0 15 1 9 13 13 1 9 9 1 11 1 11 9 1 9 3 12 9 9 2
18 3 4 13 1 0 9 9 14 1 12 9 7 1 9 9 0 9 2
7 0 9 1 9 12 13 0
6 11 11 1 9 1 11
30 9 0 9 2 9 7 9 2 0 9 1 9 7 9 9 9 1 9 2 15 13 0 9 0 9 1 9 11 11 2
34 1 9 1 0 9 4 10 9 13 2 16 0 0 9 13 3 1 12 7 12 9 2 7 16 9 1 9 9 4 13 13 12 9 2
7 13 15 9 14 3 0 2
9 0 9 1 10 9 15 3 13 2
7 9 9 12 13 0 9 2
22 16 13 0 9 2 15 13 0 13 2 3 13 9 2 3 4 15 10 9 13 9 2
21 12 7 0 9 1 9 9 2 1 9 10 9 1 0 9 2 13 1 3 0 2
13 15 13 2 16 10 9 4 13 2 3 3 2 2
14 13 15 3 3 0 9 9 16 12 7 12 9 3 2
8 13 1 0 9 7 0 9 2
11 0 9 9 13 3 0 9 1 0 9 2
24 1 10 0 9 1 10 9 13 15 2 15 13 1 9 1 9 1 15 2 3 1 12 9 2
13 13 4 1 9 10 0 9 1 12 7 12 9 2
15 13 15 13 2 16 4 15 13 1 12 9 10 9 13 2
13 1 0 9 13 3 1 9 0 9 1 9 9 2
24 13 15 3 2 16 13 10 9 1 0 2 7 15 13 2 16 9 13 0 7 13 10 9 2
12 3 13 2 16 4 13 3 1 0 9 9 2
34 13 9 2 16 15 1 0 9 13 13 1 9 2 3 13 13 9 2 7 15 15 13 1 0 9 15 2 0 9 2 9 2 9 2
10 13 2 16 13 15 0 7 3 0 2
22 13 9 2 15 10 9 13 0 9 2 13 1 15 9 2 7 3 13 0 9 3 2
11 9 15 1 9 9 3 13 3 16 9 2
19 1 0 9 11 7 9 1 10 9 13 2 7 3 1 15 7 10 9 2
5 15 15 15 13 2
7 0 9 13 3 0 9 2
20 9 15 3 13 1 9 0 9 2 0 1 0 9 2 3 3 1 9 9 2
16 15 13 9 2 3 9 9 13 7 10 9 13 1 0 9 2
12 9 1 9 0 9 10 9 9 9 11 13 2
12 13 7 9 2 16 4 10 9 13 1 0 2
4 9 13 0 9
3 1 0 9
2 11 2
21 16 1 0 9 9 1 0 9 13 11 2 11 0 0 9 2 13 13 15 13 2
24 3 3 7 13 1 9 2 16 1 9 13 9 12 9 0 9 16 9 1 9 9 1 9 2
9 13 1 15 3 9 9 11 11 2
26 9 13 1 12 9 7 3 4 13 9 9 1 9 9 1 9 1 9 12 9 1 12 9 0 9 2
20 1 11 9 13 13 1 9 13 15 0 9 7 13 15 13 9 1 9 9 2
7 13 13 7 11 7 11 2
3 9 0 9
25 13 15 9 12 2 9 9 1 9 13 11 7 3 4 13 13 11 2 1 9 9 2 7 0 2
8 11 11 2 11 2 2 9 2
27 13 4 15 2 16 4 1 9 13 3 10 11 2 3 16 4 10 9 1 9 13 1 9 9 0 9 2
24 13 4 3 0 9 1 15 2 16 4 15 13 9 11 1 10 9 13 16 9 7 0 9 2
7 1 9 11 15 13 13 2
27 13 15 13 15 2 16 15 13 1 3 0 2 7 3 0 9 2 7 3 1 11 7 15 7 1 11 2
7 10 9 13 1 11 0 2
9 1 9 9 4 13 9 0 9 2
40 11 11 2 11 2 11 2 2 9 2 13 15 2 16 4 9 11 13 0 1 9 2 16 4 15 13 0 9 1 0 2 0 9 2 7 2 3 9 9 2
9 12 2 9 13 1 15 0 9 2
10 9 11 1 9 13 3 3 0 9 2
25 13 0 2 16 7 0 0 9 13 10 9 0 2 7 16 0 13 15 3 3 2 16 13 0 2
13 13 4 15 7 3 2 16 11 13 1 9 9 2
8 11 11 2 11 2 2 9 2
20 16 13 9 1 0 0 9 2 3 13 0 2 13 2 14 3 7 9 11 2
14 7 16 15 10 9 0 9 13 2 3 1 15 13 2
6 1 9 11 4 13 2
11 13 0 2 16 4 13 13 1 15 0 2
8 11 11 2 11 2 2 9 2
11 9 13 0 9 7 11 3 10 9 13 2
11 7 15 13 2 16 4 11 13 13 13 2
9 3 3 2 16 13 9 2 2 2
8 11 11 2 11 2 2 9 2
13 13 15 1 11 2 7 13 15 3 1 10 9 2
10 13 9 2 16 4 1 15 15 13 2
8 1 11 4 1 0 3 13 2
9 15 4 3 13 3 9 1 9 2
8 11 11 2 11 2 2 9 2
7 11 4 15 3 13 13 2
20 13 0 9 13 3 7 1 1 15 2 16 9 10 9 15 13 3 1 9 2
18 13 2 16 9 4 13 1 9 9 12 9 7 1 10 9 13 9 2
9 1 10 9 13 9 9 11 0 2
10 9 0 2 0 2 11 2 13 1 9
2 11 2
45 9 0 2 0 2 11 2 2 15 13 0 9 7 13 1 9 9 0 9 2 13 1 12 2 9 12 9 9 0 1 9 0 9 1 0 9 0 7 1 9 2 0 0 9 2
14 9 0 9 9 1 15 3 13 9 9 9 11 11 2
13 9 4 13 4 13 1 0 9 1 12 2 9 2
21 1 12 2 9 13 0 2 0 2 11 2 1 11 13 0 12 9 0 9 9 2
10 14 3 13 0 9 1 9 1 9 2
24 9 13 2 16 9 13 10 9 2 16 1 15 0 2 0 2 11 2 13 1 9 0 9 2
32 16 3 13 1 3 0 9 2 0 3 0 9 2 13 0 2 0 2 11 2 16 9 1 9 0 9 0 16 12 12 9 2
14 0 9 3 3 13 3 13 10 9 1 12 0 9 2
53 2 13 1 9 2 3 0 13 0 9 13 2 16 0 13 2 2 13 11 1 9 1 9 16 9 0 9 9 2 11 2 2 15 9 7 0 9 13 2 7 0 2 0 2 11 2 2 9 2 9 2 0 2
28 9 14 1 9 13 1 9 12 9 3 2 7 3 12 12 13 0 13 1 9 9 2 16 15 9 3 13 2
22 9 9 11 11 2 11 2 13 9 1 0 9 1 1 10 0 9 1 0 9 9 2
25 9 9 11 11 13 2 16 10 0 0 9 11 11 2 15 13 1 9 9 2 13 1 0 9 2
11 2 13 15 2 13 15 9 2 2 13 2
26 16 4 1 15 13 0 9 7 0 2 0 2 11 2 1 9 13 2 13 4 4 13 0 0 9 2
10 9 14 3 3 13 0 7 0 9 2
25 11 3 3 13 2 16 9 0 9 1 9 0 9 2 1 12 2 9 2 15 13 12 9 9 2
15 9 12 4 13 1 9 9 2 0 9 1 9 0 9 2
14 9 13 13 9 12 0 2 9 2 1 9 0 9 2
14 2 15 15 1 15 13 2 2 13 9 1 9 11 2
9 9 13 1 9 1 0 9 3 0
2 11 2
26 3 1 9 9 11 2 11 7 11 1 9 0 9 13 13 9 2 16 4 13 9 0 9 0 9 2
24 2 0 2 9 9 13 12 9 11 2 9 0 9 11 11 7 9 3 2 0 9 11 11 2
38 16 1 9 9 15 13 12 9 11 2 11 11 2 11 11 2 11 11 2 15 11 2 11 2 7 11 11 2 11 2 15 3 1 12 9 9 13 2
16 11 11 2 11 2 15 13 2 12 1 12 9 9 13 0 2
32 11 2 11 2 11 2 1 9 13 2 16 10 0 9 1 9 0 2 0 0 9 1 0 9 1 12 12 9 9 13 13 2
20 13 1 0 3 13 1 9 2 15 9 13 3 1 12 9 1 0 0 9 2
32 9 9 11 11 2 11 2 13 9 10 0 9 2 16 1 9 13 13 10 9 1 15 2 2 14 15 15 9 9 13 2 2
25 9 7 9 11 11 7 13 9 0 9 1 0 2 0 9 2 0 3 3 16 12 12 9 9 2
9 9 9 1 0 9 11 13 0 9
2 11 2
32 0 9 1 9 3 12 9 9 2 15 13 0 1 9 0 9 11 2 13 3 3 0 9 2 15 7 13 1 10 9 13 2
18 0 9 15 13 0 9 12 2 9 3 2 0 9 9 9 11 11 2
20 9 0 9 13 9 9 1 0 9 9 2 15 0 9 11 13 1 0 9 2
23 9 4 13 9 13 1 0 9 10 9 7 0 9 4 13 13 13 1 12 2 9 12 2
22 0 9 3 13 1 10 9 1 0 9 13 14 12 9 9 2 12 9 3 9 13 2
12 1 11 2 11 13 0 9 9 0 0 9 2
15 1 3 0 9 15 13 1 9 0 9 9 2 9 3 2
16 14 9 0 0 9 1 0 9 13 14 1 12 7 12 9 2
13 9 9 10 0 9 3 3 3 13 9 0 9 2
14 9 9 11 13 16 0 2 13 3 13 9 0 9 2
7 0 9 11 15 13 9 9
2 11 2
16 0 9 3 0 9 1 0 9 13 9 0 0 9 11 11 2
25 16 3 13 1 10 0 9 1 9 0 7 0 9 9 2 13 1 9 0 7 0 9 7 9 2
23 2 0 2 0 7 0 9 9 2 0 1 10 9 2 13 13 9 9 11 2 2 13 2
27 9 9 11 11 1 9 9 13 2 16 9 1 9 7 9 13 7 3 13 1 0 9 13 9 1 9 2
14 3 3 15 14 13 9 1 0 0 9 2 13 11 2
32 3 0 9 2 9 2 2 15 13 13 0 9 1 9 9 0 2 14 1 11 13 9 9 7 9 9 1 12 9 1 9 2
6 9 7 13 9 9 2
15 1 11 13 10 0 9 3 0 2 16 13 10 0 9 2
17 0 9 9 13 0 2 3 15 13 9 1 9 7 9 0 9 2
22 1 0 9 13 1 11 3 12 9 9 1 15 2 16 4 13 9 13 1 0 9 2
10 9 1 11 11 2 9 9 1 0 9
28 0 9 9 13 10 9 0 9 2 15 4 15 13 13 9 1 9 7 9 9 9 1 9 1 9 7 9 2
13 3 13 10 9 0 7 15 4 3 13 1 9 2
5 10 9 13 0 2
19 13 2 14 9 9 13 1 9 3 0 9 2 13 15 13 1 9 0 2
13 0 9 7 13 13 2 13 2 14 13 1 11 2
14 3 3 15 7 13 13 9 0 9 9 1 9 11 2
18 9 1 0 9 10 9 1 9 13 3 0 2 7 10 9 9 13 2
16 1 9 9 3 13 9 0 9 7 9 1 15 9 13 9 2
12 9 4 7 3 13 2 16 9 10 9 13 2
15 9 1 9 9 4 15 3 13 13 2 3 1 9 9 2
24 9 15 13 1 15 2 16 9 0 9 13 9 7 9 9 2 3 9 2 15 13 0 9 2
5 9 11 11 13 13
3 1 0 9
2 11 2
28 2 0 9 15 13 13 2 2 13 3 9 0 0 9 11 11 2 15 15 3 3 1 0 9 13 1 9 2
23 1 9 11 7 9 4 13 3 2 16 15 1 9 9 13 1 9 9 3 1 9 9 2
18 11 13 9 9 1 10 9 13 1 15 2 16 13 15 9 9 9 2
15 1 0 9 1 9 11 15 1 10 0 9 3 15 13 2
1 3
21 2 9 0 9 2 13 3 1 0 9 1 9 9 2 15 9 1 0 9 13 2
17 0 9 4 13 3 12 9 2 9 7 9 0 2 9 9 2 2
34 0 0 7 0 9 1 9 9 2 15 4 13 13 0 9 7 9 0 9 7 9 11 2 3 13 16 9 9 0 9 11 11 11 2
26 9 9 9 1 9 1 12 2 9 9 11 11 1 9 1 9 11 15 3 13 9 1 0 0 9 2
18 9 13 0 9 2 3 2 9 2 0 9 2 9 12 7 3 11 2
6 0 9 11 13 0 9
4 11 2 11 2
24 9 13 0 9 11 2 11 2 13 3 12 9 2 15 13 1 12 5 3 16 1 9 12 2
15 1 9 9 9 1 9 11 13 0 9 1 9 0 9 2
22 0 9 1 10 0 9 13 9 0 0 7 0 9 2 15 11 13 3 1 9 9 2
24 3 13 9 9 9 11 2 11 11 2 13 9 9 9 7 0 9 2 15 13 9 0 9 2
13 15 13 9 9 13 9 9 7 9 1 0 9 2
12 13 14 1 0 9 3 0 1 15 0 9 2
19 9 13 1 10 0 9 2 0 1 9 11 2 11 0 9 2 0 9 2
23 1 0 9 1 0 0 9 2 15 13 9 1 0 9 2 13 3 9 11 12 9 9 2
13 1 15 13 9 3 9 1 9 1 9 1 11 2
5 0 9 1 9 9
2 11 2
34 3 0 0 9 2 15 13 2 1 0 9 9 13 0 0 9 2 2 13 12 2 9 1 9 9 11 9 0 0 9 1 0 9 2
21 1 0 9 2 1 9 0 9 2 14 13 1 9 1 9 11 1 11 0 9 2
19 15 15 9 4 13 1 0 0 9 7 1 0 9 1 9 1 9 3 2
24 0 9 11 13 9 0 9 7 13 15 1 0 0 9 2 1 15 15 10 9 13 9 11 2
24 0 9 13 3 1 9 9 1 0 9 2 3 15 1 0 9 9 13 1 9 1 0 9 2
18 0 9 13 1 9 9 9 9 2 1 15 15 9 13 2 9 2 2
5 0 9 13 9 9
12 0 9 2 15 4 13 12 9 2 4 13 13
2 11 2
16 0 9 9 0 9 4 3 13 1 9 9 9 1 10 9 2
22 13 15 1 9 0 9 1 0 9 7 9 2 15 3 9 13 0 9 9 1 9 2
8 0 9 13 9 0 9 9 2
17 1 0 0 9 15 13 1 12 2 7 9 10 9 13 1 12 2
19 0 9 4 13 10 9 9 13 1 9 1 9 2 3 9 13 1 9 2
13 3 0 9 4 13 13 10 9 1 9 10 9 2
12 1 9 0 9 4 9 13 13 3 12 9 2
12 9 13 2 16 9 4 13 13 1 0 9 2
28 0 0 9 1 0 2 14 12 9 2 2 0 13 3 1 12 9 2 7 3 0 3 12 7 0 0 12 2
16 10 9 4 15 14 13 9 9 1 0 12 1 12 7 12 2
25 13 15 1 15 2 16 15 15 1 9 13 9 13 2 7 7 4 15 7 13 13 3 16 12 2
22 9 9 11 11 2 11 2 13 2 16 9 13 0 2 7 1 0 9 15 14 13 2
10 13 2 16 9 9 13 12 9 3 2
19 9 3 13 2 16 4 9 1 9 9 3 1 9 13 9 12 9 9 2
10 15 4 15 4 13 1 9 9 9 2
9 3 4 15 13 9 0 9 9 2
22 9 0 9 4 1 9 13 4 1 9 0 2 15 4 13 1 9 0 9 2 13 2
39 9 0 9 0 1 9 0 9 4 4 13 1 15 9 1 1 9 9 2 3 16 9 0 9 1 9 2 16 4 3 13 7 10 9 7 10 0 9 2
20 9 15 13 2 16 4 9 13 13 7 13 9 1 9 0 9 0 0 9 2
10 0 9 4 13 0 9 13 9 9 2
7 13 9 13 0 3 3 2
7 0 9 13 1 9 12 9
2 11 2
25 1 9 7 9 0 9 1 9 11 7 9 0 0 9 13 0 9 9 1 9 3 12 9 9 2
16 1 9 9 13 3 0 0 9 2 0 9 7 0 9 9 2
35 9 7 9 0 9 10 0 9 11 11 4 9 13 1 9 0 7 0 9 2 3 0 9 0 11 11 2 0 9 1 11 7 9 11 2
16 0 9 13 11 11 1 9 9 11 2 15 9 13 0 9 2
17 2 13 4 15 13 2 0 9 4 13 0 9 2 2 13 11 2
6 0 9 4 13 0 9
2 11 2
10 0 9 4 13 1 9 13 0 9 2
12 3 15 11 13 9 0 9 9 11 11 11 2
14 9 13 14 12 9 2 1 15 3 12 9 3 0 2
18 1 9 3 13 9 1 9 2 9 2 9 2 9 7 9 1 9 2
16 9 1 3 3 0 1 0 9 13 3 1 11 11 0 9 2
31 1 9 0 9 2 3 9 11 0 11 13 9 11 2 13 11 9 9 1 9 1 12 9 2 3 15 13 9 1 9 2
15 16 4 11 11 13 13 3 0 2 13 1 9 0 9 2
20 1 9 9 9 1 11 12 15 7 13 2 16 1 0 9 1 11 13 9 2
27 1 0 9 13 0 9 7 3 0 3 1 9 9 13 2 16 13 0 9 2 3 0 9 9 0 9 2
21 11 11 1 9 9 13 2 16 1 3 0 13 0 9 9 7 2 9 9 2 2
7 1 9 13 15 1 9 2
8 0 9 9 13 1 12 9 2
12 1 0 9 11 13 1 9 9 1 9 9 2
10 1 0 9 3 0 13 1 9 9 2
4 1 9 13 9
2 11 2
11 9 0 9 1 11 4 13 9 0 9 2
23 1 9 0 9 0 9 11 11 4 1 9 0 9 2 0 9 1 11 2 13 0 9 2
6 13 3 3 9 9 2
18 11 3 13 10 0 9 2 1 15 4 9 13 1 0 16 0 9 2
21 3 0 9 2 16 9 11 13 11 2 4 13 3 3 2 16 13 9 0 9 2
18 0 9 9 1 9 15 13 1 12 2 1 0 9 13 1 0 9 2
4 3 9 10 9
2 11 2
11 0 9 4 13 9 13 3 1 0 9 2
26 13 15 1 15 9 0 0 9 1 9 9 2 9 7 9 2 15 15 3 13 7 0 7 0 9 2
11 3 4 13 9 13 9 3 1 0 9 2
27 3 15 13 1 15 2 16 4 9 1 0 12 9 9 9 1 0 9 13 3 9 1 15 7 1 9 2
16 12 9 9 15 7 13 14 10 9 2 15 13 9 0 9 2
21 15 13 1 15 2 16 9 13 1 9 15 3 9 2 15 3 1 15 9 13 2
17 9 9 15 13 2 16 3 15 0 9 13 13 9 9 1 9 2
11 3 15 13 9 9 2 15 13 3 0 2
5 0 9 4 14 13
2 11 2
19 12 0 7 0 2 0 9 13 0 9 9 1 9 1 9 1 0 9 2
7 13 15 1 0 9 9 2
17 1 9 13 4 13 9 0 9 0 1 9 0 9 15 13 9 2
17 9 9 13 9 1 9 2 16 9 13 0 7 13 0 9 9 2
20 1 0 4 3 13 9 2 15 4 13 1 9 7 13 9 1 9 0 9 2
3 15 13 9
2 11 11
9 9 0 9 1 9 13 3 9 2
14 14 3 9 15 13 11 7 10 0 9 1 0 9 2
29 14 3 9 0 9 13 0 9 15 9 2 15 1 9 0 9 9 1 11 2 11 7 3 13 9 1 0 9 2
10 3 1 9 12 12 9 13 15 15 2
14 14 15 0 9 1 0 9 13 12 7 9 9 9 2
7 13 9 2 15 13 15 2
27 16 1 0 9 1 0 9 1 11 1 9 0 9 13 9 10 3 3 0 9 2 13 15 3 10 9 2
10 10 9 13 3 3 3 1 10 9 2
16 13 7 0 2 9 1 9 12 10 0 9 10 9 15 13 2
14 13 3 9 2 16 3 1 9 11 10 9 3 13 2
11 16 4 13 15 2 15 3 13 13 15 2
3 13 3 2
16 12 1 3 3 12 9 9 9 0 9 3 3 14 13 4 2
20 9 0 9 1 0 9 7 13 3 0 7 10 9 13 7 1 9 9 9 2
16 0 9 2 11 7 11 2 15 3 14 13 2 13 0 13 2
28 1 0 9 7 13 3 3 1 15 2 16 4 9 13 1 9 0 1 9 0 11 7 1 0 9 11 13 2
21 3 13 1 0 11 2 16 3 13 1 9 9 2 16 4 13 10 9 0 9 2
12 13 9 0 9 1 0 9 9 14 7 13 2
16 15 13 2 16 10 9 4 13 9 0 9 1 9 9 13 2
23 1 9 9 1 9 9 1 9 13 13 3 13 2 16 0 9 13 0 9 9 7 9 2
18 7 15 13 10 9 7 15 15 13 2 16 13 9 7 9 15 13 2
19 1 9 9 9 2 9 10 9 13 14 1 9 0 9 3 12 9 9 2
30 13 15 1 10 9 7 3 13 10 0 9 1 15 2 16 3 13 3 14 9 15 2 15 15 1 10 9 9 13 2
4 15 13 9 2
29 15 1 0 9 7 0 9 13 1 15 2 16 4 10 9 13 3 7 15 2 16 9 13 1 0 7 1 9 2
5 7 15 13 0 2
20 15 3 13 1 9 2 16 0 0 9 4 3 13 1 9 7 9 1 9 2
22 16 9 15 1 15 13 7 13 15 9 9 1 10 9 2 13 3 1 10 0 9 2
6 9 15 13 1 3 9
10 1 9 13 9 0 9 14 12 0 9
2 11 2
17 10 9 1 0 9 13 9 1 10 9 2 16 9 10 9 13 2
9 11 15 3 13 9 10 0 9 2
20 0 0 9 2 15 1 9 9 13 7 1 0 9 2 7 9 4 13 13 2
27 16 11 13 9 9 0 9 9 9 11 11 2 13 1 9 0 9 1 9 12 1 10 9 12 0 9 2
17 9 0 9 15 9 9 9 13 2 16 10 9 9 15 13 15 2
20 1 9 1 0 9 13 0 9 9 2 15 3 13 0 9 2 12 0 9 2
19 1 9 12 9 3 13 9 9 1 0 12 9 12 9 0 9 1 9 2
23 0 0 9 13 1 0 9 11 11 14 12 9 2 3 15 10 9 13 3 1 0 9 2
18 16 7 11 13 2 1 10 9 3 13 1 0 0 9 12 0 9 2
32 9 1 9 9 13 1 10 9 13 3 0 9 0 9 2 3 10 9 7 9 1 9 0 9 3 13 1 12 9 1 0 2
20 2 3 15 13 14 1 9 9 9 2 15 15 1 15 13 2 2 13 11 2
17 3 9 9 9 1 3 0 9 11 13 7 9 10 0 0 9 2
18 1 9 9 9 13 0 9 2 15 15 13 1 3 9 2 3 13 2
23 16 11 13 11 2 11 2 13 1 0 0 9 2 16 4 15 13 2 15 10 9 13 2
12 0 4 1 0 9 13 13 9 9 0 9 2
15 3 13 1 0 9 11 2 10 9 13 7 9 0 9 2
3 9 3 13
2 11 2
29 1 3 0 9 1 0 0 9 1 11 7 11 13 3 0 9 9 7 9 9 11 11 0 9 11 1 0 9 2
33 2 16 15 13 9 2 15 13 13 2 3 13 9 1 10 9 2 2 13 11 7 13 2 16 10 9 13 1 0 9 0 9 2
34 1 9 1 10 9 11 2 11 11 13 2 16 1 0 9 4 13 1 9 0 9 9 2 0 9 2 2 15 4 13 12 5 9 2
15 10 9 4 13 1 9 0 9 2 3 1 10 0 9 2
13 1 9 9 11 13 2 16 13 9 3 10 9 2
19 1 0 9 15 4 13 9 2 3 15 15 13 7 15 4 1 15 13 2
5 0 9 13 11 9
12 13 1 9 9 1 9 9 11 2 13 9 11
2 11 2
29 2 9 9 13 1 15 0 2 16 15 1 9 9 13 7 9 11 2 13 3 13 2 7 13 1 0 9 2 2
28 3 2 3 15 13 12 2 9 12 13 1 9 11 11 0 9 9 11 11 2 0 9 9 9 9 11 11 2
12 13 15 1 9 9 2 15 15 11 13 13 2
8 9 13 1 9 7 9 9 2
36 11 2 12 2 4 1 9 9 12 3 13 16 9 1 9 0 9 11 11 11 7 3 1 12 2 9 13 9 9 9 9 1 9 9 11 2
38 9 9 9 11 11 3 11 13 2 16 1 10 9 15 13 15 2 16 13 1 9 9 1 9 9 11 11 2 7 3 13 9 13 9 9 9 11 2
19 1 15 13 1 9 2 15 13 3 0 7 9 9 3 15 13 1 9 2
14 11 13 1 11 3 1 9 1 9 9 9 0 9 2
16 2 9 1 10 9 1 9 3 13 2 2 13 0 9 11 2
23 1 15 11 4 15 13 9 0 0 9 2 1 15 13 7 0 0 9 2 9 11 11 2
23 11 3 13 2 16 11 3 13 1 0 2 0 9 2 10 9 4 13 3 1 0 9 2
23 2 9 1 9 11 1 9 11 11 1 12 9 13 9 2 15 13 0 9 0 9 9 2
17 13 13 2 15 1 10 9 11 11 13 7 13 2 2 13 11 2
6 11 2 9 15 13 0
13 2 11 13 0 9 2 15 13 13 1 0 9 2
19 9 15 13 0 2 13 15 9 0 9 2 13 15 9 1 9 0 11 2
29 9 10 9 7 10 9 0 9 13 3 9 13 3 15 2 15 15 11 13 2 16 15 2 15 15 1 15 13 2
11 13 3 7 9 9 0 9 1 0 9 2
36 13 15 15 1 9 7 9 0 1 0 9 2 1 9 0 9 16 0 0 9 11 2 2 13 9 9 11 11 1 9 1 11 1 9 12 2
5 0 9 13 0 9
2 11 2
23 0 9 13 3 0 0 9 9 7 9 0 9 9 9 0 9 11 11 1 9 0 9 2
30 0 9 9 13 1 9 9 10 0 0 9 1 12 9 9 11 11 7 10 9 1 9 12 9 0 0 9 11 11 2
11 9 0 9 13 1 11 11 9 11 11 2
16 3 16 11 11 13 15 11 11 13 10 9 14 1 9 12 2
7 11 13 9 0 0 9 2
21 1 10 9 13 10 0 0 9 9 0 9 11 11 2 15 3 1 9 11 13 2
24 15 1 9 13 3 3 1 9 7 1 0 9 2 3 13 11 9 2 15 1 9 9 13 2
17 1 9 12 15 13 1 15 2 16 4 1 11 11 3 3 13 2
4 13 9 11 11
2 11 2
22 1 9 12 9 13 1 10 9 1 11 1 0 11 0 0 9 7 0 9 11 11 2
20 10 9 1 9 0 9 4 13 1 10 9 7 13 15 9 1 9 0 9 2
1 3
17 1 12 9 13 11 10 0 9 7 1 9 3 13 9 0 9 2
27 1 9 12 4 13 9 9 9 11 0 7 10 0 9 0 0 11 7 15 13 0 9 9 9 1 11 2
34 0 9 9 11 2 11 1 9 13 2 16 13 1 9 13 1 11 9 1 9 0 9 2 16 4 13 10 0 9 0 9 1 11 2
10 9 15 13 9 3 16 12 9 9 2
8 11 2 11 15 13 1 12 9
2 11 2
25 0 9 0 9 7 0 9 11 2 11 4 1 0 9 13 1 12 0 9 11 11 7 11 11 2
10 12 0 9 4 3 13 0 9 9 2
28 9 9 13 9 1 0 9 9 7 9 9 12 9 1 9 0 9 16 1 9 0 9 2 7 7 1 9 2
14 0 9 13 15 2 16 11 15 13 3 0 16 11 2
12 10 9 1 9 11 2 11 3 13 12 5 2
22 11 11 4 13 9 11 0 11 2 11 11 2 11 0 11 2 11 11 7 11 11 2
19 1 12 9 3 13 11 9 12 9 0 9 2 9 2 12 9 9 2 2
16 11 16 9 0 9 7 9 13 1 12 9 9 12 9 9 2
21 12 0 9 9 11 2 11 1 9 0 9 11 11 4 13 4 13 1 9 9 2
8 9 11 11 13 0 0 11 2
4 9 9 15 13
8 11 13 1 12 0 9 11 2
3 0 9 9
2 11 2
28 0 9 0 9 1 9 1 0 9 14 1 0 9 3 1 11 13 11 11 11 2 0 0 9 9 1 11 2
8 1 0 9 13 9 11 12 2
19 13 3 9 1 0 9 2 16 13 0 2 7 1 0 2 0 2 9 2
17 10 0 9 13 13 9 2 7 3 1 0 0 9 13 9 9 2
20 10 0 9 11 12 13 9 11 1 9 1 9 9 1 9 1 0 9 9 2
10 1 9 13 9 13 12 7 12 9 2
17 1 15 0 2 15 13 3 1 9 1 9 9 2 13 11 0 2
12 1 0 9 13 3 13 1 0 9 7 9 2
11 0 0 9 13 13 9 14 1 12 9 2
23 3 0 9 0 9 11 15 3 1 9 0 9 7 9 1 9 12 3 13 1 0 9 2
16 1 0 9 15 13 1 9 13 15 1 0 12 9 1 9 2
19 1 0 9 7 1 11 13 10 9 1 9 12 13 9 3 12 0 9 2
12 1 0 0 9 13 1 10 9 3 13 9 2
7 9 13 13 1 11 10 9
2 11 2
28 0 9 9 0 9 13 1 11 13 10 9 2 13 3 1 9 10 10 9 1 11 11 10 0 9 11 11 2
28 7 13 9 1 9 9 2 16 9 1 9 0 11 2 3 13 0 9 1 0 9 2 13 13 3 0 9 2
23 9 9 11 11 13 2 16 9 1 9 4 13 1 9 9 2 9 7 9 1 10 9 2
12 11 0 4 0 0 9 13 9 9 1 9 2
19 11 13 2 16 11 3 13 7 13 12 0 9 7 1 12 9 0 9 2
6 3 13 14 12 9 2
20 1 11 15 13 7 1 9 1 9 0 9 2 0 12 9 3 15 4 13 2
20 11 13 9 0 9 9 11 2 11 7 11 2 3 9 1 11 10 9 13 2
10 11 2 13 9 11 1 9 11 2 2
24 10 9 13 0 0 9 2 15 13 1 9 1 0 9 2 16 9 11 13 9 1 15 13 2
11 15 1 11 13 2 16 3 4 3 13 2
15 13 15 3 13 1 0 9 2 15 13 11 1 11 13 2
15 11 13 1 12 0 9 2 15 13 9 1 9 12 9 2
24 1 11 11 2 15 0 9 3 13 2 4 1 9 9 9 13 9 9 0 9 1 0 9 2
14 11 3 13 3 9 2 9 0 9 13 13 0 9 2
13 16 4 11 13 9 2 13 4 10 9 14 3 2
33 1 0 9 1 11 15 9 13 13 2 3 13 9 13 1 15 2 16 4 1 0 9 13 9 0 9 1 9 0 0 0 9 2
5 0 9 1 0 9
2 11 2
16 0 9 1 9 7 9 13 1 0 9 13 2 0 2 9 2
25 1 9 0 9 0 11 4 10 9 13 13 3 0 0 9 1 9 1 9 9 1 9 0 9 2
21 9 13 14 12 7 12 9 0 0 9 13 2 0 2 0 9 7 13 10 9 2
20 13 1 15 2 16 10 9 13 9 1 9 0 9 7 10 9 3 9 9 2
25 9 9 13 1 0 2 16 1 0 9 13 0 0 9 7 4 15 13 1 0 9 1 10 9 2
24 7 3 2 16 15 9 13 7 13 1 0 9 2 4 10 9 13 3 1 9 10 0 9 2
20 0 9 1 9 7 9 1 10 0 9 13 0 9 1 9 9 7 0 9 2
12 0 9 0 9 13 13 14 12 9 2 9 2
6 1 11 15 13 0 9
6 0 9 13 1 0 11
2 11 2
20 0 0 11 7 0 11 0 1 11 1 9 3 13 10 0 0 9 1 11 2
29 9 11 2 0 11 2 11 2 11 2 0 2 4 13 0 9 12 9 9 2 12 9 15 1 9 13 0 9 2
17 9 4 13 12 9 2 15 4 13 0 9 9 1 9 7 9 2
24 1 9 13 13 0 0 9 2 0 9 1 0 9 7 0 9 0 2 0 7 0 0 9 2
15 9 13 3 0 1 0 9 2 9 0 9 7 9 9 2
10 11 7 0 11 3 13 3 10 9 2
16 10 9 13 13 1 0 9 1 11 2 11 2 11 7 11 2
6 9 11 13 0 9 11
2 11 2
18 0 9 11 15 13 1 9 0 9 9 0 9 1 0 9 9 11 2
22 1 0 0 9 1 15 13 0 9 9 11 11 11 7 9 0 9 9 11 11 11 2
28 9 13 13 1 0 9 9 1 9 1 0 0 9 2 9 1 15 7 1 9 1 0 9 0 7 0 9 2
29 9 10 9 2 15 4 13 3 13 9 9 2 13 13 1 3 12 9 7 10 9 13 1 12 1 12 9 9 2
23 9 9 11 13 1 11 13 1 0 9 11 11 11 2 9 11 2 9 11 7 9 11 2
4 3 13 0 9
4 1 9 0 9
10 9 11 13 13 0 9 1 0 9 2
19 1 0 9 10 9 1 9 15 1 0 9 13 2 16 13 13 0 9 2
12 15 15 9 11 13 1 0 9 15 0 9 2
23 9 9 13 1 9 12 9 2 12 9 9 13 9 9 1 9 2 3 2 0 9 2 2
25 1 1 15 2 16 0 9 3 13 9 1 9 7 9 0 9 2 0 9 9 13 3 0 9 2
32 3 15 13 0 9 2 1 15 13 1 0 9 9 13 9 9 0 9 7 9 9 0 9 1 9 2 16 4 9 13 9 2
23 9 13 3 0 13 1 0 9 9 9 0 9 2 3 16 9 9 9 1 9 9 9 2
29 3 0 9 13 9 1 0 9 2 16 4 9 13 9 1 9 7 16 3 1 0 9 13 9 1 9 10 9 2
21 1 0 9 13 0 3 9 1 9 9 1 9 7 3 7 1 9 0 9 9 2
20 1 0 9 13 9 0 13 2 10 9 7 9 9 13 1 9 9 0 9 2
39 1 0 9 15 13 15 0 9 9 2 9 9 2 0 7 0 0 9 2 9 0 9 2 9 2 1 15 4 9 13 1 0 9 7 10 0 0 9 2
26 0 0 9 1 0 9 13 9 1 15 2 16 13 9 9 1 9 2 15 4 13 9 7 0 9 2
22 1 15 13 0 9 13 7 9 1 0 9 1 9 2 16 13 9 2 9 7 9 2
16 0 9 13 1 10 9 13 7 13 9 0 9 15 15 13 2
8 13 15 13 15 7 10 9 2
11 10 9 13 1 0 9 13 3 0 9 2
36 1 15 13 9 13 7 0 9 13 0 15 9 13 1 12 9 1 9 2 3 1 15 9 13 2 7 14 3 16 12 9 1 9 0 9 2
22 9 0 9 13 13 3 9 1 9 2 9 7 0 9 2 15 13 9 1 9 9 2
11 0 9 13 9 13 13 3 1 9 9 2
9 9 1 9 13 4 3 1 11 9
2 11 2
13 1 0 9 15 1 11 3 3 16 13 9 9 2
27 0 9 9 1 9 13 12 1 0 9 0 0 9 2 1 15 3 13 1 9 7 9 10 0 0 9 2
11 9 1 15 1 3 12 9 9 3 13 2
7 10 0 9 13 0 9 2
25 1 9 12 13 1 11 12 9 2 0 9 3 12 7 1 9 12 13 9 9 1 9 12 9 2
10 3 13 1 0 9 9 12 9 9 2
17 0 3 0 9 0 9 13 12 9 2 7 1 9 13 3 0 2
41 9 0 9 13 9 11 0 1 12 9 2 9 2 2 1 15 4 13 2 0 0 9 2 1 0 9 2 7 7 0 9 7 3 3 0 2 15 4 13 13 2
10 10 9 13 14 12 9 9 9 11 2
18 3 0 0 9 15 1 9 12 13 9 0 9 7 9 1 12 9 2
21 1 9 9 13 0 9 9 12 5 2 15 13 1 0 9 12 1 0 9 9 2
11 0 9 3 13 9 2 16 13 1 9 2
3 9 2 9
23 9 9 0 7 0 9 1 9 12 2 9 13 9 2 3 13 0 0 9 1 9 9 2
33 9 9 13 13 9 3 1 9 1 12 9 2 1 9 1 9 9 2 7 1 9 1 12 9 2 1 9 3 0 0 9 2 2
15 0 9 13 13 1 9 9 1 9 7 1 0 0 9 2
13 9 7 9 9 2 12 2 9 1 11 1 11 2
28 13 2 9 9 11 2 0 12 2 12 12 11 1 11 2 9 2 2 12 2 12 2 9 2 12 2 12 2
9 9 0 9 1 9 9 7 9 2
19 9 15 13 9 0 9 2 0 9 9 7 13 0 9 1 9 0 9 2
12 9 7 9 9 2 12 2 12 2 1 11 2
34 13 2 11 2 0 12 2 11 12 2 9 2 2 12 2 12 2 2 12 2 12 2 9 2 2 12 2 12 2 2 12 2 12 2
31 0 9 9 1 9 0 9 2 0 9 9 1 9 0 9 2 0 9 9 2 12 0 9 2 15 13 0 9 0 9 2
15 9 7 9 9 2 12 2 2 12 2 7 12 2 12 2
4 13 2 11 2
4 9 0 9 2
12 9 7 9 9 2 12 2 12 2 1 11 2
4 13 2 11 2
7 0 9 2 0 0 9 2
15 9 7 9 9 2 12 2 2 12 2 12 2 1 11 2
4 13 2 11 2
6 0 9 1 11 3 13
2 11 2
24 1 9 9 9 7 0 9 13 1 0 12 2 9 12 9 9 1 0 9 3 12 0 9 2
12 1 9 1 9 12 13 1 9 1 12 9 2
13 0 9 9 1 9 9 15 7 1 9 13 3 2
17 1 9 0 9 13 9 9 1 12 9 0 16 3 1 0 9 2
24 3 15 1 9 0 9 1 9 9 13 12 9 2 15 13 1 12 3 16 1 0 0 9 2
11 1 9 0 9 4 13 12 9 1 9 2
17 1 12 2 9 12 13 9 9 1 0 9 3 12 0 0 9 2
10 1 9 13 1 12 0 9 12 9 2
5 0 9 1 0 9
2 11 2
21 1 12 9 13 1 0 9 0 2 2 0 9 2 0 0 0 9 1 0 9 2
29 1 9 0 9 13 9 0 9 1 9 1 9 0 9 1 9 2 0 9 2 9 7 0 9 7 0 0 9 2
13 9 9 13 13 1 9 0 9 7 9 1 9 2
25 9 15 1 0 9 13 16 0 9 0 9 2 0 7 0 9 2 9 0 9 7 1 0 9 2
10 3 4 13 13 3 13 13 0 9 2
16 1 0 9 15 0 9 13 0 9 3 1 10 3 0 9 2
15 15 15 13 1 0 9 2 10 9 13 3 9 0 9 2
5 11 13 7 0 9
12 0 9 13 9 3 1 3 16 12 9 1 11
2 11 2
16 0 9 11 13 1 9 0 9 12 9 9 0 9 0 11 2
17 1 0 9 12 9 0 9 15 3 13 0 0 9 0 0 9 2
24 1 0 9 13 9 11 1 9 12 1 11 2 15 3 13 1 9 0 9 13 16 3 0 2
20 1 0 9 13 9 9 1 3 16 12 0 2 0 7 0 9 1 0 9 2
8 3 9 9 3 13 12 9 2
19 9 13 1 0 0 9 3 0 7 0 9 2 0 9 0 7 0 9 2
8 0 9 3 13 1 9 9 2
9 9 9 13 1 9 0 0 9 2
18 9 11 13 0 9 2 0 9 2 9 2 9 2 9 7 0 9 2
35 13 1 15 3 0 9 11 2 0 9 2 9 9 2 0 9 1 11 2 0 9 1 11 2 0 9 11 2 0 9 11 7 0 9 2
8 9 11 13 1 9 0 9 2
21 13 15 2 16 9 1 9 13 1 9 0 9 0 2 16 9 13 12 5 9 2
17 9 1 11 13 0 1 9 2 15 13 9 1 2 0 2 9 2
10 0 9 13 3 9 9 1 0 9 2
9 1 0 9 9 11 13 9 11 2
18 9 1 10 9 13 0 9 0 9 0 9 2 9 7 0 9 9 2
21 3 15 13 2 13 15 2 16 1 9 11 15 3 13 7 13 2 7 13 9 2
2 1 9
2 11 2
21 1 9 0 9 13 9 9 1 9 11 12 5 2 15 13 12 0 9 1 9 2
7 1 10 9 13 12 9 2
29 1 0 9 0 9 13 0 0 9 12 9 1 9 2 12 9 2 2 1 15 9 13 3 16 9 2 12 2 2
23 1 0 9 0 9 13 1 9 9 9 1 11 12 9 2 1 0 9 15 13 12 9 2
15 9 0 9 15 13 1 12 1 9 12 1 0 12 9 2
7 3 9 1 9 13 0 2
17 1 9 12 13 0 9 9 12 0 9 2 1 0 0 9 12 2
3 0 11 2
27 9 9 1 0 9 13 1 9 0 9 9 1 9 0 9 1 12 5 2 15 13 3 12 9 1 9 2
16 9 13 3 13 9 7 9 0 11 2 11 2 11 7 11 2
9 1 9 1 9 13 9 7 9 2
2 11 2
14 9 9 1 0 9 13 1 0 12 2 9 12 5 2
23 9 9 1 11 1 10 9 13 12 0 2 1 15 12 9 7 12 9 1 0 0 9 2
16 1 0 9 13 1 9 12 9 1 9 2 13 15 4 12 2
9 0 9 9 13 9 2 12 2 2
15 1 9 13 3 12 0 9 7 12 0 9 15 9 9 2
9 0 9 9 13 3 12 0 9 2
9 9 15 13 13 1 12 0 9 2
10 1 0 7 0 9 13 12 0 9 2
11 9 1 0 0 9 13 13 12 0 9 2
18 9 11 1 11 13 3 3 1 12 9 9 2 15 15 13 1 9 9
4 0 9 13 9
8 9 13 1 9 2 7 1 9
11 9 1 9 15 13 9 9 7 9 1 9
11 9 9 3 13 7 10 0 9 7 9 2
26 15 15 3 9 1 0 9 13 2 7 13 15 2 16 4 15 15 1 10 0 9 7 0 9 13 2
19 0 9 13 13 9 2 16 15 13 15 9 1 0 9 1 15 1 9 2
12 3 0 0 9 9 0 9 13 9 0 9 2
17 3 13 1 9 0 9 2 9 2 9 2 2 2 2 7 9 2
16 9 13 13 9 2 0 9 2 9 2 9 0 7 0 9 2
9 1 9 9 15 9 13 10 9 2
23 9 1 9 10 9 15 13 0 9 9 3 2 13 15 0 9 9 7 3 9 0 9 2
19 0 9 1 10 9 15 13 1 11 2 7 0 13 7 1 0 0 9 2
13 3 1 0 9 13 9 0 9 1 9 10 9 2
26 9 1 0 9 13 9 1 9 9 1 9 9 2 1 15 13 0 9 7 13 10 9 1 0 9 2
20 16 13 13 9 1 9 3 0 9 2 13 9 1 0 9 13 3 10 9 2
18 9 16 3 1 0 2 0 7 0 9 13 0 13 16 9 1 9 2
5 10 9 15 13 2
10 9 15 13 3 3 13 7 13 0 2
17 0 9 15 13 7 9 1 15 13 3 15 2 15 13 9 9 2
12 0 9 9 9 9 13 1 12 7 12 9 2
19 9 1 9 9 4 9 3 13 13 0 9 2 7 15 13 3 9 9 2
32 1 9 13 3 0 3 13 0 9 1 9 1 0 9 2 13 2 16 0 9 9 13 0 9 2 1 15 15 9 3 13 2
15 0 9 3 13 0 13 9 9 2 9 7 0 0 9 2
15 1 9 9 0 9 13 13 16 1 9 2 7 7 9 2
16 10 9 13 9 7 1 9 0 9 2 15 13 9 0 9 2
21 1 9 9 4 15 13 1 10 3 0 9 2 15 15 13 1 9 2 9 2 2
9 0 9 13 13 9 1 12 9 2
12 3 15 1 9 9 13 1 9 11 7 11 2
12 9 1 0 9 0 1 0 9 13 3 0 2
20 1 9 1 9 9 12 5 12 9 7 9 12 9 13 9 1 9 12 9 2
16 16 15 9 10 9 13 1 12 9 2 9 13 1 12 9 2
23 1 0 9 2 3 2 1 9 9 5 12 12 9 7 9 12 9 3 13 12 9 3 2
14 1 9 9 1 0 9 13 9 13 3 1 12 9 2
7 9 1 15 13 3 0 2
22 1 9 12 5 12 5 12 9 13 12 9 1 9 2 1 0 9 9 13 7 9 2
11 1 9 12 9 10 9 13 3 12 9 2
13 9 0 9 13 13 1 12 9 1 9 0 9 2
8 10 9 15 9 13 1 9 2
45 9 13 12 0 9 2 1 15 0 2 12 5 2 13 0 0 9 1 12 9 2 9 12 2 7 3 2 9 12 5 12 5 12 9 2 2 1 15 0 9 13 3 12 9 2
14 1 0 2 3 0 9 13 9 13 7 9 0 9 2
8 9 1 10 9 15 13 3 2
34 3 16 12 9 9 13 11 2 15 13 9 1 11 1 11 2 11 2 11 11 2 0 9 2 11 2 0 11 2 11 7 1 11 2
11 9 13 3 0 16 3 2 1 0 9 2
11 1 9 1 9 12 9 12 13 9 12 9
17 12 9 7 1 10 0 9 1 9 12 9 12 3 12 9 3 2
20 0 9 3 13 1 3 0 9 1 0 11 7 11 9 1 11 1 0 9 2
12 9 9 15 3 1 9 9 11 11 13 13 2
46 0 9 3 13 10 9 13 1 9 9 12 5 12 5 12 9 2 7 2 3 12 9 12 2 1 0 9 12 9 2 7 1 9 12 9 1 12 9 7 9 12 9 1 12 9 2
10 1 9 0 9 13 9 9 3 9 2
19 10 9 9 15 13 9 9 2 1 12 9 1 9 15 13 12 9 3 2
15 1 9 12 9 9 13 3 12 9 2 1 12 12 9 2
19 9 9 15 1 0 9 13 13 1 12 1 12 0 9 0 9 1 9 2
17 9 12 5 12 9 13 9 9 12 2 12 2 12 7 12 9 2
12 0 13 1 12 9 7 0 1 12 9 3 2
12 3 13 9 1 0 9 9 12 7 12 9 2
7 0 9 9 13 9 11 2
20 1 0 9 12 5 12 9 15 13 13 9 12 2 12 2 12 7 12 9 2
14 1 0 9 9 13 9 1 15 0 16 1 0 9 2
23 1 0 0 9 13 9 12 9 7 9 12 9 3 2 1 0 12 3 12 9 1 9 2
36 1 0 7 0 9 2 3 15 13 7 10 9 2 15 13 9 13 3 0 9 1 9 2 15 15 13 1 9 9 14 1 0 9 12 9 2
22 0 7 0 9 13 1 9 1 0 9 12 9 2 10 9 15 3 13 1 12 13 2
23 0 12 9 1 9 12 5 12 9 7 9 12 2 12 7 12 9 13 1 9 12 9 2
22 1 9 12 9 13 12 9 2 1 12 9 12 9 7 1 12 9 12 9 1 9 2
7 0 0 4 13 12 9 2
16 0 9 15 13 1 10 9 9 13 0 9 1 11 1 11 2
13 9 9 13 13 12 9 0 1 12 1 12 9 2
33 13 0 9 1 15 1 9 11 2 0 0 9 7 0 0 7 0 9 13 1 9 10 9 0 2 7 15 13 1 9 10 9 2
15 13 2 16 15 13 9 7 13 1 9 15 0 7 0 2
31 3 3 2 16 15 13 9 2 1 0 3 13 2 2 15 3 1 9 13 2 3 1 9 9 2 3 1 9 9 11 2
6 3 1 9 16 1 9
15 1 9 15 13 3 13 10 9 2 13 7 3 3 13 9
27 1 0 9 1 11 11 9 0 9 13 1 9 9 2 16 4 1 9 1 15 13 0 9 7 0 9 2
13 9 11 11 13 15 3 2 7 9 9 13 9 2
8 3 3 9 13 3 15 13 2
19 0 9 7 7 0 9 13 1 9 3 13 15 12 2 7 3 13 9 2
22 13 13 0 9 0 1 9 9 2 3 16 0 9 2 1 15 13 9 7 0 9 2
40 16 13 9 3 1 9 2 9 13 9 2 13 0 2 2 13 0 13 2 15 13 1 9 13 2 16 0 9 2 9 2 9 2 0 9 2 9 2 2 2
20 15 13 13 2 3 0 0 9 13 2 16 13 0 9 7 3 0 0 9 2
23 0 9 15 13 3 9 2 15 13 13 0 9 2 7 1 9 13 13 9 3 7 9 2
19 1 9 9 13 13 9 7 9 1 12 9 2 3 0 9 13 0 9 2
21 7 12 9 2 1 0 9 7 9 2 15 15 1 15 13 13 2 13 0 9 2
29 13 1 9 0 9 2 7 3 1 15 2 16 9 13 9 2 9 2 2 3 0 0 9 0 3 1 0 9 2
23 1 9 15 9 2 15 13 1 9 1 9 7 0 9 2 13 1 0 7 0 1 9 2
15 0 9 13 0 0 9 1 9 2 15 15 13 1 9 2
18 16 4 13 16 3 0 9 2 13 15 1 9 2 3 1 0 9 2
30 0 0 9 1 9 1 12 9 2 10 9 1 9 1 12 9 13 0 9 2 13 0 13 2 3 15 13 1 9 2
24 1 0 9 2 3 1 9 2 15 13 13 16 0 9 9 2 13 0 9 3 3 1 9 2
24 9 1 9 13 0 0 7 0 9 2 15 13 1 9 2 7 3 15 13 3 13 1 9 2
16 9 9 3 13 13 9 9 2 16 4 0 9 13 1 9 2
21 1 0 9 15 13 1 0 9 2 3 15 10 9 3 1 9 13 1 0 9 2
37 3 1 0 9 1 9 0 9 2 1 0 9 1 0 9 14 12 5 12 5 12 9 2 0 9 3 12 9 2 13 9 9 1 3 12 9 2
10 9 10 9 15 13 12 9 1 9 2
24 9 1 9 1 0 9 12 5 12 5 12 9 2 0 9 12 9 2 13 9 14 12 9 2
5 13 1 12 9 2
14 3 1 9 9 13 2 16 1 12 15 15 3 13 2
15 12 9 13 13 0 9 7 0 9 15 13 1 0 9 2
15 16 15 9 9 13 13 1 9 2 13 13 0 0 9 2
22 1 0 9 15 7 13 7 3 13 13 9 9 1 0 9 2 13 1 0 9 2 2
7 1 15 13 3 1 9 2
27 3 16 9 1 0 9 13 9 7 13 15 0 9 7 1 9 2 12 9 13 13 7 9 0 9 3 2
7 3 3 13 3 13 9 2
11 13 15 3 1 9 2 16 15 9 13 2
44 16 13 9 0 9 2 13 15 1 9 2 15 15 1 0 0 9 13 10 9 1 9 2 3 3 1 10 9 7 0 9 2 0 9 13 3 1 9 1 12 2 9 2 2
19 15 13 3 9 9 9 1 10 9 2 13 14 1 12 1 3 12 9 2
11 3 13 1 9 3 3 2 0 0 9 2
7 9 13 1 0 9 9 2
13 10 9 13 13 3 14 15 2 16 13 3 1 9
6 9 9 3 13 12 9
2 11 2
11 7 16 13 3 9 2 13 13 3 13 2
26 13 15 13 1 9 7 13 2 16 9 2 15 4 15 3 3 13 1 9 2 13 3 7 1 15 2
19 1 0 0 9 4 1 0 9 13 12 9 1 0 9 0 12 9 9 2
20 9 1 9 15 1 10 9 13 3 12 9 7 9 1 0 9 3 12 9 2
11 13 4 12 1 15 2 3 0 12 9 2
12 0 3 13 3 9 1 9 0 12 9 9 2
28 7 16 15 9 9 1 9 12 13 1 3 16 12 9 7 9 13 1 12 2 9 13 0 1 3 16 9 2
5 9 0 9 13 0
16 16 4 13 0 2 13 13 3 9 9 2 9 7 0 9 2
13 13 9 7 0 2 3 0 9 2 9 2 9 2
11 7 15 13 13 2 9 0 2 1 9 2
12 9 10 9 13 0 9 1 9 0 0 9 2
29 1 0 9 2 15 15 13 1 12 9 2 15 9 13 1 12 9 0 9 3 2 7 1 12 9 14 12 9 2
22 1 0 9 9 2 1 0 7 0 9 2 13 9 1 12 9 0 9 1 12 9 2
22 9 15 3 13 3 12 5 9 1 0 9 1 9 1 0 9 2 15 13 13 9 2
5 9 13 0 1 9
10 9 9 9 7 9 4 13 1 0 9
2 11 2
22 1 9 0 9 4 13 4 13 0 9 12 9 9 0 0 7 0 9 9 7 9 2
12 3 1 11 15 13 9 9 0 9 11 11 2
31 1 15 15 3 13 3 1 9 0 9 10 9 2 16 9 7 9 2 15 3 13 10 9 2 4 3 13 4 13 9 2
12 0 9 4 15 13 13 14 12 9 7 9 2
37 1 9 9 1 0 11 7 1 11 11 13 2 16 9 0 9 13 9 9 0 9 7 3 3 13 4 13 0 9 1 9 12 9 9 10 9 2
10 9 1 0 9 4 13 13 0 9 2
21 1 9 9 0 9 11 7 0 9 15 0 9 3 13 2 13 7 9 3 13 2
22 1 11 2 11 13 0 2 16 4 1 9 9 13 15 0 0 9 9 1 0 9 2
9 11 1 11 13 3 0 9 11 2
15 1 9 13 10 9 1 11 12 7 13 1 0 0 9 2
20 13 12 9 2 15 13 0 9 7 9 7 13 9 1 9 7 9 0 9 2
8 0 9 9 9 1 9 1 9
2 11 2
31 9 1 9 12 9 9 13 9 1 0 9 11 11 9 9 11 11 7 9 0 11 1 0 9 0 9 1 9 0 9 2
23 9 1 11 2 11 13 2 16 0 9 12 9 15 13 1 9 1 0 9 9 0 9 2
23 9 9 13 0 9 9 2 7 9 0 9 1 12 0 9 1 0 9 3 13 0 9 2
18 0 9 13 9 3 1 9 1 9 9 0 0 9 1 0 9 9 2
18 9 3 13 9 9 11 11 1 0 9 9 1 9 9 12 9 9 2
48 10 9 13 2 16 1 1 10 0 9 13 1 0 0 9 2 11 11 13 0 9 0 9 11 0 0 11 2 15 3 13 12 9 9 9 11 11 2 2 7 7 13 13 10 0 0 9 2
27 9 13 7 9 0 0 9 2 15 4 1 0 9 9 13 9 12 12 9 1 9 1 9 0 0 9 2
13 9 3 13 2 16 1 10 9 15 0 9 13 2
20 12 0 9 13 0 13 9 1 12 9 2 3 3 15 13 13 1 0 9 2
6 11 11 9 1 12 9
3 0 11 2
30 1 3 16 9 15 3 0 9 0 9 0 9 2 11 11 2 13 1 9 9 12 12 9 2 13 9 0 11 9 2
24 7 14 1 12 9 1 0 12 9 15 15 1 9 10 9 13 13 2 16 13 1 12 9 2
17 3 15 10 9 13 1 12 3 1 0 9 9 0 1 9 9 2
24 13 15 9 9 2 15 13 2 16 15 0 0 9 13 13 9 0 9 7 3 15 13 0 2
10 3 9 9 9 13 1 11 1 9 2
13 3 3 13 1 0 9 9 1 0 9 9 9 2
16 1 9 9 4 13 0 0 9 12 12 9 13 1 9 12 2
7 11 3 1 9 12 9 9
2 11 2
22 11 2 0 0 0 9 13 1 0 9 1 12 2 9 12 9 1 9 12 9 9 2
18 0 9 9 13 1 10 9 12 9 9 2 15 13 12 9 1 9 2
28 1 12 2 12 2 12 15 11 2 0 0 2 0 0 2 0 0 7 0 0 0 9 13 1 0 0 11 2
29 0 9 9 11 2 0 0 11 13 1 12 2 9 12 9 9 2 3 12 9 1 9 7 12 9 1 0 9 2
13 9 12 9 13 1 0 9 12 2 9 12 9 2
1 3
25 0 0 9 13 1 9 9 2 15 13 0 9 9 13 9 0 9 0 9 7 10 9 1 11 2
20 0 9 3 13 9 2 15 13 1 9 0 9 1 0 9 9 3 1 9 2
13 3 7 10 9 2 16 3 0 9 2 4 13 2
5 11 9 1 0 11
2 11 2
22 9 11 2 15 13 0 9 11 3 1 0 0 11 2 15 13 1 9 1 11 11 2
12 11 13 12 1 0 0 0 9 0 0 9 2
14 1 10 9 4 1 0 9 13 1 0 9 1 11 2
9 0 9 13 0 0 9 1 11 2
25 10 9 1 12 9 13 0 0 9 1 0 11 7 13 1 0 0 9 1 12 9 0 0 9 2
8 1 0 9 15 13 0 9 2
8 13 15 9 12 0 9 0 9
4 9 1 11 2
19 9 12 0 9 0 0 9 13 13 1 0 1 9 9 9 1 0 9 2
14 13 1 0 2 0 0 9 2 9 0 7 9 0 2
18 1 9 1 9 0 9 15 13 1 9 11 11 1 9 9 0 9 2
29 0 0 9 2 3 0 0 9 4 13 13 3 12 0 9 7 10 9 4 13 1 9 11 2 11 2 0 2 2
12 13 4 15 7 3 2 9 9 9 1 9 2
21 1 9 0 2 15 4 13 3 0 2 4 13 13 9 3 1 9 0 0 9 2
44 9 0 4 13 3 0 9 2 3 2 12 7 12 9 2 2 15 4 7 3 13 1 9 9 2 7 15 13 3 2 16 15 3 13 9 1 0 9 2 13 11 2 11 2
17 1 11 13 1 9 12 0 9 2 12 0 9 7 12 0 9 2
10 1 0 0 9 15 13 3 3 12 2
21 1 9 15 1 9 0 9 13 0 9 3 0 9 7 9 2 13 11 2 11 2
5 9 12 1 0 9
2 11 2
40 9 12 3 0 9 9 13 3 1 11 0 9 2 1 15 15 1 9 1 9 0 0 9 13 13 2 3 7 10 9 15 13 9 13 1 2 0 9 2 2
22 13 15 3 2 16 1 0 7 0 9 0 9 0 1 0 9 15 13 0 0 9 2
25 0 9 15 13 2 16 9 9 2 0 9 7 9 15 13 1 2 0 9 1 12 2 9 2 2
28 0 9 9 9 12 4 3 13 13 9 9 1 0 9 2 15 13 9 7 9 9 0 9 13 0 0 9 2
6 1 9 9 15 13 9
8 9 0 9 13 9 13 0 9
8 1 0 2 9 13 13 1 9
3 1 0 9
16 0 9 2 9 9 2 11 2 12 2 9 2 11 11 2 2
27 0 7 0 9 1 9 2 9 2 9 7 0 9 0 9 2 15 3 9 3 13 16 2 9 9 2 2
6 1 0 9 11 11 2
8 9 1 11 2 11 0 11 2
2 0 9
19 0 9 11 13 10 0 9 2 9 9 11 2 7 15 13 13 10 9 2
11 0 11 15 9 13 13 3 1 0 9 2
34 7 15 13 0 9 11 2 16 4 0 11 13 7 13 15 9 2 16 13 2 16 15 1 15 0 9 1 0 9 1 9 3 13 2
17 7 11 13 0 9 10 9 7 1 0 11 15 3 13 2 2 2
40 2 0 9 1 0 9 2 13 1 0 9 0 9 10 9 7 1 0 9 15 13 9 0 9 2 13 2 16 0 11 13 1 9 9 9 1 0 9 2 2
51 3 0 0 9 1 9 2 9 7 9 13 1 0 9 9 16 3 0 7 0 9 2 16 15 10 9 1 3 0 0 9 3 3 13 0 9 7 9 2 16 9 13 0 9 9 2 1 15 13 13 2
8 12 1 9 2 11 2 12 2
8 9 1 11 2 11 0 9 2
5 9 2 11 11 2
13 13 2 11 11 2 11 11 2 11 11 7 0 2
5 0 9 1 0 9
35 0 0 0 7 0 9 1 11 1 9 0 9 11 2 9 0 11 7 0 9 9 2 0 0 11 2 3 0 9 1 0 9 3 13 2
26 1 0 9 9 13 0 7 0 0 11 2 7 15 14 3 2 16 13 0 13 1 9 1 0 9 2
39 9 0 9 0 11 15 13 1 0 0 9 2 1 9 0 9 2 0 9 2 1 9 3 0 9 9 9 14 1 9 1 9 2 9 2 2 3 2 2
45 16 9 1 15 13 1 0 2 13 15 9 11 11 1 12 9 3 2 13 2 9 2 15 3 13 13 1 10 9 1 0 9 9 0 12 9 2 2 13 2 7 2 13 2 2
25 1 0 9 10 3 0 9 15 7 13 15 9 2 15 1 9 9 0 11 13 13 9 0 11 2
17 3 9 15 3 13 7 1 0 9 9 2 13 14 0 2 15 2
22 7 3 13 9 9 1 9 0 9 1 9 0 9 7 0 9 0 9 0 9 9 2
29 9 0 9 0 11 2 0 1 0 9 2 13 3 1 0 9 7 1 3 16 0 9 13 9 3 0 10 9 2
41 13 9 1 0 9 2 3 9 13 1 0 9 2 2 15 3 13 1 9 15 0 9 2 0 9 1 9 13 15 9 14 1 9 0 9 1 0 9 0 9 2
54 0 11 13 3 0 9 2 1 15 15 15 12 9 1 9 9 7 0 9 9 3 2 13 2 1 0 9 0 9 1 0 11 2 1 0 9 1 0 9 7 0 0 9 2 1 15 4 13 7 9 2 2 2 2
24 9 2 0 0 9 15 9 9 1 3 0 9 2 15 13 3 9 14 1 0 9 0 9 2
35 16 3 16 0 7 0 9 9 13 0 11 0 9 9 2 1 15 3 13 1 9 0 9 9 2 2 13 15 1 0 9 3 13 3 2
8 0 11 2 0 11 2 11 2
11 11 2 0 9 1 9 2 12 2 9 2
7 13 9 12 2 12 11 2
3 9 9 0
30 16 9 9 0 9 1 0 9 2 9 7 0 9 3 2 4 3 1 11 13 2 3 13 1 9 9 2 3 2 2
11 13 0 2 0 2 0 9 2 0 11 2
17 9 11 11 13 10 2 9 2 2 7 15 3 1 9 11 11 2
33 13 2 2 3 15 13 13 2 13 9 14 0 9 2 7 3 0 9 2 7 10 9 13 3 10 9 2 1 15 9 13 2 2
24 13 3 11 11 16 9 7 11 11 16 11 2 1 9 9 1 15 13 3 0 11 11 11 2
11 13 15 3 16 0 9 16 16 10 9 2
35 7 16 11 10 9 13 2 0 9 14 13 1 0 9 1 9 12 2 3 13 0 11 11 0 0 11 7 11 11 13 0 7 0 11 2
21 1 0 9 13 1 9 12 9 12 9 2 0 2 11 2 7 0 2 11 2 2
38 16 0 9 4 1 12 9 13 3 2 11 11 13 11 3 1 12 1 15 2 2 11 11 15 3 13 13 1 0 9 11 11 7 10 0 0 9 2
18 16 0 11 2 7 0 11 13 9 9 9 11 2 3 14 1 11 2
8 9 9 13 9 0 9 0 2
22 11 2 11 11 2 7 11 2 11 11 2 15 13 3 0 7 13 4 3 10 9 2
23 1 12 9 15 9 3 13 11 11 2 11 2 2 13 13 3 9 11 11 2 11 2 2
12 11 11 2 11 2 14 13 0 9 1 0 2
29 15 2 15 15 13 2 1 10 9 4 13 1 9 1 0 9 0 9 2 13 3 13 0 9 9 1 10 9 2
23 9 13 10 9 2 7 1 10 9 4 9 7 13 2 9 13 7 1 9 9 0 9 2
34 11 11 13 14 9 7 11 11 16 11 2 11 11 13 0 2 13 15 9 0 11 11 2 11 2 7 0 9 11 11 2 11 2 2
23 0 9 15 1 15 13 1 11 0 11 2 0 9 7 9 0 9 1 0 9 11 11 2
42 2 7 3 3 13 2 9 9 2 11 11 7 11 11 2 15 13 1 12 9 3 9 0 9 2 11 4 15 13 3 13 2 2 2 9 9 2 3 0 0 9 2
14 0 0 9 2 0 7 0 2 0 7 0 2 2 2
39 1 0 9 15 10 9 13 3 3 2 2 15 3 14 13 9 2 2 13 4 4 2 15 3 14 13 9 2 2 3 7 2 15 4 3 13 9 2 2
16 13 15 9 2 15 13 3 10 11 2 15 15 13 13 3 2
14 16 13 0 2 16 11 15 13 9 1 9 9 9 2
26 1 12 9 15 3 3 0 9 9 13 13 15 3 3 3 3 2 16 13 14 13 2 7 7 13 2
21 7 1 0 9 15 9 13 1 9 0 9 11 2 0 15 13 9 11 7 11 2
17 0 9 11 11 15 13 2 16 0 9 1 9 13 0 1 9 2
12 13 7 14 9 0 0 9 2 15 15 13 2
12 3 13 13 9 1 15 2 16 11 3 13 2
22 14 14 3 15 15 13 10 0 9 1 10 9 2 14 2 3 15 9 15 13 2 2
21 11 7 11 13 1 15 2 7 15 3 0 9 2 15 10 9 13 7 13 13 2
5 0 9 1 15 0
27 9 1 9 2 15 15 13 0 9 2 13 3 13 1 9 2 16 1 10 9 13 10 9 1 10 9 2
22 9 9 0 9 11 11 7 13 2 16 15 10 9 13 3 13 2 0 13 9 9 2
17 1 9 1 0 9 9 9 12 13 1 9 11 13 10 0 9 2
10 13 15 2 16 13 1 9 0 9 2
8 9 13 1 10 9 10 9 2
12 3 15 13 9 2 15 15 13 0 9 13 2
29 3 4 13 0 9 2 3 9 1 9 1 9 2 9 11 1 11 7 1 11 7 0 9 1 11 7 1 11 2
14 0 9 13 9 16 9 2 9 7 9 1 11 11 2
23 9 15 3 3 7 3 13 1 0 9 1 9 7 13 9 1 10 9 2 9 7 9 2
12 3 13 1 0 9 16 9 9 2 9 9 2
25 3 16 15 9 13 1 10 9 2 4 13 13 1 0 7 0 9 2 16 13 3 9 1 9 2
14 10 9 13 1 10 9 9 9 9 2 9 7 9 2
30 11 13 0 9 2 13 3 13 2 7 3 13 10 9 1 9 1 0 9 2 3 15 9 13 2 3 1 0 9 2
8 11 15 3 13 3 1 9 2
22 1 9 15 3 13 3 2 9 1 15 13 2 7 2 1 9 15 13 2 2 2 2
5 15 13 3 9 2
14 0 9 13 13 3 1 9 9 1 9 7 1 9 2
9 9 1 0 9 13 3 0 9 2
11 3 13 15 0 9 9 2 15 13 9 2
15 13 15 3 9 7 9 2 1 15 9 1 9 3 13 2
7 13 9 1 0 0 9 2
23 1 11 13 1 9 9 0 9 1 9 2 15 15 1 10 9 13 1 0 2 0 9 2
17 1 15 10 4 15 10 9 0 13 2 7 9 3 3 13 13 2
8 10 9 9 11 13 3 0 2
23 3 15 13 9 11 11 2 7 15 15 13 13 15 2 16 9 13 0 7 13 0 9 2
17 15 15 13 2 16 0 13 9 11 11 0 9 2 9 11 11 2
20 13 15 0 9 0 9 7 9 1 9 9 2 10 0 2 0 7 0 9 2
9 1 10 9 13 1 9 10 9 2
7 3 13 3 14 3 0 2
18 9 9 11 13 13 1 9 9 0 9 2 7 13 7 1 0 9 2
20 9 1 0 9 1 0 9 13 13 9 2 15 13 2 16 0 9 13 9 2
37 1 0 9 13 3 0 2 16 15 3 13 2 16 15 3 14 13 1 0 9 2 1 9 0 2 0 2 1 9 0 7 1 0 9 7 9 2
17 0 1 0 9 1 9 13 3 0 9 1 15 0 2 1 9 2
12 9 9 0 9 1 11 7 9 9 11 11 11
5 9 11 11 2 11
5 9 2 9 7 9
52 1 9 11 11 9 9 2 9 7 9 2 13 11 2 13 9 0 9 2 15 11 11 2 12 2 2 9 0 9 1 9 2 0 9 7 0 9 0 9 0 1 9 2 13 1 11 7 1 10 0 9 2
56 13 1 15 1 0 9 0 9 2 11 2 11 7 11 2 11 2 11 2 11 2 11 2 11 2 16 9 9 0 9 2 13 10 9 1 10 9 2 1 9 9 2 15 13 11 2 2 7 0 9 15 13 1 9 2 2
8 0 9 13 1 9 11 11 2
16 16 9 4 13 10 0 9 1 9 2 15 15 13 1 9 2
10 13 4 15 11 1 9 7 13 4 2
12 13 4 11 2 9 11 2 7 13 4 15 2
6 3 15 1 15 13 2
9 13 1 9 2 16 4 15 13 2
32 16 13 3 9 16 15 0 2 13 10 9 0 9 2 7 9 0 9 1 0 2 3 7 3 0 9 2 15 13 10 9 2
21 4 15 13 13 10 9 1 9 0 7 0 9 2 16 4 15 3 13 1 9 2
4 9 11 9 0
10 13 15 0 9 2 1 15 13 9 2
4 9 7 9 2
4 9 7 9 2
4 9 7 9 2
30 1 0 10 9 15 10 9 13 9 9 1 15 2 15 15 13 1 15 7 13 15 3 2 13 1 15 10 0 9 2
26 13 15 9 2 1 15 13 13 0 9 1 0 10 9 2 3 16 9 13 9 2 1 15 15 13 2
73 13 1 15 15 0 9 2 15 9 7 15 3 15 0 9 9 2 0 9 2 9 9 9 1 9 9 2 10 9 9 7 9 2 10 9 1 0 9 7 0 9 2 1 9 13 9 7 9 13 2 9 1 9 7 9 1 9 2 9 13 9 7 9 9 7 9 2 0 9 7 0 9 2
4 13 3 15 2
20 3 15 9 10 9 2 0 7 0 2 0 1 9 9 9 2 15 13 9 2
44 0 10 9 13 1 9 2 13 9 7 9 7 13 0 9 2 13 15 3 1 9 7 13 1 9 2 16 4 3 13 1 0 9 2 15 13 9 0 0 9 2 0 9 2
13 9 0 0 9 7 13 0 9 0 2 3 0 2
15 10 0 9 13 3 10 9 7 13 15 1 10 0 9 2
14 0 1 15 13 13 2 16 4 1 15 13 10 9 2
2 15 2
5 13 11 7 11 2
7 13 11 2 15 13 11 2
5 7 11 13 11 2
24 12 9 15 7 9 13 2 16 11 13 3 7 3 2 13 10 9 7 13 15 15 1 9 2
11 13 3 9 9 2 15 13 9 2 9 2
4 7 11 13 2
3 1 9 2
8 16 4 15 13 13 2 13 2
8 1 0 9 2 1 0 9 2
9 15 15 13 2 7 10 9 11 2
15 3 14 13 0 9 2 7 16 11 3 13 2 13 9 2
15 1 9 7 1 9 12 9 15 13 1 9 1 9 11 2
42 7 3 2 1 0 9 2 15 1 11 13 3 16 15 12 9 9 2 15 15 1 9 13 2 13 9 1 9 9 7 9 1 9 7 13 15 1 9 1 9 9 2
8 3 13 9 7 13 0 9 2
11 15 13 1 9 2 9 2 9 2 9 2
9 0 7 9 15 3 13 1 9 2
7 1 9 13 0 9 9 2
9 12 7 15 9 13 9 7 9 2
48 9 15 13 9 0 2 13 1 9 1 0 9 7 9 2 13 11 0 9 2 16 15 13 7 3 13 2 7 1 9 0 9 11 13 2 16 15 2 15 15 13 15 2 15 13 7 0 2
15 16 10 9 3 13 2 10 9 15 4 13 7 1 9 2
5 3 4 13 9 2
7 0 9 15 3 13 9 2
26 4 2 14 13 13 9 2 16 4 13 9 2 4 13 13 7 10 9 1 9 7 10 9 1 15 2
13 16 11 13 2 15 9 13 10 9 2 10 9 2
20 0 9 4 13 9 0 9 2 15 2 15 13 0 2 4 13 3 7 0 2
16 3 13 0 7 0 9 2 13 4 2 13 7 13 9 3 2
5 13 15 7 9 2
8 9 13 13 2 9 15 13 2
19 9 9 2 15 13 13 9 9 2 7 13 9 11 2 4 13 2 13 2
6 13 15 15 7 9 2
3 3 3 2
12 1 9 0 9 15 13 2 16 13 3 0 2
5 7 3 3 13 2
12 13 1 9 2 16 9 13 13 0 15 9 2
12 3 4 7 13 0 2 7 0 2 9 9 2
21 3 15 11 10 9 13 2 3 15 2 15 15 13 13 9 1 9 11 7 11 2
10 1 9 13 7 13 9 7 9 9 2
13 13 3 2 16 10 9 13 7 13 0 9 0 2
10 13 3 2 16 13 3 13 16 13 2
28 13 2 15 2 15 13 15 2 2 16 1 0 9 13 9 0 13 10 0 9 1 15 0 1 15 2 13 2
12 7 15 3 13 13 10 0 9 0 0 9 2
11 0 0 9 1 9 2 15 15 13 13 2
9 7 9 9 13 15 2 15 13 2
16 9 0 1 10 0 9 1 15 13 12 1 0 9 10 9 2
16 7 10 9 13 3 0 2 16 13 14 9 2 7 7 9 2
13 9 11 11 1 11 11 2 3 0 9 0 9 11
16 9 11 1 0 9 12 2 9 2 0 3 1 9 9 11 11
25 11 11 2 9 2 2 11 11 2 11 2 7 11 11 2 11 2 1 9 0 9 1 9 1 9
4 9 1 0 9
28 1 10 0 0 9 1 9 1 9 13 9 11 11 12 0 9 2 0 9 2 11 10 10 9 7 0 9 2
20 0 12 4 9 13 2 16 4 13 0 9 1 0 9 9 2 12 1 11 2
27 0 9 0 9 15 3 13 9 9 12 2 12 2 15 1 10 3 0 0 9 3 13 7 0 0 9 2
8 1 0 9 13 9 0 9 2
29 3 1 9 0 11 11 2 9 11 11 2 2 3 11 1 9 0 11 2 11 2 11 0 9 0 9 9 9 2
15 1 9 15 13 1 9 11 2 7 3 1 0 0 9 2
22 9 0 9 13 0 9 2 13 10 3 0 2 1 15 3 0 9 13 3 7 3 2
7 11 11 7 3 13 9 2
19 16 15 1 9 16 9 13 0 0 9 2 9 15 13 1 10 0 9 2
24 9 2 11 11 2 1 3 0 9 13 1 0 9 7 1 9 0 9 13 10 3 0 9 2
14 9 13 3 0 0 9 7 3 9 7 9 0 9 2
17 9 1 9 9 13 1 9 11 7 11 12 9 3 0 0 9 2
3 9 7 9
22 0 9 15 13 1 9 2 3 15 1 0 9 1 0 9 13 11 2 11 11 2 2
30 10 0 9 1 11 2 0 1 9 15 0 0 9 2 11 11 2 2 13 9 0 9 7 10 9 13 1 0 9 2
31 9 0 9 7 0 9 15 1 0 0 9 7 9 13 2 11 15 13 1 0 9 7 9 15 13 0 9 2 13 2 2
5 2 13 9 2 2
36 1 0 9 9 13 1 9 1 11 2 9 15 1 0 7 0 9 7 0 9 13 1 0 9 2 2 0 2 3 0 0 9 9 0 9 2
10 1 9 15 1 9 0 9 3 13 2
23 0 9 7 9 13 0 9 1 9 2 9 1 0 9 13 3 0 9 7 9 0 9 2
60 0 9 13 9 9 9 2 1 0 9 2 9 0 9 11 11 2 2 3 1 15 13 3 0 9 11 11 16 3 0 9 11 2 0 9 2 1 15 11 13 10 9 13 1 0 9 7 9 0 9 2 15 1 0 9 13 9 11 11 2
2 9 9
6 0 9 0 9 13 2
24 13 15 3 1 0 9 7 0 9 0 0 9 16 1 9 0 9 9 2 9 7 0 9 2
12 9 0 9 1 0 0 9 13 3 0 9 2
8 13 15 7 9 0 0 9 2
39 1 15 13 3 0 9 13 0 9 1 0 7 0 9 13 2 13 14 9 1 9 7 9 2 15 13 10 0 9 2 2 7 3 7 1 9 7 9 2
8 15 15 13 7 0 0 9 2
17 13 2 14 11 2 9 1 9 9 1 0 9 15 13 3 0 2
10 7 15 13 14 0 9 0 0 9 2
18 3 16 1 9 13 11 7 1 9 9 1 9 0 9 1 9 9 2
9 13 15 12 9 0 9 7 9 2
22 11 11 11 2 3 10 9 2 7 3 10 3 0 9 2 10 0 2 7 0 9 2
20 7 11 11 11 2 15 13 1 3 0 9 13 3 0 9 0 9 7 9 2
14 9 1 9 2 11 2 11 2 11 2 11 2 9 2
11 9 11 11 2 9 11 11 7 11 11 2
25 9 11 11 2 9 11 2 9 11 11 2 9 11 11 2 0 9 11 11 2 0 9 11 11 2
5 9 12 2 9 2
28 11 11 2 0 2 12 2 13 1 0 9 3 3 3 1 9 12 2 3 1 0 0 9 11 13 0 9 2
24 1 10 9 0 10 9 2 16 3 1 9 0 7 3 0 2 13 0 9 9 7 0 9 2
29 1 9 0 9 15 11 11 13 0 9 9 1 9 2 16 13 1 9 2 0 1 9 9 7 9 9 11 11 2
6 11 2 11 7 9 9
9 9 0 7 0 13 1 9 0 9
21 11 11 7 11 2 11 11 13 3 0 7 3 0 9 0 9 0 12 0 9 2
6 12 13 1 0 9 2
15 0 9 3 13 13 3 0 2 7 13 3 1 15 0 2
24 0 0 9 10 9 13 2 16 13 12 1 0 9 0 9 2 3 9 2 0 1 0 2 2
14 7 3 2 0 7 0 9 13 1 9 7 0 9 2
16 10 9 13 7 3 0 2 9 12 9 15 3 3 3 13 2
43 16 1 9 13 13 9 10 9 3 9 7 9 0 9 1 0 9 2 3 1 9 13 1 1 10 0 9 9 0 3 9 0 3 9 7 9 1 0 9 7 0 9 2
33 7 3 2 15 13 13 0 16 9 0 2 3 0 2 9 1 9 1 15 2 15 9 15 1 15 13 3 2 3 1 9 0 2
9 9 7 9 13 1 9 12 9 2
10 11 15 15 7 13 3 3 16 11 2
11 9 15 13 3 1 10 0 2 0 9 2
17 9 15 15 13 9 2 14 16 15 13 2 16 15 13 1 9 2
25 1 11 13 3 9 0 1 10 9 2 16 4 3 13 1 9 2 9 7 9 13 3 3 13 2
11 11 15 13 9 2 9 2 7 3 9 2
15 0 9 2 9 7 0 9 16 4 13 1 9 0 9 2
8 9 10 9 13 13 11 11 2
15 11 13 9 7 3 9 2 7 1 10 9 13 15 13 2
14 9 7 0 9 10 3 0 9 16 4 13 1 9 2
10 10 0 9 13 0 9 1 0 9 2
16 13 0 2 16 1 9 12 1 10 9 13 13 9 9 11 2
8 11 13 1 9 9 3 0 2
20 9 10 9 2 3 16 1 11 2 13 9 2 7 13 3 9 16 9 9 2
10 3 1 10 9 3 13 9 7 9 2
8 12 10 9 13 0 9 11 2
22 13 3 3 0 2 7 3 0 2 13 0 9 3 2 3 13 15 3 1 11 11 2
19 9 1 0 9 7 9 1 9 9 2 0 9 1 9 7 9 2 2 2
13 3 3 15 13 2 7 3 13 1 9 3 0 2
18 9 4 13 2 11 9 2 2 10 9 13 9 7 0 9 10 9 2
12 0 9 13 10 9 7 15 3 7 0 9 2
11 10 9 13 13 1 10 9 1 11 11 2
27 16 4 15 15 13 13 7 3 2 13 11 3 1 9 7 9 9 13 13 2 15 13 13 9 0 9 2
15 4 3 13 1 11 7 10 9 3 13 9 1 0 9 2
9 0 0 9 15 13 7 13 3 2
19 9 1 11 13 2 16 0 9 2 0 2 7 2 0 2 13 15 0 2
16 9 2 1 15 15 13 2 13 7 0 7 13 13 1 9 2
11 13 0 13 15 2 15 4 10 9 13 2
26 1 0 9 9 2 15 13 13 9 10 9 2 13 0 3 13 2 3 15 10 9 13 3 3 0 2
26 13 4 0 13 2 16 9 0 12 9 13 0 2 16 10 9 13 9 9 2 0 9 13 1 15 2
28 13 15 13 2 16 13 1 0 9 2 0 9 4 15 7 13 13 3 7 1 3 3 3 0 9 11 11 2
13 16 4 13 9 2 13 4 13 2 16 0 13 2
20 16 4 13 9 9 2 13 16 13 15 0 9 2 14 3 0 0 9 3 2
12 9 7 9 13 13 16 9 0 9 7 9 2
25 3 0 9 2 16 0 7 0 2 9 7 9 2 13 3 13 16 9 2 16 4 0 9 13 2
9 3 2 16 10 9 13 0 9 2
9 9 13 7 3 13 9 10 9 2
27 13 15 2 16 4 0 9 0 9 13 1 15 0 2 0 2 7 3 3 13 0 15 13 1 0 9 2
16 0 9 13 3 0 9 2 3 13 9 7 9 9 9 9 2
9 0 9 13 9 7 3 15 13 2
25 9 13 3 9 9 13 7 3 15 13 2 3 0 2 9 2 10 9 13 13 7 1 9 0 2
38 0 9 14 13 2 16 13 2 14 15 2 15 9 1 15 13 16 9 2 13 3 3 2 13 15 0 9 2 9 7 9 2 15 13 13 3 0 2
4 3 9 13 3
45 3 9 13 3 14 9 9 2 13 3 1 9 2 15 13 2 7 15 13 9 2 13 0 9 2 7 13 9 0 1 10 9 2 1 9 0 9 2 0 1 10 9 7 9 2
25 7 3 2 9 2 13 13 10 9 2 16 4 0 13 10 9 2 13 7 13 2 3 13 0 2
5 6 0 9 9 2
13 15 15 13 13 2 7 15 13 15 12 1 0 2
51 7 0 9 2 3 9 0 2 9 7 9 0 2 13 9 2 1 9 15 13 2 1 10 9 15 13 2 16 4 13 0 9 2 16 4 1 9 9 13 9 15 2 15 3 1 9 13 9 0 9 2
12 1 9 9 9 2 13 11 11 2 0 9 12
2 9 9
34 16 15 11 11 13 9 10 9 9 2 15 3 13 1 0 9 2 7 15 1 15 3 13 2 13 15 15 14 9 2 7 7 9 2
68 7 14 3 1 10 9 2 1 0 4 15 3 13 2 16 1 15 1 10 0 9 4 13 2 1 0 4 15 13 9 1 9 14 0 9 9 2 15 15 13 9 1 9 2 1 0 1 15 13 0 9 2 1 15 4 15 1 15 0 2 16 3 0 2 13 16 9 2
28 7 1 0 4 15 13 13 9 1 10 9 9 3 2 3 9 11 11 9 11 11 13 0 9 1 9 9 2
17 9 1 9 15 15 13 2 16 15 15 9 7 9 13 1 9 2
20 16 15 13 2 16 4 15 13 1 9 2 16 3 13 2 13 15 10 9 2
34 7 7 15 15 13 3 3 7 0 13 2 16 15 10 13 2 16 4 15 16 12 1 9 9 7 9 1 9 13 14 3 1 9 2
26 7 3 13 2 16 16 13 15 9 2 3 3 0 9 2 1 15 3 15 13 3 12 9 3 0 2
20 1 10 9 13 10 0 9 7 9 9 9 9 7 9 1 0 9 11 11 2
30 13 15 15 12 2 13 4 0 9 7 9 7 9 1 15 2 15 15 1 15 7 1 15 2 13 2 1 0 9 2
16 0 9 15 13 2 0 9 0 2 16 4 15 13 1 9 2
42 14 4 15 1 0 0 9 13 1 9 2 15 13 13 3 16 15 2 13 3 3 16 15 2 7 3 1 15 13 9 2 9 7 9 2 15 15 3 2 13 2 2
34 14 15 15 3 13 2 16 13 9 15 2 15 15 3 3 13 11 11 7 11 11 2 16 0 9 9 7 9 1 9 13 10 9 2
16 15 15 15 13 2 3 7 1 9 9 13 3 9 0 9 2
22 15 1 15 13 2 16 13 9 1 9 2 3 13 13 9 2 7 9 2 2 9 2
11 3 1 10 9 1 9 0 9 3 13 2
42 1 9 0 9 3 13 2 16 11 13 0 9 3 9 1 0 9 1 9 7 14 3 9 2 7 0 16 9 1 9 0 9 7 9 13 15 9 1 9 7 9 2
8 7 3 13 15 1 9 9 2
10 3 1 9 4 13 7 0 1 9 2
13 3 4 7 13 2 16 1 10 9 1 9 13 2
7 16 13 15 3 0 9 2
3 7 9 2
19 16 13 0 9 13 9 1 9 2 7 14 1 9 15 2 7 0 9 2
17 13 0 7 0 2 16 4 7 15 3 13 1 15 2 16 13 2
17 7 16 15 10 9 13 9 2 16 4 11 11 13 14 1 15 2
3 9 0 9
8 11 11 15 13 1 9 12 2
10 13 9 7 9 1 0 9 1 11 2
16 1 9 15 13 0 9 7 11 11 2 0 9 7 0 9 2
19 13 9 0 9 0 9 2 3 15 3 13 10 9 2 9 11 11 2 2
13 0 7 0 13 10 9 0 0 9 2 3 9 2
6 13 15 3 7 9 2
8 10 0 9 13 0 9 9 2
8 11 13 1 9 12 1 9 2
14 11 2 11 11 15 13 1 9 9 12 1 0 11 2
10 13 9 1 0 11 7 1 0 9 2
18 13 1 0 0 9 7 3 1 11 2 1 11 2 11 7 11 2 2
18 3 1 0 11 15 13 1 0 2 7 7 0 9 0 9 0 9 2
16 11 13 9 1 11 11 11 2 15 1 10 9 13 0 9 2
7 0 0 9 13 16 0 2
24 10 0 0 9 1 10 9 13 9 0 9 2 15 15 13 1 9 0 9 2 9 7 9 2
3 1 0 9
11 11 2 11 2 11 2 9 13 9 12 2
18 0 9 9 0 9 2 9 7 9 13 0 9 0 9 1 9 0 2
8 13 0 11 1 9 11 11 2
6 11 11 2 9 11 2
20 0 9 0 9 0 9 1 11 11 1 11 11 13 1 9 0 9 7 9 2
11 13 0 9 2 13 11 11 7 11 11 2
6 11 11 2 0 9 2
24 0 9 1 9 9 1 9 9 0 0 9 2 9 11 11 2 13 13 1 11 9 0 9 2
18 0 9 11 11 2 0 0 9 4 13 9 12 2 13 11 2 9 2
8 11 11 2 0 9 7 9 2
23 0 9 7 9 0 2 0 9 13 1 9 1 0 9 0 11 2 15 13 9 11 11 2
5 2 0 2 9 13
55 0 9 1 10 9 2 0 9 0 9 0 13 2 13 15 3 2 4 13 3 1 11 9 13 1 9 11 2 13 9 2 0 9 2 9 0 9 1 11 1 9 2 13 11 11 9 2 3 1 9 3 16 9 15 2
14 15 13 7 1 9 13 3 1 9 10 9 2 2 2
38 0 9 9 9 14 0 0 0 9 2 0 15 1 11 3 0 0 7 0 9 2 13 1 11 9 1 0 7 0 0 9 1 9 0 7 0 9 2
55 1 9 0 0 9 13 9 0 7 0 2 1 15 13 0 0 9 2 1 0 9 2 15 15 16 9 13 1 0 9 7 1 15 15 1 9 1 9 2 9 11 11 13 3 13 2 13 9 1 15 0 9 2 9 2
26 9 3 7 3 13 3 16 4 13 0 9 9 0 11 2 2 13 13 1 15 2 15 4 13 2 2
4 0 0 9 2
6 9 9 7 3 0 9
14 13 15 1 9 0 1 9 12 2 3 7 3 0 2
33 13 13 2 16 13 0 9 2 15 15 13 0 9 0 9 7 1 9 0 9 1 9 0 9 7 0 9 9 1 0 9 11 2
23 0 0 9 0 0 9 10 9 1 12 9 2 15 13 9 11 11 2 3 13 9 9 2
8 1 12 9 13 1 9 0 2
18 13 15 2 16 0 9 13 13 10 0 9 1 10 9 2 3 9 2
23 9 11 9 1 0 9 13 9 0 0 9 2 11 11 1 11 2 1 12 2 12 2 2
25 13 10 9 2 1 9 0 9 11 12 2 15 13 9 2 13 13 9 2 0 9 7 12 9 2
22 0 9 2 15 15 13 2 15 13 1 9 9 11 9 7 1 9 13 13 0 9 2
13 10 9 13 1 0 9 9 9 11 7 9 9 2
20 0 9 2 9 1 9 7 1 9 2 7 11 7 15 13 9 7 13 9 2
35 7 1 9 1 11 2 3 16 1 0 9 1 9 2 1 9 2 1 9 13 9 2 7 0 9 15 1 9 9 13 1 9 1 9 2
21 1 9 1 0 0 9 1 11 2 0 1 9 12 2 13 7 0 9 3 0 2
40 13 3 10 0 2 3 0 2 9 7 3 10 9 1 9 7 11 2 11 1 15 13 1 9 14 3 2 16 13 13 15 7 10 9 7 13 13 0 9 2
41 0 9 11 11 11 13 2 16 9 11 13 9 0 9 2 15 15 1 10 9 16 0 9 13 1 9 2 0 15 1 9 1 9 2 3 13 0 9 1 15 2
4 9 1 11 2
7 13 9 11 2 11 12 2
7 13 7 9 13 11 11 2
8 12 9 2 9 7 9 13 2
3 9 7 9
32 1 9 9 11 11 13 1 0 9 9 9 1 9 2 12 2 2 1 15 9 9 7 9 11 11 13 10 0 9 0 9 2
31 9 9 2 15 13 13 1 3 0 7 3 0 9 0 0 9 11 2 9 13 1 11 9 0 9 2 0 9 0 9 2
23 9 9 13 0 9 11 11 2 15 15 13 1 9 9 1 9 1 0 9 2 2 2 2
28 0 9 9 1 9 3 13 11 11 2 9 3 0 0 9 13 0 0 0 9 1 9 9 0 9 11 11 2
22 3 0 9 2 15 13 0 9 2 9 11 11 3 2 3 3 2 13 1 0 9 2
24 11 11 15 1 9 9 3 13 7 9 13 0 9 1 9 7 9 10 9 2 15 13 3 2
15 11 11 2 3 2 7 11 11 1 9 1 9 9 1 9
19 9 7 9 11 11 2 12 2 15 0 9 13 1 9 1 9 0 9 2
59 1 10 0 9 0 9 2 12 2 13 10 0 9 2 3 0 0 9 2 0 9 9 2 12 2 1 9 11 11 2 0 9 1 0 9 9 2 12 2 2 9 1 12 9 9 1 9 2 12 2 7 9 9 9 1 9 0 9 2
2 0 9
22 10 9 13 1 0 9 16 9 1 9 2 15 15 3 13 9 11 11 1 0 11 2
21 13 15 3 0 9 2 9 15 1 15 13 1 10 9 7 3 1 9 1 9 2
43 1 0 15 13 1 9 1 15 2 16 13 9 0 15 0 9 1 9 7 16 13 10 9 2 15 13 0 9 10 9 7 15 3 13 13 2 16 1 15 13 0 9 2
14 16 9 9 0 9 1 0 13 11 2 11 9 9 2
19 13 4 15 3 1 9 2 16 0 9 7 0 9 10 9 13 0 9 2
16 0 9 2 15 4 13 1 0 2 13 15 7 9 9 13 2
13 14 1 9 4 13 9 1 11 2 11 1 11 2
21 9 15 1 15 13 2 16 4 13 9 9 2 15 15 13 1 9 2 9 2 2
9 14 2 13 3 1 10 0 9 2
8 10 9 13 12 3 0 9 2
42 13 7 2 9 1 9 9 2 9 3 2 2 2 7 3 2 9 1 9 1 9 0 9 2 2 7 2 9 3 15 0 9 1 0 9 2 7 3 2 9 2 2
14 13 0 2 16 15 3 13 0 9 0 1 0 9 2
6 13 3 1 0 9 2
11 0 9 13 14 9 1 9 2 9 3 2
18 1 0 0 9 15 13 0 9 9 2 7 13 13 14 9 0 9 2
38 9 11 2 11 13 1 0 9 2 9 2 0 9 2 7 1 15 13 9 9 0 2 1 0 3 9 2 0 2 0 9 2 2 13 2 9 2 2
13 1 0 9 13 7 0 9 2 9 2 9 2 2
19 3 15 3 13 1 9 9 2 7 11 2 11 13 1 0 9 9 9 2
22 9 13 9 1 10 2 16 0 9 9 4 13 1 0 9 2 7 13 1 0 9 2
12 1 12 2 9 2 15 3 13 9 1 9 2
21 13 4 13 1 9 2 15 13 1 9 7 9 9 2 13 2 0 9 13 2 2
15 16 13 15 3 2 9 9 7 9 3 1 10 9 13 2
19 1 0 9 2 9 3 15 0 9 2 4 9 13 1 9 2 9 2 2
14 13 15 9 1 0 0 9 13 1 9 2 13 2 2
23 13 13 2 16 9 13 1 9 3 2 9 2 7 3 13 0 9 9 2 0 9 2 2
16 3 16 1 0 9 13 9 9 13 7 1 9 1 0 9 2
9 9 1 10 9 13 1 15 9 2
20 3 0 0 9 13 9 9 2 15 13 1 9 3 1 0 9 2 13 2 2
10 13 9 9 0 1 0 9 7 9 2
13 1 0 9 2 9 2 13 9 9 1 0 9 2
22 13 0 0 9 7 13 15 3 1 0 9 9 2 3 2 13 4 1 9 9 2 2
18 4 13 1 9 2 0 11 2 7 1 9 13 1 0 9 0 9 2
19 13 15 3 14 1 9 0 9 13 9 2 1 15 13 9 1 0 9 2
25 0 9 0 9 15 3 3 13 2 16 15 9 13 13 9 13 9 2 15 13 0 9 9 13 2
11 3 3 15 1 0 0 9 13 13 9 2
18 16 9 13 9 4 13 1 0 9 2 9 1 9 9 13 1 0 2
26 1 9 9 13 2 3 15 10 9 13 10 0 9 1 0 9 7 3 15 13 1 9 0 0 9 2
7 9 0 9 2 12 2 2
15 9 1 0 9 4 3 13 7 13 15 9 9 0 9 2
21 13 14 15 2 1 15 13 9 12 9 1 0 9 7 15 13 1 0 9 0 2
11 12 9 1 9 1 9 13 9 1 9 2
28 13 15 3 3 2 16 13 9 13 1 9 2 7 16 9 3 1 9 13 13 9 9 7 9 1 9 9 2
57 1 0 9 1 9 12 13 3 1 0 9 2 0 2 9 12 9 12 9 12 9 12 9 12 9 12 2 0 2 9 12 9 12 9 12 9 12 2 0 9 1 0 9 2 7 10 9 13 0 9 7 10 9 9 3 13 2
8 0 13 1 9 7 13 12 2
12 7 1 12 9 13 0 13 7 0 13 9 2
51 9 11 2 11 1 9 12 2 0 2 9 12 9 12 9 12 9 12 9 12 9 12 2 0 2 9 12 9 12 9 12 9 12 9 12 2 2 1 15 13 0 1 9 2 13 1 9 3 2 12 2
3 7 13 2
9 1 0 9 15 10 9 13 3 2
13 9 13 9 1 9 11 2 11 11 2 11 12 2
5 0 9 13 12 2
9 0 9 0 13 3 9 0 9 2
21 0 9 7 9 15 3 3 13 2 9 13 9 1 0 9 14 1 0 9 2 2
15 1 9 11 2 11 2 11 12 2 1 9 1 9 12 2
9 2 0 9 2 0 13 9 2 2
14 0 9 2 0 9 9 12 13 7 9 12 15 13 2
4 0 15 13 2
40 9 1 9 15 13 2 11 2 11 1 11 2 9 2 11 2 11 1 0 11 2 9 2 11 2 11 1 11 11 2 11 2 11 7 11 2 11 1 11 2
2 13 2
2 13 9
9 0 9 9 12 13 0 0 9 2
16 1 9 9 4 13 1 9 7 13 15 9 0 11 2 11 2
9 1 9 13 12 2 9 10 9 2
38 9 1 9 2 0 2 9 12 9 12 9 12 9 12 9 12 9 12 2 0 2 9 12 9 12 9 12 9 12 2 13 9 2 0 1 9 13 2
7 0 13 9 1 0 9 2
16 9 15 0 9 13 1 9 9 0 9 1 12 2 9 12 2
5 9 16 9 1 9
8 2 9 12 2 12 2 12 2
25 0 9 13 1 9 1 9 9 1 0 9 7 1 15 0 7 13 10 0 2 9 1 9 2 2
13 9 9 0 1 0 9 9 13 1 9 9 9 2
30 1 0 9 9 1 10 9 13 13 0 2 13 13 10 9 9 2 1 15 3 13 10 9 0 2 0 2 0 3 2
20 1 10 9 7 1 0 9 15 3 13 7 9 10 9 2 16 13 13 0 2
30 3 7 13 9 11 1 9 1 9 10 0 9 2 0 1 0 9 9 2 7 9 9 2 15 13 3 9 0 9 2
54 1 0 9 13 13 1 11 11 1 15 2 16 4 0 9 2 0 1 0 0 9 2 15 13 9 13 9 9 2 16 3 13 1 0 0 9 2 9 0 9 2 0 9 7 15 0 2 13 9 9 1 0 9 2
23 3 13 9 0 12 9 2 13 15 3 9 0 9 2 15 15 13 0 9 9 0 9 2
5 2 2 2 2 2
46 13 2 14 3 15 1 15 1 0 9 2 13 15 3 9 2 15 13 15 1 15 2 9 9 2 15 15 13 13 12 1 0 2 13 15 9 7 9 3 2 3 15 3 9 13 2
32 9 2 1 15 15 13 9 11 2 13 3 0 7 13 9 0 9 2 3 9 13 1 9 1 9 2 15 1 15 9 13 2
48 1 0 9 13 9 15 13 1 15 2 15 13 13 1 9 0 2 7 2 15 2 1 15 13 9 9 9 2 9 7 9 0 9 2 15 9 13 1 9 2 7 3 3 13 10 0 9 2
13 13 0 2 16 3 14 15 0 15 13 3 13 2
52 13 2 14 7 3 3 9 1 9 9 9 2 3 2 1 9 9 9 1 9 0 7 0 2 13 3 3 3 1 0 9 9 0 12 9 2 3 15 1 0 9 9 13 0 0 9 1 9 0 0 9 2
14 3 3 3 13 0 9 2 10 0 0 9 13 9 2
36 9 10 9 1 9 0 13 3 0 9 1 0 9 2 7 3 7 3 0 9 9 2 0 9 1 0 9 7 2 15 13 15 2 1 9 2
50 13 2 14 3 13 9 1 0 9 10 9 2 9 2 15 4 13 7 3 13 0 9 2 13 13 9 2 3 4 13 9 13 2 15 13 1 10 9 0 2 0 2 7 15 13 0 2 0 2 2
6 9 1 9 13 9 2
7 12 9 0 2 12 9 9
8 2 9 12 2 12 2 12 2
7 9 10 9 13 3 0 2
47 1 9 15 1 0 9 7 9 13 9 2 15 13 2 16 7 13 1 9 0 2 7 3 3 13 2 7 1 0 13 0 7 0 9 7 9 2 15 15 3 13 15 2 15 0 13 2
26 15 7 13 2 3 1 0 9 9 7 9 13 9 2 3 13 9 9 7 9 7 13 15 1 9 2
41 15 13 3 0 2 16 7 0 9 0 14 0 9 1 9 7 0 9 1 9 13 15 0 9 9 13 13 2 16 3 13 2 16 9 2 9 3 2 3 13 2
21 7 13 3 0 13 9 7 13 3 0 2 16 4 1 15 13 2 0 0 9 2
4 0 9 0 9
8 2 9 12 2 12 2 12 2
12 1 9 4 15 13 9 11 11 1 11 11 2
7 13 1 9 9 1 11 2
15 13 0 2 16 15 3 13 1 15 2 3 15 3 13 2
11 3 15 4 15 1 11 11 1 9 13 2
8 1 11 4 13 9 9 12 2
7 13 15 3 12 12 9 2
14 1 10 0 9 13 0 9 2 1 15 15 13 9 2
22 15 0 4 13 0 2 14 16 13 1 9 2 7 3 3 3 2 16 13 1 9 2
13 7 3 15 3 13 9 0 2 15 13 1 9 2
28 3 7 3 1 9 4 13 9 2 1 15 4 13 0 9 2 16 4 15 13 1 9 2 1 15 13 9 2
12 7 3 4 3 13 13 15 3 1 0 9 2
13 15 0 4 13 13 16 3 3 0 9 11 11 2
23 4 4 13 13 15 3 1 10 9 2 15 15 3 13 1 10 0 9 1 9 0 9 2
13 1 10 9 15 13 1 12 7 3 9 7 9 2
7 11 11 13 3 0 9 2
11 16 13 7 3 0 7 13 3 3 13 2
16 3 3 13 13 9 2 7 13 15 3 0 9 1 0 9 2
6 10 9 4 13 0 2
18 0 9 1 15 13 2 16 3 0 7 0 9 13 9 0 7 0 2
13 3 4 13 1 15 2 16 15 3 3 13 13 2
10 0 9 13 0 9 7 0 9 0 2
8 1 9 15 15 13 3 13 2
33 1 9 12 4 13 1 9 1 11 2 7 7 1 15 13 9 2 3 4 13 13 9 9 2 15 3 10 9 7 9 15 13 2
9 13 4 9 2 16 4 15 13 2
16 1 9 4 15 13 2 16 11 11 13 1 15 3 1 11 2
5 14 13 10 9 2
25 3 2 16 1 9 13 0 10 0 9 13 15 12 2 13 15 3 1 10 0 9 1 0 9 2
5 0 9 9 7 9
8 2 11 12 2 12 2 12 2
10 3 0 13 0 9 1 9 7 9 2
31 15 0 1 11 12 2 12 2 13 1 15 3 0 2 16 3 2 16 3 15 13 10 9 1 9 1 9 0 9 0 2
15 1 9 4 3 13 2 3 13 13 0 9 9 0 9 2
76 13 2 3 13 0 9 9 9 11 2 11 2 15 4 9 13 7 1 9 10 9 15 13 1 0 9 2 7 16 13 3 0 7 15 2 13 2 13 10 9 2 2 2 2 2 2 13 15 1 15 7 12 0 9 2 7 6 2 15 15 3 13 1 10 9 2 15 2 1 10 9 2 13 3 0 2
23 10 9 13 9 7 1 9 2 1 15 4 13 2 13 9 13 1 9 1 9 9 9 2
10 0 9 1 12 9 13 3 1 9 2
39 13 15 3 3 1 9 2 7 16 15 13 10 0 9 2 3 15 9 13 3 13 2 13 3 2 13 1 9 10 0 9 9 2 15 9 11 3 13 2
46 2 2 2 2 2 7 14 1 9 2 16 13 1 9 2 1 9 15 2 10 9 1 0 9 9 3 2 2 2 1 9 9 0 9 0 2 13 3 2 2 2 2 2 9 9 2
39 0 9 15 7 13 1 0 7 7 1 0 9 2 3 9 2 2 13 9 1 9 9 2 13 6 1 9 2 2 2 2 2 15 13 13 14 1 9 2
5 2 2 2 2 2
10 7 13 3 0 0 9 2 13 9 2
26 0 9 9 13 3 3 0 2 3 3 16 1 15 0 0 9 9 2 0 0 9 2 9 2 9 2
18 1 10 0 9 15 13 1 9 9 2 15 13 9 1 9 9 3 2
31 12 9 2 15 13 9 0 0 9 1 9 1 0 9 1 9 2 15 3 13 1 11 7 13 1 9 14 1 0 9 2
27 10 3 0 0 9 7 1 10 0 9 13 2 16 1 10 9 13 0 9 1 9 9 0 9 1 9 2
24 3 3 2 16 15 13 1 9 1 9 2 7 7 15 15 13 1 10 9 7 13 15 9 2
8 3 15 13 0 9 1 11 2
35 10 0 9 2 9 0 0 0 2 3 7 0 7 1 0 9 0 9 2 15 13 1 11 9 9 7 10 9 15 13 1 0 0 9 2
35 1 9 9 9 0 9 1 0 9 13 13 0 7 9 9 11 13 1 9 9 3 3 16 10 9 0 3 1 0 0 9 1 0 9 2
10 0 9 13 9 7 13 15 9 0 2
18 15 3 13 2 15 15 13 2 0 11 2 7 2 0 9 11 2 2
20 14 13 9 9 2 7 14 9 2 7 2 16 13 13 2 7 3 0 9 2
5 9 13 9 1 9
8 2 11 12 2 12 2 12 2
10 13 3 0 2 16 9 4 3 13 2
7 13 2 16 3 13 9 2
29 13 2 14 15 2 15 13 1 0 9 3 2 9 2 16 4 15 13 9 2 3 3 13 0 9 15 15 13 2
10 13 3 9 9 2 7 3 14 0 2
37 16 4 13 1 9 12 1 9 16 0 9 7 13 0 9 2 13 10 9 3 14 12 9 7 1 15 4 13 0 0 12 9 1 2 9 2 2
20 3 3 13 0 1 0 9 2 0 9 2 2 7 2 16 9 13 1 9 2
34 3 13 1 0 9 9 9 2 7 0 3 3 13 9 0 9 9 7 1 15 15 9 13 0 9 2 3 2 9 13 12 9 2 2
12 1 10 9 13 9 12 5 7 9 12 5 2
40 3 15 13 0 9 1 9 1 9 2 9 7 9 2 7 16 0 9 0 9 13 9 0 9 9 2 1 15 15 13 2 7 15 13 1 10 9 0 9 2
3 14 9 13
12 1 0 9 13 2 3 9 2 1 11 9 2
19 1 0 9 15 15 13 2 9 1 0 9 3 13 1 0 9 0 9 2
8 9 7 9 9 13 0 9 2
5 7 3 14 0 2
14 13 2 16 11 13 1 0 9 2 1 0 0 9 2
28 13 14 9 2 16 15 15 2 15 15 13 1 9 7 9 9 2 13 2 16 10 9 13 13 15 9 3 2
10 0 9 13 1 10 9 9 3 0 2
20 3 9 9 0 0 0 9 13 3 1 9 12 1 0 0 9 2 9 9 2
12 1 0 9 3 2 13 2 15 15 0 13 2
9 9 9 13 11 16 9 1 9 2
40 15 15 15 13 2 13 15 2 16 15 1 9 9 7 12 9 13 0 9 2 3 0 1 0 9 2 1 0 9 7 1 0 9 7 0 9 1 0 9 2
30 15 15 15 13 2 13 15 1 9 1 9 9 3 7 3 0 1 9 1 0 9 2 10 9 13 0 9 0 9 2
30 0 9 13 0 9 3 3 0 9 1 12 0 9 2 11 7 0 9 7 9 1 0 9 1 0 9 1 0 11 2
18 9 2 0 9 2 7 3 13 1 9 0 9 11 11 9 0 9 2
59 1 1 0 9 9 2 3 0 9 2 0 9 7 9 1 9 2 13 9 1 9 3 0 1 0 0 9 2 9 1 0 9 1 9 1 9 7 9 11 1 0 0 9 0 0 9 2 7 13 1 9 9 12 9 1 9 7 9 2
10 1 0 0 9 1 0 11 13 9 2
11 9 2 1 0 9 1 9 7 15 9 2
17 13 3 9 9 2 16 13 11 13 1 0 7 1 3 0 9 2
14 0 9 13 10 0 9 2 7 7 3 13 9 9 2
12 2 0 9 13 9 2 1 9 13 12 9 2
26 7 7 15 3 13 9 2 2 13 11 11 2 15 3 13 11 1 9 0 3 1 9 16 1 9 2
66 1 9 13 7 9 0 1 9 2 15 3 13 10 9 16 3 9 1 0 11 2 1 11 2 2 15 0 15 1 9 14 13 1 9 2 3 16 3 0 0 9 2 15 4 3 13 1 10 9 2 2 7 1 0 9 15 13 9 0 9 0 2 0 9 2 2
41 0 2 3 0 9 2 15 13 1 0 9 7 1 0 9 10 9 2 2 3 2 3 14 3 0 9 0 1 9 2 2 13 1 0 9 14 0 9 10 9 2
10 2 15 3 3 13 2 13 15 13 2
28 1 9 7 3 3 1 0 9 2 2 13 3 0 9 9 2 15 13 13 7 3 13 1 0 9 0 9 2
36 0 9 7 0 9 2 9 15 3 16 1 11 0 11 13 11 2 13 7 9 2 16 1 2 9 2 13 1 9 9 13 9 9 1 15 2
19 9 13 0 13 1 11 7 1 0 9 2 1 9 13 13 14 0 9 2
41 2 16 15 1 9 12 9 13 7 13 9 2 13 4 0 9 15 1 9 2 2 13 15 9 11 2 15 4 1 0 9 1 9 3 15 0 9 13 14 9 2
7 13 7 2 16 15 13 2
22 1 0 9 3 15 0 9 7 9 3 1 9 3 3 13 13 14 1 0 9 9 2
6 9 9 13 9 10 9
25 3 15 3 0 9 9 13 10 9 1 9 2 16 9 13 1 9 7 9 3 3 1 0 9 2
38 9 2 3 16 9 2 9 7 0 9 0 15 9 2 13 14 3 9 1 0 9 2 2 3 13 9 9 9 2 16 9 1 9 10 9 2 2 2
13 9 1 9 13 0 2 13 9 0 7 13 9 2
10 1 9 10 9 3 13 3 7 3 2
19 13 13 1 0 0 9 2 15 13 14 0 9 1 0 9 1 10 9 2
16 9 7 9 1 15 13 15 2 13 7 13 7 3 14 15 2
6 0 0 9 13 0 2
12 3 7 15 13 10 0 9 2 3 10 9 2
13 9 13 2 16 10 3 0 0 9 13 11 11 2
2 0 9
13 0 9 0 9 16 4 15 1 0 9 13 3 2
9 0 9 9 13 3 13 12 9 2
31 9 0 1 15 13 2 16 0 9 2 1 0 3 13 9 2 3 10 9 13 2 7 10 9 15 13 1 9 0 9 2
21 9 0 0 9 3 13 1 9 15 0 9 9 2 7 9 13 13 2 15 13 2
11 9 2 3 3 15 13 2 13 3 0 2
10 9 9 13 1 9 3 9 0 9 2
10 15 3 13 1 9 1 9 10 9 2
36 13 0 9 2 13 4 1 9 0 0 9 2 13 4 15 13 9 7 9 2 13 4 15 13 0 0 7 0 9 2 0 1 9 0 9 2
15 3 4 7 13 0 9 2 0 9 7 0 9 0 9 2
4 3 9 2 9
14 9 9 0 9 13 3 13 1 9 1 9 0 9 2
21 13 1 15 2 16 4 9 13 0 2 7 1 15 2 16 13 1 9 3 13 2
44 9 9 7 9 2 3 9 2 3 7 0 9 2 3 13 10 9 0 9 7 9 2 10 9 7 13 9 2 7 15 9 2 15 4 9 13 7 15 3 4 3 7 13 2
18 9 15 4 3 13 2 13 7 3 0 9 7 13 7 1 10 9 2
22 1 10 0 9 13 3 7 0 9 1 11 7 0 9 3 3 13 10 9 13 9 2
22 0 9 13 3 1 0 9 1 9 0 9 2 15 3 3 13 1 9 1 0 9 2
32 1 0 9 13 7 3 0 9 2 15 13 3 0 9 0 9 1 12 2 2 12 2 9 2 1 15 13 13 0 9 0 2
35 1 15 15 9 9 13 3 3 2 13 13 2 16 3 0 0 9 7 9 0 9 11 13 1 0 9 1 9 11 7 13 7 9 11 2
3 9 1 9
27 1 10 0 9 10 9 13 0 9 11 11 2 15 13 0 9 1 9 1 9 0 9 1 9 0 9 2
25 15 0 0 9 13 0 9 2 1 15 13 13 9 3 1 0 9 2 15 13 3 3 9 2 2
25 1 12 2 9 15 9 2 3 16 9 2 13 0 9 9 1 10 9 1 0 9 0 0 9 2
22 0 9 7 13 9 2 12 1 11 12 2 11 0 9 2 1 0 7 1 0 9 2
12 0 9 3 3 13 9 9 2 7 0 9 2
20 13 3 1 0 9 13 1 9 2 13 15 7 3 9 13 0 1 0 9 2
2 0 9
23 0 9 15 1 9 0 9 3 13 0 0 9 2 1 15 13 0 9 9 9 2 9 2
24 3 15 3 3 13 9 0 2 1 9 2 7 2 1 9 0 2 1 0 2 1 9 2 2
20 1 9 7 0 9 13 9 1 10 9 3 0 0 9 2 15 3 13 0 9
6 2 14 2 0 9 9
16 9 2 0 7 0 9 2 15 1 9 13 1 9 7 13 2
15 0 15 2 15 13 10 9 3 13 2 7 3 3 13 2
14 7 16 3 13 9 9 11 2 9 9 15 3 13 2
12 0 9 2 9 9 7 0 9 15 14 13 2
16 9 9 1 9 1 15 13 0 9 0 1 9 9 7 9 2
14 0 7 0 9 0 9 2 15 4 3 13 9 11 2
15 13 2 13 15 3 0 7 0 0 9 13 15 14 9 2
30 0 0 9 15 3 13 15 2 15 13 0 1 9 9 2 13 0 9 7 1 10 9 13 9 1 9 0 0 9 2
19 11 11 13 13 1 9 1 9 2 0 9 2 0 9 7 3 1 9 2
22 15 13 7 9 2 11 0 11 7 11 11 2 16 3 13 9 1 0 9 1 9 2
33 7 11 11 13 9 2 16 13 0 9 1 0 9 7 3 16 0 9 2 7 0 9 1 9 9 2 9 1 9 7 0 9 2
24 11 11 3 13 9 0 0 9 7 9 0 9 2 7 3 15 13 13 1 0 9 0 9 2
37 11 11 13 13 9 2 7 1 9 2 16 4 0 9 13 9 9 2 7 11 11 2 13 2 10 9 1 0 10 9 2 15 13 9 2 2 2
7 13 2 16 0 9 13 2
36 0 9 2 0 9 2 9 2 0 9 1 9 7 0 9 0 1 9 13 3 1 0 9 2 0 9 2 0 9 7 0 9 9 9 9 2
17 3 4 3 13 7 13 10 9 7 9 13 3 2 3 13 13 2
8 7 7 3 13 9 1 9 2
18 13 15 0 9 9 2 7 16 13 9 1 9 7 0 9 1 9 2
15 13 10 0 9 9 9 13 2 7 10 0 9 3 13 2
6 15 15 15 13 9 2
6 1 0 9 7 13 2
2 9 9
9 1 9 7 9 13 13 0 9 2
13 15 13 9 1 11 2 3 13 0 9 0 9 2
14 3 9 13 10 0 9 2 2 13 0 9 11 11 2
33 0 9 0 0 9 11 2 9 9 0 0 9 0 1 0 9 2 0 9 0 9 7 3 9 9 3 0 9 7 3 7 9 2
7 15 15 13 3 0 9 2
6 9 13 0 9 9 2
12 1 10 9 15 13 0 9 7 0 0 9 2
12 9 13 0 7 13 15 13 14 0 9 9 2
13 13 7 9 16 9 7 13 0 13 3 10 9 2
23 0 9 3 1 9 9 0 9 13 1 0 9 2 7 9 9 9 2 15 15 13 13 2
19 13 15 7 3 13 0 0 9 2 13 9 15 15 1 9 1 9 9 2
27 1 9 0 9 0 9 13 2 15 13 3 9 2 7 3 3 13 1 9 9 10 9 2 14 3 9 2
11 3 13 1 9 2 15 3 2 15 3 2
33 3 15 13 2 16 9 1 9 13 1 3 0 0 9 2 9 2 15 4 7 9 13 1 0 9 2 7 14 0 9 1 9 2
14 13 1 0 9 2 1 15 10 9 1 0 9 13 2
21 10 9 13 10 9 1 9 9 1 9 2 3 13 15 9 2 15 13 3 13 2
17 1 10 9 15 13 12 3 0 9 2 9 13 2 7 3 13 2
31 0 9 13 1 0 9 2 3 0 9 13 0 2 3 0 2 14 0 2 0 1 0 9 2 3 15 13 13 9 13 2
3 9 1 9
12 1 0 0 9 11 13 1 9 12 9 3 2
17 10 9 15 13 1 9 1 12 7 12 9 2 0 9 2 9 2
15 0 9 9 9 13 3 9 9 2 9 2 9 7 9 2
26 9 3 13 2 15 0 13 1 0 9 2 0 13 7 9 9 2 9 2 7 2 0 2 0 9 2
29 9 7 9 15 13 1 9 2 9 2 9 7 3 7 1 9 13 9 10 9 2 9 2 9 7 15 0 9 2
11 0 9 13 12 9 2 0 3 13 9 2
15 13 15 3 3 9 1 15 2 16 9 15 13 13 3 2
16 3 3 14 13 9 10 0 9 2 15 15 9 13 1 9 2
24 1 0 9 0 9 2 15 15 1 0 9 13 13 0 9 1 0 9 9 2 13 3 9 2
6 10 9 15 7 13 2
20 1 0 9 13 0 7 3 0 9 2 3 15 13 1 0 2 3 7 3 2
14 9 3 0 9 1 9 9 9 15 13 1 9 9 2
11 9 1 10 9 13 7 13 0 15 13 2
27 9 0 9 11 11 7 11 11 15 1 9 9 3 13 1 11 7 1 11 2 1 11 13 0 12 9 2
4 11 16 9 9
17 2 1 15 13 9 16 9 0 9 3 1 9 2 2 13 11 2
17 2 1 11 9 10 9 13 3 3 2 16 13 1 0 9 9 2
23 16 13 0 9 2 13 3 3 13 2 16 13 9 1 11 2 13 11 7 11 2 2 2
21 13 15 9 0 9 2 15 13 0 9 0 1 9 2 3 0 9 1 0 9 2
9 10 9 15 3 13 7 1 15 2
21 7 16 15 13 3 3 2 16 3 9 3 3 3 13 2 3 15 15 13 2 2
16 7 15 14 10 9 13 10 9 13 2 3 16 13 0 9 2
28 2 13 9 2 16 4 15 9 13 13 9 9 2 1 15 13 12 9 2 7 9 2 15 3 13 1 9 2
7 3 0 13 9 0 9 2
7 15 13 1 9 3 0 2
18 13 15 9 2 15 13 9 9 2 7 7 13 7 0 12 2 2 2
10 3 7 13 15 2 15 13 9 2 2
24 1 15 0 0 9 13 1 9 9 2 13 0 9 7 9 13 1 9 2 0 1 0 9 2
18 3 1 9 2 16 1 9 4 13 10 0 9 2 3 9 13 3 2
22 1 0 9 15 9 13 9 1 9 1 9 7 15 15 13 1 9 2 16 13 0 2
20 2 10 9 2 3 1 9 2 15 13 3 13 9 2 9 7 9 1 9 2
8 3 13 2 2 13 3 11 2
27 2 1 9 13 3 0 9 7 13 15 2 16 1 9 13 0 3 3 13 9 2 16 13 10 9 2 2
19 10 9 1 9 9 2 9 7 9 1 9 1 9 15 3 3 9 13 2
10 1 0 15 3 9 1 10 9 13 2
3 9 1 9
13 0 0 2 9 15 1 9 13 1 9 0 9 2
9 10 9 3 7 13 1 10 9 2
28 9 9 2 11 2 11 1 9 1 11 3 13 2 16 10 9 15 13 1 12 9 1 11 2 7 3 3 2
10 13 15 7 1 11 2 7 1 11 2
22 1 9 1 0 9 15 9 0 0 2 9 13 1 9 2 7 14 1 10 0 9 2
23 13 15 2 16 16 15 9 15 13 2 3 13 7 9 7 9 1 12 7 12 9 13 2
11 16 13 9 13 3 3 2 9 3 13 2
12 1 15 0 0 2 9 13 10 0 0 9 2
8 0 9 15 3 10 9 13 2
42 9 0 9 7 9 9 2 11 11 13 1 0 9 9 9 2 9 0 9 1 11 3 0 0 2 9 13 1 0 9 7 13 0 9 2 7 10 9 3 3 13 2
15 9 2 11 11 13 9 9 0 9 9 0 9 1 11 2
23 1 15 15 2 1 9 1 9 0 1 9 2 9 1 9 0 0 2 9 13 3 3 2
21 2 13 15 3 9 2 7 16 13 2 7 9 1 9 9 7 9 13 3 0 2
12 13 15 3 0 9 2 9 7 0 9 2 2
14 9 13 0 0 2 9 13 9 0 9 9 0 9 2
40 3 7 13 13 9 2 16 10 9 15 13 9 2 16 13 0 9 2 16 9 13 13 3 0 9 2 16 13 9 1 15 2 16 9 9 13 13 3 9 2
8 15 15 13 0 9 0 9 2
7 13 9 2 7 7 1 9
22 1 9 11 15 9 13 13 1 9 9 7 1 12 9 2 3 7 9 15 15 13 2
10 3 13 3 2 16 4 15 9 13 2
5 9 15 13 13 2
12 9 0 1 9 13 2 7 1 9 0 9 2
31 3 0 13 9 3 0 9 2 0 13 15 1 9 9 2 15 15 9 13 3 15 7 1 9 2 16 9 9 13 0 2
28 9 2 15 13 1 9 2 13 3 9 2 15 15 13 1 9 13 2 7 3 15 13 10 9 7 1 9 2
8 3 15 9 7 10 9 13 2
34 3 15 13 13 2 16 1 9 0 9 0 9 9 13 9 9 2 16 13 15 0 9 13 14 1 12 9 2 13 1 9 0 9 2
8 14 3 13 9 9 1 9 2
21 13 9 2 1 0 9 2 9 7 9 2 2 3 10 9 3 13 0 0 9 2
16 13 15 2 16 9 13 0 9 9 7 9 9 13 0 9 2
10 10 9 15 13 3 13 3 9 9 2
15 2 9 9 13 0 0 9 2 2 13 3 9 2 11 2
17 2 9 13 13 1 15 2 16 15 4 0 9 13 3 12 9 2
10 3 7 13 9 2 15 13 9 13 2
9 0 9 13 1 3 0 9 2 2
18 3 2 15 13 9 0 2 15 13 0 10 9 7 0 0 0 9 2
21 1 3 0 9 15 13 13 2 16 9 13 13 3 3 2 3 13 3 3 13 2
19 13 14 1 15 2 3 3 15 15 13 10 0 9 2 13 1 9 2 2
13 1 0 9 15 9 13 13 1 10 9 13 3 15
3 9 1 9
13 13 9 2 15 13 9 11 2 11 1 0 9 2
18 3 15 13 0 2 16 3 3 10 9 13 2 15 0 9 15 13 2
51 11 4 13 3 1 12 9 2 7 9 10 9 3 13 1 15 3 2 16 1 0 9 2 7 1 11 3 3 13 13 2 16 9 9 13 9 2 7 15 15 1 15 13 1 9 10 12 0 9 13 2
11 9 11 7 11 13 9 9 13 1 9 2
33 1 12 9 1 15 2 15 15 1 9 3 13 9 9 2 1 0 9 1 15 2 15 15 13 7 13 0 1 9 1 0 9 2
26 1 9 4 15 13 13 11 1 11 7 11 1 11 3 7 13 15 2 15 9 13 7 15 3 13 2
19 13 15 7 2 16 16 13 9 0 0 9 2 13 7 9 3 15 13 2
21 16 1 11 2 7 1 0 9 4 3 9 13 1 0 9 2 15 13 0 9 2
14 7 10 0 9 13 0 2 16 0 2 16 10 0 2
10 0 9 15 3 13 9 9 7 9 2
17 0 9 9 3 13 1 9 3 1 10 9 2 1 15 13 9 2
10 7 15 2 1 15 13 9 2 13 2
10 7 13 9 1 9 1 9 3 0 2
32 1 11 13 10 9 2 15 15 13 9 1 0 9 7 13 13 2 16 0 9 15 11 13 3 3 2 16 4 15 13 9 2
17 3 13 11 0 9 0 7 0 2 16 10 9 13 1 0 9 2
6 15 15 1 15 13 2
31 13 3 3 0 2 16 9 13 0 9 3 1 9 2 11 11 7 11 11 13 1 9 2 15 13 3 9 2 3 3 2
15 7 0 7 0 13 9 2 1 15 4 3 13 15 15 2
23 12 1 9 9 11 13 9 9 1 9 0 9 7 9 2 7 15 1 12 9 9 11 2
23 1 9 2 16 15 11 7 11 1 15 15 3 3 13 2 3 13 2 16 13 0 9 2
7 1 0 9 15 13 15 2
23 12 9 13 0 9 2 15 15 13 1 0 9 2 12 13 9 9 2 0 0 9 13 2
9 1 12 9 13 0 9 0 9 2
32 16 9 0 2 7 7 0 15 13 1 0 9 0 9 7 13 1 9 2 1 12 15 13 7 1 0 9 7 1 0 9 2
42 3 1 11 2 16 1 11 13 0 9 2 15 4 13 9 1 9 3 2 3 1 9 1 3 0 9 9 1 9 2 1 10 0 9 2 0 9 7 9 10 9 2
3 13 9 2
38 14 1 0 9 2 7 7 1 0 9 15 13 2 16 9 13 1 0 9 10 9 2 16 1 9 3 3 0 12 9 13 13 10 9 1 9 0 2
35 13 2 16 13 15 3 10 9 1 0 9 9 2 15 15 13 0 13 2 16 10 9 13 13 15 2 3 3 7 10 9 13 0 13 2
15 7 14 3 16 11 2 11 7 16 11 2 7 16 9 2
5 15 15 13 1 9
8 9 11 11 2 0 14 0 9
27 1 0 9 13 1 9 11 7 11 1 11 9 7 0 9 2 0 9 0 9 7 3 0 9 11 11 2
21 10 9 2 15 13 0 7 0 9 9 2 4 13 13 13 14 1 0 9 9 2
3 13 11 2
2 3 2
17 10 9 13 9 2 13 1 9 2 13 0 9 7 9 9 13 2
22 3 15 2 16 4 13 0 2 13 2 13 15 0 2 7 1 0 9 13 3 9 2
9 7 3 13 3 1 15 0 9 2
26 13 4 2 16 9 11 13 1 12 9 1 9 12 10 9 1 9 2 13 4 3 1 0 0 9 2
24 9 2 16 0 9 13 9 9 2 13 14 1 9 2 7 13 0 13 2 16 15 13 9 2
36 1 9 2 3 13 15 3 16 1 15 2 3 13 2 16 9 13 12 2 12 9 2 7 15 13 1 0 9 2 7 3 13 1 12 9 2
6 15 13 1 0 9 2
15 10 0 9 13 7 1 15 2 15 13 9 9 2 2 2
8 11 13 13 3 1 15 0 2
14 1 0 9 3 13 2 16 13 0 2 16 13 9 2
19 7 3 10 9 1 0 9 13 2 3 0 9 1 9 2 1 0 9 2
15 13 1 15 3 10 9 2 15 4 13 10 0 0 9 2
18 0 13 10 0 9 7 9 13 16 15 0 2 15 15 9 3 13 2
23 7 15 13 13 0 9 2 3 13 3 9 9 7 9 2 7 0 9 13 0 0 9 2
18 3 2 11 2 7 16 10 9 13 9 9 2 13 3 3 10 9 2
19 13 4 1 15 2 16 13 1 9 1 10 9 1 0 9 1 0 9 2
24 13 15 10 0 9 9 1 9 7 9 2 0 1 9 2 13 15 13 7 15 15 3 13 2
12 13 10 9 9 10 9 9 2 7 0 9 2
9 13 2 16 13 15 0 9 9 2
11 9 9 1 9 12 13 0 7 3 13 2
15 3 13 0 9 1 0 9 2 1 0 0 9 3 0 2
14 15 13 3 1 15 2 3 15 1 15 1 9 13 2
19 16 4 9 13 0 9 2 3 4 15 13 13 3 3 2 3 2 3 2
11 13 1 0 2 16 3 13 9 1 9 2
11 13 0 9 9 7 3 13 13 0 9 2
18 9 7 13 14 1 0 9 2 16 9 7 9 13 10 9 1 9 2
8 0 9 1 9 15 15 13 2
10 13 1 12 0 9 2 13 0 9 2
13 3 13 10 9 2 15 13 1 2 0 9 2 2
12 10 9 13 10 0 9 2 15 15 13 9 2
18 7 1 15 13 7 15 15 2 15 4 13 10 9 13 1 0 9 2
11 3 13 9 1 0 2 0 7 0 9 2
18 1 15 13 0 2 16 13 9 2 13 13 2 13 13 2 15 13 2
28 15 13 14 0 9 2 0 9 13 1 11 2 11 2 1 11 2 1 0 11 2 1 0 9 7 1 11 2
8 3 13 9 9 1 0 9 2
13 15 13 16 0 9 2 1 15 9 13 14 9 2
7 13 15 3 2 7 3 2
19 1 9 2 16 9 13 3 2 16 4 13 9 2 3 4 15 13 13 2
17 7 16 4 13 2 13 0 1 0 2 2 3 13 15 3 0 2
27 10 0 9 2 3 9 9 2 13 0 9 2 0 9 9 7 13 15 1 0 9 2 0 3 9 9 2
18 15 1 9 0 9 13 9 2 0 10 9 13 1 3 0 1 9 2
13 15 4 15 13 2 13 3 1 9 9 16 9 2
16 10 9 13 3 0 1 11 2 3 13 9 1 9 7 9 2
10 0 1 15 13 1 9 3 0 9 2
13 13 15 15 2 16 10 0 9 13 0 0 9 2
19 16 15 3 13 1 0 0 9 2 13 15 2 15 4 10 0 9 13 2
12 9 15 3 13 2 7 13 3 0 0 9 2
10 3 9 2 16 13 13 1 9 9 2
3 3 13 2
39 7 13 15 0 2 16 13 15 9 7 3 13 1 9 2 7 16 15 0 9 13 1 9 7 15 15 3 13 1 0 9 7 13 0 9 1 0 9 2
5 15 7 15 13 2
20 13 3 3 0 13 2 16 9 1 9 13 2 3 3 9 2 9 13 13 2
28 1 12 1 10 9 4 0 9 13 1 9 2 15 15 13 2 16 15 13 9 0 3 10 9 1 12 9 2
13 13 15 0 9 2 13 15 3 9 9 7 9 2
5 3 9 7 9 2
19 13 9 10 9 7 9 2 15 15 13 1 0 9 1 9 1 0 9 2
19 15 10 9 13 1 3 0 2 7 15 3 13 15 2 15 15 13 9 2
26 16 0 9 13 1 9 2 7 16 13 1 0 9 2 7 13 13 0 9 2 15 3 13 9 9 2
16 7 0 9 13 1 10 9 9 15 2 3 15 13 1 9 2
17 7 15 13 2 16 0 9 13 3 0 2 7 15 3 13 9 2
17 16 15 13 1 9 0 9 2 13 0 9 1 0 9 7 9 2
9 9 13 3 3 7 3 0 9 2
12 1 15 13 7 9 13 13 10 0 0 9 2
10 1 15 9 1 9 1 9 13 0 2
18 15 2 16 9 13 15 2 16 13 15 3 0 2 13 1 3 0 2
18 3 16 0 9 1 10 2 16 15 15 3 13 2 13 1 3 0 2
21 13 15 3 2 16 9 7 9 3 15 13 2 9 9 1 10 9 13 3 0 2
12 13 9 0 9 7 9 1 2 0 9 2 2
22 13 15 0 1 9 2 1 15 1 9 13 9 2 15 4 1 9 3 3 3 13 2
14 13 2 16 0 9 13 15 2 15 1 9 9 13 2
7 15 13 15 2 15 13 2
16 3 3 15 13 2 13 7 9 0 9 2 13 3 0 9 2
11 15 13 1 9 2 15 13 1 9 0 2
12 13 4 15 13 2 0 15 13 13 10 9 2
11 13 14 1 15 2 15 15 13 10 9 2
13 13 7 9 2 16 10 9 3 3 13 1 9 2
17 3 15 13 10 9 2 16 4 15 13 13 1 15 2 15 13 2
19 3 16 15 9 13 13 2 7 13 0 1 15 13 7 3 1 15 13 2
23 15 10 0 9 3 13 1 9 1 9 2 0 7 0 9 2 0 9 3 13 10 9 2
15 15 15 13 13 1 0 9 2 7 1 10 9 3 14 2
16 9 1 10 2 15 15 13 1 0 9 9 2 13 1 0 2
28 15 10 9 13 1 9 2 15 3 13 1 10 9 3 7 1 9 2 16 13 1 9 0 11 0 2 0 2
8 13 15 9 13 14 0 9 2
10 10 9 13 3 0 7 13 3 0 2
12 0 9 13 7 0 16 10 12 12 0 9 2
22 1 9 1 9 0 9 2 16 0 0 2 13 3 0 13 2 16 15 13 15 0 2
14 3 4 13 9 0 0 9 0 15 0 9 1 15 2
16 7 15 13 2 16 1 9 9 4 13 9 1 9 7 9 2
19 9 3 13 9 2 9 7 9 2 7 9 2 9 0 9 7 0 9 2
6 10 0 9 13 9 2
16 1 15 13 2 13 2 16 0 9 13 13 1 0 0 9 2
8 3 1 9 2 9 2 9 2
13 15 3 3 13 2 1 15 13 0 9 0 9 2
12 9 13 0 13 15 2 13 2 13 3 0 2
18 0 9 1 0 9 13 1 15 2 15 13 2 9 15 13 0 9 2
9 1 9 10 9 15 7 13 9 2
23 15 4 1 9 2 15 13 1 15 13 9 0 9 2 13 10 9 13 2 13 1 15 2
3 0 9 2
2 9 2
14 9 13 2 15 13 2 7 13 1 15 3 10 9 2
8 0 9 1 9 13 3 0 2
15 3 15 13 2 16 13 15 0 9 2 7 9 13 3 2
8 13 15 3 1 9 1 9 2
13 9 13 0 9 2 7 13 15 3 13 0 9 2
25 16 4 15 9 13 3 2 16 1 15 9 4 13 1 9 7 9 2 3 13 15 3 1 9 2
17 7 16 15 13 2 16 15 3 13 0 9 2 13 1 0 9 2
21 13 4 15 3 13 9 9 1 15 2 16 4 3 3 9 13 2 13 1 15 2
9 13 4 15 13 13 7 1 9 2
11 13 3 3 0 9 1 9 2 1 9 2
9 13 15 3 1 0 2 0 9 2
17 4 13 11 9 10 0 9 2 7 15 13 0 9 16 3 11 2
17 1 9 9 9 3 13 0 9 2 16 13 0 13 10 0 9 2
15 1 12 9 13 0 2 16 15 1 0 2 0 9 13 2
19 7 13 15 3 9 1 9 3 15 0 9 3 2 3 4 15 0 13 2
22 13 1 9 2 0 9 2 3 0 9 1 0 9 2 3 13 1 0 9 12 9 2
28 13 15 15 9 2 15 1 0 9 13 9 2 16 9 13 2 3 9 1 11 1 9 1 11 2 3 3 2
20 0 9 13 0 2 13 9 9 2 15 7 1 9 1 11 13 12 12 3 2
5 15 4 11 13 2
3 0 9 2
5 9 2 9 7 3
5 9 1 9 7 9
16 11 2 3 0 0 0 9 1 9 2 3 13 12 2 9 2
12 13 15 9 1 9 12 9 0 9 1 9 2
13 13 1 9 9 7 9 1 0 9 0 0 9 2
29 13 1 15 9 9 2 0 9 9 2 9 10 9 2 9 7 0 9 2 9 9 2 9 9 3 16 0 9 2
24 1 9 1 15 11 13 9 2 15 13 1 0 2 4 15 9 13 3 2 7 15 9 13 2
8 4 9 9 13 2 7 13 2
10 3 3 13 9 9 0 0 9 9 2
5 13 1 9 9 2
6 3 4 15 13 13 2
6 3 0 13 9 9 2
8 3 15 10 0 9 13 13 2
9 3 15 9 3 13 1 0 9 2
6 3 13 9 3 9 2
14 3 13 0 9 9 1 15 2 16 4 15 13 13 2
7 3 13 0 9 3 0 2
9 13 13 9 0 9 1 10 9 2
7 13 0 13 0 9 9 2
9 9 1 10 9 13 9 1 9 2
31 13 9 9 1 0 9 13 2 15 13 2 3 4 13 2 3 13 2 10 15 13 9 7 15 13 2 7 13 2 13 2
12 0 9 4 13 3 0 9 1 15 9 9 2
18 1 9 1 12 9 2 0 7 0 2 9 11 13 9 0 0 9 2
17 10 9 15 13 1 9 9 2 0 9 2 9 2 9 7 9 2
15 13 3 0 2 16 13 9 1 9 0 9 7 0 9 2
3 7 3 2
15 9 0 9 1 10 9 13 9 1 11 2 11 7 11 2
6 3 9 13 14 12 2
17 13 0 9 1 9 7 9 2 15 13 3 12 1 10 0 9 2
23 13 9 9 2 9 2 9 2 7 3 2 13 1 12 9 9 10 9 0 9 1 11 2
12 13 15 12 9 2 1 10 3 0 9 12 2
28 1 15 13 3 9 2 16 3 13 13 10 9 1 9 12 2 12 9 2 15 4 13 15 1 10 9 13 2
16 4 2 14 1 15 13 7 13 2 14 15 1 10 9 9 2
4 7 15 0 2
15 9 2 0 9 1 15 13 3 2 13 2 14 14 9 2
13 0 13 2 16 15 3 3 13 3 0 9 9 2
2 0 9
24 0 9 13 3 0 9 0 2 16 9 13 1 12 7 12 9 9 7 1 10 9 15 13 2
9 13 1 15 9 2 15 13 9 2
9 7 13 1 10 9 0 1 9 2
7 3 9 9 9 1 9 2
21 12 1 9 9 0 9 13 2 16 9 9 1 9 13 0 1 9 0 16 0 2
11 9 0 9 7 0 9 15 13 9 9 2
20 16 4 10 9 13 0 16 12 2 9 13 1 0 9 7 9 15 3 13 2
13 16 4 13 0 16 12 2 4 15 9 13 3 2
12 0 9 9 13 2 16 15 9 13 3 12 2
15 7 9 13 2 16 15 0 9 13 1 12 9 0 9 2
17 16 4 3 13 13 10 9 9 0 9 2 3 12 9 9 13 2
14 13 15 1 0 9 2 7 15 13 2 15 15 13 2
23 13 0 2 16 4 13 13 1 9 0 1 0 9 9 9 2 15 4 9 13 0 9 2
10 0 9 3 0 9 9 4 13 0 2
22 3 9 13 2 16 9 0 9 0 1 0 9 13 13 3 12 0 1 9 0 9 2
5 13 0 9 9 2
8 7 0 7 3 0 9 9 2
5 9 15 13 10 2
17 15 13 3 0 9 2 16 15 0 0 0 2 9 9 3 13 2
3 1 9 2
5 9 2 7 9 2
12 1 11 13 9 0 9 1 0 9 1 0 9
16 9 1 11 15 1 9 13 7 3 13 2 1 12 9 12 2
26 3 4 13 1 10 9 13 9 1 9 2 16 4 15 9 13 0 0 9 11 16 10 9 0 9 2
57 10 3 0 9 13 14 3 0 13 2 0 0 9 11 11 1 11 1 0 9 1 9 2 0 9 7 9 1 15 3 13 3 3 9 16 9 1 9 9 2 15 15 13 0 9 1 0 9 1 0 9 7 9 1 0 11 2
32 1 0 2 3 0 16 0 9 1 9 11 11 15 3 1 9 13 9 9 15 9 2 0 9 2 9 11 7 9 0 11 2
33 0 9 0 9 13 13 9 2 1 15 4 15 13 3 3 9 7 15 4 15 13 12 1 9 0 0 9 9 11 1 0 9 2
27 0 9 15 13 13 3 1 12 2 0 9 9 7 9 1 0 9 13 3 16 0 7 3 13 0 9 2
6 7 13 0 15 13 2
23 9 15 7 3 13 1 15 2 3 0 7 0 13 10 9 13 7 3 15 13 15 13 2
19 9 9 13 0 9 9 0 9 2 15 13 2 1 15 1 0 9 13 2
20 0 1 9 13 1 0 9 3 1 15 2 16 10 9 4 9 1 11 13 2
33 9 9 13 9 0 9 9 9 2 16 1 9 13 1 15 2 16 15 1 9 9 13 1 9 9 9 2 14 7 1 10 9 2
11 16 10 0 9 3 13 9 9 15 0 2
29 9 11 1 10 9 13 2 16 16 4 15 0 9 9 13 13 9 0 2 3 13 9 1 9 0 9 3 0 2
38 13 2 14 3 9 1 9 10 9 2 13 1 9 9 1 15 13 2 16 4 15 3 13 9 1 9 0 0 9 7 16 4 1 15 13 10 9 2
27 9 15 10 9 3 3 13 9 13 0 0 9 2 15 13 2 16 9 9 13 3 0 1 0 9 9 2
18 9 1 9 9 13 3 13 2 7 1 10 9 13 1 11 15 0 2
42 3 15 1 15 13 1 9 7 9 0 9 1 15 2 16 0 9 13 3 0 9 2 15 3 13 2 14 0 1 9 7 16 9 13 0 13 1 0 9 0 9 2
15 9 10 9 13 7 11 11 11 2 9 0 9 0 9 2
23 10 9 13 9 10 9 7 13 2 16 15 0 9 13 2 16 0 9 13 3 3 13 2
17 9 3 0 9 1 9 9 13 3 12 1 0 9 9 1 11 2
23 3 0 13 3 0 9 9 0 9 2 15 13 1 15 2 16 7 9 13 13 0 9 2
31 13 4 3 0 13 1 10 0 9 2 15 4 13 0 9 0 9 2 15 4 3 0 0 9 13 9 1 9 9 0 2
29 1 9 0 15 0 9 0 9 13 2 7 3 1 10 9 2 7 3 0 9 1 15 2 3 13 7 13 9 2
21 3 0 9 11 13 9 10 9 2 15 13 9 0 13 9 9 14 1 9 9 2
21 0 9 3 13 0 9 0 9 0 9 1 9 9 0 7 0 9 0 0 9 2
28 9 9 15 13 1 15 2 16 4 13 3 13 1 9 7 0 9 7 13 15 1 0 9 0 9 1 11 2
41 1 0 0 9 13 0 9 0 9 11 11 9 1 15 2 16 15 13 13 1 0 9 2 13 4 13 15 0 2 3 15 2 2 1 9 2 16 13 13 15 2
21 13 1 15 9 1 9 2 15 13 13 1 9 7 13 15 13 1 9 7 9 2
12 1 9 9 13 9 3 0 2 7 2 2 2
7 7 9 13 1 0 9 2
8 3 15 13 3 1 9 9 2
18 3 3 3 13 1 9 2 7 9 13 2 16 15 15 13 3 13 2
8 13 1 15 3 14 12 9 2
2 9 11
27 15 13 13 9 2 11 11 2 9 2 13 3 7 1 9 15 3 3 13 0 9 2 16 3 3 0 2
12 13 15 0 9 12 9 2 15 13 11 11 2
5 13 9 0 9 2
9 12 5 9 11 13 0 1 9 2
7 3 0 13 14 12 5 2
21 12 5 1 15 13 9 9 11 2 9 1 9 11 3 13 2 1 12 5 2 2
11 0 9 9 11 3 13 9 1 0 9 2
15 0 9 13 3 0 2 16 14 15 15 3 13 1 9 2
33 0 2 0 9 9 2 0 1 11 2 13 3 1 11 3 1 9 11 11 0 9 2 1 15 15 13 9 1 0 7 0 9 2
26 9 9 13 9 1 0 9 2 7 3 9 1 15 2 15 1 15 2 12 9 1 9 2 3 13 2
26 13 3 9 2 1 0 9 0 7 3 2 3 1 0 9 2 7 0 2 2 9 2 9 2 9 2
24 1 10 9 13 2 16 12 0 9 13 3 0 9 2 15 7 1 0 9 13 3 0 9 2
7 9 15 1 0 0 9 2
60 0 9 13 1 0 9 3 3 2 3 7 13 1 9 0 9 7 0 9 11 11 2 0 9 7 9 11 11 2 11 7 9 7 3 0 9 11 11 2 1 9 0 1 11 7 3 0 1 11 2 13 1 12 9 9 11 3 0 9 2
4 13 15 13 0
19 1 10 9 7 9 15 13 13 9 2 14 9 2 13 9 11 2 11 2
2 11 2
17 1 9 11 11 13 1 10 9 1 9 0 9 1 9 1 9 2
5 11 15 9 13 2
16 9 15 13 12 9 2 13 15 1 15 7 1 9 13 3 2
5 9 15 13 9 2
9 11 4 13 1 0 9 9 9 2
11 13 3 2 16 10 9 13 0 9 9 2
23 0 9 2 3 9 13 9 7 15 3 13 7 13 1 15 13 2 13 1 11 10 9 2
10 13 15 9 9 11 11 2 11 2 2
15 7 15 13 13 9 1 9 9 9 0 9 1 0 9 2
16 1 3 0 9 13 9 13 2 16 10 9 13 2 0 2 2
26 11 13 13 2 16 4 15 1 2 9 2 1 9 2 16 9 4 13 1 9 7 9 2 3 13 2
19 0 9 11 11 2 9 1 9 2 1 9 9 2 9 2 1 9 13 2
17 2 13 2 15 13 9 2 13 3 0 7 3 0 2 2 13 2
34 11 11 2 9 9 0 9 1 11 7 9 9 0 9 9 2 13 15 1 9 9 2 2 13 1 15 2 16 0 9 0 9 13 2
7 2 9 13 1 9 9 2
23 1 11 3 13 0 9 2 15 4 15 13 13 9 9 16 0 7 0 2 2 13 11 2
11 0 9 9 3 14 13 0 9 7 9 2
14 2 13 15 9 9 2 7 14 9 2 2 13 11 2
8 9 11 3 13 9 6 9 2
22 13 2 16 9 2 15 1 15 13 2 15 3 9 13 2 16 4 1 15 4 13 2
18 9 2 11 15 13 2 16 3 10 9 1 9 13 9 9 0 13 2
20 11 15 7 13 2 16 1 9 9 2 15 1 15 4 13 16 1 11 2 2
11 2 0 9 3 13 13 2 2 13 11 2
17 2 1 10 9 13 9 0 9 2 9 7 9 9 1 9 12 2
4 13 15 9 2
16 13 13 9 3 2 3 13 1 12 9 2 2 13 9 11 2
1 9
25 9 15 3 13 1 3 0 9 2 15 7 3 13 0 2 16 9 13 3 7 3 3 9 0 2
35 13 15 3 0 9 3 0 9 2 1 15 15 3 0 9 9 13 1 0 2 13 15 3 1 9 0 2 0 2 1 15 0 7 0 2
8 0 9 13 9 3 0 9 2
14 1 10 9 13 3 13 0 9 2 9 7 0 9 2
24 3 15 0 2 13 2 14 3 10 9 2 13 13 15 2 15 15 13 2 3 3 7 3 2
23 16 13 2 16 13 2 7 13 3 3 2 16 0 9 9 10 9 1 0 9 3 13 2
23 3 15 7 13 13 2 16 10 0 9 10 9 13 7 1 9 15 1 15 13 10 9 2
25 13 15 2 7 15 15 3 13 2 16 4 15 15 13 1 9 2 3 10 0 0 9 3 13 2
26 15 3 13 2 16 10 9 3 13 10 0 9 2 1 15 4 13 4 1 10 9 13 1 0 9 2
6 10 9 1 15 13 2
16 13 15 3 9 9 2 7 10 9 13 13 10 3 0 9 2
28 15 1 15 13 1 9 3 3 0 9 9 2 15 15 13 15 10 9 2 15 15 3 3 13 9 0 9 2
35 16 13 2 13 7 15 2 3 13 2 9 7 9 2 16 13 1 10 9 2 16 4 15 13 1 10 9 2 1 15 15 0 9 13 2
41 9 13 9 9 0 1 15 7 13 0 9 2 16 15 3 13 15 2 15 13 0 2 15 0 13 0 9 10 3 0 9 2 15 15 3 13 1 0 9 9 2
12 13 15 3 3 2 7 3 13 15 3 0 2
11 7 13 2 13 2 14 15 1 10 9 2
20 7 13 3 10 9 9 2 16 4 3 13 2 16 15 9 9 15 9 13 2
18 9 11 7 11 13 3 1 12 9 9 1 0 9 1 11 2 11 2
24 9 11 7 11 0 7 0 13 9 1 0 9 9 1 11 7 0 0 9 9 9 5 9 2
16 1 9 15 13 3 1 9 3 1 9 7 1 9 0 9 2
24 11 11 2 9 9 2 15 0 9 13 2 2 7 1 10 9 1 9 15 13 1 15 2 2
3 9 0 9
4 11 2 11 2
15 1 9 9 15 3 1 0 9 11 13 15 10 0 9 2
25 1 9 11 13 13 9 11 7 1 0 9 0 9 11 7 0 9 11 2 15 14 1 9 13 2
21 9 11 2 15 15 1 9 13 2 1 9 13 4 2 16 4 13 14 1 9 2
18 3 13 9 7 9 11 2 15 15 1 9 9 3 13 1 9 9 2
22 0 9 13 9 11 1 9 0 9 11 2 15 1 9 13 2 7 13 9 1 9 2
2 9 9
16 13 4 3 13 2 16 4 9 1 9 13 1 9 0 9 2
10 9 11 11 1 10 9 9 9 1 9
10 10 9 13 1 15 9 13 3 0 2
14 9 11 11 1 9 1 9 9 9 9 12 2 0 9
15 16 15 13 2 15 4 15 13 7 15 4 15 13 9 2
13 0 9 9 0 9 11 11 1 10 9 9 1 11
22 13 0 9 9 9 9 2 16 15 15 15 3 13 9 1 9 1 9 1 9 0 2
11 9 11 11 11 1 9 9 11 1 9 9
5 3 3 13 9 2
12 3 7 15 2 1 15 13 2 16 13 0 2
10 9 9 11 11 11 1 10 9 1 9
18 13 4 15 2 16 15 15 13 2 7 10 0 9 13 0 2 0 2
17 15 15 13 2 15 3 3 3 13 2 9 2 7 15 3 13 2
11 9 9 11 11 1 9 9 1 9 10 9
23 0 9 13 9 1 0 9 10 9 2 9 0 1 0 9 2 9 7 0 15 0 9 2
16 1 9 0 9 0 7 0 9 1 9 1 0 9 11 11 11
22 15 13 0 9 2 16 4 13 2 16 9 11 13 1 9 0 9 0 9 7 11 2
22 7 9 1 9 2 1 10 3 13 9 2 4 15 13 4 13 7 13 9 7 13 2
31 9 0 0 9 11 2 11 11 11 1 9 9 11 2 16 9 4 13 13 14 9 2 1 10 9 4 13 13 10 0 9
5 1 9 13 0 9
16 1 0 9 15 3 13 1 9 1 9 2 13 9 11 2 11
5 0 11 2 11 2
19 0 9 0 9 11 1 0 11 4 1 0 9 13 1 0 9 0 9 2
8 11 15 13 9 9 11 11 2
31 13 2 16 1 9 2 3 1 9 0 9 2 9 0 9 11 7 9 9 1 11 13 0 9 0 9 2 15 3 13 2
24 2 0 13 7 15 2 16 9 1 0 11 4 13 1 0 9 16 0 9 2 2 13 9 2
10 0 9 4 3 13 9 9 0 9 2
36 0 9 9 1 11 4 13 1 9 9 15 0 9 1 9 11 2 9 1 0 9 4 7 1 9 3 13 1 9 2 3 9 1 9 13 2
13 7 9 1 9 13 1 9 9 1 9 1 9 2
42 9 1 9 9 0 9 11 13 7 15 2 16 9 2 15 15 13 1 11 2 9 3 13 9 2 3 7 0 9 2 16 1 9 13 2 7 3 7 1 0 9 2
12 2 13 3 13 9 10 9 2 2 13 9 2
19 16 0 9 13 1 12 2 9 9 9 9 2 11 13 9 1 0 9 2
21 2 13 15 1 9 12 2 3 15 13 2 2 13 11 9 0 9 9 11 11 2
19 0 1 15 13 2 16 4 1 9 11 7 0 9 13 3 3 0 9 2
17 11 15 13 2 16 9 0 9 1 0 9 13 13 1 10 9 2
15 2 13 3 0 2 13 0 9 2 2 13 1 10 9 2
18 9 0 9 13 14 1 0 9 9 2 7 7 1 3 0 9 9 2
21 2 14 0 2 15 4 9 13 1 9 2 13 9 1 9 9 2 2 13 11 2
3 13 0 9
8 9 9 15 1 11 13 1 9
2 11 2
31 1 9 2 15 1 0 9 0 9 15 13 13 0 0 9 2 13 11 2 15 13 1 12 9 2 9 1 11 9 11 2
19 1 9 13 11 13 7 1 0 9 2 1 9 10 9 13 9 9 11 2
24 1 0 9 13 9 0 9 11 11 0 2 2 1 1 0 0 9 4 13 9 9 1 11 2
12 0 13 9 1 11 2 16 7 9 1 11 2
8 1 0 9 4 13 9 9 2
25 9 1 11 2 12 2 12 2 9 2 9 2 2 3 13 1 9 2 7 13 1 15 9 2 2
16 9 0 9 9 13 11 9 9 2 1 9 7 15 13 9 2
24 11 0 9 9 13 1 0 9 2 11 15 9 9 13 9 2 7 7 11 13 1 9 11 2
29 2 1 9 13 0 0 9 7 3 11 15 1 0 9 13 1 9 9 1 9 0 9 9 2 2 13 0 9 2
25 0 9 11 2 12 2 9 2 12 9 2 12 9 2 12 9 2 9 12 2 12 2 12 9 2
24 13 2 11 2 11 2 2 11 2 11 2 1 9 1 11 2 12 13 1 9 1 11 2 2
14 13 2 11 2 11 2 2 11 2 0 2 11 2 2
4 9 13 3 9
7 11 14 1 0 9 9 13
2 11 2
24 1 9 13 1 9 3 1 12 9 9 3 15 13 1 0 9 0 9 9 9 11 11 11 2
9 2 9 13 3 0 2 2 13 2
29 9 0 9 1 9 0 9 2 9 1 11 2 11 11 7 9 1 0 0 2 11 11 2 7 1 9 3 13 2
22 2 0 9 13 3 0 7 0 2 16 9 4 13 3 1 9 2 2 13 0 9 2
11 0 9 11 1 0 9 13 0 0 9 2
12 7 7 13 9 9 1 9 11 1 9 9 2
6 2 3 15 15 13 2
19 16 9 13 0 9 0 7 1 9 13 3 9 1 15 2 2 13 11 2
13 1 0 0 9 1 11 13 7 0 9 0 9 2
30 1 12 0 9 4 13 11 2 11 7 0 2 13 13 11 7 1 0 0 9 15 13 9 7 11 2 9 9 9 2
7 2 13 13 3 0 9 2
12 3 16 4 15 13 1 15 2 2 13 11 2
7 0 13 7 0 9 9 2
8 9 3 3 13 1 0 9 2
6 2 9 13 0 9 2
13 7 9 1 11 3 13 2 2 13 9 11 11 2
26 0 9 9 11 2 12 2 9 2 12 9 2 12 9 2 12 9 2 9 12 2 12 2 12 9 2
12 13 2 11 7 11 2 13 1 9 9 2 2
9 13 2 11 2 9 1 11 2 2
4 1 9 1 9
7 11 13 9 0 14 1 11
2 11 2
14 3 9 2 10 9 13 1 0 0 9 9 1 11 2
7 10 0 9 3 9 13 2
29 2 16 13 9 2 13 15 7 13 3 2 13 2 2 13 3 9 0 9 11 11 11 7 0 9 11 11 11 2
15 0 0 9 9 13 3 14 1 0 9 1 0 9 9 2
9 10 0 9 15 7 1 9 13 2
18 2 13 3 13 9 2 2 13 9 0 9 7 0 9 11 11 11 2
18 12 1 0 9 0 9 13 9 9 2 0 9 3 13 7 1 9 2
24 0 13 3 12 9 2 1 9 9 1 11 15 13 11 7 11 2 1 11 3 11 7 11 2
17 0 9 1 11 11 13 1 0 9 11 2 9 13 11 7 11 2
9 2 1 0 9 15 3 13 9 2
16 0 12 9 3 13 1 0 9 2 2 13 15 9 11 11 2
19 13 13 14 9 11 11 2 15 9 1 0 2 7 3 0 0 9 13 2
22 0 9 9 3 3 13 7 1 0 0 9 15 13 13 0 9 2 0 14 1 11 2
25 0 9 11 2 12 2 9 2 12 9 2 12 9 2 12 9 2 9 12 2 12 2 12 9 2
20 13 2 11 2 11 11 2 2 11 2 11 2 2 11 2 9 1 11 2 2
32 13 2 11 2 11 2 2 11 2 12 2 11 11 2 2 11 2 9 1 11 11 2 2 11 2 1 9 9 1 11 2 2
3 9 1 9
2 11 2
19 16 3 15 1 11 13 10 0 9 2 3 13 1 9 1 9 3 12 2
28 1 12 2 12 2 15 13 12 2 9 9 11 7 13 0 9 2 13 4 15 1 15 13 3 16 1 0 2
42 3 15 7 13 1 9 9 1 9 0 11 11 2 15 15 13 1 0 9 13 12 2 12 2 7 13 15 13 1 9 0 9 0 0 11 7 1 9 1 9 11 2
32 10 9 3 13 9 9 11 2 16 10 0 9 1 0 9 13 1 9 2 7 13 15 15 9 1 0 9 1 0 0 9 2
19 1 9 0 9 7 9 9 15 9 9 11 13 10 9 13 1 0 9 2
16 1 9 12 0 9 13 3 0 2 15 1 15 13 0 9 2
5 11 3 1 11 2
2 11 11
15 1 0 0 11 13 9 9 9 0 9 9 11 1 9 2
13 11 11 3 13 1 11 11 9 12 2 12 9 2
11 10 9 11 13 1 9 11 13 3 3 2
15 1 12 9 13 0 9 7 3 1 0 13 9 1 9 2
6 13 3 12 2 12 2
13 1 9 9 9 11 15 4 13 9 11 2 11 2
46 16 15 1 0 0 9 11 1 0 0 9 11 13 2 13 0 9 0 0 9 15 2 9 11 1 11 13 1 9 9 9 11 1 9 11 7 9 13 11 1 9 1 9 9 9 2
8 4 15 13 1 9 1 11 2
10 16 13 9 2 13 15 0 9 9 2
9 11 13 7 1 10 9 0 9 2
10 1 9 11 2 11 13 9 14 0 2
15 9 9 11 1 11 13 9 9 0 9 1 9 9 11 2
16 13 15 3 13 2 16 11 13 11 7 4 13 1 11 3 2
22 13 15 15 13 13 7 11 2 7 3 4 13 13 11 1 0 9 16 9 9 11 2
13 1 15 10 0 9 13 13 0 9 7 0 9 2
30 10 9 9 9 13 15 2 1 1 10 0 0 9 15 11 11 9 9 9 13 1 15 1 9 11 2 11 2 11 2
5 9 1 9 1 9
2 11 2
29 1 0 9 9 9 9 1 0 0 9 2 15 15 13 1 9 1 11 1 11 2 4 13 11 1 12 1 9 2
24 9 11 11 7 11 11 13 1 0 11 7 11 11 15 13 1 9 9 2 15 13 9 11 2
19 0 9 1 10 9 13 11 1 9 12 7 13 1 15 15 12 0 9 2
24 1 11 15 7 11 7 3 11 3 13 2 14 11 1 0 9 13 2 16 13 9 1 9 2
6 9 1 9 13 11 2
10 11 13 11 2 11 13 3 1 15 2
7 11 15 13 11 7 11 2
12 9 11 2 11 2 11 7 11 7 13 0 2
12 1 9 13 1 0 9 11 1 9 1 11 2
3 11 1 11
2 11 2
18 0 9 0 0 0 9 11 11 15 13 0 9 0 0 9 11 11 2
37 11 13 9 1 9 9 12 7 13 1 9 15 9 11 0 2 11 2 15 9 9 11 11 1 9 13 16 0 2 9 2 1 10 0 9 9 2
5 11 13 1 0 9
23 0 9 0 0 9 13 9 11 11 2 15 1 9 13 1 0 9 1 11 9 12 9 2
9 10 9 3 13 1 12 9 3 2
27 2 13 4 2 16 4 15 13 13 7 1 12 2 16 15 0 9 1 9 1 9 13 14 3 1 12 2
26 13 7 3 1 15 0 2 2 13 9 9 11 2 15 13 2 16 15 1 0 9 11 3 13 13 2
31 2 16 13 12 2 13 0 9 2 16 4 13 4 13 1 0 9 1 11 2 2 13 10 9 9 0 0 9 11 11 2
24 11 11 3 1 0 9 13 0 9 2 2 1 12 9 4 3 13 7 13 4 9 1 9 2
14 13 4 12 9 9 2 1 15 4 15 12 9 13 2
21 3 4 15 3 13 0 9 7 16 4 13 1 9 2 3 4 15 13 0 9 2
24 16 3 4 3 1 9 13 13 2 13 0 9 9 2 16 4 1 9 13 3 1 0 9 2
7 3 15 15 7 13 2 2
22 0 0 9 13 3 12 9 2 15 7 1 15 13 2 1 1 0 9 2 14 0 2
4 11 15 13 9
7 1 9 1 11 13 0 11
2 11 2
16 1 3 0 9 13 1 0 11 0 9 9 9 9 0 9 2
30 1 15 9 13 0 9 11 2 9 13 3 9 11 7 9 0 9 1 9 11 11 2 15 13 7 13 9 0 9 2
33 7 1 9 11 7 11 13 9 11 11 2 11 2 1 9 12 9 2 14 0 9 13 10 9 11 7 11 11 1 9 9 11 2
27 0 9 1 9 13 9 9 11 11 1 11 2 1 9 12 9 15 3 13 0 9 11 11 1 0 9 2
17 9 9 0 9 13 0 9 3 12 2 9 11 11 1 0 11 2
4 13 11 11 2
3 0 11 2
15 0 9 0 9 13 11 11 11 9 0 9 1 9 9 2
51 0 0 0 9 11 2 15 13 1 10 9 0 9 11 11 2 13 2 16 15 13 13 1 9 1 0 9 12 2 2 12 2 9 1 11 1 11 0 11 11 2 15 13 1 9 0 9 9 0 9 2
6 0 13 1 9 1 9
12 11 13 11 3 13 2 16 4 13 11 7 11
2 11 2
18 1 0 0 9 2 15 13 9 11 1 11 2 13 0 9 0 9 2
8 11 3 13 1 9 0 11 2
29 9 11 11 13 0 9 2 16 1 0 11 2 11 7 11 13 11 2 0 9 2 7 9 13 7 1 9 11 2
15 2 1 9 15 9 7 3 13 0 2 2 13 15 11 2
21 1 15 2 16 4 13 11 7 11 2 15 13 1 11 2 15 13 14 1 9 2
25 0 13 1 9 1 9 9 1 0 11 1 9 7 11 2 15 13 9 1 9 2 3 1 9 2
20 2 13 4 0 2 16 4 13 0 9 12 2 12 2 2 13 9 11 11 2
8 1 9 15 13 0 12 9 2
12 9 3 9 13 3 13 3 0 11 1 11 2
9 11 4 0 13 1 9 1 11 2
14 0 0 0 9 4 13 13 9 11 11 7 11 11 2
40 2 1 9 13 7 11 2 15 13 3 1 9 3 0 9 2 7 3 3 15 13 1 9 10 9 7 13 1 9 2 2 13 15 9 2 9 2 11 11 2
19 3 7 13 2 16 1 0 9 1 0 9 1 11 13 9 1 9 11 2
12 1 0 11 13 9 0 9 1 3 0 11 2
19 0 9 2 0 1 11 2 11 7 0 9 11 7 11 2 7 13 13 2
9 11 4 0 11 13 0 0 9 2
7 0 9 13 11 1 11 2
26 11 3 13 1 9 11 2 0 7 11 2 15 13 1 0 9 2 2 11 7 11 2 12 0 2 2
10 1 9 3 13 14 12 9 2 2 2
25 1 0 9 15 13 2 3 15 11 11 2 15 15 1 0 9 13 1 9 2 13 1 11 11 2
18 2 13 2 16 15 13 0 9 2 2 13 9 2 9 2 11 11 2
19 11 1 9 13 11 12 9 7 0 9 13 10 9 7 1 0 0 9 2
29 1 9 15 3 3 13 11 2 7 16 3 11 2 15 15 1 9 13 9 1 11 2 13 3 0 7 13 13 2
11 9 12 2 9 2 15 1 12 9 2 2
8 13 15 9 2 9 2 11 11
27 11 11 2 9 0 9 7 9 11 2 15 0 9 13 9 2 1 15 15 13 4 13 1 9 9 9 2
31 0 0 9 13 0 9 11 0 11 9 9 1 12 2 9 0 9 7 9 12 9 1 9 1 9 1 9 12 2 9 2
4 11 13 10 11
7 0 0 9 1 3 12 9
2 11 2
13 1 0 9 3 12 12 9 13 0 9 0 9 2
20 0 9 11 13 1 11 10 0 9 7 13 15 12 9 1 9 12 2 12 2
6 11 11 12 11 11 12
12 13 15 1 0 9 2 15 13 7 0 9 2
8 1 9 7 13 14 1 9 2
22 3 0 9 11 13 9 1 0 9 7 11 7 1 9 1 12 2 9 3 13 11 2
28 3 3 13 11 1 12 2 9 2 11 13 1 0 9 11 2 3 1 9 3 13 7 11 13 1 9 13 2
16 11 13 1 0 9 7 0 9 2 7 12 15 15 7 13 2
20 14 1 12 2 9 11 13 11 7 11 7 11 13 1 9 1 15 14 9 2
4 13 10 9 2
9 16 9 1 0 9 13 9 0 2
32 3 13 11 2 11 15 13 1 0 9 7 1 9 3 11 9 13 2 3 11 13 0 9 9 11 7 11 13 12 2 12 2
20 3 15 13 13 9 2 1 12 9 11 13 1 12 2 12 7 0 3 13 2
21 1 12 2 9 13 11 0 9 14 9 9 2 7 0 9 13 11 1 0 9 2
8 9 0 11 15 1 0 9 13
2 11 2
9 2 11 13 0 9 1 0 9 2
22 7 15 3 13 9 9 7 9 15 3 13 2 2 13 1 9 1 11 9 11 11 2
23 3 3 16 9 1 9 13 0 9 9 2 16 9 4 13 13 9 10 9 1 0 9 2
28 15 7 13 13 9 2 15 15 13 1 9 9 12 9 1 9 7 15 4 13 0 9 2 13 1 9 2 2
11 9 9 2 9 7 9 13 9 1 9 2
26 2 9 13 0 2 16 4 1 9 13 7 3 10 9 2 13 4 15 0 2 2 13 9 11 11 2
33 1 0 9 7 10 9 1 11 2 3 3 12 9 13 2 13 0 2 2 3 4 15 15 13 13 2 16 13 9 1 9 9 2
19 13 4 15 3 13 7 15 2 16 4 1 9 13 12 14 0 9 2 2
10 12 1 9 13 1 9 9 9 11 2
14 1 9 0 9 15 13 12 9 11 1 9 12 9 2
36 2 1 0 9 13 9 13 2 2 13 1 0 9 9 11 2 7 11 1 10 9 1 12 2 12 13 9 11 2 2 11 15 3 13 2 2
20 0 9 15 13 2 2 10 9 4 3 13 2 13 2 3 15 13 9 2 2
28 1 9 15 1 9 11 3 13 2 9 2 16 4 15 13 9 2 13 1 15 2 16 15 13 0 9 9 2
38 9 11 13 9 2 2 13 15 0 9 1 0 0 9 7 1 0 9 1 15 2 2 13 1 15 7 13 2 16 3 3 11 13 16 13 1 9 2
30 9 11 11 3 3 13 2 16 10 9 13 1 10 9 3 1 9 3 2 2 3 2 16 4 13 9 13 3 3 2
11 11 2 11 7 0 15 13 10 9 2 2
1 3
34 0 9 0 3 9 13 3 13 0 9 1 0 9 9 2 12 1 11 2 3 13 3 7 3 1 9 9 9 12 1 9 1 9 2
5 9 9 11 13 0
4 11 2 11 2
19 0 9 0 0 9 15 9 11 11 15 13 1 9 12 2 9 1 9 2
23 0 0 9 2 15 13 9 9 2 13 1 9 13 3 11 11 2 11 11 7 11 11 2
38 2 1 9 7 0 9 13 15 0 2 3 4 15 13 11 11 2 9 11 2 9 2 9 2 2 2 13 3 11 11 11 2 11 2 9 0 11 2
28 11 0 9 11 2 9 7 9 0 0 9 11 2 1 9 13 1 11 2 3 1 0 9 13 1 0 11 2
5 3 1 9 11 11
17 1 9 9 1 9 11 15 13 0 9 9 11 7 9 0 11 11
23 1 9 11 11 2 0 9 9 0 9 1 9 0 11 2 4 3 16 0 9 3 13 2
22 11 4 1 9 12 1 11 3 13 0 9 7 13 1 0 9 1 0 11 1 11 2
25 3 13 9 11 7 13 15 2 1 9 9 0 0 9 7 3 16 2 0 9 2 2 10 9 2
35 16 0 9 1 10 9 15 13 1 3 0 2 0 9 3 13 2 13 0 9 11 2 11 2 11 2 15 13 1 15 9 0 9 2 2
62 10 9 7 9 1 9 9 1 9 0 9 2 11 12 2 12 2 12 2 0 9 13 3 2 12 0 9 12 9 0 9 2 0 9 9 11 11 7 9 9 0 11 2 15 4 1 9 12 13 1 9 13 9 0 0 9 7 9 2 11 11 2
5 13 9 13 3 11
25 1 9 9 12 2 3 1 9 9 9 13 11 11 2 15 3 11 13 2 3 2 13 0 9 2
34 1 0 9 1 9 7 11 11 13 3 7 10 9 4 13 14 1 9 12 2 1 9 2 3 15 9 9 11 1 10 0 9 13 2
30 15 15 15 3 13 1 0 9 9 7 9 0 0 9 2 1 12 9 1 9 4 13 7 0 12 9 13 1 9 2
11 1 9 15 3 1 9 1 0 9 13 2
22 2 1 0 9 15 13 14 3 2 13 15 10 0 9 2 2 13 3 0 11 11 2
29 2 9 13 7 1 15 0 15 2 16 15 13 10 9 2 15 4 13 1 10 9 1 11 1 9 12 7 12 2
29 1 11 15 13 0 9 9 0 9 11 11 2 15 15 1 9 13 9 0 9 2 3 15 13 1 9 9 2 2
16 15 13 9 9 9 1 11 1 9 12 7 10 15 13 9 2
9 1 10 9 4 3 3 13 9 2
13 11 13 9 1 0 11 2 13 1 9 0 9 2
9 9 9 0 4 13 3 0 9 2
25 13 1 15 9 9 9 0 11 2 15 16 9 2 10 10 9 3 4 3 13 2 9 16 9 2
20 9 9 1 11 7 13 1 10 0 9 2 16 13 10 9 3 0 7 0 2
19 13 4 15 2 16 15 15 11 13 2 16 15 9 13 10 9 2 2 2
11 13 15 2 16 11 13 1 9 0 9 2
16 15 1 15 13 2 13 15 7 3 1 0 9 11 1 15 2
10 15 9 1 11 4 7 13 1 9 2
10 0 9 1 11 13 9 11 2 11 2
28 1 0 9 13 2 16 11 3 9 9 2 13 2 1 9 11 0 9 2 15 3 4 0 3 13 2 2 2
14 13 1 15 3 14 1 9 7 1 0 9 15 0 2
21 1 10 9 2 3 1 9 12 7 12 2 4 13 1 11 1 11 7 1 11 2
15 13 7 13 2 16 11 2 11 4 3 13 1 10 9 2
21 1 9 9 13 0 2 0 9 3 13 3 0 2 13 15 9 9 0 14 9 2
10 13 4 15 15 13 7 3 2 2 2
18 16 15 13 9 1 9 2 3 13 13 1 0 9 11 1 9 12 2
15 13 4 1 0 9 2 11 2 0 9 2 9 0 9 2
11 3 4 15 13 7 3 7 13 1 9 2
12 9 9 9 11 1 11 13 3 9 10 9 2
22 3 4 4 1 3 9 13 1 9 9 0 9 1 11 2 3 15 13 9 7 9 2
11 1 9 11 2 9 11 2 4 13 11 2
20 0 9 1 11 15 3 13 10 0 9 1 0 9 11 2 0 9 7 9 2
12 1 9 12 3 0 11 13 1 11 2 2 2
21 15 15 13 2 15 1 10 9 13 3 10 0 9 3 0 9 2 3 1 11 2
7 11 13 14 9 2 2 2
3 9 1 11
26 9 9 0 11 11 11 2 0 3 1 11 1 11 2 13 1 10 9 1 0 9 13 1 0 9 2
14 1 0 9 11 3 13 14 12 9 9 9 1 9 2
37 11 13 2 16 1 10 9 13 3 1 9 9 2 15 4 2 14 3 2 13 9 1 11 2 3 15 11 13 3 1 0 0 9 1 9 2 2
18 1 9 2 15 4 1 9 13 3 9 11 2 13 3 7 11 11 2
30 2 1 9 12 14 1 0 9 4 4 13 16 9 0 9 1 0 9 0 2 9 3 0 2 2 13 11 2 11 2
19 2 13 4 12 1 10 9 9 1 0 9 2 15 4 13 13 1 9 2
60 1 0 0 9 13 9 1 11 15 1 9 9 1 11 13 11 11 2 9 0 9 7 9 0 15 9 1 3 0 9 2 7 13 15 2 16 4 13 1 9 1 12 2 1 12 2 9 12 7 16 15 13 11 11 2 3 9 0 9 2
5 3 15 3 13 2
19 2 11 3 13 0 0 9 2 15 3 11 13 13 2 9 2 9 2 2
36 10 0 0 9 4 13 13 3 1 9 12 3 1 11 11 2 16 4 15 13 1 0 9 1 11 2 3 9 1 9 9 2 11 1 9 2
15 3 4 0 9 0 9 13 1 0 0 9 0 1 9 2
20 13 9 2 16 13 11 2 16 2 9 2 9 13 2 9 13 1 12 9 2
42 13 0 9 2 16 4 10 9 13 1 11 2 9 9 1 0 9 9 2 2 3 13 11 2 7 16 4 11 13 1 0 9 10 9 9 2 2 13 11 2 11 2
4 3 14 9 2
24 13 4 3 0 2 16 4 15 0 9 13 13 9 1 0 0 9 2 0 9 7 0 9 2
27 10 10 0 7 0 9 13 1 10 9 0 9 11 11 7 11 2 15 1 10 9 13 14 1 0 9 2
13 9 11 11 1 15 10 0 9 13 12 1 15 2
24 15 2 15 11 1 10 9 3 13 2 13 13 0 0 9 2 3 9 7 0 9 0 9 2
11 3 4 15 13 1 9 13 3 0 9 2
20 0 9 3 13 9 0 9 7 10 0 7 3 0 9 1 9 9 1 11 2
14 13 9 9 9 2 15 9 13 1 9 9 1 11 2
11 13 2 16 15 13 3 14 9 2 2 2
18 9 1 9 1 11 2 0 7 0 0 0 9 2 13 9 0 9 2
20 1 9 13 3 1 9 9 2 3 7 13 9 9 11 2 11 11 2 2 2
4 2 9 3 2
16 0 9 4 3 13 1 10 0 9 9 2 0 3 15 13 2
18 0 9 9 9 13 11 11 2 0 9 0 9 3 1 9 0 9 2
4 2 9 3 2
6 0 9 1 15 9 13
11 0 9 1 0 9 13 9 11 9 9 2
15 9 9 13 13 1 0 9 7 13 1 15 3 0 9 2
19 15 2 15 13 15 3 2 13 15 3 13 15 1 15 7 1 10 9 2
7 0 9 9 9 13 9 2
20 0 2 0 2 3 15 0 9 2 1 0 9 15 3 0 1 0 0 9 2
12 9 13 3 9 2 16 9 9 11 13 9 2
27 13 15 16 9 2 13 0 9 9 9 7 3 13 7 1 9 1 9 2 16 4 15 13 9 7 3 2
16 9 11 15 16 9 13 2 13 15 9 7 3 13 13 9 2
40 1 0 9 7 1 15 2 16 9 2 9 13 13 1 9 0 9 2 4 15 1 0 13 1 9 2 11 11 1 0 9 12 2 0 9 9 0 1 11 2
12 9 9 2 13 13 9 1 0 9 7 9 2
15 9 15 13 0 9 2 3 15 2 10 9 9 3 13 2
17 1 9 2 9 2 13 0 9 7 15 2 3 9 13 15 15 2
24 0 9 16 1 9 13 1 9 2 9 7 9 2 1 9 13 1 0 15 2 1 0 9 2
9 13 0 0 9 9 1 10 9 2
14 1 15 10 9 13 2 0 13 0 9 1 0 9 2
25 0 9 9 2 15 4 3 13 2 13 1 0 9 1 11 2 12 9 13 3 1 12 12 9 2
18 13 15 3 0 9 2 15 13 1 15 2 16 9 13 3 0 9 2
23 9 9 1 0 9 3 13 3 0 2 7 9 15 1 15 3 13 7 13 14 12 9 2
28 13 7 13 2 16 13 3 3 9 2 15 0 9 13 7 15 15 13 1 15 2 16 1 9 9 4 13 2
12 1 10 9 15 13 9 13 0 9 13 9 2
21 16 13 1 0 9 2 13 15 9 13 2 16 4 16 0 13 1 10 0 9 2
39 3 3 2 3 15 9 13 13 2 9 9 13 2 16 0 0 9 1 10 9 13 1 10 9 1 9 0 9 16 0 9 0 1 9 1 0 0 9 2
14 10 9 13 9 9 9 7 3 1 15 13 3 13 2
25 0 9 9 0 9 13 0 9 2 0 9 2 0 9 7 3 7 0 9 9 1 9 1 9 2
24 1 9 9 13 13 9 0 12 9 2 16 13 0 2 16 4 13 3 0 0 7 0 9 2
29 12 1 0 9 2 3 1 3 0 9 2 13 2 16 4 1 9 13 3 12 1 9 2 3 3 15 1 9 2
15 1 9 1 0 9 15 1 0 13 0 9 1 9 9 2
10 10 9 13 1 0 9 0 0 9 2
13 0 13 2 16 4 9 1 0 9 4 3 13 2
10 1 0 9 13 9 9 9 3 0 2
21 16 15 13 0 9 2 13 1 0 9 10 0 9 2 15 3 3 13 0 9 2
6 3 13 9 0 9 2
18 13 0 9 9 2 15 1 9 9 13 1 9 2 3 13 0 9 2
7 9 11 13 1 0 9 2
11 15 1 10 9 13 1 0 9 9 0 2
22 9 9 13 1 9 9 1 9 2 3 13 3 2 7 13 15 1 0 9 10 9 2
14 16 15 9 13 2 13 4 13 1 9 1 15 15 2
10 13 15 3 1 9 0 9 3 13 2
18 3 15 1 15 0 1 9 13 2 7 3 15 1 0 9 9 13 2
12 9 15 13 2 16 15 1 15 9 13 13 2
12 1 9 9 3 13 9 2 16 15 15 13 2
17 1 10 9 13 9 9 0 7 10 9 13 13 0 9 1 9 2
9 0 7 0 9 13 3 1 9 2
14 13 0 9 15 13 2 16 4 9 13 10 9 13 2
35 13 9 9 2 15 15 13 9 1 9 2 7 15 15 13 1 9 16 9 2 13 16 9 1 9 2 16 1 15 3 10 9 4 13 2
17 1 9 9 9 4 13 13 2 16 3 9 3 13 1 0 9 2
12 0 9 3 13 3 9 16 0 9 0 9 2
11 10 9 13 13 9 7 0 9 1 9 2
12 9 9 15 13 2 16 13 13 9 1 9 2
22 13 15 2 16 4 15 15 13 9 14 3 2 16 13 9 1 9 7 15 13 9 2
22 3 0 9 9 15 10 9 13 2 16 13 1 0 9 2 7 13 13 9 1 9 2
32 1 15 15 3 3 13 9 0 7 0 2 3 15 13 1 9 9 13 2 16 10 9 13 0 13 1 0 9 1 0 9 2
45 16 1 15 15 13 2 16 13 0 9 2 7 13 1 15 0 3 13 2 13 15 1 10 9 2 7 13 1 9 2 13 15 3 9 7 9 13 2 1 10 9 4 15 13 2
5 7 9 15 13 2
4 11 13 0 9
2 11 2
24 0 9 9 11 11 3 13 3 0 0 0 0 9 2 11 2 7 13 9 1 10 0 9 2
19 9 3 13 9 1 12 9 9 7 9 11 1 0 11 7 13 10 9 2
17 11 15 13 9 0 9 11 2 13 0 0 9 7 13 1 9 2
22 1 9 9 11 11 11 1 0 9 10 9 13 9 11 2 13 15 9 2 1 11 2
13 0 2 9 2 13 13 1 9 9 2 13 2 2
15 0 9 9 3 3 13 3 0 9 0 9 2 11 2 2
22 1 9 12 2 9 13 1 11 13 7 13 3 12 3 3 0 7 0 9 7 9 2
15 11 2 0 9 7 9 13 9 0 2 15 13 1 0 9
5 11 13 9 1 9
6 11 2 11 2 11 2
28 0 9 3 13 12 9 7 12 0 0 9 7 12 9 13 1 9 1 9 11 7 11 1 0 0 9 11 2
7 13 15 0 7 0 9 2
26 9 13 12 11 1 0 9 2 1 15 9 1 11 13 1 9 9 7 15 13 0 9 7 9 13 2
14 1 0 9 1 10 9 0 9 1 9 13 12 11 2
26 1 11 2 3 1 9 0 9 13 12 0 9 2 9 13 1 9 12 0 0 9 7 12 0 9 2
30 1 11 9 1 9 13 9 13 1 0 0 9 2 15 13 9 1 9 7 9 7 15 15 3 1 9 13 9 9 2
16 1 9 15 3 1 0 9 0 0 9 9 13 1 12 11 2
7 9 3 9 1 9 13 2
24 1 1 0 9 9 1 11 7 1 0 9 0 0 9 3 0 9 1 11 3 13 0 9 2
27 1 0 9 13 1 9 12 9 7 10 9 4 13 7 1 9 2 1 15 1 0 9 13 0 0 9 2
22 0 0 9 11 3 13 11 0 9 1 0 9 2 16 11 13 13 9 1 0 11 2
50 1 9 9 11 0 9 11 11 11 1 9 9 9 1 11 13 2 16 2 0 9 9 13 3 9 13 1 0 9 1 0 11 2 4 2 14 10 9 13 7 13 7 4 2 14 13 10 9 2 2
29 1 11 1 9 11 1 9 0 9 7 1 9 9 9 13 9 2 16 4 11 3 1 0 11 13 0 0 9 2
24 0 9 0 9 1 0 11 11 11 7 3 13 2 16 15 11 13 0 9 13 1 0 9 2
5 11 2 9 9 9
2 11 2
13 0 9 11 11 13 13 9 0 9 1 9 9 2
14 13 15 1 11 1 0 0 9 1 9 9 9 9 2
14 9 15 13 9 2 9 2 0 9 7 0 9 9 2
26 1 11 14 4 10 9 13 7 14 3 9 0 9 2 16 3 2 0 9 0 9 9 1 9 2 2
27 9 11 13 2 16 9 13 1 9 9 0 9 13 1 0 9 2 15 4 1 11 13 0 9 1 11 2
40 11 3 13 2 16 13 9 1 3 0 0 9 11 2 13 2 16 13 1 0 9 0 9 2 7 13 2 16 13 2 0 9 1 9 0 0 9 11 2 2
20 3 13 2 16 1 9 1 0 9 2 10 0 9 4 13 1 9 11 2 2
4 9 13 11 9
2 11 2
49 9 1 11 11 7 9 0 9 3 1 0 11 13 0 9 3 2 16 0 9 13 12 9 9 1 9 2 15 15 13 15 2 16 13 9 9 1 9 0 11 1 11 9 0 15 1 9 11 2
41 16 13 9 11 2 9 1 0 0 9 11 11 13 0 9 7 9 1 0 0 2 15 13 2 9 0 9 2 2 2 13 9 1 9 2 7 2 9 11 2 2
19 9 9 9 13 0 9 1 9 0 9 7 13 15 1 2 9 9 2 2
14 9 3 13 1 9 9 1 9 2 16 4 13 9 2
5 0 9 1 9 9
14 0 0 0 9 0 11 13 0 9 1 9 1 12 9
15 16 0 11 4 1 10 9 13 9 2 1 15 15 13 2
13 1 9 3 13 0 9 2 9 0 2 0 9 2
15 0 9 7 13 3 1 10 0 9 9 1 3 0 9 2
29 0 0 2 9 2 1 0 9 15 3 3 13 1 9 2 1 9 13 0 0 9 11 2 0 2 0 0 11 2
14 3 1 12 9 15 13 2 16 9 10 9 13 9 2
12 10 2 9 2 9 15 13 2 7 16 13 2
24 1 9 0 9 15 3 15 13 13 2 16 15 0 9 13 1 10 2 9 2 16 9 12 2
8 3 13 9 9 1 12 9 2
14 3 15 13 13 0 2 9 2 7 13 12 9 3 2
27 9 13 2 16 9 9 7 9 0 9 1 12 9 2 15 3 13 1 9 2 3 13 0 9 10 9 2
12 11 13 2 16 9 9 4 13 12 9 9 2
15 2 10 9 13 3 9 7 0 9 2 2 13 0 9 2
13 3 3 13 14 9 12 7 12 9 9 0 11 2
17 1 9 7 9 13 1 12 0 9 1 9 1 9 12 12 9 2
10 3 13 13 12 12 9 1 12 9 2
17 1 12 2 9 2 3 13 0 9 9 2 15 9 0 13 13 2
8 1 9 9 9 3 13 9 2
8 13 7 9 2 0 11 13 2
12 13 15 9 1 0 7 0 9 1 9 12 2
7 3 13 9 2 9 2 2
10 1 11 13 0 9 3 1 9 12 2
12 1 12 9 9 13 7 0 9 1 0 9 2
11 3 12 0 9 9 13 2 16 9 13 2
14 13 15 3 2 16 9 2 0 9 2 4 3 13 2
28 2 15 3 13 2 16 4 9 13 1 9 12 9 7 9 1 15 13 1 9 2 2 13 10 9 11 11 2
12 9 13 9 9 7 9 1 12 1 0 9 2
8 1 0 9 4 13 3 9 2
30 14 15 13 1 9 2 10 9 9 1 9 9 2 7 13 10 0 9 2 13 15 0 9 9 11 11 2 11 2 2
20 2 9 9 3 3 13 2 2 13 0 9 9 0 9 1 0 9 11 11 2
17 9 13 2 16 13 3 1 9 1 9 9 2 13 7 0 9 2
15 13 1 11 2 9 9 1 9 2 13 7 9 0 9 2
15 15 3 4 13 9 0 11 2 15 0 13 9 12 9 2
8 7 15 0 13 7 0 9 2
11 0 9 9 13 13 0 2 0 9 2 2
13 9 2 9 2 3 13 0 9 1 3 0 9 2
23 16 9 13 9 2 16 1 9 13 7 3 0 9 1 0 9 13 0 16 0 9 9 2
7 3 13 1 9 0 11 2
33 1 9 0 2 0 9 13 0 9 9 11 2 0 9 9 15 13 9 9 0 9 2 1 15 13 1 11 14 9 9 9 9 2
7 0 9 3 13 0 9 11
4 11 2 11 2
18 9 0 9 7 0 9 9 15 13 1 9 1 9 1 0 9 11 2
20 1 9 15 0 9 9 0 9 13 3 1 9 13 0 9 1 0 0 9 2
32 0 9 13 2 16 0 9 0 9 0 1 9 9 11 2 0 12 9 1 11 2 3 12 9 13 9 9 1 9 0 9 2
22 9 4 13 3 1 9 11 7 11 2 3 15 13 9 0 9 2 3 16 13 11 2
20 1 10 9 0 9 1 9 0 9 3 3 10 9 13 7 4 13 3 13 2
16 11 11 13 9 2 15 13 9 0 9 1 11 1 0 9 2
20 1 9 11 13 9 9 13 0 0 9 1 0 9 10 0 9 1 0 9 2
29 0 9 0 9 13 2 16 10 9 4 13 13 9 0 9 1 0 9 7 13 10 9 14 1 9 0 0 9 2
45 0 9 11 11 3 13 9 2 16 11 3 13 0 9 11 11 2 7 13 2 16 0 9 13 1 0 9 11 2 13 13 9 1 0 0 9 7 3 13 11 9 1 9 11 2
31 9 11 9 3 13 9 9 11 2 11 1 0 0 9 9 11 11 2 15 14 1 0 13 2 16 11 13 11 12 9 2
25 9 9 9 7 9 1 9 13 9 11 1 11 11 1 11 2 15 3 4 13 1 12 2 9 2
1 3
23 9 0 9 9 11 11 1 0 9 11 13 0 0 9 1 9 10 9 13 1 0 9 2
34 3 15 7 13 2 16 1 0 9 13 0 13 7 0 9 1 9 9 1 11 2 9 0 9 1 0 9 7 9 9 1 0 9 2
19 0 9 13 1 0 9 9 12 9 3 0 9 1 9 12 9 0 9 2
20 9 0 12 9 0 9 13 1 9 1 0 11 1 12 0 0 9 1 11 2
10 9 15 1 9 13 13 12 0 9 2
16 1 0 9 4 9 13 7 11 2 15 13 0 9 9 9 2
21 9 0 9 2 15 1 9 3 13 0 9 1 0 9 2 15 1 0 9 13 2
27 9 0 9 0 0 9 0 0 9 1 9 15 3 13 13 10 9 1 9 1 11 7 0 0 9 13 2
15 9 1 9 13 1 9 1 9 0 9 1 0 0 9 2
20 9 4 13 1 12 9 3 1 0 9 1 9 9 0 2 11 1 0 9 2
30 16 3 13 0 9 0 2 11 2 12 9 13 0 9 2 15 15 13 13 0 9 1 9 9 1 9 11 2 11 2
14 0 15 15 13 3 0 9 2 15 15 13 1 9 2
28 9 0 9 0 9 11 13 1 9 1 11 1 9 1 11 0 0 9 1 11 9 0 9 0 9 11 11 2
26 13 2 16 2 9 2 16 13 0 9 1 11 2 4 13 13 2 0 9 2 9 9 1 11 2 2
4 9 11 15 13
30 9 0 2 0 2 0 7 15 0 9 13 7 9 2 0 0 9 2 2 0 3 13 2 15 13 1 9 0 7 3
20 9 9 2 9 7 9 13 9 2 1 15 13 1 9 0 9 0 0 9 2
14 9 4 13 4 13 3 3 1 9 1 0 9 9 2
9 0 9 9 13 9 9 9 9 2
33 2 0 0 9 2 2 3 3 11 9 13 2 13 1 9 0 0 9 7 9 9 3 2 1 9 7 9 14 1 9 7 9 2
15 13 1 9 3 0 2 15 15 1 0 0 9 3 13 2
14 16 13 1 9 0 2 9 4 13 1 0 9 9 2
14 10 0 2 3 2 14 0 9 7 0 9 3 13 2
22 13 3 3 0 9 1 0 9 2 0 9 9 7 0 0 9 9 1 15 9 9 2
31 9 0 2 0 2 0 7 15 0 9 13 7 9 2 0 0 9 2 2 0 3 13 2 15 13 1 9 0 7 3 2
23 9 0 9 0 9 0 9 15 3 3 13 1 9 10 0 9 2 15 3 13 0 9 2
8 0 9 9 13 3 0 9 2
25 9 1 9 0 2 0 9 2 0 1 0 9 2 3 0 9 9 2 13 1 9 0 9 11 2
17 15 7 2 3 16 1 0 9 2 13 1 0 9 1 0 11 2
29 10 9 2 1 15 0 9 13 2 3 0 9 1 0 9 9 7 0 9 1 9 0 9 2 13 3 0 9 2
8 3 3 13 1 9 0 9 2
6 13 14 1 9 9 2
20 1 0 9 7 13 9 1 0 9 1 9 9 7 0 9 0 9 0 9 2
24 1 0 9 2 3 1 9 0 9 3 13 9 9 1 9 2 13 9 0 0 9 3 9 2
10 3 13 0 13 7 9 1 0 9 2
31 0 0 0 9 2 3 0 0 9 7 0 9 13 9 1 9 1 11 13 1 0 9 1 9 7 1 9 0 0 9 2
17 0 0 9 7 1 9 9 13 3 9 2 0 9 13 9 9 2
11 0 9 13 4 13 3 1 3 0 9 2
19 9 10 9 13 2 16 1 2 0 9 2 9 1 9 0 9 3 13 2
14 0 9 10 9 2 9 2 1 9 13 0 7 9 2
19 0 9 13 3 9 2 3 14 9 1 0 9 13 11 1 9 11 13 2
24 3 16 9 1 11 13 15 0 9 1 9 9 1 9 1 9 1 2 9 9 0 9 2 2
26 0 9 13 3 13 0 9 0 9 7 9 2 14 3 1 9 9 2 0 9 7 0 3 0 9 2
8 10 9 15 13 16 3 0 2
16 3 9 13 9 9 1 9 9 1 0 9 1 9 0 9 2
10 1 0 4 15 14 13 0 0 9 2
27 9 7 13 2 3 4 15 1 10 9 2 9 2 9 0 9 13 1 10 3 0 0 9 7 0 9 2
32 9 13 10 0 9 1 9 9 11 2 15 3 3 13 9 9 0 9 1 10 9 2 9 1 0 9 7 0 9 14 13 2
12 7 1 3 0 9 13 9 9 11 0 9 2
25 1 15 2 16 4 15 11 13 0 0 9 0 9 2 7 3 13 3 10 0 9 7 0 9 2
3 9 12 9
21 1 0 9 15 1 15 0 3 13 0 9 7 9 0 9 13 13 2 1 9 2
6 3 13 13 3 15 2
30 1 0 9 2 9 7 9 2 3 3 2 13 13 2 16 1 10 9 13 3 15 2 15 4 13 2 1 0 9 2
49 9 0 9 2 0 9 0 9 7 1 0 9 9 0 9 3 2 16 15 9 1 10 9 13 9 2 13 10 0 9 7 9 1 9 3 0 9 1 0 7 0 9 1 15 2 15 15 13 2
5 3 1 0 9 2
29 9 3 4 13 10 2 7 13 15 3 9 0 2 16 13 16 0 9 13 7 13 9 2 15 4 15 13 13 2
24 13 2 14 10 9 10 9 9 1 15 2 13 0 15 13 15 2 16 10 9 4 3 13 2
32 9 2 9 2 9 2 16 3 9 3 0 2 15 3 13 13 9 13 9 0 9 7 13 2 16 4 9 4 15 15 13 2
19 3 15 3 13 3 9 2 15 10 9 1 15 13 7 1 15 3 13 2
26 1 9 7 3 12 9 9 7 9 13 13 9 9 2 13 9 9 2 13 9 7 2 3 2 13 2
9 15 15 3 15 1 10 9 13 2
13 7 9 13 2 9 13 2 0 9 13 1 9 2
46 0 0 9 2 0 9 2 13 3 0 9 13 10 0 9 2 15 3 3 7 3 13 1 10 2 0 2 9 2 15 15 16 4 3 7 13 0 2 2 16 9 13 1 9 12 2
12 13 1 9 2 16 7 10 9 13 0 13 2
25 13 2 14 7 9 15 2 16 9 9 7 3 7 0 9 4 13 0 9 2 13 15 15 13 2
23 13 9 9 0 9 7 9 2 13 9 0 9 2 13 13 2 3 10 9 0 9 13 2
35 0 7 0 9 1 10 9 13 15 2 15 15 13 1 0 0 9 2 3 15 13 7 13 9 7 15 0 15 13 1 9 1 0 9 2
24 9 1 9 2 0 9 2 0 16 0 9 2 7 15 2 16 1 0 15 9 15 13 9 2
16 0 9 2 0 1 9 1 9 9 2 0 9 7 0 9 2
9 0 9 2 9 2 9 7 9 2
2 9 2
12 9 2 3 7 9 7 0 9 1 0 9 2
6 3 0 9 0 9 2
16 9 2 9 2 9 0 9 7 3 9 1 9 0 15 9 2
3 0 2 2
6 9 7 13 0 9 2
7 9 13 9 1 0 9 2
5 9 1 9 0 2
13 7 9 13 2 9 13 2 0 9 13 1 9 2
24 0 0 9 2 13 15 9 7 9 2 2 15 3 13 9 2 0 0 9 2 2 13 3 2
22 1 9 16 1 0 9 13 0 2 0 2 3 0 2 0 2 0 2 2 9 2 2
21 13 15 9 7 10 9 13 9 2 9 2 9 2 9 2 9 7 9 1 15 2
9 13 15 7 1 15 15 13 13 2
5 13 13 3 15 2
21 1 0 9 15 1 15 0 3 13 0 9 7 9 0 9 13 13 2 1 9 2
6 3 13 13 3 15 2
14 0 9 9 12 2 2 16 4 13 3 2 13 9 2
17 9 15 13 13 2 16 13 0 7 3 0 9 7 9 15 13 2
10 1 9 3 13 2 16 9 13 2 2
16 13 0 9 2 9 4 13 1 9 2 7 1 12 9 3 2
19 9 9 10 9 1 9 0 9 13 13 15 2 16 3 13 13 3 15 2
19 3 13 15 13 1 9 2 9 15 13 7 15 13 2 0 2 10 9 2
6 10 9 3 13 0 2
27 0 9 2 0 1 9 2 15 15 13 2 15 10 0 9 3 13 2 7 1 15 13 0 9 0 9 2
4 15 3 13 2
8 9 13 3 10 9 7 9 2
15 0 9 2 9 0 9 2 15 3 13 9 0 9 9 2
17 13 2 14 15 3 3 2 13 0 9 13 3 9 9 0 9 2
6 9 0 9 1 9 2
2 0 9
23 0 9 0 9 11 11 1 0 9 9 0 9 13 2 16 9 9 13 1 11 13 9 2
18 3 16 2 0 9 2 13 7 9 9 10 9 13 2 0 9 2 2
10 9 10 0 9 13 11 1 0 9 2
16 2 0 2 9 9 11 14 13 0 9 7 1 15 7 9 2
33 1 10 9 3 13 0 9 2 16 15 3 9 4 13 9 9 11 2 15 3 4 10 9 13 13 1 9 2 1 15 15 13 2
18 3 9 9 1 0 7 0 9 1 9 9 1 9 14 13 0 9 2
22 7 11 13 1 9 0 0 9 7 13 0 9 2 10 9 4 13 13 0 9 11 2
37 13 15 2 16 11 13 0 9 0 0 9 1 0 9 2 13 2 16 9 3 15 13 9 2 7 15 2 16 15 4 13 0 9 0 0 9 2
25 13 3 2 16 9 11 1 0 9 1 11 3 13 9 2 7 16 1 9 4 15 9 13 9 2
17 0 13 9 2 16 9 0 9 0 9 13 15 13 9 10 9 2
19 11 3 0 9 13 15 2 16 9 9 11 13 0 2 16 4 13 9 2
24 13 15 2 16 4 13 15 1 9 1 9 7 15 4 15 13 9 1 12 7 13 15 9 2
19 13 4 15 15 2 16 13 9 0 7 0 2 16 4 15 13 1 9 2
5 3 3 0 9 2
9 9 13 3 9 7 9 1 9 2
16 7 9 0 9 11 13 13 3 3 1 9 16 1 9 12 2
21 13 9 2 16 9 13 11 0 9 9 2 1 15 4 13 0 9 0 0 9 2
23 9 9 2 15 15 9 13 2 13 13 9 2 15 9 9 9 9 1 9 9 11 13 2
6 9 13 3 9 9 2
32 13 3 0 1 0 9 13 15 9 10 7 15 9 2 16 3 15 1 0 9 13 2 15 15 4 15 3 13 0 9 13 2
20 7 15 2 15 4 13 1 9 2 13 3 16 9 2 10 9 15 13 13 2
26 9 13 7 0 13 14 3 2 13 2 14 15 9 2 7 9 0 1 0 9 15 13 15 13 9 2
9 10 9 15 13 1 15 0 9 2
25 14 1 11 2 7 7 1 9 2 9 7 0 9 13 13 9 1 9 0 9 7 0 9 9 2
14 10 9 15 3 13 2 16 3 1 9 13 15 0 2
7 3 15 15 13 7 11 2
18 10 1 0 9 0 9 15 7 13 0 9 2 9 2 9 2 9 2
4 9 1 0 9
25 1 9 0 0 9 3 0 9 1 0 9 7 9 13 9 1 9 9 9 1 0 9 7 9 2
32 13 3 13 2 16 0 9 13 0 2 16 3 0 3 12 9 1 12 3 0 7 3 0 9 2 7 3 15 14 15 13 2
18 0 9 3 13 9 2 0 2 9 1 0 9 7 3 1 15 13 2
5 0 9 13 0 2
23 7 15 9 3 3 13 9 2 16 4 0 9 1 0 9 13 12 9 9 1 0 9 2
9 14 13 2 16 3 10 9 13 2
26 3 15 3 15 13 13 2 1 15 4 13 13 2 16 4 1 15 1 12 9 13 3 9 9 9 2
16 4 15 3 13 13 9 7 0 0 9 2 7 15 9 13 2
5 9 13 15 0 2
21 14 15 13 0 0 9 1 9 2 15 13 13 2 13 14 13 2 7 3 13 2
18 7 10 0 9 2 9 2 9 1 9 0 1 9 1 9 0 9 2
13 9 3 13 13 1 15 2 10 9 1 15 13 2
8 15 4 0 9 13 3 13 2
15 9 7 9 9 13 13 0 9 9 9 7 10 0 9 2
7 7 13 1 9 12 9 2
19 3 13 2 1 9 2 3 0 1 10 12 9 9 7 0 1 12 9 2
11 7 3 7 15 13 3 9 13 9 3 2
15 15 3 13 13 9 1 9 2 15 13 3 14 12 9 2
12 7 1 10 0 9 15 13 13 10 0 9 2
18 9 1 0 9 15 13 1 9 11 2 15 3 10 9 13 0 9 2
22 16 15 9 13 7 13 0 2 15 1 9 13 2 13 3 9 2 9 2 1 9 2
30 0 12 2 12 2 1 9 15 0 3 12 9 15 3 4 13 13 14 0 9 2 7 3 3 9 7 0 9 9 2
7 1 11 13 9 1 9 0
2 11 2
17 0 0 9 2 15 4 13 9 9 2 13 1 0 9 0 0 2
9 13 15 3 9 1 11 11 11 2
20 0 9 13 2 16 9 1 9 13 1 9 2 3 13 9 1 0 0 9 2
10 0 9 15 1 11 13 9 1 9 2
13 2 9 9 13 1 3 3 0 9 2 2 13 2
16 9 1 15 13 3 0 0 9 7 13 14 1 9 0 9 2
6 9 11 13 1 11 9
2 11 2
17 1 9 0 9 11 11 13 9 11 11 0 13 0 9 9 9 2
31 2 15 2 15 15 3 13 2 13 9 2 1 15 9 3 13 1 9 9 2 3 9 1 9 1 9 2 2 13 11 2
20 1 9 11 4 9 11 13 1 9 7 13 7 9 2 15 13 0 9 13 2
18 2 13 7 2 16 15 1 10 9 9 3 3 13 2 2 13 11 2
8 11 13 9 2 7 15 15 2
9 9 4 3 13 1 9 1 9 2
7 10 9 13 0 0 9 2
15 11 11 2 9 0 9 2 13 4 15 12 9 0 9 2
10 12 9 15 13 1 9 9 0 9 2
11 13 4 3 0 9 7 13 4 9 9 2
9 3 1 9 4 4 13 1 9 2
11 13 7 2 16 15 3 3 13 3 15 2
17 11 11 2 9 9 7 0 9 2 1 9 9 2 1 9 9 2
21 11 11 2 9 11 2 16 9 2 15 1 12 9 13 0 0 9 2 13 9 2
22 1 9 1 9 11 2 15 13 10 9 0 9 2 4 7 3 13 1 9 9 9 2
25 11 11 2 9 11 2 13 13 2 16 4 13 10 0 0 9 16 9 7 13 4 1 15 0 2
14 3 4 15 13 9 7 15 4 13 14 1 0 9 2
17 11 11 2 9 11 2 10 0 9 13 2 7 1 9 4 13 2
21 11 11 2 0 9 11 2 16 13 15 0 0 9 2 3 13 3 3 9 9 2
20 1 10 9 15 10 0 9 13 10 9 7 13 9 2 16 3 15 7 13 2
26 11 11 2 11 2 2 9 0 9 9 2 1 0 0 9 4 15 13 1 0 9 2 3 1 9 2
24 11 11 2 11 2 2 9 0 9 9 2 13 9 7 3 13 9 9 1 3 0 0 9 2
27 13 9 13 1 9 2 13 2 16 13 0 2 16 4 16 9 13 15 1 9 1 9 7 1 9 9 2
35 11 11 2 11 2 2 9 0 9 2 13 3 0 2 16 13 14 9 1 9 7 3 4 13 13 9 0 16 10 2 15 4 15 13 2
13 16 9 9 13 9 9 3 2 3 15 15 13 2
14 11 11 2 11 2 2 9 2 13 4 9 1 9 2
12 16 9 11 13 9 2 3 13 15 1 9 2
22 11 11 2 11 2 2 9 0 9 2 13 2 16 13 9 2 7 3 13 14 9 2
21 13 15 2 16 9 4 13 16 9 2 7 0 12 9 13 15 9 2 16 13 2
5 11 1 9 10 9
10 9 9 15 13 1 11 13 1 11 11
15 3 1 9 13 1 11 11 12 2 0 9 0 0 9 2
22 1 0 9 9 7 9 1 0 9 9 13 11 9 0 0 9 1 9 12 7 12 2
43 1 9 9 11 11 13 0 9 10 9 9 9 0 9 2 0 7 0 9 2 9 9 2 9 9 2 9 9 2 9 7 9 7 3 9 0 0 9 1 9 0 9 2
11 9 9 4 15 13 13 9 0 9 9 2
14 1 9 4 1 11 13 3 2 7 9 11 11 11 2
15 9 4 1 9 13 13 0 9 9 7 12 1 12 9 2
18 0 12 13 1 9 9 3 1 9 9 0 9 9 7 9 0 9 2
8 4 3 13 3 9 10 9 2
29 9 11 11 11 3 11 13 2 16 13 2 16 1 15 4 13 9 1 9 9 2 2 13 15 3 3 0 2 2
11 13 7 2 15 4 15 13 13 10 9 2
13 9 4 15 1 10 9 13 13 0 9 9 9 2
19 13 4 14 3 13 0 9 1 0 9 2 15 4 13 14 1 0 9 2
24 9 11 11 2 11 11 7 11 11 3 11 3 13 2 16 13 13 1 11 3 13 0 9 2
16 2 9 1 10 9 4 1 0 9 4 13 16 0 9 9 2
11 7 4 9 13 3 0 2 2 13 11 2
10 13 7 2 16 9 4 3 13 3 2
24 11 13 2 16 13 2 15 4 13 13 0 9 2 7 15 1 10 9 13 15 0 7 13 2
1 3
20 9 9 11 2 11 2 11 2 4 15 13 1 9 13 9 11 11 2 11 2
23 1 9 0 9 9 11 1 11 15 3 1 9 1 0 9 13 9 9 11 11 2 11 2
10 9 11 4 3 4 13 1 12 9 2
23 11 13 3 0 9 7 9 9 9 7 1 9 12 13 1 9 11 2 11 3 1 11 2
10 0 9 4 15 14 13 13 1 0 9
2 11 2
18 1 9 0 9 11 11 4 15 0 0 0 9 13 13 1 0 9 2
31 2 15 4 15 13 9 7 3 4 10 9 13 13 1 9 2 1 15 1 0 9 13 0 9 2 2 13 11 9 11 2
15 13 3 2 16 13 10 0 9 1 9 11 7 0 9 2
35 13 15 7 2 16 0 9 0 9 1 0 9 2 15 13 0 9 2 1 9 13 7 4 13 9 2 15 4 9 0 0 9 3 13 2
18 2 13 7 0 0 9 2 16 4 15 10 9 13 2 2 13 11 2
28 9 0 9 11 11 1 9 1 0 9 13 2 16 13 0 9 0 9 2 16 13 0 9 2 7 0 9 2
15 2 1 9 10 9 1 0 9 13 3 13 7 9 11 2
10 15 4 15 3 13 2 2 13 11 2
20 9 2 16 4 9 0 9 13 0 9 2 13 1 11 9 11 9 1 11 2
17 2 3 15 9 11 13 2 10 9 13 0 9 2 2 13 11 2
29 9 0 9 11 11 13 2 16 9 1 9 9 1 11 13 11 3 2 16 13 13 9 3 3 2 16 13 9 2
20 11 11 13 1 0 9 1 9 0 9 9 10 9 2 16 4 13 1 11 2
35 0 12 9 9 1 0 0 9 9 13 3 1 9 0 9 1 11 9 0 1 9 0 9 1 11 7 1 0 9 0 2 0 9 2 2
20 13 15 3 1 9 9 0 0 9 11 11 11 2 15 13 9 9 11 11 2
35 2 15 13 3 1 11 9 7 13 1 15 2 16 4 9 1 9 13 10 9 7 9 2 2 13 0 9 0 1 0 9 0 9 0 2
4 11 9 11 13
2 11 2
21 9 9 9 11 11 13 13 9 0 9 1 0 9 9 11 1 0 2 0 9 2
24 0 9 1 9 13 9 1 9 2 7 1 15 9 13 9 1 2 0 9 0 9 9 2 2
54 0 9 13 11 1 0 2 7 13 15 7 2 16 4 15 11 13 3 13 15 9 1 15 0 2 2 15 0 13 9 3 13 7 15 0 3 13 0 13 2 1 15 9 13 7 3 13 10 9 1 10 9 2 2
34 11 3 13 2 16 4 13 0 2 16 4 15 1 9 1 9 13 13 9 10 9 1 0 9 2 15 13 13 3 1 9 1 9 2
6 9 15 13 13 1 11
2 11 2
25 0 9 11 13 1 0 9 1 0 0 9 9 7 9 0 11 7 10 9 3 13 0 0 9 2
10 13 15 3 9 0 9 11 11 11 2
20 10 9 9 9 1 9 0 9 4 14 13 14 9 9 2 7 7 0 9 2
29 3 3 13 1 11 9 3 12 9 9 7 9 2 15 13 13 9 9 9 1 12 9 1 3 12 9 0 9 2
16 1 11 1 11 0 9 3 13 2 7 9 3 13 0 9 2
26 1 9 13 0 2 16 16 13 9 2 4 9 13 10 9 7 9 2 2 16 15 13 1 9 2 2
6 9 11 2 11 2 11
6 13 9 1 9 13 0
2 11 2
16 0 9 0 9 11 2 11 2 11 3 9 13 9 9 9 2
6 10 9 13 11 11 2
24 9 9 1 0 0 0 0 9 13 0 0 9 13 1 12 2 9 0 9 9 9 7 9 2
28 9 13 13 9 7 9 9 2 10 9 2 9 2 0 9 7 9 9 2 3 7 9 9 2 9 7 9 2
21 1 0 1 3 4 13 13 9 9 0 7 0 9 1 9 2 15 4 9 13 2
17 1 0 9 1 9 13 1 12 9 2 13 15 7 3 0 9 2
14 0 0 9 13 12 2 9 7 12 2 9 0 9 2
1 3
16 9 0 9 9 1 12 5 9 11 11 13 3 9 9 11 2
61 9 13 12 9 2 0 11 11 7 0 0 11 0 2 11 3 2 0 9 13 9 2 11 2 0 2 11 2 2 0 11 5 11 11 2 2 11 0 2 11 2 2 11 11 5 0 11 5 11 2 11 2 7 11 2 0 9 5 11 2 2
6 9 9 13 14 9 2
16 1 9 13 3 9 0 9 1 0 11 11 11 2 1 11 2
10 4 13 1 0 9 9 7 9 9 2
25 9 13 1 9 3 1 0 7 0 11 13 1 0 9 0 9 2 1 15 13 2 16 13 0 2
8 13 15 3 0 7 0 9 2
22 1 0 0 9 9 1 11 4 3 1 11 11 1 15 9 13 7 0 11 1 11 2
25 15 13 0 15 2 16 2 13 9 2 7 13 0 1 11 1 11 1 12 2 9 12 2 9 2
8 3 15 13 0 0 9 11 2
4 9 11 13 11
2 11 2
17 11 13 14 0 9 2 7 0 9 2 15 15 13 1 10 9 2
21 13 15 3 9 10 0 9 11 11 1 9 9 9 1 9 1 0 9 9 11 2
17 11 15 1 11 13 0 2 9 9 2 2 0 1 9 0 9 2
22 0 9 1 9 9 10 0 0 0 9 1 0 9 13 0 9 9 2 9 2 2 2
53 1 9 0 0 0 9 1 9 9 2 9 2 2 10 9 4 3 13 2 2 13 1 0 9 0 9 1 9 14 12 5 9 11 2 12 5 11 12 2 12 5 11 12 2 12 9 9 7 12 9 0 9 2
12 0 9 9 2 15 13 9 11 2 13 9 2
18 14 9 9 13 0 2 16 12 5 0 0 9 13 0 9 9 11 2
10 11 1 9 13 3 0 7 0 9 2
7 11 13 7 1 9 11 2
23 12 12 1 15 1 9 13 3 3 11 2 12 15 3 13 1 0 0 9 2 11 12 2
10 12 9 1 9 13 14 1 0 9 9
2 11 2
14 3 1 10 9 15 0 9 13 1 0 9 0 9 2
27 9 0 9 0 9 1 9 0 9 13 2 16 15 9 13 2 1 9 13 7 9 1 12 2 12 9 2
12 1 10 9 0 9 2 9 2 13 15 0 2
11 3 1 9 2 3 13 9 3 3 15 2
20 9 9 1 11 12 11 2 11 13 2 2 0 9 13 3 13 1 0 9 2
7 9 3 13 14 12 9 2
37 16 13 1 9 12 0 9 2 13 13 12 9 2 7 13 12 9 2 16 4 13 9 1 9 1 9 9 3 2 7 13 12 9 1 12 9 2
10 13 15 2 16 0 4 13 0 9 2
8 9 9 7 3 13 0 2 2
34 9 13 9 2 16 1 0 9 1 0 9 2 3 13 9 1 9 1 0 9 9 2 13 9 3 3 3 7 9 15 1 15 13 2
13 13 1 15 0 9 2 0 9 13 1 9 9 2
20 15 3 13 13 1 0 9 1 9 2 7 9 15 13 13 2 3 9 13 2
26 9 2 16 7 1 9 4 13 0 13 3 12 9 1 12 9 16 12 1 12 2 1 10 9 13 2
32 3 9 0 9 1 0 0 9 11 11 13 2 16 9 9 13 1 15 1 15 7 1 10 9 13 3 13 1 9 10 9 2
13 3 13 2 16 9 13 3 0 14 1 0 9 2
8 13 15 13 3 9 10 9 2
12 9 3 13 9 13 1 0 9 7 1 9 2
6 3 13 1 15 9 2
7 15 3 13 9 0 9 2
27 7 7 15 3 13 2 16 9 13 3 16 10 0 2 7 15 7 3 2 16 1 9 9 13 9 3 2
10 1 11 12 1 15 13 1 0 9 2
13 13 9 2 16 13 1 10 9 1 0 9 9 2
16 1 10 9 13 15 0 9 2 3 13 0 9 0 9 13 2
7 9 11 13 1 9 11 11
1 11
29 9 0 9 11 11 7 9 0 11 11 12 13 3 1 0 9 9 0 9 1 11 2 15 13 9 1 11 11 2
14 11 15 1 9 13 1 9 0 9 9 11 7 11 2
25 3 7 13 2 16 4 0 9 1 12 2 9 13 10 9 2 1 10 9 15 11 2 11 13 2
14 9 9 3 13 1 15 13 10 9 10 9 11 11 2
20 11 2 11 13 2 16 4 1 10 9 3 13 13 0 9 9 9 1 11 2
10 9 0 0 9 4 3 13 13 11 2
19 9 0 11 1 11 12 7 3 10 9 13 9 11 1 9 1 0 9 2
25 2 13 9 1 9 7 13 15 2 16 13 0 2 16 4 12 9 13 13 10 9 2 2 13 2
14 1 15 7 0 9 0 9 13 0 9 11 1 9 2
15 10 9 15 4 13 2 9 7 13 2 16 15 13 9 2
20 1 9 3 13 9 0 11 11 2 15 13 2 16 10 9 13 12 9 11 2
20 11 2 11 4 1 0 13 1 9 0 9 7 0 9 1 0 9 0 9 2
8 2 0 9 2 13 3 7 13
9 9 13 9 0 9 7 9 10 9
2 11 2
22 1 9 13 12 9 2 15 15 13 1 9 9 13 0 9 11 3 1 12 9 9 2
13 13 1 15 7 12 0 9 9 11 7 0 9 2
13 11 15 3 13 9 9 9 1 11 12 11 11 2
28 0 9 13 12 0 2 9 2 2 1 15 12 3 1 10 9 13 0 9 1 9 2 13 1 9 0 9 2
18 9 9 11 2 11 2 15 13 1 10 9 2 0 9 11 2 11 2
18 15 15 3 13 13 2 1 10 9 1 0 9 9 11 13 0 9 2
17 1 0 9 13 3 9 0 9 11 7 9 10 9 11 2 11 2
37 0 9 13 9 0 16 2 0 9 2 1 9 2 1 15 13 11 2 11 2 2 9 1 9 12 9 1 0 9 1 0 9 1 0 0 9 2
20 9 12 2 9 3 13 3 14 9 12 9 2 1 9 3 15 13 1 9 2
14 16 4 13 9 2 13 1 9 3 9 12 12 9 2
20 1 9 9 15 9 3 13 1 9 2 3 13 9 1 11 7 12 12 9 2
8 2 3 15 13 1 0 9 2
20 3 7 13 1 11 2 13 1 9 7 15 9 13 2 2 13 11 2 11 2
15 1 12 9 15 13 1 11 2 3 1 9 7 4 13 2
13 1 0 9 13 9 12 2 9 0 9 0 9 2
19 9 13 1 9 9 9 7 9 2 0 9 3 13 1 10 9 12 9 2
13 15 12 0 13 9 9 9 1 12 1 12 9 2
13 0 1 9 13 1 0 0 9 1 9 1 11 2
19 9 3 1 0 9 13 14 12 9 9 1 9 2 10 9 7 9 9 2
7 1 0 9 15 3 13 2
15 9 1 15 15 7 9 2 15 9 9 13 2 3 13 2
23 2 12 1 9 15 3 13 2 16 3 13 14 12 9 1 9 2 2 13 11 2 11 2
16 1 15 13 10 9 0 15 2 16 0 9 13 7 13 13 2
10 3 15 3 9 9 10 9 3 13 2
6 11 2 1 9 9 13
2 11 2
15 9 9 11 15 1 9 13 13 10 0 9 7 0 9 2
19 11 15 3 1 9 1 9 0 0 0 0 9 1 11 13 9 9 11 2
16 2 13 0 9 2 16 4 15 15 15 13 2 2 13 3 2
29 1 10 9 4 15 14 9 0 9 13 13 9 0 1 0 2 0 9 2 15 1 9 9 11 13 9 7 9 2
33 2 1 10 9 3 3 14 2 16 10 9 13 14 0 9 2 1 10 9 4 15 13 13 0 9 2 15 13 2 2 13 11 2
38 13 10 9 7 9 4 1 15 13 0 3 1 9 9 2 16 14 10 9 2 7 7 3 13 3 2 9 7 9 2 13 15 3 7 13 0 9 2
5 0 9 13 13 9
2 11 2
15 0 0 9 0 1 9 7 9 13 1 10 9 13 9 2
27 13 15 3 11 1 9 1 9 0 9 2 15 1 9 0 9 9 1 0 0 9 13 0 9 0 9 2
13 1 10 9 4 9 13 0 9 9 0 0 9 2
26 0 13 0 7 0 9 7 1 9 4 13 9 9 2 13 1 11 11 11 1 0 9 0 0 9 2
28 13 2 16 1 12 7 12 9 10 9 13 0 9 2 1 0 13 13 9 0 2 7 13 2 13 9 2 2
20 9 0 9 11 11 13 2 16 13 9 1 0 9 9 1 9 7 0 9 2
5 1 11 13 9 9
2 11 2
37 0 9 11 3 1 9 11 13 2 16 4 1 9 1 9 13 4 13 9 12 0 0 9 2 15 3 4 13 1 0 0 11 3 1 0 9 2
25 1 11 7 13 0 0 0 9 2 7 9 9 2 3 4 0 9 13 9 15 9 0 0 9 2
23 1 10 9 15 3 1 9 11 13 1 9 0 9 9 1 0 0 9 1 9 1 11 2
18 11 14 13 2 16 9 0 9 1 9 0 9 13 1 10 9 0 2
11 1 9 4 1 9 3 13 1 9 9 2
1 9
23 9 12 0 9 2 11 11 1 11 7 11 11 1 11 2 4 13 4 13 1 0 9 2
30 3 3 13 9 2 3 12 9 0 13 2 16 4 13 2 0 9 2 2 3 4 15 13 0 9 0 15 12 9 2
16 14 15 3 9 12 9 3 13 1 15 2 15 13 1 9 2
19 1 9 2 15 0 9 13 7 13 2 13 2 16 3 0 9 13 0 2
37 0 9 0 7 0 9 4 15 13 13 9 1 9 2 1 15 4 9 0 11 2 15 15 3 13 1 9 0 9 2 13 0 3 9 1 9 2
21 2 15 9 2 15 9 2 2 13 3 3 0 9 2 16 15 13 13 0 11 2
21 15 15 13 1 9 2 16 9 10 0 9 1 0 9 13 0 0 9 3 9 2
44 0 9 13 13 2 16 15 0 15 13 2 16 4 11 4 3 7 3 13 2 7 16 11 9 4 13 9 9 2 3 10 2 15 4 13 9 7 9 9 0 11 1 11 2
7 6 2 0 0 9 9 2
11 9 11 13 0 2 16 0 7 3 0 2
5 3 10 0 9 2
29 1 0 9 7 10 9 13 13 9 2 15 15 1 0 0 9 2 7 3 3 3 1 0 2 0 9 2 13 2
26 0 9 0 9 1 15 13 13 9 2 1 15 13 2 11 4 13 7 9 1 11 15 1 15 13 2
85 0 9 9 2 1 15 13 9 13 2 4 7 13 0 13 7 0 9 0 2 11 15 13 13 13 2 16 15 4 13 14 9 2 7 11 4 3 13 13 1 15 2 16 15 2 0 9 2 2 15 1 9 0 9 13 11 2 13 9 2 3 15 4 13 7 3 13 1 0 9 2 10 2 15 15 15 13 2 7 1 10 9 4 0 2
35 9 2 15 15 13 1 9 3 1 9 9 11 1 11 2 7 9 11 13 10 0 9 0 9 2 13 1 9 2 15 13 0 9 3 2
19 9 9 1 11 13 9 7 9 2 16 0 9 1 9 13 9 1 9 2
28 7 14 0 9 1 9 13 2 16 16 4 1 0 9 1 9 15 13 2 13 4 0 9 13 1 0 9 2
3 3 1 9
16 11 15 13 1 12 9 9 1 15 3 16 1 0 12 9 2
3 0 0 9
3 9 13 9
13 13 9 2 15 13 9 1 9 11 2 1 9 2
34 16 9 9 9 7 11 13 2 16 1 0 0 9 13 3 0 7 0 9 2 3 13 2 16 15 1 15 13 1 3 0 9 13 2
46 2 1 9 9 7 9 9 1 0 9 1 9 9 13 3 16 12 9 9 7 15 13 13 2 16 1 10 9 13 1 9 1 9 9 2 2 13 1 9 11 0 9 11 11 11 2
17 1 10 9 13 9 9 1 9 1 9 13 3 9 1 0 9 2
27 16 1 9 9 4 3 13 9 9 2 13 13 1 9 2 3 9 1 10 9 9 13 1 9 10 9 2
21 10 9 1 0 9 13 3 15 2 15 15 13 13 0 9 1 0 9 9 11 2
20 1 9 1 9 9 4 3 1 10 9 1 0 9 12 2 9 12 13 9 2
11 9 9 11 13 0 13 3 1 0 9 2
20 1 9 0 4 13 3 12 12 9 2 1 15 15 1 0 9 13 10 9 2
15 1 9 9 9 11 11 9 13 3 1 0 9 13 9 2
8 2 13 15 9 9 0 9 2
16 9 1 9 13 13 0 2 16 1 9 9 9 2 2 13 2
20 11 2 3 16 11 2 14 13 9 2 10 0 9 0 1 0 9 9 13 2
11 12 13 2 16 9 9 4 13 0 9 2
19 1 9 0 9 0 9 11 11 11 13 9 10 9 1 9 1 0 9 2
19 0 9 10 9 13 1 9 2 16 1 9 9 4 13 13 14 0 9 2
12 11 2 11 2 11 13 0 9 1 11 7 11
2 11 2
19 9 1 0 9 0 2 0 9 3 1 11 13 9 0 9 11 2 11 2
23 13 2 16 1 9 10 0 0 9 0 9 13 3 0 3 13 0 9 7 13 1 9 2
19 1 11 2 15 13 12 1 12 0 0 9 2 3 11 11 13 0 9 2
16 13 15 1 15 9 0 0 9 11 11 2 15 13 3 9 2
26 3 13 0 9 1 3 16 12 0 9 9 2 9 7 9 9 2 1 15 15 13 1 9 0 9 2
20 13 2 16 0 9 13 3 1 0 9 0 0 9 7 0 1 9 0 9 2
22 11 3 13 0 2 16 0 9 3 13 0 9 7 13 0 9 1 11 7 0 11 2
32 1 9 0 9 11 11 13 2 16 1 9 1 9 0 9 13 9 3 0 9 9 2 16 4 15 1 15 13 1 0 9 2
5 11 13 2 0 9
2 11 2
31 2 0 9 2 0 9 9 11 11 1 0 2 0 9 13 11 11 2 0 9 0 0 9 2 11 2 9 9 11 11 2
31 9 9 11 1 0 9 2 16 2 9 2 11 1 11 13 9 2 13 11 1 9 0 9 2 16 4 15 13 1 9 2
27 2 13 7 3 9 2 16 13 3 0 3 13 0 9 2 16 15 13 0 0 9 2 2 13 9 11 2
23 11 3 13 2 16 15 1 11 3 13 15 2 15 13 7 13 1 0 9 9 0 9 2
12 10 9 3 13 0 0 9 2 13 9 11 2
9 1 9 0 9 13 0 9 0 9
2 11 2
14 9 0 11 13 1 0 9 13 0 9 12 0 9 2
11 13 15 1 9 2 15 13 11 1 9 2
36 1 0 9 9 9 12 3 13 2 16 3 10 0 9 13 0 0 9 1 0 9 9 2 15 1 0 9 13 1 9 12 1 0 0 9 2
33 16 13 1 0 9 11 2 13 1 9 9 11 10 9 9 12 9 9 2 15 4 1 9 12 2 12 13 1 0 9 7 11 2
15 0 9 11 3 9 9 12 13 14 14 12 9 9 9 2
12 0 9 15 3 3 13 13 3 1 0 9 2
25 11 13 1 0 9 9 1 3 0 9 9 0 0 9 7 9 0 9 2 3 13 16 0 9 2
38 0 9 11 13 2 16 9 11 7 9 0 0 9 0 13 1 10 9 0 9 0 9 1 0 9 11 2 15 3 13 13 1 0 9 9 7 9 2
29 16 13 1 9 11 2 10 0 9 3 2 3 1 0 9 13 9 9 1 0 9 1 0 11 1 0 0 9 2
18 1 9 2 15 13 11 1 9 2 9 9 9 13 10 0 0 9 2
35 1 12 9 2 9 2 15 4 9 1 0 9 13 2 7 4 3 13 14 9 12 1 9 9 0 1 0 9 1 9 14 12 9 9 2
11 9 0 9 13 10 0 9 1 9 12 2
18 0 9 13 3 9 9 2 15 13 9 9 2 14 1 9 0 9 2
2 9 13
2 11 2
9 1 0 9 13 3 9 0 9 2
14 9 9 13 12 9 2 9 2 9 9 9 3 13 2
18 13 9 9 12 9 13 1 12 5 7 0 9 13 1 9 12 9 2
22 9 1 0 2 9 13 12 2 9 2 3 4 1 12 9 13 9 1 0 9 9 2
4 12 12 9 2
3 1 0 9
2 11 2
25 0 12 12 9 15 13 3 9 1 0 9 1 11 2 3 9 11 11 13 0 9 2 0 11 2
27 9 0 1 0 13 9 0 0 0 9 7 13 3 13 1 15 2 15 4 13 3 0 9 1 0 9 2
16 11 13 12 2 12 9 11 7 0 1 9 12 9 0 9 2
8 11 13 3 3 1 11 13 2
19 11 13 9 1 12 9 7 1 0 9 13 7 1 0 9 12 2 9 2
25 3 0 11 2 9 0 9 0 9 0 0 9 2 3 13 0 11 2 0 9 13 1 9 3 2
4 3 1 9 12
1 3
20 0 9 3 13 9 2 15 13 1 9 0 9 1 0 9 9 3 1 9 2
14 3 7 10 9 2 16 3 2 0 9 2 4 13 2
42 0 9 0 9 1 9 1 0 9 2 15 1 9 0 9 13 9 0 9 7 13 10 0 9 1 0 9 2 13 1 0 9 13 9 1 9 1 9 12 9 9 2
3 11 13 9
2 11 2
15 0 0 9 11 3 13 0 9 7 13 12 0 9 9 2
16 1 0 9 0 11 0 9 9 1 9 12 13 12 9 9 2
14 10 1 9 0 9 13 0 9 1 9 7 0 9 2
17 11 2 15 1 12 9 13 0 9 2 3 3 13 1 0 9 2
15 15 1 15 13 9 2 16 10 0 9 11 3 13 0 2
22 9 9 11 11 13 2 16 10 0 9 2 3 0 0 9 2 13 1 9 0 9 2
20 10 9 7 13 1 0 7 13 1 15 1 0 9 0 9 1 9 0 9 2
5 0 9 13 1 9
3 0 11 2
23 0 9 0 9 3 13 1 0 9 1 0 0 0 9 1 11 2 11 2 0 9 2 2
11 0 9 1 9 13 0 9 1 0 9 2
22 1 0 0 9 3 13 10 9 9 2 11 2 2 15 15 1 11 13 9 0 9 2
25 3 9 15 13 0 0 0 9 2 9 2 0 9 11 11 2 15 15 13 13 0 9 11 11 2
15 10 9 13 11 13 1 0 9 16 0 9 1 0 9 2
15 9 4 3 13 1 9 0 9 1 0 11 3 1 9 2
5 9 11 13 0 11
2 11 2
25 16 13 3 1 0 9 9 9 11 11 11 2 13 10 9 9 1 9 0 9 1 9 11 11 2
7 0 9 13 9 9 11 2
18 1 0 9 13 13 9 1 0 9 2 13 13 9 1 9 0 9 2
7 13 3 13 9 9 9 2
15 1 9 12 2 9 13 9 2 9 0 9 2 9 3 2
14 1 9 13 0 9 7 9 2 1 15 10 9 13 2
10 15 13 15 2 16 4 1 9 13 2
12 15 4 13 4 13 3 1 9 9 0 9 2
8 9 9 13 0 1 12 9 2
4 11 13 0 9
2 11 2
12 0 9 1 9 0 7 9 13 3 11 11 2
24 9 0 12 9 9 2 9 11 2 11 7 11 11 2 13 1 12 5 1 12 9 2 9 2
17 9 0 9 1 0 9 15 13 1 12 5 1 12 9 2 9 2
15 0 9 9 13 3 12 12 2 15 13 9 1 12 5 2
23 0 0 9 9 11 0 1 9 15 13 1 12 5 7 9 13 1 0 9 1 12 5 2
14 3 15 13 9 0 9 2 1 12 9 1 12 5 2
22 7 16 11 11 3 13 0 0 9 1 0 9 12 2 13 15 1 9 9 1 9 2
23 1 0 12 9 0 9 13 9 1 9 12 9 2 9 7 0 9 13 7 1 0 9 2
13 3 0 9 0 13 9 10 0 9 7 1 11 2
12 3 15 13 1 11 7 1 11 1 12 12 2
4 9 9 15 13
9 0 9 9 1 9 13 9 0 9
22 9 9 0 9 2 15 10 9 13 0 9 2 4 1 9 9 0 9 13 1 9 2
25 0 9 4 13 13 12 9 9 1 15 2 16 15 1 15 0 9 0 9 3 13 12 2 9 2
46 9 9 2 15 4 13 1 9 0 9 2 13 1 0 9 9 9 11 1 0 9 1 0 9 1 15 2 16 3 4 13 9 1 9 9 0 1 9 0 9 1 0 7 0 9 2
24 0 0 9 10 9 9 13 9 1 9 0 0 9 1 0 7 0 1 9 0 9 1 9 2
21 3 4 13 4 13 9 9 0 0 9 2 0 0 7 0 9 1 0 0 9 2
20 10 9 4 3 13 4 13 1 9 1 15 2 16 1 15 4 13 9 9 2
14 3 1 9 0 9 7 9 4 13 0 0 0 9 2
24 15 15 3 13 0 9 9 9 1 9 0 9 7 9 0 9 7 13 9 1 0 9 9 2
10 1 0 9 9 15 13 1 0 9 2
20 1 0 9 7 0 9 4 13 9 13 1 9 1 9 9 13 0 0 9 2
37 1 10 9 2 15 13 0 9 0 9 7 9 2 13 0 9 13 9 9 3 0 7 0 1 0 0 9 2 16 0 9 10 9 3 13 0 2
19 9 7 13 13 0 9 2 15 13 9 0 7 0 9 1 0 0 9 2
12 1 0 9 9 9 4 9 13 1 9 9 2
27 3 4 0 9 9 3 13 2 13 1 9 9 9 11 1 9 9 0 9 1 9 7 1 10 0 9 2
5 0 9 13 0 9
8 9 13 0 9 3 0 9 9
2 11 2
21 0 9 0 9 13 0 9 1 9 9 2 15 4 13 0 2 0 7 0 9 2
15 9 1 9 13 12 2 9 10 9 2 13 1 9 9 2
25 9 13 0 9 0 9 9 2 9 1 9 9 7 9 10 0 9 9 9 10 9 1 0 9 2
35 9 16 3 0 9 0 9 13 9 0 9 7 9 2 3 7 13 9 2 15 13 13 1 0 9 2 0 9 9 1 9 1 0 9 2
21 9 13 0 9 9 1 0 9 7 9 2 13 7 4 0 9 1 9 7 9 2
14 9 9 1 9 4 13 9 0 9 7 0 0 9 2
23 1 9 1 0 9 4 13 9 9 0 0 9 2 9 9 9 7 9 9 1 0 9 2
26 0 9 4 13 13 10 9 7 9 2 15 15 4 13 1 9 9 9 7 1 9 9 1 10 9 2
29 9 2 10 9 15 4 13 1 9 2 4 13 13 9 9 2 16 13 1 0 9 3 0 9 9 0 9 9 2
11 3 13 13 0 0 7 0 0 9 9 2
15 9 13 13 0 9 1 9 2 13 15 9 9 1 9 2
18 3 12 9 9 7 12 9 9 13 9 0 11 1 9 9 0 11 2
20 1 0 9 4 11 13 10 9 14 0 0 9 2 7 7 0 9 7 9 2
15 1 10 9 3 11 13 1 9 2 9 7 9 0 9 2
18 0 9 9 13 2 16 0 0 9 3 13 3 3 16 1 0 9 2
4 9 13 0 9
12 16 9 3 13 0 0 9 2 9 9 3 13
33 0 9 9 2 15 13 3 0 2 13 0 2 9 9 10 0 9 2 3 13 9 13 0 0 9 9 2 3 12 9 2 9 2
21 1 0 9 2 12 9 2 13 10 9 3 3 3 2 7 7 3 13 3 0 2
18 1 9 9 3 13 0 9 9 2 15 13 3 12 0 9 1 15 2
21 9 9 12 3 13 1 12 5 10 9 1 12 2 9 2 3 4 9 3 13 2
22 9 13 1 9 12 9 2 0 12 9 1 10 0 9 1 9 12 2 9 10 9 2
15 0 9 0 9 13 0 2 3 0 1 9 9 1 9 2
20 1 12 9 0 9 14 12 13 2 3 12 13 7 0 12 2 2 2 13 2
22 3 13 9 9 11 2 0 9 10 0 9 2 7 15 1 12 5 2 1 12 9 2
19 1 9 3 13 2 0 2 9 9 0 9 1 12 5 2 1 12 9 2
30 9 9 11 13 7 1 9 9 9 12 13 3 7 9 11 2 15 13 1 12 5 2 1 15 13 9 0 12 5 2
12 13 3 1 9 2 16 9 13 3 0 9 2
14 3 1 0 9 2 7 15 3 13 9 1 0 9 2
38 9 9 0 9 13 0 2 1 3 16 12 9 13 12 0 9 2 1 15 1 0 12 9 12 2 2 2 2 9 9 3 2 14 2 1 12 5 2
15 9 13 9 11 2 15 13 1 12 5 2 1 12 9 2
18 9 1 0 9 0 9 13 3 3 16 1 9 2 7 13 0 9 2
28 1 9 0 9 0 9 13 12 9 2 1 15 3 13 14 12 2 12 2 11 11 7 0 11 12 2 11 2
18 1 0 0 9 13 9 3 0 9 2 15 15 13 1 12 9 9 2
34 13 7 9 7 0 0 9 11 2 13 4 9 0 2 16 15 15 1 0 9 2 1 0 9 7 1 0 9 2 13 3 12 9 2
13 0 9 13 3 1 9 9 11 7 12 0 9 2
1 3
31 9 9 1 11 1 9 15 1 9 13 1 12 9 1 9 1 9 0 9 2 16 1 9 13 1 0 9 1 12 9 2
25 11 13 13 0 9 0 9 1 10 9 1 0 9 12 2 9 1 11 7 12 2 9 1 11 2
17 0 9 13 9 1 0 0 9 2 3 1 9 9 7 0 9 2
15 0 9 1 0 9 7 9 13 13 9 0 9 1 9 2
9 9 0 9 3 13 12 9 9 2
19 9 0 9 1 9 1 0 9 13 1 9 1 0 9 3 1 12 9 2
15 3 12 9 0 9 13 1 0 9 0 9 1 0 9 2
5 0 9 1 9 11
2 11 2
24 0 9 11 2 15 0 9 13 12 9 9 2 13 13 0 9 1 0 9 1 0 0 9 2
23 4 13 9 0 2 0 2 12 1 9 7 9 0 2 2 9 0 2 9 7 0 9 2
9 1 9 0 9 15 13 3 3 2
40 9 1 0 9 13 1 9 12 9 2 4 2 14 13 9 1 9 12 9 7 1 9 0 9 3 12 9 2 16 0 9 0 9 9 13 3 12 9 3 2
10 11 13 1 9 1 12 7 12 9 2
20 1 9 0 0 9 15 4 13 3 1 9 9 9 2 15 13 0 0 9 2
14 9 9 4 13 3 9 9 9 2 3 3 0 9 2
9 9 9 13 1 0 9 7 11 2
5 9 12 13 0 9
11 0 9 0 1 0 9 13 3 13 0 9
32 9 1 12 0 9 9 2 0 9 7 9 0 0 7 0 9 15 1 0 9 13 1 11 2 16 4 13 1 0 0 9 2
11 9 9 13 10 0 9 1 9 0 9 2
28 1 0 9 15 13 0 0 9 2 1 15 13 13 9 2 9 7 9 7 15 3 13 9 1 9 0 9 2
23 1 9 10 7 15 9 13 15 1 10 0 0 9 7 13 10 9 3 13 0 0 9 2
27 1 0 9 2 15 13 1 0 9 1 0 9 2 15 1 9 9 13 9 0 1 14 0 12 9 9 2
46 1 0 12 9 2 15 9 9 9 12 13 1 9 9 0 9 2 13 9 0 9 2 9 9 1 0 9 2 9 0 9 1 9 2 9 0 9 1 0 9 7 9 0 0 9 2
27 0 9 13 13 0 9 9 1 10 9 2 0 9 3 0 9 7 9 0 7 0 9 1 9 0 9 2
24 1 9 2 16 4 9 13 13 9 1 9 9 7 9 2 7 13 9 2 16 10 9 13 2
14 3 0 9 15 13 3 0 0 9 2 15 13 13 2
15 16 4 13 3 0 9 2 3 4 15 13 10 0 9 2
20 13 15 2 16 1 9 9 0 0 9 9 9 3 3 13 1 9 0 9 2
25 1 0 9 15 10 9 2 3 11 7 11 2 13 2 16 1 0 9 13 0 2 3 0 9 2
18 9 13 9 1 12 0 0 9 2 10 9 15 13 1 9 10 9 2
22 13 1 15 9 0 9 0 0 9 2 9 1 3 0 9 9 7 0 9 0 9 2
24 3 3 15 13 1 9 0 9 7 9 2 9 9 0 9 7 0 9 7 9 0 9 9 2
13 13 15 3 9 15 2 3 4 0 9 13 13 2
22 16 13 4 15 1 9 13 2 13 15 1 0 9 13 0 9 9 12 1 0 11 2
6 7 1 11 9 3 13
2 11 2
23 1 0 9 13 1 0 9 11 3 12 9 2 15 13 1 12 9 3 16 1 0 9 2
28 1 9 0 0 9 1 11 1 0 9 13 1 9 9 2 3 15 9 0 9 1 9 12 13 1 12 9 2
10 1 9 9 13 9 9 1 12 9 2
17 1 0 0 9 4 3 13 1 12 9 9 3 16 1 0 9 2
4 0 11 1 9
2 11 2
24 11 13 1 9 12 9 0 9 1 9 12 9 9 1 9 1 9 12 9 9 1 9 12 2
15 1 0 9 13 3 0 9 9 2 15 13 9 0 9 2
26 0 9 13 1 0 9 0 9 9 7 3 0 9 0 9 2 15 4 15 13 13 1 12 9 9 2
13 9 9 3 13 1 12 9 7 13 12 9 9 2
12 9 15 13 1 12 9 7 13 12 9 9 2
21 15 15 13 7 9 0 9 1 9 12 9 9 1 9 12 9 9 1 9 12 2
20 1 9 13 9 0 7 0 9 2 16 1 9 13 0 9 7 9 0 9 2
5 0 9 13 1 9
8 9 9 15 1 0 9 3 13
2 11 2
30 9 1 9 1 9 0 9 1 0 0 9 13 4 13 3 1 12 2 9 1 0 9 2 3 13 0 9 0 9 2
17 16 13 9 0 9 2 13 15 10 9 1 12 2 9 0 9 2
25 0 9 13 7 13 3 3 2 4 2 14 0 0 9 1 9 13 1 9 9 3 1 9 9 2
22 1 9 1 9 3 3 10 9 13 1 9 0 9 11 2 9 13 0 9 7 9 2
17 9 13 2 16 1 2 9 2 1 0 9 13 10 9 13 3 2
23 0 0 9 13 3 2 1 9 1 0 9 2 9 1 9 9 1 9 1 9 0 9 2
35 0 9 13 0 9 1 0 9 2 15 13 1 11 0 9 7 15 1 15 13 3 12 9 1 9 7 15 0 0 0 9 13 12 9 2
33 9 1 0 9 2 3 15 2 15 13 1 9 7 0 0 9 2 13 9 1 9 2 16 10 0 0 0 0 9 13 12 9 2
17 13 15 14 9 1 9 7 0 3 0 9 2 7 7 0 9 2
21 1 9 1 0 9 15 13 3 9 1 0 9 7 9 1 9 0 9 1 9 2
29 13 15 3 9 2 9 2 9 7 0 9 1 9 1 0 9 2 16 4 13 1 9 7 9 0 2 0 9 2
18 9 15 13 3 1 9 1 9 9 7 0 9 16 7 1 0 9 2
12 3 1 9 13 13 0 9 7 9 1 9 2
12 9 13 13 15 2 15 13 9 3 1 9 2
20 15 3 9 1 9 9 13 9 1 9 7 0 9 1 15 0 9 13 15 2
24 0 9 13 1 9 13 0 9 7 9 7 3 1 0 9 9 13 13 9 14 1 12 9 2
8 0 7 0 9 13 1 9 0
2 11 2
30 9 9 9 1 9 7 9 1 9 13 9 1 3 12 9 9 15 0 9 2 15 13 1 0 0 9 0 0 9 2
13 1 9 13 1 9 9 1 0 9 12 5 9 2
14 1 9 13 12 9 2 10 9 13 3 9 0 9 2
24 0 12 5 9 13 9 9 1 12 1 12 9 7 12 9 9 1 9 1 12 1 12 9 2
11 9 1 12 5 9 1 9 1 9 13 2
21 1 0 9 2 15 13 12 5 9 9 2 15 9 1 9 7 9 1 9 13 2
18 9 13 9 1 12 5 9 2 15 13 1 15 3 16 1 0 9 2
10 13 12 9 0 3 9 0 0 9 2
9 9 1 12 9 13 1 9 9 2
3 9 9 13
4 9 1 11 2
29 16 15 13 1 9 1 0 9 13 1 0 9 10 9 2 13 0 13 0 9 9 1 9 0 9 1 0 9 2
23 16 3 13 1 9 1 0 9 0 9 1 11 1 11 2 13 9 0 9 0 0 9 2
8 10 0 9 13 1 0 9 2
19 1 9 2 3 13 9 1 0 9 13 7 10 9 13 2 13 15 0 2
19 1 0 9 0 9 13 3 2 9 9 7 9 1 9 9 9 9 9 2
32 9 11 11 2 3 2 13 3 9 0 9 11 11 2 1 0 9 13 2 16 11 13 10 0 9 0 9 2 15 13 15 2
4 9 11 13 9
2 11 2
18 0 9 0 9 11 1 0 9 13 3 12 9 9 2 3 16 3 2
14 13 15 1 9 0 9 9 11 11 1 0 9 9 2
18 9 9 3 13 1 10 9 3 1 12 9 2 1 0 12 9 9 2
29 12 9 0 0 7 0 9 2 15 13 0 9 9 2 15 13 2 3 1 3 0 9 2 0 11 7 0 9 2
22 16 3 13 11 2 11 2 0 0 9 1 11 11 7 10 9 13 9 1 9 9 2
10 15 15 1 9 13 1 12 9 9 2
22 2 13 4 0 2 16 4 9 13 13 0 9 1 10 9 9 9 2 2 13 9 2
10 9 11 4 13 1 0 9 0 9 2
21 0 9 10 9 1 0 9 4 13 1 12 9 7 1 0 2 9 1 12 9 2
4 9 13 1 9
9 11 2 11 2 11 2 11 2 2
13 1 9 0 9 13 1 11 0 9 3 0 9 2
9 3 3 13 12 7 0 9 9 2
20 11 15 13 9 9 9 9 1 9 9 11 11 2 9 9 2 0 9 2 2
23 3 10 9 13 0 9 9 1 9 7 0 9 0 9 1 0 0 9 1 11 12 11 2
10 1 9 13 0 11 0 9 1 9 2
8 0 13 9 7 3 3 9 2
8 9 7 13 1 9 9 13 2
12 1 9 15 13 1 0 7 0 9 9 11 2
17 2 9 13 1 10 9 13 2 16 15 9 9 3 13 0 9 2
19 15 13 2 1 1 9 9 2 3 0 2 3 3 0 2 2 13 11 2
27 13 3 1 0 2 0 9 2 2 3 9 12 9 13 1 9 11 9 0 11 7 13 15 1 9 13 2
7 0 11 11 11 15 13 2
12 12 1 9 4 13 1 0 0 9 9 9 2
5 0 9 4 13 2
21 9 1 9 13 15 2 16 9 1 9 11 13 13 1 0 9 2 9 7 9 2
40 11 13 1 15 2 16 7 16 13 9 3 0 0 9 1 0 9 0 2 2 10 9 7 0 9 13 1 0 9 1 0 7 0 9 7 1 9 11 2 2
23 1 9 9 2 0 9 2 13 0 9 9 10 0 9 9 9 11 7 9 1 15 0 2
6 0 13 3 3 11 2
12 9 1 0 9 1 9 11 11 2 0 0 9
14 16 0 0 9 13 3 0 2 16 15 15 13 9 2
7 13 15 1 15 0 9 2
8 0 9 0 9 7 3 13 2
11 13 2 10 0 0 9 13 1 9 9 2
21 3 13 1 0 9 9 1 9 2 7 3 9 9 7 3 3 9 9 9 13 2
34 0 9 3 13 2 3 15 15 13 7 13 3 13 2 3 15 13 2 3 15 13 13 3 2 3 2 2 3 13 1 9 3 13 2
9 7 13 15 7 1 9 0 9 2
14 15 13 13 0 9 2 7 16 15 13 10 0 9 2
15 15 0 15 3 15 13 13 2 7 13 3 13 1 9 2
15 1 9 9 13 9 0 0 9 2 7 7 15 3 13 2
12 13 15 2 16 4 3 13 13 7 0 9 2
31 13 4 3 0 2 16 4 15 13 9 10 9 2 16 4 0 10 9 13 13 14 1 15 2 16 10 9 13 7 13 2
16 1 9 3 13 15 13 14 3 2 13 2 14 9 0 9 2
17 13 15 2 7 3 15 13 2 16 4 15 13 14 3 13 9 2
14 16 13 1 9 2 15 13 1 0 9 3 0 9 2
9 1 0 9 13 9 2 13 15 2
14 13 15 0 7 0 2 16 13 9 9 2 9 9 2
15 10 0 0 9 2 15 0 9 13 9 2 13 3 0 2
11 10 9 13 9 2 1 15 9 3 13 2
15 13 1 15 0 2 7 3 13 3 1 15 9 0 9 2
22 9 15 13 13 1 15 2 16 9 13 3 2 16 13 3 0 2 3 15 13 3 2
5 15 13 3 0 2
16 15 15 13 3 2 15 3 2 15 3 2 15 13 15 12 2
10 13 15 2 16 15 3 15 3 13 2
12 3 7 10 9 13 2 16 15 13 1 9 2
8 13 0 1 10 0 9 13 2
14 15 13 9 0 9 2 15 15 13 1 10 0 9 2
21 15 15 3 3 13 2 13 15 3 13 2 16 0 0 9 13 1 15 10 9 2
15 15 13 7 0 9 9 9 7 9 9 2 13 0 13 2
47 16 15 13 1 10 9 2 15 3 13 2 13 10 0 9 2 10 9 2 10 9 2 7 16 15 10 9 13 2 16 4 15 13 3 2 13 15 1 15 3 0 2 13 15 0 9 2
19 7 3 13 13 2 16 15 1 10 9 3 13 3 3 2 16 15 13 2
13 13 15 1 15 2 1 15 13 1 0 15 13 2
23 13 15 2 16 4 15 10 9 13 0 2 16 1 15 3 13 7 9 9 7 0 9 2
21 3 13 3 3 2 15 1 0 10 9 13 10 7 15 9 7 10 7 15 9 2
15 9 3 13 2 16 13 2 15 3 13 7 10 13 9 2
28 13 15 3 7 13 15 3 2 3 15 13 2 1 9 0 9 2 0 9 7 0 9 1 15 2 15 13 2
5 0 9 13 1 11
5 11 2 11 2 2
17 12 9 13 11 11 1 11 1 0 9 1 11 9 0 0 9 2
18 3 2 1 9 2 1 9 7 3 3 2 16 13 15 1 0 9 2
31 2 3 4 13 9 7 16 3 13 1 9 13 3 2 13 4 10 9 1 0 9 1 9 9 12 2 2 13 0 9 2
15 13 14 9 2 7 3 0 9 0 0 9 1 9 12 2
13 1 0 9 13 14 12 9 2 16 13 10 9 2
22 9 1 9 2 11 13 2 2 15 1 10 9 13 1 12 1 9 1 11 1 11 2
17 1 9 9 13 9 9 1 9 2 1 15 1 9 13 0 9 2
14 9 14 12 11 3 1 9 1 9 13 13 9 9 2
14 9 11 3 13 2 16 2 0 2 11 7 3 13 2
11 3 3 3 15 9 9 13 0 9 13 2
3 2 11 2
5 11 1 9 1 9
2 11 2
26 3 3 0 9 2 0 9 2 16 9 0 2 11 13 9 2 0 1 0 9 2 9 1 9 13 2
25 13 15 1 0 0 9 1 9 9 9 0 9 11 11 1 9 9 12 1 0 0 9 1 11 2
17 1 9 11 13 2 16 15 15 13 2 16 10 9 13 0 9 2
33 13 9 9 9 2 16 1 10 9 4 13 15 2 15 13 3 3 0 7 4 15 13 13 13 1 10 9 2 13 1 11 0 2
21 1 0 9 15 9 9 13 2 16 9 13 0 9 0 9 2 3 9 9 13 2
10 13 0 0 2 0 0 9 11 2 12
3 0 11 2
44 0 0 2 0 9 11 2 12 13 9 7 1 9 9 12 9 2 7 3 2 16 13 1 0 9 1 9 9 9 1 9 2 15 13 3 0 9 0 9 0 9 1 11 2
23 1 0 0 9 0 9 15 3 1 0 9 0 9 11 1 0 11 13 9 9 11 11 2
39 13 3 0 9 9 2 7 13 12 9 2 15 13 1 15 2 16 14 11 4 13 1 2 9 0 0 9 2 2 7 7 10 9 13 1 9 0 9 2
34 10 0 0 9 0 7 0 9 13 1 9 2 15 10 9 13 1 0 9 0 0 9 2 15 15 13 1 9 0 9 2 13 11 2
20 13 4 0 2 16 4 10 9 13 13 1 0 9 3 1 9 11 2 13 2
17 9 0 9 9 0 9 11 11 13 2 16 15 9 9 4 13 2
21 1 0 7 0 9 7 0 9 9 13 7 9 9 2 15 13 0 1 9 11 2
49 0 9 11 2 12 15 1 12 2 9 1 0 0 9 11 13 12 9 12 2 9 12 2 0 9 0 0 9 0 11 7 12 9 12 2 9 12 2 0 0 9 12 2 9 0 9 9 11 2
5 11 13 0 9 9
8 1 12 2 0 9 9 9 13
6 0 11 11 13 9 9
6 11 13 9 11 11 2
8 0 9 0 9 13 3 3 2
25 3 12 0 9 7 1 15 3 12 0 2 0 9 7 11 1 11 2 13 9 1 12 2 9 2
10 9 9 13 9 11 11 1 11 11 2
21 13 15 7 9 0 9 11 2 15 15 0 9 13 9 0 0 9 1 0 9 2
22 1 11 13 1 9 1 11 7 9 0 9 10 9 11 11 2 15 3 13 1 9 2
16 11 15 9 1 11 13 1 0 9 7 13 7 9 0 11 2
37 15 3 1 0 0 9 13 11 1 10 9 2 1 9 7 0 13 0 9 7 3 9 15 13 1 9 1 9 2 16 1 9 9 13 1 9 2
13 3 13 0 12 9 2 12 9 7 12 0 9 2
26 12 9 15 9 3 13 1 9 2 16 15 13 0 0 9 1 11 2 0 0 9 2 12 2 12 2
34 9 13 1 0 11 2 11 7 11 0 1 9 2 0 0 9 1 9 13 14 11 1 12 2 9 2 2 16 9 13 0 0 9 2
10 7 12 0 9 9 15 13 1 9 2
16 11 3 13 13 10 9 9 7 11 0 9 1 0 9 11 2
21 1 0 9 15 13 3 1 12 9 7 1 9 0 11 13 11 1 12 2 12 2
18 1 12 2 9 13 11 13 10 0 9 9 2 7 9 13 0 9 2
7 9 2 12 2 7 12 2
4 9 2 11 2
26 11 11 2 9 11 2 2 1 9 4 13 0 2 7 3 15 13 1 9 2 16 13 0 9 2 2
43 11 11 2 9 11 2 2 1 9 12 2 12 4 15 13 2 16 13 9 2 11 15 1 15 13 16 9 1 9 2 7 13 15 13 2 16 3 13 9 1 9 2 2
9 2 11 2 0 11 12 11 11 12
22 0 3 13 9 2 15 13 1 12 2 9 0 9 11 2 7 9 9 13 3 0 2
26 15 13 0 13 2 13 15 3 1 9 7 3 11 13 9 15 1 9 7 1 9 2 3 7 13 2
10 1 12 2 9 15 9 3 14 13 2
9 11 13 12 9 0 7 3 13 2
13 1 9 15 0 13 0 9 2 11 7 3 13 2
4 9 2 11 2
11 3 1 9 15 3 13 11 7 11 2 2
17 11 11 2 9 11 2 2 13 0 2 0 9 13 1 15 0 2
13 3 13 9 2 0 13 1 9 7 1 9 2 2
12 2 11 2 0 0 9 1 9 13 9 9 2
11 0 0 9 7 13 1 12 2 9 0 2
10 1 0 0 9 13 0 9 9 11 2
23 1 12 9 3 13 0 9 11 7 11 1 9 1 9 13 9 1 9 2 12 2 12 2
23 13 9 1 9 1 0 9 15 0 13 14 1 0 9 9 2 7 11 3 13 0 9 2
4 9 2 11 2
17 11 11 2 9 11 2 2 1 9 7 9 13 10 9 15 13 2
12 13 15 2 16 4 13 9 1 0 9 2 2
20 11 11 2 9 11 2 2 1 0 9 15 13 0 9 1 10 0 9 2 2
26 2 11 2 3 1 9 15 0 1 10 0 9 13 2 1 0 9 7 9 13 14 1 12 2 9 2
23 15 11 13 3 0 0 9 7 11 11 13 10 9 1 9 9 1 9 2 12 2 12 2
16 9 1 9 13 9 3 1 9 11 2 16 3 9 13 11 2
33 0 9 13 3 1 12 9 2 0 15 13 14 1 12 2 9 2 3 0 11 13 9 11 7 15 15 13 13 2 12 2 12 2
24 1 0 9 15 11 1 0 9 13 1 9 2 11 15 7 13 7 1 11 15 7 9 13 2
4 9 2 11 2
9 14 2 9 15 13 1 9 2 2
27 2 11 2 9 1 15 1 9 13 11 2 16 0 11 12 9 1 9 9 1 0 9 13 0 9 11 2
20 1 0 9 13 0 0 7 9 11 1 12 2 9 13 14 0 9 9 9 2
19 1 9 9 13 9 1 9 3 9 7 1 12 2 9 2 15 13 9 2
22 1 9 13 0 9 0 9 11 2 16 1 0 12 9 13 1 9 9 0 9 11 2
4 9 2 11 2
4 9 2 12 2
23 9 1 15 1 9 13 11 2 16 0 11 12 9 1 9 9 1 0 9 13 0 9 11
30 11 11 2 9 11 2 2 13 2 16 9 4 13 0 2 7 9 3 13 15 7 9 15 3 13 1 10 9 2 2
12 11 11 2 9 11 2 2 9 3 4 13 2
15 13 15 2 16 4 13 0 9 7 9 4 15 13 2 2
15 2 9 2 9 0 9 11 13 2 16 13 1 9 11 2
11 9 1 0 9 15 9 13 14 1 9 2
15 3 0 11 2 15 15 13 1 9 2 13 3 3 3 2
18 0 3 13 9 7 11 15 1 9 11 13 1 12 2 9 1 9 2
13 3 13 12 9 13 11 2 7 15 1 9 13 2
18 11 3 13 15 9 1 9 2 11 13 7 15 3 13 1 0 9 2
14 2 9 2 3 13 9 0 9 11 12 9 1 9 2
4 9 2 11 2
23 11 11 2 9 11 2 2 9 1 9 4 3 13 9 2 7 1 15 15 13 9 2 2
23 11 11 2 9 11 2 2 11 15 1 9 7 9 2 15 3 13 15 2 13 13 2 2
19 2 11 2 1 12 2 9 0 9 3 13 0 9 7 13 3 0 9 2
22 0 9 13 14 1 12 2 9 11 2 16 13 13 15 1 9 11 7 13 15 9 2
36 1 9 3 11 13 1 12 2 12 2 1 12 2 9 0 11 13 1 12 2 12 2 7 1 0 9 12 9 7 9 11 15 13 1 9 2
10 13 14 9 1 11 7 0 9 11 2
4 9 2 11 2
14 11 11 2 9 11 2 2 9 3 13 3 0 9 2
14 9 4 3 13 2 7 3 4 15 13 1 9 2 2
15 11 11 2 9 11 2 2 13 2 15 4 1 9 13 2
6 13 13 9 9 2 2
10 2 11 2 9 11 13 1 9 12 9
15 0 9 11 13 1 9 11 2 3 13 9 9 11 7 11
5 11 2 11 2 2
15 13 3 0 2 16 1 0 9 9 13 9 9 0 9 2
38 0 9 11 11 15 7 13 2 16 4 15 1 9 10 9 12 2 12 9 11 11 13 2 2 15 15 13 1 15 2 3 15 11 1 11 13 2 2
17 11 15 13 13 2 2 11 11 13 3 0 9 2 13 2 13 2
23 9 13 2 16 1 10 9 1 9 15 3 13 11 2 7 1 10 9 2 2 13 3 2
8 0 9 15 3 13 13 11 2
15 0 9 13 9 10 9 11 2 16 15 3 13 1 9 2
17 2 1 0 9 4 13 12 9 2 3 15 1 15 13 0 9 2
25 14 4 15 3 13 0 9 2 2 13 15 11 2 15 3 13 1 15 2 16 4 15 13 9 2
18 9 1 12 2 9 7 13 9 11 3 2 3 0 11 3 13 9 2
32 2 9 15 1 15 13 2 2 13 11 2 16 9 9 11 13 3 2 2 10 9 4 13 2 2 7 9 9 13 16 0 2
31 1 0 9 0 11 11 2 3 11 2 15 11 3 13 2 7 15 14 13 9 2 3 13 1 9 12 2 12 13 9 2
18 2 1 9 4 13 13 3 1 11 11 2 7 9 4 15 13 2 2
23 16 3 13 9 2 9 0 9 13 13 3 9 9 2 7 11 15 14 1 0 9 13 2
25 2 3 15 14 13 2 16 4 13 0 2 3 15 1 12 2 9 13 9 7 3 4 13 13 2
17 9 2 16 11 13 1 11 2 9 4 13 0 7 15 4 13 2
17 3 13 3 0 9 7 15 13 13 15 1 15 2 2 13 11 2
9 9 9 13 2 16 15 11 13 9
5 11 2 11 2 2
12 3 16 1 9 13 0 9 11 12 2 12 2
17 2 16 7 13 11 1 0 9 2 3 15 13 10 9 1 9 2
19 3 15 13 2 2 13 1 9 1 9 0 9 11 11 10 9 11 11 2
13 15 15 14 13 7 13 15 2 16 13 9 0 2
10 2 1 9 13 3 0 2 2 13 2
22 11 13 12 9 2 15 4 15 13 13 9 9 2 9 11 2 9 11 7 9 11 2
7 2 11 1 9 3 13 2
20 11 13 13 10 0 9 2 10 9 13 2 7 16 12 9 13 1 9 9 2
21 11 13 0 2 2 13 11 10 9 7 13 2 2 10 9 15 3 13 7 13 2
22 16 15 3 4 13 15 2 13 15 1 9 13 3 2 16 4 15 13 7 13 2 2
16 9 13 9 1 12 2 9 2 3 11 3 13 1 9 11 2
20 0 9 15 1 9 13 9 1 9 2 13 3 9 2 7 3 15 13 11 2
12 2 13 15 15 3 2 3 15 15 13 13 2
23 1 9 15 7 9 13 2 14 15 3 13 7 13 2 2 13 11 11 1 9 1 9 2
12 2 15 13 3 1 9 2 3 13 15 0 2
12 3 2 16 13 15 14 9 7 3 1 9 2
22 9 15 3 13 2 4 13 12 9 9 7 14 1 15 13 7 13 2 2 13 11 2
14 1 11 15 1 9 13 7 11 2 15 9 13 9 2
29 2 9 2 16 4 13 3 12 9 2 2 13 0 9 2 1 15 7 9 11 13 2 11 2 2 3 0 2 2
20 1 9 15 1 0 9 13 11 7 1 9 15 3 3 1 9 13 10 9 2
34 2 13 15 9 2 3 4 13 13 3 2 2 13 15 11 11 2 15 13 2 3 16 0 9 7 9 2 10 13 9 2 12 2 2
12 11 3 13 9 2 1 0 9 13 12 9 2
11 0 0 9 13 11 2 7 1 12 9 2
14 9 11 1 0 9 1 0 11 2 3 2 7 11 2
5 3 13 9 11 2
7 11 3 13 1 9 9 12
2 11 2
19 0 0 9 3 3 13 1 9 9 0 9 9 1 0 9 2 9 12 2
21 9 13 3 9 0 0 9 2 11 2 11 11 1 0 11 0 9 9 11 11 2
22 0 9 1 9 0 9 1 9 12 13 0 9 7 11 2 16 11 3 10 9 13 2
3 1 0 9
18 3 1 9 0 9 1 0 11 1 11 13 12 0 9 11 11 11 2
12 1 9 13 10 9 7 3 15 1 9 13 2
7 3 1 9 1 9 13 2
6 9 9 4 3 13 2
13 11 11 2 9 0 11 2 15 3 13 1 9 2
9 13 15 1 9 1 0 9 11 2
14 11 13 1 9 1 0 9 1 11 11 0 9 9 2
3 0 0 9
2 11 2
23 1 9 1 9 11 11 4 1 9 13 1 9 9 0 9 0 0 9 11 11 11 11 2
24 9 3 13 9 9 7 9 9 13 9 2 16 9 13 0 13 1 0 9 9 11 1 11 2
17 9 3 1 9 1 9 13 9 2 1 9 15 7 13 1 9 2
12 11 13 0 9 2 15 11 13 1 0 9 2
10 3 3 15 13 11 11 7 11 11 2
4 0 9 13 11
7 0 9 9 11 7 9 11
5 11 2 11 2 2
13 9 11 11 7 9 11 11 13 0 9 1 9 2
11 13 1 15 0 0 9 1 11 1 11 2
12 1 0 9 13 1 9 11 12 9 1 11 2
19 0 11 3 13 1 9 0 0 9 2 7 7 14 1 9 13 9 9 2
11 2 9 13 13 9 9 3 1 10 9 2
26 13 4 2 16 13 3 3 2 7 1 9 1 9 9 15 3 13 2 2 13 1 9 9 11 11 2
14 10 9 13 9 0 9 14 1 12 9 12 2 12 2
6 0 9 13 0 9 2
11 11 1 15 3 3 13 11 12 2 12 2
20 0 9 1 9 0 9 9 2 15 13 2 13 7 9 11 3 13 0 9 2
11 1 9 13 11 1 11 2 11 7 11 2
7 7 9 9 15 15 13 2
26 13 12 2 12 2 3 3 12 2 12 2 7 11 1 0 9 9 13 1 12 2 12 1 10 9 2
34 3 13 7 0 9 2 3 9 13 1 12 2 12 1 12 2 12 7 0 12 2 12 2 7 3 3 13 9 1 9 1 0 9 2
19 2 1 0 9 7 0 9 9 4 15 9 13 2 2 13 9 9 11 2
6 15 3 1 0 9 2
18 0 9 1 9 3 13 16 0 9 2 15 15 13 7 0 10 9 2
34 1 10 9 15 1 9 9 1 9 13 9 0 9 7 3 0 9 1 11 1 11 2 1 10 9 13 1 0 9 2 13 0 9 2
6 15 3 1 0 9 2
10 1 15 4 15 13 1 9 1 11 2
38 2 9 15 1 9 13 3 2 16 4 15 13 9 1 11 2 7 3 15 13 9 2 13 2 13 4 1 15 2 2 13 9 0 9 1 11 11 2
21 1 0 9 13 9 9 11 11 2 2 13 0 2 16 9 13 3 1 9 9 2
22 3 13 0 2 16 4 15 9 13 1 9 9 2 7 1 0 9 15 3 3 13 2
11 1 0 9 15 3 13 14 12 0 9 2
19 1 0 9 15 13 1 9 12 7 1 9 9 13 1 9 3 0 9 2
8 2 9 15 13 13 9 13 2
28 9 2 15 13 1 11 2 0 9 2 9 9 2 4 15 1 15 13 13 2 2 13 9 0 9 11 11 2
8 1 9 9 3 13 9 9 2
14 2 0 9 13 9 2 9 15 3 13 14 16 9 2
8 9 13 16 9 10 0 9 2
23 13 2 16 4 9 13 13 3 2 14 3 1 0 9 14 2 2 13 9 9 11 11 2
9 9 9 11 3 13 1 9 9 2
12 2 13 12 9 2 3 15 13 1 9 9 2
28 7 9 3 13 1 15 2 16 4 11 13 3 9 0 9 9 2 7 13 0 9 1 9 9 1 9 9 2
16 0 9 11 11 2 3 2 15 13 13 11 11 1 0 11 11
3 0 9 11
7 11 11 1 0 11 11 13
3 0 11 2
28 9 0 9 0 9 0 11 11 7 9 0 9 1 11 9 0 11 11 13 0 9 0 9 0 0 0 9 2
17 11 13 9 11 11 12 2 12 2 11 13 1 11 12 2 12 2
31 1 0 9 11 11 1 0 9 11 15 13 11 7 11 2 15 13 1 12 9 2 7 3 9 11 2 15 13 12 9 2
15 1 2 9 2 13 1 0 12 1 9 11 11 7 11 2
15 11 13 12 2 12 1 11 9 9 11 1 12 2 9 2
11 1 11 13 11 7 12 9 15 13 11 2
15 1 0 11 13 9 0 11 11 0 9 10 9 1 9 2
18 11 15 13 3 2 3 15 13 11 2 15 13 1 9 7 12 9 2
20 11 15 1 0 0 9 13 7 1 9 13 1 0 11 1 11 12 2 12 2
10 10 0 9 13 11 11 1 9 11 2
18 1 11 13 1 9 0 11 12 2 12 11 9 12 9 1 0 9 2
20 13 15 1 15 11 2 15 3 3 13 11 7 15 15 3 1 0 9 13 2
27 1 11 15 13 1 0 9 11 1 0 11 2 15 13 12 0 9 7 13 3 3 1 9 10 9 11 2
17 0 9 9 0 11 11 11 4 13 1 9 0 9 1 9 9 2
2 11 11
5 11 13 0 9 9
14 9 11 1 9 1 9 14 13 1 9 1 11 14 0
9 11 2 11 2 11 2 11 2 2
43 0 9 11 2 11 2 12 2 12 2 13 3 0 1 12 9 2 7 1 12 2 9 13 3 1 11 12 9 7 13 1 12 2 9 2 15 3 13 9 1 9 14 2
26 11 13 9 3 7 12 1 0 9 9 13 13 3 12 2 9 2 3 0 9 11 11 13 0 9 2
35 2 1 9 15 13 1 12 9 0 7 1 15 13 0 2 16 15 1 10 9 13 0 9 9 11 2 2 13 9 9 0 9 11 11 2
33 1 0 12 13 0 3 0 9 12 9 7 1 15 2 16 15 9 13 14 9 9 2 13 1 9 13 1 9 9 1 0 9 2
14 2 10 9 1 9 1 9 14 13 3 1 15 0 2
21 3 13 13 1 11 7 3 7 3 1 11 2 3 3 4 13 13 1 9 11 2
12 12 9 15 3 4 13 2 2 13 11 11 2
9 3 9 0 9 13 3 14 0 2
11 2 3 13 13 2 16 13 13 0 9 2
35 0 9 13 9 2 7 3 13 3 2 7 16 1 10 9 4 1 9 12 2 12 3 13 2 16 9 13 2 2 13 0 9 11 11 2
19 10 9 13 0 12 9 3 2 7 1 11 2 1 11 7 1 11 13 2
12 3 0 13 3 9 1 11 7 3 1 11 2
25 7 1 0 9 9 4 15 9 1 9 14 13 13 14 0 9 0 9 7 11 1 0 12 9 2
41 3 0 9 2 12 2 1 9 2 15 1 9 3 13 1 9 9 2 16 3 13 12 2 12 1 11 7 13 15 3 10 0 9 1 9 2 1 15 13 3 2
10 1 10 0 9 13 7 14 0 9 2
27 2 16 13 10 9 2 16 13 11 2 11 7 11 2 13 13 2 2 13 15 1 9 0 9 11 11 2
34 10 9 2 15 1 9 9 13 10 9 9 2 13 0 9 2 3 13 1 0 0 9 7 1 9 13 0 9 9 3 1 0 11 2
8 11 13 1 11 1 9 14 9
5 11 2 11 2 2
20 1 9 9 1 9 0 9 13 0 9 1 9 11 11 11 10 0 0 9 2
31 0 9 0 12 9 1 9 0 0 9 3 13 1 9 10 9 12 2 12 7 3 15 13 10 9 1 9 1 9 14 2
28 2 1 12 9 4 1 9 3 3 13 2 2 13 0 9 11 1 9 2 1 15 15 9 10 0 9 13 2
11 2 11 1 15 13 2 7 7 13 3 2
21 15 4 15 15 13 2 7 7 15 1 9 3 13 2 2 13 9 9 11 11 2
26 15 2 16 4 9 0 1 9 14 13 13 3 14 0 9 2 13 7 9 11 2 2 15 13 0 2
11 1 11 4 13 0 9 2 7 13 4 2
7 1 11 15 13 3 3 2
12 3 15 1 10 0 9 13 9 3 3 2 2
19 15 15 13 0 7 9 11 11 11 2 2 3 1 11 15 13 0 9 2
12 13 4 3 0 7 1 15 10 9 3 13 2
11 13 15 2 16 13 1 9 14 9 2 2
23 11 7 11 15 3 13 2 16 4 15 13 13 3 15 2 15 13 10 9 1 9 14 2
21 2 1 11 13 7 0 9 2 7 15 2 15 13 1 10 0 9 9 14 3 2
41 13 9 7 7 1 0 9 13 1 9 3 15 1 11 2 2 13 11 2 15 9 3 13 7 9 11 2 2 0 9 4 3 13 2 7 13 3 0 0 9 2
16 13 0 9 7 1 10 9 15 14 3 3 13 1 9 2 2
3 9 9 9
41 0 2 11 2 11 2 12 2 12 2 2 11 11 2 9 0 2 11 2 2 13 15 0 9 2 1 0 12 4 3 13 9 2 7 3 4 13 0 9 2 2
21 11 11 2 9 11 2 2 13 15 12 0 9 2 15 13 10 9 1 0 9 2
8 15 4 13 3 7 3 2 2
33 11 2 11 2 12 2 12 2 2 11 11 2 9 11 2 2 1 9 9 4 13 9 3 2 16 16 4 15 15 13 15 13 2
16 1 12 2 9 4 3 13 7 13 13 9 2 15 13 2 2
21 11 11 2 9 11 2 2 1 9 9 4 13 2 16 12 9 13 9 14 0 2
8 13 10 0 9 7 9 2 2
22 11 2 11 2 12 2 12 2 2 11 11 2 9 11 2 2 13 4 9 0 9 2
14 13 3 1 9 2 7 13 2 16 15 15 13 2 2
15 11 11 2 9 11 2 2 15 3 13 2 13 13 0 2
16 13 15 9 0 9 2 1 9 0 9 4 13 9 1 9 2
24 13 4 2 16 16 1 9 13 14 12 9 2 9 11 2 13 4 15 1 10 9 3 12 2
16 13 15 3 9 11 11 7 1 9 11 2 11 7 11 2 2
6 1 0 9 9 3 11
26 1 0 9 0 9 13 1 9 2 15 13 1 0 9 2 0 9 13 1 0 9 0 9 11 11 2
46 1 0 9 13 0 2 1 15 13 1 12 2 9 11 11 2 11 2 2 1 12 2 11 11 2 11 2 2 1 12 2 11 11 1 11 7 1 12 2 9 9 0 11 11 11 2
29 1 9 0 1 9 13 0 9 0 9 11 11 11 2 11 11 1 11 2 2 15 13 1 0 2 0 9 0 2
16 1 0 9 13 1 0 9 3 0 2 15 3 13 0 9 2
3 2 11 2
8 11 13 9 2 16 1 9 13
2 11 2
28 11 2 15 3 1 0 9 13 10 0 9 1 0 9 1 9 1 9 2 13 1 9 1 11 10 0 9 2
28 1 9 1 9 1 9 9 2 12 13 1 12 9 3 3 2 7 16 1 0 9 1 9 13 2 3 13 2
14 11 13 0 9 7 1 0 12 9 13 12 0 9 2
9 2 13 0 9 2 3 4 13 2
7 13 4 15 0 0 9 2
7 13 4 15 1 15 3 2
33 9 2 16 1 0 9 15 9 1 9 3 13 2 13 4 13 3 3 2 2 13 11 2 15 15 1 0 9 3 13 1 9 2
10 1 0 9 13 11 2 9 9 2 2
22 13 0 7 13 9 9 12 9 2 1 0 12 9 3 2 16 0 0 2 11 11 2
10 1 0 9 13 11 1 9 12 9 2
11 0 9 15 7 13 1 9 7 13 15 2
11 7 0 0 9 15 7 1 0 9 13 2
20 11 11 2 9 0 9 2 2 1 9 13 3 0 2 3 16 15 13 11 2
12 13 12 9 1 12 0 2 7 15 13 0 2
24 9 0 13 2 9 1 9 13 0 2 1 0 9 13 9 2 16 15 13 1 0 9 2 2
16 1 0 9 1 9 13 9 0 9 1 9 1 0 12 9 2
21 9 0 0 0 9 13 1 9 9 9 11 2 15 1 9 13 0 9 11 1 11
3 11 16 0
7 9 13 0 9 9 1 11
5 0 11 2 11 2
16 11 11 13 1 0 11 1 0 9 0 11 9 0 9 9 2
30 13 15 0 9 0 9 2 15 1 12 9 3 13 1 9 7 10 9 13 1 0 9 2 1 10 9 1 0 9 2
10 0 9 13 11 1 11 7 11 11 2
16 11 11 13 3 1 0 9 1 0 9 0 9 9 1 11 2
22 13 15 10 0 0 9 2 1 9 13 1 0 9 9 1 0 9 1 11 2 11 2
19 3 16 1 11 1 9 13 9 1 11 1 0 9 13 0 0 9 9 2
17 13 7 9 2 16 15 13 3 2 15 4 13 0 9 0 9 2
11 0 9 13 11 11 2 9 0 0 9 2
2 9 9
2 11 2
22 1 0 9 9 9 1 11 13 0 9 0 9 2 16 1 9 13 11 12 2 12 2
3 9 0 9
3 9 11 2
35 11 11 2 11 2 9 0 9 1 9 11 2 15 3 13 9 0 9 11 1 9 12 1 11 11 11 2 16 15 13 1 9 10 9 2
27 11 15 10 9 1 9 1 11 13 2 16 13 9 9 9 2 7 11 15 1 9 13 0 9 1 9 2
10 11 15 13 1 9 9 1 0 9 2
20 11 2 11 2 15 11 13 12 9 2 1 10 9 13 2 7 13 15 9 2
17 10 9 13 2 7 13 9 9 2 16 15 9 1 0 9 13 2
11 3 13 9 2 16 11 13 10 9 3 2
15 2 13 15 0 9 2 15 4 1 9 13 2 2 13 2
28 9 3 13 0 0 9 2 16 4 11 13 7 9 11 13 1 0 9 1 9 2 15 15 13 1 12 9 2
12 0 11 4 13 1 0 9 1 9 15 9 2
17 3 13 0 0 9 1 9 0 9 9 1 9 11 0 0 9 2
17 9 15 13 0 9 11 2 15 13 0 2 9 2 1 0 9 2
19 0 11 11 4 1 9 1 9 13 7 9 13 9 9 9 1 0 9 2
4 0 9 1 11
6 11 15 13 16 0 9
5 9 1 9 13 15
5 11 2 11 2 2
29 12 9 1 9 1 9 2 0 9 1 12 9 9 7 12 9 9 1 9 11 13 9 0 9 11 9 1 11 2
41 0 9 1 0 9 13 1 12 9 9 12 0 9 7 11 11 13 1 9 3 16 9 9 0 2 1 10 9 13 1 0 9 2 2 15 13 3 9 12 9 2
24 9 1 0 9 9 13 9 12 9 11 11 7 16 0 9 15 13 1 0 9 13 0 12 2
14 0 9 15 15 13 1 9 12 9 0 9 11 13 2
25 9 1 12 1 0 0 9 0 9 2 10 9 13 1 0 9 0 9 2 3 13 1 0 9 2
27 3 10 9 13 1 0 9 3 3 0 9 1 12 2 2 2 9 2 1 0 9 15 1 9 13 12 2
21 2 3 4 13 2 16 4 15 13 2 16 4 13 1 0 9 1 11 3 0 2
15 3 1 9 4 13 2 16 4 13 13 2 3 13 12 2
6 3 3 13 3 0 2
24 13 4 15 2 16 16 13 9 2 3 15 3 3 13 9 2 7 3 3 13 12 9 13 2
42 13 2 16 1 9 1 11 13 1 11 0 0 9 1 0 9 2 16 4 15 15 1 9 3 3 3 13 2 2 13 9 2 1 15 13 9 0 9 1 0 9 2
48 0 9 2 12 9 2 13 3 9 11 2 15 1 0 9 13 0 9 0 9 2 2 9 4 3 13 7 9 1 9 13 2 7 16 4 13 3 0 2 16 4 13 1 0 9 3 3 2
12 0 7 13 2 16 4 13 1 9 14 12 2
17 13 4 15 1 0 9 7 13 7 13 4 15 16 0 9 2 2
36 9 10 0 9 13 0 13 0 11 11 2 9 0 9 1 12 9 9 2 2 13 14 2 16 4 1 12 3 13 1 9 0 9 11 2 2
20 1 9 13 0 9 12 9 7 13 0 2 16 13 14 12 12 1 10 9 2
28 1 0 9 9 11 11 2 15 15 3 16 12 1 0 13 0 9 9 1 9 2 15 3 3 13 0 9 2
39 1 9 1 9 7 1 9 13 9 7 0 9 13 9 9 2 2 9 1 9 13 9 2 14 1 9 4 13 9 1 0 9 7 0 9 1 9 2 2
11 0 9 13 9 7 12 13 9 1 9 2
17 0 11 15 13 1 12 7 13 1 12 9 0 11 2 12 2 2
15 2 14 4 13 9 2 3 15 0 12 9 13 0 9 2
53 9 13 3 9 1 0 9 2 1 15 15 13 3 3 2 7 1 15 2 3 15 9 11 13 1 9 1 11 2 2 13 9 11 2 10 9 2 3 16 11 2 13 0 9 1 0 9 1 12 5 12 9 2
9 0 9 15 13 1 9 0 9 2
51 1 9 13 9 1 12 9 7 1 0 9 12 9 7 0 9 2 16 13 12 0 9 2 2 13 4 15 2 16 13 9 2 7 3 15 9 11 13 2 16 13 9 1 9 2 7 16 15 13 2 2
5 9 11 2 9 11
2 11 2
28 1 9 1 9 1 0 9 1 0 11 13 11 11 11 0 9 1 9 1 12 9 9 12 9 1 12 0 2
10 11 13 1 9 7 9 1 0 9 2
9 11 11 13 1 0 9 12 9 2
22 1 0 9 15 1 12 9 13 14 12 12 9 1 9 7 1 0 9 13 0 9 2
16 0 0 9 13 3 11 11 1 9 1 0 9 9 12 9 2
13 1 9 9 13 0 9 0 9 1 11 7 11 2
2 11 13
2 11 2
11 1 0 9 13 0 0 9 12 0 9 2
14 13 15 0 9 0 9 1 9 12 1 11 11 11 2
17 3 13 2 16 0 9 0 9 1 11 13 1 12 1 12 3 2
17 9 0 0 9 13 9 2 16 0 9 13 0 9 9 1 9 2
12 1 12 1 0 9 13 9 0 0 9 11 2
7 11 2 11 13 1 9 9
3 0 11 2
37 1 9 0 12 0 9 0 11 11 2 11 4 13 0 9 11 2 11 2 15 13 9 11 1 11 2 7 7 1 15 0 13 3 12 2 12 2
39 3 13 9 0 9 11 11 13 2 2 13 15 0 2 9 13 12 0 9 9 2 3 3 13 1 11 2 11 7 15 15 10 9 13 13 2 2 13 2
13 11 3 13 1 11 7 11 2 15 13 9 9 2
18 9 11 11 11 13 11 2 11 9 9 1 12 9 7 9 12 9 2
4 11 3 1 11
5 11 2 11 2 2
33 1 0 0 9 2 9 1 9 9 2 13 1 0 9 0 9 0 9 11 11 11 2 15 3 13 0 9 14 1 9 12 9 2
31 3 13 0 9 3 1 9 2 7 3 1 15 13 9 11 11 11 11 2 16 15 1 0 9 1 11 13 13 12 9 2
39 15 15 15 3 13 2 7 16 1 0 9 1 15 13 3 2 7 3 13 0 9 1 0 9 9 12 11 11 11 2 15 3 1 11 13 1 9 3 2
22 3 1 0 9 13 3 0 9 12 2 15 1 10 9 13 0 9 0 0 0 9 2
44 2 15 12 13 1 9 2 16 4 15 10 9 13 1 9 1 0 9 2 15 13 2 2 13 1 9 9 2 15 3 2 16 15 13 13 9 2 13 0 9 1 0 9 2
40 10 0 9 13 3 13 1 9 9 1 11 2 2 3 15 15 13 2 7 3 1 0 9 13 0 9 16 0 9 1 9 0 9 2 16 3 1 15 13 2
23 3 15 3 13 3 13 2 16 16 13 9 9 2 13 1 9 13 1 9 1 12 2 2
13 1 12 9 13 11 1 11 1 0 9 11 11 2
14 2 13 3 0 9 2 7 16 13 3 0 16 15 2
14 9 15 1 9 13 3 2 16 13 0 9 1 9 2
42 1 10 9 3 13 3 3 1 0 9 2 2 13 9 9 11 11 2 15 15 13 2 16 9 1 0 9 13 3 3 7 3 1 12 9 15 4 13 1 12 9 2
25 1 9 15 13 11 11 13 2 14 16 13 10 9 1 11 2 2 3 4 13 1 9 11 9 2
18 13 4 3 11 2 7 13 15 2 16 4 15 13 13 0 9 9 2
10 0 13 3 2 7 15 13 9 2 2
4 9 11 13 9
2 11 2
33 0 0 9 9 1 11 1 9 12 9 11 13 9 9 2 16 0 9 9 1 11 11 13 7 1 0 9 1 0 15 13 9 2
30 0 9 13 1 0 7 0 9 3 12 2 12 2 3 13 11 3 9 13 2 7 13 15 2 1 0 9 3 13 2
25 1 0 9 13 1 12 2 12 7 3 1 12 2 12 2 7 11 0 9 13 9 1 10 9 2
5 0 9 1 11 11
25 0 9 15 13 0 9 1 9 11 11 1 9 11 11 9 0 9 2 0 9 1 11 11 2 2
32 13 12 9 1 9 12 2 12 0 9 0 9 2 9 2 2 15 9 12 13 0 9 7 9 11 11 2 12 2 12 2 2
13 0 9 11 11 13 3 10 9 0 9 7 9 2
22 10 9 15 11 13 3 14 9 2 7 7 9 2 1 15 1 0 9 13 10 9 2
24 9 0 9 9 11 11 15 1 9 1 9 13 1 0 1 9 11 2 11 7 11 2 11 2
11 13 15 3 1 9 0 9 1 9 0 2
26 9 0 9 9 0 9 15 13 9 0 7 0 9 9 2 9 0 9 7 11 11 11 7 11 11 2
3 2 11 2
3 9 1 9
17 9 2 0 9 3 13 15 2 15 13 1 9 3 14 0 9 2
9 13 9 9 7 0 9 0 9 2
20 3 1 0 0 0 9 9 9 13 9 7 1 0 9 13 0 9 2 2 2
34 1 9 15 15 3 3 13 2 1 12 9 1 9 11 11 0 9 1 9 2 3 9 13 1 9 15 7 11 11 13 9 9 0 2
16 1 0 9 9 11 11 15 7 11 11 3 13 1 0 9 2
24 13 15 15 15 1 9 9 11 11 2 15 15 3 13 0 9 1 10 9 2 3 0 9 2
28 9 13 3 13 2 16 9 9 13 2 1 0 0 9 7 9 2 15 15 13 13 1 9 2 13 0 9 2
6 7 13 15 9 13 2
24 3 9 0 9 2 15 13 10 0 9 13 7 13 15 1 15 2 13 9 9 0 9 9 2
36 0 9 15 14 13 2 16 3 13 1 0 9 2 0 9 11 2 1 0 3 0 0 2 9 11 7 1 3 0 0 9 1 9 11 11 2
15 0 9 9 9 0 9 11 11 13 0 0 9 0 9 2
21 15 15 1 0 9 2 7 3 3 2 1 0 9 13 1 9 0 9 1 9 2
18 11 11 1 0 9 13 7 9 0 16 15 0 9 1 11 11 3 2
17 2 3 2 0 2 11 2 3 13 12 1 0 0 9 15 9 2
32 0 9 10 0 9 1 9 3 13 7 3 0 11 1 11 2 15 1 0 9 3 13 3 0 2 0 9 1 0 0 9 2
27 0 0 9 9 11 11 2 1 9 11 2 13 3 9 0 0 9 1 9 10 0 7 0 9 2 2 2
23 0 1 0 9 0 9 1 9 0 7 0 9 13 9 0 9 1 9 2 15 13 9 2
24 13 0 9 0 9 9 1 0 9 2 3 3 0 9 3 13 1 9 10 0 9 13 9 2
9 7 14 3 2 16 15 3 13 2
27 13 2 16 3 9 9 2 15 1 0 9 13 1 3 0 9 11 7 11 2 15 10 9 13 2 2 2
6 9 2 11 2 12 2
8 9 1 11 2 11 2 11 2
14 13 2 11 11 2 11 11 2 11 1 11 7 0 2
5 9 12 2 9 2
4 0 9 0 9
26 9 3 0 9 9 0 9 12 1 0 9 0 9 7 9 4 13 12 2 9 3 1 0 0 9 2
19 1 9 13 12 12 0 9 7 9 2 3 9 9 9 2 15 9 13 2
13 12 1 9 13 7 0 9 2 0 3 1 11 2
10 9 3 13 1 12 9 3 16 3 2
14 1 9 9 11 11 15 3 3 13 9 9 3 0 2
12 0 9 4 1 0 13 1 0 7 0 9 2
17 1 12 9 4 13 3 16 12 0 9 1 9 0 1 10 9 2
10 0 9 13 9 0 9 0 0 9 2
17 1 11 13 1 9 1 9 2 16 1 0 9 4 0 9 13 2
10 2 15 15 7 13 2 2 13 11 2
15 9 13 3 3 13 1 9 7 13 1 0 9 0 9 2
9 10 0 9 7 9 3 13 9 2
24 2 13 1 15 2 16 4 10 9 13 0 2 7 7 3 15 13 9 9 2 2 13 11 2
32 2 9 9 13 13 1 0 0 9 2 2 13 7 13 2 16 0 9 0 11 11 11 13 9 11 1 9 0 9 10 9 2
22 9 0 9 9 9 13 7 9 1 9 1 0 9 2 15 13 0 9 1 0 9 2
16 9 1 0 9 13 9 0 9 0 11 0 1 9 11 11 2
20 10 9 0 15 9 0 9 13 0 9 3 1 9 1 0 9 1 9 12 2
13 0 0 9 1 9 3 13 9 9 7 9 9 2
22 2 13 7 1 9 1 3 0 7 0 9 2 2 13 9 9 9 0 9 11 11 2
18 1 9 0 9 15 1 10 9 13 13 0 9 11 7 10 0 9 2
35 11 11 1 11 2 12 1 0 9 0 9 9 9 2 9 7 9 0 2 12 2 12 2 2 13 1 9 11 11 1 10 0 1 11 2
35 9 11 13 0 9 9 10 0 9 11 11 2 12 2 12 2 2 15 1 0 9 13 1 0 12 9 13 0 11 1 0 9 11 11 2
16 1 9 9 13 3 9 9 10 0 9 7 9 0 9 0 2
5 2 11 2 9 11
3 9 1 9
33 9 2 9 2 9 2 9 2 0 9 2 9 2 9 1 9 2 0 2 3 15 13 9 2 9 13 0 2 13 9 2 2 2
20 0 9 0 9 1 9 1 10 0 9 2 9 9 1 10 0 9 2 2 2
28 7 15 13 13 0 2 3 3 0 9 9 11 11 2 0 9 2 7 13 14 13 15 3 9 9 2 2 2
17 11 13 1 10 3 0 9 3 9 0 9 2 7 1 11 11 2
14 12 3 13 0 9 2 12 15 13 1 9 0 9 2
11 3 10 9 15 10 3 0 9 3 13 2
6 7 3 13 3 9 2
12 0 9 3 3 13 9 2 16 4 13 3 2
16 13 0 9 2 16 4 1 15 0 2 3 3 1 0 9 2
22 9 13 3 1 9 9 9 2 7 7 10 0 9 15 13 1 9 14 1 0 9 2
24 9 3 2 2 2 15 3 11 13 2 0 9 2 14 1 9 12 2 3 9 1 11 2 2
17 13 15 9 2 16 11 3 13 1 10 0 9 3 10 0 9 2
15 3 4 3 13 2 16 0 0 9 3 13 1 9 0 2
8 3 9 1 0 9 3 13 2
23 1 9 1 3 2 2 2 1 15 3 7 3 0 9 13 7 1 9 3 13 14 9 2
9 16 16 4 15 11 13 2 2 2
29 3 16 3 2 7 3 15 9 15 13 15 2 1 9 7 9 1 9 7 0 9 1 0 9 14 1 0 9 2
9 2 3 1 9 15 13 9 2 2
9 0 9 16 4 3 13 0 9 2
30 7 16 4 15 13 9 2 16 0 0 9 15 9 13 7 3 2 9 9 9 13 9 0 9 7 9 0 0 9 2
13 15 13 13 2 16 11 15 0 9 10 9 13 2
21 9 1 0 9 1 15 13 0 9 2 3 9 3 13 9 1 9 10 10 9 2
27 1 10 0 9 13 11 0 9 2 7 1 9 15 3 13 10 9 2 1 15 3 10 0 9 11 11 2
18 13 7 2 16 1 15 10 0 9 1 9 13 9 11 11 3 3 2
7 3 15 2 6 2 13 2
5 11 13 9 0 9
27 1 12 2 9 9 0 9 0 9 2 15 13 1 9 1 11 1 11 2 13 0 9 11 11 1 11 2
22 1 12 0 9 1 12 9 13 9 0 9 10 0 9 1 9 13 0 9 0 9 2
11 0 7 0 9 13 9 1 11 1 11 2
11 1 9 9 13 10 9 9 0 0 9 2
31 1 11 11 1 0 9 9 7 9 2 15 13 12 1 9 2 15 0 9 13 1 9 0 9 2 0 9 7 9 9 2
5 15 2 3 2 3
12 11 11 13 3 1 9 9 11 9 0 9 2
6 13 1 12 2 9 2
37 9 9 0 9 11 11 0 9 2 9 2 9 0 2 9 2 13 11 2 13 3 2 1 12 9 2 2 1 0 9 1 9 1 9 0 9 2
30 9 11 11 7 9 11 11 4 1 0 9 2 0 12 2 11 12 2 3 1 12 9 13 10 9 13 0 2 2 2
4 13 15 11 9
32 1 9 1 0 12 2 9 0 9 3 0 7 0 9 2 0 9 7 9 11 9 11 15 3 13 12 0 7 12 0 9 2
35 0 9 1 15 1 0 9 13 12 9 2 15 15 4 1 9 12 2 7 12 2 9 13 1 9 9 9 11 7 0 9 1 0 9 2
31 1 9 0 3 0 9 15 3 1 11 13 7 9 9 1 11 2 11 2 11 2 11 2 11 2 11 2 11 7 11 2
21 1 0 9 9 0 9 7 3 13 9 9 0 9 1 0 7 0 9 9 9 2
4 15 4 3 13
4 12 13 3 2
10 0 9 13 1 0 0 9 1 11 2
8 11 11 2 9 0 9 0 9
15 9 11 13 1 9 12 1 10 11 9 3 3 0 9 2
43 11 7 11 3 13 2 16 11 2 15 3 13 1 10 2 0 2 9 2 13 1 0 9 2 10 0 9 3 9 13 2 7 1 0 9 2 15 3 13 9 0 9 2
17 1 0 2 9 2 7 1 0 9 15 7 1 12 9 13 9 2
4 0 9 0 11
22 13 15 2 16 15 9 0 9 13 1 0 9 2 2 3 14 13 13 2 11 2 2
13 9 0 9 11 11 13 0 2 2 3 3 2 2
5 0 9 0 11 9
10 9 0 9 13 16 9 9 1 9 2
8 1 10 9 15 15 15 13 2
16 3 4 15 10 2 0 2 9 13 13 7 1 0 0 9 2
4 0 0 0 9
17 15 4 15 13 2 16 4 1 9 4 13 11 2 7 0 9 2
16 9 4 3 13 9 2 3 4 7 0 9 11 13 0 9 2
7 0 9 9 13 1 9 2
6 0 0 9 9 11 11
4 11 13 9 2
8 0 9 13 10 9 1 9 2
7 7 13 9 15 1 9 2
5 3 15 15 13 2
9 0 9 7 0 9 1 9 11 11
5 2 13 15 2 2
7 9 2 2 13 15 2 2
4 11 15 13 2
11 3 2 3 13 0 9 2 13 0 9 2
11 1 9 15 13 9 2 2 13 15 2 2
8 1 9 1 9 0 9 1 11
18 16 15 3 4 13 1 15 2 13 1 11 7 13 15 3 1 9 2
7 9 0 9 2 0 1 11
4 13 0 9 2
9 13 3 13 1 15 2 13 9 2
5 13 3 10 9 2
9 0 9 11 11 2 2 12 9 2
17 13 0 2 16 10 9 13 13 9 10 9 2 16 4 13 13 2
19 9 3 9 13 7 13 1 0 9 7 3 13 1 15 3 3 16 3 2
20 9 11 11 1 9 9 11 0 0 11 1 0 9 9 0 9 1 9 1 11
9 13 0 9 9 2 7 13 9 2
8 11 11 1 9 0 0 11 11
3 11 3 9
27 13 15 9 2 13 15 3 7 13 0 9 9 9 11 1 0 9 1 0 9 1 0 9 12 0 9 2
12 2 1 10 9 13 9 11 11 2 2 13 2
11 9 0 9 13 1 9 0 11 9 9 2
13 13 9 9 12 2 10 9 1 9 9 0 9 2
17 10 9 15 13 1 11 7 1 9 13 13 10 9 2 3 13 2
8 2 13 9 13 10 9 11 2
6 15 3 13 9 9 2
19 13 4 2 16 13 3 3 13 9 1 0 9 1 9 0 2 2 13 2
24 3 15 3 1 0 9 11 13 9 11 2 9 0 1 9 0 9 1 9 11 11 12 2 2
11 1 9 12 3 13 9 11 10 0 9 2
16 0 9 1 15 13 1 9 12 14 1 0 9 1 0 9 2
5 9 13 1 9 2
14 2 13 9 14 0 13 2 3 4 15 7 15 13 2
24 9 13 3 0 2 14 2 2 13 9 9 7 13 9 3 1 9 1 9 1 12 9 9 2
10 0 9 15 1 9 13 9 9 13 2
6 1 10 9 13 9 2
20 14 9 9 1 12 2 9 7 9 0 0 9 11 11 3 13 9 3 0 2
19 1 9 13 1 9 0 0 9 2 0 9 9 2 1 9 3 0 9 2
12 0 9 3 13 0 0 0 9 7 9 9 2
21 2 15 13 0 2 16 4 13 3 2 16 4 3 3 13 9 7 14 10 9 2
7 7 3 1 15 3 13 2
21 9 3 13 2 2 13 11 2 9 1 9 2 9 2 2 7 13 3 1 9 2
16 9 12 2 9 15 13 0 9 13 0 9 1 0 9 9 2
24 1 10 9 15 15 1 9 9 9 7 9 9 1 9 9 13 13 1 9 9 0 0 9 2
10 1 10 9 13 13 0 9 0 9 2
10 1 9 9 15 0 9 9 13 13 2
9 7 7 3 13 2 13 0 9 2
4 2 1 9 2
37 9 7 9 13 1 9 2 2 13 3 9 1 0 9 7 13 9 0 9 1 0 9 9 1 0 9 7 0 9 2 0 9 1 0 9 9 2
32 0 9 0 11 13 1 9 1 9 0 9 9 2 15 13 0 13 1 12 9 2 9 0 2 9 0 9 1 9 12 2 2
15 13 0 9 2 12 9 9 0 9 2 12 9 9 2 2
7 2 15 3 13 0 9 2
20 3 15 3 2 3 16 11 2 13 2 2 13 0 9 9 1 0 0 9 2
26 1 9 9 15 3 1 10 9 1 0 9 0 0 9 13 3 7 13 9 1 9 3 0 0 9 2
18 3 13 1 9 3 0 9 11 11 1 0 0 9 1 9 0 9 2
18 2 13 15 15 2 13 15 9 2 2 13 15 0 9 12 1 0 2
19 2 13 2 16 15 15 11 13 2 16 15 13 0 2 16 15 3 13 2
13 7 11 13 14 11 2 11 13 14 9 1 11 2
17 4 15 13 3 2 7 7 1 11 4 3 13 16 1 0 9 2
12 13 15 2 13 2 2 13 7 13 1 9 2
29 1 0 9 2 15 4 1 9 9 11 13 11 7 11 2 4 3 13 0 9 2 0 15 1 11 7 0 9 2
21 1 10 9 13 1 9 14 9 9 9 2 0 9 0 9 2 9 2 0 9 2
27 2 0 9 1 15 7 0 9 1 15 2 2 13 3 7 3 1 9 1 9 2 3 3 13 9 9 2
27 2 9 15 13 2 9 15 13 2 2 13 3 0 9 1 0 9 2 13 0 15 9 7 13 0 9 2
10 13 4 1 0 9 0 9 10 9 2
12 2 0 0 9 2 2 13 7 13 15 3 2
21 2 13 0 9 2 0 9 2 2 13 1 0 2 13 9 7 13 0 9 9 2
3 9 13 2
7 2 3 13 0 3 15 2
20 11 13 0 9 9 11 1 11 11 1 11 2 3 9 0 9 11 11 11 2
25 1 9 1 15 2 16 11 0 9 3 1 9 1 9 1 9 13 2 11 10 9 13 1 9 2
15 1 9 10 9 13 0 9 3 1 11 16 1 0 9 2
9 13 15 2 16 13 10 9 0 2
14 9 1 0 9 7 1 0 9 13 12 3 0 9 2
11 9 9 10 9 13 13 2 16 13 3 2
12 9 11 4 15 13 13 3 16 9 0 9 2
14 9 0 9 1 11 13 1 0 7 0 9 3 0 2
15 10 9 4 13 0 9 13 2 16 4 15 13 9 9 2
3 1 9 2
17 9 1 9 9 9 0 11 1 9 1 9 10 9 3 3 13 2
17 3 7 13 0 3 15 2 7 15 2 16 15 11 3 4 13 2
21 1 0 9 2 15 9 13 1 9 15 0 9 2 13 13 9 9 9 1 9 2
11 1 10 9 13 7 10 9 3 15 0 2
15 13 2 16 1 9 10 9 13 13 10 9 1 9 3 2
18 9 9 1 9 4 3 13 1 15 2 16 0 9 1 9 15 13 2
10 13 4 13 2 10 9 10 9 13 2
24 1 9 9 1 9 4 15 13 13 9 7 9 9 9 9 0 7 0 11 1 9 9 11 2
11 1 15 4 13 9 10 9 1 9 0 2
18 13 2 16 9 11 2 16 15 13 7 3 2 4 13 1 9 11 2
5 13 2 16 14 2
20 11 13 7 3 0 7 0 9 2 16 1 15 9 4 13 1 10 9 13 2
5 11 1 9 0 9
52 2 3 0 9 1 0 11 2 16 13 3 3 1 9 2 15 12 12 4 13 11 2 15 13 1 9 9 2 2 13 3 9 11 2 15 13 1 9 11 2 9 11 2 7 10 9 11 1 9 12 13 2
21 9 11 1 9 11 11 13 2 16 11 3 12 9 13 1 9 2 9 7 9 2
19 9 0 9 11 2 15 4 13 1 10 9 1 9 12 2 13 9 9 2
19 7 9 0 9 15 11 3 13 1 9 9 9 2 15 13 12 2 9 2
31 2 16 9 13 2 13 0 9 16 9 2 16 4 13 9 10 0 9 2 16 1 11 13 0 9 2 2 13 9 11 2
26 2 15 0 3 4 13 7 13 15 3 2 16 10 9 13 0 13 3 2 7 14 1 12 9 2 2
37 2 3 4 13 1 9 1 0 9 2 16 15 3 13 1 9 10 0 9 1 9 9 2 2 13 10 0 9 2 10 0 9 13 13 0 9 2
30 9 11 13 3 3 1 9 1 11 2 1 10 9 13 0 9 7 10 9 7 9 13 3 0 9 0 1 0 9 2
56 9 11 11 1 10 9 13 9 9 13 0 9 10 9 2 0 0 9 2 7 0 9 9 2 15 13 3 0 7 13 15 3 3 13 1 10 9 2 13 11 11 11 2 15 13 1 0 2 2 0 9 1 9 0 9 2
38 2 13 2 16 13 0 9 16 9 2 2 13 7 13 2 16 0 13 1 15 2 16 15 4 13 3 13 1 9 2 7 13 0 15 1 9 13 2
19 1 0 2 0 9 13 14 1 0 9 1 12 9 7 12 0 4 13 2
7 1 15 13 3 12 9 2
40 2 9 1 11 13 14 9 11 2 16 15 13 7 13 7 13 1 15 9 2 16 13 0 2 7 15 15 13 1 9 13 2 2 13 0 9 9 11 11 2
20 11 2 3 13 0 9 1 11 2 16 4 15 13 13 2 16 3 13 9 2
26 10 9 13 3 7 3 3 2 16 13 15 1 15 2 16 4 13 9 11 1 11 2 2 13 11 2
26 9 7 0 11 2 13 0 9 2 7 15 9 1 9 0 11 2 2 13 0 11 11 2 9 9 2
21 2 14 14 15 13 2 7 13 2 16 15 4 13 1 15 2 15 15 13 2 2
14 12 9 1 9 9 9 13 1 11 13 10 9 9 2
11 10 9 13 1 9 1 0 9 1 9 2
1 3
25 11 3 13 9 1 11 2 15 4 13 1 9 3 2 16 4 1 0 9 13 12 1 10 9 2
31 0 9 2 1 15 4 13 9 11 2 12 1 0 9 1 9 2 4 13 1 9 1 0 9 0 9 11 11 1 11 2
13 11 4 13 1 0 9 1 11 7 1 9 11 2
19 13 15 1 11 0 0 0 9 1 9 0 9 9 0 9 9 11 11 2
23 11 13 0 9 11 1 9 0 0 9 7 13 15 1 9 9 0 0 0 9 1 11 2
37 9 0 9 0 9 2 11 2 11 11 2 12 2 4 1 9 13 0 0 9 1 9 12 9 7 9 0 9 1 9 1 9 9 1 0 11 2
21 11 15 13 15 2 16 15 13 10 0 9 0 9 7 16 13 11 3 3 13 2
26 11 11 1 10 9 1 11 13 2 9 13 9 0 1 11 2 0 9 1 9 1 11 1 9 12 2
18 13 3 11 11 2 16 4 15 13 1 9 13 2 9 1 9 2 2
18 11 13 0 9 9 7 9 2 16 4 15 13 1 9 1 0 9 2
24 9 0 11 7 11 13 3 1 11 0 9 2 15 13 13 9 1 9 1 9 0 0 9 2
29 9 13 9 9 2 15 4 13 1 9 0 9 7 1 9 0 9 2 0 1 0 0 9 1 9 1 12 9 2
27 0 0 9 13 2 16 13 1 9 11 2 15 13 1 0 9 0 9 13 0 9 0 9 3 12 9 2
27 1 9 2 15 13 9 11 9 0 0 0 9 2 11 2 2 15 13 2 16 9 1 0 9 11 13 2
20 0 0 9 13 1 11 9 11 11 2 15 13 13 0 0 9 1 12 9 2
26 10 9 2 0 1 9 12 2 7 12 2 9 0 9 11 1 11 2 13 9 9 9 1 10 9 2
30 11 13 1 9 10 9 12 9 2 12 9 7 12 9 2 1 9 2 15 15 13 12 9 2 12 9 7 12 9 2
22 1 0 9 2 15 15 13 3 12 9 2 13 1 9 1 9 1 0 0 9 11 2
22 1 10 0 7 0 9 9 13 3 0 9 0 0 9 1 0 9 0 7 0 9 2
9 14 12 9 11 13 9 11 11 2
11 13 15 3 1 12 9 3 16 1 9 2
16 13 15 1 9 0 9 2 15 9 3 13 0 0 9 11 2
17 9 1 9 3 13 12 9 1 12 0 2 9 13 7 15 13 2
4 9 1 11 13
2 11 2
18 0 9 1 0 9 13 3 1 9 1 9 1 11 2 0 9 11 2
13 1 9 15 13 9 2 7 15 7 1 0 9 2
22 0 9 13 1 15 2 7 10 9 13 3 1 9 0 7 0 9 0 1 0 9 2
9 1 9 11 13 12 9 0 9 2
15 1 0 0 9 1 9 0 9 3 13 3 1 9 11 2
20 10 9 0 11 7 0 9 7 11 15 13 1 9 11 2 15 4 15 13 2
10 9 13 1 9 9 14 12 0 9 2
16 1 9 11 13 1 9 10 9 2 15 15 3 13 1 9 2
15 9 1 11 13 3 1 0 15 9 9 9 11 1 9 2
16 0 12 9 0 9 11 1 11 13 13 11 1 12 2 9 2
13 9 0 9 2 15 15 13 0 9 1 9 1 11
5 11 15 13 1 9
2 11 2
24 0 9 11 11 13 0 9 2 16 9 1 9 3 13 7 9 7 9 13 9 13 15 9 2
33 1 9 0 0 0 9 1 11 3 11 13 1 0 9 2 0 9 0 9 2 2 1 15 15 13 10 9 3 7 3 0 9 2
18 1 9 0 9 13 11 11 2 9 0 0 0 9 1 0 0 9 2
6 11 7 11 13 0 9
9 11 13 9 1 9 1 9 0 9
2 11 2
18 0 7 0 0 9 3 13 9 1 9 9 0 9 1 9 1 11 2
13 9 3 13 9 0 9 1 0 9 1 0 9 2
26 9 1 11 13 11 11 2 15 13 1 9 0 9 2 7 1 0 9 9 9 9 11 11 2 11 2
29 2 13 15 0 9 2 3 0 7 0 2 15 13 9 0 9 7 3 13 9 1 2 0 2 9 1 0 9 2
14 11 13 1 10 9 3 0 2 2 13 11 2 11 2
39 0 9 9 11 11 2 11 3 1 11 13 9 0 2 0 9 7 13 2 16 3 2 16 4 13 9 0 9 2 4 11 13 1 0 0 9 1 11 2
24 2 11 13 3 2 7 15 13 2 16 7 3 13 2 3 0 0 9 11 2 2 13 11 2
194 0 9 3 2 13 2 2 9 0 0 9 1 9 0 9 1 9 0 9 2 1 9 0 9 0 13 1 0 9 7 13 1 9 9 2 2 9 0 2 3 0 9 2 2 15 13 12 2 9 7 1 15 15 13 9 1 9 7 9 0 1 9 0 9 2 0 9 2 0 9 7 0 9 0 0 9 2 9 7 0 9 2 2 9 0 9 1 9 9 0 9 1 0 9 1 0 9 2 2 9 0 9 1 9 0 9 7 0 9 1 0 9 2 2 9 0 9 7 3 0 9 9 1 0 9 2 3 13 0 13 9 2 2 0 9 15 9 0 9 1 11 2 2 9 9 1 9 0 0 9 1 2 0 2 9 2 1 9 15 9 0 9 0 9 1 11 2 2 9 0 9 1 9 1 9 7 9 0 2 0 2 9 1 11 7 10 9 7 9 1 0 9 9 2
34 0 9 13 2 16 9 0 9 0 9 1 0 9 2 7 15 3 1 9 0 9 2 9 7 9 2 13 0 9 3 1 9 9 2
32 1 10 9 0 9 1 9 10 9 15 12 2 9 11 13 13 1 15 9 1 11 2 15 9 13 12 9 9 2 0 9 2
6 11 13 2 1 11 9
2 11 2
17 0 9 0 11 13 1 9 1 11 10 0 12 9 1 0 9 2
12 12 9 13 1 0 9 0 9 3 12 9 2
15 0 9 9 13 9 2 14 3 10 9 13 1 9 9 2
22 2 13 3 0 2 2 13 12 0 9 3 2 16 13 1 9 1 9 10 0 9 2
17 9 1 9 0 11 1 0 9 13 9 9 1 9 9 7 9 2
33 9 0 9 9 7 9 11 11 11 11 13 10 9 1 9 0 11 1 9 7 16 9 13 2 16 15 1 9 9 13 0 9 2
5 11 13 1 9 11
2 11 2
30 11 13 0 15 0 2 0 7 0 9 1 11 2 16 4 15 13 1 11 1 0 0 9 2 7 10 9 13 0 2
9 1 11 15 13 0 9 11 11 2
30 13 1 9 1 0 9 0 0 9 1 0 9 11 7 11 0 9 14 1 0 9 11 2 0 0 12 9 1 11 2
6 11 2 9 1 9 9
5 11 2 11 2 2
7 0 9 3 13 1 11 2
20 1 0 9 11 11 15 13 0 0 7 0 9 1 10 9 1 9 0 9 2
24 9 13 2 16 3 0 9 4 13 0 0 9 1 11 2 15 7 3 13 0 9 1 9 2
24 0 9 1 11 2 11 2 11 7 0 9 2 15 15 9 13 2 13 1 9 1 9 9 2
16 3 1 12 9 9 13 3 12 9 2 3 9 13 0 9 2
19 3 15 1 9 9 13 7 9 0 0 9 11 2 0 1 9 1 11 2
37 1 0 9 2 3 13 0 13 0 9 1 0 2 13 9 0 0 9 1 11 2 9 0 9 7 9 2 16 9 9 9 4 3 13 1 9 2
5 11 13 1 9 11
2 11 2
24 0 9 3 13 9 0 0 9 11 11 2 16 4 1 15 13 3 13 1 9 1 0 11 2
25 13 2 16 9 9 11 11 1 9 1 0 11 13 9 1 9 9 1 0 0 9 2 11 2 2
23 0 9 1 0 11 11 11 1 0 9 13 2 16 1 9 9 11 4 3 13 0 9 2
5 9 2 9 7 9
15 9 13 9 9 7 9 13 12 1 9 9 9 0 9 2
23 9 11 13 11 11 3 1 9 2 16 0 9 13 13 7 13 2 16 16 4 15 13 2
37 1 0 9 2 11 7 11 1 9 1 0 9 2 13 1 0 13 7 12 9 0 9 2 0 2 15 3 3 13 9 9 0 2 7 9 0 2
26 0 2 0 2 13 11 9 7 9 15 15 2 2 13 16 9 2 2 2 2 7 16 9 2 2 2
15 10 9 2 2 2 15 7 13 2 2 0 0 11 2 2
78 1 10 9 9 1 15 13 0 2 9 2 9 3 13 4 13 16 0 9 2 9 1 0 9 2 15 2 3 15 1 9 13 2 3 1 9 13 2 15 15 3 13 2 9 2 11 11 10 9 3 13 13 2 14 3 0 9 9 2 2 3 15 13 3 1 0 9 2 7 13 10 9 3 16 9 7 9 2
42 10 9 9 13 1 0 9 2 3 1 9 9 9 0 10 9 9 7 1 10 0 0 9 1 9 0 9 2 14 0 2 7 1 10 9 13 13 3 0 0 9 2
39 2 15 3 7 3 3 3 13 0 16 9 2 2 2 15 13 3 7 3 13 2 2 13 9 9 2 11 1 9 1 9 11 1 9 12 1 9 9 2
41 3 13 2 9 3 3 13 2 16 4 3 13 13 10 9 2 15 3 13 1 0 9 7 9 2 7 16 4 13 2 16 9 13 0 1 0 10 9 0 2 2
29 1 0 12 9 4 13 9 1 9 7 9 2 15 15 3 1 0 9 16 0 9 13 9 0 3 1 0 9 2
42 13 4 0 9 9 1 9 2 9 2 7 9 2 0 9 7 9 2 0 1 15 1 9 9 0 9 9 7 1 9 2 7 1 9 2 2 15 13 1 9 0 2
34 1 0 0 9 12 0 9 2 15 13 9 7 9 2 10 9 13 1 0 9 2 15 4 3 9 13 2 3 13 1 10 9 0 2
48 0 0 9 9 13 1 9 3 0 2 16 1 0 9 0 9 9 9 7 2 9 2 2 7 2 0 9 2 3 0 7 0 9 13 2 13 7 9 9 2 16 4 13 0 9 2 13 2
15 1 0 9 9 13 0 9 0 9 0 2 0 11 11 2
20 1 9 12 4 10 9 13 3 9 9 2 2 0 9 2 2 0 11 11 2
11 1 9 0 9 13 1 9 3 0 9 2
53 9 9 9 9 11 11 1 9 9 9 13 3 0 9 2 9 0 0 9 7 9 9 2 0 2 0 2 0 2 2 7 0 9 0 9 7 9 2 9 9 7 9 2 15 13 0 1 9 7 9 10 9 2
33 0 0 9 9 9 1 9 0 9 9 7 9 9 9 1 9 9 9 15 14 13 2 7 3 1 12 9 13 1 0 0 9 2
15 9 13 9 9 7 9 13 12 1 9 9 9 0 9 2
23 9 11 13 11 11 3 1 9 2 16 0 9 13 13 7 13 2 16 16 4 15 13 2
31 10 0 2 7 3 13 13 7 0 2 9 2 0 2 9 2 2 13 15 3 2 2 7 10 0 9 3 13 0 13 2
5 12 9 0 0 9
19 1 10 9 4 13 13 12 0 0 9 2 15 3 13 0 10 0 9 2
26 3 1 9 9 12 4 1 0 9 13 0 9 2 4 13 0 9 7 4 13 0 2 0 9 9 2
28 1 10 9 15 13 12 1 0 7 3 0 0 9 7 3 3 13 1 0 9 13 2 16 15 10 9 13 2
38 10 9 4 13 2 13 0 2 9 9 2 7 15 3 13 1 0 2 0 9 2 0 1 9 7 0 15 9 2 15 1 9 1 9 0 9 13 2
36 2 13 0 9 2 15 4 9 0 15 9 2 0 1 0 9 13 1 12 9 7 15 4 13 2 16 4 15 0 9 13 9 0 0 9 2
29 2 13 15 15 9 1 10 0 9 2 0 9 1 9 1 12 9 7 13 15 10 0 9 2 1 15 13 13 2
71 2 13 0 9 2 3 0 2 0 9 2 2 15 1 9 9 1 0 2 9 0 9 9 13 2 7 1 0 9 13 3 2 9 3 3 13 7 3 9 13 9 2 15 13 0 9 0 9 2 9 13 13 2 15 13 2 7 13 15 3 2 2 7 7 0 9 9 9 0 9 2
27 13 15 3 9 0 7 13 4 10 9 1 0 0 9 7 1 3 0 0 2 3 0 7 0 2 9 2
43 16 4 13 3 13 9 16 1 10 0 0 15 9 2 16 4 13 1 3 0 9 0 9 2 7 3 1 9 2 2 3 4 3 13 13 0 9 12 9 0 0 9 2
8 1 10 9 4 13 0 9 2
26 10 0 0 15 9 10 0 9 13 2 10 9 3 13 10 0 9 2 1 15 10 0 0 9 13 2
31 7 10 3 0 9 16 11 7 11 13 10 2 16 0 2 0 2 9 1 9 7 10 3 0 9 3 13 10 9 3 2
28 0 9 13 0 9 1 15 9 0 9 2 3 7 1 0 9 2 7 15 15 10 9 13 13 7 1 9 2
24 3 13 0 2 16 13 1 12 9 3 16 1 0 9 7 16 13 0 13 1 0 9 3 2
41 13 13 0 9 9 0 9 2 13 15 10 9 3 3 13 9 1 15 9 2 7 7 9 2 15 13 1 15 13 2 13 13 9 0 9 7 13 9 0 9 2
48 10 2 3 0 7 0 9 2 16 13 15 0 2 13 13 3 2 16 4 13 1 9 0 2 0 7 0 2 2 7 7 0 2 0 7 0 2 9 2 16 4 0 9 13 13 7 3 2
30 13 1 15 2 3 3 0 9 2 0 0 9 2 0 7 3 0 0 9 2 7 3 14 3 2 0 2 0 9 2
66 13 4 13 0 2 16 15 13 13 0 9 7 16 4 15 1 10 9 3 13 2 16 4 2 13 3 0 0 9 2 0 2 0 2 9 2 13 2 16 13 1 10 0 9 0 9 2 13 0 9 0 9 2 13 0 0 2 7 7 0 2 9 10 0 9 2
42 13 2 16 7 9 2 7 9 2 7 10 0 9 4 3 10 9 13 1 9 1 0 9 7 4 13 1 15 2 16 2 3 1 10 9 2 13 15 1 0 9 2
6 9 0 2 7 0 2
10 10 9 13 3 0 9 9 1 9 2
18 1 12 9 1 0 9 2 15 13 2 4 12 13 16 0 9 9 2
22 1 0 9 2 13 15 1 9 1 9 2 0 9 2 2 13 13 9 9 1 0 2
25 9 13 3 13 16 9 9 2 7 7 16 9 1 0 9 2 15 3 12 1 9 9 9 13 2
9 9 1 9 0 9 13 3 0 2
11 0 2 0 9 1 9 13 13 0 9 2
18 9 9 1 9 2 13 0 9 9 9 1 12 9 2 7 13 0 2
37 1 0 9 9 11 11 13 9 9 12 2 9 9 2 0 1 15 2 16 9 13 13 15 2 15 4 0 7 0 9 13 0 7 0 9 9 2
9 9 0 7 0 13 14 3 0 2
13 9 1 9 1 9 13 3 0 7 3 3 0 2
15 10 9 15 13 9 0 9 2 1 9 0 13 3 9 2
22 9 1 9 7 3 13 7 9 9 13 0 7 0 2 15 13 1 3 0 0 9 2
13 9 11 1 9 9 7 9 1 11 13 3 0 2
48 0 13 3 9 2 16 0 9 13 1 0 9 2 15 13 1 9 9 0 9 3 0 7 0 2 7 16 1 15 13 3 14 10 9 1 0 9 2 9 9 3 10 0 9 3 13 2 2
12 1 10 9 13 1 9 15 9 9 1 9 2
23 0 9 15 13 15 9 0 9 2 16 0 9 9 2 1 15 4 15 13 0 9 13 2
8 0 9 7 13 13 7 3 2
35 13 3 13 2 16 9 9 13 9 13 2 16 13 15 0 13 9 0 0 9 2 7 15 3 3 13 0 9 9 1 9 1 10 9 2
35 0 0 9 13 9 2 16 7 9 13 1 9 9 2 7 13 15 7 13 9 9 0 9 1 9 2 15 4 3 13 13 7 10 9 2
18 3 15 9 1 9 13 7 3 4 10 9 9 13 2 13 3 9 2
9 3 15 13 3 9 1 0 9 2
25 16 13 13 7 0 9 9 2 13 4 10 9 13 3 2 1 15 9 9 7 1 10 0 9 2
1 9
16 1 0 9 9 0 9 13 0 9 0 11 11 2 1 11 2
29 0 13 3 1 9 12 13 10 0 9 1 10 12 0 9 2 7 7 10 9 1 0 9 13 3 12 12 9 2
29 1 12 9 2 15 15 13 1 9 11 7 3 13 1 9 11 11 2 13 1 9 1 9 1 11 9 0 9 2
14 11 13 9 13 0 9 9 1 9 9 2 3 13 2
7 3 3 13 9 12 9 2
6 9 13 1 9 7 9
2 11 2
25 9 1 12 9 13 1 3 0 9 2 15 15 1 9 0 9 13 1 0 9 1 11 1 11 2
9 13 1 15 9 2 9 7 9 2
21 1 0 9 1 0 9 15 13 9 1 9 13 1 9 0 1 9 2 15 13 2
13 3 15 2 3 1 9 2 13 1 0 9 9 2
5 9 13 1 9 9
5 11 2 11 2 2
14 1 0 9 9 4 13 12 0 11 11 2 1 11 2
27 1 0 9 13 2 16 0 1 9 1 9 12 13 1 9 9 1 11 9 1 12 9 2 15 7 13 2
34 1 9 7 1 9 12 13 3 1 9 0 11 2 12 9 2 7 1 9 7 9 1 9 9 11 2 3 15 13 9 1 12 9 2
15 9 9 3 13 7 15 9 13 1 10 0 9 1 11 2
4 0 9 13 9
5 11 2 11 2 2
16 9 12 0 9 13 0 9 9 1 11 7 0 11 1 11 2
29 16 15 12 0 9 11 2 11 2 1 11 11 13 1 9 9 2 13 1 0 9 2 13 15 1 9 7 13 2
5 9 13 1 9 2
6 9 9 13 1 9 2
8 9 13 2 9 13 0 9 2
6 9 9 13 0 9 2
11 9 0 9 1 9 9 13 14 9 1 9
2 11 2
28 9 0 9 1 9 9 13 9 1 9 2 7 9 0 9 9 9 7 9 9 16 0 9 1 9 0 9 2
11 1 0 9 9 15 13 9 9 11 11 2
28 9 0 9 9 1 9 12 9 1 0 9 1 9 13 1 11 9 2 16 1 9 13 9 1 9 7 9 2
24 13 3 1 0 9 9 2 13 9 7 13 2 16 0 9 9 13 1 9 9 1 0 9 2
31 9 0 0 9 11 11 13 2 16 9 1 9 4 3 13 7 9 9 2 13 2 2 16 4 13 1 9 9 7 9 2
13 0 9 9 1 9 13 1 10 9 3 0 9 2
33 2 13 2 14 0 9 13 7 13 2 14 15 13 0 7 0 9 9 1 9 2 13 0 9 13 7 9 2 7 9 7 9 2
16 13 15 3 1 12 9 10 9 13 3 0 2 2 13 11 2
18 9 9 1 9 1 10 9 13 15 2 16 1 15 4 13 15 9 2
21 1 9 2 1 15 13 9 13 2 13 15 3 0 9 9 1 9 2 13 11 2
39 9 11 11 1 0 9 13 2 16 15 3 0 9 1 9 9 13 7 1 15 3 9 13 2 15 3 13 0 13 10 9 1 9 10 9 1 12 9 2
25 1 10 0 9 1 9 1 9 1 9 11 15 14 11 13 3 13 2 3 10 9 13 9 9 2
6 11 13 11 1 9 11
5 11 2 11 2 2
16 9 0 9 16 0 2 3 0 0 9 13 0 9 1 9 2
15 1 9 12 2 9 9 15 13 10 3 0 9 11 11 2
11 11 13 3 12 9 7 12 9 1 9 2
21 1 0 0 9 13 11 0 9 2 15 14 13 13 14 0 9 2 7 0 9 2
11 1 9 13 11 13 3 1 9 0 9 2
10 1 9 13 7 9 1 9 10 9 2
15 11 3 13 2 16 9 13 9 9 7 13 1 0 9 2
25 0 9 9 11 11 15 10 9 1 0 9 13 1 15 2 16 15 1 9 13 13 7 0 9 2
6 11 3 13 1 0 9
6 11 11 2 11 2 2
38 3 1 9 2 16 4 0 9 13 1 9 1 9 9 7 11 1 0 9 1 9 10 0 9 2 13 0 9 13 1 0 9 0 0 9 1 9 2
9 13 1 0 9 4 7 13 0 2
27 11 15 1 9 13 9 11 11 1 9 2 15 4 15 13 13 1 9 9 11 2 15 13 12 9 9 2
36 0 9 9 11 11 1 15 13 2 16 11 15 1 9 13 13 2 13 0 0 9 2 15 1 15 1 9 12 13 0 9 1 10 9 3 2
5 11 13 1 9 9
5 11 2 11 2 2
14 2 1 0 9 13 0 2 16 9 13 1 9 0 2
37 3 1 12 9 1 15 13 9 7 0 9 13 9 1 9 7 1 0 9 2 2 13 1 9 1 0 9 11 2 11 1 11 10 9 11 11 2
44 1 9 1 9 0 9 2 15 13 1 9 9 11 11 11 9 9 2 11 1 0 11 3 13 2 16 15 13 9 2 1 15 9 13 9 2 16 1 9 13 15 1 9 2
11 9 11 13 1 10 0 9 1 9 1 11
4 11 2 11 2
32 9 11 1 0 9 7 0 2 0 9 13 0 9 0 0 9 0 9 11 1 9 3 0 0 0 9 2 11 2 1 11 2
34 1 9 11 11 11 13 10 9 0 1 0 9 9 1 0 0 9 0 9 7 13 9 0 9 9 1 0 9 1 9 0 0 9 2
17 1 0 9 13 11 9 1 0 7 0 9 7 3 9 0 11 2
27 9 0 9 11 11 11 1 11 13 2 16 11 13 0 9 1 15 2 16 4 0 9 13 3 1 11 2
10 13 9 10 9 15 1 0 9 13 2
17 2 9 1 11 4 13 15 2 11 13 3 1 11 2 2 13 2
25 9 9 11 11 11 13 2 16 1 0 9 13 3 2 1 9 1 9 0 0 9 1 9 11 2
10 9 11 11 7 10 9 13 1 9 9
5 11 2 11 2 2
27 9 0 9 3 0 11 11 13 0 9 1 9 9 2 10 9 11 11 3 7 1 9 1 9 1 9 2
28 12 13 1 0 9 9 1 9 11 11 2 15 15 1 9 1 11 2 11 12 2 9 13 1 9 11 12 2
18 9 9 11 11 11 13 9 9 1 9 7 1 9 1 9 9 13 2
18 11 12 13 0 11 11 2 2 15 13 0 9 12 9 0 0 9 2
11 12 11 15 3 10 9 13 1 0 9 2
11 11 4 13 0 9 2 15 13 9 9 2
7 1 11 11 9 13 4 2
11 9 13 9 2 1 15 9 13 11 11 2
26 1 9 11 11 2 13 10 9 0 2 7 15 0 9 13 10 0 9 1 9 1 11 1 9 9 2
11 9 2 15 13 13 2 13 1 9 0 2
13 11 13 1 10 9 1 9 9 0 2 9 2 11
7 11 2 11 2 11 2 2
24 9 13 16 9 9 7 9 0 9 9 13 15 1 0 9 2 7 15 7 1 9 1 15 2
27 1 9 1 9 11 11 2 11 2 1 9 9 0 9 11 11 11 15 13 9 9 11 11 2 11 2 2
28 11 9 13 2 16 1 10 9 13 9 9 11 11 2 11 2 2 10 9 13 4 9 1 9 0 9 13 2
21 1 9 13 3 3 9 9 11 2 3 7 13 1 10 9 7 0 9 0 9 2
19 16 15 13 11 2 9 3 13 9 13 1 0 9 1 3 0 9 11 2
17 2 0 9 13 1 9 2 7 1 9 9 9 2 2 13 9 2
11 0 9 14 13 1 9 0 2 0 9 2
21 1 9 2 16 0 2 9 2 11 13 9 11 2 11 13 2 16 1 15 13 2
11 9 1 15 13 9 9 1 9 0 9 2
20 3 9 9 11 4 1 9 9 12 13 1 9 9 7 9 2 13 9 9 2
4 1 9 1 9
12 13 0 0 9 1 0 9 1 0 9 0 2
8 13 15 3 1 10 9 13 2
24 11 11 2 11 2 2 9 9 2 3 15 13 13 2 1 15 15 13 7 9 1 0 9 2
21 15 3 13 3 7 16 13 0 2 0 9 9 2 13 2 16 13 9 1 9 2
38 3 13 0 13 2 3 15 13 1 3 0 9 2 7 15 3 4 13 7 0 9 2 1 15 15 13 14 1 0 12 9 1 9 2 7 1 12 2
6 15 13 3 3 9 2
24 11 11 2 11 2 2 9 2 15 4 13 2 16 13 12 9 10 7 15 7 16 15 13 2
28 9 13 1 10 9 15 13 2 16 1 9 0 9 7 9 13 9 9 1 0 0 9 2 0 1 0 9 2
23 3 2 15 15 13 13 7 13 13 2 16 9 13 9 0 9 7 16 15 13 0 9 2
19 3 7 4 13 9 9 2 15 3 13 2 16 13 1 0 9 7 13 2
7 3 15 1 15 3 13 2
8 3 3 15 13 3 3 9 2
26 11 11 2 0 9 2 13 15 3 9 2 7 3 3 13 13 2 3 1 9 10 9 1 9 13 2
15 14 16 13 1 9 15 2 3 15 15 13 2 7 3 2
2 13 2
15 3 16 4 15 13 14 0 12 9 2 15 4 3 13 2
26 11 11 2 0 9 2 16 4 9 13 1 15 2 3 4 15 13 10 9 7 13 4 0 15 13 2
16 11 11 2 0 9 2 13 2 16 13 10 9 9 7 15 2
13 7 13 2 16 4 15 1 15 13 10 9 9 2
15 15 1 15 13 2 16 4 15 12 9 1 9 13 13 2
5 13 9 1 9 11
5 11 2 11 2 2
45 1 9 2 16 4 9 13 0 9 3 1 0 0 9 11 2 11 11 7 9 1 9 2 3 0 0 9 11 2 2 15 1 9 11 11 1 9 13 9 11 11 2 11 2 2
16 13 14 13 2 16 9 9 13 9 2 0 9 7 0 9 2
21 3 13 2 3 11 2 11 11 13 1 9 12 1 0 9 1 9 7 12 9 2
46 9 4 1 11 13 13 2 15 15 0 9 2 16 4 9 9 7 9 0 9 2 9 7 9 2 0 1 0 9 2 13 13 9 0 9 7 13 15 1 9 9 1 0 9 2 2
7 11 13 9 2 0 9 2
5 11 2 11 2 2
19 9 11 11 11 13 1 2 3 0 2 9 11 1 9 9 1 0 9 2
18 9 4 1 11 13 13 2 16 4 15 0 0 9 13 3 13 9 2
21 2 13 0 9 2 16 13 3 1 15 9 3 9 16 10 9 2 2 13 11 2
14 9 0 4 14 3 1 11 3 0 9 13 3 3 2
19 13 3 1 9 9 2 7 1 0 9 0 9 1 9 7 9 9 9 2
20 1 0 13 11 1 10 9 7 0 9 9 1 11 2 14 12 9 9 2 2
15 13 15 14 9 15 2 3 0 9 13 0 13 10 9 2
1 3
20 2 9 13 0 2 13 9 0 9 1 9 9 7 0 9 0 9 0 9 2
21 9 13 9 9 2 15 13 1 0 0 9 11 13 2 0 3 2 0 9 2 2
21 9 11 0 2 9 2 2 0 11 11 13 2 16 4 9 1 12 2 9 13 2
14 1 9 2 16 4 13 2 13 9 9 1 0 9 2
11 9 0 9 1 9 13 1 9 1 11 2
13 10 0 0 9 13 0 9 1 9 1 0 9 2
28 1 9 9 15 9 7 9 0 9 13 13 0 7 0 9 1 9 0 9 1 9 7 11 1 9 0 9 2
9 9 13 3 2 0 9 1 11 2
16 9 1 0 9 9 13 3 3 1 9 9 9 9 2 9 2
17 0 9 13 9 13 1 9 9 2 1 9 0 12 2 11 12 2
14 0 9 4 13 1 9 11 7 1 9 0 9 9 2
23 9 0 0 9 2 9 1 9 9 7 9 2 15 13 1 9 1 0 1 11 11 11 2
18 3 16 12 9 0 9 0 7 3 0 9 13 13 1 9 12 9 2
10 9 13 0 9 9 0 0 9 11 2
6 9 13 14 3 14 3
5 11 2 11 2 2
14 3 1 12 9 1 0 9 4 3 1 9 13 9 2
13 11 15 13 9 11 11 1 0 0 9 1 11 2
12 1 15 13 15 1 9 1 0 9 3 3 2
7 0 9 3 7 4 13 2
15 9 13 3 0 9 1 0 9 9 7 9 1 10 9 2
28 1 15 4 13 9 9 9 9 7 9 1 9 2 7 15 1 11 2 0 11 2 11 2 11 7 0 9 2
11 3 15 0 9 13 3 1 0 0 9 2
10 0 0 9 13 3 0 1 0 11 2
17 13 15 7 1 0 2 15 13 3 1 11 7 11 3 0 9 2
31 1 11 11 13 3 9 3 0 9 1 9 1 11 2 3 1 11 2 3 15 9 13 1 0 9 1 11 7 1 11 2
14 1 9 3 13 9 1 15 0 9 2 3 7 3 2
25 9 9 9 13 1 11 7 0 11 2 1 0 7 0 11 7 1 11 15 13 3 7 9 9 2
5 11 13 9 1 9
5 11 2 11 2 2
18 2 15 13 9 2 15 13 0 9 2 0 1 9 0 7 0 9 2
10 9 13 9 9 11 11 2 11 2 2
22 2 3 1 9 4 3 13 1 0 9 7 13 9 2 3 13 9 7 0 0 9 2
12 13 4 13 2 16 0 9 10 9 3 13 2
20 3 13 0 2 16 10 9 13 14 0 7 0 2 2 13 0 11 2 11 2
14 3 13 0 2 0 9 2 1 0 9 13 1 9 2
18 16 13 2 1 9 13 10 0 9 1 9 13 0 9 9 11 11 2
23 2 13 4 15 2 13 4 1 15 1 9 7 13 4 15 13 16 0 3 7 3 2 2
5 9 13 9 9 2
21 1 0 9 13 3 3 0 0 9 9 9 2 7 4 7 13 1 9 0 9 2
31 1 9 1 9 13 1 9 9 3 3 0 9 9 1 0 9 2 3 0 9 0 1 0 9 9 7 3 1 9 13 2
7 0 9 13 1 11 12 12
2 11 2
24 1 10 0 9 13 1 0 9 12 0 0 9 2 1 15 15 13 3 12 7 9 9 9 2
7 3 0 13 0 0 9 2
17 3 12 9 13 12 0 9 7 12 9 13 9 12 0 0 9 2
11 12 9 0 9 7 9 13 12 0 9 2
18 0 9 15 13 7 1 9 0 9 7 12 0 0 9 13 12 9 2
8 1 11 4 9 0 9 13 2
20 10 0 3 0 0 9 4 1 0 9 13 1 0 9 7 13 3 0 9 2
10 3 7 9 9 1 9 0 9 13 2
16 9 13 0 1 0 9 2 3 15 3 13 1 12 9 3 2
8 9 9 13 9 0 9 10 9
5 11 2 11 2 2
17 9 0 9 10 9 1 9 12 13 9 9 0 9 0 12 9 2
7 13 15 1 9 9 11 2
22 0 0 0 2 12 5 2 13 2 16 0 9 10 9 13 3 0 16 1 9 12 2
18 9 13 0 0 2 12 5 2 7 9 0 0 2 12 5 2 9 2
20 1 9 3 13 2 16 1 0 9 7 0 9 9 13 9 9 9 0 9 2
23 3 9 3 13 0 9 1 12 9 2 12 5 2 7 9 1 0 9 2 12 5 2 2
12 9 13 9 11 1 9 0 9 1 12 9 2
4 9 9 13 13
3 0 11 2
18 0 9 9 9 7 0 9 11 11 1 0 9 13 9 9 1 9 2
18 1 0 9 9 9 9 0 2 11 15 1 9 13 9 11 11 11 2
22 9 0 9 11 11 10 9 13 7 13 2 16 2 1 0 9 9 13 0 9 2 2
22 9 12 13 11 1 9 0 15 9 1 3 0 1 9 9 9 1 9 7 1 9 2
21 1 9 9 13 1 10 9 3 9 0 7 0 9 1 12 9 7 9 0 9 2
18 9 9 9 13 13 0 9 1 9 3 2 15 7 1 9 13 13 2
20 11 13 1 0 2 16 4 13 9 12 7 12 9 1 9 7 12 9 9 2
20 9 9 13 1 11 12 9 2 1 15 3 9 7 13 0 9 1 0 9 2
19 0 9 11 11 2 3 2 2 9 11 11 7 0 9 11 11 2 3 2
7 9 15 13 1 9 1 9
2 11 2
17 9 0 9 1 11 1 11 15 13 1 9 11 11 1 0 11 2
16 1 12 0 13 7 9 2 11 11 1 11 2 15 13 0 2
11 9 15 13 1 12 9 1 9 12 9 2
15 1 0 12 13 9 1 9 12 9 7 13 3 12 9 2
9 0 9 15 15 1 9 9 13 2
12 3 2 1 9 9 2 15 13 9 1 9 2
10 13 15 2 15 1 0 9 13 3 2
8 9 1 9 9 13 9 0 9
2 11 2
17 9 0 9 11 11 2 11 2 13 1 0 9 1 0 9 9 2
26 13 2 16 9 13 9 1 9 9 9 0 9 2 0 9 0 2 9 2 2 16 13 0 0 9 2
18 3 13 2 16 0 9 13 9 13 15 1 9 13 1 9 3 9 2
22 1 9 9 9 9 1 9 12 0 9 0 9 0 2 9 13 0 9 3 9 9 2
11 1 10 9 3 13 9 1 0 0 9 2
16 9 4 7 1 9 1 0 9 3 13 12 9 1 0 9 2
13 1 9 1 9 0 9 0 9 15 13 0 9 2
9 9 15 9 13 1 12 9 9 2
13 9 9 13 9 2 15 9 13 1 9 0 9 2
15 13 3 1 0 9 2 1 15 4 1 11 13 0 9 2
13 0 9 1 9 9 0 2 9 4 13 1 9 2
11 1 0 9 4 13 9 13 1 9 9 2
26 11 2 11 1 9 13 3 9 9 1 0 0 9 12 11 2 15 13 13 1 0 9 1 0 9 2
3 9 1 9
35 9 2 3 13 10 9 2 13 3 1 0 9 2 16 13 9 0 2 15 14 13 2 7 3 15 13 2 7 9 0 2 0 0 9 2
5 15 13 1 9 2
29 12 1 0 9 9 13 2 16 10 9 1 0 7 0 9 2 16 3 4 15 13 15 2 13 1 9 9 13 2
23 0 9 1 9 13 3 0 7 3 15 2 0 2 0 2 0 2 0 2 0 2 0 2
17 9 13 2 13 2 13 9 2 13 2 9 13 2 13 7 13 2
17 9 9 13 9 1 9 7 0 9 13 10 0 9 1 0 9 2
32 14 3 10 9 13 10 9 3 13 7 14 3 3 3 13 10 9 1 9 13 2 16 9 3 13 3 9 13 16 9 0 2
15 3 0 0 9 11 7 13 10 0 2 13 9 1 15 2
15 13 2 16 9 13 0 2 13 2 16 13 2 16 13 2
3 16 13 2
19 9 13 10 9 7 15 13 15 10 9 13 1 15 2 16 4 15 13 2
16 3 3 13 0 9 2 13 11 11 3 1 9 1 9 11 2
24 1 0 9 13 1 9 0 9 3 0 9 2 16 12 0 4 13 1 0 9 7 0 9 2
20 1 9 2 3 15 1 0 9 13 2 13 15 14 2 3 2 3 2 3 2
15 13 15 2 16 10 9 15 15 13 7 13 1 0 0 2
19 11 11 13 2 15 1 0 9 7 9 13 9 7 15 13 1 9 9 2
18 16 0 9 13 15 0 2 16 13 9 9 2 15 15 13 9 9 2
28 3 13 1 9 9 9 0 9 2 9 0 9 2 9 7 9 2 0 9 2 15 15 13 9 0 0 9 2
23 7 3 1 10 0 9 13 9 2 9 2 15 1 0 9 13 2 16 9 15 3 13 2
11 15 11 11 13 13 15 9 9 7 9 2
20 0 4 11 3 13 7 13 2 16 9 10 3 0 9 13 3 9 10 9 2
30 13 0 13 15 2 16 10 7 15 9 13 9 2 16 13 9 7 9 2 16 4 9 13 1 9 7 13 10 9 2
16 9 15 15 13 2 15 13 13 7 10 9 13 10 9 0 2
35 10 9 13 1 0 9 2 10 9 15 13 1 9 2 10 9 13 2 15 15 13 2 7 15 2 15 10 0 0 9 13 2 15 13 2
9 7 15 15 13 2 15 4 13 2
12 15 13 9 1 9 7 11 11 15 3 13 2
25 0 11 2 0 0 9 2 13 1 11 0 9 11 11 2 0 9 11 11 7 0 9 11 11 2
10 0 9 13 9 11 11 2 3 2 2
4 0 11 9 9
2 11 2
32 11 2 0 9 0 11 2 13 1 9 16 0 9 9 0 9 9 11 11 2 15 13 9 9 0 9 1 9 11 1 9 2
22 0 0 9 4 13 11 11 1 9 1 9 9 11 7 11 11 2 9 0 9 2 2
8 1 11 13 15 3 0 11 2
23 0 9 11 15 13 9 9 11 9 11 11 2 0 0 9 9 1 11 1 12 2 9 2
21 11 11 1 0 0 9 1 9 13 11 1 11 9 11 2 11 11 1 11 11 2
21 0 0 9 13 1 10 9 1 12 9 2 15 13 11 1 0 9 1 0 9 2
16 0 0 9 15 13 0 9 12 9 7 12 9 9 11 11 2
9 9 13 11 2 15 13 12 9 9
2 11 2
13 12 9 9 13 9 1 9 1 0 9 1 11 2
12 13 1 15 9 0 9 0 9 9 11 11 2
20 9 2 15 13 1 0 9 9 14 12 9 9 2 4 13 1 9 0 9 2
14 15 1 0 9 13 9 0 9 11 2 11 2 11 2
11 9 13 1 11 0 1 0 9 0 9 2
11 1 9 1 9 13 9 0 9 9 11 2
24 0 0 11 4 9 1 11 12 13 1 9 0 9 0 9 7 9 0 7 0 9 7 9 2
13 0 4 13 1 0 9 1 9 1 9 1 9 2
13 16 4 13 0 2 13 15 12 7 12 9 9 2
12 3 4 1 9 0 9 13 3 12 9 9 2
13 13 15 0 9 10 9 0 9 1 0 12 9 2
13 1 9 12 7 12 15 13 3 1 12 9 9 2
14 1 12 9 2 0 9 2 13 0 9 1 9 12 2
8 0 9 0 3 13 9 1 11
2 11 2
30 0 9 11 11 13 0 9 10 12 0 9 1 11 1 9 0 9 11 2 16 15 9 9 4 13 13 1 0 9 2
12 13 15 1 9 1 11 9 0 9 11 11 2
48 13 3 2 16 1 10 9 3 4 3 13 2 7 0 9 15 3 1 0 9 13 13 0 9 11 11 2 16 4 13 10 9 1 9 3 12 9 9 3 2 16 10 9 12 2 9 13 2
6 3 1 11 1 9 12
5 0 9 13 1 11
2 11 2
16 1 0 0 0 9 13 3 1 0 9 0 9 11 11 11 2
16 3 15 13 13 1 9 11 11 2 1 10 9 15 9 13 2
15 13 15 3 1 9 0 9 11 11 7 1 9 11 11 2
27 9 10 9 1 11 13 7 9 11 2 3 15 13 9 11 7 13 15 1 9 0 9 7 0 9 11 2
7 3 13 11 0 0 9 2
6 9 1 11 13 12 11
4 11 2 11 2
23 3 12 0 9 13 1 9 2 16 1 9 1 0 9 0 9 11 13 3 3 0 9 2
12 13 15 9 0 9 1 11 0 1 0 11 2
15 0 9 11 3 13 1 2 0 0 0 9 2 1 11 2
16 9 9 13 2 16 1 12 9 13 14 9 9 2 3 9 2
20 2 15 3 13 1 9 9 2 7 0 13 2 16 4 13 0 2 2 13 2
6 11 7 11 13 1 9
2 11 2
18 11 7 0 9 13 9 0 15 9 0 9 7 9 9 0 0 9 2
4 9 1 9 12
8 9 11 13 0 1 10 11 9
2 11 2
23 0 9 11 11 13 0 1 10 9 1 0 9 1 0 0 9 2 0 9 11 11 11 2
21 9 3 1 9 1 0 9 1 0 11 13 2 16 10 9 15 13 3 0 9 2
31 9 0 9 0 1 11 13 1 11 0 7 4 3 3 13 1 9 2 7 7 13 0 2 16 4 0 9 13 0 9 2
13 11 7 13 13 9 11 1 10 9 1 9 9 2
26 11 11 1 9 13 2 16 15 13 9 13 0 9 2 16 15 1 9 11 11 13 1 9 0 9 2
9 11 7 11 4 15 13 13 3 2
12 1 9 0 9 11 11 4 11 13 1 9 2
24 9 9 15 13 9 0 2 0 9 1 9 2 3 4 13 0 9 9 7 3 13 10 9 2
4 0 9 0 9
2 11 2
17 0 0 9 15 1 0 9 13 1 12 9 1 9 1 9 12 2
8 1 9 4 13 3 0 9 2
13 13 15 1 9 2 15 1 9 13 0 0 9 2
25 0 9 13 1 0 9 12 9 9 2 12 9 9 2 2 15 13 1 0 9 1 12 9 3 2
20 0 9 13 1 0 9 1 12 9 2 16 1 9 12 13 9 9 12 9 2
9 9 0 9 15 13 1 12 9 2
22 9 0 9 13 3 1 12 9 2 15 13 2 16 1 11 3 13 14 12 9 9 2
11 9 9 15 1 9 12 13 1 12 5 2
10 0 0 0 9 3 13 1 12 5 2
18 0 0 9 15 13 3 1 12 5 2 3 7 13 3 1 12 5 2
32 1 0 9 13 1 9 9 2 1 10 9 13 0 0 9 9 12 9 9 2 15 13 1 12 9 9 3 16 1 0 9 2
25 9 1 0 9 13 1 9 7 9 1 0 9 2 15 1 9 9 7 9 12 13 12 9 9 2
5 0 9 7 1 9
2 11 2
31 9 1 9 0 0 9 13 9 2 16 4 0 7 0 9 1 0 9 2 1 15 15 10 9 13 2 13 7 1 9 2
11 9 10 9 13 9 13 9 1 0 9 2
36 16 13 0 9 0 11 2 1 0 9 9 15 13 3 0 9 2 16 15 3 1 9 3 3 13 9 13 0 9 0 2 3 0 2 9 2
11 0 9 9 15 13 13 14 1 9 12 2
29 0 0 9 2 15 13 3 3 0 0 0 9 1 0 9 2 1 9 13 0 9 0 9 1 11 7 1 11 2
13 9 1 0 9 4 15 13 13 1 12 1 12 2
23 3 15 3 13 1 0 9 9 0 9 2 16 1 15 4 13 9 9 1 15 0 9 2
41 9 1 0 9 2 13 1 0 11 11 11 2 0 9 0 9 2 15 13 13 0 9 1 9 0 9 7 13 15 9 0 9 2 1 15 3 0 9 3 13 2
15 3 13 9 9 13 10 9 2 16 4 13 1 9 13 2
13 9 13 1 0 12 9 7 4 13 0 0 9 2
26 9 0 9 13 0 9 1 9 2 9 2 0 9 2 0 9 7 9 2 9 2 9 7 10 9 2
37 9 7 13 0 9 2 0 15 2 16 15 1 9 12 13 1 0 9 1 9 3 2 1 10 9 15 7 9 1 9 13 9 1 0 0 9 2
4 0 9 9 9
11 9 0 9 1 0 7 0 11 4 3 13
21 0 9 0 11 13 12 2 9 0 9 0 3 0 0 9 2 0 2 0 9 2
11 0 11 13 1 15 7 13 3 12 9 2
20 1 9 13 0 3 12 9 2 9 2 3 3 13 0 0 9 0 0 9 2
23 9 10 9 13 1 9 10 9 3 3 13 2 16 0 9 3 10 9 13 1 0 9 2
30 1 9 15 4 13 13 1 15 2 16 9 3 0 13 13 1 10 0 9 2 7 15 7 1 10 9 2 3 3 2
27 0 9 13 1 0 9 3 0 2 3 3 1 15 2 15 15 13 13 0 9 0 9 1 9 0 9 2
22 1 9 13 2 16 1 0 0 9 13 3 0 9 1 9 1 9 0 7 0 11 2
18 13 1 9 2 13 15 2 16 9 13 2 2 15 13 15 1 15 2
26 1 10 9 13 0 2 11 13 13 3 2 11 3 2 11 2 0 11 7 11 3 7 0 9 3 2
33 1 0 9 13 1 9 7 3 7 1 0 9 0 0 9 2 2 3 0 0 9 0 11 11 13 0 9 1 0 0 9 2 2
26 1 0 9 9 2 1 15 13 0 9 1 0 9 2 13 13 9 0 9 1 10 0 7 0 9 2
29 14 2 1 0 9 12 9 2 3 0 9 2 15 13 12 0 2 12 0 7 0 12 4 15 13 13 1 0 2
22 1 9 13 9 10 9 2 0 9 13 9 2 0 9 13 1 9 7 0 0 9 2
18 0 0 9 13 2 16 13 13 9 9 1 0 11 1 0 0 9 2
39 7 4 0 9 13 0 9 3 3 3 16 9 2 7 1 15 0 9 0 9 11 1 11 13 3 3 0 16 9 0 0 0 9 1 9 1 0 9 2
6 0 9 13 3 0 2
17 16 15 13 2 9 1 10 0 9 13 3 0 7 1 9 9 2
7 0 14 9 2 7 7 9
19 3 13 1 0 9 9 11 9 0 1 9 9 11 12 1 9 14 9 2
18 1 0 9 10 9 9 4 13 9 13 0 9 1 10 3 0 9 2
29 3 0 9 11 12 13 0 9 0 0 9 2 7 9 1 0 9 0 9 2 9 3 13 0 9 15 12 9 2
20 9 9 11 9 0 11 11 1 9 13 2 2 9 13 13 15 0 2 0 2
16 13 4 9 1 9 7 9 2 1 15 13 13 9 3 9 2
22 3 4 13 1 0 9 2 13 15 7 7 9 0 9 2 15 7 13 0 9 2 2
12 0 9 13 0 9 1 0 9 1 0 9 2
22 9 15 3 3 13 1 9 1 9 2 7 7 7 1 11 12 13 9 0 0 9 2
8 14 16 4 15 13 1 9 2
15 3 2 1 0 9 9 7 0 9 13 9 9 3 0 2
10 9 15 7 13 13 9 7 9 9 2
16 3 0 9 1 0 9 13 2 16 15 15 10 9 13 13 2
20 1 9 4 13 0 9 0 1 11 11 9 0 9 12 9 2 12 9 2 2
21 11 12 0 0 9 13 1 10 9 3 0 9 1 12 1 12 9 1 12 9 2
21 7 1 9 0 1 9 12 9 13 0 0 9 1 0 9 7 0 0 3 0 2
11 0 9 4 13 9 2 15 13 3 0 2
16 1 0 9 13 13 12 9 1 9 2 9 13 0 0 9 2
20 1 0 9 15 13 13 0 9 0 3 0 9 2 15 9 13 3 12 9 2
16 1 10 0 9 4 13 13 0 9 1 9 7 0 9 9 2
10 11 12 13 3 0 9 0 0 9 2
25 15 15 7 13 13 1 9 1 9 13 12 9 2 3 15 1 9 9 1 0 0 9 13 4 2
15 12 1 9 1 0 15 9 1 11 13 7 9 11 11 2
15 0 0 9 13 9 12 2 9 2 15 13 3 10 9 2
13 9 13 0 9 1 9 12 9 1 9 12 9 2
17 0 9 13 12 9 2 9 1 9 1 12 1 12 1 12 9 2
4 9 16 0 9
11 9 1 0 13 1 15 0 2 7 3 0
8 0 9 1 0 9 13 9 2
15 3 15 13 1 9 1 11 13 12 2 1 15 9 13 2
18 9 1 15 0 2 16 10 9 13 4 13 9 7 0 9 13 13 2
7 13 2 16 4 4 13 2
20 9 1 9 12 9 2 9 13 9 1 0 9 7 1 0 9 1 0 9 2
24 13 0 9 1 9 2 3 0 1 9 2 15 13 0 2 16 13 15 13 1 9 1 9 2
24 1 9 9 9 0 7 0 1 0 9 1 0 9 4 16 0 9 13 1 0 9 1 9 2
22 1 0 0 9 13 1 9 0 9 13 2 16 0 9 13 13 13 10 0 0 9 2
7 15 15 13 1 9 9 2
23 1 9 1 12 9 13 1 1 3 0 9 9 7 0 9 9 0 9 9 1 9 9 2
9 1 0 9 13 3 0 0 9 2
13 0 0 9 3 9 1 12 2 12 9 3 13 2
26 1 1 0 9 9 13 9 1 9 9 13 15 3 7 1 9 1 9 13 9 9 2 9 7 9 2
12 9 13 14 9 9 1 9 7 10 0 9 2
10 9 13 2 16 0 13 13 0 9 2
9 0 13 13 15 9 9 0 9 2
10 15 4 3 13 7 13 1 10 9 2
18 1 0 9 0 13 0 15 13 9 9 7 3 13 7 9 1 9 2
10 1 15 3 13 0 9 1 9 13 2
9 13 3 1 9 9 1 0 9 2
39 13 3 7 12 9 2 16 15 10 9 1 0 9 13 1 11 3 0 7 0 9 9 1 9 9 2 15 15 13 1 9 9 3 2 3 13 10 9 2
11 15 13 9 9 1 12 9 1 0 9 2
27 0 9 13 7 1 10 9 9 7 9 9 9 2 1 15 13 3 0 9 9 2 3 9 2 1 9 2
23 0 11 2 15 15 13 10 9 3 3 2 13 9 9 1 0 9 1 0 9 9 9 2
13 10 9 13 0 9 9 1 9 15 9 7 9 2
16 0 9 13 13 15 7 13 9 9 9 1 0 0 9 9 2
19 0 13 13 9 2 16 4 15 1 9 13 7 13 3 1 0 9 9 2
33 13 4 15 3 13 2 16 16 1 15 13 10 9 9 9 2 1 0 0 9 13 9 1 9 0 7 7 0 7 1 0 9 2
3 1 0 2
4 0 9 1 11
8 11 13 2 16 15 13 9 9
41 2 12 9 4 13 9 7 3 4 15 13 1 0 9 2 2 13 15 1 10 9 11 11 2 0 9 0 9 7 1 9 9 9 11 1 9 0 7 0 11 2
20 1 0 9 2 15 15 3 13 1 9 2 15 15 13 3 2 13 2 11 2
49 1 9 2 1 15 13 1 0 9 2 1 0 9 15 3 13 2 2 15 1 0 9 3 13 0 9 9 9 2 15 11 11 13 1 11 2 0 9 2 11 2 11 2 11 2 11 7 11 2
10 2 1 9 3 1 0 11 13 15 2
20 1 9 0 9 13 1 9 9 12 1 15 3 1 11 1 12 9 1 0 2
19 7 1 12 9 13 1 11 7 0 9 1 9 2 2 13 11 2 11 2
8 9 1 11 13 9 0 9 2
13 1 0 0 9 12 9 15 9 15 13 3 9 2
8 3 3 1 10 9 13 9 2
7 1 11 15 3 13 9 2
17 0 9 12 0 9 15 1 0 9 13 13 14 1 12 9 3 2
11 11 13 3 7 1 9 1 9 0 11 2
8 7 1 9 10 9 3 13 2
11 11 2 11 13 2 2 3 15 15 13 2
17 14 15 2 7 0 9 9 0 11 4 13 1 9 9 1 11 2
15 3 4 13 1 0 9 0 0 9 1 9 1 0 9 2
22 7 13 4 3 9 7 1 10 9 0 7 0 9 13 3 9 1 9 10 9 2 2
6 9 13 13 1 11 2
19 7 7 13 11 1 0 9 1 9 0 9 1 12 7 12 9 0 9 2
25 11 2 11 13 7 3 0 2 2 1 0 4 13 1 12 9 9 2 3 15 13 1 12 9 2
27 7 1 1 15 2 16 9 13 9 3 2 16 4 13 2 13 3 9 2 3 15 13 1 9 12 2 2
1 3
13 0 9 0 9 15 13 3 1 9 9 0 9 2
25 1 9 12 13 1 0 9 13 1 12 5 0 0 9 7 1 12 9 0 9 3 16 1 9 2
4 9 9 13 9
9 9 9 0 9 13 13 1 0 9
23 9 0 9 0 9 2 15 13 0 0 9 2 13 9 9 2 9 3 0 9 9 9 2
32 1 9 11 11 11 13 9 0 9 1 3 0 9 2 15 15 13 1 9 0 9 9 1 0 9 7 9 0 9 0 9 2
28 2 9 0 0 9 4 13 3 1 3 0 9 1 9 0 9 13 1 9 2 15 13 9 9 7 10 9 2
18 3 16 1 0 9 13 1 9 2 9 7 9 7 1 10 9 9 2
26 1 10 9 4 13 13 16 9 2 0 9 2 7 7 1 0 7 0 9 2 2 13 11 2 11 2
20 9 0 9 3 16 9 0 9 13 1 10 9 13 3 9 9 1 0 9 2
23 13 3 1 9 9 0 0 9 2 9 9 9 1 0 9 7 9 0 9 1 9 9 2
29 2 3 0 9 9 11 13 1 9 1 3 0 0 9 3 0 9 2 15 13 0 9 2 2 13 11 2 11 2
32 1 0 9 3 9 2 16 10 0 9 13 0 1 9 2 11 2 11 13 2 16 9 15 13 12 9 1 0 9 7 9 2
28 2 1 9 0 9 9 7 9 1 11 7 0 9 13 13 7 9 0 9 7 9 9 2 2 13 9 11 2
48 1 0 9 1 9 0 9 1 9 12 4 0 11 2 7 3 7 11 7 11 2 13 2 16 13 9 1 0 7 0 9 14 1 9 1 12 7 3 9 2 3 1 12 7 3 9 2 2
29 9 9 10 9 1 9 9 1 9 1 12 9 1 9 12 4 7 13 9 0 0 9 9 1 0 7 0 9 2
25 2 1 0 9 10 0 7 0 9 13 1 0 9 0 0 9 1 9 0 9 0 9 7 3 2
44 11 15 13 0 10 9 7 4 15 15 3 13 2 7 1 9 15 13 1 3 0 9 2 15 3 16 1 0 9 13 0 3 13 1 0 0 9 2 2 13 11 2 11 2
5 0 9 11 1 9
2 11 2
36 0 0 9 11 1 0 0 7 0 9 1 11 13 12 2 9 0 9 9 1 0 9 7 3 0 9 1 9 9 9 7 0 9 1 9 2
17 1 11 11 1 11 13 0 0 9 3 0 2 15 4 3 13 2
23 0 0 9 13 0 9 7 13 3 1 3 0 9 9 1 0 9 2 0 9 7 9 2
20 1 0 9 4 13 4 13 3 14 12 10 9 1 0 9 1 0 9 11 2
4 9 9 1 9
2 11 2
31 9 0 9 0 9 1 9 2 0 11 2 11 2 13 9 0 9 0 9 2 15 15 1 11 13 2 1 9 0 9 2
13 1 0 9 7 9 4 13 4 13 16 0 9 2
33 3 13 9 9 1 9 9 9 11 11 2 0 9 11 13 0 9 9 9 11 1 9 12 1 9 9 0 1 9 12 1 11 2
7 9 13 1 9 11 12 2
20 15 13 14 9 9 2 7 13 3 13 7 13 9 15 9 1 9 7 9 2
22 11 2 11 13 2 16 9 0 9 9 13 9 1 0 9 0 9 1 9 2 11 2
10 1 9 4 15 13 13 9 0 9 2
17 10 9 13 9 3 1 9 0 7 9 0 2 3 3 0 9 2
11 3 13 0 13 1 0 9 7 0 9 2
19 1 11 4 13 4 1 11 13 3 0 0 0 9 0 9 2 11 2 2
14 10 0 9 13 1 9 11 1 0 9 1 0 9 2
12 9 4 13 0 9 2 9 7 0 0 9 2
1 9
14 9 0 9 1 9 1 9 13 0 0 9 1 11 2
40 9 12 2 9 13 13 9 1 9 2 12 2 9 1 9 9 2 9 7 9 2 12 2 9 1 9 0 1 0 9 7 12 2 9 1 9 7 9 9 2
23 0 9 2 9 2 0 9 12 2 12 12 11 2 9 2 2 12 2 12 2 9 12 2
27 0 9 1 0 9 13 1 12 2 2 12 2 9 9 9 11 1 9 1 9 9 9 1 11 1 11 2
18 9 13 9 15 0 9 1 9 9 9 7 9 1 9 9 0 9 2
11 9 4 13 0 9 2 0 9 13 9 2
16 0 9 12 9 1 0 9 13 9 9 1 0 9 1 9 2
37 0 9 2 9 9 11 2 9 2 9 2 0 2 2 9 12 2 0 12 2 12 12 11 1 11 2 9 2 12 2 12 2 9 12 2 12 2
4 1 0 0 9
8 11 11 11 2 13 1 9 2
14 9 9 9 9 2 9 0 11 2 12 9 2 2 2
26 9 0 0 9 13 0 9 2 3 13 9 2 3 13 1 9 1 9 7 3 15 13 0 0 9 2
17 13 15 0 9 1 9 7 9 7 13 2 3 13 9 7 9 2
29 13 7 1 9 13 9 9 1 9 1 0 9 1 9 9 1 0 9 1 0 0 2 0 2 0 7 0 9 2
15 9 13 9 0 9 1 0 9 0 9 1 0 0 9 2
14 11 11 2 9 2 9 0 11 2 12 9 2 2 2
23 0 9 0 9 13 0 9 0 7 0 9 1 9 1 0 9 14 1 9 9 1 9 2
39 13 3 15 1 15 2 15 1 9 1 0 9 13 2 7 3 15 13 1 9 2 15 13 1 9 9 0 9 9 2 9 7 9 1 0 9 9 9 2
21 9 13 0 9 1 9 9 7 1 10 9 0 1 9 2 7 1 0 9 11 2
18 7 13 9 2 15 15 13 1 0 0 9 2 3 0 7 1 9 2
11 13 9 9 2 16 3 13 7 10 9 2
3 11 1 9
1 9
2 9 2
20 9 0 0 9 9 2 11 2 3 13 2 16 1 9 15 11 13 0 9 2
28 15 2 15 1 9 13 1 15 2 13 13 1 9 2 13 1 0 0 9 11 11 2 15 13 9 9 11 2
31 0 9 0 9 0 9 0 9 9 13 2 16 0 9 13 12 9 1 12 9 2 1 15 15 1 9 13 0 9 9 2
13 11 10 9 13 9 2 2 9 13 0 9 2 2
16 9 11 13 2 16 9 11 3 13 0 9 0 9 0 9 2
11 0 9 1 12 0 9 7 3 4 13 2
14 3 1 3 12 1 12 0 9 9 13 0 0 9 2
9 0 9 13 13 1 0 9 9 2
3 3 1 11
3 0 0 9
8 9 11 16 9 1 9 0 9
17 2 2 1 9 13 12 9 2 2 13 9 0 9 1 11 2 2
23 0 9 0 9 9 11 11 7 11 11 2 3 1 9 2 15 15 13 13 9 0 9 2
6 13 1 15 0 9 2
4 9 1 12 9
26 0 9 9 2 0 9 9 2 3 3 4 13 0 13 9 10 9 3 2 16 13 1 9 0 9 2
34 9 4 13 3 1 0 9 2 9 13 1 9 9 3 14 3 2 9 9 1 15 13 3 9 9 13 2 9 1 9 13 3 9 2
9 9 13 9 7 13 13 1 15 2
2 0 9
58 1 9 4 13 10 9 9 2 3 15 0 13 13 9 9 1 9 10 9 15 2 16 13 9 9 7 9 2 3 15 3 13 1 9 0 9 13 9 9 2 13 15 11 11 2 0 0 9 0 9 11 12 2 3 9 0 9 2
10 7 15 15 1 15 3 13 15 9 2
11 15 3 13 7 0 15 13 3 1 9 2
14 9 13 0 13 9 9 2 7 13 1 15 10 9 2
10 13 13 9 7 13 15 1 10 9 2
8 1 10 9 7 13 10 9 2
9 7 13 2 14 15 9 1 9 2
4 13 15 0 2
17 9 13 9 9 9 9 2 7 13 9 2 3 15 1 15 13 2
4 13 15 13 2
3 9 13 2
14 9 13 9 9 2 15 3 1 9 0 13 7 13 2
10 9 15 13 13 7 0 9 13 3 2
7 13 9 2 3 9 13 2
5 1 9 9 1 9
21 1 11 2 11 15 3 13 1 9 2 3 15 0 13 13 0 9 1 9 9 2
9 14 1 11 12 13 15 12 9 2
12 9 13 9 0 9 2 16 9 13 9 9 2
13 1 9 15 13 13 1 15 0 0 9 1 9 2
9 15 7 1 10 9 13 3 0 2
11 11 2 11 4 14 9 1 9 0 13 2
9 1 9 15 9 1 9 3 13 2
8 10 9 9 9 15 3 13 2
18 9 2 13 0 9 1 9 0 0 9 2 15 13 9 1 9 3 2
3 15 3 2
40 2 13 4 15 1 9 2 15 4 3 9 1 9 7 9 3 13 7 13 7 0 9 9 13 9 2 13 2 14 10 9 2 16 3 13 3 1 9 0 2
9 3 15 13 1 9 1 0 9 2
20 13 7 2 16 9 13 10 9 1 3 0 2 16 4 15 15 3 13 2 2
5 15 9 0 9 2
5 15 1 15 9 2
25 1 0 9 4 13 2 16 1 0 9 13 10 9 3 0 7 3 15 1 9 13 1 3 0 2
21 12 9 13 2 16 16 9 13 1 9 9 1 10 9 2 3 3 9 13 9 2
32 1 0 9 15 15 13 13 0 9 2 0 1 11 2 11 7 11 2 11 1 11 7 11 2 11 7 11 2 11 1 11 2
19 9 13 1 9 1 9 13 3 2 11 11 13 3 1 10 9 0 9 2
2 9 9
47 11 2 11 2 15 2 16 13 0 9 2 13 0 9 2 0 9 15 13 3 2 3 2 15 7 13 2 16 1 9 13 1 9 2 15 13 13 2 13 13 2 7 3 13 0 9 2
14 9 2 9 7 9 1 12 9 0 13 1 0 9 2
20 9 3 9 1 9 15 4 1 15 13 1 0 9 14 1 12 2 12 9 2
8 1 10 0 9 13 13 9 2
39 13 15 13 1 9 2 16 4 0 9 13 9 9 2 1 15 15 3 0 9 13 1 9 9 7 0 9 2 3 9 1 9 9 13 13 3 7 9 2
15 13 3 2 1 9 9 1 12 9 9 1 9 1 9 2
24 13 4 2 16 4 15 1 9 9 13 9 9 9 2 15 4 13 0 9 1 9 1 9 2
11 13 15 1 9 1 9 9 1 0 9 2
16 13 13 1 9 2 16 4 13 1 9 3 10 10 0 9 2
44 9 9 2 15 4 12 12 9 1 10 9 13 16 0 7 0 2 4 9 3 13 1 9 2 16 4 15 15 15 13 2 13 15 3 0 9 16 0 9 2 3 13 9 2
27 13 13 15 2 16 4 15 0 9 13 2 16 4 9 13 13 3 7 16 4 15 9 13 1 0 9 2
4 1 2 9 2
15 13 4 15 13 9 2 16 15 0 9 9 13 1 9 2
26 7 0 9 1 0 0 9 15 1 9 13 1 9 2 15 3 1 9 13 9 1 9 10 0 9 2
6 1 9 4 15 13 2
2 11 11
2 9 2
3 11 7 11
2 11 2
27 11 7 0 9 4 13 0 9 1 9 1 0 9 2 15 15 13 13 12 2 2 12 2 9 1 11 2
7 13 15 3 0 9 11 2
25 11 7 11 4 3 1 11 13 0 9 0 15 0 9 2 11 7 11 4 13 9 1 9 9 2
36 0 9 15 13 1 9 11 2 11 2 11 7 0 0 2 0 9 13 7 0 0 9 2 0 11 2 11 2 11 2 11 2 11 7 0 2
21 1 1 9 1 9 11 15 13 9 2 16 15 0 9 9 4 13 3 1 11 2
14 0 9 1 11 11 11 1 9 9 7 9 9 13 2
2 15 9
2 11 2
28 9 1 0 0 9 13 1 12 2 9 12 3 9 9 1 0 9 7 0 9 2 7 15 1 9 12 9 2
20 9 2 15 13 0 9 1 9 1 0 9 2 13 9 1 9 12 9 3 2
10 15 7 13 13 0 9 1 9 11 2
15 3 15 13 9 0 0 9 1 9 12 9 3 0 9 2
13 9 13 1 0 9 1 0 9 9 1 9 12 2
1 9
2 11 2
32 0 9 1 10 0 9 12 2 9 13 9 1 9 0 1 9 9 2 9 7 9 0 9 7 9 0 1 10 9 1 9 2
26 1 9 15 3 2 13 2 16 9 1 9 13 0 13 1 9 1 9 9 9 1 12 2 9 12 2
9 0 9 13 13 7 1 10 9 2
20 9 9 1 9 9 9 0 9 1 9 11 13 0 12 2 12 12 11 12 2
5 12 9 1 9 2
2 11 2
51 1 9 9 2 3 13 0 2 16 0 9 4 13 2 13 9 1 0 9 2 13 9 0 9 9 11 11 7 13 2 13 2 16 4 10 9 4 13 9 2 16 13 2 16 15 4 13 13 1 9 2
13 0 9 11 1 0 0 9 13 14 12 9 9 2
17 0 9 2 11 7 11 13 2 16 13 9 2 15 1 15 13 2
13 9 1 9 0 9 0 0 9 7 3 13 13 2
13 9 1 0 9 13 3 0 0 9 7 0 9 2
21 1 11 2 11 4 13 0 13 15 2 16 10 9 13 0 9 1 9 0 9 2
11 1 9 2 15 13 2 4 15 13 13 2
18 9 0 0 9 2 1 9 2 13 9 0 0 9 7 13 10 9 2
10 2 9 1 11 1 12 2 9 2 2
4 9 11 2 11
9 0 9 9 13 9 1 10 9 2
8 13 15 15 7 1 9 9 2
5 9 11 11 2 11
1 0
34 0 9 3 13 10 9 2 13 1 9 9 2 13 9 7 9 0 9 2 13 15 9 1 9 7 13 2 10 9 13 9 1 9 2
17 1 0 9 13 1 11 11 1 0 9 10 9 1 11 11 11 2
34 14 3 0 9 13 1 9 7 1 9 13 11 16 15 2 15 15 13 2 7 15 13 2 16 1 9 13 13 9 2 15 15 13 2
15 3 15 1 9 3 13 2 13 13 2 16 11 13 9 2
26 6 2 10 0 11 2 13 15 2 3 3 13 1 10 9 2 12 9 0 9 2 15 13 3 0 2
19 0 0 11 1 12 2 9 13 0 9 2 13 11 2 3 13 3 3 2
6 3 1 10 0 11 2
9 13 0 7 9 3 13 0 9 2
21 0 0 9 3 13 7 13 4 15 3 1 9 13 11 2 16 4 13 3 9 2
18 13 0 2 13 11 2 16 4 0 11 13 10 0 9 1 0 11 2
12 10 9 1 11 13 13 15 1 9 0 11 2
16 3 15 13 1 0 11 1 9 9 2 9 2 9 2 9 2
11 14 11 1 9 2 0 9 2 13 3 2
17 0 9 0 0 9 13 3 3 0 9 9 9 2 9 7 9 2
27 13 3 3 0 13 2 16 11 2 11 7 11 15 13 0 9 1 15 2 16 4 3 13 1 10 9 2
15 13 3 0 9 1 15 2 16 11 3 1 15 0 13 2
7 9 0 11 13 3 0 2
16 13 1 0 9 1 15 2 15 15 1 9 13 1 0 9 2
58 11 2 11 7 11 2 10 3 0 2 7 16 3 0 9 0 11 13 2 3 15 13 2 0 9 0 9 3 16 0 9 2 3 9 9 11 2 11 11 2 11 11 7 0 0 9 0 7 0 11 1 0 9 3 3 3 13 2
11 7 1 10 9 11 2 9 2 3 13 2
4 13 7 13 2
2 11 11
5 9 13 2 13 11
2 11 2
10 0 0 9 13 1 9 9 11 11 2
26 9 9 0 9 11 11 11 1 0 9 0 9 0 2 11 13 9 2 2 16 4 13 1 9 2 2
21 11 3 13 2 16 15 10 9 0 9 0 9 11 13 1 9 1 0 0 9 2
32 0 9 1 0 11 7 9 2 0 3 1 9 9 2 13 3 1 9 1 9 0 9 1 9 1 0 9 1 9 11 11 2
5 10 9 4 13 2
7 9 1 9 9 0 9 2
6 16 13 9 2 2 2
5 11 2 11 2 2
31 0 9 1 11 4 0 9 13 9 0 9 11 1 0 9 1 9 9 0 9 0 9 9 2 5 0 11 5 11 2 2
7 9 15 7 3 3 13 2
8 9 9 11 3 13 0 9 2
14 13 3 1 9 0 0 9 2 15 13 0 0 9 2
24 2 9 4 13 2 15 13 9 13 2 2 13 9 2 11 2 11 2 9 9 9 11 11 2
20 2 3 13 13 2 16 1 0 9 13 12 9 2 16 15 9 13 13 2 2
31 9 0 9 13 2 16 0 0 9 2 13 9 10 9 13 2 2 2 4 13 3 14 13 1 9 1 9 9 11 2 2
12 3 13 2 16 9 13 3 0 9 3 13 2
29 1 0 9 1 11 12 9 9 13 1 15 2 16 4 9 13 0 9 3 10 9 2 3 13 9 9 7 9 2
23 0 9 3 13 9 1 10 9 0 9 2 1 0 9 1 9 9 2 7 1 9 9 2
10 9 7 9 13 16 2 3 0 2 2
42 10 9 1 11 12 14 13 13 0 9 1 0 9 0 9 2 1 10 9 11 13 9 2 16 15 13 3 0 13 9 9 2 1 9 0 11 3 13 2 2 2 2
23 1 9 1 9 13 1 11 3 0 9 2 16 12 1 9 9 13 9 9 11 2 11 2
17 3 2 16 0 9 13 3 13 7 13 2 3 4 7 13 3 2
21 1 0 9 2 9 2 9 9 7 0 9 1 0 9 13 13 0 9 3 0 2
24 0 9 9 7 10 9 13 2 7 1 0 9 2 15 13 9 2 16 15 9 0 9 13 2
29 16 4 3 2 9 11 13 9 0 1 9 7 0 2 9 2 0 1 0 9 2 13 4 9 13 0 9 2 2
29 3 1 9 9 9 2 11 16 9 3 3 3 13 1 9 9 9 7 9 9 2 2 2 9 1 12 9 2 2
3 1 9 2
2 11 2
23 1 10 9 13 3 0 9 1 0 11 1 0 0 9 2 1 15 15 9 13 0 9 2
40 0 9 9 11 2 15 13 9 3 12 9 9 2 3 3 13 9 0 9 9 16 1 0 9 2 3 3 12 9 2 2 14 7 0 2 3 1 0 9 2
21 0 9 2 13 2 1 0 9 3 1 11 1 9 9 3 1 9 2 2 2 2
28 0 9 3 3 13 1 9 1 10 9 1 11 2 3 15 3 13 2 7 9 3 3 13 10 9 2 2 2
2 0 9
5 11 2 11 2 2
41 2 9 13 13 3 12 7 3 12 1 15 13 0 9 1 0 9 9 2 2 13 1 0 0 9 9 2 11 9 1 0 9 9 1 9 1 9 9 1 11 2
7 1 9 4 13 0 9 2
20 9 3 13 12 0 9 9 2 15 7 13 2 16 15 1 15 13 1 9 2
20 9 9 1 9 9 13 12 0 9 2 13 3 0 2 3 13 0 0 9 2
8 9 13 7 9 7 9 9 2
22 9 15 0 9 13 12 12 9 2 1 0 9 7 1 15 13 9 13 14 3 3 2
19 13 13 2 16 1 9 4 13 13 0 9 3 1 9 2 3 1 11 2
5 13 15 11 2 11
5 11 2 11 2 2
41 9 12 2 0 9 9 1 9 2 9 7 0 9 11 7 0 9 0 9 2 9 7 9 11 2 15 15 13 1 12 2 1 12 2 9 2 13 1 0 9 2
61 9 12 0 9 4 13 9 9 0 9 2 1 0 3 2 11 2 0 9 7 9 9 1 9 2 2 11 2 0 9 2 2 11 2 9 2 2 11 2 9 2 2 1 0 3 11 2 0 0 9 11 2 9 11 2 11 11 2 11 3 2
26 1 9 9 0 9 11 9 2 11 11 13 9 2 15 15 3 13 13 16 9 2 0 9 15 13 2
3 13 1 9
2 11 2
11 9 13 9 1 9 1 3 12 9 11 2
35 13 15 1 9 0 9 2 1 15 15 1 9 9 7 9 13 9 11 1 9 1 9 1 9 0 9 0 9 11 1 10 9 1 9 2
5 11 1 11 7 11
2 0 9
2 11 2
36 9 0 9 9 7 9 10 0 9 11 11 1 0 0 9 1 11 13 2 16 9 13 13 1 9 1 9 7 0 9 7 1 0 0 9 2
17 13 3 2 16 13 1 0 0 9 2 1 9 9 11 7 11 2
29 13 1 9 1 0 9 13 0 9 1 15 2 16 15 13 1 9 15 2 15 1 9 13 9 7 13 0 9 2
3 13 15 9
3 9 1 11
5 11 2 11 2 2
19 0 9 9 13 1 0 9 9 12 13 0 0 9 1 9 0 0 9 2
14 0 9 9 4 13 9 2 0 4 13 9 0 9 2
21 1 9 10 9 13 11 9 2 9 7 9 7 9 2 15 4 13 0 9 13 2
16 9 9 13 1 9 0 9 0 0 11 7 13 0 0 9 2
18 1 9 0 9 13 11 0 9 7 9 7 13 0 9 2 3 9 2
26 9 1 9 7 9 15 13 13 1 9 0 9 9 2 0 9 2 1 9 12 2 12 12 11 12 2
15 1 9 9 13 3 0 0 0 9 3 1 0 0 9 2
21 12 9 0 9 13 0 9 0 9 11 11 7 9 11 11 1 9 12 7 12 2
18 9 9 11 1 9 1 0 12 9 13 11 7 11 0 7 11 11 2
6 9 2 11 2 11 11
22 0 9 13 12 9 1 9 12 7 12 9 1 9 1 0 9 9 1 11 1 11 2
17 0 9 13 1 9 3 12 9 1 0 9 9 1 11 1 11 2
21 0 0 9 11 13 9 9 12 1 0 2 9 2 9 1 11 1 11 1 11 2
25 9 0 9 13 1 9 3 2 1 11 9 11 11 2 15 0 0 0 9 13 1 9 0 9 2
36 12 9 0 9 1 11 15 13 12 2 0 9 0 2 15 13 0 9 1 0 11 1 9 1 12 2 9 12 1 12 2 9 12 1 11 2
16 0 0 9 0 2 15 13 1 11 2 15 13 1 12 9 2
32 0 9 1 0 9 9 7 9 9 7 0 9 13 1 9 0 9 11 11 1 0 9 0 9 9 1 9 2 0 9 11 2
19 16 9 13 9 2 16 11 2 11 13 1 12 2 9 0 9 0 9 2
23 0 9 1 0 9 13 1 0 9 1 0 9 9 0 9 1 11 1 11 1 12 9 2
18 1 0 9 13 1 11 1 0 9 0 0 9 1 9 1 0 9 2
7 13 4 15 13 12 9 2
20 0 9 9 13 3 1 0 9 3 9 11 11 11 2 11 7 9 1 9 2
18 1 9 9 7 9 13 10 9 0 0 9 9 11 11 1 0 11 2
12 13 4 3 0 0 9 2 12 9 7 9 2
28 0 9 1 9 15 13 2 16 9 10 0 9 13 1 12 7 1 12 9 1 0 9 11 2 1 11 12 2
17 0 9 9 0 9 0 9 13 3 10 9 7 9 9 11 9 2
28 2 9 2 13 0 9 16 9 0 2 13 15 1 15 0 9 2 0 9 2 9 2 0 9 7 0 9 2
18 9 1 9 7 9 2 11 9 2 0 12 2 11 12 2 12 12 2
12 0 9 13 1 9 0 9 7 9 0 11 2
24 9 1 10 9 13 3 9 9 0 9 11 11 11 2 1 9 9 2 9 0 9 11 11 2
21 9 1 11 13 11 7 3 4 13 2 9 0 9 1 0 7 0 0 9 2 2
17 0 9 0 9 9 13 2 16 13 1 9 9 7 9 0 9 2
12 0 9 0 9 9 4 13 9 2 11 11 2
23 0 9 1 9 9 0 9 0 9 2 15 15 13 1 0 9 2 13 9 12 2 9 2
15 13 0 9 2 0 9 7 9 0 9 13 13 0 9 2
7 0 9 0 9 13 0 2
2 9 9
4 2 11 2 2
21 9 13 9 9 2 13 10 9 2 13 4 16 9 12 9 1 0 9 1 9 2
7 7 9 15 15 3 13 2
22 13 4 15 1 10 9 2 16 4 1 0 9 9 11 13 0 9 2 0 9 2 2
31 1 11 3 13 1 10 9 2 14 2 1 12 9 9 9 2 0 9 2 12 9 2 7 1 0 9 13 14 12 9 2
15 1 0 9 2 15 9 13 12 2 13 3 15 1 9 2
26 7 3 9 16 1 0 9 9 13 3 9 1 0 9 9 2 3 9 0 2 3 13 9 3 0 2
14 3 13 9 13 15 1 9 1 15 0 3 12 7 2
52 3 15 15 4 10 9 13 3 0 2 7 1 9 2 15 15 3 12 9 13 1 0 9 9 7 9 1 10 2 0 2 9 7 3 1 0 9 9 0 9 2 13 0 9 0 3 14 3 0 7 0 2
11 7 15 3 7 1 15 2 3 1 9 2
3 9 9 2
5 2 9 4 13 2
5 11 2 11 13 9
5 11 2 11 2 2
56 11 11 2 9 1 0 11 2 13 12 2 9 9 2 15 13 1 12 9 12 2 9 12 2 16 15 12 2 9 0 9 11 11 11 13 2 16 15 4 3 13 2 3 13 9 9 7 9 0 0 9 1 9 2 12 2
14 16 9 10 9 13 2 13 15 11 2 11 9 13 2
85 3 13 2 16 4 11 11 3 7 1 9 13 10 9 1 12 2 12 2 12 7 16 4 0 9 2 0 7 0 2 13 13 1 10 0 9 1 12 2 12 2 12 2 7 0 9 15 3 13 2 2 7 1 0 9 0 9 0 9 11 1 12 2 12 2 12 0 2 9 2 12 2 12 9 12 2 12 13 1 9 1 0 9 2 2
36 11 2 11 13 7 1 15 2 16 15 9 13 9 2 15 13 2 7 13 2 16 4 0 9 9 9 10 0 9 3 13 7 13 0 9 2
2 0 9
5 11 2 11 2 2
13 1 12 2 9 13 1 11 0 9 0 9 11 2
33 9 13 9 9 11 7 1 9 13 9 7 9 2 15 9 13 2 7 15 2 15 15 15 13 1 9 9 1 9 9 7 9 2
16 0 9 4 9 13 2 13 0 0 9 7 13 0 0 9 2
10 1 10 9 13 7 9 0 0 9 2
2 9 11
92 0 9 2 9 7 9 2 13 2 16 15 1 0 9 13 1 10 0 9 2 15 13 1 11 1 9 12 2 7 1 10 9 2 15 13 1 9 1 0 0 9 2 14 3 0 9 2 15 15 1 9 13 0 9 2 16 0 10 9 4 15 13 7 9 2 2 0 9 9 7 9 2 0 9 0 0 9 11 0 7 9 1 9 1 0 9 2 9 7 9 11 2
16 13 15 1 0 9 3 3 0 9 1 9 10 9 7 9 2
15 3 9 2 9 7 9 1 0 9 15 13 9 0 9 2
13 9 11 2 0 12 2 12 12 11 12 2 11 12
14 9 12 2 12 2 12 2 12 2 12 9 12 2 12
4 0 9 15 13
2 11 2
16 0 9 11 15 1 9 1 9 9 1 9 1 10 9 13 2
20 10 0 9 13 2 13 3 9 0 9 0 9 7 9 9 9 9 11 11 2
18 9 0 9 13 3 1 10 9 10 9 1 10 9 1 3 0 9 2
10 0 9 3 13 14 1 0 0 9 2
2 0 9
11 1 0 0 9 13 9 11 1 0 9 2
23 9 9 15 13 1 0 9 1 0 9 1 11 9 1 11 7 13 15 9 0 0 9 2
18 1 11 1 9 11 13 1 0 9 3 9 9 9 9 1 0 9 2
14 13 0 9 2 9 2 0 9 2 9 7 0 9 2
6 9 13 9 12 9 2
22 12 2 9 13 12 0 9 1 9 12 7 12 9 1 11 11 1 11 1 9 11 2
13 1 9 3 13 0 12 9 0 9 1 11 11 2
1 9
16 1 12 9 2 3 1 9 2 13 9 2 9 0 2 11 2
12 0 9 2 15 13 9 1 9 1 0 9 2
27 13 15 0 9 2 4 13 1 11 2 3 7 1 11 7 3 1 0 9 1 11 2 3 1 9 13 2
7 1 9 13 1 0 9 2
10 1 12 9 13 1 0 9 9 12 2
19 1 9 12 13 1 12 9 0 9 13 1 0 9 1 0 9 0 9 2
9 13 15 1 11 7 13 0 9 2
24 16 0 9 11 15 13 9 1 9 2 13 10 9 7 9 2 13 9 1 9 0 9 11 2
6 15 4 13 2 13 2
18 9 1 9 15 0 9 13 1 9 11 11 7 10 9 1 0 9 2
7 15 13 10 0 0 9 2
3 2 11 2
3 9 9 13
2 11 2
25 9 9 11 1 9 0 9 11 2 15 4 13 13 9 1 0 9 11 7 11 2 13 0 9 2
31 1 0 9 13 3 9 11 7 11 2 10 9 13 3 1 3 0 9 9 3 9 9 11 2 3 9 0 9 11 12 2
27 9 9 11 11 11 3 13 2 16 13 9 9 2 15 13 0 9 2 7 3 15 15 9 0 9 13 2
31 1 0 13 2 16 15 3 13 10 9 7 16 15 13 15 13 2 16 4 15 11 13 0 0 9 0 9 0 9 9 2
4 0 9 0 9
7 0 9 11 2 11 2 2
13 0 9 13 9 7 9 1 0 0 9 1 11 2
31 0 0 9 15 3 3 13 7 1 0 9 2 9 7 9 9 11 11 15 13 1 9 0 0 9 13 7 9 3 0 2
17 16 4 3 13 1 9 2 13 4 15 1 9 1 0 0 9 2
24 2 9 10 9 3 13 2 1 9 13 10 9 2 7 13 4 0 15 1 15 13 1 0 2
22 3 0 9 13 12 7 12 9 0 9 2 14 1 9 0 1 12 9 1 9 2 2
23 10 9 15 1 0 0 9 3 13 1 9 0 9 9 2 1 9 7 0 9 0 9 2
10 3 15 9 1 10 2 9 2 13 2
16 2 13 2 7 3 13 0 9 9 13 1 10 9 3 0 2
15 0 0 9 1 0 9 13 0 13 15 1 9 1 9 2
9 13 15 1 15 2 3 3 13 2
23 13 1 9 9 2 13 3 1 9 0 7 3 0 9 2 1 9 3 13 11 11 2 2
16 0 0 9 13 3 3 1 9 9 2 7 13 15 3 2 2
5 9 1 9 7 9
2 11 2
23 0 0 9 1 0 9 1 11 0 0 0 0 2 9 13 0 9 1 0 9 9 12 2
11 9 9 13 9 1 9 9 12 7 12 2
34 1 9 13 13 3 0 0 9 9 1 12 9 2 0 9 0 9 7 0 9 9 1 0 7 0 2 15 13 14 1 0 9 0 2
26 11 13 1 12 2 12 14 1 12 2 12 9 9 7 9 2 15 13 0 9 9 2 9 2 9 2
23 1 0 9 13 13 11 11 1 0 0 9 9 7 3 14 1 12 9 9 0 9 11 2
11 9 0 0 9 13 9 1 11 7 11 2
8 3 15 4 13 0 12 9 2
22 1 0 11 4 13 0 0 9 2 15 1 9 1 0 9 13 9 7 12 0 9 2
11 1 0 9 13 3 7 9 1 0 9 2
24 1 0 9 13 13 9 9 1 9 0 9 9 1 9 2 9 9 0 11 11 7 0 9 2
22 9 3 13 0 9 1 0 9 11 11 7 9 11 11 1 0 0 11 1 0 9 2
3 9 1 11
2 11 2
34 3 13 9 9 0 9 9 1 11 9 2 11 11 2 4 12 2 9 1 12 9 13 0 9 1 9 11 1 9 11 2 0 9 2
28 1 9 13 1 10 9 9 11 1 12 9 2 15 13 0 9 1 9 9 7 13 9 1 9 3 12 9 2
14 9 1 9 7 9 3 13 7 1 9 13 9 9 2
9 9 0 12 9 13 9 10 9 2
32 14 1 15 3 1 0 9 4 13 9 0 9 2 15 15 12 0 9 2 0 9 9 12 9 7 0 0 9 13 13 11 2
16 9 13 12 1 9 13 1 9 0 9 7 7 1 9 13 2
12 1 9 13 9 2 15 13 1 9 0 9 2
18 12 1 9 15 13 3 13 2 0 7 13 1 9 13 1 12 9 2
9 15 9 13 2 7 13 4 15 2
17 1 0 9 0 1 0 9 13 0 9 9 2 0 9 1 11 2
3 3 1 9
20 1 12 9 15 13 1 0 9 2 1 12 2 9 2 3 13 0 9 11 2
24 1 10 9 13 13 7 12 9 2 15 13 1 12 9 7 12 9 2 10 9 13 13 3 2
11 0 9 0 9 0 2 0 9 1 0 9
19 0 9 0 11 13 3 3 0 9 9 11 11 2 11 11 2 9 2 2
11 9 15 1 11 13 9 0 9 11 11 2
5 9 11 11 2 11
4 1 11 13 11
4 11 1 11 2
27 0 0 9 4 1 9 2 16 4 15 3 13 9 2 13 12 9 2 15 13 3 9 1 11 1 11 2
13 1 9 10 9 15 9 11 3 13 1 12 9 2
20 1 0 9 4 15 13 11 1 12 9 2 15 13 9 1 9 1 12 9 2
33 3 13 1 0 9 9 2 15 13 3 0 9 11 1 11 1 11 2 13 0 9 0 11 2 1 15 4 3 13 12 9 9 2
8 1 9 15 13 3 12 9 2
32 0 9 1 9 13 1 11 1 11 11 2 11 2 15 3 13 1 9 13 1 12 9 9 2 3 7 3 3 1 12 9 2
3 1 9 9
2 11 2
21 3 13 0 9 1 9 0 9 1 11 2 11 2 3 15 13 10 9 12 0 2
31 1 0 9 1 9 1 15 13 9 0 1 11 2 15 1 11 13 9 9 2 7 13 15 9 1 9 7 0 0 9 2
8 3 0 0 15 13 13 9 2
6 9 2 9 2 2 2
5 11 2 11 2 2
22 9 0 9 7 9 9 13 1 9 11 1 0 9 9 1 9 9 2 9 2 9 2
25 9 15 13 13 9 9 2 0 9 2 9 1 9 0 9 2 9 2 0 9 2 9 7 9 2
28 0 9 13 0 9 2 15 13 13 3 1 9 12 7 0 15 3 13 13 1 0 9 1 9 9 9 9 2
21 9 13 13 0 9 1 12 2 9 7 13 0 2 9 0 9 13 7 1 9 2
7 1 9 1 0 9 1 11
8 2 1 9 15 13 9 2 2
33 9 1 11 9 1 11 4 13 1 9 2 9 7 9 3 3 2 3 15 13 2 7 3 13 2 2 1 12 10 9 11 11 2
31 13 4 9 0 1 0 9 1 0 7 0 0 9 1 10 9 1 9 9 1 11 1 0 9 2 1 15 13 9 9 2
31 16 1 9 4 13 2 16 3 9 2 3 14 3 15 1 0 9 11 11 9 2 2 9 15 13 2 7 3 2 13 2
9 2 2 2 2 2 13 3 3 2
8 2 13 4 15 1 0 9 2
5 2 1 0 9 2
5 2 13 3 9 2
6 2 13 3 13 9 2
7 2 13 0 9 2 9 2
4 2 0 9 2
9 2 2 2 2 2 3 13 2 2
15 11 13 0 9 9 1 0 9 2 0 1 10 9 9 2
12 3 9 2 9 2 9 2 1 9 3 9 2
11 7 9 3 1 12 9 13 1 9 9 2
15 4 3 13 9 0 9 2 15 13 7 13 13 10 9 2
39 2 3 15 1 9 15 13 2 3 1 15 13 9 1 9 2 2 13 9 11 11 2 1 10 9 1 9 9 9 1 9 12 13 15 16 10 0 9 2
4 13 0 9 2
17 1 0 9 3 13 9 9 7 9 1 9 1 12 1 12 9 2
13 3 15 3 14 13 2 16 1 9 13 12 9 2
21 13 15 2 16 9 1 9 13 3 0 2 3 1 9 1 0 0 9 2 2 2
9 7 13 3 9 7 10 0 9 2
28 3 13 9 9 13 3 2 3 7 1 0 9 2 13 13 10 9 1 9 7 3 15 7 13 9 1 15 2
14 1 15 2 3 2 2 7 2 3 1 9 2 3 2
5 9 10 9 13 2
12 1 9 15 7 9 1 0 9 9 15 13 2
8 13 15 3 16 0 0 9 2
16 7 12 9 1 0 9 15 1 0 9 3 13 3 3 3 2
17 9 9 1 10 9 13 1 9 9 2 7 15 13 3 0 9 2
17 1 9 13 9 0 9 7 2 9 2 3 13 1 10 0 9 2
7 1 15 9 13 0 9 2
26 1 9 1 15 1 0 2 9 2 13 9 7 3 7 0 9 2 15 14 13 1 15 9 0 2 2
34 2 16 3 13 0 9 2 13 4 1 15 9 2 16 4 15 9 15 9 13 2 13 15 3 3 1 9 1 9 2 2 13 15 2
14 7 3 0 9 2 2 1 9 15 13 13 9 2 2
24 1 0 9 15 13 9 9 1 10 0 9 3 3 13 2 10 9 2 9 1 3 0 9 2
5 3 13 15 3 2
10 2 13 15 9 1 9 16 0 13 2
16 7 16 13 9 3 3 1 9 2 3 14 13 15 10 9 2
15 7 3 2 16 3 3 2 13 15 9 0 9 3 2 2
10 2 7 2 3 2 2 2 2 2 2
38 3 9 0 13 9 2 3 15 7 15 2 9 3 0 7 3 3 0 2 3 13 1 10 0 2 15 10 0 9 3 7 3 2 3 7 3 13 2
18 0 9 7 9 1 3 0 9 2 16 13 15 1 11 2 13 0 2
2 11 11
4 1 10 0 9
20 9 9 11 1 10 12 2 9 13 0 9 9 0 9 2 10 9 13 9 2
24 1 0 9 9 13 0 9 13 1 9 1 9 9 2 9 9 2 7 13 15 1 9 9 2
15 9 3 13 9 13 2 9 1 9 2 15 9 9 11 2
32 10 9 13 1 9 1 9 9 11 1 9 12 2 15 9 13 13 0 9 1 9 11 7 13 3 0 9 11 1 10 9 2
12 0 9 13 13 9 9 12 9 1 9 9 2
9 10 9 4 13 3 1 0 9 2
11 3 13 0 2 16 0 9 10 9 13 2
2 11 11
23 1 0 9 1 9 13 0 9 3 3 12 2 9 1 9 9 9 9 1 11 9 9 2
13 0 9 9 9 13 9 1 9 7 13 1 9 2
4 15 4 13 2
16 1 9 2 15 1 9 13 7 1 9 9 13 2 15 13 2
2 11 11
3 13 1 9
2 11 2
38 1 3 0 9 13 13 7 13 15 2 16 4 13 1 9 12 3 13 0 9 1 0 9 0 9 1 9 12 2 13 3 9 0 9 11 11 11 2
10 1 10 9 4 13 7 10 0 9 2
9 3 13 9 1 0 3 0 9 2
11 0 9 15 13 9 0 9 1 0 9 2
33 1 9 0 9 9 11 11 11 1 10 0 9 4 13 9 0 9 11 11 13 0 0 9 0 1 0 9 9 9 11 11 11 2
10 1 11 13 4 13 9 1 9 9 2
26 1 0 0 9 3 13 0 9 2 1 15 15 9 13 2 16 15 13 0 0 9 9 1 10 9 2
12 3 7 13 0 0 9 10 0 9 9 12 2
6 9 1 11 9 11 11
3 2 11 2
15 9 11 13 0 9 0 9 1 9 0 9 12 0 9 2
15 13 15 2 16 12 1 9 10 9 13 3 9 11 11 2
23 13 1 9 11 1 15 2 16 0 9 12 1 9 7 9 1 9 13 9 10 0 9 2
13 7 13 2 14 12 15 2 13 15 13 3 15 2
30 13 15 1 10 9 13 13 15 11 2 11 2 3 15 1 9 9 3 3 13 1 9 0 9 2 15 13 3 9 2
19 3 0 9 3 13 2 7 16 13 1 9 3 2 1 10 9 3 13 2
18 3 13 0 9 1 15 0 2 7 13 9 9 7 9 1 10 9 2
42 13 2 14 15 3 9 11 13 9 0 9 2 1 10 9 15 3 3 3 13 2 13 15 2 16 1 15 13 1 0 9 3 3 3 2 3 4 15 3 3 13 2
35 13 3 13 2 16 16 4 13 0 9 9 10 2 15 15 13 1 9 0 9 2 13 4 15 9 11 13 0 9 7 1 9 9 9 2
3 2 11 2
4 1 11 13 9
2 11 2
24 0 9 13 1 9 1 9 1 9 9 1 11 2 3 15 1 0 9 13 0 9 11 11 2
10 13 15 9 9 11 1 0 0 9 2
20 9 9 13 9 9 2 15 1 9 13 0 9 7 10 9 0 1 0 9 2
20 1 9 3 13 0 9 7 3 9 0 9 0 12 9 9 15 13 1 9 2
9 7 1 0 9 15 1 11 13 2
7 0 9 15 13 1 9 2
11 0 9 15 13 3 12 0 7 9 0 2
17 9 0 0 9 13 1 9 1 9 1 9 9 0 0 9 11 2
31 1 9 4 13 10 0 9 2 1 15 7 12 1 0 9 9 11 11 2 15 4 13 1 9 9 11 11 3 1 9 2
28 12 0 0 9 2 0 3 1 9 1 0 9 2 13 9 9 1 10 9 7 10 9 13 1 2 9 2 2
3 11 1 9
1 9
2 11 2
15 0 9 9 2 11 2 13 9 1 0 0 9 1 11 2
20 1 0 0 9 13 1 0 9 12 9 2 12 9 9 2 1 12 0 9 2
34 9 9 11 11 3 13 2 16 1 3 0 9 1 12 0 9 13 1 0 9 9 13 12 0 9 1 9 2 15 13 0 9 9 2
29 0 11 13 12 9 2 12 9 2 2 9 0 9 12 9 1 9 0 3 0 9 7 0 9 0 9 12 9 2
6 12 9 13 0 9 2
2 11 2
1 11
2 0 9
2 11 2
25 0 9 7 9 4 3 13 1 9 7 10 9 1 9 1 11 4 13 2 16 11 13 10 9 2
18 9 13 9 11 1 9 11 1 0 9 13 13 1 9 9 1 9 2
15 0 9 9 0 9 13 1 0 9 7 13 1 0 9 2
13 1 9 4 13 0 9 7 14 12 0 4 13 2
10 0 0 9 13 1 9 3 1 9 2
15 1 9 0 9 13 11 1 9 12 9 7 13 3 9 2
2 9 2
3 14 1 9
2 11 2
9 9 1 11 13 13 3 0 9 2
7 13 1 15 3 0 9 2
14 9 4 13 12 9 1 9 0 9 0 9 0 9 2
14 1 0 9 13 1 9 12 11 7 12 0 4 13 2
25 0 0 9 9 4 3 13 13 0 9 2 15 13 2 16 0 0 9 11 13 0 0 9 9 2
36 1 0 9 4 1 9 13 12 9 9 0 0 9 11 11 2 9 11 11 15 13 9 9 11 11 7 9 11 11 13 9 9 9 7 9 2
23 0 0 9 0 9 11 11 13 7 3 2 1 9 10 12 2 9 2 0 10 0 9 2
21 16 10 9 4 13 3 1 11 2 15 0 9 13 1 10 9 1 11 1 9 2
21 9 9 11 1 12 0 7 0 9 1 9 3 13 3 1 9 1 0 9 11 2
19 3 16 12 0 13 1 9 2 12 9 7 4 13 2 1 15 12 3 2
20 0 9 3 2 13 2 12 2 9 0 9 1 11 9 12 9 1 9 11 2
10 12 9 3 13 7 12 0 4 13 2
14 0 12 9 9 9 2 9 13 1 0 0 9 11 2
5 13 4 12 9 2
9 0 9 11 11 13 9 1 9 2
16 13 2 16 10 9 13 13 9 0 9 7 3 3 13 9 2
18 9 15 13 9 9 9 2 0 9 2 9 9 0 9 7 0 9 2
22 1 0 9 0 1 9 11 1 11 7 11 13 3 1 0 9 0 9 9 11 11 2
21 13 1 15 9 9 0 1 0 9 1 12 9 7 9 9 9 0 7 0 9 2
28 0 9 11 11 2 11 2 15 4 13 1 12 9 1 0 11 1 0 9 2 4 13 7 13 15 1 11 2
20 1 9 13 2 16 9 1 9 2 13 0 2 2 13 0 9 7 3 13 2
12 13 15 3 13 0 9 7 13 0 0 9 2
23 9 9 13 1 9 1 9 0 0 9 11 11 11 7 10 9 11 1 9 11 1 11 2
11 1 0 9 13 7 9 2 3 0 9 2
15 15 15 3 13 1 3 0 0 9 2 3 1 0 9 2
13 0 9 13 10 0 0 9 1 11 1 12 9 2
28 13 15 3 0 9 1 9 1 0 0 2 0 9 2 1 15 9 13 1 9 1 0 9 2 0 0 9 2
23 1 11 15 3 13 1 0 11 14 12 11 1 0 12 2 13 0 9 9 11 2 11 2
13 1 9 1 0 9 13 15 0 12 9 2 13 2
13 13 3 2 16 3 11 13 1 12 9 1 11 2
17 12 9 4 13 1 9 1 0 0 9 1 9 11 7 1 11 2
5 13 15 0 9 2
20 1 15 13 1 0 9 1 9 0 0 9 7 9 9 2 15 13 9 11 2
25 0 0 0 9 11 11 13 1 9 0 9 1 11 0 9 7 1 15 3 13 7 9 0 9 2
11 13 15 3 9 0 0 9 1 0 9 2
21 0 9 1 0 9 0 9 13 12 0 9 2 15 1 10 9 9 13 0 9 2
29 10 13 10 9 9 1 9 2 13 3 0 2 7 9 2 16 13 1 11 3 0 2 13 0 9 3 0 9 2
28 9 13 1 9 1 9 2 3 15 1 12 1 9 13 0 9 2 15 0 9 3 13 7 9 2 9 13 2
18 3 13 2 16 9 1 10 9 13 9 2 7 16 15 13 0 9 2
2 0 9
2 11 2
18 1 9 0 0 9 1 9 11 0 1 12 9 13 9 9 7 9 2
21 1 10 9 13 9 2 0 9 2 1 0 9 12 2 9 7 13 9 9 0 2
19 0 9 9 7 9 13 3 12 7 12 12 9 1 9 1 0 9 9 2
27 1 9 13 1 9 0 9 13 9 3 0 9 11 2 9 9 9 11 7 0 9 0 9 7 10 9 2
25 0 9 9 2 0 9 7 1 10 9 3 0 9 13 0 9 13 0 9 14 1 9 12 9 2
20 9 11 1 11 1 0 9 11 14 2 1 0 9 0 11 2 13 11 11 2
2 11 2
1 11
2 9 13
2 11 2
25 9 0 9 11 11 15 13 13 1 9 0 9 1 11 2 16 9 11 11 13 1 9 0 9 2
41 1 9 0 9 9 7 9 11 13 2 16 9 1 0 9 7 11 2 15 13 1 15 2 16 1 9 12 0 9 11 11 13 1 11 9 2 2 4 13 2 2
2 9 11
2 13 9
2 11 2
19 11 13 13 1 9 1 9 0 11 2 0 9 1 11 2 1 0 9 2
11 13 15 1 11 0 9 11 11 2 11 2
21 13 2 16 9 11 4 15 13 7 1 9 2 15 13 13 0 9 1 0 9 2
13 0 11 1 9 13 0 9 9 0 0 9 9 2
27 9 11 13 3 9 1 9 2 0 2 9 7 13 9 2 16 10 9 15 13 9 0 9 0 0 9 2
18 1 0 9 13 1 0 0 9 11 7 1 0 9 0 11 0 9 2
4 9 1 0 9
4 11 2 11 2
25 1 0 9 1 9 0 0 9 3 0 9 13 1 9 12 0 9 2 16 13 9 0 0 11 2
27 1 0 13 0 0 9 9 11 11 11 11 2 15 3 13 2 16 4 13 1 9 1 2 0 9 2 2
12 13 15 7 1 0 9 9 0 9 1 9 2
22 1 9 2 15 15 13 1 9 2 4 13 3 0 0 0 9 11 11 7 11 11 2
29 9 1 9 7 9 9 11 2 15 1 0 0 9 13 1 0 9 1 9 1 9 2 15 13 0 12 0 9 2
10 1 9 3 13 1 9 9 12 9 2
6 1 12 9 13 9 2
21 0 9 13 0 9 9 1 9 0 9 2 3 15 1 0 9 3 3 13 11 2
15 1 9 1 11 1 9 9 13 10 9 1 0 11 9 2
11 1 9 15 3 13 0 9 12 0 9 2
3 9 1 9
3 9 1 9
2 11 2
22 3 12 9 1 9 0 2 0 9 2 13 3 1 9 11 2 11 9 0 0 9 2
21 1 11 1 0 9 13 9 11 9 0 9 2 15 13 0 9 9 10 0 9 2
10 1 9 9 4 1 12 9 15 13 2
5 15 2 3 2 3
22 11 0 2 9 9 11 1 11 2 15 13 1 10 9 11 11 1 0 9 1 11 2
25 9 2 3 12 0 9 2 15 13 1 9 11 0 9 7 13 15 1 0 9 1 9 7 9 2
2 9 9
11 9 1 0 9 7 9 0 9 11 11 11
4 13 4 15 11
19 11 11 4 13 1 0 9 1 11 2 3 13 9 9 1 9 11 9 2
16 1 9 13 9 11 11 2 7 3 4 13 1 12 1 9 2
11 3 4 13 0 9 1 0 7 0 9 2
8 15 15 7 13 3 0 9 2
13 11 11 2 1 0 9 9 11 13 1 0 9 2
11 1 11 7 0 9 7 3 13 7 13 2
14 15 13 10 9 0 9 1 9 9 14 1 9 11 2
37 1 0 9 1 9 1 0 0 9 4 1 9 12 13 1 9 1 11 9 10 9 7 3 15 1 9 9 2 16 15 13 3 10 9 2 13 2
16 0 9 13 2 16 13 0 13 9 2 7 11 14 15 13 2
7 13 4 15 2 16 13 2
23 13 4 0 7 3 0 0 9 1 11 1 11 2 3 1 11 2 7 1 11 1 11 2
14 3 4 13 9 1 9 0 0 9 2 3 1 9 2
11 13 4 12 9 7 3 3 1 9 9 2
18 13 4 1 0 0 9 1 11 2 3 4 13 13 14 1 0 9 2
16 1 12 9 4 13 1 9 9 3 0 9 2 3 3 13 2
24 13 9 2 16 3 13 7 3 3 13 2 0 0 9 4 13 1 9 0 9 1 11 2 2
8 0 12 2 9 4 13 9 2
8 1 10 9 4 15 13 13 2
14 3 15 9 13 13 0 2 13 4 13 0 9 9 2
20 1 9 13 1 9 1 10 9 7 13 3 0 2 16 15 13 1 9 3 2
18 15 15 3 13 2 16 7 3 3 0 9 1 0 9 11 13 3 2
23 11 9 15 13 1 15 2 16 15 12 9 1 9 13 9 7 13 15 13 1 10 9 2
17 1 0 12 9 4 13 1 11 11 1 12 9 7 1 10 9 2
19 9 9 9 11 13 1 15 9 7 10 9 13 3 15 1 15 3 0 2
19 0 0 9 15 13 0 9 2 15 13 9 0 0 9 7 0 9 9 2
14 3 3 2 16 13 9 9 2 13 1 15 0 9 2
9 0 9 9 11 4 13 0 9 2
11 13 15 1 9 9 0 9 0 1 9 2
16 10 9 13 2 16 4 13 13 0 2 16 4 13 13 9 2
11 16 10 9 13 2 13 15 1 15 13 2
33 13 7 2 16 4 3 16 9 13 9 2 15 4 15 1 10 9 13 3 13 2 7 7 1 10 9 4 13 3 1 0 9 2
8 13 4 3 1 9 1 11 2
16 13 15 15 7 1 9 2 16 15 4 13 3 13 1 11 2
28 0 4 15 7 13 1 10 9 7 13 0 12 9 1 11 7 9 11 2 3 4 13 1 9 12 0 9 2
20 14 1 9 4 15 13 1 11 13 9 9 1 9 9 11 7 10 0 9 2
7 13 2 16 15 15 13 2
4 11 11 2 11
4 9 9 7 9
14 0 9 9 13 1 0 9 2 0 9 9 13 0 2
17 1 9 4 13 0 9 1 0 11 1 9 7 13 9 1 15 2
27 1 11 13 3 9 2 1 9 7 9 14 13 1 9 2 15 4 1 9 13 1 9 1 9 7 9 2
32 0 0 9 12 7 9 12 9 2 2 1 9 7 9 9 12 7 9 12 9 2 2 0 0 9 12 7 12 9 2 9 2
9 1 9 13 1 9 9 0 9 2
21 1 11 13 3 2 1 9 3 3 7 13 1 9 9 1 9 2 1 9 9 2
25 0 0 9 1 12 2 1 0 9 1 9 12 9 2 2 0 0 9 12 7 12 9 2 9 2
22 1 9 7 1 9 13 1 11 0 9 7 13 7 9 9 2 1 9 9 1 9 2
35 0 9 12 7 12 9 2 9 2 1 9 12 7 12 9 2 9 2 0 9 12 7 12 9 2 9 2 1 9 1 12 9 2 9 2
13 1 9 13 9 1 12 9 7 13 1 12 9 2
11 9 13 1 12 9 7 13 1 12 9 2
37 0 9 9 12 2 9 2 1 9 2 12 1 0 11 2 2 0 9 12 9 2 9 1 9 12 2 0 9 9 12 9 2 9 1 9 12 2
10 0 0 9 13 9 12 9 2 9 2
29 0 9 12 2 9 2 9 2 12 9 2 1 9 12 2 0 2 12 1 9 12 2 9 13 12 9 2 9 2
2 9 2
10 1 0 11 15 13 1 9 0 9 2
2 9 13
29 9 10 0 9 0 9 13 3 1 0 9 9 1 9 9 9 9 11 11 9 11 11 11 0 2 1 9 2 2
7 2 16 13 2 4 13 2
34 16 15 3 13 7 15 3 13 12 9 1 0 9 2 13 4 2 16 15 1 10 9 13 2 2 13 0 2 9 2 3 1 9 2
39 0 1 9 9 9 9 9 12 11 11 15 1 0 9 1 9 13 13 7 1 9 0 9 15 13 2 2 12 2 9 15 15 1 12 9 13 9 11 2
13 0 9 4 13 1 9 2 3 4 13 0 9 2
19 3 15 13 1 9 7 12 2 9 15 13 0 9 1 9 1 11 2 2
33 1 0 9 15 1 9 13 7 0 1 9 11 11 2 15 15 1 0 9 1 0 11 13 9 2 2 3 1 15 15 13 2 2
30 16 11 11 2 0 16 9 9 11 2 13 1 9 2 3 3 13 1 11 2 3 3 2 2 15 13 16 9 2 2
16 9 1 0 13 1 9 12 2 7 16 13 3 2 2 2 2
32 9 9 4 3 13 11 11 1 0 11 2 15 1 0 9 9 12 2 12 13 9 9 1 11 7 3 15 13 1 11 9 2
14 2 0 16 13 0 9 1 11 13 0 9 1 11 2
26 7 4 1 9 13 1 0 9 2 13 12 9 9 7 3 1 10 9 13 0 9 1 0 9 2 2
20 0 9 15 11 13 7 3 2 0 9 1 11 1 9 9 15 13 13 0 2
16 7 16 2 3 1 9 13 2 3 13 1 11 13 2 2 2
3 2 11 2
3 11 13 9
3 0 11 2
21 7 1 9 0 9 7 9 9 9 9 15 13 3 0 11 11 16 0 0 9 2
12 10 9 1 15 14 3 13 10 9 11 11 2
20 15 11 1 15 13 2 2 11 13 3 16 0 1 15 2 16 4 13 0 2
9 10 9 1 15 13 12 2 12 2
5 13 3 0 2 2
13 7 0 0 9 1 11 13 3 3 1 0 9 2
30 12 2 9 1 9 9 1 11 13 1 12 9 12 12 9 0 9 11 11 7 13 3 0 0 0 0 9 1 9 2
16 2 13 3 0 9 2 15 4 15 13 2 2 13 11 11 2
16 2 13 15 15 2 16 15 13 10 9 2 15 13 0 9 2
7 15 15 13 9 9 2 2
9 1 9 15 3 13 7 0 9 2
16 10 9 9 11 13 1 15 2 16 0 0 9 15 3 13 2
30 3 13 11 11 1 12 12 9 7 1 0 9 1 10 9 13 13 2 16 4 15 10 9 13 3 1 0 12 9 2
8 3 13 0 9 3 2 1 11
5 11 1 11 9 2
24 1 0 1 15 13 9 1 9 9 0 11 2 15 13 0 9 2 9 1 0 0 9 9 2
33 1 0 9 15 13 11 2 11 2 11 1 11 11 2 7 1 0 9 13 3 14 12 9 1 3 0 0 9 9 2 1 11 2
6 13 15 11 7 11 2
47 1 0 9 7 1 0 9 11 2 11 2 11 2 11 4 1 0 9 13 3 15 2 16 11 3 13 1 0 11 2 11 7 11 13 1 9 9 7 11 3 9 1 11 11 9 13 2
20 1 9 3 0 0 9 13 3 0 9 11 7 11 2 15 13 1 12 9 2
15 1 0 9 13 3 3 11 2 3 1 11 7 12 11 2
21 1 11 13 12 9 11 7 11 2 11 2 11 2 1 12 11 2 11 7 11 2
65 1 15 13 1 12 0 9 11 2 11 12 5 2 9 2 11 2 2 11 13 12 2 11 12 2 11 2 11 2 11 2 2 3 13 1 0 9 11 2 11 2 11 2 11 2 2 9 2 11 2 11 2 11 2 7 11 2 1 11 12 5 2 11 2 2
40 1 12 9 13 1 12 9 2 11 2 11 2 2 11 2 11 2 2 0 2 11 2 11 2 2 11 2 11 2 2 11 2 11 2 7 11 2 11 2 2
24 0 9 15 13 1 9 12 9 11 11 2 15 1 10 9 13 12 9 7 13 3 0 9 2
22 11 13 3 0 9 2 15 13 10 9 13 3 1 15 2 11 13 12 0 9 2 2
10 3 13 12 0 9 13 9 12 9 2
27 1 9 12 13 1 9 11 11 2 11 2 11 2 12 13 1 11 11 2 7 11 2 11 2 11 2 2
32 1 0 15 13 1 9 12 2 3 1 0 12 9 13 11 11 2 9 11 2 11 7 15 3 13 1 12 9 2 11 11 2
8 9 0 9 10 0 9 13 2
35 3 1 9 3 13 11 11 2 9 11 2 15 13 1 0 9 12 9 2 12 11 2 11 2 11 2 11 2 7 12 11 2 11 2 2
23 11 13 7 3 1 9 9 11 11 7 11 15 13 2 3 3 13 3 13 2 11 11 2
10 0 2 9 13 1 0 9 9 3 2
36 1 9 12 15 13 1 9 1 11 11 11 9 9 7 1 9 12 2 3 4 13 9 0 9 2 13 11 11 1 0 9 2 13 11 2 2
3 2 11 2
7 1 9 15 1 11 13 9
3 16 9 9
43 13 15 9 1 9 7 13 3 0 12 2 9 11 2 15 3 13 1 11 2 13 1 0 9 1 11 2 11 2 12 2 9 1 11 7 13 12 2 12 2 1 11 2
22 14 1 10 9 1 9 15 13 0 9 1 9 1 11 2 15 13 3 1 12 9 2
16 3 1 9 0 15 9 13 9 1 9 12 9 16 9 9 2
20 1 9 11 2 11 7 11 2 15 13 1 0 9 0 9 2 15 9 13 2
28 1 0 9 9 13 13 2 9 2 1 9 0 9 1 0 9 7 1 11 2 15 1 0 9 13 11 11 2
11 15 1 11 13 7 3 13 0 7 0 2
11 1 10 9 9 13 9 1 11 3 9 2
26 7 11 11 2 9 9 7 3 9 9 2 15 13 2 16 1 0 9 9 13 7 14 15 4 13 2
21 11 13 2 16 15 1 0 9 3 13 9 7 9 0 1 0 9 2 1 9 2
31 10 9 3 13 11 11 7 1 15 13 7 11 11 2 15 1 9 0 7 0 9 9 1 9 0 1 9 13 0 9 2
37 1 10 12 9 4 13 1 11 10 9 7 13 3 0 9 9 7 0 9 2 15 3 1 11 1 11 13 2 14 16 13 1 9 9 2 2 2
20 1 0 9 1 9 13 0 9 15 1 9 2 11 2 11 2 11 2 11 2
19 3 7 13 10 0 0 11 11 2 15 9 11 7 13 0 9 2 2 2
15 1 0 9 15 15 3 3 13 2 7 1 11 13 0 2
24 11 11 15 13 9 3 1 9 11 2 15 3 13 1 11 3 0 2 7 3 15 9 13 2
18 1 11 3 3 13 2 16 0 9 4 1 1 9 13 1 9 9 2
27 12 9 15 3 1 9 13 2 7 9 12 1 11 1 0 9 3 13 9 2 16 4 13 9 1 9 2
29 1 15 15 13 2 7 16 15 13 9 0 9 11 11 2 15 15 7 1 0 9 13 1 9 9 3 3 0 2
9 1 10 9 15 7 3 13 9 2
3 2 11 2
9 11 15 13 13 7 1 9 11 2
14 0 9 13 12 9 0 9 1 0 9 1 0 9 2
2 9 11
4 15 13 9 2
2 11 2
14 15 13 12 2 9 0 9 1 9 1 11 0 9 2
21 9 13 2 16 9 9 13 13 14 12 9 1 0 9 2 3 3 15 15 13 2
32 11 2 11 11 13 2 16 0 9 0 9 4 13 13 0 11 11 2 15 9 13 1 12 9 0 9 1 9 2 0 11 2
6 0 9 13 11 11 2
26 13 1 9 11 1 0 11 2 3 15 4 13 15 1 0 9 2 16 4 15 13 1 0 9 9 2
3 11 1 9
37 7 0 9 1 9 0 11 12 2 11 7 0 9 11 13 1 0 9 9 11 11 2 9 11 2 15 13 1 9 1 11 7 13 3 13 2 2
42 0 9 11 11 7 13 2 2 15 13 1 9 9 3 2 1 9 13 11 11 2 11 1 0 11 2 9 13 1 9 1 11 2 1 9 13 7 9 11 2 2 2
11 16 4 13 9 11 2 13 15 16 9 2
19 1 11 13 3 0 9 2 1 15 13 9 0 2 7 3 15 13 13 2
12 13 15 1 9 7 1 11 13 0 9 2 2
3 2 11 2
6 9 11 2 0 2 9
3 12 0 2
23 0 9 9 11 2 0 9 1 11 1 11 2 12 9 2 1 11 15 13 12 0 9 2
21 12 9 0 9 11 2 11 2 11 4 13 1 9 0 9 1 9 9 1 11 2
45 1 12 9 13 1 9 9 9 11 2 11 2 2 11 2 1 9 12 2 12 9 2 1 11 2 11 2 2 11 2 7 12 2 12 9 2 1 11 2 11 2 2 11 2 2
7 9 13 11 11 1 11 2
21 1 9 13 11 1 11 2 11 2 13 7 9 2 2 1 9 0 9 3 13 2
2 9 13
2 11 2
14 9 9 1 9 9 11 11 15 13 9 9 1 11 2
17 12 9 0 7 12 0 9 10 9 13 7 1 9 12 7 12 2
16 1 0 9 13 9 9 1 9 11 7 0 9 1 9 11 2
20 1 9 13 1 0 9 9 9 1 0 9 11 1 9 11 7 0 9 11 2
8 9 9 15 13 0 9 9 2
2 11 13
2 11 2
34 1 12 9 1 11 1 9 11 0 11 15 13 11 11 1 0 11 2 13 1 11 11 2 7 13 15 9 9 0 15 9 0 9 2
36 9 9 1 9 9 15 7 13 9 0 0 9 2 10 9 11 2 11 13 2 2 12 1 0 9 11 13 3 2 0 2 9 1 10 9 2
10 3 3 14 13 9 13 2 2 2 2
17 9 7 11 3 13 7 13 0 9 14 1 0 9 0 0 9 2
3 11 1 11
2 11 2
26 0 9 12 2 0 9 11 11 13 1 9 9 2 12 0 11 11 11 1 0 9 11 0 2 11 2
22 2 1 9 1 11 13 13 1 11 9 0 9 2 2 13 9 0 11 11 2 11 2
23 2 13 13 2 16 13 0 9 7 1 9 12 2 12 15 13 12 9 7 12 9 2 2
2 0 9
2 11 2
27 0 0 2 0 9 9 7 9 2 1 15 3 3 1 9 13 0 9 2 13 3 1 0 9 0 9 2
41 1 0 9 9 0 2 7 0 9 4 15 13 9 0 2 9 1 12 9 13 1 12 2 1 12 9 1 11 1 0 9 4 7 13 13 1 12 9 1 11 2
11 9 9 7 9 4 3 13 1 12 9 2
4 9 7 9 11
2 11 2
18 9 11 11 11 2 11 13 1 9 1 0 11 10 0 9 1 11 2
39 3 9 1 9 0 12 13 9 11 12 2 12 2 1 12 12 9 3 13 9 1 12 2 12 7 12 9 1 0 9 9 9 13 1 9 12 2 12 2
29 11 13 9 1 12 9 1 9 2 2 3 4 13 1 9 2 3 4 9 13 1 12 9 7 3 3 13 2 2
26 2 11 11 1 0 9 13 12 9 7 0 9 12 9 15 13 1 12 2 9 9 0 9 11 2 2
2 0 0
2 11 2
38 1 9 1 0 9 13 9 9 11 2 0 9 0 9 1 0 9 2 15 13 1 11 1 11 7 13 12 9 2 1 15 12 9 13 0 0 9 2
5 9 9 9 13 2
9 0 2 7 7 0 9 9 9 11
2 0 9
5 11 2 11 2 2
18 12 9 1 9 13 0 9 10 0 0 0 9 2 12 2 11 11 2
34 1 12 9 15 9 13 1 12 9 2 0 12 9 4 13 3 0 1 0 0 9 2 16 9 13 1 9 7 9 0 1 0 9 2
24 9 2 15 13 0 9 2 15 13 9 11 7 13 1 9 1 9 1 12 2 0 0 9 2
29 9 2 15 13 1 12 2 2 12 2 9 2 13 3 0 1 0 1 9 1 9 2 1 15 13 0 12 9 2
16 1 9 1 0 9 13 9 1 9 7 9 0 1 0 9 2
13 7 1 10 9 4 13 0 9 1 0 9 9 2
25 9 0 9 13 0 9 2 15 15 13 1 9 9 1 0 9 7 1 0 9 15 3 15 13 2
13 3 10 9 3 13 1 0 11 1 0 12 9 2
26 1 0 9 2 3 13 11 2 13 11 12 9 2 3 1 12 3 16 11 2 1 0 9 12 9 2
34 15 0 1 12 2 9 1 9 11 1 9 9 13 7 0 2 7 1 9 13 3 3 9 1 9 2 3 13 3 13 2 3 0 2
14 11 11 3 16 11 13 3 1 9 9 3 10 9 2
15 9 13 0 9 11 2 15 3 13 3 1 9 1 9 2
26 0 11 11 13 0 9 1 9 2 0 12 9 13 7 13 15 15 0 9 1 9 9 1 9 9 2
23 3 7 10 9 13 1 9 2 13 13 3 9 7 13 16 0 1 0 9 1 0 9 2
20 0 13 11 2 15 9 13 9 9 2 3 12 2 15 13 3 1 15 9 2
21 0 9 13 1 0 9 9 1 0 9 2 3 16 9 13 3 1 9 0 9 2
23 0 9 0 9 1 9 0 13 3 0 9 2 9 2 15 1 0 0 9 13 0 9 2
38 1 9 1 0 9 3 13 0 9 1 11 2 7 9 9 1 0 9 13 10 9 13 3 1 9 1 9 2 1 15 7 13 1 0 9 0 9 2
36 9 9 11 2 0 11 2 11 7 11 13 1 9 1 9 3 0 9 2 16 9 11 0 15 1 0 9 1 0 12 9 13 3 1 9 2
30 1 0 9 12 9 2 9 11 2 11 13 0 2 13 0 12 7 2 12 7 15 13 9 3 7 12 7 13 9 2
18 3 13 12 9 1 9 12 2 12 2 15 13 9 12 9 1 9 2
19 4 13 12 0 9 2 12 0 2 12 0 7 12 9 13 3 1 9 2
12 9 13 12 9 2 15 13 9 12 1 9 2
12 9 9 13 1 12 9 0 9 7 0 11 2
1 9
4 15 4 13 2
31 1 12 2 9 9 13 1 0 9 12 9 1 12 9 2 1 0 12 9 1 12 9 2 1 0 12 9 1 12 9 2
51 1 12 2 9 11 13 1 12 2 9 1 0 9 12 9 12 9 2 1 0 13 12 9 1 12 9 2 1 0 12 9 1 12 9 2 1 0 12 9 1 12 9 2 1 0 12 9 1 12 9 2
46 1 12 2 9 13 1 0 9 12 9 12 9 2 1 0 13 12 9 12 9 2 1 0 13 12 9 1 12 9 2 1 0 12 9 1 12 9 2 1 0 12 9 1 12 9 2
43 1 12 2 9 0 9 12 1 12 13 1 0 9 12 9 12 9 2 1 0 13 12 9 1 12 9 2 1 0 12 9 1 12 9 2 1 0 12 9 1 12 9 2
1 9
29 1 0 9 1 11 2 12 9 2 13 11 0 12 2 12 7 11 0 12 2 12 2 13 11 11 12 2 12 2
1 9
32 1 0 9 1 0 11 13 11 11 1 0 11 0 2 11 12 2 12 7 13 11 11 12 2 12 7 11 0 12 2 12 2
3 9 2 9
23 0 9 9 12 13 1 0 9 1 9 11 11 2 9 12 9 2 0 9 11 9 12 2
22 9 15 13 13 1 9 1 9 2 9 2 0 2 9 2 9 12 2 12 12 11 2
1 3
2 0 9
22 1 0 9 11 13 11 2 11 9 11 12 2 12 7 11 9 11 11 12 2 12 2
2 1 9
6 1 1 0 2 2 2
18 1 9 11 13 11 0 12 2 12 7 1 9 15 13 1 11 11 2
17 11 11 2 0 0 9 7 9 9 11 2 15 13 9 11 11 2
6 9 13 9 1 0 9
5 13 15 11 11 2
2 11 2
24 0 9 13 2 16 1 9 1 9 1 9 0 1 0 9 3 13 0 9 0 9 11 11 2
15 11 13 9 9 11 1 11 7 13 13 12 2 9 12 2
25 9 12 2 9 12 13 2 16 15 13 9 1 0 0 9 1 9 9 9 1 9 11 1 11 2
26 0 9 0 0 9 2 9 2 3 1 0 9 1 9 11 1 11 13 2 16 0 9 13 11 11 2
35 1 0 9 9 13 2 16 2 13 9 2 16 15 13 11 11 1 11 2 2 7 3 13 9 1 11 2 15 13 13 14 12 0 9 2
16 0 0 9 9 11 13 2 16 9 13 13 0 1 0 9 2
8 13 3 1 9 7 9 9 2
29 9 9 1 0 9 1 11 2 3 13 9 13 2 13 2 16 13 1 12 9 0 2 16 13 1 11 2 11 2
21 10 9 4 13 9 0 0 9 11 11 2 15 4 13 1 9 12 1 0 11 2
23 3 13 13 11 7 11 2 1 15 15 13 2 16 13 13 1 12 9 2 0 1 9 2
32 1 9 0 9 9 13 13 12 11 2 1 15 10 9 13 9 9 11 2 15 13 13 1 11 1 9 2 0 9 7 9 2
22 3 1 9 7 9 11 11 7 11 11 13 2 16 15 13 2 16 11 13 12 9 2
34 1 9 2 15 13 0 0 9 2 0 9 1 9 2 2 11 13 0 9 2 1 15 13 0 9 11 11 2 16 4 13 9 0 2
4 9 15 13 13
38 1 11 1 12 2 12 2 13 9 1 9 11 11 0 1 9 2 1 15 15 9 0 3 1 9 11 2 11 7 11 13 1 9 9 11 2 11 2
21 9 13 9 9 10 9 2 1 15 9 0 13 2 16 4 13 4 1 9 13 2
40 12 1 9 2 15 9 11 13 9 0 2 13 3 2 2 13 3 9 2 16 4 13 10 9 1 9 12 2 9 2 15 13 7 9 9 7 9 9 2 2
12 9 11 0 2 2 15 15 3 13 10 9 2
22 16 15 15 13 2 16 4 15 13 2 7 13 2 14 6 13 9 2 15 3 13 2
11 13 2 14 15 3 2 13 15 3 13 2
8 7 1 9 15 13 13 2 2
42 10 9 9 0 9 1 9 9 2 16 15 13 9 1 9 10 9 2 13 3 0 2 16 15 7 13 9 2 16 4 15 13 1 15 2 1 15 1 9 3 13 2
10 4 13 9 1 9 1 9 12 9 2
27 11 0 16 12 1 15 15 13 15 13 7 1 15 13 15 2 15 13 2 16 4 2 3 2 13 9 2
23 14 9 0 13 2 16 10 9 13 3 14 7 14 0 9 9 2 16 1 15 13 9 2
7 7 16 15 13 0 9 2
16 11 0 13 13 2 16 1 15 15 13 2 3 2 13 9 2
11 9 1 0 9 9 13 1 9 16 9 2
32 9 9 3 13 1 15 2 16 4 1 9 13 13 2 7 9 2 15 13 1 9 9 2 3 13 2 16 1 15 9 13 2
16 1 15 15 11 0 13 13 0 15 2 16 4 13 0 9 2
22 1 15 3 15 13 13 1 15 2 16 4 13 9 2 16 10 0 9 13 0 9 2
8 3 15 4 13 3 2 2 2
42 9 2 1 0 0 9 9 12 13 2 16 3 3 2 7 16 13 2 12 4 3 7 13 2 9 9 13 1 15 2 16 4 12 9 0 0 9 1 0 9 13 2
34 16 3 1 0 9 13 1 0 0 9 2 15 13 2 13 1 0 9 13 1 15 15 0 2 16 1 9 3 15 13 14 0 9 2
8 13 15 3 7 13 15 3 2
15 3 12 3 13 9 7 1 9 2 0 3 1 0 9 2
4 9 2 11 11
4 11 11 1 11
10 9 9 2 7 15 13 2 3 2 3
18 3 15 13 9 2 15 4 3 3 7 3 13 1 15 2 16 11 2
29 16 3 2 3 1 3 2 7 3 3 2 0 9 3 13 10 9 1 9 2 2 0 9 2 15 13 11 2 2
37 1 9 13 3 13 9 7 9 2 13 15 1 9 0 9 7 9 2 16 4 15 1 15 9 7 9 13 1 0 9 1 15 2 15 3 13 2
21 16 3 2 3 15 3 13 2 16 13 15 1 3 0 9 0 7 3 0 2 2
10 9 11 11 1 0 9 13 1 9 12
6 0 9 1 9 1 9
2 0 9
28 9 13 0 9 12 2 12 2 12 1 0 9 2 3 16 9 9 2 15 11 11 13 1 0 7 0 9 2
36 9 9 1 2 0 2 9 1 9 13 14 0 9 0 9 9 1 10 9 2 7 7 9 1 9 2 15 9 9 1 9 11 11 3 13 2
37 9 13 9 1 0 9 2 9 2 11 13 1 0 9 2 15 13 1 2 0 2 9 2 9 2 9 3 2 2 7 15 15 13 0 9 13 2
27 3 15 13 1 9 0 9 2 11 2 15 1 15 13 2 16 13 9 0 9 2 7 1 9 2 2 2
31 11 15 13 0 9 9 1 9 0 9 2 15 13 1 0 9 2 16 15 3 13 2 7 3 15 13 10 9 7 9 2
33 3 7 13 1 9 2 15 13 1 10 9 1 0 9 2 9 11 2 7 9 2 7 11 11 2 2 9 3 13 9 9 2 2
34 11 2 11 11 2 13 15 15 2 9 13 15 1 9 2 3 15 13 0 9 1 9 2 0 9 9 0 9 7 9 1 9 11 2
33 1 0 2 0 9 15 13 1 0 9 2 7 2 1 1 11 11 2 9 0 0 9 2 9 12 2 2 15 11 13 9 9 2
21 1 10 0 9 13 1 9 2 7 15 15 13 2 13 9 2 13 9 9 11 2
30 13 15 2 16 13 1 9 2 15 13 1 15 2 7 1 9 13 9 1 15 15 2 16 15 13 1 2 9 2 2
16 11 9 13 1 9 11 3 3 0 2 13 1 9 7 9 2
12 3 13 9 9 1 9 0 2 13 0 9 2
69 3 13 9 1 9 2 3 13 0 9 7 1 9 2 3 11 13 1 9 9 7 13 10 9 1 15 2 3 3 15 4 13 1 9 9 2 15 11 13 1 9 7 1 9 15 13 9 9 1 10 9 2 14 2 3 9 13 11 1 10 9 2 16 15 13 10 0 9 2
60 9 11 11 15 13 1 9 9 2 7 1 1 10 9 2 11 11 2 2 15 13 1 3 16 1 0 9 0 9 2 13 1 15 1 15 0 7 0 9 0 1 0 7 0 9 9 0 9 2 15 13 15 3 0 2 16 13 0 9 2
36 11 2 11 11 2 13 0 9 9 0 15 1 9 9 2 9 7 0 0 9 1 9 2 9 2 15 15 13 3 1 9 9 10 0 9 2
43 11 2 11 11 2 13 2 3 16 11 1 9 7 11 1 9 2 0 0 9 2 15 15 13 1 10 0 9 1 9 2 15 13 1 0 9 2 7 3 4 15 13 2
15 11 11 13 9 2 1 15 13 0 2 9 2 10 9 2
19 2 3 2 16 10 2 9 2 13 9 0 9 2 15 1 9 13 2 2
83 0 9 3 0 1 0 9 2 3 2 0 2 11 11 2 9 1 9 2 9 14 0 9 11 11 1 9 11 1 0 9 2 2 9 2 11 11 2 3 0 0 2 0 7 0 9 2 9 2 11 11 2 2 10 0 9 7 9 2 1 0 9 2 13 0 15 9 2 9 7 9 2 0 15 9 9 2 15 13 9 0 9 2
43 3 16 15 1 9 11 13 1 10 9 0 9 2 7 14 1 9 0 9 2 2 13 11 9 0 9 1 9 1 9 2 13 3 0 9 0 9 1 9 2 12 2 2
30 1 0 9 1 9 11 7 9 9 4 9 2 7 1 1 9 2 15 9 9 1 11 13 2 13 1 9 14 0 2
40 3 0 0 9 2 1 9 11 7 9 15 1 9 13 3 11 11 7 11 11 2 13 3 3 2 15 13 0 2 13 15 9 0 2 0 9 2 10 9 2
4 7 9 0 2
15 15 13 13 9 2 15 13 0 9 7 13 1 0 9 2
17 9 15 13 2 9 15 3 3 13 2 7 7 4 13 2 2 2
19 1 0 9 13 12 0 9 2 15 13 9 1 9 0 9 9 1 9 2
3 11 7 2
1 0
3 11 11 2
3 9 1 11
2 11 2
29 0 9 11 11 13 3 1 12 0 9 1 11 7 11 2 15 13 1 10 9 1 9 0 9 1 0 9 11 2
14 2 0 9 1 10 9 13 0 9 2 2 13 9 2
15 12 1 9 2 3 13 0 9 11 2 13 13 0 9 2
37 2 0 0 9 9 9 13 0 12 0 9 2 2 13 11 2 15 1 10 9 13 12 0 9 0 0 9 2 15 4 13 9 13 1 0 9 2
41 9 13 2 16 4 13 9 0 9 1 0 9 2 16 2 0 9 13 0 9 2 7 0 9 13 13 1 9 9 3 0 9 2 16 13 0 9 1 9 11 2
27 0 0 9 13 3 11 2 7 0 9 4 13 1 9 11 7 0 11 2 1 15 13 11 0 0 9 2
7 11 2 0 9 2 0 9
3 3 0 9
7 0 0 9 2 0 9 2
9 1 0 9 0 9 7 0 9 2
9 15 13 9 10 9 1 10 9 2
10 11 2 7 7 0 9 13 9 9 2
9 3 0 9 13 1 11 7 11 2
15 9 1 9 3 1 11 13 3 1 9 2 13 0 9 2
13 1 0 9 13 12 9 9 2 1 0 9 12 2
14 9 1 9 7 11 13 1 9 2 3 3 15 9 2
10 9 1 11 1 11 13 1 9 0 2
8 9 13 1 9 2 1 9 2
21 2 13 10 9 2 1 9 3 13 0 9 2 2 13 15 9 0 9 11 11 2
6 2 13 1 15 9 2
17 0 9 13 1 9 9 2 1 9 4 13 0 9 1 12 9 2
5 15 13 7 3 2
12 1 9 2 15 4 3 13 2 4 9 13 2
15 1 9 15 13 3 0 9 7 12 9 1 15 13 11 2
14 13 15 1 9 1 11 2 15 13 7 9 0 9 2
18 13 2 16 9 13 3 0 7 3 15 3 13 2 2 13 9 9 2
14 1 3 0 0 9 4 15 13 13 7 1 0 9 2
17 3 2 9 11 1 0 9 2 2 13 3 3 1 12 2 9 2
9 10 9 13 9 9 1 15 2 2
16 9 1 0 2 12 9 2 1 9 1 12 9 2 12 9 2
10 3 1 9 11 13 9 3 15 9 2
19 0 9 1 0 9 11 3 1 9 13 2 7 9 13 3 0 1 9 2
17 7 1 9 9 9 2 12 9 0 1 0 2 12 9 1 9 2
26 3 0 13 7 0 9 2 7 15 2 15 2 16 13 0 9 2 13 9 9 2 16 3 0 11 2
27 7 3 0 0 9 9 1 0 9 13 2 3 0 9 1 11 4 13 14 1 9 2 9 9 1 9 2
3 7 9 2
24 1 2 9 2 16 13 9 2 12 0 9 1 9 2 3 12 9 2 3 1 9 1 9 2
16 1 0 9 13 12 2 12 9 9 2 9 0 9 13 0 2
10 10 9 13 0 7 0 9 13 13 2
9 3 13 4 9 1 11 7 11 2
21 0 9 13 3 1 11 0 2 1 12 9 1 0 14 1 12 9 1 0 9 2
15 16 15 1 9 13 0 9 2 13 9 9 0 1 9 2
16 0 9 13 13 7 13 1 15 0 12 9 9 9 1 9 2
13 9 1 9 13 2 7 9 7 9 13 3 13 2
13 3 9 11 1 11 13 12 9 13 14 1 9 2
14 1 11 1 9 13 12 9 2 0 9 7 0 9 2
15 3 3 13 0 9 13 2 7 0 9 13 3 16 3 2
15 9 11 13 15 12 9 13 14 1 9 3 1 0 9 2
9 3 1 11 13 0 9 3 0 2
9 1 9 13 1 9 9 0 9 2
28 9 0 9 1 9 11 7 0 15 13 1 12 1 12 9 2 0 1 12 9 7 0 9 13 1 12 9 2
3 2 11 2
4 9 1 0 9
29 9 0 9 15 3 1 9 1 12 9 13 9 2 16 4 15 1 9 13 1 9 7 13 15 2 16 13 9 2
9 1 10 9 15 13 9 0 9 2
34 13 0 9 9 11 2 15 2 3 13 1 0 9 1 11 2 2 13 0 9 9 0 2 9 13 0 2 2 3 7 0 9 11 2
11 13 9 11 2 3 15 13 1 9 11 2
26 13 1 9 9 11 2 15 13 2 15 1 12 3 3 0 9 13 16 0 2 9 0 7 9 0 2
18 1 0 9 9 2 14 1 9 0 0 9 2 13 9 0 15 9 2
43 7 16 15 0 9 13 1 0 9 2 13 3 15 2 15 3 1 0 9 1 0 2 0 2 0 7 0 9 7 9 13 2 0 1 9 0 9 7 0 9 2 2 2
8 0 0 9 4 13 0 9 2
20 1 0 0 9 9 12 13 1 3 0 0 9 9 7 0 9 11 11 11 2
6 13 1 9 7 9 2
16 7 13 3 3 2 16 15 9 7 9 1 9 13 1 9 2
8 13 15 2 15 15 13 13 2
26 9 13 3 10 9 2 3 3 2 16 2 0 9 2 15 1 11 13 3 0 9 9 1 0 9 2
13 9 1 0 9 13 11 1 11 7 13 15 9 2
8 1 0 9 3 13 9 9 2
30 9 11 2 3 3 9 2 2 3 16 0 1 15 2 1 15 15 0 9 13 2 13 1 9 12 1 9 2 2 2
28 3 11 1 11 2 9 7 9 2 13 2 16 1 9 9 13 12 0 9 2 9 7 9 7 9 7 9 2
5 11 13 15 0 2
15 13 7 13 2 16 9 10 9 1 9 13 13 0 9 2
19 3 4 15 13 1 0 9 2 15 0 9 1 0 9 13 9 3 13 2
20 13 4 10 9 3 0 9 1 9 0 9 7 13 4 15 15 0 9 13 2
30 1 9 1 9 0 9 7 0 9 2 3 0 9 12 13 9 2 13 9 1 0 9 3 14 0 9 2 2 2 2
32 7 2 15 13 3 13 9 1 10 9 2 0 9 2 1 15 15 1 0 9 7 3 13 13 10 0 9 2 7 0 9 2
2 11 11
3 9 1 11
3 11 13 0
2 11 2
15 1 9 9 1 0 11 13 0 9 0 9 7 0 9 2
17 7 13 0 1 11 1 9 9 9 3 13 7 13 9 0 9 2
40 13 15 0 0 9 11 11 1 0 9 0 9 1 0 9 2 15 13 1 9 9 7 9 1 9 1 9 9 9 7 3 0 0 9 0 16 2 9 2 2
12 9 9 1 0 9 13 9 9 1 0 9 2
17 11 3 13 2 16 2 2 0 9 1 11 13 0 1 9 2 2
2 11 2
1 11
3 9 1 9
2 11 2
33 3 1 0 0 9 1 9 13 10 0 9 0 11 7 0 9 11 13 0 9 1 0 9 2 1 9 2 9 7 3 0 9 2
8 13 15 0 9 11 0 11 2
19 1 9 9 13 7 0 0 9 2 0 13 9 1 9 12 7 12 9 2
25 15 13 15 2 16 0 9 0 9 2 0 14 1 9 1 0 11 2 13 13 0 9 11 11 2
32 9 13 1 12 9 2 3 4 1 0 11 13 9 9 7 13 10 9 2 12 11 2 12 11 2 12 11 7 12 9 11 2
20 0 9 15 13 2 16 0 9 1 0 9 15 13 1 0 9 0 0 9 2
26 1 9 0 11 13 3 3 12 0 0 9 2 7 1 9 1 9 0 3 14 15 13 1 0 9 2
14 9 1 0 9 1 0 9 15 13 1 12 9 9 2
2 0 9
3 0 11 2
58 0 9 11 11 11 1 11 1 9 1 0 9 11 11 2 15 13 1 0 11 2 16 4 15 13 0 9 1 9 12 9 0 0 9 1 10 9 2 13 9 2 16 9 1 0 9 4 13 3 1 15 2 16 13 1 10 9 2
32 2 13 4 15 1 9 7 9 9 0 9 11 11 7 13 4 15 1 3 0 9 1 9 1 9 2 2 13 11 1 11 2
30 2 15 9 15 13 3 3 3 2 7 3 13 13 10 9 2 2 13 0 9 11 2 15 13 0 9 1 0 9 2
33 3 16 1 9 0 9 1 11 13 11 2 11 1 11 13 13 7 1 9 1 11 1 9 7 1 0 9 15 9 1 9 11 2
4 9 1 0 9
11 1 9 0 9 1 11 4 13 9 0 9
2 9 12
4 9 1 9 9
14 15 15 4 13 2 3 2 7 15 2 1 9 2 2
2 9 12
3 11 11 2
7 9 9 2 7 15 13 3
2 9 12
5 0 9 1 0 9
2 0 11
20 1 9 13 9 11 13 10 9 1 9 0 7 0 9 2 1 15 3 13 2
20 15 3 13 2 16 3 9 2 0 9 7 0 9 1 9 3 13 9 9 2
32 1 9 12 4 1 0 9 2 13 2 10 9 2 7 9 11 4 3 3 13 1 9 2 16 9 0 9 13 13 9 0 2
34 9 0 9 7 9 4 13 10 9 0 9 2 15 15 13 1 3 0 9 0 9 1 0 9 1 0 9 7 1 0 9 0 9 2
10 7 0 9 1 11 13 1 10 9 2
15 1 9 0 9 0 9 13 13 1 12 9 9 0 9 2
27 9 1 9 7 0 9 0 9 1 0 9 13 0 2 0 2 0 7 0 0 9 1 9 9 10 9 2
10 2 0 11 2 2 9 12 0 9 2
27 15 15 3 13 2 3 0 9 7 0 9 13 1 12 2 0 9 7 9 7 13 15 9 0 0 9 2
43 0 9 13 12 1 0 0 9 0 9 2 10 9 13 0 9 9 9 0 9 7 9 9 2 9 7 9 15 4 13 1 0 9 10 0 9 2 15 13 0 0 9 2
24 13 15 1 0 9 1 9 2 1 9 7 9 2 15 7 12 1 0 9 9 13 0 13 2
29 11 11 2 0 9 1 0 9 13 2 16 0 0 9 3 13 7 1 0 9 2 3 1 11 2 11 7 11 2
26 0 0 9 2 9 9 7 0 9 13 9 0 9 3 7 13 1 0 9 0 9 9 1 0 9 2
17 11 3 3 13 2 16 0 9 13 2 7 3 3 10 9 13 2
21 0 0 9 15 3 13 3 1 9 0 0 9 7 1 0 9 0 9 7 9 2
32 1 9 1 0 9 2 0 11 2 13 9 0 0 9 11 11 2 16 2 13 13 2 16 0 9 13 0 9 1 9 11 2
21 13 9 2 16 1 11 13 9 2 1 15 4 13 2 7 10 9 15 13 13 2
45 0 9 13 9 0 9 2 9 0 9 13 0 7 0 9 0 9 7 11 2 11 7 9 15 13 13 1 0 9 9 11 2 15 13 3 0 0 9 2 15 13 10 9 2 2
22 0 7 0 0 9 13 2 16 1 12 7 12 9 15 3 13 0 9 1 0 9 2
31 11 2 11 2 11 2 11 2 0 11 2 7 1 10 0 9 13 3 0 13 7 11 2 3 13 1 9 0 0 9 2
17 10 9 11 13 13 1 0 9 15 9 3 0 2 3 0 9 2
10 11 13 1 9 1 0 9 0 9 2
15 15 9 13 4 13 1 9 2 7 3 3 1 0 9 2
18 9 0 9 7 9 1 15 13 1 3 0 9 3 0 2 3 0 2
20 9 10 0 9 13 9 7 16 15 13 3 2 13 0 13 2 3 13 0 2
25 0 9 4 3 13 13 0 9 1 9 2 15 3 13 1 15 3 0 2 0 9 1 0 9 2
26 2 3 3 13 11 13 9 1 9 9 7 1 0 9 0 9 2 2 13 9 9 0 11 11 11 2
25 2 16 4 1 9 0 9 13 0 9 2 13 10 9 1 9 3 0 2 14 2 14 0 2 2
4 11 11 2 11
24 9 0 0 0 9 11 11 3 13 12 1 0 9 1 9 1 9 9 11 11 7 0 9 2
4 9 11 2 11
4 11 2 11 2
3 9 15 13
2 11 2
31 0 2 0 9 2 1 10 9 13 9 0 9 2 3 15 0 9 1 0 9 13 2 2 13 9 0 0 9 11 11 2
27 1 0 9 0 0 11 0 9 9 13 2 16 0 9 2 3 15 13 2 7 9 1 0 9 13 2 2
35 0 9 0 11 2 9 1 9 7 1 9 2 4 13 1 9 7 13 3 0 2 13 11 1 9 2 15 13 0 0 9 9 0 11 2
18 9 1 10 9 13 3 10 0 9 2 7 16 9 13 0 11 13 2
2 9 11
2 0 9
2 11 2
20 9 1 9 1 0 11 13 11 0 0 9 1 9 2 16 4 13 1 9 2
6 13 15 0 9 11 2
12 9 13 7 0 9 2 15 13 13 1 0 2
30 3 13 1 9 1 9 15 2 9 11 2 12 2 9 9 9 2 9 7 0 9 2 15 1 0 9 16 1 9 2
11 9 9 1 0 9 13 13 9 0 9 2
2 0 9
2 0 9
2 11 2
24 2 9 9 2 15 1 9 0 9 13 9 0 9 11 11 2 16 1 0 9 13 12 9 2
8 14 1 9 3 13 11 11 2
11 0 13 11 11 2 0 9 13 11 11 2
15 0 13 9 11 11 2 9 0 9 1 9 1 0 9 2
4 0 9 1 9
17 1 9 1 9 1 11 1 11 13 12 0 9 0 9 1 9 2
11 1 12 9 15 13 1 9 3 1 9 2
19 9 7 9 9 13 2 13 9 7 1 9 12 9 13 0 12 0 9 2
9 9 9 13 9 7 13 0 9 2
19 1 9 9 9 4 12 2 9 1 12 2 9 13 12 9 7 12 9 2
11 13 1 9 12 0 9 2 15 13 9 2
20 0 9 13 2 16 9 15 13 0 9 1 15 1 0 9 11 1 0 9 2
20 13 3 3 2 16 12 9 1 9 12 7 12 9 13 12 0 9 1 9 2
29 9 1 0 9 11 9 13 1 0 9 2 15 12 2 9 3 13 1 9 1 9 1 9 11 12 9 12 9 2
17 9 13 1 9 14 1 0 9 2 3 13 12 9 1 0 9 2
17 3 13 1 0 9 9 9 7 11 7 13 9 1 9 12 9 2
2 9 9
2 11 2
24 2 9 10 9 15 1 0 9 12 13 2 2 13 9 0 2 9 2 9 11 11 2 11 2
27 2 13 15 2 16 12 9 0 9 3 13 7 4 13 1 0 9 1 12 7 1 9 1 12 9 2 2
15 9 2 15 13 9 0 9 2 7 13 0 9 0 9 2
28 1 0 0 9 13 9 10 9 0 12 7 12 9 2 16 1 0 11 15 13 9 9 1 12 7 12 9 2
28 9 11 0 13 9 16 0 9 9 2 0 9 2 1 15 15 13 0 0 9 1 0 9 12 2 9 12 2
38 1 9 2 10 9 13 1 9 12 2 13 7 0 9 1 0 9 2 13 15 3 1 9 0 9 2 0 9 2 9 0 9 7 10 0 0 9 2
3 2 11 2
5 9 11 11 2 11
4 15 13 15 2
20 1 15 3 3 13 0 0 0 9 0 1 12 9 9 11 2 11 7 11 2
45 13 3 9 0 9 2 14 3 1 9 2 11 11 2 11 0 2 11 0 2 11 11 2 11 9 0 2 2 1 9 9 2 11 11 2 11 11 2 11 11 2 11 9 0 2
18 9 15 1 0 9 13 15 0 2 7 7 10 9 7 9 13 0 2
35 13 15 1 15 13 0 2 3 15 15 15 13 2 1 0 9 13 9 9 7 9 2 7 15 15 13 1 15 2 16 13 0 9 2 2
10 3 0 13 9 0 9 7 9 9 2
29 10 9 3 13 2 3 15 0 9 13 2 3 15 13 11 2 13 15 2 7 15 2 2 7 0 15 3 13 2
22 13 7 13 0 2 13 7 15 2 15 15 13 1 11 7 13 7 9 1 15 0 2
15 0 13 2 16 13 9 2 15 13 1 9 13 1 9 2
12 0 9 13 1 9 3 0 0 7 0 9 2
2 11 11
9 9 0 9 1 11 13 3 13 2
24 0 9 9 12 7 0 9 9 0 1 15 13 14 10 9 2 7 3 9 1 11 7 11 2
12 1 9 11 13 1 9 13 9 9 0 9 2
24 9 1 9 13 1 0 9 7 10 2 3 3 0 2 9 9 13 12 2 7 12 2 9 2
16 0 9 11 1 11 13 1 0 9 0 9 1 9 2 0 2
7 0 0 9 13 0 9 2
19 0 0 9 12 9 3 4 13 2 1 9 9 1 11 2 11 7 11 2
25 0 9 9 11 11 0 1 9 10 9 11 15 13 12 2 9 12 1 0 9 0 9 1 11 2
39 9 1 9 2 1 15 13 9 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 7 11 2 11 4 13 1 9 3 0 9 2
29 9 1 0 9 1 9 0 9 4 3 3 13 9 0 7 9 0 11 2 11 1 9 0 2 11 1 0 9 2
16 1 9 9 9 0 9 11 4 13 3 9 1 0 9 3 2
24 0 9 0 2 9 7 0 0 7 0 9 0 2 0 2 11 2 4 3 13 1 9 11 2
9 3 4 3 13 0 9 0 9 2
31 0 2 9 15 1 10 9 13 9 9 7 9 0 9 2 1 9 0 2 0 2 0 2 13 9 9 13 1 0 9 2
25 12 12 9 4 13 1 0 0 9 2 0 0 0 9 2 11 2 1 10 0 9 1 0 9 2
19 10 9 13 9 9 0 9 1 3 0 9 11 12 7 9 11 0 9 2
3 0 9 12
3 9 9 0
21 0 9 13 0 9 1 0 0 9 2 1 15 9 15 1 0 9 13 9 9 2
14 1 9 0 10 9 13 13 2 16 13 1 0 9 2
21 2 3 13 3 0 9 11 2 2 13 3 1 0 9 0 9 14 1 11 12 2
34 12 9 13 0 9 1 0 7 0 9 0 2 16 4 15 3 13 9 7 0 9 2 15 3 1 0 9 0 13 1 9 0 9 2
25 9 14 1 12 9 4 13 0 9 7 0 9 2 3 13 9 1 9 2 16 15 13 9 2 2
17 3 15 0 9 13 7 13 1 9 2 13 9 1 9 7 9 2
32 1 0 9 13 0 9 2 9 15 13 1 9 7 1 0 9 15 13 0 9 0 0 9 2 16 4 2 13 1 9 2 2
29 1 0 9 13 1 15 13 9 2 3 9 2 2 7 7 10 9 2 15 15 13 1 9 0 9 3 13 9 2
18 9 1 9 7 0 9 0 13 3 3 1 9 9 2 9 7 9 2
34 0 9 13 1 9 12 10 9 9 2 1 15 7 14 10 9 9 15 13 3 0 9 2 0 9 2 9 1 9 2 9 7 9 2
26 15 0 9 13 14 0 9 2 13 3 12 9 2 15 13 9 1 0 0 9 1 9 1 0 9 2
28 16 4 13 1 9 0 9 9 2 11 2 11 2 13 4 15 13 1 12 2 3 15 1 15 13 1 11 2
2 11 11
2 9 9
1 9
2 11 2
18 9 0 9 1 9 13 10 9 7 9 9 0 9 7 9 9 0 2
40 9 13 1 15 2 16 4 9 13 13 3 2 9 0 9 2 0 7 0 9 2 9 2 9 0 7 0 2 0 7 0 9 2 9 1 9 7 1 9 2
17 9 1 9 4 1 9 13 13 0 9 9 9 7 0 0 9 2
13 0 0 9 4 3 13 13 13 3 2 0 9 2
20 9 9 3 13 2 16 9 9 15 1 10 9 13 7 13 1 9 0 9 2
3 9 13 9
3 0 11 2
18 12 7 9 9 9 9 7 0 9 13 3 0 9 0 11 1 9 2
14 13 15 0 9 1 9 10 0 9 0 9 1 11 2
14 1 1 9 9 1 0 9 15 9 13 3 1 9 2
27 9 1 0 11 15 3 3 13 1 11 2 1 0 11 2 11 2 11 2 10 9 1 0 9 7 11 2
16 3 15 13 13 2 16 1 11 4 1 9 0 9 11 13 2
31 0 9 15 1 9 9 13 3 2 0 0 9 1 9 9 2 15 13 0 9 9 9 0 7 3 9 2 16 0 9 2
4 0 9 1 11
2 0 9
7 11 2 11 2 11 2 2
40 10 9 3 4 13 1 15 2 16 2 0 0 9 2 3 3 13 9 7 16 0 10 0 9 13 13 1 9 2 14 2 14 9 9 7 9 0 0 9 2
31 3 13 1 9 2 15 15 13 3 1 9 0 7 0 0 9 7 15 1 0 9 13 2 13 1 15 1 10 9 0 2
14 1 3 0 9 15 13 2 10 13 3 9 7 9 2
14 3 14 13 7 0 9 7 1 15 7 0 0 9 2
101 1 0 9 4 13 0 9 2 16 11 1 0 2 9 2 2 0 2 9 2 14 13 13 7 13 3 2 1 9 1 11 2 3 13 11 2 11 7 11 2 7 13 7 1 11 7 1 11 2 3 13 1 9 15 2 11 1 0 9 2 13 9 0 9 2 7 13 2 16 4 0 9 7 11 13 1 0 9 9 2 1 15 15 13 2 16 9 2 0 9 2 13 1 11 1 9 2 14 0 2 2
39 16 9 9 1 9 10 9 1 10 9 7 10 9 2 13 9 2 15 4 1 0 9 13 1 9 11 2 11 2 0 9 9 11 1 0 9 9 2 2
23 9 4 3 13 1 9 2 3 1 9 2 16 9 13 10 9 0 9 2 13 1 9 2
7 0 9 11 2 11 2 11
3 9 1 11
5 11 2 11 2 2
32 9 0 9 11 2 11 15 3 13 1 12 9 9 0 0 9 2 11 2 2 15 13 1 9 0 0 9 1 11 1 11 2
14 9 7 9 9 3 1 9 13 3 9 11 11 11 2
2 0 9
5 11 2 11 2 2
2 0 9
26 0 9 1 9 11 13 1 9 9 11 1 0 9 1 11 9 1 9 12 9 7 9 1 12 9 2
14 1 9 13 1 9 9 7 1 11 9 4 13 9 2
26 0 9 13 0 9 9 1 9 9 9 1 11 2 3 13 9 2 12 9 2 12 9 7 12 9 2
14 9 3 13 9 1 0 9 2 3 3 4 13 9 2
30 0 0 9 1 9 1 9 13 1 9 3 1 9 1 0 9 1 11 9 11 2 16 4 15 13 1 11 7 3 2
10 13 1 15 13 9 1 0 9 9 2
19 1 0 9 1 9 0 9 11 1 11 13 3 0 9 3 16 12 9 2
6 11 11 1 11 1 11
4 13 4 1 15
15 1 9 4 13 1 9 0 0 9 0 9 0 11 11 2
18 10 9 13 3 3 0 2 2 0 2 2 2 16 15 13 0 13 2
35 15 1 9 2 15 4 15 3 13 2 4 7 13 3 0 1 9 1 9 2 7 1 9 2 1 0 0 9 1 12 2 12 2 12 2
18 1 10 9 13 3 9 13 4 1 15 2 15 3 13 7 1 11 2
18 3 3 13 10 0 2 9 2 1 11 11 15 16 9 9 2 2 2
14 2 13 15 2 16 0 9 11 13 9 10 0 9 2
24 13 9 11 2 15 13 3 0 9 16 9 0 9 2 9 0 9 13 1 11 10 0 9 2
15 1 0 9 4 13 15 1 0 9 1 9 1 0 9 2
17 7 15 3 1 10 9 4 13 1 0 9 2 13 9 2 2 2
14 2 13 11 1 9 3 0 2 7 3 0 1 9 2
11 15 13 1 15 9 11 1 10 0 9 2
14 11 0 10 9 2 9 7 9 13 0 0 9 9 2
23 2 13 15 1 15 2 9 11 2 16 13 9 0 0 9 11 1 0 9 7 1 11 2
36 3 15 2 9 13 13 2 2 13 2 10 13 0 9 2 7 13 15 9 2 7 16 4 15 15 13 2 4 15 13 1 10 0 0 9 2
29 0 13 13 1 12 2 7 3 15 3 13 2 10 0 9 4 13 10 0 9 13 2 16 4 15 13 13 9 2
5 13 3 9 0 2
5 13 0 15 13 2
51 1 0 9 9 9 11 4 15 3 13 13 2 16 15 10 9 13 1 0 2 7 0 9 9 7 13 10 9 3 1 10 9 0 9 2 15 2 3 13 2 2 7 2 3 7 3 13 3 0 9 2
24 7 15 13 13 1 15 9 2 3 13 9 12 2 7 16 13 9 3 0 2 7 9 12 2
44 2 13 13 0 7 0 9 0 9 2 16 4 7 15 2 15 15 13 1 9 1 11 2 13 2 3 0 13 9 0 2 3 0 2 7 0 2 0 2 9 9 2 2 2
32 13 4 9 1 12 0 9 7 13 9 2 15 4 13 2 16 4 9 0 9 2 15 13 3 0 2 15 13 1 0 9 2
13 3 13 1 0 2 0 0 9 2 15 13 13 2
9 14 10 9 15 3 13 0 9 2
14 7 3 13 9 1 0 9 2 1 0 0 0 9 2
30 15 13 9 7 3 3 7 9 2 16 4 1 0 9 3 13 2 16 10 9 15 3 13 13 3 1 11 7 11 2
2 11 11
17 9 0 11 3 13 2 16 9 11 13 2 0 9 0 9 2 2
18 1 11 9 0 9 13 2 16 2 13 13 0 9 9 1 11 2 2
35 9 1 11 2 3 0 9 13 1 0 9 0 0 9 2 13 2 16 2 9 13 2 15 13 1 15 0 2 7 3 13 10 9 2 2
16 7 1 10 9 15 7 1 0 0 9 13 9 1 0 9 2
27 0 9 9 13 2 16 16 11 13 0 9 2 3 15 0 0 9 7 9 1 0 9 4 13 13 9 2
36 0 9 0 2 11 13 2 16 9 11 13 16 2 9 2 15 13 0 11 7 13 15 13 1 0 0 7 0 9 1 11 7 1 11 2 2
24 2 15 2 16 11 3 13 1 9 0 9 0 0 9 2 13 10 9 9 1 9 0 9 2
12 0 9 15 13 2 2 13 3 0 9 11 2
24 7 13 0 9 0 9 2 16 13 9 13 15 1 12 9 9 2 15 13 0 9 0 9 2
38 1 9 0 11 1 11 13 3 0 9 0 13 15 2 16 4 0 9 13 1 0 9 9 2 13 7 2 16 4 1 0 11 13 9 1 0 9 2
34 2 13 15 9 2 15 13 0 9 2 16 4 1 12 2 9 12 13 9 0 9 9 2 16 3 0 7 0 9 2 2 13 9 2
54 2 7 15 15 13 13 2 16 4 9 0 9 2 15 16 0 3 12 9 13 2 13 9 0 9 2 4 13 7 3 9 2 16 4 13 0 9 2 16 1 0 9 13 14 12 9 0 9 2 2 13 15 9 2
36 13 12 2 9 0 9 13 1 0 9 1 9 9 0 9 0 9 11 2 11 2 0 0 9 9 13 1 9 2 15 11 1 10 9 13 2
15 1 10 9 4 13 9 13 15 9 0 0 9 7 9 2
16 3 12 9 3 1 0 11 13 1 9 1 0 3 0 9 2
27 3 9 13 13 1 0 0 9 11 2 3 1 0 9 13 1 9 12 9 2 0 9 7 13 12 0 2
11 0 9 13 1 9 1 9 9 0 9 2
9 13 15 1 9 9 11 2 11 2
29 1 9 15 13 2 16 9 13 2 16 4 13 9 13 0 9 1 0 9 7 9 9 1 9 0 0 0 9 2
24 1 9 13 1 11 13 12 9 2 1 15 3 12 0 9 11 2 11 2 9 9 0 11 2
10 4 13 12 0 9 1 0 9 11 2
5 9 9 13 0 2
12 13 3 12 2 9 0 1 11 1 9 12 2
32 1 10 9 1 9 1 9 2 15 15 13 13 1 9 2 13 3 9 9 9 1 0 9 0 0 9 11 2 11 10 9 11
15 0 9 13 1 0 9 0 9 1 9 9 1 0 11 2
15 13 15 0 0 9 7 0 9 11 2 11 1 0 9 2
23 13 2 16 11 15 13 1 3 0 9 2 16 13 13 10 9 1 11 7 0 0 9 2
11 11 13 1 0 9 3 3 1 12 3 2
42 1 9 3 13 9 2 1 15 13 0 9 3 0 9 0 12 9 2 15 15 13 1 11 7 3 3 13 7 1 10 9 15 3 12 3 1 11 13 7 13 3 2
18 0 9 2 15 15 13 1 9 0 9 2 13 13 9 3 0 9 2
12 1 0 1 12 9 13 14 1 12 0 9 2
20 0 9 13 3 14 3 1 15 2 16 9 13 13 7 1 9 1 9 9 2
16 9 9 1 9 0 11 3 13 9 1 0 11 1 12 9 2
23 1 9 0 9 15 3 1 0 9 13 12 9 9 15 9 2 1 15 3 12 9 0 2
15 1 9 1 0 9 13 1 11 0 0 9 1 0 9 2
24 1 9 9 3 13 9 0 9 2 15 13 11 1 9 9 1 9 3 1 0 9 1 11 2
27 0 9 9 1 9 2 15 3 1 9 10 9 13 0 9 1 9 1 9 0 9 2 10 9 3 13 2
19 10 9 13 3 0 2 16 13 2 16 15 1 11 3 13 16 0 9 2
28 12 9 3 7 0 0 9 15 13 12 0 9 1 11 2 15 0 9 13 1 9 10 0 9 9 1 9 2
23 0 9 13 1 9 9 9 2 9 9 1 9 10 9 9 7 13 1 9 0 0 9 2
2 9 9
2 9 9
2 11 2
15 3 0 9 9 2 3 12 2 13 1 9 1 9 12 2
25 15 13 1 0 9 2 7 0 15 13 9 0 9 2 9 7 9 2 13 1 11 0 9 9 2
38 1 9 10 0 9 0 9 15 3 0 9 13 9 0 11 2 3 13 13 12 9 2 7 11 2 3 12 9 13 1 9 9 1 0 9 9 11 2
27 9 11 11 11 13 2 16 10 9 0 9 1 11 2 13 13 3 2 7 3 2 16 13 1 9 2 2
23 0 9 1 9 13 0 11 2 3 15 3 13 12 2 1 12 1 11 7 12 1 11 2
18 12 9 13 1 9 1 0 9 7 1 9 2 15 1 15 3 13 2
7 2 9 9 13 3 0 2
15 10 9 9 13 0 2 2 13 9 0 9 11 11 11 2
42 1 0 9 0 9 13 0 9 2 15 13 1 10 9 2 1 9 13 1 0 9 9 1 0 9 2 1 12 9 2 7 1 0 0 9 1 9 2 12 9 2 2
4 9 11 2 11
2 11 11
5 0 9 2 2 2
39 1 9 2 16 15 3 2 16 3 13 11 2 13 1 11 2 11 2 7 15 0 2 0 0 9 9 13 2 2 14 13 0 9 2 7 13 15 13 2
15 13 13 2 13 15 2 1 11 7 13 15 16 1 9 2
8 9 9 13 3 0 7 0 2
23 15 2 15 13 9 1 11 2 11 2 15 1 10 9 3 13 2 10 0 9 13 2 2
50 3 15 1 10 15 13 2 16 15 11 7 0 13 13 2 16 4 1 9 13 9 7 13 1 9 9 7 9 1 9 2 13 0 0 9 9 11 11 1 9 2 15 3 13 0 9 11 0 11 2
5 0 9 13 9 9
3 9 9 13
23 9 9 15 3 13 2 13 15 9 0 9 0 9 0 0 9 7 9 9 1 0 9 2
38 0 0 9 13 9 2 16 0 9 15 1 0 12 9 13 3 1 12 9 11 2 15 13 14 9 0 9 2 15 1 9 0 9 13 9 0 9 2
28 9 0 9 7 9 15 1 0 9 13 14 1 12 2 12 9 2 7 3 1 12 9 2 3 13 10 9 2
9 9 0 9 3 13 3 3 13 2
27 9 0 9 13 13 1 0 9 2 15 13 9 0 9 1 0 9 1 9 9 1 9 9 7 9 9 2
26 0 0 9 13 9 9 13 9 7 13 9 0 9 2 15 13 1 9 9 2 13 0 9 2 2 2
5 15 9 13 1 9
10 0 9 10 0 9 13 9 1 9 2
24 7 13 15 2 16 9 9 13 3 15 0 9 2 15 15 13 13 9 7 2 13 9 2 2
6 15 15 15 3 13 2
10 0 9 0 9 13 10 9 0 9 2
20 7 1 9 0 9 10 9 13 0 9 2 0 1 9 9 9 9 9 9 2
4 7 3 9 2
11 13 15 13 1 9 9 0 0 2 9 2
32 13 14 13 2 16 9 0 7 0 9 1 0 9 2 3 15 3 0 9 13 1 9 0 0 9 9 2 3 13 9 9 2
40 10 0 9 13 13 2 9 2 16 9 13 0 15 13 1 9 2 9 7 9 2 16 9 13 0 14 1 0 9 2 9 2 16 9 7 9 15 13 15 2
13 0 9 13 9 3 13 1 9 9 7 0 9 2
34 12 0 9 2 0 1 9 1 9 2 3 13 2 16 9 2 16 15 9 13 2 3 14 15 2 16 15 1 9 3 1 15 13 2
4 13 15 9 2
15 11 7 11 13 0 2 7 13 2 16 0 2 0 9 2
8 13 15 9 2 0 0 9 2
7 14 3 2 7 1 9 2
11 7 10 9 15 13 9 1 9 0 9 2
6 3 9 11 13 0 2
12 12 2 9 15 9 13 9 9 1 0 11 2
17 1 10 9 2 15 1 0 9 13 9 3 0 2 13 9 9 2
7 1 0 9 0 12 9 2
10 3 1 9 12 0 9 3 3 13 2
16 1 11 2 9 9 2 13 9 2 0 15 3 1 0 9 2
9 13 15 9 1 9 1 0 11 2
16 12 0 9 15 13 1 9 9 2 15 15 3 13 1 11 2
7 7 3 1 3 0 9 2
11 13 1 9 9 2 13 1 9 0 9 2
15 15 13 1 0 9 2 0 9 9 7 0 9 9 9 2
10 15 3 13 9 2 15 3 3 13 2
8 13 15 9 1 9 1 9 2
14 13 15 9 9 2 15 15 13 1 0 9 0 9 2
6 3 7 3 13 13 2
20 13 13 2 16 0 9 13 9 0 7 3 0 9 13 13 0 0 0 9 2
24 1 0 9 15 1 9 13 0 0 9 2 16 3 13 9 2 0 9 3 0 1 0 9 2
27 15 13 9 2 13 2 3 0 15 4 13 9 1 0 9 2 7 3 2 16 15 4 13 0 9 9 2
13 0 9 1 9 2 0 0 2 13 3 3 0 2
22 16 9 13 10 9 2 16 15 4 13 12 9 2 13 1 9 9 1 12 9 9 2
8 13 0 1 10 9 13 9 2
6 3 9 13 1 9 2
10 1 9 9 0 9 13 13 15 0 2
12 13 0 9 9 2 15 15 13 9 9 9 2
12 13 9 1 9 7 13 15 10 0 0 9 2
16 1 15 13 9 0 3 16 1 9 1 0 11 1 0 9 2
24 3 1 0 9 2 15 15 13 1 9 1 9 0 9 2 7 1 15 2 15 12 9 13 2
5 7 9 0 13 2
17 9 9 9 13 9 1 9 0 0 9 2 0 9 9 0 9 2
19 9 1 9 7 1 9 13 13 1 9 0 9 1 0 7 0 9 9 2
11 9 12 2 13 1 9 2 9 0 9 2
23 0 9 4 13 9 2 11 11 13 9 0 9 2 7 9 1 9 7 9 4 13 9 2
18 9 4 13 2 10 9 13 2 15 13 2 16 15 4 3 13 9 2
11 9 12 2 9 3 1 15 13 9 9 2
12 7 3 15 13 13 2 15 9 13 1 9 2
10 14 1 15 13 9 3 0 7 0 2
2 11 11
10 1 9 0 9 1 11 13 9 0 9
4 9 1 0 9
33 16 0 2 11 0 2 0 9 13 12 2 9 1 11 0 9 1 12 0 9 2 13 15 1 15 0 9 2 14 9 0 9 2
13 1 0 9 0 0 0 9 15 13 15 0 9 2
33 1 0 9 1 0 9 1 0 9 14 1 0 9 2 15 7 3 4 15 13 2 15 13 3 10 9 2 15 3 0 9 3 2
16 12 9 4 7 3 13 2 9 9 10 2 15 13 9 13 2
22 3 3 0 9 0 9 9 11 15 3 1 0 9 1 9 1 0 11 13 9 13 2
16 13 15 7 7 9 1 0 9 9 0 9 15 13 13 0 2
53 11 11 2 9 11 2 1 15 15 13 2 16 4 13 11 11 2 13 7 1 9 2 14 9 1 9 2 3 13 1 9 7 3 9 9 13 15 2 16 4 15 0 9 13 1 9 1 10 9 3 0 9 2
25 10 9 14 13 2 16 1 0 9 13 15 1 9 2 7 3 3 11 13 1 9 0 9 9 2
26 1 10 9 16 4 15 9 13 13 9 7 9 1 9 13 2 16 13 1 0 9 1 0 9 9 2
19 10 9 13 3 13 1 9 0 9 7 13 0 9 9 9 9 11 11 2
29 9 3 13 9 9 2 15 1 12 9 13 9 1 9 2 16 1 9 9 13 15 1 9 2 3 7 13 9 2
29 9 2 15 15 1 11 13 1 9 3 12 9 2 13 1 0 10 9 0 9 1 9 0 9 3 1 0 9 2
12 10 9 3 13 10 9 13 15 3 13 9 2
33 3 13 3 3 2 3 10 9 3 13 2 16 13 9 9 0 1 9 2 15 3 3 15 13 2 3 3 13 9 9 0 9 2
22 10 9 3 13 7 0 9 13 9 3 2 16 4 15 13 13 0 9 0 0 9 2
4 9 13 9 2
21 0 9 15 3 13 1 0 9 2 3 13 13 7 3 7 13 2 7 13 15 2
8 3 1 9 13 1 0 9 2
25 9 13 2 16 13 3 3 3 1 9 2 16 15 7 13 15 2 1 15 13 0 9 1 9 2
19 9 11 11 3 13 0 9 2 16 13 0 9 7 9 15 13 13 9 2
10 10 9 13 2 3 7 10 9 13 2
19 1 10 9 9 13 3 0 9 7 1 9 15 13 15 9 9 0 9 2
21 0 0 9 4 13 7 9 3 13 10 3 0 9 7 1 0 9 7 9 9 2
26 15 13 9 9 2 3 9 13 2 16 15 2 15 3 3 13 0 9 2 13 0 9 7 13 9 2
21 9 9 10 9 15 13 1 9 2 3 15 7 13 1 12 0 7 0 9 0 2
16 0 7 3 0 9 9 15 13 7 1 0 11 13 0 9 2
13 0 9 3 13 9 2 16 13 9 0 0 9 2
33 9 9 1 9 9 13 9 12 9 9 11 1 9 2 9 11 11 4 13 9 9 11 11 7 9 11 11 9 9 9 7 9 2
21 9 9 13 1 9 10 0 9 2 1 0 3 0 9 9 7 0 9 11 11 2
10 10 9 15 1 10 9 13 1 9 2
34 11 11 2 15 15 13 0 9 1 0 11 13 9 0 0 9 2 7 3 1 9 13 9 1 3 0 7 3 15 13 13 1 9 2
18 1 9 0 0 9 15 15 15 13 7 3 1 9 13 1 9 9 2
28 1 10 9 3 9 13 7 0 0 9 13 2 16 15 12 9 13 1 9 1 0 9 3 0 9 9 11 2
28 15 7 13 0 12 0 9 1 9 2 3 1 9 13 9 2 1 15 15 1 9 9 3 13 2 3 13 2
13 7 1 11 13 13 9 2 9 9 2 9 0 2
2 11 11
7 9 1 9 9 11 11 9
8 10 9 9 15 4 13 9 2
15 13 15 0 9 2 1 12 9 9 1 0 9 12 9 2
22 13 4 15 0 9 2 1 12 5 1 9 0 9 7 14 1 12 5 1 0 9 2
9 13 15 15 9 7 13 0 9 2
26 13 15 2 16 1 9 13 0 9 2 15 4 3 13 1 9 9 1 9 12 2 3 3 1 9 2
11 7 4 15 13 9 15 1 0 9 13 2
26 16 3 2 3 4 1 9 13 3 2 4 13 9 0 16 3 2 14 0 3 0 9 4 3 13 2
12 13 4 3 0 7 0 9 16 1 9 12 2
12 9 0 9 15 3 13 2 16 15 9 13 2
23 15 13 0 0 9 2 9 15 13 2 13 10 9 2 15 13 0 7 15 15 13 13 2
22 13 7 1 15 2 16 4 9 9 2 2 9 9 2 13 1 15 0 9 3 0 2
43 10 9 9 15 13 7 0 9 2 9 2 16 3 9 0 7 0 9 13 13 2 16 1 0 9 1 0 9 15 10 9 13 7 0 9 9 15 1 0 9 13 13 2
18 3 15 13 13 2 16 9 0 9 13 1 9 2 7 15 13 9 2
3 2 11 2
9 12 2 11 2 15 6 2 3 2
9 3 15 13 1 0 9 2 16 2
9 2 11 2 11 7 11 2 11 2
16 12 2 16 13 3 2 13 15 1 0 2 3 0 9 3 2
9 2 11 2 11 7 11 2 11 2
4 12 2 11 2
2 11 2
5 6 15 13 9 2
2 11 2
5 2 11 2 11 2
10 12 2 13 2 13 2 3 15 13 2
9 2 11 2 11 7 11 2 11 2
4 12 2 0 2
6 7 14 1 12 9 2
9 2 11 2 11 7 11 2 0 2
4 12 2 13 2
5 2 11 2 11 2
7 12 2 0 9 2 2 2
5 15 3 13 0 2
5 2 11 2 11 2
9 2 11 2 11 7 11 2 11 2
4 12 2 11 2
8 15 13 3 1 9 2 2 2
5 2 11 2 11 2
15 9 2 11 11 2 11 11 2 11 11 2 11 11 2 11
2 15 2
3 3 2 3
25 9 0 11 13 12 2 12 2 11 9 2 12 2 12 2 0 9 7 12 2 12 2 0 9 2
9 9 9 1 9 9 1 12 9 2
7 9 0 9 13 0 9 2
40 12 2 12 2 2 12 2 11 1 0 9 7 0 9 2 12 2 12 2 12 2 12 2 0 9 1 9 11 2 11 7 11 2 11 2 13 11 11 2 2
20 11 9 2 0 12 2 11 12 2 13 9 9 0 9 2 3 1 12 2 2
38 12 2 12 2 13 11 11 2 12 2 12 2 11 11 2 11 2 12 2 12 2 11 2 11 7 11 2 11 2 12 2 12 2 11 11 2 11 2
27 11 9 7 9 11 13 9 0 9 2 9 9 7 9 10 7 0 9 2 1 12 2 12 2 1 12 2
2 12 2
13 9 13 13 0 9 1 9 2 11 7 0 9 2
20 0 0 9 11 11 13 12 2 12 2 12 1 9 11 0 9 2 12 2 2
11 1 11 13 13 9 11 11 2 11 2 2
14 9 2 9 9 2 0 9 12 2 12 12 11 12 2
2 0 9
19 1 9 0 7 1 9 0 9 15 3 3 0 0 9 13 0 7 0 2
10 3 13 0 9 7 13 15 1 15 2
11 13 9 1 0 9 2 13 1 0 9 2
17 9 2 1 9 2 15 13 1 9 2 15 13 0 16 11 11 2
21 1 0 9 1 9 2 12 1 11 1 11 13 9 0 9 2 7 7 9 0 2
21 3 13 9 9 7 1 0 9 13 0 9 9 9 1 9 7 9 9 11 12 2
19 3 2 1 12 2 9 2 13 0 13 3 9 1 0 9 1 0 13 2
18 9 12 9 13 9 1 10 9 2 7 15 7 13 13 9 0 9 2
40 0 9 7 0 9 0 9 13 11 11 2 9 9 2 12 2 2 13 15 11 11 2 0 9 13 9 11 2 9 9 2 12 2 7 0 9 13 11 11 2
12 11 11 1 0 9 10 9 13 9 10 9 2
12 1 9 0 15 15 13 13 0 9 9 0 2
17 3 0 9 11 11 13 0 0 9 11 9 0 9 12 2 9 2
27 1 15 2 16 1 0 9 13 9 2 13 9 11 11 1 10 9 1 9 2 3 7 3 3 3 2 2
14 13 9 7 13 3 13 1 9 0 9 2 7 3 2
3 2 11 2
5 9 11 11 2 11
3 13 1 11
3 9 1 9
21 3 1 9 2 12 2 12 2 2 13 1 11 0 0 9 2 3 0 0 9 2
30 1 0 9 15 13 3 10 0 9 2 9 11 2 9 11 3 2 2 2 3 7 10 9 2 3 2 9 11 2 2
15 14 10 0 9 2 14 3 0 2 13 2 3 1 9 2
22 0 9 13 0 9 1 11 2 1 3 0 11 2 2 1 0 15 13 0 11 11 2
58 13 9 0 9 2 11 2 11 2 15 13 9 1 11 1 11 12 2 16 4 3 2 13 0 0 9 0 9 7 0 9 2 1 9 0 11 2 0 1 9 2 15 13 10 0 9 7 0 2 6 2 1 3 3 0 9 2 2
14 0 9 9 3 13 0 9 2 9 9 1 0 9 2
34 11 2 11 13 3 0 9 2 11 2 11 0 7 0 9 2 9 2 0 11 2 11 2 15 13 13 1 12 2 9 9 0 9 2
27 15 13 2 16 0 7 3 2 2 7 10 9 2 2 9 7 9 13 14 3 7 10 9 13 3 0 2
40 16 13 3 0 0 9 0 9 2 9 0 9 15 3 2 13 2 2 3 3 15 11 2 11 2 11 2 7 11 2 11 2 11 2 13 1 3 0 9 2
12 3 0 9 13 3 0 9 9 7 0 9 2
46 3 0 13 11 2 11 2 11 2 2 1 0 9 13 0 7 0 9 11 2 11 2 9 2 11 2 2 3 16 0 11 2 11 2 11 2 7 0 9 11 2 11 2 11 2 2
11 11 2 11 3 13 9 9 2 11 2 2
33 1 0 9 1 9 3 13 11 2 11 2 9 2 11 2 2 11 2 11 2 11 2 7 3 3 0 11 2 11 2 11 2 2
24 0 9 13 9 0 2 0 9 2 11 0 9 2 11 2 11 13 0 9 7 0 0 9 2
7 3 0 13 3 3 2 2
14 0 9 9 13 7 0 0 9 2 7 0 15 9 2
30 1 0 9 7 9 13 9 2 0 11 2 11 2 13 15 7 3 7 9 1 9 2 9 7 9 2 13 3 0 2
55 13 2 14 13 9 11 2 11 2 9 1 9 2 2 2 2 2 2 15 15 10 9 2 13 2 2 9 2 7 13 2 16 2 2 2 2 9 2 15 3 4 13 2 1 0 9 13 2 10 9 1 9 9 2 2
29 3 2 9 15 13 13 7 13 2 2 3 11 2 2 15 15 15 14 13 14 1 9 9 1 0 9 7 9 2
7 3 1 9 13 3 9 2
2 11 11
6 11 1 11 1 10 9
2 0 9
47 1 9 3 0 9 2 15 1 15 1 0 9 13 1 11 3 11 2 3 13 9 10 9 2 11 2 9 13 3 16 12 9 0 9 0 9 11 11 11 1 11 2 11 1 11 2 2
52 7 3 3 13 1 10 9 13 9 2 1 15 12 9 0 9 13 0 9 2 9 2 9 7 9 9 2 7 0 9 0 9 2 9 2 1 15 9 9 7 9 13 3 3 3 16 0 9 1 0 9 2
46 11 1 11 13 9 1 15 2 15 13 0 9 1 9 7 15 14 9 2 1 0 9 1 0 2 1 9 9 2 15 13 0 1 0 9 13 1 10 9 2 1 9 2 15 13 2
8 0 9 13 3 9 1 9 2
30 0 9 13 10 0 9 2 15 3 13 9 7 13 10 0 13 1 9 1 0 0 9 9 1 9 7 9 11 11 2
18 10 9 9 15 7 13 0 9 2 15 10 9 13 0 9 15 3 2
39 16 15 7 7 1 0 9 1 0 9 2 1 9 3 11 2 9 1 11 3 13 0 2 3 7 3 13 9 10 2 9 2 2 9 1 9 9 13 2
19 1 9 4 7 13 9 7 9 11 2 11 11 2 2 15 10 9 13 2
15 11 15 13 13 0 0 9 1 9 7 0 9 0 9 2
42 3 1 10 9 13 7 0 2 0 9 9 2 0 9 13 13 9 0 2 15 15 13 1 9 7 1 15 9 3 3 13 13 9 7 13 15 14 0 9 0 9 2
8 9 2 3 13 1 9 0 2
16 11 1 11 2 9 2 15 13 13 2 1 10 9 3 13 2
19 13 14 2 16 15 0 0 9 13 1 15 1 9 2 1 9 9 2 2
2 11 11
2 0 9
3 3 1 9
65 12 0 0 9 1 0 9 2 1 15 3 13 0 9 9 0 2 9 2 9 2 9 2 9 1 9 11 2 11 11 2 11 2 9 11 2 11 2 1 0 9 3 0 7 0 11 2 11 2 14 0 11 2 11 1 3 0 3 0 9 9 9 7 9 2
72 2 7 12 0 9 1 0 9 2 0 0 9 0 1 0 9 2 0 0 9 0 9 2 2 3 0 9 0 9 2 7 3 0 2 9 1 0 9 2 2 9 1 9 2 0 2 7 0 2 0 9 11 2 11 2 3 0 9 11 2 11 2 1 12 1 0 9 0 11 2 11 2
27 12 9 0 9 2 10 0 2 0 9 15 13 13 3 14 9 9 1 9 2 3 0 2 3 0 2 2
8 3 15 13 12 9 3 0 2
50 13 7 1 15 14 9 0 7 0 2 13 15 3 9 9 0 2 11 13 3 1 9 1 2 9 0 9 2 2 7 0 3 0 2 3 14 3 0 9 2 7 3 3 0 9 9 1 0 9 2
96 16 3 9 9 2 9 2 9 1 9 0 9 2 0 0 9 2 0 0 9 9 3 2 2 13 9 9 2 10 0 9 9 2 6 2 9 2 2 2 2 2 2 10 9 13 3 1 9 13 2 7 2 3 1 15 13 2 3 1 3 0 9 2 15 13 1 10 0 9 7 9 3 13 1 15 9 9 2 11 13 9 16 0 0 9 3 7 3 3 2 16 13 3 0 9 2
40 3 0 2 3 0 9 0 9 13 3 9 10 9 7 10 0 9 2 13 3 0 9 1 0 2 0 0 2 9 7 3 0 9 2 9 1 9 2 13 2
27 9 2 3 3 13 9 9 2 7 3 9 0 3 1 0 9 9 0 9 15 13 3 13 10 9 3 2
21 3 13 2 0 9 4 15 1 9 11 9 3 13 0 0 9 1 0 9 9 2
18 1 0 9 15 13 0 9 2 9 15 0 2 0 9 7 0 9 2
2 11 11
5 0 9 1 9 9
3 10 0 11
7 1 9 13 9 12 9 2
78 10 0 2 1 12 2 9 10 2 9 2 2 13 9 11 11 7 9 11 11 0 9 9 9 11 11 2 13 15 1 15 1 2 9 9 1 9 3 12 2 12 2 2 3 1 0 9 2 1 9 9 2 9 9 7 9 2 1 9 9 2 7 13 1 9 3 13 2 3 9 0 9 2 2 13 9 2 2
39 9 11 2 11 1 12 2 9 13 0 9 2 1 0 7 0 9 9 2 15 13 1 0 2 2 7 13 2 4 7 13 9 1 15 13 2 2 2 2
26 13 0 9 1 3 0 7 0 9 0 7 0 9 2 15 13 9 2 3 0 9 2 3 7 13 2
32 0 9 4 13 13 9 2 3 0 9 2 1 15 0 9 13 9 9 9 7 15 4 15 13 1 12 2 9 13 0 9 2
31 13 3 9 2 15 15 3 13 9 0 9 2 0 9 2 9 3 2 2 7 13 13 9 2 15 9 11 2 11 13 2
74 0 9 1 9 9 1 0 9 2 13 9 2 16 11 2 11 13 1 2 10 0 11 2 15 13 1 0 11 3 0 7 15 15 13 2 2 2 0 9 0 7 1 0 9 2 7 9 1 12 9 2 3 3 13 13 0 9 2 2 14 3 13 1 9 3 11 2 11 2 3 11 2 11 2
26 11 2 11 7 11 2 11 9 13 1 0 9 2 1 9 0 2 2 0 9 1 0 9 1 11 2
21 10 9 13 9 1 0 9 2 15 15 0 9 13 2 13 15 1 3 12 9 2
56 9 13 2 16 11 2 11 1 9 2 3 1 9 0 9 13 2 3 13 10 0 0 9 2 7 16 2 1 9 2 9 15 13 3 16 9 9 7 1 10 9 4 13 3 13 9 2 15 9 2 1 9 2 13 2 2
48 1 9 1 13 15 11 11 7 13 0 9 2 7 9 2 15 3 3 13 9 0 9 2 0 9 9 11 2 3 1 9 12 15 13 9 13 2 2 7 7 13 0 2 7 9 0 9 2
28 13 3 13 1 0 9 0 9 2 16 15 13 9 0 9 2 1 2 0 9 2 13 2 3 2 13 2 2
25 3 13 2 0 13 1 10 9 3 9 2 16 0 2 9 2 7 0 9 3 10 0 9 13 2
3 2 11 2
21 2 0 2 9 11 11 2 10 0 2 9 2 15 13 0 9 1 9 0 9 2
10 10 0 15 13 13 2 9 11 2 2
5 9 11 11 2 11
6 11 11 1 9 0 11
3 0 9 9
20 9 9 2 3 15 13 3 13 9 0 0 9 1 9 9 0 9 11 11 2
14 9 2 15 13 0 7 0 1 10 9 7 9 9 2
12 9 2 15 3 3 1 10 9 13 1 9 2
13 9 13 7 0 0 9 7 9 0 9 11 11 2
7 13 1 9 0 11 3 2
9 9 9 13 10 9 1 0 9 2
10 3 15 13 1 0 0 9 0 11 2
13 0 11 7 10 0 9 15 13 13 16 0 9 2
7 13 15 1 0 9 9 2
15 13 9 10 9 2 15 15 1 15 1 10 9 13 13 2
4 9 13 0 2
24 12 2 9 2 2 0 9 2 2 9 2 15 7 15 2 3 13 9 2 15 13 0 13 2
22 7 15 15 13 13 14 9 3 0 0 9 2 15 15 3 13 13 0 9 1 9 2
10 13 3 0 9 1 0 9 16 15 2
8 3 10 9 13 9 1 11 2
13 0 9 3 1 11 1 11 7 0 9 1 11 2
27 12 2 9 2 9 2 0 2 0 0 9 2 15 15 3 13 1 9 2 15 13 1 0 0 9 13 2
11 3 1 9 2 3 3 1 0 0 9 2
15 1 11 15 13 9 11 2 1 11 0 9 2 2 2 2
30 12 2 9 2 0 9 2 13 10 0 7 0 9 2 9 14 3 15 0 7 3 0 2 1 9 13 0 9 9 2
22 1 9 15 13 1 9 1 9 7 15 15 2 14 1 9 2 13 10 0 0 9 2
18 0 9 15 13 3 1 15 2 13 9 2 16 4 13 13 2 2 2
7 13 9 0 9 9 9 2
23 7 13 15 0 9 9 2 15 15 13 9 9 2 9 15 9 2 9 2 9 2 2 2
4 3 13 9 2
5 9 13 0 9 2
7 0 0 9 7 15 0 2
21 0 0 9 0 2 16 9 9 2 0 9 2 2 13 7 3 3 13 2 0 2
28 9 13 2 3 15 0 9 3 13 2 9 9 7 9 13 9 9 2 3 13 13 13 0 9 9 10 9 2
16 13 15 0 1 12 9 9 7 0 9 1 9 0 9 9 2
10 10 9 7 13 3 3 1 0 9 2
10 0 9 13 0 11 7 10 0 9 2
16 13 15 15 12 0 9 7 10 2 9 2 13 12 5 9 2
21 13 3 9 9 10 9 2 9 9 1 9 7 7 9 10 9 1 0 0 9 2
6 0 9 13 7 0 2
15 7 10 9 13 3 7 1 11 2 16 13 10 0 9 2
11 0 9 7 14 14 3 13 9 1 15 2
10 13 4 13 10 9 0 9 1 11 2
11 0 9 11 15 13 0 9 1 10 9 2
10 9 13 0 2 7 9 13 3 0 2
6 9 13 9 7 9 2
6 3 11 13 9 0 2
21 1 0 9 0 13 10 9 2 1 0 3 1 15 13 14 12 0 1 0 9 2
10 7 11 13 9 1 0 7 0 9 2
8 0 9 3 13 7 13 9 2
17 9 11 3 10 9 1 15 13 2 16 0 9 13 0 0 9 2
3 15 3 2
5 15 1 15 13 2
4 3 15 13 2
6 9 15 4 13 9 2
10 3 7 2 16 11 13 9 2 9 2
30 1 11 13 9 2 16 0 9 13 9 11 1 11 7 11 1 11 2 15 4 13 1 9 9 2 9 1 9 2 2
26 13 3 7 9 0 9 2 16 0 9 0 1 0 9 2 7 15 4 4 3 0 9 2 13 2 2
11 9 7 9 2 3 15 13 2 13 10 2
24 3 2 7 15 13 2 16 13 13 13 2 15 13 1 0 9 13 3 7 1 0 9 3 2
16 3 15 13 9 9 1 10 0 0 9 2 15 15 15 13 2
24 0 9 2 15 1 0 11 13 2 13 9 0 2 13 15 9 2 15 13 0 9 2 9 2
26 13 1 10 0 9 3 15 0 1 0 7 0 9 2 7 1 3 0 9 9 1 0 9 7 9 2
15 3 1 10 0 9 15 9 3 13 7 13 0 0 9 2
15 13 15 2 16 15 15 13 7 13 1 15 3 3 0 2
40 1 9 7 1 10 9 13 2 3 3 15 3 3 13 9 11 11 2 0 9 9 2 2 15 3 13 9 10 2 9 2 9 2 3 3 13 1 9 9 2
52 10 9 13 0 9 2 0 9 3 13 10 9 9 0 9 2 9 2 11 2 2 2 2 2 7 1 9 2 3 15 1 0 9 13 12 9 9 2 11 2 2 15 13 3 7 9 13 1 9 0 9 2
17 3 0 2 3 14 2 0 2 9 2 2 7 3 9 1 9 2
20 7 1 15 15 13 0 9 3 3 13 2 16 0 9 13 15 3 3 9 2
12 3 3 13 0 2 15 13 9 7 15 14 2
10 0 9 2 12 2 3 13 0 9 2
6 12 2 3 13 0 2
17 3 13 13 15 9 2 9 2 9 2 7 13 1 15 13 9 2
7 15 15 13 1 0 9 2
43 0 10 9 2 15 2 13 2 7 2 13 2 2 3 14 1 9 12 2 13 9 2 0 2 13 14 2 15 4 15 13 1 11 2 2 7 3 15 13 1 0 9 2
13 16 13 9 0 11 2 15 3 13 1 0 11 2
19 3 2 16 15 13 1 9 10 9 7 3 15 13 1 3 0 0 9 2
39 3 13 13 2 16 9 1 11 7 11 13 7 9 0 0 9 1 9 1 9 2 7 13 0 9 0 9 2 3 2 11 5 11 5 11 2 9 2 2
7 13 15 9 9 0 9 2
12 7 3 15 13 2 3 13 9 1 9 2 2
12 10 9 13 13 9 9 2 16 4 15 13 2
5 7 3 1 15 2
11 3 3 15 10 9 9 13 3 16 9 2
3 1 11 2
2 14 2
15 7 13 15 7 9 9 15 1 0 9 2 0 9 9 2
16 1 15 13 3 14 0 9 2 7 7 0 2 0 7 0 2
15 3 3 3 13 13 0 11 1 11 2 13 4 15 9 2
9 3 15 13 0 11 1 0 9 2
10 0 9 2 15 13 0 0 0 9 2
7 14 3 1 0 11 13 2
19 3 13 9 9 9 13 1 9 9 9 2 0 2 0 2 2 2 2 2
17 1 11 13 1 10 9 0 9 2 9 2 9 2 9 2 9 2
16 13 3 0 9 0 9 7 1 15 3 3 9 3 13 9 2
31 10 9 13 1 15 0 2 16 15 13 2 16 3 9 13 3 2 16 0 2 9 2 11 2 11 2 2 2 2 2 2
10 7 9 13 9 16 0 9 1 15 2
10 3 4 3 13 1 0 9 1 9 2
35 15 15 1 10 9 13 3 3 2 2 1 15 15 13 0 2 13 1 0 9 2 10 9 13 2 9 2 2 11 13 1 15 0 9 2
13 15 13 0 9 2 15 13 15 3 0 13 2 2
7 11 2 15 13 7 9 2
2 9 2
7 9 16 9 9 9 9 2
14 3 3 13 14 12 9 7 15 15 13 3 3 13 2
12 9 1 0 9 7 0 9 0 9 13 9 2
21 0 9 15 13 3 10 0 9 13 15 7 15 1 15 15 13 16 0 1 9 2
9 7 13 15 1 15 1 0 9 2
8 9 9 11 13 0 0 9 2
12 7 3 3 2 13 2 7 0 11 1 11 2
12 1 10 9 13 9 9 16 0 9 3 13 2
8 9 11 2 3 13 15 0 2
16 13 15 3 1 9 9 7 0 9 2 15 13 13 1 9 2
10 9 15 13 13 16 9 2 0 9 2
12 9 2 9 2 9 2 9 2 9 2 2 2
8 15 4 3 13 10 0 9 2
11 1 10 9 13 9 1 9 9 13 15 2
25 1 10 9 15 13 13 11 2 0 9 2 11 2 11 2 11 2 11 2 3 13 15 0 2 2
10 15 4 3 13 10 2 0 9 2 2
14 15 1 10 0 2 15 2 15 15 13 3 1 11 2
14 1 11 13 15 3 2 1 0 9 2 9 1 9 2
21 15 15 13 1 9 2 3 13 2 3 15 13 3 0 9 2 16 13 15 15 2
20 13 1 15 2 16 9 11 13 3 0 1 0 0 11 7 7 11 16 15 2
1 11
10 9 9 2 7 15 13 2 3 2 3
19 1 9 0 0 9 13 9 1 9 2 15 13 7 3 13 1 15 0 2
21 3 2 3 15 3 13 2 13 9 1 10 0 9 0 2 16 13 1 9 9 2
27 7 14 3 15 2 1 15 7 1 15 2 13 13 2 13 9 2 9 2 16 4 15 13 1 9 9 2
26 3 10 9 15 13 2 13 3 2 16 3 3 2 16 9 15 3 3 13 2 7 3 15 3 0 2
24 3 3 11 1 0 9 13 2 16 9 15 13 10 0 9 2 10 9 1 9 9 13 0 2
18 0 9 15 13 9 2 9 2 13 15 9 2 7 16 10 0 9 2
31 1 9 12 9 13 2 3 1 9 2 15 9 9 2 1 12 7 15 9 3 1 15 13 7 9 2 7 15 15 13 2
13 0 9 1 9 9 2 13 11 2 13 0 12 2
17 7 15 15 3 7 14 13 1 9 0 9 9 0 9 10 9 2
22 7 1 10 0 9 2 0 9 2 2 9 1 0 9 7 0 0 9 1 0 9 2
19 15 15 9 7 3 13 9 12 2 3 15 13 9 7 10 9 1 11 2
44 0 3 9 1 9 13 10 3 0 9 12 2 3 13 9 2 15 3 0 9 13 9 2 1 9 7 1 9 2 0 9 2 14 16 4 1 15 9 15 13 1 0 9 2
18 15 9 0 9 2 15 0 7 0 7 2 3 13 13 2 3 0 2
4 9 13 7 13
24 7 7 0 3 0 9 0 9 15 1 9 0 9 7 15 0 2 15 13 2 13 0 9 2
52 2 13 9 9 2 2 13 12 2 2 9 14 9 2 2 13 0 2 7 0 13 1 9 2 16 9 15 13 2 1 9 9 2 2 15 4 3 13 0 9 2 0 9 2 15 3 3 4 13 9 2 2
85 14 1 12 9 3 10 9 15 13 7 13 7 13 9 2 10 0 0 9 2 2 0 9 0 1 9 15 9 2 2 13 13 9 2 15 13 0 13 2 15 3 13 2 1 0 7 3 14 3 14 0 0 9 2 1 3 0 9 2 1 0 9 9 2 16 4 15 13 14 1 10 0 9 2 15 3 9 1 9 0 13 2 7 13 2
21 1 10 9 15 13 0 2 3 0 16 0 2 9 1 9 2 15 13 9 9 2
26 9 9 13 1 9 9 0 2 7 1 9 0 9 0 2 9 1 1 9 0 0 9 0 0 9 2
30 1 10 9 13 1 9 9 12 9 1 0 9 2 1 9 10 9 2 0 1 12 9 3 0 1 0 9 0 9 2
32 7 13 15 10 9 7 10 9 2 15 1 0 9 13 2 1 10 0 7 0 9 13 9 2 0 9 1 3 0 0 9 2
27 1 9 3 7 3 13 0 2 7 3 3 0 2 9 0 9 1 9 0 7 9 0 9 7 10 9 2
6 1 9 9 13 9 2
8 2 13 4 1 0 0 9 2
34 3 7 3 13 10 9 3 13 2 2 13 0 9 11 11 7 3 13 2 2 3 13 9 2 16 0 9 13 2 7 16 13 2 2
45 9 0 0 9 0 11 13 1 9 9 12 2 2 9 3 13 1 0 2 0 7 0 9 2 16 3 13 13 16 2 9 2 2 16 2 9 2 9 3 0 2 1 9 2 2
36 2 13 4 2 13 15 7 15 3 3 11 2 1 2 0 0 9 2 0 15 9 2 16 9 7 9 13 13 14 0 2 3 0 9 2 2
4 9 9 0 9
25 13 9 2 16 4 13 2 3 15 10 9 0 9 13 2 7 3 13 1 9 7 15 1 15 2
28 13 15 13 10 9 7 9 2 15 15 15 3 3 13 1 12 0 2 0 9 1 9 11 2 3 1 15 2
2 0 2
32 14 1 15 2 16 1 15 9 7 9 15 13 3 3 7 3 2 14 15 4 13 3 7 15 13 3 2 7 15 13 3 2
4 0 2 3 2
5 15 4 13 13 2
6 0 2 7 13 15 2
10 15 1 15 13 2 15 13 15 0 2
6 10 0 2 3 3 2
12 14 16 4 1 15 2 3 1 9 2 13 2
24 7 13 0 9 2 16 13 2 15 13 2 3 1 15 0 7 0 2 16 0 9 0 9 2
10 13 15 3 9 14 0 2 7 0 2
6 1 9 2 15 13 2
9 1 9 2 10 0 9 13 9 2
8 1 0 9 2 15 15 13 2
14 1 0 9 2 16 3 1 15 3 7 3 13 0 2
60 0 9 1 9 13 1 15 0 2 13 15 3 3 12 7 3 3 0 9 0 9 2 2 16 11 2 11 2 7 7 11 13 3 9 7 9 2 9 2 9 0 9 1 11 2 13 1 9 2 13 3 13 9 2 1 2 9 2 2 2
23 3 2 13 15 0 9 2 13 15 0 9 2 7 3 15 13 0 2 3 0 7 0 2
28 9 2 0 7 0 9 0 9 2 9 0 9 2 13 1 15 13 9 9 2 14 7 9 1 0 7 0 2
11 13 15 3 1 9 2 16 4 13 13 2
20 13 15 2 15 13 9 15 2 15 13 2 1 15 13 2 15 15 15 13 2
27 13 15 1 15 15 7 1 15 2 15 13 2 1 0 9 2 15 13 3 0 9 7 4 1 15 13 2
8 3 2 13 15 1 15 13 2
48 1 0 9 2 1 0 9 7 0 9 2 1 0 9 9 2 9 7 0 0 9 2 1 0 9 2 15 15 13 2 0 9 0 15 9 0 9 2 1 0 9 0 9 9 9 2 2 2
56 7 14 16 4 2 3 3 14 1 9 2 10 15 7 0 0 13 16 0 9 0 9 1 15 2 7 3 15 2 0 2 1 9 9 2 1 15 4 4 13 7 1 15 3 15 9 7 9 0 7 14 1 3 0 9 2
21 7 3 15 13 2 16 15 1 10 0 9 4 13 3 2 16 13 1 9 0 2
5 3 3 3 15 2
32 13 15 3 3 0 9 13 1 15 2 16 16 3 2 1 9 2 1 9 2 1 9 2 13 3 3 2 3 13 3 3 2
42 7 3 15 13 13 3 2 7 3 3 1 0 0 9 0 11 7 1 0 11 7 11 2 16 4 15 13 0 9 10 0 0 2 0 2 7 7 0 7 0 9 2
7 13 0 2 7 14 0 2
6 0 2 7 14 0 2
6 13 9 2 14 9 2
8 13 0 2 7 14 1 9 2
10 15 4 15 1 0 9 13 7 13 13
2 11 11
4 7 9 13 9
22 9 0 15 1 9 9 13 9 2 11 9 2 12 2 3 13 9 2 15 13 9 2
20 13 0 9 2 13 1 10 9 3 12 9 7 13 15 13 9 1 0 9 2
16 13 2 16 15 15 13 3 2 3 4 15 13 1 0 9 2
16 10 9 13 7 9 15 2 16 7 2 0 9 13 9 2 2
8 10 3 0 9 13 0 9 2
26 15 13 2 16 4 9 13 9 2 7 2 9 0 7 0 1 0 9 2 7 3 4 15 13 9 2
28 3 15 13 2 16 9 3 13 14 10 9 2 1 15 15 13 7 1 0 9 13 0 2 16 13 9 3 2
16 16 15 3 9 2 15 3 9 2 15 3 9 1 0 9 2
18 13 15 9 2 15 15 13 1 15 9 13 3 7 13 1 15 0 2
22 3 15 15 13 10 0 9 3 13 7 3 15 1 15 13 13 7 9 1 0 9 2
17 13 2 14 15 2 16 13 0 9 13 0 9 2 3 15 13 2
19 3 3 15 13 2 13 2 14 15 2 16 9 1 0 9 13 0 9 2
9 7 3 3 13 0 9 1 9 2
9 15 9 1 0 9 15 13 3 2
25 15 15 13 2 9 13 3 3 2 9 13 0 16 15 0 7 13 2 14 0 2 13 15 15 2
4 15 1 15 2
25 3 4 15 13 13 9 0 9 2 15 4 13 9 13 9 2 15 1 0 9 9 1 9 13 2
72 7 16 1 0 9 0 9 13 3 1 12 2 12 9 2 15 13 13 15 13 1 10 9 2 16 9 15 13 3 9 9 1 0 9 2 1 15 13 1 9 3 12 9 2 1 15 15 13 1 9 0 9 2 7 0 12 7 12 12 9 15 9 13 3 2 16 15 9 13 0 9 2
12 9 9 13 13 10 2 3 0 2 0 9 2
30 3 15 13 7 3 13 2 13 15 1 15 1 9 7 13 0 0 9 2 4 2 14 15 1 15 13 13 12 9 2
26 0 9 13 9 0 0 9 2 3 15 9 15 13 9 1 0 9 2 15 13 1 10 9 3 0 2
16 9 15 13 1 0 9 2 7 13 9 2 15 9 13 9 2
22 3 4 13 9 0 9 9 7 13 2 14 0 2 1 9 13 7 13 4 7 9 2
14 3 3 13 10 0 9 2 3 4 13 0 1 0 2
8 1 9 9 2 11 11 2 0
2 0 11
4 3 13 13 2
9 1 9 2 1 9 2 1 9 2
24 3 14 13 1 9 13 9 2 3 15 7 13 1 15 2 16 4 15 13 13 9 1 9 2
18 7 3 15 13 9 2 15 13 1 9 9 2 13 15 9 2 9 2
15 7 1 9 13 9 1 10 2 9 2 7 0 9 9 2
18 13 9 2 16 1 11 15 9 13 9 2 15 13 1 0 9 0 2
5 3 3 9 13 2
30 3 2 1 3 0 11 2 1 0 0 9 2 15 1 9 13 1 12 2 12 9 2 1 9 1 12 2 12 9 2
17 1 11 13 9 1 9 3 0 2 13 15 1 12 2 12 9 2
32 1 9 2 15 9 1 0 0 9 13 2 15 13 9 1 9 0 9 2 9 1 3 0 9 0 7 0 9 2 3 9 2
25 9 0 9 2 15 3 13 9 1 9 2 15 3 7 13 2 16 13 9 9 7 10 9 13 2
28 16 15 15 13 1 9 9 13 10 0 9 7 15 7 10 9 2 4 3 13 3 3 2 16 13 15 0 2
6 1 9 11 11 2 11
3 15 9 13
6 2 11 9 2 12 2
14 13 15 13 0 9 7 13 1 0 9 9 0 9 2
34 3 9 9 15 13 2 0 9 13 3 1 11 16 1 11 2 7 7 4 9 2 11 7 11 2 3 1 0 9 13 9 0 9 2
11 1 10 9 15 3 1 11 3 3 13 2
19 1 9 9 1 11 4 13 2 16 9 9 9 13 1 9 9 0 11 2
6 14 2 9 13 0 2
20 13 12 9 2 0 13 10 9 2 10 0 9 7 3 10 9 7 10 9 2
14 9 9 13 2 16 9 0 9 13 3 1 9 11 2
27 13 15 7 16 9 0 9 2 16 4 13 9 0 9 13 0 9 1 0 9 7 15 13 9 0 9 2
16 10 9 13 15 0 1 9 2 16 15 9 11 13 7 3 2
7 1 9 11 2 11 2 11
3 9 1 9
20 13 0 9 2 0 9 7 9 0 9 7 9 15 3 13 1 10 0 9 2
5 15 15 13 3 2
24 9 4 13 1 0 9 7 9 15 13 3 2 3 2 16 16 1 9 13 2 13 1 9 2
23 9 3 13 1 0 9 2 0 9 13 0 9 2 0 0 9 15 13 1 9 1 9 2
5 7 13 15 3 2
19 9 3 13 13 2 3 15 13 9 1 0 9 2 3 15 13 1 9 2
6 3 13 3 1 9 2
25 3 15 12 9 13 0 0 9 1 9 7 11 13 1 10 0 9 1 9 7 13 1 0 11 2
27 15 13 2 12 0 9 13 1 9 0 3 2 16 4 0 1 15 13 3 10 9 1 0 9 3 11 2
8 3 15 13 2 13 7 13 2
16 0 9 2 9 11 7 9 11 13 9 7 13 7 1 9 2
5 3 2 13 9 2
5 9 15 9 13 2
4 3 7 3 2
6 16 10 0 0 9 2
4 11 9 2 11
16 2 2 2 14 2 16 4 13 9 14 16 13 0 2 2 2
3 9 11 11
3 9 1 9
21 0 9 1 9 2 10 0 9 16 0 9 2 0 9 1 9 0 1 0 9 2
74 7 9 9 1 0 0 9 2 9 2 15 10 9 13 7 15 4 15 1 15 3 13 2 2 9 1 9 0 1 0 9 15 0 1 9 9 2 16 9 15 13 1 0 9 1 9 7 9 1 9 13 9 9 1 2 9 2 7 9 1 0 1 0 9 2 2 2 13 4 15 3 3 13 2
12 0 13 2 16 1 15 13 2 16 15 13 2
13 13 10 9 2 16 1 0 9 13 1 0 9 2
22 13 4 1 15 13 1 0 9 13 2 13 7 3 15 0 13 1 10 0 0 9 2
4 11 11 2 11
3 13 15 9
6 2 11 9 2 12 2
39 9 2 16 12 9 13 3 0 9 2 15 13 14 3 2 16 4 15 13 0 9 2 7 16 15 13 2 16 9 1 11 4 15 13 15 13 9 0 2
39 13 2 14 3 9 2 1 10 0 9 9 13 2 13 4 15 15 13 1 15 0 2 6 2 9 0 2 15 10 9 2 2 7 1 10 0 9 2 2
12 3 1 9 2 16 9 13 0 9 10 9 2
31 16 2 9 13 9 2 3 9 1 10 9 2 7 9 13 1 10 9 3 0 9 2 15 13 9 1 10 9 3 13 2
11 3 13 2 13 0 7 9 0 0 9 2
7 9 13 13 9 2 6 2
7 9 9 1 15 15 13 2
16 13 15 13 9 11 7 0 0 9 2 10 9 10 9 13 2
35 13 2 14 15 3 2 3 1 0 9 13 13 2 16 1 0 9 13 15 2 15 2 13 1 15 1 15 9 2 4 3 13 10 9 2
21 13 13 2 16 0 9 1 0 9 4 15 10 9 1 2 0 2 9 13 13 2
32 0 1 15 13 2 16 15 1 9 0 2 0 7 0 9 3 13 1 15 2 1 15 3 13 2 1 9 0 9 0 9 2
7 1 9 11 11 2 11 11
2 15 13
6 2 11 9 2 12 2
28 1 0 9 1 9 0 9 0 2 9 4 13 9 2 16 0 9 0 9 10 9 13 9 9 11 7 11 2
15 2 0 9 11 7 11 14 13 2 7 7 3 13 2 2
22 15 7 10 2 0 9 2 13 10 9 1 9 2 15 3 15 9 1 9 3 13 2
28 9 9 11 11 2 11 3 13 10 9 1 9 0 2 7 3 9 9 11 7 11 9 11 10 9 3 13 2
23 13 2 16 0 9 10 9 13 3 0 2 16 9 0 3 1 0 11 7 3 1 9 2
49 1 9 9 2 16 15 13 3 1 0 0 9 2 13 0 9 2 9 0 9 11 1 9 7 1 9 2 16 9 10 9 13 3 0 1 0 9 7 10 0 9 13 9 0 9 1 15 9 2
15 13 2 16 0 9 13 9 0 7 9 11 7 11 0 2
4 11 11 2 11
3 9 16 9
8 2 11 9 2 12 2 12 2
32 9 3 13 10 0 9 9 0 9 2 15 1 10 9 13 9 9 1 9 2 15 1 10 9 13 14 0 9 10 0 9 2
15 13 15 15 2 16 14 1 10 0 9 13 13 0 9 2
21 3 3 2 16 9 13 13 1 9 0 9 2 15 13 3 13 1 0 0 9 2
28 3 13 0 13 2 16 1 12 9 1 9 12 1 15 13 13 0 9 7 1 9 2 7 1 9 0 9 2
19 3 3 15 3 3 4 13 0 9 9 0 9 2 9 7 9 0 9 2
54 3 15 13 2 16 0 9 9 13 3 13 9 10 0 9 2 15 1 9 1 3 0 9 2 13 10 9 0 9 1 10 9 2 16 1 9 1 9 13 13 1 9 0 2 3 2 3 1 15 9 13 1 9 2
4 11 11 2 11
26 9 7 9 15 3 13 0 9 2 16 4 15 13 7 13 13 3 7 3 3 2 16 1 15 13 2
5 11 11 2 0 11
1 0
30 1 9 9 11 11 13 12 9 2 15 4 15 1 15 13 13 3 9 10 0 9 2 9 10 12 9 7 0 9 2
21 13 15 2 0 2 7 16 13 13 1 12 2 9 2 13 3 16 0 7 3 2
10 2 14 12 9 15 13 2 0 2 2
4 9 7 9 2
8 0 9 15 13 14 1 9 2
4 0 9 3 2
14 3 9 13 9 2 16 4 1 15 13 10 0 9 2
16 13 2 14 15 9 3 3 2 13 15 1 0 9 1 9 2
12 13 2 14 9 9 2 13 15 1 0 9 2
11 10 9 13 0 7 13 1 15 3 9 2
7 3 15 15 13 1 9 2
8 9 13 10 0 9 0 9 2
5 13 13 0 9 2
14 13 3 11 12 13 11 12 7 13 15 1 9 13 2
24 13 0 9 13 0 9 7 13 2 16 4 15 13 9 2 16 15 13 9 9 7 0 9 2
18 13 13 0 9 1 11 7 11 2 3 15 13 0 9 1 0 9 2
18 7 13 2 14 15 3 0 9 0 9 2 13 1 15 7 9 9 2
23 14 9 15 13 2 7 0 0 2 3 0 2 7 3 0 2 9 14 13 2 7 13 2
18 3 15 13 3 0 9 2 7 14 3 2 16 4 15 13 13 3 2
20 3 15 3 3 13 0 9 2 16 4 15 13 13 7 13 1 10 0 9 2
12 13 0 13 9 2 13 2 14 3 9 9 2
13 13 0 13 0 9 2 4 2 14 3 13 9 2
22 13 2 14 1 15 2 13 9 10 9 2 10 9 2 10 9 15 3 16 9 2 2
1 13
4 11 9 2 11
25 1 9 13 1 11 3 3 2 1 0 11 7 1 11 3 3 7 9 3 3 14 0 0 9 2
37 0 9 12 7 12 9 2 9 2 2 1 12 9 3 1 9 2 0 9 1 11 12 7 12 9 2 9 2 1 11 12 7 12 9 2 9 2
17 1 9 7 1 9 13 1 11 3 9 9 2 1 9 9 3 2
12 1 9 1 9 9 14 3 7 3 0 9 2
14 0 0 9 12 7 9 12 2 1 0 9 7 0 2
19 0 9 1 9 1 9 12 7 12 2 1 9 12 7 12 9 2 9 2
25 1 0 9 13 1 9 3 2 1 9 7 9 1 9 9 3 2 9 0 9 2 3 1 9 2
28 0 9 12 7 12 9 2 9 2 1 0 9 12 7 12 9 2 9 2 0 0 12 7 12 9 2 9 2
24 0 9 12 7 12 9 2 9 2 1 9 12 7 12 9 2 9 2 1 0 0 9 9 2
11 9 9 1 9 12 9 12 9 2 9 2
29 1 9 7 1 9 13 1 11 9 7 3 2 3 1 9 9 2 1 9 1 9 7 9 9 3 7 9 9 2
36 0 9 12 7 12 9 2 9 2 1 0 9 1 12 9 2 9 2 0 9 12 7 12 9 2 9 2 1 9 12 7 12 9 2 9 2
3 9 1 9
29 3 1 0 9 13 13 1 10 9 9 7 9 2 9 2 0 9 7 9 2 7 15 1 12 3 15 0 9 2
34 1 0 9 9 15 13 9 9 1 9 2 15 13 0 9 1 0 9 2 1 0 9 1 9 14 1 0 9 7 0 9 1 0 2
9 9 10 9 13 3 10 0 9 2
24 13 9 3 1 0 9 2 3 9 7 13 3 0 9 1 9 7 9 2 3 9 0 9 2
33 0 9 2 9 1 9 2 13 9 0 0 9 0 9 2 1 3 0 9 0 0 9 1 0 9 2 14 1 0 9 7 9 2
14 1 12 9 15 13 3 1 9 9 2 3 9 9 2
33 7 1 10 0 3 13 9 7 9 10 9 2 16 1 9 1 0 0 9 3 1 15 13 9 2 15 2 3 7 3 15 13 2
19 0 13 14 9 2 15 15 13 2 7 0 13 10 9 2 3 7 3 2
37 13 15 3 0 9 15 0 9 2 15 13 1 9 9 3 0 9 2 3 9 1 9 2 0 9 2 0 9 2 3 0 9 7 0 0 9 2
3 13 13 2
5 0 9 1 9 9
12 1 0 9 13 1 10 9 0 9 9 9 2
14 3 0 2 3 1 15 0 2 7 3 1 0 9 2
15 1 9 0 9 7 9 4 13 9 9 2 9 7 9 2
9 15 9 13 1 9 9 1 9 2
10 3 1 9 13 1 0 9 9 9 2
7 13 1 9 10 0 9 2
8 1 9 9 13 7 0 9 2
8 13 9 2 15 13 15 13 2
27 10 9 1 9 13 9 9 1 9 7 9 2 10 9 13 0 9 0 9 0 3 1 9 7 1 9 2
23 13 1 9 7 3 3 13 13 1 15 2 16 13 15 3 2 7 9 1 10 9 13 2
13 13 0 13 0 1 9 0 9 0 0 12 9 2
7 13 0 13 13 7 13 2
27 13 13 14 10 0 2 15 0 9 7 13 3 0 9 2 15 0 9 0 9 13 3 1 9 1 9 2
21 15 1 10 9 13 9 1 9 9 0 1 9 15 0 0 7 0 9 0 9 2
11 15 4 13 9 2 13 9 2 13 9 2
11 13 9 7 9 2 15 13 7 13 13 2
8 13 9 2 15 13 0 13 2
33 1 12 9 10 9 13 0 9 0 0 7 3 0 9 1 9 2 3 3 3 15 9 0 13 0 0 9 7 13 15 0 9 2
8 1 9 15 7 1 9 15 2
8 14 9 9 13 1 9 9 2
10 1 15 13 0 9 9 1 0 9 2
13 9 13 0 14 9 9 2 7 7 10 0 9 2
40 13 4 7 15 15 2 15 4 3 13 2 13 2 2 2 13 0 2 7 15 3 14 13 7 0 9 2 13 2 16 1 10 9 13 0 13 3 16 9 2
11 1 15 15 13 3 3 13 16 0 9 2
12 9 2 15 3 13 7 13 9 12 1 0 2
11 9 0 10 9 13 13 7 13 0 15 2
4 9 2 11 11
7 11 1 0 9 1 0 9
5 11 13 2 11 2
2 11 2
38 0 9 9 11 2 0 9 2 0 12 9 1 9 1 9 11 2 3 3 1 9 11 2 13 11 11 11 1 9 11 7 13 3 1 9 0 9 2
17 1 9 13 0 11 11 2 1 0 9 11 11 15 7 15 13 2
22 3 15 13 10 9 2 11 1 11 13 1 0 9 2 3 0 2 2 11 13 0 2
12 11 13 0 9 1 11 12 9 7 12 9 2
9 7 1 9 9 10 9 1 0 11
5 0 9 1 9 2
9 11 11 13 1 9 3 12 9 2
13 13 7 3 0 9 1 11 11 7 13 15 15 2
12 1 9 3 9 13 1 11 11 12 2 12 2
10 11 1 9 9 13 9 1 0 9 2
24 1 9 9 1 11 13 3 1 0 9 1 0 9 7 13 12 9 1 12 9 7 12 9 2
18 1 15 13 12 0 9 11 11 7 11 2 3 11 2 11 7 11 2
16 11 13 15 12 9 9 7 13 3 0 9 2 9 12 9 2
8 13 15 2 16 7 3 13 2
33 1 11 13 3 0 0 9 9 2 15 13 7 15 2 16 4 3 3 13 1 9 15 11 1 9 0 9 1 9 0 9 11 2
19 11 11 1 0 9 13 2 2 13 15 3 7 13 15 2 16 13 9 2
12 13 4 0 9 11 2 16 4 15 15 13 2
3 7 3 2
7 9 15 13 7 9 13 2
18 13 3 7 1 9 11 2 16 13 3 9 9 13 1 9 1 9 2
5 13 3 9 2 2
26 11 9 2 15 13 1 12 9 0 16 10 9 1 9 2 13 2 2 13 4 3 0 9 1 9 2
9 1 11 13 3 1 9 3 3 2
12 13 2 16 13 0 0 12 9 1 10 9 2
11 1 15 13 3 9 2 7 3 15 13 2
10 12 9 1 9 2 14 13 0 9 2
16 7 0 13 2 16 4 9 13 0 7 13 4 15 3 3 2
17 13 3 3 0 9 2 11 13 1 0 9 9 9 2 15 13 2
8 13 3 7 3 15 15 13 2
8 1 0 9 11 11 13 9 2
11 13 15 3 1 9 0 9 1 9 11 2
7 13 3 0 16 11 11 2
11 0 9 13 7 0 2 7 10 9 9 2
29 15 13 0 2 15 13 3 1 11 13 11 9 7 11 11 2 7 15 13 1 9 2 3 15 3 15 13 2 2
18 9 0 9 11 13 7 11 1 11 2 15 13 1 0 15 12 9 2
22 7 15 7 13 2 16 11 13 3 7 13 3 0 9 12 0 9 11 1 0 9 2
20 1 9 11 1 0 11 13 3 12 9 1 9 2 12 1 15 13 11 11 2
21 9 11 2 11 13 3 9 9 11 11 7 11 11 2 1 15 13 3 0 11 2
16 1 9 11 13 10 0 9 9 11 11 2 0 9 0 11 2
28 3 1 9 13 0 9 2 13 1 11 1 9 9 2 15 15 1 9 13 1 0 9 1 3 12 9 11 2
25 11 11 2 9 9 11 11 11 11 2 15 7 13 2 16 4 10 9 13 1 9 9 0 9 2
29 2 1 10 9 10 9 13 2 7 3 15 13 2 2 13 11 2 2 16 1 9 13 9 2 1 15 13 9 2
8 9 9 13 9 3 3 13 2
8 13 15 1 0 9 1 9 2
11 3 3 13 13 9 9 7 10 9 2 2
20 15 11 11 13 10 9 1 10 9 7 13 9 1 9 9 11 9 11 11 2
6 15 15 7 13 3 2
23 2 1 15 15 0 9 3 13 7 2 9 9 2 15 3 2 7 3 2 13 9 2 2
31 13 1 9 2 16 9 13 3 11 2 1 11 11 12 2 11 2 11 2 11 2 11 7 11 2 1 11 11 7 11 2
7 0 0 2 9 13 11 2
3 9 13 9
2 11 2
28 9 1 0 9 10 0 9 1 9 9 9 1 12 9 2 0 0 9 1 0 11 2 13 1 9 3 11 2
8 10 9 13 0 9 7 13 2
3 3 3 2
6 11 2 11 12 2 12
11 3 1 9 9 13 0 2 9 0 9 2
41 1 0 9 3 3 1 0 9 13 11 7 3 11 2 7 9 13 7 12 0 2 9 2 1 15 12 2 1 12 2 9 2 2 12 2 12 13 12 2 12 2
16 0 2 9 15 1 10 0 2 0 9 13 7 12 0 9 2
19 1 9 12 1 0 9 13 11 9 2 15 1 0 2 9 3 15 13 2
21 7 1 9 0 9 9 13 3 0 2 9 9 1 9 2 7 15 1 15 13 2
31 1 12 2 9 2 13 0 9 11 9 1 9 11 1 9 2 7 9 13 7 12 1 0 9 15 13 2 12 2 12 2
26 3 1 10 9 15 13 0 2 9 2 7 15 13 9 9 2 7 16 9 13 0 12 9 3 3 2
14 9 13 3 3 9 2 15 15 13 1 9 7 9 2
19 9 11 7 11 3 13 15 13 2 7 0 9 13 3 3 3 1 9 2
25 3 3 1 11 9 1 12 9 13 0 9 3 1 0 2 9 7 0 2 9 13 3 1 9 2
16 0 9 1 12 2 9 2 13 14 9 1 9 0 2 9 2
13 2 2 1 11 11 2 0 9 0 2 9 2 9
25 1 0 12 9 0 9 1 11 15 1 0 9 9 9 1 11 13 1 9 7 12 0 11 11 2
6 15 13 9 10 9 2
15 2 11 13 9 2 15 13 3 1 9 9 9 11 11 2
22 0 9 1 0 9 1 0 0 0 9 1 11 13 0 9 1 0 9 1 11 2 2
11 13 11 9 13 7 1 0 9 1 11 2
29 2 16 15 13 1 11 1 9 1 12 9 3 1 12 2 9 2 3 4 13 7 1 0 9 9 1 0 11 2
11 3 1 10 9 13 9 9 1 0 9 2
38 11 1 10 9 13 2 15 13 2 16 16 4 13 3 3 1 11 2 3 10 9 1 0 9 13 1 0 9 9 7 4 15 3 13 0 9 2 2
13 10 9 13 9 0 2 9 2 15 13 1 11 2
40 2 3 1 0 9 13 9 2 11 2 11 7 11 3 1 9 11 1 0 11 2 3 4 13 1 0 9 0 1 15 2 1 15 13 0 9 1 0 11 2
15 10 9 15 13 3 1 11 1 11 1 0 9 0 9 2
11 0 0 9 1 9 13 13 1 11 2 2
8 0 9 15 13 1 11 2 11
3 9 0 9
20 9 13 2 2 2 2 2 2 2 2 2 2 2 2 2 2 2 2 2 2
4 11 2 11 2
40 0 9 15 1 9 3 13 1 11 1 0 9 0 11 1 11 2 11 2 3 4 9 13 1 0 9 1 0 9 9 7 3 7 1 0 9 1 0 9 2
25 9 13 13 0 9 2 9 9 4 13 14 3 2 3 3 2 16 1 11 2 11 13 0 9 2
28 16 0 7 0 11 13 3 9 0 9 0 9 2 3 0 7 3 0 11 2 11 13 0 9 0 12 12 2
15 7 3 3 7 13 1 10 9 9 3 12 0 0 9 2
32 9 1 9 15 3 13 9 1 10 0 0 0 11 2 15 3 1 9 3 13 15 13 2 7 1 0 9 13 15 0 9 2
15 1 9 3 4 3 13 12 0 9 2 15 13 0 9 2
19 9 1 10 9 13 12 0 9 1 9 1 11 2 11 2 11 7 11 2
17 13 15 4 1 0 9 1 0 9 2 10 9 13 3 12 9 2
42 0 9 13 13 1 12 0 9 2 1 15 3 12 1 0 9 13 1 9 2 12 0 3 1 9 7 12 0 15 3 13 1 9 1 12 9 2 16 0 13 9 2
22 13 15 7 1 0 9 2 0 9 12 7 1 2 0 2 9 13 9 1 9 12 2
11 0 9 13 12 7 0 1 0 9 12 2
24 0 9 0 9 11 11 15 1 10 9 3 13 2 2 13 15 0 9 1 9 1 0 9 2
15 16 13 0 9 13 2 13 3 3 13 0 9 9 2 2
11 13 9 2 3 13 11 11 1 9 3 15
10 2 2 2 7 3 4 13 10 9 2
4 16 13 9 2
15 3 4 15 13 9 2 9 13 1 15 9 2 15 13 2
12 13 7 2 16 15 10 9 13 13 1 9 2
10 7 15 3 3 2 16 15 3 13 2
8 15 3 13 14 12 1 9 2
10 3 4 15 15 13 1 9 1 11 2
6 13 4 3 15 9 2
18 3 3 4 3 13 1 9 1 11 7 15 13 1 9 1 0 9 2
10 13 4 3 3 7 13 3 1 9 2
17 7 16 4 15 13 1 9 2 3 4 13 10 9 2 2 2 2
53 9 10 3 0 9 13 11 11 2 12 0 0 9 1 11 2 0 0 9 10 0 9 2 15 15 1 0 13 13 9 2 0 2 9 9 1 0 9 7 12 0 9 1 11 2 15 13 3 0 0 9 9 2
15 1 12 9 13 0 2 3 13 7 3 13 1 0 9 2
31 3 15 15 1 0 9 3 13 2 16 1 9 13 0 12 9 2 15 13 3 1 0 9 9 12 9 1 9 1 11 2
27 2 11 13 1 0 9 9 1 0 0 9 2 3 0 16 13 3 0 9 7 9 2 2 13 11 11 2
18 2 9 3 13 13 12 0 9 2 16 4 15 13 1 10 0 9 2
13 15 13 0 3 7 1 0 9 13 15 3 0 2
27 3 4 3 13 1 0 9 1 11 14 0 7 15 13 0 9 14 1 0 9 2 7 7 1 10 9 2
19 3 4 15 15 13 7 13 1 15 2 16 3 3 15 13 13 0 9 2
18 16 4 3 13 1 11 2 11 0 2 13 4 2 16 9 3 13 2
8 7 3 13 15 3 3 2 2
8 10 9 13 9 13 3 0 2
18 10 9 11 7 3 13 2 2 15 2 13 0 9 2 15 13 9 2
22 2 9 14 13 13 1 9 2 15 13 2 7 10 9 13 13 14 0 2 7 0 2
18 7 15 1 10 9 2 16 0 9 13 12 9 2 15 13 1 9 2
34 2 16 13 2 3 9 13 10 9 2 13 3 1 9 9 9 2 2 13 15 11 2 2 7 16 13 15 3 3 12 2 15 13 2
16 16 13 2 7 13 2 3 15 3 16 3 13 13 1 9 2
7 7 3 3 13 1 15 2
12 0 12 9 1 9 13 1 9 3 15 2 2
22 11 2 3 2 13 1 0 9 0 9 7 1 2 9 2 2 9 13 3 1 9 2
24 13 15 15 3 2 16 15 9 13 1 9 7 9 1 9 13 1 9 1 0 9 3 0 2
22 11 15 13 1 9 2 7 9 1 15 3 13 15 2 15 2 9 2 13 1 9 2
13 2 1 9 11 13 15 9 2 15 3 15 13 2
27 13 15 0 2 3 15 3 13 7 13 15 13 2 16 15 13 15 0 13 2 3 10 9 13 1 9 2
6 16 1 15 13 9 2
7 9 2 2 13 3 11 2
9 2 15 13 9 2 7 9 9 2
12 7 7 1 0 9 15 9 1 9 13 13 2
20 1 9 3 13 12 9 2 9 7 9 2 1 9 15 13 7 13 2 2 2
17 7 1 9 3 3 13 9 0 9 7 2 9 2 0 9 2 2
5 13 3 1 9 2
3 2 14 2
18 16 9 4 3 13 13 1 0 9 0 9 0 9 16 11 7 11 2
15 9 13 1 11 2 11 2 11 7 3 3 1 11 2 2
4 11 11 2 11
17 11 11 0 9 11 11 1 9 0 9 1 9 11 2 0 9 2
18 7 10 9 9 15 7 13 9 0 9 2 3 12 13 3 0 9 2
3 3 1 9
18 1 9 0 9 0 9 1 11 13 9 1 11 0 9 12 2 12 2
29 2 13 4 3 0 1 0 9 7 13 4 9 9 7 0 9 13 2 16 13 3 2 2 13 1 9 11 9 2
13 2 1 10 9 13 3 0 13 13 12 1 0 2
15 13 2 16 4 13 0 9 1 9 2 2 13 11 11 2
3 11 1 9
28 9 11 7 11 13 2 0 11 2 2 9 1 0 9 9 2 15 1 9 9 9 13 0 9 11 0 9 2
2 9 9
25 12 0 7 12 0 2 15 13 0 9 9 2 1 15 13 1 9 9 1 0 11 1 9 11 2
23 10 9 1 10 9 13 3 1 9 7 3 13 12 9 10 9 2 15 13 1 0 9 2
11 3 13 1 9 1 9 7 0 9 9 2
21 1 0 9 15 13 13 3 0 9 2 12 0 1 9 9 13 7 0 15 13 2
25 12 9 10 9 13 0 9 2 3 1 9 4 3 13 1 0 9 2 16 13 0 9 2 2 2
2 0 11
22 9 11 9 11 11 3 1 0 9 13 0 9 1 9 2 16 12 9 13 0 9 2
18 1 9 13 10 9 1 0 11 12 2 12 2 16 13 0 12 9 2
36 1 0 9 13 1 9 7 11 9 2 15 13 7 13 2 2 1 0 9 1 11 15 13 0 9 2 3 13 0 2 1 12 9 3 0 2
3 3 3 2
15 13 3 16 11 11 12 9 2 7 15 13 1 9 3 2
20 2 11 13 1 10 9 12 2 12 1 11 2 10 0 9 13 0 9 11 2
13 13 7 10 9 9 2 15 13 1 9 0 9 2
5 2 11 2 11 2
4 0 9 2 2
81 0 9 0 7 0 9 0 9 1 9 11 2 11 7 11 13 1 10 9 9 12 2 12 2 12 2 16 9 9 11 9 2 0 9 12 2 12 2 12 1 11 11 11 2 7 9 11 11 2 0 12 2 12 2 12 1 11 11 11 2 13 13 1 0 0 2 9 2 13 15 0 9 7 0 9 13 12 9 0 9 2
1 9
1 9
25 0 9 2 12 2 9 0 0 9 0 9 11 15 13 1 11 1 0 9 12 2 9 1 12 2
14 0 9 4 1 0 9 1 12 13 1 9 1 11 2
29 9 13 9 9 0 0 9 2 9 7 0 9 16 9 9 1 9 0 9 2 10 13 0 7 0 9 0 9 2
3 9 2 9
18 9 11 11 11 15 1 9 0 9 13 3 1 12 9 1 0 9 2
14 0 9 0 9 15 3 13 3 13 1 0 9 9 2
1 9
10 0 9 9 1 0 9 11 2 11 2
1 9
31 9 9 9 2 15 15 13 13 1 0 9 1 0 2 9 7 13 1 0 9 2 15 13 12 2 9 1 11 2 11 2
23 4 15 13 1 9 1 9 2 15 15 4 13 12 2 9 1 11 2 11 1 9 11 2
1 9
2 11 2
1 9
11 11 2 11 3 2 1 9 1 11 11 2
14 1 12 2 0 9 15 12 9 13 9 3 1 12 2
1 9
2 0 9
3 1 0 9
2 1 11
1 9
9 0 0 9 13 1 9 1 11 2
23 1 12 2 9 13 9 3 0 0 7 0 9 3 1 0 1 0 9 1 3 0 9 2
3 9 2 9
20 9 11 11 13 9 1 0 9 9 2 11 2 2 0 0 9 11 0 9 2
10 1 9 13 11 7 1 9 9 11 2
1 9
23 0 9 2 9 9 1 0 9 1 11 2 15 13 3 3 1 12 2 9 12 1 11 2
2 0 9
2 11 2
22 3 12 9 7 14 12 9 15 13 9 9 1 0 9 1 0 0 0 9 1 11 2
22 1 9 9 9 1 9 14 9 9 13 13 1 9 0 1 0 9 1 10 0 9 2
13 9 1 9 13 0 2 1 15 10 9 7 9 2
20 1 0 9 2 15 0 9 3 13 7 13 3 12 9 2 15 3 15 13 2
32 9 9 13 9 11 1 0 11 2 3 13 3 9 0 0 9 11 2 15 15 13 1 0 9 1 9 1 9 9 1 11 2
12 3 9 9 13 9 9 0 9 7 0 9 2
12 0 0 9 13 1 15 1 9 9 9 0 2
16 13 14 9 9 7 0 9 1 11 2 7 7 0 9 9 2
5 9 11 11 2 11
12 1 12 2 9 9 15 1 2 0 2 13 2
12 11 2 11 2 11 13 2 7 15 13 2 12
13 11 2 11 2 12 2 9 9 13 1 15 2 12
8 11 2 11 2 9 9 2 12
9 11 2 11 2 0 9 9 2 12
6 15 13 9 12 2 12
9 11 2 11 2 0 13 9 2 12
11 11 2 11 2 11 0 2 9 13 2 12
11 11 2 11 2 1 9 9 0 9 2 12
7 10 9 1 9 12 2 12
14 11 2 11 2 13 15 13 0 2 9 11 9 2 12
3 1 0 9
6 0 2 9 1 11 2
2 11 2
23 12 9 11 2 12 7 0 0 9 1 11 0 1 11 4 1 9 13 1 0 9 11 2
8 13 15 3 0 9 11 0 2
20 9 3 13 2 16 0 2 9 4 9 9 13 1 0 9 1 0 9 11 2
11 13 15 14 1 0 1 9 0 0 9 2
30 1 9 0 2 13 11 11 1 0 9 2 2 15 9 3 13 1 0 9 11 2 15 3 13 0 2 9 0 9 2
31 1 9 9 9 1 9 9 1 0 9 11 11 2 11 9 9 1 0 9 13 9 1 9 9 0 0 9 1 10 9 2
3 0 0 9
12 10 0 0 9 13 1 9 13 15 1 15 2
14 3 16 10 9 9 1 11 13 3 13 9 1 9 2
17 3 4 15 1 10 9 13 13 14 1 0 9 1 9 2 13 2
39 1 1 0 9 1 15 2 16 1 0 0 9 4 13 0 12 9 0 9 7 1 0 9 13 2 13 4 15 15 13 14 1 9 0 9 1 9 9 2
9 9 9 4 3 13 3 0 9 2
11 7 3 15 13 0 7 13 0 15 13 2
8 13 4 3 13 3 7 13 2
6 13 15 3 10 9 2
8 12 2 0 9 0 9 1 9
9 12 2 9 0 9 9 1 0 9
20 12 2 9 0 9 9 11 11 9 11 2 15 15 15 13 7 9 11 13 2
9 13 15 13 9 9 10 0 9 2
18 7 2 12 2 9 15 1 9 0 0 9 13 0 9 7 13 9 2
28 3 15 13 1 0 9 11 7 11 2 2 16 15 12 9 1 9 13 2 9 15 1 9 13 2 2 2 2
22 9 2 12 2 9 15 1 9 13 0 9 7 9 9 1 9 1 9 13 9 1 9
14 9 2 11 11 13 0 0 9 11 1 0 9 9 2
19 9 9 15 7 13 13 0 9 0 2 0 9 2 7 13 15 0 9 2
13 13 15 3 9 7 13 15 9 12 0 11 11 2
9 13 7 13 2 16 10 9 13 2
12 13 15 15 1 0 9 12 9 13 0 9 2
16 3 9 2 16 9 13 13 3 12 2 13 1 0 9 9 2
14 12 9 7 12 9 4 13 3 11 11 1 0 9 2
13 9 2 15 1 15 13 2 13 13 3 3 12 2
18 7 6 2 13 2 14 3 9 12 2 13 15 13 3 11 7 11 2
2 11 11
7 0 9 12 9 0 9 2
3 12 2 9
3 15 13 9
7 2 9 9 13 9 11 2
6 13 15 0 9 2 2
19 10 12 9 13 1 0 9 2 3 1 12 9 2 9 12 0 9 9 2
21 9 13 2 16 9 13 13 1 12 9 7 13 9 13 3 12 0 9 1 15 2
43 0 9 1 9 7 13 2 16 10 9 15 4 13 14 9 0 1 0 9 2 3 0 9 9 2 15 4 13 1 0 0 9 1 9 12 7 1 12 9 1 9 12 2
23 2 13 15 2 16 10 9 13 2 15 4 9 0 13 1 9 9 7 1 0 9 2 2
19 1 9 9 13 1 0 9 0 9 9 2 1 0 0 9 0 9 9 2
42 16 4 7 0 9 13 1 9 2 13 15 0 2 7 1 0 9 7 0 9 9 2 7 3 1 9 1 0 0 9 2 7 3 1 9 9 0 9 9 12 9 2
34 3 13 1 9 13 9 0 9 2 7 15 14 1 0 0 9 2 7 7 1 9 1 0 9 7 1 9 7 9 0 9 7 9 2
16 3 16 9 15 9 13 3 13 3 0 2 0 7 0 9 2
22 16 13 1 0 9 9 2 13 15 1 12 2 9 13 9 9 7 9 13 0 9 2
25 2 15 13 2 3 4 15 13 1 0 9 2 16 4 9 13 9 0 9 3 3 2 2 2 2
48 13 0 9 13 9 3 2 13 2 14 3 16 12 9 0 2 3 16 9 11 13 13 1 0 9 2 16 13 13 9 2 13 15 1 15 2 16 0 9 9 13 13 12 9 1 9 2 2
29 13 9 7 13 0 9 13 9 1 9 2 16 15 13 1 12 9 1 9 9 9 13 9 2 15 13 9 9 2
10 1 15 2 9 2 7 9 9 13 2
25 13 2 14 3 1 9 1 10 0 9 2 13 9 0 9 1 10 0 9 9 2 1 0 9 2
17 1 9 4 3 13 9 7 13 4 1 9 7 9 0 0 9 2
29 0 0 9 15 13 1 9 0 9 3 13 1 0 2 1 9 9 2 7 9 0 9 13 9 13 0 0 9 2
24 7 7 15 3 3 13 0 9 2 7 3 13 1 9 3 3 1 0 9 13 9 0 9 2
3 2 11 2
6 13 9 9 13 9 2
3 9 0 9
18 2 9 9 7 10 0 9 13 0 13 15 2 3 13 1 9 2 2
3 11 2 11
27 16 0 9 13 3 1 9 0 9 7 9 12 0 9 9 2 9 9 7 0 9 0 9 13 0 9 2
35 9 13 1 0 9 1 0 9 9 7 9 9 2 3 0 9 1 9 9 2 9 1 9 9 2 9 0 9 0 11 9 2 9 9 2
46 2 15 13 9 2 16 4 1 0 9 1 0 9 13 7 1 10 9 1 0 12 9 13 2 4 13 9 9 14 1 12 9 7 9 9 7 0 9 2 2 13 15 1 0 9 2
47 1 0 9 15 13 2 2 9 9 14 1 12 9 4 9 13 2 13 2 14 9 1 9 12 7 12 2 9 2 9 2 2 13 1 9 3 2 9 2 3 7 1 9 3 0 2 2
33 0 9 11 9 13 9 3 1 9 9 9 2 1 15 15 1 0 13 2 2 2 2 2 13 1 0 9 0 9 1 0 9 2
47 4 15 0 10 0 9 7 0 0 9 2 1 0 9 3 9 9 0 9 7 3 16 12 9 9 1 9 2 15 10 9 13 2 11 2 0 2 11 2 11 2 11 11 7 0 2 2
22 13 15 1 9 2 1 15 13 13 13 14 15 2 15 13 9 3 7 1 3 9 2
20 1 0 9 4 13 9 13 3 1 0 9 2 16 1 9 0 0 9 2 2
54 9 9 13 9 10 9 9 12 2 1 15 15 1 0 13 2 2 15 15 13 0 7 0 9 9 2 15 13 10 9 7 0 9 15 9 2 4 13 9 9 14 1 12 9 7 0 9 1 12 9 7 0 2 2
38 2 10 9 13 1 9 0 0 9 2 16 2 9 0 9 2 2 2 13 11 11 2 15 13 1 9 1 15 2 15 13 1 9 9 1 9 9 2
35 2 3 13 9 2 16 9 13 2 9 1 0 9 2 7 2 9 1 0 9 2 2 1 15 3 13 2 16 15 1 15 13 13 9 2
9 0 9 4 3 13 9 16 9 2
26 0 9 15 3 13 9 0 9 2 9 2 0 9 1 0 9 7 7 15 2 15 9 13 1 9 2
31 16 1 15 0 9 15 13 9 0 9 2 1 15 9 13 3 1 9 0 2 13 15 3 1 9 2 15 13 9 9 2
31 11 11 3 13 9 1 11 2 3 10 9 13 1 9 0 9 2 7 16 4 3 9 13 2 4 9 13 1 12 9 2
10 1 15 4 1 0 9 13 0 2 2
9 9 9 9 3 9 0 9 13 2
11 11 13 1 0 9 13 9 1 9 9 2
2 11 11
2 9 9
5 11 2 11 2 2
19 1 0 9 9 9 0 9 13 13 0 9 1 9 0 9 7 0 9 2
21 9 2 15 0 9 13 3 1 0 9 2 13 1 0 9 0 9 0 0 9 2
11 9 13 1 9 0 9 1 9 1 11 2
9 9 10 0 9 13 3 3 13 2
19 1 10 9 13 1 0 9 1 0 9 1 0 9 13 3 16 12 9 2
5 9 13 9 11 2
5 9 1 11 13 9
3 9 1 11
4 11 2 11 2
17 11 7 0 9 1 0 9 13 9 0 9 9 1 9 1 11 2
39 0 9 13 9 9 2 1 15 15 13 2 16 2 9 11 13 2 16 9 1 9 7 9 0 2 0 2 0 7 0 9 13 3 9 9 7 9 2 2
7 9 1 9 4 13 3 3
12 1 0 9 13 1 9 9 9 2 13 7 9
2 9 9
5 11 2 11 2 2
21 0 9 3 9 4 13 4 1 9 9 9 7 0 9 13 1 0 9 0 9 2
10 10 9 4 13 3 1 9 1 9 2
6 4 13 9 7 9 2
59 13 15 2 16 4 1 9 1 12 9 13 12 9 2 3 12 9 2 2 1 9 1 9 1 12 1 12 9 12 9 2 12 9 2 2 1 12 1 12 9 12 9 2 12 9 2 7 1 12 9 4 13 12 9 2 12 9 2 2
45 0 0 9 1 0 9 4 13 1 9 13 3 1 12 9 1 9 1 9 1 12 9 0 9 7 1 12 9 1 9 2 10 9 15 13 1 9 1 12 1 12 9 0 9 2
13 0 9 4 13 4 13 1 9 9 1 12 9 2
17 9 4 13 1 9 12 9 2 15 13 1 12 9 3 16 3 2
11 13 4 7 0 9 1 9 7 9 9 2
17 1 12 1 12 9 3 1 9 7 1 12 1 12 9 1 9 2
10 1 9 4 13 9 9 9 12 9 2
22 9 0 1 0 9 4 13 4 3 13 9 12 9 2 3 1 12 9 0 16 3 2
14 13 4 13 4 3 0 2 9 7 15 1 12 9 2
18 9 9 7 0 9 1 0 0 9 13 2 16 9 3 13 13 9 2
18 2 13 7 2 16 4 15 9 0 9 13 3 13 2 2 13 9 2
8 9 9 4 13 1 12 9 2
22 1 0 0 0 9 4 13 13 1 9 2 0 9 4 15 3 13 1 9 12 9 2
14 7 1 0 0 9 4 13 1 12 9 1 10 9 2
18 1 9 9 11 4 1 0 9 9 3 13 0 9 1 9 1 9 2
7 9 4 13 3 9 3 2
12 9 1 10 9 15 3 13 3 12 9 9 2
17 3 10 9 2 7 14 0 2 2 2 3 3 15 9 9 3 13
6 1 11 1 11 0 9
5 11 2 11 2 2
20 9 1 9 9 1 9 11 1 0 0 9 4 9 11 13 1 9 9 11 2
9 0 9 0 9 13 11 0 9 2
9 13 15 3 10 9 11 2 11 2
16 1 11 10 9 11 13 9 10 9 1 11 1 11 3 3 2
7 10 9 13 11 1 0 2
6 11 2 0 9 4 13
5 11 2 11 2 2
30 9 9 1 11 12 13 1 9 2 16 4 1 9 0 9 0 9 11 2 11 2 13 9 1 9 1 11 0 9 2
9 13 15 3 9 9 9 11 11 2
6 9 7 3 3 13 2
26 1 11 15 13 2 16 9 13 1 9 11 3 16 12 9 7 9 1 9 15 3 13 13 0 9 2
25 16 0 9 13 1 9 0 9 2 13 1 11 0 9 9 9 13 2 16 13 9 1 0 9 2
21 3 4 15 13 9 2 16 4 15 13 7 3 15 13 2 16 15 1 9 13 2
4 3 1 9 12
7 0 9 4 9 13 7 9
7 11 2 11 2 11 2 2
19 9 3 13 9 0 13 0 0 9 9 2 1 15 13 1 9 0 9 2
20 1 9 13 12 9 2 12 13 1 2 12 15 15 9 13 7 12 15 13 2
12 0 2 0 2 0 9 9 7 13 10 9 2
11 9 1 10 9 13 1 0 9 1 9 2
44 1 0 9 2 3 13 9 11 2 11 0 2 2 11 2 2 4 13 9 3 10 9 2 15 1 15 13 1 9 0 9 7 10 9 4 1 1 0 9 9 1 9 13 2
18 9 11 13 2 16 4 10 9 13 7 9 0 1 9 0 7 0 2
23 1 0 9 15 7 13 9 13 2 16 4 9 0 13 9 13 14 9 2 7 7 9 2
26 13 7 4 13 2 16 4 1 12 2 9 12 13 7 4 1 15 13 0 9 7 13 9 1 9 2
11 1 10 9 13 0 9 9 1 0 9 2
4 9 1 0 9
22 9 1 9 13 9 13 1 12 9 1 12 2 9 0 9 2 3 9 13 1 9 2
9 1 0 9 13 13 1 12 9 2
11 1 12 9 13 9 7 9 0 9 13 2
17 9 13 13 1 9 0 9 2 15 13 11 2 11 2 11 2 2
28 1 15 13 9 3 2 13 2 16 15 13 0 3 0 9 9 0 1 9 9 12 7 12 7 7 9 13 2
26 3 1 9 9 1 0 9 13 11 9 9 1 9 2 15 4 13 13 0 9 7 0 2 0 9 2
9 9 13 9 9 7 10 9 13 2
31 9 11 11 2 11 2 13 3 3 13 9 1 9 1 0 9 2 16 4 13 9 0 9 3 1 9 0 1 0 9 2
13 2 13 13 0 9 1 0 2 2 13 1 11 2
5 11 13 1 9 9
10 9 11 1 11 0 1 9 11 9 13
2 9 9
7 11 2 11 2 11 2 2
20 9 9 0 9 2 11 2 15 1 10 0 9 13 9 13 9 11 11 9 2
13 3 15 13 9 9 11 7 9 1 9 11 0 2
14 13 7 3 2 16 9 13 1 9 11 0 0 9 2
9 1 9 11 13 4 9 13 3 2
23 12 9 9 11 3 3 0 9 13 1 10 9 2 1 9 13 12 9 1 0 9 2 2
25 0 0 9 4 13 1 9 1 9 2 15 13 9 9 7 0 0 9 1 9 0 9 9 11 2
28 1 9 1 9 9 4 3 12 9 9 9 13 0 9 0 0 2 15 4 16 12 1 9 13 1 0 9 2
11 1 0 9 1 9 9 7 10 9 13 2
28 11 9 10 9 13 0 9 7 13 2 16 11 13 3 2 16 9 9 13 1 0 9 2 3 7 0 0 2
24 1 9 9 9 2 1 15 4 13 9 1 9 9 2 13 2 16 0 9 4 13 1 9 2
35 15 11 13 3 0 0 9 11 11 2 15 13 2 16 3 0 9 2 15 13 9 12 1 9 2 4 13 4 1 9 1 9 9 13 2
8 15 15 1 15 7 13 4 2
19 9 0 3 13 2 16 3 13 1 9 9 2 15 4 13 0 9 13 2
22 10 9 13 13 2 16 13 1 0 9 7 0 9 9 2 7 15 13 1 15 9 2
15 11 2 11 3 13 13 15 0 9 0 11 1 9 12 2
3 3 1 9
20 9 9 13 13 0 0 9 2 2 13 11 11 2 9 9 0 9 0 9 2
3 0 0 9
13 0 9 13 1 0 9 1 9 11 1 9 11 2
13 1 9 1 9 4 1 10 9 9 1 9 13 2
2 9 11
3 9 7 9
2 11 11
15 13 4 0 9 13 0 9 3 1 0 9 7 9 9 2
15 7 13 1 10 9 13 1 10 9 3 9 2 3 9 2
18 1 10 9 15 1 0 9 13 13 9 9 7 3 7 9 0 9 2
26 0 9 1 9 13 1 9 2 16 0 9 9 7 9 1 9 4 13 13 1 0 9 0 0 9 2
25 9 7 3 3 13 9 2 1 15 0 9 2 15 1 9 13 0 9 2 13 1 9 0 9 2
11 7 1 0 9 1 9 3 9 9 3 2
16 12 9 2 0 7 9 3 0 2 13 0 9 7 10 9 2
24 13 15 9 2 3 4 10 0 9 13 13 3 3 1 15 2 15 13 1 0 9 7 9 2
25 10 0 9 4 15 3 14 13 0 9 2 3 4 9 13 0 0 9 0 9 0 1 10 9 2
22 3 1 9 2 3 4 9 3 13 13 0 9 2 3 4 15 13 9 13 10 9 2
30 1 0 9 7 15 13 13 2 16 1 9 2 3 4 13 0 9 2 4 9 7 3 13 9 1 9 1 10 9 2
7 15 13 13 3 0 9 2
14 9 13 3 0 9 9 2 7 13 13 10 0 9 2
6 15 1 15 3 13 2
29 1 9 2 3 13 3 1 0 9 10 9 2 16 10 9 13 7 3 2 13 0 2 16 15 1 15 15 13 2
4 15 13 9 2
23 9 9 1 9 13 13 0 0 9 2 9 9 3 4 13 1 10 9 13 3 0 9 2
3 7 3 2
19 7 1 9 2 16 10 0 9 4 3 1 0 9 3 13 13 10 9 2
25 3 2 9 2 15 4 3 13 0 9 0 9 2 15 3 13 1 10 9 2 15 13 1 9 2
14 9 3 13 2 16 9 4 7 3 13 1 0 9 2
15 13 2 16 0 9 13 13 0 9 9 9 2 0 9 2
14 10 9 3 4 1 0 9 13 1 10 9 1 9 2
6 9 0 11 13 0 9
5 11 2 11 2 2
46 1 9 0 9 7 9 9 15 3 9 13 9 1 0 9 9 1 9 1 15 2 16 13 1 0 7 0 9 9 7 9 1 3 12 9 0 11 2 15 15 13 13 1 0 9 2
22 2 3 4 13 9 3 2 1 11 2 11 7 11 2 2 13 15 9 9 11 11 2
15 1 0 9 9 3 13 3 12 12 0 9 0 1 9 2
18 1 11 11 13 0 9 10 0 11 2 15 1 11 13 13 1 9 2
20 3 1 15 13 9 1 0 9 2 15 1 11 4 3 13 1 0 9 3 2
9 9 9 15 1 9 13 1 11 2
28 1 10 9 9 3 13 1 9 1 11 2 4 15 13 1 9 2 9 2 9 2 9 7 3 1 0 9 2
27 9 9 1 9 7 9 1 10 9 13 10 9 1 9 1 9 1 9 7 0 9 9 9 7 9 9 2
9 9 13 3 1 0 9 0 11 2
13 9 7 15 13 2 16 4 9 1 9 13 9 2
15 9 4 15 1 11 13 13 3 1 9 14 1 12 9 2
43 9 9 15 13 2 16 1 11 4 9 0 9 13 1 0 2 0 0 9 2 15 13 9 1 0 9 2 3 15 3 13 9 1 0 9 2 15 1 11 13 9 9 2
15 9 13 9 1 9 2 16 15 9 13 0 9 7 9 2
9 13 3 7 0 9 7 9 9 2
17 11 11 4 13 2 16 0 9 4 1 0 9 13 7 0 11 2
13 10 0 4 9 13 3 2 0 4 13 0 9 2
22 9 9 1 9 7 9 7 13 1 0 9 0 9 2 1 15 15 9 3 3 13 2
26 13 2 16 9 2 3 13 1 11 13 0 9 1 9 2 15 4 13 9 9 13 2 15 3 13 2
9 9 0 9 4 13 1 9 1 9
5 11 2 11 2 2
19 9 9 7 0 9 0 9 11 11 4 13 9 9 9 0 9 1 9 2
34 1 10 9 13 9 0 9 0 9 2 15 13 11 2 0 7 0 9 2 1 9 0 9 3 16 12 12 9 1 0 9 12 9 2
9 0 9 4 13 3 1 9 9 2
22 9 9 15 15 7 13 3 13 1 12 9 1 9 2 15 4 3 13 12 9 9 2
26 9 11 11 1 9 9 15 13 2 16 3 15 1 10 9 13 3 13 2 16 9 13 3 1 9 2
16 13 7 9 2 16 1 11 2 11 4 13 7 0 0 9 2
21 11 2 11 4 13 1 9 7 3 4 15 13 2 16 4 15 1 0 9 13 2
30 2 13 2 16 4 15 1 3 0 0 9 13 1 0 9 9 2 16 15 15 13 0 9 2 15 13 0 9 9 2
26 9 0 9 13 1 9 1 0 0 0 9 9 7 0 0 9 1 9 9 9 1 9 9 0 9 2
28 0 9 9 7 0 9 13 7 9 13 0 9 1 0 9 1 11 1 9 9 0 9 1 0 0 9 2 2
13 0 9 0 9 9 9 13 1 9 1 9 11 2
14 4 13 3 2 0 2 0 7 0 9 7 9 3 2
18 0 9 11 3 13 10 9 11 11 7 9 0 9 11 9 9 11 2
14 9 1 9 11 1 9 9 1 9 13 13 1 9 2
13 13 15 3 1 9 1 11 9 0 9 11 11 2
28 1 12 9 3 2 16 13 13 0 9 1 9 9 2 4 1 12 2 9 13 9 1 0 9 9 1 11 2
4 0 9 1 11
6 0 9 2 11 2 2
21 1 0 9 1 11 1 0 9 1 9 11 4 13 1 9 3 0 9 1 9 2
12 3 15 13 13 3 0 9 2 9 7 9 2
22 11 2 15 13 3 1 9 13 15 9 0 9 14 1 0 9 2 15 13 0 9 2
20 3 13 3 9 3 13 2 7 13 1 9 13 9 1 9 1 12 2 9 2
5 9 15 13 0 9
5 11 2 11 2 2
57 0 0 9 7 11 11 2 15 13 1 9 12 7 12 1 9 1 0 9 11 7 15 4 1 9 9 9 11 11 3 13 1 9 2 15 15 13 1 0 9 2 15 3 13 10 9 1 11 2 15 13 9 1 9 0 11 2
28 11 11 13 3 1 11 3 3 13 2 7 15 3 13 9 7 0 9 9 11 11 2 9 9 1 0 9 2
14 2 11 15 13 15 13 7 9 4 15 13 3 13 2
22 9 11 13 1 15 0 9 7 16 15 13 3 13 2 3 13 0 1 9 13 3 2
29 13 9 2 16 16 11 3 13 2 13 15 16 0 9 1 9 7 9 9 9 2 2 13 3 9 11 9 11 2
8 1 11 13 1 9 3 12 9
2 9 9
5 11 2 11 2 2
18 0 9 13 1 0 9 3 12 9 2 1 15 12 15 15 13 13 2
14 1 9 1 0 9 1 9 12 13 10 9 3 0 2
33 1 0 0 0 9 13 1 10 9 1 11 2 3 4 1 10 9 1 9 13 0 11 11 2 9 9 0 11 11 11 2 11 2
20 9 13 12 0 9 1 9 1 12 9 2 15 13 9 9 12 9 1 9 2
16 1 9 13 9 0 15 2 16 1 9 9 15 13 10 9 2
10 3 9 1 9 3 12 9 3 13 2
21 9 13 2 16 3 15 13 13 9 9 2 16 7 12 1 9 13 9 1 9 2
33 3 7 9 13 13 10 9 1 15 2 16 1 0 9 9 11 13 1 10 9 2 15 15 9 13 13 2 16 4 13 0 9 2
18 9 3 16 1 9 0 9 0 11 12 2 13 7 1 9 0 9 2
29 1 9 0 9 9 11 2 11 15 7 3 13 9 2 16 4 1 11 13 9 2 15 4 15 9 1 9 13 2
42 1 0 13 3 0 9 9 1 11 2 15 4 13 1 0 9 1 9 2 9 1 9 0 9 1 0 9 7 0 9 0 9 2 15 1 10 9 13 9 0 9 2
13 15 15 3 13 1 9 7 1 9 13 10 9 2
19 1 15 2 16 9 9 13 2 13 9 0 9 9 2 1 15 3 13 2
5 9 1 12 2 9
13 0 0 9 15 13 0 9 9 13 0 9 9 2
42 2 3 15 9 9 13 2 13 4 13 1 13 1 13 2 7 13 15 2 16 12 9 0 0 9 4 13 0 9 1 0 9 9 2 2 13 0 9 9 11 11 2
5 0 9 13 14 12
5 11 2 11 2 2
14 9 0 9 9 0 2 9 2 4 3 13 1 11 2
27 9 1 9 13 9 9 9 12 2 9 7 10 9 11 2 11 13 2 16 4 13 13 13 1 12 9 2
24 1 10 9 13 1 9 9 9 2 15 13 13 14 12 2 9 10 9 7 9 1 15 13 2
17 0 9 9 13 13 1 9 11 11 9 1 9 9 0 0 9 2
40 15 13 12 1 12 9 9 2 0 13 0 9 11 2 0 9 7 11 11 0 2 9 2 2 9 11 7 9 11 0 2 9 2 2 15 13 9 9 9 2
17 1 9 2 15 9 13 2 13 1 9 3 0 9 1 0 9 2
35 1 11 2 0 0 9 2 12 2 12 9 2 9 9 7 9 1 9 13 0 9 9 9 7 9 10 9 3 1 9 0 9 1 9 2
3 9 13 9
5 11 11 2 11 11
34 1 10 9 13 0 9 2 9 9 1 11 2 2 1 15 4 1 9 0 9 3 13 9 0 9 2 11 2 7 10 9 11 9 2
25 11 13 10 0 9 2 13 15 9 9 11 0 2 2 15 13 1 9 9 9 3 0 9 13 2
20 9 2 14 15 13 0 9 1 9 2 3 1 15 9 0 9 13 1 9 2
27 12 9 9 7 13 1 9 11 9 7 13 2 16 4 15 1 10 9 13 9 2 15 1 11 13 9 2
8 1 10 9 13 9 13 3 2
9 13 4 1 15 9 12 9 9 2
16 7 9 0 9 13 9 9 2 1 15 9 1 15 13 3 2
17 9 13 9 13 3 2 16 4 15 13 16 0 9 1 0 9 2
6 9 3 3 9 13 2
25 0 9 9 13 1 0 2 7 13 1 0 9 2 7 9 11 13 2 16 15 1 9 9 13 2
4 11 13 13 9
7 11 2 11 2 11 2 2
29 1 9 9 2 10 0 9 13 0 9 13 3 1 9 2 13 4 13 0 0 9 2 1 15 0 0 9 13 2
18 13 1 0 1 9 2 9 0 9 2 9 0 9 7 9 0 9 2
37 1 9 9 1 9 0 9 2 3 9 0 9 7 9 10 9 2 13 13 1 9 9 9 9 11 2 15 13 7 9 2 1 10 9 9 13 2
15 0 9 13 0 9 11 11 2 11 11 7 0 11 11 2
19 1 9 9 11 11 13 9 0 9 9 2 1 10 9 13 0 9 11 2
13 0 9 13 13 3 1 9 11 1 0 0 9 2
7 11 2 0 9 1 0 9
5 11 2 11 2 2
21 0 9 15 13 0 0 9 0 9 2 15 13 3 1 9 0 9 2 0 9 2
17 9 9 0 9 13 3 12 1 0 9 1 0 9 7 11 0 2
41 1 9 9 9 0 9 11 11 11 0 9 0 9 2 0 1 0 9 9 2 13 9 3 2 9 2 9 7 9 0 9 11 2 15 13 9 3 1 9 9 2
11 9 4 13 1 0 0 9 12 2 9 2
5 9 9 13 7 9
2 11 2
19 0 0 9 1 9 7 0 9 13 1 9 0 0 9 1 12 2 9 2
6 15 12 13 12 9 2
8 0 9 4 1 9 3 13 2
11 0 9 1 10 9 3 0 9 9 13 2
13 10 9 15 1 9 0 9 11 11 3 13 3 2
9 1 9 13 1 11 7 10 9 2
16 9 12 2 9 13 9 9 9 2 0 1 0 9 0 9 2
8 13 13 1 0 9 9 9 2
16 1 0 9 9 9 9 13 0 9 10 0 9 7 0 9 2
5 9 14 13 9 2
26 9 9 9 11 2 11 3 13 2 16 9 13 3 9 1 9 9 11 2 16 1 15 9 13 9 2
21 0 9 11 11 3 13 0 0 0 9 2 1 0 2 11 2 1 9 1 11 2
37 0 9 2 10 9 13 9 2 9 2 0 2 11 2 1 0 2 11 2 2 13 1 0 9 0 9 11 9 10 9 9 9 1 0 12 9 2
21 9 4 13 10 0 9 3 13 1 0 9 9 9 7 3 15 15 3 13 3 2
4 9 11 11 11
19 0 9 1 9 11 11 1 0 9 1 11 4 3 13 0 9 0 9 2
15 11 13 3 12 1 0 9 1 9 2 3 1 0 9 2
9 15 13 9 1 11 1 9 12 2
16 1 9 11 13 9 11 11 2 1 9 2 1 9 0 11 2
5 9 11 11 2 11
8 9 11 3 9 9 9 13 2
13 13 7 2 16 10 9 9 3 0 9 13 9 2
4 9 1 11 13
3 11 2 11
6 2 11 2 11 2 2
26 9 9 11 11 13 2 16 9 9 11 1 9 0 0 9 1 9 0 1 11 13 9 1 0 9 2
27 2 16 4 15 3 13 13 2 3 13 9 2 16 0 9 3 13 0 9 7 9 0 9 2 2 13 2
21 3 13 2 4 13 10 0 9 2 16 10 9 13 0 7 15 15 3 4 13 2
12 2 9 9 4 3 13 2 2 13 11 11 2
20 9 0 9 13 0 9 13 1 0 0 9 1 9 11 9 9 11 11 11 2
12 1 11 15 4 13 0 2 9 2 0 9 2
12 9 0 0 9 0 9 3 13 2 13 9 2
6 0 9 13 13 3 3
5 11 2 11 2 2
15 3 13 9 2 16 4 15 9 1 9 13 1 0 9 2
15 13 15 0 9 9 13 9 0 9 9 1 9 1 9 2
24 16 4 15 9 1 0 9 1 9 1 0 2 9 13 2 0 9 4 15 3 3 13 13 2
25 9 13 9 9 13 0 9 1 9 7 1 9 2 1 15 0 9 13 9 2 10 9 9 13 2
31 11 13 9 0 9 2 16 1 9 9 13 9 3 9 2 15 13 1 12 9 9 2 7 15 7 9 10 9 1 9 2
25 1 15 2 3 13 0 9 1 9 0 9 1 9 2 15 13 13 2 16 10 9 13 3 0 2
8 13 15 3 10 9 11 11 2
17 11 2 0 2 9 2 0 9 0 9 1 12 2 9 13 4 2
22 11 2 11 2 3 0 9 9 2 3 13 2 16 1 9 13 1 9 13 9 9 2
30 1 0 9 13 2 16 9 4 13 9 9 2 7 13 2 16 9 1 9 0 9 13 14 0 9 0 9 0 9 2
14 3 1 10 9 3 9 1 0 0 9 13 9 9 2
12 9 13 0 9 0 0 9 9 2 11 2 2
32 9 2 15 13 9 2 13 1 9 12 9 2 3 9 11 2 1 9 1 0 9 1 9 9 2 15 15 13 9 12 9 2
14 9 9 7 9 1 0 9 13 1 0 0 9 0 2
11 11 3 13 9 1 10 0 9 10 9 2
14 9 11 13 1 15 2 15 4 15 13 13 2 13 2
36 9 0 9 11 1 9 3 13 2 16 1 12 9 13 1 11 1 11 12 9 9 2 15 13 3 2 0 7 0 9 2 2 15 3 13 2
22 16 15 9 9 13 1 0 9 2 13 4 0 2 16 4 15 0 9 3 3 13 2
18 13 15 9 0 0 9 11 2 11 2 15 13 0 9 1 9 9 2
24 0 11 13 9 0 9 1 0 9 1 0 9 10 0 9 2 3 1 9 9 0 0 9 2
6 9 15 13 1 0 9
5 11 2 11 2 2
12 9 0 9 15 3 13 1 9 9 1 9 2
12 1 0 0 9 11 15 13 10 9 11 11 2
28 0 0 9 13 2 16 13 9 0 2 3 13 9 2 7 16 4 13 0 2 0 9 1 9 11 2 11 2
12 15 13 1 12 9 0 9 13 12 9 3 2
42 0 9 11 2 11 2 15 4 0 9 13 2 13 1 15 2 16 1 0 0 9 15 4 13 1 12 0 9 7 1 0 9 1 12 0 9 0 1 12 0 9 2
14 3 13 0 2 10 9 4 13 9 1 0 0 9 2
15 11 13 2 16 4 15 9 0 9 13 1 9 0 9 2
7 11 13 1 11 1 0 9
2 9 9
9 9 2 11 2 11 2 11 2 2
37 1 9 3 12 9 2 9 7 9 7 1 9 2 9 7 9 1 0 2 0 7 0 11 13 9 0 0 9 2 3 0 2 0 9 11 11 2
7 9 10 9 13 9 9 2
14 1 9 0 9 1 9 7 0 9 11 13 1 9 2
10 13 15 7 13 1 10 9 11 11 2
11 15 0 13 7 13 15 7 10 0 9 2
13 9 9 0 9 1 9 0 9 13 1 9 0 2
23 0 9 1 11 0 9 1 10 9 13 2 7 9 3 13 0 9 15 0 9 7 9 2
36 11 4 0 13 3 3 2 1 0 11 11 2 11 2 0 9 11 3 2 2 1 0 11 1 0 9 0 11 1 9 2 0 9 7 9 2
20 9 13 3 1 15 2 16 3 9 11 1 11 10 9 13 3 1 9 12 2
19 0 4 15 3 13 1 11 2 15 4 13 1 9 9 1 9 0 9 2
26 1 0 9 15 3 13 1 9 9 11 11 11 11 2 15 13 12 9 9 1 11 1 9 9 12 2
31 9 9 11 13 0 9 11 1 9 9 1 9 12 2 2 16 13 1 9 0 0 9 7 13 0 9 1 0 9 2 2
29 0 9 11 13 1 9 9 1 10 9 1 9 12 3 3 2 16 11 13 1 9 9 0 9 7 13 1 9 2
6 9 11 11 9 13 2
7 7 1 9 4 13 13 9
5 11 2 11 2 2
20 9 9 15 1 9 9 1 0 9 13 3 1 9 9 7 9 3 0 9 2
17 10 9 13 3 1 9 1 9 9 11 1 11 9 9 11 11 2
25 9 3 13 2 16 9 13 1 10 9 9 13 0 9 7 13 15 1 9 0 9 1 10 9 2
25 11 9 13 1 9 1 0 9 9 11 11 12 9 1 9 0 9 7 9 2 15 4 9 13 2
5 9 9 13 9 9
2 11 2
23 0 9 9 9 1 0 9 11 11 1 9 0 9 9 4 9 9 9 2 11 2 13 2
23 7 15 3 2 16 15 13 9 9 0 9 2 15 4 3 13 1 0 9 0 0 9 2
9 9 11 15 13 1 0 0 9 2
26 2 16 15 9 13 2 3 1 0 9 13 0 13 0 9 16 13 9 2 2 13 9 11 11 11 2
18 2 3 7 13 0 9 1 15 2 16 15 15 13 9 1 9 9 2
13 1 15 15 13 9 9 7 1 9 3 13 2 2
29 9 11 13 1 9 9 0 9 2 0 11 1 0 9 4 3 13 12 9 2 15 13 1 12 9 3 16 3 2
3 11 1 9
5 11 2 11 2 2
26 9 9 11 11 13 2 16 9 9 11 1 9 0 0 9 1 9 0 1 11 13 9 1 0 9 2
27 2 16 4 15 3 13 13 2 3 13 9 2 16 0 9 3 13 0 9 7 9 0 9 2 2 13 2
23 3 13 2 4 13 10 0 9 2 16 10 9 13 0 7 15 15 1 15 3 4 13 2
12 2 9 9 4 3 13 2 2 13 11 11 2
4 11 1 0 9
5 11 2 11 2 2
26 12 1 9 2 15 13 0 9 2 11 2 13 0 9 9 2 13 15 2 9 13 0 9 1 9 2
18 2 15 13 2 16 4 9 4 13 1 0 7 3 0 0 9 2 2
21 1 9 11 4 13 0 13 0 9 0 9 16 9 2 15 4 13 14 3 0 2
29 0 9 13 1 15 2 16 4 15 9 7 10 9 13 1 9 1 9 2 13 15 7 2 16 13 0 13 9 2
29 13 4 9 7 1 0 9 2 7 1 15 2 16 4 13 0 13 1 0 9 0 9 2 3 7 1 9 9 2
8 9 11 0 1 11 13 0 13
5 11 2 11 2 2
17 0 9 1 9 0 9 1 11 7 11 13 0 9 1 12 9 2
19 10 9 13 10 9 9 9 7 0 9 1 0 9 2 15 13 1 11 2
35 9 9 7 0 9 11 11 1 10 9 3 13 2 16 0 9 13 1 15 2 16 4 0 9 4 13 1 9 2 1 15 0 9 13 2
35 0 9 10 9 9 2 15 13 10 9 1 9 2 4 3 13 2 16 4 7 1 10 9 13 2 16 10 7 15 0 9 13 0 9 2
22 0 9 4 11 13 1 10 9 1 11 2 0 9 1 9 7 0 9 11 2 11 2
21 1 9 13 13 9 1 12 9 1 9 2 15 15 13 3 1 0 7 0 9 2
14 9 11 7 11 13 3 0 2 16 13 1 0 9 2
19 11 13 13 9 1 9 1 9 7 15 3 1 9 7 9 1 12 9 2
4 9 7 0 9
22 1 9 9 4 13 13 9 1 11 14 10 0 9 2 15 13 0 0 9 1 9 2
16 3 3 13 9 1 15 2 16 3 0 9 0 9 3 13 2
26 9 13 13 7 0 2 7 13 2 16 14 0 2 9 9 0 0 9 1 0 9 1 0 9 9 2
16 1 0 9 0 9 4 9 13 2 9 9 13 0 9 2 2
16 0 9 13 14 13 14 0 9 9 2 7 7 0 0 9 2
16 13 3 3 0 9 2 15 0 9 1 0 9 0 9 13 2
17 0 15 1 10 9 13 2 14 4 15 0 4 13 3 1 15 2
12 9 4 15 13 1 15 9 2 0 7 0 2
19 3 7 13 9 0 9 1 0 9 11 11 2 9 15 1 15 13 3 2
11 13 7 13 2 1 1 10 0 2 0 2
12 14 9 2 7 9 4 13 13 9 1 9 2
13 13 10 9 4 13 13 9 2 7 9 9 9 2
8 12 0 9 3 12 0 9 2
12 11 13 0 9 3 13 7 1 15 0 9 2
9 1 0 9 15 13 13 0 9 2
24 1 9 0 0 9 13 3 3 3 0 2 16 0 2 0 9 15 1 0 9 13 3 13 2
17 0 9 9 13 1 0 9 0 2 3 3 0 2 9 7 9 2
12 13 13 9 9 2 0 9 2 0 9 0 2
26 16 13 10 9 1 9 0 9 2 9 2 0 9 2 9 9 1 9 7 15 0 2 13 3 0 2
18 0 9 3 13 13 0 9 14 1 0 0 9 2 9 0 9 2 2
6 9 0 9 9 13 2
10 13 0 1 0 9 13 3 0 9 2
17 7 10 9 4 7 13 4 1 11 13 1 9 1 0 0 9 2
20 0 9 0 0 9 2 15 13 13 9 0 9 2 13 1 9 11 7 11 2
17 0 9 9 1 0 0 9 13 0 1 0 9 13 3 1 9 2
15 3 1 9 7 13 2 10 9 13 0 9 7 0 9 2
6 9 0 9 4 13 9
5 11 2 11 2 2
10 0 9 7 9 4 1 11 13 9 2
31 9 10 0 9 13 1 0 9 2 9 1 9 9 7 10 9 7 9 1 9 9 2 9 2 0 7 0 9 3 9 2
30 13 15 1 9 1 9 1 0 9 7 9 2 15 3 12 9 13 0 9 2 12 9 13 1 2 12 15 13 2 2
18 9 13 9 13 7 1 9 2 13 15 13 3 1 9 7 0 9 2
25 9 13 9 1 0 9 1 9 3 12 7 3 12 9 9 2 16 1 9 13 3 12 9 9 2
12 1 9 1 9 7 9 15 13 9 9 9 2
21 1 9 4 9 13 13 1 9 2 16 4 13 9 0 7 0 0 9 1 9 2
7 13 15 4 0 0 9 2
26 9 1 9 2 3 9 9 1 12 12 9 1 12 9 2 13 13 14 1 9 1 9 7 9 9 2
14 1 15 4 13 13 0 9 1 9 9 2 3 9 2
18 1 1 15 2 16 9 4 9 13 2 13 10 9 13 10 0 9 2
10 9 11 13 13 9 3 0 0 9 2
9 9 13 1 9 1 9 0 9 2
23 9 13 1 0 9 9 0 9 1 3 16 12 9 9 2 3 15 13 3 3 12 9 2
19 9 7 9 13 0 13 10 9 1 9 1 9 1 12 9 1 9 9 2
5 11 2 9 1 9
4 9 9 11 11
19 2 13 0 9 2 2 13 3 3 16 3 11 11 2 0 0 0 9 2
7 13 3 0 9 2 9 2
38 7 3 9 2 13 2 14 2 16 1 0 12 9 13 13 0 0 0 9 1 11 2 16 13 1 0 12 9 2 13 1 9 2 0 9 0 11 2
6 7 16 13 13 9 2
6 7 2 13 3 13 2
34 13 14 14 13 0 9 2 13 2 0 9 0 9 2 2 3 2 13 9 0 0 9 2 3 13 9 7 0 0 9 2 2 2 2
21 3 15 13 9 0 7 0 2 13 9 11 9 1 9 11 9 2 14 9 9 2
19 1 0 9 13 9 1 0 9 7 9 2 7 3 13 3 3 0 9 2
20 3 7 9 2 3 0 1 0 9 1 9 2 13 13 1 0 9 1 9 2
21 9 9 9 13 0 9 11 11 2 0 9 1 11 11 11 2 11 11 2 2 2
5 15 1 15 13 2
15 16 0 9 13 0 9 1 11 0 9 13 1 9 0 2
11 0 10 9 13 0 9 13 0 11 12 2
16 16 15 15 9 13 2 13 13 1 9 11 12 7 11 12 2
7 15 13 10 9 2 11 2
17 9 15 7 13 3 3 13 9 1 10 9 1 0 9 0 9 2
11 15 13 9 2 3 1 11 1 9 9 2
38 3 15 13 13 7 1 0 9 2 1 9 15 13 9 0 11 2 9 11 7 11 2 0 9 11 7 11 2 16 4 15 13 2 16 15 13 9 2
10 13 13 1 12 1 9 9 9 11 2
8 13 15 0 9 1 11 0 2
13 1 9 9 15 13 9 2 0 0 13 9 11 2
17 15 2 7 14 15 2 13 1 9 11 2 3 13 0 9 11 2
13 0 9 13 13 10 9 2 13 9 0 9 9 2
16 10 0 13 2 16 4 13 9 2 13 4 15 2 7 3 2
11 0 1 10 0 9 13 9 1 9 9 2
23 9 1 11 13 9 2 3 12 2 9 9 2 13 2 7 16 10 0 9 1 15 13 2
14 1 12 9 4 13 0 13 15 9 1 12 11 9 2
6 7 13 9 7 9 2
17 10 9 7 13 2 0 2 1 0 9 2 15 15 13 0 9 2
23 3 0 9 13 0 9 2 0 9 2 2 1 15 9 9 13 9 9 0 3 1 9 2
15 2 3 15 13 13 1 15 2 2 13 0 9 10 9 2
44 13 15 3 9 9 2 15 15 1 9 0 9 1 0 12 9 13 2 9 2 0 9 13 1 9 2 1 12 9 9 2 3 12 9 9 2 2 7 3 12 0 9 9 2
48 0 11 11 2 3 1 10 0 9 2 13 9 2 2 13 0 11 1 9 2 16 4 2 13 11 2 2 3 13 2 7 16 4 15 13 13 10 3 0 0 9 2 3 13 10 9 2 2
66 16 4 13 10 9 2 16 4 13 0 9 0 9 11 11 2 7 3 16 4 13 12 9 9 2 15 15 13 9 1 0 9 2 16 13 3 2 0 2 9 2 3 3 13 11 9 9 10 9 2 12 5 9 9 11 13 1 9 7 13 15 14 0 11 11 2
14 7 1 12 9 0 9 13 0 13 15 9 1 9 2
8 13 1 15 3 16 0 9 2
4 11 13 0 9
2 11 2
25 9 11 7 9 11 15 1 9 13 1 0 9 9 9 7 13 1 15 1 0 7 0 9 11 2
34 1 9 0 9 15 13 2 16 9 13 1 9 9 11 1 9 1 9 0 9 1 11 2 10 9 13 9 11 9 9 0 9 11 2
10 11 13 1 9 1 9 7 0 9 2
16 9 1 9 0 9 1 9 2 15 13 1 0 11 2 13 2
6 11 1 9 3 13 2
5 11 13 9 1 11
3 0 11 2
28 9 11 7 11 15 13 2 3 2 2 7 3 13 13 2 3 4 13 9 9 13 13 7 13 9 1 11 2
18 1 0 11 15 13 9 0 9 1 9 9 9 9 1 11 11 11 2
18 2 0 9 2 13 9 11 1 15 9 2 3 7 1 9 0 9 2
34 1 9 1 9 13 2 16 0 9 3 13 1 9 11 7 13 2 16 10 9 15 1 9 13 13 3 3 2 16 4 3 13 9 2
5 9 1 11 7 13
2 11 2
28 3 0 9 1 9 13 1 9 1 9 9 1 0 11 13 9 1 10 0 9 1 11 1 0 7 0 9 2
34 0 9 0 9 1 0 9 11 2 11 3 13 2 16 9 1 9 9 15 13 13 2 16 0 9 7 9 0 11 14 13 0 9 2
10 9 11 1 9 9 1 9 9 1 11
4 11 2 11 2
26 12 9 0 9 13 9 0 1 9 0 9 1 11 2 16 4 3 9 13 9 15 15 13 1 11 2
26 9 13 0 9 2 16 4 13 3 0 9 0 1 11 2 7 13 15 2 16 4 13 0 9 9 2
9 9 4 13 9 11 11 1 9 2
17 9 0 11 13 0 9 2 15 11 13 1 11 7 0 9 11 2
15 13 7 0 9 1 11 2 3 15 3 3 13 0 9 2
24 2 1 0 9 1 11 4 13 15 0 9 2 3 12 2 2 13 9 9 1 11 11 11 2
20 1 11 13 7 12 1 12 9 1 11 3 13 3 2 3 15 13 9 11 2
13 1 0 9 1 11 4 1 9 13 12 0 9 2
32 9 11 1 0 11 15 13 2 0 9 2 2 3 13 0 1 9 13 0 0 9 1 1 15 2 16 0 9 9 4 13 2
12 13 15 9 0 9 11 2 11 2 11 11 2
20 1 10 9 13 1 9 14 12 9 0 9 2 3 9 13 13 3 1 9 2
4 0 9 13 9
2 11 2
18 0 9 13 12 9 7 9 0 0 9 2 15 9 4 13 9 9 2
12 11 2 11 7 11 2 11 13 13 1 9 2
12 9 15 13 2 16 4 13 1 0 9 13 2
16 9 0 9 7 9 13 3 9 9 2 16 4 13 9 13 2
23 0 0 9 2 15 9 13 13 2 15 13 1 0 9 9 0 9 0 0 0 9 11 2
36 0 9 13 10 9 2 12 0 9 9 1 11 15 13 2 0 9 2 1 12 9 2 16 4 15 13 13 1 9 9 1 9 1 9 9 2
4 9 11 2 11
8 9 11 11 12 2 15 13 9
2 11 2
26 9 11 11 12 2 2 15 15 1 9 1 9 13 9 2 15 3 1 9 13 1 0 9 11 9 2
18 13 15 9 11 2 12 1 12 9 2 1 10 9 15 9 3 13 2
23 0 9 2 15 4 3 3 13 2 13 2 16 1 9 0 0 9 13 3 1 0 9 2
23 0 9 11 11 2 11 3 13 9 10 9 2 1 15 9 1 9 7 1 15 13 9 2
5 1 11 9 0 9
2 11 2
25 9 9 1 0 9 13 3 3 1 9 11 1 0 0 9 11 2 15 13 12 1 9 9 11 2
15 13 15 3 1 9 0 9 1 9 2 16 4 13 9 2
11 9 13 0 9 1 9 2 15 13 9 2
22 1 9 0 9 15 13 9 1 0 9 2 9 0 9 9 1 9 9 11 7 11 2
22 11 13 1 9 15 9 0 9 2 7 3 13 13 10 9 9 2 15 13 0 11 2
3 9 0 9
2 11 2
13 9 11 11 11 3 13 9 1 9 9 0 9 2
18 9 1 10 9 13 2 9 11 2 2 15 1 9 13 0 9 11 2
40 1 9 1 0 0 9 1 11 11 13 2 16 0 9 13 13 1 9 0 9 0 1 9 0 0 9 2 11 2 2 0 0 9 2 9 9 7 0 9 2
33 2 9 0 9 7 9 1 9 0 9 4 13 1 9 9 0 9 2 2 13 9 11 9 9 2 15 13 13 0 9 0 9 2
26 11 13 0 0 9 2 16 4 1 12 9 13 7 13 9 2 3 4 13 0 0 9 9 9 11 2
17 0 9 13 9 2 16 4 15 0 9 0 9 13 1 0 9 2
11 10 9 13 9 11 7 9 13 7 9 2
25 9 0 9 1 0 9 11 11 2 11 2 11 7 9 10 0 9 4 1 9 3 13 9 9 2
5 13 15 0 9 2
26 1 12 9 9 13 0 9 9 11 2 11 2 0 1 9 0 0 9 1 9 0 0 9 1 11 2
25 11 4 13 3 1 9 12 9 9 7 1 9 9 1 9 3 12 9 9 2 15 13 9 11 2
37 0 9 0 0 9 4 13 9 3 2 16 9 11 13 15 2 16 9 1 9 9 9 2 15 13 10 9 2 4 13 16 0 9 0 0 9 2
10 0 9 13 9 11 11 2 11 9 2
10 1 9 15 13 9 11 11 2 11 2
15 16 9 13 9 2 1 15 13 12 9 7 1 14 12 2
14 0 9 11 13 3 9 9 7 9 9 0 11 11 2
24 10 0 9 2 0 1 0 9 11 2 11 2 13 1 9 9 9 9 1 11 7 0 9 2
31 0 0 9 9 0 2 15 13 0 10 9 1 9 9 9 11 2 13 9 1 0 9 2 16 10 9 13 0 9 11 2
8 13 15 3 0 9 0 11 2
5 9 11 13 0 11
2 11 2
19 0 9 13 9 0 9 0 11 7 13 9 1 9 0 9 0 2 11 2
27 12 9 2 15 1 9 13 9 11 2 13 9 1 15 2 16 9 11 13 1 9 0 9 0 9 11 2
33 1 9 2 15 3 13 13 9 2 15 13 9 9 0 1 0 9 1 9 12 2 15 13 11 1 0 9 9 9 0 2 11 2
28 0 9 0 11 13 1 9 0 11 7 13 13 1 11 2 9 2 11 2 11 2 11 2 0 11 7 11 2
10 9 1 10 9 13 12 9 9 3 2
8 11 7 11 13 9 1 0 9
4 11 2 11 2
35 0 9 9 11 11 7 9 0 9 11 11 11 3 1 11 13 9 2 15 13 9 1 0 9 1 11 7 0 0 9 1 11 7 11 2
40 1 3 16 12 9 0 9 15 3 11 7 11 13 13 15 1 9 0 9 1 9 9 2 9 2 9 2 9 2 9 2 9 2 0 9 7 1 0 9 2
11 9 1 9 9 9 13 0 9 11 11 2
18 12 9 13 0 9 2 16 4 13 11 1 9 0 9 0 0 9 2
16 11 13 0 0 0 9 1 11 7 11 1 0 1 0 9 2
32 2 13 0 9 7 0 9 2 16 4 3 13 13 0 9 0 9 2 15 13 13 0 9 2 2 13 11 1 0 0 9 2
10 13 2 16 11 4 13 1 0 9 2
30 0 9 0 9 13 4 1 9 13 3 1 12 2 7 14 1 12 9 9 0 9 1 9 11 7 1 0 9 11 2
9 13 15 3 0 9 9 11 11 2
50 2 13 4 15 2 1 9 1 11 1 11 2 13 11 0 9 2 15 13 3 9 7 9 7 15 13 12 9 2 3 1 9 2 3 4 13 0 9 9 2 2 13 11 1 9 1 0 0 9 2
13 0 9 9 11 11 13 1 9 1 9 1 11 2
24 13 15 1 0 9 11 11 7 13 1 15 1 0 9 11 1 11 2 15 13 1 0 9 2
14 1 9 13 0 9 9 9 11 1 9 1 0 9 2
2 9 9
20 1 9 1 12 9 13 1 0 11 0 9 0 0 9 11 11 7 11 11 2
7 12 9 13 9 0 9 2
15 0 1 9 9 2 9 11 11 13 1 11 3 1 9 2
16 1 9 1 12 1 12 2 9 13 1 9 0 9 9 9 2
13 9 11 11 13 1 11 1 11 3 1 0 9 2
20 13 13 1 9 9 2 3 16 11 11 2 15 13 1 11 3 1 9 2 2
19 12 15 13 1 0 9 1 9 2 15 13 13 1 9 1 12 1 12 2
9 3 13 1 9 9 1 0 9 2
12 1 9 4 15 12 13 13 9 1 0 9 2
32 1 10 0 9 1 11 13 9 1 3 0 11 9 9 11 2 3 0 0 9 1 11 2 9 1 0 9 9 2 7 0 2
9 13 1 9 1 0 9 3 0 2
9 12 9 3 13 9 1 0 9 2
17 9 2 15 15 13 1 9 9 2 13 9 1 9 14 12 9 2
23 1 9 13 7 13 9 1 12 9 2 9 7 0 9 1 9 2 15 13 3 1 9 2
12 9 1 9 15 4 13 1 9 1 12 9 2
10 1 9 1 11 13 10 9 12 9 2
7 13 14 1 12 0 9 2
11 3 16 9 9 13 9 3 9 0 9 2
18 9 1 9 4 13 13 9 1 9 11 11 2 10 9 13 0 9 2
2 15 2
3 3 2 3
30 0 9 1 11 11 13 3 3 2 12 2 9 9 11 1 9 1 9 11 11 2 9 11 11 2 9 11 11 2 2
19 9 9 9 13 13 3 3 1 9 11 0 9 11 11 7 0 9 11 2
20 9 1 9 13 9 2 15 4 13 1 0 9 0 9 11 1 12 2 9 2
15 0 9 11 13 3 1 12 9 0 9 1 9 11 11 2
18 9 0 9 13 3 1 12 9 9 11 11 1 12 2 9 9 9 2
19 13 11 11 2 9 2 2 11 11 2 9 2 7 11 0 2 9 2 2
20 0 9 11 13 3 3 2 12 2 9 9 11 11 9 9 1 9 11 11 2
16 9 11 11 1 9 13 9 1 9 1 0 9 1 11 9 2
3 9 1 11
2 9 2
27 1 12 9 0 1 9 2 1 11 7 1 9 1 9 2 11 2 11 2 11 3 13 0 9 11 11 2
33 3 2 1 0 9 7 1 9 0 9 0 9 11 2 10 2 9 0 9 1 9 9 0 2 2 9 1 9 2 0 9 12 2
25 9 7 9 0 0 1 9 13 1 15 2 16 11 13 3 13 9 0 9 2 0 1 0 9 2
18 9 7 9 0 9 10 9 15 13 1 10 3 0 9 1 0 9 2
29 1 9 9 1 9 11 3 3 13 2 0 9 2 2 7 3 3 16 1 9 9 13 13 1 9 1 9 9 2
27 9 1 9 9 0 9 1 9 2 10 9 2 9 7 0 9 3 13 16 0 9 1 10 9 9 9 2
17 1 11 1 0 2 1 0 9 1 9 2 1 12 11 1 11 2
8 15 1 9 1 0 0 9 2
38 0 15 15 13 13 10 9 2 3 13 9 3 13 9 7 3 13 2 1 0 9 2 0 9 2 3 0 9 2 3 13 9 0 2 0 2 9 2
30 10 9 13 7 14 9 2 7 9 3 3 13 1 0 9 7 1 9 11 11 15 15 3 13 13 9 0 0 9 2
31 1 0 9 2 1 11 0 7 0 7 1 11 0 9 2 16 3 14 0 2 15 3 3 13 9 9 2 9 10 9 2
21 15 9 1 12 10 2 0 2 9 3 13 2 13 2 14 15 9 3 2 2 2
6 13 1 10 0 9 2
15 9 2 0 9 2 9 2 10 2 9 0 2 7 13 2
4 11 11 2 11
8 10 9 1 0 11 2 2 2
2 11 11
17 0 9 9 0 11 1 15 1 9 9 0 9 13 3 0 9 2
6 3 10 0 9 13 2
25 15 3 13 13 2 9 9 1 9 2 9 0 9 1 0 9 2 7 9 0 9 9 0 9 2
19 13 3 0 2 3 3 15 11 11 13 0 9 1 9 11 2 9 9 2
24 1 0 0 0 9 11 11 11 1 9 0 9 11 11 13 10 9 13 16 12 2 9 12 2
45 0 13 15 2 16 1 9 12 2 12 13 0 9 0 0 9 2 0 0 9 11 11 2 1 9 11 11 12 1 0 0 9 2 3 13 1 9 0 9 2 7 15 0 9 2
26 0 0 7 0 9 9 0 11 13 3 0 2 3 0 0 9 13 9 9 0 2 3 16 3 0 2
15 13 3 9 2 10 9 1 0 9 13 9 0 11 3 2
17 2 16 4 13 0 9 2 0 9 9 7 3 0 0 9 2 2
13 13 3 7 9 2 10 9 13 9 16 0 9 2
12 9 13 3 10 9 2 9 13 0 9 9 2
13 13 3 14 1 9 7 1 0 0 9 0 11 2
25 13 1 15 2 16 14 13 15 2 14 15 13 2 3 13 2 14 13 15 2 13 1 0 11 2
25 13 15 15 7 10 9 2 3 10 0 9 9 7 9 2 0 15 1 3 0 9 0 0 9 2
31 9 1 9 2 9 7 9 15 3 3 3 13 2 3 16 3 0 9 9 9 1 9 3 0 9 0 0 9 11 11 2
29 9 0 11 2 15 13 11 11 3 2 13 9 9 2 7 3 15 13 1 10 0 9 2 1 15 13 3 0 2
12 9 3 13 0 1 9 9 16 0 9 9 2
21 13 9 9 1 15 10 9 7 1 10 0 9 0 9 7 9 2 7 3 9 2
16 3 1 0 9 3 15 9 13 7 15 13 3 13 2 2 2
12 3 13 9 10 9 2 3 0 9 0 11 2
13 0 7 0 9 4 13 2 7 13 15 15 15 2
7 15 13 9 7 15 9 2
12 15 13 3 2 9 7 9 9 11 11 11 2
9 1 15 15 1 9 4 13 9 2
5 9 7 9 9 2
11 0 9 9 9 13 0 9 1 9 3 2
48 9 13 9 10 9 1 0 9 2 16 15 1 0 9 9 13 0 9 0 1 0 9 7 3 13 1 9 7 9 9 0 9 2 7 0 0 0 9 2 11 0 2 11 11 7 11 11 2
22 9 2 15 15 1 3 3 9 13 0 2 7 16 0 9 2 13 3 1 9 0 2
41 9 0 3 3 1 9 2 11 11 2 11 0 2 11 9 2 3 13 13 9 7 10 9 13 1 12 9 2 0 1 9 2 7 1 0 0 9 1 0 9 2
9 1 10 9 15 7 0 9 13 2
13 3 3 9 13 9 13 15 2 7 13 15 3 2
31 3 2 3 1 0 0 9 0 9 9 2 9 0 9 11 0 2 0 16 9 7 3 3 3 0 0 2 0 9 2 2
16 3 3 1 9 0 9 9 11 11 2 0 9 9 3 3 2
23 7 3 9 11 11 2 1 15 9 9 9 1 15 13 2 10 9 10 9 13 2 2 2
17 0 7 13 9 2 9 2 1 0 9 2 0 3 1 10 9 2
29 10 9 13 0 0 9 9 9 2 15 13 1 9 13 1 3 0 9 2 16 4 13 0 9 3 13 7 13 2
26 3 7 9 13 3 1 0 0 9 7 0 0 9 13 3 1 0 9 3 2 0 2 9 11 11 2
16 11 13 1 0 9 0 2 9 2 2 1 15 10 9 13 2
6 3 2 10 0 9 2
2 11 11
5 9 11 11 0 9
18 9 2 16 10 0 9 13 1 9 0 9 2 15 3 13 0 9 2
21 9 0 9 2 0 0 9 11 11 7 0 1 12 0 0 9 2 13 9 0 2
19 3 0 9 0 9 3 13 3 3 7 3 2 16 15 13 1 0 9 2
23 13 15 13 2 3 15 9 13 3 1 9 2 0 9 2 11 11 2 15 7 3 13 2
26 9 1 9 2 1 15 15 13 9 9 1 3 0 9 7 0 9 2 15 13 9 3 1 0 9 2
28 1 9 0 9 16 4 13 3 0 0 9 7 10 9 1 2 9 1 9 2 2 1 15 15 3 3 13 2
23 9 2 15 15 9 11 13 1 9 10 3 0 9 2 11 11 2 13 13 13 0 9 2
57 0 9 2 9 2 11 11 2 7 0 9 2 9 2 11 11 2 15 1 0 9 3 13 3 16 0 9 2 3 1 9 2 1 15 0 1 9 13 1 0 9 2 2 16 16 9 2 15 15 3 13 0 9 1 0 9 2
31 13 9 7 9 2 9 13 9 3 0 2 0 0 9 2 0 9 1 0 9 1 9 2 2 15 9 15 13 1 9 2
32 13 15 7 1 9 0 9 9 7 0 9 2 0 3 16 9 0 9 2 1 9 2 2 0 1 2 0 2 9 9 0 2
22 0 0 9 15 3 3 13 1 0 9 2 13 7 1 15 2 15 13 0 2 2 2
18 0 9 11 11 7 0 0 9 9 7 9 13 1 3 16 12 9 2
18 3 1 10 9 13 1 0 9 13 0 9 2 15 15 13 0 9 2
18 13 2 14 7 13 0 9 7 3 0 9 2 0 0 9 1 9 2
14 9 11 10 9 13 9 0 9 11 11 7 11 11 2
6 12 9 13 12 9 2
45 11 2 9 2 9 2 0 2 2 11 11 12 2 12 12 11 12 2 9 2 2 12 2 12 12 12 2 12 2 12 12 12 0 9 0 9 2 11 12 2 12 12 11 1 11
3 11 11 3
24 0 9 11 11 2 9 9 0 9 2 13 10 0 9 1 9 9 1 9 9 3 1 11 2
21 2 9 13 13 7 1 9 0 9 2 7 1 9 9 2 7 1 0 0 9 2
22 3 9 13 9 2 1 15 13 13 0 9 2 15 13 1 0 9 2 2 13 11 2
12 10 9 1 0 9 13 1 9 1 12 9 2
3 2 11 2
13 9 0 0 9 11 11 2 12 2 13 9 9 2
24 3 1 0 9 1 9 0 2 11 0 13 3 11 9 2 1 15 0 7 0 9 13 9 2
28 10 9 9 7 10 9 13 1 9 11 11 7 11 11 3 0 9 1 9 2 15 1 0 9 13 0 9 2
8 1 9 13 1 12 2 9 2
5 9 11 9 2 11
4 13 3 12 9
7 11 7 11 13 1 0 9
2 9 9
19 3 1 12 9 13 1 0 11 0 9 0 0 9 11 11 7 11 11 2
6 12 9 13 0 9 2
2 11 11
15 0 1 9 9 2 9 11 11 13 1 11 3 1 9 2
14 3 1 9 1 0 9 13 1 9 0 9 9 9 2
18 13 13 1 9 9 2 3 16 11 11 2 15 13 3 1 9 2 2
16 12 15 13 1 0 9 1 9 2 15 13 13 1 0 9 2
9 3 13 1 9 9 1 0 9 2
14 1 0 9 4 15 3 12 13 13 9 1 0 9 2
32 1 10 9 1 9 1 11 13 9 1 3 0 11 9 9 11 2 0 0 9 1 11 2 9 1 0 9 9 2 7 0 2
9 13 1 9 1 0 9 3 0 2
9 12 9 3 13 9 1 0 9 2
18 9 2 15 15 1 9 13 9 2 13 9 1 9 14 12 12 9 2
22 1 9 13 13 9 1 12 9 2 9 7 0 9 1 9 2 15 13 3 1 9 2
14 9 1 9 15 4 13 3 1 12 9 1 9 11 2
17 13 14 1 12 0 9 7 1 9 1 11 10 9 13 9 9 2
11 3 16 9 9 13 9 3 9 0 9 2
19 9 1 9 4 15 13 13 9 1 9 11 11 2 10 9 13 0 9 2
13 9 11 11 1 0 9 0 9 1 9 1 0 11
2 9 11
1 9
3 0 11 2
12 0 9 12 2 9 9 14 2 11 2 0 11
26 12 2 12 2 1 9 12 2 12 2 2 11 2 11 12 2 12 2 12 2 12 2 11 13 2 2
2 11 2
14 11 12 2 12 1 9 2 2 2 12 2 12 2 2
15 9 11 2 11 12 2 12 2 12 2 12 2 2 3 2
2 11 2
59 9 11 2 12 2 9 2 11 2 11 12 2 12 2 12 2 12 2 11 2 11 12 2 12 2 12 2 12 2 11 2 11 12 2 12 2 12 2 12 2 12 2 12 2 11 2 11 12 2 12 2 12 2 12 2 12 2 12 2
36 11 2 12 2 9 2 11 2 11 12 2 12 2 12 2 12 2 2 12 2 12 2 12 2 12 2 2 12 2 12 2 12 2 12 2 2
29 9 2 11 2 11 12 2 12 2 12 2 12 2 12 2 12 2 2 11 2 11 12 2 12 2 12 2 12 2
32 11 2 9 2 11 2 11 12 2 12 2 12 2 12 2 11 2 11 2 11 12 2 12 2 12 2 12 2 12 2 12 2
17 11 2 9 2 11 2 11 2 11 12 2 12 2 12 2 12 2
31 11 2 9 2 11 2 11 12 2 12 2 12 2 12 2 12 2 12 2 11 2 1 11 12 2 12 2 12 2 12 2
14 9 9 9 1 11 2 0 9 2 11 12 2 12 2
51 9 11 9 1 0 11 2 9 7 2 11 2 0 11 12 2 12 2 0 9 2 2 11 12 2 12 2 9 9 2 11 2 11 12 2 12 2 11 2 11 12 2 12 2 11 2 11 12 2 12 2
20 9 9 1 11 2 9 2 0 9 2 12 5 12 9 2 11 12 2 12 2
19 9 2 11 2 12 2 0 9 2 1 11 2 11 2 2 12 2 12 2
5 11 12 2 12 2
7 11 2 12 11 2 12 2
3 9 0 9
2 11 2
18 0 9 11 11 13 3 0 9 9 1 9 1 9 9 1 0 9 2
24 0 11 13 3 10 9 1 0 9 2 1 15 13 1 10 9 11 11 10 0 9 1 9 2
16 4 13 3 1 9 2 3 9 13 0 9 9 1 9 9 2
2 0 9
2 11 2
13 9 0 9 11 11 15 13 3 13 9 11 11 2
16 0 9 13 13 3 12 0 9 1 11 1 0 9 1 11 2
16 11 15 1 12 9 13 1 9 1 9 1 11 1 9 12 2
18 0 9 0 9 1 0 9 7 13 9 1 10 9 7 11 15 13 2
2 11 13
2 11 2
13 0 0 9 0 9 11 11 13 9 1 0 9 2
28 0 9 2 15 1 9 1 11 13 0 7 0 9 2 13 2 16 15 13 13 9 2 9 1 9 7 9 2
6 11 11 13 13 1 11
2 11 2
4 9 13 1 9
9 11 11 13 0 2 16 13 1 9
2 9 9
32 1 0 9 0 15 3 13 9 12 10 9 11 11 7 11 11 1 11 1 11 1 11 1 11 2 3 13 9 0 9 13 2
23 3 1 0 7 1 9 13 13 9 7 9 9 11 11 7 3 13 2 16 9 13 9 2
6 11 11 2 11 1 11
22 1 9 9 0 9 13 13 1 9 11 9 9 1 9 0 2 0 9 1 0 9 2
41 1 0 9 9 1 9 1 11 1 9 1 11 1 11 13 3 11 1 11 13 1 9 0 9 0 9 11 11 2 15 13 1 0 11 7 13 2 9 2 13 2
17 16 13 1 9 2 13 2 2 13 0 2 16 13 1 9 2 2
23 0 11 3 4 1 10 9 13 0 9 11 11 1 11 7 3 13 1 0 2 0 9 2
7 13 3 3 0 9 9 2
24 0 9 11 15 3 3 3 13 0 9 2 7 3 15 3 13 13 9 1 9 1 0 9 2
28 16 15 11 11 1 11 11 13 1 9 3 1 11 2 3 13 1 9 0 11 11 2 13 1 9 0 9 2
19 9 15 13 1 9 2 9 9 13 7 13 3 9 2 16 15 9 13 2
16 0 9 9 1 11 15 13 0 9 9 11 11 7 11 9 2
18 3 0 9 9 11 11 13 3 10 0 9 2 16 15 1 9 13 2
27 3 4 15 3 13 2 9 9 4 13 3 1 9 0 9 12 2 9 9 14 11 1 11 9 1 9 2
16 16 9 13 2 13 15 9 1 9 13 1 9 3 3 3 2
34 0 9 11 11 11 2 13 0 9 1 11 2 7 11 11 2 11 0 2 11 2 15 3 13 1 11 1 11 1 9 11 2 11 2
23 11 2 15 1 11 1 11 1 9 1 11 13 2 13 13 1 9 2 14 2 11 2 2
23 11 15 13 2 16 1 9 3 13 0 0 9 2 7 1 10 9 1 0 9 13 9 2
15 9 3 13 0 9 7 13 13 2 16 1 9 13 9 2
13 11 11 13 1 9 9 10 9 1 9 0 9 2
13 10 0 9 4 15 13 1 0 9 13 11 11 2
12 3 11 11 13 1 0 9 2 3 1 11 2
13 0 0 9 13 9 1 0 11 7 9 14 13 2
12 1 10 9 13 9 3 9 11 11 11 11 2
9 2 3 13 13 2 2 13 11 2
15 1 9 0 9 13 1 11 1 11 0 9 1 0 9 2
26 1 11 11 7 0 9 11 7 11 1 15 13 7 0 9 0 9 7 9 9 1 11 12 11 9 2
30 0 9 11 11 2 12 2 2 15 1 9 13 1 11 1 0 9 11 2 13 1 0 9 9 0 9 1 0 9 2
17 1 10 9 15 3 13 1 9 9 11 2 15 15 13 1 9 2
24 0 9 13 11 2 9 9 2 1 11 11 2 9 11 11 11 2 11 11 2 7 0 11 2
4 0 9 15 2
12 4 13 1 9 3 1 11 11 7 11 11 2
17 13 15 3 0 9 9 9 7 11 2 15 3 3 3 13 3 2
4 11 1 9 9
2 11 2
33 9 0 9 0 9 11 11 3 13 2 16 4 15 0 2 9 9 0 1 0 0 9 11 7 11 13 9 1 9 12 1 11 2
41 1 9 1 9 11 11 11 11 3 13 9 10 9 2 2 11 11 4 13 2 16 16 13 1 9 11 1 9 2 9 0 1 0 0 9 15 0 9 13 2 2
3 0 9 11
2 11 2
11 0 9 9 13 3 1 9 7 12 9 2
18 1 15 0 11 13 0 9 14 1 12 2 9 2 3 15 13 11 2
12 11 1 10 9 3 3 13 14 1 0 12 2
17 1 0 9 13 0 9 0 9 11 2 16 11 13 1 0 9 2
20 1 0 9 9 9 15 11 1 10 0 9 3 13 2 7 16 13 0 9 2
16 3 1 0 12 13 7 1 9 0 13 1 12 9 12 9 2
3 9 1 9
2 11 2
17 11 11 1 11 13 1 11 0 9 9 1 0 9 1 0 9 2
8 2 13 15 10 0 9 3 2
25 13 4 0 9 1 9 11 1 9 11 7 9 9 13 1 0 9 2 2 13 0 11 2 11 2
25 1 9 4 3 13 9 1 9 9 1 11 2 15 15 4 13 1 9 12 2 2 12 2 9 2
16 9 2 11 2 11 2 11 2 11 7 11 2 11 11 2 2
3 9 11 2
1 9
12 9 2 9 0 9 9 1 0 11 4 13 2
11 1 9 1 9 13 9 1 15 0 9 2
14 0 2 0 2 3 0 9 12 7 12 9 5 9 2
19 1 9 13 9 0 9 2 3 1 9 2 15 4 1 9 13 1 0 2
19 0 9 12 7 12 9 2 9 2 0 0 9 12 7 12 9 2 9 2
30 1 9 13 3 3 2 3 9 2 0 9 9 12 7 9 12 9 2 9 2 0 0 9 12 7 12 9 2 9 2
20 1 9 13 9 1 12 7 13 1 12 2 9 13 1 12 7 13 1 12 2
26 0 9 12 2 9 2 0 9 12 9 2 9 1 9 12 2 0 9 12 9 2 9 1 9 12 2
9 0 0 9 13 12 9 2 9 2
21 1 9 0 9 13 13 0 9 9 12 0 9 2 15 13 12 9 1 0 9 2
18 0 9 1 0 9 1 9 13 3 7 3 0 2 1 9 3 0 2
15 2 11 2 0 9 9 13 3 0 2 0 9 9 0 2
3 2 11 2
6 12 9 1 9 7 9
9 11 4 13 7 13 4 1 9 3
5 11 2 11 2 2
24 9 0 9 11 13 1 0 9 12 2 7 12 2 9 9 12 9 15 13 1 0 0 9 2
10 9 0 9 4 13 15 0 0 9 2
17 1 12 0 9 1 9 12 14 3 4 0 9 13 9 1 9 2
15 1 9 12 2 12 4 15 1 9 13 11 2 7 11 2
27 0 1 0 0 9 13 12 9 1 12 9 7 12 9 2 11 13 9 12 1 12 9 7 12 0 9 2
22 13 12 9 1 9 3 3 2 13 15 11 1 12 9 2 11 4 13 1 9 3 2
10 3 4 0 9 13 1 9 1 9 2
8 3 4 13 11 1 9 12 2
27 3 13 1 9 9 1 0 0 9 1 11 2 3 4 13 1 9 3 16 0 9 7 13 4 1 9 2
15 9 4 13 3 13 1 0 9 11 1 9 12 2 12 2
42 9 1 11 3 13 1 12 9 1 12 2 9 2 1 0 9 4 13 0 2 12 9 2 7 1 15 4 13 11 2 12 2 7 11 2 12 2 0 0 9 2 2
56 0 9 13 3 0 9 2 1 9 12 2 12 4 11 1 0 9 13 11 2 7 11 2 11 2 1 9 12 4 0 11 13 9 9 11 2 7 9 11 7 1 0 0 9 2 12 2 12 2 4 1 11 13 11 11 2
12 3 0 9 4 13 0 9 0 9 0 9 2
17 11 1 12 9 4 13 1 11 2 12 2 7 11 2 12 2 2
33 9 4 15 13 14 3 2 11 4 15 13 9 1 11 2 12 2 1 12 2 2 7 11 1 9 2 12 2 1 12 2 2 2
4 11 1 0 9
6 9 11 13 11 15 13
2 9 9
5 11 2 11 2 2
38 2 11 15 14 3 13 2 16 4 15 3 13 12 9 2 2 13 1 9 9 11 2 11 2 9 9 11 2 15 3 13 9 1 9 7 1 9 2
61 1 9 9 1 9 1 11 11 13 3 1 9 9 11 2 15 9 1 9 13 3 11 2 7 1 9 9 11 15 15 13 1 11 1 9 3 1 12 9 1 9 1 11 2 0 9 3 1 9 1 12 9 2 13 15 1 12 0 9 2 2
28 12 9 13 1 0 9 9 14 3 2 11 13 13 3 14 1 0 9 2 3 15 13 9 1 9 11 2 2
40 0 9 13 14 3 1 9 0 9 11 2 15 1 0 9 9 1 9 12 2 9 11 2 11 2 12 2 12 2 13 0 9 2 15 11 13 12 2 12 2
21 1 10 9 16 4 0 11 1 9 13 9 2 1 15 0 13 1 11 1 9 2
27 9 13 13 1 0 9 11 7 9 11 2 15 1 9 9 2 9 9 1 9 2 13 9 3 13 9 2
4 0 9 1 11
8 11 13 1 0 2 11 0 9
2 11 2
23 0 9 0 9 15 14 1 0 0 9 11 2 11 13 0 3 7 11 13 3 12 9 2
11 0 9 7 13 9 0 11 1 0 11 2
17 9 13 13 3 1 9 7 9 1 0 9 13 1 12 9 9 2
13 0 2 11 4 13 0 9 0 9 11 7 11 2
6 7 11 15 13 0 2
20 1 9 4 13 11 7 1 15 2 16 13 9 2 13 9 14 1 0 9 2
15 1 9 13 11 2 0 11 4 13 3 13 14 1 9 2
9 1 9 11 13 9 12 0 9 2
20 11 15 3 1 9 13 1 11 12 9 2 7 11 1 9 9 11 3 13 2
6 0 4 13 0 11 2
26 1 0 9 1 11 7 0 1 11 15 13 11 11 13 1 11 2 15 4 13 0 9 2 9 11 2
19 11 13 11 3 1 11 2 11 7 11 2 1 15 13 0 9 7 11 2
7 11 4 13 3 0 11 2
21 9 2 15 15 1 9 1 9 13 9 9 12 9 2 13 11 3 1 0 9 2
11 1 9 9 15 3 1 0 9 13 11 2
29 11 13 1 9 1 11 3 0 9 13 15 9 1 9 2 13 15 7 4 11 2 9 2 7 11 2 9 2 2
10 9 3 3 13 0 9 11 1 11 2
24 1 9 0 4 0 13 7 0 9 11 2 11 7 11 2 7 3 3 13 9 9 1 9 2
23 9 4 1 3 0 11 2 11 7 11 2 11 13 7 0 9 11 2 12 0 9 2 2
52 9 12 2 9 2 9 2 12 2 11 2 11 2 9 12 2 11 2 11 2 12 2 11 2 11 2 0 2 11 2 11 2 9 2 11 2 11 2 11 11 2 2 11 2 11 2 12 2 11 2 11 2
18 13 1 11 2 0 9 9 2 9 10 9 11 11 1 9 9 1 9
5 1 0 9 11 11
4 9 13 9 2
4 9 13 9 2
6 9 13 1 0 9 2
5 9 9 13 9 2
4 9 9 13 2
5 13 2 16 13 2
5 1 9 7 9 2
5 13 14 10 9 2
5 0 9 0 9 2
9 9 3 1 15 13 1 0 9 2
7 0 9 13 3 0 9 2
14 15 15 13 2 16 4 13 2 15 10 0 9 13 2
18 16 4 15 13 9 2 13 4 15 0 7 15 4 13 13 3 3 2
8 16 4 15 13 9 2 3 2
11 7 0 9 1 9 13 2 3 0 9 2
7 15 13 2 15 13 15 2
20 7 3 1 12 0 9 1 9 0 9 0 9 9 13 2 9 1 9 2 2
8 1 9 9 2 9 2 9 2
24 9 2 1 0 9 2 13 3 0 9 1 0 9 2 0 9 9 7 9 9 1 0 9 2
9 9 1 15 13 1 0 0 9 2
31 7 3 0 9 13 9 9 2 10 0 9 7 9 0 9 1 9 13 9 1 0 9 9 13 10 9 3 1 10 9 2
9 7 1 9 13 9 1 0 9 2
27 3 0 13 1 9 1 0 9 9 9 7 9 2 15 15 1 0 9 9 9 3 13 7 13 9 0 2
7 7 1 15 13 0 9 2
33 0 3 0 9 3 13 10 9 3 3 3 3 7 15 0 3 13 2 16 13 3 13 0 9 2 7 15 13 0 9 0 9 2
13 9 13 1 3 0 9 3 0 9 0 9 9 2
15 9 1 9 10 0 9 3 0 9 0 9 7 0 9 2
16 0 9 13 3 7 0 9 1 15 2 15 13 15 0 9 2
18 3 15 1 15 9 1 3 15 9 0 9 15 3 0 9 3 13 2
22 3 3 3 1 15 13 12 9 2 15 15 15 3 13 7 13 2 0 7 0 9 2
28 3 15 1 11 3 3 13 1 15 9 9 13 1 15 2 15 13 3 1 10 10 9 9 0 9 2 2 2
7 9 13 9 3 1 9 2
4 9 16 0 9
5 11 2 11 2 2
22 9 2 16 9 13 2 0 9 2 2 13 1 0 9 9 1 9 9 7 0 9 2
17 10 9 13 3 13 10 9 1 10 9 2 16 13 0 13 15 2
10 13 7 14 3 13 2 15 15 13 2
35 9 1 9 0 9 9 2 9 0 2 9 9 2 7 9 2 9 2 13 9 1 9 9 7 0 9 1 12 2 0 9 11 1 11 2
20 13 1 15 1 0 9 2 15 3 13 13 1 0 9 7 3 13 10 9 2
39 1 9 0 9 2 1 15 0 4 1 9 13 2 15 9 1 9 9 7 0 9 13 2 16 10 9 1 9 13 10 0 9 2 1 15 10 9 13 2
21 2 1 3 0 13 2 16 4 1 15 13 3 9 2 2 13 11 11 1 9 2
9 10 9 1 15 13 1 9 13 2
28 2 13 3 13 1 15 2 15 9 10 3 0 9 13 2 16 15 13 1 10 9 2 2 13 11 2 11 2
24 10 10 9 15 1 15 13 1 0 9 9 14 1 3 0 9 2 7 0 9 15 13 13 2
25 9 9 15 13 3 1 15 2 16 9 0 9 9 9 3 13 0 7 0 7 13 0 15 13 2
5 0 9 13 0 9
6 0 11 2 11 2 2
27 12 9 2 9 2 12 0 9 7 0 9 9 13 9 0 9 9 0 9 1 9 12 0 9 1 11 2
23 15 2 3 1 9 13 2 3 13 10 9 1 0 9 1 11 1 9 13 15 1 9 2
58 1 0 0 9 1 9 9 1 11 2 15 13 9 0 9 2 13 9 12 9 2 12 0 9 2 0 9 2 9 2 12 9 2 12 9 2 12 9 2 12 9 2 14 12 9 9 7 0 9 9 1 9 2 15 1 0 9 2
32 13 15 3 1 0 9 2 15 13 2 3 9 13 2 1 0 9 0 0 9 2 1 15 13 7 9 9 2 15 3 13 2
24 9 1 11 10 10 9 1 10 2 9 2 3 13 2 16 4 13 15 0 1 10 0 9 2
28 12 13 13 1 0 9 0 9 2 0 0 13 3 1 9 2 0 4 13 7 9 1 9 1 9 4 13 2
16 1 9 2 15 4 13 2 13 9 9 1 10 9 1 9 2
5 11 2 11 2 2
22 0 9 0 9 9 11 7 9 11 11 11 3 4 13 2 16 9 3 13 0 9 2
12 11 15 13 9 9 9 9 11 11 2 11 2
29 1 11 2 11 13 0 9 0 9 9 11 1 15 2 16 13 9 0 9 7 0 0 9 1 9 12 9 9 2
9 15 9 13 9 0 10 0 9 2
12 1 10 9 4 1 11 2 11 13 0 9 2
14 13 15 7 9 2 16 11 2 11 15 13 1 9 2
6 15 13 12 2 9 2
3 10 9 2
2 9 9
2 11 11
36 0 9 13 1 9 9 9 2 7 1 15 13 15 3 10 0 9 2 15 13 7 13 14 9 2 7 16 15 13 2 3 13 15 0 9 2
17 13 15 9 9 12 2 9 1 12 0 9 1 11 1 11 12 2
19 12 9 3 3 3 13 1 9 9 11 11 2 15 13 0 9 2 2 2
35 13 7 9 2 16 13 1 2 10 9 2 3 15 3 13 7 13 2 2 7 1 10 9 9 7 9 2 3 2 13 10 0 9 2 2
63 3 9 15 13 2 16 0 9 13 9 9 7 9 9 2 3 13 2 13 9 2 13 9 2 13 9 7 9 2 2 9 9 2 9 2 3 2 13 3 9 2 2 3 15 13 1 9 1 9 1 9 7 13 15 2 0 9 2 1 9 7 9 2
27 12 9 13 1 15 2 16 0 9 13 9 1 9 2 15 2 13 7 0 9 7 0 0 0 9 2 2
42 11 11 13 7 15 2 16 1 0 9 2 15 1 9 13 1 9 2 13 15 1 9 9 2 7 13 9 2 15 15 0 13 2 7 7 13 1 0 9 1 9 2
15 2 7 3 3 10 9 13 9 2 2 13 15 11 11 2
21 1 9 2 1 9 0 9 0 0 9 1 0 9 2 1 9 9 15 13 15 2
28 14 1 12 9 2 15 15 10 9 3 13 2 16 10 9 2 13 9 2 2 16 2 13 15 10 9 2 2
4 0 11 13 9
2 9 9
11 9 0 11 13 3 0 9 1 0 9 2
14 13 7 0 13 0 9 7 2 13 2 15 0 9 2
24 15 13 9 0 9 9 3 12 9 0 9 7 9 2 15 15 13 1 11 2 11 7 11 2
2 11 11
7 9 13 3 10 0 9 2
23 0 9 2 0 9 9 1 0 9 2 13 9 1 0 9 11 1 9 12 9 1 11 2
27 1 15 12 9 15 3 13 7 0 9 1 9 7 9 1 9 7 9 9 7 1 0 9 1 0 9 2
28 0 9 11 9 3 13 1 0 9 0 11 1 9 1 9 0 9 2 3 0 9 2 9 9 7 0 9 2
11 9 15 13 0 9 1 11 7 1 11 2
22 11 15 3 13 9 1 9 0 9 1 0 9 0 11 1 9 1 12 9 2 9 2
23 3 13 11 1 11 9 7 9 1 0 9 12 9 2 9 2 1 9 13 1 0 9 2
10 0 9 13 1 9 0 9 1 11 2
30 0 2 9 2 11 3 13 9 1 9 1 0 9 11 7 13 7 0 9 1 9 9 1 9 7 0 9 1 11 2
14 4 13 3 9 1 9 12 9 1 0 9 0 11 2
15 9 9 2 0 3 1 9 12 2 3 13 0 0 9 2
12 0 9 11 13 1 11 9 1 0 0 9 2
11 9 1 10 9 7 13 3 0 0 9 2
21 1 0 0 9 12 9 2 1 15 15 13 12 9 2 13 11 9 1 12 9 2
23 1 11 13 11 0 9 3 1 9 2 9 11 1 11 3 13 3 12 9 2 3 1 12
3 9 1 9
11 9 11 9 1 9 11 11 1 9 9 2
5 9 11 11 2 11
6 9 0 1 9 1 9
13 0 9 9 0 13 3 0 16 9 1 0 9 2
22 9 11 11 2 0 10 0 9 0 9 2 13 1 9 2 16 9 13 3 10 9 2
10 7 13 2 16 0 9 9 3 13 2
22 2 16 15 11 13 9 7 13 0 13 10 0 9 2 13 3 9 9 2 2 13 2
51 9 11 11 11 1 0 9 1 9 9 1 10 9 9 0 9 1 9 3 13 9 9 7 13 2 16 9 0 9 13 9 1 12 12 9 0 9 0 9 1 9 0 9 2 7 15 15 15 13 13 2
4 13 0 9 2
22 10 9 13 13 9 9 2 15 15 13 2 13 15 7 3 13 9 9 2 13 11 2
28 16 13 1 9 2 13 2 16 13 1 9 0 9 2 3 16 13 1 9 0 9 2 1 15 15 13 9 2
16 13 3 9 9 1 0 9 2 15 15 1 9 9 9 13 2
14 13 2 16 9 13 9 1 0 0 7 0 0 11 2
23 0 9 3 13 2 16 1 9 0 0 9 0 0 9 9 2 11 2 13 0 9 9 2
31 3 13 9 11 11 2 9 11 11 2 12 1 9 11 2 13 1 12 9 0 1 9 2 15 13 1 9 1 9 13 2
7 0 9 13 9 0 9 2
19 1 9 1 9 11 1 0 11 4 13 0 9 2 9 7 0 9 9 2
24 1 9 13 0 9 12 2 9 12 9 9 12 2 1 9 0 9 2 0 0 9 11 12 2
4 11 13 9 9
4 11 13 9 9
41 0 9 0 9 1 0 9 2 11 2 2 1 15 13 1 11 3 11 2 11 7 11 2 15 3 1 11 13 1 9 9 0 9 9 1 12 2 9 0 9 2
4 11 9 2 11
39 1 0 9 2 15 1 0 9 0 9 11 13 9 9 2 13 1 12 2 9 13 9 3 1 12 12 1 3 0 9 7 1 12 12 1 3 0 9 2
17 3 15 13 9 0 9 1 9 1 9 1 11 2 11 7 11 2
19 1 0 9 0 9 15 3 4 1 9 11 13 3 1 9 0 9 3 2
12 0 9 13 13 3 1 9 9 1 0 9 2
23 9 13 1 12 2 9 12 9 1 0 9 14 1 10 9 1 3 0 9 13 1 9 2
16 3 1 0 9 0 9 13 13 9 14 1 9 12 7 12 2
17 1 9 1 9 9 11 3 1 9 1 11 13 1 0 9 9 2
13 1 9 9 13 0 9 1 0 1 9 0 9 2
27 3 1 9 9 13 0 9 9 7 9 11 11 2 0 9 9 1 9 1 12 9 9 4 13 9 9 2
34 0 9 9 11 11 1 9 1 9 11 13 2 16 15 9 9 1 12 2 9 12 13 13 2 7 7 1 10 9 4 13 9 9 2
11 1 0 9 1 15 13 7 1 9 12 2
17 11 4 13 1 9 12 1 11 7 13 13 1 12 2 9 12 2
38 1 0 9 3 1 9 13 13 13 0 9 1 9 0 9 9 1 10 9 1 0 12 1 12 9 2 3 1 12 2 9 12 2 1 0 9 12 2
15 1 0 9 4 3 13 10 9 9 2 9 7 0 9 2
13 1 9 1 11 7 11 1 15 13 3 9 11 2
3 13 1 15
10 0 9 13 1 0 9 1 10 9 2
46 1 9 15 3 3 13 0 9 1 0 11 2 16 1 9 3 13 0 9 1 9 0 9 7 1 0 9 15 13 7 9 1 11 1 11 7 1 11 2 3 15 13 0 0 9 2
52 9 1 0 0 9 9 13 1 0 9 1 11 0 9 0 9 2 15 15 13 1 0 0 9 2 3 15 3 2 13 11 11 2 11 2 2 9 9 2 11 2 2 11 2 11 2 7 9 2 11 2 2
9 1 15 9 15 13 1 12 9 2
3 2 11 2
3 9 1 9
2 9 2
20 9 7 2 11 2 12 9 2 2 11 2 11 2 12 2 11 2 0 11 2
21 1 0 9 9 9 15 11 1 10 0 9 3 13 2 7 16 0 9 13 15 2
16 3 1 0 12 13 7 1 9 0 13 1 12 9 12 9 2
21 1 9 7 0 9 11 3 13 0 9 7 13 14 1 9 11 1 12 2 9 2
7 3 7 11 1 9 13 2
17 9 2 11 2 11 2 2 2 11 2 11 2 12 11 2 2 2
6 9 2 12 2 12 2
6 9 2 12 2 12 2
7 1 9 2 12 2 12 2
4 9 2 12 2
14 12 2 12 2 12 2 12 2 12 2 12 2 12 2
2 1 9
2 11 11
21 3 2 7 3 2 13 4 15 13 3 2 16 0 9 13 9 9 1 0 9 2
29 15 2 1 3 12 9 0 9 7 0 0 9 2 13 9 2 16 4 11 13 13 9 2 1 15 15 13 9 2
27 9 2 15 3 0 9 9 1 0 0 9 0 9 13 2 13 7 10 9 2 16 1 9 13 0 9 2
14 1 0 9 13 13 3 14 9 2 16 9 3 13 2
14 10 9 13 0 9 3 9 2 10 9 13 0 9 2
38 16 11 2 1 10 9 13 0 9 0 15 3 9 3 2 3 0 9 2 7 9 9 9 1 9 13 9 9 1 9 2 1 9 11 13 15 0 2
18 9 9 9 11 11 13 1 0 9 2 15 0 0 9 9 9 13 2
28 1 0 4 13 9 2 16 9 13 9 14 1 9 2 15 13 1 9 1 0 2 3 7 0 7 0 9 2
28 10 9 13 1 9 1 0 9 3 0 7 1 9 9 13 13 14 9 0 2 7 7 13 9 1 0 9 2
21 3 2 13 15 1 9 0 9 1 9 0 1 0 9 1 0 9 13 1 9 2
35 2 0 9 13 13 3 16 9 1 0 9 2 2 13 1 10 9 9 11 11 11 2 12 1 10 9 11 2 15 1 0 9 13 9 2
32 9 15 3 3 13 1 9 2 16 3 13 1 9 0 9 2 15 3 7 3 13 0 9 7 13 16 12 1 9 1 9 2
8 7 3 15 13 9 1 9 2
6 13 15 7 9 0 2
23 9 2 7 13 13 16 7 9 11 2 2 0 1 0 9 2 15 13 13 1 0 9 2
18 10 9 4 13 4 13 0 9 16 0 9 1 9 0 9 9 12 2
16 3 15 13 2 1 9 11 11 11 2 9 9 1 0 9 2
14 0 0 9 0 9 15 1 0 9 13 13 16 9 2
27 14 1 9 9 2 7 16 9 9 9 2 15 13 1 9 9 9 0 13 0 9 7 0 9 0 9 2
6 11 2 9 1 9 9
5 11 2 11 2 2
26 0 9 9 2 16 15 9 13 9 0 13 9 9 2 2 13 10 9 0 9 9 1 0 9 2 2
15 9 11 15 3 13 9 9 11 11 2 11 2 11 2 2
20 0 9 9 0 9 12 2 9 1 15 13 9 2 15 9 9 0 9 13 2
34 11 13 2 16 9 11 11 13 1 9 9 9 2 1 15 9 9 3 0 13 4 13 3 7 9 1 0 9 1 9 9 1 9 2
17 3 1 0 0 9 1 0 9 3 1 15 13 0 9 0 9 2
16 2 13 3 9 9 2 9 7 0 2 0 9 2 2 13 2
27 1 9 9 11 2 11 13 3 9 11 2 11 9 9 2 9 7 9 0 0 9 11 11 2 11 2 2
5 9 11 11 2 11
7 9 1 11 13 0 0 9
2 11 2
20 11 7 11 3 1 11 3 13 10 9 1 9 0 9 11 11 0 0 9 2
13 11 13 11 1 9 9 0 0 9 1 9 12 2
28 11 3 13 11 1 3 0 9 2 9 0 9 9 0 9 1 0 9 9 7 1 9 0 9 1 0 9 2
14 9 4 3 13 2 16 9 1 9 12 13 3 0 2
17 1 0 9 15 12 9 13 3 2 16 15 9 13 1 0 9 2
13 0 0 9 13 3 0 9 9 0 9 0 9 2
31 9 9 3 1 10 9 0 0 9 13 14 15 2 16 15 13 1 0 9 7 16 1 9 9 12 9 3 13 12 9 2
11 11 7 11 13 2 16 15 9 9 13 2
18 13 7 1 9 3 0 2 3 15 15 13 10 9 7 9 9 9 2
12 0 0 9 15 1 15 13 3 1 9 12 2
5 11 13 9 1 9
2 11 2
33 0 9 9 11 11 3 13 2 16 4 11 13 9 0 2 0 9 1 11 7 11 1 3 0 9 9 1 9 10 0 0 9 2
32 10 9 13 9 2 16 1 9 15 13 0 9 7 0 9 7 16 10 9 4 15 13 13 9 0 9 1 0 11 7 9 2
23 1 9 15 13 9 0 11 2 15 15 1 9 11 13 1 0 9 0 9 1 9 11 2
8 3 1 0 11 1 9 12 2
5 11 15 13 0 9
38 1 11 9 2 0 9 1 9 1 11 2 15 13 1 0 9 0 2 0 9 13 1 0 9 2 13 3 0 0 9 2 16 4 15 13 0 9 2
13 1 0 15 9 9 9 1 9 1 0 9 13 2
2 9 11
6 9 11 13 9 0 9
5 11 2 11 2 2
11 1 9 1 9 13 9 11 12 9 9 2
16 1 9 15 13 9 11 2 15 13 10 9 0 0 9 11 2
21 0 9 0 9 1 10 0 9 13 12 9 2 9 2 11 7 13 3 12 9 2
16 1 0 9 0 9 9 11 15 3 13 0 9 11 11 11 2
30 1 10 9 9 9 9 13 11 1 9 9 0 0 11 2 3 10 9 13 0 9 11 11 11 1 9 0 9 11 2
23 10 9 13 3 2 1 10 0 9 9 11 7 11 15 13 7 0 0 9 1 9 11 2
31 9 0 9 11 11 11 2 15 13 1 0 9 1 9 0 9 2 3 13 2 16 11 2 13 1 0 9 7 9 2 2
18 1 11 2 11 0 9 9 11 13 1 9 0 9 9 0 0 9 2
22 3 3 13 0 9 9 11 11 2 13 0 9 0 9 1 0 9 11 9 11 13 2
17 11 3 13 11 1 15 2 16 0 9 11 1 0 9 3 13 2
25 16 9 13 0 9 2 15 1 9 0 9 3 13 10 9 1 11 1 9 3 12 9 2 9 2
14 9 0 9 11 11 15 10 9 7 13 2 7 13 2
23 11 11 3 13 9 1 15 2 16 1 9 0 9 1 9 11 2 11 4 3 13 9 2
20 1 9 2 15 13 11 1 9 2 9 3 13 9 7 9 3 4 13 9 2
19 3 4 3 1 11 13 2 4 13 9 11 13 10 9 1 0 0 9 2
8 0 9 13 11 3 1 9 2
16 11 11 3 3 9 11 1 0 0 9 1 0 9 3 13 2
31 1 9 1 9 10 9 1 9 12 1 9 1 9 11 13 2 16 13 3 13 0 9 2 15 0 0 9 1 9 13 2
19 9 11 1 9 3 13 2 16 3 13 9 1 9 1 0 0 0 9 2
19 13 3 2 16 3 1 0 9 13 1 0 9 9 0 9 1 0 9 2
35 2 13 15 3 10 9 2 13 4 13 1 9 2 2 13 11 12 9 1 15 2 16 1 0 9 13 9 16 0 0 9 1 9 11 2
7 15 13 9 2 15 13 9
5 11 2 11 2 2
16 1 0 9 0 9 13 9 1 11 7 11 9 9 0 9 2
17 1 12 9 9 7 0 9 13 12 2 0 3 9 7 9 2 2
11 1 9 9 7 0 9 13 3 0 0 2
15 13 15 15 3 0 9 1 11 7 9 0 9 1 11 2
6 13 0 9 0 9 2
10 1 9 13 3 9 7 9 1 15 2
6 15 9 13 1 9 2
8 3 9 1 9 4 13 3 2
22 1 9 9 0 0 9 1 11 13 9 1 0 9 1 9 9 0 9 7 9 0 2
6 0 12 9 13 0 2
25 13 15 1 0 9 0 9 2 15 15 3 0 9 3 13 2 7 3 13 3 0 9 1 15 2
16 2 3 13 15 0 9 2 3 9 13 2 2 13 11 11 2
23 1 9 13 0 9 13 0 9 9 1 9 12 7 12 12 2 9 12 7 12 12 9 2
12 1 0 9 0 9 4 13 3 12 0 9 2
8 9 0 9 13 9 1 0 9
5 11 2 11 2 2
19 1 9 13 0 9 9 1 9 9 11 11 1 9 0 9 1 9 11 2
19 1 9 9 0 2 9 0 2 9 11 13 2 16 13 1 9 1 9 2
13 11 11 13 9 2 16 3 13 1 9 12 9 2
19 9 0 2 9 7 13 1 9 9 2 16 4 9 13 3 1 12 9 2
32 15 15 1 9 2 16 0 9 0 9 13 0 7 9 9 1 0 9 0 9 4 13 9 0 9 7 13 15 0 0 9 2
30 0 9 1 11 1 0 9 7 0 9 13 1 0 9 9 9 2 13 9 2 9 2 11 11 1 0 9 0 9 2
21 0 9 13 3 1 9 9 1 9 2 3 9 0 0 9 13 7 13 0 9 2
17 1 11 13 9 3 0 9 3 2 1 9 0 9 1 0 9 2
11 0 9 13 1 9 1 10 0 0 9 2
17 1 9 3 13 13 0 9 2 3 2 0 9 7 3 0 9 2
20 1 11 11 15 13 3 0 0 9 0 9 1 11 2 3 3 13 0 9 2
32 0 13 7 9 1 0 9 2 3 3 13 1 9 9 1 9 12 1 3 0 9 2 15 9 1 0 9 1 11 3 13 2
18 9 9 11 11 13 1 9 0 9 2 3 13 0 9 1 0 9 2
5 9 11 11 2 11
1 13
15 0 9 9 2 12 9 1 9 2 7 3 6 1 15 2
11 0 9 1 9 1 9 13 3 1 9 2
8 1 9 15 13 2 7 15 2
21 3 13 0 2 16 4 1 0 9 13 1 9 1 9 2 7 15 13 9 9 2
7 13 15 9 2 7 9 2
6 9 1 15 13 9 2
4 9 13 9 2
14 0 9 9 13 9 13 9 7 9 1 9 0 9 2
6 9 13 1 10 9 2
9 13 9 2 3 4 15 13 9 2
4 0 9 3 0
5 11 2 11 2 2
28 9 4 13 13 1 9 9 9 11 11 9 13 1 0 9 9 0 9 2 16 4 10 9 13 0 9 9 2
29 0 0 9 2 11 2 13 0 13 1 15 2 16 3 2 9 2 15 13 9 2 15 4 13 13 9 1 9 2
19 3 4 1 9 11 11 11 13 0 2 16 4 9 9 13 13 3 9 2
30 11 2 11 13 2 16 3 9 1 0 9 0 9 2 10 9 3 9 13 2 4 3 13 0 0 9 1 9 9 2
26 1 0 9 9 13 3 0 9 0 9 13 2 3 2 13 2 7 15 9 13 0 9 1 0 9 2
27 11 13 2 16 12 9 9 2 15 13 9 0 9 0 1 0 9 2 13 0 13 1 9 0 9 9 2
19 9 13 13 1 9 3 2 9 9 2 10 9 2 1 0 9 0 9 2
26 9 4 13 3 2 0 12 9 13 2 16 15 13 10 9 3 2 2 16 4 15 4 9 3 13 2
22 16 13 1 0 9 2 1 9 11 2 11 15 0 9 11 13 1 9 1 10 9 2
5 13 9 3 0 2
5 11 2 11 2 2
18 9 1 9 9 2 15 13 9 1 9 0 9 2 13 3 1 9 2
24 9 3 3 2 3 1 0 0 9 1 9 2 13 2 16 0 9 13 13 1 9 9 0 2
15 1 9 2 11 2 11 1 11 15 13 1 9 0 9 2
23 1 11 13 3 2 9 0 14 1 12 9 9 2 1 12 9 15 7 13 3 12 5 2
10 13 3 10 9 2 15 13 10 9 2
16 3 9 13 0 9 13 15 1 15 9 2 3 13 10 9 2
11 9 13 2 16 9 3 13 13 1 9 2
12 13 3 1 0 9 9 2 15 9 9 13 2
5 9 1 11 13 9
5 11 2 11 2 2
13 9 0 9 9 9 1 0 9 1 11 13 9 2
18 1 0 9 13 1 9 9 9 7 3 15 9 9 13 1 12 9 2
24 0 9 7 1 15 9 13 7 1 9 13 3 0 9 0 9 2 3 15 0 13 9 13 2
27 11 11 2 9 9 0 9 2 9 11 13 2 16 9 9 2 9 11 2 3 1 9 13 15 1 9 2
10 3 9 0 9 4 1 0 9 13 2
11 1 12 2 9 13 0 13 3 0 9 2
4 9 9 15 13
5 11 2 11 2 2
16 0 9 10 9 13 13 0 9 9 2 9 11 1 0 9 2
22 0 9 0 9 13 1 9 9 9 11 11 9 15 9 3 1 9 0 7 0 9 2
23 9 9 13 13 1 10 9 0 9 9 2 0 0 9 2 0 9 4 13 1 9 9 2
16 2 13 13 9 11 7 11 2 13 13 0 2 2 13 11 2
29 3 9 16 9 4 13 9 7 9 2 15 13 9 1 9 10 0 9 11 11 2 13 9 1 9 1 9 2 2
22 1 0 9 13 3 13 0 9 7 0 9 1 9 11 2 15 13 12 0 9 9 2
6 9 1 9 2 0 2
29 9 15 1 0 9 13 1 0 9 2 16 1 0 9 13 10 0 0 9 2 1 15 13 3 2 7 0 9 2
11 1 0 9 13 9 9 9 0 1 9 2
28 1 9 10 9 4 13 9 9 14 12 0 9 2 3 0 9 9 13 0 2 13 15 7 1 9 1 9 2
4 9 11 13 9
7 11 2 11 2 11 2 2
30 7 0 9 1 0 9 13 1 0 9 0 9 1 0 9 11 2 11 1 9 1 9 0 9 1 0 9 1 11 2
12 9 11 1 15 13 11 11 1 9 1 11 2
28 3 3 13 2 9 13 0 9 1 9 2 15 13 1 9 0 9 9 1 0 9 2 15 0 9 3 13 2
29 2 0 9 13 1 0 9 13 1 0 9 2 16 15 7 0 9 13 2 7 10 9 3 13 2 2 13 11 2
31 1 0 9 11 13 9 9 11 11 2 16 9 9 13 9 1 9 1 12 9 7 1 10 9 13 0 9 7 0 9 2
24 1 11 13 0 0 7 0 9 1 9 12 9 0 9 2 1 15 12 13 13 2 12 13 2
6 9 1 11 13 13 9
5 11 2 11 2 2
25 7 1 9 9 7 9 0 0 9 13 0 9 9 9 1 12 0 9 7 12 9 0 0 9 2
10 0 9 1 0 11 13 0 9 9 2
19 1 9 0 0 9 11 2 11 13 3 11 0 9 0 13 0 0 9 2
21 15 13 13 1 9 9 2 13 9 2 2 15 15 11 13 1 0 9 1 9 2
29 0 9 9 11 15 3 3 13 2 1 0 9 1 9 0 9 1 0 9 1 9 0 9 1 9 9 0 9 2
14 13 15 1 0 9 7 9 0 0 9 7 0 9 2
12 1 0 0 9 13 9 11 9 11 2 11 2
30 11 11 2 0 1 9 0 2 15 1 9 12 2 9 13 1 0 9 1 11 2 11 2 3 3 13 9 1 11 2
9 13 15 0 9 0 9 11 11 2
22 0 2 3 3 0 11 11 1 11 0 13 1 9 1 0 9 1 0 0 0 9 2
12 10 0 0 9 13 2 16 11 13 9 9 2
21 13 15 7 9 2 16 15 1 9 0 9 3 13 0 9 7 9 1 9 9 2
12 9 1 11 13 2 16 4 11 13 13 9 2
6 9 15 13 1 9 9
2 11 2
34 3 16 0 9 9 1 0 9 7 9 0 9 7 9 9 1 11 15 1 9 1 9 9 1 11 13 1 9 1 11 7 0 11 2
12 13 1 15 0 0 9 2 15 10 9 13 2
13 9 13 1 9 12 16 9 1 9 0 0 9 2
28 13 9 1 11 2 15 15 13 2 16 0 9 13 13 3 1 9 2 7 13 9 1 9 0 9 1 9 2
14 9 13 1 15 2 16 4 15 1 9 13 9 9 2
5 13 1 12 9 2
27 1 0 9 7 9 9 0 9 1 0 9 13 9 11 11 1 0 0 9 9 9 7 0 9 11 11 2
6 9 1 11 13 1 11
2 11 2
11 9 9 1 11 11 11 13 11 1 12 9
2 9 9
5 11 2 11 2 2
12 3 1 9 13 11 0 9 1 9 9 12 2
15 11 11 15 3 13 1 11 9 9 11 11 7 11 11 2
35 2 3 4 13 9 1 9 2 7 9 13 1 0 9 1 9 1 3 16 12 9 7 3 16 1 10 0 9 13 9 9 2 2 13 2
22 2 11 13 0 9 2 13 15 1 9 7 15 4 13 1 10 0 9 14 1 9 2
7 1 9 11 3 15 13 2
25 16 9 13 12 9 2 15 13 1 10 9 3 3 2 13 15 13 2 3 9 13 9 13 9 2
14 16 4 15 13 1 9 9 2 13 15 13 3 3 2
12 1 9 3 4 13 1 11 11 1 9 11 2
8 13 2 16 3 13 13 9 2
29 2 16 13 1 9 9 1 11 2 11 2 11 13 2 16 9 12 15 3 13 3 7 3 1 3 0 9 2 2
6 0 9 13 9 0 2
8 11 7 11 15 7 13 9 2
16 1 9 1 9 12 3 1 9 13 0 9 0 0 9 2 2
19 9 0 11 11 11 3 13 0 9 2 16 0 11 3 9 9 9 13 2
27 9 9 1 11 7 0 9 1 0 11 13 11 2 16 4 13 9 2 15 4 13 0 9 1 0 9 2
12 0 9 0 9 11 11 11 13 3 1 11 2
31 1 15 4 13 0 9 2 0 1 9 11 2 11 7 11 2 15 15 0 9 13 13 9 1 0 9 7 9 0 11 2
17 10 9 9 4 13 9 9 1 11 7 0 9 9 11 1 11 2
35 9 0 9 9 0 9 4 13 15 2 16 0 11 13 9 1 9 1 11 2 13 3 0 9 11 11 1 9 1 9 9 11 2 11 2
26 9 0 9 13 1 9 0 9 0 9 2 1 15 4 1 0 9 13 11 13 12 9 1 3 12 2
9 11 2 11 2 9 13 9 0 9
2 9 9
14 9 13 1 10 9 9 9 9 1 9 0 0 9 2
17 1 10 9 13 1 0 9 11 11 2 9 0 9 1 0 9 2
15 11 11 9 13 9 2 16 15 9 0 9 13 3 3 2
12 9 11 13 9 9 0 9 1 0 9 3 2
5 15 15 13 15 2
40 9 2 15 9 13 9 9 1 9 0 9 2 13 9 2 16 13 1 9 0 9 2 16 4 15 9 0 9 13 2 13 2 16 4 0 9 13 3 3 2
13 16 4 13 0 9 2 13 4 15 15 9 13 2
22 9 9 2 10 9 7 9 1 10 9 13 3 9 12 9 2 15 15 3 13 3 2
4 9 1 9 12
4 9 1 9 12
11 3 13 2 16 4 9 13 13 9 9 2
28 13 4 9 9 11 11 2 15 1 10 9 13 0 9 2 16 9 7 0 0 9 13 1 9 9 9 11 2
15 16 3 13 0 9 2 13 9 1 9 0 9 0 9 2
22 7 13 9 2 16 4 2 14 1 15 13 9 7 0 9 2 3 4 9 13 3 2
9 13 1 10 9 3 14 15 0 2
23 13 0 9 2 9 0 9 2 15 13 1 12 9 9 0 9 2 13 0 9 0 9 2
13 9 9 2 9 7 9 13 12 1 9 0 9 2
38 16 4 15 3 13 1 0 9 2 1 0 9 0 9 7 9 2 3 9 13 1 9 9 2 13 12 0 9 2 13 4 15 1 9 7 1 9 2
21 13 9 2 16 4 15 9 7 11 13 13 1 9 0 9 2 3 0 1 9 2
23 13 1 0 9 0 9 9 7 10 9 9 2 1 15 13 2 16 10 9 4 15 13 2
15 13 9 1 0 9 0 9 2 1 10 9 0 1 9 2
19 15 13 9 2 0 9 13 9 0 12 2 9 2 3 0 12 2 9 2
13 13 2 16 9 1 15 3 13 2 15 13 9 2
12 13 15 2 16 4 15 9 0 9 3 13 2
23 16 15 13 1 15 2 16 4 13 1 11 7 11 2 3 13 15 9 1 9 0 9 2
12 1 9 9 13 11 7 11 2 13 0 9 2
22 9 13 9 9 13 15 3 1 9 10 0 9 7 9 9 10 9 13 9 1 9 2
29 13 2 16 0 9 13 2 1 15 15 1 9 13 2 7 16 3 0 0 9 13 2 15 13 14 9 0 9 2
6 1 11 13 3 14 9
5 11 2 11 2 2
14 1 0 9 4 15 9 0 9 13 13 1 0 9 2
13 1 0 0 9 11 15 13 10 9 11 2 11 2
20 0 9 13 15 2 16 11 4 13 3 13 9 2 15 13 4 13 0 9 2
15 15 11 13 1 9 1 9 2 15 11 13 1 9 12 2
6 9 1 9 1 0 11
2 11 2
19 13 1 9 1 0 9 10 9 13 9 0 0 9 1 9 11 7 15 2
22 1 12 2 1 12 2 9 15 13 1 9 0 9 9 11 2 13 9 9 11 11 2
20 1 11 4 15 13 9 13 9 11 11 2 9 11 11 7 9 9 11 11 2
32 9 3 13 0 9 11 11 2 9 9 11 11 11 7 11 11 11 2 0 9 11 1 0 9 11 1 0 11 7 0 9 2
8 1 9 11 15 15 9 3 13
5 11 2 11 2 2
34 0 9 2 15 1 0 9 9 2 3 13 1 9 0 9 1 9 1 0 9 7 9 2 13 13 9 1 9 2 13 9 0 9 2
25 9 3 13 2 16 9 13 3 10 9 2 15 1 9 13 12 9 9 2 3 15 13 12 9 2
6 11 13 3 12 9 2
24 3 1 0 9 15 13 0 9 2 11 2 2 9 9 11 7 11 7 9 9 1 0 9 2
20 1 9 13 9 1 9 1 12 9 9 2 1 9 9 0 1 9 12 2 2
11 3 9 13 3 12 9 1 0 0 9 2
23 10 9 13 3 2 3 1 9 7 3 2 1 9 0 9 1 9 2 0 1 0 9 2
34 3 15 13 9 0 2 7 0 9 0 9 13 2 16 1 0 9 2 12 7 12 9 9 2 15 1 0 9 13 3 9 9 9 2
50 11 3 4 1 9 13 12 9 9 2 11 12 9 2 2 11 12 9 2 2 11 7 11 2 11 1 12 9 2 2 11 12 9 2 2 11 7 11 1 12 9 2 2 11 2 11 12 9 9 2
10 9 0 9 1 9 9 3 13 11 2
31 15 2 16 1 11 2 11 15 1 9 0 1 9 9 13 1 3 0 9 11 2 4 15 13 3 9 9 1 0 9 2
18 3 13 0 9 2 11 2 0 9 7 9 0 2 3 12 9 9 2
8 0 0 9 11 13 9 16 0
5 11 2 11 2 2
9 0 0 9 11 13 9 16 0 2
15 13 15 1 9 0 0 9 1 9 12 2 15 13 9 2
9 1 0 9 0 9 13 9 9 2
22 9 9 0 9 0 9 13 3 12 9 2 1 15 13 1 9 0 9 13 12 9 2
28 1 9 13 9 0 9 1 12 9 2 0 1 12 9 2 2 0 9 1 12 9 2 7 9 1 12 9 2
15 3 1 9 9 13 9 9 2 1 12 9 1 9 12 2
22 1 0 9 15 3 13 2 1 0 15 13 1 0 12 2 1 9 13 1 12 9 2
15 9 9 15 13 1 9 7 1 9 13 9 1 9 13 2
16 9 9 13 1 9 12 9 2 1 12 3 16 1 9 12 2
7 0 9 9 13 12 9 2
17 9 9 12 13 1 0 9 12 9 2 1 12 3 16 1 9 2
6 13 15 7 9 9 2
14 0 9 15 1 9 7 9 3 13 1 9 7 9 2
14 1 9 7 9 13 12 9 9 2 1 9 12 9 2
8 1 9 4 3 13 0 9 2
19 1 0 9 13 12 9 0 9 2 15 13 3 16 1 0 7 0 9 2
12 0 9 9 13 1 12 2 0 1 12 9 2
19 0 9 9 2 1 9 1 12 9 2 1 9 12 2 9 13 0 9 2
14 0 9 13 9 1 9 12 9 7 9 13 12 9 2
7 13 3 3 16 0 9 2
74 9 13 2 16 4 12 9 4 13 1 9 0 7 0 9 2 3 1 9 11 2 11 2 0 11 7 11 2 12 9 4 13 4 13 1 0 2 9 2 0 9 16 9 9 1 0 9 2 12 9 4 13 13 1 9 9 9 7 9 9 7 9 11 7 12 9 1 9 9 1 9 0 9 2
8 11 15 1 11 13 9 0 9
5 11 2 11 2 2
33 9 9 1 9 0 9 1 9 2 15 13 11 11 2 11 2 2 4 1 9 11 11 2 11 13 0 9 0 9 0 9 12 2
39 9 3 13 1 9 11 2 3 11 13 1 9 0 9 2 15 9 13 1 9 9 3 9 2 15 13 1 9 1 9 0 2 7 14 1 0 7 0 2
18 2 11 13 0 13 1 9 0 9 1 15 2 16 4 13 0 9 2
21 13 4 9 10 9 7 13 4 2 16 0 9 4 13 1 9 9 0 0 9 2
15 7 12 1 15 13 3 0 9 2 2 13 11 2 11 2
22 1 15 13 9 3 10 0 0 9 0 0 9 2 3 13 9 0 9 1 9 0 2
16 2 1 10 9 15 3 4 13 2 15 13 9 7 15 14 2
20 7 9 15 4 13 15 2 15 4 13 3 1 0 9 2 2 13 9 11 2
18 1 15 15 3 13 9 0 9 2 15 13 1 0 9 3 9 11 2
3 9 1 9
5 11 11 2 11 11
15 9 11 11 15 3 13 1 0 9 11 2 11 7 11 2
12 1 12 9 13 10 9 3 9 9 11 11 2
27 13 2 14 9 9 9 11 11 1 11 1 9 9 2 13 10 0 9 1 0 9 3 12 3 0 9 2
17 13 15 3 2 16 9 13 1 0 13 9 10 9 9 1 9 2
7 15 13 9 10 0 9 2
15 11 11 13 1 11 9 1 0 9 9 7 9 1 9 2
22 10 9 13 0 9 12 9 13 0 9 7 13 15 9 0 9 14 1 9 0 9 2
19 3 3 13 0 9 1 9 9 0 9 13 1 11 2 3 3 1 11 2
24 1 9 11 9 9 11 11 13 2 16 9 1 0 9 4 13 13 9 0 9 1 0 9 2
8 0 9 15 13 9 1 11 2
22 1 0 9 9 13 9 1 9 7 0 9 1 0 9 2 16 15 3 13 0 9 2
34 0 9 13 7 9 9 9 2 7 15 3 13 14 12 3 0 9 1 0 9 9 0 9 7 13 15 13 9 1 0 9 0 9 2
14 13 2 14 3 13 1 9 2 13 15 13 9 0 2
10 13 7 13 1 9 0 9 1 9 2
23 13 13 2 13 2 13 9 2 15 13 3 1 9 9 11 0 9 10 9 1 0 11 2
34 15 4 13 13 2 16 0 13 11 1 10 9 3 1 9 0 2 1 0 9 13 11 12 1 0 0 9 0 9 2 3 11 2 2
7 13 0 13 0 7 0 2
26 0 9 13 3 0 9 2 1 1 15 2 16 0 9 0 9 13 13 0 9 9 0 9 7 11 2
16 13 15 1 10 9 13 7 13 0 2 16 15 13 3 0 2
35 1 0 9 13 15 0 13 12 2 1 15 9 13 9 0 9 0 9 2 9 2 7 9 15 1 15 2 3 0 9 1 12 0 9 2
12 9 0 9 1 9 11 11 13 15 14 9 2
9 9 0 9 13 7 7 0 9 2
16 11 11 13 0 9 2 15 4 3 9 1 0 11 13 13 2
4 11 13 0 9
5 11 2 11 2 2
32 13 0 9 9 0 0 9 0 9 4 13 0 3 3 2 16 4 15 13 2 3 0 9 2 15 4 9 9 13 9 2 2
16 1 11 15 3 13 9 9 0 7 9 0 9 11 11 11 2
11 2 1 9 15 7 3 13 2 2 13 2
12 9 9 11 1 15 3 13 2 7 3 3 2
13 3 0 9 1 9 13 11 1 2 3 0 2 2
27 0 9 11 13 1 15 15 2 16 0 0 9 13 0 9 7 13 15 9 1 9 1 0 9 10 9 2
9 1 9 9 13 9 2 13 11 2
15 0 9 9 11 11 3 1 11 13 1 10 0 9 11 11
5 9 11 11 2 11
4 9 15 13 9
5 11 2 11 2 2
20 1 0 9 9 9 11 2 11 1 11 13 4 11 13 0 9 1 0 9 2
29 13 15 3 0 9 11 2 11 1 9 9 1 0 9 1 9 0 9 9 11 2 15 15 13 1 9 0 9 2
11 2 9 0 13 2 2 13 11 9 11 2
5 0 9 1 11 13
2 11 2
26 9 1 0 9 7 0 0 9 2 15 1 0 9 13 0 9 1 9 12 2 13 9 0 0 9 2
6 13 15 3 9 9 2
20 0 9 1 0 9 13 9 1 0 9 1 9 13 10 9 1 0 0 9 2
6 11 13 1 9 1 9
2 11 2
21 0 11 13 9 13 1 9 0 1 9 9 2 15 1 9 12 13 0 0 9 2
12 1 10 9 15 3 13 9 9 11 1 11 2
28 3 0 9 11 11 2 11 3 13 2 16 0 11 13 1 0 9 1 9 1 11 2 11 2 10 0 9 2
22 1 9 0 9 15 11 3 13 13 9 1 9 0 9 2 15 4 13 7 0 9 2
3 3 1 9
28 1 0 9 16 1 12 9 1 9 13 3 12 0 9 1 9 9 11 1 11 2 15 15 13 3 0 9 2
19 9 13 0 12 9 7 0 0 9 13 9 2 15 13 3 1 12 9 2
24 10 9 13 9 9 15 2 16 11 13 3 0 9 1 9 1 9 0 9 2 3 9 13 2
16 9 0 0 9 1 9 3 1 11 9 13 1 2 0 2 2
26 9 3 9 3 13 1 15 2 16 13 0 9 9 1 0 9 9 2 15 13 1 0 9 0 9 2
5 0 2 0 0 9
2 11 2
17 9 1 0 9 13 3 9 9 11 7 11 11 11 7 11 11 2
36 2 10 0 9 15 13 15 9 2 15 1 9 13 2 7 13 3 0 2 16 13 1 0 9 2 2 13 9 11 1 0 0 9 1 11 2
21 13 2 16 9 12 9 1 1 10 0 9 13 2 3 0 16 1 0 9 2 2
34 0 9 9 11 11 13 1 10 9 9 2 16 1 9 12 9 13 10 9 10 2 16 4 15 0 0 2 0 9 13 7 9 0 2
5 1 9 11 2 11
2 9 9
7 0 9 11 1 11 11 11
17 9 9 11 7 11 2 15 15 13 1 9 3 2 13 0 9 2
13 11 15 13 10 0 9 0 9 1 9 0 9 2
73 3 13 9 1 11 0 9 0 0 0 9 2 11 2 2 11 11 2 1 15 15 1 0 11 7 1 11 13 9 0 9 11 11 2 9 9 0 9 2 11 2 1 9 9 11 11 15 13 0 9 2 9 9 2 11 11 7 11 11 7 1 11 13 7 9 0 9 2 11 2 11 11 2
20 9 11 15 13 1 9 1 9 0 9 1 11 7 13 15 9 1 0 9 2
11 9 11 15 1 9 1 11 13 3 3 2
45 11 2 11 3 1 11 13 2 16 11 4 1 11 13 2 7 0 9 2 7 10 0 9 11 11 2 9 0 9 9 2 13 2 16 1 11 13 2 0 7 0 0 9 2 2
10 1 10 9 15 0 9 1 11 13 2
7 0 9 15 13 1 9 2
11 1 15 11 7 11 15 13 1 9 11 2
41 3 15 13 1 9 9 0 9 1 11 2 3 7 13 2 16 13 2 14 15 1 9 2 13 15 2 16 4 1 0 2 0 2 0 9 2 4 13 9 9 2
44 0 9 13 1 10 9 3 3 7 3 2 3 3 2 7 3 2 15 1 11 13 2 16 15 13 14 14 13 0 9 1 0 9 2 15 14 2 13 2 1 0 0 9 2
11 7 13 9 11 13 9 1 9 1 11 2
18 1 0 0 9 13 3 0 9 1 9 9 9 2 0 11 7 11 2
16 1 15 13 3 13 9 0 9 2 16 2 13 2 11 11 2
20 7 13 11 0 13 15 7 1 9 11 2 13 2 16 13 9 1 9 9 2
38 11 7 10 9 13 13 2 3 7 13 2 13 2 14 15 13 0 9 0 0 9 2 15 3 1 9 1 0 2 0 9 13 9 1 9 0 9 2
12 2 11 15 3 9 13 0 9 1 11 2 2
31 7 3 15 9 11 2 11 3 13 2 3 15 13 1 10 9 2 7 16 13 12 9 1 9 9 2 13 15 1 9 2
6 9 13 2 7 0 2
29 0 9 13 10 9 2 9 15 1 15 13 1 15 7 1 15 2 13 15 1 15 10 9 2 13 15 0 9 2
23 15 13 12 2 11 15 1 11 13 13 1 9 9 2 11 13 13 1 9 0 0 9 2
14 1 0 9 2 16 9 0 0 9 2 4 13 9 2
28 0 9 1 0 0 9 7 1 3 0 9 9 11 4 13 9 7 12 9 13 9 13 2 16 0 9 2 2
10 3 15 0 2 3 7 9 0 9 2
31 3 15 2 15 12 9 13 2 11 13 2 16 14 0 9 2 7 7 15 13 1 14 13 0 2 0 9 1 0 9 2
14 11 13 2 16 13 9 1 9 1 15 0 0 9 2
13 9 13 2 15 1 15 11 7 11 1 9 13 2
44 1 0 9 12 9 1 9 0 9 2 0 12 9 1 9 2 15 13 0 9 0 9 2 13 12 2 9 2 9 9 2 9 0 9 2 15 13 13 12 2 12 5 9 2
28 0 14 13 9 0 9 2 0 9 0 9 7 3 1 0 9 13 0 0 0 9 1 3 12 2 12 5 2
7 9 11 13 0 9 10 9
2 9 11
5 9 1 11 9 9
2 11 2
31 3 12 9 0 0 9 13 7 0 12 4 13 1 0 9 1 9 2 1 10 9 15 13 9 9 1 0 9 1 11 2
16 13 15 3 9 0 9 11 1 11 2 11 2 7 0 9 2
27 3 12 0 9 13 1 9 3 1 9 9 0 9 2 3 15 13 3 16 12 9 3 1 0 9 11 2
14 9 11 13 2 16 13 0 13 2 15 13 9 9 2
5 0 9 11 15 13
2 11 2
26 1 9 3 12 9 15 1 0 0 9 1 0 9 13 0 9 0 0 9 2 11 2 0 11 11 2
10 9 11 7 3 13 0 12 9 9 2
29 1 9 0 0 9 2 15 4 13 1 9 12 1 0 12 9 0 9 2 15 1 11 3 13 3 12 9 9 2
25 1 0 9 13 0 9 9 1 11 1 12 9 9 13 0 9 9 11 2 11 2 1 12 9 2
20 0 0 0 9 13 3 3 9 12 9 2 7 1 10 9 15 13 0 9 2
29 0 0 9 2 15 1 9 9 1 9 13 1 0 9 1 9 2 1 0 0 9 13 1 0 9 14 0 9 2
32 0 9 9 3 0 9 2 10 0 9 1 9 2 11 11 2 1 12 9 13 0 9 1 9 2 13 14 12 9 0 9 2
48 3 13 3 0 9 2 3 3 0 13 11 1 9 0 11 2 3 13 3 12 9 1 12 9 9 0 9 7 1 9 0 2 11 2 3 1 9 3 1 12 9 9 13 11 9 9 11 2
29 0 9 13 2 16 11 15 13 1 9 0 2 11 14 0 9 0 9 9 2 7 3 0 9 7 9 0 9 2
4 9 4 13 3
2 11 2
32 0 7 0 9 3 1 11 13 9 2 16 9 1 0 9 4 3 13 2 3 16 4 15 13 0 13 1 0 9 1 9 2
36 1 11 7 13 9 2 16 13 11 1 14 13 9 1 0 9 3 2 16 15 0 9 13 1 9 11 7 1 9 11 2 13 3 9 11 2
4 9 1 0 9
8 3 13 12 9 1 0 9 2
15 13 9 0 9 2 1 15 1 0 9 13 1 0 9 2
18 12 2 9 0 9 0 0 9 0 9 9 1 0 11 2 11 2 2
18 13 9 2 13 0 9 7 0 9 2 15 9 9 13 2 13 13 2
16 12 2 13 12 1 9 0 9 1 0 0 9 2 11 2 2
4 13 12 9 2
16 12 2 1 9 9 13 0 0 9 1 11 2 0 11 2 2
4 12 9 13 2
13 12 2 9 1 9 0 9 1 11 2 11 2 2
7 0 9 13 0 9 9 2
21 12 2 9 0 9 0 0 9 2 11 2 2 13 15 9 9 1 0 9 2 2
5 13 1 9 9 2
5 9 13 3 9 2
12 12 2 13 0 9 0 0 9 2 11 2 2
9 1 9 9 0 9 13 12 9 2
17 12 2 9 0 9 0 11 11 1 11 2 11 2 9 11 2 2
9 3 13 9 9 2 9 0 9 2
8 0 0 9 13 1 0 9 2
9 12 9 13 2 14 12 9 13 2
8 0 0 9 1 9 0 9 2
22 12 2 1 0 9 0 0 11 2 9 11 12 2 11 2 13 12 9 0 0 9 2
4 12 9 13 2
23 2 9 0 9 1 0 9 1 9 11 2 11 2 13 0 9 9 0 9 1 9 11 2
10 12 9 13 2 0 9 9 1 9 2
15 2 9 12 9 0 9 1 0 9 11 2 0 11 2 2
4 13 12 9 2
17 2 9 0 0 9 1 0 9 1 11 2 11 2 9 11 2 2
6 0 9 13 12 9 2
16 12 2 13 0 0 9 1 0 9 0 0 9 2 11 2 2
6 0 9 13 9 11 2
13 12 2 9 1 0 9 0 0 9 2 11 2 2
17 1 9 0 9 9 1 9 12 9 13 1 9 2 3 13 9 2
3 12 0 2
24 12 2 1 0 9 1 11 2 11 2 9 11 2 15 13 9 9 9 0 1 9 0 9 2
15 12 9 13 2 12 9 13 2 1 0 9 0 9 9 2
21 12 2 9 7 0 9 12 1 12 9 0 9 1 11 2 11 2 3 11 2 2
24 3 3 12 0 7 12 0 2 3 12 9 13 2 13 12 9 0 9 1 0 9 12 9 2
18 1 9 12 13 1 0 9 3 1 12 9 9 2 1 10 12 9 2
20 1 9 12 13 0 9 9 2 16 9 0 9 13 1 9 12 7 12 12 2
10 1 11 13 13 1 12 9 9 9 2
11 1 12 9 7 9 13 1 12 9 9 2
9 1 0 9 4 13 3 12 9 2
10 1 9 12 13 1 9 9 12 9 2
17 12 2 1 0 9 11 2 11 2 13 1 9 12 9 9 9 2
14 13 14 10 0 9 2 7 9 9 13 9 0 9 2
16 12 2 9 1 0 9 0 9 0 11 1 11 2 11 2 2
8 13 1 0 9 9 2 11 2
4 9 13 0 11
12 11 13 11 7 10 0 9 2 3 9 1 11
2 9 9
2 11 11
42 16 9 1 11 0 9 3 13 9 0 9 11 11 7 10 9 9 11 11 1 9 13 2 3 15 11 13 1 0 9 1 0 11 2 13 9 9 11 11 1 11 2
47 11 9 1 0 11 7 1 11 13 0 9 2 13 9 0 9 1 0 0 9 7 1 10 9 13 2 3 3 2 7 1 15 3 2 9 0 9 2 1 15 4 15 1 9 13 13 2
11 10 9 0 9 10 0 2 9 2 13 2
11 1 9 11 11 4 15 13 2 16 0 2
20 2 13 1 3 2 3 0 9 2 2 13 11 1 0 0 9 3 1 9 2
20 11 2 13 11 1 15 3 2 2 13 13 9 2 16 4 13 0 9 2 2
17 1 0 9 0 9 13 15 0 9 2 3 3 1 9 0 9 2
18 14 2 15 1 9 15 13 2 16 0 11 3 3 12 0 9 13 2
24 1 10 9 15 13 7 0 9 9 0 11 2 9 11 11 11 2 7 0 9 9 11 11 2
24 0 2 7 0 11 13 1 9 0 9 0 9 1 9 0 9 2 7 3 0 0 0 9 2
32 11 13 2 3 13 2 1 0 9 1 9 13 1 11 3 0 9 16 2 0 2 9 1 11 0 3 2 3 2 0 9 2
26 16 11 10 9 1 0 0 9 13 1 0 9 2 13 9 2 15 1 10 9 13 0 0 9 11 2
39 2 13 1 0 0 9 2 15 13 13 9 1 0 9 1 0 9 7 13 13 0 9 2 2 3 13 11 1 9 2 15 11 13 0 9 1 0 11 2
33 11 2 15 13 1 11 13 9 0 9 13 3 1 0 11 0 9 0 11 2 13 7 1 9 0 0 9 0 7 13 1 9 2
40 0 11 3 1 9 1 9 13 2 16 13 9 1 0 9 1 0 9 2 11 2 2 16 4 13 0 9 0 9 1 0 9 1 11 2 11 15 7 13 2
25 2 1 0 9 4 13 0 11 13 1 0 9 3 3 3 9 1 12 7 12 9 2 2 13 2
18 1 0 9 9 13 9 11 1 9 9 3 0 2 7 3 14 0 2
14 13 11 10 9 13 2 16 4 9 1 0 9 13 2
11 1 10 9 13 1 0 13 3 11 9 2
51 1 9 2 16 11 7 0 11 13 3 1 0 9 1 11 1 9 9 1 0 11 7 9 4 1 10 9 13 2 3 2 13 11 2 13 9 1 0 9 2 16 4 15 13 3 15 2 9 9 2 2
17 9 2 15 15 1 0 0 0 9 13 3 2 13 13 1 9 2
9 7 3 7 1 10 9 13 9 2
12 1 9 1 11 13 11 1 0 9 13 0 2
4 11 13 0 9
8 0 9 11 1 11 11 11 11
13 3 3 0 9 13 3 13 1 9 0 0 9 2
23 1 9 3 0 9 11 11 11 1 0 2 11 11 11 11 13 9 1 0 9 0 11 2
9 0 9 0 9 13 9 10 9 2
25 11 1 11 11 11 11 11 2 9 9 11 2 13 1 9 10 0 0 9 7 13 3 1 11 2
22 0 9 4 1 9 11 13 1 9 12 9 7 3 15 13 0 9 2 9 1 11 2
14 11 13 0 0 9 2 1 10 9 15 3 13 9 2
7 13 15 3 9 12 9 2
23 0 1 9 2 15 13 1 9 0 9 2 15 1 0 9 1 12 9 13 9 0 9 2
8 3 9 13 9 0 9 9 2
21 9 0 9 4 13 2 0 9 2 2 1 15 15 1 9 0 9 13 15 9 2
3 11 1 9
6 9 1 0 9 9 13
2 9 9
2 11 11
22 2 3 13 13 1 0 9 0 9 2 2 13 1 9 3 0 0 9 11 11 11 2
35 10 0 9 13 9 0 9 12 1 9 0 0 0 9 2 11 2 2 15 15 3 13 16 9 0 9 9 0 9 11 11 2 11 2 2
14 11 15 13 1 0 0 9 12 1 0 9 0 9 2
12 9 0 9 15 3 13 10 9 11 7 11 2
22 11 7 0 9 15 3 13 13 9 0 9 7 9 0 9 2 15 13 12 2 9 2
14 1 15 3 13 11 2 13 11 2 0 1 0 9 2
12 13 15 7 1 9 2 15 13 1 0 9 2
27 7 3 13 13 0 9 2 1 15 13 12 0 9 2 11 11 11 2 11 2 7 11 11 2 11 2 2
11 10 9 15 13 0 9 7 13 0 9 2
16 11 11 13 1 9 12 9 9 2 11 13 7 9 10 9 2
28 15 15 13 2 13 3 1 9 0 9 9 11 11 11 2 2 13 0 0 9 7 15 1 15 13 13 2 2
13 11 11 15 13 1 9 13 14 1 0 0 9 2
17 10 9 13 12 9 1 0 9 2 15 10 9 13 12 2 9 2
6 11 13 12 12 9 2
21 3 3 13 0 9 0 9 9 11 11 11 2 2 12 9 15 13 13 13 2 2
12 11 11 4 13 3 1 9 0 2 9 9 2
21 3 4 7 13 1 12 1 15 2 15 1 0 9 13 13 9 1 9 1 9 2
16 1 15 2 15 13 0 9 2 13 3 0 9 9 0 9 2
15 0 13 9 9 7 13 16 12 1 0 0 9 0 9 2
13 13 15 13 2 16 9 1 11 13 3 1 9 2
26 9 13 9 13 15 1 0 9 3 3 2 16 15 0 9 13 1 9 9 7 2 0 9 2 11 2
9 2 10 9 15 3 13 13 2 2
10 9 1 0 9 4 13 13 0 9 2
13 9 3 13 7 9 1 9 15 13 1 0 9 2
13 9 1 9 7 1 9 1 11 7 3 3 13 2
7 0 9 2 7 0 9 2
8 2 11 12 2 12 2 12 2
36 13 4 1 15 3 13 9 1 0 9 2 1 0 9 14 1 9 2 15 4 13 9 7 3 9 10 9 13 3 7 3 1 9 0 9 2
48 1 9 0 9 2 15 1 15 3 13 2 13 3 9 9 7 13 15 2 16 13 14 14 13 9 2 15 13 0 1 9 0 7 3 0 9 1 9 7 9 7 9 10 3 3 0 9 2
12 0 9 1 9 15 3 13 9 11 7 11 2
9 3 15 2 16 15 3 13 9 2
12 9 15 3 13 2 16 9 9 13 1 9 2
40 3 15 13 0 9 2 15 3 2 3 2 1 9 11 11 2 3 13 2 7 16 3 10 9 3 3 2 3 7 3 2 13 2 15 0 2 15 0 2 2
33 9 7 9 1 15 13 9 3 2 3 7 3 15 13 9 13 2 13 9 9 2 3 4 15 13 13 15 0 3 1 0 9 2
23 13 3 1 0 9 1 9 3 0 7 9 9 2 15 4 13 13 0 0 9 12 9 2
22 3 3 15 13 9 2 3 2 3 7 3 15 1 12 9 13 15 0 2 3 0 2
19 13 0 2 16 15 15 13 3 3 3 7 1 9 2 3 7 1 9 2
11 1 15 13 15 2 16 13 10 3 15 2
6 3 15 9 13 3 2
7 13 0 9 1 10 9 2
63 3 2 16 3 3 13 0 10 0 2 0 9 7 13 10 9 14 1 15 2 16 13 3 13 2 3 13 2 13 15 9 1 9 2 7 10 9 15 13 7 15 2 16 13 0 13 0 7 16 13 13 0 15 2 15 13 2 16 4 15 13 15 2
25 0 9 2 15 3 13 2 3 0 9 2 2 13 3 0 2 7 1 9 15 1 15 14 13 2
11 7 3 4 1 15 13 1 10 0 9 2
41 7 3 9 1 10 9 2 3 4 13 13 2 0 9 2 2 13 1 9 11 2 16 13 1 10 2 0 9 2 7 3 1 10 9 3 0 1 9 7 9 2
4 11 11 2 11
4 1 0 9 13
30 1 9 11 15 3 14 12 9 9 13 9 9 10 9 1 9 15 2 16 0 9 13 0 9 1 9 9 0 9 2
14 9 1 9 1 9 0 9 9 7 9 9 3 13 2
29 1 0 9 0 9 4 3 3 9 0 9 13 2 3 13 2 7 16 4 1 0 9 9 0 9 13 0 9 2
23 1 9 2 16 3 13 1 9 9 7 3 0 2 15 1 0 9 9 9 13 7 9 2
34 13 15 3 1 9 2 16 9 13 0 0 9 16 9 9 1 9 7 0 9 9 13 13 3 12 9 2 16 10 9 4 13 13 2
5 9 13 7 0 2
19 0 9 1 0 9 9 7 9 7 1 0 9 4 3 3 13 0 9 2
19 9 9 1 10 0 9 3 4 1 9 13 9 2 1 0 9 0 9 2
8 3 3 13 0 3 3 13 2
25 1 0 9 13 10 9 0 9 1 9 7 9 9 2 9 9 2 3 3 0 9 1 0 9 2
33 9 2 15 4 13 1 0 9 13 3 0 9 2 7 15 3 7 15 2 15 15 3 13 7 15 15 3 13 2 13 3 0 2
34 0 9 1 0 9 13 3 9 2 16 4 13 1 9 3 15 2 16 3 3 0 0 9 0 9 13 9 2 15 13 0 0 9 2
6 1 9 11 11 2 11
14 9 1 9 1 9 9 2 11 12 2 12 2 12 2
16 13 4 9 11 2 11 2 16 4 13 3 9 1 0 9 2
18 7 3 3 1 0 9 1 11 2 3 1 0 1 11 2 0 9 2
11 3 15 13 13 1 9 9 7 14 9 2
11 3 1 0 3 7 3 1 0 1 9 2
15 13 2 16 15 13 3 6 2 16 13 9 0 7 3 2
23 3 2 16 4 13 0 2 13 3 2 16 9 13 0 2 7 1 9 13 3 3 13 2
14 3 13 1 9 12 9 2 15 15 13 13 1 9 2
21 3 3 14 0 9 1 0 7 13 1 11 2 3 13 3 9 1 9 7 9 2
11 13 2 16 9 13 9 2 13 15 9 2
29 7 16 13 2 9 11 2 9 1 9 2 13 15 9 9 2 3 1 9 2 6 1 9 7 6 1 9 2 2
4 11 11 2 11
5 0 0 9 11 2
5 12 2 0 9 2
4 12 2 0 9
5 0 9 4 13 3
7 11 11 9 0 9 9 9
31 1 11 13 12 2 9 9 2 9 2 9 9 7 9 9 2 2 15 9 13 11 11 2 9 9 9 9 9 9 11 2
30 1 9 13 3 3 13 9 9 9 9 9 0 9 1 9 9 1 9 2 0 9 0 9 9 12 2 9 10 9 2
24 10 9 7 9 0 1 9 2 3 0 2 13 3 0 9 1 9 2 16 3 13 14 3 2
40 0 9 2 1 15 10 9 13 2 13 2 16 0 0 9 1 9 13 0 9 0 9 7 13 15 9 1 0 2 3 0 2 9 2 1 9 7 9 9 2
43 1 10 9 13 0 15 13 2 7 9 1 9 2 9 0 9 7 9 2 16 7 9 9 9 13 2 16 0 9 15 1 0 9 13 1 9 12 2 12 9 9 9 2
12 15 13 3 9 2 9 9 2 7 15 0 2
7 1 9 9 13 10 9 2
39 1 9 12 2 3 4 13 9 9 2 15 13 3 2 15 9 13 1 3 0 9 16 3 2 7 9 0 9 13 3 3 7 9 3 3 0 16 3 2
29 1 9 9 9 0 9 1 0 7 0 9 13 2 16 1 12 9 9 13 3 12 9 0 9 1 9 0 9 2
6 7 3 9 3 13 2
21 1 9 12 13 1 9 0 9 2 7 9 9 0 7 0 9 13 3 9 9 2
30 12 9 0 0 9 3 0 9 13 3 12 9 7 0 9 13 12 9 1 12 9 1 9 2 3 12 5 10 9 2
34 9 9 7 0 9 3 13 2 16 0 9 1 0 9 13 12 2 12 5 10 9 2 7 12 2 12 9 2 9 3 1 0 9 2
10 9 9 7 3 10 9 13 1 15 2
32 13 15 13 15 2 16 1 10 9 15 13 3 0 9 9 2 15 13 1 9 12 9 2 9 1 0 9 0 9 12 9 2
14 13 3 1 0 9 2 15 13 1 0 9 15 0 2
30 13 15 3 1 0 9 2 1 15 13 2 16 0 9 4 1 9 10 9 3 13 1 9 12 2 12 5 0 9 2
26 0 9 9 0 9 15 7 13 1 0 9 2 10 9 1 9 7 9 0 0 9 13 7 13 0 2
8 7 13 0 9 0 9 0 2
31 1 15 13 0 13 1 9 2 16 1 0 9 13 0 9 9 1 0 9 13 2 7 9 0 9 13 0 16 0 9 2
15 0 9 0 9 0 9 7 9 10 9 15 4 3 13 2
28 0 9 15 15 13 2 16 3 4 1 9 13 9 0 9 7 0 9 9 0 1 9 2 13 1 0 9 2
8 9 9 9 13 7 13 9 2
4 9 13 9 9
26 1 0 9 2 15 13 9 1 0 9 1 9 1 9 0 9 9 2 15 0 9 3 13 1 9 2
37 1 9 0 9 13 0 9 9 1 9 1 0 9 2 16 1 0 9 13 9 9 1 11 12 5 7 13 3 3 0 16 1 0 9 9 0 2
29 10 9 9 1 0 9 13 7 1 9 2 16 0 9 13 1 9 2 16 15 1 10 9 3 13 10 0 9 2
29 1 9 9 7 13 0 0 9 2 11 2 2 7 3 9 1 9 3 13 3 13 1 12 9 1 0 12 9 2
25 12 1 0 9 9 9 13 9 9 9 7 9 1 0 9 2 15 13 0 9 1 9 0 9 2
14 9 13 7 9 1 9 0 0 9 11 1 0 9 2
10 15 3 13 3 3 2 16 15 13 2
23 9 9 13 0 9 2 16 4 1 10 9 13 1 0 0 9 7 9 3 9 11 13 2
27 13 3 3 2 7 0 9 13 1 0 9 9 1 9 12 9 1 9 2 15 4 13 3 3 1 9 2
41 0 9 0 9 2 7 16 0 2 4 13 9 9 0 9 1 0 9 2 7 1 0 9 4 13 0 9 9 9 2 16 4 3 13 9 0 9 1 9 0 2
28 0 9 9 11 11 15 13 2 16 11 1 9 9 9 13 15 7 16 13 2 16 15 1 15 0 9 13 2
23 9 7 9 13 9 9 3 13 2 16 1 0 9 9 13 9 9 13 0 9 0 9 2
27 3 1 9 13 9 9 13 9 1 15 2 16 9 9 13 1 11 1 9 7 16 13 9 0 0 9 2
14 15 4 13 9 9 0 1 9 9 2 16 3 9 2
35 1 9 4 13 9 9 7 1 10 9 7 13 15 2 16 15 1 15 4 13 1 0 9 9 9 9 12 1 9 9 9 1 10 9 2
3 2 11 2
6 13 0 9 1 0 9
5 11 2 11 2 2
15 0 9 0 9 2 11 2 3 13 0 9 1 9 9 2
18 1 0 9 4 13 2 16 1 9 9 13 4 13 3 12 12 9 2
12 16 4 10 9 13 2 0 9 4 3 13 2
13 1 0 9 9 13 12 9 2 1 0 12 9 2
14 1 9 0 9 9 1 0 9 9 13 12 0 9 2
44 7 13 9 9 9 14 1 12 2 9 2 3 4 3 13 3 12 12 9 1 0 12 12 9 2 7 3 4 13 0 9 9 12 9 0 9 2 9 12 9 1 9 2 2
31 9 13 2 16 9 2 15 13 9 13 2 13 1 9 1 0 9 9 13 3 12 9 9 1 9 3 12 9 1 9 2
4 11 13 0 9
5 11 2 11 2 2
31 0 9 11 11 13 13 9 0 11 11 13 3 1 0 7 0 9 3 16 12 9 2 3 1 12 3 16 1 0 9 2
17 0 11 13 13 1 0 0 9 9 16 13 11 12 7 11 11 2
17 9 4 1 9 2 0 9 12 9 2 13 13 7 9 1 9 2
29 15 13 1 0 9 3 0 2 0 2 9 13 13 2 2 0 9 7 0 2 15 13 0 9 7 9 13 13 2
19 9 15 3 1 0 9 13 1 0 9 7 13 15 15 3 13 7 13 2
30 11 11 13 9 1 10 9 1 9 10 9 7 14 3 1 0 9 9 2 7 3 9 2 2 7 9 1 0 9 2
5 11 7 11 13 9
5 11 2 11 2 2
15 1 0 9 1 0 9 12 9 13 0 9 12 9 9 2
9 13 1 15 1 9 0 9 9 2
17 9 1 9 9 13 9 2 15 13 9 9 11 12 2 9 12 2
10 9 4 13 9 9 1 12 2 9 2
19 9 10 0 0 9 13 3 0 9 12 9 2 9 2 3 12 9 2 2
13 0 9 11 15 13 1 12 1 12 9 2 9 2
27 9 1 9 9 13 1 12 1 12 9 2 9 2 0 9 1 9 15 13 1 12 1 12 9 2 9 2
16 0 9 11 2 9 0 9 1 3 0 9 2 13 12 5 2
15 9 0 9 1 0 9 15 3 13 1 12 1 12 5 2
18 0 9 11 13 1 0 9 1 0 9 9 2 0 9 7 4 13 2
12 0 9 1 0 9 13 3 0 7 0 9 2
8 11 13 9 1 9 0 9 2
11 1 12 0 9 11 3 13 12 9 9 2
26 3 4 3 1 11 13 2 9 1 9 9 13 9 2 15 13 9 9 11 9 12 2 12 2 12 2
8 9 9 4 13 12 2 9 2
17 1 0 9 9 11 7 11 13 9 11 3 0 9 12 9 9 2
28 0 9 9 0 9 13 1 9 12 12 9 2 9 2 0 9 13 12 9 7 0 9 13 12 9 2 9 2
9 9 0 2 0 9 13 12 5 2
31 1 12 2 12 2 12 13 11 9 1 0 7 0 9 1 9 12 9 2 9 2 15 13 3 3 3 16 9 9 12 2
21 0 9 11 1 0 9 13 1 3 16 0 0 9 7 1 0 9 0 9 9 2
24 0 9 3 13 0 0 9 9 11 1 0 9 3 12 9 2 9 7 1 9 1 12 9 2
17 0 0 9 12 9 4 3 13 1 12 12 9 7 12 12 9 2
5 9 9 1 0 9
2 11 2
26 9 1 9 0 0 9 13 9 9 1 0 9 2 15 13 0 9 9 2 0 0 0 9 2 3 2
22 1 0 9 15 7 4 9 10 9 1 0 9 1 0 9 13 1 9 9 1 9 2
8 13 15 1 0 9 9 11 2
25 0 9 9 1 9 13 1 12 9 2 16 1 9 13 1 12 9 1 12 9 1 9 0 9 2
13 9 10 9 13 9 10 9 1 12 7 12 9 2
19 0 9 9 9 13 0 0 9 9 2 1 15 13 9 3 9 16 3 2
25 1 11 11 2 0 9 11 2 13 1 9 3 3 9 2 15 4 1 0 9 13 1 0 9 2
17 1 9 13 1 11 3 9 9 7 10 0 9 3 4 13 13 2
4 9 1 9 9
2 11 2
11 3 0 9 13 0 9 13 9 9 9 2
19 3 9 13 2 16 4 13 0 0 9 9 13 2 0 9 2 7 9 2
16 0 9 13 3 13 9 9 2 13 9 0 0 9 0 9 2
11 0 9 13 7 0 9 7 0 0 9 2
24 9 12 0 9 3 13 12 9 2 16 0 9 12 7 12 9 1 9 4 9 13 1 0 2
16 9 3 13 3 12 0 9 7 1 15 0 9 12 9 9 2
11 3 1 9 12 4 13 14 1 12 9 2
11 9 0 0 9 7 13 9 0 0 9 2
9 12 0 9 13 0 9 0 9 2
18 0 9 13 0 9 0 11 1 0 11 1 12 2 7 12 2 9 2
12 13 15 3 9 0 0 9 1 9 7 9 2
19 9 13 9 12 2 9 2 3 15 1 11 1 9 0 9 13 0 9 2
4 0 0 2 11
21 0 9 1 9 0 9 1 9 12 9 9 13 1 9 1 11 9 0 2 11 2
31 9 0 9 0 2 11 11 2 11 2 13 0 2 11 2 11 7 11 1 0 0 9 2 13 7 13 9 1 0 9 2
15 10 9 13 13 1 0 9 2 3 9 1 12 9 9 2
28 12 9 9 1 9 9 11 4 13 1 11 7 12 9 9 2 15 15 13 1 9 2 13 3 1 0 9 2
16 11 4 13 1 9 12 16 0 0 9 1 0 9 1 11 2
3 2 11 2
4 9 13 14 11
5 11 2 11 2 2
20 9 1 9 12 12 9 1 12 9 13 1 9 0 9 0 9 0 9 11 2
7 0 9 15 9 9 13 2
26 0 0 9 0 9 11 2 0 2 9 2 2 2 11 2 13 12 9 9 2 0 9 12 9 9 2
10 0 9 0 0 9 13 12 9 9 2
17 0 9 12 9 9 13 1 9 9 7 12 9 9 1 9 9 2
15 1 9 9 13 9 12 9 7 1 0 9 12 9 9 2
13 3 15 9 11 13 1 9 12 1 12 9 9 2
8 0 9 9 13 12 9 9 2
14 0 9 9 13 12 9 2 1 15 12 1 0 9 2
12 9 1 9 1 0 9 13 0 12 9 9 2
20 1 9 13 11 3 12 9 9 2 15 13 1 12 5 3 16 1 9 12 2
38 1 0 9 11 1 0 9 13 9 9 9 12 1 9 1 11 7 11 2 9 11 2 9 0 11 1 11 2 0 9 11 11 7 0 9 11 11 2
26 0 0 9 2 16 13 9 9 1 0 9 11 7 9 0 9 11 2 11 2 13 11 1 10 9 2
4 9 13 9 9
20 3 0 9 9 1 0 9 13 1 0 9 9 2 1 15 15 13 15 13 2
9 9 15 13 7 1 9 0 9 2
24 1 2 0 2 9 13 1 10 9 7 0 9 7 1 10 0 9 13 10 9 7 0 9 2
15 10 9 7 9 15 1 15 3 1 9 0 9 13 13 2
22 9 0 1 9 9 1 9 9 3 13 2 7 15 1 9 1 9 7 1 0 9 2
24 1 11 15 3 9 1 9 12 13 1 9 12 5 2 7 3 1 9 12 15 13 12 5 2
19 9 13 1 12 9 0 9 9 7 1 9 0 0 15 9 9 0 9 2
17 9 9 1 0 9 1 9 13 7 1 0 9 3 3 3 0 2
22 13 15 0 9 9 1 9 1 0 9 2 9 12 9 1 9 7 12 9 1 9 2
14 1 11 13 3 13 0 9 1 12 9 1 12 9 2
23 1 0 0 9 13 3 0 9 1 0 9 2 1 15 3 3 9 13 1 9 3 3 2
13 15 15 3 13 13 9 7 3 13 1 0 9 2
18 1 9 0 9 13 0 9 9 9 3 0 9 2 10 9 3 13 2
18 9 4 13 13 0 9 0 0 9 2 15 13 7 9 3 0 9 2
19 3 15 3 13 0 9 2 13 9 9 0 9 2 15 13 13 9 9 2
18 10 9 4 7 3 3 13 0 9 7 1 0 9 15 13 3 0 2
3 2 11 2
4 11 13 1 9
5 11 2 11 2 2
23 1 0 9 13 1 0 2 0 9 2 0 2 9 2 11 14 9 9 2 9 7 9 2
33 9 1 0 9 10 9 11 11 13 2 16 1 0 0 0 2 0 9 13 9 9 0 9 2 0 9 2 0 9 7 0 9 2
23 0 9 0 9 15 1 9 0 0 9 13 2 13 2 2 13 0 9 0 1 0 9 2
20 0 9 0 9 9 0 0 2 9 2 11 15 13 1 9 2 0 9 2 2
14 3 13 1 9 11 1 9 9 0 9 11 1 11 2
20 0 0 9 11 13 12 2 9 9 1 11 2 11 2 15 13 14 12 9 2
47 16 15 1 10 9 13 1 0 9 9 1 9 2 0 0 9 13 14 12 9 9 2 2 13 1 9 14 12 9 2 15 13 0 9 9 2 14 12 9 4 13 9 1 0 9 11 2
15 1 0 9 12 9 11 10 9 1 9 9 13 1 12 2
26 0 9 11 13 1 9 9 3 12 9 2 9 2 7 0 9 4 9 13 1 0 9 0 2 9 2
2 11 2
18 13 4 3 9 1 9 9 0 9 1 0 11 1 9 12 2 12 2
26 9 4 13 0 9 9 2 0 9 12 9 2 9 2 0 9 0 2 9 2 12 9 2 9 2 2
18 11 13 3 9 0 9 2 0 9 13 11 2 12 9 2 9 2 2
13 1 0 0 9 13 9 1 11 12 9 2 9 2
12 3 13 0 1 9 13 9 12 9 2 9 2
50 10 9 15 3 13 9 0 9 2 12 9 3 2 2 9 15 13 13 1 9 1 0 9 2 3 1 12 9 13 9 2 7 13 13 7 9 9 1 0 9 9 2 1 10 13 9 3 1 11 2
8 0 9 13 9 9 1 11 2
8 0 9 11 13 9 1 12 9
2 11 2
20 0 9 0 9 11 1 0 9 13 12 9 9 1 0 9 14 12 9 9 2
9 13 1 15 0 9 9 9 11 2
22 9 9 13 1 12 9 1 3 12 9 9 7 0 0 9 9 13 3 12 9 9 2
21 9 9 13 1 12 9 9 2 1 15 1 11 11 13 9 1 0 12 9 9 2
22 9 1 9 13 1 9 0 9 3 12 9 9 2 1 15 1 9 9 14 12 9 2
11 9 9 13 1 10 9 3 12 9 9 2
13 1 0 9 0 9 13 1 0 9 0 9 11 2
8 0 9 9 13 12 9 9 2
10 0 9 9 4 13 1 12 9 9 2
19 1 0 9 0 9 13 13 12 9 9 2 15 13 12 9 15 9 9 2
51 0 9 4 13 4 13 1 11 2 11 3 2 12 9 4 13 13 11 9 2 9 2 0 2 2 12 9 11 11 2 12 9 0 9 2 12 9 4 13 13 1 0 9 7 9 4 13 11 7 11 2
20 9 0 9 0 9 11 13 3 12 9 2 15 13 12 9 1 0 9 9 2
11 9 9 1 9 9 12 13 12 9 9 2
15 1 0 9 7 9 0 9 13 1 3 16 12 9 9 2
32 1 9 13 9 1 0 9 7 1 0 9 12 9 2 1 15 13 12 9 1 0 9 2 12 9 1 9 7 12 9 9 2
14 0 9 9 13 3 12 9 7 9 1 9 12 9 2
12 0 0 9 9 13 3 9 0 12 9 9 2
26 11 0 2 9 2 15 13 1 9 0 9 2 0 9 2 0 9 2 9 7 0 9 1 0 9 2
15 3 13 0 9 9 9 2 11 2 11 2 9 7 9 2
9 3 9 13 9 9 7 0 9 2
21 9 9 9 1 9 12 15 13 1 12 2 1 12 2 9 3 1 11 7 11 2
12 0 9 9 1 12 9 3 13 11 7 11 2
16 13 1 15 9 0 0 9 2 11 2 1 10 9 1 11 2
4 11 13 0 9
2 11 2
30 1 0 0 9 0 9 11 11 1 9 12 13 9 9 1 9 1 9 12 9 9 2 9 9 7 9 0 0 9 2
13 9 9 9 0 9 4 13 3 13 12 9 9 2
29 3 13 0 9 0 9 11 11 11 2 13 1 0 9 13 0 9 1 12 12 9 2 7 13 15 13 9 9 2
9 1 0 9 9 13 3 0 9 2
12 3 0 9 13 9 9 2 9 7 0 9 2
20 1 15 9 9 13 1 0 12 9 9 12 9 9 7 9 9 12 9 9 2
11 13 15 2 16 13 1 9 2 0 9 2
13 0 9 15 13 9 1 12 9 7 13 1 9 2
16 1 9 13 0 9 3 9 7 13 0 9 1 9 0 9 2
7 13 15 10 0 9 9 2
28 1 9 12 9 1 0 0 0 11 13 9 14 9 0 9 7 9 0 1 0 9 9 13 10 3 9 9 2
7 2 13 0 2 2 13 2
7 2 13 15 1 15 2 2
7 0 9 1 11 0 9 2
2 9 2
2 9 2
3 0 9 2
11 15 13 9 0 9 2 15 13 0 9 2
20 16 13 10 0 9 2 9 13 9 9 1 9 1 9 7 9 1 0 9 2
31 14 1 9 12 13 1 0 11 2 9 2 9 1 0 9 1 12 5 7 13 4 1 12 5 3 9 7 9 10 9 2
15 1 0 9 1 11 13 3 1 0 9 7 12 9 0 2
23 13 0 2 16 9 1 9 0 9 13 14 3 0 2 3 16 15 13 1 11 0 9 2
26 1 10 9 2 7 2 3 1 12 9 2 4 0 9 10 9 13 2 7 3 10 9 3 3 13 2
22 3 13 3 3 16 9 2 15 13 1 0 9 3 0 9 7 13 3 3 1 9 2
11 0 9 13 3 3 0 7 0 16 3 2
14 1 0 9 0 9 13 3 12 2 12 9 0 9 2
12 3 13 1 9 9 0 14 12 9 0 9 2
24 9 13 3 3 0 2 16 15 2 15 15 13 2 15 3 13 1 2 9 2 9 7 9 2
8 1 9 15 13 14 0 9 2
9 9 0 9 9 13 3 0 9 2
20 7 3 15 2 16 0 9 13 1 10 9 3 0 2 13 10 0 15 9 2
22 2 0 1 9 2 1 9 13 1 3 9 2 15 3 9 9 13 4 9 9 13 2
21 9 0 9 13 0 2 2 13 9 2 11 11 2 11 1 0 0 9 1 11 2
35 2 9 3 13 9 13 3 0 9 1 0 9 2 13 15 15 2 7 3 13 0 9 2 15 4 15 3 13 13 13 1 9 7 9 2
11 7 15 1 0 2 3 0 2 13 2 2
35 0 9 9 0 1 9 13 3 0 1 15 2 16 4 15 13 9 7 9 9 0 9 2 16 0 9 2 0 2 9 15 3 3 13 2
33 0 9 1 0 11 15 3 3 13 1 10 0 0 9 2 2 13 4 15 3 0 9 0 9 7 9 7 13 4 13 0 2 2
22 1 12 9 3 15 10 9 13 3 9 9 2 13 0 9 0 9 7 9 2 2 2
23 0 9 13 10 9 2 16 0 0 9 15 3 13 1 9 9 7 13 15 3 0 9 2
3 7 9 2
15 3 1 9 4 10 9 13 1 0 9 2 13 15 9 2
36 2 16 13 15 2 15 13 0 9 11 11 2 13 11 11 7 13 9 11 11 2 13 0 2 16 3 13 9 2 2 13 9 0 0 9 2
31 15 15 13 9 13 15 15 1 11 2 0 0 9 2 15 13 13 10 2 9 2 14 3 3 2 16 4 13 9 9 2
19 11 3 13 1 12 9 1 11 11 2 15 13 1 9 0 9 0 9 2
10 0 0 9 3 3 13 1 10 9 2
11 11 13 2 16 9 15 0 9 3 13 2
21 2 13 4 13 0 9 2 13 3 7 9 2 15 13 2 16 4 13 1 9 2
15 13 0 2 3 15 10 9 13 0 9 3 16 9 2 2
6 1 0 9 13 11 11
4 9 1 9 9
2 9 9
6 1 10 0 9 13 2
30 13 0 0 9 7 15 2 15 4 13 1 10 9 2 13 2 16 1 0 9 11 1 11 13 3 1 15 3 9 2
4 13 4 13 2
16 11 11 13 1 9 16 9 7 1 15 15 13 12 0 9 2
9 3 3 15 13 12 7 12 9 2
3 13 9 2
17 9 7 9 2 15 13 1 15 2 15 3 13 2 13 7 13 2
14 9 13 9 13 7 9 15 15 3 7 3 13 13 2
10 3 2 10 9 9 13 3 0 9 2
7 9 2 0 13 0 9 2
2 11 11
10 11 11 13 0 0 9 2 12 9 2
14 13 9 7 3 15 0 9 13 1 9 1 10 9 2
10 1 10 9 13 9 0 7 0 9 2
31 12 1 9 2 11 2 0 2 11 11 2 3 11 2 13 1 12 9 0 0 9 1 9 2 1 9 12 13 0 9 2
9 9 11 11 13 1 0 1 9 2
11 9 11 13 2 16 9 1 15 11 13 2
9 16 13 9 9 2 11 14 9 2
5 15 1 15 13 2
8 1 0 9 13 9 7 9 2
19 15 13 15 0 2 3 15 0 2 7 9 13 2 16 0 9 13 11 2
9 9 9 13 2 16 15 3 13 2
6 16 13 15 0 9 2
12 9 2 15 13 7 3 2 16 15 13 9 2
8 3 4 1 15 13 0 9 2
5 13 0 7 9 2
9 13 4 11 2 3 13 1 9 2
10 0 4 13 2 16 4 4 13 9 2
13 16 9 9 9 2 9 2 2 2 1 15 3 2
10 9 4 14 1 10 9 13 13 0 2
12 13 15 2 16 11 12 9 1 9 3 13 2
8 7 9 13 1 15 3 15 2
10 11 11 13 3 9 2 9 7 9 2
8 2 13 2 16 9 13 2 2
4 2 13 9 2
8 13 4 13 1 9 7 13 2
8 15 13 3 0 9 1 9 2
18 7 9 4 15 13 13 3 1 9 7 14 1 0 9 1 9 2 2
13 2 10 9 4 13 2 16 4 13 1 9 2 2
4 2 3 0 2
10 3 4 15 13 2 16 15 13 9 2
18 3 4 13 12 2 9 12 1 9 13 9 1 11 7 13 4 15 2
10 1 10 9 15 3 7 3 13 9 2
5 1 9 15 13 2
6 16 13 2 9 2 2
11 16 16 15 3 13 9 2 15 3 13 2
5 7 1 10 9 2
24 3 13 12 9 9 9 2 13 0 2 16 15 9 13 13 2 16 4 13 0 9 1 9 2
10 7 14 2 16 13 9 14 0 2 2
9 2 0 9 13 1 15 3 2 2
6 2 1 10 9 14 2
13 15 15 3 3 13 2 10 4 0 13 9 9 2
16 9 1 10 9 7 9 13 2 2 2 13 2 15 13 9 2
9 9 13 0 2 0 9 1 9 2
13 3 9 13 2 16 4 3 13 2 16 9 13 2
3 3 13 2
18 10 9 1 15 13 3 3 0 2 16 3 15 3 13 2 16 13 2
8 7 13 1 15 2 16 13 2
4 13 3 9 2
7 14 13 0 13 0 9 2
23 15 2 16 15 15 0 13 7 13 2 3 4 13 9 1 9 2 15 1 15 3 13 2
5 13 0 13 9 2
18 3 15 3 13 2 16 13 1 0 9 2 3 13 9 2 13 9 2
6 7 9 15 1 15 2
7 13 15 9 7 15 9 2
17 16 4 0 13 2 1 10 13 9 2 2 2 3 15 3 14 2
5 13 4 13 0 2
7 16 4 13 13 3 9 2
6 15 4 13 1 9 2
10 0 9 11 13 0 9 1 0 9 2
12 13 2 16 4 15 1 0 9 13 0 9 2
5 16 13 1 9 2
12 13 15 2 16 7 15 13 15 13 9 9 2
8 7 13 2 16 1 0 2 2
8 2 3 4 15 13 9 2 2
19 2 1 9 12 4 13 1 9 3 1 9 11 11 2 0 9 0 9 2
7 15 0 13 9 1 11 2
22 13 1 15 3 3 2 16 15 0 9 1 0 9 4 3 13 2 16 4 15 13 2
7 3 4 15 13 0 9 2
15 9 15 12 13 1 9 2 13 10 9 7 9 15 13 2
17 13 15 3 2 3 4 13 7 13 15 1 12 12 10 9 2 2
12 2 13 15 2 16 9 13 0 2 2 2 2
8 2 11 15 13 13 15 9 2
11 3 4 15 13 2 3 13 0 1 9 2
5 13 15 0 9 2
18 16 13 0 2 1 15 9 13 15 2 15 13 0 13 1 0 9 2
4 9 13 0 2
4 0 7 0 2
5 13 1 0 9 2
11 13 15 1 15 3 7 13 15 15 13 2
11 13 0 13 3 2 3 4 15 15 13 2
6 13 1 15 13 9 2
11 13 15 9 2 9 2 0 16 15 2 2
16 2 16 4 13 1 9 2 3 4 13 0 7 14 0 9 2
8 2 2 13 15 0 2 0 2
13 3 2 16 13 15 0 1 9 2 1 15 13 2
7 1 9 4 13 10 9 2
10 10 9 15 3 13 1 9 16 13 2
5 16 4 13 0 2
4 15 15 13 2
4 13 4 15 2
7 1 9 3 13 0 9 2
14 9 2 9 9 2 15 4 13 0 2 9 2 2 2
6 13 4 15 1 9 2
10 7 3 13 9 2 16 13 15 9 2
4 14 0 9 2
7 13 4 1 15 15 2 2
8 2 1 9 15 15 13 2 2
4 2 3 13 2
17 16 4 15 13 1 0 2 13 9 0 2 15 15 13 1 9 2
7 13 4 15 7 1 9 2
16 12 10 0 9 2 9 2 15 13 3 1 9 13 0 9 2
5 13 1 15 9 2
10 3 15 15 13 1 10 9 1 9 2
10 13 3 10 10 9 9 1 11 3 2
4 7 1 9 2
8 14 3 15 15 13 1 11 2
11 3 4 13 1 0 9 15 0 7 0 2
5 0 9 12 9 2
5 7 13 7 9 2
28 3 2 16 13 9 7 13 1 11 9 1 9 2 13 1 15 13 9 2 3 15 13 13 9 2 2 2 2
7 2 7 13 15 9 2 2
5 2 15 3 14 2
15 7 1 15 2 3 15 13 10 9 2 13 9 1 9 2
25 13 0 3 1 15 2 16 4 15 12 1 9 13 1 9 2 13 0 9 7 13 1 9 2 2
10 2 3 4 13 13 9 7 9 2 2
10 2 9 15 0 13 9 2 15 13 2
16 3 3 2 16 1 12 4 15 13 13 1 12 9 0 9 2
5 3 15 13 0 2
15 13 9 2 15 2 16 3 15 1 15 13 2 0 13 2
18 3 15 13 1 9 2 2 2 7 13 3 15 2 15 13 0 2 2
8 9 2 11 2 11 2 11 2
4 0 9 13 9
9 0 9 15 13 13 9 7 0 9
2 9 9
7 9 1 9 13 13 9 2
23 0 9 2 15 15 3 13 14 1 10 9 1 9 2 4 13 3 1 9 9 3 13 2
9 9 13 13 2 3 15 9 13 2
16 13 13 9 13 10 9 3 1 9 3 9 2 15 13 3 2
9 9 0 9 3 15 1 15 13 2
15 9 7 9 15 3 13 1 0 9 2 1 0 0 9 2
2 11 11
26 2 15 15 15 13 10 9 13 2 2 13 15 11 11 2 15 13 1 0 9 11 1 0 9 11 2
10 13 9 2 16 9 15 13 10 9 2
40 3 13 1 9 9 2 3 15 13 9 1 9 7 9 2 15 3 13 10 9 2 16 4 10 9 13 10 9 2 16 13 0 9 7 13 1 15 15 13 2
19 3 7 9 9 13 13 9 13 10 9 2 1 9 1 9 13 10 9 2
34 11 13 3 3 3 0 1 10 9 2 15 4 3 13 3 0 9 2 7 9 2 15 13 10 9 1 0 9 2 3 13 7 3 2
3 0 0 9
23 2 1 9 13 1 10 9 12 9 2 7 10 9 3 15 1 9 1 10 9 3 13 2
10 1 9 13 1 9 11 14 12 9 2
7 0 12 13 1 0 9 2
19 0 9 15 4 13 13 7 15 2 15 1 15 4 13 2 13 13 3 2
13 0 9 13 13 0 9 2 2 13 15 11 11 2
6 9 13 0 0 9 2
24 1 9 12 9 1 9 0 9 15 13 9 1 9 12 3 2 1 0 9 13 9 1 9 2
16 1 9 9 1 9 9 13 0 9 0 1 9 1 0 9 2
29 1 0 0 7 0 9 15 13 13 7 1 0 2 3 9 9 2 9 9 7 3 9 2 15 13 3 0 9 2
12 0 9 15 3 13 9 1 0 0 0 9 2
20 0 9 2 15 13 9 2 1 15 4 13 1 9 2 13 9 9 7 9 2
27 9 15 13 2 3 13 9 1 9 2 15 13 1 10 9 2 13 15 13 9 7 0 9 3 1 9 2
31 9 4 3 13 9 13 3 1 15 2 3 15 1 9 13 2 10 4 1 15 13 9 2 15 15 1 10 9 13 3 2
23 9 7 10 9 13 1 9 1 9 0 2 7 1 10 9 15 13 2 16 13 0 9 2
5 9 1 9 1 9
11 12 9 1 0 9 4 13 3 0 9 2
17 1 9 13 9 1 10 9 2 15 13 3 7 13 15 1 9 2
14 2 13 15 1 15 15 13 2 3 7 1 0 9 2
6 10 9 13 1 9 2
15 9 15 3 1 9 13 1 0 9 2 15 13 10 9 2
9 12 9 4 13 9 0 1 0 2
17 9 10 9 7 1 15 13 2 13 3 13 2 2 13 11 11 2
6 0 0 9 13 3 2
7 9 7 9 15 9 13 2
16 9 9 4 1 12 9 13 1 0 9 2 0 9 13 9 2
17 9 9 1 9 13 0 9 1 0 9 2 1 0 14 1 0 2
14 3 13 1 15 3 0 9 2 3 1 9 13 0 2
23 13 15 3 1 9 0 9 2 9 0 9 2 9 9 0 9 2 9 2 9 1 9 2
10 1 9 1 9 13 7 9 1 9 2
14 13 7 9 1 15 2 15 15 13 13 1 9 9 2
22 13 0 2 16 4 13 0 13 9 1 0 9 2 3 1 9 2 15 15 9 13 2
4 1 9 9 2
32 1 9 7 9 0 9 15 3 3 13 7 0 0 9 2 15 13 1 15 9 7 15 15 3 13 13 1 9 9 1 9 2
24 1 0 9 13 4 3 12 1 12 0 9 1 9 9 13 2 1 0 4 13 10 0 9 2
27 9 2 15 13 9 1 0 9 2 13 2 16 13 9 2 3 13 9 2 15 15 13 7 1 0 9 2
8 1 10 9 13 13 7 9 2
19 7 9 0 1 9 9 11 3 13 9 1 0 0 9 1 0 9 9 2
23 15 14 16 4 15 15 13 10 9 1 9 0 9 7 13 1 15 14 1 0 0 9 2
5 0 9 1 0 9
16 0 11 13 10 0 9 3 2 16 1 15 13 7 0 9 2
18 1 9 1 15 13 2 7 1 9 1 9 1 9 15 0 9 13 2
12 0 11 3 3 13 1 9 16 1 0 9 2
18 13 15 9 7 9 2 16 15 12 9 13 1 9 0 1 0 9 2
9 11 13 1 9 3 1 0 9 2
10 15 1 9 9 13 10 9 1 9 2
12 11 15 13 2 13 14 0 9 7 13 9 2
5 9 9 13 9 2
16 13 1 0 9 2 0 9 13 9 7 13 1 0 15 11 2
10 1 0 12 9 11 13 1 0 9 2
18 11 4 13 1 12 7 12 9 7 13 15 9 1 0 9 1 11 2
2 11 11
24 15 15 1 0 9 13 14 1 9 2 3 11 9 13 2 16 9 1 9 13 3 1 9 2
22 3 0 0 9 1 0 9 2 16 4 15 1 15 13 0 9 3 0 1 0 9 2
16 11 13 3 3 1 0 0 9 1 9 0 1 9 0 9 2
15 0 9 10 9 9 3 13 13 1 9 1 3 0 9 2
23 7 9 13 3 10 9 7 13 13 13 1 10 0 9 2 3 15 13 1 9 10 9 2
58 1 15 4 13 15 0 2 16 4 13 9 1 0 9 2 15 15 3 13 1 9 2 13 12 9 1 9 1 0 9 2 7 1 15 15 9 3 13 2 16 0 9 13 13 1 15 3 2 0 2 2 15 1 0 9 13 15 2
42 1 9 1 0 9 9 0 9 15 9 1 0 9 9 13 1 10 9 2 16 10 0 9 1 0 9 1 11 1 11 13 1 9 1 0 9 1 0 11 0 9 2
38 9 13 9 9 1 9 2 1 0 9 2 1 0 9 2 1 9 1 9 1 0 0 9 11 7 11 2 15 15 9 1 0 9 14 3 13 13 2
10 3 15 13 0 9 1 9 0 9 2
4 10 0 9 2
11 15 0 13 9 2 15 0 15 13 13 2
16 9 1 12 9 3 13 9 2 1 9 2 1 0 0 9 2
62 2 0 9 3 15 13 9 13 2 13 2 9 2 2 13 4 3 9 1 9 1 0 9 7 10 9 1 9 1 0 9 2 2 16 4 15 15 13 2 13 4 3 9 1 9 2 16 4 15 13 2 13 4 12 9 2 7 15 4 3 13 2
24 2 9 13 2 16 16 4 11 13 11 2 7 12 1 15 4 13 9 1 9 1 0 9 2
29 0 9 11 15 3 13 13 1 0 9 9 1 9 1 9 9 2 15 4 9 0 9 13 1 0 0 9 0 2
24 2 14 15 9 2 16 3 15 13 13 2 13 9 1 0 9 2 15 4 3 1 9 13 2
11 3 15 13 2 3 3 15 1 9 13 2
5 1 0 9 13 9
13 1 0 11 0 9 13 12 2 9 0 0 9 2
16 12 1 9 9 1 9 0 9 13 3 9 0 9 11 11 2
2 11 11
22 16 13 9 0 0 9 9 0 2 3 13 2 16 0 9 15 3 13 7 9 0 2
20 3 0 9 1 11 2 1 9 12 2 13 0 9 1 9 12 9 1 9 2
18 1 0 12 9 4 13 0 0 9 7 9 2 9 2 9 2 2 2
32 1 9 12 13 0 9 0 0 9 1 0 0 0 9 2 3 4 0 9 13 12 9 1 9 0 9 0 9 2 9 11 2
5 3 10 9 13 2
25 2 1 0 9 2 3 13 7 10 9 0 9 2 13 9 3 9 0 9 2 2 13 11 11 2
30 2 7 15 3 1 9 2 13 3 9 1 10 9 16 11 11 2 11 2 11 11 7 11 11 2 2 3 1 9 2
20 9 13 0 9 0 9 11 2 15 16 10 0 9 1 9 13 0 11 11 2
15 13 15 9 9 3 3 3 2 1 10 9 7 3 3 2
16 2 15 1 9 2 15 3 1 11 13 2 13 1 10 9 2
25 2 3 4 13 13 0 9 0 9 2 0 0 9 1 9 9 11 7 1 0 9 1 9 11 2
12 3 13 3 9 9 11 1 0 9 11 11 2
14 15 13 0 0 9 1 0 9 2 2 13 9 11 2
12 2 1 9 10 9 1 0 3 13 13 9 2
25 3 9 1 9 2 15 1 11 13 0 7 0 9 2 15 13 0 9 7 0 0 15 9 13 2
22 16 13 1 9 2 0 11 2 9 9 9 15 13 1 0 9 2 7 13 0 9 2
26 0 9 10 10 9 15 15 7 13 0 2 3 9 1 11 11 7 9 2 16 15 3 13 11 11 2
9 1 0 9 15 3 13 3 13 2
9 1 0 0 9 13 9 0 9 2
28 9 13 1 15 2 16 0 9 9 13 1 9 10 10 9 7 1 0 9 7 9 13 0 2 2 13 11 2
10 15 2 3 2 3 12 2 12 2 2
26 0 9 11 13 3 3 2 12 2 9 0 9 11 11 11 1 9 11 11 7 1 0 9 11 11 2
24 3 4 1 9 12 2 9 0 7 0 9 9 13 9 13 15 9 0 1 9 1 9 9 2
21 1 0 13 3 2 11 11 2 11 11 11 11 2 11 11 2 9 9 7 0 2
7 9 13 1 12 2 9 2
12 9 9 12 4 13 1 9 9 11 1 11 2
6 13 1 12 2 9 2
20 0 9 1 9 9 1 9 13 13 1 0 0 9 1 11 1 12 2 9 2
12 9 7 9 13 1 0 9 0 9 11 11 2
7 9 13 1 12 2 9 2
19 0 9 0 9 11 11 2 12 2 4 3 13 1 0 9 1 0 11 2
22 11 15 13 3 0 9 2 1 15 13 12 1 0 2 9 11 2 12 2 12 2 2
5 2 11 2 9 11
7 1 0 9 4 13 0 9
31 1 0 0 9 4 1 9 3 13 12 0 9 1 0 0 9 0 2 0 7 0 9 2 0 7 0 1 9 0 9 2
8 10 9 13 9 9 3 3 2
9 9 15 3 13 0 9 10 9 2
2 11 11
31 0 9 15 1 9 1 15 13 3 0 9 0 1 9 0 2 0 9 7 9 7 1 9 9 11 11 15 9 9 13 2
22 1 9 1 9 9 9 2 15 4 13 3 0 9 9 2 13 0 9 0 0 9 2
9 15 3 13 1 0 9 9 11 2
7 9 0 9 13 7 0 2
20 13 2 16 9 2 9 9 7 13 3 9 9 2 0 1 0 9 10 9 2
9 1 9 12 0 9 13 9 0 2
24 1 10 9 13 9 9 0 9 1 0 9 2 1 15 13 12 7 12 9 1 0 1 9 2
19 1 12 0 9 0 1 0 9 9 9 13 0 9 2 12 9 2 12 2
10 1 15 4 1 9 13 3 12 9 2
31 0 13 2 16 0 9 15 13 3 1 0 9 2 7 13 15 0 9 1 9 0 0 9 2 15 13 1 0 9 9 2
17 13 3 1 9 2 16 0 0 7 0 9 13 0 9 0 9 2
43 2 15 15 13 2 16 0 9 13 15 2 16 15 3 4 13 1 0 0 9 2 16 13 1 3 1 0 9 11 2 16 13 11 2 7 11 2 16 13 1 11 11 2
28 3 15 9 3 13 7 13 15 15 2 15 15 15 13 1 9 1 9 2 2 13 11 11 1 9 0 9 2
47 1 0 9 1 9 0 9 15 13 0 2 0 9 1 0 9 2 7 15 1 9 10 3 0 9 7 9 2 11 0 11 2 9 11 11 2 9 11 11 2 9 11 11 0 2 2 2
17 16 4 9 9 13 2 16 9 13 0 9 3 1 0 0 9 2
10 0 9 13 7 0 9 7 0 9 2
12 1 9 11 11 15 13 11 11 7 11 11 2
25 9 11 7 10 0 9 9 2 15 13 9 1 9 2 7 13 2 16 0 9 13 3 1 9 2
9 9 2 11 11 13 1 0 0 9
5 9 11 11 2 11
4 9 13 1 9
27 9 2 12 1 9 0 9 0 9 13 13 9 13 15 1 0 9 1 9 15 2 15 13 3 1 9 2
26 0 9 11 11 7 11 11 1 0 11 2 1 9 1 9 11 11 1 0 9 2 10 9 3 13 2
19 9 13 3 2 1 0 9 7 9 9 3 13 9 0 0 9 1 9 2
18 9 11 11 13 3 0 10 3 0 9 1 15 9 7 0 0 9 2
15 9 13 9 0 7 0 2 14 15 9 15 7 13 3 2
26 0 0 0 7 0 9 13 1 0 9 7 10 9 13 14 9 9 2 7 3 7 0 9 0 9 2
29 3 15 13 9 2 1 9 9 2 2 7 0 7 0 9 0 9 2 15 1 15 3 13 13 10 0 0 9 2
24 9 11 11 13 3 16 0 9 9 9 0 9 2 7 13 0 2 16 3 13 3 1 15 2
13 9 13 0 9 0 1 0 9 2 9 7 9 2
18 3 0 13 7 0 9 2 0 1 10 2 3 16 1 0 2 9 2
27 3 10 9 1 10 9 13 0 9 2 1 15 15 1 9 9 13 0 0 9 2 15 13 3 1 15 2
72 9 9 13 3 9 0 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 2 13 7 7 9 0 2 11 2 11 2 11 2 11 2 11 2 7 0 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 2
5 9 13 0 9 2
12 0 9 3 13 2 16 0 0 9 13 9 2
26 0 9 2 3 3 15 13 11 11 2 13 10 0 9 3 1 9 2 3 1 3 0 0 9 9 2
25 0 9 2 0 3 9 0 9 9 1 9 2 13 3 0 9 9 1 0 2 7 0 2 9 2
27 0 0 9 15 1 15 13 1 10 9 3 2 16 9 9 9 2 3 1 9 0 9 2 9 11 2 2
35 15 3 13 9 7 1 9 0 9 7 3 15 3 13 0 9 1 9 0 9 2 3 2 14 3 0 9 2 9 9 2 0 9 2 2
2 11 11
19 11 11 7 11 11 4 13 0 9 3 1 0 9 0 2 11 7 11 2
21 9 0 9 0 9 2 11 2 9 0 2 4 13 1 9 9 9 1 0 9 2
20 9 13 1 9 1 9 11 2 1 11 7 1 9 9 7 1 9 10 9 2
5 9 1 9 7 9
24 9 0 9 1 9 2 9 2 11 11 13 1 12 2 7 12 2 9 1 0 0 9 11 2
16 12 2 9 13 3 3 9 9 1 0 9 0 9 1 11 2
36 1 9 4 13 3 0 9 0 0 9 2 3 0 9 0 9 2 13 4 9 1 0 9 9 0 9 2 0 9 13 11 1 9 12 2 2
24 9 4 13 9 0 0 9 0 9 2 15 13 12 2 9 1 9 7 4 13 14 1 11 2
23 1 9 1 0 9 15 9 13 1 9 14 1 11 2 3 13 0 0 9 1 0 9 2
10 13 4 1 0 9 0 9 7 11 2
7 9 9 4 13 0 9 2
11 9 13 9 2 13 11 2 7 0 9 2
13 9 11 11 1 9 0 9 13 0 2 11 9 2
39 0 0 9 15 4 13 1 0 0 9 2 0 0 9 2 0 9 2 7 9 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 7 0 2 2
7 3 1 15 13 7 9 2
29 9 4 13 1 9 9 9 10 9 7 9 1 9 1 0 9 2 12 2 9 2 13 1 9 9 9 1 9 2
3 2 11 2
4 11 1 11 2
21 1 9 0 9 0 11 1 9 11 11 15 1 9 13 0 9 1 0 9 11 2
12 3 4 13 4 1 0 9 0 9 3 13 2
19 1 9 13 9 11 11 7 0 9 2 15 16 0 0 9 13 11 11 2
16 9 11 4 13 1 9 2 7 9 0 9 13 9 0 9 2
16 16 1 10 9 13 9 16 1 9 0 9 2 13 7 9 2
16 9 3 13 14 1 0 9 2 16 4 15 15 13 1 9 2
3 2 11 2
6 0 9 13 9 11 11
9 0 9 0 9 13 2 9 9 2
2 9 9
2 11 11
14 9 2 0 2 12 2 13 0 9 2 13 1 9 0
26 1 9 2 16 2 13 9 13 9 2 2 13 0 0 9 0 9 2 16 13 2 9 10 9 2 2
20 1 15 13 0 9 2 1 15 13 9 0 0 0 9 0 9 1 9 12 2
9 1 0 0 9 15 13 9 9 2
9 3 3 4 0 9 0 9 13 2
6 13 15 3 1 9 2
39 1 0 9 9 15 1 15 13 0 9 2 13 9 0 9 2 9 1 0 9 9 13 2 3 13 12 9 2 3 12 2 1 15 9 0 12 7 12 2
19 0 0 9 7 13 9 0 0 9 1 9 0 9 2 0 9 0 9 2
46 1 0 9 2 12 9 1 9 12 2 12 2 2 3 1 9 13 0 9 7 9 2 3 9 0 1 9 1 12 9 13 1 9 1 12 2 2 9 7 3 0 9 13 1 9 2
23 9 3 13 0 0 9 2 0 9 1 0 9 2 10 9 13 9 2 0 9 0 9 2
22 3 3 15 1 9 0 9 13 15 2 0 2 2 15 9 9 13 9 0 0 9 2
11 9 7 13 0 9 2 0 0 0 9 2
17 0 13 3 0 9 9 2 15 15 13 1 9 2 9 7 9 2
23 16 0 9 1 9 9 12 9 2 9 1 9 13 3 12 9 2 7 0 9 13 9 2
34 0 9 15 1 9 9 13 1 9 9 7 0 9 0 9 2 1 15 15 13 0 9 2 3 13 9 1 9 2 0 1 0 9 2
25 1 9 9 13 3 13 14 9 0 1 12 2 12 9 9 7 0 1 9 7 3 0 1 9 2
8 0 9 0 9 13 1 9 2
22 10 9 1 9 9 9 0 9 9 11 2 11 7 1 0 0 9 13 1 0 9 2
33 9 0 1 0 9 0 9 2 1 15 9 3 13 9 2 0 9 7 9 2 15 7 1 9 13 9 0 9 1 9 11 11 2
17 9 14 0 13 9 3 0 9 11 11 1 12 2 9 10 9 2
25 9 13 13 0 9 0 1 3 0 0 2 0 7 0 9 1 9 9 7 9 0 9 7 9 2
20 1 12 9 13 4 13 1 9 9 1 9 2 1 9 13 9 9 0 9 2
24 9 13 1 9 13 16 0 9 0 7 0 9 2 10 9 16 12 1 0 9 0 9 9 2
28 1 0 15 0 9 9 15 13 0 0 0 9 2 15 0 9 13 13 1 0 0 9 0 0 9 1 9 2
15 1 9 2 15 13 0 9 2 15 9 9 0 9 13 2
39 3 3 13 9 0 9 2 1 15 13 1 0 7 9 1 9 10 9 2 11 2 11 7 0 2 2 15 1 9 9 2 15 14 3 3 0 2 13 2
10 1 0 9 15 7 13 13 9 0 2
34 16 4 1 0 9 9 13 1 0 9 0 7 0 2 1 15 1 11 13 9 11 11 2 11 2 0 10 9 1 11 7 0 11 2
20 9 9 9 2 0 9 9 9 13 12 3 0 9 1 9 0 9 9 11 2
33 1 0 9 13 9 0 1 0 3 9 2 3 0 9 12 9 2 9 1 0 9 7 9 2 9 0 9 7 0 9 1 11 2
18 0 9 9 13 3 9 9 2 16 13 0 9 13 3 16 0 9 2
43 9 0 0 9 0 9 13 9 1 3 0 9 0 9 10 9 2 11 11 2 9 11 11 11 11 2 2 11 11 2 9 11 11 2 7 11 11 2 9 11 11 2 2
15 9 0 12 13 1 0 0 9 2 15 3 13 9 9 2
25 12 9 11 11 2 11 2 7 11 11 2 11 2 0 9 13 10 0 9 3 1 0 0 9 2
19 11 3 3 13 0 9 2 1 15 7 13 0 0 9 2 13 9 2 2
30 9 0 9 11 11 13 3 12 2 9 2 12 2 2 0 9 1 9 2 12 2 7 9 1 9 11 2 12 2 2
35 0 9 2 0 9 2 0 9 11 7 0 9 2 7 9 2 11 11 2 11 11 7 11 11 2 13 9 0 7 0 9 0 0 9 2
14 3 0 9 4 13 1 9 0 7 0 9 11 11 2
41 9 0 1 9 12 2 12 7 0 1 9 12 2 12 2 3 0 9 2 1 11 11 7 11 11 2 7 0 9 2 13 7 0 7 15 1 15 10 0 9 2
19 9 1 0 9 7 0 9 13 3 1 0 9 7 0 9 1 0 9 2
16 9 1 9 2 9 7 9 13 1 0 9 9 12 0 9 2
40 9 15 13 1 9 7 9 2 7 13 1 9 3 2 14 3 16 9 7 9 7 1 0 2 3 15 0 9 2 9 2 11 11 2 9 2 11 11 2 2
22 0 9 9 13 11 2 0 9 1 0 0 9 2 15 13 9 0 9 7 0 9 2
29 9 0 9 7 11 3 3 3 13 0 9 12 9 1 0 9 1 0 9 11 11 1 9 12 2 9 9 2 2
30 3 0 7 3 0 0 9 3 13 0 11 1 9 2 0 9 2 7 12 0 9 2 6 6 2 2 9 7 0 2
2 11 11
5 9 16 0 1 9
8 9 13 0 9 2 13 11 11
2 9 9
30 9 11 11 2 12 2 3 13 1 12 9 2 3 3 9 1 9 1 9 0 9 13 9 7 9 11 11 1 9 2
11 0 9 15 13 9 9 9 1 0 11 2
2 11 11
6 3 4 10 9 13 2
25 13 4 15 3 13 2 16 4 15 1 10 9 13 3 2 16 1 0 9 13 0 9 1 11 2
13 7 11 13 1 15 2 15 3 13 2 0 9 2
15 1 15 15 13 1 0 9 9 9 7 9 9 15 15 2
19 1 10 9 13 3 0 0 9 2 3 3 16 1 10 9 2 1 9 2
16 9 13 1 9 0 9 7 13 4 2 16 4 10 9 13 2
28 7 15 4 13 2 16 4 15 9 3 13 2 16 4 2 3 13 11 2 13 9 9 2 7 10 0 9 2
7 16 4 1 15 13 9 2
20 16 4 13 1 9 2 9 7 3 7 1 0 9 2 15 15 3 3 13 2
11 10 0 9 13 2 16 4 13 0 9 2
6 3 2 3 7 3 2
31 3 1 12 1 11 12 13 9 10 0 9 9 13 10 9 2 0 11 11 2 9 2 10 9 13 9 7 9 2 2 2
16 3 15 13 2 16 9 7 0 9 13 9 16 0 1 9 2
18 9 15 13 13 2 13 13 7 3 15 15 13 1 9 9 0 9 2
10 16 9 0 9 4 13 15 0 9 2
33 13 4 15 13 1 9 2 16 10 0 9 2 15 4 15 13 3 1 9 2 13 1 9 7 13 9 0 1 0 9 3 9 2
33 0 9 13 3 10 2 14 12 2 7 15 15 13 13 2 3 15 6 15 13 2 16 13 9 7 3 1 10 9 13 1 9 2
17 1 0 9 11 9 1 0 9 13 14 0 2 7 7 0 9 2
7 3 15 10 0 9 13 2
31 16 4 3 13 7 13 9 0 9 2 13 4 1 9 9 13 2 16 13 3 0 0 9 2 1 15 0 2 1 9 2
11 1 15 15 7 13 1 9 3 9 9 2
10 7 15 3 2 3 14 1 0 9 2
15 16 13 0 9 10 9 2 3 13 1 10 9 3 0 2
15 13 3 2 10 0 9 2 9 7 9 15 1 15 13 2
18 16 13 13 10 9 1 9 9 2 13 15 0 9 9 1 9 0 2
23 7 16 15 0 13 1 15 0 2 13 13 9 9 1 15 2 9 7 9 2 3 9 2
4 9 2 11 11
4 9 11 11 2
4 0 11 1 11
23 9 2 0 9 1 11 11 13 1 9 9 11 1 9 1 0 9 11 11 1 9 12 2
18 9 9 13 9 9 11 11 2 1 9 11 11 9 13 9 11 11 2
27 11 1 9 13 1 9 0 9 0 9 7 13 3 1 0 11 9 2 15 0 0 9 13 1 0 9 2
19 0 9 13 0 0 9 1 0 9 2 0 0 9 2 0 15 1 9 2
31 15 13 13 9 0 9 9 2 9 7 0 0 9 2 1 15 15 13 9 9 2 15 11 13 1 10 0 9 1 11 2
20 10 9 3 3 13 1 9 3 0 1 9 9 2 3 0 2 3 3 0 2
32 9 9 2 1 15 15 9 7 9 13 3 3 2 16 13 0 2 13 3 1 9 9 0 1 9 7 9 0 1 9 9 2
14 13 15 0 9 2 9 3 0 0 7 0 9 9 2
7 0 9 13 3 1 9 2
22 15 15 2 3 15 13 2 1 9 9 13 7 10 9 13 9 9 7 0 0 9 2
31 1 0 9 15 13 1 9 0 9 2 1 0 11 11 16 9 11 2 13 11 11 2 7 3 1 11 11 1 0 9 2
29 10 3 0 11 13 0 9 0 9 1 3 0 9 0 9 7 10 0 9 13 1 0 9 16 9 3 0 9 2
35 9 0 0 9 3 13 3 0 9 2 3 11 11 16 0 11 2 11 11 16 11 11 2 0 0 9 2 7 11 11 16 0 9 11 2
23 0 9 13 3 15 0 9 2 0 1 9 1 9 10 0 9 11 11 2 11 11 2 2
22 0 9 9 2 15 10 9 7 0 9 13 9 1 0 9 2 13 0 9 11 11 2
27 9 7 0 9 13 9 7 9 3 3 0 2 16 3 1 0 9 3 13 10 0 9 2 9 3 0 2
19 15 13 7 14 0 9 2 15 13 13 0 0 9 1 0 7 0 9 2
2 11 11
28 9 2 11 11 2 3 16 11 11 2 2 11 11 2 9 11 2 7 11 11 2 11 2 1 9 11 1 9
3 9 11 11
5 9 1 9 13 11
8 0 9 11 1 11 13 11 11
7 11 1 11 2 11 2 2
27 9 1 0 0 9 1 11 2 15 13 1 0 9 1 9 9 1 11 2 13 11 11 1 9 11 11 2
9 9 0 9 13 11 11 1 11 2
6 3 13 9 0 9 2
29 0 9 13 0 9 2 1 15 13 0 13 9 2 15 15 1 9 11 7 0 9 13 3 1 12 1 12 9 2
13 1 9 3 4 13 0 9 2 3 1 0 9 2
4 9 1 0 9
12 11 13 1 2 9 2 7 1 0 11 15 13
2 9 9
5 11 2 11 2 2
36 3 13 0 9 11 11 1 9 9 11 1 11 11 2 16 4 3 3 13 1 0 9 1 9 1 0 11 2 10 0 9 13 12 2 12 2
27 1 0 9 15 13 2 16 13 1 9 9 2 7 1 11 0 11 1 9 9 2 3 1 0 0 9 2
28 2 13 4 13 9 7 13 9 2 16 4 1 9 13 3 1 0 9 2 2 13 3 10 9 11 2 11 2
17 13 15 1 0 2 16 3 0 9 9 15 3 1 12 9 13 2
22 9 2 1 15 13 0 9 1 9 7 9 12 9 2 13 3 1 12 9 1 9 2
24 12 13 0 9 9 7 14 12 15 1 9 1 12 9 13 1 9 0 9 9 9 1 9 2
35 9 0 9 9 1 9 2 15 15 13 13 12 2 7 12 2 12 2 1 0 9 2 13 0 9 2 9 11 2 1 0 9 1 9 2
3 3 1 9
5 9 9 2 11 2
8 12 9 2 2 11 2 11 2
7 0 11 1 9 1 0 11
2 9 11
2 11 11
2 9 9
1 9
3 0 11 2
11 0 9 12 2 9 9 14 2 0 11 2
1 9
7 9 2 12 2 7 12 2
4 11 2 12 2
4 11 2 12 2
2 11 2
3 9 11 2
11 9 2 11 2 11 2 11 2 11 2 2
26 11 2 11 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 11 2 11 2
26 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2
12 0 9 2 12 2 9 2 11 2 11 0 2
4 11 2 12 2
4 11 2 12 2
5 11 11 2 12 2
4 11 2 12 2
4 11 2 12 2
4 11 2 12 2
4 11 2 12 2
2 11 2
1 9
9 9 1 9 1 9 2 9 9 2
2 12 2
4 9 13 11 2
3 13 4 2
5 0 9 1 9 13
3 0 11 2
50 3 0 9 0 11 11 2 15 13 1 12 2 9 9 14 0 11 1 9 11 12 2 12 1 9 2 13 1 0 9 0 9 1 11 11 12 2 12 7 13 15 1 9 0 9 9 12 2 12 2
27 1 0 9 15 13 3 0 9 11 11 2 15 13 1 12 2 9 0 9 2 7 1 9 9 15 13 2
19 1 0 11 13 11 11 12 2 12 2 16 15 13 1 9 1 0 9 2
16 1 12 2 12 13 3 1 9 0 9 11 11 7 11 11 2
10 1 0 9 13 3 14 13 11 11 2
22 1 0 9 1 0 11 13 0 9 11 11 2 15 13 12 1 12 0 9 0 11 2
5 0 9 13 0 9
6 9 1 11 13 9 2
7 0 13 9 2 13 11 11
2 9 9
9 11 2 11 2 11 2 11 2 2
10 2 9 13 3 0 7 13 15 9 2
15 10 9 13 0 9 7 13 0 2 16 15 15 0 13 2
19 2 3 9 2 0 2 9 9 12 11 11 1 0 9 0 9 0 11 2
25 0 9 9 7 9 10 9 13 11 0 11 2 16 1 0 9 13 9 11 7 13 1 0 9 2
23 1 0 0 9 11 11 11 15 9 1 11 13 0 9 7 1 11 4 13 0 0 9 2
36 0 9 13 3 0 2 0 11 11 11 13 1 9 11 1 9 12 3 1 0 9 2 11 11 11 13 9 9 2 1 15 4 1 9 13 2
11 2 13 4 2 16 11 13 13 14 9 2
12 16 9 9 12 1 15 7 9 13 3 13 2
19 1 9 7 9 13 14 0 9 2 2 13 1 0 9 1 9 11 11 2
13 2 13 4 15 3 13 2 16 4 13 1 9 2
26 13 15 3 0 2 3 4 3 3 3 1 9 13 2 2 13 11 2 3 1 9 13 3 1 9 2
36 15 11 15 13 9 9 13 7 1 0 9 11 1 11 15 13 1 9 9 2 14 13 1 11 1 0 9 1 0 9 9 1 9 10 9 2
50 2 10 11 2 11 13 0 9 2 13 3 7 0 11 4 13 14 13 2 2 13 15 1 9 11 7 13 15 1 0 9 1 9 2 2 0 9 7 9 11 15 13 2 16 1 0 9 13 9 2
6 0 0 9 3 13 2
45 2 0 9 13 1 9 7 11 11 2 0 9 11 2 2 13 4 1 11 7 1 0 9 4 15 13 2 16 10 9 1 10 9 3 13 9 2 1 9 3 15 3 13 2 2
20 9 1 9 0 9 13 3 2 1 9 9 9 9 15 13 0 9 11 11 2
23 1 9 11 13 11 3 0 9 2 7 1 9 3 1 9 13 9 12 9 1 0 9 2
16 3 0 9 13 13 1 9 0 9 2 15 13 13 0 9 2
19 9 13 3 9 2 16 11 2 16 4 15 13 9 2 3 13 10 9 2
27 0 9 9 11 11 11 15 3 3 16 11 11 11 13 1 9 2 16 1 11 4 15 3 3 13 13 2
9 9 4 3 3 3 9 9 13 2
31 3 15 9 13 13 1 0 9 1 0 9 2 9 0 9 2 9 2 15 15 13 7 1 9 11 1 11 1 0 11 2
13 11 3 16 9 9 1 11 15 3 1 9 13 2
34 15 3 13 7 0 9 9 11 11 2 15 1 9 9 11 3 1 9 11 11 13 2 16 3 13 1 9 0 1 9 1 9 9 2
13 2 9 13 3 3 0 2 16 15 13 10 9 2
22 9 4 15 15 13 13 3 2 7 15 15 13 2 2 13 15 11 2 0 0 9 2
12 12 15 1 9 13 1 9 7 13 15 9 2
28 3 11 4 15 13 13 9 9 9 2 1 15 3 1 9 1 9 1 9 1 9 11 13 11 11 3 11 2
7 2 9 3 1 15 13 2
23 13 13 2 16 9 1 11 13 0 9 2 7 13 9 9 12 2 7 0 9 13 9 2
13 9 4 15 13 13 3 7 13 4 15 13 11 2
35 2 3 16 11 13 7 11 1 0 9 9 2 2 9 1 15 13 3 10 9 9 2 13 15 1 15 2 16 4 4 10 9 3 13 2
61 3 13 1 15 9 9 2 9 13 1 0 9 0 9 9 2 15 4 3 13 7 13 13 0 9 9 2 2 13 15 11 7 13 15 1 10 0 9 2 2 9 12 13 3 0 9 7 9 15 13 3 13 9 2 16 15 13 3 10 9 2
8 3 13 3 0 9 2 14 2
9 11 13 0 9 2 15 4 13 2
11 13 0 7 13 1 9 0 9 3 15 2
20 2 1 0 9 0 9 13 0 9 11 11 9 0 9 1 9 9 0 9 2
27 12 9 4 1 11 1 15 0 9 1 9 9 13 0 9 7 15 0 0 2 0 7 0 9 4 13 2
43 9 11 3 13 9 12 0 9 9 7 13 9 0 9 1 11 2 16 4 0 9 4 3 3 13 1 10 0 9 2 15 4 13 13 13 3 3 3 1 3 0 9 2
21 2 1 11 13 15 0 9 2 13 9 0 9 2 2 13 0 0 9 11 11 2
3 11 13 13
6 9 1 11 0 0 9
2 9 9
7 11 1 11 2 11 2 2
71 2 13 0 1 15 2 16 4 13 3 0 9 2 7 13 0 2 16 15 3 13 13 1 9 9 7 13 15 3 9 7 13 2 2 13 0 9 11 11 2 9 11 11 2 15 15 16 0 1 0 0 9 13 1 9 9 0 9 1 11 1 9 12 2 1 9 1 11 1 11 2
27 9 13 1 9 0 9 1 0 9 1 11 11 3 12 2 12 1 9 2 7 0 12 9 13 1 9 2
18 2 0 9 1 15 15 11 7 13 1 9 14 2 7 13 0 9 2
9 13 15 1 0 9 1 0 9 2
10 16 15 4 13 7 15 7 11 11 2
4 15 13 0 2
14 13 3 3 3 12 9 2 9 3 13 7 1 15 2
24 3 4 7 13 1 10 9 1 0 9 2 3 4 13 10 9 2 7 1 9 14 0 2 2
25 11 11 13 1 9 13 15 1 11 11 2 15 13 3 3 2 16 3 1 15 9 1 9 13 2
6 2 15 3 13 9 2
10 9 13 9 2 13 3 9 1 15 2
23 3 3 13 13 9 2 0 9 7 9 9 9 11 11 11 11 2 9 2 9 2 2 2
38 2 11 13 1 0 9 1 11 1 11 1 11 1 11 7 1 12 9 0 9 9 1 11 1 11 2 12 12 12 9 1 0 9 10 9 1 11 2
10 2 13 4 15 13 2 3 4 13 2
9 7 3 13 13 2 3 15 13 2
7 13 1 9 2 2 2 2
3 9 1 9
5 11 2 11 2 2
30 1 9 11 15 13 0 0 9 0 0 9 3 0 9 9 11 2 1 15 13 13 9 12 2 7 12 2 0 9 2
17 3 0 0 9 13 9 12 9 9 9 0 9 12 2 12 9 2
33 11 11 2 9 0 9 9 12 2 3 13 2 16 1 9 9 13 2 2 13 9 2 15 15 13 9 7 1 10 9 4 13 2
12 13 15 0 2 16 4 3 15 11 13 2 2
3 9 13 11
4 11 1 11 2
33 1 9 13 13 10 9 0 9 1 11 2 9 4 1 9 13 2 2 16 11 1 9 12 2 12 1 11 15 3 13 1 9 2
15 1 15 15 13 13 0 9 2 15 13 12 2 12 11 2
17 16 3 13 11 3 1 12 9 0 11 2 13 3 1 9 11 2
4 11 2 12 2
4 11 2 12 2
4 11 2 12 2
4 11 2 12 2
2 11 2
17 9 2 11 2 11 2 12 11 2 2 2 11 2 11 2 2 2
4 11 2 12 2
4 11 2 12 2
4 11 2 12 2
2 11 2
4 11 2 12 2
4 11 2 12 2
4 11 2 12 2
4 11 2 12 2
4 11 2 12 2
4 11 2 12 2
2 11 2
14 1 9 1 11 0 9 13 1 9 1 11 12 2 12
2 9 9
29 0 0 9 13 1 10 0 9 1 0 9 1 12 2 9 9 1 11 1 11 1 0 9 1 11 12 2 12 2
22 15 13 1 15 2 16 1 0 9 13 1 9 1 12 9 1 11 2 9 9 9 2
18 0 9 13 2 11 2 11 2 11 2 11 7 11 2 11 2 11 2
22 1 9 4 13 11 1 0 1 0 9 11 2 0 11 2 11 13 1 9 9 2 2
9 0 9 11 1 11 1 11 11 11
31 10 9 0 12 15 13 2 16 11 11 2 9 1 15 13 1 0 9 2 13 3 1 9 1 10 9 0 9 1 11 2
25 9 0 9 0 9 13 7 0 9 1 12 2 9 2 3 11 13 1 0 9 9 1 9 11 2
21 1 12 9 3 13 10 9 9 13 2 7 11 1 11 13 1 15 0 0 9 2
9 2 9 2 1 11 7 13 3 2
18 1 9 13 13 2 1 0 9 0 11 13 0 9 1 0 0 9 2
23 1 9 13 7 9 9 2 13 4 1 0 9 7 1 9 1 0 9 3 13 1 9 2
37 9 1 9 12 3 13 9 1 0 9 7 16 1 12 2 9 13 11 1 9 1 11 13 1 9 1 9 9 2 13 11 3 1 12 2 12 2
15 0 9 13 1 9 1 0 12 9 13 3 0 9 9 2
17 1 15 7 13 14 11 0 9 7 3 0 9 1 9 11 11 2
10 0 9 3 3 1 0 9 13 11 2
4 11 2 12 2
4 11 2 12 2
4 11 2 12 2
4 11 2 12 2
2 11 2
8 9 2 11 2 11 2 2 2
12 11 2 11 2 11 2 11 2 11 2 11 2
6 11 2 11 2 11 2
18 0 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2
2 11 2
4 11 2 12 2
2 11 2
2 11 2
2 11 2
4 9 2 11 2
4 11 2 12 2
2 11 2
13 0 9 9 13 0 2 0 9 9 13 3 0 2
3 2 9 2
21 1 9 0 9 13 3 0 9 9 12 0 9 2 15 13 12 9 1 0 9 2
10 1 9 13 1 11 3 2 3 9 2
23 0 9 12 7 12 9 2 2 1 0 9 7 0 2 0 0 12 7 12 9 2 9 2
11 1 12 9 1 9 1 12 9 2 9 2
4 0 0 9 2
15 1 9 7 1 9 13 3 3 2 3 9 9 1 9 2
22 0 0 9 1 9 12 7 12 9 2 9 2 2 1 9 12 7 12 9 2 9 2
13 0 0 9 1 12 9 12 7 12 9 2 9 2
12 9 13 1 9 1 12 7 13 1 12 9 2
10 9 13 1 12 7 13 1 12 9 2
26 0 9 12 2 9 2 0 9 12 9 2 9 1 9 12 2 0 9 12 9 2 9 1 9 12 2
9 0 0 9 13 12 9 2 9 2
9 9 1 0 11 13 9 0 9 2
9 1 10 9 13 0 9 1 9 2
13 4 13 0 7 0 9 12 7 12 9 2 9 2
5 0 11 2 0 11
11 9 11 15 1 9 4 13 3 1 12 9
2 9 9
6 0 11 2 11 2 2
19 9 12 2 12 1 9 0 11 13 11 10 9 0 0 9 12 2 12 2
31 1 9 15 13 0 9 1 0 11 7 1 0 0 9 15 1 0 12 9 2 3 13 14 12 1 11 2 13 12 9 2
6 2 3 13 15 0 2
32 1 9 15 13 13 2 16 1 0 12 9 13 3 11 7 13 1 11 2 2 13 9 11 11 1 9 9 1 9 0 9 2
28 1 9 10 9 13 7 0 2 2 1 9 4 1 1 9 11 7 11 13 9 2 1 12 13 3 3 0 2
16 1 9 2 15 4 1 12 2 9 13 2 4 15 9 13 2
26 2 1 9 9 15 13 3 1 12 2 9 2 16 0 11 1 9 12 2 12 3 13 0 0 9 2
21 2 10 9 15 3 13 7 13 4 14 3 1 9 9 2 2 13 0 9 11 2
13 2 13 1 11 13 10 9 2 7 15 13 13 2
10 14 4 15 0 9 9 1 9 13 2
21 1 11 7 11 13 10 9 0 2 7 1 9 0 9 4 3 1 9 13 2 2
4 3 9 9 13
2 9 9
5 11 2 11 2 2
28 3 1 0 0 9 16 1 15 0 14 13 9 11 7 11 2 15 13 0 9 14 1 3 0 11 7 11 2
9 3 13 1 9 2 1 15 13 2
15 11 13 9 12 2 12 1 11 1 11 1 3 0 9 2
24 0 9 9 2 15 15 13 1 9 2 13 0 12 9 2 16 15 3 13 9 11 7 11 2
5 9 15 13 13 2
17 2 3 1 0 9 4 13 3 7 10 9 4 15 13 3 15 2
28 13 4 13 14 1 9 2 16 4 15 9 13 1 9 2 15 4 14 13 9 2 2 13 3 0 9 11 2
23 1 0 9 15 11 13 1 11 1 0 9 2 15 3 1 9 13 2 12 2 12 2 2
36 9 11 2 11 2 11 2 11 2 11 4 13 3 1 9 2 9 12 9 2 7 13 15 1 15 0 11 2 11 7 9 2 1 15 13 2
11 2 13 4 15 2 16 4 13 9 0 2
23 14 15 1 9 9 13 0 2 16 4 13 1 9 9 2 2 13 9 2 9 2 11 2
30 1 11 15 3 13 9 1 0 9 2 7 1 0 9 15 13 9 9 1 0 9 2 15 13 0 9 13 1 11 2
12 3 13 4 3 9 13 9 11 11 11 11 2
20 2 1 11 13 3 1 11 1 12 12 9 2 3 4 13 1 12 12 3 2
15 1 9 13 9 1 0 9 11 2 2 13 9 11 11 2
3 11 15 13
5 11 2 11 2 2
28 0 9 11 1 11 1 12 2 0 9 13 1 9 7 9 0 11 11 2 15 15 1 9 13 0 9 9 2
26 2 13 4 1 15 1 11 7 13 15 11 2 2 13 0 9 2 15 15 1 10 9 13 1 9 2
19 2 3 0 9 3 1 9 15 13 1 9 7 13 4 1 9 9 13 2
26 2 3 11 13 9 2 1 12 9 4 13 13 1 9 7 1 0 12 9 3 3 1 9 1 9 2
29 2 1 9 15 13 14 1 9 2 3 13 3 9 13 15 3 10 9 2 9 9 11 2 9 2 9 2 2 2
22 2 3 7 11 13 2 0 9 13 16 10 9 11 2 1 9 13 14 3 2 2 2
9 11 11 13 0 9 11 14 1 9
5 9 11 11 2 11
4 9 12 2 9
18 1 9 13 9 9 11 11 1 9 12 2 9 1 0 9 1 11 2
3 2 11 2
3 0 0 9
7 9 1 9 9 15 13 9
2 9 9
9 11 2 11 2 11 2 11 2 2
36 9 1 9 9 9 1 11 13 11 0 9 2 3 13 0 9 2 9 7 9 2 2 13 0 9 1 0 9 7 13 15 1 0 9 11 2
20 1 0 9 2 3 0 9 11 2 13 3 11 1 11 2 3 13 7 0 2
37 11 15 3 1 0 9 13 13 1 9 0 9 11 7 11 2 15 13 13 7 3 11 15 3 3 13 2 16 13 9 1 10 9 3 3 0 2
23 3 3 15 13 10 0 9 1 11 1 0 9 9 2 1 15 13 9 0 9 1 11 2
9 9 1 11 11 2 0 9 0 9
32 3 13 0 9 11 11 2 9 1 11 11 7 9 1 11 2 7 0 9 0 9 1 9 1 9 1 9 11 11 1 11 2
10 2 3 4 15 13 1 9 1 11 2
26 1 0 9 15 13 12 2 11 2 11 2 11 2 11 2 11 2 11 7 11 2 1 11 13 9 2
21 11 15 15 3 13 2 7 3 13 1 15 12 9 7 13 15 4 14 1 9 2
11 3 13 2 15 13 1 9 0 7 0 2
14 2 10 0 9 3 13 11 2 15 13 1 0 9 2
23 2 1 11 11 13 1 11 1 9 0 9 2 3 1 11 13 0 11 2 15 3 13 2
16 11 13 0 9 2 7 13 15 1 9 7 3 13 3 9 2
12 2 13 15 9 11 2 11 7 9 1 9 2
21 2 3 4 9 0 9 1 11 13 12 9 2 7 3 11 3 13 1 0 9 2
19 9 13 1 15 0 2 11 13 3 0 9 7 11 1 10 9 3 13 2
12 2 3 4 13 1 0 9 1 9 1 11 2
16 2 13 13 0 9 1 10 9 2 16 9 15 13 4 2 2
3 2 11 2
13 3 1 11 2 9 0 9 2 11 11 2 0 9
7 0 9 13 1 0 9 9
5 11 2 11 2 2
21 1 0 9 0 9 15 12 3 0 9 9 0 9 0 9 13 11 13 9 9 2
9 13 4 15 3 13 3 10 9 2
9 11 15 3 13 9 9 11 11 2
20 1 10 0 9 3 9 13 2 16 15 9 9 9 13 9 11 13 0 9 2
8 9 4 15 13 13 9 9 2
23 2 0 4 15 1 9 13 9 0 9 2 16 15 13 0 16 9 2 2 13 9 11 2
11 9 13 9 1 9 0 9 1 12 9 2
16 9 9 15 1 9 2 1 0 9 9 2 13 1 12 9 2
12 13 2 14 15 7 0 2 13 13 7 3 2
19 9 15 7 13 13 3 7 9 9 1 9 9 13 2 16 13 7 3 2
10 2 3 0 0 9 13 7 1 9 2
20 9 3 13 3 2 13 15 1 0 9 2 2 13 11 2 11 1 9 9 2
9 0 9 13 14 12 9 1 12 9
5 11 2 11 2 2
15 1 9 1 9 1 0 9 1 11 13 7 3 0 9 2
30 3 1 0 9 11 1 11 15 15 13 12 2 1 0 1 0 0 9 12 2 1 0 9 0 9 1 11 3 12 2
27 3 4 1 9 9 11 7 11 13 0 9 2 1 10 9 13 13 12 9 1 0 9 3 1 9 0 2
16 0 9 0 1 0 9 13 0 7 3 2 3 7 4 13 2
22 0 9 1 11 2 15 13 3 0 9 2 15 4 13 9 1 11 7 1 11 13 2
6 9 9 13 9 15 2
27 0 0 9 4 13 1 12 9 7 12 9 12 9 2 3 9 2 15 13 1 12 0 9 1 0 9 2
33 1 12 2 0 9 13 0 9 2 15 3 13 1 0 9 2 12 7 1 0 9 15 10 9 13 14 3 2 3 1 12 9 2
23 15 2 15 13 1 0 9 1 0 9 12 2 12 2 7 1 9 13 12 7 12 12 2
33 9 9 3 1 9 9 1 12 9 3 13 14 3 0 9 2 7 7 0 0 9 2 16 13 9 7 9 1 9 9 0 9 2
18 3 15 13 13 2 16 4 12 2 0 13 0 9 1 9 0 9 2
7 15 3 13 12 9 3 2
9 1 0 9 1 11 7 9 13 2
18 9 3 9 13 12 9 3 7 1 0 9 4 13 13 7 0 9 2
17 3 3 1 0 9 11 13 1 0 9 3 16 1 0 0 9 2
14 16 4 13 2 13 12 7 12 12 9 3 1 9 2
8 11 2 11 2 1 11 4 13
2 9 9
7 11 2 11 2 11 2 2
39 9 11 11 3 13 9 9 2 16 1 9 1 9 9 11 11 7 9 9 11 11 13 0 9 1 9 9 9 9 0 9 2 11 2 11 11 1 9 2
5 2 13 1 9 2
17 9 11 1 15 10 1 15 13 2 2 13 0 0 9 11 11 2
9 11 13 4 13 1 0 9 9 2
23 1 10 9 9 11 13 2 16 9 9 13 3 10 0 9 1 9 11 2 7 11 13 2
50 1 10 9 1 9 0 9 11 2 11 2 11 2 11 7 11 2 11 15 13 2 16 11 2 11 13 1 9 2 16 12 9 9 11 2 15 3 0 9 13 0 9 1 10 9 2 13 0 9 2
12 9 10 9 9 3 13 1 0 9 11 13 2
69 9 9 0 0 9 11 13 2 9 9 11 2 11 2 9 2 2 10 9 11 11 2 9 9 9 11 11 2 9 9 9 7 9 11 11 2 9 0 0 9 11 11 2 9 9 9 11 11 2 9 11 11 2 11 2 0 9 0 9 11 11 11 7 11 11 1 9 9 2
10 1 9 9 11 13 12 9 9 9 2
10 0 9 11 1 9 9 13 9 9 2
5 9 11 15 9 13
2 11 2
31 3 12 9 9 13 0 9 1 9 9 0 9 1 0 0 0 9 1 0 9 2 15 13 3 1 11 7 11 1 11 2
17 13 15 3 0 9 1 0 9 2 9 0 9 0 9 11 11 2
37 1 9 13 0 9 12 12 9 2 1 9 12 9 2 1 9 12 9 7 1 9 12 9 9 2 7 15 2 3 1 0 9 2 2 13 11 2
13 13 15 3 1 15 0 9 0 12 2 9 12 2
11 0 9 7 11 10 9 1 9 11 13 2
13 11 13 2 16 15 12 0 9 13 1 0 9 2
18 3 3 3 4 0 9 9 1 0 0 9 13 2 3 3 13 13 2
5 0 0 9 13 9
2 11 2
27 0 9 0 9 11 11 15 13 16 9 0 9 7 9 2 15 13 3 0 1 15 0 16 0 1 15 2
15 1 9 1 9 0 9 1 0 11 15 3 13 9 11 2
47 1 9 1 9 9 2 10 9 13 2 16 10 9 13 3 0 2 11 1 10 9 2 15 1 11 13 1 9 9 1 11 2 9 13 10 9 7 10 0 9 7 13 2 16 13 0 2
20 13 2 0 9 9 2 0 9 2 9 7 0 9 9 2 9 7 9 2 2
24 1 0 9 0 11 13 2 16 4 3 13 9 7 16 3 13 1 9 9 2 15 3 13 2
21 16 9 13 15 2 16 15 1 9 12 1 0 9 13 1 11 11 16 10 9 2
21 11 13 2 16 15 13 13 2 15 15 13 1 15 13 1 9 0 9 16 9 2
22 3 15 13 11 2 16 10 0 9 1 9 13 1 9 2 16 0 1 0 9 2 2
15 3 11 10 9 13 2 2 11 7 15 4 3 3 13 2
25 2 0 9 13 2 16 0 9 13 1 11 11 2 15 3 1 9 3 1 11 13 9 0 9 2
21 1 0 9 13 11 2 0 9 1 10 9 2 1 9 12 2 16 13 0 9 2
22 10 9 13 1 9 7 3 1 0 9 1 9 0 9 2 1 15 13 3 12 9 2
38 11 3 13 2 16 10 0 9 13 9 7 10 9 1 15 2 16 1 0 2 0 9 13 4 13 0 9 2 13 0 9 2 15 13 1 0 9 2
28 0 9 0 9 13 9 2 16 1 11 13 9 7 9 7 16 13 15 3 9 9 16 9 2 13 9 11 2
34 0 9 13 0 9 2 16 1 0 9 0 0 9 1 9 12 13 7 10 9 7 9 2 15 15 10 9 1 9 13 1 0 9 2
28 9 0 9 11 11 11 13 16 0 7 0 9 7 13 2 16 10 9 13 2 16 0 9 13 0 1 9 2
14 0 9 11 13 1 10 0 9 11 7 9 11 11 2
38 10 9 13 7 9 0 0 9 11 11 7 10 2 0 9 2 2 7 3 9 15 13 0 0 0 0 9 11 11 2 15 13 16 0 7 0 9 2
19 12 9 1 0 9 1 9 3 12 9 9 13 3 3 1 11 1 11 2
26 9 0 9 1 9 7 9 2 11 2 1 9 13 12 9 9 2 0 9 7 9 1 9 9 11 2
5 9 11 11 2 11
6 12 12 0 9 1 9
2 11 2
17 1 11 13 3 1 9 12 12 0 9 2 10 9 13 9 9 2
12 1 0 9 1 11 15 13 9 9 11 11 2
10 13 2 16 13 13 9 0 0 9 2
20 2 1 10 9 2 15 13 3 9 2 15 3 13 1 15 13 2 2 13 2
18 11 13 2 16 9 9 3 13 9 9 2 15 13 1 0 0 9 2
17 10 9 13 9 0 9 7 9 1 9 13 2 16 13 1 9 2
21 1 0 9 14 12 9 0 9 1 9 0 9 13 9 1 0 9 12 9 9 2
10 15 13 9 0 9 7 9 0 9 2
19 2 9 1 0 9 13 3 13 9 9 7 0 9 9 2 2 13 11 2
25 13 2 16 9 9 9 13 13 3 7 13 13 1 9 0 9 1 9 1 0 9 1 0 9 2
7 11 2 9 15 13 1 9
2 11 2
34 9 9 0 1 0 9 11 15 1 0 9 13 7 1 12 2 12 9 13 1 9 11 1 11 2 15 13 3 12 9 1 0 9 2
23 9 2 15 3 13 3 3 1 0 9 7 13 0 9 2 13 1 0 9 1 12 9 2
18 13 1 15 11 11 1 0 9 0 9 7 13 2 16 13 9 9 2
33 0 15 0 9 13 1 11 11 2 9 9 14 2 15 13 0 9 2 0 9 0 9 1 9 9 9 1 0 9 1 0 9 2
9 0 9 9 15 1 15 3 13 2
4 0 0 9 2
15 1 9 7 1 9 13 3 9 2 3 9 9 1 9 2
13 0 0 9 1 9 12 7 12 2 9 2 9 2
13 0 0 9 1 12 9 12 7 12 9 2 9 2
12 9 13 1 9 1 12 7 13 1 12 9 2
10 9 13 1 12 7 13 1 12 9 2
26 0 9 12 2 9 2 0 9 12 9 2 9 1 9 12 2 0 9 12 9 2 9 1 9 12 2
9 0 0 9 13 12 9 2 9 2
21 1 9 9 13 2 15 13 1 10 9 2 7 7 15 13 3 10 9 2 2 2
8 9 1 9 9 1 9 13 0
2 11 2
29 10 0 9 1 9 10 12 0 9 1 0 9 2 15 15 13 0 9 1 9 2 3 1 9 9 9 3 13 2
10 13 15 3 9 9 0 9 11 11 2
7 9 10 9 13 1 0 2
13 1 10 9 13 3 0 15 1 10 9 3 13 2
20 2 16 9 13 9 1 9 1 9 2 3 15 4 10 9 13 2 2 13 2
17 9 0 0 9 4 15 1 11 9 13 13 3 9 1 0 9 2
38 13 2 16 3 13 0 2 15 15 13 2 7 13 2 16 9 9 11 11 13 1 9 2 3 15 13 9 13 2 3 1 11 1 9 9 0 9 2
5 0 2 9 1 0
5 11 2 11 2 2
18 0 9 7 9 1 10 0 9 0 1 0 0 9 13 13 9 0 2
16 16 13 10 9 11 9 2 0 15 7 1 9 13 1 9 2
15 2 13 15 13 1 9 0 9 1 0 9 2 2 13 2
26 9 4 13 1 9 1 9 12 3 0 1 9 0 12 9 9 2 16 4 10 9 13 3 12 9 2
32 1 0 9 1 9 9 0 13 2 16 15 1 15 2 13 9 2 7 16 7 0 9 13 1 15 9 13 10 10 0 9 2
22 15 4 15 0 1 0 9 3 1 0 9 3 0 9 13 13 9 9 1 9 9 2
4 11 13 0 9
2 11 2
19 1 11 15 3 13 0 9 2 1 15 15 13 9 9 1 0 0 9 2
26 1 0 9 15 13 1 0 9 2 0 9 13 13 1 12 1 12 9 7 9 15 13 3 1 9 2
10 13 15 0 9 9 1 9 0 9 2
15 9 11 11 13 2 16 0 9 4 13 1 12 2 9 2
8 13 1 0 9 1 0 9 2
9 9 9 13 11 11 3 9 11 2
19 0 9 0 9 2 16 13 0 9 0 9 2 4 13 1 12 2 9 2
14 3 0 0 9 15 13 3 10 9 7 13 10 9 2
7 9 1 9 1 9 12 2
5 9 13 3 7 3
5 11 2 11 2 2
22 0 9 9 9 0 0 9 2 1 9 12 2 13 0 9 1 9 0 9 3 3 2
7 13 1 12 9 0 9 2
17 0 9 11 13 1 0 9 7 3 13 2 16 15 15 13 13 2
19 9 3 3 13 9 12 0 0 9 2 7 15 1 11 7 1 9 11 2
17 9 9 3 0 9 13 2 16 1 9 0 9 15 3 9 13 2
12 3 13 3 3 9 2 16 13 0 0 9 2
5 9 1 0 9 2
8 9 13 7 1 9 0 9 2
7 1 0 9 13 3 0 2
16 9 13 13 0 9 2 1 15 4 0 9 0 9 13 9 2
15 0 9 4 13 13 9 1 9 9 9 1 9 0 9 2
21 0 0 9 13 1 12 1 0 2 9 2 2 15 13 9 9 9 11 0 9 2
6 13 13 0 0 9 2
18 9 15 13 3 9 0 9 7 9 11 2 0 0 7 0 9 2 2
23 13 13 9 11 0 9 1 15 2 16 4 13 13 0 9 2 15 4 13 16 0 9 2
4 0 9 15 13
5 11 13 0 0 9
2 9 9
5 11 2 11 2 2
31 0 9 13 3 10 9 13 1 0 9 2 16 9 2 1 15 13 13 9 2 15 13 3 7 13 15 9 1 9 9 2
16 13 15 1 9 2 15 3 13 1 9 1 11 0 0 9 2
32 11 2 11 2 9 0 9 11 0 9 0 9 13 2 16 1 9 9 13 1 0 9 0 9 2 15 13 7 9 9 11 2
11 15 4 13 13 7 0 9 0 9 11 2
20 0 9 13 0 9 9 0 9 2 7 7 13 4 10 0 9 13 0 9 2
18 16 13 11 2 11 2 0 9 3 13 10 9 1 0 9 1 9 2
25 9 9 13 13 0 2 0 9 0 12 9 2 0 16 9 9 1 0 9 7 0 1 0 9 2
18 0 9 13 13 7 0 9 0 9 2 15 13 13 3 9 0 9 2
5 0 9 1 0 9
10 1 11 13 3 4 13 0 2 0 9
2 9 9
4 11 2 11 2
21 15 9 0 0 9 0 9 1 0 9 1 11 7 11 13 3 1 9 1 11 2
40 0 9 11 11 7 9 9 11 11 13 3 3 1 0 9 9 11 11 2 15 1 0 9 13 0 9 7 3 15 13 1 9 0 2 0 9 1 9 9 2
17 10 0 9 11 11 2 15 15 3 13 9 2 13 1 15 3 2
18 13 2 14 15 1 9 2 13 11 7 11 9 3 1 12 9 9 2
17 9 13 15 1 15 13 0 9 1 9 0 9 1 9 0 9 2
24 11 13 2 16 1 12 9 1 9 13 13 10 9 2 3 7 3 13 10 9 1 10 9 2
21 1 9 4 13 13 1 11 7 11 13 0 9 2 15 13 13 9 1 0 9 2
7 3 13 9 3 1 0 9
5 13 15 0 9 2
25 0 9 2 15 15 13 13 13 2 13 11 2 16 2 15 13 13 11 1 9 1 0 9 2 2
16 0 0 9 9 11 7 13 2 16 13 1 2 0 9 2 2
15 1 10 9 13 15 9 0 9 9 11 7 9 11 11 2
9 1 9 10 9 13 9 9 0 2
2 11 2
3 9 1 11
3 9 9 12
20 9 9 11 11 13 3 3 0 2 1 9 0 9 13 2 1 0 9 2 3
5 9 11 9 2 11
3 9 9 9
5 11 2 11 2 2
23 0 9 2 15 13 9 2 7 2 9 3 0 1 13 9 2 13 1 9 0 9 11 2
30 1 0 9 1 0 9 2 15 3 13 1 11 2 13 9 2 11 11 1 11 2 16 9 9 1 10 9 3 13 2
44 16 1 9 12 0 9 3 2 3 2 0 9 9 2 2 13 1 9 2 12 9 2 9 0 12 5 15 9 13 1 0 9 2 2 3 4 1 9 9 13 3 12 9 2
21 1 0 9 15 3 13 0 9 13 9 7 3 15 13 2 16 15 9 13 9 2
25 1 11 3 13 13 2 3 15 9 13 7 3 1 9 7 3 15 0 9 2 9 2 3 13 2
9 0 9 1 11 1 9 9 13 2
27 0 9 9 9 11 0 13 2 16 1 9 2 15 1 9 13 2 4 3 13 3 9 9 7 9 9 2
30 9 4 13 13 3 0 2 16 15 9 1 9 13 1 2 0 2 0 9 2 2 10 9 7 13 13 1 0 9 2
7 3 15 13 14 9 0 2
31 1 9 0 9 13 15 3 1 9 9 1 12 9 2 9 1 0 9 2 9 9 2 1 9 1 9 7 1 9 3 2
5 0 11 13 3 9
5 11 2 11 2 2
17 0 9 0 9 15 1 0 9 9 1 12 9 13 1 9 9 2
16 16 1 9 12 13 12 9 2 9 0 9 3 15 13 12 2
17 16 13 1 9 0 0 9 0 9 2 1 0 9 13 11 3 2
20 1 9 12 13 0 9 12 9 2 1 9 1 0 9 12 7 1 0 12 2
23 3 15 1 11 13 12 7 9 9 9 2 15 13 3 1 12 12 3 16 1 9 12 2
10 13 12 12 9 7 9 9 9 13 2
4 13 12 9 2
8 0 9 9 15 13 1 9 2
16 1 9 11 9 15 1 0 9 13 13 1 9 11 0 9 2
26 16 4 13 14 1 3 0 2 13 4 10 9 1 0 9 1 9 12 1 9 12 9 3 16 3 2
19 0 9 7 13 13 7 1 0 0 9 2 3 9 9 1 0 9 9 2
12 7 1 9 3 9 9 13 7 3 15 13 2
32 2 0 2 15 13 2 13 9 1 9 2 2 13 11 2 11 7 13 2 16 13 9 9 1 11 7 3 3 1 0 9 2
5 11 13 9 0 9
5 11 2 11 2 2
32 9 1 9 7 9 9 0 9 2 11 2 13 1 9 12 9 9 9 9 0 9 9 9 11 11 2 15 9 13 0 9 2
10 11 1 15 3 13 9 11 11 9 2
26 9 13 13 11 11 2 15 13 1 9 12 1 9 1 0 9 16 9 9 0 9 1 0 9 9 2
13 1 9 12 11 11 2 11 13 7 13 1 9 2
19 9 9 2 11 13 9 12 2 9 1 9 0 9 9 1 11 1 11 2
10 0 9 9 11 11 11 13 1 9 2
16 1 9 12 15 13 9 2 11 13 1 9 7 3 1 11 2
24 10 9 11 15 13 1 11 0 9 1 0 9 1 9 2 15 13 13 1 9 1 9 9 2
32 11 13 3 1 9 9 9 11 2 1 15 15 3 13 2 1 9 10 9 7 3 13 7 9 1 11 7 3 14 1 11 2
28 11 13 3 2 16 13 9 9 2 10 9 7 9 9 2 7 16 0 11 15 13 1 9 1 9 9 11 2
13 0 0 9 15 3 13 10 9 13 9 0 9 2
25 9 2 16 11 11 2 2 13 1 12 9 1 11 1 9 9 2 15 15 15 13 1 9 12 2
15 11 15 13 1 9 7 3 13 9 2 16 10 9 13 2
17 1 9 10 9 15 1 11 13 1 10 0 9 14 1 9 12 2
29 10 9 1 11 2 11 13 7 9 9 11 11 2 7 13 1 9 2 16 13 1 9 9 2 7 1 0 9 2
35 11 13 9 3 1 10 0 9 2 3 13 11 1 0 9 13 9 0 9 2 7 7 15 13 1 9 1 9 2 16 4 13 1 9 2
2 9 9
5 11 2 11 2 2
27 1 0 9 10 0 9 1 9 0 9 1 11 13 3 1 0 9 9 9 9 11 2 11 2 11 2 2
35 1 12 2 9 9 9 11 2 11 1 9 1 0 9 13 2 16 1 9 2 3 9 13 9 1 9 2 13 1 9 15 1 0 9 2
37 3 0 9 2 15 13 0 2 9 2 11 7 9 9 0 9 1 9 9 9 1 9 11 2 13 0 0 9 1 9 9 11 11 3 1 0 2
38 1 9 3 7 9 0 9 1 0 9 2 11 2 13 2 16 9 9 9 2 16 9 9 9 7 9 1 9 0 9 2 4 1 9 11 3 13 2
23 1 9 11 15 1 9 3 13 0 9 7 0 0 9 11 0 2 9 2 13 3 0 2
50 1 0 9 13 1 11 7 10 9 1 9 2 16 9 0 9 1 0 9 2 11 2 7 9 9 11 3 13 2 16 4 10 9 13 9 0 9 9 12 13 0 9 2 15 13 9 1 9 9 2
28 9 11 13 9 1 15 2 16 9 13 13 2 0 1 9 2 2 7 9 2 16 4 13 0 13 0 9 2
12 1 0 9 13 13 3 0 9 9 2 9 2
7 9 13 1 9 2 9 9
2 11 2
20 9 0 9 1 12 1 12 9 9 13 9 7 3 2 13 10 0 9 2 2
10 3 9 0 9 1 10 9 15 13 2
15 13 15 1 9 2 15 13 9 9 1 9 1 9 11 2
17 1 0 9 12 12 0 9 1 12 1 12 9 13 9 0 9 2
9 9 1 15 3 13 3 16 9 2
10 9 1 9 9 7 1 0 9 13 2
50 9 1 9 7 9 9 11 13 0 2 15 13 1 9 9 9 0 9 7 10 9 1 0 9 2 16 4 15 13 1 0 9 1 9 2 11 11 2 0 9 9 2 12 2 11 2 12 12 11 12
20 0 9 0 9 15 9 4 13 1 9 9 0 9 13 1 9 12 2 9 2
4 9 13 0 2
16 1 9 1 0 9 0 9 13 1 12 2 9 9 12 9 2
19 9 4 13 13 1 9 12 9 7 0 0 9 4 13 13 13 1 9 2
6 1 11 13 9 12 9
7 11 2 11 2 11 2 2
16 9 13 1 9 1 0 9 1 9 1 0 9 1 12 9 2
21 16 15 10 9 3 14 13 13 0 9 2 9 0 9 15 3 13 14 1 11 2
13 1 9 9 13 13 2 16 15 9 4 3 13 2
25 9 1 0 9 13 13 7 9 9 9 2 7 9 0 9 4 13 3 0 9 9 1 0 9 2
20 1 11 1 1 15 15 15 0 7 0 9 13 3 1 9 2 3 1 9 2
18 1 9 1 11 15 1 9 13 14 12 9 7 1 9 1 12 9 2
7 9 1 0 9 7 13 2
7 9 3 3 13 9 9 2
20 16 11 13 0 9 0 0 9 11 11 2 11 2 15 13 13 1 0 9 2
19 15 2 15 13 9 1 9 7 0 9 2 3 13 9 1 9 10 9 2
12 13 15 3 15 13 2 3 1 15 13 9 2
9 2 1 10 0 9 1 9 13 2
12 13 15 3 1 9 2 2 13 11 2 11 2
2 11 2
30 9 0 9 11 11 2 9 12 11 2 13 9 10 9 2 15 15 1 12 2 1 12 2 9 13 1 0 9 9 2
28 9 1 0 9 2 9 1 9 0 9 7 9 2 0 0 9 7 0 0 9 11 2 12 1 15 13 3 2
13 12 1 0 9 13 1 0 0 9 11 3 13 2
9 13 1 9 11 2 9 7 11 2
14 13 15 4 3 3 1 12 2 12 7 9 13 0 2
5 13 9 1 9 9
7 11 2 11 2 11 2 2
24 1 9 0 9 1 11 13 1 9 3 0 11 2 11 2 10 1 9 0 9 2 9 9 2
22 9 2 15 13 3 13 1 0 9 2 13 1 12 0 9 3 0 9 9 12 9 2
10 1 9 13 0 9 13 7 13 9 2
6 9 9 13 3 0 2
39 0 9 13 9 0 9 1 11 2 16 4 0 9 0 9 11 1 11 13 9 11 2 7 13 9 1 0 9 7 1 9 7 9 0 9 1 10 9 2
15 16 4 11 13 1 9 9 2 13 15 9 1 11 13 2
8 11 13 2 0 9 2 0 9
7 11 2 11 2 11 2 2
28 1 9 9 0 9 2 16 4 13 9 9 0 9 0 9 9 2 13 10 9 9 11 11 3 12 9 13 2
27 1 10 9 4 13 0 9 9 1 0 9 13 9 11 11 7 13 0 2 16 15 1 0 9 13 15 2
27 9 0 9 9 11 0 2 11 11 2 7 9 9 11 11 2 11 2 13 2 16 0 9 13 13 9 2
19 1 10 9 11 2 11 2 11 7 11 4 9 12 0 9 13 13 9 2
16 9 0 9 15 1 9 0 9 13 9 0 9 11 11 0 2
4 2 11 2 2
8 1 10 9 13 1 12 9 2
15 1 11 13 14 10 9 9 2 7 9 0 9 7 9 2
8 1 0 9 13 1 9 0 9
5 11 2 11 2 2
14 0 9 13 0 9 1 9 1 0 9 1 0 9 2
18 1 9 0 9 0 9 0 9 1 11 15 3 13 10 9 11 11 2
28 3 1 9 13 9 0 9 0 0 2 9 15 13 1 15 0 9 2 3 15 9 13 3 1 10 0 9 2
24 3 3 1 0 7 0 11 13 0 9 3 3 7 1 0 9 2 16 1 11 2 13 11 2
12 11 15 1 15 3 13 1 0 9 1 9 2
28 11 2 15 13 3 10 9 13 1 9 3 1 11 2 15 7 3 13 13 1 0 9 0 11 1 0 9 2
14 2 7 11 13 3 13 1 0 9 2 2 13 9 2
12 9 15 1 9 1 9 7 1 0 9 13 2
19 13 7 9 1 12 0 9 1 9 7 1 0 9 9 1 0 0 9 2
20 11 3 13 1 9 1 9 9 7 13 2 16 4 1 10 9 4 13 9 2
33 9 2 15 13 1 9 0 0 12 9 2 13 1 11 0 9 2 16 15 13 9 1 15 0 9 1 11 7 11 1 13 11 2
17 3 3 13 9 1 15 2 16 4 1 9 4 13 0 9 11 2
33 9 9 11 2 15 13 9 1 11 9 2 13 3 11 2 16 2 9 13 3 0 2 7 16 15 1 9 13 9 1 0 9 2
10 9 14 13 1 0 9 9 9 11 2
17 9 0 0 9 0 1 9 11 3 13 0 9 0 0 0 9 2
9 13 15 0 9 1 0 9 11 2
24 12 9 13 0 11 7 13 15 9 1 9 0 9 2 16 15 3 13 1 2 0 9 2 2
6 13 15 3 0 9 2
21 0 9 2 15 4 13 1 0 9 1 9 2 4 13 13 1 15 3 12 9 2
19 13 15 3 1 0 9 9 9 11 1 15 2 16 9 3 0 9 13 2
6 0 9 1 9 7 9
2 9 9
5 11 2 11 2 2
40 9 13 15 13 9 2 7 2 9 7 9 2 13 12 1 9 0 9 1 9 0 0 0 9 2 9 2 2 10 9 9 0 9 13 7 13 1 9 9 2
16 9 4 13 1 9 11 13 0 9 9 1 9 0 9 11 2
10 0 9 3 13 0 7 0 9 9 2
27 1 9 10 9 4 15 13 9 13 9 2 10 9 4 13 14 0 9 2 7 13 4 13 1 0 9 2
24 10 9 13 9 1 9 1 9 2 0 9 9 1 9 0 0 9 7 1 9 1 13 9 2
13 9 0 9 13 9 1 0 9 2 9 7 9 2
17 0 9 13 3 13 1 9 9 9 7 9 9 1 3 0 9 2
42 1 9 9 13 9 9 9 1 9 12 9 1 0 2 1 9 9 9 7 0 9 2 2 0 9 7 10 9 3 13 13 15 0 9 2 7 1 9 9 9 2 2
33 1 9 9 1 9 15 13 0 9 10 0 9 7 9 2 15 13 9 1 9 10 9 7 15 13 0 9 2 0 1 10 9 2
16 3 4 1 9 13 9 2 1 15 13 10 0 9 9 9 2
28 13 1 9 12 2 7 12 2 9 2 0 9 2 9 2 9 2 9 2 0 9 2 9 2 9 9 3 2
27 1 9 9 13 9 0 9 13 0 9 0 0 9 7 9 2 1 0 9 13 3 13 7 0 0 9 2
15 3 15 13 7 1 9 9 2 0 9 2 9 7 9 2
29 0 0 9 4 13 13 0 9 1 0 9 2 1 0 9 4 9 9 13 4 13 9 0 7 9 9 0 9 2
5 0 2 9 1 0
5 11 2 11 2 2
2 9 0
2 11 11
14 9 0 9 11 13 2 16 0 9 0 9 13 9 2
11 0 0 0 9 13 1 9 9 7 9 2
7 13 15 13 14 0 9 2
10 13 13 0 9 7 13 1 0 9 2
5 4 13 0 9 2
13 10 9 13 9 1 9 9 12 1 9 0 9 2
20 15 3 13 2 16 4 1 0 9 1 9 12 13 13 0 9 0 9 0 2
24 9 13 7 1 0 9 10 10 9 1 10 10 9 2 0 0 9 1 9 2 15 13 15 2
20 1 9 9 12 13 9 1 0 13 1 9 2 16 4 13 9 1 13 9 2
32 9 10 9 3 7 13 2 13 15 7 1 9 3 0 9 7 0 9 2 1 15 15 9 0 0 9 10 0 9 13 3 2
21 9 1 9 13 9 1 9 9 16 0 2 10 9 15 3 13 1 9 0 9 2
10 9 13 1 0 9 13 9 10 9 2
6 3 3 13 13 0 2
16 9 13 1 10 9 9 9 0 9 1 9 0 0 0 9 2
5 11 13 14 13 2
15 9 11 13 3 3 9 2 16 9 1 9 13 3 3 2
11 0 9 15 13 3 0 9 0 9 9 2
16 10 9 13 2 16 9 15 1 9 0 9 0 9 13 3 2
47 9 0 0 9 11 11 3 13 2 16 4 13 1 9 1 9 7 9 2 7 13 2 16 0 2 9 2 2 16 13 9 9 7 9 1 10 9 2 13 13 3 0 9 7 3 9 2
12 1 0 9 13 9 7 9 13 1 0 9 2
19 13 10 9 0 9 13 3 0 2 16 7 0 9 4 13 13 0 9 2
9 1 0 9 13 9 3 0 9 2
12 1 9 0 9 13 0 13 9 7 0 9 2
5 15 13 9 0 2
18 1 9 7 9 9 3 4 13 9 7 9 9 1 0 9 0 9 2
9 13 3 2 9 0 9 13 13 2
16 9 14 13 7 3 13 14 1 15 13 3 9 0 0 9 2
19 3 2 9 13 0 9 9 7 3 3 14 9 0 0 9 1 10 9 2
5 13 15 4 9 2
21 13 2 14 15 9 7 9 1 10 0 9 2 13 15 3 0 9 10 0 9 2
7 9 1 0 9 13 16 9
5 11 2 11 2 2
19 9 0 9 7 9 9 7 9 13 3 9 3 13 1 0 15 0 9 2
25 10 9 13 14 9 11 1 9 2 7 7 9 10 0 9 2 15 13 9 13 1 0 9 9 2
28 9 0 9 3 0 15 9 9 1 0 9 13 0 9 1 9 2 15 15 13 9 9 1 0 9 7 9 2
28 9 2 16 4 9 13 1 0 9 9 0 9 2 11 11 13 2 16 15 13 2 16 11 4 9 9 13 2
22 11 13 1 0 0 9 3 13 9 12 9 7 0 4 13 9 0 12 9 0 9 2
15 9 11 7 13 2 16 1 10 9 13 0 13 0 9 2
24 10 9 13 1 0 9 2 0 9 9 7 9 2 11 2 11 7 13 7 0 9 1 11 2
27 1 0 9 15 11 13 3 2 7 1 11 15 13 0 2 1 3 0 9 3 13 10 9 12 9 9 2
8 15 9 11 13 13 0 9 2
6 0 9 13 1 0 9
2 11 2
23 9 2 16 4 0 9 13 9 1 9 0 9 1 9 0 9 2 4 13 1 12 9 2
16 13 15 3 9 11 11 2 11 2 2 15 13 9 0 9 2
39 9 1 0 9 9 11 11 0 2 11 2 13 1 9 9 1 0 9 9 2 1 15 15 9 0 9 13 3 1 9 0 9 1 9 9 12 7 12 2
29 1 0 9 13 0 9 14 1 10 9 9 2 7 7 1 9 0 9 7 9 7 1 0 9 2 15 11 13 2
28 9 2 0 0 9 2 13 4 13 0 9 14 1 9 2 3 9 9 13 1 9 2 12 2 9 12 2 2
9 0 9 13 4 3 13 12 9 2
22 11 13 2 16 10 9 4 13 1 1 15 2 16 1 0 9 15 13 12 9 9 2
10 1 9 0 9 1 9 3 3 15 13
5 11 2 11 2 2
10 0 9 1 9 3 3 3 15 13 2
23 14 1 9 12 15 13 9 1 9 12 9 0 9 2 15 3 3 1 10 9 3 13 2
22 3 1 9 0 0 9 7 3 9 0 13 0 9 7 9 7 7 9 3 0 9 2
24 0 9 1 9 4 15 13 13 3 9 9 7 10 9 1 0 9 2 9 9 7 10 9 2
13 13 3 0 13 9 1 9 2 0 9 2 9 2
22 0 9 1 0 9 7 9 13 1 15 2 16 4 0 9 1 9 13 0 3 3 2
9 3 7 10 9 13 9 10 9 2
16 3 3 13 9 9 7 0 9 2 4 15 13 9 11 11 2
30 2 0 9 9 7 0 9 13 9 9 7 15 15 13 1 15 2 16 9 9 7 0 9 4 13 13 9 10 9 2
18 9 2 15 4 13 10 0 9 13 2 13 1 10 9 3 12 9 2
12 9 13 1 9 9 2 9 2 1 9 2 2
27 9 11 13 2 16 13 9 9 9 11 11 7 9 9 11 11 1 9 2 1 15 15 13 1 0 9 2
12 9 1 0 9 13 9 14 1 12 9 9 9
7 11 2 11 2 11 2 2
31 13 9 0 0 9 2 9 2 7 9 16 0 9 1 0 9 13 9 0 9 9 1 9 7 9 10 0 9 7 9 2
9 9 9 13 1 10 9 9 9 2
11 1 10 9 13 0 9 1 9 9 0 2
22 1 3 0 9 9 1 9 13 1 9 14 3 0 9 9 9 1 9 12 9 9 2
6 9 4 15 13 13 2
34 0 9 4 13 1 9 9 13 9 9 0 9 1 15 0 7 0 9 2 15 13 0 9 1 9 7 3 15 3 13 16 0 9 2
14 3 1 10 9 1 9 15 9 13 13 3 0 9 2
9 9 9 1 10 9 13 3 0 2
38 1 0 9 13 9 0 9 1 0 9 7 9 10 9 7 9 2 3 15 2 15 10 9 13 1 9 7 13 15 16 0 9 2 3 7 10 9 2
32 16 7 10 9 13 0 0 9 0 16 0 9 2 13 9 0 9 0 9 2 15 3 13 13 9 9 1 10 9 0 9 2
24 0 9 4 13 13 9 7 9 0 9 7 9 9 1 10 9 2 12 7 12 9 9 2 2
11 10 9 4 15 13 13 9 1 12 9 2
5 1 0 0 9 3
2 11 2
24 9 0 0 9 4 13 13 11 11 2 15 4 3 13 9 0 0 9 16 9 0 0 9 2
17 9 11 3 13 9 11 2 13 15 1 15 13 3 0 0 9 2
11 11 13 1 11 9 9 1 9 1 9 2
6 13 9 10 0 9 2
16 1 9 2 15 15 3 13 1 0 9 2 13 1 9 12 2
18 9 9 0 0 9 2 15 13 1 11 2 13 1 12 2 9 13 2
8 9 1 11 11 2 9 9 11
18 13 9 2 16 1 0 9 1 9 9 13 9 0 9 1 9 0 2
14 3 13 1 15 2 16 3 3 4 13 0 9 13 2
11 13 0 9 1 0 13 3 9 3 0 2
12 15 3 3 3 13 9 7 13 1 9 0 2
28 16 13 1 0 0 9 2 13 13 9 0 0 9 2 0 0 9 1 9 2 15 4 13 13 0 9 9 2
10 7 1 15 14 15 3 0 9 13 2
8 0 9 0 9 13 0 9 2
24 9 1 9 15 13 2 16 15 3 15 13 2 7 15 4 13 2 9 15 13 13 7 13 2
12 7 13 15 2 16 3 4 3 13 9 13 2
5 3 4 15 13 2
34 14 4 13 2 16 13 0 13 1 15 2 16 15 2 15 15 4 13 1 0 9 2 13 0 9 1 15 2 15 15 3 13 9 2
9 3 1 0 9 0 9 9 13 2
3 2 11 2
8 11 2 11 1 9 1 0 9
5 11 2 11 2 2
11 9 11 11 13 3 1 9 9 1 9 2
28 1 3 0 9 9 11 11 7 1 9 9 11 11 13 1 9 9 1 0 9 7 10 9 1 0 0 9 2
12 9 1 0 9 1 0 9 13 13 0 9 2
9 11 13 1 9 2 9 1 9 13
4 11 2 11 2
16 1 9 0 2 0 0 9 4 1 9 1 9 13 0 9 2
43 0 9 9 7 9 0 2 0 0 9 13 2 16 1 9 0 9 9 2 15 13 0 11 7 15 13 0 9 1 0 9 1 0 9 1 11 2 3 13 9 0 9 2
15 0 11 7 10 9 13 7 3 13 1 0 9 0 9 2
20 0 9 1 9 1 9 4 15 13 13 0 9 1 3 12 9 0 0 9 2
22 9 0 9 4 3 3 13 7 13 9 0 9 14 1 11 2 7 7 1 0 11 2
21 9 13 3 0 9 1 11 2 15 13 1 10 9 13 0 9 1 11 7 11 2
24 0 9 0 9 11 1 0 11 11 11 3 13 9 1 0 0 2 0 9 1 11 7 11 2
10 13 15 3 1 11 9 9 11 11 2
49 2 0 9 9 13 9 1 0 9 11 7 11 2 2 13 9 2 0 9 2 2 1 15 15 11 3 1 0 9 13 1 0 0 2 0 9 11 11 7 1 0 11 1 9 0 11 11 11 2
22 11 13 9 9 11 13 9 1 11 2 13 3 11 11 1 9 1 0 9 11 11 2
27 11 7 9 11 13 2 16 4 3 13 9 1 9 1 11 2 3 15 13 0 11 13 7 1 0 9 2
24 2 0 0 9 2 1 10 9 13 2 13 1 11 2 2 13 9 0 9 1 9 1 11 2
20 1 9 11 1 0 0 9 0 2 0 9 2 15 3 13 1 12 0 9 2
4 11 13 0 9
4 11 2 11 2
34 0 9 13 3 1 0 9 3 9 2 1 15 9 13 13 0 9 2 15 13 13 0 9 9 7 15 13 13 14 1 9 0 9 2
18 9 9 13 3 9 1 0 9 1 11 2 15 13 1 0 0 9 2
24 9 2 16 1 11 13 9 13 0 9 1 3 0 1 0 2 13 3 1 11 9 9 11 2
28 13 1 10 9 9 9 9 11 11 2 15 13 1 9 0 9 2 16 11 3 13 2 3 13 9 10 9 2
16 11 11 1 0 9 13 1 11 7 13 15 3 1 11 11 2
27 9 0 9 13 1 9 1 9 1 0 11 2 16 4 15 13 13 0 9 2 15 3 13 3 12 9 2
11 1 9 7 9 4 13 3 12 9 9 2
4 9 11 2 9
4 11 13 9 9
2 11 2
15 0 9 9 11 11 13 10 0 9 1 0 9 9 9 2
43 9 1 9 13 15 11 2 16 1 9 1 9 0 13 2 16 1 9 9 11 1 0 9 2 9 2 0 9 11 2 7 1 15 0 9 9 4 13 3 0 0 9 2
32 1 0 9 9 0 11 9 10 0 9 13 2 2 16 4 9 3 3 13 4 13 2 13 15 9 9 2 7 3 9 2 2
22 1 0 9 13 0 9 9 14 1 9 15 1 2 0 0 9 2 7 15 9 13 2
9 11 15 13 1 2 9 2 1 11
2 11 2
24 11 13 13 13 0 0 9 3 0 9 11 2 16 4 10 9 13 1 11 12 0 0 9 2
6 13 15 9 0 9 2
14 1 0 9 13 0 9 9 11 2 15 13 1 11 2
10 9 11 7 14 9 1 0 9 13 2
24 13 1 11 12 9 9 2 9 11 2 0 7 0 9 2 12 9 7 12 9 7 9 9 2
5 9 1 11 13 9
4 11 2 11 2
12 9 1 0 0 9 3 3 13 0 9 11 2
7 1 9 13 1 9 9 2
12 9 9 13 1 9 1 11 2 11 7 11 2
9 9 15 13 1 0 9 1 9 2
30 9 0 9 11 13 2 16 9 1 0 11 2 1 15 15 13 1 12 9 2 13 0 9 16 9 2 9 7 9 2
4 0 9 13 9
2 11 2
23 14 12 0 0 9 2 10 0 9 1 0 9 0 9 13 0 9 2 4 13 0 9 2
31 1 0 13 0 0 9 11 2 11 7 11 2 11 2 0 9 11 2 11 2 11 7 0 0 9 0 9 11 2 11 2
23 9 3 13 1 9 9 2 16 4 4 9 13 7 0 0 9 9 7 9 11 2 11 2
6 9 11 1 11 2 11
2 11 2
26 9 0 9 0 9 11 11 2 11 2 1 9 0 0 9 13 3 1 11 0 0 9 2 11 2 2
25 10 9 13 2 16 0 9 11 2 15 13 4 11 13 2 13 9 10 9 1 9 1 0 11 2
17 11 2 15 1 11 13 2 15 13 1 9 0 9 1 0 9 2
24 13 3 9 0 9 7 13 1 15 9 2 15 13 12 9 1 0 9 0 9 9 1 11 2
6 9 13 15 3 3 9
2 11 2
27 0 9 0 9 1 0 9 1 9 13 12 9 9 7 9 7 0 9 3 15 1 15 13 3 0 9 2
12 13 3 1 3 0 9 2 9 0 9 2 2
33 13 15 9 0 9 9 11 11 1 0 9 9 0 1 11 0 9 9 7 9 9 2 15 15 13 7 9 1 10 9 0 9 2
18 11 13 2 16 9 2 9 9 2 9 9 1 0 9 13 0 9 2
19 9 13 3 0 9 1 9 7 1 0 9 2 7 9 0 9 0 9 2
29 9 3 13 2 16 1 0 9 15 13 0 9 3 0 0 9 2 7 15 1 9 2 3 0 9 0 9 2 2
4 0 9 1 9
6 11 2 11 2 11 2
23 0 9 3 13 9 7 13 2 16 0 9 13 13 12 9 0 0 9 7 9 1 9 2
36 11 11 2 15 13 0 9 1 9 0 0 9 2 11 2 2 13 1 11 2 16 0 9 1 11 7 0 9 4 13 1 9 3 0 9 2
38 11 2 1 15 13 13 3 9 9 11 2 13 2 16 0 9 2 15 4 13 9 9 1 0 9 9 11 11 7 1 15 13 9 11 2 13 0 2
14 1 0 9 11 3 13 0 9 1 0 9 7 9 2
28 0 9 0 9 3 13 2 16 1 9 11 1 9 9 4 1 9 13 12 9 7 12 0 9 0 0 9 2
25 1 0 9 11 13 15 3 1 12 9 9 1 11 2 16 3 4 9 10 9 13 1 0 9 2
14 9 1 9 1 11 15 1 0 9 13 3 12 0 2
32 0 9 9 11 11 1 9 13 9 1 0 9 11 2 15 4 13 0 9 1 11 2 7 13 0 9 2 7 1 9 9 2
14 13 15 1 9 2 15 3 13 9 0 0 11 11 2
12 0 9 13 1 0 9 1 12 9 1 11 2
7 3 13 1 0 0 9 2
18 9 11 1 0 9 1 11 13 2 16 13 1 9 1 9 0 9 2
21 0 9 11 2 11 13 1 9 9 1 11 7 11 2 15 13 1 10 9 0 2
13 13 15 1 11 1 9 0 9 0 9 1 9 2
18 0 9 13 1 9 1 9 9 0 9 9 1 9 1 9 0 9 2
13 10 9 13 0 10 9 1 10 9 1 12 9 2
29 9 11 9 11 3 9 0 9 11 11 13 2 16 4 4 13 9 1 9 1 9 0 1 9 9 7 0 9 2
22 9 9 11 11 3 13 2 16 0 0 9 11 4 13 0 9 1 9 1 0 9 2
23 9 0 0 9 4 1 9 13 1 0 11 1 9 1 11 2 16 0 9 13 10 9 2
11 13 15 9 11 1 9 1 0 0 9 2
19 1 9 0 9 13 3 1 9 12 9 7 12 4 13 1 9 10 9 2
9 13 15 3 0 9 9 1 9 2
27 1 0 9 13 1 9 0 12 9 2 1 15 15 13 1 9 13 2 16 15 9 13 1 9 0 9 2
17 11 3 13 12 0 9 2 15 3 1 9 13 9 1 9 11 2
16 13 15 0 0 9 1 15 2 16 9 15 13 1 0 9 2
16 0 0 0 9 9 1 9 0 11 13 9 3 14 9 9 2
7 13 15 3 0 9 11 2
13 9 9 11 1 11 7 13 10 9 13 7 13 2
32 9 9 9 2 15 15 13 12 2 7 12 2 9 13 9 0 9 12 2 4 1 0 9 13 1 12 2 7 12 2 9 2
11 13 15 3 0 9 11 2 11 2 11 2
27 3 12 9 13 7 3 16 12 13 13 1 0 9 11 7 0 9 2 15 1 9 1 9 13 0 9 2
15 13 15 9 11 1 9 1 0 9 0 9 7 0 9 2
5 1 11 13 9 9
2 11 2
20 1 12 9 0 9 13 1 0 9 1 9 13 9 1 0 12 9 0 9 2
32 9 0 0 0 9 13 2 16 0 0 9 11 11 13 1 12 9 9 1 0 9 11 1 11 2 15 3 13 12 9 9 2
26 1 0 9 13 3 0 9 9 11 11 11 1 12 9 7 1 0 0 9 0 9 1 12 9 9 2
17 0 9 13 0 9 1 0 11 2 15 15 3 13 0 9 9 2
31 1 9 12 12 0 9 13 1 0 11 1 0 9 1 9 1 0 9 3 12 9 9 2 16 0 0 9 14 12 9 2
15 1 9 4 15 13 1 0 9 13 0 9 0 1 9 2
22 10 9 13 13 0 0 9 2 9 9 9 2 15 15 13 9 0 0 9 11 11 2
13 1 9 9 13 4 13 12 9 7 9 0 9 2
7 15 12 13 1 9 9 2
17 3 0 9 15 13 9 3 3 2 16 15 3 13 9 11 11 2
13 15 15 13 1 11 12 2 9 2 13 9 11 2
25 1 11 15 3 13 0 9 9 11 11 1 0 9 11 1 11 2 16 4 3 13 9 0 9 2
26 9 0 0 9 9 11 11 11 3 13 2 16 9 11 1 9 13 13 0 1 15 7 13 13 9 2
38 1 9 1 9 13 2 16 0 9 13 11 0 9 2 15 13 1 15 1 2 0 9 0 2 16 13 9 2 16 13 9 2 16 4 15 13 2 2
4 11 13 15 15
2 11 11
19 15 2 15 15 1 9 13 2 15 13 13 14 1 15 2 15 13 9 2
13 10 9 13 0 9 11 11 0 9 1 0 11 2
30 9 2 15 13 1 0 12 9 2 3 1 0 9 13 9 11 11 2 13 0 9 7 13 1 0 1 0 12 9 2
21 0 9 0 9 2 15 3 1 0 11 7 11 13 9 2 3 13 0 9 9 2
24 1 0 2 0 9 1 0 9 7 0 0 0 9 2 11 2 3 13 1 12 12 12 9 2
35 14 1 0 9 13 1 0 11 12 9 2 15 9 0 9 11 1 9 2 11 2 13 1 2 0 7 0 9 2 2 15 3 11 13 2
20 0 9 13 0 7 13 1 15 3 15 2 0 9 7 9 13 7 9 13 2
28 0 9 10 9 1 12 2 9 13 9 9 0 9 11 1 11 2 11 2 1 0 9 2 12 9 2 2 2
19 1 9 11 2 1 9 7 9 9 15 3 13 0 9 7 9 3 0 2
20 0 9 13 1 9 9 0 9 2 9 2 9 7 2 14 2 9 2 2 2
30 3 0 2 0 9 0 2 0 2 11 1 0 0 11 7 1 11 1 9 0 9 13 1 3 0 9 9 7 9 2
34 1 11 9 2 9 0 9 0 0 11 2 0 0 9 3 13 12 2 9 1 9 2 3 4 13 2 9 2 9 1 9 9 11 2
9 1 9 3 13 15 1 0 9 2
33 0 0 9 2 13 15 3 11 2 2 0 0 2 9 2 2 13 13 1 0 9 1 2 9 9 2 7 13 9 1 0 9 2
15 12 9 3 13 9 1 9 9 11 7 13 1 15 13 2
42 9 15 13 7 13 15 0 9 2 0 1 9 2 3 11 2 11 7 9 0 0 9 13 1 11 10 9 2 4 2 14 9 13 15 15 2 15 0 15 3 13 2
16 9 15 3 2 16 3 15 2 13 1 9 7 0 9 9 2
23 1 9 9 13 0 9 11 7 9 0 0 9 2 1 12 0 9 13 9 11 11 12 2
31 9 9 13 1 9 1 9 9 2 15 3 13 9 1 10 9 2 16 3 1 11 15 13 2 9 2 0 9 0 9 2
30 0 9 11 13 13 2 16 9 2 15 13 9 11 13 2 3 13 9 9 9 2 7 13 13 9 0 9 2 2 2
24 15 9 13 3 0 2 16 10 9 13 3 13 13 1 11 0 9 9 1 9 10 0 9 2
11 1 12 9 0 9 1 11 3 13 0 2
8 11 4 13 15 15 2 2 2
4 9 9 1 11
10 0 9 7 9 13 9 1 12 9 9
2 9 9
7 0 9 11 1 11 11 11
15 13 2 14 15 15 1 9 2 3 15 13 3 10 9 2
21 15 13 7 9 9 1 9 11 11 2 15 0 9 13 1 0 9 12 9 9 2
15 0 12 10 9 13 0 9 2 0 7 0 0 0 9 2
9 7 3 10 9 15 13 1 9 2
20 13 0 0 7 3 0 9 2 16 4 9 13 1 9 7 9 0 0 9 2
18 9 2 15 1 0 9 13 9 2 13 3 0 2 16 13 14 3 2
6 7 2 15 13 9 2
23 15 12 9 9 13 9 7 9 11 11 7 10 9 11 16 9 9 3 1 12 0 9 2
9 0 9 13 9 1 9 12 9 2
19 7 16 0 9 13 9 2 0 0 0 9 3 13 7 13 3 0 9 2
4 15 13 9 2
21 3 3 15 13 0 0 9 2 0 9 13 3 9 9 0 0 0 9 1 11 2
27 1 9 10 9 4 3 12 1 0 9 13 13 0 2 16 0 9 13 9 0 9 2 15 13 0 9 2
21 1 15 2 16 15 13 9 2 13 13 2 16 7 12 9 9 0 9 13 9 2
17 9 2 7 1 0 9 0 9 2 13 0 9 7 9 9 11 2
19 15 13 0 9 9 2 15 13 16 9 1 0 9 2 7 9 9 13 2
22 1 13 9 13 12 9 9 2 16 0 9 15 13 1 12 9 7 9 13 12 9 2
27 9 9 2 0 10 9 9 1 9 0 9 1 11 2 13 11 16 12 0 9 2 1 9 3 12 2 2
20 1 9 0 9 1 10 9 2 15 15 13 12 9 9 2 13 9 12 9 2
6 1 9 2 0 9 2
11 1 9 15 1 0 9 13 9 12 9 2
14 1 0 9 13 11 12 9 16 9 1 9 0 9 2
8 1 9 15 13 3 12 9 2
16 10 15 15 13 1 9 0 9 9 2 15 0 9 13 13 2
5 0 9 7 0 9
18 11 11 3 9 13 2 16 9 13 7 9 0 9 7 9 0 9 2
4 15 3 13 2
15 9 7 13 2 3 9 7 9 13 2 3 13 2 13 2
15 0 9 13 9 3 0 9 2 16 0 9 15 3 13 2
21 9 11 2 0 11 13 7 3 0 2 16 7 9 9 13 9 13 16 3 0 2
18 7 3 10 9 2 0 9 2 9 0 9 2 13 2 7 3 3 2
26 1 15 13 7 0 13 2 16 10 9 3 0 9 16 0 11 13 2 7 16 9 0 9 4 13 2
19 13 15 2 16 11 13 3 0 9 2 16 0 9 13 3 3 16 3 2
14 3 13 9 9 0 9 2 1 15 0 9 13 2 2
12 13 13 3 0 9 10 9 7 0 9 3 2
6 15 3 9 3 13 2
25 3 3 13 9 2 16 0 9 9 0 9 3 9 10 9 13 9 0 9 7 13 9 1 9 2
7 11 11 7 13 3 9 2
31 13 9 2 15 13 0 9 0 9 2 9 1 0 9 2 0 0 0 9 2 0 9 2 7 7 9 9 1 3 0 2
16 13 0 0 9 2 13 9 2 13 9 3 0 9 2 2 2
5 0 13 9 7 9
25 3 11 13 1 9 13 9 2 13 9 2 16 9 1 0 9 1 9 13 1 0 9 1 11 2
7 3 3 9 1 10 9 2
27 16 2 16 15 9 9 13 2 16 4 13 2 1 9 2 2 13 13 9 1 9 12 7 12 9 9 2
20 15 2 13 2 1 10 0 9 3 3 2 16 1 15 0 9 13 13 9 2
10 13 3 3 0 16 11 7 11 11 2
14 1 9 0 9 13 3 0 9 9 1 3 0 9 2
30 13 1 9 2 0 2 10 9 9 9 2 15 0 9 9 9 13 1 15 2 16 0 9 2 15 13 2 3 13 2
9 1 0 9 13 7 0 0 9 2
23 12 0 0 9 13 0 9 9 12 0 9 2 0 9 11 11 7 0 9 11 11 11 2
19 2 9 13 3 7 2 16 4 15 9 1 15 13 2 2 2 11 2 2
22 2 0 2 15 15 9 1 9 13 2 13 2 16 15 1 9 13 2 2 2 11 2
17 13 3 1 0 9 2 16 4 13 2 15 1 15 12 13 9 2
2 9 11
30 9 0 9 15 13 9 11 11 7 0 9 9 9 11 11 1 9 9 12 2 9 1 9 2 4 11 13 2 2 2
6 13 15 3 9 9 2
47 9 0 9 13 2 16 2 10 9 3 0 9 1 11 7 10 0 9 11 2 15 3 3 3 13 9 1 9 0 9 2 4 13 1 12 7 12 9 13 0 9 1 9 10 9 2 2
30 9 3 13 0 9 9 2 16 4 13 10 9 2 1 15 1 9 1 0 9 13 0 9 0 9 7 9 10 9 2
3 2 11 2
2 11 2
3 9 1 11
13 9 11 1 9 9 7 0 9 9 9 7 0 9
2 11 11
27 9 11 13 2 16 0 9 2 0 1 11 9 0 9 7 9 2 13 3 3 3 9 0 9 0 9 2
28 3 15 13 2 16 0 9 15 9 1 9 0 9 13 13 3 7 14 3 2 16 13 13 1 0 9 9 2
16 0 7 0 0 9 1 9 7 11 10 9 13 11 9 12 2
13 9 0 11 2 0 7 3 0 11 2 13 0 2
24 9 9 9 0 9 1 11 15 13 9 1 0 0 9 2 15 15 3 13 0 9 9 9 2
43 1 0 9 0 9 2 3 15 13 1 11 7 3 3 1 0 9 2 13 1 0 9 0 9 1 9 7 9 7 9 0 9 7 9 0 9 13 9 11 7 0 9 2
21 1 9 0 9 13 0 9 1 0 0 9 9 7 0 9 3 13 13 0 9 2
21 9 9 9 1 10 9 15 13 2 16 7 1 9 0 9 4 13 13 1 9 2
17 1 0 9 15 3 13 0 9 1 0 9 7 13 15 0 9 2
4 7 7 3 2
24 15 3 0 9 13 2 15 0 13 9 0 9 11 7 15 0 13 9 9 0 9 0 9 2
20 11 3 0 9 13 10 9 1 9 9 7 3 0 9 9 9 7 0 9 2
47 7 16 4 13 3 0 2 15 13 1 11 9 2 9 11 11 13 9 11 1 9 7 9 0 9 1 15 2 16 15 15 13 1 15 9 7 1 9 1 11 13 13 1 9 0 9 2
20 13 15 15 13 2 16 9 15 1 10 9 13 13 0 9 1 10 0 9 2
45 9 7 11 3 1 2 3 0 2 9 9 1 11 13 0 9 2 0 7 0 9 1 0 9 2 16 4 13 0 9 11 7 11 2 13 10 9 7 13 9 9 7 0 9 2
12 11 3 3 13 13 1 9 2 16 13 15 2
23 0 9 15 13 10 9 2 7 3 4 15 13 13 10 9 1 9 1 9 11 7 11 2
16 13 15 0 16 11 2 16 0 9 15 13 13 2 16 13 2
19 0 9 3 7 13 0 9 2 16 4 4 13 9 1 9 9 1 11 2
5 11 15 13 13 2
10 10 9 13 3 0 2 7 3 0 2
26 13 15 13 2 16 1 0 9 13 14 0 11 2 0 0 7 0 9 7 9 11 2 11 7 11 2
22 9 13 13 7 0 9 15 13 2 16 13 13 0 2 16 0 9 0 9 15 13 2
5 3 13 9 13 2
11 7 3 13 2 16 15 15 13 0 9 2
5 11 4 13 9 2
7 3 15 4 13 0 9 2
18 1 9 11 0 9 3 3 13 9 9 0 9 7 0 9 1 11 2
12 11 2 9 2 11 7 11 14 13 13 9 2
5 16 11 1 11 2
7 9 1 12 9 13 13 0
8 11 11 2 9 2 13 1 11
14 1 0 0 9 13 14 12 9 9 1 0 0 9 2
25 0 12 9 2 3 11 2 15 13 7 13 1 11 2 4 0 13 9 0 2 7 13 13 0 2
36 9 1 0 0 9 13 14 1 11 2 7 7 1 11 7 1 11 7 2 16 9 10 9 13 2 16 4 10 9 13 7 13 0 0 9 2
25 9 9 13 0 9 0 9 1 11 7 0 9 13 9 9 2 15 4 1 11 13 0 0 9 2
45 10 9 13 0 9 2 15 3 13 3 1 0 9 1 0 9 2 13 1 12 7 1 3 9 9 11 7 1 9 12 13 3 1 0 0 9 2 13 3 0 0 9 7 9 2
13 13 1 9 0 9 13 1 11 3 3 3 0 2
24 0 0 9 3 1 0 9 0 9 2 15 15 13 0 0 9 2 0 9 13 7 3 13 2
36 7 9 13 2 16 0 0 2 7 0 2 9 2 15 13 9 11 7 1 9 12 13 1 0 2 15 1 3 0 9 13 1 11 3 9 2
33 1 0 9 13 0 0 9 1 0 0 9 1 9 2 3 3 13 0 0 9 2 13 0 0 9 0 9 2 9 7 0 9 2
51 1 11 4 3 13 16 9 2 15 4 2 16 15 11 13 2 13 2 16 4 15 13 2 3 15 13 13 7 9 0 1 11 2 3 13 0 9 1 9 7 9 2 7 4 15 13 13 1 10 9 2
51 0 9 13 7 9 0 2 7 14 1 9 2 0 9 13 13 2 15 1 0 0 2 0 9 13 3 9 11 2 15 3 2 13 1 12 9 2 2 16 10 9 10 10 9 1 0 9 3 3 13 2
38 13 15 7 3 9 2 16 11 2 9 15 1 9 7 9 1 9 1 0 0 9 1 9 13 9 2 7 0 0 9 15 13 12 2 0 7 0 2
42 1 11 13 9 9 1 3 3 0 9 2 0 0 9 2 3 0 9 11 2 13 1 9 0 9 0 0 0 9 2 0 0 9 7 0 9 2 15 13 0 9 2
26 16 4 0 9 13 13 9 1 9 2 15 15 0 9 13 2 13 15 3 13 9 1 12 0 9 2
31 7 16 13 0 10 9 7 9 9 2 15 3 7 3 1 9 13 0 9 2 0 15 1 10 9 3 7 3 3 13 2
2 0 9
7 9 2 11 11 9 0 9
3 2 11 2
41 11 9 11 15 13 1 9 9 9 2 16 4 9 7 9 13 13 7 1 0 9 1 3 0 9 2 1 15 15 13 1 11 2 2 2 7 0 9 0 11 2
43 7 16 9 10 9 13 2 13 3 12 1 0 9 2 0 9 1 9 0 9 2 15 4 13 3 2 16 9 1 9 2 13 15 1 9 2 7 7 1 15 13 9 2
10 10 9 1 0 9 13 1 0 9 2
20 9 10 0 9 13 9 9 3 0 9 2 1 15 13 9 7 3 7 9 2
24 13 15 3 9 10 0 9 10 9 0 1 0 9 13 14 3 0 2 16 13 1 0 9 2
62 7 16 4 13 2 9 9 13 1 9 9 2 15 13 0 2 1 9 2 7 15 1 10 9 2 16 3 13 0 9 2 7 3 15 1 0 9 13 1 0 9 2 16 4 13 9 9 2 7 15 9 1 9 0 1 9 0 9 7 9 9 2
22 10 9 15 3 1 9 13 2 9 2 7 7 1 0 9 1 9 13 13 0 9 2
17 13 7 1 10 0 0 9 2 15 4 13 10 9 1 10 9 2
48 3 7 16 4 1 9 13 13 0 9 2 13 15 13 0 9 2 3 15 1 12 13 9 9 2 15 4 3 13 0 9 7 15 13 0 2 16 4 15 2 3 13 2 13 0 0 9 2
41 16 15 3 3 9 0 1 9 9 13 1 9 9 9 7 1 15 15 1 0 9 13 1 10 9 1 9 13 0 9 2 3 13 0 0 9 13 7 10 9 2
14 1 3 0 7 13 9 13 1 9 1 9 0 9 2
47 9 1 0 9 2 0 9 7 0 9 9 13 13 1 0 0 7 3 0 2 16 0 9 9 2 16 1 9 1 9 13 3 10 9 2 0 0 9 2 9 2 9 7 9 0 9 2
24 15 4 3 13 13 1 15 2 16 13 9 1 10 9 0 7 16 13 3 13 1 0 9 2
19 13 0 13 1 0 9 2 16 3 13 2 10 9 13 0 9 3 13 2
19 13 1 9 13 9 9 13 0 7 0 3 13 2 16 9 9 3 13 2
17 16 9 1 9 9 13 3 0 2 7 7 15 1 15 3 13 2
21 15 1 15 2 16 15 13 0 9 7 16 15 13 1 0 16 9 9 7 9 2
32 15 4 13 1 15 2 16 13 13 9 9 0 12 7 12 12 9 2 7 3 3 13 2 14 1 9 0 10 3 0 9 2
26 16 13 9 9 1 15 0 16 1 0 9 2 13 4 3 13 2 15 13 9 10 9 7 10 9 2
16 9 0 9 4 15 3 13 13 7 13 1 10 9 0 9 2
25 7 3 1 9 2 16 13 0 13 1 10 9 0 0 9 2 16 14 2 13 0 9 3 13 2
16 1 9 1 15 2 10 9 15 15 13 13 1 9 0 9 2
4 0 9 13 9
9 0 9 15 13 13 9 7 0 9
2 9 9
7 9 1 9 13 13 9 2
23 0 9 2 15 15 3 13 14 1 10 9 1 9 2 4 13 3 1 9 9 3 13 2
29 1 0 0 7 0 9 15 13 13 7 1 0 2 3 9 9 2 9 9 7 3 9 2 15 13 3 0 9 2
23 9 7 10 9 13 1 9 1 9 0 2 7 1 10 9 15 13 2 16 13 0 9 2
5 9 1 9 1 9
11 12 9 1 0 9 4 13 3 0 9 2
7 0 9 13 13 7 1 9
2 9 9
20 1 0 9 15 3 3 13 2 16 10 9 0 9 13 0 0 9 16 0 2
14 13 15 13 10 9 2 0 9 2 9 0 9 3 2
24 1 15 2 10 9 15 10 9 13 9 9 2 4 13 1 9 9 11 11 9 2 11 2 2
17 11 11 1 9 9 13 1 9 0 2 9 0 9 1 0 9 2
18 10 9 15 10 9 13 13 16 4 13 1 0 9 9 1 0 9 2
15 2 0 9 2 3 13 0 9 2 13 13 0 0 9 2
21 13 1 15 2 15 1 11 13 2 15 9 13 13 1 9 7 9 9 0 9 2
17 13 0 9 9 9 2 9 9 2 9 2 9 7 9 0 9 2
19 3 13 9 2 3 13 13 0 9 2 16 1 15 13 1 0 9 9 2
16 13 0 9 13 7 3 2 16 15 13 13 7 1 9 0 2
11 1 15 2 15 13 13 2 0 9 13 2
20 9 0 9 2 15 15 1 0 9 13 13 2 13 1 15 2 16 13 9 2
9 1 10 9 13 9 9 0 2 2
4 13 13 0 2
24 2 3 10 9 13 0 0 7 0 9 2 15 9 9 3 13 2 7 13 9 1 0 9 2
13 3 13 0 9 9 2 0 1 0 7 0 9 2
20 1 15 15 3 13 3 9 2 15 13 1 9 11 2 11 2 11 7 11 2
18 13 1 9 2 16 11 15 13 7 4 3 13 3 0 9 16 3 2
13 3 3 13 1 9 0 9 10 9 1 0 9 2
5 15 15 3 13 2
20 9 3 13 15 2 16 1 15 4 13 0 0 9 2 9 2 0 9 3 2
11 16 4 13 2 4 1 9 3 13 9 2
36 7 0 9 3 13 2 16 16 13 13 1 9 7 13 9 2 13 3 13 3 9 0 9 7 15 15 3 13 3 3 2 16 10 9 13 2
10 15 1 15 3 3 13 0 9 2 2
23 10 0 9 1 0 9 13 1 15 2 16 0 9 15 13 13 1 0 11 7 0 11 2
3 13 9 2
13 2 3 1 9 13 2 16 9 0 9 13 0 2
11 15 13 13 3 2 0 9 2 9 3 2
9 1 10 9 15 13 3 0 9 2
11 12 1 9 0 9 13 13 10 0 9 2
24 7 14 15 2 16 4 15 1 0 9 13 0 9 2 15 4 1 15 13 16 1 0 9 2
12 13 15 13 9 9 2 7 3 0 9 9 2
12 13 3 10 9 1 11 3 0 16 1 11 2
18 2 13 15 2 16 15 3 13 1 10 0 9 2 15 13 3 0 2
18 13 15 2 16 11 13 1 15 2 16 4 13 3 3 0 16 11 2
13 3 13 2 16 4 13 13 0 7 13 0 9 2
20 3 13 9 2 16 1 0 9 13 1 9 0 3 0 0 9 16 14 11 2
30 3 11 2 13 15 2 16 13 14 0 2 7 1 10 9 3 0 7 13 10 9 7 16 15 13 9 0 9 2 2
21 7 1 10 9 2 3 1 9 11 2 11 7 0 11 2 13 3 3 0 9 2
13 13 15 2 16 7 15 13 0 9 13 3 0 2
8 2 10 9 4 13 0 9 2
22 16 3 7 3 4 1 15 13 0 9 9 16 3 2 9 1 10 9 13 0 9 2
12 3 13 14 1 15 2 16 4 4 3 13 2
17 13 0 2 16 4 0 9 1 9 1 9 9 13 10 0 9 2
13 13 13 2 16 1 15 13 3 9 2 7 14 2
12 7 13 15 9 2 15 9 3 13 13 2 2
13 7 13 10 0 9 1 10 9 0 2 7 14 2
3 2 13 2
22 1 9 9 7 0 9 4 13 0 9 2 1 15 4 15 9 1 10 9 3 13 2
21 0 9 4 13 0 9 1 9 0 9 7 9 1 10 9 3 1 9 3 13 2
13 15 13 13 2 16 9 13 3 0 7 3 0 2
23 3 14 9 0 9 9 2 15 4 0 9 13 0 9 10 9 2 15 9 3 13 2 2
15 10 9 15 13 1 9 1 9 0 0 9 0 2 11 2
16 3 3 3 9 13 9 2 16 13 9 1 9 10 9 0 2
13 13 15 2 16 9 1 10 0 9 13 3 13 2
8 2 9 13 3 13 0 9 2
23 13 9 2 16 1 9 15 3 15 13 13 9 2 16 13 4 15 13 3 7 0 9 2
11 3 3 13 1 15 2 16 3 13 4 2
8 7 15 13 9 2 15 13 2
13 15 13 1 15 0 0 9 2 3 1 9 9 2
32 3 15 1 15 13 2 3 15 13 2 12 9 15 1 10 9 13 7 3 3 15 13 9 1 15 2 16 4 13 13 3 2
12 1 0 9 11 2 0 15 15 13 0 2 2
12 15 3 15 1 10 9 4 1 0 9 13 2
59 2 1 1 15 2 16 9 0 0 9 15 1 9 1 0 9 13 0 0 9 2 13 9 1 9 10 9 1 12 2 12 9 1 9 1 9 9 2 12 2 12 1 9 9 1 9 11 1 11 2 9 1 11 2 9 11 7 11 2
16 0 9 1 9 0 1 9 0 9 9 13 13 1 9 11 2
25 13 9 9 9 1 9 11 7 0 4 13 1 9 9 9 2 15 13 9 12 2 9 0 9 2
14 9 0 9 13 0 9 11 2 10 9 13 9 9 2
16 0 9 9 9 1 9 11 3 13 13 7 13 1 0 9 2
26 9 9 1 0 9 13 7 9 0 9 0 9 7 9 11 2 15 0 9 3 4 13 12 2 9 2
15 0 9 9 9 0 0 9 13 7 9 0 3 0 9 2
11 9 0 9 4 13 1 9 0 9 11 2
18 0 9 1 11 7 0 13 13 7 13 2 3 13 9 10 9 2 2
3 9 11 11
11 9 9 2 1 9 1 9 12 7 1 9
11 0 9 0 0 9 0 11 1 9 1 11
2 9 11
19 0 0 9 1 12 9 13 0 0 9 16 9 15 1 9 0 0 9 2
4 4 3 13 2
12 3 3 15 13 0 9 1 11 1 0 9 2
14 0 0 9 15 13 9 9 1 9 7 4 3 13 2
15 3 1 10 12 2 9 15 0 9 13 9 1 0 9 2
14 13 15 2 3 15 3 3 13 7 13 0 0 9 2
24 4 1 0 0 7 0 9 7 9 3 13 16 9 1 0 9 9 7 9 0 9 1 9 2
19 9 2 13 9 1 0 0 9 2 15 13 13 9 14 1 12 2 9 2
12 9 13 7 1 0 9 10 9 2 3 0 2
17 14 1 9 12 15 13 13 2 16 0 9 4 13 7 13 9 2
11 15 13 9 2 13 15 9 0 2 0 2
18 13 4 15 2 3 1 9 12 13 0 0 9 10 0 9 1 9 2
25 13 4 15 2 16 1 9 12 4 13 9 9 1 0 11 2 16 13 10 9 2 7 3 15 2
29 0 9 10 12 9 2 3 15 9 13 0 9 2 4 13 14 0 9 0 9 2 15 3 11 1 12 9 13 2
19 1 9 9 15 13 11 2 9 2 11 2 9 2 9 7 9 15 9 2
10 13 1 3 12 9 10 12 0 9 2
10 10 15 0 7 0 13 0 13 9 2
10 9 13 9 11 7 0 9 1 9 2
12 0 9 13 3 1 11 2 7 3 13 13 2
13 0 9 13 1 11 2 1 11 7 1 0 9 2
14 0 9 3 13 0 9 7 13 9 13 10 0 9 2
12 0 0 9 9 1 11 13 9 9 1 9 2
23 3 0 9 2 13 15 14 1 12 12 2 13 9 9 7 9 12 0 0 9 1 9 2
14 13 15 9 7 9 12 0 9 0 9 7 10 9 2
6 1 9 9 11 2 11
5 9 9 1 9 12
4 9 11 2 9
14 3 2 16 13 15 13 2 11 12 2 12 2 12 2
7 3 3 15 9 11 13 2
15 13 13 9 3 0 1 9 1 0 9 0 9 0 9 2
27 13 1 9 2 12 9 2 15 15 1 9 7 12 9 13 2 7 16 3 3 2 13 4 3 0 9 2
21 9 9 12 4 13 3 1 9 7 9 13 3 14 1 0 9 16 0 9 9 2
25 9 13 7 0 13 3 1 9 1 0 9 2 16 4 3 13 1 9 3 2 16 0 9 13 2
70 0 9 1 0 9 9 2 9 7 9 13 13 12 2 9 2 13 15 3 13 0 2 16 1 9 7 9 13 0 2 7 16 9 13 2 16 15 13 7 3 2 9 9 12 9 2 1 12 2 0 9 2 13 7 9 1 15 4 13 13 2 13 3 0 9 2 1 0 9 2
31 14 9 2 9 15 13 1 9 2 7 3 13 2 16 13 13 3 16 13 2 7 3 1 9 15 13 9 15 3 13 2
10 1 0 9 15 7 13 13 9 0 2
12 1 9 9 15 15 13 3 1 9 2 13 2
15 1 15 15 13 0 2 16 9 13 13 1 12 2 9 2
47 4 3 0 9 13 0 9 2 3 13 1 10 9 13 1 10 9 3 2 13 4 3 13 13 3 15 7 3 15 15 9 4 13 2 16 1 0 9 13 10 0 9 2 13 0 9 2
3 9 9 2
11 0 9 15 9 13 2 15 15 13 9 2
39 1 15 2 16 4 1 9 7 0 9 1 9 13 2 13 13 9 1 0 9 7 3 9 1 9 3 2 16 15 1 0 9 10 9 13 1 12 9 2
3 3 0 2
21 1 10 9 7 0 9 13 13 2 7 0 15 13 1 0 9 2 4 13 13 2
25 6 2 16 15 13 2 3 15 13 3 1 0 0 9 2 3 0 9 13 1 0 9 3 3 2
8 1 9 9 4 13 9 9 2
7 13 9 9 7 9 3 2
18 1 9 4 1 15 13 9 2 11 11 12 15 1 15 3 13 9 2
6 1 9 11 11 2 11
14 3 2 16 13 15 13 2 11 12 2 12 2 12 2
7 3 3 15 9 11 13 2
21 9 9 12 4 13 3 1 9 7 9 13 3 14 1 0 9 16 0 9 9 2
15 7 9 4 13 1 9 9 2 11 12 2 12 2 12 2
6 13 3 0 9 0 2
14 9 1 9 1 9 12 13 12 5 0 0 0 9 2
20 1 0 9 13 0 2 16 15 0 9 13 1 12 2 12 5 0 0 9 2
15 0 0 9 13 0 9 9 7 1 10 9 13 10 9 2
18 9 13 3 1 15 2 16 9 13 0 1 0 9 7 1 0 9 2
16 16 4 1 9 9 4 13 3 2 13 13 9 10 0 9 2
7 0 9 13 3 10 0 2
28 1 0 0 9 4 13 1 9 1 15 12 5 9 1 9 13 9 11 7 15 13 0 9 1 0 0 9 2
20 9 13 1 9 9 1 9 0 9 0 1 0 9 2 0 9 7 0 9 2
30 3 13 3 3 0 2 16 13 0 9 2 16 1 9 9 4 13 0 9 11 2 7 15 3 7 1 0 0 9 2
20 0 7 0 9 0 9 13 9 0 9 7 3 3 14 9 1 9 2 12 2
27 9 13 3 14 12 9 1 9 2 15 13 9 0 0 9 9 2 7 13 9 1 9 9 9 7 9 2
27 3 1 10 9 13 0 2 16 9 1 10 9 13 3 3 0 9 0 9 2 15 13 2 7 13 15 2
18 3 3 15 13 2 16 9 1 9 0 9 13 1 0 9 9 9 2
33 9 0 9 7 9 2 15 0 9 3 3 13 2 13 3 0 2 16 15 15 3 7 3 13 9 2 15 13 1 0 0 9 2
17 13 4 0 13 2 16 0 0 9 9 9 1 0 9 3 13 2
16 16 15 15 3 13 2 13 15 3 13 9 9 7 0 9 2
6 1 9 11 11 2 11
4 1 0 9 9
14 1 0 9 10 9 4 13 12 0 9 7 1 9 2
23 13 1 0 11 7 11 2 15 15 13 13 9 7 13 2 16 15 1 15 13 15 13 2
7 13 1 9 2 1 9 2
17 13 12 9 0 3 0 2 3 3 0 9 2 7 15 15 13 2
16 13 15 1 0 9 7 3 15 13 7 13 2 13 0 9 2
9 10 9 13 9 1 9 1 9 2
11 12 10 9 7 13 9 9 3 1 9 2
15 9 13 1 9 2 13 1 9 7 3 15 13 1 9 2
26 7 6 2 11 3 13 2 0 2 9 2 15 3 3 3 10 0 9 13 2 15 13 1 0 9 2
53 16 15 3 13 1 9 2 13 9 7 13 9 7 13 2 16 15 13 10 9 2 9 7 0 2 16 15 3 13 13 15 16 9 0 9 0 9 0 9 3 2 3 13 13 9 0 2 13 13 1 10 9 2
44 16 4 13 1 9 9 3 9 9 11 2 3 4 15 9 9 13 2 16 1 9 0 2 15 1 9 7 1 9 15 13 2 13 0 13 3 0 9 0 2 15 13 0 2
65 13 2 14 9 11 1 9 2 1 15 9 2 3 1 9 2 2 16 15 13 9 10 0 9 2 13 15 2 16 4 1 10 9 13 1 0 9 2 13 13 1 9 2 16 4 13 2 16 10 0 9 13 1 9 9 2 9 9 7 9 1 9 3 0 2
17 15 13 9 2 16 4 3 7 3 13 13 1 9 2 1 9 2
35 10 9 9 13 13 1 9 2 16 4 13 3 1 9 0 9 2 1 15 2 16 15 13 0 2 3 2 16 13 1 0 7 0 9 2
21 16 4 9 9 11 15 13 2 16 13 1 15 9 2 3 4 15 13 1 9 2
18 15 15 7 7 10 0 9 3 13 7 13 15 2 16 13 15 0 2
20 3 15 15 3 13 2 16 9 2 9 2 10 9 13 1 9 9 1 9 2
30 13 15 2 1 10 9 13 1 15 2 16 4 15 1 9 13 0 0 9 2 7 1 9 0 9 7 1 0 9 2
27 7 13 9 2 16 0 9 13 3 2 15 15 13 2 3 14 13 3 13 2 15 15 13 15 3 0 2
32 3 13 9 2 16 13 0 15 3 13 2 16 9 0 0 9 13 0 7 15 13 2 16 10 9 13 0 2 0 2 0 2
32 3 15 15 13 2 16 13 1 10 0 9 2 7 15 4 15 13 13 13 1 9 2 15 4 13 2 16 13 1 9 0 2
18 13 4 15 13 2 16 4 13 9 2 1 9 2 15 13 1 9 2
11 3 15 1 10 9 3 13 2 7 15 2
18 13 3 13 0 9 9 7 13 15 1 9 9 9 3 2 9 3 2
6 13 2 16 15 13 2
8 11 11 2 11 13 9 2 11
12 15 13 1 9 2 11 12 2 12 2 12 2
19 13 15 2 16 16 9 13 9 13 15 3 1 9 15 2 15 4 13 2
17 7 3 1 15 13 2 16 4 13 1 9 9 2 0 9 2 2
19 1 9 2 0 2 15 13 15 7 3 15 13 2 2 3 13 9 2 2
21 13 0 2 16 3 13 0 1 0 9 7 3 9 1 0 9 7 9 15 13 2
8 13 3 13 9 9 16 9 2
6 1 9 11 11 2 11
2 13 9
14 3 14 10 9 15 13 10 9 9 2 16 9 0 2
22 10 9 15 13 3 1 9 1 0 9 0 9 7 13 3 1 9 13 15 10 9 2
29 1 0 1 15 15 10 0 7 0 9 13 9 9 7 0 9 7 9 15 15 13 7 1 9 13 7 13 15 2
30 1 15 15 7 7 15 13 1 9 0 1 0 9 7 10 9 3 13 2 12 1 0 9 13 3 9 0 0 9 2
31 3 7 13 1 10 9 9 9 0 7 12 1 12 9 0 0 9 0 2 1 15 15 13 9 7 9 9 1 0 11 2
19 9 10 0 9 13 1 0 9 10 9 7 4 3 13 1 10 0 9 2
14 0 2 1 9 3 0 0 9 13 3 1 9 12 2
34 13 7 15 2 15 13 0 9 10 0 9 7 13 4 13 1 10 9 2 16 4 15 3 3 13 1 0 9 1 10 3 0 9 2
29 7 15 2 15 15 9 13 13 2 7 3 4 13 10 10 0 9 13 2 0 9 9 3 13 9 0 9 9 2
12 0 0 9 2 0 2 9 2 9 12 2 11
34 15 2 3 2 3 12 2 12 2 2 0 9 1 0 11 13 3 2 12 2 1 9 9 11 11 11 1 9 11 11 13 2 9 2
28 0 9 13 3 3 2 12 2 9 0 0 9 1 9 11 11 13 2 9 2 7 1 11 11 1 0 9 2
25 9 1 9 11 11 13 1 9 1 0 9 11 1 11 2 0 9 2 2 1 12 2 9 2 2
22 0 0 9 13 3 2 12 2 0 1 10 9 1 9 11 2 15 13 9 11 9 2
8 9 13 0 9 9 9 11 2
25 0 9 9 2 9 0 9 11 11 0 9 7 0 9 11 13 1 0 0 9 1 9 0 9 2
19 3 15 13 1 3 0 0 9 9 2 16 4 13 1 9 12 0 9 2
21 1 15 3 13 0 0 9 11 11 7 9 11 11 2 1 10 9 15 9 13 2
18 1 9 1 0 4 2 3 1 0 9 11 11 2 13 9 9 11 2
8 3 15 9 13 1 0 9 2
26 15 4 3 13 1 0 9 2 1 9 2 9 2 11 0 2 7 2 0 2 9 2 11 11 2 2
18 10 9 9 13 1 0 9 0 9 0 1 3 0 9 2 9 9 2
11 2 1 9 0 9 2 9 11 11 2 2
14 1 15 15 13 9 2 9 2 0 9 2 3 9 2
28 9 9 2 10 9 7 9 2 13 11 15 0 9 2 3 0 0 7 0 9 1 9 0 2 7 3 0 2
30 9 0 9 2 3 0 9 7 0 9 13 3 13 1 0 9 9 7 9 2 7 1 0 9 9 13 15 3 0 2
12 3 15 15 13 1 0 9 1 9 11 11 2
25 15 15 3 13 3 1 9 0 9 10 9 2 3 7 15 15 13 2 16 2 9 13 9 2 2
30 0 9 2 0 9 13 9 13 9 2 0 2 2 0 2 11 13 1 9 9 2 16 4 13 2 15 15 7 13 2
16 11 13 1 9 3 12 1 0 9 2 13 9 10 0 9 2
34 9 0 1 15 2 16 4 4 9 13 2 16 2 9 2 4 0 3 2 1 0 9 7 1 9 13 15 0 9 2 13 0 9 2
27 0 2 3 0 9 0 13 9 7 11 11 16 11 2 10 0 9 2 9 1 9 2 13 0 9 9 2
14 1 0 9 9 7 3 15 13 1 0 9 0 9 2
13 9 0 9 3 13 3 7 3 3 10 0 9 2
30 10 0 9 13 11 11 1 9 2 3 4 13 13 9 0 9 0 7 15 13 12 1 0 9 1 0 9 0 9 2
7 13 15 1 15 3 9 2
21 11 11 9 2 11 11 7 11 11 1 9 0 9 7 0 9 11 1 0 9 9
3 9 11 11
34 11 2 0 3 2 9 9 2 12 1 3 0 0 0 9 9 2 0 11 2 0 2 13 1 9 3 1 0 9 11 1 0 11 2
8 9 13 0 9 0 9 11 2
10 1 11 13 9 2 9 7 0 9 2
40 9 11 11 1 12 9 9 9 13 1 12 1 0 9 0 0 9 2 3 7 0 9 2 7 16 4 15 3 13 2 11 15 1 15 3 13 0 9 9 2
20 0 9 1 9 13 0 9 9 11 10 13 11 2 0 9 0 1 9 11 2
17 3 3 0 0 9 11 13 1 9 1 9 0 9 2 0 11 2
18 9 10 9 16 16 4 15 13 1 9 12 2 3 13 10 0 9 2
16 0 0 9 11 13 3 0 2 16 3 1 9 0 2 9 2
52 10 9 3 13 7 9 0 9 9 2 7 16 13 9 2 16 9 9 2 0 3 13 3 0 7 1 0 9 11 11 2 9 2 2 11 11 2 9 2 7 9 11 2 0 2 10 0 0 9 13 9 2
20 7 0 9 9 2 9 11 11 13 1 9 3 14 1 9 2 7 2 2 2
43 1 9 1 9 2 11 2 0 2 13 1 15 2 11 3 2 9 3 13 3 3 7 3 7 10 9 9 13 15 2 3 2 2 15 2 15 13 0 9 3 0 9 2
12 13 15 3 9 2 7 9 2 13 2 14 2
43 13 2 16 9 9 2 0 13 9 0 9 0 9 2 4 13 0 2 7 3 1 11 15 9 13 13 2 1 15 3 9 7 2 9 2 13 1 9 3 3 0 11 2
15 0 9 2 15 15 9 12 1 0 13 2 3 13 15 2
51 0 1 9 15 3 9 2 0 3 13 1 10 0 2 2 0 2 9 2 15 13 11 9 2 3 1 11 11 2 7 9 10 13 1 15 2 15 13 3 0 9 9 2 3 1 11 0 16 0 9 2
13 3 1 11 13 0 9 2 0 2 9 2 2 2
2 11 9
6 9 9 2 9 3 13
20 9 9 2 9 13 1 9 12 9 11 11 2 9 11 11 7 9 11 11 2
25 3 1 15 13 3 12 0 9 7 4 13 1 12 9 2 0 15 3 0 0 9 7 0 9 2
39 16 10 0 9 13 9 2 9 3 2 11 12 2 12 2 0 9 9 1 9 1 9 9 2 9 2 11 11 2 2 0 9 1 9 0 9 1 11 2
33 11 11 0 9 9 9 2 9 3 13 0 0 9 9 11 11 2 1 9 13 1 12 2 3 3 1 11 9 3 1 11 12 2
27 2 10 9 13 9 9 2 0 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 11 2 9 2
13 3 13 2 3 15 9 10 9 13 7 15 2 2
15 3 0 0 9 11 9 1 9 12 1 10 0 0 9 2
11 2 7 3 15 13 13 3 1 9 0 2
11 13 2 16 4 15 9 10 9 13 9 2
26 10 9 3 13 1 9 13 3 3 2 16 0 3 0 9 2 2 13 9 9 11 2 11 11 11 2
7 2 3 13 1 9 9 2
36 10 9 15 3 13 1 0 0 9 2 1 0 9 4 13 9 1 0 9 2 15 10 9 3 13 2 1 0 11 9 4 13 9 2 2 2
16 1 9 10 0 9 13 1 9 9 9 0 9 2 2 13 2
7 7 15 9 2 9 13 2
36 2 11 11 13 9 1 0 7 0 7 1 15 2 16 12 7 0 13 9 2 11 11 15 13 1 12 9 13 1 9 10 9 1 0 9 2
29 11 9 13 0 2 0 9 2 2 11 11 3 13 9 10 9 1 9 7 3 9 2 15 15 13 1 0 9 2
19 11 11 13 0 9 1 9 7 9 0 0 9 2 2 13 11 11 11 2
23 9 11 11 0 9 16 13 15 1 9 2 0 9 1 11 3 13 7 15 15 3 13 2
13 3 13 2 3 2 16 1 9 13 9 3 0 2
18 3 15 13 13 9 10 9 2 15 15 9 10 9 3 13 0 9 2
13 16 13 0 9 2 13 15 15 1 0 9 9 2
11 1 0 9 13 10 9 3 0 0 9 2
13 1 0 0 9 4 1 9 3 13 0 9 9 2
16 13 15 0 9 12 9 2 11 11 2 11 11 7 11 11 2
31 9 4 13 13 9 1 0 9 7 3 0 0 9 2 14 12 9 0 2 2 3 15 4 13 0 0 7 0 0 9 2
14 9 15 9 9 13 1 9 2 7 15 1 0 9 2
18 9 9 13 2 16 4 3 13 13 9 0 9 2 3 3 13 9 2
14 9 1 9 13 9 1 9 0 9 1 10 0 9 2
17 0 9 15 13 13 14 1 0 9 7 1 9 9 13 0 9 2
18 1 11 4 3 13 7 0 9 2 7 4 9 9 13 13 3 0 2
6 9 9 13 3 0 2
22 12 9 9 13 2 16 0 9 13 0 13 9 7 13 15 7 13 1 0 0 9 2
20 9 4 13 13 7 0 9 9 11 11 2 12 2 2 9 0 9 0 9 2
12 11 13 1 9 2 15 13 10 9 0 9 2
23 3 13 1 11 11 1 0 9 1 9 2 1 0 9 15 13 0 9 1 11 7 9 2
10 13 9 9 3 0 0 9 1 11 2
24 0 9 9 4 13 0 9 2 0 1 9 1 9 9 2 13 15 1 15 9 0 9 11 2
29 9 13 9 3 9 0 0 0 9 2 3 3 13 3 2 11 0 2 11 11 2 11 11 2 11 11 7 0 2
15 0 9 1 15 9 13 4 2 10 9 4 10 9 13 2
9 1 9 13 7 0 9 1 9 2
21 3 13 9 10 3 9 7 15 0 1 0 9 1 9 2 3 3 13 0 9 2
3 0 9 13
7 3 9 13 1 11 7 11
20 0 9 9 9 0 11 11 13 10 9 0 9 1 9 9 7 9 0 9 2
17 1 0 9 13 1 0 9 1 9 0 0 9 13 12 12 9 2
10 9 13 12 9 0 3 1 12 9 2
27 2 0 9 2 0 16 0 9 10 0 9 2 13 1 0 9 12 9 2 15 4 13 1 12 9 2 2
10 0 9 3 13 12 9 1 12 9 2
25 0 9 2 12 12 2 13 1 0 9 0 9 11 11 2 15 1 0 9 9 13 9 11 11 2
12 0 9 13 3 1 9 11 11 7 11 11 2
22 2 3 13 0 9 2 16 0 9 13 9 3 2 2 13 10 9 9 9 11 11 2
19 2 7 13 16 12 1 9 15 2 16 13 9 1 9 7 0 9 2 2
28 0 0 9 2 12 12 2 13 1 9 9 0 9 9 11 11 2 15 15 3 13 0 0 9 2 0 9 2
29 9 11 13 11 11 2 3 9 9 2 3 16 11 11 7 3 11 11 2 9 0 9 2 15 13 12 9 2 2
27 2 16 9 13 9 2 1 15 13 15 1 10 9 13 2 1 9 13 3 1 9 13 2 2 13 11 2
21 2 9 0 9 2 1 15 4 15 9 14 13 13 2 13 3 13 2 2 2 2
9 15 1 0 9 13 1 0 9 2
32 3 3 11 2 9 9 4 15 13 13 9 9 9 2 15 15 13 7 13 3 3 2 11 11 2 11 2 9 12 12 2 2
24 1 1 0 9 9 0 9 13 9 3 7 9 11 9 1 11 2 11 2 9 12 12 2 2
3 2 11 2
3 9 0 9
26 9 0 7 0 9 9 2 12 11 1 11 13 1 15 1 12 9 3 12 9 7 10 0 0 9 2
23 1 9 1 0 9 2 15 15 13 1 9 12 7 13 3 0 2 13 15 0 3 0 2
4 11 11 2 11
25 13 15 3 1 15 2 16 9 0 9 13 9 9 9 7 9 2 7 3 15 13 1 9 9 2
27 2 13 4 1 0 9 9 7 10 9 13 13 10 9 0 9 2 2 13 0 9 0 0 9 11 11 2
9 2 9 9 13 1 10 0 9 2
12 13 1 0 9 2 7 3 1 9 0 9 2
16 13 4 15 2 16 4 0 9 13 0 9 3 0 9 2 2
21 0 9 13 0 9 1 9 0 9 2 7 3 16 1 0 15 15 13 0 9 2
22 2 13 15 7 15 2 15 13 15 9 2 16 4 15 15 3 13 2 2 13 11 2
15 2 1 15 4 13 2 16 4 9 13 9 3 1 11 2
13 12 9 1 9 12 9 2 15 13 13 0 9 2
24 11 13 12 12 9 7 0 9 15 3 13 3 3 1 9 1 3 16 12 12 9 2 2 2
14 13 10 9 1 9 13 9 9 2 15 13 10 9 2
12 7 16 4 13 0 2 15 4 1 15 13 2
16 0 9 2 10 13 0 9 2 0 9 1 12 9 9 13 2
11 2 0 9 9 13 9 7 9 0 9 2
10 0 9 4 15 0 13 3 16 9 2
36 0 9 15 7 1 11 13 3 2 16 9 11 15 13 1 3 0 9 2 15 13 9 9 3 1 0 9 2 0 1 0 9 1 9 0 2
19 1 15 13 9 9 0 9 2 15 4 15 13 13 1 9 0 9 9 2
13 1 15 1 9 13 3 0 9 0 0 9 9 2
3 0 9 11
5 9 13 9 1 11
2 9 9
23 2 9 11 2 11 9 2 11 11 2 11 11 2 13 10 0 9 1 0 11 0 11 2
28 13 1 0 9 7 13 1 15 1 0 9 13 9 14 12 2 15 9 2 7 13 1 15 2 0 13 2 2
12 1 10 0 9 13 0 9 11 12 0 9 2
22 9 13 11 11 2 15 3 13 3 1 11 11 2 11 2 11 11 2 11 2 11 2
10 2 1 11 13 3 12 9 9 11 2
13 0 12 9 13 0 7 0 9 9 1 0 11 2
40 1 9 0 9 1 0 9 2 1 15 13 1 9 9 9 11 11 9 3 7 3 0 16 1 9 0 2 13 14 11 11 13 3 7 2 13 15 9 2 2
22 16 11 15 13 0 10 9 1 9 2 9 11 13 9 10 9 7 13 15 1 9 2
10 3 15 13 2 16 13 14 0 9 2
19 11 15 13 2 16 0 16 0 9 13 9 2 1 15 3 3 13 13 2
32 1 10 9 13 0 9 9 11 1 0 7 0 9 2 15 13 3 12 2 9 1 11 7 13 4 13 12 2 9 1 11 2
32 0 9 0 1 12 2 9 1 9 11 4 3 13 1 0 0 9 1 9 7 4 3 13 3 0 9 7 9 1 0 9 2
41 9 11 13 12 7 12 9 7 1 9 9 13 3 3 7 9 11 11 2 1 0 9 13 3 1 9 9 2 7 1 9 11 11 2 3 14 9 11 7 9 2
13 1 0 9 1 11 7 11 15 13 1 12 9 2
8 3 13 10 9 1 9 9 2
15 2 13 4 1 9 7 10 9 15 13 2 2 13 11 2
19 2 13 4 1 11 2 16 4 13 13 1 9 2 15 1 15 13 2 2
3 2 11 2
2 11 2
17 0 9 0 11 2 11 13 1 0 9 1 11 9 1 0 9 2
23 1 9 15 0 0 9 13 1 11 2 3 15 9 9 2 9 2 13 1 9 0 9 2
24 0 9 13 3 9 11 7 9 10 9 15 1 9 13 1 0 1 9 0 9 11 2 11 2
20 11 13 3 1 11 7 0 1 9 13 1 9 0 9 11 2 11 2 11 2
26 1 9 15 15 1 9 1 11 13 9 2 15 13 1 0 9 1 9 2 3 11 7 11 2 11 2
20 1 9 11 2 11 13 0 9 0 9 1 12 9 2 3 1 9 11 12 2
20 3 0 9 1 0 12 0 9 15 4 13 1 9 1 11 12 1 12 9 2
21 11 11 1 11 11 9 11 13 0 9 1 0 9 9 0 9 11 1 0 11 2
16 11 11 1 9 11 11 9 11 15 13 0 9 11 1 9 2
6 14 9 1 0 9 13
16 9 0 0 9 11 11 13 3 3 9 13 15 2 15 15 13
2 9 9
56 2 15 15 15 13 1 10 9 2 2 2 13 15 15 10 0 9 9 1 0 9 1 9 0 9 2 11 12 2 12 2 3 9 9 11 11 0 1 9 3 13 2 16 15 0 9 10 9 13 9 1 0 9 1 11 2
35 0 9 11 1 11 1 11 11 11 13 9 3 3 0 1 0 9 2 7 10 0 9 13 15 15 2 16 3 3 3 3 3 13 13 2
28 13 15 2 16 11 11 7 11 0 13 3 3 14 10 0 9 1 0 9 2 15 15 3 15 1 15 13 2
15 10 9 13 1 0 9 9 1 11 1 11 3 0 9 2
19 1 3 0 9 1 9 1 11 2 12 2 12 2 13 3 0 9 9 2
22 3 13 9 12 9 1 11 2 1 0 9 4 13 12 9 7 13 12 2 12 2 2
38 3 3 4 13 1 11 2 12 2 12 2 2 15 15 1 9 0 9 9 0 9 13 1 9 1 9 3 3 16 3 3 2 7 3 15 15 13 2
14 9 7 0 9 13 9 1 11 2 12 2 12 2 2
12 3 1 15 15 1 10 9 13 9 1 9 2
27 16 9 1 0 11 3 13 1 9 7 0 9 2 9 9 11 0 13 9 1 2 3 0 2 2 2 2
46 9 1 9 2 0 13 9 1 12 9 1 0 9 9 7 15 2 15 0 9 7 0 9 13 1 0 9 9 13 1 0 9 7 10 0 9 9 9 2 15 3 13 1 0 9 2
29 13 9 3 0 11 11 2 16 1 0 9 1 0 9 3 13 10 9 7 1 9 2 15 15 1 11 13 13 2
43 2 16 13 9 11 11 2 13 2 2 13 15 1 10 0 9 2 3 15 13 2 16 15 16 0 13 9 11 1 9 9 1 9 12 1 11 13 1 0 9 1 9 2
16 13 2 16 4 10 9 13 7 10 0 9 10 0 9 2 2
25 9 0 9 4 15 7 7 1 10 9 2 3 9 0 9 3 13 2 13 3 13 1 0 9 2
25 1 1 9 0 9 4 13 13 0 9 9 2 1 15 13 9 16 0 7 0 9 14 0 9 2
40 13 13 3 0 1 9 2 16 15 13 0 9 13 2 16 13 9 13 0 0 9 7 13 15 3 1 9 2 15 2 1 9 2 13 9 0 9 1 9 2
30 14 13 11 11 13 10 0 7 0 9 2 0 1 0 9 2 13 4 13 2 16 9 7 9 1 9 3 15 13 2
22 1 9 2 1 9 0 0 0 9 2 13 3 7 9 9 7 0 9 13 1 9 2
18 1 9 7 13 2 16 13 1 9 9 2 9 15 15 1 9 13 2
8 11 11 15 3 3 13 13 2
12 13 15 13 2 7 13 15 2 15 15 13 2
9 13 1 9 16 9 2 2 2 2
6 13 10 3 0 9 2
20 13 13 1 15 2 3 13 2 7 12 9 1 15 13 7 3 13 1 11 2
10 13 1 9 1 9 2 13 15 9 2
18 16 13 2 15 13 9 2 15 13 9 2 7 13 1 15 13 9 2
4 13 15 13 2
2 15 2
5 11 11 2 9 11
5 9 11 1 0 9
16 9 1 9 13 9 2 7 1 9 1 0 11 11 13 3 3
2 9 9
14 9 0 0 9 1 9 11 11 13 0 9 0 9 2
19 3 15 1 11 13 9 1 9 7 13 9 1 15 13 3 1 0 9 2
6 11 11 2 11 1 11
21 1 0 9 1 0 9 0 9 2 15 1 9 12 13 0 9 2 13 3 13 2
34 0 9 9 7 15 3 13 1 11 11 2 12 2 14 1 15 2 16 9 0 11 13 9 7 0 7 0 9 1 9 13 1 9 2
22 1 9 12 1 15 0 9 1 9 12 1 11 3 13 13 9 3 2 16 13 3 2
33 1 12 9 0 0 9 0 9 13 3 16 9 11 11 2 15 15 1 9 12 13 1 9 0 9 16 0 9 1 9 9 9 2
27 3 1 11 1 9 9 9 3 13 11 3 1 0 9 0 11 12 2 12 7 1 9 9 13 7 9 2
5 0 11 15 13 2
40 0 9 1 9 13 12 9 1 11 2 11 7 11 2 7 16 1 0 13 9 10 9 14 0 9 2 13 4 3 11 0 13 1 15 1 9 1 0 9 2
5 0 9 13 0 2
22 9 13 12 2 9 7 9 0 9 13 13 1 0 11 1 12 2 2 12 2 12 2
6 2 13 4 13 9 2
17 14 2 1 9 15 13 13 2 2 13 11 11 1 9 1 11 2
38 1 0 0 9 1 11 12 2 12 15 15 13 2 2 13 4 15 13 2 13 9 7 15 3 13 1 0 9 7 13 15 2 2 13 1 0 9 2
35 2 1 11 15 13 1 9 10 9 2 2 13 15 13 9 9 11 11 2 12 1 9 0 11 2 15 13 1 0 9 1 0 0 9 2
17 2 9 1 12 0 9 13 0 2 9 1 12 9 13 3 0 2
14 9 15 1 9 4 13 13 10 0 9 1 0 9 2
10 2 1 9 1 15 13 0 9 9 2
20 1 9 13 0 9 11 12 2 12 2 0 9 0 9 11 11 12 2 12 2
29 3 15 12 13 9 9 0 11 7 0 9 15 13 0 11 11 7 9 1 11 4 13 0 9 16 0 0 9 2
2 11 11
3 9 11 9
1 9
3 0 11 2
4 11 1 11 2
5 11 2 11 2 2
27 9 0 0 9 11 11 15 13 15 2 16 4 0 13 1 10 0 9 11 2 15 13 1 0 0 9 2
20 9 9 1 15 13 9 11 11 2 10 9 7 3 1 0 9 11 3 13 2
11 2 9 13 1 11 9 0 2 7 0 2
13 13 13 0 9 2 7 9 13 3 1 0 9 2
25 1 9 9 15 9 13 2 3 13 11 12 0 9 1 0 7 0 0 9 2 2 13 11 11 2
3 9 1 11
5 11 2 11 2 2
17 0 9 9 11 11 15 3 13 11 9 2 10 9 13 11 11 2
33 9 13 1 11 1 9 12 2 12 2 1 10 9 3 1 11 11 7 11 11 13 1 9 11 11 7 9 13 1 12 2 9 2
7 3 13 12 9 1 11 2
8 9 1 11 13 1 12 9 2
5 13 7 9 9 11
6 1 9 13 9 9 2
4 9 1 9 2
7 9 9 11 2 11 2 2
22 9 1 11 4 1 9 13 0 0 9 9 2 15 15 3 13 14 1 9 0 9 2
15 0 9 15 13 3 12 0 9 2 16 15 4 13 12 2
18 2 3 15 13 2 16 3 13 11 7 11 2 1 15 4 3 13 2
19 1 0 9 3 13 11 7 1 9 9 11 2 2 13 9 9 11 11 2
27 11 7 11 13 14 9 3 2 3 9 9 1 12 9 3 13 1 9 2 16 9 4 0 13 0 9 2
17 13 4 7 7 0 9 2 11 2 11 2 11 7 0 0 9 2
37 13 3 0 9 2 0 7 0 9 1 9 1 11 2 11 7 11 2 0 1 11 2 11 2 13 15 0 9 11 11 11 2 2 11 7 11 2
32 9 11 11 11 3 3 13 9 10 9 2 15 15 13 13 0 0 9 2 3 1 9 9 13 0 9 11 2 11 2 11 2
32 1 9 13 2 11 11 2 11 11 2 12 11 11 2 2 11 11 2 11 11 2 11 11 7 11 11 2 15 11 11 2 2
14 9 1 9 9 13 11 11 2 11 0 7 11 9 2
13 0 9 1 9 12 11 9 13 13 1 9 9 2
13 0 9 9 13 0 2 16 3 2 13 12 9 2
15 0 9 13 11 2 3 9 13 9 1 9 12 9 9 2
12 9 13 12 9 7 1 9 13 3 0 9 2
19 11 9 2 3 13 9 12 2 9 3 2 13 13 9 1 12 9 9 2
6 11 3 13 1 9 9
9 1 9 9 0 9 15 13 0 9
2 9 9
2 11 2
34 9 0 9 9 1 9 9 9 12 11 11 2 15 1 9 3 13 1 9 1 11 2 15 13 1 9 3 1 9 11 1 0 11 2
20 11 11 11 2 15 13 0 9 2 4 13 1 11 1 0 9 1 9 9 2
21 9 1 9 0 9 13 4 1 10 0 9 13 1 9 1 9 0 9 1 11 2
16 11 3 3 13 9 2 0 0 9 2 15 13 9 0 9 2
36 15 9 11 11 2 15 0 9 13 0 0 9 2 0 9 1 9 1 3 2 1 0 9 1 10 0 9 11 11 13 1 9 9 0 9 2
25 9 2 11 11 13 1 9 1 11 9 0 9 2 15 4 13 13 9 1 9 0 9 0 9 2
6 10 9 3 13 13 2
32 3 12 9 2 11 11 7 11 11 2 13 0 2 0 9 2 3 0 9 0 1 9 9 12 7 0 15 9 1 10 9 2
17 9 12 9 15 4 13 7 0 9 11 1 10 0 9 1 11 2
33 9 11 11 11 15 3 13 9 2 16 4 9 0 9 1 9 9 12 2 1 15 15 0 9 13 2 13 9 0 9 1 11 2
12 13 3 9 2 16 4 9 1 11 13 0 2
10 7 15 13 1 9 0 9 0 9 2
17 3 15 13 2 16 11 13 1 0 12 9 0 9 0 0 9 2
30 3 7 2 16 9 1 11 11 2 1 15 15 13 12 2 9 0 0 9 2 13 13 1 3 0 7 7 3 0 2
17 13 13 2 16 4 10 9 1 9 0 9 11 13 1 11 13 2
18 11 11 3 13 1 9 10 9 9 2 16 13 1 0 9 0 9 2
8 3 13 15 0 9 10 11 2
29 7 16 0 9 11 11 2 15 13 3 13 1 9 1 9 2 15 3 13 1 9 2 10 9 13 7 3 0 2
8 9 9 12 7 7 9 13 2
14 9 11 11 3 13 9 1 9 2 15 13 11 11 2
22 10 9 4 15 13 13 0 11 11 11 2 1 15 11 13 14 1 0 9 0 9 2
5 0 9 13 11 2
11 11 15 1 12 9 13 1 0 9 0 9
2 9 9
4 11 9 2 11
32 12 9 13 3 14 1 9 7 0 9 1 9 9 11 1 11 9 9 0 0 9 11 7 13 15 13 0 9 0 0 9 2
8 3 15 13 1 12 2 13 2
63 1 12 1 12 1 12 13 9 11 11 7 10 9 11 11 2 16 0 9 13 9 11 1 9 12 2 15 13 2 16 0 9 1 11 1 9 12 2 13 2 0 0 9 11 2 7 9 9 11 11 2 16 0 9 13 12 2 9 12 13 11 2 2
35 3 14 1 12 0 13 1 9 11 2 9 11 11 7 10 9 11 11 2 10 9 13 9 1 9 1 9 9 1 12 2 9 12 2 2
9 13 9 13 3 13 0 9 0 2
13 1 0 9 13 1 0 9 13 0 9 12 9 2
45 0 9 0 11 13 3 1 9 1 9 2 11 0 1 11 11 11 2 7 3 1 9 1 9 2 11 11 11 2 7 13 9 3 1 0 9 2 7 7 1 9 9 10 9 2
14 9 3 13 1 9 2 0 9 0 9 1 0 9 2
32 7 1 0 0 9 0 9 13 0 1 9 13 3 9 1 15 2 15 13 0 9 2 13 2 1 0 0 9 1 9 12 2
29 1 15 3 13 9 2 1 15 15 9 1 3 0 9 13 13 1 9 0 9 11 0 9 0 9 11 11 11 2
15 1 15 9 11 9 11 11 2 2 9 13 1 15 11 2
13 11 13 10 0 9 7 1 0 9 15 3 13 2
16 0 13 1 15 9 11 2 15 13 2 16 9 13 11 2 2
28 3 10 9 1 9 11 9 2 11 11 13 1 9 1 0 9 0 13 2 16 10 9 13 1 9 11 11 2
4 9 0 2 11
2 11 2
8 11 2 11 2 2 2 12 2
7 9 9 2 11 0 9 2
2 11 2
2 11 2
3 0 9 2
2 11 2
11 9 9 2 15 13 9 1 11 2 4 13
22 1 9 1 9 1 11 4 13 9 9 9 11 2 15 13 9 1 11 2 11 11 2
12 1 0 9 13 11 0 16 9 9 12 9 2
18 9 13 13 1 9 2 16 9 1 11 13 1 9 12 9 0 9 2
26 0 9 3 1 9 0 9 13 10 9 2 7 0 9 11 13 2 16 9 13 0 9 9 1 9 2
17 1 0 9 14 13 11 1 9 1 3 0 0 9 7 1 9 2
24 1 9 15 13 7 0 9 9 11 11 1 11 2 2 13 2 16 9 1 11 4 3 13 2
12 9 9 12 13 0 16 0 9 1 11 2 2
1 9
3 11 11 2
3 0 11 2
3 11 3 13
5 11 2 11 2 2
27 9 11 15 1 0 9 1 9 1 11 2 12 2 12 2 13 1 0 9 0 9 1 0 9 1 9 2
33 0 9 9 13 9 11 1 9 11 2 15 13 3 1 0 9 0 9 7 1 0 9 1 9 1 11 4 10 9 1 9 13 2
20 1 9 11 13 3 0 9 9 12 0 9 2 15 13 12 9 1 0 9 2
16 1 0 9 1 9 9 0 9 9 0 9 3 13 0 9 2
16 1 9 1 0 9 1 0 9 13 7 0 13 0 0 9 2
12 1 9 13 9 7 13 2 3 9 7 9 2
16 0 9 12 7 12 9 2 0 0 12 7 12 9 2 9 2
13 1 9 13 9 2 3 14 3 2 3 3 9 2
15 0 9 12 7 12 9 2 2 0 12 7 12 9 11 2
20 1 9 13 9 1 12 7 13 1 12 2 9 13 1 12 7 13 1 12 2
26 0 9 12 2 9 2 0 9 12 9 2 12 1 9 12 2 0 9 12 9 2 12 1 9 12 2
9 0 0 9 13 12 9 2 9 2
16 0 9 1 0 9 1 9 13 3 3 0 2 1 9 0 2
3 2 11 2
13 9 2 0 9 0 1 0 11 1 9 4 13 2
8 9 1 9 13 13 0 9 2
11 4 13 0 9 12 7 12 9 2 9 2
21 9 1 11 11 2 0 9 1 0 9 9 1 11 10 13 9 1 0 0 9 2
17 2 3 13 1 11 2 3 15 1 9 13 1 11 10 0 9 2
15 13 7 3 1 9 2 16 1 9 4 13 14 12 9 2
23 7 7 4 13 13 0 13 9 1 0 9 1 11 2 12 9 2 9 2 9 2 2 2
12 1 0 12 9 15 13 0 9 1 0 11 2
29 9 9 15 1 11 13 9 0 9 7 1 9 2 16 13 3 1 9 11 11 2 13 11 1 9 1 0 9 2
22 16 15 15 13 13 15 1 9 7 9 2 13 1 0 9 1 11 13 1 0 9 2
22 1 0 9 15 15 1 9 13 0 9 11 2 15 13 3 10 9 2 2 2 9 2
2 11 9
2 11 2
13 1 9 9 14 1 0 9 13 12 2 9 9 2
24 0 9 13 11 11 9 2 15 1 0 9 13 12 9 1 9 2 12 2 9 7 0 9 2
14 1 9 15 13 1 9 0 0 9 11 11 1 11 2
12 1 0 9 4 13 9 11 11 7 11 11 2
3 9 1 9
7 12 9 0 9 11 2 11
2 9 9
5 11 2 11 2 2
30 9 0 0 9 11 2 11 2 12 2 12 2 1 9 13 14 1 12 2 9 7 1 15 13 3 9 1 0 9 2
27 0 9 4 1 9 13 0 9 9 11 7 11 9 2 1 9 9 3 13 9 11 1 9 0 9 11 2
39 2 9 2 16 1 9 13 9 2 13 4 0 0 9 2 2 13 9 11 11 2 2 1 9 0 13 3 0 2 7 15 4 1 15 13 13 9 2 2
22 0 9 13 1 12 2 9 2 3 0 11 13 0 9 7 13 1 15 0 0 9 2
15 12 1 0 9 13 1 9 7 9 15 1 10 9 13 2
18 3 1 0 9 0 9 13 11 0 9 2 16 0 13 9 1 9 2
11 2 13 0 9 2 0 15 13 1 9 2
11 0 9 2 0 2 2 13 15 9 11 2
8 9 11 1 0 9 3 13 2
21 1 0 9 13 7 1 0 9 11 2 15 13 1 9 2 15 14 13 3 9 2
11 9 3 1 9 13 9 9 3 1 11 2
31 0 9 13 9 9 7 9 3 1 9 7 1 10 0 9 4 13 9 0 9 9 11 7 11 2 15 3 9 13 2 2
12 2 16 13 1 9 2 3 13 1 9 9 2
11 13 4 0 2 16 4 3 13 10 9 2
21 1 9 13 9 9 11 2 15 12 9 7 9 2 2 13 15 9 0 9 11 2
6 9 11 13 11 9 9
7 11 2 11 2 11 2 2
15 12 0 9 9 1 0 9 1 9 1 12 2 9 13 2
28 11 13 11 2 12 2 12 2 2 11 13 12 9 1 11 2 12 2 12 2 1 9 13 1 0 9 2 2
22 12 9 3 13 9 11 2 12 2 12 2 2 15 13 9 1 11 1 12 2 9 2
11 0 9 1 9 3 13 9 1 9 11 2
19 2 1 15 2 16 13 0 9 10 9 2 13 15 0 16 9 1 9 2
55 1 9 13 3 2 9 15 3 3 13 2 7 7 15 13 13 9 0 9 2 15 15 13 1 9 1 9 1 0 9 2 2 13 9 9 11 11 7 13 3 9 2 16 0 13 7 2 16 4 9 9 2 13 2 2
13 2 13 4 3 13 9 1 9 2 7 13 15 2
11 11 3 13 3 2 7 7 13 14 13 2
15 13 13 2 16 3 13 2 2 13 11 0 9 9 11 2
29 0 9 11 15 13 2 16 1 9 9 4 13 1 11 13 10 9 2 16 9 9 2 1 9 1 9 1 9 2
21 11 13 9 11 1 12 2 9 2 7 9 11 15 3 13 1 0 9 10 9 2
23 11 13 1 9 12 2 12 1 11 0 9 11 2 10 9 1 0 9 3 13 0 11 2
20 11 13 13 0 9 2 16 4 3 13 11 2 7 9 9 11 13 0 9 2
12 9 12 2 9 9 2 12 2 12 2 12 2
12 13 13 11 2 11 2 7 11 2 11 2 2
8 13 0 9 1 0 0 9 2
21 9 10 9 1 9 15 1 0 13 1 0 11 3 0 7 13 13 10 0 9 2
11 0 9 13 1 11 7 3 13 9 0 2
5 3 3 1 11 2
11 1 11 13 9 0 2 7 9 15 13 2
8 11 13 3 3 1 9 1 2
18 13 7 0 9 2 16 16 15 0 13 1 2 13 15 13 7 11 2
10 13 10 9 1 9 10 9 1 9 2
20 13 3 13 1 15 2 16 10 0 9 9 13 0 9 1 0 9 1 9 2
9 14 15 2 3 15 9 0 13 2
11 16 10 0 9 4 3 1 9 9 13 2
12 13 15 2 16 9 1 9 13 1 9 13 2
14 15 1 10 9 2 7 0 9 3 2 13 0 9 2
19 13 15 7 2 16 9 13 13 13 1 10 9 1 0 9 1 9 12 2
8 9 1 9 13 1 11 9 2
9 16 10 9 13 2 13 9 0 2
19 4 10 9 13 3 1 0 9 2 7 7 2 13 2 1 9 0 9 2
7 13 15 13 1 0 9 2
5 13 15 3 9 2
11 7 3 3 13 1 9 2 7 1 9 2
13 13 15 1 9 9 9 1 9 2 11 2 0 2
6 0 0 9 13 0 2
14 15 15 13 15 0 1 11 7 0 9 3 3 13 2
7 15 3 13 7 1 11 2
10 16 13 1 11 13 0 9 1 11 2
11 2 0 9 15 13 1 9 1 11 2 2
22 11 13 2 16 15 2 15 15 13 2 13 3 1 9 1 9 9 9 9 1 11 2
20 1 0 9 1 9 2 11 2 1 11 4 13 0 9 7 13 15 15 13 2
22 1 9 9 0 0 7 0 9 15 13 13 3 1 0 9 1 9 1 0 9 9 2
26 9 0 7 0 0 9 2 0 7 0 2 2 9 2 9 9 7 9 13 1 9 1 12 2 9 2
3 2 11 2
9 9 2 9 2 9 2 9 11 11
27 1 0 0 9 13 9 2 16 0 2 0 2 0 9 7 9 2 16 7 9 7 9 2 13 0 9 2
42 1 11 2 1 11 7 1 11 10 9 9 7 0 9 0 7 0 9 3 9 1 0 9 13 0 3 15 2 16 15 1 9 13 1 9 1 9 2 15 13 9 2
38 16 4 1 11 13 0 9 2 3 15 3 3 13 2 16 9 2 15 13 1 11 7 3 3 2 3 13 1 9 2 13 0 9 3 1 0 9 2
17 0 15 13 1 9 2 15 13 9 13 1 9 1 9 0 9 2
12 9 13 3 0 9 9 2 3 0 7 0 2
66 15 9 2 9 2 9 2 3 9 0 12 9 2 15 13 1 9 2 16 4 15 1 15 15 13 2 16 4 15 15 13 2 7 16 4 15 1 9 2 11 7 11 13 10 9 2 7 13 15 2 16 4 15 9 2 11 7 11 13 9 13 7 0 9 9 2
11 7 3 3 1 9 1 9 0 0 9 2
33 9 9 1 9 9 0 2 11 15 1 9 9 13 1 9 0 9 2 16 15 1 0 7 3 1 0 9 13 2 3 16 9 2
12 0 10 9 1 9 9 0 2 11 13 0 2
28 15 0 15 13 7 9 0 9 2 15 13 9 2 7 0 9 2 15 15 13 3 13 16 2 9 9 2 2
144 16 4 9 9 1 0 11 2 3 1 11 14 1 11 13 10 9 0 2 3 7 0 9 0 9 2 9 7 9 2 16 13 0 2 11 2 13 9 1 9 13 15 9 0 11 1 11 1 11 2 1 9 12 2 12 9 1 0 2 11 1 11 9 9 2 9 1 11 2 3 1 9 12 4 13 12 0 9 2 16 4 15 13 13 0 11 2 0 0 2 11 2 9 0 2 11 1 11 2 9 0 11 1 11 2 9 1 11 2 9 1 11 2 10 11 1 11 3 2 3 2 2 3 4 15 13 1 9 2 1 15 0 9 13 9 0 9 1 9 7 9 0 9 2
6 9 1 11 13 9 2
19 1 12 9 9 11 4 13 12 9 2 1 15 2 14 2 1 12 13 2
30 1 9 9 4 1 12 9 2 1 15 13 3 12 9 9 2 13 12 9 2 2 13 9 0 9 1 0 9 11 2
22 2 1 0 9 13 0 9 0 9 2 15 13 13 0 9 2 1 15 15 9 13 2
12 13 15 0 9 2 9 1 0 9 2 9 2
17 9 1 11 13 0 9 2 9 2 0 9 2 2 13 9 11 2
11 0 9 1 9 1 11 13 13 0 9 2
25 9 9 9 9 9 1 9 2 15 13 9 1 11 9 1 9 2 13 1 0 9 12 2 12 2
25 3 1 11 2 9 13 3 1 9 2 13 11 11 9 1 0 9 1 11 11 1 9 1 0 12
7 9 11 2 1 9 0 9
4 11 11 2 11
23 3 12 0 9 13 3 3 1 9 0 9 1 11 9 1 9 9 0 15 9 0 9 2
31 9 9 0 9 13 3 0 1 15 2 16 4 11 2 11 2 11 7 11 13 1 9 0 9 13 1 0 2 9 2 2
20 1 9 2 15 10 9 13 1 0 9 3 2 9 10 9 13 3 0 9 2
18 2 13 2 16 15 0 9 13 1 0 9 2 0 15 7 13 13 2
17 9 9 0 9 2 15 13 1 9 9 2 15 13 13 1 9 2
29 1 10 9 15 13 2 16 9 4 13 3 0 9 2 2 13 15 1 15 3 1 11 0 9 9 11 11 11 2
45 1 9 9 11 11 13 0 9 0 9 9 9 1 9 15 2 16 12 1 0 9 2 0 9 0 9 1 0 9 2 9 9 1 9 13 7 13 9 1 10 9 1 12 9 2
20 9 7 13 3 0 9 1 15 2 16 4 9 9 1 9 9 2 13 2 2
29 9 0 9 0 9 11 3 13 10 0 9 7 7 12 13 0 9 1 9 1 9 2 1 15 4 0 9 13 2
26 10 9 13 3 13 9 2 16 4 15 1 10 9 13 1 9 0 9 1 9 3 3 2 13 2 2
5 2 9 1 11 13
2 11 2
27 9 9 0 9 2 9 2 3 13 9 9 9 2 16 4 13 0 9 7 0 12 0 9 9 0 9 2
26 9 9 2 0 9 10 0 0 9 1 9 1 0 9 2 4 1 9 0 9 13 1 9 1 11 2
23 11 2 11 2 11 2 11 2 11 2 11 7 12 0 9 13 3 1 9 14 9 9 2
15 0 9 9 0 7 0 11 1 11 13 3 11 7 11 2
4 11 13 9 9
2 11 2
20 0 9 3 13 9 0 9 2 15 13 13 11 9 11 9 1 9 1 11 2
20 9 3 13 9 9 9 0 9 2 16 15 1 9 9 13 9 9 12 9 2
20 13 13 3 9 9 1 9 2 15 13 9 9 0 9 7 9 1 0 9 2
7 9 9 3 13 9 9 2
33 9 9 7 9 1 0 9 13 1 0 9 9 0 0 9 7 13 7 12 1 9 2 1 15 15 11 13 1 9 1 9 11 2
17 0 9 1 9 7 9 2 0 1 0 9 2 10 9 3 13 2
36 1 9 9 11 11 4 13 9 9 13 10 0 9 7 9 3 2 16 13 15 0 1 10 0 9 2 3 0 9 1 9 1 9 2 9 2
3 13 9 9
9 9 0 9 1 11 11 11 1 11
2 9 9
4 11 11 11 11
24 1 9 1 9 9 0 9 1 9 0 9 13 3 1 11 10 9 9 0 0 9 11 11 2
8 13 9 1 9 1 0 9 2
9 10 9 13 1 0 9 0 9 2
18 13 7 13 9 1 11 2 10 0 9 13 1 9 1 11 0 9 2
11 3 3 13 0 9 1 9 0 0 9 2
15 9 11 11 15 13 3 1 9 1 9 1 0 0 9 2
16 1 9 2 3 15 13 2 13 2 2 13 1 15 12 9 2
12 13 15 2 16 13 10 0 9 1 10 9 2
15 1 0 9 15 13 2 16 4 15 11 13 13 0 9 2
19 9 4 15 3 13 7 13 4 15 0 7 1 11 2 7 1 11 2 2
4 9 1 9 12
11 3 1 9 3 0 9 2 9 9 11 11
2 0 12
2 9 12
10 3 2 16 4 15 1 9 9 13 2
5 3 7 15 13 2
3 9 11 11
5 0 9 13 9 11
4 11 11 2 11
24 1 0 9 13 3 3 1 11 9 0 9 0 9 9 9 1 9 0 9 1 0 12 9 2
14 1 9 9 13 13 3 12 9 9 1 0 9 12 2
12 3 3 15 13 9 2 15 13 1 9 9 2
35 1 9 0 2 9 2 4 3 1 10 9 15 13 1 15 2 16 4 15 1 9 0 9 13 11 2 11 2 11 7 11 10 0 9 2
20 3 3 13 14 15 2 16 4 9 1 9 13 3 9 0 9 1 0 9 2
13 11 1 15 4 13 9 16 0 2 3 1 9 2
11 0 9 13 0 2 15 13 0 0 9 2
13 1 10 0 9 15 3 9 13 14 1 0 9 2
17 3 3 13 3 0 2 16 9 1 0 9 15 1 10 9 13 2
31 3 7 15 3 9 9 13 13 9 2 16 4 3 0 9 1 9 0 9 1 9 4 13 14 1 0 9 9 1 9 2
11 9 1 9 9 4 3 13 3 0 9 2
4 9 1 0 9
30 2 16 13 9 0 9 1 9 3 2 13 15 1 9 9 2 2 13 3 3 9 0 2 0 9 11 2 11 11 2
45 9 3 13 9 2 16 13 1 9 2 16 16 4 9 4 1 12 2 9 13 2 13 4 1 0 9 0 2 16 4 15 11 2 11 2 11 7 11 13 1 9 1 0 9 2
15 0 9 4 15 3 1 9 10 9 13 3 16 1 9 2
8 11 13 1 9 9 11 7 11
2 11 2
42 0 9 11 11 3 13 2 16 0 9 11 11 13 1 0 7 0 9 2 15 4 13 11 13 15 1 9 9 1 0 9 1 9 11 7 1 11 1 0 9 11 2
38 2 13 9 1 3 0 9 9 0 0 9 2 7 3 15 13 2 16 9 9 1 9 11 13 3 12 7 12 9 2 7 11 1 15 3 13 13 2
15 3 15 13 2 2 13 11 1 9 9 1 0 0 9 2
16 10 9 7 0 9 15 13 2 16 10 9 9 1 15 13 2
18 13 3 0 9 9 2 15 13 10 9 2 7 0 9 0 0 9 2
10 9 11 9 9 13 9 3 9 9 2
7 13 15 1 10 10 9 2
2 14 2
10 13 15 3 2 0 9 13 1 15 2
17 0 9 9 0 9 11 13 0 0 9 1 9 0 1 0 9 2
7 7 3 15 1 15 13 2
26 1 11 4 15 13 1 0 9 7 13 4 2 16 9 9 13 1 15 2 15 13 13 1 0 9 2
5 13 4 9 9 2
19 9 11 7 9 13 9 1 15 2 16 4 15 13 2 15 13 1 0 2
8 7 15 13 7 9 0 9 2
23 9 0 9 11 11 2 11 13 2 16 13 2 3 13 13 9 11 7 3 9 0 9 2
16 3 15 13 13 3 1 12 9 2 16 15 9 1 9 13 2
18 7 10 9 13 13 3 1 12 1 10 9 9 2 15 4 3 13 2
3 3 9 2
9 1 11 7 0 0 9 7 13 2
18 10 9 2 3 2 9 11 7 9 11 2 7 7 0 2 15 13 2
20 11 1 15 14 13 9 10 0 9 7 13 15 3 2 13 3 9 9 11 2
13 13 2 16 0 2 0 9 1 9 10 9 13 2
13 1 15 3 1 15 13 9 9 1 9 9 11 2
18 10 9 13 13 2 16 9 13 1 15 0 16 1 12 1 9 9 2
13 3 11 13 3 14 15 2 15 15 13 9 9 2
33 9 13 1 15 2 16 9 9 3 13 3 4 13 10 9 2 16 9 15 13 1 9 7 10 9 15 13 2 16 3 15 13 2
10 7 1 11 3 10 9 13 9 3 2
16 3 13 3 0 9 2 11 15 13 9 1 0 9 2 3 2
11 7 16 11 13 14 2 9 1 15 13 2
9 13 3 13 1 0 9 3 13 2
19 0 13 2 7 9 13 2 16 1 9 9 1 10 9 15 13 3 13 2
10 16 13 7 9 3 11 2 3 13 2
23 13 4 7 2 16 15 1 9 13 9 7 9 2 15 15 3 13 1 3 3 0 9 2
12 15 3 13 2 16 9 13 0 9 9 9 2
5 11 2 11 2 2
23 9 9 3 13 12 0 0 9 1 0 9 12 9 7 3 13 13 0 9 1 0 11 2
24 1 9 9 2 0 13 0 12 9 2 9 13 1 15 1 12 0 0 9 1 9 12 9 2
25 1 9 11 13 2 16 1 9 12 13 9 9 1 9 1 11 1 9 12 1 3 16 9 9 2
6 9 13 9 1 11 2
18 9 2 15 3 11 13 0 9 2 13 2 16 0 9 4 3 13 2
7 9 13 3 9 1 11 2
22 0 9 13 9 2 3 1 11 13 0 9 0 9 3 2 16 1 9 13 15 9 2
19 0 9 2 15 13 1 9 2 15 13 9 2 0 9 7 9 1 11 2
20 1 9 9 15 9 9 13 1 0 9 1 0 11 1 11 7 13 10 9 2
20 3 15 13 1 9 1 3 0 9 2 15 1 9 1 9 13 3 0 9 2
10 15 7 13 1 11 9 1 9 9 2
3 9 12 2
21 16 1 9 12 13 1 11 1 9 9 12 9 1 11 2 3 15 13 3 12 2
5 9 11 11 2 11
15 10 9 1 10 0 9 3 2 13 2 1 9 9 11 2
26 9 1 9 7 9 0 9 1 9 1 12 2 9 12 13 0 0 9 1 0 9 0 11 7 11 2
20 1 0 9 7 11 3 1 11 13 12 9 2 3 13 9 11 13 0 9 2
5 12 9 1 0 9
2 11 2
12 3 1 9 4 13 11 11 13 13 0 9 2
23 15 1 15 13 1 15 2 3 15 0 0 9 13 9 2 0 13 9 0 16 12 9 2
21 15 9 15 1 11 13 1 0 9 1 0 0 9 2 0 0 9 7 0 9 2
18 11 2 11 2 15 14 3 13 0 9 2 13 3 13 1 12 9 2
8 15 13 13 7 0 9 0 2
18 9 4 13 9 2 9 11 2 7 13 15 13 11 2 0 0 9 2
11 9 11 13 1 9 9 3 1 0 9 2
6 9 13 1 9 12 2
5 9 9 15 4 13
5 11 2 11 2 2
30 9 9 1 9 15 3 13 1 12 5 1 9 1 12 5 1 9 2 15 13 1 9 1 9 1 12 9 3 9 2
15 9 9 13 1 9 9 7 7 1 15 3 13 0 9 2
34 1 9 11 11 1 0 9 9 7 9 13 0 2 16 0 9 13 13 0 9 3 13 2 16 15 13 12 1 0 9 2 3 9 2
11 0 9 0 9 13 2 16 9 15 13 2
17 3 15 9 13 1 12 2 7 12 2 9 2 9 7 3 13 2
17 9 13 1 9 2 11 0 7 0 0 9 13 2 13 15 9 2
14 14 3 7 1 11 13 0 9 0 9 1 9 9 2
28 1 10 9 13 0 9 11 2 11 12 9 2 7 15 9 0 9 2 15 3 1 10 9 16 1 0 13 2
9 0 9 13 13 1 9 1 0 9
4 11 2 11 2
14 1 12 9 10 9 13 1 3 2 0 7 0 9 2
33 1 9 0 9 1 9 1 12 1 12 9 1 9 9 12 7 12 15 13 1 9 9 9 1 12 9 3 16 1 0 0 9 2
14 1 11 15 1 0 9 9 10 9 1 12 9 13 2
31 12 1 12 9 10 9 13 13 0 2 0 9 2 13 0 2 13 0 0 9 2 4 1 15 13 9 7 0 9 9 2
37 13 15 3 9 1 0 9 11 11 1 12 2 0 9 11 1 9 1 9 11 2 15 13 1 12 2 1 12 2 9 1 9 1 9 1 11 2
14 1 9 13 3 1 12 9 0 13 0 9 0 9 2
31 1 9 11 4 13 9 0 9 2 0 9 2 0 9 2 3 0 9 7 0 9 2 15 13 1 0 9 9 3 13 2
21 9 2 15 13 13 7 1 9 2 15 13 3 16 12 9 7 9 3 1 11 2
19 13 3 7 0 9 2 15 13 9 3 1 9 9 9 7 9 0 9 2
5 11 2 11 2 2
24 13 9 0 7 0 9 1 0 9 0 13 3 1 0 9 9 9 11 2 11 2 11 2 2
15 2 13 15 9 2 15 15 15 13 2 2 13 10 9 2
22 1 9 1 9 9 1 0 9 11 3 13 13 0 9 1 9 1 9 11 2 11 2
28 13 1 9 0 9 9 0 9 1 11 2 11 2 11 7 0 9 3 9 9 11 2 11 2 11 2 13 2
31 2 13 9 7 1 11 2 0 9 7 3 13 13 2 2 13 0 9 0 9 1 9 0 9 11 2 11 2 11 2 2
20 9 3 13 2 16 13 0 2 16 4 0 9 13 9 10 9 1 9 9 2
18 1 11 2 11 2 11 2 4 10 9 13 4 13 16 0 9 9 2
9 7 0 9 9 3 13 2 13 2
23 0 9 0 9 7 11 13 4 13 1 0 0 2 0 9 2 15 1 9 13 10 9 2
6 11 11 1 9 13 4
5 11 2 11 2 2
11 0 0 9 13 0 9 1 9 0 9 2
14 16 15 4 1 10 9 13 2 13 1 9 0 9 2
15 1 10 9 7 9 13 11 11 2 3 15 1 9 13 2
8 9 0 9 3 11 13 13 2
23 1 9 11 11 15 9 3 13 13 0 9 2 15 15 13 9 1 11 7 1 0 9 2
25 3 2 3 15 15 13 2 15 13 1 0 9 0 2 1 15 13 3 13 3 9 7 0 9 2
16 16 15 0 9 13 1 9 1 0 9 2 9 4 15 13 2
37 11 13 3 3 9 9 2 0 9 1 9 11 13 0 13 2 2 3 2 1 11 11 2 0 11 2 0 11 2 11 7 1 12 0 9 11 2
13 3 1 9 16 1 0 9 13 1 12 9 9 2
17 9 9 13 1 0 9 11 3 13 2 3 14 7 1 0 9 2
16 13 15 15 0 9 1 9 9 7 9 9 1 9 0 9 2
17 9 9 1 0 9 11 13 3 3 2 16 4 13 13 10 9 2
10 9 1 9 0 9 0 9 1 9 2
5 11 2 11 2 2
19 9 4 13 13 9 13 1 9 0 9 1 9 7 9 9 7 9 9 2
20 10 9 9 1 9 13 3 12 9 1 9 1 10 9 0 1 9 0 9 2
15 9 7 3 13 0 13 9 2 15 4 13 9 1 9 2
17 10 9 3 1 9 0 9 13 9 11 11 2 11 2 1 9 2
21 9 9 13 13 9 2 1 15 4 15 9 13 9 9 13 1 9 0 9 3 2
10 0 9 4 13 9 13 1 0 9 2
25 1 9 13 9 7 9 9 0 13 9 2 16 9 15 10 9 1 12 9 13 9 0 0 9 2
5 15 13 12 9 2
4 0 9 13 3
2 11 2
29 9 15 12 9 2 15 13 0 9 2 15 1 0 0 9 9 7 0 9 13 1 9 10 9 7 9 1 9 2
11 1 9 11 13 10 9 3 13 10 9 2
13 1 0 0 9 15 13 9 0 9 11 11 11 2
23 0 9 13 11 2 11 2 0 9 2 9 0 2 0 9 2 9 9 7 0 9 9 2
18 1 11 4 9 3 2 13 0 9 9 7 13 15 1 10 9 2 2
12 13 15 3 0 7 0 9 2 9 7 9 2
5 11 13 9 1 11
2 11 2
20 13 9 2 16 4 13 9 1 9 9 1 0 0 9 11 2 4 9 11 2
19 1 0 0 9 11 15 13 10 9 11 11 2 15 13 3 9 0 9 2
16 9 11 1 15 13 1 0 9 1 9 9 7 0 0 9 2
16 13 2 16 11 7 11 13 9 2 7 11 9 13 12 9 2
10 7 3 13 0 9 0 1 0 9 2
18 9 0 0 9 11 11 13 1 9 11 2 13 2 14 9 1 9 2
2 13 2
14 11 4 13 1 9 13 2 13 15 9 9 1 9 2
7 13 15 1 10 0 9 2
2 13 2
16 13 0 9 7 0 9 1 0 11 2 11 2 11 2 11 2
11 13 15 11 13 2 16 4 13 0 9 2
9 9 1 11 13 1 9 9 0 2
6 1 0 11 13 9 2
13 3 2 12 9 1 9 2 3 13 13 0 9 2
8 13 9 9 0 9 1 11 2
18 14 2 7 13 15 2 16 3 13 10 9 2 3 1 11 2 13 2
13 7 9 15 4 13 13 3 2 16 4 13 9 2
18 1 9 1 0 9 15 13 1 15 2 16 4 9 13 13 11 13 2
13 9 1 15 3 13 2 7 14 3 15 3 13 2
9 13 15 3 13 0 9 0 9 2
4 15 13 9 2
18 1 0 9 15 15 13 2 1 12 2 1 15 12 13 1 0 11 2
6 3 1 12 12 9 2
7 13 9 2 16 9 13 2
7 3 13 2 7 13 0 2
14 1 9 12 13 1 10 9 0 2 3 10 9 13 2
8 9 1 11 11 2 0 0 9
24 3 1 9 9 13 1 15 2 16 12 1 0 9 0 9 13 9 9 1 0 9 7 9 2
7 13 3 13 10 0 9 2
17 15 13 3 1 0 9 2 13 15 3 0 9 2 9 1 9 2
19 9 13 0 7 1 10 9 3 13 9 0 0 9 7 13 1 10 9 2
24 0 9 13 1 10 9 0 0 9 7 9 2 16 0 9 9 13 1 15 9 9 7 9 2
3 2 11 2
8 0 9 1 0 9 1 0 9
5 11 2 11 2 2
17 1 9 9 9 13 3 9 1 9 0 0 9 9 2 11 11 2
28 9 11 11 13 9 2 16 10 9 4 1 0 9 13 7 16 15 3 1 0 9 10 0 9 13 0 9 2
23 3 3 9 13 9 9 9 1 9 9 7 9 7 1 10 9 2 15 13 9 0 9 2
25 9 1 9 13 2 16 13 13 1 3 0 9 7 16 9 9 1 15 0 13 3 0 0 9 2
13 9 3 13 7 9 9 9 7 9 1 9 12 2
20 1 2 0 9 0 9 2 13 1 11 2 0 9 2 3 1 10 0 9 2
17 3 9 13 9 11 9 9 9 9 2 1 15 9 4 9 13 2
14 9 3 13 1 0 9 0 9 11 1 9 0 9 2
18 9 13 1 12 2 9 13 9 2 1 15 13 0 9 1 0 9 2
23 11 11 3 13 9 9 9 0 9 7 9 0 9 0 9 2 0 15 9 9 0 9 2
20 2 13 4 0 2 16 4 15 15 13 13 9 0 0 9 2 2 13 9 2
11 9 0 9 9 9 13 0 9 11 11 2
37 0 0 9 10 9 13 13 13 11 3 3 16 0 0 9 2 7 2 3 3 2 16 0 9 2 15 1 0 9 1 0 9 13 13 7 9 2
12 9 11 2 13 11 2 13 0 13 1 9 2
25 15 2 16 13 1 9 9 11 2 13 1 15 2 15 15 15 13 3 3 13 2 13 0 9 2
27 13 1 0 9 7 13 11 2 16 4 15 13 9 15 2 15 13 2 4 3 11 13 3 3 1 9 2
10 14 4 15 3 13 0 9 0 9 2
19 11 15 3 13 13 0 9 2 15 3 2 3 3 3 2 13 1 11 2
23 0 9 0 9 11 1 11 3 13 2 16 1 9 0 9 13 16 0 13 0 9 0 2
6 15 1 10 9 13 2
10 3 0 9 0 15 1 9 1 11 2
14 10 9 2 1 0 9 1 9 0 9 2 3 13 2
3 11 13 9
6 11 2 11 2 11 2
24 0 0 9 2 11 2 3 13 2 16 13 10 9 1 0 9 9 9 1 9 0 2 11 2
26 11 11 13 9 9 11 2 16 13 9 1 9 0 2 11 2 3 12 9 13 1 9 1 0 9 2
22 9 13 1 9 1 9 13 0 9 9 2 3 3 2 16 4 13 3 13 1 9 2
5 9 13 3 3 2
29 1 9 0 9 2 15 15 13 4 13 2 13 9 11 1 9 11 11 0 9 1 9 1 0 9 0 0 9 2
47 0 9 1 9 3 16 12 9 15 9 13 2 16 11 1 0 9 13 3 0 12 9 9 2 16 0 11 13 12 9 7 1 9 0 0 9 2 11 2 11 11 2 1 11 12 9 2
13 2 0 9 13 1 9 0 9 7 9 0 9 2
19 1 0 4 13 3 0 9 0 1 9 12 2 15 13 3 9 0 9 2
37 3 2 1 9 9 1 9 1 9 2 13 9 2 16 4 0 9 13 13 1 0 0 9 2 2 13 3 1 0 9 1 11 0 9 11 11 2
12 0 9 11 11 13 3 13 9 11 0 9 2
28 1 9 1 0 9 0 9 11 11 1 11 11 13 2 16 4 13 13 3 1 12 9 9 1 0 12 9 2
5 0 9 14 13 9
2 11 2
23 0 0 9 3 13 2 16 1 9 0 9 0 1 9 1 0 9 0 1 9 13 9 2
15 9 0 0 11 13 10 9 1 15 2 15 10 9 13 2
8 13 14 2 16 13 0 9 2
12 15 4 3 1 9 13 7 15 13 1 9 2
12 1 9 2 16 13 1 11 2 13 9 13 2
13 0 9 3 1 9 13 2 16 0 9 13 11 2
7 0 0 9 13 0 9 2
33 0 9 3 13 9 11 11 2 16 13 1 9 13 9 2 7 13 9 1 15 2 16 4 15 1 9 0 0 9 13 0 13 2
8 9 15 13 2 3 2 2 2
37 9 1 9 9 9 2 1 12 9 2 13 13 9 12 9 1 0 11 2 15 15 0 9 13 0 9 13 9 1 0 9 1 9 12 1 15 2
19 3 3 13 0 9 2 9 13 3 1 9 1 9 13 0 9 0 9 2
17 9 13 1 9 7 13 9 1 9 2 3 15 0 9 9 13 2
19 1 9 2 16 9 13 9 2 7 9 3 13 1 9 9 3 1 9 2
18 9 2 1 15 13 14 9 2 7 7 9 2 16 0 9 13 3 2
4 11 13 0 9
2 11 2
24 13 1 9 1 0 9 13 0 9 11 11 1 9 2 16 15 1 9 10 9 13 0 9 2
24 2 13 2 16 1 10 9 4 13 3 15 0 9 2 2 13 9 1 0 9 1 9 11 2
18 11 13 2 16 13 0 9 2 16 12 1 9 9 13 9 1 9 2
10 2 3 15 13 13 9 2 2 13 2
16 13 3 2 16 1 9 13 14 12 7 12 9 1 9 9 2
5 0 9 1 9 9
23 11 13 2 16 0 11 13 9 2 0 9 2 1 9 2 16 15 13 13 9 1 9 2
18 0 11 0 9 13 2 16 15 3 13 1 0 9 1 9 1 11 2
36 0 9 9 0 0 9 13 1 9 1 9 0 9 1 9 9 1 0 9 1 9 9 2 15 13 1 9 9 9 9 1 9 9 9 9 2
13 9 9 11 11 13 2 16 1 10 9 15 13 2
29 0 9 11 11 3 1 0 9 11 13 0 0 9 2 15 15 0 0 9 16 0 9 13 1 9 9 1 9 2
23 11 3 13 3 15 0 9 11 2 12 2 15 1 9 12 9 13 1 9 0 0 9 2
12 13 15 1 11 9 0 9 9 9 11 11 2
15 0 9 4 13 11 3 7 3 16 0 0 9 11 11 2
29 13 15 1 10 0 9 2 9 9 2 0 0 9 0 9 11 11 2 15 3 11 1 9 12 13 1 0 9 2
20 3 9 9 0 0 15 3 13 0 9 1 9 1 0 9 0 9 0 9 2
8 13 15 9 0 0 9 11 2
38 9 1 0 9 2 15 1 9 12 13 9 0 9 1 0 9 2 11 2 2 13 0 9 11 1 9 0 9 1 11 1 12 2 1 12 2 9 2
18 1 9 11 2 15 4 13 1 11 2 13 9 0 9 9 0 9 2
42 0 9 11 11 2 15 4 1 9 13 1 11 7 3 13 11 2 13 2 3 2 3 1 0 9 7 13 1 0 9 2 15 15 7 3 4 13 14 1 10 9 2
13 11 15 13 9 1 0 9 2 15 15 9 13 2
52 0 9 4 3 13 0 9 0 0 0 0 0 9 2 11 2 1 9 1 0 9 0 9 1 9 1 11 2 1 15 15 13 0 9 2 7 1 9 1 9 0 9 2 15 13 0 9 9 11 11 11 2
13 1 0 9 1 0 2 0 11 4 13 10 9 2
20 3 3 13 9 2 4 12 9 1 9 1 9 13 0 9 7 9 0 13 2
11 12 3 12 9 0 0 9 9 3 13 2
39 0 11 11 11 2 15 4 1 9 1 9 13 0 9 1 12 9 9 2 4 13 9 2 1 9 9 0 9 11 11 11 4 13 3 13 14 12 9 2
9 9 2 15 13 9 2 3 1 9
23 9 2 15 4 1 9 1 9 1 9 1 12 9 1 11 13 2 4 3 13 1 9 2
24 14 0 2 12 9 0 9 4 3 1 10 0 9 1 0 9 1 11 13 1 0 0 9 2
9 10 9 1 9 13 9 1 9 2
15 9 2 15 9 13 2 13 1 9 1 9 13 1 9 2
9 0 9 9 13 7 13 1 9 2
13 0 9 7 13 2 16 1 9 13 1 0 9 2
22 0 9 11 15 1 11 1 0 9 13 1 0 9 9 2 15 4 1 0 9 13 2
15 1 9 13 1 0 9 14 12 3 0 9 7 10 9 2
28 0 9 7 1 10 9 13 7 9 15 13 2 16 13 12 1 3 9 2 15 15 13 9 1 11 1 11 2
3 2 11 2
4 9 11 13 0
7 11 13 1 9 11 1 9
2 9 9
5 3 0 0 9 2
18 1 11 15 9 1 9 13 0 9 2 1 15 4 15 13 0 9 2
17 9 7 3 13 7 0 9 13 0 9 7 1 10 9 1 9 2
24 1 9 15 9 13 9 7 10 9 3 13 0 9 2 16 13 0 9 0 13 1 0 9 2
10 3 1 9 2 14 1 11 2 2 2
4 11 9 9 13
2 9 9
4 11 11 2 11
17 9 0 9 13 10 0 9 2 15 13 9 0 9 1 0 9 2
34 0 0 9 13 0 9 11 9 1 9 11 1 9 11 2 0 9 12 0 9 2 15 3 4 1 12 9 13 7 3 13 1 11 2
46 13 0 12 9 9 2 16 13 0 13 9 2 3 13 9 1 9 2 2 9 0 7 0 9 7 9 1 9 2 0 1 9 0 2 9 0 9 2 12 2 12 2 1 11 2 2
9 0 2 7 10 0 9 0 9 2
28 13 3 2 16 0 0 0 9 13 13 9 11 1 9 2 10 9 9 2 7 13 9 0 9 1 0 9 2
15 1 0 9 11 2 1 11 2 3 0 9 13 9 11 2
27 13 15 9 9 1 9 10 9 7 3 13 1 15 2 15 3 13 9 13 2 16 0 9 13 0 9 2
24 10 9 13 11 0 9 2 0 9 2 2 15 13 9 2 0 9 2 9 11 1 11 11 2
19 9 0 0 9 1 11 13 0 9 0 9 7 9 10 9 1 0 9 2
9 13 9 2 15 3 13 0 13 2
19 9 0 9 7 9 9 1 9 9 1 0 9 7 9 15 13 0 9 2
13 13 15 7 13 14 3 2 16 15 13 0 9 2
16 1 0 9 15 13 1 10 9 1 9 0 0 7 0 9 2
13 1 9 0 0 9 15 3 13 9 13 11 9 2
44 11 11 2 10 0 11 13 3 1 0 0 9 2 7 3 10 0 9 11 11 13 1 9 10 9 0 9 2 3 0 9 0 9 11 2 16 9 1 9 7 9 13 0 2
26 9 0 9 11 1 9 1 0 9 13 0 3 0 9 0 1 11 1 9 9 1 9 1 0 9 2
12 3 13 2 16 0 11 13 13 0 16 0 2
25 1 11 15 7 9 3 2 13 2 9 11 7 10 2 0 9 2 13 16 9 1 9 0 9 2
28 9 1 2 9 2 1 0 9 2 15 15 13 3 1 11 2 13 1 9 2 15 1 0 9 13 1 11 2
26 1 9 1 0 9 1 11 11 15 3 16 12 5 0 11 13 2 16 0 9 10 9 13 1 0 2
20 11 15 13 1 9 1 9 1 9 2 15 13 1 12 9 1 9 0 9 2
12 9 1 0 9 1 9 9 9 13 0 9 2
26 11 11 2 0 9 0 0 9 7 9 0 9 2 0 9 2 2 0 1 0 9 2 13 0 9 2
21 9 2 13 2 9 13 1 9 0 9 16 9 7 9 1 9 2 9 1 9 2
41 0 11 2 13 3 9 0 11 2 15 3 13 3 1 9 2 3 1 9 2 7 15 1 0 9 2 13 9 7 9 1 9 7 13 15 9 1 9 7 9 2
18 7 10 9 15 1 0 9 13 13 1 11 1 9 7 1 9 0 2
19 1 0 9 4 11 13 10 0 9 7 13 4 15 0 1 9 0 9 2
19 0 11 13 1 9 2 15 13 9 1 9 0 7 0 9 2 3 0 2
37 3 0 7 0 9 7 9 0 0 9 2 15 13 13 0 9 0 9 7 15 13 9 1 10 0 9 2 15 1 0 0 9 13 16 0 9 2
42 0 9 1 11 7 9 0 0 9 1 0 9 1 9 2 1 0 9 9 1 0 1 0 9 2 3 13 2 16 9 0 9 7 9 9 13 1 11 1 9 9 2
10 0 0 9 0 9 9 0 9 0 11
12 11 2 0 7 11 2 12 2 12 2 12 2
13 1 10 9 4 13 3 9 9 0 9 1 9 2
15 13 15 15 9 11 2 11 2 11 7 3 15 15 13 2
27 9 13 1 11 11 1 11 2 11 2 11 2 15 15 13 1 2 12 9 2 2 7 3 15 13 9 2
8 1 15 15 3 13 9 11 2
7 9 13 3 1 10 9 2
28 7 16 15 15 13 2 3 9 10 9 15 13 9 9 2 7 3 9 2 15 11 13 7 13 1 10 9 2
4 11 11 2 11
3 14 1 9
5 6 2 9 11 2
28 13 4 3 0 9 9 2 11 12 2 12 2 12 2 2 15 3 13 9 2 13 0 9 1 9 7 9 2
14 3 13 13 0 2 16 10 9 9 1 0 13 0 2
21 13 15 13 9 1 10 9 1 9 1 10 2 3 13 0 2 0 2 9 0 2
32 1 0 9 0 2 3 4 13 9 1 9 13 2 16 4 13 10 0 9 2 13 4 1 15 10 9 2 16 15 9 13 2
44 0 9 2 0 9 1 9 2 12 2 4 13 9 2 16 13 14 1 9 9 2 15 13 9 9 3 1 0 0 9 7 1 0 9 2 7 13 14 3 1 9 0 9 2
29 3 9 9 2 9 2 0 9 2 9 2 0 9 7 0 9 13 1 11 2 0 13 12 2 7 12 2 9 2
21 9 7 9 15 3 13 12 2 12 9 1 9 1 11 7 0 12 9 1 11 2
12 9 2 9 7 9 13 13 12 9 1 9 2
14 3 15 7 9 11 7 9 13 1 12 9 1 9 2
48 13 0 12 9 2 13 15 1 0 9 0 2 0 2 9 1 9 0 7 1 0 9 2 7 1 0 9 11 13 0 9 1 0 9 1 0 9 2 1 0 9 7 9 1 9 7 9 2
20 4 13 2 16 1 0 9 13 0 9 1 0 9 2 16 0 9 3 13 2
8 0 15 13 7 1 0 9 2
26 0 0 9 13 0 7 1 0 9 11 2 3 9 9 13 0 9 1 9 9 7 13 0 9 9 2
11 7 1 9 0 0 9 13 0 13 9 2
16 13 14 9 1 0 9 2 13 4 13 9 1 0 9 9 2
20 7 13 0 13 0 9 1 9 9 1 9 7 1 0 9 9 1 0 9 2
17 0 9 4 13 1 9 1 9 13 1 11 7 3 13 0 9 2
16 0 0 9 1 9 0 9 1 0 9 13 3 0 9 9 2
15 1 9 13 9 10 0 9 7 9 0 9 1 0 9 2
1 9
11 1 11 13 12 0 0 9 7 12 9 2
18 14 1 0 9 11 13 3 16 12 9 2 1 0 9 1 12 3 2
7 13 9 2 16 13 9 2
4 9 0 9 13
2 11 2
9 0 9 13 3 1 10 0 9 2
18 1 0 9 0 9 13 0 0 9 1 0 9 0 9 1 12 9 2
17 1 0 9 9 13 9 0 9 1 0 9 0 9 1 12 9 2
21 0 9 15 13 1 12 9 2 16 9 13 13 1 3 16 12 12 15 0 9 2
7 9 9 13 1 12 9 2
11 3 13 13 9 9 2 0 7 0 9 2
12 0 9 13 3 1 0 9 2 9 7 9 2
9 0 0 0 9 1 9 1 0 9
5 11 2 11 2 2
26 0 7 0 9 13 9 9 7 9 2 9 2 1 9 10 0 9 9 2 15 15 13 10 0 9 2
14 1 9 1 9 13 1 10 9 13 1 0 0 9 2
26 9 3 13 9 9 9 1 0 9 2 13 9 2 9 7 13 9 0 9 1 9 1 15 0 9 2
23 3 13 3 3 9 0 9 1 9 1 0 9 7 9 3 0 2 3 15 9 3 13 2
16 14 1 11 3 3 13 0 9 1 9 9 1 12 0 9 2
12 9 13 1 10 9 14 12 9 2 9 3 2
41 0 0 0 0 0 9 13 9 12 0 9 2 9 7 9 1 9 11 2 0 7 0 0 0 7 0 11 2 1 11 2 15 15 13 12 2 2 12 2 9 2
20 13 1 0 9 2 3 15 13 9 9 1 12 9 2 3 0 7 0 11 2
8 3 16 9 9 13 1 11 2
8 1 11 13 1 11 12 9 2
15 9 1 9 13 0 9 0 9 7 13 1 9 0 9 2
20 1 0 9 13 7 12 9 2 0 7 11 2 0 9 0 9 7 11 9 2
18 0 9 1 0 9 2 1 5 2 1 11 0 1 12 2 12 2 12
3 9 2 11
7 1 0 9 13 9 1 9
5 11 2 11 2 2
17 3 12 9 0 9 12 9 15 13 1 0 0 9 11 2 9 2
21 1 0 9 9 1 9 12 9 2 9 4 13 12 9 1 9 7 12 1 9 2
13 9 1 15 3 13 0 9 1 0 7 0 9 2
11 1 9 1 0 9 15 3 13 12 9 2
14 0 9 0 0 9 13 1 12 1 12 9 1 9 2
14 3 13 9 1 9 9 2 3 3 13 1 10 9 2
28 9 9 0 9 13 1 3 16 12 9 1 12 9 2 3 3 15 13 7 1 0 9 2 16 13 12 9 2
18 13 15 7 2 16 15 9 0 9 1 3 0 9 0 9 3 13 2
14 9 9 1 0 12 0 9 13 3 1 12 9 9 2
19 13 7 0 13 2 16 13 9 9 1 0 9 2 0 12 1 12 9 2
14 0 0 9 11 2 9 15 13 1 9 12 2 9 2
5 0 9 2 9 9
31 0 9 0 0 9 2 11 2 2 15 15 13 1 11 2 13 0 0 9 11 11 9 2 16 11 13 0 9 13 0 2
21 9 2 15 4 13 13 0 9 1 9 10 9 2 15 13 1 11 13 0 9 2
15 15 13 1 9 10 9 1 9 9 13 1 0 9 11 2
14 3 10 9 13 1 10 9 13 7 13 1 0 9 2
26 9 0 9 2 9 7 0 9 1 9 9 15 13 13 3 9 1 11 7 0 9 13 1 0 9 2
21 9 15 3 13 13 1 11 13 9 2 7 10 9 2 14 1 9 12 12 9 2
20 1 0 9 13 11 9 2 15 13 0 1 10 0 9 3 1 12 0 9 2
15 1 0 9 13 9 11 3 13 9 11 7 1 10 9 2
18 0 9 1 0 9 13 0 9 2 3 0 9 7 9 1 0 9 2
3 0 9 9
7 9 0 11 15 13 1 9
3 0 11 2
13 9 9 13 3 1 0 9 3 9 0 11 11 2
24 1 12 9 1 10 9 1 9 11 13 7 3 1 0 9 1 12 2 9 9 14 1 11 2
25 9 13 13 9 1 9 9 2 3 13 9 12 2 12 2 7 1 10 9 13 1 9 9 11 2
21 1 12 2 7 12 2 9 13 9 11 7 11 7 15 4 1 3 0 9 13 2
8 1 9 15 13 9 0 11 2
16 1 0 11 13 3 3 11 11 2 7 16 3 14 1 9 2
24 0 3 13 12 2 12 2 16 1 12 1 9 13 11 11 2 7 9 13 1 12 2 12 2
21 9 15 3 13 12 9 1 9 11 2 7 1 10 0 9 13 1 9 9 11 2
3 11 13 9
2 11 2
15 1 0 9 11 1 11 13 11 11 12 9 1 0 9 2
26 1 15 4 13 4 13 9 1 10 0 0 9 2 15 4 15 13 3 1 12 2 12 9 1 9 2
16 9 0 0 4 13 4 13 1 0 9 7 3 3 9 9 2
15 2 1 9 1 9 9 13 1 11 9 9 1 0 9 2
16 9 9 14 1 9 4 13 13 9 0 9 1 0 9 2 2
25 1 9 9 0 0 13 9 9 1 12 0 9 13 2 2 3 3 13 9 1 9 3 0 2 2
26 11 3 13 1 0 9 2 2 13 0 2 16 0 9 4 13 1 0 7 0 9 1 9 3 13 2
12 9 13 11 11 2 11 11 7 11 11 2 2
1 9
9 0 9 9 9 1 0 0 9 2
6 11 13 9 9 1 11
3 0 11 2
17 9 11 11 1 11 0 11 4 13 0 9 11 9 12 2 12 2
21 11 13 12 9 1 12 0 7 10 0 9 11 11 1 9 11 11 15 13 12 2
9 0 0 9 13 11 11 1 11 2
30 9 0 9 11 2 12 9 2 13 1 0 9 0 9 12 9 1 9 2 3 12 0 9 2 12 9 7 12 9 2
45 11 13 0 9 11 2 15 13 1 12 9 13 9 9 9 2 12 2 2 12 0 9 2 12 2 2 12 9 2 12 2 2 12 9 2 12 2 7 12 0 9 2 12 2 2
23 1 0 12 9 15 15 13 3 12 9 2 11 11 2 3 11 11 7 11 11 2 11 2
1 9
5 13 9 9 11 2
2 11 2
4 0 9 1 11
6 11 9 2 11 2 2
24 0 0 9 1 9 11 1 9 9 13 0 9 9 11 2 15 15 3 13 9 0 9 9 2
9 11 13 3 13 14 1 0 9 2
10 1 0 12 3 13 3 0 0 9 2
5 13 0 9 11 2
10 9 11 11 11 13 9 2 15 13 9
2 9 9
50 1 0 9 1 0 9 9 11 2 11 2 12 2 12 2 4 13 2 16 0 9 11 11 2 12 9 2 9 11 11 11 2 1 0 9 0 9 1 11 1 11 1 11 2 12 2 12 2 13 2
4 11 11 2 11
38 1 10 9 4 13 9 9 7 0 0 9 15 1 0 9 13 9 1 12 2 12 2 12 2 13 1 11 2 2 9 9 13 13 1 12 2 12 2
24 11 15 3 13 3 12 9 1 0 9 2 9 1 9 7 10 9 7 9 0 9 15 13 2
17 2 11 15 13 9 11 2 15 13 1 9 13 1 0 0 9 2
6 13 2 16 13 9 2
14 9 9 1 11 15 3 13 2 2 13 9 11 11 2
15 9 9 13 2 16 11 13 13 1 0 9 14 16 9 2
24 3 15 13 13 11 11 2 11 2 2 15 15 7 1 9 13 7 4 13 1 9 1 9 2
22 1 0 12 0 9 1 0 0 9 2 1 9 12 2 15 12 1 15 13 0 9 2
14 13 7 3 3 0 2 16 11 15 1 9 3 13 2
30 1 9 14 3 3 13 1 9 12 9 7 1 9 1 0 9 2 16 11 13 9 9 2 15 13 7 9 0 9 2
9 11 13 0 9 9 16 10 9 2
18 1 12 9 2 1 15 12 9 2 15 1 12 9 13 3 12 9 2
21 3 7 11 11 2 15 13 1 9 11 1 11 11 14 1 0 9 2 3 13 2
20 9 9 12 0 9 13 7 13 2 16 10 3 0 9 3 13 3 1 9 2
35 2 13 4 15 13 1 9 2 7 13 4 15 13 1 9 2 16 4 10 0 7 0 9 13 1 15 13 9 9 2 2 13 11 11 2
33 0 9 3 13 2 16 10 9 3 13 9 2 1 15 11 3 13 1 11 2 16 4 1 9 13 13 1 11 7 14 1 11 2
30 2 13 2 16 0 15 3 4 13 2 16 1 11 2 14 4 13 10 9 2 15 4 13 3 15 0 2 2 13 2
23 9 11 11 0 9 1 0 9 13 7 1 9 9 13 9 2 16 9 13 10 0 9 2
3 11 3 13
2 11 2
19 7 1 9 0 9 1 9 13 1 0 9 11 7 1 0 9 11 11 2
13 9 0 0 9 1 15 13 9 1 9 9 12 2
27 1 9 15 7 13 13 2 16 4 11 13 4 3 13 1 9 7 16 1 10 9 13 11 11 1 11 2
3 13 4 2
2 11 2
3 0 9 11
2 11 2
16 0 0 9 1 12 2 9 11 9 13 1 11 11 11 11 2
11 1 9 1 12 9 13 1 9 12 9 2
28 0 13 11 11 11 9 1 12 9 0 2 13 7 0 9 1 9 2 16 13 1 9 9 1 9 12 9 2
7 9 15 13 11 11 11 2
20 1 0 9 13 11 11 1 9 7 9 0 9 7 1 0 9 13 0 9 2
13 1 0 9 1 12 9 13 0 0 9 11 11 2
16 3 0 9 13 11 9 11 11 2 9 15 13 11 11 11 2
15 0 9 11 11 13 0 0 9 7 1 0 9 0 9 2
3 11 3 13
15 0 9 13 3 7 0 0 9 2 15 3 13 1 11 2
29 9 11 11 11 1 0 9 13 2 16 13 0 9 3 13 9 1 9 9 1 9 2 1 15 3 13 1 9 2
15 0 9 13 7 9 9 9 2 15 4 13 9 1 9 2
22 1 9 13 3 9 13 9 2 1 15 4 13 1 9 13 1 9 9 7 9 9 2
5 0 9 13 13 2
13 10 9 4 13 13 3 1 11 11 12 2 9 2
5 9 1 9 15 13
14 9 11 13 9 11 1 11 12 2 12 7 13 3 9
2 9 9
7 0 9 11 1 11 11 11
20 9 11 13 1 9 9 9 9 1 9 11 12 2 12 7 13 3 0 9 2
22 16 4 11 13 0 2 13 4 15 3 0 9 1 9 2 15 11 13 3 1 9 2
5 12 9 13 3 2
29 3 0 11 13 3 1 9 1 9 1 9 14 9 2 1 0 9 3 11 3 13 1 7 1 9 11 13 9 2
17 1 12 2 9 7 13 9 1 0 9 2 11 1 9 13 9 2
31 0 11 3 3 11 13 1 10 9 2 15 7 3 13 13 9 7 3 9 11 13 14 1 12 2 9 11 9 1 9 2
13 9 11 3 13 12 9 2 7 11 15 0 13 2
27 1 0 9 2 12 9 2 15 9 9 3 13 1 9 11 2 7 0 9 14 3 13 1 0 0 9 2
19 11 3 14 3 13 9 7 16 11 1 12 2 9 13 1 2 13 13 2
5 11 2 13 4 0
23 9 0 9 9 11 11 1 9 13 2 16 10 9 13 16 3 2 2 13 4 0 2 2
17 3 13 14 0 2 16 15 3 1 15 13 1 11 14 1 9 2
23 0 9 9 11 11 14 13 0 9 7 13 2 16 11 3 13 1 12 1 0 9 11 2
16 2 3 4 15 7 13 2 16 1 9 2 2 13 1 9 2
20 1 9 11 13 3 0 9 9 12 0 9 2 15 13 12 9 1 0 9 2
21 1 9 7 1 9 13 1 11 3 7 3 2 3 2 3 1 0 9 9 9 2
30 0 0 9 1 9 12 7 12 9 2 9 2 1 9 12 7 12 9 2 9 2 0 0 12 7 12 9 2 9 2
24 1 9 13 9 1 12 7 13 1 12 9 2 9 13 1 9 1 12 7 13 1 12 9 2
10 0 9 1 0 9 1 9 13 0 2
2 9 3
2 11 2
4 11 0 9 9
11 1 11 13 3 9 16 1 12 9 0 9
2 9 9
5 11 2 11 2 2
19 1 0 0 9 0 0 9 13 11 11 1 0 9 11 3 12 2 12 2
11 0 2 16 0 9 13 1 9 11 11 2
21 9 0 9 11 3 13 1 12 2 9 1 9 12 2 12 9 1 0 9 11 2
34 2 9 13 1 10 9 0 9 16 0 9 2 2 13 11 1 0 9 2 3 11 13 12 2 12 1 3 0 9 2 15 3 13 2
6 0 9 13 9 13 2
17 2 1 9 4 13 0 9 2 7 11 1 9 13 15 0 13 2
15 1 12 2 9 13 11 2 15 4 15 13 1 9 13 2
21 16 4 7 13 2 16 9 13 1 15 3 3 7 13 1 10 9 2 13 4 2
25 7 11 15 1 15 3 13 2 13 7 15 4 13 0 0 9 7 3 7 0 2 2 13 11 2
12 3 1 0 0 9 13 11 0 9 2 2 2
17 2 7 3 3 4 15 13 2 1 0 9 4 13 12 9 2 2
15 11 13 3 1 0 0 9 3 1 9 3 16 0 9 2
23 15 11 13 0 9 2 2 16 4 15 3 13 2 13 4 13 1 0 12 9 3 9 2
18 1 11 15 15 13 2 7 9 9 13 2 16 1 9 15 3 13 2
13 15 13 3 0 16 11 2 1 15 13 1 9 2
12 3 9 13 10 9 2 15 13 3 3 15 2
11 9 1 0 9 15 3 13 1 9 2 2
8 7 1 9 15 3 13 15 2
25 9 13 9 7 1 9 13 12 12 9 2 15 13 3 16 1 15 0 9 1 12 0 9 2 2
22 1 9 0 0 9 9 2 11 13 1 11 2 11 1 11 2 13 7 9 0 11 2
18 2 16 15 13 2 3 13 9 3 1 9 2 16 13 2 13 0 2
16 7 3 13 15 0 2 13 9 2 7 3 15 13 13 15 2
13 15 3 13 9 2 7 3 3 1 15 9 13 2
15 1 9 9 7 4 13 7 13 0 9 2 2 13 11 2
2 11 11
5 9 11 11 2 11
9 1 9 11 13 3 9 16 1 11
11 1 0 11 15 1 0 11 3 3 13 4
2 9 9
5 11 2 11 2 2
18 0 0 9 2 11 2 13 9 9 9 7 9 15 13 7 0 9 2
19 0 9 1 9 1 9 7 3 13 3 13 2 13 15 9 1 0 9 2
34 9 9 2 11 2 15 13 12 0 9 2 1 15 13 9 0 3 2 1 0 12 9 15 4 13 12 2 7 12 2 9 1 9 2
14 0 9 4 13 9 9 7 3 12 9 1 0 9 2
15 11 13 12 9 9 2 0 7 0 7 3 13 1 0 2
33 15 13 2 16 3 1 11 4 11 13 0 0 9 2 16 0 11 2 16 13 9 2 13 9 0 0 9 2 15 13 0 9 2
37 0 12 0 9 13 0 9 7 1 15 4 1 0 9 1 0 0 9 13 7 11 2 13 2 14 9 2 0 0 9 13 1 9 9 0 2 2
21 9 11 15 13 0 9 9 2 1 15 13 12 0 9 2 3 3 16 1 11 2
32 7 3 12 0 9 2 15 15 1 9 3 1 9 9 13 2 7 3 0 1 9 0 9 13 9 2 13 2 1 9 11 2
27 1 10 9 4 13 11 14 12 9 7 2 4 2 14 13 11 9 11 7 13 2 14 2 13 7 15 2
23 13 7 3 0 2 16 9 2 15 15 13 1 9 9 2 13 9 0 9 2 7 3 2
32 3 11 1 9 0 9 4 15 1 9 9 13 2 7 13 9 2 16 1 15 4 13 9 9 7 0 0 9 2 2 2 2
10 10 9 15 11 4 13 14 1 9 2
26 9 9 15 13 13 0 2 7 9 13 1 9 2 3 0 9 13 0 2 7 1 9 9 15 13 2
27 9 13 2 16 9 2 15 15 13 1 11 2 4 13 1 9 11 2 7 11 13 3 0 9 2 2 2
19 7 10 9 15 4 11 13 14 1 9 7 9 9 15 13 1 0 9 2
8 0 9 13 13 1 0 9 2
29 1 12 9 1 9 11 15 3 4 13 1 0 1 9 9 1 0 9 9 2 12 9 4 13 13 1 0 11 2
13 7 15 15 7 13 0 9 2 3 15 3 13 2
3 11 1 0
2 11 2
31 0 9 9 0 11 1 12 2 0 9 13 1 0 9 11 11 7 11 11 2 15 13 0 0 9 11 9 7 11 11 2
15 11 13 1 0 9 3 1 11 11 1 0 9 9 11 2
10 9 0 9 13 9 1 12 2 9 2
18 0 13 9 0 11 7 11 11 7 13 1 10 9 12 9 9 11 2
4 11 13 1 9
5 11 2 11 2 2
11 9 9 11 3 13 9 7 13 14 0 2
23 9 11 2 11 13 9 2 7 1 9 15 1 9 11 2 11 13 1 10 3 0 9 2
38 2 9 9 1 9 2 13 9 1 9 9 11 7 11 2 1 15 15 13 7 9 2 7 0 0 9 0 9 11 2 15 13 3 2 7 11 2 2
18 9 2 3 9 3 13 1 9 1 11 9 7 11 2 9 11 2 2
29 9 4 15 0 13 3 1 10 9 2 7 4 13 2 1 10 9 13 1 0 9 0 7 15 4 1 11 13 2
6 11 13 12 9 5 9
2 11 2
42 11 11 2 0 9 11 1 0 9 13 13 0 0 0 0 9 2 15 13 9 3 12 9 5 9 7 15 13 1 9 11 2 11 11 1 9 12 1 9 1 11 2
18 2 13 13 0 3 0 9 2 3 9 1 9 2 3 1 0 9 2
20 15 3 13 1 11 9 9 11 2 15 13 0 13 14 9 12 9 5 9 2
22 3 9 12 9 5 9 4 0 1 0 9 13 2 2 13 12 0 9 7 0 9 2
5 14 11 2 7 11
5 11 2 11 2 2
22 0 9 10 0 9 1 9 1 9 9 13 11 2 3 4 3 15 13 2 7 11 2
13 1 9 13 0 9 1 9 15 0 9 1 11 2
31 2 13 15 2 14 4 1 9 12 2 3 13 3 12 9 0 2 3 13 1 9 2 2 13 10 9 9 9 11 11 2
15 1 11 4 9 9 11 13 1 9 12 2 9 1 11 2
32 9 1 9 2 9 1 9 1 11 13 2 13 1 0 9 2 3 4 13 3 2 1 12 10 7 0 9 1 0 0 9 2
32 0 0 2 0 9 15 13 13 9 1 0 9 2 15 1 3 0 9 13 3 0 9 0 9 2 0 9 2 0 11 3 2
10 3 0 9 4 13 0 9 1 11 2
18 3 0 9 9 13 9 1 9 1 11 2 3 15 13 9 1 9 2
8 2 11 2 9 11 11 2 11
13 3 1 11 2 0 9 13 1 0 9 2 0 9
10 0 9 13 1 9 3 0 9 1 9
2 11 2
23 0 9 1 0 9 1 11 4 3 13 13 9 2 10 9 1 9 3 13 1 0 9 2
19 9 0 9 1 0 9 11 7 0 0 9 0 9 13 9 3 12 9 2
12 3 15 13 9 0 9 11 2 9 11 11 2
29 9 9 1 0 9 2 15 13 13 1 12 2 9 13 0 9 0 1 11 2 13 1 12 9 3 1 12 9 2
21 1 0 9 1 11 13 3 0 9 10 9 7 13 3 7 12 0 9 1 9 2
18 9 11 13 2 2 16 15 13 15 2 16 0 9 10 9 13 2 2
22 0 9 13 1 9 1 12 2 9 3 12 0 9 11 9 0 9 1 9 1 9 2
22 1 9 0 9 3 13 13 7 12 9 2 15 4 13 0 9 2 13 11 2 11 2
5 0 9 1 9 9
2 11 2
26 0 9 11 11 3 1 11 13 3 13 0 0 9 9 2 16 10 9 13 0 9 1 9 9 11 2
40 11 15 13 13 10 9 9 7 13 1 10 9 0 9 1 9 0 9 9 12 2 12 3 0 9 9 2 1 11 2 13 11 1 9 1 0 9 11 11 2
12 3 13 2 16 1 11 13 9 11 1 11 2
19 13 0 2 16 4 11 13 9 11 0 9 1 0 0 9 2 13 11 2
15 11 13 13 9 1 9 1 11 2 15 13 12 9 9 2
21 1 9 1 11 15 13 9 0 0 9 7 0 9 2 3 1 9 9 7 9 2
9 0 9 11 2 11 7 11 2 11
4 11 2 11 2
29 9 11 7 11 11 11 7 11 11 13 12 2 9 1 0 11 0 9 9 1 9 9 9 2 9 2 11 2 2
14 13 15 3 1 11 7 1 11 0 9 9 12 9 2
49 0 9 13 12 13 1 10 3 0 9 1 0 9 7 9 7 1 15 2 16 11 7 11 15 13 13 1 0 0 9 7 3 15 13 1 9 14 10 9 2 7 7 9 0 0 7 0 11 2
27 9 0 9 9 13 2 16 11 11 13 9 10 9 1 0 9 7 13 2 16 15 1 0 11 3 13 2
13 13 4 15 1 10 9 1 11 1 0 0 9 2
38 2 9 13 9 0 9 12 9 2 10 9 7 0 9 2 15 15 13 9 9 7 0 9 0 0 9 2 2 13 3 11 0 9 0 9 11 11 2
23 0 9 1 15 13 3 9 12 9 1 9 1 9 1 10 9 7 9 13 1 10 9 2
17 12 9 15 13 1 9 2 15 13 0 1 15 9 1 9 9 2
7 11 2 11 13 1 9 9
2 11 2
26 0 9 1 11 11 11 3 13 1 11 1 9 0 9 11 2 11 7 1 9 0 9 11 2 11 2
18 13 1 9 0 9 9 0 9 11 2 11 2 11 2 11 7 11 2
7 0 9 2 11 13 3 0
2 11 2
37 1 0 9 0 0 9 1 0 9 2 15 15 13 13 9 0 0 11 11 2 13 1 0 9 11 1 12 9 1 12 2 0 7 0 2 9 2
20 1 0 9 11 15 1 10 0 9 2 15 13 1 9 2 13 0 9 11 2
38 9 13 2 0 9 11 2 0 9 11 2 15 13 1 9 12 1 9 2 13 0 1 9 2 7 7 13 0 9 9 1 0 9 2 2 13 11 2
31 1 0 9 0 9 9 9 1 11 3 13 2 16 9 9 2 0 16 0 2 15 1 9 12 1 9 12 3 16 13 2
4 3 0 16 9
7 9 13 3 0 0 9 2
5 9 13 13 9 9
7 13 9 2 13 2 13 2
6 13 10 0 9 0 2
19 0 9 3 0 9 1 9 11 12 2 1 9 12 2 13 3 12 9 2
17 1 9 15 9 13 0 9 12 9 11 12 1 12 7 12 9 2
35 1 9 15 3 13 3 9 2 16 9 9 3 13 1 9 0 9 16 1 9 9 2 7 7 3 13 9 9 9 3 3 0 16 9 2
19 3 3 13 0 9 2 13 13 9 2 9 2 9 2 9 0 9 3 2
35 0 9 9 1 0 9 2 3 15 3 13 9 2 1 15 3 13 2 13 3 0 9 1 9 10 9 2 7 13 1 0 9 0 9 2
37 16 9 9 13 13 13 15 15 1 9 9 1 10 9 2 13 0 3 3 13 2 3 13 0 10 9 2 0 1 9 2 13 14 16 0 9 2
36 16 4 13 9 1 0 9 3 0 2 13 0 0 9 11 0 9 1 9 11 12 2 15 15 13 1 0 9 0 9 2 15 13 9 0 2
16 9 2 9 9 0 9 1 0 9 2 13 3 13 1 9 2
13 1 0 9 7 0 9 13 10 9 16 1 9 2
15 1 15 7 9 13 7 15 9 1 9 9 13 10 9 2
16 16 9 13 3 2 13 9 9 3 3 2 16 9 13 3 2
21 3 15 7 3 13 13 2 16 0 2 0 9 1 9 13 0 9 14 1 9 2
22 7 15 13 13 1 15 3 9 1 9 2 15 13 1 0 9 9 2 0 0 9 2
36 9 2 0 10 9 2 13 0 9 1 9 2 3 0 9 2 7 1 9 9 1 9 13 9 0 9 3 3 2 16 13 15 9 13 3 2
31 0 9 15 15 3 13 1 9 9 1 9 2 15 13 9 1 0 9 9 2 16 15 2 15 4 3 13 2 13 0 2
19 0 9 0 9 0 9 9 3 13 2 7 7 3 13 9 3 0 9 2
32 13 15 15 2 16 1 9 13 10 9 13 1 9 2 15 13 1 15 10 9 2 0 1 0 9 2 7 1 12 9 3 2
10 3 15 13 2 16 4 15 9 13 2
31 13 4 2 16 13 9 1 9 2 7 10 9 13 1 3 0 2 16 9 13 13 1 9 2 15 13 1 15 1 9 2
17 3 15 1 10 9 13 9 9 3 2 16 13 1 15 3 9 2
26 1 0 9 13 7 0 1 9 9 13 14 1 0 9 1 0 9 2 7 7 1 9 1 0 9 2
10 0 9 9 13 9 9 1 0 9 2
23 12 9 11 12 0 9 13 14 12 9 2 16 4 13 1 9 12 2 12 7 12 9 2
27 1 0 9 13 14 1 12 5 0 2 7 7 15 1 9 0 9 13 7 1 15 2 10 9 9 13 2
12 0 9 9 13 13 1 9 1 9 12 9 2
10 9 0 9 13 10 9 1 9 9 2
5 3 13 0 9 2
24 13 15 15 3 13 2 16 1 9 2 15 13 1 9 1 9 2 15 1 9 13 9 0 2
15 7 7 1 0 9 1 0 0 9 3 3 13 10 9 2
30 10 9 13 2 16 15 13 9 2 3 3 0 2 15 13 9 0 2 9 7 0 9 7 13 1 0 7 0 9 2
38 12 9 10 9 13 0 12 9 2 7 3 13 13 1 15 2 16 12 9 1 9 0 9 2 1 9 1 9 3 12 9 2 13 1 12 9 3 2
30 1 9 2 15 13 0 9 9 2 3 0 16 0 2 15 3 13 0 9 2 7 0 9 13 12 7 12 12 9 2
13 9 9 1 12 9 15 13 1 12 7 12 12 2
23 9 9 0 0 9 13 7 3 0 16 1 0 9 7 9 9 13 3 1 0 9 0 2
34 9 10 9 13 3 13 14 16 9 2 7 3 7 16 0 9 2 7 15 7 3 1 9 0 9 2 15 4 1 9 13 1 9 2
13 1 0 9 13 13 9 0 9 9 1 0 9 2
22 13 13 1 12 9 9 13 14 12 9 7 9 0 9 4 4 13 14 1 12 9 2
17 9 9 1 12 9 4 13 13 3 1 12 12 9 9 0 9 2
25 10 9 4 15 13 13 7 1 10 9 1 0 9 2 7 3 1 9 13 7 13 7 13 9 2
17 1 10 9 9 13 0 9 9 0 9 2 9 3 2 0 9 2
12 7 15 1 9 9 13 3 13 10 0 9 2
12 1 9 10 9 13 13 10 9 2 7 15 2
5 2 9 9 9 2
7 3 13 15 1 9 12 2
10 0 9 9 9 13 14 1 9 9 2
12 16 15 13 3 9 2 13 10 9 0 9 2
18 1 15 0 9 9 9 13 3 15 1 0 9 2 15 13 9 3 2
4 2 9 9 2
7 13 9 7 3 0 9 2
5 15 13 0 9 2
13 10 9 15 13 9 3 2 1 0 4 13 3 2
4 2 0 9 2
21 13 2 1 10 9 15 13 3 2 15 13 1 9 9 9 2 12 9 0 9 2
14 0 9 13 12 9 1 9 2 0 12 9 1 9 2
14 3 0 9 2 12 9 1 9 2 13 14 10 9 2
9 0 9 13 3 12 9 1 9 2
16 9 0 0 9 3 13 9 9 7 9 2 7 3 13 9 2
16 16 15 13 3 1 9 9 2 3 13 3 0 12 9 9 2
11 13 9 2 15 13 0 9 7 13 3 2
24 0 9 13 9 1 9 0 9 2 7 3 13 1 12 0 9 13 3 9 2 3 7 9 2
13 1 10 9 13 0 15 13 9 2 0 1 9 2
12 15 0 9 13 2 16 13 9 2 7 9 2
14 15 3 0 9 13 0 1 9 2 16 13 0 9 2
16 3 0 13 9 9 0 9 2 7 15 1 9 10 9 13 2
12 1 9 13 7 9 2 9 2 9 7 9 2
10 3 0 9 0 9 4 15 13 13 2
26 9 2 0 3 2 16 15 1 15 13 15 3 13 2 16 4 9 13 0 9 2 13 13 3 0 2
14 10 9 13 13 3 0 9 2 15 15 13 0 9 2
24 10 9 13 1 9 13 0 9 7 13 9 9 7 9 2 3 13 4 13 9 7 9 9 2
9 9 15 3 13 7 1 10 9 2
19 13 15 13 1 9 9 2 3 15 13 0 9 1 9 2 3 1 9 2
30 16 4 13 10 9 2 13 4 15 0 9 2 16 13 9 14 1 9 2 15 4 13 2 13 2 1 10 0 9 2
17 3 15 12 9 0 9 2 3 1 9 2 13 9 1 0 9 2
9 13 15 1 10 9 1 9 9 2
25 0 15 13 13 1 9 1 9 1 9 3 9 0 9 2 0 9 9 2 9 9 7 9 0 2
12 1 10 9 15 9 7 9 1 9 9 13 2
12 0 9 0 2 9 13 4 13 7 1 9 2
27 13 9 1 9 2 7 13 9 0 7 0 10 0 9 2 16 4 3 13 1 9 1 0 9 0 9 2
15 13 15 2 16 13 1 9 2 15 13 9 0 9 13 2
34 1 0 11 13 3 0 9 1 9 9 2 15 4 13 15 2 16 15 1 9 9 13 9 2 0 1 9 2 15 4 1 15 13 2
16 9 13 0 9 1 0 9 7 9 7 1 15 13 0 9 2
11 9 13 13 7 13 14 9 1 0 9 2
40 3 13 15 9 2 15 9 15 13 2 7 15 13 1 15 2 16 9 2 0 2 16 13 9 7 1 0 9 9 2 13 1 15 9 1 9 7 3 3 2
28 16 13 1 9 2 15 15 9 7 9 13 2 3 4 15 13 13 0 9 2 3 10 2 1 15 3 13 2
26 3 13 0 9 1 9 2 15 1 9 9 7 9 13 3 7 13 15 2 16 4 15 15 15 13 2
2 11 11
10 15 13 13 1 0 9 1 0 9 2
18 2 0 9 3 1 12 7 12 9 1 12 9 11 12 0 9 11 2
10 2 3 12 9 9 2 9 7 3 2
5 2 12 9 9 2
4 2 9 9 2
13 2 9 1 0 9 1 9 1 9 3 12 9 2
12 2 9 1 9 9 1 9 2 3 12 9 2
7 2 9 9 1 0 9 2
9 3 0 2 7 3 0 0 9 13
10 2 0 9 9 2 0 0 9 2 2
7 2 12 7 12 9 9 2
13 2 12 9 9 2 9 2 3 2 3 3 2 2
6 2 0 9 0 9 2
17 2 9 1 9 1 0 9 9 16 12 7 1 9 2 0 2 2
14 2 0 9 9 1 0 7 0 9 2 9 9 3 2
19 2 9 9 1 0 9 1 0 9 9 2 1 0 9 2 7 1 9 2
5 2 9 0 9 2
10 2 9 3 1 12 0 9 11 12 2
17 2 9 0 9 3 12 9 12 9 7 12 7 3 9 12 9 2
8 2 0 9 9 0 0 9 2
12 2 9 0 9 9 1 0 9 0 0 9 2
4 2 9 2 2
12 2 9 9 9 1 3 9 1 0 9 9 2
8 9 9 2 9 4 3 13 13
13 2 0 9 1 9 9 7 9 1 9 0 9 2
6 2 9 9 0 9 2
4 9 1 9 2
10 2 9 4 13 1 0 9 0 9 2
24 2 0 9 9 9 0 9 2 7 2 0 9 1 0 9 2 4 1 10 9 13 9 9 2
10 2 1 9 13 9 9 1 9 9 2
9 13 3 1 0 9 11 12 11 2
2 9 2
3 9 3 0
10 1 9 3 13 1 12 9 9 1 9
36 9 9 12 4 13 9 1 9 2 15 13 2 1 9 14 9 2 7 7 0 0 7 0 9 2 13 0 9 9 9 2 15 15 3 13 2
13 3 7 1 15 13 7 3 1 0 9 7 13 2
2 11 11
22 15 13 3 9 9 0 9 9 11 1 0 7 0 9 2 1 15 15 0 9 13 2
17 3 13 9 11 11 2 9 13 10 9 1 0 9 7 9 9 2
24 13 1 0 9 9 2 7 13 7 0 9 9 2 15 13 2 16 15 15 9 13 7 14 2
14 3 0 9 13 9 2 15 3 9 2 15 3 2 2
9 9 13 9 10 9 9 0 9 2
17 9 13 9 9 7 15 13 0 9 9 2 9 13 7 9 0 2
4 12 2 12 3
22 13 15 15 13 9 1 0 9 9 2 1 15 13 9 13 2 0 9 2 9 9 2
19 1 9 9 11 11 11 13 1 0 9 3 13 1 12 9 9 1 9 2
10 9 10 9 13 7 13 0 9 9 2
26 7 15 13 2 3 0 2 0 2 15 13 2 16 9 13 1 9 3 12 2 12 9 9 1 9 2
32 13 14 13 2 16 1 12 2 9 12 2 3 1 9 2 13 2 3 12 9 2 13 0 14 9 9 9 3 1 12 9 2
4 15 1 15 11
37 1 0 9 1 11 2 11 2 11 2 9 7 1 0 11 4 15 13 2 16 3 15 0 9 1 9 15 13 3 0 2 3 3 0 0 9 2
5 7 15 15 0 2
27 2 1 9 0 9 9 7 9 9 11 4 15 13 2 16 13 1 15 0 0 9 3 15 13 1 9 2
18 1 9 13 9 9 9 11 11 2 15 1 0 0 9 9 13 9 2
16 15 13 3 0 9 7 13 1 15 2 3 13 9 0 9 2
10 10 9 1 9 9 9 3 3 13 2
21 9 13 2 16 0 9 13 13 10 0 9 7 3 13 3 13 1 10 0 9 2
18 9 9 9 15 13 12 0 9 2 0 9 2 0 9 7 0 9 2
11 10 9 3 13 0 9 0 0 0 9 2
36 13 7 0 13 2 16 15 3 3 1 12 9 7 1 12 12 9 13 0 9 1 15 2 16 10 7 0 0 9 2 9 2 0 9 13 2
2 9 9
27 9 9 2 9 2 7 3 2 13 3 1 9 9 13 3 3 2 16 1 9 9 2 9 7 0 9 2
25 16 9 13 3 14 9 2 7 3 9 1 0 9 2 13 9 2 16 4 4 9 13 1 9 2
52 7 15 3 13 1 9 2 16 7 1 9 9 2 15 13 7 9 2 7 9 1 15 2 15 9 13 1 9 9 9 14 1 9 2 16 13 9 2 15 13 1 9 13 2 3 9 2 9 7 3 2 2
21 13 2 14 3 1 0 9 1 10 9 2 13 0 2 16 0 9 9 3 13 2
12 9 15 3 13 2 7 9 0 9 13 0 2
1 3
3 0 0 9
22 9 2 16 9 16 9 0 1 9 9 7 9 13 1 10 9 13 2 13 3 0 2
24 7 15 3 13 15 0 2 16 0 0 9 2 15 1 0 9 0 9 7 13 2 7 13 2
2 11 11
42 10 9 3 13 9 12 2 9 2 3 0 0 9 13 2 16 1 0 0 9 1 11 13 9 1 9 0 7 0 9 2 1 15 1 9 0 9 13 0 0 9 2
23 10 9 3 13 9 11 11 11 9 2 16 9 0 9 11 1 0 9 13 9 0 9 2
30 16 9 1 0 9 0 9 13 2 16 1 9 9 13 15 0 9 2 3 7 15 0 2 13 0 9 1 12 9 2
31 1 9 0 0 9 4 15 13 2 16 10 9 1 9 0 7 0 9 3 13 1 15 2 3 13 12 0 9 1 9 2
41 9 3 13 9 0 9 1 9 2 3 1 15 3 13 9 1 9 9 9 2 15 4 13 0 9 1 0 1 9 0 0 0 9 1 9 0 9 1 0 9 2
32 13 2 14 9 2 16 0 7 0 9 4 13 1 9 2 3 15 15 13 1 9 9 2 16 13 0 9 9 1 0 9 2
20 10 9 1 0 9 13 12 9 9 2 0 7 13 9 3 1 12 9 9 2
19 1 9 0 9 4 7 3 3 13 7 2 13 2 0 2 3 0 9 2
24 1 11 11 7 13 2 16 4 9 0 7 0 9 13 13 0 9 1 9 0 0 0 9 2
15 15 15 13 0 9 2 3 15 13 3 1 0 9 3 2
28 0 9 2 15 13 10 0 9 1 9 0 9 2 2 13 2 13 9 9 2 16 9 10 9 13 3 9 2
43 13 2 14 15 7 2 16 0 0 9 1 0 9 3 13 0 9 9 2 13 3 2 16 0 9 9 0 7 0 1 3 0 0 9 13 15 3 3 13 1 10 9 2
8 9 13 1 9 2 7 1 9
8 11 11 13 9 9 1 0 9
10 9 4 13 2 13 2 14 9 9 2
6 3 13 9 11 11 2
37 0 9 9 9 2 0 1 9 12 2 9 0 9 2 0 9 0 9 7 0 9 15 13 9 2 3 9 0 9 13 10 0 9 1 0 9 2
63 1 9 2 0 9 9 9 9 2 15 15 3 13 9 3 13 9 1 3 0 9 2 11 11 13 9 2 16 1 0 13 2 16 9 13 3 13 9 0 9 2 1 10 9 0 1 10 9 9 7 9 10 9 2 15 4 13 0 9 0 0 9 2
21 13 2 16 13 14 1 0 9 1 3 0 9 9 2 7 3 9 0 0 9 2
30 16 4 9 13 1 0 9 2 15 0 9 2 0 1 9 3 13 2 13 0 9 3 1 0 9 0 9 3 0 2
30 1 9 2 1 10 9 2 10 0 9 4 13 13 15 0 0 9 9 3 7 1 9 2 4 15 13 10 9 9 2
19 11 9 2 9 0 9 0 9 2 10 9 13 1 15 16 9 14 3 2
15 1 9 15 15 13 2 7 3 3 3 2 3 7 3 2
36 16 13 1 0 9 2 13 4 13 14 3 0 2 16 9 13 0 7 9 9 13 14 14 1 9 2 15 4 15 13 13 1 9 1 9 2
18 3 15 15 7 4 13 0 9 2 16 15 13 13 13 9 10 9 2
30 12 9 13 0 2 11 13 0 0 9 7 1 10 0 9 13 0 9 7 9 1 9 3 2 15 3 13 3 13 2
37 13 0 9 2 15 0 9 4 13 10 9 2 7 15 15 3 13 14 9 2 7 15 2 2 1 15 0 0 9 4 15 13 16 10 9 13 2
27 13 1 9 14 0 9 2 7 3 9 2 3 0 9 13 9 2 15 13 1 9 2 9 1 0 9 2
21 9 2 16 13 1 0 9 9 2 13 3 1 9 0 9 2 0 7 1 9 2
20 16 13 2 16 15 15 10 0 2 0 9 2 3 13 2 14 13 3 9 2
31 13 2 16 13 9 9 2 3 15 0 9 13 9 3 1 9 2 3 3 15 0 9 1 9 13 13 1 10 0 9 2
8 7 3 1 15 13 13 0 2
54 11 11 2 0 9 0 9 2 0 2 9 2 2 11 2 11 2 13 0 2 16 3 15 13 1 15 2 16 9 1 9 0 9 15 13 1 9 1 0 9 9 9 2 7 0 9 1 0 9 9 7 10 9 2
44 10 9 4 15 3 13 13 2 16 15 15 0 9 13 2 16 1 0 9 13 3 12 9 9 0 9 2 15 13 1 9 1 10 9 2 9 2 1 0 9 3 0 9 2
35 16 4 15 7 13 9 9 1 9 12 2 3 13 13 0 9 2 9 9 0 9 3 3 13 2 7 13 9 9 2 3 15 3 13 2
28 16 13 9 2 15 13 1 9 3 16 15 2 16 0 9 2 3 10 9 13 2 13 13 15 9 9 9 2
30 1 15 3 13 0 0 9 2 3 0 9 9 9 2 7 0 9 2 13 0 9 1 0 9 7 9 0 9 9 2
56 16 7 13 1 9 13 0 9 0 9 9 2 3 3 13 2 16 15 13 13 3 0 9 3 9 2 14 3 13 1 9 10 9 2 2 3 13 2 16 3 13 10 9 2 2 3 1 0 9 1 9 7 10 0 9 2
40 13 10 9 2 16 0 9 13 3 3 2 1 9 13 1 9 10 9 2 7 16 15 13 13 2 3 13 7 0 9 7 10 9 1 9 3 0 0 9 2
3 9 1 9
7 15 15 13 2 13 9 2
9 13 2 3 3 2 2 13 9 2
6 11 1 11 1 12 9
13 7 1 0 0 9 9 12 13 0 9 1 0 0
18 1 9 0 9 13 1 9 11 11 9 0 9 1 9 1 11 11 2
39 13 15 15 1 9 2 3 9 10 9 0 9 13 9 12 9 9 2 1 9 0 9 15 3 13 9 7 13 15 7 9 1 9 10 9 1 0 9 2
6 13 11 11 7 11 11
40 9 3 1 9 12 2 12 3 1 0 9 11 13 1 9 0 9 2 9 0 2 9 0 3 1 15 2 3 13 9 1 9 11 2 1 15 15 11 13 2
6 13 3 10 0 9 2
26 3 11 11 13 0 9 1 10 9 1 0 9 0 9 11 2 15 1 11 11 13 13 1 0 9 2
15 13 4 3 9 2 15 0 9 13 1 0 9 1 0 2
42 7 16 3 13 9 2 1 15 13 13 0 9 9 0 0 9 2 9 1 0 9 9 7 0 9 11 11 11 11 2 1 9 2 4 13 9 0 15 1 0 9 2
21 2 3 4 13 0 1 9 1 9 1 9 9 0 9 7 9 9 9 0 9 2
7 13 15 15 13 0 9 2
13 13 15 9 9 9 7 3 4 13 0 0 9 2
11 2 13 15 7 3 2 16 4 3 13 2
18 14 2 9 4 13 7 0 9 13 14 1 9 9 2 1 9 9 2
35 13 2 16 15 13 3 7 2 16 15 13 0 9 10 9 1 10 0 9 1 11 7 3 1 10 9 2 1 15 4 13 1 0 9 2
15 13 15 15 15 13 9 2 15 15 1 10 9 3 13 2
15 2 3 4 13 0 9 3 1 0 9 2 3 1 0 2
12 13 15 9 2 7 0 9 13 0 15 13 2
9 0 9 4 3 13 1 12 9 2
15 0 13 1 15 2 16 13 3 9 13 15 1 9 11 2
28 0 9 13 10 9 2 16 9 9 2 3 0 9 15 13 13 2 7 3 3 13 0 9 0 1 0 9 2
5 9 13 0 9 2
12 0 9 13 3 3 13 2 13 9 13 9 2
6 3 3 1 15 13 2
15 13 0 9 9 1 11 2 15 4 13 7 1 10 9 2
17 2 16 0 9 4 15 13 9 9 9 2 0 9 7 0 9 2
8 13 2 16 9 9 15 13 2
6 3 13 15 1 0 2
12 16 4 13 2 13 1 11 3 16 12 9 2
10 1 9 10 9 4 13 3 12 9 2
6 2 15 13 0 9 2
5 3 15 13 0 2
20 15 15 2 15 12 9 2 13 0 1 15 2 3 3 4 13 0 9 9 2
11 16 4 13 3 2 13 15 13 7 9 2
14 4 2 14 13 3 2 13 0 13 1 0 9 9 2
10 15 13 2 16 15 15 13 13 9 2
5 7 9 13 10 2
8 2 1 10 9 4 13 9 2
21 13 4 1 9 13 10 9 9 2 15 13 1 9 9 2 1 15 13 13 9 2
25 13 4 15 3 13 15 0 9 2 13 0 0 9 9 7 13 3 2 16 4 10 9 13 13 2
9 2 13 4 3 3 9 0 11 2
11 13 4 1 15 1 9 9 3 0 9 2
22 10 9 1 9 9 9 13 13 9 0 2 16 0 9 2 7 3 13 0 0 9 2
15 3 4 13 9 10 0 9 2 16 4 15 13 0 9 2
22 13 13 0 9 1 15 0 9 7 13 3 1 0 9 2 15 4 13 16 10 9 2
26 13 7 13 2 16 4 15 0 9 13 1 0 9 1 9 9 1 0 9 2 15 4 13 0 9 2
24 13 4 3 2 16 10 9 2 3 9 2 15 4 13 1 0 9 7 1 11 2 4 13 2
14 15 2 16 4 13 0 9 2 13 4 15 10 9 2
12 2 13 12 1 9 9 9 3 9 9 9 2
13 3 4 13 0 9 1 9 2 15 13 1 9 2
17 13 15 3 2 7 9 13 13 9 10 9 7 10 9 1 9 2
15 1 15 4 3 13 9 2 7 13 15 14 1 0 9 2
25 3 13 13 3 1 0 7 0 9 2 7 15 3 2 16 4 15 13 13 9 9 2 15 13 2
17 2 16 11 13 1 11 2 13 3 9 9 2 15 9 9 13 2
7 13 3 1 9 0 9 2
6 3 13 15 1 15 2
18 7 15 4 13 9 1 9 2 15 11 1 0 9 7 0 9 13 2
7 13 9 1 10 0 9 2
21 1 15 4 13 0 9 1 9 9 1 10 9 7 3 4 13 9 1 10 9 2
11 9 10 0 9 13 0 2 7 13 0 2
25 3 4 13 0 9 2 16 4 13 0 9 1 9 9 7 3 13 1 10 9 1 10 0 9 2
7 2 1 9 9 13 9 2
18 1 9 11 15 13 15 2 16 9 0 9 13 7 0 2 7 0 2
3 15 13 2
12 13 0 9 1 9 1 9 1 10 0 9 2
14 13 2 16 13 11 9 1 0 9 7 15 13 0 2
11 13 4 15 2 16 15 13 1 0 9 2
5 13 2 16 14 2
12 16 1 0 13 3 2 13 15 1 0 9 2
7 7 3 1 15 3 13 2
20 13 4 2 14 13 9 1 0 9 2 7 3 3 13 0 13 1 0 9 2
18 13 15 2 16 10 9 13 3 1 9 7 16 1 15 13 15 13 2
5 13 1 9 9 2
16 7 13 13 2 16 4 11 13 3 0 9 16 0 0 9 2
18 2 7 16 9 13 9 15 2 15 0 9 2 13 15 9 13 9 2
16 7 1 9 13 0 2 16 9 0 9 13 0 16 9 9 2
15 7 1 10 15 4 13 13 11 1 9 2 15 13 0 2
18 13 2 14 9 9 2 13 15 3 3 13 11 1 9 11 1 11 2
17 1 15 4 13 9 0 13 0 0 9 7 1 10 9 4 13 2
8 2 13 9 1 3 0 11 2
5 13 3 1 11 2
21 7 3 13 9 1 0 9 2 16 4 13 2 16 13 9 1 9 1 0 9 2
8 1 15 15 13 1 15 0 2
15 13 11 2 16 4 13 9 9 10 10 9 1 9 11 2
15 2 0 1 10 0 9 13 13 1 11 1 9 0 9 2
7 1 10 9 15 15 13 2
2 3 2
6 13 1 9 10 9 2
13 1 9 11 13 3 9 2 16 13 1 10 9 2
19 3 15 9 13 2 16 15 0 9 2 15 0 13 0 9 7 9 9 2
10 13 4 15 3 0 1 9 10 9 2
9 13 4 0 0 9 1 10 9 2
15 3 3 0 1 9 0 9 13 9 0 9 1 9 9 2
16 1 9 3 13 9 2 13 2 14 15 0 2 16 4 13 2
14 2 16 4 13 1 11 2 3 13 10 10 0 9 2
5 3 3 13 9 2
2 14 2
5 4 13 0 9 2
15 1 15 13 0 9 2 1 15 4 13 10 7 15 9 2
14 0 0 9 10 0 9 13 13 10 9 1 0 9 2
18 3 4 13 9 1 0 9 2 16 4 1 10 9 13 0 0 9 2
24 1 0 12 9 4 13 9 1 9 1 11 2 11 2 11 2 11 7 1 12 0 9 13 2
19 13 3 0 0 9 1 11 7 1 0 9 13 9 1 0 9 1 11 2
10 2 11 13 0 9 1 12 9 3 2
14 13 15 7 2 16 3 0 9 9 3 13 0 13 2
20 3 4 13 0 9 1 9 0 9 2 16 4 13 13 0 9 1 0 9 2
16 16 4 13 13 7 13 3 12 9 1 9 2 13 0 9 2
15 7 13 0 9 13 3 12 9 3 2 14 2 14 3 2
12 16 4 15 13 13 2 3 4 15 13 13 2
18 16 15 13 13 9 1 3 9 2 13 9 9 1 0 9 7 13 2
9 2 3 2 15 13 0 9 11 2
8 15 12 9 3 15 3 13 2
14 15 13 2 16 1 12 9 7 15 12 12 13 0 2
16 11 15 3 13 13 0 9 1 9 1 9 2 3 13 9 2
7 9 10 9 15 13 13 2
12 13 1 9 9 10 9 3 1 0 9 0 2
15 2 13 4 2 16 11 13 0 1 9 3 12 9 3 2
7 3 7 13 1 12 3 2
6 14 2 7 13 0 2
15 2 13 2 14 1 10 9 2 13 3 9 2 7 9 2
21 3 2 16 4 3 3 13 2 4 13 2 16 13 9 9 1 9 12 9 3 2
27 16 4 7 13 13 1 15 2 16 4 13 9 3 1 9 2 15 13 0 13 2 9 9 15 13 13 2
15 12 1 10 9 13 13 1 10 9 9 2 15 13 9 2
27 3 3 13 7 13 2 13 3 9 2 7 13 9 3 2 16 4 13 0 1 9 3 16 12 9 3 2
9 13 2 16 15 15 13 13 9 2
13 2 16 4 13 1 11 2 0 13 9 9 11 2
10 1 3 3 13 10 9 1 15 13 2
9 3 4 15 13 13 9 1 9 2
13 9 13 0 9 1 9 2 1 9 7 1 9 2
9 2 3 13 9 0 9 0 11 2
7 13 3 13 9 10 9 2
14 3 15 13 2 16 4 13 2 3 3 13 0 9 2
8 7 3 13 13 9 7 9 2
9 2 13 15 1 10 0 0 9 2
7 13 0 9 1 9 12 2
19 13 4 9 2 16 9 9 12 13 13 15 1 10 0 9 2 3 13 2
10 11 4 13 13 9 9 2 10 13 2
8 3 0 9 1 9 1 9 2
6 3 13 0 10 9 2
16 7 1 15 4 13 13 9 2 3 13 9 7 1 0 9 2
6 2 7 15 0 9 2
8 3 4 15 13 10 0 9 2
12 3 14 2 1 15 4 13 13 1 10 9 2
18 13 13 9 2 15 13 13 1 0 9 2 16 4 15 10 9 13 2
8 15 4 13 1 0 0 9 2
21 2 1 10 9 3 13 2 16 9 0 9 1 11 2 3 1 11 13 0 9 2
3 15 13 2
19 13 3 13 9 2 13 0 9 7 9 1 9 0 9 13 1 9 9 2
7 13 3 0 13 10 9 2
27 2 1 15 13 10 9 1 11 0 7 1 15 15 13 1 9 2 1 15 4 15 13 1 9 1 11 2
6 9 12 9 13 0 2
12 3 15 13 2 16 1 12 9 15 3 13 2
12 0 9 11 13 2 16 15 13 0 0 9 2
11 15 4 13 2 7 1 9 4 13 15 2
8 1 15 11 13 3 0 9 2
15 0 9 13 1 15 2 16 9 11 13 3 0 16 11 2
22 13 0 13 0 9 9 1 9 9 1 11 2 16 3 13 3 9 7 3 10 9 2
20 2 1 15 15 1 3 16 12 9 9 1 11 13 10 9 7 1 15 14 2
16 13 15 1 15 2 16 9 13 3 3 0 2 3 4 13 2
14 1 15 13 4 2 16 0 7 0 9 11 13 0 2
18 7 13 15 2 16 13 15 3 0 2 16 3 3 13 0 9 9 2
7 3 3 7 13 1 9 2
29 2 3 13 0 9 9 1 15 2 16 9 1 0 11 13 2 16 4 15 13 0 9 15 12 1 0 0 9 2
6 10 9 15 3 13 2
11 16 15 13 2 3 13 10 9 1 11 2
17 1 10 9 4 13 1 10 0 9 2 1 10 9 2 1 11 2
6 2 3 15 13 3 2
9 1 0 9 13 15 9 1 11 2
15 13 7 3 13 2 16 1 0 9 13 3 13 10 9 2
27 2 15 13 10 9 13 1 12 9 9 11 2 15 13 1 9 2 16 9 1 0 9 1 11 4 13 2
8 13 1 15 16 1 0 9 2
3 13 1 9
11 16 9 9 3 13 2 1 9 13 3 3
17 1 9 0 9 13 0 0 9 7 1 15 14 0 9 9 9 2
11 13 15 2 16 0 9 3 13 13 0 2
12 7 3 13 12 1 0 9 1 9 1 11 2
4 15 15 13 2
2 9 2
23 15 10 9 1 9 13 13 2 16 15 2 0 3 2 14 2 7 15 13 9 9 11 2
2 11 11
13 9 9 9 13 0 9 9 9 7 9 0 9 2
11 9 9 1 0 0 9 13 9 10 9 2
12 13 10 9 2 7 13 15 3 0 0 9 2
7 1 15 15 13 9 9 2
22 9 1 10 9 4 1 12 5 13 9 9 2 10 9 1 0 9 1 0 9 13 2
29 3 0 9 13 9 9 2 14 12 5 2 2 9 2 14 12 5 2 2 7 9 7 9 2 1 12 5 2 2
10 9 15 1 0 9 13 3 12 9 2
22 13 2 14 15 3 0 9 9 1 12 9 9 2 12 9 1 10 13 1 9 9 2
2 13 15
35 7 16 4 9 0 9 13 3 1 9 2 13 15 15 3 3 13 1 9 9 0 1 9 2 7 3 3 14 1 0 9 1 0 9 2
3 15 3 2
10 0 9 1 9 9 0 9 13 9 2
14 0 9 13 3 9 0 9 1 9 1 0 0 9 2
11 9 11 13 9 1 9 12 9 1 9 2
61 1 9 1 9 13 2 0 9 2 14 12 5 2 2 9 2 12 5 2 2 0 9 2 12 2 12 5 2 2 0 9 2 12 2 12 5 2 2 0 0 9 2 12 2 12 5 2 2 0 0 9 2 12 5 2 7 16 0 9 9 2
18 1 3 0 9 1 0 9 1 0 9 13 9 13 3 3 1 15 2
9 1 9 15 9 13 1 12 5 2
3 9 1 9
12 13 9 0 9 9 1 9 12 7 9 12 2
12 1 12 9 9 15 13 12 9 0 9 11 2
18 1 10 9 13 9 9 12 9 1 9 12 7 12 9 1 9 12 2
9 1 10 9 15 13 13 0 9 2
18 15 13 1 9 0 9 1 11 12 9 2 16 3 1 9 12 9 2
12 0 9 1 9 13 12 5 9 1 0 9 2
17 15 13 1 0 0 9 12 9 7 1 9 9 12 3 12 9 2
23 0 9 9 11 0 1 9 1 9 12 3 13 12 9 1 9 2 3 1 9 12 9 2
28 0 9 13 7 0 9 3 9 2 16 15 7 1 10 9 13 0 9 1 9 1 12 1 12 9 1 9 2
17 9 9 13 0 2 13 11 9 2 9 0 9 9 2 9 11 2
13 1 9 9 13 2 15 4 13 9 1 10 9 2
13 13 3 1 10 9 2 3 3 13 0 9 13 2
10 9 3 13 1 9 3 1 0 9 2
2 9 13
12 0 9 13 3 3 0 16 9 0 1 11 2
10 9 9 1 0 9 13 14 12 9 2
11 7 13 15 13 7 9 2 9 7 9 2
13 1 9 15 9 0 9 13 1 12 9 1 9 2
15 9 1 9 11 3 13 0 9 1 0 0 9 1 15 2
8 16 15 13 9 1 9 9 2
17 3 9 7 9 2 15 15 13 1 10 9 2 15 1 9 13 2
12 0 0 9 13 1 9 0 9 9 9 9 2
9 9 3 13 9 1 0 0 9 2
11 1 12 2 9 12 7 7 10 9 13 2
8 9 9 11 13 0 9 13 2
20 13 15 3 9 13 2 16 10 9 13 3 0 9 2 0 9 7 0 9 2
13 1 10 9 13 9 1 9 1 0 9 7 9 2
13 15 13 2 16 1 9 9 4 13 10 0 9 2
26 9 9 15 7 13 3 13 2 1 1 15 2 16 0 9 3 3 1 9 9 11 13 9 0 9 2
29 13 2 14 7 11 3 1 10 0 9 1 0 7 14 3 0 9 2 13 0 9 16 15 13 1 0 0 9 2
15 3 15 13 9 9 1 9 14 1 12 9 1 9 9 2
20 0 9 7 4 13 1 9 9 0 9 2 15 1 11 13 1 0 1 11 2
28 1 9 15 4 1 0 13 13 2 3 13 9 0 2 16 9 1 9 4 15 13 13 1 0 7 0 9 2
24 1 9 2 16 4 15 0 9 13 1 0 0 9 9 9 2 13 15 9 1 9 0 9 2
36 13 2 14 15 1 9 2 13 4 0 9 13 1 9 0 9 2 3 4 13 13 13 0 12 9 11 2 15 4 13 13 3 0 0 9 2
2 9 2
11 9 9 2 0 1 9 11 1 9 12 2
7 0 9 9 1 9 12 2
7 9 9 9 1 9 12 2
4 0 9 7 15
2 0 11
15 0 9 0 11 2 11 2 13 1 0 7 0 1 9 2
21 16 13 0 9 3 1 9 12 2 13 15 9 9 2 15 13 3 1 0 9 2
20 11 13 3 16 12 9 7 13 0 9 1 12 9 9 1 9 1 12 9 2
24 1 9 9 9 11 11 13 11 1 12 9 1 12 9 0 9 7 3 13 1 12 9 9 2
19 0 9 1 0 9 0 9 13 1 9 11 3 1 0 9 1 0 9 2
16 3 16 3 0 0 0 9 13 13 1 0 9 9 1 9 2
11 1 11 13 11 9 3 3 16 12 9 2
25 3 15 1 11 1 11 13 3 3 3 2 1 9 12 15 9 9 13 14 1 0 12 9 3 2
8 3 11 13 12 9 12 0 2
12 9 9 11 1 11 15 7 13 13 1 12 2
19 1 9 0 9 13 11 9 1 11 9 0 9 0 11 1 9 1 11 2
36 9 2 0 11 2 0 9 2 12 2 12 2 12 12 11 12 2 9 2 2 2 12 2 12 12 12 2 9 2 2 12 2 12 12 12 2
3 9 1 9
18 9 1 9 7 0 9 13 0 9 9 2 10 9 13 9 0 9 2
12 15 4 13 0 9 1 9 7 9 1 11 2
17 9 1 9 1 9 13 0 9 0 9 1 0 9 7 0 9 2
30 1 9 1 0 9 13 3 13 9 7 13 0 9 1 9 12 9 1 9 2 12 9 1 9 7 12 9 1 9 2
11 1 9 9 4 0 13 1 12 0 9 2
28 9 13 0 9 1 11 7 3 1 9 2 0 3 9 1 0 11 7 3 0 9 1 3 0 9 1 11 2
24 9 9 13 1 9 2 0 9 15 13 12 2 2 12 2 9 7 0 9 13 1 9 9 2
6 0 9 13 1 9 2
30 9 2 9 1 9 7 0 9 2 0 12 2 12 12 11 12 2 9 2 7 9 2 2 12 2 12 12 2 12 12
5 1 9 15 9 13
4 0 9 1 9
19 1 9 9 4 1 9 12 13 12 9 12 0 9 2 11 2 1 11 2
21 1 10 9 4 13 12 5 12 9 5 12 5 12 5 2 7 2 3 12 9 2
15 10 9 12 5 13 1 9 0 9 9 3 0 0 9 2
18 9 15 3 3 13 7 9 9 2 15 4 13 1 10 9 1 9 2
21 1 9 12 13 0 9 2 15 13 2 16 9 1 9 12 2 12 15 4 13 2
14 13 4 15 7 7 0 9 2 3 0 9 2 13 2
46 13 4 9 0 9 1 9 2 3 15 0 9 13 2 16 1 0 2 0 9 13 10 9 13 2 7 1 0 2 13 15 9 1 9 2 10 9 9 7 9 13 1 0 11 13 2
18 13 7 13 2 16 1 0 9 13 13 7 1 9 2 7 1 9 2
2 9 2
20 2 13 9 3 3 7 13 15 1 9 13 15 3 2 16 15 1 15 13 2
12 2 1 9 9 1 0 9 13 3 10 9 2
26 9 0 9 2 16 13 2 9 2 1 15 13 13 2 2 3 1 9 0 9 13 13 14 3 0 2
4 11 11 2 11
22 9 0 1 10 9 2 0 1 0 9 9 2 4 3 13 7 3 13 9 12 9 2
10 4 3 13 1 0 9 1 12 9 2
19 13 15 1 15 2 10 9 4 15 1 9 13 7 10 1 15 13 9 2
2 9 9
11 0 9 1 9 13 1 0 9 0 9 2
23 1 9 9 9 2 9 12 3 0 1 0 9 7 15 11 13 10 9 2 1 12 5 2
19 11 1 0 9 13 12 9 2 7 15 13 3 3 3 1 9 1 0 2
12 0 9 9 0 9 1 9 12 13 3 0 2
18 0 9 13 3 1 0 9 12 9 7 10 0 9 9 13 12 9 2
4 2 0 9 2
4 13 15 9 2
6 13 2 15 3 13 2
10 13 15 15 2 16 0 9 13 3 2
8 13 15 0 10 9 0 9 2
9 13 3 1 15 13 9 0 9 2
7 10 9 13 1 10 9 2
2 0 9
17 13 15 13 2 1 10 0 9 13 1 0 9 9 1 0 9 2
4 11 9 2 11
15 13 1 9 9 3 9 2 9 2 9 2 9 7 3 2
53 13 15 9 9 1 9 0 9 2 9 0 9 1 0 9 2 13 15 9 9 0 9 1 12 9 2 13 13 1 9 9 2 13 0 9 2 9 2 9 2 0 9 2 9 2 0 9 2 9 2 9 3 2
16 7 9 13 9 7 13 13 15 0 2 16 9 10 0 9 2
2 11 11
20 9 2 0 12 2 12 12 11 12 2 9 2 2 2 12 2 12 12 12 2
3 9 13 9
25 9 9 2 15 4 1 9 13 0 9 2 3 13 1 15 2 16 4 9 1 10 9 13 0 2
14 9 9 7 1 10 9 13 7 13 9 9 0 9 2
2 3 2
2 11 11
55 9 9 1 9 9 13 3 0 2 13 9 9 11 11 11 2 16 9 2 15 1 15 13 3 9 2 7 3 13 7 3 13 3 0 2 15 1 9 13 1 15 2 16 4 1 15 13 9 0 1 9 7 9 9 2
21 10 9 13 1 0 7 9 9 9 2 15 1 0 12 9 9 11 13 1 9 2
35 3 15 13 11 11 2 1 9 12 13 9 11 1 12 0 9 7 3 13 1 9 3 12 9 2 15 13 1 12 9 7 12 0 9 2
15 7 15 3 9 2 15 0 13 9 9 1 9 9 9 2
51 1 0 9 2 16 13 9 0 9 2 9 1 9 9 2 9 2 9 7 9 2 10 9 1 9 2 9 7 0 9 9 7 7 9 0 9 2 13 9 9 3 9 0 9 2 15 1 15 15 13 2
19 1 1 0 0 9 0 0 9 13 9 1 10 9 7 9 3 16 3 2
24 9 9 13 9 16 0 0 2 13 3 10 9 2 7 1 10 9 13 13 10 9 3 0 2
30 7 16 3 9 11 14 1 12 9 2 3 13 1 9 0 9 9 2 13 9 13 1 9 2 0 9 7 9 9 2
26 1 9 0 9 15 11 13 12 7 12 9 1 9 2 7 15 1 15 2 16 13 1 9 0 9 2
16 3 13 14 9 2 3 13 15 12 9 1 1 0 9 9 2
37 1 0 9 13 1 9 12 9 1 9 7 3 1 9 11 12 13 15 1 9 14 12 9 1 0 9 1 9 2 16 13 1 9 7 0 9 2
17 1 10 9 1 9 11 11 4 9 13 7 1 9 9 1 9 2
25 9 9 15 13 1 9 2 1 15 13 12 9 1 9 9 2 15 13 9 13 14 1 9 9 2
22 1 0 9 1 0 9 13 2 16 9 13 1 0 9 0 9 2 3 3 3 15 2
7 10 9 15 3 3 13 2
26 16 4 9 1 9 0 9 13 16 3 0 2 13 9 11 1 10 9 3 12 0 7 12 0 9 2
11 13 7 0 9 9 0 2 0 0 9 2
20 1 0 9 13 0 9 9 2 9 9 0 9 7 9 0 3 0 0 9 2
18 9 2 11 2 9 2 1 9 2 0 2 2 1 9 12 2 12 2
2 10 9
5 1 9 13 12 9
8 2 9 9 2 12 2 12 2
26 1 0 9 15 1 9 9 1 9 0 9 2 0 9 0 9 2 13 1 0 9 9 7 0 9 2
15 16 13 1 10 9 0 9 2 1 9 13 3 0 9 2
11 12 1 10 9 13 0 9 9 10 9 2
33 16 9 13 0 9 2 0 1 10 0 0 9 13 7 3 0 9 2 15 13 3 9 0 9 7 3 2 13 10 9 10 9 2
21 0 0 9 2 15 13 1 0 9 0 9 2 3 3 13 9 9 9 10 9 2
11 13 15 3 0 9 9 9 1 0 9 2
11 13 3 3 10 9 1 9 7 0 9 2
10 3 15 9 9 13 0 9 0 9 2
5 15 15 3 13 2
13 13 1 9 9 9 0 9 1 9 3 0 9 2
22 1 10 0 9 2 15 3 13 9 2 15 9 10 9 13 16 9 1 9 0 9 2
16 10 9 4 15 13 13 0 9 9 2 9 1 9 9 2 2
13 3 0 2 15 13 9 1 9 9 2 13 9 2
4 11 11 2 11
5 13 15 13 3 0
8 2 9 9 2 12 2 12 2
18 16 4 13 3 0 15 13 2 14 4 9 13 0 9 2 16 13 2
13 7 16 9 15 9 13 2 16 15 3 13 13 2
34 9 13 1 15 2 16 16 15 13 1 10 0 9 14 1 9 2 13 0 9 7 13 3 13 1 9 2 7 15 1 15 0 13 2
16 9 16 9 9 10 9 15 14 13 1 0 9 7 1 15 2
21 13 9 15 13 13 0 9 3 1 9 3 0 9 2 16 3 13 3 0 9 2
24 10 9 2 15 9 13 2 15 7 13 2 16 3 15 1 9 13 2 3 15 1 9 13 2
18 0 4 13 2 16 4 15 9 7 9 3 13 1 0 9 13 3 2
7 3 4 13 9 7 9 2
27 7 16 15 1 10 9 13 2 3 7 3 2 16 13 0 9 2 3 13 3 9 2 15 1 9 13 2
13 9 13 7 13 9 9 2 1 9 15 13 3 2
14 7 1 15 2 15 9 7 0 9 13 2 9 13 2
15 1 9 9 7 1 0 9 15 3 3 13 7 13 15 2
4 15 13 9 2
11 0 9 9 13 14 0 1 12 0 9 2
15 3 0 7 13 2 16 3 15 3 13 9 0 0 9 2
4 11 11 2 11
6 9 1 9 1 0 9
8 2 9 9 2 12 2 12 2
8 3 4 15 13 10 9 9 2
5 13 3 1 9 2
16 13 4 15 2 16 1 9 15 3 3 13 2 7 15 3 2
13 13 1 9 2 15 13 3 0 2 3 13 9 2
21 9 1 9 0 1 9 9 15 15 3 13 7 1 0 9 15 3 14 4 13 2
7 0 0 9 4 3 13 2
7 4 15 13 3 1 9 2
31 13 1 15 13 0 9 2 10 1 9 0 0 9 2 15 1 9 2 0 9 1 0 9 9 2 0 9 3 2 2 2
14 1 15 3 15 15 9 1 9 13 1 0 12 9 2
26 16 13 7 1 0 9 2 7 1 0 9 2 13 2 16 9 1 15 13 7 1 0 0 9 0 2
14 3 0 4 15 3 2 1 0 9 2 13 3 3 2
10 9 15 3 3 13 7 13 0 9 2
4 11 11 2 11
7 9 2 9 2 9 7 15
8 2 9 9 2 12 2 12 2
29 9 2 1 15 15 10 0 0 9 1 0 9 13 13 9 7 9 1 15 0 0 9 2 13 3 1 0 9 2
35 7 16 9 7 9 15 3 3 1 0 9 13 1 0 9 2 13 15 3 1 0 9 10 9 15 2 16 4 13 10 0 2 9 2 2
82 10 9 13 13 7 1 0 9 2 3 1 12 9 13 0 9 0 7 0 1 0 9 2 15 1 9 0 9 13 9 7 9 13 1 9 1 3 0 0 9 2 7 1 0 9 2 3 3 3 1 15 2 13 0 9 2 1 15 15 15 0 0 9 3 16 9 7 9 13 9 2 15 9 15 13 2 7 13 1 15 9 2
19 3 3 13 12 1 9 10 9 2 13 0 9 1 10 9 0 9 0 2
28 9 15 13 9 1 10 2 16 1 0 9 13 9 0 0 9 1 9 9 7 4 15 1 15 13 0 9 2
28 3 3 13 13 9 9 7 9 1 9 9 1 9 7 13 15 1 15 9 0 1 10 9 2 3 9 0 2
41 0 0 9 13 2 16 16 4 3 1 9 0 13 9 7 9 2 13 15 1 10 9 0 9 2 3 9 1 9 2 16 10 0 9 7 13 1 10 9 13 2
19 1 2 9 2 9 7 9 1 0 9 13 7 3 13 16 1 9 0 2
24 1 0 9 1 15 7 10 9 13 9 0 1 9 0 1 9 2 7 15 3 9 9 0 2
7 11 11 2 9 9 0 9
3 9 2 12
9 9 2 9 2 11 9 2 9 12
4 9 9 2 9
10 0 9 2 2 11 12 2 9 2 12
7 0 9 2 2 9 2 14
10 9 2 2 9 2 12 5 12 5 12
6 9 2 2 9 2 12
2 9 2
5 9 1 0 9 2
9 13 13 9 9 1 9 12 9 2
9 12 9 1 9 2 0 9 2 2
8 12 9 9 2 9 9 9 2
11 9 0 9 12 0 9 2 0 9 9 2
8 9 1 9 7 9 1 9 2
2 9 2
5 9 1 0 9 2
6 9 9 7 16 9 2
10 12 9 9 9 13 13 0 9 9 2
3 9 2 12
8 9 2 9 2 11 11 2 12
4 9 9 2 9
10 0 9 2 11 12 2 9 2 2 12
7 0 9 2 9 2 2 14
10 9 2 9 2 2 12 5 12 5 12
6 9 2 9 2 2 12
2 9 2
11 9 0 1 9 7 1 9 13 0 9 2
11 9 1 12 9 2 1 15 12 0 9 2
6 9 9 1 0 9 2
10 0 9 0 0 9 2 9 1 9 2
10 9 9 1 9 9 1 9 0 9 2
16 1 0 9 9 9 1 0 0 9 7 1 9 1 9 9 2
3 0 9 2
3 9 9 2
8 12 9 9 2 12 9 9 2
8 9 12 9 2 0 9 9 2
8 0 9 9 2 9 2 9 2
7 9 12 9 1 12 9 2
4 9 0 9 2
23 9 1 0 9 3 2 1 9 9 1 9 1 0 9 7 9 1 12 9 7 1 9 2
17 9 9 12 2 12 7 9 1 12 5 2 3 9 1 12 5 2
2 9 2
21 0 9 9 2 3 15 0 9 2 3 13 7 9 1 0 9 1 0 0 9 2
3 9 2 12
9 9 2 9 2 11 9 11 2 12
4 9 9 2 9
10 0 9 2 2 11 12 2 9 2 12
10 9 2 2 9 2 12 5 12 5 12
7 9 2 2 9 2 12 12
2 9 2
9 0 9 0 1 9 1 0 9 2
10 15 13 7 10 9 12 9 3 9 2
9 0 9 0 16 1 0 0 9 2
21 1 9 2 16 0 9 13 0 7 1 9 2 3 13 9 11 2 12 0 3 2
2 9 2
15 9 2 15 13 7 1 9 1 9 13 7 13 0 9 2
14 13 15 3 9 2 13 0 9 2 15 3 13 9 2
3 9 2 12
8 9 2 9 2 11 11 2 12
4 9 9 2 9
10 0 9 2 2 11 12 2 9 2 12
7 0 9 2 2 9 2 14
10 9 2 2 9 2 12 5 12 5 12
6 9 2 2 9 2 12
2 9 2
5 9 0 1 9 2
18 9 1 12 9 2 1 15 12 1 0 9 7 12 1 0 0 9 2
6 9 9 3 7 3 2
8 12 9 9 2 12 9 9 2
4 0 9 9 2
5 9 9 1 9 2
10 9 1 12 9 1 9 1 9 9 2
5 9 9 16 9 2
5 9 9 0 9 2
11 9 9 0 0 9 1 0 9 1 9 2
2 9 2
16 9 1 3 0 9 1 9 0 9 2 3 13 13 3 13 2
3 9 2 12
6 9 2 9 2 11 12
4 9 9 2 9
10 0 9 2 11 12 2 9 2 2 12
7 0 9 2 9 2 2 14
10 9 2 9 2 2 12 5 12 5 12
6 9 2 9 2 2 12
2 9 2
12 9 0 1 9 7 1 0 9 1 0 9 2
12 9 9 13 1 3 12 9 7 13 12 9 2
13 0 9 9 13 9 1 12 9 1 0 0 9 2
8 9 1 12 0 9 11 12 2
17 9 12 9 2 1 15 12 1 0 9 7 12 1 0 0 9 2
7 12 9 9 2 0 9 2
18 0 7 3 0 9 9 13 2 16 7 0 9 15 13 1 11 12 2
5 12 0 0 9 2
4 0 9 9 2
8 9 9 1 0 7 0 9 2
16 0 9 1 9 0 9 9 14 1 12 9 7 1 10 9 2
7 9 1 9 7 9 9 2
6 9 9 9 9 9 2
2 9 2
10 9 1 0 9 1 0 7 0 9 2
11 13 13 1 9 1 0 9 1 9 9 2
3 9 2 12
9 9 2 9 2 11 11 11 2 12
5 9 9 2 9 9
10 0 9 2 11 12 2 9 2 2 12
7 0 9 2 9 2 2 14
10 9 2 9 2 2 12 5 12 5 12
6 9 2 9 2 2 12
2 9 2
10 9 0 1 9 1 9 1 9 9 2
7 12 9 9 13 12 9 2
6 13 0 7 0 9 2
13 9 9 1 12 9 1 9 9 1 0 12 9 2
17 0 9 9 9 2 9 1 9 0 9 1 0 9 1 9 9 2
10 0 9 12 9 2 0 9 12 9 2
6 0 9 0 0 9 2
3 0 9 2
8 9 0 1 12 9 11 12 2
7 0 9 12 5 12 9 2
8 9 9 9 1 9 0 9 2
11 0 9 9 1 12 9 7 1 9 9 2
14 0 9 9 0 9 1 0 9 2 7 1 9 9 2
9 0 9 2 9 2 1 9 9 2
6 12 0 9 1 9 2
8 0 9 1 9 9 0 9 2
2 9 2
25 0 0 9 0 9 7 3 0 9 7 9 9 13 10 9 1 9 3 0 1 0 9 0 9 2
3 9 2 12
8 9 2 9 2 11 11 12 9
4 9 9 2 9
10 0 9 2 11 12 2 9 2 2 12
7 0 9 2 9 2 2 14
10 9 2 9 2 2 12 5 12 5 12
6 9 2 9 2 2 12
2 9 2
8 9 1 9 1 12 9 9 2
8 9 1 12 9 7 9 9 2
12 1 15 12 1 0 9 2 12 1 0 9 2
10 0 9 15 1 0 9 13 1 9 2
19 0 9 9 7 9 9 1 9 0 9 13 1 9 9 7 9 0 9 2
6 0 9 9 0 9 2
10 0 9 7 3 9 14 1 12 9 2
3 0 9 2
8 9 9 0 9 1 9 9 2
4 9 1 9 2
6 0 9 13 0 9 2
4 12 9 9 2
4 0 9 9 2
6 0 9 1 0 9 2
7 0 9 9 1 12 9 2
8 9 0 9 9 1 0 9 2
2 9 2
20 9 1 3 0 9 1 0 9 13 9 0 9 1 9 2 15 3 13 9 2
3 9 2 12
7 9 2 9 2 11 9 12
4 9 9 2 9
10 0 9 2 11 12 2 9 2 2 2
7 0 9 2 9 2 2 14
10 9 2 9 2 2 12 5 12 5 12
6 9 2 9 2 2 12
2 9 2
11 9 0 1 9 7 1 9 9 0 9 2
20 1 9 2 16 13 9 1 0 9 2 3 13 1 9 2 3 13 0 9 2
10 1 10 9 0 0 9 13 10 9 2
16 12 0 9 2 1 15 12 1 0 9 2 9 1 0 9 2
7 0 0 9 0 0 9 2
12 9 9 0 9 7 9 9 7 1 10 9 2
8 12 9 9 7 12 9 9 2
14 9 9 2 12 9 7 12 9 1 9 9 7 9 2
6 0 9 9 1 9 2
2 9 2
20 9 3 3 0 9 2 0 1 9 0 9 7 1 9 2 15 13 9 3 2
4 9 2 0 9
1 9
15 9 0 9 13 1 9 9 2 9 1 0 9 0 9 2
21 10 9 13 1 11 0 1 9 12 1 9 9 11 11 16 9 1 9 0 9 2
10 0 0 9 4 13 9 1 9 12 2
6 13 3 0 9 9 2
9 3 13 12 9 9 12 9 9 2
7 0 9 13 1 3 0 2
11 1 9 11 15 3 9 9 1 9 13 2
23 16 1 9 12 15 13 9 1 0 12 9 2 9 0 9 15 13 1 12 9 1 9 2
7 9 1 11 13 3 0 2
24 1 9 15 3 0 9 13 1 12 9 2 1 0 9 15 13 12 9 7 1 9 12 9 2
14 0 9 13 1 0 9 2 3 15 13 1 12 9 2
51 0 9 3 13 1 2 2 12 9 9 1 12 9 2 2 12 9 9 1 12 2 2 12 9 0 9 2 12 9 2 1 12 9 2 2 9 9 11 14 12 9 2 2 12 9 0 9 14 12 9 2
12 1 12 9 3 13 0 1 9 13 3 15 2
18 3 0 9 13 1 12 9 2 9 1 9 1 11 1 12 9 3 2
4 9 1 9 2
11 9 9 9 1 9 1 9 12 2 12 2
4 7 9 13 9
7 9 9 13 15 9 0 9
14 13 9 2 1 10 9 15 0 13 3 10 0 9 2
18 15 3 3 15 2 16 0 9 1 10 9 13 13 1 9 3 9 2
6 13 15 7 1 9 2
21 12 1 10 9 1 9 13 7 11 11 2 9 9 9 9 1 11 1 11 12 2
23 9 1 15 13 1 15 2 10 0 9 13 2 10 9 2 16 9 2 13 1 10 9 2
13 2 13 15 1 15 2 16 13 3 13 10 9 2
14 15 15 1 15 2 7 1 9 1 9 3 2 13 2
4 13 14 9 2
8 13 0 9 1 9 7 3 2
20 16 13 15 1 9 2 13 15 0 7 13 15 1 0 2 7 13 3 13 2
8 13 4 15 13 14 0 9 2
8 13 15 2 16 9 13 15 2
12 1 0 9 4 13 13 0 9 9 7 9 2
13 13 9 1 0 9 7 1 9 0 1 9 9 2
21 10 9 7 0 0 9 1 10 9 13 13 2 3 7 1 9 2 16 1 15 2
4 15 13 9 2
11 1 9 15 13 3 2 16 9 1 15 2
15 2 3 4 15 3 13 2 15 3 13 13 9 0 9 2
21 9 9 2 15 1 9 2 1 9 13 15 3 3 1 12 1 9 1 0 9 2
11 15 1 15 1 9 13 0 9 1 9 2
6 13 15 10 9 9 2
12 1 10 9 7 10 0 9 13 3 3 0 2
10 16 0 9 2 13 7 15 0 9 2
10 15 7 13 13 0 1 9 1 9 2
11 2 13 4 1 0 9 2 15 15 13 2
20 9 4 13 13 0 2 9 13 13 2 15 15 1 15 13 7 15 4 13 2
22 16 9 13 2 13 1 9 2 16 4 15 13 2 3 3 1 10 9 13 13 13 2
15 13 1 15 2 16 4 3 13 9 7 3 9 13 9 2
6 15 15 1 15 13 2
18 2 1 10 9 15 10 9 1 0 9 0 9 13 1 9 10 9 2
12 9 2 3 15 15 13 3 2 15 3 13 2
16 9 13 1 9 2 16 4 13 9 2 1 15 3 13 13 2
13 1 9 15 15 3 3 13 13 7 13 15 0 2
9 9 3 13 9 9 2 15 13 2
13 1 0 9 2 3 13 0 2 9 2 1 9 2
6 9 9 13 0 9 2
13 1 15 13 0 0 9 13 3 3 3 12 9 2
7 3 13 10 9 7 9 2
30 13 15 15 3 0 2 16 13 2 14 13 9 2 13 13 0 9 9 2 7 15 3 3 1 0 2 0 2 9 2
19 1 10 0 9 2 15 13 0 9 9 2 13 9 1 10 9 7 9 2
7 2 15 15 13 1 9 2
17 13 2 16 4 9 7 9 15 9 1 9 13 0 9 7 9 2
11 7 15 13 1 15 9 7 1 9 9 2
41 10 9 13 1 9 7 3 0 2 9 15 3 15 13 2 13 1 0 9 7 1 15 2 16 13 16 9 2 0 9 7 3 16 0 9 2 15 10 9 13 2
9 1 15 12 1 0 13 15 13 2
18 1 0 9 13 7 0 9 7 9 15 2 9 2 9 7 0 9 2
17 13 9 10 9 13 7 0 9 9 2 15 13 1 9 7 3 2
19 13 15 9 7 9 13 10 9 1 15 7 13 13 1 0 9 9 0 2
10 15 13 9 9 2 15 10 9 13 2
10 13 15 15 3 7 0 9 10 9 2
5 11 11 2 11 11
4 9 1 9 2
4 9 1 9 2
23 7 3 13 13 9 2 15 10 9 7 9 13 10 9 1 0 9 7 0 9 0 9 2
3 9 1 9
8 0 9 9 1 0 9 1 11
22 0 9 7 9 13 1 0 0 9 7 3 1 0 9 2 15 13 1 9 0 9 2
27 13 3 0 2 16 4 15 13 2 16 1 0 9 1 0 9 9 2 9 7 9 1 9 15 13 3 2
19 3 1 0 9 7 0 0 9 13 13 7 9 9 2 3 16 0 9 2
17 10 9 3 13 9 2 13 9 9 1 0 7 0 9 1 11 2
9 0 9 13 12 0 9 0 9 2
37 0 9 2 3 9 2 0 9 7 0 9 2 13 12 5 2 9 0 7 0 9 12 5 2 9 9 7 0 9 12 5 7 9 12 5 9 2
16 1 12 5 4 13 9 0 9 7 12 5 13 0 0 9 2
7 1 9 9 13 0 9 2
7 9 10 9 13 3 13 2
42 1 10 9 15 13 1 9 2 16 13 0 9 0 9 2 0 9 2 1 15 13 0 9 2 7 0 9 0 0 9 2 9 2 7 3 9 2 9 7 0 9 2
21 10 9 15 3 1 10 9 13 2 16 10 0 9 13 0 9 7 13 0 9 2
8 0 9 13 3 9 7 9 2
3 9 15 13
25 1 9 13 9 7 9 3 13 10 0 9 2 3 13 9 7 9 7 13 0 9 1 9 3 2
16 9 13 13 10 0 9 2 13 9 2 13 9 9 7 9 2
10 0 9 13 3 13 9 7 0 9 2
24 9 1 0 9 13 3 0 2 7 2 3 13 9 1 11 7 11 2 0 7 3 15 13 2
29 9 1 11 13 2 16 9 15 13 13 1 9 10 9 0 9 2 0 9 7 9 0 9 1 9 7 10 9 2
6 0 9 13 0 9 2
14 1 0 9 9 13 1 11 9 9 0 9 1 9 2
14 7 3 13 13 2 16 0 0 2 9 13 7 0 2
3 13 15 9
56 9 9 7 0 9 15 13 1 9 2 16 13 0 3 1 9 0 9 1 0 9 13 9 9 10 9 2 13 15 1 9 1 0 9 2 0 9 2 0 9 2 9 2 7 13 15 13 15 0 9 7 13 0 0 9 2
25 7 13 1 0 9 1 0 9 1 11 2 1 9 9 0 9 2 13 0 0 9 9 1 9 2
7 13 13 1 12 0 9 2
8 1 0 13 9 7 0 9 2
22 1 0 9 13 0 9 0 9 2 0 9 2 13 15 1 9 7 0 9 0 9 2
7 0 9 13 7 13 0 2
32 1 0 15 9 13 1 0 9 2 0 9 0 2 9 2 9 2 9 7 0 0 9 0 1 9 9 7 1 9 1 9 2
17 13 4 3 9 7 0 9 7 9 13 13 1 0 9 10 9 2
16 1 0 9 4 13 0 9 7 1 9 13 7 1 0 9 2
14 9 7 9 15 13 13 1 10 0 9 7 10 9 2
12 16 13 13 15 2 13 13 9 15 15 9 2
18 3 0 13 7 13 3 0 0 9 7 1 9 0 9 13 0 9 2
24 0 13 13 15 0 9 3 2 16 4 15 1 15 13 7 0 9 1 0 9 7 0 9 2
2 11 11
16 2 9 2 0 9 1 11 2 0 12 2 12 12 11 2 2
4 9 1 9 2
3 0 9 2
11 0 0 9 7 9 13 9 13 1 9 2
7 9 15 13 10 9 13 2
1 9
7 9 11 11 1 9 9 2
19 1 10 9 1 11 13 9 9 1 12 9 7 12 9 9 1 12 9 2
12 7 1 12 9 7 0 9 9 13 0 9 2
35 9 1 9 2 0 9 2 9 0 9 2 4 13 2 16 1 9 4 13 9 0 9 12 2 3 12 9 1 0 9 9 9 12 9 2
6 15 4 9 13 13 2
13 9 0 9 1 0 9 3 13 1 9 10 9 2
3 0 11 12
32 11 11 2 12 2 0 0 9 9 2 9 2 0 9 2 9 2 0 9 7 9 1 10 9 2 12 2 2 12 2 12 2
25 11 2 11 2 11 11 2 12 2 9 9 2 9 7 0 0 9 2 12 2 2 12 2 12 2
21 0 2 11 2 11 2 9 2 2 0 0 9 9 2 12 2 2 12 2 12 2
21 11 2 11 2 12 2 0 0 9 0 9 7 9 2 12 2 2 12 2 12 2
16 11 2 12 2 0 9 1 9 2 12 2 2 12 2 12 2
18 12 2 9 0 0 9 0 1 0 9 2 12 2 2 12 2 12 2
23 11 2 12 2 0 0 9 1 0 7 0 9 1 0 9 2 12 2 2 12 2 12 2
23 9 2 12 2 0 0 9 1 0 9 2 0 9 7 9 2 12 2 2 12 2 12 2
13 11 2 0 9 9 2 12 2 2 12 2 12 2
22 11 2 12 2 0 9 0 7 0 9 1 0 0 9 2 12 2 2 12 2 12 2
21 0 2 11 2 11 2 9 2 2 0 0 9 9 2 12 2 2 12 2 12 2
22 11 2 11 2 12 2 0 0 9 0 9 7 9 12 2 12 2 2 12 2 12 2
24 11 2 11 2 0 0 9 9 2 9 2 0 9 7 0 9 2 12 2 2 12 2 12 2
24 11 2 0 0 9 9 1 0 9 2 9 2 9 7 0 9 2 12 2 2 12 2 12 2
19 9 12 11 2 12 2 0 0 9 0 9 2 12 2 2 12 2 12 2
19 11 11 2 9 1 9 0 9 0 0 9 2 12 2 2 12 2 12 2
30 11 2 12 2 0 0 9 9 2 9 2 9 2 9 7 9 1 0 0 7 0 9 2 12 2 2 12 2 12 2
27 11 11 2 12 2 0 0 9 2 9 2 9 2 9 2 0 9 7 9 2 12 2 2 12 2 12 2
29 11 2 12 2 0 0 9 0 9 1 9 2 9 2 9 7 9 9 1 0 9 2 12 2 2 12 2 12 2
20 11 2 12 2 0 0 9 0 0 9 7 9 2 12 2 2 12 2 12 2
2 12 2
23 11 5 11 2 0 9 1 9 1 9 0 0 9 2 12 2 12 2 2 12 2 12 2
53 9 2 9 11 11 11 2 11 5 11 2 9 2 9 2 0 2 2 9 2 11 11 2 0 9 12 2 12 12 11 2 9 2 2 2 12 2 12 12 2 12 2 9 2 2 9 2 2 12 2 12 12 2
4 9 2 9 9
6 9 1 12 2 9 9
18 9 9 13 1 10 9 1 9 2 16 4 15 1 15 9 13 13 2
15 9 1 0 9 13 1 9 9 7 13 9 2 9 9 2
8 9 13 1 9 1 0 9 2
1 9
3 9 0 9
27 9 9 0 9 2 15 13 9 11 2 13 9 0 9 9 0 9 11 11 2 11 7 11 11 2 11 2
44 13 0 9 2 7 3 7 3 13 9 0 9 2 7 2 0 9 9 1 9 9 2 9 7 9 9 2 9 7 9 9 7 3 7 10 9 2 9 9 7 0 9 9 2
28 13 15 7 9 3 0 2 9 7 9 0 9 7 0 9 1 9 2 9 0 9 2 9 7 9 0 9 2
7 0 9 13 13 0 9 2
10 9 13 3 0 9 0 9 0 9 2
27 9 13 13 3 1 9 0 9 2 0 9 2 9 0 9 2 3 16 1 9 9 1 0 7 0 9 2
37 2 9 2 11 2 1 9 12 2 12 12 11 12 2 9 2 2 2 12 2 12 2 2 12 2 12 12 2 9 2 2 12 2 12 12 2 2
2 0 9
8 9 1 9 13 3 16 14 9
24 0 0 9 12 2 12 2 2 12 2 12 2 12 2 15 4 13 1 9 9 9 2 9 2
20 13 3 10 9 1 0 7 0 9 1 11 13 10 9 1 0 7 0 9 2
18 0 9 1 0 9 13 1 9 3 0 1 11 2 1 11 7 11 2
12 0 0 9 9 13 0 9 0 7 0 11 2
6 15 15 3 4 13 2
32 3 9 7 9 2 16 0 9 2 9 2 0 9 2 0 9 2 9 2 9 2 9 2 0 9 2 0 9 2 7 3 2
10 15 13 3 0 9 1 9 1 15 2
5 7 15 13 0 2
24 0 1 9 11 2 11 13 0 9 1 9 2 9 2 0 9 2 9 2 9 2 9 9 2
41 13 15 2 16 9 9 15 4 13 3 1 9 7 0 9 9 0 9 3 1 0 0 9 2 15 13 0 9 7 9 2 7 0 9 1 10 9 1 0 9 2
14 9 1 11 4 15 13 13 16 9 3 1 0 9 2
8 0 9 13 1 9 13 9 2
19 1 9 13 0 9 2 0 9 7 0 9 1 9 12 9 2 9 12 2
14 9 0 0 9 15 3 13 1 12 9 2 9 12 2
23 1 11 15 13 13 3 12 9 2 16 1 12 13 9 14 12 9 12 1 9 0 9 2
9 1 9 13 7 9 1 9 9 2
8 9 9 7 13 13 14 0 2
12 7 1 9 13 1 9 0 9 9 2 9 2
21 0 9 7 13 10 9 7 9 7 1 11 2 3 13 0 0 9 1 0 9 2
2 11 9
31 9 2 11 2 9 12 2 9 12 2 12 12 11 12 2 9 2 2 2 12 2 12 12 12 12 2 12 12 12 12 2
1 9
5 9 2 9 2 9
22 2 9 2 9 2 9 2 0 9 0 9 2 9 9 2 0 9 9 1 0 9 2
31 9 2 12 2 2 12 2 12 2 2 12 2 2 12 2 12 2 12 2 9 12 2 12 2 7 12 2 12 2 12 2
34 9 2 11 2 9 2 0 12 2 12 12 11 12 2 9 11 2 9 2 2 2 12 2 12 12 2 9 2 2 12 2 12 12 2
33 2 9 2 0 9 9 9 2 0 9 0 9 2 9 9 1 0 7 0 9 2 9 2 9 2 9 2 9 9 7 0 9 2
8 9 2 12 2 12 2 12 2
34 9 2 11 2 9 2 0 12 2 12 12 11 12 2 9 11 2 9 2 2 2 12 2 12 12 2 9 2 2 12 2 12 12 2
27 2 9 2 0 9 9 2 0 9 1 0 9 0 9 2 9 2 9 2 9 2 9 9 2 9 3 2
11 9 2 12 2 2 12 2 12 2 12 2
43 9 2 11 2 11 2 9 2 2 9 2 9 2 0 2 2 0 9 11 2 0 12 2 2 12 2 12 2 12 12 11 12 2 9 2 5 9 2 2 12 2 12 2
9 2 9 2 9 2 0 9 9 2
38 9 2 12 2 2 12 2 12 2 2 12 2 2 12 2 12 2 2 12 2 2 12 2 12 2 12 2 12 0 9 2 9 0 9 1 11 2 2
38 9 2 9 9 9 2 0 9 2 9 2 11 11 2 1 9 12 2 12 12 11 12 2 9 2 2 2 12 2 12 2 9 2 2 12 2 12 2
24 2 9 2 9 7 9 9 2 0 9 9 0 9 0 1 9 2 9 9 2 0 9 3 2
8 9 2 12 2 12 2 12 2
37 9 2 11 2 9 2 11 11 2 0 12 2 12 12 11 12 2 9 2 2 2 12 2 12 12 2 9 2 5 9 2 2 12 2 12 12 2
28 2 9 2 0 9 1 0 9 2 9 9 7 0 2 15 0 9 13 9 9 7 0 9 1 9 1 9 2
18 9 2 12 5 3 9 2 9 1 0 0 9 1 0 9 1 11 2
36 9 2 11 2 11 2 9 2 9 2 0 2 2 11 12 2 12 12 11 12 2 9 2 2 2 12 2 12 2 12 2 12 2 9 12 2
11 2 9 2 9 1 9 0 9 3 9 2
9 9 2 9 12 2 7 9 12 2
25 9 2 9 9 11 11 2 0 12 2 12 12 11 11 2 9 2 5 9 2 2 12 2 12 2
24 2 9 2 0 9 11 1 9 2 0 9 7 9 2 0 9 2 9 2 9 2 9 9 2
18 9 2 12 2 12 2 2 12 2 12 2 2 12 2 12 2 12 2
31 9 2 9 2 11 2 0 12 2 12 12 11 11 2 9 2 2 2 12 2 12 12 2 9 2 2 12 2 12 12 2
12 2 9 2 9 15 13 7 9 1 0 9 2
11 9 2 12 2 2 12 2 12 2 12 2
32 9 2 11 2 9 2 9 2 0 2 2 0 12 2 12 12 11 12 2 9 2 5 9 2 2 12 2 12 12 2 12 2
37 2 9 2 9 7 15 2 9 9 9 1 9 1 9 12 2 9 1 0 9 7 0 9 1 9 7 9 9 2 9 9 2 9 9 2 9 2
32 9 2 11 2 9 2 9 2 0 2 2 0 12 2 12 12 11 12 2 9 2 5 9 2 2 12 2 12 12 2 12 2
52 2 9 2 0 9 2 9 1 9 1 0 9 2 0 9 9 3 3 0 2 9 9 9 1 9 1 0 9 2 9 1 0 2 7 0 2 9 7 9 1 9 1 0 9 2 9 1 9 7 0 9 2
31 9 2 12 2 2 12 2 12 2 2 12 2 12 2 2 12 2 12 2 2 12 2 12 2 2 12 2 12 2 12 2
32 9 2 11 2 9 2 9 2 0 2 2 0 12 2 12 12 11 12 2 9 2 5 9 2 2 12 2 12 12 2 12 2
48 2 9 2 9 9 2 9 9 7 9 0 9 1 9 2 9 1 9 2 9 0 9 2 9 0 9 2 0 9 2 9 2 0 9 2 9 7 9 2 0 9 2 9 7 9 1 9 2
32 9 2 11 2 9 2 9 2 0 2 2 0 12 2 12 12 11 12 2 9 2 5 9 2 2 12 2 12 12 2 12 2
29 2 9 2 0 9 2 3 3 13 2 9 9 1 9 2 9 1 9 2 9 9 2 0 9 2 9 0 9 2
2 12 2
32 9 2 11 2 9 2 9 2 0 2 2 0 12 2 12 12 11 12 2 9 2 5 9 2 2 12 2 12 12 2 12 2
63 2 9 2 9 9 12 2 2 9 12 9 2 0 9 7 0 2 9 2 9 7 9 0 2 9 2 9 9 9 2 0 9 9 2 9 0 9 2 3 13 0 9 1 9 2 0 9 9 9 2 0 9 9 7 0 9 2 9 9 1 9 9 2
32 9 2 11 2 9 2 9 2 0 2 2 0 12 2 12 12 11 12 2 9 2 5 9 2 2 12 2 12 12 2 12 2
57 2 9 2 9 1 9 2 11 9 1 9 2 11 11 2 9 2 9 12 2 11 12 2 9 2 11 12 2 12 2 12 1 11 2 9 2 0 2 11 1 9 2 9 2 11 12 2 9 12 2 9 12 2 9 2 0 2
32 9 2 11 2 9 2 9 2 0 2 2 0 12 2 12 12 11 12 2 9 2 5 9 2 2 12 2 12 12 2 12 2
6 9 1 9 1 12 9
9 1 9 9 1 9 13 9 0 9
19 13 4 15 2 16 13 0 9 3 2 16 4 13 0 9 2 13 0 2
7 9 7 9 0 9 13 2
15 9 9 11 2 15 15 1 15 13 2 7 13 15 0 2
23 16 3 13 15 9 1 9 2 13 0 9 1 9 2 16 13 1 9 2 3 1 9 2
8 3 0 13 9 1 10 9 2
6 13 13 14 12 9 2
2 11 11
21 0 9 9 15 13 1 9 2 0 2 16 13 0 0 9 1 9 9 7 9 2
2 12 2
2 0 9
13 3 9 10 9 13 13 1 9 9 0 9 11 2
9 1 9 0 9 13 1 9 9 2
24 0 1 9 13 3 0 0 9 2 0 9 11 2 7 1 9 9 7 9 9 9 9 11 2
14 10 9 15 13 7 0 9 0 9 1 9 9 9 2
8 0 1 9 13 0 9 11 2
15 13 1 3 0 9 2 1 15 3 12 13 9 0 9 2
17 13 3 13 15 0 2 13 11 0 2 9 9 2 1 9 2 2
5 0 9 3 13 2
2 12 2
2 0 9
16 16 9 10 9 13 2 13 0 9 2 1 15 13 9 3 2
18 13 15 13 9 2 16 4 13 2 16 1 10 9 13 9 7 3 2
39 13 2 16 0 9 13 9 1 9 2 15 13 2 9 13 2 13 9 2 13 9 1 9 1 0 9 2 0 9 13 9 12 9 9 2 2 13 9 2
11 0 0 9 1 9 13 9 7 3 13 2
18 1 9 0 9 13 0 9 2 13 0 9 7 9 1 9 9 2 2
8 1 0 9 13 3 14 9 2
66 3 2 16 9 9 0 9 1 9 9 13 0 2 13 3 14 0 9 7 13 9 1 9 9 2 2 9 1 0 9 13 0 9 9 2 15 4 1 9 13 13 0 9 1 9 9 2 12 9 2 1 0 9 7 14 15 13 1 9 2 3 13 15 1 9 2
2 0 9
33 9 15 13 1 10 9 2 16 9 1 9 13 3 9 2 7 3 9 2 7 15 7 1 9 0 9 2 3 3 0 9 13 2
4 13 12 9 2
16 12 2 0 9 1 0 9 2 1 11 2 3 15 15 13 2
14 7 3 1 11 4 13 0 0 9 2 13 11 0 2
16 16 4 13 2 15 15 13 2 3 4 15 1 9 7 13 2
7 3 13 0 9 1 9 2
5 9 13 9 9 2
11 13 4 0 9 2 0 9 2 0 9 2
10 7 10 9 13 3 0 16 1 9 2
14 15 7 13 0 16 9 7 9 15 3 13 1 9 2
15 16 4 13 9 13 2 13 4 1 9 2 13 11 0 2
4 15 13 15 2
9 13 9 1 9 7 9 13 0 2
13 1 1 12 0 9 9 7 13 13 1 9 3 2
19 0 9 4 15 13 13 0 9 2 3 13 1 9 2 7 3 1 9 2
15 1 9 2 16 15 13 2 13 1 9 2 10 13 9 2
6 3 15 15 13 3 2
24 9 13 9 1 9 16 9 1 15 2 16 13 0 13 9 2 16 1 9 13 9 0 9 2
6 13 3 3 0 9 2
39 1 1 15 2 16 9 1 9 13 1 9 9 9 12 2 13 15 9 1 0 9 2 16 13 4 13 1 9 7 14 1 9 1 9 13 1 9 12 2
12 7 9 13 1 9 13 3 1 9 9 12 2
16 0 9 13 1 0 13 15 10 9 14 1 0 9 1 11 2
22 13 15 0 2 7 16 4 13 0 9 2 3 4 10 9 13 2 13 15 11 0 2
1 2
25 1 9 1 9 7 9 13 9 9 12 2 12 9 2 2 1 9 1 9 1 9 12 2 9 2
8 9 9 1 11 7 13 0 2
20 1 9 11 1 0 9 11 2 1 15 7 9 11 13 2 13 3 0 9 2
12 3 13 9 13 2 16 13 1 9 7 9 2
14 3 13 2 13 2 14 15 10 9 2 13 1 9 2
20 9 2 9 11 2 9 11 2 0 12 2 9 2 2 2 12 2 12 12 2
5 9 1 9 2 2
4 0 0 9 2
9 3 9 2 3 9 2 3 9 2
5 0 9 13 2 13
10 0 9 0 9 15 13 12 2 9 12
25 0 9 2 9 0 9 1 0 9 13 1 9 9 12 2 0 10 9 13 12 2 9 9 12 2
9 9 12 15 13 0 9 0 9 2
11 3 15 13 9 3 1 12 9 2 9 2
13 1 15 13 14 12 9 2 9 1 9 1 9 2
7 15 15 3 3 13 13 2
2 11 11
9 9 9 12 13 13 0 0 9 2
12 1 11 4 12 2 9 12 3 13 10 9 2
25 13 1 15 7 9 2 15 13 10 9 2 7 1 9 1 9 0 9 7 10 9 15 13 9 2
34 13 15 14 1 12 7 12 0 9 2 7 13 15 2 16 4 4 15 13 2 13 11 11 2 9 9 1 9 0 9 7 10 9 2
2 9 3
11 10 9 13 9 1 9 9 12 7 12 2
16 1 9 12 0 9 13 2 15 15 13 1 0 9 9 9 2
17 1 12 2 9 9 12 13 1 10 9 14 1 12 1 12 9 2
36 1 1 9 9 10 0 9 1 9 9 1 9 0 9 7 10 9 11 1 9 0 9 11 7 1 0 9 11 9 9 12 13 10 9 3 2
9 1 0 12 9 13 3 14 12 2
57 1 0 9 4 9 3 13 9 1 0 9 1 12 0 9 2 14 12 9 2 2 9 9 1 9 2 7 13 16 0 9 9 1 9 0 9 7 10 9 1 0 9 2 0 9 2 9 1 9 12 2 12 9 2 7 3 2
14 13 15 3 3 1 9 12 9 1 9 9 1 9 2
11 13 2 14 9 1 9 2 13 15 13 2
25 13 15 13 7 0 9 2 0 9 2 9 1 9 2 0 9 2 2 7 3 3 1 9 9 2
39 9 13 9 7 1 15 2 16 4 15 13 1 9 1 0 0 9 12 9 12 2 12 9 2 2 15 13 2 16 13 9 1 9 13 14 1 9 9 2
8 3 15 9 13 1 0 9 2
18 3 1 9 9 4 13 1 12 9 2 3 15 4 10 9 3 13 2
21 1 15 13 7 3 13 9 1 10 9 2 16 9 1 9 13 13 10 0 9 2
16 3 13 1 9 2 16 9 13 0 9 9 2 3 0 9 2
10 12 1 0 9 9 13 9 15 9 2
18 10 9 4 13 4 13 1 0 9 2 15 13 3 0 9 1 9 2
11 9 2 1 15 9 13 2 13 0 9 2
7 3 15 15 3 3 13 2
10 3 3 0 9 13 1 9 0 9 2
1 9
17 15 9 0 0 9 15 13 1 9 1 9 0 9 7 10 9 2
21 3 4 1 12 2 12 2 12 13 12 9 1 12 9 9 2 13 15 14 12 2
24 0 9 1 15 2 12 9 9 2 13 13 1 9 7 9 13 1 9 0 9 9 1 9 2
17 12 1 0 9 13 0 0 9 9 2 13 1 12 9 9 2 2
47 3 0 0 9 15 4 3 13 9 1 9 9 9 1 9 2 7 2 13 2 14 0 2 9 1 9 9 1 9 12 9 12 2 12 9 2 2 3 15 13 1 9 2 3 3 13 2
10 15 7 1 9 2 1 15 15 13 2
8 1 11 11 13 10 9 10 2
39 16 15 13 1 0 9 2 13 15 1 0 9 9 1 9 2 7 4 2 14 13 0 9 2 13 1 12 5 0 9 2 15 3 13 12 5 0 9 2
2 0 9
7 3 15 13 3 0 9 2
6 9 15 13 0 9 2
12 16 15 13 2 7 13 3 2 13 15 9 2
12 9 15 7 3 13 2 16 0 9 3 13 2
25 13 12 9 2 13 11 11 2 9 9 9 9 7 9 9 1 9 1 9 0 9 7 10 9 2
30 7 15 13 9 1 9 7 0 9 13 1 9 13 7 13 0 9 2 1 9 1 9 12 9 9 12 2 12 9 2
35 13 2 14 15 1 9 2 7 3 13 10 9 2 13 1 9 0 9 2 1 15 13 9 13 9 2 1 9 12 9 12 2 12 2 2
16 15 2 15 13 2 7 13 3 0 0 9 2 13 0 9 2
27 16 13 9 2 16 13 1 9 9 2 13 4 10 9 13 9 14 1 12 5 0 9 2 14 0 2 2
18 1 0 9 3 9 1 9 0 9 7 10 9 13 7 13 0 9 2
27 9 15 13 9 2 15 13 3 2 7 16 1 15 13 2 3 15 15 1 15 13 0 9 1 9 9 2
16 1 9 12 9 12 2 12 9 2 13 10 9 13 3 9 2
44 0 9 13 3 1 15 2 16 15 9 2 13 2 13 9 0 7 3 1 9 9 12 2 12 9 2 2 7 16 9 13 1 9 9 2 1 15 4 3 13 2 15 13 2
18 1 0 9 13 3 0 9 0 9 2 15 4 13 1 0 9 9 2
22 3 15 13 9 0 0 9 9 1 9 2 13 3 13 9 2 15 4 3 3 13 2
27 13 2 14 15 1 9 1 12 9 1 9 9 2 13 4 13 0 9 2 15 4 13 9 9 1 9 2
16 3 0 2 3 0 13 2 16 13 9 7 13 1 0 9 2
14 3 4 13 0 9 7 9 7 13 13 1 0 9 2
22 16 15 15 13 3 2 13 9 13 1 0 9 7 13 1 9 2 16 4 13 9 2
2 9 13
8 9 0 9 13 14 1 9 2
7 3 9 9 13 10 9 2
12 16 9 13 2 13 15 9 13 1 0 9 2
16 13 15 13 2 16 9 9 13 1 9 0 9 1 15 0 2
7 3 13 2 16 13 3 2
9 0 15 13 2 16 1 15 13 2
12 3 13 13 1 10 0 9 2 13 11 11 2
25 13 3 3 9 0 1 9 2 13 1 9 0 9 1 12 7 12 1 12 9 2 7 4 13 2
9 13 3 3 0 9 2 13 0 2
6 0 9 13 0 9 2
34 16 4 15 7 9 9 13 2 13 15 9 2 13 15 1 0 9 13 1 9 2 0 1 15 4 13 1 0 9 2 13 11 11 2
27 13 7 2 16 1 9 14 1 12 5 7 1 9 1 3 3 12 5 13 1 9 15 2 15 15 13 2
4 0 9 13 2
12 16 0 9 13 10 9 2 1 15 15 13 2
10 12 2 9 12 15 15 7 13 0 2
2 9 9
12 13 0 2 16 4 15 0 9 13 9 9 2
23 11 9 13 9 1 9 0 11 2 16 4 13 13 15 9 2 15 1 9 0 11 13 2
17 0 9 9 13 13 1 9 0 0 9 7 0 3 13 0 9 2
16 13 15 1 9 0 9 9 2 0 9 9 2 9 1 9 2
11 9 4 3 13 9 9 2 15 13 9 2
25 9 2 9 1 9 0 11 2 9 9 12 2 12 12 11 2 9 2 7 9 2 2 12 2 12
1 9
37 1 0 7 0 0 9 15 0 9 13 3 3 13 2 16 4 15 3 13 1 0 3 0 0 9 1 0 9 9 7 15 2 15 1 15 13 2
23 13 15 2 16 10 9 1 15 13 13 9 2 15 13 0 9 1 0 0 9 7 9 2
22 15 2 16 0 7 0 9 2 13 13 7 3 16 0 9 1 0 0 9 1 11 2
10 11 11 2 11 2 0 9 11 2 11
3 9 13 9
11 1 9 13 3 0 9 2 3 7 0 9
12 1 9 9 9 3 13 9 11 1 0 9 2
13 1 9 1 10 9 7 13 0 9 2 3 0 2
25 7 15 9 1 10 0 0 9 13 7 1 0 9 9 1 0 9 7 3 3 0 9 1 9 2
13 13 15 15 3 9 13 1 0 12 7 12 9 2
2 11 11
32 0 9 2 16 4 9 3 0 9 2 3 13 9 9 2 1 15 4 3 9 3 15 13 2 13 2 13 3 3 1 15 2
12 13 4 15 3 3 3 2 16 16 13 9 2
21 15 7 13 2 16 13 13 10 9 7 15 15 13 9 2 16 15 13 3 0 2
2 9 9
6 9 13 1 12 9 2
9 1 15 14 0 12 13 0 9 2
38 0 9 2 15 15 3 13 1 9 9 2 13 0 2 9 1 9 13 13 9 1 0 9 7 1 0 9 13 13 1 9 7 0 0 9 0 9 2
13 0 9 9 13 2 7 1 12 9 15 3 13 2
30 7 3 2 16 0 9 9 1 9 9 1 0 9 13 0 1 0 9 2 0 14 3 0 9 15 1 0 9 13 2
7 0 9 13 1 0 9 2
16 0 9 15 9 13 13 15 0 9 7 13 15 1 15 15 2
19 1 9 2 9 7 0 0 9 1 9 2 0 1 9 2 13 3 9 2
3 9 15 13
29 9 9 1 10 9 7 9 1 15 15 13 3 3 1 15 2 3 15 13 1 9 7 9 2 16 1 0 9 2
14 15 15 13 10 9 2 0 9 15 13 1 0 9 2
40 3 15 15 13 2 13 13 1 9 9 2 1 15 2 16 15 14 3 13 7 3 3 13 2 0 13 1 15 0 9 2 2 3 13 0 15 13 7 15 2
32 9 9 2 15 13 13 1 9 2 1 9 9 15 9 11 13 3 3 2 3 4 13 13 0 9 1 9 1 0 9 9 2
11 0 9 1 9 13 7 1 9 9 3 2
7 9 13 3 0 9 9 2
12 1 0 9 0 12 9 15 15 14 12 13 2
20 1 15 9 13 13 0 9 3 1 0 9 1 0 9 2 9 2 9 2 2
10 3 15 7 9 0 9 13 0 9 2
8 13 1 9 7 1 9 9 2
6 1 0 13 15 0 2
20 1 15 13 13 7 15 15 15 4 1 3 13 2 3 13 0 9 9 9 2
24 16 9 13 12 7 12 5 0 9 2 15 15 13 1 0 9 2 13 15 13 9 3 0 2
2 9 9
13 9 1 9 11 13 0 0 9 12 7 12 9 2
10 13 0 9 2 1 15 9 13 9 2
8 15 13 0 1 12 0 9 2
24 9 15 3 13 1 9 1 9 1 9 7 0 9 2 9 13 13 1 9 9 0 9 9 2
7 9 15 3 1 9 13 2
5 9 13 9 9 2
26 13 1 9 0 9 7 0 9 0 0 9 2 3 1 9 3 7 1 9 0 9 1 10 10 9 2
7 9 13 1 0 0 9 2
14 13 9 1 9 10 9 2 9 9 7 0 9 9 2
3 9 1 9
15 0 1 9 13 1 0 7 9 2 1 15 13 9 9 2
8 15 13 3 16 9 1 9 2
31 9 15 3 13 13 9 2 15 13 3 13 0 9 9 1 0 9 2 16 4 15 13 0 9 9 7 9 15 3 13 2
21 3 4 13 2 16 4 1 10 9 13 3 14 12 9 2 7 14 12 16 3 2
12 3 4 15 3 13 2 13 4 15 10 9 2
24 13 1 15 13 0 9 9 9 7 9 1 1 0 9 9 2 7 1 9 1 0 9 9 2
38 1 0 9 9 13 7 1 9 0 9 2 16 13 9 1 12 9 2 16 4 13 9 9 7 1 0 9 3 13 9 2 15 3 13 1 9 9 2
36 9 2 11 2 9 2 9 2 0 2 2 1 9 12 2 12 12 11 2 9 2 2 2 12 2 12 12 2 9 2 2 12 2 12 12 2
5 2 9 1 9 2
5 7 9 13 13 2
10 13 2 16 1 15 13 9 7 9 2
5 1 9 13 9 9
10 9 0 7 0 9 7 13 9 0 9
13 11 2 9 0 7 0 9 2 13 1 0 11 2
17 9 0 9 1 0 9 13 9 13 10 9 0 3 0 0 9 2
6 1 0 9 13 2 9
11 13 9 0 0 9 7 11 15 3 13 2
18 9 13 3 0 2 7 10 9 15 13 2 13 15 9 9 11 11 2
9 1 9 1 0 9 13 9 0 2
21 13 0 9 1 9 1 9 7 0 7 0 9 15 13 0 9 14 1 10 9 2
7 11 13 14 12 0 9 2
13 0 9 1 15 9 13 14 9 0 9 9 9 2
6 9 9 3 13 9 2
21 0 1 15 13 0 9 7 9 15 1 9 13 1 9 7 9 1 0 9 9 2
13 14 9 9 15 13 3 1 9 2 9 0 9 2
16 9 9 13 13 7 1 0 0 9 1 11 7 1 0 9 2
19 11 11 2 1 0 9 13 3 13 12 9 0 9 2 3 13 0 9 2
19 3 1 9 1 9 13 14 1 0 9 2 0 9 2 0 9 7 9 2
2 0 9
14 13 0 9 9 13 12 1 10 0 9 2 13 9 2
13 13 3 2 16 15 13 10 10 9 1 9 3 2
23 9 7 9 2 7 7 9 0 9 2 13 10 9 3 14 12 9 7 9 1 10 9 2
9 3 1 12 12 9 13 1 0 2
9 9 7 13 15 9 3 2 3 2
19 13 2 14 11 13 1 9 2 13 15 1 0 9 7 0 9 1 15 2
5 15 9 3 13 2
4 13 2 15 13
17 1 12 9 9 13 0 9 9 2 15 15 3 13 7 1 9 2
13 9 15 13 3 2 3 1 0 9 3 7 9 2
16 9 13 1 9 1 9 2 3 13 9 1 0 9 9 9 2
7 9 7 13 9 9 3 2
8 13 15 3 0 9 1 9 2
15 16 9 3 13 2 13 14 2 15 13 13 2 13 9 2
17 11 13 1 9 1 12 1 12 5 3 1 0 9 7 10 9 2
20 1 11 11 15 3 13 1 0 9 7 3 0 9 2 3 1 9 0 9 2
19 1 9 9 4 1 12 9 13 12 9 2 3 3 15 13 12 9 9 2
18 0 9 15 13 3 12 12 9 7 1 9 13 1 9 10 9 9 2
10 13 9 2 9 9 7 9 2 2 2
8 0 9 1 9 9 13 9 2
23 3 1 0 9 9 1 15 13 12 5 1 9 9 7 9 15 13 13 1 15 7 3 2
15 9 13 13 12 1 9 0 9 2 15 13 1 0 9 2
2 11 0
39 9 2 11 2 9 0 7 0 9 2 9 2 9 2 0 2 2 12 12 0 11 2 9 2 2 2 12 2 12 2 12 2 9 2 2 12 2 12 2
1 11
34 9 11 2 9 2 9 2 0 2 2 1 9 1 9 11 2 15 13 14 10 9 9 1 0 2 7 3 9 1 9 9 0 9 2
18 3 1 9 1 11 2 9 9 2 15 9 13 0 9 0 0 9 2
30 9 9 3 1 0 9 1 9 2 1 15 15 13 3 9 9 2 3 13 3 1 9 0 9 13 9 1 0 9 2
17 9 2 11 2 9 2 9 2 0 2 2 0 12 2 12 12 11
17 9 11 2 15 13 1 9 1 0 9 9 1 0 9 0 11 2
16 9 13 1 14 12 9 0 9 0 0 9 2 0 9 9 2
10 9 9 1 0 9 13 0 7 0 2
30 9 2 11 2 0 2 9 2 2 0 12 2 12 12 11 2 9 2 2 2 12 2 12 2 9 2 2 12 2 12
22 9 11 2 9 9 2 1 9 7 9 9 9 2 9 7 0 9 2 1 9 2 2
20 3 0 9 0 9 2 0 0 0 9 7 9 0 9 2 13 0 0 9 2
18 15 13 0 0 9 1 0 9 2 15 15 9 13 3 1 0 11 2
32 9 2 11 2 9 9 2 11 11 12 2 12 12 0 11 2 9 2 2 2 12 2 12 12 2 9 2 2 12 2 12 12
5 2 14 2 0 9
18 12 10 9 2 9 2 13 2 16 13 15 13 2 7 13 15 13 2
30 1 10 0 9 15 13 7 1 10 9 9 2 15 2 15 13 1 9 2 3 1 9 2 9 14 1 2 9 2 2
34 1 0 9 15 3 13 9 2 16 4 3 3 13 0 9 2 16 3 13 2 16 7 9 15 13 13 0 2 3 13 0 2 9 2
28 1 15 2 16 13 9 7 9 2 4 15 13 1 9 1 0 9 2 1 15 15 13 0 9 10 0 9 2
26 1 9 13 7 7 9 1 0 9 7 0 9 2 15 13 9 2 9 7 9 0 1 9 1 9 2
19 1 9 15 9 13 1 9 9 2 9 2 9 7 9 1 0 0 9 2
22 1 10 9 2 3 13 13 13 9 2 7 13 1 0 9 1 9 2 13 7 9 2
12 13 4 1 15 1 9 9 2 12 2 12 2
9 1 9 1 10 9 1 9 13 2
7 3 13 3 1 15 0 2
15 3 15 4 13 13 2 16 10 9 4 4 9 3 13 2
6 1 15 4 13 13 2
13 1 0 9 13 9 1 12 1 12 9 9 9 2
10 1 9 0 9 13 0 9 3 0 2
24 3 7 1 9 1 9 15 9 13 14 1 12 9 9 9 2 16 9 9 13 1 0 9 2
42 0 9 13 2 16 1 0 9 0 9 1 12 2 1 0 9 2 2 7 12 2 1 9 1 9 2 13 3 2 16 13 0 9 9 7 0 9 1 9 3 9 2
27 9 15 3 13 15 9 2 15 4 1 9 13 16 9 7 9 7 13 1 15 2 16 13 0 7 0 2
14 13 3 7 9 9 2 16 3 9 2 9 2 9 2
17 7 9 2 9 13 13 14 1 0 9 2 7 3 1 0 9 2
2 16 2
16 0 9 7 0 9 15 2 15 13 9 15 2 15 15 13 2
2 11 0
4 1 9 1 9
13 0 9 2 15 1 15 13 1 9 7 15 1 9
18 9 2 0 9 2 15 13 1 10 9 7 1 9 1 9 7 9 2
9 3 1 9 1 10 9 3 13 2
4 13 15 0 2
26 3 13 0 13 1 9 9 2 16 0 9 15 0 13 2 16 1 9 13 1 0 9 1 0 9 2
20 3 15 10 9 0 13 2 16 0 9 13 0 9 7 4 13 0 9 9 2
13 15 3 13 2 16 13 0 13 14 9 3 0 2
14 13 13 7 9 2 15 13 0 9 2 7 9 0 2
18 0 13 7 0 1 9 2 15 0 9 1 9 9 13 2 0 13 2
35 16 0 10 9 13 7 1 9 9 0 9 13 2 13 15 9 2 16 0 4 13 9 2 15 0 1 9 10 9 1 9 0 9 13 2
3 1 15 13
31 1 9 0 1 9 2 16 0 9 4 13 1 0 9 1 10 9 9 2 13 9 0 9 2 0 1 9 0 7 0 2
26 0 9 13 9 2 1 15 0 13 1 15 2 16 9 2 15 13 0 2 13 0 1 0 9 9 2
33 10 9 0 13 7 1 9 2 1 0 9 2 2 7 1 9 1 0 7 0 2 3 0 9 0 2 3 1 9 0 9 2 2
12 1 0 9 3 13 0 9 1 0 7 0 2
43 16 15 1 0 9 2 10 9 13 3 9 9 0 2 13 1 0 9 9 2 13 0 13 1 0 9 0 1 9 7 0 13 0 10 9 0 1 9 1 0 9 13 2
26 9 10 9 13 7 13 9 9 2 3 0 0 9 0 2 2 7 9 2 13 2 14 1 0 9 2
13 0 9 13 1 9 1 9 1 9 0 7 0 2
72 13 2 14 1 9 0 2 13 0 13 2 12 2 0 9 9 2 12 2 9 0 9 7 0 9 2 12 2 9 9 7 13 13 1 9 2 16 15 0 9 13 1 9 3 2 3 7 13 13 1 0 9 10 9 2 2 7 16 0 9 13 0 9 9 2 3 3 12 0 9 2 2
15 13 2 14 1 9 0 2 13 0 13 1 0 0 9 2
20 12 2 9 1 9 9 7 9 1 9 13 2 16 0 9 13 0 9 9 2
17 12 2 9 1 0 9 1 9 2 16 13 9 13 7 1 9 2
3 9 1 9
14 9 9 0 9 13 13 3 0 1 9 9 9 0 2
48 16 13 1 9 0 9 0 10 9 9 2 3 0 9 13 13 14 1 9 10 9 1 9 2 16 0 13 9 1 9 3 1 12 9 1 9 9 7 3 7 3 13 1 9 9 0 9 2
17 9 0 9 13 0 13 3 1 0 2 1 15 4 0 9 13 2
30 13 2 14 7 0 2 3 1 0 9 2 13 1 9 0 9 2 13 0 9 1 9 1 9 0 1 9 0 9 2
10 0 13 0 13 10 9 1 0 9 2
11 0 9 13 1 0 9 9 0 0 9 2
12 2 13 2 14 1 9 0 9 2 12 9 2
11 2 13 2 14 1 9 9 2 12 9 2
11 2 13 2 14 1 9 9 2 12 9 2
13 2 13 2 14 1 9 0 9 2 3 12 9 2
13 0 0 9 13 0 0 9 13 2 3 7 13 2
2 11 11
4 9 1 9 2
3 0 9 2
10 13 1 15 12 9 0 7 0 9 2
3 1 0 9
15 13 9 2 15 13 9 0 9 1 9 1 11 7 11 2
31 1 15 2 15 15 15 13 1 9 3 0 9 7 3 3 13 9 7 9 7 9 2 15 13 1 0 9 1 0 9 2
7 9 13 13 14 0 9 2
13 7 15 1 9 2 16 13 9 1 10 9 13 2
17 3 1 15 2 15 13 13 9 1 9 12 2 12 0 9 9 2
19 11 13 0 1 0 2 7 3 0 9 2 15 15 13 13 10 0 9 2
26 10 9 15 1 10 9 13 7 1 0 9 7 9 2 1 15 15 13 9 9 9 2 15 11 13 2
11 9 13 1 0 9 7 3 3 0 9 2
11 0 9 0 9 13 9 9 9 9 9 2
14 13 15 15 13 1 9 9 1 0 9 9 9 12 2
9 3 15 3 13 9 2 0 9 2
2 0 9
30 3 0 9 1 9 9 0 9 0 7 0 9 2 3 15 13 9 2 15 15 13 12 2 9 1 0 9 1 11 2
20 4 13 0 9 3 0 9 1 0 7 0 9 7 0 9 1 9 0 9 2
31 9 2 9 0 9 2 9 3 0 9 2 1 9 12 9 2 12 12 11 12 2 11 2 9 2 2 2 12 2 12 12
5 9 2 9 7 15
2 9 9
12 13 4 9 1 9 2 15 4 15 15 13 2
19 3 4 4 9 13 2 16 4 9 13 1 9 2 15 13 1 9 0 2
5 13 9 9 0 2
6 11 2 11 2 2 11
25 9 13 3 2 7 1 12 2 9 12 0 0 9 2 11 2 13 13 9 2 15 13 9 13 2
30 3 13 13 1 9 0 2 10 9 13 13 2 15 15 13 2 10 9 15 13 2 15 13 2 13 13 13 7 13 2
28 9 13 4 13 1 0 9 9 7 9 3 2 16 4 12 9 13 1 9 7 16 4 0 9 13 12 9 2
51 1 10 0 9 13 9 13 2 1 12 9 2 12 11 2 9 2 9 7 9 9 2 0 9 2 7 9 7 9 0 9 2 2 9 0 9 2 9 9 7 1 9 13 13 0 2 15 15 9 13 2
26 1 9 0 13 9 3 13 0 9 0 9 7 9 1 15 2 16 15 1 9 13 13 1 0 9 2
18 13 7 10 9 2 16 4 9 9 13 7 1 0 9 9 9 13 2
27 13 2 16 9 15 13 1 9 9 9 1 12 9 2 12 11 2 16 4 1 0 9 9 13 7 13 2
2 0 9
15 1 9 10 9 1 9 4 13 13 2 16 9 3 13 2
8 7 4 1 10 9 13 9 2
9 1 15 4 13 1 9 0 9 2
8 13 0 15 1 10 9 13 2
7 11 2 11 2 2 0 11
34 1 9 9 1 9 9 2 15 15 4 3 13 2 15 13 13 1 12 9 1 9 9 1 0 9 1 9 2 15 13 1 9 13 2
6 9 13 0 3 13 2
3 9 15 9
10 1 9 9 1 9 4 15 13 9 2
16 1 9 3 4 15 0 9 13 7 13 4 15 1 9 13 2
5 13 3 10 9 2
6 11 2 11 2 2 11
27 9 15 13 13 3 1 9 1 9 2 15 13 3 10 9 2 7 0 9 0 9 2 15 1 9 13 2
11 3 13 2 16 9 9 15 9 13 0 2
30 13 4 3 13 2 16 9 15 9 4 13 1 9 0 0 9 9 14 3 2 13 2 14 15 9 15 0 0 9 2
26 4 2 14 9 13 3 2 7 3 2 13 9 0 9 14 3 2 13 2 14 9 0 1 0 9 2
2 0 9
12 1 9 4 15 14 0 9 13 1 0 9 2
12 9 15 13 0 9 2 15 4 13 13 3 2
23 16 13 2 16 9 13 3 2 13 4 15 2 16 13 10 0 9 3 15 13 10 9 2
6 11 2 11 2 2 9
8 3 13 1 9 9 0 9 2
12 13 15 9 1 9 15 2 0 1 0 9 2
11 0 9 13 13 1 9 12 7 12 11 2
37 9 9 13 0 9 13 7 1 0 9 9 7 1 9 9 2 13 2 14 1 9 13 9 1 9 0 9 7 13 2 14 15 1 9 0 9 2
40 1 0 9 13 9 13 2 16 4 1 12 9 1 9 0 9 13 0 9 3 9 9 2 7 16 4 1 10 9 13 1 9 2 15 0 9 13 2 9 2
15 0 9 13 4 13 9 1 0 9 2 0 9 13 13 2
23 16 13 0 9 13 1 0 9 7 14 12 1 9 2 9 9 15 9 13 1 0 9 2
11 1 10 9 13 4 9 13 1 9 0 2
25 13 2 14 13 9 1 0 9 3 2 13 15 15 0 9 1 0 9 7 9 9 3 13 9 2
38 0 9 13 13 2 13 2 14 1 9 2 1 15 13 13 7 13 9 2 7 13 2 14 0 9 9 2 7 16 4 13 4 0 9 13 1 9 2
14 13 2 14 1 0 9 13 9 2 13 9 0 9 2
17 3 0 9 2 1 9 12 9 0 1 9 9 2 9 9 13 2
3 9 1 9
16 13 1 0 9 7 13 4 13 9 1 9 9 0 9 9 2
13 13 0 9 7 13 4 13 9 1 9 12 9 2
7 7 15 13 1 15 15 2
8 13 15 4 9 0 9 13 2
6 11 2 11 2 2 11
42 9 12 11 13 2 16 4 1 9 9 9 9 13 9 3 7 3 1 0 9 2 13 2 14 15 9 9 7 13 2 14 1 0 7 3 0 9 2 7 9 9 2
25 1 9 9 9 9 1 0 9 13 0 3 0 7 0 9 9 7 3 9 0 9 7 9 9 2
17 7 13 0 9 13 2 1 10 9 2 9 1 9 9 1 9 2
14 9 13 2 11 11 2 9 9 0 9 1 11 12 2
5 13 9 9 2 12
15 1 0 9 0 9 10 9 13 9 9 2 0 11 11 2
6 0 9 2 9 11 2
13 16 13 12 9 2 13 1 15 0 7 11 11 2
10 13 9 9 2 16 1 11 13 9 2
9 15 13 9 9 9 1 9 9 2
16 2 9 1 11 2 11 2 11 2 1 9 2 15 13 13 2
11 12 1 3 0 9 13 13 9 11 9 2
13 3 3 9 9 1 9 1 11 9 13 1 15 2
15 2 1 0 9 11 11 13 7 3 13 2 15 13 3 2
1 9
8 2 0 9 7 9 9 9 2
34 9 2 11 2 9 2 0 12 2 12 12 11 12 2 9 11 2 9 2 2 2 12 2 12 12 2 9 2 2 12 2 12 12 2
9 2 0 9 2 0 9 1 9 2
15 9 2 9 2 9 12 2 9 7 9 12 2 12 9 2
32 9 2 11 2 9 2 0 2 7 0 9 2 9 9 2 11 9 12 2 12 12 11 12 2 9 2 2 2 12 2 12 2
23 2 9 1 0 9 2 1 2 0 2 0 2 9 7 9 1 9 13 0 2 9 2 2
32 9 2 11 2 9 2 0 2 7 0 9 2 9 9 2 11 9 12 2 12 12 11 12 2 9 2 2 2 12 2 12 2
23 2 0 9 1 0 9 2 0 0 9 1 9 2 9 2 3 9 1 9 0 9 2 2
32 9 2 11 2 9 2 0 2 7 0 9 2 9 9 2 11 9 12 2 12 12 11 12 2 9 2 2 2 12 2 12 2
13 2 0 9 2 9 9 2 0 9 0 1 11 2
25 9 2 13 9 1 9 1 0 9 3 2 16 4 13 0 9 7 13 3 13 1 9 9 9 2
9 9 2 12 2 9 2 9 12 2
26 9 2 9 9 11 11 2 0 12 2 12 12 11 11 2 9 2 5 9 2 2 12 2 12 12 2
21 2 0 9 1 11 2 9 1 9 7 0 9 0 1 9 9 1 11 1 9 2
9 9 2 12 2 9 2 9 12 2
26 9 2 9 9 11 11 2 0 12 2 12 12 11 11 2 9 2 5 9 2 2 12 2 12 12 2
33 2 9 1 9 0 9 2 9 9 1 9 1 9 7 9 1 0 9 9 2 9 2 9 7 9 2 1 0 9 9 7 9 2
5 9 2 9 12 2
26 9 2 9 9 11 11 2 0 12 2 12 12 11 11 2 9 2 5 9 2 2 12 2 12 12 2
10 2 0 9 2 1 0 9 0 9 2
9 9 2 12 2 9 2 9 12 2
26 9 2 9 9 11 11 2 0 12 2 12 12 11 11 2 9 2 5 9 2 2 12 2 12 12 2
17 2 0 7 0 9 2 9 7 0 9 0 1 9 9 1 9 2
32 9 2 11 2 9 2 9 2 0 2 2 0 12 2 12 12 11 12 2 9 2 5 9 2 2 12 2 12 12 2 12 2
4 2 9 9 2
13 9 2 12 2 12 2 2 12 2 12 2 12 2
2 9 2
22 11 2 9 2 9 2 0 2 2 0 12 2 12 12 11 12 2 9 2 5 9 2
8 2 12 2 12 12 2 12 2
39 2 0 9 2 9 9 2 3 13 1 9 7 1 9 2 3 13 9 10 7 9 9 2 9 1 0 7 0 9 9 2 0 9 7 9 9 1 9 2
32 9 2 11 2 9 2 9 2 0 2 2 0 12 2 12 12 11 12 2 9 2 5 9 2 2 12 2 12 12 2 12 2
13 2 0 9 2 0 9 1 9 1 9 0 9 2
12 9 9 2 9 2 0 9 7 9 1 9 2
11 9 2 12 2 2 12 2 12 2 12 2
32 9 2 11 2 9 2 9 2 0 2 2 0 12 2 12 12 11 12 2 9 2 5 9 2 2 12 2 12 12 2 12 2
27 2 0 11 2 9 9 1 9 2 9 0 9 2 9 0 9 2 9 1 9 2 0 9 9 0 9 2
2 12 2
32 9 2 11 2 9 2 9 2 0 2 2 0 12 2 12 12 11 12 2 9 2 5 9 2 2 12 2 12 12 2 12 2
8 2 0 9 2 9 9 9 2
14 12 0 9 2 0 9 9 7 0 9 7 0 9 2
32 9 2 11 2 9 2 9 2 0 2 2 0 12 2 12 12 11 12 2 9 2 5 9 2 2 12 2 12 12 2 12 2
3 9 1 9
8 12 9 3 13 1 10 9 2
3 0 9 13
15 9 10 9 3 1 11 9 13 9 1 0 9 0 9 2
10 9 9 10 9 3 13 12 2 9 2
47 1 1 15 2 16 13 1 15 2 13 2 10 9 9 2 1 9 2 13 10 0 9 1 0 9 2 7 0 9 1 9 0 9 4 3 3 13 2 13 7 10 9 1 10 9 13 2
12 1 10 9 13 9 1 9 3 12 12 9 2
15 9 7 13 7 0 3 0 9 2 1 15 13 1 3 2
13 0 9 13 0 9 7 1 0 9 13 3 9 2
24 15 1 10 9 7 9 15 13 13 10 0 9 13 2 14 13 10 9 2 3 13 0 9 2
4 9 2 9 12
12 9 1 11 11 2 9 0 7 0 9 11 9
17 0 9 7 0 9 1 10 9 1 15 13 9 7 0 9 9 2
6 15 15 15 13 13 2
33 0 9 13 9 7 3 14 10 9 1 0 9 7 9 2 7 16 4 1 9 12 13 9 1 9 7 13 13 1 9 11 11 2
11 1 15 4 15 13 9 10 9 7 9 2
40 13 4 15 1 9 0 9 2 3 1 9 9 1 0 11 7 9 1 10 9 7 9 13 14 3 3 2 16 15 1 15 13 3 13 10 9 2 16 0 2
26 15 13 1 9 7 3 2 3 13 1 9 11 2 11 2 11 7 9 11 9 0 9 10 0 9 2
7 13 2 16 15 13 9 2
45 16 15 1 15 3 13 2 3 15 13 2 16 9 7 9 13 7 1 0 9 2 16 13 0 9 7 16 4 15 13 3 13 2 13 4 13 11 1 0 9 15 13 1 9 2
10 3 0 13 7 9 13 2 16 3 2
5 14 15 13 3 2
16 1 9 1 9 2 0 9 7 0 9 15 1 15 13 13 2
7 13 3 1 15 13 9 2
13 13 3 1 0 9 7 13 15 4 15 3 13 2
14 3 4 15 13 1 0 9 1 9 2 3 1 9 2
9 13 15 1 0 9 2 1 9 2
24 1 9 15 13 2 7 0 9 7 0 9 13 13 2 7 16 15 13 3 1 9 1 9 2
20 1 15 2 16 4 9 13 13 15 2 15 13 7 3 13 2 13 13 9 2
15 15 13 10 9 7 1 9 0 9 10 9 9 11 11 2
3 9 9 2
27 3 13 0 11 7 15 14 3 14 3 2 16 10 9 13 1 11 7 10 9 1 0 9 11 2 11 2
20 13 4 15 13 9 9 7 9 11 2 11 2 11 2 11 2 11 2 11 2
7 15 13 0 7 0 9 2
10 15 15 13 13 9 1 0 10 9 2
10 1 15 7 13 13 12 2 9 2 2
17 3 4 13 9 9 1 11 2 13 9 7 13 15 3 13 9 2
25 12 4 1 9 13 1 9 12 9 0 9 2 10 7 14 9 13 1 11 13 7 13 15 13 2
9 15 4 15 13 1 15 1 9 2
15 14 12 9 4 15 7 13 1 9 2 0 4 13 9 2
8 14 15 9 7 0 9 13 2
3 9 9 13
21 3 0 13 13 9 0 9 3 0 11 11 2 16 10 9 11 14 13 10 9 2
16 0 0 9 9 7 9 3 3 1 0 9 13 9 1 9 2
10 13 3 9 2 1 15 7 15 13 2
13 9 13 2 9 13 1 15 2 9 0 9 3 2
15 1 0 9 1 0 9 1 11 13 14 13 7 13 15 2
9 3 15 2 3 3 2 3 13 2
23 11 11 4 13 1 9 2 3 15 13 9 11 7 9 11 2 12 9 2 12 9 2 2
10 11 11 15 3 2 1 9 2 13 2
4 13 4 1 9
21 15 3 13 9 11 11 2 11 3 2 16 13 0 9 1 9 9 1 9 9 2
15 1 9 7 12 15 3 3 13 10 9 1 9 9 11 2
29 15 15 13 1 10 9 1 0 0 9 2 15 15 13 14 1 11 1 10 10 3 0 9 2 13 1 9 9 2
20 1 9 9 11 3 13 13 15 7 13 1 10 9 7 16 4 15 13 15 2
24 7 15 3 13 2 16 9 2 15 4 10 9 13 2 15 13 1 9 2 7 16 13 0 2
10 1 15 13 3 9 3 16 0 9 2
2 0 9
29 3 14 3 0 9 2 3 3 0 2 4 13 13 2 16 0 0 9 1 9 9 11 11 7 11 11 13 9 2
23 3 3 13 7 9 15 13 2 16 3 1 11 11 13 1 9 2 1 9 2 10 9 2
17 13 9 13 2 3 0 2 0 0 7 13 0 0 7 0 9 2
18 0 15 3 3 13 9 11 7 11 2 15 13 9 9 1 0 9 2
16 9 1 9 13 11 11 3 1 0 9 3 15 13 0 9 2
5 9 7 1 15 2
3 9 3 13
15 13 3 1 0 9 2 15 0 1 15 13 9 11 11 2
29 10 9 1 0 9 11 11 3 9 1 0 9 3 3 13 2 7 9 9 1 15 2 15 15 13 2 3 13 2
18 13 15 7 13 1 9 11 2 3 13 0 9 2 16 13 10 9 2
6 1 10 9 15 13 2
11 13 4 16 9 1 9 2 13 15 0 2
11 3 15 13 1 0 9 1 9 0 9 2
7 3 14 0 9 1 12 2
2 0 9
8 13 9 9 1 9 11 11 2
14 1 0 9 1 10 9 13 9 2 9 7 9 9 2
9 13 3 2 3 15 14 3 13 2
7 1 0 9 2 1 9 2
21 13 4 15 13 2 16 15 13 0 9 1 9 7 9 2 7 1 9 1 9 2
8 1 15 15 13 9 7 9 2
9 0 9 15 11 11 3 13 9 2
9 7 9 9 7 0 9 15 13 2
4 12 9 13 9
10 1 12 9 9 15 13 1 0 9 2
7 0 9 2 0 9 7 9
12 1 0 12 9 13 9 0 9 1 12 9 2
10 13 15 1 0 9 1 0 9 9 2
32 9 4 15 13 13 3 3 2 3 9 13 0 9 0 9 7 9 9 2 15 15 3 13 1 0 12 5 9 1 0 9 2
2 11 9
19 0 9 13 1 9 11 0 3 3 2 16 15 4 13 1 9 0 9 2
33 13 2 16 9 13 0 0 2 7 0 9 9 0 9 1 9 1 9 11 11 2 7 0 9 2 15 13 1 11 0 12 9 2
26 0 0 9 13 9 1 0 9 1 11 2 15 1 9 0 9 1 0 9 13 3 14 12 5 11 2
2 0 9
9 0 9 13 9 0 9 7 9 2
34 9 11 2 15 13 0 10 9 1 11 2 13 1 0 9 3 9 2 16 3 1 9 12 13 9 12 9 2 0 9 2 9 2 2
27 13 1 15 9 0 9 2 0 0 9 0 9 7 9 9 2 15 13 0 0 9 0 9 1 0 9 2
24 0 9 15 9 13 13 1 12 9 1 12 9 2 9 2 3 1 9 9 9 7 9 9 2
18 11 3 13 1 9 9 9 3 1 9 9 2 3 0 7 0 9 2
18 13 15 2 16 9 9 1 12 9 13 9 9 1 12 9 2 9 2
21 16 4 9 13 9 9 1 12 9 2 9 4 15 13 3 1 12 9 9 9 2
32 3 15 13 7 0 0 9 0 9 7 0 9 11 2 15 13 1 0 9 9 1 9 12 9 9 1 12 9 9 1 9 2
23 9 13 0 0 9 2 15 9 13 13 9 1 10 9 2 3 1 9 0 7 0 9 2
18 11 3 3 13 1 12 9 2 9 9 1 0 0 9 1 0 11 2
21 1 9 0 9 13 3 0 13 0 9 1 0 9 2 16 3 1 3 0 11 2
25 9 1 9 9 0 9 1 11 13 13 1 12 1 12 9 2 16 1 11 4 13 14 12 9 2
24 7 15 9 0 9 1 11 13 13 7 3 15 13 9 0 9 2 1 10 9 15 13 9 2
3 9 13 9
20 11 7 11 2 15 13 1 11 1 0 9 2 13 1 0 12 9 0 9 2
17 3 9 0 9 11 15 1 9 12 2 12 13 1 12 1 12 2
6 9 13 12 9 9 2
12 1 9 9 7 9 9 13 9 12 9 9 2
20 9 4 3 13 1 12 9 2 3 13 12 9 2 3 14 9 1 0 9 2
14 13 15 15 3 13 9 9 9 12 1 3 16 12 2
9 1 0 9 13 1 11 0 9 2
25 1 0 12 9 9 12 13 11 9 12 9 9 2 16 1 0 9 3 13 0 9 12 9 9 2
8 13 3 3 1 0 9 9 2
20 12 9 1 0 9 13 3 9 0 9 2 15 13 1 9 14 12 5 9 2
3 9 9 2
11 0 9 3 13 0 0 9 2 0 9 2
21 16 1 9 12 13 1 11 10 9 3 0 2 1 0 12 9 13 1 0 9 2
21 0 9 9 9 7 0 9 13 9 0 9 2 16 13 1 9 1 9 12 9 2
17 12 5 9 1 3 0 9 13 1 9 1 0 9 1 0 9 2
18 0 9 2 15 13 0 1 9 9 2 3 13 3 0 9 0 9 2
35 1 0 12 9 9 0 9 13 1 9 2 3 1 9 1 0 9 2 12 9 9 7 1 0 12 9 9 13 9 13 1 0 12 9 2
24 9 13 13 9 9 0 9 2 15 3 13 14 12 5 9 7 3 13 13 1 12 5 9 2
18 0 9 0 9 13 0 9 2 15 3 13 1 9 12 1 12 5 2
9 10 9 15 13 14 1 0 9 2
4 9 13 1 5
7 2 2 9 1 12 2 9
7 9 1 9 2 0 9 2
8 13 1 9 1 0 0 9 2
11 1 9 9 1 9 15 13 3 13 9 2
5 9 2 0 9 2
2 9 2
3 0 9 2
1 9
5 9 2 9 2 9
39 13 0 2 0 2 0 2 0 11 2 9 2 9 2 0 2 2 12 12 11 12 2 11 2 11 1 11 12 2 9 2 2 9 2 2 12 2 12 2
22 9 2 11 1 11 2 0 11 12 2 1 9 2 11 2 9 2 11 2 0 9 2
24 9 0 9 1 0 9 11 12 2 9 2 9 2 9 2 9 7 15 2 15 1 15 13 2
29 9 12 2 9 2 9 2 9 2 9 2 9 2 9 2 9 0 7 0 2 12 2 2 12 2 12 2 12 2
46 13 9 11 2 9 2 9 2 0 2 2 12 12 11 2 0 9 2 11 12 2 9 2 2 2 12 2 12 12 2 12 2 9 12 2 9 2 2 9 2 2 12 2 12 12 2
71 9 2 11 2 0 9 2 11 1 11 2 11 2 9 11 2 11 2 11 2 0 9 2 0 11 2 9 2 11 2 9 11 9 2 11 2 9 0 9 2 9 2 0 9 2 11 2 9 2 11 2 11 2 9 2 11 1 11 2 11 1 11 2 9 11 2 11 2 0 9 2
3 0 9 2
23 11 2 9 11 2 1 12 9 2 2 11 2 11 2 9 1 11 2 1 12 9 2 2
49 9 12 2 12 2 0 11 2 11 2 9 2 11 2 9 0 9 2 11 2 0 9 0 9 2 11 2 9 0 9 2 11 1 11 2 11 2 9 1 9 2 9 1 11 2 9 9 9 2
17 0 9 2 9 2 9 2 9 1 0 12 2 1 12 9 2 2
5 9 12 2 12 2
27 13 0 9 2 12 12 11 12 2 11 2 9 12 2 9 12 2 9 2 2 9 2 2 12 2 12 2
16 9 2 0 9 2 11 2 9 2 11 1 11 2 9 11 2
17 0 9 2 11 12 2 0 9 2 0 9 2 1 0 9 9 2
5 9 12 2 12 2
34 13 11 2 9 1 9 7 9 2 12 12 11 12 2 0 9 12 2 9 2 2 2 12 2 12 12 2 12 2 9 2 12 12 2
21 9 2 11 2 2 0 9 2 11 1 11 2 11 2 9 11 2 11 2 11 2
5 9 12 2 12 2
40 13 11 2 9 2 9 2 0 2 2 0 9 2 12 12 11 12 2 0 12 2 9 2 2 2 12 2 12 2 12 2 9 2 2 12 2 12 2 12 2
14 11 12 2 9 2 0 9 2 9 12 2 0 9 2
22 12 2 9 0 0 7 0 9 9 7 0 9 2 12 2 2 12 2 12 2 12 2
39 13 11 2 9 1 9 9 7 9 2 12 12 11 12 2 9 2 0 9 12 2 9 2 2 2 12 2 12 2 12 12 2 9 2 2 12 2 12 2
11 9 2 11 2 0 9 2 11 2 9 2
16 0 9 2 11 12 2 0 9 2 0 9 1 0 9 9 2
7 9 1 9 9 7 9 2
10 9 15 1 9 9 7 0 9 13 2
14 9 13 7 0 9 2 9 11 15 3 13 9 9 2
3 1 0 9
10 0 9 1 9 2 7 1 9 15 13
27 0 9 0 9 2 3 0 9 11 2 3 13 1 0 0 9 3 12 9 9 7 13 15 12 9 9 2
11 9 9 13 0 9 7 9 9 0 9 2
2 11 9
14 9 7 13 9 10 0 9 2 7 9 13 3 13 2
17 3 13 0 2 9 2 13 1 9 7 9 3 12 9 9 3 2
14 3 12 9 9 13 9 7 12 9 9 9 0 9 2
16 0 12 9 9 15 3 13 13 1 0 9 2 3 0 9 2
7 9 9 4 3 13 9 2
27 0 9 13 12 9 1 12 9 2 15 13 3 2 16 1 15 15 1 11 13 2 13 0 9 11 11 2
3 9 1 9
6 0 9 13 13 9 2
24 3 3 13 9 2 11 2 12 9 9 9 1 0 9 2 3 4 13 13 1 9 7 9 2
18 13 15 7 13 3 0 9 1 10 9 7 13 1 15 9 0 9 2
22 1 10 9 3 13 9 9 1 9 9 2 13 9 9 0 2 9 2 11 11 9 2
9 9 1 0 9 13 3 12 9 2
15 3 3 15 4 13 9 9 2 7 16 1 9 9 13 2
13 1 0 9 9 9 3 13 2 16 9 9 13 2
17 3 0 9 13 0 9 2 1 15 13 13 9 9 1 0 9 2
19 16 15 9 1 9 13 2 13 0 9 2 3 0 1 12 7 12 9 2
17 16 13 1 0 0 9 7 13 9 1 9 2 13 13 9 9 2
3 1 0 9
20 13 15 2 16 13 1 3 0 9 2 15 7 13 0 9 1 9 0 9 2
9 9 0 7 0 9 15 3 13 2
14 16 4 13 0 9 3 13 2 13 0 9 0 9 2
10 9 4 13 13 1 9 1 0 9 2
11 13 4 15 7 13 0 9 7 0 9 2
19 13 15 2 16 15 3 13 9 2 7 13 0 0 9 2 13 11 11 2
22 3 15 9 13 0 9 1 9 9 1 12 9 7 0 9 1 10 9 7 9 9 2
2 1 9
12 9 1 9 9 15 13 1 12 7 12 9 2
12 0 9 15 13 13 2 7 15 1 9 13 2
13 3 9 10 9 2 0 9 2 13 9 0 9 2
9 7 13 9 13 1 9 0 9 2
10 1 9 13 4 13 0 9 0 9 2
11 0 9 13 0 13 7 9 0 9 9 2
25 13 15 13 9 3 3 1 9 3 0 7 0 9 2 12 7 12 9 2 2 9 1 0 9 2
11 9 13 1 9 0 9 7 0 0 9 2
11 9 0 9 13 3 0 9 9 0 9 2
20 9 13 1 0 9 2 12 2 12 9 1 12 9 2 2 16 13 0 9 2
8 7 9 15 13 9 9 9 2
14 0 13 2 16 3 7 3 4 7 9 1 9 13 2
35 9 2 0 9 2 0 2 9 2 2 11 12 2 12 12 11 11 2 9 2 2 2 12 2 12 12 2 9 2 2 12 2 12 12 2
11 9 2 1 9 13 9 0 9 1 9 2
1 11
15 11 9 13 0 9 9 11 2 15 13 1 0 9 9 2
10 13 1 9 9 2 9 7 9 9 2
5 11 11 2 11 11
14 9 13 1 9 1 9 2 15 4 13 1 0 9 2
23 0 9 11 13 9 1 0 11 1 12 0 9 2 3 1 15 13 0 1 0 0 9 2
23 9 13 9 1 11 11 1 0 9 1 9 12 2 15 4 15 1 9 13 13 1 9 2
17 1 0 9 13 11 2 1 0 9 14 12 9 9 2 12 9 2
16 1 9 0 11 13 7 0 9 9 11 2 0 1 9 12 2
48 3 9 0 9 11 11 2 15 15 1 9 10 9 2 13 1 9 12 2 13 1 9 10 0 9 2 13 9 2 7 13 10 0 9 2 1 15 7 0 9 11 2 2 13 9 0 9 2
33 9 1 9 13 15 2 15 1 0 9 13 2 0 9 2 0 9 7 3 10 9 13 0 9 2 11 11 2 7 0 0 9 2
16 3 0 9 9 2 0 2 9 2 9 2 13 3 0 9 2
40 9 0 9 2 1 15 9 11 13 9 11 2 15 3 13 7 10 9 9 13 2 2 13 9 9 0 2 1 15 13 1 9 9 9 7 9 11 13 9 2
4 7 14 15 2
14 0 9 10 9 13 3 9 1 9 2 9 1 9 2
16 11 9 15 3 3 13 9 9 2 15 13 0 7 0 9 2
64 7 3 2 16 9 13 0 9 2 11 9 13 3 3 3 13 3 1 0 11 2 2 15 4 15 13 2 0 2 1 0 9 2 13 15 13 7 15 2 15 15 13 1 10 0 9 0 9 13 3 2 9 13 3 10 9 2 16 7 0 3 13 9 2
14 1 9 4 3 13 9 0 9 9 1 0 9 9 2
51 16 15 3 13 13 0 9 1 9 2 7 13 0 9 1 9 2 1 9 0 9 1 11 13 9 11 3 9 2 2 13 11 9 13 16 0 9 1 10 9 2 15 1 15 1 0 9 13 9 9 2
16 16 7 13 1 9 2 0 2 9 13 1 9 1 0 9 2
10 12 9 9 4 1 15 13 3 3 2
5 9 1 9 2 2
13 9 11 2 9 2 9 7 9 2 15 13 13 2
3 9 0 9
3 9 3 0
3 13 9 9
4 1 9 0 9
18 1 10 9 15 14 1 9 12 2 9 0 9 13 0 9 0 9 2
18 1 0 9 9 2 15 13 4 13 9 1 9 2 13 12 0 9 2
12 1 9 4 0 9 13 14 1 12 9 9 2
33 0 9 4 1 0 9 0 1 12 2 9 12 13 13 9 9 11 2 0 2 9 2 2 10 9 13 0 13 7 1 0 9 2
19 13 9 2 3 4 13 1 9 0 0 9 12 9 1 9 1 0 9 2
16 0 0 9 13 0 0 0 9 7 11 2 0 2 9 2 2
11 9 4 13 1 15 9 9 1 0 9 2
21 10 9 13 1 0 9 9 2 15 1 9 1 0 9 4 1 0 9 3 13 2
6 0 9 9 2 9 2
22 10 9 7 4 13 9 9 2 1 15 15 4 3 13 7 9 0 9 7 9 9 2
12 0 9 0 9 1 9 11 13 3 12 9 2
15 0 9 9 0 9 1 0 9 9 4 13 0 9 11 2
14 1 0 0 9 0 11 4 3 13 9 9 10 9 2
22 9 9 13 9 9 0 9 0 0 9 2 15 15 13 1 0 0 2 9 2 11 2
24 10 9 13 0 9 9 1 0 9 11 2 0 2 9 2 7 3 1 0 9 1 0 9 2
8 13 7 9 2 15 15 13 2
33 1 0 9 4 0 9 1 9 13 3 1 9 9 2 9 2 3 2 9 0 9 2 7 9 9 7 9 9 9 1 0 9 2
3 9 0 9
18 1 9 12 13 1 0 9 1 10 9 3 14 9 11 7 9 11 2
14 10 9 13 3 7 1 9 0 9 0 9 0 9 2
15 7 1 9 9 9 12 9 15 3 13 9 0 0 9 2
21 0 9 9 10 9 13 1 9 9 3 1 9 0 1 0 9 15 9 1 9 2
40 15 2 15 13 1 9 10 9 7 13 10 9 1 9 2 13 1 9 0 9 9 12 2 12 2 12 2 3 16 9 0 9 2 15 10 9 13 9 9 2
15 0 9 9 0 0 9 13 3 9 9 0 16 1 9 2
15 1 0 9 1 9 15 7 9 11 7 9 11 3 13 2
14 13 15 3 3 0 0 9 1 9 0 9 9 9 2
23 0 9 11 1 0 9 15 3 3 13 1 9 1 0 9 1 9 9 2 3 12 5 2
2 0 9
9 9 13 1 0 9 0 9 9 2
47 0 9 9 10 9 2 0 1 9 7 1 0 9 2 13 1 9 1 0 9 3 0 2 12 9 3 9 11 2 7 15 1 15 15 9 0 9 13 1 0 3 16 11 1 9 9 2
18 3 7 3 15 9 1 9 3 13 1 9 0 1 15 2 0 0 2
12 9 9 10 9 15 3 13 1 9 10 9 2
35 9 7 9 0 9 10 9 2 0 9 2 3 7 1 0 9 13 10 9 1 9 9 9 2 15 13 9 9 7 13 15 3 3 9 2
25 13 0 2 16 1 9 9 9 15 15 0 9 7 9 4 13 13 9 15 0 9 1 10 9 2
9 15 13 1 9 9 9 0 9 2
24 10 9 13 3 0 1 9 2 15 13 1 0 9 7 13 1 0 2 7 0 9 9 9 2
25 0 9 4 13 13 1 9 0 2 0 2 9 9 9 1 0 9 7 15 13 2 3 4 13 2
2 11 11
3 11 2 11
37 9 2 0 0 9 2 0 2 9 2 2 11 12 2 12 12 11 12 2 9 2 2 2 12 2 12 12 2 9 2 2 12 2 12 12 12 2
3 13 0 9
1 11
9 2 11 2 9 2 9 2 0 2
27 9 2 0 12 2 12 12 11 12 2 9 2 2 2 12 2 12 12 2 9 2 2 12 2 12 12 2
6 2 9 2 9 12 2
6 2 9 9 2 12 2
26 2 9 2 0 2 0 9 1 9 9 2 9 1 9 0 9 2 0 9 0 2 3 0 2 9 2
22 2 9 2 9 0 1 9 0 9 2 0 9 2 0 9 1 9 2 9 0 9 2
4 2 9 9 2
6 1 0 9 12 13 2
22 2 9 2 2 1 9 2 2 3 1 9 2 9 9 15 13 1 12 1 12 9 2
5 12 3 0 9 2
25 2 1 0 9 13 2 16 4 15 9 9 13 1 12 2 13 9 9 11 11 2 1 9 2 2
16 3 1 10 9 13 0 9 9 2 0 9 1 15 7 9 2
30 13 3 14 1 1 15 0 0 9 2 7 1 0 9 1 9 7 0 9 0 9 2 1 15 15 9 15 9 13 2
8 13 13 9 2 7 0 9 2
24 7 3 13 13 0 9 7 9 1 9 2 7 13 7 9 9 2 9 0 9 1 0 9 2
19 13 3 0 9 1 9 0 0 9 7 1 9 9 2 3 13 10 9 2
2 9 9
2 11 11
19 0 9 7 0 9 13 0 2 9 13 1 9 7 9 2 15 3 13 2
20 2 13 15 12 2 9 12 1 11 2 13 9 0 9 9 0 2 9 9 2
7 13 0 2 13 12 9 2
6 2 9 0 9 11 2
40 2 1 9 10 0 9 13 16 9 2 3 13 16 0 9 2 9 2 3 15 13 0 9 9 9 1 9 9 1 9 7 9 1 0 12 1 0 0 9 2
13 1 9 12 13 9 0 9 7 13 15 10 9 2
20 13 1 9 0 9 11 2 15 13 0 9 9 9 7 13 15 10 0 9 2
6 2 13 0 9 9 2
20 13 0 0 9 2 0 9 9 7 9 1 9 2 9 9 7 9 2 9 2
28 10 9 1 0 9 0 11 13 1 0 9 9 1 9 0 1 9 11 2 0 0 9 1 12 1 12 9 2
19 2 13 0 9 0 2 0 7 0 2 13 1 10 9 1 9 7 9 2
14 13 15 15 2 15 15 13 13 7 9 13 16 9 2
18 13 13 2 16 1 9 10 9 13 16 9 0 9 2 9 9 2 2
8 1 9 13 2 16 13 3 2
21 11 11 13 3 0 2 7 2 0 9 2 0 15 1 9 13 15 1 9 0 2
3 9 13 11
8 0 9 2 14 1 0 9 2
3 13 0 9
9 0 9 13 0 13 1 0 9 2
26 1 0 11 9 13 14 1 9 9 0 7 0 9 2 15 15 13 3 9 9 2 9 7 0 9 2
21 13 4 15 15 1 15 1 0 9 2 7 3 1 0 9 1 9 1 0 9 2
21 11 11 2 9 2 11 2 14 3 4 13 0 9 1 9 2 15 13 1 0 2
16 9 9 9 1 11 4 13 12 0 9 2 15 13 0 9 2
33 9 0 0 9 2 15 0 9 3 13 1 0 11 7 1 0 11 2 13 16 0 16 9 9 2 15 4 13 1 11 7 11 2
5 3 9 13 0 2
26 3 1 9 3 13 1 0 9 7 4 2 14 15 9 13 2 13 2 16 15 1 10 0 9 13 2
24 11 11 2 11 0 2 9 2 2 11 2 1 11 4 3 3 13 0 9 2 3 0 9 2
20 1 0 9 13 0 9 1 9 0 9 7 9 2 3 3 0 9 1 9 2
14 0 9 13 9 9 2 16 10 9 15 13 1 12 2
23 16 15 1 9 13 3 9 1 9 1 9 9 2 3 4 15 13 3 1 0 9 3 2
20 1 11 15 13 1 0 9 13 9 0 9 11 2 15 4 13 13 9 9 2
19 0 9 4 13 2 16 4 10 0 0 9 4 3 3 13 1 0 9 2
14 13 15 0 0 9 1 11 2 1 9 9 7 3 2
18 3 4 15 13 3 9 13 9 2 13 0 9 13 9 1 0 9 2
17 13 4 15 9 0 9 2 15 13 0 2 13 4 15 3 9 2
16 11 11 2 11 2 11 2 0 9 4 3 3 13 3 3 2
14 13 0 9 1 9 0 0 9 2 3 13 3 0 2
13 13 15 15 3 1 9 9 2 3 1 9 9 2
14 1 0 9 13 13 10 0 9 1 9 0 9 9 2
14 3 1 9 1 12 9 15 13 9 3 1 12 9 2
11 13 3 14 1 12 0 9 1 11 3 2
21 13 4 15 1 9 0 9 2 15 4 13 13 14 1 11 2 7 3 1 11 2
16 10 9 13 3 3 0 7 3 9 0 9 1 0 9 13 2
20 11 11 2 11 2 12 2 11 2 3 4 13 0 9 3 1 11 7 11 2
16 13 4 9 1 9 0 9 1 11 2 7 9 13 3 0 2
20 0 0 9 13 3 0 13 3 1 0 9 1 0 9 2 3 1 12 9 2
7 9 13 3 1 9 9 2
24 16 15 0 9 3 13 2 13 12 9 9 3 7 1 9 9 13 4 13 3 9 1 9 2
9 13 15 7 13 1 0 0 9 2
20 3 4 13 2 16 13 0 9 1 9 2 15 13 3 1 9 7 1 9 2
19 13 15 15 15 1 0 0 9 2 3 0 9 1 0 13 14 3 0 2
13 1 15 9 1 0 9 4 13 10 9 1 9 2
14 3 1 11 13 3 0 9 9 2 9 13 3 0 2
4 0 11 2 9
4 13 0 9 2
5 1 0 9 3 13
18 14 12 9 1 11 1 11 1 11 13 0 9 1 9 0 9 11 2
21 1 0 9 13 1 9 14 12 0 9 2 0 9 1 12 9 1 11 1 11 2
3 11 7 9
17 1 11 11 2 9 9 2 13 1 9 9 0 9 7 0 9 2
10 9 13 3 2 3 15 13 0 9 2
8 1 9 11 13 9 10 9 2
4 2 0 9 2
14 9 13 1 9 1 0 9 7 9 15 13 0 9 2
41 7 1 9 0 9 2 0 15 1 12 2 12 5 2 13 9 9 3 1 0 9 16 1 9 2 16 4 15 15 7 13 13 3 9 3 7 14 1 10 9 2
4 2 0 9 2
8 13 0 16 9 0 0 9 2
9 0 9 13 1 9 12 0 9 2
21 15 13 1 9 14 14 12 0 9 2 7 9 13 1 10 9 13 12 12 9 2
25 3 13 9 0 9 12 9 2 15 0 9 2 1 15 13 0 9 9 2 14 1 12 9 3 2
4 2 0 9 2
6 11 13 9 14 3 2
18 3 1 9 2 3 13 0 13 9 9 1 9 7 9 1 0 9 2
20 3 13 3 3 13 9 1 9 2 16 4 13 0 9 9 7 0 0 9 2
14 13 3 1 9 0 2 15 9 9 13 3 0 9 2
4 2 9 9 2
10 0 9 13 1 9 12 2 12 5 2
16 10 9 13 1 0 9 7 1 9 2 15 15 13 1 9 2
6 1 0 9 13 9 2
17 1 0 9 12 5 2 0 12 5 13 9 13 2 16 13 3 2
9 0 9 13 9 1 9 0 9 2
10 1 9 13 13 2 13 15 9 11 2
11 13 1 0 9 9 7 13 15 13 9 2
1 9
7 9 9 13 9 1 9 2
23 9 13 13 1 15 2 16 15 15 1 15 1 0 9 3 9 13 2 7 1 15 13 2
15 9 9 15 9 9 0 11 1 0 9 13 12 9 9 2
13 1 0 9 15 13 0 9 2 13 15 9 11 2
14 7 16 13 1 15 0 9 2 13 9 10 9 13 2
16 13 13 7 10 9 10 2 16 4 15 13 10 0 0 9 2
7 9 9 13 3 7 3 2
10 0 9 1 9 0 9 13 0 9 2
22 13 4 15 1 0 9 2 16 4 1 9 1 9 13 1 0 9 2 13 15 9 2
10 0 9 13 2 13 7 1 0 9 2
11 9 1 9 7 10 0 9 15 15 13 2
14 3 7 9 15 4 1 0 9 10 9 13 0 9 2
2 11 11
22 9 2 11 2 9 0 9 2 0 12 2 12 12 11 2 9 2 2 2 12 2 12
5 2 9 1 9 2
4 13 3 13 2
5 13 9 7 13 2
10 10 3 0 9 13 13 13 9 9 2
24 1 9 2 16 15 13 1 9 2 13 9 1 0 7 0 9 7 10 9 13 1 0 9 2
9 0 9 13 0 3 1 10 9 2
4 9 1 0 9
10 1 9 12 4 13 1 9 1 9 2
24 1 9 9 1 11 1 11 1 15 13 2 16 4 15 13 0 9 7 13 10 9 1 11 2
13 13 4 9 1 0 9 2 9 15 7 13 13 2
9 3 15 1 11 13 9 0 9 2
15 13 4 1 15 2 7 4 13 1 9 0 9 1 11 2
12 3 4 15 13 2 16 4 1 9 13 13 2
7 9 1 9 9 7 13 2
4 13 15 13 2
5 13 9 1 9 2
4 9 9 2 12
47 1 1 15 2 16 4 13 1 9 0 9 1 9 2 4 4 7 13 1 0 9 0 9 9 1 0 1 9 9 9 2 7 10 9 13 1 9 9 1 9 3 3 0 9 0 9 2
13 1 0 9 4 15 1 15 13 9 1 0 9 2
36 16 4 10 9 13 1 9 1 0 9 13 2 13 4 3 2 16 4 13 14 0 2 7 3 0 9 2 7 13 7 0 9 1 9 11 2
17 3 13 1 10 9 2 9 9 4 3 13 2 9 9 7 14 2
8 1 10 9 4 13 0 9 2
12 1 0 7 0 9 1 0 9 15 13 13 2
6 9 2 9 2 11 11
25 9 2 0 7 3 0 9 2 0 12 2 11 12 2 9 2 5 9 2 2 12 2 12 12 2
3 11 13 13
5 9 3 13 9 2
5 11 15 1 11 13
11 1 12 9 13 3 13 9 0 11 11 2
13 1 9 2 15 13 12 12 9 2 13 15 3 2
22 10 0 9 13 1 9 12 0 9 2 15 13 12 9 2 7 0 9 12 9 11 2
10 1 9 13 9 2 1 9 9 9 2
2 11 11
14 9 15 3 0 9 13 2 7 10 9 13 3 0 2
12 1 0 9 4 11 3 13 9 1 0 9 2
8 0 9 13 14 12 9 3 2
14 9 1 0 9 13 1 12 2 12 9 9 1 11 2
2 3 11
10 9 15 3 1 11 13 3 1 11 2
10 1 0 9 3 13 12 5 15 9 2
18 9 15 14 3 13 1 9 0 9 2 1 15 13 1 9 0 9 2
10 13 3 11 2 15 13 0 0 9 2
16 1 0 12 9 0 9 13 1 11 3 16 12 9 0 9 2
9 1 0 9 11 15 13 12 9 2
11 9 9 1 9 0 11 3 13 12 5 2
13 1 0 9 15 7 13 13 14 12 9 9 3 2
18 0 9 13 9 2 16 3 0 9 9 1 12 9 13 9 3 13 2
10 13 10 9 2 16 15 15 3 13 2
28 0 9 13 1 11 11 2 12 5 2 2 3 13 11 7 9 2 1 12 5 2 7 11 2 12 5 2 2
11 0 9 1 11 1 0 9 13 0 9 2
20 1 9 2 3 13 9 9 2 13 1 0 9 13 1 0 9 9 7 9 2
3 9 7 9
9 9 0 9 4 3 3 3 13 2
23 9 9 1 9 12 9 2 15 1 9 12 13 12 9 1 9 2 13 1 9 15 13 2
12 0 9 13 0 9 2 15 13 3 10 9 2
18 0 9 9 13 3 1 9 1 12 9 2 9 9 1 9 3 12 2
25 1 9 9 13 9 1 0 9 1 12 9 3 16 12 9 2 1 9 3 3 1 12 9 3 2
9 0 9 13 9 1 9 0 9 2
13 9 11 13 1 9 9 9 3 1 9 7 9 2
16 9 9 1 9 1 0 9 7 1 0 9 13 14 12 5 2
8 1 0 9 13 12 9 9 2
19 0 13 1 0 9 2 0 13 1 0 9 7 0 13 1 0 0 9 2
13 15 13 1 9 1 12 9 1 9 1 12 9 2
3 15 9 13
13 1 9 9 13 1 11 0 0 9 1 12 9 2
7 3 13 15 1 9 3 2
6 3 15 3 13 3 2
37 16 1 0 9 9 13 9 1 11 1 9 12 7 12 1 12 9 3 2 1 9 12 2 3 4 13 3 10 9 2 15 13 3 16 12 9 2
18 0 9 2 15 13 1 9 14 12 9 2 13 9 3 1 12 9 2
8 9 4 15 13 1 0 9 2
16 0 0 9 13 1 9 9 3 12 9 1 9 1 0 9 2
15 13 15 10 9 7 9 9 13 13 3 1 9 0 9 2
13 1 10 9 13 1 11 15 9 1 9 0 9 2
12 3 1 0 9 13 3 13 0 9 9 11 2
9 0 9 13 1 9 9 12 9 2
13 9 1 11 15 13 13 7 13 9 1 12 9 2
1 9
19 1 9 0 9 13 1 9 0 9 9 0 9 1 9 1 0 0 9 2
18 1 9 4 1 11 13 3 16 12 9 2 0 1 0 9 12 9 2
16 15 9 2 15 13 0 12 5 0 9 2 4 13 0 9 2
8 9 0 9 13 13 1 9 2
30 13 15 1 0 9 0 9 2 7 1 15 7 1 0 9 2 16 9 11 13 1 3 0 9 0 11 7 0 11 2
4 0 2 11 2
13 7 1 0 9 9 13 3 10 0 9 3 13 2
9 9 2 9 9 1 11 1 0 9
15 9 1 9 0 2 1 9 1 9 13 4 0 9 3 2
5 9 2 13 4 13
2 9 9
10 9 1 15 13 9 1 9 0 9 2
11 3 15 2 9 2 13 1 15 10 13 2
5 11 11 2 0 11
30 0 9 15 1 9 2 0 9 0 9 2 2 7 3 7 1 0 9 2 1 9 13 9 2 15 13 9 3 13 2
8 9 7 9 13 13 0 9 2
12 9 13 1 9 2 10 9 1 9 4 13 2
9 0 9 13 1 0 9 9 9 2
27 3 13 9 15 2 16 13 9 2 1 0 15 13 7 9 1 0 9 13 0 0 9 2 3 0 9 2
20 9 13 13 7 0 9 10 9 2 0 0 9 1 0 7 0 9 7 3 2
16 0 9 0 9 13 0 9 2 9 2 9 2 9 9 2 2
27 9 9 13 0 0 9 9 2 1 15 14 12 1 0 12 9 9 1 12 9 7 9 4 1 9 13 2
27 1 9 9 3 13 2 16 15 1 15 2 16 13 9 13 2 13 2 13 1 15 9 2 7 0 9 2
17 9 2 0 0 9 7 0 9 13 4 1 9 11 13 1 9 2
38 13 2 14 15 13 9 1 9 1 9 0 9 2 13 4 13 3 9 0 7 0 0 9 0 9 1 0 11 2 7 9 1 9 7 9 1 11 2
29 13 15 15 2 13 2 14 15 1 9 2 9 2 9 9 2 13 4 13 13 1 0 9 7 0 0 9 2 2
31 3 15 13 13 1 9 2 16 13 9 13 0 0 9 2 15 4 13 7 9 13 2 16 13 1 3 0 7 0 9 2
2 11 11
5 1 9 15 9 13
4 9 1 0 9
6 13 1 0 0 9 2
9 1 0 9 15 9 3 13 13 2
13 7 15 13 2 16 15 12 9 13 9 3 12 2
9 12 1 15 13 0 2 0 3 2
21 9 10 0 9 3 13 15 2 16 13 7 13 3 9 2 15 15 10 9 13 2
9 13 4 9 7 13 15 1 9 2
19 0 9 4 13 2 3 3 13 0 2 1 9 0 2 0 9 1 15 2
4 7 9 9 2
13 9 9 2 10 0 9 3 13 0 9 0 9 2
11 13 13 2 13 9 2 13 7 4 13 2
26 3 14 2 7 1 15 2 15 3 13 3 7 3 0 0 9 2 13 9 1 9 15 3 0 9 2
18 3 2 1 9 1 0 0 9 7 9 13 9 3 2 7 3 0 2
2 9 2
16 2 13 15 13 0 9 2 1 15 13 13 9 3 0 9 2
28 2 13 2 14 9 1 9 10 0 2 1 9 2 9 2 13 10 9 3 3 2 16 13 9 3 0 9 2
5 11 11 2 0 11
22 9 0 1 10 9 2 0 1 0 9 9 2 4 3 13 7 3 13 9 12 9 2
10 4 3 13 1 0 9 1 12 9 2
19 13 15 1 15 2 10 9 4 15 1 9 13 7 10 1 15 13 9 2
2 9 9
15 3 12 12 9 9 11 13 1 0 9 1 9 0 9 2
33 13 15 1 1 0 9 9 1 0 9 9 2 9 0 9 2 12 9 1 9 12 2 2 7 7 9 9 9 3 1 9 9 2
24 0 9 13 13 10 9 13 2 16 1 0 9 3 1 0 9 9 13 1 9 7 10 9 2
13 9 0 9 1 0 9 15 3 13 1 12 12 2
4 9 7 9 9
8 0 9 0 9 1 0 0 9
21 1 9 0 9 9 13 9 9 0 0 9 2 11 2 1 11 0 9 0 9 2
34 3 12 9 9 2 9 9 2 0 7 0 9 7 9 15 13 12 9 3 0 1 9 2 9 9 9 7 9 0 7 3 0 9 2
2 11 11
21 1 9 13 3 1 9 9 0 9 2 3 1 9 9 2 1 15 15 9 13 2
17 9 13 16 0 9 0 9 0 1 0 9 2 9 2 0 9 2
37 9 7 9 2 15 13 1 9 0 9 9 9 2 13 3 13 1 0 9 2 9 15 1 10 9 9 13 1 9 2 14 3 1 9 0 9 2
15 16 15 3 9 2 13 2 2 13 3 1 9 0 9 2
6 9 13 1 9 9 2
21 0 9 9 13 3 0 7 7 3 3 0 2 3 9 0 9 7 9 0 9 2
31 10 9 3 13 9 0 9 2 3 0 2 13 9 13 9 9 1 0 9 2 1 9 9 9 13 9 2 13 1 9 2
6 9 15 13 0 9 2
39 13 9 2 16 13 15 9 9 1 12 9 13 0 9 2 7 13 0 13 15 15 7 1 0 9 2 7 15 13 9 2 1 15 15 4 9 3 13 2
25 16 9 1 9 9 9 1 9 13 0 9 9 2 13 15 3 9 13 1 15 2 3 13 0 2
15 1 9 13 9 2 0 9 2 15 7 9 9 3 13 2
25 1 9 1 9 0 7 3 0 9 13 9 2 16 9 13 9 9 7 9 1 0 9 0 9 2
6 13 15 3 16 0 2
15 7 9 13 1 9 1 0 9 3 1 9 9 7 9 2
11 7 3 3 3 13 1 9 7 9 9 2
18 1 9 13 13 3 0 9 13 15 1 9 2 15 13 9 3 9 2
14 13 15 2 16 9 10 9 13 7 9 1 0 9 2
43 13 3 12 0 9 2 1 12 9 15 13 9 2 15 13 7 13 10 9 13 2 3 9 13 1 9 7 9 1 9 2 2 1 0 9 9 9 1 0 9 3 13 2
15 0 4 3 13 0 9 9 1 9 2 3 1 0 9 2
22 9 4 13 7 3 13 9 0 0 7 0 9 2 15 13 1 9 0 7 0 9 2
34 9 2 0 0 9 2 15 2 12 2 9 12 2 12 12 11 2 9 2 2 2 12 2 12 2 12 2 9 2 2 12 2 12 2
5 12 2 7 12 2
20 1 9 9 9 2 12 1 9 1 9 0 9 13 16 0 9 9 12 9 2
19 1 0 9 9 7 4 13 1 12 9 2 13 15 10 9 1 0 9 2
5 13 15 7 15 2
37 16 3 13 3 7 0 2 13 2 16 9 12 9 13 0 9 13 14 1 9 12 1 9 0 9 1 9 12 2 7 1 9 12 13 12 9 2
2 10 9
2 9 9
8 2 9 9 2 12 2 12 2
12 16 9 9 13 0 2 13 15 15 3 0 2
25 7 15 13 12 9 9 2 15 4 13 10 0 9 2 16 4 15 1 0 9 13 1 0 9 2
17 13 15 2 10 9 2 10 9 2 2 13 4 15 14 0 9 2
16 7 15 3 13 2 16 15 9 13 9 2 16 4 15 13 2
11 13 4 15 3 13 2 13 10 0 9 2
15 13 4 9 1 0 0 9 7 3 4 9 13 0 9 2
24 13 15 9 7 0 9 2 7 16 13 1 0 9 0 1 0 9 2 13 15 0 9 9 2
15 0 9 4 3 13 1 9 9 1 9 2 9 0 9 2
16 9 1 9 2 2 9 7 11 2 2 13 2 9 7 11 2
33 13 0 2 16 0 9 9 1 10 9 3 13 2 7 13 13 2 16 15 13 1 0 0 9 3 2 16 15 13 13 9 9 2
6 7 15 13 9 9 2
5 9 13 13 9 2
8 11 7 11 11 2 11 1 11
2 0 9
8 2 9 9 2 12 2 12 2
9 13 1 9 14 12 9 1 9 2
5 13 3 0 9 2
38 1 0 9 7 1 0 9 1 9 9 1 0 0 9 7 0 9 1 15 1 0 9 2 7 15 0 9 9 9 4 15 1 10 9 13 0 9 2
24 16 4 13 9 9 2 13 4 1 0 9 1 0 9 12 9 12 3 12 0 9 0 9 2
23 1 9 1 9 1 10 9 4 13 13 1 9 9 0 9 1 9 12 2 12 2 9 2
39 1 9 10 12 9 2 13 2 14 0 9 9 1 0 9 2 13 1 9 0 9 7 1 9 9 12 9 9 9 12 9 2 0 9 4 3 13 2 2
21 9 2 15 13 0 9 1 0 0 9 2 10 9 13 7 3 13 3 0 9 2
11 3 4 1 0 9 13 1 9 0 9 2
12 13 9 0 9 2 15 15 13 0 9 9 2
17 0 9 13 9 9 1 3 0 9 2 3 3 1 9 9 9 2
21 1 0 9 15 15 13 2 16 9 13 0 1 9 2 1 15 15 9 13 13 2
18 3 13 9 13 9 9 2 15 15 13 13 14 9 2 14 3 9 2
8 3 13 9 13 3 1 9 2
18 15 13 3 0 2 16 9 15 13 2 7 1 9 1 9 0 9 2
11 0 9 4 14 13 7 1 9 7 9 2
21 13 15 7 13 3 0 9 1 0 9 2 3 13 3 9 2 1 9 1 9 2
7 0 9 13 0 0 9 2
15 16 13 13 0 9 2 13 9 13 7 3 13 1 9 2
22 16 13 10 9 9 1 9 0 2 13 1 15 1 0 9 0 7 13 1 15 0 2
5 11 11 2 0 11
3 3 7 3
8 2 9 9 2 12 2 12 2
7 13 0 9 1 11 3 2
10 3 15 13 14 3 0 2 13 3 2
15 10 9 15 3 13 2 3 15 13 9 7 3 7 9 2
8 3 1 0 9 13 0 9 2
18 16 15 13 14 3 0 9 2 9 15 13 3 0 7 13 15 0 2
29 0 9 13 9 9 15 2 16 0 13 3 1 0 9 7 13 13 7 9 1 9 1 0 9 7 9 1 9 2
19 1 15 3 15 13 2 3 3 15 3 13 2 16 4 15 0 13 3 2
23 13 4 1 9 9 2 12 1 9 1 9 2 13 9 2 13 2 1 9 7 15 15 2
4 9 13 0 2
10 13 4 15 1 0 7 9 15 13 2
6 14 0 13 1 9 2
33 0 9 15 7 13 2 16 0 13 0 1 15 2 16 9 3 13 2 7 7 13 15 9 1 9 2 16 1 15 9 3 13 2
39 7 13 15 12 2 16 15 1 0 9 13 2 3 15 13 2 3 15 1 15 13 12 9 7 3 1 15 13 9 2 7 0 9 15 13 1 0 9 2
4 11 11 2 11
7 13 4 15 15 2 3 9
8 2 9 9 2 12 2 12 2
19 1 10 9 15 9 9 13 0 9 2 15 13 14 1 9 9 1 9 2
22 0 9 1 9 1 9 15 2 9 2 13 9 7 9 0 9 2 7 3 0 9 2
17 13 10 9 10 9 13 2 7 15 13 2 16 0 9 13 3 2
8 3 3 0 0 9 0 9 2
10 0 9 9 13 9 2 9 9 3 2
11 7 15 3 13 14 10 9 2 3 3 2
13 9 9 13 2 16 9 10 9 13 3 14 9 2
5 7 15 13 9 2
35 10 0 9 13 0 7 13 7 10 0 9 2 15 9 13 3 3 1 9 7 3 2 9 1 15 3 13 0 9 1 9 10 12 9 2
5 0 3 13 13 2
21 15 2 15 15 13 0 9 13 2 13 14 13 2 16 4 1 10 9 3 13 2
11 7 15 10 9 3 13 13 1 12 9 2
10 13 1 15 3 0 2 3 7 0 2
16 13 3 2 16 9 13 2 15 1 15 4 13 7 15 13 2
9 13 9 14 1 9 13 3 0 2
12 14 4 3 3 13 1 9 7 9 1 9 2
4 11 11 2 11
3 9 11 3
34 3 9 9 15 13 1 0 0 9 9 11 2 15 1 0 9 9 13 1 9 12 2 2 12 2 9 9 1 9 9 7 9 11 2
9 9 4 13 1 12 0 0 9 2
27 0 13 0 7 0 9 2 16 9 0 9 2 9 1 9 9 2 9 1 0 9 2 9 9 7 3 2
9 0 13 13 1 9 3 0 9 2
29 1 0 9 9 11 13 3 9 0 9 1 0 9 2 3 9 3 0 9 2 1 15 13 9 9 0 9 11 2
5 11 11 2 9 2
14 11 2 11 5 11 2 9 2 9 2 0 2 2 11
11 1 0 9 1 11 4 15 13 3 3 2
13 9 11 13 1 9 9 7 9 0 1 0 11 2
14 10 9 13 7 0 0 9 1 0 9 9 0 9 2
26 1 9 0 9 13 3 7 0 9 9 11 10 0 9 0 9 2 9 9 0 9 7 0 0 9 2
13 0 11 4 15 16 9 13 1 0 9 10 9 2
8 12 9 15 13 3 3 13 2
22 9 1 11 15 13 1 2 16 0 9 9 7 9 1 9 15 15 13 13 3 3 2
12 1 9 13 1 9 1 9 0 9 3 0 2
26 13 0 2 16 1 9 9 11 13 2 16 13 1 15 2 3 15 13 9 7 3 15 13 9 2 2
22 1 10 9 0 0 9 9 13 1 10 9 7 13 15 2 16 9 13 15 1 15 2
6 3 13 9 0 9 2
9 1 10 9 13 11 13 0 9 2
10 1 0 9 9 13 1 11 3 0 2
14 13 4 15 7 2 16 4 9 9 9 13 0 0 2
17 3 13 1 15 9 2 15 15 13 2 16 13 13 14 1 9 2
15 16 13 1 9 13 15 1 9 9 2 7 15 3 13 2
21 3 9 9 13 2 16 1 0 9 13 1 0 9 2 15 4 13 1 10 9 2
22 7 16 0 13 7 9 1 9 2 16 10 9 13 0 2 7 15 14 2 13 2 2
12 13 13 9 2 15 15 1 15 13 1 9 2
13 13 9 2 16 15 2 0 11 2 13 15 13 2
19 15 3 12 9 13 12 10 9 0 9 2 16 1 15 0 9 15 13 2
7 3 7 14 10 0 9 2
10 9 13 0 9 2 16 13 0 9 2
18 15 13 13 1 11 0 7 0 9 2 1 15 4 13 9 12 9 2
32 0 9 15 3 13 2 7 9 13 3 1 9 2 1 15 15 3 3 13 2 7 1 15 2 15 13 1 0 9 0 9 2
7 13 15 0 9 0 9 2
16 9 1 0 9 1 0 9 7 9 1 9 13 7 10 9 2
20 1 0 9 15 13 2 16 10 0 9 13 0 9 9 2 1 15 13 0 2
9 13 15 7 9 9 7 9 9 2
12 3 13 13 9 7 9 9 1 9 0 9 2
3 9 1 9
9 0 9 2 9 13 3 0 9 9
29 1 0 9 12 13 9 1 9 0 9 1 9 9 0 3 0 9 1 9 2 7 0 7 16 9 0 0 9 2
29 1 15 2 16 1 10 9 9 9 13 3 7 0 9 2 13 9 0 9 11 2 1 9 0 9 13 0 9 2
2 11 11
15 11 15 13 9 0 9 2 0 9 7 0 9 1 15 2
27 0 9 2 15 13 13 0 1 9 9 2 13 1 9 13 0 9 0 1 9 2 13 9 9 1 15 2
14 7 1 9 13 7 0 9 2 13 13 0 9 9 2
2 0 9
11 1 15 9 9 3 12 5 12 9 13 2
10 3 2 9 9 13 13 14 1 9 2
24 13 13 7 13 10 9 2 9 9 2 15 13 7 3 13 0 9 2 3 13 4 9 13 2
21 0 9 2 1 10 9 7 9 0 9 15 11 13 2 13 13 9 7 1 9 2
13 3 4 13 12 9 0 9 2 0 1 0 9 2
14 0 13 3 0 13 3 2 1 0 9 1 12 9 2
20 0 9 13 13 15 2 15 13 3 0 7 13 12 9 2 7 13 12 9 2
7 0 13 0 9 12 9 2
11 15 9 9 13 9 0 9 1 11 3 2
7 15 13 0 9 9 9 2
9 3 7 1 10 9 13 9 9 2
5 15 1 15 13 2
9 9 0 9 13 9 9 0 9 2
12 13 15 3 3 13 9 9 9 1 10 9 2
11 13 3 9 13 9 15 9 1 10 9 2
23 13 9 2 16 13 15 3 3 15 13 2 7 16 9 9 1 12 9 13 1 9 9 2
24 9 15 13 2 16 13 13 9 2 13 1 0 9 3 9 1 9 7 0 9 7 13 9 2
18 3 1 9 15 13 7 1 9 2 0 15 1 9 2 13 3 9 2
19 7 9 13 13 9 2 16 15 1 9 3 13 2 16 15 13 1 9 2
11 9 15 3 13 13 1 0 9 0 9 2
24 13 9 2 16 3 4 13 13 0 2 16 13 0 0 9 2 16 4 15 13 10 0 9 2
11 3 15 7 13 13 1 9 7 0 9 2
23 12 1 9 13 1 9 9 0 1 9 1 9 0 9 2 15 13 9 10 0 0 9 2
23 13 15 7 0 9 1 10 9 2 7 15 13 13 1 10 9 7 9 9 1 9 9 2
3 9 1 9
16 0 9 9 13 9 2 15 15 7 13 9 7 0 9 9 2
28 3 15 3 13 10 0 9 1 10 9 2 7 3 9 13 1 10 9 3 14 3 1 10 0 2 9 2 2
10 1 0 9 13 9 9 7 9 9 2
10 1 0 9 7 9 0 9 9 9 2
19 3 0 9 1 0 9 13 1 0 9 9 2 1 15 4 13 13 9 2
17 9 4 3 13 0 9 9 2 15 13 3 3 13 1 9 9 2
10 7 1 10 0 9 13 9 0 9 2
12 3 13 9 9 2 13 0 9 9 1 15 2
24 3 1 0 0 9 9 10 9 13 9 3 0 9 1 0 9 9 7 1 9 13 1 9 2
8 7 3 10 9 13 9 9 2
9 1 11 13 3 9 9 0 9 2
12 0 9 13 10 9 2 15 13 13 1 9 2
7 15 13 0 9 9 9 2
18 9 3 13 3 9 3 3 10 9 2 9 9 13 2 10 9 13 2
12 13 3 2 16 15 1 9 13 1 9 13 2
17 9 3 13 13 2 16 9 13 1 9 9 2 7 13 13 9 2
41 7 16 3 9 9 9 13 0 9 1 0 9 2 13 3 3 13 1 9 2 0 9 13 13 12 1 9 0 3 9 1 0 7 0 2 3 7 10 0 9 2
14 3 0 9 13 13 0 2 7 16 3 0 2 9 2
32 9 2 11 2 0 12 2 12 12 11 12 2 9 2 2 2 12 2 12 12 2 9 2 5 9 2 2 12 2 12 12 2
4 9 1 9 2
4 9 7 9 2
22 14 15 1 9 9 13 13 2 16 10 9 13 0 7 1 9 0 3 1 9 9 2
9 7 1 15 9 1 0 9 13 2
5 12 11 1 0 9
12 1 0 13 1 9 9 2 0 9 13 1 9
16 12 11 1 0 9 2 3 12 0 0 9 2 13 0 9 2
20 12 13 1 0 9 2 3 15 13 0 9 10 2 3 3 0 2 0 9 2
16 12 15 3 13 1 9 0 0 9 1 0 0 7 0 9 2
25 11 11 2 9 0 9 1 0 9 2 13 1 15 3 2 16 10 0 0 9 1 11 1 11 2
19 1 0 9 1 9 12 7 12 15 13 1 9 7 13 3 0 0 9 2
8 1 15 0 15 13 0 9 2
18 3 1 9 11 13 9 0 9 2 3 13 12 5 9 2 0 9 2
9 3 3 12 9 13 16 13 9 2
4 11 3 1 9
19 1 0 12 9 13 0 9 0 9 2 0 0 9 2 10 9 9 9 2
12 9 13 12 9 2 1 15 13 12 0 9 2
15 1 0 9 15 13 9 1 9 15 2 7 15 3 9 2
10 13 3 9 2 9 7 9 0 9 2
11 0 9 1 0 12 9 13 9 1 0 2
19 1 9 12 3 13 12 9 2 12 9 7 0 9 1 3 12 9 9 2
7 0 9 13 12 9 9 2
14 3 15 13 12 9 7 0 9 13 1 12 9 9 2
16 13 15 2 10 13 9 2 16 15 3 3 13 1 0 9 2
8 9 13 9 11 11 11 11 2
8 13 15 0 9 2 7 13 2
27 13 2 14 13 1 0 2 7 3 3 0 9 2 13 15 13 0 0 9 7 3 15 1 0 9 13 2
21 16 13 1 0 9 2 16 9 0 9 13 1 10 9 1 9 3 2 3 13 2
19 0 9 13 9 7 0 10 9 13 9 0 9 1 9 1 0 0 9 2
27 0 9 13 11 2 11 2 11 2 11 7 3 11 2 13 15 13 9 1 9 0 0 9 7 1 11 2
12 1 9 10 9 3 13 14 12 9 0 9 2
15 0 0 9 3 13 0 9 7 9 1 9 10 0 9 2
4 3 13 9 2
9 3 3 1 9 13 1 9 9 2
8 9 1 9 9 13 10 9 2
9 3 13 1 0 9 3 3 12 2
29 0 9 0 9 11 11 13 9 12 9 7 11 11 1 9 11 11 2 9 9 9 2 9 12 9 12 12 9 2
21 9 9 1 9 0 9 7 10 9 13 9 13 11 11 11 2 11 7 10 9 2
9 15 7 3 13 12 1 9 9 2
20 10 9 13 3 0 9 1 9 12 9 2 15 9 11 13 1 9 0 9 2
26 11 11 15 13 1 9 3 1 9 1 9 0 9 7 10 9 2 7 16 3 13 2 3 1 9 2
8 15 13 1 0 9 9 13 2
14 9 0 9 3 13 1 11 11 7 9 2 0 9 2
5 1 11 1 9 9
11 0 9 13 9 1 9 2 7 14 1 9
14 3 0 9 13 1 12 9 3 1 11 11 1 11 2
17 1 9 0 9 13 9 0 9 1 12 12 9 9 3 1 12 2
9 1 9 13 1 12 0 12 9 2
23 14 15 3 10 9 13 1 9 2 0 9 7 3 15 13 9 1 9 7 3 13 9 2
10 3 15 10 9 13 1 12 9 9 2
17 1 10 9 15 13 3 1 12 9 2 0 1 10 0 0 9 2
13 3 15 13 13 9 9 7 13 13 9 1 9 2
27 13 0 9 1 11 2 13 15 13 15 9 0 9 7 13 15 3 3 13 2 7 16 3 1 9 9 2
18 9 9 13 0 9 2 11 2 11 2 7 1 9 15 13 0 9 2
18 15 4 3 13 1 9 9 9 1 0 9 7 13 1 0 0 9 2
5 0 9 2 0 9
14 1 9 1 0 9 4 13 9 0 9 11 11 9 2
11 2 1 10 9 13 1 9 1 0 9 2
33 0 9 13 9 7 15 0 15 9 13 9 1 10 2 16 13 3 13 11 14 16 15 2 7 3 1 11 7 0 9 11 11 2
15 11 15 3 13 15 1 9 11 7 15 13 1 9 15 2
17 1 9 12 4 13 0 9 11 2 15 13 0 9 9 0 11 2
7 9 9 13 9 0 9 2
14 3 13 3 0 9 7 9 16 13 0 9 7 3 2
9 2 3 13 0 9 10 0 9 2
13 13 15 2 16 3 14 1 10 9 13 0 9 2
26 1 9 15 13 0 9 1 9 3 15 13 7 3 4 3 1 12 9 13 10 9 12 1 12 9 2
20 13 9 12 1 0 2 9 0 9 2 7 7 0 9 1 9 12 9 0 2
11 10 9 4 13 4 13 1 9 3 3 2
7 2 13 3 1 0 9 2
10 3 13 9 0 9 7 9 9 11 2
5 4 13 0 9 2
13 9 0 9 13 9 2 1 15 10 9 4 13 2
13 13 4 13 9 0 9 2 3 15 0 9 13 2
9 13 7 2 16 4 13 10 9 2
5 3 4 13 9 2
6 2 15 13 0 9 2
5 4 13 0 9 2
21 1 0 13 9 11 11 2 15 1 9 0 11 13 11 16 9 1 0 0 9 2
14 2 13 1 15 0 9 10 0 9 1 9 0 9 2
5 9 13 1 9 2
15 10 0 9 13 13 9 1 9 2 3 1 0 0 9 2
23 0 9 4 11 13 1 0 9 2 0 9 13 13 9 1 9 7 3 3 1 0 9 2
19 1 9 7 13 2 16 13 3 0 13 1 11 1 0 9 0 0 9 2
15 7 0 9 7 0 0 9 13 13 1 9 3 0 9 2
15 13 2 16 0 9 13 13 9 3 2 16 4 13 0 2
3 0 9 9
14 1 12 9 15 3 3 13 9 10 9 1 0 9 2
8 13 3 9 7 9 1 9 2
40 1 0 0 9 13 3 15 1 9 2 3 7 13 0 9 7 9 1 0 9 9 2 9 7 9 2 1 9 9 2 15 1 10 9 0 7 0 9 13 2
7 1 9 7 0 9 13 2
29 9 11 2 0 9 9 2 2 9 2 9 2 0 2 2 15 13 10 9 1 11 1 0 11 2 3 1 9 2
67 0 9 9 7 9 1 9 7 0 0 9 13 9 9 2 1 0 9 9 13 7 9 1 0 9 2 16 13 10 9 9 2 13 15 15 2 3 2 0 9 2 3 2 2 7 3 9 2 15 13 9 9 0 9 2 13 13 7 1 9 1 0 9 10 9 13 2
17 7 3 2 16 0 9 13 0 9 9 13 3 16 1 12 9 2
4 9 2 9 9
8 0 9 2 12 2 12 2 9
11 9 1 10 9 13 9 3 1 0 9 2
15 9 13 1 9 1 9 0 9 0 1 9 9 10 9 2
3 0 7 0
18 9 9 7 9 9 1 9 0 9 1 11 1 11 13 1 0 9 2
19 1 9 0 9 13 9 0 9 0 9 11 11 2 15 4 13 1 9 2
17 2 13 3 0 9 2 15 13 9 1 12 9 9 1 0 9 2
9 13 1 15 7 0 9 16 0 2
13 13 13 2 16 10 9 13 7 0 9 10 9 2
14 3 13 4 0 0 9 13 1 0 9 3 1 9 2
8 3 15 13 1 9 0 9 2
38 0 9 1 11 4 13 0 9 1 9 9 2 16 4 13 0 9 9 2 9 2 3 0 9 2 0 7 3 3 0 9 2 9 9 9 7 3 2
10 2 3 13 9 1 10 9 9 9 2
22 9 13 1 0 9 12 9 9 9 2 15 13 1 9 0 9 9 1 12 12 9 2
9 9 7 13 1 9 3 1 9 2
12 15 13 2 16 1 0 0 9 4 9 13 2
17 2 9 13 1 9 3 3 2 16 13 1 0 0 9 0 9 2
9 9 1 9 3 13 3 9 9 2
16 13 7 13 2 16 0 9 13 0 0 9 7 9 0 9 2
8 3 2 0 9 13 0 9 2
17 0 9 3 13 13 1 9 7 9 2 15 13 0 1 9 9 2
16 9 0 0 9 7 9 1 9 0 9 15 3 13 1 9 2
5 10 9 4 13 2
25 2 13 15 1 15 2 16 9 0 9 2 0 9 0 11 2 13 0 9 1 11 13 0 9 2
6 13 15 1 0 9 2
16 13 13 9 1 0 9 1 0 12 9 1 12 7 12 5 2
13 13 3 0 9 1 11 7 10 0 9 13 13 2
23 13 3 2 16 1 0 11 15 13 9 9 9 2 15 1 0 0 9 13 7 0 9 2
12 9 9 13 13 9 2 15 13 13 15 9 2
7 3 13 10 9 12 5 2
6 2 13 0 9 9 2
13 13 9 2 16 1 0 9 15 3 13 9 9 2
24 1 0 9 7 13 13 9 1 0 7 0 9 2 9 7 0 9 2 15 4 13 0 9 2
9 3 13 9 10 9 3 1 9 2
3 9 1 9
5 9 9 7 9 2
4 9 13 0 9
21 9 11 15 3 13 2 1 9 2 10 0 9 7 13 15 1 9 13 0 9 2
12 1 0 9 7 0 9 7 13 7 0 9 2
17 0 9 2 9 7 9 15 13 10 9 14 1 9 9 7 9 2
22 9 9 11 0 15 13 13 0 9 1 10 9 2 15 15 9 10 0 9 3 13 2
2 11 11
23 1 0 12 9 2 15 1 11 2 11 13 1 3 0 9 2 9 13 1 9 14 3 2
15 13 0 9 1 0 9 7 3 13 0 9 10 0 9 2
3 9 1 9
15 1 15 0 3 13 13 9 9 7 9 2 13 11 9 2
6 15 13 9 1 9 2
22 0 9 2 15 3 9 9 13 2 13 2 13 15 2 9 2 9 9 15 13 13 2
22 13 1 15 3 0 9 9 1 9 7 3 9 9 9 2 9 9 7 0 0 9 2
9 9 11 13 3 1 10 9 3 2
12 9 13 13 1 9 2 0 1 15 13 9 2
17 0 9 7 9 2 15 13 2 15 13 1 0 9 9 7 9 2
19 9 1 10 9 7 10 9 3 13 2 7 15 13 13 13 7 1 9 2
15 13 3 1 10 9 2 1 9 9 13 9 13 0 9 2
9 0 9 13 1 0 9 0 9 2
13 1 12 9 15 9 13 3 1 12 9 1 9 2
26 0 9 7 9 15 13 9 2 1 15 4 13 9 1 9 9 1 9 2 0 9 7 0 0 9 2
13 1 15 7 1 9 13 9 2 9 1 9 2 2
5 15 15 15 13 2
20 15 2 3 13 9 0 13 2 16 1 15 9 13 9 7 1 10 0 9 2
21 3 13 0 2 16 14 13 2 16 15 15 9 13 2 7 15 13 15 1 15 2
6 9 10 9 13 13 2
17 1 0 0 9 13 1 0 9 0 9 2 10 9 9 13 3 2
3 0 0 9
28 9 9 3 13 2 16 9 13 9 1 9 3 1 15 2 10 1 9 13 9 2 15 1 15 9 13 3 2
17 9 1 9 9 2 0 9 0 9 7 0 9 2 15 13 9 2
35 1 0 9 13 9 13 9 9 9 3 7 3 1 9 2 3 15 0 9 13 1 10 9 9 2 13 1 9 0 0 9 3 1 9 2
7 10 9 4 9 13 3 2
14 13 2 14 9 0 0 9 2 9 15 13 0 9 2
8 3 13 7 9 9 7 3 2
21 1 0 9 2 3 0 2 13 9 9 1 9 7 1 9 15 13 7 0 9 2
12 1 0 9 1 0 9 9 13 9 0 9 2
15 1 0 0 0 0 9 7 0 9 1 9 13 0 9 2
11 13 2 14 15 15 2 13 13 9 9 2
11 13 15 2 16 1 9 9 13 10 9 2
17 1 9 9 4 15 3 13 1 9 12 7 12 9 1 12 9 2
9 15 4 7 0 9 9 13 13 2
7 7 13 3 15 9 13 2
15 10 9 2 9 0 7 0 9 2 13 0 1 9 9 2
17 7 0 9 1 9 9 13 0 0 9 2 15 1 15 13 9 2
6 3 13 9 14 0 2
23 3 2 16 1 0 9 9 13 9 9 9 7 13 9 0 9 2 13 9 1 10 9 2
16 16 7 16 3 0 9 13 0 9 2 9 3 13 0 9 2
3 2 9 2
8 0 9 2 3 13 2 13 2
19 9 15 3 13 13 14 1 9 0 7 0 9 7 13 9 1 0 0 9
6 2 9 1 9 2 2
15 0 0 9 13 2 3 0 13 0 9 7 9 1 9 2
8 0 9 1 0 9 9 13 2
37 9 2 11 2 9 2 9 2 0 2 2 0 12 2 12 12 11 12 2 9 2 2 2 12 2 12 12 12 2 9 2 2 12 2 12 12 12
3 9 2 9
3 9 1 9
9 7 12 5 9 13 13 9 0 9
20 9 1 9 9 4 13 13 0 9 2 16 15 13 9 2 16 15 0 13 2
22 0 9 4 15 3 13 13 1 9 0 9 2 3 10 2 15 13 9 9 0 9 2
40 15 15 13 9 9 0 9 11 2 11 7 11 7 9 0 0 9 11 2 11 11 2 15 4 13 2 16 4 13 9 2 15 4 13 13 0 9 0 9 2
26 15 13 0 9 1 15 2 16 4 9 1 10 0 9 2 3 15 13 10 9 2 13 9 1 9 2
31 1 0 9 13 0 2 16 4 0 9 13 0 9 1 9 15 1 9 2 3 13 9 2 3 13 1 9 9 7 3 2
7 7 15 13 3 0 9 2
17 1 9 2 15 13 9 9 11 2 13 9 9 0 9 3 0 2
25 3 0 9 1 9 9 9 13 12 12 12 9 7 1 0 0 9 7 13 14 12 7 9 9 2
30 13 2 14 9 9 3 9 9 2 3 9 0 9 2 15 15 13 1 12 7 12 9 2 13 12 7 12 12 9 2
12 16 4 9 13 12 9 2 13 12 9 3 2
31 7 9 3 13 13 15 9 2 15 13 9 9 2 9 2 9 9 7 3 1 9 15 13 13 9 9 2 3 9 13 2
22 7 15 0 13 9 9 2 15 3 15 13 13 13 0 9 1 9 1 0 0 9 2
22 13 15 13 3 2 16 10 9 13 3 1 9 0 9 2 16 15 15 15 3 13 2
18 1 15 2 16 13 13 1 9 2 15 1 10 9 13 0 9 9 2
15 3 0 0 9 1 9 7 9 9 1 9 1 0 9 2
9 13 15 7 3 1 0 9 13 2
21 16 13 1 0 9 7 15 9 1 15 0 2 13 15 15 13 7 13 9 15 2
15 1 9 15 1 9 0 9 13 3 12 5 1 0 9 2
21 13 1 10 0 9 11 9 2 13 2 14 15 2 16 9 4 13 7 9 9 2
5 15 0 15 13 2
13 10 9 13 13 14 15 2 15 13 13 0 9 2
15 1 0 9 1 9 11 15 13 3 12 9 1 9 0 2
17 16 15 13 13 9 0 9 1 9 9 2 13 15 13 10 9 2
7 13 3 1 9 1 9 2
26 13 15 13 0 9 2 0 9 2 9 1 9 9 2 13 2 14 15 1 9 2 2 3 0 9 2
12 3 15 13 13 0 9 7 9 1 9 9 2
14 9 13 13 0 12 9 7 13 15 1 15 0 9 2
30 16 9 10 0 9 13 2 13 15 15 1 15 13 2 7 13 13 1 15 2 16 0 9 9 10 9 13 12 9 2
21 0 9 2 3 0 9 2 13 0 7 13 1 0 9 2 15 15 13 3 3 2
12 1 3 3 15 13 0 9 13 3 0 9 2
16 13 2 14 15 1 9 2 3 13 15 12 9 7 12 9 2
4 3 12 9 2
26 13 2 14 7 1 10 9 2 13 15 9 2 16 9 4 3 13 7 13 1 9 9 1 10 9 2
20 13 15 7 9 2 3 0 9 13 9 1 9 2 16 13 1 0 0 9 2
26 9 4 15 13 13 13 2 3 13 0 9 13 7 15 1 15 13 13 2 16 4 15 13 3 3 2
20 9 0 9 13 13 0 9 1 9 9 7 9 9 2 3 4 13 0 13 2
39 1 9 2 15 13 3 9 9 2 1 15 15 9 3 13 7 0 9 2 1 15 4 15 4 13 1 10 9 2 15 3 13 1 9 1 3 0 9 2
1 9
5 9 2 9 2 9
10 2 9 2 0 9 7 9 9 9 2
33 9 2 11 2 9 2 0 12 2 12 12 11 12 2 9 11 2 9 2 2 2 12 2 12 12 2 9 2 2 12 2 12 12
16 2 9 2 0 9 9 7 9 9 2 3 1 9 7 9 2
13 9 2 12 2 12 2 2 12 2 12 2 12 2
8 2 9 2 3 0 9 9 2
13 9 2 12 2 12 2 2 12 2 12 2 12 2
8 9 2 12 2 12 2 12 2
32 9 2 11 2 9 2 9 2 0 2 2 0 12 2 12 12 11 12 2 9 2 5 9 2 2 12 2 12 12 2 12 2
45 2 9 2 0 9 2 9 9 9 2 0 9 9 2 9 0 9 2 0 9 2 0 9 9 9 2 0 9 9 7 0 9 2 9 9 1 9 9 2 0 9 7 0 9 2
2 12 2
32 9 2 11 2 9 2 9 2 0 2 2 0 12 2 12 12 11 12 2 9 2 5 9 2 2 12 2 12 12 2 12 2
6 9 1 9 0 9 2
3 0 0 9
3 0 0 9
4 0 9 7 15
2 11 11
22 9 0 9 11 11 13 1 9 0 9 2 3 13 11 11 1 11 9 1 0 9 2
36 1 9 15 13 1 0 0 9 2 15 13 3 0 0 9 2 0 9 2 1 0 9 7 0 9 2 7 0 9 2 3 0 9 7 9 2
13 1 9 1 12 9 9 13 9 9 1 12 5 2
12 13 12 9 7 10 9 13 1 12 9 9 2
20 1 0 9 13 11 2 0 11 7 11 2 1 15 9 13 12 5 15 9 2
14 1 0 11 1 11 13 9 11 11 1 9 0 9 2
16 1 9 1 11 13 9 12 9 9 11 7 11 7 9 11 2
25 3 15 1 0 9 13 0 9 7 9 11 7 11 2 15 15 13 13 1 0 9 7 0 9 2
42 1 0 12 9 13 1 0 9 0 12 7 12 9 2 15 13 0 0 9 2 3 3 13 9 7 9 2 13 11 11 2 9 11 11 1 0 11 2 1 9 2 2
13 9 13 1 12 9 13 1 0 9 3 9 9 2
34 9 2 11 11 11 11 2 0 12 2 12 12 11 12 2 9 2 2 2 12 2 12 12 12 2 9 2 2 12 2 12 12 12 2
4 9 2 0 9
3 3 13 9
20 9 3 13 0 2 7 1 1 15 2 16 13 9 3 0 2 13 0 9 2
11 9 1 10 9 7 9 13 3 3 0 2
16 16 13 13 0 9 7 9 9 2 13 9 13 7 3 3 2
14 13 4 15 1 9 2 1 15 15 13 9 1 9 2
15 1 9 13 0 0 9 7 15 13 0 9 0 0 9 2
16 3 1 9 13 0 9 2 9 2 3 7 9 7 0 9 2
11 13 15 9 0 2 0 2 0 7 0 2
16 9 15 3 13 2 0 9 13 0 9 2 3 15 3 13 2
21 16 4 1 9 13 9 2 13 4 1 14 0 9 2 1 9 1 9 0 9 2
8 3 4 9 13 1 0 9 2
16 15 13 9 13 2 3 1 9 13 0 9 13 7 13 0 2
6 11 11 2 11 1 11
14 0 9 0 1 10 9 13 3 0 9 7 0 9 2
11 4 3 12 3 13 1 9 1 12 9 2
26 13 14 9 2 15 4 13 1 10 0 9 2 7 7 10 2 1 15 15 9 2 9 13 16 9 2
3 0 16 9
9 0 11 13 0 9 1 0 9 11
15 9 1 0 11 13 1 11 11 0 9 2 7 0 9 2
13 1 9 0 7 0 9 13 0 9 7 0 9 2
9 13 15 7 13 3 3 0 9 2
2 11 9
27 1 0 9 1 10 0 9 7 9 13 0 9 1 0 9 0 9 1 0 9 2 0 9 11 11 9 2
29 1 9 4 1 11 13 0 9 11 9 2 1 15 13 9 12 9 2 0 12 9 4 13 1 11 1 0 9 2
2 13 9
23 11 2 11 2 11 2 11 7 0 0 9 13 0 9 7 7 13 9 1 11 1 9 2
6 0 9 7 11 13 2
17 13 9 13 15 15 2 15 9 3 13 2 1 0 9 0 9 2
10 1 15 4 10 9 7 9 13 0 2
6 9 15 13 15 9 2
11 3 4 13 1 9 9 1 0 9 9 2
20 9 13 9 9 9 1 9 13 9 1 9 11 12 2 13 0 9 11 9 2
8 0 15 13 9 0 0 9 2
19 11 13 3 1 9 0 9 1 9 7 9 9 2 3 16 1 10 9 2
13 7 15 13 13 9 1 9 9 14 1 0 9 2
11 3 4 9 13 9 1 9 7 1 9 2
12 3 15 13 1 9 9 0 9 9 0 9 2
11 9 13 13 0 0 9 7 9 0 9 2
10 1 0 9 13 9 13 7 13 9 2
30 1 9 9 13 3 3 13 0 9 2 15 10 9 3 13 7 13 9 1 9 14 1 9 1 0 9 1 0 9 2
2 9 13
9 0 9 10 0 9 15 3 13 2
10 9 13 9 9 9 1 3 0 9 2
23 1 9 13 14 0 9 2 7 7 0 9 1 9 7 3 9 1 3 0 9 9 11 2
23 12 9 9 15 3 3 0 9 13 2 1 0 13 0 9 2 3 0 7 9 7 9 2
9 13 4 13 9 9 1 9 9 2
16 9 15 1 10 9 13 3 0 9 7 9 2 13 11 9 2
15 1 11 1 9 3 13 2 7 3 15 13 9 15 9 2
10 9 3 13 0 9 1 9 0 9 2
19 13 0 9 1 9 9 2 9 2 0 9 7 13 0 9 1 10 9 2
19 13 9 2 16 1 9 9 11 4 1 0 9 13 3 3 7 1 9 2
23 9 13 2 16 3 12 9 9 11 13 1 0 9 2 15 13 3 3 16 1 12 9 2
33 9 2 11 2 0 2 9 2 2 0 12 2 12 12 11 2 9 2 2 2 12 2 12 12 2 9 2 2 12 2 12 12 2
9 9 2 13 13 9 9 1 9 9
3 9 13 9
8 9 9 13 0 9 7 9 9
8 9 1 11 11 13 3 0 2
16 7 12 9 1 12 9 1 0 0 9 13 9 1 9 13 2
10 15 1 9 15 13 2 7 13 15 2
16 13 13 9 0 0 9 1 9 2 16 4 13 9 1 9 2
2 11 11
6 9 3 13 0 9 2
13 1 9 13 1 0 9 1 11 3 12 9 9 2
6 9 3 13 1 9 2
10 0 9 7 0 9 3 13 1 9 2
16 13 9 2 0 9 9 2 0 9 1 9 1 11 7 11 2
9 13 15 7 3 1 11 15 13 2
8 16 13 0 0 9 9 9 2
4 13 0 9 2
7 1 11 15 13 14 3 2
7 13 13 3 1 9 9 2
5 2 14 2 1 9
18 1 0 9 11 11 13 9 11 11 9 1 0 9 1 9 9 12 2
19 1 0 9 2 16 3 13 9 2 16 1 9 15 13 2 15 13 0 2
10 9 14 13 10 9 1 9 1 9 2
4 15 13 15 2
15 7 2 9 2 13 15 0 13 1 9 7 13 3 3 2
4 13 15 3 2
9 15 3 13 1 9 2 0 9 2
7 9 15 7 13 0 9 2
5 13 2 13 0 2
15 16 9 13 2 16 1 9 11 13 0 0 9 15 9 2
15 14 15 0 2 9 2 12 9 2 9 2 9 7 9 2
17 13 0 0 9 2 1 0 9 9 2 15 13 0 1 0 9 2
18 9 10 9 1 15 13 2 7 3 13 14 1 9 15 9 7 9 2
53 13 3 9 1 9 2 0 9 9 2 9 9 1 9 9 9 2 9 1 0 9 2 0 9 2 15 4 15 13 1 9 9 2 9 1 9 0 9 1 9 2 0 9 1 9 9 7 0 9 1 9 9 2
2 13 9
11 9 9 7 13 2 0 9 1 15 9 2
12 1 0 9 1 9 9 15 13 1 11 13 2
15 9 11 15 13 7 15 3 13 2 13 11 11 2 9 2
10 16 9 3 9 11 13 13 0 9 2
6 1 9 15 3 13 2
11 7 13 2 15 13 0 7 13 15 13 2
18 7 3 13 2 3 13 0 9 13 7 10 13 13 1 9 9 9 2
9 9 0 9 13 0 3 1 9 2
7 1 9 1 11 13 9 2
6 9 1 9 9 13 2
6 15 13 1 0 9 2
14 1 9 9 4 13 3 9 9 9 2 13 11 11 2
11 1 0 9 11 2 11 13 12 5 9 2
2 0 9
9 0 9 13 13 3 1 0 9 2
11 1 9 15 9 13 0 13 0 0 9 2
25 9 1 0 0 9 0 11 1 11 2 15 0 9 3 12 9 13 2 13 9 1 0 9 9 2
16 11 13 1 2 7 13 2 16 4 11 1 15 13 14 9 2
13 3 2 16 15 15 13 9 1 11 2 15 13 2
5 3 13 0 9 2
8 13 3 13 1 10 0 9 2
7 15 3 13 0 9 9 2
21 13 9 12 0 9 9 7 0 0 9 2 15 13 3 0 9 0 9 1 9 2
3 15 13 13
6 0 13 1 9 9 2
11 1 9 9 12 15 9 13 3 1 9 2
6 9 9 15 7 13 2
18 3 13 9 1 11 3 12 0 9 2 12 5 9 13 9 3 15 2
6 3 15 13 9 9 2
9 0 9 13 1 12 9 12 9 2
9 1 11 1 9 9 13 3 15 2
5 15 3 3 13 2
18 1 9 11 11 15 1 9 12 9 13 1 9 3 1 12 9 9 2
22 1 9 12 9 9 1 9 12 2 1 12 5 9 2 15 0 13 1 12 9 9 2
7 3 15 3 13 0 9 2
12 1 0 9 1 12 9 9 13 3 12 9 2
8 1 15 13 14 12 1 9 2
30 9 2 11 2 11 11 2 0 12 2 12 12 11 2 9 2 2 2 12 2 12 12 2 9 2 2 12 2 12 12
14 9 2 13 4 13 13 0 9 2 15 13 0 9 2
4 9 1 9 2
6 9 13 1 12 9 2
20 0 9 11 2 0 9 0 9 7 0 0 9 15 0 2 15 12 9 13 2
1 11
3 1 0 9
19 11 2 0 2 9 2 11 2 10 0 9 13 1 9 11 1 3 0 2
9 9 13 3 13 9 1 9 9 2
12 0 9 9 7 0 9 15 13 1 12 9 2
13 9 13 1 12 9 7 9 9 3 13 0 9 2
22 9 2 11 2 0 2 9 2 11 2 12 12 11 2 9 2 9 2 2 12 2 12
1 11
3 1 0 9
10 9 1 11 2 10 9 13 0 9 2
24 1 0 9 13 3 3 12 0 9 2 3 10 9 1 9 2 7 7 9 0 7 1 9 2
17 1 9 1 12 1 12 9 15 3 1 12 9 13 1 12 9 2
19 9 9 13 0 9 9 7 3 0 9 2 1 15 13 1 9 3 9 2
12 15 13 7 0 9 1 9 7 9 0 9 2
25 9 2 1 11 2 12 12 11 2 9 2 2 2 12 2 12 2 9 2 2 12 2 12 12 12
1 11
3 1 0 9
21 9 3 2 0 11 2 10 9 1 9 7 9 15 13 1 0 9 11 7 9 2
21 9 0 9 1 3 0 9 11 15 15 13 13 1 10 9 1 9 9 9 9 2
12 1 11 13 0 9 3 1 0 9 1 11 2
13 9 9 13 0 9 7 9 9 14 1 9 9 2
39 9 2 3 2 0 11 2 9 2 11 12 2 12 12 11 12 2 9 2 2 2 12 2 12 12 12 2 12 12 12 2 9 2 2 12 2 12 12 12
1 11
3 1 0 9
24 9 11 2 9 2 9 2 9 2 9 2 0 2 2 15 13 1 0 9 0 9 0 9 2
19 9 13 1 0 0 9 7 13 0 9 0 9 2 15 13 14 0 9 2
17 1 0 9 15 9 13 3 3 2 1 15 13 9 0 9 9 2
38 9 2 11 2 9 2 9 2 0 2 2 0 12 2 12 12 11 2 9 2 2 2 12 2 12 12 12 12 2 9 2 2 12 2 12 12 12 12
1 11
3 1 0 9
22 9 11 2 9 9 2 1 9 7 9 9 9 2 9 7 0 9 2 1 9 2 2
20 3 0 9 0 9 2 0 0 0 9 7 9 0 9 2 13 0 0 9 2
18 15 13 0 0 9 1 0 9 2 15 15 9 13 3 1 0 11 2
32 9 2 11 2 9 9 2 11 11 12 2 12 12 0 11 2 9 2 2 2 12 2 12 12 2 9 2 2 12 2 12 12
4 2 9 13 2
4 9 7 0 9
11 9 9 9 11 1 0 9 1 9 13 2
15 1 0 9 13 3 2 3 1 15 2 9 7 0 9 2
11 9 9 13 13 9 1 12 2 9 12 2
16 13 3 9 1 15 2 16 4 9 7 9 13 1 10 9 2
2 11 11
16 1 0 9 13 9 1 0 9 0 0 9 0 7 0 9 2
18 0 9 13 13 3 13 0 9 0 9 2 15 15 13 1 0 9 2
24 1 9 0 9 13 9 9 9 2 16 1 0 9 4 13 14 0 9 1 9 0 9 9 2
19 1 9 3 0 0 9 15 13 0 1 15 7 10 9 13 15 0 9 2
14 9 4 13 10 9 13 9 7 9 9 1 0 9 2
23 0 0 9 13 1 11 11 2 0 9 9 9 11 2 0 9 2 15 13 3 0 9 2
21 0 9 1 9 4 13 4 13 9 0 9 2 1 0 9 3 1 12 9 3 2
15 0 9 13 1 9 9 1 9 7 9 9 9 7 9 2
21 9 15 13 14 1 9 0 7 0 9 2 7 7 1 9 9 0 9 7 9 2
5 13 15 13 12 2
24 3 0 9 4 13 13 3 9 1 15 2 16 15 3 13 9 2 16 4 0 9 13 0 2
6 2 14 2 0 9 2
30 1 9 3 13 0 9 1 9 9 1 0 9 2 7 13 12 2 16 1 0 7 0 2 15 15 9 13 1 9 2
19 3 13 13 1 9 2 15 13 9 9 2 0 9 2 0 7 0 9 2
4 13 15 9 2
23 16 9 15 13 2 15 4 13 13 1 0 0 7 0 9 2 3 15 9 9 3 13 2
10 7 4 15 13 9 9 7 0 9 2
19 10 9 7 13 0 2 16 0 9 15 13 10 9 1 0 9 7 9 2
12 13 4 1 15 7 1 9 9 12 2 12 2
35 16 10 9 13 1 10 9 0 2 3 13 0 13 1 9 2 3 15 1 9 13 2 16 4 3 13 1 9 9 1 9 9 1 9 2
25 3 15 13 12 9 0 9 2 2 9 9 7 9 9 2 9 7 9 9 2 2 0 9 9 2
21 1 0 9 13 0 9 1 9 0 9 1 11 7 11 7 10 9 1 10 9 2
15 0 9 15 1 9 3 13 7 3 15 4 13 9 9 2
22 7 3 13 13 2 14 15 10 0 7 0 9 13 7 13 1 9 2 1 0 9 2
15 13 7 13 1 9 9 3 2 1 0 9 1 12 9 2
9 1 0 9 9 13 1 0 9 2
47 7 13 0 2 15 15 13 15 0 3 13 1 9 2 16 4 13 1 9 12 0 9 2 1 15 13 15 0 9 9 2 1 9 15 2 15 13 1 0 9 3 0 1 9 1 9 2
13 3 1 12 9 13 13 2 9 13 10 9 9 2
7 15 13 3 13 16 9 2
23 0 9 15 1 9 9 7 9 13 2 7 15 4 13 13 2 16 15 13 9 1 9 2
26 7 13 0 15 1 0 0 9 1 9 13 2 16 13 1 9 2 7 1 9 9 2 3 1 9 2
6 0 2 15 2 13 2
2 11 11
3 9 1 9
10 9 9 1 2 10 9 2 13 13 9
17 13 0 15 13 9 1 0 9 2 3 3 2 16 13 3 13 2
6 14 3 15 15 13 2
7 7 1 15 13 0 9 2
18 1 10 9 9 13 0 3 13 2 16 13 1 9 2 15 3 13 2
14 9 13 7 0 7 0 9 0 2 7 0 9 9 2
26 3 9 10 9 1 2 10 9 2 4 15 13 13 1 0 9 7 15 15 13 0 9 1 0 9 2
18 1 10 9 13 0 9 9 12 7 12 0 9 2 0 9 1 9 2
1 9
23 9 1 9 15 13 0 9 2 0 1 9 2 16 0 1 9 0 9 9 13 7 13 2
15 2 15 13 3 1 9 0 0 9 2 9 2 9 2 2
9 0 9 13 9 13 1 0 9 2
12 16 3 13 2 13 9 3 13 0 9 0 2
23 1 9 10 0 9 13 13 12 0 9 0 1 15 2 16 0 9 1 0 13 7 3 2
31 12 2 16 0 9 13 2 13 9 9 0 1 10 9 2 0 1 0 2 3 0 2 9 2 16 10 9 13 7 13 2
21 16 15 0 2 15 9 13 2 13 13 9 10 9 2 13 10 9 13 3 0 2
10 3 10 0 9 0 13 9 0 9 2
38 12 2 1 0 9 2 16 0 13 13 1 9 0 9 2 13 3 9 0 3 2 7 2 0 13 13 0 9 2 16 4 0 13 2 16 9 13 2
14 9 15 7 13 2 16 0 13 3 2 16 9 13 2
23 9 0 9 13 3 9 9 0 2 1 10 9 7 9 13 2 16 0 9 13 7 3 2
3 13 1 9
14 16 15 0 9 1 0 13 2 13 1 10 9 9 2
19 1 9 7 13 0 9 9 1 9 2 7 0 13 3 13 9 0 9 2
15 13 3 0 9 1 0 2 16 1 10 9 13 3 9 2
12 0 9 13 15 2 16 0 1 0 9 13 2
6 15 13 9 0 9 2
16 0 13 1 0 9 0 9 7 13 9 9 9 1 10 9 2
41 9 9 0 2 0 1 0 9 2 13 9 9 0 2 7 1 10 9 7 9 13 2 16 3 0 0 9 13 7 16 10 9 4 13 3 7 1 9 0 9 2
9 13 1 9 0 2 3 15 13 2
37 16 13 13 7 3 9 0 9 2 15 13 1 15 2 13 2 16 13 0 9 13 2 16 4 9 13 2 7 15 3 13 9 1 9 10 9 2
24 1 0 9 2 13 2 14 0 13 9 0 9 2 13 1 0 9 13 0 2 16 9 13 2
16 10 9 13 0 13 1 10 9 2 1 15 15 1 0 13 2
29 16 0 13 0 9 1 10 9 0 13 2 13 3 9 10 9 13 2 1 9 1 15 2 16 0 9 3 13 2
20 10 9 0 13 9 9 2 16 9 9 1 15 13 9 9 9 1 0 9 2
2 11 11
27 13 0 9 11 2 0 2 0 12 9 2 12 12 11 12 2 11 2 9 2 2 2 12 2 12 12 12
4 9 1 9 2
5 13 9 1 9 2
12 15 13 1 9 9 9 1 2 10 9 2 2
5 9 2 9 7 15
3 9 1 9
11 13 0 9 7 9 10 9 13 1 9 2
22 13 2 16 4 15 13 0 9 7 13 13 1 15 2 16 13 1 9 1 0 9 2
6 11 2 11 2 2 11
36 1 0 9 13 9 9 9 12 2 12 9 2 2 1 9 0 0 9 7 0 9 1 9 1 0 7 9 0 0 9 7 1 9 1 9 2
17 1 10 0 9 13 13 0 0 9 2 1 15 13 13 9 13 2
28 1 0 9 7 13 2 16 9 0 1 9 13 9 1 0 9 1 9 2 16 9 1 9 13 3 12 9 2
2 9 9
14 16 15 10 0 0 9 13 2 13 4 15 9 0 2
27 3 2 1 9 12 9 7 12 9 2 13 2 16 7 15 13 0 7 13 15 15 3 2 3 4 13 2
6 7 4 13 9 13 2
4 13 15 0 2
9 1 3 3 15 3 13 13 9 2
6 11 2 11 2 2 11
21 16 9 0 9 13 3 9 1 9 0 9 7 0 0 9 1 9 7 0 9 2
11 13 7 13 1 0 9 1 0 0 9 2
10 10 9 7 13 13 12 1 12 9 2
24 16 4 10 0 9 13 1 12 9 2 13 1 9 9 13 1 9 2 16 0 0 9 13 2
2 0 9
11 10 9 13 13 1 0 9 1 9 12 2
20 3 4 15 13 2 16 1 0 9 13 1 0 9 13 1 0 9 0 9 2
12 1 9 9 9 13 3 12 9 12 9 0 2
4 13 15 0 2
13 3 15 13 13 2 16 3 0 9 10 9 13 2
6 11 2 11 2 2 11
12 0 9 9 13 13 0 1 0 9 0 9 2
31 1 0 9 13 1 9 1 0 9 0 0 9 9 0 9 2 16 10 9 13 1 10 9 7 1 9 0 1 0 9 2
11 1 0 9 13 1 9 9 0 9 9 2
28 1 15 13 2 16 9 2 15 13 0 1 0 9 3 2 13 13 10 0 9 2 7 9 9 13 3 0 2
34 1 0 9 15 2 15 13 13 1 10 9 0 9 0 9 2 13 15 1 0 9 13 2 16 4 15 10 9 13 7 13 0 9 2
14 3 13 13 0 9 2 15 13 4 13 7 1 9 2
34 1 15 13 2 16 15 13 13 1 9 7 13 2 16 4 0 9 4 13 13 15 9 10 0 9 2 3 10 0 9 13 9 0 2
2 9 9
23 13 9 0 9 7 1 9 13 1 15 2 16 12 1 15 15 3 13 7 13 15 9 2
19 16 13 12 3 13 2 4 13 7 15 4 7 13 2 16 0 9 13 2
27 3 4 15 13 2 16 0 9 1 15 13 9 9 2 15 15 13 1 9 15 2 16 13 13 9 9 2
3 13 3 2
6 11 2 11 2 2 11
35 0 9 13 9 1 9 9 1 0 9 2 16 0 9 1 9 3 7 3 0 0 9 2 1 9 10 0 0 9 1 9 0 0 9 2
23 1 15 13 0 2 16 1 0 9 13 9 13 1 15 2 15 13 15 0 9 2 9 2
2 9 9
26 13 15 1 9 1 0 9 7 9 9 13 7 9 9 1 15 2 16 13 1 0 9 0 1 9 2
18 13 4 15 2 16 10 9 4 13 13 2 7 13 13 0 0 9 2
7 11 2 11 2 2 0 11
37 1 9 1 0 0 9 9 3 7 3 0 0 9 13 9 2 9 7 0 9 0 1 0 9 0 9 7 1 9 0 9 2 15 13 0 9 2
15 15 13 2 16 9 9 4 13 1 10 9 13 1 15 2
6 9 2 9 2 11 11
25 9 13 2 0 7 0 9 2 0 12 2 11 12 2 9 2 5 9 2 2 12 2 12 12 2
5 9 2 10 0 9
1 11
24 0 9 1 11 7 11 13 3 1 12 9 2 9 2 16 0 9 13 1 12 9 2 9 2
15 1 9 12 13 0 9 1 12 5 7 9 1 12 5 2
22 0 9 0 9 13 9 7 0 9 2 12 5 2 2 9 2 0 9 7 0 9 2
26 1 0 9 15 13 9 2 12 5 2 2 9 2 12 5 2 7 9 7 0 9 2 12 5 2 2
16 3 15 13 9 0 9 2 16 13 9 9 7 13 9 9 2
17 1 11 13 9 0 9 7 0 9 1 12 0 2 3 0 9 2
47 9 1 9 2 15 13 1 11 14 12 9 9 2 4 13 3 1 9 2 9 2 3 9 7 11 2 2 9 2 11 0 2 2 7 7 0 9 2 11 2 7 0 9 2 11 2 2
20 1 11 13 0 9 0 9 2 15 4 13 1 0 9 2 11 2 11 2 2
1 9
14 1 0 9 1 12 9 13 9 11 3 0 0 9 2
9 1 10 9 7 13 1 11 13 2
18 1 0 0 9 13 13 9 0 9 9 2 15 13 1 9 0 9 2
20 1 9 15 13 13 0 0 9 2 15 13 1 9 0 9 2 3 0 9 2
12 11 13 0 9 1 9 0 9 1 0 9 2
14 13 13 3 0 9 2 15 15 13 9 1 9 13 2
4 9 0 9 2
13 3 13 0 9 1 11 1 12 0 9 0 9 2
25 13 15 9 2 13 9 0 7 0 9 2 14 1 9 1 0 9 2 15 13 7 13 0 9 2
22 13 1 15 7 0 9 1 9 0 0 9 2 15 0 9 9 0 9 13 7 13 2
25 0 9 13 1 9 3 9 12 9 9 2 1 15 13 0 9 1 9 0 9 1 9 7 9 2
43 9 2 0 9 1 9 11 2 0 15 2 12 2 11 12 2 1 9 0 12 2 2 9 2 2 2 12 2 12 12 12 12 2 9 2 2 12 2 12 12 12 12 2
1 9
9 2 0 9 2 0 9 1 9 2
3 9 1 9
19 9 9 2 1 15 13 3 1 9 1 12 9 2 3 3 13 10 9 2
31 13 15 1 15 1 3 12 9 10 9 2 15 15 13 10 9 2 10 9 9 13 10 9 1 0 9 9 9 0 9 2
17 16 3 13 0 0 9 2 13 13 15 2 15 13 0 9 3 2
16 10 9 7 13 0 9 2 15 9 1 10 9 7 9 13 2
19 4 2 14 13 0 9 10 9 2 13 15 3 1 9 1 3 0 9 2
20 12 1 15 13 3 9 11 11 2 0 9 7 0 9 2 15 13 0 9 2
4 9 9 9 13
10 1 0 9 1 0 9 13 9 9 0
21 1 0 9 0 9 13 0 0 9 10 9 9 2 15 15 3 13 0 0 9 2
30 1 15 2 1 10 9 13 0 0 9 1 0 9 2 10 9 1 10 9 13 2 4 13 1 10 0 9 11 9 2
2 11 11
13 2 1 9 0 0 0 9 13 3 16 9 9 2
15 3 13 9 0 9 10 9 1 0 9 9 1 0 9 2
30 13 15 15 13 1 0 9 2 16 2 7 15 1 9 2 13 9 9 9 2 3 13 0 9 2 0 16 0 9 2
16 3 0 15 13 1 9 7 1 9 2 3 15 13 3 9 2
12 13 1 0 9 9 2 7 0 15 3 13 2
7 2 13 15 3 10 9 2
13 16 13 2 3 1 9 1 9 12 4 3 13 2
10 3 15 3 13 2 9 9 13 0 2
19 13 15 7 9 14 3 0 9 2 7 3 0 9 1 9 1 0 9 2
27 13 2 16 0 9 2 15 9 1 9 12 9 9 1 9 9 13 3 9 7 0 9 2 15 3 13 2
18 0 13 2 16 10 9 13 1 9 2 7 1 0 16 0 9 9 2
12 2 15 13 2 16 3 0 9 13 9 9 2
4 7 3 9 2
23 0 9 13 0 9 7 0 9 2 15 13 13 9 1 0 12 9 9 7 13 15 9 2
20 13 3 0 9 0 9 2 7 3 10 9 2 3 1 15 9 1 15 0 2
13 7 3 10 9 1 9 13 0 1 9 0 9 2
17 2 13 15 13 3 2 16 1 0 9 13 9 13 9 0 9 2
5 13 15 3 0 2
41 13 3 9 0 0 9 1 9 2 7 3 15 9 2 15 13 0 1 9 9 9 7 15 13 9 9 7 9 9 1 10 9 2 10 9 13 3 13 7 13 2
19 3 3 2 16 13 0 9 7 9 9 2 3 13 9 3 1 0 9 2
4 2 15 13 2
43 13 2 16 4 13 13 9 1 9 12 1 12 9 12 9 2 7 15 4 13 13 1 15 2 16 4 3 1 0 0 9 13 3 13 0 0 7 0 9 1 0 9 2
22 7 9 10 9 13 9 3 0 9 9 9 2 3 13 9 2 3 9 10 0 9 2
23 3 7 13 2 16 13 1 0 9 7 0 9 2 3 13 1 10 9 9 1 0 9 2
25 2 3 13 9 10 9 1 0 9 2 10 0 9 2 10 9 9 0 9 7 10 9 1 9 2
3 3 3 2
22 13 3 1 15 2 16 9 13 12 0 9 7 15 2 15 1 15 13 2 3 13 2
33 1 0 9 9 15 13 12 9 9 0 9 2 15 13 9 1 0 9 9 9 9 2 15 4 13 3 1 9 13 1 12 9 2
22 16 13 1 9 0 14 0 9 2 3 13 0 2 16 3 0 0 9 9 4 13 2
17 2 13 15 2 16 10 9 0 9 13 0 9 1 9 9 9 2
16 14 2 7 7 4 1 0 0 9 13 7 0 7 0 9 2
14 10 9 13 9 0 7 0 9 2 0 13 0 9 2
32 9 3 13 2 16 9 10 0 9 13 0 9 9 2 15 13 3 0 2 9 15 13 1 9 3 14 12 9 7 12 9 2
23 2 0 9 2 0 0 0 9 2 15 4 0 3 13 2 13 13 9 0 9 3 0 2
27 13 1 15 2 16 9 9 13 2 1 9 1 9 2 1 0 9 0 9 2 16 13 1 9 9 9 2
13 7 1 9 9 15 13 9 0 9 1 12 9 2
17 13 15 0 16 1 9 9 1 9 2 3 3 13 1 9 9 2
23 1 9 11 7 11 4 9 9 3 13 3 2 16 4 3 13 0 9 16 9 0 9 2
27 16 15 13 1 9 2 3 15 13 16 9 2 16 9 13 0 9 2 16 1 9 15 10 9 3 13 2
14 1 10 0 9 15 7 13 13 7 1 9 7 3 2
10 13 7 3 0 9 2 0 0 9 2
28 13 15 2 16 0 9 13 1 0 9 3 2 7 14 0 13 3 0 2 16 4 15 13 0 9 3 13 2
14 2 13 4 15 13 3 1 12 9 2 0 0 9 2
19 13 9 2 16 1 15 0 9 1 9 7 14 12 9 13 12 9 9 2
17 13 4 3 0 9 1 0 9 0 9 2 14 1 12 9 9 2
29 9 13 2 16 16 4 13 15 9 2 15 4 13 3 1 9 2 3 3 13 0 9 13 7 13 15 13 9 2
33 9 1 12 9 2 1 15 13 9 9 2 13 0 2 7 1 1 0 9 13 0 2 16 3 3 3 15 1 15 13 0 9 2
7 2 3 15 10 9 13 2
24 1 9 13 3 3 0 9 3 0 9 2 1 15 15 0 9 1 9 13 2 15 1 0 2
11 1 0 2 9 3 14 13 3 1 9 2
40 13 15 7 1 10 9 3 9 2 16 1 12 9 9 2 7 0 9 2 15 3 13 14 12 9 2 13 13 2 3 13 2 9 1 3 0 9 0 9 2
20 13 1 15 13 3 0 9 3 0 9 2 3 13 1 0 9 13 0 9 2
10 2 15 4 15 13 3 1 0 9 2
18 1 10 9 1 9 0 13 1 15 9 0 12 2 13 1 9 9 2
8 0 9 13 2 3 15 13 2
28 9 15 15 13 3 0 2 16 1 9 0 2 7 15 3 2 16 9 9 13 3 3 3 0 2 16 3 2
26 1 0 9 3 13 9 1 9 12 9 9 9 1 0 9 2 13 1 15 2 16 3 13 0 9 2
25 7 1 9 15 13 7 15 13 4 15 13 13 12 2 0 0 9 7 13 15 3 16 9 0 2
46 15 13 2 16 3 13 9 15 2 7 0 9 7 9 2 7 13 13 1 10 0 9 2 15 15 14 3 13 1 9 1 10 9 0 9 7 15 13 7 0 0 9 1 0 9 2
2 9 2
17 9 0 0 9 1 9 13 0 3 2 16 13 0 9 10 0 9
3 0 9 9
9 7 1 10 9 13 13 0 9 9
18 1 10 9 15 4 1 9 12 2 9 0 9 13 0 9 0 9 2
18 1 0 9 9 2 15 13 4 13 9 1 9 2 13 12 0 9 2
25 1 0 9 12 9 0 1 12 2 9 0 9 13 12 5 1 9 2 10 9 9 13 12 9 2
33 1 12 5 13 1 9 1 0 9 0 9 2 1 15 15 13 0 9 9 2 3 2 0 9 11 2 11 11 2 11 11 2 2
79 1 0 9 3 1 9 0 2 0 2 0 2 0 9 2 3 2 0 9 11 2 9 9 2 9 11 2 11 2 13 13 9 0 9 1 9 0 2 0 2 0 2 11 11 2 9 0 11 2 9 11 2 11 11 2 7 9 0 2 3 1 0 9 7 9 2 11 11 2 11 11 2 9 11 1 2 11 2 2
36 1 9 2 15 7 1 0 9 9 1 0 9 3 13 3 16 12 0 0 9 0 9 2 15 1 9 12 13 3 15 9 0 1 9 9 2
3 13 0 9
5 9 13 0 9 2
17 3 15 1 0 9 13 0 9 0 9 2 15 13 3 3 13 2
15 15 0 9 13 9 0 0 9 7 0 9 1 0 9 2
26 0 0 9 13 9 3 1 9 0 2 0 7 0 9 2 15 14 3 13 13 10 3 0 0 9 2
15 7 1 10 9 13 7 13 15 3 0 16 9 0 9 2
24 1 0 2 0 7 3 0 9 7 1 9 2 15 13 1 9 0 9 0 2 13 9 0 2
23 10 9 15 13 13 0 9 1 0 0 9 7 3 15 13 1 0 0 9 7 9 9 2
27 10 9 13 14 9 1 10 9 2 7 3 7 3 0 9 2 15 15 13 3 15 13 1 0 0 9 2
19 13 7 3 7 10 9 2 15 15 9 0 9 10 9 13 0 9 13 2
22 10 9 13 0 9 9 2 13 3 0 2 13 13 1 0 9 2 3 0 9 9 2
22 10 9 2 1 0 9 1 9 2 15 13 13 9 2 3 13 7 3 15 13 9 2
3 9 0 9
38 1 9 9 0 9 1 9 12 1 0 9 13 10 0 9 12 9 2 15 13 12 5 0 0 9 9 15 9 1 0 9 0 9 2 12 9 2 2
21 9 1 9 13 2 16 0 9 9 9 9 13 0 7 0 0 9 4 13 9 2
35 16 15 9 9 15 9 13 1 12 2 9 12 1 12 5 1 12 9 2 9 0 9 13 3 3 2 1 12 5 7 13 9 12 9 2
14 1 10 9 9 1 9 3 2 1 0 9 2 13 2
22 1 12 2 12 0 9 9 0 9 13 12 9 2 15 13 7 14 12 5 0 9 2
20 13 15 2 1 10 0 9 13 1 0 9 0 9 0 9 2 13 7 0 2
23 13 3 3 3 13 0 9 2 9 7 9 10 9 2 0 9 10 9 2 10 0 9 2
21 1 9 1 12 2 9 13 0 15 13 1 9 10 9 7 1 9 3 0 9 2
10 1 9 13 3 13 0 9 0 9 2
22 9 13 0 2 7 13 2 14 3 2 13 13 7 1 9 9 0 9 0 0 9 2
5 11 9 2 11 0
34 9 2 0 0 9 2 0 2 9 2 2 11 12 2 12 12 11 12 2 9 2 2 2 12 2 12 12 2 9 2 12 12 12 2
8 13 2 13 2 2 13 1 9
10 3 13 0 9 11 9 13 9 11 11
20 1 9 9 1 0 9 11 1 9 0 9 12 5 9 11 3 3 13 9 2
8 3 12 3 13 0 12 9 2
24 11 15 3 13 9 13 7 1 15 2 3 13 0 1 9 9 2 15 13 0 9 1 11 2
18 2 3 0 2 13 12 9 2 12 9 7 13 10 2 0 9 2 2
2 11 11
11 9 9 2 3 13 1 11 11 0 15 2
33 13 2 7 16 4 15 13 13 2 16 9 9 10 9 13 0 0 9 0 9 1 9 7 9 1 9 0 9 1 10 0 9 2
15 3 0 9 15 3 13 7 3 15 1 15 0 9 13 2
14 3 15 13 2 16 0 9 9 0 0 9 3 13 2
11 13 15 3 1 13 3 0 9 1 9 2
50 7 11 11 13 0 12 2 0 9 2 15 13 1 0 9 9 12 9 9 9 2 15 1 0 9 13 1 0 12 0 0 0 9 1 0 9 12 9 1 12 0 9 2 1 15 12 0 0 9 2
7 1 15 13 9 10 9 2
7 13 3 1 12 9 9 2
23 13 15 3 7 3 15 13 0 9 2 7 9 3 0 7 3 0 9 13 3 0 9 2
6 3 13 3 0 9 2
49 0 9 2 12 9 9 2 13 1 9 9 1 0 9 2 0 0 9 7 0 9 1 9 7 9 2 9 9 0 12 0 9 9 9 7 9 0 9 3 0 0 0 9 16 0 9 11 11 2
16 3 3 15 13 3 9 0 0 9 1 0 9 0 0 9 2
25 3 13 3 13 15 2 16 10 0 9 15 1 10 9 13 16 0 9 3 1 12 7 12 9 2
30 15 15 13 0 9 1 0 9 2 0 0 9 7 0 9 1 9 7 9 2 3 15 15 4 13 3 3 1 9 2
13 13 15 3 1 12 9 9 2 15 7 3 13 2
28 13 15 2 16 0 9 4 3 13 10 9 1 9 2 10 9 13 0 3 1 9 0 0 9 2 0 9 2
14 1 10 9 15 2 1 9 9 2 3 13 11 11 2
26 9 0 9 4 15 1 0 9 13 1 0 0 9 2 1 15 13 9 9 0 9 1 12 9 9 2
31 9 13 13 3 2 12 9 9 13 13 1 0 9 0 9 2 12 9 13 0 0 0 9 7 12 9 0 0 0 9 2
25 1 9 9 11 1 9 12 13 1 10 9 9 9 1 0 0 9 1 9 12 13 1 12 9 2
13 15 15 7 13 2 3 13 2 12 2 9 12 2
9 13 2 15 15 13 13 9 15 2
24 15 12 9 13 3 13 7 13 9 1 0 9 2 7 15 15 13 13 7 13 1 0 9 2
5 13 14 1 15 2
23 13 15 2 16 9 10 0 0 9 2 15 13 9 9 11 2 13 1 10 9 3 0 2
19 10 9 4 3 13 2 7 16 13 9 2 16 10 9 3 13 9 9 2
12 3 0 9 13 13 9 1 15 9 3 9 2
19 1 1 15 2 16 10 9 13 1 0 9 2 13 15 0 7 0 9 2
30 1 0 0 9 4 7 13 4 3 13 10 9 7 9 1 9 2 1 15 4 15 13 1 0 9 2 15 15 13 2
14 13 3 9 2 16 13 1 9 0 9 0 0 9 2
6 15 13 3 0 9 2
29 13 2 14 15 14 3 1 2 9 2 2 16 13 9 7 13 9 2 13 13 1 0 9 1 9 0 9 9 2
46 1 10 9 13 3 13 2 16 11 11 15 13 13 0 0 9 2 15 13 0 13 9 9 9 1 9 10 9 2 3 1 9 2 16 9 15 13 0 0 9 1 9 1 10 9 2
19 15 13 1 0 9 2 15 4 13 4 13 3 0 12 9 9 11 11 2
6 0 9 2 9 2 9
3 9 0 9
9 9 1 12 9 13 9 14 9 9
25 3 3 16 9 13 9 9 9 2 3 13 1 0 13 2 3 13 13 0 9 1 9 0 9 2
21 9 13 0 9 1 9 0 9 7 13 2 16 3 14 15 0 9 0 9 13 2
15 10 0 9 13 3 9 13 9 9 9 1 9 0 9 2
16 0 9 13 3 9 9 2 7 0 9 4 14 13 3 0 2
20 9 3 13 13 0 9 7 13 15 13 2 16 13 0 9 1 15 1 9 2
9 13 15 16 1 0 9 0 9 2
16 3 13 1 9 9 2 0 13 3 9 9 0 1 9 9 2
9 13 7 14 1 0 9 0 9 2
9 0 13 7 0 9 1 10 9 2
13 13 0 13 2 15 1 10 9 13 7 15 14 2
32 10 9 13 0 9 2 0 3 2 7 7 15 13 3 13 1 0 9 7 7 1 15 13 3 0 0 9 1 10 0 9 2
6 3 9 13 0 9 2
4 13 9 9 2
3 9 0 9
4 0 9 1 9
8 0 0 9 9 11 1 0 9
19 1 3 12 9 9 0 9 1 12 9 0 9 13 3 0 15 2 2 2
26 14 1 12 0 2 15 0 2 15 3 13 9 0 2 0 0 9 2 7 15 13 0 9 12 9 2
38 1 9 15 13 2 16 7 16 4 3 3 13 11 2 16 9 13 0 2 3 4 15 3 1 9 0 9 13 3 13 10 9 1 9 1 0 11 2
2 11 11
34 1 9 9 1 0 9 7 9 15 7 13 2 16 9 3 0 0 9 1 11 7 11 4 13 3 13 3 9 0 9 7 15 0 2
29 0 9 4 3 13 1 9 3 0 12 9 2 7 3 7 3 2 2 7 1 9 13 0 9 9 9 0 9 2
2 13 9
26 9 1 10 9 13 0 9 9 11 2 15 15 13 13 3 1 9 0 0 0 9 1 9 0 9 2
40 16 13 1 10 9 0 9 2 16 9 9 2 2 1 0 9 7 13 16 0 0 9 9 2 15 15 13 3 0 0 9 13 0 9 1 0 9 1 11 2
18 1 9 9 13 10 9 13 3 1 9 12 9 7 3 1 0 9 2
30 10 9 7 15 13 1 9 2 16 0 9 7 9 4 13 3 0 9 1 9 9 1 9 10 0 9 1 0 9 2
4 9 1 0 9
26 3 10 9 13 3 0 2 16 0 9 0 9 1 0 9 15 13 3 9 9 1 9 7 0 9 2
29 10 9 15 13 13 1 9 0 9 1 9 2 9 7 9 2 11 11 2 9 1 0 9 9 0 9 1 11 2
17 1 0 9 2 15 4 13 3 13 1 9 1 12 2 9 13 2
51 12 2 1 12 2 9 13 1 0 9 9 1 9 11 11 7 11 11 2 1 10 9 0 9 2 0 9 2 13 1 9 9 0 9 7 9 9 9 11 1 11 11 9 1 9 9 7 1 9 11 2
14 12 2 1 12 2 9 4 11 11 9 0 9 13 2
27 10 9 13 1 0 0 9 2 11 2 0 0 7 0 9 2 2 15 4 13 1 9 0 9 0 9 2
27 12 2 3 0 9 1 9 9 9 13 7 10 9 13 1 11 13 7 3 2 7 1 9 0 9 11 2
20 12 2 9 9 11 13 9 15 9 0 1 9 9 0 0 9 13 11 11 2
13 13 15 1 9 9 12 1 9 12 2 9 12 2
9 1 10 9 13 13 7 0 9 2
16 12 2 0 0 9 4 13 1 0 0 9 0 9 7 9 2
10 10 9 15 13 1 9 9 0 9 2
35 12 2 9 9 10 9 13 1 9 9 9 12 0 9 12 2 12 9 2 2 0 1 9 12 9 12 1 9 9 9 12 2 12 9 2
28 12 2 1 15 9 13 1 12 2 9 9 2 16 4 1 9 0 9 13 9 13 9 7 0 9 9 11 2
16 12 2 0 9 16 1 0 9 4 11 13 7 1 9 0 2
3 9 1 9
10 16 13 0 9 3 13 9 0 9 2
9 6 1 15 2 13 15 15 13 2
6 7 9 13 3 0 2
3 9 13 9
5 0 9 0 9 2
6 0 0 11 15 13 13
19 9 1 0 0 9 13 0 9 11 11 11 1 0 9 0 0 9 9 2
17 1 10 9 2 15 13 1 9 15 0 9 2 13 9 1 9 2
18 0 9 1 9 3 3 9 9 13 9 0 9 7 13 3 1 9 2
8 9 11 15 9 13 1 9 2
2 11 11
15 0 9 13 2 16 15 0 0 9 9 13 1 0 9 2
19 0 9 13 3 2 12 1 15 13 9 2 13 15 11 11 2 9 9 2
15 1 9 15 13 7 1 15 2 13 15 7 10 0 9 2
18 13 4 15 13 0 0 9 1 9 7 3 13 9 2 3 9 13 2
4 9 0 7 0
15 0 9 4 13 0 9 2 7 9 3 1 9 9 13 2
15 2 0 9 13 13 3 3 1 9 9 1 9 9 2 2
9 0 0 9 13 9 13 0 9 2
21 3 13 10 9 2 14 9 13 9 0 9 2 1 0 9 7 13 15 1 9 2
17 16 13 7 13 9 9 13 2 13 1 9 9 0 1 0 9 2
12 15 9 13 7 1 0 9 0 9 7 9 2
9 0 9 7 13 1 0 0 9 2
14 14 3 15 1 0 9 13 11 11 11 1 0 9 2
11 15 13 0 9 2 11 2 11 2 9 2
11 1 0 9 2 9 3 0 7 0 9 2
18 9 9 7 9 15 1 9 9 3 13 9 9 11 11 1 9 3 2
13 9 15 13 7 9 2 9 0 0 9 1 15 2
19 9 0 9 2 0 7 0 2 13 10 9 2 13 15 1 15 9 9 2
10 13 15 3 13 0 9 1 0 9 2
20 1 9 9 15 0 2 0 2 11 13 1 0 9 7 9 0 9 7 9 2
12 13 13 1 9 0 9 1 0 7 0 9 2
53 1 9 13 3 1 9 9 2 0 3 14 1 11 2 7 1 10 0 9 0 2 7 0 9 2 1 0 9 2 0 9 2 0 9 1 9 7 9 2 7 3 7 1 9 0 0 9 2 7 3 0 9 2
15 13 15 2 16 0 9 0 0 9 13 0 16 10 9 2
2 0 9
20 1 0 9 13 9 13 0 0 9 3 7 3 2 3 3 15 9 13 13 2
26 13 15 1 15 11 2 9 0 2 0 2 0 2 0 9 2 7 3 7 9 1 0 7 0 11 2
13 9 15 13 3 15 0 9 7 13 7 9 0 2
8 13 1 9 9 1 0 9 2
17 1 15 3 1 0 9 13 1 9 0 9 2 3 1 12 9 2
21 9 9 13 1 15 10 9 1 9 7 3 15 15 13 7 9 13 9 0 9 2
25 1 15 2 16 9 9 11 11 11 13 0 2 13 7 10 0 0 9 1 9 1 0 0 9 2
38 9 2 11 11 11 2 0 9 12 2 12 12 11 12 2 9 2 2 2 12 2 12 12 12 2 12 12 12 2 9 2 2 12 2 12 12 12 2
16 9 11 11 11 4 1 9 1 9 0 9 13 9 9 12 2
5 2 9 1 9 2
4 13 3 13 2
5 13 9 7 13 2
10 10 3 0 9 13 13 13 9 9 2
24 1 9 2 16 15 13 1 9 2 13 9 1 0 7 0 9 7 10 9 13 1 0 9 2
9 0 9 13 0 3 1 10 9 2
2 0 9
21 13 4 15 2 16 13 1 9 0 0 9 13 7 1 9 9 1 9 1 9 2
4 11 11 2 11
38 13 2 14 13 1 9 9 1 0 0 9 2 13 15 15 9 0 7 0 9 1 9 2 7 15 14 1 9 9 0 1 10 9 1 9 0 9 2
8 9 1 0 0 9 13 13 2
20 13 7 13 1 15 2 16 9 0 1 9 13 3 0 16 9 1 0 9 2
7 9 4 13 13 13 15 2
15 7 13 13 15 1 9 9 7 9 1 9 0 0 9 2
6 9 2 9 2 11 11
24 9 2 0 7 3 0 9 2 0 12 2 11 12 2 9 2 5 9 2 2 12 2 12 12
3 1 9 9
17 13 9 7 13 4 13 2 16 0 9 13 7 0 9 1 9 2
4 11 11 2 9
42 9 9 1 10 9 1 9 13 13 9 9 12 2 12 9 2 1 9 0 9 2 9 9 12 2 12 9 2 2 12 2 12 9 2 7 12 2 12 9 2 2 2
15 9 0 9 13 1 9 13 0 1 9 0 9 0 9 2
4 15 15 13 2
17 9 13 9 0 1 9 2 9 2 1 9 12 9 7 12 9 2
25 13 15 15 1 9 0 1 9 2 9 2 9 2 9 2 9 2 9 1 9 2 9 7 3 2
17 9 13 9 2 9 7 0 9 2 15 4 13 9 3 12 9 2
3 0 9 2
37 1 9 4 13 9 1 9 12 2 15 13 0 9 11 12 7 3 16 9 13 9 9 9 9 2 9 9 13 13 9 9 12 1 9 12 2 2
16 1 9 13 4 1 9 13 7 0 9 2 9 7 3 2 2
18 0 9 15 13 14 1 9 2 7 9 15 13 1 9 9 2 9 2
2 9 2
19 1 9 9 13 0 9 2 15 13 7 1 0 9 0 9 0 0 9 2
6 1 9 13 0 13 2
14 9 2 1 12 9 2 3 0 7 0 1 12 9 2
6 9 9 1 0 9 2
14 16 13 1 9 0 7 9 2 13 15 7 10 9 2
7 9 9 3 1 0 9 2
14 1 0 9 13 0 13 0 0 9 2 0 9 2 2
15 9 1 9 1 9 2 3 7 10 9 1 9 7 9 2
30 9 0 9 1 9 9 2 15 13 9 10 9 2 9 9 7 9 9 2 13 1 9 2 9 0 9 7 3 2 2
16 0 9 9 2 1 0 9 15 9 2 1 9 10 0 9 2
27 2 13 2 14 10 9 1 9 2 13 9 9 13 7 1 9 9 13 2 16 9 13 0 0 9 2 2
15 0 9 1 9 0 11 2 11 2 16 13 1 9 2 2
6 0 9 1 15 13 2
19 16 7 9 13 9 9 7 9 1 0 9 2 13 0 9 13 7 13 2
16 9 0 9 13 1 9 12 9 2 16 9 13 15 9 2 2
9 9 1 9 15 13 9 0 9 2
14 1 0 9 15 13 1 9 1 12 9 1 12 9 2
11 9 13 13 9 9 1 9 7 9 9 2
28 9 13 2 9 9 2 1 10 9 15 13 2 3 4 13 2 1 3 13 7 3 15 7 1 15 4 13 2
15 9 13 0 2 0 9 7 9 13 13 9 0 1 15 2
27 9 1 9 2 0 9 2 3 15 9 13 13 2 16 9 4 13 2 13 13 15 13 9 9 1 9 2
8 11 11 2 0 0 9 2 11
41 9 2 0 0 9 2 0 9 12 2 1 9 12 2 12 12 11 12 2 11 2 9 2 2 2 12 2 12 12 2 9 2 2 12 2 12 12 2 12 12 2
5 1 9 15 9 13
6 15 13 2 13 1 12
13 13 4 12 2 15 4 13 0 9 1 9 9 2
15 1 9 4 15 13 13 0 0 9 1 9 3 12 9 2
12 9 9 15 13 9 10 12 9 13 0 9 2
7 13 1 0 7 0 9 2
5 13 4 12 9 2
23 7 15 13 1 0 9 16 9 9 2 7 2 0 7 0 2 7 13 0 1 0 9 2
11 13 4 9 0 9 1 9 1 0 9 2
16 10 9 1 9 2 0 9 2 1 10 9 13 9 9 0 2
10 7 0 9 13 9 1 12 9 3 2
8 15 4 13 13 9 0 9 2
25 1 9 0 9 13 10 9 2 15 13 3 0 2 13 7 13 1 12 9 2 0 7 0 9 2
25 16 9 13 1 0 9 2 13 0 13 0 7 0 9 2 7 3 13 0 13 9 9 7 9 2
11 3 13 12 9 2 7 3 13 3 0 2
8 1 0 9 4 15 13 13 2
11 1 12 9 0 9 13 9 3 1 9 2
22 9 2 0 9 10 9 2 15 7 13 1 9 2 7 9 13 9 1 12 9 12 2
11 1 0 9 9 13 7 9 1 9 9 2
15 1 12 9 15 13 3 2 16 3 14 14 13 0 9 2
13 7 14 3 16 9 9 2 7 3 1 0 9 2
11 9 3 13 9 2 16 13 1 0 9 2
2 9 2
23 2 3 13 0 3 13 2 16 0 9 10 9 12 9 15 1 9 9 13 1 0 9 2
17 2 9 13 0 9 2 7 13 0 15 13 1 0 9 7 9 2
6 11 2 11 2 0 11
22 9 0 1 10 9 2 0 1 0 9 9 2 4 3 13 7 3 13 9 12 9 2
10 4 3 13 1 0 9 1 12 9 2
19 13 15 1 15 2 10 9 4 15 1 9 13 7 10 1 15 13 9 2
3 9 9 12
17 0 9 0 4 13 0 9 9 1 0 9 1 9 12 9 9 2
25 9 9 4 13 12 9 9 2 12 9 9 4 13 1 9 9 7 0 9 4 13 1 9 9 2
18 10 9 7 9 15 1 0 9 13 2 7 3 10 9 10 9 13 2
33 1 9 9 9 11 4 3 1 9 9 13 1 0 9 0 12 9 9 2 7 2 15 13 1 0 9 0 2 2 13 10 9 2
13 0 9 13 10 0 0 9 9 1 9 12 9 2
23 12 9 10 0 0 9 1 0 9 0 9 13 9 2 0 0 9 13 1 9 7 9 2
4 9 2 0 9
3 9 1 9
24 9 13 9 10 9 2 7 9 15 13 9 15 2 16 10 9 4 0 0 9 13 1 9 2
7 0 9 1 15 3 13 2
21 16 0 9 13 1 9 0 0 0 9 9 15 2 15 13 9 2 13 0 9 2
7 11 11 2 2 9 9 2
2 10 9
3 9 1 9
8 2 9 9 2 12 2 12 2
33 1 9 2 0 1 9 9 1 0 9 2 15 15 13 9 1 9 9 1 9 2 13 2 16 15 13 1 9 1 0 0 9 2
33 7 4 1 9 9 13 9 1 9 3 2 16 4 9 9 13 13 0 9 1 9 1 12 1 12 9 7 1 12 1 12 9 2
12 9 1 12 1 12 9 13 13 1 9 9 2
31 0 9 13 13 3 1 0 9 0 9 2 7 1 10 9 13 0 9 1 11 1 9 1 0 9 13 1 9 9 9 2
27 1 9 9 15 13 13 9 13 9 9 1 9 1 9 0 9 2 7 16 9 3 0 9 3 3 13 2
33 3 4 9 3 0 9 13 1 15 2 16 1 1 9 1 0 9 4 0 9 1 12 1 12 9 1 12 2 12 2 12 13 2
20 3 4 3 13 7 9 1 9 9 2 15 4 13 9 7 9 0 9 0 2
19 13 3 9 1 9 1 12 1 12 9 7 0 9 1 12 1 12 9 2
11 11 11 2 9 9 2 11 0 2 9 2
4 1 9 1 9
8 2 9 9 2 12 2 12 2
11 13 3 14 13 1 9 1 0 9 9 2
16 13 15 13 7 1 10 9 2 16 0 9 3 13 1 9 2
20 0 9 13 0 0 9 1 0 9 2 15 4 3 1 15 13 1 0 11 2
22 1 0 9 13 1 0 9 0 9 2 9 4 13 7 3 13 2 16 15 15 13 2
8 15 13 0 9 1 0 9 2
19 1 0 9 13 0 9 2 3 7 13 15 2 15 4 1 0 9 13 2
8 3 4 13 15 13 9 9 2
21 1 10 9 13 13 9 2 16 0 0 9 13 9 3 3 9 2 15 9 13 2
24 13 9 2 16 9 0 9 7 9 9 13 13 10 9 2 15 9 13 7 15 13 13 9 2
26 7 15 13 15 9 2 7 9 0 9 7 9 2 13 4 1 15 2 13 0 9 1 0 9 13 2
12 13 1 15 1 9 0 0 9 1 10 9 2
4 11 11 2 11
4 15 13 0 9
8 2 9 9 2 12 2 12 2
18 1 9 10 9 4 1 9 0 9 13 9 2 15 13 13 10 9 2
24 13 2 0 2 9 3 1 2 0 2 9 2 16 13 10 9 3 12 1 9 10 0 9 2
19 0 2 15 9 13 13 2 13 13 9 9 3 12 0 9 1 10 9 2
24 1 9 10 12 9 13 9 1 9 1 0 9 2 15 3 13 2 3 7 9 13 0 9 2
32 15 4 7 13 13 1 10 9 2 13 12 2 9 2 2 16 10 9 13 1 9 12 2 15 13 3 1 12 9 12 9 2
14 7 4 9 10 9 13 3 13 2 9 1 0 2 2
6 11 7 11 0 2 11
5 13 1 15 1 9
8 2 9 9 2 12 2 12 2
21 13 3 0 2 10 9 1 9 13 9 2 3 1 0 0 9 2 0 15 9 2
8 0 13 7 2 16 13 0 2
24 10 0 9 7 13 9 1 10 9 2 16 0 9 1 0 9 13 1 12 7 12 9 9 2
28 1 9 7 9 13 9 3 0 2 16 15 15 13 13 14 15 2 1 15 13 9 10 9 1 10 9 0 2
31 9 1 9 13 9 1 0 1 0 9 2 9 1 9 2 16 13 9 2 0 9 2 9 2 9 2 9 2 9 3 2
21 13 15 2 16 0 0 9 1 10 9 3 13 1 0 9 2 7 3 13 9 2
17 0 0 9 3 13 1 9 1 9 13 2 16 15 1 15 13 2
14 3 13 9 13 15 1 9 1 0 9 9 0 9 2
4 11 11 2 11
1 12
34 13 4 15 2 15 14 13 2 0 2 9 1 9 2 9 7 9 2 15 13 1 0 9 12 2 0 9 2 10 0 9 0 9 2
23 1 0 9 4 10 9 1 0 9 13 3 7 13 4 15 12 9 1 0 9 0 9 2
2 11 2
13 13 4 15 2 13 1 9 7 0 9 13 0 2
9 13 4 7 13 2 0 9 2 2
24 3 4 13 9 1 12 9 0 9 2 16 13 3 13 12 9 1 3 0 9 1 9 9 2
6 11 11 2 11 2 11
6 9 0 9 1 0 9
8 2 9 9 2 12 2 12 2
10 3 10 9 13 0 0 9 1 11 2
42 7 1 0 9 3 1 9 13 14 9 9 2 16 9 15 0 13 3 1 9 2 3 13 10 9 1 9 1 0 9 2 16 15 1 3 0 9 13 13 9 3 2
11 9 13 9 9 7 1 0 9 7 9 2
22 1 1 15 2 16 9 3 13 4 1 9 13 9 9 7 0 9 2 13 3 0 2
34 9 9 3 13 7 10 9 2 15 15 13 9 9 2 3 9 7 0 9 15 3 13 9 1 9 2 15 15 1 9 9 3 13 2
12 16 15 9 9 15 13 2 13 15 9 13 2
20 9 13 15 2 15 13 2 16 9 10 0 9 4 13 13 9 0 0 9 2
4 11 11 2 11
3 12 0 9
13 9 9 4 15 13 13 3 2 16 1 0 9 2
47 1 0 9 0 9 2 3 2 1 1 0 9 0 9 2 0 9 16 7 0 9 0 0 9 2 1 0 2 0 7 0 9 2 2 9 9 1 9 12 2 12 3 13 1 9 9 2
26 0 9 7 9 15 7 13 9 9 9 1 12 5 9 9 12 1 12 2 12 5 1 9 0 9 2
1 2
22 9 0 9 0 9 1 9 13 3 3 12 9 2 9 2 7 2 3 12 5 9 2
42 7 16 3 7 0 9 13 0 13 1 9 9 9 7 9 9 9 2 13 2 16 9 3 13 0 1 9 12 2 12 9 2 9 3 2 12 2 12 5 9 2 2
16 15 4 13 3 13 0 9 11 2 0 1 9 0 9 9 2
11 9 1 9 2 1 9 9 7 0 2 2
2 9 2
8 3 0 9 0 9 3 3 2
11 13 15 0 9 2 16 13 9 1 0 9
2 0 2
9 9 9 2 13 13 2 9 13 2
6 9 13 1 9 3 3
5 13 9 7 10 9
11 1 9 0 9 15 9 13 3 9 9 13
50 13 15 3 9 2 7 9 13 2 16 1 0 9 3 3 13 0 9 2 14 1 12 5 2 3 2 1 9 9 1 9 9 9 1 12 5 2 2 7 9 9 15 13 1 9 9 0 0 9 2
2 9 2
2 9 2
6 7 12 2 7 0 2
22 0 9 4 3 13 9 0 9 2 15 7 1 9 0 9 1 11 13 1 12 5 2
28 1 9 1 10 7 0 9 13 13 9 0 9 1 0 9 9 9 1 12 2 12 0 9 0 1 9 9 2
3 9 13 9
33 0 9 2 13 0 9 0 9 7 0 9 9 2 4 13 13 1 15 3 16 9 2 7 9 0 0 9 4 13 13 3 0 2
16 1 0 9 4 1 9 9 3 13 9 9 1 12 5 3 2
10 1 0 9 9 9 4 3 3 13 2
20 3 0 9 0 9 13 3 7 3 9 1 11 2 7 1 3 0 9 9 2
27 9 1 11 15 3 3 3 13 2 7 10 9 4 15 13 13 14 1 9 12 1 1 0 9 0 9 2
13 9 0 9 0 9 3 13 3 2 0 9 9 2
21 15 15 13 1 0 9 13 7 1 9 9 1 11 2 3 1 9 9 9 2 2
3 0 0 9
28 9 7 9 9 11 2 0 9 9 0 9 2 4 13 13 1 9 0 9 3 9 0 9 1 0 9 9 2
16 9 0 9 7 9 9 9 4 7 9 9 3 0 9 13 2
11 0 0 9 15 1 9 13 1 12 5 2
22 1 9 12 7 4 9 0 9 3 13 2 15 15 13 9 9 1 3 12 0 9 2
29 9 0 0 9 4 1 9 9 3 13 2 7 7 13 0 13 0 9 0 0 9 1 9 3 12 2 12 9 2
29 10 9 7 13 0 0 9 13 14 1 12 2 12 5 2 7 1 9 12 13 3 13 9 9 12 2 12 5 2
33 9 0 9 2 7 1 9 7 9 9 1 0 9 2 3 13 1 0 9 1 15 3 2 15 13 13 7 1 9 12 2 12 2
22 3 0 9 3 13 0 9 0 9 9 1 11 2 15 15 3 13 14 1 12 5 2
25 1 9 12 13 9 0 0 9 0 16 9 9 2 16 0 9 15 1 9 13 1 3 12 5 2
4 13 1 9 9
37 0 9 1 9 1 9 1 9 2 1 9 1 9 0 9 9 2 13 1 11 3 0 14 1 9 1 0 0 9 2 7 7 1 11 7 11 2
61 10 0 2 9 2 2 3 16 0 9 1 0 9 9 1 9 10 0 9 2 13 3 0 9 2 15 1 0 9 2 9 2 12 9 13 3 14 1 9 12 2 3 1 9 12 1 15 9 2 15 15 3 13 2 13 3 3 9 9 2 2
26 7 13 1 9 1 10 7 0 9 13 0 9 0 9 2 0 1 9 9 9 1 12 2 12 9 2
7 2 13 15 2 2 2 2
14 13 9 1 9 2 9 2 9 2 9 2 7 3 2
12 13 13 2 3 13 0 2 0 7 0 9 2
8 13 13 9 1 0 9 9 2
7 3 1 15 13 10 9 2
10 10 9 13 1 9 0 9 1 11 2
3 9 2 9
11 13 4 13 10 9 13 9 9 7 9 2
6 3 13 9 1 9 2
4 11 11 2 11
25 1 9 10 9 4 15 13 13 3 2 16 0 9 9 1 0 9 7 0 9 13 1 9 9 2
5 3 3 13 9 2
16 1 0 9 13 1 9 2 15 13 9 13 7 1 10 9 2
16 9 1 9 7 13 13 9 2 3 9 2 15 9 9 13 2
35 1 10 9 13 10 9 1 11 12 1 9 0 2 1 11 12 1 9 9 2 3 13 7 9 9 1 9 7 1 11 12 2 9 0 2
32 0 9 7 13 1 9 0 9 1 0 9 2 15 13 0 2 0 9 1 11 12 2 15 13 1 11 12 2 1 0 9 2
9 9 1 9 4 13 7 0 9 2
2 11 11
16 9 2 0 2 0 9 1 11 12 2 0 12 2 11 12 2
15 9 0 9 1 9 2 9 9 12 2 12 12 11 12 2
3 9 1 11
31 1 9 0 9 4 13 0 0 9 2 11 2 1 9 1 0 9 9 1 11 2 0 11 2 12 9 3 1 11 2 2
16 0 0 9 13 0 9 1 9 7 9 9 2 9 7 9 2
8 9 13 13 7 9 2 9 2
9 9 13 0 13 3 1 9 9 2
53 9 2 0 11 9 2 9 2 11 11 2 9 2 11 11 2 9 12 2 11 2 12 11 9 2 0 2 11 2 9 2 2 2 12 2 2 12 2 12 2 12 2 9 2 2 12 2 2 12 2 12 2 12
4 0 9 1 9
6 13 15 9 1 0 9
10 1 9 4 13 0 9 1 10 9 2
9 13 15 7 1 9 13 13 3 2
10 1 9 15 13 2 16 4 15 13 2
3 9 13 2
5 13 13 3 3 2
12 13 1 0 0 9 2 3 13 15 0 9 2
2 11 11
10 1 9 0 9 11 13 9 7 9 2
9 9 3 13 9 9 9 1 9 2
13 1 9 13 2 1 9 13 9 0 7 13 9 2
2 13 9
8 0 9 9 13 1 12 9 2
15 16 15 13 7 1 9 2 13 15 13 14 12 12 9 2
21 9 13 13 7 2 13 2 2 13 9 2 2 13 2 14 13 7 15 3 13 2
8 13 0 9 9 3 13 9 2
11 10 9 13 1 9 3 0 9 9 9 2
14 1 11 7 13 9 0 9 1 0 0 9 1 11 2
17 9 2 15 13 9 1 9 9 2 13 9 0 9 9 0 9 2
24 3 13 0 13 12 2 12 5 0 9 9 16 0 9 7 3 3 13 12 7 12 12 9 2
5 9 13 7 3 2
17 9 2 9 1 0 9 1 0 9 13 9 13 9 3 1 11 2
19 1 0 9 1 0 9 0 9 7 11 13 2 15 13 1 10 9 13 2
16 16 13 1 9 0 2 1 0 9 7 9 9 2 7 3 2
2 9 9
16 1 9 9 12 15 1 9 1 9 9 0 9 3 13 9 2
16 11 3 13 12 0 9 2 1 15 12 1 12 0 9 9 2
14 9 15 1 9 9 0 9 7 0 9 13 1 15 2
13 3 13 7 9 9 1 0 9 1 9 0 9 2
11 9 9 13 1 11 3 1 0 0 9 2
10 15 13 1 0 9 12 9 14 9 2
19 0 9 13 1 9 12 9 0 9 2 15 9 13 1 11 7 1 9 2
17 0 9 13 12 9 2 10 9 4 13 3 1 9 0 9 9 2
2 9 3
23 0 0 9 13 9 9 1 9 9 2 9 9 7 0 9 2 0 15 1 9 10 9 2
17 9 15 13 2 3 0 0 9 2 0 9 7 0 9 9 9 2
17 9 15 13 3 13 2 7 3 1 10 9 7 1 9 0 9 2
10 13 15 0 1 9 7 9 0 9 2
7 3 4 15 9 13 9 2
25 7 3 1 0 9 15 13 11 13 15 9 2 0 1 9 2 7 1 11 15 13 14 0 9 2
2 9 0
19 11 13 1 9 1 9 11 1 12 9 2 1 15 13 0 9 0 9 2
11 0 9 13 2 16 9 13 9 0 9 2
18 10 9 13 0 1 9 9 2 10 9 2 9 9 7 0 0 9 2
6 15 9 0 9 13 2
19 13 2 14 0 9 11 0 9 12 12 9 2 9 1 9 13 12 9 2
16 9 13 1 0 9 9 2 9 10 9 13 7 1 0 9 2
17 16 15 13 9 9 13 7 13 1 9 0 2 9 13 10 9 2
22 15 9 3 13 2 16 4 13 0 2 3 15 3 13 9 0 9 7 3 10 9 2
19 16 11 13 9 9 1 9 9 2 13 9 9 2 7 15 13 9 3 2
6 3 15 15 7 13 2
35 9 2 11 2 9 2 9 2 0 2 2 0 12 2 12 12 0 11 2 9 2 2 2 12 2 12 12 2 9 2 2 12 2 12 12
10 9 2 11 11 2 9 2 11 0 11
2 9 2
3 0 9 2
8 13 0 9 7 0 0 9 2
4 9 2 0 9
4 9 0 9 13
15 9 9 13 9 2 15 1 9 1 9 13 7 0 9 2
7 13 15 1 15 9 9 2
15 13 4 1 0 9 1 11 11 1 9 9 9 7 9 2
24 2 13 9 9 1 9 9 2 15 13 0 0 9 1 9 1 9 0 9 1 9 7 9 2
13 10 9 3 3 13 2 10 9 15 13 1 9 2
6 14 16 13 1 9 2
11 13 9 2 7 15 13 0 10 9 13 2
15 7 3 13 7 13 13 1 9 7 9 9 2 15 13 2
7 10 9 15 1 15 13 2
21 13 9 9 0 9 2 15 15 13 13 0 2 7 9 10 0 9 13 3 0 2
19 2 16 15 13 3 13 2 16 9 13 9 1 0 9 7 13 15 9 2
2 14 2
4 15 13 13 2
11 2 13 0 13 9 1 9 1 0 9 2
6 0 9 15 3 13 2
20 13 15 3 1 9 2 3 13 15 9 13 1 9 2 3 1 9 0 9 2
9 9 0 9 13 13 16 0 9 2
13 2 13 3 9 3 3 13 2 16 13 9 0 2
10 9 0 9 7 0 9 13 15 13 2
8 9 9 15 9 9 13 3 2
10 13 15 9 2 7 13 15 3 0 2
18 2 3 16 1 0 9 9 3 7 1 9 13 0 7 3 0 9 2
19 3 4 13 9 13 2 16 15 13 1 9 2 3 13 3 13 1 9 2
14 13 4 15 13 3 15 2 16 13 9 3 0 9 2
9 16 13 3 0 9 2 3 9 2
15 10 9 13 9 3 10 9 2 16 0 9 1 0 9 2
6 15 13 15 9 9 2
23 9 2 15 15 7 9 13 14 1 0 9 2 1 9 7 9 2 9 13 10 9 13 2
7 7 3 0 9 3 13 2
16 2 1 15 3 4 13 13 13 9 2 15 15 13 13 9 2
32 13 2 14 9 2 15 13 0 0 9 2 13 4 0 15 13 1 9 2 16 13 3 2 9 9 2 1 11 2 9 9 2
16 13 3 0 9 2 3 15 3 3 13 11 7 3 15 13 2
22 9 13 13 3 3 0 7 16 15 15 13 2 13 15 1 10 9 2 9 7 9 2
10 2 13 9 9 13 3 1 0 9 2
18 16 13 1 0 9 2 13 0 9 2 16 4 13 1 9 0 9 2
16 1 15 15 3 3 13 1 9 2 7 1 9 15 3 13 2
25 3 13 3 3 0 9 2 16 4 15 15 0 13 13 3 1 9 2 16 15 3 13 9 9 2
5 13 9 1 9 2
8 9 1 9 0 9 0 0 9
13 0 0 9 15 13 0 9 16 9 0 9 9 2
18 10 0 9 0 9 1 3 16 9 9 13 1 9 9 1 9 9 2
24 10 9 13 0 2 1 0 9 2 1 9 1 0 9 2 14 1 9 1 0 9 10 9 2
18 1 9 9 13 2 16 13 13 1 0 9 1 0 9 0 0 9 2
24 1 12 5 15 7 13 1 9 12 2 12 9 2 3 1 9 2 3 9 13 9 10 9 2
3 9 13 9
44 10 9 2 0 15 1 9 9 1 0 7 0 9 2 13 2 16 3 0 9 13 2 15 15 13 9 7 9 1 0 9 1 9 0 9 2 3 0 1 10 9 1 9 2
12 9 1 0 9 15 13 7 10 9 0 9 2
22 3 13 10 9 9 0 12 9 2 15 9 0 9 13 3 13 10 0 7 0 9 2
25 3 14 12 5 9 13 0 13 1 12 9 1 9 0 9 7 1 0 0 9 14 1 12 9 2
36 13 1 15 9 2 16 9 2 0 9 0 9 2 15 3 3 13 7 13 2 16 4 13 0 13 1 9 7 10 9 9 1 10 0 9 2
19 1 0 0 9 13 1 10 9 12 5 9 7 15 1 9 0 0 9 2
11 12 9 13 9 2 9 7 0 0 9 2
17 12 9 13 9 0 9 2 9 13 9 1 9 7 9 0 9 2
3 9 7 9
42 9 13 1 9 9 1 12 5 9 1 0 9 10 9 7 0 9 10 0 9 2 1 12 5 1 9 0 9 2 7 15 13 1 9 2 15 13 1 9 7 9 2
17 1 0 9 13 9 1 9 1 0 9 7 0 0 7 0 9 2
44 0 0 9 15 7 13 14 1 9 9 1 9 7 9 9 1 10 9 2 7 13 0 9 9 1 9 7 9 9 2 1 15 9 13 13 9 1 10 0 9 7 1 9 2
12 13 15 3 0 9 0 1 9 1 0 9 2
19 1 0 9 13 9 9 2 9 7 9 2 15 13 9 9 14 0 9 2
31 9 15 15 13 2 16 1 9 0 0 9 13 0 9 9 1 9 2 0 9 7 0 9 2 3 2 3 7 3 0 2
38 9 9 0 0 9 1 12 2 9 12 13 2 16 9 9 1 0 9 13 9 3 1 0 9 2 1 0 9 15 15 13 9 1 9 7 0 9 2
5 11 11 2 9 11
30 9 2 0 0 9 2 0 12 2 12 12 11 12 2 9 2 2 2 12 2 12 12 2 9 2 2 12 2 12 2
4 9 1 9 2
8 9 1 9 13 1 0 9 2
18 9 3 4 13 3 3 1 10 9 13 7 10 9 9 1 10 9 2
3 9 0 9
4 3 0 0 9
8 0 9 13 3 3 16 0 9
18 1 10 9 15 4 1 9 12 2 9 0 9 13 0 9 0 9 2
17 1 0 9 9 2 15 13 4 13 1 9 2 13 12 0 9 2
14 9 12 9 7 12 9 13 1 0 9 9 1 0 2
22 13 15 1 9 2 3 15 3 13 9 0 9 7 9 1 9 0 9 2 3 11 2
25 0 9 1 9 12 2 12 13 3 3 1 0 9 7 13 1 0 9 9 1 9 1 10 9 2
10 0 9 13 1 9 0 9 3 0 2
21 3 7 3 2 16 3 0 9 9 13 1 0 9 9 9 9 7 0 9 9 2
2 0 9
17 9 9 9 1 9 0 9 13 1 0 9 1 0 9 3 0 2
21 1 0 9 4 9 13 13 9 13 1 12 9 2 1 0 9 1 0 9 2 2
28 1 0 9 13 3 9 0 9 9 7 11 2 9 7 9 1 11 7 0 11 2 0 9 11 7 9 11 2
23 1 0 9 13 0 9 9 14 12 9 2 9 2 7 14 9 1 0 9 1 0 9 2
2 9 9
34 3 16 9 1 9 0 9 0 9 7 9 9 1 9 9 9 1 0 0 9 13 0 2 16 0 9 1 9 10 9 13 0 13 2
22 9 9 13 0 9 1 0 9 1 9 2 16 0 9 9 13 13 0 9 0 9 2
12 0 9 0 9 15 1 0 12 9 3 13 2
25 9 9 13 9 9 0 9 2 1 0 9 3 2 16 3 1 9 12 13 1 0 9 7 9 2
2 9 9
9 0 9 13 3 0 9 0 9 2
14 9 12 13 0 9 1 0 9 9 0 9 0 9 2
30 0 9 13 1 9 9 2 3 9 4 0 9 13 1 9 0 9 9 7 13 9 1 9 9 0 9 1 0 9 2
16 0 9 9 0 0 2 9 7 0 9 13 0 9 3 3 2
12 3 0 9 0 9 13 0 9 16 1 9 2
3 9 15 13
24 9 2 7 3 3 9 2 13 0 9 0 9 7 0 9 2 0 7 0 9 7 0 9 2
15 1 9 1 9 13 9 13 0 9 0 1 0 12 9 2
13 0 9 15 13 1 9 0 9 0 9 0 9 2
27 9 13 10 0 9 3 3 2 1 9 12 0 9 11 7 11 11 0 9 2 2 1 0 9 7 12 2
4 9 1 0 9
17 9 9 9 9 7 0 9 13 3 0 1 0 9 16 1 9 2
12 0 0 9 0 9 1 0 9 13 3 0 2
21 13 15 13 3 0 9 2 7 9 0 1 9 15 3 13 3 1 0 9 9 2
29 9 0 9 13 1 9 0 9 9 2 16 9 13 13 1 0 9 9 2 1 10 0 9 13 9 3 9 2 2
22 0 9 13 13 1 15 2 16 13 3 9 9 1 9 7 16 0 9 13 3 0 2
5 11 11 2 11 11
36 9 2 0 0 9 2 0 2 9 2 2 11 12 2 12 12 11 12 2 9 2 2 2 12 2 12 12 2 9 2 2 12 2 12 12 2
4 9 2 9 9
6 9 1 12 2 9 9
31 13 9 11 2 9 2 1 9 12 2 12 12 11 2 9 2 2 2 12 2 12 2 12 2 9 2 2 12 2 12 2
38 13 0 9 7 9 2 0 2 9 2 2 0 9 2 0 12 2 12 12 11 12 2 9 2 2 2 12 2 12 2 9 2 2 12 2 12 12 2
37 13 11 0 11 2 0 7 0 9 2 0 9 12 2 12 12 11 12 2 9 2 2 2 12 2 12 12 2 9 2 2 12 2 12 12 12 2
23 13 11 2 0 12 2 12 12 11 12 2 9 2 2 2 12 2 12 12 2 12 12 2
27 13 9 11 2 1 9 12 2 12 12 2 11 12 2 9 2 9 2 2 9 2 2 12 2 12 12 2
36 13 11 2 9 2 9 2 0 2 2 0 9 2 0 12 2 12 12 11 12 2 9 2 2 2 12 2 12 2 9 2 2 12 2 12 2
36 13 9 0 11 2 9 2 9 2 0 2 2 0 12 2 12 12 11 12 2 9 2 2 2 12 2 12 2 9 2 2 12 2 12 12 2
37 13 0 2 0 2 11 2 0 11 2 9 2 9 2 0 2 2 11 1 11 12 2 12 12 11 12 2 9 2 2 9 2 2 12 2 12 2
10 13 0 2 0 2 11 2 0 11 2
9 9 1 10 9 13 0 9 9 2
7 13 1 0 9 0 9 2
12 9 13 1 9 2 1 15 1 9 9 13 2
3 15 0 9
9 13 1 0 9 2 13 15 1 9
12 0 0 9 13 0 9 9 1 9 0 9 2
12 3 9 13 11 11 2 9 9 11 1 11 2
5 15 13 0 3 2
2 11 11
24 9 1 9 0 9 4 0 0 9 13 16 9 9 2 15 13 0 1 9 7 9 0 9 2
14 9 13 13 9 1 0 9 7 9 2 1 0 9 2
9 0 9 4 13 9 1 10 9 2
9 12 1 15 15 13 9 0 9 2
25 9 4 13 13 9 2 15 13 1 0 9 0 9 2 14 16 9 2 9 7 0 9 0 9 2
14 0 9 4 13 13 3 0 9 7 13 3 12 9 2
30 7 15 13 0 2 9 13 13 15 2 9 2 0 9 2 9 9 2 9 7 3 15 2 15 13 13 1 10 9 2
7 9 15 13 13 3 15 2
11 7 3 15 13 1 9 9 3 16 15 2
17 9 4 13 4 13 3 1 12 2 9 12 1 0 0 9 11 2
34 9 2 11 2 9 2 12 2 9 12 2 12 12 11 2 9 2 2 2 12 2 12 2 12 2 12 2 9 2 2 12 2 12 2
1 9
3 13 1 9
21 9 13 1 9 2 15 13 9 9 11 2 13 11 11 1 0 9 1 9 9 2
7 3 13 1 9 13 13 2
8 15 13 10 9 1 0 9 2
13 0 9 13 13 16 9 1 15 2 15 3 13 2
39 13 15 1 9 3 7 0 9 13 0 9 2 7 3 13 1 0 9 2 1 15 15 9 13 13 2 1 9 7 9 2 15 1 9 10 9 13 13 2
32 0 9 3 13 1 0 9 2 1 9 2 1 9 7 9 2 1 9 9 2 9 9 2 0 9 2 7 7 9 1 9 2
25 16 11 11 13 0 9 2 1 0 13 2 0 9 15 13 2 2 15 13 2 16 4 13 2 2
15 0 9 13 2 2 15 13 9 7 15 13 0 9 2 2
22 0 9 13 2 2 15 13 9 2 15 13 9 2 15 13 1 0 9 10 9 2 2
13 16 13 10 9 2 4 15 13 16 9 1 9 2
28 9 2 9 11 2 0 12 2 12 12 11 12 2 9 2 2 2 12 2 12 2 9 2 2 12 2 12 2
6 0 9 7 9 1 9
18 9 0 9 13 15 9 1 9 9 2 9 7 9 1 0 9 13 2
19 10 9 13 1 9 11 11 0 9 7 9 1 9 2 15 13 9 11 2
6 13 13 1 12 9 2
12 1 0 15 13 0 7 0 9 7 10 9 2
16 0 13 13 9 2 10 9 2 9 1 15 2 7 0 9 2
13 0 3 13 1 9 9 7 3 13 0 0 9 2
7 9 13 13 3 1 9 2
31 9 15 13 13 15 3 2 16 4 15 15 1 9 13 13 0 2 15 13 9 13 0 9 1 0 9 7 9 1 9 2
33 9 2 11 2 1 9 12 2 12 12 11 12 2 9 2 2 2 12 2 12 12 2 12 12 2 9 2 2 12 2 12 12 2
4 13 0 9 2
9 9 9 7 9 1 9 7 9 9
22 9 9 2 7 3 15 1 0 9 3 13 0 9 2 13 1 9 1 9 3 3 2
13 15 0 2 0 3 2 15 0 2 0 3 0 2
15 7 3 15 2 9 7 9 2 13 15 0 2 15 13 2
12 9 4 15 13 13 9 9 0 9 7 9 2
5 15 3 3 13 2
4 7 2 2 2
2 11 11
13 1 0 9 13 9 2 15 13 13 1 10 9 2
28 12 1 9 2 15 13 10 9 13 1 9 2 13 11 11 2 9 9 0 9 2 9 0 7 0 9 11 2
15 9 1 15 13 1 15 2 15 13 13 9 9 0 9 2
11 2 13 1 9 9 9 0 9 7 9 2
2 3 2
18 3 3 2 16 1 15 15 13 10 9 2 15 13 0 7 0 9 2
24 15 15 3 13 7 16 15 9 10 9 13 7 13 15 3 13 2 3 15 1 0 9 13 2
24 1 9 15 3 13 0 9 2 15 13 9 9 7 9 1 9 2 13 9 7 3 15 13 2
4 9 3 13 2
10 15 13 3 9 2 3 15 0 9 2
18 7 12 1 0 9 9 13 13 9 7 9 9 2 15 13 10 9 2
20 2 13 1 9 0 9 2 15 4 13 9 7 13 1 10 0 9 1 9 2
7 0 13 3 9 13 9 2
18 1 9 9 13 1 9 9 1 0 9 2 15 13 13 9 1 9 2
23 3 15 2 16 1 9 0 9 4 9 13 0 9 9 2 16 13 15 1 0 0 9 2
26 13 3 13 9 9 2 16 4 9 13 2 16 9 9 13 12 7 1 9 13 14 12 7 7 3 2
6 1 9 3 13 13 2
19 1 9 9 9 15 3 13 7 0 9 0 1 10 9 2 3 7 9 2
9 2 9 15 3 13 3 1 9 2
14 9 4 13 9 9 2 16 3 13 0 9 7 9 2
9 7 3 4 13 9 13 1 9 2
6 3 13 7 0 9 2
18 9 2 15 15 13 0 9 2 3 13 2 3 1 9 1 15 13 2
26 7 4 9 13 1 0 13 2 3 1 9 13 2 15 13 0 9 2 3 15 13 7 3 15 13 2
19 2 15 13 3 0 1 0 9 2 7 1 0 9 13 9 7 0 9 2
8 4 3 9 13 7 0 9 2
2 3 2
27 9 4 13 3 13 9 2 10 9 13 2 15 15 13 2 15 1 9 13 1 10 9 7 9 14 0 2
38 13 7 1 9 9 9 9 2 3 4 13 15 0 9 2 15 10 9 13 2 1 10 9 15 13 2 10 9 10 9 13 2 3 16 9 10 9 2
43 9 2 0 9 2 9 2 9 2 0 2 2 0 12 2 12 12 11 2 9 2 2 2 12 2 12 12 2 12 12 2 9 2 12 2 9 2 2 12 2 12 12 2
4 9 2 0 9
2 0 9
15 9 0 0 9 13 3 10 2 16 9 1 15 13 9 2
15 3 15 7 1 15 13 9 2 15 15 1 0 15 13 2
15 1 9 11 13 9 11 1 9 1 11 9 0 0 9 2
42 1 0 9 2 15 10 9 3 13 2 7 9 13 7 0 9 1 0 2 10 0 9 9 13 2 3 15 13 2 1 10 9 15 13 13 16 9 2 3 15 13 2
8 13 4 15 0 9 7 13 2
9 1 0 9 7 1 10 9 13 2
19 13 14 1 15 13 2 16 9 2 15 9 13 9 0 9 2 13 0 2
22 0 9 4 3 9 13 2 0 9 7 9 13 7 0 13 1 9 9 3 0 9 2
4 11 0 2 11
14 0 9 0 1 10 9 13 1 0 9 7 0 9 2
11 4 3 12 3 13 1 9 1 12 9 2
26 13 14 9 2 15 4 13 1 10 0 9 2 7 7 15 2 1 15 15 9 2 9 13 16 9 2
2 9 13
14 0 9 1 0 9 1 11 13 3 0 0 0 9 2
33 13 1 0 11 12 2 12 0 9 1 9 9 7 9 2 0 0 9 2 1 0 9 2 1 9 9 2 0 9 7 1 9 2
20 10 9 15 13 3 2 3 1 9 1 0 9 2 9 13 13 1 0 9 2
15 16 9 0 9 13 3 0 2 13 0 9 1 10 9 2
31 1 15 13 9 1 0 9 2 11 2 9 2 12 2 12 2 12 2 12 2 0 9 12 7 13 0 9 1 10 9 2
5 9 7 1 0 9
6 9 1 0 9 15 13
10 3 13 3 0 9 16 1 0 9 2
17 3 7 3 13 7 3 7 1 9 13 9 9 1 9 0 9 2
13 14 15 0 1 15 13 13 10 9 2 10 9 2
30 3 0 9 11 2 9 2 9 2 0 2 2 13 1 12 9 2 3 13 12 9 7 1 9 13 10 9 3 13 2
11 1 9 9 15 13 3 1 9 0 9 2
17 1 15 2 1 15 13 10 9 2 13 9 1 10 9 11 11 2
14 3 1 9 9 9 13 15 9 1 0 7 0 9 2
6 13 15 1 10 9 2
17 16 13 1 9 2 11 13 1 10 9 1 9 2 15 3 13 2
19 13 1 0 9 11 2 15 1 0 0 9 7 0 9 13 3 0 9 2
11 9 13 3 1 9 9 13 1 9 9 2
18 15 3 1 9 13 1 9 2 15 13 3 3 1 10 9 3 9 2
21 15 2 15 15 13 10 0 9 2 7 10 9 13 7 13 15 0 9 1 9 2
20 0 9 13 13 0 9 11 1 0 0 9 2 13 15 15 3 9 7 9 2
4 9 7 1 9
9 1 9 0 9 4 7 9 13 2
18 7 1 0 0 9 13 3 10 9 2 15 13 0 7 0 1 9 2
11 1 0 9 13 15 0 9 0 9 9 2
10 1 9 9 4 1 9 13 3 3 2
20 1 10 9 13 9 9 0 9 1 0 0 9 7 9 9 0 9 1 9 2
16 9 15 13 9 1 0 9 2 16 4 13 0 13 0 9 2
8 3 11 13 9 10 9 9 2
17 7 15 7 1 10 0 9 2 7 3 1 9 7 1 9 9 2
22 3 1 0 9 13 0 9 9 10 0 9 1 9 11 2 15 13 1 0 12 9 2
2 9 9
14 0 9 13 1 0 9 3 9 0 2 0 2 11 2
10 9 11 11 15 13 3 1 0 9 2
11 11 11 3 13 9 9 7 13 15 13 2
14 3 13 9 2 15 13 14 1 0 9 0 9 9 2
14 1 15 13 13 0 9 2 15 13 1 9 3 3 2
65 1 9 10 0 9 2 0 7 0 9 9 2 9 9 1 0 9 2 3 2 3 3 7 1 10 9 9 3 13 2 9 2 3 3 3 13 2 9 2 3 3 13 7 3 2 13 1 9 9 9 0 9 9 1 15 9 1 0 9 1 9 1 0 9 2
25 16 15 13 2 16 1 9 0 9 13 7 13 1 15 9 2 13 9 3 9 1 0 9 9 2
33 1 0 9 2 15 13 3 1 9 2 7 9 13 3 13 2 13 1 9 9 1 9 9 2 1 9 0 9 7 9 1 9 2
6 11 15 13 9 11 2
11 10 0 11 13 3 11 13 1 9 9 2
2 0 9
18 1 9 11 13 9 2 0 3 0 2 3 0 9 1 9 7 9 2
11 3 13 15 9 0 9 11 7 0 11 2
14 3 3 13 0 9 0 1 9 2 9 1 0 9 2
25 11 11 13 10 9 7 13 15 3 0 9 2 10 9 13 9 13 15 2 0 9 7 9 9 2
8 3 13 11 13 9 0 9 2
25 13 9 7 3 7 13 9 0 9 2 9 2 9 2 9 2 9 2 9 2 0 9 2 9 2
12 9 9 1 9 13 9 1 9 0 0 9 2
15 3 13 1 15 2 16 4 15 13 0 9 1 9 11 2
30 11 11 13 7 0 9 15 15 13 2 16 16 4 13 3 15 13 0 9 9 2 13 0 1 15 13 0 9 9 2
2 11 11
29 9 2 11 2 9 2 9 2 0 2 2 0 12 2 12 12 11 12 2 9 2 7 9 2 2 12 2 12 2
3 9 2 9
8 13 0 9 1 9 1 9 13
17 1 9 13 13 1 9 2 7 3 16 1 9 15 1 9 15 13
18 13 4 10 9 7 16 13 0 9 2 13 4 15 13 9 0 9 2
13 3 4 13 1 9 7 10 9 15 15 3 13 2
13 13 15 9 9 1 12 2 9 2 9 3 13 2
9 10 9 1 9 13 7 3 0 2
16 15 4 13 13 2 16 4 13 2 16 4 15 13 3 13 2
10 13 3 0 9 1 9 1 0 9 2
6 11 11 2 11 1 11
7 10 0 9 9 11 13 2
17 1 0 9 15 13 13 0 9 1 2 13 9 2 3 0 9 2
18 3 0 9 11 11 13 3 1 12 12 2 3 15 1 12 3 13 2
13 0 9 1 15 12 9 2 15 13 9 1 0 2
4 0 13 7 0
42 1 11 11 2 15 13 9 0 9 12 2 9 1 0 9 1 11 2 15 13 13 0 3 0 9 1 9 15 2 16 9 2 1 15 13 3 9 2 13 10 9 2
16 3 0 9 9 13 2 16 1 15 1 9 13 13 0 9 2
21 1 9 15 7 3 13 0 9 1 9 1 9 9 2 9 2 9 7 0 9 2
20 3 9 1 9 1 9 13 0 2 7 9 10 9 7 9 9 13 9 0 2
42 15 4 15 3 1 9 12 13 2 16 1 0 12 9 0 0 9 2 15 10 9 3 13 9 2 0 9 1 0 15 9 2 2 4 1 12 9 13 1 12 9 2
3 9 13 0
10 1 9 9 4 13 3 0 9 9 2
15 0 2 7 0 9 0 9 13 3 3 0 16 0 11 2
8 0 9 13 0 1 0 9 2
11 3 3 0 13 9 11 11 7 11 11 2
7 1 9 15 7 3 13 2
11 7 13 0 13 2 15 4 13 13 9 2
10 13 2 14 9 2 13 15 15 13 2
15 9 7 1 9 15 9 3 13 2 16 15 13 3 3 2
14 3 4 14 13 0 9 2 7 3 10 9 3 13 2
41 1 12 2 9 2 12 2 9 2 3 15 13 0 0 9 2 13 3 9 3 1 10 9 2 9 7 9 11 2 11 2 11 2 11 2 11 2 11 2 11 2
50 1 12 2 9 2 12 2 9 13 3 13 0 2 9 0 9 2 1 15 13 3 11 2 11 2 11 2 11 2 11 7 3 0 9 12 2 9 16 11 2 11 2 11 2 11 2 11 2 11 2
2 0 9
30 9 0 9 15 13 1 9 12 2 3 4 13 0 9 2 7 1 0 7 0 9 13 11 2 11 2 11 7 0 2
13 9 10 9 13 1 9 7 3 15 13 1 9 2
10 1 9 0 9 13 3 3 0 9 2
11 0 9 9 1 15 13 1 12 12 9 2
15 0 7 3 3 0 13 9 9 9 11 2 0 2 9 2
36 1 15 13 1 3 0 11 7 11 2 3 3 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 7 0 2
13 3 1 11 15 10 0 9 13 13 1 12 12 2
8 9 9 7 13 14 1 9 2
4 9 3 1 9
5 13 3 9 9 2
23 0 13 9 2 13 9 7 9 2 14 1 9 0 16 9 13 13 9 7 9 10 9 2
27 13 2 14 1 9 11 1 0 9 1 11 0 0 9 12 12 2 1 10 0 9 3 13 3 1 12 2
18 0 9 2 14 12 5 12 9 2 10 9 9 9 13 1 12 9 2
3 14 0 9
8 0 9 9 13 3 9 9 2
5 13 3 13 9 2
6 10 9 13 3 9 2
13 3 1 9 2 1 15 15 3 13 10 9 9 2
16 9 7 9 13 2 3 4 9 13 2 1 9 7 9 9 2
8 0 11 13 3 0 16 0 2
28 9 3 13 1 9 2 13 2 14 9 9 1 15 2 16 13 13 1 9 2 7 4 13 1 9 7 9 2
14 9 2 9 7 9 1 9 1 9 3 13 9 9 2
28 7 15 13 0 1 9 2 3 13 1 9 10 9 2 16 7 0 9 15 13 3 13 2 16 13 9 0 2
24 1 9 15 13 9 2 16 1 10 9 1 11 13 11 11 7 13 2 9 10 9 4 13 2
3 9 1 9
21 0 2 15 15 13 13 9 2 4 15 13 3 13 9 2 1 10 13 9 9 2
4 13 12 9 2
17 15 0 2 15 3 13 1 0 9 2 13 0 9 1 0 9 2
18 3 3 0 13 9 1 0 9 2 1 0 9 2 15 13 7 0 2
12 0 9 13 3 9 1 0 9 2 16 0 2
16 3 0 9 13 2 13 2 14 9 1 0 9 7 3 0 2
13 13 1 9 2 15 13 1 0 9 13 0 9 2
21 10 9 3 13 2 14 1 9 2 7 0 9 3 13 1 9 12 2 12 9 2
9 0 2 0 9 13 3 9 0 2
11 13 7 9 2 3 13 9 0 16 9 2
15 3 15 2 3 13 9 0 2 13 15 13 9 0 9 2
21 7 13 3 13 15 2 16 3 13 0 9 7 0 9 2 16 0 1 0 9 2
3 9 1 9
25 9 11 4 3 13 9 2 15 3 13 9 9 2 16 13 1 10 9 15 0 2 3 9 9 2
14 9 13 13 1 9 2 9 2 1 9 7 1 9 2
12 10 9 15 10 9 9 13 3 3 1 9 2
8 9 15 1 7 10 9 13 2
29 7 13 1 9 3 3 3 0 9 1 9 2 7 13 0 13 15 1 9 9 1 9 9 7 13 1 9 9 2
21 7 13 3 0 13 2 3 15 13 2 16 9 13 3 15 15 0 2 3 0 2
3 9 1 9
13 1 0 9 13 1 9 0 9 12 12 0 9 2
25 3 15 13 2 16 13 15 2 15 4 13 9 3 1 11 7 15 15 15 13 13 1 0 9 2
32 1 9 9 9 9 11 11 2 15 15 13 12 2 9 12 2 4 0 9 2 12 5 12 9 2 13 1 0 9 12 9 2
11 3 4 15 13 13 3 3 1 12 12 2
12 0 7 13 2 16 7 1 9 15 13 9 2
8 0 1 9 13 3 0 9 2
22 3 15 13 2 16 15 9 13 2 3 13 1 9 0 2 16 1 15 15 9 13 2
17 1 12 2 9 9 11 11 1 12 9 15 13 12 9 1 12 2
14 9 9 11 13 12 5 7 13 15 0 1 0 9 2
24 0 9 2 15 4 15 10 9 13 13 2 13 9 11 12 2 9 1 9 9 1 12 9 2
12 1 9 15 13 12 9 7 9 13 3 12 2
18 10 9 1 9 13 0 15 9 0 1 9 13 1 0 9 1 9 2
10 0 9 1 10 9 13 14 1 9 2
31 1 9 1 9 13 0 13 1 15 2 16 15 13 3 2 3 1 0 9 2 7 1 10 9 13 0 13 9 12 9 2
19 1 9 9 1 11 13 0 9 0 2 9 2 9 9 1 12 2 9 2
11 9 13 12 9 2 12 9 13 1 9 2
9 9 13 0 13 12 9 1 9 2
4 1 9 10 9
8 1 9 7 9 13 13 3 2
13 13 1 15 2 16 13 13 7 13 7 3 3 2
38 3 13 13 0 9 2 3 1 0 9 11 1 0 9 1 11 7 1 11 1 9 2 3 13 3 1 9 11 1 9 7 0 9 13 3 0 9 2
10 13 4 12 0 9 1 0 0 9 2
23 9 9 1 9 13 9 9 1 0 9 2 16 10 0 9 13 0 16 12 9 2 9 2
15 13 1 0 9 2 1 12 1 3 0 9 1 0 9 2
6 13 15 1 0 9 2
7 13 1 0 9 12 5 2
23 0 9 11 11 2 14 12 5 12 2 2 9 2 4 3 13 9 9 13 1 12 9 2
29 1 15 0 9 10 9 2 14 12 5 12 2 2 3 0 9 2 13 1 0 9 1 9 11 1 9 12 9 2
27 3 13 13 2 16 9 0 9 9 15 1 11 13 1 12 7 12 9 16 1 11 1 12 7 12 9 2
4 1 9 1 15
5 15 0 13 9 2
5 0 9 3 13 2
14 16 4 10 9 13 1 11 9 13 2 13 12 9 2
34 7 15 13 3 9 2 7 13 9 1 0 2 9 7 9 3 3 13 9 7 13 15 0 12 5 9 7 12 5 9 1 0 9 2
10 9 15 1 10 9 15 13 0 9 2
23 13 2 14 15 1 10 9 9 1 12 9 2 9 13 13 9 14 1 12 5 9 0 2
23 13 2 14 9 1 10 9 2 13 15 9 3 7 13 0 9 12 5 1 0 9 9 2
3 3 15 13
23 9 11 1 9 13 0 7 10 9 13 1 9 15 2 16 15 13 1 3 0 9 9 2
9 0 9 15 3 13 14 12 9 2
4 7 13 9 2
10 9 13 3 1 12 0 16 1 11 2
11 7 3 13 0 9 1 9 7 0 9 2
36 1 9 2 15 13 1 9 2 15 13 1 9 14 12 5 2 9 13 11 7 13 1 9 14 1 12 2 12 5 0 2 16 13 9 0 2
7 9 1 0 9 9 13 2
9 0 9 1 0 9 13 12 5 2
20 3 12 9 15 1 9 13 7 13 15 9 2 15 13 10 0 7 0 9 2
27 13 2 14 9 9 2 13 9 9 3 1 9 2 7 13 15 3 2 16 1 15 4 13 9 1 9 2
17 13 15 3 9 1 9 2 16 9 2 15 9 13 2 13 0 2
2 13 9
18 13 2 14 9 9 0 9 2 1 15 4 13 2 13 13 0 9 2
17 7 13 3 13 1 9 2 13 2 14 15 2 16 13 1 9 2
15 7 13 15 13 2 4 2 14 15 13 9 1 0 9 2
22 9 9 13 9 9 9 3 7 3 0 2 13 1 15 2 16 0 9 13 10 9 2
32 3 14 15 0 9 13 9 7 1 0 9 3 13 0 2 16 4 9 1 9 13 1 9 2 3 3 13 15 1 9 0 2
20 10 9 4 15 13 13 0 9 7 13 15 1 9 2 15 15 13 13 9 2
11 9 0 9 13 1 9 1 0 0 9 2
3 9 13 2
25 3 0 9 2 13 2 14 1 9 11 11 2 3 7 13 13 0 9 2 16 10 9 13 9 2
4 9 1 9 2
15 3 15 13 7 1 9 12 1 9 13 0 9 11 11 2
5 9 2 9 2 9
13 1 0 9 9 13 3 9 3 12 9 0 0 9
19 0 7 0 9 13 10 9 1 0 9 7 1 9 7 10 9 3 13 2
15 10 9 3 13 9 9 11 11 1 9 2 15 13 9 2
2 11 11
33 3 13 3 1 9 13 2 0 9 1 9 0 7 0 9 13 13 3 1 0 0 9 2 0 0 9 7 0 9 9 0 9 2
3 3 9 9
28 1 9 3 13 2 16 1 9 12 4 3 1 9 3 0 7 0 9 13 1 0 9 3 16 12 9 9 2
22 3 15 1 15 13 9 9 9 11 2 7 15 9 0 9 1 9 3 12 9 9 2
32 0 9 4 13 9 9 2 3 12 9 9 2 9 9 7 0 9 2 1 12 9 9 2 7 9 9 2 14 12 9 9 2
21 3 3 9 13 1 3 0 9 0 7 0 9 3 12 2 12 5 0 0 9 2
2 0 9
23 1 9 0 9 13 9 0 7 0 9 0 0 9 7 0 9 7 3 7 9 0 9 2
15 0 7 13 2 16 9 0 7 0 9 13 0 0 9 2
14 0 9 1 3 0 9 13 13 0 9 7 0 9 2
35 9 0 7 0 9 7 3 13 1 9 1 9 3 0 0 9 2 7 9 2 2 0 0 9 2 3 3 3 0 9 1 3 0 9 2
18 9 10 9 13 13 1 9 11 11 3 0 9 9 16 0 9 9 2
4 9 1 9 12
32 9 9 9 11 1 0 9 13 2 16 1 1 0 9 9 9 1 9 9 15 3 13 7 10 9 1 9 0 9 1 9 2
26 9 13 0 9 9 1 0 9 2 3 9 2 15 9 9 13 1 9 9 9 0 0 7 0 9 2
33 9 11 11 2 1 1 0 9 7 0 9 2 15 13 1 9 1 0 9 2 4 1 0 9 9 9 1 9 12 13 0 9 2
4 1 9 2 2
22 1 9 9 9 7 11 4 13 9 9 1 9 9 1 12 2 12 5 1 9 12 2
4 1 9 2 2
19 4 13 9 1 9 0 9 1 9 9 1 9 1 12 9 1 12 9 2
4 1 9 2 2
17 4 13 3 0 9 1 9 1 0 9 7 13 1 0 9 9 2
4 1 9 2 2
14 4 13 9 1 9 9 1 0 9 1 9 9 9 2
24 9 0 9 13 9 9 1 9 0 9 9 1 0 9 1 3 0 9 1 9 0 9 12 2
20 13 7 0 3 13 2 16 1 9 13 0 9 7 13 15 14 1 9 9 2
3 3 12 9
9 1 9 12 4 13 3 12 9 2
11 1 0 9 13 15 0 9 9 7 9 2
30 9 4 7 13 13 9 9 9 1 9 15 9 1 9 12 2 7 15 1 9 9 0 9 1 15 9 1 0 9 2
28 9 11 11 1 15 13 2 9 4 13 1 9 0 1 0 9 0 9 1 9 12 1 0 9 12 9 9 2
35 9 9 1 9 0 9 1 0 0 9 13 3 1 9 9 1 3 0 9 1 9 12 3 12 9 9 2 15 4 13 1 3 0 9 2
26 0 9 3 3 13 0 9 1 0 9 2 3 9 9 1 0 9 9 2 7 9 9 1 0 9 2
20 13 1 0 9 0 9 2 15 0 9 9 2 15 3 0 9 1 0 9 2
19 13 2 16 15 13 12 1 0 9 9 10 9 0 9 7 10 0 9 2
7 2 9 2 9 2 7 9
17 1 0 9 15 13 13 3 2 3 1 15 13 9 10 0 9 2
5 9 13 3 0 2
14 0 9 7 9 13 2 3 13 2 1 0 9 9 2
28 16 4 9 13 9 9 2 3 13 9 2 16 1 9 9 1 9 15 13 9 13 7 3 13 10 9 3 2
20 16 9 3 13 7 0 9 7 0 0 9 1 9 9 2 9 7 9 9 2
11 15 15 13 13 2 13 1 10 9 15 2
24 13 9 1 9 2 15 13 9 0 2 9 0 13 1 9 0 0 9 9 2 11 7 11 2
54 9 1 9 7 9 1 11 3 1 0 13 2 16 1 9 9 13 1 9 0 9 2 16 15 13 0 9 9 7 9 2 15 13 0 9 2 13 0 0 9 2 3 13 1 0 9 2 0 9 2 9 7 9 2
11 9 1 9 9 13 13 7 9 1 9 2
33 11 13 9 2 13 2 9 2 9 2 2 1 12 9 2 11 3 1 12 9 7 11 15 10 2 14 2 9 13 1 12 9 2
13 3 0 9 13 1 9 9 1 0 7 0 9 2
34 3 1 0 9 13 1 9 0 9 1 9 1 12 9 2 0 1 12 7 12 9 2 7 11 15 10 9 1 9 13 1 12 9 2
30 15 13 13 9 1 0 9 2 9 7 9 1 9 2 16 13 0 13 1 0 9 3 2 16 15 13 1 0 9 2
18 1 9 0 9 9 13 7 1 9 0 9 9 9 9 7 0 9 2
35 0 9 15 7 13 7 15 2 15 13 9 15 2 16 15 13 1 9 2 7 15 13 1 0 9 1 9 9 7 3 13 10 0 9 2
28 9 1 0 9 1 9 9 13 3 0 2 7 13 0 3 13 1 9 2 16 7 3 13 9 1 9 9 2
11 9 9 15 7 13 13 7 13 3 13 2
14 15 4 13 1 9 1 9 9 0 9 13 1 9 2
20 2 13 3 1 9 9 0 9 7 9 1 0 9 2 3 15 13 1 9 2
34 2 13 1 15 2 16 9 1 0 2 9 2 9 13 3 0 2 16 9 0 9 13 13 14 1 0 9 2 15 13 1 9 9 2
18 2 13 15 13 1 0 9 1 9 9 2 16 15 4 15 3 13 2
14 2 13 9 1 9 1 9 2 15 3 9 3 13 2
7 13 7 13 2 13 0 2
2 11 11
2 9 9
4 1 9 9 2
3 13 0 9
5 1 9 15 13 2
23 15 3 13 0 9 9 2 15 15 13 10 0 9 1 9 7 0 9 7 13 10 9 2
15 1 15 13 9 7 9 13 2 1 15 4 15 13 13 2
11 0 0 9 4 13 13 15 9 13 9 2
35 3 15 13 1 9 1 9 1 9 9 2 16 15 13 14 12 0 9 0 9 7 15 13 2 3 1 0 9 2 9 9 10 9 13 2
14 9 4 13 3 13 9 9 7 9 9 0 9 9 2
16 7 3 13 1 2 0 9 2 2 7 1 12 0 9 9 2
1 9
29 1 0 9 13 13 0 9 9 9 7 9 2 1 9 1 15 2 16 13 1 9 0 7 0 9 2 7 9 2
9 7 4 13 9 13 9 7 9 2
12 9 1 0 1 0 9 13 13 1 9 9 2
19 15 13 0 9 1 9 0 9 9 9 2 15 13 13 0 9 9 9 2
16 9 13 2 16 9 9 9 1 9 9 1 9 9 9 13 2
9 3 13 4 10 9 13 0 9 2
7 9 9 13 9 0 9 2
14 15 13 2 16 1 12 9 13 4 9 13 15 0 2
18 1 9 0 9 13 9 9 0 9 2 15 15 13 1 12 0 9 2
1 9
13 9 9 9 15 1 9 9 1 0 9 15 13 2
25 1 9 12 9 2 12 0 9 2 16 13 1 9 9 1 0 9 2 13 9 1 0 9 9 2
8 13 7 3 13 0 0 9 2
31 13 15 7 13 2 16 0 9 15 4 13 13 9 3 2 16 4 13 0 9 2 15 1 15 4 13 0 9 0 9 2
9 7 4 13 1 9 0 9 9 2
21 0 9 15 1 9 0 9 13 1 9 12 9 2 12 13 9 9 1 9 9 2
9 3 13 13 1 15 1 10 9 2
24 9 2 9 13 9 1 15 2 9 2 10 9 2 9 2 9 7 9 2 10 9 7 9 2
30 9 2 16 9 13 13 9 2 1 15 13 9 0 9 13 2 7 9 13 9 1 0 9 2 15 4 10 9 13 2
22 9 2 16 9 7 15 2 15 1 15 13 2 1 0 9 3 13 0 9 1 9 2
35 9 2 16 9 3 13 10 9 2 0 1 9 9 2 3 15 2 16 13 9 7 9 1 9 0 1 9 9 1 9 0 16 12 9 2
44 9 2 13 2 14 0 1 9 0 9 1 9 7 1 9 13 3 2 16 9 13 13 2 7 13 2 14 9 7 9 9 2 1 10 9 13 0 9 7 9 0 9 13 2
33 9 2 13 2 14 1 9 2 15 13 3 1 9 0 1 9 9 7 0 0 9 7 9 7 9 10 0 9 13 10 9 13 2
28 9 2 13 2 14 9 12 7 3 9 2 1 9 2 16 1 15 13 3 13 2 16 4 13 3 12 9 2
11 9 2 13 2 14 9 9 1 0 9 2
18 1 9 13 13 2 16 9 4 13 3 9 1 9 10 9 1 9 2
23 3 4 13 0 0 9 13 9 13 7 14 9 9 2 3 10 9 7 0 9 1 9 2
15 15 4 13 9 9 2 16 4 15 2 13 2 0 9 2
8 3 1 9 0 9 0 9 2
5 11 11 2 0 9
4 9 1 9 2
17 9 9 2 13 3 9 2 3 16 9 15 13 16 0 1 9 2
2 9 9
18 1 9 13 0 10 9 2 3 1 3 0 9 13 0 9 0 9 2
18 1 12 9 10 9 13 0 9 0 9 12 1 0 9 1 9 9 2
19 9 1 9 2 10 11 2 4 13 2 16 13 1 9 12 0 1 11 2
7 9 3 13 1 0 9 2
7 0 9 13 10 12 9 2
13 9 13 1 9 9 3 16 12 0 9 7 9 2
14 13 1 15 7 12 2 15 4 15 13 3 1 9 2
6 0 9 13 10 9 2
8 15 13 13 10 9 9 13 2
21 0 9 7 9 1 11 13 1 0 9 9 2 16 13 0 9 1 9 9 9 2
15 10 9 13 2 16 9 13 0 3 12 9 7 7 0 2
23 7 10 9 4 13 9 1 9 12 13 0 9 2 15 9 13 1 9 1 12 12 9 2
11 9 15 3 13 9 2 15 13 1 9 2
18 15 13 9 1 9 0 9 7 13 1 9 2 16 15 13 1 11 2
8 9 13 3 3 2 3 3 2
14 7 9 2 15 13 13 9 0 9 2 13 0 9 2
13 9 13 13 0 9 1 9 7 13 15 1 9 2
8 11 4 13 1 0 0 9 2
24 1 9 15 13 2 16 9 0 4 13 2 13 0 7 0 9 2 15 15 13 13 10 9 2
13 0 9 1 9 13 9 2 16 9 13 0 9 2
31 1 9 2 3 15 13 9 2 15 1 9 9 9 13 11 11 2 4 0 7 0 9 13 7 13 9 13 3 9 9 2
17 10 9 13 7 0 7 13 15 14 2 13 2 14 1 0 9 2
3 1 0 9
21 12 15 13 3 0 7 3 13 9 1 9 7 13 13 2 7 10 9 15 13 2
8 3 0 9 13 13 0 9 2
3 15 3 2
6 15 13 1 10 9 2
11 16 13 15 13 7 13 0 9 0 9 2
10 1 15 13 15 0 2 11 7 11 2
29 9 13 0 2 7 12 1 0 9 13 9 2 16 0 9 12 9 13 3 0 1 1 0 9 0 7 0 9 2
5 15 1 15 13 2
6 9 13 1 9 12 2
9 13 2 15 13 13 1 9 9 2
18 13 1 15 2 16 7 3 13 2 1 15 15 10 9 9 3 13 2
13 9 15 13 2 3 13 7 1 10 0 9 13 2
8 9 13 1 0 9 0 9 2
12 3 15 13 2 16 4 11 13 1 12 9 2
9 3 15 9 13 1 12 9 9 2
14 7 3 15 12 1 0 7 0 9 13 1 0 9 2
18 3 15 15 13 2 15 15 13 1 0 7 3 0 9 9 12 9 2
5 9 2 9 7 15
2 9 9
19 1 9 12 4 13 1 9 1 9 12 9 2 7 10 9 14 12 9 2
6 7 3 13 9 0 2
12 3 13 10 9 13 2 16 15 13 16 0 2
24 13 4 13 2 3 13 1 10 9 13 9 9 1 9 0 0 9 2 3 10 13 13 9 2
6 11 2 11 2 2 11
8 0 9 13 13 1 9 9 2
30 3 7 13 13 2 16 0 9 1 0 2 0 9 9 13 3 1 0 9 2 1 15 4 13 4 10 9 3 13 2
57 1 9 2 16 4 0 9 9 13 2 13 0 9 13 1 9 0 9 2 1 9 2 16 9 13 13 7 1 10 9 1 9 0 9 7 16 13 7 3 13 9 1 0 9 7 1 0 9 1 9 2 1 15 13 0 9 2
21 16 15 10 9 13 16 0 2 13 12 1 9 2 3 9 13 2 0 9 9 2
16 10 9 9 1 9 0 0 9 13 13 1 10 9 9 9 2
35 16 15 9 13 1 9 0 0 9 1 0 9 9 2 7 9 2 9 7 9 1 0 9 2 7 9 1 3 9 2 13 9 0 9 2
27 1 10 9 3 13 13 0 2 9 9 2 15 15 13 9 9 9 1 10 9 7 9 9 1 10 9 2
31 1 10 9 13 0 13 2 16 0 0 9 13 1 10 9 0 10 9 7 3 9 13 9 1 9 9 9 0 7 0 2
33 1 10 9 15 13 13 2 16 9 9 4 13 9 7 1 9 2 7 1 9 2 15 7 15 2 7 7 1 9 7 9 3 2
9 9 9 13 13 1 12 0 9 2
19 9 9 13 0 2 0 9 2 15 13 13 3 9 0 2 3 9 0 2
13 1 10 9 15 3 9 0 0 9 13 0 9 2
29 2 3 15 1 0 0 9 13 9 15 9 2 15 13 0 9 2 0 1 9 3 13 3 3 9 10 9 2 2
12 2 3 15 9 0 9 13 1 9 0 9 2
35 1 9 2 16 4 3 0 9 13 7 1 9 9 9 2 13 15 0 9 10 9 7 0 9 15 3 13 1 0 9 1 3 0 9 2
8 1 9 15 9 13 0 9 2
14 13 13 2 16 9 9 1 0 9 13 9 1 9 2
35 10 9 9 9 2 15 13 13 1 12 0 9 2 13 7 3 0 9 7 1 9 12 10 0 9 13 0 9 13 9 0 9 3 3 2
14 0 9 13 0 13 14 1 0 9 0 9 0 9 2
2 9 9
11 1 9 9 4 13 9 1 3 0 9 2
14 12 1 9 13 2 7 13 2 16 15 0 9 13 2
17 16 4 1 15 13 9 2 3 15 13 2 16 1 15 13 9 2
3 13 9 2
7 3 13 10 9 13 3 2
7 11 2 11 2 2 0 11
26 10 9 13 13 9 12 0 9 1 0 9 2 3 0 9 9 7 9 13 13 1 9 12 7 12 2
14 1 10 9 13 1 10 9 9 1 0 9 3 0 2
16 15 13 2 16 15 13 13 9 10 9 1 9 9 0 9 2
17 10 9 15 7 13 9 13 3 7 3 1 10 9 13 0 9 2
32 1 9 13 2 16 0 9 13 9 1 9 2 9 7 9 1 9 7 9 1 3 0 0 9 2 15 13 3 0 0 9 2
31 1 9 12 0 9 10 9 0 9 3 0 9 13 2 13 2 14 1 0 9 2 15 13 9 2 7 15 4 3 13 2
2 11 11
29 9 13 0 9 11 2 11 2 0 12 9 2 12 12 11 12 2 11 2 9 2 2 2 12 2 12 12 12 2
5 13 9 9 2 12
8 15 13 13 11 3 7 3 2
8 9 0 13 9 1 0 9 2
18 0 9 11 11 13 3 2 16 4 13 3 13 2 15 13 1 9 2
4 9 9 13 2
7 2 9 1 9 3 13 2
10 1 10 0 0 9 15 11 11 13 2
16 2 11 11 2 0 9 7 9 1 11 2 3 0 13 15 2
6 2 9 12 9 0 11
13 2 0 9 1 9 2 2 9 13 16 0 9 2
5 2 9 11 11 2
4 9 2 0 9
6 9 9 9 9 1 9
2 9 2
4 0 9 2 12
4 0 9 2 12
12 9 9 2 9 0 9 2 9 2 0 9 2
4 0 9 2 12
4 0 9 2 12
17 9 0 9 2 0 7 9 0 9 2 0 9 2 0 9 9 2
8 0 9 2 12 2 12 9 2
8 0 9 2 12 2 12 9 2
27 9 13 13 9 9 2 1 0 7 0 9 7 9 2 9 9 1 9 7 9 9 1 0 2 0 9 2
7 10 9 4 13 9 9 2
20 13 13 15 1 0 9 0 9 2 15 4 13 0 7 10 9 1 9 9 2
10 0 9 1 9 13 13 9 13 9 2
38 1 9 13 15 0 2 16 1 15 13 0 9 2 9 2 1 15 15 13 1 12 9 2 4 15 3 13 13 2 13 11 11 1 0 9 0 9 2
3 9 13 9
18 1 9 12 13 0 0 9 11 1 11 10 9 3 3 7 9 3 2
21 9 13 1 12 9 9 2 15 13 1 9 9 7 9 3 3 16 1 12 9 2
17 1 0 9 11 11 4 13 1 15 2 15 15 1 10 9 13 2
10 2 3 9 13 1 9 0 0 9 2
16 13 4 3 1 15 2 1 9 13 14 15 2 15 3 13 2
9 15 13 3 9 9 9 11 11 2
16 7 15 4 1 9 9 13 9 0 9 2 3 3 13 9 2
19 7 1 0 0 9 4 13 9 2 16 9 1 9 13 3 3 16 9 2
18 7 4 13 1 9 2 0 9 2 0 9 2 0 9 7 0 9 2
11 2 1 15 13 2 16 1 15 13 0 2
5 0 9 13 9 2
8 0 9 15 1 15 13 13 2
15 9 3 13 13 13 9 0 0 9 2 7 0 9 13 2
8 0 9 9 13 9 1 9 2
19 3 10 0 9 13 0 9 12 9 2 15 15 13 13 7 10 0 9 2
15 13 4 15 3 9 11 7 13 13 10 0 9 1 9 2
11 0 9 11 15 13 1 11 1 10 9 2
9 2 13 15 9 3 9 7 9 2
7 13 4 15 13 0 9 2
16 3 4 13 1 9 14 13 9 9 9 7 1 9 15 13 2
5 3 13 9 0 2
6 7 4 13 0 9 2
14 13 4 3 9 0 9 2 13 9 0 9 7 9 2
18 1 9 15 4 3 13 9 1 9 0 9 2 16 0 9 13 0 2
18 13 4 12 9 9 1 9 0 9 2 13 9 7 9 0 9 13 2
9 2 1 10 9 13 9 0 9 2
5 3 4 13 9 2
11 3 4 1 9 12 3 13 1 15 0 2
15 9 11 13 1 0 9 2 16 15 13 1 0 0 9 2
15 10 0 9 13 0 9 2 15 1 0 9 13 0 9 2
10 15 13 1 9 9 1 12 9 9 2
10 0 12 9 0 13 9 1 0 9 2
17 1 0 13 9 13 3 2 7 16 0 9 13 1 9 0 9 2
15 10 9 13 2 16 1 0 9 11 15 9 13 1 9 2
11 13 7 9 1 9 9 1 10 0 9 2
2 11 0
7 3 13 9 2 3 13 9
7 9 9 13 0 9 1 9
24 0 9 1 9 9 7 9 13 1 15 2 16 4 15 13 3 13 0 0 9 1 0 9 2
16 13 7 9 7 0 0 9 2 9 2 9 2 9 2 9 2
8 1 9 4 3 13 13 9 2
14 0 0 9 13 3 13 2 3 15 3 3 10 13 2
20 0 9 1 9 13 1 0 9 3 1 9 9 9 12 11 2 9 2 11 2
2 11 11
13 0 9 1 9 1 9 13 13 0 9 0 9 2
17 1 9 15 3 13 13 3 2 1 0 9 15 9 9 3 13 2
34 13 2 14 3 1 0 9 1 11 7 11 1 9 12 7 12 9 3 2 13 15 3 1 9 9 14 12 9 12 7 12 0 9 2
5 7 15 13 9 2
32 1 10 9 15 3 13 13 9 2 9 7 9 3 2 16 3 1 11 7 0 1 0 11 2 3 13 12 9 1 12 9 2
9 0 0 9 9 13 1 9 12 2
12 1 0 12 9 15 7 1 0 9 13 9 2
16 7 15 1 9 0 9 13 0 9 1 9 7 1 10 9 2
2 0 9
13 15 13 0 9 9 9 1 9 12 1 9 12 2
13 1 0 9 1 11 2 3 11 2 13 9 9 2
8 3 9 13 15 9 1 11 2
16 3 1 0 0 9 9 9 3 13 2 3 16 1 0 11 2
26 3 13 13 9 9 7 1 0 9 9 3 1 0 11 2 13 11 11 2 9 9 9 0 9 11 2
5 9 13 0 9 2
18 1 0 9 13 0 9 11 2 11 2 11 2 11 2 11 2 11 2
14 9 15 3 13 1 0 9 1 11 2 3 3 13 2
14 3 1 0 9 1 11 13 9 9 14 1 0 9 2
3 0 12 9
23 1 9 0 9 13 9 9 2 9 12 7 12 2 1 9 9 9 7 9 1 9 12 2
21 0 9 13 1 11 11 0 7 13 1 10 9 1 9 12 9 9 1 9 12 2
12 1 10 9 4 13 4 13 15 0 9 9 2
14 9 1 0 9 4 13 4 13 1 12 7 12 5 2
16 13 15 1 9 0 9 2 16 3 13 3 0 2 3 13 2
22 3 15 13 3 3 1 11 2 15 13 1 10 9 1 9 0 9 1 0 9 9 2
14 1 0 9 4 3 14 13 13 3 9 0 1 9 2
41 1 9 4 15 13 13 1 11 14 1 0 11 2 1 9 12 3 13 0 9 1 9 11 2 9 2 13 4 13 4 7 9 9 12 1 11 1 11 1 11 2
25 9 9 12 11 2 11 11 4 15 13 13 14 1 11 7 9 9 12 11 2 11 14 1 11 2
45 1 9 4 13 4 13 9 0 11 2 11 2 9 1 11 2 9 9 2 12 2 2 3 9 9 1 11 2 11 2 0 11 2 11 2 9 2 12 2 7 11 11 2 11 2
22 13 2 14 0 9 9 0 9 1 15 2 15 13 13 1 9 12 2 3 15 13 2
18 13 7 9 1 9 2 3 13 13 0 9 2 13 13 3 0 9 2
7 13 9 9 15 3 13 2
2 12 0
38 1 9 11 13 1 9 12 9 9 7 12 9 9 2 1 10 13 12 9 9 12 2 9 2 12 9 9 12 2 9 7 12 9 9 12 2 9 2
10 0 9 13 12 9 0 0 0 9 2
12 9 0 9 9 13 1 0 9 9 12 9 2
18 0 9 2 3 13 1 0 9 3 9 0 9 2 13 9 12 9 2
10 1 10 9 13 1 9 3 0 9 2
40 1 9 9 7 13 14 12 9 9 7 9 1 9 9 0 16 12 9 1 9 2 16 1 0 9 9 13 9 14 12 9 1 9 2 1 9 12 9 3 2
34 1 0 9 9 9 0 9 3 13 2 16 1 9 12 1 9 1 9 12 13 9 3 1 12 5 7 1 0 9 3 1 12 5 2
12 9 1 9 13 7 0 9 14 1 0 9 2
22 1 9 0 9 13 12 9 1 9 0 0 9 1 0 12 9 9 1 11 7 11 2
56 13 2 14 1 9 2 16 4 15 15 1 10 9 13 2 7 1 11 3 13 0 9 9 7 10 9 13 2 2 1 9 0 9 13 3 0 2 16 0 9 13 1 9 7 9 9 2 3 0 0 9 7 9 0 9 2
13 7 3 10 9 13 13 10 9 1 9 7 9 2
5 9 13 1 9 2
8 9 13 1 9 9 1 0 9
30 13 15 2 16 9 2 0 9 9 0 9 1 9 0 2 13 0 9 2 9 0 9 13 7 3 7 3 3 13 2
15 7 9 0 9 2 0 9 9 1 12 9 2 13 0 2
31 0 9 3 13 9 1 3 9 9 2 16 0 11 3 2 11 3 2 11 3 2 11 3 7 9 9 3 14 3 3 2
2 11 11
22 13 7 7 0 2 0 9 2 7 3 16 0 9 13 12 1 12 9 0 0 9 2
16 3 7 9 2 16 9 3 13 2 13 1 0 9 13 3 2
29 3 0 0 9 9 1 9 13 14 3 13 0 9 2 16 13 1 9 3 3 3 2 7 3 14 1 0 9 2
34 0 9 2 16 13 1 9 9 9 7 9 1 3 3 0 9 2 13 3 0 10 9 13 2 16 3 7 3 15 1 15 3 13 2
20 13 15 7 1 15 2 15 0 15 1 10 0 0 9 1 0 3 9 13 2
49 0 2 16 10 9 2 15 13 13 0 9 1 9 2 13 15 7 15 2 0 9 2 2 3 1 9 9 4 13 9 9 2 3 9 9 7 3 9 0 9 2 15 1 0 3 0 9 9 2
21 13 3 2 16 0 0 9 15 2 1 15 9 7 9 2 1 9 1 12 13 2
23 1 9 1 15 12 0 9 2 0 0 9 13 3 9 0 9 9 2 3 0 9 9 2
9 9 13 2 3 13 10 9 0 2
2 9 9
51 0 9 2 10 9 0 9 2 13 7 13 1 3 0 9 2 15 13 9 7 9 9 1 10 9 3 1 9 2 3 1 9 2 3 12 0 0 9 2 1 15 13 12 0 9 1 0 2 9 9 2
26 7 3 13 2 16 15 13 0 11 3 9 2 0 3 9 0 9 2 3 16 9 0 9 1 0 2
34 3 15 13 0 9 2 0 9 2 3 15 13 9 9 2 3 0 9 2 1 12 1 0 12 2 12 5 1 0 12 12 9 2 2
37 7 3 13 0 2 16 3 7 3 4 13 13 1 0 9 1 9 1 9 2 3 15 1 0 9 9 0 0 9 4 13 3 13 3 3 9 2
35 16 15 13 0 9 0 9 2 7 9 2 2 7 9 9 0 2 16 0 9 1 9 9 2 13 1 10 9 1 0 9 0 14 3 2
29 13 3 0 9 3 0 9 1 0 9 2 7 3 3 15 13 9 0 9 16 9 1 9 3 0 2 7 0 2
21 9 2 15 1 0 9 13 0 9 2 4 1 0 9 3 3 13 2 3 3 2
3 1 9 9
47 9 2 0 9 1 0 9 1 9 12 2 9 7 1 0 12 9 2 3 1 0 9 11 9 13 1 12 5 1 9 3 2 2 13 2 13 15 2 1 0 9 12 2 9 3 13 2
38 0 9 1 12 7 12 5 0 0 0 9 9 15 13 13 10 9 2 15 13 1 0 9 13 0 9 9 1 0 9 2 3 16 13 0 9 9 2
37 3 15 15 13 2 16 0 9 1 9 2 7 3 1 9 2 13 0 9 1 3 0 9 0 9 0 9 9 0 9 1 10 0 7 0 9 2
26 9 15 3 13 2 7 9 1 0 9 0 9 2 3 7 3 0 9 1 0 9 9 3 13 9 2
22 14 0 9 13 2 16 13 3 0 9 2 16 15 1 0 9 13 3 0 9 9 2
15 9 2 3 0 0 9 4 13 0 9 2 13 14 0 2
2 9 9
21 0 9 2 0 1 0 9 13 9 1 9 9 7 9 2 13 0 9 0 9 2
30 13 13 2 16 9 2 3 13 1 0 9 1 9 0 9 2 3 7 3 3 10 2 0 9 2 13 1 9 9 2
15 3 2 1 9 0 9 2 13 1 9 1 9 0 9 2
25 9 2 16 0 9 13 10 0 2 15 13 9 13 1 9 9 2 3 1 0 9 13 0 9 2
3 9 9 2
4 9 0 9 2
6 15 12 9 13 13 3
12 2 0 9 11 12 2 12 2 9 1 9 2
2 9 2
17 0 11 1 11 1 12 2 12 2 0 2 11 2 2 0 11 12
6 11 0 11 9 2 12
4 9 2 9 9
2 13 0
25 9 9 0 0 9 11 13 1 9 12 2 3 0 9 9 0 0 1 11 13 9 1 9 11 2
15 3 15 9 2 9 9 2 9 2 9 2 13 1 0 2
25 9 1 10 9 3 13 0 9 2 9 9 2 9 0 9 2 0 9 7 9 9 7 0 9 2
23 16 15 0 9 7 9 9 3 13 2 14 1 0 12 9 3 2 13 15 7 9 9 2
32 15 3 13 1 9 0 9 7 9 7 9 0 9 7 9 1 11 7 0 11 2 7 7 9 7 9 9 1 11 7 11 2
18 13 7 9 2 3 15 13 0 0 0 9 2 9 2 9 2 9 2
18 3 0 9 9 13 7 9 9 0 9 7 0 9 1 9 7 9 2
10 0 9 9 9 13 9 9 7 9 2
27 9 2 9 0 0 9 11 2 0 12 2 11 12 12 2 9 2 7 9 2 2 12 2 12 2 12 2
3 9 0 9
13 9 13 1 0 0 9 0 9 1 9 12 2 12
39 1 9 11 7 9 1 0 9 11 13 0 0 9 2 15 13 0 7 0 9 9 9 1 0 9 7 9 2 3 3 9 0 0 9 3 7 1 9 2
34 13 15 14 1 0 0 9 1 0 9 9 0 9 2 7 13 13 1 9 7 10 0 9 2 3 9 9 10 0 0 9 2 11 2
12 0 9 3 1 0 9 13 3 1 0 9 2
9 1 10 9 3 13 3 12 9 2
27 2 9 7 9 10 9 2 1 9 0 0 9 2 3 14 9 2 4 7 13 3 9 0 7 0 9 2
35 2 0 9 9 13 1 0 2 7 0 9 13 1 9 9 9 0 9 2 14 3 13 1 9 2 7 9 2 2 0 3 1 9 9 2
3 3 3 9
28 1 10 0 9 13 13 2 16 3 15 13 9 9 2 15 9 15 13 3 14 14 1 9 9 1 0 9 2
27 1 0 9 1 9 2 15 13 10 0 0 9 2 9 0 2 9 7 0 9 0 9 15 0 9 13 2
20 3 3 13 0 0 9 2 3 1 12 2 9 2 2 16 4 13 0 9 2
21 15 1 0 9 1 9 9 9 7 9 13 1 12 2 9 3 1 3 0 9 2
11 13 3 3 12 9 2 15 4 3 13 2
29 1 9 9 9 12 1 9 0 13 0 13 0 9 1 0 9 9 2 15 15 13 7 13 3 0 9 0 9 2
39 13 1 0 7 0 9 0 2 1 9 9 1 10 9 3 2 7 0 9 2 16 7 9 1 11 1 15 9 9 12 2 1 0 9 9 0 15 9 2
25 0 9 9 12 3 13 9 3 0 9 14 1 12 2 9 12 2 7 3 7 1 0 9 12 2
5 3 3 7 3 2
14 1 9 12 2 12 15 13 0 9 0 9 0 9 2
18 9 0 0 9 11 2 1 11 2 4 13 1 9 1 9 7 9 2
11 0 9 9 0 2 9 4 3 3 13 2
51 3 13 7 0 13 0 9 0 9 2 3 9 0 9 7 0 9 0 9 1 11 1 11 2 7 0 9 1 0 9 13 15 1 9 1 9 0 0 9 14 9 2 2 1 0 9 1 9 9 11 2
15 0 9 4 15 1 10 9 13 13 0 9 1 9 9 2
20 3 9 0 9 4 3 13 2 3 7 4 13 0 9 9 7 9 0 9 2
27 0 9 1 9 1 0 9 13 3 0 2 16 0 9 1 9 1 0 9 0 9 4 13 13 3 0 2
29 9 0 9 0 9 0 9 7 9 0 9 0 9 13 3 0 9 2 1 15 15 13 10 0 9 9 9 9 2
24 15 4 15 13 1 0 9 13 9 12 2 12 5 7 1 0 9 9 14 12 2 12 5 2
29 15 13 0 9 2 1 15 15 3 13 9 1 9 9 9 2 9 7 0 9 0 9 0 9 1 0 12 9 2
7 11 11 2 0 0 9 2
8 11 11 2 9 1 0 9 11
9 9 9 9 9 1 9 12 2 12
5 0 9 1 12 9
10 11 13 1 9 0 9 13 1 0 9
14 0 9 11 11 13 1 0 9 0 9 3 1 9 2
8 1 10 0 9 1 15 13 2
2 11 11
9 0 9 11 13 1 12 9 9 2
30 0 9 13 2 16 12 5 9 13 9 0 9 2 12 5 13 1 9 2 12 5 1 0 7 12 5 0 0 9 2
6 0 9 15 13 9 2
13 1 9 9 4 15 3 13 13 3 1 9 12 2
8 9 11 1 9 12 13 0 2
13 9 13 1 12 9 9 2 9 13 1 12 9 2
9 9 1 9 13 1 12 9 9 2
3 9 1 9
28 13 13 2 16 1 0 9 2 15 3 13 1 0 9 2 13 9 7 1 9 0 9 13 1 10 9 9 2
26 0 9 9 11 7 13 3 13 1 15 2 16 9 13 1 9 12 9 13 9 7 15 9 13 13 2
8 0 9 3 13 1 0 9 2
21 1 9 10 9 13 0 12 12 9 9 2 7 15 9 1 15 12 5 9 13 2
28 0 9 3 13 2 12 5 9 0 9 2 12 5 0 9 2 12 5 0 7 0 9 2 12 5 0 9 2
28 15 13 3 13 0 9 9 2 15 13 9 3 1 9 12 13 9 0 9 7 13 0 9 1 9 0 9 2
9 15 15 13 9 14 12 9 9 2
19 9 3 3 4 13 7 9 1 9 2 1 9 15 13 7 1 9 9 2
4 15 13 9 2
10 1 10 9 13 0 9 3 3 13 2
8 13 3 7 0 7 10 9 2
5 3 15 13 9 2
22 9 9 11 11 11 15 3 13 15 2 16 13 13 13 1 9 0 9 0 0 9 2
24 3 4 13 0 9 13 1 0 9 0 9 0 9 2 15 13 0 9 7 4 13 0 9 2
13 11 13 1 0 2 0 9 9 3 13 10 9 2
21 3 13 2 13 0 9 9 0 9 2 7 7 13 3 0 0 9 1 0 9 2
38 3 13 2 9 13 9 1 0 9 0 0 9 2 7 13 15 9 1 15 2 15 13 0 9 9 2 3 0 9 2 7 9 1 0 7 0 9 2
22 16 13 0 9 13 9 1 0 9 2 13 3 13 14 0 2 7 0 9 1 9 2
17 3 16 4 13 14 1 0 9 2 13 3 13 9 9 14 3 2
7 10 9 4 13 3 9 2
20 4 15 7 3 13 1 9 2 15 13 3 9 2 7 15 7 0 7 0 2
23 3 13 13 2 16 13 9 3 1 9 0 0 9 2 3 7 0 0 9 7 0 9 2
25 11 4 15 3 13 13 9 0 9 2 1 0 2 2 1 9 2 10 0 0 9 10 9 13 2
20 13 4 9 13 7 13 0 9 2 16 4 1 9 13 7 4 13 3 0 2
9 3 4 3 7 15 13 13 9 2
14 15 4 3 13 7 9 1 10 9 1 9 0 9 2
26 1 0 9 2 7 16 4 9 2 15 4 13 2 13 2 13 13 9 11 1 9 0 9 3 0 2
4 9 1 0 9
5 9 13 3 9 2
5 9 13 13 0 9
20 9 9 0 9 11 1 0 9 15 13 0 9 11 2 11 2 11 7 11 2
25 0 9 15 1 9 11 7 11 13 1 9 9 0 9 7 0 9 7 15 1 0 7 0 9 2
27 1 15 13 0 9 3 1 0 0 9 2 15 13 0 10 9 2 9 7 0 9 2 13 9 11 11 2
3 9 1 9
21 1 11 13 1 9 0 2 7 15 7 3 2 16 7 3 13 1 0 9 9 2
31 16 1 9 12 15 13 12 2 15 13 9 9 9 14 1 12 7 12 9 2 3 1 0 9 4 15 13 13 3 12 2
27 3 2 16 1 15 2 16 4 15 3 3 13 9 9 2 15 15 3 13 13 2 4 0 0 9 13 2
7 0 9 3 13 9 9 2
16 0 15 3 13 2 16 9 10 9 13 13 1 9 0 9 2
34 15 4 13 9 1 0 9 2 7 15 7 3 2 16 9 13 1 0 9 14 3 3 2 16 13 9 1 0 9 1 9 0 9 2
19 9 9 15 3 13 2 16 0 9 13 13 14 0 2 3 0 9 9 2
11 1 0 9 13 3 1 9 0 9 9 2
17 13 1 15 9 2 16 9 0 0 9 13 1 11 14 12 9 2
2 0 9
15 9 9 11 13 2 16 1 0 9 13 0 9 1 0 2
9 13 1 9 12 9 1 12 9 2
22 1 10 9 2 3 7 9 1 9 0 9 2 13 1 11 0 9 1 15 0 9 2
13 9 13 13 15 2 16 4 15 3 9 3 13 2
26 15 4 13 2 1 9 9 9 2 13 3 0 9 7 9 2 3 7 0 9 2 15 10 9 13 2
19 0 9 13 2 16 4 15 11 13 0 0 9 1 0 9 9 0 9 2
28 16 4 9 1 0 9 13 9 1 15 2 3 13 1 9 1 0 9 2 3 1 9 1 9 9 9 3 2
22 3 4 13 13 15 13 7 0 9 2 7 15 4 3 13 1 9 2 13 11 11 2
21 0 9 2 3 13 9 2 13 7 0 2 0 9 10 9 2 15 13 3 13 2
3 9 1 9
12 3 15 3 1 9 13 1 0 9 1 9 2
7 0 9 15 7 3 13 2
16 10 0 9 15 13 13 1 12 9 2 7 3 1 12 9 2
8 7 15 9 9 11 13 1 2
16 1 9 1 0 9 15 13 13 9 10 0 9 1 10 9 2
13 13 1 12 2 12 2 12 9 2 13 0 9 2
12 13 15 3 1 9 9 7 13 1 0 9 2
19 1 10 9 15 13 2 16 15 1 15 3 0 9 13 9 2 7 3 2
28 1 9 9 7 9 9 13 1 11 13 10 9 7 1 0 9 2 3 1 9 0 9 2 3 1 0 9 2
2 0 9
21 1 0 9 13 13 0 9 2 3 15 13 0 0 9 1 0 9 9 0 9 2
16 7 16 13 14 1 0 9 2 13 15 15 15 1 0 9 2
35 9 2 9 11 1 11 2 0 2 9 2 2 0 9 2 11 12 2 12 12 11 2 9 2 12 2 12 2 9 2 12 2 12 12 2
2 9 2
11 0 9 13 13 14 0 2 3 0 9 9
3 9 9 2
3 3 15 13
7 1 9 9 3 9 3 13
9 9 9 13 1 9 12 3 3 2
13 1 12 2 12 2 12 13 9 12 9 1 9 2
8 1 9 0 9 3 12 9 2
29 1 12 2 9 12 13 1 9 12 0 13 12 9 1 0 9 2 1 9 0 1 9 1 9 12 9 2 9 2
2 11 11
4 9 13 13 2
5 9 9 13 3 2
7 9 9 1 9 14 13 2
15 1 9 13 9 2 9 9 2 10 9 7 1 9 9 2
2 0 9
9 9 1 9 13 1 9 9 0 2
9 0 9 3 9 9 9 9 13 2
3 13 0 2
32 1 0 9 1 11 2 11 13 13 2 16 1 9 12 9 1 9 7 0 9 13 1 9 1 9 7 9 1 12 12 9 2
11 0 9 1 9 15 3 13 12 9 9 2
11 12 9 1 9 3 9 13 14 1 9 2
7 1 0 9 15 13 0 2
19 9 13 9 9 1 9 7 13 15 3 13 2 16 10 9 3 13 9 2
15 9 13 1 0 9 2 16 1 10 9 1 9 13 0 2
2 0 9
13 0 9 2 0 15 3 9 2 13 1 12 5 2
18 13 0 13 2 16 13 9 9 9 2 0 10 9 4 3 3 13 2
9 7 3 0 9 4 13 1 9 2
22 16 4 15 3 9 1 9 13 3 2 13 4 3 1 10 9 13 7 1 12 5 2
14 9 1 9 9 15 13 1 9 1 12 9 1 9 2
19 7 13 9 9 2 15 15 13 1 12 9 2 0 3 14 1 12 9 2
5 7 13 0 13 2
5 3 13 7 9 2
8 3 0 9 13 3 3 3 2
18 9 9 1 0 9 13 9 2 16 4 15 10 0 9 1 9 13 2
17 7 3 15 3 13 3 9 2 16 4 13 1 0 9 15 13 2
14 9 9 13 3 2 16 15 13 7 13 1 0 9 2
11 1 0 9 1 9 15 13 3 13 13 2
14 0 9 9 13 2 16 9 15 13 7 9 13 0 2
9 0 9 13 1 10 9 1 0 2
15 13 13 2 16 3 9 1 9 1 0 9 1 9 13 2
10 13 4 9 9 3 13 7 3 13 2
16 7 7 10 9 1 9 9 1 9 13 3 0 2 13 0 2
13 13 1 9 12 2 12 2 0 9 9 9 9 13
2 9 2
4 13 0 9 2
5 3 13 3 0 2
11 0 15 13 1 10 9 1 9 1 9 2
8 15 13 1 12 0 9 9 2
18 16 4 15 15 13 2 3 15 3 16 0 9 4 1 9 13 9 2
4 0 9 7 15
20 0 9 11 13 14 1 12 9 2 3 15 13 13 9 9 1 9 0 9 2
16 1 9 13 1 12 9 7 13 0 9 12 7 12 9 9 2
13 3 13 1 12 9 7 13 1 3 16 12 9 2
8 9 13 1 11 1 9 11 2
16 9 3 13 9 1 9 2 0 9 7 9 1 9 0 9 2
11 0 9 13 0 0 9 7 0 0 9 2
17 9 0 9 13 9 0 9 2 15 13 0 9 1 12 9 9 2
29 13 15 3 1 9 0 9 1 12 1 12 9 2 0 9 1 12 1 12 9 7 0 9 1 12 1 12 9 2
8 1 11 9 13 1 9 12 2
42 1 0 0 9 4 3 13 9 1 9 0 7 0 9 7 0 9 1 0 9 11 1 12 9 9 9 2 13 11 11 2 0 9 11 0 11 9 2 9 2 0 2
19 0 9 3 13 11 1 0 0 9 1 11 7 3 15 13 1 9 11 2
42 9 2 11 0 0 11 9 2 9 2 0 2 2 0 12 2 12 12 11 12 2 9 2 2 2 12 2 12 12 12 12 2 9 2 2 12 2 12 12 12 12 2
4 9 1 0 9
14 1 9 13 1 9 9 1 9 1 9 7 0 1 9
12 1 0 9 13 1 9 9 14 12 9 9 2
34 3 12 9 9 13 0 2 12 9 0 2 12 9 0 2 12 9 0 9 13 0 0 9 2 7 3 2 12 9 2 13 0 9 2
2 11 11
42 13 7 0 9 2 16 1 12 2 9 15 10 0 9 3 13 2 7 15 9 9 9 9 1 9 1 9 7 0 9 2 15 1 9 12 2 9 13 9 9 11 2
18 1 0 9 15 3 13 2 16 1 0 9 4 13 3 12 0 9 2
18 1 9 0 9 9 0 9 1 0 9 3 3 13 9 9 0 9 2
12 13 15 7 1 9 1 0 9 0 0 9 2
4 12 2 0 9
35 9 2 9 9 15 13 9 2 9 1 9 0 9 4 9 13 2 15 13 2 16 1 9 15 13 3 0 9 0 0 7 0 9 2 2
37 9 2 1 9 15 4 13 7 9 2 16 10 9 15 13 9 2 9 1 9 0 9 9 1 9 2 1 15 13 0 0 9 2 9 13 2 2
34 9 2 9 13 1 9 9 10 9 2 7 10 0 0 9 2 3 15 13 2 16 1 9 9 15 13 9 9 2 3 7 9 2 2
27 9 2 0 9 9 13 13 3 0 0 9 2 9 7 13 9 9 2 16 4 0 9 13 1 9 2 2
42 9 2 13 2 14 15 9 2 16 9 13 2 13 15 13 0 9 9 2 13 15 2 16 9 13 10 0 9 3 1 12 12 7 9 15 13 3 1 10 9 2 2
36 9 2 9 13 12 9 1 15 2 16 4 15 1 9 9 1 9 9 13 2 16 15 13 2 1 9 10 9 13 9 13 9 15 0 2 2
46 9 2 13 2 14 9 1 9 1 9 12 9 2 13 3 1 9 0 12 9 3 13 9 1 9 2 1 15 13 0 9 2 3 4 13 3 0 0 9 2 9 15 7 13 2 2
37 9 2 13 2 14 15 9 2 16 9 13 2 13 3 10 9 2 13 13 4 3 1 9 0 9 2 16 10 9 0 1 0 9 13 13 2 2
18 9 2 9 9 15 13 9 0 9 1 9 1 9 1 9 10 9 2
37 9 2 9 2 9 7 9 0 9 13 9 2 0 7 0 9 2 15 13 9 9 2 0 9 9 13 1 10 9 13 0 9 1 0 9 2 2
4 12 2 0 9
18 9 2 9 11 7 11 13 13 14 1 9 9 2 1 0 9 2 2
18 9 2 9 15 13 2 13 15 1 9 2 16 13 1 9 9 2 2
27 9 2 9 0 9 2 7 7 9 7 9 15 13 3 2 15 7 13 9 13 9 9 0 1 9 2 2
42 9 2 1 9 2 16 9 3 1 9 13 9 1 9 9 2 7 3 13 1 12 2 9 12 2 13 9 9 13 1 15 3 1 12 2 9 12 9 1 9 9 2
26 9 2 1 9 9 13 9 9 2 15 4 13 1 0 0 9 9 7 1 0 9 9 1 0 9 2
35 9 2 9 9 1 9 13 9 1 9 2 9 0 9 9 7 13 13 3 0 0 9 7 9 9 13 1 12 9 13 0 0 9 2 2
36 9 2 1 9 13 9 9 9 1 0 9 2 15 15 13 16 9 1 15 9 9 1 0 0 9 7 9 13 4 13 3 1 12 9 2 2
27 9 2 1 12 2 9 12 13 0 9 13 1 0 9 1 9 7 9 0 9 2 3 0 9 9 2 2
6 9 9 2 2 9 2
4 9 13 1 9
32 9 1 0 9 0 9 2 9 0 9 1 15 9 2 9 9 9 0 7 0 9 2 15 13 9 2 1 15 9 3 13 2
13 1 9 1 0 9 13 1 10 9 0 0 9 2
17 7 4 15 10 9 9 13 2 15 15 3 13 7 15 13 13 2
6 11 11 2 11 11 2
12 13 15 9 9 13 1 9 0 9 0 9 2
24 13 1 15 2 16 1 0 9 13 9 2 16 13 9 2 15 4 13 1 0 9 9 9 2
15 15 13 7 9 1 0 9 2 3 1 12 0 9 9 2
22 7 13 3 1 9 0 9 2 16 13 0 9 2 1 9 9 2 3 13 9 0 2
6 15 4 15 13 13 2
6 11 11 2 11 11 2
6 13 15 0 0 9 2
19 13 15 2 16 13 0 2 16 0 9 13 1 9 2 15 13 1 9 2
19 1 15 4 13 4 13 1 15 9 2 7 7 15 0 13 9 7 9 2
27 3 4 15 13 12 9 2 16 1 3 0 9 9 4 0 9 13 13 0 2 16 4 15 13 3 9 2
11 13 4 15 7 3 9 1 9 0 9 2
6 11 11 2 9 11 2
13 3 4 15 13 13 0 7 0 9 1 12 9 2
9 13 4 15 3 9 1 15 0 2
13 13 4 7 9 1 9 2 15 3 13 1 9 2
6 11 11 2 11 11 2
15 15 16 9 3 13 9 1 9 2 15 13 9 3 13 2
9 3 1 9 9 3 13 0 9 2
22 3 1 0 9 4 1 12 13 12 9 1 0 9 2 7 9 10 12 9 15 13 2
4 15 13 0 2
2 0 9
18 9 9 0 9 11 11 16 0 1 9 13 9 9 9 1 11 12 2
28 15 13 0 9 2 3 4 13 10 9 11 11 2 9 10 9 2 1 10 0 9 13 3 0 9 0 9 2
10 2 15 15 13 1 0 9 0 9 2
10 0 9 9 1 9 13 9 9 9 2
5 1 15 13 13 2
18 16 4 15 13 2 13 4 13 1 10 9 7 10 9 7 0 9 2
15 3 13 9 12 9 9 7 4 13 3 9 1 0 9 2
16 0 9 13 0 2 7 3 0 12 9 9 13 1 0 9 2
23 15 2 16 15 15 13 13 0 9 1 0 9 11 2 13 4 1 9 13 0 0 9 2
19 3 4 13 12 9 9 7 12 9 9 9 13 3 2 3 15 9 13 2
9 3 3 15 13 9 9 11 12 2
7 13 4 15 3 12 9 2
14 3 4 13 1 0 9 13 3 9 9 7 15 9 2
7 1 9 12 4 9 13 2
7 9 7 3 3 13 9 2
15 13 1 9 2 15 13 13 2 16 1 9 13 0 9 2
13 1 0 9 13 15 9 2 16 13 9 0 9 2
8 2 15 15 13 1 0 9 2
26 3 4 13 9 13 1 15 2 15 9 9 9 9 13 7 15 1 10 9 13 0 1 10 9 13 2
5 1 9 13 9 2
9 2 3 4 15 3 13 9 9 2
18 13 4 1 0 9 7 13 15 2 4 13 3 16 4 13 1 9 2
14 9 9 3 13 2 16 4 9 3 3 13 0 9 2
14 16 13 0 9 2 13 9 7 4 9 13 1 9 2
6 15 13 13 0 9 2
17 7 3 13 15 0 1 0 9 2 15 13 2 16 15 15 13 2
10 2 3 15 9 9 9 13 1 9 2
12 0 13 13 15 3 2 16 4 13 0 9 2
7 9 9 13 1 0 9 2
13 3 4 15 13 2 10 9 4 1 0 9 13 2
22 3 13 13 0 9 2 3 4 13 15 0 9 2 9 2 9 2 9 9 7 3 2
21 0 13 13 9 0 9 1 9 7 0 9 1 9 2 16 4 9 13 0 9 2
8 3 4 13 12 9 0 9 2
11 13 15 9 2 16 15 15 3 3 13 2
9 7 1 9 4 15 9 13 3 2
6 9 2 0 9 7 15
1 11
16 0 9 1 0 9 13 3 1 9 12 9 9 11 1 11 2
19 13 7 9 2 16 1 9 13 0 9 0 9 7 9 1 9 9 11 2
10 0 9 9 15 13 1 12 9 9 2
21 0 9 9 13 9 2 16 1 0 12 12 9 13 9 9 14 1 12 9 9 2
18 9 0 9 13 3 2 13 9 9 2 9 1 0 12 1 12 9 2
28 0 7 0 9 2 9 7 0 9 4 13 3 1 0 9 2 14 12 5 2 7 0 9 2 12 5 2 2
7 9 13 3 1 0 9 2
32 1 0 9 4 13 12 9 9 1 9 9 1 9 0 9 7 0 9 2 13 11 11 2 3 0 9 11 2 1 9 2 2
24 9 9 2 15 13 1 0 9 1 11 1 11 7 4 13 1 12 9 2 13 3 1 9 2
13 3 3 15 7 0 9 13 1 11 1 0 9 2
9 4 13 3 1 11 7 0 11 2
8 3 15 13 7 1 0 9 2
41 9 2 0 9 11 2 2 12 2 9 11 2 9 12 2 11 11 2 0 2 11 2 11 9 12 11 12 9 12 2 9 2 2 2 12 12 2 12 12 12 2
13 9 9 9 1 9 10 9 1 9 9 7 9 2
6 9 9 13 12 9 2
29 10 9 13 1 15 0 9 9 12 2 12 2 12 2 12 2 0 9 11 12 2 0 12 2 0 9 12 12 2
22 1 9 13 3 9 1 9 10 9 2 9 0 9 9 9 7 9 1 0 9 2 2
16 13 13 3 1 9 1 0 9 9 1 0 12 2 11 12 2
13 9 13 16 0 12 2 3 12 9 1 0 9 2
21 9 1 0 9 13 0 1 0 9 3 1 0 9 2 7 15 1 9 12 5 2
45 12 9 13 11 11 2 9 2 12 2 12 12 12 2 12 12 12 2 12 12 12 2 12 12 12 2 12 12 12 2 12 12 12 9 12 2 9 2 2 12 2 12 12 12 2
4 13 13 7 13
5 9 13 0 9 2
6 13 9 9 9 7 9
8 13 4 3 3 2 0 13 2
22 3 13 11 11 2 9 1 11 2 0 9 1 9 2 16 15 13 0 9 9 12 2
24 10 9 13 1 9 9 11 11 2 11 11 2 11 11 7 9 9 2 0 0 9 1 11 2
9 1 0 9 9 15 13 7 9 2
2 11 11
9 11 11 13 1 9 9 0 9 2
11 3 13 1 9 9 10 9 2 3 9 2
9 10 9 2 15 13 1 11 9 2
15 1 15 13 9 0 9 2 16 15 13 9 0 1 9 2
10 1 9 13 1 9 1 11 2 11 2
11 1 9 2 7 13 15 1 15 1 9 2
10 13 0 9 0 7 13 1 0 9 2
6 3 15 13 9 9 2
11 13 15 1 15 9 2 13 13 1 9 2
9 1 9 12 15 13 7 13 13 2
10 13 2 16 14 3 13 13 10 9 2
12 2 16 4 15 13 0 2 13 1 15 2 2
9 1 0 9 15 13 9 7 9 2
10 13 0 2 16 9 15 3 3 13 2
6 9 4 13 15 9 2
12 3 1 9 4 3 13 0 9 9 1 9 2
9 12 0 9 2 13 2 9 9 2
9 2 3 0 13 9 1 0 9 2
7 13 4 3 2 15 13 2
6 13 4 10 0 9 2
10 13 4 9 9 2 15 4 15 13 2
10 13 4 13 9 2 16 15 13 9 2
7 13 7 0 2 13 4 2
14 9 13 14 9 2 9 1 9 1 9 7 0 9 2
21 3 13 9 2 15 13 3 3 12 9 0 9 3 2 13 12 9 1 9 11 2
6 3 13 3 9 9 2
6 3 2 9 13 9 2
9 2 7 0 9 1 9 1 11 2
4 15 13 0 2
10 13 4 15 3 2 16 3 15 13 2
6 10 0 9 4 13 2
13 3 0 9 1 9 9 2 3 13 0 3 13 2
14 7 9 2 3 15 13 1 9 2 15 13 3 0 2
9 3 15 15 13 13 1 0 9 2
5 3 4 3 13 2
11 13 4 1 9 0 9 2 3 1 9 2
15 13 15 9 2 16 16 15 13 9 7 1 9 13 9 2
7 9 13 0 7 3 0 2
6 9 13 0 0 9 2
8 2 3 3 1 15 2 2 2
6 3 3 13 9 13 2
15 7 13 0 7 7 9 13 0 2 16 4 13 0 9 2
13 1 9 13 0 13 15 9 7 3 1 9 13 2
11 10 9 13 0 13 2 4 0 3 13 2
18 7 13 13 3 1 12 2 13 0 13 0 9 7 1 0 15 13 2
5 2 3 15 13 2
8 13 4 2 13 2 16 9 2
12 9 13 1 9 2 15 15 12 9 1 15 2
16 3 4 13 13 7 3 13 1 0 9 2 15 4 15 13 2
11 7 13 4 9 13 7 13 3 13 0 2
6 2 16 0 9 13 2
10 1 9 13 1 0 7 13 1 9 2
6 3 13 1 9 3 2
15 9 13 1 12 0 9 9 2 9 2 9 2 1 0 2
11 3 4 3 13 0 9 2 13 4 15 2
9 15 15 13 1 9 2 1 9 2
8 2 9 13 3 3 10 9 2
10 9 13 9 1 12 7 12 9 3 2
12 3 13 0 9 2 16 4 13 0 9 1 2
6 10 9 1 0 9 2
8 13 13 12 3 2 3 3 2
10 1 9 11 7 11 13 9 10 9 2
5 3 13 9 3 2
9 7 1 0 9 2 16 15 13 2
8 13 0 9 7 9 13 0 2
7 2 1 15 13 9 13 2
8 13 1 9 9 9 1 9 2
14 13 9 2 16 3 13 0 9 2 0 3 7 3 2
9 9 4 13 13 0 9 2 9 2
8 0 9 0 9 2 0 9 2
8 15 13 9 1 9 0 9 2
11 0 9 13 15 2 0 9 4 13 9 2
10 9 13 13 0 9 7 1 15 9 2
7 2 10 9 15 13 0 2
12 9 9 3 13 2 9 15 13 1 9 9 2
26 14 3 1 15 13 0 2 7 15 1 10 9 13 1 9 0 9 2 1 0 9 2 1 0 9 2
4 9 15 13 2
12 13 14 13 2 15 13 1 10 3 0 9 2
5 9 9 13 3 2
17 7 7 0 9 2 1 15 13 9 2 4 13 14 12 0 9 2
13 0 9 12 7 12 9 9 0 7 1 9 0 2
11 3 13 2 15 9 13 2 7 3 13 2
12 1 9 13 7 1 9 2 15 13 0 9 2
11 2 3 13 2 3 13 10 9 1 9 2
7 1 9 0 9 0 9 2
9 14 1 9 2 7 1 0 9 2
7 9 13 0 1 12 9 2
5 9 13 13 9 2
9 13 15 15 3 9 1 9 9 2
5 2 3 0 9 2
8 13 15 2 16 1 15 13 2
22 0 10 9 15 13 13 7 13 1 9 1 11 2 15 4 13 1 9 1 9 9 2
7 2 1 0 9 13 9 2
5 13 15 13 15 2
14 3 2 3 15 9 0 13 1 12 2 13 1 0 2
10 12 9 1 9 9 13 9 1 9 2
2 3 2
7 2 15 15 3 14 13 2
2 3 2
15 1 10 9 15 13 1 0 9 9 2 9 7 9 9 2
6 9 4 13 0 9 2
9 13 9 1 11 7 13 3 3 2
5 13 15 1 9 2
16 13 15 1 9 2 9 2 9 2 9 2 9 2 9 9 2
5 13 1 10 9 2
9 1 9 13 7 9 1 9 9 2
7 15 13 10 0 0 9 2
5 9 13 14 9 2
8 13 9 2 16 1 9 13 2
5 2 7 9 0 2
20 16 15 1 11 13 1 0 9 2 3 4 13 7 13 2 16 0 14 13 2
4 9 15 13 2
12 13 15 0 9 2 7 0 9 3 1 9 2
8 13 15 15 2 3 0 9 2
40 9 2 9 11 2 12 2 9 12 2 12 12 11 12 2 9 2 9 2 2 12 2 12 12 12 2 9 0 9 1 11 12 2 9 2 2 2 12 2 12
7 9 2 9 11 1 11 2
7 9 3 13 0 9 9 2
4 7 3 13 2
2 9 2
8 9 13 3 0 9 2 7 0
2 9 9
1 12
18 0 9 1 9 9 2 15 13 13 9 2 13 13 9 1 0 9 2
10 0 9 1 0 0 9 3 4 13 2
13 10 9 13 10 9 1 10 0 9 1 9 12 2
25 13 9 9 9 1 9 0 9 9 9 1 0 9 2 16 9 4 13 1 10 9 13 12 9 2
4 2 0 9 2
4 13 15 9 2
6 13 2 15 3 13 2
10 13 15 15 2 16 0 9 13 3 2
8 13 15 0 10 9 0 9 2
9 13 3 1 15 13 9 0 9 2
7 10 9 13 1 10 9 2
3 9 7 9
29 13 4 2 16 9 0 9 13 9 13 9 1 0 9 2 15 13 10 9 1 0 9 7 13 15 1 15 9 2
18 13 15 15 0 2 16 1 0 0 9 3 9 9 13 13 0 9 2
4 11 11 2 11
4 13 15 0 2
14 16 15 13 1 15 0 2 13 13 0 9 12 9 2
2 11 11
27 9 2 9 2 9 2 0 9 2 0 12 2 12 12 11 12 2 9 2 2 2 12 2 12 12 12 2
2 10 9
6 3 3 15 13 1 9
8 2 9 9 2 12 2 12 2
48 9 0 9 0 9 1 0 9 4 1 9 0 9 3 13 0 9 2 16 3 1 11 2 7 15 9 0 0 9 2 12 9 2 7 9 0 9 1 9 2 12 5 12 5 12 9 2 2
42 0 9 2 13 2 14 0 9 2 3 11 12 9 3 2 3 12 9 3 2 13 0 0 9 2 7 2 1 0 9 2 15 4 1 15 3 13 14 12 9 3 2
15 1 15 15 1 0 9 0 9 1 11 13 0 9 9 2
40 16 4 13 0 9 2 16 4 13 9 0 9 1 11 2 0 2 1 9 9 1 9 7 1 9 2 2 4 0 9 13 3 0 12 2 7 3 12 9 2
4 11 11 2 11
18 9 9 2 0 9 13 2 3 13 0 1 9 13 3 0 9 9 2
15 9 4 13 1 0 0 9 7 13 4 1 15 0 9 2
9 15 3 10 9 13 1 0 9 2
4 1 9 0 9
8 2 9 9 2 12 2 12 2
11 9 1 0 9 4 15 13 1 0 9 2
4 7 9 9 2
17 9 9 7 9 1 9 13 13 9 2 15 13 9 1 0 9 2
29 1 0 0 9 2 7 13 15 13 15 0 2 9 3 1 9 7 9 13 9 1 15 9 2 9 7 9 9 2
8 0 9 13 1 9 3 13 2
15 7 9 2 15 0 9 13 2 15 13 1 9 9 13 2
16 13 0 13 2 3 15 3 1 15 9 13 1 0 0 9 2
4 11 11 2 11
4 0 9 1 9
8 2 9 9 2 12 2 12 2
12 13 15 9 2 3 10 9 13 10 9 9 2
18 3 1 9 9 2 7 16 15 13 2 16 3 9 3 13 16 13 2
13 7 15 13 0 2 16 15 4 13 1 15 13 2
24 1 0 9 1 10 9 2 1 9 2 7 9 1 0 9 2 3 13 0 9 1 0 9 2
19 0 9 3 13 2 10 9 13 1 0 9 3 9 10 9 1 0 9 2
17 14 15 1 15 13 9 0 9 2 3 3 9 2 3 3 9 2
19 13 9 9 2 7 13 15 2 15 13 15 2 15 13 15 0 9 9 2
27 7 1 0 9 13 1 15 3 9 10 2 16 0 0 9 13 10 9 3 1 9 0 1 0 9 9 2
8 13 15 13 9 1 10 9 2
4 11 11 2 11
2 0 9
8 2 9 9 2 12 2 12 2
14 16 0 9 13 0 9 0 9 7 0 9 0 9 2
24 9 13 13 9 1 10 9 7 3 13 10 9 3 2 7 14 13 3 7 13 9 0 9 2
10 9 0 9 15 0 9 3 13 13 2
24 7 16 4 13 2 3 1 9 0 2 9 0 9 2 13 13 2 3 7 10 9 13 3 2
42 3 13 0 9 2 15 13 3 1 9 1 9 2 7 0 9 13 13 1 9 9 3 2 16 3 13 2 3 3 7 10 9 4 13 0 9 1 0 9 1 9 2
19 3 4 9 9 7 9 9 9 2 3 7 1 9 0 9 9 2 13 2
22 7 10 9 15 13 1 9 2 3 13 13 1 9 9 9 2 7 9 9 1 9 2
21 16 13 9 1 9 3 0 2 3 13 0 13 9 1 9 2 7 3 13 9 2
9 0 9 9 15 3 9 3 13 2
20 13 15 2 16 0 9 4 1 0 9 10 9 13 13 9 1 9 3 0 2
16 1 15 2 15 13 3 1 9 2 13 0 9 1 9 0 2
21 1 0 9 13 7 0 0 9 2 7 16 4 15 13 16 9 1 9 10 9 2
11 3 0 13 13 7 9 9 11 7 11 2
5 11 11 2 0 11
5 9 13 9 7 9
8 2 9 9 2 12 2 12 2
23 13 3 10 0 0 9 1 9 2 3 13 9 3 0 2 16 1 9 7 13 0 9 2
16 13 4 7 9 2 16 9 1 9 1 9 1 9 13 13 2
9 3 1 15 1 9 3 13 0 2
12 13 3 0 2 7 3 15 15 1 15 13 2
14 13 2 16 1 0 9 13 3 2 7 16 13 3 2
4 11 11 2 11
6 12 15 13 2 0 14
11 0 9 1 11 7 11 9 1 9 11 2
10 12 13 9 1 9 2 0 1 0 9
10 9 11 13 0 9 11 16 0 9 2
29 1 0 9 0 2 11 13 1 11 3 0 9 9 16 1 11 2 15 15 3 13 1 0 9 9 1 0 9 2
2 11 11
23 16 15 9 3 13 1 0 9 9 0 9 14 1 12 0 9 2 0 13 12 0 9 2
19 1 0 9 13 9 1 11 2 15 9 0 9 13 0 9 2 3 0 2
3 11 1 11
18 9 9 2 15 15 0 9 13 1 0 9 2 13 0 9 0 9 2
20 0 9 9 10 0 9 3 13 1 11 2 3 13 0 9 7 0 0 9 2
17 11 13 0 9 2 9 2 0 9 2 9 0 9 9 3 13 2
17 1 11 15 13 0 0 9 2 15 13 0 9 11 7 0 9 2
12 1 11 13 3 9 11 3 0 16 1 9 2
10 3 15 3 13 1 9 9 7 9 2
25 3 13 9 2 3 13 11 13 1 9 1 11 1 9 2 16 3 13 0 9 0 1 0 11 2
17 1 11 2 15 13 9 11 12 2 9 2 3 13 1 12 11 2
20 0 1 15 4 13 9 11 11 2 15 3 10 9 13 16 2 0 9 2 2
4 0 7 0 9
36 0 9 13 1 9 1 0 9 1 3 0 9 9 2 0 0 9 1 9 7 9 1 12 5 1 0 0 9 1 0 9 9 1 0 9 2
18 13 15 15 13 12 5 9 9 1 11 9 1 11 7 0 0 9 2
22 1 0 9 9 13 3 9 0 9 11 1 9 14 12 9 9 3 2 13 0 9 2
16 11 13 0 9 2 16 4 13 0 9 1 9 13 1 11 2
7 9 4 13 0 9 11 2
20 9 11 15 13 9 9 1 11 1 12 9 9 1 9 12 1 12 9 3 2
15 1 9 0 9 7 0 9 0 9 3 3 13 0 9 2
12 13 1 15 3 9 1 9 0 9 0 9 2
29 0 9 3 0 9 1 0 9 13 0 9 2 3 9 9 13 12 5 2 13 15 0 9 2 3 13 0 9 2
19 15 3 13 0 9 2 9 9 1 9 15 13 2 13 9 0 2 11 2
16 0 9 11 13 9 9 2 9 2 0 0 9 2 9 3 2
8 0 9 4 13 0 9 11 2
8 7 9 0 9 13 1 11 2
3 9 1 9
9 0 9 0 9 13 7 0 9 2
9 0 9 9 13 9 1 0 9 2
19 13 9 1 0 7 0 9 2 1 9 7 9 2 1 0 9 7 9 2
17 3 2 16 13 9 3 3 0 2 3 13 2 16 13 0 9 2
6 3 13 9 0 9 2
24 0 9 1 9 13 1 9 3 12 9 9 2 16 1 0 9 13 15 9 2 13 0 9 2
31 0 9 13 3 9 2 15 15 13 0 9 7 9 2 15 4 3 13 9 2 3 1 0 1 15 13 9 3 0 9 2
23 3 0 9 13 3 11 2 3 13 9 13 12 5 7 9 9 13 12 7 12 0 9 2
10 1 9 1 11 3 3 13 0 9 2
13 16 0 15 13 9 1 0 9 7 0 0 9 2
13 12 9 13 1 9 0 9 13 1 0 0 9 2
3 15 13 2
9 1 0 9 1 9 11 13 11 2
13 1 0 9 7 0 9 13 0 7 1 12 9 2
17 15 1 15 13 3 13 10 0 7 0 9 15 13 1 9 11 2
22 9 0 9 3 13 2 16 15 1 0 0 0 9 1 11 13 3 0 9 1 11 2
14 1 0 9 1 11 3 15 13 16 1 2 9 2 2
12 3 11 7 11 3 13 2 16 9 13 0 2
8 13 15 7 1 0 0 9 2
24 1 11 3 13 13 1 0 9 9 1 0 9 2 7 12 9 15 12 3 13 1 0 11 2
4 9 1 9 2
17 1 9 13 15 16 1 9 2 12 13 2 1 0 13 0 9 2
4 2 0 9 2
4 9 11 1 9
14 1 9 7 9 9 0 0 0 9 15 13 0 9 2
16 3 9 11 2 15 9 13 9 7 13 15 9 7 0 9 2
14 3 15 0 9 3 10 9 13 1 9 3 0 9 2
2 11 11
35 0 10 9 13 13 9 7 9 2 16 10 9 13 0 2 13 15 2 3 7 1 15 13 13 2 13 11 11 2 9 0 0 9 11 2
2 0 9
27 1 0 9 9 13 0 9 2 0 9 0 9 2 15 13 13 1 0 9 1 9 7 13 0 2 9 2
6 0 9 13 0 9 2
30 0 0 9 13 13 10 9 7 9 1 9 2 15 4 13 1 12 9 2 9 2 9 2 9 2 1 12 9 9 2
24 0 9 9 1 9 13 13 15 0 9 2 1 15 15 13 9 9 1 0 0 7 0 9 2
32 1 9 1 0 9 0 2 11 11 13 3 9 9 1 10 9 1 9 11 12 9 1 11 1 9 0 2 0 7 0 9 2
14 10 9 3 13 9 1 9 1 11 2 11 7 11 2
31 9 13 9 9 13 15 0 0 9 2 13 10 9 9 0 9 1 11 7 0 0 11 11 2 0 9 1 9 9 2 2
14 1 9 1 10 9 13 13 1 11 0 9 7 9 2
2 9 0
12 0 9 1 9 13 0 1 2 11 9 9 2
18 13 0 1 9 9 1 9 2 9 2 7 7 1 9 9 1 9 2
14 0 9 9 13 9 1 9 0 2 0 2 7 0 2
18 9 13 1 9 1 9 9 7 9 2 15 13 9 1 3 0 9 2
53 13 2 14 15 2 13 3 1 9 9 11 2 0 11 2 2 11 2 11 2 7 11 2 11 2 2 15 13 9 10 12 9 2 15 1 9 13 0 9 2 7 13 0 13 10 9 7 9 10 9 7 9 2
34 9 1 11 13 7 1 9 11 7 13 9 9 1 9 9 1 9 9 2 13 9 9 7 13 0 13 0 9 1 9 10 0 9 2
4 9 13 1 9
11 1 9 0 9 2 0 9 13 3 0 9
20 12 1 9 0 9 11 4 0 1 9 0 0 9 1 0 9 1 0 9 2
21 1 0 9 4 1 9 1 10 9 3 13 1 9 2 15 13 9 1 9 9 2
17 0 13 7 0 9 2 16 0 9 13 0 9 2 15 13 10 9
30 1 9 9 1 10 9 15 13 1 9 0 9 2 3 4 13 9 13 15 1 9 9 2 15 15 13 13 10 9 2
3 9 1 9
12 13 1 15 9 0 7 0 2 7 7 0 2
9 3 0 9 7 13 2 9 2 2
48 13 15 1 9 2 15 1 0 9 13 9 7 9 7 1 9 15 15 13 9 2 15 3 3 13 0 9 2 15 11 13 3 0 2 0 2 0 2 2 2 2 7 3 3 0 2 0 2
25 13 15 1 9 2 16 15 15 13 14 9 2 15 13 15 13 2 7 13 3 2 13 15 13 2
12 13 3 1 9 2 16 9 13 9 1 9 2
24 7 3 15 3 3 3 13 3 0 9 1 9 2 13 0 9 7 3 3 13 15 7 15 2
33 1 0 9 2 1 9 2 1 0 9 1 9 9 2 15 4 13 4 3 13 13 0 9 2 15 15 15 1 9 0 9 13 2
5 7 3 13 3 2
13 3 3 0 2 0 7 0 13 9 1 10 9 2
20 15 0 13 10 9 1 9 2 15 4 13 13 2 15 0 13 10 0 9 2
12 7 9 3 0 2 7 3 4 15 3 13 2
5 7 3 9 13 2
6 13 3 2 7 3 2
3 0 13 3
11 1 9 7 13 13 0 2 3 0 9 2
10 10 9 1 15 1 0 9 3 13 2
10 13 9 9 2 9 7 0 0 9 2
29 13 15 13 2 16 0 9 2 0 10 9 2 13 10 9 1 9 9 7 3 2 15 13 0 2 1 0 9 2
25 3 3 0 9 15 13 2 16 10 9 13 3 0 2 3 0 13 9 2 15 1 15 4 13 2
29 16 15 13 2 15 13 9 1 9 9 2 13 2 16 3 16 0 0 13 9 0 9 2 9 9 7 0 9 2
23 13 15 7 13 2 16 3 0 9 0 9 13 0 9 1 9 9 2 1 15 4 13 2
40 13 15 2 16 0 9 3 13 0 9 2 15 4 13 13 2 7 13 15 1 9 10 0 9 2 1 0 9 9 7 1 9 2 15 4 1 15 13 13 2
13 13 13 9 0 9 7 13 9 1 9 9 0 2
21 0 9 15 3 3 13 13 1 0 9 1 9 0 9 2 16 13 2 16 13 2
11 1 9 15 13 7 9 1 0 9 9 2
31 13 15 7 9 2 3 9 0 1 0 0 9 0 1 11 2 1 3 0 9 2 13 0 13 1 0 2 0 0 9 2
7 7 15 1 3 0 9 2
17 9 13 3 9 0 2 3 0 0 9 2 15 1 0 9 13 2
2 11 11
35 9 2 11 2 0 2 9 2 2 1 9 12 2 12 12 11 12 2 9 2 2 2 12 2 12 12 2 9 2 2 12 2 12 12 2
4 9 1 9 2
16 14 13 13 2 9 1 0 9 13 13 3 2 16 0 9 2
3 3 1 9
15 0 9 9 11 13 1 12 2 12 2 1 12 2 12 2
22 0 9 1 0 0 9 1 11 15 3 3 13 7 1 0 9 0 2 0 0 9 2
39 9 9 11 11 1 10 9 12 2 9 3 13 2 16 9 1 0 0 7 0 9 4 0 0 9 13 3 1 12 2 9 2 7 3 1 12 2 9 2
52 0 9 0 9 2 15 9 13 0 9 11 11 13 9 0 9 1 9 2 3 13 9 0 0 9 2 7 7 13 0 9 2 7 15 9 0 0 2 0 9 0 2 0 9 1 9 2 9 7 0 9 2
5 7 9 0 9 2
12 1 12 2 9 13 11 13 1 9 0 9 2
54 9 9 9 11 2 15 15 9 0 9 1 9 3 13 2 13 0 2 1 0 9 13 13 3 0 0 9 2 3 4 12 9 3 13 9 0 1 12 2 9 12 2 16 4 13 4 0 0 7 0 9 13 9 2
31 1 10 9 7 9 9 11 11 13 2 15 13 9 3 1 9 9 0 9 2 15 4 15 10 9 13 13 7 10 9 2
30 9 2 15 13 13 1 11 0 1 15 3 2 16 0 9 0 9 13 1 9 0 9 1 0 0 0 7 0 9 2
20 0 9 7 9 15 15 3 13 9 1 3 0 9 7 9 9 1 0 9 2
2 11 11
4 9 2 9 9
5 11 2 11 2 11
1 11
27 0 2 11 2 12 2 12 2 0 7 0 9 9 0 9 2 11 2 12 2 2 12 2 12 2 12 2
42 13 11 9 11 9 2 12 12 11 2 11 12 2 9 2 2 2 12 2 12 12 2 12 12 2 12 12 2 12 2 9 2 2 12 2 12 12 2 9 2 12 2
15 9 2 11 2 12 2 12 2 2 12 2 12 2 12 2
41 13 11 11 2 12 12 11 2 0 12 2 9 2 2 2 12 2 12 12 2 12 12 2 12 2 12 12 2 9 2 2 12 2 12 12 2 9 2 12 12 2
21 11 2 9 0 0 9 2 11 2 9 11 2 12 2 2 12 2 12 2 12 2
41 13 11 11 2 0 2 9 2 2 12 12 11 2 1 11 12 2 9 2 2 2 12 2 12 2 12 12 2 12 2 9 2 2 12 2 12 12 2 12 12 2
28 11 2 0 9 9 2 9 2 9 2 9 7 0 9 0 9 2 11 2 12 2 2 12 2 12 2 12 2
6 13 11 11 2 11 2
20 11 2 12 2 0 3 0 9 2 11 2 12 2 2 12 2 12 2 12 2
47 13 9 2 0 2 9 2 2 12 12 11 2 11 11 12 2 12 2 9 2 2 2 12 2 12 2 12 2 12 12 2 12 2 9 2 2 12 2 12 12 2 9 2 12 2 12 2
20 9 2 9 7 9 1 9 7 9 2 11 12 2 2 12 2 12 2 12 2
5 13 11 2 11 2
1 11
1 11
16 11 2 0 9 0 9 2 12 2 2 12 2 12 2 12 2
19 11 2 9 9 7 0 9 2 11 2 12 2 2 12 2 12 2 12 2
20 9 2 0 9 9 2 9 7 0 9 2 12 2 2 12 2 12 2 12 2
16 11 2 0 9 0 9 2 12 2 2 12 2 12 2 12 2
17 0 0 9 2 12 2 9 2 12 2 2 12 2 12 2 12 2
18 11 2 0 9 0 9 7 9 2 12 2 2 12 2 12 2 12 2
12 9 9 2 12 2 2 12 2 12 2 12 2
31 9 1 11 13 0 11 0 2 0 12 2 12 2 12 11 2 9 2 2 2 12 2 12 2 9 2 12 9 0 2 11
16 9 11 2 0 9 9 2 12 2 2 12 2 12 2 12 2
15 11 2 0 9 9 2 12 2 2 12 2 12 2 12 2
18 11 2 9 2 0 9 0 9 2 12 2 2 12 2 12 2 12 2
22 11 2 9 0 9 2 0 2 0 7 0 9 2 12 2 2 12 2 12 2 12 2
32 9 2 11 2 9 2 9 2 0 2 2 0 12 2 12 12 11 2 0 9 2 9 2 2 9 2 2 12 2 12 12 2
1 11
26 11 2 0 0 9 9 9 2 9 2 9 7 0 9 2 11 2 12 2 2 12 2 12 2 12 2
18 11 2 0 9 1 9 2 11 2 12 2 2 12 2 12 2 12 2
22 11 2 0 9 9 9 2 9 2 9 2 11 2 12 2 2 12 2 12 2 12 2
21 11 2 12 2 0 0 9 2 11 2 12 2 12 2 2 12 2 12 2 12 2
35 9 1 11 13 11 2 0 2 9 2 9 12 2 9 2 12 11 2 9 2 2 2 12 2 12 12 2 9 2 2 12 2 12 12 2
1 9
3 1 0 9
53 0 9 9 12 1 0 9 1 11 2 15 3 13 1 15 2 16 9 0 9 15 3 3 13 2 7 15 1 12 2 9 0 9 2 3 1 0 9 4 13 1 9 2 1 9 13 0 9 9 1 9 9 2
26 1 10 9 15 9 13 13 0 9 9 9 1 0 9 7 14 9 9 9 9 3 0 1 0 9 2
4 1 9 13 9
8 9 9 9 2 0 9 13 9
41 9 1 9 0 7 3 0 9 2 15 13 9 9 9 11 2 13 9 9 9 9 0 7 0 9 9 0 7 0 9 2 9 2 1 9 13 15 1 0 9 2
27 3 1 0 9 0 9 1 9 4 15 13 0 9 9 9 11 11 11 2 15 13 10 9 1 0 9 2
26 2 13 15 2 16 9 9 0 7 0 9 4 13 0 13 3 1 12 2 9 12 2 3 15 13 2
18 7 16 9 1 10 9 13 2 13 15 13 2 16 9 13 0 9 2
16 1 0 9 9 13 0 0 9 0 9 0 1 9 0 9 2
4 3 13 13 2
25 3 9 1 9 1 9 12 13 12 9 7 1 9 12 13 1 12 9 2 3 13 15 12 9 2
10 3 13 1 0 9 0 1 0 9 2
13 2 9 3 13 9 13 3 9 2 3 7 9 2
5 13 13 0 9 2
10 0 9 9 0 9 13 0 0 9 2
13 13 3 13 9 3 2 16 4 0 9 13 0 2
8 9 13 3 13 1 0 9 2
10 0 0 9 13 1 15 3 16 9 2
15 3 3 13 0 13 2 3 1 9 1 9 0 9 13 2
19 13 3 1 9 7 9 9 1 9 1 9 2 15 13 10 9 12 9 2
11 16 0 9 7 9 13 0 3 1 9 2
6 13 3 7 0 9 2
13 1 0 9 4 9 7 0 9 13 13 0 9 2
16 0 9 13 1 9 7 9 7 7 13 13 3 1 0 9 2
20 14 16 15 13 2 16 10 9 15 13 15 9 2 13 0 1 15 13 13 2
32 2 7 16 15 15 4 3 13 0 9 9 2 9 3 13 13 1 0 2 9 9 2 1 0 7 0 9 9 1 0 9 2
7 15 4 15 13 1 9 2
5 13 1 0 9 2
5 0 9 13 0 2
29 13 7 0 13 3 3 2 16 15 4 13 0 9 1 9 0 9 1 15 2 16 9 0 9 4 13 0 9 2
31 1 9 9 0 12 0 9 2 0 9 9 0 2 13 0 9 2 16 9 9 4 13 13 0 9 9 9 1 0 9 2
14 9 16 15 4 15 13 3 13 2 3 1 12 9 2
12 3 15 15 7 13 1 9 9 2 13 9 2
14 16 4 9 13 2 13 4 9 0 9 9 1 9 2
15 7 13 0 3 13 2 10 9 4 1 9 9 13 13 2
19 7 1 9 1 0 9 13 2 16 13 3 13 0 9 10 9 1 9 2
29 2 9 1 0 13 13 0 9 1 0 9 1 15 9 0 9 2 3 14 1 15 2 15 13 10 9 1 9 2
11 15 4 13 0 0 9 1 9 2 13 2
11 13 15 2 16 4 15 4 13 0 9 2
19 0 0 9 13 1 9 0 9 2 1 15 15 13 9 1 9 1 9 2
27 16 4 1 15 13 15 9 0 0 9 2 1 9 1 15 4 15 13 13 0 0 9 1 10 9 9 2
15 15 0 4 13 13 1 10 9 1 9 3 12 9 9 2
19 2 0 9 2 15 9 13 2 3 13 3 1 9 1 10 9 0 9 2
8 4 9 13 1 10 0 9 2
2 14 2
10 1 0 9 4 13 9 0 9 9 2
8 15 13 9 0 9 0 9 2
18 13 2 16 3 13 3 1 9 2 3 0 0 9 1 9 9 13 2
16 0 9 13 4 2 7 10 9 13 1 0 0 9 16 9 2
18 13 15 3 0 16 0 9 2 7 13 13 3 2 16 1 15 13 2
12 13 4 2 16 0 9 9 9 13 0 9 2
19 10 9 1 0 9 13 1 15 2 3 3 15 4 10 9 1 9 13 2
15 13 4 3 0 1 0 9 7 9 3 3 13 0 9 2
6 0 9 13 1 9 2
11 13 1 9 0 9 9 9 11 11 11 2
14 0 9 9 4 1 10 9 9 0 7 0 9 13 2
5 1 10 9 13 2
2 9 12
1 9
6 9 1 9 7 0 9
9 1 9 12 4 13 0 0 9 2
11 3 1 15 15 13 7 0 9 1 9 2
15 15 13 9 13 10 9 9 7 13 3 10 9 9 3 2
42 1 3 0 9 13 7 1 0 9 2 15 13 3 9 9 9 1 9 9 9 2 9 1 9 1 9 2 9 9 7 9 9 9 9 0 15 9 9 2 0 9 2
25 13 9 9 1 9 13 15 1 10 9 13 9 9 1 9 7 0 9 2 15 13 0 9 11 2
43 1 9 0 9 13 0 9 9 1 9 1 9 1 9 7 9 0 9 9 2 12 2 12 9 2 2 16 9 7 9 4 13 0 9 2 2 13 3 9 9 0 9 2
23 9 2 9 11 2 0 12 2 12 12 11 2 9 2 5 9 2 2 12 2 12 12 2
3 9 0 9
32 0 0 9 7 1 15 0 9 9 15 13 1 0 9 9 0 9 2 3 15 13 7 0 9 1 0 3 9 1 0 9 2
18 11 11 2 9 9 9 0 9 2 15 10 9 13 13 1 0 9 2
7 13 9 7 9 0 9 2
34 9 10 9 13 3 3 3 1 9 2 9 0 9 0 9 13 0 9 1 0 9 2 1 9 1 9 7 9 2 0 15 0 9 2
17 3 3 13 9 9 0 9 7 0 9 13 1 9 3 3 3 2
18 1 0 9 15 0 9 3 13 11 13 7 13 15 3 9 2 2 2
12 0 9 7 9 13 13 13 15 3 16 11 2
13 7 3 3 13 1 9 9 10 0 9 2 2 2
31 0 9 1 0 9 13 3 3 13 11 2 13 3 0 9 10 0 9 2 7 3 2 3 13 2 2 13 10 9 2 2
17 3 13 13 0 9 1 9 1 15 0 1 15 2 16 4 13 2
13 9 2 0 11 2 0 12 2 12 12 11 12 2
4 13 9 9 13
7 9 0 9 13 9 16 0
15 13 9 2 16 0 13 10 9 2 15 0 13 1 9 2
23 3 3 13 13 0 9 1 9 2 15 13 0 3 2 16 3 13 0 9 3 0 9 2
35 1 15 2 3 3 0 0 9 2 15 13 9 9 2 9 1 9 9 3 13 13 15 1 0 9 2 4 13 1 10 0 9 11 11 2
2 11 11
8 2 13 1 15 12 9 9 2
17 1 0 13 2 1 0 2 0 1 0 9 9 2 3 7 13 2
21 16 0 7 0 13 9 9 2 13 15 2 16 15 4 15 13 1 0 9 9 2
3 13 15 2
20 1 10 9 13 13 0 9 2 7 1 0 9 9 3 10 9 3 13 13 2
11 1 15 4 13 7 0 2 16 0 9 2
11 2 3 1 0 9 2 15 3 3 13 2
14 15 13 0 9 2 15 15 13 13 2 7 14 3 2
35 13 1 9 2 16 4 13 2 10 9 7 9 13 0 2 7 1 15 15 1 15 7 13 2 15 1 15 13 10 0 9 1 12 9 2
21 3 1 15 13 0 9 2 7 1 0 9 9 13 1 2 7 3 9 7 9 2
19 2 16 13 3 9 0 9 0 2 3 0 9 13 3 1 0 0 9 2
13 10 0 0 9 9 13 3 0 7 1 0 9 2
24 9 13 7 1 10 9 14 1 12 9 2 13 1 9 9 12 2 12 2 9 2 9 2 2
22 1 0 7 0 9 9 3 13 2 16 13 9 0 0 9 7 3 13 10 0 9 2
13 2 13 4 13 2 16 9 13 7 13 3 0 2
14 1 9 0 9 3 13 9 13 10 9 13 3 3 2
9 7 0 9 9 2 0 0 9 2
15 9 3 13 1 15 2 16 14 2 7 14 2 7 3 2
21 2 15 3 13 2 16 9 2 1 15 13 9 9 7 9 2 9 0 9 13 2
27 13 3 15 9 2 7 12 13 0 2 3 3 13 0 9 2 0 9 7 0 0 9 1 9 1 9 2
20 3 15 3 13 2 13 1 9 0 9 2 15 4 3 13 1 9 0 9 2
18 0 9 0 9 3 7 13 16 9 0 9 7 15 0 9 3 13 2
7 7 9 13 9 7 3 2
18 2 1 9 9 13 13 0 9 1 0 9 7 0 11 7 0 11 2
22 0 9 13 3 3 0 2 3 3 1 9 2 7 3 13 2 7 13 3 7 3 2
12 9 13 3 1 15 2 16 4 13 10 9 2
8 9 13 3 0 0 9 9 2
8 15 16 9 2 9 2 2 2
32 2 2 2 2 1 15 7 13 0 9 1 11 2 11 2 11 2 11 2 11 2 7 10 0 11 2 13 15 3 1 11 2
38 7 15 13 9 9 9 1 0 9 2 7 16 13 1 11 2 9 13 9 1 12 0 9 2 15 13 9 7 13 2 15 4 13 0 15 3 13 2
25 2 15 3 13 1 9 2 16 15 1 9 10 9 13 9 9 7 1 0 9 2 3 1 9 2
16 0 9 9 9 1 9 13 9 10 9 2 3 1 0 9 2
8 0 7 13 9 0 9 13 2
8 7 3 1 15 15 9 13 2
37 2 13 3 2 16 16 15 13 2 16 14 9 0 9 15 13 1 0 9 2 3 9 9 9 1 3 0 9 13 1 0 9 0 9 0 9 2
14 3 2 3 13 0 7 0 9 2 13 7 10 9 2
6 7 9 13 3 0 2
33 16 15 13 3 0 9 9 2 3 13 0 9 9 2 9 9 0 0 9 7 0 0 9 2 15 9 14 13 2 3 9 9 2
23 2 3 1 9 0 9 2 16 13 0 0 0 9 0 9 13 2 4 13 3 0 9 2
23 1 0 7 3 0 9 15 13 13 2 7 3 15 13 13 2 15 15 13 1 9 9 2
17 16 4 13 7 0 9 2 3 3 9 13 7 4 13 15 13 2
12 0 9 15 9 3 13 7 14 15 15 13 2
21 2 15 13 9 2 15 10 9 13 14 3 13 9 0 0 7 0 9 2 2 2
17 2 2 2 7 3 15 1 15 13 9 0 9 9 9 2 2 2
14 2 2 2 2 7 9 7 3 13 3 1 9 9 2
42 3 13 0 13 12 9 2 9 10 9 2 15 13 0 9 2 7 7 3 13 9 0 9 0 9 2 7 3 9 0 9 2 3 3 3 13 3 9 1 0 9 2
7 2 4 3 13 0 9 2
18 13 7 3 0 9 9 1 0 9 13 1 9 1 9 2 0 11 2
12 13 1 9 2 15 13 9 1 9 0 9 2
39 10 9 15 14 13 9 0 9 7 13 9 1 0 9 2 7 3 13 0 9 2 16 1 9 9 15 13 4 13 9 1 9 2 16 9 0 0 9 2
6 2 3 13 9 9 2
13 1 9 2 14 0 7 0 2 7 1 0 9 2
59 13 2 16 9 1 9 13 1 0 9 13 0 15 0 2 16 0 9 9 9 2 3 15 2 16 15 13 9 13 15 3 9 7 9 1 10 0 9 2 3 13 0 9 3 2 16 4 9 7 9 9 9 7 9 13 1 0 9 2
12 2 15 3 13 9 1 9 1 0 9 13 2
17 13 15 3 10 9 10 9 2 16 13 0 0 9 7 9 9 2
22 1 15 15 9 4 13 13 2 13 9 2 16 13 0 3 13 1 0 9 9 9 2
21 16 15 3 13 16 9 1 9 9 7 9 9 9 9 2 13 15 1 10 9 2
2 9 2
11 9 3 13 9 9 1 9 1 0 9 9
4 13 1 0 9
11 3 1 12 0 9 13 0 9 0 9 2
9 13 15 1 9 1 10 0 9 2
7 0 9 13 12 2 9 2
17 13 15 1 0 9 0 9 2 0 9 0 2 0 7 0 9 2
15 0 9 0 12 2 12 2 4 1 0 13 9 12 9 2
4 9 2 0 9
2 9 3
22 1 9 0 9 2 0 1 10 9 2 4 1 0 9 9 7 9 13 3 15 3 2
18 0 0 9 0 9 1 11 1 0 9 9 7 9 0 1 9 9 2
16 0 9 1 9 11 7 0 9 9 13 1 0 9 0 9 2
19 1 9 0 9 2 9 2 9 2 3 13 0 9 16 10 0 0 9 2
14 0 9 2 3 9 2 13 0 13 3 1 0 9 2
21 9 1 9 12 9 13 9 1 9 10 12 2 9 3 1 9 9 9 7 9 2
6 9 13 3 12 9 2
13 9 2 15 4 13 1 9 2 13 1 12 9 2
12 1 9 1 9 13 1 10 9 7 9 9 2
17 9 0 9 7 1 0 9 7 9 13 3 10 2 10 2 9 2
8 0 0 9 13 3 9 11 2
9 13 15 2 16 4 13 7 0 2
4 11 11 2 9
14 0 9 0 1 10 9 13 1 0 9 7 0 9 2
11 4 3 12 3 13 1 9 1 12 9 2
26 13 14 9 2 15 4 13 1 10 0 9 2 7 7 15 2 1 15 15 9 2 9 13 16 9 2
3 13 10 9
8 11 15 13 1 0 7 0 9
27 16 4 1 9 9 9 2 12 2 12 13 9 0 9 2 13 4 15 1 9 9 9 7 0 0 9 2
20 9 1 9 9 7 9 1 10 9 9 9 3 1 3 0 9 13 9 11 2
22 1 10 9 3 10 3 0 9 13 2 3 1 9 9 11 13 3 12 1 0 9 2
2 11 11
40 1 9 2 3 4 15 13 0 9 9 11 2 9 2 3 15 3 13 13 0 9 2 16 3 0 9 2 3 13 0 2 13 11 11 2 12 1 9 9 2
11 13 4 2 16 15 4 13 1 0 9 2
17 1 9 1 9 1 9 9 7 9 15 7 10 0 0 9 13 2
12 9 1 0 9 0 9 1 15 3 3 13 2
16 7 4 15 1 0 9 13 13 3 7 1 0 7 0 9 2
9 13 15 0 9 2 7 13 9 2
2 9 9
21 11 15 13 2 16 3 3 13 3 0 7 0 9 2 15 1 9 13 10 9 2
26 3 1 15 13 0 9 11 11 2 15 15 13 3 0 9 2 0 9 1 0 9 2 3 0 9 2
19 0 9 9 13 10 9 0 9 2 16 4 9 13 13 3 0 9 9 2
20 16 13 15 1 9 2 10 9 13 11 15 2 7 13 10 9 1 0 9 2
17 1 15 13 3 1 9 3 0 9 2 15 13 1 9 9 9 2
45 10 9 13 0 7 0 9 2 15 3 13 9 2 7 3 13 0 13 1 0 9 1 0 9 9 2 10 9 7 9 2 13 9 9 0 9 2 7 13 9 1 9 0 9 2
17 10 9 0 0 0 2 9 2 4 13 9 0 9 16 9 9 2
11 3 1 9 9 1 0 9 13 3 3 2
9 13 3 7 9 1 9 0 9 2
3 3 1 9
17 3 3 13 9 13 2 16 1 9 13 3 10 0 7 0 9 2
20 9 0 9 7 0 9 13 3 16 14 9 1 0 9 2 9 1 0 9 2
14 0 9 1 9 0 9 13 9 7 0 7 0 9 2
10 0 9 3 13 2 3 15 13 9 2
9 9 13 1 9 0 9 3 13 2
13 3 0 9 13 9 2 3 3 3 13 10 9 2
12 15 13 9 2 0 15 1 9 9 0 9 2
9 0 3 13 1 9 9 0 9 2
13 13 1 0 13 7 13 9 9 9 7 10 9 2
28 16 4 9 1 9 13 1 9 2 13 1 0 9 9 1 9 11 13 9 9 1 10 9 0 9 1 9 2
4 13 2 15 13
31 0 9 13 2 16 9 15 13 9 1 0 9 7 13 15 2 16 15 13 13 7 1 0 9 2 1 15 3 3 13 2
15 3 13 1 9 9 9 2 3 15 1 10 9 13 13 2
22 3 13 13 9 9 0 9 3 2 7 3 14 0 9 9 1 0 9 3 0 9 2
9 0 13 15 3 1 0 9 11 2
13 9 15 15 13 3 1 0 0 9 2 15 13 2
27 9 7 13 13 3 0 9 0 7 3 0 9 2 13 3 0 0 9 1 9 7 10 9 1 9 9 2
15 13 13 9 9 9 1 0 9 2 13 3 0 0 9 2
16 1 9 13 11 0 9 2 7 15 3 2 7 7 1 9 2
21 1 0 0 9 2 15 15 13 1 10 9 9 2 13 11 3 0 9 7 9 2
10 13 15 3 1 9 7 9 2 9 2
12 3 15 9 1 10 9 9 9 12 3 13 2
15 0 9 12 9 15 7 13 9 2 15 4 3 13 13 2
22 11 11 15 13 2 16 3 4 13 1 10 9 2 9 13 2 15 3 9 3 13 2
39 9 2 11 2 9 2 9 2 0 2 2 0 12 2 12 12 11 12 2 9 2 2 12 2 12 2 12 2 12 2 12 2 9 2 2 12 2 12 2
2 9 2
3 1 9 2
3 3 14 2
4 1 10 9 2
5 1 0 3 14 2
3 1 9 2
5 15 1 10 9 2
3 9 1 9
10 3 3 3 3 9 13 1 9 10 9
1 9
19 0 9 1 11 4 13 13 0 1 0 9 2 1 15 13 10 0 9 2
17 0 9 15 13 0 9 2 15 13 0 9 0 9 1 0 9 2
10 16 3 0 9 13 13 9 9 9 2
8 10 9 16 10 15 13 13 2
17 13 15 7 0 9 2 15 13 9 0 0 9 2 0 12 9 2
17 13 0 7 1 9 0 9 2 15 13 13 0 9 1 0 9 2
12 11 11 2 11 2 9 9 7 9 2 11 9
9 1 9 7 1 9 2 3 1 9
27 1 9 4 13 1 9 10 0 9 2 3 4 13 13 0 9 2 16 4 13 3 3 7 13 3 3 2
63 1 9 9 4 13 2 15 4 13 13 3 1 9 2 16 4 15 13 13 1 9 2 16 4 4 3 1 9 0 9 13 1 0 0 9 7 3 16 15 4 13 1 9 0 9 13 0 9 9 1 3 0 9 16 4 15 13 9 1 9 0 9 2
45 9 4 13 13 15 1 0 0 2 0 9 2 1 15 4 13 0 0 9 2 9 0 9 7 9 9 9 9 7 13 4 4 3 1 9 0 9 7 0 9 1 0 0 9 2
6 1 9 15 13 9 2
14 1 9 11 11 2 9 9 9 9 1 0 9 13 2
33 9 1 9 4 1 9 13 2 7 1 9 9 0 0 9 13 0 9 2 16 0 13 1 0 0 9 0 0 9 7 3 9 2
22 1 9 9 15 1 0 9 4 15 0 0 13 13 9 1 0 9 1 9 12 5 2
18 1 9 9 13 3 13 0 9 2 10 9 13 0 1 9 9 9 2
13 1 0 9 4 13 3 12 5 7 3 12 5 2
32 13 2 14 3 10 9 1 9 12 9 2 4 1 9 13 1 9 9 1 9 12 2 12 9 7 1 9 1 9 12 9 2
9 12 10 9 15 13 1 0 9 2
13 1 9 4 13 2 9 1 9 15 1 9 13 2
4 1 0 9 2
29 1 9 4 13 3 1 9 9 2 3 1 0 9 2 1 15 4 13 10 9 2 16 4 15 13 1 9 13 2
26 1 9 4 15 14 1 9 1 0 9 1 11 13 2 9 15 1 9 1 9 9 13 3 1 9 2
27 9 9 0 7 0 9 15 13 2 16 10 9 4 13 1 15 2 15 13 0 9 2 16 10 9 13 2
11 13 15 1 10 9 2 0 9 4 13 2
11 9 1 0 9 1 9 0 9 3 13 2
50 10 9 2 15 4 13 0 9 1 12 9 1 0 9 12 9 1 0 9 12 9 2 4 15 13 3 13 1 0 12 9 1 12 9 3 2 3 4 15 4 13 7 1 9 1 0 9 1 12 2
14 3 4 3 13 1 9 2 1 0 9 2 12 9 2
16 9 9 15 3 13 2 16 4 13 9 1 9 9 9 9 2
12 9 0 9 9 13 9 1 9 0 0 9 2
13 3 13 13 2 14 3 15 9 13 3 0 9 2
17 1 9 0 9 15 1 10 9 13 16 0 13 15 1 9 11 2
1 11
3 1 0 9
16 9 11 1 9 9 0 9 2 15 4 13 1 0 0 9 2
18 9 13 12 9 7 1 12 9 1 3 0 9 2 15 4 13 9 2
14 0 9 7 0 9 9 9 13 1 9 3 1 9 2
11 1 9 9 0 9 13 9 7 9 0 2
30 9 2 11 2 0 2 9 2 2 0 12 2 12 12 11 2 9 2 2 2 12 2 12 2 9 2 2 12 2 12
31 9 11 9 11 2 7 11 11 2 15 13 12 0 0 9 0 9 11 7 0 0 9 1 9 3 3 16 12 9 9 2
25 9 4 3 3 3 13 1 9 2 16 4 13 3 13 1 9 7 9 9 1 9 10 0 9 2
34 9 2 11 11 2 0 2 9 2 2 0 12 2 12 12 11 12 2 9 2 2 2 12 2 12 12 2 9 2 2 12 2 12 12
21 9 11 9 2 15 13 1 0 9 13 9 0 9 9 0 9 2 0 9 9 2
17 15 13 9 12 0 9 2 15 4 13 3 0 12 9 1 11 2
11 0 9 13 12 9 2 0 12 9 9 2
20 9 13 3 0 14 1 9 11 2 7 3 15 13 7 1 0 9 1 11 2
39 9 2 11 9 2 0 2 9 2 2 9 0 9 2 1 9 12 2 12 12 11 12 2 9 2 2 2 12 2 12 12 2 9 2 2 12 2 12 12
4 9 7 9 2
4 9 7 9 9
13 9 9 0 9 13 3 1 9 2 15 13 3 2
33 0 9 3 13 2 16 10 0 9 13 9 7 15 7 0 9 9 7 9 0 9 9 2 1 15 3 13 9 1 9 7 9 2
17 7 4 13 9 13 0 9 1 10 0 9 2 3 1 0 9 2
2 11 11
12 13 15 3 3 2 1 15 15 13 9 13 2
19 13 15 14 1 0 9 9 2 7 7 1 0 9 1 0 7 0 9 2
22 1 15 2 15 9 3 13 2 4 3 13 1 11 11 1 11 2 15 13 1 9 2
34 16 13 1 10 9 1 15 0 9 2 1 12 9 9 15 15 13 13 9 2 16 1 10 9 1 15 13 2 15 13 3 3 12 2
24 13 15 3 2 16 1 10 9 3 10 9 2 3 15 16 10 9 13 1 9 7 9 15 2
5 1 9 10 7 0
5 3 13 1 9 2
13 13 15 14 15 12 9 2 15 13 1 10 9 2
23 1 9 0 9 2 9 2 0 9 2 9 2 9 7 9 2 13 3 7 1 0 9 2
16 15 3 3 13 1 9 9 2 7 7 10 9 3 13 9 2
26 0 13 7 15 2 3 9 13 7 3 1 9 9 1 9 2 15 13 0 9 7 1 9 0 9 2
8 13 4 15 13 7 0 9 2
23 7 15 1 10 9 11 0 13 2 10 9 1 0 9 10 9 15 13 9 2 3 9 2
4 0 13 12 9
33 1 10 0 9 1 11 15 13 1 15 2 16 1 0 9 13 9 1 9 1 9 3 0 2 3 7 1 9 12 7 12 9 2
28 13 15 2 16 1 15 4 15 13 13 1 9 9 1 10 9 2 7 13 9 1 12 9 4 13 3 0 2
24 16 1 12 0 9 13 9 11 11 12 9 2 3 1 12 0 9 4 15 13 1 12 9 2
17 13 4 13 3 7 9 0 7 0 9 2 3 7 9 0 9 2
17 9 10 9 4 3 13 1 0 0 9 2 7 15 13 1 0 2
16 13 15 2 16 9 4 13 13 1 9 3 1 12 1 15 2
12 9 4 15 15 13 13 0 9 7 3 9 2
3 9 1 9
23 16 9 13 0 9 7 9 3 2 13 15 15 1 9 0 7 9 10 9 9 9 11 2
10 9 13 3 12 9 9 1 0 9 2
25 1 9 15 9 0 7 0 9 13 9 0 7 0 9 2 9 2 1 9 13 15 1 0 9 2
13 1 9 15 1 15 13 13 9 0 7 0 9 2
4 9 1 9 2
17 9 16 9 2 1 12 9 13 1 0 7 1 0 1 0 9 2
18 1 15 3 15 12 3 13 2 13 4 3 13 14 1 12 1 15 2
7 13 1 9 12 7 12 2
6 1 0 9 15 3 13
5 9 2 9 2 9
10 13 15 0 7 0 9 1 0 9 2
8 15 13 9 7 15 13 9 2
6 10 13 1 15 9 2
24 3 15 13 2 16 0 9 13 13 9 9 7 9 2 16 0 9 7 9 9 15 3 13 2
24 1 0 9 13 9 1 10 9 7 9 7 3 13 1 9 3 0 7 0 2 1 0 9 2
17 13 9 9 2 9 2 9 2 9 2 0 9 9 7 9 9 2
9 3 15 13 2 16 13 1 9 2
11 13 9 9 2 9 2 0 9 2 9 2
21 3 3 13 13 2 7 1 9 9 13 1 9 2 16 7 10 9 13 13 9 2
18 13 9 9 2 9 1 0 0 9 2 9 2 9 1 0 9 9 2
26 9 15 13 2 16 1 10 9 3 13 1 9 2 7 9 2 15 13 13 16 9 7 0 9 9 2
13 15 15 13 2 15 13 1 9 1 9 7 9 2
22 13 15 13 0 9 2 15 4 1 0 9 1 3 0 9 13 1 0 9 0 9 2
8 2 9 9 13 3 3 0 2
10 13 15 9 1 9 0 2 0 9 2
33 9 13 9 16 9 2 9 2 9 2 7 1 9 9 0 9 13 0 13 2 16 9 9 13 9 13 9 9 7 3 13 9 2
18 2 13 13 0 15 9 2 15 13 13 2 13 7 3 13 1 9 2
13 10 9 13 1 9 9 9 1 0 7 0 9 2
20 2 9 0 9 13 0 3 13 3 9 7 3 13 0 2 7 3 0 9 2
13 2 13 4 13 1 9 9 10 9 7 9 9 2
9 7 13 0 13 0 9 7 9 2
13 3 0 9 13 1 10 9 0 9 1 10 9 2
22 7 10 9 15 4 13 13 9 1 9 9 1 10 9 1 10 9 2 9 2 9 2
10 16 2 13 2 15 13 15 0 9 2
2 11 11
6 9 2 14 2 13 9
9 0 9 7 0 9 2 12 2 2
17 9 0 9 13 0 9 7 13 9 1 9 0 0 9 7 9 2
23 10 9 3 13 4 13 7 9 2 15 9 1 15 13 3 1 0 9 2 9 7 9 2
6 3 13 3 3 0 2
30 0 9 0 11 13 3 1 9 12 9 2 1 15 11 2 11 13 9 9 2 15 13 0 9 1 9 9 1 9 2
33 10 3 0 9 13 13 1 9 1 9 2 16 1 9 12 15 1 15 7 1 9 13 9 9 0 15 3 9 0 9 0 9 2
13 15 13 9 13 15 1 9 9 2 9 7 9 2
18 7 13 0 13 15 1 10 9 7 3 3 3 13 0 9 0 9 2
19 1 0 9 13 9 2 1 15 13 9 13 9 1 9 13 1 12 9 2
2 0 9
14 13 15 0 2 3 0 2 7 13 0 1 15 13 2
15 2 9 7 9 0 9 2 0 9 0 9 1 0 9 2
11 2 9 2 15 3 13 0 9 0 9 2
9 2 9 9 7 9 1 0 9 2
4 2 0 9 2
10 2 9 2 9 7 9 0 0 9 2
5 2 9 9 9 2
9 2 9 0 9 2 0 7 9 2
2 0 9
22 1 15 4 15 13 13 16 4 15 13 2 15 13 1 9 9 1 15 7 10 9 2
5 1 15 3 13 2
21 12 2 9 1 9 0 9 0 1 9 2 16 15 3 0 9 13 13 0 9 2
12 12 2 0 9 1 9 0 9 1 0 9 2
14 12 2 3 0 9 1 9 9 2 9 0 9 3 2
24 12 2 0 9 9 9 9 1 0 9 10 9 2 16 0 9 13 13 1 10 9 0 9 2
20 12 2 0 9 1 0 9 0 1 9 9 1 9 9 1 15 1 10 9 2
9 12 2 9 0 9 1 9 9 2
13 12 2 9 9 0 9 1 9 13 1 15 9 2
8 12 2 0 9 0 9 9 2
11 12 2 9 9 2 7 0 9 0 9 2
17 12 2 9 9 2 7 10 9 2 1 9 7 0 9 0 9 2
10 12 2 0 9 7 0 9 1 9 2
13 12 2 9 9 2 9 2 9 3 2 1 9 2
9 12 2 9 7 0 0 9 9 2
3 15 13 9
18 10 0 9 1 0 9 13 13 0 9 9 1 9 0 9 0 9 2
19 1 12 0 9 4 13 0 9 9 0 9 2 15 13 13 9 0 9 2
13 1 10 9 15 3 0 9 9 13 1 0 9 2
28 16 1 15 13 2 16 13 9 2 13 15 1 0 9 0 9 0 15 9 2 15 13 9 2 13 10 9 2
18 16 7 9 13 9 1 0 9 2 13 3 0 9 2 7 0 9 2
5 11 11 2 0 9
4 11 11 2 2
17 14 2 7 3 0 0 9 2 1 15 15 13 13 9 1 9 2
4 3 13 0 9
10 9 2 9 7 9 13 1 0 9 2
25 9 1 9 3 13 13 2 15 13 0 9 10 10 0 9 1 10 10 9 2 7 3 13 9 2
28 3 3 13 0 9 9 2 12 2 12 1 9 10 0 9 2 15 4 13 1 9 1 9 9 1 9 12 2
20 7 10 9 1 15 9 3 13 1 9 12 7 1 10 9 13 1 0 9 2
9 0 9 4 13 1 9 0 9 2
16 0 0 9 9 7 1 9 0 9 10 0 9 13 0 9 2
22 13 1 15 3 9 2 15 15 1 3 0 9 13 2 7 10 0 9 13 3 0 2
18 1 9 9 10 9 15 13 3 13 0 9 2 15 13 9 7 9 2
13 1 9 0 9 13 9 9 9 3 1 9 12 2
21 10 9 13 4 13 1 0 9 0 1 0 11 2 15 15 7 9 9 3 13 2
24 16 4 3 13 1 9 9 9 2 13 0 9 11 9 0 9 0 9 1 9 0 9 9 2
13 15 15 13 3 13 9 0 9 0 9 1 9 2
24 16 13 7 0 9 9 1 0 9 0 2 13 3 3 0 13 0 9 1 15 9 1 9 2
19 3 15 13 2 16 9 9 1 0 9 11 13 0 16 9 0 1 11 2
20 1 9 11 13 3 9 9 2 16 4 13 1 9 13 2 1 15 13 13 2
15 15 15 13 13 15 9 9 2 15 13 0 9 0 9 2
14 10 9 9 2 7 9 9 2 7 3 13 13 9 2
24 1 10 9 4 15 13 13 1 9 1 9 9 2 15 15 7 13 13 3 16 1 12 9 2
20 16 4 15 13 0 9 13 3 2 4 13 3 14 16 0 9 9 0 9 2
12 7 3 15 13 2 16 9 1 0 9 13 2
7 3 1 0 9 13 9 2
22 13 15 3 12 9 0 9 2 15 3 1 9 12 13 1 0 9 1 0 9 9 2
32 3 3 3 13 10 9 1 10 0 9 2 16 15 1 9 0 9 11 11 11 13 2 16 3 10 9 13 9 9 2 2 2
13 9 2 0 9 3 13 7 0 15 3 13 13 2
2 11 11
3 1 9 2
7 13 9 0 9 1 9 2
17 3 15 13 2 16 15 15 1 15 1 9 13 13 9 0 9 2
3 1 0 9
4 9 0 13 2
2 3 2
26 9 13 3 0 9 2 16 13 2 9 13 0 9 2 7 3 3 0 0 0 9 2 4 13 9 2
19 13 2 14 13 0 9 13 15 0 9 7 3 13 0 9 0 9 9 2
3 9 9 2
12 13 15 3 1 0 10 0 9 2 13 9 2
5 7 3 2 2 2
22 1 9 0 2 7 7 0 9 9 1 10 0 9 13 2 16 13 10 0 9 13 2
4 13 0 9 2
7 13 15 10 9 3 0 2
18 3 16 1 3 14 2 7 1 9 0 3 13 0 9 9 0 9 2
22 15 13 1 10 9 9 7 10 9 0 2 15 15 13 1 9 12 7 12 9 12 2
7 11 10 9 1 0 9 2
15 3 13 13 9 2 15 13 1 0 2 0 9 0 9 2
6 0 9 2 9 7 15
3 9 1 9
18 1 9 4 13 9 9 2 7 15 1 15 13 3 7 1 10 9 2
6 13 4 15 7 3 2
18 15 15 7 13 0 9 2 15 15 12 13 2 15 15 1 9 13 2
12 13 15 9 13 3 7 13 13 9 1 9 2
4 11 11 2 11
31 1 9 12 0 9 15 9 13 13 9 9 2 16 15 0 13 1 15 7 1 9 10 9 3 2 16 15 13 0 9 2
27 1 9 1 10 9 4 15 0 9 13 13 10 9 7 13 3 0 9 1 9 0 9 2 15 13 9 2
14 1 10 9 4 4 10 9 1 9 9 1 9 13 2
35 10 9 7 13 3 1 9 2 16 4 3 10 9 2 13 2 2 15 13 2 16 0 9 13 3 10 0 9 7 13 9 0 9 9 2
35 1 9 2 16 0 9 13 1 0 9 9 2 3 1 10 9 1 15 7 10 9 13 2 7 12 13 3 0 9 1 9 1 10 9 2
5 2 9 2 1 9
25 1 0 0 9 4 13 0 13 15 1 9 9 2 16 1 9 9 4 4 13 7 9 13 13 2
7 3 15 13 1 9 13 2
13 3 2 16 13 1 9 2 13 0 9 1 9 2
29 15 15 3 13 1 9 7 0 9 2 16 3 4 13 7 13 1 9 13 10 9 2 1 15 13 3 9 0 2
4 13 15 13 2
4 11 11 2 11
20 9 9 13 1 0 9 9 3 13 0 9 1 9 0 9 2 13 9 12 2
28 3 4 7 10 9 13 9 9 13 9 3 1 12 9 0 9 0 9 1 9 7 9 1 9 3 12 9 2
8 10 9 15 13 1 0 9 2
27 16 15 3 0 9 1 9 13 0 9 9 2 13 15 13 1 10 9 0 9 3 0 7 0 9 0 2
12 0 0 9 4 15 7 13 1 9 10 9 2
27 13 1 15 2 16 4 13 2 3 1 0 9 7 0 9 2 3 1 9 1 9 0 9 7 0 9 2
2 9 9
12 13 9 1 0 9 2 3 3 13 0 9 2
24 3 13 12 0 7 0 9 7 13 1 15 2 16 1 9 1 15 0 9 13 1 9 9 2
7 15 1 15 7 9 13 2
17 13 9 2 16 13 13 0 9 2 16 4 13 13 14 0 9 2
6 4 13 13 0 9 2
4 11 11 2 11
11 13 15 2 16 4 10 0 9 3 13 2
48 1 0 0 9 2 15 4 1 15 0 9 13 2 7 1 15 4 15 13 9 9 2 4 13 3 3 13 2 16 1 9 2 16 7 9 13 9 13 2 13 3 1 9 1 9 0 9 2
33 13 0 2 16 9 13 0 13 2 16 3 9 13 3 3 7 1 0 9 7 9 1 15 0 9 13 1 10 9 3 10 9 2
2 9 9
28 1 0 0 9 4 15 13 1 15 2 16 9 1 10 9 15 13 13 3 3 2 16 12 9 2 0 9 2
26 9 9 4 7 4 13 2 16 10 9 10 9 3 1 9 13 9 2 16 4 13 0 0 0 9 2
5 13 9 9 9 2
4 11 11 2 11
35 1 1 15 2 16 13 3 0 9 2 15 15 13 1 9 2 0 9 2 7 9 4 13 1 15 0 9 2 13 15 15 0 9 13 2
11 9 0 1 3 0 9 4 13 0 9 2
14 0 9 13 0 9 9 2 11 11 2 11 1 11 2
23 9 2 11 2 1 9 9 12 2 12 12 11 1 11 2 9 2 2 2 12 2 12 2
2 9 9
11 3 13 3 9 2 3 13 0 15 13 2
28 1 9 0 9 13 9 2 3 13 10 9 2 10 9 15 13 2 3 13 1 0 9 2 7 1 0 9 2
20 0 9 2 1 15 0 9 2 1 0 9 14 3 13 9 2 13 3 3 2
3 15 13 2
9 9 13 1 10 9 9 1 9 2
24 1 10 9 2 15 15 13 1 9 1 12 2 9 2 13 0 9 2 9 7 0 9 9 2
14 9 1 10 9 13 12 2 9 1 9 12 10 9 2
3 9 0 9
3 9 13 9
8 9 15 3 13 0 9 0 9
19 1 10 9 15 13 0 9 0 9 2 15 13 1 12 2 9 0 9 2
14 1 9 9 2 0 9 1 9 2 13 12 0 9 2
27 9 4 13 14 1 3 0 9 9 9 2 7 13 7 0 9 2 15 1 9 0 9 13 1 10 9 2
32 1 10 12 0 9 1 9 0 9 7 12 9 2 9 2 13 1 15 9 0 9 1 10 9 2 15 15 3 13 0 9 2
2 0 9
20 0 0 9 13 9 0 9 1 0 9 2 9 0 9 7 9 0 0 9 2
21 9 1 0 0 9 7 9 13 0 9 13 1 9 2 15 13 0 9 7 9 2
18 13 15 0 9 2 3 13 0 9 2 9 7 3 13 9 0 9 2
10 0 9 15 3 3 13 1 0 9 2
13 9 7 13 7 0 9 1 9 0 7 0 9 2
15 9 0 9 15 3 13 9 2 15 13 0 1 0 9 2
8 3 15 13 7 9 0 9 2
7 0 9 13 9 7 9 2
11 0 9 9 15 13 9 7 9 0 9 2
21 3 15 13 13 9 0 9 1 0 9 2 3 1 9 9 2 9 2 0 9 2
24 1 0 9 15 13 0 9 0 9 9 0 0 9 2 3 1 9 2 9 7 0 9 2 2
2 9 9
41 3 13 1 9 9 0 9 2 3 1 0 9 2 9 9 9 2 3 0 9 0 9 2 9 9 0 9 1 9 2 9 0 9 9 7 3 0 9 1 9 2
16 1 12 2 9 4 13 3 12 0 9 1 9 12 9 9 2
36 1 9 0 9 13 1 9 0 1 9 0 9 3 2 0 9 2 10 0 0 9 2 0 9 11 2 11 2 11 2 15 0 9 3 2 2
15 10 9 7 4 3 13 7 3 4 13 14 0 9 9 2
17 13 3 1 11 2 11 2 0 9 2 0 9 11 2 11 11 2
29 1 9 0 9 13 1 12 2 9 9 0 15 9 9 2 9 2 9 2 0 9 2 9 2 9 7 0 9 2
3 9 0 9
32 1 9 0 0 9 2 3 2 9 7 9 2 13 0 9 2 15 9 0 9 9 7 0 9 0 9 13 0 9 1 9 2
14 9 13 4 13 1 3 0 9 7 9 1 0 9 2
11 13 13 9 0 9 7 1 12 2 9 2
15 0 0 9 9 0 9 1 9 15 13 1 9 12 9 2
24 9 0 9 13 1 9 9 0 9 12 9 2 15 13 1 12 5 3 16 9 9 15 9 2
10 3 4 13 9 14 1 9 9 12 2
13 1 10 9 13 0 0 9 9 9 1 12 9 2
5 11 11 2 11 11
32 9 2 0 0 9 2 11 12 2 12 12 11 12 2 9 2 2 2 12 2 12 12 2 9 2 2 12 2 12 12 12 2
3 0 9 9
24 1 9 12 1 9 9 9 13 9 9 9 1 0 0 9 2 15 13 1 12 2 9 12 2
42 1 9 13 2 16 1 9 1 12 2 12 2 12 13 9 11 11 1 9 9 1 9 0 9 9 7 13 13 1 9 9 7 1 15 3 9 1 9 12 5 9 2
35 10 9 4 13 7 1 9 12 2 9 2 12 9 7 1 9 12 9 9 2 12 2 12 9 2 2 1 9 1 9 1 9 0 9 2
15 1 9 2 16 15 9 13 0 9 2 13 15 1 9 2
3 9 3 9
10 9 1 3 16 12 9 13 9 7 9
13 0 9 3 13 3 7 3 3 16 1 12 9 2
15 13 3 1 9 7 13 2 16 4 15 13 3 1 9 2
13 10 9 15 3 13 1 10 0 9 7 11 11 2
18 9 3 13 1 9 9 2 15 15 3 1 10 9 7 9 7 13 2
2 11 11
11 13 1 9 2 3 0 9 13 12 9 2
17 13 1 0 9 2 16 9 1 0 0 9 1 11 13 3 9 2
2 13 9
20 16 9 1 9 13 1 9 10 2 0 0 9 13 14 1 10 0 9 3 2
15 9 9 13 3 3 3 0 16 3 2 13 11 2 11 2
7 1 9 15 15 3 13 2
3 13 0 2
14 0 2 15 1 9 13 13 2 13 0 9 1 9 2
29 16 13 13 2 16 9 15 13 3 3 7 9 9 13 0 9 2 3 14 13 0 9 1 9 9 1 0 9 2
11 13 15 15 7 0 9 7 9 1 9 2
3 9 1 9
13 1 10 9 13 3 0 2 16 9 13 2 13 2
11 13 14 10 9 7 9 2 15 9 13 2
6 3 0 15 7 13 2
18 1 0 9 9 13 0 9 9 1 9 9 2 9 9 7 9 9 2
11 3 13 0 9 2 9 2 9 2 9 2
11 15 13 0 9 2 3 12 12 15 9 2
6 15 13 1 0 9 2
12 9 1 9 1 0 9 1 11 2 11 13 2
22 9 13 0 9 2 7 16 14 15 3 2 2 13 0 15 13 1 0 7 0 9 2
14 13 7 0 9 9 2 7 3 15 1 0 9 13 2
6 9 13 3 3 0 2
9 9 13 7 1 9 9 1 9 2
18 3 4 13 9 3 2 7 1 0 0 9 0 9 2 16 15 13 2
8 7 15 4 15 3 13 9 2
18 16 13 9 0 1 9 7 0 9 2 13 0 9 1 0 9 0 2
23 0 0 9 1 0 9 9 1 9 9 13 9 2 15 15 1 0 9 13 14 12 9 2
11 9 9 13 1 9 11 2 11 1 9 2
16 3 13 9 1 0 9 1 0 9 2 14 1 10 9 3 2
25 9 13 3 0 2 7 1 0 9 0 9 15 13 9 0 2 9 2 2 15 3 13 16 9 2
22 3 15 13 9 1 9 2 3 1 9 13 3 12 9 2 7 1 9 9 15 13 2
9 1 9 13 13 7 1 0 9 2
8 9 1 9 13 3 0 9 2
8 0 9 13 3 0 2 0 2
17 0 7 0 3 3 2 7 3 0 9 15 13 1 9 7 9 2
11 1 9 13 9 0 2 3 1 9 9 2
11 0 9 13 9 9 7 13 3 1 9 2
7 1 9 9 13 0 9 2
15 9 13 1 9 2 3 13 9 3 2 13 1 0 9 2
3 13 15 3
6 9 13 1 9 3 2
12 15 13 9 2 15 15 11 2 11 3 13 2
12 15 2 15 3 13 2 15 13 0 9 13 2
15 9 2 15 3 13 9 14 3 2 13 3 9 2 13 2
17 13 15 0 9 2 1 15 13 9 7 1 9 2 7 1 9 2
11 1 9 0 9 3 13 7 9 9 9 2
11 9 15 1 15 0 9 13 1 12 9 2
18 1 0 9 1 9 3 9 13 1 12 9 2 1 9 9 12 9 2
18 3 13 3 9 9 7 9 2 7 3 3 9 15 13 9 7 13 2
5 15 13 3 0 2
25 11 11 13 2 16 9 15 3 13 3 2 16 4 13 14 10 12 9 2 7 3 3 0 9 2
23 7 3 10 0 9 13 2 16 4 15 9 13 1 9 3 2 16 13 1 15 9 13 2
18 15 7 13 9 15 2 9 13 3 0 7 9 3 13 7 3 13 2
15 9 2 9 9 2 11 11 2 0 12 2 12 12 11 12
4 9 1 9 2
15 3 15 13 2 3 0 9 13 7 1 0 9 15 0 2
1 9
12 1 9 9 15 13 9 9 13 1 0 9 2
9 9 9 1 9 9 12 1 9 12
4 9 9 9 9
1 11
1 11
7 11 2 0 0 2 9 2
2 0 11
1 11
1 11
1 11
7 11 2 0 9 2 9 2
2 9 2
9 0 9 2 9 2 0 9 2 9
7 9 2 9 2 9 2 9
5 9 12 2 12 2
30 11 12 2 9 9 2 0 0 11 2 9 12 2 12 2 0 9 9 7 9 2 12 2 2 12 2 12 2 12 2
39 13 11 2 9 2 9 2 0 2 2 0 9 2 12 12 11 12 2 11 12 2 9 2 2 2 12 2 12 12 2 9 2 2 12 2 12 2 12 2
46 11 2 9 0 9 2 9 12 2 12 2 9 0 7 0 9 1 9 7 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 12 2 2 12 2 12 2 12 2
43 13 9 11 2 9 2 9 2 0 2 2 12 12 11 2 0 9 2 11 12 2 9 2 2 2 12 2 12 12 2 12 2 9 2 2 9 2 2 12 2 12 12 2
44 9 2 9 2 9 7 9 12 2 0 0 9 0 9 2 9 9 2 0 9 2 9 1 9 9 2 9 7 9 1 9 7 0 9 2 12 2 2 12 2 12 2 12 2
45 13 11 2 0 2 9 2 2 9 9 7 9 2 12 12 11 12 2 9 12 2 9 12 2 9 2 2 2 12 2 12 12 2 9 2 2 12 2 12 12 2 9 2 12 2
5 9 12 2 12 2
50 9 2 11 2 11 2 11 1 11 2 11 2 9 11 2 2 11 2 11 2 0 11 2 11 2 9 2 11 2 9 1 11 2 11 2 0 2 11 2 11 1 11 2 11 1 11 2 0 9 2
22 0 9 2 11 2 9 9 2 2 11 12 2 11 2 9 11 2 1 12 9 2 2
25 0 9 2 11 2 9 11 1 12 9 2 2 11 2 9 2 9 1 11 2 1 12 9 2 2
5 9 12 2 12 2
20 11 2 9 2 11 2 0 9 0 9 2 12 2 2 12 2 12 2 12 2
49 13 0 9 7 9 2 0 2 9 2 2 12 12 11 12 2 9 12 2 0 2 9 2 9 12 2 9 2 2 2 12 2 12 12 2 9 2 2 12 2 12 12 2 12 12 2 12 12 2
28 11 2 9 2 11 2 0 9 9 2 0 9 2 9 1 9 7 9 2 12 2 2 12 2 12 2 12 2
6 13 0 9 7 9 2
26 11 2 9 2 11 2 0 9 9 1 9 2 9 7 0 9 2 12 2 2 12 2 12 2 12 2
6 13 0 9 7 9 2
35 11 2 9 2 9 2 0 9 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 12 2 2 12 2 12 2 12 2
6 13 0 9 7 9 2
27 11 2 9 2 9 2 11 2 0 9 0 9 2 9 7 0 9 2 12 2 2 12 2 12 2 12 2
6 13 0 9 7 9 2
21 11 2 9 2 0 11 2 0 0 9 9 2 12 2 2 12 2 12 2 12 2
6 13 0 9 7 9 2
37 9 2 0 11 2 11 2 11 2 9 11 2 11 2 11 2 11 2 0 9 2 2 11 1 11 2 11 2 9 1 9 2 2 9 1 11 2
16 0 9 2 9 2 9 2 9 2 0 12 2 1 12 2 2
5 9 12 2 12 2
31 11 12 2 0 9 1 9 2 9 0 9 2 12 2 12 2 12 2 12 2 9 12 2 12 2 12 1 12 9 2 2
29 13 0 9 9 2 12 12 2 11 12 2 0 12 2 9 2 2 2 12 2 12 2 9 2 2 12 2 12 2
14 9 2 0 9 2 11 2 9 2 2 11 1 11 2
17 0 9 2 11 12 2 0 9 2 1 0 9 9 1 0 9 2
5 9 12 2 12 2
41 11 12 2 9 2 11 2 11 12 2 0 9 0 9 7 9 2 0 9 7 0 0 7 0 9 0 9 9 9 7 9 2 12 2 2 12 2 12 2 12 2
46 13 11 2 0 2 9 2 2 12 12 11 12 2 11 2 9 2 9 2 2 9 2 2 12 2 12 2 12 12 2 9 2 2 2 12 2 12 12 2 9 2 2 12 2 12 2
31 11 12 2 9 2 9 9 12 2 0 9 2 0 9 2 0 9 2 0 9 2 2 12 2 2 12 2 12 2 12 2
31 13 9 9 1 0 9 2 11 11 2 11 2 12 12 11 12 2 11 2 0 12 2 9 2 2 2 12 2 12 12 2
10 9 2 11 2 11 1 11 2 11 2
18 0 9 2 11 12 2 11 2 11 2 1 11 2 1 12 9 2 2
2 9 2
10 9 2 11 2 11 2 11 2 11 2
2 9 9
15 9 0 9 13 4 13 15 9 9 2 3 7 0 9 2
19 1 0 9 13 13 7 9 0 9 13 3 0 9 2 3 9 9 9 2
9 1 15 13 1 0 9 0 9 2
7 12 2 10 9 15 13 2
17 12 2 3 3 15 13 2 16 9 9 1 9 13 9 10 9 2
7 15 13 0 9 10 9 2
16 12 2 1 9 7 9 13 7 3 0 13 1 10 9 13 2
6 1 15 13 9 9 2
6 15 13 1 9 9 2
19 12 2 13 13 2 13 13 15 7 0 7 13 10 9 7 9 1 15 2
8 1 15 13 13 13 9 9 2
5 10 9 9 13 2
38 12 2 16 4 9 9 3 13 7 13 1 10 9 13 2 13 3 13 15 2 16 3 3 16 1 15 2 3 7 1 10 9 13 9 13 0 9 2
4 15 15 13 2
6 9 1 9 0 9 2
19 12 2 0 9 13 13 9 2 9 7 9 2 15 13 0 1 0 9 2
20 0 13 3 13 10 0 2 3 2 0 9 2 15 4 13 9 7 9 9 2
4 12 2 14 2
8 0 9 13 0 9 0 9 2
9 12 2 9 9 13 9 0 9 2
14 12 2 0 9 13 2 16 2 4 13 9 0 9 2
8 9 0 9 4 13 3 3 2
5 0 9 13 0 2
7 1 0 9 4 13 0 2
4 13 0 9 2
13 12 2 3 0 9 4 13 1 9 1 9 9 2
51 9 2 11 2 0 0 9 2 11 9 2 9 2 9 2 0 2 2 0 2 9 2 9 2 0 9 2 12 2 12 12 11 12 2 9 2 2 2 12 2 12 12 2 9 2 2 12 2 12 12 2
6 9 1 9 9 11 2
19 9 2 9 2 9 2 13 9 0 2 3 3 0 2 3 0 0 9 2
5 9 7 9 5 9
6 9 15 13 1 9 2
4 0 9 13 9
7 9 9 7 9 3 13 2
11 15 2 15 13 13 2 3 13 0 9 2
13 13 9 7 1 15 13 3 2 15 15 13 13 2
14 13 3 9 2 16 9 13 14 15 2 15 3 13 2
12 3 1 9 0 9 15 13 0 9 0 11 2
2 11 11
15 9 11 11 2 1 9 2 13 9 3 1 9 1 11 2
7 9 3 13 1 12 9 2
10 13 9 2 9 9 7 0 0 9 2
2 0 9
18 1 9 9 13 9 3 3 2 16 13 9 2 1 15 15 13 13 2
5 9 9 13 0 2
7 0 1 9 13 13 9 2
11 1 15 13 13 14 14 13 7 0 9 2
10 13 15 9 0 9 7 3 0 9 2
33 13 15 3 1 15 2 16 4 0 9 13 9 2 15 13 1 9 2 0 9 1 9 2 9 0 9 3 2 0 0 9 9 2
14 1 12 1 9 9 13 2 16 9 0 9 15 13 2
17 16 9 13 9 1 0 9 13 2 13 15 3 7 13 0 9 2
6 13 9 13 1 9 2
10 3 2 1 9 13 3 16 9 9 2
6 13 4 3 10 9 2
15 0 9 13 3 3 13 9 2 15 15 13 7 13 4 2
16 9 9 13 7 13 1 15 9 9 9 7 0 9 2 9 2
4 1 9 15 13
14 1 0 9 2 15 9 13 2 13 0 9 9 9 2
7 13 15 1 0 0 9 2
13 3 0 11 13 9 13 1 12 7 12 5 9 2
19 15 0 9 2 15 3 13 9 9 3 2 16 13 0 9 13 0 9 2
24 3 3 13 9 1 9 9 2 9 15 3 13 1 0 9 1 9 9 9 7 9 0 9 2
11 10 9 13 14 0 9 2 13 9 11 2
16 1 0 9 15 13 0 9 2 0 1 12 7 12 9 3 2
6 3 15 9 3 13 2
15 3 0 9 13 0 9 1 9 9 2 10 9 13 9 2
21 3 15 13 1 9 1 0 9 2 1 9 12 15 13 9 1 0 9 1 9 2
12 13 9 2 13 9 2 7 1 9 1 9 2
5 9 13 3 0 2
2 0 9
14 3 0 13 13 1 9 9 2 13 9 1 0 9 2
9 9 15 1 0 9 13 7 13 2
5 0 15 13 13 2
9 0 9 13 1 11 14 12 9 2
34 1 11 15 13 9 2 15 13 9 1 12 9 2 3 9 2 15 13 1 12 12 0 9 9 2 2 3 0 9 2 15 13 9 2
9 1 10 9 13 13 14 0 9 2
7 0 11 13 3 9 0 2
12 9 3 13 2 16 13 1 0 9 9 9 2
4 11 15 13 2
14 15 0 9 13 0 2 16 15 13 1 15 0 9 2
15 16 0 11 13 13 0 9 2 3 13 0 9 1 9 2
24 9 13 7 9 0 9 1 0 9 7 1 9 9 2 1 15 13 9 13 7 1 0 9 2
16 15 13 0 1 9 9 1 9 0 9 2 3 13 9 9 2
20 1 15 2 16 4 15 13 9 9 2 10 0 9 3 13 2 13 9 11 2
12 0 11 3 13 9 13 0 9 3 1 9 2
17 0 9 3 15 13 2 7 9 15 1 9 9 13 1 0 9 2
12 0 11 13 10 9 1 0 9 0 9 9 2
1 9
9 13 0 12 13 2 16 3 13 2
4 9 1 9 2
7 9 0 9 13 13 0 2
13 1 9 9 1 12 9 15 0 11 13 1 0 2
6 1 0 9 15 3 13
12 9 1 9 7 0 9 4 15 13 13 0 9
15 9 0 7 0 9 13 1 9 9 1 9 7 0 9 2
35 9 7 9 3 13 2 16 15 13 14 1 9 9 9 2 7 7 1 0 9 9 9 2 15 4 1 15 13 13 0 9 1 0 9 2
9 3 4 13 13 1 9 1 9 2
3 13 11 11
34 1 0 9 4 9 0 9 13 12 9 2 9 1 9 1 0 9 2 7 9 1 0 9 9 2 7 9 1 9 1 0 0 9 2
25 7 16 15 1 0 9 13 10 9 3 13 2 13 0 15 3 13 1 12 7 13 15 0 9 2
11 13 1 9 9 1 9 2 15 9 13 2
21 1 9 10 0 9 3 13 1 9 2 15 13 13 1 0 9 3 1 12 9 2
44 13 3 1 9 14 9 9 2 7 7 9 7 9 15 1 9 2 3 9 9 1 9 7 9 9 2 13 0 9 9 9 11 11 11 2 15 4 13 1 9 9 10 9 2
2 9 9
10 9 3 13 13 9 0 9 7 9 2
25 13 15 2 16 9 4 13 13 9 1 15 2 16 9 1 10 9 13 13 1 9 10 0 9 2
31 3 4 15 12 0 9 9 2 7 2 1 0 9 2 0 9 2 1 9 7 1 9 2 13 12 9 1 0 9 9 2
12 1 0 9 15 13 2 3 4 15 14 13 2
10 9 9 1 10 9 13 12 9 3 2
13 1 15 13 9 3 12 9 2 15 15 15 13 2
8 9 1 15 13 12 9 3 2
11 9 13 12 9 7 0 9 13 12 9 2
8 0 9 13 13 9 12 9 2
18 1 9 4 13 9 0 9 12 9 7 3 13 9 1 9 12 9 2
5 3 15 15 13 2
3 9 9 2
1 3
2 1 9
3 0 9 12
4 9 2 9 12
3 0 9 12
4 0 9 12 12
2 0 9
15 9 3 13 3 3 13 0 9 1 9 9 7 0 9 2
9 0 4 15 13 13 1 0 9 2
13 13 4 15 13 9 1 10 0 9 2 3 9 2
20 0 9 4 15 13 3 1 15 2 16 4 15 1 0 9 13 0 0 9 2
20 3 13 7 9 9 1 9 1 9 0 0 9 7 3 0 0 7 0 9 2
22 13 4 15 13 9 9 2 16 4 15 3 9 3 13 1 9 9 2 9 7 9 2
16 1 9 1 0 9 13 0 7 0 9 0 9 1 0 9 2
23 3 2 16 15 3 0 9 13 3 0 0 9 2 4 15 13 1 0 9 2 13 2 2
10 13 4 15 0 0 9 1 0 9 2
21 3 7 0 9 1 9 1 9 9 9 2 7 9 3 3 0 2 13 11 11 2
4 9 12 9 3
24 1 9 3 0 9 1 9 9 1 9 0 9 13 9 9 0 9 2 1 15 15 13 9 2
29 1 9 0 9 2 15 13 15 0 16 9 9 2 4 13 13 7 3 0 9 9 2 7 2 15 1 15 2 2
18 3 15 13 13 2 16 3 1 9 1 12 9 3 15 9 13 4 2
14 3 4 15 9 0 9 13 1 0 9 7 1 9 2
20 9 13 1 15 2 16 1 9 1 9 1 0 9 13 0 0 9 0 9 2
2 9 9
21 1 0 0 9 4 15 3 1 12 2 12 2 12 13 9 0 9 1 0 9 2
26 9 1 10 9 13 1 0 9 0 9 2 7 1 15 2 16 4 9 1 0 9 13 9 0 9 2
15 0 9 1 9 0 9 4 15 13 13 1 9 9 9 2
20 3 4 13 4 13 0 2 9 0 9 1 9 2 9 7 0 1 0 9 2
14 13 1 15 0 16 1 9 2 16 15 13 16 9 2
8 1 0 9 9 13 9 9 2
5 13 15 9 9 2
10 13 15 2 15 13 9 1 0 9 2
15 1 9 0 9 4 15 13 1 0 9 9 12 9 9 2
17 15 4 15 13 3 13 1 9 9 7 3 1 0 7 1 9 2
17 1 15 10 0 0 9 4 15 13 15 13 7 9 2 7 9 2
17 1 0 0 7 2 0 2 9 4 15 13 13 0 9 7 9 2
11 9 3 13 2 7 16 14 1 9 9 2
16 0 9 13 7 3 2 0 2 9 13 1 9 9 1 9 2
2 9 9
37 7 16 15 15 0 9 9 0 7 0 9 2 9 2 4 3 13 2 9 3 13 7 0 9 0 9 1 0 7 0 9 1 9 1 0 9 2
5 15 13 12 9 2
16 3 13 2 16 4 13 1 0 9 9 1 9 1 0 9 2
19 0 1 9 13 2 16 13 3 9 1 9 10 9 1 0 1 0 9 2
22 3 9 9 9 9 1 0 9 13 1 9 9 2 3 1 2 9 2 9 1 9 2
3 0 9 9
16 1 9 1 9 13 1 9 9 0 13 1 0 9 9 9 2
13 1 0 9 13 1 12 9 7 0 1 12 9 2
20 2 0 9 2 1 9 3 12 9 4 13 13 9 1 9 12 7 12 9 2
16 3 4 13 13 1 0 9 1 0 9 1 0 9 10 9 2
26 0 9 13 7 9 9 9 9 9 1 0 0 0 9 7 0 9 9 13 0 9 0 9 1 9 2
18 9 0 0 9 3 13 9 2 16 4 15 0 9 13 1 15 9 2
17 1 0 9 9 0 1 9 13 1 9 9 11 10 3 0 9 2
15 9 13 1 0 9 9 2 7 7 13 13 14 0 9 2
4 9 1 9 2
13 3 15 15 3 3 13 2 9 7 9 3 13 2
19 16 4 3 1 15 13 9 1 0 7 0 9 2 13 4 15 13 3 2
4 13 15 0 9
8 0 9 9 9 11 3 13 9
21 1 0 9 13 0 2 9 2 9 9 1 12 9 9 9 11 2 9 1 11 2
19 16 7 9 1 9 13 2 13 15 1 0 0 9 1 9 3 0 9 2
2 11 11
10 1 9 9 11 15 7 13 0 9 2
18 9 11 3 13 3 0 0 9 2 15 15 3 1 10 9 3 13 2
30 1 9 0 0 9 1 9 12 2 15 3 13 1 12 0 9 0 9 7 0 9 2 15 1 9 13 0 0 9 2
2 0 9
9 1 12 9 13 0 9 13 9 2
15 7 15 9 13 1 9 14 1 9 2 7 7 1 9 2
18 9 13 1 11 9 1 9 2 13 0 9 1 11 2 11 7 3 2
9 1 0 9 15 1 15 13 9 2
20 13 9 2 16 1 9 13 9 1 9 0 9 0 0 2 0 7 0 9 2
18 1 0 9 13 12 9 9 9 9 11 2 9 13 13 1 0 9 2
24 0 9 9 11 11 13 0 0 9 2 13 4 12 0 9 2 15 4 13 0 9 1 9 2
3 1 0 9
19 0 9 9 9 9 11 13 2 1 15 7 9 2 3 15 9 13 9 2
6 3 13 12 0 9 2
30 1 0 0 9 13 9 1 9 9 12 7 12 9 2 7 3 13 7 9 1 0 9 2 14 16 4 9 13 9 2
11 16 4 13 1 9 2 13 9 7 9 2
17 1 9 13 9 1 12 9 9 7 9 9 2 13 11 2 11 2
10 1 9 12 13 9 10 9 1 12 2
24 13 15 3 13 9 1 9 2 3 4 13 1 9 2 0 2 9 2 15 3 2 15 3 2
9 3 3 13 0 9 1 9 9 2
18 13 15 2 16 13 9 14 12 2 12 9 9 2 7 3 7 0 2
5 3 15 13 3 2
17 3 4 9 9 13 14 1 9 9 2 16 1 10 9 9 13 2
19 3 15 9 13 14 12 7 12 9 2 7 15 13 3 16 12 0 9 2
5 0 13 9 9 2
11 9 13 1 0 9 2 1 9 7 9 2
15 13 15 14 9 9 1 3 0 9 2 7 7 9 9 2
15 0 9 15 3 1 0 9 13 9 1 12 9 9 3 2
13 13 2 14 9 9 1 12 2 13 9 10 9 2
2 13 9
11 1 9 9 9 13 0 9 1 10 9 2
11 13 9 0 9 13 9 2 16 13 0 2
10 13 15 2 16 7 0 9 3 13 2
20 7 15 9 4 13 14 9 9 2 7 7 0 9 2 3 0 9 1 9 2
5 7 3 13 9 2
15 13 4 15 13 0 9 2 0 9 3 12 9 0 9 2
18 13 13 3 15 2 16 4 13 0 9 7 9 2 13 11 2 11 2
29 9 7 13 3 1 9 0 9 2 9 7 9 1 0 9 7 13 13 7 16 0 9 2 15 13 0 0 9 2
15 9 1 9 2 12 1 9 9 13 9 0 9 1 11 2
5 3 13 10 9 2
2 9 9
14 11 13 1 12 9 3 1 12 0 9 1 12 9 9
2 9 2
15 9 2 15 2 13 2 3 9 0 9 2 7 3 9 2
24 3 1 0 9 2 3 9 0 1 10 9 13 3 0 9 2 15 15 13 1 2 9 2 2
22 3 3 2 10 9 13 1 9 7 9 0 9 1 15 13 3 1 9 9 1 9 2
2 11 11
25 1 9 0 9 9 13 2 16 1 9 0 9 2 9 7 9 13 9 3 0 1 9 9 9 2
45 16 1 15 13 9 0 0 9 1 9 2 9 2 1 9 7 9 2 3 13 2 16 1 9 0 9 2 3 1 9 10 9 9 1 9 15 1 0 9 7 9 13 9 9 2
3 0 9 9
8 0 9 3 13 3 9 9 2
10 3 15 7 3 13 2 7 3 13 2
44 7 3 13 2 16 3 1 0 9 7 9 1 9 12 13 13 9 2 9 9 7 9 2 2 10 9 13 1 9 12 13 12 9 1 0 9 2 7 15 13 3 14 9 2
29 1 9 15 13 7 0 2 9 2 2 1 15 13 2 1 9 9 2 1 9 12 1 9 1 9 9 10 9 2
33 10 9 4 7 3 13 2 16 1 9 13 3 13 9 2 16 1 12 9 0 9 13 11 1 12 9 0 0 9 7 0 9 2
14 7 16 9 10 9 13 2 9 10 0 9 3 13 2
42 13 1 15 1 0 9 2 16 1 12 9 0 9 13 9 12 9 2 12 9 2 12 9 2 12 9 2 12 9 2 12 9 2 12 9 2 12 9 7 12 9 2
5 0 9 2 9 2
37 1 9 9 0 9 11 13 0 9 0 9 0 0 9 2 15 13 9 1 9 7 4 13 1 0 9 2 15 13 0 0 9 7 0 0 9 2
22 0 9 13 9 2 16 13 1 9 2 16 9 13 1 0 9 1 9 12 1 12 2
6 0 9 15 13 9 2
17 0 9 2 9 13 7 9 9 13 2 13 3 13 7 3 13 2
25 0 9 13 9 7 9 2 9 15 13 2 16 1 9 1 9 2 3 1 9 7 1 0 9 2
7 9 3 13 7 9 9 2
43 9 0 9 1 9 13 7 3 0 2 7 15 2 1 2 12 9 2 7 0 9 0 9 2 7 7 15 2 16 1 9 4 13 7 0 9 9 1 11 1 0 9 2
2 0 9
33 1 0 9 2 9 9 11 7 9 0 9 11 2 13 1 9 12 1 0 9 13 7 1 9 13 0 9 12 2 12 0 9 2
13 3 0 9 13 3 0 9 1 9 13 7 13 2
10 3 0 9 9 15 13 7 13 9 2
28 1 15 13 7 0 9 2 3 15 9 1 9 9 0 9 13 1 0 12 9 3 13 7 3 13 1 9 2
5 12 9 1 15 2
47 16 0 9 13 1 9 0 9 9 1 9 2 1 15 0 9 13 9 9 11 1 11 2 13 1 0 12 9 2 12 9 0 2 12 9 2 12 11 1 9 7 10 9 3 0 9 2
2 9 9
14 1 10 0 9 15 13 3 9 2 7 7 0 9 2
16 9 0 9 1 0 9 11 0 2 0 9 9 13 3 9 2
24 7 15 1 15 13 3 13 0 9 2 3 9 1 0 9 2 15 13 3 1 9 1 9 2
19 1 9 0 13 3 3 3 13 9 7 3 15 3 13 1 9 1 9 2
20 10 7 15 0 9 15 13 3 1 9 16 13 9 2 9 2 9 7 9 2
13 15 3 13 0 9 2 15 13 3 13 7 13 2
13 15 15 13 0 9 2 3 15 13 3 0 9 2
17 1 15 1 15 3 13 1 9 2 16 15 13 1 12 12 9 2
24 13 15 3 1 9 2 16 4 13 3 1 9 2 7 3 13 9 2 16 4 15 13 3 2
28 1 0 0 9 4 3 1 0 9 3 9 13 7 3 15 13 15 13 2 16 3 13 15 0 9 3 0 2
3 3 3 2
18 1 10 9 13 3 13 2 16 3 13 9 1 9 2 0 10 9 2
32 7 13 3 10 9 3 4 2 16 10 9 2 15 4 1 9 0 9 13 9 9 11 2 13 3 0 9 7 4 3 13 2
45 0 9 3 13 1 9 2 16 9 13 3 3 13 1 9 0 0 9 1 9 15 2 15 0 0 9 2 14 3 9 9 11 2 3 13 15 1 0 9 2 13 1 0 9 2
36 1 9 0 9 15 3 3 13 9 9 0 0 9 7 9 7 9 9 1 9 9 7 9 2 0 0 7 0 0 9 0 9 7 0 9 2
17 15 0 3 13 0 0 9 9 7 9 10 9 2 15 13 9 2
60 1 0 9 3 0 9 9 2 9 7 9 2 13 2 14 3 0 0 9 1 9 0 7 0 9 2 9 1 12 9 13 7 10 9 2 15 13 2 13 9 0 9 11 1 9 0 9 2 1 0 0 0 9 1 12 9 10 0 9 2
4 9 1 9 2
7 9 9 1 9 1 0 9
5 2 12 2 12 2
5 0 9 9 1 9
5 2 1 9 9 2
8 2 9 2 9 9 11 11 2
4 9 1 9 2
14 9 15 13 7 10 2 9 2 13 0 9 9 1 9
4 14 15 3 13
7 0 9 13 9 1 9 2
5 0 9 13 13 0
8 12 9 13 9 10 9 13 2
23 13 1 15 13 7 0 9 9 9 0 0 7 0 9 1 11 2 11 2 11 7 11 2
21 9 15 13 9 0 9 1 0 9 0 9 7 9 7 3 0 9 13 10 9 2
20 11 11 2 9 9 9 7 9 11 2 0 0 9 13 3 1 12 9 9 2
9 1 15 15 13 9 9 12 9 2
21 1 0 9 13 10 7 0 9 3 1 9 9 9 7 9 1 9 7 0 9 2
18 1 0 9 3 13 9 1 9 0 9 7 9 1 9 7 0 9 2
13 11 11 2 11 11 2 0 9 13 14 12 9 2
21 13 3 1 0 9 7 0 7 0 9 1 10 9 1 10 9 0 9 1 9 2
21 13 1 0 9 9 1 9 0 9 2 15 15 13 1 9 0 9 9 7 9 2
11 9 1 0 9 13 7 1 15 3 0 2
17 15 1 11 13 3 12 9 2 15 15 1 15 13 9 7 12 2
33 11 11 2 9 9 0 9 9 11 2 10 10 9 13 2 16 0 9 13 1 0 11 3 0 9 2 15 3 13 1 0 9 2
19 13 15 15 3 1 0 9 1 9 0 1 9 2 7 7 1 0 9 2
16 1 1 0 9 1 0 9 13 13 13 3 7 1 0 9 2
16 3 10 0 9 3 13 9 9 2 15 13 1 9 0 9 2
7 13 1 15 7 0 9 2
38 11 11 2 0 9 1 9 11 1 11 2 0 9 2 16 4 15 0 9 13 13 1 0 9 2 13 0 0 9 1 0 9 2 3 9 7 9 2
17 9 2 15 13 1 11 13 2 13 13 0 9 9 1 10 9 2
15 0 9 13 9 2 15 4 13 15 0 0 9 7 9 2
23 1 9 1 0 9 7 9 1 15 13 9 0 9 2 15 13 9 13 7 13 1 0 2
13 9 9 13 0 2 1 0 9 14 1 0 9 2
22 11 11 2 0 9 11 7 11 2 0 9 4 15 13 1 11 13 3 3 16 3 2
21 13 0 2 16 4 15 13 0 9 9 9 0 9 2 1 9 1 9 0 9 2
18 1 0 9 13 9 13 15 0 9 2 15 15 3 13 1 0 11 2
13 0 9 13 3 1 0 9 2 9 7 0 9 2
16 11 11 2 0 9 11 2 13 1 11 10 0 0 0 9 2
18 3 9 11 1 0 11 0 1 0 9 9 1 9 0 7 0 9 2
11 9 9 13 3 0 7 9 13 3 0 2
25 3 16 13 3 0 9 0 9 1 11 7 11 2 13 9 13 3 2 7 0 9 1 15 13 2
5 0 9 1 0 9
6 0 9 9 13 9 2
7 13 13 3 1 9 1 11
24 1 0 9 1 11 4 13 9 16 0 0 9 13 0 0 9 0 0 9 9 11 2 11 2
29 9 13 1 15 0 2 16 1 0 9 13 9 2 15 1 0 9 13 1 9 1 9 1 0 9 0 0 9 2
7 9 15 13 7 0 9 2
3 13 11 11
20 9 0 9 1 9 11 2 11 13 1 9 12 7 12 1 3 16 12 9 2
22 9 9 15 1 0 9 13 1 12 1 12 7 9 1 12 9 9 1 12 9 9 2
10 7 13 1 0 9 9 0 9 13 2
18 9 13 1 0 9 0 9 2 15 1 9 13 13 7 3 3 13 2
3 9 1 0
29 1 9 1 0 9 0 9 11 2 11 4 13 1 9 0 9 2 0 9 7 0 9 2 15 13 13 1 9 2
10 9 3 13 3 1 9 14 1 9 2
13 0 0 9 2 15 15 3 13 0 2 13 0 2
24 3 15 13 9 1 0 9 2 15 13 1 9 13 7 0 9 2 3 9 0 1 9 9 2
13 0 9 13 7 9 9 2 15 9 13 1 9 2
31 1 0 9 9 1 9 15 13 1 10 0 9 2 1 15 4 0 7 0 9 13 1 0 9 1 0 9 7 0 9 2
9 9 9 3 13 1 9 12 9 2
8 0 9 1 15 13 12 9 2
30 0 9 13 9 12 9 1 9 1 9 0 9 0 9 9 2 13 15 0 7 13 0 9 7 13 15 0 0 9 2
31 0 9 15 0 9 2 15 13 12 7 12 9 2 1 15 2 15 13 9 1 0 7 0 9 2 13 9 13 1 9 2
13 9 0 9 15 3 0 9 13 13 1 0 9 2
8 9 0 9 13 1 0 9 2
11 0 9 1 9 11 2 11 13 3 0 2
27 3 1 9 9 9 0 0 9 15 15 13 2 16 15 15 13 13 9 9 9 1 9 14 1 12 5 2
37 9 3 0 9 15 13 1 12 9 1 0 12 9 2 1 0 9 15 13 9 9 1 0 9 1 12 1 12 9 7 9 1 12 1 12 9 2
19 3 13 3 0 9 2 3 9 13 10 3 0 9 2 13 12 1 9 2
27 1 9 9 15 13 2 16 4 9 9 13 13 3 9 3 2 15 1 9 13 1 10 9 0 9 0 2
15 3 12 9 1 9 9 13 0 3 0 0 9 1 9 2
18 1 12 9 0 9 9 13 1 0 9 1 9 0 9 1 12 5 2
8 13 1 15 7 0 9 9 2
23 1 9 13 1 9 11 2 11 1 0 2 7 3 0 9 2 15 3 13 9 1 9 2
13 13 4 15 2 16 13 9 9 0 1 0 9 2
17 9 15 0 9 9 3 13 2 16 15 3 2 3 13 9 9 2
3 14 1 11
15 1 9 13 9 9 11 2 11 14 3 13 1 0 9 2
17 1 9 12 13 1 11 1 0 9 0 3 16 12 5 0 9 2
13 3 15 10 9 13 13 1 12 5 1 0 9 2
24 3 1 0 11 15 13 1 0 9 1 12 1 12 5 7 1 11 1 12 5 1 12 5 2
19 9 15 13 13 0 9 1 9 0 0 9 1 12 1 12 5 0 9 2
21 13 15 15 9 1 0 9 2 0 9 0 0 2 15 3 13 12 5 0 9 2
16 1 9 11 2 11 13 0 9 7 9 1 0 7 0 11 2
3 9 1 11
17 0 9 13 9 1 11 7 0 9 13 3 1 9 1 0 9 2
30 13 2 16 13 1 15 0 9 0 9 7 13 0 9 2 13 11 11 2 1 9 9 2 3 13 1 9 3 11 2
22 1 11 13 0 9 13 1 0 9 9 9 12 2 16 4 13 3 9 9 1 9 2
23 13 15 15 2 16 13 13 9 0 9 1 0 9 2 15 13 1 10 9 16 3 0 2
34 1 9 2 16 11 2 11 13 1 9 1 0 0 7 0 9 2 13 13 11 13 7 13 3 9 1 3 0 9 16 1 0 11 2
27 11 2 11 13 3 1 11 11 1 9 0 0 9 2 15 4 13 3 1 0 9 7 13 13 12 9 2
11 9 13 3 0 0 9 0 0 0 9 2
18 13 3 1 10 0 9 2 15 4 13 1 9 11 11 0 9 13 2
4 9 1 9 2
3 9 2 12
2 9 9
8 9 1 9 2 9 1 9 2
5 13 16 0 9 2
15 15 15 15 13 3 2 13 9 13 1 0 9 7 13 2
3 3 0 9
6 0 9 13 12 9 2
7 9 3 1 9 1 12 9
9 9 0 9 1 11 15 3 13 2
18 0 9 1 0 9 4 13 3 0 9 2 1 0 9 1 12 9 2
26 3 15 15 13 2 16 4 13 9 2 16 15 13 9 13 1 9 2 3 15 15 15 13 1 11 2
12 3 9 12 2 9 7 13 0 9 0 9 2
16 9 13 1 9 9 3 2 13 15 2 9 0 9 13 0 2
8 0 0 9 15 13 0 9 2
12 9 3 13 12 9 9 1 0 9 11 3 2
20 3 1 15 13 0 0 9 1 11 0 9 0 9 2 15 4 13 9 13 2
3 9 1 9
12 0 0 9 13 0 9 0 14 9 0 9 2
33 3 13 9 12 12 9 7 3 16 12 9 9 2 15 13 9 1 0 11 2 13 11 11 2 9 0 0 9 2 1 9 2 2
19 10 9 9 13 9 7 9 13 1 15 9 7 1 9 3 1 9 9 2
21 1 9 15 3 13 2 16 9 1 9 13 9 7 9 13 1 9 1 0 9 2
16 1 9 13 7 3 9 2 15 13 1 0 9 1 0 11 2
15 13 15 13 9 9 1 9 2 16 15 0 9 13 0 2
2 0 9
21 9 0 1 9 13 3 13 0 9 2 15 13 0 9 1 9 1 9 0 9 2
29 1 12 9 0 9 4 9 7 9 13 1 9 7 4 13 1 9 2 15 15 13 1 9 2 7 1 0 9 2
25 0 9 13 9 9 1 9 2 15 4 13 1 9 7 13 3 2 16 4 3 13 0 9 9 2
13 1 9 9 13 9 1 15 2 16 15 9 13 2
26 9 15 13 2 16 15 0 9 13 1 12 9 2 14 12 5 15 13 1 9 3 0 7 0 9 2
9 3 15 13 1 9 10 12 9 2
13 1 15 9 3 14 12 9 9 13 1 9 3 2
16 13 15 15 9 9 9 2 15 13 7 0 2 7 0 9 2
21 3 15 3 13 1 12 9 11 2 7 9 2 15 3 7 3 13 1 9 9 2
11 7 3 0 9 0 0 9 3 12 13 2
33 13 3 13 0 9 0 9 2 15 13 3 1 0 9 7 9 3 2 16 13 0 0 9 13 14 9 2 7 3 7 0 9 2
14 15 15 13 9 9 7 9 9 3 1 0 0 9 2
7 9 1 9 2 0 9 2
9 13 9 9 3 1 9 1 9 2
2 3 2
2 13 2
19 1 12 9 9 1 11 13 1 9 0 9 9 9 11 1 0 9 9 2
18 1 0 15 13 0 9 2 0 12 9 12 7 9 1 12 12 9 2
13 9 13 0 9 1 12 9 9 1 11 2 11 2
18 12 9 1 9 2 3 13 9 13 10 9 2 15 13 13 0 9 2
5 13 15 0 9 2
8 16 4 9 13 9 7 3 2
2 9 9
6 9 13 1 0 9 2
11 9 1 9 13 1 9 7 3 13 13 2
9 9 1 9 13 9 7 9 13 2
17 3 13 7 9 3 1 9 13 12 9 9 12 9 9 12 9 2
19 13 7 7 9 2 15 1 0 9 9 13 2 16 0 9 13 3 9 2
13 9 13 10 9 13 1 9 1 0 9 7 9 2
2 9 1
21 1 9 9 2 15 13 1 9 11 11 2 13 9 9 12 1 9 9 0 9 2
10 15 15 13 1 12 9 1 9 11 2
14 1 9 13 9 13 1 9 0 9 11 12 1 11 2
8 0 9 9 1 10 9 13 2
7 0 9 1 9 9 13 2
24 2 0 9 2 15 13 9 1 12 9 2 13 3 0 7 13 9 9 9 1 0 9 9 2
34 2 0 9 9 13 0 9 1 0 9 2 13 15 9 12 9 2 7 1 0 9 7 9 12 5 12 2 3 2 12 5 12 9 2
14 2 9 1 9 12 13 13 0 1 9 1 0 9 2
21 2 0 9 9 13 0 3 3 13 1 0 9 1 9 2 1 9 9 7 3 2
4 15 13 1 2
22 9 1 9 9 0 9 11 13 9 1 12 9 9 7 0 0 9 13 12 9 9 2
22 9 1 9 1 11 2 11 13 1 12 2 9 12 1 9 0 9 14 12 9 12 2
6 13 15 7 3 3 2
17 10 0 9 15 13 2 13 11 11 2 0 9 2 1 9 2 2
10 3 13 2 1 15 1 0 9 13 2
17 2 9 0 9 13 2 14 3 13 1 9 7 9 1 0 9 2
13 0 9 13 3 9 13 2 3 15 1 15 13 2
15 1 0 9 9 13 9 0 2 16 13 1 12 9 9 2
13 2 0 9 13 0 13 1 9 9 7 0 9 2
17 3 7 13 13 0 9 2 9 13 9 13 7 13 15 1 15 2
15 2 0 13 0 9 1 9 2 15 9 7 9 9 13 2
13 9 1 9 13 0 3 1 9 0 7 0 9 2
8 1 9 15 13 7 13 3 2
8 3 3 2 16 13 9 3 2
9 16 4 13 9 2 13 15 0 2
2 11 11
34 9 2 9 2 0 2 9 2 2 11 12 2 12 12 11 2 9 2 2 2 12 2 12 12 12 2 9 2 2 12 2 12 12 12
3 9 2 12
3 9 2 11
7 9 2 11 2 9 2 11
8 0 9 2 9 0 11 1 11
6 9 1 9 9 2 12
4 9 9 2 12
5 9 2 13 1 9
9 9 2 9 2 13 13 1 9 2
7 9 12 2 12 2 12 2
27 9 2 9 11 13 1 0 9 3 12 9 1 0 2 11 2 15 3 3 13 1 0 9 1 11 11 2
8 1 9 13 9 7 0 9 2
7 12 0 9 13 1 9 2
15 0 9 1 9 13 13 9 2 16 13 0 0 9 9 2
8 9 13 1 12 7 12 9 2
13 1 9 13 1 9 9 7 9 7 9 1 9 2
10 1 9 13 9 2 9 7 9 9 2
4 9 1 9 2
3 9 2 12
4 9 2 11 11
5 9 2 11 2 11
5 0 9 2 0 9
6 9 1 9 9 2 12
4 9 9 2 12
4 9 2 14 9
3 9 2 0
18 9 2 9 1 0 9 2 0 9 7 9 9 4 13 1 9 9 2
12 9 13 13 1 9 11 2 1 9 9 11 2
9 1 9 13 9 0 7 0 9 2
15 9 1 0 9 1 9 9 2 1 9 1 0 0 9 2
21 1 9 13 9 1 12 9 1 0 0 9 2 0 9 2 0 9 7 0 9 2
28 1 9 9 1 9 1 0 9 2 9 7 9 1 9 2 4 9 1 9 13 12 9 7 1 9 12 9 2
8 13 0 13 9 9 1 9 2
3 9 2 12
3 9 2 11
5 9 2 11 2 11
5 0 9 2 9 11
6 9 1 9 9 2 12
9 9 2 1 12 9 3 9 7 9
11 9 2 1 9 9 13 9 12 9 1 9
10 9 2 0 2 9 11 2 9 11 2
16 9 2 9 13 14 12 9 1 11 1 9 11 1 0 9 2
16 9 9 1 11 2 11 2 9 11 7 9 1 9 0 11 2
17 11 2 12 9 1 2 9 2 2 11 2 12 9 1 2 9 2
13 9 1 0 2 0 7 0 9 1 0 0 9 2
6 0 9 1 0 9 2
10 1 9 13 0 9 7 3 0 9 2
5 1 9 13 9 2
7 1 9 13 0 15 13 2
9 13 0 13 1 9 9 9 9 2
3 9 2 12
4 9 2 11 11
5 9 2 9 2 11
9 0 9 2 0 0 11 2 2 2
6 9 1 9 9 2 12
4 9 9 2 12
3 9 2 9
16 9 2 3 2 9 1 11 3 1 9 2 13 12 2 12 2
22 9 2 0 9 13 1 0 9 11 2 14 10 9 1 9 2 7 3 3 0 9 2
11 9 4 1 0 9 13 7 13 0 9 2
18 1 9 9 13 9 0 11 2 9 2 9 0 9 7 9 1 9 2
9 0 0 9 1 9 2 12 9 2
12 1 9 13 9 2 1 9 2 7 0 9 2
13 1 9 13 12 9 2 9 1 9 7 0 9 2
9 1 9 1 0 9 9 7 9 2
15 9 13 9 2 9 2 9 2 9 7 9 1 0 9 2
9 9 13 1 0 9 7 0 9 2
3 9 2 12
3 9 2 11
7 9 2 11 2 11 2 11
9 0 9 2 9 0 9 2 2 2
6 9 1 9 9 2 12
18 9 2 1 12 1 12 9 3 2 1 12 1 12 9 12 5 9 2
4 9 2 9 2
11 9 2 3 1 11 12 2 12 2 12 2
11 9 2 11 15 13 1 9 0 9 11 2
14 1 9 13 9 9 11 2 0 9 7 0 0 9 2
7 13 9 9 7 0 9 2
15 9 11 2 3 13 9 2 13 1 11 13 14 12 9 2
10 0 9 13 9 2 15 13 1 9 2
7 1 9 13 9 0 9 2
7 13 13 3 0 0 9 2
8 1 9 13 1 9 12 9 2
9 0 9 1 9 7 9 1 9 2
15 1 9 13 9 2 12 9 2 9 2 0 9 7 9 2
13 9 2 9 9 0 9 7 9 1 12 0 9 2
10 9 1 0 9 13 0 14 1 9 2
23 1 9 13 13 9 1 9 2 15 15 13 1 9 1 9 7 13 12 9 7 12 9 2
3 9 2 12
3 9 2 11
6 9 2 11 2 0 9
8 0 9 2 9 11 2 2 2
6 9 1 9 9 2 12
12 9 9 2 12 2 1 12 9 14 9 1 12
3 9 2 9
8 9 2 3 12 2 12 2 12
19 9 2 0 9 15 13 1 0 9 11 2 9 11 13 10 9 0 9 2
16 0 9 1 11 13 0 9 2 0 9 13 13 7 1 11 2
18 1 0 0 9 13 0 13 9 1 11 2 11 2 11 2 11 3 2
26 9 13 13 14 12 9 1 0 9 2 1 9 0 9 11 1 10 9 2 9 7 9 1 0 9 2
7 9 2 3 9 7 9 2
7 3 13 1 9 10 9 2
14 9 13 0 7 0 1 9 2 9 2 9 7 9 2
8 9 2 9 9 9 7 9 2
3 9 2 12
3 9 2 11
5 9 2 11 2 11
10 0 9 2 9 11 2 9 2 9 2
6 9 1 9 9 2 12
4 9 9 2 12
3 9 2 9
15 9 2 9 1 11 12 9 1 9 1 12 2 12 2 12
18 9 2 9 11 13 13 1 0 9 0 14 12 9 9 9 1 11 2
13 1 0 9 13 0 0 7 0 9 0 0 9 2
20 1 0 9 13 9 9 2 9 2 9 2 9 2 9 2 9 9 7 9 2
5 9 9 0 9 2
8 1 9 7 1 9 0 9 2
9 15 9 13 13 0 9 7 9 2
9 9 1 9 9 0 9 7 9 2
8 9 0 9 1 9 12 9 2
3 9 2 12
4 9 2 0 11
7 9 2 11 2 11 1 11
9 0 9 2 9 11 11 2 2 2
9 9 1 9 9 2 9 12 2 12
9 9 9 2 1 12 9 9 12 5
11 9 2 9 2 9 1 9 12 9 1 9
3 9 2 0
18 9 2 9 13 13 1 9 11 1 11 2 1 9 11 1 0 9 2
25 13 3 12 9 0 0 9 2 15 15 3 13 1 9 2 15 13 0 3 1 9 1 0 9 2
12 9 13 3 12 9 1 9 0 14 0 9 2
10 1 9 13 3 1 9 9 7 9 2
8 0 9 1 9 9 1 9 2
8 0 9 2 0 9 1 9 2
8 9 1 9 2 9 7 9 2
6 1 9 13 14 9 2
9 1 9 9 7 9 1 0 9 2
7 9 0 2 0 7 0 2
4 9 1 9 2
5 9 2 13 4 13
3 1 9 9
14 1 9 9 1 9 1 0 9 15 3 13 9 9 2
13 3 13 15 1 9 1 9 2 15 13 1 9 2
4 11 11 2 11
42 9 2 1 3 13 9 9 2 13 7 13 0 9 1 9 1 9 2 3 7 3 15 13 13 7 3 15 13 0 9 2 13 9 9 12 1 9 1 9 9 2 2
41 1 10 0 0 9 13 13 9 3 0 9 0 1 9 2 15 13 1 9 1 0 9 2 9 12 9 12 9 9 12 2 12 9 2 2 1 9 0 9 2 2
7 1 9 9 13 0 9 2
4 12 2 9 2
14 1 9 2 1 15 15 13 9 9 2 13 13 9 2
6 1 9 3 0 13 2
9 9 2 9 0 3 16 1 9 2
8 9 2 9 0 1 9 9 2
5 12 2 0 9 2
8 1 0 9 3 13 0 9 2
18 0 9 2 1 15 4 9 13 2 13 13 2 9 12 0 9 2 2
18 2 9 1 9 2 10 0 9 2 9 7 9 9 2 0 0 9 2
7 2 0 9 1 10 9 2
5 2 0 9 9 2
6 2 9 7 9 9 2
5 2 9 9 9 2
4 2 9 9 2
6 2 9 1 9 3 2
4 2 9 9 2
5 2 9 9 3 2
21 9 2 1 15 10 9 13 2 7 13 0 15 3 13 2 13 4 0 9 13 2
17 1 0 0 9 2 9 1 0 2 15 9 0 9 13 13 15 2
16 12 2 9 13 1 10 0 9 9 2 9 12 0 9 2 2
22 9 3 0 9 0 1 9 2 0 14 3 3 1 9 1 9 9 2 13 12 9 2
19 0 9 13 1 12 2 9 9 9 0 16 9 12 2 9 1 9 9 2
21 0 9 15 9 2 15 13 16 9 9 13 1 12 9 1 10 9 1 0 9 2
10 12 2 9 1 9 15 1 9 13 2
12 13 15 7 13 1 9 9 1 9 12 9 2
3 2 2 2
4 9 1 9 2
35 0 9 2 15 15 0 9 1 9 9 9 13 2 13 0 9 2 9 1 9 1 9 9 12 2 12 9 2 2 1 9 0 9 2 2
9 1 9 15 13 9 0 0 9 2
8 11 11 2 0 9 11 2 9
5 1 9 15 9 13
5 3 0 1 9 13
18 12 9 13 1 9 0 9 1 9 11 1 0 9 14 12 9 9 2
13 1 12 1 0 0 9 13 9 1 9 10 9 2
30 9 4 15 13 1 9 0 9 12 9 2 15 7 13 0 9 7 10 9 13 1 9 2 16 0 9 13 15 15 2
16 9 2 0 13 1 9 0 9 12 9 9 2 15 3 13 2
16 16 0 13 3 0 9 2 4 0 9 3 1 12 9 13 2
20 9 13 3 0 13 9 9 1 9 0 9 3 1 9 9 9 1 0 9 2
47 0 9 13 9 1 9 1 9 9 2 0 1 9 9 2 9 1 15 13 3 0 9 2 1 15 2 16 13 2 13 9 2 3 2 16 4 0 9 13 1 9 13 1 9 0 9 2
8 9 13 10 9 13 0 9 2
9 15 2 3 15 3 13 2 13 2
5 0 9 3 13 2
8 0 9 15 13 13 0 9 2
49 13 15 7 2 16 0 9 9 13 2 1 0 9 2 1 9 12 9 9 13 9 2 13 7 0 9 2 15 1 9 1 9 13 1 9 0 9 14 12 9 2 7 1 0 9 13 0 9 2
31 1 9 0 9 0 9 13 3 9 1 9 2 7 3 1 12 5 9 1 0 9 2 15 13 14 12 5 1 9 9 2
12 3 13 15 0 2 16 13 0 9 0 9 2
6 15 13 13 3 3 2
9 9 13 9 1 9 1 12 9 2
7 1 9 15 13 15 13 2
2 9 2
14 2 7 0 9 9 13 9 13 15 1 9 10 9 2
23 2 13 2 14 0 9 2 13 9 1 0 9 2 3 16 13 1 0 7 3 0 9 2
4 11 11 2 11
22 9 0 1 10 9 2 0 1 0 9 9 2 13 3 13 7 3 13 9 12 9 2
10 4 3 13 1 0 9 1 12 9 2
19 13 15 1 15 2 10 9 4 15 1 9 13 7 10 1 15 13 9 2
2 9 9
2 12 5
24 1 0 12 9 0 9 13 12 9 9 1 0 9 1 0 9 2 1 9 7 0 2 9 2
18 1 0 7 0 9 11 12 15 13 11 11 2 9 9 1 0 9 2
32 0 9 13 1 9 3 1 9 9 0 9 7 13 0 9 2 16 15 3 1 9 13 0 9 2 15 9 13 15 1 9 2
32 1 0 0 9 15 13 7 0 2 15 13 3 3 7 3 0 16 1 0 9 7 1 10 9 13 0 9 14 12 9 9 2
23 7 16 13 9 9 1 9 0 2 13 15 1 9 0 9 7 13 4 0 10 9 13 2
4 2 0 9 2
3 9 9 9
11 1 9 12 10 0 9 13 9 12 9 2
12 13 4 9 9 0 7 9 9 9 1 9 2
3 9 13 2
32 13 15 2 16 9 2 15 13 13 1 0 9 2 13 13 9 1 9 9 9 1 9 0 9 1 9 12 9 1 9 12 2
11 7 1 9 12 10 9 13 9 12 9 2
11 13 9 13 9 1 9 9 1 9 12 2
4 11 11 2 11
36 1 3 9 1 9 12 3 13 13 2 1 9 12 1 10 9 0 9 13 9 2 15 7 13 13 0 7 0 9 1 9 0 9 7 9 2
19 16 4 7 1 0 9 13 0 7 9 1 9 2 13 15 1 15 3 2
11 1 9 9 15 0 9 9 9 13 13 2
4 10 0 9 2
2 0 9
24 0 9 1 0 9 7 11 15 13 3 13 14 1 9 12 2 16 0 9 13 1 9 12 2
24 1 0 9 13 0 9 1 0 12 9 0 9 9 12 9 0 9 2 14 12 9 9 2 2
15 13 15 14 1 12 5 3 16 1 0 9 1 9 12 2
21 1 0 9 15 3 13 9 7 0 9 2 0 9 2 9 7 9 2 3 9 2
18 0 9 15 3 3 13 1 9 11 2 9 2 9 2 9 7 9 2
11 1 0 9 13 0 9 9 1 0 9 2
3 9 15 13
17 9 0 9 1 0 9 13 3 0 16 1 9 0 9 0 9 2
13 1 0 9 13 0 9 1 11 3 12 9 9 2
23 13 15 3 7 3 2 16 1 11 13 9 14 0 7 0 9 2 15 1 9 3 13 2
21 1 0 12 7 12 9 13 2 3 1 9 9 2 11 13 12 7 12 9 9 2
17 3 15 13 9 0 9 1 0 11 2 13 15 9 1 9 9 2
3 9 0 9
33 0 9 0 9 13 9 0 9 2 15 13 13 7 13 0 9 2 1 11 2 3 13 13 1 0 9 2 15 13 13 0 9 2
19 13 3 9 0 9 0 9 2 15 13 9 2 9 2 3 1 0 9 2
1 9
16 1 0 9 1 11 0 12 9 13 0 9 3 0 0 9 2
15 1 0 0 9 13 9 13 0 9 1 0 9 1 11 2
13 13 13 9 0 9 2 15 15 13 0 9 13 2
17 0 9 13 0 0 9 13 3 9 1 11 2 15 1 9 13 2
35 9 2 9 0 9 2 1 0 9 12 2 12 12 11 12 2 9 2 2 2 12 2 12 12 12 2 9 2 2 12 2 12 12 12 2
2 10 9
3 9 1 9
8 2 9 9 2 12 2 12 2
15 16 9 9 13 0 1 0 9 13 9 1 0 0 9 2
19 7 1 0 9 15 3 3 9 9 13 13 9 1 9 10 9 1 9 2
23 13 9 1 10 9 12 9 1 9 9 9 1 9 2 7 3 14 1 9 9 0 9 2
30 1 1 15 2 16 9 9 13 9 1 9 2 7 7 1 9 2 13 15 3 2 16 3 0 9 13 3 1 9 2
22 13 15 7 13 14 1 9 7 9 2 3 1 0 9 9 13 3 12 7 12 9 2
25 16 9 3 0 9 13 13 1 12 9 9 2 15 13 15 0 2 2 3 13 16 9 9 13 2
21 7 13 15 13 1 9 2 16 9 15 13 12 2 12 9 1 9 9 1 9 2
29 13 15 2 16 13 0 9 2 15 4 9 13 2 16 4 13 1 10 9 0 12 9 1 9 9 9 0 9 2
24 10 0 9 7 0 9 13 2 16 13 9 2 15 13 0 9 7 13 15 9 1 0 9 2
12 3 13 3 0 2 16 9 0 9 13 0 2
25 7 0 9 1 10 9 13 9 1 9 9 2 16 0 9 1 9 15 13 13 1 15 2 9 2
5 11 11 2 0 11
3 9 1 9
9 2 9 9 9 2 12 2 12 2
41 1 0 7 0 9 4 15 13 9 2 15 4 13 3 9 9 9 2 12 2 12 9 2 2 15 13 9 9 2 12 2 12 9 2 2 1 9 9 7 9 2
22 10 9 1 9 12 13 9 13 0 0 9 1 0 0 9 1 12 2 12 2 12 2
17 3 1 9 9 1 9 9 4 13 13 9 13 1 9 9 9 2
60 1 9 9 9 3 13 12 9 2 9 9 2 12 2 12 9 2 2 1 9 0 9 2 1 15 15 1 9 12 13 1 0 2 16 9 9 11 13 1 9 9 3 7 3 13 9 9 2 7 2 0 9 2 7 1 9 9 9 9 2
34 1 9 1 12 9 2 3 9 9 13 9 9 2 12 2 12 9 2 9 9 2 0 9 2 1 9 10 9 1 9 12 9 3 2
52 9 1 9 9 13 0 3 1 9 2 16 9 4 13 9 1 9 1 9 2 13 2 14 0 0 9 0 16 0 9 2 13 0 13 9 1 12 2 12 2 7 9 1 9 9 13 0 1 12 2 12 2
6 11 11 2 11 2 11
4 9 1 9 2
20 13 1 9 2 16 9 9 2 9 7 9 0 9 1 9 1 9 13 0 2
15 13 15 9 9 0 9 1 0 9 0 0 9 11 11 2
23 13 15 2 16 0 9 13 3 1 0 0 0 9 2 15 15 13 0 9 7 0 9 2
15 0 9 13 1 9 9 2 7 3 1 9 1 9 9 2
22 3 9 1 9 0 0 9 13 1 3 0 9 9 2 16 1 9 0 9 7 9 2
4 11 11 2 11
3 9 7 9
54 16 0 0 7 0 9 1 11 13 3 9 2 7 13 4 15 3 7 3 15 2 15 4 13 0 13 9 0 7 0 9 3 2 16 4 13 0 1 9 13 14 1 10 9 7 3 0 9 1 0 9 13 3 2
33 13 15 14 0 9 2 7 13 15 1 15 9 2 16 15 3 13 9 0 13 0 9 1 0 9 9 2 7 3 7 1 0 2
28 16 13 1 9 10 9 7 10 9 2 13 15 13 7 0 9 2 3 7 3 2 16 13 9 1 0 9 2
18 13 0 9 2 15 0 9 13 7 3 15 7 9 9 0 9 13 2
11 13 15 3 1 0 9 1 3 0 9 2
4 11 11 2 11
3 0 9 2
5 1 11 3 1 9
8 2 9 9 2 12 2 12 2
32 0 9 0 15 3 9 1 0 9 13 9 2 16 14 9 2 7 3 10 9 15 13 13 2 16 10 0 9 13 0 13 2
15 1 11 15 15 13 9 0 1 9 7 10 9 1 9 2
19 13 15 15 0 2 7 13 0 9 9 13 1 0 3 0 7 0 9 2
21 14 2 9 13 9 2 15 13 9 7 3 9 2 7 1 15 13 13 0 9 2
16 1 15 13 0 3 3 13 2 16 3 0 9 15 3 13 2
6 11 11 2 11 1 11
6 9 2 0 9 7 15
1 11
11 10 0 0 0 9 13 13 1 9 12 2
7 13 9 9 1 0 9 2
18 1 9 13 1 0 0 9 9 2 9 2 9 7 0 9 1 9 2
13 9 13 12 9 7 13 0 9 1 12 9 9 2
13 1 0 9 11 13 11 2 11 2 11 7 11 2
9 1 0 9 13 9 14 12 9 2
15 1 9 13 3 1 9 9 2 1 9 13 15 0 9 2
16 14 12 5 9 13 11 1 9 2 0 12 5 13 3 9 2
10 1 9 13 0 9 1 11 3 13 2
14 13 4 1 9 9 7 1 9 0 9 13 0 9 2
31 1 9 9 2 15 13 13 9 0 9 2 13 1 9 0 9 2 13 11 11 2 0 9 11 9 2 1 9 2 0 2
5 2 1 9 2 2
21 9 13 1 11 1 0 9 9 7 1 9 0 9 9 7 9 7 1 11 9 2
35 9 2 11 9 2 1 9 2 0 2 2 0 12 2 12 12 11 12 2 9 2 2 9 2 2 12 2 12 12 12 2 12 12 12 2
4 2 0 9 2
12 0 9 11 13 0 9 2 0 1 9 9 2
21 13 9 9 1 0 9 9 2 9 1 0 9 2 0 2 0 9 11 7 3 2
12 3 13 1 0 9 1 3 3 12 9 9 2
23 9 0 9 13 3 9 13 1 9 0 9 7 9 2 3 1 9 13 9 1 0 9 2
16 3 0 9 13 0 9 0 9 2 15 13 14 1 9 9 2
26 1 0 9 13 9 9 1 0 0 9 1 11 2 11 2 11 2 11 2 7 1 11 2 11 2 2
27 1 9 9 2 9 13 1 9 1 9 0 9 2 9 0 0 9 0 1 0 9 2 7 0 0 9 2
2 11 11
39 9 2 0 9 2 0 9 11 2 0 12 2 12 12 11 12 2 9 2 2 12 2 12 12 2 12 12 2 9 2 5 9 2 2 12 2 12 12 2
1 9
2 0 9
16 3 0 0 9 0 0 9 1 0 9 13 1 0 0 9 2
9 3 15 13 13 12 9 9 9 2
20 1 0 9 10 0 9 13 0 9 1 11 2 11 2 11 7 9 9 11 2
35 0 9 15 13 13 1 0 9 9 2 15 13 13 1 9 12 14 1 12 0 2 7 3 9 2 7 7 0 9 13 1 0 9 9 2
30 0 9 13 0 0 9 15 0 9 9 7 0 9 2 16 4 13 9 10 9 1 0 9 0 9 0 11 1 11 2
3 1 0 9
15 9 9 13 1 10 9 11 2 11 2 11 11 0 11 2
17 3 10 0 9 13 1 9 12 9 9 0 9 1 12 9 9 2
15 0 9 0 7 0 9 13 1 0 9 0 9 0 9 2
10 9 13 1 9 3 16 12 9 9 2
26 0 0 9 15 13 1 11 2 11 2 1 0 9 7 0 11 2 13 15 7 1 9 0 0 9 2
2 9 11
15 0 9 11 13 3 9 1 10 9 1 11 1 0 11 2
20 1 0 0 9 13 12 9 9 0 11 2 11 2 13 9 1 12 9 9 2
15 1 0 9 9 13 12 9 11 0 11 9 12 9 9 2
27 1 0 9 9 13 12 9 7 9 1 0 9 9 11 2 9 9 2 9 9 2 9 9 7 0 9 2
4 3 11 13 9
10 9 1 9 2 13 15 2 15 13 9
10 9 7 9 15 1 10 9 13 3 2
13 14 13 15 15 2 16 3 9 13 3 1 9 2
8 9 0 9 11 15 7 13 2
22 3 2 1 0 9 2 12 9 9 2 15 13 13 2 16 10 9 9 1 9 13 2
26 9 1 9 2 3 11 13 9 7 0 9 1 9 0 9 2 13 0 9 9 11 11 1 12 9 2
12 12 2 13 15 0 16 9 2 1 0 9 2
14 12 2 16 0 3 2 1 0 9 9 7 9 9 2
3 3 15 13
38 13 9 9 2 15 1 15 13 1 9 9 7 1 15 3 13 0 9 2 9 1 0 9 2 7 3 1 0 0 9 2 13 15 9 11 9 11 2
7 13 15 0 9 1 9 2
7 9 11 13 1 12 9 2
8 1 9 1 15 13 0 9 2
20 13 15 15 14 1 0 9 2 7 15 2 16 15 13 0 9 1 0 9 2
17 7 9 3 13 9 7 0 7 13 1 0 9 2 13 10 9 2
21 16 13 15 9 2 13 9 7 9 2 13 9 1 0 9 7 1 0 0 9 2
16 3 3 13 0 9 7 13 1 9 9 2 1 15 3 13 2
12 16 2 15 1 15 2 15 10 0 9 13 2
19 11 3 13 1 9 9 13 1 9 9 1 9 2 15 15 3 3 13 2
19 9 9 13 7 16 9 0 9 13 1 15 0 7 3 0 16 0 9 2
18 3 3 13 1 9 3 3 0 0 9 1 0 9 1 9 0 9 2
13 7 1 10 9 13 0 11 1 9 1 9 13 2
5 3 13 15 0 2
20 1 0 9 4 9 1 9 13 13 15 2 9 0 9 13 2 13 9 9 2
8 13 7 1 15 13 9 9 2
10 10 9 2 7 9 3 15 3 13 2
16 15 2 15 13 13 10 0 9 2 3 1 15 13 0 9 2
5 1 9 3 9 2
2 0 9
32 16 4 13 1 10 9 13 3 0 9 16 9 1 0 9 2 13 4 15 13 1 12 2 12 9 3 2 13 15 9 11 2
12 13 4 15 1 0 9 7 13 4 15 3 2
11 16 13 0 9 2 13 1 0 9 9 2
16 7 3 13 7 11 13 1 15 2 16 0 9 15 13 3 2
14 14 0 0 9 13 7 0 2 13 9 9 9 9 2
11 10 9 15 13 1 0 9 1 9 9 2
23 9 9 2 1 9 3 0 9 9 2 7 9 0 0 9 1 3 0 2 13 9 13 2
7 3 7 1 9 10 9 2
10 1 0 9 15 0 9 13 0 9 2
14 13 15 15 13 3 1 0 11 2 13 15 9 11 2
6 13 3 0 0 9 2
9 1 0 9 13 3 0 9 0 2
27 3 15 10 9 13 9 3 14 1 10 9 2 0 3 13 9 0 9 1 9 2 16 15 9 13 15 2
13 3 1 0 9 15 3 3 13 0 9 1 9 2
23 1 9 1 11 13 9 7 9 2 16 0 9 13 0 0 9 2 12 9 1 9 9 2
17 9 0 7 0 9 13 1 0 9 1 0 9 13 0 0 9 2
20 1 11 13 1 15 2 16 4 9 9 13 0 0 9 1 9 0 9 9 2
13 1 0 9 13 7 12 9 2 13 15 9 11 2
30 3 2 3 9 13 12 9 2 13 0 9 3 2 1 9 9 7 9 13 2 16 13 0 9 1 12 9 1 9 2
2 11 11
33 9 2 11 11 2 9 2 9 2 9 2 0 12 2 12 2 12 12 11 12 2 9 2 2 9 2 2 12 2 12 2 12 2
11 11 13 1 0 11 2 3 13 0 0 9
2 9 9
3 9 1 9
4 11 2 11 2
33 9 2 11 11 2 0 0 9 9 2 9 2 0 7 0 9 2 12 2 2 12 2 12 2 12 2 0 9 11 9 2 9 2
30 0 11 9 2 12 2 0 0 9 9 2 0 7 0 9 2 12 2 2 12 2 12 2 12 2 0 9 11 9 2
32 11 2 0 9 9 9 2 9 2 9 7 0 9 2 12 2 2 12 2 12 2 12 2 0 9 11 9 2 9 2 9 2
30 11 2 0 0 9 9 2 9 2 0 9 7 0 9 2 12 2 2 12 2 12 2 12 2 0 9 11 2 9 2
4 11 2 11 2
33 9 2 12 2 0 0 9 2 0 9 2 0 7 0 9 2 9 2 9 9 2 0 9 2 12 2 2 12 2 12 2 12 2
20 11 2 12 2 0 9 9 7 0 9 2 12 2 2 12 2 12 2 12 2
56 0 9 0 11 2 0 2 0 2 2 11 1 11 7 11 0 11 2 9 2 9 2 0 2 2 9 11 11 2 12 12 11 2 0 12 2 9 2 2 2 12 2 12 2 12 2 9 2 2 12 2 12 2 12 12 2
4 11 2 11 2
19 9 2 12 2 0 0 7 0 9 2 12 2 2 12 2 12 2 12 2
39 9 1 11 2 9 2 12 12 11 1 11 2 0 9 12 2 9 2 2 2 12 2 12 12 2 12 12 2 12 12 2 9 2 2 12 2 12 12 2
4 11 2 11 2
17 9 2 12 2 9 5 9 2 12 2 2 12 2 12 2 12 2
21 11 2 12 2 0 9 9 7 9 1 9 2 12 2 2 12 2 12 2 12 2
36 11 2 12 2 0 9 9 2 9 2 9 2 9 2 9 2 9 2 9 7 9 1 0 7 0 9 2 12 2 2 12 2 12 2 12 2
55 9 11 11 1 11 2 11 11 2 11 2 2 9 2 9 2 0 2 2 12 12 11 2 9 12 2 9 12 2 9 2 2 2 12 2 12 12 2 12 12 2 12 12 2 9 2 2 12 2 12 12 2 12 12 2
4 11 2 11 2
11 0 9 2 0 9 2 9 2 0 9 2
7 9 2 0 9 7 9 2
5 9 7 0 9 2
13 0 0 9 2 12 2 2 12 2 12 2 12 2
38 9 9 1 11 2 0 11 2 11 2 9 12 11 2 12 11 9 2 2 9 2 2 2 12 2 12 2 12 2 12 2 9 2 2 12 2 12 2
23 9 2 9 0 9 2 9 2 2 2 12 2 12 12 2 9 2 2 12 2 12 12 2
1 9
22 9 9 11 2 9 2 9 2 0 2 2 15 1 9 9 11 13 1 9 1 11 2
24 1 9 12 2 9 13 9 0 9 1 0 9 1 9 1 9 2 7 3 1 15 3 0 2
17 10 9 2 15 10 0 9 13 2 13 13 9 1 9 9 9 2
7 0 9 1 0 0 9 2
1 9
3 14 7 14
12 10 9 1 9 15 13 16 0 2 0 9 2
19 9 14 7 14 2 1 9 9 1 9 1 0 9 2 1 15 3 13 2
47 13 9 0 9 2 15 15 13 1 9 7 1 9 2 3 0 9 7 0 9 2 1 0 9 1 9 9 2 16 4 15 3 3 2 3 16 7 9 9 2 13 3 7 3 15 13 2
22 13 15 3 13 2 9 2 2 3 0 7 0 9 9 2 14 2 7 2 14 2 2
28 9 14 7 14 13 13 15 2 15 15 15 13 2 13 15 1 0 9 2 13 13 0 9 2 9 7 9 2
59 9 9 11 11 15 13 2 1 10 9 9 4 13 15 2 15 2 3 13 2 13 7 15 1 9 10 9 2 0 9 2 3 13 2 3 13 2 14 2 15 2 15 13 1 15 0 2 7 2 14 2 15 2 15 13 1 15 0 2
28 9 2 9 11 2 0 12 2 12 12 11 12 2 9 2 2 2 12 2 12 2 9 2 2 12 2 12 2
3 9 1 9
51 9 11 11 2 11 9 1 9 2 9 1 12 2 9 2 15 13 9 9 11 2 13 9 1 9 7 9 2 15 9 13 1 9 12 2 12 1 0 9 16 3 11 2 11 11 11 7 0 11 11 2
24 1 15 15 13 13 9 13 2 9 9 2 15 3 13 2 15 13 3 3 3 1 15 2 2
25 9 2 15 13 13 1 0 7 0 9 2 1 9 7 13 15 1 9 2 15 3 13 0 9 2
39 3 1 0 9 9 0 9 13 3 1 15 11 11 13 2 0 9 13 0 9 1 12 0 9 0 1 0 7 0 9 2 9 2 9 7 9 0 9 2
21 0 9 15 4 3 3 13 1 15 2 15 9 2 9 7 9 3 13 1 0 2
16 3 0 15 13 9 1 9 16 0 9 0 0 9 2 2 2
28 9 2 9 11 2 0 12 2 12 12 11 12 2 9 2 2 2 12 2 12 2 9 2 2 12 2 12 2
4 9 2 0 9
3 9 1 9
20 1 0 9 9 15 7 10 9 13 0 9 2 10 9 1 0 7 0 9 2
26 1 9 2 1 15 15 0 9 13 2 13 0 9 0 1 0 9 2 3 13 3 10 9 1 9 2
11 9 9 1 9 13 0 3 1 10 9 2
12 9 13 9 9 7 13 1 9 0 0 9 2
17 9 13 10 9 7 13 9 2 15 4 3 1 9 1 9 13 2
17 16 15 9 13 2 13 0 2 16 15 9 10 9 1 9 13 2
30 16 13 1 9 2 3 9 1 15 3 13 2 16 15 1 9 1 9 13 13 0 9 7 9 1 9 13 3 0 2
5 11 11 2 11 12
14 0 9 0 1 10 9 13 1 0 9 7 0 9 2
20 13 14 9 1 0 0 9 2 7 7 15 2 1 15 15 9 13 16 9 2
3 9 7 9
32 1 0 9 4 13 16 0 0 9 10 9 2 9 13 0 13 1 9 9 15 9 2 1 15 13 0 7 0 9 7 9 2
6 15 3 2 15 3 2
14 1 0 9 13 0 2 1 0 13 15 9 7 9 2
12 15 15 13 9 0 9 0 9 11 11 11 2
2 11 11
26 0 2 15 4 13 1 10 9 13 1 0 9 9 2 13 9 7 10 9 2 13 15 13 11 11 2
15 3 3 13 0 9 1 0 7 13 2 16 15 9 13 2
14 13 4 15 13 2 16 4 15 13 10 9 0 9 2
18 15 15 13 9 7 15 13 13 1 9 7 13 2 10 9 4 13 2
18 13 3 2 4 13 0 2 15 1 10 9 13 3 0 7 0 9 2
54 0 10 9 13 2 16 15 13 1 9 0 9 2 0 9 13 1 12 5 2 9 1 0 9 9 13 2 3 0 9 0 9 7 0 9 2 3 0 9 2 0 9 9 2 0 9 0 9 2 3 0 0 9 2
53 3 15 13 1 0 0 9 9 1 0 9 2 3 13 1 9 9 2 2 3 12 0 9 1 15 2 13 9 9 2 2 3 13 1 0 9 9 2 16 13 15 13 7 13 0 2 10 9 13 7 15 14 2
14 10 9 7 9 4 13 1 10 9 2 13 11 11 2
31 15 13 1 0 9 13 9 1 15 2 15 13 13 15 7 3 2 15 13 13 0 7 3 7 15 13 3 13 1 9 2
18 1 15 9 15 13 0 2 16 13 13 1 0 9 7 9 0 9 2
5 7 13 4 15 2
10 0 9 13 2 13 0 3 13 9 2
16 0 13 7 13 9 9 1 12 7 12 9 7 3 13 9 2
15 9 15 13 13 2 16 0 9 13 15 2 15 15 13 2
14 1 0 9 13 3 0 9 2 15 13 13 0 9 2
20 0 9 13 0 9 2 16 15 15 13 2 3 15 13 7 1 0 9 13 2
17 15 3 3 13 2 3 15 13 0 9 2 15 9 13 1 9 2
32 13 4 13 10 9 2 16 13 13 3 7 1 9 9 2 13 11 11 7 13 2 13 15 2 15 1 15 13 14 1 9 2
10 15 15 15 3 13 2 7 3 13 2
39 13 3 1 9 0 9 2 15 15 13 2 9 13 2 9 10 7 10 9 13 1 9 0 9 2 16 1 0 9 13 9 7 10 9 1 15 4 13 2
15 7 13 15 15 13 7 1 12 9 15 15 0 9 13 2
26 9 2 0 9 0 2 9 2 1 0 9 12 2 12 12 11 2 9 2 12 12 2 9 2 12 12
3 9 2 9
14 9 2 15 1 15 13 0 9 2 3 13 0 9 2
16 9 13 1 9 2 1 15 3 13 9 7 0 9 1 9 2
17 9 9 13 2 16 9 13 9 13 0 9 2 15 9 13 13 2
16 13 3 0 9 9 2 15 13 9 9 7 9 3 9 13 2
28 13 15 9 0 2 7 0 7 0 2 1 9 1 0 1 11 2 3 15 0 13 13 15 2 9 7 9 2
9 11 11 2 9 0 0 9 9 9
1 11
3 1 0 9
15 9 11 11 1 9 7 9 0 9 0 9 2 3 0 2
21 1 12 9 9 9 13 12 5 9 9 1 9 7 9 9 3 3 13 9 9 2
35 9 2 11 11 2 9 2 9 2 0 2 2 0 12 2 12 12 11 2 9 2 2 2 12 2 12 12 2 9 2 2 12 2 12 12
1 11
3 1 0 9
15 11 1 9 9 0 9 2 15 4 13 1 0 0 9 2
4 15 13 11 9
10 9 11 11 13 1 11 9 1 9 9
20 1 10 9 0 9 0 9 9 10 9 11 11 13 9 13 9 1 0 9 2
2 11 11
5 10 9 13 3 2
24 3 13 1 9 1 11 2 15 13 1 0 9 1 9 12 2 15 9 13 3 12 9 9 2
21 3 13 3 9 2 15 15 13 1 9 0 9 9 12 1 9 14 12 9 9 2
21 0 9 13 9 10 9 2 15 13 1 9 9 9 1 0 0 9 1 9 12 2
30 1 9 1 0 9 4 0 12 9 13 1 9 12 1 12 7 1 9 0 9 1 15 2 15 13 9 9 1 11 2
24 9 13 9 0 9 1 11 1 9 14 12 9 9 2 16 1 0 9 13 14 12 9 9 2
4 15 15 13 2
20 0 9 13 2 16 13 1 9 9 12 7 12 13 13 9 9 9 9 9 2
41 9 9 13 1 15 2 15 15 13 2 13 15 9 9 7 9 9 9 9 7 9 11 11 2 15 13 9 9 2 15 10 9 3 13 1 11 9 9 11 11 2
19 0 9 1 9 13 2 16 4 9 13 13 9 9 2 15 0 9 13 2
28 13 3 1 15 2 16 4 15 13 13 3 0 9 1 9 2 3 0 9 2 16 3 9 1 9 7 3 2
20 1 12 2 9 12 4 13 13 13 9 2 15 4 15 13 13 9 0 9 2
18 3 4 13 13 9 1 9 0 0 9 1 9 9 7 9 1 11 2
2 0 9
24 1 15 2 10 9 4 0 9 13 2 15 13 3 9 9 2 3 1 10 9 4 13 13 2
39 0 9 4 13 2 16 4 1 9 0 9 9 13 13 13 0 0 9 2 16 13 9 1 9 0 9 2 3 7 9 9 0 9 2 3 13 11 11 2
29 13 1 10 0 9 2 3 4 15 13 13 9 0 10 0 9 2 15 9 9 4 0 13 0 9 1 10 9 2
23 9 9 0 9 1 9 1 12 9 13 7 9 9 1 9 9 1 9 0 9 1 11 2
39 1 9 10 9 15 15 13 2 16 4 13 13 1 10 9 0 2 7 0 9 15 1 10 9 13 0 9 2 16 4 13 3 3 10 9 10 9 13 2
26 7 13 4 13 9 13 10 9 2 15 4 1 9 10 0 9 13 13 2 7 13 2 13 11 11 2
3 9 13 9
22 9 0 0 9 13 7 9 1 9 9 1 0 9 0 9 0 9 1 10 0 9 2
12 13 3 7 9 9 1 0 9 1 9 12 2
12 10 9 13 7 9 9 2 15 12 9 13 2
19 1 0 9 13 1 9 2 16 13 9 7 9 2 1 0 1 0 9 2
20 0 9 13 9 3 1 9 2 0 9 2 0 9 7 0 9 1 0 9 2
28 16 13 1 0 9 0 7 0 9 2 13 15 13 3 2 16 4 0 9 13 10 9 2 7 9 1 15 2
13 0 9 15 13 13 13 7 13 15 15 13 13 2
29 9 13 2 16 0 9 13 0 0 9 2 15 9 13 13 0 9 1 15 2 15 4 13 13 1 0 9 0 2
6 9 2 15 13 0 2
8 13 15 9 0 0 9 7 9
17 0 9 9 1 9 1 9 0 9 9 12 4 13 12 2 9 2
10 9 13 0 13 1 12 2 9 12 2
2 11 11
33 1 0 9 9 1 9 0 9 2 15 13 0 0 9 11 2 0 9 11 11 2 11 2 0 7 0 9 2 15 13 7 9 2
16 9 4 13 16 9 1 9 2 15 13 0 9 1 0 9 2
13 13 9 13 9 2 0 9 2 9 7 0 9 2
27 0 9 13 0 13 14 1 11 11 2 7 3 1 9 0 9 2 0 9 7 1 15 0 9 1 9 2
44 9 4 13 9 2 1 15 13 11 11 2 10 9 2 11 11 2 9 9 11 2 11 11 2 11 2 9 0 0 9 7 11 11 2 9 9 11 7 0 9 9 0 9 2
26 0 9 9 13 0 13 3 1 12 2 9 2 16 0 9 13 1 9 7 0 9 9 13 1 9 2
8 3 4 13 9 7 0 9 2
41 9 2 11 2 0 9 2 9 2 12 2 9 12 2 12 12 11 2 9 2 2 2 12 2 12 12 2 12 12 2 9 2 2 12 2 12 12 2 12 12 2
4 2 9 13 2
2 0 9
17 0 9 9 9 11 13 10 9 3 0 9 9 2 9 7 9 2
31 3 13 1 0 9 9 1 9 1 0 9 7 9 2 13 15 3 7 7 9 1 0 9 1 0 9 7 1 0 9 2
28 1 9 9 0 0 9 1 0 0 0 11 2 0 9 1 0 9 0 11 2 13 10 9 0 9 1 11 2
37 13 1 9 2 15 1 0 9 13 9 9 7 9 11 2 11 0 9 7 11 0 11 7 1 0 9 0 9 11 1 9 11 7 11 0 11 2
24 0 9 15 1 9 13 13 1 9 9 0 9 1 11 7 1 0 9 1 9 1 10 9 2
24 3 0 2 7 1 10 9 3 0 9 2 13 9 9 2 10 9 15 13 1 11 3 13 2
18 0 9 1 0 13 0 9 1 0 9 1 9 13 0 7 0 9 2
10 9 9 13 9 0 1 9 0 9 2
27 0 13 3 0 9 9 2 9 12 7 12 9 2 9 1 9 7 9 9 7 9 1 0 7 0 9 2
11 0 9 13 1 11 12 9 1 12 9 2
2 11 11
27 9 2 9 9 11 2 0 12 2 12 12 11 12 2 9 2 2 2 12 2 12 12 12 12 2 12 2
2 0 9
26 3 0 9 13 1 15 2 16 9 2 3 3 1 15 2 13 0 9 2 3 7 3 13 1 15 2
14 10 7 0 9 2 9 2 9 9 13 13 3 3 2
19 16 13 0 0 0 9 1 9 7 9 2 3 13 1 10 9 3 0 2
19 15 7 13 13 0 9 1 9 2 7 1 10 9 13 1 9 0 9 2
41 13 4 15 15 7 1 9 0 9 2 0 9 1 0 2 9 2 9 2 3 2 2 9 2 3 13 9 1 2 0 9 2 7 2 0 9 1 9 12 2 2
18 13 1 9 2 15 15 13 16 9 7 13 1 15 0 9 1 12 2
5 13 1 15 13 2
26 2 9 13 9 2 15 9 13 7 13 1 9 2 9 7 9 0 9 0 9 0 10 9 13 9 2
26 2 9 13 7 9 7 9 0 9 1 9 2 9 7 9 0 9 2 16 13 0 10 9 13 9 2
19 0 9 7 13 2 4 2 14 9 1 10 9 9 13 2 0 9 2 2
12 9 0 9 2 9 3 13 13 3 0 9 2
9 1 15 15 3 1 15 3 13 2
31 13 15 3 2 16 1 9 1 0 9 9 13 10 9 2 0 0 9 9 7 9 0 9 12 9 2 0 9 13 9 2
18 9 0 9 13 9 1 9 2 9 7 9 0 9 2 15 13 0 2
21 13 2 16 0 9 13 9 0 7 0 9 2 16 9 9 9 13 9 9 9 2
10 3 9 13 1 9 2 0 9 2 2
25 13 15 3 2 16 13 3 13 2 3 16 9 2 15 15 10 9 13 1 0 9 7 1 9 2
23 13 15 13 14 0 2 7 7 0 9 2 9 2 2 0 9 7 9 2 3 7 3 2
11 9 7 13 13 13 1 9 13 0 9 2
20 9 9 9 15 13 1 0 9 9 2 15 13 7 0 9 2 9 0 13 2
28 3 13 2 13 2 14 15 2 16 10 9 13 0 7 0 2 3 3 13 2 16 9 0 13 0 7 0 2
18 0 9 15 1 15 3 3 13 2 7 3 2 16 15 9 9 13 2
10 1 10 9 7 13 0 9 1 9 2
17 7 13 14 9 9 2 3 15 13 1 10 9 0 9 1 9 2
2 11 11
3 0 9 9
6 7 9 13 1 9 2
5 9 7 1 10 9
12 1 0 9 9 15 1 15 13 1 0 9 2
15 1 11 7 3 13 2 13 9 2 15 13 9 0 9 2
7 13 15 10 9 7 15 2
18 1 9 4 15 13 13 1 0 9 9 1 0 0 9 11 2 11 2
30 0 9 1 0 11 13 0 9 11 13 9 12 9 9 1 9 9 11 11 11 2 16 3 13 9 10 3 0 9 2
3 1 15 13
20 11 15 13 3 0 9 9 9 12 9 11 2 15 13 13 9 1 9 9 2
23 0 9 0 1 0 9 9 3 11 13 1 9 0 11 1 0 9 10 9 11 2 11 2
24 9 11 1 11 13 1 9 2 16 15 13 12 1 0 9 2 3 9 2 13 1 9 2 2
11 3 9 9 13 1 0 9 3 0 9 2
13 0 9 3 13 7 3 1 9 0 9 0 9 2
38 0 9 3 13 9 9 2 16 7 0 7 15 0 9 1 9 13 0 9 9 7 0 9 1 9 3 13 9 9 1 9 0 7 0 9 0 9 2
19 13 1 9 2 16 1 0 15 9 0 9 15 0 9 13 7 1 15 2
20 7 13 0 13 2 15 13 0 0 9 9 0 9 2 1 9 1 0 9 2
1 9
11 13 15 1 0 9 2 15 13 0 9 2
9 9 0 9 13 9 9 0 9 2
9 13 1 12 0 9 13 10 9 2
25 2 13 1 9 0 2 0 7 0 9 2 15 13 0 7 3 0 9 2 14 0 7 0 9 2
11 2 10 9 13 1 0 0 9 3 0 2
15 2 9 13 9 1 9 10 9 7 10 9 0 9 13 2
40 1 9 0 9 2 15 4 13 4 13 1 0 9 2 13 13 3 9 0 7 0 2 0 9 2 9 7 9 0 9 2 0 9 2 9 2 9 9 3 2
19 1 9 0 9 0 0 9 13 0 13 0 9 2 0 9 2 9 3 2
35 1 9 0 9 2 15 13 13 16 0 9 15 13 13 0 9 2 0 9 2 9 2 9 0 9 2 0 7 0 9 2 0 9 3 2
2 9 9
14 0 2 15 13 0 9 13 1 0 9 2 13 9 2
43 15 3 13 13 2 10 9 13 13 16 9 13 7 3 7 13 2 7 15 3 13 3 2 13 2 2 16 15 3 0 9 7 9 13 1 0 0 9 0 7 3 0 2
5 11 11 2 0 9
1 9
3 9 1 9
37 9 13 10 9 1 9 3 1 9 2 16 13 15 0 0 9 2 0 9 7 9 2 13 1 0 9 7 0 0 9 2 9 2 7 0 9 2
15 13 15 2 1 15 15 13 1 9 15 1 10 9 13 2
4 11 11 2 11
13 0 9 13 10 9 1 0 9 1 9 3 3 2
7 13 7 1 9 9 9 2
15 0 9 13 0 1 10 9 13 0 9 7 1 9 9 2
16 9 3 13 13 3 0 2 16 4 10 9 13 13 9 9 2
7 9 3 13 3 13 3 2
22 1 10 9 2 13 2 14 15 1 9 1 0 9 2 13 13 1 9 9 7 9 2
14 0 9 13 13 7 0 2 7 1 9 16 0 9 2
26 1 9 1 15 13 13 1 9 2 16 1 15 13 0 9 3 3 13 2 1 0 9 7 0 9 2
6 13 3 1 9 9 2
25 7 9 9 13 14 0 2 13 0 9 2 3 9 7 1 9 13 9 7 13 1 15 0 9 2
7 0 1 9 13 0 9 2
18 13 15 1 9 1 9 9 2 13 0 7 1 9 1 9 7 9 2
22 13 2 14 1 9 15 9 2 9 13 2 13 15 2 9 2 2 2 7 13 15 2
11 9 13 0 1 9 7 9 15 3 13 2
30 0 9 13 2 16 7 0 9 13 13 0 9 2 15 13 14 12 5 0 9 2 15 13 0 9 9 0 1 9 2
14 1 9 9 0 9 13 3 1 9 9 7 10 9 2
20 16 10 12 9 4 13 2 9 13 0 1 9 7 0 0 9 15 3 13 2
9 1 9 9 13 3 0 3 13 2
5 13 13 3 0 2
25 2 0 9 9 2 16 4 15 13 3 3 1 0 9 2 7 1 0 2 15 13 7 0 9 2
11 16 9 13 13 9 11 11 11 2 11 2
12 2 9 0 9 2 15 13 0 9 1 9 2
9 16 9 1 9 13 3 0 9 2
5 2 15 13 9 2
38 0 2 3 16 0 7 0 9 13 13 1 9 11 1 0 9 7 9 1 10 9 13 9 11 2 10 9 13 9 1 9 14 0 9 3 0 9 2
4 2 9 9 2
40 13 0 13 15 9 1 10 10 9 2 13 2 16 13 9 1 9 2 13 15 9 15 0 9 2 7 7 3 15 13 0 9 2 15 13 0 9 1 0 2
7 10 0 9 13 3 0 2
2 11 11
20 9 2 11 12 2 12 12 11 12 2 9 2 5 9 2 2 12 2 12 2
1 9
4 9 1 12 9
9 9 1 9 9 13 3 12 9 9
18 7 16 0 9 0 9 3 3 13 2 1 9 0 9 3 3 13 2
9 13 2 16 10 9 0 9 13 2
16 13 15 7 15 9 2 1 15 4 13 2 16 15 4 13 2
20 1 15 2 3 13 9 14 0 2 9 13 1 11 11 2 9 9 0 9 2
5 11 11 2 11 11
20 2 9 9 0 0 9 3 13 10 9 2 7 15 15 3 13 1 10 9 2
3 13 13 2
20 9 9 0 9 13 9 2 3 3 13 9 9 2 15 13 1 9 1 9 2
37 13 3 1 3 12 9 9 9 1 9 9 2 7 3 15 13 2 14 1 0 9 2 14 16 9 0 2 7 3 0 2 7 3 16 9 0 2
6 2 15 15 13 13 2
9 16 0 9 13 0 2 13 0 2
13 7 13 9 1 12 9 13 1 9 0 9 0 2
5 13 13 9 9 2
22 9 1 9 7 3 13 7 10 0 9 2 13 9 10 9 1 9 9 1 0 9 2
14 2 1 15 15 3 3 13 1 0 9 1 9 12 2
19 3 1 15 13 12 9 9 2 7 3 2 7 1 9 2 9 7 3 2
12 15 2 16 3 13 0 9 2 13 1 0 2
11 9 7 13 2 16 15 0 9 3 13 2
37 9 15 1 9 7 3 2 16 12 9 9 15 13 2 13 15 1 9 3 13 7 3 3 13 15 2 15 1 10 3 0 9 3 13 16 0 2
24 2 4 13 9 9 7 1 9 2 3 15 13 9 14 3 2 16 10 9 13 3 0 9 2
10 10 9 1 9 9 4 13 1 0 2
12 7 3 13 3 9 2 15 13 7 0 9 2
11 3 9 15 13 7 9 10 9 13 9 2
8 3 15 13 9 13 9 3 2
18 15 4 13 1 0 2 3 1 0 9 2 7 3 10 9 3 13 2
13 9 0 9 13 13 9 2 7 13 13 0 9 2
24 3 15 13 2 16 4 15 1 10 9 13 0 1 11 13 2 3 15 3 13 1 10 9 2
7 2 3 10 9 13 3 2
17 1 9 2 3 15 13 0 9 2 1 15 7 3 4 15 13 2
16 9 13 14 15 10 2 7 15 15 1 15 0 13 3 13 2
15 1 10 0 9 13 7 9 7 3 1 10 9 13 9 2
32 1 10 9 1 10 0 9 10 9 13 9 2 15 13 2 7 9 2 16 0 9 0 9 2 4 1 15 1 0 9 13 2
19 2 3 7 3 12 9 9 9 2 15 13 9 1 9 2 13 3 9 2
8 15 13 9 1 9 0 9 2
19 16 9 13 2 7 13 14 1 12 0 0 9 2 13 9 9 10 9 2
19 13 9 2 15 13 3 14 12 9 2 7 13 0 9 1 9 0 9 2
6 4 15 13 1 12 2
24 2 3 13 9 2 16 4 3 13 1 9 1 9 9 7 13 2 3 15 13 1 0 9 2
5 3 1 15 0 2
40 3 13 3 13 2 16 9 9 13 3 0 2 3 16 15 9 13 1 9 9 2 15 15 15 13 3 13 2 13 9 2 1 15 15 13 9 2 7 3 2
19 7 3 13 9 1 9 2 3 13 3 13 9 13 9 9 1 0 9 2
36 2 13 15 3 1 9 2 16 9 7 0 9 13 15 2 15 13 3 0 9 2 7 3 2 16 13 13 9 7 1 9 2 13 1 9 2
39 13 1 9 9 2 3 9 2 15 15 13 0 9 2 1 15 13 9 13 7 15 1 15 2 15 13 7 13 14 3 1 0 2 0 9 1 0 9 2
6 15 13 3 9 11 2
28 0 13 10 9 1 0 9 2 3 15 15 13 13 9 9 7 13 9 3 1 3 0 7 3 0 0 9 2
26 3 4 10 9 13 3 1 9 1 9 2 16 15 1 10 9 3 13 2 16 1 0 9 3 13 2
24 9 13 2 7 16 13 0 7 0 9 13 2 3 9 13 4 2 7 13 15 0 1 9 2
8 2 10 9 15 3 13 3 2
7 1 0 12 9 9 9 2
11 3 12 9 15 15 3 13 1 0 9 2
14 3 13 0 9 2 9 1 9 2 9 7 0 9 2
13 2 1 9 2 15 13 1 9 2 15 3 13 2
27 16 13 0 1 9 2 16 15 3 0 9 2 0 9 7 9 1 9 0 9 3 3 3 13 1 9 2
28 13 4 3 13 0 9 1 9 2 15 13 15 0 1 10 0 0 9 2 7 3 15 13 9 7 13 9 2
9 2 4 1 9 13 7 10 9 2
24 14 2 7 15 1 9 2 16 4 9 13 13 1 0 9 1 0 9 2 0 1 0 9 2
10 0 15 13 1 9 2 3 13 9 2
12 2 7 1 0 9 13 3 9 9 9 9 2
16 15 13 3 9 2 0 1 0 9 2 3 1 9 1 9 2
32 13 15 0 9 2 12 13 9 2 1 0 9 0 12 15 13 9 2 7 13 1 9 7 3 0 12 9 0 15 3 13 2
13 2 3 15 13 1 9 9 13 1 3 0 9 2
11 13 2 16 4 13 13 1 9 9 12 2
13 13 3 9 7 9 2 7 15 3 13 13 9 2
9 15 13 13 9 3 1 9 9 2
24 2 0 9 1 9 9 1 10 9 0 11 13 9 9 9 7 9 2 3 12 7 15 9 2
26 13 15 3 1 15 1 9 2 16 1 0 9 13 1 10 9 9 9 2 16 4 15 3 3 13 2
7 10 9 13 3 0 9 2
20 15 13 7 11 2 7 11 2 3 13 1 0 9 9 0 9 1 9 0 2
21 1 15 13 3 1 0 2 16 0 9 2 7 1 15 13 9 9 1 0 9 2
34 16 1 15 15 9 13 3 16 15 13 3 2 3 15 3 3 13 13 9 2 3 15 10 9 2 7 0 9 1 9 13 3 9 2
14 13 4 7 3 1 9 2 15 4 13 9 1 9 2
3 9 1 9
11 13 15 13 9 2 3 15 10 9 13 9
3 9 1 9
6 0 9 13 0 0 9
10 0 9 13 3 3 0 7 0 9 2
19 10 9 9 2 14 13 1 0 2 0 9 7 0 9 2 13 0 9 2
17 3 12 12 9 0 9 13 1 9 0 7 0 9 7 9 9 2
20 1 9 4 7 13 13 3 0 9 0 0 9 2 0 9 7 9 0 9 2
3 1 0 9
12 0 9 13 1 10 9 3 13 9 0 9 2
14 10 9 3 13 9 9 11 12 3 16 9 9 9 2
17 1 0 2 0 9 13 9 9 2 3 13 7 0 9 0 9 2
10 1 9 9 3 9 13 9 1 11 2
8 0 9 13 0 9 0 9 2
11 10 9 13 9 13 2 7 13 15 9 2
20 3 4 9 0 9 1 12 9 13 12 9 9 2 7 13 13 14 12 9 2
17 7 1 0 9 13 1 0 9 2 13 0 9 0 9 11 11 2
14 0 12 9 9 15 13 9 9 7 9 9 1 9 2
3 9 1 9
8 9 13 7 0 9 1 9 2
13 3 1 11 15 13 0 9 1 9 13 0 9 2
20 0 9 13 0 9 1 0 0 9 1 11 2 11 7 13 9 0 0 9 2
24 13 7 13 3 1 9 7 9 9 1 0 9 2 7 3 1 9 9 1 9 9 2 9 2
23 10 9 3 13 9 1 10 0 9 2 15 13 9 0 9 1 10 9 7 1 0 9 2
31 0 9 13 2 16 16 9 1 0 9 3 13 1 0 9 0 9 13 2 0 9 3 13 9 3 1 0 7 0 9 2
10 0 9 13 13 13 0 9 15 9 2
2 9 11
10 0 9 13 9 3 1 9 0 9 2
10 13 13 11 0 9 1 9 0 9 2
26 1 10 9 13 0 0 9 12 9 2 11 13 12 9 2 2 15 4 13 0 9 7 1 9 11 2
11 0 9 13 3 13 3 0 9 0 9 2
14 9 15 7 13 2 16 0 9 13 1 10 0 9 2
18 7 13 13 3 0 0 9 2 15 1 9 13 7 0 9 2 9 2
6 13 13 1 0 9 2
28 13 15 14 0 9 2 7 3 9 0 9 2 15 4 13 9 1 9 7 9 0 0 9 2 13 11 11 2
35 9 2 0 9 2 0 2 9 2 2 0 12 2 12 12 11 12 2 9 2 2 2 12 2 12 12 2 9 2 2 12 2 12 12 2
8 9 1 0 2 9 2 0 9
8 9 2 1 9 2 9 2 12
8 9 2 1 9 2 9 2 12
2 9 12
3 13 15 9
7 9 13 13 1 15 9 2
3 9 9 9
16 15 13 15 2 16 9 0 7 0 9 1 0 11 3 13 2
10 9 1 10 9 1 9 12 3 13 2
15 1 9 9 11 2 11 2 11 1 9 12 13 15 3 2
14 0 9 13 1 12 9 9 1 12 9 7 3 13 2
15 1 0 9 9 13 9 0 9 3 1 9 0 0 9 2
10 1 9 2 9 2 9 2 9 9 2
5 0 9 3 13 2
2 9 9
11 9 3 13 9 10 9 1 9 9 9 2
7 0 9 13 13 7 3 2
22 9 9 13 9 9 9 9 1 9 3 1 9 2 1 0 9 2 9 7 1 9 2
9 13 9 13 7 0 9 9 9 2
18 9 1 12 12 15 13 2 13 11 11 2 2 1 9 2 2 9 2
6 15 13 1 9 0 2
14 9 0 9 13 15 7 9 9 9 13 15 0 9 2
13 15 15 1 0 9 13 1 12 9 7 13 0 2
33 9 13 0 13 7 9 1 12 9 0 2 13 2 14 1 9 1 0 9 2 3 1 9 9 1 9 2 15 13 0 1 9 2
6 7 15 13 14 9 2
13 9 7 3 13 9 1 9 14 12 9 5 9 2
14 13 1 0 9 7 9 9 13 3 2 16 13 9 2
14 13 9 2 16 1 9 13 9 7 13 15 0 9 2
2 13 9
14 0 9 13 2 16 1 9 0 9 9 13 9 9 2
4 3 13 15 2
16 9 9 13 1 12 9 12 5 2 3 4 13 13 12 5 2
16 9 15 13 1 0 9 2 15 15 13 0 9 1 0 9 2
13 0 9 13 13 0 0 9 7 1 10 9 13 2
12 1 0 9 13 1 11 12 7 3 9 3 2
9 0 9 13 13 9 9 1 11 2
12 9 3 13 7 13 0 13 1 9 0 9 2
8 9 7 13 9 7 9 13 2
22 0 9 13 9 9 9 7 9 2 15 15 13 1 12 2 12 1 0 12 2 12 2
9 3 1 0 9 13 3 12 9 2
19 3 13 12 9 2 15 13 3 3 12 9 3 2 7 4 3 3 13 2
3 9 1 9
9 3 13 15 4 2 13 9 11 2
6 0 9 13 3 0 2
10 7 16 4 3 9 13 2 15 3 2
14 9 1 9 7 9 12 13 1 9 12 9 1 9 2
9 9 13 0 2 16 15 3 13 2
6 0 9 13 12 9 2
10 9 13 7 15 2 16 13 9 9 2
9 1 9 13 3 9 1 0 9 2
8 0 1 15 13 13 0 9 2
12 16 15 15 15 13 2 13 1 12 5 9 2
19 9 7 13 9 2 0 9 2 7 1 10 9 13 3 13 0 0 9 2
3 9 16 9
11 3 3 9 1 12 9 13 1 0 9 2
10 9 7 9 9 15 3 13 7 13 2
9 9 13 1 9 13 7 9 13 2
17 1 0 0 9 13 9 13 13 9 1 0 9 1 12 9 9 2
6 13 15 9 3 0 2
10 7 9 13 3 0 2 13 9 11 2
14 1 0 9 13 9 2 7 16 13 1 9 3 0 2
13 3 1 9 1 9 9 9 13 10 9 1 11 2
6 1 9 15 13 9 2
10 3 13 7 13 2 7 3 3 13 2
12 12 9 13 0 13 2 16 13 9 13 9 2
18 13 0 13 9 9 7 0 9 2 1 15 9 4 15 13 0 9 2
12 3 15 12 9 13 3 9 9 7 13 3 2
40 9 2 11 2 11 2 11 2 9 2 9 2 0 2 2 0 12 2 12 12 11 2 9 2 2 2 12 2 12 12 12 2 9 2 2 12 2 12 12 12
15 9 2 0 9 2 0 9 2 15 9 1 11 13 3 2
5 13 9 9 2 12
22 9 15 13 13 2 13 1 9 3 0 0 0 9 1 9 11 11 2 9 11 11 2
16 1 9 9 11 13 0 11 0 9 1 9 12 0 0 9 2
13 9 3 13 0 9 9 2 3 3 13 0 9 2
6 0 9 3 13 0 2
11 13 2 14 15 1 9 9 2 13 9 2
6 13 12 9 1 9 2
13 2 1 0 0 9 13 2 0 9 2 2 2 2
4 3 15 9 2
4 9 11 11 2
4 9 2 10 9
3 11 11 13
14 0 11 2 15 13 11 11 2 15 3 13 3 13 2
13 1 0 9 1 0 9 15 13 15 0 2 9 2
3 13 15 2
7 0 9 13 11 9 11 2
2 11 11
15 0 9 1 0 9 13 14 3 0 2 3 1 0 9 2
22 1 9 13 9 1 9 9 2 9 13 2 13 15 3 9 0 9 2 9 7 9 2
12 0 9 1 0 0 9 15 13 1 0 9 2
20 13 15 2 16 15 13 9 2 15 13 0 0 9 13 1 0 2 0 9 2
17 0 9 11 3 13 0 9 1 9 1 9 9 9 11 0 9 2
15 2 9 2 15 13 3 2 16 13 12 2 9 2 13 2
14 1 0 9 0 9 7 13 1 0 9 3 0 9 2
24 9 9 13 0 9 11 9 11 11 15 9 9 11 1 0 9 1 9 1 0 7 0 9 2
24 3 16 9 0 7 0 9 4 13 1 9 0 9 7 1 10 9 15 13 7 0 0 9 2
14 1 9 0 9 13 9 7 0 9 0 9 11 11 2
13 15 13 1 11 9 1 9 0 9 1 9 9 2
8 13 0 9 1 9 0 9 2
40 3 13 13 7 13 2 16 0 9 7 3 9 11 11 13 16 12 1 0 9 11 7 7 3 2 16 15 16 15 9 1 9 13 9 7 13 1 9 0 2
7 12 7 3 3 13 0 2
38 9 1 9 1 0 0 9 2 9 0 9 2 9 0 9 1 0 9 7 3 9 1 0 0 9 1 9 0 9 13 0 9 2 15 4 13 13 2
5 9 1 11 15 13
11 1 11 13 0 9 7 9 1 9 0 9
21 9 0 2 7 1 0 9 2 0 7 0 9 0 11 2 13 3 9 0 9 2
13 3 1 9 3 0 9 13 10 9 13 0 9 2
11 9 0 9 15 13 0 3 1 9 12 2
20 9 15 9 13 9 1 9 9 1 0 9 2 9 13 9 2 15 4 13 2
11 11 13 1 9 3 0 2 3 15 13 2
7 9 1 0 11 15 13 2
3 9 1 9
19 1 0 0 9 1 9 13 0 9 1 0 9 0 7 3 15 0 9 2
11 13 1 15 0 12 9 9 1 0 9 2
6 15 13 9 1 11 2
27 1 9 9 2 9 0 9 1 9 9 7 9 0 0 9 4 13 10 0 9 1 9 0 9 1 11 2
8 1 9 9 15 9 3 13 2
19 4 13 9 0 9 2 15 9 9 0 7 0 9 1 10 9 3 13 2
8 13 15 3 0 9 1 11 2
29 0 9 1 9 1 9 13 3 9 0 9 2 3 9 2 7 0 0 9 0 9 0 9 1 0 7 0 9 2
2 3 13
12 9 13 3 12 1 9 2 15 13 0 9 2
9 13 3 7 0 9 7 0 9 2
10 1 0 9 3 13 9 9 0 9 2
19 1 9 0 9 7 4 13 14 10 9 2 10 9 13 13 1 0 9 2
26 1 0 9 13 1 11 12 5 9 3 16 12 9 7 3 14 12 5 13 1 10 9 1 12 9 2
17 1 9 13 3 9 1 0 9 2 15 13 13 3 16 0 9 2
12 0 9 0 9 13 3 1 0 9 7 9 2
7 3 3 0 9 13 3 2
14 9 3 13 9 1 11 2 15 15 13 1 9 0 2
12 3 0 9 9 13 1 11 3 12 7 3 2
25 0 9 13 9 9 1 11 7 11 2 15 13 1 9 13 7 13 1 11 1 12 7 12 9 2
2 9 9
16 9 9 1 0 7 0 11 13 1 9 0 9 9 0 9 2
15 3 13 0 0 9 2 3 9 0 0 9 2 9 3 2
10 1 0 9 15 13 13 7 9 9 2
13 1 9 13 1 9 1 0 9 1 11 12 9 2
15 13 3 14 12 0 0 9 2 3 1 9 7 0 9 2
10 0 12 9 13 1 0 9 0 9 2
2 0 9
13 11 13 13 9 9 1 0 9 2 9 7 9 2
22 3 13 0 13 0 0 9 2 1 9 0 1 0 9 2 9 9 2 0 9 3 2
10 3 15 1 9 10 9 15 3 13 2
23 13 15 13 7 15 2 16 3 13 0 9 1 9 9 9 2 15 15 10 9 3 13 2
16 13 15 13 0 0 9 1 9 0 9 2 15 4 13 9 2
29 10 9 9 0 9 4 15 13 1 9 9 2 1 9 7 9 9 7 9 0 9 2 9 2 9 7 0 9 2
9 9 13 13 9 9 1 10 9 2
3 3 13 9
19 9 9 13 2 16 1 0 12 9 15 9 1 9 13 3 1 12 5 2
10 9 0 9 1 11 7 13 0 9 2
19 1 0 9 11 13 0 0 9 2 0 9 2 0 0 9 1 0 9 2
22 13 15 0 3 13 3 1 9 9 2 9 7 9 2 9 13 1 9 7 9 9 2
8 3 7 1 9 9 13 9 2
6 0 0 9 13 0 2
13 13 15 9 1 0 2 15 15 1 0 9 13 2
10 9 9 9 3 13 13 7 9 9 2
13 3 3 9 0 9 9 0 9 0 9 3 13 2
16 0 9 9 1 9 13 13 14 3 2 16 15 13 0 9 2
16 1 10 9 3 13 0 9 2 15 15 4 13 3 1 9 2
2 11 0
12 9 1 0 9 1 11 2 9 2 0 2 2
8 9 1 9 2 0 0 9 2
13 13 0 9 1 9 2 15 13 0 7 0 9 2
3 9 1 9
9 1 0 9 11 13 2 9 2 9
30 1 0 9 2 15 13 11 2 15 15 13 13 1 10 9 7 9 0 9 2 13 15 0 9 1 11 1 12 9 2
18 0 9 0 9 13 9 11 12 9 11 11 11 1 3 9 12 9 2
19 13 7 13 7 0 1 9 2 0 9 2 0 0 9 7 0 0 9 2
18 15 15 13 13 1 9 0 9 11 2 15 1 0 9 10 9 13 2
18 3 13 3 13 9 1 9 7 9 13 3 0 1 10 9 7 9 2
34 16 15 0 9 13 2 13 15 7 3 10 9 7 9 2 7 13 10 9 2 3 15 13 0 9 1 10 0 0 9 1 0 9 2
9 13 2 16 1 11 15 9 13 2
3 3 0 9
7 0 9 13 0 9 7 9
17 1 10 9 15 1 9 12 2 9 0 9 13 0 9 0 9 2
15 1 9 9 2 15 4 13 1 9 2 13 12 0 9 2
33 9 7 0 9 9 13 2 16 4 7 1 0 9 4 10 9 13 7 13 9 2 0 9 2 9 9 2 0 9 3 2 2 2
11 10 9 7 13 13 2 3 9 0 9 2
22 13 15 7 9 1 0 11 2 3 15 15 13 13 9 9 7 9 0 7 0 9 2
3 14 9 3
23 9 13 1 12 2 9 0 9 9 1 3 12 9 9 2 15 13 3 12 10 0 9 2
15 0 9 13 3 1 9 9 2 15 13 3 1 9 9 2
24 9 13 3 13 12 0 7 0 9 2 0 11 11 1 9 12 9 9 2 7 0 0 9 2
6 1 9 9 15 13 2
19 9 15 13 12 9 1 0 0 9 9 2 0 1 12 2 9 1 9 2
14 1 0 7 0 9 13 3 1 0 9 1 0 9 2
34 9 0 9 15 1 9 12 13 1 9 12 1 3 16 9 7 10 0 9 9 9 3 2 9 2 0 9 2 0 9 3 2 2 2
14 1 9 1 0 9 7 13 10 9 3 0 7 0 2
2 0 9
19 16 9 0 9 9 13 1 3 0 9 2 3 0 7 0 13 0 9 2
22 1 0 9 13 1 0 9 1 9 9 12 0 9 2 1 0 0 9 1 9 12 2
15 9 0 9 15 3 13 7 13 9 9 12 3 12 12 2
20 0 0 9 1 9 0 9 13 12 9 2 15 13 1 0 9 9 1 9 2
22 0 9 9 13 3 9 9 2 7 1 15 15 0 9 13 0 0 9 7 0 9 2
22 7 4 13 0 9 0 1 9 0 0 9 2 15 15 13 9 3 1 12 9 9 2
25 1 15 4 1 9 12 13 13 14 12 0 9 1 12 9 2 3 12 9 9 4 13 13 9 2
25 1 9 1 0 9 13 3 1 0 9 2 1 9 12 13 0 9 0 9 12 2 12 9 2 2
10 1 0 9 13 9 9 1 0 9 2
2 0 9
14 1 9 7 9 15 1 12 2 9 13 0 9 9 2
19 13 1 9 1 0 2 0 2 9 1 0 9 7 3 1 3 0 9 2
21 15 4 15 13 1 10 9 13 7 0 9 9 2 9 2 7 15 7 9 9 2
33 1 11 13 7 0 13 1 9 2 16 9 4 1 9 9 3 13 2 7 3 0 9 0 9 4 13 3 1 9 9 7 9 2
9 7 9 9 13 1 10 9 13 2
25 1 0 9 13 3 0 9 16 1 9 2 0 9 15 13 7 13 13 1 0 9 7 9 9 2
21 1 12 2 9 13 7 9 0 9 11 2 15 4 3 13 3 1 12 2 9 2
13 3 1 11 15 3 13 1 9 0 0 0 9 2
22 10 9 2 15 13 3 0 9 9 1 9 2 13 0 9 7 4 1 15 13 9 2
3 11 11 2
2 11 11
31 9 2 0 0 9 2 11 12 2 12 12 11 12 2 9 2 2 12 2 12 12 2 9 2 2 12 2 12 12 12 2
11 15 13 11 1 12 9 9 2 1 9 2
3 0 11 2
19 2 9 9 2 9 2 2 2 9 7 9 2 2 13 1 9 12 2 2
5 1 9 4 15 13
9 11 13 10 9 1 0 9 7 9
21 3 2 16 13 1 9 12 0 9 11 2 13 11 11 1 9 1 12 9 9 2
12 9 3 13 12 9 9 7 9 13 12 9 2
33 3 13 12 9 0 1 9 1 11 3 12 9 2 0 9 13 3 1 12 9 9 7 9 1 15 12 9 13 1 9 12 9 2
15 10 9 4 13 0 1 0 9 7 1 0 9 12 9 2
2 11 11
7 16 0 13 9 12 9 2
14 0 13 9 10 0 9 2 16 4 13 3 0 9 2
27 0 13 9 10 0 9 2 15 4 1 9 0 9 13 13 3 0 9 1 15 9 9 7 13 3 9 2
2 12 9
14 11 13 1 9 1 9 1 9 10 12 9 0 9 2
11 9 9 2 9 2 0 9 7 0 9 2
5 15 13 13 0 2
9 7 9 13 9 1 0 0 9 2
22 13 1 15 7 0 9 2 7 1 9 9 0 9 2 9 1 0 9 2 0 9 2
13 1 12 9 13 0 0 11 2 0 9 0 11 2
8 0 13 1 12 7 12 9 2
19 11 13 0 9 0 9 1 9 1 9 11 2 16 0 13 0 0 9 2
16 11 13 9 0 15 1 9 0 0 7 0 9 2 0 9 2
10 3 13 16 0 9 0 1 0 9 2
22 11 1 0 11 15 13 1 9 7 9 0 7 0 9 2 1 0 13 0 0 9 2
12 11 1 11 15 13 1 9 7 9 0 9 2
12 1 0 0 9 1 11 1 15 13 0 9 2
8 11 11 13 9 9 1 11 2
17 7 11 13 1 15 9 7 0 0 9 2 0 9 7 0 9 2
15 3 4 13 13 0 9 1 11 7 11 0 15 0 9 2
21 15 9 13 0 2 13 1 15 1 0 9 2 13 15 3 1 9 0 0 9 2
12 0 9 13 0 9 2 15 1 15 13 11 2
17 1 9 11 15 13 3 3 3 2 16 9 4 13 1 10 9 2
30 1 15 15 13 3 3 7 9 1 9 2 9 7 3 2 16 13 0 3 13 9 9 0 9 7 3 13 0 9 2
4 1 9 0 11
13 1 11 3 13 1 0 9 0 9 1 9 9 2
10 15 15 7 13 2 16 13 0 9 2
11 7 11 11 13 9 9 3 1 0 9 2
23 13 0 9 2 1 9 15 1 15 13 1 0 9 7 3 15 13 10 9 1 9 9 2
5 3 13 9 11 2
14 13 13 9 3 12 7 3 3 15 13 1 10 9 2
17 3 13 0 13 0 9 2 0 9 2 0 0 9 1 10 9 2
7 0 13 1 9 0 9 2
6 13 9 9 1 9 2
14 16 15 9 3 13 2 13 15 11 13 7 0 9 2
21 3 15 13 1 0 9 11 7 15 13 9 1 10 9 1 10 0 7 0 9 2
14 14 15 9 13 13 2 16 15 13 13 13 1 9 2
11 3 3 15 7 1 15 10 9 13 13 2
19 7 11 11 15 1 0 9 0 9 13 13 0 9 9 1 9 1 11 2
36 9 2 11 2 9 2 9 2 0 2 2 0 12 2 12 12 11 12 2 9 2 2 2 12 2 12 12 2 9 2 2 12 2 12 12 2
4 9 1 9 2
11 9 13 0 2 1 0 9 15 7 13 2
3 16 3 13
7 0 9 13 1 9 9 2
6 9 1 9 1 0 9
19 1 0 9 4 13 0 9 9 7 0 9 1 0 0 9 1 0 9 2
19 3 1 0 9 4 13 0 9 2 3 13 9 1 9 1 9 7 9 2
11 13 1 10 9 2 16 13 9 1 9 2
23 1 0 9 9 1 11 2 11 7 11 4 3 13 2 16 4 13 1 10 0 0 9 2
18 9 13 0 2 1 0 9 7 9 1 9 9 14 1 0 0 9 2
3 9 1 9
34 1 9 3 15 2 16 15 1 11 13 1 0 9 7 0 9 2 15 15 13 9 1 0 9 2 15 3 2 13 1 9 9 12 2
26 1 9 9 13 3 0 9 2 3 0 9 2 13 11 2 11 11 2 9 9 11 2 1 9 2 2
12 0 9 13 0 9 1 0 9 9 2 13 2
26 1 0 9 4 15 15 13 13 9 9 2 3 1 0 9 11 13 1 0 12 9 1 12 9 9 2
22 1 11 7 0 9 13 1 9 0 9 2 9 7 0 9 3 3 1 0 9 9 2
17 1 9 15 13 0 9 7 3 0 9 13 9 1 9 3 0 2
10 9 1 9 15 13 1 0 9 3 2
5 1 9 15 13 13
13 1 9 2 15 0 9 13 2 15 13 11 0 2
10 3 15 13 0 9 0 9 7 9 2
21 11 13 10 0 0 9 2 7 15 13 13 0 7 0 9 0 9 7 9 9 2
24 1 11 15 1 9 13 3 0 0 9 2 15 13 9 9 7 1 0 9 7 0 9 0 2
23 1 9 9 13 0 9 2 1 0 9 13 0 0 9 9 2 10 0 9 13 0 9 2
25 13 15 0 9 1 9 0 9 0 2 11 1 9 2 13 15 1 0 9 7 1 0 0 9 2
18 9 2 9 2 9 7 9 1 9 15 13 1 9 0 9 9 9 2
7 1 9 3 13 11 11 2
9 9 9 13 1 9 1 0 9 2
16 9 9 2 15 13 13 0 9 2 3 13 0 9 1 9 2
12 1 9 9 1 9 13 13 9 9 0 9 2
10 1 9 0 9 13 0 9 7 9 2
10 1 0 15 13 9 13 0 0 9 2
20 1 0 9 13 9 9 9 2 9 7 9 2 15 13 13 1 0 0 9 2
25 9 9 15 13 13 0 9 1 0 9 9 2 16 3 1 0 9 13 9 9 9 7 0 9 2
9 9 1 9 2 0 9 1 11 2
8 1 9 13 3 0 0 9 2
4 9 14 12 9
8 0 9 9 9 1 9 1 11
37 15 13 1 9 0 9 1 0 9 0 0 9 11 2 15 15 1 0 13 7 1 9 9 0 2 3 0 9 1 0 9 1 0 9 1 11 2
23 10 9 3 13 9 9 11 9 12 9 1 9 9 9 0 9 1 12 0 9 1 11 2
2 11 11
9 9 11 13 0 9 1 0 9 2
22 3 15 13 9 9 9 9 9 9 11 11 11 2 9 4 13 1 9 0 9 9 2
1 9
49 9 13 13 1 0 0 7 0 9 1 9 9 1 12 9 1 0 7 0 9 1 9 0 9 2 9 2 9 2 9 2 0 9 7 0 9 2 0 9 7 9 2 9 1 9 7 0 9 2
2 0 9
11 9 4 13 1 0 9 3 1 12 9 2
6 9 9 13 7 13 2
10 12 9 15 0 9 13 13 3 3 2
41 1 9 13 4 13 0 9 2 9 1 0 9 2 9 9 1 0 9 2 0 9 0 9 2 9 0 1 0 9 7 9 1 0 9 2 9 2 9 7 3 2
15 1 9 0 7 13 4 13 9 0 1 9 7 9 9 2
14 9 9 1 0 9 1 12 9 13 12 9 1 9 2
28 11 7 10 9 13 3 9 2 15 4 13 1 0 9 2 0 9 2 0 9 9 2 0 9 7 0 2 2
2 0 9
16 1 0 9 7 9 0 13 13 1 9 9 9 0 0 9 2
13 9 2 11 11 11 2 12 2 2 12 2 12 2
27 2 9 13 13 1 0 9 2 0 9 2 9 2 9 1 9 2 0 9 2 0 9 7 0 9 2 2
10 11 11 2 12 2 2 12 2 12 2
15 2 9 9 13 9 7 0 9 1 9 1 0 9 2 2
11 11 11 1 11 2 12 2 2 12 12 2
18 2 13 15 4 9 1 0 2 0 7 0 9 2 0 9 7 9 2
21 1 9 10 9 15 13 9 1 9 11 2 15 13 13 1 9 9 1 9 2 2
8 11 11 1 11 2 9 12 2
40 2 9 15 13 1 0 9 2 9 2 0 9 2 9 2 0 9 2 9 2 9 1 9 2 0 7 0 9 2 9 2 9 2 0 9 2 0 9 2 2
19 9 9 1 9 1 0 9 13 1 9 1 9 9 11 7 1 9 11 2
20 0 9 3 1 0 9 13 3 13 3 1 12 2 9 12 1 9 9 11 2
17 9 4 13 1 0 9 1 11 11 7 1 9 4 0 9 13 2
19 9 2 9 9 11 2 9 9 9 2 0 9 12 2 12 12 11 12 2
36 7 2 9 11 2 1 11 12 2 0 2 9 2 9 2 12 2 12 12 11 12 2 9 2 2 2 12 2 12 2 9 2 12 2 12 2
5 2 9 1 9 2
2 9 9
27 3 13 13 1 9 9 2 15 4 13 0 0 9 1 9 0 9 7 9 9 15 1 10 9 3 13 2
18 13 13 10 9 0 9 16 9 7 10 9 13 10 9 1 9 13 2
6 11 2 11 2 2 11
22 3 13 3 13 2 16 4 13 0 0 9 2 3 9 3 1 9 1 0 0 9 2
32 16 14 2 13 9 13 7 1 9 12 7 9 12 9 9 2 7 15 3 1 9 1 9 9 0 9 7 9 0 0 9 2
6 9 2 9 2 11 11
24 9 2 0 7 3 0 9 2 0 12 2 11 12 2 9 2 5 9 2 2 12 2 12 12
5 9 2 13 4 13
3 3 1 9
20 16 4 15 13 13 16 9 9 1 0 9 2 13 15 0 9 9 0 9 2
12 13 9 9 13 15 2 0 9 2 15 10 2
5 11 11 2 0 11
16 9 13 9 0 9 0 9 16 2 9 9 2 14 3 13 2
33 9 1 9 1 0 9 2 9 12 2 12 9 2 2 1 9 0 9 2 9 12 2 7 13 0 9 13 9 9 9 0 9 2
3 3 0 9
10 0 9 13 0 2 3 0 9 9 2
43 1 9 9 0 9 13 7 3 0 2 16 4 9 0 9 3 13 0 9 2 16 4 3 3 13 9 9 1 9 2 9 9 12 2 12 9 2 1 9 0 9 2 2
6 3 1 10 0 9 2
27 0 9 7 9 1 10 0 9 13 13 9 9 0 9 0 13 7 13 1 0 9 7 9 1 0 9 2
2 9 9
9 0 9 10 9 13 14 12 9 2
18 10 9 13 0 0 9 7 1 0 9 15 13 13 1 10 9 0 2
19 1 0 9 13 1 0 0 9 3 0 9 9 7 9 9 0 0 9 2
17 9 9 4 15 3 13 7 9 0 9 1 9 4 9 3 13 2
19 0 9 1 9 1 0 9 7 13 9 9 13 0 9 1 9 0 9 2
24 9 9 13 0 9 1 0 9 2 9 9 12 2 12 9 2 2 1 9 9 7 9 2 2
34 16 15 13 2 13 0 13 2 3 4 13 0 9 2 9 12 9 12 2 12 9 2 2 7 0 9 9 0 9 2 0 9 2 2
15 1 9 3 9 13 7 9 2 1 15 15 10 9 13 2
17 1 9 9 1 9 13 2 16 15 13 13 3 1 9 9 12 2
3 11 9 2
5 0 9 11 2 9
5 1 9 15 9 13
4 9 15 3 13
13 13 4 15 1 9 1 9 0 9 1 0 9 2
23 1 12 9 13 3 0 7 0 9 2 1 0 13 0 9 9 2 9 1 9 7 3 2
24 16 3 3 13 7 9 7 3 1 9 13 2 13 3 3 9 0 9 7 3 15 15 13 2
14 1 9 9 4 7 13 9 2 15 1 15 13 9 2
17 13 4 2 16 9 13 3 13 7 13 15 13 9 1 0 9 2
15 7 4 13 0 9 7 13 0 9 0 9 1 0 9 2
18 13 4 2 16 1 9 1 9 7 1 0 0 9 1 15 13 9 2
7 7 1 0 9 13 0 2
7 7 15 13 15 16 4 2
7 9 15 3 13 3 13 2
20 7 16 15 13 9 1 9 2 13 15 10 9 13 2 3 13 1 12 9 2
21 9 1 9 13 7 0 9 7 1 0 9 15 13 15 2 15 13 0 16 0 2
13 1 9 15 0 13 1 0 7 15 3 13 0 2
11 7 15 3 13 2 3 13 13 9 9 2
6 15 9 3 15 13 2
29 10 9 4 3 1 0 9 13 9 2 0 15 14 13 2 16 1 9 1 9 4 13 1 15 3 2 7 13 2
23 9 2 2 13 15 13 0 9 1 9 3 0 9 9 1 10 9 2 16 13 0 9 2
15 2 9 1 2 0 2 9 15 13 13 15 2 15 9 2
12 3 1 0 9 9 15 3 13 1 10 9 2
5 11 11 2 0 11
22 9 0 1 10 9 2 0 1 0 9 9 2 13 3 13 7 3 13 9 12 9 2
10 4 3 13 1 0 9 1 12 9 2
19 13 15 1 15 2 10 9 4 15 1 9 13 7 10 1 15 13 9 2
2 9 9
2 12 5
13 9 0 9 1 0 0 9 13 3 12 12 9 2
10 3 1 9 12 13 10 9 0 9 2
33 13 1 15 3 9 1 9 0 9 2 15 4 13 11 1 12 2 9 12 13 2 16 13 1 10 9 1 11 13 10 0 9 2
39 1 9 1 11 1 11 4 13 9 0 9 2 15 13 2 16 9 1 3 0 9 4 13 12 9 10 0 9 7 12 9 1 0 9 1 3 0 9 2
33 0 9 4 13 10 10 0 9 16 13 9 7 9 2 1 9 4 9 13 1 12 2 9 12 7 1 9 1 12 2 9 12 2
16 1 0 9 2 15 13 1 0 0 9 2 4 13 0 9 2
4 11 13 1 9
14 9 9 2 9 2 15 1 9 13 7 0 9 1 9
10 9 0 11 13 1 15 14 9 9 2
12 1 0 9 15 1 15 0 9 10 9 13 2
16 3 9 9 7 13 9 2 15 15 13 1 9 10 9 13 2
2 11 11
15 0 7 0 9 0 11 11 13 10 9 14 1 12 9 2
8 13 15 3 1 9 0 9 2
16 12 9 11 2 12 11 2 7 1 12 9 0 7 0 9 2
21 11 13 1 0 9 3 7 3 1 9 2 3 15 9 13 1 9 9 1 9 2
4 13 15 0 2
30 15 3 2 16 11 2 10 9 13 11 1 10 0 9 2 13 1 0 9 9 3 0 2 16 15 14 12 9 13 2
12 3 1 0 12 9 13 9 0 9 12 9 2
13 9 15 7 13 1 9 2 15 11 10 9 13 2
26 3 4 3 13 1 9 7 0 9 2 13 4 15 3 13 1 9 9 2 13 15 9 9 11 11 2
8 0 9 4 13 1 9 9 2
17 3 4 15 13 2 16 3 9 13 2 16 15 13 10 9 13 2
28 1 0 0 9 9 11 7 13 9 1 9 0 7 0 9 16 13 9 9 7 11 2 1 0 7 0 9 2
9 0 9 13 9 0 0 9 11 2
15 13 15 3 13 0 9 7 13 1 15 3 1 10 9 2
39 1 9 0 9 1 0 9 9 13 9 11 0 9 2 13 9 9 2 0 9 2 7 0 9 2 16 4 1 9 9 13 1 9 3 14 12 9 11 2
12 1 0 9 0 9 3 13 9 9 1 9 2
14 9 3 1 12 2 12 9 0 9 13 0 9 13 2
13 13 15 0 9 9 2 13 15 1 15 9 11 2
14 1 9 1 9 13 9 13 9 16 12 1 10 9 2
8 11 13 1 10 9 1 9 2
16 1 0 12 9 15 15 13 13 14 12 0 9 2 3 9 2
19 3 15 13 7 1 10 0 9 2 16 13 9 9 2 11 2 11 11 2
18 1 9 0 9 13 9 11 9 13 3 10 9 1 12 7 12 5 2
7 1 10 9 15 13 9 2
2 12 2
3 13 9 2
25 1 9 2 16 1 15 11 3 13 2 13 9 9 1 12 0 9 0 9 7 14 12 0 9 2
2 12 2
5 1 9 13 9 2
4 13 0 9 2
18 9 13 1 9 9 0 9 2 0 1 0 9 7 9 1 10 9 2
23 0 12 4 13 3 3 13 1 11 2 0 1 0 0 9 13 10 9 3 1 0 9 2
2 12 2
3 13 9 2
27 11 13 0 9 1 9 11 7 0 0 9 9 2 9 2 9 2 0 7 0 9 0 11 7 9 2 2
13 4 13 7 16 9 0 9 3 1 9 7 11 2
14 10 0 9 0 9 13 2 13 15 1 9 9 9 2
12 13 15 1 9 13 10 9 2 15 3 13 2
34 9 2 0 11 11 2 9 2 9 2 0 2 2 0 12 2 12 12 11 12 2 9 2 2 9 2 2 12 2 12 12 12 12 2
4 2 0 9 2
3 9 0 9
10 9 13 13 1 10 9 1 9 12 2
15 9 1 9 4 13 2 7 0 9 15 13 3 0 9 2
14 9 2 16 13 13 1 9 2 4 13 16 0 9 2
11 1 9 12 4 3 13 0 9 14 12 2
17 1 9 12 13 1 0 9 9 7 3 13 9 15 13 0 9 2
11 1 9 12 9 13 3 1 0 0 9 2
32 13 0 13 9 7 0 9 1 9 12 1 12 9 2 7 13 9 15 13 0 9 3 15 2 15 13 0 9 1 9 12 2
4 11 11 2 11
25 13 9 13 3 3 15 2 15 13 0 9 2 0 9 13 1 10 9 3 7 3 9 9 2 2
24 1 10 9 7 13 2 16 10 9 3 13 13 0 0 9 2 7 16 1 9 12 3 13 2
3 11 13 0
9 1 0 9 13 0 11 3 0 2
3 3 13 2
9 9 7 13 13 7 1 0 9 2
10 0 9 11 11 13 9 1 0 9 2
13 1 12 9 9 7 9 13 9 1 9 9 11 2
25 0 13 9 1 0 9 11 2 0 1 11 2 15 1 9 13 1 11 9 9 2 9 7 9 2
40 1 9 12 13 0 9 11 11 2 15 13 7 13 1 0 9 9 7 0 9 2 9 2 9 1 9 2 9 2 0 9 7 0 0 9 2 15 9 11 2
2 13 9
9 11 13 1 9 0 9 3 0 2
16 11 11 13 10 9 3 0 9 7 9 13 9 0 9 9 2
23 9 15 0 9 13 2 1 9 2 2 16 11 15 3 13 7 13 1 0 9 1 11 2
16 1 11 11 2 1 15 13 9 13 1 9 14 1 10 9 2
23 9 4 13 7 1 9 9 2 15 3 13 12 9 7 15 13 7 9 3 1 12 9 2
24 10 9 0 9 9 13 7 13 0 9 2 13 11 11 2 1 9 2 2 0 9 11 11 2
2 0 9
9 1 9 9 11 13 3 0 9 2
20 11 11 2 13 9 0 0 9 9 1 11 2 3 13 1 9 13 11 11 2
10 0 9 4 13 3 1 0 0 9 2
24 1 0 9 13 1 9 7 9 9 1 0 9 1 11 2 11 2 3 4 13 15 9 11 2
35 0 15 1 9 9 13 13 15 9 1 0 9 2 15 3 13 2 15 3 13 1 9 2 2 15 13 12 1 9 3 0 9 0 9 2
42 9 2 11 11 2 0 2 9 2 2 0 12 2 0 2 9 2 9 12 2 12 12 11 2 9 2 2 2 12 2 12 12 12 2 9 2 2 12 2 12 12 12
4 9 2 0 9
2 0 9
12 0 0 9 13 1 9 12 1 9 11 12 2
6 2 12 2 12 2 2
11 13 1 0 9 9 7 13 9 9 0 2
7 3 15 13 1 12 9 2
17 1 9 12 2 3 4 1 11 13 0 9 2 13 9 12 9 2
11 3 1 9 9 13 3 0 9 7 9 2
14 1 9 13 9 1 3 0 2 7 0 9 0 9 2
28 13 15 3 9 0 0 9 11 2 16 15 3 1 9 12 2 12 13 0 9 7 9 1 10 9 1 9 2
18 11 13 1 3 0 9 1 0 9 2 15 15 3 13 1 12 5 2
13 1 9 0 9 13 7 10 0 9 1 0 9 2
22 1 9 15 0 9 13 3 1 12 9 2 16 3 1 9 12 15 13 1 12 9 2
9 3 9 1 11 13 12 9 3 2
16 16 9 13 1 9 1 12 9 2 9 14 1 12 5 3 2
9 3 0 9 13 1 0 0 9 2
25 16 0 1 12 1 12 9 13 13 1 9 1 12 9 3 2 9 1 12 9 13 1 12 9 2
15 3 0 9 9 1 12 1 12 9 13 1 12 0 9 2
53 11 13 1 9 14 12 5 9 2 9 7 9 12 5 2 9 1 12 5 2 9 2 9 7 0 0 9 12 5 2 1 9 7 0 9 1 12 5 2 1 9 14 12 5 2 1 9 3 16 12 5 3 2
10 11 13 1 2 12 9 9 14 12 9
9 2 12 9 9 1 12 2 12 9
10 2 12 9 0 9 14 12 2 12 9
9 2 12 9 0 9 12 2 12 9
8 2 12 9 0 9 14 12 9
9 1 12 9 15 10 13 15 13 2
12 10 9 13 13 9 9 7 10 9 0 9 2
10 3 0 9 13 1 12 1 12 9 2
4 9 1 9 2
5 9 0 9 0 9
4 0 9 7 15
2 0 11
10 0 0 0 9 4 13 1 9 12 2
25 1 9 13 9 13 12 9 9 11 2 15 13 11 11 1 0 11 2 11 2 0 9 7 11 2
35 3 13 14 12 9 9 7 13 9 1 12 9 9 2 13 11 11 2 1 9 2 2 0 9 0 11 1 11 2 11 2 11 7 11 2
10 1 15 13 12 9 9 1 0 9 2
17 3 0 9 1 15 13 9 9 2 3 15 13 1 12 9 9 2
9 1 9 9 12 13 3 1 11 2
25 1 0 9 13 15 12 7 1 0 3 3 2 13 11 11 2 0 9 0 11 1 11 7 11 2
12 3 9 13 12 11 2 1 15 14 12 9 2
14 13 3 1 9 0 0 9 2 15 13 9 1 11 2
12 1 0 7 0 9 15 13 3 1 0 9 2
18 13 9 1 0 9 2 3 9 1 9 2 9 2 0 7 0 9 2
39 9 2 0 11 11 11 0 2 2 0 9 12 2 12 12 11 12 2 9 2 2 2 12 2 12 12 12 12 2 9 2 2 12 2 12 12 12 12 2
3 9 13 9
10 1 9 1 11 4 15 13 11 11 13
24 0 9 0 9 9 2 9 2 9 7 0 9 0 9 1 15 9 9 11 7 11 13 0 2
5 9 3 13 9 2
11 15 9 9 9 13 2 7 13 0 9 2
9 3 9 9 13 1 0 9 0 2
8 9 7 13 0 13 1 9 2
11 1 9 9 12 2 12 13 11 0 9 2
12 1 0 9 13 1 12 9 2 9 10 0 2
7 9 15 1 15 3 13 2
8 3 13 9 3 16 13 13 2
1 13
11 3 12 2 12 9 13 1 9 12 0 2
13 9 9 13 1 0 0 9 0 9 9 7 9 2
8 7 0 9 7 13 13 9 2
9 1 0 9 9 13 0 13 3 2
22 13 2 3 13 9 9 2 13 9 2 13 9 7 9 2 3 13 9 7 0 9 2
7 0 9 13 11 3 10 2
8 9 15 3 13 1 0 9 2
16 15 13 10 9 16 0 9 7 10 9 13 1 15 3 9 2
5 3 15 13 9 2
9 1 15 13 9 9 7 0 9 2
11 13 15 0 9 2 9 2 9 1 15 2
4 7 0 9 2
4 15 14 13 2
1 9
20 1 11 13 2 16 4 15 9 9 1 11 7 1 9 1 12 9 3 13 2
11 7 9 3 1 9 13 1 9 1 11 2
17 0 12 9 7 12 9 13 1 9 1 0 9 2 16 13 11 2
12 13 0 9 7 10 9 13 12 5 0 9 2
27 1 9 13 3 16 0 9 2 15 1 15 13 1 9 9 2 13 11 11 2 1 9 2 2 0 9 2
12 1 9 13 10 9 3 0 7 3 7 0 2
14 0 9 13 3 0 9 2 1 15 13 9 0 9 2
18 0 9 1 11 1 15 13 15 16 0 9 3 2 3 7 9 13 2
7 9 1 11 13 1 9 2
9 13 0 0 9 7 0 0 9 2
6 0 13 1 15 9 2
18 16 3 3 15 0 9 13 2 13 1 9 3 3 2 16 13 13 2
15 9 0 9 15 1 9 1 9 1 12 9 2 13 2 2
12 3 0 11 13 1 0 9 1 12 7 12 2
8 10 0 15 13 1 0 9 2
3 13 3 2
19 9 11 13 9 2 16 11 3 13 15 7 16 1 10 9 13 10 9 2
17 0 0 9 13 1 9 12 9 12 9 2 1 9 0 12 9 2
7 13 15 1 9 0 9 2
9 1 0 9 9 13 9 7 3 2
6 0 9 9 13 15 2
11 0 9 13 3 0 2 15 13 0 9 2
14 0 9 13 9 2 10 9 13 1 12 2 12 5 2
19 7 7 12 5 9 13 1 9 3 9 2 7 16 13 15 1 9 9 2
12 1 12 2 12 5 9 9 13 0 0 9 2
15 15 15 1 9 9 13 2 13 1 9 13 0 7 0 2
2 11 13
34 9 2 11 2 0 2 9 2 2 0 12 2 12 12 11 2 9 2 2 2 12 2 12 2 9 2 2 12 2 12 12 2 12 12
6 9 2 9 7 9 2
6 4 15 13 15 13 2
5 16 13 9 1 9
9 7 9 13 1 9 13 1 0 9
21 9 13 9 2 1 15 13 9 2 0 13 13 0 9 2 13 1 9 10 9 2
7 10 0 9 13 10 9 2
39 7 16 15 13 13 9 3 3 2 12 1 9 13 2 3 13 9 1 9 0 9 2 0 1 9 9 7 1 9 2 7 13 3 0 9 3 1 9 2
11 7 0 9 1 9 7 9 0 0 9 2
2 11 11
23 9 13 15 1 10 0 9 0 9 3 1 10 9 13 3 0 9 2 7 13 10 9 2
47 16 13 3 9 1 10 9 7 1 9 9 2 3 13 3 0 9 2 16 10 9 15 13 2 0 2 7 2 0 2 9 2 7 15 1 9 13 1 0 9 2 15 13 3 13 3 2
8 12 0 9 7 13 13 0 2
3 0 1 0
12 9 9 3 3 3 13 2 3 13 1 9 2
26 16 13 1 9 0 9 2 14 15 13 15 1 0 9 9 2 15 15 13 13 3 15 2 13 2 2
12 11 11 2 9 9 9 2 13 7 0 9 2
22 9 15 13 13 9 2 3 13 3 15 2 3 15 15 13 1 9 7 9 9 9 2
10 1 9 9 13 1 15 3 0 9 2
25 9 9 3 1 9 9 13 1 9 7 9 9 2 16 4 13 3 0 9 9 2 0 15 9 2
22 1 15 15 13 13 9 1 9 1 9 13 9 2 15 4 13 1 9 10 9 13 2
12 3 3 4 15 13 9 1 0 9 10 9 2
17 3 4 13 9 1 9 2 1 10 9 13 15 9 9 0 9 2
23 1 9 2 15 13 4 15 1 9 13 0 1 9 2 10 0 9 2 9 2 9 9 2
25 3 4 3 13 1 9 1 9 2 13 15 9 1 9 7 9 2 13 1 10 9 1 9 9 2
16 1 9 4 3 13 1 9 2 16 13 0 9 3 10 9 2
27 7 13 4 7 9 15 1 9 2 3 4 13 3 1 0 9 0 9 7 9 2 13 10 9 10 9 2
17 1 9 13 3 9 13 2 16 13 13 1 0 9 2 7 3 2
8 7 9 13 13 7 0 9 2
11 13 0 9 3 9 2 7 9 7 9 2
22 1 0 1 9 13 13 3 2 7 13 3 2 15 1 15 13 13 2 3 4 13 2
16 0 13 15 7 1 9 2 13 13 2 10 9 1 15 13 2
3 9 1 9
6 14 0 13 3 9 2
7 7 13 13 7 0 9 2
15 10 9 2 3 13 0 9 3 13 7 0 9 11 11 2
6 3 9 13 1 9 2
24 1 9 13 3 0 13 1 9 2 1 15 2 15 13 3 13 2 15 15 13 7 15 14 2
12 7 3 14 15 9 13 13 1 9 1 9 2
14 1 15 13 0 15 13 0 9 2 16 14 1 9 2
5 7 0 13 9 2
9 10 0 9 3 13 2 13 9 2
6 7 13 15 1 15 2
10 16 13 9 0 2 13 1 9 15 2
14 15 15 13 1 0 9 2 15 15 3 13 10 9 2
26 13 15 1 9 13 3 10 9 2 13 15 9 2 7 3 13 9 9 1 10 0 9 1 0 9 2
13 14 1 9 1 11 13 10 9 3 12 9 3 2
7 12 0 0 9 13 13 2
27 14 13 3 13 2 16 1 0 9 9 9 13 2 16 10 0 0 9 13 1 9 3 10 9 10 9 2
2 9 9
4 0 9 1 9
17 9 1 0 9 2 0 9 2 11 2 12 2 2 12 2 12 2
32 13 9 11 2 9 12 2 9 12 2 12 12 11 12 2 11 2 9 2 2 2 12 2 12 2 9 2 2 12 2 12 2
28 9 7 10 9 2 12 2 9 9 9 2 0 9 7 0 9 1 9 2 11 2 12 2 2 12 2 12 2
46 13 11 11 2 9 2 9 2 0 2 12 2 9 12 2 12 12 11 12 2 9 2 2 2 12 2 12 12 2 12 12 2 12 12 2 9 2 2 12 2 12 12 2 12 12 2
15 9 2 0 9 9 2 11 2 12 2 2 12 2 12 2
4 13 11 11 2
16 11 2 0 9 0 9 2 11 2 12 2 2 12 2 12 2
47 13 0 9 7 9 2 0 2 9 2 2 9 12 2 12 12 11 2 9 2 2 2 12 2 12 12 2 9 2 2 12 2 12 12 2 12 12 2 12 12 2 9 2 12 12 9 2
41 9 2 11 2 9 2 0 7 0 9 0 7 0 9 7 9 2 9 0 9 7 0 9 9 2 9 7 9 1 0 9 2 11 2 12 2 2 12 2 12 2
35 13 11 11 2 9 2 9 2 0 2 2 9 12 2 12 12 11 2 9 2 2 2 12 2 12 12 2 9 2 2 12 2 12 12 2
13 9 0 9 2 11 2 12 2 2 12 2 12 2
37 13 9 9 11 2 9 2 9 2 0 2 2 0 9 12 2 9 2 2 2 12 2 12 12 2 12 12 12 2 9 2 2 12 2 12 12 2
18 11 12 2 9 2 0 9 9 2 11 2 12 2 2 12 2 12 2
41 13 11 2 9 1 9 9 7 9 2 0 9 12 2 12 12 11 12 2 9 2 2 2 12 2 12 12 2 12 12 2 12 2 9 2 2 12 2 12 12 2
19 11 2 0 0 9 0 9 7 9 2 11 2 12 2 2 12 2 12 2
4 13 11 11 2
20 11 12 2 0 9 9 2 9 2 9 2 11 2 12 2 2 12 2 12 2
50 13 11 2 0 2 9 2 2 9 9 7 9 2 9 12 2 9 12 2 12 12 11 12 2 9 2 2 2 12 2 12 2 12 12 2 12 12 2 9 2 2 12 2 12 12 2 9 2 12 2
41 11 9 2 12 2 0 7 0 9 9 7 9 1 9 7 9 2 11 2 12 2 2 12 2 12 2 12 2 9 2 12 2 2 12 2 12 2 12 2 9 2
36 13 9 11 9 2 0 12 2 9 9 2 12 12 11 12 2 9 2 2 2 12 2 12 12 2 9 2 2 12 2 12 12 2 12 12 2
15 9 7 9 12 2 0 11 2 12 2 2 12 2 12 2
28 13 9 9 2 12 12 0 11 2 0 12 2 9 2 2 2 12 2 12 2 9 2 2 12 2 12 12 2
43 9 7 9 2 0 9 2 0 7 0 9 2 0 7 0 9 2 9 2 0 9 2 9 2 9 0 9 9 1 9 7 9 2 0 11 2 12 2 2 12 2 12 2
7 13 9 9 2 0 11 2
26 11 12 2 12 2 9 0 9 0 9 7 9 1 15 9 9 2 11 2 12 2 2 12 2 12 2
33 13 0 0 9 2 0 12 2 12 12 11 2 9 2 2 2 12 2 12 12 2 12 12 2 12 2 9 2 2 12 2 12 2
16 0 11 2 0 9 9 2 9 2 12 2 2 12 2 12 2
5 13 0 11 9 2
21 9 12 2 12 2 0 0 7 0 9 9 2 11 2 12 2 2 12 2 12 2
38 13 0 9 7 9 2 0 2 9 2 2 0 9 2 12 12 11 2 0 12 2 9 2 2 2 12 2 12 12 2 9 2 2 12 2 12 12 2
6 15 13 2 15 13 2
6 15 13 2 15 15 13
11 0 9 13 12 0 9 2 15 13 15 2
13 3 9 13 9 1 2 15 11 2 15 9 2 2
9 13 15 1 15 11 2 15 9 2
4 6 13 14 2
14 1 0 9 1 9 12 3 3 13 9 3 1 9 2
2 11 11
61 9 2 15 13 3 14 1 0 9 0 9 1 9 9 1 12 9 15 0 11 11 2 15 15 1 12 9 1 9 1 9 13 2 7 3 15 14 13 2 16 13 13 10 0 11 1 0 3 9 9 12 9 9 2 9 7 9 2 7 14 2
28 10 9 1 0 9 13 13 9 9 2 3 9 1 10 9 2 3 4 15 15 13 1 12 12 1 12 9 2
26 9 13 3 1 0 15 0 9 0 9 1 15 15 2 15 15 13 13 9 2 7 13 15 13 15 2
2 0 9
20 9 9 10 3 0 13 3 1 9 2 7 15 3 2 13 1 9 3 0 2
20 7 15 13 2 3 2 7 16 3 3 3 2 15 4 0 9 13 3 3 2
50 7 15 2 16 0 0 9 13 3 12 0 0 3 9 2 16 9 2 16 3 3 13 13 2 14 3 2 7 3 1 0 9 3 9 9 13 2 7 3 13 2 16 4 3 13 13 15 0 9 2
103 13 7 9 2 16 15 1 9 9 13 9 9 1 9 1 9 2 15 10 9 3 13 2 16 9 0 7 0 2 0 2 3 3 10 2 1 15 9 13 2 7 0 2 1 15 13 14 15 2 16 15 3 7 3 13 2 16 13 15 2 7 13 9 1 9 7 9 3 1 12 9 2 7 1 9 9 15 3 13 2 16 13 0 9 7 1 0 9 13 0 2 3 3 13 0 2 15 15 3 7 3 13 2
17 15 13 15 3 9 3 0 2 16 9 0 9 13 1 15 0 2
25 7 16 7 15 1 9 13 3 1 15 0 9 2 7 15 3 0 9 2 13 4 15 13 3 2
29 1 0 9 1 0 9 7 1 15 2 3 1 15 13 2 4 15 13 9 2 1 15 13 2 16 10 9 13 2
7 13 1 9 12 2 12 2
5 1 0 9 12 9
4 9 1 9 2
18 13 15 7 13 15 2 13 13 2 7 13 0 9 2 7 3 15 2
1 9
3 9 0 9
32 3 1 9 10 9 9 0 9 2 9 7 9 11 11 2 11 13 10 9 2 0 9 13 7 9 2 7 9 7 7 13 2
7 10 9 13 0 0 9 2
9 0 9 13 9 9 1 9 9 2
30 10 9 13 0 9 2 9 2 15 15 15 13 2 0 9 7 9 2 1 15 13 0 0 9 2 3 0 0 9 2
13 7 13 10 9 0 9 2 16 3 0 0 9 2
42 9 1 15 15 1 0 9 0 13 15 9 2 16 4 13 1 9 2 15 13 7 11 11 2 0 9 15 13 2 16 13 9 3 3 2 16 13 1 0 0 9 2
21 13 15 2 16 15 13 13 3 13 9 1 10 9 2 16 4 15 13 10 9 2
17 13 15 0 2 16 13 9 2 16 4 15 13 13 1 10 9 2
26 9 15 3 13 13 3 10 0 9 2 10 9 13 7 9 9 1 9 1 9 2 15 13 0 9 2
28 9 2 9 11 2 0 12 2 12 12 11 12 2 9 2 2 2 12 2 12 2 9 2 2 12 2 12 2
5 9 1 9 7 9
37 9 9 1 9 7 9 13 1 9 13 0 9 1 15 2 15 15 1 9 15 13 2 7 3 0 9 1 15 2 15 1 15 3 13 3 3 2
22 1 0 9 13 9 9 9 2 10 9 7 9 2 9 9 2 3 13 9 0 9 2
18 1 0 9 13 1 0 7 0 7 0 9 9 2 1 0 0 9 2
40 1 9 13 13 3 0 7 9 2 1 15 13 3 9 9 0 1 9 0 9 11 2 0 0 9 0 9 2 9 2 0 9 2 0 2 0 7 0 9 2
13 13 3 9 0 0 9 0 9 1 9 0 9 2
33 9 2 11 2 1 9 12 2 12 12 11 12 2 9 2 2 2 12 2 12 12 2 12 12 2 9 2 2 12 2 12 12 2
4 0 9 1 9
11 9 9 13 0 9 9 1 9 1 0 9
31 1 3 16 0 9 9 9 12 2 12 9 2 2 1 0 9 15 13 2 16 9 10 9 15 3 13 7 13 9 9 2
17 7 3 3 1 9 4 13 2 16 10 3 0 0 9 4 13 2
104 9 9 0 9 2 10 0 9 4 13 9 9 9 0 9 2 15 13 3 1 2 2 9 0 7 0 9 9 9 2 2 9 0 9 9 9 2 2 9 9 0 9 2 2 9 9 0 9 2 9 10 9 7 9 1 9 2 2 9 9 2 0 15 9 7 9 9 1 9 2 2 9 9 0 9 0 9 1 9 0 9 2 2 9 0 9 7 2 9 0 9 7 9 9 1 9 1 0 9 7 1 9 9 2
4 0 9 1 9
40 16 13 1 0 0 9 0 9 2 13 0 13 3 1 0 9 0 7 0 9 9 9 1 15 9 0 9 2 15 13 1 0 7 0 2 0 7 0 9 2
15 9 13 16 0 9 15 2 15 13 0 9 1 9 9 2
27 0 9 2 15 10 9 13 2 4 1 0 9 13 1 9 7 9 0 9 1 9 13 9 1 9 9 2
21 13 15 3 0 9 0 9 2 3 1 9 9 2 15 13 12 1 0 9 9 2
29 9 3 4 3 1 10 9 13 2 16 10 0 9 13 9 1 0 9 7 9 0 9 1 0 9 1 9 9 2
20 4 13 10 9 2 9 9 10 9 2 9 0 9 2 0 9 7 15 0 2
19 0 9 13 3 1 9 9 3 0 2 16 0 9 1 0 9 0 9 2
23 9 9 0 7 0 9 13 7 9 9 0 9 0 9 2 0 10 0 9 1 10 9 2
19 1 12 9 13 1 0 9 9 9 1 15 0 9 7 3 9 9 9 2
4 1 9 0 9
13 0 0 9 0 9 13 9 9 0 9 9 9 2
44 13 1 0 9 2 0 0 9 9 9 0 7 0 9 7 0 9 0 9 1 0 9 1 15 2 16 0 9 0 0 9 2 9 7 9 2 3 0 9 1 15 13 9 2
20 3 15 3 13 9 0 9 7 9 15 13 9 9 10 9 1 3 0 9 2
4 9 1 0 9
10 0 9 13 7 0 9 9 0 9 2
22 13 15 9 0 9 14 1 9 2 7 7 1 0 9 7 9 15 3 13 9 9 2
38 0 1 0 9 2 0 15 9 0 9 2 13 10 9 1 9 2 1 0 9 3 13 2 16 1 0 9 4 10 9 3 13 15 1 9 0 9 2
24 13 15 3 0 9 2 0 1 15 2 16 15 9 0 9 13 3 9 0 1 9 0 9 2
14 3 15 13 7 9 9 2 0 15 9 1 0 9 2
19 3 4 9 13 1 0 9 13 9 1 9 0 9 1 9 9 1 15 2
2 0 9
29 0 4 3 13 1 0 9 1 9 0 9 9 7 0 0 9 2 15 3 13 3 3 0 9 1 9 0 9 2
20 9 9 13 0 9 9 9 2 0 15 3 1 0 9 9 0 7 0 9 2
28 1 0 9 13 1 9 3 9 2 10 9 13 13 1 9 7 9 0 9 0 9 2 0 1 0 0 9 2
38 1 9 0 3 13 1 9 2 1 15 0 9 1 9 1 0 9 0 9 13 9 0 0 9 2 0 0 9 2 7 9 0 9 1 0 9 9 2
9 3 15 3 13 9 9 1 9 2
2 9 9
22 9 3 13 0 9 0 0 9 1 15 2 16 3 13 9 9 15 0 9 1 9 2
19 3 13 0 9 2 16 0 9 13 4 13 2 16 13 1 9 1 9 2
16 0 9 9 0 9 7 13 7 1 9 9 0 2 0 9 2
26 13 3 1 9 9 0 9 2 3 0 9 7 10 9 1 0 9 7 10 9 1 0 9 0 9 2
29 10 9 15 1 0 9 13 3 13 3 1 0 9 1 0 7 0 9 2 3 16 13 1 0 9 9 7 9 2
21 13 15 13 9 9 3 15 0 9 1 0 9 2 9 7 3 7 9 10 9 2
28 0 9 2 15 13 0 1 0 9 13 2 13 9 9 0 9 2 14 13 1 10 9 2 3 1 0 9 2
30 0 0 9 9 1 0 7 0 0 9 2 3 1 0 9 7 9 13 3 0 9 9 0 9 16 9 0 0 9 2
29 9 13 3 14 13 2 16 9 9 0 9 4 1 9 13 9 11 2 1 9 4 15 1 15 13 13 9 11 2
25 16 15 13 1 9 2 0 9 1 9 0 9 4 13 1 0 9 13 1 9 1 9 0 9 2
9 11 11 2 9 0 9 9 9 11
4 9 1 9 2
9 0 9 0 9 13 13 3 1 9
3 9 1 9
25 9 2 0 9 13 2 13 9 1 9 2 13 15 9 10 9 13 7 13 15 3 3 1 9 2
1 9
3 1 0 9
24 0 9 1 11 12 2 11 1 10 0 9 1 9 2 15 13 13 1 9 0 9 1 11 2
25 0 2 9 2 9 2 15 4 3 13 1 9 0 0 9 1 9 12 2 3 3 10 9 13 2
30 0 0 9 3 14 13 0 9 15 2 9 11 13 7 0 9 13 2 15 13 2 3 0 9 4 13 2 7 13 2
4 9 2 0 9
4 1 9 1 9
12 13 9 9 2 15 13 13 9 3 1 9 2
2 3 2
12 9 10 9 13 9 1 9 3 1 0 9 2
21 0 9 13 10 0 9 7 16 13 2 13 15 10 9 7 0 9 1 0 9 2
16 3 9 13 9 1 0 9 1 9 15 0 9 7 1 9 2
32 9 9 2 1 15 15 0 9 3 13 2 0 9 13 3 1 0 9 1 0 9 2 2 4 3 13 1 9 0 12 9 2
33 9 13 0 9 0 9 7 10 9 2 9 0 9 7 0 2 3 0 9 2 1 15 15 9 13 2 3 12 2 12 5 9 2
22 9 2 9 13 0 1 9 2 15 13 7 1 0 9 13 1 9 2 13 0 9 2
18 3 13 13 0 9 7 9 2 9 1 9 3 13 1 9 9 2 2
15 9 1 9 2 13 9 1 9 9 2 9 7 9 9 2
24 9 1 9 2 0 9 2 3 0 9 2 1 10 9 7 1 10 9 13 1 0 9 9 2
4 11 0 2 11
14 0 9 0 1 10 9 13 1 0 9 7 0 9 2
4 9 1 9 9
9 1 0 9 13 1 9 7 0 9
16 1 9 13 0 9 1 0 9 2 0 3 1 9 0 9 2
20 1 15 3 0 0 9 0 9 2 0 3 3 2 16 15 13 13 1 9 2
21 3 0 9 11 2 15 13 7 13 0 7 15 3 3 7 0 9 1 0 9 2
2 11 11
10 9 9 13 10 9 7 9 11 11 2
13 13 2 16 15 3 13 1 0 9 1 10 9 2
11 9 9 3 0 7 0 9 13 3 0 2
10 0 9 7 9 0 9 13 3 9 2
17 0 9 9 2 0 1 9 2 3 15 13 13 2 7 3 13 2
10 9 9 1 9 3 13 13 3 0 2
3 9 13 9
19 16 4 15 9 13 2 13 9 13 0 9 7 13 9 2 15 13 9 2
20 10 9 13 3 0 9 2 15 15 1 0 9 13 1 9 2 9 7 9 2
12 9 4 15 13 2 16 4 13 1 9 3 2
26 13 14 12 9 2 16 10 0 15 1 15 3 3 13 2 16 13 1 3 0 9 2 4 13 9 2
20 9 13 0 9 1 0 0 9 2 15 0 9 13 2 7 3 9 13 9 2
9 0 9 1 0 9 13 12 9 2
11 9 15 13 13 3 2 9 4 13 0 2
9 13 13 0 0 9 12 9 9 2
2 0 9
19 3 16 0 9 1 9 13 9 9 7 3 0 9 1 0 7 0 9 2
23 9 13 0 9 2 15 13 1 9 0 9 3 1 9 7 9 9 2 3 1 0 9 2
13 9 13 16 0 0 9 2 1 15 15 13 9 2
6 12 13 13 1 0 2
20 13 15 13 0 9 7 15 3 13 9 9 2 9 0 9 2 9 2 9 2
9 9 15 13 13 7 0 0 9 2
11 1 0 0 9 13 9 1 9 11 11 2
22 13 9 14 3 1 9 1 0 9 2 16 15 3 3 3 9 13 2 13 0 9 2
11 13 15 10 9 2 3 13 3 1 15 2
15 13 15 2 16 15 3 13 9 9 2 13 11 2 11 2
2 9 9
18 9 13 12 9 1 9 7 0 12 9 1 0 9 2 9 7 9 2
15 1 12 9 9 3 13 0 9 2 15 13 1 9 9 2
14 1 9 13 9 7 9 2 1 9 1 9 0 9 2
20 16 15 1 0 9 13 2 15 13 2 2 13 1 9 2 13 11 2 11 2
11 16 9 13 13 10 9 2 3 15 13 2
25 16 13 1 15 9 2 13 3 2 13 0 2 0 15 1 15 13 13 2 9 15 1 15 13 2
14 9 13 9 9 7 9 2 7 13 9 1 0 9 2
13 3 13 9 2 16 4 13 9 1 9 2 13 2
18 7 16 1 0 9 12 12 9 13 9 1 0 9 3 9 3 13 2
8 1 10 9 10 9 9 13 2
20 9 2 15 9 13 3 0 9 3 2 10 9 13 7 3 15 13 9 13 2
34 9 9 9 1 0 9 13 9 1 15 2 16 4 15 9 13 3 13 0 9 2 7 1 9 1 0 9 13 0 9 1 0 9 2
39 9 2 11 2 9 2 9 2 0 2 2 0 12 2 12 2 12 12 11 12 2 9 2 2 2 12 2 12 12 12 2 9 2 2 12 2 12 12 12
1 9
15 0 9 9 15 1 9 11 13 12 9 2 9 1 9 2
13 13 13 9 2 0 9 1 9 7 0 1 9 2
3 9 2 9
11 0 0 9 13 9 1 0 9 0 9 2
20 1 9 0 9 1 15 13 1 10 9 13 0 9 0 9 7 9 0 9 2
26 13 9 13 1 0 9 2 15 13 3 3 13 9 7 9 0 9 2 3 13 9 0 9 1 9 2
27 3 1 9 9 0 11 15 13 1 9 9 13 14 12 7 0 9 9 16 13 15 1 9 1 0 9 2
6 11 11 2 0 0 9
2 13 13
14 9 1 0 9 2 0 9 2 13 0 9 0 9 2
21 13 0 15 2 16 15 9 13 0 0 9 7 15 13 12 0 9 1 12 9 2
17 13 15 2 16 1 0 9 13 0 13 1 9 9 3 12 9 2
22 3 1 15 15 4 1 9 9 13 0 9 1 10 0 7 9 3 13 9 0 9 2
29 1 0 9 13 2 16 9 9 2 15 13 12 2 9 2 13 12 2 9 7 9 0 9 13 0 12 2 9 2
20 3 15 0 9 13 12 9 2 1 0 9 15 13 12 2 3 0 13 12 2
20 1 0 9 15 13 3 1 9 1 9 12 9 2 9 7 9 13 12 9 2
3 2 13 2
27 1 9 12 2 9 15 13 0 9 2 9 9 1 0 9 9 1 0 9 7 9 1 0 9 1 9 2
67 1 9 12 2 9 13 9 1 9 9 7 9 0 9 2 9 2 9 1 9 9 2 10 0 0 9 13 9 12 9 2 9 2 9 0 9 1 9 9 2 10 0 0 9 13 9 12 9 7 13 9 12 9 2 9 2 9 0 9 1 9 1 9 0 0 9 2
35 3 15 13 9 7 13 9 1 0 9 2 7 2 9 1 12 2 9 9 1 0 0 9 2 9 2 9 1 9 9 1 0 0 9 2
5 2 9 7 9 2
29 2 1 0 9 15 13 9 1 9 12 0 2 2 9 2 15 13 13 9 0 0 2 2 9 7 0 0 9 2
16 9 10 9 1 9 0 9 9 13 1 2 0 9 2 9 2
30 15 13 1 9 3 2 2 9 1 9 2 7 13 15 3 13 1 9 2 2 9 2 0 1 0 9 0 11 11 2
43 16 9 3 1 12 9 13 2 9 14 13 2 2 0 9 2 1 9 9 13 10 0 9 2 2 16 9 0 9 9 14 13 3 0 2 2 2 16 3 0 0 9 2
2 9 2
23 3 3 13 9 7 9 9 1 15 2 3 1 0 9 13 2 16 4 15 13 0 9 2
21 16 7 9 1 9 13 15 2 3 15 13 15 1 0 9 13 3 15 1 15 2
1 11
3 1 0 9
14 9 11 1 9 3 0 9 11 7 10 9 9 11 2
14 9 13 1 0 9 7 9 0 0 9 1 0 9 2
15 9 9 1 9 9 7 9 9 13 0 9 9 1 9 2
38 9 2 11 2 9 2 9 2 0 2 2 12 12 11 9 2 12 2 9 2 2 2 12 2 12 12 12 2 9 2 9 2 2 12 2 12 12 12
1 11
24 9 11 11 1 0 9 9 1 9 0 9 2 1 15 13 0 9 0 9 2 9 7 9 2
16 9 13 0 9 3 1 9 1 0 9 7 0 9 1 9 2
7 9 15 13 7 9 9 2
39 9 2 11 11 2 9 2 9 2 0 2 2 0 12 2 12 12 11 12 2 9 2 2 2 12 2 12 12 12 2 9 2 2 12 2 12 12 12 2
3 9 0 9
25 3 15 15 7 15 1 9 2 0 9 7 9 13 2 16 13 1 9 7 9 0 9 0 9 2
35 3 15 15 13 13 2 16 14 3 2 1 0 9 2 13 1 10 9 9 9 0 10 0 9 1 0 9 7 1 9 7 9 10 9 2
5 3 13 15 0 2
9 3 15 10 9 13 7 13 9 2
19 10 9 13 13 0 2 7 14 3 13 3 1 10 0 9 13 0 9 2
20 15 3 13 2 16 15 15 13 9 7 0 9 13 1 0 9 2 0 9 2
17 0 7 13 9 2 3 9 13 7 13 7 9 0 1 0 9 2
14 1 10 9 13 1 9 9 1 15 2 3 9 13 2
30 1 9 4 13 13 1 9 0 1 9 0 9 2 3 3 9 0 15 1 9 2 9 2 9 2 0 9 2 9 2
14 3 15 13 2 16 9 0 9 15 13 13 1 9 2
16 1 10 9 7 13 1 0 9 2 1 15 13 12 0 9 2
27 1 10 9 13 3 2 16 15 13 3 3 2 16 1 9 9 9 13 9 2 15 4 13 1 0 9 2
56 15 4 13 2 9 2 10 9 13 2 14 15 15 3 3 13 2 9 13 3 2 0 2 7 2 0 13 9 1 9 1 0 9 2 9 7 0 9 9 1 10 9 2 2 15 9 12 9 2 12 9 0 9 7 9 2
12 13 15 2 1 9 2 3 1 12 0 9 2
5 13 1 15 13 2
33 12 2 15 3 13 7 13 9 1 0 0 1 9 1 9 0 9 2 4 13 9 9 14 1 12 9 7 9 9 7 0 9 2
35 12 2 3 4 13 2 15 9 1 0 2 0 1 9 1 9 10 9 2 9 7 9 13 7 13 2 7 15 13 0 9 0 9 9 2
19 3 13 13 2 0 9 4 13 13 1 10 9 9 0 7 2 0 2 2
2 11 11
4 1 9 1 9
8 15 13 9 7 9 9 7 9
9 1 0 9 9 2 9 13 9 2
9 1 9 7 13 0 13 7 9 2
22 0 7 0 15 1 9 13 15 2 7 14 3 13 10 9 1 9 1 0 0 9 2
8 3 7 1 15 13 0 9 2
19 0 9 13 1 0 9 9 1 9 3 9 0 2 0 9 9 1 9 2
36 1 15 13 2 2 9 9 1 9 0 9 2 2 9 9 1 9 9 1 9 9 2 2 9 9 1 9 1 0 9 2 15 13 0 13 2
49 0 0 9 0 1 0 9 2 0 9 9 1 9 2 3 10 9 1 9 1 0 9 2 15 13 0 13 2 13 1 9 12 7 12 9 9 2 12 2 12 9 2 2 9 9 1 9 9 2
44 3 13 13 2 16 9 2 15 1 9 9 1 0 9 13 10 9 1 0 9 2 1 9 2 16 1 9 2 15 13 9 0 13 2 13 9 2 13 1 3 0 9 9 2
4 9 1 0 9
15 9 10 9 9 9 13 9 1 0 9 1 9 7 9 2
42 15 15 13 3 1 10 9 2 15 13 9 9 7 9 2 13 3 1 9 1 9 7 0 9 7 3 3 1 9 2 3 2 10 9 2 2 15 4 9 9 13 2
12 10 9 13 4 13 3 3 2 3 13 0 2
16 3 10 9 13 4 13 14 1 9 2 15 13 12 9 9 2
2 9 9
56 1 12 9 9 13 9 1 10 9 13 1 9 2 16 4 13 1 0 9 2 13 1 0 9 2 13 2 7 1 9 2 16 9 1 9 1 12 9 1 9 0 9 13 9 1 0 9 2 15 13 0 9 1 0 9 2
42 1 9 2 3 15 13 9 1 0 0 9 1 9 1 3 9 3 2 13 9 1 10 0 9 13 2 16 4 1 9 13 0 9 7 4 13 0 9 7 10 9 2
8 10 9 13 9 13 9 3 2
14 7 3 2 9 1 0 9 13 3 9 9 0 9 2
1 9
28 13 13 2 16 1 9 2 9 12 2 12 2 13 3 2 16 4 10 9 4 3 13 3 9 2 3 9 2
32 1 9 9 13 0 0 9 1 0 9 1 9 2 16 1 0 9 9 0 13 1 9 2 13 13 3 9 2 9 2 9 2
23 10 9 1 0 9 13 12 1 9 9 9 1 9 1 0 9 2 15 13 9 0 13 2
42 1 9 2 16 4 13 9 7 13 0 7 1 9 13 9 2 13 9 15 0 2 16 13 1 9 1 12 9 9 7 13 1 9 0 9 1 0 9 9 1 9 2
32 1 10 9 13 13 1 9 0 0 9 9 1 9 0 9 2 7 1 0 9 1 15 2 7 9 13 3 0 13 0 9 2
2 11 11
28 13 0 9 11 2 0 2 0 12 9 2 12 12 11 12 2 11 2 9 2 2 2 12 2 12 12 12 2
4 9 1 9 2
18 9 13 9 2 1 9 9 7 13 3 13 1 9 2 7 7 9 2
1 9
4 13 15 9 9
9 10 9 15 13 1 0 0 9 2
10 13 4 1 15 0 9 2 13 9 2
15 13 0 9 2 0 9 2 9 9 7 9 13 3 0 2
5 13 4 1 15 2
4 11 11 2 11
27 14 13 0 9 2 13 15 3 0 9 7 16 0 3 13 9 10 9 2 9 1 9 0 9 7 9 2
12 13 15 7 1 9 10 9 2 9 2 9 2
14 3 3 13 10 9 2 3 15 4 3 13 1 9 2
7 7 15 13 7 0 9 2
13 9 0 15 0 9 4 13 13 0 7 0 9 2
3 13 0 2
5 16 14 2 3 2
8 7 13 3 3 0 2 0 2
6 13 7 13 0 9 2
15 13 15 9 1 9 3 2 3 7 13 3 3 3 0 2
18 1 9 13 9 2 7 13 3 9 11 1 0 9 14 13 10 0 2
10 13 1 9 2 9 7 9 0 9 2
25 9 15 3 1 15 3 3 13 13 3 7 3 2 7 3 15 4 13 3 13 0 9 1 9 2
8 13 4 7 3 13 10 9 2
8 3 4 13 1 15 13 9 2
19 15 13 14 10 9 2 15 15 13 0 9 13 3 1 0 9 7 9 2
11 3 13 0 13 10 9 13 9 7 9 2
14 3 0 9 15 13 15 13 1 0 9 2 15 13 2
16 1 3 0 9 4 13 9 2 16 4 13 3 10 0 9 2
9 13 15 1 10 9 13 9 9 2
19 1 9 7 9 0 0 9 13 3 3 7 1 3 9 13 0 0 9 2
14 0 9 7 0 0 9 13 0 9 3 0 9 9 2
3 11 11 2
3 9 11 12
35 9 2 11 12 2 0 15 2 12 2 12 12 11 12 2 9 2 2 2 12 2 12 12 2 9 2 5 9 2 2 12 2 12 12 2
3 1 0 9
12 13 13 1 15 7 14 7 14 15 15 13 2
2 15 2
2 9 2
25 13 14 15 0 2 7 3 7 9 2 15 13 3 0 7 13 1 9 9 3 3 16 15 9 2
9 3 13 15 3 1 9 1 15 2
20 13 15 15 1 0 9 7 3 9 12 7 12 0 2 3 0 2 9 9 2
4 13 7 13 2
7 3 13 13 2 3 3 2
8 7 3 15 3 15 13 13 2
24 7 3 1 15 0 9 1 9 2 15 13 13 2 16 0 1 0 9 2 0 9 0 9 2
4 13 0 9 2
7 0 9 1 9 12 9 2
17 15 13 9 1 15 2 15 15 9 1 0 9 13 1 0 9 2
8 1 0 9 1 9 0 9 2
6 3 13 9 1 9 2
13 1 15 9 13 1 0 9 1 0 9 10 9 2
7 9 9 1 11 3 13 2
9 13 15 2 15 13 3 3 13 2
7 7 1 0 9 13 9 2
27 1 15 15 13 7 3 13 10 2 9 2 9 2 1 15 15 13 1 0 7 0 9 0 9 10 9 2
2 9 9
5 13 15 3 13 2
7 3 15 13 13 9 10 9
2 12 2
17 13 3 1 12 2 9 7 1 9 2 16 15 13 1 9 9 2
2 12 2
20 9 0 9 1 0 9 3 3 13 9 9 9 2 7 3 9 0 9 9 2
2 12 2
12 13 1 0 9 13 3 9 1 9 0 9 2
2 12 2
22 13 1 0 9 13 3 9 1 0 9 7 10 9 15 13 3 13 16 9 9 0 2
2 12 2
28 13 2 14 0 9 1 9 2 15 10 9 3 13 2 13 1 15 2 7 15 3 2 13 15 15 1 15 2
2 12 2
13 1 9 1 9 7 10 9 13 2 0 9 2 2
12 15 13 7 1 9 1 9 2 13 3 13 2
2 12 2
21 16 3 13 13 1 0 9 2 13 1 9 2 15 13 3 2 9 3 15 13 2
11 7 13 2 16 16 0 9 15 15 13 2
2 12 2
12 16 13 1 9 14 12 9 2 3 9 13 2
11 13 1 12 9 1 12 9 13 0 9 2
2 12 2
10 13 15 1 9 9 9 1 0 9 2
20 7 3 15 13 3 0 9 1 0 9 2 16 10 0 9 3 13 9 0 2
2 12 2
26 13 9 1 9 2 15 13 1 9 2 13 13 3 0 2 1 9 0 9 3 1 9 3 15 13 2
5 9 2 9 7 15
3 9 1 9
12 13 0 9 2 15 1 9 12 9 13 9 2
37 16 4 13 1 0 9 2 16 13 1 9 13 0 9 2 9 2 9 2 9 2 13 9 2 16 1 9 1 12 9 13 12 9 9 9 11 2
17 9 9 15 3 13 13 1 10 0 9 2 15 1 9 13 9 2
13 13 10 9 0 7 1 10 9 15 0 9 13 2
7 11 2 11 2 2 0 11
23 1 9 1 9 9 15 13 2 16 4 15 13 1 0 9 2 15 13 0 9 0 9 2
75 16 13 1 0 9 1 9 0 7 0 9 2 3 0 9 1 0 9 2 4 13 9 9 12 2 12 9 2 2 1 9 2 0 9 2 7 9 11 9 2 12 2 12 9 2 2 1 0 9 1 0 9 2 15 7 4 13 9 9 2 12 2 12 9 2 2 7 9 9 2 12 2 12 9 2
3 9 7 9
16 1 9 1 9 15 2 12 9 2 4 13 9 1 9 9 2
19 12 1 15 13 14 1 12 9 1 9 0 0 9 16 0 9 7 9 2
32 1 9 9 4 15 3 13 2 16 9 13 9 1 0 9 1 15 2 16 15 4 13 1 9 9 9 10 9 16 0 9 2
8 13 15 0 13 1 0 9 2
6 11 2 11 2 2 11
17 16 4 1 9 9 13 9 2 13 3 10 9 13 3 0 9 2
10 1 15 13 13 2 16 9 13 0 2
20 7 13 3 15 13 9 2 16 1 10 9 13 0 13 9 9 1 0 9 2
11 9 13 3 13 3 1 0 9 1 9 2
4 9 1 0 9
7 1 9 15 4 13 9 2
16 13 7 1 3 0 9 2 16 1 9 2 3 15 4 13 2
10 13 0 13 3 10 9 1 0 9 2
6 11 2 11 2 2 11
50 1 10 9 15 13 1 9 3 3 2 7 0 9 13 13 2 3 13 13 2 16 4 13 0 9 0 1 9 9 2 12 2 12 9 2 2 1 9 9 9 2 12 2 12 9 2 7 0 9 2
21 1 10 9 13 9 9 0 9 9 2 9 1 9 9 0 1 9 2 2 2 2
12 1 15 4 9 9 1 9 0 9 13 3 2
37 2 9 15 13 3 1 9 2 3 10 0 9 1 9 4 1 9 9 11 13 1 12 2 9 12 2 3 1 15 3 3 4 13 7 1 9 2
14 2 9 13 13 0 9 9 9 9 1 9 0 9 2
15 10 9 13 13 9 2 15 4 13 9 9 1 0 9 2
5 13 1 10 9 2
21 2 9 0 9 2 16 0 9 13 1 9 9 3 9 2 1 15 4 13 9 2
14 2 9 2 15 13 2 16 4 9 13 1 0 9 2
31 0 9 9 9 1 9 9 2 3 0 9 2 13 0 9 2 0 9 2 2 2 2 7 15 13 7 1 9 9 9 2
10 15 3 13 9 9 1 0 9 9 2
3 9 0 9
19 13 3 9 2 7 1 1 9 13 3 0 9 2 16 13 9 10 9 2
10 13 7 9 13 16 9 1 9 9 2
20 10 9 4 13 1 10 9 9 0 1 9 9 9 2 3 0 7 0 9 2
6 11 2 11 2 2 11
63 0 0 9 13 9 0 9 1 10 9 2 2 1 9 0 9 2 2 1 9 0 9 7 9 1 0 9 2 2 1 9 0 9 2 3 9 2 9 2 0 9 2 9 3 2 2 2 2 16 0 9 1 9 0 9 1 9 1 9 3 0 9 2
22 3 3 13 2 16 0 9 13 13 1 0 7 15 0 9 7 10 9 4 13 9 2
17 13 0 7 3 7 0 2 16 13 3 13 2 10 9 13 0 2
21 1 15 4 13 3 2 13 2 0 9 1 9 9 9 2 3 0 7 0 9 2
20 3 13 2 16 1 9 9 0 9 13 1 0 0 9 9 9 7 9 9 2
31 3 4 9 13 9 2 3 9 7 9 2 1 9 1 9 2 9 13 2 7 3 0 0 9 13 3 9 9 1 9 2
10 1 9 0 9 13 0 13 0 9 2
30 9 13 0 9 11 2 11 2 9 2 0 9 12 2 12 12 11 12 2 9 2 5 9 2 2 12 2 12 12 2
5 13 9 9 2 12
13 11 2 0 0 9 9 2 15 13 1 10 9 2
25 13 4 0 0 9 7 1 9 4 13 14 9 0 2 0 2 13 15 1 0 9 9 11 11 2
13 0 0 9 13 0 9 0 9 7 3 7 9 2
15 13 15 2 16 1 0 15 0 9 13 7 9 1 9 2
14 9 1 11 15 13 0 9 2 1 15 9 15 13 2
11 1 9 9 11 13 7 0 9 1 11 2
7 9 11 2 11 2 11 2
4 9 1 0 9
6 9 13 9 1 0 9
22 13 9 1 15 2 16 9 10 9 13 9 1 15 3 0 9 2 13 3 0 9 2
27 16 4 15 10 9 13 11 11 13 2 13 13 1 0 9 2 3 15 10 7 0 9 1 0 9 13 2
23 1 0 9 15 3 15 13 2 16 4 1 10 0 9 11 13 9 9 0 9 0 9 2
24 2 2 2 2 2 2 2 2 2 2 2 2 2 2 2 2 2 2 2 2 2 2 2 2
2 11 11
23 2 2 2 2 2 2 2 2 2 2 2 2 2 2 2 2 2 2 2 2 2 2 2
20 1 9 15 13 14 9 9 2 11 15 13 7 1 0 9 1 9 11 11 2
2 0 9
57 10 0 0 9 2 0 1 9 9 2 7 0 1 0 9 9 2 0 1 9 2 0 1 9 7 0 1 10 0 9 2 15 1 9 1 0 9 9 0 9 13 9 9 7 13 1 9 9 9 2 15 13 1 0 9 0 2
18 1 15 15 3 3 13 2 1 10 9 2 10 9 7 10 9 13 2
24 7 16 1 0 9 15 13 9 13 1 9 2 13 15 3 9 9 2 3 1 15 3 13 2
20 0 9 2 15 11 13 1 9 2 15 13 9 0 9 1 9 1 0 9 2
36 16 1 0 0 9 13 13 0 9 2 0 9 4 3 3 13 7 9 15 3 13 0 9 9 2 7 15 1 9 1 10 9 7 0 9 2
28 13 15 2 16 15 2 7 3 0 9 0 9 1 0 9 2 4 15 13 13 9 1 9 7 0 9 9 2
6 0 9 13 9 9 2
2 9 13
49 4 2 14 13 2 16 1 0 9 3 15 11 11 13 1 9 0 9 2 13 3 13 10 9 15 2 16 3 15 3 15 13 1 15 2 16 4 13 1 9 9 9 2 15 1 10 9 13 2
22 0 9 9 1 9 13 11 11 2 9 9 0 11 2 15 13 1 10 9 0 9 2
20 1 0 9 15 1 15 11 11 13 2 16 0 1 15 4 13 16 0 9 2
17 0 11 15 13 9 7 9 9 2 11 9 0 9 7 0 9 2
15 1 15 2 16 1 9 7 0 9 15 4 13 1 9 2
13 7 9 13 2 16 13 0 13 0 9 0 9 2
12 7 15 3 13 13 2 16 15 10 9 13 2
11 3 4 15 13 13 7 10 9 1 9 2
2 13 9
8 0 9 9 13 3 9 9 2
23 13 15 0 2 16 13 1 3 0 9 2 3 13 0 0 9 13 1 10 9 7 9 2
12 1 9 9 1 9 13 9 3 1 0 9 2
25 1 0 9 2 15 13 13 9 9 3 14 9 1 9 0 0 9 2 13 11 11 1 9 9 2
7 0 13 9 1 0 9 2
21 3 1 9 1 0 11 15 11 13 13 9 1 0 9 7 0 9 9 1 9 2
10 1 10 0 9 13 9 1 9 9 2
25 1 1 15 2 16 1 9 13 1 9 2 15 13 1 9 7 1 0 9 2 13 15 9 9 2
20 7 13 2 16 15 4 13 9 1 9 0 9 9 7 16 13 7 9 9 2
2 11 11
30 9 2 11 2 0 12 2 12 12 11 2 9 2 2 2 12 2 12 2 9 2 2 9 2 2 12 2 12 12 2
11 9 1 9 2 9 13 13 1 9 9 2
3 9 1 9
11 9 1 9 2 9 2 9 7 0 9 9
14 13 1 10 9 9 2 15 10 9 13 13 0 9 2
21 3 13 0 13 15 1 0 9 9 1 9 0 9 2 1 15 15 13 7 9 2
2 11 11
28 1 9 0 0 0 9 11 13 13 9 2 15 13 1 0 9 0 9 2 16 9 2 9 7 0 9 9 2
25 13 7 2 16 1 9 9 13 2 16 9 4 13 13 3 0 9 7 3 15 13 3 12 9 2
41 16 9 9 4 1 0 9 2 15 13 1 9 1 11 11 2 9 0 9 2 0 9 7 1 15 0 9 1 9 2 13 9 2 9 7 9 2 9 7 9 2
47 1 0 9 9 9 13 2 2 0 9 1 9 9 7 9 9 2 2 9 3 13 2 2 9 1 9 9 2 9 2 9 7 9 2 2 9 9 2 2 0 0 9 9 9 1 9 2
20 9 9 1 9 13 1 9 2 7 9 13 0 13 14 1 12 2 9 12 2
41 9 2 11 2 0 9 2 15 2 12 2 9 12 2 12 12 11 2 9 2 2 2 12 2 12 12 2 12 12 2 9 2 2 12 2 12 12 2 12 12 2
8 0 9 0 9 1 12 2 9
8 2 9 1 12 2 9 12 2
3 2 9 2
8 9 2 9 11 7 9 11 9
51 0 9 9 13 0 9 1 9 9 9 1 0 9 0 9 2 9 3 1 0 12 9 13 12 9 0 0 9 10 9 1 0 0 9 12 12 9 1 12 0 9 2 7 10 0 9 13 1 0 9 2
16 15 13 3 2 13 3 10 9 13 1 9 1 12 12 9 2
19 14 14 12 9 9 13 1 15 9 0 9 1 3 2 16 9 12 9 2
3 9 0 9
4 2 9 12 2
3 11 11 11
4 9 2 9 11
4 0 9 1 9
8 9 13 13 2 14 2 0 2
5 3 10 9 13 2
4 0 9 13 2
8 9 9 1 9 15 3 13 2
4 9 13 9 2
9 9 15 1 0 9 13 0 9 2
7 1 10 0 15 13 9 2
10 9 15 13 9 2 15 13 13 9 2
13 9 7 13 13 2 13 15 2 16 9 13 3 2
2 11 11
13 0 9 2 0 1 9 0 9 2 13 0 9 2
10 1 9 9 13 3 2 13 15 9 2
11 9 13 3 1 9 2 7 9 7 13 2
13 9 2 0 1 0 9 0 9 2 13 13 9 2
8 9 9 1 9 9 13 9 2
1 13
11 1 9 12 13 9 1 9 1 12 9 2
9 1 9 15 13 12 2 12 9 2
12 9 13 12 9 7 10 9 12 9 1 9 2
16 13 13 2 0 2 9 2 13 12 2 12 9 1 9 2 2
16 0 0 9 13 10 9 9 1 9 7 9 9 1 12 9 2
13 13 15 3 7 1 9 1 9 13 0 1 9 2
20 13 1 15 9 9 2 9 1 12 9 2 7 9 2 9 1 12 9 2 2
5 9 13 3 0 2
20 3 13 11 11 2 9 0 9 1 11 2 13 15 15 12 2 12 5 0 2
3 15 13 2
14 3 3 15 13 7 9 9 1 9 12 2 12 9 2
9 9 9 1 9 9 15 3 13 2
18 16 9 3 13 12 0 9 2 16 9 9 13 0 9 2 13 9 2
9 9 2 9 2 9 7 3 9 2
5 13 9 7 9 2
12 1 9 15 3 13 9 2 15 13 9 0 2
2 3 13
13 9 7 9 13 3 13 2 16 9 13 10 9 2
10 1 9 15 9 2 9 7 9 13 2
10 1 0 9 15 15 13 9 9 3 2
24 9 3 13 10 9 1 9 9 2 15 1 0 9 2 13 2 0 9 0 2 3 0 9 2
6 1 9 13 13 9 2
10 7 15 15 2 9 2 3 3 13 2
13 9 15 13 1 9 1 0 9 7 9 0 9 2
12 3 16 4 15 10 9 3 13 2 13 15 2
4 0 13 9 2
12 1 9 13 15 3 0 2 7 7 3 0 2
14 0 9 13 1 9 13 1 9 9 2 9 15 13 2
13 9 1 10 9 13 0 2 13 15 1 15 3 2
23 9 13 9 7 9 10 0 9 13 0 16 9 7 9 2 13 0 9 2 13 0 9 2
7 9 15 1 15 3 13 2
19 9 15 13 1 9 2 13 15 9 2 0 9 0 9 9 1 9 9 2
28 1 10 9 15 3 3 13 2 16 15 3 13 13 2 16 9 4 13 9 0 7 0 2 7 16 15 13 2
12 9 3 15 13 2 7 15 15 15 13 13 2
14 9 2 9 2 9 2 9 2 9 2 9 2 2 2
3 1 9 9
18 9 1 9 13 3 9 1 9 1 9 0 9 2 15 1 9 13 2
14 1 9 15 1 0 9 10 9 3 13 1 15 0 2
9 10 9 2 10 9 2 10 9 2
9 9 9 1 9 10 9 3 13 2
20 9 2 0 9 7 9 2 15 3 13 1 10 0 9 7 13 1 9 3 2
7 10 9 13 13 1 9 2
7 9 13 1 9 0 9 2
6 9 9 1 9 13 2
5 13 10 0 9 2
7 7 3 13 15 1 0 2
17 9 4 13 13 2 16 4 13 9 2 1 15 13 3 1 9 2
9 7 15 0 9 13 3 1 15 2
10 15 13 13 2 16 4 1 9 13 2
11 13 1 0 9 9 7 15 13 13 15 2
8 9 15 13 2 7 16 3 2
12 3 4 13 15 1 15 7 13 15 0 9 2
3 13 13 2
6 1 9 13 15 0 2
13 3 2 13 4 13 9 2 15 13 3 10 9 2
13 9 13 2 9 2 7 15 1 15 3 15 13 2
8 1 0 9 13 9 3 3 2
11 9 1 15 13 13 3 1 9 1 9 2
7 10 9 13 7 2 2 2
11 0 9 7 0 9 9 15 13 1 9 2
15 3 4 0 9 13 0 9 1 9 9 14 1 9 9 2
11 10 9 15 3 4 13 13 7 15 3 2
8 16 9 4 13 0 9 3 2
8 16 13 3 0 9 7 13 2
6 13 2 13 3 9 2
8 7 1 9 13 3 13 9 2
9 9 7 9 9 1 15 3 13 2
1 9
5 9 9 15 13 2
6 13 13 7 1 9 2
14 0 9 13 3 3 0 2 7 13 10 2 9 2 2
6 7 13 13 0 9 2
7 3 2 9 13 1 9 2
13 13 0 15 13 2 16 9 13 10 9 1 9 2
12 13 4 15 1 15 2 7 13 3 1 9 2
5 7 9 13 0 2
14 9 2 16 9 13 9 14 3 1 9 2 13 0 2
3 9 1 9
1 9
2 9 12
5 12 5 0 9 12
6 12 5 9 1 9 12
4 12 5 9 12
7 12 5 9 1 12 9 12
4 12 5 9 12
2 9 12
4 9 1 9 12
7 9 1 9 1 12 9 12
2 9 12
5 0 9 7 9 12
4 12 5 9 12
4 12 5 9 12
2 3 12
3 9 1 9
1 9
2 9 12
2 9 12
4 12 5 9 12
4 12 5 9 12
2 9 12
2 9 12
4 12 5 9 12
4 12 5 9 12
5 12 5 9 9 12
8 9 1 9 2 12 5 2 12
4 9 1 9 12
4 9 1 9 12
6 9 1 9 9 7 9
3 1 0 12
2 9 12
2 3 12
16 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 12
18 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 12
4 13 15 13 2
18 7 13 1 15 2 16 15 13 1 3 0 2 16 4 13 1 9 2
9 7 13 2 9 2 9 7 13 2
9 0 9 2 9 2 0 9 2 9
7 0 2 11 2 9 16 9
5 9 12 2 12 2
25 11 12 2 0 9 1 9 2 0 12 2 15 1 9 7 9 9 2 12 2 2 12 2 12 2
40 13 0 9 7 9 2 0 2 9 2 2 0 9 11 2 12 12 11 12 2 0 12 2 9 2 2 2 12 2 12 12 2 9 2 2 12 2 12 12 2
20 11 2 9 2 11 2 0 9 0 7 0 9 2 12 2 2 12 2 12 2
48 13 0 9 7 9 2 0 2 9 2 2 12 12 11 12 2 9 12 2 9 2 2 2 12 2 12 12 2 9 2 2 12 2 12 12 2 12 12 2 12 12 2 9 2 12 12 9 2
33 11 2 9 9 11 2 10 9 2 10 9 2 9 2 9 2 9 2 0 9 2 9 2 0 9 2 12 2 2 12 2 12 2
29 13 9 11 2 12 12 11 2 1 9 12 2 9 2 2 2 12 2 12 2 12 2 9 2 2 12 2 12 2
23 11 2 0 9 7 0 9 2 12 2 0 0 7 0 9 2 12 2 2 12 2 12 2
21 13 0 9 9 11 2 12 12 11 2 0 12 2 9 2 2 2 12 2 12 2
5 9 12 2 12 2
67 9 2 11 2 11 1 11 2 11 2 11 1 0 9 2 11 2 11 2 11 2 9 11 2 11 2 11 2 0 11 2 11 2 9 11 9 2 11 2 0 9 2 9 2 11 2 11 12 2 9 2 11 2 11 2 11 2 11 2 9 2 11 1 11 2 11 2
29 0 9 2 11 2 9 9 2 11 2 11 2 9 1 9 2 11 12 2 11 2 9 11 2 1 12 9 2 2
5 9 12 2 12 2
66 9 2 11 1 11 2 0 11 2 11 2 9 2 11 2 9 0 9 2 9 11 2 11 2 11 2 11 2 9 0 9 2 11 2 0 9 2 11 12 2 9 2 11 1 11 2 11 2 11 2 9 1 9 2 11 2 11 1 11 2 9 9 9 2 11 2
5 9 12 2 12 2
17 11 12 2 9 9 2 0 9 0 9 12 2 2 12 2 12 2
38 13 11 11 2 11 2 11 2 9 11 5 11 2 9 2 0 2 9 2 9 12 2 12 12 11 12 2 9 2 2 9 2 2 12 2 12 12 2
3 9 12 2
24 11 12 2 9 9 2 9 7 9 2 12 2 9 0 9 2 9 2 9 2 9 9 2 2
34 13 0 11 11 2 12 12 11 12 2 0 12 2 9 2 2 2 12 2 12 2 12 2 9 2 2 9 2 2 12 2 12 12 2
1 11
17 0 9 0 9 1 9 7 9 9 1 0 9 13 1 9 12 2
25 13 1 9 12 9 7 13 9 12 9 9 2 13 11 11 2 9 0 9 11 2 1 9 2 2
29 0 9 9 13 1 0 11 1 11 2 0 9 13 9 1 11 2 0 0 11 2 11 2 7 11 2 11 2 2
23 3 16 12 5 9 13 1 9 2 3 1 0 9 0 2 11 2 1 0 7 0 9 2
19 1 11 13 0 9 9 11 1 9 12 9 0 0 9 2 9 2 0 2
32 9 9 7 9 9 2 15 13 0 3 1 9 2 15 13 1 11 1 12 9 9 1 9 12 1 12 9 9 1 0 9 2
35 1 12 1 9 9 0 0 11 11 13 0 9 13 9 9 7 0 9 2 3 0 9 11 12 7 11 12 2 0 9 1 11 7 0 2
21 0 9 13 9 1 11 3 13 2 16 13 0 9 1 0 9 16 1 0 9 2
35 9 2 0 0 9 2 9 2 0 2 2 9 2 11 2 11 12 2 12 2 12 12 11 12 2 9 2 2 9 2 2 12 2 12 2
5 9 13 1 0 9
11 1 9 3 16 1 9 2 10 3 0 9
42 1 10 9 9 11 13 3 3 1 9 2 13 15 11 1 9 7 13 15 2 10 9 2 7 7 15 3 3 13 10 9 7 9 13 14 1 9 2 15 15 13 2
26 0 9 15 3 3 15 13 1 15 1 9 7 9 2 16 9 13 3 0 7 0 2 16 9 13 2
9 9 4 3 13 1 0 9 9 2
6 13 1 15 7 3 2
2 11 11
13 9 13 2 16 14 12 9 10 0 9 13 0 2
13 1 15 13 1 9 10 9 1 9 0 9 11 2
7 13 15 7 14 1 11 2
25 1 9 11 11 2 9 0 9 11 2 11 2 9 13 2 16 10 9 13 0 7 1 0 9 2
45 13 15 3 2 16 1 0 0 9 2 15 13 12 9 2 13 0 9 12 9 2 0 2 0 9 12 9 7 9 2 3 9 9 2 7 7 9 1 9 1 9 2 12 9 2
17 13 15 2 3 13 9 2 13 0 9 2 3 13 9 0 9 2
3 16 9 13
6 13 15 0 0 9 2
14 3 0 9 13 3 9 9 2 13 1 9 2 13 2
23 9 2 16 10 9 13 3 2 15 3 13 13 13 9 2 13 2 13 9 2 13 9 2
35 13 3 1 12 9 1 0 2 3 15 13 1 9 7 9 2 3 13 9 2 16 15 13 7 15 13 13 3 2 3 15 3 9 13 2
11 7 3 1 0 9 13 13 9 1 9 2
27 3 9 13 13 2 9 2 9 2 9 2 13 7 1 0 9 16 9 7 9 2 1 15 13 13 3 2
9 16 10 9 13 1 9 15 0 2
3 7 13 2
3 7 3 2
16 7 1 9 13 0 0 9 16 1 9 2 3 10 0 9 2
58 0 13 7 9 2 0 9 2 9 2 15 13 1 10 9 0 9 7 9 9 2 7 13 3 0 9 2 2 0 9 7 0 0 9 2 1 10 9 9 2 2 0 0 9 2 0 9 2 15 15 4 15 13 2 2 0 9 2
50 9 1 9 13 2 3 15 15 1 10 9 1 0 0 9 13 2 0 9 2 9 2 12 5 2 0 9 7 0 0 9 12 5 2 0 9 12 5 2 0 0 9 12 5 2 0 9 12 5 2
20 3 0 9 15 13 3 13 7 15 13 2 16 3 0 9 7 0 0 9 2
3 9 14 9
15 2 0 9 2 1 9 13 15 2 15 15 1 15 13 2
11 7 9 0 9 3 1 10 10 9 13 2
6 0 9 13 0 9 2
26 0 13 1 9 1 9 2 0 3 9 15 9 7 9 2 9 1 9 2 9 0 9 9 7 3 2
47 0 13 0 9 9 2 16 3 15 13 9 2 0 13 0 9 2 9 15 13 9 3 13 2 7 15 9 1 15 3 13 2 9 13 13 7 13 9 2 15 13 1 9 13 15 0 2
23 1 0 9 13 13 7 13 7 15 2 1 15 15 13 9 2 3 13 1 0 9 0 2
31 3 9 9 0 9 2 1 15 13 12 12 9 0 9 2 3 3 1 15 9 13 2 7 13 10 9 2 15 15 13 2
25 0 0 9 13 2 16 12 5 0 0 9 13 12 5 9 2 16 12 5 9 13 12 5 9 2
23 3 12 5 9 9 13 0 9 2 9 16 3 9 9 2 15 7 13 14 12 5 9 2
11 15 9 13 3 3 13 9 1 0 9 2
24 9 13 0 9 10 9 13 0 9 2 15 1 15 13 3 9 0 9 2 9 9 2 9 2
16 3 3 9 4 13 13 9 2 7 16 3 15 15 13 13 2
5 15 13 7 9 2
61 9 11 13 2 16 0 0 9 13 13 3 2 12 9 0 9 2 0 2 2 12 9 0 2 9 1 0 9 2 2 12 9 9 2 9 2 9 2 9 0 9 2 0 9 2 2 12 5 9 2 9 9 2 9 9 7 9 3 2 2 2
21 0 9 2 1 9 2 2 1 15 15 13 9 0 0 9 2 13 12 5 9 2
30 0 12 5 13 0 9 2 1 15 15 13 3 9 0 1 9 2 1 9 2 1 9 2 7 7 9 3 15 13 2
2 9 9
21 9 10 9 1 9 0 7 0 9 13 13 0 9 2 0 2 7 3 15 15 2
19 13 15 13 2 16 13 13 14 3 1 9 0 9 7 16 0 10 9 2
25 1 15 13 3 13 9 2 13 15 9 2 15 13 13 15 0 2 15 9 13 0 9 7 9 2
15 15 7 13 13 9 2 15 13 13 2 10 13 13 9 2
21 7 13 1 9 2 15 15 13 9 13 3 2 16 4 13 0 2 0 2 0 2
25 11 11 7 11 11 1 10 9 9 13 1 0 2 7 7 0 9 13 2 0 9 7 0 9 2
6 0 7 3 0 9 2
8 0 9 2 3 13 15 0 2
6 9 2 9 7 9 2
6 0 9 7 0 9 2
3 0 9 2
5 13 15 0 9 2
15 7 1 9 9 7 10 0 9 1 0 7 13 3 13 2
18 3 3 2 15 13 1 15 2 10 9 15 9 13 7 3 15 13 2
26 11 11 1 11 2 11 13 2 16 1 9 10 9 13 13 3 9 1 9 1 9 1 14 9 9 2
9 1 10 9 13 13 3 10 9 2
22 9 3 13 2 16 9 15 1 15 4 13 3 2 16 15 13 9 2 9 7 9 2
13 7 3 15 15 4 1 10 9 13 7 13 9 2
18 9 9 13 2 16 15 9 2 7 1 15 7 10 9 2 13 3 2
13 9 0 9 1 0 3 13 15 0 9 7 9 2
46 13 15 3 13 2 16 0 9 13 3 13 14 1 15 2 3 3 2 3 1 0 9 2 13 2 7 1 15 2 3 3 13 13 10 9 7 13 0 9 0 9 1 3 0 9 2
3 9 1 9
11 0 9 1 9 2 9 9 1 15 13 9
17 9 0 0 7 0 9 7 3 0 9 9 9 11 13 9 9 2
30 9 15 3 13 2 16 13 10 9 1 9 2 7 15 3 3 2 16 13 9 2 16 9 1 9 3 13 13 3 2
2 11 11
26 16 15 3 13 9 3 0 0 9 2 13 4 15 10 12 9 2 0 9 0 0 9 7 0 11 2
3 0 15 13
9 13 11 11 2 0 9 2 11 2
10 2 3 13 9 12 9 14 10 9 2
7 13 1 10 9 0 9 2
34 3 1 9 1 0 9 0 9 1 0 7 0 9 15 13 2 16 1 9 13 0 9 0 9 7 13 1 0 9 1 0 9 13 2
7 10 9 13 1 0 9 2
22 3 13 9 9 2 15 2 16 4 15 13 0 9 2 13 10 9 1 9 13 9 2
12 15 15 7 1 9 1 9 1 0 9 13 2
9 2 13 4 0 9 10 9 9 2
6 3 2 7 13 9 2
16 15 13 1 9 1 9 0 7 0 9 2 0 1 0 9 2
24 13 1 15 0 9 12 9 9 2 7 0 4 13 0 9 10 0 9 7 3 1 15 13 2
13 15 7 13 0 2 10 9 4 0 9 3 13 2
2 14 2
13 13 2 14 15 13 3 3 2 13 3 0 9 2
29 10 9 0 9 4 3 0 13 1 0 9 2 7 13 1 15 14 9 9 7 3 15 15 13 0 9 13 9 2
12 2 1 10 9 9 11 13 9 1 9 3 2
17 9 13 1 0 9 16 1 9 2 15 13 9 9 1 10 9 2
19 9 0 7 0 9 9 3 3 13 2 16 1 15 9 1 9 13 9 2
8 3 13 1 9 9 7 9 2
34 1 11 15 13 15 0 2 15 13 9 9 2 13 1 15 3 2 13 0 9 2 7 3 13 3 1 9 2 16 1 3 0 9 2
26 7 13 9 2 1 9 15 9 2 0 7 0 2 15 3 3 9 13 13 2 16 1 10 9 13 2
13 2 3 1 10 9 13 13 9 9 9 16 9 2
20 7 13 0 9 2 16 4 15 13 13 1 0 7 0 2 0 7 0 9 2
9 9 9 1 3 0 9 3 13 2
17 13 15 0 15 2 16 16 15 3 13 2 15 15 13 14 9 2
17 2 2 2 2 13 1 9 2 15 15 2 14 2 13 1 9 2
23 9 0 9 7 9 2 16 15 2 9 2 13 15 1 12 9 2 3 3 13 3 3 2
18 7 13 3 9 0 0 9 7 0 0 9 2 13 3 1 0 9 2
10 0 2 15 15 13 2 13 9 9 2
24 1 9 9 13 0 2 16 9 9 9 1 0 9 4 13 3 3 13 0 2 16 0 9 2
45 7 13 9 2 16 12 0 9 13 0 9 1 9 9 7 0 12 9 15 13 2 13 10 9 0 2 16 1 9 12 1 12 9 2 3 0 9 2 4 9 3 13 3 15 2
2 0 9
32 15 13 9 9 0 9 2 0 3 3 15 2 16 9 10 9 13 9 13 0 9 9 11 2 16 1 15 3 13 15 0 2
10 7 9 10 0 9 11 11 13 0 2
7 2 3 13 9 0 9 2
22 9 9 1 11 13 0 9 2 15 13 9 9 7 9 1 9 1 9 15 3 13 2
18 0 9 1 11 13 3 0 2 7 15 2 15 13 2 3 13 9 2
14 13 13 3 0 9 2 3 10 9 2 15 13 9 2
19 2 9 13 2 16 3 15 3 13 1 15 2 15 15 3 0 9 13 2
13 15 15 15 13 16 9 9 2 0 1 9 9 2
14 3 15 13 16 9 3 1 9 2 7 15 13 9 2
4 2 13 15 2
28 16 3 4 13 12 12 9 2 0 1 9 7 10 9 4 15 13 0 9 13 2 7 3 1 10 9 13 2
29 15 13 3 9 0 9 1 9 2 3 12 0 9 13 1 0 9 0 9 9 7 9 1 15 7 0 15 13 2
8 2 10 9 10 9 13 13 2
18 1 0 9 13 13 14 1 9 9 1 10 9 2 15 10 9 13 2
21 7 15 13 9 2 3 13 0 10 9 3 13 7 0 0 9 0 0 9 13 2
10 3 14 9 13 0 9 9 7 9 2
20 15 0 4 13 3 9 1 15 2 16 13 0 9 7 7 3 0 0 9 2
5 9 2 13 4 13
3 1 0 9
18 0 9 15 13 0 9 0 9 2 16 13 15 2 15 13 1 9 2
8 1 15 13 13 9 10 9 2
9 9 0 9 9 13 0 0 9 2
25 3 1 0 9 13 9 12 12 2 12 7 10 9 12 2 12 2 12 2 12 2 12 2 12 2
28 1 15 15 13 9 0 2 0 9 2 9 2 9 2 9 2 0 0 0 9 2 0 9 2 9 7 9 2
7 9 13 1 15 10 9 0
3 0 9 2
5 0 9 13 13 2
2 0 2
20 0 2 15 13 0 9 7 9 2 0 2 0 2 1 9 9 7 9 2 2
8 0 9 2 1 0 9 2 2
18 0 2 0 9 7 0 9 9 1 2 9 0 9 1 9 9 2 2
11 1 0 0 9 2 1 0 9 7 9 2
18 1 0 9 3 9 13 9 2 1 15 15 0 9 13 1 0 9 2
1 3
3 0 9 2
8 1 9 15 13 1 12 9 2
35 1 12 2 9 15 13 9 0 3 0 0 9 2 16 13 0 2 1 0 9 2 1 9 0 1 0 9 2 3 0 2 1 0 9 2
15 0 9 13 13 7 3 0 1 9 9 1 9 1 9 2
14 1 9 2 9 2 9 2 13 13 3 14 12 9 2
18 1 0 2 0 7 0 9 1 9 1 12 9 13 13 9 3 0 2
26 1 12 2 9 15 13 9 0 0 9 2 0 2 13 13 7 3 0 9 7 0 9 9 9 9 2
11 9 13 13 7 3 0 2 14 7 0 2
14 13 15 0 9 3 0 1 9 9 1 9 1 9 2
15 1 0 2 0 7 0 9 13 13 9 3 0 2 0 2
29 1 12 0 9 13 2 16 0 0 9 13 13 9 9 2 9 7 9 1 9 0 9 2 9 7 0 13 13 2
9 9 15 13 3 12 9 1 9 2
25 1 0 9 15 1 0 9 13 1 12 2 9 9 3 12 9 2 1 12 2 9 3 12 9 2
18 0 9 0 13 13 1 12 2 7 1 12 2 9 9 3 12 9 2
33 1 9 1 0 9 2 7 1 0 9 2 15 13 1 12 2 9 3 12 5 9 9 9 7 9 7 9 0 1 12 2 9 2
30 1 0 9 15 13 3 12 5 9 9 0 0 9 2 7 9 0 2 7 9 9 14 1 12 5 0 16 13 13 2
2 11 11
5 1 9 15 9 13
3 16 13 9
15 1 9 4 15 13 1 12 0 9 0 0 9 1 9 2
26 10 0 9 13 1 9 2 16 15 1 9 0 9 9 13 2 16 9 13 9 1 9 0 9 13 2
15 13 15 3 1 9 9 1 9 2 15 9 9 3 13 2
25 16 4 15 3 3 13 2 16 9 13 1 9 1 9 0 2 13 15 0 9 1 9 7 9 2
13 1 10 9 4 15 1 9 9 9 13 0 9 2
21 13 4 9 2 16 9 3 13 10 9 1 0 0 9 2 16 10 9 13 0 2
11 0 0 0 9 13 0 2 3 7 15 2
17 9 1 9 3 13 7 13 15 1 0 9 1 9 1 0 9 2
21 10 9 4 15 13 7 13 9 13 13 0 0 9 1 0 9 7 1 0 9 2
28 7 16 4 15 1 15 13 2 3 14 4 15 3 13 2 16 10 9 13 1 0 9 2 7 1 0 9 2
7 9 9 15 13 3 13 2
12 10 10 9 1 9 13 14 1 9 7 9 2
17 1 0 9 7 1 9 13 9 0 2 1 9 1 9 3 15 2
42 7 3 4 15 13 0 9 2 16 4 15 3 13 2 3 13 13 0 9 0 0 9 2 16 9 2 0 9 7 9 1 0 7 0 9 1 0 9 2 9 9 2
22 7 3 15 2 15 15 15 1 9 13 1 0 9 2 15 3 13 9 7 0 9 2
2 9 2
18 2 13 2 16 0 9 13 1 9 1 15 2 3 4 9 9 13 2
15 2 1 9 1 9 13 0 13 0 9 7 9 0 9 2
7 11 2 11 2 2 0 11
23 9 2 0 1 10 9 2 0 1 0 9 9 2 4 3 13 7 3 13 9 12 9 2
10 4 3 13 1 0 9 1 12 9 2
17 13 15 2 15 9 4 15 1 9 13 7 10 1 15 13 9 2
2 9 9
25 1 0 9 9 9 1 9 13 0 9 2 12 5 9 2 1 9 0 9 9 2 9 7 9 2
17 0 0 9 13 9 1 9 7 0 9 2 15 13 3 12 5 2
15 9 1 9 2 7 2 9 2 9 2 9 13 12 5 2
19 1 0 0 9 2 15 9 13 2 15 13 1 0 0 9 9 12 9 2
4 2 0 9 2
2 9 9
11 1 9 12 4 13 13 1 9 0 9 2
15 1 0 9 1 9 12 4 13 1 12 5 9 9 9 2
20 14 1 9 12 4 13 0 9 2 1 15 15 15 13 14 12 5 9 9 2
18 4 15 13 2 16 1 9 12 7 12 4 13 9 1 9 1 9 2
19 13 15 2 16 0 9 1 9 9 9 13 2 16 0 9 13 0 9 2
19 0 9 4 13 1 9 2 16 9 13 1 9 7 9 0 9 4 13 2
4 11 11 2 11
14 9 1 9 9 9 1 9 12 5 13 1 10 9 2
46 16 4 1 9 12 13 0 9 1 3 0 9 9 2 12 2 12 9 2 1 9 1 9 9 2 13 2 1 2 0 2 9 2 13 0 9 9 2 16 4 13 9 1 0 9 2
26 9 2 11 11 2 0 9 2 0 12 2 12 12 11 12 2 9 2 2 2 12 2 12 12 12 2
3 9 2 9
5 9 1 9 1 11
15 9 3 13 12 12 9 1 9 0 9 7 1 10 9 13
6 3 4 13 3 9 2
14 0 4 15 13 7 13 3 2 16 4 15 13 9 2
20 13 15 2 16 4 1 15 13 13 3 9 2 16 3 3 14 13 0 9 2
4 11 9 2 11
2 11 11
22 9 0 1 9 13 3 13 1 9 2 16 10 9 4 13 1 0 9 1 0 9 2
15 7 13 3 9 2 16 1 9 13 0 9 0 0 9 2
7 13 15 7 7 1 15 2
2 3 13
7 9 1 9 9 13 0 2
18 1 9 13 15 9 9 1 9 1 0 9 2 0 9 2 0 9 2
34 3 0 9 7 9 13 13 0 9 1 9 0 9 2 16 0 9 2 15 13 1 9 9 0 9 3 13 1 9 2 13 13 9 2
24 0 9 9 1 9 13 3 0 11 2 0 0 11 2 0 11 2 0 0 11 2 0 11 2
13 3 13 13 2 0 9 2 1 11 7 1 11 2
5 9 2 1 9 2
26 13 4 0 13 1 0 9 1 9 1 9 2 7 13 10 9 2 3 4 10 9 0 9 13 13 2
10 7 13 3 2 16 0 9 15 13 2
16 3 13 1 9 7 13 15 9 13 0 7 1 0 0 9 2
14 9 1 10 0 9 13 14 9 7 13 15 1 0 2
25 0 9 0 2 9 2 1 0 9 3 13 7 12 15 1 15 13 2 15 7 10 9 3 13 2
6 0 11 2 11 2 9
48 0 9 2 0 1 9 2 4 9 11 13 0 9 16 3 11 2 12 1 10 0 9 13 1 9 1 9 2 7 0 11 9 2 9 2 0 2 2 1 10 9 1 0 9 1 11 2 2
15 9 13 3 7 9 9 11 2 0 9 2 3 11 2 2
27 10 9 4 3 2 13 13 7 1 9 2 3 13 9 9 9 11 2 15 13 7 13 9 0 1 11 2
20 13 4 15 13 2 16 10 9 2 3 0 9 2 3 13 9 2 3 9 2
4 7 3 9 2
6 1 9 15 3 13 2
17 13 15 0 9 12 9 2 15 3 13 9 1 9 0 0 9 2
16 1 10 0 9 3 13 12 0 9 7 13 15 9 1 9 2
30 16 15 0 13 0 2 16 15 0 9 13 2 16 9 13 9 2 13 3 2 16 1 0 9 15 9 13 9 13 2
24 9 13 1 15 2 16 0 9 0 9 13 9 9 2 16 9 13 15 0 2 16 9 9 2
25 16 1 9 15 0 9 2 15 1 12 2 9 13 9 11 2 13 13 9 7 13 13 1 9 2
4 1 9 7 9
34 9 1 10 9 13 0 2 13 14 3 2 3 13 9 2 3 9 1 9 9 2 15 13 13 9 7 9 0 9 1 9 0 9 2
21 7 13 13 15 2 16 15 2 15 13 1 9 0 16 0 9 2 15 3 13 2
9 9 15 1 10 9 9 9 13 2
36 3 0 9 2 16 13 9 2 13 1 9 2 3 9 13 0 1 0 9 3 1 9 2 1 15 13 9 12 1 12 3 0 9 0 9 2
19 0 13 3 0 9 11 2 0 11 1 9 2 2 10 9 13 1 9 2
8 0 13 0 9 11 7 11 2
9 1 0 9 13 9 0 0 9 2
20 10 9 9 15 3 13 0 7 4 13 1 0 9 7 16 15 13 0 9 2
18 16 2 0 2 9 4 13 12 5 2 1 0 4 13 12 5 9 2
18 1 9 4 9 11 9 1 0 9 1 11 9 13 11 7 0 11 2
15 3 0 9 4 13 14 12 9 1 9 1 9 12 9 2
6 1 0 9 15 13 2
3 9 12 9
20 0 9 13 9 2 16 1 9 13 13 12 9 2 15 4 13 3 0 9 2
10 13 7 0 9 7 9 1 9 9 2
28 0 9 13 0 2 12 9 2 9 2 9 2 2 9 2 9 2 2 9 2 9 2 7 9 2 9 2 2
9 13 15 9 2 15 13 9 9 2
30 13 15 13 14 0 9 2 15 1 15 13 3 0 9 2 7 7 3 13 9 2 3 1 0 9 2 3 0 9 2
4 0 13 1 9
12 1 0 9 15 13 1 0 9 9 10 9 2
31 0 9 7 0 9 2 9 2 13 9 0 9 2 3 1 9 1 9 1 12 7 0 9 13 13 10 9 1 10 9 2
23 9 2 9 2 0 2 9 13 9 2 15 13 9 1 9 2 15 15 13 1 9 9 2
14 9 13 9 1 10 9 2 10 9 13 13 0 9 2
6 9 9 3 13 3 2
3 0 13 0
6 3 15 13 9 0 2
14 9 13 3 15 2 16 0 13 9 7 13 1 0 2
12 0 9 13 1 9 0 2 0 7 3 0 2
15 9 2 15 4 13 1 9 3 0 2 15 3 9 13 2
10 3 13 3 3 0 9 2 9 2 2
20 0 9 9 7 1 9 13 10 9 2 7 9 9 13 2 3 13 9 0 2
16 0 9 13 1 15 3 0 2 16 10 9 13 0 13 3 2
8 0 9 13 1 0 9 0 2
20 1 9 9 2 9 13 0 9 9 2 0 2 0 2 0 2 0 2 0 2
3 0 13 0
9 9 15 13 1 9 1 12 9 2
8 9 1 12 3 15 13 3 2
29 9 9 0 9 2 9 2 9 12 2 3 0 9 2 1 9 12 9 15 3 13 1 12 2 12 9 2 9 2
11 9 13 2 16 1 9 9 13 9 3 2
6 13 4 13 10 9 2
10 9 9 9 5 9 12 9 5 9 12
15 3 12 0 9 4 3 13 12 2 12 5 12 12 2 2
26 9 13 3 0 2 12 0 9 0 9 13 1 0 0 9 11 7 9 1 9 14 12 9 2 9 2
22 13 15 13 15 2 16 1 9 1 0 9 13 9 2 15 15 13 2 13 0 9 2
4 3 0 1 9
29 1 9 9 7 9 9 14 15 2 16 10 9 13 9 1 12 1 12 9 2 3 0 2 0 2 0 2 0 2
28 4 13 9 9 10 9 2 7 4 15 13 3 0 2 3 0 7 1 9 2 15 15 13 9 9 3 0 2
4 11 13 0 9
20 1 9 15 1 9 13 1 9 2 15 15 13 1 15 1 0 3 0 9 2
12 12 1 15 13 3 11 2 15 13 12 3 2
26 1 15 13 9 9 1 0 9 1 12 9 1 12 9 2 9 0 9 13 0 2 1 15 9 9 2
16 11 7 0 11 13 1 11 1 9 0 9 9 1 0 9 2
25 1 11 13 13 2 16 0 9 9 9 1 0 9 13 1 9 9 14 1 12 0 9 1 9 2
9 9 0 9 0 9 13 3 0 2
23 9 1 10 9 0 2 16 13 11 2 13 9 0 9 7 3 3 0 9 13 0 11 2
2 9 9
24 3 13 9 9 9 2 10 9 2 15 4 13 9 9 2 16 4 15 13 13 1 0 11 2
22 0 9 2 9 9 7 9 9 12 2 3 1 0 9 2 13 1 0 11 12 9 2
18 1 9 2 16 13 1 9 1 9 11 2 13 12 5 9 12 9 2
45 0 9 2 10 9 1 9 11 11 1 0 11 13 1 9 9 2 1 0 9 13 13 12 5 7 1 0 3 14 12 5 2 2 1 10 9 13 12 5 2 3 14 12 9 2
20 13 15 1 12 9 7 13 0 9 1 0 9 2 12 5 9 2 12 9 2
22 13 2 14 9 12 9 1 9 2 10 9 4 13 1 9 2 13 9 7 12 9 2
12 1 11 4 9 9 13 0 9 1 15 3 2
40 13 4 1 15 14 12 9 2 9 2 13 2 14 15 1 9 4 15 9 13 14 12 9 2 2 16 1 9 9 13 1 11 12 5 9 1 15 9 2 2
23 11 13 9 1 11 1 12 5 9 2 16 15 9 2 0 9 7 9 13 1 0 9 2
20 3 10 9 13 3 0 9 2 7 10 9 2 3 0 13 14 13 1 9 2
13 3 3 15 1 15 13 9 1 9 1 12 9 2
36 1 11 3 13 12 0 9 2 9 9 2 3 0 7 0 9 7 9 9 12 2 1 9 12 9 2 1 9 9 15 13 1 12 9 2 2
41 0 9 13 3 14 12 5 2 7 13 3 13 15 2 16 11 15 13 13 1 9 11 16 15 2 15 9 13 2 3 9 0 9 13 2 13 3 9 7 9 2
5 9 7 9 3 1
31 10 9 13 3 9 1 15 2 3 4 13 13 2 7 0 13 7 0 9 9 2 15 15 13 2 4 2 14 13 13 2
10 9 1 12 9 13 11 1 0 9 2
11 1 0 9 7 13 2 16 4 13 9 2
25 3 1 15 13 1 9 9 2 1 15 15 13 2 7 1 9 2 7 13 15 10 9 1 9 2
14 13 2 14 9 9 3 2 13 15 13 1 9 0 2
15 11 13 9 2 1 15 13 0 9 13 3 1 0 9 2
15 1 0 11 4 9 13 1 0 9 1 11 0 0 9 2
19 3 9 2 0 9 7 9 2 15 13 9 1 9 2 13 9 13 3 2
25 15 2 15 4 15 0 11 1 9 13 2 4 13 1 0 9 0 2 16 4 9 9 3 13 2
20 1 9 4 7 13 0 13 1 0 9 2 16 4 13 0 9 9 0 9 2
45 16 3 1 0 0 9 9 1 12 9 1 9 4 10 9 13 9 2 15 13 1 12 9 2 1 12 7 9 9 13 1 12 9 2 12 5 12 5 12 7 13 1 9 2 2
7 7 9 0 13 3 0 2
34 1 0 9 13 7 13 2 16 3 2 16 13 13 0 9 2 4 13 7 1 15 13 1 9 1 9 2 3 13 9 9 7 9 2
19 3 13 0 1 0 9 2 1 0 0 9 2 13 9 9 9 1 9 2
21 10 9 4 13 13 2 16 0 0 9 13 2 15 13 2 7 13 0 9 9 2
22 16 13 0 9 2 16 13 15 1 9 2 3 4 9 9 9 1 9 13 13 0 2
13 3 1 0 0 9 2 7 3 16 9 1 9 2
5 9 7 9 0 9
12 13 15 1 9 2 13 4 15 7 3 7 13
17 16 0 1 10 9 1 9 0 9 13 1 9 9 9 0 9 2
11 16 4 15 13 2 13 13 1 0 9 2
13 0 9 9 1 11 13 1 9 0 9 1 9 2
10 1 10 9 15 7 13 3 3 13 2
2 11 11
22 1 0 9 1 9 0 9 13 9 9 10 9 2 13 9 2 13 9 1 0 9 2
9 0 9 13 0 9 1 0 9 2
13 1 15 13 1 9 9 9 2 15 13 10 9 2
14 2 0 0 9 1 0 9 13 9 7 13 15 9 2
11 3 9 13 9 1 0 9 1 10 9 2
8 15 13 0 9 1 9 9 2
10 15 15 13 1 11 9 7 13 0 2
11 10 9 13 10 9 1 10 9 0 9 2
19 9 9 13 1 9 2 3 3 13 1 10 9 13 10 0 9 1 9 2
12 15 15 13 13 3 14 1 9 9 1 9 2
2 0 9
30 2 1 9 9 15 13 1 10 9 9 2 1 9 15 13 1 15 13 9 2 13 9 1 9 7 13 0 9 9 2
18 1 9 9 9 11 9 13 2 1 0 9 12 9 4 13 13 9 2
5 3 13 12 9 2
4 13 12 9 2
18 7 3 9 13 9 2 7 1 0 3 12 9 15 9 3 13 12 2
12 9 1 15 13 2 7 3 3 13 1 9 2
29 16 13 1 9 7 3 13 7 0 9 2 9 7 0 0 9 7 0 9 1 9 2 13 15 3 9 10 9 2
7 11 9 13 2 13 9 2
4 14 15 13 2
6 13 4 1 15 9 2
25 13 3 9 1 15 2 3 13 9 2 13 9 2 13 3 9 2 3 13 9 7 13 0 9 2
12 2 9 0 9 13 1 9 0 9 0 9 2
14 13 15 13 9 2 15 1 0 9 2 3 0 9 2
16 0 13 3 2 1 9 2 13 1 0 9 7 13 0 9 2
20 1 10 9 13 0 2 16 4 13 0 9 3 3 16 12 5 9 9 9 2
3 13 15 9
30 1 0 9 1 9 0 9 13 9 7 1 0 0 9 2 1 9 0 9 1 9 9 2 0 9 1 0 0 9 2
7 15 13 7 3 0 9 2
35 1 9 2 15 11 13 2 7 1 9 2 15 13 2 3 15 13 3 1 0 9 13 2 3 12 2 2 13 0 13 14 12 9 3 2
25 13 4 2 16 13 9 13 15 12 9 2 16 0 0 9 12 13 2 7 13 4 9 15 13 2
26 2 16 4 15 1 0 9 13 1 9 3 9 2 13 0 13 9 2 7 2 13 1 9 9 2 2
13 1 9 0 9 4 3 13 0 10 9 3 13 2
5 0 9 13 9 2
25 9 13 2 16 1 9 9 9 13 3 7 15 2 16 3 13 13 9 1 0 9 1 0 9 2
9 0 15 7 13 0 9 1 15 2
17 1 9 0 0 9 1 9 13 2 0 9 13 13 9 12 9 2
22 1 9 3 13 2 16 13 4 13 15 2 9 13 1 9 13 2 7 0 9 13 2
8 3 0 9 13 14 0 9 2
7 1 0 9 10 9 3 2
11 2 3 0 9 13 1 3 0 9 9 2
18 1 10 9 15 13 0 2 3 13 9 2 0 15 1 9 1 9 2
3 9 13 9
19 16 4 15 13 2 16 0 9 13 1 9 0 9 2 13 15 3 9 2
35 16 9 11 9 13 1 9 13 1 9 12 9 9 1 9 1 9 7 1 9 2 16 9 13 3 9 2 13 15 2 9 13 0 9 2
14 13 0 9 2 7 15 13 0 9 7 13 15 13 2
29 3 13 9 13 2 16 13 14 1 0 9 2 16 4 11 13 9 2 3 13 13 9 7 9 2 16 13 9 2
16 3 13 1 9 0 9 2 16 13 2 16 13 3 0 9 2
6 9 7 9 0 9 2
3 5 2 2
7 2 0 9 1 0 9 2
5 2 3 0 9 9
9 2 0 9 2 1 9 2 9 2
5 2 2 9 9 9
6 2 3 0 9 2 2
2 9 9
6 2 1 9 9 0 2
16 2 1 9 9 9 1 9 3 1 0 9 2 9 9 9 10
2 2 9
5 2 2 3 15 0
4 2 9 1 9
5 2 2 9 9 2
5 9 1 9 2 2
14 9 1 9 2 1 0 9 15 13 0 1 10 9 2
2 10 9
8 15 15 13 2 0 2 2 2
8 2 9 9 2 12 2 12 2
30 1 9 9 0 9 13 13 2 16 2 1 9 9 9 0 7 0 9 15 13 3 13 9 0 9 1 9 9 2 2
14 13 13 2 16 15 4 13 0 9 9 1 0 9 2
38 14 3 3 0 9 7 0 9 13 9 1 9 0 9 1 9 11 1 0 9 9 7 9 0 13 9 0 9 1 9 12 2 9 2 12 0 9 2
37 9 9 1 0 9 1 9 0 9 4 13 7 9 9 1 9 9 9 2 12 2 12 2 15 1 10 9 13 7 9 0 9 1 9 9 13 2
10 9 1 0 9 4 3 3 13 10 2
27 1 9 9 0 9 1 0 9 4 13 9 9 1 9 0 9 2 15 7 9 1 9 1 10 9 13 2
37 9 4 13 7 1 10 9 0 2 16 4 1 0 9 4 13 1 0 9 2 7 2 13 13 9 1 9 7 9 1 0 9 14 1 9 11 2
39 7 1 0 9 15 13 13 2 16 13 13 9 12 2 9 2 12 0 9 2 1 15 9 13 13 1 10 9 1 0 9 7 1 0 9 16 0 9 2
4 11 13 2 11
3 13 15 9
17 13 1 0 9 1 0 9 7 13 2 16 15 15 1 9 13 2
5 3 15 9 13 2
6 13 1 9 0 9 2
24 9 13 2 16 13 0 2 3 15 15 13 7 13 2 16 9 13 13 2 16 15 13 9 2
18 13 2 16 3 10 9 15 1 10 9 15 15 1 9 13 1 9 2
7 15 4 13 13 2 13 2
15 13 9 15 13 7 13 1 9 2 16 3 3 3 13 2
13 1 0 9 2 3 0 2 13 1 0 9 3 2
14 9 15 1 0 9 1 9 1 9 7 9 9 13 2
11 7 15 13 2 16 4 13 10 10 9 2
6 11 11 2 9 1 11
4 9 1 0 9
8 2 9 9 2 12 2 12 2
35 1 0 9 4 13 9 1 10 9 2 0 9 4 1 0 9 1 11 13 1 12 9 2 15 13 3 0 9 1 0 7 0 9 0 2
19 9 13 3 2 1 9 7 9 13 2 16 13 1 9 0 9 0 9 2
26 1 9 1 11 2 11 1 0 9 13 15 9 2 15 13 1 9 0 9 7 9 0 9 1 9 2
11 1 10 9 13 1 9 9 1 12 9 2
15 0 4 1 9 9 1 0 9 13 0 9 7 0 9 2
12 15 0 15 13 2 16 4 9 13 3 3 2
12 1 9 2 15 0 9 9 13 2 15 13 2
3 11 11 2
7 3 0 9 0 9 2 11
4 9 1 11 13
8 2 9 9 2 12 2 12 2
11 9 0 9 13 3 1 9 15 0 9 2
17 0 7 0 9 2 15 13 9 10 9 1 0 9 2 13 9 2
15 1 9 15 13 1 15 7 9 9 2 9 2 9 9 2
17 1 15 15 13 9 2 16 3 1 15 10 9 1 3 0 13 2
19 3 7 3 2 16 3 1 10 9 1 9 15 1 0 9 13 0 9 2
24 3 13 0 9 0 1 0 9 1 0 9 15 2 3 13 3 0 9 13 9 9 1 9 2
22 3 3 0 9 7 9 3 13 2 16 1 0 7 3 0 9 13 10 9 13 3 2
21 9 0 9 13 13 16 9 2 16 9 1 9 15 14 13 2 7 7 13 9 2
4 1 9 13 9
8 2 9 9 2 12 2 12 2
23 0 9 2 3 15 13 9 13 7 15 9 13 2 16 13 3 9 9 2 13 3 0 2
14 13 15 3 9 1 0 9 1 9 0 9 1 9 2
15 3 1 9 2 9 15 13 7 0 9 7 3 15 13 2
17 10 0 9 2 15 13 9 7 3 7 10 9 2 13 3 9 2
37 9 13 1 15 2 16 9 13 0 7 9 1 0 0 9 2 15 15 15 14 1 9 13 2 7 0 3 0 9 1 0 9 2 13 3 0 2
4 11 11 2 11
3 9 7 9
8 2 9 9 2 12 2 12 2
16 1 0 9 13 0 9 2 15 13 13 1 9 9 2 9 2
17 16 4 15 13 13 9 1 12 9 2 15 3 4 1 9 13 2
12 13 15 7 2 16 9 0 9 13 0 3 2
23 16 13 10 0 2 15 9 1 0 9 13 2 13 0 0 9 1 9 13 1 0 9 2
4 11 11 2 11
4 2 0 9 2
4 11 13 1 0
8 0 9 15 13 9 1 9 2
25 1 12 0 15 13 7 0 9 2 15 13 12 2 9 12 3 16 0 9 0 0 7 0 9 2
20 12 1 0 9 9 3 15 9 2 7 3 7 0 2 13 9 9 1 9 2
21 0 9 2 9 2 9 9 1 0 0 9 2 0 9 2 15 15 3 0 13 2
43 12 1 0 9 13 7 11 2 0 11 12 2 0 1 9 1 0 9 1 0 9 0 11 2 11 2 15 15 13 12 2 7 12 2 12 2 12 1 9 9 1 11 2
30 13 15 3 0 7 0 9 1 9 9 2 9 2 0 7 0 9 2 9 2 9 2 9 2 9 0 9 7 0 2
20 9 9 13 7 0 9 1 9 2 9 7 9 2 9 0 9 2 0 9 2
14 12 1 0 9 0 9 11 15 13 1 9 1 9 2
17 13 1 9 2 9 2 1 10 9 13 7 9 1 9 7 9 2
25 1 0 9 13 9 0 13 0 9 1 9 0 9 1 11 2 3 9 0 1 9 9 1 11 2
14 3 1 9 0 9 13 9 9 1 9 9 1 11 2
17 1 9 10 9 13 9 1 9 13 1 10 9 9 1 9 9 2
21 10 9 13 9 1 15 9 1 9 15 2 3 15 13 9 9 12 7 9 12 2
13 3 9 13 9 9 1 9 2 15 4 3 13 2
16 9 3 13 9 13 9 1 9 0 9 2 15 15 13 9 2
18 9 9 13 0 13 0 9 9 9 1 0 9 2 9 2 7 3 2
24 0 0 9 13 13 1 9 11 1 2 11 2 15 13 0 0 9 1 11 7 13 3 13 2
24 9 1 0 9 1 9 13 10 9 2 9 9 2 0 9 2 9 9 2 9 2 9 9 2
23 1 15 9 13 13 0 9 1 9 2 1 0 9 7 10 9 2 1 9 9 7 9 2
2 11 0
37 9 2 0 0 9 11 2 0 12 2 12 12 11 12 2 9 2 2 2 12 2 12 2 12 2 12 2 12 2 9 2 2 12 2 12 12 2
3 9 13 9
10 0 9 13 3 7 15 13 7 13 9
30 1 9 1 12 1 9 1 0 9 12 2 9 13 0 9 2 16 1 9 0 9 0 9 13 9 3 3 0 9 2
7 9 13 1 9 9 9 2
14 9 15 3 9 3 7 13 2 13 15 0 11 11 2
9 0 7 13 2 16 13 1 9 2
19 3 13 9 0 9 7 9 15 13 1 9 2 13 2 15 3 3 13 2
18 9 9 15 13 3 14 14 1 12 9 2 7 3 13 9 0 9 2
3 1 9 9
26 1 9 9 4 0 13 13 2 15 15 13 1 9 13 3 1 9 7 1 9 7 15 1 0 9 2
21 1 9 9 15 13 0 9 0 9 2 0 3 7 1 9 1 9 7 1 9 2
13 1 10 9 3 13 1 0 9 9 1 0 9 2
10 7 3 0 9 2 3 3 1 9 2
8 1 9 13 1 9 9 9 2
11 15 1 9 2 7 9 13 0 13 3 2
15 0 2 0 1 9 3 1 9 2 15 13 13 7 3 2
19 0 1 0 13 1 10 9 0 2 9 1 9 15 13 13 1 3 9 2
6 9 13 3 3 0 2
6 0 9 13 0 9 2
13 3 13 3 13 15 2 15 4 1 15 13 9 2
20 9 13 9 2 10 9 13 13 1 9 2 1 9 2 1 9 2 7 9 2
14 3 13 9 2 10 13 9 2 15 15 13 2 13 2
15 1 9 13 0 9 7 1 0 9 2 3 1 0 9 2
5 13 15 0 0 2
20 0 9 13 7 1 15 15 13 0 2 15 1 0 9 2 3 9 7 9 2
3 9 15 13
20 7 1 9 15 0 9 9 9 2 3 9 2 9 2 9 2 13 9 9 2
7 15 3 13 1 9 9 2
18 13 1 15 9 9 0 7 0 9 7 9 9 1 0 9 7 9 2
7 9 7 9 13 0 9 2
7 7 15 7 13 0 9 2
12 0 9 3 13 14 12 2 7 3 12 9 2
12 1 0 9 9 9 13 2 3 15 13 13 2
19 16 12 9 13 1 0 9 9 1 9 9 2 0 13 13 1 15 12 2
8 3 15 15 13 7 10 9 2
5 9 2 9 2 9
9 7 1 9 15 13 13 1 9 2
11 1 15 9 11 13 9 1 9 0 9 2
12 3 13 15 10 9 2 3 9 7 0 9 2
13 13 15 13 3 1 9 9 2 15 0 9 13 2
24 3 15 15 15 13 3 2 16 9 1 0 9 2 9 11 15 9 13 2 13 3 1 9 2
6 13 1 9 0 9 2
7 13 9 2 7 14 3 2
7 13 0 13 0 0 9 2
11 1 9 2 15 13 3 9 2 13 9 2
16 3 1 9 13 1 9 1 9 12 2 9 0 9 10 9 2
14 15 2 1 15 15 13 9 9 2 3 13 1 9 2
16 13 0 13 15 3 7 1 9 0 9 2 16 13 0 9 2
11 0 9 4 13 0 9 7 9 1 9 2
13 1 0 9 0 9 13 7 1 0 9 0 9 2
20 3 0 0 2 0 9 15 13 0 9 9 1 9 7 3 1 15 13 9 2
9 9 15 7 13 3 1 0 9 2
8 3 3 9 13 0 0 9 2
11 13 1 3 0 9 2 15 15 3 13 2
12 13 3 4 13 9 9 7 10 9 1 9 2
2 11 0
25 9 2 9 2 9 2 9 12 2 9 2 12 12 11 12 2 9 2 2 2 12 2 12 12 2
3 9 1 12
16 3 9 9 13 9 1 9 0 9 1 9 0 9 9 9 2
29 3 13 1 9 2 3 13 0 7 0 9 2 3 1 9 7 9 9 13 0 9 2 15 13 9 7 13 9 2
15 1 0 9 4 1 9 12 1 9 0 9 13 12 9 2
11 0 1 9 13 1 0 9 13 0 9 2
18 1 0 9 4 1 10 9 13 15 9 1 9 1 0 9 12 9 2
19 13 1 15 9 11 11 1 11 2 9 9 0 1 9 9 12 2 12 2
4 9 2 0 9
2 0 9
13 10 9 15 13 13 10 9 1 0 9 0 9 2
9 15 3 0 15 13 3 0 9 2
5 15 7 9 9 2
19 3 15 13 13 2 16 1 0 9 13 1 9 13 9 2 1 0 15 2
10 1 12 1 0 9 15 9 13 3 2
6 0 9 13 0 9 2
24 3 14 9 10 9 13 0 9 7 3 15 9 13 1 0 9 9 9 13 1 15 3 0 2
27 0 9 13 3 9 2 15 3 3 3 13 2 7 14 0 1 0 13 0 13 15 0 9 1 0 9 2
6 11 11 2 11 1 11
14 0 9 0 1 10 9 13 1 0 9 7 0 9 2
26 13 14 9 2 15 4 13 1 0 0 9 2 7 7 15 2 1 15 15 9 2 9 13 16 9 2
3 9 13 9
8 1 10 9 2 9 9 1 9
11 0 9 13 1 9 15 0 2 15 13 2
6 3 7 0 9 13 2
38 7 3 2 16 1 0 9 13 0 9 2 15 15 13 9 9 1 9 2 13 15 13 2 16 1 11 3 13 0 9 0 0 9 2 9 7 9 2
12 7 3 0 9 3 13 9 2 3 3 13 2
7 0 9 13 1 0 9 2
43 1 9 1 0 9 11 13 9 0 9 2 1 0 9 13 9 2 15 13 9 2 14 3 1 9 0 9 1 0 9 2 7 1 9 9 2 9 3 15 13 7 3 2
28 9 2 15 15 1 10 9 13 7 13 1 9 2 16 15 13 1 9 2 15 13 2 13 1 10 9 9 2
14 1 0 9 0 9 13 13 9 7 13 15 1 9 2
10 13 10 9 2 15 4 13 0 9 2
6 13 1 9 2 12 2
3 13 10 9
5 9 13 9 2 9
3 13 10 9
10 0 9 2 9 1 0 9 7 9 9
15 13 0 9 13 9 13 9 9 2 15 13 9 10 9 2
21 13 15 3 13 0 2 15 13 1 9 0 15 10 9 2 9 2 9 7 9 2
5 1 10 9 13 2
26 3 15 13 0 0 9 2 9 7 9 2 9 1 9 0 9 2 9 9 9 2 0 7 0 9 2
11 9 13 13 3 13 7 15 2 15 13 2
36 7 1 10 9 1 9 9 4 13 3 13 10 9 1 0 9 2 1 10 9 9 13 9 2 1 3 0 9 13 13 2 10 0 9 13 2
10 0 9 13 3 13 7 10 0 9 2
11 7 3 12 1 9 15 13 0 9 9 2
27 0 2 15 13 0 1 10 9 13 2 13 15 13 1 9 2 9 11 11 2 7 1 10 9 15 13 2
17 9 2 15 13 2 13 0 7 4 1 10 9 13 10 0 9 2
11 9 2 0 12 9 13 9 1 9 9 2
10 2 1 9 7 12 9 13 1 11 2
5 13 10 0 9 2
12 2 13 4 0 9 11 2 9 9 7 9 2
21 1 9 12 4 3 13 9 0 9 9 2 0 1 0 9 2 9 7 0 9 2
5 13 15 0 9 2
10 13 9 1 9 9 2 9 7 9 2
24 13 4 3 9 1 9 0 0 0 9 1 12 9 2 0 1 9 9 7 9 9 3 9 2
8 13 4 3 9 1 9 9 2
22 2 3 13 9 7 9 9 7 9 2 13 0 9 9 2 15 13 0 3 15 13 2
13 13 10 9 1 9 1 9 7 9 1 9 9 2
10 9 1 0 9 13 3 1 0 9 2
14 13 4 9 9 1 0 9 1 9 9 0 0 9 2
13 1 9 13 0 13 1 9 11 7 10 0 9 2
15 13 9 0 3 13 2 13 15 7 1 0 9 7 9 2
23 2 9 13 13 3 2 16 1 0 4 13 9 2 13 15 3 3 13 7 13 0 9 2
9 2 13 9 13 1 0 0 9 2
5 13 0 0 9 2
8 3 13 9 1 9 0 9 2
6 0 13 1 0 9 2
9 3 13 0 7 0 13 1 9 2
20 2 13 3 0 9 2 16 4 13 3 0 2 1 15 13 7 1 15 14 2
9 3 1 15 7 3 0 0 9 2
7 9 9 13 1 15 0 2
14 13 7 0 9 10 0 9 2 16 0 1 0 9 2
15 0 15 3 13 2 7 0 3 1 9 9 10 9 13 2
25 2 1 0 9 13 0 0 9 2 1 15 15 4 3 13 2 7 3 13 13 15 2 15 13 2
25 2 0 9 13 1 15 13 1 15 9 9 2 13 0 9 0 9 2 9 15 0 7 0 9 2
10 2 13 0 9 12 2 12 12 9 2
2 0 9
11 13 9 1 9 9 2 7 9 7 9 2
10 2 13 1 11 2 13 10 0 9 2
10 2 13 4 0 9 9 0 1 11 2
18 1 9 12 2 12 4 13 9 9 7 9 1 11 11 1 0 11 2
48 12 9 4 13 1 9 9 2 3 3 1 9 9 9 2 9 9 4 13 0 1 12 9 1 11 2 12 9 9 7 9 1 0 9 1 11 2 1 9 1 11 16 0 0 9 0 9 2
11 1 0 0 9 4 13 12 7 12 9 2
18 2 3 9 7 9 13 9 2 9 7 9 2 0 9 13 1 9 2
12 1 9 1 0 9 4 13 9 11 7 11 2
4 0 9 13 2
11 13 0 13 3 1 9 2 3 1 9 2
14 13 1 9 1 11 3 0 13 2 7 13 9 14 2
34 2 13 15 13 9 2 15 4 15 3 3 13 2 13 14 9 2 7 3 9 2 16 15 2 15 13 2 1 15 13 2 13 9 2
7 2 0 0 9 15 13 2
24 13 3 3 7 1 0 9 13 1 9 2 7 15 3 3 9 2 3 1 9 2 0 9 2
6 13 3 0 0 9 2
6 13 15 9 0 9 2
12 13 15 3 0 2 0 9 2 16 0 9 2
19 9 9 2 1 15 13 13 2 13 0 2 7 9 4 13 0 7 0 2
28 2 13 9 1 9 10 0 9 2 7 15 16 0 9 2 7 16 0 0 9 1 9 9 7 9 2 9 2
11 2 13 2 16 0 9 13 9 1 9 2
14 2 10 9 7 9 13 9 12 2 12 12 9 3 2
41 9 2 11 2 0 2 9 2 2 1 9 12 2 12 12 11 12 2 9 2 2 2 12 2 12 12 2 9 12 2 9 2 5 9 2 2 12 2 12 12 2
4 9 1 9 2
13 9 9 2 1 9 15 9 13 13 10 0 9 2
1 9
14 9 0 7 0 9 13 1 0 9 3 14 3 0 2
6 3 7 13 9 9 2
12 13 0 13 9 0 9 7 3 13 0 9 2
18 3 15 13 2 16 9 13 1 0 9 2 7 0 9 13 3 0 2
17 0 9 2 3 13 11 13 2 13 0 9 2 7 9 0 9 2
19 0 9 0 7 0 9 13 13 3 0 2 15 15 13 3 9 7 9 2
9 11 11 2 9 0 9 11 2 11
3 0 9 9
6 0 9 9 1 0 9
59 16 0 9 1 9 9 9 11 11 11 1 9 1 9 0 9 13 2 16 9 9 9 1 0 9 4 2 13 2 1 9 2 13 3 3 2 16 9 7 3 9 11 15 1 0 9 13 13 1 0 9 9 0 7 3 0 9 9 2
28 13 0 9 2 16 0 0 9 2 16 3 14 1 9 9 2 15 13 1 9 9 1 0 2 0 2 9 2
36 10 9 13 0 2 3 7 9 9 2 16 7 0 0 9 13 13 15 2 16 4 0 9 4 13 1 9 2 15 13 1 10 9 15 0 2
2 9 9
20 1 9 1 10 9 9 13 2 16 3 9 9 1 0 9 0 9 9 13 2
35 13 15 3 1 9 0 0 9 2 1 15 9 13 15 0 16 9 1 0 7 0 9 0 7 3 0 9 7 0 9 1 9 0 9 2
21 0 9 9 13 3 13 15 2 16 1 0 9 13 9 10 9 3 9 12 12 2
28 1 15 13 3 13 3 16 12 0 9 2 15 4 1 9 0 9 3 13 16 0 9 9 1 3 0 9 2
34 7 1 10 9 7 13 10 9 2 16 9 0 1 0 9 4 1 9 9 1 12 7 12 9 13 1 9 0 9 7 1 0 9 2
24 3 9 2 3 3 12 2 12 9 9 13 13 16 0 7 0 9 15 2 15 15 3 13 2
4 9 2 9 2
32 9 1 0 9 13 3 0 7 3 2 16 4 3 4 13 0 9 2 1 15 15 13 1 9 15 0 0 0 7 0 9 2
55 0 0 9 9 9 9 3 13 10 0 9 1 9 2 15 4 13 13 0 9 9 2 16 4 13 3 13 9 2 10 0 9 13 0 9 2 7 9 0 3 0 2 0 7 15 0 3 0 7 9 7 9 0 9 2
2 11 11
4 11 13 3 0
9 14 1 12 2 9 1 9 1 11
6 2 0 0 9 13 9
15 11 13 3 0 9 14 1 0 2 7 7 0 9 9 2
26 1 10 9 13 9 9 1 0 9 7 9 2 11 2 1 9 1 0 9 7 9 9 10 0 9 2
23 1 9 9 0 11 13 13 1 9 2 0 9 7 9 1 9 14 11 1 0 0 9 2
13 1 9 0 9 15 16 0 9 0 0 11 13 2
40 0 9 0 0 9 15 13 3 2 16 13 9 9 0 9 12 0 9 11 1 0 0 9 1 9 2 16 4 13 9 1 9 1 0 9 9 1 0 9 2
4 14 1 0 9
14 1 9 9 9 11 1 0 9 13 3 0 9 0 2
23 10 0 0 9 1 9 13 3 1 12 5 9 0 11 7 1 12 5 9 0 0 9 2
24 1 0 9 13 11 1 11 2 15 1 0 9 13 0 9 2 7 3 13 1 11 7 11 2
13 0 11 15 13 3 1 11 14 1 12 2 9 2
18 13 15 12 5 1 11 2 7 3 1 11 2 11 2 11 7 11 2
18 11 4 3 13 7 11 2 16 3 13 1 11 2 0 11 7 11 2
37 1 11 13 13 14 0 9 2 16 11 2 15 15 1 9 3 1 11 13 1 0 9 1 11 2 13 1 9 0 0 9 14 1 12 2 9 2
2 3 0
24 16 11 3 13 1 0 9 11 2 13 15 15 3 3 0 9 2 13 12 1 0 9 9 2
37 1 9 9 1 12 3 0 9 9 13 1 9 1 11 0 3 11 2 1 12 5 2 2 11 2 1 12 5 2 7 11 2 1 12 5 2 2
9 1 0 12 9 11 15 13 3 2
44 9 9 7 9 13 3 1 9 0 1 0 11 2 1 12 5 2 2 1 0 9 0 2 1 12 5 2 2 1 11 2 1 12 5 2 7 1 11 2 1 12 5 2 2
13 1 15 15 3 13 0 9 0 9 1 0 9 2
15 1 9 0 11 13 0 9 7 0 9 0 9 1 9 2
33 9 7 13 13 3 0 2 16 1 15 9 15 9 1 0 9 11 13 3 7 1 10 9 4 15 13 13 1 9 0 0 9 2
3 1 9 13
19 9 0 0 9 13 1 0 0 9 1 9 12 12 5 7 3 12 5 2
17 3 13 1 9 0 11 10 0 9 3 3 1 0 0 9 3 2
18 13 10 9 1 0 11 1 12 5 7 1 0 0 9 1 12 5 2
41 0 0 9 7 13 2 16 9 0 11 1 0 0 9 3 13 7 1 0 9 0 9 15 13 1 12 5 1 12 9 9 2 1 12 5 1 0 9 9 12 2
27 0 9 0 9 1 0 0 9 13 3 1 0 9 9 2 3 9 13 1 0 9 0 9 1 12 5 2
8 9 1 9 13 1 12 5 2
23 0 13 2 16 0 9 1 0 9 11 13 3 1 9 1 0 9 0 3 1 12 5 2
28 3 1 0 9 0 9 13 1 9 7 9 1 9 12 9 2 15 13 12 5 9 0 9 1 0 0 9 2
4 9 1 12 9
22 13 15 2 16 9 1 0 0 9 13 3 7 1 0 9 1 12 7 12 5 3 2
12 7 3 15 4 3 13 0 9 9 7 9 2
22 15 13 15 2 16 0 9 3 13 7 0 9 2 15 13 3 0 1 9 0 9 2
20 9 13 2 16 0 0 9 15 1 0 9 13 0 0 9 3 1 9 12 2
2 11 0
14 9 9 1 9 1 9 12 2 0 11 5 12 5 2
8 9 1 9 2 9 1 9 2
10 3 1 0 9 13 3 0 7 0 2
9 13 15 7 1 0 0 9 11 2
1 11
3 1 0 9
16 9 11 1 9 7 9 0 9 7 0 9 1 9 0 9 2
6 9 13 1 0 9 2
15 9 7 0 9 9 13 0 2 16 9 9 13 1 9 2
30 9 2 11 2 0 12 2 12 12 11 2 9 2 2 2 12 2 12 12 2 12 2 9 2 2 12 2 12 12 2
1 11
3 1 0 9
15 9 0 11 1 9 7 9 0 9 0 9 2 3 0 2
21 1 12 9 9 9 13 12 5 9 9 1 9 7 9 9 3 3 13 0 9 2
12 9 13 3 13 9 9 7 3 15 15 13 2
35 9 2 0 11 2 9 2 9 2 0 2 2 0 12 2 12 12 11 2 9 2 2 2 12 2 12 12 2 9 2 2 12 2 12 12
1 11
3 1 0 9
15 11 1 9 9 0 9 2 15 4 13 1 0 0 9 2
3 9 9 11
40 16 15 13 1 0 9 2 9 2 1 9 7 9 2 3 15 13 2 16 3 13 4 3 13 13 0 9 2 0 15 9 9 2 9 7 3 9 10 9 2
50 16 15 15 3 13 2 16 9 2 9 7 3 9 1 9 13 9 7 9 7 3 13 2 16 9 13 0 14 1 9 2 15 13 9 0 0 9 2 15 15 13 1 9 2 13 14 1 9 11 2
10 3 1 9 10 9 13 9 1 9 2
13 0 9 7 9 13 13 7 1 9 1 0 9 2
15 7 3 2 13 13 9 1 9 7 9 1 9 1 15 2
17 15 13 13 2 16 13 15 0 2 7 7 10 9 13 0 13 2
13 7 9 9 3 13 15 1 9 7 9 1 9 2
33 3 13 0 13 2 16 9 13 9 13 1 0 2 16 4 15 1 9 13 1 9 9 7 9 9 9 2 7 13 15 0 9 2
31 3 4 3 13 13 1 9 2 16 0 9 2 7 1 0 3 9 13 2 13 13 1 9 0 0 9 7 0 0 9 2
13 7 3 13 1 15 2 16 13 1 9 7 9 2
48 9 2 9 7 9 2 0 7 0 9 2 4 15 13 13 1 9 2 16 13 13 9 9 1 12 9 0 0 9 7 9 1 9 9 9 1 9 2 16 4 13 1 9 1 9 12 9 2
23 3 3 13 0 13 9 2 16 4 4 13 9 0 9 2 7 1 9 1 12 9 9 2
33 3 13 2 13 0 13 3 0 9 2 0 7 0 9 2 16 9 13 9 13 0 2 16 4 15 2 13 2 0 9 1 9 2
9 3 3 13 13 0 7 0 9 2
10 0 9 13 13 9 9 0 7 0 2
16 3 7 13 10 10 9 7 9 2 3 15 15 4 13 9 2
2 11 11
24 13 0 7 3 0 9 2 0 12 2 11 12 2 9 2 5 9 2 2 12 2 12 12 2
4 9 14 1 9
8 1 9 9 13 0 9 9 9
33 9 2 9 2 9 2 9 2 9 0 7 1 12 0 9 1 0 11 2 11 7 3 13 9 9 7 9 2 15 13 9 11 2
18 9 15 13 16 0 9 1 9 1 0 7 0 9 2 1 10 9 2
2 11 11
15 9 9 11 7 11 0 13 9 1 0 0 9 1 9 2
9 0 9 9 4 7 10 9 13 2
7 13 15 3 1 0 9 2
2 13 9
9 9 9 13 14 9 15 9 9 2
13 1 9 9 13 0 13 3 0 2 3 0 9 2
16 13 14 1 12 0 16 0 9 2 7 13 9 3 10 9 2
15 3 15 3 13 2 3 13 9 3 0 2 10 13 9 2
22 9 9 1 0 9 3 13 3 12 5 2 16 9 1 0 9 13 3 12 5 9 2
2 13 9
13 1 9 9 3 13 9 0 9 1 9 1 9 2
5 3 13 0 9 2
6 11 15 13 10 9 2
8 7 15 13 1 0 9 9 2
33 3 13 0 0 9 2 15 0 7 0 9 13 3 1 9 0 9 2 7 13 15 1 9 2 9 9 2 3 0 9 0 9 2
32 3 13 0 13 15 2 1 9 15 3 3 13 3 0 9 1 0 9 9 1 9 2 7 13 9 3 9 9 1 0 9 2
29 15 9 9 11 7 13 1 0 0 9 7 13 1 15 14 0 9 9 2 9 7 9 2 7 3 7 0 9 2
10 1 0 9 15 13 9 0 9 9 2
9 7 3 15 2 3 10 9 13 2
9 1 9 9 13 3 12 9 9 2
11 1 10 9 13 1 9 7 1 0 9 2
7 3 13 0 9 1 9 2
6 15 7 1 9 13 2
11 0 0 9 13 3 7 3 13 9 9 2
9 0 9 13 1 9 1 10 9 2
10 13 0 0 9 2 9 0 9 9 2
9 3 9 0 9 13 9 9 9 2
11 0 9 13 2 16 1 15 13 9 9 2
12 3 13 13 1 9 1 0 0 9 7 9 2
3 9 13 0
10 1 11 13 1 0 9 12 0 9 2
7 13 1 15 13 0 9 2
16 0 9 3 13 9 7 9 2 1 0 9 13 13 1 9 2
5 9 13 0 9 2
15 1 0 9 1 15 13 2 16 4 15 13 13 10 9 2
13 13 4 1 0 9 14 12 5 2 13 11 11 2
10 1 9 4 13 3 11 2 3 9 2
33 15 15 13 0 3 1 9 1 9 9 2 1 0 9 2 1 9 1 9 9 2 7 10 9 15 13 7 1 9 9 1 11 2
24 16 9 9 4 15 13 3 13 0 9 2 0 1 0 9 2 16 1 15 4 15 13 9 2
12 15 4 13 1 9 1 0 9 9 1 0 2
19 0 9 4 13 7 1 9 9 2 16 3 9 13 9 1 9 0 9 2
2 0 9
18 10 9 9 13 1 9 9 16 9 9 2 15 3 13 0 9 9 2
11 9 1 9 1 9 7 9 10 9 13 2
19 13 7 9 1 9 7 0 9 7 9 9 2 1 9 2 1 10 9 2
12 9 1 15 13 11 3 13 1 9 0 9 2
44 9 2 11 2 9 2 9 2 0 2 2 1 9 12 2 12 2 12 12 11 12 2 9 2 2 2 12 2 12 12 12 2 12 12 12 2 9 2 2 12 2 12 12 12
2 9 2
11 9 9 7 9 2 9 13 7 0 9 2
1 9
5 0 9 13 9 9
4 9 7 0 9
6 0 9 7 10 9 2
4 14 7 1 9
16 1 0 9 0 9 15 0 9 13 0 9 0 9 7 9 2
7 4 7 13 9 7 9 2
22 13 10 0 9 2 14 13 7 13 2 1 10 9 2 13 9 9 2 12 2 12 2
10 13 7 0 13 10 9 7 0 9 2
23 0 9 13 0 9 1 15 2 16 9 0 9 7 9 1 11 13 1 9 11 1 11 2
3 9 1 11
10 16 3 0 0 9 13 9 11 11 2
21 15 15 1 9 12 13 1 9 1 9 2 16 4 15 3 1 11 13 0 9 2
12 16 15 13 1 9 2 0 0 9 3 13 2
25 13 1 10 9 0 0 9 1 9 2 1 10 9 11 1 9 12 13 11 1 9 1 11 12 2
28 12 1 9 9 13 2 16 11 3 1 9 0 9 13 15 2 16 4 15 0 13 9 2 9 7 9 15 2
11 14 1 9 13 0 0 9 1 10 9 2
24 0 0 9 13 11 11 2 15 15 13 13 9 9 2 15 13 10 9 1 11 7 1 11 2
20 9 9 12 15 13 13 0 0 9 7 3 13 9 1 0 9 7 0 9 2
24 1 9 9 13 11 2 15 0 9 9 0 9 13 1 9 1 0 2 0 9 1 9 12 2
11 0 9 0 9 13 10 9 1 9 3 2
2 10 9
12 0 9 13 13 16 9 2 7 16 0 9 2
27 13 2 16 1 0 0 9 0 9 13 1 9 0 9 9 0 9 0 1 9 12 1 0 9 0 9 2
11 13 1 9 12 0 9 2 9 0 9 2
32 1 9 1 9 15 13 15 2 15 0 9 3 13 2 13 2 1 15 7 1 0 13 0 9 2 15 13 13 13 1 9 2
10 16 13 2 16 0 15 1 9 13 2
63 9 2 15 2 16 15 4 9 13 7 15 3 13 0 2 3 1 0 9 2 9 2 9 2 9 2 9 2 9 2 9 2 1 9 15 0 9 1 9 2 7 1 9 0 9 1 15 2 3 1 9 9 9 2 1 15 4 9 7 0 9 13 2
10 9 2 0 7 0 9 0 15 9 2
34 9 0 15 2 3 7 3 2 9 0 9 13 13 9 9 2 9 2 9 2 3 15 0 2 15 4 9 9 13 7 15 13 0 2
18 3 7 15 2 15 1 9 9 1 9 0 1 0 9 13 1 9 2
17 9 9 10 9 13 1 15 2 16 0 4 13 9 13 0 9 2
2 9 9
6 9 9 9 13 0 2
15 13 13 0 2 0 2 13 7 0 9 7 9 1 9 2
17 9 13 7 1 10 9 2 16 13 9 13 9 2 9 7 9 2
26 9 9 13 4 13 14 1 9 9 0 7 0 9 2 1 10 9 15 0 1 0 7 0 9 13 2
11 15 4 0 9 9 0 9 4 3 13 2
16 9 4 13 13 3 3 2 16 13 0 9 9 1 9 9 2
20 10 0 9 13 3 15 2 16 15 0 9 13 3 0 3 2 16 9 9 2
12 0 9 13 2 16 9 13 13 13 1 9 2
13 9 2 13 2 13 2 16 13 0 9 10 9 2
12 9 7 13 13 3 0 1 9 1 9 0 2
5 11 11 2 0 9
4 9 1 9 2
8 13 9 2 9 3 3 13 2
10 9 1 9 2 7 3 6 1 15 2
20 1 10 9 13 1 0 9 0 9 9 1 0 9 9 1 9 9 7 9 2
34 1 0 9 12 7 12 15 3 1 0 13 7 15 2 15 13 0 2 3 3 0 2 9 1 9 0 0 9 1 0 9 0 9 2
8 1 9 15 13 2 7 15 2
21 3 13 0 2 16 4 1 0 9 13 1 9 1 9 2 7 15 13 9 9 2
13 15 7 13 3 3 2 15 13 9 10 0 9 2
4 13 15 13 2
8 13 13 0 9 9 9 12 2
6 13 15 9 7 9 2
24 9 1 15 13 2 15 9 4 15 13 3 13 2 7 15 3 9 2 3 7 10 0 9 2
21 13 3 14 13 0 9 10 9 1 10 0 9 2 3 15 13 9 12 7 12 2
4 9 13 9 2
6 9 13 1 0 9 2
18 13 3 9 0 7 0 9 2 15 13 9 2 16 1 15 15 13 2
12 7 15 2 1 15 13 0 1 0 9 13 2
5 13 1 9 12 2
5 9 2 9 7 15
3 9 1 9
13 13 0 13 0 0 9 1 9 1 0 9 9 2
5 15 13 0 13 2
6 11 2 11 2 2 11
17 9 13 3 9 9 2 12 2 12 9 2 2 2 0 9 2 2
26 1 12 9 2 12 0 9 15 9 13 0 9 0 3 9 0 9 7 1 0 9 1 9 9 9 2
22 0 9 15 3 13 14 9 0 2 7 10 9 13 4 13 7 3 2 3 9 9 2
27 1 12 9 2 12 0 9 13 0 9 2 3 7 0 2 0 2 9 2 2 0 9 0 1 9 9 2
13 0 9 1 9 12 3 13 9 7 9 0 9 2
65 1 9 12 10 0 9 13 9 1 9 0 9 7 9 2 15 13 0 9 13 1 9 9 7 10 9 1 0 2 16 1 0 12 9 15 13 0 9 7 4 13 9 9 2 15 13 0 9 1 3 16 12 9 7 9 1 9 0 16 12 9 13 10 9 2
36 16 15 1 0 9 9 0 0 9 1 0 9 3 13 1 9 9 1 0 0 9 2 4 13 1 9 3 9 9 9 1 3 16 0 9 2
40 3 13 1 9 9 1 9 9 9 13 7 0 9 2 3 0 9 2 9 0 9 7 0 9 2 3 3 9 2 15 13 0 9 2 3 9 7 9 9 2
27 1 10 9 13 1 12 9 2 12 9 2 9 2 0 0 9 0 0 9 2 1 10 9 13 9 9 2
29 3 0 9 15 4 13 9 2 3 9 4 13 15 1 9 2 15 13 13 1 0 9 16 9 9 7 9 9 2
29 13 4 13 2 16 1 12 9 2 12 13 9 1 9 1 9 9 13 9 1 9 9 2 1 15 4 9 13 2
19 1 10 9 7 13 0 9 7 13 1 9 9 2 16 15 13 7 3 2
35 9 13 0 13 2 16 1 0 2 9 0 2 0 2 9 2 1 9 15 9 13 3 0 9 9 0 9 1 9 7 0 9 10 9 2
3 9 7 9
13 0 9 13 1 9 0 9 9 1 12 0 9 2
13 0 9 15 3 13 7 1 10 9 0 9 13 2
9 15 13 3 0 2 13 12 9 2
10 10 9 13 1 9 1 9 9 0 2
20 13 4 15 2 16 15 9 13 13 16 9 0 1 9 2 16 1 15 13 2
7 11 2 11 2 2 0 11
24 0 9 2 15 13 1 9 10 0 9 1 9 1 9 1 9 2 13 1 9 1 9 13 2
38 9 1 9 1 9 4 1 12 9 9 2 12 2 12 9 2 13 3 2 16 13 3 13 0 9 9 2 3 9 9 2 2 1 15 15 9 13 2
32 9 0 1 9 9 0 9 1 9 1 9 13 1 9 1 9 13 2 15 13 2 16 9 9 1 10 9 9 1 9 13 2
3 9 1 9
23 13 0 13 9 9 1 9 2 16 0 9 13 13 0 9 2 0 9 7 9 1 9 2
19 3 4 9 2 9 2 15 3 1 10 9 13 2 7 9 1 9 13 2
6 11 2 11 2 2 11
29 1 9 2 10 9 13 1 9 0 9 0 9 3 13 2 1 9 2 0 0 9 3 2 2 15 0 9 13 2
10 0 9 10 9 13 12 9 0 9 2
32 16 13 7 9 7 9 1 9 9 0 9 7 13 7 1 0 9 9 9 2 13 1 9 9 1 9 1 9 9 10 9 2
2 11 11
28 13 0 9 11 2 0 2 0 12 9 2 12 12 11 12 2 11 2 9 2 2 2 12 2 12 12 12 2
3 9 9 2
5 1 9 7 1 11
13 3 15 0 9 3 3 13 1 0 9 7 0 9
13 13 9 16 9 2 14 0 7 3 1 0 9 2
32 13 4 15 1 15 3 2 16 15 10 0 9 13 1 9 0 9 2 16 12 13 13 3 0 9 7 0 0 2 3 0 2
8 10 9 13 3 3 3 13 2
2 11 11
46 9 13 3 3 13 2 16 1 15 16 4 13 1 10 9 2 3 9 1 15 13 0 9 7 9 0 9 2 0 9 7 9 0 9 2 13 0 2 6 2 7 13 13 0 9 2
5 13 15 10 0 9
32 9 9 1 9 2 3 1 10 0 9 13 3 3 3 0 2 16 1 9 9 0 9 15 1 9 13 16 1 10 0 9 2
27 9 9 1 11 12 11 11 2 9 14 16 13 15 0 9 3 2 7 0 1 15 15 1 9 7 13 2
12 10 9 15 3 3 13 1 12 7 0 9 2
32 16 4 13 9 13 15 2 3 3 3 1 15 2 13 2 9 1 9 11 2 9 7 10 9 13 15 10 0 9 2 2 2
22 12 9 1 0 9 15 1 9 0 9 1 0 9 11 2 9 1 9 3 13 9 2
34 3 0 13 7 0 9 2 9 1 9 2 15 15 1 9 0 9 3 13 2 3 16 1 9 2 7 1 0 11 2 9 0 9 2
3 9 7 9
30 1 0 9 15 3 13 13 2 16 9 10 0 9 2 13 2 9 9 1 9 9 2 7 1 9 2 15 15 13 2
15 1 9 0 3 3 13 2 16 9 13 15 2 10 13 2
49 9 2 3 1 0 9 1 0 9 2 3 3 7 1 10 0 9 13 0 9 1 0 9 2 15 13 3 15 2 7 1 9 2 0 9 1 9 2 7 1 9 2 15 0 13 3 0 9 2
2 9 9
10 13 15 3 9 2 7 2 2 2 2
9 1 9 13 9 1 0 9 9 2
39 13 10 9 2 13 0 0 9 1 15 3 3 16 15 2 9 2 15 13 1 0 9 2 15 13 1 10 9 1 9 0 9 2 3 0 2 14 0 2
40 16 3 0 9 13 2 13 9 9 9 0 9 0 0 9 7 1 15 0 9 1 9 15 2 3 2 3 7 3 15 13 13 3 10 0 2 0 9 2 2
8 13 1 9 2 12 2 12 2
3 9 1 0
3 12 0 9
4 9 1 9 2
22 9 9 2 9 15 9 13 2 16 9 2 13 9 1 9 3 3 9 2 13 9 2
2 0 2
3 11 15 13
12 0 9 13 14 9 2 7 7 9 1 0 9
15 0 0 9 13 2 16 9 0 9 15 1 9 9 13 2
23 15 1 15 13 2 16 1 9 15 9 13 2 13 1 0 9 2 7 3 15 7 13 2
20 13 15 1 9 1 10 0 9 3 1 10 0 9 2 3 15 9 13 3 2
2 11 11
26 1 15 2 16 4 15 13 9 0 9 2 3 0 9 3 9 13 2 2 13 0 13 3 12 9 2
39 3 13 0 9 0 0 9 2 15 13 0 15 1 0 9 2 1 9 0 9 2 13 1 10 9 3 2 16 13 9 0 9 7 13 15 1 10 9 2
43 1 0 13 1 0 9 10 0 9 2 3 15 13 0 0 9 2 14 1 9 2 13 1 15 2 16 0 2 7 1 12 9 2 2 7 1 0 13 15 9 1 9 2
4 9 15 13 12
57 16 13 9 1 0 9 10 9 1 9 3 1 15 2 14 13 2 16 1 9 9 3 13 2 16 3 13 1 9 0 9 12 0 9 2 3 16 15 0 9 3 13 2 2 13 15 13 2 3 15 13 1 0 9 1 9 2
17 13 3 2 16 10 9 13 3 12 2 1 3 0 9 4 13 2
27 13 15 7 12 10 9 2 16 0 2 7 3 3 0 2 9 15 13 0 9 2 3 1 9 0 9 2
2 0 9
31 13 9 2 3 15 9 0 9 13 0 9 2 7 15 3 1 9 1 9 13 2 7 7 15 13 1 9 9 7 9 2
34 0 9 0 9 2 7 0 1 9 2 1 0 9 2 1 0 2 1 0 9 1 12 2 12 9 13 13 3 1 12 7 12 9 2
27 9 1 0 9 11 2 1 15 3 0 2 3 16 0 0 0 9 0 9 13 1 12 5 7 3 0 2
16 3 13 9 2 10 9 15 13 0 9 3 2 16 9 9 2
27 10 0 11 2 11 11 12 7 11 12 2 2 15 3 13 0 0 0 9 2 13 1 12 1 12 9 2
39 0 9 9 1 9 9 1 9 2 3 1 0 9 0 9 2 0 9 9 2 13 0 9 13 9 0 9 2 7 13 15 2 16 0 0 9 13 9 2
32 0 7 0 9 2 3 1 0 9 9 1 0 9 2 3 16 9 1 0 9 9 2 13 3 3 1 9 0 2 16 0 2
3 13 15 12
16 0 9 13 13 1 12 9 2 7 3 13 0 9 13 12 2
107 1 15 13 9 1 0 2 9 0 0 9 2 9 2 12 7 12 9 2 2 9 2 12 7 12 9 2 2 9 2 0 9 1 12 7 12 9 2 0 0 7 9 2 2 9 2 3 1 12 9 2 9 0 9 14 1 9 2 0 14 1 12 9 2 2 9 2 6 12 9 2 9 14 12 9 2 7 9 9 2 16 13 9 2 9 2 9 2 9 9 2 9 1 9 9 2 15 15 13 15 1 0 12 7 12 9 2
38 9 2 15 13 9 2 16 0 9 13 3 1 15 2 1 10 0 9 1 9 0 9 2 13 9 2 16 0 2 7 0 2 9 13 3 3 3 2
20 3 13 7 0 9 1 9 2 9 7 9 13 2 12 2 7 3 3 12 2
5 15 0 15 13 2
14 0 2 7 3 3 0 2 13 9 1 9 7 9 2
50 13 3 9 2 9 0 3 1 12 9 2 0 13 1 12 2 16 15 7 3 13 2 2 0 1 9 1 9 12 2 12 2 7 3 0 9 2 9 1 12 7 12 9 2 2 7 9 7 9 2
30 3 13 9 14 13 1 9 2 16 1 9 13 15 16 1 9 2 15 13 2 15 13 2 7 15 13 2 15 13 2
59 9 2 16 13 1 9 0 9 2 9 2 9 14 1 12 9 2 13 3 2 3 9 1 12 9 2 0 7 0 1 9 13 0 9 2 2 7 9 0 9 2 12 9 1 9 2 16 15 13 13 15 1 9 1 9 1 9 2 2
2 9 9
76 9 2 15 13 14 1 10 0 9 2 3 13 13 0 9 2 3 15 3 13 2 16 1 15 2 16 4 1 0 2 9 2 1 0 9 7 9 1 9 13 1 15 2 13 15 1 0 9 14 12 9 1 9 9 1 9 13 1 9 1 9 15 9 3 12 2 16 9 1 15 4 13 0 12 9 2
30 13 1 9 2 9 1 9 2 1 9 0 9 2 15 15 11 13 2 15 13 0 13 7 1 10 3 3 0 9 2
19 1 15 13 3 9 2 7 14 1 9 2 16 4 10 0 9 3 13 2
25 16 9 1 9 13 9 1 9 1 0 9 2 3 3 1 15 2 15 3 3 3 13 1 9 2
3 9 2 9
4 3 13 9 3
4 9 1 9 2
19 10 9 1 15 2 15 15 1 9 13 14 3 13 2 7 0 9 13 2
34 1 9 9 9 12 9 1 9 1 9 1 9 12 2 12 1 0 9 9 2 9 2 2 13 13 3 1 9 2 3 13 1 9 2
4 15 13 3 2
1 9
14 0 9 9 1 0 7 0 9 2 1 12 2 12 2
7 9 9 9 9 9 0 9
6 9 0 12 12 12 11
7 9 0 12 12 12 11 12
7 9 0 12 12 12 0 9
8 9 0 12 12 12 11 12 9
7 9 9 12 12 12 11 12
9 9 9 12 12 12 11 12 2 12
6 9 0 12 12 12 9
8 9 0 12 12 12 11 12 9
7 9 0 12 12 12 11 12
6 9 0 12 12 12 11
7 9 0 12 12 12 11 12
6 9 0 12 12 12 11
6 9 0 12 12 12 11
7 9 0 12 12 12 11 12
5 0 0 9 13 9
8 13 1 9 9 9 11 11 11
32 16 9 9 7 10 9 13 0 9 3 13 2 1 9 1 9 1 9 9 9 11 4 15 1 9 13 1 9 11 11 11 2
11 2 3 13 1 0 9 0 13 9 0 2
3 3 3 2
19 9 0 0 9 13 3 3 2 16 15 0 9 1 0 13 13 1 9 2
13 1 10 9 2 16 1 9 4 10 9 13 9 2
7 0 9 3 3 13 9 2
19 3 13 9 0 9 13 3 9 2 7 3 0 2 16 15 13 0 9 2
19 2 3 13 13 1 0 9 0 13 1 0 9 2 3 1 0 9 9 2
2 3 2
15 1 15 13 0 9 2 15 9 13 13 7 13 0 9 2
16 13 0 9 1 9 0 4 1 10 9 13 13 15 10 9 2
41 16 15 13 10 0 9 2 15 15 4 3 13 9 2 13 15 1 15 0 2 16 16 4 15 13 16 10 9 2 13 1 15 9 7 13 1 15 9 0 9 2
9 3 15 13 1 0 7 0 9 2
12 0 0 9 16 0 9 13 1 15 0 9 2
24 2 13 15 2 16 1 9 12 0 9 2 0 7 0 7 11 2 13 0 9 1 10 9 2
17 1 0 7 0 3 14 2 3 13 1 15 2 15 13 0 9 2
14 1 11 13 9 9 10 9 2 16 3 0 9 13 2
7 15 4 10 9 13 13 2
6 3 15 13 9 11 2
6 7 15 4 15 13 2
5 13 15 0 9 2
9 7 1 15 4 0 13 3 13 2
13 11 13 10 9 7 15 15 13 13 9 1 9 2
12 2 3 15 13 2 16 15 10 9 3 13 2
28 3 7 3 2 16 0 9 2 3 15 2 1 9 13 9 13 15 9 2 16 9 1 15 13 9 0 9 2
10 7 0 9 13 3 0 9 1 9 2
8 2 10 9 1 9 9 11 2
4 0 15 9 2
26 3 15 3 13 2 16 13 1 0 9 2 16 3 15 13 10 0 0 9 2 15 3 13 13 0 2
3 13 12 9
9 1 9 13 0 11 9 9 9 3
23 10 0 9 2 1 0 9 3 12 7 12 9 9 9 13 1 10 9 0 0 0 9 2
13 7 1 9 4 13 13 1 9 9 1 0 9 2
19 11 13 0 7 0 9 2 9 2 9 2 9 2 9 2 9 7 9 2
29 13 15 9 2 3 15 3 0 9 1 12 9 9 3 3 13 1 0 9 2 3 15 15 13 1 15 0 9 2
2 0 9
13 1 9 0 0 9 1 9 12 9 13 0 9 2
22 9 0 9 4 3 13 1 9 0 9 2 0 2 0 2 0 7 0 9 3 9 2
26 3 0 9 2 9 0 7 9 2 13 13 3 1 9 9 2 3 1 9 9 2 9 7 0 9 2
8 0 9 3 13 0 9 11 2
32 10 0 9 1 9 0 9 13 1 9 1 0 9 2 15 1 0 9 13 1 9 0 9 2 13 12 1 10 9 11 11 2
13 13 9 2 16 0 9 3 13 13 1 0 9 2
10 3 13 1 9 14 1 10 0 9 2
17 0 9 7 13 1 9 2 3 4 13 13 7 1 3 0 9 2
11 10 0 9 13 7 13 1 0 0 9 2
10 9 13 3 1 9 1 9 10 9 2
9 3 4 1 9 13 13 0 9 2
13 7 4 3 13 9 0 0 9 2 13 11 11 2
3 9 1 9
12 3 9 0 0 9 13 13 9 16 0 9 2
22 1 1 0 0 9 13 1 12 0 9 13 7 13 2 15 13 9 10 7 15 9 2
27 1 10 9 11 13 1 9 0 9 0 9 1 3 16 12 7 9 9 9 2 15 4 13 7 9 11 2
15 3 1 15 4 13 9 0 0 9 7 0 9 1 9 2
13 12 9 13 13 0 9 11 7 0 7 0 9 2
29 1 0 0 9 11 13 9 0 9 1 0 1 0 9 7 9 0 9 2 15 4 13 9 0 0 9 1 11 2
8 10 0 9 7 13 15 0 2
11 1 9 0 9 13 3 9 9 9 9 2
15 13 4 13 1 11 0 9 16 0 9 1 11 7 11 2
20 3 13 1 15 13 1 9 9 11 0 9 2 15 13 2 16 13 0 9 2
15 1 10 9 13 15 9 0 9 7 9 2 13 11 11 2
22 3 1 12 9 15 13 11 13 7 1 0 0 9 1 9 7 13 2 0 2 9 2
32 9 2 11 2 0 2 9 2 2 12 12 11 2 11 2 9 2 2 2 12 2 12 12 2 9 2 2 12 2 12 12 2
6 9 0 2 9 2 11
5 9 2 1 9 2
5 9 2 1 9 2
7 9 9 0 9 12 9 2
1 9
5 9 2 10 0 9
6 0 9 1 0 2 11
19 1 9 12 13 0 0 9 1 0 9 7 0 9 1 0 2 11 0 2
27 1 0 12 9 15 0 9 13 1 12 9 9 1 9 12 2 3 3 1 11 2 1 0 12 9 9 2
8 0 9 13 3 0 16 9 2
19 10 0 9 13 0 0 9 2 9 1 9 7 0 9 7 9 1 9 2
19 0 9 15 13 3 1 0 9 2 3 9 2 9 7 0 0 9 9 2
15 0 2 11 3 13 0 9 9 2 15 15 13 0 9 2
14 14 12 15 4 13 1 9 2 0 0 9 13 9 2
21 0 9 1 9 9 1 0 9 0 2 11 13 14 1 12 9 9 0 9 11 2
12 1 0 9 1 9 9 0 9 13 11 11 2
12 1 0 9 13 3 13 9 1 9 1 11 2
20 0 7 0 9 13 1 11 7 0 9 1 9 3 0 9 1 9 0 9 2
17 9 1 0 9 13 12 9 9 1 9 0 7 0 0 0 9 2
16 1 0 9 10 9 3 13 0 9 2 15 13 1 9 11 2
22 0 0 7 0 9 1 11 13 0 9 13 9 1 0 9 2 9 7 9 0 9 2
24 13 1 0 9 1 0 7 0 9 3 2 7 9 9 1 9 0 9 7 9 0 0 9 2
1 9
26 1 0 9 1 0 2 11 1 12 9 13 9 11 9 2 15 4 13 1 12 9 1 9 12 9 2
10 13 13 1 9 13 1 0 12 9 2
23 1 0 0 9 13 0 9 13 9 9 0 0 9 1 0 0 9 2 3 9 7 9 2
37 9 2 11 0 7 0 11 2 0 12 2 12 12 11 12 2 9 2 2 2 12 2 12 12 12 12 2 9 2 2 12 2 12 12 12 12 2
5 9 2 9 2 9
5 9 12 2 12 2
21 11 12 2 0 9 1 9 2 11 2 9 0 0 9 12 2 2 12 2 12 2
2 12 2
30 13 9 9 2 12 12 11 12 2 0 9 12 2 9 2 2 9 2 2 12 2 12 2 9 2 2 12 2 12 2
33 11 12 2 9 9 2 9 7 9 2 12 2 9 0 9 9 7 9 2 9 9 7 10 0 9 2 12 2 2 12 2 12 2
34 13 0 11 11 2 12 12 11 12 2 0 12 2 9 2 2 2 12 2 12 2 12 2 9 2 2 9 2 12 2 2 12 12 2
40 11 12 2 9 2 9 9 2 0 7 0 9 2 9 2 9 2 9 2 9 1 9 2 9 2 9 2 9 15 9 2 9 2 12 2 2 12 2 12 2
2 12 2
32 13 11 2 9 2 9 2 0 2 2 12 12 11 12 2 0 12 2 9 2 2 9 2 2 12 2 12 12 2 12 12 2
25 11 12 2 0 9 2 11 2 0 9 9 2 9 2 9 2 9 2 12 2 2 12 2 12 2
2 12 2
40 13 11 11 7 11 2 9 2 0 9 2 12 12 11 12 2 0 9 12 2 9 2 2 2 12 2 12 12 2 12 12 2 9 2 12 12 2 12 12 2
33 11 2 9 2 9 12 2 0 7 0 9 14 1 0 2 9 7 9 2 9 2 9 2 9 2 2 12 2 2 12 2 12 2
2 12 2
33 13 11 2 12 12 11 12 2 0 12 2 9 2 12 12 2 12 12 2 12 12 2 9 2 2 9 2 2 12 2 12 12 2
24 11 2 9 2 11 11 11 2 0 9 0 7 0 9 7 9 2 12 2 2 12 2 12 2
2 12 2
22 13 11 11 2 12 12 11 2 0 12 2 9 2 2 9 2 2 12 2 12 12 2
40 11 2 9 0 9 2 0 9 2 0 9 2 0 9 9 2 9 2 9 7 9 2 9 2 9 2 0 7 0 9 2 9 2 12 2 2 12 2 12 2
2 12 2
56 13 9 9 2 12 12 11 2 0 9 2 0 9 12 2 9 2 2 9 2 2 12 2 12 12 7 9 2 9 2 9 2 0 2 2 12 12 11 2 0 9 2 11 12 2 9 2 2 9 2 2 12 2 12 12 2
32 11 2 9 0 9 2 11 12 2 0 0 0 9 2 9 7 9 1 9 9 7 9 1 9 2 12 2 2 12 2 12 2
2 12 2
11 13 9 9 11 1 9 1 9 9 11 2
20 9 2 9 2 11 12 2 12 2 0 0 9 2 12 2 2 12 2 12 2
2 12 2
25 13 11 2 0 2 9 2 2 12 12 9 2 11 12 2 9 2 2 9 2 2 12 2 12 2
5 9 12 2 12 2
5 9 12 2 12 2
5 9 12 2 12 2
23 11 2 11 2 9 9 7 9 2 9 12 2 0 9 9 2 12 2 2 12 2 12 2
2 12 2
42 13 11 2 9 2 9 2 0 2 2 0 9 2 12 12 11 12 2 0 12 2 9 2 2 2 12 2 12 2 12 2 12 2 9 2 2 12 2 12 2 12 2
13 9 2 0 9 2 11 2 11 2 11 1 11 2
5 9 12 2 12 2
8 12 2 12 2 12 9 2 2
35 13 9 11 2 12 12 11 12 2 9 2 11 11 12 2 9 2 2 2 12 2 12 12 2 9 2 2 9 2 2 12 2 12 12 2
36 11 2 9 11 2 11 11 2 0 9 0 9 2 9 2 9 2 9 0 9 7 9 1 0 7 3 0 9 2 12 2 2 12 2 12 2
2 12 2
37 13 9 0 11 2 9 2 9 2 0 2 2 12 12 11 12 2 0 12 2 9 2 2 2 12 2 12 12 2 9 2 2 12 2 12 12 2
5 9 12 2 12 2
38 11 12 2 9 9 2 0 0 9 7 9 9 2 12 2 9 2 13 15 3 1 12 2 0 0 9 7 9 9 11 1 11 2 12 2 2 12 2
2 12 2
38 13 0 2 0 2 11 2 2 0 11 2 9 2 9 2 0 2 2 12 12 11 12 2 11 1 11 12 2 9 2 2 9 2 2 12 2 12 2
3 13 9 2
4 0 9 0 9
27 13 3 0 9 7 9 3 13 1 9 9 14 9 2 7 0 9 2 14 3 1 9 2 7 0 9 2
20 7 0 9 2 15 1 10 9 13 9 1 9 1 0 0 9 2 13 0 2
34 0 9 4 13 9 13 15 7 13 3 12 1 12 0 9 2 9 2 9 7 9 9 2 9 7 9 9 9 2 7 0 9 2 2
21 9 13 1 9 0 0 9 1 12 2 9 12 2 0 13 9 1 0 9 2 2
9 9 13 0 9 9 9 2 11 2
4 9 0 9 2
2 12 2
21 10 9 13 0 9 1 9 9 2 13 0 9 2 1 15 13 1 9 9 13 2
2 12 2
12 13 9 0 9 2 0 9 1 0 0 9 2
2 12 2
17 13 9 0 9 2 9 2 9 2 9 3 2 2 1 9 9 2
2 12 2
9 13 0 9 0 9 2 9 2 2
2 12 2
7 15 13 1 9 0 9 2
6 9 1 9 0 9 2
19 12 2 7 15 13 9 7 9 9 1 9 2 7 9 1 9 0 9 2
2 12 2
29 9 9 13 3 0 9 2 0 7 0 9 2 0 9 9 2 9 9 7 9 2 9 9 7 9 1 9 9 2
11 1 10 13 0 9 0 2 0 2 9 2
2 12 2
9 9 13 9 1 9 7 9 9 2
2 12 2
22 11 2 9 2 0 2 2 9 2 0 2 2 9 2 0 2 7 9 2 0 2 2
26 11 2 9 2 0 7 0 2 2 9 2 0 9 2 0 9 2 2 9 2 0 2 0 9 2 2
15 11 2 9 2 9 13 9 3 2 2 9 2 3 2 2
2 12 2
23 9 9 2 9 7 9 2 9 9 2 9 7 9 2 9 9 7 0 9 2 9 9 2
50 9 2 11 2 0 0 9 2 11 9 2 9 2 9 2 0 2 2 0 2 9 2 9 2 0 9 12 2 12 12 11 12 2 9 2 2 2 12 2 12 12 2 9 2 2 12 2 12 12 2
17 0 9 2 9 13 2 13 15 7 13 0 0 9 1 0 9 2
4 9 2 0 9
2 9 9
6 10 9 13 3 3 0
16 1 10 9 1 9 9 1 9 1 0 9 4 1 9 13 2
2 9 2
30 13 4 15 13 2 16 13 9 1 9 15 0 2 9 9 0 9 11 11 2 15 9 1 9 4 1 9 9 13 2
11 2 9 1 9 0 9 13 7 9 9 2
11 3 4 15 13 9 1 9 13 0 9 2
11 1 9 1 9 13 9 13 1 10 9 2
37 7 4 13 13 1 9 9 1 9 2 3 1 9 9 1 0 9 7 0 9 2 9 9 1 0 9 7 9 9 16 9 9 1 9 0 9 2
6 2 3 15 3 13 2
6 14 9 13 3 0 2
4 9 13 3 2
11 9 1 9 13 1 15 0 7 3 0 2
21 13 2 14 0 9 2 0 7 0 9 2 3 0 9 2 3 9 2 13 9 2
11 2 13 3 9 1 0 9 3 3 0 2
12 3 3 2 7 10 9 13 1 10 9 13 2
19 1 9 13 3 9 16 1 9 1 0 9 9 7 1 9 9 0 9 2
18 1 9 15 15 13 0 0 0 9 7 9 2 0 9 2 0 9 2
12 3 15 13 7 1 0 9 2 3 0 9 2
11 2 13 15 1 9 9 9 1 0 9 2
16 0 9 9 16 9 9 3 13 1 1 0 9 7 9 9 2
22 3 2 13 2 13 9 0 9 2 3 1 9 2 3 4 15 13 13 1 0 9 2
33 13 15 2 3 0 9 4 13 1 9 2 16 4 9 9 0 9 13 7 9 4 1 9 10 9 13 9 13 1 0 0 9 2
32 9 1 9 1 9 13 3 0 2 13 1 15 2 16 9 0 15 3 7 3 9 1 9 4 13 13 0 0 7 0 9 2
6 0 9 2 1 7 1
9 9 11 4 1 9 13 3 7 3
16 1 9 9 11 4 13 0 9 16 1 9 9 1 9 11 2
13 13 15 2 16 9 4 1 9 13 3 7 3 2
16 13 1 15 12 1 12 0 9 11 1 0 9 2 0 3 2
11 10 0 9 9 13 9 7 9 9 11 2
42 0 9 13 9 11 11 2 2 16 13 10 9 2 13 13 2 16 13 15 0 0 9 2 15 4 13 1 11 1 0 9 7 15 13 1 9 7 9 3 10 9 2
17 13 9 2 9 2 9 2 13 9 9 2 9 7 9 1 9 2
27 2 0 9 9 13 1 10 9 0 2 7 0 9 14 1 9 9 0 7 0 13 9 7 9 1 9 2
11 0 9 0 9 4 13 3 9 0 9 2
13 3 13 2 11 13 0 7 0 9 7 1 9 2
44 2 16 15 10 9 2 15 15 13 1 0 9 9 2 10 9 13 2 13 0 13 9 9 0 1 9 9 0 7 13 15 2 16 3 15 13 0 2 13 15 1 0 9 2
19 2 11 2 11 3 13 9 1 15 2 16 11 4 15 13 13 0 9 2
36 7 13 9 0 9 1 15 2 16 13 1 9 9 11 7 11 2 7 1 9 9 2 9 0 9 1 0 9 7 9 7 9 9 9 11 2
33 1 9 1 9 11 11 13 9 2 1 15 13 2 9 0 7 13 15 15 9 7 0 9 7 15 9 0 15 1 10 9 2 2
16 1 9 1 9 0 7 0 9 13 2 16 9 13 9 11 2
7 9 3 13 9 0 9 2
31 2 13 15 9 7 9 9 1 0 9 2 7 15 13 2 16 9 4 13 1 9 9 2 1 9 7 9 0 9 2 2
5 9 1 9 2 12
15 2 3 4 15 13 13 12 9 2 2 13 3 11 11 2
40 0 9 11 2 11 2 11 2 15 13 0 7 0 9 2 15 1 9 9 13 1 0 9 2 0 0 9 13 13 1 9 2 3 2 1 9 9 1 11 2
3 2 11 2
4 9 2 11 2
2 11 11
6 0 9 13 2 9 13
16 1 0 0 9 13 9 3 1 0 9 2 16 1 0 9 2
29 3 15 3 9 11 3 13 2 9 13 3 9 1 9 2 9 7 0 9 0 9 16 1 9 0 9 1 9 2
3 9 1 9
9 9 1 9 0 7 0 9 1 9
21 0 9 1 0 9 13 10 9 0 0 9 11 2 11 2 11 1 11 1 11 2
27 9 2 15 13 0 7 0 9 2 3 3 13 1 0 9 2 13 15 7 1 9 2 7 3 1 9 2
24 0 9 0 9 15 7 9 2 0 9 9 16 0 0 9 1 9 0 9 2 1 9 13 2
20 0 9 9 7 9 13 1 0 9 2 15 9 9 13 1 0 9 1 9 2
24 1 10 9 7 9 2 9 1 9 1 0 9 9 2 3 9 13 2 16 9 10 9 13 2
8 2 9 9 4 13 13 9 2
36 1 1 15 2 16 0 9 1 10 9 13 12 9 9 2 9 0 9 11 2 11 2 11 4 13 13 7 1 0 9 3 1 12 0 13 2
36 13 15 2 16 9 13 13 0 9 7 9 4 13 13 10 9 3 16 1 9 1 9 9 2 2 13 15 0 0 9 9 9 9 2 11 2
45 9 3 13 2 16 1 9 9 13 9 0 9 13 12 9 3 2 16 4 3 13 12 0 9 2 16 4 2 3 16 0 0 9 2 13 1 9 0 9 13 9 1 10 9 2
6 15 13 9 2 13 3
1 9
6 15 13 9 2 13 3
48 11 11 1 0 9 0 9 9 15 3 1 9 9 1 9 1 9 13 2 2 1 9 9 13 9 9 9 1 10 9 2 1 15 4 15 13 1 9 9 1 0 9 1 12 2 9 12 2
12 1 9 0 13 3 0 9 16 1 9 9 2
27 16 13 1 9 0 9 1 9 2 0 9 1 9 0 7 9 9 4 15 13 1 9 0 9 13 2 2
6 3 4 9 9 13 2
14 2 9 9 4 13 9 1 9 9 2 11 7 9 2
19 1 0 9 13 1 1 9 9 9 0 2 16 15 13 9 7 9 9 2
22 9 7 13 11 13 0 9 2 15 13 13 1 0 9 2 16 4 9 9 13 2 2
13 11 4 13 2 16 4 13 9 1 0 0 9 2
7 15 13 7 9 0 9 2
22 2 10 9 2 15 13 3 1 9 2 13 0 9 7 13 15 13 0 9 16 11 2
25 7 15 2 15 13 0 9 11 2 4 1 15 3 1 0 9 13 9 1 9 0 1 0 9 2
22 9 13 13 3 2 3 9 13 0 9 3 3 2 16 15 13 1 9 13 9 2 2
6 0 0 9 2 2 2
1 9
6 0 0 9 2 2 2
39 1 9 9 15 0 9 9 11 11 13 15 2 3 13 1 9 9 2 3 1 0 9 13 1 9 9 1 9 2 3 13 0 9 2 16 15 13 9 2
26 0 9 9 11 11 3 13 1 10 9 2 0 9 9 3 4 13 2 7 3 15 1 15 13 9 2
26 1 9 10 0 9 1 9 13 9 9 7 9 0 9 2 1 15 0 13 2 7 14 1 0 9 2
14 3 3 13 9 9 1 0 9 2 15 15 9 13 2
42 0 0 9 13 7 1 9 2 15 4 13 9 9 0 9 2 7 1 0 9 2 15 13 1 2 9 2 7 3 1 9 0 9 2 3 3 0 9 13 0 9 2
18 7 1 15 13 9 9 9 2 10 9 0 3 7 1 9 0 9 2
21 1 10 9 13 3 13 9 2 16 0 9 15 13 2 7 3 9 13 0 9 2
28 10 9 13 0 13 0 9 9 12 9 9 2 7 1 9 1 15 13 13 9 7 13 2 3 13 0 9 2
11 0 9 3 13 0 9 1 9 0 9 2
9 13 9 2 9 15 3 13 9 2
23 10 9 15 1 10 9 13 0 2 7 12 9 13 3 0 9 1 9 7 9 1 9 2
18 7 1 9 1 9 9 2 0 9 7 9 15 13 1 9 7 9 2
61 1 9 9 9 2 15 4 13 15 1 9 9 0 9 2 1 9 2 1 10 0 9 1 9 1 9 2 1 9 13 9 9 9 0 9 1 12 1 12 2 0 9 2 2 15 1 1 9 9 13 1 9 0 9 7 9 9 9 1 15 2
17 13 9 2 16 13 9 3 0 13 9 0 9 1 0 9 9 2
24 16 4 13 0 3 13 9 0 9 7 3 9 9 3 13 1 9 1 10 9 1 0 9 2
19 1 0 0 9 13 9 9 1 0 0 9 2 15 3 3 13 10 9 2
11 0 9 1 0 9 7 0 9 1 9 2
3 11 11 2
2 11 11
5 0 0 9 13 13
13 11 15 13 13 9 9 2 1 9 7 11 7 11
15 9 0 9 13 1 9 12 9 9 2 15 13 0 9 2
23 1 0 12 9 0 9 13 0 9 12 9 9 2 16 1 0 9 3 13 14 12 9 2
13 0 9 11 3 3 13 0 9 0 9 1 9 2
15 1 9 10 2 9 1 9 2 3 13 0 9 0 9 2
15 3 1 9 13 12 9 9 2 3 13 0 12 9 9 2
24 9 1 9 13 0 9 0 0 9 2 9 2 2 0 9 12 0 9 2 1 0 12 9 2
30 0 9 9 13 2 16 9 9 1 9 13 1 0 9 2 12 2 0 1 9 9 7 13 15 10 9 1 0 9 2
15 0 13 7 9 0 2 0 2 9 2 9 7 0 9 2
22 13 0 2 16 11 2 11 7 11 13 13 13 0 9 2 16 4 13 9 10 9 2
32 3 9 0 9 9 9 9 0 9 13 2 16 15 13 0 13 7 16 2 9 13 13 7 3 0 9 9 0 0 9 2 2
14 0 9 4 13 1 9 2 15 13 13 0 9 9 2
32 9 9 1 9 7 0 9 1 0 12 9 13 13 0 0 9 1 11 2 7 3 9 10 9 1 0 9 0 7 0 9 2
14 1 9 9 1 9 13 9 0 9 11 11 1 11 2
17 0 9 11 11 13 9 11 7 13 10 9 1 9 0 0 9 2
31 1 9 13 2 16 11 10 0 9 13 9 9 1 0 9 2 16 4 9 1 11 13 1 9 9 1 11 1 10 9 2
4 9 1 0 9
7 9 9 13 0 9 1 9
29 1 9 13 1 9 3 13 3 9 1 9 3 12 9 9 2 15 13 14 1 12 3 16 3 2 12 9 2 2
23 10 0 9 1 0 9 13 9 2 13 9 7 9 7 1 9 9 13 1 0 9 3 2
7 1 15 15 3 13 9 2
16 9 10 9 13 0 9 7 9 2 1 15 9 9 3 13 2
18 13 1 9 1 0 9 1 0 9 9 2 15 0 9 13 0 9 2
33 1 9 0 9 2 3 16 3 2 13 0 0 9 9 9 11 11 2 3 13 2 3 13 9 9 1 0 9 7 9 11 2 2
19 1 15 13 2 16 9 4 3 13 2 13 9 7 13 3 12 9 13 2
18 16 13 3 16 12 9 9 2 13 1 9 9 0 0 9 9 9 2
9 1 0 9 13 0 9 1 11 2
25 13 0 9 2 3 0 9 1 9 13 0 9 13 9 1 9 9 2 16 3 3 12 9 13 2
19 9 13 9 1 9 7 9 2 15 13 9 2 16 9 1 9 3 13 2
24 3 15 13 2 16 16 0 9 9 13 2 13 0 9 3 1 9 9 7 3 15 3 13 2
19 3 0 9 13 13 1 9 1 12 9 9 2 1 0 9 13 9 9 2
27 9 9 9 7 9 9 11 11 13 2 16 3 0 9 13 9 1 9 0 9 2 9 9 9 7 9 2
13 13 1 0 9 2 0 9 13 1 9 0 9 2
26 16 3 1 9 15 0 9 13 2 3 13 9 1 15 2 16 4 15 1 9 1 9 3 13 13 2
33 1 9 1 9 13 9 2 16 1 12 9 13 9 13 3 14 12 9 0 9 7 1 9 2 16 1 15 13 2 13 9 9 2
17 1 0 11 7 1 11 9 9 13 3 2 9 0 9 7 9 2
21 0 9 1 9 13 0 9 2 7 3 9 9 2 3 16 13 9 2 3 13 2
11 10 9 13 1 0 9 13 7 1 15 2
4 9 1 0 9
27 0 9 0 9 13 0 9 1 9 1 9 0 9 7 0 9 1 9 12 9 9 2 12 9 9 2 2
30 13 1 12 9 0 0 9 11 7 13 15 2 16 1 9 12 9 1 9 15 1 10 9 13 9 9 1 12 9 2
19 1 9 9 9 15 1 12 9 9 13 0 9 2 3 9 9 7 9 2
15 1 10 9 4 12 9 13 1 9 9 1 0 0 9 2
10 9 15 3 13 13 0 9 1 9 2
12 0 12 9 9 4 13 1 9 1 0 9 2
13 12 9 9 9 9 13 13 1 9 9 0 9 2
26 9 3 13 13 0 9 15 2 16 9 1 9 1 9 0 1 9 0 9 15 13 1 12 9 9 2
12 1 12 9 15 13 9 1 0 7 0 9 2
10 0 9 13 13 9 9 1 9 9 2
13 1 0 9 13 0 9 9 9 7 9 0 9 2
11 0 9 2 15 13 9 2 4 3 13 2
13 9 9 13 13 9 0 9 2 15 13 0 13 2
18 1 9 12 0 9 4 13 9 9 0 0 0 9 11 11 7 11 2
15 12 9 15 4 13 9 0 9 9 11 7 9 11 11 2
3 9 1 9
39 2 0 0 9 2 0 9 0 9 2 4 13 2 2 13 3 0 9 9 11 11 1 9 2 15 4 13 9 0 9 0 9 1 0 9 1 0 9 2
28 2 9 0 9 4 3 3 13 7 9 2 16 4 11 13 13 0 0 9 2 4 13 2 2 13 9 11 2
6 9 15 3 13 1 9
14 3 7 3 1 9 9 13 1 9 9 10 9 7 9
15 1 9 10 9 13 0 13 1 9 10 9 9 7 9 2
11 9 0 9 9 13 13 1 12 0 9 2
14 1 0 13 1 9 7 9 0 9 9 1 9 9 2
20 1 9 13 1 0 9 14 12 9 9 2 3 13 1 9 9 2 9 3 2
26 0 9 9 9 2 15 15 7 9 16 0 9 13 3 2 13 9 10 3 0 0 9 9 1 9 2
6 9 7 0 9 0 9
12 9 9 13 0 9 1 2 9 2 0 9 2
21 9 9 1 12 2 9 12 4 1 9 13 3 9 3 0 9 2 3 9 3 2
14 1 9 9 13 3 0 9 0 9 2 9 7 9 2
32 10 9 4 13 3 1 9 0 7 0 9 2 7 15 7 0 9 9 2 7 9 9 2 3 10 9 2 9 1 9 0 2
22 16 13 3 1 0 9 2 13 15 10 9 1 9 0 3 2 7 3 7 3 3 2
11 7 1 0 9 15 13 0 9 0 9 2
9 9 10 9 13 13 9 0 9 2
25 3 1 9 9 3 0 9 9 13 3 0 9 7 3 9 1 0 9 9 1 9 15 13 13 2
23 10 9 1 9 13 14 0 9 2 3 9 1 9 0 9 2 10 9 13 1 9 3 2
21 3 4 3 15 13 2 9 0 1 12 2 9 15 13 3 9 2 9 7 9 2
11 1 9 9 13 1 10 9 1 0 9 2
5 9 9 13 9 9
13 3 1 0 0 9 9 15 13 1 0 9 9 2
37 0 9 9 9 7 3 7 9 0 9 9 11 9 3 13 2 16 9 15 1 0 9 13 10 9 2 16 13 0 0 9 9 1 0 9 13 2
36 9 9 1 9 15 3 1 9 12 9 9 1 9 13 14 12 9 2 1 9 0 9 1 9 14 12 9 7 1 9 0 9 14 12 9 2
38 16 1 9 9 13 9 9 9 2 10 9 15 1 12 2 9 13 3 1 9 2 1 15 1 9 2 1 0 9 0 2 9 2 9 2 13 9 2
19 7 1 10 9 1 9 13 10 9 3 0 7 14 3 13 12 9 9 2
18 14 3 15 3 13 13 2 16 4 13 1 10 9 0 9 9 13 2
23 9 3 13 9 9 11 1 12 9 2 1 9 0 12 9 13 3 0 9 14 12 9 2
23 1 0 9 9 13 0 9 9 3 12 9 7 3 13 1 9 2 16 4 9 9 13 2
35 3 15 13 13 2 16 1 0 9 9 1 12 9 2 15 13 9 3 0 9 16 12 9 1 0 9 2 13 9 1 9 14 12 9 2
23 1 15 0 9 15 13 13 1 0 9 2 15 1 10 9 13 13 0 9 1 0 9 2
26 1 0 9 13 3 0 0 9 9 2 7 15 1 12 9 1 9 1 0 7 1 12 9 1 0 2
20 9 1 12 9 0 9 13 1 12 9 2 1 9 9 13 3 1 12 9 2
3 9 7 9
15 0 9 9 2 15 15 3 3 13 3 2 13 0 9 2
21 1 9 9 9 9 12 2 12 15 1 0 9 13 0 9 9 7 9 1 9 2
63 0 9 2 15 0 9 3 2 3 13 0 9 1 9 0 9 7 9 0 9 2 13 13 2 13 1 9 12 9 1 9 0 0 9 2 1 0 9 12 9 2 7 1 9 2 9 0 1 9 2 0 9 3 12 9 2 1 12 9 1 9 0 2
28 9 7 13 0 2 16 3 2 16 13 9 9 7 9 13 1 10 9 0 9 2 13 13 9 1 15 9 2
7 7 15 13 3 3 9 2
10 1 9 9 13 13 1 9 0 9 2
38 1 12 2 12 2 12 13 3 1 9 0 9 9 2 15 13 15 9 2 0 9 4 3 13 9 2 7 13 0 9 2 3 2 4 9 13 9 2
9 3 1 9 9 4 3 7 13 2
26 13 15 3 9 12 0 9 2 9 12 9 2 1 0 9 1 9 9 2 12 9 1 0 0 9 2
74 1 10 9 4 3 2 1 3 2 13 0 9 1 11 2 12 9 0 9 2 12 0 2 12 0 2 12 1 0 9 2 12 1 9 7 9 2 2 0 9 13 7 1 9 9 12 9 1 0 9 2 12 9 1 9 7 9 2 7 0 9 2 1 12 9 1 9 1 12 9 1 9 2 2
14 13 0 2 16 9 0 9 15 13 7 1 0 9 2
24 1 9 15 3 13 9 0 7 0 9 1 0 0 9 2 7 15 3 1 12 7 12 9 2
15 1 1 9 9 15 7 0 9 13 13 14 1 9 9 2
7 15 15 13 12 2 9 12
7 15 3 0 0 9 9 2
44 13 4 7 3 0 9 2 1 15 0 3 3 3 13 9 2 15 13 10 0 9 1 9 1 0 9 0 9 2 3 3 9 2 10 9 1 9 4 13 3 1 9 2 2
32 0 9 13 13 3 1 9 0 9 0 0 9 1 0 9 7 1 9 9 9 9 9 9 2 7 10 9 9 3 7 13 2
39 1 0 9 10 9 4 13 13 14 9 0 9 2 7 15 1 9 0 9 1 12 9 7 13 4 3 7 0 9 2 7 15 1 9 14 1 12 9 2
30 1 9 3 13 1 9 0 0 9 2 15 13 0 9 9 2 7 7 3 2 9 2 12 5 9 1 0 9 2 2
12 9 9 0 0 9 1 9 15 7 3 13 2
17 10 9 13 3 12 0 9 0 9 2 0 13 14 1 12 9 2
16 13 4 15 9 2 11 0 2 1 0 9 0 0 9 11 2
15 13 15 2 16 1 9 9 9 9 13 9 1 0 9 2
24 2 15 13 13 12 9 12 9 1 0 9 2 15 3 1 9 9 1 12 9 1 9 13 2
17 15 4 1 0 12 9 13 1 11 3 9 16 1 0 0 9 2
18 9 13 7 1 0 9 7 13 2 16 1 9 3 13 1 12 9 2
16 3 2 16 9 4 1 15 3 13 2 7 1 9 9 13 2
19 13 15 2 16 9 13 9 1 9 9 9 7 13 2 3 9 13 2 2
28 10 3 7 3 0 9 13 1 9 2 11 2 15 2 12 2 9 12 2 12 12 11 9 2 2 9 3 3
1 12
2 9 2
8 9 13 2 0 7 0 9 2
18 11 2 0 2 0 9 0 1 9 11 1 11 1 9 7 9 9 2
26 12 9 1 12 9 1 12 9 1 9 13 9 0 9 1 12 2 12 9 1 9 2 0 9 9 2
20 0 9 2 13 1 0 2 9 2 13 15 1 0 9 2 13 0 9 9 2
10 3 0 15 2 12 9 1 12 9 2
20 12 0 9 13 9 2 9 7 9 1 9 2 9 2 9 9 7 9 9 2
7 13 7 13 9 9 11 2
20 1 9 1 9 13 9 2 9 2 0 2 9 2 9 12 2 12 12 11 12
47 9 2 0 9 11 13 2 2 9 2 9 2 9 2 9 2 9 2 0 2 9 2 9 0 2 9 2 9 2 2 0 9 2 0 9 2 2 9 1 9 2 9 2 9 2 2 9
7 0 0 9 1 11 2 11
6 0 9 13 0 9 2
12 9 2 2 12 2 12 12 12 2 12 12 12
1 12
4 0 9 1 11
5 11 2 11 2 2
31 1 0 9 0 9 13 1 9 2 1 9 0 9 10 9 1 0 9 2 9 9 11 11 1 9 0 9 0 0 9 2
14 10 9 3 13 9 3 2 0 15 13 3 3 3 2
10 3 3 4 13 13 0 9 9 0 2
31 13 15 2 16 0 9 0 0 9 11 2 15 4 13 13 0 9 2 13 13 9 0 0 9 1 9 1 0 9 11 2
11 13 4 15 11 11 2 9 0 0 9 2
41 9 11 11 11 1 9 1 0 9 1 0 13 2 16 9 9 2 15 15 13 1 11 11 2 7 10 9 2 3 1 0 9 7 1 9 9 11 2 13 0 2
30 2 16 4 10 9 13 0 9 1 11 2 13 4 15 0 2 0 7 0 9 11 1 15 0 9 2 2 13 3 2
8 13 4 10 9 9 11 13 2
33 2 13 2 3 9 9 11 13 9 1 10 9 9 11 2 15 15 13 1 11 11 2 7 15 3 10 9 1 0 9 3 13 2
31 13 1 15 13 2 7 3 15 13 13 2 16 15 15 16 9 0 0 9 1 10 2 0 9 2 7 15 0 13 2 2
1 9
2 0 9
32 9 1 11 7 11 13 0 9 1 0 9 9 11 2 15 4 15 13 13 9 0 9 2 10 9 13 1 0 0 9 11 2
16 13 12 9 2 16 4 13 2 16 10 10 9 3 13 4 2
2 9 2
22 9 3 13 0 12 9 9 1 0 9 2 16 4 9 12 9 11 13 4 3 13 2
15 1 9 15 3 1 9 12 0 9 13 3 9 1 11 2
39 1 15 7 15 9 2 16 9 11 13 3 13 1 12 2 9 2 16 1 10 9 13 9 11 13 0 9 0 15 3 0 9 2 15 9 13 9 2 2
23 11 15 3 13 13 2 16 9 11 7 11 13 0 2 7 9 1 9 0 9 13 9 2
10 7 11 2 7 11 7 15 10 13 2
36 3 2 14 15 15 15 13 7 13 2 1 9 12 0 0 9 2 15 4 1 0 9 1 11 13 0 9 10 9 2 13 1 9 7 9 2
24 13 2 14 15 7 3 9 13 0 9 11 9 9 1 9 9 0 2 4 13 10 0 9 2
3 9 13 9
9 9 9 9 9 0 9 1 0 9
27 9 7 9 9 9 2 3 13 0 9 0 9 0 9 11 2 3 10 9 7 9 2 0 9 11 11 2
66 13 9 0 9 9 9 2 0 0 9 0 9 9 12 2 9 1 15 9 2 1 9 2 9 2 9 7 9 1 9 2 9 2 9 14 1 0 9 2 2 2 2 2 2 2 7 3 7 9 9 0 2 3 15 2 15 4 13 1 9 2 2 13 11 11 2
40 2 13 0 2 16 0 9 13 3 0 2 7 13 15 1 9 9 7 0 9 2 15 4 13 9 7 13 2 16 15 7 15 15 13 14 14 16 0 0 2
41 12 2 12 9 13 3 0 2 13 4 13 3 12 2 9 9 11 11 2 7 13 14 1 9 12 2 16 14 3 13 9 0 0 9 2 7 1 0 13 9 2
56 13 4 9 3 0 2 0 7 0 2 3 2 11 2 11 2 11 2 11 2 11 2 0 2 11 2 11 2 11 2 11 2 11 2 1 15 2 16 0 13 3 13 2 10 9 2 2 9 9 2 15 4 0 3 13 2
38 13 3 3 0 9 2 16 13 15 12 9 3 1 15 13 9 1 11 11 2 13 15 2 16 10 9 13 1 10 0 0 2 9 2 3 3 2 2
22 9 2 9 2 15 7 1 11 3 3 13 3 3 2 16 0 9 3 0 2 2 2
8 2 13 2 7 13 15 0 2
24 7 0 0 9 15 10 9 13 2 13 15 15 2 7 0 9 3 1 0 9 13 9 3 2
25 9 13 13 2 0 2 7 1 10 9 13 0 9 2 9 0 9 2 9 2 9 2 7 9 2
23 3 14 2 7 9 13 9 2 3 2 3 1 0 9 15 13 13 7 13 3 15 15 2
22 13 15 3 2 7 14 3 4 13 9 0 9 7 9 13 3 10 0 3 0 9 2
12 13 7 2 16 13 1 0 9 7 0 9 2
32 0 9 13 2 12 9 1 0 9 7 9 15 2 3 13 2 13 2 1 15 13 10 9 2 3 15 2 15 1 9 13 2
19 7 9 13 0 12 9 2 3 2 1 9 2 3 9 0 0 0 9 2
11 15 9 10 0 0 9 3 13 1 9 2
11 0 9 13 0 9 2 13 3 1 9 2
28 9 15 3 13 2 3 4 3 13 9 2 15 4 13 13 1 0 9 9 2 3 1 9 10 0 9 3 2
34 9 3 13 1 15 9 2 13 15 2 16 0 2 7 0 2 16 13 1 0 9 0 9 1 9 2 9 15 1 15 13 13 3 2
30 3 7 1 9 13 15 9 2 3 9 0 9 11 11 2 15 15 13 2 16 0 9 13 0 2 2 1 9 2 2
8 13 1 10 9 0 9 13 2
42 13 15 10 9 2 3 9 0 0 9 1 0 0 9 2 7 0 9 2 13 15 3 2 16 4 9 3 0 9 13 1 9 2 1 9 2 2 3 1 0 9 2
15 3 15 13 2 16 3 1 9 9 1 9 15 9 13 2
7 13 0 2 0 2 9 2
26 3 3 14 2 14 15 2 16 1 0 11 11 4 13 11 11 2 10 9 15 13 1 9 13 15 2
2 0 11
19 16 15 13 0 9 9 12 2 9 0 9 13 2 3 15 15 13 1 2
9 0 0 9 11 15 7 3 13 2
20 13 1 0 2 3 0 9 2 3 14 9 0 9 2 15 15 3 3 13 2
9 1 0 9 13 7 9 11 0 2
16 9 0 9 9 13 3 3 0 2 7 13 15 0 0 9 2
19 1 15 15 3 13 9 9 1 3 0 9 9 2 11 7 9 2 11 2
27 0 9 3 13 0 11 7 0 9 13 1 9 11 11 1 9 11 11 11 2 15 15 3 1 9 13 2
16 3 0 13 7 9 0 9 2 15 13 7 1 3 0 11 2
36 7 16 0 3 13 1 9 2 16 0 9 3 13 9 2 3 13 11 10 0 9 2 1 15 1 9 13 7 0 9 7 3 3 0 9 2
20 9 9 12 15 13 14 9 0 9 2 7 3 9 0 9 1 0 9 9 2
2 9 3
10 9 2 11 11 2 0 9 2 9 2
19 2 0 0 9 11 11 13 11 1 9 1 9 0 9 7 0 0 9 2
35 9 2 11 11 2 1 0 9 1 11 13 0 9 9 0 9 11 11 2 12 7 12 2 2 15 4 1 10 9 13 1 0 0 9 2
9 14 1 9 13 13 9 0 9 2
16 9 2 11 2 11 2 11 11 11 13 12 1 0 0 9 2
7 13 1 11 7 11 11 2
18 1 12 2 9 13 0 9 7 10 0 9 3 13 9 11 1 11 2
4 1 15 9 9
34 1 0 9 9 2 0 9 12 2 2 15 13 1 0 9 1 0 9 1 0 7 3 0 9 2 13 1 9 13 9 9 11 11 2
41 1 1 15 2 16 10 9 13 3 16 12 1 0 9 2 1 12 9 13 1 10 9 3 14 12 2 2 2 0 9 2 13 13 9 3 1 10 9 1 9 2
11 11 13 3 9 2 10 9 15 3 13 2
53 0 9 2 9 0 9 2 1 15 9 13 9 2 9 7 10 0 9 1 9 0 14 1 15 9 2 12 1 0 9 13 13 1 9 9 1 0 9 9 9 11 2 3 4 13 16 9 9 9 7 9 2 2
31 7 9 2 15 13 1 9 12 2 1 10 9 13 2 7 13 15 1 15 1 10 9 13 16 1 0 0 9 1 9 2
11 13 15 0 9 2 15 13 16 0 9 2
6 11 11 13 9 9 2
4 0 2 3 2
20 13 15 13 1 15 9 2 3 3 2 7 3 3 3 2 1 0 0 9 2
7 13 15 2 16 9 13 2
4 15 15 13 2
11 15 2 15 3 13 2 13 1 9 3 2
14 1 9 15 13 3 0 9 2 0 15 1 0 9 2
7 9 0 10 0 0 9 2
11 9 1 9 2 15 15 13 1 0 9 2
10 13 15 10 0 9 0 1 10 9 2
12 11 11 13 2 16 3 14 15 13 1 9 2
8 15 9 3 1 9 9 13 2
8 9 13 13 1 12 2 9 2
10 9 13 11 11 2 9 9 12 2 12
10 2 1 0 9 13 10 9 0 9 2
12 3 10 9 13 1 12 9 11 11 1 9 2
22 3 1 9 2 12 2 2 13 11 3 9 2 15 15 3 12 13 2 0 11 11 2
12 4 13 1 3 0 9 9 9 11 1 11 2
42 9 0 9 4 15 13 13 9 9 11 14 3 7 9 12 12 2 9 2 7 3 1 15 11 13 9 2 1 15 13 3 3 2 12 2 9 4 13 13 0 11 2
4 9 1 9 9
28 11 2 11 2 11 13 11 1 11 15 2 16 15 13 1 0 9 9 0 7 13 3 9 9 7 9 9 2
29 1 11 9 13 0 9 1 9 0 9 11 7 9 9 7 9 9 2 1 15 15 1 9 13 0 7 0 9 2
30 14 12 9 9 13 1 0 0 9 9 9 1 0 9 2 3 15 13 13 0 9 9 9 11 7 0 9 0 9 2
16 2 2 10 9 13 11 2 2 13 12 1 9 1 10 9 2
38 0 9 11 1 11 13 1 9 10 10 9 0 2 9 2 0 9 7 0 9 2 9 1 9 2 0 9 7 0 9 2 0 9 7 9 1 9 2
19 1 9 11 11 15 13 0 9 9 1 9 1 0 9 0 9 2 2 2
18 9 15 13 1 0 7 0 9 1 9 1 9 1 9 7 3 3 2
32 0 9 9 9 1 9 9 9 7 9 9 7 3 9 11 11 1 0 9 1 0 2 13 1 9 9 2 13 1 9 9 2
34 0 3 13 0 9 1 9 11 11 1 0 9 13 3 9 7 13 15 0 13 7 9 13 1 9 2 15 1 9 0 9 11 13 2
16 9 0 2 1 15 13 7 9 0 9 7 9 9 2 2 2
25 9 9 2 1 15 15 13 9 11 1 9 0 9 2 1 0 9 7 1 9 9 9 7 9 2
6 2 0 9 2 13 3
11 16 9 11 13 9 2 9 11 3 13 9
26 3 9 1 9 13 3 1 0 9 1 11 0 9 9 2 0 9 2 2 3 15 13 0 0 9 2
20 9 3 13 9 1 11 2 16 9 9 11 13 14 0 9 1 0 9 11 2
18 3 1 0 15 0 9 13 1 11 1 9 1 9 9 2 0 9 2
36 1 9 1 9 4 13 13 15 0 9 3 9 11 2 9 11 2 9 11 2 9 1 11 7 9 11 2 15 15 13 1 9 1 12 9 2
25 1 9 10 0 9 13 1 9 0 9 9 1 10 0 9 11 2 16 4 15 13 1 0 9 2
32 13 15 15 0 2 3 14 15 2 16 0 13 2 16 7 1 0 0 9 9 13 9 1 0 9 2 1 15 15 3 13 2
14 16 4 3 13 1 15 2 16 4 1 0 9 13 2
59 1 9 15 1 0 9 13 9 0 9 9 11 2 3 3 1 0 9 2 7 1 9 1 9 2 13 2 1 9 0 9 2 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 9 0 11 2 11 2 11 2 1 11 2 2
14 3 0 9 13 9 2 2 14 2 13 15 2 13 2
11 1 0 9 13 0 13 9 1 0 9 2
11 7 15 16 15 3 13 14 9 1 9 2
15 13 1 15 9 2 10 9 13 2 13 2 15 15 13 2
9 10 9 1 0 9 3 13 2 2
20 13 10 9 1 10 9 2 16 3 2 16 1 9 1 11 4 15 13 13 2
21 1 9 1 9 4 13 3 0 2 0 9 1 9 9 4 13 1 9 0 9 2
11 9 13 3 1 0 9 2 7 2 2 2
18 2 13 0 13 14 1 12 9 2 4 15 13 13 15 1 12 2 2
23 0 2 9 15 3 13 3 2 3 7 3 1 11 2 1 12 9 13 0 0 0 9 2
11 1 9 1 9 11 9 11 9 3 13 2
38 13 15 2 16 1 9 13 11 2 1 9 4 13 1 0 13 9 1 0 9 11 1 15 2 16 9 0 1 0 9 4 13 13 9 1 9 9 2
30 0 9 4 3 13 1 9 2 11 2 9 2 11 2 11 2 9 2 11 2 11 2 11 2 11 2 0 2 11 2
30 11 10 9 13 2 7 13 2 16 3 1 9 9 11 13 2 2 1 9 3 13 9 2 7 13 15 14 1 9 2
23 13 10 9 1 9 1 9 7 1 9 2 3 16 13 15 2 13 15 10 0 9 2 2
39 1 9 11 3 2 3 13 1 0 9 2 1 15 15 9 13 1 9 9 2 9 11 13 2 2 13 1 3 0 9 2 16 13 15 3 1 0 9 2
12 3 3 15 14 1 9 13 9 10 9 2 2
3 0 9 9
5 11 2 11 2 2
26 1 0 9 4 3 1 9 9 11 12 11 11 1 0 9 13 0 0 0 9 1 0 7 0 9 2
15 3 15 13 10 9 11 11 2 4 9 13 1 12 9 2
18 1 0 9 13 13 12 9 2 15 4 15 13 13 9 1 0 9 2
21 2 3 4 13 13 1 3 0 0 9 1 3 7 3 0 2 2 13 11 11 2
28 0 9 13 3 16 9 1 9 1 3 0 7 0 9 2 1 9 9 1 15 3 13 9 9 1 0 9 2
2 9 3
2 11 2
19 10 9 11 4 0 9 9 13 2 7 10 9 1 0 9 13 3 0 2
9 13 15 3 0 9 11 11 11 2
16 1 10 9 13 10 0 9 1 0 9 0 9 1 9 9 2
18 0 9 1 9 10 9 13 1 11 2 11 13 9 9 9 0 9 2
13 1 10 9 1 10 9 13 0 9 9 9 11 2
44 9 3 11 2 9 0 9 1 9 1 11 7 1 11 2 3 4 1 0 7 1 0 9 13 9 1 10 9 9 2 13 1 9 0 9 1 11 9 2 11 9 1 9 2
15 1 0 9 15 1 9 1 0 9 13 0 9 1 11 2
9 9 9 0 9 7 3 4 13 2
28 1 9 9 9 15 1 9 9 1 11 2 11 2 11 7 1 11 13 13 0 9 1 9 3 12 9 9 2
11 7 0 9 13 3 9 1 9 9 2 12
3 9 1 9
3 11 11 2
34 0 11 11 2 15 13 1 9 1 9 1 3 0 9 1 11 11 2 3 15 13 0 9 9 9 1 9 2 13 1 9 9 13 2
10 13 7 13 2 16 15 10 9 13 2
13 13 15 3 9 0 0 9 1 11 11 11 11 2
17 11 11 15 1 3 0 9 13 3 3 2 16 13 0 9 9 2
28 0 1 0 2 0 9 2 3 4 13 2 13 1 9 2 3 1 9 2 7 13 15 3 13 1 0 9 2
13 1 9 13 1 9 2 3 13 2 1 0 9 2
12 1 9 0 9 13 1 9 2 7 1 9 2
14 0 9 1 0 13 0 9 1 0 9 9 0 9 2
14 11 11 13 3 3 0 0 2 15 1 10 9 13 2
6 9 1 11 1 11 2
2 11 2
36 9 0 11 11 11 1 0 9 13 1 9 0 9 11 11 11 14 13 1 11 2 7 3 0 0 9 13 13 12 9 1 9 1 0 9 2
9 2 11 11 13 0 9 1 11 2
26 13 3 12 9 2 3 15 9 2 3 9 2 13 1 0 9 7 3 13 9 2 2 13 11 11 2
33 11 7 11 15 1 10 9 1 9 9 11 3 4 13 9 1 9 1 0 9 2 7 1 9 2 9 7 3 15 3 13 4 2
13 11 11 15 13 13 1 15 0 9 9 11 11 2
6 9 1 11 13 0 9
7 11 2 11 2 11 2 2
31 0 0 9 2 15 1 9 13 1 9 11 1 11 1 0 9 9 9 12 3 11 2 15 3 1 0 9 3 13 13 2
15 0 9 3 3 13 1 10 9 14 12 9 9 0 9 2
23 1 9 9 13 0 9 7 10 9 13 9 2 0 9 4 3 13 14 1 12 9 9 2
33 9 3 10 9 9 2 9 0 9 7 9 9 2 3 0 0 9 2 13 1 9 7 0 9 2 1 15 15 9 13 0 9 2
14 0 9 13 3 1 0 9 1 9 0 9 7 11 2
39 3 2 16 13 3 9 13 2 9 12 2 12 11 2 11 1 9 9 12 2 12 1 12 9 7 9 0 9 12 2 12 1 11 1 11 13 3 13 2
26 0 9 15 1 0 9 13 1 0 11 2 1 9 11 7 3 0 9 2 3 9 13 12 9 9 2
19 1 9 11 2 3 15 9 13 14 1 9 9 2 13 4 9 13 9 2
10 9 15 13 7 1 9 0 0 9 2
3 9 1 9
7 11 1 11 2 11 2 2
30 0 9 1 9 1 9 9 0 1 11 0 0 9 13 1 9 0 9 0 9 1 12 2 9 13 9 1 0 9 2
20 1 9 13 3 14 12 9 9 0 9 2 1 9 14 1 12 5 1 9 2
17 9 13 9 14 1 12 5 0 9 2 9 13 9 13 1 9 2
23 9 13 3 13 12 5 9 0 9 2 0 9 7 9 13 14 1 9 12 5 0 9 2
13 0 0 9 1 12 9 13 9 1 11 0 9 2
26 9 0 7 0 9 0 9 11 1 11 1 11 13 2 16 1 9 4 9 13 3 12 9 9 3 2
3 9 0 9
2 11 2
44 1 0 9 9 9 11 11 11 9 0 9 9 1 9 0 0 9 1 9 9 1 0 9 13 1 9 2 16 4 9 13 13 0 9 7 3 13 13 1 0 9 9 9 2
21 0 9 9 3 13 7 1 0 9 7 0 9 13 13 16 0 7 0 0 9 2
7 9 1 9 3 11 13 0
2 0 9
2 9 9
3 9 9 9
9 9 1 9 9 0 9 1 11 3
46 1 11 3 13 16 1 9 2 7 3 15 1 9 11 2 3 4 1 0 9 13 0 9 0 15 1 9 11 2 11 2 11 2 13 13 14 0 9 7 0 9 13 9 7 9 2
19 0 0 9 7 0 9 1 0 9 3 13 13 1 0 0 9 0 9 2
27 0 13 1 9 0 9 0 0 0 9 2 15 9 9 11 11 13 1 9 9 1 11 1 0 9 11 2
27 0 12 9 0 0 9 1 0 7 0 9 1 11 13 14 0 9 0 0 9 2 15 7 3 14 13 2
36 1 9 9 2 1 15 13 12 9 1 9 1 12 9 2 1 11 2 0 9 7 11 2 2 13 0 9 1 0 9 11 7 11 2 11 2
49 3 13 3 3 0 9 2 10 0 9 13 1 9 0 12 9 2 16 0 11 9 12 2 15 13 11 11 2 13 14 1 12 2 9 1 9 12 9 1 0 11 12 5 9 2 11 11 11 2
36 11 7 13 14 3 0 9 2 13 3 0 7 0 9 15 1 15 13 2 2 7 3 0 9 2 15 1 9 0 10 0 9 13 10 9 2
56 9 13 12 2 1 12 0 9 11 12 11 7 12 0 11 12 2 1 12 0 9 13 1 0 9 12 12 5 12 11 11 11 2 15 13 3 12 0 9 0 9 1 9 12 5 12 2 12 9 11 7 12 0 9 11 2
16 0 0 9 13 16 3 9 11 2 11 2 15 13 12 9 2
28 0 15 13 13 0 0 9 9 12 11 2 12 1 15 2 9 0 9 11 2 11 2 11 3 13 9 9 2
20 10 11 2 11 7 11 1 2 9 2 11 12 13 0 9 1 9 12 9 2
24 1 0 7 3 3 0 9 13 11 11 0 2 7 3 0 9 7 13 15 9 1 0 9 2
27 9 0 9 7 1 9 13 7 0 9 1 11 2 15 13 3 0 9 9 7 3 3 7 3 0 9 2
16 3 3 15 13 13 2 15 4 13 3 1 0 9 7 9 2
4 9 11 7 11
6 9 11 15 13 1 9
24 0 0 9 1 9 9 1 0 9 7 0 9 13 1 9 1 9 1 11 11 11 1 11 2
12 13 0 9 9 2 7 13 15 3 0 9 2
16 9 13 0 9 1 0 9 11 11 2 15 1 0 9 13 2
6 1 0 9 13 9 2
17 15 0 15 13 11 11 2 15 1 10 9 13 3 1 9 12 2
19 1 9 13 11 11 1 12 2 12 2 12 7 12 1 0 12 9 2 2
19 9 1 9 1 0 9 15 13 2 0 2 1 0 9 1 9 11 11 2
20 1 9 9 0 1 9 1 12 9 13 1 9 0 9 7 1 12 9 13 2
49 13 15 11 2 9 2 2 2 11 2 13 2 2 2 11 2 11 2 2 2 11 2 9 2 2 2 11 2 11 2 2 2 11 2 11 2 2 2 11 2 11 2 7 11 2 11 2 2 2
18 1 9 9 0 2 9 11 7 11 13 1 0 9 7 13 1 9 2
4 9 2 12 2
9 11 2 11 2 2 12 2 12 2
9 11 2 11 2 2 12 2 12 2
8 11 2 11 2 12 2 12 2
9 11 2 11 2 2 12 2 12 2
9 11 2 9 2 2 12 2 12 2
7 11 2 11 2 2 12 2
5 9 9 2 12 2
12 11 2 11 2 11 2 2 12 9 2 12 2
5 11 2 11 12 2
3 11 1 11
29 9 11 11 11 1 11 13 1 9 0 9 1 11 0 9 7 13 12 1 0 9 2 16 11 13 14 11 11 2
12 15 3 13 1 0 9 11 1 11 7 11 2
15 11 2 0 2 11 2 2 12 2 12 2 12 2 12 2
12 11 2 11 2 12 2 12 2 12 2 12 2
15 11 2 0 2 11 2 2 12 2 12 2 12 2 12 2
12 9 11 0 1 9 0 2 9 13 1 15 13
15 11 11 2 0 0 9 1 11 2 13 9 9 0 9 2
12 1 11 1 11 13 9 0 13 9 12 9 2
10 10 9 13 0 9 1 9 1 9 2
32 7 16 3 13 7 0 9 9 11 3 1 11 2 13 15 9 0 9 2 3 0 9 1 9 2 15 13 12 9 12 9 2
26 1 9 9 1 11 15 11 13 1 3 0 9 11 1 11 2 15 13 9 12 9 2 7 3 13 2
4 9 1 9 9
16 15 13 3 10 9 1 0 9 1 0 0 9 9 1 11 2
8 11 9 2 2 13 15 9 2
12 9 13 3 16 15 2 15 4 15 13 13 2
7 11 13 0 3 0 9 2
8 0 9 13 1 10 9 2 2
12 11 11 2 2 13 4 15 13 3 0 9 2
13 11 4 3 13 13 9 2 15 4 15 13 2 2
23 11 11 2 2 13 15 2 16 4 13 13 9 2 16 4 15 3 1 9 1 11 13 2
23 3 1 0 9 4 15 1 9 0 9 13 3 3 2 16 12 1 12 9 13 9 13 2
11 7 1 11 4 13 3 9 0 9 2 2
19 11 11 2 2 1 0 9 3 1 9 13 12 9 2 7 3 14 12 2
22 1 11 13 3 11 11 7 1 10 9 15 13 3 12 1 12 0 9 0 0 9 2
15 13 0 9 2 1 9 13 15 2 13 13 9 7 13 2
14 4 3 13 1 15 2 3 15 15 15 13 13 2 2
21 3 3 13 0 9 1 11 1 11 2 1 11 2 3 2 7 1 0 11 13 11
1 9
5 0 11 2 11 2
9 11 12 2 12 2 12 2 12 2
12 11 13 1 12 9 0 0 9 1 10 9 2
26 11 2 0 9 11 11 1 9 14 1 9 13 11 9 12 2 12 2 12 2 12 2 12 2 12 2
14 9 9 2 11 2 11 12 2 12 2 12 2 12 2
26 0 11 2 1 9 0 9 11 15 13 0 9 2 15 9 4 13 9 11 11 1 9 1 9 9 2
14 3 0 2 10 0 0 9 15 13 9 1 9 9 2
33 11 1 9 1 9 11 11 13 2 3 16 11 2 11 11 2 11 2 11 2 11 2 11 2 9 9 11 7 0 9 11 11 2
26 11 2 0 9 0 0 9 1 0 9 11 11 2 12 2 13 3 13 1 10 9 7 1 0 9 2
10 13 1 15 9 9 9 0 0 9 2
33 0 9 11 11 2 12 2 2 15 1 9 1 9 0 9 3 13 1 9 2 13 2 16 15 1 9 9 4 13 7 0 9 2
25 11 11 2 11 15 9 1 9 1 0 11 13 3 3 2 3 15 7 13 1 0 9 0 9 2
7 0 9 3 13 1 11 2
14 16 9 11 9 13 2 10 9 9 11 15 13 1 9
21 13 9 12 2 9 9 2 9 0 12 2 7 12 2 9 2 7 13 10 9 2
15 11 11 13 9 1 0 11 1 9 12 2 12 2 12 2
16 1 9 13 0 11 1 11 1 9 12 2 12 2 12 9 2
16 0 9 11 11 1 12 9 2 13 14 12 9 2 2 12 2
16 11 2 11 11 2 7 11 2 11 2 12 12 9 2 12 2
8 11 2 11 2 12 2 12 2
7 11 2 11 12 2 12 2
8 11 2 12 11 11 2 12 2
4 9 2 12 2
6 11 11 12 2 12 2
6 11 11 12 2 12 2
3 11 12 2
35 0 9 13 9 11 11 11 1 9 1 0 9 11 1 9 1 0 12 2 12 7 9 1 0 2 11 11 2 11 2 2 12 2 12 2
19 9 1 11 12 2 12 15 0 2 0 9 13 1 9 1 9 1 9 2
15 1 0 9 15 13 10 9 12 2 9 0 9 1 11 2
2 1 9
35 1 9 1 11 12 2 12 2 12 2 12 2 13 0 2 11 1 0 9 9 1 9 12 1 0 9 2 3 11 2 11 2 11 2 2
30 11 2 0 9 11 2 13 9 1 9 11 1 0 9 12 2 12 2 12 2 12 2 1 10 9 1 9 0 9 2
15 0 9 2 11 2 11 12 2 12 2 12 2 12 2 2
13 3 1 15 15 13 11 9 0 11 1 12 9 2
33 9 1 11 2 11 2 11 12 2 12 2 12 2 12 2 2 1 12 2 9 2 11 2 11 12 2 12 2 12 2 12 2 2
4 3 1 12 12
10 0 9 11 2 11 2 11 12 2 12
19 3 1 12 12 13 3 1 9 0 2 9 1 10 0 9 1 9 11 2
10 1 11 13 1 12 9 1 12 9 2
7 12 9 13 1 9 3 2
9 0 9 15 13 3 1 12 9 2
13 1 0 9 1 12 9 13 7 9 9 11 0 2
16 13 15 3 1 3 0 9 2 11 2 0 2 11 2 11 2
13 7 3 10 9 15 13 1 9 1 12 2 9 2
14 1 9 13 9 11 2 11 3 13 9 7 11 13 2
19 9 15 1 0 9 10 9 13 1 9 2 7 3 9 13 1 10 9 2
11 1 0 9 15 13 11 1 9 7 13 2
14 1 11 0 9 3 1 9 2 3 13 1 0 9 2
13 3 0 11 13 1 0 9 0 9 7 4 13 2
43 9 11 2 11 2 11 2 11 2 11 2 11 2 9 2 11 2 0 2 11 2 11 2 9 2 11 2 11 2 11 2 11 11 2 11 11 2 11 2 11 2 11 2
7 9 2 12 2 7 12 2
4 11 2 12 2
4 11 2 12 2
4 0 2 12 2
4 11 2 12 2
4 11 2 12 2
2 11 2
7 9 2 11 2 11 2 2
6 9 2 12 2 12 2
6 9 2 12 2 12 2
6 9 2 12 2 12 2
4 9 2 12 2
14 12 2 12 2 12 2 12 2 12 2 12 2 12 2
6 9 3 13 2 2 2
13 1 0 11 15 3 1 9 13 1 0 7 0 2
14 1 15 15 13 13 2 1 10 9 15 3 15 13 2
9 11 0 13 0 9 3 0 9 2
13 13 9 2 16 4 1 15 1 10 10 9 13 2
10 0 13 2 13 13 2 13 2 13 2
10 1 9 15 7 3 1 0 9 13 2
21 3 15 3 0 9 11 2 11 2 11 13 2 16 10 9 0 9 15 3 13 2
35 2 13 3 0 0 9 1 15 2 16 4 9 13 9 7 10 9 9 2 2 13 10 0 9 1 11 0 0 9 2 3 9 11 11 2
16 3 4 9 11 13 2 16 13 1 9 0 9 1 0 9 2
9 6 2 13 1 0 9 2 2 2
4 1 9 15 13
9 0 11 2 1 9 0 13 14 12
18 11 11 11 13 3 0 9 0 9 11 2 15 3 13 1 0 11 2
15 3 13 1 10 9 1 9 12 2 16 3 13 3 3 2
26 7 1 9 13 12 1 0 9 0 0 9 9 3 2 1 9 12 2 9 2 3 13 10 0 9 2
27 10 9 13 1 9 1 9 0 11 0 0 9 11 2 15 1 0 0 9 1 0 11 13 0 12 9 2
25 1 0 9 0 9 13 2 11 2 2 3 4 11 13 2 14 1 9 2 3 13 10 9 11 2
18 1 9 7 13 12 9 1 9 12 2 12 2 12 2 12 7 12 2
32 3 13 11 1 0 11 12 9 2 1 15 1 12 13 1 9 3 7 3 13 9 13 9 11 11 2 15 3 13 12 7 2
11 0 9 13 13 0 9 1 9 0 9 2
12 13 0 2 16 3 15 13 3 1 0 9 2
13 1 9 13 12 1 9 0 9 3 0 9 11 2
36 1 0 9 0 2 11 2 0 13 1 9 13 11 2 11 2 11 2 11 2 11 11 2 11 7 1 9 9 11 2 11 2 11 7 11 2
10 9 0 9 13 1 0 9 0 9 2
15 3 1 9 11 2 15 15 13 1 9 0 9 11 11 2
5 3 9 1 11 2
20 4 13 0 0 9 2 1 15 1 9 13 1 11 1 0 9 1 0 11 2
9 3 15 1 15 13 10 0 9 2
34 1 0 9 0 9 4 13 9 11 11 2 13 16 9 2 12 2 7 11 11 2 15 1 11 13 11 1 12 9 7 13 0 9 2
16 11 15 13 9 3 13 7 1 9 1 0 11 15 11 13 2
13 13 3 0 2 3 15 13 11 11 2 12 2 2
20 1 0 9 2 3 1 9 7 9 1 9 9 13 11 7 11 2 13 3 2
10 1 3 0 9 3 13 7 0 9 2
18 7 3 1 9 15 13 11 11 11 7 15 13 13 0 14 1 9 2
13 1 9 9 4 13 1 15 13 0 0 11 11 2
15 1 0 9 1 11 13 2 16 13 1 0 9 0 9 2
7 11 13 1 9 9 11 2
18 3 15 13 1 0 11 7 1 9 0 9 3 13 1 0 0 11 2
15 1 9 3 13 3 0 9 0 2 9 2 9 7 11 2
8 9 2 11 2 11 2 2 2
6 15 15 13 1 9 9
6 11 15 13 1 11 2
21 0 9 1 0 11 0 0 9 13 2 16 13 9 7 1 0 9 1 0 9 2
24 11 11 2 0 9 2 13 1 9 11 11 0 9 1 11 12 2 12 9 9 11 7 11 2
15 1 9 3 1 9 13 1 9 9 9 0 9 11 11 2
21 0 9 0 9 0 9 13 2 16 9 11 13 9 9 11 2 11 2 9 11 2
25 9 7 13 2 11 15 13 1 11 7 1 9 13 1 9 2 1 12 2 9 15 13 13 11 2
12 13 15 2 16 0 9 9 13 13 0 9 2
15 3 2 1 9 13 7 10 9 16 11 2 11 7 11 2
5 11 13 1 9 2
15 1 11 13 1 0 9 11 11 7 1 9 1 0 9 2
19 1 9 12 2 12 13 9 9 0 9 11 2 15 13 1 9 1 11 2
17 11 11 2 15 15 13 1 9 1 11 2 13 3 14 1 9 2
11 0 9 7 13 2 16 1 9 13 0 2
17 15 9 9 9 7 13 2 16 13 9 1 9 1 9 9 13 2
12 3 3 9 0 1 9 0 9 11 1 9 2
18 0 15 13 2 16 1 0 9 13 9 9 1 9 1 3 0 9 2
13 9 13 1 9 1 9 7 9 13 0 1 9 2
5 9 13 1 11 2
13 1 0 9 13 9 1 0 9 11 1 11 11 2
15 1 9 2 1 15 9 13 1 0 9 2 15 9 13 2
12 13 9 0 9 2 1 15 13 7 9 9 2
3 11 13 2
27 0 9 13 1 9 11 11 0 9 11 11 2 7 3 2 16 3 13 15 2 16 1 9 13 1 11 2
24 1 0 9 10 9 13 3 1 9 1 11 14 0 9 2 1 0 15 1 9 11 3 13 2
1 3
3 9 13 9
28 11 13 12 1 0 9 9 2 13 3 9 1 9 12 2 0 0 0 9 2 15 15 13 1 10 0 9 2
29 9 0 9 11 0 0 13 13 7 13 0 0 9 1 9 3 2 16 4 15 13 0 9 0 11 0 1 11 2
6 0 9 2 1 7 1
45 1 9 9 2 15 13 10 9 0 9 9 2 11 2 11 13 2 16 13 0 2 16 4 9 11 2 1 15 4 9 11 13 13 0 2 13 9 1 0 9 7 0 0 9 2
12 1 0 9 15 1 9 9 13 9 0 9 2
9 0 9 13 9 9 11 11 11 2
12 1 15 3 0 9 13 9 1 9 0 9 2
19 3 13 0 9 9 9 2 3 9 13 9 9 3 15 13 1 0 9 2
26 7 9 11 13 9 2 16 4 11 13 0 9 1 0 7 0 9 11 2 15 4 13 0 0 9 2
12 1 9 1 9 0 9 9 13 3 0 9 2
31 1 9 2 15 13 1 9 1 9 11 1 9 11 11 2 15 1 9 10 9 3 13 0 9 11 7 9 11 11 11 2
13 2 10 9 1 9 13 7 13 3 1 0 9 2
9 13 15 13 7 13 14 0 9 2
22 15 9 13 1 15 1 10 9 0 7 0 9 1 9 1 0 0 9 13 9 9 2
55 2 1 9 1 9 2 15 15 13 2 16 9 2 13 10 9 2 7 10 0 9 2 2 11 11 13 2 16 2 9 13 9 9 9 0 9 2 9 7 9 7 1 0 9 13 9 0 9 1 9 0 0 9 2 2
55 3 13 9 2 1 15 14 9 15 9 13 13 1 15 2 16 9 2 15 13 2 13 9 9 1 9 2 7 10 9 13 9 0 9 0 9 11 11 2 2 9 0 9 13 3 0 9 2 16 13 9 10 9 2 2
5 3 4 9 13 2
1 9
13 9 0 9 0 9 13 3 1 9 11 0 9 2
12 1 10 9 4 13 0 0 9 1 9 11 2
12 1 9 4 15 13 2 15 1 15 14 13 2
16 3 2 13 3 9 7 9 9 2 15 3 13 10 0 9 2
31 7 13 1 15 13 7 15 0 2 15 13 11 9 2 9 1 12 9 2 9 0 9 2 9 0 9 7 9 2 2 2
15 3 9 13 2 16 1 10 9 13 7 0 9 0 9 2
4 9 13 13 0
10 1 9 9 11 11 1 9 11 11 11
3 2 11 2
19 13 4 13 9 2 15 0 9 13 9 11 11 1 9 0 9 9 11 2
17 2 1 0 9 13 3 1 9 9 10 9 2 15 13 3 0 2
12 13 15 3 9 1 3 0 9 9 7 3 2
10 1 10 9 9 13 3 1 9 12 2
22 3 15 15 13 13 3 3 2 7 15 14 1 9 0 9 11 2 15 4 13 9 2
16 9 9 15 7 13 7 1 0 9 2 3 0 15 11 2 2
18 11 11 15 13 15 2 16 9 13 0 13 9 2 3 15 15 13 2
18 2 1 0 9 13 0 9 0 13 15 10 9 9 2 1 15 13 2
15 1 9 2 15 4 13 2 15 1 10 9 1 9 13 2
23 16 1 15 3 13 15 3 2 1 9 15 15 13 2 16 13 0 11 1 9 0 9 2
30 11 11 1 0 0 9 13 0 9 11 9 2 1 15 13 2 16 15 0 9 13 13 3 2 3 15 1 15 13 2
10 13 4 7 2 16 0 9 13 9 2
21 1 9 1 10 9 13 9 3 0 7 0 3 1 9 2 9 2 0 9 2 2
15 0 9 0 0 9 3 13 2 16 13 0 9 10 9 2
18 7 15 11 11 13 1 15 2 16 10 9 3 13 9 9 7 9 2
16 2 1 15 15 13 2 13 1 15 13 14 3 1 0 9 2
22 0 9 1 0 0 9 13 9 9 0 9 1 9 2 15 15 3 13 13 0 9 2
15 10 9 7 3 13 1 0 0 9 7 13 3 0 2 2
11 1 0 9 9 1 11 9 11 11 13 2
5 15 13 9 9 2
6 2 1 9 3 13 2
11 9 7 0 9 13 1 10 3 0 9 2
32 10 9 11 3 13 1 15 9 2 7 13 15 1 9 2 3 3 3 2 16 11 11 13 0 9 0 9 11 11 11 2 2
21 3 13 9 11 11 2 16 15 13 2 0 9 2 1 9 0 0 9 1 9 2
17 2 15 0 13 2 3 16 4 15 1 10 9 13 1 0 9 2
22 3 15 1 0 0 9 13 1 9 9 3 0 0 9 7 10 9 1 9 11 11 2
32 11 11 13 2 16 4 13 4 11 11 13 2 7 16 13 9 9 11 2 1 15 15 13 9 1 0 9 7 3 1 15 2
8 10 10 9 7 3 13 2 2
4 11 13 9 9
6 11 11 1 0 9 9
2 11 2
54 15 0 9 7 9 13 13 1 9 2 16 16 13 1 9 9 0 0 0 9 2 11 2 2 13 2 16 4 15 1 10 9 13 0 9 9 2 2 13 3 11 11 2 15 4 1 10 9 13 4 13 9 11 2
29 1 9 1 11 11 3 13 10 0 9 2 16 11 4 15 13 13 1 0 9 2 15 13 1 0 9 0 9 2
11 2 13 4 15 13 9 2 15 9 13 2
22 15 13 9 2 9 2 0 9 7 9 9 9 3 7 3 2 2 13 11 2 11 2
13 0 9 11 15 1 15 13 13 1 9 0 9 2
18 10 9 13 3 7 9 9 1 11 2 15 15 16 9 11 4 13 2
18 3 2 3 13 2 13 0 13 1 9 7 9 9 11 1 0 9 2
32 1 9 2 16 11 13 0 9 1 11 11 2 3 3 13 10 0 9 9 11 11 2 13 2 16 13 13 1 9 10 9 2
19 2 16 9 0 9 0 9 1 11 4 1 10 9 13 9 2 2 13 2
19 1 9 11 13 1 0 9 9 9 11 11 11 2 11 2 7 0 9 2
25 3 13 1 0 9 1 9 0 9 0 9 2 13 1 9 9 13 0 0 0 9 7 0 9 2
28 1 9 11 2 11 4 13 9 0 9 1 9 9 13 10 9 9 11 2 3 4 7 13 13 1 0 9 2
17 13 2 16 1 9 2 3 4 13 11 2 13 0 7 0 9 2
19 11 2 11 3 13 2 16 1 0 9 15 13 7 3 1 9 9 11 2
13 0 9 1 9 0 9 4 7 13 13 1 9 2
17 11 2 11 13 2 16 13 3 2 0 7 9 9 9 0 9 2
30 1 10 9 4 1 9 0 9 0 9 13 13 9 9 1 0 9 2 0 9 0 9 3 2 2 9 9 1 9 2
15 1 9 0 9 9 4 13 1 10 9 13 3 0 9 2
19 1 0 9 4 3 13 13 0 7 0 9 2 0 9 7 9 0 9 2
2 11 13
2 11 2
26 1 9 2 16 4 0 9 13 9 0 9 9 7 3 15 13 2 13 13 9 0 9 11 0 11 2
12 13 15 3 1 9 9 0 9 0 9 11 2
28 1 10 9 15 3 13 2 16 2 16 15 13 9 13 9 2 13 3 13 0 9 11 1 9 10 9 2 2
26 9 13 1 0 0 0 9 0 9 0 1 0 9 11 1 0 11 2 1 15 14 12 9 13 0 2
19 13 2 16 16 0 9 13 0 9 3 13 2 13 0 0 7 0 9 2
9 9 1 9 0 11 2 11 2 2
23 1 0 2 0 9 15 3 13 9 12 0 0 9 7 9 0 7 0 9 1 0 11 2
28 12 9 2 0 9 1 12 9 13 3 12 9 9 2 1 0 9 15 4 10 9 13 3 3 1 0 9 2
26 0 9 1 9 12 12 9 1 9 13 3 1 9 9 9 0 9 7 9 12 0 9 7 12 9 2
35 0 9 1 9 0 9 7 9 13 9 0 2 0 9 2 15 13 9 9 2 0 9 11 2 0 9 0 11 2 0 9 7 9 9 2
13 1 9 11 9 13 1 9 0 9 0 13 9 2
12 12 9 7 9 3 9 13 0 0 9 0 2
3 9 1 9
5 11 2 11 2 2
16 0 9 1 0 9 0 7 0 9 13 3 1 11 9 11 2
33 3 13 3 9 9 11 9 2 13 15 1 0 0 9 1 9 0 9 2 1 15 9 13 0 0 9 1 9 0 7 0 9 2
14 1 9 13 0 9 2 1 0 9 4 13 12 9 2
12 9 13 9 0 13 1 9 9 7 0 9 2
3 9 1 9
6 0 11 2 11 2 2
22 0 0 9 13 12 9 0 9 1 9 0 11 9 1 9 1 11 7 0 9 11 2
25 13 15 1 9 9 0 2 9 2 11 0 11 7 9 0 1 9 7 9 1 9 13 9 11 2
8 3 15 1 9 13 12 9 2
6 9 4 13 1 9 2
2 9 13
5 11 2 11 2 2
18 9 0 9 13 1 9 1 11 12 0 9 1 11 7 12 10 9 2
12 0 9 9 13 2 9 13 1 11 1 11 2
12 16 9 0 9 13 11 2 13 3 9 0 2
19 9 13 1 9 12 1 15 2 13 1 0 9 2 1 15 13 0 9 2
7 1 9 4 13 0 9 2
3 9 1 9
5 11 2 11 2 2
19 0 9 1 11 13 1 0 0 9 1 9 1 9 11 1 9 9 11 2
12 1 9 1 9 1 9 13 1 0 9 9 2
7 9 15 3 13 1 9 2
9 3 15 3 13 0 1 0 9 2
8 1 9 9 13 1 0 9 2
3 9 1 9
7 11 1 11 2 11 2 2
36 9 2 15 13 1 9 7 13 1 9 2 13 9 0 0 9 1 0 9 9 2 12 1 11 2 13 4 1 15 12 2 12 2 12 2 2
28 9 9 11 2 11 2 1 11 1 0 2 9 2 13 3 2 16 13 1 9 7 13 15 3 1 0 9 2
20 1 0 9 12 9 13 1 9 12 0 9 1 11 7 0 12 9 4 13 2
1 9
3 13 9 2
19 1 9 1 0 9 0 9 1 9 13 12 0 7 12 0 9 1 11 2
18 1 0 9 13 1 0 9 9 7 0 1 15 13 0 9 1 9 2
4 9 9 3 13
5 11 2 11 2 2
22 3 0 0 9 13 0 9 9 11 9 0 9 9 2 11 11 1 9 0 9 11 2
31 1 9 2 3 3 4 13 9 0 9 1 0 9 0 9 2 15 3 3 13 9 0 9 0 9 0 9 0 1 11 2
18 1 9 0 9 9 15 3 13 13 9 1 9 9 1 9 12 9 2
15 0 9 4 13 13 9 2 3 3 13 3 1 10 9 2
8 0 9 13 0 9 3 12 2
24 13 0 9 2 16 9 1 9 1 11 15 1 9 13 9 11 2 7 1 11 13 9 9 2
3 9 13 9
24 0 9 1 12 9 0 9 13 1 0 9 1 11 9 0 9 11 1 0 11 9 11 11 2
9 3 1 12 9 14 13 0 9 2
49 12 9 0 9 13 2 16 1 9 9 15 1 9 2 16 13 0 9 3 2 0 9 3 13 1 15 1 9 2 3 15 13 13 2 10 15 13 9 1 9 2 7 3 15 13 9 1 9 2
10 13 7 1 9 9 1 9 7 9 2
14 12 0 9 13 0 9 1 0 9 1 0 0 9 2
17 12 1 15 3 3 13 1 12 9 2 0 13 0 9 1 9 2
6 12 13 9 7 9 2
10 3 15 1 0 0 9 13 1 9 2
18 2 12 9 3 13 9 2 2 13 15 3 12 1 0 9 1 11 2
21 2 12 15 3 13 12 9 7 13 15 13 2 0 3 13 9 1 0 11 2 2
15 0 9 0 9 1 9 3 13 2 16 15 13 7 13 2
5 2 13 15 9 2
22 16 4 15 13 9 2 14 4 15 9 13 15 2 2 13 15 12 1 9 0 9 2
21 2 9 13 9 9 7 0 9 13 7 1 15 2 2 13 10 9 9 9 11 2
15 2 9 0 9 13 3 0 9 16 3 7 13 15 13 2
15 13 15 3 9 2 1 9 7 1 9 15 13 9 9 2
17 3 15 13 0 9 2 10 9 13 1 0 9 2 0 1 0 2
20 9 9 13 0 9 2 7 13 7 0 9 9 1 0 9 7 1 9 2 2
10 0 0 9 15 9 1 11 4 13 2
17 3 7 13 0 2 3 13 9 2 7 13 1 9 13 0 9 2
2 0 9
16 0 9 15 1 15 1 9 0 9 13 0 9 1 12 9 2
24 1 9 13 9 12 9 2 9 13 9 12 1 9 12 2 1 9 9 12 9 12 10 9 2
34 0 0 9 2 0 0 9 2 4 13 1 9 2 3 1 0 11 13 9 3 14 1 12 9 2 16 11 13 3 12 9 2 9 2
20 0 0 9 3 1 0 9 13 1 10 9 9 3 0 9 0 9 1 11 2
17 1 0 0 7 0 9 13 13 9 0 9 1 9 1 0 9 2
44 1 10 9 15 13 9 2 1 9 9 7 13 1 9 2 3 7 9 2 0 9 12 7 12 2 0 9 12 7 12 2 9 9 3 9 2 3 7 1 12 9 2 9 2
8 9 1 0 9 0 0 9 2
16 9 2 13 15 2 13 3 9 2 3 3 9 1 9 13 2
28 9 0 9 13 1 0 13 10 9 2 3 0 9 11 4 4 13 2 7 13 1 9 0 9 7 0 9 2
19 13 15 15 1 9 9 0 9 0 9 2 9 2 9 2 9 7 9 2
2 0 9
2 0 9
2 0 9
12 3 1 0 9 15 3 13 1 0 0 9 2
15 13 9 1 9 2 9 2 13 15 0 9 7 0 9 2
54 0 13 2 16 15 13 1 9 1 15 2 16 10 10 0 9 1 0 9 13 1 9 1 9 2 1 15 15 13 1 0 9 2 7 1 9 0 9 13 9 9 2 13 9 7 9 1 9 7 13 9 0 9 2
24 1 10 9 3 9 9 7 15 2 15 15 13 2 13 9 10 9 7 13 3 7 0 9 2
25 13 15 3 13 2 16 1 0 0 9 13 9 9 7 9 16 15 0 9 7 9 1 15 0 2
14 10 0 0 9 13 13 10 9 13 7 13 10 9 2
17 9 0 0 9 2 16 13 9 7 13 3 13 2 13 9 9 2
10 1 10 9 13 7 0 9 0 9 2
33 16 4 15 1 9 13 2 13 15 3 9 1 0 9 9 0 9 1 2 12 0 2 9 2 2 16 4 10 9 4 13 3 2
40 7 16 9 0 9 13 9 2 15 1 15 13 1 0 7 0 9 2 13 3 9 16 10 0 9 7 2 13 2 14 2 16 9 1 9 7 9 0 9 2
19 9 0 0 9 13 9 9 2 9 9 7 9 9 9 2 15 15 13 2
34 1 10 9 13 13 13 1 9 9 0 9 2 16 15 15 2 15 15 15 13 2 13 2 16 9 15 13 2 7 13 1 15 9 2
13 10 9 4 13 13 13 16 9 1 0 9 9 2
33 9 1 0 9 7 9 2 15 13 0 2 4 3 13 4 13 16 9 0 9 7 10 0 9 1 9 1 9 16 9 0 9 2
19 1 9 0 9 4 9 0 9 13 9 2 16 13 13 1 9 0 9 2
38 13 2 16 13 1 9 0 7 0 2 15 13 0 1 10 9 7 13 15 13 0 15 2 15 13 7 15 3 2 7 15 15 3 2 16 13 9 2
33 7 7 15 2 15 4 15 0 0 9 1 10 9 13 2 4 13 1 9 2 7 4 4 13 3 1 10 9 9 1 0 9 2
9 0 0 9 15 10 9 13 4 2
19 13 15 7 13 2 16 3 13 13 2 16 4 15 13 9 1 10 9 2
22 3 13 15 3 13 2 15 4 15 13 13 2 16 4 15 7 0 9 13 15 0 2
27 9 13 7 0 2 13 2 14 15 2 16 13 1 15 10 9 2 13 15 1 9 7 0 0 0 9 2
8 13 15 2 14 2 7 14 2
5 9 13 9 0 9
11 0 9 9 12 13 7 3 9 0 9 2
4 13 13 9 2
14 1 11 3 13 9 2 3 4 1 10 9 9 13 2
21 6 2 15 13 0 9 13 9 2 15 15 2 1 10 9 7 9 2 13 9 2
14 7 15 14 9 0 9 2 7 3 7 9 0 9 2
20 15 2 16 13 3 1 9 9 10 9 14 0 9 2 13 3 0 9 9 2
26 10 0 0 9 3 13 9 13 0 9 2 16 15 13 13 2 3 1 9 2 16 9 13 3 13 2
8 16 9 15 10 9 13 13 2
12 13 7 9 2 16 0 9 1 9 13 0 2
21 13 3 9 1 9 1 9 2 15 13 3 12 1 9 1 0 9 1 9 9 2
18 0 9 4 13 1 9 9 2 15 4 1 12 0 9 13 0 9 2
6 7 16 9 9 13 2
17 3 13 9 0 9 2 16 4 13 9 9 2 15 4 9 13 2
12 13 2 14 15 0 2 13 4 13 0 9 2
8 15 13 0 9 1 9 9 2
17 1 9 13 0 3 13 12 9 2 2 0 9 2 2 0 9 2
7 11 13 13 12 0 9 2
26 15 13 2 16 1 11 13 13 12 9 2 12 0 2 12 0 7 12 0 2 7 3 12 7 12 2
25 10 9 13 3 1 9 0 9 2 13 2 14 16 0 9 0 9 11 2 3 13 0 9 13 2
15 13 12 0 9 2 7 15 7 9 1 9 7 9 9 2
52 1 0 9 2 16 13 9 9 1 9 2 13 9 1 15 2 16 2 9 7 11 13 9 1 0 11 2 2 11 11 2 2 9 2 13 15 15 2 2 13 0 9 7 0 9 1 15 3 13 0 9 2
19 13 2 14 9 9 1 12 0 9 2 3 13 1 9 9 0 1 11 2
33 1 0 9 13 3 12 9 2 9 7 13 0 2 16 4 15 12 9 13 1 10 9 2 9 2 9 2 1 0 9 13 15 2
22 9 4 13 9 1 9 9 2 7 4 13 0 0 9 1 0 9 0 1 9 9 2
15 9 2 13 15 0 9 9 2 9 9 2 9 0 11 2
10 9 2 13 13 9 1 0 9 9 2
10 15 15 13 9 2 13 9 3 0 2
29 11 2 7 0 0 0 9 2 13 2 16 13 1 10 9 1 0 9 2 15 13 1 11 1 9 9 1 11 2
4 15 15 13 2
32 9 2 16 4 1 11 13 13 0 9 2 7 2 0 9 2 2 1 15 11 13 2 13 9 0 9 13 3 0 0 9 2
31 11 13 2 16 9 11 13 9 1 9 0 9 2 0 9 13 0 16 12 9 0 0 9 7 0 9 13 12 9 9 2
10 3 15 13 9 9 2 0 9 3 2
16 15 13 3 0 9 2 16 0 9 1 0 0 9 13 0 2
5 15 1 15 13 2
9 9 9 4 13 3 3 0 9 2
18 0 9 9 7 4 3 13 1 15 2 10 0 0 9 4 9 13 2
27 1 9 9 2 15 13 9 1 11 2 13 13 9 9 3 15 2 15 4 13 1 0 2 0 9 2 2
22 3 0 9 1 0 9 2 9 9 9 1 12 9 1 0 13 13 1 9 9 9 2
17 13 15 9 3 12 9 2 7 9 0 9 13 9 1 0 9 2
39 9 0 9 2 12 1 0 0 9 11 11 13 2 16 0 9 0 11 13 0 9 2 0 9 15 3 13 3 13 9 0 9 16 0 9 1 0 9 2
24 3 2 16 9 1 0 7 0 9 13 15 2 16 0 9 1 9 10 9 13 13 0 9 2
17 3 1 10 9 4 3 13 0 9 0 0 9 1 0 0 9 2
16 7 7 0 9 1 11 13 0 9 7 0 9 9 7 9 2
9 0 9 13 0 13 1 0 9 2
23 0 9 2 9 1 2 0 9 2 13 13 3 1 9 2 4 2 14 11 13 0 9 2
18 9 15 13 3 13 1 10 0 9 1 10 9 7 9 1 0 9 2
3 13 9 2
18 14 2 16 1 3 0 9 2 16 13 9 9 2 13 13 3 9 2
5 13 13 1 9 2
11 14 2 16 15 15 9 1 9 13 13 2
12 9 13 13 11 2 16 4 13 9 10 9 2
5 13 0 9 9 2
10 14 2 7 16 15 1 9 13 9 2
12 9 3 13 0 9 2 3 15 15 3 13 2
4 15 1 9 2
19 9 0 9 13 13 0 9 1 15 2 15 13 9 1 0 7 0 9 2
4 13 0 9 2
10 3 13 9 1 9 1 11 7 11 2
5 15 15 13 13 2
5 9 7 9 9 2
16 9 0 1 0 9 13 0 9 2 14 15 15 13 7 14 2
23 2 9 13 9 0 9 2 3 13 9 11 7 13 15 3 15 0 2 0 0 9 2 2
1 9
1 11
2 11 12
4 11 11 1 9
28 0 9 11 11 0 15 3 16 11 11 1 0 9 13 3 3 1 12 1 10 11 7 9 9 1 0 9 2
3 0 9 9
2 11 2
2 9 2
2 11 2
38 9 1 9 0 9 11 7 0 9 15 13 0 9 0 9 0 9 1 11 2 15 15 1 9 13 1 0 9 11 7 1 0 9 2 15 15 13 2
11 13 3 14 0 9 2 16 9 9 13 2
30 0 9 0 1 9 13 2 0 2 7 14 0 2 2 16 13 0 9 3 0 2 13 1 11 0 9 9 15 11 2
9 11 4 13 13 1 9 9 9 11
5 13 15 9 11 9
2 11 2
26 2 16 9 0 11 4 13 9 0 9 0 0 9 2 3 13 10 9 1 9 11 0 7 0 9 2
11 11 13 13 3 7 1 9 10 9 2 2
20 13 15 9 9 9 11 9 1 9 1 0 9 9 0 9 11 11 1 11 2
6 9 13 9 0 9 2
27 13 9 2 16 16 4 11 13 11 16 0 2 13 4 15 2 0 9 1 9 10 10 9 1 11 2 2
24 2 0 9 15 13 13 3 3 7 15 15 13 13 10 9 1 0 9 2 2 13 11 9 2
15 9 9 13 3 9 1 9 0 9 1 0 9 3 7 9
38 9 1 0 9 0 9 7 9 0 9 3 0 9 2 15 4 13 1 9 9 2 13 12 1 0 9 9 0 9 1 11 1 9 1 0 0 11 2
17 3 13 1 9 0 9 3 2 16 4 10 9 13 3 0 9 2
11 3 4 1 0 9 1 9 13 0 9 2
27 10 9 13 0 9 9 9 0 9 13 9 1 0 9 2 15 14 1 9 12 13 1 9 12 9 0 2
14 1 12 1 0 9 3 3 0 11 13 0 9 9 2
16 1 9 9 4 3 9 13 1 0 9 1 9 7 9 9 2
20 9 9 3 13 0 12 9 2 16 4 3 7 1 9 13 9 1 10 9 2
33 13 3 0 0 9 1 9 0 9 1 9 9 2 15 4 13 9 12 9 3 0 9 2 9 2 9 7 3 3 7 0 9 2
22 10 9 13 0 9 9 13 9 9 7 13 9 9 2 15 3 1 9 0 9 13 2
16 1 0 9 13 9 7 0 9 3 9 0 9 1 0 9 2
24 13 15 2 16 15 9 11 11 3 13 9 0 9 11 1 11 2 16 4 10 0 9 13 2
31 0 9 9 13 3 1 0 0 9 14 1 0 9 9 1 9 7 13 10 0 9 2 3 1 9 1 0 9 1 11 2
23 16 3 9 1 9 13 3 7 14 2 3 13 9 2 16 13 1 9 0 9 1 9 2
5 1 11 15 3 13
5 11 13 9 1 9
2 11 2
19 11 7 11 15 3 3 13 1 9 9 2 15 13 1 9 13 1 9 2
19 11 13 2 16 0 0 9 13 3 9 1 10 9 1 9 11 3 11 2
9 11 7 13 2 16 9 13 11 2
28 0 9 15 3 13 1 0 9 1 9 1 9 9 2 15 4 1 11 13 0 9 0 9 1 9 0 9 2
14 9 13 0 9 1 2 9 0 7 0 9 11 2 2
11 1 10 9 13 11 1 9 3 0 11 2
20 9 11 1 11 15 13 3 9 0 9 2 15 1 9 13 9 1 10 9 2
24 0 9 13 9 12 1 0 9 2 15 15 1 9 1 9 13 13 9 9 1 9 1 11 2
12 9 15 1 10 9 3 1 0 9 13 9 9
8 0 9 2 9 14 1 0 9
22 16 15 1 9 0 2 0 9 3 13 9 2 4 13 9 16 0 11 2 3 11 2
28 11 15 3 1 9 1 11 3 1 9 13 0 9 0 9 2 3 1 9 0 0 9 7 1 9 0 9 2
13 0 1 0 0 9 13 2 7 3 11 11 13 2
23 9 1 9 9 0 9 15 13 3 2 3 16 11 1 0 9 1 0 9 13 15 14 2
38 3 1 10 9 13 3 0 9 2 2 13 2 1 0 13 11 1 11 15 7 0 12 0 9 3 13 1 0 9 9 2 0 9 2 1 15 2 2
7 3 13 7 1 9 11 2
14 1 15 13 1 0 9 13 2 3 14 15 13 2 2
54 7 3 15 2 3 1 11 2 13 1 9 12 2 7 12 2 9 1 0 9 9 11 1 11 7 9 11 11 0 9 0 9 15 2 16 13 13 0 9 9 7 9 2 2 0 2 9 10 9 1 12 0 9 2
29 11 7 11 13 0 9 14 1 11 1 12 9 2 7 3 3 1 11 2 16 13 0 9 0 9 10 0 9 2
32 9 2 0 1 9 0 9 2 1 15 4 12 2 9 13 1 0 9 13 11 15 14 3 11 2 13 1 11 9 0 9 2
5 15 13 0 9 2
23 3 13 2 14 1 0 9 2 16 1 0 2 0 9 13 0 9 0 11 13 14 3 2
47 3 7 3 0 9 1 12 9 11 10 9 13 0 2 9 2 2 16 11 14 13 9 1 0 11 2 3 15 3 13 3 1 9 1 0 9 9 7 1 9 0 9 9 1 9 9 2
17 1 0 9 13 7 3 0 9 2 1 15 13 1 9 7 9 2
14 3 1 0 0 7 0 9 13 13 14 3 0 9 2
19 13 1 15 2 16 9 1 9 11 13 0 16 0 9 1 0 0 9 2
21 3 1 0 9 10 9 15 3 13 0 9 2 15 13 3 0 0 9 0 9 2
14 3 15 13 3 0 9 3 0 9 7 9 0 9 2
36 1 0 0 9 2 1 9 1 11 7 11 2 4 3 10 9 13 3 16 9 9 1 0 9 2 2 7 3 15 9 3 13 2 2 2 2
31 15 3 2 16 0 0 9 13 9 1 9 2 0 9 2 2 15 4 13 4 9 12 13 16 9 1 9 0 0 9 2
24 9 11 7 11 1 0 9 4 1 0 2 3 7 3 0 11 3 13 1 2 0 9 2 2
16 0 1 15 3 13 1 12 2 9 12 1 11 1 0 9 2
37 13 13 9 2 16 7 0 9 9 4 13 2 9 9 2 2 7 9 0 9 1 0 9 13 3 0 2 1 15 15 13 7 0 9 1 9 2
40 13 2 16 9 1 9 0 0 9 1 12 2 9 12 2 15 4 3 13 3 1 12 9 7 15 4 1 9 13 9 9 3 11 2 9 0 9 3 13 2
15 1 15 13 1 9 0 9 2 15 4 13 14 0 9 2
15 0 9 2 1 15 11 13 3 3 2 13 3 3 0 2
15 13 2 16 3 2 16 4 15 13 13 7 0 9 9 2
5 0 9 13 1 11
8 13 15 3 3 3 1 9 12
2 11 2
15 11 13 13 13 15 10 0 9 1 0 9 1 0 9 2
13 13 15 9 0 9 9 2 15 15 13 4 13 2
24 10 9 13 13 0 9 11 11 1 9 1 9 0 9 11 2 15 4 13 1 12 2 9 2
29 1 9 2 16 11 4 1 10 0 9 13 2 13 15 9 1 0 9 1 11 7 11 2 13 9 0 9 9 2
8 13 0 9 9 2 7 9 2
11 1 9 11 15 3 13 12 7 9 9 9
7 11 2 1 10 9 2 2
15 2 13 2 16 1 9 13 15 2 15 15 13 10 9 2
13 7 15 13 2 13 7 4 13 14 1 9 2 2
36 13 15 1 0 0 9 0 9 11 11 1 11 2 12 2 2 9 2 15 3 10 9 13 9 0 9 1 0 9 2 1 15 13 3 13 2
34 9 0 9 2 15 4 1 0 9 13 0 9 2 13 9 11 11 2 16 13 10 9 1 0 9 2 15 1 9 13 9 1 9 2
23 0 9 10 9 13 9 0 9 1 11 11 11 2 9 0 9 2 15 13 0 0 9 2
31 11 14 1 0 9 13 9 9 2 1 0 9 0 11 3 12 9 9 2 1 9 0 9 2 0 9 7 14 0 9 2
20 1 10 9 9 13 1 9 0 9 11 11 2 10 9 2 9 7 0 9 2
15 1 9 0 9 15 3 3 13 3 12 7 9 9 9 2
47 2 15 9 2 15 4 13 1 11 11 11 2 10 9 7 9 1 9 0 9 2 13 3 0 7 15 14 13 2 16 0 9 13 3 3 9 0 9 16 9 2 2 13 1 15 9 2
37 9 3 13 3 2 7 11 4 3 3 3 13 2 16 4 15 9 13 2 3 13 0 9 2 1 10 9 13 0 0 9 1 15 7 10 9 2
7 15 7 11 3 13 13 2
15 0 9 3 13 1 9 7 9 2 1 15 13 0 9 2
33 1 10 9 3 0 9 2 11 11 2 12 2 2 13 3 16 9 9 2 14 12 9 2 1 0 0 9 2 15 1 9 13 2
35 0 0 9 13 1 0 9 13 2 15 2 16 13 10 9 2 13 9 9 2 15 4 13 1 15 2 16 13 9 13 9 2 7 14 2
19 1 0 9 13 7 9 0 0 9 2 15 3 3 13 9 1 0 9 2
25 1 15 3 13 0 9 2 16 13 13 14 1 9 7 13 9 1 0 9 1 9 10 0 9 2
26 13 3 0 2 7 13 14 0 9 2 1 15 15 13 13 1 10 2 1 9 3 0 2 0 9 2
33 9 0 9 15 13 1 15 2 16 9 3 13 9 1 9 2 16 4 13 1 10 9 2 15 13 0 13 0 9 1 12 9 2
25 3 0 9 13 1 9 11 2 14 2 12 9 2 3 1 12 3 2 16 13 1 9 9 0 2
12 1 9 4 3 1 9 1 9 13 12 9 2
8 1 0 9 15 4 13 1 9
5 3 3 13 11 11
2 11 2
26 1 9 0 11 4 3 13 9 13 9 0 9 11 11 2 16 1 0 0 9 3 3 13 0 9 2
18 9 1 9 1 10 9 13 12 9 0 0 9 7 10 9 0 9 2
10 9 0 11 13 1 9 3 12 9 2
13 1 9 11 11 1 9 9 13 3 12 12 9 2
13 9 1 11 1 9 11 10 9 4 14 13 9 11
2 11 2
27 9 0 0 9 13 13 0 9 12 0 9 11 2 7 4 15 1 10 9 13 9 11 1 10 9 9 2
12 13 15 9 0 0 9 1 9 11 2 11 2
24 0 9 15 1 11 3 13 2 16 9 9 11 11 13 9 1 9 0 1 0 9 1 9 2
21 13 9 3 1 15 2 16 10 9 13 13 9 0 9 1 11 1 9 0 9 2
36 0 2 0 9 1 0 9 2 15 3 13 0 9 0 9 7 9 0 9 1 12 9 2 13 13 9 9 0 9 11 1 11 1 9 9 2
24 1 9 9 10 9 4 1 10 9 1 0 9 13 0 9 9 11 2 15 13 3 1 11 2
26 11 2 15 1 9 9 13 0 0 9 2 3 13 2 16 9 0 0 9 11 15 1 10 9 13 2
9 9 11 13 1 9 1 11 3 11
5 9 9 1 11 13
4 11 2 11 2
14 1 9 0 9 1 11 7 11 13 9 3 0 9 2
14 13 15 15 1 9 11 2 15 4 3 13 1 11 2
28 9 2 15 13 0 0 9 11 11 1 10 0 9 0 11 2 13 1 9 0 9 2 15 4 13 0 9 2
19 1 9 13 9 2 16 0 2 0 9 15 13 3 1 0 9 0 11 2
24 0 9 4 3 13 7 1 9 9 2 16 0 9 7 9 1 9 13 0 2 13 9 9 2
27 13 15 3 1 15 2 16 4 9 11 13 9 13 1 9 0 9 7 16 4 3 13 9 1 0 9 2
12 11 13 2 16 9 13 1 9 15 0 9 2
8 0 9 9 7 13 0 9 2
14 9 9 0 9 0 11 1 11 13 1 10 9 13 2
24 13 15 7 13 1 0 9 2 15 13 13 11 7 9 1 11 7 11 2 13 15 1 9 2
27 0 9 11 2 15 13 13 3 3 1 11 0 3 10 9 11 2 13 3 13 9 1 9 1 10 9 2
27 1 9 9 13 1 11 12 2 9 3 0 9 1 0 9 2 15 3 13 1 10 9 3 16 0 9 2
6 9 1 9 13 0 2
5 9 11 1 9 11
2 11 2
25 0 9 7 9 2 0 3 1 0 2 0 2 9 0 0 9 2 13 1 0 9 3 1 9 2
26 16 15 13 1 9 13 11 7 11 2 3 4 13 11 7 11 2 15 13 3 0 9 9 0 11 2
41 15 2 15 15 13 1 11 2 13 1 0 0 9 0 9 2 13 3 0 9 0 11 7 13 2 16 9 1 9 9 2 15 13 3 1 9 2 13 1 9 2
10 11 13 13 2 7 16 15 10 9 13
2 11 2
14 11 13 9 1 9 0 9 1 11 7 10 0 9 2
25 13 15 0 9 9 7 0 9 11 11 1 9 0 9 0 11 2 15 3 13 1 11 1 11 2
26 2 0 9 9 11 1 0 9 15 7 1 10 0 9 1 0 2 0 9 13 2 2 13 0 9 2
23 0 9 13 9 2 16 9 11 7 0 9 1 11 15 4 13 9 0 11 1 9 13 2
22 13 3 0 9 0 9 1 0 9 2 15 9 9 1 0 9 0 9 2 13 2 2
7 1 11 13 3 10 9 9
5 13 15 3 1 11
2 11 2
18 1 12 0 9 7 12 11 4 13 1 9 1 9 1 9 0 11 2
7 13 15 1 9 0 9 2
30 1 10 9 15 1 9 13 3 9 11 1 9 11 2 15 13 1 9 0 11 2 0 9 2 15 13 3 1 11 2
24 12 9 4 13 7 12 0 13 1 0 0 9 0 2 3 1 9 2 2 15 13 0 9 2
4 9 9 13 0
4 0 9 1 11
2 11 2
17 9 9 0 0 9 11 1 9 11 13 7 9 1 0 9 0 2
21 1 9 9 11 3 9 0 9 2 10 9 13 9 2 3 13 1 9 0 9 2
24 9 2 15 15 13 1 10 3 7 3 0 9 2 4 1 0 9 13 0 9 1 0 9 2
27 10 9 13 4 13 0 9 1 1 10 0 0 9 2 1 0 9 15 13 0 9 0 9 9 0 9 2
29 1 0 9 13 9 11 1 9 1 9 14 12 9 2 1 15 9 13 9 1 9 7 1 9 1 0 9 9 2
22 9 11 11 13 1 9 0 9 2 16 4 13 1 9 9 9 7 13 0 0 9 2
7 9 9 4 13 13 12 2
19 1 11 9 13 3 12 9 7 13 0 9 1 9 12 7 12 9 9 2
18 9 2 15 13 12 1 0 9 1 9 11 2 13 1 9 12 9 2
4 9 1 11 2
30 12 9 4 13 7 12 0 13 1 9 1 9 1 0 9 9 1 0 0 9 2 1 15 13 0 0 9 0 9 2
5 13 15 0 9 2
4 0 9 13 2
28 0 9 11 2 0 0 9 1 9 9 1 10 9 7 9 2 13 1 9 9 0 9 11 11 1 10 9 2
7 9 1 9 13 1 0 11
2 11 2
31 1 12 9 3 0 9 1 11 15 1 9 1 9 13 13 9 9 1 9 2 1 15 3 13 1 12 9 1 12 9 2
13 9 13 0 9 7 13 0 9 9 7 0 9 2
13 9 13 10 0 9 2 1 15 12 13 7 13 2
17 12 1 0 9 13 0 9 1 9 3 2 16 13 13 0 9 2
19 1 3 0 9 15 9 13 13 9 1 0 9 0 9 9 1 0 9 2
6 12 9 0 9 13 2
11 11 9 9 2 9 1 0 11 0 9 13
2 11 2
11 0 9 3 3 13 0 9 0 11 11 2
13 1 0 9 4 1 9 13 12 7 12 0 9 2
8 0 9 15 13 12 9 13 2
15 9 15 13 0 9 2 7 9 0 7 0 3 13 0 2
26 3 1 9 13 13 1 9 9 9 2 1 15 15 13 0 9 1 11 2 11 9 9 11 7 11 2
31 9 13 1 0 9 3 1 0 2 0 9 2 3 1 0 11 2 0 9 1 0 9 2 15 13 9 7 9 0 9 2
5 1 11 15 3 13
7 13 3 1 9 3 12 9
2 11 2
14 1 0 9 1 11 7 0 9 11 4 13 12 11 2
23 13 15 3 1 0 9 0 9 2 15 15 13 1 0 0 9 11 2 10 9 11 11 2
24 13 3 2 16 0 9 13 13 15 1 15 2 16 4 4 13 0 9 9 1 10 0 9 2
28 1 10 9 13 3 0 2 16 4 11 13 9 9 0 9 11 2 15 15 13 2 0 9 2 7 13 9 2
30 0 9 9 13 2 16 1 12 2 9 2 3 1 9 13 9 2 13 1 9 12 9 0 9 7 0 12 4 13 2
4 9 9 4 13
2 11 2
4 9 9 4 13
2 11 2
16 9 9 0 9 0 9 11 3 1 0 9 13 1 0 9 2
15 9 13 9 9 7 16 9 13 9 0 9 7 12 9 2
13 1 9 7 13 0 2 16 15 9 13 1 9 2
29 1 9 13 9 1 0 7 11 2 0 9 1 9 9 2 3 15 1 0 9 13 9 1 0 0 7 0 9 2
12 1 0 9 1 9 13 9 1 0 0 9 2
7 1 9 4 13 7 11 2
4 11 13 1 9
2 11 2
2 11 2
2 11 2
39 3 0 9 0 9 1 11 13 2 16 12 5 11 13 13 2 14 2 7 12 5 2 14 2 1 9 2 15 12 2 9 13 1 9 0 9 1 11 2
17 12 9 0 9 3 13 9 0 9 0 9 1 0 9 0 9 2
24 9 13 9 1 0 0 9 7 9 9 13 1 9 2 16 9 9 4 13 11 1 9 11 2
22 2 13 0 13 0 11 2 16 0 11 2 2 13 15 2 3 2 7 2 3 2 2
20 9 11 11 3 13 2 16 13 2 14 2 4 13 1 9 1 11 7 11 2
8 11 13 9 1 0 9 1 11
8 4 1 15 13 7 1 0 9
2 11 2
15 11 13 9 1 9 0 9 1 11 2 7 10 0 9 2
51 1 9 1 0 9 9 11 1 0 9 0 9 2 0 9 2 11 11 13 9 10 0 9 15 2 16 9 13 9 1 9 1 0 11 2 1 15 11 13 1 9 0 9 1 9 0 1 9 1 11 2
26 13 3 0 9 0 9 1 0 9 2 15 9 9 1 0 0 9 1 0 9 0 9 2 13 2 2
7 11 11 13 9 0 9 2
2 11 2
7 11 11 13 9 0 9 2
2 11 2
16 12 1 0 9 0 11 11 11 13 1 0 9 9 0 9 2
12 13 15 9 10 9 1 0 0 9 11 11 2
16 0 9 0 0 0 9 7 1 9 1 0 9 10 9 13 2
34 11 11 1 9 1 0 9 0 9 11 13 2 16 1 0 9 1 0 9 15 13 1 10 9 0 9 2 9 0 0 9 11 11 2
14 9 1 9 15 3 13 1 2 9 0 9 11 2 2
7 3 13 9 2 13 13 2
24 1 9 0 0 9 11 11 2 0 1 9 1 11 1 0 0 11 2 13 3 0 0 9 2
9 3 12 0 9 3 13 1 9 2
7 13 9 15 13 0 9 2
14 1 10 2 9 2 15 13 9 1 9 0 0 9 2
9 3 15 0 9 13 10 12 9 2
15 9 0 9 1 0 9 0 11 1 0 12 9 3 13 2
15 1 0 9 0 1 0 9 13 3 1 12 9 9 3 2
10 3 10 15 15 13 1 0 9 12 2
28 1 15 0 13 3 1 12 9 7 3 15 10 2 0 0 9 2 13 13 1 9 0 12 2 0 9 2 2
12 3 9 2 15 1 0 9 13 2 13 0 2
29 3 3 13 0 9 9 0 2 1 0 9 15 13 1 0 9 1 0 0 9 0 0 9 2 3 3 0 9 2
18 1 9 10 9 13 9 3 13 2 7 3 15 1 9 13 13 9 2
21 3 1 15 13 1 9 0 2 7 16 15 1 0 13 9 2 3 13 0 9 2
10 1 0 9 15 3 10 9 3 13 2
27 3 13 1 9 1 9 0 11 0 9 11 11 2 9 13 1 9 1 9 9 2 9 13 7 9 13 2
38 3 16 13 9 2 15 0 9 13 0 9 3 7 3 2 7 16 3 13 1 9 2 13 15 0 9 1 0 9 1 9 2 1 15 13 3 13 2
22 9 0 9 15 1 0 9 13 1 10 9 2 16 15 15 3 13 13 7 0 9 2
27 11 7 11 2 9 2 1 10 9 13 1 0 9 9 2 3 3 13 9 1 9 1 9 0 0 9 2
23 9 1 10 9 13 7 0 9 0 9 7 0 9 12 9 2 15 13 3 1 10 9 2
22 1 9 0 9 9 13 9 2 9 0 9 11 7 11 13 0 9 1 0 9 2 2
25 1 9 9 13 1 0 9 7 9 9 0 9 2 15 13 12 9 1 0 9 1 0 0 9 2
29 4 3 13 0 9 1 15 2 16 4 9 2 1 10 9 1 0 9 13 2 13 1 0 9 1 9 13 9 2
24 1 0 9 4 7 1 9 9 13 13 7 10 9 2 15 0 9 1 9 0 9 13 3 2
21 9 13 3 15 2 16 0 9 1 10 9 9 9 1 1 9 9 3 7 13 2
19 11 13 2 16 9 1 9 1 0 9 13 7 0 9 0 15 0 9 2
34 15 13 10 9 7 13 10 9 3 15 2 16 13 7 13 9 1 0 9 12 9 7 1 9 15 1 9 13 2 1 9 0 9 2
8 10 9 13 3 3 3 0 2
53 16 15 0 0 9 13 3 13 7 15 9 0 0 9 13 9 9 2 4 9 9 0 15 10 9 15 3 3 13 1 9 10 0 9 2 13 9 2 2 2 0 9 0 2 13 9 2 2 1 9 9 11 2
13 1 0 9 0 9 1 0 11 13 3 12 2 9
14 3 15 14 11 1 9 10 0 9 13 0 9 11 2
19 9 13 1 11 11 11 2 0 0 9 2 15 4 9 9 13 12 0 9
3 9 1 11
5 11 2 11 2 2
19 1 9 0 9 4 1 0 9 13 9 0 0 9 1 9 0 9 11 2
13 11 13 1 0 7 0 9 9 1 0 0 9 2
18 16 0 3 13 0 9 1 9 1 9 2 15 13 0 9 0 9 2
13 2 9 2 1 15 4 13 2 3 13 1 11 2
18 3 13 9 2 13 14 2 16 0 9 0 9 13 0 12 9 9 2
11 13 4 12 9 1 11 13 1 0 9 2
19 0 9 13 9 2 15 15 3 13 2 2 13 15 0 9 11 11 11 2
1 9
3 9 15 13
34 13 9 0 0 9 7 3 3 13 9 2 16 9 11 7 0 9 11 11 15 13 13 9 0 9 9 0 9 16 0 1 0 9 2
27 3 2 3 3 15 13 3 1 10 0 9 1 9 0 9 2 7 7 3 2 16 13 3 12 9 9 2
5 13 15 1 0 2
17 0 9 15 13 2 16 16 4 13 10 9 1 0 9 0 9 2
32 13 15 0 9 2 16 9 0 3 3 13 13 3 3 2 16 4 15 0 9 13 2 16 15 3 15 13 7 13 0 9 2
14 0 9 15 3 13 3 0 7 13 0 9 0 9 2
17 9 10 9 11 1 10 9 13 1 9 15 0 0 9 0 9 2
12 10 9 15 13 3 13 0 9 9 1 11 2
16 15 15 3 13 9 15 0 9 2 15 13 0 9 9 9 2
17 1 10 0 9 15 15 13 9 1 9 9 1 0 7 0 9 2
16 1 0 9 15 13 9 9 0 2 0 9 0 9 9 11 2
32 12 1 15 13 3 9 9 11 11 11 2 11 2 15 1 0 9 11 11 7 11 11 13 0 9 2 7 2 1 9 11 2
7 13 7 11 0 1 9 2
10 15 1 15 13 0 9 2 4 13 2
14 16 7 1 10 9 13 0 9 1 9 7 0 9 2
24 1 0 7 0 9 13 15 3 0 9 2 0 9 7 9 9 1 0 9 1 2 0 2 2
11 10 9 3 13 1 0 9 0 0 9 2
18 3 3 2 16 15 13 9 0 9 0 0 9 1 9 9 0 9 2
17 9 3 10 2 16 4 1 0 9 0 9 13 4 9 3 13 2
2 11 11
3 1 0 9
50 2 0 9 13 3 9 9 1 9 11 7 13 3 13 7 1 15 2 2 3 3 13 1 0 9 3 1 0 9 2 9 13 15 2 12 1 0 9 9 2 9 11 7 9 0 9 0 11 11 2
31 13 3 1 12 1 9 9 2 16 7 0 9 1 9 1 9 11 13 1 9 9 2 7 3 13 1 0 2 0 9 2
42 13 14 0 2 16 0 9 9 9 9 0 9 13 7 3 0 9 0 0 9 1 9 0 9 2 16 3 9 9 9 11 2 11 7 11 1 9 9 1 0 11 2
39 3 1 0 9 11 11 15 13 0 9 1 15 2 15 13 13 11 11 2 0 9 15 3 13 10 9 0 9 7 13 1 9 0 11 1 3 0 9 2
23 13 3 10 9 2 16 15 9 10 9 3 13 1 9 2 16 15 11 11 13 1 9 2
21 1 9 9 9 4 3 3 0 7 0 9 13 3 13 10 0 9 1 0 9 2
33 10 9 7 13 9 12 0 9 2 3 0 9 13 0 9 0 0 9 7 13 15 13 3 1 0 2 16 0 9 1 0 9 2
21 7 3 3 3 0 0 9 1 11 3 13 1 9 13 0 9 1 0 15 9 2
22 9 9 10 9 13 3 0 2 7 3 1 0 9 7 3 0 11 4 13 13 9 2
47 7 3 13 9 9 2 3 3 9 11 2 11 2 11 2 3 13 1 0 9 11 7 11 9 12 0 9 1 9 2 16 4 3 9 9 11 11 13 9 7 9 9 0 9 1 0 2
27 16 13 15 13 2 13 15 3 9 11 2 15 3 13 1 11 0 9 2 16 15 3 13 9 0 9 2
24 7 3 15 13 2 16 0 0 9 1 0 0 9 15 13 13 1 9 3 1 9 0 9 2
19 3 4 10 0 9 13 1 15 0 16 0 7 0 9 0 9 0 9 2
2 11 11
7 9 9 11 2 11 2 2
25 9 1 9 2 15 13 9 1 11 11 2 1 11 2 13 3 1 0 9 13 0 9 1 11 2
18 1 9 13 11 11 2 12 9 9 9 2 15 1 15 13 1 9 2
30 0 15 13 2 16 9 2 15 15 1 15 13 3 1 9 3 7 1 0 9 15 13 9 2 13 1 9 1 9 2
9 3 13 9 2 16 4 13 9 2
16 1 9 13 13 2 16 9 11 11 2 13 13 1 0 9 2
14 1 9 13 13 2 16 9 11 11 2 13 13 1 0
4 0 9 4 13
8 9 0 9 1 9 13 0 9
16 9 12 1 12 13 3 1 0 0 9 9 0 9 9 11 2
9 1 12 0 15 12 9 13 9 2
52 1 9 0 9 15 1 0 13 2 2 15 2 9 0 2 2 2 2 3 1 9 0 9 7 0 9 1 9 0 9 0 2 2 2 2 3 15 2 9 0 9 2 13 15 2 2 2 1 10 9 2 2
33 3 1 9 9 0 9 11 11 13 9 2 1 15 15 13 2 16 9 1 0 9 13 1 15 0 2 7 7 1 15 13 13 2
16 13 2 16 0 9 1 9 9 13 1 9 1 9 9 9 2
7 1 9 11 13 11 11 2
25 13 2 16 1 9 13 0 9 7 16 9 13 10 0 9 2 16 10 9 13 13 0 0 9 2
17 13 2 16 0 9 15 10 9 13 1 0 9 1 1 0 9 2
8 1 10 9 3 13 11 11 2
26 0 9 11 11 2 11 2 13 9 2 16 15 15 9 9 13 1 9 2 15 4 13 9 1 9 2
31 11 11 1 9 1 9 12 0 9 13 2 16 13 3 13 14 9 9 2 7 7 9 9 2 15 9 11 7 11 13 2
14 1 0 9 13 3 9 0 9 7 11 1 0 9 2
22 0 9 1 10 9 13 9 11 2 15 13 9 9 16 0 7 1 9 0 9 9 2
18 13 2 16 11 13 9 7 13 15 3 2 16 13 9 3 12 9 2
34 1 9 9 4 13 1 10 9 11 13 9 9 2 15 15 1 12 2 9 12 13 9 12 0 9 7 9 12 2 9 12 9 9 2
9 0 9 10 9 13 9 0 9 2
26 13 15 2 16 10 9 13 14 3 2 16 13 11 2 7 3 2 16 13 15 0 9 0 9 9 2
8 2 9 9 13 1 10 9 2
21 3 13 15 7 9 2 7 0 9 7 9 13 9 2 9 7 9 0 9 2 2
22 13 2 16 15 9 0 9 3 13 2 7 9 2 15 13 11 1 11 2 15 13 2
23 1 10 9 13 2 16 10 9 13 9 1 11 7 11 2 13 9 9 9 9 1 11 2
10 1 9 9 11 13 0 9 0 9 2
15 1 9 15 9 11 11 13 1 9 1 9 3 0 9 2
8 9 13 9 11 2 11 2 2
22 14 9 13 3 3 0 0 9 2 15 1 9 13 14 12 9 9 3 11 1 11 2
26 2 3 1 9 13 1 9 12 2 7 0 9 2 2 13 3 11 11 2 9 0 0 9 1 11 2
13 2 1 9 13 1 9 12 9 1 0 0 9 2
16 9 1 9 7 13 3 0 2 16 13 1 10 9 9 13 2
13 16 4 13 13 2 13 4 9 0 7 3 2 2
10 3 3 3 13 1 9 14 0 0 9
5 9 9 1 9 2
18 0 9 1 9 0 9 4 13 1 9 1 9 9 1 9 0 11 2
19 9 3 13 9 1 11 2 11 2 2 0 2 16 9 13 9 0 9 2
12 4 13 1 0 9 9 1 9 1 9 9 2
4 9 1 9 2
9 12 0 9 13 1 9 0 9 2
11 9 13 7 13 9 1 9 12 12 9 2
12 3 1 9 4 13 12 0 2 12 1 11 2
14 2 11 2 1 9 4 13 12 0 2 12 1 11 2
4 0 9 13 9
5 11 2 11 2 2
9 0 0 0 9 1 11 13 9 2
18 13 1 11 3 1 9 7 13 13 1 9 9 2 13 0 0 9 2
11 9 1 0 9 7 3 13 14 12 9 2
6 10 9 3 13 9 2
18 2 9 1 0 0 9 2 15 13 13 0 10 9 2 13 3 0 2
29 9 2 3 4 13 12 9 2 13 0 2 2 13 15 1 9 3 0 9 1 9 0 9 0 11 11 11 11 2
31 9 3 13 1 9 0 0 9 11 2 16 3 7 9 13 3 9 1 15 2 15 3 9 0 9 13 2 7 15 14 2
38 13 4 15 9 2 11 11 2 0 9 0 9 9 2 11 2 2 0 9 13 1 9 9 9 1 9 0 9 2 9 9 15 3 13 1 9 0 2
10 13 9 9 2 15 3 13 0 9 2
15 2 0 9 2 15 13 12 1 0 9 9 2 13 9 2
9 9 4 13 9 9 0 1 15 2
10 13 0 9 9 0 9 1 0 9 2
20 0 9 1 10 9 4 13 2 16 0 2 15 15 13 1 9 2 4 13 2
29 1 10 0 9 13 13 15 2 13 15 7 1 9 9 7 9 1 9 2 13 9 1 9 1 9 0 0 9 2
9 1 9 0 1 9 3 13 2 2
3 1 9 9
23 1 10 9 13 7 1 9 2 1 15 13 9 9 2 7 1 15 2 15 13 0 9 2
2 1 9
25 1 10 9 4 13 1 9 1 15 2 3 15 10 0 0 3 13 0 9 7 13 3 1 9 2
23 14 2 13 15 13 0 9 2 16 9 13 13 1 0 7 13 15 10 9 9 7 9 2
27 3 2 16 1 10 9 13 9 11 2 0 9 9 7 9 1 11 1 11 2 13 9 1 0 0 9 2
4 13 15 9 2
16 9 9 13 12 9 9 2 7 1 9 15 0 9 13 13 2
23 13 3 3 13 7 9 1 11 11 2 7 15 2 9 9 11 11 2 7 9 1 9 2
7 0 9 13 3 0 9 2
14 3 15 2 15 13 10 9 1 11 0 1 0 9 2
25 3 2 1 9 1 11 1 11 2 13 10 9 2 16 13 3 2 11 2 11 2 11 7 0 2
8 3 15 13 13 2 13 9 2
12 13 15 2 16 4 15 13 1 9 9 13 2
5 13 15 7 0 2
10 10 2 9 9 2 3 13 10 9 2
30 15 4 15 15 13 2 16 4 9 13 2 7 3 13 0 1 15 2 3 13 13 1 10 9 2 7 13 0 9 2
13 7 3 9 13 7 13 7 15 13 13 2 2 2
19 3 4 15 14 13 9 2 15 3 13 0 9 2 7 15 15 13 9 2
33 3 4 15 13 2 16 4 15 10 9 13 15 2 15 4 13 9 11 13 1 15 2 16 0 16 13 10 9 13 13 0 9 2
4 0 9 9 9
51 0 9 9 0 2 9 2 9 1 9 2 0 2 11 1 9 13 1 9 12 9 2 3 14 12 9 2 1 9 1 9 0 9 2 2 1 0 9 1 0 9 3 12 9 2 3 1 12 9 2 2
18 1 3 0 9 11 13 0 0 9 12 9 7 15 1 0 12 9 2
19 9 1 9 0 9 9 13 3 1 12 7 12 9 0 1 9 1 9 2
30 1 10 9 15 0 2 9 2 9 13 3 13 9 9 9 2 0 9 1 9 13 12 9 2 0 13 12 9 2 2
14 1 9 1 12 9 3 0 9 13 3 1 12 9 2
24 9 9 9 4 9 9 13 1 12 9 2 1 9 15 7 13 1 9 10 9 1 12 9 2
30 3 4 1 9 13 9 9 1 9 2 15 0 2 9 2 9 13 1 12 9 2 1 9 7 3 3 1 12 9 2
26 1 9 1 15 9 2 15 3 13 7 0 9 1 9 2 7 1 9 9 9 2 13 3 0 9 2
11 0 9 9 9 1 0 9 13 9 7 9
20 0 9 9 1 0 9 0 2 9 2 9 11 9 13 1 9 9 10 9 2
26 3 1 0 9 9 1 9 2 0 1 0 9 3 1 12 2 9 2 13 10 9 3 0 9 9 2
38 1 0 9 0 2 9 2 11 9 2 15 15 15 3 13 13 1 9 9 3 11 11 11 2 13 0 9 12 9 0 9 11 0 9 9 12 9 2
32 1 10 9 13 13 3 9 9 9 2 1 12 9 1 10 9 2 2 3 7 0 0 9 12 9 1 12 9 9 1 9 2
12 0 9 9 2 1 0 9 2 13 12 9 2
44 1 0 9 9 15 13 2 16 0 9 15 1 0 9 1 12 9 2 15 13 7 3 0 7 13 15 15 13 3 14 0 9 2 4 1 9 11 13 1 12 9 1 9 2
31 0 9 3 1 12 9 9 11 1 0 9 1 9 14 12 9 2 7 15 13 3 0 2 13 1 0 9 1 12 9 2
2 1 9
3 0 9 9
24 9 0 0 9 2 11 2 13 1 0 9 0 9 12 0 9 2 1 10 4 13 12 9 2
9 13 15 3 0 9 11 11 0 2
26 0 9 4 13 1 9 1 12 9 1 12 9 9 2 16 3 1 0 9 13 9 1 9 12 9 2
24 9 4 13 3 1 9 9 2 9 7 0 9 7 9 0 9 2 3 4 13 0 0 9 2
22 3 11 1 0 9 0 9 13 7 13 1 9 9 9 0 9 1 9 12 9 9 2
10 13 12 9 1 9 3 12 9 9 2
32 13 4 15 9 2 11 11 2 1 0 9 0 0 9 11 2 10 9 4 13 9 11 13 13 0 9 9 11 1 12 9 2
10 13 15 2 16 11 13 13 10 9 2
15 2 15 13 9 10 9 1 0 9 2 13 3 9 9 2
23 11 13 9 0 9 7 3 9 9 13 0 2 16 1 9 13 3 12 7 12 9 2 2
5 0 2 7 3 0
11 12 9 1 0 9 1 12 2 9 0 9
15 13 0 9 1 9 2 15 13 1 0 9 1 0 9 2
12 0 9 13 0 9 1 0 9 12 2 12 2
8 9 11 0 9 0 2 9 2
15 0 0 9 1 0 9 13 0 9 1 0 9 0 9 2
9 9 9 1 12 9 13 12 9 2
23 0 0 9 0 9 15 13 1 12 5 2 1 9 2 9 2 9 2 3 1 12 5 2
11 9 15 3 13 1 9 1 9 9 9 2
18 1 0 9 15 1 10 0 9 13 12 2 0 9 9 9 1 11 2
11 1 9 13 0 9 2 9 7 9 9 2
32 9 13 13 9 1 11 11 1 11 7 1 9 9 9 11 9 13 1 0 9 9 1 10 9 1 9 0 7 0 0 9 2
4 0 9 11 2
23 0 9 1 3 12 9 13 0 9 2 15 13 0 7 0 9 1 9 0 7 0 9 2
18 9 15 13 14 1 0 9 2 7 13 15 7 10 9 3 1 11 2
15 1 10 9 13 0 9 1 11 0 0 9 1 0 9 2
20 1 11 11 2 9 9 9 2 4 13 9 1 0 9 13 9 12 9 9 2
3 11 11 2
16 0 9 1 12 9 15 13 0 9 0 7 3 7 0 9 2
16 1 0 9 13 9 3 12 9 1 9 0 9 7 0 9 2
18 1 9 9 11 11 0 9 4 1 0 9 13 13 3 12 9 9 2
14 10 0 9 13 9 13 1 9 9 7 9 0 9 2
7 13 0 1 9 3 0 2
7 9 1 9 9 13 9 9
14 1 12 2 9 15 13 9 9 1 9 1 0 9 2
6 3 13 9 0 9 2
15 13 3 0 2 16 1 0 9 13 1 0 9 0 9 2
15 9 11 7 9 7 4 1 9 14 12 9 13 0 9 2
32 13 1 15 9 2 15 1 9 9 1 9 13 1 0 9 2 1 0 9 10 9 4 0 9 9 13 1 9 1 9 2 2
25 13 15 2 16 0 9 9 1 9 1 9 9 1 0 9 13 9 9 14 1 12 9 1 9 2
38 9 0 9 9 3 13 2 16 3 0 9 4 13 9 2 15 13 1 12 2 12 2 12 1 9 0 0 9 2 0 9 7 9 1 0 9 2 2
18 1 10 9 0 9 1 0 9 4 9 9 9 13 13 14 12 9 2
13 1 10 9 3 9 9 9 1 9 13 0 9 2
8 1 9 0 13 7 9 0 2
10 10 0 9 15 1 9 9 3 13 2
16 0 0 9 1 9 12 9 13 13 3 0 9 9 1 9 2
46 1 10 9 4 9 9 0 1 9 0 1 12 2 9 12 2 3 0 9 12 9 13 0 2 13 13 3 12 2 12 9 2 3 1 9 2 16 0 0 9 9 13 1 9 13 2
18 1 9 9 1 9 7 13 1 9 0 9 9 0 2 14 12 2 2
17 13 2 14 15 9 2 12 1 9 13 13 7 9 13 10 9 2
23 13 4 15 7 9 9 9 9 0 2 9 2 11 11 11 2 16 1 9 13 1 9 2
22 2 9 13 3 2 7 16 1 11 13 0 9 1 0 9 9 2 2 13 11 11 2
14 2 1 12 2 12 2 3 9 9 13 13 0 9 2
7 13 15 0 9 7 9 2
16 0 0 9 3 1 9 1 9 0 9 13 9 9 9 13 2
8 7 1 10 9 15 15 13 2
10 9 13 0 7 0 9 13 0 2 2
3 10 9 9
1 9
3 10 9 9
11 9 0 9 9 1 9 13 1 9 3 2
8 13 15 9 2 9 7 9 2
6 15 3 4 13 9 2
38 3 3 4 15 13 2 0 9 12 9 15 13 1 12 9 1 0 9 1 9 2 1 12 9 1 0 9 1 9 7 3 1 12 9 1 0 9 2
5 15 13 9 9 2
20 1 0 9 13 7 3 0 9 0 9 9 1 11 2 0 2 9 2 9 2
34 16 13 9 0 9 9 2 3 1 9 13 9 12 9 11 1 12 9 1 12 9 2 1 9 9 2 15 13 3 9 2 1 12 2
12 3 0 13 7 10 0 9 2 9 9 9 2
31 14 3 13 0 2 9 2 9 13 2 16 4 10 9 13 3 1 0 9 2 3 0 9 13 9 1 9 9 1 9 2
22 1 9 1 9 13 9 3 14 12 9 2 9 1 0 9 13 3 14 1 15 3 2
7 7 9 13 15 3 0 2
41 14 3 3 1 9 7 9 0 0 9 1 0 9 2 15 1 15 13 13 1 0 9 2 1 12 2 9 0 9 13 1 9 0 0 9 2 15 9 3 13 2
41 3 16 3 1 0 9 9 9 2 3 9 9 13 1 9 13 9 9 2 13 1 12 2 9 0 0 9 13 2 16 10 9 9 13 9 1 9 1 0 9 2
28 13 0 13 2 16 0 9 13 1 9 9 0 9 1 0 9 13 9 9 1 0 9 2 15 9 3 13 2
30 9 2 13 16 0 9 0 2 9 2 9 2 4 3 13 13 0 9 9 0 0 9 0 9 7 3 3 0 9 2
35 3 1 0 9 9 1 0 0 9 7 4 0 0 9 2 3 9 1 0 9 2 1 10 9 3 3 13 9 2 2 13 1 0 9 2
34 13 0 7 0 9 2 1 15 0 13 3 13 0 0 0 9 2 3 3 2 16 3 1 9 0 9 13 0 9 0 9 3 3 2
8 7 3 7 1 0 9 9 2
17 1 9 0 0 9 13 2 16 0 9 0 9 3 0 9 13 2
11 1 10 9 15 7 13 13 0 0 9 2
21 3 3 13 2 16 3 13 1 11 7 1 0 9 0 11 2 3 1 0 11 2
26 3 3 15 7 9 13 1 9 9 2 15 7 10 9 13 2 15 13 13 9 9 1 9 0 9 2
9 9 9 0 15 4 1 9 13 2
3 9 2 12
3 9 1 9
24 12 9 0 1 0 9 15 9 9 13 2 16 9 13 1 0 9 11 13 3 9 9 9 2
14 3 0 9 0 9 0 0 9 13 7 0 0 9 2
15 3 1 12 9 0 4 13 13 9 14 1 12 1 9 2
18 3 3 9 13 1 15 2 16 1 0 9 13 9 13 11 7 11 2
22 14 12 9 15 7 13 2 16 9 0 9 13 13 1 9 9 2 1 11 7 11 2
11 0 9 4 15 3 13 0 12 9 9 2
7 9 13 3 0 9 0 2
39 16 15 13 2 16 9 11 7 11 4 3 1 0 9 16 0 13 0 9 0 9 2 7 7 1 10 12 9 13 9 1 9 0 9 3 1 0 11 2
27 3 2 16 3 1 0 0 9 9 11 7 11 2 15 13 1 0 9 9 2 4 0 9 13 13 3 2
26 0 0 9 7 13 2 16 9 0 9 13 3 14 9 9 1 0 9 2 7 7 1 0 0 9 2
15 13 14 7 14 1 15 9 0 9 13 11 13 3 0 2
2 9 9
21 1 12 9 12 2 9 13 1 9 9 1 9 9 12 0 9 0 9 11 11 2
18 10 9 11 12 11 13 3 1 9 7 13 1 9 2 3 15 13 2
15 11 2 11 2 15 10 9 13 15 2 13 0 0 9 2
10 9 15 1 0 9 9 9 9 13 2
14 9 13 1 9 10 0 9 2 1 9 1 0 9 2
22 11 2 11 3 13 2 16 3 2 13 2 2 7 1 9 15 13 1 0 9 9 2
16 1 9 12 2 9 10 9 13 1 11 9 9 11 11 11 2
22 3 2 16 4 13 0 9 2 13 1 9 1 0 9 10 9 11 7 13 1 9 2
7 9 4 1 9 3 13 2
11 9 13 9 0 9 7 9 0 0 9 2
21 3 1 9 13 1 9 3 3 12 9 1 9 10 9 2 15 15 13 0 9 2
9 3 4 11 2 11 13 1 9 2
2 0 9
22 9 2 15 3 13 1 0 11 1 0 9 0 9 11 2 13 13 3 0 0 9 2
21 9 9 13 13 0 9 2 16 4 3 13 9 0 9 9 7 13 15 15 13 2
13 16 4 3 13 2 13 15 1 15 0 0 9 2
9 9 0 9 1 11 13 10 9 2
42 1 0 9 1 0 9 1 0 9 2 0 0 9 9 2 15 9 0 9 13 1 10 9 1 0 0 9 7 0 9 14 1 9 1 9 2 3 2 0 9 2 2
11 3 15 3 3 0 9 13 10 9 13 2
9 7 3 15 13 3 1 10 9 2
39 13 3 14 9 3 0 9 2 7 3 15 1 15 13 1 9 0 9 13 15 9 3 2 16 15 13 9 2 7 3 13 2 3 15 1 15 9 13 2
13 3 15 13 1 9 3 0 9 9 11 14 3 2
20 13 7 13 2 16 10 0 9 1 0 9 13 0 9 0 9 10 9 13 2
1 9
48 9 9 0 7 9 11 11 11 2 15 13 11 11 2 11 16 0 9 1 12 2 9 9 2 3 13 2 16 10 9 1 9 10 9 2 0 1 0 0 9 11 2 15 10 9 3 13 2
22 13 2 16 16 13 1 9 10 9 2 13 1 9 9 1 1 9 12 0 0 9 2
21 2 1 1 0 9 9 15 15 13 13 0 2 7 3 15 0 13 2 2 13 2
18 3 15 13 9 1 9 2 15 13 0 9 1 0 9 9 9 11 2
33 3 2 16 4 15 15 3 3 13 2 7 13 15 1 10 9 9 12 0 9 2 13 2 15 4 13 2 13 2 15 4 13 2
10 10 9 0 9 2 15 13 7 13 0
8 9 13 9 0 7 3 0 2
13 13 0 7 0 9 3 0 9 1 9 3 0 2
20 13 10 9 13 2 13 2 7 1 15 13 2 3 7 9 13 1 10 9 2
19 13 7 9 0 3 1 10 9 2 9 2 9 2 9 2 9 2 2 2
14 1 0 9 4 13 16 15 0 2 3 7 3 0 2
46 1 0 9 13 15 13 9 2 7 16 13 1 0 0 9 2 14 1 9 9 11 11 0 3 13 2 16 4 15 9 7 9 13 2 16 16 4 3 3 13 2 13 16 2 15 2
6 11 11 13 0 9 2
22 13 7 9 2 16 3 15 15 13 2 13 2 0 9 0 9 2 0 15 0 9 2
25 1 0 9 7 2 13 0 9 0 11 2 15 13 12 9 9 2 0 3 3 2 3 13 0 2
37 13 1 9 1 0 9 9 2 3 1 0 9 2 0 2 3 0 9 2 9 7 9 15 13 13 9 2 9 0 0 9 3 16 0 0 9 2
24 11 2 1 0 7 9 0 9 9 0 2 13 9 0 9 2 9 2 7 7 0 0 9 2
28 7 10 9 9 13 3 1 9 2 1 0 9 1 0 9 2 1 9 7 9 2 15 13 7 15 15 13 2
25 13 1 9 2 1 15 15 7 9 13 3 0 9 2 7 13 15 2 15 3 13 7 13 9 2
37 3 13 3 3 2 16 4 9 13 1 15 2 16 3 10 9 3 1 11 2 9 2 11 7 11 13 2 3 13 13 1 9 9 9 2 9 2
35 13 15 15 3 3 2 3 1 9 7 9 9 13 3 9 15 2 3 3 15 9 13 15 2 16 13 2 7 3 13 2 2 3 13 2
7 11 11 13 14 9 0 2
12 3 15 9 0 2 9 2 13 9 0 9 2
17 13 15 9 1 9 0 9 7 1 10 0 2 7 0 2 9 2
25 9 0 9 0 9 0 0 0 9 15 13 1 0 0 0 9 1 9 12 2 2 12 2 9 2
41 1 9 2 1 12 9 2 13 3 2 0 9 9 11 2 11 0 9 2 0 11 7 9 1 11 7 9 9 11 2 11 12 9 2 10 9 15 9 3 13 2
23 1 0 9 1 11 13 1 9 14 1 12 2 9 1 11 9 12 2 9 0 0 9 2
35 1 9 0 2 11 15 13 9 1 11 2 11 2 11 2 11 7 11 2 15 13 9 11 2 11 2 11 2 11 2 11 7 0 9 2
31 9 9 1 9 2 0 1 12 2 9 9 11 2 11 2 11 2 13 1 0 0 9 1 0 9 13 1 12 2 9 2
26 0 9 0 9 2 0 9 11 11 13 1 10 9 12 2 9 1 12 9 2 1 0 9 0 9 2
2 0 9
51 1 10 9 1 9 7 9 2 1 11 2 11 7 0 9 2 15 15 3 3 1 10 9 13 2 7 1 15 3 2 13 1 0 9 2 2 1 2 9 2 3 1 9 13 9 7 9 2 2 2 2
14 1 15 15 13 9 2 1 15 3 13 7 13 0 2
31 13 9 2 9 1 9 0 9 2 3 1 9 11 11 2 13 9 12 1 0 0 9 0 9 7 0 9 2 11 11 2
46 9 14 2 16 9 2 15 7 3 13 1 9 2 1 15 11 13 1 0 9 2 1 9 11 11 2 7 1 10 9 1 11 11 2 0 7 3 0 9 2 2 13 3 9 0 2
19 15 3 13 9 9 0 7 13 3 0 9 10 0 0 9 7 0 9 2
12 0 3 0 0 9 13 7 7 3 3 0 2
13 3 13 9 1 0 9 1 9 10 9 7 9 2
19 1 9 1 0 11 3 1 11 9 4 9 13 9 9 11 12 0 9 2
3 13 15 2
28 9 2 11 11 2 0 9 2 0 0 9 9 3 3 0 2 0 9 0 7 0 9 2 13 1 0 9 2
44 9 2 11 11 2 9 13 9 2 0 9 0 9 1 10 0 2 0 9 2 1 9 9 2 1 15 15 13 2 9 1 0 9 2 2 3 1 12 1 9 9 12 2 2
27 9 2 11 11 2 0 9 2 11 11 1 0 9 0 0 9 2 1 15 13 1 0 9 9 0 9 2
8 1 9 1 10 9 9 11 2
4 1 9 2 3
13 9 9 0 9 11 11 3 13 9 9 10 9 2
18 13 15 13 3 1 9 0 9 7 1 0 9 2 15 13 9 3 2
17 13 15 7 13 0 9 2 7 4 9 13 13 0 1 0 9 2
10 9 9 4 3 13 13 1 9 9 2
11 1 9 15 13 9 13 9 0 0 9 2
5 13 13 0 9 2
10 15 9 4 13 4 13 1 0 9 2
8 13 4 7 4 3 3 13 2
11 3 4 15 13 13 9 9 3 0 9 2
24 15 15 13 0 9 2 11 11 13 9 1 9 10 0 9 13 1 0 9 9 9 7 9 2
22 13 1 9 2 7 16 13 9 2 3 13 2 1 9 0 9 2 0 9 13 9 2
28 9 4 15 13 13 14 1 0 9 2 7 7 1 0 9 11 11 2 15 13 9 1 0 9 13 0 9 2
14 15 13 13 0 9 2 7 13 13 9 9 0 9 2
11 13 13 7 0 7 0 9 1 0 9 2
3 12 9 3
14 9 2 9 7 9 11 11 1 9 9 1 0 0 9
3 0 9 2
60 3 15 13 12 1 9 9 9 2 9 0 9 7 9 3 2 9 3 2 9 7 9 0 9 9 13 15 1 9 2 9 0 0 9 2 3 3 0 11 1 0 9 11 11 10 11 15 13 2 3 2 3 15 13 3 16 12 9 3 2
32 2 3 2 13 9 0 9 1 9 11 2 13 15 9 1 0 9 2 7 3 15 1 0 9 13 2 16 13 9 0 9 2
13 16 13 9 2 13 15 1 9 10 0 11 2 2
21 12 9 3 2 16 13 2 13 1 9 11 11 9 1 9 9 1 0 0 9 2
14 2 14 2 0 0 9 15 13 2 3 3 15 13 2
19 16 9 13 0 0 9 2 13 4 1 12 0 9 2 7 3 15 13 2
14 14 2 13 3 2 13 1 3 0 9 2 3 9 2
17 3 4 7 13 0 9 7 2 9 2 12 9 9 2 2 2 2
3 15 13 2
11 0 9 15 7 13 2 1 15 15 13 2
31 2 13 4 15 0 9 2 2 9 1 15 2 16 15 13 13 7 1 0 9 2 2 7 15 4 13 2 7 7 13 2
17 9 13 15 1 9 13 1 9 2 15 15 13 13 0 2 0 2
6 13 15 1 9 9 2
33 9 9 9 1 0 0 9 15 13 13 1 9 0 9 7 9 2 7 0 9 2 0 9 2 15 13 13 3 7 3 1 9 2
14 3 3 9 13 1 9 0 0 9 7 13 1 9 2
6 9 13 9 1 9 2
14 1 15 13 0 2 16 4 13 10 9 10 0 9 2
22 2 7 2 13 3 1 9 2 16 9 7 9 10 9 2 3 2 13 1 9 2 2
4 2 3 13 2
20 10 9 13 2 16 3 13 3 2 1 9 13 9 2 16 13 3 3 3 2
24 7 16 4 13 0 2 1 9 4 12 0 9 13 9 1 9 2 9 2 12 2 2 9 2
35 1 10 9 4 13 7 1 9 2 7 1 9 2 3 2 16 15 1 11 13 7 15 13 2 16 3 13 3 3 2 13 1 15 9 2
31 2 0 9 10 9 13 1 12 9 2 12 13 9 9 2 1 0 9 2 0 9 7 0 9 13 15 3 15 12 9 2
5 15 15 13 13 2
6 9 2 9 2 9 2
11 2 13 2 15 15 15 13 15 2 2 2
40 9 2 9 2 9 2 9 1 9 2 0 9 7 3 0 9 1 9 9 2 16 15 13 2 1 9 0 11 11 2 11 11 2 0 9 0 9 2 2 2
6 2 13 9 2 2 2
11 13 4 15 1 9 9 13 9 0 9 2
13 2 7 2 9 13 10 0 9 1 9 9 9 2
6 13 4 15 3 0 2
9 9 15 1 15 13 13 0 9 2
15 0 9 2 3 15 3 13 2 13 2 16 4 13 13 2
9 9 3 13 12 9 7 13 15 2
9 1 9 3 15 7 9 13 9 2
4 13 15 15 2
9 14 13 9 1 2 0 9 2 2
28 13 4 7 0 9 7 13 4 3 0 9 1 9 11 2 1 15 4 13 3 0 9 2 0 9 7 9 2
32 13 2 16 1 9 9 1 0 0 9 15 13 15 2 7 7 15 13 2 9 15 9 2 1 9 10 9 2 13 15 2 2
2 11 11
3 9 2 9
10 9 13 11 11 2 9 9 0 9 2
41 2 3 3 15 1 0 9 13 0 9 1 9 7 0 9 2 15 13 0 9 1 9 1 0 11 2 15 13 0 9 1 12 9 3 12 0 9 1 0 9 2
15 13 15 3 1 0 7 0 9 7 1 9 13 0 9 2
20 13 2 16 13 0 13 10 9 2 1 15 13 7 9 0 9 2 10 9 2
38 3 13 3 3 0 9 2 7 3 11 9 1 11 2 9 2 15 13 1 15 0 3 1 9 7 9 2 7 0 11 1 9 0 9 11 11 2 2
4 9 9 1 9
5 11 2 11 2 2
35 0 0 9 2 15 13 1 11 13 13 1 12 2 9 0 9 2 4 13 4 2 16 9 3 13 9 0 9 2 3 1 10 9 13 2
29 1 0 9 0 9 9 4 13 9 0 9 2 1 15 15 0 9 0 9 2 9 7 9 0 7 0 4 13 2
16 3 4 13 2 1 0 9 2 1 9 9 9 3 0 9 2
21 13 15 13 7 9 2 15 13 1 9 13 1 0 9 3 0 9 1 0 9 2
13 9 9 9 0 9 13 4 13 1 0 0 9 2
9 9 4 13 1 9 9 0 9 2
9 0 9 0 9 11 2 11 2 2
18 0 9 0 0 9 1 11 15 3 13 11 9 2 0 9 10 9 2
12 9 13 0 0 9 3 1 0 9 0 9 2
23 2 1 9 9 13 3 0 9 15 9 0 0 0 9 2 2 13 11 9 1 10 9 2
3 9 0 9
8 13 4 7 13 9 1 0 9
35 1 0 9 2 3 1 9 13 9 1 9 3 0 12 0 7 12 0 9 2 15 13 1 15 2 16 1 0 9 4 13 9 3 9 2
16 9 1 0 9 13 1 15 3 3 0 2 7 7 0 2 2
13 1 9 1 9 1 0 9 13 9 7 10 9 2
21 3 1 9 1 11 2 11 13 3 9 1 0 0 9 12 9 0 9 1 9 2
7 7 3 13 3 0 9 2
7 1 9 13 9 7 9 2
19 9 1 9 9 1 10 9 3 7 13 3 0 2 3 15 9 9 13 2
23 0 9 1 9 9 0 9 1 9 1 11 13 0 9 14 1 9 2 3 13 9 9 2
17 1 11 11 2 9 9 2 4 15 13 9 7 10 9 3 13 2
12 0 9 1 0 9 13 7 0 9 1 11 2
5 2 11 2 11 2
10 9 0 9 13 4 7 13 9 1 0
35 1 0 9 2 3 1 9 13 9 1 9 3 0 12 0 7 12 0 9 2 15 13 1 15 2 16 1 0 9 4 13 9 3 9 2
26 2 0 9 15 13 13 9 1 9 7 1 0 9 2 2 13 15 9 11 11 1 12 2 0 9 2
17 2 10 9 7 13 3 7 9 2 15 13 1 9 9 1 9 2
16 9 1 0 9 13 1 15 3 3 0 2 7 7 0 2 2
13 1 9 1 9 1 0 9 13 9 7 10 9 2
22 2 0 9 13 1 9 9 7 9 1 15 13 9 1 0 9 2 2 13 11 11 2
19 3 1 12 0 9 13 3 7 12 0 9 7 12 9 1 9 0 9 2
19 1 9 11 15 9 1 9 3 13 7 9 2 15 15 1 9 13 13 2
15 12 3 0 9 13 3 1 9 12 2 0 9 0 9 2
35 1 0 9 9 9 3 3 9 13 0 0 9 2 9 2 0 9 1 0 9 2 9 13 1 0 9 9 7 13 15 1 12 0 9 2
23 9 1 9 13 13 9 9 2 7 3 1 0 9 15 3 3 1 10 9 4 13 0 2
13 0 12 13 12 2 0 9 13 1 9 9 9 2
21 3 1 9 1 11 2 11 13 3 9 1 9 12 9 0 9 1 0 0 9 2
4 0 9 13 9
5 11 2 11 2 2
17 0 0 0 9 13 1 11 3 1 9 7 13 13 1 9 9 2
11 9 1 0 11 7 3 13 14 12 9 2
18 2 9 1 0 0 9 2 15 13 13 10 0 9 2 13 3 0 2
29 9 2 3 4 13 12 9 2 13 0 2 2 13 15 1 9 3 0 9 1 9 0 9 0 11 11 11 11 2
3 11 3 13
21 0 9 0 9 7 9 11 11 11 13 3 1 9 0 9 9 2 9 7 9 2
30 0 11 12 2 15 13 1 11 1 9 9 11 2 13 1 12 9 1 12 2 9 9 9 12 3 11 1 0 9 2
21 2 13 0 13 9 9 1 9 9 2 2 13 3 9 11 11 1 0 0 9 2
11 9 7 1 10 9 13 13 14 0 9 2
21 1 9 13 1 3 0 0 9 2 3 13 1 9 13 9 1 12 9 1 9 2
13 1 0 9 13 9 0 11 9 1 9 9 9 2
21 1 10 9 13 13 1 9 0 9 9 3 1 9 2 3 12 9 1 9 9 2
21 0 9 11 11 7 11 11 2 15 13 13 1 0 9 2 4 13 9 1 9 2
10 2 9 1 9 13 1 0 9 3 2
14 9 0 9 1 9 13 13 2 2 13 15 11 11 2
14 0 1 9 13 3 0 9 2 1 10 9 13 9 2
7 1 11 3 13 7 9 2
40 16 1 9 9 0 9 9 1 11 4 11 11 1 9 0 13 1 9 7 10 0 9 13 3 0 2 1 9 9 1 0 9 1 11 15 10 9 3 13 2
20 9 13 1 9 0 9 9 2 11 2 11 3 0 2 16 9 13 13 9 2
16 2 9 11 1 15 3 1 9 13 2 3 7 13 1 9 2
15 1 0 9 15 13 0 0 9 2 3 9 1 0 9 2
12 9 3 13 1 9 2 2 13 15 9 11 2
17 9 13 13 1 0 9 1 9 7 1 0 9 9 1 0 9 2
18 9 1 9 1 0 9 13 1 0 9 0 9 11 11 1 11 13 2
8 2 13 9 9 9 2 12 2
28 0 0 11 2 1 15 15 1 9 3 3 3 13 11 11 2 4 1 9 9 13 1 0 9 9 1 11 2
9 9 13 1 9 9 7 0 9 2
2 9 13
2 11 2
16 9 9 1 11 7 11 1 9 11 2 9 15 3 13 13 2
15 13 13 7 13 9 1 9 9 12 1 9 11 2 11 2
22 1 9 12 2 9 2 3 9 13 2 15 1 10 9 13 10 9 0 9 7 9 2
15 9 4 13 9 1 9 1 12 9 7 9 14 12 9 2
13 1 9 11 7 11 9 13 1 12 9 0 9 2
1 9
4 13 1 9 2
15 9 13 1 9 12 0 9 1 11 1 9 11 2 9 2
17 13 7 0 9 2 16 3 4 13 1 0 9 9 1 0 9 2
3 0 9 2
21 9 1 9 9 9 13 9 2 15 15 3 0 9 13 1 0 9 9 1 11 2
8 13 15 3 3 9 0 9 2
3 3 13 2
11 9 2 3 13 1 11 3 2 3 9 2
19 9 1 9 12 7 12 9 2 9 2 1 9 12 7 12 9 2 9 2
20 1 11 3 7 3 2 0 9 12 7 12 2 0 12 7 12 9 2 9 2
16 9 13 1 9 1 12 2 12 7 13 1 12 2 12 9 2
16 9 13 1 9 1 12 2 12 2 13 1 12 2 12 9 2
19 9 9 2 0 9 12 9 2 9 1 9 12 2 0 12 1 9 12 2
9 0 0 9 13 12 9 2 9 2
12 0 9 2 0 9 13 0 2 0 9 0 2
5 0 9 2 11 2
1 9
2 0 9
9 1 9 13 3 0 0 9 9 2
12 1 9 1 15 3 7 3 2 1 0 9 2
16 15 13 0 9 1 9 0 9 2 13 9 9 16 0 9 2
8 1 9 0 9 3 13 9 2
10 15 13 13 3 13 0 9 1 9 2
13 1 0 9 9 9 13 7 13 15 15 4 13 2
23 16 15 11 13 4 13 11 2 13 15 2 16 9 13 1 9 10 0 9 9 2 13 2
12 9 3 4 13 9 1 10 0 9 7 9 2
31 0 7 13 2 16 0 9 1 9 2 1 15 4 13 2 7 3 7 1 9 2 15 4 13 2 13 13 9 0 9 2
14 13 15 3 2 16 1 0 9 13 3 3 0 9 2
28 1 9 0 0 9 15 3 4 3 0 9 0 9 11 11 13 13 0 7 0 0 9 2 15 13 3 13 2
3 11 13 9
5 11 2 9 9 13
2 11 2
34 2 13 1 15 0 2 16 4 11 0 3 13 0 9 2 2 13 11 3 3 1 9 11 1 9 1 11 1 9 1 0 0 9 2
28 1 10 9 13 1 9 2 15 9 13 0 2 9 2 13 15 9 9 1 0 9 7 4 13 1 0 9 2
29 2 13 9 0 9 3 0 1 9 11 13 3 0 2 2 13 1 0 9 1 9 0 9 11 11 2 11 2 2
8 2 3 15 3 13 0 9 2
37 13 4 15 1 9 2 16 4 4 13 0 9 2 15 13 1 9 0 0 9 2 2 13 7 13 2 2 14 15 2 15 13 0 2 13 0 2
11 15 13 13 3 1 0 11 1 9 2 2
16 10 10 9 3 1 9 13 1 0 9 11 11 2 11 2 2
19 2 7 0 9 0 11 13 3 9 1 0 9 16 9 11 2 2 13 2
33 15 3 10 9 13 9 2 2 13 4 15 13 2 16 9 9 13 12 2 12 2 12 2 7 7 3 15 9 0 11 13 2 2
2 0 9
3 9 9 9
8 11 1 11 1 0 9 1 11
20 15 14 13 10 0 9 11 11 2 3 2 2 11 11 1 0 0 9 11 2
10 9 11 2 11 9 9 9 1 12 9
36 0 9 1 9 1 12 9 11 11 13 1 11 2 16 13 13 15 13 1 9 0 9 1 10 9 11 11 1 0 9 12 2 9 1 11 2
16 10 9 13 0 9 0 9 9 2 15 13 3 12 12 9 2
13 2 13 0 9 2 7 13 3 3 13 10 9 2
25 15 1 15 13 2 16 13 0 9 2 7 16 13 9 2 9 2 11 3 13 2 3 13 2 2
19 12 9 4 13 1 0 9 9 2 12 7 13 1 0 9 13 9 9 2
22 11 1 9 1 11 3 3 3 13 11 11 2 11 1 11 13 0 1 10 9 11 2
8 11 3 13 0 9 9 0 9
22 1 9 3 15 1 9 9 11 13 9 1 9 0 9 7 13 1 15 9 0 11 2
40 0 9 4 13 1 9 11 9 1 0 0 0 9 2 2 9 9 11 1 9 13 0 1 1 10 0 9 2 15 15 13 0 0 9 1 0 9 9 2 2
14 0 13 2 16 1 0 9 15 9 13 3 1 11 2
17 7 10 9 2 1 15 15 0 9 1 9 1 9 0 3 13 2
23 1 9 9 15 15 13 11 1 11 7 9 10 9 13 12 0 2 12 0 7 12 0 2
9 9 11 9 2 11 3 1 12 2
23 2 1 9 15 1 15 13 9 11 2 13 14 14 1 0 0 9 2 15 9 3 13 2
14 3 3 11 3 13 2 15 3 4 1 15 3 13 2
30 13 4 0 2 16 4 15 1 15 13 10 9 2 13 13 2 16 15 3 13 2 16 15 1 11 13 1 10 9 2
49 2 0 0 9 3 9 13 2 7 0 9 4 3 13 1 9 2 16 1 3 0 9 13 1 0 9 2 0 9 1 0 0 9 11 2 2 15 13 9 0 7 15 15 13 10 9 1 9 2
2 9 3
21 9 9 0 9 11 11 1 0 0 9 1 11 13 3 0 9 1 9 12 9 2
8 9 9 13 3 0 12 9 2
11 9 15 13 13 1 11 11 1 11 11 2
4 11 13 0 9
8 9 11 3 1 12 2 9 11
4 11 13 0 9
8 1 0 9 1 11 13 3 3
19 0 12 9 13 13 1 0 0 9 2 7 3 13 13 1 0 7 0 2
28 15 3 2 16 1 0 9 13 9 0 9 2 13 15 1 12 2 0 9 2 16 15 13 2 16 3 13 2
26 1 10 9 13 0 9 1 11 2 9 1 0 9 2 15 3 1 0 9 13 14 1 12 2 9 2
19 3 13 3 1 9 2 0 1 0 9 7 1 0 9 0 9 2 12 2
33 1 15 9 9 2 11 2 2 10 9 3 13 16 9 2 11 1 11 2 11 1 11 7 11 1 11 11 13 1 12 9 12 2
23 13 4 15 7 12 2 7 13 2 16 15 9 11 1 11 7 9 11 1 11 3 13 2
30 3 13 0 9 11 2 13 0 9 2 7 1 9 12 2 12 1 15 13 12 0 9 2 9 7 3 9 0 11 2
7 7 3 12 2 12 2 2
9 3 3 13 1 9 3 1 11 2
32 11 15 13 1 0 9 7 1 0 9 1 0 9 2 1 0 11 13 3 10 9 16 3 2 7 13 15 9 12 2 12 2
29 9 13 9 11 2 2 13 9 11 15 13 2 3 4 15 13 1 9 12 2 12 7 3 1 9 12 2 12 2
17 7 3 1 9 13 13 2 16 9 13 0 9 1 3 0 9 2
6 3 4 15 13 15 2
23 3 1 9 15 9 13 9 2 1 9 15 4 13 11 2 1 0 9 13 0 9 9 2
15 7 1 12 9 13 0 9 9 2 1 9 1 9 2 2
13 3 15 13 7 0 9 11 1 0 9 1 11 2
11 2 13 15 9 2 3 1 9 4 13 2
20 14 15 10 9 13 9 2 16 13 1 9 9 16 9 2 7 3 3 13 2
17 3 13 9 2 3 13 11 9 2 7 9 15 1 0 9 13 2
3 13 0 2
17 14 1 9 4 13 9 2 7 3 15 13 11 0 0 9 2 2
17 12 9 12 2 9 13 0 9 2 11 1 11 7 11 1 11 2
27 9 13 9 9 9 11 11 2 2 13 1 9 1 9 9 11 2 16 4 15 0 13 3 3 1 9 2
14 16 13 9 2 13 0 9 1 0 9 7 9 9 2
19 3 3 13 11 11 2 11 2 11 2 11 7 11 9 2 11 0 9 2
16 3 1 9 0 1 10 9 2 3 1 9 0 1 12 9 2
11 16 4 15 15 13 2 16 13 13 2 2
7 3 1 11 2 11 2 11
9 9 1 0 4 10 9 13 15 12
26 3 12 1 0 12 0 9 1 0 9 4 13 1 11 1 11 2 1 12 9 2 12 2 9 12 2
34 13 10 0 9 2 16 10 9 4 15 10 0 9 3 13 13 2 13 4 3 12 2 12 7 1 9 3 0 9 15 13 12 9 2
29 3 2 1 9 0 11 7 11 2 1 0 9 9 7 9 14 9 1 9 2 13 9 11 13 1 0 12 12 2
27 1 15 3 13 3 9 15 9 2 15 13 9 11 13 1 10 0 9 1 9 1 0 9 12 1 11 2
28 1 3 0 0 9 15 3 3 1 0 9 13 11 2 15 3 13 0 9 7 0 9 15 2 13 2 3 2
26 1 9 0 9 7 9 13 0 2 16 0 9 1 11 13 13 13 2 1 15 13 0 9 7 9 2
18 0 9 13 0 2 3 13 9 15 0 2 16 9 13 1 9 9 2
23 9 11 2 2 16 4 13 13 0 9 1 11 1 0 9 2 15 4 14 3 13 13 2
20 14 2 14 2 11 13 1 15 2 13 2 16 1 11 15 9 13 3 3 2
11 13 15 0 0 9 2 15 15 7 13 2
16 11 13 0 9 2 7 3 1 9 2 7 15 15 13 2 2
36 1 0 9 13 10 9 3 15 2 16 2 0 9 9 7 9 11 4 13 3 2 7 14 3 2 16 4 1 15 10 9 13 3 3 2 2
10 3 7 3 11 9 1 0 9 13 2
14 3 15 7 13 13 9 2 16 9 9 13 3 11 2
13 2 16 13 2 3 3 1 9 9 2 2 2 2
36 1 9 0 0 9 10 9 3 13 13 2 13 15 15 3 14 3 0 2 2 13 13 1 15 2 16 11 13 1 9 2 15 9 11 13 2
34 7 16 1 0 9 15 0 13 2 16 13 1 9 2 3 3 7 13 0 9 11 7 1 11 7 1 10 9 13 11 7 11 2 2
23 1 9 4 3 1 12 9 13 12 9 1 0 9 2 1 12 3 15 0 1 0 9 2
22 1 0 9 9 13 3 0 9 9 1 0 9 2 15 1 0 9 9 13 13 9 2
38 9 9 13 13 1 12 2 13 15 0 9 11 2 15 15 13 1 9 12 9 9 1 9 1 11 1 11 2 13 4 12 2 12 9 1 9 2 2
40 1 9 13 9 9 0 9 1 9 10 7 0 3 0 9 1 11 2 11 7 11 2 9 15 3 13 1 0 9 11 2 1 9 9 1 0 9 13 11 2
3 0 0 9
26 12 9 1 0 0 9 11 2 11 4 1 0 9 9 13 0 9 1 11 7 0 9 11 11 11 2
37 9 9 0 9 9 2 11 11 7 0 9 0 2 9 2 11 11 4 13 2 16 0 2 9 1 9 9 2 3 9 7 9 2 13 0 9 2
55 9 9 13 3 2 3 1 9 2 7 1 9 9 14 1 9 9 12 2 0 0 9 2 1 15 1 0 9 12 9 11 7 0 12 0 11 2 3 13 0 0 9 0 9 2 15 13 3 0 0 9 2 9 3 2
22 9 13 0 1 9 0 0 9 2 7 13 0 2 16 10 9 13 12 9 1 9 2
3 11 1 9
9 0 9 11 11 13 3 1 9 2
24 1 9 1 11 13 1 10 9 9 0 9 11 2 15 13 1 9 0 9 1 12 9 9 2
31 11 13 9 9 11 9 7 0 9 15 13 1 9 7 0 9 11 2 15 13 1 9 9 7 9 9 1 9 0 9 2
16 2 9 13 3 1 9 11 2 2 13 11 2 9 9 11 2
4 9 13 1 11
7 11 2 1 10 9 2 2
32 1 3 0 9 0 9 7 9 2 0 1 0 9 10 9 2 13 1 9 3 1 0 9 9 0 9 11 2 11 2 11 2
52 11 11 11 1 0 9 11 11 12 15 16 0 13 1 9 0 9 2 7 1 0 0 9 0 1 11 1 9 1 11 2 7 3 1 0 9 13 1 9 12 9 0 0 9 0 1 11 7 11 1 11 2
45 1 11 13 12 0 9 2 1 15 3 3 16 9 0 9 7 9 2 1 15 12 0 11 12 2 2 9 2 9 11 2 11 2 9 7 2 9 2 9 11 2 11 2 11 2
50 1 12 9 0 9 2 15 15 13 0 9 1 12 3 2 0 9 13 9 0 1 12 2 2 4 13 12 0 11 12 12 5 12 2 1 15 15 0 9 13 3 0 9 2 15 13 11 11 11 2
87 3 1 9 13 11 11 9 15 2 15 1 0 11 2 7 3 1 11 7 12 0 9 11 2 13 1 9 7 13 9 0 0 9 2 3 16 0 9 2 15 1 0 9 3 13 9 9 1 15 2 16 4 0 13 14 13 1 11 1 9 0 2 7 0 2 0 0 9 2 7 7 13 12 2 9 3 1 11 1 9 2 3 1 0 0 9 2
38 11 13 7 3 3 3 2 3 0 9 13 11 2 3 13 1 9 1 9 0 9 2 1 9 3 2 7 1 0 12 9 3 2 13 0 9 11 2
5 11 1 11 1 9
36 1 0 9 9 1 9 9 1 0 9 1 0 11 13 0 2 9 11 11 7 11 11 1 0 9 11 2 11 12 2 12 7 13 1 9 2
3 13 0 9
6 9 9 13 10 9 11
33 1 12 7 12 9 1 11 4 13 1 10 9 1 0 11 2 13 11 11 2 0 9 0 9 10 9 3 1 0 9 1 11 2
35 13 3 3 16 9 11 11 0 2 9 0 0 2 9 1 9 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 7 11 2
30 11 13 2 16 4 13 13 3 9 2 15 13 0 7 0 9 2 7 2 3 13 2 2 1 11 13 3 9 2 2
13 0 9 13 2 16 4 13 0 13 0 2 9 2
26 11 13 0 9 2 7 16 4 4 13 1 10 0 2 0 9 2 2 13 4 15 0 7 1 11 2
39 9 1 9 11 7 13 1 0 2 16 11 13 13 1 0 9 2 7 1 0 9 15 13 9 0 9 2 16 4 4 13 9 1 0 9 1 0 9 2
12 2 15 4 7 13 9 3 2 2 13 11 2
37 1 9 15 13 0 9 1 0 9 1 0 2 9 2 9 11 2 13 11 1 9 2 2 13 9 2 16 13 15 1 11 7 15 1 11 2 2
25 1 0 9 4 13 0 9 11 2 12 0 11 11 2 3 0 1 0 9 9 1 9 11 11 2
16 13 9 1 12 9 7 1 11 7 13 1 9 9 9 11 2
18 3 4 13 10 9 2 7 1 0 9 0 9 15 13 2 16 13 2
3 9 11 13
12 9 0 0 2 9 11 11 15 13 10 9 2
24 12 0 0 2 9 11 11 7 11 9 15 13 0 9 9 9 1 11 1 9 0 9 9 2
12 1 0 9 10 9 13 11 9 1 0 9 2
56 0 9 1 9 1 0 0 9 1 0 9 11 11 13 0 9 2 13 9 9 9 1 9 9 11 7 11 7 11 4 13 9 16 0 3 0 9 1 9 9 12 9 11 2 16 13 1 0 9 1 0 11 1 9 9 2
27 9 3 13 1 9 2 16 1 0 9 11 2 15 13 0 9 2 13 9 0 2 9 10 9 1 9 2
26 2 13 15 0 0 9 2 2 13 9 0 2 9 11 1 0 9 1 11 2 7 9 10 9 13 2
15 2 13 3 1 11 2 11 2 11 2 9 2 12 2 2
2 11 13
25 0 0 9 11 13 2 16 13 13 9 0 9 11 11 11 1 0 9 0 9 9 11 11 11 2
22 11 4 13 9 9 1 0 12 9 0 9 1 15 2 16 9 9 13 1 11 13 2
28 11 3 13 1 9 1 0 9 1 11 11 2 1 15 13 1 0 9 12 9 2 7 3 4 9 11 13 2
9 0 9 1 11 9 0 11 13 2
2 1 9
2 11 2
17 11 13 1 12 9 2 1 0 9 13 11 7 0 0 11 9 2
3 11 11 2
24 1 9 1 0 9 1 0 11 13 0 2 9 11 0 9 9 12 9 1 0 11 1 11 2
17 9 0 9 11 1 9 1 11 13 0 9 1 11 12 2 12 2
30 0 0 9 1 9 11 11 1 11 15 13 9 0 0 0 9 2 10 9 13 13 9 9 1 9 12 1 0 9 2
18 0 9 0 11 1 11 13 11 11 1 0 9 11 2 11 7 11 2
7 11 15 13 9 1 0 9
29 11 11 2 15 1 11 13 1 11 2 15 3 4 1 10 0 9 13 1 12 9 2 15 15 3 11 11 13 2
29 9 9 13 2 16 11 1 9 10 9 13 9 7 13 3 1 9 1 9 2 15 3 13 3 9 2 15 13 2
12 11 11 13 0 9 1 0 0 9 11 11 2
19 9 2 15 1 9 0 9 13 1 11 11 2 13 13 1 9 0 9 2
15 0 9 0 0 11 11 15 13 12 0 9 11 11 11 2
11 0 9 13 1 0 9 0 12 9 9 2
27 9 9 1 11 1 11 2 15 13 12 9 7 10 9 1 9 2 13 1 3 0 9 9 1 0 9 2
13 9 13 0 2 12 9 13 7 0 12 13 9 2
23 0 9 9 13 1 9 9 9 1 11 11 2 11 2 15 15 13 12 2 9 1 11 2
19 0 0 9 13 9 1 12 9 2 3 9 2 11 2 15 13 3 12 2
3 9 1 9
13 9 9 1 9 9 7 0 9 13 1 0 11 2
26 0 9 11 7 11 15 13 1 9 12 2 12 1 0 9 11 2 11 1 9 2 3 13 1 11 2
23 0 9 9 1 0 9 9 1 12 9 15 13 11 11 2 16 13 1 0 9 11 11 2
4 9 13 11 2
23 11 11 13 1 9 12 5 12 9 1 0 9 2 16 0 13 11 11 7 0 11 11 2
6 11 7 11 2 0 9
5 15 15 1 15 13
6 11 7 11 2 0 9
20 1 0 9 13 1 0 9 7 0 9 0 9 0 9 2 11 2 11 11 2
18 9 1 10 0 9 0 9 13 9 2 7 3 13 2 1 9 9 2
15 7 7 1 11 15 0 9 13 13 9 1 11 7 11 2
10 3 13 7 7 1 9 0 7 0 2
44 2 9 3 13 3 1 9 2 2 13 15 9 11 2 2 3 1 0 9 13 14 3 3 9 1 11 2 3 13 9 3 9 1 9 2 11 13 9 3 1 0 9 2 2
22 11 11 15 13 15 2 16 0 9 11 2 1 9 11 2 4 15 13 3 0 9 2
24 2 3 0 9 2 16 13 15 7 15 2 3 3 13 12 0 9 0 9 1 0 12 2 2
26 13 3 14 1 15 14 10 0 9 2 15 4 15 9 7 9 9 12 0 9 1 3 0 11 13 2
21 15 13 3 3 3 13 2 13 0 7 0 9 2 0 13 1 9 3 1 9 2
14 13 3 3 0 13 1 0 9 9 9 1 10 9 2
30 3 7 0 0 9 2 1 10 0 9 3 7 1 9 1 11 0 1 9 9 11 2 13 0 13 2 15 13 3 2
5 9 7 9 1 11
29 9 9 7 9 9 4 1 9 1 9 13 1 0 9 1 0 0 9 10 9 1 15 2 9 11 11 2 12 2
20 1 12 9 2 0 1 9 9 2 4 15 13 13 12 9 0 0 0 9 2
28 7 1 15 7 0 2 9 2 1 9 12 11 11 7 11 9 2 1 9 12 11 11 2 15 1 11 2 2
27 1 9 4 13 10 0 9 2 15 3 3 13 9 1 0 9 7 9 10 9 1 9 4 13 3 0 2
22 9 9 11 13 3 9 9 2 15 15 4 13 1 0 9 9 7 1 9 11 11 2
26 13 7 3 0 0 9 11 11 2 15 15 1 9 13 0 9 7 10 9 14 13 1 9 3 3 2
2 0 9
33 1 9 0 9 0 0 13 3 0 0 9 1 0 9 1 9 10 9 3 2 3 4 15 13 1 0 9 11 11 1 11 11 2
4 11 7 11 2
4 11 7 11 2
4 0 9 9 0
2 11 2
30 9 11 7 9 12 9 9 3 13 9 1 9 0 9 9 9 7 9 9 2 15 4 15 13 13 0 0 9 11 2
20 9 13 10 9 0 9 11 2 11 2 11 2 11 2 11 2 11 7 11 2
26 9 12 9 15 3 1 9 3 13 2 13 7 2 16 4 9 13 13 3 2 7 15 3 0 9 2
1 3
3 9 13 11
19 0 9 1 11 4 1 10 0 9 13 3 12 9 2 9 13 3 12 2
24 1 0 9 13 12 9 2 1 0 0 9 7 9 12 9 7 12 0 9 13 0 0 9 2
38 9 0 9 16 9 3 0 3 13 1 12 9 9 11 2 9 3 3 13 0 9 13 12 9 10 9 2 13 15 1 0 9 9 1 9 0 9 2
2 0 9
38 9 1 11 11 7 11 11 15 13 9 11 11 9 2 16 4 13 2 16 4 9 0 0 9 13 0 1 11 13 0 9 11 11 1 9 9 11 2
20 16 13 1 0 0 9 2 9 12 9 0 9 13 9 11 11 1 9 9 2
29 9 0 0 9 1 9 1 11 13 9 11 1 2 0 2 7 1 9 1 0 0 9 13 2 9 0 9 2 2
28 1 0 9 11 1 0 9 11 9 13 2 16 13 10 9 11 2 7 7 15 15 2 3 13 1 9 2 2
3 2 11 2
32 9 0 9 11 11 11 13 11 1 0 9 2 7 1 0 9 1 9 1 0 9 0 9 2 13 3 0 9 11 11 11 2
24 9 11 2 7 7 0 9 1 9 0 9 11 13 1 10 9 11 11 2 1 0 9 2 2
12 13 1 9 2 10 9 13 1 0 9 11 2
41 9 9 11 2 11 1 9 3 0 9 11 13 1 15 0 2 7 13 2 1 10 10 9 13 2 13 3 1 11 9 2 9 11 11 11 2 11 2 11 2 2
29 13 15 1 9 2 16 1 12 9 11 1 11 13 12 0 2 12 9 0 0 9 7 12 13 1 0 9 9 2
3 2 11 2
7 15 2 9 0 2 2 2
4 0 9 1 11
2 11 2
10 9 1 9 9 11 1 11 3 13 2
37 9 13 9 0 9 2 1 15 13 1 9 9 9 9 2 15 2 9 0 2 2 2 2 1 0 9 2 15 2 9 0 9 2 2 2 2 2
15 13 3 9 9 1 15 2 16 0 9 13 0 9 11 2
12 1 0 9 13 9 2 16 9 13 0 9 2
17 3 9 13 9 2 1 15 4 9 9 13 4 13 14 0 9 2
18 1 9 9 13 9 2 16 9 9 13 0 1 0 9 13 9 11 2
10 1 9 9 10 9 9 1 9 13 2
25 1 0 9 13 11 11 2 11 2 2 16 13 0 7 0 9 0 9 9 11 1 0 9 9 2
30 2 13 9 0 9 3 0 1 9 11 13 3 0 2 2 13 7 13 2 16 2 9 9 13 12 2 9 12 2 2
25 9 11 11 2 9 2 13 2 16 9 16 15 13 13 9 9 2 15 13 1 9 10 0 9 2
20 2 13 15 2 16 4 13 12 9 2 2 13 10 9 11 11 2 11 2 2
23 9 9 0 9 1 9 7 10 9 1 9 13 1 10 9 7 9 11 11 2 11 2 2
19 13 2 16 2 16 15 13 13 1 11 2 13 0 15 13 0 9 2 2
12 10 9 13 0 9 9 1 9 11 7 11 2
7 15 2 9 0 2 2 2
34 0 9 11 11 1 10 9 1 9 9 13 9 0 9 7 9 2 16 13 9 1 11 7 11 7 13 15 1 9 0 9 1 11 2
30 3 3 13 2 13 15 9 11 11 11 2 1 15 10 9 13 2 16 3 13 9 2 16 4 11 13 0 9 11 2
18 2 1 11 13 15 15 0 1 9 7 9 2 2 13 11 2 11 2
35 13 3 9 9 1 0 9 7 0 9 1 9 1 0 9 7 13 2 2 10 9 2 15 13 11 1 11 2 13 15 13 11 3 2 2
22 9 11 11 2 11 2 13 3 9 11 2 11 16 2 0 7 0 2 7 13 15 2
23 2 15 13 9 2 16 15 15 13 2 13 15 15 2 9 9 2 2 13 11 2 11 2
20 11 2 11 13 1 0 2 16 4 9 11 13 9 9 10 9 7 14 3 2
23 9 11 15 1 15 12 9 13 10 9 7 9 2 7 13 15 3 9 0 9 1 15 2
25 13 9 2 16 3 1 9 9 4 1 11 13 9 9 9 1 0 9 7 9 1 11 7 11 2
10 9 0 9 13 4 3 13 1 9 2
3 0 9 11
2 11 2
30 1 9 9 11 13 3 10 9 11 0 9 2 11 11 9 0 0 0 9 2 11 2 1 9 1 12 2 9 12 2
18 9 2 11 11 2 13 12 2 1 9 12 7 12 13 0 9 11 2
28 1 12 2 9 14 1 9 12 13 9 9 0 9 9 11 11 7 1 9 12 13 9 0 9 11 1 11 2
28 1 9 12 7 12 13 9 0 9 11 1 0 11 7 1 9 12 15 13 9 0 9 0 9 11 1 11 2
3 13 9 9
5 9 1 9 2 12
41 0 0 9 2 12 0 7 12 0 9 2 12 0 9 2 12 0 9 7 12 0 9 2 4 13 1 12 9 9 7 1 12 2 9 12 15 15 9 13 13 2
24 13 15 10 0 9 2 7 2 3 15 3 13 9 11 2 13 15 7 1 0 9 1 9 2
13 13 15 3 0 9 2 9 0 13 1 9 3 2
20 0 9 2 3 2 9 9 12 7 9 11 2 12 2 1 0 9 13 4 2
18 1 0 11 15 1 9 13 10 9 12 7 1 0 9 3 12 9 2
11 9 1 9 7 9 0 9 13 12 9 2
24 9 9 0 2 9 9 11 11 13 3 13 1 15 2 1 15 9 0 9 0 2 9 13 2
34 4 13 1 9 2 1 15 15 13 13 0 9 1 0 9 2 7 7 1 15 2 16 15 13 9 2 3 2 1 0 9 7 9 2
23 1 0 0 0 9 3 13 0 9 1 9 0 0 0 9 2 15 13 0 13 1 9 2
13 12 10 9 4 1 9 13 1 0 9 1 11 2
6 0 9 2 13 9 11
5 11 2 11 2 2
20 3 3 4 15 13 3 1 9 0 9 11 2 13 13 9 0 15 10 9 2
8 11 11 7 1 15 13 13 2
28 3 2 1 10 9 1 9 0 2 9 11 9 11 13 2 16 10 0 9 15 4 0 9 13 1 0 9 2
12 13 2 16 13 9 1 10 0 9 1 9 2
25 2 4 15 3 13 7 13 7 15 2 7 9 0 9 0 9 10 0 9 2 2 13 11 11 2
42 3 13 2 16 10 9 1 11 0 15 13 9 11 1 9 0 7 0 2 7 3 9 0 11 1 3 0 0 0 9 0 9 7 9 2 15 13 3 1 0 9 2
15 1 10 9 1 3 0 9 13 9 11 11 12 0 9 2
34 1 0 2 3 7 3 14 13 9 2 16 4 13 2 0 9 2 11 16 0 9 7 16 4 13 10 9 1 9 3 7 3 13 2
22 0 7 13 3 0 9 2 9 3 11 11 13 13 3 3 0 9 0 0 0 9 2
20 13 15 15 2 16 0 9 11 1 9 1 11 13 10 0 9 11 0 9 2
13 11 11 15 13 1 0 9 11 11 2 11 2 2
28 9 0 9 11 1 0 11 13 9 2 15 4 1 9 0 9 9 2 11 11 13 9 1 9 12 9 9 2
28 1 11 13 10 9 13 9 0 9 2 1 15 15 0 9 13 3 2 16 3 13 9 10 9 1 0 9 2
27 1 9 15 13 7 3 0 9 9 2 16 1 0 9 13 1 0 9 1 9 7 9 1 9 9 11 2
15 3 4 3 13 2 10 9 13 9 0 9 1 0 11 2
26 9 13 9 0 9 2 16 1 9 4 1 11 13 14 12 9 2 16 9 0 9 15 3 13 12 2
18 1 9 1 10 9 13 9 9 1 9 9 0 2 9 2 11 11 2
22 9 11 2 12 1 12 9 1 11 2 15 13 9 9 9 2 13 9 1 11 13 2
28 1 0 9 10 9 11 11 9 13 9 1 10 2 16 4 11 13 0 9 1 9 9 7 0 9 1 11 2
3 9 0 9
6 13 3 9 10 9 13
5 11 2 11 2 2
26 16 9 0 0 9 11 11 13 1 0 9 9 9 0 1 9 9 2 0 9 1 9 13 15 13 2
22 9 9 0 9 4 3 13 0 0 9 11 11 7 1 9 1 0 9 13 13 9 2
28 2 15 15 15 13 2 16 15 1 10 9 13 12 9 2 15 9 1 9 13 2 2 13 15 3 11 11 2
26 3 4 3 13 2 9 13 3 2 16 12 9 11 11 2 11 11 7 11 11 13 9 1 11 11 2
21 1 0 9 13 10 9 2 15 3 2 13 2 16 11 13 0 9 1 0 9 2
34 9 9 1 9 9 13 1 0 9 1 0 9 9 7 1 9 2 15 13 9 1 15 2 16 3 1 9 13 9 0 9 13 9 2
13 16 15 9 13 7 11 11 2 9 0 9 13 2
9 3 3 13 9 0 0 9 13 2
7 3 3 13 9 0 0 9
12 0 9 1 9 11 13 13 0 9 9 1 9
36 9 1 9 2 9 7 0 0 9 1 0 9 9 12 13 1 9 3 9 11 0 9 3 0 9 2 15 13 13 0 2 0 7 0 9 2
14 0 9 13 1 0 11 7 11 0 0 9 1 9 2
13 10 9 1 12 9 1 0 9 13 7 3 0 2
23 1 0 9 1 11 7 9 13 12 9 0 9 2 9 0 9 7 0 0 9 12 9 2
26 1 9 13 2 16 15 3 0 9 9 1 11 13 1 9 1 9 7 3 13 13 1 9 0 9 2
8 1 9 15 13 14 12 9 2
9 1 9 13 3 1 0 9 9 2
19 9 9 13 1 0 9 9 1 0 9 7 9 11 11 11 1 9 9 2
11 11 13 1 9 1 0 9 9 9 9 2
13 13 9 1 15 2 16 1 10 13 9 3 9 2
32 9 2 1 15 15 1 9 13 0 9 7 13 3 1 9 2 13 4 13 1 0 9 9 0 9 1 9 9 1 12 9 2
27 2 13 15 9 2 16 9 13 2 7 13 15 13 1 0 9 2 2 13 9 0 9 9 9 11 11 2
21 1 9 13 9 0 9 13 3 1 9 9 9 11 2 11 2 11 7 10 9 2
30 1 9 13 12 9 1 0 9 1 0 9 2 9 9 1 11 7 0 9 1 9 1 9 1 12 9 9 1 11 2
10 0 9 1 9 0 9 13 1 9 11
5 11 2 11 2 2
15 9 12 0 11 1 0 9 1 0 9 11 15 3 13 2
32 2 3 9 13 12 9 7 1 0 12 9 3 13 13 2 2 13 15 3 9 11 11 1 9 11 2 9 0 9 1 11 2
21 2 0 13 2 16 9 13 9 12 11 2 1 15 15 3 13 0 9 9 2 2
27 10 9 13 2 16 9 15 13 1 0 0 9 3 2 16 15 11 13 9 7 13 1 15 13 1 9 2
16 0 9 15 3 13 2 10 9 3 1 9 13 13 7 11 2
15 1 15 9 11 11 2 2 9 13 1 9 9 3 0 2
19 0 9 13 2 16 11 13 1 9 0 9 1 9 7 0 9 1 9 2
9 1 9 9 9 13 1 9 9 2
11 15 13 0 9 2 15 15 3 13 2 2
23 0 2 12 0 9 1 11 2 4 13 14 3 7 1 0 0 9 4 1 0 9 13 2
4 9 3 1 9
5 11 2 11 2 2
42 0 9 1 9 0 0 0 9 11 1 11 7 11 1 11 2 1 15 13 1 9 12 0 11 11 7 0 12 11 4 3 13 2 13 1 0 9 1 9 1 11 2
34 3 15 9 0 9 2 15 3 13 1 11 2 13 3 2 16 4 12 9 9 2 3 1 11 7 11 2 13 1 0 9 3 13 2
27 1 9 4 13 12 0 1 9 1 12 1 12 9 2 1 15 12 9 13 1 9 9 0 11 11 11 2
22 0 9 0 9 4 13 1 0 9 9 0 9 2 9 0 9 2 9 7 0 9 2
7 9 11 11 2 11 2 2
17 0 9 7 9 2 0 0 9 11 11 4 13 1 11 10 9 2
10 15 13 9 0 0 9 1 0 9 2
19 3 3 12 2 9 4 1 9 13 9 11 11 7 0 3 0 9 9 2
20 9 13 3 13 9 0 9 9 11 11 11 2 15 13 12 0 9 7 9 2
13 0 0 9 13 13 1 9 0 0 7 0 9 2
4 9 1 9 9
5 9 1 9 3 0
5 11 2 11 2 2
34 9 0 9 4 1 11 13 9 1 0 9 0 0 9 1 9 11 11 2 15 1 0 9 1 3 12 9 9 1 9 13 0 9 2
33 1 0 12 9 15 13 12 9 1 9 0 9 2 9 2 1 3 0 9 2 15 3 13 1 10 9 7 0 0 7 0 9 2
24 2 10 0 9 13 10 0 9 1 9 9 1 0 9 2 2 13 15 3 9 9 11 11 2
26 2 0 13 13 15 1 0 9 2 15 13 1 9 2 7 1 0 9 15 13 9 7 3 13 9 2
13 13 9 0 9 2 15 9 7 3 3 13 2 2
27 1 0 9 9 15 1 9 13 3 12 3 0 9 7 1 0 9 13 9 1 12 9 0 9 1 9 2
18 10 12 9 13 0 9 0 9 2 15 15 13 1 9 9 1 9 2
3 9 0 9
5 11 2 11 2 2
26 12 9 1 9 7 0 9 1 0 9 3 12 9 13 3 1 11 11 11 12 9 1 3 0 9 2
12 9 0 9 15 13 1 0 9 0 9 11 2
23 9 9 4 13 9 1 0 9 1 11 2 0 12 13 0 9 1 9 7 0 1 11 2
23 1 3 0 9 12 9 3 13 9 0 11 1 9 0 9 9 1 0 9 1 12 9 2
3 9 1 9
6 0 11 2 11 2 2
22 1 0 13 3 9 9 0 9 1 0 0 9 9 0 9 0 9 0 11 11 11 2
33 2 13 15 15 0 9 2 9 2 7 7 3 9 2 0 9 7 9 7 0 9 2 1 15 15 3 1 15 13 14 14 12 2
35 3 15 0 9 2 15 13 10 0 9 2 13 3 0 1 12 2 9 13 0 9 9 0 9 0 9 2 15 4 13 9 0 9 2 2
9 9 1 9 0 9 13 12 9 2
21 13 9 2 16 15 2 15 1 10 9 13 2 4 13 9 0 9 0 9 13 2
4 0 9 13 9
8 1 9 9 15 13 13 1 9
6 0 11 2 11 2 2
13 0 0 0 9 13 3 13 1 0 0 0 9 2
7 13 9 11 7 11 0 2
7 1 9 9 15 13 13 2
10 2 3 4 13 9 1 12 9 9 2
9 3 9 1 9 1 9 9 13 2
20 16 4 15 13 1 9 2 3 1 12 7 12 9 2 2 13 9 2 11 2
14 12 9 13 1 0 9 2 7 15 13 13 0 9 2
14 13 2 16 1 15 13 9 14 12 9 10 0 9 2
19 1 9 1 9 4 3 13 7 0 9 2 16 15 15 10 9 4 13 2
14 2 3 13 3 1 0 9 2 9 1 9 4 13 2
24 13 4 15 3 1 9 13 0 9 2 15 13 0 9 1 9 7 9 4 15 13 9 2 2
8 13 13 7 9 9 1 9 2
17 1 0 11 13 14 0 2 7 15 3 13 9 1 9 0 9 2
8 9 1 9 11 2 11 2 2
25 9 1 12 9 3 0 0 9 11 11 11 1 11 13 9 9 1 9 2 0 9 11 11 9 2
21 0 9 0 7 0 9 9 1 10 9 9 13 9 0 9 2 0 1 0 9 2
15 1 9 3 13 13 9 1 9 7 9 0 9 1 9 2
30 2 9 13 1 0 9 2 1 10 0 0 9 13 0 9 9 2 9 7 0 9 2 2 13 15 9 9 11 11 2
4 9 0 9 2
19 1 9 7 9 1 9 12 9 13 1 9 3 0 9 9 11 1 11 2
10 9 15 1 10 9 13 1 9 9 2
3 13 9 2
10 12 0 9 13 9 1 11 1 11 2
17 9 13 9 2 9 2 9 7 0 9 1 9 1 12 12 9 2
4 9 1 9 2
15 9 9 0 9 0 9 13 9 0 9 1 0 1 11 2
7 1 9 9 13 12 9 2
4 0 9 3 0
5 11 2 11 2 2
17 1 12 9 0 0 9 7 0 9 13 3 1 11 1 12 9 2
34 0 0 9 13 0 0 2 9 2 11 9 11 7 11 2 1 15 13 12 2 12 2 12 13 7 3 0 12 2 7 12 2 9 2
11 9 9 9 7 3 13 1 9 0 9 2
6 9 13 3 0 9 2
26 1 0 9 13 3 12 9 1 0 11 7 13 15 1 15 2 13 2 14 9 7 9 2 12 9 2
22 1 0 0 9 13 9 1 12 0 9 3 9 9 1 15 7 1 12 0 9 3 2
16 9 0 0 9 13 0 9 12 9 7 9 0 9 12 9 2
13 1 15 13 9 1 9 9 1 9 9 7 9 2
13 9 13 13 3 0 9 2 16 4 15 3 13 13
4 9 13 0 9
7 9 13 9 7 13 9 9
19 3 1 9 13 0 2 9 0 0 9 2 9 2 2 0 1 11 11 2
29 11 11 2 0 2 9 2 2 9 0 9 9 2 3 1 12 2 9 13 9 0 9 2 15 15 13 0 13 2
27 2 11 11 15 1 0 9 13 9 9 2 9 9 13 3 0 9 1 12 9 2 0 9 1 9 12 2
17 13 15 2 16 15 3 13 9 2 2 13 0 9 11 11 11 2
26 1 15 11 2 0 7 0 0 7 0 9 2 13 1 0 9 0 7 13 15 1 0 9 3 13 2
24 9 7 13 0 2 0 9 9 2 1 0 9 2 2 7 13 3 9 13 1 9 0 9 2
27 11 15 7 13 13 0 9 7 9 13 1 0 9 2 7 16 1 12 2 12 2 13 9 1 9 13 2
15 1 0 9 7 9 13 0 9 2 3 9 1 12 9 2
39 1 9 9 9 11 11 1 12 2 9 9 11 13 2 16 2 13 1 0 0 9 13 9 0 1 9 0 9 7 13 9 0 1 9 1 0 9 2 2
14 9 3 13 15 13 9 9 2 7 13 1 10 9 2
19 9 11 7 11 11 15 1 9 12 2 9 1 11 3 13 9 9 9 2
27 11 13 15 2 16 1 9 9 9 1 9 9 13 9 0 9 7 3 9 13 0 9 1 0 9 9 2
27 9 9 9 15 3 13 13 1 9 9 0 9 9 2 12 2 12 9 0 9 0 2 9 1 9 12 2
14 16 0 9 9 13 1 0 9 2 13 15 13 9 2
17 1 0 9 1 9 7 9 9 0 0 9 13 3 13 0 9 2
4 9 1 9 13
5 11 2 11 2 2
31 0 9 1 9 12 0 9 1 9 1 12 2 9 13 2 16 1 9 11 1 11 15 13 0 0 9 0 9 1 9 2
24 1 0 9 9 9 0 9 1 0 9 1 9 1 9 3 1 12 9 1 9 13 1 11 2
9 1 9 13 7 0 9 1 9 2
19 1 9 7 9 13 12 9 9 12 9 0 9 1 9 14 1 12 9 2
26 1 0 9 0 9 9 0 9 9 11 2 9 13 12 3 0 9 1 9 12 2 12 7 12 9 2
20 15 13 1 11 7 9 7 1 12 1 15 9 13 12 9 2 0 1 9 2
34 1 9 0 9 0 0 9 11 11 13 1 3 0 2 7 0 7 0 9 2 10 9 15 1 0 9 13 1 12 9 7 12 9 2
20 9 9 9 3 13 7 13 2 16 9 13 1 0 9 0 0 9 1 9 2
4 0 9 1 9
5 11 2 11 2 2
15 12 9 0 9 1 11 4 13 0 2 9 2 9 11 2
18 1 3 0 9 1 9 9 11 1 11 4 13 13 3 12 2 9 2
16 1 15 9 13 3 1 0 11 1 9 0 9 9 1 11 2
18 0 0 9 2 15 1 11 13 9 2 15 13 3 1 9 0 9 2
22 0 9 9 1 0 9 7 0 9 7 13 2 16 9 3 13 3 12 2 12 9 2
26 9 1 11 2 1 15 0 1 11 3 1 9 13 2 4 13 9 3 1 9 9 2 3 1 9 2
34 16 4 7 1 15 3 13 9 1 10 9 2 1 15 15 1 9 0 9 13 13 12 7 12 9 3 2 13 9 1 0 9 13 2
3 9 1 9
6 0 11 2 11 2 2
15 9 9 7 0 9 13 1 9 9 9 1 10 0 9 2
21 9 15 13 13 0 9 2 0 9 2 9 2 0 0 9 7 0 9 7 9 2
21 0 9 13 9 1 9 0 9 9 2 9 9 9 2 0 9 9 7 9 3 2
12 9 1 9 13 3 3 16 12 9 7 9 2
31 9 4 13 1 9 9 13 9 0 11 1 15 9 1 9 7 1 9 15 13 13 0 0 9 9 7 0 9 1 11 2
3 9 1 9
5 11 2 11 2 2
34 9 1 9 12 7 12 9 13 1 9 3 9 0 9 9 11 1 0 9 2 16 3 1 0 9 13 1 9 1 11 1 0 9 2
17 0 9 1 9 13 2 0 13 1 0 9 1 9 1 0 9 2
18 9 3 1 9 9 13 2 7 3 3 15 1 0 9 13 1 9 2
5 9 9 1 12 9
17 9 1 0 9 3 0 9 13 3 1 9 9 1 0 15 9 2
14 1 0 9 9 15 1 3 0 9 13 13 0 9 2
18 1 0 9 9 2 3 16 9 13 3 1 9 2 3 13 0 9 2
10 9 1 9 3 13 1 9 1 9 2
11 16 7 13 9 2 13 9 1 0 9 2
7 0 9 3 13 1 9 2
5 9 13 1 9 2
14 0 9 0 9 15 15 3 13 13 9 1 9 9 2
5 9 13 3 3 2
6 9 13 7 3 13 2
11 1 0 15 9 0 9 13 9 1 9 2
16 13 3 1 12 9 2 2 1 9 13 6 3 1 10 9 2
3 7 9 2
5 15 13 3 3 2
7 13 15 15 3 3 3 2
14 2 1 9 9 15 13 0 9 9 0 9 0 11 2
15 3 3 13 2 16 0 9 4 1 12 9 13 1 9 2
8 1 9 9 13 3 1 9 2
5 3 3 1 0 2
8 3 1 9 1 9 1 9 2
7 2 0 9 13 12 9 2
22 3 15 7 13 9 0 9 2 15 13 3 1 12 12 2 2 13 9 9 11 9 2
11 1 9 0 0 9 13 7 0 0 9 2
16 1 9 13 10 9 13 1 12 9 7 9 1 9 3 3 2
11 1 15 13 0 3 13 0 9 0 9 2
9 9 1 9 13 12 2 3 12 2
11 1 12 7 3 9 3 15 9 13 9 2
11 9 2 9 2 9 9 2 9 2 9 2
23 2 7 13 15 7 15 2 2 2 2 13 15 1 0 9 1 9 12 9 9 1 9 2
13 3 13 0 9 1 9 7 9 15 13 1 9 2
4 9 15 13 2
11 9 15 13 1 9 7 13 16 0 9 2
14 1 9 9 3 13 2 0 9 16 3 13 1 9 2
18 0 9 9 1 9 1 9 13 1 15 9 0 7 3 13 0 9 2
9 2 9 13 12 9 1 9 12 2
11 1 9 0 9 4 3 3 13 13 9 2
24 12 11 11 2 12 1 12 12 9 4 13 3 1 15 2 16 15 13 1 12 9 12 12 2
15 12 1 15 1 15 13 9 2 2 13 0 9 11 9 2
8 12 9 13 1 10 9 9 2
21 9 0 11 13 1 9 9 1 9 9 3 9 2 0 9 2 9 9 2 9 2
14 9 9 15 3 3 3 13 1 0 9 0 0 9 2
7 3 15 3 13 12 9 2
7 2 3 15 3 13 9 2
12 13 2 16 10 9 1 15 4 13 7 3 2
14 15 15 4 13 9 2 2 13 0 9 0 11 9 2
10 1 0 9 13 9 1 9 0 9 2
23 0 0 9 1 11 1 11 13 3 12 0 9 2 0 11 2 9 2 11 7 11 11 2
13 9 3 13 0 0 9 2 7 0 9 3 13 2
5 14 9 0 9 2
27 16 13 1 12 9 1 9 1 9 3 12 9 2 13 15 15 9 1 15 2 3 15 15 2 13 2 2
11 1 9 13 3 15 12 9 3 1 9 2
21 9 9 13 0 9 2 9 13 7 1 0 9 15 1 9 13 1 9 7 9 2
3 3 13 2
19 1 9 0 9 9 13 0 9 1 9 0 9 2 9 2 9 7 9 2
13 1 10 9 3 3 13 7 0 0 9 2 2 2
8 1 9 13 11 1 0 9 2
4 13 0 9 2
4 3 15 13 2
6 9 9 3 13 9 2
8 1 9 13 9 2 9 2 2
12 9 9 0 0 0 9 15 1 9 9 13 2
12 11 13 0 3 13 1 0 9 1 9 9 2
9 1 11 9 2 1 0 0 9 2
9 2 3 15 13 3 1 9 9 2
10 13 7 0 9 7 1 0 0 9 2
39 1 9 13 13 9 1 9 7 9 2 3 3 7 0 0 9 2 7 3 4 13 9 13 3 0 9 9 11 2 12 2 2 13 9 0 11 11 11 2
13 1 12 9 0 9 13 3 15 9 1 9 15 2
18 0 13 1 15 3 0 0 9 2 1 15 13 0 9 1 0 9 2
8 3 13 9 13 1 0 9 2
17 2 7 16 3 15 13 1 9 2 0 9 15 1 12 9 13 2
20 3 7 1 15 9 13 14 0 9 7 1 0 9 13 2 3 15 15 13 2
28 16 13 9 0 0 9 9 2 7 3 13 15 1 9 10 9 3 0 9 2 2 13 1 9 9 11 9 2
16 12 1 0 9 13 9 7 13 15 2 0 9 0 9 2 2
6 0 9 7 3 13 2
13 9 2 15 3 13 9 9 1 9 2 13 3 2
11 1 9 9 3 1 0 9 13 0 9 2
14 9 0 11 15 1 9 13 13 1 0 9 9 11 2
2 11 11
3 9 2 9
8 9 2 1 9 12 2 11 12
35 9 1 9 0 0 9 11 2 11 2 11 3 12 2 9 2 2 1 15 4 15 13 2 16 12 9 13 9 3 3 1 9 0 9 2
15 4 13 0 9 1 9 2 11 11 2 9 0 9 11 2
36 9 13 2 16 9 11 2 15 1 12 7 12 9 10 9 13 1 9 9 9 1 9 0 9 2 15 13 7 9 2 15 13 1 11 9 2
25 2 3 4 13 9 1 12 2 9 9 2 12 2 9 9 7 9 2 16 0 9 1 12 9 2
12 1 0 9 1 15 13 0 9 1 10 9 2
11 12 10 9 13 1 9 1 9 0 9 2
19 0 9 9 2 0 7 0 9 2 13 3 1 9 2 3 16 0 9 2
22 0 9 1 12 2 9 9 13 1 15 1 9 1 12 9 7 0 9 1 12 9 2
24 9 11 1 12 2 9 4 3 3 13 2 7 1 1 9 0 9 4 15 13 15 3 13 2
12 1 15 13 1 9 0 9 0 1 12 9 2
21 13 15 3 2 16 9 0 2 3 0 9 11 9 9 13 2 16 4 13 15 2
14 16 4 13 9 2 13 0 0 9 2 15 13 13 2
28 3 3 3 4 13 3 1 9 1 12 2 9 2 1 15 4 3 13 9 1 11 2 11 7 1 0 11 2
26 16 15 13 9 1 12 2 9 2 13 4 1 9 9 12 9 1 9 9 1 0 9 1 12 9 2
16 15 13 9 1 0 2 0 9 1 9 12 14 1 9 12 2
8 15 9 13 1 9 9 9 2
19 15 9 15 13 9 9 7 9 9 11 1 9 12 2 12 12 12 2 2
1 9
2 11 12
6 12 9 2 9 2 9
4 12 9 2 9
3 12 9 9
2 12 9
2 12 9
5 12 0 9 9 11
3 12 9 9
4 12 0 9 0
3 12 9 9
7 12 11 13 2 13 2 13
7 12 0 9 2 12 2 2
3 12 0 9
3 12 9 0
4 12 9 13 9
4 12 9 1 0
5 12 1 9 0 11
6 12 0 9 12 1 12
4 12 0 9 9
6 12 1 10 9 7 9
2 12 9
3 12 9 9
2 12 11
3 12 10 9
3 12 0 9
5 12 1 9 1 9
4 12 9 7 15
3 12 9 9
5 9 1 12 1 12
3 12 9 11
2 12 9
3 12 10 9
4 12 9 0 9
3 12 9 11
5 12 0 9 2 9
4 12 11 2 11
19 2 0 9 9 2 9 1 9 1 9 12 1 9 2 1 9 2 9 11
3 0 2 11
14 12 9 13 13 1 0 0 9 1 9 9 0 11 2
5 2 14 12 9 2
13 13 15 3 7 13 15 2 2 3 10 9 2 2
47 3 2 9 13 13 15 3 2 3 3 2 16 1 10 9 13 1 15 0 2 10 9 13 1 9 11 11 2 0 9 2 15 4 1 10 0 9 1 0 0 13 1 0 1 10 9 2
9 0 9 3 7 13 3 0 9 2
21 11 11 2 12 7 12 2 3 13 12 2 9 10 9 2 13 0 9 0 9 2
6 0 9 15 3 13 2
14 16 0 13 2 16 3 12 1 15 13 3 11 9 2
28 9 9 11 13 3 11 11 11 2 7 1 10 9 15 13 3 1 12 9 2 3 15 13 9 9 0 9 2
16 13 15 1 0 9 0 7 1 10 9 2 15 3 11 13 2
25 2 3 2 16 2 9 2 1 0 9 9 13 7 1 0 9 11 11 1 11 1 12 9 2 2
19 9 9 13 3 11 7 11 2 11 1 9 11 9 7 0 11 1 11 2
26 9 13 0 9 3 0 9 2 3 0 9 13 9 1 9 1 9 13 0 9 9 0 15 1 9 2
14 7 3 2 13 15 3 0 9 2 15 13 0 9 2
27 1 9 4 13 9 2 1 15 4 9 13 2 9 9 14 3 9 13 2 7 13 0 9 1 10 9 2
9 9 13 13 14 1 12 2 9 2
8 11 11 2 0 2 11 1 11
7 11 2 9 13 2 0 2
2 11 2
27 1 2 0 2 13 9 0 11 11 11 0 9 1 11 7 11 2 13 2 14 15 11 16 9 0 9 2
24 7 1 9 2 16 4 9 3 13 2 7 13 11 1 0 13 1 0 9 1 0 0 9 2
29 2 16 13 1 11 7 0 9 1 0 9 2 13 15 9 13 15 1 0 9 7 13 0 0 9 2 2 13 2
7 1 0 11 13 9 1 9
24 1 0 9 0 9 0 9 0 9 11 11 13 0 9 1 0 9 11 1 0 9 0 9 2
21 16 7 13 0 9 2 13 15 1 9 3 0 9 9 0 0 9 2 11 2 2
16 1 0 9 0 9 1 0 11 3 9 13 3 12 2 9 2
28 14 1 9 12 2 3 1 11 3 13 0 9 1 9 7 9 2 13 0 9 1 11 12 9 1 12 9 2
9 1 9 12 15 3 13 12 9 2
11 1 12 9 15 15 3 12 13 1 9 2
23 13 9 2 16 1 0 9 13 9 1 15 1 9 1 11 9 2 15 13 3 15 13 2
19 1 12 9 0 0 9 15 0 12 9 1 0 9 13 1 0 9 9 2
24 1 0 9 13 9 0 0 9 2 11 2 2 15 13 9 7 9 1 9 0 9 7 9 2
12 1 9 12 13 12 9 1 0 9 1 9 2
24 16 13 7 13 1 3 0 0 9 2 13 3 9 10 9 1 9 7 13 14 1 0 9 2
19 9 11 1 9 0 9 13 1 9 9 0 9 1 9 2 3 13 9 2
26 9 1 11 13 3 0 2 16 13 10 9 1 9 3 1 0 9 2 15 13 2 16 9 13 11 2
11 0 0 9 13 2 16 11 13 14 9 2
33 2 0 11 13 0 9 9 2 3 15 13 3 7 3 13 2 2 13 11 9 2 0 1 9 1 0 11 1 9 1 0 11 2
17 2 13 1 0 9 2 2 13 7 1 9 1 9 9 0 9 2
40 2 13 15 13 2 15 15 13 2 13 1 9 7 13 1 1 9 0 0 9 2 2 13 9 9 11 11 1 11 2 15 13 1 11 3 16 9 1 9 2
29 9 9 13 14 1 12 2 9 2 3 0 9 11 12 2 1 9 0 9 3 13 9 0 9 0 7 0 9 2
18 16 1 9 12 13 0 9 9 2 0 9 13 1 9 1 0 9 2
17 0 3 12 9 13 9 9 3 3 3 2 15 13 1 9 9 2
20 9 9 13 1 9 2 13 15 1 0 0 9 7 1 10 9 1 0 9 2
13 0 9 0 9 13 9 7 1 0 9 0 9 2
17 1 9 0 9 7 0 9 15 9 13 0 9 16 0 0 9 2
25 1 9 0 9 7 3 13 9 1 9 11 1 0 9 7 9 1 11 2 1 15 9 3 13 2
10 9 1 9 12 7 13 0 9 9 2
24 1 9 13 0 9 7 9 9 7 9 0 9 15 13 0 9 0 9 9 1 9 7 9 2
20 0 9 9 15 13 9 0 0 9 1 9 2 3 15 11 13 3 1 9 2
19 0 9 11 15 13 3 0 1 9 9 2 15 15 0 7 0 9 13 2
25 3 12 0 13 7 9 1 0 11 3 3 1 9 7 1 12 9 0 7 0 9 13 3 9 2
2 11 9
6 9 13 9 11 1 11
9 7 9 13 13 2 9 1 9 2
6 13 15 7 9 1 9
2 11 2
35 9 9 0 1 0 9 11 13 3 1 10 0 0 9 1 9 3 14 9 2 16 10 0 9 1 11 13 9 15 0 9 9 11 11 2
43 16 0 11 11 1 0 11 13 9 0 9 1 9 11 7 13 2 16 13 13 1 12 1 0 9 16 0 9 2 13 15 9 0 9 7 9 1 9 1 0 12 9 2
13 1 0 9 13 3 9 9 1 0 9 13 9 2
20 0 11 15 7 13 0 9 7 0 9 0 15 13 1 9 1 10 0 9 2
34 9 13 9 1 0 0 9 2 9 0 9 1 9 0 9 13 9 1 9 11 1 9 1 0 9 7 0 9 15 13 1 9 9 2
18 15 0 11 3 13 7 13 15 13 1 11 0 12 9 2 16 9 2
7 3 11 13 9 1 0 9
4 1 11 13 9
21 9 0 11 2 10 0 7 0 2 3 13 1 0 11 2 13 3 3 0 9 2
9 7 0 9 13 1 9 3 0 2
27 1 0 2 14 2 1 9 3 14 11 13 15 2 14 2 2 3 10 9 1 9 3 1 9 13 11 2
30 16 1 11 13 1 9 13 0 9 2 1 10 9 2 3 9 9 4 7 4 13 1 9 9 2 13 9 3 0 2
39 13 15 7 9 11 2 3 9 0 9 13 9 0 9 2 3 7 1 9 2 16 2 9 9 2 2 9 9 2 13 3 0 16 9 0 9 7 9 2
27 1 11 7 10 9 11 13 9 1 11 9 0 9 2 3 15 3 13 1 9 0 9 1 0 0 9 2
20 16 4 11 3 13 9 0 9 2 13 1 0 9 9 10 9 1 9 0 2
19 13 15 3 1 9 1 9 9 9 1 9 12 2 3 13 10 9 12 2
20 15 13 1 9 2 16 4 15 9 9 0 9 0 1 11 13 13 0 9 2
24 10 0 9 9 13 2 16 9 3 13 1 9 10 9 2 3 13 2 16 9 4 9 13 2
18 1 9 9 4 13 13 1 0 9 2 1 15 7 13 9 0 9 2
33 16 13 1 9 1 0 9 2 7 2 1 12 2 9 2 3 13 9 1 9 0 2 16 9 0 9 15 3 13 7 1 9 2
33 13 1 15 2 10 9 4 13 0 0 2 14 2 1 0 0 9 2 15 4 15 3 3 2 0 9 2 13 16 9 1 9 2
39 0 9 13 1 11 3 0 2 7 3 3 2 3 3 11 13 0 0 9 2 3 4 3 2 13 10 0 9 1 12 5 1 12 5 1 9 0 2 2
27 0 2 14 2 4 1 0 9 13 3 0 9 7 13 4 1 9 1 9 2 13 15 2 15 13 2 2
4 1 0 9 2
13 0 9 1 11 14 13 2 7 9 9 15 14 13
1 9
13 0 9 1 11 14 13 2 7 9 9 15 14 13
3 13 9 9
33 1 11 7 0 9 11 3 3 13 3 9 9 1 0 9 12 9 2 9 1 0 9 1 10 9 0 11 15 7 3 3 13 2
47 16 15 3 13 13 0 7 0 9 9 2 9 1 10 9 11 15 3 13 1 0 0 9 2 15 4 13 9 0 9 1 9 11 2 3 16 13 15 3 10 9 1 0 9 1 11 2
14 13 15 7 3 0 9 2 7 16 1 9 9 13 2
8 0 9 11 1 11 15 13 2
34 11 3 13 1 12 9 9 2 7 13 15 15 13 7 0 9 1 0 9 9 1 11 2 15 13 3 9 1 0 0 9 3 11 2
17 1 11 13 13 9 3 14 10 0 9 2 16 13 11 7 11 2
27 9 7 11 2 15 1 11 13 1 11 0 9 2 13 3 1 0 0 9 2 16 4 13 9 9 13 2
31 7 16 11 3 1 9 13 0 0 9 2 13 15 15 2 15 15 13 2 3 3 2 13 1 9 0 9 1 9 9 2
18 9 0 11 11 3 13 2 16 13 13 13 1 9 11 10 0 9 2
32 0 9 4 13 9 13 10 9 7 13 15 2 16 11 3 13 9 13 0 2 7 3 13 1 2 9 2 0 7 0 9 2
24 13 15 2 16 15 4 3 13 1 15 2 3 3 15 0 9 13 1 0 9 7 9 9 2
11 3 15 9 11 13 7 13 1 11 13 2
16 0 9 0 9 1 9 13 7 13 9 15 7 3 13 13 2
28 16 15 10 9 2 3 0 1 0 0 2 13 2 4 11 13 0 9 2 7 3 7 9 9 7 0 9 2
6 7 9 9 15 13 2
17 4 13 1 0 9 1 0 9 2 7 1 0 7 0 0 9 2
7 9 1 11 15 13 0 9
14 2 10 9 13 3 0 9 2 7 3 13 9 2 2
19 3 3 13 1 9 11 1 11 0 9 9 11 11 1 0 9 0 9 2
38 0 9 1 2 0 9 2 11 7 11 2 3 3 1 9 11 2 13 1 9 1 9 0 9 1 9 9 9 12 2 0 9 1 9 11 1 11 2
25 0 11 15 13 1 3 0 11 13 2 1 10 0 9 2 2 3 16 0 11 1 0 11 2 2
28 3 1 15 13 13 0 9 0 2 0 9 2 1 15 15 0 9 3 3 3 13 0 9 2 0 9 2 2
31 0 9 4 3 13 13 2 16 0 0 9 13 3 0 7 1 9 1 11 2 7 0 9 13 1 0 9 1 9 12 2
10 3 3 13 15 9 2 3 0 2 2
24 0 9 3 1 11 3 1 0 12 9 13 3 2 0 11 2 2 7 0 2 0 11 2 2
41 11 15 1 9 10 0 0 9 2 3 1 9 12 2 12 9 1 9 0 11 2 13 1 0 9 2 7 3 13 0 13 1 9 7 9 2 16 9 13 3 2
10 11 13 3 14 0 2 7 3 0 2
11 13 15 13 1 0 9 7 1 0 9 2
34 14 1 12 9 0 9 3 13 2 1 9 0 7 0 9 2 1 10 0 9 7 3 3 0 11 3 3 13 9 9 11 7 9 2
11 11 16 0 0 9 13 3 1 10 9 2
27 1 9 12 15 13 12 9 9 0 9 2 15 13 1 0 9 13 2 0 1 9 12 2 0 12 2 2
22 3 13 1 9 12 0 9 2 0 2 0 7 0 1 12 9 11 2 11 7 11 2
11 13 15 7 15 3 0 9 9 1 9 2
18 0 0 9 11 13 1 0 9 13 2 16 2 9 13 0 9 2 2
23 1 12 9 13 9 1 9 10 0 9 7 1 0 7 0 9 2 3 9 13 0 9 2
29 3 1 12 9 15 9 13 9 12 2 3 4 9 13 2 3 16 13 15 1 0 0 9 2 0 9 1 9 2
11 3 15 13 9 11 2 15 13 0 9 2
32 0 9 1 0 9 13 9 9 3 3 1 0 9 2 9 9 2 2 7 2 10 10 0 9 2 2 15 1 15 13 2 2
15 7 15 14 11 1 9 10 0 9 13 10 0 9 11 2
16 7 11 13 3 3 15 0 9 3 3 3 16 0 15 11 2
9 13 1 11 7 11 13 1 15 2
12 11 3 13 7 3 13 0 9 2 1 11 2
6 3 0 2 7 0 2
8 9 3 3 3 13 1 9 2
8 3 7 1 3 3 0 9 2
23 0 9 4 13 1 9 9 2 15 15 3 10 9 13 1 9 1 9 1 11 1 11 2
12 9 13 9 2 15 13 13 0 0 9 9 2
3 11 13 13
7 2 14 2 9 1 11 0
2 11 2
32 9 9 11 11 11 13 2 16 13 1 9 2 16 11 1 0 9 13 0 9 1 0 0 2 0 7 0 9 1 9 11 2
20 2 1 10 9 4 13 1 9 9 2 2 13 1 9 1 0 9 11 12 2
38 9 9 11 10 9 13 1 0 9 0 9 1 11 2 1 15 13 9 9 7 9 9 3 13 7 9 9 0 1 12 2 9 13 3 1 9 13 2
5 13 12 2 9 0
10 13 12 2 9 0 13 4 11 7 11
2 11 2
12 1 11 3 13 12 2 0 9 9 0 9 2
26 9 15 13 9 12 0 9 10 9 2 15 13 12 9 7 1 15 4 1 10 9 13 11 7 11 2
7 9 13 9 0 9 11 2
25 13 2 16 0 9 4 15 1 9 13 15 1 9 13 13 1 0 9 2 7 14 14 1 9 2
33 10 9 1 9 13 2 16 11 2 0 9 9 2 13 0 1 0 9 1 0 12 9 1 0 9 0 0 9 1 9 0 9 2
28 1 9 1 11 13 2 16 4 0 9 11 13 0 9 1 9 9 2 15 9 14 13 2 7 3 3 13 2
7 9 9 0 13 1 9 2
7 1 0 11 13 9 1 9
7 9 1 9 2 9 3 13
2 11 2
16 1 0 0 11 13 1 9 1 9 9 1 9 9 1 9 2
11 3 0 9 13 9 9 1 11 1 11 2
5 3 4 15 13 2
24 1 0 9 13 3 9 1 11 2 15 15 1 11 13 1 9 2 1 9 0 9 1 11 2
19 0 9 13 3 1 0 9 1 11 2 0 9 7 0 9 1 9 13 2
25 3 1 0 11 15 13 1 0 12 9 13 0 9 0 9 1 0 9 9 14 1 0 9 9 2
9 1 11 4 13 3 9 1 11 2
6 11 13 3 2 16 13
6 1 9 13 12 12 9
2 11 2
15 9 0 9 13 3 2 16 3 13 2 13 3 9 11 2
19 1 12 9 9 13 9 0 16 9 2 16 9 13 14 12 9 0 9 2
15 0 9 15 13 9 1 9 2 9 2 9 7 0 9 2
11 14 12 9 9 13 1 9 1 0 9 2
11 0 0 9 1 11 13 3 14 12 9 2
14 0 9 1 9 0 9 1 9 12 13 14 12 9 2
4 11 1 0 9
5 0 9 9 13 9
2 11 2
24 0 0 9 15 1 0 9 0 9 1 9 11 7 3 13 9 1 9 2 9 7 0 9 2
28 0 9 13 1 0 9 1 9 11 7 0 11 1 0 9 1 11 2 16 0 9 13 0 9 1 9 11 2
11 14 1 11 13 1 12 9 7 12 0 2
20 0 9 2 15 3 3 13 1 9 9 1 0 9 0 9 2 13 0 9 2
10 1 0 9 13 9 7 0 0 9 2
11 9 13 13 1 0 9 1 9 1 9 2
12 9 13 0 9 2 15 13 0 9 0 9 2
17 0 9 13 9 9 11 2 3 13 9 0 9 7 0 9 9 2
7 9 13 7 1 9 11 2
21 1 15 13 13 13 7 9 9 11 1 0 9 2 15 13 13 3 1 9 3 2
12 7 0 2 7 0 9 15 7 13 13 9 2
19 9 9 9 13 2 16 0 9 15 13 1 11 7 11 2 3 1 11 2
18 1 11 2 3 15 1 9 1 9 13 0 9 2 13 13 0 9 2
26 9 0 11 11 1 9 1 11 13 2 16 10 9 13 11 1 2 0 12 7 12 9 2 0 9 2
35 11 0 9 1 0 9 1 11 13 2 16 10 0 9 4 2 1 12 9 2 13 11 7 3 13 1 12 0 9 7 13 1 0 9 2
20 1 11 13 9 0 9 11 1 0 9 11 11 2 15 13 13 3 9 9 2
26 1 15 13 13 11 7 11 7 3 13 1 9 10 9 0 9 2 15 15 13 3 1 9 1 11 2
7 11 2 0 2 0 7 0
11 1 0 11 15 14 3 13 2 15 13 15
15 1 15 9 0 0 9 0 2 0 9 2 9 11 2 2
20 7 3 1 9 3 0 7 3 2 3 15 1 10 9 13 2 9 1 9 2
34 11 2 1 9 14 1 3 0 16 11 2 13 3 0 9 13 15 0 2 0 9 2 2 0 3 1 11 2 1 11 7 1 11 2
23 13 3 3 9 2 3 0 2 3 0 2 15 4 13 0 9 13 0 9 0 9 9 2
29 16 1 10 0 0 0 9 3 9 13 9 2 3 2 3 7 3 1 10 9 2 16 4 11 13 13 7 13 2
16 11 2 15 3 4 0 9 13 1 9 2 13 14 12 9 2
13 3 13 1 11 2 16 15 3 13 0 0 9 2
20 13 15 2 7 3 2 16 4 15 1 0 9 13 13 9 0 7 0 9 2
23 0 9 2 3 0 9 13 1 0 9 1 0 9 11 7 13 9 2 13 14 3 0 2
16 3 7 0 13 13 2 16 11 13 9 1 0 0 0 11 2
8 3 13 9 2 3 13 9 2
18 7 9 13 1 0 11 9 3 3 0 2 3 3 1 9 3 0 2
36 1 0 9 9 13 1 11 0 0 9 2 13 15 14 12 9 9 2 7 3 15 13 14 9 16 15 2 7 7 9 0 1 9 7 9 2
36 16 13 0 9 9 1 0 9 9 1 9 9 11 11 1 0 9 2 1 11 0 9 0 0 9 2 16 9 9 1 9 2 4 13 0 2
21 9 1 0 11 13 15 0 9 7 13 10 9 2 3 15 1 0 9 13 9 2
22 14 3 15 13 13 2 16 11 13 3 3 13 2 7 16 10 0 9 13 3 13 2
15 1 0 9 3 13 2 9 2 2 15 15 14 3 13 2
7 15 13 3 2 3 13 2
6 7 11 3 13 11 2
18 9 3 13 0 9 1 9 2 7 13 3 0 2 10 13 0 9 2
16 9 3 2 3 13 9 7 1 0 0 0 9 2 13 15 2
28 13 15 7 1 0 0 9 7 13 1 15 9 2 15 4 13 0 9 2 15 4 15 13 13 0 9 11 2
15 3 15 9 2 0 3 0 9 2 13 9 13 0 9 2
11 0 9 13 9 0 9 0 9 0 9 2
26 1 12 9 14 2 10 2 9 13 13 10 9 1 0 9 9 2 16 4 13 9 1 9 1 9 2
5 0 0 9 4 13
2 11 2
5 0 0 9 4 13
2 11 2
31 0 0 0 9 1 0 9 2 15 0 0 9 13 1 0 9 1 9 11 2 15 0 9 7 9 13 3 13 1 9 2
12 9 13 1 12 12 9 9 3 1 9 11 2
32 1 9 9 2 15 15 13 1 12 9 7 9 2 1 12 0 9 2 3 12 9 7 7 9 9 0 9 2 13 12 9 2
14 9 9 13 9 7 9 9 13 4 13 1 10 9 2
9 9 3 1 11 13 12 9 9 2
4 0 9 1 9
5 0 9 7 9 9
17 1 0 9 0 9 9 9 13 0 9 1 10 9 3 0 9 2
29 0 9 7 0 9 13 2 16 0 9 13 1 12 9 2 1 9 12 1 9 12 1 12 1 0 9 9 2 2
8 0 9 13 1 0 12 9 2
12 10 0 9 13 9 1 0 9 1 9 9 2
46 0 9 2 0 9 9 1 9 2 9 1 9 3 9 7 0 0 9 0 0 9 1 9 11 7 0 9 0 11 13 9 1 0 0 9 1 9 9 11 11 1 9 1 9 12 2
8 9 1 9 13 7 9 0 2
17 9 13 1 9 7 3 1 9 0 9 13 2 16 9 9 13 2
9 3 3 13 0 9 1 10 9 2
5 9 13 9 9 2
24 9 13 9 0 9 1 11 2 15 13 0 9 9 2 16 2 0 9 9 13 3 0 2 2
19 13 0 9 1 0 9 2 16 16 9 10 9 13 2 0 9 13 9 2
4 11 11 2 11
4 9 1 9 2
19 9 1 12 9 1 9 2 15 13 1 0 11 2 3 13 1 0 9 2
5 12 9 9 13 2
5 0 9 1 9 2
12 12 0 0 9 15 13 1 9 1 0 9 2
11 13 15 9 0 9 0 0 9 9 11 2
11 1 0 9 15 13 1 9 0 0 9 2
4 9 1 9 2
20 3 12 0 7 12 0 15 13 9 9 1 9 1 9 11 1 9 0 11 2
9 9 4 13 1 9 0 1 9 2
16 13 15 3 9 9 9 9 2 15 13 1 9 0 0 9 2
3 9 13 2
19 9 0 9 0 9 13 3 9 1 9 1 2 0 0 9 9 9 2 2
5 9 13 13 1 9
2 11 2
5 9 13 13 1 9
3 11 11 2
12 3 12 0 9 1 0 9 13 3 1 9 2
25 1 9 9 15 13 9 2 15 13 13 0 9 2 16 4 0 9 1 9 0 9 13 3 9 2
20 14 12 9 1 0 9 15 13 1 0 9 9 11 2 3 13 13 13 9 2
17 0 9 7 9 13 9 9 1 0 9 0 7 0 9 1 11 2
24 9 13 2 16 3 0 0 9 13 0 9 16 0 0 9 2 15 13 14 1 12 12 3 2
11 9 11 1 9 9 2 9 15 13 1 9
2 11 2
21 0 9 0 9 11 11 2 10 1 9 13 0 9 1 11 2 13 3 0 9 2
21 1 10 9 13 3 14 12 9 0 0 9 2 1 0 12 9 7 9 0 9 2
9 9 9 3 3 13 9 1 9 2
13 9 15 1 3 0 9 13 1 0 9 0 9 2
23 0 9 1 9 13 7 9 9 13 1 0 9 1 9 9 2 3 13 9 9 0 9 2
18 9 2 15 13 1 9 0 9 2 13 3 13 1 12 9 9 9 2
8 1 9 9 3 13 15 0 2
16 0 9 13 0 9 7 13 15 0 9 1 9 2 16 13 2
7 9 13 13 0 0 9 2
13 1 11 15 1 0 9 13 1 12 9 9 9 2
22 9 0 0 9 11 11 3 13 0 9 1 9 7 9 2 7 13 9 1 10 9 2
21 9 0 9 2 0 1 9 9 2 3 13 2 16 13 13 9 7 13 0 9 2
12 1 0 9 9 13 9 9 0 9 11 11 2
14 9 2 15 3 13 9 11 2 13 1 0 9 9 2
12 1 0 9 3 13 0 9 0 7 0 9 2
4 11 13 0 9
4 9 9 15 13
2 11 2
22 0 9 9 3 3 13 9 2 16 15 0 9 0 1 11 13 1 9 1 0 9 2
14 0 9 1 11 3 13 9 7 0 0 9 3 9 2
25 16 15 1 10 9 4 13 0 9 2 13 0 9 9 7 1 9 13 2 13 15 1 9 9 2
40 11 3 13 1 0 9 9 0 0 9 11 2 15 1 9 1 9 0 9 1 11 13 2 16 1 0 9 0 9 1 0 9 3 1 11 4 10 11 13 2
28 11 3 13 2 16 10 9 4 13 13 10 0 9 1 0 9 11 2 1 15 15 13 13 1 9 1 11 2
5 0 9 1 9 9
4 9 13 7 13
2 11 2
10 11 2 0 9 9 2 13 0 9 2
10 0 9 3 13 3 3 16 12 9 2
28 0 9 9 11 11 13 13 0 9 1 9 12 9 9 7 1 12 2 9 9 11 13 15 12 9 0 9 2
11 3 4 3 13 1 12 9 9 10 9 2
10 0 9 4 13 9 2 9 13 9 2
17 9 9 7 0 13 1 9 1 11 1 0 9 1 0 9 9 2
17 9 13 7 13 2 16 4 9 13 9 7 3 4 13 0 9 2
11 3 0 13 1 11 0 7 0 9 9 2
16 9 1 15 3 13 0 9 7 3 2 7 14 1 0 9 2
15 0 9 1 9 13 3 7 9 0 1 0 9 1 11 2
10 9 7 9 7 10 9 3 13 13 2
5 9 11 15 13 13
8 1 9 11 15 4 13 1 9
4 11 2 11 2
23 0 0 9 2 15 3 12 9 13 1 9 11 2 13 3 0 9 0 9 13 10 9 2
21 0 9 15 1 9 9 13 13 1 11 3 1 9 11 7 3 1 9 9 11 2
12 1 12 9 13 1 9 11 7 13 15 13 2
19 1 0 9 15 0 9 13 0 9 2 7 1 0 9 1 0 9 13 2
22 1 0 9 4 1 9 13 7 9 1 0 9 2 7 1 0 9 15 9 3 13 2
29 0 9 9 13 2 16 0 9 1 11 13 13 9 1 9 9 2 15 4 13 13 0 9 9 12 9 7 9 2
16 0 9 4 13 3 1 9 11 2 15 13 3 13 0 9 2
26 1 0 9 13 7 3 13 11 9 9 0 9 11 1 9 2 15 1 0 9 13 1 9 0 9 2
7 1 11 13 9 0 9 2
13 9 1 9 9 11 11 15 13 3 14 1 9 2
14 10 9 3 13 4 9 13 9 9 1 9 0 9 2
33 9 0 9 11 11 11 15 3 1 9 1 11 3 13 3 1 0 11 2 3 13 9 0 9 0 9 11 1 11 2 9 2 2
33 0 9 11 1 10 9 13 0 2 9 1 9 2 15 1 0 9 13 2 7 13 9 2 16 10 0 9 1 9 11 13 0 2
4 11 13 0 9
6 0 9 2 12 9 9
2 11 2
20 9 0 9 0 0 9 11 12 9 3 13 0 9 1 0 11 1 0 11 2
13 10 9 13 7 9 10 9 7 9 0 0 9 2
24 1 9 10 9 13 0 0 9 0 9 9 11 11 2 15 4 1 9 13 1 9 1 9 2
12 11 13 10 9 1 10 9 14 12 9 9 2
26 0 9 9 2 16 13 9 7 9 2 13 9 0 9 11 1 0 9 11 11 2 11 9 1 9 2
16 1 3 0 9 11 13 0 9 1 9 7 9 9 0 9 2
5 9 11 13 1 11
5 9 0 9 13 0
2 11 2
25 1 0 9 0 9 1 11 3 13 0 9 1 0 9 7 9 11 11 9 0 0 0 0 9 2
33 1 0 9 1 0 7 0 9 13 2 16 0 9 1 9 0 1 0 0 9 13 3 13 7 13 0 15 13 3 1 0 9 2
27 1 0 9 1 0 9 13 0 9 9 1 0 7 0 9 2 15 7 2 3 13 2 13 0 0 9 2
35 0 9 1 0 9 13 11 2 11 1 0 2 7 3 9 1 9 13 1 10 9 0 16 1 0 9 0 9 7 13 15 7 0 9 2
5 1 0 11 3 9
2 11 2
5 1 0 11 3 9
2 11 2
20 1 0 11 2 11 2 13 1 9 1 0 9 9 0 9 12 9 1 9 2
26 1 10 9 2 15 9 9 11 11 13 1 2 9 1 9 2 2 15 3 13 10 0 9 1 11 2
17 13 1 0 0 9 2 15 13 13 2 3 10 9 13 9 9 2
21 1 9 13 13 3 3 0 0 0 9 2 3 3 13 0 9 12 9 1 9 2
4 9 15 13 2
20 0 9 13 1 9 1 9 9 2 15 15 13 1 9 9 1 9 0 11 2
15 13 15 15 13 2 16 9 13 0 9 7 13 0 9 2
10 3 10 9 15 9 1 9 9 13 2
7 1 9 15 3 13 3 2
4 3 15 13 2
12 13 15 1 15 0 11 2 11 2 1 11 2
3 13 9 2
20 3 9 0 9 1 11 1 9 11 4 13 12 9 9 11 1 9 9 9 2
13 13 15 15 3 3 0 9 2 15 15 13 13 2
6 9 15 13 0 0 9
5 11 2 11 2 2
38 2 14 11 2 7 11 13 9 0 9 1 11 1 0 9 2 2 13 3 1 0 9 11 11 2 0 9 11 1 11 7 9 9 9 11 2 11 2
31 9 11 2 15 15 1 11 13 2 13 1 9 9 1 0 15 9 0 9 9 1 0 0 9 2 15 13 1 0 11 2
15 2 12 2 9 12 15 13 1 11 13 10 12 2 9 2
11 13 1 15 3 9 2 15 1 11 13 2
41 1 9 15 13 1 0 9 10 9 7 13 1 15 7 9 11 2 2 13 9 11 2 15 9 11 11 11 13 2 16 15 1 9 0 1 0 9 13 0 9 2
17 1 0 0 9 2 15 4 13 3 1 12 9 2 13 13 9 2
27 11 11 1 9 13 3 0 9 1 9 1 11 7 0 9 11 2 3 13 12 1 0 0 9 1 9 2
3 9 1 9
6 0 9 1 9 12 9
6 0 11 2 11 2 2
33 9 9 0 0 9 9 1 11 1 0 11 1 9 1 0 11 7 1 11 13 3 9 12 12 9 7 9 1 9 10 0 9 2
20 1 0 9 15 13 9 0 9 9 12 1 0 11 1 11 7 11 1 11 2
32 2 13 9 1 9 12 2 13 15 1 15 2 16 4 3 0 9 13 3 3 0 2 2 13 9 0 9 1 11 11 11 2
16 9 0 9 13 2 16 1 9 9 1 9 13 13 0 9 2
13 1 9 3 13 9 2 16 11 9 9 12 13 2
25 1 15 3 9 11 11 11 13 2 2 9 15 13 9 9 2 13 3 1 3 0 9 9 9 2
13 0 0 9 13 9 9 1 0 9 1 9 11 2
16 1 0 9 9 1 0 11 15 13 0 9 0 9 0 9 2
3 11 1 9
8 0 9 1 11 3 13 1 11
5 11 2 11 2 2
19 1 0 9 13 11 11 0 2 9 2 12 0 9 11 2 11 12 9 2
17 9 1 0 9 9 13 0 9 3 1 9 13 1 3 0 9 2
12 2 15 13 1 0 9 2 15 15 3 13 2
39 14 12 9 9 15 13 1 9 1 9 10 0 9 1 0 9 7 12 9 13 1 9 1 9 2 2 13 15 11 11 2 0 9 11 11 0 2 9 2
8 12 11 13 1 12 9 9 2
7 3 13 4 9 13 3 2
15 3 15 11 13 13 1 0 9 9 1 9 12 9 9 2
9 9 13 3 1 9 13 1 11 2
19 2 1 0 9 13 1 9 9 7 9 1 9 2 3 13 13 0 9 2
14 3 3 3 7 3 4 15 13 13 3 1 10 9 2
8 1 12 9 13 1 0 9 2
20 3 3 13 9 1 9 9 2 0 9 9 2 9 7 9 2 13 11 11 2
10 10 9 11 13 1 9 11 3 13 2
16 13 15 2 16 1 9 0 0 11 11 4 13 1 11 0 2
14 0 9 13 1 9 11 3 0 7 3 0 16 11 2
24 3 0 11 13 9 11 2 11 1 9 0 11 2 15 13 0 9 1 0 9 7 0 9 2
3 1 9 9
23 1 10 9 13 7 1 9 2 1 15 13 9 9 2 7 1 15 2 15 13 0 9 2
9 1 0 9 9 0 9 11 0 11
38 0 9 2 1 9 12 2 9 12 13 9 10 9 9 11 11 9 11 3 1 9 2 16 15 1 9 13 3 3 0 0 9 11 3 2 2 14 2
7 9 1 15 13 15 0 2
18 15 15 13 1 15 2 16 4 0 9 13 2 16 4 13 9 9 2
16 13 9 2 3 1 15 13 0 9 2 16 9 13 0 2 2
19 3 13 2 16 13 9 0 9 0 9 2 15 1 9 11 11 7 11 2
23 10 0 9 14 3 13 0 9 10 9 7 10 0 9 1 9 2 15 2 3 2 13 2
26 9 7 9 10 9 13 3 1 0 9 3 0 2 16 3 15 13 9 11 2 7 7 7 10 9 2
55 13 1 15 2 16 15 3 13 9 9 2 15 15 13 13 13 12 9 7 3 1 0 9 11 2 7 0 9 9 10 9 13 2 7 1 9 0 13 4 2 16 10 9 3 13 2 0 2 0 9 7 1 0 9 2
12 13 1 9 9 9 2 9 2 9 2 2 2
58 13 2 16 1 0 9 13 14 3 3 13 1 10 0 9 2 7 16 3 1 15 13 7 9 0 9 7 9 1 9 0 9 2 13 3 1 0 9 9 2 1 15 1 9 13 9 0 9 10 9 2 7 9 9 7 9 9 2
7 11 2 11 2 11 2 11
1 9
3 9 1 9
12 0 0 9 15 13 1 9 1 9 7 9 2
12 1 0 9 10 1 9 0 9 13 1 9 2
12 3 2 9 15 13 2 7 16 3 2 13 2
6 9 9 13 3 0 2
14 1 12 2 9 13 1 9 9 1 9 1 0 9 2
23 10 9 13 13 3 3 7 1 9 7 9 1 9 3 3 2 16 13 0 9 0 9 2
28 1 10 9 4 10 0 9 13 14 9 9 0 1 9 0 0 9 2 7 7 3 0 9 0 1 0 9 2
30 0 9 7 9 15 1 9 13 1 12 2 9 13 0 13 1 9 1 9 7 1 9 9 13 0 9 0 0 9 2
42 9 9 1 15 2 16 9 13 7 9 2 13 3 0 9 2 7 1 1 0 9 2 3 15 3 1 10 9 13 13 2 15 3 1 12 2 9 13 13 1 9 2
23 7 16 4 3 4 0 9 3 13 2 13 9 2 15 4 13 10 0 9 1 9 9 2
25 2 0 2 0 9 3 13 3 1 10 9 1 9 7 9 4 13 9 9 1 9 9 1 9 2
5 15 1 10 9 2
12 9 3 13 10 0 9 2 15 13 10 9 2
20 7 16 4 10 9 3 13 1 9 9 2 0 2 9 2 15 13 3 13 2
23 3 13 0 15 13 2 16 1 9 0 0 9 13 9 2 15 15 13 3 14 3 13 2
12 0 9 13 1 0 9 1 9 9 11 11 2
20 7 13 3 0 9 2 16 9 1 0 15 9 9 9 1 9 3 3 13 2
6 7 15 13 0 9 2
25 7 3 0 9 3 13 9 0 9 2 15 15 13 2 16 4 9 13 13 1 0 9 9 9 2
23 0 9 15 13 3 1 12 9 1 0 9 2 15 4 13 13 0 9 9 1 9 9 2
2 11 11
3 0 0 9
15 9 11 13 3 0 9 0 9 2 1 0 0 9 2 2
18 7 1 9 12 2 12 2 12 15 13 0 9 0 9 9 1 9 2
18 1 0 9 9 15 13 2 16 1 10 9 4 13 9 1 0 9 2
16 13 15 3 9 1 0 9 1 0 9 7 0 9 9 11 2
26 1 1 10 9 4 13 0 13 2 16 9 2 0 2 9 15 13 1 9 0 9 7 13 0 9 2
5 9 13 7 0 2
19 9 12 2 15 13 1 9 9 13 13 9 2 1 15 13 2 9 13 2
26 9 12 3 13 9 9 2 1 15 9 13 9 2 16 4 15 2 13 2 10 9 3 1 10 9 2
17 10 9 4 14 3 13 9 0 9 2 7 1 9 3 13 9 2
15 0 9 4 3 13 13 1 10 9 15 10 9 7 9 2
28 9 12 3 13 0 7 0 9 13 15 9 10 9 1 9 2 15 1 15 9 13 2 16 15 15 3 13 2
14 1 9 12 13 13 9 3 2 0 9 7 0 9 2
39 9 2 15 4 13 9 0 9 2 4 3 13 13 14 10 9 2 7 3 2 1 9 9 2 7 9 15 2 15 15 9 1 0 9 3 2 13 2 2
25 9 2 16 1 0 2 9 13 1 9 0 9 9 2 9 7 0 2 13 14 3 14 3 0 2
18 3 2 1 0 2 9 2 0 2 13 9 13 1 10 9 7 9 2
27 1 0 9 9 4 15 3 9 13 13 1 9 2 1 15 4 15 1 0 9 13 9 9 1 9 9 2
16 10 9 0 9 4 3 3 13 9 1 9 0 9 0 9 2
24 0 9 9 9 2 15 15 13 9 9 2 9 2 1 9 0 0 9 2 13 10 0 9 2
12 1 9 12 13 3 2 13 1 9 0 9 2
10 14 3 13 13 2 15 15 15 13 2
15 13 3 2 9 1 9 9 1 11 1 0 9 0 9 2
18 7 13 3 3 9 9 9 2 13 2 14 10 9 1 9 1 9 2
24 0 15 3 13 9 12 2 15 13 9 9 13 0 9 0 9 2 13 2 14 15 0 9 2
12 1 2 0 2 9 13 3 9 3 0 9 2
27 3 9 12 2 15 3 2 13 2 16 4 9 9 13 0 7 0 9 7 0 9 1 3 16 12 9 2
10 10 9 3 3 13 9 1 0 9 2
24 9 12 2 16 9 0 9 2 13 9 9 2 7 13 7 1 9 1 9 0 9 7 9 2
12 0 9 9 13 12 1 0 9 1 9 9 2
15 0 9 2 1 0 0 9 2 13 0 13 1 10 9 2
22 1 9 2 16 4 15 9 13 1 0 9 2 13 4 15 1 0 2 9 3 9 2
13 9 9 13 7 0 1 9 0 7 0 9 13 2
2 11 11
11 13 4 15 11 11 2 9 9 0 9 11
32 1 9 9 0 9 0 9 2 0 2 9 2 2 11 11 4 9 13 7 1 9 9 2 15 13 0 9 11 1 15 9 2
6 13 10 9 3 0 2
3 3 13 2
21 9 9 2 3 9 9 2 13 1 9 1 10 9 3 9 13 3 0 0 9 2
16 9 9 1 9 2 9 9 7 0 0 9 13 1 9 0 2
2 0 9
7 13 4 13 3 0 9 2
8 9 7 13 13 1 9 9 2
21 9 3 13 13 2 3 15 13 12 0 9 2 15 4 13 1 9 10 9 2 2
6 11 2 11 2 2 11
11 1 9 9 15 13 9 13 1 9 9 2
13 1 10 9 13 13 2 16 4 1 9 3 13 2
23 13 2 14 9 1 0 9 9 1 9 9 2 13 9 1 9 9 9 13 9 9 9 2
3 2 11 2
30 0 9 9 7 1 0 9 1 9 2 7 3 0 9 9 1 9 2 13 9 9 7 9 0 9 12 1 0 9 2
22 0 9 3 13 1 3 0 9 1 9 7 3 0 9 0 9 13 0 9 0 9 2
27 1 0 9 3 1 9 7 9 15 13 0 7 0 9 0 9 9 2 3 15 10 9 13 16 9 0 2
16 1 0 9 15 9 0 9 13 1 12 7 13 12 9 9 2
13 1 9 12 15 13 9 14 1 12 9 9 3 2
18 9 9 13 7 0 9 2 3 1 0 9 0 11 7 9 0 11 2
13 9 1 10 9 13 0 1 9 7 13 0 9 2
12 3 13 9 3 0 9 2 3 9 1 9 2
10 0 9 11 4 13 0 9 1 11 2
26 10 0 9 2 1 9 12 9 2 9 2 7 13 9 1 11 1 0 9 2 15 13 13 0 9 2
22 1 0 9 13 7 11 2 7 3 15 13 1 9 0 9 1 9 9 1 0 9 2
16 0 9 11 2 11 13 9 1 11 7 13 9 0 0 9 2
20 9 0 9 1 9 13 9 2 7 1 9 0 9 1 9 9 13 0 9 2
23 1 12 3 0 9 3 11 7 11 13 9 0 9 0 9 2 11 12 9 15 9 2 2
20 1 9 15 3 13 3 12 9 9 2 1 15 1 0 9 13 14 12 9 2
21 0 9 1 9 13 0 1 0 11 1 0 9 12 9 9 7 9 12 9 9 2
19 9 10 9 15 3 13 1 0 0 9 1 11 2 1 9 7 0 11 2
16 9 13 3 9 0 9 2 1 10 9 13 7 11 1 11 2
19 1 0 11 15 3 13 9 2 16 13 0 9 1 0 9 0 9 9 2
3 9 9 13
17 11 11 13 12 2 9 1 9 9 9 7 0 9 0 0 9 2
8 4 15 3 3 13 1 11 2
9 13 15 3 0 9 1 0 9 2
36 16 9 9 9 9 13 2 16 9 15 1 10 0 9 9 1 0 9 1 9 1 0 9 13 1 9 9 2 2 15 13 9 9 9 2 2
28 10 9 13 9 9 9 11 11 1 9 2 2 0 15 15 16 9 9 1 9 9 2 2 13 15 1 9 2
5 0 9 1 11 11
14 9 9 12 9 9 11 11 4 13 9 3 12 9 2
41 13 15 1 12 9 1 9 11 1 11 2 12 1 9 9 7 9 2 12 7 12 1 0 9 2 12 1 9 0 9 7 1 0 7 12 9 1 9 0 9 2
19 3 15 7 13 9 1 9 1 11 2 3 1 9 9 1 0 0 9 2
30 1 0 9 3 13 0 9 12 9 2 1 15 13 13 0 12 9 9 7 9 2 1 10 9 15 13 3 1 9 2
23 1 9 9 9 0 2 9 2 11 11 11 13 7 1 9 0 13 3 15 9 1 0 9
36 15 13 1 9 1 9 9 9 1 0 9 2 1 15 0 9 13 2 16 15 9 13 9 9 7 9 11 11 2 15 13 1 9 12 9 2
20 13 3 9 2 16 15 9 9 13 13 9 1 9 7 13 15 1 9 9 2
23 2 9 0 9 9 3 13 3 0 2 2 13 15 3 9 9 9 7 9 11 11 11 2
38 2 3 7 13 2 16 9 9 15 1 0 9 2 13 1 9 2 13 3 3 7 3 3 1 9 9 2 3 4 15 0 9 3 13 3 0 2 2
27 11 11 3 13 10 9 2 15 13 9 11 11 1 9 13 9 1 0 9 2 7 13 3 10 0 9 2
16 10 9 3 13 2 2 9 16 9 9 9 3 13 10 9 2
22 0 9 9 2 1 15 15 13 9 0 9 2 13 7 1 0 9 16 1 9 2 2
18 13 15 1 9 11 9 7 11 11 2 1 15 15 13 0 9 11 2
14 10 9 0 9 13 2 16 0 9 9 11 11 13 2
11 0 9 1 9 9 13 3 0 0 9 2
38 4 13 0 0 9 9 2 0 9 15 13 13 14 1 0 9 7 1 9 0 1 0 9 1 15 2 16 13 0 3 13 1 0 0 9 0 9 2
12 9 9 13 14 1 9 0 9 1 0 9 2
15 0 9 13 14 1 9 9 3 0 0 9 0 0 9 2
20 1 9 10 9 11 11 1 9 12 9 4 1 9 9 13 9 1 0 9 2
18 1 9 1 9 0 9 1 11 15 1 0 9 13 9 1 9 9 2
9 11 7 9 1 9 0 9 13 2
16 0 9 11 11 13 12 9 9 2 15 13 0 9 12 9 2
32 1 0 9 13 9 9 11 2 12 9 9 2 11 11 2 12 9 2 11 11 2 12 9 7 11 9 11 2 12 9 9 2
14 9 0 9 0 9 13 12 9 7 9 12 9 9 2
20 1 9 9 7 0 9 9 4 7 13 13 0 0 9 9 7 10 0 9 2
11 7 1 9 9 9 9 1 10 9 13 2
26 0 13 3 0 9 1 9 0 2 11 11 2 9 11 2 0 9 11 2 9 7 0 9 11 11 2
8 11 11 2 11 11 2 11 11
12 9 11 1 0 11 13 0 11 12 9 9 2
8 2 13 15 3 7 1 9 2
10 9 13 0 7 1 10 9 3 0 2
19 1 0 9 15 3 13 2 2 13 15 3 11 11 2 0 9 9 11 2
22 9 10 9 1 9 3 13 12 9 9 2 15 13 2 3 9 9 2 12 9 9 2
23 13 9 15 1 10 9 13 7 1 0 12 3 0 9 2 10 0 9 3 13 1 9 2
26 1 0 9 0 9 1 0 9 13 0 9 2 3 1 12 9 13 9 1 11 14 1 3 0 9 2
24 15 4 13 9 0 9 9 1 0 11 1 9 0 9 2 15 10 0 9 13 3 3 13 2
3 2 11 2
7 9 11 2 11 1 9 13
17 0 9 9 1 9 10 9 9 1 0 9 13 1 9 1 11 2
24 10 9 0 9 9 0 0 9 0 9 0 9 11 11 15 13 13 9 1 12 1 12 9 2
32 2 13 3 1 0 9 10 9 2 2 13 9 11 2 2 3 1 9 1 0 9 13 1 0 9 13 12 9 1 0 12 2
14 9 10 9 1 0 9 13 3 3 1 10 9 13 2
7 1 10 9 4 15 13 2
23 13 3 1 0 9 2 0 9 2 9 2 0 0 9 2 9 2 9 2 9 7 9 2
27 2 9 1 9 1 9 1 9 0 9 13 1 9 0 9 1 9 7 9 2 9 2 0 9 1 9 2
16 1 0 9 13 1 9 9 9 1 11 1 9 12 7 12 2
11 3 13 9 0 9 1 0 0 9 11 2
17 1 9 9 7 13 4 1 9 0 2 0 9 13 0 0 9 2
18 9 11 13 7 9 2 16 15 13 3 10 9 9 9 1 0 9 2
36 2 1 10 9 4 13 3 1 12 2 9 0 13 15 9 1 9 1 11 2 2 13 9 11 2 2 7 15 13 12 1 3 0 9 2 2
18 1 9 11 11 4 1 9 9 1 0 9 7 11 13 13 1 9 2
9 3 0 9 15 13 9 0 9 2
18 13 15 9 0 9 1 9 12 2 12 2 3 4 13 1 9 9 2
21 2 9 13 10 2 1 10 9 13 0 2 16 4 0 9 13 15 2 15 0 2
13 3 0 9 13 3 1 9 2 2 13 9 11 2
3 0 9 13
36 9 0 2 0 9 0 0 9 2 11 2 11 11 3 13 1 11 11 2 16 4 13 0 0 9 9 2 7 13 3 13 9 1 0 9 2
32 1 0 9 1 9 9 0 9 11 11 13 2 16 0 9 1 11 13 2 3 0 2 2 16 1 11 13 2 3 0 2 2
21 0 0 9 3 13 2 16 1 0 9 13 0 0 9 1 0 12 1 12 9 2
19 13 15 0 9 0 9 7 9 0 0 9 1 9 1 0 9 0 9 2
48 0 9 9 1 0 9 1 9 0 9 4 13 13 0 0 9 2 9 2 3 2 7 13 15 14 2 16 9 13 3 13 9 2 16 3 15 13 0 9 2 13 3 1 9 0 0 11 2
12 9 13 2 16 3 0 9 9 13 0 9 2
15 9 2 15 13 1 0 9 2 13 3 13 15 10 9 2
9 1 0 9 15 13 9 0 9 2
13 2 7 9 3 3 13 1 9 2 2 13 9 2
12 3 13 3 1 11 2 16 4 13 0 9 2
22 9 2 0 1 9 1 11 7 11 2 4 13 13 0 9 1 9 0 9 0 9 2
8 0 9 13 1 15 3 0 2
20 16 9 13 0 9 2 3 1 9 0 9 13 10 9 13 2 13 0 11 2
11 9 3 1 0 9 13 1 3 16 9 2
20 1 9 13 1 0 0 9 11 1 0 9 9 1 9 0 9 7 0 9 2
43 1 9 11 11 2 9 1 0 11 11 2 2 4 1 9 13 0 0 9 11 1 9 9 2 16 4 13 13 1 0 9 0 9 2 7 9 4 13 2 1 15 13 2
8 0 9 11 14 13 9 9 2
8 9 13 1 12 2 12 9 2
11 9 9 15 3 13 7 1 9 1 11 2
19 1 9 0 9 13 0 9 1 0 9 1 9 9 0 9 7 0 9 2
12 9 1 11 13 1 9 1 12 5 12 9 2
4 11 13 10 9
38 9 1 0 9 9 15 3 3 13 10 9 1 9 0 9 9 13 2 0 0 9 2 1 0 9 9 0 1 0 9 1 11 2 11 7 0 11 2
23 13 15 0 9 1 9 14 12 0 9 0 11 1 0 9 9 9 1 11 7 0 9 2
28 0 9 9 9 0 2 9 1 0 9 11 3 13 9 1 9 9 1 11 1 12 5 1 9 1 0 9 2
21 1 9 13 3 1 9 1 9 1 9 2 3 9 0 2 9 13 9 0 9 2
22 15 4 3 13 9 1 11 2 14 3 1 10 9 2 7 3 1 12 2 12 9 2
26 9 9 0 2 0 9 7 0 9 1 9 9 2 16 13 1 0 9 2 3 13 9 0 9 11 2
29 9 0 9 3 15 13 1 15 2 16 11 2 7 11 7 11 2 4 3 13 1 9 9 16 9 1 0 9 2
12 13 1 15 0 0 9 0 1 12 2 9 2
12 0 9 4 13 1 9 0 9 1 0 9 2
33 1 9 10 9 13 0 2 16 16 4 1 10 9 13 2 13 4 7 11 2 11 3 11 0 1 9 7 9 2 0 9 2 2
35 10 9 4 15 3 13 1 0 9 10 9 7 3 4 15 13 1 9 2 16 9 10 9 15 13 3 12 7 12 9 2 3 3 2 2
30 2 0 0 9 2 2 3 1 12 9 2 4 3 13 9 9 7 3 4 3 13 10 9 9 9 1 11 1 11 2
38 0 9 11 1 9 0 2 9 4 13 0 9 0 9 11 2 11 2 15 15 13 1 9 12 2 7 12 2 9 1 0 9 0 9 2 11 2 2
4 11 13 10 9
8 3 4 13 9 1 0 2 9
16 0 9 13 9 11 2 16 4 13 13 9 9 9 1 11 2
42 13 4 13 1 9 2 0 9 2 1 0 9 2 15 4 13 9 11 12 2 9 1 9 9 0 0 9 1 11 1 11 2 11 7 11 2 1 15 0 9 11 2
32 0 9 10 9 13 9 2 3 9 9 2 15 0 2 9 13 3 13 1 0 12 9 2 4 1 15 13 1 0 9 11 2
28 3 3 13 1 9 9 1 9 0 2 9 1 15 9 11 7 14 1 11 2 11 7 11 2 13 0 13 2
12 0 9 0 9 3 13 9 1 9 9 11 2
36 0 9 2 1 10 9 7 0 9 9 2 1 9 13 0 1 2 0 9 2 2 15 13 10 9 9 11 2 16 9 13 9 1 0 9 2
33 13 0 2 16 1 9 9 11 1 9 0 2 9 9 1 12 0 9 15 13 3 0 9 2 15 3 13 1 0 9 0 9 2
25 9 9 0 9 7 9 0 9 11 1 9 9 9 13 2 16 1 9 13 3 1 9 10 9 2
20 11 15 13 13 1 0 0 9 0 9 0 9 2 0 9 2 1 0 9 2
8 13 15 0 9 0 9 0 2
12 0 9 13 0 9 0 9 7 9 0 9 2
8 11 11 13 13 9 7 10 9
5 11 2 11 2 2
46 2 13 13 2 16 9 9 13 15 2 15 4 13 2 2 13 1 10 0 0 9 1 9 9 11 11 2 0 2 9 2 2 9 11 2 11 7 11 0 9 9 7 9 11 11 2
28 16 3 13 2 1 10 9 13 9 3 1 12 9 3 13 0 9 9 1 9 1 9 1 0 7 0 9 2
16 9 9 13 9 15 13 1 0 0 9 7 13 9 10 9 2
11 9 11 3 13 9 0 0 9 9 9 2
32 1 9 9 0 0 9 2 15 15 13 3 1 9 0 9 2 13 1 9 9 0 13 9 9 1 0 9 1 0 9 9 2
24 1 11 11 0 9 1 10 9 13 2 7 1 9 7 13 2 0 9 13 1 9 0 9 2
17 1 9 1 9 9 3 13 1 9 7 0 9 4 13 13 9 2
24 16 13 1 0 9 0 9 1 0 9 11 2 9 11 4 13 0 0 9 1 10 0 9 2
41 1 0 9 1 9 11 11 11 13 2 16 1 9 9 13 13 9 9 1 12 9 1 15 2 16 3 16 12 0 9 13 1 0 2 0 9 1 0 9 9 2
21 9 11 13 2 16 16 4 0 9 13 2 13 13 0 0 9 1 9 0 9 2
5 0 9 9 13 9
33 0 0 9 2 0 9 2 3 0 0 9 2 10 15 13 11 2 3 2 0 9 0 0 9 1 9 9 9 9 0 0 9 2
7 15 1 9 10 9 9 2
26 15 10 0 9 2 15 13 9 7 1 0 0 9 2 15 1 0 9 3 13 7 13 1 9 11 2
11 15 1 12 9 2 4 13 3 0 9 2
36 1 0 9 9 15 7 13 7 0 0 9 7 9 2 3 2 0 2 9 2 7 9 2 3 4 13 14 9 2 7 3 9 11 13 9 2
11 0 9 13 1 9 1 9 0 0 9 2
23 15 3 13 15 2 16 4 1 9 9 7 1 9 11 13 0 9 13 0 16 0 9 2
6 3 15 10 9 13 2
23 13 15 1 15 2 16 4 9 11 13 4 13 0 9 2 16 4 1 15 13 9 3 2
21 16 4 15 13 2 0 9 13 7 1 10 9 7 3 0 0 9 13 15 13 2
2 0 9
22 0 9 7 9 11 11 13 1 9 11 12 2 15 13 1 9 12 2 3 0 9 2
9 13 15 15 7 3 13 1 11 2
46 11 12 1 15 13 14 1 10 9 2 3 13 1 9 9 7 9 11 11 2 11 1 9 0 0 9 2 3 3 1 0 9 9 7 3 1 11 2 1 0 0 9 1 9 12 2
26 11 13 1 9 1 9 2 13 15 9 3 2 0 2 7 13 9 16 0 9 2 15 13 10 9 2
16 1 10 9 13 0 9 13 16 9 1 9 9 7 0 9 2
20 0 9 7 9 1 0 9 0 1 15 9 2 9 10 9 2 13 0 9 2
42 9 1 0 0 9 2 9 0 0 9 2 9 2 9 2 9 0 0 9 2 9 9 2 0 9 1 9 9 2 0 9 2 9 2 9 2 9 7 9 2 2 2
14 0 2 0 15 3 13 1 0 9 1 9 0 9 2
25 9 9 15 13 2 0 9 13 2 0 9 2 9 1 11 2 0 9 10 7 10 9 1 15 2
22 2 11 15 16 0 9 13 2 16 4 9 13 10 9 2 2 13 11 11 2 11 2
12 2 0 9 4 13 2 16 15 13 10 9 2
7 0 0 9 13 3 0 2
23 3 15 7 13 13 2 16 13 9 1 15 0 9 7 3 3 3 4 11 12 13 2 2
3 9 3 0
26 0 0 7 0 9 2 15 15 13 1 11 7 10 9 13 13 1 9 11 2 4 1 9 3 13 2
37 0 1 15 13 7 9 9 1 9 9 11 11 2 2 1 12 3 4 13 9 9 2 16 4 15 13 13 2 16 9 13 13 1 12 1 9 2
5 13 7 0 9 2
12 9 12 9 9 13 9 7 0 9 1 9 2
5 9 13 9 9 2
19 3 15 9 13 13 2 16 4 15 10 9 13 3 13 0 9 9 2 2
23 9 13 13 0 9 11 11 2 2 9 0 9 13 9 1 9 1 9 1 9 0 9 2
5 1 9 13 9 2
7 9 1 15 13 9 9 2
13 3 0 9 1 1 12 13 1 12 9 1 9 2
21 1 9 9 2 16 0 9 15 1 9 13 13 2 13 7 10 9 1 9 2 2
9 1 9 15 3 13 9 0 9 2
40 1 9 9 13 11 11 2 2 1 9 15 13 1 12 9 3 2 9 15 7 1 9 0 9 3 13 2 16 13 1 15 3 2 16 4 13 13 0 9 2
14 3 7 9 13 9 2 15 9 13 1 12 0 2 2
19 0 9 13 9 0 9 9 7 0 11 11 11 1 12 7 12 9 9 2
6 1 11 9 7 1 9
14 9 1 0 9 15 1 0 9 1 9 9 3 13 2
35 1 9 13 10 9 2 1 9 0 9 7 1 9 9 2 3 15 13 9 0 9 11 11 2 15 13 13 1 12 2 12 2 0 9 2
14 9 7 13 9 3 1 9 1 9 3 12 2 12 2
34 1 9 4 13 11 2 11 2 2 9 9 13 3 9 12 9 2 15 13 9 3 0 1 1 15 2 15 9 13 7 10 13 9 2
32 1 0 9 2 3 9 13 1 12 9 1 9 2 1 0 12 12 2 2 15 4 13 9 7 9 2 13 3 9 12 9 2
21 9 1 9 9 13 15 2 16 4 10 9 13 1 12 9 3 2 16 4 13 2
19 13 7 0 9 2 13 15 15 3 13 9 0 9 7 13 1 0 9 2
10 1 0 9 3 1 9 13 0 9 2
22 0 9 13 1 0 9 3 7 13 15 2 16 3 15 1 9 13 7 0 9 2 2
3 15 1 15
38 1 9 15 13 7 9 0 9 11 11 2 2 9 11 1 9 2 12 13 9 1 0 9 2 1 15 3 12 9 13 9 7 9 3 1 0 9 2
26 12 13 2 16 9 9 2 3 9 2 3 0 9 2 13 13 9 0 0 9 3 1 9 9 9 2
22 9 2 3 13 0 9 2 13 3 1 9 7 9 0 1 9 0 2 2 2 9 2
16 1 0 9 2 13 1 9 1 9 11 2 4 3 9 13 2
39 9 9 13 1 9 0 7 1 9 7 0 9 2 7 2 9 2 13 2 16 9 13 9 2 7 1 15 13 9 2 15 4 13 13 7 9 10 9 2
32 1 9 13 0 2 16 4 4 13 9 9 2 1 9 7 9 13 0 9 2 9 13 13 0 9 7 13 15 3 0 9 2
18 2 1 10 9 13 9 11 1 9 0 9 12 7 9 9 9 3 2
12 13 0 2 16 1 0 9 3 10 9 13 2
3 0 11 0
17 9 0 9 0 11 15 1 9 1 9 0 9 0 9 13 0 2
25 1 12 9 4 9 13 13 1 11 7 1 9 10 9 9 9 13 10 0 9 0 2 9 0 2
25 1 9 9 1 11 2 3 4 13 12 2 9 1 11 2 13 3 0 9 0 2 0 2 11 2
27 0 1 10 9 3 13 2 16 9 3 13 9 7 9 2 7 10 9 3 1 9 11 11 13 15 9 2
7 15 13 3 0 7 0 2
20 13 1 15 7 9 1 0 9 7 0 9 2 14 1 0 0 9 13 9 2
33 9 15 1 9 0 9 9 13 1 9 2 7 1 10 9 2 15 13 13 7 3 13 10 9 2 13 14 9 9 7 0 9 2
10 3 9 10 9 13 9 0 0 11 2
18 13 15 3 1 9 0 9 2 9 9 2 9 0 7 0 0 9 2
14 0 9 1 0 0 9 9 13 11 11 14 1 11 2
8 7 0 9 13 0 9 9 2
14 0 13 0 11 2 15 13 0 1 0 0 0 9 2
9 3 1 15 13 7 0 9 9 2
9 1 10 9 13 0 7 9 9 2
16 12 1 9 10 0 9 13 13 1 0 9 9 1 0 11 2
18 0 9 1 10 9 13 3 0 9 2 3 1 9 12 1 15 9 2
25 1 12 9 7 13 1 0 9 2 7 0 9 9 1 0 9 2 16 4 15 13 13 1 9 2
34 3 0 9 3 13 3 0 16 0 2 9 0 2 13 7 3 0 7 13 9 2 15 4 15 13 13 10 0 9 0 1 0 9 2
16 1 9 13 0 9 2 3 15 0 9 13 0 9 11 11 2
17 7 9 13 11 11 2 0 1 12 1 0 0 9 2 1 9 2
3 9 16 9
23 3 16 9 15 9 11 11 9 2 0 1 9 1 9 11 1 9 11 11 2 13 13 2
11 0 9 0 9 13 1 9 9 7 9 2
19 9 15 13 2 16 13 10 9 2 15 3 3 13 2 3 13 10 9 2
10 3 3 15 13 9 0 9 1 9 2
17 0 9 9 13 3 0 9 0 9 11 11 2 15 13 15 3 2
13 9 13 0 7 0 3 15 2 16 15 15 13 2
23 11 11 2 3 16 0 9 2 13 1 9 9 9 2 11 11 15 3 16 10 9 13 2
11 9 13 13 1 9 2 16 15 13 13 2
26 3 15 13 7 3 13 2 16 9 13 9 0 9 2 9 15 13 1 9 2 7 9 9 9 9 2
9 9 13 1 0 9 11 11 12 2
6 9 3 9 11 11 2
38 9 0 0 9 2 10 9 2 9 11 2 11 2 4 3 13 9 0 0 9 0 0 9 2 9 2 12 2 2 13 0 9 11 3 1 12 9 2
18 9 0 9 1 0 2 11 1 11 2 9 11 13 9 0 0 9 2
31 9 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 7 11 2 11 13 1 9 0 9 0 2 11 11 11 2
5 0 9 0 9 2
20 1 10 9 15 13 1 0 9 0 9 2 15 13 1 10 9 3 0 9 2
7 9 13 1 12 2 9 2
25 9 9 9 2 9 7 9 12 0 11 11 11 7 11 11 0 0 9 3 13 1 0 9 9 2
6 13 1 12 2 9 2
18 0 0 9 9 11 2 15 13 0 13 3 1 12 9 1 9 11 2
19 9 11 11 13 10 0 9 0 9 9 3 1 12 9 1 0 9 11 2
21 1 9 9 11 2 11 2 9 13 3 1 0 9 0 9 0 0 7 0 9 2
28 3 9 1 0 9 3 13 1 9 9 2 15 1 10 9 13 12 1 9 1 0 9 0 9 1 0 9 2
24 1 12 9 1 12 9 9 3 1 9 0 9 9 9 14 1 9 13 10 0 7 0 9 2
3 2 11 2
4 9 11 0 11
4 2 11 2 2
25 1 12 9 0 7 0 9 0 0 2 9 2 11 7 10 0 9 13 0 9 1 0 0 9 2
24 1 9 0 9 9 11 11 4 0 9 2 15 15 9 10 0 0 9 13 2 10 9 13 2
29 0 9 11 4 13 13 0 9 1 0 9 16 0 0 11 2 16 0 9 1 11 13 0 16 0 9 9 11 2
18 3 13 11 11 2 9 1 11 13 13 0 9 3 1 0 0 9 2
3 9 1 11
5 11 2 11 2 2
18 9 13 9 0 9 0 9 11 1 9 9 13 1 10 9 9 9 2
18 3 13 9 11 11 2 9 1 0 9 4 15 13 13 7 3 13 2
25 9 9 4 13 4 13 3 2 1 9 2 0 9 11 2 9 9 2 9 9 9 7 0 9 2
19 1 0 9 4 0 9 13 7 1 9 4 9 13 9 0 0 0 9 2
26 1 12 2 9 12 4 1 0 12 9 9 1 9 0 9 13 9 7 4 13 1 0 9 12 9 2
12 0 9 2 1 0 9 0 2 13 12 9 2
2 13 0
2 11 2
25 1 9 0 9 0 9 1 11 2 12 0 11 11 2 2 15 13 12 0 11 11 2 1 11 2
11 16 0 1 0 9 9 4 13 1 9 2
18 13 2 14 15 9 0 2 13 15 9 9 9 1 12 1 12 9 2
6 9 9 9 3 13 2
26 1 9 1 9 1 0 9 13 1 9 12 2 9 3 3 0 9 10 9 2 12 0 9 11 11 2
26 10 0 9 2 0 1 0 9 2 13 9 1 9 9 2 3 13 2 3 1 9 1 12 2 9 2
16 9 0 9 3 13 0 9 2 16 9 9 13 0 0 9 2
2 9 3
5 11 2 11 2 2
28 1 9 0 9 1 0 0 9 1 9 1 12 2 12 2 3 13 1 9 11 7 11 1 9 1 0 9 2
11 13 15 9 12 2 12 2 12 2 12 2
21 1 9 11 2 11 2 11 2 9 9 2 0 2 0 9 4 13 0 0 9 2
25 16 0 13 9 1 0 0 9 13 3 0 9 2 3 3 13 9 1 0 9 7 1 0 9 2
16 1 0 9 15 9 13 1 0 9 2 1 0 15 3 13 2
2 0 9
2 11 2
21 9 0 9 13 0 0 7 0 9 2 11 2 1 12 9 9 9 9 0 9 2
12 4 13 9 9 7 9 1 0 9 7 9 2
15 1 0 9 15 13 13 3 0 9 0 9 2 9 0 2
5 9 1 11 1 9
39 9 0 9 11 11 2 11 2 1 0 11 13 10 0 9 13 1 9 9 0 9 1 9 11 11 2 11 2 2 15 13 1 0 9 9 0 0 9 2
26 1 9 2 15 15 9 11 13 1 9 2 13 9 11 13 12 1 0 9 1 0 9 1 0 11 2
34 0 9 1 10 9 13 13 7 10 9 0 0 9 2 0 0 9 2 15 3 13 1 12 9 9 2 7 10 9 13 3 11 11 2
5 9 1 11 1 9
25 2 13 2 16 1 0 9 13 9 0 9 2 7 13 3 0 9 2 15 15 3 13 1 9 2
9 13 15 9 2 2 13 11 11 2
29 9 0 9 13 1 9 3 0 9 9 11 1 11 2 15 16 0 9 13 1 0 9 0 0 9 1 0 11 2
23 0 9 15 1 9 9 1 10 9 13 2 16 15 1 0 9 3 15 0 13 9 13 2
46 2 0 9 13 0 2 7 3 15 0 9 1 0 11 2 1 15 4 13 1 9 10 9 7 9 10 9 2 11 7 0 9 2 13 7 10 0 9 0 9 2 2 13 9 11 2
23 2 0 0 9 13 9 2 1 9 4 3 13 3 3 2 16 4 15 3 13 10 9 2
29 9 13 2 16 12 1 12 9 9 15 13 1 9 11 1 9 0 11 2 7 1 15 15 10 9 3 13 2 2
34 11 11 13 2 16 15 1 15 1 9 1 10 9 13 3 11 1 0 11 2 3 7 0 9 9 1 9 11 7 3 3 9 11 2
43 16 9 9 1 0 0 9 13 9 11 1 9 3 14 3 2 16 0 9 13 1 0 7 0 9 2 13 15 1 0 9 0 9 1 11 2 15 4 13 0 9 13 2
8 9 1 9 11 2 11 2 2
10 9 12 9 9 13 0 9 1 11 2
20 1 9 13 9 10 9 2 13 9 2 9 2 13 1 9 2 13 0 9 2
7 1 0 9 9 15 13 2
15 1 0 9 10 9 13 9 1 9 9 3 1 12 9 2
17 9 13 12 9 2 9 0 12 9 2 12 9 15 13 15 9 2
20 1 0 9 2 3 15 9 13 1 0 0 9 2 4 0 3 13 10 9 2
14 14 1 0 9 7 9 13 1 9 9 12 9 9 2
22 0 9 3 13 1 12 2 9 0 0 9 1 9 9 2 9 1 9 9 7 13 2
21 16 9 13 3 3 0 9 2 4 13 13 9 9 2 13 10 9 2 13 9 2
8 9 1 0 9 13 3 0 2
14 0 0 9 4 13 14 12 9 15 9 1 9 9 2
21 9 2 15 4 13 0 9 9 2 7 13 9 0 9 0 10 9 2 3 13 2
16 9 13 3 1 3 0 9 7 3 4 13 9 1 9 9 2
14 9 1 12 9 15 13 1 12 7 12 9 1 9 2
13 0 9 9 1 9 13 1 9 12 7 12 9 2
9 0 9 4 7 13 0 9 9 2
27 0 9 1 9 10 9 2 10 9 7 9 9 15 13 3 1 9 9 2 13 1 10 9 1 9 9 2
8 9 4 3 9 13 3 9 2
8 0 9 9 9 3 13 0 2
15 9 13 13 1 0 9 2 15 4 13 4 12 9 13 2
8 9 9 0 9 9 3 13 2
12 1 9 9 1 9 0 9 7 9 15 13 2
5 9 1 9 0 9
5 11 2 11 2 2
20 9 0 9 4 1 0 9 11 0 9 11 11 13 10 0 0 9 11 11 2
25 9 11 11 0 9 11 13 15 2 16 13 10 9 1 9 1 9 2 15 15 13 0 0 9 2
12 9 13 9 9 9 3 1 9 1 10 9 2
3 11 9 13
10 16 9 13 9 3 2 13 1 0 9
7 11 2 11 2 11 2 2
37 1 9 13 1 11 12 0 9 15 1 9 9 0 9 0 9 0 1 9 9 1 9 0 9 11 11 13 1 9 9 11 7 0 9 11 11 2
21 9 11 13 1 9 0 0 9 1 9 13 3 2 16 4 9 13 1 0 9 2
19 13 15 3 9 1 9 9 3 1 11 2 3 15 15 3 13 9 13 2
19 3 9 9 1 11 11 15 13 2 16 1 12 9 15 13 9 11 13 2
32 11 11 2 9 9 0 2 9 2 11 11 0 15 3 9 7 9 9 2 15 13 2 2 1 9 9 1 11 13 15 0 2
16 1 10 10 7 0 9 4 13 9 7 13 15 7 3 2 2
15 1 9 0 0 9 11 11 3 15 13 3 1 9 9 2
10 2 1 15 0 9 13 3 10 9 2
22 16 15 2 3 13 2 13 3 0 9 11 7 15 0 2 3 13 1 0 9 2 2
2 0 9
2 9 9
3 9 9 9
4 9 12 12 12
4 9 12 12 12
4 9 12 12 12
7 9 2 9 2 12 12 12
6 0 2 9 12 12 12
6 0 2 9 12 12 12
3 2 9 2
3 12 12 12
7 9 2 9 2 12 12 12
4 9 12 12 12
21 13 9 12 2 9 9 2 9 0 12 2 7 12 2 9 2 7 13 10 9 2
10 12 2 0 2 11 2 11 11 12 12
6 12 2 11 2 11 12
6 12 2 11 2 11 12
7 12 2 11 2 11 12 12
7 12 2 11 2 11 11 12
17 12 2 11 11 2 2 0 2 11 12 2 15 12 2 0 9 2
6 12 2 11 2 11 12
6 12 2 11 2 11 12
8 12 2 11 2 0 2 11 12
6 12 2 11 2 11 12
7 12 2 11 2 11 12 12
6 12 2 11 2 11 12
12 12 2 11 2 11 12 2 15 0 0 9 2
4 0 9 0 9
41 2 9 0 9 1 11 15 13 2 16 2 0 2 9 11 13 3 9 1 0 9 1 11 1 0 9 11 2 11 2 16 15 13 1 9 0 9 1 0 9 2
39 1 0 9 15 13 2 16 0 9 13 9 2 1 15 13 7 9 1 9 3 12 9 1 9 2 0 11 2 1 0 0 9 2 2 13 0 9 11 2
25 1 9 1 0 9 9 13 2 16 1 9 0 2 0 9 13 13 0 9 2 0 0 9 2 2
49 1 0 9 2 15 13 4 13 2 0 9 2 3 1 0 9 15 3 13 1 9 9 11 2 7 10 9 1 9 0 9 3 13 2 7 15 15 13 9 9 1 3 3 0 7 0 9 2 2
5 9 13 1 12 9
8 3 1 0 9 9 1 0 11
15 0 9 9 2 0 9 12 9 2 15 1 0 9 13 2
33 9 1 9 15 12 3 0 9 11 2 12 2 1 9 11 2 1 11 2 12 2 2 13 0 9 7 1 9 13 9 0 9 2
40 1 9 15 7 3 13 1 9 1 12 0 9 2 15 3 13 3 11 7 11 2 16 12 13 1 0 2 0 9 13 11 11 1 9 1 0 0 9 11 2
42 9 9 11 11 1 0 9 2 2 13 2 16 0 9 9 13 1 15 2 16 1 9 1 9 4 12 0 9 2 0 0 9 0 9 7 0 9 2 13 10 9 2
30 1 9 9 9 2 11 4 15 7 3 13 2 16 16 9 13 0 9 2 3 9 1 10 9 0 9 13 2 2 2
23 16 15 3 1 9 11 1 0 9 13 3 2 3 4 9 13 9 2 16 15 9 13 2
18 7 15 13 1 15 2 16 9 1 0 9 15 14 10 0 9 13 2
15 2 3 0 2 11 3 1 9 13 1 12 2 9 9 2
10 3 9 13 11 0 0 2 9 0 2
24 2 15 13 2 7 13 3 9 9 2 15 4 13 13 9 13 2 3 15 13 1 0 9 2
17 0 9 13 2 16 0 9 3 0 9 15 13 2 16 15 13 2
24 0 2 16 9 13 1 9 0 9 2 15 13 1 9 1 15 2 1 15 15 13 1 15 2
29 2 13 15 7 13 2 16 16 9 1 9 1 11 13 2 13 15 0 9 9 7 13 15 10 9 1 9 13 2
7 7 15 4 13 1 9 2
15 7 3 9 9 10 9 9 2 11 1 10 0 9 13 2
15 9 0 9 13 9 12 9 2 15 13 3 9 9 9 2
10 1 9 9 7 4 13 3 12 9 2
17 11 0 2 2 9 1 10 9 9 13 0 9 1 9 10 9 2
28 13 3 0 9 0 0 9 2 9 9 9 2 9 2 9 2 9 2 9 2 9 9 2 15 10 15 13 2
26 11 7 11 1 15 15 3 13 2 15 13 9 10 0 0 9 11 11 2 1 15 4 12 9 13 2
11 0 9 13 1 9 3 13 11 11 2 2
12 0 11 0 9 2 12 2 11 2 12 2 11
20 1 0 11 1 0 2 0 2 7 3 0 9 15 13 0 9 9 1 9 2
26 7 1 10 9 13 9 3 2 11 2 0 1 9 2 10 0 9 13 2 11 13 14 1 9 11 2
15 1 9 15 7 11 1 0 9 13 9 7 13 1 9 2
22 11 3 0 9 13 9 7 3 15 1 9 1 0 9 13 0 9 2 3 13 0 2
22 1 9 13 3 1 11 1 0 9 7 1 3 16 12 2 7 12 2 9 15 13 2
19 3 11 7 11 13 0 7 0 9 1 0 9 9 2 11 13 1 0 2
67 9 11 2 12 2 11 2 11 2 2 2 12 2 11 2 11 2 2 12 2 11 2 11 2 2 15 11 2 2 12 2 11 2 11 2 2 11 2 2 12 2 11 2 11 2 2 11 2 2 12 2 11 2 11 2 11 2 2 12 2 11 2 11 2 11 2 2
34 0 9 9 2 12 2 11 12 2 12 2 11 12 2 12 2 11 12 2 12 2 11 12 2 12 2 11 12 2 12 2 11 12 2
6 3 12 2 9 0 9
17 9 0 9 11 2 11 13 1 0 12 2 9 0 9 0 9 2
18 11 13 3 13 2 3 1 11 13 0 9 2 15 3 13 7 9 2
13 10 0 0 9 13 1 2 9 2 12 0 11 2
23 2 13 1 15 3 1 10 9 7 9 0 9 1 11 7 11 2 2 13 0 9 11 2
17 9 9 2 3 15 13 11 13 1 0 9 12 2 12 1 11 2
25 2 1 10 0 9 2 3 4 13 15 12 9 2 10 9 13 0 7 13 15 9 1 0 9 2
17 3 0 9 13 3 13 7 13 0 9 2 2 13 9 11 11 2
36 11 1 9 3 13 9 2 15 3 1 11 4 3 13 2 2 13 4 15 0 9 1 11 2 3 4 13 0 9 2 2 13 0 9 11 2
23 1 11 13 2 0 2 11 2 1 9 1 9 0 12 9 1 12 9 2 12 13 11 2
18 9 11 11 2 2 16 4 3 13 2 13 13 1 9 9 1 9 2
6 11 13 9 0 9 2
8 13 9 7 13 1 15 2 2
63 9 0 12 2 9 2 1 12 2 11 2 11 2 9 11 2 2 11 2 11 2 11 2 2 11 2 11 2 11 2 2 11 2 11 2 11 2 2 11 2 11 2 11 2 2 12 2 11 2 0 2 11 2 9 2 2 11 2 11 2 11 2 2
23 9 11 7 11 11 11 2 3 2 7 11 11 13 10 9 1 11 0 9 2 9 9 13
2 0 9
10 9 11 13 13 13 10 9 1 11 11
42 2 13 13 1 9 9 2 15 13 7 13 2 16 4 13 9 1 9 2 1 15 13 1 10 12 9 2 2 13 1 9 1 11 3 9 0 9 9 11 11 11 2
19 13 15 1 0 9 10 9 2 9 9 11 11 1 9 11 11 0 11 2
24 11 13 1 11 9 2 15 4 13 1 9 1 11 7 0 2 9 13 14 9 12 0 9 2
27 2 14 1 12 9 0 9 11 7 1 12 9 9 11 11 2 11 4 13 10 9 2 2 13 9 11 2
34 2 13 4 1 15 2 16 11 13 1 11 0 9 7 13 9 1 9 1 9 1 11 14 1 9 2 16 4 13 9 1 9 9 2
18 7 16 11 13 15 9 2 16 4 7 13 9 2 7 9 3 2 2
18 1 10 9 15 11 13 2 3 13 10 9 2 9 0 9 11 11 2
23 2 9 11 13 11 2 16 4 13 9 2 1 15 13 3 13 2 16 11 13 10 9 2
15 16 15 13 2 13 15 0 9 2 3 13 10 9 13 2
35 11 13 2 16 11 9 13 13 2 7 9 11 15 13 2 16 13 9 2 7 1 10 9 7 9 9 11 13 11 1 9 10 9 2 2
28 9 11 13 0 9 1 0 9 11 1 9 2 3 4 13 2 16 4 13 9 1 0 9 11 11 1 11 2
32 2 11 13 0 15 9 9 1 11 13 2 7 3 11 13 9 11 1 11 2 3 4 15 1 9 13 2 2 13 9 11 2
21 13 2 16 11 11 1 10 9 13 10 9 1 9 7 13 13 11 1 12 9 2
11 13 15 7 13 2 16 11 13 1 9 2
29 2 15 10 9 13 1 10 9 9 2 16 13 13 10 9 1 9 11 7 10 9 9 11 2 2 13 9 11 2
9 0 0 9 9 11 13 0 9 2
37 2 13 15 1 15 2 16 1 0 9 9 11 13 0 0 9 1 9 9 2 13 10 9 2 13 1 0 9 2 0 9 2 2 13 0 9 2
16 2 9 9 11 15 3 13 0 9 2 7 13 15 14 9 2
15 13 3 10 9 2 15 4 13 9 11 15 10 9 13 2
12 16 15 13 2 13 15 1 15 9 9 2 2
20 9 11 13 2 16 13 1 9 9 1 11 7 10 9 2 15 0 9 13 2
19 2 13 4 1 0 9 7 15 15 13 2 15 13 1 10 9 0 2 2
20 1 9 2 3 15 13 11 11 2 9 11 13 2 2 11 13 1 15 0 2
20 1 0 9 15 13 9 1 12 9 2 7 3 4 0 1 11 13 2 2 2
14 13 15 2 16 1 9 9 1 11 4 15 15 13 2
3 2 14 2
19 7 16 13 11 0 9 2 12 9 12 9 9 13 12 9 12 9 9 2
7 1 0 9 15 13 2 2
17 11 13 13 3 11 2 7 9 11 2 15 13 0 1 9 9 2
17 2 15 15 3 13 2 13 9 10 0 9 2 2 13 9 11 2
22 2 1 11 1 9 9 1 12 9 13 0 1 12 9 2 15 13 1 0 9 2 2
4 13 15 9 9
7 0 9 11 2 3 9 2
8 16 9 2 3 1 12 9 2
14 2 13 3 1 9 2 3 13 3 0 9 13 2 2
34 15 13 11 11 2 0 9 0 2 9 0 7 0 9 2 11 2 1 10 9 1 9 1 9 12 2 15 3 3 13 0 9 11 2
9 2 1 3 13 9 9 0 9 2
6 2 1 9 10 9 2
16 9 3 13 9 1 9 11 2 3 3 1 9 9 2 2 2
8 1 10 9 15 9 9 13 2
11 2 15 1 15 15 13 3 13 10 9 2
8 3 15 7 13 13 9 9 2
48 7 16 1 10 9 9 13 7 3 2 4 13 1 15 2 16 0 9 4 13 1 10 0 9 1 11 3 9 2 7 1 1 10 0 0 9 4 13 9 7 1 9 3 1 9 2 2 2
10 7 11 16 9 4 1 10 13 9 2
14 2 10 9 1 11 13 13 1 9 9 12 2 2 2
23 4 15 9 9 13 9 12 2 12 2 3 3 2 3 13 15 13 1 0 7 0 9 2
22 2 7 1 9 15 4 1 15 9 13 12 2 12 7 3 15 13 3 1 10 9 2
13 7 9 15 4 13 9 1 10 0 9 2 2 2
14 3 13 13 0 9 2 3 0 0 9 2 3 11 2
22 2 13 2 16 4 9 13 1 9 10 9 2 3 15 13 2 3 1 9 0 9 2
26 9 13 1 11 10 9 2 16 15 9 2 0 3 1 0 9 2 4 3 13 1 0 9 2 2 2
8 10 13 0 9 1 9 9 2
20 2 13 15 3 13 9 1 9 2 9 2 9 2 9 7 10 9 7 9 2
10 7 3 3 3 0 0 9 2 2 2
8 10 9 13 9 9 1 9 2
22 2 15 2 15 1 9 13 2 15 13 14 12 9 2 7 3 7 15 9 0 9 2
31 16 7 15 1 9 2 15 9 13 2 13 1 0 9 2 13 10 9 2 16 4 15 1 0 9 13 13 16 0 15 2
15 10 15 7 3 13 1 0 9 2 15 13 13 2 2 2
11 10 13 1 15 9 9 11 1 10 9 2
8 2 1 9 9 13 1 9 2
16 1 0 9 13 9 9 2 15 13 0 13 10 9 1 9 2
24 13 3 3 1 0 9 1 0 7 0 9 1 0 9 2 16 4 15 0 9 13 2 2 2
17 4 13 0 9 0 9 16 0 9 0 9 9 13 1 0 9 2
24 2 13 13 10 9 2 9 9 9 2 3 3 14 0 7 0 9 2 13 1 0 0 9 2
27 13 7 2 16 13 9 7 16 15 9 9 15 4 13 1 0 9 2 15 13 3 9 0 9 2 2 2
6 13 15 13 9 9 2
26 2 15 4 3 13 2 7 14 0 9 13 9 1 12 9 2 16 1 0 9 15 13 1 12 9 2
7 7 14 13 1 9 9 2
10 13 7 13 2 16 1 9 15 13 2
8 1 9 9 13 3 1 9 2
3 7 9 2
11 3 2 3 14 2 7 1 12 9 2 2
5 0 9 2 11 13
8 11 15 1 11 13 9 1 11
25 14 1 0 9 2 7 3 3 1 9 15 10 0 9 13 3 1 10 0 0 9 1 0 9 2
33 11 3 13 1 9 3 1 11 2 3 15 13 1 11 7 3 3 1 10 9 13 3 0 9 11 2 11 2 11 1 9 9 2
64 1 0 9 11 4 13 12 9 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 2 0 2 11 2 15 13 1 9 1 11 2 0 12 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 1 0 9 11 2 11 13 1 11 2
7 0 9 13 1 0 11 2
41 1 9 13 9 11 2 15 9 11 9 2 11 7 9 11 13 2 16 10 0 9 1 0 9 1 11 15 1 0 9 13 0 9 2 4 1 15 13 11 2 2
36 11 11 3 13 9 9 11 2 9 0 9 2 2 3 13 2 16 11 13 10 0 9 2 7 1 3 0 0 9 3 13 9 15 13 2 2
35 0 11 13 1 9 9 1 10 9 2 0 13 9 11 2 12 9 2 12 5 1 9 2 2 0 9 9 11 2 15 13 9 0 11 2
42 1 15 12 13 1 9 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 7 11 2
19 2 1 0 9 15 13 9 2 7 13 1 12 0 9 9 12 2 12 2
18 7 13 2 16 3 3 3 9 13 2 2 13 15 3 13 9 11 2
18 3 7 13 3 10 11 2 2 3 13 0 9 2 16 4 15 13 2
9 13 2 16 1 10 9 15 13 2
29 13 15 1 15 2 16 15 13 2 16 13 9 12 2 12 2 16 13 13 3 9 7 3 3 15 13 3 2 2
16 11 2 2 11 13 9 2 16 1 10 9 0 9 3 13 2
20 13 15 2 16 1 9 11 3 13 1 0 9 7 13 13 13 3 0 9 2
9 7 15 13 2 16 3 13 2 2
18 9 9 11 11 2 2 1 0 9 4 3 1 11 13 2 13 0 2
15 7 3 15 1 11 3 13 0 9 2 13 2 16 13 2
18 7 11 15 3 13 3 13 2 3 10 9 2 9 7 9 13 9 2
6 13 13 1 15 2 2
3 11 3 13
38 0 12 9 0 9 9 11 2 11 2 11 1 11 1 11 13 12 9 11 11 2 12 2 11 2 12 2 11 2 2 9 7 13 3 1 9 11 2
26 0 9 11 13 1 9 0 14 12 2 12 9 2 1 11 2 7 13 15 3 9 1 9 0 9 2
37 3 10 0 9 11 11 2 11 11 2 13 13 12 9 1 9 0 9 1 0 9 2 1 9 13 3 16 9 7 3 13 14 1 12 2 9 2
26 1 0 11 13 3 11 0 9 12 2 12 2 12 9 2 1 0 11 3 12 2 12 2 12 9 2
29 1 9 13 1 0 9 0 11 2 3 7 3 13 11 1 12 2 12 9 2 1 11 2 12 11 11 12 2 2
55 1 9 9 15 3 13 0 9 11 2 12 2 11 2 12 2 11 2 2 11 1 11 12 12 5 12 13 1 9 0 1 9 12 2 12 9 2 1 9 2 11 1 0 9 12 13 0 2 12 2 12 9 2 2 2
20 1 9 13 0 0 12 9 0 9 1 0 9 2 12 9 2 1 9 11 2
5 9 9 1 11 2
76 11 2 11 2 2 11 2 12 2 12 2 12 9 2 12 2 11 2 11 2 11 2 12 2 12 2 12 9 2 12 2 11 2 11 2 2 11 2 12 2 12 2 12 9 2 12 2 11 2 11 2 11 2 12 2 12 2 12 9 2 12 2 11 2 11 2 2 11 2 12 2 12 2 12 9 2
9 11 1 11 1 0 9 1 9 2
8 1 9 1 11 13 14 11 2
5 9 13 2 9 13
4 0 9 1 11
41 2 9 0 9 1 11 15 13 2 16 2 0 2 9 11 13 3 9 1 0 9 1 11 1 0 9 11 2 11 2 16 15 13 1 9 0 9 1 0 9 2
28 0 9 13 9 2 1 15 13 7 0 9 1 9 2 0 11 2 1 0 0 9 2 2 13 0 9 11 2
16 1 9 0 2 0 9 13 13 0 9 2 0 0 9 2 2
12 1 9 1 9 11 15 13 7 1 0 9 2
13 3 9 9 11 11 13 9 1 3 0 7 0 2
17 1 9 0 9 13 2 16 13 9 2 16 4 13 9 9 9 2
23 3 13 2 16 2 0 0 9 2 1 15 1 11 13 2 15 4 13 1 0 9 2 2
30 9 0 9 2 15 15 13 9 7 13 2 16 9 1 9 9 1 9 13 9 1 9 11 11 2 13 9 1 9 2
26 0 13 7 0 9 1 11 1 9 9 12 2 9 2 10 9 13 13 2 0 0 9 1 11 2 2
12 4 15 3 13 0 9 11 9 0 9 11 2
20 2 13 10 9 9 7 13 15 1 0 9 0 9 2 2 13 15 1 9 2
14 2 1 0 9 2 15 13 1 9 2 4 13 9 2
19 4 13 2 7 9 10 9 2 3 1 12 9 2 2 13 3 1 9 2
36 1 9 9 13 2 16 4 9 11 13 1 0 9 1 11 2 16 15 13 9 14 0 9 9 12 2 9 2 7 0 9 1 15 13 9 2
2 1 9
18 9 9 2 12 2 11 12 2 12 2 11 12 2 12 2 11 12 2
18 11 11 2 11 2 7 11 11 2 11 2 13 1 12 9 9 9 2
17 11 11 2 0 0 2 0 9 2 9 11 12 2 13 3 9 2
2 13 2
2 9 9
8 0 2 11 2 11 2 2 2
40 0 2 0 9 1 9 9 1 9 2 11 2 12 2 12 2 11 2 12 2 3 2 2 9 1 12 9 2 12 2 11 2 11 2 2 2 12 2 11 2
1 9
2 11 2
45 9 11 2 12 2 11 2 12 2 11 2 12 2 11 2 12 2 11 2 12 2 11 2 12 2 11 2 12 2 11 2 11 2 11 2 2 2 12 2 11 2 12 2 11 2
77 9 11 2 12 2 11 2 12 2 11 2 12 2 11 2 12 2 11 2 12 2 11 2 12 2 11 2 12 2 11 2 12 2 11 2 12 2 11 2 12 2 11 2 2 2 12 2 11 2 12 2 11 2 12 2 11 2 12 2 11 2 12 2 11 2 12 2 11 2 12 2 11 2 12 2 11 2
2 11 2
57 9 12 2 9 9 11 11 2 12 9 2 9 11 2 2 11 2 11 11 2 12 2 12 2 12 2 12 2 12 2 12 2 11 2 12 9 2 9 11 2 2 11 2 11 2 12 2 12 2 12 2 12 2 12 2 12 2
2 11 2
16 9 9 9 11 2 11 2 11 12 2 12 2 12 2 12 2
3 0 11 2
21 1 9 11 4 13 2 16 9 9 9 15 4 13 1 9 12 9 0 0 9 2
3 3 0 9
5 15 15 1 15 13
3 3 0 9
24 9 9 11 13 9 1 0 9 1 9 1 11 15 2 1 9 11 15 11 1 10 9 13 2
14 7 13 7 0 2 16 9 9 13 11 10 0 9 2
12 1 3 0 9 7 13 9 1 9 0 9 2
8 15 15 15 3 1 9 13 2
31 9 11 9 11 15 13 2 16 15 15 13 0 2 7 16 13 3 1 9 1 9 2 16 4 0 0 9 10 9 13 2
13 13 7 10 10 9 2 15 3 1 0 9 13 2
25 13 1 10 0 9 2 15 15 13 13 1 10 9 1 9 1 0 0 9 7 13 11 0 9 2
17 6 2 9 11 13 0 7 15 1 15 13 3 1 15 3 9 2
15 1 9 13 7 3 7 11 11 2 9 3 2 0 2 2
16 15 3 13 13 2 16 4 15 10 2 9 2 1 9 13 2
4 7 3 13 2
2 1 9
42 11 1 11 2 12 9 2 2 1 11 11 13 0 9 9 1 9 1 11 2 12 2 11 2 11 2 9 11 2 12 2 12 2 11 2 9 2 11 2 2 12 2
41 0 2 0 9 2 9 2 11 2 11 11 12 2 12 2 9 11 2 11 11 12 2 12 2 0 11 2 11 11 12 2 12 2 11 11 2 11 12 2 12 2
23 1 9 2 12 2 7 12 2 12 2 2 15 13 2 11 2 11 2 0 11 2 11 2
8 9 3 0 9 13 1 11 2
65 1 9 2 0 9 9 2 1 12 2 9 2 11 2 11 12 2 12 2 9 2 9 2 12 2 11 2 11 2 12 2 2 2 12 2 11 12 9 2 9 2 11 2 11 12 2 12 2 12 2 12 2 2 11 2 11 12 2 12 2 12 2 12 2 2
6 0 2 9 13 13 2
57 9 9 1 9 0 9 1 11 2 12 9 2 2 12 2 11 2 11 2 11 2 14 2 11 2 12 2 12 2 12 2 12 2 11 12 2 12 2 11 12 2 12 2 11 2 11 2 11 2 11 2 9 2 12 2 12 2
21 11 2 0 11 12 2 12 2 1 9 1 0 9 11 7 11 1 9 0 9 2
5 13 0 2 11 2
27 9 9 11 13 9 1 9 0 9 1 9 9 11 2 11 7 13 0 9 1 0 0 9 1 0 9 2
23 0 9 3 2 11 2 9 11 2 12 2 11 2 2 0 2 11 2 11 2 12 2 2
25 0 9 11 11 15 3 1 0 9 2 1 12 2 1 12 2 2 12 2 9 1 9 13 9 2
4 1 11 3 11
64 1 12 2 9 2 12 1 12 0 9 2 0 9 13 3 9 11 2 11 2 11 2 2 12 2 12 2 12 9 2 12 2 11 2 11 2 11 2 2 15 11 9 2 12 2 12 9 2 12 2 11 2 11 2 11 2 2 11 11 2 12 2 12 2
5 11 0 1 0 11
16 1 0 11 2 1 0 9 9 2 15 1 10 9 9 13 2
18 1 9 11 13 2 7 9 9 13 9 2 9 13 7 11 7 11 2
17 1 9 13 1 0 9 7 13 3 14 12 2 7 12 2 9 2
14 3 11 7 11 13 0 7 0 9 1 0 9 9 2
69 9 1 11 2 12 2 11 2 11 2 2 2 12 2 11 2 11 2 2 2 12 2 11 2 11 2 2 15 11 2 2 12 2 11 2 11 2 2 11 2 2 12 2 11 2 11 2 2 11 2 2 12 2 11 2 11 2 11 2 2 12 2 11 2 11 2 11 2 2
34 0 9 9 2 12 2 11 12 2 12 2 11 12 2 12 2 11 12 2 12 2 11 12 2 12 2 11 12 2 12 2 11 12 2
4 11 1 0 11
5 9 11 13 0 9
26 11 11 2 0 2 0 9 2 3 9 11 7 11 1 11 2 4 13 1 0 0 11 1 0 11 2
53 9 10 9 11 11 2 9 0 9 1 11 12 2 15 13 1 9 2 1 15 13 7 9 2 16 3 11 1 9 3 4 3 1 11 0 13 2 16 3 13 10 9 2 0 9 11 2 11 2 11 2 3 2
31 2 7 3 4 15 1 11 13 7 13 4 15 2 16 16 15 13 1 11 2 3 13 9 16 9 11 2 16 15 13 2
9 7 1 15 13 1 9 1 11 2
10 11 15 13 2 16 1 9 13 13 2
16 4 13 1 9 0 1 0 9 2 10 0 9 1 15 13 2
34 13 15 2 16 3 4 13 13 16 9 1 11 7 11 1 12 9 2 7 3 16 15 9 1 15 16 0 13 2 2 13 0 9 2
5 11 3 2 13 2
19 0 9 11 13 10 0 9 2 15 13 1 0 9 11 2 3 9 11 2
22 13 3 3 1 0 9 9 2 13 1 0 9 9 9 0 2 9 2 11 11 11 2
20 1 9 1 11 13 3 14 12 9 15 0 9 2 1 15 13 7 9 9 2
11 3 1 9 15 13 12 9 1 9 9 2
36 11 2 2 0 9 12 9 13 3 3 2 16 4 1 15 0 13 9 2 15 13 1 9 2 7 16 4 13 9 1 0 9 1 9 2 2
18 11 1 0 12 7 9 9 9 3 2 13 2 1 0 0 0 0 2
16 7 9 0 9 1 9 7 10 9 9 9 1 11 13 0 2
11 3 11 16 0 0 9 11 9 11 13 2
3 13 4 15
4 13 9 16 9
22 9 9 11 1 9 2 9 2 9 2 9 2 13 11 11 2 12 2 1 9 11 2
24 15 13 1 0 9 9 2 7 1 9 9 1 9 13 1 1 9 7 9 3 13 16 9 2
25 10 9 15 7 13 9 1 0 9 2 0 9 13 1 0 11 7 3 1 11 13 9 12 9 2
10 1 0 9 13 13 1 11 0 9 2
23 3 0 9 13 0 1 9 11 11 2 12 2 2 15 13 1 9 16 9 1 0 9 2
14 9 9 1 9 1 9 13 1 15 2 16 13 9 2
3 0 0 9
33 11 2 0 9 0 0 9 9 9 2 7 3 3 11 1 11 13 9 12 0 2 7 3 0 9 0 0 9 11 11 11 11 2
18 0 9 1 11 1 0 9 13 1 3 0 13 1 9 9 0 9 2
22 0 9 4 1 9 10 9 11 9 2 11 11 13 1 0 7 1 9 9 11 11 2
22 9 2 11 15 13 1 0 9 13 2 16 4 15 1 3 0 9 3 13 3 13 2
5 11 1 11 3 0
17 1 0 9 7 12 9 0 9 13 3 11 11 2 11 9 2 2
31 1 0 9 15 13 1 11 11 2 11 9 2 12 2 12 9 2 2 11 11 2 11 11 2 12 2 12 9 2 2 2
1 3
3 9 13 11
15 0 9 11 11 13 3 3 11 11 0 9 1 11 11 2
14 1 9 1 10 9 13 9 9 0 9 11 11 11 2
27 1 9 9 0 1 9 0 9 13 1 0 9 1 11 2 9 11 1 11 2 0 9 2 0 9 9 2
13 1 9 9 1 10 0 9 1 9 0 9 13 2
5 0 9 1 9 9
2 11 2
26 0 9 13 0 9 2 16 15 0 9 13 0 9 2 13 3 1 10 9 1 11 0 9 11 11 2
47 3 13 2 0 0 9 2 15 1 0 9 1 11 13 2 13 9 15 2 16 0 9 1 9 12 9 13 13 1 0 9 0 9 1 9 2 16 0 9 1 0 9 11 13 3 0 2
21 0 9 1 11 1 10 9 1 10 0 0 9 0 2 9 2 15 1 9 13 2
13 1 10 9 3 13 9 9 1 10 9 1 9 2
26 16 9 0 9 13 1 0 9 2 3 2 1 9 0 9 9 9 2 9 0 0 9 13 15 9 2
14 9 13 2 15 3 0 9 11 4 1 9 9 13 2
5 2 14 2 0 11
2 11 2
33 9 9 0 9 11 3 13 9 9 0 9 2 13 3 0 9 0 9 11 11 16 9 1 0 9 9 9 7 9 11 11 11 2
33 15 13 2 16 0 9 9 0 9 11 13 2 16 9 2 3 11 4 13 1 9 1 0 9 2 4 1 15 13 13 11 11 2
36 9 11 13 1 0 9 9 11 2 1 15 15 9 1 0 9 1 9 0 9 1 11 3 13 2 15 4 13 14 1 0 0 7 0 9 2
2 0 9
31 1 11 2 11 15 15 13 13 1 11 0 9 2 16 0 9 13 3 1 15 3 2 13 3 1 11 9 11 11 11 2
57 10 9 1 15 3 13 2 16 15 11 2 11 16 0 9 3 13 1 12 9 2 2 13 3 0 9 2 16 13 1 9 9 1 11 7 11 7 9 0 9 0 11 1 11 2 7 15 3 13 0 2 2 13 11 2 11 2
8 0 9 0 9 15 13 11 2
18 9 11 11 11 13 2 16 11 13 9 9 1 9 1 9 0 9 2
37 9 0 9 9 0 13 11 11 2 15 13 9 1 10 9 1 9 9 0 9 2 16 4 3 13 9 1 9 11 11 2 11 1 9 9 11 2
37 9 0 9 9 0 3 13 1 9 1 0 9 3 0 9 2 15 13 11 9 7 15 15 13 1 9 11 2 11 2 11 1 9 0 2 9 2
13 13 0 2 16 4 15 13 1 9 9 9 9 2
35 1 9 9 0 9 11 11 2 11 2 15 1 15 3 13 9 9 1 0 11 2 0 0 9 2 11 2 7 3 0 9 2 11 2 2
6 9 13 2 0 9 2
9 9 11 11 2 11 2 1 0 9
15 1 0 9 13 9 11 1 9 9 0 9 1 0 9 2
7 15 13 1 10 0 9 2
10 2 0 9 9 13 9 0 9 9 2
17 0 9 13 3 0 9 2 0 9 9 13 15 3 7 3 13 2
5 2 1 15 3 2
15 2 9 13 9 13 9 2 1 0 9 13 13 10 9 2
17 16 9 13 0 9 3 1 9 2 9 7 9 13 10 0 9 2
24 9 13 0 9 13 3 9 2 7 3 1 9 9 2 0 9 13 1 9 1 15 0 9 2
18 9 4 1 10 9 3 13 9 7 1 0 9 2 15 12 4 13 2
15 10 9 2 0 1 9 0 9 2 13 3 1 0 9 2
13 9 13 2 16 13 3 13 7 0 9 0 9 2
6 15 0 9 13 2 2
3 9 9 12
5 11 2 11 2 2
18 9 9 9 2 11 12 1 0 9 13 12 0 9 11 11 1 11 2
13 0 9 15 13 3 0 9 11 11 1 0 11 2
18 1 0 0 9 4 1 9 1 9 10 9 13 1 0 9 3 3 2
30 1 9 0 9 13 12 0 9 7 0 9 0 9 13 1 9 10 0 9 2 9 2 7 7 0 9 7 3 9 2
30 3 4 13 0 9 1 9 9 9 11 2 15 15 1 0 9 12 9 13 12 0 11 11 1 0 11 2 9 9 2
1 9
3 9 13 2
30 9 1 9 9 12 9 13 1 9 1 9 1 9 0 9 1 11 13 10 0 9 12 0 9 1 9 11 2 9 2
12 0 9 15 13 7 1 9 4 13 1 9 2
3 0 9 2
17 9 9 1 9 12 9 13 1 9 11 1 11 13 12 0 11 2
12 13 2 16 9 13 1 10 9 2 0 9 2
3 9 9 2
12 1 12 0 9 13 1 9 9 1 0 11 2
24 1 11 15 13 9 11 11 9 1 9 12 9 2 1 11 1 0 9 11 11 1 12 9 2
15 0 9 2 12 13 0 9 9 11 12 0 1 0 9 2
1 9
3 9 1 9
33 3 3 13 0 9 0 9 16 0 9 1 15 2 3 13 7 3 13 4 13 9 2 9 2 9 2 15 2 15 13 9 9 2
39 3 7 4 11 13 0 9 0 9 2 15 1 0 13 10 9 2 3 2 9 0 9 1 0 9 7 0 9 2 13 1 0 9 1 0 9 7 9 2
47 11 11 2 9 1 10 0 9 2 10 9 1 0 9 13 2 16 2 9 7 9 12 9 2 3 0 2 13 13 9 0 9 0 0 9 2 7 16 0 9 4 3 3 13 0 9 2
16 1 0 9 13 1 10 9 0 12 9 2 0 2 0 9 2
25 9 13 9 0 9 2 1 15 2 3 2 10 9 13 1 9 1 12 9 3 16 9 1 9 2
33 3 3 13 1 9 11 2 16 13 2 16 4 15 2 15 4 16 0 9 13 1 0 9 10 9 2 13 1 15 3 0 9 2
3 9 13 9
8 0 9 2 13 2 12 9 9
5 11 2 11 2 2
22 0 0 0 9 1 9 0 9 2 9 1 9 2 9 2 9 7 9 13 0 9 2
30 3 15 3 13 9 11 2 11 1 0 9 2 9 12 9 13 1 9 3 9 0 9 1 0 9 14 12 9 9 2
28 9 13 9 7 9 12 0 9 15 13 1 9 2 3 1 0 11 2 2 12 9 3 13 7 13 1 11 2
20 0 9 7 9 1 0 9 9 1 9 13 3 3 2 16 9 13 14 9 2
24 1 0 2 0 7 0 11 15 3 13 1 9 2 9 7 9 7 1 11 13 9 1 9 2
9 9 13 3 0 1 9 1 9 2
15 1 9 9 13 12 9 2 12 9 7 0 0 9 9 2
13 9 9 2 15 13 1 0 9 2 13 3 13 2
12 0 9 9 7 9 4 13 9 13 9 9 2
7 9 9 11 2 11 2 2
49 0 9 2 9 1 9 2 9 0 9 1 11 7 11 2 9 11 1 9 1 0 9 2 9 1 9 7 9 1 0 9 7 0 2 9 1 0 9 13 3 1 11 9 0 11 7 0 9 2
17 1 12 9 2 15 13 13 9 2 13 9 9 7 9 1 9 2
13 12 0 15 3 13 1 0 9 0 9 9 0 2
25 2 1 0 9 13 1 9 16 0 2 9 12 10 9 2 2 13 15 11 11 2 9 9 11 2
17 2 1 0 11 13 9 3 0 9 2 0 9 13 7 1 11 2
9 3 13 9 1 9 1 11 2 2
1 9
3 13 0 2
12 0 9 0 9 15 13 12 0 9 1 11 2
19 3 1 9 15 1 9 1 11 13 9 11 12 7 3 15 1 11 13 2
14 9 2 9 2 9 7 0 9 0 1 11 15 13 2
6 9 13 9 1 11 2
9 1 9 13 0 9 9 1 11 2
6 9 13 2 0 9 2
7 3 4 10 9 13 13 2
41 2 13 4 3 9 2 16 0 9 13 3 9 0 9 2 7 14 9 9 0 9 2 9 9 13 3 3 1 9 2 3 4 9 13 2 7 3 4 13 0 2
35 9 4 13 7 9 0 9 2 10 9 4 15 13 14 1 0 9 2 7 7 1 9 0 9 7 3 2 3 13 13 0 13 0 9 2
11 2 0 13 7 9 1 0 9 7 9 2
5 15 13 10 9 2
22 2 1 9 9 0 9 4 13 0 9 13 12 9 2 15 4 15 13 1 0 9 2
27 9 9 4 13 13 13 7 0 9 2 13 2 16 15 1 0 9 9 13 2 13 15 10 0 9 2 2
17 0 9 0 9 13 7 9 0 0 9 1 9 0 9 2 2 2
17 2 9 3 13 1 9 2 16 9 7 0 9 4 13 13 0 2
16 1 9 4 15 7 13 2 16 15 13 13 1 0 0 9 2
20 15 15 13 13 0 0 9 2 3 1 0 9 13 0 9 1 9 0 9 2
21 1 15 13 1 15 3 3 0 9 13 2 1 0 9 0 9 1 9 0 9 2
21 3 1 9 0 0 9 4 1 10 9 13 13 7 12 9 2 15 0 9 13 2
16 1 0 9 13 3 0 2 16 0 9 10 9 9 3 13 2
15 2 0 9 1 9 9 13 1 9 1 0 7 0 9 2
11 3 4 15 1 15 10 9 13 3 13 2
20 2 1 9 0 9 4 15 10 9 13 13 9 11 11 11 1 9 11 11 2
19 3 3 3 15 9 0 9 1 9 13 2 7 13 15 10 9 3 13 2
11 13 9 2 16 13 2 0 9 9 2 2
13 0 9 4 7 13 0 9 13 1 0 9 2 2
2 9 3
7 11 1 11 2 11 2 2
22 9 9 1 0 9 7 0 9 1 11 1 0 9 15 13 1 0 9 3 1 9 2
21 1 9 9 3 0 0 9 13 7 12 0 9 7 1 9 4 13 7 0 9 2
9 1 0 9 13 9 9 0 9 2
23 16 15 10 0 9 13 2 13 4 4 13 14 1 11 7 3 7 1 9 1 0 11 2
4 15 13 0 9
8 1 9 9 1 9 13 9 9
41 1 9 9 0 9 7 9 0 9 11 11 7 11 11 1 12 2 9 1 9 9 1 0 9 13 12 9 3 13 9 9 11 12 2 12 1 9 9 7 9 2
9 9 15 13 3 9 12 7 12 2
29 9 0 9 13 0 9 0 9 0 9 2 7 13 2 16 4 1 0 9 0 9 13 9 9 9 9 0 9 2
50 2 16 9 11 1 9 13 2 13 15 3 13 9 9 1 9 0 9 11 7 10 9 2 15 1 0 13 1 9 0 9 9 2 1 9 0 0 9 1 0 2 7 7 1 9 3 0 0 9 2
39 13 7 1 9 2 9 1 9 9 2 16 0 2 1 11 3 3 13 14 0 9 9 9 9 1 9 10 9 2 2 13 9 0 9 1 9 9 9 2
28 13 2 16 9 0 9 2 1 10 9 9 9 7 13 2 15 13 3 1 0 11 2 1 11 7 1 11 2
23 1 9 9 0 9 11 1 11 11 11 15 9 13 1 9 1 9 9 7 9 0 9 2
26 2 0 9 13 0 9 0 9 7 1 9 9 13 1 9 13 0 9 2 10 9 0 9 3 13 2
20 1 10 9 15 13 3 1 1 0 9 0 9 1 0 2 7 0 9 11 2
16 3 1 0 9 9 11 13 0 9 11 0 9 1 9 11 2
8 9 9 13 13 10 0 9 2
21 9 0 9 10 9 13 0 12 9 9 0 9 7 13 4 15 0 9 9 2 2
22 2 10 0 9 1 0 9 13 9 1 9 0 9 1 9 0 9 1 9 9 11 2
34 16 0 9 13 9 13 1 10 9 2 13 1 15 3 0 9 12 2 9 2 2 13 15 11 11 1 0 9 0 9 1 9 9 2
23 2 1 9 1 9 9 1 0 9 4 13 1 0 9 7 13 15 1 0 7 3 0 2
6 13 14 1 9 9 2
8 0 9 3 13 9 0 9 2
40 13 7 7 0 2 16 4 9 0 9 1 10 9 13 2 15 15 13 2 1 9 9 15 13 9 7 3 15 15 13 2 2 13 15 3 9 9 11 11 2
23 2 7 15 9 13 2 16 9 0 9 4 13 9 0 9 2 13 0 9 7 13 15 2
22 1 9 0 9 11 9 9 9 13 16 9 9 1 9 2 16 0 9 9 13 2 2
9 1 9 1 11 13 14 9 1 9
5 11 2 11 2 2
24 0 9 1 9 11 11 13 1 0 9 0 2 13 3 1 11 9 2 15 13 10 9 13 2
13 13 15 9 9 11 1 9 7 0 9 11 11 2
18 1 0 9 11 2 11 13 2 2 13 0 2 16 9 9 13 0 2
12 13 0 13 0 9 7 13 15 9 13 2 2
29 1 9 9 13 2 2 13 2 16 15 1 12 0 9 0 0 9 13 3 7 13 7 15 2 15 15 15 13 2
15 3 15 13 3 2 16 1 0 9 3 13 15 0 2 2
29 11 11 13 2 16 9 4 15 1 9 7 9 13 2 16 15 13 9 7 16 3 2 15 0 13 9 13 2 2
15 9 1 15 2 16 4 13 7 9 1 9 2 3 13 2
19 3 13 2 13 9 9 1 9 0 14 1 9 2 16 9 0 9 13 2
39 2 13 7 9 2 16 15 12 0 9 3 2 16 4 10 9 13 9 1 9 2 13 9 7 3 13 12 9 7 12 0 9 2 2 13 11 2 11 2
8 9 1 9 11 2 11 2 2
47 1 9 7 9 1 9 13 0 9 9 11 2 11 2 2 12 2 2 15 13 1 9 12 1 0 9 1 12 9 13 0 11 1 0 9 0 11 1 0 11 2 3 4 13 1 9 2
16 13 1 9 1 11 2 11 2 3 16 9 9 11 11 11 2
41 12 1 9 11 2 11 2 2 12 2 2 0 1 11 1 9 16 9 2 13 1 9 1 9 1 0 9 0 9 7 1 9 13 1 0 9 1 11 1 11 2
22 13 15 3 11 2 11 2 2 12 2 1 11 2 15 1 11 11 2 13 9 9 2
3 9 1 9
5 11 2 11 2 2
11 0 9 0 9 15 13 0 9 11 9 2
21 1 9 3 9 13 13 9 0 11 11 12 9 2 11 7 11 11 12 9 11 2
37 12 9 13 3 0 16 0 9 9 1 0 0 9 7 13 9 0 0 9 0 2 9 2 11 0 11 7 0 2 9 2 11 11 2 9 11 2
12 9 9 1 12 9 9 13 12 7 12 9 2
5 0 9 1 9 12
5 11 2 11 2 2
18 1 12 7 12 9 4 11 1 9 0 9 13 13 9 13 0 9 2
12 10 0 9 4 13 3 1 9 9 0 9 2
21 9 13 7 4 13 0 9 11 2 15 13 9 9 11 11 7 11 0 9 11 2
32 1 9 10 9 2 15 13 0 9 2 13 0 9 1 11 9 1 15 2 16 15 9 13 9 0 1 9 0 7 0 9 2
9 14 0 9 13 13 9 9 12 2
3 9 1 9
5 11 2 11 2 2
19 1 9 0 9 11 0 9 9 1 11 13 0 0 9 1 9 12 9 2
19 0 0 9 13 0 9 9 11 2 15 13 9 1 0 0 9 7 9 2
6 9 13 1 12 9 2
12 9 3 13 9 11 0 1 9 1 9 9 2
9 10 9 4 3 13 3 0 9 2
14 0 9 13 1 11 3 9 0 15 1 9 0 9 2
16 1 2 9 2 13 3 11 2 11 2 11 2 11 7 11 2
43 9 11 11 1 0 9 3 3 13 1 9 10 9 2 15 1 10 0 9 13 1 0 9 7 9 0 9 2 9 2 7 3 7 9 2 15 13 3 9 1 0 9 2
6 11 13 13 1 9 11
5 2 9 2 12 2
4 1 11 1 9
6 1 0 9 0 0 9
10 9 11 11 1 0 9 13 3 0 2
20 10 0 11 3 13 10 9 2 15 1 0 9 1 0 9 13 3 15 0 2
4 7 14 3 2
6 0 11 2 0 9 2
4 3 9 13 2
9 13 1 0 9 2 13 0 9 2
25 3 13 15 2 15 4 13 13 2 0 9 7 9 7 9 1 0 9 7 0 9 7 2 2 2
21 13 3 3 2 1 0 9 2 1 15 15 13 13 9 1 9 1 0 7 9 2
13 13 9 2 13 15 2 1 9 15 13 0 9 2
18 13 9 2 9 3 13 1 9 0 7 0 2 9 10 0 9 13 2
3 13 15 2
7 13 1 15 16 2 9 2
15 16 4 15 9 1 15 13 2 16 13 2 13 15 3 2
3 1 9 2
7 10 9 15 13 0 9 2
25 1 0 2 0 0 9 2 15 13 13 1 0 9 2 9 3 1 9 9 2 9 7 13 9 2
9 15 15 7 1 9 13 1 9 2
19 7 3 3 2 9 13 12 2 1 15 3 0 0 9 1 9 0 9 2
29 9 13 9 1 9 1 11 7 11 1 15 3 13 9 10 0 0 9 2 15 13 16 3 1 11 2 7 11 2
7 7 15 13 3 1 9 2
31 1 9 2 13 2 14 0 15 12 7 12 9 13 9 0 9 2 1 0 9 3 0 2 13 13 1 12 2 9 9 2
6 1 9 3 0 9 2
17 7 3 9 1 9 2 11 11 13 16 9 9 1 11 1 9 2
23 2 16 4 15 3 13 7 13 2 13 4 15 3 2 16 4 15 13 1 9 2 2 2
18 9 13 0 9 2 13 15 3 13 2 7 13 2 16 13 3 0 2
12 13 1 9 13 7 3 2 4 13 0 9 2
13 0 9 2 13 4 2 16 3 13 15 1 9 2
13 7 16 15 9 13 2 13 15 13 7 3 2 2
6 3 13 9 1 0 9
3 11 11 2
12 3 2 0 1 0 9 2 1 9 0 0 9
1 9
6 12 9 2 9 2 9
4 12 9 2 9
3 12 9 9
3 12 0 9
4 12 9 1 9
3 12 9 9
3 12 9 9
12 12 1 9 1 9 2 11 11 2 11 11 2
2 12 9
4 12 11 0 9
3 12 10 9
5 12 0 9 1 11
2 12 9
4 12 9 2 9
2 12 11
2 12 9
2 12 11
5 12 9 1 0 9
9 12 0 9 2 9 9 9 9 2
3 12 9 9
5 9 1 12 1 12
4 12 14 1 11
3 12 15 2
3 12 9 11
2 12 11
4 12 9 1 11
8 12 3 12 9 2 12 2 2
9 12 9 7 9 2 2 2 2 2
3 12 9 9
5 12 1 0 0 9
4 12 0 9 11
3 12 0 0
4 12 11 0 11
4 12 9 1 9
2 12 11
4 12 11 2 11
5 12 11 2 0 9
6 12 9 2 12 2 2
3 12 9 9
4 12 9 1 11
4 12 11 0 9
3 12 9 11
4 12 0 9 12
4 9 11 1 9
5 11 2 11 2 2
43 2 11 15 1 0 9 3 13 7 4 13 9 7 0 9 9 2 2 13 0 9 9 11 11 2 11 2 2 16 1 9 0 9 9 11 13 1 9 3 0 9 9 2
30 3 3 11 2 11 13 2 11 4 13 9 9 9 1 9 9 11 2 0 9 9 1 9 7 9 7 0 0 9 2
11 10 9 3 9 11 7 11 1 9 13 2
7 1 10 9 13 9 9 2
21 9 9 11 11 2 11 2 13 2 16 9 13 9 9 1 9 9 1 12 9 2
11 9 7 0 9 13 1 11 3 0 9 2
13 9 1 9 13 1 9 9 1 9 1 9 11 2
4 11 7 0 9
5 11 14 13 0 9
2 11 2
18 11 13 3 0 13 0 9 0 9 1 9 1 9 11 1 9 12 2
9 13 15 3 0 9 0 2 11 2
57 1 15 7 0 9 1 11 2 3 3 13 0 7 0 9 0 9 0 9 1 11 2 11 2 11 7 0 0 2 0 9 2 13 0 13 1 9 0 9 1 0 9 2 16 11 13 1 0 9 0 1 0 9 1 12 9 2
29 9 11 7 11 15 13 1 9 9 1 11 3 0 9 1 0 9 2 15 1 9 0 9 13 9 1 0 9 2
21 0 2 0 9 0 9 15 13 1 9 0 2 11 13 3 1 0 9 1 11 2
3 9 13 9
2 11 2
3 9 13 9
2 11 2
20 0 9 13 9 9 7 0 9 13 10 9 3 2 13 1 9 9 11 11 2
36 13 2 16 10 9 15 13 1 15 9 2 7 13 2 16 4 1 11 13 9 2 3 1 0 9 13 1 9 2 7 7 1 9 0 9 2
35 13 2 16 1 11 13 0 0 9 1 0 7 0 11 2 7 7 1 9 13 13 10 9 7 9 2 15 4 1 10 9 13 13 9 2
25 13 9 2 16 1 0 9 13 13 3 15 2 15 1 0 9 13 3 3 2 3 3 0 9 2
10 11 13 0 9 2 10 9 13 7 0
1 9
10 11 13 0 9 2 10 9 13 7 0
4 13 1 0 9
14 9 1 9 0 0 9 3 13 9 1 9 0 9 2
21 13 9 9 2 13 13 1 10 0 9 2 7 13 1 15 15 2 15 3 13 2
7 3 0 2 7 0 11 2
22 9 0 9 2 0 0 9 1 0 9 7 3 0 9 0 9 9 15 13 11 0 2
33 3 13 9 2 3 13 0 9 2 3 15 13 9 2 3 13 9 0 9 2 3 12 7 9 9 0 0 9 13 1 0 9 2
9 11 15 1 9 13 7 13 15 2
19 1 9 0 9 15 3 13 15 2 15 13 9 2 15 3 13 3 13 2
17 15 3 15 7 11 13 2 15 3 9 2 3 15 13 2 13 2
18 9 1 9 7 9 2 11 2 13 1 0 9 13 9 9 3 0 2
23 7 3 0 0 9 2 15 13 3 11 2 13 9 7 9 3 13 1 0 9 1 11 2
28 1 9 2 7 15 14 1 9 7 9 0 0 7 0 11 2 15 9 15 13 1 0 9 7 10 0 9 2
24 9 2 16 3 3 13 0 7 0 9 0 9 1 0 0 9 2 7 13 9 1 10 9 2
10 1 0 9 0 9 14 1 9 11 2
14 11 16 9 3 3 13 0 9 1 0 7 0 9 2
12 9 0 9 13 7 3 0 16 1 0 9 2
12 13 16 13 2 16 0 9 13 1 15 0 2
19 13 7 7 13 9 2 16 15 4 1 9 3 13 1 0 9 0 9 2
4 9 3 1 15
2 11 2
4 9 3 1 15
2 11 2
26 9 0 0 7 0 9 3 3 13 1 9 11 0 0 0 9 3 2 16 13 9 0 0 0 9 2
21 9 11 0 0 0 9 7 11 0 0 11 0 13 10 9 1 0 7 0 9 2
19 9 9 9 13 2 16 0 9 13 9 9 2 9 0 9 7 9 13 2
4 3 3 1 9
2 11 2
4 3 3 1 9
2 11 2
18 12 9 13 1 9 1 11 9 9 2 1 0 15 3 13 12 9 2
18 1 9 1 9 0 9 2 3 9 2 13 15 7 1 0 9 0 2
14 3 7 13 15 3 3 2 16 15 1 9 13 3 2
25 9 9 4 13 1 9 9 9 11 11 1 0 9 2 15 13 0 9 9 9 7 0 0 9 2
35 16 3 1 0 9 13 9 9 12 7 12 9 2 12 7 12 9 1 9 2 2 13 15 3 1 3 3 2 16 13 9 1 0 9 2
5 11 13 0 9 11
9 9 1 9 9 7 9 1 12 9
2 11 2
21 1 9 9 7 9 1 12 9 13 0 9 1 11 9 9 7 0 9 11 11 2
33 1 9 11 13 2 16 15 2 15 15 13 2 4 13 1 2 9 9 2 2 4 1 15 13 9 2 4 13 7 1 9 13 2
20 9 9 13 9 1 9 3 2 3 15 9 1 9 9 13 7 1 0 9 2
21 1 0 9 15 1 0 9 11 3 13 9 1 9 0 9 11 11 7 10 9 2
11 1 0 9 15 13 1 9 3 10 9 2
9 0 9 13 1 9 11 2 11 2
28 0 9 9 11 11 13 1 12 2 9 0 9 11 13 2 16 4 4 1 0 9 13 0 9 1 9 11 2
16 10 9 4 7 13 3 9 0 9 9 0 9 2 11 2 2
6 13 15 3 9 11 2
17 1 9 0 9 11 13 3 1 0 9 7 0 0 9 11 11 2
10 9 3 10 9 13 16 9 0 9 2
18 0 0 9 13 1 9 2 15 1 10 9 13 0 9 1 9 0 9
4 0 9 1 11
7 1 11 13 13 2 2 2
8 2 10 9 4 13 2 14 2
16 3 13 9 11 0 9 7 13 1 0 9 0 9 0 2 2
14 9 9 11 1 11 2 9 0 1 0 9 10 9 2
10 7 9 12 1 0 9 0 9 3 2
19 0 9 9 1 11 13 0 9 7 0 9 2 7 9 15 13 3 3 2
26 16 9 13 9 1 9 12 9 1 0 0 9 7 3 13 2 16 13 2 16 1 15 11 4 13 2
20 13 15 2 9 13 2 14 2 2 1 11 13 1 10 0 9 7 13 9 2
13 1 0 9 1 11 1 0 9 13 9 3 0 2
30 11 11 2 15 13 1 10 9 9 12 2 16 9 0 9 2 7 0 1 0 9 2 2 13 10 9 1 0 9 2
20 1 0 9 4 13 1 9 2 16 4 11 13 2 14 2 1 9 1 9 2
18 16 10 0 0 9 2 9 9 7 9 0 9 2 4 9 3 13 2
26 11 3 13 10 9 2 13 15 15 2 16 14 1 9 9 2 13 2 9 2 1 9 0 0 9 2
15 13 13 0 2 16 0 9 2 15 15 13 2 4 13 2
9 3 4 13 1 9 13 16 9 2
14 1 9 1 1 11 2 15 1 10 0 9 13 13 2
8 13 9 2 16 15 11 13 2
13 16 0 2 9 13 1 9 11 1 15 13 13 2
23 12 1 10 9 13 0 9 1 9 3 2 2 13 15 0 9 2 15 13 2 2 2 2
20 15 3 13 7 1 11 4 15 3 13 2 16 3 13 1 9 10 0 9 2
9 7 14 16 4 9 1 9 13 2
18 11 1 9 13 9 0 9 2 1 15 9 15 7 13 13 0 9 2
12 15 4 15 13 2 16 4 1 11 9 13 2
7 9 10 9 13 0 9 2
12 3 13 2 15 15 13 1 9 9 1 9 2
23 9 13 2 16 9 0 9 4 15 13 2 14 4 13 0 13 0 0 9 2 0 9 2
9 3 7 2 16 15 7 15 13 2
25 3 13 0 2 16 16 4 3 9 9 9 13 2 13 4 15 9 0 11 9 14 0 9 9 2
29 7 3 3 2 1 9 4 15 13 13 10 9 2 16 3 1 9 4 11 13 1 0 9 2 0 9 7 9 2
27 9 2 16 9 1 11 13 0 9 2 4 0 9 13 1 15 2 16 4 13 3 13 7 13 0 9 2
16 15 4 7 13 9 0 9 9 2 0 9 9 7 9 9 2
27 13 4 15 3 3 3 2 16 4 15 15 1 0 9 13 2 7 3 2 16 4 1 15 13 9 9 2
11 9 13 0 7 13 15 1 9 1 11 2
22 16 9 0 9 13 3 9 0 9 2 1 10 9 15 9 13 9 1 9 0 11 2
10 9 3 0 9 13 4 11 3 13 2
26 16 0 9 13 2 16 1 0 0 9 13 13 2 13 15 15 2 1 9 1 11 2 13 1 9 2
21 3 15 7 13 2 16 10 9 13 3 0 2 7 3 15 4 1 9 13 15 2
7 7 11 1 9 3 13 2
16 7 16 4 9 1 9 13 1 0 9 2 9 4 13 0 2
14 3 4 11 13 3 3 0 2 13 4 15 3 0 2
12 16 0 4 9 0 9 13 13 11 7 11 2
28 12 9 13 3 3 0 2 16 4 15 13 13 13 1 0 9 2 13 7 10 9 2 16 4 13 0 9 2
11 3 7 13 7 9 13 15 1 0 9 2
32 11 2 0 0 9 0 9 7 0 9 0 9 2 4 15 13 1 9 7 13 4 15 1 0 9 0 9 9 1 15 9 2
9 11 4 15 13 3 1 0 11 2
19 7 11 2 3 15 0 13 0 9 2 4 3 13 2 16 13 0 9 2
41 9 4 13 9 0 9 1 0 9 1 9 2 1 15 7 4 13 0 13 2 4 13 9 9 2 9 9 7 9 11 1 9 2 15 4 0 9 13 1 9 2
22 9 13 2 16 4 3 11 13 1 0 15 11 13 7 13 15 0 9 3 1 15 2
17 0 9 4 13 11 13 0 9 2 16 4 15 13 3 1 11 2
17 16 4 15 11 13 1 10 0 9 13 2 15 7 3 1 11 2
4 11 2 11 2
16 9 9 11 11 11 13 1 9 1 11 2 3 13 9 11 2
13 3 2 13 1 12 2 0 9 11 1 0 11 2
5 1 9 9 9 2
21 9 1 0 9 11 11 11 4 13 13 1 9 0 9 9 0 9 12 2 9 2
9 13 15 1 0 9 9 0 9 2
3 0 9 2
25 9 0 15 13 1 9 1 11 7 11 1 0 9 9 1 0 2 0 9 0 11 1 0 11 2
4 1 11 13 9
4 9 0 0 9
2 11 2
22 9 0 9 0 9 9 9 1 11 13 9 11 7 11 2 16 4 13 0 0 9 2
25 1 3 0 9 13 2 16 1 0 9 1 11 13 9 2 13 9 2 13 9 7 13 15 9 2
19 0 2 0 9 2 0 9 11 3 13 9 0 9 0 0 11 11 11 2
32 13 1 15 2 16 0 9 1 0 0 9 1 11 13 0 9 9 0 9 11 2 15 2 13 1 9 9 7 9 0 2 2
12 1 0 9 0 1 12 2 9 13 9 11 2
10 13 15 3 9 0 0 9 11 11 2
20 1 9 2 16 15 9 13 2 2 13 1 9 9 7 4 13 0 9 2 2
12 11 13 2 16 1 10 9 13 1 10 9 2
8 1 11 13 7 9 2 7 0
6 13 15 3 9 10 9
8 11 2 1 10 0 9 2 2
38 11 2 16 10 9 0 11 2 13 1 0 9 10 9 1 0 9 2 12 9 1 9 0 9 0 0 9 2 9 2 0 3 0 9 9 2 1 2
26 3 3 13 15 2 15 9 11 13 1 10 9 2 16 1 10 9 13 2 7 9 2 7 0 2 2
24 3 2 13 15 3 7 15 1 9 2 14 2 15 13 13 3 0 9 7 13 15 1 9 2
18 15 0 2 14 2 2 0 1 9 2 13 3 15 2 15 11 13 2
23 0 9 2 3 16 12 9 2 13 9 10 9 7 15 2 16 13 9 11 1 0 9 2
34 15 2 16 9 2 13 2 2 11 13 9 7 3 13 3 10 0 9 2 16 9 2 15 15 13 1 9 0 9 2 13 3 0 2
30 1 9 13 3 0 9 2 7 15 0 2 1 15 2 15 4 13 13 1 9 9 1 0 0 9 1 9 0 9 2
55 1 15 9 2 16 13 1 9 9 2 0 9 7 9 9 11 2 11 3 13 10 0 9 2 9 9 7 0 9 1 15 13 9 9 10 7 15 9 2 7 9 2 1 15 15 0 13 2 16 13 3 1 0 9 2
25 13 2 14 11 16 9 10 0 9 2 11 2 15 15 15 13 2 15 3 13 2 3 13 0 2
13 11 0 1 9 7 9 1 9 9 3 3 13 2
20 7 1 15 3 15 13 0 9 2 1 0 9 7 0 2 1 15 0 9 2
28 1 0 7 0 11 2 15 13 2 14 2 2 1 11 1 12 5 2 2 7 0 9 2 3 9 0 9 2
37 9 13 14 9 2 7 3 9 2 9 13 2 16 9 1 9 2 15 15 13 11 2 13 0 1 0 0 9 2 3 0 15 13 1 0 9 2
33 11 15 3 3 13 1 9 2 1 9 2 15 15 0 9 13 2 7 0 9 2 15 4 2 3 15 13 2 3 13 1 0 2
7 10 15 13 3 0 9 2
17 9 9 2 7 14 3 0 2 13 7 2 16 15 13 15 13 2
23 3 13 9 1 0 9 2 3 3 3 13 4 13 9 1 15 2 15 15 1 9 13 2
8 11 3 1 15 7 1 15 2
23 15 2 15 15 3 13 2 2 1 9 2 2 13 3 13 13 9 1 9 10 0 9 2
27 7 9 11 2 3 0 7 0 2 2 15 1 15 13 1 9 1 0 9 2 15 1 10 9 3 13 2
6 9 7 9 1 0 9
10 0 2 14 2 2 0 9 13 13 3
2 11 2
16 1 9 13 0 9 0 9 0 9 1 0 9 1 0 9 2
14 3 13 7 1 10 9 13 9 1 0 9 0 9 2
20 9 11 11 13 1 0 2 16 14 0 9 11 2 0 9 2 0 0 9 2
16 11 3 13 1 15 2 16 4 0 9 13 1 9 1 9 2
19 9 9 11 11 13 1 2 9 2 2 15 4 13 1 0 9 1 11 2
16 9 13 2 16 2 0 9 13 3 2 2 13 9 0 9 2
16 1 2 10 9 1 9 2 13 0 9 11 9 9 11 11 2
21 9 1 0 0 9 1 0 9 1 15 13 9 9 9 2 3 16 7 1 11 2
36 0 9 11 11 3 13 9 0 9 1 0 9 1 0 9 7 13 2 16 10 9 11 13 2 9 9 1 9 2 15 4 3 3 13 2 2
18 1 9 9 11 13 3 9 9 11 11 11 9 0 9 1 0 9 2
26 9 9 0 9 2 11 2 11 11 1 9 1 9 0 0 9 1 0 9 3 13 0 9 10 9 2
20 0 9 0 9 13 3 1 11 9 2 1 15 13 9 0 9 1 0 9 2
39 0 9 11 2 15 3 13 1 9 0 9 0 9 2 13 9 9 1 0 11 1 0 9 3 1 9 1 15 2 16 1 9 0 9 13 3 0 13 2
22 0 9 9 11 11 13 3 2 16 9 0 9 4 13 4 1 0 7 0 9 13 2
11 1 10 9 15 7 13 0 9 9 9 2
13 0 0 9 13 0 9 0 9 1 9 1 0 2
23 10 9 4 3 13 13 3 16 3 2 16 11 13 10 9 1 9 2 13 9 11 11 2
17 0 9 13 13 1 9 2 16 15 15 12 0 9 0 9 13 2
22 13 7 13 1 9 1 12 2 9 2 3 3 2 16 4 9 11 13 2 13 11 2
4 11 3 1 11
2 11 2
14 1 0 9 1 0 9 13 1 0 9 12 9 9 2
7 13 15 3 0 9 9 2
10 9 13 3 12 9 2 1 13 12 2
6 0 9 13 12 9 2
23 0 9 4 13 1 9 9 1 0 9 7 9 11 2 3 15 0 9 13 1 12 9 2
50 1 9 1 0 9 9 9 1 9 9 11 11 1 0 0 9 13 2 16 11 15 12 2 9 14 13 9 2 13 9 7 13 9 1 3 0 9 9 2 7 3 13 2 16 13 3 0 13 11 2
31 13 2 16 9 9 13 0 11 2 7 2 3 13 2 1 9 13 10 11 7 16 9 2 7 16 0 2 16 13 3 2
55 9 0 0 9 13 10 9 1 0 9 2 9 9 2 16 3 1 0 7 0 9 2 15 1 9 13 1 9 2 16 11 1 9 13 1 9 0 9 2 9 13 0 9 7 1 10 9 13 9 9 9 2 14 2 2
28 9 9 0 9 11 1 0 9 1 0 9 1 0 9 4 1 0 9 11 13 1 0 9 2 3 7 9 2
10 0 9 13 2 16 0 9 13 13 2
25 0 9 11 11 2 15 1 0 9 13 0 9 2 1 9 13 1 9 9 9 0 9 0 9 2
13 0 9 11 15 4 13 3 12 2 9 1 11 2
16 13 15 3 1 0 11 9 0 9 1 9 9 9 9 11 2
43 9 9 0 9 7 9 0 9 13 1 9 1 9 1 11 9 0 9 1 0 9 7 13 9 0 0 9 2 9 2 2 15 4 13 1 9 0 0 9 2 11 2 2
4 0 9 1 11
4 0 9 1 9
2 9 2
40 0 0 9 2 0 9 11 11 2 3 1 9 0 11 13 2 16 1 9 9 12 2 12 9 1 9 0 0 9 2 13 1 9 11 9 1 9 0 9 2
23 13 2 16 1 9 1 0 0 9 13 1 12 0 9 1 9 11 11 9 0 0 9 2
21 2 13 4 1 9 0 0 9 2 0 9 7 0 0 9 2 2 13 9 11 2
17 9 10 9 13 0 9 2 16 4 13 11 1 9 1 0 9 2
17 0 9 15 1 11 13 1 9 12 2 3 3 2 16 11 13 2
13 10 9 15 7 13 13 7 13 9 1 0 9 2
13 0 0 2 9 2 15 13 1 9 12 2 9 2
6 9 11 1 0 9 11
6 9 9 0 9 0 9
3 0 11 2
28 0 9 13 1 0 9 9 9 11 2 15 4 15 13 9 9 9 0 9 13 0 9 2 13 15 7 13 2
23 13 15 3 1 0 11 0 9 11 11 1 9 9 0 9 1 12 2 9 0 9 11 2
21 9 11 1 15 13 9 2 16 4 13 0 9 15 0 9 2 15 13 0 9 2
34 11 11 13 9 0 9 11 11 11 2 11 2 16 4 0 9 13 0 2 3 0 9 0 3 3 13 1 9 9 9 3 1 9 2
25 1 10 9 13 0 9 9 11 1 9 9 11 7 13 0 9 2 16 4 15 1 10 9 13 2
43 1 11 2 11 13 0 9 7 11 3 1 12 0 9 2 13 0 9 7 13 0 9 2 13 9 9 0 9 7 13 9 1 15 1 9 9 0 9 7 9 0 9 2
4 1 9 15 13
2 11 2
4 1 9 15 13
2 11 2
21 1 9 9 7 9 1 12 9 13 0 9 1 11 9 9 7 0 9 11 11 2
10 11 13 9 0 9 1 2 0 9 2
16 1 0 9 0 9 13 0 0 9 12 9 2 11 7 11 2
27 9 11 11 1 15 2 16 0 9 13 0 9 2 13 13 1 0 12 2 12 2 15 13 2 16 3 2
16 16 9 4 9 13 2 13 0 2 16 9 1 10 9 13 2
14 11 11 7 11 11 15 13 7 7 4 13 13 9 2
18 3 16 3 15 13 13 2 16 4 4 11 13 16 0 9 0 9 2
23 4 3 13 1 10 9 2 16 0 9 13 3 1 9 0 9 7 3 3 0 9 13 2
21 16 13 9 1 9 10 9 2 13 13 2 16 9 13 1 0 9 1 0 9 2
32 11 13 9 0 9 1 2 0 9 2 7 1 15 2 16 9 1 11 13 1 15 2 16 4 11 13 0 9 10 0 9 2
17 1 0 9 13 0 9 2 16 0 9 13 1 0 2 14 2 2
17 9 1 9 0 9 1 0 11 13 3 0 2 16 0 9 13 2
5 11 13 12 9 2
23 13 13 1 9 9 0 2 16 11 15 13 13 1 9 1 0 0 9 7 1 0 9 2
9 15 7 1 11 3 13 0 9 2
29 0 9 0 9 2 15 13 0 9 2 13 0 1 0 0 9 11 2 7 4 13 3 9 9 1 9 0 9 2
25 3 13 9 2 16 0 9 4 13 0 9 15 2 1 15 0 9 13 2 12 0 9 9 11 2
14 0 2 14 2 9 13 9 2 7 9 13 3 3 13
4 13 0 0 9
3 11 11 2
4 13 0 0 9
2 11 2
28 9 0 9 0 9 1 9 13 0 0 9 11 11 1 9 2 15 13 10 9 2 0 0 9 9 11 11 2
22 11 13 10 9 2 16 2 9 0 9 1 10 9 13 4 3 13 0 9 9 2 2
23 10 0 9 7 9 13 1 12 1 0 9 10 9 7 9 0 9 9 13 0 9 9 2
20 11 11 3 13 2 16 11 13 1 10 9 1 9 9 7 9 3 3 15 2
24 3 15 11 2 11 13 1 11 2 11 7 11 16 1 10 9 1 9 1 9 9 1 9 2
5 9 11 1 0 9
5 9 1 9 9 11
2 11 2
43 2 9 0 9 13 0 2 0 9 2 7 9 0 9 7 9 13 9 1 9 2 2 13 1 9 2 9 9 2 2 15 1 10 9 13 1 11 2 0 9 11 11 2
37 0 9 13 1 9 7 10 9 2 10 9 4 13 10 9 1 9 9 1 11 12 2 9 12 7 12 13 1 0 9 2 3 13 0 12 9 2
13 1 9 0 7 0 9 13 13 13 1 0 9 2
19 10 0 0 9 2 15 13 0 9 2 4 13 1 9 9 9 11 11 2
3 11 13 9
2 11 2
3 11 13 9
2 11 2
18 1 0 0 9 1 11 13 7 12 1 12 9 3 16 12 9 9 2
30 1 0 0 9 13 3 9 1 12 0 2 0 9 9 11 11 2 12 9 0 9 2 7 11 11 2 12 9 2 2
14 9 15 13 3 12 9 2 15 13 12 9 0 9 2
2 9 9
6 11 11 2 11 2 2
26 0 9 1 11 13 3 1 9 12 9 0 1 9 0 9 2 1 15 13 1 9 1 11 2 11 2
18 10 9 13 9 3 2 16 9 11 11 2 13 2 16 15 9 13 2
18 9 13 0 1 9 2 1 0 9 13 0 2 16 13 1 0 9 2
6 9 9 13 3 0 2
13 3 4 1 0 11 7 1 11 13 3 12 9 2
3 13 1 11
5 11 2 11 2 2
16 9 3 13 0 1 9 0 9 0 1 9 9 1 0 11 2
9 13 1 15 1 9 12 2 9 2
23 0 9 16 9 13 12 0 9 1 11 7 12 1 11 2 15 15 1 10 0 9 13 2
13 12 4 1 0 9 13 1 9 9 3 1 9 2
13 1 15 4 13 9 7 0 9 4 13 1 11 2
3 1 9 9
23 1 10 9 13 7 1 9 2 1 15 13 9 9 2 7 1 15 2 15 13 0 9 2
4 4 9 13 2
20 1 9 9 13 2 15 10 9 2 2 11 3 12 2 12 2 2 13 13 2
5 3 13 13 15 2
3 15 3 2
16 9 13 2 15 15 13 7 15 15 1 15 4 13 0 9 2
11 13 9 2 16 9 9 13 11 7 11 2
25 9 7 13 2 16 15 9 11 13 2 7 15 13 9 0 11 1 9 0 9 2 9 7 9 2
16 3 13 13 9 11 1 9 9 9 9 1 12 9 7 9 2
12 15 15 13 1 9 2 13 15 3 3 13 2
9 15 0 15 13 9 1 9 11 2
11 13 2 16 13 0 0 9 13 1 9 2
39 13 7 2 16 1 9 11 4 13 0 9 2 1 11 15 3 13 13 0 9 1 0 9 7 0 9 7 0 9 2 16 4 11 13 13 1 9 11 2
7 13 0 13 3 7 13 2
17 7 15 2 13 15 2 11 7 9 11 13 16 0 9 2 2 2
15 3 15 13 2 16 15 13 13 9 7 9 1 0 9 2
11 3 9 2 11 2 9 2 9 2 2 2
14 7 13 9 7 9 1 0 9 15 13 1 9 9 2
14 13 0 2 16 4 13 2 16 15 1 15 13 9 2
54 3 7 9 7 9 13 13 1 9 2 16 1 0 9 2 9 0 9 9 1 15 7 1 0 9 2 1 0 3 0 2 7 3 0 9 9 7 9 13 1 0 9 9 9 1 9 1 12 0 9 10 0 9 2
23 11 2 11 2 13 15 2 16 4 10 9 13 13 2 16 4 3 13 10 0 0 9 2
31 0 9 1 9 11 11 2 11 3 12 2 12 2 2 4 13 9 1 3 0 0 9 11 2 11 7 11 16 0 9 2
11 0 4 13 1 0 9 1 9 0 9 2
18 1 9 11 4 13 1 9 0 9 0 9 7 9 11 13 3 0 2
5 11 11 2 11 12
3 9 1 9
5 11 2 11 2 2
24 9 0 9 12 9 0 9 13 13 2 16 4 9 9 13 9 0 9 9 1 9 7 9 2
11 13 15 1 9 0 2 0 0 9 9 2
18 9 11 4 3 13 2 16 4 4 13 1 9 9 0 9 1 9 2
35 15 4 13 13 0 9 3 2 16 9 1 9 9 9 1 9 7 9 2 3 13 13 1 0 9 2 12 2 9 2 2 13 3 0 2
22 9 13 9 2 16 4 15 13 9 0 9 0 9 9 7 3 3 9 10 0 9 2
5 11 13 9 1 9
16 0 9 3 13 9 1 0 9 0 9 1 9 2 11 2 2
24 9 4 13 9 9 1 10 0 7 0 9 0 9 1 0 7 0 9 7 0 9 7 9 2
13 3 2 16 9 13 12 0 9 2 13 9 3 2
19 9 0 9 4 1 0 9 13 1 0 11 0 9 0 9 2 11 2 2
30 0 0 9 1 9 13 10 9 1 9 7 1 1 15 2 16 1 9 4 13 9 11 2 13 0 13 3 0 9 2
46 11 4 13 9 2 15 13 9 0 1 9 9 2 3 9 0 7 0 9 2 15 13 0 13 2 7 13 15 9 2 3 4 13 4 13 9 1 9 9 2 9 2 9 7 9 2
17 0 9 9 13 3 9 1 0 9 11 7 9 1 0 9 9 2
5 3 10 9 1 11
8 4 13 9 1 9 12 9 9
20 11 13 9 13 15 1 0 0 9 0 12 9 9 2 14 12 9 9 2 2
31 10 1 9 0 9 0 9 0 13 0 9 0 9 2 1 0 9 12 13 0 9 9 12 9 9 2 7 9 0 9 2
22 11 13 3 1 9 11 13 1 9 0 9 12 9 9 2 3 7 13 3 12 9 2
18 10 0 9 1 11 3 13 12 9 9 2 3 12 9 2 9 2 2
49 1 11 11 1 0 9 9 4 9 13 1 11 7 11 1 9 1 9 10 0 9 1 11 2 7 14 1 9 2 16 15 12 0 9 1 11 13 1 0 9 1 9 2 15 15 3 13 0 2
27 16 4 1 0 9 13 2 13 4 12 9 3 1 9 13 2 7 1 9 9 9 11 3 13 15 9 2
36 9 9 10 0 9 2 7 3 7 9 2 15 4 13 9 9 2 7 0 9 12 9 2 0 0 9 2 0 9 2 0 9 3 2 2 2
12 1 9 9 9 1 15 9 9 13 9 11 2
19 0 9 4 13 13 0 1 9 9 2 16 1 10 9 13 0 9 9 2
5 9 9 13 1 9
12 1 11 11 3 13 3 0 2 15 13 1 9
57 16 15 1 9 1 0 9 15 13 1 9 2 16 1 9 0 9 9 13 1 0 9 3 12 9 7 0 3 12 4 13 1 0 9 13 0 9 2 3 3 13 1 15 9 0 2 15 3 7 1 10 9 15 0 9 13 2
12 2 1 0 9 15 1 9 1 9 3 13 2
34 3 13 2 16 9 13 1 12 2 9 7 12 2 9 2 7 3 13 12 9 2 16 4 9 1 9 13 13 12 7 12 9 9 2
36 9 2 15 13 9 1 0 9 3 3 1 12 2 9 2 13 12 9 2 2 13 15 0 9 0 2 9 2 11 2 9 2 11 11 0 2
26 2 13 2 16 4 9 1 0 0 2 9 2 11 4 13 3 2 16 4 1 15 9 13 0 9 2
32 15 13 2 16 13 2 16 4 3 1 9 13 0 9 7 3 14 12 9 2 2 13 9 0 0 9 9 0 9 11 11 2
17 2 9 9 3 13 9 3 3 13 2 15 15 13 1 9 9 2
4 13 9 9 2
29 16 15 13 13 9 7 1 9 2 14 15 15 13 3 2 14 13 9 13 1 12 9 7 13 15 0 9 2 2
24 1 9 0 9 1 9 9 15 3 13 1 9 2 16 1 0 9 3 13 1 12 0 9 2
16 2 3 9 11 13 9 3 1 12 9 2 2 13 11 0 2
12 2 0 9 15 7 13 13 2 16 9 13 2
9 1 9 13 12 9 0 9 2 2
5 9 9 13 1 9
25 1 9 0 9 1 9 15 9 9 0 11 13 1 12 1 12 7 0 9 9 15 1 9 13 2
18 3 7 1 9 9 1 11 13 1 0 9 1 0 9 9 0 9 2
38 0 9 9 2 15 13 9 2 1 12 3 0 13 15 3 12 9 9 7 9 2 1 10 9 15 13 3 1 9 9 2 3 13 9 1 0 9 2
21 2 1 11 13 1 10 9 1 12 9 0 9 7 3 0 13 3 9 1 9 2
6 9 1 9 7 13 2
25 3 4 3 0 9 3 1 0 9 13 0 9 13 2 2 13 9 9 9 9 1 11 11 11 2
12 2 3 1 9 9 13 1 9 9 10 9 2
15 4 13 2 16 4 15 9 1 9 13 3 3 13 2 2
2 11 11
45 2 15 10 9 2 15 13 13 13 7 3 13 9 2 13 3 1 12 0 9 2 9 7 9 1 9 7 9 2 2 13 3 1 11 0 9 7 9 9 9 11 11 11 0 2
26 1 9 3 13 1 0 12 9 2 9 11 7 13 2 16 1 9 9 4 13 13 9 1 9 0 2
13 11 11 13 9 0 9 9 3 1 9 1 9 2
46 16 4 13 3 0 9 2 13 1 10 9 1 9 0 9 0 9 2 2 13 7 1 10 0 9 2 16 0 9 13 3 13 7 13 4 4 13 1 12 2 9 2 2 13 11 11
4 2 2 11 2
14 9 9 1 9 9 9 7 9 9 0 9 13 0 2
9 13 15 3 0 9 9 11 11 2
24 1 9 0 9 9 9 9 2 15 13 13 1 11 2 13 2 16 9 10 9 13 15 13 2
21 9 11 13 9 9 2 7 16 13 1 10 9 1 9 2 0 7 0 9 9 2
18 2 7 2 0 9 13 9 2 15 4 13 13 10 9 1 0 9 2
15 0 9 1 9 10 9 7 3 13 2 2 13 11 11 2
3 11 13 9
39 3 1 12 9 2 10 9 15 3 13 1 0 7 0 9 0 9 2 13 0 2 16 4 9 0 0 9 13 1 9 0 9 9 1 9 1 0 9 2
10 13 15 1 0 9 9 11 7 11 2
21 13 1 10 0 2 9 2 2 1 15 9 13 1 12 12 9 2 12 9 2 2
27 7 10 9 13 13 1 0 11 2 15 4 13 12 2 9 9 13 9 2 15 1 15 9 1 9 13 2
35 3 4 9 13 10 9 13 9 9 7 10 0 9 3 1 15 2 16 15 9 0 2 9 2 13 3 2 3 1 9 0 9 0 9 2
39 1 0 9 11 13 9 2 16 0 9 4 13 13 7 1 9 2 3 13 1 0 7 0 9 14 0 9 7 11 3 3 13 12 9 0 9 1 9 2
13 11 7 1 0 9 13 0 9 1 9 10 9 2
29 9 9 13 7 9 13 9 1 0 9 10 11 3 1 0 9 2 3 0 12 12 9 13 3 9 9 7 11 2
2 1 9
3 9 3 13
35 1 0 0 9 1 11 2 11 2 13 1 0 0 9 0 9 2 15 4 3 13 1 9 12 9 1 0 9 1 12 9 1 0 9 2
26 1 9 11 11 11 15 0 9 9 9 13 3 7 3 13 2 16 1 11 13 0 9 1 9 9 2
9 9 0 9 1 11 13 3 0 2
18 3 4 13 12 9 9 2 16 0 9 1 0 9 13 12 9 9 2
4 9 2 11 3
5 9 2 0 0 9
19 9 0 9 1 0 9 3 13 2 15 9 13 1 0 9 9 9 3 2
18 0 13 10 9 1 11 2 3 15 13 3 13 3 3 1 9 9 2
3 11 1 11
17 12 1 0 0 9 9 2 9 11 2 13 1 11 9 10 9 2
27 13 1 0 0 0 9 2 15 1 11 2 3 13 0 9 3 1 9 0 0 9 2 4 13 10 9 2
28 9 4 1 10 0 9 13 13 12 2 1 11 3 9 13 12 9 2 7 13 15 1 15 4 7 0 9 2
21 11 4 1 11 13 9 0 9 2 1 15 13 0 9 0 11 7 0 9 11 2
12 9 11 3 1 11 13 12 9 7 12 9 2
19 1 9 9 11 11 7 4 13 1 9 7 1 0 9 7 1 9 9 2
8 0 9 1 9 4 13 1 0
36 0 0 0 9 0 9 1 9 9 9 1 11 13 1 9 12 11 11 2 0 2 9 2 2 1 9 2 15 13 1 9 1 0 9 11 2
7 9 13 9 12 9 9 2
20 16 9 9 1 9 9 1 0 9 13 11 3 0 9 1 11 1 15 9 2
5 11 2 0 0 9
5 2 9 2 12 2
2 9 3
7 11 11 2 9 9 12 2
15 16 1 0 9 13 11 12 9 2 0 13 1 0 9 2
23 1 9 11 2 15 13 3 0 9 1 0 9 2 13 0 9 0 9 1 9 11 9 2
5 0 9 9 11 2
27 9 11 2 11 7 11 11 15 13 0 9 2 9 1 9 2 9 3 3 0 2 1 9 10 0 9 2
18 1 0 9 11 11 15 13 3 7 3 1 12 9 1 9 1 0 2
6 0 9 2 9 9 2
8 0 9 0 0 9 13 11 2
21 9 15 13 1 0 11 2 4 13 1 0 9 9 2 16 9 4 13 11 11 2
1 9
31 9 11 2 11 7 11 2 11 13 3 1 9 9 11 2 11 2 9 1 9 9 2 11 7 0 2 11 0 1 11 2
13 11 11 11 13 1 9 3 1 0 9 11 11 2
18 11 11 2 9 2 11 1 0 11 3 13 1 12 9 1 9 9 2
13 0 9 11 7 11 11 13 3 1 0 9 9 2
2 0 9
14 3 13 1 0 9 2 13 15 12 1 10 0 9 2
38 3 0 0 9 1 0 2 0 2 9 2 0 9 11 1 0 9 9 0 2 1 9 0 0 9 11 1 11 2 1 9 7 1 0 9 0 9 2
12 11 11 13 7 3 2 3 15 13 0 9 2
16 1 0 9 15 13 1 0 9 9 11 2 15 15 3 13 2
16 9 9 9 9 11 11 13 10 9 1 0 9 9 1 9 2
40 9 11 11 13 3 0 0 2 9 2 2 11 11 2 11 2 3 3 2 0 1 0 9 7 9 7 11 11 2 11 2 16 0 9 2 15 13 1 9 2
35 1 9 0 9 15 3 13 11 9 2 7 7 10 11 2 15 1 10 9 13 1 0 9 2 13 10 0 9 1 9 0 2 9 2 2
4 9 2 11 2
2 11 11
2 9 13
5 11 11 2 9 2
42 3 4 15 13 1 12 2 0 9 0 9 1 11 1 11 2 3 4 13 1 10 9 9 1 9 12 9 2 0 9 7 9 11 2 15 13 0 9 1 0 9 2
33 1 15 15 9 13 1 0 9 2 11 2 11 2 11 2 13 15 3 3 2 16 13 1 9 2 16 4 15 13 1 12 9 2
26 3 10 0 9 1 9 13 2 7 3 1 15 1 11 3 1 9 13 16 1 2 9 0 9 2 2
11 3 15 13 2 16 9 0 9 13 9 2
16 16 4 13 13 2 16 15 1 0 0 9 13 0 0 9 2
3 9 1 11
30 1 0 9 10 9 13 9 12 1 9 1 0 0 9 1 11 2 3 3 13 3 16 9 11 2 0 9 0 9 2
16 0 9 4 13 0 9 9 0 11 2 11 7 11 1 0 2
2 11 2
16 3 13 0 0 9 2 0 2 0 2 0 2 7 0 11 2
24 1 9 15 13 9 13 1 11 2 11 7 12 9 2 0 9 3 4 13 11 7 0 9 2
11 9 0 9 12 9 9 12 9 1 9 9
22 10 9 1 0 9 0 9 15 13 9 12 0 9 7 0 9 1 0 7 0 9 2
7 11 9 2 9 0 9 2
12 1 0 9 1 9 11 15 13 13 0 9 2
27 16 11 13 10 9 14 1 9 0 9 2 13 3 9 11 9 1 10 9 7 9 9 0 9 1 9 2
18 1 9 4 13 1 9 11 2 11 7 9 11 1 0 7 0 9 2
11 1 11 15 13 0 9 0 2 0 9 2
33 0 9 2 0 9 2 13 13 12 0 9 7 1 9 9 12 2 0 1 9 3 3 2 13 4 1 9 13 7 0 0 9 2
24 13 7 1 9 0 9 1 9 0 7 0 9 2 15 15 4 1 9 1 10 0 9 13 2
29 1 10 9 15 13 13 7 11 3 0 9 7 0 0 0 9 2 3 9 2 15 4 9 1 9 0 9 13 2
18 0 9 4 13 14 0 9 2 0 4 13 2 3 2 7 1 11 2
16 7 3 0 9 2 9 0 9 4 15 13 13 1 10 9 2
23 15 13 9 14 1 9 9 11 7 10 9 2 1 9 9 15 13 1 0 9 0 9 2
7 11 11 2 9 0 9 2
24 13 15 2 16 4 1 11 13 4 13 0 9 0 9 3 2 3 15 13 1 0 9 11 2
50 15 13 2 16 4 1 12 9 13 0 9 16 0 9 1 9 2 1 9 0 7 9 0 9 2 2 0 2 3 0 9 2 7 1 9 0 3 9 0 2 0 2 15 4 13 1 9 0 9 2
55 13 15 2 16 1 11 4 13 4 13 12 0 9 2 0 11 7 0 9 9 12 2 2 16 4 13 1 9 13 9 2 0 2 0 2 0 2 0 9 7 12 0 9 1 9 9 13 3 2 16 4 15 3 13 2
21 0 2 0 9 12 2 7 0 9 2 3 0 9 4 4 13 1 0 0 9 2
39 1 0 9 11 7 11 4 15 0 13 2 16 12 13 0 0 9 1 9 9 2 1 9 11 2 2 15 13 9 0 7 0 9 7 3 13 9 9 2
25 1 15 3 3 13 1 9 12 2 3 13 3 0 9 9 2 7 1 15 0 9 0 9 13 2
12 11 11 2 9 0 9 1 0 7 0 9 2
15 9 13 9 11 7 0 2 9 1 9 9 9 1 0 2
24 1 9 0 9 9 9 15 13 1 9 0 9 2 7 15 7 0 9 9 9 0 0 9 2
50 13 3 2 16 4 0 0 9 13 9 1 0 9 3 1 9 9 9 0 9 2 15 13 9 2 7 16 4 15 9 1 9 9 7 9 13 3 2 16 4 4 3 0 9 13 9 7 9 9 2
13 15 15 13 0 9 2 0 9 7 3 15 13 2
27 1 2 0 2 9 15 13 2 16 0 9 3 13 2 3 0 9 9 13 2 7 1 9 9 3 13 2
33 1 9 11 11 11 7 9 0 0 9 13 15 3 2 9 13 3 1 12 2 9 13 0 9 2 3 13 0 13 0 0 9 2
59 7 16 9 0 9 4 13 2 2 0 2 13 15 2 16 1 0 9 0 11 4 13 4 13 9 3 1 0 9 7 16 3 13 13 1 9 2 13 2 14 2 4 2 14 13 13 2 3 13 2 0 9 12 7 14 0 9 12 2
9 7 9 0 9 13 7 3 13 2
21 13 15 3 3 2 16 9 11 0 1 0 0 9 9 10 2 9 2 3 13 2
20 13 1 0 9 2 1 9 9 2 7 1 3 0 9 2 15 13 0 9 2
32 9 7 13 3 0 2 9 3 11 2 13 1 9 12 0 9 0 11 0 11 11 2 2 9 15 13 11 2 0 2 9 2
8 0 9 7 13 1 9 0 2
23 13 3 0 9 9 2 15 3 13 0 2 9 2 7 2 9 2 1 9 7 9 9 2
19 1 9 2 3 13 0 9 0 2 13 3 9 9 13 0 9 2 2 2
13 7 3 15 3 9 1 0 9 13 1 0 9 2
61 7 7 16 4 2 1 9 9 2 11 11 3 13 9 12 2 0 0 9 2 2 7 16 4 11 11 16 9 9 13 3 9 3 13 2 13 4 15 13 9 2 7 1 0 9 3 0 9 4 13 0 0 9 2 15 4 15 11 3 13 2
39 1 10 0 9 1 0 9 13 3 0 0 9 2 16 3 3 2 1 9 0 9 3 13 0 9 7 9 9 2 1 15 15 3 9 9 13 2 2 2
51 13 15 2 1 0 9 0 0 9 2 7 3 13 0 0 9 2 0 9 0 9 1 9 9 2 0 9 1 9 11 2 2 3 13 0 9 9 2 13 0 9 2 2 1 9 2 3 1 9 12 2
4 2 3 11 2
17 14 3 2 16 15 15 13 2 14 2 2 13 11 3 0 9 2
21 6 2 9 0 2 0 2 0 0 0 9 3 3 16 11 9 1 9 1 9 2
2 0 9
25 0 0 9 11 11 4 3 1 11 13 11 11 1 9 9 9 7 11 11 1 9 0 9 9 2
33 9 11 2 11 2 0 3 1 9 0 9 2 13 9 9 12 1 11 1 9 12 1 9 9 0 0 2 9 0 9 1 9 2
21 13 1 15 13 4 0 7 0 0 9 0 1 0 12 9 1 11 7 1 9 2
4 11 16 9 2
9 11 11 13 1 11 1 9 12 2
35 12 9 3 2 1 15 12 2 13 1 0 0 9 9 10 0 9 9 9 2 12 2 15 3 13 1 0 2 9 1 9 0 9 11 2
99 9 9 2 12 13 0 9 11 1 9 9 0 2 9 0 9 9 2 9 0 9 7 0 9 2 9 9 2 0 9 2 0 0 9 3 2 13 11 11 9 0 9 2 1 10 0 9 2 3 1 9 2 15 13 0 9 11 2 0 9 2 15 3 3 13 1 10 0 9 2 3 7 3 3 13 15 0 0 9 10 0 2 9 2 2 0 9 2 9 7 9 2 9 2 0 2 2 2 2
27 13 15 11 0 3 7 3 2 1 10 9 2 14 3 3 2 7 15 3 1 9 9 3 13 9 9 2
18 0 9 13 0 9 2 10 9 13 3 0 7 3 15 13 0 9 2
32 0 9 9 1 9 13 0 9 0 9 2 16 7 0 11 13 9 2 10 9 15 9 13 7 10 9 15 1 0 9 13 2
11 1 9 2 7 1 9 2 15 4 13 2
4 9 2 9 2
2 0 9
6 13 12 9 12 0 9
25 13 0 2 0 2 9 1 11 2 12 9 12 2 0 2 9 2 0 9 1 0 9 9 2 12
7 9 2 2 12 2 12 12
4 9 1 9 2
5 0 9 1 9 11
12 9 1 9 0 9 2 0 9 7 0 9 9
3 9 12 13
5 11 2 11 2 2
17 0 0 7 0 9 9 9 9 2 12 13 3 1 0 9 9 2
34 9 2 15 13 0 9 11 11 7 11 0 1 9 1 0 9 0 11 9 2 9 2 0 2 2 13 3 1 11 0 9 11 11 2
10 9 13 3 0 11 11 12 11 12 2
10 12 9 13 1 10 9 10 9 11 2
18 1 0 9 13 9 0 11 2 0 2 9 1 0 9 0 9 11 2
35 3 3 0 9 9 12 0 9 9 9 2 15 4 13 13 3 16 9 12 9 2 15 1 9 1 9 9 13 2 3 4 13 13 3 2
4 0 9 15 13
10 1 9 9 12 2 9 9 13 10 9
35 1 1 9 1 9 1 11 4 1 9 0 2 9 1 11 11 11 13 0 2 16 4 10 9 1 0 9 11 2 11 1 11 3 13 2
21 2 3 15 13 15 13 2 7 10 9 4 13 13 3 3 2 2 13 11 11 2
30 3 15 3 13 2 0 9 13 1 0 9 13 2 2 13 15 1 0 0 9 3 1 9 2 3 7 1 10 9 2
17 3 15 13 7 1 9 0 9 0 9 1 0 9 3 1 9 2
17 16 4 7 10 9 13 13 3 2 4 13 1 0 9 13 2 2
21 3 9 0 1 9 0 9 12 2 9 13 11 11 1 0 9 3 3 0 9 2
9 9 9 13 1 11 11 3 0 2
19 9 1 15 13 15 9 2 15 15 13 9 1 9 11 2 7 10 9 2
25 2 10 0 9 1 9 12 2 9 2 1 15 13 4 13 3 10 9 9 2 7 0 9 13 2
14 9 3 3 13 7 1 9 1 15 15 15 13 2 2
24 1 9 9 11 11 11 4 1 9 1 0 9 1 0 9 2 11 13 0 7 0 9 2 2
35 2 1 9 9 2 15 4 13 0 9 2 13 4 13 14 9 2 7 9 0 9 2 15 13 13 9 9 2 2 13 3 11 2 11 2
14 9 0 9 13 1 0 2 3 16 0 7 0 9 2
13 2 10 9 15 13 9 2 16 0 9 13 9 2
17 13 15 13 9 1 0 9 1 0 9 2 2 13 1 10 9 2
18 9 0 9 13 1 11 2 11 0 7 13 15 15 3 3 0 9 2
3 9 1 11
5 11 2 11 2 2
30 9 0 0 9 2 10 9 13 9 7 9 0 7 0 0 9 2 4 3 13 1 9 1 11 2 0 9 2 12 2
33 10 9 2 0 9 11 2 0 11 2 11 7 11 0 11 2 15 10 9 13 1 9 0 0 7 0 9 1 9 0 9 11 2
21 9 4 13 1 9 2 16 0 9 4 3 13 4 13 1 9 7 0 0 9 2
29 9 4 1 9 9 9 2 11 11 2 15 13 1 9 0 9 2 13 1 9 9 9 1 11 7 0 0 9 2
11 0 0 9 2 1 9 9 13 13 9 2
13 0 1 9 0 0 9 13 3 0 9 0 9 2
18 1 9 1 0 9 1 0 9 9 13 0 9 1 12 0 9 9 2
17 9 9 15 13 1 11 7 1 9 13 2 16 15 13 13 9 2
12 2 9 2 4 3 13 1 0 9 0 9 2
27 1 0 7 0 13 0 15 0 2 9 2 0 9 9 9 1 9 7 9 0 9 0 2 11 11 11 2
15 2 9 15 13 9 9 13 3 2 3 3 13 9 13 2
24 13 3 9 13 2 16 15 2 15 15 15 13 1 9 2 13 3 0 9 2 7 14 9 2
11 3 4 15 3 13 13 1 9 0 9 2
34 16 4 13 9 7 13 15 1 9 7 9 7 9 7 9 15 13 1 9 7 9 13 2 13 4 15 1 9 2 2 13 11 11 2
19 3 9 0 0 9 11 11 13 2 16 3 15 9 9 13 9 0 9 2
26 2 9 7 10 9 13 13 1 9 12 7 9 12 9 0 9 9 9 11 9 2 12 2 12 9 2
18 9 9 13 0 3 1 9 2 16 13 1 0 9 7 1 0 9 2
13 1 0 9 7 13 13 9 2 2 13 9 11 2
22 9 2 16 9 4 13 3 2 4 1 9 0 9 1 0 9 0 9 9 11 13 2
21 2 1 15 13 0 13 3 3 3 10 0 9 2 1 15 13 1 9 13 9 2
25 1 9 0 9 7 13 0 9 2 16 15 15 13 9 1 9 13 0 9 2 2 13 9 11 2
29 1 0 9 0 9 9 13 2 9 2 9 2 3 3 15 13 0 0 9 2 14 2 0 9 1 9 9 2 2
25 2 13 3 0 13 15 2 15 13 1 0 9 2 9 7 13 15 3 1 9 9 1 0 9 2
9 3 16 13 1 9 0 13 9 2
12 0 3 13 13 2 7 16 14 0 2 9 2
14 7 15 15 2 16 15 13 2 0 0 9 13 2 2
4 9 9 9 13
5 11 2 11 2 2
18 9 9 11 3 1 9 13 13 9 9 11 9 2 11 2 11 2 2
24 1 9 13 12 9 2 3 1 11 2 11 2 11 2 11 2 1 13 12 2 13 15 12 2
21 1 13 7 9 9 11 2 7 15 7 3 2 16 0 7 0 9 13 13 1 2
26 0 9 1 11 12 2 15 13 1 11 9 0 9 1 9 9 9 7 10 9 2 1 15 13 11 2
29 9 9 15 0 9 13 13 3 1 9 2 3 1 9 1 9 9 13 0 9 11 11 1 9 2 9 7 9 2
10 1 0 9 0 9 13 9 1 9 2
9 1 9 15 0 11 11 13 9 2
19 0 9 9 3 13 2 16 11 9 13 4 3 3 1 0 0 9 13 2
28 9 11 9 1 0 0 9 11 3 13 2 16 0 7 0 9 9 9 11 13 2 16 4 4 13 0 9 2
11 1 10 0 0 9 15 4 3 13 9 2
6 1 11 7 11 0 9
7 9 0 9 11 15 3 13
22 0 9 0 11 11 11 11 7 11 11 13 1 9 0 9 0 1 0 9 1 11 2
27 0 0 9 2 0 1 12 0 9 2 13 1 11 12 0 9 2 1 12 9 1 11 13 9 12 9 2
12 1 0 9 13 0 9 9 1 11 12 9 2
24 3 0 9 1 11 13 9 11 2 15 13 1 0 2 0 9 1 11 2 13 15 12 3 2
16 11 2 13 1 11 2 13 12 2 3 13 2 3 2 12 2
21 0 9 1 11 15 13 3 0 9 11 11 2 15 15 13 1 12 1 12 3 2
11 0 1 11 13 9 11 1 9 12 9 2
35 0 9 11 13 3 1 11 12 9 2 1 11 15 13 3 12 2 3 1 9 2 7 1 12 9 4 15 10 9 13 13 14 1 12 2
12 3 14 12 9 1 11 13 1 12 9 3 2
19 12 1 15 13 0 9 11 2 1 11 7 3 13 0 9 1 12 9 2
6 0 2 9 2 9 13
6 9 1 12 2 9 11
13 0 2 9 2 9 13 0 9 1 11 1 0 9
31 0 9 4 13 0 9 2 0 9 11 2 11 1 0 12 9 13 1 0 9 3 12 9 3 0 9 2 1 0 9 2
9 3 11 3 1 0 9 3 13 2
14 7 1 9 13 11 0 7 9 1 12 9 13 0 2
13 0 9 0 13 0 9 11 2 0 9 1 9 2
16 14 12 9 1 9 15 13 1 0 9 0 9 0 11 13 2
23 1 9 0 9 11 2 0 9 2 2 12 9 13 3 0 2 1 0 9 13 9 2 2
16 1 11 13 3 9 9 1 0 11 11 11 2 9 0 9 2
35 9 9 13 10 0 9 2 0 9 7 13 0 2 9 13 0 7 0 9 2 9 11 2 11 2 9 11 7 1 9 7 0 0 9 2
34 13 3 0 9 3 13 2 3 13 1 9 3 1 9 9 11 7 11 1 11 11 2 1 11 3 11 13 2 16 9 13 3 13 2
13 12 9 13 0 9 2 0 9 13 9 0 9 2
34 9 11 11 2 2 13 0 9 2 13 1 9 1 0 9 2 13 9 7 1 9 9 2 1 12 2 9 4 1 9 13 12 2 2
9 11 11 15 3 13 1 9 11 2
25 1 11 13 14 1 9 0 9 11 11 1 0 0 9 2 0 3 13 9 7 1 9 13 11 2
24 7 1 11 3 13 9 1 2 9 2 2 10 0 9 2 13 9 2 13 2 3 13 3 2
26 3 3 2 16 9 1 10 0 2 9 2 2 3 0 9 0 1 0 9 1 11 2 1 11 13 2
10 3 9 9 2 7 0 9 2 2 2
29 9 12 0 9 2 13 13 0 11 2 0 9 2 7 0 11 2 11 3 1 12 2 9 2 12 9 1 9 2
4 0 9 0 9
12 11 13 9 9 2 0 2 9 13 15 13 9
27 1 0 0 9 2 1 10 9 14 12 9 9 2 13 0 2 0 9 13 9 0 9 1 0 9 9 2
13 13 15 1 9 0 9 9 11 11 1 11 3 2
19 0 9 1 9 11 13 0 9 9 2 9 0 9 1 11 7 13 9 2
31 2 9 4 13 0 2 1 9 2 7 13 3 9 0 9 2 12 9 1 9 2 12 9 1 11 2 2 13 9 11 2
24 2 0 0 9 13 1 9 9 1 9 2 3 4 3 1 9 13 2 16 9 15 13 13 2
16 2 13 2 16 15 13 7 0 9 1 0 9 1 9 13 2
15 1 12 0 9 2 16 15 13 2 13 3 9 12 9 2
14 0 13 1 15 2 16 4 15 13 3 15 13 2 2
18 2 15 15 3 13 2 7 13 15 2 16 9 13 3 1 9 9 2
10 2 9 13 1 11 12 0 0 9 2
23 7 3 1 15 13 0 9 2 15 13 0 13 2 16 1 9 9 9 12 9 13 2 2
10 2 3 1 15 13 1 9 12 9 2
26 2 10 9 7 10 9 2 1 15 13 11 9 2 13 1 9 2 7 3 14 13 1 0 9 2 2
12 2 13 15 15 2 16 9 9 15 3 13 2
5 9 13 9 9 2
21 2 15 4 13 0 2 16 4 13 9 3 13 2 7 1 10 9 13 3 13 2
10 3 13 3 1 9 10 9 9 2 2
7 2 13 3 3 2 2 2
16 2 16 4 12 0 9 13 2 13 4 15 9 12 9 2 2
8 2 3 3 9 13 2 2 2
18 2 4 13 1 15 2 10 9 15 3 1 9 7 9 13 13 2 2
11 2 13 1 9 1 11 7 9 3 13 2
15 2 9 4 13 1 11 7 9 2 9 1 15 13 2 2
7 2 15 13 3 0 9 2
9 2 9 15 13 1 12 9 2 2
13 2 13 0 0 9 9 3 3 13 1 9 9 2
12 2 0 9 9 13 12 9 7 13 13 0 2
11 13 4 13 2 1 10 9 9 13 2 2
2 0 9
28 0 9 2 0 12 2 9 0 9 1 12 9 0 0 9 2 15 13 7 1 9 0 11 1 9 1 11 2
21 1 9 15 13 12 2 9 9 11 2 11 2 15 13 0 9 11 1 0 9 2
14 9 13 1 12 2 9 1 11 2 9 1 0 11 2
32 9 15 13 1 9 1 12 1 12 9 2 1 9 11 2 1 9 12 2 11 12 7 1 9 1 12 9 1 9 11 11 2
3 9 13 9
25 9 1 9 2 3 13 9 12 9 0 0 9 2 11 11 7 11 11 2 15 13 9 11 3 2
19 13 1 15 1 0 2 16 14 3 13 13 1 10 9 1 9 0 9 2
14 16 3 1 10 9 15 13 2 13 15 9 2 9 2
8 7 10 9 1 9 3 13 2
11 9 1 9 15 1 0 9 13 9 9 2
18 12 9 3 13 2 16 1 9 0 9 15 13 3 0 9 2 9 2
18 7 16 15 10 9 13 13 1 9 9 2 13 4 10 0 9 13 2
17 9 11 7 11 7 13 2 16 1 0 15 9 1 9 13 15 2
13 13 1 9 2 15 15 13 13 2 15 13 13 2
28 1 9 13 9 2 16 9 13 13 10 9 1 10 9 3 3 3 2 16 4 13 3 2 3 7 1 9 2
3 11 13 14
3 11 13 11
18 9 0 0 9 11 11 13 1 9 11 11 1 11 1 12 9 9 2
8 13 15 3 1 11 9 11 2
16 1 9 0 9 13 11 12 9 9 1 9 7 9 1 9 2
15 1 9 1 11 11 2 9 9 1 11 1 11 7 0 11
22 0 0 0 9 1 15 0 1 9 13 1 9 0 9 7 9 10 9 9 11 11 2
14 13 1 0 9 1 0 9 10 0 9 1 9 9 2
5 2 13 0 9 2
25 3 4 1 9 9 11 11 2 9 1 11 1 11 2 13 3 9 0 11 11 1 0 0 9 2
6 9 7 13 1 9 2
6 13 4 3 0 9 2
17 9 3 13 2 16 10 0 9 13 3 3 0 9 16 0 9 2
19 9 10 0 9 9 4 13 9 2 3 9 1 0 9 3 13 0 9 2
24 14 1 9 2 16 9 10 0 9 1 9 13 2 9 15 1 9 3 13 1 0 9 2 2
3 11 13 9
16 1 9 13 9 11 2 11 12 9 0 9 1 11 1 11 2
38 3 13 9 11 11 2 12 2 11 2 12 2 11 2 2 0 9 13 11 2 11 11 2 2 15 13 3 12 2 1 9 12 2 12 9 1 11 2
9 1 9 3 13 11 2 11 2 2
55 1 9 9 3 13 9 11 2 12 2 11 2 12 2 11 2 2 11 1 11 12 12 5 12 13 1 9 12 2 2 2 12 2 12 9 2 2 11 1 9 12 12 5 12 13 12 2 2 2 12 2 12 9 2 2
3 11 1 11
20 3 13 1 9 1 12 0 9 1 11 2 11 13 11 11 1 9 1 11 2
12 2 9 2 13 13 9 10 9 1 9 9 2
13 3 3 1 0 9 2 3 11 13 1 9 11 2
3 11 13 9
7 11 11 15 13 1 11 2
14 3 15 1 15 13 9 0 9 11 11 7 11 11 2
24 1 9 1 11 11 2 15 1 15 11 13 7 9 1 0 12 9 9 2 13 13 1 11 2
21 3 7 1 15 13 3 7 9 11 13 13 2 11 3 13 9 11 1 0 9 2
3 11 13 14
2 11 13
18 9 0 0 9 11 11 13 1 9 11 11 1 11 1 12 9 9 2
8 13 15 3 1 11 9 11 2
16 1 9 0 9 13 11 12 9 9 1 9 7 9 1 9 2
5 2 13 3 13 2
18 13 3 0 2 16 15 3 13 2 2 13 1 9 1 9 11 11 2
8 9 1 11 13 3 12 9 2
21 11 3 1 11 3 13 12 9 9 2 16 11 13 9 1 9 12 2 12 9 2
3 9 15 13
1 9
16 1 9 11 2 11 2 1 11 13 0 7 9 0 9 11 2
12 13 15 3 13 1 9 9 1 11 1 11 2
24 0 9 9 9 12 1 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2
3 9 15 13
22 9 0 3 9 16 0 9 13 1 0 12 0 9 9 0 11 2 15 13 11 9 2
18 1 9 0 0 9 2 0 0 1 12 2 9 2 11 13 1 9 2
18 9 1 0 9 13 11 10 9 1 0 9 2 3 15 13 9 9 2
24 0 9 0 7 9 1 0 9 15 13 0 9 11 2 13 15 7 14 12 2 12 2 12 2
33 11 3 13 1 12 9 9 2 12 2 12 2 1 9 15 13 0 9 2 3 9 1 0 9 1 9 15 11 13 9 1 9 2
7 13 15 3 3 13 11 2
25 3 11 13 1 0 9 1 10 0 7 0 9 7 0 9 9 11 1 12 0 9 1 0 9 2
4 9 13 9 2
8 9 13 1 9 9 0 11 2
29 0 13 9 2 13 12 9 7 1 12 2 9 2 13 12 2 12 1 0 9 0 2 11 7 9 11 1 0 2
8 0 13 9 2 1 9 2 2
12 1 9 0 12 13 2 7 0 13 9 11 2
21 1 0 9 11 13 11 0 9 2 16 4 3 11 7 11 13 1 12 2 12 2
10 1 9 3 14 9 13 1 0 9 2
17 0 13 3 2 1 9 1 12 9 13 9 7 0 12 9 13 2
19 1 0 9 13 0 9 0 2 10 9 13 13 1 0 9 1 0 9 2
16 0 9 11 3 13 9 9 2 3 7 1 12 9 3 13 2
21 9 13 9 2 13 1 9 2 7 16 0 1 12 2 9 13 1 12 2 12 2
25 1 12 9 3 9 13 9 2 7 1 12 2 9 13 2 16 4 11 9 13 1 12 2 12 2
17 1 0 9 7 9 13 9 2 15 12 9 1 9 13 0 9 2
10 1 0 9 13 9 14 1 0 9 2
18 11 1 9 1 0 9 13 1 9 7 1 12 9 13 9 1 9 2
14 15 15 13 1 9 2 13 9 7 13 0 12 9 2
20 0 12 15 13 0 2 7 0 2 9 2 13 0 11 1 9 7 0 9 2
11 1 0 9 9 1 0 9 15 0 13 2
15 3 1 0 9 13 1 0 9 9 7 0 11 15 13 2
15 1 12 2 9 13 3 1 12 9 1 9 11 7 11 2
18 1 0 9 3 11 11 13 2 7 9 9 3 13 11 1 0 9 2
18 16 11 1 12 9 0 12 13 3 9 2 13 1 0 9 9 3 2
13 13 0 7 0 1 9 2 3 15 3 13 11 2
12 9 16 9 2 1 15 9 13 0 0 9 2
10 0 13 0 9 2 7 13 1 9 2
7 7 9 11 11 13 0 2
19 9 0 12 13 9 9 2 12 1 0 11 7 14 12 1 11 2 11 2
13 12 9 3 13 1 9 7 13 15 13 0 9 2
23 0 0 9 11 7 13 7 0 9 2 0 9 13 11 2 11 7 11 13 1 0 9 2
22 3 3 11 2 11 13 0 9 0 9 2 3 13 9 2 7 9 15 3 13 3 2
16 9 7 3 13 0 9 7 11 12 9 1 12 9 13 9 2
18 11 3 13 15 1 0 2 3 15 13 0 11 2 7 13 14 9 2
28 0 12 13 1 9 0 9 1 9 9 2 12 2 0 2 9 1 9 12 9 2 7 13 15 12 2 12 2
24 1 0 0 0 9 2 12 9 1 9 2 13 11 1 9 9 2 7 9 1 9 13 3 2
11 9 11 11 13 0 9 1 9 11 1 11
2 1 9
16 0 9 1 0 9 1 9 1 9 1 11 13 0 2 9 2
12 11 1 0 9 2 9 2 13 14 1 9 2
19 1 9 1 9 4 13 1 11 9 9 9 11 11 2 11 2 12 2 2
13 1 9 13 9 10 9 7 13 15 10 0 9 2
31 1 11 1 0 2 9 15 13 9 9 0 0 9 11 12 0 9 7 0 9 9 1 9 0 1 12 9 9 11 11 2
21 0 9 11 3 0 1 9 7 9 15 13 1 9 1 9 1 0 9 1 11 2
32 9 11 2 15 16 0 9 1 9 12 13 1 11 1 11 0 0 9 2 13 1 11 9 2 16 15 3 13 13 9 0 2
30 0 9 11 2 15 13 1 12 9 0 9 7 13 12 9 1 9 0 9 2 15 3 13 1 9 9 1 0 11 2
18 11 11 2 0 9 9 9 12 13 2 16 4 13 13 1 9 11 2
16 3 10 0 9 11 11 15 3 3 1 9 1 9 12 13 2
27 11 11 13 0 9 0 0 9 2 15 1 9 11 11 13 0 9 3 1 10 9 9 11 1 12 9 2
20 1 11 15 1 11 13 11 11 7 11 2 11 11 2 9 11 7 11 11 2
31 14 9 13 1 15 2 16 0 0 9 11 11 2 11 2 1 11 2 10 0 9 2 13 3 13 0 0 0 9 11 2
17 0 0 9 1 15 13 7 13 1 3 0 9 1 0 0 9 2
24 9 11 13 1 9 12 0 9 0 11 2 15 13 13 1 9 10 9 1 9 11 1 11 2
30 9 9 1 12 9 2 11 2 11 12 2 12 2 12 2 12 2 2 11 2 11 12 2 12 2 12 2 12 2 2
5 3 7 3 13 9
5 15 15 1 15 13
5 3 7 3 13 9
23 16 9 1 9 0 9 7 9 13 9 0 2 9 11 11 0 9 10 9 1 0 9 2
29 2 1 0 9 13 0 9 0 0 9 7 0 9 1 12 9 0 9 7 15 15 13 2 15 13 2 2 13 2
19 10 9 15 13 1 0 9 2 3 7 2 3 0 2 12 9 3 13 2
22 2 13 1 0 9 2 9 13 13 13 1 9 9 2 15 13 13 1 9 15 0 2
24 13 3 13 3 9 9 2 16 4 1 12 9 3 15 3 13 3 1 9 2 2 13 9 2
31 9 1 9 2 15 13 0 0 9 1 9 2 3 9 2 10 9 15 13 1 0 9 1 9 0 7 0 9 2 9 2
16 13 2 16 10 9 13 9 2 7 1 0 0 9 15 13 2
22 0 9 13 0 9 1 0 9 2 7 3 15 13 2 1 9 9 3 3 3 13 2
30 16 9 13 1 9 9 9 9 2 3 1 9 15 13 13 9 7 9 2 3 3 0 2 1 0 9 1 10 9 2
32 3 1 9 1 9 7 9 2 1 9 7 9 2 13 13 0 9 2 16 7 14 9 2 7 7 9 7 9 13 0 9 2
5 12 9 1 12 9
11 9 0 9 11 15 13 1 2 9 2 11
24 16 10 9 1 12 1 9 0 9 11 3 3 13 2 15 15 1 0 9 13 14 1 0 2
14 0 9 14 13 7 16 15 13 2 3 1 9 13 2
22 7 15 1 15 9 1 0 9 13 0 9 0 9 2 9 11 11 11 2 12 2 2
29 2 1 9 12 2 16 4 13 1 9 1 9 1 11 2 4 13 9 1 11 2 15 4 3 13 12 2 12 2
17 3 13 7 1 11 7 3 1 11 13 3 3 12 9 2 2 2
14 2 13 2 16 12 9 1 15 12 13 1 11 15 2
8 1 11 13 1 3 0 9 2
10 0 13 0 3 1 12 7 12 9 2
11 15 13 2 16 1 11 3 15 3 13 2
10 13 0 2 10 9 1 15 13 9 2
7 15 3 13 0 9 2 2
6 2 16 1 9 13 2
6 2 13 1 9 2 2
9 2 9 9 2 7 1 10 0 2
13 2 3 13 13 10 9 2 16 13 15 0 2 2
14 2 14 13 0 2 16 1 11 13 9 11 2 2 2
6 2 3 15 15 13 2
15 1 9 1 9 2 15 13 0 11 2 4 15 3 13 2
20 13 2 10 4 15 1 15 13 9 2 16 4 15 13 9 9 1 0 9 2
26 1 11 13 7 11 2 11 7 9 2 15 13 1 11 1 11 2 9 9 11 2 14 2 11 2 2
12 2 13 4 9 2 15 1 9 13 1 9 2
10 13 1 9 2 7 15 13 0 9 2
14 2 16 15 13 12 2 13 4 15 1 9 1 9 2
14 1 9 15 9 13 2 16 4 13 15 16 0 9 2
11 14 15 13 13 1 10 9 16 0 9 2
7 3 4 15 13 0 9 2
17 15 7 9 4 13 9 9 2 7 3 3 15 15 3 13 2 2
12 2 10 4 10 9 9 1 10 12 9 13 2
21 2 4 15 13 2 7 13 15 3 15 0 2 15 4 15 13 1 0 9 2 2
17 2 7 1 0 9 1 11 1 11 4 1 9 15 13 2 2 2
17 2 1 9 15 9 13 15 13 2 15 13 3 0 9 10 9 2
11 3 4 15 15 1 0 9 3 13 2 2
11 2 13 4 15 1 9 2 15 13 0 2
15 2 13 4 15 3 1 9 2 7 16 3 13 0 9 2
10 13 2 1 15 15 15 3 13 2 2
8 2 3 3 15 9 13 9 2
17 2 9 3 1 15 13 9 7 9 15 1 10 9 3 13 2 2
6 2 13 0 0 9 2
3 2 0 2
14 13 1 9 1 9 9 2 13 3 1 0 9 2 2
13 2 13 1 0 0 9 1 0 9 0 10 9 2
11 2 13 2 13 0 9 7 3 0 9 2
13 13 15 2 7 16 4 15 13 12 2 12 2 2
5 2 10 13 9 2
5 2 14 3 9 2
9 7 13 2 16 13 0 9 2 2
3 9 2 9
5 9 12 2 9 2
7 9 1 11 14 1 0 9
2 11 2
24 0 9 13 1 15 2 16 4 9 9 1 0 9 0 9 11 4 3 13 14 1 9 11 2
48 2 0 9 1 15 13 13 14 1 9 2 16 4 13 9 15 0 9 1 0 9 2 2 13 9 9 11 11 11 2 15 3 9 11 13 16 9 9 9 11 1 9 1 0 9 1 11 2
21 11 2 11 13 2 16 1 9 1 11 13 0 15 13 1 0 0 9 1 11 2
2 11 2
30 0 9 9 1 0 9 11 7 0 9 9 9 11 7 11 3 1 9 11 13 9 0 7 0 0 9 7 0 9 2
14 1 0 0 9 15 13 1 0 9 9 9 11 11 2
47 1 0 9 2 9 0 9 1 0 9 11 11 0 2 7 0 9 13 1 9 1 0 9 9 3 0 9 2 15 13 1 15 2 16 3 0 2 0 7 0 9 13 1 0 9 0 2
3 9 1 11
5 11 2 11 2 2
18 12 9 2 9 1 0 0 9 0 9 2 4 13 9 0 0 9 2
7 13 1 15 3 10 9 2
43 13 3 3 2 16 0 9 9 10 9 3 3 13 3 0 0 9 0 9 2 9 11 2 11 2 11 7 11 2 11 2 1 15 13 4 9 1 0 9 1 11 13 2
19 9 11 11 11 13 2 16 4 0 9 13 1 9 9 13 10 0 9 2
12 9 15 7 13 13 9 9 1 11 3 3 2
15 1 0 12 13 3 11 12 9 2 1 12 0 13 9 2
7 3 0 9 13 0 9 2
12 10 9 13 9 0 9 13 10 9 1 9 2
14 9 0 9 3 1 9 4 13 13 0 9 9 11 2
14 1 15 13 9 13 9 0 2 15 4 13 0 9 2
2 0 9
2 11 2
21 9 9 0 9 0 3 11 2 11 7 11 4 13 4 13 2 0 2 9 11 2
12 13 15 3 9 0 9 11 1 11 11 11 2
14 1 15 4 10 12 9 10 9 3 13 7 1 9 2
2 0 9
24 9 1 11 7 11 1 0 9 13 0 2 13 1 0 9 9 9 11 11 11 1 0 9 2
44 9 13 2 16 12 9 15 1 0 9 1 11 13 2 16 1 9 1 0 9 4 13 2 16 4 13 0 9 2 15 4 13 0 13 0 9 9 1 0 9 7 0 9 2
11 2 10 9 13 2 2 13 11 2 11 2
12 1 9 9 11 13 13 10 0 9 11 9 2
26 2 13 15 2 16 13 0 13 0 9 2 15 4 4 13 9 2 15 13 12 9 2 2 13 3 2
15 0 9 1 11 13 1 15 1 0 9 10 9 0 9 2
32 9 1 0 9 13 3 7 3 7 13 1 9 9 0 9 2 13 15 1 0 9 0 9 11 2 15 15 13 1 0 9 2
15 0 9 11 13 0 9 1 0 7 1 0 9 0 9 2
3 9 11 11
2 11 2
21 9 9 2 3 13 13 1 0 9 0 9 2 1 11 11 1 9 13 10 9 2
16 0 0 2 9 15 3 13 1 9 1 11 7 0 2 9 2
33 13 2 16 9 1 15 2 16 4 13 1 10 9 1 9 9 11 2 13 2 16 4 15 9 9 9 1 9 13 10 0 9 2
9 2 13 13 9 0 15 1 9 2
15 13 1 15 2 7 1 9 9 9 2 2 13 11 11 2
32 13 2 16 15 1 9 9 9 13 1 15 2 16 4 9 13 4 13 12 9 9 2 16 1 9 9 4 13 14 0 9 2
14 2 1 10 9 13 0 0 9 0 9 9 7 9 2
16 9 4 13 14 1 0 9 7 10 9 2 2 13 11 11 2
2 9 9
7 11 1 11 2 11 2 2
40 0 9 2 1 15 1 0 12 9 4 1 9 0 9 13 1 0 11 12 9 7 13 12 0 9 2 12 9 7 12 0 9 2 13 1 9 9 0 9 2
16 3 3 13 9 0 9 9 11 11 11 2 9 4 3 13 2
19 9 13 13 0 0 9 0 9 1 11 2 15 1 9 13 3 1 12 2
15 1 0 9 3 13 1 12 9 9 1 9 12 9 9 2
3 0 0 9
6 9 1 0 2 9 2
9 11 11 2 9 9 1 11 9 11
5 11 2 11 2 2
15 1 0 0 9 1 9 0 9 13 11 11 3 0 9 2
42 1 0 9 0 9 1 9 0 9 4 13 9 11 11 1 0 2 9 2 11 11 2 10 0 9 4 13 0 9 11 11 2 7 0 0 9 9 11 0 9 9 2
11 10 9 9 13 0 0 9 0 12 9 2
8 10 0 0 0 9 13 4 2
29 3 13 13 2 16 1 9 1 0 2 9 2 11 11 15 13 10 9 9 1 9 13 1 0 2 9 2 11 2
25 0 9 0 9 2 7 2 12 0 9 2 1 12 0 9 13 9 9 0 12 9 1 10 9 2
14 3 15 13 1 3 12 9 1 11 7 12 1 9 2
8 12 0 9 4 13 1 11 2
21 1 0 9 11 11 11 11 11 13 14 0 2 16 0 9 0 9 13 1 11 2
38 1 10 9 13 7 15 2 16 14 11 3 13 0 9 1 10 3 0 0 9 7 9 1 0 9 2 15 4 13 1 9 13 9 0 9 11 11 2
6 9 9 1 9 0 9
17 0 9 0 0 9 1 0 9 13 1 9 9 11 10 0 9 2
20 3 3 2 16 9 4 13 1 9 9 9 2 9 9 0 9 10 9 13 2
16 9 9 11 11 11 2 11 2 15 13 2 16 3 9 13 2
26 3 0 9 11 9 11 9 2 11 2 13 2 16 15 15 9 13 2 7 13 3 1 9 0 9 2
33 3 4 15 3 13 2 15 0 9 9 0 9 11 9 1 9 13 7 13 15 14 3 2 16 15 15 13 2 7 10 9 2 2
40 0 0 9 15 13 2 16 2 0 0 9 2 2 0 0 0 9 2 15 10 9 13 7 13 1 11 1 0 9 2 2 16 4 15 9 13 15 13 2 2
15 10 9 11 4 15 3 13 2 15 9 0 9 3 13 2
16 11 11 2 11 2 2 2 9 0 0 9 15 15 13 0 2
6 13 10 3 0 9 2
19 3 0 9 9 2 9 1 9 9 7 0 9 1 9 0 7 0 9 2
16 13 15 2 16 4 10 9 13 2 16 4 4 3 13 2 2
16 13 4 15 11 0 2 9 9 11 2 9 11 2 11 2 2
18 1 3 0 9 9 11 4 13 4 3 13 9 0 9 11 1 11 2
19 15 4 4 13 9 10 9 1 0 9 11 7 3 4 13 1 10 9 2
20 13 15 3 2 3 2 16 4 4 13 9 9 11 2 9 1 0 9 13 2
23 2 9 1 0 9 11 4 15 13 3 1 10 9 2 7 15 9 9 11 11 11 11 2
22 16 13 2 13 15 1 9 9 2 16 9 1 15 2 16 4 15 13 9 2 13 2
25 15 13 3 9 2 16 7 9 9 9 11 11 13 2 16 1 10 9 13 9 11 11 1 11 2
15 13 15 1 15 7 1 0 9 2 3 2 1 0 9 2
22 13 2 16 9 11 13 9 7 11 2 7 13 1 15 2 3 1 9 0 1 11 2
8 13 9 11 2 15 13 2 2
3 15 1 11
1 9
3 15 1 11
17 3 0 9 1 9 0 0 9 1 11 4 13 13 1 0 9 2
30 0 0 9 2 11 2 0 9 13 2 16 0 9 9 1 0 9 13 2 16 11 13 4 13 1 9 1 0 9 2
19 3 11 13 2 16 16 9 0 9 9 1 11 4 13 0 0 9 11 2
33 13 15 3 3 0 2 13 1 0 9 11 4 13 3 0 9 2 15 4 1 15 3 13 13 7 9 1 9 0 1 10 9 2
15 9 3 13 2 7 9 0 9 2 3 9 9 2 13 2
28 0 9 13 3 0 9 9 7 9 11 11 2 15 1 9 1 9 0 9 13 2 16 9 9 0 9 13 2
36 0 9 9 1 11 13 2 3 7 1 9 0 0 9 11 2 15 13 2 16 10 9 13 0 13 15 1 0 0 9 2 16 3 3 0 2
28 2 0 9 7 13 3 13 2 3 1 9 4 3 1 0 9 11 9 9 13 0 9 1 9 2 2 2 2
12 0 9 4 9 11 13 3 9 9 9 9 2
18 7 3 7 1 15 13 9 2 13 3 14 0 13 1 0 0 9 2
8 11 13 1 10 9 0 9 2
19 10 0 9 3 11 1 10 0 9 3 13 1 9 9 2 15 13 9 2
14 14 9 3 13 13 2 10 9 1 9 10 9 13 2
10 7 3 13 9 13 3 12 0 9 2
31 0 9 3 0 9 13 7 13 1 9 2 3 4 13 3 0 2 3 0 9 9 2 13 4 15 4 9 0 9 2 2
26 13 3 2 16 11 2 3 3 0 2 15 3 1 9 9 13 13 1 3 0 0 9 1 0 9 2
22 7 3 0 9 0 9 15 3 13 10 0 9 2 7 9 3 3 13 1 10 9 2
36 7 15 13 1 0 9 9 9 2 12 1 15 13 7 1 0 11 2 2 3 13 0 9 9 2 7 3 0 9 13 10 9 1 0 9 2
6 14 16 15 13 11 2
12 9 3 1 9 3 13 3 1 0 0 9 2
16 1 9 11 4 7 0 9 13 3 13 7 9 1 15 0 2
5 0 9 1 9 9
5 11 2 11 2 2
32 16 13 3 9 0 9 9 12 2 0 1 9 9 1 9 0 9 0 0 9 1 0 11 2 0 9 15 13 13 10 9 2
14 13 15 15 3 9 9 9 1 11 1 11 11 11 2
20 1 15 15 9 13 7 9 13 7 0 9 2 9 9 1 9 1 9 9 2
15 1 11 3 13 12 0 9 9 7 0 13 13 12 9 2
9 9 1 15 1 9 9 12 13 2
37 3 15 13 9 9 0 9 1 11 11 11 2 9 1 15 13 3 0 7 0 2 2 13 15 13 2 16 4 15 1 9 9 13 9 9 2 2
5 11 11 13 1 11
36 9 9 11 11 2 0 1 0 9 9 2 13 3 1 9 9 1 9 1 9 11 2 11 2 2 15 4 13 13 11 0 9 1 0 9 2
25 9 13 9 3 13 2 16 0 9 13 13 7 9 9 1 12 9 9 13 13 14 1 12 9 2
10 13 15 15 3 0 9 11 11 11 2
29 1 15 13 9 9 1 9 1 9 0 9 1 11 11 2 0 9 11 2 2 1 11 13 9 9 11 11 11 2
25 13 7 13 0 9 9 1 0 9 7 13 9 1 9 2 1 15 4 13 14 12 1 12 9 2
13 15 0 1 10 9 13 2 2 13 15 11 11 2
3 9 1 9
5 11 2 11 2 2
28 1 9 1 9 0 9 13 1 9 12 9 1 12 1 12 9 2 15 13 1 0 9 9 1 11 1 11 2
17 9 2 13 1 9 9 9 2 1 0 9 13 9 9 1 9 2
24 9 13 1 9 2 13 9 2 13 9 7 1 0 9 13 0 9 1 15 13 9 12 9 2
19 12 1 0 9 15 1 9 13 3 1 9 3 1 0 9 1 0 9 2
21 16 15 1 9 1 9 13 9 9 2 9 13 0 0 9 7 13 9 1 9 2
6 9 16 0 0 9 2
5 11 2 11 2 2
19 0 9 9 0 9 11 7 11 1 9 11 15 13 3 3 1 9 11 2
23 13 15 1 15 1 9 0 9 3 1 9 1 9 9 9 7 0 9 2 15 9 13 2
29 9 11 11 11 15 1 9 13 2 16 11 7 11 13 0 3 13 1 0 9 9 1 9 2 7 1 15 13 2
21 16 13 1 12 0 9 2 11 7 11 15 13 2 7 1 9 1 15 4 13 2
29 11 11 3 13 2 2 4 3 13 9 11 11 11 2 16 13 2 16 4 15 13 2 16 13 0 13 9 9 2
19 15 4 14 13 3 2 16 13 0 13 9 2 3 15 13 1 0 9 2
19 7 3 4 15 1 11 13 1 15 2 16 16 9 13 2 13 13 2 2
21 9 11 2 11 7 11 13 3 1 15 2 16 13 9 0 9 9 10 9 9 2
8 3 7 10 9 11 3 13 2
3 9 1 9
6 0 11 2 11 2 2
15 3 0 9 0 9 9 11 13 3 9 11 1 0 11 2
21 3 4 1 11 13 12 10 9 2 15 1 9 9 11 0 13 9 13 1 9 2
14 0 9 13 7 3 1 9 7 9 4 13 3 13 2
2 9 9
6 0 11 2 11 2 2
16 0 0 9 1 0 11 13 1 0 9 10 9 9 9 9 2
13 9 9 13 0 9 1 12 0 9 1 0 11 2
26 2 1 9 13 1 10 9 1 9 12 2 2 12 2 9 2 2 13 3 9 9 0 11 11 11 2
24 2 1 0 9 3 13 9 0 9 2 7 7 3 13 3 13 9 9 2 15 13 9 9 2
10 9 4 14 1 9 0 9 13 2 2
21 1 9 9 0 9 0 9 1 0 11 11 11 4 1 9 13 12 9 1 9 2
24 2 13 4 3 7 0 9 2 7 13 13 2 16 15 10 9 15 13 3 1 10 12 9 2
18 13 0 9 1 12 12 0 11 2 7 7 13 9 7 1 0 9 2
14 3 15 7 3 13 9 9 1 0 9 9 9 2 2
3 9 4 13
5 11 2 11 2 2
16 9 9 0 9 11 2 9 4 7 1 0 9 0 9 13 2
15 0 9 12 9 9 13 9 13 1 0 0 7 0 9 2
54 9 2 11 11 1 0 9 3 13 2 16 1 9 9 15 13 13 9 2 16 0 9 0 2 0 11 2 13 0 13 0 9 0 9 9 2 2 3 0 9 9 11 2 2 15 13 3 0 9 1 9 0 9 2
36 1 10 9 2 1 15 13 13 1 0 9 9 0 9 9 0 9 2 13 10 9 9 2 11 11 3 9 2 0 7 0 9 2 10 9 2
3 3 13 2
2 9 2
9 1 11 13 3 2 3 3 9 2
14 0 9 12 7 12 2 0 0 12 7 12 9 11 2
7 2 1 11 3 7 3 2
14 0 9 12 7 12 2 0 12 7 12 9 11 2 2
15 1 9 9 13 1 12 2 12 7 13 1 12 2 12 2
15 9 13 1 9 1 12 2 12 7 13 1 12 2 12 2
3 9 9 2
16 0 9 12 9 11 13 1 9 12 2 0 12 1 9 12 2
8 0 0 9 13 12 9 11 2
3 0 9 2
10 0 9 13 0 2 0 2 9 0 2
5 0 9 2 11 2
5 1 0 9 14 9
5 11 2 11 2 2
14 12 9 0 9 0 9 0 9 9 11 11 3 13 2
17 1 9 12 0 9 0 1 0 9 15 14 1 9 0 9 13 2
18 9 9 2 16 13 1 9 1 0 9 2 13 0 9 1 12 9 2
20 3 0 9 3 13 2 16 15 13 3 0 9 7 9 2 1 10 0 9 2
24 13 15 3 14 13 2 16 13 1 0 9 0 9 2 15 1 9 13 3 1 9 10 9 2
34 11 2 15 4 1 9 9 13 1 9 1 9 2 15 3 13 2 16 4 15 13 1 11 2 3 13 9 9 9 2 0 0 9 2
2 11 3
5 11 2 11 2 2
34 0 9 1 12 0 9 13 12 0 9 1 11 1 0 9 1 11 1 11 7 13 2 16 3 10 9 13 1 0 0 9 11 11 2
24 9 13 7 1 0 9 0 11 3 3 13 0 9 1 9 2 15 13 1 0 12 0 9 2
19 9 3 13 1 9 13 12 9 7 10 9 15 3 13 0 9 1 11 2
1 9
7 7 13 15 9 2 2 2
16 0 9 11 3 13 9 11 13 0 9 9 1 11 7 9 2
24 1 3 2 0 2 13 0 13 9 2 15 15 1 15 13 7 15 13 1 9 0 9 11 2
9 1 9 4 13 4 13 9 11 2
28 7 16 7 9 13 0 7 13 15 9 9 11 2 16 9 13 10 9 1 9 13 2 9 3 13 3 3 2
9 9 11 3 1 0 9 3 13 2
11 13 15 15 2 15 13 9 1 9 9 2
5 15 15 3 13 2
8 1 9 15 13 13 10 9 2
11 3 13 9 2 7 9 1 15 4 13 2
19 1 0 9 9 1 11 10 0 9 3 13 0 9 10 9 1 9 9 2
28 15 2 16 10 9 0 9 13 2 15 13 13 14 0 9 9 11 2 15 3 3 3 0 9 1 9 13 2
2 11 13
5 11 2 11 2 2
36 9 11 11 11 2 11 2 13 9 2 3 4 13 10 9 9 11 11 1 9 9 11 2 16 15 1 0 9 11 1 9 11 2 11 13 2
13 11 2 11 13 3 0 9 1 0 9 9 9 2
5 0 9 1 12 9
9 9 0 2 13 3 7 3 13 13
5 11 2 11 2 2
25 2 13 3 7 3 13 13 2 13 13 7 3 13 3 2 3 15 13 0 2 13 0 0 9 2
7 10 9 13 0 9 13 2
7 0 9 13 0 9 2 2
24 10 9 13 1 9 11 9 11 0 2 11 2 2 16 3 13 0 9 9 11 1 0 9 2
17 0 9 3 13 12 9 9 2 15 9 13 9 1 10 0 9 2
33 13 15 1 0 9 9 1 12 2 1 12 0 2 0 9 1 15 2 16 0 4 1 12 2 9 13 7 10 9 13 1 9 2
14 10 2 0 2 9 13 1 11 2 11 1 9 9 2
13 9 2 15 15 9 13 2 3 3 13 0 9 2
14 9 1 9 9 9 4 13 13 0 9 9 0 9 2
16 0 9 2 1 15 13 0 9 9 2 4 13 1 12 9 2
36 13 1 15 14 1 9 3 9 9 2 15 3 13 9 9 2 0 9 9 9 0 7 0 9 1 10 9 7 13 1 0 9 11 7 11 2
17 9 11 11 1 9 9 11 13 9 9 1 9 9 1 0 9 2
22 1 15 4 11 13 1 9 13 2 16 4 1 12 2 9 13 9 15 9 9 11 2
25 11 4 13 3 13 2 16 4 1 12 2 9 11 9 13 9 9 9 1 0 7 0 9 9 2
18 1 12 2 9 4 3 9 13 13 9 9 12 9 1 9 10 9 2
23 9 1 11 11 11 1 0 9 9 1 9 13 2 2 13 2 16 3 13 9 13 9 2
16 15 3 4 4 1 11 13 3 2 16 4 13 0 9 11 2
25 16 15 15 13 2 16 4 4 13 3 2 16 4 13 9 0 11 2 3 15 15 15 13 2 2
27 9 9 15 3 3 13 1 9 9 1 9 9 9 7 12 0 9 1 9 1 9 0 0 0 9 9 2
19 16 15 9 4 0 9 9 13 2 13 9 1 9 9 1 9 10 9 2
9 1 9 9 10 9 9 11 13 2
6 9 0 2 9 13 9
7 9 13 9 1 0 9 9
5 11 2 11 2 2
57 9 9 0 9 7 0 9 1 9 0 9 11 2 7 15 3 1 9 0 9 2 9 2 0 2 0 2 0 2 0 9 2 3 2 7 0 9 0 9 2 9 2 9 7 9 9 2 13 0 9 0 9 1 12 2 9 2
34 1 12 2 9 11 9 3 13 9 11 9 9 9 1 0 7 0 9 9 7 1 0 9 9 9 1 9 1 9 1 9 0 9 2
31 10 9 0 9 11 11 1 9 11 13 9 9 2 15 9 13 1 9 10 0 0 9 1 9 9 1 9 1 0 9 2
22 9 13 11 9 1 0 9 9 11 0 12 2 9 2 15 4 13 1 9 0 9 2
37 3 9 11 0 2 11 2 9 13 2 16 2 13 3 7 3 13 13 2 13 13 7 3 13 3 2 3 15 13 0 2 13 0 0 9 2 2
10 3 13 2 10 9 13 0 9 13 2
6 0 9 13 0 9 2
17 13 15 3 1 12 9 9 2 15 9 13 9 1 10 0 9 2
33 13 15 1 0 9 9 1 12 2 1 12 0 2 0 9 1 15 2 16 0 4 1 12 2 9 13 7 10 9 13 1 9 2
2 9 12
2 9 12
2 12 9
2 0 9
1 9
4 12 2 9 12
2 0 9
4 11 3 1 11
3 9 2 12
2 0 9
4 9 13 0 9
9 3 12 9 1 9 11 13 0 9
15 1 11 3 4 12 2 12 2 13 9 0 9 1 9 2
26 13 4 1 15 1 9 9 0 11 11 2 15 13 3 2 16 4 13 1 0 9 0 9 1 11 2
27 1 9 0 9 13 2 16 9 9 11 13 0 7 0 13 7 9 2 15 15 1 0 9 13 10 9 2
11 9 11 11 13 9 1 9 9 1 9 2
26 3 12 2 12 2 12 4 13 0 9 0 9 11 2 11 2 7 9 9 2 0 9 11 2 11 2
19 9 4 13 1 9 0 9 1 0 9 1 11 2 3 7 13 9 9 2
13 3 13 7 0 9 2 3 15 9 13 1 9 2
17 9 13 13 1 0 9 1 11 2 0 1 11 7 0 9 11 2
13 15 13 9 12 2 9 2 3 4 13 0 9 2
58 16 0 9 0 9 0 9 2 11 9 13 1 0 9 2 16 11 2 11 2 9 9 12 2 12 2 12 13 0 9 0 9 1 9 9 0 0 9 2 16 1 0 9 0 9 11 2 15 0 9 13 0 0 2 11 2 11 2
15 3 15 13 2 16 9 0 9 13 15 9 0 9 11 2
32 1 9 9 11 10 9 13 9 2 16 4 0 9 13 13 1 9 0 9 0 9 1 3 0 2 7 15 1 10 0 9 2
20 9 11 13 9 2 16 15 1 10 9 13 1 9 7 13 15 1 0 9 2
18 3 4 15 13 2 0 9 3 13 7 9 13 1 0 9 1 11 2
44 9 1 9 1 9 9 4 1 9 11 9 2 9 0 9 1 11 13 3 0 9 11 2 16 9 13 13 9 0 7 0 9 2 16 3 0 9 13 9 1 9 15 2 2
31 1 1 15 2 16 9 9 11 11 15 1 9 13 13 10 9 2 13 4 15 3 1 9 9 1 11 9 2 11 11 2
26 13 15 2 3 9 13 3 1 0 9 7 3 3 3 1 11 13 2 16 15 9 13 1 0 9 2
17 2 9 11 3 13 9 13 2 7 0 9 13 1 9 0 9 2
24 1 0 9 15 13 9 1 9 2 3 15 9 13 1 15 2 1 9 0 9 1 12 9 2
9 10 9 4 13 9 1 9 2 2
8 1 9 11 11 13 12 9 2
13 0 9 9 13 3 1 11 7 9 13 0 9 2
12 1 10 9 4 15 13 9 12 7 12 9 2
24 13 15 7 13 7 9 2 16 11 11 4 1 10 9 13 9 1 9 9 1 9 0 9 2
10 3 4 15 13 9 0 9 3 13 2
9 1 0 9 15 13 0 0 9 2
15 0 9 13 9 0 9 7 13 1 9 9 1 0 11 2
12 0 9 4 1 11 11 13 13 1 12 9 2
18 1 10 9 4 13 14 0 11 2 11 2 2 7 7 0 9 0 2
7 13 7 2 15 4 13 2
18 3 4 15 13 1 11 2 0 9 13 9 9 15 9 9 1 11 2
15 1 9 9 9 9 2 11 11 7 13 13 1 9 9 2
21 15 13 13 14 0 9 2 7 14 1 9 9 1 11 2 3 3 3 13 9 2
13 1 10 0 0 2 9 9 11 13 9 1 9 2
10 13 2 16 0 9 13 1 12 9 2
21 2 7 9 15 13 3 12 9 7 3 1 0 9 3 13 3 1 0 9 2 2
36 9 9 0 9 15 9 9 11 11 13 3 2 2 2 1 0 9 3 15 13 0 9 9 7 13 13 2 16 1 0 9 4 13 3 3 2
10 7 4 13 9 1 9 0 9 2 2
21 11 11 2 9 9 0 11 1 11 2 7 10 9 11 3 13 9 9 3 11 2
36 0 9 2 9 1 11 1 12 9 2 13 11 2 11 1 11 2 0 9 9 11 11 11 2 11 1 11 7 0 9 11 2 11 1 11 2
1 9
2 9 12
6 12 9 2 9 2 9
4 12 9 2 9
3 12 9 9
5 12 13 15 2 13
2 12 9
4 12 1 9 9
2 12 11
3 12 9 9
5 9 1 12 1 12
3 12 9 9
6 12 11 1 2 0 9
7 1 9 2 9 2 9 9
3 12 0 9
7 12 11 13 2 13 2 13
6 12 9 2 9 2 9
3 12 0 9
4 12 13 2 13
2 12 9
3 12 9 11
7 12 11 11 2 12 2 2
4 12 9 1 0
7 12 13 2 15 15 13 2
2 12 9
4 12 9 2 9
6 12 0 9 12 1 12
5 12 3 3 13 15
2 12 9
3 12 9 9
1 11
2 12 9
3 12 13 15
3 12 9 0
5 12 1 0 0 9
4 12 9 7 15
5 9 1 12 1 12
3 12 9 11
2 12 9
6 12 0 2 0 2 11
4 12 9 0 9
5 12 0 9 2 9
3 12 9 11
3 12 9 11
3 12 13 15
8 12 0 9 11 2 12 2 2
4 12 9 1 9
2 12 9
4 12 9 9 11
3 12 9 11
3 12 9 11
3 12 9 9
2 9 12
3 12 9 11
2 12 9
3 12 9 11
3 12 0 0
6 12 3 13 2 13 9
3 12 11 9
3 12 9 11
4 12 11 0 11
3 12 9 11
2 12 11
4 12 0 9 11
3 12 9 11
2 12 11
4 12 0 9 11
4 12 9 1 9
3 12 0 9
3 12 9 9
10 12 9 2 9 2 13 15 2 2 2
4 12 11 2 11
5 12 11 2 0 9
2 12 11
3 12 9 11
2 12 11
2 12 9
2 12 9
3 12 9 11
3 12 11 9
6 12 9 2 12 2 2
4 12 11 12 2
4 12 9 11 11
6 12 9 7 9 1 11
4 12 0 9 9
3 12 0 9
4 12 11 2 11
4 12 0 9 11
3 12 9 11
4 12 0 9 11
3 12 9 11
5 3 9 1 9 2
13 2 13 1 0 9 13 9 9 9 1 9 9 2
29 3 1 10 9 13 1 0 9 0 9 3 1 9 0 0 9 7 11 2 2 13 15 3 0 9 9 11 11 2
11 9 4 3 13 13 13 9 9 1 15 2
31 3 4 15 13 13 9 2 3 3 13 3 0 9 3 2 0 2 9 9 1 0 9 0 0 9 1 0 2 0 9 2
7 11 4 3 13 9 9 2
17 0 9 13 3 9 0 11 2 15 15 13 13 1 15 1 11 2
31 2 16 4 0 9 1 10 9 13 3 14 0 9 7 13 15 0 2 13 4 15 3 13 0 2 0 9 7 3 13 2
18 7 13 9 9 13 7 13 4 1 10 9 3 2 2 13 9 11 2
12 1 9 9 1 11 7 11 13 7 0 9 2
30 2 1 9 2 16 11 0 9 3 13 2 13 7 1 9 3 2 2 13 9 9 9 0 9 7 0 9 11 11 2
14 0 9 4 1 9 9 13 3 13 9 1 0 9 2
10 1 0 9 0 11 3 10 9 13 2
10 9 9 13 11 13 1 2 9 9 2
2 11 2
26 1 9 12 2 3 13 0 9 2 15 0 11 0 1 11 13 1 2 9 9 2 3 1 9 11 2
18 9 9 2 0 3 1 2 9 2 0 11 2 13 9 1 0 9 2
8 9 1 0 0 9 13 9 2
21 9 7 13 0 9 16 9 0 9 7 1 15 7 0 9 2 0 2 0 9 2
15 1 9 9 15 13 1 11 9 9 9 1 11 1 9 2
34 13 15 2 9 2 2 15 0 9 1 9 1 11 1 11 13 7 13 15 3 1 3 12 0 0 9 1 0 9 1 3 0 9 2
16 3 1 9 3 1 11 13 13 9 1 12 9 3 0 9 2
39 12 9 3 13 1 11 9 2 16 10 9 13 3 3 2 3 15 13 0 9 7 13 1 9 1 0 9 1 0 9 16 11 2 3 7 1 0 9 2
33 0 9 0 0 9 1 11 11 11 13 2 16 1 9 0 9 9 0 2 9 2 0 3 1 12 2 13 2 7 3 15 13 2
18 9 13 0 9 7 9 0 9 1 9 1 9 9 9 7 9 9 2
25 0 9 13 1 11 9 0 1 0 9 2 15 15 3 13 14 11 2 7 7 11 7 0 11 2
14 3 15 13 3 13 2 7 13 15 13 3 1 9 2
17 3 13 3 0 7 16 15 1 15 13 2 13 15 0 0 9 2
13 15 7 13 13 1 0 9 1 9 10 12 9 2
18 0 9 13 0 9 0 1 9 9 1 0 9 7 9 1 0 9 2
18 1 9 12 13 1 0 9 9 1 11 16 12 1 9 9 0 9 2
23 3 11 1 10 9 13 12 9 2 16 14 9 9 13 1 11 7 1 12 9 1 11 2
42 3 9 1 0 9 13 1 9 1 0 9 2 7 9 13 3 0 7 13 9 1 9 11 7 9 10 9 2 16 9 13 3 1 0 9 12 7 12 9 1 9 2
20 0 9 7 0 9 15 3 13 9 2 3 10 9 13 7 3 13 0 9 2
20 9 13 1 9 0 0 9 2 7 3 1 3 0 0 9 2 15 13 11 2
12 0 0 9 3 4 3 3 13 2 3 3 2
26 11 11 1 0 9 1 0 11 13 1 0 9 0 9 0 0 9 2 15 13 1 0 9 9 13 2
14 0 9 9 7 0 9 1 0 9 13 9 7 9 2
19 2 0 2 0 9 2 16 13 1 9 9 2 3 3 9 0 9 13 2
23 0 9 13 0 9 7 13 1 9 3 9 2 15 3 13 7 1 0 9 2 13 11 2
20 9 1 9 13 7 9 2 16 15 1 0 7 0 9 13 0 9 9 9 2
8 0 9 9 11 1 0 9 2
7 13 15 1 11 9 11 2
19 13 3 1 9 2 10 9 7 13 1 0 2 0 2 9 1 0 9 2
11 9 1 0 9 9 13 7 0 9 7 9
2 11 2
5 13 15 0 9 2
3 13 9 2
5 4 13 1 9 2
25 3 13 13 10 9 0 9 2 15 13 1 0 9 0 9 1 12 9 9 0 9 1 0 9 2
9 0 9 13 9 10 12 0 9 2
13 9 13 4 13 9 9 2 1 9 1 0 0 9
19 2 0 2 9 13 3 9 2 9 2 0 9 2 9 9 7 0 9 2
8 9 15 13 1 9 13 9 2
22 1 9 4 13 7 9 7 9 2 9 7 1 15 13 4 13 9 7 3 0 9 2
4 9 0 9 2
3 0 9 2
20 1 10 9 4 11 13 1 9 12 13 0 9 2 15 4 13 0 0 9 2
3 0 9 2
19 9 11 4 13 13 0 0 7 0 9 2 15 4 15 13 1 9 9 2
12 1 9 12 4 11 13 13 13 0 0 9 2
3 0 9 2
28 1 9 0 9 9 4 11 13 0 9 1 9 9 2 9 2 9 2 9 9 2 9 1 9 9 7 9 2
3 0 9 2
12 10 9 4 1 9 0 9 13 7 0 9 2
4 9 1 9 2
15 4 13 0 9 1 9 9 1 9 2 15 13 9 11 2
8 9 9 1 9 11 13 0 2
2 9 2
24 0 9 9 13 0 9 9 1 15 0 9 7 1 9 12 7 0 9 7 9 13 1 9 2
5 1 11 13 14 15
4 11 2 9 9
15 0 0 9 1 11 13 0 7 3 9 2 16 0 9 2
16 13 1 15 2 16 1 15 4 13 3 14 12 12 0 9 2
25 9 13 3 13 14 9 1 0 9 2 3 15 2 15 3 13 1 9 12 2 7 10 9 2 2
29 9 11 2 16 0 9 15 13 3 11 3 3 2 0 2 1 11 7 3 2 13 0 7 3 4 13 0 9 2
19 13 14 1 11 2 1 15 12 0 9 15 13 13 1 9 9 1 9 2
25 11 13 1 11 3 12 9 2 11 1 11 14 9 2 16 1 0 9 9 13 11 1 9 2 2
16 3 2 13 2 13 11 2 3 13 11 7 11 1 12 9 2
19 11 1 11 13 0 1 0 9 1 9 2 3 15 7 13 13 0 9 2
3 13 15 2
5 3 15 9 13 2
9 14 2 15 9 15 13 14 3 2
27 7 13 13 14 1 11 2 11 3 13 1 9 0 9 1 11 2 16 15 11 13 9 1 0 0 9 2
41 13 4 0 2 7 3 0 2 16 4 15 11 2 15 15 13 0 9 1 10 9 1 9 2 13 12 9 13 9 9 0 9 1 11 2 1 11 7 1 11 2
25 3 4 15 1 0 9 2 15 11 13 1 9 1 9 11 1 0 0 9 2 13 3 0 9 2
3 11 13 4
2 11 2
3 11 13 4
2 11 2
16 9 13 0 0 9 11 0 9 13 9 0 0 9 11 11 2
23 1 9 1 9 11 13 2 16 2 13 10 9 9 0 0 9 11 2 13 0 0 9 2
27 0 9 13 11 2 15 15 13 1 0 9 1 12 9 2 3 1 9 2 16 1 15 9 13 0 9 2
7 0 9 13 1 0 11 0
22 0 0 9 9 0 9 13 0 9 2 15 4 13 1 9 13 13 3 1 9 12 2
18 15 7 13 13 3 1 9 2 16 1 9 0 9 13 0 0 9 2
17 9 10 9 2 16 10 9 13 4 2 3 13 9 1 0 9 2
15 1 9 0 0 9 1 15 9 7 13 11 3 3 3 2
12 9 13 3 1 0 0 9 7 1 9 9 2
20 16 3 4 13 10 9 2 1 11 1 9 4 3 13 1 3 0 0 9 2
13 11 13 7 10 9 3 13 9 1 3 0 9 2
16 15 13 0 13 9 11 2 15 4 3 13 1 9 0 9 2
33 1 9 2 15 13 11 2 4 10 0 9 13 1 0 12 9 9 2 12 9 13 3 12 9 2 13 1 9 12 1 12 12 2
21 0 9 13 3 0 9 10 10 9 2 11 3 13 3 12 9 2 11 12 9 2
24 1 15 0 11 2 1 15 13 0 12 9 2 13 9 1 0 9 2 15 1 0 9 13 2
19 13 7 3 0 2 16 15 11 13 1 9 12 13 0 9 13 15 11 2
46 1 0 15 0 9 7 0 9 1 0 9 2 3 15 9 9 1 9 13 3 9 2 13 3 7 0 9 3 3 0 13 0 9 7 13 3 0 9 1 9 10 0 9 1 11 2
8 2 0 11 13 1 0 9 2
8 15 4 15 13 13 1 9 2
20 7 16 13 13 9 11 2 3 3 13 0 2 2 13 3 0 9 11 11 2
22 0 9 9 3 3 0 7 9 0 9 13 7 9 0 0 9 2 11 2 0 9 2
28 1 9 2 3 4 11 13 2 10 0 9 11 7 11 13 2 16 0 9 13 15 1 0 0 7 0 9 2
24 15 7 3 1 9 1 0 9 1 11 13 1 9 2 15 9 13 9 0 9 1 10 9 2
3 7 9 2
33 9 1 9 9 0 11 3 7 3 13 4 2 9 15 7 3 13 13 0 9 2 15 4 9 1 9 13 1 9 1 9 9 2
29 9 0 11 1 9 4 13 13 0 9 9 7 9 13 1 0 9 1 3 0 9 2 3 0 0 2 14 2 2
10 0 9 13 0 2 14 9 13 3 0
1 9
25 11 13 1 9 14 0 9 7 15 2 14 2 13 2 16 15 13 2 13 16 2 3 14 2 2
29 16 7 13 3 0 3 7 9 2 15 0 11 1 9 1 9 13 7 3 13 2 13 15 3 9 9 1 9 2
8 9 13 3 0 9 1 9 2
25 13 7 2 7 16 15 13 9 16 0 9 2 13 3 3 1 15 13 7 9 2 1 15 13 2
15 9 9 13 2 16 9 9 9 13 0 2 7 3 0 2
23 7 0 13 3 9 2 1 15 0 9 13 10 9 1 9 2 7 9 2 3 3 13 2
17 11 13 13 9 1 9 3 1 9 2 3 1 15 13 0 9 2
31 9 0 9 2 1 15 9 13 0 9 2 7 0 0 0 9 13 9 13 15 3 0 9 7 3 13 1 9 9 9 2
25 9 1 0 9 13 3 12 9 0 9 1 9 2 0 9 2 9 7 9 2 9 1 15 9 2
33 0 0 9 13 1 9 2 11 13 0 9 1 9 1 9 12 2 7 15 13 13 3 2 13 15 7 1 9 0 9 1 11 2
24 0 0 9 15 3 13 3 7 1 15 2 16 13 11 1 10 9 2 7 16 13 9 0 2
27 15 15 7 13 14 1 0 2 1 0 0 9 13 13 0 9 2 1 15 13 9 13 2 0 7 0 2
10 13 15 2 16 0 13 15 9 9 2
13 16 15 1 15 9 0 9 13 2 13 9 13 2
14 16 9 1 9 4 13 3 1 0 9 2 13 0 2
19 0 13 2 16 4 9 13 9 0 11 2 15 3 10 9 7 9 13 2
4 11 13 0 9
2 11 2
2 11 2
10 9 0 9 3 13 9 1 0 9 2
21 1 0 9 13 1 9 2 0 9 0 9 1 9 9 9 1 9 0 9 2 2
9 13 15 2 16 13 1 0 9 2
17 11 3 13 13 0 0 9 2 16 4 13 0 9 1 0 9 2
19 11 13 9 14 10 9 2 15 13 1 9 1 9 12 2 7 10 9 2
8 9 0 9 1 9 9 1 11
36 1 15 9 1 9 9 1 11 7 1 9 9 2 16 15 1 11 13 9 0 9 2 13 13 1 0 9 2 1 10 9 13 9 11 0 2
36 13 14 1 15 13 11 9 2 16 4 3 3 13 10 0 9 1 0 11 2 7 3 1 15 13 0 9 1 0 11 2 15 13 3 0 2
21 0 9 11 9 1 10 0 9 1 9 9 13 2 16 9 0 9 13 3 0 2
23 1 9 9 9 3 13 9 0 9 7 0 0 9 0 9 2 3 0 0 9 10 9 2
2 0 11
10 11 3 13 12 9 2 7 14 9 2
18 10 9 1 0 9 11 13 2 16 4 15 0 9 13 3 1 9 2
31 13 15 7 0 2 3 3 13 9 9 2 15 13 13 9 2 16 4 13 0 9 3 3 2 13 2 14 11 10 9 2
29 9 12 0 9 0 9 15 1 10 0 0 9 4 13 14 13 1 10 0 9 2 7 4 15 13 3 3 13 2
23 9 0 9 15 13 3 13 0 0 9 1 9 1 0 11 2 7 15 9 0 9 11 2
2 0 11
16 0 9 0 9 0 9 13 1 9 0 9 3 9 1 9 2
31 0 9 1 0 9 7 9 7 3 1 15 0 9 11 3 13 2 3 0 13 1 15 9 11 9 3 0 9 1 9 2
10 0 9 0 9 3 13 3 3 13 2
18 0 13 2 16 4 13 0 9 2 7 9 13 9 9 1 10 9 2
18 16 0 11 0 9 0 9 13 2 10 3 0 9 15 13 10 9 2
18 3 13 9 2 7 3 0 9 2 7 16 12 9 13 1 0 9 2
9 0 9 9 7 3 10 9 13 2
1 11
6 2 0 9 13 0 2
4 11 13 10 9
2 11 2
26 15 9 1 9 0 9 1 11 1 9 12 13 1 15 0 0 9 11 11 7 0 0 9 11 11 2
14 3 15 3 13 9 0 9 2 15 15 13 0 9 2
22 11 7 13 2 16 13 7 3 13 2 16 0 9 13 0 7 13 9 1 0 9 2
19 2 16 9 1 15 13 9 7 9 2 14 15 13 1 15 2 2 13 2
8 1 9 0 9 13 14 3 11
2 11 2
14 2 0 9 13 1 0 9 7 13 15 14 0 9 2
7 1 15 13 10 9 13 2
17 13 15 0 9 1 9 2 0 9 1 0 0 9 2 11 11 2
19 2 11 3 13 10 0 9 7 1 9 10 9 13 11 2 2 13 9 2
40 0 0 9 3 3 13 2 16 13 1 0 9 11 1 9 0 9 9 11 1 0 9 2 1 15 13 10 9 1 11 11 11 13 9 1 0 9 1 11 2
38 1 0 16 1 0 11 13 9 0 9 1 11 9 0 9 7 0 0 0 9 2 11 2 11 11 1 9 2 15 13 13 1 0 9 0 9 11 2
13 13 7 2 16 0 9 2 13 9 0 9 2 2
4 9 13 0 9
2 11 2
3 0 11 2
33 14 1 9 13 1 0 9 3 1 0 11 11 2 15 13 12 9 1 9 2 15 15 13 9 7 3 15 13 13 9 7 9 2
19 1 9 13 3 1 9 2 16 9 13 1 0 9 2 16 13 0 9 2
11 1 11 13 9 9 11 11 1 9 3 13
2 11 2
28 1 9 9 12 0 9 2 1 3 0 11 2 13 3 1 0 11 9 3 0 9 1 9 1 9 9 11 2
8 9 13 0 9 9 11 11 2
18 1 9 9 11 1 9 1 9 9 13 0 9 9 9 9 1 11 2
18 10 9 13 13 9 1 9 1 9 9 2 9 7 9 9 7 9 2
38 9 9 11 2 11 7 11 13 0 9 2 1 15 13 1 0 9 9 0 9 13 1 9 0 9 3 1 0 11 7 13 0 7 0 9 0 9 2
24 1 0 9 0 9 9 13 3 9 0 9 11 11 2 15 13 3 1 0 9 1 9 11 2
5 9 1 9 2 2
37 3 0 9 9 1 9 9 13 1 0 9 9 1 0 0 9 2 16 1 9 1 11 13 1 12 1 0 12 9 9 1 9 3 12 9 9 2
4 9 1 9 2
20 3 16 9 9 1 0 9 13 3 3 9 2 16 1 0 0 9 13 9 2
9 0 9 15 13 1 12 9 9 2
5 1 11 13 12 9
5 0 9 3 13 4
2 11 2
24 16 1 0 9 13 1 11 1 9 1 9 0 9 2 0 9 13 1 0 9 0 9 11 2
19 1 9 0 9 15 3 13 9 11 7 9 2 15 13 1 9 0 9 2
17 0 9 1 9 1 0 9 3 13 13 0 9 1 9 0 9 2
18 0 9 4 13 3 1 9 11 1 9 9 0 11 2 9 7 11 2
28 0 9 13 2 16 1 0 0 9 0 9 13 1 11 12 9 7 16 4 13 9 1 9 9 2 9 2 2
15 0 9 9 3 13 1 9 12 0 9 3 0 9 11 2
5 11 11 13 1 11
7 9 1 9 13 2 11 13
3 0 11 2
43 0 9 13 0 9 9 9 11 1 9 9 0 9 11 2 0 9 1 9 1 11 7 9 9 1 0 7 0 9 1 0 11 13 0 9 0 12 2 9 0 9 11 2
11 0 9 3 13 1 10 9 1 10 9 2
32 11 11 15 13 13 9 1 0 0 9 1 9 0 9 1 0 9 9 9 11 2 0 9 2 11 2 11 2 11 7 11 2
27 9 1 9 7 1 0 7 0 9 13 9 2 1 15 13 0 9 2 16 4 0 11 1 0 9 13 2
9 11 13 2 16 13 3 1 9 2
22 0 9 11 1 9 4 1 9 13 3 13 9 9 11 2 3 13 0 9 9 9 2
27 3 12 1 15 2 11 2 11 7 11 2 4 15 1 15 1 11 13 0 13 2 16 3 13 10 9 2
16 0 9 9 11 13 2 16 4 4 11 13 1 15 9 11 2
25 0 9 9 11 11 13 0 11 1 0 7 0 9 15 2 3 0 9 13 3 3 7 3 3 2
5 1 9 1 0 11
20 16 0 11 13 9 1 9 0 9 2 1 9 1 0 9 15 13 0 9 2
6 15 13 0 7 0 2
8 9 1 0 11 15 13 0 2
19 11 7 11 15 13 13 9 2 15 3 13 11 1 0 0 7 0 9 2
24 9 0 9 0 3 15 0 9 1 9 0 11 1 11 7 0 9 0 11 13 9 1 11 2
11 0 9 1 0 9 4 13 9 0 9 2
37 13 15 7 11 2 0 7 0 1 12 0 9 2 15 13 1 0 9 1 0 9 1 9 12 2 9 2 3 13 1 10 0 9 1 0 9 2
8 3 13 3 1 9 1 0 2
21 1 9 0 9 15 13 2 16 11 4 13 0 9 1 9 2 9 7 0 9 2
9 0 9 9 9 13 0 0 9 2
19 9 11 11 15 7 13 13 0 0 9 0 0 9 7 10 9 9 9 2
37 9 13 1 9 0 7 0 9 2 1 15 13 13 0 9 0 9 2 13 1 9 0 9 7 13 0 7 0 9 7 0 0 9 2 11 2 2
14 9 10 9 13 11 16 0 9 13 9 7 10 9 2
49 10 9 13 1 11 1 0 9 1 9 0 9 2 13 9 1 0 9 0 1 0 9 7 13 2 16 9 13 0 13 0 9 1 0 12 9 0 0 9 1 10 9 1 12 9 1 9 0 2
5 9 9 0 9 13
17 9 0 11 13 0 9 1 10 0 9 1 3 16 12 9 9 2
30 1 0 10 12 9 0 9 2 10 9 15 3 13 1 12 2 3 3 13 3 0 9 1 9 0 7 3 7 0 2
24 3 7 13 9 2 7 1 15 7 3 0 9 1 15 2 16 13 0 9 3 3 3 0 2
25 0 9 3 1 10 3 1 9 3 0 9 9 13 3 0 9 2 15 4 3 13 13 9 9 2
9 7 1 15 13 3 0 9 9 2
15 9 2 15 15 9 13 2 4 1 0 9 13 3 0 2
26 10 0 9 2 16 1 15 13 2 7 13 0 2 16 9 9 2 15 9 1 9 13 2 3 13 2
10 3 3 15 13 13 1 9 0 9 2
30 1 10 0 9 4 15 13 13 3 1 0 9 2 7 3 13 4 13 3 1 9 12 2 3 4 11 13 0 9 2
29 1 9 7 13 10 9 0 3 1 9 2 16 1 9 0 9 13 0 0 9 2 0 7 0 9 2 9 3 2
16 1 9 9 1 13 15 11 7 11 7 13 11 3 3 3 2
26 16 4 10 10 9 13 4 2 1 11 2 15 1 9 12 13 13 9 2 4 13 3 0 0 9 2
16 9 13 13 9 2 15 13 11 3 13 0 9 0 9 11 2
20 9 0 9 13 3 0 10 9 2 11 3 13 3 12 9 2 11 12 9 2
15 0 11 3 13 9 1 0 9 2 15 1 0 9 13 2
19 9 0 9 7 13 0 9 9 2 16 15 13 9 1 11 3 0 13 2
36 1 9 15 3 13 13 0 9 9 2 15 3 7 3 13 0 9 0 11 2 11 7 11 2 7 15 3 13 0 13 10 0 9 1 9 2
7 2 9 11 13 0 9 2
14 1 15 13 9 1 11 2 2 13 12 1 0 9 2
8 2 0 11 13 1 0 9 2
8 15 4 15 13 13 1 9 2
19 7 16 13 13 9 11 2 3 3 13 0 2 2 13 0 9 11 11 2
44 1 10 9 3 1 9 0 9 13 4 13 9 3 0 2 15 3 13 0 9 11 7 11 1 0 0 9 2 1 15 9 13 3 3 7 1 15 13 0 9 7 0 9 2
14 3 7 9 1 9 9 0 11 3 7 3 13 4 2
21 9 15 7 3 13 13 0 9 2 15 4 9 1 9 13 1 9 1 9 9 2
26 9 0 11 4 13 13 0 9 9 7 13 1 0 9 1 3 0 9 2 3 0 0 2 14 2 2
5 0 9 13 1 9
2 11 2
2 11 2
22 11 11 2 12 0 9 0 0 9 11 11 2 13 1 9 1 0 1 0 9 11 2
19 1 9 15 13 3 3 2 16 15 13 1 0 9 7 13 9 1 9 2
11 1 9 13 12 9 3 1 9 7 9 2
7 11 7 11 15 13 1 9
2 11 2
2 11 2
20 0 9 0 0 9 11 11 13 11 7 11 2 16 4 13 9 10 0 9 2
22 1 9 0 9 11 3 13 1 9 0 9 0 9 2 15 4 13 13 1 9 9 2
14 0 9 4 13 4 13 3 2 16 4 9 13 0 2
18 1 0 9 0 9 0 0 9 13 9 9 2 13 15 1 9 2 2
5 11 13 1 9 9
2 11 2
2 11 2
29 11 3 1 12 2 0 9 0 9 1 0 9 2 11 2 13 1 9 0 9 2 15 4 1 9 9 11 13 2
24 3 13 9 0 9 1 9 11 11 11 2 11 3 13 2 15 10 9 2 0 1 9 11 2
16 1 0 9 13 1 11 1 9 9 3 12 9 0 12 9 2
5 11 11 13 1 11
3 11 9 13
3 0 11 2
16 0 9 0 9 13 7 0 9 0 9 12 2 9 11 11 2
14 9 12 9 0 9 13 11 7 0 9 9 11 11 2
29 15 13 1 9 9 11 3 1 9 1 9 3 13 9 9 2 15 4 13 0 9 0 9 1 9 0 9 11 2
10 13 15 2 16 9 1 9 13 3 2
21 1 9 15 13 2 16 0 9 11 7 0 9 13 4 13 1 0 9 0 11 2
17 11 13 7 1 9 1 11 13 7 9 15 13 13 9 11 11 2
18 0 9 9 15 3 1 10 9 13 1 11 3 1 0 9 1 11 2
28 13 2 16 11 13 9 3 0 2 7 0 9 9 2 15 15 1 10 9 9 1 9 0 9 13 1 9 2
26 1 9 11 0 1 9 1 0 9 15 13 2 16 9 13 13 13 0 15 9 1 0 7 0 11 2
29 0 9 15 3 13 1 3 0 0 9 11 2 7 3 1 9 11 1 9 2 15 4 13 13 9 3 1 11 2
4 11 13 0 9
4 11 13 1 9
2 11 2
22 11 3 13 2 16 13 9 9 9 11 9 2 12 1 9 15 9 0 9 1 11 2
11 13 15 9 9 11 1 0 9 11 11 2
27 13 2 16 0 9 13 10 0 9 7 3 13 1 0 9 0 1 9 0 9 15 9 9 1 9 11 2
27 0 0 9 1 9 1 11 3 1 11 13 2 16 13 13 0 9 2 3 13 0 9 1 9 0 9 2
38 2 13 1 15 0 9 2 7 0 13 13 7 13 2 3 1 15 11 13 7 1 15 15 13 2 2 13 9 0 9 11 11 1 9 9 1 11 2
29 9 0 9 11 11 13 2 16 11 13 13 13 1 10 0 0 9 2 3 7 13 9 1 10 9 1 0 9 2
4 11 13 9 11
5 9 13 1 0 9
2 11 2
27 9 13 0 9 0 9 1 11 7 0 9 1 0 0 9 11 13 9 0 9 1 0 9 11 1 11 2
15 9 12 9 15 13 1 9 0 2 0 7 0 9 11 2
15 13 3 9 1 9 9 0 9 0 9 9 1 12 9 2
15 1 0 12 9 4 13 1 11 13 12 1 9 0 9 2
14 0 9 13 3 9 1 11 7 3 13 13 0 9 2
21 0 9 13 9 15 0 9 1 11 7 13 0 9 13 0 9 7 9 0 9 2
3 9 13 2
28 1 0 9 0 9 15 13 9 9 1 11 7 11 1 12 9 9 2 16 1 0 9 12 13 12 9 9 2
4 9 1 11 2
22 11 13 13 13 9 1 9 9 1 0 9 2 15 4 13 0 0 9 1 0 9 2
9 11 13 13 9 1 9 13 3 9
2 11 2
49 0 9 7 9 0 0 9 0 9 11 11 13 10 9 1 0 9 0 9 2 1 15 13 9 3 12 9 7 0 9 1 9 3 16 12 9 9 2 7 13 13 13 9 0 0 9 10 9 2
13 3 13 3 0 9 1 0 9 0 9 0 9 2
15 11 3 3 13 9 2 1 15 15 13 10 0 0 9 2
27 1 9 4 13 3 12 9 2 1 15 11 11 2 0 9 9 11 2 13 1 0 9 1 0 9 9 2
7 1 9 13 11 10 9 2
5 1 9 3 11 13
5 7 0 9 13 0
2 11 2
32 9 11 15 1 12 9 13 13 9 11 12 11 2 15 15 3 1 9 13 1 0 9 1 9 12 9 2 14 12 9 2 2
19 9 0 9 13 0 9 15 2 16 7 9 9 11 7 9 11 13 0 2
9 13 2 16 10 9 13 3 0 2
15 2 13 2 16 4 15 3 13 3 16 0 13 9 2 2
8 9 0 11 11 13 1 9 9
11 2 13 9 11 2 9 11 11 11 2 2
12 2 13 15 2 9 2 13 11 11 11 2 2
10 2 3 1 9 15 13 2 3 13 2
11 7 3 9 13 1 15 2 2 13 9 2
7 2 13 4 14 12 9 2
14 13 4 13 2 9 2 16 9 13 1 0 11 2 2
25 3 13 0 9 0 11 9 12 0 9 0 9 1 9 12 2 1 9 12 2 9 1 9 11 2
53 1 12 9 9 11 2 0 9 2 0 3 1 9 16 1 9 0 9 9 1 9 2 11 2 2 1 9 0 9 2 9 1 0 9 2 0 11 11 11 2 9 0 9 2 3 0 0 9 1 9 0 11 2
42 1 10 9 1 9 13 0 9 0 9 9 11 11 2 11 2 16 15 13 13 14 1 9 7 0 9 1 11 11 1 11 7 16 15 11 13 13 0 0 9 9 2
21 1 12 9 9 9 15 13 1 12 12 9 2 7 14 2 10 9 3 13 0 2
7 9 11 13 1 0 9 2
11 13 1 15 7 9 9 2 7 9 9 2
6 9 13 0 9 9 2
46 3 1 11 13 1 9 9 3 11 11 2 10 9 7 9 2 9 3 16 2 9 11 2 2 11 11 2 2 9 11 2 2 0 0 9 2 15 15 14 1 9 13 1 9 9 2
12 7 3 9 9 7 10 9 2 9 11 11 2
19 1 10 9 2 15 15 13 1 9 11 9 2 15 9 13 11 1 9 2
15 13 15 0 9 2 3 0 9 7 9 9 11 1 9 2
27 15 13 2 16 4 15 11 13 2 16 11 2 2 9 2 2 9 2 13 0 14 12 9 9 2 11 2
27 15 15 13 3 1 0 9 1 2 9 2 2 1 9 12 7 9 12 2 3 7 1 15 13 14 9 2
20 7 16 9 13 9 1 9 2 15 1 9 13 11 2 13 15 9 3 0 2
21 0 9 11 2 9 2 9 2 9 2 12 1 0 9 9 2 13 3 1 9 2
21 10 2 0 9 2 13 12 2 9 12 2 3 15 1 11 2 9 11 2 13 2
7 1 9 0 9 7 9 2
28 3 15 15 13 13 9 7 9 1 0 9 2 9 13 9 2 1 0 9 9 2 7 2 0 0 9 2 2
26 1 10 0 9 3 13 3 0 9 2 15 15 13 7 15 2 16 1 10 9 13 1 0 9 11 2
31 1 9 12 15 13 1 0 9 1 11 11 0 11 2 1 15 15 3 13 2 9 9 2 1 12 1 0 9 9 9 2
27 1 9 3 13 11 3 1 11 2 3 3 13 3 2 2 7 11 15 13 9 1 2 0 0 9 2 2
18 7 3 13 9 0 9 9 1 11 7 3 15 13 9 1 9 9 2
11 15 3 13 0 9 1 9 1 9 12 2
23 10 9 9 9 9 13 16 2 0 9 9 2 7 13 16 9 9 2 15 13 9 9 2
13 10 9 13 9 0 9 2 15 13 13 9 9 2
9 13 3 0 2 16 9 13 0 2
14 9 11 11 7 3 13 9 10 0 9 7 0 9 2
6 16 15 9 13 3 3
6 7 9 13 13 1 9
3 11 0 2
22 10 9 3 13 0 9 2 15 13 1 9 1 11 1 9 0 9 1 9 1 9 2
28 1 9 3 3 13 9 13 1 9 2 16 4 1 15 13 10 9 2 3 16 4 15 13 9 1 0 9 2
13 3 15 12 9 13 1 9 7 13 9 12 9 2
5 9 13 9 1 9
2 11 2
2 11 2
24 1 11 15 3 13 0 9 1 0 0 9 2 15 4 13 9 1 0 7 0 9 1 9 2
16 9 9 11 13 9 2 16 4 15 13 1 0 9 1 9 2
16 1 0 9 11 3 13 0 9 7 13 2 16 0 9 13 2
12 9 1 9 0 0 9 13 10 9 0 9 2
3 13 1 9
1 9
13 1 0 9 1 9 7 9 13 10 0 0 9 2
20 11 11 3 1 11 2 15 15 13 1 11 2 15 1 9 13 1 11 11 2
11 9 11 0 2 2 3 13 1 9 9 2
7 13 15 1 10 9 13 2
9 3 13 2 16 15 13 1 11 2
7 3 2 16 13 0 9 2
25 0 13 9 11 2 15 13 9 1 9 2 0 2 15 13 0 0 9 2 7 9 13 0 9 2
6 14 3 13 13 11 2
12 16 15 13 9 11 2 13 4 1 0 9 2
14 9 9 9 2 3 1 15 13 2 13 3 1 15 2
15 16 15 9 1 15 13 2 13 3 1 0 9 9 2 2
22 11 11 11 1 9 1 11 1 9 12 2 9 13 3 1 9 1 11 1 11 11 2
20 9 11 11 2 2 13 1 15 12 0 9 2 0 1 11 7 0 1 11 2
27 1 9 3 13 0 9 1 11 2 3 4 13 12 2 12 2 7 1 0 12 9 4 15 13 7 13 2
10 13 13 3 2 7 16 13 11 9 2
8 0 13 13 1 9 7 9 2
14 9 3 13 3 0 15 2 15 15 13 1 11 2 2
20 11 1 9 1 12 9 13 11 11 2 15 1 0 9 13 11 11 12 9 2
12 9 9 11 11 2 2 1 10 9 13 9 2
15 13 7 2 15 15 13 2 13 15 13 0 9 1 9 2
7 10 9 15 3 13 9 2
8 0 9 13 11 7 0 11 2
18 3 0 1 0 9 1 11 2 15 4 13 12 2 12 2 13 11 2
6 9 10 9 13 0 2
12 3 3 7 11 2 15 13 0 9 1 9 2
17 10 9 7 13 2 13 3 10 0 9 7 13 9 1 9 2 2
2 0 9
8 9 13 9 1 9 7 9 2
13 11 11 3 13 1 0 11 2 1 9 13 11 2
14 9 11 11 2 2 7 12 1 9 13 1 10 9 2
26 1 0 9 3 1 11 2 15 7 13 3 0 9 2 15 13 2 16 10 9 13 7 1 9 11 2
17 13 3 13 3 9 12 9 1 0 9 3 1 0 0 9 2 2
18 11 1 0 9 3 1 12 9 13 11 2 1 9 15 13 1 11 2
19 9 11 11 2 2 1 9 9 4 13 2 16 13 9 0 9 16 3 2
19 13 15 2 16 13 3 13 0 2 16 1 9 9 0 9 13 14 11 2
17 13 15 1 9 9 7 0 15 3 13 9 13 2 15 13 0 2
7 1 10 15 13 13 9 2
18 16 13 1 11 2 3 15 13 15 13 1 0 9 1 9 9 14 2
11 0 4 3 13 2 16 1 15 13 2 2
4 0 13 1 9
12 11 11 15 13 1 9 7 13 15 9 0 9
17 7 14 1 9 9 15 1 10 9 1 9 11 3 13 11 11 2
8 1 11 15 13 16 9 9 2
15 2 1 9 4 13 3 9 2 13 15 7 7 7 3 2
14 3 3 13 13 1 9 3 2 2 13 10 0 9 2
8 2 3 13 0 9 2 13 2
21 0 9 1 9 3 1 11 13 1 15 2 16 11 13 3 1 9 9 1 9 2
18 2 14 4 13 0 2 10 0 9 1 9 7 1 15 1 11 13 2
17 7 13 2 16 15 1 10 9 1 11 13 3 3 16 9 3 2
10 13 15 2 16 1 12 2 9 13 2
22 1 9 9 4 15 13 3 1 9 2 0 9 13 1 0 9 2 15 15 3 13 2
9 13 15 15 1 11 3 2 2 2
10 3 15 2 13 4 3 1 0 9 2
22 2 1 10 9 15 15 13 2 7 0 4 9 7 12 13 7 13 15 1 9 2 2
12 2 13 4 2 16 15 15 13 2 15 3 2
19 2 9 1 11 13 1 10 0 9 1 9 2 7 3 15 13 15 0 2
9 13 10 9 2 15 15 15 13 2
7 3 15 7 13 15 2 2
18 2 15 15 13 1 15 2 16 3 3 0 9 13 1 10 9 3 2
29 11 11 7 11 13 1 11 2 0 9 13 9 2 15 13 1 11 13 9 1 3 16 9 7 3 13 1 9 2
8 2 13 9 2 16 3 13 2
24 7 1 0 9 4 10 0 9 13 13 0 0 9 2 15 4 15 1 9 0 9 13 3 2
16 12 4 9 3 13 2 7 3 13 3 0 1 9 2 2 2
8 13 4 15 1 0 0 9 2
21 15 4 3 1 10 9 13 13 0 0 9 9 2 15 3 3 1 9 13 9 2
17 2 9 15 13 2 16 13 9 2 7 3 3 13 0 0 9 2
9 15 3 13 3 0 3 0 9 2
5 15 7 9 13 2
12 0 9 4 1 15 13 13 12 7 12 9 2
13 15 2 16 13 9 9 2 4 15 13 3 13 2
14 13 7 2 16 3 1 11 1 15 3 13 9 9 2
17 3 15 7 13 13 2 16 0 9 13 1 0 9 3 13 2 2
12 2 1 10 9 11 4 13 3 1 9 13 2
13 2 15 13 15 12 2 0 13 13 15 3 2 2
10 9 2 0 12 2 11 12 2 12 12
23 1 10 9 13 7 1 9 2 1 15 13 9 9 2 7 1 15 2 15 13 0 9 2
19 1 9 1 0 9 1 11 1 9 1 9 1 9 13 11 9 1 11 2
17 2 13 15 0 2 3 14 13 0 9 7 1 15 15 13 9 2
10 13 4 15 7 1 9 12 1 9 2
25 2 13 15 3 3 2 3 4 3 15 2 11 2 10 9 1 0 7 3 13 13 1 9 2 2
8 15 13 9 2 3 15 13 2
16 1 9 9 12 4 13 1 9 7 10 9 1 9 1 11 2
13 13 4 1 9 1 11 2 14 12 9 1 11 2
17 13 4 15 2 16 15 13 7 13 0 2 0 9 1 9 11 2
18 13 4 7 13 2 13 1 9 2 13 7 1 9 9 13 1 11 2
18 1 9 4 15 13 1 9 9 1 11 2 15 13 0 9 16 15 2
17 1 9 2 3 4 4 13 2 13 1 15 1 0 9 0 12 2
7 12 1 15 13 1 9 2
19 3 2 16 4 15 13 3 2 16 4 15 13 14 3 2 1 0 11 2
6 15 13 1 9 3 2
24 15 4 4 1 9 13 1 9 1 9 9 2 9 0 9 2 1 10 9 4 13 1 9 2
20 1 0 9 11 4 3 13 13 9 2 13 4 0 2 13 9 1 12 9 2
14 13 4 15 13 9 2 16 4 13 13 1 9 9 2
16 13 1 10 9 0 2 3 3 2 9 15 13 1 9 13 2
13 3 15 7 3 13 0 9 2 13 0 1 9 2
8 0 13 2 0 13 1 9 2
30 7 13 2 7 14 1 9 10 9 2 15 15 3 3 13 1 2 0 7 0 2 9 0 9 2 2 13 9 9 2
24 1 9 2 15 13 1 9 1 9 9 9 2 13 11 11 1 11 2 9 0 9 9 9 2
45 2 13 15 3 12 9 2 16 9 9 9 13 9 0 9 7 11 11 2 16 4 13 0 9 2 1 0 9 13 9 0 9 7 13 0 9 1 9 9 7 9 9 0 9 2
20 1 10 9 15 13 3 15 2 16 11 13 0 9 2 7 1 10 0 9 2
16 9 7 9 9 15 3 13 2 7 15 15 13 1 0 9 2
45 7 3 13 9 9 1 0 9 1 9 0 9 2 1 15 1 0 13 9 9 2 9 7 9 0 9 1 12 2 12 2 12 2 9 9 7 9 9 0 1 9 7 0 9 2
17 0 0 9 13 1 9 3 3 0 0 9 2 15 13 0 9 2
7 3 3 13 9 7 9 2
15 9 3 13 7 9 9 2 9 2 7 3 1 9 9 2
19 1 11 3 3 13 0 9 7 9 2 13 9 2 9 13 1 9 9 2
18 1 0 9 4 9 1 10 9 13 1 0 9 2 7 9 13 0 2
19 16 15 9 9 7 9 1 9 13 0 2 13 7 15 9 1 9 9 2
7 9 9 13 1 9 9 2
29 9 13 13 1 0 0 9 9 9 1 11 12 2 1 9 0 12 2 0 2 9 2 12 2 2 13 9 11 2
13 1 9 1 11 9 2 9 9 9 11 11 11 2
16 0 11 2 15 13 9 0 9 9 2 4 3 13 1 9 2
12 1 0 9 15 7 0 9 1 10 9 13 2
19 2 1 11 13 3 0 9 2 16 3 13 1 9 7 9 9 1 9 2
9 3 7 1 15 13 9 10 9 2
15 15 13 1 0 9 2 15 13 1 9 0 0 1 15 2
15 1 0 9 4 0 13 2 7 13 15 13 3 0 9 2
21 3 7 4 13 0 9 9 1 12 9 2 1 15 4 15 0 13 13 1 9 2
24 13 3 3 1 9 11 1 11 2 11 1 12 9 7 3 15 0 9 1 9 13 13 2 2
4 9 13 11 11
2 1 9
37 0 0 9 11 11 11 11 2 15 13 1 10 9 7 9 1 9 11 2 11 7 3 13 1 9 9 11 2 11 2 13 10 9 11 1 9 2
30 9 11 9 2 15 13 1 11 1 11 2 3 1 9 13 1 9 11 1 11 9 2 3 13 13 9 1 0 9 2
15 2 3 3 7 3 13 2 2 13 15 9 11 11 11 2
3 11 1 9
5 11 2 11 2 2
45 9 12 0 9 2 2 2 2 7 9 13 2 2 2 3 2 2 2 2 2 2 9 1 9 1 9 2 7 2 2 2 2 7 3 13 13 0 9 2 13 3 0 9 11 2
29 9 2 15 13 0 9 11 11 2 13 1 9 9 9 0 9 0 9 1 9 0 9 7 9 1 9 10 9 2
16 13 1 9 1 9 0 9 11 2 10 0 9 7 9 9 2
3 9 1 9
5 9 1 0 9 2
13 9 0 12 9 13 1 12 0 9 1 0 9 2
11 13 15 3 7 3 16 0 9 9 11 2
11 1 11 9 1 0 9 13 0 0 9 2
28 3 1 12 9 13 0 9 9 2 9 13 3 1 12 9 7 0 9 4 13 13 1 9 1 12 2 9 2
4 9 13 1 9
5 11 2 11 2 2
25 0 9 1 11 3 13 0 9 1 11 11 2 2 0 2 16 1 9 12 13 1 11 0 9 2
7 9 13 9 9 1 9 2
11 9 9 13 0 9 1 9 1 9 9 2
8 13 0 7 3 0 0 9 2
8 3 1 10 9 13 10 9 2
21 9 16 0 13 3 0 11 11 2 2 15 3 13 1 9 2 3 4 9 13 2
18 15 3 13 16 9 2 7 13 2 16 3 1 0 9 13 0 9 2
25 1 9 0 9 7 4 13 9 1 10 9 2 1 9 11 11 2 9 13 9 0 1 9 9 2
4 0 9 13 2
3 9 1 9
23 1 0 9 9 1 11 13 1 9 0 9 12 9 0 9 0 9 2 15 13 0 9 2
12 9 9 15 13 0 9 1 9 1 0 9 2
10 1 12 2 9 13 0 9 1 9 2
32 1 9 1 0 9 1 0 7 0 0 9 15 1 9 9 0 9 11 11 3 13 9 2 15 13 0 0 9 13 1 11 2
15 1 0 9 13 12 9 13 2 16 0 9 13 1 15 13
2 9 9
18 0 9 1 9 0 0 9 4 1 12 2 9 13 1 0 9 11 2
25 13 3 1 11 7 11 1 11 1 0 9 1 9 2 15 4 13 0 9 9 0 1 0 9 2
8 2 13 0 0 9 1 9 2
27 9 1 9 2 9 2 9 7 0 0 9 4 13 9 2 9 2 9 7 0 0 9 3 1 12 9 2
10 15 15 13 13 9 1 10 0 9 2
7 3 13 13 0 0 9 2
18 4 3 13 0 9 10 9 2 2 13 9 0 9 0 9 11 11 2
12 9 13 0 9 2 9 15 13 13 3 3 2
3 13 1 11
16 9 11 11 11 13 1 9 12 2 9 9 11 1 9 3 2
22 1 9 0 9 9 11 9 1 11 13 9 1 11 2 1 15 15 3 13 1 11 2
7 3 13 1 12 9 9 2
21 1 0 9 13 9 1 9 13 1 12 9 0 2 15 13 1 12 9 10 9 2
20 2 9 1 9 7 1 10 9 12 2 12 13 3 0 2 2 13 11 11 2
11 9 11 15 3 1 11 3 13 16 3 2
28 1 10 9 13 7 14 0 2 2 3 4 1 9 13 10 9 2 7 3 7 7 15 13 1 15 0 9 2
19 0 9 13 3 0 16 3 0 2 16 15 9 13 2 3 3 13 2 2
4 9 1 9 13
7 1 0 0 9 3 13 9
5 0 9 13 9 2
14 9 1 15 1 0 9 1 11 1 11 13 3 0 2
10 13 15 2 16 15 15 1 9 13 2
16 9 9 9 2 12 4 13 0 9 2 9 0 0 9 13 2
26 3 13 9 12 1 10 0 1 9 2 7 15 3 1 0 9 2 15 15 1 0 9 13 3 13 2
29 2 15 15 4 13 0 9 2 13 2 2 13 15 9 0 9 7 3 9 9 9 11 11 11 1 11 11 11 2
11 2 1 9 0 9 3 13 0 9 13 2
17 0 9 2 1 15 15 15 13 3 12 9 2 13 3 13 13 2
18 14 9 9 4 13 12 9 7 3 15 13 14 9 1 15 12 9 2
12 0 9 1 9 1 9 9 13 1 9 12 2
14 13 15 9 9 9 2 1 10 9 4 13 3 15 2
13 3 0 9 15 1 0 9 3 13 12 9 2 2
15 9 13 0 9 0 13 1 9 9 7 1 9 1 9 2
15 12 9 1 9 13 0 9 12 9 2 0 12 9 2 2
17 12 9 15 3 3 13 11 2 7 3 13 0 12 9 3 13 2
23 3 15 13 0 9 2 15 7 3 13 3 1 9 0 9 2 15 15 13 1 12 9 2
10 1 15 3 13 2 2 13 9 11 2
32 15 13 3 1 11 11 2 1 15 9 1 0 9 1 9 12 4 9 13 2 9 9 1 9 0 9 0 1 9 1 9 2
17 1 9 11 11 2 11 9 1 9 13 12 9 9 1 0 9 2
7 3 15 13 1 12 9 2
19 1 0 9 7 9 11 13 0 13 9 2 7 3 9 1 12 9 13 2
16 10 9 1 9 1 0 9 9 13 9 0 9 13 12 9 2
19 0 9 3 13 1 9 9 2 15 4 13 13 1 0 9 1 0 9 2
12 0 9 4 1 0 9 13 3 3 12 9 2
6 0 9 2 0 9 2
7 0 9 0 9 1 0 9
22 2 13 0 9 16 9 9 1 0 9 2 3 3 4 1 9 9 13 13 0 9 2
19 7 13 15 1 9 1 9 9 9 1 9 0 9 1 0 7 0 9 2
35 9 13 2 16 1 0 9 3 4 9 13 1 9 2 7 1 9 9 2 2 13 15 15 1 9 9 0 9 1 11 2 11 11 11 2
21 0 9 3 3 13 0 12 12 7 1 9 1 9 0 15 13 13 7 1 9 2
52 9 0 9 0 0 9 0 9 2 0 9 12 5 2 0 12 5 7 0 12 5 1 9 1 9 0 2 13 14 0 9 7 9 0 9 2 7 7 9 11 2 15 15 1 15 1 2 0 2 9 13 2
25 3 3 13 9 0 9 0 0 9 1 0 12 1 12 9 2 16 15 3 13 1 9 0 9 2
13 13 4 15 0 9 0 9 9 9 2 11 11 2
16 2 9 2 16 9 0 9 15 3 3 13 2 13 3 0 2
36 9 9 3 13 0 9 7 13 9 2 16 4 0 9 13 13 1 10 9 2 7 1 9 9 9 1 0 0 9 7 9 3 13 9 0 2
22 9 10 9 3 13 2 7 16 15 13 13 2 13 2 16 13 0 9 0 9 13 2
20 3 15 13 9 9 2 16 15 10 9 2 3 0 9 0 9 2 13 13 2
38 13 7 1 9 13 15 7 3 12 9 0 9 2 16 15 1 0 9 0 9 7 0 9 0 9 1 9 9 13 3 9 9 1 0 9 9 2 2
13 13 0 9 7 3 9 0 2 16 13 0 9 2
34 2 15 13 0 9 2 3 15 15 0 9 9 1 9 0 9 13 3 0 2 16 9 1 0 7 0 9 15 1 10 9 3 13 2
34 1 9 9 15 3 3 13 12 9 2 7 16 4 13 0 9 3 0 2 7 7 9 13 9 3 3 1 9 7 9 1 9 9 2
32 0 13 3 1 9 9 0 2 7 7 1 9 13 15 3 3 2 15 0 9 9 1 9 2 15 0 9 1 15 9 2 2
49 13 15 2 16 9 2 15 15 13 0 0 0 9 2 4 13 1 9 1 9 13 3 2 16 3 13 1 9 0 7 0 2 1 9 7 1 0 9 2 9 3 13 10 9 1 9 15 9 2
24 3 3 3 13 1 9 12 7 12 9 1 15 2 16 4 15 9 9 13 1 9 0 9 2
34 2 9 13 0 9 2 16 3 10 9 13 1 9 1 12 9 2 7 13 12 0 9 2 16 9 9 13 1 12 10 9 3 0 2
11 9 9 9 1 9 3 7 13 3 3 2
23 3 13 9 2 16 1 0 9 13 9 0 9 7 1 0 9 4 7 3 13 0 9 2
35 16 15 7 3 13 12 9 2 13 10 9 2 9 9 1 9 13 0 7 9 0 0 9 2 3 13 15 9 0 2 13 0 9 3 2
25 13 7 1 0 13 9 15 2 16 13 15 3 3 2 7 13 3 7 15 9 9 1 9 2 2
11 3 13 9 9 1 9 0 7 0 9 2
23 2 13 4 14 1 0 9 2 1 0 9 15 10 9 13 3 14 1 9 0 9 9 2
26 1 0 9 15 3 3 13 13 9 2 15 4 9 9 9 13 7 13 3 0 9 1 9 1 15 2
33 1 1 15 2 16 0 9 13 0 3 13 7 3 3 13 10 0 9 2 13 9 9 14 1 0 0 9 2 3 1 9 12 2
11 7 16 15 4 9 0 9 14 13 2 2
17 1 9 9 0 9 13 13 2 9 15 15 13 13 1 0 9 2
12 9 0 9 9 1 9 3 13 3 3 9 2
26 0 9 2 15 0 9 13 9 2 13 9 2 16 9 0 13 1 9 12 9 0 9 1 9 0 2
26 7 0 9 14 13 9 2 16 3 3 13 9 1 0 9 7 0 0 9 2 15 4 13 0 9 2
2 11 11
4 9 2 11 2
2 11 11
1 9
5 0 9 0 16 9
14 10 9 15 1 9 0 9 13 1 9 1 0 9 2
15 3 9 9 2 9 9 7 0 0 9 13 13 0 9 2
11 1 0 9 13 3 0 0 9 0 9 2
8 1 9 9 1 15 13 9 2
9 13 1 0 9 0 9 1 9 2
12 13 15 3 9 2 15 13 3 1 0 9 2
15 1 12 2 9 13 1 9 0 9 1 11 7 0 9 2
14 13 0 9 0 9 1 9 10 0 9 1 9 9 2
11 3 3 0 9 9 7 9 13 0 9 2
15 13 15 7 2 16 1 11 3 13 2 3 0 9 13 2
12 11 3 4 3 7 3 3 13 1 9 9 2
8 10 9 13 1 9 1 9 2
31 9 3 9 13 2 16 0 9 13 9 13 2 3 7 13 2 16 13 9 13 2 3 13 13 2 15 7 1 10 9 2
9 1 10 9 9 4 13 1 9 2
6 13 4 9 0 9 2
12 11 2 11 7 11 7 1 9 9 9 13 2
11 13 1 9 2 16 10 9 13 10 9 2
10 13 15 1 9 11 9 13 0 9 2
21 3 15 13 2 16 7 10 9 2 15 3 9 13 2 15 1 15 4 13 13 2
18 0 9 9 1 9 13 2 16 9 15 13 3 13 9 1 9 9 2
19 13 4 13 0 10 9 1 9 9 3 13 7 13 2 3 9 0 9 2
22 1 0 9 7 13 9 2 16 4 9 1 0 9 13 1 0 9 14 0 0 9 2
11 3 2 1 0 15 3 13 3 0 9 2
13 7 1 0 9 10 0 9 13 1 3 0 9 2
14 1 9 0 9 10 9 1 9 11 13 7 12 9 2
17 7 9 9 3 13 13 2 16 9 9 13 3 1 9 0 9 2
2 11 11
3 0 9 13
19 12 1 9 0 9 0 0 9 1 9 9 13 10 3 0 9 1 15 2
17 1 0 0 9 9 0 9 13 7 9 9 15 13 1 0 9 2
15 15 2 13 2 14 13 9 9 2 4 13 13 0 9 2
8 9 13 12 9 2 9 0 2
29 11 13 1 9 9 1 10 9 2 15 13 9 12 1 0 9 3 0 9 1 11 1 0 9 1 9 0 9 2
7 9 3 4 13 12 9 2
18 3 13 9 1 9 7 9 9 2 15 13 0 9 0 9 11 11 2
19 15 13 1 15 1 0 9 13 9 7 0 7 0 9 0 11 7 9 2
17 9 0 9 13 13 12 9 12 0 9 7 9 0 9 1 9 2
5 9 7 9 13 2
13 0 9 13 3 0 9 1 9 0 9 1 9 2
20 3 9 1 9 9 0 9 4 13 0 9 2 15 3 13 7 0 0 9 2
24 0 9 0 9 1 9 0 9 15 1 0 7 0 0 9 13 1 2 0 2 9 0 9 2
13 15 13 2 16 9 13 1 10 9 7 0 9 2
8 0 9 15 7 13 0 9 2
14 13 0 13 9 0 9 16 9 7 9 0 0 9 2
7 10 9 15 13 2 13 2
17 1 0 9 3 13 7 0 9 2 15 9 9 13 7 13 9 2
11 7 0 9 0 0 9 3 9 9 13 2
19 0 9 4 13 14 3 2 16 9 13 9 9 1 9 7 9 0 9 2
23 15 13 3 7 0 0 9 7 13 15 2 3 13 13 9 15 2 15 13 13 15 0 2
19 3 2 16 13 9 13 9 9 1 0 9 2 15 4 13 3 0 9 2
7 7 3 12 9 13 0 2
15 9 15 2 3 16 1 0 0 9 2 13 1 0 9 2
9 7 15 13 1 0 9 10 9 2
2 11 11
6 9 2 1 15 4 13
22 1 0 11 3 13 0 9 9 2 0 9 7 0 9 1 0 9 2 9 7 9 2
26 1 0 9 9 1 10 9 13 12 9 1 12 9 2 7 3 15 11 13 1 0 0 9 1 11 2
22 4 13 1 9 2 13 7 4 1 12 0 9 9 1 9 7 3 12 9 1 11 2
32 1 9 13 7 9 0 9 11 11 2 9 0 9 11 1 11 2 9 11 2 11 2 11 11 2 0 11 2 11 7 11 2
17 10 9 15 13 13 14 1 0 9 2 13 3 7 0 0 9 2
8 13 0 13 2 3 15 13 2
19 11 11 2 9 0 9 11 1 12 9 2 13 9 9 2 9 7 9 2
11 2 1 0 11 4 13 0 9 1 11 2
13 1 0 9 15 15 13 0 11 2 16 13 0 2
10 1 11 3 3 1 10 9 13 2 2
16 1 9 1 9 0 7 9 9 0 9 15 13 9 11 11 2
24 1 0 9 7 9 15 3 9 2 16 13 3 2 13 13 0 9 2 9 9 7 0 9 2
23 1 9 2 10 9 15 1 9 1 12 9 13 2 13 0 9 11 11 11 2 16 12 2
12 15 7 13 10 9 2 13 14 13 7 12 2
22 2 1 9 13 12 9 10 9 0 9 11 7 9 2 2 13 15 13 9 11 11 2
17 1 9 0 11 13 9 1 9 9 2 9 7 9 9 9 11 2
10 9 13 3 14 3 0 0 9 11 2
32 0 9 13 1 9 0 9 11 11 1 12 9 11 2 15 15 13 1 9 7 9 1 11 2 15 15 13 1 9 7 9 2
18 11 2 9 2 1 9 2 0 2 2 13 1 9 10 0 0 9 2
26 13 12 9 3 11 11 2 11 13 2 7 9 15 13 13 2 16 3 13 13 9 2 2 2 2 2
22 9 9 11 11 2 2 13 15 3 11 2 15 13 9 1 9 2 11 3 1 11 2
11 11 15 13 9 7 13 1 15 10 9 2
19 13 2 16 15 15 13 13 10 9 1 11 2 10 9 13 1 0 2 2
4 0 9 1 9
36 16 0 9 13 9 1 9 9 1 11 0 2 3 2 2 9 1 11 7 11 13 3 0 9 1 0 0 9 2 15 13 13 9 0 9 2
40 7 13 9 9 9 12 0 7 0 9 1 12 2 0 0 9 1 11 2 15 3 13 2 3 12 0 9 2 10 9 1 0 9 13 1 9 0 9 9 2
11 13 15 15 11 11 1 0 9 7 9 2
24 9 1 9 1 11 13 14 10 0 9 1 3 0 9 2 7 7 9 9 2 0 0 9 2
16 1 0 9 15 13 9 1 11 1 0 9 3 13 0 9 2
3 9 1 11
5 11 2 11 2 2
32 12 9 0 9 11 13 9 13 0 0 9 0 9 7 13 15 2 3 1 0 0 0 9 11 11 7 11 9 2 0 9 2
10 1 9 1 9 9 11 1 11 13 2
40 9 9 9 1 9 0 2 9 2 11 2 9 2 11 11 11 15 13 2 16 11 4 1 11 13 13 9 1 9 2 9 2 0 9 7 0 9 0 9 2
20 9 9 9 11 13 14 9 1 0 0 9 2 1 15 15 0 0 9 13 2
5 9 11 1 0 9
15 1 9 9 11 7 11 13 3 1 9 9 13 0 9 2
29 12 9 7 13 13 9 13 0 9 2 3 4 15 9 13 0 2 13 3 1 11 9 9 7 9 11 11 11 2
22 12 9 13 13 0 0 9 1 9 7 13 9 2 15 9 0 9 4 13 1 11 2
14 13 4 7 13 0 7 0 9 2 15 13 0 11 2
19 1 0 9 13 13 9 2 3 3 0 9 13 2 13 1 9 12 9 2
28 9 1 9 0 9 13 1 9 1 11 2 11 7 0 2 0 9 2 3 16 12 9 13 9 10 9 13 2
4 0 9 0 9
13 9 0 9 15 1 9 13 1 0 12 9 9 2
7 13 15 1 9 9 9 2
26 3 3 13 0 2 16 1 0 9 12 2 13 12 2 9 2 13 9 1 9 7 9 11 0 9 2
27 1 0 12 9 0 0 9 13 0 9 12 9 9 2 16 3 15 13 1 0 9 12 2 12 9 9 2
11 1 0 0 0 9 13 9 12 9 9 2
18 0 9 13 2 16 1 9 0 0 9 15 9 13 1 12 9 9 2
12 0 0 0 9 11 13 3 16 12 9 9 2
18 3 9 1 0 9 13 0 7 0 9 2 9 7 9 1 9 11 2
14 15 3 13 1 0 9 0 9 3 16 0 9 9 2
30 1 0 12 9 0 0 9 13 9 1 9 0 9 12 9 9 2 16 0 9 1 9 13 1 0 9 12 9 9 2
19 0 9 7 0 9 13 2 16 9 0 9 15 13 3 0 9 0 9 2
13 9 0 0 9 0 9 0 9 2 12 2 0 9
31 1 9 0 9 0 9 13 0 9 1 9 0 9 1 0 9 11 12 2 9 1 11 11 7 3 9 9 1 11 9 2
51 1 1 15 2 16 0 0 9 1 9 12 0 9 2 12 2 12 2 12 1 12 9 2 4 3 15 13 2 13 7 1 0 9 0 7 0 9 2 15 15 13 4 13 2 0 9 13 1 3 0 2
19 15 15 13 3 0 9 11 9 2 1 15 9 15 9 1 9 3 13 2
46 3 15 3 13 2 3 1 9 0 2 9 1 9 0 9 2 2 11 11 12 2 12 2 12 7 11 9 12 2 12 2 12 2 4 1 0 11 13 0 9 7 13 0 0 9 2
19 1 9 7 0 7 0 9 13 2 16 13 0 9 1 9 0 9 13 2
22 9 9 11 11 7 9 11 3 13 2 16 0 9 13 9 0 9 1 12 0 9 2
16 3 0 9 13 1 9 0 2 1 9 11 9 0 12 9 2
43 1 10 9 7 13 3 0 2 16 0 9 13 1 9 12 0 9 1 9 0 9 9 7 3 1 1 9 1 9 12 9 3 0 1 0 11 7 0 9 0 9 11 2
2 1 9
3 9 0 9
42 1 9 9 1 0 9 15 1 0 9 0 0 9 2 9 2 9 2 0 0 9 2 9 2 11 13 1 0 9 1 12 9 7 1 0 9 0 9 1 12 9 2
16 11 3 13 12 2 12 0 9 9 2 0 1 0 0 9 2
5 0 9 13 1 9
24 1 9 13 9 1 9 13 3 0 9 0 9 0 1 12 7 12 9 1 12 1 12 9 2
9 0 9 13 3 1 0 13 9 2
19 9 9 15 3 13 3 0 9 0 0 9 2 15 13 12 9 1 9 2
27 9 9 3 13 3 0 9 0 0 9 1 9 2 15 13 9 12 9 9 1 9 12 9 9 1 9 2
36 9 9 7 0 9 11 7 11 3 1 0 9 13 2 16 4 13 1 9 0 0 9 2 11 2 7 4 13 1 0 9 2 15 11 13 2
24 3 13 2 16 13 9 13 0 9 1 9 7 9 2 7 0 9 13 0 0 9 12 9 2
14 3 1 9 9 13 9 9 1 9 1 12 1 12 2
15 0 9 13 1 9 0 9 9 13 0 0 9 0 9 2
21 13 15 2 16 14 1 9 13 1 0 9 1 0 9 9 0 15 12 9 9 2
25 16 4 4 0 9 13 2 13 9 2 16 15 0 9 0 9 2 14 12 9 9 2 3 13 2
34 16 4 9 13 0 9 2 0 9 7 0 9 7 13 2 13 4 15 0 9 0 0 9 7 1 15 0 0 9 9 1 9 11 2
19 0 0 9 3 13 9 0 9 2 16 1 9 0 9 3 13 9 9 2
25 1 0 9 13 0 9 2 15 13 9 0 9 2 13 0 9 1 0 0 9 1 9 1 9 2
20 1 9 13 1 0 9 2 0 0 9 11 2 15 13 0 9 1 12 9 2
30 0 9 4 0 9 1 9 0 0 9 2 9 2 13 1 12 9 7 3 15 1 0 9 3 13 1 0 9 9 2
24 11 2 15 0 9 13 10 9 1 11 2 1 9 13 13 0 0 9 1 12 1 12 9 2
17 0 11 1 11 13 1 0 9 13 10 0 9 9 1 0 9 2
12 13 1 0 0 9 0 9 1 9 9 12 2
11 9 0 0 9 13 15 12 0 0 9 2
12 0 9 13 13 0 9 7 9 1 0 9 2
3 11 7 11
21 11 13 9 11 2 3 0 9 9 1 9 7 9 9 1 9 9 0 9 9 2
12 0 9 9 4 3 13 3 13 0 9 9 2
18 13 15 1 9 0 9 11 9 11 1 9 1 9 11 13 1 11 2
12 9 1 9 9 13 12 9 15 0 9 11 2
32 1 0 9 11 1 11 11 13 1 0 9 12 0 9 1 9 12 9 2 9 9 3 2 3 12 9 2 9 9 3 2 2
7 9 0 9 1 11 7 11
11 1 9 13 15 0 9 1 11 7 11 2
26 13 15 3 3 2 3 9 0 0 9 11 11 1 9 0 9 13 2 16 9 4 13 9 1 11 2
10 1 9 15 4 13 7 0 0 9 2
20 11 13 2 16 15 1 11 1 11 13 9 2 7 9 9 11 13 0 9 2
13 1 9 0 9 9 14 13 9 11 1 0 9 2
8 0 9 13 9 0 9 11 2
23 1 10 9 3 11 12 2 9 13 1 0 9 9 2 15 13 9 1 12 9 3 13 2
9 15 4 13 9 0 9 1 11 2
33 1 0 9 13 1 0 9 9 7 0 9 2 7 0 9 1 9 0 9 0 9 15 1 0 9 13 9 1 9 12 9 9 2
12 0 9 13 13 1 9 9 1 11 7 11 2
5 11 2 1 9 9
49 2 0 9 4 13 1 0 0 9 7 0 9 11 11 9 1 9 2 15 13 1 9 0 9 0 7 0 9 1 0 9 11 1 0 9 11 2 2 13 3 9 11 11 2 9 11 11 11 2
24 3 3 13 2 9 1 0 9 3 4 13 9 9 11 2 15 15 13 1 9 10 9 13 2
13 12 1 0 9 9 13 9 9 1 0 12 9 2
20 1 10 9 1 9 11 13 0 0 9 2 3 4 9 1 9 13 4 13 2
29 16 13 1 0 9 0 9 2 10 9 13 1 12 9 9 2 9 11 15 13 2 16 9 9 3 4 3 13 2
21 13 7 13 2 16 1 0 9 4 15 9 0 1 9 13 9 3 0 0 9 2
5 9 11 13 0 9
5 11 13 11 1 9
5 11 2 11 2 2
28 0 9 1 10 0 9 13 9 9 0 9 1 9 1 9 2 15 4 13 1 9 13 9 1 12 0 9 2
31 0 9 11 11 1 15 1 9 10 9 13 2 16 9 0 7 0 9 4 15 13 13 3 3 1 9 1 9 7 11 2
19 1 10 9 4 9 11 13 13 1 10 9 3 2 9 1 9 0 9 2
18 9 3 13 9 1 15 2 16 9 11 13 9 9 1 9 0 9 2
29 3 15 13 1 9 10 9 13 0 9 11 2 15 4 13 13 1 10 9 3 0 9 9 1 9 9 0 9 2
18 1 0 9 0 0 9 13 11 11 0 2 0 7 3 0 9 11 2
13 9 0 9 11 11 11 3 13 0 9 10 9 2
15 3 13 2 9 0 0 9 13 13 0 9 1 10 9 2
12 3 0 9 1 11 7 0 9 1 0 9 2
20 1 3 0 13 0 9 9 11 1 9 2 15 13 3 2 11 7 0 11 2
5 9 11 1 0 9
5 11 2 11 2 2
14 9 1 9 9 0 9 1 9 15 3 13 0 9 2
25 1 10 9 1 11 7 11 4 13 13 1 9 9 1 9 12 2 12 2 13 9 9 11 0 2
18 4 15 13 0 9 2 7 0 7 0 9 15 4 13 1 0 9 2
20 9 13 9 0 9 2 1 15 9 13 1 10 9 2 1 10 9 15 13 2
23 9 9 11 11 15 1 15 13 2 16 9 7 9 0 9 7 0 9 15 13 9 11 2
29 9 10 9 4 1 9 13 3 1 0 9 1 9 9 12 2 12 7 3 2 16 4 1 9 13 13 10 9 2
30 9 3 3 13 2 16 9 9 7 9 9 15 4 13 1 0 9 16 15 0 2 3 15 13 10 2 0 9 2 2
3 13 0 9
5 11 2 11 2 2
10 9 0 9 0 9 13 3 9 11 2
20 1 15 15 13 9 9 7 0 9 2 9 1 0 9 7 9 7 9 9 2
15 1 10 9 15 13 3 0 9 9 7 9 9 7 9 2
25 2 1 0 9 4 3 1 0 9 13 11 11 16 9 9 7 11 11 16 9 9 7 9 2 2
16 4 3 13 9 1 9 7 0 9 0 9 2 0 9 9 2
17 9 3 13 0 9 2 16 4 13 9 9 9 7 9 9 11 2
20 1 9 1 10 9 9 0 9 13 9 2 16 1 10 9 9 13 9 9 2
11 13 4 15 11 11 2 9 11 1 11 2
14 0 9 13 0 2 9 0 9 1 9 10 9 9 2
21 13 4 15 7 2 16 10 9 4 13 2 7 15 13 9 1 0 9 0 9 2
11 13 4 15 15 3 1 10 9 0 9 2
34 2 13 4 15 3 1 3 0 9 0 9 2 16 4 10 9 4 13 1 9 2 1 15 4 13 2 15 13 1 9 7 9 9 2
35 13 15 2 16 16 4 4 9 9 3 0 0 9 13 1 0 9 2 3 4 1 15 13 13 9 3 0 2 16 13 9 10 9 2 2
2 1 9
3 9 1 9
14 1 9 9 11 11 11 4 1 0 9 13 0 9 2
15 1 9 9 3 13 1 9 9 2 9 9 7 9 9 2
23 9 1 0 0 9 13 2 16 9 1 9 15 2 3 2 13 14 1 12 9 0 9 2
18 7 13 1 15 0 0 9 2 3 13 9 11 9 13 1 9 9 2
5 11 1 9 1 11
5 11 2 11 2 2
29 9 11 1 11 11 11 2 15 0 9 13 1 10 9 2 3 13 9 0 9 11 1 9 10 0 9 1 11 2
31 1 10 0 9 13 13 14 0 9 2 7 7 0 9 1 9 9 11 1 12 9 7 13 3 0 9 1 12 0 9 2
3 0 9 9
12 9 9 9 9 13 1 0 0 3 0 9 2
24 0 9 13 9 1 0 9 11 11 2 15 13 1 0 9 0 9 2 15 13 16 3 0 2
20 13 9 0 9 7 9 7 15 13 2 16 0 9 3 13 9 1 0 9 2
25 0 9 10 9 2 15 1 12 9 3 13 11 2 13 15 9 1 15 2 16 4 13 0 9 2
20 1 10 9 15 3 13 9 0 7 0 1 9 1 0 9 7 9 11 11 2
29 15 1 0 9 0 9 13 1 0 9 0 11 11 2 9 13 3 3 0 11 11 2 11 2 9 0 11 11 2
11 0 9 13 0 0 9 1 9 11 9 2
23 1 0 9 1 9 15 10 9 13 7 3 0 0 9 1 9 9 7 0 9 0 9 2
3 1 9 9
5 0 0 11 1 9
32 13 15 2 16 7 9 12 2 11 1 0 11 15 13 13 1 9 9 7 13 2 16 15 13 1 9 0 2 9 9 2 2
29 1 9 15 7 13 2 16 15 1 9 2 15 4 1 0 9 9 13 2 4 13 1 9 0 9 11 7 11 2
31 3 3 3 9 11 11 2 11 11 7 15 2 7 16 3 0 9 11 12 2 9 0 9 0 9 13 9 7 0 9 2
27 3 0 9 0 2 7 0 9 13 9 9 2 9 7 0 9 2 10 9 11 11 2 11 13 0 9 2
35 0 11 11 2 11 15 1 9 11 11 13 1 10 2 9 0 9 10 9 2 2 3 3 2 7 14 3 3 0 0 9 7 0 9 2
27 0 9 15 13 0 0 9 9 0 9 2 9 11 2 11 2 2 0 9 1 0 9 0 11 7 9 2
39 7 3 14 3 13 3 0 9 9 9 0 2 0 9 2 0 3 1 11 2 7 9 11 11 2 1 15 13 0 9 11 11 2 11 0 9 1 11 2
1 9
14 9 2 9 1 9 3 0 2 15 1 15 9 13 2
17 3 1 0 9 13 3 1 12 9 1 0 9 1 11 1 11 2
26 9 11 11 7 10 9 2 11 11 7 9 11 11 2 4 13 3 1 12 1 0 0 9 1 11 2
22 11 11 13 10 9 0 7 3 0 9 3 1 12 9 1 9 11 1 0 0 9 2
19 9 13 11 11 2 0 9 9 9 1 9 7 9 9 0 9 1 11 2
10 11 11 13 0 9 9 2 9 9 2
9 15 12 15 4 13 1 12 9 2
33 11 11 13 9 9 9 9 2 0 9 0 9 7 0 11 2 1 9 0 0 9 2 3 15 15 0 9 13 7 9 9 9 2
16 11 11 7 10 3 2 0 2 9 3 0 9 13 2 2 2
36 9 1 9 13 9 2 16 4 1 11 0 2 15 13 9 1 0 11 2 1 9 13 9 1 0 9 2 10 9 15 13 3 12 9 9 2
17 9 1 9 9 1 9 3 0 9 13 1 9 9 1 9 12 2
15 3 1 11 11 7 1 9 2 10 0 9 1 0 9 2
4 9 0 16 9
34 9 9 1 11 1 15 9 0 9 0 0 11 2 0 15 1 0 9 2 14 13 2 7 9 9 11 1 0 9 3 13 1 9 2
34 9 11 4 1 15 13 13 3 3 1 11 2 3 13 3 1 0 9 0 15 1 9 0 7 0 9 2 15 13 3 0 9 9 2
8 1 0 9 15 11 13 9 2
16 10 9 13 0 9 9 7 9 2 15 3 13 0 0 9 2
12 9 2 9 7 3 0 9 15 7 13 3 2
12 15 13 7 1 9 2 15 13 9 11 15 2
22 11 13 1 9 7 11 2 15 3 15 9 13 2 14 1 9 2 7 3 1 9 2
9 3 13 9 0 0 16 0 9 2
25 9 1 9 13 0 9 2 1 15 13 9 0 7 13 15 0 9 2 15 15 13 1 0 9 2
22 1 9 9 2 3 9 13 9 2 15 3 13 9 0 9 2 7 15 1 9 13 2
14 1 0 9 13 0 9 2 1 15 4 15 13 9 2
5 15 14 13 9 2
11 3 13 9 1 0 9 7 1 9 0 2
16 0 13 15 1 0 15 0 0 9 2 3 15 9 13 13 2
10 0 9 7 9 11 13 1 15 9 2
2 9 3
28 9 11 13 10 9 2 9 1 9 0 0 9 2 3 1 0 9 1 0 0 2 13 11 3 1 12 9 2
15 11 11 11 2 9 9 9 1 0 9 7 12 0 9 2
15 16 0 11 13 10 9 1 9 2 13 15 9 7 9 2
11 11 15 13 1 9 0 9 7 9 0 2
8 11 11 2 9 1 0 9 2
15 11 13 0 9 0 0 9 2 10 9 3 13 10 9 2
5 9 1 9 7 9
7 12 9 1 9 7 9 9
29 2 15 3 0 2 0 7 0 10 9 3 13 2 2 2 13 1 9 9 9 1 9 9 11 2 11 11 2 2
22 9 0 0 9 13 1 9 2 16 13 9 11 11 3 3 0 0 9 7 11 9 2
31 10 9 2 9 2 1 15 13 9 9 11 11 2 9 11 11 13 1 0 9 7 0 9 2 3 7 9 9 3 13 2
17 9 11 11 13 3 3 2 16 16 4 13 0 9 1 0 9 2
12 9 9 13 3 0 2 16 10 9 13 13 2
21 0 9 11 11 13 0 9 13 9 2 15 13 3 1 9 9 16 9 7 9 2
24 13 15 7 9 9 1 0 9 2 9 3 13 7 9 15 13 7 9 2 7 9 0 9 2
14 3 9 2 3 11 0 9 13 9 9 0 2 13 2
49 1 10 9 3 13 1 9 9 9 9 9 11 7 11 2 1 15 11 11 11 13 3 12 0 9 7 9 11 11 13 1 12 9 1 0 9 11 11 2 9 11 2 7 11 11 2 11 2 2
32 11 7 11 13 1 0 9 11 2 3 0 7 3 0 11 11 11 2 7 9 15 13 1 11 14 1 9 11 7 3 3 2
22 0 9 15 13 1 0 9 0 9 2 13 0 2 0 7 3 0 2 7 3 0 2
22 1 0 9 13 1 9 10 9 2 1 9 9 2 15 0 13 1 9 0 15 15 2
23 11 11 13 14 3 0 2 0 1 15 2 1 10 9 2 16 4 3 3 13 10 9 2
51 9 1 0 7 0 9 13 9 7 1 0 0 0 9 2 3 0 7 3 0 16 0 9 11 11 2 0 2 3 0 2 7 3 10 9 0 11 11 13 2 7 3 0 7 3 0 9 11 11 11 2
26 1 0 7 0 9 2 9 7 9 15 13 0 9 0 2 0 9 2 0 9 2 9 11 11 2 2
16 13 1 9 7 9 2 1 9 7 9 2 1 9 7 9 2
9 9 1 3 0 9 1 0 0 9
27 1 0 9 1 9 0 0 9 1 0 11 15 9 9 13 9 0 0 9 7 13 3 1 9 0 9 2
11 1 9 13 9 11 1 11 12 0 9 2
18 1 9 13 0 9 1 3 0 9 7 1 9 2 1 9 13 9 2
14 13 15 0 9 10 9 1 9 0 9 1 0 11 2
28 1 9 15 13 3 1 12 9 2 7 3 1 0 9 9 11 2 15 13 1 0 9 2 13 1 0 9 2
18 9 13 0 9 7 3 2 16 10 9 13 1 12 9 0 16 0 2
15 3 0 9 15 12 9 13 1 0 9 3 12 9 9 2
19 0 9 1 11 13 0 9 1 0 9 7 1 9 12 13 3 0 9 2
42 2 0 9 2 1 15 13 1 9 2 9 13 1 9 2 15 13 3 0 0 9 2 2 13 11 11 2 0 9 1 9 9 11 9 2 9 2 0 2 1 11 2
17 1 9 1 9 0 9 7 9 11 13 9 0 9 9 0 9 2
12 9 1 0 9 13 13 3 16 12 0 9 2
9 1 0 9 3 13 9 0 9 2
18 1 11 11 13 10 9 9 3 1 0 9 7 9 13 1 0 9 2
34 2 0 9 13 10 9 2 16 13 0 13 1 0 0 9 1 10 9 2 2 13 11 11 2 13 9 0 9 1 0 9 1 11 2
13 2 0 9 15 9 13 1 0 9 1 9 9 2
21 15 4 13 2 16 13 1 15 9 2 15 15 13 3 9 9 1 0 9 2 2
10 9 0 9 11 11 11 13 0 9 2
10 2 0 9 4 13 1 9 0 9 2
12 0 3 13 0 2 16 9 1 0 9 13 2
9 9 13 2 13 15 3 0 9 2
17 13 13 1 9 2 15 13 1 9 7 15 13 1 0 9 2 2
14 1 15 15 0 9 13 1 0 9 1 9 0 9 2
4 2 15 13 2
13 1 0 9 15 0 9 13 2 2 13 11 9 2
31 2 1 9 1 9 4 13 0 9 7 0 9 2 15 13 9 13 2 2 13 9 9 0 9 0 9 1 11 11 11 2
13 2 1 0 9 16 13 9 9 7 9 13 13 2
14 12 1 9 9 11 1 0 9 13 9 0 9 2 2
23 9 0 9 7 9 11 11 1 9 11 9 2 9 2 0 2 1 11 13 0 9 3 2
17 3 13 3 13 9 1 10 9 2 1 15 15 1 0 9 13 2
19 13 15 3 1 0 9 0 7 0 9 7 1 9 0 9 1 0 9 2
18 2 3 9 13 13 9 1 9 7 9 4 13 13 10 9 1 9 2
17 3 4 10 9 13 3 1 10 9 7 9 2 2 13 11 11 2
3 3 0 9
1 9
3 3 0 9
30 0 9 1 11 13 0 9 13 9 1 9 1 12 9 1 11 2 15 13 3 0 16 9 7 13 9 9 1 11 2
20 0 9 1 11 15 13 3 1 12 7 12 9 1 9 2 0 13 1 9 2
20 9 3 0 1 9 1 9 2 1 15 13 13 14 12 9 2 15 3 13 2
15 1 0 9 1 11 4 3 3 13 9 1 0 9 9 2
10 7 15 13 3 3 0 16 1 9 2
13 3 13 2 16 13 3 3 14 9 9 1 9 2
19 1 9 9 9 1 9 13 4 13 3 2 16 9 13 3 10 0 9 2
11 3 13 13 2 16 15 1 9 15 13 2
24 14 9 2 7 7 9 2 9 7 9 13 2 16 9 13 1 9 9 13 2 0 4 13 2
10 9 9 1 9 4 3 13 1 9 2
61 9 9 1 9 13 2 15 13 2 13 7 13 9 1 9 2 16 4 15 3 13 0 9 1 0 2 4 13 1 12 7 12 9 9 2 1 12 7 12 9 1 9 2 16 3 13 16 9 0 9 7 13 1 9 7 1 9 0 12 9 2
19 0 9 15 7 13 9 2 15 4 9 13 1 9 0 1 9 10 9 2
25 3 4 0 13 0 9 13 1 9 2 13 2 13 1 9 7 1 10 0 9 13 1 0 9 2
10 3 3 4 15 13 1 9 1 9 2
18 0 9 7 13 9 13 3 3 7 13 0 2 16 7 3 13 4 2
15 9 9 1 9 15 3 13 13 1 10 0 9 3 0 2
26 3 2 16 3 13 0 7 0 9 9 2 15 9 1 9 2 1 15 13 0 0 0 9 2 13 2
19 0 9 2 12 9 9 1 0 11 13 3 3 1 0 9 11 3 3 2
30 10 9 13 9 2 15 13 2 16 4 15 0 9 13 1 10 9 7 3 2 16 4 15 13 9 9 1 10 9 2
11 3 13 12 9 1 9 0 11 11 3 2
34 13 15 2 16 9 0 9 13 1 0 9 3 3 0 0 9 1 9 9 2 3 0 9 1 0 11 7 11 9 7 12 0 9 2
42 3 10 9 13 2 16 4 13 0 0 9 2 1 15 15 15 4 13 1 0 1 15 2 15 15 15 1 10 9 13 2 15 15 1 15 13 2 1 15 13 0 2
14 13 4 10 9 2 16 4 15 3 3 13 9 9 2
10 13 13 9 2 15 15 3 3 13 2
7 0 9 1 9 7 1 9
11 0 9 9 9 2 15 3 13 9 11 2
19 0 9 15 15 7 13 2 7 3 0 9 13 9 1 0 9 0 9 2
39 1 9 7 9 11 11 2 15 13 1 10 9 2 13 9 11 11 2 9 2 2 11 11 2 9 2 2 11 11 2 9 2 7 11 11 2 0 2 2
11 1 10 9 4 13 1 9 0 0 9 2
10 1 0 9 13 1 15 13 14 3 2
2 3 2
12 2 3 2 1 9 12 2 15 15 3 13 2
14 15 4 13 15 9 0 0 9 7 0 9 13 9 2
9 13 4 9 2 15 15 15 13 2
12 3 0 0 9 2 11 13 13 2 11 11 2
10 10 9 13 0 9 2 7 14 9 2
10 10 9 15 1 15 13 1 9 11 2
11 16 4 15 15 13 2 13 15 1 9 2
16 7 11 11 15 15 13 1 9 11 11 7 10 9 13 3 2
18 9 15 15 13 2 16 15 13 14 3 2 16 4 13 0 11 12 2
16 3 4 13 10 0 9 1 9 2 0 9 7 9 0 9 2
5 3 13 9 2 2
7 15 0 2 11 2 13 2
10 2 1 9 4 13 9 1 0 11 2
4 15 15 13 2
5 11 11 13 9 2
6 13 15 10 0 9 2
10 13 4 0 9 7 13 4 1 9 2
8 9 1 15 13 1 9 15 2
8 9 13 0 1 9 7 9 2
6 3 3 13 15 0 2
12 13 1 15 9 0 11 7 0 0 9 2 2
8 3 7 1 15 13 10 9 2
17 2 9 1 11 15 13 2 16 4 15 13 3 1 0 9 9 2
5 15 13 1 9 2
8 1 11 13 3 1 9 9 2
24 1 9 9 11 11 3 13 3 0 9 2 7 13 4 15 2 16 15 13 1 15 1 9 2
9 3 15 13 9 10 9 11 11 2
7 7 11 11 3 13 9 2
14 1 9 15 12 2 9 13 9 7 9 9 9 2 2
6 9 4 13 12 9 2
4 13 15 9 2
19 2 15 15 13 2 16 12 7 9 9 1 12 9 7 12 9 13 3 2
13 13 4 15 9 2 16 4 1 15 13 0 9 2
7 11 11 13 0 9 2 2
17 13 15 9 1 0 11 7 0 0 0 9 2 3 11 7 9 2
13 10 9 11 11 15 1 9 14 3 13 11 11 2
12 2 16 13 0 9 2 15 13 3 3 9 2
10 13 1 15 2 16 0 13 16 11 2
5 3 13 9 11 2
11 9 9 0 9 13 1 11 1 0 12 2
15 1 15 15 9 13 9 2 16 13 15 11 7 11 2 2
4 1 15 13 2
8 2 9 13 3 1 0 9 2
15 13 3 10 9 14 13 7 13 9 2 14 15 15 13 2
9 9 13 9 9 2 9 7 9 2
8 15 3 4 13 13 0 9 2
25 10 9 13 2 16 4 15 9 1 9 13 2 13 15 7 3 13 13 1 15 2 15 13 2 2
3 13 0 2
10 2 14 2 7 13 15 1 10 9 2
4 13 15 9 2
7 0 15 13 14 0 9 2
10 13 10 9 2 7 1 9 13 2 2
17 3 13 16 0 9 10 9 1 15 2 15 13 1 0 9 15 2
5 2 13 3 0 2
11 13 9 2 15 15 13 7 1 0 9 2
5 3 13 3 0 2
9 9 1 9 15 1 15 13 2 2
12 13 15 2 16 11 13 0 9 1 10 9 2
4 2 3 14 2
36 3 16 4 13 2 7 3 15 13 0 9 7 15 13 1 9 2 15 13 13 9 7 9 2 1 15 15 13 7 13 2 1 15 15 13 2
6 3 3 13 15 0 2
12 13 2 16 0 0 9 13 1 15 3 0 2
16 11 7 11 2 11 2 11 2 11 7 0 13 15 9 2 2
2 11 11
4 15 13 15 2
2 11 11
5 9 0 9 1 11
5 13 1 0 9 2
11 13 9 7 9 1 0 9 9 1 11 2
7 1 11 13 9 0 9 2
10 1 9 12 13 16 9 3 1 9 2
15 1 0 9 1 9 12 4 1 10 9 13 1 0 9 2
7 3 13 9 10 0 9 2
14 2 10 9 1 9 9 13 0 2 2 13 11 11 2
9 2 13 4 1 10 0 9 13 2
17 3 4 15 7 13 2 16 0 9 4 13 13 3 0 0 9 2
10 9 7 9 13 1 9 9 0 2 2
19 1 9 1 9 0 9 13 15 0 9 0 0 9 2 16 13 0 9 2
16 9 9 4 1 15 13 0 13 3 7 0 9 15 3 13 2
11 0 9 11 11 13 9 7 9 0 9 2
15 2 13 15 1 9 7 13 1 9 2 3 4 9 13 2
9 1 9 4 13 1 9 0 9 2
12 1 9 4 1 15 13 9 2 2 13 9 2
7 1 9 13 3 1 9 2
14 2 13 4 1 9 9 2 9 0 1 0 0 9 2
10 13 15 9 9 2 15 4 15 13 2
15 1 9 4 15 1 15 3 13 2 7 3 15 13 2 2
2 11 11
4 9 2 11 11
3 9 1 9
1 9
3 9 1 9
11 3 3 13 9 0 9 1 9 0 9 2
10 9 10 9 13 13 9 10 0 9 2
17 3 1 9 7 12 0 9 13 1 9 13 1 9 1 0 9 2
27 3 15 9 0 9 9 0 9 13 2 16 16 15 4 13 2 15 15 1 9 9 1 10 9 9 13 2
12 1 9 3 3 14 4 13 13 1 12 9 2
19 1 12 13 3 12 9 2 1 0 9 2 15 3 13 1 10 9 9 2
15 9 4 13 1 11 12 2 9 3 7 3 1 12 9 2
2 0 9
5 11 2 11 2 2
19 1 9 4 3 13 9 0 9 0 2 0 9 1 12 0 9 7 9 2
15 0 9 13 9 9 9 1 0 9 1 0 9 1 11 2
19 0 9 13 3 9 9 0 0 9 2 15 13 13 9 1 11 1 11 2
36 9 2 15 13 10 9 13 0 9 7 9 1 0 9 2 15 13 1 0 9 1 11 1 0 9 13 1 9 12 2 7 9 12 2 9 2
2 0 9
5 11 2 11 2 2
27 1 0 9 4 13 1 9 9 0 9 0 9 0 9 1 3 16 12 9 9 1 0 9 1 0 11 2
21 1 15 15 0 9 9 13 0 9 16 9 9 13 1 0 9 7 3 16 9 2
11 0 9 0 9 11 13 12 9 9 9 2
15 9 9 13 3 1 9 2 0 9 7 0 9 0 9 2
22 15 4 13 13 9 1 2 0 2 9 2 15 4 3 13 13 0 13 1 0 9 2
8 0 9 3 13 0 0 9 2
15 9 13 1 9 0 9 1 9 9 1 9 1 0 9 2
3 9 12 13
6 0 9 13 9 1 9
5 11 2 11 2 2
37 0 9 9 12 1 0 9 0 12 12 9 3 10 9 2 9 9 9 1 11 2 3 1 9 3 13 1 9 9 9 2 12 1 0 9 9 2
24 3 0 9 13 3 9 11 12 2 1 15 3 9 11 12 2 2 15 3 13 0 9 9 2
20 9 0 9 2 9 9 12 2 13 9 9 11 1 9 12 9 2 0 9 2
11 3 3 15 1 15 1 11 13 10 9 2
26 0 7 13 0 9 3 1 9 2 9 2 2 3 1 15 2 16 13 3 9 13 9 12 12 9 2
20 16 0 9 13 3 0 9 2 10 9 13 3 7 13 10 9 1 0 9 2
13 9 9 9 7 13 2 16 1 9 15 3 13 2
24 1 10 9 13 9 9 12 12 9 9 12 2 13 4 15 3 13 13 1 0 9 0 9 2
11 1 9 9 9 7 7 3 9 3 13 2
22 0 0 9 11 2 9 11 11 2 11 11 7 11 11 15 1 0 9 13 0 11 2
16 9 0 11 13 0 11 2 12 9 2 1 9 12 12 9 2
12 1 9 15 7 13 7 1 3 0 0 9 2
24 3 15 3 13 9 9 11 2 13 15 3 0 9 1 0 3 0 11 11 1 12 9 9 2
3 3 13 2
23 9 2 1 9 1 9 13 1 11 3 3 2 1 0 9 11 3 7 3 2 3 9 2
21 0 9 12 7 12 2 1 9 3 2 1 11 3 14 3 1 9 2 3 9 2
32 0 9 12 7 12 2 1 12 9 1 12 2 0 7 0 9 12 7 12 9 2 9 15 4 1 11 1 9 13 1 0 2
15 2 3 13 1 11 3 7 3 2 1 9 3 3 2 2
29 1 9 9 13 1 12 2 12 7 13 1 12 2 12 2 9 13 1 9 12 2 12 7 13 1 12 2 12 2
20 9 9 2 0 9 12 1 9 12 2 0 12 9 2 9 2 1 9 12 2
4 0 9 12 2
15 0 9 2 0 9 3 0 2 0 9 13 2 9 2 2
3 9 1 9
5 11 2 11 2 2
38 9 0 9 9 1 9 2 3 4 9 1 9 12 2 12 13 1 12 9 2 13 3 1 12 0 3 1 9 0 9 12 0 9 1 12 2 9 2
17 9 1 0 9 12 12 9 13 3 3 0 0 9 1 12 9 2
10 12 0 9 4 13 1 12 12 9 2
5 13 0 7 0 9
8 2 0 9 9 13 0 9 2
39 1 9 0 9 0 9 9 2 16 9 9 2 3 3 15 13 0 0 9 2 13 14 2 0 9 1 9 9 2 1 0 11 3 13 9 9 11 11 2
9 2 10 9 13 3 0 7 0 2
24 0 4 13 9 10 9 1 9 12 7 12 9 1 9 3 3 0 0 9 1 0 0 9 2
14 15 13 1 0 9 1 12 9 2 1 0 0 9 2
30 0 9 4 15 13 13 1 15 2 10 13 7 13 9 1 9 9 7 9 7 3 13 7 13 9 9 1 11 2 2
18 11 11 3 13 1 15 2 16 0 9 9 13 13 16 9 0 9 2
14 2 9 7 10 9 4 13 1 9 0 9 0 9 2
11 15 0 9 9 13 9 1 3 0 9 2
18 1 10 9 4 9 3 13 1 9 7 9 9 2 2 13 11 11 2
60 3 11 11 1 9 11 11 15 13 2 16 16 4 1 9 0 7 0 9 3 13 2 16 2 9 2 16 13 13 7 13 3 1 0 9 7 1 9 0 2 4 13 16 0 9 2 2 13 1 0 9 1 10 9 9 0 10 0 9 2
29 2 1 0 9 4 13 2 16 0 2 9 2 13 1 9 0 11 0 9 2 15 15 4 13 1 9 0 11 2
10 3 0 13 0 9 13 0 1 0 2
28 1 11 3 13 0 0 9 1 9 15 1 0 9 0 2 16 13 9 2 9 2 9 7 3 0 9 9 2
21 1 9 10 9 2 3 0 1 0 9 2 4 9 9 13 2 2 13 11 11 2
31 1 1 0 9 1 9 9 13 1 11 11 0 13 0 7 0 9 15 0 9 1 15 2 16 13 0 13 0 0 9 2
31 2 13 4 3 13 1 9 0 9 2 3 4 13 4 3 2 13 9 0 7 0 7 9 9 2 1 15 13 13 2 2
3 9 0 9
22 9 12 2 9 9 9 1 0 9 2 15 13 0 1 0 11 2 13 3 1 11 2
22 9 1 9 9 13 9 11 11 12 2 2 15 15 3 13 3 0 9 1 10 9 2
14 1 12 0 9 13 7 10 9 16 3 9 11 11 2
18 7 3 13 10 0 9 2 15 13 12 9 2 1 0 1 0 11 2
11 1 9 9 13 3 9 1 0 0 9 2
19 0 9 9 12 2 15 13 9 9 9 13 1 12 9 2 4 3 13 2
13 13 1 9 11 12 1 0 9 2 0 11 12 2
13 13 15 3 1 11 1 9 11 1 9 12 9 2
16 0 9 7 2 16 15 13 2 3 3 1 9 13 0 9 2
6 0 11 1 10 9 2
5 11 2 11 2 2
11 2 9 9 0 1 9 13 0 9 13 2
36 9 13 9 9 2 7 9 13 10 9 9 9 2 2 13 15 3 1 9 0 9 1 9 9 1 10 9 11 11 1 9 9 7 9 9 2
21 13 2 16 9 4 13 3 1 9 9 1 9 2 7 9 1 15 3 13 13 2
33 1 9 0 9 2 0 9 1 0 9 9 2 15 13 9 9 2 7 0 9 15 3 13 13 1 0 9 2 15 13 0 9 2
22 1 9 1 9 9 9 1 9 0 9 13 3 0 0 0 9 0 9 11 1 11 2
17 1 9 3 13 9 1 9 2 10 3 0 9 4 13 1 9 2
30 1 9 0 9 15 1 9 0 9 13 9 1 12 7 12 9 2 1 11 2 11 2 11 7 10 0 9 1 15 2
8 9 13 1 0 9 1 11 2
11 9 1 0 9 9 1 0 11 1 11 2
15 9 9 9 1 9 1 10 9 13 1 9 0 9 9 2
6 1 11 1 9 11 2
27 0 9 11 3 1 9 9 11 11 13 10 9 9 12 2 12 13 1 11 1 9 11 11 2 11 11 2
33 3 13 11 11 2 9 9 0 9 11 11 2 9 11 1 0 9 13 1 10 9 12 9 1 0 9 12 9 1 9 1 11 2
15 2 0 9 15 7 13 9 13 2 2 13 11 2 11 2
18 3 13 2 16 1 0 9 4 1 11 9 11 13 12 0 9 11 2
25 2 16 9 4 11 13 1 9 7 2 15 13 9 0 9 2 13 9 9 11 9 9 13 2 2
20 9 9 0 0 9 11 11 1 9 13 1 0 9 11 11 11 11 10 9 2
31 2 0 9 2 15 13 1 9 1 10 9 2 15 13 9 11 11 2 13 9 1 10 2 16 4 4 13 1 0 9 2
11 13 15 7 9 0 10 9 1 11 2 2
4 9 13 10 9
7 11 2 11 2 11 2 2
38 3 3 13 0 9 13 7 3 7 13 9 0 2 9 1 11 2 16 0 9 13 0 9 2 15 14 13 13 9 0 2 9 1 0 9 0 11 2
16 9 9 4 3 13 7 9 9 10 9 1 0 9 1 11 2
12 3 1 10 0 9 13 3 9 0 0 9 2
28 1 10 9 15 0 2 0 9 1 11 11 11 13 2 16 0 9 9 11 1 9 11 13 1 0 9 13 2
28 9 15 13 3 13 1 11 2 7 16 13 3 9 11 2 4 9 13 1 9 11 2 15 13 7 0 9 2
22 1 9 12 2 9 2 15 3 13 10 9 1 9 2 13 9 9 11 10 0 9 2
24 2 13 9 9 2 16 4 9 9 7 10 9 13 2 2 13 15 0 9 11 11 11 11 2
6 9 11 13 4 1 15
23 1 0 0 9 11 2 3 13 7 0 0 9 2 13 1 9 1 0 9 1 0 9 2
8 13 15 1 15 1 9 11 2
8 1 0 13 1 9 1 11 2
15 3 15 13 13 9 2 7 16 9 13 1 10 0 9 2
10 1 9 1 11 15 3 13 0 9 2
7 15 15 14 13 1 9 2
11 15 15 7 3 13 13 2 15 13 9 2
9 9 13 9 9 7 3 14 13 2
6 1 9 13 3 0 2
7 7 3 13 10 9 13 2
22 13 15 7 13 9 1 9 2 2 0 15 13 7 1 0 9 2 16 13 1 9 2
6 13 1 0 9 2 2
16 13 15 3 1 0 9 2 1 15 15 13 3 1 9 11 2
11 13 14 1 0 0 9 0 9 9 11 2
10 3 15 13 9 2 0 9 13 2 2
8 13 15 9 7 13 1 9 2
21 2 10 9 13 3 3 7 1 0 2 3 15 13 13 2 2 13 9 9 11 2
16 2 0 13 15 1 9 2 15 13 0 3 1 0 9 2 2
14 9 9 13 3 3 1 9 2 16 4 13 1 9 2
16 16 10 9 13 3 0 9 2 3 9 13 7 9 1 9 2
19 1 0 13 1 11 2 9 7 1 0 9 1 11 13 10 12 0 9 2
18 16 15 13 1 10 9 2 1 9 13 0 9 9 2 3 15 13 2
3 9 7 9
4 3 7 1 15
3 9 7 9
22 13 4 0 7 0 9 2 16 4 13 9 12 9 0 9 7 12 9 0 9 9 2
20 11 2 11 2 9 0 2 0 9 9 9 2 9 12 9 2 9 12 9 2
17 0 9 2 9 0 2 9 11 2 9 12 9 2 9 12 9 2
15 11 2 9 0 2 9 11 2 9 12 2 9 12 9 2
18 11 2 0 9 2 0 9 9 11 2 9 12 9 2 9 12 9 2
16 11 2 9 0 2 9 11 2 9 12 9 2 9 12 9 2
20 11 2 11 2 9 0 2 0 9 9 11 2 9 12 9 2 9 12 9 2
7 3 15 13 1 0 9 2
13 13 15 13 9 7 9 2 10 0 9 15 13 2
2 9 0
9 9 9 0 9 11 2 11 11 11
10 2 12 1 9 10 9 13 0 9 2
20 16 15 13 9 9 1 0 11 7 0 9 2 13 9 1 10 9 14 11 2
6 3 9 3 13 0 2
25 9 1 0 9 15 13 9 14 1 15 2 16 15 0 9 13 9 1 0 9 12 9 1 9 2
20 1 0 9 2 3 15 9 13 13 9 14 12 9 1 9 2 13 7 9 2
22 0 0 9 15 1 9 9 13 3 13 7 13 0 2 16 4 13 0 9 13 2 2
2 13 9
3 9 1 9
2 13 9
14 12 9 13 1 0 9 0 9 0 9 1 0 11 2
11 9 2 15 13 2 3 3 13 1 9 2
8 13 15 2 14 15 13 9 2
2 13 2
7 13 15 13 7 13 9 2
11 13 15 14 12 9 9 2 9 2 9 2
12 1 9 13 13 9 9 9 2 15 13 3 2
6 7 1 15 13 9 2
16 16 3 15 13 2 16 15 13 2 13 15 9 1 0 9 2
16 3 0 9 12 9 13 1 9 9 7 13 2 16 15 13 2
7 0 7 3 13 9 13 2
14 9 15 13 2 16 4 15 15 13 3 13 1 9 2
16 1 12 0 9 15 12 9 13 9 13 7 9 13 13 9 2
16 12 1 9 4 13 2 15 13 10 0 2 15 9 13 13 2
5 0 10 9 13 2
19 12 1 15 1 9 13 13 2 0 15 13 7 9 13 3 16 0 9 2
7 1 9 7 10 9 13 2
15 13 2 16 15 13 14 3 2 16 4 13 1 9 9 2
21 13 13 2 16 1 0 9 13 1 9 1 9 7 3 1 9 9 3 13 9 2
19 7 1 10 9 9 12 9 13 1 0 9 9 2 9 7 9 0 9 2
22 11 11 2 2 15 13 3 3 0 2 0 9 1 11 13 1 12 7 12 9 9 2
10 10 9 11 11 2 13 1 9 3 2
15 12 15 1 9 13 2 0 9 7 1 0 9 9 13 2
2 0 9
9 13 9 10 0 9 0 2 9 2
9 11 11 1 12 2 9 9 12 2
13 9 13 13 7 9 0 9 7 9 1 0 9 2
6 12 2 9 1 0 9
21 9 9 2 9 2 0 9 2 9 0 9 2 9 2 9 2 9 7 0 9 2
6 12 2 9 1 0 9
22 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 7 0 2
4 12 2 0 9
24 9 9 2 0 9 2 9 0 9 3 2 0 9 2 9 1 0 9 9 9 2 7 0 2
6 12 2 9 1 0 9
37 9 9 2 12 2 7 12 2 9 2 9 9 2 9 2 0 9 9 2 9 9 2 9 1 9 2 9 9 2 9 9 2 9 9 7 0 2
6 12 2 9 2 0 9
5 9 2 9 2 9
9 12 2 9 2 0 9 2 0 9
44 9 9 0 9 2 9 0 9 2 9 9 2 9 1 9 9 2 9 0 9 2 9 2 9 2 9 9 2 9 2 9 2 9 2 9 1 9 2 9 2 9 7 0 2
14 0 9 13 1 0 9 7 1 0 9 0 2 9 2
11 11 2 9 12 2 12 2 12 2 12 2
21 0 0 9 2 15 1 9 9 1 9 0 11 1 9 0 9 3 13 1 9 11
32 1 11 13 1 11 11 1 9 1 10 0 9 0 0 0 9 11 11 12 2 12 7 0 1 9 0 0 9 0 9 9 2
18 13 15 3 0 9 9 2 0 2 9 2 15 3 13 3 0 9 2
21 16 0 9 11 3 1 9 3 1 11 11 13 2 13 10 9 9 12 9 9 2
3 2 11 2
3 11 13 9
13 9 11 15 13 1 2 9 9 2 1 0 11 2
34 9 1 15 2 16 11 13 9 13 11 2 16 4 13 9 12 9 7 9 0 1 12 9 1 9 1 0 9 2 13 1 0 2 2
19 15 13 11 11 7 3 13 2 16 15 13 1 12 1 10 9 0 9 2
7 1 9 15 13 9 9 2
21 3 3 2 12 9 2 13 11 2 13 11 2 11 11 2 11 2 11 2 11 2
8 3 13 10 9 0 0 9 2
17 11 13 1 9 11 11 2 0 9 11 7 12 2 9 0 9 2
24 15 0 15 13 13 3 1 2 9 9 2 2 3 4 13 0 9 11 1 11 1 0 11 2
18 2 1 10 9 11 4 13 3 2 16 4 15 13 9 1 15 13 2
4 3 14 3 2
12 16 4 3 13 2 10 9 4 15 11 13 2
17 2 13 15 12 2 3 13 2 16 3 1 11 2 7 0 9 2
8 13 4 15 1 9 1 11 2
14 2 13 4 2 16 1 15 2 11 7 11 4 13 2
12 3 1 11 2 11 2 11 4 15 3 13 2
15 7 3 7 1 0 9 1 0 9 1 0 9 0 9 2
7 3 1 10 0 9 2 2
12 13 15 13 2 3 4 9 11 1 11 13 2
7 2 11 13 13 10 9 2
11 16 13 1 9 1 9 2 11 15 13 2
8 7 13 3 0 9 1 9 2
16 11 3 13 3 13 1 15 2 16 9 4 13 14 12 9 2
31 2 11 4 13 9 1 0 9 1 12 9 0 2 15 13 1 0 9 1 12 9 3 2 16 16 4 13 1 0 9 2
4 13 15 11 2
7 2 11 13 9 12 9 2
14 1 10 9 13 0 9 3 2 16 1 9 13 3 2
14 4 1 15 13 7 1 11 2 7 1 15 0 2 2
11 1 9 10 9 4 13 11 13 0 9 2
7 2 3 1 9 1 9 2
16 7 3 7 1 11 2 7 15 4 13 4 10 9 13 3 2
12 3 4 15 13 13 1 0 9 12 9 9 2
6 3 4 13 13 3 2
14 14 1 9 2 3 1 9 2 7 3 1 0 9 2
10 12 9 1 0 9 4 3 13 15 2
7 3 9 1 15 13 2 2
13 3 0 13 13 2 3 2 9 9 2 3 13 2
23 0 13 14 15 2 16 9 15 13 13 1 9 1 9 9 9 9 7 0 3 13 3 2
2 11 11
4 9 2 11 2
2 11 11
5 1 0 9 1 9
7 11 1 11 1 0 9 11
16 3 0 9 0 0 9 13 1 9 9 11 2 11 1 11 2
26 13 15 1 9 7 0 9 11 11 13 1 9 1 11 7 11 2 1 9 4 13 11 7 11 11 2
24 0 9 11 13 3 1 0 9 0 0 11 2 15 13 1 9 7 3 1 11 7 1 9 2
13 11 13 9 9 0 9 11 2 1 15 13 11 2
20 1 9 13 0 9 9 2 16 0 11 13 13 1 11 0 9 1 0 0 2
13 3 0 9 11 2 11 13 0 9 1 0 9 2
15 13 15 1 11 1 3 0 0 9 0 9 11 2 11 2
18 1 9 13 0 9 2 0 9 9 12 9 4 1 15 12 9 13 2
23 0 9 11 2 11 2 15 1 9 3 13 11 2 3 1 0 9 2 2 7 13 9 2
48 13 15 7 9 1 9 1 0 9 9 1 0 9 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 0 11 2 11 2 11 7 11 2 0 11 2
2 11 13
21 11 3 13 1 9 12 0 9 11 2 3 15 7 4 13 1 15 3 9 13 2
5 11 13 0 9 2
12 3 3 3 9 9 13 1 9 1 0 9 2
7 0 9 11 13 9 11 2
19 11 3 1 9 1 0 2 11 3 13 2 7 3 10 9 9 11 13 2
29 0 12 9 0 9 9 11 2 11 1 9 1 0 11 13 11 11 2 11 11 2 1 11 11 1 11 7 11 2
14 3 3 13 11 2 11 11 2 1 9 12 2 2 12
24 1 9 13 3 0 9 11 2 12 2 11 2 12 2 11 2 2 0 13 11 2 11 2 2
23 10 11 7 11 2 12 11 2 13 1 9 0 7 0 9 7 3 13 0 7 0 9 2
3 9 1 11
15 2 13 0 1 9 13 2 3 15 11 11 13 1 9 2
8 13 15 13 10 9 7 9 2
28 13 7 2 16 1 15 13 4 13 0 0 9 2 2 13 1 0 9 1 0 11 9 11 11 1 0 9 2
16 1 9 9 0 9 11 15 9 13 0 9 1 0 9 9 2
14 9 1 15 1 9 13 9 2 15 11 3 13 9 2
19 11 2 2 1 0 9 13 15 3 3 3 2 16 16 4 13 1 9 2
16 1 0 9 15 13 13 2 1 9 7 13 3 7 9 2 2
5 11 3 1 9 13
3 9 1 9
12 11 3 1 9 13 11 2 2 1 10 9 2
15 0 11 13 0 9 1 0 9 12 1 9 12 2 9 2
13 9 13 1 9 9 12 2 3 4 13 0 9 2
12 16 0 9 15 4 13 1 9 3 9 9 2
8 7 10 3 13 9 1 11 2
17 0 7 13 2 16 1 9 9 15 13 9 13 1 11 3 12 2
15 7 1 0 9 1 0 9 15 9 1 9 11 13 3 2
21 2 11 11 15 3 13 16 0 9 1 9 2 2 13 0 9 11 11 11 11 2
17 9 11 11 13 1 11 1 11 2 3 4 3 1 11 13 2 2
9 13 12 9 2 13 10 0 9 2
5 15 1 15 11 2
9 2 7 15 13 9 2 7 9 2
10 12 9 13 1 9 0 2 2 2 2
11 1 11 13 1 11 0 0 9 11 11 2
15 9 11 13 2 1 0 9 11 11 2 9 1 9 0 2
10 1 9 13 7 11 11 2 11 2 2
13 0 9 11 11 13 9 1 9 0 9 11 11 2
9 1 0 9 1 11 13 12 9 2
10 1 9 7 13 1 9 2 15 13 2
12 13 2 16 1 0 9 13 1 12 12 9 2
18 2 1 11 1 11 13 3 12 7 9 9 9 1 9 2 2 2 2
9 1 11 13 9 9 9 11 11 2
14 2 13 13 9 2 2 13 0 9 7 0 9 11 2
15 0 3 13 2 16 11 13 1 9 9 1 9 1 11 2
10 2 3 10 9 13 2 2 13 11 2
17 1 11 13 2 16 11 11 15 1 11 3 13 2 13 7 3 2
13 13 15 2 16 9 9 11 4 11 13 3 3 2
13 3 15 9 0 9 1 0 9 13 9 1 11 2
12 3 3 11 13 9 1 11 12 3 9 9 2
10 11 3 13 1 9 1 9 13 2 2
2 9 0
13 11 11 7 11 11 15 13 9 0 2 9 9 2
13 13 1 15 0 2 9 9 1 9 0 0 9 2
28 0 0 9 11 7 0 9 11 13 1 9 11 11 16 0 0 3 13 9 7 13 9 1 9 12 1 11 2
12 11 2 1 9 13 1 9 0 9 1 9 2
54 1 9 15 13 1 9 11 2 11 2 11 2 11 2 11 2 11 2 2 11 2 11 2 11 2 11 2 1 0 11 2 9 1 9 2 7 1 3 0 9 11 2 11 2 11 2 2 11 2 11 2 11 2 2
16 13 15 7 0 12 9 1 9 1 0 9 9 1 0 9 2
4 9 2 2 2
13 11 2 2 13 4 10 9 2 9 1 0 9 2
15 10 0 9 13 2 16 4 3 1 0 9 13 12 9 2
16 9 1 0 12 9 9 13 0 9 10 9 1 3 0 9 2
11 0 13 1 12 9 2 9 13 13 0 2
12 3 15 13 11 2 10 0 9 13 11 2 2
8 11 2 2 9 9 13 9 2
8 1 15 9 2 16 9 13 2
6 9 13 9 10 9 2
12 3 7 13 13 2 16 0 9 13 0 2 2
5 2 2 2 7 9
20 11 2 2 1 0 9 13 3 10 9 2 15 15 3 13 3 1 9 2 2
18 11 2 2 3 4 13 1 0 9 2 16 15 13 14 12 2 12 2
9 1 10 9 9 1 9 13 2 2
15 11 2 2 0 9 15 1 15 13 2 3 4 15 13 2
18 3 15 7 13 9 1 9 7 15 2 16 4 15 13 1 0 9 2
11 3 3 15 13 1 10 0 9 0 2 2
12 9 1 0 9 13 1 9 9 9 0 9 11
2 1 9
19 0 9 1 11 11 11 15 13 1 9 1 11 9 9 1 9 9 9 2
19 11 1 9 1 9 4 13 3 9 11 7 9 11 2 3 13 1 11 2
25 11 11 2 12 2 2 0 0 9 9 1 9 2 15 1 12 9 13 1 0 9 1 0 11 2
11 3 0 2 13 15 1 9 0 0 9 2
17 1 0 9 15 7 1 15 13 9 0 9 2 9 9 7 9 2
28 9 11 2 11 11 0 11 2 15 1 0 9 1 0 11 1 0 9 1 9 13 9 7 12 9 4 13 2
19 0 13 2 16 15 3 13 3 3 2 3 1 9 9 13 1 0 9 2
62 9 13 9 0 9 2 0 9 9 2 9 2 2 12 2 9 0 9 2 1 9 13 7 11 11 2 11 11 2 11 11 2 11 11 7 11 11 2 11 2 12 9 13 1 11 1 12 9 2 2 0 9 2 1 11 1 9 1 12 9 2 2
33 9 0 9 9 11 11 2 0 11 11 2 2 13 1 0 9 9 9 1 11 11 11 2 0 9 11 15 13 9 0 9 2 2
16 1 9 11 11 2 0 9 0 9 2 15 13 3 12 9 2
14 1 12 0 9 15 13 10 0 9 3 16 12 9 2
4 11 2 11 2
9 11 2 11 2 2 11 2 11 2
17 11 2 11 2 2 9 2 0 2 0 2 2 2 11 2 11 2
1 11
9 0 0 0 9 13 12 2 9 2
7 0 9 13 1 9 0 2
3 9 1 9
18 9 11 7 11 2 12 0 9 2 3 13 12 2 9 0 0 9 2
18 3 13 1 11 2 3 13 3 1 9 0 11 7 11 1 0 11 2
4 11 11 2 2
3 11 11 2
2 1 9
14 11 13 3 1 9 11 1 0 0 9 1 11 11 2
14 9 15 9 0 11 2 11 2 13 9 9 11 11 2
8 9 13 1 0 9 3 0 2
8 9 1 9 1 0 0 9 2
29 11 2 12 2 9 2 13 1 11 1 10 9 1 12 2 9 12 2 12 7 12 9 1 9 3 12 2 12 2
10 3 3 9 3 13 1 12 2 12 2
14 0 11 13 9 11 11 2 12 2 0 1 9 11 2
5 9 13 9 1 9
30 9 2 1 9 11 2 11 2 15 1 9 13 1 9 1 9 9 1 9 0 9 2 7 0 9 13 16 1 9 2
8 1 11 11 3 13 7 9 2
25 12 2 9 2 11 2 11 2 11 12 2 12 2 9 11 11 13 1 12 2 9 2 9 11 2
2 9 2
4 13 9 1 11
24 3 13 4 9 9 11 11 11 11 2 12 2 1 3 0 9 1 11 2 12 2 12 2 2
14 2 13 2 3 15 3 0 9 3 13 2 2 13 2
32 1 9 9 2 15 13 1 0 12 0 9 1 9 3 1 11 7 1 11 2 13 2 2 4 13 13 12 9 1 9 2 2
7 1 15 3 13 9 9 2
9 2 9 13 15 7 15 13 15 2
21 16 9 1 15 13 2 16 15 13 9 7 16 4 13 13 2 3 15 15 13 2
9 1 9 15 13 7 13 15 9 2
9 15 7 1 9 1 11 13 2 2
9 10 4 3 13 0 9 1 9 2
22 2 1 0 9 13 1 9 12 12 9 2 1 15 15 13 13 12 9 7 12 9 2
16 11 1 11 13 12 9 2 13 9 2 13 12 9 9 2 2
7 15 13 3 15 2 2 2
31 2 7 0 9 13 15 7 9 1 9 2 15 13 12 9 7 9 2 15 13 9 7 9 13 2 13 3 12 9 9 2
17 7 9 1 9 2 15 13 1 9 2 13 3 12 9 9 2 2
15 11 11 16 0 9 13 0 9 2 13 15 3 0 9 2
23 2 15 13 9 1 0 9 2 3 13 11 1 9 2 7 11 4 3 13 13 1 15 2
13 3 11 13 2 16 15 13 13 2 15 7 13 2
17 13 9 9 2 15 15 13 9 7 9 9 13 9 1 9 2 2
17 10 13 9 1 0 9 9 1 11 7 3 1 0 9 1 9 2
9 2 10 0 9 10 9 3 13 2
11 13 15 15 2 16 15 3 13 0 9 2
35 15 15 3 1 9 13 2 14 13 15 9 11 2 14 13 15 11 7 0 9 2 15 3 9 1 9 13 7 14 15 13 1 10 9 2
9 13 15 3 1 9 7 13 9 2
29 14 1 0 9 13 3 11 2 7 16 15 3 13 3 0 9 2 15 3 13 1 0 9 2 3 13 15 9 2
13 3 15 13 1 9 10 9 11 1 0 11 11 2
28 2 9 11 2 15 13 1 11 2 13 0 9 7 13 13 11 2 16 13 9 2 1 15 15 13 1 9 2
17 10 9 11 0 13 7 3 15 2 15 13 9 11 11 2 13 2
11 3 13 9 7 15 15 13 1 9 2 2
15 3 15 13 1 11 11 2 15 15 15 13 1 11 11 2
32 2 16 4 4 13 2 16 11 13 3 9 1 11 2 16 4 3 13 9 2 3 15 9 11 13 3 2 16 13 1 11 2
15 13 15 1 9 1 0 0 9 2 7 13 13 3 0 2
14 15 15 15 3 13 7 15 15 13 13 1 0 9 2
12 10 9 13 0 7 1 9 15 15 13 2 2
6 13 0 9 10 9 2
17 2 3 2 13 4 15 0 9 0 9 7 13 9 1 0 9 2
11 13 13 9 2 15 4 1 11 13 9 2
12 15 11 13 0 1 15 2 16 3 13 2 2
8 16 7 13 10 9 2 2 2
7 2 15 13 2 10 9 2
20 1 0 9 13 3 1 0 9 0 9 2 15 13 0 9 7 13 13 2 2
2 0 9
7 9 2 12 2 2 12 2
9 9 2 12 2 9 12 1 9 2
35 9 2 12 2 11 2 11 2 2 12 2 11 2 11 2 2 12 2 11 2 11 2 2 12 2 11 2 11 2 7 11 2 11 2 2
6 12 9 13 12 9 2
20 9 1 9 2 11 2 11 2 7 0 2 11 2 2 12 1 12 2 9 2
23 9 2 12 5 12 9 2 12 5 12 9 2 2 12 5 12 9 2 12 5 1 9 2
9 9 2 12 2 9 12 1 9 2
21 1 9 1 9 11 11 2 12 2 2 15 1 10 0 0 9 13 1 11 1 11
9 3 4 16 15 0 13 1 9 2
15 2 3 15 13 11 2 3 4 13 2 7 11 15 13 2
11 3 4 13 1 0 9 2 1 9 13 2
16 3 13 13 2 16 16 13 0 9 2 11 15 0 9 13 2
2 9 2
13 9 13 15 3 4 13 2 7 13 4 13 9 2
9 13 3 3 9 2 3 1 9 2
9 12 9 1 12 9 13 15 2 2
2 9 9
2 11 2
7 11 12 2 12 2 2 2
12 11 2 11 2 2 2 2 3 4 13 9 2
9 9 13 9 11 7 9 11 2 2
12 11 2 11 2 2 2 2 13 4 1 9 2
4 3 13 9 2
8 1 3 13 1 12 9 2 2
2 11 2
7 11 12 2 12 2 2 2
21 11 2 0 2 2 2 2 11 13 0 0 9 1 0 9 2 13 15 9 11 2
10 10 0 1 0 9 13 13 3 2 2
16 11 2 9 2 2 2 2 0 13 9 1 12 10 9 2 2
2 11 2
9 0 2 11 12 2 12 2 2 2
25 11 2 0 2 2 2 2 1 0 0 12 2 3 15 1 9 13 9 2 3 4 13 10 9 2
14 9 15 13 0 11 9 2 15 13 1 15 9 2 2
19 11 2 0 2 0 2 2 2 2 0 9 1 9 9 1 0 9 13 2
12 3 15 13 9 1 0 9 2 3 0 9 2
26 1 9 1 11 15 14 11 1 0 11 13 2 1 11 7 0 11 11 15 13 3 12 2 12 2 2
2 11 2
7 11 12 2 12 2 2 2
21 11 2 0 2 2 2 2 12 12 4 13 1 9 2 14 1 9 15 15 13 2
6 9 4 13 0 2 2
20 11 2 11 2 2 2 2 1 12 9 13 9 2 16 13 9 1 0 9 2
18 3 13 11 2 1 9 9 13 9 11 2 15 13 1 9 11 2 2
3 13 4 15
20 0 9 0 9 9 11 2 11 2 9 12 2 12 7 9 11 1 0 9 2
19 1 10 9 0 9 13 0 9 2 9 9 15 13 12 9 11 7 11 2
13 3 7 13 9 0 9 2 13 9 1 10 9 2
6 1 9 13 12 9 2
18 16 11 13 1 9 9 2 13 4 14 0 13 1 9 14 1 9 2
3 9 1 9
6 13 9 9 11 11 11
9 2 13 4 9 12 3 0 9 2
24 1 0 9 13 1 9 9 0 12 2 12 2 3 12 2 12 7 0 12 13 12 2 12 2
5 15 13 3 9 2
14 0 11 13 0 9 16 3 2 9 3 13 7 13 2
17 7 3 10 0 9 1 11 2 3 11 13 0 9 12 2 12 2
27 7 3 15 13 3 0 9 2 1 0 12 14 12 2 12 7 1 0 13 11 1 12 9 12 0 9 2
17 3 15 15 13 2 3 9 3 0 9 13 7 10 9 13 13 2
12 15 13 1 10 9 3 0 2 9 0 9 2
5 0 9 3 13 2
14 15 7 13 9 3 0 7 0 9 7 0 9 9 2
9 1 15 13 3 11 13 12 9 2
24 0 9 13 1 0 9 9 1 0 9 2 3 13 13 0 0 9 7 13 0 9 9 2 2
1 9
4 9 1 0 9
35 0 0 9 9 0 9 1 11 2 11 2 11 7 11 13 2 16 9 9 11 13 3 3 0 2 3 15 13 9 9 1 11 7 11 2
22 1 9 9 11 1 11 11 11 15 9 0 9 13 13 9 9 0 9 1 0 9 2
15 15 4 15 13 13 3 9 1 0 9 0 7 0 9 2
19 9 15 13 1 9 0 0 9 2 15 4 13 1 9 10 9 13 15 2
24 2 3 4 13 1 15 2 16 4 13 13 1 9 1 0 9 1 11 2 2 13 11 11 2
20 16 0 9 0 9 1 9 0 9 7 11 13 0 2 3 13 0 9 11 2
13 1 9 0 0 2 0 9 15 3 13 0 9 2
24 9 13 1 15 2 16 13 9 11 11 13 3 0 9 7 13 9 1 0 11 1 0 9 2
18 7 15 4 13 1 0 9 0 2 7 9 4 13 13 0 0 9 2
13 3 15 2 15 13 0 9 1 0 9 1 9 2
2 9 9
2 13 4
2 9 9
10 9 13 9 2 9 13 1 0 9 2
32 0 9 11 11 13 9 1 9 7 9 2 15 13 13 9 9 2 15 1 10 9 13 3 2 3 2 2 3 4 13 13 2
6 10 9 13 14 11 2
16 0 9 13 1 10 0 9 13 7 13 9 1 9 9 9 2
24 9 7 13 2 16 4 15 12 9 9 2 0 0 9 11 7 11 2 3 13 1 9 9 2
28 13 15 9 1 15 2 16 2 0 2 13 13 9 1 9 2 1 15 9 13 9 13 9 9 1 9 9 2
30 10 0 9 3 11 7 11 13 13 9 9 9 2 1 9 3 0 9 7 13 3 0 9 2 7 3 7 9 9 2
14 0 9 1 11 7 11 7 13 9 7 1 15 3 2
23 11 2 15 10 9 1 2 0 0 9 2 11 9 9 13 2 13 3 13 3 3 0 2
30 1 0 9 15 11 13 3 7 0 9 2 0 0 9 2 0 9 9 2 7 3 0 9 2 3 1 9 0 9 2
17 15 13 3 0 9 2 15 1 11 11 7 10 11 3 13 9 2
4 10 9 1 11
2 11 2
21 1 9 9 9 11 4 1 10 9 11 11 13 10 9 2 15 4 13 0 9 2
14 3 3 13 2 9 7 9 13 1 9 0 9 9 2
42 11 2 11 3 13 1 9 0 9 1 9 0 9 1 0 0 9 11 11 2 15 1 9 13 2 16 2 11 3 13 10 0 9 7 1 9 10 9 13 11 2 2
30 2 13 1 15 2 16 16 4 15 1 11 10 9 13 2 11 11 4 1 15 9 3 13 2 2 13 11 2 11 2
4 3 13 9 9
1 9
4 3 13 9 9
13 1 9 13 0 9 11 1 9 9 9 1 11 2
24 0 9 9 9 11 11 11 4 15 13 2 15 13 9 1 9 11 2 15 13 3 11 13 2
13 2 1 10 9 13 2 16 4 15 13 13 11 2
16 15 15 13 0 2 16 4 1 9 9 11 13 9 9 11 2
16 13 15 7 9 9 7 1 9 15 1 15 3 4 13 2 2
14 9 0 9 7 9 11 3 13 13 15 1 9 9 2
26 2 10 9 13 10 9 2 9 1 9 7 9 3 13 2 16 4 9 13 1 9 9 11 9 11 2
8 1 15 4 9 13 4 13 2
14 3 15 13 9 9 2 16 9 13 10 9 13 2 2
5 0 9 1 11 13
5 11 2 11 2 2
27 0 9 1 0 9 0 11 11 3 1 9 1 9 0 9 11 13 2 16 10 9 1 9 11 13 0 2
29 12 1 9 13 9 0 2 0 9 2 7 15 7 1 9 2 16 1 11 13 3 12 9 9 0 7 0 9 2
13 9 1 9 13 2 1 10 9 2 10 0 9 2
22 9 3 13 9 0 9 2 9 0 9 1 0 2 9 7 13 3 9 10 0 9 2
20 1 14 3 0 9 10 9 13 11 2 11 9 9 1 9 0 9 1 11 2
18 9 11 3 13 2 16 1 9 12 4 9 1 11 3 3 3 13 2
32 11 2 11 1 9 10 9 3 13 2 16 7 1 9 9 0 9 1 0 9 4 13 10 0 9 1 3 0 9 16 3 2
11 11 11 7 13 13 9 10 9 11 11 2
19 1 9 16 0 13 1 9 11 11 9 1 11 9 11 11 2 11 2 2
27 13 2 16 9 13 9 1 11 2 11 3 0 7 16 13 3 9 0 9 2 15 13 7 1 0 9 2
2 0 9
35 1 9 1 9 11 2 11 7 11 1 11 1 0 9 9 0 0 9 7 1 0 9 12 9 13 3 1 11 9 0 9 11 1 11 2
26 9 11 1 11 11 11 1 15 13 2 16 0 9 1 0 9 13 9 0 9 2 7 7 9 0 2
42 1 9 0 9 0 1 11 15 1 9 9 0 9 13 1 0 9 9 9 11 11 11 13 2 9 7 9 7 13 10 9 2 16 0 4 15 3 13 1 11 2 2
3 9 1 9
26 0 9 2 15 13 3 0 9 1 9 11 7 11 1 11 2 4 13 13 0 9 0 1 0 11 2
24 12 0 9 1 9 3 12 9 7 12 0 9 3 1 9 13 9 1 0 9 11 5 11 2
15 1 9 4 9 13 13 1 9 14 1 0 9 1 11 2
16 9 0 7 0 9 1 12 10 9 13 11 1 12 9 9 2
21 1 9 0 9 13 13 9 9 3 1 12 12 2 15 15 13 3 1 0 9 2
30 0 9 1 0 9 0 3 15 3 13 9 0 0 9 2 7 2 1 9 9 11 11 2 13 13 9 1 9 11 2
9 9 13 9 1 0 2 2 0 9
5 11 2 11 2 2
11 0 0 9 0 9 1 11 13 0 9 2
27 3 15 13 9 9 0 9 1 11 9 2 11 11 2 1 9 13 1 9 11 1 9 12 0 0 9 2
19 9 13 0 9 2 15 15 1 11 13 1 9 1 9 1 9 9 9 2
9 13 15 15 13 14 1 12 9 2
14 11 11 3 13 2 10 7 15 9 9 15 9 13 2
13 11 13 12 9 0 9 1 10 9 1 0 9 2
20 1 0 9 10 7 0 9 4 13 2 16 15 1 15 0 13 1 10 9 2
17 0 9 9 1 11 15 12 0 9 9 9 13 3 12 2 9 2
24 13 0 9 7 9 3 13 9 7 13 9 7 14 1 9 13 0 9 1 0 9 0 9 2
8 9 13 2 9 9 13 9 9
3 2 9 2
5 13 9 0 4 13
9 11 3 13 1 0 9 11 11 11
9 15 3 3 13 2 15 15 13 2
10 2 10 9 13 0 2 16 4 13 2
42 13 10 9 1 9 2 1 15 9 13 2 7 15 13 2 10 9 1 0 9 10 9 2 0 9 7 9 0 0 9 2 1 9 1 9 7 9 2 9 2 9 2
27 0 9 13 1 9 2 16 13 3 0 9 2 7 3 1 15 13 13 7 15 3 13 7 1 15 13 2
33 9 1 10 9 15 3 13 2 7 3 15 3 13 15 2 16 4 16 9 13 1 10 0 9 2 1 15 4 13 16 9 2 2
17 10 9 15 1 9 13 1 9 2 15 16 0 13 0 15 9 2
27 7 13 15 3 9 9 2 0 9 13 7 10 9 11 11 2 16 15 13 9 13 9 1 9 9 9 2
5 15 13 10 9 2
30 2 9 9 15 13 3 2 16 15 1 9 13 2 1 0 7 3 2 16 4 13 2 16 4 15 9 13 1 12 2
11 13 15 15 2 16 13 9 9 10 9 2
23 13 0 9 0 9 2 0 0 9 0 2 7 7 9 3 0 2 15 15 3 13 13 2
6 3 4 15 15 13 2
13 11 11 13 0 9 2 13 3 1 3 0 9 2
29 3 15 13 2 16 13 2 14 9 9 2 4 13 3 15 13 2 14 3 13 9 2 7 13 3 10 0 9 2
9 13 10 10 9 2 7 13 15 2
25 13 3 1 9 10 9 2 13 15 7 2 16 0 9 13 3 15 0 2 15 4 15 13 13 2
22 7 7 16 4 15 15 13 1 15 10 13 2 3 14 3 1 9 0 9 0 9 2
28 13 15 9 2 15 3 1 0 9 13 9 11 7 3 13 2 16 1 9 9 4 13 13 9 1 9 11 2
26 13 3 9 2 16 13 2 14 15 13 15 13 2 3 15 15 15 4 3 13 1 0 9 9 2 2
4 9 9 0 13
8 1 11 14 2 1 11 0 9
21 9 0 9 1 10 9 11 13 7 13 9 9 0 9 0 9 1 11 2 11 2
44 9 9 2 9 0 9 11 1 11 1 11 2 11 2 13 3 12 9 1 9 12 9 1 11 2 12 1 11 2 11 7 12 1 9 12 9 1 0 9 11 1 0 9 2
14 9 1 9 12 9 4 1 0 9 13 1 0 9 2
29 0 9 1 9 12 9 1 11 2 11 7 11 13 1 9 1 9 7 4 15 1 9 9 1 0 9 9 13 2
7 13 15 0 9 1 11 2
22 9 1 0 9 1 0 9 4 13 0 9 13 1 9 1 9 9 1 0 9 9 2
17 15 4 13 13 0 9 11 2 15 9 13 15 9 9 1 9 2
18 9 9 4 7 13 0 9 11 2 11 1 0 9 3 1 9 12 2
42 11 11 1 9 0 9 9 0 9 11 2 2 0 9 1 11 2 11 15 1 9 9 13 3 2 16 4 14 10 9 13 9 7 9 7 10 9 4 13 9 9 2
37 15 15 13 2 16 13 1 3 0 9 7 13 15 15 0 16 9 9 1 0 9 13 9 9 2 16 10 9 1 0 9 1 11 13 0 2 2
26 0 9 0 9 0 9 11 2 11 11 11 13 2 16 10 0 9 13 14 3 2 16 4 13 9 2
17 2 9 7 9 13 9 1 0 9 7 13 10 9 1 0 9 2
12 3 9 9 1 9 0 9 1 11 4 13 2
13 0 9 1 11 2 11 7 11 4 13 9 3 2
13 9 7 9 15 1 9 13 2 2 13 11 11 2
19 1 15 13 0 9 13 3 2 16 9 2 15 13 2 13 13 1 9 2
24 9 2 16 13 0 13 15 1 0 9 2 15 4 3 9 13 2 3 1 9 0 9 13 2
15 2 9 13 13 9 9 1 9 2 3 13 3 9 9 2
12 10 0 9 15 13 1 0 9 9 0 9 2
41 16 4 10 9 13 7 13 2 13 4 3 1 0 0 9 9 0 9 2 7 9 1 9 2 2 13 15 11 11 2 9 9 0 0 9 11 1 11 1 11 2
18 9 9 0 9 0 9 1 11 2 11 13 9 12 0 9 1 11 2
18 1 15 13 1 0 9 2 3 9 4 13 3 2 7 13 0 9 2
23 9 12 0 9 1 0 9 7 1 9 9 1 11 15 3 13 3 1 0 16 0 9 2
38 2 16 4 13 2 16 0 9 11 13 9 0 9 13 2 13 4 15 15 3 13 1 2 2 13 15 11 11 1 9 0 9 0 9 1 0 11 2
14 9 0 9 7 13 9 0 9 2 15 3 9 13 2
23 1 0 9 4 9 13 13 0 12 9 2 16 0 1 9 4 13 13 9 14 12 9 2
8 9 10 9 13 1 0 11 2
10 14 1 9 9 13 3 0 9 0 2
21 9 9 0 11 3 13 9 0 12 9 1 9 2 15 13 9 11 3 1 9 2
29 2 1 0 9 13 13 1 9 9 9 2 15 4 0 9 9 13 2 2 13 15 1 15 9 0 11 11 11 2
8 2 13 13 9 1 9 2 2
17 9 9 3 13 1 9 9 0 9 2 3 7 13 0 0 9 2
5 13 9 0 4 13
6 3 4 3 3 13 2
26 2 9 1 15 2 16 7 0 9 1 9 9 0 9 2 13 4 13 2 16 4 15 3 15 13 2
25 16 4 13 2 10 9 4 13 2 16 4 15 13 1 9 2 16 4 1 9 1 9 13 9 2
22 16 4 4 13 2 13 4 9 1 9 2 15 13 0 15 9 2 3 1 9 2 2
14 1 9 1 0 9 13 9 10 9 1 9 3 3 2
28 16 3 1 9 12 15 13 0 13 15 9 11 2 15 15 13 3 0 2 1 9 12 13 9 9 9 13 2
5 3 15 15 13 2
5 2 9 13 3 2
24 12 1 15 13 3 0 9 2 16 9 13 9 2 7 10 9 1 0 9 13 7 10 9 2
23 7 10 9 13 13 3 7 15 2 16 3 10 9 13 9 1 0 9 3 1 10 9 2
23 15 13 3 3 2 15 4 15 13 1 9 2 16 4 13 13 7 13 1 12 9 2 2
16 10 0 9 1 9 13 11 2 15 15 3 13 1 10 9 2
32 0 9 13 10 9 7 15 2 16 9 1 9 2 0 9 2 4 0 1 9 11 11 1 9 12 7 1 10 0 9 11 2
9 13 4 13 10 9 1 10 9 2
30 2 1 9 9 11 4 13 15 0 2 3 2 3 4 15 3 13 9 1 10 2 16 4 1 10 9 13 3 13 2
27 13 4 15 1 3 0 9 7 13 4 2 16 10 10 9 1 15 4 13 13 14 7 14 0 0 9 2
15 16 4 13 15 0 1 0 9 9 11 2 13 0 9 2
17 9 11 13 3 3 9 13 3 10 0 9 2 15 15 13 13 2
20 0 9 13 2 16 15 9 9 11 11 13 3 0 2 16 9 9 9 11 2
16 7 15 13 3 10 9 2 15 4 3 13 1 10 0 9 2
27 13 3 9 7 9 2 16 4 13 10 9 7 13 15 10 0 9 13 9 0 9 2 13 15 0 2 2
17 11 11 3 13 2 16 4 1 10 0 9 3 13 10 0 9 2
18 7 7 3 0 0 7 0 9 13 10 9 16 9 1 10 0 9 2
10 3 13 1 10 10 9 1 9 9 2
29 2 9 2 3 9 11 7 11 13 2 16 4 4 13 9 2 13 0 7 0 2 13 1 15 3 14 0 9 2
31 1 10 9 4 13 9 1 15 2 15 13 0 2 15 13 9 7 15 13 0 0 2 0 7 0 9 1 10 0 9 2
12 16 15 9 11 13 1 15 2 13 10 9 2
13 9 15 1 15 3 13 2 16 15 13 10 9 2
16 15 4 1 0 9 13 13 1 10 0 9 7 1 15 13 2
7 13 4 3 13 0 9 2
9 13 15 2 16 15 13 10 9 2
13 13 15 3 4 13 13 9 2 15 13 10 9 2
9 1 15 4 7 10 9 13 2 2
23 1 0 9 10 0 9 3 13 1 9 0 9 2 15 4 15 15 3 3 7 3 13 2
12 13 4 1 15 1 0 9 3 9 10 9 2
17 2 9 4 4 13 9 1 9 2 3 4 1 15 3 3 13 2
9 3 15 15 13 13 1 9 3 2
14 15 7 3 7 10 9 13 3 13 2 7 1 15 2
30 11 3 2 16 4 13 0 9 2 13 1 11 0 9 2 16 0 2 15 14 13 15 2 15 0 0 9 3 13 2
27 13 15 13 2 16 4 15 1 9 13 13 11 7 0 9 0 9 1 15 2 16 4 13 1 15 0 2
10 7 1 15 4 13 1 9 13 11 2
40 7 4 13 2 16 13 13 0 9 2 15 13 3 4 13 2 16 15 15 3 0 0 9 13 2 7 4 13 2 16 13 9 2 1 15 3 16 3 13 2
10 13 4 3 1 0 9 7 0 9 2
10 13 2 10 9 4 10 9 13 2 2
11 3 1 10 9 13 9 9 9 0 9 2
7 13 1 15 9 0 9 2
7 2 13 1 9 0 9 2
15 10 9 13 3 0 9 2 7 15 10 9 13 0 9 2
15 9 13 1 0 9 3 13 1 10 9 7 3 7 3 2
18 13 1 10 9 2 15 13 1 9 1 0 9 7 10 9 13 4 2
18 1 9 3 0 4 3 13 0 13 9 10 9 1 0 9 1 9 2
19 15 15 7 13 2 16 13 3 10 9 15 1 0 9 13 1 10 9 2
75 11 13 3 2 3 2 2 10 0 9 3 13 3 3 2 16 9 9 3 13 1 15 9 2 15 4 13 10 9 7 15 4 15 13 3 10 9 2 15 4 13 10 0 15 9 2 13 2 14 7 9 0 2 0 9 13 9 9 1 11 2 16 0 9 2 13 3 9 9 2 13 13 15 2 2
22 16 13 1 9 1 12 9 2 13 0 3 1 9 0 9 2 10 9 15 14 13 2
41 13 1 0 9 12 9 2 16 4 9 13 3 2 1 9 9 2 16 4 12 0 9 13 9 0 7 16 4 10 0 9 13 13 9 2 0 9 7 0 9 2
26 11 13 9 1 9 2 11 13 13 10 9 1 9 7 13 15 1 11 13 2 3 15 15 3 13 2
27 13 1 15 0 9 1 9 0 9 15 13 3 3 0 2 9 1 9 15 3 13 3 13 3 0 9 2
37 1 0 9 7 13 13 2 16 4 15 11 3 13 9 2 16 4 13 14 1 9 0 7 13 9 0 10 9 14 1 9 2 3 9 3 13 2
11 13 2 14 15 3 2 13 4 15 15 2
27 7 15 13 2 9 11 2 3 11 2 15 3 13 1 9 9 2 15 13 3 1 11 7 3 0 2 2
14 2 9 4 13 9 9 0 9 2 2 2 2 2 2
29 2 16 4 15 3 13 2 0 9 4 15 13 16 9 7 13 4 15 15 2 2 13 4 1 9 1 0 9 2
8 13 3 9 1 9 0 9 2
15 2 15 3 15 10 9 13 13 2 16 15 1 9 13 2
14 3 4 0 9 10 9 13 2 15 15 13 14 9 2
25 7 16 13 2 16 9 13 3 3 0 2 3 15 13 2 16 15 0 9 4 13 1 9 0 2
10 13 2 14 15 3 2 15 3 2 2
19 16 4 1 9 13 1 11 11 2 13 4 9 2 0 9 0 9 2 2
24 13 15 2 16 1 9 0 0 9 7 9 1 10 0 9 13 3 0 13 0 9 0 9 2
26 2 0 9 7 9 13 3 9 1 10 9 7 9 2 7 3 1 15 2 16 4 15 15 13 2 2
36 14 2 15 13 9 2 7 1 9 10 9 3 1 0 9 2 13 9 1 11 7 0 9 1 9 1 9 12 2 13 3 0 9 7 9 2
7 13 3 15 10 0 9 2
18 2 3 2 16 10 9 1 9 1 9 0 9 13 3 1 10 9 2
17 7 7 15 13 0 13 7 3 7 3 13 1 0 0 0 9 2
15 13 9 2 16 9 2 0 9 2 13 7 0 9 2 2
18 15 1 15 2 10 0 9 4 15 3 13 13 9 13 0 9 9 2
22 2 9 9 2 9 2 9 7 3 9 13 3 0 2 16 13 3 0 1 15 13 2
8 7 4 3 3 13 9 9 2
28 12 1 9 9 2 3 15 2 13 2 16 13 1 9 3 9 0 2 15 13 3 16 1 9 0 9 2 2
21 0 0 9 4 1 15 13 13 0 0 9 2 15 4 13 9 2 14 9 9 2
18 13 15 3 1 10 9 1 11 11 2 15 9 13 9 10 0 9 2
17 7 11 3 13 2 16 14 1 0 9 11 13 0 9 0 9 2
6 13 3 1 0 9 2
51 2 11 13 3 0 2 10 9 9 2 15 13 1 0 9 2 15 13 2 9 13 0 7 15 4 3 3 13 2 16 13 9 15 13 1 15 0 9 7 15 9 0 9 7 13 10 0 9 3 3 2
10 9 0 9 13 1 15 10 0 9 2
44 3 13 9 2 15 13 10 0 9 2 0 9 1 9 2 13 13 9 7 3 13 2 7 13 15 15 0 13 1 10 9 9 1 9 7 13 15 15 13 2 13 15 0 2
30 9 9 13 9 0 9 2 9 2 9 0 9 7 9 0 9 2 13 15 15 15 4 13 13 15 9 0 9 2 2
26 13 15 13 2 16 1 11 13 9 15 2 16 10 0 9 4 13 7 13 9 15 13 7 9 13 2
14 2 13 4 2 16 0 0 9 13 0 7 0 9 2
23 3 13 9 13 9 0 0 9 9 0 9 7 13 9 2 3 15 3 13 0 9 13 2
25 3 13 3 0 0 9 13 1 0 9 1 2 9 2 2 2 9 2 7 2 0 9 2 2 2
24 13 9 2 16 15 15 3 9 11 2 7 7 0 9 13 13 2 16 4 13 1 10 9 2
11 13 3 0 9 13 1 0 9 0 9 2
16 2 7 1 15 13 3 0 9 7 3 9 1 0 9 0 2
38 13 2 14 13 9 12 13 9 10 0 9 2 3 4 15 13 13 15 2 15 13 3 2 9 0 2 2 10 0 9 2 15 15 3 1 9 13 2
12 10 9 4 13 13 3 14 9 0 7 0 2
19 13 15 2 7 13 4 15 13 2 9 2 15 13 3 0 1 15 12 2
28 7 3 15 13 13 10 9 1 15 2 16 4 13 7 13 15 1 0 0 0 9 2 3 1 9 10 9 2
41 1 10 9 7 2 3 15 0 9 3 3 13 7 3 13 0 9 2 3 4 10 0 9 3 13 2 14 13 2 15 15 13 2 16 15 13 3 0 9 13 2
10 15 4 14 13 14 1 0 0 9 2
34 13 15 15 2 16 3 3 13 9 3 0 2 0 1 9 3 3 0 0 0 7 0 9 2 3 9 3 0 1 10 0 0 9 2
5 15 13 9 0 2
31 16 13 1 15 3 2 13 9 1 10 9 13 7 15 13 2 7 13 15 7 2 16 4 10 9 13 1 10 0 9 2
11 3 4 3 10 0 0 9 3 3 13 2
21 3 13 15 2 16 4 10 9 1 10 0 9 13 2 16 13 9 3 3 0 2
15 9 10 9 1 15 7 9 0 9 15 3 3 13 2 2
15 9 0 9 15 13 1 0 9 1 0 0 9 11 11 2
29 3 15 15 2 15 13 9 3 1 3 0 9 9 2 13 1 9 2 15 1 10 9 13 1 9 3 0 9 2
13 2 13 2 16 3 7 15 13 3 3 13 2 2
37 16 3 13 1 11 11 2 1 9 15 13 9 1 15 2 16 9 13 1 9 12 0 9 13 0 9 9 11 1 3 3 0 9 9 0 9 2
5 13 10 9 0 2
16 2 16 15 13 0 9 11 7 11 2 13 15 1 0 9 2
44 13 15 1 15 0 2 1 0 9 2 7 15 15 13 2 16 1 10 9 9 15 9 11 7 11 3 13 2 16 4 1 11 11 13 1 9 2 16 4 13 9 0 9 2
45 13 15 1 9 2 3 9 9 13 1 0 13 9 1 9 7 13 15 1 0 0 9 2 7 15 15 13 2 16 10 9 4 13 3 13 3 9 3 0 2 15 13 11 11 2
8 9 13 7 7 0 0 9 2
9 13 3 7 1 9 7 1 9 2
35 15 1 15 1 11 11 3 14 13 2 13 4 3 1 15 2 7 13 4 1 15 1 15 1 9 0 9 2 14 3 10 2 9 2 2
22 1 9 9 15 13 2 16 13 3 2 16 11 11 13 9 9 7 11 11 9 9 2
24 7 1 0 9 15 3 13 0 9 2 3 7 15 2 15 15 1 9 13 16 3 0 2 2
6 13 15 3 1 9 2
16 13 14 0 13 15 15 2 16 4 13 13 9 0 0 9 2
15 13 15 7 13 2 1 10 9 4 3 0 9 13 13 2
8 2 9 4 13 3 2 13 2
18 3 4 13 13 9 2 16 4 1 9 10 9 13 3 0 0 9 2
44 13 15 2 16 4 13 10 9 3 13 2 16 4 3 13 14 1 0 9 9 7 14 1 12 9 7 16 4 15 0 13 1 9 7 14 3 2 16 4 3 10 9 13 2
29 3 7 1 0 9 4 13 0 2 16 4 13 15 2 16 15 13 0 13 9 2 15 15 13 3 1 0 9 2
60 3 4 13 13 9 2 15 9 13 0 0 9 7 15 13 14 1 15 2 16 4 1 9 1 9 13 9 2 13 9 1 9 2 13 0 9 1 9 7 13 0 9 9 2 9 2 1 15 4 15 13 13 1 0 9 3 3 1 9 2
37 15 4 10 9 3 1 9 13 2 7 15 13 3 0 9 2 0 2 16 3 13 2 13 1 15 2 16 13 15 0 13 1 0 9 7 9 2
11 13 14 3 9 0 4 14 3 13 2 2
17 7 0 9 2 3 15 4 3 13 2 16 13 2 10 9 2 2
13 13 1 9 13 9 9 7 13 10 9 7 9 2
10 2 13 4 15 15 2 7 14 3 2
9 13 4 15 3 2 7 3 3 2
29 13 15 9 1 0 9 2 15 4 15 13 14 1 12 9 2 16 4 15 3 3 13 1 15 0 7 0 9 2
8 2 10 0 9 13 3 2 2
31 16 4 4 1 10 0 9 1 11 2 3 15 15 3 14 2 13 2 2 13 2 15 1 15 13 2 3 4 15 13 2
5 13 15 10 9 2
28 13 4 3 1 10 9 7 9 11 11 2 15 13 10 10 0 9 3 2 7 1 9 9 2 15 15 13 2
29 13 1 15 9 2 16 13 10 0 9 1 9 9 7 9 2 15 1 9 0 9 2 1 15 13 13 10 9 2
22 7 9 1 10 9 13 1 10 9 7 13 15 15 1 15 7 15 15 1 15 13 2
29 1 15 15 7 13 2 13 1 9 10 0 9 7 15 13 3 0 9 1 9 1 0 9 2 15 9 15 13 2
10 3 2 16 13 10 9 2 16 0 2
7 13 7 0 2 7 0 2
64 16 4 15 3 13 1 15 2 16 2 13 10 9 2 2 13 4 1 9 1 0 9 13 2 3 15 1 0 9 13 1 0 9 2 13 15 2 9 9 15 13 7 13 2 3 15 1 0 9 7 0 9 3 13 7 3 0 9 3 13 7 3 13 2
5 15 15 4 13 2
53 13 3 7 10 0 9 1 15 2 3 4 15 13 3 1 10 9 13 2 3 0 9 3 13 2 3 0 9 13 2 3 13 1 0 9 2 13 10 9 1 0 9 2 1 9 0 9 7 1 9 0 9 2
13 13 3 2 3 1 10 9 3 13 9 7 9 2
55 3 7 0 2 16 0 9 1 9 7 9 0 0 9 2 13 15 0 2 9 1 0 9 0 9 2 1 15 4 10 9 13 13 2 1 9 7 9 0 9 2 15 4 15 13 13 2 1 9 2 15 4 13 13 2
42 15 15 3 13 2 7 13 4 9 2 16 4 15 1 15 13 2 7 13 3 1 10 0 7 15 0 0 9 1 9 9 2 3 4 15 13 13 1 0 0 9 2
48 13 2 10 2 9 2 13 15 0 2 16 9 1 9 2 15 4 0 3 13 2 1 0 0 9 2 15 1 10 9 13 2 7 1 9 2 3 1 10 0 9 10 9 7 9 13 2 2
4 9 2 11 2
2 11 11
1 9
2 9 12
5 9 1 12 1 12
5 9 1 12 1 12
1 11
1 3
3 9 13 11
29 11 9 2 9 9 11 2 15 13 2 16 3 0 9 9 9 4 13 9 9 0 9 2 3 9 12 0 9 2
11 13 15 1 0 9 11 1 9 1 11 2
21 9 1 11 2 11 15 13 7 13 4 14 3 1 9 9 9 2 15 9 13 2
30 9 10 9 7 0 9 13 1 0 9 0 1 11 7 13 2 16 1 10 9 13 3 13 1 0 9 15 9 13 2
25 9 9 0 12 2 9 1 12 9 7 12 9 11 13 3 0 0 9 1 9 1 9 9 9 2
19 9 15 13 12 9 0 9 2 15 13 12 9 9 7 12 9 0 9 2
26 9 9 0 12 9 9 0 9 0 0 9 0 9 1 11 13 3 9 9 11 11 9 11 11 11 2
28 1 0 9 0 9 1 0 13 9 11 1 9 0 7 9 0 1 15 2 16 11 4 13 0 9 0 9 2
20 0 9 13 1 9 11 11 11 14 0 9 11 2 7 3 7 10 0 9 2
5 9 11 15 3 13
2 11 2
5 9 11 15 3 13
2 11 2
28 9 0 9 11 11 1 9 0 0 9 11 11 13 9 2 16 4 15 11 13 3 13 1 9 1 0 9 2
25 11 2 12 2 3 13 2 16 15 1 9 13 9 2 16 15 9 1 0 9 1 0 9 13 2
25 0 9 11 13 11 2 11 2 15 13 3 0 9 0 9 2 16 0 9 15 13 1 0 9 2
16 12 9 15 1 15 13 2 16 1 9 9 4 1 9 13 2
19 14 1 12 9 10 9 13 1 11 1 11 0 9 11 11 1 10 0 9
10 0 9 1 9 9 0 9 11 7 11
2 11 2
15 0 0 9 2 11 2 15 0 9 13 1 11 0 9 2
6 13 15 3 9 11 2
17 0 9 15 1 9 1 9 13 1 9 11 1 11 9 0 9 2
37 9 1 0 9 1 0 9 2 0 9 11 11 2 9 11 13 2 16 15 11 7 0 9 13 0 9 1 9 1 9 9 2 0 9 7 9 2
10 0 9 1 9 1 11 15 4 13 9
12 1 0 0 9 15 1 0 0 9 13 9 2
27 1 0 9 4 13 12 9 9 2 14 12 9 2 3 7 1 0 9 12 9 9 2 12 9 2 3 2
19 9 4 13 2 16 10 9 13 14 12 9 9 0 1 9 1 0 9 2
27 1 9 1 15 15 1 9 9 13 13 9 1 9 9 1 0 9 2 1 15 4 15 9 3 13 9 2
8 13 11 9 11 9 1 9 2
2 11 2
14 11 4 13 1 11 1 9 15 0 9 9 1 9 2
9 13 15 3 0 9 9 11 11 2
14 13 1 3 0 9 0 9 2 15 4 13 9 12 2
24 11 2 11 13 2 2 13 15 2 16 4 13 13 9 1 11 3 1 9 2 7 13 9 2
17 13 9 2 16 4 15 15 13 13 9 2 7 13 15 13 2 2
17 9 1 0 9 0 9 1 0 9 11 11 3 3 13 1 9 2
20 1 0 9 1 9 0 9 3 7 0 9 13 9 0 9 0 1 10 9 2
15 2 13 9 11 11 13 1 0 2 0 9 9 2 12 2
9 9 11 11 13 1 0 2 0 9
2 11 2
17 0 9 9 11 11 13 3 1 9 0 2 0 9 1 0 9 2
41 2 13 2 16 13 10 9 2 7 13 2 16 10 9 13 0 2 2 13 9 0 9 1 9 1 9 2 15 13 9 1 9 1 9 11 11 7 9 11 11 2
29 2 13 15 2 16 3 13 9 2 16 4 15 13 9 11 1 15 9 1 9 11 1 15 9 2 2 13 11 2
3 0 11 2
19 11 4 13 1 2 0 9 2 1 11 2 13 3 0 9 9 11 11 2
30 2 13 0 13 1 0 9 1 0 9 1 0 9 2 2 13 9 9 11 3 1 9 9 1 10 0 9 11 11 2
6 2 10 9 13 0 2
15 13 15 13 11 2 15 15 13 2 2 13 11 2 11 2
2 11 2
2 9 2
11 0 0 9 3 13 9 0 11 11 9 2
5 13 15 0 9 2
2 11 2
2 9 2
14 9 0 9 11 11 15 3 3 13 12 2 0 9 2
9 9 1 10 9 13 9 11 11 2
10 3 15 13 2 16 4 13 0 9 2
4 11 1 11 2
18 1 9 9 0 9 11 11 13 3 3 1 11 9 0 9 11 11 2
4 9 13 0 9
2 11 2
8 9 13 0 9 11 2 11 2
18 9 1 3 0 9 2 12 4 13 1 9 0 0 9 1 0 11 2
8 13 15 3 9 11 2 11 2
16 9 13 1 9 9 2 1 15 9 9 1 9 1 9 13 2
20 9 1 9 1 0 9 13 1 9 2 16 9 15 13 9 3 13 1 9 2
14 9 10 9 15 1 0 9 13 1 10 9 12 9 2
18 1 3 0 9 0 9 13 9 2 16 9 3 13 2 15 3 13 2
26 16 9 13 2 3 0 9 2 15 1 15 13 2 4 13 0 9 1 15 0 3 2 13 0 9 2
9 11 13 1 11 2 9 0 7 0
1 9
9 11 13 1 11 2 9 0 7 0
17 11 2 3 10 0 0 2 0 9 2 4 13 1 9 0 9 2
20 13 15 3 7 3 3 7 3 9 2 15 13 13 0 9 1 9 10 9 2
40 11 13 1 9 1 2 0 9 2 2 16 4 15 7 3 13 1 9 2 7 14 1 10 0 9 0 1 9 2 3 1 9 9 13 10 10 9 3 0 2
35 16 9 0 9 0 0 9 1 9 13 2 16 3 3 15 14 13 7 1 0 0 9 2 11 15 4 13 3 13 9 1 9 1 11 2
15 3 1 0 9 0 9 13 2 16 15 3 3 15 13 2
25 3 0 7 0 9 1 15 2 7 3 1 0 0 7 0 9 2 13 2 13 7 13 0 9 2
31 0 9 9 1 9 0 9 3 13 4 3 13 3 3 3 14 3 2 16 11 13 14 9 1 0 0 0 7 0 9 2
24 13 13 3 16 9 2 9 7 15 9 0 9 9 2 16 13 3 3 1 9 0 9 9 2
25 11 13 3 3 3 1 9 0 9 2 3 3 3 2 16 11 13 1 0 9 1 11 7 11 2
31 16 13 3 3 9 2 10 10 9 13 2 7 11 13 3 3 13 10 9 1 2 9 2 0 9 2 7 3 0 9 2
9 3 3 3 13 16 13 0 9 2
7 7 16 1 3 0 9 2
18 9 11 1 11 15 13 9 2 9 2 9 2 7 13 15 7 9 2
23 13 14 0 9 0 2 15 13 10 9 13 1 9 0 9 2 9 9 7 9 1 11 2
4 0 9 1 11
2 11 2
48 0 9 1 11 0 11 2 9 1 10 0 9 11 0 11 13 3 0 9 9 11 11 1 0 11 9 9 1 9 9 2 15 13 3 0 1 9 11 1 9 1 9 0 9 1 11 11 2
27 2 0 9 4 13 7 10 9 9 11 7 7 9 3 13 9 12 0 9 1 11 2 2 13 9 11 2
9 9 1 11 13 4 13 9 11 11
2 11 2
31 11 13 0 9 11 11 11 9 2 1 15 15 13 2 16 4 13 0 7 0 9 1 3 0 0 9 1 9 12 9 9
14 13 15 1 9 3 1 11 9 0 9 0 11 11 2
36 1 0 9 1 9 11 1 11 2 3 15 13 0 9 0 0 9 7 0 9 2 11 13 2 16 1 11 13 0 9 2 15 13 3 9 2
4 9 1 9 13
7 9 9 7 11 15 3 13
2 11 2
27 0 9 7 0 0 9 2 11 2 15 3 13 13 9 0 9 0 9 9 1 11 1 9 11 11 11 2
46 1 0 9 4 0 9 1 0 9 11 11 11 7 9 0 9 11 11 13 7 1 9 2 16 4 13 3 0 9 13 3 1 0 0 9 11 7 11 2 15 9 11 13 0 9 2
21 9 9 13 0 9 1 9 1 9 1 11 1 11 2 15 15 13 9 9 0 9
22 9 1 9 1 0 2 11 15 13 3 1 9 2 16 0 11 13 0 9 0 1 9
5 9 2 11 2 11
12 9 1 11 13 0 9 1 2 0 9 2 11
6 10 9 13 1 0 9
2 11 2
29 11 2 11 2 11 2 11 7 11 2 15 13 9 9 7 9 2 15 15 3 13 1 2 0 9 2 1 11 2
29 1 0 9 0 9 13 12 9 1 11 2 9 1 0 9 13 12 2 11 12 2 11 12 7 9 1 11 12 2
32 1 9 11 0 11 13 0 9 1 11 13 9 1 0 9 2 7 3 4 15 3 13 0 9 0 9 7 3 13 15 13 2
39 9 9 13 3 0 2 9 9 7 3 9 12 2 12 9 9 2 3 12 2 12 12 9 2 1 10 9 7 1 9 9 7 2 9 1 0 9 2 2
6 2 9 9 2 1 9
8 13 15 9 11 2 11 2 11
2 11 2
15 9 0 9 11 2 11 2 11 4 3 3 13 1 11 2
37 12 9 0 0 9 0 1 11 7 11 2 15 1 11 13 1 11 2 3 13 9 10 9 1 3 12 0 0 9 1 9 1 0 1 0 9 2
15 9 9 13 3 1 0 9 12 0 9 7 10 0 9 2
6 9 9 13 12 9 2
19 0 2 7 16 0 9 1 9 11 7 11 13 3 1 9 12 11 0 2
12 7 3 0 9 13 7 9 2 9 9 2 2
2 0 2
4 7 3 0 9
4 13 15 9 9
2 11 2
2 9 2
4 13 15 9 9
2 11 2
32 1 9 7 9 2 15 1 9 7 1 9 1 9 13 0 11 2 7 7 11 7 11 2 13 1 9 7 4 13 9 9 2
21 1 3 0 9 11 2 11 2 13 1 0 9 12 9 7 12 15 13 3 0 2
13 9 9 3 13 9 7 9 2 4 13 10 9 2
7 9 13 9 1 9 9 2
2 9 9
2 11 11
2 9 9
15 1 12 9 9 15 13 1 0 11 1 9 0 0 9 2
10 0 9 7 14 13 1 9 0 9 2
7 3 15 13 9 0 9 2
16 1 9 1 0 9 13 1 0 9 9 1 0 11 7 11 2
3 3 1 9
20 11 11 15 13 2 16 13 13 9 9 7 3 4 15 15 1 9 9 13 2
8 3 15 16 9 0 9 13 2
33 0 9 9 9 13 0 2 13 1 0 9 7 1 9 2 0 9 1 9 11 7 11 13 1 9 0 0 9 9 1 9 9 2
17 1 15 15 1 0 0 9 0 9 9 1 0 11 13 9 9 2
39 0 9 13 1 2 9 1 9 2 7 1 15 2 16 15 9 2 11 13 2 16 0 9 4 13 1 0 9 7 3 15 13 10 9 1 9 2 2 2
28 13 13 7 9 0 9 11 2 15 0 9 13 13 9 1 9 9 7 1 9 9 11 15 1 10 9 13 2
19 16 3 13 9 9 9 1 9 0 2 9 13 2 16 1 15 9 13 2
27 13 15 3 13 2 16 15 15 9 13 3 3 2 16 4 15 9 9 13 13 9 1 12 9 0 9 2
10 0 9 0 9 9 9 11 11 13 0
25 2 9 0 9 13 1 9 0 9 13 1 0 0 9 2 2 13 9 9 0 9 9 11 11 2
17 1 9 9 15 13 9 2 7 0 0 9 15 13 0 0 9 2
37 9 9 0 9 0 9 2 11 2 11 11 15 7 13 2 16 9 9 13 9 9 0 9 9 0 9 15 2 16 13 9 0 9 1 12 9 2
16 15 3 0 9 13 2 13 1 9 13 1 9 10 9 3 2
21 2 0 9 13 3 13 2 13 1 9 2 16 9 13 3 2 2 13 11 11 2
21 2 16 13 3 0 2 16 1 9 11 13 0 9 0 9 11 10 9 13 2 2
15 2 0 9 13 13 3 1 0 9 2 9 2 9 2 2
15 9 0 9 13 7 0 9 0 9 2 15 13 9 9 2
30 15 3 13 7 13 9 0 9 2 13 3 2 13 0 9 2 2 3 13 1 9 9 2 12 2 12 9 1 9 2
29 9 9 0 9 9 11 11 2 2 13 9 9 13 2 13 3 1 9 15 2 10 9 15 1 15 3 13 2 2
3 9 2 11
4 9 2 11 3
13 9 0 9 4 13 1 0 2 0 7 0 9 2
15 13 1 0 9 0 9 2 15 4 13 9 1 10 9 2
12 4 13 9 1 0 0 9 7 9 0 9 2
7 13 1 9 12 0 9 2
3 2 11 2
2 0 11
31 0 9 0 0 9 11 1 9 0 9 15 1 0 12 9 0 9 13 1 0 9 12 1 12 9 2 1 12 9 9 2
10 1 15 1 0 11 13 12 9 9 2
23 0 9 9 1 0 9 7 1 11 13 9 11 0 9 10 9 1 11 2 11 7 11 2
23 3 13 0 9 11 2 13 11 3 13 10 9 1 12 9 9 11 7 11 1 0 12 2
28 11 13 1 9 12 10 9 1 11 1 0 12 9 1 12 9 7 1 0 12 9 13 13 14 12 9 9 2
13 0 9 9 4 15 3 13 13 1 12 9 3 2
20 9 13 2 16 16 3 13 0 9 9 12 9 9 2 3 3 4 13 9 2
15 3 13 1 9 12 9 7 1 11 13 12 11 7 11 2
5 0 9 13 1 9
17 2 9 9 7 13 1 0 9 12 9 9 2 2 13 11 11 2
10 0 9 9 13 0 9 9 1 9 2
11 0 9 13 7 1 9 7 9 1 9 2
22 7 2 3 13 9 11 2 9 11 13 9 15 0 9 0 9 1 3 12 9 9 2
23 9 11 11 13 3 9 9 1 0 9 2 15 4 13 1 9 9 1 9 9 7 9 2
26 2 0 9 13 9 9 1 9 1 9 7 1 9 2 2 13 1 0 9 9 11 11 2 11 2 2
12 13 2 16 1 10 9 13 0 9 0 9 2
19 0 0 9 13 1 9 9 9 11 1 9 0 9 11 1 0 9 12 2
26 13 9 11 2 16 4 3 13 9 2 15 13 9 1 0 9 0 9 2 3 1 9 9 1 9 2
16 9 13 3 1 0 9 13 9 1 9 0 9 1 0 9 2
12 3 3 13 9 0 9 0 9 11 11 11 2
32 9 13 7 0 0 9 13 13 2 3 2 7 3 3 3 2 2 16 0 9 11 11 13 2 16 15 9 1 15 3 13 2
23 0 0 9 3 13 2 16 1 9 13 0 9 0 15 1 0 9 2 9 1 12 9 2
5 13 15 0 9 2
4 0 9 1 9
5 9 10 9 3 13
17 0 9 0 9 11 2 11 4 3 13 2 16 9 13 1 9 2
17 11 13 9 9 2 15 13 9 0 9 1 11 2 11 7 11 2
46 2 10 9 13 3 0 9 9 2 16 9 13 1 1 0 9 3 0 2 2 13 9 9 0 0 9 9 0 9 11 11 7 13 2 2 13 4 2 16 4 13 9 7 0 9 2
20 0 9 2 15 15 9 11 13 2 13 3 13 7 13 14 1 0 9 2 2
17 1 9 11 9 13 9 2 16 4 1 15 9 0 9 13 11 2
14 9 9 13 2 16 4 15 13 0 9 9 1 11 2
19 9 11 3 13 3 2 16 13 9 1 15 2 16 4 1 11 15 13 2
18 13 15 7 1 9 2 16 1 9 0 9 13 9 1 0 9 11 2
24 9 15 3 13 14 1 12 9 2 16 15 1 10 9 13 9 11 1 11 7 0 0 9 2
9 2 3 0 0 9 13 1 9 2
26 0 9 13 13 1 9 9 2 7 13 2 16 13 1 9 2 3 1 9 9 2 2 13 9 11 2
4 0 9 11 12
8 9 1 11 13 9 9 9 12
14 9 0 9 11 12 13 4 13 1 12 2 9 12 2
20 9 0 9 11 11 11 11 13 2 16 1 0 9 4 13 14 12 9 9 2
17 2 13 15 4 3 3 2 16 15 4 13 2 2 13 9 11 2
7 3 9 13 12 0 9 2
12 13 15 12 2 9 13 9 1 0 9 2 2
11 0 9 13 12 9 2 13 15 4 12 2
13 0 9 2 9 11 12 2 12 2 13 12 9 2
15 9 0 9 13 3 14 12 9 9 1 0 9 11 12 2
11 0 9 15 1 9 11 13 1 12 9 2
7 0 9 13 9 0 9 2
8 15 13 3 12 9 0 9 2
6 1 9 13 12 9 2
47 16 0 9 0 11 12 2 9 0 0 9 0 1 0 0 9 2 13 3 9 7 9 9 13 1 9 0 9 2 1 9 2 3 3 13 9 1 0 9 2 13 9 0 9 9 13 2
40 1 9 12 4 13 12 9 2 12 9 9 2 2 1 9 12 13 9 12 9 2 12 9 0 9 2 2 1 9 12 4 13 12 9 2 12 9 9 2 2
20 1 9 12 3 13 9 1 9 14 12 9 7 1 9 3 3 3 12 9 2
10 0 9 9 13 1 9 0 0 9 2
32 11 7 1 0 9 13 9 3 1 11 2 11 2 0 3 0 9 2 0 11 2 11 2 0 9 2 11 2 11 7 11 2
12 2 13 15 13 3 3 2 2 13 9 11 2
11 2 1 0 9 7 9 13 4 3 13 2
16 1 0 9 4 13 0 0 9 2 7 15 3 13 3 13 2
13 1 12 2 9 4 13 9 1 0 9 7 9 2
8 4 13 3 7 0 9 2 2
8 9 1 9 1 0 9 13 2
16 1 9 11 15 7 11 13 2 16 1 10 9 3 4 13 2
6 3 0 9 1 9 9
24 9 14 1 9 12 9 9 13 15 9 2 15 15 3 13 9 7 4 1 9 13 1 9 2
24 9 12 2 9 2 1 9 0 7 0 2 7 12 2 9 13 3 9 15 3 0 0 9 2
17 3 13 1 9 9 15 0 9 1 9 13 0 9 1 0 9 2
43 1 0 9 13 1 9 2 1 10 9 2 13 3 9 3 0 0 9 2 3 15 0 9 2 2 16 1 9 9 1 0 9 13 3 9 1 9 13 1 9 0 9 2
9 7 10 9 3 13 13 0 9 2
11 2 1 0 0 9 13 3 1 0 9 2
20 1 11 13 1 0 9 13 14 12 12 0 9 2 16 9 13 13 12 12 2
18 7 3 2 16 4 15 9 13 3 1 9 2 13 1 3 0 9 2
45 3 13 9 0 9 9 2 3 0 9 4 13 3 2 7 1 9 2 7 1 10 9 13 13 7 1 9 2 2 13 15 11 11 2 9 0 9 0 9 0 2 9 2 11 2
17 3 0 9 1 0 9 13 13 3 3 3 0 9 12 0 9 2
9 15 13 0 9 0 9 1 9 2
45 3 16 12 9 9 7 13 1 3 9 9 2 7 16 0 9 4 13 1 0 9 3 2 7 1 0 9 15 3 3 13 12 7 12 9 2 2 10 9 13 1 9 15 9 2
7 9 7 13 9 13 3 2
15 2 10 9 13 7 0 9 2 1 15 15 13 9 13 2
18 3 3 13 1 15 9 0 9 7 1 9 9 15 15 3 13 13 2
22 13 1 15 2 16 4 0 9 10 9 13 7 9 13 2 1 9 0 9 7 13 2
35 9 4 15 13 13 1 9 1 0 9 7 3 13 9 2 16 15 3 3 13 13 2 1 0 4 15 15 13 9 2 2 13 11 11 2
3 9 1 9
5 11 2 11 2 2
9 9 9 11 13 9 0 0 9 2
40 9 9 11 11 13 3 1 10 9 2 16 11 11 13 2 1 9 1 0 9 2 3 1 0 9 1 0 9 0 9 3 1 9 11 7 9 0 0 9 2
28 3 3 11 2 11 13 2 0 0 9 15 3 13 2 10 9 15 4 13 1 9 9 7 9 0 9 9 2
10 0 13 3 9 1 9 0 2 9 2
20 2 0 9 0 9 9 4 1 0 9 13 1 0 7 0 0 9 0 9 2
20 1 10 9 4 13 1 11 1 9 9 0 0 9 2 2 13 11 2 11 2
14 0 7 0 9 4 15 1 15 13 13 1 0 9 2
12 9 0 2 9 15 4 13 1 9 10 9 2
18 0 9 9 9 11 11 13 2 16 0 9 0 9 13 3 12 9 2
16 3 3 2 3 13 2 11 11 13 1 9 13 0 0 9 2
3 11 1 11
5 11 2 11 2 2
27 9 0 9 11 11 2 11 2 13 1 0 0 9 11 9 11 11 11 1 0 9 0 9 1 0 9 2
22 10 9 3 1 0 9 11 2 11 13 9 2 3 13 11 13 10 9 1 0 9 2
28 11 11 3 13 2 16 12 7 12 9 0 9 1 0 9 3 13 1 11 2 16 13 0 1 9 0 9 2
2 9 11
17 9 11 7 10 9 1 0 9 13 1 0 9 7 1 9 9 2
8 13 1 9 2 3 1 11 2
32 2 1 9 9 12 4 13 0 9 2 2 13 9 9 11 11 2 2 7 3 4 3 13 7 3 15 13 2 16 3 13 2
17 13 4 15 15 2 14 16 15 9 3 13 2 15 3 13 2 2
5 3 15 11 13 2
13 3 13 1 10 9 11 10 0 9 9 1 15 2
6 1 0 13 3 0 2
22 9 13 3 3 0 2 7 0 9 7 9 1 9 0 9 9 15 13 13 1 9 2
6 0 9 3 13 9 2
15 9 13 0 2 15 13 0 1 9 15 15 15 3 13 2
6 1 9 13 0 11 2
26 9 1 0 9 15 7 9 13 1 9 14 3 7 7 9 2 9 2 9 13 1 15 13 3 0 2
8 11 15 3 3 13 1 9 2
18 3 9 13 9 0 0 9 2 15 4 13 13 7 1 0 0 9 2
22 2 1 15 15 3 13 7 1 0 9 12 9 3 2 15 13 2 2 13 11 11 2
11 9 10 9 9 0 11 11 3 13 1 9
9 16 9 13 2 15 13 14 3 2
4 13 1 0 2
19 1 9 11 11 2 11 13 0 0 9 11 11 1 9 10 9 11 11 2
11 9 11 13 1 0 9 2 1 0 9 2
16 9 13 13 0 9 9 2 15 15 13 1 9 1 0 9 2
19 11 13 1 9 10 0 9 9 1 0 9 9 12 1 9 0 11 11 2
12 1 9 13 3 1 9 0 13 1 0 9 2
16 3 13 1 11 9 9 2 15 1 9 12 13 0 0 9 2
22 15 0 0 15 13 1 12 0 9 2 10 9 9 13 13 3 12 9 1 12 9 2
4 15 13 15 2
18 11 15 13 1 12 1 9 13 0 9 2 15 3 3 13 9 9 2
23 3 13 10 9 2 3 15 9 13 11 11 1 9 9 1 9 2 2 2 13 15 0 2
24 0 9 1 10 9 3 3 13 0 2 3 13 7 13 9 9 2 9 2 9 7 0 9 2
7 13 13 14 12 0 9 2
17 12 2 9 1 9 9 9 1 0 9 0 9 15 13 1 9 2
7 12 2 0 0 1 11 2
10 15 13 9 7 13 15 15 3 13 2
33 7 2 13 2 14 15 3 10 9 7 9 13 9 1 0 16 3 0 9 2 13 15 0 9 2 16 9 15 13 2 1 0 2
10 9 11 11 2 11 13 1 10 9 2
20 11 13 1 9 0 9 1 9 2 16 9 15 13 3 2 3 1 15 13 2
6 13 3 1 15 0 2
36 9 13 3 3 1 11 11 2 9 9 11 11 2 2 9 0 9 11 2 15 13 9 1 9 0 9 0 15 13 9 1 0 9 1 11 2
15 10 0 9 1 9 9 13 0 2 0 9 1 0 9 2
32 0 9 13 3 11 11 2 15 13 0 9 1 9 9 2 1 15 15 13 2 9 2 1 0 11 2 3 9 2 3 9 2
5 7 13 9 0 2
29 13 15 15 3 13 9 9 1 9 2 0 9 13 0 2 1 0 9 15 9 13 2 16 13 15 10 0 9 2
10 7 3 4 13 13 1 9 1 9 2
6 15 9 2 15 9 2
22 9 1 9 3 13 7 1 11 1 9 0 0 9 1 9 9 2 1 15 15 13 2
13 11 11 13 11 11 1 0 0 9 1 9 11 2
22 1 9 13 15 9 1 12 2 9 2 3 13 9 9 12 9 1 12 9 0 9 2
7 3 2 16 13 1 15 2
10 9 1 9 12 0 9 0 2 9 9
9 9 0 13 10 9 1 0 9 2
32 13 15 10 9 2 3 0 2 13 3 0 13 1 0 9 7 0 9 2 9 2 9 7 0 9 15 13 2 14 9 13 2
7 0 9 3 13 9 12 2
14 15 1 15 13 3 12 2 9 2 7 3 0 9 2
49 7 15 9 12 13 1 11 9 12 2 0 11 13 13 1 9 12 2 9 9 15 13 1 9 12 7 0 11 7 11 13 1 9 9 2 1 10 9 2 2 3 2 1 0 9 2 2 2 2
6 7 11 9 13 9 2
15 9 9 15 1 9 12 13 1 0 11 1 9 2 12 2
10 1 15 15 7 9 3 13 2 2 2
21 1 9 13 1 9 0 9 2 11 11 2 2 0 1 9 9 1 12 2 9 2
25 1 9 7 0 2 9 2 13 2 15 13 13 0 9 1 0 2 0 2 9 2 0 11 9 2
24 3 13 1 9 14 0 9 11 11 1 9 0 9 2 9 11 7 11 11 16 9 0 9 2
11 1 0 2 16 0 9 0 9 3 13 2
14 16 0 0 9 7 9 13 2 3 1 0 0 9 2
21 0 2 9 0 7 1 9 2 11 9 12 15 13 1 9 2 9 9 7 9 2
17 3 15 13 10 0 0 9 2 7 1 9 13 9 2 9 0 2
28 11 13 9 2 13 10 9 0 9 1 9 7 0 9 13 9 0 9 1 10 9 2 9 9 9 11 11 2
23 1 9 9 3 9 2 9 2 9 2 3 2 0 2 9 2 0 9 2 9 2 2 2
44 11 11 16 2 9 2 1 9 11 11 13 3 1 15 2 16 4 1 3 0 9 7 0 9 13 0 9 2 13 15 3 9 0 9 2 3 13 0 9 7 0 0 9 2
28 3 2 0 2 13 9 2 12 9 0 2 3 0 2 3 0 7 0 2 0 15 1 9 7 9 2 2 2
7 13 2 16 15 13 13 2
24 0 9 1 11 15 3 13 1 9 15 9 2 16 16 4 15 1 15 0 3 2 13 2 2
15 15 13 9 2 0 9 7 9 2 3 15 13 1 15 2
20 7 0 13 9 9 1 9 13 9 2 1 15 4 7 0 9 13 0 9 2
2 0 9
24 13 15 13 0 0 9 1 9 9 1 9 2 3 15 9 11 2 11 11 2 13 9 9 2
43 7 9 9 9 2 10 9 13 3 9 11 2 13 9 11 11 7 9 11 11 2 3 7 3 2 2 7 7 15 1 12 2 3 0 2 0 9 2 13 2 13 15 2
52 3 0 9 2 0 9 7 9 2 3 9 1 0 9 2 1 0 9 3 15 0 9 1 9 9 0 2 0 1 9 7 3 0 2 7 3 7 9 0 9 2 16 3 3 15 1 0 9 3 13 13 2
41 1 0 2 3 7 0 9 14 2 7 13 3 0 9 1 9 2 3 9 13 9 2 10 0 9 13 1 9 7 1 0 9 3 13 2 15 1 15 13 2 2
22 16 13 7 10 9 1 9 7 9 1 10 0 0 9 2 3 13 16 1 9 13 2
2 9 3
2 11 2
33 0 0 9 9 11 11 2 1 0 0 9 9 9 0 9 1 0 9 9 1 11 2 11 2 11 2 13 1 9 0 9 9 2
4 11 11 11 2
36 0 0 9 2 1 15 0 3 1 9 11 2 9 11 7 9 1 11 2 13 1 9 1 12 9 1 0 9 9 1 9 1 9 11 11 2
7 12 9 1 2 2 2 2
36 1 0 9 3 0 0 9 2 12 1 9 12 2 13 11 11 2 1 0 9 2 0 9 10 0 9 2 13 0 9 11 11 1 0 9 2
1 9
9 0 14 9 15 13 3 1 11 2
15 13 9 0 7 11 1 9 11 2 11 7 11 2 11 2
17 1 0 0 9 1 11 13 3 7 3 11 1 9 1 9 9 2
13 0 9 11 13 3 1 9 9 9 9 9 11 2
22 0 9 1 9 11 11 13 3 1 9 9 11 2 11 2 9 1 0 9 0 9 2
7 0 9 13 1 10 0 9
7 11 2 11 2 11 2 2
12 0 9 13 3 1 12 0 1 9 0 9 2
26 0 11 11 0 2 11 13 1 10 9 1 11 12 2 11 12 9 1 9 7 12 1 0 0 9 2
22 1 9 2 15 13 0 9 7 13 1 9 2 13 9 0 9 2 0 1 0 9 2
7 1 9 13 9 9 11 2
19 0 9 13 1 9 9 9 9 12 1 9 2 15 4 13 1 9 11 2
16 1 9 13 9 2 1 15 10 0 9 13 12 2 9 11 2
16 11 4 0 0 9 13 1 0 0 9 2 3 4 3 13 2
19 0 9 9 3 13 15 2 16 13 1 9 1 9 9 10 1 0 9 2
16 9 9 1 0 9 13 1 9 3 9 7 9 1 0 9 2
3 3 13 2
28 9 2 3 13 1 11 3 7 3 2 1 11 3 2 1 11 14 3 2 1 3 0 9 9 7 7 9 2
26 0 9 12 7 12 9 2 9 2 0 12 7 12 9 2 9 2 1 12 9 1 12 9 2 9 2
4 0 0 9 2
17 1 9 7 1 9 13 1 11 3 3 2 3 1 9 3 9 2
14 0 9 12 7 12 2 0 12 7 12 9 2 9 2
10 2 1 11 13 3 3 7 3 2 2
30 1 9 13 9 1 12 2 12 7 13 1 12 2 12 2 9 13 1 9 1 12 2 12 7 13 1 12 2 12 2
10 9 9 2 0 9 12 9 2 9 2
8 0 9 13 12 9 2 9 2
5 0 9 2 11 2
5 0 9 1 0 9
13 13 0 2 16 9 9 9 3 13 1 9 15 2
10 2 14 2 7 3 4 1 15 13 2
17 9 1 9 1 15 3 3 13 2 3 15 13 1 9 9 13 2
14 3 13 1 9 7 1 9 9 2 1 9 4 13 2
16 1 15 2 15 15 1 9 13 2 4 0 9 9 13 9 2
13 7 9 1 11 1 10 9 13 3 0 0 9 2
20 2 1 9 13 13 0 9 9 2 15 13 1 9 9 13 14 0 0 9 2
9 16 15 9 12 13 2 4 13 2
13 9 9 9 14 13 2 16 2 9 13 13 2 2
14 9 13 13 7 0 9 2 15 13 0 9 9 12 2
14 9 7 13 2 16 13 15 4 14 9 1 9 3 2
12 9 13 3 13 9 1 9 1 15 0 9 2
27 3 4 7 3 13 2 7 1 0 9 11 1 11 1 11 2 7 1 0 7 0 9 1 9 9 13 2
10 9 1 9 1 9 3 13 13 0 2
21 9 1 9 9 12 13 3 13 0 9 12 9 7 1 15 3 12 9 0 9 2
11 9 13 10 9 1 0 0 9 1 11 2
21 9 9 2 7 9 9 2 13 9 1 9 9 7 13 1 0 9 1 9 9 2
20 1 15 9 13 9 9 9 1 9 9 2 1 9 9 1 0 9 9 2 2
12 9 9 13 13 7 13 3 16 0 9 9 2
9 1 9 7 9 9 13 10 9 2
27 2 10 9 1 10 9 13 1 10 9 9 2 13 2 15 13 1 9 2 2 13 15 0 9 9 9 2
13 0 9 12 4 15 13 13 1 0 9 0 9 2
25 1 9 15 13 2 16 9 0 15 1 9 2 13 9 9 1 3 16 9 9 1 9 10 9 2
22 10 9 9 9 1 9 9 13 2 16 0 9 2 4 1 9 9 9 13 9 2 2
9 15 13 1 1 0 0 9 0 2
13 1 10 9 0 9 13 13 0 9 7 0 9 2
20 15 7 3 0 9 9 9 13 2 2 1 10 0 9 13 2 15 13 2 2
14 13 9 2 16 0 9 13 12 12 9 1 0 9 2
15 9 9 3 1 10 9 13 1 0 9 9 9 9 9 2
21 1 0 0 9 13 10 9 0 3 1 0 0 9 13 0 9 1 12 9 9 2
30 0 9 13 1 9 9 9 2 12 1 0 9 9 9 9 12 2 15 13 0 9 9 9 13 1 0 9 12 9 2
16 3 4 7 3 13 2 9 12 7 9 10 9 13 10 9 2
23 16 9 9 3 13 3 16 0 0 9 1 9 1 9 2 13 3 7 1 9 10 9 2
3 9 1 9
5 11 2 11 2 2
30 9 9 9 2 0 3 9 9 9 7 9 9 1 9 9 9 2 13 9 2 16 1 9 13 13 1 9 0 9 2
26 3 16 9 0 2 0 0 9 2 13 15 0 2 9 9 2 9 2 1 10 0 9 1 0 9 2
9 0 9 1 15 13 13 1 9 2
26 2 3 7 13 1 9 2 15 13 2 16 0 9 13 9 2 2 13 15 1 9 9 9 11 11 2
14 2 9 9 0 9 7 9 13 13 9 9 7 9 2
10 9 13 13 7 3 0 9 3 9 2
13 1 9 13 1 0 9 0 0 7 0 9 2 2
18 9 9 15 1 9 13 3 1 0 0 9 7 0 9 1 9 9 2
10 16 13 0 0 9 2 13 3 0 2
6 1 9 7 3 13 2
8 9 9 1 15 4 3 13 2
34 0 0 9 11 2 15 13 9 1 0 9 9 9 2 3 13 2 16 0 9 0 1 11 1 9 9 13 13 1 15 1 10 9 2
19 2 1 11 4 3 13 7 0 9 2 2 13 9 11 2 9 9 11 2
25 1 11 13 7 1 2 0 9 1 0 9 1 9 10 9 2 7 4 9 13 1 9 3 2 2
17 0 0 9 2 3 0 9 9 2 13 3 9 1 0 9 9 2
11 0 9 15 13 1 0 9 1 0 9 2
4 0 9 13 9
2 11 2
24 9 1 9 12 0 9 1 11 4 13 4 13 1 9 2 15 3 13 9 9 0 9 11 2
35 0 9 2 15 4 13 13 0 9 1 9 1 9 11 2 4 13 3 13 9 0 9 1 0 0 9 2 15 10 9 1 0 9 13 2
33 3 3 13 2 1 9 1 15 2 1 15 1 12 9 4 9 13 2 4 13 9 9 2 7 15 1 12 2 12 7 12 9 2
10 0 9 13 3 13 1 0 0 9 2
16 9 4 13 3 1 15 2 15 13 13 0 9 1 10 9 2
19 1 9 0 9 1 9 4 9 13 9 0 9 1 9 0 15 0 9 2
23 9 3 3 13 13 14 12 9 9 1 9 0 0 9 2 16 4 13 4 13 10 9 2
28 0 9 2 9 0 9 1 9 0 9 9 2 15 3 4 1 12 9 13 0 9 2 4 3 3 13 9 2
27 9 13 9 9 2 16 4 13 0 9 1 9 15 2 16 1 12 2 9 13 9 0 9 1 9 9 2
13 0 9 1 0 9 9 9 12 3 7 13 1 9
29 10 9 15 3 1 0 9 9 9 13 9 1 9 1 9 9 12 2 15 13 1 12 9 13 0 9 9 9 2
16 13 7 0 2 16 15 9 3 3 1 0 9 1 11 13 2
26 13 15 13 2 16 9 12 4 13 1 9 1 0 2 9 7 0 9 15 13 14 9 9 9 9 2
32 0 9 16 0 9 9 3 13 13 1 9 1 9 0 9 1 0 9 7 9 13 0 9 2 9 2 9 2 15 13 13 2
27 9 9 9 2 15 15 13 13 13 2 15 3 13 2 16 9 3 1 9 13 7 13 15 1 0 9 2
11 15 13 9 9 9 0 9 1 9 9 2
5 13 15 7 9 2
23 2 9 9 1 9 3 13 2 2 13 3 1 10 9 11 11 1 9 1 9 11 11 2
17 2 13 2 14 9 9 13 2 13 13 2 16 13 0 2 9 2
12 13 15 2 16 10 9 1 9 9 13 2 2
10 1 11 11 13 9 9 1 9 9 2
22 3 3 7 13 13 9 9 7 9 9 2 15 15 3 13 9 1 12 1 12 9 2
3 9 3 11
2 11 2
27 1 0 9 4 0 9 1 0 9 1 12 2 12 2 12 13 0 9 11 2 15 9 13 1 9 12 2
14 9 9 2 3 9 2 0 1 9 11 2 13 11 2
22 1 0 9 7 9 13 0 9 0 0 9 1 9 9 2 15 4 3 13 4 13 2
16 9 11 2 10 9 13 3 1 11 2 13 9 1 9 12 2
8 9 0 9 12 2 9 1 11
5 11 1 9 0 9
7 11 2 11 2 11 2 2
15 0 7 0 9 15 13 1 0 9 12 2 9 1 11 2
17 13 15 3 0 9 11 11 9 1 0 9 9 0 9 0 9 2
23 11 13 2 16 0 9 9 12 9 13 9 0 9 2 0 9 7 0 9 1 0 9 2
22 2 13 1 0 9 1 9 2 16 15 13 0 9 7 13 15 1 9 12 1 12 2
40 1 0 0 9 15 13 9 9 2 9 9 7 9 9 2 7 16 4 15 13 2 13 15 9 2 2 13 11 1 9 2 15 13 10 9 1 0 0 9 2
22 0 9 9 9 4 1 10 9 13 9 0 9 2 15 4 1 11 13 9 1 9 2
17 13 9 2 16 9 4 13 13 13 1 9 9 7 13 1 9 2
21 11 3 13 2 16 11 1 9 0 9 12 2 9 12 13 11 9 0 0 9 2
43 9 0 9 11 11 1 15 7 9 13 2 16 9 1 0 9 11 13 3 1 10 9 2 16 9 3 13 7 13 14 1 0 9 2 3 15 13 1 12 0 9 11 2
11 2 13 2 15 13 15 1 9 0 9 2
10 3 4 1 15 13 2 2 13 11 2
21 11 2 11 2 11 2 9 1 0 9 2 1 9 13 1 9 0 9 9 9 9
24 0 9 11 11 7 10 9 0 9 11 11 15 13 1 0 9 9 9 0 9 0 9 1 11
3 13 0 9
7 1 11 11 1 9 3 11
27 9 3 11 2 15 3 1 11 7 11 2 11 13 0 9 9 0 9 2 13 1 0 9 11 1 9 2
16 13 4 15 7 12 1 9 9 2 9 0 9 11 11 11 2
24 3 3 13 9 1 9 11 11 7 11 11 1 12 9 7 15 1 9 0 1 0 7 0 2
7 2 15 13 3 0 9 2
19 9 7 3 9 4 15 3 13 13 2 16 9 13 1 0 9 0 9 2
21 9 1 0 9 11 7 10 0 9 13 3 13 9 9 2 15 3 13 1 9 2
13 13 3 1 9 2 7 1 9 15 1 0 9 2
24 9 10 9 4 13 13 7 9 0 1 0 9 9 7 9 2 15 4 13 0 9 11 2 2
14 13 1 9 0 9 2 15 4 13 13 0 9 11 2
16 2 1 9 13 3 13 1 9 13 0 0 9 1 12 9 2
24 1 15 4 13 13 10 2 0 9 2 2 15 13 3 9 11 7 4 13 1 0 9 9 2
22 10 0 9 7 9 9 7 13 13 9 10 0 9 2 7 0 0 9 1 10 9 2
19 1 0 9 13 9 0 1 0 0 9 2 15 4 13 3 1 0 9 2
20 3 11 3 3 13 2 16 13 9 0 2 1 15 13 9 7 0 9 9 2
11 7 0 9 1 0 9 13 0 0 9 2
26 13 1 9 15 13 2 15 15 3 13 2 15 13 3 13 7 1 10 9 4 13 1 11 0 2 2
16 13 15 2 16 4 0 13 11 16 0 0 9 1 15 3 2
18 2 11 15 13 13 3 9 0 1 0 9 7 3 0 9 1 9 2
31 13 13 3 9 0 2 7 13 0 13 9 9 3 2 16 4 13 0 14 1 15 0 7 0 9 2 7 7 1 9 2
15 3 3 3 2 3 15 13 1 9 0 7 0 9 2 2
20 13 15 9 2 16 13 13 0 7 0 11 1 9 0 1 9 1 0 9 2
19 2 7 15 2 7 15 0 1 9 11 4 1 9 1 9 9 3 13 2
17 13 1 9 3 7 9 1 9 2 1 15 11 13 16 9 0 2
43 13 3 1 9 1 0 9 9 2 7 1 15 13 3 0 9 2 2 1 9 9 2 9 9 9 2 7 15 14 1 9 7 7 9 2 0 9 7 1 0 9 2 2
15 10 9 15 13 1 0 9 11 2 15 13 0 9 9 2
15 13 3 1 0 2 3 0 11 0 0 9 9 1 9 2
24 2 13 15 13 2 16 11 2 0 1 9 9 0 9 2 15 4 15 3 13 0 9 9 2
32 7 3 15 3 13 0 0 9 1 11 2 15 4 15 13 13 16 0 0 9 2 0 1 0 9 7 0 9 0 9 2 2
17 13 15 2 16 9 13 0 10 0 9 1 15 7 11 3 13 2
21 2 16 15 10 9 2 3 13 2 13 1 0 9 7 9 11 2 3 3 14 2
34 13 2 16 11 4 13 9 13 0 9 9 2 9 7 0 9 0 1 15 2 16 4 15 9 13 1 9 10 9 3 2 3 3 2
54 7 13 9 2 13 2 14 13 0 9 16 9 0 9 2 13 15 3 3 13 0 9 1 0 9 2 15 9 13 2 0 9 2 0 9 2 9 0 9 2 0 9 1 9 1 0 9 2 0 9 9 7 3 2
17 15 15 13 1 9 13 9 1 0 0 7 0 9 0 10 9 2
16 13 3 1 10 9 1 9 7 3 2 7 1 9 3 2 2
19 10 10 0 9 7 13 2 16 4 3 3 13 1 0 9 11 1 11 2
7 13 4 1 15 13 9 2
13 2 13 13 2 16 11 13 13 16 0 0 9 2
24 7 15 3 13 13 15 1 0 9 2 15 4 13 9 13 1 9 3 16 3 1 9 2 2
14 13 15 2 16 0 9 1 11 13 13 1 9 9 2
11 2 15 15 13 7 3 13 10 9 2 2
4 13 15 11 11
4 9 2 11 2
2 11 11
2 0 9
3 11 13 9
5 9 4 13 3 13
25 1 9 9 13 9 11 11 13 1 15 2 16 0 9 13 12 9 7 1 9 13 9 9 9 2
7 13 15 0 0 9 11 2
15 3 1 9 13 9 9 11 9 0 0 9 1 12 9 2
19 9 15 13 13 1 3 16 12 9 2 7 1 9 13 9 1 12 9 2
21 1 0 12 0 0 9 15 9 9 13 1 0 9 2 15 13 12 9 0 9 2
17 9 3 0 9 9 15 13 1 0 12 9 7 3 13 7 9 2
17 1 3 0 9 9 13 9 9 9 12 9 1 3 0 12 9 2
29 9 15 13 13 9 1 9 0 9 7 0 9 13 13 1 12 9 7 13 12 9 9 2 12 9 2 9 2 2
15 13 15 3 9 9 1 0 9 16 0 9 7 0 9 2
11 1 0 9 13 13 9 1 9 1 9 2
17 16 9 9 2 9 7 3 0 9 4 13 13 1 3 0 9 2
3 9 1 9
24 9 12 9 0 0 9 1 11 7 11 13 0 9 1 9 2 15 13 13 1 0 0 9 2
14 10 9 13 1 9 12 9 2 16 9 13 12 9 2
30 9 0 9 11 11 1 9 1 9 9 13 2 16 9 0 9 13 9 1 0 9 7 13 15 1 0 9 0 9 2
13 1 10 9 4 15 0 9 13 2 13 11 11 2
8 1 11 0 0 9 11 11 11
3 0 9 11
2 11 2
5 2 1 10 9 2
24 9 0 11 11 13 3 0 9 9 9 0 9 1 0 11 1 0 9 0 11 12 2 12 2
8 11 13 0 11 3 0 9 2
14 0 9 2 11 2 11 2 11 2 2 12 2 12 2
5 0 9 1 0 9
9 11 13 3 16 9 9 0 9 9
16 0 9 11 2 9 9 2 13 0 0 0 9 9 12 9 2
19 13 15 3 1 0 9 1 0 9 9 9 9 1 9 1 9 11 11 2
17 9 13 9 11 2 15 13 3 0 0 1 11 2 0 9 11 2
40 2 11 15 15 16 9 3 13 7 9 1 15 13 0 2 2 13 9 9 11 11 2 2 7 9 12 0 9 11 12 9 13 1 9 0 0 16 0 2 2
39 1 11 13 13 7 9 9 11 11 11 2 15 1 9 13 2 2 9 10 9 1 10 9 13 3 12 9 7 3 13 13 2 16 13 10 9 13 2 2
28 1 9 11 3 2 3 3 13 9 7 15 15 1 9 9 13 2 13 9 11 2 16 9 13 9 0 9 2
27 11 11 2 9 9 11 11 2 15 11 13 2 13 2 16 10 9 15 13 13 9 3 1 9 0 9 2
11 11 7 11 13 1 0 7 0 12 9 2
21 9 1 0 2 1 12 2 9 12 9 2 1 0 12 2 1 0 12 2 3 2
18 9 11 2 15 13 9 0 9 2 13 0 9 1 9 3 1 9 2
7 13 1 15 3 3 3 2
23 1 9 2 3 13 1 15 9 13 2 13 9 11 2 2 13 4 15 15 2 7 9 2
9 13 4 0 15 1 15 13 2 2
13 1 9 13 4 0 9 1 9 7 0 0 9 2
54 3 4 13 0 9 0 2 1 15 13 12 9 2 3 2 10 0 9 11 1 9 1 11 2 0 11 2 0 11 7 11 2 0 0 11 2 0 11 1 11 7 11 2 15 13 1 11 0 0 9 1 9 12 2
18 1 1 0 9 0 9 1 9 13 3 9 0 2 0 13 7 9 2
21 1 9 12 1 9 13 4 7 9 0 0 11 11 2 15 3 1 11 15 13 2
17 13 15 1 15 2 16 4 13 11 2 7 0 9 11 13 3 2
22 12 2 9 0 0 2 1 0 0 9 11 0 0 2 15 13 1 9 12 2 9 2
33 1 9 3 13 3 2 10 0 9 13 3 0 0 9 1 12 1 0 0 9 7 1 10 9 1 10 9 15 3 13 10 9 2
3 9 1 9
11 2 13 15 3 0 2 3 4 15 13 2
5 13 4 0 9 2
32 1 12 9 3 1 9 7 3 3 13 1 9 2 2 2 2 2 13 9 1 9 3 1 0 11 0 9 11 11 11 11 2
15 9 11 1 9 0 9 11 11 13 0 9 1 0 9 2
16 10 0 9 13 12 9 1 12 2 9 15 15 13 12 9 2
8 13 15 13 0 9 2 2 2
23 7 2 9 11 12 2 12 15 13 1 12 2 12 2 11 3 13 2 7 9 3 13 2
18 9 15 13 1 12 2 16 15 13 0 9 2 1 15 9 9 13 2
20 11 11 14 3 13 1 9 2 2 9 9 2 1 9 15 15 15 13 2 2
7 0 9 0 9 1 11 2
15 3 9 2 12 1 10 0 0 9 2 15 13 1 9 2
27 13 13 9 1 9 1 0 9 1 0 11 2 7 2 1 9 15 1 9 9 9 12 2 12 2 13 2
13 15 3 2 16 0 9 0 9 13 9 1 11 2
16 16 13 9 9 15 9 3 12 2 12 2 4 13 3 9 2
28 1 9 13 1 0 9 1 11 2 9 9 2 11 1 11 11 11 2 2 12 15 13 9 7 0 13 1 2
38 11 2 2 9 13 13 1 0 7 0 2 9 10 9 13 0 2 16 15 15 3 13 2 14 13 7 9 9 11 11 2 14 15 13 13 9 2 2
18 9 2 1 9 4 13 9 3 0 9 1 11 1 0 0 1 11 2
29 1 11 0 11 13 9 1 11 7 11 2 15 15 13 13 2 16 4 13 1 11 2 7 15 13 2 3 2 2
29 11 3 13 13 2 13 15 7 1 9 13 2 11 7 11 1 11 3 13 2 7 3 4 0 9 13 1 9 2
28 15 13 3 9 1 11 7 11 1 9 12 2 12 2 1 9 7 9 12 2 12 2 1 9 12 2 12 2
7 0 9 15 13 7 9 2
20 3 9 11 2 15 13 11 2 3 13 9 9 9 11 7 11 9 9 11 2
7 12 13 13 9 1 11 2
19 9 11 7 11 15 13 1 9 9 13 2 16 1 10 9 1 9 13 2
3 11 3 0
71 1 0 12 9 0 9 9 11 2 11 1 9 1 11 15 3 13 11 1 0 11 12 2 1 0 9 13 0 0 9 2 14 1 12 2 12 2 3 2 12 2 12 9 2 1 12 9 11 2 12 2 11 2 12 2 11 2 7 1 0 9 9 15 13 0 9 1 0 11 11 2
25 0 0 9 2 11 11 2 11 2 2 13 1 9 0 2 1 12 2 12 9 2 1 10 9 2
30 11 1 0 11 12 13 12 2 9 2 12 2 12 9 2 2 7 1 10 0 0 9 15 13 9 0 0 9 11 2
19 9 9 7 9 15 13 2 3 13 11 2 11 2 7 11 2 11 2 2
2 11 13
22 0 9 11 11 15 1 10 0 9 11 11 13 0 9 7 3 1 9 13 0 9 2
23 0 9 13 2 16 11 13 1 0 0 9 7 13 13 1 9 1 0 9 1 11 11 2
18 1 10 9 4 13 4 13 7 9 1 12 9 1 9 1 0 9 2
22 0 9 2 15 11 1 9 13 2 4 13 2 7 0 9 13 1 12 9 9 3 2
12 9 1 9 1 11 15 1 0 9 13 3 2
3 9 2 9
1 9
24 11 2 11 11 3 13 2 16 10 0 9 13 12 0 11 11 11 2 15 3 13 11 11 2
5 11 2 0 9 2
18 0 9 11 11 13 3 1 11 0 0 9 1 0 9 9 12 9 2
12 13 3 11 11 2 12 9 2 1 0 9 2
11 9 13 1 12 1 0 9 2 12 9 2
10 1 12 13 11 1 9 1 11 11 2
13 1 9 9 13 0 2 9 1 12 12 9 3 2
6 3 15 13 1 9 2
14 1 12 9 13 0 2 0 9 13 7 13 1 9 2
27 2 16 4 11 13 3 12 12 2 13 4 15 9 2 2 13 15 11 11 7 13 2 2 13 3 0 2
6 3 15 3 13 4 2
17 3 15 4 13 13 2 16 4 13 3 10 9 3 1 9 2 2
6 9 11 13 1 9 2
11 3 7 12 9 2 12 9 9 7 9 2
12 7 13 7 1 0 9 9 1 9 12 9 2
9 11 13 0 9 7 3 13 0 2
8 12 9 3 13 1 0 9 2
15 1 12 9 2 1 9 1 12 9 13 11 3 13 9 2
7 9 11 15 13 0 9 2
9 1 9 0 9 13 0 12 9 2
7 12 9 13 0 12 9 2
15 1 9 1 12 9 13 1 0 9 9 12 2 12 9 2
10 1 12 11 13 1 9 3 1 11 2
22 11 13 1 9 9 9 1 10 9 2 7 0 9 12 2 12 13 12 9 7 9 2
3 9 15 13
4 0 9 0 9
27 12 0 9 2 3 2 0 9 11 2 13 1 11 1 0 9 1 9 2 15 15 13 1 9 1 9 2
24 9 9 15 7 13 1 15 2 16 1 9 9 15 13 13 2 15 13 9 1 9 10 9 2
17 3 15 4 9 13 3 1 9 2 3 13 0 9 7 9 9 2
18 0 9 13 1 9 12 2 1 9 13 9 11 2 11 7 0 9 2
2 0 11
56 0 9 2 1 9 9 0 9 9 2 15 0 9 11 11 13 1 9 11 1 11 11 7 3 15 3 1 0 9 3 13 10 0 0 9 2 3 15 3 11 3 13 2 1 0 9 11 13 12 2 7 11 12 2 2 2
16 2 0 9 4 15 13 2 16 1 11 13 2 2 13 11 2
9 2 7 15 13 3 14 0 9 2
10 7 3 15 13 1 10 9 15 0 2
8 3 15 13 13 10 9 2 2
9 3 15 11 3 13 1 0 11 2
24 2 0 13 2 16 15 3 3 13 1 9 0 0 2 2 9 9 11 9 2 0 9 9 2
19 3 1 12 9 15 13 2 16 4 3 13 13 2 7 3 15 15 13 2
16 13 15 15 14 3 2 16 3 13 12 9 1 0 9 2 2
10 3 0 9 2 10 0 9 1 9 2
11 2 3 14 2 0 9 13 0 9 2 2
5 9 1 9 1 9
12 9 9 9 12 11 11 13 1 0 9 1 9
42 2 16 15 13 2 3 13 15 1 15 9 7 13 15 1 15 9 2 2 13 15 11 11 2 12 2 2 12 1 0 10 9 15 9 2 1 0 9 0 9 11 2
26 9 9 9 12 15 3 16 0 9 13 1 9 1 0 9 2 15 1 12 0 9 13 3 12 9 2
17 2 15 15 13 1 15 12 9 9 2 15 3 10 9 3 13 2
20 1 0 9 7 0 9 4 7 13 10 9 7 9 2 16 4 15 13 13 2
11 3 10 10 9 4 13 2 2 13 11 2
11 2 1 12 9 15 7 3 14 3 13 2
27 15 16 15 13 3 1 9 0 9 0 11 2 11 1 0 9 2 1 15 4 13 0 0 9 10 9 2
14 7 11 4 3 13 13 10 9 3 7 13 4 15 2
22 7 3 15 13 2 16 4 15 13 13 2 7 16 15 3 13 2 13 15 9 2 2
10 1 10 0 9 13 11 3 14 0 2
11 1 9 12 9 9 9 13 9 9 12 2
21 2 7 15 13 10 9 2 14 7 14 13 9 2 3 4 15 15 3 13 2 2
15 15 7 9 13 2 1 9 0 9 3 1 9 9 12 2
21 2 13 4 3 12 1 10 9 2 16 4 13 13 1 10 9 3 12 9 9 2
7 15 14 13 2 13 15 2
11 3 9 1 15 15 13 3 1 9 2 2
14 1 0 9 2 15 11 13 2 13 0 9 12 9 2
15 2 13 15 9 2 10 9 7 3 10 9 2 9 11 2
20 13 4 15 15 1 9 7 13 15 12 9 2 16 4 15 13 1 12 9 2
8 13 1 15 3 0 9 9 2
19 13 3 0 9 2 13 4 15 1 9 7 3 4 15 1 15 13 9 2
11 13 4 15 2 13 7 13 1 9 2 2
22 11 13 1 0 9 1 9 7 3 13 14 3 9 2 15 15 1 9 13 1 11 2
8 7 3 1 10 9 13 9 2
23 2 10 9 2 15 13 1 9 16 9 2 15 12 9 1 9 13 1 9 7 3 13 2
12 16 4 1 15 1 9 13 3 3 9 2 2
17 0 9 2 3 0 9 7 0 9 2 15 1 10 9 3 13 2
13 13 1 0 9 7 3 3 15 13 1 9 11 2
13 2 15 3 2 16 4 13 1 9 2 2 13 2
3 1 9 9
39 12 1 9 2 0 1 9 1 11 2 9 11 11 1 11 2 15 13 13 0 9 1 0 9 2 1 11 13 7 3 15 13 9 9 9 1 12 9 2
37 11 11 15 13 0 9 2 1 15 13 2 2 1 9 12 2 12 2 4 4 13 9 1 0 9 2 15 13 13 9 2 11 1 9 0 9 2
10 9 9 4 1 9 9 13 9 9 2
5 3 4 15 13 2
36 1 9 15 13 9 2 11 1 0 9 2 16 4 15 1 9 13 1 9 2 3 0 9 2 15 4 15 13 1 9 1 2 0 2 9 2
13 13 4 3 3 9 1 9 9 1 9 10 9 2
25 3 15 13 7 9 9 9 11 2 16 4 15 1 0 9 1 11 13 2 16 15 15 3 13 2
34 3 1 9 4 7 13 13 1 9 2 16 10 9 13 13 2 16 15 13 13 1 0 9 7 16 4 13 1 9 13 12 2 9 2
11 1 9 0 9 4 13 1 9 2 11 2
16 1 15 13 0 9 2 16 14 9 13 0 13 7 1 9 2
27 3 4 15 13 2 16 13 1 0 9 2 15 13 9 1 9 2 7 16 9 13 0 14 1 12 9 2
37 15 7 13 2 16 9 13 2 16 4 13 3 2 0 2 2 0 2 9 2 9 2 2 2 0 2 16 13 4 13 12 2 7 12 2 9 2
9 3 4 15 13 9 10 9 11 2
11 15 13 9 2 16 13 13 15 13 9 2
15 15 3 15 2 13 2 9 7 13 4 15 1 0 9 2
13 1 9 4 13 9 1 9 0 9 1 9 9 2
16 1 9 4 3 13 0 9 9 0 9 7 13 15 1 9 2
16 15 9 13 3 1 0 9 2 7 13 13 2 16 1 0 2
10 13 4 13 0 9 9 1 10 9 2
7 3 1 15 13 13 9 2
13 7 15 13 16 0 9 1 0 9 0 9 2 2
4 3 11 11 2
44 13 2 16 0 2 0 9 2 0 2 1 0 0 9 2 16 4 15 13 0 0 9 1 9 2 15 3 3 13 13 2 3 0 9 14 2 7 15 1 15 0 0 9 2
4 12 9 9 13
8 7 9 0 9 13 10 0 9
18 0 0 9 1 15 13 0 9 1 9 1 9 1 9 12 1 11 2
37 0 9 3 1 11 1 0 9 13 2 7 0 2 15 13 10 9 13 2 13 0 9 2 15 15 0 2 9 1 12 2 9 1 10 9 13 2
32 13 2 14 15 3 0 12 9 0 9 2 7 9 15 10 0 9 3 13 13 2 3 1 10 0 0 9 13 9 1 9 2
23 1 9 9 0 2 9 13 13 15 0 2 10 0 9 2 15 4 13 1 0 9 9 2
30 1 9 10 9 13 14 3 0 0 9 2 9 1 9 9 0 2 0 9 2 9 9 0 9 2 9 0 9 9 2
19 0 9 2 11 0 9 1 0 9 11 13 9 2 4 1 10 9 13 2
31 16 0 9 1 0 9 2 0 9 13 15 3 1 1 9 2 0 0 9 1 9 7 3 2 15 15 4 13 0 9 2
13 13 9 7 9 2 1 0 7 0 9 7 13 2
10 0 9 1 9 13 9 0 1 9 2
23 3 15 1 9 13 1 15 2 3 3 15 13 1 0 9 2 1 15 15 0 9 13 2
18 13 15 1 15 3 9 2 15 3 13 1 9 1 9 10 0 9 2
19 13 1 9 2 16 15 13 9 0 2 15 3 15 1 0 9 9 13 2
28 7 13 3 2 16 1 9 1 11 7 11 2 0 9 13 12 2 3 2 12 9 2 4 15 13 3 3 2
34 7 16 4 1 0 9 13 9 2 15 13 0 2 2 3 3 0 9 4 13 13 2 16 10 0 9 13 1 0 0 9 9 3 2
20 0 9 10 9 13 2 16 9 15 3 13 13 1 0 9 0 9 0 9 2
50 13 2 10 9 2 1 15 13 13 11 2 11 2 11 2 9 2 11 2 11 2 11 2 11 7 0 2 13 1 0 9 0 9 2 1 9 1 9 0 2 11 2 1 9 1 12 7 12 9 2
11 0 10 9 3 13 3 0 1 0 9 2
31 9 14 13 2 16 1 9 15 1 15 15 13 14 3 7 3 2 1 0 9 7 9 9 2 3 2 11 7 0 2 2
17 9 9 4 15 7 3 13 9 1 9 13 1 10 9 16 3 2
40 9 1 0 9 1 0 9 13 13 3 16 0 9 2 16 0 0 9 4 13 1 9 1 0 7 16 12 1 10 0 9 15 3 1 10 9 13 3 3 2
6 9 13 1 9 11 2
20 0 9 11 11 15 13 0 9 1 9 2 15 13 1 9 0 0 0 9 2
24 13 15 3 1 0 9 9 11 11 11 1 0 2 0 9 2 1 15 11 13 12 2 12 2
6 11 13 0 0 12 2
17 1 9 13 12 0 9 2 3 3 13 2 12 13 12 2 12 2
18 0 9 11 11 11 13 2 16 0 9 1 9 9 13 9 1 9 2
5 9 13 12 9 2
22 11 13 9 1 12 9 7 13 9 0 9 2 15 3 13 9 1 9 1 0 9 2
8 3 13 1 12 9 0 9 2
2 11 13
14 9 11 7 9 11 13 13 0 9 9 11 11 11 2
20 15 3 13 1 0 9 12 9 9 7 3 13 13 0 9 1 12 9 0 2
21 1 9 15 13 3 14 12 0 9 2 12 1 12 9 7 12 1 12 0 9 2
5 1 9 11 0 9
14 11 2 11 2 11 4 13 9 2 0 9 12 2 9
5 11 2 11 2 2
14 9 1 9 9 9 4 9 13 1 9 12 2 9 2
16 13 1 15 9 1 9 3 0 12 2 9 11 12 0 9 2
16 13 4 12 0 9 2 15 13 13 9 9 1 9 1 9 2
40 1 9 9 1 9 9 13 15 9 0 9 2 15 13 2 16 4 9 1 9 9 4 13 9 9 2 3 16 4 9 1 9 9 4 3 1 10 9 13 2
28 11 11 2 11 2 13 2 16 4 15 1 9 1 9 9 9 13 3 2 16 4 15 9 13 13 0 9 2
14 1 10 9 7 13 0 13 14 1 15 9 9 9 2
15 9 15 3 13 2 16 3 1 10 9 13 9 0 9 2
10 0 9 0 9 9 13 9 9 11 2
28 0 9 1 12 2 9 13 1 9 9 11 11 2 11 2 11 11 11 2 9 0 9 0 9 2 0 9 2
44 1 0 9 1 15 13 1 9 9 3 12 9 2 13 15 12 2 2 1 0 9 9 9 12 9 2 13 15 12 2 7 1 0 9 11 11 12 9 2 13 15 12 2 2
16 1 0 9 13 2 7 11 11 9 11 2 11 2 11 13 2
30 3 1 9 13 9 12 1 0 9 11 11 2 11 2 2 16 4 15 9 9 13 2 7 1 10 9 13 9 9 2
30 1 9 9 9 9 13 3 12 1 9 11 11 11 2 11 2 11 2 2 15 13 1 9 7 9 1 9 10 9 2
26 11 2 11 13 2 16 2 9 9 4 15 3 13 13 9 2 16 4 1 15 13 9 7 9 2 2
22 1 9 0 9 15 4 0 9 9 9 13 12 2 9 2 3 3 1 10 9 11 2
18 0 9 4 13 2 16 4 3 3 13 2 16 13 0 13 0 9 2
29 9 0 9 11 11 3 1 9 11 11 7 11 11 13 3 1 11 1 9 1 9 0 9 9 9 0 9 0 9
2 0 9
2 11 2
48 11 11 15 3 13 1 10 0 9 2 13 3 0 9 0 0 9 11 11 1 9 11 1 9 1 9 9 11 11 11 2 11 2 11 2 2 16 11 11 13 9 0 9 1 11 1 11 2
23 0 9 11 11 13 0 0 9 7 0 9 0 0 2 9 11 11 15 13 1 3 0 2
26 13 3 1 15 2 16 1 9 1 9 1 0 9 13 11 11 13 3 13 9 1 9 1 9 9 2
47 1 9 1 9 11 3 11 11 13 2 16 13 9 2 16 15 11 11 1 11 13 1 9 1 9 2 13 1 0 9 11 2 1 15 13 16 9 0 9 1 9 9 11 1 9 11 2
4 9 11 7 11
2 11 2
35 9 9 11 11 11 3 13 2 16 1 0 0 9 0 9 2 11 2 11 13 0 9 2 7 9 0 9 11 13 9 0 9 1 9 2
32 2 0 9 13 2 16 10 9 13 1 9 11 2 15 15 13 1 11 2 2 13 11 2 11 1 9 2 15 3 13 11 2
44 11 11 1 10 9 13 2 16 0 9 9 11 15 13 2 3 9 0 9 9 0 9 2 2 7 13 2 16 2 0 0 9 4 13 1 0 9 1 0 9 1 11 2 2
4 9 1 0 9
1 9
4 9 1 0 9
19 0 9 13 0 9 9 2 15 4 1 0 9 13 13 1 9 0 9 2
38 0 0 9 13 1 0 0 9 0 9 3 2 16 1 9 3 2 3 0 9 0 9 13 10 9 3 13 1 0 0 9 2 3 13 9 3 0 2
10 16 1 9 13 0 9 2 3 13 2
19 3 14 15 1 9 10 9 13 2 16 15 1 11 15 2 0 2 13 2
58 0 9 0 2 9 2 11 2 9 2 11 2 7 13 2 3 1 9 12 2 9 3 7 1 0 9 1 9 13 13 2 10 9 7 3 15 3 1 12 2 9 9 9 13 2 13 9 1 9 2 15 15 1 10 9 13 3 2
21 2 9 13 0 2 2 13 3 2 11 11 2 0 9 9 1 3 16 12 9 2
36 15 1 9 15 3 3 13 1 0 9 2 16 9 9 13 0 9 9 2 3 7 1 9 2 15 4 1 11 7 1 9 13 9 0 0 2
40 1 9 2 16 9 1 0 9 7 1 9 1 9 1 11 13 1 9 1 9 1 9 2 15 1 0 9 13 13 9 2 16 0 7 0 9 9 13 9 2
33 9 10 9 13 0 9 2 1 0 9 9 1 9 4 15 3 13 2 16 2 1 9 13 1 0 9 0 13 3 15 9 2 2
23 9 2 13 0 0 9 2 9 9 13 12 9 7 0 3 12 9 1 9 13 0 9 2
11 16 3 14 9 9 2 3 14 9 9 2
24 0 13 7 9 2 16 0 1 15 2 15 3 1 9 13 13 3 2 1 15 3 3 13 2
35 1 15 15 1 9 11 13 0 9 2 3 2 3 13 9 3 2 13 3 1 9 2 7 1 9 1 10 9 15 1 9 13 2 2 2
17 15 3 13 1 15 2 16 0 0 9 15 13 1 9 3 0 2
17 7 0 9 13 3 1 9 1 0 9 16 1 9 9 3 13 2
6 9 9 11 13 1 11
39 2 13 2 16 0 9 3 13 1 15 2 16 4 0 0 9 13 12 2 9 12 2 2 13 15 9 9 1 0 9 7 9 11 11 11 2 11 2 2
13 1 10 9 13 7 0 9 13 7 1 10 9 2
29 0 0 9 7 13 9 1 9 0 0 9 0 9 2 9 11 2 3 1 9 10 9 2 3 1 10 0 9 2
40 9 1 9 9 11 13 13 1 9 11 11 13 1 0 9 11 10 9 3 3 2 16 15 0 9 13 1 15 2 16 13 13 0 9 13 9 2 7 9 2
17 13 3 2 16 9 0 9 13 1 0 0 9 3 1 9 9 2
32 11 7 3 9 1 9 11 13 1 9 2 7 10 9 13 1 12 2 9 12 2 3 4 13 0 9 13 10 9 1 9 2
8 9 11 1 11 11 13 3 2
26 9 13 1 0 7 0 9 1 9 12 2 12 7 0 2 0 9 15 13 10 9 2 15 15 13 2
38 1 10 9 2 16 15 1 9 11 13 9 1 9 0 9 11 2 15 1 9 12 13 1 0 9 9 2 11 11 13 2 16 15 1 15 3 13 2
13 2 9 1 9 9 11 13 1 10 9 0 9 2
18 10 9 4 13 1 9 0 9 13 0 9 1 0 9 2 2 13 2
52 9 9 1 0 9 7 9 11 11 11 2 11 2 1 9 9 1 9 9 11 13 2 16 13 0 15 3 13 3 1 10 9 2 16 4 1 0 9 11 1 12 2 12 2 12 13 0 9 10 0 9 2
22 1 10 9 0 9 3 13 1 15 2 16 4 0 2 9 12 2 9 10 9 13 2
40 1 10 9 2 3 4 13 9 0 0 2 0 9 2 16 13 9 1 0 9 7 9 1 11 7 0 9 2 11 11 13 2 16 15 13 1 3 0 9 2
22 2 13 15 0 9 9 2 15 14 13 13 2 16 4 13 3 1 12 7 0 9 2
16 13 0 13 9 7 0 9 2 7 9 14 3 2 2 13 2
23 0 4 1 10 9 13 2 16 4 15 12 1 9 13 13 10 0 9 1 9 3 3 2
28 1 10 9 13 2 16 0 2 0 9 13 3 1 9 11 7 16 15 0 0 9 0 9 13 1 12 9 2
28 0 9 9 11 11 2 15 9 1 0 9 7 9 3 13 2 15 13 2 16 10 9 3 13 10 0 9 2
14 1 9 10 9 13 1 10 9 0 9 1 12 9 2
1 9
2 13 9
9 0 9 13 1 10 9 1 11 2
33 3 13 1 9 0 9 3 0 0 9 9 11 11 2 16 15 2 15 15 1 11 13 2 13 13 9 7 13 13 0 9 3 2
45 3 0 9 13 7 9 11 7 9 11 11 11 2 16 9 13 2 16 11 16 0 9 4 15 13 2 16 4 13 1 0 9 2 3 2 0 13 1 10 9 2 9 13 2 2
14 1 2 9 2 10 9 13 2 16 3 13 1 9 2
16 3 13 15 0 2 16 16 4 13 9 13 9 10 9 9 2
11 3 15 13 2 16 4 13 10 9 13 2
23 12 9 4 15 3 13 13 7 13 2 16 0 2 15 15 3 13 2 13 9 7 13 2
10 9 1 0 9 11 11 2 13 4 9
2 11 2
34 9 9 11 11 11 13 2 16 13 1 9 1 9 0 9 0 9 10 0 9 2 15 13 13 1 9 2 3 9 13 16 9 11 2
19 13 15 1 9 2 15 15 1 0 9 13 1 11 2 11 0 9 11 2
13 2 1 10 0 9 4 13 2 13 7 13 4 2
30 15 9 0 1 0 9 4 1 0 9 13 7 13 15 3 9 0 1 10 9 2 2 13 9 9 11 7 9 11 2
24 0 9 9 11 2 11 2 16 1 9 9 9 13 0 9 2 13 1 15 3 0 7 0 2
36 2 0 9 1 0 9 4 13 1 9 9 12 7 12 7 13 1 9 12 2 3 4 13 13 2 16 4 1 9 13 9 9 2 2 13 2
34 0 9 0 9 13 1 11 2 11 15 0 9 7 4 3 0 9 13 3 9 9 2 3 0 9 9 11 2 7 3 9 9 11 2
14 2 3 4 3 13 9 9 2 14 9 1 9 2 2
14 9 12 2 9 12 4 11 2 11 13 9 0 9 2
24 2 3 4 13 10 9 2 16 1 9 9 0 9 15 13 13 7 13 10 9 2 2 13 2
25 3 0 9 1 0 9 0 9 15 11 2 11 1 10 9 13 2 16 2 3 13 2 15 13 2
11 2 15 9 4 13 1 3 0 9 2 2
45 3 11 11 13 3 2 2 0 3 0 9 13 0 9 13 1 9 9 0 9 1 11 7 11 9 11 7 10 9 7 3 13 9 7 0 9 7 13 0 9 1 0 9 2 2
4 0 9 3 13
5 11 2 11 2 2
19 1 0 9 3 16 12 9 0 9 11 13 3 3 13 14 12 9 9 2
37 10 9 13 3 1 9 0 9 11 1 11 2 15 3 1 0 9 13 0 9 12 9 11 11 0 15 0 9 1 0 9 9 12 2 9 12 2
28 1 9 0 9 15 9 0 9 11 11 11 13 2 16 9 1 0 9 9 1 0 9 13 1 9 10 9 2
13 2 9 1 0 9 3 4 13 1 0 9 9 2
22 1 10 9 1 12 0 9 4 13 1 12 0 9 2 16 10 9 13 2 7 3 2
28 15 3 13 1 15 0 9 2 16 0 9 15 15 13 2 10 9 13 9 7 15 3 2 2 13 11 11 2
18 9 0 9 11 13 9 2 16 15 1 9 3 3 13 9 0 9 2
4 9 0 9 11
5 11 2 11 2 2
30 12 12 9 9 11 2 12 0 9 7 10 9 13 0 9 0 9 1 0 9 2 15 13 1 9 1 11 2 11 2
20 0 11 4 13 1 9 12 2 13 3 0 0 9 2 16 13 0 0 9 2
20 3 1 10 9 13 1 0 9 1 11 9 12 9 2 0 2 11 12 9 2
19 9 13 2 16 13 15 9 11 0 2 13 15 7 13 1 1 0 9 2
1 9
4 9 1 9 2
20 12 9 13 1 11 12 0 11 9 2 15 13 1 0 9 9 10 0 9 2
11 11 13 2 16 4 9 13 9 7 13 2
8 3 4 13 1 9 1 9 2
4 9 1 9 9
5 11 2 11 2 2
25 9 1 3 16 12 9 9 3 3 13 1 0 9 9 2 15 13 12 9 7 9 1 0 11 2
35 3 0 10 9 9 13 1 11 1 11 2 3 1 9 0 2 11 11 3 0 9 13 0 9 9 2 9 7 0 9 3 1 0 9 2
3 0 9 9
6 0 11 2 11 2 2
15 0 9 9 9 11 1 11 15 3 13 11 11 1 11 2
18 1 9 13 9 11 13 9 1 0 9 3 1 12 9 1 0 9 2
15 1 0 12 12 0 9 13 13 1 0 9 0 12 9 2
7 3 9 13 9 9 9 2
13 1 9 0 9 4 15 3 9 11 13 13 12 2
32 2 1 0 9 13 13 3 12 9 2 2 13 3 9 9 11 11 2 2 13 1 15 9 0 9 2 10 9 13 13 3 2
11 2 1 11 4 13 3 7 0 0 9 2
13 1 0 9 9 9 13 13 9 7 1 0 9 2
6 3 13 15 3 0 2
11 1 0 9 1 11 13 3 12 9 3 2
10 3 13 9 13 0 9 14 12 9 2
14 13 15 7 1 11 2 11 2 11 2 11 7 11 2
3 11 13 9
5 11 2 11 2 2
26 3 7 3 13 11 1 9 0 9 7 13 15 1 0 9 15 1 9 0 9 11 13 11 7 11 2
30 1 0 9 9 1 9 9 9 3 9 11 11 13 2 16 13 1 0 9 0 1 0 9 1 10 0 7 0 9 2
11 9 11 13 7 0 1 9 10 9 13 2
25 9 7 13 2 16 4 10 9 13 9 9 1 9 2 9 1 9 9 7 9 0 9 12 9 2
25 9 11 11 11 13 9 0 9 2 15 13 1 9 9 11 11 7 13 3 2 13 9 0 9 2
1 3
3 9 13 11
30 11 4 1 9 11 11 11 13 1 9 0 9 1 0 9 7 11 2 16 11 13 9 11 1 0 9 1 9 9 2
3 9 1 9
5 11 2 11 2 2
14 9 9 13 1 9 1 9 1 9 1 11 0 9 2
19 3 13 9 9 1 9 1 9 1 9 11 7 13 2 16 13 1 9 2
11 10 9 13 9 2 15 12 0 9 13 2
17 1 12 0 9 13 9 9 1 0 9 7 9 0 7 0 9 2
9 9 3 13 0 9 7 0 9 2
11 13 4 15 11 11 2 9 11 7 9 11
18 13 15 2 16 0 9 1 0 7 0 9 13 14 1 9 0 9 2
28 2 16 13 9 0 7 13 15 2 16 13 0 2 3 15 13 13 16 9 1 11 2 15 13 9 9 9 2
10 1 10 9 4 7 13 13 9 11 2
14 9 0 9 13 1 9 0 9 13 15 15 1 9 2
16 14 3 13 1 9 9 1 9 2 16 1 15 13 0 9 2
32 1 9 13 0 7 13 3 2 11 3 13 0 9 1 9 9 0 9 2 16 4 13 9 1 9 9 1 10 0 9 2 2
1 9
4 1 11 1 11
13 3 12 9 1 9 0 9 13 1 9 9 11 2
12 1 9 11 11 4 15 13 1 9 3 3 2
17 1 0 9 2 1 9 10 1 0 0 9 14 1 0 0 9 2
17 3 0 0 9 13 1 9 9 2 16 9 9 9 15 13 9 2
31 3 15 13 7 9 2 16 10 0 9 10 9 0 9 2 9 2 9 13 7 9 4 15 13 13 1 9 9 0 9 2
10 7 9 15 7 13 13 2 15 13 2
12 13 15 3 3 12 9 2 15 9 9 13 2
8 12 1 15 13 3 9 0 2
19 15 2 0 2 3 9 3 13 3 2 16 1 0 12 9 13 0 9 2
15 13 15 3 3 2 16 1 0 0 13 0 9 10 9 2
17 0 9 1 9 9 7 13 13 0 9 1 9 1 0 0 9 2
14 10 0 9 4 10 0 9 13 3 16 10 0 9 2
36 1 0 9 13 3 1 9 9 2 16 10 9 4 1 9 13 13 3 9 7 0 9 7 13 9 2 15 1 9 2 16 0 2 13 9 2
13 1 9 9 1 11 1 11 15 3 3 3 13 2
3 9 1 9
6 0 11 2 11 2 2
21 3 1 0 9 3 3 13 1 9 1 9 11 1 0 11 9 1 0 0 9 2
13 3 13 0 9 1 9 11 7 13 15 1 9 2
11 1 12 9 13 13 3 1 0 0 9 2
8 0 0 9 13 9 2 2 2
12 3 14 0 9 13 9 0 11 2 9 11 2
17 10 9 7 9 13 9 9 1 9 12 9 0 9 1 9 9 2
29 0 9 3 15 13 1 0 9 2 3 11 11 13 9 2 15 13 9 11 1 9 0 9 1 0 9 0 9 2
27 1 9 15 13 7 11 11 1 0 9 0 9 1 0 9 7 0 2 9 2 11 11 2 9 0 9 2
17 1 0 9 13 1 9 0 11 12 0 0 9 2 3 3 12 2
7 0 11 7 11 2 9 9
5 0 9 1 0 9
7 0 11 7 11 2 9 9
22 9 12 2 7 12 2 9 10 9 15 13 1 0 9 11 3 1 10 9 9 9 2
13 9 10 9 13 7 0 9 2 3 0 0 9 2
35 10 9 15 13 3 1 0 9 1 0 9 0 9 9 2 13 15 7 1 9 10 0 9 7 13 15 3 3 1 15 9 9 0 9 2
27 3 15 10 9 15 1 0 0 9 11 13 7 1 9 1 0 0 9 7 1 9 10 1 15 1 9 2
25 3 13 9 2 15 13 9 9 7 1 9 1 3 0 9 3 13 7 9 7 9 0 0 9 2
25 1 9 0 11 7 11 13 3 1 0 9 10 0 2 16 3 0 2 7 3 14 3 0 9 2
3 14 0 9
38 9 12 2 9 13 1 0 9 11 0 1 0 9 0 9 2 15 13 3 0 0 9 9 9 2 12 2 7 0 0 9 2 12 2 1 0 9 2
36 0 0 9 0 4 3 1 0 9 1 9 12 1 9 13 2 3 13 13 1 15 1 0 9 9 2 13 7 3 1 3 0 9 1 9 2
12 3 15 13 0 9 9 1 0 2 0 9 2
23 15 1 12 0 9 15 7 13 9 10 9 7 13 13 3 7 3 10 9 13 7 13 2
16 9 0 9 13 3 0 7 9 10 9 13 0 9 7 9 2
23 3 0 2 0 0 9 9 12 2 9 13 0 9 7 1 9 1 0 0 9 3 3 2
12 13 15 2 16 0 9 13 3 1 12 9 2
17 3 15 7 13 7 9 1 9 2 1 9 2 1 0 9 3 2
16 7 3 4 13 0 0 9 2 16 13 9 2 9 2 9 2
21 7 15 13 1 0 9 13 1 0 9 0 9 2 0 1 0 9 3 0 11 2
7 9 9 3 13 3 0 2
26 0 9 2 7 16 14 3 0 2 13 14 0 9 9 1 9 1 9 0 2 3 13 3 0 9 2
20 1 15 0 9 13 2 16 1 9 0 11 13 1 9 0 9 1 0 9 2
6 15 0 9 14 13 2
4 9 1 9 9
22 9 1 0 9 9 13 1 9 7 1 0 9 9 0 11 1 11 7 1 0 9 2
28 9 3 13 14 0 9 2 3 10 9 13 2 7 14 13 7 9 0 9 2 15 4 13 1 9 0 9 2
42 15 3 13 9 0 0 9 0 13 1 9 9 2 13 10 9 1 0 9 7 3 13 9 1 9 7 0 9 9 2 15 13 3 1 9 12 1 0 9 1 9 2
18 13 1 0 3 0 9 0 2 11 2 7 0 0 9 2 11 2 2
29 10 12 9 13 9 0 11 2 3 13 1 0 9 1 11 7 13 3 0 9 1 3 0 0 9 1 0 11 2
8 15 13 1 9 11 3 0 2
24 1 0 13 12 9 0 9 1 9 0 9 1 0 9 2 16 13 3 2 9 0 9 3 2
32 1 9 9 12 1 15 13 9 11 2 15 1 0 13 9 11 2 15 13 0 9 3 0 9 11 2 11 2 0 11 11 2
36 0 2 9 15 3 13 1 0 9 0 9 2 1 10 9 13 3 9 15 11 1 0 0 9 2 13 7 13 9 11 7 3 0 0 9 2
30 1 9 1 12 9 15 4 13 9 0 1 9 2 9 1 0 9 0 9 7 9 9 7 9 1 9 9 1 9 2
3 1 0 9
9 9 9 12 13 11 1 11 9 2
10 15 13 0 9 1 9 0 0 9 2
20 3 15 3 13 0 2 0 9 7 7 9 9 9 11 11 13 1 10 9 2
10 3 0 9 0 11 1 15 13 9 2
14 0 0 9 15 1 10 9 13 9 0 9 0 11 2
51 13 15 7 9 0 9 1 0 9 9 2 1 0 9 1 0 9 0 2 9 1 0 9 2 0 9 2 7 1 9 0 0 9 14 1 9 0 9 0 3 0 9 0 9 2 15 15 13 1 11 2
17 1 9 9 11 13 13 0 9 2 9 9 11 13 3 0 9 2
21 9 0 9 1 0 9 0 11 13 3 0 2 16 0 2 9 13 13 10 9 2
13 3 15 13 9 9 12 0 9 2 11 7 11 2
14 10 9 7 13 0 7 13 15 0 0 9 1 9 2
23 9 0 0 9 13 2 16 4 10 9 13 7 3 1 0 9 13 0 2 3 0 9 2
13 0 9 9 13 3 2 1 15 15 13 0 9 2
11 0 0 9 1 11 13 1 10 0 9 2
4 9 9 1 9
31 12 9 1 9 1 12 9 1 12 9 13 1 9 9 1 0 9 1 0 11 2 11 1 9 1 12 1 12 0 9 2
9 16 9 13 2 13 13 1 9 2
8 9 0 9 13 3 1 9 2
8 0 9 15 7 13 1 9 2
15 9 2 1 15 13 0 9 2 3 13 4 13 9 9 2
29 16 9 12 2 9 13 9 0 0 9 1 0 11 0 9 12 9 1 15 2 13 0 9 14 1 12 9 9 2
8 3 9 12 9 13 3 9 2
21 9 15 13 15 9 2 15 1 0 9 1 9 12 2 9 13 9 1 9 12 2
34 2 15 3 13 9 1 9 2 15 3 15 4 13 3 13 9 2 2 13 11 11 2 9 0 9 2 3 3 13 3 16 12 9 2
35 2 3 1 9 4 15 3 13 1 0 9 0 9 1 9 0 0 9 2 13 15 7 13 1 9 9 7 9 9 2 2 13 11 11 2
20 12 9 13 3 9 10 0 9 1 9 2 15 1 10 9 13 7 9 0 2
34 1 12 1 9 0 0 9 2 1 10 9 13 3 0 9 11 11 2 13 1 10 9 0 0 9 0 12 9 2 9 7 10 9 2
20 9 1 9 2 0 9 13 1 3 16 12 9 9 2 13 0 9 1 9 2
15 2 9 13 3 9 9 1 0 2 15 13 0 0 9 2
15 13 7 2 16 4 1 9 13 13 2 2 13 11 11 2
17 9 13 0 0 9 7 9 1 9 0 9 1 10 9 1 9 2
37 9 2 15 1 12 2 9 13 9 9 9 1 9 2 15 1 9 9 3 13 13 1 9 2 9 2 15 3 13 0 9 2 16 15 13 9 2
17 1 0 11 13 3 9 3 10 9 2 3 15 3 13 12 9 2
7 1 9 13 0 12 9 2
24 1 9 13 3 9 1 0 9 1 9 2 3 13 3 1 9 13 9 2 16 15 3 13 2
21 0 9 1 0 9 13 1 9 11 11 2 15 1 12 9 13 1 9 9 9 2
14 13 0 9 2 15 1 0 9 13 9 0 0 9 2
9 2 3 4 15 13 13 15 9 2
23 13 4 1 15 3 0 9 2 7 13 15 10 9 7 13 4 1 15 13 2 2 13 2
20 2 3 4 15 1 9 13 1 0 9 0 9 1 11 2 2 13 11 11 2
17 2 13 4 2 3 13 0 9 1 15 2 16 3 4 13 9 2
14 13 3 3 0 9 9 1 9 2 3 1 0 9 2
14 13 15 9 9 1 0 9 2 16 13 9 1 9 2
10 1 10 9 4 15 3 0 13 2 2
3 1 9 9
23 1 10 9 13 7 1 9 2 1 15 13 9 9 2 7 1 15 2 15 13 0 9 2
2 0 9
3 2 2 2
29 1 9 11 11 2 11 3 12 2 12 2 2 4 13 9 1 3 0 0 9 11 2 11 7 11 16 0 9 2
11 0 4 13 1 0 9 1 9 0 9 2
18 1 9 11 4 13 1 9 0 9 0 9 7 9 11 13 3 0 2
5 11 11 2 11 12
37 2 2 2 9 0 9 4 15 3 13 7 9 1 0 9 2 1 9 3 0 0 9 0 9 2 0 9 11 2 13 4 13 3 9 9 2 2
41 7 0 9 2 13 2 14 15 0 9 2 11 2 9 11 2 4 10 9 3 13 1 15 2 15 15 0 9 9 0 0 9 7 0 9 3 13 1 0 9 2
6 4 3 13 11 11 2
4 2 9 2 2
5 11 2 11 2 11
3 2 2 2
26 1 0 9 2 0 2 15 13 12 9 2 0 3 0 9 2 7 15 2 9 2 7 2 9 2 2
22 13 7 2 16 4 0 0 0 9 1 0 0 9 13 0 16 0 2 7 2 11 2
37 10 9 9 1 0 0 9 13 0 9 0 9 2 3 2 11 2 11 2 2 11 2 11 2 2 11 2 11 2 2 11 2 11 2 2 2 2
19 3 0 7 0 9 16 11 2 11 2 11 3 2 4 15 13 13 3 2
27 1 9 2 16 4 15 10 9 13 2 13 15 9 0 9 2 0 9 2 0 9 9 1 0 9 3 2
15 13 1 15 0 9 9 7 13 15 3 3 3 3 3 2
22 1 0 9 0 9 1 9 9 11 15 13 1 0 9 3 0 9 16 1 0 9 2
27 13 15 10 9 2 16 0 9 3 0 9 13 3 2 7 15 3 1 11 2 3 1 11 7 1 11 2
42 13 4 15 7 0 0 0 9 3 13 0 9 7 13 4 15 13 9 7 9 0 9 1 10 0 9 10 9 2 3 15 15 13 10 0 7 0 2 0 9 2 2
24 7 16 15 1 15 13 1 11 2 0 1 11 7 0 1 11 2 3 14 13 7 13 3 2
21 3 3 4 15 13 13 0 9 0 9 2 1 15 15 3 13 7 4 13 3 2
6 9 2 11 11 2 11
3 9 1 9
5 11 2 11 2 2
7 2 13 15 3 1 0 2
32 0 9 1 9 13 9 2 1 15 13 14 3 10 9 3 0 2 2 13 15 3 9 2 11 11 2 9 0 9 0 9 2
20 3 1 11 11 2 9 9 9 2 13 1 0 9 0 9 9 3 1 9 2
16 0 9 10 0 7 1 15 0 9 13 9 1 0 9 9 2
23 0 9 9 2 0 9 7 9 13 1 9 9 7 9 1 9 1 0 9 9 1 9 2
1 9
1 7
1 9
23 9 0 9 11 11 7 11 11 1 9 13 2 16 9 15 13 9 9 1 0 0 9 2
26 13 15 2 16 9 13 1 11 16 11 1 0 9 2 13 2 1 9 9 11 2 9 1 0 9 2
25 3 0 13 2 15 9 9 1 9 13 2 13 15 3 9 0 9 11 11 7 10 9 11 11 2
11 13 3 1 9 0 12 2 9 3 13 2
21 9 14 9 0 2 7 3 3 1 0 9 0 9 0 2 15 13 1 0 9 2
14 0 1 15 13 3 15 2 16 1 10 9 3 13 2
34 16 15 13 9 1 9 9 2 15 3 13 1 9 1 12 12 9 9 13 9 0 9 7 0 9 1 2 0 9 1 0 9 2 2
6 13 15 1 10 9 2
17 15 15 14 13 10 9 9 2 1 9 0 9 2 1 10 9 2
25 16 9 13 9 0 13 9 0 9 2 7 7 16 13 0 15 1 9 3 0 9 13 1 9 2
24 16 11 3 13 2 13 15 2 0 9 1 9 11 2 16 15 15 4 13 9 7 0 9 2
6 0 13 7 9 12 2
25 1 15 13 2 0 7 0 9 2 9 1 9 9 1 0 9 7 9 2 15 15 15 3 13 2
38 9 10 9 15 13 9 1 9 2 1 0 1 0 9 0 0 9 9 2 9 2 9 7 9 2 1 10 9 4 13 9 2 15 15 15 3 13 2
26 14 3 1 15 2 1 9 12 13 4 0 9 7 9 9 9 2 9 3 2 1 0 9 9 13 2
13 1 10 9 4 15 9 3 13 1 9 1 9 2
11 9 10 9 13 1 0 2 13 7 0 2
7 13 9 1 9 9 12 2
14 1 0 9 0 9 15 9 13 1 0 9 1 9 2
6 15 13 3 10 9 2
25 10 9 3 13 1 9 9 2 7 13 2 16 9 13 10 0 9 0 9 2 13 2 0 9 2
12 13 2 16 9 13 9 7 9 7 9 9 2
21 9 15 9 13 1 15 2 1 15 4 15 13 9 2 16 4 13 1 15 9 2
10 9 13 15 3 0 2 13 15 15 2
35 13 9 0 0 2 9 9 0 9 11 3 13 2 16 15 15 9 13 2 3 13 13 9 9 1 0 9 2 16 15 0 13 9 9 2
26 1 10 0 9 13 12 9 2 7 13 9 2 7 13 2 7 13 2 16 4 15 9 1 15 13 2
37 1 9 1 9 9 13 2 16 15 13 2 16 4 9 11 13 1 9 0 0 9 0 2 7 9 15 15 3 7 13 2 14 15 9 9 13 2
16 13 7 9 2 16 9 0 15 0 9 4 10 9 3 13 2
3 15 13 2
11 9 13 9 2 7 16 4 9 9 13 2
23 3 3 9 13 2 10 0 9 2 2 16 15 13 0 9 2 15 13 1 9 15 0 2
15 13 13 9 1 9 2 13 1 9 7 1 9 15 13 2
1 9
1 11
2 11 12
2 11 12
1 11
1 12
1 12
6 15 13 1 9 11 2
2 13 4
6 15 13 1 9 11 2
36 9 1 9 9 1 11 13 1 9 2 16 16 0 0 9 11 11 9 11 13 2 9 1 9 9 13 0 9 11 11 7 0 9 11 11 2
27 9 11 7 11 13 1 9 9 1 12 9 0 2 16 13 0 1 11 2 1 15 13 0 9 0 11 2
32 9 15 13 2 3 0 7 0 9 12 0 7 1 15 0 0 9 13 2 16 11 11 13 9 1 3 2 0 9 1 11 2
14 11 2 11 1 0 9 13 1 12 9 7 12 9 2
34 11 2 11 2 15 15 13 0 9 11 2 13 13 9 1 0 9 1 9 2 16 15 11 2 11 13 0 9 2 16 4 13 9 2
31 11 2 11 13 0 9 11 2 11 7 13 2 16 13 1 0 2 14 16 0 9 13 2 16 13 13 13 1 9 11 2
59 11 2 11 15 3 13 2 16 15 13 7 16 11 2 11 1 9 13 1 0 9 2 15 3 13 2 16 4 13 13 1 10 9 1 9 0 9 11 11 2 15 1 1 0 9 1 11 7 0 9 0 0 9 13 13 3 0 9 2
9 9 11 3 13 15 2 15 13 2
14 0 9 1 11 2 11 13 13 2 3 13 9 9 2
8 3 13 7 0 7 11 11 2
24 0 7 0 9 1 0 9 13 12 0 9 7 13 15 2 16 4 13 0 9 1 0 11 2
17 11 2 11 7 15 0 15 13 2 16 4 15 13 13 0 9 2
26 16 9 9 12 0 9 13 2 16 9 13 1 9 2 13 12 0 9 2 1 15 12 13 13 9 2
17 13 7 15 2 16 4 10 9 13 2 7 3 4 1 9 13 2
14 7 3 13 1 10 0 9 2 7 15 15 13 9 2
29 16 13 9 0 9 2 13 13 2 16 13 9 0 9 2 13 1 10 9 1 11 0 9 0 0 9 11 11 2
10 12 2 12 2 12 2 0 0 11 11
2 9 9
2 11 2
10 2 9 12 2 9 12 1 11 2 2
15 9 12 9 13 1 9 9 7 9 2 9 2 12 12 2
25 12 9 1 12 2 2 9 13 1 9 10 9 7 9 2 9 2 12 12 2 9 2 12 12 2
28 12 9 1 12 9 13 1 9 9 2 12 12 2 9 2 12 12 2 9 2 12 12 2 9 2 12 12 2
15 12 9 1 12 9 13 1 15 9 1 9 9 2 12 2
17 12 9 1 12 9 13 1 15 9 1 9 9 2 12 2 12 2
14 12 9 1 12 2 2 9 13 1 9 0 9 12 2
20 12 9 1 12 2 2 9 13 1 9 0 9 12 2 12 2 12 2 12 2
14 12 9 1 12 2 2 9 13 1 9 0 9 12 2
20 12 9 1 12 2 2 9 13 1 9 0 9 12 2 12 2 12 2 12 2
16 12 9 1 12 2 2 9 13 1 9 0 9 12 7 12 2
11 0 9 11 13 12 2 9 12 1 11 2
4 0 9 1 9
6 1 11 15 14 13 3
2 11 2
37 12 9 11 13 13 2 16 15 15 1 9 0 9 13 3 16 3 2 1 12 9 13 9 3 3 0 7 3 9 0 9 13 0 9 1 11 2
14 13 15 1 9 0 9 2 15 3 13 9 0 9 2
29 16 1 9 0 9 1 9 2 16 2 11 13 0 9 2 2 13 14 12 9 0 2 3 1 9 3 12 9 2
31 9 13 10 0 9 15 2 16 0 9 15 3 13 9 1 9 2 7 13 15 10 9 2 16 4 13 3 13 0 9 2
21 1 9 0 1 9 7 0 9 2 7 16 3 0 2 7 3 13 9 1 9 2
27 1 9 1 9 2 16 2 9 13 0 9 2 2 3 13 12 9 0 7 2 3 13 2 12 9 0 2
10 14 12 9 9 9 10 9 3 13 2
5 0 9 9 13 13
2 11 2
2 11 2
5 0 9 9 13 13
2 11 2
38 16 9 0 9 11 11 7 3 16 9 0 9 9 1 11 4 13 9 0 9 0 9 11 7 9 10 0 9 11 2 11 2 0 7 1 0 9 2
23 11 4 13 9 9 9 0 9 11 11 11 2 0 1 9 2 9 2 9 7 0 9 2
13 11 4 13 1 0 9 0 0 9 1 9 0 2
13 13 15 9 11 7 11 9 1 9 1 0 9 2
1 9
13 13 15 9 11 7 11 9 1 9 1 0 9 2
5 9 9 13 7 11
27 2 1 11 7 11 13 14 10 9 16 1 0 9 7 0 9 2 2 13 11 11 1 0 9 1 11 2
27 13 2 14 15 13 2 16 11 11 16 9 3 13 0 9 1 0 9 2 13 15 1 15 1 9 9 2
10 11 13 1 9 3 13 10 0 9 2
13 10 9 15 3 13 9 1 9 0 2 0 9 2
40 16 9 1 11 11 7 0 0 2 0 9 13 3 1 12 9 3 2 7 15 3 14 1 0 9 11 2 1 9 1 11 7 11 4 13 13 3 0 9 2
21 11 13 1 0 0 9 0 9 2 16 13 9 0 9 1 0 0 9 1 11 2
16 3 13 9 1 11 7 11 3 1 10 9 9 9 3 13 2
12 3 13 0 9 1 0 9 2 1 9 0 2
14 10 9 1 11 7 11 13 0 1 0 9 1 9 2
18 0 9 1 9 7 11 11 2 16 1 15 3 13 2 3 13 13 2
21 16 15 11 1 11 13 13 2 13 3 1 9 2 16 4 13 13 1 0 9 2
20 9 9 1 12 9 13 1 9 1 11 2 15 11 13 1 9 1 9 12 2
10 11 13 1 10 9 3 3 1 9 2
15 9 11 13 0 9 3 3 0 9 2 16 13 15 3 2
31 13 3 2 16 10 0 9 13 1 9 0 9 1 11 14 1 0 0 9 2 1 15 3 13 0 9 0 9 0 9 2
9 11 11 0 9 1 9 3 13 2
17 3 0 9 9 1 10 9 1 12 9 7 13 1 0 0 9 2
18 0 9 1 0 9 3 13 13 2 16 13 9 11 1 11 1 9 2
15 13 7 3 0 9 7 13 2 16 10 9 3 13 9 2
29 1 0 9 9 0 9 1 11 13 0 0 9 11 11 2 1 9 3 2 7 0 9 11 11 11 11 2 3 2
21 9 7 9 2 15 13 13 1 12 1 12 0 9 1 9 0 0 0 9 11 2
17 13 1 9 1 9 2 3 9 1 9 9 13 0 0 9 11 2
7 0 9 11 9 9 0 9
2 11 2
23 11 3 13 2 0 9 2 1 11 2 16 15 1 0 9 13 1 10 9 15 0 9 2
27 0 0 9 15 13 13 0 0 9 2 16 4 13 1 11 15 0 0 0 9 2 13 9 9 11 11 2
23 9 1 11 13 1 15 2 16 7 0 9 0 0 9 1 9 1 9 1 11 15 13 2
24 1 0 9 1 9 9 11 13 0 9 1 0 9 2 0 0 9 7 9 9 0 0 9 2
3 9 15 13
5 11 2 11 2 2
30 1 0 9 0 9 11 1 0 11 13 0 9 9 11 11 9 1 15 2 16 10 9 11 11 13 1 9 1 9 2
31 9 13 2 16 15 3 13 11 2 11 13 1 9 10 9 7 16 15 13 3 3 2 16 10 9 1 9 13 0 9 2
22 9 11 3 15 3 3 13 1 11 2 11 2 15 13 2 16 15 2 9 13 2 2
15 1 10 9 9 1 9 2 15 9 9 13 9 2 13 2
14 13 2 16 11 2 11 13 0 9 0 1 12 9 2
32 1 9 1 9 3 13 2 16 15 2 13 13 1 9 2 15 3 0 9 13 2 7 13 15 15 2 3 10 9 13 2 2
28 1 10 9 1 0 9 4 13 9 11 1 9 13 9 7 1 0 0 9 9 2 7 13 1 10 0 9 2
12 1 11 7 11 3 13 0 9 13 12 0 9
2 11 2
21 1 0 9 11 7 11 4 1 9 13 12 0 0 9 0 9 11 2 9 2 2
10 1 3 9 11 7 11 3 13 9 2
22 0 9 15 1 0 9 3 13 1 0 9 9 1 11 7 1 9 11 1 0 11 2
9 0 9 13 1 11 0 0 9 2
14 0 7 0 9 7 3 13 1 0 9 9 0 9 2
15 0 9 13 2 16 0 9 13 1 11 13 1 12 9 2
27 9 11 7 11 7 11 1 9 1 9 1 9 11 13 2 16 15 13 13 0 9 1 9 9 1 11 2
43 9 0 9 1 11 11 11 7 9 11 15 13 2 16 3 13 11 0 0 9 0 11 2 16 4 3 7 1 9 13 0 9 2 15 13 2 9 0 9 0 9 2 2
7 11 7 9 15 13 1 9
2 11 2
17 11 7 9 15 13 1 9 0 9 9 0 0 9 1 0 9 2
30 9 1 9 1 9 0 9 1 9 1 11 11 2 11 13 2 16 11 13 1 9 10 9 1 9 0 0 9 11 2
18 0 2 0 9 1 9 9 0 0 9 13 1 9 1 0 9 11 2
7 11 2 1 2 11 0 9
2 11 2
18 0 0 9 11 2 1 2 11 4 13 1 0 0 9 9 0 9 2
17 0 9 11 2 1 2 11 4 13 0 9 1 0 9 3 3 2
7 1 9 9 13 0 9 2
24 1 9 13 9 1 10 0 9 1 0 9 9 1 9 11 2 11 2 11 2 12 2 9 2
10 9 9 4 13 1 3 16 12 9 2
6 9 9 9 1 11 2
2 11 2
33 0 9 2 15 13 1 9 1 11 2 3 13 13 9 1 9 9 0 9 1 0 2 11 2 16 15 3 0 9 13 0 9 2
24 0 9 3 13 2 16 1 0 9 9 2 3 15 9 13 2 13 13 9 2 15 13 13 2
5 9 9 9 13 2
11 0 0 9 3 13 2 16 9 3 13 2
4 0 0 9 13
2 11 2
35 9 2 15 1 9 13 1 0 9 11 0 9 0 9 1 9 1 9 10 9 11 11 2 3 13 10 9 2 15 4 1 9 9 13 2
16 0 9 1 0 9 11 2 12 9 3 1 11 2 3 13 2
15 1 12 9 9 1 9 13 13 7 3 9 9 3 13 2
10 9 0 7 0 11 1 11 1 0 9
2 11 2
36 0 9 13 13 0 7 1 9 9 1 0 9 2 7 10 9 13 13 9 0 0 9 2 13 3 1 0 9 0 9 0 9 9 11 11 2
17 13 2 16 0 9 0 9 11 15 13 12 2 9 1 0 11 2
22 13 15 1 9 0 9 1 0 9 7 11 7 1 0 9 1 9 0 7 0 11 2
27 13 2 16 0 9 15 13 1 9 0 9 2 16 11 2 15 15 1 0 9 13 2 13 10 0 9 2
14 13 9 0 9 2 15 13 1 9 1 0 9 9 2
21 1 0 9 0 9 0 9 13 0 9 2 0 9 2 0 9 7 0 0 9 2
15 1 9 9 7 0 0 9 13 11 9 1 0 0 9 2
8 10 9 1 2 0 2 11 2
2 11 2
42 9 0 9 11 11 3 13 9 2 16 11 11 7 0 9 11 11 1 10 0 9 13 9 0 2 0 2 11 2 15 4 13 13 0 9 2 10 9 13 0 9 2
16 9 11 11 13 10 9 0 1 9 0 11 1 0 7 0 2
9 3 10 9 3 13 9 0 9 2
39 0 11 1 9 1 0 9 1 11 13 2 16 1 10 0 9 1 11 15 11 7 11 13 13 9 11 2 11 7 9 9 2 11 2 11 7 11 2 2
15 9 10 9 13 1 9 9 1 0 9 1 11 7 11 2
27 2 11 2 11 7 9 9 4 16 3 0 9 0 9 13 1 10 9 13 0 7 0 9 1 9 12 2
21 0 9 4 13 9 13 1 10 9 2 16 15 1 15 4 13 2 2 13 9 2
8 9 0 9 0 9 11 7 11
2 11 2
21 1 9 9 9 7 9 9 0 1 11 13 3 1 11 0 9 0 9 0 9 2
18 9 15 1 0 13 0 0 9 11 2 11 7 0 9 11 2 11 2
25 9 15 13 1 9 0 9 9 9 11 2 11 2 13 0 9 11 11 2 15 9 13 1 11 2
16 12 1 0 9 13 9 1 0 9 2 0 9 7 0 9 2
24 1 11 15 1 1 0 9 9 13 3 1 15 2 10 9 13 1 12 1 10 9 2 11 2
18 2 13 15 15 2 7 9 2 2 13 0 9 11 2 9 2 12 2
10 11 13 9 1 11 9 9 11 7 11
2 11 2
39 0 9 0 9 1 9 2 9 7 9 7 0 9 0 9 1 9 0 2 2 0 9 13 9 0 9 0 9 11 11 1 9 0 9 11 11 1 11 2
16 11 13 1 15 9 1 0 11 2 13 1 9 9 11 11 2
12 13 9 0 9 2 1 15 15 1 9 13 2
17 1 0 13 9 1 11 7 13 9 12 9 13 1 10 9 9 2
11 1 11 0 9 4 13 0 9 1 11 2
1 3
2 13 9
30 1 9 9 9 9 2 11 2 1 9 13 9 9 9 2 0 15 0 9 0 9 2 15 4 13 0 9 7 9 2
14 13 1 0 9 11 7 11 2 13 9 9 11 11 2
2 11 2
1 0
27 9 9 1 11 1 0 0 9 1 11 2 15 13 9 0 9 11 2 4 0 2 9 11 13 1 9 2
6 13 15 1 9 11 2
2 0 9
14 0 9 0 0 0 9 1 9 11 13 3 1 11 2
18 1 9 9 15 13 0 7 0 9 2 15 4 13 3 11 2 11 2
3 11 3 13
39 11 2 11 15 3 13 1 0 9 2 13 9 0 9 11 2 11 1 9 1 9 9 11 11 2 11 2 11 2 2 16 11 13 9 0 9 1 11 2
4 11 1 0 9
36 9 9 11 11 2 11 13 2 16 1 9 0 9 2 11 2 11 13 0 9 2 7 15 1 9 2 16 9 0 9 11 13 9 0 9 2
9 9 9 11 11 0 9 1 0 11
2 11 2
20 1 9 9 0 9 1 9 0 9 11 11 13 3 3 11 11 2 12 2 2
35 1 0 9 15 13 1 0 9 0 0 9 1 15 2 16 13 9 1 9 9 12 1 0 9 9 1 9 11 2 15 10 9 13 9 2
20 1 9 0 1 9 9 13 9 13 9 7 9 2 15 4 15 13 3 13 2
9 9 7 13 2 16 13 0 9 2
27 1 9 1 11 15 13 1 15 2 16 4 1 9 9 13 9 0 9 2 15 13 10 0 9 0 9 2
22 9 11 11 13 1 9 2 3 12 1 0 9 13 0 0 9 1 9 11 1 11 2
9 11 11 13 0 7 13 12 9 2
17 13 0 1 9 0 9 0 1 0 0 9 2 15 13 1 9 2
5 0 9 13 11 13
10 11 13 9 2 15 15 13 1 9 2
27 9 10 9 13 1 10 9 3 0 2 13 9 13 9 0 3 2 16 9 9 13 10 9 12 0 9 2
16 1 0 9 15 13 3 12 2 12 2 9 7 12 2 9 2
25 12 2 16 3 3 7 3 2 13 1 0 11 2 3 1 9 11 1 0 0 9 2 9 2 2
31 1 0 9 15 4 13 1 15 2 16 13 10 0 9 13 12 9 0 9 1 9 0 9 1 9 0 2 11 7 11 2
54 0 0 9 3 3 13 13 9 0 9 1 9 2 15 13 13 9 1 9 1 0 9 2 11 2 2 3 7 13 0 9 9 2 1 9 2 13 9 1 9 1 11 2 7 1 9 1 9 13 0 0 9 2 2
14 1 9 1 11 3 11 13 2 16 13 10 0 9 2
27 1 9 12 7 12 2 3 4 15 11 13 2 3 2 13 9 11 2 4 0 9 3 13 4 3 13 2
19 9 2 12 1 9 0 11 7 0 1 11 2 4 7 0 9 3 13 2
27 1 0 9 4 15 3 13 13 0 13 1 15 9 2 3 16 0 9 1 0 9 13 9 12 9 9 2
30 0 9 13 7 0 2 11 3 3 13 2 16 1 11 3 13 2 7 16 7 3 13 0 13 0 9 7 13 11 2
26 9 15 3 1 9 13 2 1 0 9 7 13 0 9 1 9 9 0 7 0 9 2 15 9 13 2
29 0 9 13 3 3 1 9 1 9 1 0 0 9 9 1 9 1 15 2 16 15 13 1 9 1 0 0 9 2
16 3 3 4 0 9 2 16 13 2 7 13 2 3 13 9 2
14 15 15 4 13 12 2 9 2 7 9 3 13 0 2
23 16 4 3 11 9 1 9 13 2 13 4 15 14 1 0 9 9 3 16 12 0 9 2
27 9 2 15 13 1 0 11 2 4 15 3 13 13 7 0 9 7 9 2 15 4 13 3 1 10 9 2
30 14 3 3 2 11 4 1 0 9 13 7 1 10 9 13 15 1 9 9 7 4 15 3 13 13 1 10 0 9 2
54 7 16 9 9 13 1 15 2 16 0 11 13 3 3 13 0 9 1 9 0 11 2 15 4 3 13 1 9 1 11 7 11 13 12 1 12 9 0 9 2 13 9 0 11 9 2 15 13 1 9 11 3 0 2
32 13 15 2 16 11 2 9 0 10 0 9 1 9 9 2 4 13 13 10 9 9 9 1 15 9 0 7 3 7 0 11 2
21 3 13 10 0 9 14 14 0 9 7 1 0 9 4 15 1 10 9 14 13 2
35 1 0 9 7 13 1 9 1 0 9 1 12 9 2 12 9 3 2 2 7 0 0 9 1 9 0 13 3 4 3 2 13 9 2 2
27 0 9 13 7 9 7 0 9 2 10 0 2 7 3 0 9 4 14 14 3 13 1 9 1 0 9 2
32 7 3 16 11 7 11 13 3 7 11 9 2 16 4 10 9 2 9 9 7 9 9 2 13 13 9 7 10 0 0 9 2
22 0 9 13 7 7 9 1 15 2 16 4 15 9 0 9 13 1 9 13 10 9 2
45 13 7 9 2 16 1 9 2 15 3 3 12 9 13 3 0 7 0 9 2 13 11 3 0 9 7 1 9 1 15 13 3 3 3 9 16 10 10 9 2 15 13 9 11 2
15 1 0 9 9 15 7 9 13 10 9 0 9 7 9 2
31 11 11 1 10 9 13 2 16 1 10 9 1 9 13 16 2 9 2 15 15 13 13 1 9 2 7 13 3 0 2 2
27 7 1 3 0 9 2 3 1 9 2 11 14 2 7 14 2 2 4 9 11 13 9 7 1 0 9 2
7 0 9 11 13 9 1 11
11 10 9 13 0 0 9 1 0 10 9 2
16 9 11 11 15 3 13 1 0 9 9 7 1 15 3 13 2
9 13 15 16 0 11 13 10 9 2
8 1 11 13 3 10 0 9 2
9 10 9 13 10 9 1 0 9 2
9 13 0 2 7 9 11 13 13 2
11 7 15 1 9 2 15 13 9 0 9 2
3 15 13 2
5 15 3 13 13 2
15 13 3 2 1 9 7 1 10 9 2 1 9 10 9 2
4 13 15 15 2
14 15 4 15 3 10 9 13 3 2 15 4 15 13 2
11 3 12 9 13 1 0 9 11 1 9 2
15 3 13 0 7 0 9 2 15 0 13 7 3 15 0 2
8 13 4 15 9 11 13 3 2
13 16 15 15 3 13 2 15 15 13 13 0 9 2
8 13 15 15 1 10 0 9 2
13 11 4 15 13 3 3 2 15 13 15 3 0 2
23 13 3 3 9 2 16 4 15 9 2 0 9 7 9 13 3 1 10 9 13 7 13 2
17 13 2 16 9 2 15 13 0 9 0 9 2 13 13 1 9 2
31 16 4 7 1 12 9 13 10 0 9 2 13 4 15 9 1 9 7 13 4 9 2 16 4 1 10 9 9 15 13 2
16 3 3 13 1 9 9 10 9 2 7 13 3 3 1 9 2
16 1 9 10 9 13 1 10 9 9 0 9 1 9 0 9 2
24 16 2 9 0 9 2 2 15 4 13 1 0 9 1 11 2 15 15 3 13 13 7 13 2
19 9 1 11 15 13 14 3 2 16 4 15 1 15 13 1 9 0 9 2
17 13 3 1 0 0 9 1 10 9 7 1 10 9 2 1 9 2
18 0 9 13 3 9 2 16 0 9 3 13 2 16 0 9 3 13 2
27 13 15 0 9 11 2 16 1 9 1 11 13 2 2 13 13 14 0 9 2 7 7 0 0 9 2 2
18 11 11 13 12 0 9 2 7 3 15 2 16 13 3 3 0 9 2
17 3 1 15 13 9 0 9 2 16 4 13 9 1 9 0 9 2
5 13 1 15 0 2
18 1 15 4 15 13 3 13 1 9 15 9 7 3 3 1 0 9 2
14 13 15 11 11 1 11 2 9 15 7 13 16 11 2
17 15 1 15 3 13 1 0 9 2 16 16 4 13 1 15 0 2
12 1 15 3 3 13 2 1 11 7 1 11 2
6 3 2 16 1 11 2
10 15 13 0 2 1 11 14 1 11 2
10 11 13 0 16 0 2 11 7 9 2
9 11 3 13 2 7 11 13 0 2
9 13 9 0 9 15 9 3 9 2
3 6 14 2
20 13 3 1 9 11 11 2 1 15 4 3 13 7 3 13 3 9 10 9 2
29 3 15 13 7 3 15 0 9 13 2 3 2 3 13 15 2 4 13 13 0 9 2 15 13 7 1 12 9 2
7 7 3 13 3 16 0 2
16 13 4 12 9 9 9 7 0 9 2 13 9 7 16 9 2
10 13 3 10 9 2 15 4 13 13 2
13 13 3 0 1 15 2 16 4 13 1 0 9 2
12 10 0 9 13 12 9 2 13 15 16 9 2
10 3 13 15 3 3 13 1 10 9 2
8 13 15 3 3 9 16 11 2
10 3 14 2 16 10 9 3 13 9 2
7 9 0 9 11 13 9 9
23 9 0 11 1 9 0 9 2 11 2 4 13 15 2 16 11 3 13 9 2 15 13 2
25 7 9 11 7 11 13 0 9 1 9 1 11 2 16 15 11 13 9 0 9 2 13 0 9 2
18 0 9 13 15 2 1 10 9 13 9 9 13 1 0 9 11 11 2
15 9 9 0 9 3 13 9 9 2 15 4 3 13 3 2
18 3 4 10 9 13 1 0 9 2 0 9 2 7 15 1 9 9 2
21 15 0 0 9 1 0 11 1 9 11 13 4 1 9 11 2 15 9 3 13 2
23 0 0 0 9 1 9 9 13 9 0 9 11 11 2 16 4 9 11 13 9 0 9 2
22 13 4 0 13 1 0 11 1 0 9 2 15 4 13 13 1 10 9 9 0 9 2
12 9 11 13 2 16 10 9 13 13 3 9 2
25 7 13 15 3 9 2 15 4 13 0 9 13 2 16 15 7 3 13 13 11 1 9 7 11 2
3 0 9 9
1 9
3 0 9 9
33 16 13 1 9 12 1 0 9 0 9 0 0 9 9 11 2 13 15 13 10 9 11 2 16 4 15 13 9 1 9 7 9 2
15 3 13 1 9 12 9 7 10 9 13 12 9 1 9 2
25 11 15 3 10 9 14 13 2 15 4 7 3 1 9 9 0 0 9 13 1 9 12 2 12 2
19 7 1 9 9 3 13 0 9 1 9 7 9 13 2 13 15 1 9 2
14 11 15 3 13 9 9 2 15 15 11 13 3 3 2
15 7 11 3 13 1 9 16 12 1 9 0 9 2 2 2
3 7 9 2
23 16 1 0 9 15 13 9 0 9 1 9 13 16 0 9 2 3 13 3 1 0 9 2
31 9 9 15 9 13 1 11 7 1 9 0 9 0 11 3 1 9 9 2 3 15 13 12 7 1 0 9 3 12 9 2
30 1 1 15 2 16 3 0 9 15 9 13 1 12 9 2 13 15 2 16 15 1 12 9 0 9 13 3 1 12 2
12 9 15 3 13 1 12 1 12 0 0 9 2
8 3 11 3 13 0 0 9 2
21 1 15 13 15 3 0 2 0 9 12 1 12 15 10 9 13 1 12 1 12 2
17 13 1 9 1 9 0 9 2 9 0 9 0 9 9 3 13 2
12 7 13 9 2 16 15 10 9 3 13 13 2
7 1 0 9 15 3 13 2
4 9 9 13 0
2 11 2
4 9 9 13 0
2 11 2
12 3 1 11 13 9 1 0 0 7 0 9 2
26 9 13 2 16 0 9 0 9 4 13 13 14 12 9 2 15 7 4 13 1 9 9 1 0 9 2
13 1 0 9 13 1 12 9 0 0 9 0 9 2
11 0 9 0 9 13 13 1 12 9 9 2
17 15 1 0 12 9 2 15 15 9 13 2 4 13 13 12 9 2
5 12 0 9 15 13
2 11 2
44 1 9 4 3 13 12 0 0 9 2 9 9 1 0 9 11 7 11 2 15 13 10 9 1 0 9 2 7 9 9 1 0 9 2 9 1 11 7 11 2 0 0 9 2
7 9 15 13 1 10 9 2
6 11 11 13 3 1 9
2 11 2
14 0 9 11 11 2 9 0 9 2 13 3 3 0 2
11 11 4 3 13 1 12 9 1 0 11 2
6 9 9 3 13 0 2
6 1 9 13 9 9 13
5 11 2 11 2 2
17 9 0 9 13 9 13 9 9 2 16 15 0 9 13 13 9 2
21 9 0 9 7 13 9 10 9 1 9 1 9 0 9 13 7 13 15 9 13 2
20 9 15 3 1 9 13 3 1 10 9 2 15 13 1 10 10 9 3 13 2
8 13 15 15 9 9 11 11 2
31 9 9 3 13 9 1 9 0 9 0 9 3 15 2 16 1 15 3 13 0 9 2 15 4 15 13 13 1 0 9 2
20 15 1 9 7 1 10 0 9 13 0 0 0 9 1 9 0 9 1 9 2
11 13 15 15 9 0 9 9 9 11 11 2
10 0 9 13 1 0 9 7 9 9 2
15 1 9 1 0 9 13 1 0 9 9 10 0 0 9 2
11 9 13 7 0 13 9 1 9 0 9 2
14 15 13 9 9 2 15 13 9 3 0 7 0 9 2
18 9 0 7 0 9 13 3 1 9 3 0 0 9 9 9 7 9 2
29 0 9 13 2 16 4 1 0 9 0 9 1 9 9 4 13 0 9 9 9 0 1 9 0 9 1 0 9 2
7 9 13 16 9 2 13 11
5 11 2 11 2 2
18 1 10 9 14 13 1 9 9 1 0 9 1 9 1 0 9 9 2
13 13 13 1 0 9 2 9 15 0 9 7 3 2
19 13 15 3 1 9 1 2 9 0 9 9 2 9 11 11 2 11 2 2
28 1 15 15 0 9 2 15 3 0 9 13 1 9 2 13 7 9 7 0 9 2 1 15 15 13 0 9 2
17 3 1 9 13 2 16 10 9 13 0 9 7 9 2 13 11 2
18 9 13 0 9 2 10 9 4 13 13 0 0 2 0 7 0 9 2
13 0 9 4 9 13 4 1 11 1 0 9 13 2
6 9 13 7 9 11 2
8 13 15 13 16 0 0 9 2
15 0 9 13 7 0 9 11 2 15 15 9 13 3 13 2
47 15 0 9 3 3 3 1 10 9 1 0 9 13 2 16 3 13 9 2 16 4 1 9 10 9 7 9 13 15 7 2 15 0 2 1 0 9 3 10 9 2 15 15 13 0 9 2
5 9 9 1 9 12
5 11 2 11 2 2
20 9 2 9 7 9 9 0 9 13 1 0 9 3 13 1 12 2 9 12 2
17 3 1 9 0 9 13 13 9 9 2 1 15 13 10 9 13 2
16 9 9 0 9 13 13 9 9 9 9 2 15 3 13 9 2
19 0 1 9 0 0 9 2 0 2 9 2 4 13 1 12 2 9 12 2
9 1 9 13 12 9 1 0 9 2
8 1 9 13 11 13 0 9 2
19 9 0 9 4 13 4 3 13 9 2 9 13 9 0 0 9 9 2 2
16 9 7 9 13 3 0 13 1 0 9 9 0 9 12 9 2
10 9 1 9 9 13 12 7 12 9 2
12 9 9 11 13 9 1 9 9 1 10 9 2
23 13 2 16 1 9 9 13 1 9 1 12 12 0 9 1 9 1 12 7 12 9 9 2
37 9 11 11 2 11 2 2 12 1 9 9 2 15 1 9 1 9 11 13 2 16 1 9 9 13 0 13 1 9 10 9 12 9 7 0 9 2
11 0 9 16 9 13 7 9 9 0 9 2
19 1 11 10 9 13 3 9 1 9 9 2 15 13 4 13 1 9 12 2
19 9 13 2 16 9 0 9 1 9 15 10 9 13 14 1 14 12 9 2
12 0 9 13 9 1 12 7 12 9 2 13 2
11 11 2 0 0 9 1 11 1 12 2 9
7 11 2 11 2 11 2 2
15 0 0 9 1 9 1 11 13 0 9 1 12 2 9 2
24 9 9 11 11 3 13 2 16 0 9 1 9 13 13 2 16 3 15 0 9 13 7 13 2
21 11 13 2 16 1 0 9 9 4 13 0 9 2 0 12 9 0 9 1 9 2
16 0 9 1 0 9 4 13 9 9 1 0 9 7 0 9 2
23 3 4 13 2 16 13 0 13 0 9 7 16 13 9 1 9 1 10 9 2 13 11 2
28 0 2 0 0 9 2 15 13 1 11 2 3 13 9 2 15 13 9 0 9 0 9 1 9 0 9 11 2
20 9 0 9 1 9 11 11 13 2 16 12 9 4 3 13 0 9 1 9 2
12 1 0 0 9 13 11 3 0 9 7 11 2
24 9 9 0 9 1 9 11 11 15 13 2 16 0 9 4 15 13 13 1 12 7 12 9 2
10 9 13 14 1 12 9 9 9 9 2
1 11
16 1 9 2 15 13 1 9 2 13 9 2 15 13 15 1 9
5 9 0 7 0 9
7 15 15 13 1 9 9 2
7 9 13 9 0 9 1 0
7 11 2 11 2 11 2 2
16 9 9 13 1 9 9 9 0 9 1 0 2 16 13 0 2
20 3 3 9 0 13 0 9 1 0 7 0 7 3 3 0 7 0 16 0 2
14 0 9 4 13 1 0 2 14 16 13 1 10 9 2
16 13 15 1 9 9 1 9 0 9 1 0 0 9 0 9 2
27 9 15 13 13 2 15 15 9 13 1 9 9 7 10 9 3 13 9 2 16 13 1 0 7 0 9 2
27 1 3 15 9 2 12 9 2 13 0 9 9 7 16 3 0 15 13 7 10 9 2 1 12 9 9 2
20 0 9 15 13 1 0 9 9 2 7 16 7 15 13 1 9 12 12 9 2
10 0 9 9 13 0 1 12 9 0 2
15 3 12 12 9 15 13 2 16 13 1 0 7 0 9 2
25 1 1 15 2 16 0 1 9 13 9 7 9 9 2 13 13 2 16 9 13 9 3 0 9 2
15 9 1 9 0 9 3 13 3 0 2 13 1 15 11 2
5 9 1 9 1 11
2 11 2
24 9 0 9 0 9 1 0 9 0 9 9 11 11 1 11 1 9 11 15 4 13 0 9 2
23 9 9 15 13 9 1 9 7 9 9 1 10 9 7 3 15 13 13 7 15 9 11 2
21 9 9 0 9 1 11 11 11 3 13 2 16 0 9 3 13 1 9 0 9 2
19 1 15 15 7 13 0 9 0 11 2 1 10 9 4 9 9 13 13 2
14 1 9 1 9 2 13 1 9 2 2 13 11 11 2
25 1 11 11 1 0 9 0 11 13 9 0 9 1 9 1 9 9 2 15 15 1 10 9 13 2
11 1 9 4 9 13 0 9 1 0 9 2
14 9 4 13 3 1 15 13 9 9 1 9 0 9 2
32 9 13 0 9 1 0 9 2 15 4 13 9 1 0 9 2 0 1 9 1 9 1 9 14 1 9 7 3 1 0 9 2
14 3 3 15 0 9 1 11 3 13 0 0 0 9 2
16 0 9 15 13 1 11 1 9 0 9 7 13 15 0 9 2
11 9 1 0 9 1 11 3 1 9 9 13
6 9 15 3 13 14 13
5 11 2 11 2 2
11 9 0 9 0 9 13 2 13 9 9 2
26 3 7 9 9 9 9 9 11 11 13 2 16 1 9 0 9 15 15 1 9 13 1 0 9 13 2
17 0 0 9 13 4 13 1 9 0 9 2 15 3 13 0 9 2
20 9 13 13 0 9 2 13 9 9 7 13 9 2 7 15 1 0 9 9 2
18 0 9 13 13 9 2 9 15 13 1 0 9 7 0 9 9 13 2
17 11 11 13 2 16 9 9 13 9 9 9 0 9 0 1 9 2
38 10 9 13 3 12 2 1 11 1 11 1 11 1 9 12 9 2 0 9 1 11 1 11 1 11 7 0 9 1 0 11 1 0 11 0 12 9 2
10 1 9 15 10 9 13 1 11 9 2
17 2 3 15 9 13 2 16 9 3 4 13 2 2 13 9 11 2
28 1 15 13 9 1 0 12 9 13 2 3 4 0 9 1 9 13 7 3 1 0 9 13 0 9 0 9 2
10 3 4 15 7 9 13 13 0 9 2
17 10 9 15 13 2 16 9 4 13 14 13 9 7 4 13 9 2
26 1 11 11 0 9 13 1 9 0 9 13 2 16 13 13 7 13 9 2 13 9 7 9 0 9 2
4 11 13 13 9
5 11 2 11 2 2
12 0 9 15 7 1 9 13 13 0 0 9 2
11 9 9 7 13 9 0 9 1 9 9 2
16 9 3 13 1 9 9 2 3 9 0 9 13 0 0 9 2
25 1 0 9 9 11 11 4 0 9 1 12 9 13 3 1 12 9 9 2 3 3 4 13 9 2
16 16 15 9 4 13 2 13 1 9 1 0 9 7 0 9 2
7 9 4 13 13 1 9 2
8 9 13 1 9 12 9 9 2
15 1 0 0 9 4 15 1 1 9 1 9 9 13 13 2
11 9 4 3 13 1 9 9 1 0 9 2
12 1 11 11 4 15 9 13 13 1 12 9 2
6 9 0 9 13 13 3
5 11 2 11 2 2
11 9 0 9 13 1 9 10 9 0 9 2
10 3 9 13 16 9 9 0 9 12 2
15 1 10 9 13 12 9 2 16 3 13 3 12 9 9 2
25 9 0 9 2 15 1 9 9 13 3 1 9 2 13 2 16 15 15 3 13 9 9 0 9 2
22 1 9 13 7 3 13 9 1 3 0 2 15 4 1 0 9 9 13 1 0 9 2
12 9 3 0 7 9 9 4 13 1 0 9 2
11 9 9 13 9 2 9 9 13 0 9 2
22 12 9 1 0 9 12 9 13 0 9 11 2 11 2 0 0 9 1 11 7 11 2
13 1 9 9 4 3 13 12 9 1 9 0 9 2
14 1 9 0 9 11 11 4 9 0 9 3 13 9 2
25 9 13 1 9 0 9 10 9 1 9 9 13 0 9 7 9 9 2 13 7 0 9 9 13 2
16 9 3 13 1 9 15 12 9 2 15 13 1 9 0 9 2
5 9 3 13 9 9
4 9 4 13 9
7 1 11 13 9 9 1 9
2 11 2
15 0 0 9 0 9 1 9 0 11 13 1 0 9 11 2
17 0 9 1 9 4 13 9 2 15 13 9 13 0 9 1 0 2
12 9 1 0 9 13 1 9 1 0 9 0 2
18 0 9 9 13 1 9 9 9 0 9 9 7 9 2 15 13 9 2
7 15 13 9 1 10 9 2
16 9 9 1 15 13 9 3 0 2 16 4 15 13 13 9 2
23 9 13 15 0 9 2 13 7 0 9 7 3 13 9 9 2 1 15 15 0 9 13 2
14 1 0 9 0 9 1 9 3 4 13 12 9 9 2
14 9 4 13 7 1 9 2 16 9 13 3 1 9 2
29 1 11 13 0 9 1 12 9 2 1 0 9 15 13 16 0 13 0 9 1 11 1 11 7 3 11 1 11 2
19 9 0 9 13 1 10 9 9 0 9 7 13 3 9 1 11 7 11 2
15 9 13 13 3 3 0 9 11 0 9 1 3 0 9 2
6 2 9 13 9 9 2
5 1 9 14 9 11
5 11 2 11 2 2
33 0 9 0 9 15 4 13 13 14 9 11 2 15 13 1 10 9 0 9 7 13 3 1 0 9 9 1 9 0 9 12 9 2
10 13 1 15 9 2 15 13 0 9 2
16 0 9 4 13 13 9 2 9 7 9 9 0 1 0 9 2
31 0 0 9 2 1 15 13 4 0 9 3 13 2 7 13 2 13 2 16 3 0 0 9 13 0 1 10 9 3 13 2
3 9 13 0
5 11 2 11 2 2
13 9 3 13 9 12 0 0 0 0 9 1 11 2
24 0 9 1 10 0 9 1 9 2 9 7 9 13 1 9 3 1 9 9 9 9 9 11 2
22 0 2 15 1 0 9 13 2 9 13 0 9 1 9 7 13 15 3 1 9 9 2
14 1 9 13 7 0 11 12 2 7 9 13 1 9 2
15 12 0 9 13 0 12 2 9 0 0 9 1 0 11 2
5 9 1 9 1 9
5 11 2 11 2 2
25 1 9 0 0 9 4 3 13 0 9 1 0 0 9 1 9 7 0 9 1 11 7 1 11 2
16 9 4 13 0 9 2 16 3 1 0 9 13 13 0 9 2
16 9 9 0 9 4 13 13 9 9 9 7 12 9 3 9 2
33 1 9 13 0 15 13 1 12 2 9 1 0 9 9 9 2 11 1 0 9 12 1 11 7 1 11 1 0 9 12 1 11 2
22 1 0 9 4 9 13 1 9 0 0 9 1 0 9 2 1 11 1 11 1 0 2
24 9 9 7 9 4 13 0 9 0 1 0 9 2 1 0 9 15 13 1 0 7 0 9 2
6 0 9 3 13 13 9
2 11 2
19 13 3 16 0 2 16 10 0 9 7 9 13 9 0 9 1 9 9 2
19 13 15 3 9 9 9 0 9 7 0 9 1 11 2 11 2 11 11 2
13 0 9 13 1 15 0 9 0 9 2 3 0 2
27 9 0 9 3 13 0 9 13 1 15 0 9 2 16 9 4 13 13 1 10 9 3 14 1 9 9 2
7 0 9 14 4 1 11 13
5 11 2 11 2 2
30 9 0 1 0 11 1 11 2 1 15 0 9 13 9 1 9 1 9 7 9 2 4 1 0 9 13 3 1 11 2
10 13 15 3 9 0 0 9 11 11 2
7 13 15 1 12 0 9 2
16 1 11 4 1 11 1 0 9 1 0 9 13 3 12 9 2
25 9 1 9 7 9 13 1 9 11 13 7 0 9 15 13 9 15 2 16 3 13 9 0 9 2
17 0 9 13 1 9 10 9 1 9 9 13 2 7 13 1 11 2
34 1 9 13 7 9 0 9 9 15 0 9 1 11 2 15 13 12 2 9 11 11 9 0 9 9 9 0 11 11 2 11 2 11 2
34 13 1 15 3 2 16 12 9 3 13 9 9 1 9 7 9 2 7 0 13 7 13 13 2 16 15 4 1 9 7 9 3 13 2
12 9 1 10 9 13 3 13 7 1 0 9 2
17 9 4 13 1 9 9 11 11 2 15 15 1 11 1 11 13 2
9 0 9 0 1 12 2 12 2 12
2 9 9
8 9 9 9 9 9 9 9 9
13 11 9 2 2 12 9 2 1 0 2 9 11 2
4 15 1 12 9
6 9 12 2 12 2 12
1 9
1 9
1 9
3 11 12 12
4 0 9 12 12
3 11 12 12
4 0 9 12 12
4 0 9 12 12
8 0 9 1 9 2 0 1 9
7 11 2 11 2 11 2 2
22 1 11 13 1 9 9 9 0 7 11 1 9 14 1 12 9 0 16 1 0 9 2
20 11 2 15 3 13 1 11 12 9 2 15 1 11 13 1 12 7 12 9 2
20 0 9 13 3 1 12 7 12 9 2 1 11 1 9 11 1 12 9 2 2
18 9 1 9 11 15 13 1 9 3 2 1 12 7 12 9 1 9 2
28 9 1 0 9 13 1 10 9 1 9 13 7 10 9 2 15 13 1 9 1 11 1 11 7 1 0 11 2
10 13 13 3 0 9 1 0 0 9 2
35 12 1 15 13 1 9 0 0 9 11 7 9 11 1 9 11 3 1 9 1 11 2 0 3 1 9 3 1 0 11 1 9 1 11 2
17 1 9 9 15 3 1 12 9 13 1 9 1 12 1 12 9 2
13 1 0 9 13 3 0 9 3 0 16 1 15 2
22 9 15 1 0 9 3 13 2 1 0 9 7 1 9 0 9 13 3 1 9 0 2
22 1 11 13 1 15 1 9 9 1 12 2 9 1 12 9 2 12 9 2 1 9 2
31 0 9 2 15 0 9 13 0 9 7 9 2 0 2 1 9 7 0 2 2 13 1 9 0 9 0 16 9 1 9 2
8 3 0 9 13 1 0 11 2
19 16 1 11 7 11 13 9 0 2 12 9 2 2 1 11 15 13 13 2
22 3 1 11 7 1 0 11 13 1 9 9 7 1 11 15 9 13 14 1 0 9 2
10 9 15 3 13 1 12 1 12 9 2
7 9 13 13 9 1 12 9
5 11 2 11 2 2
12 9 0 0 9 13 9 9 1 0 12 9 2
18 0 9 4 1 10 9 13 1 9 0 9 2 15 0 9 9 13 2
14 9 13 3 9 0 9 3 13 0 9 1 10 9 2
11 13 9 1 9 9 0 9 1 0 9 2
13 16 0 13 9 0 13 11 9 13 0 0 9 2
23 0 1 9 2 0 0 9 2 15 13 3 16 9 9 2 13 9 9 1 9 7 9 2
19 0 9 11 2 1 15 13 9 14 12 9 2 13 9 9 1 9 9 2
13 9 0 9 0 9 13 10 9 3 1 9 9 2
29 3 1 12 2 9 2 3 9 1 9 9 1 9 9 1 0 9 2 13 9 13 9 2 15 13 9 10 9 2
30 9 13 11 0 0 9 7 9 12 11 2 15 15 16 0 1 0 9 12 0 9 13 9 1 0 9 12 2 9 2
32 2 12 9 13 9 9 2 9 9 9 13 1 10 9 13 1 12 2 2 3 12 2 9 2 2 13 15 9 11 11 11 2
7 9 1 11 13 1 9 9
5 11 2 11 2 2
19 9 1 9 9 15 1 9 9 13 12 1 0 9 3 12 9 0 9 2
8 13 15 3 9 9 0 9 2
11 15 4 1 15 3 13 0 9 0 9 2
10 0 9 13 1 9 9 9 9 9 2
22 16 15 9 13 1 10 9 2 4 13 3 1 11 7 1 12 2 12 2 12 13 2
19 10 9 15 7 9 13 2 1 9 0 9 4 7 13 13 0 9 11 2
7 9 4 2 13 2 0 9
2 11 2
19 0 9 1 9 0 0 9 2 0 1 12 9 0 9 2 13 3 9 2
18 0 9 13 13 3 2 9 9 2 9 10 9 7 9 1 9 9 2
13 13 7 13 13 0 9 7 13 1 0 9 9 2
7 9 1 9 13 9 1 9
5 11 2 11 2 2
17 0 9 1 0 9 2 15 13 9 1 0 9 2 13 3 9 2
38 1 9 1 12 9 15 13 12 9 2 1 9 1 12 7 12 9 12 9 2 1 9 1 12 1 12 9 12 9 7 1 9 1 12 9 12 9 2
6 9 4 13 1 9 2
6 9 15 13 1 9 9
5 11 2 11 2 2
24 9 1 9 9 0 9 15 1 0 9 1 9 9 13 12 1 0 9 3 12 9 0 9 2
12 13 15 3 9 9 0 9 7 9 0 9 2
15 15 4 1 10 9 1 0 9 3 13 0 9 0 9 2
18 10 0 9 2 15 15 9 13 3 2 15 13 1 9 9 9 9 2
23 16 15 9 13 1 0 9 9 2 4 3 13 1 9 12 9 1 9 1 9 10 9 2
29 1 9 2 16 15 15 9 1 9 10 9 13 2 9 4 13 3 1 9 0 9 7 1 12 2 9 12 13 2
15 9 15 7 10 9 13 2 0 13 9 1 9 1 9 2
14 1 9 0 9 4 7 13 13 0 9 9 0 9 2
28 9 2 15 13 9 0 0 9 2 15 1 9 4 13 13 3 3 12 7 12 9 2 16 9 13 0 9 2
4 0 9 13 9
5 11 2 11 2 2
18 0 9 13 1 12 2 9 0 0 9 1 12 9 1 12 9 3 2
34 0 0 9 3 13 1 0 9 1 12 9 2 1 12 2 2 0 1 12 9 2 1 12 2 7 0 1 12 9 2 1 12 2 2
19 13 15 3 0 9 1 9 1 9 9 1 12 9 1 9 1 12 9 2
12 0 9 4 3 13 0 9 12 7 12 9 2
16 9 1 0 9 2 0 2 0 9 2 4 3 13 12 9 2
5 9 13 1 12 9
2 11 2
14 9 9 1 12 9 1 0 9 3 13 0 0 9 2
25 10 9 11 11 11 13 9 0 9 0 9 1 0 12 9 0 9 7 9 3 12 9 2 9 2
9 3 13 15 3 0 9 0 9 2
9 0 7 0 9 9 1 0 9 9
2 9 9
3 9 0 2
3 9 0 2
4 11 11 12 12
4 11 11 12 12
3 11 12 12
5 11 11 11 12 12
5 11 0 11 12 12
5 0 0 11 12 12
3 11 12 12
3 11 12 12
4 11 11 12 12
4 11 11 12 12
8 0 2 0 2 9 11 12 12
3 11 12 12
4 11 11 12 12
3 9 12 12
5 11 0 11 12 12
4 9 11 12 12
3 11 12 12
5 9 11 11 12 12
6 11 11 0 11 12 12
5 0 9 11 12 12
4 9 11 12 12
4 0 9 12 12
4 0 9 12 12
5 9 11 11 12 12
3 11 12 12
4 0 9 12 12
6 11 2 11 11 12 12
5 3 0 9 12 12
4 11 11 12 12
3 11 12 12
6 0 9 13 1 9 9
15 0 0 9 9 9 13 12 9 2 3 0 9 0 9 2
4 0 9 13 9
20 3 0 0 9 4 3 13 0 9 12 9 2 0 12 9 7 0 12 9 2
18 0 0 9 4 13 0 9 12 9 2 0 12 9 7 0 12 9 2
12 0 9 4 3 13 0 9 12 7 12 9 2
32 9 1 0 9 2 0 2 0 9 2 13 1 9 12 9 7 9 1 9 1 0 9 13 13 14 12 9 3 1 0 9 2
3 0 9 9
12 3 0 9 13 9 0 9 1 9 0 9 2
26 9 4 13 9 13 1 9 2 4 13 13 2 16 15 13 1 0 9 1 9 0 9 1 0 9 2
10 7 9 13 13 1 9 9 7 9 2
8 9 15 3 13 0 0 9 2
19 12 10 9 13 16 0 9 2 0 9 13 1 9 1 9 0 9 9 2
25 3 4 9 13 1 9 2 16 15 9 13 0 7 0 9 2 7 7 13 0 9 2 9 13 2
6 13 1 3 0 9 2
7 9 13 9 16 0 0 2
25 9 2 16 4 13 10 9 7 13 9 13 9 2 3 13 2 16 15 13 9 9 7 9 9 2
27 10 9 13 0 13 3 16 9 1 0 9 1 9 0 1 9 7 1 0 9 2 3 16 9 0 9 2
20 0 9 3 13 1 15 2 16 4 13 0 9 9 2 15 1 15 9 13 2
5 9 9 3 13 2
5 13 15 15 13 2
10 9 9 9 1 0 9 9 13 0 2
11 3 13 9 3 0 2 16 15 13 13 2
11 3 7 10 0 9 1 0 9 3 13 2
5 13 0 13 0 2
22 0 9 9 0 9 11 11 2 11 2 3 1 9 13 2 16 13 0 13 0 9 2
8 9 3 13 9 3 1 9 2
14 9 7 9 1 9 0 9 13 1 10 9 3 9 2
25 9 2 15 13 1 0 9 2 4 3 13 13 9 10 9 1 9 2 16 13 1 9 7 9 2
11 13 3 1 9 2 7 3 3 1 9 2
7 1 9 11 4 15 13 13
2 11 2
24 1 3 0 9 4 15 13 0 0 9 2 11 2 1 10 9 11 11 13 14 1 12 9 2
15 2 13 9 9 7 9 9 2 2 13 1 0 0 9 2
25 16 3 13 2 9 13 1 2 0 2 9 1 10 9 2 3 3 2 1 9 2 9 7 9 2
18 1 9 11 2 11 4 9 13 13 9 1 9 2 7 1 0 9 2
26 9 11 15 13 1 15 2 16 4 15 1 0 9 13 2 16 4 11 1 9 13 1 9 0 9 2
13 13 15 3 1 15 9 2 1 15 13 0 9 2
6 9 0 9 1 0 9
1 9
2 0 9
2 11 9
1 11
3 12 9 12
3 12 9 12
4 11 13 9 9
2 11 2
11 0 0 9 13 2 16 4 13 13 9 2
28 0 9 3 13 9 0 0 9 11 11 11 2 0 2 1 15 2 13 3 0 13 1 9 0 9 2 9 2
19 0 9 10 9 3 3 13 2 13 7 0 2 13 1 10 9 9 2 2
27 9 13 7 14 0 9 1 9 2 16 4 15 13 13 0 9 1 9 2 3 11 13 9 12 9 9 2
12 9 9 1 9 13 1 9 3 12 1 12 2
3 9 0 9
21 9 11 3 1 0 9 13 2 16 13 10 9 9 1 9 9 9 9 11 11 2
30 4 3 13 0 9 0 9 11 2 15 0 9 13 9 1 0 9 9 2 11 1 9 7 13 9 9 10 0 9 2
16 9 0 9 3 3 13 1 9 2 3 15 15 3 13 13 2
40 13 13 2 16 1 0 9 0 9 13 9 1 0 9 11 11 11 2 15 4 1 0 9 13 1 10 0 9 1 9 1 9 9 1 9 0 9 11 11 2
43 13 3 0 9 11 2 16 10 10 9 13 9 13 10 9 1 3 0 9 7 3 2 16 0 9 11 13 10 9 2 15 4 13 0 9 1 0 9 1 9 11 11 2
51 1 15 7 0 13 1 9 2 16 0 0 9 11 13 0 9 13 1 9 11 11 2 16 4 13 9 1 0 9 2 1 15 0 9 13 3 9 2 7 15 3 14 1 10 9 2 7 3 1 9 2
24 3 0 9 2 15 13 9 11 7 0 9 2 13 2 0 9 2 9 9 0 9 1 9 2
21 1 11 11 3 13 0 11 3 0 9 2 16 4 1 15 13 9 1 0 9 2
20 16 9 1 10 9 10 9 13 2 3 14 3 3 2 16 13 10 0 9 2
6 3 7 4 9 13 2
19 1 9 13 9 7 1 2 0 9 2 4 13 4 13 7 10 9 11 2
14 3 3 15 13 9 1 0 9 11 11 7 11 11 2
21 7 7 15 3 11 11 13 15 2 16 3 4 13 13 1 3 0 9 0 9 2
3 0 0 9
8 11 7 11 13 1 11 1 9
7 11 2 11 2 11 2 2
14 1 0 9 9 11 15 13 1 0 11 0 9 11 2
14 13 3 9 0 0 9 2 15 13 1 12 2 9 2
20 10 9 13 9 0 9 0 9 12 9 9 7 9 1 3 12 9 0 9 2
33 0 9 0 9 2 9 7 9 11 11 2 15 0 9 2 1 0 0 9 2 3 13 13 9 9 9 2 14 1 9 3 0 2
43 14 3 2 16 13 7 13 15 9 12 9 9 2 9 9 2 11 2 13 3 11 2 10 9 3 13 0 7 0 9 9 0 1 9 3 0 2 7 3 3 3 0 2
7 9 0 9 13 0 0 9
7 11 2 11 2 11 2 2
22 9 9 11 11 2 15 12 2 9 13 0 0 9 2 9 0 9 2 13 3 13 2
11 1 10 9 4 13 16 9 1 9 9 2
28 9 9 11 11 15 13 2 16 15 1 10 9 13 15 11 11 2 16 9 13 10 9 1 9 9 11 9 2
27 2 9 0 9 4 13 3 12 9 1 9 9 0 9 2 13 4 7 3 10 9 2 2 13 9 11 2
30 0 9 9 9 11 11 15 13 2 16 9 13 2 9 9 7 13 9 7 9 13 0 9 2 15 13 7 13 9 2
21 2 13 13 10 9 1 10 9 2 16 0 2 7 0 2 2 13 11 2 11 2
5 9 1 9 2 12
7 13 15 12 2 11 1 11
21 9 0 9 13 15 12 2 0 0 9 11 11 2 13 12 2 9 9 11 11 2
30 13 4 15 15 2 16 15 3 13 0 9 2 2 0 9 4 13 1 9 11 2 15 1 10 9 13 0 0 9 2
22 9 9 4 13 1 9 2 3 9 0 9 2 1 15 15 9 13 1 0 9 2 2
5 15 13 0 9 2
35 2 1 0 9 15 1 9 9 11 11 13 11 11 7 11 11 2 0 9 13 11 11 2 0 9 11 1 9 4 13 11 11 2 2 2
28 13 2 16 4 13 0 9 2 7 1 0 0 9 13 2 16 15 10 9 13 2 9 11 2 11 2 2 2
8 1 15 13 0 2 9 2 2
7 13 15 15 1 15 2 2
2 9 3
8 0 11 2 3 1 0 9 2
11 0 9 15 13 1 9 9 1 0 9 2
16 15 13 7 9 0 9 0 1 9 11 2 15 13 9 11 2
11 0 0 9 13 9 0 9 7 9 9 2
22 9 9 13 0 9 2 1 0 13 9 2 1 0 12 12 9 1 0 9 7 9 2
5 0 9 9 13 2
3 2 11 2
5 9 1 0 9 2
27 12 1 0 9 1 9 0 0 9 13 9 11 11 1 9 12 2 0 9 0 9 13 1 12 9 3 2
19 0 0 9 13 7 1 9 9 2 16 2 0 2 9 13 13 0 9 2
7 13 11 12 1 12 9 2
3 2 11 2
25 11 11 12 13 0 9 0 9 2 15 1 9 12 9 9 13 1 11 7 0 12 9 0 11 2
10 13 15 9 0 1 11 12 2 9 2
15 0 9 9 13 1 12 9 1 0 9 0 9 11 11 2
14 9 9 11 1 9 1 11 13 13 1 12 2 9 2
3 11 1 9
25 13 1 0 0 9 1 11 9 4 13 9 2 16 4 15 7 13 7 13 1 9 0 0 9 2
42 9 11 2 15 3 1 9 1 9 13 0 9 3 13 0 2 7 7 1 12 9 9 13 13 3 16 0 0 9 2 0 9 7 0 9 2 1 0 9 3 0 2
19 13 0 0 9 2 7 13 0 9 1 0 0 9 1 3 0 0 9 2
19 13 1 9 9 2 7 1 9 2 15 1 9 13 0 9 3 1 9 2
3 0 9 9
15 3 2 11 2 13 10 9 9 11 11 7 9 11 11 2
5 13 0 0 9 2
31 9 0 9 13 0 2 0 9 2 0 9 15 0 2 0 2 1 15 13 0 9 2 7 3 3 9 0 9 1 11 2
25 13 15 9 0 2 1 0 0 9 2 16 3 13 0 1 9 9 11 2 15 1 15 13 11 2
20 0 9 3 13 9 11 7 11 2 3 3 13 0 9 2 3 2 0 2 2
15 16 9 13 9 2 15 3 1 9 13 2 13 0 9 2
24 16 4 12 9 13 13 14 1 0 9 2 10 0 9 13 3 0 2 13 4 9 1 9 2
4 9 9 7 9
19 2 9 4 13 9 3 2 16 4 15 13 3 2 2 13 3 11 11 2
22 11 11 2 15 3 13 1 9 11 0 1 10 9 2 9 2 13 10 9 1 15 2
17 3 16 13 10 9 3 0 9 2 13 10 9 2 0 2 9 2
13 3 16 0 9 13 15 16 9 0 9 9 9 2
26 1 9 1 9 0 9 13 11 1 0 9 0 14 1 9 9 9 7 9 2 15 7 3 13 0 2
26 13 1 15 0 9 9 7 3 3 0 9 1 9 2 2 0 9 15 13 2 3 1 15 3 13 2
16 13 15 0 9 2 2 2 13 15 1 10 9 3 3 2 2
12 10 9 3 16 0 9 13 0 7 3 0 2
11 13 0 9 14 1 10 9 7 9 9 2
11 3 16 9 9 13 9 9 7 9 9 2
9 3 0 2 13 3 14 3 0 2
25 0 3 0 9 13 0 9 15 2 16 14 1 0 2 7 7 1 0 9 13 0 9 0 13 2
21 0 13 7 0 9 7 9 0 9 1 0 9 7 9 9 13 1 0 9 9 2
14 0 0 9 15 13 9 1 2 0 2 9 1 9 2
17 13 16 9 0 9 2 16 4 15 9 13 7 15 13 13 3 2
11 0 9 13 1 9 13 1 0 9 1 9
5 11 2 11 2 2
18 0 9 13 1 12 2 9 0 9 1 9 0 1 9 1 0 9 2
23 0 1 0 9 2 15 3 9 13 3 1 11 7 11 2 13 1 9 9 3 12 9 2
22 1 0 9 1 9 13 9 1 9 1 11 13 1 12 9 2 1 0 9 12 9 2
14 9 10 9 13 9 9 2 15 13 13 0 9 9 2
37 1 9 1 9 0 9 13 0 9 9 9 1 9 1 0 9 1 12 2 9 1 0 9 1 12 9 1 12 2 1 0 1 12 1 12 9 2
14 1 0 0 9 15 1 10 9 13 12 9 1 9 2
19 0 9 11 11 2 15 3 16 11 3 13 1 11 2 9 1 9 13 2
27 0 9 9 1 11 7 11 13 1 11 12 9 1 9 7 0 9 2 0 9 1 11 11 13 12 9 2
6 0 9 13 9 13 9
5 11 2 11 2 2
16 1 0 0 9 3 13 1 9 9 11 7 0 11 1 11 2
18 0 9 13 13 0 9 11 11 2 15 3 13 13 0 9 1 11 2
11 9 0 9 1 9 1 9 13 7 0 2
20 0 9 1 11 15 3 13 3 0 9 1 0 9 2 15 3 13 0 9 2
26 2 13 4 0 9 1 11 2 16 4 15 1 0 9 13 9 1 9 2 2 13 0 9 11 11 2
14 0 0 9 11 15 3 13 1 9 13 1 9 9 2
16 1 15 13 0 9 13 2 16 13 13 7 1 9 3 13 2
16 2 13 15 1 9 2 16 0 9 13 13 1 9 0 9 2
17 1 9 13 1 15 3 16 9 1 9 2 15 13 15 1 9 2
11 13 4 1 15 2 7 15 15 13 2 2
13 9 1 11 7 0 11 13 1 9 1 12 9 2
13 13 3 12 9 2 1 15 13 0 7 0 9 2
31 2 13 15 13 7 1 0 9 1 0 11 3 2 16 3 13 1 9 7 9 2 0 9 7 9 2 2 13 11 11 2
19 2 9 13 7 1 9 9 2 14 3 13 1 9 15 2 15 13 2 2
5 11 13 14 0 9
5 11 2 11 2 2
24 0 9 13 9 1 0 9 0 0 0 9 7 0 9 0 9 11 11 3 1 9 0 9 2
11 13 15 15 3 0 9 1 0 0 9 2
13 11 4 13 1 9 9 0 9 7 9 0 9 2
14 0 9 15 13 1 9 9 9 0 0 9 11 11 2
24 9 15 13 1 9 2 7 1 0 9 9 2 7 16 11 11 3 13 2 16 15 11 13 2
25 11 15 2 3 13 2 13 9 9 9 3 2 16 11 13 2 16 15 3 7 9 2 13 2 2
12 11 11 13 9 9 9 1 12 1 12 9 2
9 9 1 9 2 3 3 7 3 2
19 0 0 9 12 7 12 9 2 9 2 0 0 12 7 12 9 2 9 2
10 9 1 12 9 1 12 9 2 9 2
18 3 4 13 0 0 2 3 0 7 0 9 12 7 12 9 2 9 2
23 9 7 9 2 1 9 13 3 7 3 2 9 9 1 9 1 11 3 1 9 7 9 2
25 0 9 12 7 12 9 2 9 2 0 12 7 12 9 2 9 2 1 11 14 12 9 2 9 2
29 1 9 13 9 7 9 1 9 2 3 7 9 2 9 12 7 12 9 2 9 2 1 11 14 12 9 2 9 2
17 9 2 9 9 1 0 9 1 10 9 13 12 5 1 0 9 2
11 9 2 0 9 0 2 0 9 3 0 2
35 1 9 13 9 1 12 2 12 7 13 1 12 2 12 2 9 13 1 9 1 12 2 12 7 13 1 9 1 12 2 12 9 0 9 2
22 9 9 2 0 9 12 9 9 13 1 9 12 2 0 12 9 2 9 1 9 12 2
9 0 0 9 2 12 9 2 9 2
2 0 9
2 9 2
15 11 2 3 2 9 9 12 2 9 9 12 9 2 11 2
8 11 0 2 3 12 2 12 2
9 0 9 2 3 3 12 2 12 2
8 11 2 3 3 12 2 12 2
7 11 2 3 12 2 12 2
9 11 2 11 2 3 12 2 12 2
7 11 2 3 12 2 12 2
7 11 2 3 12 2 12 2
8 11 2 3 3 12 2 12 2
9 11 2 11 2 3 12 2 12 2
8 11 2 3 3 12 2 12 2
10 11 2 11 2 3 3 12 2 12 2
9 11 2 11 2 13 12 2 12 2
3 9 1 9
6 11 2 9 12 2 12
6 11 2 3 12 2 12
6 11 2 9 12 2 12
6 11 2 3 12 2 12
6 11 2 3 12 2 12
6 11 2 9 12 2 12
6 11 2 3 12 2 12
6 11 2 3 12 2 12
6 11 2 9 12 2 12
6 11 2 3 12 2 12
6 11 2 9 12 2 12
6 11 2 3 12 2 12
6 11 2 3 12 2 12
6 11 2 3 12 2 12
7 0 11 2 3 12 2 12
6 11 2 9 12 2 12
6 11 2 3 12 2 12
6 11 2 3 12 2 12
6 11 2 3 12 2 12
6 11 2 3 12 2 12
9 9 1 0 9 13 1 9 3 13
5 11 2 11 2 2
22 1 0 0 9 2 15 13 1 0 0 9 1 0 9 2 13 1 9 3 13 9 2
32 9 4 13 14 1 12 2 9 1 9 9 1 0 9 13 9 1 9 3 1 0 1 12 9 2 1 9 13 0 12 9 2
23 9 9 13 2 16 4 13 1 0 9 1 0 9 11 2 1 11 7 1 11 7 11 2
18 1 9 9 0 0 9 11 4 13 9 2 16 13 1 0 9 9 2
9 3 13 13 3 9 9 1 9 2
20 1 0 9 13 13 0 9 2 15 13 1 0 9 1 9 7 13 0 9 2
23 0 9 13 0 9 1 9 0 2 0 2 0 2 0 2 1 0 0 9 7 1 9 2
12 9 7 13 13 1 9 9 7 13 3 9 2
22 3 3 13 1 0 9 9 9 1 9 3 0 2 9 1 11 15 13 0 9 9 2
8 1 0 9 15 13 0 9 2
24 1 0 9 0 9 11 11 15 9 13 1 9 3 2 16 9 1 11 13 1 10 9 0 2
8 11 13 2 16 13 0 9 9
5 11 2 11 2 2
19 10 9 11 13 11 11 2 16 1 9 9 9 13 0 9 0 9 11 2
32 1 0 9 11 13 9 0 7 0 9 11 11 11 2 16 13 9 0 9 0 9 0 9 11 11 11 1 9 1 0 9 2
8 11 11 3 4 13 9 11 2
13 10 9 15 13 0 9 7 0 7 0 9 11 2
24 1 9 2 15 4 13 1 9 0 9 11 2 13 2 16 9 1 9 0 9 11 13 4 2
33 9 0 7 0 9 11 11 11 12 2 9 12 13 2 16 9 13 15 2 15 4 13 9 1 9 11 7 9 0 9 1 11 2
11 9 13 0 9 7 13 0 11 7 11 2
48 0 9 11 13 3 12 2 9 12 1 9 2 16 15 1 9 11 13 9 13 1 15 2 16 11 10 9 13 7 13 9 0 9 11 1 12 2 9 12 2 15 15 13 13 0 9 9 2
27 3 0 9 2 15 10 9 13 2 13 1 9 9 7 0 9 10 9 2 15 7 1 10 0 9 13 2
28 0 9 13 2 16 9 0 7 0 9 2 16 11 11 13 9 10 9 2 13 9 13 7 9 0 9 13 2
32 0 9 11 3 12 2 9 13 9 1 0 9 11 11 1 9 9 9 9 7 13 9 11 11 2 16 4 9 13 10 9 2
12 11 11 13 7 3 9 0 9 11 1 11 2
33 9 0 9 11 11 11 3 1 11 13 2 16 0 9 3 13 9 11 1 9 9 9 9 2 13 15 7 10 9 1 0 9 2
7 9 9 9 13 3 9 11
7 11 2 11 2 11 2 2
16 0 9 9 9 13 3 0 9 0 9 11 11 2 11 2 2
18 9 11 11 3 13 2 16 3 0 9 1 10 9 13 3 9 9 2
23 11 3 3 13 1 9 0 9 0 9 11 11 2 15 9 13 0 9 11 12 2 9 2
13 11 11 13 1 9 9 0 9 9 9 1 9 2
11 1 0 9 9 9 9 15 3 13 13 2
16 1 11 4 10 9 13 4 13 1 10 0 9 1 0 9 2
25 1 10 9 2 3 13 9 1 9 9 9 9 2 11 11 13 2 2 1 9 13 0 3 13 2
26 10 9 13 13 1 0 9 9 2 7 16 13 10 9 13 2 13 0 2 16 4 1 9 13 2 2
17 1 9 2 16 13 1 11 11 1 10 0 9 2 13 9 3 2
16 9 15 3 1 9 11 1 9 1 9 13 1 9 9 9 2
21 15 3 1 9 13 0 9 7 13 3 1 9 7 1 15 2 16 4 15 13 2
22 10 9 13 1 15 0 2 16 3 13 10 2 0 9 2 13 9 1 2 9 2 2
11 1 0 9 9 13 0 9 14 12 9 2
19 1 15 15 7 13 7 1 9 9 9 1 9 9 2 15 13 0 9 2
3 2 11 2
6 9 2 11 2 11 11
8 0 9 0 9 13 9 9 9
5 11 2 11 2 2
31 0 9 9 0 0 9 11 11 13 9 1 9 9 1 0 0 9 16 9 0 0 0 9 7 1 9 9 9 11 11 2
29 11 3 16 9 0 9 13 1 9 0 9 9 2 1 15 13 1 9 0 0 9 2 15 13 0 9 11 11 2
28 11 11 15 13 1 0 9 16 9 0 0 9 1 0 9 9 1 9 0 9 13 0 9 9 9 0 9 2
22 3 1 15 13 0 9 1 9 1 10 0 9 7 9 0 0 0 9 11 2 11 2
36 11 1 10 9 3 2 13 9 0 9 2 1 15 11 2 11 2 1 9 1 15 0 9 11 11 13 1 9 12 0 9 1 0 9 11 2
11 10 9 7 4 1 9 1 0 9 13 2
29 15 1 0 9 12 13 0 9 1 0 9 2 16 1 0 9 4 3 1 9 1 9 12 13 3 16 12 9 2
21 9 13 1 9 13 11 2 11 2 7 11 15 13 2 16 4 1 15 13 9 2
12 0 0 9 1 0 11 0 9 11 11 13 2
10 3 4 10 9 13 0 9 1 11 2
4 0 9 13 9
5 11 2 11 2 2
13 9 7 9 0 0 9 3 13 1 9 11 11 2
28 1 9 9 13 1 9 9 11 11 2 11 2 7 10 9 15 13 11 11 2 11 2 2 12 0 9 11 2
17 1 9 13 2 16 16 15 13 0 2 13 10 9 1 0 9 2
11 16 7 13 2 9 13 13 9 1 9 2
8 0 9 9 11 13 12 9 2
12 9 13 3 10 9 1 0 9 2 3 9 2
11 11 13 9 1 0 9 7 9 9 9 2
5 11 11 7 10 9
12 9 2 9 2 9 2 9 2 7 11 3 13
2 11 2
26 0 9 1 9 11 11 15 1 0 9 13 1 10 9 11 11 1 0 9 1 9 1 11 2 11 2
17 3 13 1 0 9 1 11 11 1 0 9 1 9 9 1 11 2
11 4 15 3 13 10 9 10 0 0 9 2
24 3 9 11 2 9 11 2 9 11 2 9 1 9 2 7 3 0 9 11 2 3 0 9 2
12 0 0 9 0 1 0 9 1 11 13 9 2
6 15 3 1 15 13 2
30 9 0 11 2 15 0 9 7 13 11 11 2 1 15 13 2 2 0 9 13 11 2 9 7 0 9 15 13 11 2
24 3 13 3 12 0 9 2 15 15 1 9 13 2 9 11 2 9 1 9 11 7 9 11 2
10 13 4 2 3 0 13 13 0 9 2
11 15 10 15 3 13 15 0 9 1 0 2
9 1 9 4 13 1 9 14 9 2
17 14 7 10 0 9 13 11 11 7 9 1 9 1 9 11 11 2
13 15 13 1 11 2 7 3 13 12 9 1 11 2
7 13 10 9 10 9 13 2
16 10 9 13 0 9 2 15 15 3 13 3 14 1 0 9 2
11 1 10 9 3 4 13 9 13 3 2 2
27 1 9 2 16 9 11 2 3 15 11 13 2 13 3 9 9 2 9 13 2 2 15 3 13 1 9 2
8 1 12 9 4 13 14 9 2
5 15 3 3 13 2
8 9 1 15 13 14 9 9 2
9 9 1 0 9 13 3 0 2 2
18 11 15 13 2 16 1 15 9 10 9 15 13 0 9 13 7 3 2
19 2 13 2 16 4 9 13 3 2 7 15 15 15 4 13 1 0 9 2
14 13 10 9 9 1 0 9 4 7 13 3 0 2 2
19 1 9 12 15 11 11 13 2 16 1 9 10 9 13 3 12 9 9 2
23 2 16 4 7 13 15 13 7 2 16 13 2 13 4 13 3 12 9 2 2 13 11 2
13 2 7 15 13 7 9 1 15 2 15 13 2 2
34 0 0 9 11 11 1 15 13 2 2 13 4 0 2 16 4 15 3 13 13 14 7 14 1 0 9 2 16 0 4 13 0 9 2
6 7 3 13 9 2 2
29 11 11 15 3 1 9 10 9 13 1 9 9 2 12 2 1 10 0 9 1 9 9 7 0 9 11 2 11 2
23 0 9 1 9 9 11 2 7 3 7 1 9 9 1 11 2 7 13 1 0 9 0 2
10 1 9 15 13 13 7 10 0 9 2
33 2 3 13 2 2 13 1 15 11 2 2 3 15 13 3 14 13 2 16 4 1 11 13 3 3 2 16 3 13 11 2 11 2
3 14 13 2
5 13 15 16 9 2
9 16 13 13 0 2 3 13 0 2
15 7 16 15 13 15 1 0 9 2 13 13 9 9 2 2
24 9 11 11 1 10 0 9 2 9 1 12 5 12 9 2 1 15 1 9 11 13 1 0 9
4 3 1 9 9
2 11 2
17 1 9 13 3 12 0 9 2 10 9 15 4 13 9 0 9 2
22 1 11 13 11 11 1 11 11 2 1 3 0 0 9 15 13 11 11 7 11 11 2
18 9 9 11 2 16 0 2 13 1 0 9 0 0 9 2 11 2 2
17 1 15 15 13 7 0 9 11 11 7 11 1 0 9 12 13 2
20 9 13 1 9 3 13 1 0 12 1 9 9 2 9 9 11 7 11 11 2
12 12 9 4 13 3 0 9 12 9 0 9 2
15 1 0 9 15 7 2 16 0 2 13 3 11 11 11 2
3 11 13 9
5 11 2 11 2 2
23 14 1 0 0 11 2 7 3 1 9 9 3 13 11 11 1 9 0 9 11 0 11 2
24 2 9 13 1 9 0 2 15 3 1 0 9 3 13 2 2 13 0 0 9 1 10 9 2
19 0 0 9 13 0 0 9 9 0 9 1 9 1 9 12 9 0 9 2
24 0 0 13 0 9 11 11 1 11 11 7 3 11 11 2 9 0 9 1 9 12 2 12 2
24 16 15 12 3 13 2 1 0 9 13 13 9 9 2 15 13 1 11 2 13 0 9 2 2
88 9 2 9 2 9 2 11 2 11 12 2 12 2 12 2 12 2 11 2 11 2 11 12 2 12 2 12 2 12 2 11 2 11 12 2 12 2 12 2 12 2 11 2 11 2 12 2 12 2 12 2 12 2 12 2 9 2 9 2 11 2 11 12 2 12 2 12 2 12 2 12 2 12 2 11 2 11 2 12 2 12 2 12 2 12 2 12 2
5 9 1 0 2 11
6 0 11 2 11 2 2
10 1 12 0 9 4 13 9 0 11 2
28 0 9 0 9 13 9 0 11 1 12 9 2 3 1 12 0 9 13 7 9 2 15 3 13 1 10 9 2
26 9 13 3 9 11 1 9 11 2 0 9 13 7 11 2 11 2 7 3 15 0 11 2 11 2 2
17 1 9 13 3 12 9 1 9 1 0 9 7 9 1 12 9 2
5 9 1 12 9 2
11 10 9 2 11 2 11 2 11 2 11 2
6 11 2 11 2 11 2
3 9 2 9
20 9 12 1 12 2 12 2 12 2 12 2 12 2 12 2 0 9 2 12 2
6 15 15 1 11 3 13
3 0 11 2
20 0 9 11 11 0 9 1 0 12 9 13 1 10 9 1 0 9 9 11 2
13 1 0 9 15 1 0 9 13 0 11 11 11 2
13 0 9 2 0 12 9 2 13 10 9 0 9 2
22 7 12 0 9 15 7 15 13 2 9 13 14 0 9 2 16 0 9 15 3 13 2
19 1 12 2 9 13 9 11 2 1 11 2 11 2 11 2 11 7 11 2
16 10 9 15 3 1 15 13 9 1 0 0 9 7 12 0 2
15 3 15 1 9 13 11 2 11 7 11 7 16 0 11 2
18 1 9 1 11 13 3 0 11 2 7 7 15 15 3 13 1 9 2
18 0 9 15 13 11 2 15 13 1 12 2 9 7 3 13 0 9 2
13 9 13 14 1 0 12 9 7 15 3 13 3 2
13 9 2 12 2 9 2 0 2 12 9 2 12 2
3 11 9 9
5 0 9 15 13 13
7 11 2 1 10 9 2 2
17 1 0 9 1 0 9 15 13 0 11 11 9 9 1 0 9 2
13 0 9 10 9 13 2 16 13 1 9 0 9 2
21 9 10 9 13 9 0 9 7 15 0 0 9 11 2 3 9 10 2 13 15 2
3 9 9 11
7 11 1 11 11 3 0 9
5 11 2 11 2 2
40 3 9 15 9 11 11 13 1 0 9 2 1 9 7 1 9 1 2 0 2 9 15 13 9 11 11 2 11 2 15 4 11 2 13 2 1 0 2 11 2
27 2 3 13 1 3 0 9 1 0 11 2 16 1 0 0 0 9 13 14 1 0 9 2 2 13 11 2
40 2 10 0 9 13 2 7 3 7 4 13 9 0 9 7 13 2 16 9 11 2 11 2 9 2 15 4 13 1 9 7 13 1 11 13 2 1 15 13 2
28 1 10 9 1 0 0 9 3 1 11 4 15 1 10 9 13 2 13 3 9 13 2 15 1 15 13 2 2
41 1 9 13 0 1 0 9 1 0 11 2 1 10 9 3 12 2 9 13 0 0 9 1 11 11 2 1 9 1 15 13 3 1 12 2 9 2 1 0 11 2
5 0 9 1 9 11
2 11 2
35 9 0 0 9 11 11 2 15 13 1 9 12 1 9 1 9 9 1 9 0 9 9 11 11 2 13 12 9 9 1 9 1 10 9 2
15 9 4 13 9 11 11 2 15 0 9 9 13 1 9 2
16 9 9 4 13 1 0 9 1 11 2 1 15 11 11 13 2
4 9 13 0 9
2 11 2
29 0 9 11 2 15 15 13 0 9 11 2 11 2 13 10 0 9 2 10 9 13 1 0 9 9 0 0 9 2
16 9 13 7 9 2 16 4 13 0 9 2 16 4 9 13 2
26 9 7 9 9 11 11 2 15 9 11 1 9 13 2 13 2 16 13 1 9 13 9 7 15 3 2
3 0 0 9
8 0 0 9 9 0 1 9 9
8 11 2 1 10 0 9 2 2
40 3 2 3 1 0 9 9 2 12 13 9 9 9 1 0 9 3 9 9 11 1 0 9 2 13 11 11 10 9 2 13 0 9 2 7 9 3 13 13 2
8 4 1 15 13 12 0 9 2
19 13 15 15 1 0 9 0 9 0 9 7 13 15 0 9 1 0 9 2
16 2 11 13 9 1 9 7 13 9 2 2 13 9 11 11 2
6 2 13 15 15 2 2
10 2 13 15 9 2 15 13 3 3 2
9 13 15 9 2 2 13 0 9 2
19 0 9 13 1 0 9 3 12 0 9 2 13 3 3 12 9 1 9 2
21 1 0 9 4 13 12 9 1 12 9 2 11 13 12 2 11 7 11 1 12 2
11 11 13 3 16 0 7 13 1 15 11 2
25 2 16 4 13 2 16 13 11 9 3 1 0 9 2 13 4 2 16 15 3 13 2 2 13 2
7 0 9 15 13 0 9 2
11 2 13 4 1 9 2 2 13 9 11 2
16 2 13 15 2 16 16 1 9 13 0 9 2 13 15 0 2
11 0 4 13 2 16 4 13 12 0 9 2
14 11 13 1 9 0 7 10 9 3 14 13 3 2 2
9 11 11 13 9 3 7 1 9 2
20 1 12 9 15 13 9 9 2 1 15 10 0 9 13 13 9 9 9 9 2
34 2 16 4 15 15 3 13 3 12 0 9 2 15 3 13 3 15 2 2 13 11 2 9 2 15 13 1 10 9 7 9 3 0 2
10 0 9 9 13 1 9 1 0 9 2
24 1 9 1 9 15 1 9 9 13 1 0 12 15 12 0 9 2 11 2 11 1 0 9 2
18 1 9 9 13 1 12 9 11 1 12 2 7 11 1 12 2 9 2
2 11 2
2 11 2
18 0 9 11 11 13 1 0 9 1 11 0 0 9 1 12 9 9 2
2 1 9
29 1 0 0 9 1 11 13 0 9 0 9 1 9 12 5 12 9 2 12 2 12 2 0 9 1 12 0 9 2
11 12 9 13 1 0 9 1 11 0 9 2
22 11 13 12 9 0 9 9 12 2 12 2 11 13 0 1 0 9 1 12 2 12 2
20 0 9 0 9 11 7 11 13 11 11 1 11 1 11 2 15 13 0 9 2
21 0 9 11 0 11 11 2 15 9 13 3 0 11 11 2 13 9 1 0 9 2
15 11 13 13 0 9 1 9 0 9 1 9 7 1 9 2
21 0 9 0 0 9 1 9 12 4 13 0 9 12 9 7 0 9 1 0 9 2
15 9 11 13 0 9 9 12 1 11 7 9 12 1 11 2
10 0 9 0 9 13 9 12 9 9 2
1 9
9 11 11 2 0 11 12 2 12 2
9 0 9 1 0 9 1 0 11 2
14 1 9 13 9 1 0 11 7 0 9 13 1 9 2
9 0 9 13 0 9 11 7 11 2
20 1 0 9 15 13 9 12 0 9 2 9 9 2 9 2 11 7 9 11 2
7 11 9 9 1 12 9 2
12 11 2 11 12 2 12 2 12 2 12 2 2
13 11 13 1 9 2 3 15 13 1 11 1 11 2
4 11 13 1 9
11 11 2 9 2 11 2 11 2 11 2 2
5 0 9 13 9 2
5 11 13 15 7 13
2 11 2
30 11 11 11 13 9 1 9 0 9 7 13 0 9 0 9 11 1 11 2 15 13 1 11 1 11 7 13 12 9 2
3 11 1 9
2 11 2
15 9 0 0 0 0 9 11 11 1 9 1 11 13 13 2
31 0 0 9 1 9 1 11 13 1 9 9 2 9 0 9 2 1 9 1 9 9 0 9 0 9 7 13 15 13 9 2
9 0 9 4 13 13 1 0 9 2
5 0 9 12 3 0
6 13 12 2 9 9 11
6 0 11 2 11 2 2
27 0 12 2 9 9 11 2 9 0 1 9 12 1 0 9 9 11 2 13 3 1 12 9 1 0 11 2
16 0 9 13 3 14 3 1 9 2 9 15 13 1 9 9 2
17 0 9 12 2 3 0 1 9 0 11 9 11 2 7 13 13 2
10 11 3 13 13 0 9 1 11 9 2
18 0 2 9 2 3 13 0 9 9 11 11 2 2 9 2 0 11 2
16 1 9 13 7 0 0 9 2 11 2 11 2 11 2 3 2
10 9 9 13 0 0 9 0 9 9 2
29 1 11 13 0 9 11 11 10 9 2 12 11 2 12 11 2 12 11 2 1 9 13 7 9 1 11 7 11 2
27 9 9 11 13 3 7 9 11 11 1 11 9 12 2 11 11 1 11 7 11 1 11 1 11 11 11 2
11 0 13 7 0 9 1 9 1 9 11 2
7 11 13 3 0 9 9 2
24 9 11 13 0 12 9 7 13 12 0 9 2 12 9 2 2 1 9 12 2 1 9 12 2
15 1 9 1 0 11 13 0 9 1 9 1 12 2 9 2
3 13 4 15
2 16 11
24 0 9 11 11 10 0 9 1 12 2 9 0 9 1 11 13 3 9 11 1 9 11 12 2
12 3 4 11 1 9 13 7 16 9 13 11 2
7 7 15 15 13 9 11 2
20 9 11 11 15 3 3 13 1 9 16 9 2 14 3 2 3 11 11 13 2
37 9 9 11 11 13 0 9 7 1 0 9 9 11 1 9 1 11 2 3 0 9 13 15 2 15 15 13 1 9 2 15 4 1 11 3 13 2
3 2 11 2
2 0 9
18 9 11 15 13 1 9 10 0 9 1 11 2 11 11 2 1 11 2
18 13 7 1 10 9 2 15 13 1 9 3 1 9 1 3 0 9 2
3 14 3 2
22 13 1 0 9 13 1 9 3 3 2 13 2 7 1 9 9 15 13 14 1 9 2
20 12 0 9 1 15 13 0 9 2 3 16 15 13 2 1 9 2 9 11 2
11 9 15 13 2 9 9 1 0 9 13 2
10 0 9 3 13 0 9 1 15 3 2
3 2 11 2
6 1 11 13 9 12 9
5 0 9 13 1 9
2 11 2
25 0 11 13 1 9 2 10 9 4 13 1 12 9 9 2 7 13 15 9 9 7 3 7 9 2
28 9 15 13 1 9 2 16 1 9 13 1 11 11 11 1 12 9 9 2 16 13 1 9 3 1 9 9 2
24 2 9 1 11 13 12 9 2 2 13 0 9 11 2 16 13 1 3 0 9 1 12 9 2
10 3 1 11 13 13 13 1 0 11 2
13 0 9 15 13 1 9 13 9 11 1 11 11 2
20 0 9 1 9 12 9 9 3 13 2 1 0 7 13 9 1 9 1 11 2
19 1 9 11 11 1 0 0 13 2 7 11 13 0 13 10 0 0 9 2
22 9 11 13 3 1 9 1 9 3 16 12 12 9 2 15 13 7 14 9 1 9 2
17 9 9 11 11 2 0 9 7 9 9 2 7 3 3 13 9 2
19 2 1 0 0 9 11 13 1 12 9 7 4 13 1 9 2 2 13 2
5 10 9 13 1 11
5 11 2 11 2 2
27 1 9 1 0 9 2 15 15 13 1 9 12 2 2 12 2 9 1 11 2 15 4 13 1 0 9 2
26 10 9 13 9 11 11 11 11 11 2 15 15 13 2 2 11 13 7 0 0 9 2 7 9 0 2
5 0 9 15 13 2
9 7 4 1 15 13 9 15 2 2
19 1 11 13 3 12 9 1 0 11 2 11 2 11 1 11 7 1 11 2
24 11 13 9 2 12 9 1 9 2 2 0 9 7 0 9 2 3 12 9 1 9 12 9 2
20 0 9 13 1 9 3 7 3 2 9 15 3 3 13 3 1 9 9 9 2
5 0 9 3 3 0
6 9 11 1 9 13 9
2 11 2
26 11 11 2 0 9 2 15 13 9 2 16 15 1 9 0 9 9 1 9 9 1 0 9 13 9 2
16 13 1 12 9 3 2 16 13 0 0 9 9 2 12 9 2
5 15 13 13 9 2
16 1 0 0 9 13 9 3 1 12 7 3 1 12 9 3 2
10 0 9 3 13 9 0 9 11 11 2
21 2 9 2 2 13 2 2 10 9 13 13 3 0 9 2 16 4 13 3 13 2
8 7 16 3 13 2 2 2 2
4 11 15 13 2
22 2 16 13 9 0 2 13 12 9 2 7 16 13 0 2 12 9 2 2 13 11 2
15 2 15 4 13 2 16 15 1 15 1 9 3 13 2 2
4 15 15 13 2
16 11 13 1 0 9 13 9 0 9 2 7 15 13 1 9 2
12 13 1 9 0 9 1 9 12 7 12 9 2
13 2 13 15 1 0 9 1 9 9 2 2 13 2
16 0 9 1 0 9 2 1 0 9 9 1 9 2 13 3 2
22 2 0 9 15 3 13 3 2 16 13 3 0 2 7 15 3 13 1 9 1 9 2
14 10 0 9 13 2 7 16 4 15 13 14 12 9 2
13 7 7 13 1 0 2 2 13 0 9 11 11 2
13 2 15 15 3 13 0 13 0 9 1 12 9 2
13 7 16 15 1 12 9 13 2 0 15 13 2 2
12 0 9 13 13 9 2 13 0 9 7 9 2
6 7 13 10 9 9 2
12 1 9 11 15 11 13 2 7 7 9 13 2
16 2 13 15 9 2 9 2 7 15 4 13 2 2 13 11 2
9 1 0 9 13 3 13 10 9 2
6 13 13 13 3 9 2
18 10 0 9 15 3 13 2 10 0 0 9 13 13 1 9 1 9 2
10 0 9 1 10 9 9 13 0 9 2
4 13 9 11 2
18 2 15 13 10 7 0 9 2 13 15 1 0 9 2 2 13 11 2
13 13 3 0 9 2 15 1 10 9 13 10 9 2
24 11 11 13 1 9 1 9 9 11 11 7 9 11 13 0 9 1 10 0 9 1 0 9 2
10 13 15 1 11 9 9 0 9 11 2
13 2 15 15 13 13 2 7 3 15 12 9 13 2
6 13 9 2 7 13 2
15 13 1 9 2 7 1 15 13 13 2 2 13 9 11 2
24 1 0 9 13 9 0 9 2 1 15 13 13 3 1 10 9 2 1 9 2 9 2 9 2
23 0 9 13 3 1 12 12 9 2 1 0 9 2 0 11 7 0 11 2 13 3 0 2
14 9 11 16 0 9 13 1 10 0 9 11 7 11 2
12 2 0 9 1 11 13 2 2 13 11 11 2
12 2 9 4 15 13 2 7 0 9 13 2 2
18 2 15 15 15 13 2 2 13 11 11 2 2 7 15 15 13 13 2
13 1 9 13 16 9 12 0 7 12 0 9 2 2
36 12 1 0 9 1 9 9 13 0 0 9 2 1 15 11 11 11 2 0 11 2 15 15 1 11 13 2 7 11 11 13 0 9 1 9 2
14 11 12 2 0 1 0 9 2 13 1 12 0 9 2
4 11 13 1 9
6 0 9 9 0 0 9
2 11 2
20 9 9 7 3 0 9 9 2 15 13 0 9 2 15 13 1 9 0 9 2
25 13 15 2 16 15 0 9 13 12 9 7 12 9 1 12 9 2 0 9 7 13 14 12 9 2
7 9 13 0 13 1 9 2
23 9 9 11 13 9 1 9 12 9 0 9 1 9 1 9 2 15 1 10 0 9 13 2
11 0 9 1 0 9 13 11 12 2 12 2
4 1 0 9 2
23 11 2 11 12 2 12 2 11 2 11 12 2 12 2 0 9 2 2 11 12 2 12 2
7 9 0 9 13 0 9 2
14 9 0 9 13 9 1 9 2 3 1 15 13 9 2
22 1 12 9 9 13 9 9 9 13 1 9 11 2 7 9 9 11 1 10 9 13 2
7 9 3 13 1 0 9 2
19 9 9 11 11 2 11 2 7 9 9 11 11 2 11 2 1 0 9 9
8 9 13 0 9 0 9 11 11
5 11 2 11 2 2
39 0 0 9 9 2 12 9 0 1 0 9 11 11 4 13 3 1 9 0 9 13 0 9 11 2 12 2 11 2 12 2 11 2 12 7 9 2 12 2
11 13 15 3 9 9 7 0 9 11 11 2
18 1 15 4 9 1 9 12 13 12 7 12 0 9 9 2 12 9 2
11 11 11 3 9 13 3 0 9 0 9 2
17 9 3 13 1 9 0 9 2 16 0 0 9 1 0 9 13 2
17 9 9 2 12 9 4 9 13 1 0 9 9 1 11 2 11 2
21 3 4 15 13 13 13 7 1 0 9 9 2 12 9 2 15 4 13 0 9 2
10 9 0 9 13 13 9 1 11 11 2
16 11 13 7 9 9 9 2 12 9 1 9 0 9 0 0 2
12 10 9 13 0 9 9 7 14 3 0 9 2
27 3 13 13 2 16 9 4 1 9 13 12 9 2 9 7 9 2 7 14 9 1 10 9 9 2 12 2
7 9 12 0 1 9 3 0
5 11 2 11 2 2
27 1 0 0 9 2 1 15 12 9 13 7 12 4 3 13 2 13 1 9 1 9 1 9 11 1 11 2
17 1 9 11 1 0 0 9 7 11 12 15 12 9 13 7 13 2
13 9 11 15 13 13 7 1 0 9 13 1 9 2
17 9 0 9 9 2 15 13 1 0 9 2 15 1 9 13 13 2
4 0 9 13 9
7 11 1 11 2 11 2 2
27 9 0 0 9 1 11 1 11 13 1 9 0 9 11 0 11 1 11 2 15 13 9 1 9 0 9 2
29 9 13 0 7 0 9 2 9 7 9 7 13 0 9 1 12 0 9 2 16 9 13 13 9 9 0 0 9 2
22 11 13 0 9 0 9 13 9 1 11 2 1 15 13 0 9 1 0 9 3 0 2
21 11 2 3 0 0 9 2 13 9 13 0 0 9 1 0 11 1 0 0 9 2
8 9 1 12 9 14 13 1 9
6 0 11 2 11 2 2
24 12 9 0 9 2 9 1 3 12 9 9 15 3 1 9 13 1 9 11 1 11 1 11 2
8 9 3 13 1 9 0 9 2
23 1 9 3 3 0 11 11 2 1 11 1 2 11 2 13 2 16 0 9 13 1 9 2
18 1 9 11 13 12 0 11 11 2 1 9 12 10 3 3 0 9 2
13 11 11 2 7 11 11 2 7 9 3 13 13 2
8 9 13 3 1 9 1 11 2
10 1 9 1 9 3 13 13 12 9 2
17 10 9 11 11 2 13 1 9 3 1 11 9 12 7 12 9 2
19 1 0 11 15 1 9 1 11 13 0 12 9 1 9 7 12 1 9 2
9 3 3 13 9 1 12 12 9 2
5 13 9 2 13 11
6 0 11 2 11 2 2
15 9 1 11 15 13 0 11 1 9 1 9 1 0 11 2
27 13 13 3 3 2 7 16 15 3 1 12 9 13 1 9 2 3 13 9 1 12 9 9 2 13 15 2
5 9 1 9 13 9
5 11 2 11 2 2
14 9 2 15 13 0 0 9 1 11 2 13 9 9 2
21 9 13 13 2 1 10 9 15 4 13 1 9 2 0 9 0 9 0 0 9 2
15 9 9 0 0 9 0 13 1 0 9 1 11 9 9 2
9 0 9 4 1 9 13 1 9 2
5 0 9 13 1 11
5 11 2 11 2 2
32 0 9 0 11 13 1 9 11 1 11 3 3 12 9 1 0 11 2 3 0 9 7 13 2 7 13 3 0 16 1 11 2
12 0 9 11 1 11 15 13 1 12 12 9 2
28 9 9 1 11 13 0 9 9 2 16 1 15 4 9 1 11 0 9 9 1 0 9 7 0 0 9 13 2
13 0 9 0 11 13 3 1 9 3 12 9 9 2
13 0 9 13 1 11 1 9 7 13 3 1 9 2
12 1 9 13 3 3 1 9 1 9 9 3 2
23 9 1 0 9 13 0 9 11 2 15 1 0 12 9 13 1 9 11 3 12 9 9 2
10 10 9 13 1 0 0 9 0 9 2
17 1 11 11 2 9 1 9 11 1 11 2 0 9 10 9 13 2
4 0 9 13 9
6 0 11 2 11 2 2
24 1 9 9 2 9 0 9 2 9 0 9 13 3 0 9 1 0 11 0 9 11 0 11 2
26 9 13 3 0 9 1 0 9 1 11 9 1 9 2 15 13 9 0 9 2 7 1 9 11 13 2
15 0 9 1 10 9 13 3 9 2 9 2 9 7 9 2
26 1 0 9 0 9 3 13 3 9 11 11 2 9 11 2 0 9 2 9 11 1 11 7 11 11 2
5 9 9 1 11 13
6 0 11 2 11 2 2
45 0 9 0 9 1 0 9 2 15 3 3 13 9 1 11 2 4 13 1 0 0 0 9 1 11 2 3 15 1 12 2 9 1 12 2 9 13 1 12 9 0 7 0 9 2
14 1 9 9 11 11 0 9 13 1 9 1 9 9 2
5 3 3 1 9 9
12 9 9 1 9 0 9 9 9 13 10 9 2
20 13 15 7 13 10 0 9 7 15 13 1 0 2 0 9 1 0 10 9 2
18 9 10 9 14 13 10 0 9 15 2 16 1 9 13 10 0 9 2
6 13 3 9 0 9 2
17 12 2 9 2 7 13 1 0 9 2 13 1 9 12 3 3 2
31 3 3 3 1 9 9 1 0 9 2 14 1 15 2 16 4 15 13 0 9 2 14 1 15 2 16 13 14 9 10 2
21 9 13 3 1 15 2 15 9 16 9 7 15 0 9 2 3 2 2 3 13 2
16 13 2 14 3 2 16 15 13 2 13 13 15 0 16 9 2
21 15 13 9 1 10 9 7 16 13 2 15 1 9 0 9 15 3 7 13 13 2
42 12 2 1 0 2 0 2 3 0 9 2 0 1 3 0 7 0 0 9 7 1 0 2 3 0 2 9 2 13 10 0 9 9 7 13 9 0 9 9 10 9 2
19 7 15 4 15 13 2 3 10 0 0 9 2 15 10 9 7 9 13 2
23 9 13 1 15 2 16 1 10 9 13 0 9 1 15 2 16 4 9 13 13 0 9 2
18 13 2 14 10 9 2 13 15 1 0 0 2 3 0 9 10 9 2
33 9 15 13 3 2 9 9 13 2 9 13 9 0 9 10 9 2 9 15 13 3 2 9 13 3 9 1 9 2 3 2 3 2
40 3 13 0 9 2 13 2 16 15 15 10 9 13 2 13 15 1 9 0 9 2 13 1 0 9 15 0 9 2 7 1 10 0 9 0 0 9 3 13 2
23 9 3 13 2 7 16 15 9 2 3 1 0 9 10 9 2 13 2 13 10 0 9 2
32 9 15 13 3 3 2 16 15 13 13 3 0 9 1 0 7 0 9 2 9 2 15 13 9 1 9 9 7 1 9 9 2
5 7 15 13 13 2
19 3 9 9 1 0 0 9 7 1 9 15 2 16 13 3 0 7 0 2
35 0 9 4 13 2 16 4 13 2 16 3 2 13 2 0 2 15 13 9 1 9 12 1 9 12 1 3 16 0 2 1 15 0 9 2
17 15 4 13 9 7 13 4 15 9 3 1 0 0 9 0 9 2
4 3 15 13 2
24 16 9 1 9 12 13 1 10 0 9 3 16 3 2 13 9 13 1 0 9 16 9 1 9
11 13 9 11 7 0 0 9 2 3 14 2
17 9 2 15 13 9 3 1 12 5 2 13 13 9 1 12 5 2
5 13 15 9 15 2
33 1 15 13 15 0 9 15 9 2 16 4 15 2 15 13 9 1 12 5 7 9 1 12 5 2 13 9 2 16 15 13 3 2
25 9 9 11 1 11 2 16 15 3 9 15 3 13 7 16 15 13 0 13 1 9 2 13 0 2
22 3 15 13 2 3 15 15 3 13 2 3 13 9 13 15 1 9 0 9 1 9 2
7 7 7 15 3 13 15 2
11 13 2 16 13 9 10 0 9 13 9 2
16 16 13 3 2 0 0 9 2 15 13 9 14 1 0 9 2
10 7 9 3 13 9 7 13 0 9 2
41 16 4 15 4 13 2 13 0 10 9 3 12 0 9 2 15 13 2 16 3 0 9 13 13 9 0 9 14 3 2 16 9 0 7 0 9 9 13 12 5 2
14 7 10 0 9 13 10 9 2 9 2 7 9 9 2
9 1 9 7 1 0 9 13 2 16
9 13 2 16 15 9 10 15 13 2
33 14 2 14 2 13 4 0 2 16 4 13 1 10 9 7 9 2 7 14 3 1 9 0 2 9 3 7 1 0 9 0 9 2
7 16 9 9 13 1 0 9
19 9 13 2 9 13 2 9 13 2 9 13 2 0 9 13 2 9 13 2
9 1 10 9 13 0 9 0 9 2
17 3 2 7 13 3 2 16 3 3 2 13 1 15 9 0 9 2
14 13 15 2 16 15 13 1 0 9 9 1 0 9 2
9 13 0 9 7 13 1 9 9 2
18 13 9 10 0 9 2 16 1 15 15 9 1 0 9 3 13 3 2
5 15 13 0 9 2
8 1 0 9 13 15 10 9 2
26 14 2 16 15 15 13 3 2 7 3 2 16 15 13 0 9 2 1 15 13 2 13 7 13 9 2
5 9 15 3 13 2
19 9 15 13 1 9 0 9 0 9 1 0 9 0 10 9 1 0 9 2
12 9 2 3 15 13 2 13 2 15 7 3 2
7 1 9 1 11 2 11 2
5 7 3 1 9 2
16 13 15 2 16 13 9 1 9 1 9 7 9 4 3 13 2
11 9 9 2 7 15 15 13 2 13 9 2
13 0 14 13 9 3 1 15 2 16 1 9 13 2
21 1 10 0 9 13 15 15 2 15 15 3 13 16 3 1 11 2 7 1 9 2
28 1 9 1 11 3 15 13 2 1 15 2 15 14 13 9 2 7 1 9 15 13 2 16 15 13 3 0 2
14 0 1 0 9 7 13 15 2 15 13 0 9 3 2
14 3 0 0 9 3 13 1 10 9 9 1 0 9 2
25 1 9 0 9 1 9 7 9 1 9 14 15 15 13 9 3 0 9 2 7 10 9 13 0 2
33 0 15 13 2 1 15 13 1 10 9 2 16 1 9 13 0 16 10 0 2 1 10 9 2 16 9 1 9 13 3 1 9 2
8 7 16 4 13 3 14 0 2
19 1 10 0 1 0 9 0 9 15 3 14 13 1 9 9 0 1 9 2
50 3 1 9 2 3 9 9 11 11 13 10 0 9 2 1 15 3 13 2 16 15 3 13 1 9 2 7 7 9 1 15 13 2 15 13 2 16 0 9 9 13 13 2 7 10 9 13 13 9 2
7 16 15 3 1 15 13 2
18 16 16 4 9 1 9 13 2 13 15 2 14 13 2 14 13 2 2
5 7 3 1 15 2
19 13 3 7 9 0 9 2 3 14 2 9 2 15 13 0 9 1 9 2
24 13 10 0 9 2 16 15 1 15 3 13 0 12 9 2 13 4 1 9 3 3 1 9 2
14 9 13 3 3 14 9 2 2 2 13 15 2 9 2
11 13 15 3 0 2 16 15 3 3 13 2
4 12 7 13 2
17 16 4 13 13 9 1 9 2 13 15 15 1 9 9 0 9 2
4 13 15 15 2
4 13 15 15 2
10 13 15 15 15 2 15 13 1 9 2
37 13 15 1 11 9 1 12 2 16 4 13 7 13 2 16 15 9 4 13 2 7 13 15 15 2 14 1 0 9 9 2 0 1 9 0 9 2
11 11 2 3 2 7 11 3 1 9 1 9
4 9 13 9 9
5 11 2 11 2 2
14 1 9 9 9 15 3 1 9 0 9 13 0 9 2
19 1 9 9 13 9 3 2 16 9 9 9 13 14 9 2 7 7 9 2
25 9 1 10 9 3 13 0 9 7 13 3 1 9 7 1 15 2 16 4 1 10 9 15 13 2
22 10 9 13 7 1 15 0 2 16 3 13 2 0 9 2 13 9 1 2 9 2 2
14 1 0 9 9 3 13 0 9 1 9 14 12 9 2
13 13 3 9 9 1 9 9 2 15 13 0 9 2
7 9 13 9 1 11 0 9
5 11 2 11 2 2
24 0 9 13 9 1 0 9 0 0 0 9 7 0 9 0 9 11 11 3 1 9 0 9 2
11 13 15 15 3 0 9 1 0 0 9 2
13 11 4 13 1 9 9 0 9 7 9 0 9 2
14 0 9 15 13 1 9 9 9 0 0 9 11 11 2
24 9 15 13 1 9 2 7 1 0 9 9 2 7 16 11 11 3 13 2 16 15 11 13 2
26 11 15 2 16 15 13 2 13 9 9 9 3 2 16 11 13 2 16 15 3 7 9 2 13 2 2
12 11 11 13 9 9 9 1 12 1 12 9 2
6 1 9 13 9 1 9
5 11 2 11 2 2
30 0 9 1 0 9 13 12 0 9 9 0 9 11 11 11 2 1 10 12 0 9 11 11 2 2 9 9 1 9 2
24 13 15 1 9 1 10 0 9 1 11 7 13 2 16 15 13 2 16 3 13 9 7 9 2
8 13 3 13 10 0 0 9 2
16 3 13 7 9 2 7 10 9 2 15 1 15 13 1 9 2
21 1 9 11 11 2 13 10 9 1 9 2 15 3 13 2 13 15 7 13 9 2
9 9 3 11 11 2 13 1 9 2
1 9
2 11 12
3 12 9 12
4 12 1 9 9
4 12 9 1 15
3 12 9 9
7 12 0 9 2 12 2 2
9 12 9 13 2 0 9 1 9 12
8 12 13 9 9 2 13 9 9
2 12 11
8 12 9 1 9 2 12 2 2
10 12 9 2 7 9 2 2 2 2 2
3 12 9 9
2 12 9
4 12 9 1 9
5 12 9 1 12 9
7 12 9 0 9 2 0 9
9 12 9 1 0 9 2 12 2 2
2 12 9
2 12 9
6 12 0 2 0 2 11
4 12 12 9 9
9 12 0 9 1 9 2 12 2 2
12 12 9 0 9 2 12 2 2 2 0 0 9
2 12 9
6 12 9 2 9 2 9
12 12 0 9 2 12 2 2 2 0 0 0 9
6 12 11 2 12 2 2
6 12 9 2 9 2 9
3 12 9 11
10 12 9 1 0 9 2 0 0 2 9
2 12 9
7 12 9 2 9 2 11 11
9 12 12 2 0 2 0 9 11 12
6 12 0 2 0 2 11
2 11 12
4 12 9 2 9
11 12 1 9 1 9 2 11 11 2 11 11
6 12 9 9 1 0 9
3 12 9 9
2 12 9
3 12 9 12
3 12 0 9
3 12 11 3
2 12 9
8 12 9 0 9 2 9 9 0
2 12 9
9 12 11 9 7 9 2 12 2 2
3 12 9 9
4 12 3 3 3
5 12 9 2 7 0
3 12 1 12
3 12 9 11
5 12 0 11 2 9
3 12 9 9
2 12 9
3 12 0 9
2 12 9
4 12 0 1 11
9 12 9 1 9 2 0 0 9 9
5 12 9 9 2 9
8 12 9 1 9 2 12 2 2
3 12 9 12
6 12 3 1 11 2 11
5 12 12 9 1 9
3 12 9 11
2 11 12
4 12 0 11 9
3 12 0 11
4 12 0 11 9
3 12 0 11
2 12 9
3 12 0 9
4 12 0 11 9
3 12 11 9
2 12 9
3 12 0 9
3 12 0 9
3 12 0 9
3 12 11 11
6 12 9 9 2 12 9
6 12 9 9 2 12 9
4 12 9 1 9
12 12 0 9 9 2 12 2 2 2 0 9 9
2 12 9
4 12 9 1 9
4 12 0 9 9
2 12 3
2 12 9
3 12 11 3
2 12 9
6 12 9 2 12 2 2
3 12 9 12
4 12 9 1 11
3 12 0 9
2 12 9
4 12 11 9 3
1 9
2 11 12
1 12
3 11 11 12
2 11 12
2 9 9
36 12 9 11 2 11 2 0 9 2 12 0 9 2 0 9 2 12 0 11 2 12 2 9 2 12 0 9 2 12 9 1 9 2 12 9 3
2 9 9
44 12 11 2 12 9 2 12 11 2 12 11 2 12 11 2 0 9 2 12 9 2 12 0 9 2 9 2 12 12 9 2 9 2 12 9 2 12 12 3 1 0 11 2 9
13 1 0 9 15 3 1 11 13 9 2 15 13 9
7 11 13 9 1 9 1 11
7 11 2 11 2 11 2 2
27 9 13 9 11 11 1 9 0 9 2 16 9 11 11 2 11 2 3 13 9 2 16 11 13 1 11 2
21 11 13 13 16 9 0 9 2 1 11 7 1 9 0 9 1 9 9 3 13 2
20 11 15 3 13 11 13 1 9 9 12 2 9 2 3 15 13 16 0 9 2
13 13 15 1 9 2 1 15 9 13 9 9 11 2
30 11 13 2 16 11 3 1 0 9 11 11 11 13 1 9 9 12 2 10 9 13 11 1 10 9 2 9 1 11 2
9 11 9 1 10 9 1 11 13 2
12 13 2 16 1 11 13 1 12 9 9 9 2
8 13 15 3 7 1 0 9 2
12 11 13 2 16 1 11 13 9 1 9 9 2
16 9 1 9 11 13 12 9 2 9 14 1 9 10 9 13 2
7 9 11 2 13 0 0 9
2 11 2
26 0 9 13 0 9 9 0 9 2 0 9 11 2 10 0 9 13 11 7 15 13 9 12 9 0 2
12 9 13 2 16 10 9 13 3 13 0 9 2
27 1 9 0 0 9 7 9 13 2 16 9 9 13 9 15 2 16 11 13 0 9 0 9 1 9 9 2
10 16 11 13 1 11 2 0 9 15 13
1 9
18 9 1 15 2 16 11 4 13 0 9 16 3 11 2 15 13 13 2
23 0 2 7 3 0 2 0 9 15 1 9 13 0 9 2 0 0 9 15 13 13 11 2
20 0 9 15 9 11 13 0 9 2 3 11 13 7 3 13 1 9 0 9 2
13 3 15 13 11 1 0 9 2 3 13 9 9 2
26 3 15 13 0 9 2 0 11 2 2 15 13 9 2 16 10 9 7 9 1 0 9 13 0 9 2
28 1 0 9 13 1 9 9 7 9 7 1 10 0 2 9 2 1 0 9 13 10 9 2 3 0 9 13 2
12 3 1 10 9 1 9 9 13 11 7 11 2
21 3 1 10 0 9 13 11 14 0 9 2 3 13 10 9 2 14 3 3 13 2
19 13 0 2 16 0 7 0 13 9 10 9 2 15 13 1 9 0 9 2
19 13 2 3 4 13 13 1 0 3 0 3 0 2 16 13 1 9 0 2
31 9 1 9 13 0 0 9 11 2 7 16 3 1 11 2 0 11 2 13 1 9 1 10 0 9 3 3 1 12 9 2
28 1 9 0 9 1 9 0 9 13 7 9 2 16 0 9 13 1 3 0 9 0 9 16 3 3 0 9 2
19 7 3 2 0 2 9 2 15 13 13 9 1 11 7 15 15 13 9 2
30 0 9 11 2 15 3 13 1 11 1 9 0 9 1 9 1 3 0 0 9 2 4 13 1 3 0 9 3 9 2
12 16 4 13 16 11 2 13 15 16 3 13 2
6 9 11 13 12 9 9
2 11 2
41 9 1 11 2 12 2 2 15 15 3 1 9 13 1 9 11 2 12 2 7 13 1 9 9 1 9 2 13 12 9 9 2 16 4 13 13 10 0 0 9 2
14 0 9 9 1 11 13 0 9 14 1 9 9 9 2
23 9 11 13 3 1 10 0 9 1 0 9 2 16 11 13 16 9 9 11 1 9 11 2
23 9 1 9 1 0 0 9 13 2 16 9 9 7 9 1 11 13 1 0 9 1 9 2
19 9 11 2 16 4 15 13 13 9 2 4 15 1 9 9 13 3 13 2
13 9 9 11 13 12 9 2 1 12 9 0 9 2
9 10 9 13 14 1 12 9 3 2
16 3 12 9 9 3 13 11 1 9 2 9 2 9 7 9 2
24 9 12 9 9 13 13 1 9 0 0 9 1 0 11 7 0 12 9 1 10 9 0 9 2
6 1 11 13 12 0 9
2 11 2
23 1 12 9 9 0 9 3 13 1 0 9 11 1 9 0 9 7 9 11 1 0 9 2
38 10 9 4 13 1 0 0 9 2 15 13 13 1 0 9 1 9 1 9 1 9 2 16 9 11 4 13 9 1 9 0 9 9 1 0 0 9 2
28 9 9 11 13 2 16 11 13 0 9 13 9 7 13 0 9 0 1 12 9 0 0 9 1 0 0 9 2
32 0 0 9 13 2 16 9 9 13 15 0 1 0 9 9 1 0 9 1 11 7 1 9 13 9 0 0 9 11 11 11 2
29 3 3 7 13 9 9 0 9 11 11 11 1 9 9 12 0 9 9 12 2 16 1 0 9 11 13 12 9 2
24 9 0 0 9 13 9 0 9 1 9 11 2 15 13 1 9 2 3 3 10 9 13 0 9
14 1 11 13 11 1 12 9 7 11 3 1 12 9 2
7 11 13 13 1 12 9 2
8 9 13 9 11 1 12 9 2
37 3 9 13 1 11 0 2 9 2 11 2 15 13 1 0 9 1 0 9 2 11 1 12 2 11 1 12 2 11 1 12 7 9 1 12 9 2
5 11 13 9 7 9
2 11 2
30 16 1 9 9 9 1 0 9 11 13 3 12 9 9 2 0 9 13 13 14 1 0 9 7 9 13 1 0 9 2
26 1 9 0 11 2 15 3 9 13 13 9 0 11 1 9 2 13 4 0 0 9 11 13 0 9 2
33 2 11 13 3 1 0 9 15 2 15 3 3 13 1 0 9 2 2 13 3 9 11 11 2 0 9 0 0 9 2 11 2 2
34 13 2 16 1 9 2 3 13 9 1 15 2 15 13 3 9 0 9 2 13 9 2 2 15 11 7 9 1 0 0 9 13 2 2
22 9 2 15 13 1 9 3 12 9 9 1 9 7 9 2 13 13 9 1 0 9 2
8 3 13 13 9 9 7 9 2
13 7 3 9 13 1 9 15 2 15 4 9 13 2
28 2 9 13 3 2 3 0 2 2 13 9 2 11 11 2 9 7 0 0 9 2 15 3 13 1 9 11 2
17 2 13 9 3 1 10 9 2 3 13 10 9 3 1 9 2 2
23 9 0 9 2 0 1 0 9 2 0 9 7 0 9 2 3 11 13 9 2 3 13 2
15 16 4 15 9 11 13 1 9 9 2 13 13 0 9 2
39 0 9 15 3 13 1 15 2 16 10 9 15 13 13 9 1 9 9 0 9 2 7 15 3 2 16 11 4 13 11 1 12 1 12 2 0 9 2 2
5 9 1 9 2 12
8 9 1 11 2 3 0 9 9
2 11 2
22 0 9 2 0 9 7 9 1 11 2 9 11 7 11 7 0 2 0 9 0 9 2
4 9 7 9 2
17 15 13 11 2 0 0 9 9 2 15 0 9 13 13 9 9 2
18 13 1 11 13 3 0 2 1 11 7 11 7 13 0 15 3 13 2
52 3 1 9 2 7 3 2 16 11 13 10 9 1 9 3 13 2 1 11 13 0 15 13 9 2 7 15 13 14 3 9 2 7 3 3 9 2 0 0 9 1 0 9 2 7 3 2 3 13 13 9 2
34 1 0 0 9 4 1 9 12 2 0 2 1 15 13 9 1 9 2 12 9 0 9 13 2 3 3 1 9 1 9 1 0 9 2
38 16 13 3 9 9 9 7 13 9 0 9 2 13 3 9 1 9 1 11 3 13 2 0 9 13 7 0 13 9 9 0 2 16 13 14 0 9 2
22 1 9 7 9 13 0 2 7 0 9 13 2 16 4 1 9 1 11 13 0 9 2
34 0 9 7 11 13 9 1 0 9 9 0 9 2 7 7 4 15 13 13 2 16 13 0 13 0 9 2 15 13 1 11 3 0 2
12 9 3 3 13 9 2 16 13 9 1 9 2
30 0 9 1 9 13 9 1 15 12 7 12 9 2 0 0 9 1 12 7 12 2 9 1 0 9 1 9 3 3 2
44 9 0 0 9 1 9 1 9 3 13 3 0 2 3 13 0 9 2 7 13 0 13 1 3 0 9 2 15 9 3 13 2 7 13 3 0 2 15 15 0 9 13 13 2
16 15 7 2 15 15 10 15 13 2 15 11 13 16 0 9 2
27 1 15 0 0 9 7 1 9 1 15 13 0 9 2 3 3 0 9 2 9 2 0 9 2 15 3 2
35 13 15 1 15 13 2 13 15 13 1 9 7 1 9 2 7 3 15 13 0 9 1 9 1 9 1 9 7 1 9 1 9 7 9 2
23 3 13 3 13 9 1 0 9 0 9 1 10 9 1 9 1 9 3 16 1 0 9 2
27 16 13 1 9 2 1 9 13 13 3 3 0 9 2 3 0 9 13 1 9 1 9 12 7 12 9 2
19 9 13 3 1 9 2 1 9 7 9 2 9 13 3 3 0 16 9 2
33 3 9 9 2 9 7 9 2 2 9 1 9 1 9 2 13 1 0 2 3 1 12 9 0 9 15 10 9 13 1 12 9 2
32 9 13 3 13 13 2 7 3 13 11 0 9 2 1 2 0 2 2 16 0 9 14 1 3 0 7 0 9 1 0 9 2
12 0 13 3 13 15 1 9 1 3 0 9 2
35 7 1 0 9 13 9 2 3 15 1 9 9 0 0 9 9 9 13 2 7 13 3 15 15 13 9 1 0 9 7 1 9 0 9 2
30 1 9 1 11 7 13 13 9 0 9 2 11 2 11 2 11 7 11 2 1 0 2 3 16 15 13 9 1 9 2
24 1 0 0 9 13 1 11 3 0 0 2 0 7 0 9 2 1 9 13 0 0 0 9 2
23 3 13 7 1 1 9 3 0 15 13 9 2 15 13 3 1 9 7 1 0 0 9 2
10 1 9 1 11 13 1 11 13 9 2
18 13 15 3 12 9 1 9 7 3 3 2 1 9 1 9 2 2 2
3 0 9 2
5 11 13 9 7 9
5 9 1 9 2 12
26 11 11 2 12 1 9 9 11 2 13 3 1 9 2 16 9 9 1 0 9 13 3 1 12 9 2
30 7 9 15 13 2 15 15 13 1 9 1 9 7 1 9 2 10 0 9 13 0 1 9 2 16 15 9 13 3 2
23 2 15 13 9 1 15 2 2 13 9 2 11 11 2 16 13 1 12 9 1 0 9 2
18 0 9 3 4 13 1 0 9 9 2 16 4 3 3 13 1 9 2
16 9 4 1 0 9 2 3 13 9 2 13 3 16 12 9 2
24 9 11 7 11 13 2 16 3 13 13 7 13 9 9 1 9 7 13 2 16 15 13 9 2
11 1 15 13 0 7 9 9 9 7 9 2
12 13 9 9 1 0 9 2 16 4 13 9 2
20 0 9 0 9 4 13 0 9 9 9 7 9 1 9 13 0 1 9 9 2
21 13 14 13 1 0 9 7 10 9 2 3 1 9 13 3 16 12 9 7 9 2
13 16 13 9 9 7 9 9 2 9 7 9 13 2
28 2 13 2 16 15 3 13 15 13 9 1 12 12 9 2 9 15 3 13 1 10 9 2 2 13 9 11 2
16 2 3 15 13 16 1 0 9 2 3 13 1 9 12 9 2
8 7 13 15 3 1 9 2 2
7 9 9 11 1 9 15 13
21 0 9 2 0 0 9 1 0 3 1 0 9 2 13 3 3 9 16 9 9 2
17 14 7 15 13 1 9 0 9 15 2 15 13 13 1 0 9 2
29 3 13 15 12 9 2 3 4 1 11 11 13 9 0 9 2 11 2 16 9 9 0 9 3 0 9 9 11 2
27 0 9 11 13 13 1 9 0 9 7 9 1 9 1 0 9 2 13 9 0 9 7 0 9 1 9 2
25 1 10 3 0 9 4 9 7 9 9 11 1 0 9 7 0 9 13 0 3 0 7 0 9 2
21 3 1 9 13 9 0 9 14 0 1 9 9 2 7 13 9 1 15 7 13 2
22 3 3 3 0 9 4 13 10 0 9 7 0 9 13 13 1 0 0 9 1 9 2
46 0 0 7 0 9 2 0 0 0 9 7 0 9 2 3 1 0 0 9 2 1 12 9 1 9 2 7 0 0 7 0 9 0 9 13 1 11 10 0 9 1 3 3 0 9 2
46 0 11 13 3 0 0 9 2 3 0 7 0 9 0 9 1 9 0 0 9 0 9 9 7 1 0 9 9 9 2 15 3 13 10 0 9 1 9 9 9 7 1 15 0 9 2
31 13 7 3 9 2 16 9 0 9 15 3 2 16 3 13 13 15 15 2 16 3 13 9 1 0 9 2 3 1 9 2
26 14 0 9 2 0 9 0 9 2 7 0 9 2 9 0 9 9 7 0 9 2 15 3 3 13 2
20 12 2 3 7 0 9 1 9 2 0 9 2 13 9 1 0 9 0 9 2
49 0 9 1 10 9 13 9 0 0 9 1 9 9 0 2 0 9 1 9 2 15 15 13 13 9 1 9 9 0 7 0 9 9 2 15 15 0 9 13 1 0 9 7 2 9 9 2 11 2
26 0 9 7 9 0 0 7 3 0 9 2 15 3 13 0 9 2 13 3 0 9 9 9 0 9 2
28 1 15 13 0 2 16 4 11 13 0 9 7 3 13 0 7 0 0 9 2 15 13 0 9 1 0 9 2
29 3 1 15 15 13 3 13 0 9 0 9 1 11 16 1 3 0 7 2 3 0 2 9 2 0 1 9 0 2
45 0 9 9 2 1 9 1 0 9 0 9 2 15 13 3 0 1 9 0 0 9 2 4 15 13 13 1 9 0 9 0 9 9 9 0 9 2 15 4 13 1 9 0 9 2
30 14 3 15 3 13 2 2 13 9 9 7 13 15 1 12 9 2 13 15 13 0 9 7 13 15 1 0 9 2 2
16 9 11 13 3 0 7 10 0 7 0 9 13 3 16 0 2
32 1 9 1 15 2 15 15 10 9 13 2 16 2 0 9 2 13 9 0 9 2 13 1 0 9 2 15 13 1 0 9 2
2 11 11
4 9 13 9 9
6 9 9 1 11 12 9
2 11 2
31 0 9 0 0 9 2 15 1 9 13 16 0 9 0 9 9 1 0 9 1 0 11 2 4 7 4 13 12 0 9 2
14 1 9 4 7 4 13 9 2 9 2 9 7 9 2
15 10 9 4 13 1 9 1 11 2 11 2 11 7 11 2
4 11 13 9 11
2 11 2
19 12 9 3 13 1 9 1 11 2 16 11 13 0 9 2 15 13 9 2
8 13 15 0 9 0 9 9 2
18 1 10 9 9 13 1 9 11 2 0 9 1 11 2 15 13 11 2
6 0 9 3 9 13 2
7 0 9 15 13 1 9 11
2 11 2
37 0 9 11 1 11 11 11 11 3 13 1 0 9 11 2 16 4 15 13 1 9 0 11 11 11 2 15 15 3 1 0 0 9 13 0 9 2
20 12 9 13 13 9 9 9 2 15 13 3 1 9 1 11 2 9 9 2 2
4 12 0 9 13
2 11 2
29 1 0 9 3 4 13 12 0 9 0 0 9 1 0 9 1 0 9 7 9 1 9 2 15 9 13 13 9 2
16 13 15 0 9 9 0 1 11 1 0 9 1 0 0 9 2
5 11 13 13 0 9
3 0 11 2
17 9 11 13 13 12 0 0 9 2 16 3 11 13 9 0 9 2
9 13 15 3 1 0 11 9 11 2
14 9 13 4 13 2 16 4 11 13 13 9 0 9 2
5 9 0 9 1 11
2 11 2
32 9 0 0 9 13 15 0 9 7 0 9 2 15 13 1 9 0 9 2 16 4 13 9 0 0 7 0 9 1 10 9 2
15 13 15 3 0 9 11 2 11 1 9 1 3 0 9 2
38 9 9 0 9 13 3 2 16 0 9 1 9 1 10 9 13 0 0 9 11 11 2 0 1 9 9 1 0 0 9 11 1 0 9 11 2 9 2
14 3 15 1 11 2 11 13 7 13 2 0 2 9 2
38 0 9 1 9 1 3 0 9 3 13 2 16 9 0 9 13 13 3 1 9 1 0 9 1 9 9 9 0 9 7 9 9 2 15 13 1 9 2
22 1 0 9 3 1 9 11 2 11 13 0 9 11 2 0 9 11 7 9 0 9 2
7 11 7 11 13 1 11 11
2 11 2
31 11 7 11 2 15 16 0 9 1 0 0 9 4 13 3 1 11 2 4 13 10 9 1 9 9 1 9 9 0 9 2
27 13 15 3 1 11 0 9 9 11 11 2 15 15 1 9 11 11 13 9 12 0 9 2 9 12 2 2
16 1 0 9 12 9 13 11 1 9 1 10 0 9 11 11 2
11 9 15 1 10 9 13 1 0 0 9 2
25 2 11 13 9 1 9 9 2 15 13 10 9 2 7 15 13 3 12 2 2 13 11 1 9 2
21 13 2 16 11 15 13 1 11 2 13 7 13 2 2 7 2 3 15 13 2 2
23 11 1 9 11 3 13 0 9 11 7 11 1 9 9 2 16 11 7 11 13 3 9 2
51 11 3 13 1 15 2 16 4 0 9 1 10 0 9 1 11 4 1 9 9 12 0 3 1 9 1 11 13 2 7 13 2 16 0 9 9 12 2 1 15 15 13 1 9 10 9 2 13 1 9 2
18 1 9 10 9 13 9 0 9 9 11 11 2 16 15 1 9 13 2
22 0 9 11 11 3 13 1 11 2 16 4 15 13 1 9 0 9 12 0 9 9 2
6 11 13 1 9 9 2
21 1 0 9 9 9 12 15 13 11 13 3 3 2 3 0 9 9 12 3 13 2
11 1 9 11 15 1 9 1 11 3 13 2
28 12 1 9 9 13 1 0 9 9 11 11 9 2 16 9 9 12 14 13 11 0 9 1 9 12 9 9 2
10 9 13 4 13 1 9 0 0 9 2
31 10 9 4 13 13 1 12 9 0 9 1 9 12 2 12 9 1 0 9 7 12 9 1 0 9 7 0 0 0 9 2
19 0 12 9 4 13 0 9 0 0 9 1 9 9 9 1 9 10 9 2
20 11 1 9 13 9 12 9 1 9 7 0 9 7 12 9 9 1 0 9 2
10 9 9 12 13 1 11 13 0 9 11
2 11 2
42 0 9 12 0 0 9 9 2 9 12 2 15 3 1 10 0 9 13 1 9 0 9 11 7 13 2 16 13 10 9 9 1 11 2 15 4 4 13 1 9 9 2
17 1 0 0 9 3 13 11 2 11 7 11 1 9 0 9 9 2
16 9 9 12 1 15 3 13 9 1 9 13 1 11 0 9 2
30 15 4 13 13 9 9 9 9 2 12 2 1 15 13 4 1 0 9 1 11 13 12 9 2 0 9 0 9 11 2
10 9 9 12 13 1 9 9 9 9 2
13 10 9 13 9 11 7 11 1 9 1 10 9 2
21 0 9 1 9 9 4 12 9 13 0 9 2 15 4 13 10 0 9 1 9 2
12 2 13 11 7 11 2 2 2 9 2 12 2
7 0 9 13 1 11 7 11
2 11 2
23 0 9 0 9 11 11 7 10 0 0 9 11 11 3 13 1 11 0 9 1 9 9 2
16 11 11 13 2 16 10 9 13 1 0 0 9 0 1 11 2
22 9 13 2 16 4 9 0 1 11 1 11 4 13 1 11 2 16 3 1 11 13 2
42 1 9 2 16 15 4 9 13 1 9 11 2 11 2 11 13 2 16 4 3 13 4 13 0 9 1 11 2 7 13 9 2 16 15 13 0 9 13 7 1 11 2
6 0 9 1 9 1 9
2 11 2
14 0 9 3 13 2 16 3 13 1 9 1 9 9 2
15 13 9 2 15 1 0 9 13 13 9 9 2 0 9 2
11 13 7 2 16 9 3 13 1 9 15 2
16 9 4 13 1 12 0 9 2 1 15 15 4 9 9 13 2
25 0 9 13 9 2 15 9 13 9 7 13 3 1 0 9 2 0 9 9 2 3 13 0 9 2
3 0 9 9
3 9 1 9
3 0 9 9
26 1 9 2 15 13 10 9 0 13 9 9 2 13 7 9 2 1 9 0 1 0 9 1 0 9 2
15 9 13 7 9 9 2 1 9 13 9 9 1 0 9 2
15 13 0 1 9 2 7 13 3 9 1 9 0 0 9 2
23 13 15 13 7 16 0 9 1 9 2 13 1 9 9 9 7 9 2 0 7 0 9 2
14 16 4 15 0 9 1 9 13 2 13 9 3 13 2
19 0 13 1 15 0 9 7 0 2 0 7 0 9 1 9 1 12 9 2
25 9 15 13 13 1 9 1 0 9 2 0 7 0 2 16 15 1 15 13 1 9 13 0 9 2
24 13 15 9 13 0 2 13 15 1 0 9 7 9 2 7 13 9 15 13 1 10 0 9 2
10 0 9 1 12 2 1 12 2 12 2
15 13 2 14 1 9 7 9 13 3 2 9 1 12 9 2
11 9 4 13 1 9 2 1 9 1 9 2
1 9
55 0 9 11 13 0 0 9 1 9 9 0 9 1 9 9 9 2 0 9 2 9 7 9 0 9 2 9 2 9 1 0 9 11 1 0 9 12 2 12 12 11 2 0 9 1 0 9 4 13 3 1 12 2 9 2
1 9
2 11 2
6 9 12 2 12 2 12
12 11 11 1 0 9 0 9 11 2 13 11 2
4 0 1 9 2
5 1 12 2 12 2
24 9 9 7 9 2 0 9 1 9 7 1 9 1 9 11 11 2 11 2 1 12 2 12 2
1 9
2 11 2
18 0 9 2 9 2 9 2 0 9 2 2 0 9 1 0 9 0 9
2 11 2
29 12 9 2 12 9 7 0 9 1 0 9 1 9 11 11 2 0 9 2 12 2 12 2 1 12 2 12 2 2
2 11 2
15 11 11 1 9 11 11 9 9 2 1 12 2 12 2 2
2 11 2
13 9 11 11 1 9 9 2 1 12 2 12 2 2
2 11 2
21 9 1 9 1 9 9 2 11 11 2 11 11 2 2 2 1 12 2 12 2 2
2 11 2
36 9 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 7 11 2 11 2 11 1 9 1 0 9 2 1 12 2 12 2 2
2 11 2
14 1 0 0 9 1 9 9 2 1 12 2 12 2 2
2 11 2
16 0 9 0 11 1 0 9 0 9 2 1 12 2 12 2 2
2 11 2
36 1 9 7 9 2 9 0 9 1 9 12 7 12 2 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 2 1 12 2 12 2 2
4 11 1 11 2
21 9 2 9 11 2 11 7 11 2 11 1 9 1 9 2 1 12 2 12 2 2
4 11 1 11 2
18 9 7 9 1 9 11 1 9 9 2 11 2 1 12 2 12 2 2
4 11 1 11 2
15 9 11 11 1 9 9 2 11 2 1 12 2 12 2 2
5 0 9 1 11 2
6 9 12 2 12 2 12
24 11 11 2 9 2 9 2 9 1 0 9 2 0 9 11 11 2 2 1 12 2 12 2 2
5 0 9 1 11 2
8 9 9 2 0 9 1 0 9
5 0 9 1 11 2
20 9 1 11 2 0 9 1 0 9 2 11 2 11 2 11 2 11 0 2 2
5 0 9 1 11 2
29 0 9 2 9 2 9 2 9 11 11 2 11 11 2 11 11 7 11 11 1 0 9 2 1 12 2 12 2 2
5 0 9 1 11 2
14 11 11 2 9 1 0 9 2 1 12 2 12 2 2
6 0 11 2 11 2 2
19 11 11 7 9 0 9 7 9 9 1 9 9 2 1 12 2 12 2 2
4 11 1 11 2
48 0 9 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 1 9 1 9 2 1 12 2 12 2 2
2 11 2
25 9 12 2 12 2 9 9 11 11 2 9 1 9 1 9 9 0 9 2 1 12 2 12 2 2
2 11 2
20 11 11 2 0 9 1 0 9 12 2 9 0 9 2 1 12 2 12 2 2
2 11 2
13 0 9 0 9 7 9 12 2 9 1 9 0 9
2 0 9
2 11 2
18 13 1 0 9 1 3 0 0 9 9 11 2 1 12 2 12 2 2
2 11 2
14 13 9 0 9 1 9 11 2 1 12 2 12 2 2
4 9 1 11 2
14 0 9 2 0 2 0 9 9 1 9 1 9 0 9
2 11 2
6 9 12 2 12 2 12
24 11 11 2 0 9 1 9 9 1 0 9 2 0 9 11 11 2 2 1 12 2 12 2 2
3 0 11 2
9 0 0 9 1 9 2 1 9 2
2 11 2
22 9 1 9 2 9 9 2 11 11 11 11 13 1 9 9 2 1 12 2 12 2 2
1 9
2 11 2
13 12 9 0 9 1 9 2 1 12 2 12 2 2
2 11 2
23 11 7 9 2 9 7 9 9 9 12 2 12 1 0 9 0 0 9 2 9 2 9 2
2 11 2
17 9 0 11 2 0 9 9 1 0 9 2 1 12 2 12 2 2
2 11 2
14 9 0 0 9 1 0 9 2 1 12 2 12 2 2
2 11 2
16 9 9 9 1 0 9 0 0 9 2 1 12 2 12 2 2
2 11 2
29 0 11 1 0 9 0 9 9 9 11 2 0 9 0 9 2 9 11 2 11 2 2 2 1 12 2 12 2 2
2 11 2
15 9 1 9 9 0 1 0 9 2 1 12 2 12 2 2
2 11 2
18 0 9 1 0 9 2 0 9 2 0 9 2 0 9 2 0 9 2
2 11 2
25 11 2 11 7 12 2 9 0 0 9 1 11 1 9 12 1 9 11 2 1 12 2 12 2 2
4 11 1 11 2
15 9 1 9 0 9 1 0 9 2 1 12 2 12 2 2
4 11 1 11 2
25 13 15 15 1 9 1 0 9 2 1 12 2 9 9 9 11 2 2 2 1 12 2 12 2 2
2 11 2
26 9 9 0 9 0 12 2 1 9 2 1 9 9 0 9 1 11 2 2 2 1 12 2 12 2 2
2 11 2
12 0 0 9 1 9 2 1 12 2 12 2 2
3 0 11 2
16 0 9 1 9 11 2 11 2 11 2 1 12 2 12 2 2
3 0 9 2
19 9 11 1 0 9 1 0 9 2 1 0 9 2 1 12 2 12 2 2
3 0 9 2
14 9 1 0 9 1 0 9 2 1 12 2 12 2 2
2 0 9
2 11 2
6 9 12 2 12 2 12
10 11 11 1 9 0 9 2 13 11 2
2 11 2
6 9 12 2 12 2 12
29 9 9 2 1 0 9 1 0 9 1 0 9 11 2 9 1 11 1 12 2 12 2 1 9 9 0 9 12 2
2 11 2
6 9 12 2 12 2 12
21 9 1 11 2 9 9 0 0 9 1 0 9 11 2 1 0 9 1 0 9 2
1 11
6 9 12 2 12 2 12
11 3 14 2 9 0 0 9 1 0 9 11
2 11 2
5 0 9 2 11 2
8 0 9 12 1 9 1 9 2
6 9 12 2 12 2 12
2 11 11
8 11 2 1 11 1 11 2 2
10 9 9 11 12 1 0 9 9 9 2
6 9 12 2 12 2 12
4 9 1 0 11
6 9 12 2 12 2 12
3 9 1 11
3 9 0 9
26 11 12 2 12 2 9 1 9 7 9 2 9 11 2 11 2 0 12 2 12 12 11 12 2 9 2
10 11 11 2 13 15 2 9 2 2 2
5 2 9 11 2 11
12 11 11 2 11 2 9 1 9 2 12 2 2
4 2 11 11 2
29 9 2 0 9 2 9 2 12 2 11 11 2 11 2 2 9 2 9 2 9 2 1 0 9 12 2 12 12 11
26 9 9 2 9 1 9 7 0 9 2 9 2 12 2 11 11 2 2 9 2 0 12 2 11 12 2
8 11 11 2 9 2 9 11 2
8 11 11 2 9 2 11 11 2
9 9 0 0 9 2 0 9 11 2
9 11 1 0 9 2 0 9 11 2
10 9 11 1 0 9 2 0 9 11 2
1 9
6 0 9 1 0 9 2
17 9 13 1 9 2 11 3 2 0 12 2 12 2 12 12 11 2
23 13 13 14 9 2 15 4 1 0 9 13 1 9 2 7 2 12 9 1 0 9 9 2
5 0 9 2 9 11
6 9 12 2 12 2 12
2 11 12
33 9 11 9 9 1 0 9 9 11 9 2 11 1 0 9 9 2 1 10 9 9 13 1 9 11 2 11 1 9 9 1 11 2
6 9 12 2 12 2 12
2 11 12
18 9 2 13 7 13 2 0 9 2 9 9 2 0 9 1 0 9 2
6 9 12 2 12 2 12
2 11 12
5 11 9 2 2 2
12 2 1 9 0 9 1 9 2 12 1 9 2
6 9 11 11 2 12 9
3 0 9 2
12 12 7 12 9 1 0 9 2 9 2 9 2
4 12 2 12 12
6 9 2 9 2 9 2
15 12 0 9 2 9 2 9 2 2 9 1 0 9 1 11
3 12 0 9
10 12 2 12 0 9 2 9 2 9 2
4 12 2 12 9
10 12 0 9 2 9 2 9 2 9 2
11 12 2 12 4 15 13 2 9 0 9 2
9 12 9 1 9 2 9 1 9 2
4 9 0 9 2
1 9
4 9 0 9 2
49 0 9 2 16 0 9 13 9 9 1 9 2 7 7 4 9 1 9 7 9 2 15 13 3 0 9 2 13 2 15 1 9 9 0 9 0 9 11 1 9 0 9 1 0 9 13 13 0 2
7 0 9 9 13 12 5 2
52 3 3 13 9 0 9 2 1 12 5 2 2 16 3 1 15 13 0 12 5 9 2 7 15 14 1 9 1 11 7 0 11 2 7 13 15 9 9 0 9 1 12 5 2 15 15 13 1 9 12 5 2
13 1 12 5 13 7 9 9 2 15 13 9 9 2
6 7 9 13 3 0 2
42 1 0 9 3 4 1 9 13 9 1 11 2 7 16 15 13 3 14 0 2 13 15 3 9 9 2 15 15 7 1 11 13 9 9 2 15 13 12 0 0 9 2
11 13 3 9 11 2 9 0 9 4 13 2
45 3 13 9 0 9 14 1 9 0 0 9 1 9 0 11 2 11 1 12 5 2 11 1 12 5 2 2 1 11 2 11 7 9 0 11 2 1 0 9 7 1 9 0 9 2
32 1 0 9 13 9 0 2 11 12 5 2 11 12 5 2 1 11 12 5 2 2 0 13 14 1 11 2 11 7 1 11 2
17 1 0 11 2 11 2 11 2 11 2 11 7 11 3 9 13 2
20 1 0 9 14 11 7 0 9 1 11 13 9 0 1 0 11 9 9 9 2
15 3 3 15 7 0 9 13 13 9 1 9 2 13 9 2
25 9 9 13 2 7 13 1 9 1 0 9 2 15 3 13 14 1 0 0 9 2 3 13 3 2
9 7 0 9 13 0 13 0 9 2
4 9 16 0 9
13 2 1 9 0 9 2 9 11 11 1 9 1 9
2 11 2
33 9 2 9 7 9 11 11 2 12 2 1 15 13 3 1 0 9 11 2 2 2 9 1 0 9 1 11 9 14 1 11 9 2
21 0 0 9 1 0 9 2 9 11 11 11 2 15 1 9 0 9 13 0 9 2
32 2 1 0 9 15 13 2 16 15 1 9 13 3 0 9 2 1 0 2 16 13 1 9 2 2 13 0 9 11 2 11 2
22 7 3 1 0 9 0 9 11 11 15 13 9 13 1 9 9 1 0 9 0 9 2
32 11 13 7 1 9 0 9 11 7 1 9 1 9 2 3 3 13 9 1 11 2 11 2 11 2 13 1 0 9 0 9 2
8 1 12 13 0 9 0 9 2
8 13 15 3 12 1 10 9 2
22 2 13 4 15 1 9 0 9 2 1 15 13 13 2 16 15 3 15 4 13 13 2
17 13 15 13 10 9 3 3 2 13 9 9 7 9 9 1 9 2
8 3 2 1 10 9 3 13 2
11 16 4 15 3 13 13 9 15 0 2 2
14 13 15 2 16 15 9 9 13 16 3 0 9 13 2
10 2 13 2 16 15 13 9 9 2 2
15 10 9 2 3 10 0 9 2 4 15 13 9 0 9 2
7 13 3 1 9 0 9 2
3 2 13 2
28 1 9 13 3 9 2 15 15 13 2 16 4 15 13 13 2 2 16 16 2 15 13 1 15 15 1 15 2
17 10 9 13 1 15 1 9 0 2 9 4 13 9 1 9 2 2
9 1 15 15 1 9 10 9 13 2
20 2 0 4 13 1 9 9 11 11 2 11 2 11 2 11 7 11 11 2 2
13 13 1 15 11 9 2 15 9 13 2 7 13 2
14 2 13 11 3 3 12 9 2 10 9 4 15 13 2
12 13 7 3 0 2 16 13 1 0 9 2 2
8 15 15 3 1 9 9 13 2
17 2 9 13 0 9 9 2 15 15 1 0 9 13 3 15 13 2
33 13 15 7 9 9 9 2 13 1 10 9 2 13 1 9 2 9 2 15 15 2 13 2 14 0 7 0 2 3 13 1 9 2
20 9 3 13 1 9 9 7 13 2 3 13 3 0 9 2 14 2 14 2 2
8 0 13 10 9 7 9 9 2
9 13 15 2 16 13 9 16 15 2
21 2 9 13 3 2 16 13 15 3 2 16 13 15 2 15 13 2 13 7 13 2
10 13 15 2 3 3 15 13 9 9 2
19 16 4 13 2 3 10 0 9 13 9 13 2 13 4 15 1 9 15 2
20 1 12 9 1 10 0 9 15 12 3 13 0 9 2 3 0 12 9 9 2
12 13 15 15 0 2 3 3 13 15 1 9 2
24 13 4 15 1 15 9 9 11 2 0 7 0 9 10 0 9 2 7 15 15 15 13 2 2
1 9
25 9 1 9 2 0 9 1 9 11 11 2 13 9 0 9 1 0 9 1 11 1 12 2 9 2
6 9 9 1 12 9 2
11 9 11 11 1 0 9 13 1 12 9 2
22 9 11 11 0 9 4 13 1 12 9 1 0 9 1 11 7 13 1 12 2 9 2
5 9 3 11 11 2
18 11 2 0 0 9 1 9 2 0 9 0 9 2 4 13 9 12 2
20 9 0 1 9 2 9 7 9 2 0 1 9 0 9 2 13 1 9 9 2
19 9 1 15 13 7 11 11 2 15 11 13 9 12 1 0 9 0 9 2
15 1 10 9 0 0 9 13 2 2 2 10 9 13 11 2
3 2 11 2
12 0 9 2 9 2 6 9 2 0 9 2 2
36 2 0 9 0 9 13 1 11 1 0 9 1 12 2 9 9 2 15 1 9 7 0 9 11 2 11 2 11 13 9 11 2 11 2 11 2
16 9 13 1 15 2 1 15 15 11 13 13 1 9 10 9 2
20 9 1 9 1 0 9 9 2 7 9 7 9 1 9 0 9 13 0 9 2
6 9 13 1 12 9 2
3 2 11 2
6 9 11 2 13 3 11
33 1 0 2 3 0 9 0 0 9 11 0 9 1 0 9 1 9 4 15 10 9 13 2 15 13 9 1 0 9 7 9 9 2
11 2 15 2 11 13 3 0 0 9 2 2
7 4 3 13 0 0 9 2
7 2 3 2 1 0 9 2
4 13 3 11 2
17 1 10 0 9 4 13 12 0 0 9 2 7 1 0 9 2 2
7 13 1 0 9 0 13 2
8 2 3 0 2 13 0 9 2
10 1 11 3 13 2 16 13 3 2 2
3 9 1 11
2 11 2
19 0 9 11 11 13 3 1 9 0 0 9 9 1 9 0 9 11 11 2
13 1 12 2 9 13 9 3 16 3 1 12 9 2
26 0 9 1 12 9 2 0 9 2 0 0 9 7 9 13 1 12 1 0 2 15 15 3 3 13 2
16 9 11 15 13 11 11 2 0 11 9 10 0 9 11 11 2
4 9 7 0 9
7 0 9 11 11 1 0 9
29 0 10 9 4 3 13 2 7 11 11 13 12 1 10 2 15 13 10 9 13 0 9 7 3 13 9 0 9 2
20 13 15 3 7 1 9 10 0 0 9 0 2 15 3 13 1 0 9 11 2
16 9 15 1 15 13 0 12 9 2 15 13 1 9 0 14 2
23 1 9 3 13 9 9 1 0 9 1 9 0 9 11 2 7 3 0 9 0 9 13 2
33 0 3 13 3 0 16 0 7 0 0 9 1 9 0 7 0 9 2 7 9 0 9 7 0 9 1 0 9 15 13 1 15 2
23 0 9 13 1 9 9 13 0 13 13 1 15 1 13 1 13 0 14 1 0 0 9 2
29 7 13 15 14 0 9 2 7 3 0 9 1 13 1 13 15 7 0 9 9 1 0 1 0 9 7 3 15 2
35 1 9 0 1 9 13 0 3 9 12 0 9 0 9 0 9 2 11 11 7 11 11 2 15 1 9 13 2 3 9 1 9 1 9 2
23 10 15 7 13 14 9 1 9 2 15 13 0 0 9 2 3 0 2 3 3 3 0 2
34 13 0 9 2 13 0 11 1 9 14 2 7 1 9 9 9 1 11 3 13 2 14 13 3 2 14 11 11 13 11 11 2 11 2
44 9 15 7 12 0 13 2 13 2 14 0 0 9 2 0 9 1 3 15 13 0 9 0 3 1 9 7 9 0 9 2 16 1 9 0 1 0 9 3 13 9 14 9 2
27 9 13 9 1 0 9 2 16 13 0 13 15 9 0 0 13 0 9 7 0 1 0 9 1 0 9 2
15 13 3 7 9 1 0 9 2 0 15 13 1 9 9 2
16 15 0 1 15 13 2 7 3 13 15 0 9 1 0 9 2
2 0 9
4 0 9 11 11
28 12 0 0 9 0 9 15 1 9 0 9 13 0 9 11 11 7 1 10 9 13 12 9 1 0 9 9 2
48 15 0 2 9 12 9 2 15 13 1 0 9 7 1 9 12 3 1 0 0 9 2 3 3 11 13 10 0 9 9 0 9 2 0 1 0 9 12 0 0 9 1 10 0 9 1 11 2
26 11 1 9 13 1 0 9 9 2 3 0 1 0 0 9 2 3 7 10 9 13 13 3 0 9 2
57 0 0 2 3 3 3 0 9 11 13 1 0 11 15 9 7 9 2 3 15 15 1 9 13 10 2 0 2 2 0 9 2 1 15 13 16 9 1 9 3 0 2 7 1 0 9 1 0 9 1 9 7 9 13 3 9 2
9 3 7 15 13 3 3 2 2 2
34 9 13 1 0 9 13 0 2 3 0 9 0 0 9 2 15 13 1 9 7 1 0 9 13 1 15 0 0 2 9 0 9 2 2
9 14 15 13 3 9 1 0 9 2
24 0 0 9 13 0 9 1 9 2 7 13 1 9 0 16 0 2 0 3 1 9 7 9 2
3 11 13 11
2 11 2
23 0 9 0 9 0 9 11 13 0 9 11 11 2 12 2 2 0 2 9 2 9 12 2
43 7 16 11 13 1 9 1 0 9 2 3 15 13 12 2 9 11 1 11 1 0 9 2 13 1 10 0 11 1 0 9 1 0 11 1 11 7 0 11 11 1 11 2
17 15 15 1 0 9 13 1 0 9 1 9 12 9 3 1 11 2
2 0 9
4 12 2 12 2
5 11 12 2 12 2
3 11 12 2
4 9 1 12 9
2 11 2
34 9 11 11 2 0 9 9 9 12 7 0 9 0 9 0 9 11 4 13 1 11 1 9 1 12 9 2 15 13 1 9 12 9 2
14 9 13 0 9 1 3 9 9 2 16 15 3 13 2
12 9 9 1 0 9 13 10 9 1 12 9 2
10 9 13 13 9 2 16 4 9 13 13
5 11 2 11 2 2
45 16 4 13 13 9 0 9 9 11 0 0 2 0 9 9 12 9 2 2 0 9 9 2 13 3 9 1 9 7 9 9 11 11 1 9 11 11 7 1 0 9 13 13 9 2
20 2 9 15 3 13 1 9 2 1 9 9 13 9 3 2 2 13 9 11 2
9 2 15 15 3 13 2 13 9 2
27 1 12 12 9 15 3 13 3 12 0 9 2 11 2 11 7 11 2 7 1 9 1 15 13 0 2 2
21 9 13 1 11 13 2 16 1 11 13 0 9 2 3 4 13 13 2 16 13 2
7 15 13 7 9 0 9 2
27 2 9 4 13 1 0 9 2 7 7 4 13 13 9 1 12 9 1 9 2 15 13 1 11 0 9 2
15 7 10 9 7 13 1 9 9 0 9 2 2 13 11 2
12 0 2 9 2 13 1 0 9 12 0 9 2
16 13 15 7 1 9 2 7 4 13 1 11 13 9 1 9 2
10 1 15 15 1 9 13 9 13 9 2
33 9 3 13 9 2 16 9 15 9 13 2 16 4 15 0 9 3 13 1 15 2 16 1 11 1 0 9 13 1 9 2 2 2
13 0 9 11 0 0 13 3 0 9 1 12 9 2
5 9 1 0 2 11
3 0 11 2
19 0 0 0 9 0 9 0 13 1 9 1 0 11 2 0 9 10 9 2
17 0 9 13 11 0 9 2 9 0 11 2 0 9 7 1 11 2
31 13 13 0 9 1 0 9 2 15 15 1 0 11 13 1 0 9 2 7 15 4 9 13 1 0 9 1 9 12 9 2
20 1 0 9 13 13 1 9 2 9 2 0 9 11 2 0 0 0 9 11 2
12 9 9 13 12 2 0 12 7 0 12 9 2
3 9 1 9
3 0 11 2
16 0 9 11 2 0 1 9 1 9 9 11 2 15 13 9 2
18 9 15 13 2 16 12 2 9 13 11 12 9 2 16 15 13 13 2
12 0 9 4 11 13 1 9 1 9 9 11 2
8 9 3 13 11 3 1 9 2
26 0 9 9 13 9 2 1 15 0 9 0 9 1 9 13 2 16 11 1 9 9 13 9 0 9 2
6 15 15 13 1 9 0
5 15 15 1 15 13
6 15 15 13 1 9 0
12 0 12 2 9 11 13 13 0 9 0 9 2
20 13 7 9 2 16 15 10 0 9 3 3 13 1 0 9 14 3 1 9 2
18 9 9 1 9 13 13 14 0 9 2 7 3 9 0 9 0 9 2
8 14 11 13 1 0 9 12 2
6 13 7 11 16 11 2
18 15 0 2 15 15 1 9 9 13 0 2 0 2 11 2 13 0 2
8 7 3 0 11 3 3 13 2
11 13 7 14 1 9 7 9 1 9 9 2
13 3 15 13 2 16 3 0 13 7 9 1 9 2
38 7 3 16 11 13 1 0 9 3 3 2 16 13 14 12 0 9 7 13 1 0 9 13 9 2 9 11 13 12 9 7 0 1 9 11 3 12 2
19 3 0 9 2 15 3 2 16 15 13 1 0 9 2 13 7 11 11 2
19 15 3 3 13 1 9 7 1 12 3 0 0 9 11 9 12 1 9 2
17 9 11 13 16 9 1 0 9 9 9 2 0 9 9 9 9 2
13 7 7 0 7 0 9 7 0 9 3 13 15 2
10 0 13 3 9 2 3 1 0 9 2
42 3 9 9 11 11 11 11 14 13 9 1 9 2 3 13 9 3 9 11 2 10 9 1 0 9 10 9 13 7 15 14 7 10 15 3 13 2 15 13 0 9 2
10 15 13 2 16 15 13 3 1 9 2
15 3 1 9 3 13 3 3 2 9 9 12 13 3 3 2
23 12 0 7 3 14 3 0 0 9 2 11 7 11 2 3 3 13 10 9 12 14 3 2
9 13 11 11 1 0 9 1 11 2
2 11 2
22 0 0 9 1 0 11 15 13 9 2 16 0 9 11 2 12 2 13 13 1 11 2
29 3 1 0 9 1 0 2 11 11 3 13 0 9 1 0 9 7 1 9 9 9 7 9 13 1 0 0 9 2
21 9 0 9 1 9 13 2 16 15 1 15 13 2 16 4 11 13 1 11 9 2
42 3 1 9 11 11 2 9 0 0 9 1 9 2 3 15 1 11 1 9 13 2 7 16 11 13 2 2 16 13 10 9 1 9 2 4 15 3 13 1 9 2 2
21 9 0 9 11 11 13 2 2 9 1 9 13 2 16 4 15 3 13 1 9 2
17 16 13 11 13 1 11 2 13 3 13 0 9 2 3 3 2 2
19 1 9 0 9 13 0 0 9 2 15 15 13 1 10 9 2 9 11 2
7 13 1 0 9 1 9 2
1 9
12 11 2 9 9 2 11 2 11 2 11 2 2
18 11 2 9 2 9 9 2 11 2 11 2 2 2 11 2 11 2 2
4 9 1 11 13
6 11 11 3 13 0 9
2 11 2
18 11 11 2 12 2 2 9 0 11 15 13 3 1 10 0 0 9 2
15 12 15 13 1 11 2 12 1 11 7 12 1 0 11 2
11 1 0 0 9 13 1 9 0 12 9 2
13 3 1 10 0 0 9 13 9 1 0 0 9 2
31 2 13 13 0 16 0 9 7 3 15 13 2 16 13 1 9 2 15 13 1 10 9 0 7 15 13 3 1 0 9 2
28 16 15 13 9 2 0 9 4 15 13 1 11 2 3 4 13 9 13 0 9 2 15 13 15 16 3 15 2
20 13 2 3 3 11 2 1 11 7 1 11 13 3 9 2 15 13 9 2 2
10 9 1 11 1 0 9 1 11 13 2
6 2 15 1 10 9 2
19 13 4 3 7 10 0 9 2 7 11 15 13 1 9 2 3 13 13 2
13 1 11 13 9 11 2 11 1 15 3 13 9 2
22 3 15 15 13 0 9 11 9 11 1 9 11 2 16 4 13 9 13 15 1 11 2
20 13 4 2 16 9 15 13 1 0 9 9 9 2 7 3 4 15 3 13 2
14 10 9 13 7 9 2 16 0 9 13 13 1 9 2
19 3 13 11 15 13 1 15 2 16 15 1 9 13 13 15 1 0 9 2
18 3 13 2 16 4 13 3 3 1 0 9 2 3 1 9 9 2 2
12 10 13 9 1 0 9 9 1 0 9 11 2
8 2 15 9 13 0 9 3 2
11 13 15 2 16 0 0 9 9 3 13 2
14 3 1 0 9 4 13 2 3 9 13 1 0 9 2
20 11 3 15 13 1 15 2 10 0 9 15 13 7 1 15 7 15 13 3 2
9 13 3 1 10 9 3 0 9 2
17 7 0 4 2 16 4 15 15 13 2 16 9 11 13 15 3 2
13 13 3 0 0 9 2 15 13 1 9 9 2 2
15 1 11 4 13 7 0 9 1 0 9 1 11 3 15 2
22 2 13 9 2 16 9 11 15 1 15 13 2 16 4 13 0 13 9 1 9 11 2
23 13 4 10 9 1 9 7 12 2 9 1 9 1 11 4 13 2 16 15 1 15 13 2
12 3 4 15 13 2 13 15 14 9 1 9 2
10 7 3 3 15 11 13 1 9 11 2
21 0 2 15 15 3 13 2 13 2 16 11 15 3 13 2 7 3 15 13 3 2
21 3 15 15 13 9 9 9 11 7 9 4 13 2 3 4 15 1 10 9 13 2
18 9 4 13 2 13 4 15 3 2 16 15 3 13 0 0 9 2 2
11 13 10 9 10 9 1 9 11 2 11 2
6 2 13 4 15 15 2
21 15 15 3 13 2 16 15 13 10 9 7 16 15 10 0 9 13 1 0 9 2
11 16 1 15 13 15 2 3 13 13 2 2
9 1 3 3 15 3 13 16 9 2
7 2 3 4 13 3 3 2
17 16 15 13 10 9 7 13 15 9 2 4 15 13 13 3 3 2
9 7 3 15 3 4 13 0 9 2
12 7 3 2 16 13 2 3 13 9 0 9 2
17 12 9 1 15 9 13 2 7 1 10 9 15 13 13 13 2 2
12 13 2 16 4 13 13 7 3 16 1 11 2
14 2 7 16 9 11 4 13 3 2 0 9 3 13 2
23 16 15 9 11 4 13 2 3 1 11 13 3 16 10 12 9 2 1 10 13 9 2 2
5 9 0 7 0 9
10 1 9 15 3 13 2 16 11 13 11
4 11 2 11 2
31 9 9 11 2 11 11 1 9 1 11 3 13 9 0 9 0 0 9 11 11 1 0 9 1 0 9 0 7 0 9 2
17 9 15 13 10 9 1 9 1 9 1 0 0 9 1 0 11 2
11 2 3 13 0 2 1 3 0 9 13 2
20 1 0 9 13 13 7 1 9 2 16 11 13 0 1 0 15 0 9 13 2
16 13 2 14 15 0 9 0 2 4 13 1 9 13 11 11 2
11 0 9 13 1 9 3 2 2 13 11 2
26 3 1 9 15 1 9 9 13 9 11 2 11 11 7 11 11 2 1 9 3 13 9 3 11 11 2
27 9 9 11 7 11 15 13 13 1 0 9 3 2 3 1 9 1 11 7 11 13 11 11 1 11 11 2
9 10 9 13 11 11 1 11 11 2
41 9 9 11 2 11 7 11 13 1 9 1 0 9 1 0 9 1 9 9 2 9 9 1 9 7 9 13 0 9 1 12 2 9 2 0 9 13 1 12 9 2
14 1 9 1 9 1 0 9 15 13 1 11 3 11 2
24 10 0 9 11 11 15 3 13 13 9 0 0 9 2 1 15 13 1 0 12 9 0 9 2
9 7 4 1 9 1 0 11 13 2
26 9 0 9 11 11 13 2 16 9 1 11 13 11 11 2 15 4 13 3 1 11 11 13 1 9 2
11 1 9 11 13 1 11 11 7 11 11 2
3 9 0 9
2 11 2
31 0 9 1 9 0 9 13 1 12 2 9 9 1 0 9 1 11 9 11 1 9 11 2 11 2 9 2 11 2 11 2
11 9 9 15 1 10 9 13 11 1 11 2
10 1 9 1 9 1 9 13 11 0 2
3 9 3 0
14 9 11 11 13 2 15 15 13 1 0 9 2 2 2
5 11 2 11 2 2
40 9 2 15 13 0 9 11 11 2 9 1 9 2 0 2 2 7 15 13 9 9 11 11 0 9 1 0 0 9 3 0 1 9 11 2 3 3 13 9 2
23 9 11 11 11 9 11 3 13 2 15 0 9 13 2 16 9 13 9 2 15 13 9 2
41 2 14 2 9 11 15 1 10 9 13 3 3 3 2 1 9 15 3 1 0 9 13 2 16 9 10 9 13 2 2 13 11 11 2 9 0 9 11 11 11 2
19 2 9 10 9 1 9 11 13 0 9 2 16 13 13 0 9 1 9 2
24 3 7 13 2 16 15 4 13 13 1 0 9 2 7 16 9 0 9 15 3 14 13 2 2
2 11 9
3 11 11 2
18 11 11 1 0 9 15 13 9 9 1 9 1 9 1 0 11 11 2
16 12 0 9 1 9 9 13 0 11 2 0 11 7 0 11 2
18 1 0 9 15 9 11 13 1 9 9 2 15 13 1 11 7 11 2
2 13 3
14 0 9 13 1 0 9 2 7 1 9 9 13 13 3
8 11 2 1 10 0 9 2 2
19 0 9 1 0 9 9 13 0 0 9 1 9 9 16 9 9 10 9 2
19 13 15 15 12 0 7 12 0 9 2 15 15 13 1 0 9 1 9 2
40 1 9 2 15 15 13 3 9 9 1 10 9 2 3 0 16 13 0 9 2 7 15 13 9 1 9 0 9 1 10 0 9 2 13 15 9 0 0 9 2
7 0 9 13 3 13 3 2
24 10 9 13 13 3 2 9 15 13 1 0 9 2 7 0 9 9 15 13 13 0 0 9 2
26 9 11 11 13 1 0 9 12 9 1 9 7 0 9 1 9 11 11 13 1 9 9 9 0 9 2
14 10 9 4 13 7 9 9 9 2 3 0 1 9 2
21 13 15 13 1 9 7 9 2 16 0 9 9 11 1 0 9 1 9 9 13 2
15 10 9 2 0 3 1 0 9 2 13 1 0 0 9 2
16 10 0 9 2 16 0 3 1 9 2 3 3 1 9 13 2
18 9 0 9 13 0 2 13 15 14 9 9 2 0 3 1 0 9 2
33 9 10 9 15 1 9 11 13 2 16 10 9 9 2 0 2 0 2 7 1 9 3 0 2 13 1 0 9 9 13 1 0 2
19 10 10 0 9 1 9 13 3 15 15 2 3 10 9 9 9 1 9 2
28 13 2 16 1 0 9 9 1 0 9 13 9 2 12 0 9 2 7 1 0 9 13 12 9 2 12 2 2
16 3 3 13 9 11 0 9 0 9 11 7 11 1 9 9 2
13 1 15 13 9 7 3 13 7 1 0 9 9 2
26 11 11 3 13 14 16 9 2 7 7 16 9 0 9 10 0 9 2 12 0 11 7 12 0 11 2
26 9 0 2 11 7 11 2 16 1 0 9 9 0 2 15 3 0 2 15 0 2 13 3 1 9 2
33 10 0 9 13 9 0 9 7 13 3 0 2 16 1 10 0 9 1 9 7 1 9 15 13 3 3 9 2 15 3 13 11 2
20 1 9 13 1 9 9 2 0 9 12 15 13 2 7 12 1 15 13 9 2
16 0 9 11 13 0 2 0 9 11 0 2 0 9 11 0 2
14 0 0 9 13 14 0 9 1 9 2 15 15 13 2
15 1 9 9 12 1 0 11 9 3 13 14 0 9 11 2
5 9 9 1 9 2
7 14 12 9 13 0 9 2
4 11 3 1 0
4 11 1 11 2
22 11 11 15 13 9 12 2 9 0 9 11 1 11 2 7 13 3 0 9 0 9 2
10 1 0 11 13 9 12 2 12 9 2
33 0 9 11 13 9 1 12 9 7 9 0 0 9 11 15 13 1 9 12 2 12 9 2 1 12 1 10 0 9 11 1 11 2
2 9 2
6 11 2 11 2 2 12
6 11 2 11 2 2 12
6 11 2 11 2 2 12
2 0 9
2 11 2
18 11 11 2 0 0 9 13 0 9 1 9 0 9 1 0 0 9 2
40 11 13 1 9 0 9 11 2 11 2 12 2 12 2 12 9 2 15 15 3 13 11 1 11 1 9 12 1 9 9 9 11 2 11 2 12 2 12 2 2
5 9 2 11 2 11
3 11 11 12
88 12 1 9 1 0 11 2 12 11 2 12 2 9 2 12 0 9 2 12 11 11 2 12 0 2 12 0 9 12 2 0 2 9 2 12 11 7 10 9 2 12 11 2 12 3 2 16 13 9 2 12 9 2 12 11 2 12 15 2 12 2 9 0 2 9 2 12 0 9 2 0 2 9 2 12 9 7 0 9 1 9 2 0 2 0 2 9 2
2 11 12
29 12 0 9 2 9 2 12 13 9 2 12 15 15 13 2 13 2 12 11 2 12 9 1 9 2 12 9 7 9
2 11 12
93 12 9 2 12 9 7 9 2 12 9 1 9 2 12 9 11 2 12 0 2 12 15 13 0 9 2 12 0 9 2 12 11 2 12 9 9 2 12 11 2 12 9 9 2 12 0 9 2 12 0 9 2 12 12 9 1 9 9 2 12 9 7 9 2 12 3 1 9 2 12 9 11 2 12 0 9 2 12 0 9 2 12 9 1 9 2 12 0 9 2 12 0 9
1 12
118 12 9 2 12 9 1 9 2 12 0 9 2 12 9 1 9 2 12 11 2 12 0 9 2 12 9 2 12 9 1 9 2 12 1 0 9 11 2 12 9 1 11 2 12 9 2 12 9 11 11 2 12 9 2 11 2 12 9 1 11 2 12 0 9 2 12 9 2 12 9 12 2 9 2 12 9 1 11 2 12 10 9 2 12 9 2 12 9 2 12 9 9 2 12 11 11 2 12 0 9 2 12 9 2 12 9 2 12 9 15 0 2 12 0 9 2 12 9
4 0 9 9 13
5 11 2 11 2 2
17 0 9 7 1 9 1 3 12 12 9 13 9 1 11 1 11 2
13 9 0 0 9 15 13 0 9 1 9 1 11 2
11 0 9 13 2 16 9 13 3 1 11 2
14 1 9 1 10 9 15 13 0 9 7 13 0 9 2
8 0 9 0 9 13 13 11 2
4 0 9 1 11
5 11 2 11 2 2
27 1 12 9 1 9 7 1 0 1 9 13 1 9 9 0 12 0 9 1 10 9 1 11 9 1 11 2
5 0 9 9 13 2
10 1 9 13 9 9 2 15 9 13 2
15 0 9 13 2 16 9 9 13 9 9 1 0 0 9 2
11 9 9 13 3 0 2 9 1 9 13 2
4 9 1 9 13
7 11 2 11 2 11 2 2
23 9 9 3 13 1 3 0 0 9 1 0 9 11 1 0 9 1 9 1 9 9 13 2
24 0 0 9 13 1 12 9 9 1 0 9 14 1 11 1 9 1 9 12 9 1 0 9 2
13 11 13 1 0 9 3 1 0 9 0 12 9 2
14 9 9 15 0 9 0 9 13 1 12 7 12 3 2
10 1 9 3 13 9 9 1 0 9 2
10 1 0 9 4 13 9 0 9 9 2
15 1 9 9 0 9 13 0 9 1 12 2 9 9 9 2
27 0 9 2 15 4 11 1 12 9 1 0 9 13 2 4 3 13 1 0 9 16 1 3 0 0 9 2
15 3 4 13 7 9 9 2 15 1 15 13 3 1 11 2
13 1 9 0 9 15 13 1 0 9 11 0 9 2
18 15 12 9 11 1 9 12 7 12 9 15 13 9 1 0 9 11 2
23 1 9 9 1 10 9 1 12 9 7 3 0 0 9 4 1 12 9 13 0 9 13 2
15 1 0 0 9 2 3 11 3 13 9 2 13 9 0 2
8 10 9 4 13 3 1 9 2
8 9 0 9 2 9 13 0 9
1 9
2 11 12
3 12 9 12
8 12 9 9 2 9 11 2 11
3 12 9 9
8 12 9 1 9 2 12 2 2
5 12 13 9 1 9
7 12 16 13 9 2 0 9
3 12 9 9
9 12 0 9 1 9 2 12 2 2
4 12 9 1 9
3 12 0 9
2 12 9
3 12 1 12
2 12 9
6 12 9 9 2 12 11
3 12 0 9
2 12 9
6 12 9 2 12 2 2
12 12 0 9 1 9 9 2 12 2 2 0 9
2 12 9
6 12 0 2 0 2 11
4 12 9 1 9
7 12 1 9 2 12 2 2
2 12 9
6 12 9 2 9 2 9
6 12 0 9 2 0 9
5 12 11 2 9 11
6 12 9 2 9 2 9
2 12 11
14 12 9 9 2 9 9 2 0 9 1 9 12 2 9
2 12 9
12 12 11 2 11 2 11 2 9 2 12 2 2
6 12 0 2 0 2 11
2 11 12
4 12 9 2 9
2 12 9
2 12 11
3 12 9 9
3 12 9 12
3 12 0 9
3 12 11 9
2 12 9
7 12 9 9 1 0 2 9
3 12 9 11
3 12 9 9
2 12 0
4 12 9 1 9
4 12 9 1 9
2 12 11
3 12 9 12
2 12 9
3 12 0 9
2 12 9
4 12 11 0 9
10 12 13 0 9 2 2 1 3 0 9
10 12 16 9 1 9 2 9 1 11 11
13 12 0 9 2 1 9 9 2 11 2 11 2 11
3 12 9 9
4 12 9 7 9
4 12 9 11 11
2 11 12
3 12 0 9
4 12 0 11 9
3 12 11 9
2 12 9
4 12 0 11 9
3 12 0 11
4 12 0 11 9
3 12 0 11
3 12 9 9
3 12 0 11
3 12 9 9
3 12 0 11
3 12 9 11
3 12 11 11
3 12 11 12
3 12 9 3
3 12 9 11
3 12 9 3
3 12 11 11
2 12 9
3 12 0 9
6 12 9 2 12 2 2
2 12 9
7 12 9 11 2 0 2 9
6 12 0 9 2 9 11
8 12 9 2 0 2 9 1 9
4 12 11 2 12
3 12 0 9
2 12 9
3 12 9 3
2 9 9
42 12 0 9 2 12 0 9 2 0 9 2 12 9 9 2 9 2 12 0 9 11 2 9 2 12 0 9 2 9 11 2 12 9 1 9 2 12 9 3 2 0 9
2 9 9
53 12 9 0 9 1 9 2 12 9 2 12 0 9 2 12 11 2 9 2 12 11 2 0 9 2 12 9 2 12 0 9 2 12 11 2 11 2 9 2 12 9 9 2 9 2 12 9 2 12 9 9 2 9
5 9 9 1 0 9
5 11 2 11 2 2
23 9 3 1 12 12 9 13 9 2 15 13 0 9 7 0 9 1 0 9 9 1 11 2
19 9 9 15 13 2 9 3 13 2 16 3 1 9 15 1 0 9 13 2
5 1 9 9 13 2
4 13 7 13 9
7 11 1 11 2 11 2 2
16 0 9 1 9 12 9 13 1 9 1 11 1 11 12 9 2
17 13 1 9 1 9 7 16 12 13 9 9 2 0 15 3 13 2
19 1 9 9 1 9 15 9 1 10 9 13 12 9 2 12 9 7 9 2
8 9 13 0 9 1 0 9 2
4 9 0 1 9
5 11 2 11 2 2
14 0 9 13 1 0 9 1 9 11 1 11 0 9 2
17 13 1 9 2 9 13 1 9 2 13 1 15 7 13 15 13 2
9 0 15 3 13 9 13 7 13 2
4 13 9 0 9
5 11 2 11 2 2
19 0 9 1 0 9 1 0 9 1 9 11 13 12 0 0 9 0 9 2
16 1 9 2 16 9 0 9 15 13 9 2 9 1 9 13 2
21 1 11 1 9 13 1 9 2 13 1 11 7 3 15 9 13 1 12 9 9 2
13 1 10 9 13 0 9 13 7 1 10 9 13 2
6 1 0 9 13 13 9
2 11 2
22 0 9 13 0 9 1 9 9 9 0 9 11 11 13 1 9 10 9 0 0 9 2
23 13 3 1 9 0 9 1 9 0 9 2 1 15 4 9 1 9 3 9 9 13 13 2
31 9 9 13 0 0 9 2 14 1 0 0 9 2 15 4 1 12 9 13 0 9 2 4 13 0 9 1 9 7 9 2
19 1 15 13 13 3 12 9 0 9 7 1 9 9 9 2 9 7 9 2
26 3 15 13 9 11 11 11 2 9 9 15 13 2 16 9 2 15 13 2 4 13 14 1 0 9 2
23 1 15 1 12 9 13 1 9 1 10 9 0 0 9 7 1 0 9 9 13 9 9 2
27 9 0 9 2 15 10 9 13 1 9 2 13 13 9 1 0 9 2 7 3 13 1 0 11 0 9 2
10 1 9 4 13 13 9 3 12 9 2
36 9 1 0 9 2 15 13 13 13 1 9 12 2 13 12 9 9 7 1 10 9 4 3 14 12 9 13 2 16 4 13 0 9 7 9 2
22 1 9 9 13 10 9 11 11 2 2 13 4 13 9 9 2 15 15 13 15 13 2
14 13 15 13 15 9 1 12 0 9 7 12 0 9 2
8 0 9 13 1 9 3 12 2
12 0 0 9 15 13 13 1 0 9 0 2 2
18 0 7 3 12 1 0 9 9 9 13 14 0 0 9 1 0 9 2
12 9 1 9 0 0 0 9 3 9 9 13 2
4 9 9 13 9
23 11 11 13 2 16 10 9 13 9 0 9 0 1 9 1 0 9 1 11 1 11 11 2
10 9 15 13 1 9 1 9 0 9 2
9 9 4 13 12 9 1 10 9 2
6 0 9 0 9 13 2
27 3 13 9 11 2 16 4 1 9 9 13 1 9 11 0 9 2 3 1 9 9 9 13 4 9 13 2
13 9 2 1 9 2 7 4 13 14 12 2 9 2
26 10 9 15 9 1 0 9 11 13 1 9 11 11 2 9 9 11 2 9 0 9 11 7 0 9 2
19 11 11 13 2 16 1 0 9 13 15 9 1 9 1 0 9 1 9 2
11 9 4 3 13 0 9 9 11 11 11 2
19 0 9 13 0 9 2 15 13 2 16 13 0 7 0 2 7 0 9 2
15 1 9 11 11 1 12 2 9 1 9 1 9 15 13 2
20 15 15 7 13 1 12 2 9 2 3 13 9 1 0 9 2 11 11 13 2
28 11 11 2 0 9 9 0 9 2 15 13 2 16 15 3 15 14 1 9 0 9 1 0 9 1 9 13 2
17 1 9 9 13 13 10 9 2 7 7 9 1 0 9 13 13 2
6 3 15 13 0 9 2
9 1 9 3 3 9 13 0 9 2
21 1 9 0 9 15 1 9 11 13 0 9 11 11 1 9 9 7 9 0 9 2
9 9 13 9 9 7 13 9 9 2
18 1 0 9 4 15 3 13 7 14 1 12 9 13 1 9 0 9 2
3 9 13 2
7 1 9 13 4 13 0 9
2 11 2
15 9 0 9 3 13 0 13 15 13 1 0 9 0 9 2
10 13 15 9 0 9 9 9 11 11 2
17 9 1 0 9 1 0 0 9 13 9 1 9 9 0 10 9 2
15 16 9 0 9 13 10 9 2 4 15 3 10 9 13 2
11 9 1 10 9 13 9 0 2 0 9 2
13 0 0 9 3 13 1 9 2 1 15 4 13 2
23 3 3 9 7 9 13 1 9 1 9 2 16 4 13 1 0 9 13 0 9 0 9 2
8 12 1 9 1 9 0 9 13
7 11 2 11 2 11 2 2
12 1 10 9 9 0 9 13 9 2 11 11 2
18 0 9 9 9 9 3 13 2 16 11 11 13 9 1 9 11 11 2
11 9 11 13 9 13 1 9 3 10 9 2
30 11 11 2 0 1 0 9 0 9 1 11 2 13 12 1 12 9 2 1 10 9 1 9 13 0 9 9 9 9 2
12 11 11 15 1 0 9 13 1 0 0 9 2
10 13 7 3 13 1 9 2 3 13 2
9 9 10 9 13 9 9 9 9 2
10 1 0 9 11 11 13 10 9 0 2
11 9 7 10 9 15 4 13 2 13 11 2
28 0 9 3 13 13 2 16 0 9 13 9 0 9 0 9 2 15 13 9 1 0 9 1 9 12 7 12 2
6 9 9 13 9 1 9
2 11 2
17 9 9 3 1 9 13 1 9 9 9 1 0 9 11 11 0 2
20 13 12 0 9 0 9 3 1 9 2 7 0 13 7 9 0 1 9 12 2
26 2 1 10 9 13 9 2 16 4 1 15 13 1 9 0 2 16 13 12 9 3 2 2 13 11 2
23 9 15 1 11 13 1 9 9 2 1 9 9 2 2 1 15 4 13 4 9 13 3 2
15 1 9 9 1 12 2 9 4 9 13 4 13 1 9 2
11 0 9 4 13 13 1 0 9 12 9 2
8 9 13 13 9 1 9 0 9
2 11 2
17 1 9 0 9 1 0 11 13 1 9 0 9 9 13 9 9 2
11 13 15 9 9 1 9 0 9 11 11 2
17 1 15 15 1 15 4 13 3 0 9 13 3 1 10 9 9 2
7 9 13 0 9 0 9 2
18 9 0 9 2 14 12 0 9 2 13 7 3 2 3 1 0 9 2
31 3 3 13 11 2 9 15 13 14 3 2 16 0 9 13 9 0 0 9 7 1 9 1 0 0 9 13 0 9 9 2
24 15 13 1 9 0 9 2 1 9 0 9 2 1 0 9 1 9 13 0 9 1 9 11 2
30 9 4 3 13 14 1 9 2 3 14 1 9 1 9 9 0 9 2 2 3 1 10 9 13 3 0 9 10 9 2
7 3 13 1 11 0 9 2
11 1 0 10 9 13 0 9 12 12 9 2
13 11 2 11 3 3 13 9 1 9 1 0 9 2
18 13 3 1 9 0 9 2 3 9 2 10 9 4 13 1 0 9 2
9 1 0 9 1 11 13 0 9 9
5 11 2 11 2 2
32 1 0 9 9 0 0 2 0 9 13 9 11 11 11 9 9 14 1 9 0 9 7 9 2 7 3 1 9 0 9 9 2
21 2 1 12 9 13 0 9 1 0 9 1 0 9 13 2 2 13 3 1 11 2
15 1 0 9 4 1 15 13 4 13 0 9 0 0 9 2
21 9 11 11 2 11 2 13 9 0 7 0 9 1 0 0 7 0 9 1 0 2
17 3 13 9 1 9 13 0 9 1 9 0 9 1 9 10 9 2
5 9 4 3 13 9
7 11 2 11 2 11 2 2
17 15 9 2 15 1 9 13 3 9 2 13 0 3 0 9 13 2
8 13 15 15 0 9 11 11 2
22 9 13 0 9 13 2 16 3 9 13 1 9 0 9 0 9 9 7 1 0 9 2
23 10 0 9 13 9 9 11 11 2 15 13 1 9 12 9 11 7 12 11 2 1 9 2
11 11 3 12 1 9 3 13 1 10 9 2
12 11 1 15 13 2 16 1 10 9 4 13 2
27 2 3 7 13 2 16 1 10 9 15 9 9 9 7 9 13 2 9 15 7 13 2 2 13 0 9 2
17 11 11 2 15 13 3 0 0 9 2 0 9 1 9 3 13 2
14 2 1 9 9 4 13 10 0 9 2 2 13 11 2
13 13 2 16 13 13 9 1 15 12 0 9 13 2
13 2 3 4 7 1 9 13 0 9 2 2 13 2
35 7 1 0 0 9 0 9 15 0 9 1 9 7 9 1 0 9 13 3 1 9 2 15 4 13 9 0 9 7 0 9 9 0 9 2
26 0 9 11 11 11 2 11 2 13 1 0 9 1 10 9 2 0 1 9 1 9 9 9 0 9 2
19 9 2 15 13 2 4 13 1 0 2 0 9 2 15 13 1 0 9 2
21 0 9 15 13 1 9 11 11 2 9 1 9 2 0 9 2 9 7 12 9 2
11 1 11 4 9 13 16 9 1 0 9 2
21 1 0 2 0 9 4 9 13 3 1 9 2 1 15 4 9 13 1 9 11 2
6 9 1 9 13 9 9
23 9 4 1 10 9 1 0 9 13 3 1 9 0 9 2 9 0 9 7 9 9 9 2
13 11 15 13 2 16 4 9 9 13 13 15 0 2
29 2 7 13 9 1 9 7 9 2 15 15 13 2 13 2 7 14 7 3 3 15 3 13 15 13 2 2 13 2
15 9 13 1 9 0 9 9 13 1 9 2 7 13 9 2
31 9 9 15 13 2 16 10 9 13 4 13 7 1 0 9 1 9 3 0 9 1 12 2 9 2 1 1 10 0 9 2
14 9 0 9 11 3 13 0 9 9 1 14 9 9 2
5 2 13 10 9 2
15 15 13 0 3 13 7 13 2 2 13 9 11 11 11 2
19 9 13 1 15 1 9 9 1 9 0 9 0 2 16 13 10 0 9 2
25 1 0 13 2 16 4 0 9 13 13 14 1 9 9 9 2 3 1 9 12 2 3 13 9 2
7 2 9 13 4 13 3 2
10 15 7 10 9 13 2 2 13 11 2
16 9 13 10 3 0 0 9 4 13 3 13 0 7 0 9 2
31 2 0 9 1 9 9 10 0 9 7 9 0 9 1 9 1 0 0 9 13 1 9 9 2 2 13 9 9 11 11 2
23 9 9 11 11 15 13 2 16 4 15 3 13 3 13 9 9 2 0 1 9 0 9 2
17 2 9 3 13 2 16 4 1 0 0 9 13 4 9 3 13 2
27 13 3 13 9 9 1 9 1 9 2 7 13 2 16 15 3 13 10 9 10 0 9 2 2 13 11 2
6 9 1 9 1 0 9
13 2 11 11 13 14 9 7 9 2 7 3 9 2
14 10 9 3 13 14 9 7 9 2 7 3 9 2 2
27 10 9 13 1 10 9 1 9 11 11 9 0 0 9 2 10 3 3 0 9 13 1 0 9 1 11 2
31 10 9 13 14 9 1 9 2 15 7 1 9 13 14 1 11 2 7 3 9 9 0 9 2 3 0 0 9 0 11 2
31 0 7 0 0 9 13 9 2 16 3 0 9 9 0 9 2 15 13 11 11 2 1 15 13 7 0 0 7 0 9 2
44 15 9 13 1 0 9 0 0 9 0 9 1 12 2 9 2 3 16 12 1 9 3 3 0 9 12 13 9 9 0 9 2 14 1 0 9 0 9 1 9 1 9 0 2
27 0 9 13 0 9 9 1 0 9 1 9 12 2 1 15 13 9 1 9 0 2 0 0 0 9 9 2
43 1 0 11 13 2 16 13 3 0 9 9 0 9 1 15 2 15 13 0 9 1 9 1 9 2 12 7 3 3 0 9 9 1 9 2 12 2 7 9 2 12 2 2
28 1 0 9 0 9 7 1 9 0 13 0 0 9 1 0 9 2 15 3 1 0 9 0 9 13 10 9 2
20 3 0 9 13 0 9 1 0 9 0 9 2 1 10 9 1 9 0 9 2
23 2 1 9 15 2 15 13 9 2 15 15 3 13 1 0 9 2 2 13 9 1 9 2
33 9 11 11 13 14 9 12 0 9 0 9 2 7 3 0 9 1 9 13 1 9 2 1 15 13 9 13 7 1 15 3 13 2
2 9 9
17 11 15 13 0 9 0 7 0 9 2 3 15 1 0 9 13 2
29 7 9 13 2 9 7 9 13 2 0 7 0 9 7 0 7 0 9 13 14 0 9 7 9 13 3 2 2 2
12 13 9 10 9 1 3 0 9 13 7 9 2
15 13 1 0 0 9 11 2 7 1 0 9 15 9 13 2
22 7 3 13 0 9 13 9 0 9 0 9 2 0 9 9 11 1 9 12 2 9 2
23 13 15 1 9 0 0 9 2 1 15 13 14 13 2 7 7 13 9 1 0 0 9 2
23 9 13 0 9 9 14 1 0 9 7 10 9 2 7 7 1 0 9 11 1 12 9 2
33 9 13 10 9 1 0 9 0 0 9 15 13 9 0 9 7 1 9 0 10 9 1 9 7 0 0 9 0 2 11 2 11 2
16 9 10 3 16 0 9 13 12 0 9 9 0 9 7 9 2
34 10 0 0 9 4 13 3 0 9 2 7 7 9 1 9 9 15 13 1 15 7 13 15 13 9 9 11 1 0 9 1 0 9 2
30 9 13 1 9 14 0 0 9 7 0 9 2 7 7 0 9 9 2 15 9 9 13 0 9 1 9 7 0 9 2
4 0 9 11 11
17 3 1 0 9 10 9 13 0 9 11 11 2 13 15 9 9 2
5 9 13 10 9 2
30 7 15 15 1 10 9 2 0 12 9 9 2 13 2 3 15 13 1 9 11 11 2 16 15 13 3 1 10 9 2
33 13 15 3 3 16 12 9 9 2 16 13 9 9 2 13 1 0 9 2 0 9 0 9 1 9 0 9 2 11 15 13 2 2
18 15 13 3 2 1 0 9 9 2 9 1 9 0 9 0 0 9 2
11 7 10 9 15 13 13 7 13 0 9 2
13 14 2 13 15 0 9 1 9 9 1 10 9 2
30 10 15 13 9 2 10 9 2 16 15 1 9 9 9 2 10 0 2 13 1 9 9 2 16 15 13 1 9 9 2
17 13 4 1 9 10 0 9 2 1 10 9 2 13 4 10 9 2
2 3 2
12 16 15 13 9 3 3 2 16 4 13 9 2
9 0 9 11 11 15 13 2 13 2
9 11 7 1 10 9 1 9 13 2
23 9 15 13 13 9 1 0 0 9 7 15 13 9 1 9 2 13 15 1 15 16 9 2
18 15 4 7 13 3 3 2 16 15 9 11 10 9 3 7 3 13 2
16 7 13 2 7 16 4 3 13 1 9 1 9 13 1 9 2
11 3 15 3 3 13 13 3 0 0 9 2
12 7 3 15 13 9 7 13 3 1 9 9 2
12 9 11 15 13 9 2 9 2 9 2 9 2
4 3 3 3 2
19 11 2 13 2 13 4 9 2 3 4 15 13 2 7 13 15 3 3 2
5 13 15 2 13 2
19 7 3 4 1 9 13 9 0 2 3 0 9 2 2 11 15 13 2 2
9 13 4 15 1 0 9 0 9 2
16 9 11 13 2 16 13 9 2 0 2 1 9 0 2 0 2
13 9 15 13 15 12 2 9 2 10 9 7 9 2
5 13 15 9 9 2
13 7 15 13 10 0 9 2 15 13 13 0 9 2
19 13 15 2 16 9 13 12 0 9 2 16 3 13 9 2 3 13 9 2
10 16 0 13 9 1 0 11 16 9 2
2 11 11
9 9 12 0 9 13 3 2 9 2
9 10 9 13 3 9 9 7 9 2
7 15 0 13 3 3 3 2
5 14 7 15 0 2
10 2 13 7 1 9 7 13 15 3 2
7 14 3 13 0 9 2 2
5 0 9 0 9 9
12 13 12 7 13 2 16 0 9 13 1 9 2
7 9 9 13 1 10 9 2
19 13 15 7 10 0 9 2 3 3 2 13 9 0 0 9 9 11 11 2
7 3 9 7 3 1 15 2
28 2 13 15 0 9 0 2 15 13 1 9 9 10 9 9 9 3 1 9 7 3 1 0 9 2 15 13 2
9 13 15 7 0 9 0 9 9 2
7 13 9 7 0 9 9 2
22 0 9 13 9 2 16 9 13 9 0 0 9 2 15 9 1 9 9 13 0 9 2
18 0 9 1 9 7 9 13 0 0 9 1 15 7 13 15 1 9 2
25 10 9 13 0 2 13 4 2 16 4 9 2 15 1 15 1 9 13 2 13 0 0 9 2 2
16 9 7 9 3 2 13 15 13 2 13 0 9 13 1 9 2
7 13 3 0 9 1 9 2
12 2 13 15 3 2 16 15 9 0 9 13 2
6 10 9 1 15 13 2
12 1 0 9 13 9 2 15 2 15 15 13 2
7 1 9 13 1 10 9 2
6 1 15 13 9 9 2
13 1 0 15 3 0 9 15 9 13 10 9 13 2
6 9 13 7 9 2 2
4 3 13 9 2
5 2 3 2 3 2
13 9 13 1 9 2 1 9 13 15 1 9 2 2
8 1 9 0 4 13 9 0 2
13 2 3 13 9 0 2 0 2 15 15 13 3 2
8 15 15 13 0 0 2 9 2
14 12 9 15 3 13 2 11 0 9 11 7 0 11 2
16 13 15 7 15 0 2 13 3 9 2 15 10 9 3 13 2
11 15 2 15 13 2 13 3 3 0 2 2
7 13 0 10 9 1 9 2
11 2 13 2 15 3 9 1 0 0 9 2
4 2 3 13 2
4 1 0 9 2
9 13 9 7 9 2 15 3 13 2
13 13 2 14 7 13 1 15 2 3 13 7 13 2
11 13 15 9 3 0 9 16 10 9 2 2
17 13 15 0 9 2 9 2 3 15 13 3 2 16 4 3 13 2
10 2 0 9 7 9 13 14 0 9 2
9 1 9 1 10 9 15 3 13 2
24 0 13 2 16 4 15 13 1 9 7 13 1 15 2 15 4 13 13 9 7 9 10 9 2
15 3 13 9 2 7 3 4 13 1 9 1 0 0 9 2
18 16 15 1 10 9 13 2 4 13 3 9 2 3 15 1 15 13 2
15 3 4 15 13 13 1 9 2 3 4 13 15 15 2 2
33 9 16 0 2 3 11 11 2 9 2 2 11 11 2 0 9 2 9 2 2 3 11 11 2 9 2 2 11 11 2 0 9 2
4 0 9 1 9
4 9 1 9 9
14 12 1 0 9 1 9 9 13 3 1 11 11 11 2
28 11 13 2 9 2 0 9 3 0 0 9 11 11 7 11 11 2 1 0 9 2 15 15 3 3 13 9 2
24 0 9 2 15 3 3 13 7 1 9 9 2 13 10 0 9 0 9 3 7 3 3 3 2
22 12 9 4 13 1 9 2 15 3 13 1 0 9 0 9 2 3 15 0 13 9 2
24 9 1 0 9 1 9 11 13 0 9 9 2 9 2 11 2 9 2 9 9 9 7 9 2
17 0 9 13 1 9 9 3 1 9 2 7 1 3 0 9 9 2
5 0 9 15 13 2
28 13 13 9 1 0 9 2 0 0 9 2 0 9 2 1 15 7 3 1 10 9 3 0 1 15 3 13 2
57 3 0 13 0 9 1 9 2 3 15 1 9 13 0 0 9 0 9 2 15 9 11 11 13 9 13 10 9 16 9 9 1 0 9 2 15 3 7 2 10 9 13 2 7 13 15 1 9 11 11 1 9 12 2 9 2 2
32 9 7 9 2 11 11 2 13 3 3 0 9 9 2 15 15 7 1 0 13 13 1 11 11 7 10 9 1 9 1 9 2
22 9 15 13 11 11 11 2 1 15 4 1 10 9 13 1 9 7 0 9 1 9 2
13 0 9 3 13 9 0 7 0 9 1 9 9 2
14 0 9 4 13 0 9 11 11 7 0 9 11 11 2
24 0 9 2 15 0 9 13 9 7 9 11 11 2 9 7 9 11 11 7 9 11 11 0 2
4 9 1 9 13
5 11 2 11 2 2
17 1 12 12 9 3 13 3 1 9 0 9 1 0 9 0 9 2
11 0 9 2 3 12 9 2 13 0 9 2
12 9 1 15 13 3 7 9 9 1 0 9 2
34 9 3 13 13 14 1 9 2 7 13 1 15 13 7 12 9 3 2 7 13 1 12 9 2 9 1 12 2 0 9 1 0 9 2
34 1 9 9 1 0 9 2 0 2 9 2 2 11 11 13 10 9 7 3 13 0 9 1 10 9 3 1 9 9 2 15 13 9 2
20 3 3 4 13 0 9 0 9 2 7 15 15 13 0 9 0 9 0 9 2
4 13 9 7 9
5 11 2 11 2 2
35 1 12 2 9 2 3 1 0 9 1 9 13 1 9 7 13 15 3 2 13 9 1 12 0 0 9 0 9 12 1 9 9 11 11 2
17 0 9 13 1 15 1 9 9 7 13 15 13 9 0 0 9 2
28 11 11 13 1 0 9 7 13 0 2 12 9 0 9 2 0 0 9 7 1 0 9 9 0 9 9 9 2
4 1 9 13 2
13 3 13 1 15 0 9 2 0 9 7 0 9 2
21 1 9 13 0 9 1 9 9 2 1 0 9 13 7 0 0 9 7 0 9 2
30 9 15 13 13 1 0 0 9 2 1 9 12 2 7 1 12 2 9 0 9 1 11 2 9 2 12 2 12 12 2
9 15 4 15 13 1 0 9 9 2
2 9 9
9 15 4 15 13 1 0 9 9 2
18 1 0 9 9 4 15 13 13 0 9 9 11 1 0 9 1 9 2
5 11 2 11 2 11
13 1 0 9 9 4 15 13 9 10 7 10 9 2
5 11 2 11 2 11
7 16 4 15 9 3 13 2
10 16 4 15 13 0 7 13 3 0 2
10 16 4 15 15 13 1 9 1 15 2
6 16 4 13 0 9 2
5 11 2 11 2 11
8 0 9 9 0 9 2 2 2
5 11 2 11 2 11
42 3 0 7 1 9 15 3 3 13 9 2 4 2 14 13 2 16 10 9 13 1 9 2 15 15 3 13 9 0 2 0 2 0 7 0 16 9 2 9 7 9 2
29 16 16 9 13 1 0 9 2 13 2 16 3 3 10 0 9 1 9 13 7 13 13 0 7 1 9 1 9 2
5 11 2 11 2 11
5 1 9 13 14 9
7 11 2 11 2 11 2 2
25 0 9 11 11 2 2 11 13 3 0 9 2 15 13 0 0 9 1 0 9 1 11 2 9 2
16 1 0 0 9 13 0 9 1 9 7 9 9 4 13 9 2
23 9 1 9 0 9 13 12 9 7 3 9 9 1 0 9 13 3 0 16 1 0 9 2
38 9 0 0 11 1 9 1 15 13 1 9 1 0 9 1 12 9 2 7 16 9 13 1 9 0 2 9 1 9 4 15 13 13 1 9 12 9 2
24 0 0 9 2 0 1 0 0 0 9 1 0 9 1 11 2 3 13 1 12 9 0 9 2
10 10 9 9 1 9 0 9 13 13 2
20 1 9 11 11 2 9 9 11 0 11 2 13 1 15 3 12 0 0 9 2
18 1 0 7 0 9 13 3 2 9 0 9 1 11 7 1 0 9 2
11 0 9 1 11 1 11 10 9 13 9 2
17 1 9 0 9 13 7 9 9 1 9 1 0 0 7 0 9 2
22 9 1 9 9 3 13 9 0 0 9 2 15 4 16 0 1 15 1 10 9 13 2
21 11 13 3 1 12 0 9 3 1 9 1 9 0 9 2 0 9 13 7 11 2
5 0 0 1 12 9
7 11 2 11 2 11 2 2
25 0 9 1 9 9 0 0 13 3 0 0 9 1 9 0 9 7 0 9 9 0 9 1 9 2
8 13 15 3 9 9 11 11 2
9 9 3 13 13 15 3 0 9 2
16 13 15 4 7 1 9 9 1 0 9 7 1 9 0 9 2
14 0 9 13 9 9 1 0 7 0 9 0 1 9 2
16 0 9 1 0 9 9 4 13 13 9 0 1 9 7 9 2
26 9 0 0 4 13 0 7 0 9 1 9 11 1 9 1 12 9 2 1 9 9 0 9 13 0 2
10 0 9 4 9 13 1 12 2 9 2
16 0 9 1 9 9 4 13 13 0 16 12 9 1 9 9 2
21 9 9 4 13 1 9 0 1 9 12 9 9 9 9 2 15 9 13 9 13 2
6 1 9 0 9 1 9
7 11 2 11 2 11 2 2
22 0 9 0 9 1 12 9 13 1 0 9 13 9 9 0 9 7 13 10 0 9 2
8 13 15 3 9 9 11 11 2
11 13 7 2 1 10 9 4 13 9 13 2
36 2 1 10 9 13 3 2 16 4 15 13 1 0 9 7 0 9 2 2 13 9 11 2 15 13 3 9 9 0 9 0 1 11 7 11 2
14 2 13 9 2 3 15 0 9 13 1 9 0 9 2
27 9 9 1 9 4 13 9 9 0 9 1 0 9 10 9 2 16 4 15 10 9 13 2 2 13 11 2
20 0 9 7 0 9 0 9 15 13 3 13 3 2 1 9 0 11 1 11 2
15 10 0 9 13 0 0 9 9 1 0 9 14 12 9 2
7 13 15 9 9 11 11 2
23 2 9 0 9 13 1 15 0 2 2 13 3 11 11 2 9 9 9 11 11 1 11 2
14 9 1 11 3 13 2 13 7 3 0 9 0 9 2
19 2 16 1 9 4 3 13 9 9 2 9 0 9 14 13 2 2 13 2
10 9 0 9 1 11 4 13 13 13 2
14 13 15 9 0 9 0 2 9 2 0 9 11 11 2
8 10 9 3 13 10 9 9 2
25 9 2 15 15 13 13 13 2 13 2 16 9 0 9 1 11 4 3 13 7 1 9 0 9 2
27 15 13 3 13 12 9 7 0 9 13 1 10 9 3 13 9 10 9 1 12 9 2 15 4 13 9 2
19 1 10 0 9 9 9 1 11 1 9 9 11 11 11 11 1 9 13 2
21 2 1 9 9 9 13 9 1 12 9 7 13 2 16 9 3 13 0 9 2 2
17 9 9 1 0 9 1 0 7 0 9 13 7 1 0 9 0 2
11 3 0 9 7 9 9 13 1 0 9 2
10 13 15 7 0 9 1 9 1 11 2
22 2 9 4 13 1 9 2 9 15 13 3 0 9 2 2 13 9 9 11 11 11 2
8 0 9 13 1 9 1 12 9
5 11 13 9 13 9
7 11 2 11 2 11 2 2
20 0 0 9 3 13 9 9 1 0 9 1 9 9 1 9 1 12 9 3 2
20 1 9 15 3 13 9 9 2 15 7 13 10 9 1 9 1 3 0 9 2
30 9 15 15 3 13 3 1 10 0 9 1 9 3 1 0 9 2 9 9 3 1 9 1 12 9 13 2 13 2 2
19 1 0 9 13 0 9 1 0 1 9 0 9 0 0 9 12 9 9 2
20 13 15 1 3 0 0 9 2 1 15 15 13 9 0 1 0 12 2 9 2
23 1 0 9 2 15 13 9 1 9 0 1 0 9 2 13 11 9 0 1 12 9 9 2
18 16 15 10 9 13 13 1 0 9 2 4 3 13 13 9 10 9 2
9 13 15 3 9 9 11 11 11 2
15 1 10 9 13 13 9 0 9 1 0 14 1 12 9 2
29 16 4 0 9 7 9 13 10 9 2 13 4 15 9 0 9 13 1 0 9 9 0 9 1 11 2 13 11 2
7 9 0 9 13 3 14 13
7 11 2 11 2 11 2 2
25 0 0 9 13 2 16 12 7 12 9 0 0 9 7 9 15 13 1 9 1 0 9 10 9 2
12 13 15 15 11 11 2 9 9 0 9 11 2
30 1 3 12 9 0 0 9 15 3 3 13 14 12 9 9 2 15 4 1 9 9 13 2 13 7 15 15 9 13 2
15 0 9 4 13 0 9 0 7 0 0 9 1 10 9 2
24 13 3 3 1 9 0 9 2 9 0 9 13 1 11 3 0 16 12 9 1 10 0 9 2
37 9 1 3 0 9 9 1 9 7 9 0 7 13 0 13 14 1 9 2 3 12 0 9 9 3 13 1 0 9 2 3 16 3 13 0 9 2
8 10 9 13 12 2 9 12 2
29 3 1 10 9 13 3 0 13 0 9 2 10 9 13 3 12 2 9 2 0 9 2 2 9 2 7 9 2 2
40 0 9 1 10 9 13 0 1 0 9 13 3 1 12 2 9 7 9 1 9 12 2 12 7 12 9 2 10 9 13 12 2 9 2 3 1 12 2 9 2
21 1 11 11 13 11 3 14 12 12 9 1 9 0 9 1 9 3 12 9 9 2
6 11 1 11 13 3 9
2 11 2
29 9 11 15 13 3 0 9 1 0 9 9 2 7 16 1 0 9 13 10 9 1 9 1 12 9 1 12 9 2
24 1 11 13 0 9 1 3 0 9 1 11 0 9 11 1 12 9 2 3 12 9 2 2 2
45 13 11 11 1 12 9 2 12 9 2 2 2 9 11 2 11 1 12 9 2 12 9 2 2 2 11 1 12 9 2 12 9 2 2 7 11 1 12 9 2 12 9 2 2 2
17 9 0 9 1 9 13 1 11 3 1 12 9 1 12 9 9 2
4 9 9 13 9
2 11 2
21 9 0 9 1 9 1 9 0 0 9 12 2 9 13 9 1 0 9 0 9 2
11 3 15 7 13 2 16 4 10 9 13 2
8 3 15 9 13 13 0 9 2
12 9 4 13 1 9 0 9 1 9 0 9 2
21 0 9 9 11 11 11 13 2 16 9 1 9 13 2 16 4 15 1 15 13 2
14 2 13 4 9 1 10 9 7 15 4 15 3 13 2
11 3 4 3 13 9 1 9 2 2 13 2
15 9 0 9 13 4 12 2 9 12 13 1 9 0 9 2
18 16 7 9 2 15 15 13 13 2 13 9 2 13 0 9 1 9 2
14 2 1 10 9 15 13 3 15 0 2 2 13 11 2
18 2 3 15 13 2 16 14 15 9 4 13 3 2 3 4 13 13 2
12 10 9 13 0 2 13 15 3 3 0 2 2
27 9 9 13 7 11 11 2 9 0 9 2 15 13 1 9 9 12 9 13 9 0 9 1 0 9 11 2
17 2 16 4 15 13 1 0 9 2 3 4 15 13 2 2 13 2
19 11 7 0 9 0 9 11 11 13 0 9 0 9 1 0 9 1 0 2
13 13 15 7 13 2 15 7 3 13 1 9 13 2
10 2 9 11 3 13 2 2 13 11 2
14 9 13 0 9 0 0 9 2 1 15 0 9 13 2
21 13 1 15 7 9 1 9 9 2 1 9 9 9 2 7 15 7 9 0 9 2
4 0 9 1 11
7 11 2 1 10 9 2 2
7 9 0 9 13 1 9 2
23 9 12 9 1 0 9 2 9 2 9 7 9 15 13 1 12 0 9 2 0 1 9 2
8 2 13 4 9 7 13 15 2
22 14 2 11 2 14 2 2 13 0 9 11 1 0 11 0 0 9 0 9 11 11 2
13 9 2 12 9 7 9 2 13 9 0 9 11 2
10 1 9 3 15 13 9 7 0 9 2
5 9 1 9 13 2
7 3 3 4 13 10 9 2
41 2 13 4 1 9 11 12 12 9 2 7 3 4 13 10 9 16 1 9 12 2 9 1 9 7 1 9 3 2 16 4 13 13 10 9 2 2 13 11 11 2
14 2 13 16 1 9 1 10 9 3 1 0 9 2 2
10 1 11 7 0 11 13 0 13 9 2
11 9 13 2 16 1 12 9 13 12 9 2
9 9 0 9 7 13 1 9 9 2
43 2 16 4 15 13 10 0 9 2 13 4 13 1 0 9 2 0 1 15 13 0 16 12 9 2 7 13 15 2 9 2 9 7 9 1 9 0 9 2 2 13 11 2
18 2 13 9 2 16 3 13 3 11 2 2 13 1 15 12 1 15 2
29 2 10 9 2 2 13 11 2 2 13 2 16 13 15 1 9 0 9 2 16 13 15 7 10 9 15 15 13 2
24 10 9 13 0 1 0 9 1 11 2 14 13 2 3 3 13 2 16 9 13 16 9 2 2
5 9 1 9 2 12
4 0 9 13 11
2 11 2
17 0 9 1 9 12 9 0 9 13 3 0 9 11 7 9 11 2
9 13 3 0 9 9 7 0 13 2
18 1 0 9 4 9 9 13 1 0 9 9 14 12 9 3 1 11 2
33 1 0 9 11 4 12 7 12 9 13 1 9 9 1 0 9 9 11 2 0 12 9 4 13 7 9 13 1 9 0 0 9 2
12 0 9 9 11 11 1 0 0 9 1 0 9
2 1 9
7 9 4 13 1 9 1 9
3 9 2 12
9 9 0 9 4 13 1 12 12 9
3 9 2 12
2 1 9
7 1 11 4 13 10 0 9
3 9 2 12
1 9
9 9 9 0 0 4 13 1 12 9
3 9 2 12
9 10 9 13 0 2 13 9 11 11
5 11 2 11 2 2
26 12 1 9 3 1 9 1 0 9 11 11 1 9 0 9 13 2 9 15 13 15 2 15 15 13 2
6 13 1 9 0 9 2
11 13 4 15 11 11 2 16 13 10 9 2
7 2 10 0 9 9 13 2
18 3 13 10 9 3 13 1 12 0 2 16 4 15 13 16 9 9 2
19 10 9 15 3 3 13 1 12 2 9 12 2 3 4 15 13 0 9 2
19 13 15 13 10 9 1 9 9 2 13 0 13 10 9 2 9 7 9 2
14 13 3 12 9 1 0 7 10 0 9 13 3 0 2
12 1 15 3 13 0 9 0 9 10 9 2 2
8 11 13 10 9 0 9 0 9
2 11 2
24 11 13 0 0 9 0 9 3 2 16 9 11 13 9 2 16 15 11 13 13 12 0 9 2
22 0 9 1 9 3 13 1 9 11 2 16 4 2 13 3 7 13 0 0 9 2 2
23 9 9 11 11 11 1 9 13 9 9 2 16 15 13 9 2 15 13 13 1 0 9 2
10 9 9 0 9 13 1 2 0 2 2
35 0 9 11 11 13 1 9 3 1 0 9 3 3 2 16 15 9 11 11 13 13 2 16 0 0 0 9 1 3 16 12 9 13 0 2
21 2 2 2 2 11 13 13 2 16 15 13 13 1 0 9 2 2 13 11 11 2
24 0 9 9 11 11 3 13 2 16 0 9 13 13 1 9 9 2 16 11 4 13 0 9 2
4 9 11 13 9
5 11 2 11 2 2
26 0 9 9 11 11 2 15 13 1 0 9 1 0 9 2 15 3 13 1 0 9 1 9 11 11 2
16 9 9 13 1 0 9 9 0 7 0 11 1 9 0 9 2
16 11 3 3 13 1 9 11 7 12 9 13 1 9 9 11 2
13 0 9 13 9 10 9 1 9 11 1 0 9 2
24 0 9 10 9 13 9 9 2 15 13 9 9 1 9 9 7 9 2 1 9 9 0 9 2
41 16 13 1 0 2 0 9 2 1 0 9 2 3 1 9 2 2 13 3 1 0 9 9 11 1 9 2 16 3 1 15 11 13 3 3 0 9 2 16 13 2
8 9 9 13 9 1 0 9 9
5 11 2 11 2 2
21 10 9 0 9 13 9 2 16 9 9 1 9 9 13 15 1 15 13 1 9 2
32 9 2 15 1 9 13 9 2 3 13 9 7 9 9 13 0 9 1 9 9 7 1 15 2 16 4 15 13 1 9 9 2
19 9 9 9 0 9 11 11 13 2 16 13 0 9 9 1 9 12 9 2
11 1 9 13 15 1 15 1 12 9 3 2
16 0 9 3 13 13 9 1 0 9 2 7 0 9 3 13 2
12 9 13 12 0 9 0 9 1 0 14 12 2
26 2 16 4 9 13 13 15 9 2 13 15 9 9 0 1 9 7 13 15 9 2 2 13 11 11 2
19 13 2 16 1 0 9 13 9 9 9 2 7 15 1 15 3 13 9 2
20 9 0 9 9 7 9 11 11 3 13 2 16 4 9 13 1 9 0 9 2
26 0 0 9 4 15 1 15 13 13 1 9 7 1 9 0 0 9 4 15 9 7 9 13 13 3 2
9 2 16 9 9 13 2 2 13 2
11 9 1 0 9 13 3 13 1 9 1 9
7 11 2 11 2 11 2 2
17 9 1 0 9 4 13 1 12 2 9 13 1 9 3 1 9 2
16 0 9 13 13 14 1 9 2 7 15 3 1 9 9 9 2
20 13 15 1 9 2 15 13 9 9 16 0 9 0 9 7 15 13 0 9 2
15 9 13 9 7 1 9 15 13 9 1 9 0 1 9 2
32 9 1 15 2 16 4 9 1 9 3 13 1 9 2 13 9 9 9 9 7 9 2 3 0 9 13 2 7 3 0 9 2
11 9 1 9 3 3 13 9 9 1 9 2
14 9 0 9 13 2 16 13 13 14 1 9 1 9 2
38 0 9 1 11 3 3 13 9 9 1 9 9 2 3 9 1 9 9 0 9 1 12 9 13 7 13 0 0 9 1 9 1 9 7 13 0 9 2
8 0 9 13 3 7 0 9 2
12 0 9 15 3 13 13 10 9 9 1 9 2
19 13 1 9 1 0 9 9 13 0 9 0 9 7 9 1 9 0 9 2
8 11 11 13 1 12 9 9 9
5 11 2 11 2 2
24 9 7 9 2 0 9 11 11 13 3 13 2 16 1 9 2 15 15 3 13 2 13 9 2
8 9 4 13 13 13 12 9 2
5 11 13 12 9 2
18 9 13 3 1 0 9 2 0 9 13 9 9 9 7 0 12 9 2
9 9 13 9 9 9 1 9 11 2
7 15 3 13 3 0 9 2
10 0 9 11 13 9 1 12 12 9 2
15 11 13 1 9 9 12 9 12 9 9 2 9 7 9 2
6 13 3 1 0 9 2
12 1 9 9 11 11 13 11 0 0 9 9 2
10 9 7 13 0 9 1 9 9 9 2
14 13 15 11 13 1 9 0 15 1 9 0 0 9 2
14 3 1 10 9 15 9 1 11 13 7 1 0 9 2
11 0 9 13 1 0 9 9 0 0 9 2
10 10 9 13 1 12 9 3 16 11 2
21 16 1 9 12 11 13 3 12 9 9 9 2 3 9 13 12 7 12 9 9 2
14 11 11 13 0 9 0 9 1 9 1 9 0 9 2
13 0 9 13 1 9 9 1 0 12 1 12 9 2
13 12 15 13 0 9 7 12 9 13 1 0 9 2
19 1 9 13 11 1 10 9 0 9 7 9 15 13 7 1 9 7 9 2
4 0 9 1 11
7 9 1 11 2 11 2 2
24 0 9 0 9 11 11 13 3 1 9 1 9 1 11 1 0 9 11 9 1 9 0 9 2
24 9 0 9 9 13 7 9 9 9 1 9 2 15 13 9 9 1 9 9 9 0 9 11 2
15 9 1 11 15 13 3 9 9 1 10 0 9 1 11 2
10 1 10 9 1 15 13 12 0 9 2
12 1 9 1 9 0 9 3 13 12 0 9 2
7 9 4 13 3 1 9 11
5 11 2 11 2 2
19 1 0 7 0 9 0 2 0 9 13 0 9 0 9 16 1 0 11 2
17 10 9 9 13 9 0 9 2 15 1 9 1 9 13 0 9 2
24 1 9 0 0 9 1 0 7 0 9 1 9 11 9 11 11 13 15 13 9 7 0 9 2
11 0 9 13 3 9 0 9 9 0 9 2
29 2 9 2 15 13 1 11 1 9 0 9 2 13 3 1 9 13 1 9 9 9 0 9 2 2 13 11 11 2
13 2 13 10 9 1 9 4 13 13 1 10 9 2
31 13 15 3 13 2 16 3 4 0 1 9 1 9 9 1 0 9 13 1 15 2 15 1 15 13 1 0 0 9 2 2
18 3 16 1 0 0 9 15 13 13 9 1 0 9 7 11 1 9 2
19 15 13 1 9 14 10 9 2 1 15 0 9 13 0 13 0 9 9 2
15 13 15 13 9 1 9 9 7 9 1 9 9 0 9 2
13 2 9 4 1 10 9 13 1 0 7 0 9 2
27 3 7 1 9 9 0 1 9 4 13 13 2 16 4 1 9 13 3 0 9 9 2 2 13 11 11 2
5 9 1 9 13 9
2 11 2
32 1 9 0 9 2 15 13 1 0 7 0 9 1 9 2 15 13 3 3 9 7 9 13 1 0 9 1 0 7 0 9 2
9 1 9 3 7 15 0 9 13 2
18 2 15 3 13 2 3 15 1 9 13 2 2 13 9 9 11 11 2
13 9 13 1 0 9 3 9 0 1 9 1 9 2
17 0 2 0 9 13 9 9 1 9 2 15 4 13 1 0 9 2
11 9 13 9 11 7 11 0 1 0 11 2
11 9 2 15 3 3 13 9 2 13 11 2
8 1 0 11 3 13 12 9 2
15 2 1 9 9 13 3 9 9 2 2 13 15 9 11 2
19 2 1 0 0 9 15 3 13 3 9 2 15 13 1 11 7 0 9 2
5 3 3 13 2 2
9 3 0 9 15 1 9 13 3 2
17 3 1 9 1 9 13 14 12 9 2 3 14 9 13 1 12 2
9 1 9 13 3 9 0 9 9 2
6 13 13 1 12 9 2
16 12 9 13 0 0 9 2 9 1 11 2 10 9 1 11 2
15 9 13 1 9 9 1 0 9 1 11 2 9 1 11 2
9 9 13 13 1 0 9 1 11 2
6 9 1 9 13 1 11
5 11 2 11 2 2
24 1 0 0 9 1 9 11 1 0 11 13 3 9 12 9 1 9 0 0 9 11 7 11 2
30 10 9 1 15 13 0 9 1 0 9 7 1 10 9 9 9 7 15 9 0 1 9 1 11 13 0 0 9 11 2
19 9 4 13 1 9 9 9 7 9 2 16 1 9 15 13 9 7 9 2
18 3 15 13 9 0 9 11 11 2 11 2 13 4 13 10 9 0 2
7 9 13 1 9 10 0 9
5 11 2 11 2 2
8 9 10 9 15 13 3 13 2
15 3 1 9 7 9 13 13 3 1 0 9 0 0 9 2
18 0 0 9 13 1 11 11 1 0 0 9 1 10 9 1 9 0 2
20 1 9 10 9 13 0 0 9 2 14 3 4 10 9 13 9 0 9 9 2
9 2 13 1 9 9 1 0 9 2
13 16 13 9 9 3 3 2 13 15 9 0 9 2
8 9 13 1 0 9 3 3 2
36 0 9 4 15 3 13 13 3 7 3 2 15 13 0 9 3 1 0 9 2 2 13 11 11 2 10 0 9 1 0 9 3 13 3 3 2
21 1 0 9 2 16 1 9 13 4 0 9 1 12 9 11 2 9 3 13 9 2
5 2 13 15 0 2
8 0 9 4 13 14 9 9 2
19 15 7 13 2 16 0 9 4 1 9 13 2 14 9 9 13 0 2 2
9 13 13 15 9 1 12 2 9 2
19 9 13 2 16 13 2 14 1 0 11 2 13 15 1 0 7 0 9 2
14 7 0 9 3 13 2 16 15 9 13 2 9 13 2
2 13 9
15 0 9 13 9 9 2 16 13 9 9 3 2 16 13 9
5 11 2 11 2 2
8 3 9 9 9 13 0 9 2
10 0 9 13 3 9 2 16 13 9 2
12 0 9 1 9 9 15 13 7 1 0 9 2
39 9 0 0 9 1 11 2 15 13 9 9 1 9 11 2 0 9 2 11 2 11 7 11 3 1 2 0 2 9 13 10 9 1 9 1 12 12 9 2
19 9 0 9 9 9 7 9 13 3 0 7 3 14 3 0 16 9 9 2
20 9 3 13 2 16 9 13 0 9 2 3 9 2 15 13 7 4 3 13 2
13 1 0 9 9 3 9 13 7 10 9 15 13 2
10 3 0 0 9 9 13 12 9 9 2
13 1 9 9 9 4 0 9 13 1 0 0 9 2
3 9 1 9
2 11 2
29 12 9 1 11 2 15 9 13 1 9 1 9 3 11 11 1 9 13 0 9 0 0 9 2 13 3 1 9 2
29 0 9 2 15 13 1 12 9 2 4 13 1 0 9 9 7 9 9 7 13 15 9 9 9 12 7 12 9 2
17 9 2 15 0 9 3 13 16 3 0 2 4 13 1 0 9 2
27 9 13 1 15 12 0 9 2 15 15 13 13 1 9 12 9 1 12 9 2 7 2 12 9 1 9 2
6 3 15 13 1 9 2
17 1 0 11 13 15 1 0 12 9 3 0 9 9 2 13 9 2
3 9 9 13
5 11 2 11 2 2
13 9 9 1 9 15 3 13 13 1 9 7 9 2
17 3 3 13 1 0 9 2 15 1 0 9 13 1 10 0 9 2
13 0 9 3 13 1 0 9 7 9 13 1 9 2
15 10 9 13 1 0 13 7 16 9 15 2 15 13 9 2
10 2 13 2 13 3 9 9 0 9 2
8 0 9 13 7 9 10 9 2
10 0 0 9 13 7 0 9 0 9 2
21 3 13 7 1 0 9 2 3 0 9 13 1 0 9 1 0 9 1 0 9 2
7 0 1 9 0 9 13 13
8 0 9 13 1 12 9 9 9
5 11 2 11 2 2
25 1 9 1 9 0 9 7 0 9 10 9 1 9 3 1 11 12 13 9 1 9 3 12 9 2
19 0 11 11 2 13 1 9 1 0 9 1 9 11 11 0 9 11 11 2
17 0 9 7 10 9 3 13 2 16 13 0 9 7 9 10 9 2
20 9 9 15 15 3 9 1 9 1 9 9 12 9 13 2 3 2 3 13 2
15 1 9 0 9 12 9 15 13 0 9 9 2 11 11 2
10 1 10 9 13 13 12 9 9 9 2
17 9 1 9 13 0 9 2 15 1 10 9 13 9 12 9 9 2
14 9 9 13 0 9 11 11 2 2 15 9 3 13 2
22 11 11 2 13 9 1 9 2 0 0 9 15 4 13 1 9 7 9 1 0 9 2
9 1 15 13 9 9 1 9 9 2
19 12 1 0 9 2 15 13 3 0 1 9 9 2 7 9 13 1 9 2
18 1 9 13 13 2 16 4 13 0 9 2 15 4 1 9 9 13 2
10 1 9 9 13 1 9 3 12 9 2
4 9 1 9 2
10 3 7 3 13 1 9 2 3 9 2
19 0 0 9 12 7 12 9 2 9 2 0 0 12 7 12 9 2 9 2
10 9 1 12 9 1 12 9 2 9 2
11 0 7 0 9 12 7 12 9 2 9 2
4 9 7 9 2
14 3 1 9 2 3 7 9 2 1 9 13 1 9 2
31 0 0 9 1 9 12 7 12 9 2 9 2 1 9 12 7 12 9 2 9 2 0 0 9 12 7 12 9 2 9 2
17 9 2 9 9 1 0 9 1 10 9 13 12 5 1 0 9 2
11 9 2 0 9 0 2 0 9 3 0 2
33 1 9 13 9 1 12 2 12 7 13 1 12 2 12 2 9 13 1 9 1 12 2 12 7 13 1 12 2 12 9 0 9 2
3 9 9 2
20 0 9 12 9 2 9 13 1 9 12 2 0 12 9 2 9 1 9 12 2
8 0 0 9 12 9 2 9 2
3 9 1 9
3 11 1 11
2 11 2
22 0 9 12 2 0 9 11 11 13 12 9 1 9 0 9 11 11 1 0 11 11 2
19 9 12 9 13 9 0 0 9 11 2 15 13 3 1 12 2 11 11 2
3 9 1 11
2 11 2
25 1 0 9 0 9 1 0 9 1 11 13 9 0 9 1 11 12 2 12 2 12 2 12 2 2
8 9 12 9 0 9 13 11 2
29 13 15 1 0 9 2 0 9 1 3 0 9 1 15 9 13 0 9 1 0 9 2 3 3 13 1 10 9 2
15 1 9 9 13 10 9 1 9 1 9 1 9 1 11 2
5 1 9 1 0 9
8 0 11 13 12 2 9 1 11
2 11 2
23 1 9 0 9 0 11 1 0 11 4 3 13 1 9 12 9 0 12 2 9 10 9 2
19 9 9 11 13 12 2 9 0 9 0 9 1 0 9 1 11 1 11 2
14 0 9 12 2 9 13 0 9 1 9 2 0 11 2
4 0 0 9 2
35 0 9 13 1 12 0 9 0 9 9 7 9 2 9 9 2 11 2 11 2 11 2 11 2 1 11 2 11 2 7 1 10 0 9 2
11 1 11 13 13 1 9 3 12 0 9 2
21 9 0 9 13 1 0 9 11 9 12 0 9 7 0 9 1 9 12 0 9 2
11 3 13 9 9 0 9 3 12 0 9 2
19 1 9 4 13 0 9 0 9 1 11 2 0 16 12 1 0 1 9 2
24 9 1 9 9 9 1 11 4 1 0 9 13 1 9 12 1 9 0 0 9 2 11 2 2
3 9 11 11
5 0 0 9 15 13
14 15 2 15 13 1 9 2 9 11 2 2 13 0 9
2 11 2
27 1 9 0 9 11 0 1 9 9 15 13 7 0 9 0 0 9 2 15 15 0 9 13 1 0 9 2
41 0 9 13 9 9 11 13 9 1 15 9 9 12 2 9 11 7 3 9 9 0 9 11 2 15 7 9 11 13 3 1 12 9 3 2 9 2 9 2 2 2
35 1 0 9 11 11 13 9 11 11 1 9 9 9 7 1 0 9 11 2 13 9 9 11 11 11 1 0 9 1 9 9 0 9 11 2
68 0 9 11 3 1 0 9 13 9 1 9 1 15 9 9 9 2 15 13 1 9 1 9 9 11 13 1 9 9 9 12 2 9 2 3 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 7 11 11 2 15 0 9 3 13 9 7 1 9 9 9 2
37 1 10 9 0 9 13 13 3 13 9 0 9 7 10 9 13 0 9 0 0 9 1 12 2 12 2 12 2 3 7 1 12 2 12 2 12 2
4 1 9 13 9
11 10 0 9 1 9 13 1 9 10 9 2
19 15 2 16 13 0 7 9 3 13 9 0 9 1 9 2 15 13 9 2
21 0 0 9 3 13 13 14 9 9 1 11 2 7 7 0 9 1 9 0 9 2
17 1 0 9 1 9 7 9 2 11 2 13 0 9 13 0 9 2
15 13 15 2 16 9 13 13 1 0 9 0 16 1 0 2
31 15 2 16 9 9 1 9 4 3 13 0 9 12 9 7 10 10 9 13 1 0 9 14 12 9 2 13 10 9 13 2
11 9 13 2 16 3 1 10 9 13 13 2
25 7 13 0 2 16 16 13 9 0 9 2 15 13 10 9 2 13 4 9 13 13 3 0 9 2
23 9 13 0 0 9 1 9 2 15 13 1 0 9 9 7 0 1 15 2 15 9 13 2
8 13 3 1 0 7 0 9 2
14 9 4 15 3 13 13 9 13 0 9 1 0 9 2
15 9 2 15 13 9 7 1 0 9 2 13 3 3 13 2
20 14 3 13 7 9 13 2 16 13 9 0 9 2 15 10 0 9 13 9 2
18 1 9 9 13 15 2 16 1 9 9 1 0 9 13 0 0 9 2
28 16 9 13 13 0 9 1 9 2 15 13 2 7 0 1 9 0 2 13 15 9 2 15 10 9 3 13 2
6 10 9 9 3 13 2
10 9 15 7 13 13 1 9 13 3 2
10 3 9 0 9 2 7 0 0 9 2
19 9 10 0 9 3 13 9 0 7 3 0 2 7 15 10 9 3 13 2
3 9 9 13
36 9 0 9 2 1 15 9 9 0 3 0 9 13 9 0 9 2 13 3 0 7 0 9 2 1 15 4 9 0 13 9 0 9 0 9 2
24 7 9 2 0 1 15 2 3 9 7 9 13 2 0 1 0 9 2 15 1 9 13 13 2
23 1 0 9 15 3 3 13 14 9 9 2 3 3 9 9 2 15 4 9 13 1 9 2
14 13 0 9 0 9 0 9 13 1 0 0 9 0 2
25 0 9 1 15 2 15 3 13 2 13 2 1 9 9 2 3 9 13 1 0 2 9 1 9 2
10 3 13 0 9 13 7 10 9 13 2
30 10 9 4 13 3 1 0 9 7 3 2 13 2 14 10 9 9 2 16 4 3 3 13 9 13 2 3 4 13 2
11 1 0 9 7 1 9 1 9 15 13 2
17 9 1 9 0 9 0 9 11 1 0 9 0 9 13 10 9 2
19 1 9 4 13 13 9 1 9 9 2 3 0 1 0 9 1 7 1 2
12 9 2 3 0 10 9 2 15 13 1 9 2
4 9 0 9 13
7 9 13 2 13 7 13 2
9 9 13 15 13 3 13 1 9 2
22 3 1 3 0 9 0 9 16 0 9 13 0 2 16 13 3 3 0 16 9 15 2
14 9 15 3 1 9 9 13 3 3 0 7 3 0 2
24 1 10 0 9 13 16 0 9 9 2 0 9 15 3 13 7 3 15 13 9 1 9 9 2
4 9 13 15 2
15 9 7 9 0 9 2 9 0 9 7 0 9 0 9 2
13 13 15 9 0 9 7 0 9 9 2 1 0 2
46 1 12 2 9 12 15 1 0 11 13 0 2 16 0 9 13 0 2 3 7 9 2 16 4 13 0 0 9 2 7 3 9 9 2 15 15 13 9 1 0 9 2 13 16 9 2
23 1 0 9 10 9 3 13 2 16 0 9 13 14 0 9 2 7 3 9 1 0 9 2
23 9 1 11 3 1 9 0 0 7 9 13 9 0 9 2 15 3 1 3 0 0 9 2
11 1 12 2 9 7 10 9 13 0 9 2
16 9 1 10 9 13 9 0 9 7 9 7 0 9 0 9 2
15 0 9 13 3 0 9 2 0 3 14 1 0 0 9 2
14 1 10 9 13 14 1 0 9 11 12 7 12 9 2
32 13 15 14 0 9 1 0 9 7 9 1 9 2 7 7 9 1 9 7 9 0 7 0 9 2 15 13 16 9 1 9 2
15 0 9 0 9 9 13 1 0 9 1 0 7 0 11 2
31 9 1 10 9 13 2 0 9 0 9 3 13 9 9 2 7 3 15 9 7 9 1 9 10 9 13 13 2 3 13 2
24 0 1 9 13 9 11 1 11 2 1 9 15 13 7 11 2 15 3 13 0 9 0 9 2
31 9 13 7 1 0 9 2 7 3 7 1 0 9 2 15 15 9 9 11 11 3 1 10 9 1 9 13 13 2 3 2
27 3 0 2 0 9 3 13 9 10 0 9 2 15 13 13 9 2 3 7 0 9 2 16 15 9 13 2
29 13 15 10 9 9 2 16 14 9 2 7 7 9 9 3 13 2 16 15 13 1 15 13 15 1 9 13 9 2
12 1 9 1 9 13 9 13 2 3 13 9 2
11 13 15 3 1 9 2 3 7 1 9 2
43 16 9 13 0 9 13 3 0 2 16 9 1 0 9 13 3 0 9 1 0 9 2 13 15 9 2 16 0 9 2 16 13 0 9 0 9 2 1 0 9 0 13 2
10 9 13 0 13 2 16 13 15 13 2
8 16 13 9 2 13 7 9 2
6 7 9 15 13 3 2
7 9 0 9 13 7 1 9
3 9 13 9
32 11 11 2 9 0 0 9 2 15 1 9 12 13 0 9 1 0 9 14 1 0 9 11 2 13 1 10 9 1 9 9 2
23 9 11 13 2 16 1 9 0 9 13 0 3 13 2 11 13 9 2 7 7 13 13 2
17 9 13 3 0 9 9 2 3 0 16 0 9 7 9 1 11 2
25 1 9 2 15 13 3 0 16 10 10 2 13 9 9 7 9 0 2 15 15 1 0 9 13 2
20 1 10 0 9 13 15 2 16 13 9 9 9 2 3 16 12 9 3 0 2
12 3 0 0 9 7 9 11 13 9 0 9 2
37 1 12 2 9 3 13 9 9 2 15 1 9 3 13 2 1 0 0 9 15 7 2 3 13 9 0 9 2 9 9 1 0 9 13 1 9 2
16 9 1 15 13 0 9 2 15 13 0 9 1 9 0 9 2
15 11 11 13 1 9 2 16 13 0 9 0 9 0 9 2
47 1 0 9 1 9 11 2 3 15 7 1 9 13 2 16 13 0 9 2 16 9 2 13 2 1 3 0 9 2 1 9 10 9 2 3 0 9 11 13 3 3 7 3 2 16 13 2
6 9 4 13 0 9 2
7 15 9 13 3 3 13 2
21 9 9 13 3 13 2 16 9 4 3 13 3 1 0 7 0 9 7 0 9 2
17 3 9 13 1 9 1 15 2 16 9 13 10 9 2 3 3 2
20 16 9 7 9 13 13 9 0 9 7 9 2 0 9 13 13 1 9 9 2
4 9 13 0 9
24 9 1 3 0 9 13 0 9 1 0 7 0 9 0 9 7 0 9 1 9 0 0 9 2
19 9 9 9 7 9 9 0 1 9 0 9 7 9 0 9 15 13 3 2
20 12 2 0 9 0 0 9 3 1 0 9 9 2 3 7 1 10 0 9 2
19 0 9 15 9 13 14 3 7 3 2 3 3 1 9 0 9 0 9 2
21 12 2 0 9 9 1 0 9 7 0 9 9 3 0 9 9 1 9 0 9 2
16 12 2 9 1 9 7 9 0 9 1 9 9 1 0 9 2
42 1 0 9 13 13 7 12 0 9 2 1 0 9 13 0 9 7 0 0 9 12 9 7 3 0 0 9 2 3 2 16 10 0 9 3 3 13 0 9 7 9 2
10 12 2 0 9 0 9 1 0 9 2
31 13 13 9 9 0 1 9 0 9 2 9 9 1 0 9 0 7 0 0 9 13 13 2 16 4 15 13 10 0 9 2
18 12 2 9 9 1 0 2 0 7 0 9 7 9 1 10 0 9 2
53 9 7 9 13 9 2 16 14 0 9 0 9 1 0 11 2 1 11 2 1 11 7 3 2 0 1 0 0 7 0 9 0 9 7 1 0 9 1 9 2 9 2 7 9 0 9 2 13 13 9 1 9 2
23 0 9 1 9 9 0 9 13 10 9 9 1 0 9 2 15 13 0 0 9 0 9 2
39 12 2 9 0 9 0 1 9 0 9 2 9 0 9 7 9 0 9 2 9 1 3 0 0 9 2 1 0 9 9 9 7 9 9 1 9 9 9 2
17 13 0 13 1 9 2 16 9 0 9 4 3 13 1 9 0 2
38 12 2 9 0 9 0 1 0 9 1 9 0 9 2 1 9 12 1 12 9 1 9 1 0 9 7 13 2 14 1 9 9 2 3 3 3 2 2
24 12 2 9 0 9 0 1 9 1 0 9 7 1 9 9 3 0 9 1 0 7 0 9 2
44 12 2 0 9 9 0 9 2 10 0 9 1 9 7 0 9 1 9 0 9 2 15 15 13 3 2 15 2 16 0 9 9 13 11 14 1 12 2 9 9 0 9 2 2
36 11 3 9 9 1 9 0 9 13 1 0 9 0 3 3 13 0 0 9 7 13 9 9 0 2 9 10 9 1 9 9 15 13 9 9 2
47 12 2 0 0 9 10 0 9 2 1 9 9 2 2 15 13 2 7 3 13 9 9 0 9 0 9 7 3 13 9 0 9 9 0 1 0 2 0 7 0 9 9 7 9 0 9 2
52 0 9 0 9 9 7 9 1 0 9 13 3 0 2 15 13 14 1 0 9 9 0 9 2 3 0 9 9 9 2 2 7 3 1 9 0 9 0 3 1 0 9 9 7 0 9 9 0 1 9 9 2
21 13 7 3 13 1 15 2 16 9 1 0 9 13 13 0 9 9 0 0 9 2
24 9 9 0 0 9 1 9 9 7 9 0 9 1 9 7 10 0 9 13 9 10 0 9 2
19 0 9 2 0 9 7 0 9 2 1 9 0 2 3 13 10 9 9 2
8 7 0 9 13 9 7 9 2
16 13 2 16 15 10 9 13 7 10 0 9 1 0 9 13 2
9 9 9 0 0 4 13 1 12 9
8 9 13 13 15 3 0 9 2
15 13 15 4 7 1 9 9 1 0 9 7 9 0 9 2
28 9 0 0 4 13 0 7 0 2 9 1 9 11 1 9 2 1 12 9 2 1 9 9 0 9 13 0 2
10 0 9 4 9 13 1 12 2 9 2
16 0 9 1 9 9 4 13 13 0 16 12 9 1 9 9 2
21 9 9 4 13 1 9 0 1 9 12 9 9 9 9 2 15 9 13 9 13 2
4 9 1 9 0
20 9 13 1 0 9 9 9 11 11 0 9 9 9 7 9 0 7 0 9 2
7 1 9 15 13 12 9 2
33 0 9 0 9 7 9 13 12 9 9 2 1 15 1 0 9 4 13 9 7 9 1 12 9 9 7 1 11 1 12 9 9 2
20 0 0 9 9 1 11 15 3 13 1 12 9 7 1 11 1 12 9 9 2
27 2 16 15 1 0 9 3 12 9 0 0 9 13 3 12 13 2 13 15 1 9 2 2 13 11 11 2
32 2 1 12 9 9 0 0 9 13 9 9 1 0 9 12 9 1 12 9 9 0 9 2 15 13 3 0 9 2 2 13 2
7 1 11 13 9 12 9 2
19 1 11 15 1 9 13 12 9 2 15 13 3 12 9 1 12 12 9 2
11 10 9 13 1 9 9 1 12 9 9 2
20 1 3 0 9 0 9 0 9 1 9 9 9 4 1 9 9 13 12 9 2
3 9 13 9
2 11 2
19 9 0 7 0 9 2 9 2 13 0 9 1 9 0 0 7 0 9 2
10 3 1 0 9 15 13 9 11 11 2
26 13 2 16 0 12 9 0 9 7 9 11 2 15 9 13 2 1 9 0 9 4 13 13 0 9 2
33 0 9 13 2 16 9 1 0 0 9 12 9 9 4 13 1 9 2 1 0 12 9 9 15 13 14 3 1 9 1 9 12 2
9 9 13 9 1 11 1 9 12 2
35 0 9 12 9 1 0 9 12 9 1 0 9 0 2 9 13 1 0 9 12 9 2 1 0 9 4 0 9 13 1 12 7 12 9 2
4 1 11 0 9
2 11 2
18 9 13 1 11 1 9 1 9 9 1 12 9 2 12 9 2 3 2
14 0 9 3 13 9 1 0 9 1 12 1 12 9 2
32 9 0 9 2 12 9 2 4 13 1 12 9 2 14 12 9 2 2 0 9 0 9 1 9 12 9 2 14 12 9 2 2
22 0 9 13 13 13 12 2 9 7 4 15 13 14 1 12 9 2 14 12 9 2 2
29 1 11 13 0 9 0 1 0 9 3 0 9 2 11 2 11 2 16 1 0 9 2 9 2 11 2 11 2 2
8 11 2 11 7 11 13 0 9
2 11 2
19 9 12 0 9 0 9 2 11 2 11 7 11 2 13 9 1 0 9 2
39 13 2 16 1 12 2 9 0 9 4 13 9 2 1 9 0 9 2 2 1 15 15 4 13 13 7 0 0 0 9 7 15 4 1 9 13 0 9 2
19 9 15 12 9 13 2 16 9 11 2 11 7 11 13 9 0 0 9 2
18 13 15 1 9 15 9 1 0 0 7 0 9 7 1 9 0 9 2
16 13 1 0 13 1 9 9 2 0 9 7 0 7 0 9 2
6 1 11 1 9 0 9
2 11 2
11 9 13 3 0 1 9 1 0 0 9 2
9 0 9 15 3 13 1 11 3 2
26 1 9 15 9 9 13 1 12 9 2 14 12 9 2 7 1 9 1 12 9 2 0 12 9 2 2
5 0 9 3 1 9
7 11 2 11 2 11 2 2
26 0 9 2 11 2 13 1 0 9 2 3 15 13 0 9 2 1 9 9 9 1 9 12 9 9 2
15 9 15 1 9 13 1 9 0 9 7 0 7 0 9 2
6 13 1 9 0 9 2
17 1 0 9 9 1 0 2 9 4 13 12 9 11 1 12 9 2
29 0 9 2 1 10 9 13 13 9 1 0 9 2 13 13 1 12 7 12 9 1 12 9 1 0 9 12 9 2
4 0 9 1 11
2 11 2
19 1 11 4 13 13 0 7 0 9 2 15 4 13 0 9 7 13 9 2
18 13 13 0 9 12 9 9 2 13 7 3 0 2 15 15 15 13 2
21 13 4 13 9 9 0 0 11 2 10 9 4 13 1 9 0 0 7 0 9 2
9 0 9 0 1 12 2 12 2 12
2 9 9
8 9 9 9 9 9 9 9 9
4 15 1 12 9
6 9 12 2 12 2 12
3 9 9 9
4 15 1 12 9
6 9 12 2 12 2 12
12 9 9 1 0 9 13 13 0 9 7 0 9
2 11 2
20 14 1 12 9 4 15 13 13 0 0 9 7 9 2 0 9 7 0 9 2
19 13 15 1 9 9 1 9 1 0 9 2 15 12 2 9 13 1 9 2
8 0 9 4 13 13 1 9 2
9 3 13 1 9 9 2 3 9 2
15 9 3 10 9 13 1 9 9 0 12 9 1 9 0 2
45 1 15 4 3 1 9 13 3 0 9 2 0 9 2 9 1 9 2 0 2 0 2 0 7 0 9 2 9 0 9 7 9 2 9 7 9 1 9 9 7 0 9 7 9 2
17 3 9 7 9 0 9 15 13 1 9 12 9 1 9 12 9 2
16 9 7 3 7 9 13 1 10 9 1 9 3 1 0 9 2
22 9 0 9 2 3 1 9 0 9 2 7 13 3 1 0 0 7 0 9 16 3 2
15 10 9 3 10 9 13 16 9 1 2 3 0 9 2 2
8 1 15 0 9 12 9 13 2
22 7 9 13 2 16 9 10 9 1 0 9 13 0 3 1 0 9 0 9 1 15 2
36 0 9 3 9 7 9 13 0 0 9 1 9 2 9 7 0 0 9 7 9 9 1 0 9 2 15 13 9 1 0 9 1 3 0 9 2
27 1 12 1 12 9 15 3 7 13 7 9 2 15 1 0 9 13 13 2 3 0 9 2 9 7 9 2
13 3 15 9 1 9 1 9 0 9 13 3 0 2
18 1 9 12 9 1 0 13 3 13 9 7 9 1 0 9 7 9 2
22 13 1 15 3 13 0 9 2 15 3 13 9 12 9 2 1 9 1 9 7 9 2
23 9 4 1 0 9 13 9 9 1 0 9 14 1 12 2 9 0 9 1 9 0 9 2
8 3 15 13 1 12 2 9 2
21 0 9 3 4 13 3 1 10 9 13 9 1 0 9 14 12 7 12 9 9 2
23 9 9 1 9 1 0 9 3 13 9 0 9 2 15 13 0 0 9 0 1 9 9 2
14 13 9 13 0 9 1 12 9 1 9 9 0 9 2
19 3 13 7 3 13 9 9 0 0 9 1 9 0 9 1 9 1 0 2
13 10 9 13 0 1 9 1 9 12 9 1 9 2
28 1 10 9 13 4 3 13 9 9 9 2 13 0 13 9 9 1 9 2 9 7 9 9 0 7 0 9 2
33 3 1 0 9 2 3 0 9 13 9 0 1 9 9 1 0 9 0 9 2 13 9 0 3 1 0 9 9 9 1 0 9 2
22 0 15 13 1 12 9 2 1 12 9 2 2 0 1 12 9 2 1 12 9 2 2
28 10 9 13 0 9 1 0 9 2 3 13 3 9 0 9 0 9 9 3 0 2 12 9 13 1 9 0 2
5 11 2 11 2 2
24 0 9 1 0 9 9 2 9 2 2 1 15 15 0 0 9 13 3 0 0 9 2 13 2
27 1 9 1 12 9 2 12 9 7 12 9 2 0 1 9 2 13 9 9 1 9 9 12 7 12 9 2
17 9 13 1 0 9 9 2 15 15 1 9 13 1 12 2 9 2
23 1 10 9 3 0 0 9 3 2 13 0 9 9 9 2 15 1 15 13 13 3 13 2
23 16 9 1 9 13 3 0 9 2 13 4 9 9 13 1 9 9 2 1 15 13 9 2
8 9 9 7 9 13 1 11 3
7 1 9 15 13 12 9 2
26 2 1 12 9 9 0 0 9 13 9 9 12 9 1 12 9 9 0 9 2 15 13 3 0 9 2
8 2 1 11 13 9 12 9 2
19 1 11 15 1 9 13 12 9 2 15 13 3 12 9 1 12 12 9 2
11 10 9 13 1 9 9 1 12 9 9 2
22 1 3 0 9 0 9 0 9 1 9 12 9 9 4 1 9 9 13 12 9 9 2
19 9 0 9 9 1 3 0 9 13 1 12 9 0 9 0 1 12 9 2
6 0 7 0 9 13 9
2 11 2
19 9 0 7 0 9 2 9 2 13 0 9 1 9 0 0 7 0 9 2
11 1 0 0 9 15 13 10 9 11 11 2
32 1 10 9 13 1 9 2 16 0 12 9 0 9 7 9 11 2 15 9 13 2 3 1 9 0 9 4 13 13 0 9 2
21 0 9 13 2 16 9 1 0 0 9 1 9 12 9 9 4 13 1 0 9 2
17 1 0 12 9 9 9 15 4 13 14 3 1 9 1 9 12 2
10 9 9 13 9 1 11 1 9 12 2
31 3 0 0 9 13 7 3 12 9 9 9 2 1 9 12 0 9 13 12 9 9 7 3 12 9 9 13 12 0 9 2
16 12 9 9 4 13 1 9 7 0 3 12 9 13 3 13 2
35 0 9 12 9 1 0 9 12 9 1 0 9 0 2 9 13 1 0 9 12 9 2 1 0 9 13 0 9 13 1 12 7 12 9 2
16 0 0 9 13 0 9 1 9 9 1 9 12 1 0 9 2
19 1 9 13 0 9 1 12 1 12 9 2 13 15 7 13 7 0 9 2
7 13 9 12 2 12 12 2
32 0 9 1 0 12 1 11 13 1 12 2 12 2 1 0 0 9 9 9 1 9 3 1 9 2 15 13 9 1 0 9 2
12 0 13 13 0 9 9 0 9 1 12 9 2
18 0 0 9 1 9 9 0 9 1 11 13 1 0 0 0 9 1 9
3 9 1 9
5 11 2 11 2 2
14 9 0 9 0 0 9 13 1 9 9 1 0 9 2
19 0 9 0 9 1 15 13 9 1 0 11 1 0 0 9 1 0 9 2
10 1 9 13 1 9 0 9 9 12 2
23 9 13 9 1 9 0 11 1 0 9 7 0 9 1 9 2 13 13 3 0 0 9 2
16 1 0 11 15 1 0 9 13 1 9 9 0 0 9 11 2
31 1 11 11 1 0 9 7 0 9 11 7 9 3 13 0 9 1 9 2 16 9 0 9 3 4 13 1 0 0 9 2
7 9 11 13 9 1 0 9
5 11 2 11 2 2
16 0 9 1 9 0 9 1 11 13 1 12 1 10 0 9 2
30 9 9 9 9 7 0 12 3 0 9 13 9 11 11 11 1 0 9 1 9 2 15 1 9 3 13 1 0 9 2
8 13 15 3 1 0 0 9 2
12 10 9 13 9 0 0 9 9 2 11 11 2
26 1 15 13 1 9 1 9 0 0 9 7 4 13 7 0 9 2 16 4 15 3 3 13 9 9 2
12 9 13 0 2 7 16 13 0 9 7 9 2
14 1 11 2 11 13 0 3 9 1 0 0 9 9 2
28 3 13 2 13 11 1 9 3 0 9 1 9 0 9 7 9 9 2 7 0 9 12 12 9 13 3 0 2
18 2 9 15 13 3 12 12 9 2 7 13 3 3 2 16 13 9 2
10 1 9 4 3 13 2 2 13 9 2
17 11 13 16 9 1 9 2 0 2 1 9 0 1 0 9 0 2
20 1 9 13 1 3 16 9 9 2 1 15 15 1 9 0 9 13 0 9 2
16 15 3 13 9 1 0 9 2 15 13 9 1 9 7 9 2
5 11 13 9 1 9
38 9 12 2 9 1 0 9 3 3 13 9 0 9 7 9 2 1 10 9 3 9 11 11 13 1 9 1 9 11 0 2 0 9 0 9 11 12 2
17 0 9 3 13 0 2 7 0 9 15 15 13 3 3 7 3 2
27 0 9 7 9 13 13 3 1 9 3 2 10 9 1 9 3 12 9 2 15 13 1 0 0 11 13 2
24 1 9 2 15 13 1 0 9 1 0 9 2 15 1 0 9 1 9 13 9 7 0 9 2
7 1 9 9 3 13 11 2
53 3 16 12 9 1 10 0 9 13 3 9 1 11 0 16 0 9 3 2 13 15 9 1 9 12 2 3 9 11 1 9 13 9 1 0 11 13 1 9 0 9 9 2 15 13 11 0 9 1 9 10 9 2
18 9 3 15 13 2 3 13 1 9 9 2 16 15 11 13 1 9 2
31 3 10 9 2 16 13 1 11 3 9 2 1 15 15 13 3 3 9 2 1 0 9 3 13 2 7 13 3 3 0 2
21 1 0 12 9 13 11 0 9 11 1 0 9 2 1 15 13 0 9 1 11 2
28 3 2 3 15 9 11 13 3 3 9 7 9 1 15 11 7 14 3 1 11 2 7 3 7 10 9 13 2
10 2 15 13 15 3 1 10 11 2 2
37 2 3 4 15 13 13 0 9 2 15 1 0 9 1 11 2 15 9 15 1 9 0 13 7 12 0 9 2 13 1 9 9 1 9 0 11 2
30 0 0 9 1 9 7 0 9 1 11 10 9 3 13 2 3 1 1 0 9 2 1 15 15 11 3 0 9 13 2
14 11 15 3 13 9 2 15 13 13 1 0 9 0 2
12 11 0 9 13 1 10 0 9 12 9 9 2
27 9 0 9 1 11 13 11 3 12 9 9 2 14 1 0 9 4 1 9 9 0 9 13 12 9 9 2
16 9 15 13 7 1 12 9 2 15 13 13 9 1 0 11 2
21 11 15 13 13 2 13 3 2 3 0 2 0 7 3 0 16 3 1 9 2 2
18 10 9 13 9 9 3 7 0 9 0 9 1 11 9 9 11 11 2
30 3 3 0 9 3 13 9 1 9 1 9 2 1 15 11 13 12 0 9 16 9 14 1 15 2 16 13 0 9 2
18 11 13 0 2 16 0 9 11 12 2 13 1 9 0 0 9 11 2
16 10 9 2 11 12 2 2 13 1 0 9 10 0 0 9 2
6 15 10 9 3 13 2
24 1 0 9 15 15 1 9 1 0 9 13 3 3 2 3 1 0 9 2 15 1 15 13 2
17 13 3 3 13 2 16 13 0 16 11 2 0 1 10 0 9 2
24 0 9 15 13 2 16 15 3 3 13 2 16 13 2 14 12 9 2 4 0 3 3 13 2
28 3 15 7 11 15 10 9 3 13 2 7 0 9 13 13 0 9 2 16 15 13 3 0 9 3 0 9 2
22 9 1 11 3 3 3 13 9 1 9 2 15 15 1 9 9 9 1 11 3 13 2
2 11 11
27 0 9 15 1 10 9 9 13 2 7 3 3 0 13 2 13 2 14 15 3 1 9 7 9 1 9 2
7 13 15 1 9 0 9 2
2 11 11
3 9 2 9
4 0 9 1 11
19 0 9 9 15 13 1 9 1 11 1 0 9 2 3 4 13 9 9 2
33 0 9 1 9 0 9 2 3 15 13 2 13 9 0 9 2 15 13 1 9 12 2 9 9 2 3 13 3 9 0 9 11 2
39 0 9 1 9 2 15 15 4 13 14 1 9 0 9 2 15 13 13 3 3 7 13 3 10 9 2 16 13 14 9 2 16 4 13 1 0 0 9 2
8 0 9 11 3 13 9 1 9
40 13 15 0 2 7 7 1 3 12 9 9 0 9 15 13 0 9 11 11 11 13 10 0 7 0 9 2 16 0 7 0 9 1 10 9 15 3 3 13 2
36 0 9 11 1 0 9 1 11 13 11 1 9 2 15 13 3 2 11 7 11 2 3 0 9 7 0 9 3 7 3 13 0 7 0 9 2
15 9 11 1 10 3 0 0 9 13 3 0 9 16 3 2
35 13 0 9 2 3 13 0 9 2 7 1 9 1 9 9 7 3 0 0 9 13 0 9 2 15 13 1 9 13 9 2 0 9 2 2
31 3 0 9 7 10 9 11 11 4 10 9 13 1 0 9 2 3 13 13 10 0 0 9 2 16 1 15 13 0 9 2
15 4 15 3 13 9 1 0 7 3 0 9 1 0 9 2
13 15 11 11 4 3 13 0 0 9 1 10 9 2
18 13 15 3 2 16 0 11 15 13 1 0 9 1 9 9 0 9 2
38 1 11 1 15 13 7 9 1 11 2 3 4 3 13 9 11 3 1 9 2 3 15 11 11 1 11 13 13 9 1 0 9 0 9 7 0 9 2
45 16 13 1 11 2 7 0 0 9 0 0 9 9 1 9 7 0 9 2 15 3 13 9 1 9 2 7 0 9 0 9 3 13 0 0 9 9 7 9 0 9 9 10 9 2
41 3 15 13 2 16 11 13 0 0 9 13 1 15 2 16 4 15 13 9 0 9 7 0 9 9 7 9 13 9 0 7 0 9 7 1 15 7 9 0 9 2
7 0 9 13 2 0 13 3
10 9 0 0 9 15 9 13 1 9 2
27 10 9 0 1 9 1 0 0 9 7 9 1 0 9 15 7 3 13 1 9 2 0 0 15 9 9 2
33 0 9 2 1 15 15 1 0 9 13 7 13 0 0 9 2 4 13 9 7 1 9 9 12 2 9 12 3 13 1 12 9 2
19 3 9 0 9 13 1 0 0 9 9 1 14 10 9 9 0 0 9 2
26 3 1 11 2 3 13 1 9 13 9 0 9 2 13 7 10 9 7 13 3 1 9 2 1 9 2
10 15 10 7 1 10 9 1 9 13 2
11 14 9 15 7 0 9 1 12 2 9 2
14 9 11 3 13 1 12 9 9 2 0 1 10 9 2
20 9 1 15 3 13 7 9 13 15 3 14 0 9 1 10 9 1 0 9 2
23 3 2 16 15 13 11 2 7 3 7 0 11 2 13 11 3 0 3 0 9 1 9 2
30 0 9 13 2 16 12 11 13 9 9 12 9 1 9 2 13 15 1 9 9 7 1 0 9 9 1 9 1 9 2
12 7 3 3 2 3 9 13 2 3 3 13 2
24 9 2 15 9 13 1 9 0 9 2 13 0 9 2 16 3 0 9 0 9 13 10 9 2
37 9 3 13 13 11 1 11 2 16 13 1 3 0 0 2 0 2 0 7 0 9 2 7 7 10 9 13 3 0 16 10 2 15 13 9 11 2
24 16 15 14 11 13 1 9 9 2 3 4 15 10 9 13 1 9 12 9 1 12 9 9 2
14 16 11 11 2 11 13 3 2 13 15 1 3 0 2
8 3 1 12 9 9 2 2 2
13 10 9 3 15 13 7 7 13 1 0 9 4 2
27 0 9 15 7 1 10 9 9 13 7 3 3 0 13 2 13 2 14 15 3 1 9 7 9 1 9 2
7 13 15 1 9 0 9 2
28 1 9 1 9 7 1 0 9 0 3 0 9 12 0 9 15 3 0 9 1 9 3 3 13 0 0 9 2
13 1 10 9 0 11 13 10 9 0 0 9 11 2
8 13 15 15 3 16 0 9 2
11 3 0 9 4 13 3 3 3 3 13 2
17 16 7 13 0 0 9 1 12 2 9 2 13 15 10 9 0 2
12 0 9 1 9 9 1 11 15 7 13 3 2
18 3 15 13 0 9 1 11 9 2 1 15 13 3 0 7 3 13 2
4 9 9 13 11
2 11 2
20 1 12 9 0 9 1 0 11 4 13 9 0 2 15 15 3 13 3 13 2
13 13 15 11 11 2 9 9 9 9 0 9 9 2
24 1 10 9 13 0 9 3 1 9 0 11 2 3 4 0 9 13 1 12 9 9 7 9 2
21 1 0 9 13 3 9 12 9 2 3 0 9 9 13 14 12 9 1 9 0 2
12 9 13 3 1 9 9 7 13 15 3 9 2
24 1 10 9 13 0 13 1 15 0 9 2 7 0 9 7 0 9 13 1 10 9 0 9 2
30 9 9 7 13 9 1 9 3 12 9 9 2 3 12 9 9 2 1 0 9 2 16 4 15 13 3 15 0 9 2
39 1 9 3 1 12 9 2 3 1 12 9 15 9 13 7 3 15 1 0 9 9 13 3 0 9 2 3 13 15 9 7 13 1 9 9 1 0 9 2
14 9 0 9 1 9 1 15 13 10 14 12 0 9 2
31 1 9 0 11 15 0 9 1 0 9 11 13 13 10 9 7 9 1 0 9 0 9 0 9 2 15 13 7 3 0 2
5 1 11 13 9 9
2 11 2
19 9 9 0 9 1 0 0 0 9 1 11 13 9 0 0 9 0 9 2
25 1 9 2 15 13 9 3 16 0 9 2 13 12 9 9 2 1 13 12 7 12 15 9 13 2
40 9 11 11 1 0 9 13 9 1 9 9 0 9 1 0 9 9 7 13 2 16 1 0 9 9 0 9 13 13 9 9 3 0 7 0 7 13 15 0 2
15 13 1 10 9 7 9 2 7 1 9 9 2 13 11 2
15 0 0 9 2 9 9 11 11 15 3 9 0 9 13 2
15 10 9 4 3 13 0 0 9 1 9 0 9 1 11 2
27 11 13 1 0 9 9 9 9 9 9 7 13 3 9 2 16 9 0 0 9 13 0 0 9 10 9 2
31 1 9 0 1 9 3 0 9 13 0 0 9 0 1 0 9 2 15 1 0 13 1 9 7 9 9 1 9 10 9 2
32 0 0 9 1 10 9 13 2 16 1 9 9 13 9 2 9 7 9 1 0 9 3 0 7 1 10 9 13 13 7 9 2
9 9 0 9 13 1 11 7 1 11
2 11 2
18 9 1 9 2 0 9 7 9 2 4 3 13 1 0 7 0 9 2
12 13 15 3 1 9 1 0 7 0 0 9 2
30 0 9 13 1 9 0 11 7 11 2 0 9 4 13 1 11 2 11 2 11 2 11 2 11 2 11 7 0 11 2
8 0 9 0 9 11 13 1 11
2 11 2
22 0 9 0 0 9 2 0 0 0 0 0 9 1 9 0 11 2 13 3 1 11 2
38 3 12 9 0 9 15 13 1 9 12 0 9 2 15 1 11 13 1 0 9 2 7 1 0 12 9 0 9 11 1 11 2 15 13 3 3 13 2
11 0 12 0 9 13 1 11 12 2 9 2
18 0 9 9 11 13 13 9 0 9 2 15 3 13 12 0 0 9 2
32 11 13 3 3 0 2 7 13 7 9 2 16 1 0 9 1 10 9 0 11 4 13 4 13 7 0 11 2 11 7 11 2
48 0 0 9 0 9 11 13 2 16 11 15 4 13 13 15 9 1 12 9 2 7 1 0 9 15 13 2 16 9 7 9 0 9 13 0 9 4 13 13 10 9 1 9 1 9 0 9 2
6 11 2 9 1 9 13
2 11 2
21 0 9 11 11 3 13 9 1 9 2 10 0 9 9 13 9 1 11 7 11 2
6 9 3 13 1 9 2
37 9 1 0 13 2 16 10 9 11 2 15 1 12 9 13 1 0 9 2 7 13 9 10 9 2 4 13 1 9 7 4 13 13 9 1 9 2
22 9 9 3 13 3 10 9 2 15 13 9 0 11 1 9 12 2 7 10 0 9 2
28 11 2 15 13 1 9 1 12 2 7 12 2 9 7 13 3 12 1 12 9 9 2 13 7 1 9 13 2
17 9 11 1 0 9 1 9 11 13 2 16 9 13 0 0 9 2
21 11 13 1 9 2 16 13 9 0 0 9 7 16 12 9 0 11 13 9 9 2
11 11 1 9 9 1 10 9 13 3 3 2
19 9 11 15 13 1 0 7 13 0 9 1 9 9 2 9 7 0 9 2
12 0 9 13 13 9 9 0 0 9 1 11 2
38 9 11 7 9 11 2 1 15 15 11 13 1 9 1 9 2 13 1 9 2 16 9 13 3 1 9 1 9 9 0 9 2 13 7 13 0 9 2
21 13 1 15 10 9 2 1 15 0 9 13 3 0 0 9 0 9 2 9 2 2
15 9 2 15 13 2 13 14 0 7 1 9 9 15 13 2
8 11 13 10 9 0 9 0 9
24 11 13 0 0 9 0 9 3 2 16 9 11 13 9 2 16 15 11 13 13 12 0 9 2
6 13 15 3 9 11 2
38 0 9 9 11 11 3 13 2 16 0 9 13 13 1 9 9 2 16 11 4 13 9 1 9 1 9 1 0 9 0 3 2 9 0 9 0 9 2
7 0 9 0 9 13 1 9
1 9
7 0 9 0 9 13 1 9
14 0 9 1 9 11 7 11 15 13 3 7 1 9 2
48 16 0 9 3 13 15 2 16 4 10 0 9 0 9 13 13 0 9 2 9 7 12 1 9 9 2 0 9 0 3 0 0 9 2 15 13 2 16 4 11 13 3 3 13 16 0 9 2
37 9 3 3 13 9 11 7 11 2 1 0 9 7 7 15 13 1 9 3 0 7 0 9 0 9 2 16 3 13 1 0 9 11 9 0 9 2
29 10 9 0 9 9 2 1 15 4 13 13 15 12 9 2 3 11 2 11 7 9 2 0 9 2 15 3 13 2
20 3 0 9 13 13 10 9 7 13 13 2 16 11 7 11 13 3 3 13 2
14 9 1 15 3 13 13 2 16 1 10 9 13 9 2
29 7 3 1 9 0 2 15 15 7 0 13 2 13 0 11 7 11 2 16 15 1 15 13 1 9 12 0 9 2
30 13 2 14 1 9 2 16 3 3 13 1 12 9 0 9 2 3 1 15 13 2 16 14 10 9 13 10 9 13 2
32 9 15 13 3 13 2 16 1 15 4 13 2 16 15 7 13 1 9 10 9 13 15 0 9 2 4 15 13 3 10 9 2
16 11 7 11 3 13 13 2 16 15 15 15 13 2 7 3 2
16 0 9 3 4 2 13 15 2 3 13 0 9 10 0 9 2
7 0 9 3 1 15 13 2
35 7 4 13 1 9 11 2 7 3 15 13 1 9 1 9 2 7 15 13 1 9 2 7 15 3 13 9 1 9 9 1 0 9 9 2
11 0 9 1 10 0 9 13 16 13 3 2
9 9 1 11 13 13 3 3 3 2
7 11 13 0 2 7 13 9
32 11 11 13 0 9 9 9 11 7 9 0 9 1 0 9 2 1 15 15 1 0 9 0 9 13 0 9 0 1 0 9 2
19 1 0 9 15 13 1 11 1 11 9 0 2 7 0 9 1 0 9 2
8 1 10 9 15 13 0 9 2
5 13 11 0 9 2
7 11 15 13 0 9 13 2
19 9 7 13 2 1 10 9 13 3 0 2 16 4 15 0 9 3 13 2
15 1 10 9 4 1 15 13 0 13 3 16 12 9 9 2
13 1 0 9 13 9 1 0 7 0 9 9 9 2
18 13 3 7 7 0 9 2 7 15 2 16 11 13 9 1 9 13 2
20 3 13 9 15 2 16 7 13 9 1 0 9 2 15 15 13 1 10 9 2
21 15 13 9 0 9 9 0 9 2 7 7 1 10 9 13 11 13 1 0 9 2
34 1 15 2 15 4 13 2 13 0 2 16 16 4 15 13 13 0 9 2 13 4 13 0 9 9 2 16 4 15 0 9 13 9 2
20 13 4 0 13 3 0 9 0 9 2 9 1 9 0 9 2 15 3 13 2
13 3 13 3 13 2 16 9 9 0 9 11 13 2
8 3 9 3 13 9 9 12 2
11 0 9 15 9 9 12 3 0 9 13 2
11 1 9 10 9 4 7 13 0 9 9 2
17 1 9 10 9 4 3 13 9 1 9 12 9 9 2 15 13 2
8 13 0 13 9 10 9 11 2
19 1 0 9 13 0 13 0 9 9 2 7 3 3 13 9 10 9 13 2
29 1 15 13 3 7 9 9 1 9 0 1 9 2 1 15 13 16 9 7 0 9 2 7 9 1 10 0 9 2
10 7 1 15 15 15 1 11 13 13 2
8 3 0 9 13 7 0 9 2
24 11 15 13 13 3 0 9 9 2 7 7 13 9 15 13 2 3 4 1 9 13 10 9 2
16 1 11 13 1 0 9 0 9 7 11 13 1 15 0 9 2
10 0 9 13 9 1 0 9 0 11 2
6 15 13 3 0 9 2
53 1 9 13 0 9 1 0 9 9 9 2 15 13 3 0 9 7 1 9 4 13 1 9 2 1 15 15 10 9 13 2 16 1 10 9 4 11 13 7 0 9 2 7 0 9 2 7 13 4 9 0 9 2
31 3 15 13 1 15 2 16 4 10 9 4 11 13 14 9 10 0 9 2 7 16 4 15 13 0 3 0 7 0 9 2
12 13 15 2 16 4 13 0 9 7 1 11 2
16 14 2 9 2 15 4 1 11 13 2 15 1 0 9 13 2
9 13 7 9 1 9 0 9 11 2
15 0 9 3 0 9 13 0 9 11 7 9 1 9 11 2
16 9 0 9 0 15 11 13 9 2 15 13 15 9 0 9 2
5 13 14 1 15 2
30 9 13 9 1 0 0 9 2 16 3 4 13 0 9 1 11 2 3 15 13 13 11 2 11 2 7 7 0 9 2
13 3 3 3 13 2 3 13 1 0 9 10 9 2
9 11 7 11 3 13 9 1 0 9
2 11 2
27 11 7 9 1 9 11 13 0 9 1 0 9 1 9 13 1 0 9 12 9 0 0 2 0 0 9 2
7 13 15 3 0 9 11 2
46 0 0 9 11 13 10 9 1 9 0 9 1 11 2 1 15 15 0 9 13 1 9 0 9 2 10 9 15 3 1 0 9 1 9 0 9 13 0 9 1 11 7 0 9 13 2
17 9 13 9 3 7 1 9 11 11 7 9 0 9 11 11 11 2
16 0 9 1 9 9 13 2 16 0 0 9 11 11 15 13 2
8 13 7 2 15 15 15 13 2
42 0 2 0 9 15 13 1 0 9 1 0 9 1 0 9 0 9 1 0 9 11 7 1 9 11 7 1 9 0 11 2 1 15 15 13 9 3 9 2 3 9 2
6 0 9 13 11 10 9
2 11 2
18 9 0 9 0 9 3 13 2 16 13 1 11 12 9 1 9 9 2
6 13 15 3 9 9 2
34 13 13 2 15 1 12 9 13 9 0 9 11 11 11 2 11 1 9 1 9 0 2 0 9 2 1 10 9 15 3 13 9 9 2
9 1 0 9 1 11 12 9 13 3
2 11 2
15 3 0 9 13 3 0 7 0 9 1 0 9 1 11 2
46 1 0 9 15 0 9 13 13 10 0 9 1 11 2 16 0 9 13 2 16 13 3 15 9 1 9 2 0 9 1 15 2 7 16 10 9 13 13 3 14 12 9 1 10 9 2
29 0 9 0 0 9 3 13 0 9 0 9 11 0 11 2 1 15 1 9 11 13 3 12 9 0 1 11 9 2
20 13 3 2 16 15 3 3 13 13 0 9 2 15 13 1 9 11 2 11 2
27 3 3 1 12 9 13 4 13 9 1 9 7 9 7 1 12 9 4 14 13 9 2 15 13 11 9 2
16 0 9 7 13 2 16 9 3 13 2 13 7 13 0 9 2
26 9 1 11 7 10 0 9 11 13 3 1 9 3 2 16 0 9 13 11 1 9 9 1 0 9 2
20 1 10 9 13 3 1 9 11 7 1 0 9 2 16 10 9 13 0 9 2
27 0 9 15 13 1 9 1 0 0 9 11 1 9 10 9 2 15 13 1 0 9 1 0 9 7 0 9
22 1 10 9 11 1 9 7 1 9 1 9 15 13 11 11 1 1 11 2 9 9 11
6 9 0 0 9 13 13
2 11 2
19 9 9 0 9 1 0 0 0 9 1 11 13 9 0 0 9 0 9 2
40 9 11 11 1 0 9 13 9 1 9 9 0 9 1 0 9 9 7 13 2 16 1 0 9 9 0 9 13 13 9 9 3 0 7 0 7 13 15 0 2
6 11 13 0 9 0 9
2 11 2
24 0 9 9 11 11 13 2 16 3 1 9 10 9 4 15 11 13 13 1 9 10 0 9 2
19 1 9 1 9 11 13 2 16 2 3 15 15 13 7 15 4 13 2 2
29 1 0 9 13 2 16 1 10 9 2 4 15 13 11 13 0 9 1 9 2 3 15 3 13 0 12 9 2 2
19 1 0 9 4 1 11 13 2 3 0 13 15 1 9 1 0 9 2 2
11 9 9 0 9 1 11 13 2 0 2 9
2 11 2
26 9 9 0 9 1 11 11 11 11 13 1 9 9 1 0 9 2 0 2 0 9 1 9 0 9 2
37 2 16 4 1 15 13 1 15 2 16 4 13 0 9 13 2 13 15 2 16 13 9 9 7 13 15 2 2 13 15 9 9 0 9 11 11 2
11 10 9 13 10 9 9 1 9 11 11 2
21 2 3 1 0 9 13 3 14 9 2 13 9 7 15 15 15 1 9 13 2 2
22 16 11 11 13 0 9 3 2 13 11 11 1 9 0 9 2 1 15 0 9 13 2
33 9 1 0 9 13 2 13 2 16 9 1 0 9 1 9 13 2 0 9 1 9 11 2 10 9 3 13 2 13 3 1 9 2
15 15 2 16 13 2 0 2 9 2 14 13 1 10 9 2
12 11 11 3 13 9 0 9 1 0 0 9 2
8 0 9 15 1 9 14 13 2
14 2 15 13 0 2 9 15 3 2 13 2 9 2 2
9 1 11 3 3 13 9 0 9 2
7 0 9 9 15 13 9 2
21 3 7 1 0 2 0 9 2 15 13 3 10 9 13 2 2 0 2 9 13 2
18 9 11 11 1 0 11 13 1 9 2 0 2 9 9 12 12 9 2
12 9 1 11 1 11 13 1 0 9 1 9 2
12 2 15 9 0 9 13 3 2 1 12 9 2
15 9 4 15 7 0 9 1 9 7 13 13 15 1 9 2
8 0 11 15 13 1 12 9 2
7 3 13 1 15 3 3 2
11 0 9 13 14 12 2 2 13 11 11 2
24 2 15 13 9 0 1 11 2 2 13 15 1 15 11 11 2 16 15 1 15 13 13 9 2
22 1 9 2 16 15 13 13 0 9 2 15 13 2 16 14 2 16 13 1 15 9 2
8 9 15 13 2 16 13 12 9
7 11 2 11 2 11 2 2
20 9 9 1 11 2 11 13 1 9 3 9 1 0 0 9 1 9 10 9 2
15 11 2 11 2 2 12 2 13 13 1 9 3 12 9 2
28 9 13 1 10 9 1 0 9 1 9 1 9 1 9 9 0 9 2 10 9 13 9 1 0 9 9 9 2
17 1 10 9 13 0 1 10 9 12 9 7 9 13 1 0 9 2
19 3 1 9 0 9 9 13 1 0 9 1 11 9 0 1 10 0 9 2
13 9 13 1 3 0 12 0 11 2 11 2 9 2
19 1 12 9 15 13 1 15 2 16 13 13 0 9 9 7 0 0 9 2
26 3 15 3 13 9 2 15 15 9 13 2 12 9 13 3 0 9 2 15 13 1 3 0 9 0 2
9 10 9 13 9 7 0 0 9 2
7 1 9 13 9 9 9 2
9 1 9 13 1 11 12 11 0 2
9 9 13 1 9 2 0 1 9 2
23 9 3 13 0 9 9 9 2 10 9 4 0 0 9 13 1 10 9 1 11 2 11 2
4 9 1 9 13
5 11 2 11 2 2
14 1 9 15 13 12 7 9 9 9 0 9 1 11 2
5 3 1 9 13 2
17 1 9 1 12 9 1 9 15 1 11 2 0 9 13 0 9 2
17 1 9 0 15 9 13 1 9 2 13 1 15 7 3 15 13 2
3 9 13 9
5 11 2 11 2 2
14 1 9 0 9 9 13 0 0 9 1 11 1 11 2
18 1 0 0 9 9 13 1 9 13 9 1 3 16 12 9 12 9 2
14 13 3 0 9 2 9 7 13 9 1 10 0 9 2
12 9 13 1 0 9 1 9 1 9 1 9 2
6 1 9 13 1 9 9
5 11 2 11 2 2
21 12 3 0 9 1 9 12 7 12 9 1 11 13 3 1 9 0 9 1 9 2
15 12 0 9 13 13 9 1 12 9 7 9 9 11 11 2
7 13 0 7 1 0 9 2
8 13 9 14 1 9 9 9 2
16 9 1 15 13 3 9 1 9 2 15 13 1 10 0 9 2
4 1 9 7 9
2 11 11
44 9 11 11 2 9 2 9 0 9 2 7 10 9 9 11 11 2 9 9 2 3 7 3 13 12 1 0 9 0 9 0 9 1 9 2 7 9 1 0 9 2 7 3 2
33 9 0 9 13 1 15 1 9 12 2 15 13 9 9 2 9 2 0 9 7 9 1 10 9 2 15 2 15 13 0 0 9 2
28 9 12 13 9 2 15 4 9 13 0 9 2 9 0 9 2 1 15 9 2 9 2 9 2 9 7 9 2
7 9 12 13 9 0 9 2
48 9 11 2 15 15 9 0 9 3 13 2 13 1 9 15 0 9 2 1 9 1 10 9 7 9 2 15 9 9 2 9 2 0 9 2 0 9 3 16 9 2 0 9 3 16 0 9 2
11 15 12 9 15 3 3 13 7 13 15 2
15 9 12 13 1 9 12 1 0 9 2 3 3 1 9 2
57 10 9 7 9 13 14 3 1 9 9 2 7 1 0 9 9 1 12 0 9 2 16 9 12 9 7 9 2 3 0 9 13 2 15 1 15 13 13 9 9 12 10 9 2 3 9 7 15 0 9 1 9 2 9 2 9 2
15 16 4 9 1 9 13 2 13 4 9 2 15 13 3 2
28 13 1 15 2 16 15 2 15 15 13 9 9 7 9 2 13 9 9 7 13 15 3 2 3 3 7 3 2
23 3 10 9 12 1 9 13 7 13 2 15 13 1 0 9 12 1 9 12 7 9 12 2
32 3 15 13 13 2 16 3 1 9 2 7 3 15 3 3 1 9 3 9 12 2 7 9 12 2 15 13 9 2 15 13 2
6 13 1 9 3 12 2
11 1 0 13 0 9 2 1 0 11 11 2
25 10 9 12 15 13 9 9 2 16 13 0 13 0 9 2 15 4 15 1 0 9 13 15 0 2
32 13 2 16 13 1 15 3 16 9 0 9 12 2 15 15 1 15 13 2 7 13 15 13 2 1 15 13 2 3 1 9 2
18 0 9 1 9 13 2 16 15 13 9 0 9 2 15 15 3 13 2
25 1 15 13 3 10 9 2 16 13 13 0 2 16 15 1 15 13 2 7 0 2 16 15 13 2
7 16 9 10 9 1 9 2
32 13 15 1 9 2 3 15 13 9 9 2 3 13 1 9 2 16 4 13 2 16 13 9 1 9 2 13 7 13 3 3 2
29 16 13 9 1 10 9 9 0 9 2 0 0 2 3 0 9 0 9 2 3 13 3 1 9 7 13 15 9 2
13 13 15 3 3 2 16 13 3 0 2 3 0 2
27 16 4 13 0 3 2 13 4 15 9 2 10 9 13 13 0 14 1 0 9 2 16 15 13 9 9 2
31 15 2 15 13 1 9 2 15 13 1 9 9 2 13 15 15 13 2 1 0 9 13 13 7 9 2 7 9 7 3 2
39 16 3 13 13 9 0 9 2 1 15 2 7 2 16 15 2 2 13 13 7 9 0 9 2 1 15 2 2 13 2 14 15 1 15 1 3 0 9 2
45 10 9 12 13 2 16 4 15 15 3 13 2 16 15 13 1 9 13 16 1 0 9 2 15 15 13 13 2 13 2 16 4 13 2 15 13 2 7 7 15 3 14 15 13 2
23 7 15 13 13 2 16 9 13 3 1 9 2 15 13 3 3 3 0 2 7 3 0 2
31 9 12 2 15 15 0 9 13 3 2 13 1 0 3 2 16 15 9 1 0 9 10 9 13 3 2 7 16 3 3 2
42 16 15 3 13 2 16 9 13 2 13 1 15 13 10 0 9 2 15 4 15 9 2 13 9 0 2 0 7 0 9 2 3 13 2 16 4 15 15 13 1 15 2
19 9 4 13 13 9 2 3 4 15 1 10 9 3 10 0 9 3 13 2
3 7 3 2
17 16 4 13 2 16 9 2 13 4 1 15 0 7 0 11 9 2
35 13 15 2 16 4 13 0 9 15 2 3 3 13 2 16 13 7 3 2 3 3 13 2 7 16 15 0 13 2 16 4 3 13 13 2
22 16 3 13 15 2 16 3 13 2 13 13 2 16 0 9 13 12 1 0 9 3 2
15 9 10 9 13 0 9 2 0 9 7 9 13 0 9 2
10 1 0 9 9 3 13 0 7 0 2
23 9 12 9 9 7 9 3 13 1 15 2 16 4 15 10 9 12 3 13 1 15 0 2
32 9 13 2 16 13 7 13 0 9 1 9 7 9 2 3 13 3 0 2 16 13 0 2 13 15 0 7 1 9 1 9 2
16 3 4 3 13 0 2 16 4 10 9 13 3 2 3 13 2
31 1 10 9 15 15 13 13 2 16 4 0 9 13 1 9 9 0 2 3 3 2 16 4 1 10 9 3 13 10 9 2
28 1 0 9 10 9 12 3 13 2 16 13 1 0 9 2 16 9 2 1 15 13 9 9 2 13 9 9 2
23 0 13 2 16 4 15 3 13 0 7 13 10 0 9 3 2 16 4 10 9 0 13 2
18 3 16 15 10 0 0 9 13 2 16 13 3 0 9 9 9 9 2
27 16 15 7 10 9 12 13 9 12 1 9 0 9 0 9 2 13 2 16 4 13 13 1 0 0 9 2
25 16 4 13 1 9 3 0 2 3 4 13 15 13 7 13 2 1 9 2 16 13 0 7 0 2
13 7 14 16 13 3 0 9 10 0 9 0 9 2
13 9 9 7 0 0 9 13 9 9 1 9 9 2
13 9 0 0 9 9 13 9 0 9 9 9 9 2
10 0 9 13 0 9 1 9 12 9 2
18 9 0 9 7 10 9 2 1 15 13 10 9 2 13 0 9 9 2
6 0 13 0 2 2 2
33 9 0 9 13 3 9 9 9 1 0 9 0 15 7 9 0 9 2 1 0 9 7 9 10 9 2 15 13 13 0 3 9 2
20 15 13 2 16 9 13 3 0 2 7 16 15 13 13 2 14 1 0 9 2
10 1 0 9 9 7 9 13 0 9 2
21 3 16 13 15 12 1 9 2 3 13 0 9 3 3 13 9 9 0 9 9 2
17 7 14 16 15 3 13 0 9 9 0 3 0 9 10 0 9 2
24 13 3 3 3 0 9 9 0 9 2 13 3 0 9 0 9 2 1 15 0 9 9 13 2
43 7 15 10 3 0 9 9 1 9 7 9 1 9 2 7 3 2 1 15 2 3 15 13 9 7 0 9 2 1 9 1 9 7 9 0 9 2 15 15 13 13 9 2
25 14 16 4 13 9 1 0 0 7 0 9 2 15 4 15 15 13 3 2 16 13 9 9 9 2
46 1 10 9 13 2 13 7 13 0 9 0 9 3 0 2 1 9 1 0 9 2 1 15 2 16 15 15 13 7 13 2 1 9 1 9 2 15 3 13 7 15 15 7 10 9 2
9 13 9 9 2 10 9 13 3 2
27 7 13 1 9 9 0 9 3 0 2 15 1 9 12 15 13 1 0 9 12 7 15 15 3 3 13 2
23 7 15 1 9 0 9 12 13 1 9 12 13 2 7 15 3 13 3 2 3 1 9 2
30 13 3 0 9 2 16 9 13 12 1 9 10 9 2 16 13 2 16 13 2 0 9 2 15 13 0 9 9 0 2
54 7 15 3 13 16 9 10 0 9 2 15 15 13 1 9 0 9 9 9 7 13 1 10 9 1 12 9 2 16 3 13 2 16 15 15 13 9 2 7 16 4 15 9 13 2 13 2 16 15 1 15 15 13 2
31 10 9 12 3 13 2 16 15 1 15 10 13 1 9 0 2 0 2 7 0 0 9 2 7 4 1 9 7 9 13 2
15 13 2 16 4 10 9 1 15 13 9 2 7 3 3 2
13 3 4 15 13 7 13 4 1 15 1 15 9 2
9 7 1 15 0 13 3 11 11 2
6 13 15 15 2 13 2
25 13 1 9 9 1 0 9 1 9 7 13 15 2 15 13 9 2 13 15 1 9 9 2 2 2
18 16 1 15 13 2 13 2 2 3 2 3 13 2 13 0 9 2 2
22 7 16 15 13 2 13 2 2 3 2 3 13 2 13 9 1 11 3 1 9 2 2
48 12 9 0 0 9 9 2 9 9 2 0 11 2 9 11 2 11 11 2 9 2 1 15 15 13 2 16 13 0 9 2 11 2 11 2 11 2 9 0 2 9 2 9 2 9 2 2 2
25 0 0 9 2 15 4 13 13 1 9 7 13 9 1 9 2 2 13 15 1 15 2 2 2 2
14 3 1 9 0 2 0 9 1 10 9 13 10 9 2
6 13 15 9 10 9 2
15 15 13 9 1 9 9 9 9 1 9 0 9 9 12 2
8 13 2 14 2 3 15 13 2
7 13 13 10 9 0 9 2
10 7 13 14 1 0 9 9 0 9 2
16 13 2 16 4 15 1 15 9 1 0 0 9 15 3 13 2
30 13 15 13 9 2 3 4 15 13 13 2 16 9 9 9 13 0 9 2 7 13 3 0 2 16 9 13 10 9 2
14 13 2 14 15 2 13 4 15 2 16 4 15 13 2
11 9 9 9 1 0 0 9 4 13 0 2
11 9 9 9 13 9 7 15 2 15 13 2
24 7 0 13 14 1 9 2 1 15 13 0 7 0 2 1 9 2 16 15 15 13 15 13 2
7 13 15 10 9 9 13 2
2 13 2
2 3 2
5 3 7 1 15 2
5 13 9 0 9 2
3 13 9 2
9 10 9 9 13 3 14 0 9 2
10 13 2 14 15 2 13 1 9 15 2
7 13 15 3 7 3 13 2
5 13 15 0 9 2
13 13 2 14 15 2 3 1 9 14 13 15 3 2
3 12 2 12
3 0 9 9
17 1 0 0 9 1 9 10 0 9 2 9 2 15 3 3 13 2
15 16 0 9 15 13 9 2 9 9 2 0 1 0 9 2
9 7 13 15 9 2 15 15 13 2
13 1 9 10 9 15 13 13 0 0 9 0 9 2
24 9 9 2 15 13 9 1 0 9 2 13 13 3 0 2 7 3 14 14 13 15 1 9 2
18 7 13 1 0 9 2 0 9 2 7 2 0 9 2 14 13 0 2
13 1 9 9 15 7 1 0 9 13 12 0 9 2
12 13 1 15 11 1 12 2 9 10 2 9 2
30 9 3 0 0 9 1 0 9 2 3 0 9 0 9 1 0 9 2 1 10 9 3 13 0 9 12 0 0 9 2
16 13 15 2 16 9 13 9 10 9 1 9 1 12 9 9 2
33 0 9 2 0 9 1 9 11 11 13 9 1 12 0 9 2 3 15 13 1 9 9 2 15 2 13 0 9 16 0 9 2 2
25 9 13 2 16 9 13 14 9 10 9 1 10 0 9 2 7 16 13 3 9 9 1 10 9 2
9 1 10 9 13 1 0 9 9 2
14 13 1 9 2 3 1 9 2 16 4 10 9 13 2
21 10 9 2 3 2 0 11 2 13 1 9 2 16 4 9 13 1 10 0 9 2
5 15 15 13 9 2
34 7 2 7 1 15 15 1 0 9 13 2 0 9 0 9 2 1 15 13 9 1 9 9 0 9 2 13 3 9 1 9 0 9 2
18 0 9 13 3 0 2 7 3 9 1 15 7 0 9 13 3 0 2
38 0 9 1 9 1 9 2 12 13 14 9 1 9 0 9 2 7 3 1 0 9 0 9 2 3 9 1 9 10 0 9 16 9 13 3 1 9 2
18 9 1 9 10 0 9 2 16 13 9 11 2 4 13 3 3 2 2
26 3 10 9 15 13 2 15 13 14 1 15 2 7 3 1 11 2 2 13 15 13 1 9 0 9 2
46 13 2 16 1 15 4 13 9 2 9 2 9 1 9 2 13 0 9 3 1 10 9 1 9 7 9 2 7 2 16 1 15 13 1 9 2 16 13 1 15 1 10 0 9 3 2
4 9 2 11 11
3 12 2 12
47 2 2 2 1 9 9 11 2 11 2 0 7 0 9 2 2 9 12 2 12 2 12 2 12 2 15 3 1 9 3 3 13 9 2 3 13 1 9 2 2 2 2 0 2 2 2 2
16 13 15 12 1 0 9 9 9 2 1 15 3 1 15 13 2
3 2 2 2
43 13 3 1 9 11 2 15 1 9 15 9 10 0 9 3 13 7 13 2 2 3 13 13 2 16 15 11 13 2 16 4 3 13 2 16 2 13 1 9 11 2 2 2
10 10 0 9 13 1 10 0 9 9 2
9 2 1 9 13 1 9 9 2 2
10 2 1 0 9 13 1 9 9 2 2
6 3 15 10 9 13 2
30 13 9 3 0 2 13 1 15 3 15 2 13 15 1 15 10 9 0 0 7 15 15 1 0 9 9 13 3 13 2
22 3 4 3 13 13 9 3 9 2 16 4 14 3 2 7 7 3 13 3 1 9 2
5 9 2 11 2 11
10 10 9 15 13 1 0 9 10 9 2
1 9
2 9 9
2 11 11
8 9 9 15 13 3 1 9 2
5 3 13 9 0 2
18 9 13 13 0 9 2 15 15 13 2 16 15 13 2 3 13 9 2
18 13 0 7 3 0 2 16 15 1 9 13 13 9 1 0 1 0 2
19 4 3 13 2 16 0 9 3 13 2 13 2 14 1 10 9 0 9 2
9 7 15 15 9 9 13 1 9 2
9 9 7 1 9 13 7 0 9 2
25 7 3 0 2 7 0 2 13 13 2 16 16 9 13 7 13 1 9 2 7 15 1 15 13 2
15 3 15 13 9 2 7 13 7 13 2 16 13 15 3 2
9 10 7 0 9 4 15 3 13 2
9 13 3 3 0 9 2 0 9 2
6 7 13 15 3 3 2
20 13 9 2 16 15 13 9 9 7 9 1 9 2 1 15 15 13 13 9 2
12 0 13 15 3 1 9 2 1 15 3 13 2
18 9 9 15 13 2 16 4 13 2 16 12 9 13 13 0 9 9 2
15 13 7 3 1 0 9 0 9 2 0 9 7 0 9 2
32 3 0 13 15 1 15 2 15 13 3 0 9 1 10 9 2 7 13 15 2 16 0 0 9 13 13 14 1 2 9 2 2
14 1 10 9 15 9 13 13 9 7 13 13 1 9 2
30 2 0 9 4 1 0 9 13 1 12 0 9 2 9 7 9 2 7 12 13 0 2 2 13 11 11 2 0 9 2
10 14 2 3 0 9 4 3 13 9 2
18 3 15 3 13 1 9 2 16 9 13 13 3 1 9 9 7 9 2
39 7 9 0 9 1 10 9 13 1 0 9 1 3 0 9 9 2 7 1 0 0 2 0 9 9 15 13 0 9 2 9 7 9 2 3 0 1 0 2
16 3 15 1 9 0 1 0 0 9 13 1 10 0 9 0 2
22 7 13 9 0 3 1 0 9 7 0 9 2 15 13 13 1 9 0 7 0 9 2
37 9 2 12 13 11 11 1 11 2 2 0 9 2 15 15 13 3 13 9 9 2 16 15 1 15 13 9 2 15 3 13 13 3 0 9 9 2
29 13 13 2 16 1 9 13 3 3 16 1 9 2 1 9 3 16 1 9 2 1 9 3 16 1 9 2 2 2
24 3 13 13 2 16 1 0 9 9 15 1 0 9 13 15 2 15 13 13 1 0 9 2 2
8 13 7 3 1 9 10 9 2
12 2 13 2 16 9 0 9 15 13 1 9 2
30 7 0 9 10 9 13 2 16 9 9 13 3 13 1 9 10 9 9 7 9 2 2 13 11 2 11 9 2 12 2
15 11 2 11 7 9 2 2 9 9 2 9 7 9 1 9
39 9 2 9 2 11 2 11 2 9 2 2 1 0 9 0 1 11 13 1 9 12 3 0 9 2 0 1 0 9 9 12 0 0 9 1 10 0 9 2
15 3 12 9 13 1 0 9 0 12 9 1 0 0 9 2
22 1 9 7 1 9 9 0 9 11 15 7 13 13 9 2 15 13 1 10 9 9 2
44 1 0 9 15 13 1 9 0 9 2 3 9 2 9 2 9 7 9 2 3 15 13 9 10 9 1 0 9 2 1 0 9 7 0 9 14 1 9 0 7 3 0 9 2
56 3 15 3 9 13 9 10 0 9 1 9 1 9 2 0 9 7 0 9 2 13 15 1 9 1 9 2 1 0 9 0 9 1 0 9 7 10 9 7 12 9 9 4 13 7 9 9 0 9 1 0 9 1 9 9 2
28 0 9 13 9 1 9 2 9 7 9 7 3 3 13 0 9 2 0 0 2 0 7 0 9 0 0 9 2
12 9 13 9 1 9 7 0 9 0 0 9 2
88 0 9 15 13 13 3 0 9 2 15 13 1 9 0 2 9 9 1 9 9 1 9 7 9 2 9 9 1 0 0 9 2 9 0 9 9 1 9 2 9 9 1 9 7 1 0 9 2 9 9 9 2 9 2 0 9 2 10 9 1 9 10 7 0 2 0 9 1 9 2 10 9 1 0 0 9 1 9 7 9 14 1 9 9 3 2 2 2
45 9 13 12 9 2 2 0 1 12 9 13 0 9 3 2 3 13 1 3 16 12 9 2 7 4 3 13 14 9 7 9 0 9 2 7 3 9 2 0 7 0 9 7 9 2
38 13 4 15 13 0 9 9 2 15 13 1 9 7 9 2 10 0 9 13 9 0 9 0 7 0 9 3 7 3 3 15 2 10 9 13 9 9 2
35 9 1 9 10 9 13 13 2 3 0 9 2 12 9 2 7 0 9 2 12 9 2 1 1 0 9 0 9 3 3 13 9 0 9 2
2 11 11
6 2 13 1 9 9 2
11 1 0 9 4 15 13 3 3 0 9 2
13 3 15 13 1 2 0 2 7 2 0 2 9 2
20 12 1 0 9 9 15 13 1 9 2 3 13 1 9 0 2 2 2 2 2
39 1 9 0 9 13 3 0 2 0 9 3 2 0 9 13 1 5 0 2 0 2 9 7 9 13 2 13 2 13 5 0 2 0 9 1 0 2 0 2
9 3 7 13 1 10 9 3 3 2
27 1 9 1 9 0 11 4 3 13 12 9 0 10 7 0 9 2 7 13 3 0 1 0 9 0 9 2
12 13 13 9 7 3 13 10 0 9 7 9 2
62 9 10 9 7 9 13 2 3 13 2 16 15 9 2 15 15 3 13 0 9 2 13 1 12 9 2 0 2 0 0 2 0 9 2 7 0 2 0 0 0 9 2 2 13 9 2 13 2 13 9 2 9 2 2 9 13 2 13 1 9 9 2
40 2 1 0 9 13 1 9 9 9 2 1 0 1 10 9 2 2 9 9 1 10 9 13 1 9 2 16 13 0 2 3 0 7 16 13 1 0 9 9 2
2 7 2
2 12 2
28 1 9 16 13 0 9 2 13 9 2 13 9 2 13 9 2 13 1 9 0 2 9 0 9 13 3 0 2
2 12 2
30 9 0 9 13 3 9 0 2 3 1 9 2 7 13 15 15 3 1 9 0 2 0 9 2 13 1 9 0 9 2
8 13 4 1 0 9 0 9 2
10 9 9 13 1 9 9 9 0 9 2
12 10 9 15 13 9 1 0 9 1 0 9 2
7 3 13 9 0 12 9 2
46 3 15 4 13 9 2 9 13 13 9 1 0 9 9 2 2 7 3 4 3 15 13 13 1 9 1 9 2 13 3 13 13 9 1 10 9 2 2 13 3 1 0 2 0 9 2
2 12 2
34 0 9 13 3 0 2 7 16 9 13 3 9 0 2 13 9 9 3 2 0 3 1 15 2 16 15 1 15 13 9 1 0 9 2
14 2 1 15 9 13 0 9 7 13 0 9 2 2 2
14 2 0 9 2 3 13 0 9 2 13 0 9 2 2
16 10 9 3 13 9 10 9 1 9 2 3 13 1 9 0 2
2 12 2
26 0 9 9 0 9 13 10 9 2 16 2 1 9 1 9 0 2 13 2 16 4 4 13 9 9 2
29 7 3 0 9 2 9 4 13 3 2 13 13 9 9 2 7 0 9 2 2 15 1 9 1 9 13 0 13 2
20 3 13 15 1 9 16 4 13 9 2 9 2 9 2 13 9 2 13 9 2
2 12 2
21 9 0 9 2 0 3 2 0 9 1 0 9 2 2 13 7 10 9 0 9 2
56 7 3 2 9 2 10 9 1 9 0 9 15 13 0 9 2 13 13 9 9 2 9 2 16 9 1 0 9 9 0 2 2 10 9 2 2 7 13 7 9 9 2 0 9 2 9 2 2 15 9 0 9 13 15 13 2
24 16 4 15 13 3 13 2 13 2 16 15 0 3 2 0 9 13 13 7 13 3 7 3 2
36 7 13 3 0 13 2 16 7 1 0 9 13 3 9 13 15 3 2 7 3 2 1 9 2 15 7 13 1 0 0 9 2 1 9 9 2
21 9 1 12 9 1 9 15 3 13 2 1 9 10 9 13 1 9 0 9 9 2
12 3 9 13 10 9 2 16 2 2 2 2 2
45 9 10 9 13 13 2 16 13 0 9 0 9 13 3 0 2 3 7 0 2 7 13 9 2 16 9 10 9 13 13 1 15 3 0 7 0 2 13 1 3 0 9 0 9 2
36 3 1 10 9 2 3 16 1 0 2 15 7 13 0 13 1 9 2 13 10 0 2 0 2 9 7 0 9 2 1 15 15 15 3 13 2
7 7 1 15 3 3 3 2
1 11
36 9 2 12 11 11 2 11 0 2 9 9 1 11 1 11 2 13 9 10 12 9 2 1 15 4 2 1 10 9 2 13 4 13 0 11 2
41 10 9 4 13 1 0 9 2 0 9 2 15 13 0 11 13 2 2 1 15 15 13 13 2 16 10 9 13 9 1 0 9 2 7 7 1 0 9 1 9 2
66 9 13 9 2 9 2 0 9 2 0 9 7 0 9 1 9 1 0 0 9 2 16 11 2 12 2 11 2 12 2 0 9 2 14 1 3 0 2 16 11 2 11 2 11 2 12 2 11 2 9 11 2 9 2 9 2 2 9 1 11 2 7 0 9 2 2
52 0 9 13 0 14 3 2 16 13 9 15 13 9 0 9 2 15 4 13 4 9 3 13 2 7 2 15 13 0 2 3 2 16 13 9 2 10 9 9 13 3 2 16 4 15 9 13 13 1 10 9 2
27 12 9 2 15 0 9 13 1 9 2 15 13 4 13 1 12 9 2 13 9 0 9 9 0 1 9 2
20 13 15 1 12 5 7 13 3 2 9 16 9 2 0 9 7 0 9 9 2
14 15 3 13 0 9 9 1 0 9 1 0 12 9 2
29 3 2 9 15 13 3 0 2 16 3 13 1 0 9 16 1 0 9 2 16 3 14 9 2 0 9 16 9 2
31 0 9 1 0 9 15 1 9 13 3 1 9 3 1 12 2 0 9 2 3 13 9 9 13 1 9 1 9 3 9 2
44 9 2 12 0 9 1 9 2 11 2 2 0 9 2 10 0 9 13 9 0 7 0 9 2 13 13 0 9 1 9 13 9 9 2 1 15 15 13 9 1 9 7 9 2
12 9 2 12 9 13 9 2 0 0 9 9 2
37 16 4 0 9 13 0 9 1 9 1 9 7 9 2 13 9 9 11 1 0 9 1 12 7 12 9 9 1 12 7 3 1 12 12 9 9 2
26 13 0 9 10 9 15 2 16 15 13 13 9 1 9 2 1 9 7 1 9 1 15 9 1 0 2
28 3 9 1 0 9 1 9 2 12 13 9 9 2 9 7 0 9 13 9 9 1 9 9 7 9 0 9 2
12 1 10 9 4 1 12 9 13 10 9 9 2
35 15 2 15 13 16 9 13 3 9 7 9 2 3 13 2 3 1 9 10 9 2 1 9 13 15 9 7 9 3 0 9 9 7 9 2
21 9 15 3 13 0 9 9 0 7 0 9 1 0 9 7 1 0 3 0 9 2
26 16 10 9 9 13 1 9 13 9 0 1 0 9 2 0 9 15 13 9 0 0 9 1 0 9 2
29 7 0 9 3 13 1 15 2 16 9 4 13 13 9 9 0 9 7 9 0 4 13 13 3 4 13 10 9 2
15 13 1 9 7 9 9 7 9 10 0 9 15 13 0 2
52 3 9 13 1 10 1 9 0 9 2 1 0 9 2 1 9 1 9 2 1 9 2 0 16 13 1 12 9 2 7 0 9 9 7 9 2 15 13 9 10 9 2 13 1 15 0 16 13 3 1 9 2
33 1 10 0 9 2 3 7 1 0 0 9 2 13 3 9 0 9 2 15 13 10 9 1 9 2 16 13 9 0 9 7 9 2
33 9 13 2 16 13 3 0 9 9 2 16 16 13 15 9 3 0 2 13 0 15 3 13 1 0 9 7 13 0 3 13 9 2
10 0 9 4 15 7 13 13 0 9 2
23 1 0 10 9 13 0 0 9 9 0 9 2 3 3 2 7 1 10 9 15 9 13 2
41 7 2 3 15 15 13 13 0 2 13 0 9 2 7 13 1 15 2 3 3 4 13 2 1 0 1 0 9 2 1 0 9 7 1 0 9 13 3 0 9 2
41 3 0 2 0 9 9 1 10 9 13 3 13 2 3 0 0 9 13 0 1 9 0 9 2 1 9 0 7 0 0 9 7 1 9 1 9 1 3 0 9 2
29 9 3 13 4 1 9 13 7 13 4 13 0 9 7 0 9 2 15 15 13 0 2 7 1 0 16 0 9 2
9 15 13 1 9 1 9 0 9 2
22 16 13 0 7 3 0 9 2 13 0 13 2 16 3 0 9 13 15 1 12 9 2
29 1 12 9 13 15 9 7 9 2 15 13 9 2 0 9 7 9 1 0 9 1 10 9 1 0 7 0 9 2
33 10 9 13 13 0 2 13 2 16 1 15 2 16 4 13 15 0 2 13 3 16 4 13 0 13 9 7 13 9 1 0 9 2
30 7 13 4 13 0 3 7 1 9 13 2 3 7 0 9 2 2 3 15 13 1 9 1 9 0 15 1 10 9 2
31 13 1 10 9 15 1 15 4 13 4 13 1 0 2 15 13 2 16 10 9 13 3 0 7 3 16 13 10 9 0 2
28 0 9 13 15 2 15 13 11 2 9 2 15 15 13 0 9 0 9 2 3 3 2 3 0 9 0 9 2
8 3 15 9 9 13 3 0 2
17 12 9 13 9 1 9 7 1 9 13 7 13 15 3 13 9 2
20 3 0 9 7 13 13 15 0 9 10 9 7 13 0 15 13 1 0 9 2
13 13 4 13 9 1 0 9 9 7 9 10 9 2
17 16 9 9 13 0 9 13 3 0 9 10 9 2 0 9 0 2
25 1 12 9 13 9 11 2 11 2 11 2 16 9 1 10 9 4 13 13 0 1 9 0 9 2
61 1 0 9 13 1 3 0 9 13 3 16 13 2 16 0 9 13 12 1 0 9 1 9 2 7 16 13 2 16 9 13 3 13 1 9 0 1 9 0 7 16 13 1 15 0 13 1 9 2 16 9 1 9 13 13 2 7 9 13 0 2
17 10 9 3 16 13 0 9 0 9 2 7 13 3 9 16 9 2
13 15 9 9 13 9 2 9 2 9 7 0 9 2
21 3 4 0 9 13 1 0 16 0 2 15 13 2 16 0 9 9 3 13 0 2
6 7 15 9 0 9 2
27 13 4 0 9 13 2 16 9 13 9 9 9 7 16 3 0 9 13 2 16 9 13 9 1 0 9 2
41 7 3 2 16 9 9 13 1 0 2 9 9 2 15 15 13 13 9 2 7 3 9 2 15 13 1 9 9 0 9 2 7 13 15 9 1 0 0 9 2 2
5 3 15 13 13 2
30 13 13 1 3 0 9 2 16 13 2 16 0 9 15 13 2 16 4 13 9 0 9 2 16 3 13 1 0 9 2
20 16 7 1 0 9 9 0 9 0 7 9 9 1 9 7 9 1 9 13 2
77 7 3 13 3 3 9 2 1 15 13 2 16 15 3 0 9 13 13 2 3 0 9 13 9 1 9 9 2 3 15 10 9 13 1 0 9 3 1 15 0 7 0 9 2 1 9 9 2 1 0 9 9 2 1 9 9 2 7 3 15 13 0 9 2 13 0 1 0 2 15 15 15 13 13 3 0 2
21 9 13 1 15 2 16 1 9 0 9 13 1 3 2 16 13 0 13 0 9 2
9 9 16 0 9 13 4 13 3 2
20 9 2 3 13 1 0 9 7 9 2 13 0 2 13 2 14 13 0 9 2
17 12 1 0 9 2 1 15 13 0 9 13 2 13 10 0 9 2
23 3 2 1 9 10 9 7 9 13 15 3 10 9 2 15 9 13 1 0 9 0 9 2
6 9 13 9 0 9 2
11 13 13 2 16 11 13 3 0 16 11 2
30 13 15 1 9 11 11 2 16 13 3 16 0 2 7 2 13 1 9 9 2 7 13 9 9 0 9 1 0 9 2
26 16 1 12 12 9 4 3 13 3 9 0 9 2 3 3 12 12 9 13 1 9 0 9 0 3 2
16 14 13 2 10 9 1 10 9 13 1 9 2 13 0 9 2
30 1 9 0 9 13 0 9 9 1 9 0 11 11 2 11 7 11 11 2 11 0 1 10 9 0 9 1 9 0 2
24 9 13 9 2 15 9 13 1 9 0 9 2 7 13 7 9 3 3 0 16 13 0 9 2
11 3 13 1 10 9 3 16 12 9 0 2
37 16 0 9 9 15 1 10 12 9 3 13 2 0 9 1 10 9 13 9 1 15 2 15 10 9 0 9 13 16 0 7 15 15 13 1 9 2
11 7 13 10 9 13 2 16 10 9 13 2
24 7 16 4 13 4 13 9 1 9 2 13 4 1 9 1 9 0 9 0 2 3 0 9 2
18 12 1 0 13 1 15 2 16 9 2 15 3 13 9 2 15 13 2
27 3 13 0 13 9 1 0 9 3 1 9 7 9 2 1 9 2 9 7 9 3 15 1 12 9 13 2
18 3 13 3 12 1 10 9 2 16 9 15 13 3 7 3 3 0 2
16 7 3 2 1 0 0 9 7 9 0 9 13 3 0 9 2
22 1 0 9 13 10 15 0 2 16 7 1 0 9 13 4 13 1 0 14 10 9 2
35 0 9 9 9 2 15 13 9 2 4 1 10 9 13 9 2 9 2 9 2 9 2 9 0 9 2 9 2 9 7 0 9 0 9 2
22 1 0 9 9 13 10 9 12 2 12 9 9 2 9 2 9 2 2 1 11 2 2
17 3 1 3 0 9 13 0 13 16 3 0 3 16 12 9 11 2
14 3 13 15 2 16 3 0 9 4 1 9 9 13 2
13 16 15 13 3 3 0 2 3 15 13 3 13 2
15 10 9 13 2 16 15 9 2 9 7 9 13 9 9 2
31 3 7 13 2 16 9 9 7 9 13 10 0 9 1 0 9 2 7 16 10 9 0 9 3 13 2 15 13 0 9 2
36 13 15 0 2 16 0 9 0 9 9 1 11 13 2 16 12 9 15 13 2 16 9 4 13 4 13 3 1 0 9 16 0 9 9 9 2
29 10 9 13 3 0 2 15 13 0 9 2 7 1 9 9 9 12 2 9 4 3 13 13 2 16 15 13 3 2
41 9 1 9 2 12 2 12 2 12 2 12 2 12 2 12 13 1 9 11 11 2 0 9 0 9 13 14 13 2 0 9 9 2 9 12 2 9 2 12 2 12
7 9 2 11 11 2 9 2
11 2 2 12 2 13 9 1 0 9 11 2
14 1 9 9 7 9 10 9 15 13 0 7 0 9 2
7 9 2 11 11 2 9 2
9 2 2 12 2 13 0 9 11 2
10 13 1 0 9 7 13 15 1 9 2
7 9 2 11 11 2 9 2
11 2 2 12 2 13 0 9 11 1 11 2
15 13 15 0 9 1 0 9 12 2 0 9 11 1 11 2
7 9 2 11 11 2 9 2
11 2 2 12 2 13 0 9 11 1 11 2
21 1 9 0 0 9 9 0 9 11 15 13 9 0 9 0 9 7 9 0 9 2
15 9 2 11 11 2 2 12 2 13 0 9 11 1 11 2
9 1 9 9 1 11 15 13 9 2
9 9 2 9 2 11 11 2 9 2
10 2 2 12 2 13 11 11 1 11 2
11 1 9 9 0 9 11 15 13 9 9 2
7 9 2 11 11 2 9 2
17 2 2 12 2 13 9 2 9 7 9 1 0 9 11 1 11 2
14 1 0 9 1 11 15 13 9 0 9 7 9 11 2
7 9 2 11 11 2 9 2
13 2 2 12 2 13 9 0 9 1 11 1 11 2
13 1 9 0 9 1 9 15 13 9 9 0 9 2
14 11 11 2 2 12 2 13 9 1 0 9 1 11 2
15 4 13 1 9 9 11 1 11 7 13 15 9 7 9 2
21 9 2 9 2 11 0 2 9 2 2 2 2 12 2 13 0 9 11 1 11 2
23 13 9 9 0 7 0 9 2 13 15 9 9 2 9 2 9 7 13 9 0 9 9 2
14 9 2 11 11 2 2 12 2 13 0 9 1 11 2
12 1 0 9 10 9 15 13 9 0 0 9 2
5 9 9 0 9 2
21 14 4 15 13 15 1 9 0 9 2 14 4 13 3 7 13 1 9 14 3 2
7 3 13 3 3 0 9 2
25 15 9 13 1 9 7 9 1 9 7 13 9 1 9 2 3 13 2 7 0 9 15 13 9 2
16 15 13 9 0 1 9 9 7 9 2 1 9 11 11 2 2
35 1 9 0 2 0 2 0 7 0 9 9 13 9 0 2 0 2 9 9 7 9 2 7 2 16 13 11 2 9 4 13 9 1 9 2
15 7 1 0 9 2 0 2 0 7 0 2 13 9 9 2
29 7 9 3 0 15 1 10 9 13 2 0 9 2 0 9 2 9 9 13 1 9 7 3 7 9 13 3 0 2
9 3 9 7 9 13 3 1 9 2
10 13 3 10 9 9 2 13 0 9 2
14 13 15 15 2 16 9 11 11 13 9 9 0 9 2
9 14 7 14 1 9 9 0 9 2
8 10 9 13 3 0 7 0 2
20 13 3 1 12 1 0 9 9 2 1 11 2 1 9 14 0 2 7 0 2
37 1 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 7 3 1 0 0 9 2 9 7 9 9 2
22 13 15 3 9 1 0 9 2 13 15 9 7 9 9 2 15 13 2 13 7 13 2
18 7 13 15 9 0 0 9 7 13 9 2 16 0 2 0 7 0 2
19 7 13 15 15 2 16 11 11 13 10 9 3 2 16 15 13 10 9 2
14 0 13 9 1 0 9 7 9 2 0 13 9 9 2
24 0 0 9 7 9 13 16 9 9 2 9 2 0 9 2 0 1 9 7 0 9 0 9 2
12 9 7 9 11 11 13 3 13 1 0 9 2
16 15 13 2 3 0 1 10 9 13 9 9 2 9 0 9 2
19 1 9 9 11 11 1 11 1 11 13 0 9 2 3 3 0 10 9 2
19 15 1 15 13 2 15 13 2 7 0 9 13 1 15 3 0 9 9 2
11 1 9 13 9 0 9 0 1 9 9 2
7 7 1 15 13 0 9 2
13 11 15 13 9 1 9 2 15 13 2 3 2 2
21 13 15 7 15 2 13 7 2 16 0 9 3 13 2 16 3 14 1 0 9 2
4 13 14 13 2
8 3 9 0 1 0 9 13 2
9 7 3 15 15 1 0 13 0 2
2 11 11
3 0 9 2
4 13 15 0 9
4 1 9 0 9
5 1 9 9 0 2
2 11 11
16 0 9 4 13 7 13 3 0 9 1 10 9 1 0 9 2
26 9 1 0 9 15 13 1 9 3 0 9 0 9 7 0 9 7 9 4 13 1 0 9 7 9 2
24 7 14 13 9 2 16 0 9 16 0 9 3 13 2 7 3 3 2 16 13 7 0 9 2
34 0 9 4 13 7 9 9 2 7 3 9 9 2 15 15 13 2 7 0 0 9 7 0 0 9 2 1 15 9 1 10 9 13 2
24 0 9 13 0 9 16 0 0 9 2 0 9 2 2 7 2 13 15 13 9 1 0 9 2
13 13 15 7 1 9 0 9 2 9 9 0 9 2
10 7 3 13 0 0 9 0 0 9 2
20 0 7 0 9 13 1 0 9 14 0 10 0 9 2 7 3 7 1 15 2
41 10 3 0 9 13 1 9 2 16 0 9 13 14 3 0 9 2 10 9 13 0 9 1 9 2 7 0 9 13 3 14 3 0 9 2 10 9 13 0 9 2
24 16 4 13 9 0 2 13 0 15 13 3 1 0 0 9 2 15 1 9 12 9 3 13 2
36 7 1 3 0 0 9 13 9 9 2 15 1 0 7 0 9 1 9 9 9 13 9 2 1 10 9 1 9 13 3 9 0 16 9 0 2
20 3 13 0 9 1 9 10 9 0 9 7 13 9 9 1 9 9 0 9 2
46 3 13 1 10 9 3 3 3 2 16 13 13 0 9 9 1 9 1 9 1 9 11 2 1 0 9 2 16 1 10 9 13 13 1 9 0 3 1 0 9 2 3 1 12 9 2
63 1 9 13 3 0 9 9 2 15 13 0 0 9 1 0 9 7 9 2 1 15 1 0 9 13 2 16 1 9 9 9 9 9 2 12 1 12 2 9 0 0 9 2 3 0 0 9 2 15 13 1 0 9 9 1 9 12 16 9 1 9 12 2
57 1 0 9 3 1 12 9 0 7 14 0 9 3 13 3 0 9 0 9 2 16 1 9 9 9 9 9 2 12 1 12 2 9 0 0 9 2 3 0 0 9 2 15 13 1 0 9 9 1 9 12 16 9 1 9 12 2
13 10 9 13 0 9 1 9 0 9 16 0 9 2
37 1 1 15 2 16 9 13 9 1 9 0 9 2 7 3 13 0 9 1 9 1 10 9 2 13 0 3 0 9 16 0 9 1 9 3 0 2
11 15 15 7 3 3 3 13 1 10 9 2
39 7 0 9 2 15 9 13 2 13 3 10 0 1 9 9 2 7 7 0 9 2 15 9 1 10 9 13 2 13 3 3 9 0 9 16 9 0 9 2
8 0 9 13 9 9 0 0 9
13 3 0 9 13 3 0 9 9 16 9 0 9 2
7 0 13 3 9 1 9 2
25 16 0 9 9 2 9 7 9 13 13 0 9 3 9 9 2 0 9 13 3 9 7 9 9 2
23 15 13 0 9 3 2 1 9 9 9 0 9 2 9 2 15 13 0 9 0 9 9 2
10 0 9 7 3 13 0 7 7 0 2
29 0 13 2 16 1 0 9 3 0 9 13 3 1 9 13 2 16 13 3 0 2 7 2 16 13 9 10 9 2
15 10 9 15 1 9 9 13 9 0 0 9 2 9 2 2
22 0 9 0 9 13 0 9 2 9 0 9 1 10 9 9 2 15 13 10 0 9 2
10 10 9 13 9 9 1 9 0 9 2
27 16 1 10 9 13 1 10 9 1 9 1 9 2 3 3 1 9 12 9 0 2 13 13 3 12 9 2
21 1 9 9 3 7 3 15 9 0 9 2 9 2 2 9 0 0 9 2 13 2
19 1 3 0 9 3 13 15 9 0 9 7 1 9 13 3 9 0 9 2
8 1 10 9 13 1 9 9 2
47 16 13 9 12 9 7 12 9 2 3 0 9 2 1 9 9 0 2 15 13 1 9 2 1 9 15 9 0 9 0 9 1 0 9 2 0 9 1 12 9 2 1 12 1 0 9 2
31 2 1 0 3 13 1 0 9 0 9 1 9 0 9 2 1 9 9 7 9 10 9 2 0 9 2 13 10 9 2 2
27 16 15 1 0 9 10 9 13 0 9 2 3 1 9 12 2 12 13 1 3 0 9 9 1 10 9 2
20 1 9 12 2 12 4 3 0 9 3 7 3 13 2 15 9 0 9 13 2
29 16 4 13 0 9 3 0 2 13 4 1 9 0 9 1 3 0 9 2 1 9 0 0 0 9 4 15 13 2
16 16 4 13 9 9 3 3 0 2 13 4 9 9 3 0 2
12 1 3 0 9 7 3 13 3 3 0 9 2
27 15 13 1 9 2 16 1 9 0 9 13 3 0 9 2 0 1 9 9 0 9 7 0 1 9 9 2
67 16 15 13 1 10 9 0 9 7 16 13 1 9 2 16 9 9 0 9 13 1 9 3 12 5 12 2 12 1 9 7 9 7 9 0 0 9 16 13 3 12 5 12 12 9 9 2 3 13 2 16 1 12 0 9 2 1 12 9 2 13 13 9 14 12 9 2
25 15 13 2 16 9 3 0 0 9 1 9 2 10 9 15 13 2 13 3 1 9 12 0 9 2
25 16 13 12 9 3 0 9 2 7 2 1 10 9 13 1 9 2 13 15 1 0 9 0 9 2
49 16 13 1 0 9 0 7 0 9 1 3 0 9 0 2 16 13 15 3 1 9 9 1 9 0 9 2 13 9 9 0 9 2 15 13 0 9 0 2 13 2 1 10 9 15 0 9 13 2
30 16 4 3 13 2 16 1 9 9 13 1 15 9 0 9 2 7 16 13 0 0 9 2 13 3 13 9 0 9 2
17 9 0 9 9 15 7 13 13 16 0 9 0 13 9 0 9 2
15 13 0 13 2 16 4 14 3 13 1 9 9 3 0 2
27 1 15 15 1 9 13 7 9 2 15 3 0 13 2 15 10 9 2 3 7 3 2 13 9 10 9 2
20 9 10 9 13 0 9 2 9 0 9 2 7 0 9 2 16 9 9 0 2
18 3 13 3 0 2 3 0 9 9 13 3 0 7 3 0 3 0 2
10 3 15 13 2 16 0 9 3 13 2
26 1 0 9 13 0 2 16 13 9 1 9 0 13 1 3 0 9 2 7 15 1 3 12 5 9 2
5 3 15 7 13 2
39 16 15 3 9 13 1 9 9 0 9 2 7 16 13 1 0 9 2 9 2 15 15 13 9 12 9 1 9 1 0 2 3 3 3 13 1 9 0 2
42 16 7 13 0 9 1 9 9 9 1 0 9 2 3 4 13 0 13 3 0 0 7 3 0 9 2 16 4 13 13 2 16 0 9 13 2 7 13 9 0 9 2
15 9 1 3 0 7 3 0 9 13 1 9 9 3 0 2
31 16 1 0 9 13 2 16 9 0 9 1 12 9 2 9 7 9 13 9 10 0 9 2 1 9 3 0 10 9 13 2
28 9 0 3 0 9 3 13 3 3 9 0 9 2 15 4 0 9 7 9 13 2 16 9 10 0 0 9 2
15 1 9 3 0 9 15 3 13 1 9 0 7 0 9 2
34 16 12 9 9 13 1 0 9 2 4 13 0 0 9 2 3 13 10 9 3 3 2 13 15 1 15 0 0 9 7 0 9 9 2
32 7 1 9 2 16 15 3 13 1 9 0 2 13 3 1 10 0 9 2 9 13 0 9 2 13 15 12 0 3 3 13 2
21 16 9 0 9 15 3 13 9 9 2 9 7 9 7 9 10 9 7 0 9 2
17 3 9 13 3 3 0 1 9 2 9 7 9 16 1 0 9 2
21 3 9 13 2 3 1 9 13 2 3 0 1 9 2 9 7 9 16 1 9 2
24 16 4 15 7 13 13 10 9 1 9 0 9 2 15 4 13 13 9 7 9 1 0 9 2
22 4 15 13 15 2 16 12 10 9 13 1 9 3 0 9 2 12 13 3 0 9 2
13 4 7 13 0 0 9 2 16 10 9 13 3 2
16 9 15 13 13 0 7 0 9 1 9 9 2 3 9 9 2
29 9 9 13 0 9 2 9 2 15 13 9 9 0 9 9 2 7 2 9 0 9 0 9 9 1 0 0 9 2
18 1 9 0 9 3 13 1 0 9 0 9 2 13 15 3 10 9 2
58 13 14 0 1 10 9 13 2 16 9 9 13 15 0 1 9 2 0 9 2 15 4 1 9 3 13 7 1 9 9 2 13 9 12 2 12 2 12 2 12 2 12 2 12 2 12 2 12 2 12 2 12 2 12 2 12 2 2
11 9 0 9 0 9 13 3 15 3 0 2
18 13 3 9 9 9 7 4 7 13 2 7 13 2 0 7 0 9 2
8 13 7 0 9 1 9 9 2
38 1 15 9 0 2 3 0 7 0 2 13 1 10 9 3 3 0 2 7 13 2 14 15 13 1 9 9 2 13 0 1 15 13 1 0 0 9 2
25 0 9 7 13 3 3 0 9 1 9 0 9 9 2 9 9 7 9 9 2 2 1 9 9 2
34 9 13 3 13 16 9 0 9 2 9 9 7 9 0 9 2 7 2 0 7 0 9 3 9 9 2 0 1 9 9 9 1 9 2
21 1 9 9 15 0 9 9 13 2 12 1 0 15 3 13 2 13 2 13 15 2
21 9 2 1 15 1 0 9 13 2 13 4 13 3 0 9 2 7 7 0 9 2
19 13 0 2 16 9 9 2 9 0 9 2 4 1 9 9 13 0 9 2
22 1 0 9 9 0 2 3 9 15 15 13 1 9 9 2 4 13 3 3 0 9 2
21 1 9 0 9 7 0 9 13 0 13 1 9 12 9 0 9 2 9 7 9 2
38 3 9 9 15 13 13 2 10 9 15 0 9 1 9 9 13 2 7 3 9 9 15 13 9 2 10 0 9 13 0 13 7 3 3 10 9 13 2
26 16 13 1 15 3 9 9 9 2 13 1 15 3 13 2 16 4 13 0 9 9 13 1 0 9 2
43 16 7 13 3 1 9 7 9 1 9 1 0 0 9 2 9 1 9 7 0 9 0 9 9 2 13 3 0 2 16 9 13 0 1 9 9 13 7 13 15 0 9 2
8 13 2 1 9 13 2 2 2
35 1 9 4 13 3 0 9 0 9 1 9 0 9 2 9 9 2 15 4 13 9 0 9 7 3 13 7 13 1 9 0 9 9 0 2
10 1 9 15 3 13 3 13 9 9 2
22 1 0 9 13 1 0 9 9 13 2 16 15 9 1 0 9 3 3 13 1 0 2
47 9 10 0 9 13 9 0 3 0 9 2 0 0 9 2 9 0 7 1 10 9 3 1 0 9 9 2 0 0 9 2 13 3 9 12 2 12 2 12 2 12 2 12 2 12 2 2
29 10 9 3 13 9 3 15 3 0 9 7 13 14 9 9 2 16 3 3 13 7 9 0 2 0 7 0 9 2
19 9 13 2 1 0 2 13 7 13 3 0 9 9 0 1 0 9 9 2
29 13 3 3 0 2 16 13 13 7 1 3 0 9 9 2 15 13 13 1 0 9 2 3 12 9 7 12 9 2
24 0 9 3 13 13 1 0 9 0 2 16 13 0 3 13 3 9 9 0 1 0 0 9 2
17 0 7 14 13 2 16 13 1 9 3 0 2 0 0 0 9 2
25 9 9 0 1 3 0 9 7 0 1 0 0 9 15 3 3 13 9 1 9 1 9 3 0 2
26 10 9 3 13 2 16 9 13 13 0 9 1 9 0 9 3 2 3 3 13 2 1 9 9 0 2
20 9 9 0 13 3 0 9 9 2 15 0 9 1 0 9 13 9 0 9 2
1 9
2 9 9
3 0 9 2
3 11 2 9
2 11 11
8 9 1 2 9 9 9 2 9
2 11 11
5 9 9 0 9 11
5 11 11 2 11 11
3 0 9 2
2 11 11
4 9 1 0 9
2 11 11
8 9 2 9 2 7 0 9 2
2 11 11
5 9 0 9 0 9
2 11 11
7 11 11 2 9 9 7 9
2 11 11
2 11 11
8 9 9 1 9 9 7 9 9
2 11 11
5 0 9 13 15 9
2 11 11
2 0 9
2 11 11
7 2 0 2 7 2 0 2
2 11 11
3 1 9 9
3 9 7 9
2 9 9
1 9
5 9 2 9 7 9
3 9 1 9
11 11 11 2 9 9 2 9 7 9 1 9
4 9 1 10 9
1 9
4 1 9 7 9
3 9 7 9
3 9 1 9
4 13 4 1 9
1 9
3 0 0 9
7 9 9 1 9 9 1 11
2 0 9
1 9
7 2 9 2 9 9 9 9
5 9 9 13 0 9
6 1 0 9 2 2 2
9 3 13 9 0 9 1 0 2 9
2 0 9
6 0 9 2 14 0 9
2 0 9
6 2 13 1 9 9 2
2 0 9
7 11 11 2 9 9 0 9
7 11 11 2 9 1 9 9
1 11
1 9
6 9 1 12 9 9 9
7 9 1 2 9 9 9 2
2 11 11
31 1 15 2 3 4 13 1 9 0 9 1 0 9 1 0 9 1 11 2 4 3 13 2 9 12 2 12 2 12 2 2
19 9 4 3 13 1 0 9 9 2 0 9 1 9 9 2 9 9 0 2
5 3 13 9 0 2
5 13 15 3 9 2
48 9 9 2 12 11 2 11 7 11 2 11 1 0 9 2 11 2 13 1 9 11 2 12 2 12 2 12 2 9 2 1 15 13 0 9 0 2 3 13 13 0 0 9 9 1 9 13 2
27 9 2 16 4 15 10 9 13 13 12 0 9 2 15 13 1 12 2 12 9 14 1 12 2 12 9 2
29 1 9 9 4 15 7 13 14 3 2 16 4 15 9 1 15 3 3 3 13 2 16 13 9 1 0 2 9 2
20 15 13 1 3 0 0 2 9 2 1 0 0 9 1 15 9 0 1 9 2
19 14 1 11 7 13 0 0 9 0 1 2 0 2 2 3 15 0 9 2
19 3 13 1 15 9 2 3 15 9 1 9 13 10 0 9 1 0 9 2
23 3 9 1 0 0 9 13 7 0 9 1 0 9 13 4 13 3 1 12 7 12 9 2
31 13 3 9 2 16 4 15 3 14 13 13 9 1 0 9 2 15 4 3 13 3 3 2 16 4 0 13 4 3 13 2
15 16 4 10 9 13 2 13 9 9 1 9 1 9 13 2
20 2 13 4 15 15 13 3 7 9 11 2 13 9 12 2 12 2 12 2 2
10 0 9 4 13 14 12 2 12 9 2
38 1 0 9 11 4 13 9 0 9 11 2 11 1 9 1 11 2 11 2 7 11 2 11 2 11 1 0 9 2 11 2 2 15 1 0 9 13 2
35 13 3 0 0 9 9 0 9 0 9 1 12 9 2 7 7 9 0 15 9 0 9 2 9 2 9 2 12 2 9 9 3 2 2 2
8 9 0 9 15 1 15 13 2
31 3 3 1 0 9 12 9 13 2 16 9 9 10 9 15 3 7 3 13 1 0 9 2 15 4 3 3 13 3 13 2
16 0 9 13 2 16 9 3 9 13 3 0 16 1 9 3 2
27 0 0 9 13 0 0 9 2 15 13 0 9 0 1 0 9 2 7 10 9 13 1 9 1 0 9 2
7 3 4 15 3 15 13 2
12 4 1 15 13 14 12 0 9 1 0 9 2
5 7 15 13 9 2
33 0 9 15 13 1 0 9 2 3 3 9 9 9 13 4 1 9 13 16 3 0 7 13 13 9 2 16 15 15 3 13 9 2
17 3 4 15 13 13 2 16 4 13 9 9 9 1 0 9 3 2
29 3 9 11 7 11 4 3 3 3 1 0 9 13 1 12 9 1 11 7 13 13 1 9 1 9 7 0 9 2
13 9 9 9 9 3 13 9 7 13 1 15 13 2
20 10 9 1 11 4 13 7 9 4 13 9 1 0 9 2 0 1 0 9 2
13 11 7 11 10 9 13 1 2 9 1 9 2 2
14 7 16 12 9 1 9 9 13 2 13 15 0 9 2
29 1 0 9 13 7 9 1 0 9 0 1 9 11 2 0 9 15 9 7 9 2 11 12 2 12 2 12 2 2
19 13 15 3 13 7 7 15 13 14 12 9 2 1 15 15 13 0 9 2
18 9 15 13 1 9 9 9 7 13 15 9 0 9 9 11 7 11 2
7 13 15 2 15 13 2 2
13 15 9 9 13 0 9 0 9 1 9 2 12 2
13 2 7 15 3 3 13 2 3 15 3 13 2 2
19 9 0 9 9 9 13 3 10 0 9 1 9 2 15 15 9 9 13 2
14 9 0 9 13 0 2 11 12 2 12 2 12 2 2
52 0 13 2 16 1 9 2 13 2 3 2 1 15 0 9 11 2 11 2 11 1 0 9 1 0 11 2 11 2 2 15 1 9 13 9 9 1 0 9 2 0 9 1 0 9 12 2 12 2 12 2 2
5 13 3 0 9 2
7 0 9 15 13 1 11 2
21 13 0 2 16 15 10 9 13 1 9 1 9 2 12 2 15 3 13 15 9 2
15 4 1 15 2 3 2 13 0 9 3 1 0 9 9 2
24 1 0 9 4 1 9 11 13 7 13 0 9 7 1 10 9 4 13 0 9 1 9 9 2
21 0 9 15 3 13 13 15 2 16 4 13 12 9 9 0 9 7 9 3 13 2
16 13 15 0 9 2 15 15 13 1 9 13 1 9 0 9 2
28 15 4 7 13 1 9 13 0 9 9 1 9 1 0 9 7 1 9 0 9 2 15 4 1 9 9 13 2
14 3 4 1 11 13 9 2 15 13 9 9 1 9 2
18 13 7 13 14 9 1 0 9 7 9 0 1 9 2 15 4 13 2
17 1 10 9 15 13 13 7 7 9 9 2 15 13 1 9 13 2
6 7 9 13 1 9 2
21 9 0 9 0 9 9 3 7 13 0 9 7 13 15 1 0 9 1 0 9 2
48 9 9 1 15 3 3 1 9 2 3 13 0 1 15 2 13 2 16 9 0 9 13 1 9 13 2 7 9 7 13 1 10 0 9 1 9 3 2 11 12 2 12 7 12 2 12 2 2
26 3 15 15 7 9 0 9 1 0 9 3 7 3 13 7 3 15 10 9 3 2 13 2 10 9 2
24 7 0 9 1 11 2 11 1 9 1 11 15 3 13 13 0 9 2 15 13 10 0 9 2
19 13 15 1 15 9 1 9 1 9 0 7 9 1 9 9 3 0 9 2
24 9 9 15 13 1 0 2 9 2 13 9 12 2 12 2 12 2 12 2 12 2 12 2 2
13 1 9 1 0 7 0 9 9 13 9 9 0 2
13 2 0 7 0 9 13 3 9 1 10 9 2 2
18 7 15 3 0 9 7 9 13 3 13 1 9 3 0 9 0 9 2
55 11 2 11 2 11 1 9 1 11 2 3 10 9 2 15 13 1 0 9 9 11 7 11 1 9 2 12 2 13 9 12 2 12 2 12 2 7 13 0 9 2 13 1 10 9 1 10 9 1 3 0 7 0 9 2
27 0 9 2 9 9 9 2 13 9 1 9 3 0 9 1 0 0 9 0 9 2 1 0 2 0 9 2
7 3 15 13 7 13 9 2
21 10 9 4 13 0 9 12 7 3 9 0 0 9 2 0 3 2 12 9 2 2
32 16 0 9 13 3 0 9 0 9 9 2 0 9 13 3 7 13 13 2 1 10 9 15 0 9 0 9 1 0 9 13 2
8 3 3 4 13 9 0 9 2
34 0 0 9 13 9 0 9 0 2 7 0 9 15 13 15 0 2 3 3 0 9 2 1 15 15 3 13 9 9 1 0 0 9 2
22 10 9 3 13 15 2 16 15 0 9 13 9 3 15 0 2 9 2 1 12 9 2
19 16 3 3 13 9 9 2 13 4 15 10 9 3 13 2 0 9 2 2
13 9 13 3 1 9 2 7 13 9 1 0 9 2
41 13 2 14 15 3 10 9 2 3 1 9 2 1 15 4 1 0 9 13 9 9 1 9 2 15 1 15 3 13 1 0 9 2 11 12 2 12 2 12 2 2
29 7 16 9 13 1 9 1 9 9 1 10 2 0 9 2 2 13 15 3 10 3 0 9 2 9 9 9 2 2
15 10 9 4 13 1 0 9 2 1 15 13 9 0 9 2
23 2 0 9 2 3 13 1 9 10 0 9 1 0 9 7 15 7 1 9 0 9 9 2
33 7 9 10 9 4 3 1 9 9 13 13 13 9 1 0 2 9 0 2 2 15 13 0 7 0 9 0 9 11 9 2 12 2
5 11 2 0 9 2
10 9 9 1 9 0 9 10 9 0 2
12 9 9 2 9 4 13 1 9 9 7 13 2
19 10 9 0 9 13 9 2 16 13 13 2 16 9 13 1 9 0 9 0
1 12
2 12 2
4 9 9 9 2
15 1 0 9 15 13 0 9 0 9 1 12 3 0 9 2
33 1 0 15 9 0 9 13 1 9 12 9 0 9 2 9 0 1 12 7 0 9 9 2 0 1 15 9 9 2 15 13 13 2
15 1 0 9 1 9 9 2 9 13 0 9 1 9 0 2
30 16 9 13 13 9 9 1 0 9 7 13 13 0 9 9 3 1 12 9 2 13 1 9 3 1 9 0 0 9 2
14 1 0 9 7 0 15 0 9 13 2 13 9 12 2
32 1 0 9 15 9 9 0 9 13 2 16 1 12 9 15 9 0 15 3 1 9 1 0 9 13 14 3 2 12 12 7 2
10 11 2 9 1 2 9 9 9 2 2
11 9 9 9 3 0 9 2 0 9 2 2
12 9 1 9 7 9 0 13 13 1 9 9 2
7 9 1 9 13 0 7 0
10 11 2 11 2 9 9 2 2 2 2
29 9 9 9 1 0 9 2 12 2 9 2 12 2 0 9 0 1 9 9 2 12 2 0 9 0 1 0 9 2
23 9 1 0 9 13 0 2 2 0 2 2 7 4 13 7 13 7 9 0 9 2 0 2
9 12 2 9 2 0 9 0 0 9
19 9 0 9 0 9 2 0 9 2 7 3 0 0 9 2 0 9 2 2
29 0 0 9 3 0 0 9 2 15 15 3 13 1 0 9 9 2 13 9 9 0 0 9 7 9 10 0 9 2
14 2 9 1 3 0 9 13 0 9 0 1 0 9 2
22 16 1 0 9 13 9 3 0 9 9 9 2 13 0 9 0 9 1 12 9 0 2
2 11 2
8 13 15 3 2 13 4 13 2
3 9 11 11
8 11 2 0 9 13 15 9 2
19 9 0 9 7 9 0 9 1 0 7 0 9 2 11 7 0 2 12 2
20 9 2 1 15 13 0 9 3 0 9 9 2 4 13 1 9 9 1 9 2
17 9 13 2 16 0 9 13 0 9 2 7 13 3 0 1 9 2
33 9 0 7 0 0 9 2 1 9 9 7 1 9 0 9 1 9 9 9 2 13 9 1 9 0 1 9 7 9 0 1 9 2
13 2 9 9 4 13 9 9 1 9 1 9 2 2
17 9 9 9 9 1 0 9 13 1 3 0 9 9 9 0 9 2
21 0 9 13 0 9 9 2 2 0 9 2 2 1 0 9 7 13 7 0 9 2
13 2 9 9 4 13 9 9 1 9 1 9 2 2
22 9 9 9 7 0 9 1 0 9 2 15 13 1 0 9 1 9 1 12 9 9 2
17 9 9 4 13 1 9 2 1 15 15 13 9 9 1 0 9 2
12 1 9 9 15 13 9 9 9 0 0 9 2
11 0 9 1 9 13 9 2 3 4 13 9
5 11 2 0 9 2
3 0 9 2
13 11 11 2 0 2 12 2 12 2 12 1 11 2
13 1 9 12 2 12 13 1 9 0 9 1 11 2
11 1 9 2 12 13 9 1 9 0 9 2
8 2 0 2 7 2 0 2 2
2 11 11
24 13 3 3 13 2 16 13 15 15 13 1 9 0 9 2 3 3 2 16 1 9 9 15 2
1 12
28 9 2 0 2 7 2 0 2 2 7 2 0 2 7 2 0 2 4 13 1 0 9 9 2 9 7 9 2
22 9 9 0 9 13 1 9 1 9 0 13 0 9 0 3 1 2 9 2 0 9 2
21 13 15 7 9 9 7 0 9 9 3 13 2 3 13 10 9 0 7 3 0 2
48 3 15 7 13 2 16 15 1 9 9 9 13 2 16 9 1 9 2 1 9 1 0 9 2 13 13 9 2 16 9 0 9 13 14 9 0 0 9 2 1 15 3 13 9 0 1 0 2
8 0 2 0 2 9 13 9 2
32 13 2 14 9 7 9 2 9 0 2 2 13 15 0 9 2 1 9 2 1 9 9 2 15 15 3 13 16 2 0 2 2
6 10 13 1 15 9 2
17 9 9 7 9 13 2 16 0 9 4 13 1 9 0 9 9 2
17 13 15 3 0 0 9 2 15 13 9 1 9 9 1 9 9 2
17 9 13 9 0 2 16 9 9 13 1 9 1 3 0 9 9 2
38 0 9 13 13 0 7 0 9 1 9 7 1 0 9 7 13 15 13 14 1 9 0 9 7 0 9 2 0 9 13 1 15 10 9 3 0 2 2
6 9 9 3 3 13 2
14 10 15 13 1 0 9 13 3 3 1 0 9 9 2
28 9 9 13 7 3 0 9 9 2 7 13 3 10 0 9 16 9 9 2 7 7 13 13 9 15 1 9 2
41 9 4 3 13 15 2 16 0 9 13 1 9 1 9 2 3 9 1 9 13 13 2 16 0 2 3 0 9 15 3 13 1 15 2 16 4 3 1 9 13 2
20 7 12 9 9 13 13 16 2 0 2 2 7 0 13 10 9 1 15 13 2
16 1 0 9 15 3 13 2 16 0 0 9 13 0 16 0 2
24 0 9 2 16 0 9 13 9 13 1 10 0 9 7 13 15 1 9 2 15 13 16 0 2
43 3 15 13 3 3 13 2 16 0 9 4 3 13 1 10 9 1 9 13 2 0 2 2 0 9 2 15 13 9 14 0 2 15 15 3 13 13 0 9 9 7 9 2
22 16 9 13 1 9 2 13 15 9 0 9 2 3 9 2 15 15 13 1 0 9 2
35 3 1 12 9 9 13 1 9 0 9 0 9 1 0 11 1 0 9 0 9 1 0 11 7 1 0 9 0 9 9 0 2 1 9 2
6 0 9 13 3 9 2
14 13 7 10 9 0 9 3 0 2 3 15 3 13 2
14 1 0 9 13 9 1 0 11 14 3 3 0 9 2
4 13 3 0 2
12 9 9 3 13 13 9 9 14 1 0 9 2
13 7 9 13 3 1 9 2 15 15 13 13 0 2
8 13 7 13 1 0 9 0 2
20 1 0 0 9 0 9 0 13 3 3 0 2 3 7 3 13 9 0 9 2
41 9 15 13 1 2 0 2 7 2 0 2 7 1 0 9 2 9 2 9 7 9 13 0 2 15 15 3 13 1 0 9 2 16 9 7 9 13 0 2 0 2
30 9 13 1 10 0 9 3 2 0 2 16 9 2 7 10 0 9 15 13 1 0 9 1 12 14 1 12 9 9 2
32 9 7 13 13 0 9 1 9 2 3 13 10 9 7 3 4 0 9 2 1 15 9 1 10 0 0 9 2 3 13 9 2
6 3 13 15 1 9 2
25 3 0 0 9 15 3 1 0 9 11 13 1 9 2 16 9 3 13 3 9 16 3 0 9 2
30 16 9 13 9 0 9 1 9 9 2 13 9 0 9 2 7 0 9 1 9 0 9 13 10 9 1 9 0 9 2
22 9 4 1 3 0 9 13 1 0 7 0 9 2 0 14 0 9 7 0 0 9 2
47 1 0 9 2 3 0 9 2 15 13 2 16 9 13 14 0 0 9 2 10 9 4 13 3 1 9 0 9 10 9 2 7 13 13 0 9 7 9 0 9 2 9 9 9 9 2 2
47 1 9 0 9 1 9 2 9 7 0 9 13 13 7 1 9 1 9 2 3 1 10 9 2 7 1 0 9 0 9 13 3 13 9 2 16 9 0 9 15 13 1 9 9 3 9 2
36 9 0 9 0 1 3 0 9 3 3 13 1 9 2 7 15 1 0 9 2 16 13 3 3 13 15 2 16 10 9 13 2 15 13 9 2
35 0 9 2 3 0 9 2 16 9 13 1 9 1 3 2 0 2 9 2 13 2 7 12 9 13 1 15 1 9 0 16 12 9 9 2
43 0 9 13 1 0 10 3 0 9 14 3 0 9 1 2 9 9 2 7 9 13 3 1 10 9 2 15 15 3 13 9 2 7 0 9 2 1 10 9 15 13 9 2
34 1 0 9 9 13 0 9 1 0 9 9 2 0 2 0 3 0 9 9 9 2 0 2 2 7 1 10 9 13 9 1 0 9 2
27 9 3 13 2 16 9 2 0 2 7 2 0 2 13 3 9 0 9 1 0 9 2 16 3 0 9 2
52 15 15 13 14 9 7 9 2 7 3 10 0 9 2 16 3 2 9 7 9 2 9 13 3 2 7 4 1 9 9 13 0 9 0 9 2 16 9 3 13 0 9 2 7 15 3 14 1 0 9 2 2
43 3 4 13 7 0 9 2 16 9 13 2 0 2 9 16 9 2 7 0 9 0 9 13 9 1 0 9 2 9 0 9 7 0 9 9 7 9 15 1 0 9 13 2
22 9 2 15 15 13 2 13 0 9 9 2 1 15 4 13 0 12 9 13 1 0 2
22 16 9 3 10 9 13 2 13 1 9 1 0 9 14 3 0 2 7 7 3 0 2
7 15 15 13 7 11 11 2
50 1 9 10 9 15 3 13 2 16 1 10 9 13 9 3 3 0 9 11 11 2 9 1 0 0 9 1 9 2 2 15 13 3 9 12 2 9 4 13 14 3 7 13 15 3 0 9 9 2 2
30 1 10 9 11 13 9 2 3 13 0 9 2 0 2 7 2 0 2 2 3 13 9 2 0 2 7 2 0 2 2
6 0 9 2 14 0 9
12 1 9 1 0 9 13 3 13 11 3 3 2
13 13 2 16 1 10 9 13 9 9 1 15 9 2
44 0 0 9 1 11 13 2 16 9 9 9 13 1 12 9 2 1 9 12 9 2 2 9 0 1 12 2 1 12 9 2 7 0 0 9 15 13 1 9 1 12 9 3 2
11 0 3 13 3 0 9 9 9 1 9 2
2 11 11
3 12 2 12
3 9 0 9
40 9 0 9 3 13 2 7 2 16 4 13 9 9 0 1 9 9 2 2 15 13 0 9 9 2 2 13 1 10 9 9 9 2 2 0 1 0 9 9 2
2 0 9
9 1 9 15 13 1 9 2 10 2
31 3 15 9 1 0 13 9 9 2 16 9 9 2 1 9 9 2 9 2 2 9 7 9 9 2 9 9 9 13 0 2
7 13 3 9 2 5 9 2
6 0 9 12 2 2 2
6 0 9 12 2 2 2
6 0 9 12 2 2 2
6 0 9 12 2 2 2
6 0 9 12 2 2 2
4 9 0 9 2
20 0 9 13 9 0 9 7 0 9 2 0 9 13 9 0 9 7 0 9 2
4 9 0 9 2
13 16 4 13 0 9 13 2 13 9 13 1 9 2
11 3 2 0 9 13 10 9 1 0 9 2
41 16 0 9 7 13 3 9 13 15 1 9 12 2 12 2 12 2 12 2 12 2 12 7 12 2 13 15 15 9 0 16 12 7 0 1 12 7 1 12 2 2
36 7 16 13 9 9 3 13 2 13 15 9 13 1 9 9 9 7 9 2 15 4 13 14 0 9 9 9 2 15 13 1 0 9 3 0 2
8 9 2 9 2 7 0 9 2
2 11 11
30 1 9 9 4 9 2 9 2 13 3 1 0 2 3 0 7 0 9 2 10 9 13 0 13 1 0 0 0 9 2
40 1 0 9 7 1 3 0 9 15 13 2 9 2 1 15 0 0 9 2 7 16 15 1 9 13 3 1 9 0 9 2 1 0 0 11 7 1 0 11 2
19 1 10 9 0 0 9 4 1 15 13 9 9 2 0 3 1 9 0 2
13 10 9 13 9 1 9 9 9 9 7 10 9 2
22 13 3 15 0 1 9 9 2 9 2 7 1 2 9 2 2 13 14 0 9 9 2
30 0 9 7 3 9 9 1 11 13 9 9 7 9 2 15 13 1 9 9 9 2 9 2 7 2 9 2 3 3 2
18 1 9 13 2 9 2 0 9 0 9 9 2 0 2 2 9 2 2
15 10 9 4 1 9 0 9 0 9 13 1 12 1 0 2
21 13 15 3 3 2 3 10 2 0 2 9 9 2 9 2 7 2 9 2 13 2
13 9 9 2 9 2 13 0 3 3 12 9 9 2
16 1 0 7 3 2 0 9 15 13 9 2 12 11 2 11 2
27 1 10 9 2 9 7 9 2 2 1 9 0 0 9 7 9 2 15 13 1 0 9 0 7 0 11 2
18 2 12 9 0 9 9 13 9 9 2 15 2 16 13 2 15 13 2
33 13 15 2 16 10 9 13 9 10 9 7 15 3 13 2 13 7 13 9 2 10 9 2 16 13 2 13 10 9 2 2 2 2
15 10 10 9 3 13 11 2 11 9 2 15 13 15 9 2
21 12 1 10 0 9 15 13 9 2 1 15 13 2 16 1 0 9 13 10 9 2
27 16 1 10 9 13 7 13 1 9 9 2 13 2 16 13 7 16 1 9 13 9 2 15 13 10 9 2
23 11 13 10 9 9 2 2 13 10 9 7 9 9 0 9 2 13 9 7 13 1 9 2
22 16 15 13 2 13 1 10 9 2 7 9 4 13 0 9 2 15 15 3 13 9 2
26 16 15 3 0 9 13 2 13 2 16 9 2 10 0 2 15 15 13 2 3 13 10 9 2 2 2
22 9 13 9 2 13 9 13 13 2 10 9 15 13 2 3 3 4 13 2 2 2 2
5 0 9 13 0 2
31 9 7 9 12 2 9 13 0 9 9 1 9 9 1 0 11 2 1 15 15 3 13 7 9 1 11 2 11 7 11 2
38 0 9 7 13 1 0 11 7 7 15 1 0 9 13 9 9 0 2 7 2 2 9 2 2 7 1 15 0 9 2 9 2 7 2 0 9 2 2
2 0 9
50 9 1 9 9 2 9 2 7 2 9 2 2 3 4 13 0 9 12 2 9 2 13 11 2 11 2 11 2 15 13 15 1 0 9 2 9 2 2 0 9 1 9 7 9 2 12 2 12 2 2
22 1 10 9 13 1 9 1 9 9 2 0 9 7 9 0 1 0 9 7 0 9 2
25 10 9 13 1 0 2 2 9 2 2 0 9 9 9 1 0 9 9 0 11 7 1 0 9 2
31 11 13 1 9 2 16 9 13 0 13 1 0 9 16 9 0 1 9 9 7 16 13 15 0 9 9 2 15 9 13 2
24 1 10 9 4 9 13 3 1 9 2 3 9 13 9 9 2 1 15 10 9 13 10 9 2
22 9 10 0 9 2 0 1 0 9 0 9 2 3 13 7 9 9 0 9 7 9 2
33 0 9 1 9 7 9 7 13 0 9 9 11 11 2 9 7 9 2 2 12 2 7 11 11 11 2 0 9 2 2 12 2 2
25 10 9 7 10 9 13 0 2 0 2 9 9 16 0 9 0 9 2 15 13 13 3 10 9 2
14 9 2 0 9 13 7 13 15 1 0 9 0 9 2
27 16 13 0 1 9 2 0 2 9 13 0 9 2 3 13 15 9 2 16 7 10 9 13 9 0 9 2
19 9 2 1 0 9 13 0 3 0 9 9 7 15 13 0 7 0 9 2
19 9 2 9 4 13 1 9 7 3 2 9 13 4 13 1 9 10 9 2
31 9 13 3 0 9 7 13 1 15 0 9 16 1 0 0 9 2 7 2 3 9 1 9 7 9 2 9 0 9 3 2
25 9 2 1 0 13 2 16 15 0 9 0 0 9 15 13 1 15 13 2 16 4 13 3 0 2
11 13 9 9 0 9 2 9 10 9 3 2
36 1 9 10 9 2 16 1 0 0 9 2 1 0 9 2 9 2 15 3 13 9 9 0 9 2 0 2 9 2 7 16 3 4 13 13 2
20 9 2 0 9 4 13 7 9 9 1 9 13 13 7 1 0 7 0 9 2
2 9 9
22 1 0 9 7 9 2 9 2 16 9 15 9 12 2 9 13 7 9 9 10 9 2
41 13 15 7 13 2 16 15 9 0 9 9 1 9 15 13 1 0 9 0 0 0 7 0 9 2 15 13 13 1 10 9 9 2 16 14 1 10 9 9 9 2
28 0 9 1 2 9 2 7 2 9 2 7 9 12 2 7 12 2 9 13 1 9 0 1 0 12 9 9 2
52 9 10 9 3 3 13 2 16 13 1 9 0 1 12 2 7 12 2 9 10 2 9 2 13 1 9 3 2 1 12 2 7 12 2 9 1 2 10 2 9 2 2 7 16 14 2 3 14 1 9 9 2
15 13 15 3 2 1 10 9 1 9 0 9 13 0 9 2
4 9 13 10 2
22 9 2 9 2 16 9 0 9 13 9 2 13 1 9 9 10 1 2 0 9 2 2
20 10 9 13 0 9 2 15 1 9 10 9 13 1 9 2 1 9 9 15 2
14 9 2 9 13 7 13 9 2 15 15 13 10 9 2
15 9 2 9 15 13 1 9 1 9 9 0 9 1 9 2
22 9 2 0 9 10 9 13 9 2 16 9 9 4 13 1 9 1 2 0 9 2 2
31 1 10 9 13 9 2 16 0 9 13 10 9 2 16 12 1 15 2 0 2 2 0 9 2 2 4 13 1 0 9 2
20 9 0 9 2 0 9 2 4 3 3 13 1 9 0 9 2 9 0 9 2
13 9 7 9 9 15 13 1 9 7 9 0 9 2
20 9 2 9 13 1 9 0 0 0 7 0 9 2 3 3 3 13 0 9 2
18 9 2 9 13 1 9 9 9 13 0 9 7 9 1 9 7 9 2
18 7 4 13 9 9 0 9 7 9 7 15 4 1 9 13 0 9 2
11 9 2 9 9 13 1 9 9 7 9 2
24 9 9 0 9 7 9 2 10 9 3 2 13 13 3 1 9 0 9 7 1 9 0 9 2
7 13 15 3 9 0 9 2
20 9 2 9 13 1 9 1 0 9 9 9 2 13 2 1 9 9 0 9 2
25 9 2 9 13 1 9 2 3 15 13 0 9 3 7 3 9 13 10 9 1 9 10 0 9 2
23 10 9 15 9 13 1 10 9 7 13 10 9 7 9 2 15 13 1 10 9 0 9 2
21 1 10 0 9 13 13 7 13 7 3 0 9 15 13 13 9 7 10 0 9 2
23 13 15 7 1 9 7 9 12 2 7 12 2 9 2 10 9 7 9 13 13 3 3 2
29 3 3 15 13 2 16 0 0 9 0 9 4 13 1 0 9 7 16 13 0 9 16 0 9 9 3 3 13 2
3 9 0 9
16 0 9 9 2 0 16 9 2 4 1 0 12 9 13 9 2
13 1 0 9 9 13 0 13 3 11 11 2 11 2
15 9 13 3 2 3 0 0 2 9 2 9 9 7 9 2
47 13 15 2 16 9 12 2 9 2 15 14 3 13 0 9 1 9 7 1 10 9 15 3 13 1 9 9 2 9 7 0 9 2 13 1 10 9 1 0 9 2 1 0 9 1 9 2
7 0 9 13 7 0 9 2
20 9 2 9 2 4 13 1 9 7 13 9 7 9 10 9 2 3 3 9 2
29 13 9 2 16 0 9 0 9 2 9 7 9 2 13 0 9 2 7 10 9 13 15 0 1 0 9 10 9 2
48 1 9 0 9 11 2 15 13 1 9 12 2 7 1 9 12 2 9 1 11 2 13 0 11 10 0 9 9 2 16 1 0 9 9 13 10 9 10 9 0 2 13 3 0 7 0 9 2
18 10 9 2 1 15 15 9 7 9 13 2 4 7 13 1 0 9 2
50 0 9 7 9 9 0 9 7 9 13 1 9 10 9 2 13 7 13 0 9 2 16 3 15 13 2 7 13 1 0 0 9 0 1 9 2 9 2 2 15 13 1 0 9 2 9 2 15 0 2
23 9 11 2 11 2 15 13 3 9 15 0 9 9 2 9 2 3 13 12 9 1 12 2
9 9 2 9 13 0 9 0 9 2
15 9 2 9 1 0 9 7 9 2 15 13 13 0 9 2
13 15 9 0 11 2 11 2 11 2 9 2 12 2
3 0 9 9
26 0 9 0 7 0 9 2 3 3 16 9 0 9 2 7 13 2 16 1 0 9 13 7 9 0 2
15 10 9 13 4 13 9 2 9 9 2 3 10 0 9 2
18 3 0 7 0 9 13 2 16 9 13 13 9 12 2 0 7 0 2
22 16 1 9 12 9 7 9 13 0 12 7 12 0 9 2 3 0 9 13 1 9 2
25 9 0 9 3 13 2 16 9 2 9 2 13 9 1 9 2 0 1 0 9 16 2 9 2 2
41 9 10 9 13 9 2 16 1 0 0 9 2 7 3 1 9 2 9 7 1 0 9 2 1 10 9 2 4 13 9 2 15 13 9 1 0 9 13 10 9 2
34 9 13 1 10 9 2 9 9 7 9 10 9 2 1 9 2 3 13 9 7 9 2 13 15 9 0 2 9 2 9 3 2 2 2
23 3 0 13 9 2 16 0 9 13 10 9 2 1 15 14 12 4 13 1 9 7 9 2
38 15 9 10 9 2 0 9 2 9 2 9 2 13 1 0 9 7 1 9 9 15 3 12 1 15 13 1 0 2 9 2 2 7 2 1 0 9 2
29 9 2 15 13 1 9 2 15 13 9 7 9 0 9 2 9 2 15 15 3 13 1 10 9 2 10 9 13 2
24 1 9 1 2 0 2 9 13 7 13 1 10 9 7 9 2 15 15 13 3 2 1 9 2
28 9 13 0 9 0 9 9 7 9 2 16 7 2 0 2 9 15 1 9 9 13 1 9 0 7 0 9 2
11 9 1 9 3 13 13 1 0 9 9 2
14 13 15 13 16 0 9 9 2 0 1 0 9 9 2
20 13 15 13 16 9 9 0 9 0 0 0 9 7 9 1 2 0 2 9 2
18 13 15 3 13 16 9 0 9 1 9 7 10 9 1 9 2 9 2
57 1 9 9 13 13 2 9 2 1 9 0 9 2 0 9 10 0 9 2 7 15 1 9 1 10 0 9 2 13 2 13 0 2 16 13 9 0 2 0 2 0 7 0 2 3 2 13 9 1 9 9 2 9 3 2 2 2
11 1 9 10 9 13 9 0 15 1 9 2
22 3 16 9 9 2 4 7 9 7 0 9 13 1 9 7 9 9 7 1 0 9 2
12 9 13 3 9 15 9 0 1 0 9 9 2
43 13 4 15 13 2 16 16 9 7 9 1 15 0 13 9 9 0 1 0 7 0 0 9 2 7 9 13 15 7 9 0 9 2 1 9 2 1 0 7 0 0 9 2
13 9 13 3 3 0 9 16 9 2 7 13 0 2
4 9 16 0 9
51 1 9 0 9 1 9 7 1 10 9 1 9 13 13 3 12 0 9 2 15 13 10 9 1 9 2 1 0 9 2 3 2 1 9 9 1 9 7 3 2 7 1 9 1 9 1 9 7 0 9 2
9 0 13 16 0 2 0 16 0 2
19 0 9 13 9 1 9 9 7 9 2 10 9 15 1 10 0 9 13 2
24 13 0 2 16 4 13 9 9 7 3 2 9 7 3 15 1 10 0 9 16 1 9 13 2
30 9 0 10 9 13 0 9 7 3 3 13 1 10 9 2 9 2 3 16 0 0 9 2 3 13 2 1 9 2 2
18 1 9 15 3 13 9 9 2 9 2 9 7 0 9 7 0 9 2
20 9 13 3 9 2 15 13 9 2 7 2 9 15 10 9 1 12 0 9 2
35 1 0 9 13 9 10 2 0 2 9 9 9 0 16 9 2 3 16 3 4 13 9 1 9 2 3 0 1 9 9 2 9 9 2 2
19 9 0 0 9 15 13 1 0 9 9 13 1 9 2 9 2 9 0 2
26 1 10 9 13 10 0 9 2 9 13 0 2 2 13 9 2 9 2 9 1 10 2 0 9 9 2
25 9 13 9 9 7 0 9 2 13 15 13 2 7 2 13 13 10 9 7 9 1 0 9 9 2
13 9 3 1 9 9 3 13 2 7 14 1 9 2
20 10 0 9 15 13 14 1 9 7 13 14 1 9 9 11 2 11 7 11 2
17 4 13 3 3 7 1 9 2 9 7 0 9 1 9 0 9 2
9 9 9 0 13 0 9 0 9 2
21 1 10 0 9 4 9 13 16 9 0 9 2 13 3 3 2 16 4 15 13 2
43 3 1 9 0 9 2 11 2 15 13 10 9 2 2 2 2 2 9 13 9 2 16 4 13 10 9 2 13 15 2 16 4 13 9 0 2 16 9 7 9 15 13 2
16 7 9 15 13 7 13 15 2 13 7 13 15 7 13 9 2
23 13 15 7 13 1 0 9 2 1 0 9 2 1 15 0 2 15 15 13 1 9 2 2
17 3 13 1 9 9 9 1 9 2 9 2 7 3 9 1 15 2
19 0 9 4 13 16 9 9 2 3 15 0 2 16 9 1 2 9 2 2
16 9 0 9 9 13 1 9 9 2 9 2 1 9 0 9 2
31 9 13 14 9 9 0 1 12 2 0 2 9 2 16 0 0 9 4 13 0 2 0 2 9 1 0 2 0 2 9 2
16 1 10 9 4 9 13 15 1 9 1 0 9 9 0 9 2
18 9 9 4 13 7 1 9 1 0 9 7 3 1 9 1 9 0 2
17 9 1 9 9 0 15 13 9 0 9 3 1 9 0 0 9 2
22 3 15 3 3 13 9 9 1 10 9 2 13 2 3 2 9 2 9 0 2 2 2
16 0 9 13 3 9 9 1 9 2 7 3 9 9 1 9 2
11 9 3 13 1 0 9 2 13 15 3 2
14 13 3 9 0 14 1 0 9 2 3 2 9 2 2
13 13 3 15 13 1 12 3 0 0 9 1 9 2
14 12 2 0 2 15 13 0 9 2 13 9 1 9 2
27 0 2 0 2 15 13 9 7 0 9 2 9 1 9 13 7 1 9 2 15 13 9 2 13 0 9 2
36 9 1 15 4 13 9 0 0 9 2 7 2 2 0 2 7 2 0 2 9 2 7 0 9 9 2 7 3 0 9 1 9 16 9 0 2
5 9 0 9 0 9
4 2 0 9 2
2 11 11
15 0 9 7 9 9 13 9 9 1 9 2 15 13 9 2
16 9 1 15 13 1 9 9 9 9 9 1 0 9 0 9 2
17 12 1 3 0 9 13 9 1 9 0 9 0 9 2 9 2 2
19 9 0 9 13 13 9 10 0 9 7 0 9 2 15 15 1 15 13 2
6 15 15 13 0 9 2
23 13 1 0 0 2 0 7 0 9 0 0 9 9 2 3 13 3 16 12 9 9 2 2
16 1 9 9 4 13 12 9 2 1 15 12 15 3 3 13 2
21 3 9 9 1 9 2 7 9 2 0 9 2 0 9 13 3 1 9 0 9 2
19 0 1 9 9 1 9 2 0 1 0 9 0 9 7 12 1 0 9 2
16 0 15 13 13 9 0 9 1 9 0 9 1 9 7 9 2
12 15 4 7 13 1 0 9 0 7 0 9 2
23 1 0 15 13 9 2 10 9 9 2 9 2 1 15 9 13 1 9 2 13 12 9 2
22 13 3 9 9 9 1 9 7 1 9 2 7 7 13 0 10 9 0 3 3 13 2
19 9 15 3 13 1 0 0 9 2 16 13 9 2 0 9 2 0 9 2
10 4 7 13 7 0 7 0 0 9 2
1 13
7 1 0 9 13 9 0 2
13 13 15 3 13 12 9 2 13 2 13 2 13 2
15 10 9 13 0 9 7 10 9 4 13 3 0 9 9 2
22 0 9 4 13 9 1 9 9 2 7 3 15 9 13 1 9 9 9 1 9 12 2
15 3 13 15 9 2 9 0 7 0 9 2 9 7 9 2
24 0 9 13 9 9 9 9 0 9 1 0 9 2 1 9 2 15 13 9 7 9 0 9 2
10 13 15 9 3 1 9 0 7 0 2
21 16 0 9 15 13 9 2 0 9 2 10 9 7 1 0 9 9 7 0 9 2
31 9 9 13 1 0 9 13 2 15 9 13 10 9 1 0 7 0 9 10 9 2 15 13 9 9 1 0 9 9 9 2
39 9 9 0 9 13 1 9 9 0 9 7 13 15 1 0 9 9 1 10 9 14 1 9 12 9 2 13 9 12 2 2 2 2 2 2 2 12 2 2
23 1 0 9 0 9 9 1 0 9 15 13 3 13 1 9 2 15 4 10 0 9 13 2
2 0 9
15 9 0 9 0 9 1 9 1 9 4 13 16 0 9 2
22 4 13 1 9 9 0 9 1 3 0 2 0 2 0 7 3 0 0 7 0 9 2
16 0 9 13 0 2 9 9 2 15 13 3 0 9 10 9 2
35 0 9 13 9 2 9 2 9 7 9 2 10 9 13 0 9 1 10 9 2 0 9 2 14 1 9 9 2 0 9 1 0 9 2 2
18 0 9 13 0 9 0 9 2 3 0 2 15 13 13 0 9 9 2
50 0 7 0 0 9 13 0 2 0 7 0 9 2 0 2 0 2 0 2 2 10 9 13 13 0 9 9 2 15 13 1 0 9 0 9 15 2 16 13 13 9 7 13 15 1 9 1 0 9 2
19 15 0 9 15 13 1 0 9 2 7 0 9 9 0 9 13 0 9 2
35 15 13 13 9 9 2 13 13 0 0 9 2 9 0 1 0 9 2 13 13 3 0 2 16 4 15 13 0 3 13 7 13 2 3 2
19 1 0 9 13 15 1 15 13 0 9 9 1 15 0 7 0 9 9 2
17 0 0 9 13 13 3 2 16 9 9 13 13 0 9 9 9 2
23 1 9 15 13 2 16 16 10 9 13 0 9 2 16 4 13 2 10 9 13 9 0 2
28 3 2 13 2 14 9 13 3 3 2 13 0 2 0 9 2 15 15 0 9 0 9 13 10 0 0 9 2
21 3 4 15 13 1 9 0 9 2 3 15 13 1 9 0 1 9 0 9 9 2
21 1 1 9 0 9 13 0 9 9 0 9 0 9 9 2 15 13 1 9 13 2
12 9 0 9 13 0 9 0 1 9 0 9 2
21 15 4 13 3 0 9 0 1 9 9 9 2 15 1 9 7 10 9 13 13 2
38 13 15 9 2 15 13 2 9 2 9 2 16 13 9 2 0 9 2 0 0 9 9 7 9 2 0 2 0 7 0 9 9 2 0 9 2 0 2
12 0 9 9 9 13 9 0 9 1 0 9 2
53 15 4 13 1 9 0 9 1 0 9 7 1 9 0 9 2 16 13 9 9 7 9 1 0 9 2 9 0 9 2 9 2 2 9 9 1 9 1 0 9 2 3 2 1 0 0 9 2 11 1 11 2 2
28 0 9 0 9 13 0 9 0 0 9 2 15 15 13 1 9 7 0 9 9 2 1 15 13 4 9 13 2
27 0 0 9 13 3 0 9 0 7 0 9 2 9 2 15 13 13 1 9 9 1 9 7 1 9 9 2
31 1 0 9 13 9 9 2 9 0 9 2 9 0 9 2 9 9 1 9 0 3 1 9 2 9 9 1 10 9 3 2
29 13 15 1 15 0 9 2 15 13 9 0 0 9 7 13 15 1 15 2 15 0 9 13 9 2 0 9 2 2
6 15 13 0 9 9 2
22 3 15 0 9 9 13 9 9 1 9 9 1 9 2 15 13 1 0 9 0 9 2
36 13 15 0 9 2 13 15 9 9 9 2 13 15 9 9 0 0 9 2 9 2 9 2 9 2 7 3 13 15 9 1 9 9 15 9 2
10 9 9 9 13 3 0 9 0 9 2
34 15 0 9 13 13 0 0 0 9 2 13 15 3 0 0 0 9 12 9 2 15 13 9 1 9 13 2 0 9 13 3 0 2 2
29 9 15 7 13 1 0 9 9 2 15 13 10 9 7 1 0 9 15 13 3 1 12 1 12 2 9 1 9 2
12 15 15 13 9 1 0 9 9 1 0 9 2
45 1 0 0 9 0 9 12 5 9 2 9 2 12 13 1 0 1 9 7 13 0 1 9 0 1 0 9 7 1 9 9 7 13 3 12 5 9 1 0 9 0 1 0 9 2
9 13 3 9 1 0 9 0 9 2
10 1 0 9 4 13 0 9 0 9 2
18 15 2 15 13 0 9 9 1 0 9 2 13 4 13 1 0 9 2
17 15 13 9 9 0 1 9 0 9 7 9 1 11 7 1 11 2
23 0 9 1 0 9 7 0 9 3 4 13 1 0 0 9 12 7 12 9 1 9 9 2
6 10 9 3 4 13 2
9 10 9 13 1 9 1 0 9 2
46 0 9 9 13 13 0 1 12 2 12 9 2 15 13 9 2 1 15 13 1 0 9 13 0 9 2 9 2 0 9 2 7 1 15 13 0 13 7 13 0 0 9 0 0 9 2
27 16 13 9 0 9 1 9 9 9 2 13 15 1 9 0 9 9 1 15 2 7 3 1 9 0 9 2
51 7 4 9 1 0 9 13 1 9 2 7 15 13 0 9 1 0 7 0 9 2 9 9 7 15 7 9 9 0 9 1 9 2 7 3 9 9 9 0 9 1 9 2 16 4 9 1 9 9 13 2
19 13 13 2 16 9 0 1 0 9 0 9 4 1 10 9 13 1 9 2
35 15 15 9 13 3 1 15 0 0 9 2 1 0 9 2 3 4 13 9 1 15 0 2 15 1 15 3 13 2 13 15 3 1 9 2
9 13 3 0 13 9 0 9 9 2
52 1 0 9 2 7 0 7 0 2 13 2 13 10 9 2 16 4 9 9 9 13 3 0 2 3 13 0 2 2 15 13 1 9 9 2 7 0 7 3 0 2 2 13 9 2 15 13 3 0 2 2 2
26 4 3 13 2 16 1 9 0 9 13 9 9 7 9 0 16 13 9 9 1 9 9 9 1 9 2
14 7 15 13 9 2 15 15 3 10 0 9 13 13 2
26 1 0 9 13 3 13 9 1 9 9 0 9 1 15 2 16 3 13 9 1 0 9 7 0 9 2
14 13 2 7 9 15 13 1 15 2 3 15 7 13 2
5 0 9 13 9 2
28 9 0 9 4 13 3 3 16 12 9 9 7 3 3 3 15 13 2 16 1 10 9 13 3 0 0 9 2
18 15 3 13 7 1 0 0 9 2 16 0 9 9 0 9 13 9 2
37 1 9 15 2 16 0 9 13 13 0 7 1 9 9 2 9 3 3 13 15 0 9 9 9 0 9 7 13 9 2 15 4 10 9 3 13 2
30 3 2 1 11 1 12 9 0 0 9 1 0 9 11 13 9 0 9 1 11 2 15 13 15 9 1 9 0 9 2
25 15 3 7 13 13 2 7 10 9 13 3 13 2 16 15 1 10 9 9 9 0 10 9 13 2
12 0 9 13 0 9 13 1 12 7 12 9 2
28 15 2 16 10 9 7 9 4 13 1 11 1 12 9 2 13 9 10 9 2 7 9 0 9 1 0 9 2
39 0 0 9 13 9 2 16 3 13 1 9 0 9 13 9 2 7 0 9 13 3 13 2 13 9 10 9 1 9 2 12 1 15 13 1 0 11 2 2
30 3 13 0 2 16 1 0 9 9 13 1 0 9 9 7 9 9 2 15 13 9 0 1 0 9 9 7 9 9 2
30 7 3 0 9 2 0 1 0 2 13 2 16 3 4 13 1 15 2 16 13 0 13 0 9 2 7 15 3 13 2
17 1 0 9 13 3 0 2 16 7 12 1 12 9 13 0 9 2
7 13 15 3 3 9 0 2
13 0 9 9 16 0 2 7 0 13 0 0 9 2
31 13 4 15 13 2 16 9 9 1 0 9 0 9 0 9 4 13 1 9 7 16 9 10 0 9 13 1 10 9 9 2
18 13 15 10 9 0 2 7 0 9 13 15 2 15 0 9 13 3 2
22 3 13 3 0 9 2 15 13 12 1 0 9 9 2 9 13 15 3 1 0 9 2
3 14 2 13
13 9 9 2 1 9 15 13 1 0 9 0 9 2
26 16 13 1 12 2 3 2 13 15 3 1 10 0 9 1 9 11 2 9 2 12 2 12 7 12 2
27 13 4 9 7 9 7 13 4 7 3 9 13 15 1 9 2 13 3 1 15 2 3 15 1 15 13 2
6 13 15 1 0 9 2
3 9 0 2
4 9 9 0 9
7 9 2 0 9 2 0 9
13 2 9 9 1 9 12 2 12 9 1 9 1 9
4 2 9 1 9
11 2 9 7 9 9 1 9 1 9 12 9
7 2 9 1 9 1 0 9
6 2 9 9 1 0 9
6 2 9 9 2 3 2
4 2 9 1 9
3 2 0 9
6 9 1 7 1 0 9
2 1 2
7 2 0 0 0 9 1 9
15 2 0 9 9 1 0 9 2 7 1 0 9 1 0 9
8 2 9 9 0 9 0 1 9
16 2 9 9 4 13 1 11 2 3 1 9 1 9 1 0 9
5 2 0 9 1 9
15 2 9 13 3 1 0 9 2 7 3 1 9 0 1 9
19 2 12 2 12 5 9 9 1 0 9 2 12 2 12 5 1 0 9 2
2 1 2
22 2 0 9 13 1 10 0 9 13 2 7 0 9 13 0 9 9 2 3 9 7 9
7 2 0 9 1 9 15 13
4 2 3 0 9
30 2 9 13 0 9 0 9 2 1 11 12 9 9 1 9 2 12 2 7 2 12 0 9 2 9 14 12 9 12 2
6 2 13 1 9 9 9
9 2 9 0 9 13 9 1 0 9
22 1 0 9 13 12 9 2 11 2 11 2 11 2 11 7 11 2 0 1 0 9 2
12 15 12 9 13 12 5 9 0 9 0 9 2
6 9 2 9 2 0 9
13 2 9 9 1 9 12 2 12 9 1 9 1 9
8 2 9 1 9 7 1 0 9
4 1 9 3 0
8 2 9 9 1 9 7 0 9
2 2 9
13 2 9 0 0 9 1 9 10 9 12 9 1 9
9 2 9 0 9 2 15 13 0 9
10 2 0 9 9 1 12 5 9 0 9
4 2 9 0 9
5 9 1 7 1 9
2 1 2
4 2 3 0 9
28 2 1 9 9 13 0 9 1 9 1 9 9 1 0 9 2 1 9 11 7 11 0 14 1 9 2 12 2
16 2 9 0 9 13 9 7 13 9 1 9 0 9 1 0 9
15 2 9 2 1 9 2 13 10 0 9 1 9 9 0 9
9 2 0 9 13 0 9 1 0 9
14 2 9 0 9 2 12 5 1 9 7 12 5 1 9
6 2 9 1 0 9 9
2 1 2
11 2 9 1 9 13 0 13 1 0 9 2
18 1 9 15 3 13 1 9 9 1 0 9 2 7 7 1 0 9 9
7 2 9 9 13 13 0 9
9 2 9 1 9 9 13 3 3 0
15 2 1 0 9 13 9 9 1 9 0 9 1 9 2 12
13 2 9 13 9 1 9 1 0 9 7 3 15 13
7 9 12 12 12 12 12 12
7 9 2 9 0 9 1 11
15 12 12 0 9 1 9 12 13 1 11 2 0 1 11 2
18 13 13 9 0 9 1 1 0 9 9 1 9 9 12 7 9 12 2
11 9 0 1 9 0 9 9 13 1 9 2
17 7 1 0 9 13 1 9 2 12 9 0 9 3 12 9 9 2
2 11 11
6 9 1 12 9 9 9
6 1 9 9 1 9 2
22 1 9 2 15 13 0 0 9 9 2 13 15 2 16 0 2 0 9 2 9 0 2
36 9 1 9 0 11 13 9 2 16 10 9 0 1 9 13 3 3 3 0 9 9 0 2 15 15 7 3 3 13 16 9 3 0 7 0 2
22 9 9 0 13 15 4 3 3 13 2 16 13 1 9 2 16 4 13 0 9 9 2
18 7 9 0 9 0 1 9 13 3 0 16 9 9 0 2 0 3 2
45 15 13 14 0 7 3 3 0 9 9 2 7 9 15 13 15 3 3 7 13 15 3 1 9 2 0 1 10 9 2 15 7 1 9 9 13 1 9 0 9 1 9 7 9 2
34 9 9 0 1 9 2 15 3 1 0 9 13 0 2 13 15 1 0 9 0 9 10 9 2 16 3 3 0 9 0 13 9 9 2
28 9 0 2 0 0 9 0 2 13 0 9 9 7 1 10 9 2 1 15 1 9 0 13 7 9 2 2 2
9 9 12 2 9 12 2 9 2 12
3 9 9 2
12 9 0 13 15 3 10 9 0 9 1 9 2
19 1 0 9 2 13 0 9 2 0 2 11 0 2 2 13 10 0 9 2
31 9 0 13 15 9 2 7 9 2 15 13 13 2 13 15 1 9 10 2 16 15 3 0 9 16 0 3 1 15 13 2
29 9 0 2 9 9 2 13 15 3 0 9 2 7 9 0 2 0 0 9 9 2 13 1 9 2 13 0 9 2
21 0 9 9 0 7 2 14 9 2 9 0 2 13 15 2 7 13 3 10 9 2
9 9 12 2 9 12 2 9 2 12
4 9 9 0 9
2 11 11
2 11 0
13 0 9 0 9 13 7 3 1 9 16 0 0 2
21 16 0 9 13 3 1 9 9 2 0 9 0 0 0 9 3 13 15 9 0 2
8 9 9 13 1 15 9 0 2
31 1 10 0 2 15 1 9 13 9 7 13 0 7 13 2 13 0 9 2 15 9 13 3 0 2 3 2 0 0 9 2
23 13 7 1 15 2 16 4 13 0 2 0 9 1 9 9 2 7 16 4 13 0 9 2
11 0 7 0 9 15 13 1 15 0 9 2
12 0 0 9 3 13 0 0 9 1 0 9 2
18 3 13 2 10 9 13 9 13 2 16 10 13 9 1 0 9 9 2
15 3 16 9 0 0 9 13 0 9 0 9 1 10 9 2
19 13 2 16 0 9 13 13 9 7 1 3 0 7 0 0 9 0 9 2
4 9 0 9 2
18 0 9 4 13 3 1 3 0 9 2 15 13 9 14 1 9 9 2
8 13 0 9 0 9 0 9 2
9 9 10 9 0 9 13 0 9 2
19 15 13 3 11 2 11 2 7 9 9 13 3 9 9 7 0 0 9 2
3 0 9 9
20 1 9 15 13 10 9 2 15 15 3 13 0 9 2 9 9 7 9 9 2
14 0 13 0 9 11 2 15 13 12 9 1 0 9 2
17 9 11 7 11 13 12 9 2 16 11 13 0 7 11 0 9 2
14 1 0 9 13 0 9 11 2 0 3 9 12 11 2
12 0 0 9 15 13 1 0 9 7 0 9 2
8 0 9 13 0 9 7 9 2
12 0 9 13 9 1 9 2 3 16 0 9 2
14 1 9 2 0 1 0 9 1 9 2 4 13 9 2
10 9 4 13 1 9 1 0 9 9 2
15 0 9 13 0 9 1 0 7 13 15 1 0 9 9 2
17 3 13 10 9 9 2 9 2 9 7 9 2 13 9 12 2 2
24 1 0 9 4 13 9 9 2 1 9 4 13 9 0 9 2 9 9 4 13 9 0 9 2
13 0 9 9 2 9 7 9 15 13 0 0 9 2
14 13 1 9 9 0 9 7 9 0 9 1 0 9 2
10 9 7 0 9 13 0 9 0 9 2
17 9 9 7 9 15 13 9 1 0 0 9 13 15 0 0 9 2
22 1 9 4 0 9 3 13 1 0 0 9 2 16 4 13 4 3 13 1 0 9 2
8 3 13 13 7 13 1 9 2
6 0 9 13 0 9 2
3 0 9 2
8 0 9 9 13 13 9 9 2
18 0 9 2 0 0 0 9 2 13 3 0 16 9 1 9 0 9 2
7 3 13 9 3 0 9 2
8 9 15 13 1 9 7 9 2
9 15 13 0 9 9 2 9 2 2
12 9 7 9 4 13 1 3 0 9 10 9 2
12 9 12 9 13 3 0 7 13 15 1 9 2
14 9 15 1 9 13 1 0 9 2 15 15 13 9 2
9 15 3 13 0 9 7 0 9 2
20 4 1 9 9 13 1 2 0 9 2 1 9 7 1 10 9 13 9 9 2
19 0 9 13 15 9 1 9 9 2 15 9 13 9 1 0 9 1 9 2
17 1 9 0 9 15 13 0 2 0 9 2 0 13 0 9 9 2
13 3 0 9 13 0 9 1 0 9 2 0 9 2
20 9 9 7 9 9 2 9 2 9 3 2 13 0 0 9 0 1 9 9 2
28 1 10 0 9 15 13 0 9 2 9 1 9 2 9 2 9 2 9 9 2 9 7 9 9 3 2 2 2
13 0 13 7 0 9 2 9 0 9 9 2 9 2
29 9 0 9 15 13 1 12 9 2 9 1 9 1 9 2 0 0 2 7 9 1 9 1 9 2 0 0 2 2
14 0 9 13 0 1 10 9 2 0 1 10 9 9 2
20 3 13 0 1 0 9 1 9 7 3 3 3 9 13 2 15 13 10 9 2
14 0 7 0 9 0 9 13 0 9 9 1 0 9 2
12 15 13 7 0 13 2 14 16 13 0 9 2
8 9 0 9 1 0 7 0 9
19 0 9 0 9 13 3 13 1 12 9 1 0 9 9 9 1 0 9 2
15 9 0 9 13 1 9 9 1 0 0 9 1 0 9 2
16 0 9 1 0 9 4 13 1 0 9 1 9 0 0 9 2
26 9 0 9 13 1 0 9 0 0 9 2 3 2 9 2 9 9 2 7 1 15 13 0 0 9 2
24 1 0 9 0 9 15 13 9 9 2 15 13 13 1 12 9 3 1 0 2 7 0 9 2
16 1 0 9 1 12 0 9 15 9 13 3 3 9 7 9 2
15 0 9 9 0 9 13 1 0 9 1 0 9 9 9 2
17 12 9 15 1 9 9 13 2 7 3 3 0 9 13 15 0 2
8 10 0 9 10 9 13 3 2
25 16 0 9 13 0 0 9 2 13 4 15 1 9 0 9 0 9 0 1 0 9 3 0 9 2
11 0 9 1 0 9 7 10 9 1 0 9
14 0 9 13 16 9 9 1 9 12 9 7 12 9 2
12 14 1 0 9 1 11 9 13 9 9 0 2
22 9 9 7 0 9 2 0 0 0 9 2 13 0 9 1 0 9 1 9 0 9 2
27 3 1 11 9 15 0 9 9 0 9 7 0 9 13 1 0 7 0 9 1 0 9 7 9 0 9 2
4 9 9 0 9
11 1 0 9 13 0 9 9 12 0 9 2
18 0 15 13 0 9 2 16 0 9 13 3 0 9 9 1 0 9 2
14 0 9 13 9 1 9 9 7 0 9 13 10 9 2
12 9 9 1 0 9 13 9 1 0 9 9 2
19 0 9 0 9 2 0 9 2 13 9 9 1 9 9 1 0 0 9 2
11 9 1 9 0 9 15 13 1 9 9 2
22 16 9 9 9 9 4 13 9 9 2 13 9 10 9 1 9 3 12 2 12 9 2
15 12 10 9 2 0 7 0 2 15 1 0 9 9 13 2
17 1 9 0 9 13 0 3 9 2 0 1 0 9 1 9 9 2
7 9 15 13 1 9 9 2
36 16 0 9 0 9 0 9 13 3 3 0 2 13 1 9 1 9 1 0 9 0 9 2 2 13 9 9 1 9 1 9 7 1 9 9 2
12 1 0 9 15 1 9 9 13 3 0 9 2
11 9 9 0 0 9 13 0 1 9 9 2
15 1 9 9 13 9 9 2 7 3 15 13 7 10 9 2
20 13 7 0 13 2 16 9 13 1 9 12 9 9 9 2 7 9 9 9 2
4 9 9 0 9
10 9 9 0 9 15 13 16 9 9 2
16 9 9 4 13 16 9 9 1 9 0 9 7 9 10 9 2
18 0 0 9 13 0 0 9 0 9 2 15 13 13 1 0 9 9 2
5 10 0 9 13 2
11 13 14 9 10 9 2 15 13 9 9 2
11 0 9 13 0 0 9 2 0 12 9 2
16 9 1 0 9 4 13 1 0 0 9 0 9 0 0 9 2
5 9 9 1 0 9
30 0 9 13 1 0 9 1 9 1 0 9 3 0 0 9 2 1 10 9 1 3 12 9 2 13 9 2 12 2 2
19 9 9 13 1 9 10 9 3 3 2 3 16 1 9 0 9 0 9 2
10 13 0 9 2 7 9 13 3 0 2
10 7 13 4 1 0 9 13 0 9 2
17 9 9 13 14 1 9 0 9 2 7 3 1 9 0 0 9 2
5 0 9 7 0 9
11 9 1 9 9 1 9 9 13 10 9 2
11 1 9 9 0 9 9 13 13 0 9 2
19 1 9 0 9 13 0 0 0 9 0 9 0 9 2 3 12 5 2 2
13 9 0 9 0 9 13 0 7 0 9 0 9 2
17 0 1 9 13 0 0 9 1 9 9 16 9 0 1 0 9 2
19 13 15 1 9 1 9 11 2 3 0 9 13 9 0 3 3 1 9 2
12 1 0 9 0 9 13 0 9 0 9 13 2
2 0 9
12 3 9 9 9 1 0 9 13 1 9 9 2
17 9 15 1 0 9 9 13 0 9 7 13 15 1 9 0 9 2
12 7 1 9 9 13 1 9 13 9 0 9 2
20 9 9 9 0 1 9 9 2 0 9 2 13 7 3 0 16 1 3 0 2
16 9 9 1 9 13 9 2 7 7 1 9 13 0 0 9 2
24 13 0 9 9 2 7 7 9 2 15 15 3 13 13 7 13 0 2 13 1 0 9 9 2
4 9 7 0 9
13 9 13 14 1 9 9 2 7 3 1 0 9 2
17 9 4 13 3 9 2 7 7 1 3 0 13 9 9 0 9 2
2 9 9
22 1 0 9 0 9 4 13 9 9 2 0 0 9 9 2 9 9 2 1 0 9 2
11 0 9 13 0 9 1 11 7 1 9 2
16 15 3 13 2 15 13 9 0 9 2 13 13 14 15 0 2
14 1 9 0 0 9 13 9 0 9 2 7 0 9 2
15 1 0 9 9 13 9 16 9 2 9 2 9 7 3 2
13 10 1 3 0 9 0 9 13 0 1 3 0 2
26 3 1 9 15 13 13 0 9 9 2 3 2 9 2 9 9 2 9 2 0 7 0 9 2 9 2
11 1 9 9 13 0 9 16 9 1 9 2
18 3 10 0 13 0 13 10 9 1 9 2 0 2 9 2 0 9 2
21 10 0 9 13 9 1 0 9 1 0 9 2 15 15 13 1 9 1 9 2 2
10 0 9 13 9 0 9 1 0 9 2
11 12 3 13 0 9 2 9 2 0 9 2
18 13 15 3 2 16 9 13 0 13 7 3 13 3 0 9 1 9 2
22 16 15 13 13 14 12 9 9 2 15 13 13 2 13 9 0 9 1 0 0 9 2
9 3 4 9 13 3 1 0 9 2
17 1 9 1 9 15 13 0 9 2 3 1 9 1 9 0 9 2
28 0 9 9 0 9 13 0 13 3 3 2 7 9 2 16 0 0 9 3 13 0 0 9 2 15 3 13 2
18 7 1 9 15 13 10 0 9 2 7 3 9 1 3 0 0 9 2
11 0 9 3 3 13 0 0 9 9 9 2
23 9 0 7 13 2 16 15 13 0 9 2 1 15 15 1 0 9 10 9 0 9 13 2
7 1 9 15 13 0 9 2
9 1 3 0 15 15 1 9 13 2
7 9 13 1 10 0 9 2
1 9
15 11 2 11 7 9 2 2 0 9 9 0 9 1 9 2
3 0 0 11
14 0 9 13 14 9 2 7 7 9 2 9 7 3 9
2 11 11
19 0 9 13 0 0 9 9 11 1 0 9 1 9 2 0 0 9 3 2
16 3 9 13 3 0 9 9 2 10 9 2 9 7 9 9 2
7 15 15 3 0 9 13 2
2 9 9
18 1 0 9 0 9 7 9 1 9 9 13 0 9 3 0 10 9 2
39 0 9 13 15 2 1 3 0 7 0 9 0 9 1 9 9 13 9 2 10 0 9 13 13 9 0 3 1 0 9 7 13 15 13 0 9 0 9 2
26 9 2 13 9 0 9 2 13 0 2 13 7 13 0 9 9 7 9 2 9 9 7 9 0 9 2
29 9 2 3 0 0 9 9 9 2 0 2 9 0 9 0 9 2 0 9 1 0 9 1 0 2 3 0 9 2
2 9 9
38 0 9 10 9 2 3 0 2 15 13 9 2 12 7 13 15 9 2 11 11 2 11 1 9 11 11 1 11 2 11 2 1 9 11 11 11 11 2
9 9 13 3 0 16 0 11 11 2
17 1 0 9 15 13 2 1 9 10 9 2 1 9 0 11 11 2
24 1 10 9 13 9 16 2 0 2 0 2 14 2 0 9 2 2 0 9 1 9 13 9 2
31 0 0 9 13 9 9 2 9 1 0 9 2 2 1 15 13 1 12 9 15 0 9 9 2 15 13 11 1 10 9 2
27 10 9 13 12 2 10 9 13 9 10 9 16 0 0 11 2 2 11 11 2 0 11 7 11 0 11 2
16 3 13 9 9 12 9 0 0 9 2 15 4 3 13 9 2
16 9 0 9 1 0 9 4 13 1 9 16 10 9 1 9 2
29 9 13 1 10 9 0 9 2 9 1 11 2 2 15 13 12 9 2 0 9 4 13 12 0 9 1 0 9 2
13 15 13 1 9 0 9 2 3 3 15 13 9 2
8 1 0 0 9 13 9 9 2
2 0 9
28 9 0 9 4 13 3 12 9 2 13 13 1 9 0 9 2 15 13 3 1 9 9 2 1 9 9 2 2
20 15 3 0 13 13 0 9 3 9 9 2 15 15 3 13 0 7 0 9 2
33 9 9 2 15 15 3 13 2 13 7 13 3 9 0 9 2 7 13 1 9 0 9 1 0 9 7 13 15 0 9 1 9 2
31 13 2 14 9 13 2 4 13 9 9 2 15 3 13 1 9 7 9 0 9 2 9 9 1 9 7 9 7 9 0 2
23 1 9 0 9 13 9 0 9 10 9 7 13 2 16 15 13 13 0 9 1 0 9 2
22 16 13 0 9 2 4 13 9 0 9 7 0 9 4 13 9 1 10 9 1 9 2
25 1 0 9 15 9 13 3 1 0 0 9 1 9 12 9 0 15 1 9 0 11 7 0 11 2
15 9 1 0 9 15 13 13 0 9 7 3 1 12 9 2
33 1 0 9 15 13 3 12 9 2 0 0 9 9 7 9 1 0 9 7 0 9 1 0 9 7 10 9 2 16 9 7 9 2
4 9 7 9 9
38 16 4 9 9 13 2 13 3 1 9 9 7 15 9 9 2 16 4 13 9 0 9 1 9 3 3 13 9 9 7 13 15 1 10 0 0 9 2
27 0 9 13 2 16 15 9 13 0 2 2 14 0 9 2 2 7 16 15 9 13 3 3 13 10 9 2
44 1 9 9 4 13 10 0 9 2 3 1 9 9 15 15 9 9 13 2 16 9 0 0 9 1 9 9 4 13 1 10 10 0 9 7 16 1 9 9 15 13 0 9 2
18 15 9 15 13 0 9 9 0 1 9 13 7 13 3 1 0 9 2
32 1 9 9 3 0 1 9 15 13 9 1 9 0 9 2 9 9 0 1 10 9 7 9 9 0 2 3 7 3 0 9 2
21 9 13 3 0 0 9 1 0 9 7 13 1 15 0 9 4 13 7 0 9 2
9 9 15 13 3 1 9 1 9 2
20 9 4 13 9 2 9 4 3 13 3 16 9 9 7 16 9 1 0 9 2
19 1 0 0 9 3 13 0 9 1 9 2 15 15 3 13 3 1 9 2
38 9 13 0 2 0 3 0 9 2 7 3 15 3 13 1 0 9 12 9 2 15 15 3 3 3 13 2 7 3 3 13 0 9 11 1 0 9 2
32 9 9 0 9 4 13 1 3 12 2 9 0 13 9 2 9 3 2 13 9 2 9 1 9 9 1 0 12 9 2 2 2
23 15 2 1 15 15 13 2 1 10 9 13 15 3 16 9 0 2 2 4 13 16 9 2
14 0 0 9 13 0 7 0 1 15 9 1 0 0 2
45 13 15 2 16 15 9 13 1 9 1 0 9 10 9 2 4 3 13 1 12 9 1 0 9 7 3 15 13 2 3 16 13 0 9 3 2 16 4 15 13 7 13 13 9 2
63 9 7 9 1 0 9 9 13 0 9 1 9 0 1 15 0 3 15 0 9 1 0 9 0 3 7 3 0 9 1 9 2 0 9 1 9 9 13 10 9 12 9 2 13 13 3 1 9 7 9 2 7 3 3 15 0 9 13 3 14 1 9 2
17 9 9 0 9 9 13 3 13 1 0 9 1 12 0 1 0 2
17 15 0 15 13 15 0 9 7 9 1 9 13 1 10 9 0 2
5 15 13 1 9 2
35 9 1 0 9 13 7 0 9 2 3 1 9 2 1 15 9 9 1 9 3 13 9 2 3 13 1 0 9 13 2 16 4 13 0 2
69 9 13 14 0 9 0 2 1 9 15 3 13 1 9 2 15 15 1 9 13 3 14 1 12 9 2 2 7 13 7 0 7 0 9 2 0 9 2 1 15 3 13 2 0 9 13 14 9 2 7 7 9 2 9 7 3 9 2 16 0 9 2 15 13 9 0 1 9 2
3 9 1 9
9 1 15 15 13 1 9 7 1 15
3 9 11 11
23 1 9 9 0 9 4 3 3 13 9 11 11 2 3 9 3 0 9 11 11 2 11 2
16 13 1 9 2 16 15 10 0 9 13 9 10 9 0 9 2
17 7 16 0 9 11 2 9 11 13 0 13 1 2 9 2 2 2
26 10 9 1 9 2 12 13 9 1 0 9 3 1 9 0 9 2 13 9 12 2 12 2 12 2 2
14 1 0 9 1 0 11 4 13 3 11 0 9 9 2
18 13 15 9 0 9 11 11 1 10 9 1 0 0 9 1 10 9 2
4 9 10 9 2
9 0 9 2 3 13 9 3 2 2
16 1 11 0 9 13 3 0 9 9 2 9 1 9 2 2 2
17 9 1 9 13 9 11 11 2 3 3 1 0 12 9 9 9 2
31 7 1 10 9 4 13 13 1 10 9 2 1 0 9 9 2 15 15 13 13 9 2 13 9 0 9 2 7 15 0 2
12 13 3 3 0 2 16 0 9 9 9 9 2
16 9 1 9 13 11 11 1 9 0 2 9 2 2 0 9 2
25 13 0 13 2 16 1 9 9 15 1 11 13 1 9 3 10 9 2 0 1 9 0 9 3 2
13 11 13 0 7 12 1 9 13 10 9 1 11 2
19 9 11 11 1 9 15 13 11 11 2 9 1 12 0 9 0 9 9 2
15 1 9 12 2 12 13 12 9 2 3 0 12 9 12 2
7 13 4 7 9 1 9 2
20 13 15 15 9 0 0 9 2 15 1 9 9 1 12 9 15 3 2 13 2
12 9 15 3 4 13 1 0 0 9 1 9 2
4 0 9 1 9
16 9 3 13 3 9 7 9 1 9 0 9 1 0 9 11 2
35 11 11 11 1 0 9 7 11 11 1 0 9 1 11 13 9 2 15 4 13 9 1 11 11 12 2 7 12 2 9 7 12 2 9 2
18 13 1 9 2 12 9 13 1 0 9 0 9 3 1 9 2 12 2
15 0 9 13 9 12 9 7 10 9 13 3 9 9 11 2
17 0 9 11 11 3 13 9 16 0 1 9 1 9 9 0 9 2
11 0 9 13 9 1 9 0 0 9 9 2
27 9 13 13 2 16 1 0 2 0 9 9 1 0 9 1 9 13 3 0 2 0 9 3 1 9 11 2
12 3 4 13 13 0 9 2 1 15 7 0 2
10 7 1 9 3 13 13 0 0 9 2
32 11 11 1 0 9 13 9 0 9 2 12 3 2 7 13 2 16 3 13 0 9 7 9 2 15 15 3 13 1 0 9 2
17 9 0 9 7 9 2 9 2 9 7 9 9 12 13 3 0 2
23 1 0 9 9 15 11 13 13 7 9 1 9 0 2 15 13 1 0 9 0 0 9 2
18 9 13 14 0 9 11 13 14 14 9 7 13 7 3 3 10 9 2
31 9 0 9 3 13 10 0 9 2 15 13 3 10 0 9 2 3 2 0 2 0 9 2 2 7 3 13 0 9 9 2
6 15 15 13 13 13 2
6 0 9 13 3 9 2
24 16 13 9 11 0 9 0 9 2 13 1 9 2 15 13 3 13 16 13 15 1 9 9 2
17 7 15 13 1 10 0 9 10 0 9 2 3 0 9 13 3 2
20 7 15 10 9 13 1 0 9 3 3 1 9 7 4 10 0 9 13 3 2
5 3 9 1 9 2
25 12 0 9 1 0 9 9 2 11 11 7 11 11 13 0 9 2 15 13 9 1 9 2 9 2
12 13 15 1 9 1 9 0 9 1 0 9 2
11 9 4 13 1 9 9 2 9 7 9 2
23 0 9 15 9 3 13 2 16 9 13 3 0 9 2 16 4 13 13 1 9 9 9 2
8 9 13 1 11 16 0 9 2
18 1 0 9 13 3 9 1 9 9 2 13 0 0 0 9 1 11 2
21 10 9 13 1 10 9 13 16 9 2 7 13 4 13 3 0 0 9 7 9 2
22 3 2 9 2 12 4 1 11 13 1 12 9 9 9 1 9 9 9 0 1 9 2
10 9 9 9 4 3 13 1 12 5 2
3 13 15 2
6 1 9 9 15 13 2
24 3 2 16 4 9 13 2 3 2 12 5 2 3 4 14 1 11 13 1 9 0 12 9 2
29 7 15 13 3 2 13 9 9 2 13 3 9 11 2 11 1 9 2 12 1 10 9 2 9 2 9 2 2 2
18 1 0 9 13 9 9 9 2 3 15 13 9 1 11 1 0 11 2
22 9 7 1 9 13 0 9 13 9 1 0 0 9 0 1 10 9 16 3 0 9 2
15 3 0 9 1 0 9 13 9 9 2 3 9 7 9 2
20 1 9 15 13 9 9 1 9 12 2 12 9 1 9 2 15 3 13 12 2
32 0 0 9 0 9 2 15 4 13 10 0 3 0 9 2 13 3 1 15 3 3 2 3 1 12 5 1 15 15 13 9 2
7 10 9 13 1 9 9 2
28 9 3 13 1 9 1 9 2 3 0 9 13 3 9 13 2 16 4 13 3 0 9 2 15 13 9 9 2
30 9 3 13 1 12 9 2 16 15 9 9 13 13 0 9 9 0 9 9 2 7 16 1 15 13 9 0 2 2 2
14 0 2 0 9 13 3 1 9 1 9 1 0 9 2
31 9 15 13 0 0 9 7 13 15 2 16 1 15 9 15 13 12 9 1 9 2 12 13 0 9 9 2 0 9 9 2
10 7 10 9 15 13 3 10 9 9 2
5 3 9 13 1 9
19 9 15 13 9 1 9 12 9 9 2 9 0 2 2 15 13 1 9 2
11 1 9 1 9 13 9 7 13 2 2 2
30 1 9 2 3 9 13 9 0 9 1 12 9 2 13 1 9 9 7 15 10 9 15 3 13 15 9 3 1 9 2
15 13 1 9 2 14 1 9 15 13 2 16 4 15 13 2
13 13 13 15 0 2 16 15 9 13 1 12 9 2
12 2 15 13 7 9 9 9 0 9 2 2 2
23 3 13 7 15 9 13 7 13 15 1 9 2 7 16 0 0 2 9 2 13 3 0 2
15 3 9 13 10 9 9 2 15 3 13 3 0 7 0 2
15 9 13 2 16 13 7 0 9 1 0 9 9 2 9 2
22 15 13 1 9 0 1 9 2 7 1 12 9 7 15 2 13 2 7 13 1 9 2
13 7 9 15 3 13 3 9 16 9 10 0 9 2
5 3 15 11 13 9
24 0 9 13 9 9 1 9 7 9 1 9 2 12 1 12 5 2 1 0 9 12 9 9 2
15 9 13 9 0 9 7 9 9 2 1 12 5 3 2 2
21 9 9 13 1 12 5 3 2 9 9 13 1 9 11 7 0 9 11 12 2 2
20 3 13 7 0 9 2 9 1 12 5 2 2 7 9 2 7 12 5 2 2
27 1 0 9 9 1 9 13 3 11 1 12 5 0 9 1 0 9 2 7 3 1 11 2 11 7 11 2
3 9 0 9
17 0 9 13 9 2 12 0 0 9 0 9 1 9 0 0 9 2
13 13 1 3 0 9 2 10 0 0 9 3 13 2
42 16 15 3 1 11 9 2 12 13 2 0 9 15 1 15 13 3 3 7 3 15 13 2 16 11 13 3 3 1 15 2 1 0 9 13 1 15 9 0 0 9 2
41 9 2 15 13 13 0 9 9 9 7 0 9 9 1 0 9 2 7 13 0 9 7 15 0 2 9 2 9 2 0 9 2 9 2 13 1 12 5 2 11 2
20 3 13 3 2 16 4 9 10 9 13 9 0 0 9 2 7 15 13 3 2
16 3 11 13 2 16 4 9 4 13 3 7 3 3 0 9 2
22 2 13 3 0 9 0 15 2 16 9 0 1 0 9 13 0 9 13 2 2 2 2
16 3 3 3 10 9 2 1 9 0 7 1 11 3 3 0 2
6 1 15 11 3 13 2
7 3 13 10 9 7 9 2
21 13 15 2 16 1 10 10 0 9 13 3 13 2 7 13 9 10 9 7 9 2
32 1 0 9 9 11 4 13 13 0 9 10 9 2 13 9 1 0 9 9 13 10 0 0 9 2 9 7 9 1 0 9 2
17 16 4 15 13 13 3 0 9 7 1 9 7 9 2 13 0 2
17 9 13 1 0 9 0 1 9 1 9 13 13 3 3 0 9 2
7 0 2 9 2 1 0 9
29 3 16 9 0 0 9 13 3 7 0 11 2 13 15 1 0 9 7 9 10 9 11 2 11 2 11 7 11 2
17 1 0 9 13 0 13 2 16 10 9 13 1 10 9 3 0 2
18 1 9 0 9 3 13 1 9 0 11 13 1 12 0 9 7 9 2
26 3 13 1 10 9 1 12 3 0 9 14 1 9 12 9 2 12 5 1 15 1 9 0 11 2 2
18 13 15 0 9 1 0 0 9 7 9 1 11 2 11 7 0 11 2
31 3 2 1 9 0 9 13 1 9 1 0 9 7 0 9 0 9 9 2 1 9 7 9 1 0 0 9 7 0 9 2
34 9 11 0 1 11 2 9 9 11 2 13 3 12 9 1 0 9 11 2 11 7 11 7 13 0 12 9 1 9 1 9 0 9 2
5 9 7 9 0 9
16 1 10 9 15 15 13 2 16 0 9 0 9 13 0 9 2
10 3 0 0 0 9 13 7 3 0 2
12 3 3 13 0 9 10 9 1 9 2 12 2
34 0 9 11 11 2 11 2 11 13 2 16 9 13 1 15 12 0 9 2 0 9 2 9 1 0 9 2 0 9 7 1 0 9 2
4 9 7 9 2
18 13 0 9 2 16 4 15 9 1 0 9 3 13 12 2 12 7 2
30 13 1 0 0 9 0 2 16 4 3 2 1 3 0 0 9 13 9 3 12 5 7 0 9 15 13 1 0 9 2
19 0 0 9 13 3 13 9 9 12 2 0 9 7 9 9 9 2 9 2
17 1 9 0 9 15 4 13 0 0 9 11 14 1 9 2 12 2
17 13 15 1 15 2 16 1 15 4 3 13 12 9 1 0 9 2
13 9 2 12 4 13 4 13 0 9 2 11 12 2
11 9 0 9 1 11 13 11 9 2 12 2
20 1 9 2 12 15 13 1 9 12 11 1 11 7 3 7 9 0 0 9 2
9 3 16 11 3 13 1 10 9 2
7 13 15 0 9 1 11 2
28 11 15 3 13 1 9 1 0 9 0 11 2 1 0 9 11 2 16 0 11 13 0 9 1 0 9 9 2
18 7 16 9 2 16 11 15 13 3 1 0 9 0 9 2 13 0 2
5 13 11 0 9 2
18 1 11 15 13 12 2 0 0 9 0 9 9 3 0 0 0 9 2
11 9 11 13 3 1 0 9 0 0 9 2
22 1 0 7 3 0 9 1 9 12 9 13 7 1 9 1 9 1 10 9 7 9 2
8 10 9 13 13 1 9 9 2
19 9 13 7 12 9 2 3 0 2 9 2 15 4 1 10 9 3 13 2
35 0 0 9 15 3 13 7 15 7 1 10 9 2 16 1 9 13 1 10 9 9 2 3 9 13 1 9 9 1 9 12 2 12 9 2
21 13 15 2 16 1 0 12 9 12 5 15 9 0 1 0 9 13 9 12 9 2
44 9 11 7 3 13 0 2 3 3 0 9 1 0 9 9 2 12 1 15 2 16 4 9 1 0 9 13 1 0 9 11 2 9 4 13 1 9 7 12 9 13 10 9 2
42 0 9 0 9 11 2 11 2 11 13 2 16 15 13 1 10 9 1 10 9 2 1 9 2 3 2 2 14 1 9 2 16 4 7 11 13 0 0 9 16 11 2
26 0 4 7 1 10 9 13 3 0 9 2 0 15 2 1 15 13 0 9 2 11 2 11 7 11 2
23 12 0 9 4 13 13 11 7 13 9 11 2 15 4 16 0 9 13 0 0 9 11 2
11 15 13 0 13 1 9 12 2 12 9 2
29 11 2 11 13 2 16 16 13 0 9 2 12 9 9 2 1 9 9 2 12 2 2 13 0 9 1 12 9 2
12 13 1 0 9 0 9 10 9 13 7 0 2
18 3 16 15 10 9 13 13 0 7 0 9 2 15 13 1 9 11 2
12 9 2 15 13 11 2 13 1 9 1 9 2
29 13 2 16 15 1 15 3 13 11 7 11 2 15 1 9 1 11 7 11 13 1 0 9 16 11 1 9 11 2
8 9 13 3 13 9 10 9 2
34 13 15 7 11 3 13 14 1 9 2 7 7 1 11 2 3 15 13 9 11 2 7 1 11 2 1 15 9 15 7 9 11 13 2
18 13 15 2 16 0 9 0 1 9 1 9 2 13 0 9 1 9 2
22 0 9 2 15 4 13 0 13 12 9 2 4 13 7 13 0 14 1 12 9 3 2
8 7 15 3 13 9 0 11 2
7 15 15 4 13 2 2 2
11 0 9 13 1 10 9 3 0 0 9 2
14 13 15 3 3 1 9 2 15 13 0 9 7 11 2
11 13 1 9 1 0 9 7 1 9 9 2
9 1 0 9 9 13 1 12 9 2
13 3 4 0 9 13 1 9 12 1 9 0 9 2
14 1 10 9 13 13 12 9 2 11 11 7 11 11 2
20 11 3 13 1 9 0 9 7 1 10 9 13 2 7 13 2 9 0 9 2
8 3 13 9 9 9 9 9 2
17 12 0 11 13 1 9 3 7 13 13 16 12 1 0 0 9 2
13 1 9 4 15 12 13 13 1 0 9 1 11 2
20 1 0 9 1 9 12 2 12 13 0 9 1 0 9 11 9 1 9 11 2
16 3 15 1 15 13 0 9 2 1 10 9 15 13 1 9 2
20 13 0 2 16 1 0 9 13 7 0 0 9 0 9 1 0 9 1 11 2
7 9 1 9 9 13 0 2
14 9 2 12 13 1 10 9 0 9 1 12 0 9 2
17 13 13 2 16 15 13 3 2 7 16 1 9 11 7 3 13 2
15 9 1 9 0 0 9 7 11 7 4 1 0 9 13 2
18 10 0 9 15 13 2 16 15 13 3 7 13 1 0 9 0 9 2
25 11 1 10 9 13 1 9 1 11 3 9 16 0 9 1 0 9 2 16 9 11 13 3 13 2
15 13 15 9 2 16 7 11 1 11 13 3 3 2 2 2
10 6 10 9 7 9 0 9 2 2 2
2 11 11
7 2 9 2 9 9 9 9
47 1 0 3 0 9 1 0 9 0 9 13 2 16 9 10 9 9 3 0 0 9 13 15 3 0 2 7 15 1 0 0 2 16 13 3 2 9 9 0 2 14 1 0 9 1 9 2
22 3 1 10 0 9 15 13 1 0 9 9 0 0 0 9 2 15 13 0 0 9 2
32 10 3 0 9 13 3 2 0 9 7 0 2 2 0 2 0 2 9 2 9 2 15 1 10 2 0 2 9 13 9 2 2
20 13 15 1 14 3 0 9 1 15 0 9 2 10 9 4 13 3 0 9 2
17 0 13 15 3 9 1 9 9 2 0 1 10 0 9 2 9 2
26 11 2 11 2 1 9 11 12 2 12 2 12 2 13 1 0 9 2 15 4 1 10 9 13 13 2
19 0 9 0 9 13 1 9 1 9 2 9 2 0 9 1 9 0 9 2
28 10 3 0 0 0 9 7 14 10 0 0 9 15 13 1 9 1 0 9 2 7 2 1 0 12 9 9 2
19 0 9 15 13 1 9 3 10 0 9 2 1 9 10 0 2 0 9 2
21 0 9 9 2 3 2 0 2 9 0 9 2 15 13 1 0 9 0 9 9 2
22 1 9 13 3 0 9 9 3 0 9 1 9 3 0 9 1 9 9 2 10 9 2
8 0 9 4 13 9 0 9 2
12 0 9 13 15 7 13 9 0 0 9 9 2
2 11 11
13 1 9 2 0 9 11 11 1 9 12 7 12 2
12 1 9 11 11 9 2 9 2 7 0 9 2
25 0 0 9 2 9 2 9 9 2 2 15 1 0 9 11 11 1 11 1 11 1 9 9 13 3
2 9 13
38 0 9 11 2 11 2 11 11 2 11 12 2 12 2 12 2 12 2 13 1 11 9 9 2 9 0 2 7 0 0 9 2 9 2 9 0 2 2
25 13 9 9 12 2 9 9 1 9 9 12 9 2 7 13 15 1 9 1 9 12 9 1 9 2
10 1 12 9 15 1 9 9 9 13 2
24 13 15 2 16 9 7 0 0 9 13 12 5 9 7 0 1 15 13 1 10 9 1 9 2
9 9 9 13 0 9 1 9 9 2
6 15 15 13 7 3 2
24 1 0 9 4 13 9 7 9 9 13 13 1 9 2 9 13 2 16 4 15 13 9 9 2
18 0 9 13 1 3 0 9 3 15 2 1 10 0 9 15 13 9 2
12 0 9 13 15 7 12 5 1 15 13 9 2
17 9 13 9 14 1 9 9 2 7 10 9 13 1 10 9 0 2
24 10 0 9 9 13 2 7 9 1 15 13 2 11 12 2 12 2 12 2 12 2 12 2 2
18 9 9 2 9 14 3 13 3 0 9 2 0 9 13 9 13 9 2
13 1 0 0 9 15 2 0 9 2 13 3 3 2
27 1 9 15 13 1 15 2 16 9 13 0 0 9 2 9 13 9 2 7 13 3 0 9 1 0 9 2
17 9 4 3 13 2 16 3 0 9 2 1 9 2 13 0 9 2
29 9 13 7 3 3 2 0 9 15 3 13 9 9 7 10 9 1 9 9 13 13 9 2 15 13 3 0 9 2
18 13 0 13 3 3 2 7 1 15 9 13 9 7 9 13 1 9 2
15 3 0 13 9 1 0 9 0 0 9 2 13 9 0 2
9 9 7 9 9 11 11 2 9 2
11 3 2 0 9 0 11 1 9 12 2 9
18 3 2 9 11 1 9 9 0 0 9 13 1 9 1 9 2 12 2
8 1 9 0 9 2 9 11 11
42 3 2 0 9 1 9 2 9 11 2 11 2 13 0 12 9 7 13 3 2 1 0 11 2 0 9 0 9 0 11 2 2 9 2 0 1 9 9 0 1 15 2
19 1 9 11 11 2 9 7 9 0 9 2 9 2 12 2 11 2 11 12
13 3 2 0 9 11 1 0 11 13 9 7 9 2
18 1 9 0 0 0 9 2 11 11 2 11 11 11 12 2 9 2 12
13 9 0 11 1 9 0 9 2 9 12 2 9 2
8 1 9 0 9 2 9 11 11
51 9 13 11 11 2 9 12 2 12 2 12 2 12 2 12 2 7 13 2 14 10 0 9 2 13 2 2 2 2 2 13 1 15 2 15 15 3 3 0 9 13 1 9 0 9 0 0 9 2 2 2
19 1 9 13 13 15 2 7 15 7 0 0 9 0 9 9 2 2 2 2
29 0 9 3 13 9 9 2 10 9 13 3 14 0 2 4 3 3 1 0 9 13 9 1 9 2 9 1 9 2
13 9 12 13 0 3 3 16 9 15 1 10 9 2
27 1 9 13 1 9 2 7 1 9 9 2 15 4 13 9 9 2 14 3 0 0 9 9 2 2 2 2
4 9 11 2 11
3 11 11 2
4 0 7 0 2
26 9 9 13 7 3 0 9 9 7 13 3 10 0 9 16 9 9 7 7 13 13 9 15 1 9 2
41 9 4 3 13 15 2 16 0 9 13 1 9 1 9 2 3 9 1 9 13 13 2 16 0 2 3 0 9 15 3 13 1 15 2 16 4 3 1 9 13 2
26 9 11 7 11 0 2 0 11 2 9 12 2 9 2 12 2 1 9 11 11 1 9 2 12 7 12
24 3 0 0 9 9 15 3 1 0 9 11 13 1 9 2 16 13 3 9 16 3 0 9 2
30 16 9 13 9 0 9 1 9 9 2 13 9 0 9 2 7 0 9 1 9 0 9 13 10 9 1 9 0 9 2
15 9 11 7 11 0 2 0 11 2 9 12 2 9 2 12
38 3 2 9 9 9 9 2 15 13 1 11 9 0 0 9 2 1 9 0 0 9 2 11 11 2 11 2 11 2 11 0 11 2 0 2 0 11 12
38 3 2 9 1 0 9 9 9 9 0 2 11 2 1 2 11 2 1 9 9 2 15 13 0 1 0 9 7 13 3 13 1 0 11 3 0 9 2
17 15 9 13 1 0 9 2 9 2 1 9 9 2 9 1 11 2
21 12 0 9 13 0 9 9 12 2 12 2 12 0 13 0 9 9 12 2 12 2
3 9 11 11
34 9 11 11 2 0 9 2 1 0 9 9 11 1 0 0 11 1 11 2 3 16 0 0 9 13 1 9 12 7 12 9 0 0 9
24 0 9 0 9 0 9 9 0 2 11 2 0 1 9 11 11 1 0 9 1 0 11 1 11
12 9 0 9 9 0 2 11 2 1 10 9 2
9 9 9 1 9 2 12 13 11 11
20 9 9 9 1 9 11 11 1 9 9 9 1 9 7 9 12 2 9 11 11
20 11 11 2 11 2 12 2 12 2 0 9 9 2 9 12 9 2 9 11 11
32 11 11 2 9 2 12 2 9 2 9 2 12 5 12 5 12 9 2 9 1 9 9 1 9 1 0 9 9 2 9 11 11
7 9 9 1 9 9 1 11
50 0 9 11 11 2 11 2 11 2 11 2 13 9 0 2 9 1 0 7 0 9 2 2 1 15 15 13 2 16 9 0 9 1 9 9 9 1 9 9 15 1 9 2 12 13 1 12 9 9 2
28 9 13 0 9 10 9 1 12 9 9 1 9 3 0 9 2 7 0 0 9 1 9 0 9 7 0 9 2
46 3 15 13 2 16 9 1 9 9 0 9 13 3 12 2 12 9 1 9 2 1 9 1 12 2 12 9 1 9 1 9 9 9 7 12 7 3 9 1 9 1 9 9 1 9 2
15 3 0 9 13 0 1 10 9 0 2 0 7 0 9 2
9 1 11 13 0 9 12 0 9 2
10 3 12 5 10 9 15 13 1 9 2
25 1 15 13 3 12 9 2 15 4 13 1 9 0 12 9 7 3 15 3 1 9 0 9 13 2
23 0 9 9 15 13 1 9 3 0 2 3 1 0 9 2 9 0 9 7 0 9 9 2
34 16 12 1 9 9 0 9 1 9 0 9 15 1 9 13 9 9 0 1 9 9 1 9 0 9 11 11 1 0 9 1 9 12 2
31 3 13 1 3 12 9 9 13 0 9 1 9 12 9 2 0 0 11 12 2 12 2 9 2 12 2 9 2 12 2 2
2 11 11
3 12 2 12
5 9 9 13 0 9
44 9 0 9 2 3 9 1 9 9 0 1 9 0 9 7 9 9 2 3 13 1 0 9 7 13 13 0 9 0 9 0 9 1 0 9 2 11 12 2 12 2 12 2 2
45 11 11 2 11 1 0 9 7 10 9 13 2 16 0 9 0 9 13 0 0 9 9 0 0 9 1 12 7 12 9 1 0 9 2 15 13 0 1 0 9 9 0 0 9 2
18 0 9 13 9 12 9 2 0 9 0 0 9 7 9 0 9 9 2
20 1 9 1 10 0 9 13 0 9 1 9 0 9 7 13 13 3 10 9 2
9 1 10 9 15 13 10 9 3 2
32 3 15 13 2 16 9 0 9 13 1 0 0 9 14 0 9 2 0 2 7 0 2 11 12 2 12 2 12 2 12 2 2
2 11 11
6 1 0 9 2 2 2
59 9 2 12 9 0 9 1 9 1 12 0 9 9 13 0 9 1 0 9 2 0 0 0 9 2 2 13 0 0 9 7 3 13 3 12 9 2 1 9 9 2 16 13 9 0 9 2 13 9 12 2 12 2 12 2 14 12 9 2
39 0 13 15 2 16 15 13 9 2 15 3 13 9 2 16 4 9 9 10 9 13 2 7 3 13 0 2 13 0 0 9 2 1 10 9 13 9 9 2
10 13 10 9 2 15 9 3 2 13 2
11 9 1 9 13 13 0 2 16 13 9 2
7 9 3 3 4 13 9 2
39 0 9 9 15 13 1 9 0 9 7 13 2 3 9 13 4 13 1 9 2 3 15 9 13 13 1 0 9 9 9 2 3 15 9 13 13 9 3 2
16 9 2 12 9 13 12 9 9 7 13 3 13 12 9 9 2
26 9 13 9 0 9 2 7 3 13 0 9 1 0 9 1 9 2 13 15 7 9 2 3 1 15 2
16 10 15 4 13 1 2 0 0 9 2 2 0 11 1 11 2
26 7 3 3 2 1 12 2 9 2 12 2 1 9 12 13 13 2 0 9 11 1 0 9 9 2 2
20 2 3 13 0 9 2 9 2 7 3 13 9 9 0 2 9 2 7 0 2
8 2 3 13 9 2 3 0 2
11 16 13 0 9 1 9 0 2 13 0 2
6 2 0 9 13 3 2
24 2 16 0 9 13 2 13 2 16 13 4 13 1 9 1 12 2 9 7 1 12 2 9 2
3 13 9 2
11 2 16 13 3 0 9 2 3 15 13 2
24 2 3 13 9 0 9 1 0 2 3 2 13 13 0 9 1 9 2 3 4 13 0 2 2
30 2 13 15 9 3 2 3 1 9 1 0 9 7 0 9 2 1 9 1 9 2 9 2 7 3 9 2 2 2 2
22 2 13 0 9 0 2 3 15 3 13 2 16 9 13 13 3 0 7 13 2 2 2
12 2 13 0 9 1 9 2 9 7 0 9 2
8 2 13 14 0 7 0 9 2
2 11 11
15 9 2 1 15 13 0 9 2 7 9 13 13 2 9 2
15 3 13 1 0 11 9 2 2 2 2 2 1 0 9 2
24 16 15 9 1 0 9 13 1 9 2 13 2 9 2 9 9 2 15 15 1 9 13 13 2
16 0 9 13 0 9 2 10 9 1 0 9 4 13 13 9 2
26 3 15 7 13 2 16 10 9 2 9 9 2 13 0 9 9 9 1 9 15 2 16 13 9 9 2
14 3 13 9 0 9 2 3 0 2 1 9 0 9 2
22 1 10 9 1 3 0 9 13 7 13 12 5 9 2 11 12 2 12 2 12 2 2
27 1 0 9 1 9 13 16 15 1 9 13 1 9 9 1 9 7 14 7 0 9 9 0 9 0 9 2
20 1 9 4 3 13 0 7 0 9 2 1 15 7 1 1 9 13 0 9 2
18 3 7 1 15 13 9 2 7 16 0 9 13 2 0 9 0 9 2
1 11
2 0 9
11 9 13 0 9 0 0 9 1 10 9 2
13 13 15 9 0 9 2 3 0 0 7 0 9 2
6 10 9 9 13 9 2
14 13 9 0 9 7 9 7 10 9 13 3 0 0 2
39 13 0 3 16 9 7 3 1 9 15 13 0 0 9 2 3 0 9 2 1 0 2 2 0 0 9 2 2 0 9 9 2 1 15 13 0 0 13 2
15 13 0 9 0 2 0 0 9 2 7 13 15 9 2 2
11 1 15 13 0 9 1 9 3 16 9 2
12 3 1 9 2 7 1 9 13 9 13 3 2
12 13 15 2 16 9 13 9 9 0 0 9 2
39 0 9 13 9 1 3 0 9 9 0 15 0 9 2 0 9 13 0 9 0 9 2 0 9 7 0 9 7 13 9 2 1 15 13 2 13 2 9 2
18 9 0 9 13 0 9 0 15 1 9 9 7 9 2 1 0 9 2
43 1 0 9 4 1 0 9 0 9 13 9 0 9 2 15 13 3 0 3 1 9 9 0 9 2 9 2 7 1 0 2 0 2 9 2 11 12 2 12 2 12 2 2
20 13 15 2 16 13 1 9 2 10 9 13 0 1 0 9 0 9 0 9 2
21 3 0 0 9 0 9 1 9 0 9 13 0 2 16 7 13 0 1 0 9 2
15 9 15 3 13 1 0 9 9 7 9 0 9 0 9 2
25 0 9 9 0 9 0 9 3 13 1 0 0 9 10 14 3 0 2 0 7 10 9 0 9 2
2 11 11
3 0 0 9
19 9 0 9 1 0 9 0 0 9 15 3 13 0 7 3 0 9 9 2
51 1 9 1 0 9 15 13 3 12 0 0 9 7 15 13 13 14 1 0 9 2 7 3 1 0 9 9 2 9 7 9 2 1 9 9 13 9 2 16 0 9 13 0 2 13 1 2 9 9 2 2
25 0 3 0 9 0 9 1 0 9 13 2 0 9 2 2 9 0 9 2 0 1 9 2 12 2
21 0 9 1 0 9 11 4 13 11 2 11 2 1 9 0 7 1 9 0 9 2
16 4 13 11 7 11 14 1 9 2 12 2 3 4 13 11 2
30 1 2 0 9 2 13 9 0 2 0 9 2 7 15 13 9 1 11 0 2 0 9 0 2 7 11 2 9 11 2
15 10 9 15 3 13 9 12 2 9 7 9 15 13 3 2
15 13 0 9 2 7 13 3 7 11 7 10 9 13 0 2
16 11 13 10 9 13 1 9 9 9 2 16 4 13 10 9 2
9 7 13 13 1 9 2 13 9 2
19 9 15 11 2 13 10 9 2 13 1 9 1 9 0 1 9 0 9 2
14 9 13 3 13 7 13 7 15 13 1 9 11 0 2
9 13 13 1 9 1 9 9 11 2
5 15 1 15 13 2
14 13 15 9 1 9 9 10 9 2 16 3 13 3 2
15 7 3 2 9 9 13 13 3 0 2 16 9 0 9 2
19 15 13 2 16 9 15 13 3 13 2 13 7 3 2 16 15 13 9 2
1 11
5 1 9 0 7 0
22 3 15 3 13 9 1 15 2 3 13 0 2 0 9 7 3 13 9 1 9 9 2
25 0 4 13 12 9 2 7 16 15 3 10 9 1 9 3 13 2 13 2 16 13 0 0 9 2
8 1 9 9 15 13 10 9 2
24 10 0 7 0 13 7 9 9 2 15 16 9 13 2 13 2 7 1 15 3 3 13 4 2
45 13 3 10 9 2 7 15 13 0 9 2 16 10 9 13 14 3 3 13 1 0 9 2 13 0 9 7 0 0 9 2 7 3 13 1 9 2 13 2 7 13 1 0 9 2
48 13 15 3 7 0 2 9 0 9 13 3 13 3 2 13 15 3 1 9 7 13 15 1 10 9 7 9 13 7 0 2 2 16 4 3 13 9 2 16 9 13 9 7 4 13 10 9 2
19 14 7 0 0 9 13 0 9 9 0 9 2 1 15 13 14 12 9 2
8 9 15 7 13 13 3 0 2
40 13 15 9 0 0 9 2 1 15 15 13 9 9 9 9 1 9 9 2 7 1 9 9 2 2 3 0 1 9 9 2 7 9 13 0 7 0 9 9 2
36 7 9 15 3 13 13 1 9 9 7 1 10 9 9 2 16 4 3 3 13 1 15 2 16 0 13 7 13 0 13 0 9 1 0 9 2
52 3 15 3 3 13 9 2 11 11 2 9 2 2 9 9 2 12 2 12 2 9 2 12 2 2 1 15 15 13 13 2 16 4 7 13 1 15 2 16 7 1 10 9 13 10 9 2 15 10 9 13 2
7 13 15 7 3 3 0 2
38 13 1 9 1 15 2 16 7 9 2 0 0 9 2 13 13 0 2 16 15 2 15 3 3 3 13 16 9 9 9 0 9 2 3 13 1 9 2
26 3 3 1 3 0 9 9 15 13 13 10 3 0 2 9 0 9 2 3 3 2 16 1 9 0 2
54 13 7 0 9 2 16 7 1 10 0 9 4 3 13 9 2 10 9 9 3 14 13 2 7 15 2 1 15 9 7 3 3 13 10 0 9 2 7 1 15 3 13 3 0 9 7 2 13 2 0 9 10 9 2
40 7 15 7 3 2 16 0 13 2 16 7 16 15 9 7 9 3 13 1 0 9 2 15 3 13 0 9 1 9 9 7 15 3 10 9 9 1 0 9 2
43 1 15 4 7 13 13 2 15 13 10 0 9 2 0 3 3 1 10 9 2 3 1 9 13 2 7 3 7 3 13 1 9 3 0 9 2 3 13 9 1 9 9 2
43 7 15 3 3 13 2 16 3 9 13 3 9 2 1 15 13 10 9 2 1 1 9 10 0 9 2 14 3 0 2 13 3 2 9 12 2 12 2 12 2 12 2 2
20 3 2 7 3 3 2 3 13 13 1 15 9 1 9 2 0 9 2 11 2
53 9 2 15 13 0 9 9 1 0 9 7 13 10 9 3 0 0 9 2 3 13 10 9 1 9 1 0 9 10 9 2 16 10 9 2 15 13 1 0 9 1 10 0 9 2 13 1 9 2 0 0 9 2
52 7 9 2 15 1 10 9 13 1 0 9 2 14 2 0 0 9 7 9 2 13 3 0 9 13 3 0 9 2 16 9 2 15 15 10 9 13 1 9 13 14 1 15 2 7 3 3 7 1 0 9 2
28 16 13 1 9 0 9 2 13 1 15 3 13 15 10 0 9 2 15 3 3 13 2 3 13 1 0 9 2
44 13 10 9 2 1 10 9 2 15 13 9 2 2 15 13 15 3 7 15 3 2 16 13 10 9 1 10 9 1 0 15 9 2 0 3 0 9 12 9 2 1 0 9 2
66 7 15 1 9 0 9 3 0 2 0 15 9 9 1 0 9 7 0 9 2 7 0 2 0 1 9 0 9 2 0 9 13 7 3 15 13 1 0 9 2 1 0 9 1 15 2 1 9 2 0 2 9 9 1 9 2 14 1 9 9 9 2 3 7 13 2
37 9 2 15 15 1 10 9 13 1 9 2 15 3 3 13 1 0 0 9 3 1 10 9 2 3 0 9 0 9 7 9 13 15 1 0 9 2
48 15 2 15 15 15 13 2 7 1 0 9 13 2 3 13 15 2 3 2 13 10 0 9 7 13 15 0 9 0 0 9 2 15 13 9 2 7 3 9 1 0 9 9 2 0 2 9 2
31 16 7 2 3 13 9 2 11 2 13 15 2 15 3 0 9 13 2 16 4 15 1 10 9 13 7 13 15 10 9 2
32 0 9 2 9 0 9 1 9 9 13 1 10 9 13 3 1 9 2 3 0 2 2 16 1 9 2 1 15 1 9 13 2
18 13 13 2 16 9 15 9 13 7 13 15 1 0 9 3 0 13 2
16 16 13 1 0 9 7 9 9 2 13 15 3 1 15 13 2
52 7 3 13 10 0 9 2 3 9 1 9 1 0 9 2 16 4 15 13 13 0 9 7 16 4 1 15 0 9 9 13 13 0 2 7 16 3 0 2 9 1 0 9 2 7 10 0 9 1 10 9 2
22 16 15 1 15 10 13 2 13 1 15 1 10 9 3 13 0 9 1 9 9 9 2
8 9 15 13 9 9 1 9 2
62 15 13 13 9 2 16 3 3 3 2 7 0 9 9 7 9 9 0 9 2 9 2 7 3 9 2 7 3 9 0 9 2 9 7 0 9 2 3 9 9 1 9 9 7 9 2 16 1 9 9 10 9 2 1 9 1 9 2 9 3 13 2
13 7 3 1 9 3 13 3 9 9 9 10 9 2
28 14 4 15 3 13 13 1 0 9 2 16 15 13 3 0 7 14 3 13 1 9 0 9 13 9 15 0 2
28 1 0 1 15 4 13 13 9 2 7 3 9 1 9 2 7 15 1 3 0 9 7 3 2 7 3 9 2
27 15 4 13 4 13 0 9 9 2 7 15 7 3 2 1 0 9 2 3 15 0 9 1 15 3 13 2
37 7 13 4 3 0 13 1 3 0 16 0 9 9 2 0 9 9 2 2 3 0 2 2 2 9 2 0 9 2 2 15 3 13 10 0 9 2
28 15 1 9 1 9 2 11 2 1 10 0 2 2 3 0 0 9 1 0 9 2 9 9 2 2 3 13 2
32 13 7 1 10 9 2 16 0 9 9 1 0 9 13 0 9 7 16 4 15 10 9 13 13 2 9 0 2 3 0 2 2
28 13 4 7 13 9 3 1 10 9 2 15 13 10 0 9 2 1 0 9 2 0 1 0 0 9 10 9 2
7 9 2 11 11 2 9 2
20 2 9 2 9 7 9 7 0 1 0 9 2 2 9 12 2 12 2 12 2
35 9 2 11 2 11 13 9 7 9 1 9 9 2 1 15 13 1 9 13 2 7 3 9 2 1 15 13 2 7 15 15 13 1 9 2
41 2 13 1 15 2 16 4 9 2 7 2 9 0 1 2 9 1 0 9 2 2 4 13 15 2 3 3 9 13 1 0 9 2 3 2 0 1 0 9 2 2
24 13 10 9 13 3 3 0 2 7 13 15 9 0 9 1 0 1 9 9 2 0 9 2 2
29 13 0 9 3 0 9 2 15 13 0 9 7 1 0 9 0 9 2 3 3 2 16 4 10 0 9 13 0 2
20 13 3 0 9 2 15 1 9 13 3 13 2 14 1 9 9 0 9 2 2
25 0 2 3 0 9 0 11 2 15 1 0 0 9 13 3 2 16 13 0 0 9 1 0 9 2
46 1 0 9 2 16 0 9 13 10 0 9 1 2 9 0 9 2 2 3 2 16 13 14 3 0 2 13 9 10 9 0 1 9 1 10 9 2 7 3 15 13 9 10 0 9 2
15 13 2 0 9 2 9 7 0 9 9 13 3 9 0 2
28 13 14 2 16 0 9 13 1 9 9 0 9 7 9 9 1 9 9 9 1 0 0 9 13 1 9 0 2
22 2 13 1 15 2 16 12 9 13 3 13 3 2 3 2 3 16 12 2 0 9 2
47 7 16 15 4 13 14 9 7 9 2 7 9 10 9 2 16 13 3 7 13 9 9 1 9 2 4 13 0 0 9 7 0 2 16 0 2 9 1 9 2 7 9 13 14 12 9 2
10 9 10 9 13 1 15 13 10 9 2
11 13 7 2 16 3 10 9 13 12 9 2
22 1 10 9 13 7 1 15 2 16 0 9 13 13 16 9 0 0 9 1 0 9 2
17 9 9 2 3 1 0 9 2 7 0 2 13 0 9 9 9 2
24 13 4 9 2 16 4 1 9 9 13 13 10 9 1 9 7 13 13 15 13 1 0 9 2
16 13 4 3 13 1 0 7 0 9 2 15 10 9 3 13 2
7 9 2 11 11 2 9 2
21 1 9 9 2 11 2 11 1 9 2 11 11 2 9 12 2 12 2 12 2 2
34 2 2 2 9 2 11 1 9 2 12 2 12 13 9 7 9 1 0 0 9 1 0 9 1 11 12 7 1 0 9 3 3 13 2
27 13 7 0 9 2 1 0 9 4 9 2 12 1 0 9 13 0 0 0 9 2 0 9 3 1 11 2
23 13 4 15 15 13 2 16 3 2 13 4 3 14 0 9 9 9 7 9 9 13 9 2
22 16 0 1 9 9 2 12 15 9 2 11 13 11 11 2 9 1 0 0 9 2 2
5 9 2 11 2 11
11 3 7 3 13 0 9 2 1 9 10 9
11 2 2 2 3 3 13 1 9 0 9 2
21 1 0 9 2 16 13 0 9 7 9 2 15 13 2 16 3 13 1 0 9 2
16 1 0 9 15 3 3 13 16 1 9 1 9 1 10 9 2
12 10 9 16 9 0 9 15 13 3 1 9 2
33 1 0 9 15 7 0 9 13 1 10 9 2 1 15 0 0 9 13 15 13 2 16 9 9 1 0 9 13 13 15 1 15 2
33 9 0 9 13 4 7 13 3 2 16 4 13 0 9 3 15 2 15 3 1 0 9 1 9 13 2 0 9 2 9 2 9 2
39 13 3 13 0 0 9 1 9 9 2 1 0 9 7 1 10 9 1 9 2 16 4 13 2 2 15 15 0 9 13 2 1 10 9 13 9 0 2 2
50 13 2 14 0 9 1 9 9 9 1 9 10 9 2 1 9 0 9 7 0 9 9 2 4 13 3 2 2 11 11 13 7 13 7 13 15 9 2 7 10 9 9 7 9 13 1 9 1 12 2
7 7 3 9 13 13 2 2
19 0 9 15 13 3 0 3 2 3 15 1 15 13 9 9 0 0 9 2
24 15 15 13 15 1 0 9 1 9 2 15 13 9 1 0 9 2 15 13 0 7 0 9 2
34 15 3 15 13 1 0 9 9 2 15 3 13 1 9 9 2 16 2 9 15 13 1 9 13 2 16 4 9 9 13 0 9 2 2
26 0 9 4 14 13 9 15 2 15 3 13 0 9 1 9 0 9 2 7 16 15 13 13 0 9 2
36 0 9 15 13 13 14 1 0 9 2 7 7 1 9 9 2 7 9 7 9 2 13 3 1 10 9 2 15 1 10 9 13 1 0 9 2
11 10 9 7 13 0 9 0 1 9 9 2
11 1 15 13 0 13 3 9 7 0 9 2
20 3 0 0 9 4 3 3 13 7 10 9 2 15 13 1 9 3 0 9 2
5 0 9 13 9 2
23 3 1 0 9 15 13 1 9 10 9 13 0 0 9 2 16 13 9 2 9 7 9 2
24 0 9 15 13 13 3 10 9 1 9 2 16 4 13 2 3 13 0 13 9 0 9 3 2
19 10 9 3 13 4 13 14 1 9 2 7 3 1 0 9 2 2 2 2
9 9 2 9 2 11 11 2 9 2
12 0 9 2 9 12 2 12 2 12 2 12 2
3 2 2 2
15 11 2 11 13 0 9 1 9 7 9 9 10 9 9 2
33 9 2 1 15 13 15 0 2 13 3 3 0 2 7 9 13 0 9 9 0 9 2 16 15 0 13 13 2 3 3 2 0 2
19 3 0 0 9 13 9 2 15 15 13 0 0 9 10 9 7 0 9 2
34 3 4 13 9 1 9 9 7 9 2 9 13 9 2 0 9 0 9 2 15 0 3 13 7 13 13 1 0 9 14 1 0 9 2
21 9 9 13 0 9 2 7 3 15 3 1 10 9 3 13 2 9 13 3 0 2
32 0 9 16 9 9 2 9 0 0 9 2 2 9 2 7 7 9 9 2 9 7 3 0 9 13 3 14 0 7 0 9 2
37 0 7 0 9 13 1 10 9 9 3 0 9 9 3 1 0 9 2 3 9 9 13 1 0 9 0 9 2 7 7 1 9 0 9 10 9 2
13 2 0 0 11 1 11 12 2 12 2 12 2 2
2 11 11
14 1 9 1 9 2 9 12 2 12 2 12 2 12 2
7 13 4 13 3 12 9 2
12 2 1 9 13 14 9 2 15 0 13 9 2
14 14 1 9 7 1 9 2 7 1 15 4 13 9 2
13 0 1 9 2 1 9 2 1 0 13 9 2 2
4 2 11 11 2
6 9 2 11 11 2 11
23 1 0 9 13 3 0 0 9 13 3 1 9 12 0 9 1 9 2 9 15 13 0 2
7 11 11 2 3 0 9 2
9 0 9 2 11 12 2 9 2 12
3 0 9 11
21 3 1 12 2 7 12 2 9 12 13 11 11 9 10 9 11 2 11 2 11 2
7 12 9 15 1 9 13 2
19 13 15 2 15 13 3 3 15 0 9 1 9 7 3 13 1 10 9 2
35 12 7 0 13 1 9 10 9 3 0 9 2 16 13 1 9 10 9 9 0 9 2 15 1 10 9 13 0 9 7 13 15 7 11 2
12 10 9 13 2 7 3 1 10 0 9 13 2
28 9 0 9 13 1 15 2 16 0 7 0 3 9 13 2 16 13 9 10 9 2 3 2 14 13 15 13 2
33 7 9 13 13 0 2 13 2 14 15 13 3 0 9 9 7 13 2 14 15 16 9 13 0 0 9 7 15 0 13 0 9 2
27 13 15 15 2 16 0 9 1 9 13 3 9 7 9 9 10 9 2 7 3 0 9 2 1 15 13 2
58 9 0 9 2 7 3 3 9 2 2 15 15 13 9 16 14 1 9 2 3 3 1 9 1 9 1 15 2 15 13 9 0 9 0 9 9 7 1 9 0 9 2 13 15 1 15 2 16 1 9 13 9 2 13 9 7 9 2
66 3 4 7 13 13 1 9 0 9 1 0 9 7 0 0 9 2 15 13 3 3 2 16 13 1 9 9 0 2 3 0 1 9 0 9 2 7 13 15 0 9 2 16 4 13 2 3 15 13 9 10 7 15 9 2 10 9 2 0 9 7 9 9 1 9 2
28 7 13 2 14 15 9 10 9 1 0 2 7 9 1 15 10 9 13 2 2 13 15 0 9 0 16 9 2
22 10 9 13 3 13 15 15 2 15 13 0 9 2 7 13 15 10 9 13 0 9 2
27 13 9 9 9 2 1 15 10 9 15 13 2 1 15 13 13 0 9 2 16 7 9 13 13 15 0 2
12 3 15 0 9 13 7 1 0 9 2 2 2
29 0 9 2 15 15 9 13 9 9 2 13 1 15 2 16 9 13 0 9 2 13 2 1 15 13 0 9 9 2
14 7 2 13 15 0 9 2 15 13 3 0 9 0 2
34 13 1 15 2 16 1 9 1 9 9 7 0 9 13 3 1 9 9 2 3 3 16 9 2 13 15 15 0 13 13 1 9 9 2
56 7 9 13 1 15 2 16 1 9 13 9 3 10 9 2 15 13 3 13 1 9 2 7 7 15 9 3 13 10 9 2 16 9 13 9 2 15 13 13 3 9 9 9 2 7 7 9 0 2 7 7 15 13 3 13 2
8 1 10 9 15 13 15 13 2
17 14 9 0 9 13 7 13 2 3 15 13 15 7 0 0 9 2
11 9 9 13 13 9 1 9 0 9 9 2
22 15 13 7 1 9 13 1 0 9 9 2 9 9 7 9 13 9 9 0 10 9 2
14 0 9 13 1 10 9 9 9 7 1 15 13 0 2
26 1 0 9 13 3 13 1 0 9 2 7 10 9 13 1 0 9 14 3 7 3 15 13 0 9 2
4 13 11 2 11
15 2 2 11 13 0 9 2 1 15 15 11 13 10 9 2
15 1 9 1 10 9 4 13 14 3 1 11 9 2 12 2
28 3 0 9 4 13 3 3 1 9 2 11 2 11 2 9 7 9 2 2 13 9 2 9 9 2 12 2 2
8 2 13 7 9 13 11 9 2
4 1 9 1 9
6 9 12 2 12 2 12
50 1 9 9 2 12 0 9 1 9 2 12 13 11 2 11 2 11 9 11 2 11 2 11 7 11 2 11 9 1 9 2 9 2 15 13 0 9 1 9 16 0 11 9 2 3 9 1 9 2 2
24 9 3 13 9 0 9 7 9 2 7 15 15 13 10 9 2 15 15 13 9 7 9 9 2
47 7 3 9 2 16 0 9 4 13 1 9 2 3 1 0 9 2 13 3 0 2 3 15 9 13 9 2 9 2 9 2 15 13 0 13 1 0 9 2 7 16 15 13 10 9 13 2
14 16 10 9 13 0 2 13 9 9 2 3 10 9 2
45 3 3 0 13 7 1 9 9 9 2 3 9 3 0 7 0 14 1 11 7 9 0 0 9 2 3 13 9 0 0 9 2 16 4 15 15 13 13 3 1 11 7 1 11 2
43 13 14 13 2 3 13 10 9 9 9 1 0 9 9 0 11 2 7 3 9 2 16 9 0 0 9 0 9 2 0 9 9 11 11 2 15 13 1 9 3 13 3 2
66 9 10 9 2 0 1 0 9 1 15 9 2 13 14 11 2 9 2 0 9 7 9 9 0 9 2 13 1 9 1 15 1 0 9 2 15 15 13 0 9 2 16 15 3 13 1 0 7 0 9 2 13 15 3 1 10 9 2 7 3 1 15 13 13 0 2
30 1 0 9 3 1 10 9 13 0 9 11 11 7 9 15 13 9 3 13 10 9 1 0 9 2 15 13 3 13 2
6 7 13 1 0 9 2
73 13 2 14 11 1 9 2 16 11 9 13 11 2 7 16 15 11 15 15 0 13 2 7 16 0 1 9 13 10 0 9 2 16 15 13 9 2 10 9 13 3 13 3 2 16 16 10 9 13 9 0 9 1 0 9 2 2 3 10 12 9 13 2 16 7 1 0 9 13 9 9 0 2
23 1 9 13 1 0 9 2 0 13 3 2 1 9 2 7 3 15 13 3 1 0 9 2
26 11 2 11 2 11 15 13 3 2 7 13 15 1 11 2 1 11 3 2 1 0 9 0 9 11 2
6 0 9 13 16 9 2
19 1 9 15 13 2 1 9 13 7 3 3 1 9 15 13 1 9 0 2
68 3 13 0 1 11 2 11 2 11 2 11 2 1 0 9 1 15 13 11 11 2 1 0 9 1 15 13 11 11 2 13 15 1 11 2 11 2 1 9 0 2 1 11 2 11 2 11 2 11 11 2 1 9 2 1 11 1 11 2 7 3 1 15 4 13 11 11 2
56 1 10 9 13 0 13 2 16 9 2 12 13 11 2 11 2 11 2 2 0 9 9 0 13 4 9 10 2 1 0 9 13 15 4 9 1 9 10 7 13 9 9 10 2 4 3 13 1 0 9 0 2 2 2 2 2
40 9 1 0 9 2 15 13 11 1 9 2 13 13 7 0 7 0 2 0 0 9 13 0 7 1 9 9 0 2 16 13 1 0 9 3 9 9 11 11 2
41 1 15 13 3 0 0 9 11 0 9 2 7 0 9 3 13 2 16 1 0 9 13 1 9 13 13 2 1 9 7 9 0 9 2 7 3 13 10 9 3 2
2 11 11
3 11 11 2
4 9 1 11 2
8 9 0 9 1 3 0 11 2
9 0 9 2 9 11 2 11 2 12
16 9 2 11 11 13 9 9 7 9 1 0 9 11 1 11 2
23 1 9 2 12 13 1 9 9 9 1 0 9 11 7 1 0 9 13 0 9 0 9 2
16 9 13 0 1 0 9 0 9 1 9 0 9 7 9 11 2
24 0 9 13 10 0 0 0 9 2 9 0 9 2 2 15 9 2 12 13 3 1 9 11 2
18 13 15 2 16 0 9 3 1 10 9 13 2 15 13 15 9 9 2
19 9 3 4 0 9 7 7 3 13 3 3 1 0 9 7 1 0 9 2
32 13 9 2 16 15 3 0 9 13 2 15 3 15 1 9 13 2 7 16 13 0 13 0 9 2 16 0 9 13 15 0 2
16 0 9 0 9 7 1 0 0 9 0 9 13 13 0 9 2
19 13 15 13 0 0 9 2 9 0 9 2 9 0 9 0 1 0 9 2
37 7 13 15 3 13 9 0 9 2 10 0 7 0 9 7 3 1 0 9 3 0 9 16 13 9 7 9 9 1 9 1 9 0 7 0 9 2
15 1 9 9 0 0 9 15 11 2 11 13 9 1 11 2
25 1 0 9 9 11 2 15 13 3 1 0 9 12 2 9 2 13 1 9 7 9 9 3 15 2
10 13 12 1 10 0 9 3 0 9 2
8 13 1 9 0 11 1 11 2
15 3 13 10 9 2 3 13 1 0 9 7 1 0 9 2
24 3 2 3 7 3 3 13 11 2 11 9 2 1 15 13 2 10 0 9 2 9 0 9 2
16 13 2 10 9 13 1 9 2 15 13 7 13 0 0 9 2
21 9 0 9 7 1 0 13 1 9 0 9 1 9 2 1 9 7 1 0 9 2
14 1 9 0 9 13 13 9 9 1 9 7 0 9 2
15 0 9 1 10 3 0 7 0 9 13 3 0 16 0 2
33 1 9 15 3 13 0 9 7 3 1 0 9 10 0 2 9 2 15 9 3 13 2 1 10 9 7 1 10 9 13 9 13 2
35 1 9 2 12 13 0 9 3 1 9 9 2 7 3 1 9 9 2 0 2 13 0 2 9 2 7 1 9 0 7 0 9 9 9 2
13 3 3 15 1 15 13 9 2 9 7 9 9 2
27 1 10 9 13 11 2 11 1 9 9 0 9 9 9 2 11 11 2 7 13 3 3 0 7 0 9 2
20 13 14 9 2 16 1 10 0 9 1 9 13 1 9 9 3 3 0 9 2
2 11 11
20 2 1 9 9 13 13 1 10 0 9 7 9 2 7 3 15 13 0 9 2
18 10 9 13 3 3 9 7 0 9 2 7 16 4 13 0 0 9 2
24 15 3 13 1 0 9 2 16 13 1 15 9 2 15 13 13 10 9 1 9 1 0 9 2
31 16 7 15 13 12 9 7 13 0 2 16 13 3 1 9 1 0 9 2 3 3 13 9 0 7 13 15 1 9 2 2
5 11 2 1 9 11
7 9 9 1 0 9 9 2
43 1 9 15 13 1 12 9 7 9 1 9 0 9 1 9 11 11 1 11 2 16 4 13 9 0 9 1 9 9 2 1 0 9 1 9 7 9 1 9 2 0 9 2
28 9 0 9 15 13 7 1 9 10 9 2 3 9 12 9 11 11 2 1 0 0 2 9 2 9 2 2 2
38 9 2 11 11 1 10 9 15 13 1 0 9 10 9 2 3 13 2 16 10 9 1 9 15 1 9 13 9 2 0 2 9 10 0 9 2 2 2
13 9 13 1 9 9 7 0 0 9 1 0 9 2
42 13 15 1 9 9 9 0 9 2 1 9 1 0 9 2 1 15 2 16 15 9 1 9 13 0 9 0 1 9 2 1 9 0 9 1 9 1 0 9 2 2 2
4 1 9 1 9
72 9 9 2 13 11 2 11 2 9 12 2 12 2 12 2 12 2 12 2 1 0 0 9 2 15 13 9 9 7 1 15 13 9 9 15 0 9 2 13 1 0 9 1 9 3 0 9 1 0 9 9 2 16 4 15 1 15 2 1 9 2 9 7 10 9 1 0 9 3 13 13 2
49 7 16 4 15 9 13 0 2 13 11 2 11 9 2 0 2 11 2 12 2 9 12 2 9 12 2 12 2 1 9 2 16 9 2 15 13 9 9 2 13 14 3 0 2 16 13 0 9 2
19 0 0 0 9 2 15 4 13 1 9 9 2 13 1 0 9 3 0 2
27 15 4 13 2 16 9 1 9 0 9 13 3 0 2 16 3 13 9 9 2 7 3 9 9 3 0 2
6 11 12 2 12 2 12
5 9 9 1 9 2
16 1 0 0 9 3 9 0 13 15 9 1 9 9 1 9 2
24 3 4 13 12 9 9 1 3 10 9 2 1 15 12 7 1 9 7 14 1 3 1 9 2
21 3 13 15 3 2 15 3 3 3 13 13 2 16 13 9 9 1 9 3 0 2
7 9 9 13 15 1 9 2
8 15 9 14 1 0 13 0 2
11 1 12 13 9 3 1 9 2 2 2 2
9 9 12 2 9 12 2 9 2 12
3 9 7 9
2 11 11
16 1 10 0 9 9 2 12 13 9 1 11 0 9 0 9 2
18 0 9 10 9 3 13 0 9 9 2 1 15 9 0 11 3 13 2
32 1 9 15 3 13 0 9 7 0 9 2 0 9 7 9 1 9 9 7 9 0 2 9 7 0 9 1 9 7 0 9 2
33 1 9 0 0 0 9 13 10 9 3 0 2 0 9 13 0 9 1 9 2 0 2 1 2 0 2 2 16 15 13 9 0 2
27 15 13 9 7 15 9 2 15 9 7 15 9 15 13 14 3 7 14 1 0 9 2 3 13 1 9 2
20 9 0 9 13 7 14 3 3 9 13 1 9 15 14 1 9 9 0 9 2
30 3 3 12 1 0 13 3 13 1 9 9 7 9 9 2 0 11 3 3 13 9 9 7 9 7 13 15 1 15 2
37 16 13 0 9 1 9 7 9 13 3 0 9 13 3 1 9 0 2 15 2 15 15 13 2 14 16 9 11 1 9 2 9 9 7 9 9 2
11 0 9 9 13 3 10 0 9 0 9 2
27 15 15 1 0 9 1 0 9 13 7 0 0 9 3 16 9 0 9 13 9 0 2 0 7 3 0 2
22 1 0 0 9 13 15 7 3 2 3 0 9 13 13 1 9 2 0 9 7 3 2
25 3 0 9 9 13 3 9 7 9 7 9 2 0 9 15 2 16 12 9 1 0 9 13 3 2
18 0 13 13 15 1 0 9 1 9 0 9 2 3 1 10 0 9 2
24 0 9 7 9 2 3 7 9 9 2 15 1 12 2 2 12 2 9 13 0 9 7 9 2
30 16 13 13 1 9 10 9 2 0 9 3 1 9 13 7 3 12 9 2 2 13 13 7 0 9 1 0 9 0 2
24 7 0 9 4 3 13 3 1 9 9 2 13 1 0 9 1 0 9 7 0 9 0 9 2
14 3 9 12 2 9 13 0 9 0 0 9 0 9 2
50 1 9 0 9 15 13 0 9 0 0 9 2 15 13 0 9 11 1 10 9 2 13 15 1 0 9 9 2 0 9 7 9 2 9 3 2 16 7 1 0 9 2 3 1 9 13 9 9 2 2
43 0 9 10 1 0 9 3 0 9 13 12 0 9 2 1 9 13 9 0 9 2 16 3 0 9 9 2 7 0 9 1 9 0 9 2 9 0 1 9 7 0 9 2
21 3 0 9 0 9 13 9 9 3 0 2 0 7 0 1 9 3 16 1 9 2
19 1 9 9 0 11 15 13 9 2 16 13 3 15 13 1 0 9 15 2
25 13 3 3 0 9 2 9 0 9 0 9 13 3 0 7 0 2 0 7 0 2 3 3 0 2
18 3 0 9 0 9 9 0 11 13 3 11 2 11 1 10 9 9 2
6 15 16 10 9 13 2
17 13 3 0 13 9 2 16 0 9 9 1 10 9 9 13 0 2
28 7 1 9 10 0 9 4 0 2 0 0 9 13 13 1 9 10 0 9 2 0 2 16 15 13 3 9 2
7 9 7 2 0 2 0 9
2 11 11
32 9 1 0 9 0 16 2 0 2 9 4 13 0 9 2 9 0 9 2 0 7 0 9 2 3 2 0 9 0 9 2 2
27 0 9 1 9 7 3 13 1 0 9 1 9 7 1 0 9 0 2 0 2 7 3 14 3 0 9 2
39 10 2 0 2 9 0 9 13 9 0 2 2 0 9 2 2 9 12 2 12 2 12 2 2 3 2 7 9 0 2 2 0 9 2 2 0 0 9 2
14 2 9 2 13 0 0 9 2 0 1 9 7 9 2
9 1 11 15 3 13 1 0 9 2
30 0 0 9 13 9 1 0 9 7 1 9 2 9 0 2 15 13 9 0 9 2 9 2 9 2 9 7 9 9 2
11 3 13 0 3 0 9 0 9 10 9 2
29 9 1 9 9 7 9 0 9 0 9 1 9 0 13 3 0 9 7 9 2 11 2 11 2 11 2 11 2 2
33 0 9 1 9 11 2 12 2 12 2 12 2 13 1 9 1 9 2 9 2 2 15 15 13 9 2 12 2 11 2 11 2 2
21 13 7 0 9 1 0 9 9 2 12 2 11 2 7 9 2 12 2 11 2 2
18 0 9 0 1 9 9 0 13 9 9 9 2 7 2 3 0 9 2
4 12 2 12 2
21 9 13 1 9 3 3 2 13 0 9 2 13 9 0 9 7 9 9 1 9 2
18 13 1 9 12 0 0 9 2 1 0 2 9 2 7 1 0 9 2
26 13 1 9 16 9 2 13 3 10 9 2 5 9 2 3 9 2 13 9 12 2 12 2 12 2 2
26 0 9 1 9 2 0 3 13 9 9 2 13 3 7 1 9 10 9 3 1 9 9 1 9 9 2
26 0 9 0 9 4 13 1 9 15 9 9 0 14 3 1 9 2 9 2 9 2 9 2 9 2 2
45 1 15 15 13 12 2 2 16 1 0 0 9 13 9 9 2 3 2 9 1 9 2 9 2 2 1 0 9 0 2 7 2 16 4 13 9 2 16 4 4 3 13 0 9 2
12 1 9 9 9 9 1 9 13 3 0 9 2
22 1 9 9 1 9 2 0 1 9 15 13 3 9 1 0 9 2 1 9 7 9 2
47 12 9 0 9 13 1 9 2 9 2 16 1 9 2 3 4 13 0 9 9 1 9 2 0 1 0 9 9 0 2 15 10 9 2 13 15 9 2 13 9 9 1 0 0 9 9 2
13 3 0 13 9 1 9 9 2 9 2 1 9 2
16 7 13 0 3 13 1 9 0 1 0 9 7 9 3 0 2
26 3 2 11 7 0 2 12 2 13 2 16 0 9 0 9 1 0 9 13 1 12 9 9 1 9 2
34 3 4 13 0 9 0 9 2 9 1 9 7 0 0 9 2 7 9 0 9 9 2 9 9 7 9 2 9 15 13 0 0 9 2
12 13 0 9 9 7 9 4 13 9 9 9 2
14 10 9 13 3 0 2 0 9 1 9 2 2 2 2
14 9 13 9 7 1 9 2 7 3 9 9 4 13 2
17 1 15 0 9 1 9 7 9 13 0 13 2 16 9 13 3 2
49 13 2 14 15 11 2 0 0 11 2 11 2 13 11 2 12 2 9 1 9 9 2 1 9 9 2 7 16 3 1 9 0 9 2 13 13 3 1 9 3 0 0 9 2 0 1 9 9 2
23 13 9 1 0 9 9 2 3 2 9 1 9 9 2 9 2 2 7 9 13 3 0 2
22 1 9 0 9 2 15 13 3 0 9 2 13 14 9 2 9 2 0 9 10 9 2
24 0 9 2 0 1 9 0 2 9 0 2 13 9 1 0 9 1 9 1 2 0 2 9 2
13 13 16 0 9 3 7 3 2 7 13 3 0 2
45 3 0 0 9 2 15 10 9 7 9 3 13 0 0 9 2 13 0 0 9 7 13 15 7 1 9 9 2 15 13 9 2 15 13 0 9 9 2 7 13 3 1 9 0 2
34 1 10 9 9 0 1 9 2 12 2 12 2 12 2 13 13 1 9 1 2 0 2 9 3 0 2 3 4 15 1 0 9 13 2
30 0 9 12 9 0 5 13 1 9 2 0 2 9 14 9 2 7 7 10 0 9 2 11 12 2 12 2 12 2 2
39 0 9 1 0 9 9 1 11 9 2 12 13 3 0 7 3 4 3 13 3 10 0 9 2 3 9 2 15 15 10 9 3 3 13 1 0 0 9 2
29 10 9 2 7 2 9 9 9 1 9 0 0 9 2 9 2 9 2 13 13 1 0 9 3 1 9 0 9 2
13 11 13 1 9 9 3 9 3 0 0 9 11 2
34 0 9 9 1 9 9 2 9 2 13 0 9 9 2 15 1 9 0 9 2 3 13 9 1 9 0 0 0 9 2 13 13 0 2
24 1 9 1 9 2 12 13 1 11 1 12 9 9 2 9 2 1 0 9 12 9 9 3 2
19 9 0 9 15 1 10 9 13 14 14 12 2 7 15 3 1 0 9 2
16 3 13 9 2 0 2 7 0 9 2 13 0 9 7 9 2
24 1 9 0 9 7 1 0 9 9 15 13 1 9 1 12 9 0 9 1 12 9 0 9 2
38 1 9 0 9 2 15 13 3 0 3 1 0 9 2 13 0 9 12 7 0 7 1 9 12 9 15 13 9 9 1 12 9 9 9 2 9 2 2
24 9 1 9 11 13 3 3 7 13 9 1 0 9 2 9 2 1 9 1 0 9 0 9 2
25 13 0 13 2 3 15 9 1 0 9 2 11 2 13 1 0 9 9 1 9 9 1 9 9 2
1 9
2 9 11
7 0 9 7 0 9 9 9
2 11 9
20 1 9 15 9 13 13 7 13 9 9 9 9 0 1 15 0 7 0 9 2
18 13 2 14 0 9 0 2 13 3 3 1 9 3 0 9 0 9 2
23 0 9 1 9 9 2 1 9 10 0 9 1 10 0 9 2 13 9 2 3 2 9 2
25 9 0 9 2 10 9 7 9 15 13 9 2 3 10 9 13 7 3 15 10 9 1 9 13 2
35 3 9 9 0 9 13 1 9 2 3 7 3 10 9 13 7 3 15 13 1 0 9 2 3 3 3 1 9 9 2 15 13 10 9 2
14 9 9 9 2 15 13 9 0 9 2 15 13 0 2
20 15 13 9 9 1 10 0 9 2 0 9 2 1 14 12 2 12 9 9 2
9 1 11 3 13 0 9 10 9 2
27 1 9 9 0 2 9 0 2 13 1 3 16 12 9 9 1 0 9 0 9 1 11 1 0 0 9 2
22 0 9 1 0 9 13 1 9 10 0 9 2 15 13 3 7 13 1 15 0 9 2
22 3 7 13 0 9 9 0 1 15 2 16 4 15 9 13 1 9 16 12 0 9 2
34 1 9 0 9 9 2 9 0 2 13 1 0 9 3 7 3 1 0 9 9 2 16 15 1 10 9 13 3 3 0 0 0 9 2
15 0 9 3 3 13 10 0 9 7 16 12 9 13 3 2
37 1 10 9 15 7 1 9 13 0 9 2 3 9 9 9 9 2 9 2 2 9 2 1 15 13 13 15 9 0 1 9 7 9 9 16 9 2
22 1 9 9 13 0 9 2 9 2 2 15 2 16 9 13 2 13 13 7 13 15 2
14 10 9 13 1 9 3 0 7 3 0 1 0 9 2
29 1 9 9 9 13 13 0 9 2 13 11 2 9 12 2 12 2 12 2 2 15 13 0 9 1 0 9 9 2
31 9 9 1 11 2 11 2 11 13 9 0 1 0 9 9 2 15 13 0 15 2 16 4 1 9 13 3 1 0 9 2
30 9 2 9 7 9 2 13 1 10 9 3 9 1 9 2 1 9 2 2 16 9 1 9 2 1 9 2 15 13 2
16 9 3 10 9 7 1 15 0 9 2 9 2 13 0 9 2
29 9 13 9 3 12 9 0 9 7 9 0 9 7 1 0 9 11 2 0 9 0 9 2 1 15 13 0 9 2
27 9 13 13 1 9 0 9 2 7 2 13 15 13 0 9 1 0 9 1 3 0 9 9 2 9 2 2
4 9 2 12 2
31 13 12 0 9 2 0 9 1 9 13 1 9 0 9 2 13 2 2 16 10 9 13 0 2 7 13 3 13 3 9 2
18 3 12 1 12 0 9 0 9 13 3 1 11 2 9 2 12 2 2
23 15 13 2 16 0 0 9 2 3 2 9 2 10 9 13 0 0 9 2 13 1 11 2
12 3 0 9 7 13 9 2 3 0 9 13 2
36 3 4 15 13 2 16 9 9 9 13 3 0 7 16 15 13 13 0 9 2 1 0 9 15 13 12 2 12 5 0 9 1 12 9 9 2
20 3 4 7 0 9 9 2 3 0 0 11 2 13 1 0 12 2 12 9 2
10 0 9 1 9 13 3 0 12 5 2
55 4 15 13 3 2 16 1 0 9 13 1 11 3 0 9 9 0 2 15 13 3 13 0 9 9 9 3 1 11 2 7 3 7 1 0 9 0 9 2 3 13 9 0 0 9 9 0 1 11 3 10 9 12 9 2
20 1 10 9 13 3 0 2 16 1 9 13 15 0 9 9 7 3 13 9 2
10 1 10 0 0 9 3 13 12 9 2
32 13 15 2 16 1 12 9 13 1 11 14 12 9 0 9 2 7 3 1 12 1 10 9 13 15 0 9 2 1 9 2 2
29 4 13 3 10 3 2 0 9 10 9 7 15 15 13 3 1 0 9 2 3 7 1 9 9 2 3 9 13 2
8 1 10 9 15 13 3 9 2
26 9 3 13 2 16 13 10 9 2 15 4 13 9 0 9 1 11 7 9 0 9 1 14 12 9 2
29 3 1 9 0 9 2 0 0 0 9 1 0 9 2 3 2 11 2 2 13 0 9 0 9 9 1 0 9 2
20 3 9 2 16 4 3 0 13 10 9 3 1 9 2 13 1 9 3 0 2
17 1 15 1 10 9 13 3 7 3 15 9 3 3 13 7 13 2
21 13 3 7 0 9 2 16 0 9 4 1 11 0 9 3 13 7 13 9 0 2
44 3 13 10 0 9 7 1 3 0 9 1 0 9 7 9 7 13 9 2 16 13 3 1 9 10 12 0 9 2 1 15 3 13 1 0 9 1 0 9 10 0 9 9 2
50 9 9 9 7 13 2 16 1 9 9 9 4 3 1 0 9 2 3 4 0 9 1 11 13 2 3 3 2 3 2 1 0 11 2 2 13 13 1 0 9 10 9 9 3 0 16 0 12 9 2
9 0 9 0 9 7 15 15 13 2
11 0 9 9 15 13 0 0 9 0 9 2
31 1 0 9 9 13 1 9 9 13 15 0 0 9 7 13 15 1 0 9 9 2 15 7 13 7 10 9 0 9 2 2
21 9 15 1 0 9 13 3 0 9 2 3 2 0 9 7 15 13 1 9 0 2
15 13 0 2 16 10 9 13 1 3 0 9 0 9 9 2
27 7 13 0 2 16 10 9 13 1 0 9 0 9 9 0 2 14 3 15 2 15 13 1 0 9 9 2
10 3 3 3 13 0 0 9 0 9 2
33 1 9 0 9 7 13 1 0 9 0 9 9 1 15 2 13 1 9 0 16 1 0 9 7 3 0 16 1 0 7 0 9 2
10 0 9 15 13 9 2 0 2 9 2
49 13 0 2 16 16 4 9 9 9 13 1 14 12 2 12 7 0 0 9 1 0 12 2 12 5 9 1 9 9 2 13 4 15 9 9 9 1 12 14 1 12 9 9 7 13 4 1 9 2
29 13 4 9 0 9 1 11 7 9 4 3 13 9 9 0 2 15 1 10 9 3 13 11 7 13 9 0 9 2
34 9 7 1 9 13 0 9 9 9 2 9 7 0 9 2 15 3 3 13 9 16 0 0 9 10 9 9 2 1 15 15 13 9 2
12 3 3 3 13 0 9 9 10 9 1 9 2
32 13 3 1 0 9 9 9 0 2 1 15 3 13 15 10 0 9 2 7 13 1 9 0 1 0 9 9 0 9 0 9 2
7 3 13 9 3 0 9 2
23 13 0 15 3 2 13 2 16 9 10 9 1 0 9 15 13 7 13 1 10 0 9 2
25 9 0 9 10 9 7 9 10 9 3 13 1 9 0 7 3 13 9 0 9 2 9 10 9 2
32 13 0 15 13 2 16 1 0 9 9 2 12 9 4 13 13 3 2 12 9 2 4 13 10 0 9 3 13 1 0 9 2
17 3 0 9 9 9 4 13 9 0 9 0 9 10 3 0 9 2
19 13 4 15 3 9 0 9 2 16 0 9 9 4 13 9 15 0 9 2
25 16 1 11 15 1 9 13 0 9 2 1 0 11 4 13 7 1 9 0 9 0 9 1 11 2
23 3 4 15 13 9 0 0 9 1 0 9 7 10 9 1 9 0 2 3 13 0 9 2
17 10 9 4 13 9 1 9 9 7 10 9 3 13 1 9 9 2
15 3 10 9 7 13 9 2 16 9 13 1 3 0 9 2
17 10 2 9 9 2 0 1 9 12 0 9 13 3 13 1 9 2
23 13 15 3 2 12 2 9 12 9 2 1 15 0 13 12 9 2 9 13 1 9 2 2
21 10 12 9 9 13 1 0 9 2 10 9 13 3 2 13 9 9 7 9 9 2
16 9 13 1 9 0 9 7 12 2 0 2 13 9 0 9 2
12 0 1 15 13 3 12 9 7 9 15 13 2
17 1 0 9 9 3 13 2 1 10 9 1 12 2 9 3 13 2
10 13 0 2 16 13 3 15 3 0 2
19 1 0 9 9 2 9 3 13 9 0 1 0 1 12 9 12 2 9 2
16 13 10 2 9 9 2 9 2 3 1 9 0 9 9 13 2
4 9 2 9 2
13 0 9 1 9 9 0 1 9 13 13 0 9 2
16 3 0 13 9 0 9 0 9 2 15 13 9 0 0 9 2
26 0 9 0 0 9 15 13 1 0 9 2 15 13 3 0 2 16 13 0 15 13 7 1 9 9 2
14 9 10 9 1 9 3 13 0 9 1 9 0 9 2
12 9 0 9 0 0 9 15 13 9 2 9 2
11 9 9 15 13 0 9 0 1 9 9 2
18 9 0 9 13 1 9 12 2 12 9 2 13 3 1 9 3 0 2
13 0 9 9 0 3 0 9 13 12 2 12 9 2
20 1 9 9 9 15 9 0 9 13 3 1 9 1 9 2 1 15 4 13 2
25 9 13 9 0 3 0 9 3 1 0 9 2 3 7 1 10 9 2 15 3 13 9 0 9 2
39 1 0 9 7 1 0 9 9 13 0 9 0 9 2 7 2 9 0 9 1 9 0 2 0 1 10 9 1 0 9 2 1 9 7 1 0 9 9 2
16 1 9 10 9 15 13 1 9 9 9 0 9 1 9 9 2
6 0 9 9 2 2 2
40 3 10 9 13 1 0 9 2 9 15 0 15 13 1 9 0 9 2 15 13 0 9 9 9 1 0 0 9 2 0 9 15 9 2 15 13 9 13 2 2
14 1 10 9 15 13 2 16 4 13 0 0 0 9 2
26 1 0 0 9 13 0 0 9 0 9 9 2 0 9 9 1 9 1 9 2 16 10 9 13 0 2
12 16 13 1 9 3 0 9 2 13 9 0 2
11 0 9 0 0 9 13 9 0 0 9 2
20 9 0 9 15 7 13 1 9 9 3 0 2 7 1 3 0 0 0 9 2
90 15 13 3 12 9 2 13 3 1 0 9 2 0 9 0 9 13 3 0 0 9 9 2 7 10 0 9 13 1 0 9 1 0 9 2 0 2 9 2 2 15 13 3 9 0 9 7 15 13 13 3 0 2 3 0 2 9 2 1 0 0 9 15 9 13 1 0 9 2 15 3 13 13 3 3 0 9 2 7 13 14 3 0 9 15 0 9 9 2 2
30 1 9 10 9 13 7 0 0 9 3 13 2 10 9 7 13 1 9 16 1 0 9 2 7 1 0 9 10 9 2
19 3 13 0 9 0 9 13 3 2 3 15 7 13 10 0 9 0 9 2
3 9 7 9
2 11 11
2 11 11
2 11 11
39 2 2 2 7 16 16 13 9 1 15 2 15 13 2 15 0 9 13 2 2 2 2 13 15 9 0 9 9 1 0 9 7 1 0 9 2 2 2 2
7 11 11 11 2 1 11 9
13 2 9 12 2 2 9 12 2 2 13 2 11 11
5 3 13 10 9 2
7 10 9 13 9 1 9 2
19 3 13 0 9 2 3 0 11 13 9 7 9 9 2 15 1 9 13 2
26 3 7 1 9 9 0 9 2 7 3 1 9 0 9 4 13 0 9 9 1 0 7 0 9 9 2
15 13 2 16 9 13 9 0 9 7 9 9 7 9 9 2
13 13 2 1 15 15 13 2 13 10 0 0 9 2
21 13 2 16 0 9 9 9 9 13 0 9 2 9 2 15 9 13 14 12 12 2
19 13 2 16 9 13 10 0 9 2 13 10 9 2 9 7 9 1 15 2
8 13 2 3 9 1 15 13 2
26 13 2 16 9 0 9 4 3 7 3 13 1 0 9 0 9 7 15 3 1 9 0 1 0 9 2
25 13 4 0 1 9 9 2 13 3 2 2 16 9 0 7 0 13 13 1 0 0 2 0 9 2
20 13 2 16 9 13 10 0 9 1 9 9 2 7 0 7 3 3 0 9 2
17 7 13 3 7 15 0 2 0 9 1 9 4 3 13 0 9 2
16 13 4 0 13 9 7 13 2 16 3 13 1 9 3 15 2
18 1 9 7 0 9 13 9 2 1 9 15 3 3 13 2 16 13 2
25 1 15 15 13 3 3 13 2 13 2 14 15 10 0 9 2 15 0 9 9 9 13 3 13 2
8 3 2 2 15 13 9 9 2
39 15 15 13 2 16 3 3 1 9 13 2 16 10 9 2 3 2 9 2 13 2 7 3 2 7 3 13 13 9 2 16 15 10 2 0 2 9 13 2
5 15 13 9 9 2
5 15 13 9 9 2
16 3 10 0 9 13 13 12 9 3 2 16 0 9 13 12 2
6 3 13 1 0 9 2
15 3 9 3 9 13 9 0 9 7 9 16 0 0 9 2
8 1 10 10 9 3 13 13 2
14 10 9 1 9 15 3 2 7 3 7 3 2 13 2
26 0 9 4 9 13 16 1 9 0 9 2 3 0 9 13 0 9 9 9 2 15 2 7 15 2 2
23 3 3 4 13 9 0 9 2 15 1 9 13 2 7 9 0 9 1 0 9 0 9 2
21 9 15 1 9 9 9 1 3 0 9 7 9 1 0 9 13 0 9 10 9 2
26 0 9 4 15 3 13 2 16 9 9 1 9 13 0 9 2 13 4 0 9 1 10 7 15 9 2
13 3 13 0 2 16 3 0 0 9 13 0 9 2
30 0 9 3 13 2 16 9 13 0 9 2 7 2 3 16 9 10 0 9 2 15 0 0 0 9 13 12 1 0 2
28 3 1 0 9 15 13 2 16 9 9 13 3 0 9 2 7 2 16 1 9 9 13 0 9 10 9 3 2
34 9 9 13 3 10 9 2 9 2 0 9 2 2 1 9 2 1 15 10 9 13 11 2 11 2 11 2 15 13 1 9 9 9 2
32 10 9 1 0 9 9 9 13 2 7 3 7 1 0 9 13 9 2 16 9 7 9 0 0 9 9 13 2 3 9 13 2
20 0 7 0 9 0 9 4 15 3 13 3 13 7 1 9 9 0 0 9 2
33 9 0 1 0 9 7 13 15 0 2 14 16 1 10 9 13 13 2 7 0 9 3 0 0 9 15 1 9 1 15 7 13 2
26 1 2 9 0 9 2 3 0 11 13 15 9 0 1 0 9 2 3 3 13 1 9 9 0 9 2
12 1 15 4 13 13 10 9 10 9 1 9 2
23 3 3 15 13 2 16 9 0 7 0 9 9 13 3 0 9 2 9 0 9 9 9 2
15 10 9 13 1 9 9 9 3 3 0 2 13 7 0 2
18 13 3 7 0 9 9 2 15 0 9 0 0 9 13 3 0 9 2
43 10 9 4 15 1 0 9 3 13 2 7 4 1 9 13 3 1 15 2 16 4 15 10 9 13 13 2 2 10 9 4 3 13 7 1 9 15 1 15 13 3 15 2
22 13 15 3 2 16 13 15 3 10 9 2 15 13 1 9 9 0 1 9 3 0 2
14 9 0 9 0 9 3 3 13 10 9 1 0 9 2
34 1 9 9 7 9 2 3 2 9 2 13 2 16 9 1 9 13 9 2 15 4 1 0 9 13 0 2 13 1 15 0 9 9 2
25 9 13 9 10 9 7 13 7 0 9 13 2 16 0 9 0 9 13 3 0 16 0 0 9 2
27 9 10 9 4 3 0 9 13 1 2 0 2 2 15 4 13 1 0 9 1 10 9 1 9 0 9 2
19 1 0 9 13 2 16 1 9 0 9 0 9 13 13 7 0 9 9 2
32 0 9 1 2 9 2 15 13 3 1 9 2 15 15 3 13 9 0 9 7 15 13 10 9 1 9 10 0 9 2 2 2
30 9 2 15 4 3 13 1 9 2 15 15 3 2 3 1 9 1 9 11 2 11 2 11 2 13 0 9 10 9 2
25 0 9 2 15 15 13 1 9 9 0 9 2 4 1 0 9 13 0 9 2 15 13 1 9 2
8 3 15 3 13 1 9 0 2
20 3 16 15 13 10 9 2 15 7 13 1 15 2 3 13 9 0 9 13 2
19 3 15 3 13 0 9 2 1 15 9 7 9 9 9 9 0 9 13 2
4 0 1 0 9
24 9 0 9 9 15 13 1 12 2 9 10 9 2 3 11 11 16 0 13 0 9 10 9 2
15 13 3 0 9 13 3 13 10 0 0 9 2 0 9 2
15 15 13 3 13 1 9 9 0 0 9 9 0 0 9 2
27 10 9 13 3 9 2 7 2 9 2 15 15 1 9 13 7 10 9 13 0 1 9 0 9 16 9 2
15 1 0 9 13 0 1 0 9 1 9 9 10 9 13 2
25 0 0 9 9 15 10 9 13 3 0 9 9 2 10 9 1 15 0 9 7 9 0 9 13 2
13 9 0 0 9 13 3 1 0 9 3 0 9 2
47 3 1 9 0 9 4 1 9 13 0 9 2 15 13 1 9 2 16 0 9 0 1 9 13 0 9 2 9 3 2 0 9 1 0 9 7 9 4 1 10 0 9 13 3 0 9 2
30 13 3 1 9 0 13 0 9 9 9 2 13 0 3 0 9 13 0 9 2 16 1 0 9 7 0 0 9 13 2
22 0 0 9 13 1 10 9 0 9 0 9 0 2 3 0 0 9 0 1 0 9 2
9 9 10 9 13 7 3 0 9 2
25 7 0 9 9 9 1 0 9 4 3 1 9 0 13 3 0 9 2 4 0 9 9 13 3 2
19 10 9 13 13 1 9 0 9 0 9 2 15 4 1 0 9 3 13 2
32 15 13 1 0 9 9 0 1 9 10 0 9 2 1 9 9 0 13 2 1 10 9 13 1 9 13 0 9 1 0 9 2
28 1 0 9 0 9 15 3 3 13 9 9 1 9 0 0 9 1 9 7 0 9 13 3 9 0 9 9 2
37 7 3 2 16 9 9 0 9 13 10 9 0 3 1 9 2 1 0 9 13 13 3 2 9 0 9 2 2 10 0 9 15 1 10 9 13 2
16 10 9 13 3 2 3 13 0 9 9 9 7 13 10 9 2
9 10 9 13 2 16 13 0 9 2
16 1 3 0 0 9 13 13 15 1 0 9 1 9 0 9 2
8 3 7 13 9 9 0 9 2
11 9 15 13 3 1 9 0 9 0 9 2
24 1 1 3 0 9 0 9 13 7 0 13 0 9 0 9 2 15 13 3 2 1 0 9 2
20 0 0 9 13 7 14 9 0 9 2 10 9 15 13 3 1 9 0 9 2
23 1 10 9 9 13 3 0 9 2 7 9 3 0 2 13 15 0 9 0 0 9 2 2
23 10 0 2 9 2 15 13 3 0 9 1 9 0 9 7 0 9 0 9 1 0 9 2
14 13 15 2 3 3 10 9 13 1 9 11 11 9 2
10 13 2 16 12 12 9 15 3 13 2
12 1 0 0 9 13 0 13 9 0 0 9 2
11 9 15 3 13 9 0 1 12 0 9 2
24 7 16 3 0 0 9 13 3 1 9 0 2 13 1 0 13 0 3 1 9 9 0 9 2
4 9 9 0 9
25 1 9 9 9 15 13 0 2 9 9 2 15 0 0 9 0 9 13 3 12 7 3 15 9 2
30 0 9 1 9 9 13 10 9 9 2 15 13 3 13 1 0 9 2 16 4 13 0 9 2 15 4 0 9 13 2
11 10 9 9 13 0 1 0 9 0 9 2
14 4 3 13 3 2 16 4 13 0 9 0 9 9 2
23 12 1 3 0 9 9 13 1 10 0 9 2 7 3 1 0 9 2 9 0 0 9 2
36 15 13 9 9 1 0 9 2 7 2 9 2 3 15 3 15 13 2 2 15 13 13 1 3 0 2 7 3 1 10 9 1 2 0 2 2
23 1 0 9 1 0 9 2 3 9 3 0 2 16 13 9 0 2 13 0 9 9 12 2
24 3 1 0 9 2 3 1 3 0 7 1 10 9 2 0 2 9 2 13 0 9 1 9 2
40 13 2 14 2 16 1 10 9 13 9 0 9 0 7 3 0 16 9 2 13 15 10 9 1 10 9 1 9 2 3 12 9 13 0 9 7 0 0 9 2
33 0 9 13 1 0 9 13 0 9 2 13 2 14 10 9 1 0 0 0 9 2 13 0 9 9 2 15 13 0 9 3 13 2
16 1 10 9 3 13 9 0 9 1 9 9 0 9 0 9 2
17 13 2 14 3 9 0 2 0 2 2 13 10 0 9 3 0 2
41 0 9 7 14 13 2 13 2 14 2 16 0 9 10 9 13 0 2 13 15 3 1 15 2 16 10 9 0 13 13 2 7 13 13 1 0 9 7 0 2 2
24 13 7 0 9 9 2 3 2 0 9 2 2 15 13 13 1 0 7 0 9 1 12 9 2
3 0 9 9
44 0 0 9 9 9 15 13 7 1 0 0 2 7 0 9 0 9 9 2 1 9 0 1 0 9 11 13 0 2 0 9 0 9 3 12 5 7 0 9 3 12 5 2 2
24 3 16 0 9 0 9 13 3 9 9 2 7 2 9 0 9 1 9 1 3 0 0 9 2
6 9 13 13 14 3 2
14 9 0 9 9 1 0 9 13 1 9 12 2 12 2
15 1 9 1 0 9 13 3 0 16 1 9 1 9 0 2
17 1 0 9 2 15 13 9 2 9 0 9 13 1 12 2 12 2
15 1 11 9 13 10 9 3 0 9 1 9 1 0 9 2
14 1 0 9 9 9 0 9 3 13 1 12 2 12 2
19 13 2 16 9 0 9 0 9 13 9 9 2 15 13 0 9 3 13 2
18 0 9 0 9 9 3 13 2 16 0 9 0 9 4 13 13 0 2
15 14 2 3 4 3 13 2 10 9 13 13 1 0 9 2
27 13 3 13 3 9 10 0 9 9 2 3 2 0 9 2 2 16 4 13 9 0 9 13 1 3 0 2
9 9 9 13 13 16 9 1 9 2
8 10 13 9 9 1 9 9 2
31 13 15 2 16 9 0 1 0 9 15 13 7 1 0 9 2 7 16 3 9 0 1 9 4 13 3 13 16 9 0 2
25 13 2 16 15 13 7 15 2 16 0 0 7 0 9 9 13 1 0 9 0 9 3 0 9 2
11 3 15 3 4 13 2 3 13 15 3 2
8 10 9 13 9 1 9 9 2
8 10 9 3 13 13 3 0 2
15 3 3 14 15 13 0 9 1 9 15 9 7 9 9 2
21 3 7 13 9 7 0 9 0 9 3 0 9 2 16 0 9 13 13 10 9 2
28 0 9 3 13 2 13 15 7 13 3 1 9 0 2 7 1 10 9 2 16 15 3 13 1 0 9 9 2
14 12 1 0 9 9 13 3 13 9 15 0 15 9 2
23 0 9 10 9 13 3 13 9 0 9 10 9 2 16 4 9 13 0 2 0 2 9 2
27 9 13 13 3 3 0 2 16 4 13 9 9 3 3 2 13 3 1 9 13 1 3 0 9 0 9 2
27 1 0 9 7 13 13 3 3 0 2 7 0 9 0 9 13 13 9 1 0 0 9 9 0 1 9 2
30 3 10 9 13 0 9 10 0 9 1 0 9 7 10 9 13 15 1 0 9 0 0 9 2 9 2 1 0 9 2
20 0 9 0 9 13 13 3 0 1 9 0 9 1 0 9 15 9 0 9 2
28 15 13 2 16 9 0 9 4 13 13 9 2 15 9 13 0 13 1 10 9 1 0 9 7 9 9 9 2
47 10 9 13 13 10 9 10 9 7 9 2 3 9 2 11 2 11 2 9 2 2 9 2 11 2 11 7 9 2 11 2 11 1 0 9 11 2 1 10 9 4 10 9 3 13 13 2
70 13 4 3 9 2 9 2 11 2 11 2 9 2 2 1 10 0 9 2 9 2 9 2 11 2 11 2 9 2 2 7 9 2 11 2 11 2 9 2 2 1 0 9 11 1 9 9 0 9 7 9 2 11 2 11 2 9 2 2 7 9 2 11 2 11 1 0 9 9 2
3 12 2 12
4 9 1 9 2
25 9 2 12 2 2 9 9 0 9 1 9 9 1 0 9 1 9 1 0 9 7 1 0 9 2
20 13 2 16 16 0 9 0 9 13 3 0 2 10 9 1 9 9 13 0 2
20 9 2 12 2 2 9 9 9 0 9 1 9 9 1 0 9 7 1 9 2
34 1 12 9 4 9 13 1 9 9 1 0 9 2 13 15 0 0 9 1 0 9 1 0 7 0 9 2 0 9 13 0 9 2 2
5 9 0 9 7 9
3 0 9 11
11 13 16 9 1 9 2 12 7 9 2 12
3 9 0 9
26 3 13 1 0 7 0 9 2 1 9 9 0 9 13 0 14 0 9 9 2 7 7 10 0 9 2
16 3 0 9 9 9 13 0 2 9 9 2 0 2 9 2 2
21 10 9 13 13 1 0 9 0 1 9 1 3 9 0 9 0 9 1 9 9 2
40 1 9 0 9 0 9 1 0 9 2 16 10 9 13 3 13 3 1 9 2 3 13 13 9 2 15 1 9 0 9 13 9 10 9 0 15 9 1 9 2
16 0 9 15 3 13 0 9 7 9 9 9 15 0 9 13 2
10 13 9 9 9 0 9 1 9 9 2
28 9 10 9 2 15 13 12 1 9 0 9 11 1 9 9 9 7 9 0 9 2 13 9 2 12 7 12 2
24 12 9 3 13 9 2 15 13 1 9 9 0 1 0 9 9 1 0 0 9 7 1 9 2
20 0 9 13 2 16 9 1 9 9 9 9 1 9 9 0 9 13 13 0 2
7 3 7 10 9 13 13 2
37 9 0 9 3 13 3 9 16 9 3 0 2 7 2 1 9 3 0 0 9 9 3 1 9 3 1 0 9 2 15 0 9 0 9 3 13 2
2 9 9
4 9 2 11 9
20 9 2 11 11 2 9 2 2 2 12 2 13 0 2 0 9 11 1 11 2
17 1 9 9 9 7 9 1 11 15 13 9 9 7 9 0 9 2
19 9 2 11 11 2 9 2 2 2 12 2 13 9 1 11 11 1 11 2
14 1 0 9 1 11 15 13 9 0 9 1 9 9 2
9 3 13 1 9 9 9 9 12 2
16 9 2 11 11 2 2 12 2 13 9 1 11 11 1 11 2
14 1 0 9 1 11 15 13 9 0 9 1 9 9 2
14 1 0 9 13 1 9 11 2 11 1 9 1 11 2
14 9 2 11 11 2 2 12 2 13 11 11 1 11 2
14 1 0 9 1 11 15 13 9 0 9 1 9 9 2
13 1 0 9 13 1 0 9 1 0 9 1 11 2
19 9 2 11 11 2 9 2 2 2 12 2 2 13 9 12 2 12 2 12
27 9 2 9 2 11 11 2 9 2 2 2 12 2 13 1 11 9 1 11 7 1 0 9 11 1 11 2
19 1 9 0 9 9 9 0 9 7 9 1 11 15 13 0 7 0 9 2
16 9 2 11 11 2 2 12 2 13 9 1 11 11 1 11 2
15 1 0 9 0 9 1 11 15 13 9 2 3 0 9 2
4 11 11 2 11
4 11 11 2 11
7 15 1 9 2 9 7 9
21 15 2 15 15 13 13 2 15 13 10 12 9 0 2 13 16 15 0 9 13 2
23 1 10 0 9 1 9 11 1 10 9 9 13 10 9 3 2 3 0 13 13 9 9 2
20 3 0 13 9 9 1 9 3 0 2 0 2 7 9 10 9 1 0 9 2
24 3 15 3 13 2 16 9 1 0 9 13 0 9 2 16 13 0 9 2 9 2 3 2 2
22 7 1 9 13 9 3 0 2 10 3 0 9 0 13 9 9 0 2 0 2 0 2
48 13 3 9 9 2 1 0 9 15 13 3 15 2 15 9 9 2 1 10 0 9 2 2 7 2 10 9 10 9 2 9 7 9 2 15 13 3 3 0 1 9 2 9 2 9 7 9 2
33 2 13 0 2 16 9 9 2 1 9 1 0 0 9 2 13 3 0 1 0 7 0 9 1 9 2 9 2 9 2 9 2 2
21 16 9 15 13 13 10 9 3 3 0 2 3 16 9 0 7 14 3 3 0 2
23 7 16 13 3 1 9 15 2 15 13 9 0 2 13 9 9 1 9 0 9 3 0 2
26 13 15 3 1 9 0 9 11 2 1 9 11 2 10 9 2 9 2 9 2 1 9 9 9 3 2
46 0 9 10 0 0 9 13 1 0 7 0 9 2 3 9 13 9 2 7 2 0 9 1 9 2 3 0 9 2 2 1 9 16 9 9 2 9 2 9 9 2 9 0 9 0 2
42 7 1 0 9 15 13 9 9 1 0 9 3 3 2 3 15 13 1 0 9 16 13 15 1 10 9 2 7 15 3 13 2 13 15 1 9 9 2 13 9 9 2
14 13 3 3 7 10 9 11 2 1 15 15 13 11 2
37 10 9 13 3 13 3 2 3 1 9 2 3 2 2 1 10 0 9 2 15 13 3 9 2 16 9 2 3 9 11 2 13 1 15 0 9 2
28 7 3 3 13 9 9 0 9 9 2 0 9 2 13 3 1 0 9 9 10 9 2 0 1 9 9 3 2
33 7 15 3 3 13 2 1 0 9 9 2 16 13 1 9 11 2 16 4 3 13 10 0 9 9 9 1 0 7 0 9 9 2
24 15 2 16 9 13 1 15 2 16 15 10 9 13 1 0 9 2 4 15 13 3 16 9 2
28 10 0 9 7 9 15 13 1 0 0 9 2 13 2 14 0 1 15 1 9 2 13 0 9 1 9 2 2
35 7 14 15 13 9 2 9 13 3 2 9 0 12 9 2 1 15 0 13 0 2 2 7 7 10 9 1 10 9 1 15 3 13 2 2
86 13 15 3 2 16 0 9 10 9 15 13 3 0 2 3 7 0 2 7 10 9 2 16 3 1 9 13 9 10 0 9 9 9 2 7 10 9 2 0 9 9 1 9 0 3 2 2 0 1 9 15 0 2 0 2 3 2 0 7 1 0 0 9 2 15 13 3 3 3 13 2 3 3 16 1 9 9 10 0 9 1 15 0 2 0 2
13 7 1 9 0 9 2 13 9 9 2 7 14 2
14 13 2 14 15 0 9 2 13 15 2 16 3 13 2
16 14 1 9 15 9 13 9 3 9 9 2 7 15 3 0 2
31 14 2 7 13 2 1 13 10 9 9 1 9 3 13 2 16 13 3 10 9 2 7 13 15 0 9 1 9 2 9 2
24 3 15 3 2 3 4 15 9 13 12 0 9 2 7 3 14 9 2 1 15 0 15 13 2
1 11
6 9 9 3 1 9 9
2 11 11
29 1 10 9 15 13 1 0 9 9 11 9 1 9 2 11 11 2 15 1 9 13 9 9 9 2 9 0 9 2
32 1 0 9 13 1 0 9 1 9 1 9 0 9 1 9 1 10 9 7 10 9 2 0 9 2 13 10 9 3 3 3 2
32 13 15 2 16 9 9 13 3 0 2 16 4 15 13 3 13 2 15 13 1 0 9 13 3 0 9 10 9 2 9 9 2
30 15 9 0 9 7 10 9 1 0 9 7 9 9 15 3 13 13 2 13 15 3 1 0 9 2 15 13 9 9 2
39 7 3 2 15 13 13 2 3 2 1 10 9 2 3 14 1 15 9 2 9 2 1 0 9 2 13 1 0 9 2 2 15 3 9 13 7 13 9 2
7 15 13 10 0 9 9 2
7 10 9 13 9 0 9 2
24 13 15 2 16 0 9 9 12 2 15 9 13 2 13 3 3 3 16 15 2 1 15 13 2
17 13 9 9 9 3 3 1 15 2 16 15 0 9 13 1 9 2
17 7 3 3 13 3 0 9 2 3 15 2 15 13 9 2 13 2
11 10 0 9 15 3 3 13 1 9 13 2
21 3 15 7 13 2 10 9 4 13 13 9 2 9 2 15 4 13 1 9 13 2
12 10 9 2 16 1 9 0 0 9 2 13 2
15 7 3 1 0 9 3 0 9 2 13 9 3 9 9 2
6 13 3 10 0 9 2
50 1 12 2 0 9 1 9 1 11 2 15 15 13 3 16 12 9 2 15 13 14 1 12 9 2 1 0 9 14 12 9 0 9 9 1 9 2 2 3 1 9 1 9 4 13 7 9 1 9 2
11 15 15 13 3 7 9 1 11 2 11 2
25 1 9 0 9 1 0 9 1 0 9 1 9 9 4 7 3 10 9 3 13 0 13 1 9 2
14 1 12 9 0 9 11 2 11 10 9 3 3 13 2
18 13 2 16 4 9 13 13 1 9 2 16 4 3 13 13 0 9 2
32 3 13 2 16 9 9 15 2 16 13 2 1 0 9 2 3 3 10 0 9 2 13 3 3 13 10 0 2 0 2 9 2
14 0 9 15 1 9 13 0 7 1 0 0 9 9 2
30 1 0 9 13 11 2 11 3 2 1 9 2 12 2 1 10 9 2 16 9 9 13 9 2 7 15 9 0 9 2
17 9 2 0 9 9 2 9 2 13 9 0 2 3 0 0 9 2
12 1 0 15 13 15 2 16 13 0 0 9 2
14 4 13 1 9 7 9 7 13 15 0 14 12 9 2
30 0 1 9 13 12 9 2 0 13 9 2 9 2 9 0 9 9 2 0 15 13 1 0 2 0 9 7 1 9 2
17 9 13 13 9 2 15 13 0 9 9 9 9 9 1 9 9 2
26 1 11 2 11 9 0 9 1 11 1 9 12 2 9 13 9 0 9 9 2 15 13 0 1 9 2
6 9 3 13 1 11 2
23 1 9 11 2 11 13 9 9 3 2 16 15 9 7 9 13 1 15 2 3 1 11 2
25 3 7 13 9 2 3 13 11 2 7 14 11 2 9 1 3 0 9 9 9 2 12 5 2 2
28 1 9 9 0 9 0 12 7 3 9 15 13 2 16 9 13 1 11 0 3 1 15 2 16 15 13 9 2
11 7 7 15 3 9 9 1 10 9 13 2
8 3 15 7 13 9 16 3 2
10 3 9 10 2 9 14 1 9 9 2
19 9 3 9 2 7 15 2 2 1 9 9 9 15 7 13 3 3 0 2
3 9 1 9
5 9 1 9 11 11
2 11 11
34 16 4 15 15 1 15 13 9 0 9 1 9 9 2 13 4 13 9 2 16 15 15 15 3 13 7 13 15 7 4 3 15 13 2
25 1 9 4 15 13 1 9 9 2 3 3 3 13 11 11 1 9 9 7 9 2 15 13 9 2
19 7 16 0 9 3 13 2 3 2 9 1 0 0 9 7 0 9 0 2
17 9 2 12 1 11 13 9 0 9 7 9 11 11 7 11 11 2
22 0 7 3 0 9 2 1 15 1 10 9 13 0 9 3 3 1 0 9 13 9 2
6 13 15 12 0 9 2
16 10 9 7 9 15 3 7 3 1 0 9 13 2 13 0 2
13 0 1 15 13 3 3 2 0 9 9 7 9 2
28 9 11 11 13 13 9 15 2 3 15 10 0 9 1 0 9 7 9 13 13 1 9 2 15 9 13 3 2
35 9 2 11 1 9 1 0 7 0 9 1 11 13 1 0 9 1 9 11 2 16 4 15 13 10 9 2 1 15 13 3 1 12 9 2
12 9 2 15 13 15 3 2 7 15 2 9 2
14 3 13 1 11 7 13 1 9 16 9 9 1 9 2
22 3 1 11 2 11 7 11 2 11 13 9 9 1 9 2 15 13 1 10 0 9 2
30 10 0 9 13 7 9 0 9 2 7 16 15 13 13 3 0 2 3 3 15 3 1 0 9 1 15 10 9 13 2
13 9 2 11 13 3 12 2 9 12 1 0 9 2
22 16 4 15 10 9 2 1 15 3 16 9 1 15 13 2 13 7 1 9 10 9 2
10 13 13 1 9 1 9 1 0 9 2
17 7 16 15 13 1 11 9 12 2 9 12 2 13 15 12 9 2
2 0 9
5 9 9 1 0 9
2 11 11
20 11 2 0 9 2 15 15 13 1 0 9 2 13 9 9 3 1 0 9 2
18 1 0 12 7 12 9 9 15 0 9 3 13 1 0 9 0 9 2
12 3 15 13 10 9 0 9 7 9 0 9 2
19 0 9 11 13 14 0 0 9 1 10 9 2 7 7 9 10 0 9 2
11 14 3 1 0 0 9 15 13 1 11 2
8 10 9 13 1 11 3 0 2
15 13 15 3 1 9 7 9 2 15 13 3 0 7 0 2
18 9 9 7 9 11 13 10 1 9 9 0 9 9 1 0 9 9 2
23 11 15 3 13 10 0 9 3 3 3 0 9 2 10 9 13 3 0 1 0 9 11 2
19 9 9 11 15 13 1 9 1 9 9 7 9 2 3 1 12 9 9 2
16 3 0 0 9 11 13 14 1 0 9 0 1 0 9 11 2
24 9 0 7 0 9 3 13 13 15 1 9 1 0 9 0 11 2 11 2 0 11 7 11 2
19 0 9 3 9 9 0 9 13 7 9 0 9 0 7 0 9 7 9 2
15 3 15 1 15 13 9 0 0 9 1 0 9 0 9 2
26 13 15 3 1 0 9 1 0 9 2 1 9 11 1 11 1 0 11 2 1 0 9 7 1 0 11
3 0 0 9
24 0 9 0 9 1 0 9 4 13 9 9 1 9 1 9 0 9 7 3 1 0 0 9 2
13 1 0 9 4 0 9 11 13 1 9 0 9 2
14 1 0 0 9 0 11 15 13 0 0 2 0 9 2
15 16 1 0 9 11 13 0 9 2 11 13 9 0 9 2
10 13 15 1 0 9 0 9 9 9 2
15 10 9 1 0 9 9 13 0 10 0 9 1 0 9 2
17 13 15 13 0 9 7 9 0 9 2 3 16 0 9 9 9 2
29 1 9 9 10 9 13 0 13 9 9 1 0 9 1 9 0 0 0 9 7 9 0 9 0 3 0 0 9 2
10 0 9 13 3 13 1 0 0 11 2
3 0 0 9
20 1 9 15 9 1 0 9 13 14 3 7 0 9 3 3 13 0 9 11 2
16 1 0 9 3 13 9 9 0 9 1 0 0 9 9 9 2
12 1 10 9 13 7 9 2 9 7 9 9 2
7 9 13 0 9 9 11 2
9 13 15 0 9 2 9 7 9 2
15 0 9 15 12 9 13 0 0 9 9 2 0 0 9 2
14 9 9 13 3 0 2 1 10 9 14 1 12 9 2
10 9 9 13 0 9 16 9 0 9 2
13 1 0 9 15 13 9 2 15 13 9 0 9 2
13 1 0 2 7 3 1 0 9 13 9 0 9 2
21 9 10 0 9 13 0 9 1 0 9 7 13 13 9 10 9 1 0 0 9 2
15 0 1 15 13 3 0 1 9 7 9 9 9 1 9 2
19 1 0 9 13 13 0 9 1 9 9 2 1 10 9 13 13 0 9 2
13 0 9 13 3 1 9 9 1 9 9 7 9 2
7 13 15 0 9 0 9 2
3 0 0 9
18 9 9 13 1 0 9 7 9 9 11 2 0 1 9 0 0 9 2
21 0 9 0 9 13 0 9 9 9 2 0 3 0 0 9 7 3 0 0 9 2
15 1 9 15 3 13 9 2 9 7 3 0 9 7 9 2
12 1 9 9 15 9 3 13 2 13 0 9 2
7 10 9 15 13 7 9 2
11 9 13 9 9 2 9 9 7 9 9 2
15 0 7 3 0 9 9 1 9 9 13 0 9 9 9 2
18 13 0 9 2 15 13 1 0 9 2 15 9 13 9 0 0 9 2
20 9 13 1 9 9 1 9 2 3 16 1 0 9 2 7 13 0 0 9 2
19 9 13 2 16 10 9 13 3 0 0 9 2 3 0 9 9 0 9 2
5 9 0 9 7 9
21 1 9 3 13 0 7 0 9 2 15 13 1 0 9 0 9 2 9 7 9 2
9 10 10 9 13 1 9 14 3 2
22 1 11 13 0 1 10 9 3 0 9 7 9 1 9 1 9 11 1 0 0 11 2
23 1 0 0 9 1 10 9 13 1 9 9 7 9 9 2 9 2 9 0 1 11 3 2
9 9 13 0 7 9 0 9 9 2
12 0 9 13 3 0 2 7 7 4 13 9 2
3 0 0 9
14 0 0 0 9 1 9 4 13 1 9 9 9 0 2
23 1 10 9 2 1 12 9 9 2 13 1 0 9 1 9 9 7 1 9 9 0 9 2
15 1 9 2 3 15 11 13 13 2 13 15 0 0 9 2
11 1 0 11 15 3 3 13 1 15 9 2
3 11 15 13
35 1 9 2 3 15 11 13 13 1 9 0 11 7 11 7 13 15 13 0 9 2 1 14 12 9 2 9 2 2 13 15 9 0 9 2
17 1 0 9 15 13 9 7 1 9 9 15 13 0 9 7 11 2
15 9 11 13 2 16 9 0 9 15 13 13 3 7 3 2
17 1 0 9 13 0 9 0 9 2 3 0 1 3 3 0 9 2
19 1 9 9 15 13 10 9 0 3 1 0 9 2 3 2 9 7 9 2
15 1 9 0 11 2 9 7 11 15 13 0 2 0 9 2
25 1 0 11 13 7 1 9 0 9 0 15 2 15 13 1 11 1 9 9 2 1 12 9 9 2
10 13 15 0 9 0 2 0 7 0 2
11 9 10 0 9 13 3 0 2 16 11 2
22 1 3 16 12 9 9 15 3 13 9 0 9 2 13 9 2 15 13 1 0 9 2
10 9 0 9 15 3 13 1 9 9 2
15 9 0 2 9 2 7 3 9 0 0 9 13 3 0 2
7 11 13 7 7 0 9 2
15 13 3 9 0 0 9 2 15 14 3 3 13 0 9 2
19 3 0 9 13 3 3 13 1 9 11 2 15 4 13 16 0 0 9 2
17 3 15 9 13 3 1 9 0 9 2 0 0 9 1 0 9 2
7 0 0 9 13 0 11 2
20 0 9 0 7 0 3 1 9 0 11 13 9 0 0 9 0 7 0 9 2
5 0 9 0 0 9
13 1 9 9 7 9 15 9 1 11 13 0 9 2
25 13 15 3 10 0 9 2 3 15 7 13 0 9 0 9 2 12 5 9 7 12 5 9 2 2
22 3 1 9 9 7 9 15 1 0 9 13 1 10 9 9 2 15 13 7 1 9 2
29 1 10 9 13 0 9 9 2 15 1 9 13 1 11 2 1 0 11 2 0 11 2 0 11 7 1 0 11 2
14 0 9 9 13 7 12 1 0 9 0 9 2 0 2
12 0 7 0 9 0 9 13 9 9 2 9 2
15 13 12 9 1 0 0 9 14 1 0 9 0 0 9 2
23 1 9 7 9 0 9 13 9 9 9 2 9 7 9 2 9 2 15 13 3 1 11 2
10 3 15 3 13 0 9 9 0 11 2
11 1 0 0 9 13 9 2 9 7 9 2
23 3 0 9 0 1 0 9 2 1 10 0 9 2 13 9 0 2 3 2 9 9 2 2
13 1 11 13 9 10 9 0 2 0 7 0 9 2
17 13 13 1 9 1 0 9 2 3 13 9 0 2 0 2 9 2
9 1 0 9 9 0 13 9 9 2
25 10 9 15 3 13 0 9 2 16 1 9 7 9 9 1 9 13 9 2 16 4 4 13 9 2
23 1 9 11 13 0 0 2 9 2 9 9 2 15 3 13 0 9 2 2 0 9 2 2
10 3 10 9 13 13 1 9 0 9 2
10 4 3 13 2 16 9 10 9 13 2
3 0 0 9
14 0 0 9 13 1 9 3 0 2 0 7 0 9 2
10 10 0 9 13 0 9 1 9 0 2
9 1 9 9 9 13 9 0 9 2
11 15 13 0 0 9 0 9 9 7 9 2
17 1 10 9 15 0 11 7 11 3 13 7 3 15 7 3 13 2
9 10 9 13 1 11 0 9 9 2
29 13 0 2 16 9 0 0 9 0 1 11 1 9 13 3 0 16 9 0 2 0 9 0 15 3 1 0 11 2
10 1 12 9 9 15 13 1 11 9 2
11 3 9 2 12 4 7 11 13 1 11 2
16 11 15 7 3 1 0 9 1 10 9 13 2 9 9 2 2
15 1 9 11 2 11 2 11 2 12 2 0 9 1 11 2
3 3 11 2
2 11 11
32 13 1 0 9 0 9 13 15 3 1 10 0 9 2 13 10 9 7 1 9 13 3 0 9 2 15 1 15 1 15 13 2
20 13 4 15 2 16 10 9 3 13 9 7 13 9 2 7 14 15 3 13 2
7 9 1 9 15 13 3 2
31 15 15 13 13 7 3 7 13 3 2 15 2 15 13 0 9 2 3 13 9 2 0 2 2 13 2 14 1 9 11 2
14 15 7 3 13 2 1 15 13 1 10 9 3 9 2
15 13 3 9 9 11 3 10 9 2 7 16 2 3 15 2
16 13 15 3 1 9 2 16 15 13 10 2 16 3 13 15 2
26 13 3 3 2 13 4 15 9 0 9 13 2 15 15 14 3 9 13 7 3 15 15 3 13 11 2
14 7 12 7 0 13 3 0 2 3 4 15 3 13 2
37 1 0 9 15 13 3 13 1 9 3 0 2 7 3 3 0 2 3 3 2 16 13 9 0 7 0 9 2 0 9 2 0 9 7 3 2 2
22 3 1 9 2 15 13 0 2 7 3 14 0 2 13 3 1 9 2 3 9 13 2
17 9 3 0 7 0 16 9 11 13 9 1 9 9 3 16 3 2
48 14 3 7 1 9 1 9 2 9 9 0 7 9 9 0 2 3 9 9 1 0 9 7 9 9 9 1 9 7 9 0 9 11 2 7 3 9 9 0 7 0 1 9 0 7 0 9 2
19 15 15 15 13 13 1 9 7 1 0 9 2 7 7 15 15 13 15 2
8 7 9 11 13 13 1 0 15
11 13 1 9 14 0 9 2 7 7 9 2
6 7 16 2 3 15 2
25 13 11 4 13 14 0 2 7 15 11 2 11 2 7 11 2 16 3 11 4 13 3 1 11 2
15 7 13 0 13 14 9 9 2 7 7 0 9 0 9 2
12 15 15 13 13 0 9 1 9 7 9 9 2
6 13 7 14 0 9 2
21 1 9 13 13 9 11 10 0 9 2 7 16 14 14 15 1 11 7 11 2 2
22 1 9 15 3 13 0 9 0 9 9 1 9 1 10 9 2 1 9 3 15 0 2
13 10 9 11 13 7 0 9 2 3 3 1 9 2
39 1 9 11 1 11 4 3 13 1 9 9 0 0 9 1 9 2 1 9 13 1 0 9 0 9 2 2 3 13 4 0 9 13 0 0 9 7 9 2
12 9 11 13 3 13 3 0 9 0 0 9 2
19 13 15 15 1 0 2 1 3 0 0 9 15 10 9 3 3 3 13 2
19 0 1 15 13 10 0 9 14 11 2 7 9 3 2 3 15 13 3 2
32 16 3 13 9 9 1 9 9 3 1 0 9 2 13 15 14 0 9 7 9 9 7 1 9 15 13 13 9 1 0 9 2
32 0 9 0 0 9 9 2 3 4 2 14 13 9 9 2 15 1 15 13 13 2 13 3 3 0 2 7 3 3 3 0 2
25 1 15 3 13 2 13 15 2 16 4 15 10 2 9 11 2 13 9 9 7 9 9 7 9 2
17 16 15 15 13 2 13 15 10 9 1 9 3 3 9 3 3 2
7 3 15 13 2 15 15 13
2 11 11
9 9 0 9 13 1 9 10 9 2
18 9 1 9 15 1 9 13 2 15 15 16 9 13 1 15 7 15 2
17 9 7 9 9 13 2 3 3 2 3 3 2 7 9 13 3 2
21 3 2 7 16 14 3 2 13 0 9 7 9 1 15 2 3 13 0 7 0 2
25 9 15 13 2 16 9 13 3 7 13 7 0 9 13 2 15 15 15 15 1 10 9 3 13 2
26 13 13 7 15 2 15 4 1 15 7 10 0 7 13 2 7 13 13 2 16 9 1 0 9 13 2
7 13 3 13 7 1 15 2
5 6 2 14 13 2
37 9 2 13 15 15 7 3 0 9 4 13 10 9 13 3 9 2 7 9 15 3 13 13 7 13 7 1 9 2 3 15 13 1 10 0 9 2
6 15 15 1 9 3 13
28 0 10 9 0 9 2 16 3 13 1 0 9 2 9 1 9 7 9 0 9 2 15 13 1 12 0 9 2
24 1 15 0 15 2 9 2 9 2 9 0 9 2 13 2 16 4 13 13 9 9 1 10 2
27 13 15 2 1 15 15 3 13 9 13 2 7 3 1 9 2 13 2 16 3 1 9 2 13 0 9 2
40 0 9 9 13 3 1 9 0 9 7 9 2 13 3 1 0 9 2 14 1 0 2 9 2 2 3 9 13 12 9 7 10 0 9 13 16 9 9 2 2
15 10 9 13 0 9 9 1 0 9 7 9 3 0 9 2
17 13 0 9 2 3 1 0 0 9 2 7 9 13 1 0 9 2
7 15 3 13 0 9 9 2
12 1 15 4 0 9 9 13 2 13 7 13 2
8 15 1 10 9 13 1 9 2
18 16 15 1 15 15 0 13 2 13 15 3 2 3 0 9 9 13 2
22 13 15 15 2 16 15 13 0 9 1 0 9 2 7 15 13 13 0 7 1 15 2
3 3 13 9
44 15 2 16 9 2 15 13 13 2 15 15 10 9 13 2 4 15 15 13 13 2 7 16 16 13 0 13 15 15 2 13 4 15 13 3 15 2 13 9 14 3 3 3 2
32 9 2 7 14 14 9 2 1 0 9 2 15 1 9 13 1 9 2 13 15 7 13 2 13 0 10 9 7 3 0 9 2
24 9 7 9 3 13 9 0 9 7 15 2 16 4 13 2 13 3 2 16 4 3 13 3 2
11 13 15 13 1 9 7 16 0 3 3 2
17 1 0 9 15 13 9 0 9 1 0 9 3 3 9 0 9 2
28 13 15 1 15 3 9 2 3 10 0 9 7 0 9 0 0 9 13 2 16 15 3 0 2 15 0 9 2
6 3 15 15 7 13 2
12 0 9 2 3 0 2 13 9 9 2 12 2
54 3 3 13 11 2 11 2 11 7 9 0 9 2 0 11 3 2 13 9 1 10 9 2 0 9 15 13 9 1 9 0 9 1 0 11 2 1 12 9 13 9 9 3 1 12 12 9 2 13 1 11 3 3 2
20 1 9 0 9 0 0 9 13 9 10 0 9 3 0 11 2 11 2 11 2
27 13 15 12 9 2 13 0 9 0 9 7 1 9 9 0 10 9 9 13 0 9 1 12 2 12 5 2
6 0 13 2 16 13 2
19 1 9 13 0 9 1 10 9 7 14 15 1 15 13 7 9 1 9 2
28 0 9 13 14 1 9 2 15 13 11 9 2 1 3 12 5 2 2 11 0 9 7 10 9 3 0 9 2
6 1 15 13 10 9 2
25 11 13 1 15 2 16 0 9 2 1 0 9 9 0 9 2 13 13 7 3 0 2 16 0 2
19 0 9 9 2 13 2 14 1 0 9 2 14 3 13 9 1 9 9 2
15 13 1 15 2 16 4 9 13 0 9 16 0 0 9 2
44 0 9 2 16 9 2 12 1 11 13 2 13 2 12 5 9 11 3 0 0 9 1 9 1 9 1 12 2 12 9 2 3 3 1 0 13 13 12 5 9 1 0 9 2
16 16 0 0 13 9 11 7 11 2 15 3 13 9 0 9 2
8 9 9 9 2 12 13 0 2
13 9 0 9 7 9 0 9 13 1 0 0 9 2
15 3 4 15 13 2 3 10 9 13 3 0 9 0 9 2
8 7 9 9 2 12 13 0 2
28 0 9 13 3 0 0 9 7 9 2 15 13 1 9 0 9 2 13 3 2 3 3 1 9 2 1 9 2
14 0 0 9 15 1 15 13 0 9 2 7 15 13 2
19 0 0 9 0 1 0 9 2 9 2 9 2 3 2 2 13 13 9 2
23 15 15 11 13 7 0 0 9 0 9 3 1 0 9 9 9 13 0 9 0 0 9 2
24 9 0 2 7 0 9 2 15 13 0 9 1 9 9 0 9 2 13 1 9 1 9 3 2
24 1 0 9 2 15 13 13 3 1 9 0 7 0 9 2 4 3 13 1 3 0 0 9 2
17 13 13 1 9 2 3 15 0 2 16 3 7 13 2 15 13 2
17 15 4 13 9 0 9 13 7 13 1 10 9 0 9 0 9 2
38 1 0 9 13 3 0 7 3 2 0 9 13 2 16 16 15 9 13 3 2 16 13 9 1 9 9 7 9 0 9 2 9 9 3 13 15 0 2
18 13 1 9 2 9 9 7 0 9 2 15 15 4 2 9 2 13 2
18 0 0 9 0 9 7 9 9 4 1 9 13 1 12 9 1 9 2
21 9 4 13 9 2 13 1 2 7 1 2 2 2 1 9 2 1 15 13 2 2
20 13 0 2 16 0 9 9 1 9 13 2 9 2 1 2 14 3 13 2 2
13 15 4 15 7 13 1 9 9 14 1 9 9 2
37 9 0 9 13 3 2 3 13 2 13 3 2 3 13 2 7 13 2 14 15 15 3 13 2 13 4 15 13 2 15 15 10 9 13 3 13 2
6 3 15 13 13 9 2
10 9 9 4 15 3 13 1 12 9 2
16 1 15 1 15 4 1 3 0 9 13 13 0 9 0 9 2
21 1 0 15 7 13 2 9 2 9 2 9 2 7 3 0 9 2 10 9 13 2
16 1 9 9 13 14 0 9 10 9 7 3 0 9 15 0 2
45 9 2 13 1 9 9 2 2 13 3 0 2 7 2 13 0 9 2 2 3 3 2 1 9 2 1 9 2 1 9 2 15 15 13 13 2 7 15 13 3 9 13 2 2 2
27 9 2 15 15 13 1 9 2 2 2 1 9 16 13 1 9 2 9 7 9 2 13 3 9 0 9 2
21 3 0 9 13 1 10 9 9 2 16 3 13 10 0 9 1 10 3 0 9 2
31 1 9 15 9 9 13 0 9 13 2 7 1 0 9 9 9 2 9 2 9 13 0 9 13 1 9 9 1 0 9 2
11 9 1 9 9 1 0 9 13 3 0 2
20 1 9 13 1 9 3 0 2 1 0 9 3 0 9 2 3 0 0 9 2
24 13 15 1 15 14 1 0 9 2 9 1 9 7 0 9 0 9 13 1 9 9 0 9 2
20 13 2 14 15 9 13 0 0 9 2 13 4 15 13 2 1 15 0 2 2
17 15 7 3 13 9 2 16 9 13 3 1 10 0 2 0 2 2
36 13 2 14 15 10 0 9 1 9 9 1 9 2 13 15 3 2 7 13 9 1 9 1 0 9 2 9 0 7 9 2 3 10 1 9 2
25 13 2 14 9 2 13 15 10 0 9 1 0 9 9 1 0 9 2 0 9 7 9 10 9 2
19 0 9 9 13 10 9 2 1 9 9 9 14 1 9 9 13 9 9 2
30 13 4 13 1 9 0 9 7 9 10 0 9 2 9 9 2 9 1 0 9 9 2 7 9 0 9 13 10 9 2
8 1 9 9 4 15 3 13 2
22 7 1 0 9 3 13 15 1 9 9 2 1 0 9 13 7 10 9 9 0 9 2
11 9 0 0 9 4 7 13 13 3 0 2
65 3 15 2 16 9 1 9 2 0 9 9 2 13 14 0 9 2 9 2 13 15 12 9 1 9 1 9 7 1 0 9 2 13 13 1 0 9 1 15 2 16 15 4 13 1 10 0 9 2 1 9 2 3 1 9 2 2 15 13 1 0 9 3 0 2
31 9 13 7 15 2 16 4 9 13 9 2 7 13 3 2 15 0 13 1 9 0 9 9 2 15 13 0 15 13 2 2
19 1 0 9 13 7 1 0 9 9 2 10 9 2 9 7 3 7 9 2
41 13 1 0 0 9 9 2 13 15 1 10 9 1 9 9 1 9 9 2 2 2 7 3 1 0 9 15 0 9 15 2 16 15 9 13 9 7 13 9 15 2
13 0 7 0 9 0 9 13 1 9 0 9 0 2
15 7 1 0 9 2 1 9 7 9 9 2 13 3 9 2
16 3 4 15 13 1 0 9 2 15 13 13 1 0 9 9 2
13 13 3 7 3 0 9 2 1 15 15 3 13 2
30 13 9 0 1 0 9 1 0 0 9 2 3 15 9 7 0 0 9 2 13 3 0 7 13 15 0 9 0 9 2
11 0 9 13 3 0 9 1 10 9 9 2
63 3 13 2 16 12 5 0 13 1 0 9 0 0 9 2 13 1 15 13 2 16 1 0 2 0 2 9 2 7 2 1 0 9 9 2 4 1 9 15 9 9 13 0 9 0 9 0 2 13 15 1 12 7 12 5 2 15 15 13 9 9 2 2
33 15 0 9 9 1 0 0 9 15 1 9 9 13 2 15 0 13 9 2 16 3 13 0 2 0 2 9 0 9 1 0 9 2
3 7 3 2
27 9 1 9 7 9 9 13 1 9 9 2 7 1 9 10 9 7 12 9 0 9 15 13 14 3 3 2
9 16 0 9 13 0 9 3 13 2
21 1 9 9 3 0 1 9 0 9 13 1 0 9 9 9 9 1 3 12 5 2
32 3 3 13 9 2 7 16 3 0 2 16 4 1 9 9 13 9 7 7 1 9 15 9 4 3 3 13 1 15 0 9 2
22 10 9 13 7 3 0 7 1 9 1 9 9 13 0 13 15 1 0 0 9 9 2
3 3 13 0
26 13 4 15 2 7 16 3 16 4 13 0 9 1 15 10 9 2 3 14 10 0 9 0 9 13 2
15 16 15 10 9 3 13 2 13 3 2 10 9 13 13 2
22 3 2 7 15 3 1 0 9 2 13 0 2 16 10 0 13 0 2 16 15 13 2
4 15 15 13 2
24 16 13 7 0 9 1 3 0 9 1 10 9 2 3 7 0 9 0 9 2 13 13 3 2
13 3 13 1 10 9 13 0 9 9 7 9 9 2
14 1 15 15 13 13 2 3 3 2 1 9 0 9 2
16 13 15 7 13 1 0 7 0 9 9 7 1 9 0 9 2
19 3 13 2 14 9 1 10 0 9 1 9 2 13 1 10 9 15 0 2
24 13 1 15 2 15 3 13 13 9 1 9 2 16 1 0 2 7 1 15 0 2 9 13 2
16 15 7 13 10 9 1 9 9 7 3 15 15 13 9 13 2
27 0 9 2 1 15 4 13 13 2 13 15 2 16 1 9 9 0 9 7 9 0 9 3 13 15 9 2
32 1 0 0 9 15 3 13 13 10 9 2 15 10 9 1 0 9 13 3 2 16 3 13 1 9 9 2 7 3 9 9 2
26 13 3 3 7 9 2 16 7 14 0 2 16 15 9 13 1 15 7 13 9 0 9 3 0 9 2
9 13 15 1 15 2 13 15 15 2
39 1 3 0 9 4 0 9 13 2 16 4 9 3 13 2 1 0 9 7 9 1 0 9 3 3 0 2 14 1 12 2 12 9 9 1 9 2 9 2
22 16 7 3 4 13 9 2 13 3 14 12 2 9 15 13 7 15 4 15 15 13 2
10 7 7 15 4 15 13 14 3 13 2
30 11 11 11 2 12 2 12 2 12 2 12 2 12 2 12 2 2 9 2 10 9 15 13 3 0 1 9 0 9 2
21 14 1 9 2 12 13 1 0 9 2 0 2 0 11 2 0 7 0 9 2 2
12 9 2 12 13 3 0 9 1 9 0 9 2
30 3 2 13 9 9 0 9 1 9 2 12 2 2 0 0 0 9 2 9 9 2 0 9 9 2 12 2 7 0 2
2 9 12
5 0 9 7 0 9
55 9 1 0 9 0 1 0 9 7 0 9 0 1 9 1 0 9 4 3 13 1 9 11 2 11 2 9 1 9 2 2 9 12 2 12 2 12 2 12 2 2 3 15 13 9 1 9 0 1 9 1 12 0 9 2
18 2 9 2 3 13 2 3 16 3 1 0 9 2 9 0 9 9 2
34 16 13 0 0 9 7 0 13 0 2 13 9 2 9 13 0 9 2 2 13 2 14 15 3 2 13 9 2 9 13 0 9 2 2
15 13 2 14 12 3 2 13 9 2 13 2 3 13 2 2
9 0 1 9 13 13 0 0 9 2
16 9 0 0 9 13 13 16 2 9 2 0 9 0 0 12 2
34 13 2 14 7 0 9 1 10 2 9 2 2 9 13 9 9 9 1 0 9 3 2 1 9 9 2 9 1 2 9 2 3 13 2
41 1 9 2 3 3 13 9 9 1 0 0 7 3 9 9 1 0 0 9 7 1 0 9 9 9 1 12 9 0 2 4 15 9 9 9 1 9 1 9 13 2
29 16 4 15 9 13 1 0 9 2 13 4 7 1 3 0 12 9 14 12 1 15 7 9 0 4 10 9 13 2
8 9 1 9 4 15 3 13 2
34 0 9 13 1 0 9 13 1 2 9 9 2 3 2 16 9 0 9 13 9 9 2 0 2 2 9 0 9 13 9 2 0 2 2
28 0 9 3 13 2 16 13 3 0 2 16 15 9 13 1 9 1 2 0 2 9 2 7 2 9 9 2 2
19 0 9 15 13 7 15 2 3 1 0 9 15 7 9 13 1 0 9 2
22 13 2 14 15 2 16 9 13 1 15 3 0 2 9 0 1 12 9 4 3 13 2
33 0 9 1 9 13 3 2 9 2 12 9 2 7 10 9 15 4 13 3 3 7 9 9 1 0 9 13 1 9 1 0 9 2
17 0 9 13 10 0 9 2 0 9 2 9 1 9 2 0 9 2
25 15 13 9 0 9 3 2 16 0 9 0 0 7 0 9 13 3 2 0 2 2 4 3 13 2
17 12 9 15 4 7 13 3 3 2 3 16 9 0 1 0 9 2
12 1 10 9 13 0 9 1 0 9 1 0 2
25 15 7 13 15 1 15 2 16 14 1 9 9 13 3 12 9 2 3 16 1 9 13 12 9 2
2 11 11
2 9 12
7 13 0 9 2 15 13 2
7 13 15 2 16 15 9 13
8 13 2 14 3 2 16 9 12
6 13 3 0 9 12 2
6 7 16 15 15 13 2
1 9
3 0 9 2
9 15 3 13 2 1 15 10 9 2
7 15 13 3 3 1 9 2
5 7 7 10 9 12
8 13 3 2 7 16 15 13 2
3 7 15 13
2 3 15
1 9
37 0 9 11 11 2 12 2 12 2 2 9 11 2 2 0 16 9 9 9 2 1 9 11 9 13 2 9 9 2 11 11 2 12 2 12 2 2
26 13 15 3 1 10 0 9 2 3 7 13 10 9 1 9 9 7 9 1 9 0 9 0 1 9 2
28 11 9 7 13 1 9 0 9 0 9 2 10 9 13 13 1 2 0 2 9 2 16 0 9 4 13 9 2
20 4 13 9 13 0 9 2 15 13 2 13 2 14 9 2 9 2 13 9 2
54 0 9 1 9 13 1 15 2 2 16 9 12 13 3 0 9 12 2 7 16 15 15 13 2 2 7 9 3 9 2 16 9 0 9 13 9 2 13 13 9 2 2 13 13 4 13 2 1 9 2 0 9 2 2
18 1 0 9 13 0 9 1 9 2 9 12 2 14 1 9 0 9 2
29 1 9 2 7 16 1 0 9 13 9 2 16 1 15 13 2 3 0 2 13 13 9 3 2 2 9 12 2 2
25 13 2 14 15 13 9 2 13 13 2 16 9 13 0 2 4 2 14 13 2 16 16 13 4 2
33 7 1 9 2 0 2 9 2 16 2 0 9 2 13 0 9 2 9 2 7 9 0 9 3 0 9 2 3 10 2 9 2 2
17 15 7 13 1 9 2 1 15 13 0 9 3 2 0 2 9 2
28 7 16 13 0 9 0 9 2 13 0 3 13 9 9 1 0 9 1 0 9 2 16 3 0 7 0 9 2
2 11 11
2 9 12
18 13 4 13 9 2 16 0 9 1 9 9 0 9 13 14 9 0 2
35 0 9 2 9 2 3 13 3 2 1 9 0 9 2 16 13 0 9 0 9 2 7 2 0 9 9 2 1 0 9 0 9 13 0 2
38 9 13 14 0 2 7 7 0 9 7 9 0 9 15 13 13 7 9 0 9 3 2 16 3 1 9 10 9 13 10 9 14 3 0 7 0 9 2
2 11 11
12 15 13 15 3 13 2 13 0 7 15 15 2
31 1 9 0 9 2 9 2 9 7 9 2 0 9 2 9 9 2 2 15 1 9 11 11 13 0 9 2 12 2 9 2
3 9 1 9
4 11 11 2 11
4 11 11 2 11
6 11 11 2 1 0 9
12 11 0 2 9 2 2 12 9 2 2 12 5
13 11 11 2 11 2 11 2 0 9 2 9 7 9
3 0 11 2
6 11 11 2 0 0 9
10 2 11 2 9 2 7 0 0 9 2
12 0 11 1 11 11 2 12 9 2 2 12 5
23 1 12 9 13 1 9 0 9 0 9 0 9 11 11 0 9 0 16 2 0 9 2 2
23 13 15 9 0 1 0 9 3 1 0 9 2 0 9 0 9 2 9 7 9 1 9 2
23 9 13 13 3 2 16 1 9 9 0 9 0 9 13 9 2 9 13 9 7 13 9 2
18 9 13 2 3 13 9 9 1 9 9 2 16 4 15 13 1 9 2
8 1 0 9 15 9 13 0 2
13 0 9 13 2 16 9 13 7 0 2 7 0 2
8 9 15 7 13 2 7 13 2
20 7 0 9 15 3 13 1 2 0 2 9 0 9 2 1 15 13 9 0 2
31 1 0 9 9 13 10 9 3 0 2 16 15 13 9 2 15 1 0 9 13 13 9 7 13 2 3 1 15 9 13 2
22 1 10 9 2 2 1 9 2 0 9 7 0 9 13 13 7 13 2 2 13 11 2
16 0 9 2 16 9 13 2 13 0 9 7 0 2 7 0 2
19 11 15 13 2 16 10 0 9 13 2 16 1 0 9 13 15 3 0 2
25 7 15 0 2 16 10 9 13 1 10 0 9 1 9 2 1 0 9 2 15 13 9 2 12 2
24 0 9 2 0 9 0 9 2 13 9 0 9 9 2 9 2 9 2 1 0 9 1 9 2
23 1 9 0 9 4 10 9 13 16 10 9 9 2 0 9 2 7 16 9 1 0 9 2
10 0 9 7 13 15 3 9 10 9 2
16 3 13 0 1 2 0 2 9 13 0 9 7 0 9 9 2
13 16 13 9 0 9 9 2 1 15 13 10 9 2
13 15 13 9 2 15 13 9 3 1 9 0 9 2
58 9 10 0 9 9 4 3 13 9 11 11 2 15 13 2 16 9 0 9 13 2 0 2 9 2 7 13 9 2 1 15 13 0 9 1 9 0 0 9 9 2 3 2 9 2 16 0 9 13 4 13 1 9 9 1 9 9 2
24 16 0 9 9 13 10 9 9 15 10 0 9 9 2 3 2 9 15 0 9 1 15 0 2
30 16 9 13 9 2 0 9 2 13 2 2 15 0 9 14 1 12 4 13 7 9 13 1 0 9 1 9 7 9 2
10 1 9 0 0 9 13 9 3 0 2
21 0 9 13 14 9 0 9 2 7 0 9 2 0 9 2 9 2 9 7 9 2
56 16 9 13 9 2 0 9 2 15 13 9 12 0 9 2 12 2 1 15 15 9 3 13 7 9 13 3 1 9 2 7 0 2 1 15 15 3 13 7 9 15 13 1 9 2 2 13 7 9 13 7 0 2 7 0 2
21 13 15 13 2 16 1 0 9 7 1 9 9 13 9 9 13 15 3 3 0 2
18 9 13 1 9 1 15 2 3 13 9 2 16 4 15 13 9 9 2
25 9 2 15 10 9 13 2 13 2 16 13 0 9 2 16 13 9 7 0 9 2 16 13 9 2
20 10 0 9 13 14 15 2 16 13 0 9 7 9 9 2 9 9 9 3 2
10 16 4 15 13 2 13 4 9 13 2
12 10 9 1 9 3 13 10 9 10 0 9 2
17 7 9 1 0 9 13 0 9 2 3 3 13 0 9 11 11 2
35 1 9 12 1 0 9 1 11 2 1 11 2 11 13 2 16 0 9 13 0 2 16 3 13 13 3 2 16 15 13 0 13 0 9 2
22 16 9 13 9 7 16 0 9 13 2 9 13 0 9 2 3 2 9 7 9 2 2
16 10 9 2 15 13 0 9 0 9 2 13 9 1 0 9 2
18 16 3 9 9 13 9 2 16 4 13 2 9 13 1 10 0 9 2
7 3 2 11 0 9 13 2
8 13 2 16 0 9 13 0 2
45 13 13 0 9 2 2 0 0 2 2 2 15 2 16 4 13 2 13 9 13 9 0 9 3 3 16 9 1 9 2 4 3 13 0 0 9 2 4 3 13 9 9 0 9 2
15 11 13 7 12 9 13 9 9 2 16 4 12 0 13 2
28 1 9 13 10 0 9 2 3 16 15 13 13 10 9 1 0 9 1 9 2 15 13 13 0 1 9 10 2
18 13 2 16 13 9 1 12 1 12 0 9 2 13 11 9 2 12 2
34 16 13 2 16 13 0 9 2 16 9 13 1 12 7 0 9 2 13 15 0 9 2 16 9 13 3 1 12 2 7 1 0 9 2
21 3 15 9 13 3 2 16 0 9 13 2 16 9 13 0 9 9 1 12 9 2
10 13 3 3 1 12 9 2 7 13 2
28 2 7 16 13 1 0 9 2 13 13 2 16 9 13 3 0 2 7 0 2 2 13 15 1 15 3 11 2
5 11 15 7 13 2
34 13 2 16 9 1 12 9 2 9 1 9 2 9 1 12 1 9 2 13 1 9 13 15 1 9 2 15 0 9 13 0 0 9 2
27 0 9 1 9 9 15 3 13 1 9 2 15 3 2 3 13 9 7 13 0 9 9 2 16 13 9 2
39 1 9 9 10 0 9 13 4 13 1 9 0 9 9 2 9 9 2 9 2 1 15 13 9 2 10 9 1 10 0 9 2 15 13 0 9 7 9 2
7 10 9 4 13 3 9 2
14 7 1 0 9 2 1 0 9 2 13 3 0 9 2
5 9 13 9 9 2
9 0 9 13 4 3 13 1 9 2
11 7 9 13 3 9 0 7 0 2 2 2
36 0 9 10 9 13 1 9 2 9 2 2 15 9 2 3 2 9 0 9 2 13 9 0 9 7 13 0 9 0 2 13 1 9 3 9 2
30 14 16 15 11 1 10 9 13 3 13 2 15 7 15 13 15 2 9 2 2 10 0 9 13 3 0 16 10 9 2
12 0 9 9 2 9 2 13 13 1 9 9 2
14 1 0 9 15 0 9 13 2 16 15 13 1 9 2
21 9 9 2 15 13 9 2 13 9 0 9 2 7 7 13 1 9 7 9 9 2
25 1 10 9 13 14 0 9 1 9 2 16 9 9 13 1 9 2 16 1 9 9 13 0 9 2
28 15 4 15 13 2 16 9 1 10 0 9 2 3 0 9 13 3 0 2 4 13 13 0 9 3 0 9 2
38 1 9 9 0 9 0 9 13 9 3 0 9 7 1 0 9 3 3 0 9 2 15 13 0 9 1 0 9 7 13 15 9 1 0 9 7 9 2
30 10 3 0 9 13 0 9 9 2 15 1 0 9 13 2 16 9 12 2 9 13 9 2 0 9 2 9 0 9 2
21 13 15 2 16 11 7 10 9 3 16 0 0 0 0 2 11 13 9 9 0 2
58 3 0 13 9 2 16 13 9 1 0 9 7 0 0 9 2 9 2 15 13 9 1 9 11 11 2 9 2 10 9 13 2 16 2 9 0 9 13 0 9 0 9 2 2 16 0 9 13 9 9 2 3 13 2 16 13 9 2
33 3 2 9 13 9 0 9 0 1 9 1 12 2 9 2 16 0 9 13 0 9 2 0 2 7 0 9 2 0 2 16 9 2
11 13 15 2 16 9 9 3 13 1 9 2
13 3 15 3 13 2 16 9 9 13 1 0 9 2
21 11 13 2 16 0 2 9 7 10 0 9 2 13 9 2 7 7 9 15 9 2
38 11 11 2 15 13 9 2 3 13 9 0 9 11 11 9 2 15 13 9 2 0 9 2 9 2 12 1 0 9 16 2 2 9 0 9 13 0 2
14 14 13 10 9 2 7 1 0 9 15 7 13 2 2
20 11 13 2 16 13 10 9 2 16 9 13 0 7 0 9 2 3 15 13 2
44 3 16 13 9 9 0 9 2 13 2 13 4 15 13 1 15 2 16 15 9 13 1 0 9 2 2 1 0 9 2 1 9 9 7 9 2 15 13 10 0 9 1 9 2
13 2 0 9 2 9 0 9 13 9 1 0 9 2
35 0 9 9 2 0 9 11 11 9 2 13 0 9 3 9 11 11 11 2 15 9 2 9 0 0 9 2 3 13 9 2 0 9 2 2
16 11 11 2 0 9 7 9 9 2 9 7 0 0 9 2 2
16 7 11 2 15 13 11 1 9 9 2 9 1 0 9 2 2
34 10 9 13 0 0 9 2 0 9 15 13 2 1 0 9 2 15 15 0 9 7 0 9 13 13 1 10 9 2 9 9 2 2 2
19 13 15 2 16 15 13 1 9 9 2 16 7 9 13 15 0 16 9 2
15 16 9 7 9 15 13 13 12 0 0 2 9 2 2 2
5 9 10 9 13 2
12 1 0 13 9 11 11 2 1 0 9 2 2
44 11 2 9 12 9 2 13 0 9 1 9 2 9 1 9 2 2 9 2 9 2 2 0 9 2 0 9 2 9 7 9 2 15 13 0 9 2 16 13 1 9 10 9 2
18 10 9 13 3 3 9 2 16 15 15 13 13 1 15 7 1 15 2
23 11 13 2 13 15 1 0 9 2 1 15 2 3 13 2 3 3 13 13 9 1 0 2
9 13 9 0 9 2 16 13 9 2
6 3 13 9 9 9 2
12 3 13 11 0 9 1 13 1 9 0 9 2
39 9 2 12 0 9 11 11 13 2 16 16 0 9 7 9 2 0 1 10 9 13 9 2 13 9 0 9 2 3 13 10 9 13 0 9 1 0 9 2
30 1 0 9 13 13 2 3 16 0 9 2 11 2 15 13 15 0 2 10 9 2 2 16 13 9 0 2 7 0 2
12 1 0 9 13 3 0 9 9 9 9 13 2
24 7 15 3 2 16 15 13 0 9 1 9 2 3 0 12 9 13 4 3 13 1 9 9 2
64 3 13 9 11 11 7 11 11 2 10 9 13 0 9 2 9 9 13 13 1 15 2 16 15 13 3 0 2 2 16 15 9 9 15 9 2 15 3 13 7 4 13 2 15 9 2 15 3 13 7 15 13 2 4 3 13 1 12 0 9 0 9 2 2
18 16 2 0 9 2 13 10 9 2 13 10 9 0 9 9 9 0 2
27 16 11 3 9 13 2 7 13 2 16 10 9 13 2 16 15 11 13 2 11 15 13 1 10 0 9 2
20 13 2 16 2 0 9 9 2 13 15 2 13 3 1 3 0 9 0 9 2
38 13 3 2 9 9 13 3 1 9 3 1 15 2 15 13 2 1 2 7 3 1 15 2 15 13 3 1 9 9 2 2 15 13 0 9 1 9 2
24 1 10 9 13 1 0 1 1 12 0 9 1 0 1 0 9 0 0 9 13 15 7 14 2
17 11 13 3 3 1 9 9 13 15 1 0 9 16 13 1 9 2
53 2 10 0 9 9 13 2 16 9 15 13 13 1 0 7 0 9 7 16 0 9 9 2 16 13 9 2 13 15 0 16 0 9 0 15 9 2 15 15 3 13 7 13 3 13 15 15 1 0 9 9 2 2
19 10 9 13 9 9 0 15 13 9 0 9 1 9 1 9 7 1 9 2
6 3 9 15 13 13 2
33 0 2 7 16 3 0 9 9 13 9 0 9 12 2 9 2 13 0 7 0 9 11 11 2 2 0 9 2 9 7 9 2 2
17 1 9 0 9 15 11 13 1 9 2 13 15 15 1 9 2 2
42 13 1 9 2 16 3 2 7 16 9 13 9 9 11 11 2 9 0 9 2 15 9 13 9 0 9 2 10 9 2 16 13 9 9 1 9 7 9 3 0 9 2
25 11 13 1 9 15 2 15 15 13 2 0 9 2 2 9 0 9 1 0 9 0 9 0 9 2
8 2 13 9 9 1 0 9 2
14 0 9 1 0 9 13 0 1 9 7 1 9 2 2
38 3 13 2 11 13 2 16 0 0 9 1 0 9 2 1 9 1 9 2 4 13 0 9 7 16 7 15 3 0 2 16 13 9 2 0 9 13 2
30 0 9 1 0 9 13 3 9 1 0 9 2 10 16 0 9 0 9 7 0 9 10 9 0 1 9 1 0 9 2
15 9 0 9 1 10 9 13 0 9 2 16 13 3 0 2
26 15 13 1 9 2 16 9 15 13 1 9 0 9 2 14 16 13 13 1 9 9 2 3 0 9 2
24 16 0 9 13 1 9 0 2 15 2 3 11 13 2 13 1 9 2 15 3 13 0 9 2
10 1 12 9 9 13 0 9 1 0 2
14 16 15 0 9 1 0 0 9 13 2 13 0 9 2
24 0 9 2 0 9 13 0 9 2 7 7 0 9 2 15 13 3 0 9 2 13 3 0 2
7 9 13 3 1 12 9 2
12 13 0 2 16 3 15 15 13 2 7 3 2
32 7 15 2 16 15 9 1 0 9 13 1 0 7 9 1 0 9 1 0 2 13 11 7 11 13 12 0 9 0 9 9 2
12 1 0 2 3 13 9 1 0 7 0 9 2
19 12 9 4 13 0 9 2 7 3 13 15 1 12 2 12 2 12 9 2
15 1 0 2 13 0 9 9 15 2 7 13 15 9 15 2
14 16 9 13 1 10 0 2 0 0 9 2 13 0 2
6 16 14 2 15 13 2
13 9 15 13 13 10 0 9 1 9 10 0 9 2
8 3 14 15 13 0 9 9 2
21 9 13 11 11 2 9 9 9 0 0 9 2 11 2 9 2 7 0 0 9 2
15 0 9 0 9 15 13 9 0 9 0 0 9 0 9 2
23 0 9 13 3 2 0 16 9 2 0 9 15 13 1 0 9 2 3 0 9 10 9 2
12 9 10 9 13 0 2 16 3 13 10 9 2
8 0 9 1 15 4 13 9 2
16 13 2 16 9 0 9 1 9 13 15 2 15 15 13 13 2
8 0 9 13 3 9 0 9 2
12 9 0 9 13 0 2 16 3 13 9 9 2
26 11 13 12 10 0 9 7 13 0 9 2 0 0 9 2 1 15 15 13 13 9 9 1 0 9 2
15 10 9 13 0 2 2 16 15 13 2 13 1 15 2 2
9 7 11 3 13 1 0 0 9 2
49 13 15 1 9 13 0 0 9 7 13 1 3 0 9 9 0 9 2 1 15 13 3 0 9 0 9 13 3 2 16 4 15 9 13 9 0 9 7 16 4 13 2 3 15 9 1 9 13 2
13 9 2 3 15 15 11 13 2 13 0 2 2 2
21 3 2 13 14 10 0 9 2 7 0 9 0 9 2 16 4 3 13 10 9 2
28 15 1 10 9 0 9 13 3 2 0 2 2 1 15 2 16 1 0 9 15 1 15 10 9 9 13 13 2
17 7 1 9 13 15 2 15 15 13 2 3 0 9 15 9 9 2
19 16 15 9 13 3 0 9 2 13 15 9 9 1 9 7 0 9 13 2
15 3 0 9 13 3 3 3 16 0 9 2 15 13 13 2
18 3 13 0 9 3 0 1 9 7 9 2 3 13 3 0 1 9 2
9 7 1 15 13 15 1 10 9 2
24 10 9 1 9 15 13 2 16 0 9 7 10 9 0 9 13 0 3 3 2 16 13 0 2
41 10 9 4 2 13 2 1 9 11 11 2 0 9 9 2 9 7 9 2 2 1 15 9 13 9 0 1 9 0 9 7 9 0 9 2 9 9 12 9 2 2
52 11 15 3 2 13 2 2 13 15 14 9 9 2 16 9 13 2 0 2 9 1 9 9 7 9 13 2 0 2 9 1 9 9 3 7 12 9 13 1 15 2 16 2 13 2 13 13 9 9 2 2 2
4 11 13 14 2
22 0 9 13 4 13 9 2 7 3 13 9 1 9 0 9 9 7 1 3 0 9 2
15 10 9 13 0 9 2 13 0 9 2 7 7 15 13 2
19 9 1 9 1 0 9 13 2 3 15 13 0 9 2 15 13 4 13 2
13 13 9 2 15 13 4 13 2 16 13 9 13 2
17 0 9 13 3 9 2 3 9 13 10 9 13 0 9 7 9 2
58 0 9 13 2 16 0 9 13 3 0 7 0 14 3 2 16 2 3 15 0 0 9 13 2 9 13 9 2 7 3 2 16 13 9 2 1 0 9 2 1 0 9 14 1 0 9 2 15 2 13 15 13 2 13 13 16 9 2
19 0 0 9 13 0 9 9 3 3 16 0 9 2 0 9 9 0 9 2
36 11 13 2 16 9 2 16 0 9 13 0 9 2 13 13 9 0 2 7 9 13 9 1 0 9 4 3 13 0 9 2 7 4 13 3 2
29 1 9 0 2 16 2 9 13 9 2 2 13 9 0 9 1 9 2 7 0 9 15 13 10 9 1 9 0 2
14 1 9 13 9 10 0 9 3 2 16 15 11 13 2
14 13 14 1 9 0 2 3 9 13 9 1 9 9 2
15 1 10 9 15 9 3 13 1 15 7 9 15 3 13 2
20 1 0 9 13 3 12 9 1 9 2 10 9 13 0 7 10 9 3 13 2
28 1 0 2 10 0 9 2 9 7 9 13 0 9 2 10 0 9 13 13 9 0 9 1 12 9 1 0 2
8 3 13 15 0 9 1 9 2
20 3 13 11 2 13 0 0 9 2 15 13 9 9 7 9 9 13 1 9 2
18 11 7 0 9 9 15 3 13 13 10 9 2 16 4 10 9 13 2
33 7 13 15 2 16 10 9 4 13 10 0 9 2 10 13 0 9 2 15 2 3 15 13 2 13 2 16 9 9 13 10 9 2
26 13 2 16 4 4 13 2 16 1 9 0 9 9 2 9 2 4 3 13 1 10 0 9 1 9 2
7 11 13 10 9 3 3 2
36 2 1 15 10 0 9 3 0 7 0 9 13 1 15 2 16 13 1 9 16 1 0 0 9 2 1 15 15 9 13 0 0 2 9 2 2
8 7 15 13 3 16 14 9 2
42 9 0 9 13 2 16 1 15 9 3 13 9 7 2 2 2 9 2 16 13 9 0 9 9 2 13 0 2 16 15 13 1 9 9 2 15 3 3 13 2 2 2
17 13 0 2 16 0 1 0 0 9 4 13 9 2 9 7 9 2
28 9 2 16 0 9 13 3 0 9 9 7 0 9 2 2 2 2 13 13 0 0 9 1 9 10 9 2 2
41 1 10 9 13 13 2 16 4 13 1 9 0 9 2 15 15 13 2 16 4 1 15 0 2 3 3 2 16 9 1 10 9 2 0 9 2 13 3 0 2 2
14 9 3 13 10 9 7 7 0 9 13 0 1 9 2
19 16 0 9 13 2 16 0 9 13 0 2 15 15 13 1 0 0 9 2
5 10 9 13 0 2
36 9 2 12 12 0 9 2 11 11 2 11 11 7 11 11 2 13 9 0 9 2 15 3 13 9 2 1 15 15 13 13 2 0 9 2 2
25 3 13 2 10 9 13 0 9 9 2 15 13 9 2 16 0 9 13 3 2 16 4 13 9 2
26 16 7 9 9 13 3 0 2 13 9 2 16 15 15 13 10 0 9 1 0 9 2 3 3 0 2
8 13 13 3 1 9 9 9 2
34 15 13 2 16 9 13 0 0 9 1 0 9 1 9 13 0 2 16 0 9 13 0 9 0 0 9 2 0 9 2 9 9 3 2
24 7 0 9 2 9 7 0 9 2 13 9 9 9 2 15 13 1 9 13 9 1 0 9 2
27 9 10 9 13 15 2 15 1 0 9 13 2 7 3 9 10 9 15 13 13 3 1 0 2 0 9 2
21 16 13 9 10 9 0 2 13 2 3 13 0 9 9 9 13 1 9 0 9 2
11 9 13 0 9 9 1 0 7 0 9 2
19 13 2 16 13 9 2 3 0 9 13 1 0 1 9 3 1 0 9 2
15 9 15 13 7 9 2 9 13 3 7 0 2 7 0 2
20 7 3 2 1 9 1 0 0 9 7 0 0 9 2 13 10 9 0 9 2
9 9 9 13 13 1 9 9 0 2
15 3 9 13 9 0 9 2 16 0 9 13 3 1 9 2
17 13 15 3 2 16 0 0 9 4 13 0 9 3 1 0 9 2
31 7 13 2 14 1 9 0 9 1 0 9 2 3 13 0 2 16 16 9 13 9 0 9 0 2 13 15 9 15 0 2
28 3 2 9 9 0 9 2 15 9 13 10 0 0 9 2 13 13 2 10 9 9 7 9 3 13 1 15 2
5 2 13 11 11 2
1 9
4 11 2 11 2
16 9 1 9 2 0 11 9 2 9 12 2 9 2 12 2 12
4 9 1 10 9
8 9 12 2 12 2 12 2 12
8 9 12 2 12 2 12 2 12
55 0 9 2 7 16 15 15 0 13 2 13 14 3 0 0 9 2 7 3 3 7 9 9 2 9 7 0 9 2 3 15 15 13 9 9 7 9 2 15 13 1 3 0 9 0 9 7 13 7 1 0 9 9 2 2
44 13 9 2 16 0 0 9 13 3 12 9 7 12 9 2 15 13 0 13 2 3 16 9 13 2 16 0 9 13 3 12 0 9 2 15 13 7 13 1 9 0 9 2 2
41 2 0 9 2 0 9 13 0 2 0 9 7 9 4 3 13 1 0 9 2 7 16 15 0 13 2 9 9 3 13 9 10 9 2 16 13 1 9 0 9 2
36 0 13 7 2 0 2 9 0 9 2 1 0 9 15 1 9 13 9 2 1 0 9 9 0 7 3 15 1 9 13 9 7 0 9 2 2
47 1 0 9 1 9 9 2 0 9 13 3 0 1 9 0 9 2 3 13 7 9 2 0 2 2 13 2 14 1 15 15 2 15 3 3 13 0 0 9 2 7 13 13 9 1 9 2
7 7 13 7 9 0 9 2
10 15 2 10 0 9 15 3 7 13 2
38 3 15 2 16 15 2 3 0 2 0 9 2 16 13 3 0 9 9 2 0 7 9 9 9 2 1 15 10 9 0 9 3 13 13 10 0 9 2
57 3 4 15 13 13 1 9 2 0 2 7 1 0 9 3 3 3 7 1 9 2 16 1 0 2 0 9 2 2 15 3 13 7 13 10 3 0 9 1 9 7 0 9 2 7 13 2 16 13 1 9 0 9 1 15 3 2
37 3 3 7 0 9 3 13 9 2 16 9 2 0 13 2 3 2 13 9 9 1 0 9 3 2 16 4 13 14 15 2 15 15 13 0 9 2
60 13 1 9 2 16 0 9 2 9 0 2 7 2 0 2 9 3 1 3 0 9 13 4 13 3 1 3 16 12 9 2 7 3 13 1 0 9 14 9 2 12 2 13 9 3 0 9 11 2 11 2 15 10 9 3 13 9 1 9 2
48 1 0 9 7 0 0 9 15 3 13 10 9 2 15 13 13 2 0 2 9 1 0 0 9 9 2 15 15 0 9 13 2 13 11 2 11 2 0 11 12 2 12 2 12 2 12 2 2
27 15 1 10 9 13 3 0 2 9 3 13 7 13 1 15 9 2 16 3 13 0 13 15 1 3 0 2
28 0 2 9 1 9 2 0 15 13 3 3 2 16 0 9 0 9 1 9 13 9 2 15 3 13 1 11 2
50 1 9 0 0 9 0 9 2 1 9 9 11 2 9 2 13 1 9 10 2 0 2 9 2 3 3 0 9 9 7 9 13 1 0 9 2 16 9 2 9 1 9 13 3 10 2 9 9 2 2
41 13 15 9 0 9 15 1 15 2 13 3 3 9 0 2 1 0 9 9 2 16 2 0 2 9 13 3 3 0 2 7 1 9 9 9 9 13 3 0 9 2
29 13 7 13 0 9 9 0 9 2 7 0 0 9 2 9 15 1 0 0 0 9 13 13 9 0 2 0 9 2
56 13 1 15 9 1 0 9 7 9 1 12 1 0 3 0 9 2 11 7 9 2 2 11 12 2 12 2 12 2 12 2 2 7 3 0 9 2 16 15 3 3 0 0 9 13 13 1 0 9 0 9 3 9 0 9 2
53 7 3 0 9 1 9 0 9 2 1 15 1 15 13 9 2 15 15 13 1 9 1 9 2 16 2 15 2 3 3 3 13 1 9 7 16 0 9 3 13 1 9 2 16 0 9 13 9 2 7 0 9 2
20 13 1 9 2 16 9 1 0 9 9 2 9 13 2 7 13 2 3 9 2
17 7 1 0 9 13 3 10 9 1 0 9 2 7 0 9 13 2
29 13 3 2 3 4 13 2 9 9 13 14 9 9 2 7 3 9 2 9 2 9 2 9 7 0 9 0 9 2
11 7 1 0 9 4 15 3 14 14 13 2
48 7 3 15 12 3 0 0 9 1 9 12 3 0 9 3 13 2 16 1 0 0 9 13 1 10 0 9 14 9 2 7 3 9 2 7 3 9 2 9 2 1 15 4 10 9 13 9 2
4 9 2 11 11
1 9
2 9 11
3 11 9 12
7 3 15 13 2 15 15 13
3 11 11 12
3 9 7 9
9 11 11 2 11 11 2 11 11 12
2 0 9
3 9 11 12
2 0 9
3 11 11 12
5 9 7 0 0 9
3 11 11 12
3 0 0 9
3 11 11 12
3 9 1 9
10 11 11 2 11 2 11 11 2 11 12
3 11 11 12
4 1 9 9 12
3 9 7 9
1 12
6 13 15 2 13 0 12
7 9 9 3 1 9 9 12
4 9 1 9 12
3 9 1 9
6 11 11 2 9 9 12
11 11 2 11 2 9 1 9 7 1 9 12
8 11 11 2 9 12 2 9 12
12 11 2 11 2 11 2 9 2 9 7 9 12
1 9
3 9 9 12
5 9 1 10 9 12
3 0 9 12
1 9
3 9 11 12
3 9 9 12
4 9 1 9 12
5 13 4 1 9 12
1 9
2 9 12
4 9 1 9 12
8 9 11 2 9 11 7 9 12
4 9 0 9 12
6 9 9 1 9 13 12
6 0 9 9 0 9 12
3 0 9 12
6 0 9 7 0 9 12
5 0 9 0 9 12
5 3 3 7 3 12
3 9 11 12
2 0 9
8 15 1 9 2 9 7 9 12
2 0 9
8 11 11 2 1 9 1 15 12
5 11 11 12 2 12
2 9 9
2 11 11
18 2 11 11 7 11 11 2 1 9 1 15 15 1 9 0 9 13 2
25 0 9 13 0 9 2 16 0 0 9 13 7 1 3 3 0 9 9 10 3 0 9 7 9 2
27 0 9 13 3 0 1 9 7 9 2 9 9 0 1 9 7 9 2 9 7 9 0 1 9 7 9 2
19 0 9 13 13 7 1 9 2 0 9 2 2 3 1 9 9 0 9 2
30 10 9 2 15 13 9 13 0 9 7 11 2 13 1 3 0 9 2 16 12 9 13 15 1 3 0 9 3 0 2
17 14 9 2 9 7 0 9 1 9 2 7 7 15 0 7 0 2
31 1 0 9 15 13 2 16 0 9 0 15 1 9 1 9 0 7 0 9 13 0 9 9 16 9 0 7 1 9 0 2
25 0 9 7 0 9 13 0 9 1 0 9 2 0 0 9 0 9 16 9 7 9 14 0 9 2
21 16 0 9 13 13 3 15 0 9 1 9 2 13 0 9 1 0 11 3 0 2
41 1 9 0 7 0 2 3 3 1 0 0 7 0 9 2 15 13 9 0 9 2 15 2 15 15 13 1 0 11 2 3 13 0 0 9 13 1 0 9 9 2
25 9 13 3 0 7 0 0 9 15 13 14 1 9 2 15 15 3 13 2 16 0 1 0 9 2
46 13 3 16 0 0 9 15 2 15 4 13 13 2 9 2 1 0 16 0 0 9 9 2 0 9 15 13 1 15 2 15 3 13 2 16 3 13 1 0 9 0 9 2 7 9 2
62 1 9 0 9 2 0 7 0 2 3 13 0 15 9 1 0 9 13 3 2 15 13 0 9 9 2 0 3 2 9 2 2 3 1 10 0 9 2 9 15 13 15 2 15 3 13 2 3 2 13 0 9 2 1 9 1 9 9 7 0 9 2
30 1 0 9 13 0 3 0 9 10 9 2 1 11 15 3 13 2 9 2 3 0 2 13 0 2 1 0 0 9 2
32 0 9 2 16 0 2 0 2 2 2 0 2 2 9 13 2 3 16 15 9 0 2 9 3 1 9 9 1 9 3 3 2
41 9 10 9 3 13 9 2 9 7 9 2 3 3 1 9 13 0 9 0 9 0 9 2 16 4 15 1 15 13 0 2 9 13 1 9 2 14 1 9 2 2
21 0 9 1 9 3 0 13 7 10 0 9 2 3 3 0 9 0 1 9 9 2
44 13 3 0 2 16 1 3 0 9 13 0 3 0 9 2 16 15 13 0 7 0 9 2 9 0 9 3 13 9 1 0 9 2 7 1 0 0 9 9 15 0 0 9 2
25 1 10 9 3 13 1 9 0 9 9 0 16 0 7 1 9 1 9 7 0 9 15 3 0 2
27 12 0 9 0 9 15 1 9 3 13 7 13 15 3 1 3 0 9 2 3 3 13 1 9 3 9 2
25 3 13 0 1 15 13 7 13 15 9 0 9 2 3 0 1 9 3 0 9 2 3 0 9 2
10 9 9 13 3 0 14 1 0 9 2
9 11 2 12 2 12 2 12 2 12
10 11 2 12 2 12 2 12 2 12 2
8 11 2 12 2 12 2 12 2
2 12 2
13 11 1 0 7 0 11 2 12 2 12 2 12 2
6 13 9 1 0 9 2
4 9 1 9 2
19 1 9 0 9 11 1 11 13 13 12 0 9 9 0 9 12 7 12 2
21 12 1 15 13 1 9 14 12 9 13 1 15 9 2 0 15 9 1 0 9 2
23 13 9 0 1 0 9 0 9 7 1 0 11 1 10 0 9 0 9 1 0 9 0 2
9 9 12 2 9 12 2 9 2 12
8 1 0 9 9 1 9 0 2
28 1 1 9 2 15 4 13 1 9 1 9 2 13 15 13 0 2 13 0 9 3 1 0 9 0 2 2 2
23 1 9 10 13 3 1 3 2 16 9 0 13 9 1 15 9 0 2 3 0 9 0 2
22 16 4 9 10 13 0 2 13 3 2 16 4 9 0 3 13 13 2 15 3 0 2
17 1 0 9 9 2 16 0 9 9 13 13 15 0 9 9 9 2
33 3 13 15 9 10 2 15 13 0 9 0 2 9 2 16 4 13 0 9 0 7 0 1 10 9 2 16 1 9 2 9 9 2
15 1 15 13 9 2 13 3 3 13 2 3 9 3 0 2
23 1 0 9 1 9 9 13 13 2 16 9 1 0 2 0 2 9 1 9 0 3 13 2
9 9 12 2 9 12 2 9 2 12
4 9 9 0 2
41 9 0 2 15 3 15 2 3 1 9 12 0 2 3 13 2 13 1 0 12 9 3 9 10 9 2 7 13 10 9 1 0 9 3 9 16 2 14 1 9 2
12 15 13 9 1 9 2 15 15 13 13 9 2
47 7 9 0 1 0 9 13 15 1 9 0 9 2 9 2 0 1 11 2 9 0 13 2 15 15 3 3 13 13 2 16 9 13 1 0 2 0 9 7 14 0 9 1 9 15 13 2
15 9 0 13 1 15 3 13 1 0 9 2 16 13 0 2
9 9 12 2 9 12 2 9 2 12
4 9 7 9 2
23 16 9 9 1 9 15 13 2 13 1 15 0 0 9 11 2 16 9 13 0 2 2 2
32 9 2 11 13 9 15 0 10 9 9 9 1 9 9 1 9 9 7 0 9 10 2 3 9 2 15 15 3 13 2 2 2
9 9 12 2 9 12 2 9 2 12
8 0 9 2 9 2 7 9 2
2 11 11
23 0 9 11 11 1 11 2 3 11 2 15 3 13 2 16 15 9 0 9 13 1 9 2
16 1 15 13 2 16 9 13 0 7 0 9 7 1 0 9 2
30 13 3 0 9 2 9 2 7 11 2 0 15 3 1 15 0 9 2 15 13 0 9 1 9 9 16 9 0 9 2
28 9 2 15 13 0 9 13 1 9 0 9 2 15 13 2 16 0 9 0 9 2 9 7 3 13 0 9 2
23 13 15 9 9 2 9 0 2 2 9 9 2 9 0 2 7 9 0 2 9 0 2 2
26 3 1 10 9 15 13 2 16 0 9 13 13 0 9 7 1 9 7 13 15 1 15 0 0 9 2
14 10 9 13 9 0 2 15 4 1 9 13 9 0 2
8 9 13 3 3 0 9 13 2
29 7 15 13 9 9 2 15 15 13 1 15 9 0 7 4 13 1 0 0 9 2 9 2 9 2 9 0 2 2
10 9 9 13 2 7 16 13 0 9 2
9 9 15 15 13 15 3 3 13 2
13 13 3 0 2 16 9 13 10 9 0 0 9 2
21 0 13 2 16 13 1 9 1 9 2 0 2 16 13 15 9 0 0 9 9 2
15 11 11 13 1 9 9 1 0 9 2 11 3 12 2 2
12 9 13 14 0 9 2 15 15 0 9 13 2
8 13 15 3 14 9 0 9 2
32 15 15 13 9 1 9 9 2 0 1 0 9 2 2 12 2 9 13 10 9 2 15 13 9 13 1 9 0 9 7 9 2
15 2 12 2 9 1 9 4 3 13 9 0 9 2 9 2
19 2 12 2 0 9 13 13 3 1 10 9 2 15 13 1 9 0 9 2
11 1 9 0 0 9 4 13 1 12 9 2
17 1 9 2 1 15 4 9 13 2 15 9 9 13 1 9 9 2
8 9 3 3 13 0 9 9 2
21 0 9 1 9 4 13 3 2 16 9 4 13 0 9 2 7 9 1 9 9 2
10 1 11 13 0 9 1 9 9 9 2
17 9 15 13 0 9 9 7 1 9 0 1 9 9 13 0 9 2
14 1 0 9 4 9 13 1 9 1 9 1 0 9 2
6 0 9 15 13 9 2
20 9 2 9 0 9 9 2 13 3 3 3 9 7 9 9 7 1 9 9 2
12 4 3 13 9 9 7 9 2 15 15 13 2
8 0 9 9 3 13 7 13 2
17 3 7 13 1 10 0 9 7 1 10 9 15 13 3 7 3 2
25 11 11 2 9 9 0 9 13 2 16 13 1 9 9 1 9 9 2 15 13 1 11 3 13 2
19 1 15 15 9 13 12 9 2 9 0 2 9 2 0 7 9 2 0 2
18 10 9 9 13 2 7 13 15 9 1 0 9 7 3 15 3 13 2
10 9 10 0 9 13 3 0 7 0 2
23 9 1 9 13 9 2 16 9 0 1 0 9 1 9 13 3 0 9 9 1 0 9 2
24 0 9 1 10 9 15 15 13 3 3 1 9 9 7 9 2 3 3 1 0 9 0 9 2
21 1 10 9 13 11 9 2 16 7 1 9 13 10 9 0 9 2 10 0 9 2
25 9 4 13 9 2 16 9 0 3 13 13 0 9 2 15 15 13 13 1 9 0 9 0 9 2
13 1 9 9 0 0 9 13 11 0 9 11 11 2
4 9 13 0 2
18 1 9 13 0 9 0 9 0 9 2 9 2 3 0 1 0 9 2
14 11 13 2 16 9 2 9 13 0 0 7 0 9 2
18 13 3 2 16 3 0 9 13 0 1 9 7 13 3 0 0 9 2
18 9 13 7 0 9 2 0 9 13 0 9 2 7 15 1 0 9 2
11 7 3 10 9 7 1 10 9 13 9 2
7 9 2 9 2 11 11 13
21 9 12 2 12 2 12 13 1 9 12 9 9 11 2 0 0 0 9 10 9 2
54 9 11 1 9 12 2 12 13 1 0 9 9 2 11 7 9 2 11 1 11 2 1 9 12 2 12 13 9 12 2 0 9 9 11 2 3 13 9 9 0 9 7 9 11 2 3 9 9 0 7 0 9 11 2
9 13 15 1 9 0 9 1 11 2
29 13 15 1 9 9 9 7 3 1 15 2 16 4 3 13 9 10 9 2 13 0 9 1 10 9 9 0 9 2
16 0 9 0 9 9 2 11 13 7 1 0 9 1 9 9 2
33 13 9 10 9 2 15 13 1 10 9 7 13 15 0 9 9 9 2 9 1 10 3 0 9 2 7 3 9 1 9 7 9 2
42 1 10 9 13 9 9 11 1 3 0 9 7 13 2 3 3 2 9 1 9 2 15 13 0 2 16 13 3 2 9 0 2 9 2 9 2 9 7 13 15 3 2
26 15 7 3 13 1 9 10 9 2 3 13 2 16 0 2 2 0 2 2 9 15 3 3 3 13 2
31 3 3 1 9 9 7 9 2 14 15 0 9 3 13 9 2 0 9 1 0 9 2 2 9 12 2 12 2 12 2 2
28 13 9 10 9 2 2 11 13 0 9 2 15 15 13 1 10 9 2 1 10 9 2 1 10 9 13 2 2
15 15 13 9 11 11 2 9 2 11 15 15 7 3 13 2
8 13 2 16 13 0 15 13 2
2 11 11
11 9 2 11 11 2 9 1 9 7 1 9
27 9 2 11 5 11 2 11 12 2 12 9 2 9 2 9 13 2 1 9 9 0 9 12 2 2 2 2
20 16 4 0 9 13 1 9 2 0 10 9 13 13 2 15 15 3 9 13 2
9 13 2 16 10 9 9 9 13 2
29 1 0 0 9 2 11 2 11 12 2 4 9 13 2 7 13 3 9 2 2 9 9 2 16 10 9 13 0 2
7 9 9 2 13 9 2 2
65 15 15 3 13 2 7 1 9 0 9 4 1 0 9 1 10 2 15 15 15 1 9 9 1 9 13 2 13 1 10 9 2 9 13 9 9 7 9 2 15 9 13 7 13 3 2 3 7 3 10 9 2 9 2 9 7 9 3 0 2 3 7 0 9 2
14 9 3 3 13 7 13 1 9 2 3 16 0 9 2
32 9 3 2 1 15 3 3 2 13 0 2 0 2 0 7 0 9 7 0 15 2 3 0 2 13 9 13 7 13 10 9 2
16 3 4 9 7 9 13 1 9 2 16 4 15 3 3 13 2
49 1 0 9 9 0 9 7 9 15 2 15 4 0 13 1 10 9 2 9 2 9 2 9 2 9 2 0 9 2 0 9 2 9 0 9 2 9 7 9 1 0 9 2 13 1 0 0 9 2
41 3 10 9 9 2 9 0 0 9 2 3 3 13 15 14 2 7 0 9 7 0 0 2 4 15 0 1 15 1 10 9 13 13 2 16 1 15 13 3 3 2
18 1 10 9 7 13 2 16 9 3 13 7 13 0 9 0 0 9 2
2 11 11
11 10 9 0 1 9 12 15 13 3 7 3
45 3 2 16 15 13 15 2 15 13 3 4 13 1 9 12 2 16 3 15 13 0 9 9 2 0 9 9 2 0 9 2 0 9 7 9 7 3 0 0 0 9 3 3 0 2
16 3 15 13 0 9 16 0 0 9 2 15 3 13 0 9 2
34 3 15 7 13 1 9 2 0 1 9 12 2 2 16 4 0 1 9 3 3 2 16 3 1 0 2 12 11 9 0 7 1 9 2
7 15 13 2 13 15 13 2
26 7 1 10 0 9 13 12 9 2 15 9 3 3 13 2 7 15 1 9 2 16 13 2 3 13 2
35 1 15 13 3 3 13 9 2 7 0 9 13 13 15 1 9 2 15 13 1 15 1 9 0 7 1 9 0 3 0 7 14 3 0 2
19 11 11 2 9 12 2 9 2 11 2 9 2 12 2 9 2 11 11 2
28 11 2 11 2 11 2 9 2 9 7 9 2 11 2 11 2 12 2 9 2 11 11 2 9 11 11 2 2
22 0 1 15 13 0 9 15 9 0 0 9 1 0 9 9 2 0 9 7 0 9 2
20 0 13 3 1 10 0 10 0 9 0 13 0 9 9 10 0 7 0 9 2
9 11 13 12 2 9 16 9 9 2
19 9 9 13 15 2 3 15 9 13 2 16 13 3 2 16 1 9 13 2
15 9 0 9 2 0 1 0 9 2 10 0 9 3 13 2
2 11 11
6 11 11 2 9 9 2
16 11 11 12 2 12 9 2 12 9 2 2 9 11 2 11 2
3 12 2 9
13 11 11 2 12 2 12 2 13 1 0 0 9 2
6 13 9 11 2 11 2
6 13 15 3 0 9 2
46 3 13 12 9 3 3 0 9 2 15 13 11 11 2 12 2 2 9 1 9 11 9 2 12 2 2 0 9 2 12 2 2 0 0 9 7 10 0 9 2 12 2 7 15 0 2
14 9 2 12 4 13 1 9 7 1 12 9 9 13 2
21 3 4 13 2 7 0 9 15 9 2 12 13 9 13 1 0 9 11 1 11 2
8 1 9 12 13 3 1 9 2
17 1 10 12 9 3 0 9 1 12 0 9 13 11 2 11 9 2
5 13 13 1 9 2
10 13 15 9 2 15 13 13 0 9 2
23 1 0 9 15 13 9 2 16 9 0 1 9 9 9 9 15 13 9 1 9 0 9 2
34 1 0 9 9 1 2 0 9 2 9 2 9 7 9 2 7 3 9 7 9 13 11 2 11 13 9 7 10 9 3 1 15 0 2
14 13 3 1 0 9 2 9 7 9 2 7 1 15 2
10 13 15 13 9 9 2 10 0 9 2
6 13 1 9 7 9 2
8 9 1 9 13 10 0 9 2
15 13 15 2 16 1 10 0 9 13 3 0 2 3 0 2
9 13 0 2 0 7 10 9 0 2
26 13 3 1 0 9 10 9 2 7 7 1 9 2 3 15 13 1 11 2 11 7 13 12 9 9 2
40 10 2 9 2 2 9 9 1 9 2 13 9 0 12 9 0 9 9 2 11 11 7 11 11 2 7 13 9 1 9 2 15 13 2 13 1 15 15 0 2
31 9 0 9 13 12 0 9 1 9 2 15 15 15 13 16 2 9 2 15 13 1 9 9 2 7 9 9 7 9 2 2
90 13 15 1 15 10 0 9 9 7 10 0 9 2 3 2 0 9 7 9 9 2 11 1 9 0 9 2 9 9 2 9 9 2 9 9 1 9 7 9 2 9 7 9 9 2 9 1 0 9 2 9 1 9 16 9 9 2 0 9 0 0 9 2 11 11 16 12 1 0 0 9 0 9 7 0 9 2 15 15 13 3 9 1 9 16 0 9 1 9 2
20 13 15 0 9 2 10 9 3 13 0 9 11 9 7 0 9 9 11 11 2
2 11 11
8 9 9 2 3 1 9 1 9
8 9 12 2 12 2 12 2 12
18 1 12 2 9 9 13 11 11 7 9 11 1 11 9 9 1 9 2
21 1 10 9 7 9 4 14 13 1 9 13 10 9 1 9 7 3 0 9 9 2
32 12 2 9 9 2 9 13 3 10 0 9 2 1 15 2 3 2 1 0 9 2 3 2 13 15 16 2 3 2 7 3 2
8 3 15 13 13 9 9 9 2
8 3 13 9 13 3 1 9 2
47 0 0 9 2 0 9 2 13 10 2 9 2 2 15 2 15 9 3 13 13 2 1 9 13 2 7 3 13 15 0 1 15 2 16 15 1 10 9 0 9 13 7 9 13 1 9 2
18 3 0 9 15 3 13 2 1 0 7 0 9 7 3 1 9 0 2
33 12 2 0 9 2 4 2 14 3 1 11 9 0 9 13 9 9 2 3 9 15 15 16 1 0 9 2 3 13 10 9 0 2
7 9 4 3 13 9 9 2
6 9 1 15 13 0 2
16 9 3 13 9 1 3 0 0 9 2 15 4 15 13 13 2
17 1 10 9 15 9 1 9 13 1 0 9 9 2 0 9 2 2
25 9 13 1 0 9 14 3 16 11 1 9 2 15 13 3 0 9 9 7 3 15 13 13 2 2
8 13 15 13 15 7 1 9 2
23 12 10 9 3 2 16 15 13 1 0 9 2 13 2 3 15 13 2 1 9 1 11 2
19 7 3 2 9 1 15 13 2 9 15 13 2 15 3 13 3 0 9 2
25 15 15 13 1 9 2 1 9 7 14 15 1 15 13 2 2 15 13 3 2 16 13 1 11 2
11 16 4 13 3 2 15 4 13 9 2 2
19 7 3 3 1 9 2 1 15 11 13 2 13 15 1 10 0 0 9 2
19 9 13 0 7 0 9 2 15 0 9 13 7 13 15 13 15 1 15 2
6 10 0 13 0 9 2
50 3 15 13 7 1 10 0 0 9 2 3 13 3 0 2 7 3 14 3 0 2 13 2 14 15 15 13 9 10 9 2 7 15 16 0 9 7 2 3 13 2 9 0 9 13 0 9 10 9 2
17 12 2 0 9 2 13 3 0 1 9 2 15 13 1 0 9 2
22 13 1 15 9 9 7 13 1 0 9 9 0 9 4 13 13 0 7 14 0 9 2
10 13 3 0 13 2 10 15 9 13 2
17 13 15 3 13 3 1 9 1 0 9 7 9 15 3 0 13 2
33 2 9 2 7 2 9 2 2 12 9 0 16 0 2 0 4 13 9 2 3 3 13 13 1 9 2 13 2 14 1 15 0 2
23 3 3 0 9 13 2 7 9 13 3 15 0 1 9 2 16 9 3 13 1 9 15 2
11 14 12 13 13 2 0 9 13 3 0 2
18 13 15 13 1 0 9 7 1 0 9 2 13 9 7 14 15 3 2
28 13 15 13 0 7 13 15 13 0 2 13 15 3 0 2 7 3 15 1 15 15 10 9 13 2 15 13 2
11 0 13 2 16 15 15 13 2 1 9 2
20 12 2 9 7 9 2 9 1 9 13 0 7 13 9 13 1 10 10 9 2
10 3 13 15 10 9 0 7 0 9 2
11 13 15 7 3 13 7 9 1 15 13 2
7 3 16 1 10 0 9 2
2 11 11
3 0 9 2
8 9 12 2 12 2 12 2 12
31 1 9 2 9 0 9 2 15 11 11 2 13 3 3 2 13 9 2 15 13 14 0 9 7 3 15 1 15 13 13 2
14 13 15 0 9 9 9 2 15 15 13 1 0 11 2
29 13 3 13 1 0 9 2 2 12 1 0 9 0 9 1 9 0 0 9 13 3 0 9 9 0 9 9 2 2
33 9 10 9 2 7 2 9 0 15 1 0 2 0 3 2 2 9 9 2 13 1 0 9 2 7 2 9 1 10 9 2 0 2
10 1 10 9 15 13 3 13 0 9 2
25 9 15 13 2 16 2 9 9 1 9 0 9 13 3 9 10 2 0 2 9 9 2 2 2 2
27 7 13 2 14 3 4 9 0 9 13 1 0 12 2 9 2 0 3 2 7 0 9 1 9 9 2 2
9 15 13 1 9 0 9 0 9 2
34 2 13 15 9 9 2 9 7 0 9 2 15 7 15 15 3 13 13 2 2 2 7 3 2 3 4 1 0 0 9 13 13 2 2
27 3 13 10 9 9 2 0 0 9 2 9 2 9 2 9 2 13 9 10 10 9 7 3 15 13 2 2
15 16 4 9 13 1 9 2 3 1 15 3 13 15 9 2
42 16 13 9 2 0 9 2 3 2 16 1 15 13 3 9 0 0 7 0 9 1 9 2 2 2 2 2 7 15 15 3 13 13 2 2 2 3 13 15 9 0 2
5 15 13 3 9 2
6 3 13 2 9 13 2
15 7 10 9 13 9 0 9 1 9 1 9 13 3 0 2
33 9 0 9 13 1 9 10 7 15 0 9 2 16 13 3 2 9 7 9 9 2 9 0 9 2 0 9 2 0 9 2 0 2
9 7 7 0 9 13 0 9 3 2
13 15 9 13 16 9 0 9 7 0 9 1 9 2
13 0 9 13 3 10 9 2 15 15 3 13 13 2
22 12 9 13 13 0 9 7 0 9 1 9 0 7 0 9 1 9 9 9 7 9 2
30 1 10 9 13 10 9 13 9 9 9 7 9 2 13 15 13 3 16 9 9 2 2 15 15 13 7 13 1 9 2
12 3 13 10 9 0 2 7 1 9 3 13 2
12 3 13 3 7 9 2 15 3 13 16 0 2
10 0 9 7 0 9 13 3 3 15 2
27 1 9 3 13 14 12 9 2 3 0 9 2 9 0 2 3 9 2 0 9 0 1 9 1 9 2 2
19 0 9 13 3 11 11 2 3 15 9 13 2 12 2 9 2 12 2 2
37 11 13 2 16 1 9 9 2 15 9 13 0 9 2 15 3 13 0 9 2 2 9 4 3 1 10 0 9 14 1 0 9 13 7 13 2 2
52 7 13 11 11 2 0 9 1 9 2 12 2 2 15 12 9 3 13 2 9 2 12 2 2 2 7 16 13 1 0 0 9 2 13 11 3 15 0 2 15 13 1 9 13 2 9 13 9 0 9 2 2
17 7 13 2 2 0 1 15 13 9 2 15 15 1 10 9 13 2
32 15 15 13 9 9 1 15 2 15 13 1 10 9 13 15 1 9 2 13 10 7 15 0 9 2 13 1 0 9 2 3 2
52 16 3 2 10 0 9 13 0 9 7 9 2 1 15 1 0 9 12 0 2 0 7 0 9 1 0 9 13 0 9 2 3 15 13 15 0 16 9 1 10 9 1 9 2 16 4 3 13 13 0 9 2
42 16 9 13 1 10 0 9 2 16 4 13 0 9 10 0 9 7 3 1 9 13 2 16 15 10 9 7 0 9 15 3 13 2 3 13 15 9 1 10 9 2 2
43 7 3 13 2 2 9 13 0 9 9 2 3 3 15 3 3 13 2 3 2 10 9 2 16 4 0 9 2 0 9 2 0 9 2 9 2 9 3 2 2 3 13 2
49 1 9 1 15 2 16 9 3 13 0 9 2 0 9 13 1 0 2 9 1 9 7 9 1 10 0 9 2 10 15 13 0 9 2 16 15 0 13 13 2 10 15 13 0 2 2 2 2 2
16 2 0 9 13 3 3 2 16 15 13 16 9 9 13 0 2
24 16 9 1 9 2 15 15 0 9 13 1 9 0 0 9 2 15 13 10 3 0 9 2 2
22 9 13 9 2 0 9 1 9 2 2 7 3 9 1 9 2 9 2 3 0 9 2
30 3 4 15 13 1 0 9 2 16 4 13 2 16 0 9 3 13 0 10 9 2 1 15 15 3 1 0 9 13 2
26 15 4 15 13 2 16 4 3 13 13 9 2 1 10 9 15 13 7 1 15 15 3 15 15 13 2
16 13 14 2 16 13 15 1 15 3 7 16 15 15 13 13 2
12 3 4 15 3 13 1 9 2 15 4 13 2
10 13 4 15 1 0 2 7 1 0 2
15 1 9 15 1 15 13 1 10 9 2 16 4 13 9 2
14 13 4 15 1 0 2 7 4 15 13 13 7 13 2
9 0 9 13 0 9 2 3 0 2
7 10 9 2 7 9 9 2
13 0 9 13 4 13 3 3 2 16 4 15 13 2
21 13 2 14 15 9 1 9 9 1 0 9 9 2 3 15 13 9 9 1 9 2
17 9 9 15 14 13 9 2 9 13 9 2 9 2 0 9 3 2
18 15 13 7 1 0 0 9 2 15 9 2 15 9 2 15 9 3 2
9 0 9 4 13 3 14 0 9 2
14 1 15 15 13 10 9 2 16 10 13 3 9 0 2
10 14 15 13 2 1 15 13 3 0 2
22 9 2 15 13 16 9 2 13 3 9 7 15 2 15 13 2 13 1 9 10 9 2
17 1 9 2 15 15 13 2 15 15 13 9 2 0 9 7 9 2
15 9 0 9 15 13 1 0 9 2 3 1 9 16 15 2
29 3 15 13 0 9 7 9 2 0 9 7 0 9 0 9 2 3 2 9 2 2 15 1 9 13 2 15 13 2
10 9 0 9 13 7 13 1 0 9 2
10 13 15 3 9 9 7 9 1 0 2
19 9 16 0 9 2 0 9 2 0 9 7 0 9 13 3 13 0 9 2
40 13 9 2 7 13 15 13 2 16 1 9 9 1 12 2 9 2 7 3 3 3 10 9 3 2 15 13 10 9 0 9 13 1 10 9 7 13 15 0 2
20 1 9 9 9 13 13 0 9 9 9 2 7 13 7 9 2 13 15 0 2
17 9 1 10 9 13 1 9 2 15 13 0 9 7 0 0 9 2
16 9 9 13 2 16 9 9 13 1 9 3 9 15 1 9 2
14 9 15 1 0 9 13 3 0 1 9 16 1 9 2
15 16 9 13 9 7 13 2 3 13 1 9 0 9 9 2
9 15 7 13 9 1 9 0 9 2
40 1 9 13 1 9 9 2 1 9 9 1 9 9 9 1 15 7 9 9 2 9 2 1 15 13 2 3 2 2 9 4 13 3 7 9 3 13 0 9 2
19 13 7 1 9 9 2 16 9 13 0 9 2 3 13 2 16 3 13 2
5 15 13 7 9 2
30 7 13 3 1 9 10 9 1 0 9 2 15 15 13 13 2 7 0 9 2 7 16 10 0 9 13 3 13 9 2
29 1 9 9 7 0 9 13 3 2 13 9 7 1 9 3 13 2 16 16 13 9 3 3 2 3 0 9 13 2
27 0 9 1 10 9 1 9 13 1 0 9 3 11 2 13 2 14 1 0 9 9 1 9 7 0 9 2
23 1 0 9 13 2 16 9 0 9 4 13 1 12 2 9 2 7 3 1 10 9 13 2
28 9 1 9 0 9 13 3 2 1 3 16 12 9 0 9 11 1 11 2 15 13 1 0 9 11 16 9 2
26 13 1 9 2 16 9 0 9 1 11 1 0 9 13 0 9 16 1 11 7 9 13 14 12 2 2
24 13 2 16 9 9 1 9 13 3 0 2 7 16 3 0 9 13 1 11 7 1 11 0 2
25 13 1 10 9 13 7 3 13 1 9 2 16 9 13 13 9 9 2 7 13 0 13 9 9 2
15 13 15 0 9 15 1 0 9 7 9 9 1 10 9 2
51 3 3 2 16 13 13 9 7 13 9 2 16 4 15 13 9 1 11 7 11 2 7 3 3 2 16 13 2 3 3 13 12 3 0 9 0 0 9 1 0 9 1 0 9 2 13 1 10 9 15 2
21 0 9 1 9 9 13 9 14 1 10 9 3 2 13 2 14 1 0 0 9 2
13 9 2 0 9 2 13 3 0 9 1 2 15 3
3 9 9 2
42 13 13 1 0 9 2 2 2 2 1 9 0 9 0 2 11 2 11 2 11 12 2 13 9 2 9 2 0 0 9 0 0 9 1 0 9 9 7 9 2 2 2
12 16 13 1 9 3 0 1 9 2 13 3 2
12 2 0 0 11 2 11 12 2 9 2 2 2
9 3 15 13 7 9 1 0 9 2
17 13 1 0 2 0 0 9 2 1 10 9 2 15 13 13 9 2
14 1 9 2 3 16 1 0 9 13 13 1 9 0 2
15 3 13 9 0 2 7 2 1 9 13 9 1 0 9 2
53 2 13 2 14 4 9 1 9 0 9 2 7 1 15 2 16 13 1 15 0 7 1 15 0 2 13 2 16 15 4 0 9 1 10 9 13 0 9 10 9 2 7 13 1 10 9 9 0 1 0 9 2 2
13 9 9 13 13 0 2 0 2 13 1 9 9 2
28 13 1 10 9 2 16 13 9 2 13 2 2 2 13 2 2 15 2 13 2 2 2 13 15 9 2 3 2
25 9 9 13 10 9 7 9 16 9 0 3 3 7 0 9 2 13 10 9 16 2 0 9 2 2
37 1 15 2 16 1 9 13 1 0 9 7 3 1 9 9 2 13 7 9 0 9 3 13 2 3 3 16 13 0 9 13 0 9 7 0 9 2
19 9 3 13 13 9 2 3 7 9 2 7 15 3 0 2 0 0 9 2
27 0 9 13 1 10 9 3 0 2 3 1 9 2 15 15 13 2 14 15 13 2 3 0 0 9 2 2
16 9 15 3 3 13 1 15 2 16 0 9 15 13 13 9 2
12 16 9 13 1 0 9 9 2 13 0 9 2
40 4 1 15 13 12 9 0 7 0 9 11 11 2 0 9 1 0 9 2 9 0 2 11 2 12 2 0 15 3 9 0 2 13 2 9 2 2 2 2 2
5 15 1 15 13 2
9 1 2 0 9 2 15 3 13 2
18 7 4 13 13 9 0 2 7 4 15 14 13 13 7 1 10 9 2
8 7 3 4 13 13 9 9 2
9 13 15 2 16 10 9 3 13 2
3 9 1 9
39 16 4 13 9 2 3 13 0 0 0 9 9 2 9 0 2 2 13 15 13 2 3 10 9 13 1 0 9 2 9 12 2 12 7 12 2 12 2 2
27 1 0 9 7 10 9 13 9 0 2 7 9 2 3 0 7 0 0 9 1 0 9 11 11 1 11 2
29 11 2 11 2 11 1 0 9 2 11 2 1 0 9 0 9 13 2 16 12 1 12 0 9 13 3 13 9 2
11 2 3 13 1 10 9 0 12 9 2 2
19 3 9 9 13 0 2 0 14 12 0 7 14 12 5 13 0 0 9 2
6 13 3 7 0 9 2
20 16 1 12 9 13 9 2 9 0 9 13 9 0 9 7 13 16 1 9 2
8 3 15 3 13 13 10 9 2
19 10 0 7 3 0 9 13 9 1 0 3 0 7 0 9 9 1 9 2
10 13 4 7 9 2 16 9 13 9 2
16 16 13 10 0 9 2 13 4 15 7 9 3 10 9 13 2
10 3 13 13 9 0 1 11 7 3 2
20 9 10 9 4 15 7 14 13 1 0 9 2 11 12 2 12 2 12 2 2
2 11 11
3 12 2 12
7 9 11 2 9 11 7 9
13 9 11 13 0 0 9 2 9 9 7 9 0 2
26 1 0 9 2 1 0 0 9 2 12 2 15 13 2 16 13 11 0 11 1 0 9 0 1 9 2
12 11 2 9 0 2 4 13 1 3 0 9 2
22 9 4 13 1 12 9 2 15 4 13 1 9 2 0 9 2 9 11 7 0 9 2
40 0 9 13 0 9 0 15 1 9 9 1 0 9 2 7 0 9 7 0 9 13 0 9 2 10 9 13 1 9 1 9 10 9 1 12 2 9 0 9 2
10 0 9 4 13 11 11 9 2 12 2
17 1 0 9 9 2 12 4 13 7 4 1 15 13 10 0 9 2
24 10 9 13 0 0 9 1 0 9 2 15 13 1 9 12 9 0 9 9 11 1 0 9 2
23 9 13 3 16 9 2 16 9 13 0 0 9 0 9 1 9 3 1 9 1 0 9 2
35 0 9 13 0 9 7 15 15 3 13 2 15 4 0 9 3 13 0 7 0 9 2 3 2 16 9 9 15 13 9 1 0 0 9 2
11 9 0 9 13 7 0 9 0 7 0 2
29 9 3 3 13 2 16 0 2 2 9 2 4 1 9 13 1 9 3 0 9 9 11 7 3 0 9 11 11 2
17 0 9 3 13 0 9 0 9 2 15 9 13 0 16 12 9 2
22 9 13 0 2 0 9 7 0 9 13 3 0 0 9 2 15 4 3 13 7 13 2
12 12 9 13 1 0 9 9 1 9 1 9 2
14 15 15 0 9 9 11 1 0 9 3 13 0 9 2
43 9 0 9 7 13 10 0 9 2 16 9 13 3 9 2 7 3 9 2 16 3 3 9 9 15 9 13 13 1 9 0 9 7 3 1 9 9 13 3 0 0 9 2
31 7 3 1 9 0 7 0 9 0 7 3 0 0 9 0 15 1 0 9 9 13 2 16 0 9 13 1 9 0 13 2
11 3 15 13 0 9 2 13 13 0 9 2
3 7 3 2
1 9
19 11 11 2 12 2 2 0 9 1 0 11 2 9 1 0 0 2 9 2
9 11 12 2 12 2 12 2 12 2
2 11 11
3 12 2 12
4 9 7 0 9
18 1 0 2 0 2 9 9 9 15 1 9 9 1 9 9 13 9 2
25 3 1 9 13 0 9 13 1 0 9 9 7 1 0 9 13 3 1 10 9 1 9 9 9 2
40 9 13 9 9 2 15 1 0 13 0 9 1 9 9 9 7 13 15 0 2 16 10 0 9 2 15 7 13 13 3 0 9 2 4 13 3 13 9 9 2
51 1 15 13 9 2 16 3 2 1 9 2 15 13 0 0 9 2 0 9 0 0 9 2 15 15 13 1 0 3 0 9 9 7 9 2 13 3 1 9 0 0 9 0 14 1 12 5 1 9 9 2
31 9 9 1 9 1 9 7 0 9 2 9 2 12 2 9 2 12 2 12 2 13 13 0 9 0 9 9 0 0 9 2
26 16 4 15 9 1 0 9 7 9 13 13 2 13 4 15 3 1 9 9 0 9 1 10 0 9 2
2 11 11
3 12 2 12
3 9 0 9
20 1 9 0 9 9 7 9 9 13 0 2 16 15 10 9 9 1 9 13 2
12 13 1 15 13 0 9 2 15 15 13 9 2
33 1 0 9 9 13 3 9 2 12 0 9 11 2 11 3 16 12 0 9 2 15 3 1 15 13 13 1 0 9 14 10 9 2
28 0 9 7 10 9 1 9 4 3 0 10 9 13 1 15 0 2 3 15 0 9 13 3 13 9 7 9 2
25 3 1 0 9 15 13 2 16 1 9 13 15 3 2 0 9 13 3 12 1 0 2 9 2 2
66 13 3 9 2 16 15 1 9 7 3 3 2 3 1 9 2 0 9 0 9 3 13 2 7 1 9 0 7 0 9 3 13 10 0 7 0 9 2 3 7 3 2 2 16 7 9 10 9 2 15 13 13 1 9 2 13 15 7 13 9 1 9 0 0 9 2
27 1 9 4 13 0 9 12 1 10 9 9 2 0 2 9 2 0 9 2 11 12 2 12 2 12 2 2
23 9 0 9 0 9 15 3 3 13 1 9 3 2 10 10 9 2 15 13 9 1 9 2
30 11 2 11 2 11 7 11 2 11 13 0 9 0 9 1 0 9 9 1 0 9 2 15 2 15 13 9 1 9 2
14 7 13 2 16 15 0 0 9 13 1 9 9 0 2
7 1 15 13 10 9 0 2
20 1 9 0 0 9 13 3 1 9 13 1 9 9 0 9 0 9 0 9 2
2 11 11
3 12 2 12
2 0 9
13 16 13 9 9 2 13 15 15 3 0 2 0 2
19 9 9 1 11 2 11 2 11 11 7 13 9 2 15 13 13 0 9 2
14 13 1 9 9 0 2 7 16 0 14 1 12 9 2
19 13 15 1 0 9 9 0 9 2 9 2 2 0 1 0 9 1 11 2
21 3 15 13 2 16 13 1 10 0 9 2 7 3 13 0 2 16 13 10 9 2
21 13 15 3 0 9 2 0 9 13 0 9 2 3 7 9 9 9 1 0 9 2
11 15 3 13 1 0 9 1 9 9 9 2
22 3 9 2 12 4 13 9 9 3 0 9 2 3 0 1 9 9 1 0 9 2 2
14 1 9 9 15 3 13 0 9 2 15 10 9 13 2
20 7 10 0 9 9 2 15 2 15 13 7 13 9 2 7 9 2 9 2 2
29 9 0 9 15 13 2 16 10 9 13 0 9 9 7 13 1 10 9 16 9 2 11 12 2 12 2 12 2 2
2 11 11
3 12 2 12
3 9 1 9
74 9 2 9 1 9 2 2 15 13 1 10 9 2 15 13 9 2 15 4 15 1 0 13 3 9 12 2 9 2 3 13 1 9 2 3 1 9 2 2 15 15 13 1 0 7 0 9 0 9 2 3 2 1 9 0 9 2 7 13 3 0 0 9 2 3 2 9 1 0 9 7 0 9 2
17 11 3 13 2 16 13 2 14 0 9 0 2 3 13 9 0 2
18 2 13 9 2 2 13 0 9 11 2 11 2 2 9 13 0 2 2
16 9 3 16 4 3 13 9 1 0 9 9 16 9 0 9 2
22 14 13 13 9 2 13 2 15 15 1 9 15 13 7 1 15 15 13 0 9 9 2
12 9 13 9 2 16 15 1 10 9 13 9 2
19 1 0 9 3 2 9 13 2 3 15 15 9 13 13 1 10 0 9 2
78 13 2 3 1 15 1 9 2 3 4 0 13 1 9 1 9 1 0 9 2 14 7 1 9 1 15 2 3 14 9 3 13 0 2 0 7 0 9 2 11 2 11 2 11 2 11 12 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 7 0 2
46 3 15 13 2 3 15 10 0 9 11 2 15 13 1 9 10 9 2 13 9 11 2 11 1 0 9 2 0 9 11 11 9 2 7 1 0 9 2 0 9 1 0 0 9 2 2
22 1 9 11 13 2 2 13 9 2 16 13 15 0 2 7 13 15 0 9 2 2 2
14 10 9 15 1 11 11 14 13 2 13 15 3 9 2
9 13 15 15 3 0 2 3 0 2
17 2 9 9 2 13 4 15 16 0 11 2 2 15 13 15 2 2
10 13 15 9 2 7 13 15 1 9 2
9 0 9 2 3 0 2 7 0 2
19 9 1 0 9 15 3 13 2 1 15 15 13 3 0 2 0 2 0 2
13 13 15 7 7 9 2 3 14 15 13 3 0 2
22 3 15 13 7 9 2 7 16 15 1 15 1 10 9 2 11 2 11 2 13 3 2
9 0 1 10 9 13 1 9 9 2
16 15 4 3 7 13 2 15 13 3 2 13 4 15 15 14 2
14 3 4 13 2 16 1 0 9 4 13 1 0 9 2
6 15 4 15 13 13 2
4 12 13 0 2
30 10 9 13 0 2 0 9 1 9 7 1 0 0 9 2 9 2 9 2 9 2 0 9 2 9 1 9 2 9 2
11 13 15 1 15 2 13 1 10 0 9 2
18 3 4 15 13 1 9 3 3 7 2 3 2 2 7 9 1 9 2
25 1 9 2 15 13 2 9 9 2 2 7 1 9 2 10 9 2 9 7 9 13 9 0 9 2
36 2 9 2 15 13 10 3 1 9 2 15 1 11 3 13 1 9 13 9 10 9 2 1 15 4 15 13 9 2 0 9 2 2 0 9 2
17 9 3 13 14 1 9 2 3 3 15 13 9 7 9 0 9 2
17 0 0 9 13 1 9 9 0 1 9 1 0 9 7 0 9 2
17 2 3 13 1 0 9 0 1 15 2 0 2 9 9 2 2 2
19 16 0 9 2 13 4 3 15 1 12 9 3 0 9 0 9 12 9 2
13 2 3 13 9 7 13 15 0 9 7 9 2 2
19 13 2 16 15 13 0 9 9 2 15 13 13 1 9 2 7 1 9 2
44 13 15 2 16 4 15 13 1 0 9 11 11 2 0 9 9 11 2 11 2 11 2 7 16 4 13 10 9 9 16 15 2 16 4 13 1 10 9 2 10 9 7 9 2
16 13 15 1 15 2 16 4 10 9 13 1 9 10 0 9 2
10 3 3 9 9 2 7 9 0 9 2
14 3 15 13 3 10 0 9 2 15 13 0 0 9 2
4 11 11 2 11
42 12 1 9 2 3 15 13 2 15 13 2 16 11 11 2 9 7 9 2 15 1 15 3 13 2 13 12 2 12 2 12 2 3 9 1 9 2 0 0 9 2 2
9 0 9 9 2 11 11 2 9 2
3 9 0 9
1 11
22 0 9 9 2 13 15 1 9 7 1 9 0 9 9 2 10 4 13 0 9 9 2
22 1 9 13 9 0 1 9 1 0 9 2 1 10 9 3 7 1 9 1 10 9 2
54 9 13 1 15 0 2 16 3 13 14 1 0 9 2 7 3 1 9 9 2 1 15 0 7 0 9 13 4 13 1 9 2 0 9 10 0 9 2 1 0 9 3 1 9 0 16 0 0 0 9 9 1 11 2
30 13 1 0 9 2 15 4 13 3 13 1 9 3 0 0 9 7 15 4 15 3 13 3 3 3 7 3 13 3 2
32 7 13 10 9 7 9 0 0 9 7 13 2 16 9 2 15 13 2 13 3 10 9 2 15 13 1 0 0 9 3 0 2
4 1 9 10 9
4 11 11 2 11
2 9 9
28 1 9 9 1 9 9 1 9 12 2 12 2 3 4 15 1 9 9 0 9 13 13 9 2 9 7 9 2
20 2 13 15 9 2 1 15 4 13 9 2 16 13 9 9 1 9 12 3 2
3 9 9 2
18 2 2 2 2 2 9 1 0 9 13 3 3 9 1 9 10 9 2
21 9 15 13 13 3 9 0 9 2 0 2 0 2 1 0 9 2 2 2 2 2
33 15 3 9 10 9 13 2 15 3 13 10 0 9 7 3 3 13 9 10 9 2 0 15 15 3 13 2 13 2 13 2 13 2
24 0 2 0 2 0 1 9 1 9 7 1 15 3 0 1 0 9 1 15 2 2 2 2 2
26 9 3 16 1 9 9 2 1 0 9 13 1 9 2 1 9 15 16 0 9 9 2 9 2 9 2
18 0 9 4 15 13 3 3 13 9 9 7 9 2 16 9 0 9 2
25 10 9 4 3 13 3 0 9 2 7 3 0 7 0 9 13 1 10 9 0 16 3 0 9 2
26 13 2 16 1 9 13 13 1 9 7 1 9 0 2 10 9 0 9 2 7 3 15 13 9 0 2
16 1 0 9 2 0 0 9 7 0 9 0 9 3 13 9 2
19 7 3 13 2 16 9 2 9 0 2 15 13 7 16 2 9 0 2 2
2 11 11
7 12 2 0 9 11 2 11
25 9 13 3 0 13 9 1 9 2 13 0 9 0 0 9 1 9 9 2 13 9 9 12 9 2
11 1 10 9 7 9 13 3 7 9 9 2
28 9 7 13 13 9 9 1 0 9 2 7 13 9 0 1 9 2 7 13 9 9 0 9 2 2 2 2 2
22 2 2 2 2 2 9 1 9 0 9 0 4 14 13 9 10 2 0 2 9 0 2
22 1 10 9 15 13 13 9 2 9 2 9 2 9 2 7 13 1 15 13 0 15 2
2 11 11
5 0 9 11 2 11
17 9 2 11 11 2 2 12 2 13 9 1 0 9 11 1 11 2
20 1 0 9 15 1 0 9 1 11 13 9 9 9 1 9 7 9 0 9 2
21 3 3 15 13 2 16 10 0 7 0 9 1 15 1 0 9 0 9 3 13 2
9 13 3 14 1 9 9 2 2 2
18 3 0 9 15 13 2 16 9 7 0 9 10 0 9 13 1 9 2
31 0 15 15 13 13 3 0 2 16 1 9 1 0 9 13 3 10 9 9 3 13 9 7 3 15 3 13 9 0 9 2
16 9 2 3 13 0 9 2 1 15 7 3 13 9 7 9 2
11 15 3 13 15 0 7 0 1 9 9 2
9 10 9 13 15 2 16 0 9 2
25 13 3 15 2 15 11 13 2 0 9 0 9 2 7 13 9 1 0 9 2 15 13 0 9 2
37 9 3 13 3 3 2 16 0 9 2 15 4 3 13 0 9 2 7 14 4 1 15 13 3 16 1 9 2 0 9 2 16 16 1 0 9 2
24 10 0 9 13 0 7 1 10 0 9 7 3 13 15 2 15 15 13 1 2 9 9 2 2
42 13 1 15 2 16 0 9 4 13 2 16 4 9 3 13 0 9 7 9 2 15 13 9 0 0 9 2 7 16 4 4 13 1 0 9 1 9 2 10 9 13 2
18 16 3 0 9 13 2 13 3 0 15 1 15 1 10 9 3 13 2
165 7 1 9 2 15 13 2 15 13 2 15 13 9 2 9 2 7 13 15 1 9 9 0 1 9 0 9 9 2 1 9 2 10 9 1 0 9 9 13 15 13 2 13 3 9 9 16 2 9 2 2 2 9 2 2 2 9 2 2 2 9 2 2 15 15 4 13 1 10 9 1 0 9 7 9 2 15 1 9 10 9 13 2 2 1 9 2 15 13 9 1 15 2 15 13 15 0 9 7 13 2 1 15 13 10 9 2 16 9 13 1 9 2 1 9 2 10 0 9 9 7 9 9 9 13 1 15 2 16 13 1 9 3 9 2 1 10 9 13 3 3 1 0 9 0 2 7 3 0 13 9 2 16 4 15 3 13 13 7 3 13 0 0 9 2
35 16 15 7 3 13 2 1 15 13 0 9 2 15 13 13 2 16 4 13 13 3 7 3 1 0 9 2 14 15 15 1 15 4 13 2
16 10 9 1 0 9 7 3 13 9 9 2 15 13 4 13 2
27 7 16 15 9 7 9 9 3 1 10 9 13 2 10 9 13 0 9 7 9 7 9 0 9 2 2 2
25 1 9 2 15 15 13 2 16 9 13 2 13 9 1 9 2 7 9 2 9 2 2 9 2 2
14 1 9 13 9 2 16 4 13 9 0 9 7 9 2
22 7 9 7 9 15 7 13 2 16 0 9 13 7 9 7 9 2 7 3 13 9 2
18 0 9 0 9 2 7 7 9 7 9 13 0 9 1 9 10 9 2
32 13 2 16 15 9 2 9 2 3 13 16 9 0 9 2 2 9 2 7 2 9 2 9 2 7 10 9 2 13 9 9 2
45 15 15 13 2 16 11 3 13 13 1 9 7 9 9 2 16 13 10 0 9 2 16 15 2 16 3 15 13 3 2 15 13 9 13 2 13 7 9 1 9 7 9 1 9 2
23 7 3 16 3 9 7 9 0 9 9 13 3 9 1 15 2 3 3 9 2 13 2 2
9 11 11 2 11 2 9 1 0 9
14 0 2 9 2 0 2 9 12 2 12 2 12 2 12
21 13 3 3 9 2 3 4 3 13 13 10 9 15 2 15 4 13 13 2 2 2
36 0 0 7 0 9 0 9 13 13 9 1 10 0 0 9 2 2 2 16 4 13 1 9 9 0 13 2 13 7 13 10 9 3 2 2 2
25 1 9 1 9 9 1 9 9 7 9 13 1 0 9 3 1 9 1 9 9 1 9 7 9 2
28 10 9 13 1 10 9 2 9 2 9 1 9 0 9 1 0 7 0 9 7 13 1 9 0 9 10 9 2
16 13 3 2 16 3 15 13 9 2 0 2 7 2 0 2 2
10 13 15 15 2 16 15 13 0 9 2
21 0 9 0 9 4 3 13 0 13 2 13 15 7 2 16 4 15 0 9 13 2
13 7 0 0 9 3 13 2 13 15 2 2 2 2
17 0 7 0 9 9 0 0 9 13 9 2 15 15 13 9 9 2
20 16 1 15 4 1 9 0 9 9 13 0 9 9 7 9 2 10 9 13 2
32 10 9 13 14 3 2 16 9 13 7 13 2 16 9 13 3 0 9 1 9 7 16 13 1 3 0 9 16 10 0 9 2
24 14 3 13 0 2 16 15 1 15 3 7 3 13 9 2 15 13 9 3 13 1 10 9 2
9 11 11 2 11 2 9 1 0 9
14 0 2 9 2 0 2 9 12 2 12 2 12 2 12
14 11 11 2 11 13 9 1 0 0 9 1 0 11 2
15 11 11 2 11 13 9 9 1 9 0 9 0 0 9 2
16 9 1 15 15 13 10 9 2 7 3 0 10 9 13 9 2
24 0 9 7 9 7 13 3 3 13 7 1 9 9 2 2 2 7 7 1 9 0 2 2 2
26 9 13 13 3 9 2 15 13 9 1 10 9 2 3 9 9 2 15 13 3 0 2 7 0 9 2
16 13 13 0 9 2 15 15 13 13 9 1 0 9 2 2 2
29 3 4 0 13 1 10 0 9 7 0 0 9 2 15 3 13 13 14 0 9 2 7 3 10 9 13 13 9 2
13 9 13 0 9 3 1 0 2 3 7 0 9 2
34 7 9 9 2 13 2 14 1 10 9 1 9 2 13 2 16 13 1 9 10 9 13 3 7 3 2 16 13 3 1 10 9 0 2
31 7 9 9 2 0 0 9 2 13 9 2 15 0 13 15 2 2 4 13 3 3 2 16 1 10 9 9 3 3 13 2
17 11 11 7 11 11 2 9 0 9 7 9 2 11 2 11 2 12
2 9 11
29 9 0 10 9 3 1 9 0 15 1 9 13 3 14 1 9 1 2 0 2 9 13 10 0 9 1 9 0 2
18 7 9 15 13 1 10 9 7 10 9 1 15 1 15 13 10 9 2
11 9 0 9 7 9 13 1 9 3 0 2
15 16 15 13 9 2 13 15 7 3 1 9 2 3 9 2
44 3 1 9 2 12 13 1 11 3 3 0 9 0 15 16 2 0 11 11 2 2 1 3 1 9 0 9 9 0 2 0 1 11 2 2 15 15 13 1 9 13 15 0 2
33 7 14 9 2 7 15 9 3 2 3 7 9 2 9 2 9 2 9 3 2 2 7 3 7 9 2 9 2 0 9 7 9 2
7 3 0 1 0 10 9 2
10 3 9 2 12 13 14 10 9 9 2
26 3 15 10 9 13 3 1 9 2 13 0 9 7 13 1 0 9 2 11 12 2 12 2 12 2 2
19 9 0 0 9 9 13 0 0 0 9 11 2 11 2 11 1 0 9 2
21 16 0 9 15 9 13 9 10 9 16 9 2 7 15 3 9 0 9 7 9 2
17 13 15 15 3 2 11 2 15 9 13 1 10 2 9 0 2 2
18 9 9 1 9 7 15 13 2 7 3 10 9 13 13 14 1 9 2
18 1 15 3 1 9 9 9 2 13 3 9 12 2 12 2 12 2 2
22 15 7 1 0 9 13 9 0 2 7 3 0 9 2 13 9 1 9 2 12 2 2
2 11 11
3 12 2 12
4 3 3 7 3
37 3 3 7 3 13 9 1 0 9 14 12 9 0 9 0 9 2 9 0 2 2 15 13 1 15 13 16 0 9 3 0 1 9 1 9 3 2
10 0 9 13 0 1 10 9 10 9 2
50 10 0 9 2 15 15 13 1 10 3 0 9 9 2 13 3 1 9 0 9 2 9 0 9 2 2 0 0 9 2 2 1 15 9 13 11 2 11 2 11 0 9 2 16 15 13 0 9 9 2
25 0 9 2 0 7 0 0 9 3 3 13 2 7 3 13 1 0 9 2 0 1 15 0 2 2
18 3 0 9 13 1 0 9 9 13 3 1 0 0 9 16 1 0 2
6 3 15 0 9 13 2
28 15 13 9 3 0 0 0 7 0 9 2 7 3 13 9 2 15 13 1 9 1 0 9 2 9 3 0 2
22 1 10 0 9 15 3 13 3 2 9 0 9 2 16 4 15 13 3 1 9 9 2
11 3 15 1 10 9 13 9 1 0 9 2
17 9 13 12 10 9 2 11 2 11 2 12 2 12 2 12 2 2
15 12 1 15 13 0 0 9 7 0 0 2 3 0 9 2
13 0 13 13 14 0 9 2 16 13 0 3 13 2
24 1 9 2 15 13 13 12 9 2 4 13 0 9 9 0 7 0 9 1 12 9 1 0 2
20 0 9 2 1 0 3 0 9 2 13 15 0 3 2 2 9 10 9 13 2
19 0 0 9 3 13 13 0 9 1 9 7 3 7 0 2 3 0 9 2
2 11 11
3 12 2 12
2 0 9
5 9 0 9 1 9
20 12 1 0 9 0 9 2 15 13 2 13 9 12 2 12 2 12 2 12 2
10 1 10 9 15 13 0 9 0 9 2
16 0 9 2 13 3 0 0 9 16 9 0 7 15 9 3 2
22 13 2 14 0 9 9 1 0 9 1 10 9 2 13 0 0 9 16 9 0 9 2
43 0 9 13 0 9 10 0 9 2 16 13 15 1 0 9 9 13 3 3 15 13 1 9 0 9 2 9 7 1 9 2 3 3 1 10 0 7 3 0 9 0 9 2
25 0 9 7 9 15 3 13 9 0 9 2 15 13 0 9 2 1 10 9 13 3 1 9 9 2
39 9 0 2 10 0 9 1 9 9 13 2 12 2 0 9 0 9 1 0 9 12 2 15 4 13 1 9 1 9 9 2 9 9 7 9 7 0 9 2
11 12 2 9 9 7 9 2 9 0 9 2
6 12 2 9 0 9 2
9 12 2 0 9 9 12 1 9 2
5 12 2 0 9 2
8 9 0 13 0 0 9 9 2
20 1 9 0 10 9 13 2 1 0 9 10 9 13 2 13 9 2 12 2 2
18 10 9 4 13 3 2 7 2 16 0 9 9 12 13 9 0 9 2
39 13 7 0 2 16 9 13 3 0 2 9 9 9 13 0 9 9 12 2 15 3 13 9 0 9 2 1 15 13 1 9 0 9 7 0 9 9 12 2
30 9 9 7 9 0 9 13 1 9 2 12 1 0 9 9 9 12 1 9 2 1 9 2 12 1 0 0 9 9 2
5 3 13 10 9 2
12 9 9 12 13 1 0 9 7 0 13 9 2
14 9 9 12 15 1 9 13 3 1 12 2 12 9 2
26 9 2 10 0 9 13 0 9 2 0 9 2 0 9 1 9 9 2 9 9 2 9 9 7 9 2
17 9 2 12 13 9 12 2 12 9 9 2 3 13 14 12 9 2
25 9 9 2 13 15 3 1 9 9 12 9 2 13 7 1 9 2 7 1 9 2 15 13 9 2
15 0 9 9 12 9 13 3 12 9 2 0 1 12 9 2
19 9 2 7 0 2 0 9 13 0 9 9 2 15 13 3 1 0 9 2
14 1 9 15 13 3 3 1 9 9 7 0 9 9 2
7 13 0 9 1 0 9 2
6 13 0 7 3 0 2
23 9 9 12 2 13 13 1 9 0 9 0 0 9 7 10 9 1 9 1 9 9 12 2
24 0 9 15 13 2 10 9 0 4 13 3 2 16 4 13 0 0 9 16 15 10 9 3 2
13 3 2 9 13 12 7 3 0 9 16 9 12 2
15 9 9 13 3 12 7 7 12 7 3 9 16 9 12 2
15 9 0 9 13 1 9 9 12 2 3 1 9 0 9 2
9 0 7 0 9 9 1 0 12 9
31 1 9 0 9 13 9 9 9 12 12 9 2 9 2 12 3 12 9 7 9 12 9 4 3 13 1 9 12 2 12 2
13 1 0 12 9 4 13 12 5 9 9 9 12 2
11 0 9 9 1 0 9 3 13 1 15 2
19 3 4 1 0 12 9 13 9 0 9 2 16 4 13 13 9 1 9 2
21 2 3 15 13 13 0 2 16 10 9 1 0 9 9 13 0 2 14 0 9 2
30 3 2 14 3 13 10 9 16 0 7 0 9 2 16 13 0 11 7 11 7 3 16 13 0 7 0 9 12 9 2
8 0 9 15 13 9 10 9 2
19 2 1 0 9 4 13 1 0 9 13 1 9 9 3 1 12 2 9 2
10 0 9 13 0 2 3 14 3 0 2
9 9 9 15 13 1 9 2 12 2
16 1 9 12 2 12 13 0 9 0 2 3 3 13 1 9 2
24 9 0 9 1 0 9 13 1 9 2 7 0 9 13 0 7 13 2 16 13 1 0 9 2
15 2 0 9 15 13 3 16 0 2 3 1 0 12 9 2
18 0 9 13 1 9 7 9 9 0 1 0 9 7 0 1 9 0 2
11 9 13 0 9 1 9 7 0 1 9 2
11 9 4 15 13 13 2 7 9 13 9 2
7 0 9 1 9 13 0 2
14 9 7 0 9 13 1 9 0 9 7 9 0 9 2
10 2 0 9 13 1 9 7 0 9 2
20 1 0 9 13 1 9 9 1 12 2 12 5 7 3 1 3 0 9 9 2
13 1 9 9 1 9 2 12 13 3 1 0 9 2
16 0 9 13 1 9 2 12 3 0 9 9 2 3 1 9 2
16 1 9 2 12 15 13 0 7 0 9 9 7 1 0 9 2
24 16 0 9 1 0 9 13 0 1 0 9 2 13 1 0 9 1 0 2 0 9 0 9 2
18 0 0 9 2 3 11 2 13 3 9 2 0 9 13 3 1 9 2
43 2 1 9 9 9 9 9 12 7 0 9 9 15 9 2 11 13 2 16 9 2 12 2 3 13 1 9 9 9 12 1 9 1 9 1 0 9 2 13 10 0 9 2
11 2 9 13 1 12 2 9 7 1 15 3
11 2 9 13 14 1 12 5 7 3 7 9
5 2 13 15 9 9
7 2 9 9 15 13 14 3
17 3 15 3 13 1 9 2 7 1 15 10 9 13 0 9 9 2
23 12 1 15 0 13 0 9 9 2 0 1 9 7 9 9 2 15 3 13 1 0 9 2
8 0 0 9 13 9 0 9 2
8 9 9 1 11 1 0 12 9
9 0 9 13 14 12 5 9 9 2
9 13 3 1 9 0 9 0 9 2
8 3 13 12 1 0 0 9 2
20 0 9 11 13 1 0 0 9 16 11 2 16 0 9 13 3 0 0 9 2
10 1 0 12 9 4 13 10 0 9 2
9 12 2 9 13 10 3 0 9 2
12 13 3 7 1 9 13 2 16 11 15 13 2
19 1 0 9 13 1 9 12 2 9 1 9 12 2 12 13 3 1 9 2
8 13 15 9 0 7 0 9 2
11 0 9 15 13 2 0 9 15 3 13 2
10 3 13 0 9 3 0 16 0 9 2
2 12 2
17 3 16 1 9 9 13 1 0 9 9 2 1 9 1 12 5 2
17 9 4 13 3 1 9 7 9 2 9 7 9 3 13 0 9 2
2 12 2
29 9 9 13 9 7 0 9 2 3 13 3 0 9 0 1 9 1 9 0 9 2 15 15 13 3 1 9 11 2
8 1 11 3 13 10 0 9 2
10 9 9 13 9 2 7 13 3 0 2
8 13 15 13 0 9 0 9 2
5 9 2 7 9 2
8 0 9 1 9 7 9 0 9
2 11 11
49 0 9 2 15 15 1 10 9 1 9 11 2 11 2 11 3 13 1 10 9 13 0 9 3 0 9 9 1 0 10 9 12 9 2 13 3 0 9 1 10 0 9 2 7 3 10 0 9 2
35 0 1 15 13 9 11 11 2 11 2 12 2 2 2 0 0 9 2 0 9 1 0 9 2 2 15 13 1 0 11 11 1 0 11 2
23 9 2 11 1 0 12 9 9 13 9 3 3 12 0 9 0 15 0 9 7 9 9 2
28 1 0 9 2 1 15 15 13 9 10 0 9 2 3 1 9 0 11 0 0 9 2 4 13 9 0 9 2
13 1 0 9 7 3 1 9 9 0 13 10 9 2
2 0 9
27 0 9 13 9 2 15 9 0 9 7 10 0 9 1 9 13 3 1 9 9 0 9 7 15 15 13 2
25 9 2 0 9 2 15 3 3 13 1 9 0 9 9 0 0 9 0 1 9 0 2 0 9 2
29 13 15 0 2 7 3 0 9 2 9 9 1 9 4 13 9 7 9 0 9 2 7 9 9 0 9 0 9 2
24 14 1 9 12 2 9 13 9 3 0 9 9 1 9 2 0 15 3 1 0 9 0 9 2
28 9 12 2 9 13 11 2 11 2 11 9 0 0 9 2 15 13 1 9 1 0 9 9 7 9 9 0 2
12 9 4 13 0 9 2 10 9 13 9 3 2
16 3 13 1 11 10 0 9 2 15 13 9 1 0 0 9 2
18 0 9 13 2 16 13 13 12 1 10 0 9 1 0 9 2 9 2
6 9 13 0 9 0 2
10 9 7 9 13 0 9 1 9 9 2
14 7 3 1 10 9 15 13 2 0 9 2 0 9 2
26 10 9 7 13 0 7 3 13 9 1 0 9 2 13 0 9 2 13 0 9 7 13 0 0 9 2
16 9 12 2 9 15 0 9 3 13 7 9 0 13 13 0 2
18 1 10 9 15 1 0 9 13 13 0 3 3 0 9 1 0 9 2
8 3 3 13 1 9 0 9 2
10 2 9 2 13 14 1 9 9 12 2
32 9 12 2 9 2 3 0 9 7 9 0 9 2 13 11 11 2 9 0 9 1 9 9 1 11 2 0 9 1 9 9 2
13 1 0 9 0 15 0 9 13 15 10 0 9 2
7 0 9 15 13 1 9 2
12 12 2 9 10 9 13 3 13 0 0 9 2
21 9 13 9 9 3 1 9 1 9 9 2 9 9 2 9 9 7 0 0 9 2
35 9 13 3 13 2 3 13 2 16 10 9 2 3 2 11 2 11 2 11 12 2 13 2 16 0 9 0 9 13 9 0 16 0 9 2
6 13 15 2 9 2 2
21 3 12 2 9 12 13 0 9 1 0 9 3 0 1 0 9 2 1 12 9 2
19 9 11 13 9 12 9 2 9 1 0 9 1 11 7 13 15 1 9 2
7 10 9 13 3 1 11 2
20 9 1 9 0 9 13 9 1 9 0 9 3 1 15 2 16 13 0 9 2
16 15 2 15 15 3 13 2 13 3 9 0 9 2 16 9 2
2 9 12
9 9 9 2 0 9 0 9 10 9
35 3 13 9 2 16 15 1 10 9 13 9 7 9 2 16 1 0 9 0 2 0 7 0 9 10 9 15 3 13 0 7 0 0 9 2
18 9 2 11 13 2 3 15 9 13 1 9 1 0 9 1 12 9 2
42 1 12 9 9 13 9 9 2 9 2 9 2 9 2 0 7 0 9 2 15 13 9 0 9 7 9 9 7 13 3 0 9 16 1 10 9 2 3 13 9 0 2
19 1 0 9 13 10 9 2 10 9 7 9 7 3 10 0 7 0 9 2
17 10 9 13 2 16 9 9 0 0 9 13 0 2 7 3 0 2
20 13 2 16 13 1 9 9 15 2 16 3 13 0 9 2 7 0 15 13 2
14 13 9 0 9 7 0 9 9 12 1 9 0 9 2
18 13 15 7 2 16 9 9 13 3 16 9 0 9 0 16 9 11 2
44 3 3 7 3 3 15 13 9 9 2 11 2 11 2 16 2 9 1 0 9 3 13 10 0 0 0 9 2 3 2 9 1 0 9 7 0 9 7 1 9 7 9 2 2
28 2 13 15 2 15 4 15 13 2 16 4 0 9 13 9 1 9 0 9 3 2 2 13 15 11 2 11 2
20 13 4 1 2 9 2 11 2 1 10 9 2 1 9 10 0 7 0 9 2
17 13 4 4 13 9 1 9 9 7 9 2 1 15 15 13 9 2
40 13 0 2 15 4 13 1 9 2 15 13 0 1 0 9 9 2 7 3 4 13 9 1 0 9 2 16 4 13 0 9 13 15 1 0 9 10 0 9 2
17 7 15 15 4 15 13 1 9 0 9 1 9 3 0 0 9 2
9 0 9 1 0 9 2 9 9 9
15 1 10 0 9 13 3 0 13 15 9 7 9 0 9 2
4 3 13 0 2
15 13 9 9 7 9 1 9 1 12 2 9 13 3 0 2
18 9 13 13 3 2 3 1 0 9 15 13 0 9 9 1 0 9 2
27 0 9 15 3 13 14 3 3 2 7 3 2 16 9 13 1 9 2 7 3 2 16 15 1 15 13 2
13 0 9 0 9 7 13 13 0 16 9 0 9 2
24 10 0 9 13 13 1 9 0 9 2 16 9 0 9 13 13 16 9 9 2 3 9 9 2
18 9 3 3 13 0 9 2 15 13 0 1 15 0 9 1 0 9 2
7 3 3 15 13 9 9 2
13 3 13 15 3 9 9 0 1 0 9 0 9 2
12 3 15 13 9 9 0 1 0 7 0 9 2
9 11 13 0 9 2 16 11 0 2
20 13 3 1 0 9 9 13 0 9 2 7 13 2 1 10 9 4 9 13 2
5 0 9 13 9 2
22 9 0 9 13 0 9 2 7 10 9 1 9 9 7 10 9 9 13 3 0 9 2
5 9 12 2 9 12
10 0 0 9 2 3 13 2 3 13 2
19 11 2 11 2 11 2 12 2 13 1 11 9 0 9 0 15 0 9 2
38 0 12 5 9 2 1 15 15 13 0 9 7 0 13 0 0 9 2 2 1 0 9 2 13 1 0 12 2 12 9 0 9 2 15 13 0 9 2
17 1 9 15 13 2 16 3 0 9 11 13 1 9 12 2 12 2
10 1 9 12 7 13 1 3 0 9 2
23 7 15 12 5 3 3 0 7 0 9 4 3 1 0 9 13 10 9 1 9 1 9 2
30 0 9 13 7 1 0 9 7 3 0 9 13 10 0 9 2 1 15 13 9 2 15 13 9 7 4 13 9 9 2
32 0 9 1 0 9 7 13 3 0 2 7 16 15 15 13 2 9 13 7 13 13 0 9 9 2 7 16 4 3 13 9 2
42 13 2 14 15 0 12 9 9 0 9 7 9 9 2 16 4 15 13 1 9 9 2 13 15 9 12 9 9 9 12 2 15 3 13 9 0 9 1 12 2 9 2
7 10 9 3 13 3 0 2
25 3 15 13 3 3 2 1 9 12 2 12 13 1 0 9 0 9 0 9 16 1 0 12 9 2
13 13 15 7 2 16 0 9 13 0 9 0 9 2
18 3 15 13 9 0 0 9 2 15 15 1 0 9 3 3 3 13 2
23 7 13 13 9 0 9 2 1 15 3 15 13 2 3 16 4 1 10 9 13 0 9 2
67 7 1 15 9 1 9 9 2 1 9 10 9 7 9 10 9 2 15 3 13 2 16 10 3 0 9 13 3 14 0 2 16 9 9 0 15 1 9 0 0 9 7 3 3 0 16 0 9 9 9 7 9 15 9 0 9 2 16 13 0 9 3 13 10 0 9 2
29 9 9 13 1 15 2 16 13 11 2 11 2 11 2 16 4 9 13 7 15 15 1 15 13 16 9 1 9 2
3 0 9 2
46 0 9 2 3 0 1 0 9 13 9 14 12 0 9 7 12 9 9 2 0 9 2 2 0 11 0 11 2 12 2 0 11 11 2 2 15 13 3 0 9 10 9 1 9 9 2
40 10 9 13 1 12 0 9 2 9 16 0 9 2 9 12 2 12 2 12 2 12 2 7 9 7 9 0 1 9 2 9 12 2 12 2 12 2 12 2 2
3 9 1 9
3 11 11 2
3 9 9 2
8 0 9 1 0 9 0 9 2
4 11 7 9 2
3 11 12 2
39 0 0 9 2 15 15 13 9 0 9 2 13 10 0 9 1 9 0 7 13 15 9 9 0 2 15 1 12 2 9 2 1 2 10 2 9 2 13 2
6 0 9 13 10 9 2
25 13 1 9 1 0 9 2 1 9 0 9 2 0 9 2 9 9 2 1 9 7 9 0 9 2
40 15 10 0 7 0 9 1 15 3 3 13 2 13 15 3 0 1 0 7 13 3 0 9 9 2 15 1 12 2 9 2 10 2 9 2 13 1 0 9 2
9 0 9 10 9 3 13 0 9 2
26 9 0 9 13 1 9 0 7 9 0 9 1 0 9 0 9 2 9 0 0 9 7 9 11 0 2
11 13 15 9 0 9 1 0 0 9 9 2
20 9 13 0 7 0 9 0 9 0 0 9 1 0 0 9 2 9 7 9 2
30 13 15 1 9 0 1 9 9 2 15 13 1 0 9 2 1 9 0 9 7 9 2 7 1 9 0 9 0 9 2
4 11 11 2 11
7 13 0 9 1 0 9 2
2 11 0
16 0 9 2 9 0 9 7 9 2 13 0 3 0 0 9 2
13 10 9 15 1 0 0 9 13 1 12 9 3 2
29 0 9 10 9 1 0 9 2 14 7 3 1 15 2 4 3 13 9 1 0 9 10 9 7 9 0 0 9 2
11 0 9 1 9 0 9 15 13 3 9 2
16 0 9 4 13 12 9 2 9 0 9 7 9 9 0 9 2
44 3 3 15 13 9 1 9 1 9 1 0 9 0 9 1 9 1 0 2 0 2 15 7 13 7 15 2 9 9 2 9 15 10 0 9 4 13 7 0 9 9 0 9 2
56 9 9 0 9 4 13 3 3 0 9 2 0 9 9 2 7 2 3 16 12 5 0 0 9 2 4 13 7 0 9 0 9 2 7 9 9 0 9 1 9 9 3 0 9 0 10 0 9 13 10 0 0 9 1 0 2
15 10 9 0 9 15 3 13 1 0 2 0 9 0 9 2
26 3 15 7 13 9 2 16 9 9 13 1 10 0 9 2 0 3 3 16 9 9 2 9 7 9 2
41 0 9 2 3 2 1 15 0 9 15 3 13 1 0 9 13 3 3 2 13 2 14 1 9 2 1 15 3 13 0 9 9 2 0 9 0 2 0 0 9 2
34 13 15 2 16 1 0 9 13 0 3 0 9 1 0 2 0 9 2 15 9 1 0 9 0 9 7 9 9 13 0 9 0 9 2
26 1 9 9 0 9 15 7 3 13 13 9 2 10 9 15 13 13 16 0 2 0 9 0 9 9 2
25 9 9 13 13 0 9 9 1 0 0 9 7 13 0 2 16 9 1 15 13 16 9 0 9 2
44 1 9 1 3 0 9 7 0 9 13 0 9 2 7 0 9 9 0 1 0 9 2 7 3 9 1 0 9 2 9 0 1 9 0 9 7 9 0 3 1 9 0 9 2
25 1 0 9 15 3 3 13 3 1 9 9 3 0 9 2 1 10 9 13 1 9 0 9 9 2
45 0 9 1 10 9 13 9 0 9 2 9 2 11 7 0 2 0 9 2 12 2 15 13 1 9 0 9 1 9 9 7 1 0 9 12 1 3 0 0 9 2 0 0 9 2
42 9 2 0 0 9 2 7 2 1 0 0 9 9 9 2 13 3 3 0 2 16 4 13 9 0 2 9 2 9 7 0 0 0 9 2 15 13 0 9 0 9 2
12 1 10 9 1 0 9 4 9 0 9 13 2
22 13 3 0 2 16 1 9 0 9 13 13 0 10 0 9 2 0 1 9 9 9 2
25 0 9 3 13 2 16 15 10 9 13 14 1 3 0 9 2 7 7 1 9 0 0 9 9 2
18 1 9 9 0 9 15 13 13 0 9 9 1 10 9 7 0 9 2
10 13 15 3 13 0 9 1 10 9 2
21 3 3 4 13 2 16 10 9 13 1 9 9 7 0 0 9 9 0 0 9 2
16 0 13 1 15 14 0 9 9 2 7 1 0 9 9 9 2
8 9 4 3 13 9 0 9 2
13 9 9 0 0 9 13 1 15 0 7 3 0 2
30 9 0 9 15 3 13 1 9 0 1 0 9 2 1 9 9 1 12 1 12 12 9 15 13 9 3 1 9 2 2
22 9 0 9 13 3 3 0 2 3 7 7 3 1 10 9 9 0 9 1 9 13 2
66 1 0 9 10 9 13 0 9 7 0 9 0 9 2 3 0 9 13 1 9 2 1 0 9 3 13 9 2 9 2 9 7 3 0 9 2 3 0 9 10 9 4 13 2 2 7 9 0 9 2 3 1 0 9 2 9 2 9 2 9 2 9 2 9 2 2
46 0 13 2 16 0 9 13 13 14 1 0 9 2 3 2 1 10 0 9 2 7 7 1 9 0 1 9 2 15 13 0 9 9 0 9 9 2 3 9 7 13 7 9 9 9 2
32 1 9 0 9 13 0 13 15 14 3 0 0 9 1 0 9 2 0 2 9 2 9 2 9 2 9 2 9 7 9 2 2
15 3 4 3 13 12 9 2 13 15 7 9 14 12 9 2
40 0 9 2 3 3 0 9 2 13 3 1 0 0 9 2 7 16 4 9 0 9 13 4 13 16 0 9 0 9 2 13 4 10 9 3 12 1 0 9 2
40 7 0 9 9 1 15 2 0 9 9 0 12 9 9 2 13 3 3 0 16 9 0 9 10 0 9 2 16 3 2 9 9 12 7 0 2 9 2 9 2
31 0 0 9 2 15 13 9 13 1 9 9 3 0 0 9 2 13 1 9 9 12 0 2 3 9 0 0 0 9 3 2
28 10 9 7 1 10 9 13 13 9 10 9 2 3 3 2 16 0 9 0 9 1 9 9 9 13 3 0 2
29 1 9 1 9 2 15 4 4 13 1 0 0 9 1 9 0 9 7 0 9 2 15 1 9 13 13 3 3 2
40 7 16 10 0 0 9 13 0 13 9 0 9 2 0 9 9 2 0 9 2 0 2 7 0 9 2 0 0 9 13 0 7 13 0 0 9 1 0 9 2
27 9 9 9 1 0 9 13 3 2 16 15 14 3 0 9 13 0 13 0 9 1 9 7 9 12 9 2
29 4 13 3 9 1 9 0 9 2 9 0 2 9 2 9 2 9 2 2 7 7 9 9 2 9 7 0 9 2
12 1 10 0 9 13 3 13 7 9 0 9 2
10 13 15 7 0 9 0 7 0 9 2
10 0 0 9 13 3 3 0 0 9 2
38 1 9 9 1 0 9 13 3 9 3 0 9 2 16 15 13 13 9 1 0 9 2 7 13 0 2 16 13 9 0 9 10 9 1 9 1 0 2
15 1 0 9 0 0 9 1 0 9 13 3 14 10 9 2
17 13 15 2 16 0 9 13 13 13 9 1 9 10 9 9 3 2
45 1 15 2 16 0 9 13 1 3 0 9 0 1 0 9 2 13 7 9 2 16 1 10 9 1 9 13 0 13 12 2 12 9 9 2 16 4 4 13 9 0 1 10 9 2
21 9 10 9 1 9 7 13 0 2 7 1 0 9 13 7 0 0 9 7 9 2
27 16 3 0 9 3 0 9 0 9 1 9 13 0 2 1 15 0 13 9 10 9 1 0 9 0 9 2
37 3 3 9 0 2 9 9 2 7 2 0 0 9 0 9 7 9 10 9 1 9 2 4 13 13 0 9 7 13 10 9 7 0 9 1 9 2
34 1 15 3 0 9 13 3 0 2 16 0 0 9 13 9 1 0 0 9 2 15 13 0 13 1 9 1 9 9 9 1 0 9 2
16 0 13 3 9 9 2 15 15 10 9 13 0 9 1 9 2
23 1 9 9 0 9 7 9 10 9 13 0 9 2 16 15 0 9 13 1 0 2 9 2
46 13 15 3 2 16 10 9 15 13 13 14 1 10 0 9 1 9 2 1 15 15 13 9 0 9 2 3 0 0 9 0 1 9 9 12 2 3 2 1 10 9 9 12 9 12 2
26 10 9 2 0 3 1 0 9 2 7 0 7 1 0 9 7 9 2 15 3 13 1 9 0 9 2
39 10 0 9 13 0 13 9 9 9 0 1 9 1 9 2 9 2 0 9 0 2 2 2 15 1 9 1 0 7 0 9 13 1 9 9 10 0 9 2
33 13 3 1 9 2 16 1 9 13 13 7 9 0 0 9 2 15 3 2 3 1 0 9 2 13 13 10 0 9 1 0 9 2
38 0 9 9 9 12 13 7 9 14 1 9 2 7 7 1 9 0 9 7 15 2 16 13 9 0 7 0 2 13 1 9 0 2 3 3 0 9 2
16 0 0 9 13 3 1 9 9 0 9 7 3 0 0 9 2
14 13 15 2 16 0 0 9 13 3 0 0 0 9 2
18 0 9 1 9 7 0 9 9 13 3 0 9 1 9 0 0 9 2
29 13 3 1 9 0 0 9 2 3 2 3 0 0 9 9 7 9 9 1 9 2 2 16 3 1 9 9 13 2
25 1 9 9 13 0 13 2 16 1 0 0 9 9 15 1 9 0 9 13 7 0 9 0 9 2
25 0 9 0 9 13 3 2 9 2 9 2 1 12 2 0 2 9 2 15 13 0 0 0 9 2
13 10 9 4 3 13 1 9 9 0 3 0 9 2
21 1 0 3 0 9 13 3 13 0 9 10 9 1 9 0 9 7 0 0 9 2
34 13 3 2 16 1 0 9 0 9 1 9 13 14 10 9 1 9 2 7 3 10 9 1 9 2 15 3 13 7 1 0 9 9 2
34 1 10 9 13 7 0 9 2 10 9 13 3 1 9 7 9 0 9 1 9 2 1 9 0 9 1 9 7 1 9 3 0 9 2
28 13 0 2 16 1 0 0 9 13 0 9 10 9 1 9 3 13 2 13 7 0 13 10 9 0 0 9 2
26 13 7 3 13 0 2 9 2 15 13 9 10 9 0 7 0 9 0 9 13 7 7 13 0 9 2
16 0 9 4 3 3 13 2 3 3 2 9 1 3 0 9 2
11 3 0 7 0 9 13 0 13 10 9 2
30 1 10 0 9 15 13 9 9 1 9 2 9 0 2 9 2 1 0 9 2 9 2 0 9 2 14 1 0 9 2
20 10 9 13 13 9 0 9 1 9 9 0 9 2 7 15 13 10 0 9 2
24 0 9 15 13 7 1 9 0 9 2 1 15 13 1 9 0 9 1 9 1 0 0 9 2
12 13 15 3 1 0 0 9 10 0 0 9 2
20 15 10 9 13 3 0 7 13 10 9 1 0 9 1 0 9 1 9 9 2
11 13 7 9 0 9 3 0 9 1 9 2
19 13 1 10 9 13 3 0 2 13 2 14 9 9 9 1 9 3 0 2
19 1 9 9 1 9 15 13 1 0 0 9 9 2 10 9 7 9 9 2
38 1 12 9 3 13 0 0 7 0 9 10 9 7 0 2 1 9 0 9 2 1 0 9 3 10 3 0 9 1 9 7 0 9 0 9 0 9 2
20 0 9 9 13 13 0 9 1 0 9 9 7 1 10 9 1 9 0 9 2
19 3 3 13 10 9 3 12 1 10 9 0 1 9 9 7 9 0 9 2
56 1 9 0 9 13 7 0 0 9 10 9 13 7 13 10 9 13 15 3 0 9 7 0 9 2 9 0 9 2 9 0 9 2 0 9 2 1 9 0 0 9 1 9 2 7 16 9 10 9 4 0 13 14 1 9 2
1 9
1 9
1 9
2 0 9
2 0 9
5 0 9 9 9 12
14 9 13 1 9 10 9 2 16 4 15 15 13 0 2
24 7 3 0 9 7 9 2 15 1 9 13 0 9 2 13 1 12 12 3 9 9 0 9 2
14 14 13 15 2 16 9 13 10 9 7 0 9 13 2
16 9 9 13 3 0 2 13 9 2 16 9 9 13 9 0 2
7 9 13 3 1 9 9 2
19 9 7 9 13 3 3 9 2 16 13 1 9 7 13 15 3 13 9 2
25 3 13 2 3 1 9 9 3 13 15 9 1 0 9 2 7 9 0 3 13 1 9 0 9 2
12 9 15 3 9 13 7 3 15 1 9 13 2
6 9 2 9 2 11 2
6 11 2 9 2 11 12
16 1 9 12 13 1 9 11 9 11 11 2 9 1 9 2 2
21 1 12 9 3 3 13 10 2 0 9 1 9 2 2 9 9 9 7 9 2 2
29 12 9 13 3 0 3 15 2 15 13 1 0 9 3 3 0 0 0 9 1 0 2 0 9 9 0 1 11 2
15 0 13 1 9 1 10 9 7 9 1 0 9 0 9 2
26 3 13 1 9 13 1 9 0 2 3 0 9 0 9 2 15 15 13 9 0 9 1 9 0 9 2
13 13 15 9 1 0 9 3 0 7 1 9 0 2
3 2 11 2
23 3 2 15 15 13 2 16 9 2 9 2 9 7 9 4 13 9 2 9 7 10 9 2
18 13 3 9 1 9 2 3 9 7 9 1 9 2 3 9 1 9 2
15 3 13 1 15 9 15 2 7 16 4 13 0 1 15 2
21 1 15 2 0 0 0 13 13 9 1 9 7 13 2 16 4 13 2 3 13 2
14 9 3 1 10 9 13 13 7 3 3 16 3 3 2
10 13 9 15 15 2 13 9 15 15 2
10 10 2 9 15 2 13 9 10 9 2
7 11 9 2 9 2 9 2
5 12 2 9 2 12
20 2 1 15 2 16 4 1 15 13 2 13 3 3 0 2 16 4 15 13 2
21 10 9 4 4 10 9 3 0 13 13 2 16 10 9 13 2 16 1 15 13 2
18 2 13 0 9 13 3 9 9 2 15 15 3 7 3 13 1 9 2
20 3 0 9 3 13 2 7 13 14 15 1 9 7 0 9 3 13 7 13 2
4 11 2 11 2
2 11 2
5 9 2 9 7 9
7 15 1 15 2 15 2 15
77 0 9 2 7 3 3 9 2 13 10 9 2 16 0 2 9 0 2 9 2 0 2 2 2 7 2 15 2 15 2 15 2 15 2 15 2 15 2 15 2 15 13 1 15 3 12 0 9 2 15 2 15 2 15 2 15 15 13 16 10 9 1 9 2 16 13 1 12 2 2 12 2 7 12 2 9 2
24 13 15 9 2 15 13 2 1 10 9 13 1 9 9 10 7 3 15 13 9 0 2 0 2
24 2 12 2 2 11 13 1 9 10 2 15 2 15 2 15 2 15 2 15 2 15 9 2 2
12 2 12 2 2 11 13 1 9 10 9 2 2
44 9 2 12 2 3 13 2 16 9 0 2 9 2 0 2 2 10 13 3 2 16 9 2 15 0 9 2 2 9 2 2 13 2 13 0 1 9 2 15 13 13 9 9 2
15 3 9 9 2 0 2 7 2 16 0 15 3 1 9 2
66 13 3 13 2 16 9 9 2 0 13 0 9 2 16 4 15 13 2 3 4 1 9 2 12 2 13 1 9 14 9 1 9 9 2 12 2 2 7 2 2 11 13 1 9 10 9 2 2 2 3 13 15 1 9 2 3 9 2 0 2 1 10 9 13 2 2
23 10 9 4 7 13 0 2 1 9 4 13 0 2 16 15 3 9 2 10 13 1 11 2
48 9 1 9 9 2 0 2 0 2 7 13 2 3 0 2 13 2 2 13 7 1 15 2 2 2 13 7 1 15 2 2 13 2 16 4 13 2 3 0 7 10 9 1 9 3 13 9 2
6 13 13 7 7 11 2
33 7 3 2 1 9 2 9 15 13 7 1 9 9 7 9 9 10 9 2 13 0 13 9 2 10 9 0 2 2 10 9 2 2
19 13 7 13 2 16 1 10 9 1 0 9 13 9 10 0 9 3 0 2
42 3 11 2 11 1 10 9 1 9 0 9 13 2 16 9 9 2 13 15 13 10 9 2 13 0 2 13 0 2 16 13 15 9 2 10 2 7 2 15 2 2 2
26 13 1 9 2 1 15 13 13 12 9 2 2 13 7 2 13 2 2 2 10 9 7 9 13 0 2
17 1 10 9 15 13 13 3 0 9 2 0 2 15 2 15 2 2
20 1 10 9 15 13 3 2 3 2 2 13 15 1 9 1 10 0 9 2 2
20 16 7 0 9 13 3 1 10 9 3 0 2 9 12 9 9 1 15 13 2
26 13 12 9 2 2 9 2 11 13 9 13 1 10 9 0 1 10 9 2 2 2 3 13 0 9 2
25 7 9 1 15 4 14 13 9 9 1 9 2 0 2 3 2 2 2 2 0 1 10 9 2 2
3 3 14 2
32 1 9 15 13 1 12 9 2 2 9 2 2 10 9 13 9 2 7 2 9 9 2 2 10 9 13 9 2 11 2 2 2
26 9 9 13 3 9 2 11 2 2 15 13 0 1 9 9 2 3 10 0 9 9 2 0 2 10 2
37 13 7 1 9 0 2 9 2 11 2 13 9 9 0 9 2 13 2 2 2 16 1 9 13 0 9 2 3 9 13 3 9 9 2 0 10 2
45 13 3 2 16 16 4 1 0 9 0 13 0 9 0 2 15 13 2 2 2 2 2 3 4 13 1 9 9 2 0 10 1 1 0 9 10 0 9 2 9 2 11 2 2 2
10 7 15 13 2 3 13 10 9 0 2
3 12 2 12
27 1 9 9 1 9 9 1 9 12 2 12 2 3 4 15 1 9 9 0 9 13 13 9 9 7 9 2
35 2 2 2 3 13 3 7 3 13 9 7 9 2 15 13 0 9 0 2 3 16 9 13 13 1 0 9 14 1 0 9 7 0 9 2
6 15 13 9 1 9 2
38 9 7 4 13 1 0 9 0 9 7 9 1 9 2 2 9 9 2 2 2 9 9 12 2 2 2 9 9 2 2 2 9 0 9 2 2 3 2
6 15 4 13 3 0 2
45 1 9 9 0 13 2 16 13 1 0 12 9 10 9 2 16 13 1 11 2 11 2 7 3 1 0 9 2 3 4 10 9 1 9 13 7 4 2 14 15 3 3 13 13 2
53 7 3 13 0 9 9 1 9 7 9 2 15 13 3 0 7 0 9 9 13 0 1 15 7 13 0 9 9 2 15 4 13 15 2 16 13 1 10 9 15 13 7 15 3 1 10 9 13 7 3 3 13 2
43 1 0 9 13 3 0 9 9 9 2 9 7 9 2 16 4 0 9 13 1 9 2 15 15 13 2 13 7 13 7 13 13 9 2 15 13 2 16 15 13 1 9 2
27 14 1 9 9 7 0 9 15 13 9 13 1 0 9 7 13 15 7 3 9 1 9 7 9 2 2 2
2 11 11
2 12 2
4 9 11 2 11
3 12 2 12
42 2 2 2 2 0 9 9 4 13 13 0 7 0 9 0 9 2 9 15 9 7 9 2 0 9 9 2 13 3 2 0 11 1 9 12 2 7 9 9 1 9 2
44 0 9 13 7 0 0 0 9 2 9 0 2 0 7 1 9 0 9 2 1 9 3 9 9 0 9 7 0 9 2 3 13 13 9 2 2 0 9 4 13 0 13 3 2
17 9 7 9 4 3 13 13 1 9 0 9 7 9 9 0 9 2
31 9 4 13 1 9 7 9 13 0 9 9 7 0 9 1 9 2 7 3 15 13 1 0 9 7 9 2 2 2 2 2
30 2 2 2 2 2 16 9 9 3 13 2 13 2 13 2 0 9 2 16 15 15 4 1 9 13 2 2 2 2 2
2 11 11
5 0 9 11 2 11
3 12 2 12
23 9 4 13 13 0 13 2 1 15 13 9 9 0 9 7 0 9 15 13 1 0 9 2
31 9 13 10 0 9 2 16 4 13 1 9 0 9 2 15 1 9 0 7 13 9 14 10 9 2 7 7 10 0 9 2
24 3 9 4 13 13 0 0 9 1 15 2 16 4 13 3 0 13 0 9 7 3 15 13 2
21 9 9 4 1 15 13 13 0 2 7 13 4 15 3 13 3 1 9 1 9 2
32 9 2 15 13 13 1 15 2 16 4 10 0 9 13 7 13 1 10 9 9 9 2 13 3 13 13 9 10 7 0 9 2
2 11 11
5 0 9 11 2 11
3 12 2 12
19 16 4 9 2 9 7 9 13 9 0 9 2 13 0 9 9 1 9 2
10 7 10 2 0 9 2 13 9 9 2
10 7 9 13 9 9 7 9 13 9 2
2 11 11
5 0 9 11 2 11
3 12 2 12
3 2 2 2
32 3 9 1 10 0 9 2 9 2 9 13 13 9 9 2 15 15 1 15 3 3 13 2 15 7 3 3 13 3 3 9 2
21 9 7 13 3 13 2 7 15 1 15 3 13 2 15 13 0 7 15 13 0 2
22 9 2 10 9 13 13 3 0 9 2 15 7 13 1 9 9 7 10 9 16 9 2
15 9 2 15 15 3 13 13 7 13 10 0 9 7 9 2
19 9 13 0 9 2 14 7 15 2 1 9 0 1 9 1 9 10 9 2
16 13 2 16 4 13 13 3 0 1 9 0 9 1 0 9 2
18 3 4 13 4 0 9 3 1 9 13 1 9 0 9 9 2 2 2
22 9 15 13 2 16 3 3 13 1 9 9 0 2 0 7 0 2 15 7 13 9 2
29 13 3 1 15 2 16 1 9 10 12 2 9 2 13 13 15 15 2 7 13 2 14 1 9 2 13 3 9 2
2 11 11
3 9 2 11
3 12 2 12
35 2 2 2 1 15 1 0 9 13 16 0 9 2 15 13 0 13 2 16 4 15 15 1 10 9 13 3 2 13 3 14 1 9 9 2
34 10 0 9 4 13 13 9 0 9 1 0 15 2 16 1 15 4 13 0 9 9 2 15 13 0 9 9 9 2 0 9 2 3 2
15 13 4 3 13 1 9 9 7 0 9 13 1 0 9 2
18 0 9 9 10 9 4 15 3 13 1 9 9 0 9 1 10 9 2
25 1 9 0 9 13 3 0 9 13 0 9 3 0 9 2 0 1 15 1 15 2 2 2 2 2
2 11 11
4 9 11 2 11
3 12 2 12
29 9 1 9 2 3 4 15 1 9 9 9 13 13 9 2 9 7 9 2 13 3 10 9 2 12 2 12 2 2
15 1 9 3 13 2 7 9 9 15 3 2 13 9 9 2
18 13 4 3 3 13 10 9 9 2 7 15 7 0 2 0 9 2 2
7 13 15 3 15 1 15 2
4 7 3 9 2
32 15 0 13 9 2 15 15 3 13 14 1 15 2 7 13 1 9 2 13 13 1 0 9 7 3 15 1 9 13 1 9 2
10 7 15 9 13 1 9 1 9 9 2
39 7 10 0 9 13 1 10 9 1 0 9 2 15 13 7 1 9 1 11 11 7 1 11 15 13 2 3 15 13 9 9 1 9 7 0 9 2 2 2
19 2 2 2 9 15 13 9 1 9 2 9 1 9 2 3 13 9 9 2
21 13 2 16 13 0 9 2 9 7 9 13 3 3 0 2 9 11 2 11 2 2
2 11 11
1 11
3 12 2 12
27 2 2 2 9 13 1 9 0 2 16 9 13 9 15 9 10 9 2 13 2 14 0 0 9 2 2 2
14 3 9 0 7 0 1 9 9 13 3 13 1 9 2
23 7 7 9 0 13 13 0 9 2 16 10 9 13 2 13 7 13 15 15 13 2 2 2
2 11 11
5 0 9 11 2 11
11 9 2 9 2 2 9 1 9 4 13 2
3 12 2 12
3 9 1 9
2 11 11
22 3 0 13 9 7 9 9 2 13 9 9 9 9 7 9 0 9 9 2 3 9 2
34 9 7 9 0 9 2 1 0 0 9 14 1 0 0 9 2 13 10 9 3 9 9 7 0 9 10 9 7 1 15 0 0 9 2
31 9 9 0 1 10 9 3 13 9 0 9 2 15 15 13 1 9 15 1 9 9 7 9 2 0 9 7 0 0 9 2
25 13 15 7 3 2 7 2 3 2 3 1 9 7 9 2 13 9 2 7 7 15 13 16 0 2
11 1 0 9 13 7 9 1 0 9 9 2
12 15 7 13 2 16 13 9 15 1 15 13 2
32 10 10 9 2 13 16 9 7 9 2 13 13 0 7 1 9 0 9 2 15 3 13 0 1 9 2 10 9 13 13 15 2
34 10 9 13 9 9 2 9 9 13 3 0 9 16 9 2 7 0 9 2 1 15 9 1 9 13 2 15 1 0 9 3 13 9 2
30 13 0 9 13 10 9 13 9 0 9 16 9 0 9 1 9 9 2 15 3 15 1 9 13 2 15 13 9 9 2
22 7 1 0 9 9 13 0 9 9 13 7 1 1 0 9 13 4 13 16 0 9 2
17 1 10 9 3 13 7 4 3 13 10 9 0 9 9 7 9 2
13 9 2 16 1 9 9 0 9 13 2 13 9 2
19 0 13 3 9 2 16 10 9 13 3 10 0 9 0 2 0 9 2 2
18 1 3 0 9 3 16 9 13 9 9 2 7 7 7 15 15 13 2
20 0 9 1 9 10 9 13 3 2 9 2 16 9 1 9 13 10 0 9 2
14 10 9 15 13 1 9 0 9 0 15 9 0 9 2
16 1 9 0 9 13 0 9 3 0 9 2 1 15 3 13 2
18 1 0 9 4 13 2 16 1 9 7 9 1 9 13 0 9 9 2
22 3 15 7 10 9 13 3 2 16 9 7 9 1 9 13 3 13 9 7 9 9 2
33 10 9 13 7 1 9 1 9 7 1 10 9 13 9 2 16 1 9 7 9 9 13 3 0 9 2 9 7 9 1 9 9 2
12 13 15 9 0 9 13 2 16 15 3 13 2
37 13 2 14 0 9 14 3 2 16 4 9 13 0 9 2 7 3 1 15 2 16 4 13 0 0 9 2 13 1 10 9 9 7 9 13 0 2
14 15 4 1 10 9 13 9 10 0 9 7 0 9 2
19 13 14 1 9 2 0 9 2 9 2 3 2 2 7 1 9 0 9 2
11 7 9 9 1 9 12 0 9 13 13 2
25 4 3 13 0 9 2 7 10 9 1 9 2 15 13 2 13 0 2 7 2 9 13 0 9 2
13 3 2 1 9 13 13 0 9 0 9 7 3 2
14 15 13 1 9 9 7 9 9 2 15 13 0 9 2
10 9 9 0 15 0 9 13 7 0 2
5 9 13 0 9 2
25 13 2 16 9 1 0 9 13 3 0 2 7 0 9 15 13 2 16 1 0 9 13 0 9 2
18 15 4 13 7 1 9 1 9 2 16 4 0 9 13 0 9 9 2
16 9 0 9 13 3 0 7 0 9 9 1 0 9 0 9 2
15 1 9 9 13 15 10 0 9 2 0 9 2 11 3 2
29 9 9 0 9 13 3 0 9 2 7 7 14 15 9 13 0 2 7 3 9 1 0 0 9 13 1 15 9 2
18 1 9 15 13 2 16 7 3 0 9 16 9 9 13 9 9 9 2
9 1 10 9 9 13 0 9 9 2
16 1 9 3 0 9 13 9 9 2 16 0 13 2 3 0 2
31 13 0 2 16 9 9 9 13 3 0 1 9 2 9 2 7 3 0 13 2 16 3 13 13 7 1 9 7 0 9 2
24 1 9 9 2 15 13 9 9 7 9 1 9 2 13 14 3 15 2 15 13 3 0 9 2
12 3 1 0 9 13 1 0 9 13 10 9 2
16 3 3 13 10 0 9 1 9 9 2 15 13 9 0 9 2
30 0 9 3 2 12 9 1 15 7 0 9 1 0 9 1 9 7 0 9 1 9 13 13 0 9 0 9 0 9 2
31 9 1 2 0 2 9 4 3 13 0 9 7 2 9 2 9 1 9 0 2 0 7 0 13 3 9 0 9 12 9 2
41 9 3 13 0 9 2 0 7 0 9 2 7 7 0 9 1 9 9 2 15 1 0 9 13 0 9 7 15 7 9 9 2 13 13 0 9 1 9 0 9 2
33 0 9 0 9 1 0 9 13 0 0 9 2 15 13 13 2 16 1 9 9 9 13 9 1 0 9 9 1 2 0 2 9 2
20 3 9 0 9 13 9 2 15 13 3 9 2 7 7 0 9 9 0 9 2
25 3 3 0 9 2 9 2 7 0 9 13 9 2 3 13 13 0 9 1 0 9 7 9 9 2
33 10 9 3 0 9 13 2 7 9 2 15 13 3 1 9 9 13 1 9 9 7 3 13 3 13 9 1 0 9 9 1 9 2
46 13 3 0 2 16 4 3 9 7 0 9 15 10 9 13 2 16 1 0 9 13 9 2 7 3 7 9 9 2 7 3 0 9 3 2 3 4 9 1 9 13 1 0 0 9 2
24 1 9 13 2 9 2 2 15 13 1 9 7 1 9 15 0 16 9 9 0 1 0 9 2
20 13 9 1 15 2 16 9 9 0 9 13 1 0 9 3 0 9 1 9 2
16 3 3 1 9 7 9 2 3 1 9 2 9 7 0 9 2
35 13 14 9 2 3 15 13 10 9 2 16 1 9 1 0 9 0 9 4 1 15 0 9 9 9 1 9 7 9 13 3 14 1 9 2
5 3 13 9 12 2
6 0 9 1 9 7 9
2 11 9
19 0 9 0 9 7 0 9 15 3 13 9 0 9 2 0 2 7 0 2
15 10 9 3 13 3 3 3 16 9 1 9 7 1 9 2
12 3 7 14 1 3 3 0 9 13 1 0 2
50 7 16 11 11 13 9 2 12 1 11 9 1 9 2 0 9 7 1 9 9 11 2 2 13 10 9 0 9 9 9 1 9 9 0 9 7 1 9 0 9 2 15 3 13 1 9 10 12 9 2
26 3 11 11 3 13 2 16 0 9 1 0 9 1 9 2 12 13 3 2 0 2 0 0 9 2 2
25 9 9 1 0 9 13 3 0 2 13 4 2 3 0 9 9 1 9 13 0 2 3 3 0 2
10 7 15 15 4 13 1 0 12 9 2
38 13 3 2 16 9 13 0 0 9 2 7 3 13 0 13 9 2 3 13 0 9 1 9 1 9 0 9 2 15 13 9 2 9 2 9 7 9 2
16 3 2 3 13 9 0 0 9 0 2 13 9 1 0 9 2
19 7 9 1 0 9 15 13 0 9 2 15 1 15 13 9 7 0 9 2
27 1 10 9 3 13 0 9 0 9 0 1 15 2 16 4 15 1 9 0 9 13 7 13 9 7 9 2
41 0 9 1 11 13 15 0 2 7 13 12 9 2 0 9 13 3 3 1 0 9 2 16 10 0 9 2 3 15 9 13 3 3 2 13 1 9 3 0 9 2
28 3 0 1 10 9 13 9 9 2 11 2 12 2 3 0 1 0 9 1 0 9 1 0 9 1 9 9 2
13 3 15 15 13 9 2 3 3 9 7 0 9 2
5 14 15 13 9 2
37 15 4 1 15 3 13 7 10 0 9 2 7 9 2 7 9 2 3 14 3 0 9 2 14 16 16 15 1 9 13 9 2 15 4 3 13 2
6 7 13 15 0 9 2
18 3 15 13 2 16 15 1 9 13 2 15 3 13 3 3 1 9 2
17 1 9 9 13 10 9 2 16 13 3 3 16 9 12 1 11 2
15 13 3 1 0 0 9 10 9 1 9 14 12 0 9 2
11 3 13 15 3 0 9 16 10 1 11 2
28 0 9 13 1 9 1 0 9 15 0 2 7 0 9 1 0 9 13 0 9 1 9 12 7 12 0 9 2
17 3 0 9 13 15 1 9 1 9 12 0 9 2 12 2 2 2
17 3 4 15 1 15 13 13 14 12 9 9 2 16 13 10 9 2
34 7 10 9 13 3 2 3 14 1 9 9 9 2 3 4 13 9 9 7 9 9 2 0 14 12 9 9 2 14 3 0 0 9 2
27 0 9 13 1 15 1 0 9 9 14 12 9 2 9 7 1 15 13 9 2 3 15 3 9 13 3 2
5 13 15 0 9 2
13 0 9 13 3 9 9 2 1 10 9 15 13 2
23 1 9 1 0 15 9 1 12 9 15 9 3 13 9 2 16 15 15 13 13 9 9 2
8 13 15 2 9 1 9 2 2
19 16 13 1 10 9 1 9 2 0 9 2 13 0 9 2 9 1 9 2
23 7 3 2 13 1 9 2 16 3 2 14 3 2 13 9 9 1 12 9 0 0 9 2
36 11 11 7 11 11 2 15 1 10 9 13 7 0 13 1 2 0 9 2 2 13 2 16 1 9 9 13 3 13 1 0 9 7 9 9 2
23 0 9 13 9 1 0 0 9 7 9 0 0 9 2 15 3 3 3 13 1 9 11 2
12 15 15 13 3 2 16 9 1 9 9 13 2
20 15 15 3 13 0 7 0 9 0 11 2 11 2 1 9 9 2 11 2 2
22 0 9 9 13 1 9 9 7 9 10 0 2 7 0 0 9 1 12 9 3 9 2
34 0 9 13 3 3 0 1 0 9 2 1 0 9 1 9 1 0 11 13 0 9 3 10 9 2 16 7 0 9 4 3 13 9 2
18 10 9 13 7 0 2 7 9 13 0 9 7 9 9 1 15 0 2
17 9 2 1 9 1 0 0 9 9 2 13 1 9 9 0 9 2
21 0 13 0 9 3 9 7 1 15 13 0 9 2 0 10 9 9 0 9 9 2
15 13 1 15 12 0 9 0 9 9 7 12 9 9 9 2
14 0 0 9 9 13 3 0 2 3 13 9 1 11 2
23 0 9 15 0 9 13 3 13 2 15 15 13 3 10 0 9 2 7 7 9 1 15 2
12 9 9 13 0 7 0 9 9 1 15 9 2
22 3 15 3 3 13 1 9 1 0 9 15 2 15 13 1 3 0 9 3 1 9 2
5 13 15 0 9 2
11 15 3 0 9 13 13 0 9 7 9 2
15 13 7 2 16 3 9 3 13 0 9 2 1 15 13 2
13 0 9 15 13 3 13 10 9 1 9 7 9 2
21 3 10 0 7 0 9 15 13 1 0 9 2 3 13 9 2 1 15 15 13 2
20 13 3 9 2 16 15 7 15 9 3 13 13 2 16 15 13 3 1 9 2
18 3 0 0 9 4 15 3 13 1 9 2 7 9 15 15 15 13 2
11 7 10 9 13 14 13 2 3 13 13 2
21 7 9 13 1 9 12 0 0 9 2 3 15 3 13 1 0 9 0 7 0 2
24 0 9 3 13 3 9 2 7 0 9 9 9 9 1 9 13 0 9 7 9 0 9 9 2
16 3 15 0 9 3 13 1 9 9 3 0 16 9 1 9 2
41 0 9 10 0 9 0 9 13 11 2 3 3 9 2 12 11 11 13 12 0 9 2 0 16 15 9 9 3 13 1 9 1 0 0 9 0 9 1 0 9 2
15 10 0 0 9 13 7 0 7 13 14 12 9 9 0 2
18 10 0 9 13 9 7 0 9 1 9 9 12 2 14 9 9 0 2
20 7 16 13 2 1 15 3 13 0 9 2 0 15 3 1 9 1 0 9 2
19 9 1 2 0 9 2 1 9 7 13 15 3 9 0 1 9 0 9 2
15 1 9 0 9 13 9 2 15 13 0 3 7 0 9 2
23 13 15 9 0 2 9 0 2 7 13 15 9 3 1 9 2 3 13 9 7 0 9 2
4 9 13 9 2
8 2 9 1 9 15 13 2 2
10 16 9 13 1 9 2 3 0 13 2
22 9 13 3 0 14 12 2 12 2 12 9 2 2 2 2 7 0 12 2 12 9 2
31 16 13 0 9 9 1 9 1 9 2 9 13 0 9 9 2 1 15 13 9 0 9 7 13 13 1 9 9 0 9 2
25 15 15 1 9 13 9 9 2 1 15 15 13 2 13 7 13 16 10 0 9 15 1 9 13 2
17 1 9 3 0 9 1 12 9 13 7 1 9 15 15 3 13 2
15 1 10 9 15 3 0 7 3 0 9 13 3 1 9 2
30 10 9 13 3 13 1 0 9 11 2 11 7 1 12 9 11 2 1 9 1 9 0 11 2 1 9 11 7 11 2
17 3 15 1 9 13 0 2 0 9 0 2 9 1 2 9 2 2
28 16 9 1 9 1 9 13 10 9 2 13 15 1 0 9 7 3 2 3 13 16 15 0 13 1 9 3 2
39 10 9 4 1 9 3 13 0 9 7 7 2 3 2 10 9 15 13 2 16 10 9 13 1 15 3 0 2 16 15 9 1 0 9 13 3 9 9 2
23 2 14 3 10 9 7 9 0 2 16 15 3 13 2 13 9 12 2 12 2 12 2 2
36 1 9 12 4 1 0 9 0 9 7 15 0 9 0 9 2 0 9 7 0 0 9 13 9 0 9 10 9 1 9 0 1 9 9 12 2
17 13 15 2 3 2 16 4 15 1 15 13 13 14 1 10 9 2
22 1 0 9 0 0 9 4 9 13 3 9 2 12 7 1 11 3 2 9 2 12 2
27 1 0 12 9 4 13 7 1 0 11 7 1 11 7 3 3 2 7 11 2 11 2 11 2 11 3 2
18 1 3 0 13 0 2 16 0 9 1 9 13 9 0 9 1 9 2
11 15 7 13 1 10 9 1 3 9 0 2
17 7 7 16 7 3 13 9 9 3 2 10 9 15 3 3 13 2
13 3 13 3 0 0 9 9 7 0 9 1 9 2
10 0 7 0 9 9 3 13 9 9 2
20 7 7 15 1 9 13 9 13 1 9 9 2 15 4 15 9 1 9 13 2
14 1 0 9 10 9 13 15 3 2 3 15 9 13 2
20 16 1 0 9 13 9 9 1 11 1 9 10 0 9 2 13 1 0 9 2
30 0 9 15 13 1 11 7 16 1 9 9 13 14 1 12 9 2 3 1 0 9 0 9 2 9 2 13 3 0 2
9 15 7 13 0 9 1 9 9 2
15 15 15 3 3 13 15 2 15 15 13 3 3 10 9 2
20 16 15 2 15 1 15 13 7 15 15 1 15 3 13 2 1 10 9 13 2
6 16 13 15 2 9 2
11 2 0 11 9 2 12 2 12 2 12 2
6 7 15 15 3 13 2
13 14 16 15 15 13 3 2 3 4 1 11 13 2
8 15 1 15 2 9 9 2 2
9 1 9 13 3 12 3 0 9 2
18 16 4 15 13 2 14 2 9 2 13 9 12 2 12 2 12 2 2
2 11 11
3 12 2 12
3 9 13 9
4 0 9 13 11
2 11 11
32 3 7 3 13 9 9 2 15 15 13 13 1 10 9 3 1 9 1 12 9 2 10 9 13 13 1 0 9 7 11 2 2
10 13 1 0 11 7 13 15 9 9 2
25 13 13 11 3 10 0 2 0 2 9 7 13 14 1 0 9 0 1 3 0 2 0 9 2 2
22 1 9 0 9 7 3 3 14 1 11 13 9 9 0 2 0 3 3 16 9 0 2
26 0 13 3 12 9 2 0 3 0 2 14 9 13 3 0 1 0 9 7 1 9 13 12 0 9 2
6 10 0 9 13 0 2
16 16 4 15 13 1 0 9 2 13 4 15 2 9 0 2 2
38 13 3 1 9 9 2 10 9 4 1 0 9 3 13 1 2 9 2 2 15 13 2 2 2 16 4 3 4 13 1 2 0 2 9 1 9 9 2
45 13 15 3 9 10 9 9 0 2 15 13 0 0 9 1 0 9 7 9 2 15 1 0 9 13 9 15 2 16 13 0 9 1 9 1 9 2 3 9 13 3 9 1 9 2
9 9 15 13 3 16 2 9 2 2
4 3 3 14 2
7 10 9 14 13 10 9 2
19 16 10 9 15 13 13 9 1 0 9 2 0 9 13 9 1 0 9 2
11 3 1 0 9 0 9 7 3 7 9 2
8 1 9 1 15 13 9 9 2
16 9 15 13 1 9 7 9 9 7 15 13 1 0 9 9 2
25 9 4 13 7 9 1 0 9 2 0 9 0 9 2 3 7 3 0 9 1 9 9 7 9 2
15 3 0 9 16 9 2 0 9 9 7 9 13 9 9 2
19 1 9 15 3 13 9 2 15 15 3 13 1 0 9 2 15 15 13 2
6 13 7 0 0 9 2
15 16 0 9 13 0 9 1 9 2 13 9 13 9 9 2
4 15 13 3 2
16 1 10 9 9 13 12 9 2 13 9 7 1 9 15 13 2
11 1 0 9 13 0 0 9 3 12 9 2
13 9 1 0 9 4 13 1 10 9 9 9 3 2
28 1 0 12 9 15 7 9 13 1 10 9 3 13 7 15 0 9 2 15 15 3 13 3 14 1 10 9 2
22 9 10 9 4 3 3 13 2 16 13 0 15 3 7 1 0 9 13 1 0 9 2
5 10 9 9 3 2
31 1 9 4 3 13 3 0 9 2 15 4 3 1 9 13 9 2 15 13 10 9 1 9 2 7 13 2 16 13 0 2
23 1 9 15 13 1 0 9 7 13 3 1 3 10 0 9 9 2 15 13 0 9 13 2
27 3 15 10 9 13 1 0 9 1 9 11 7 11 1 9 11 7 3 15 10 9 13 7 1 0 9 2
18 3 4 1 11 10 9 3 13 7 0 9 15 13 7 1 0 9 2
12 1 0 9 9 1 12 9 15 3 13 3 2
21 1 11 1 9 12 13 1 11 1 11 2 11 2 13 0 9 9 9 10 9 2
9 0 9 9 3 3 3 15 13 2
11 9 13 4 3 13 1 9 0 1 11 2
45 1 9 0 9 4 13 0 12 9 2 15 1 0 9 13 1 15 12 3 7 15 14 1 9 2 9 2 9 2 9 2 9 2 9 2 7 7 9 7 9 7 3 14 9 2
22 3 1 0 9 13 13 3 1 12 9 9 9 9 2 15 13 3 14 9 0 9 2
20 0 13 1 9 1 12 9 1 12 9 7 4 1 15 13 12 7 12 9 2
14 0 12 5 13 9 1 12 9 2 7 15 3 0 2
18 13 15 9 2 16 9 2 15 15 0 9 1 9 13 2 9 13 2
32 9 10 9 15 0 9 13 1 9 0 9 1 9 7 9 2 11 2 2 16 15 1 0 12 9 13 0 9 16 1 11 2
23 1 10 9 4 13 9 12 9 9 2 13 9 1 11 7 11 7 13 4 13 0 9 2
12 0 9 13 3 13 7 13 9 9 1 9 2
14 13 3 1 15 2 15 4 4 0 13 1 0 9 2
27 7 1 9 2 3 4 9 13 2 15 0 9 1 15 2 16 10 9 13 3 0 9 2 13 13 0 2
9 0 9 1 10 9 15 15 13 2
39 9 9 13 13 1 3 12 9 0 2 7 3 0 9 1 9 2 0 15 1 9 1 11 1 9 11 7 13 15 2 16 0 9 13 1 10 9 0 2
1 9
3 9 1 9
18 9 3 0 2 3 0 2 7 1 9 0 9 9 15 3 3 13 2
48 13 15 3 1 0 0 9 2 3 15 13 3 1 9 16 9 0 2 2 9 9 9 2 2 7 15 3 1 9 2 9 7 9 2 9 12 2 12 2 12 7 12 2 12 2 12 2 2
32 9 9 0 11 2 11 2 11 1 0 9 1 9 2 11 2 15 3 1 10 9 13 13 2 16 1 0 0 9 13 9 2
17 9 0 2 9 0 2 13 3 3 1 0 7 0 9 0 9 2
21 16 13 3 1 9 2 0 9 15 13 1 2 9 2 2 0 2 0 9 2 2
19 3 3 7 13 2 14 9 13 1 9 9 7 9 3 0 9 1 9 2
27 1 9 10 9 13 3 12 9 9 0 9 2 16 13 9 0 2 3 10 9 0 1 0 9 0 9 2
21 10 9 13 1 15 2 16 15 15 1 9 13 13 9 1 9 0 9 9 9 2
10 13 4 15 13 0 9 0 0 9 2
23 13 2 16 10 0 9 13 0 9 16 9 9 1 9 2 11 12 2 12 2 12 2 2
2 11 11
3 12 2 12
8 9 2 3 14 9 1 9 2
28 1 9 9 15 13 9 2 16 9 9 7 9 13 2 7 13 4 13 16 9 1 9 2 7 3 3 13 2
9 3 15 9 13 3 1 0 9 2
18 15 0 4 15 13 13 16 11 1 10 9 2 0 9 1 9 2 2
40 9 2 9 2 15 13 13 3 2 0 11 12 2 12 2 12 2 7 13 0 9 1 0 9 2 7 14 2 1 9 12 2 12 9 2 3 10 0 9 2
7 9 9 13 3 0 9 2
59 0 9 9 13 10 0 9 13 2 0 9 13 1 12 15 9 1 9 2 12 2 7 9 13 14 12 2 7 9 13 13 12 0 7 12 0 9 2 15 15 1 10 9 13 13 2 1 0 9 0 15 12 9 2 0 2 9 2 2
33 0 13 9 9 1 11 2 0 0 0 9 13 13 3 9 2 7 9 9 1 9 9 9 7 9 1 9 15 13 1 0 9 2
19 0 9 13 1 0 2 0 2 9 2 3 0 9 15 1 10 9 13 2
33 4 15 0 9 13 0 9 2 7 15 4 13 0 9 7 15 0 2 1 0 9 2 4 13 2 7 13 1 9 2 3 3 2
2 11 11
3 12 2 12
4 1 9 1 9
10 1 9 11 2 11 2 1 9 2 2
8 9 12 2 12 2 12 2 12
8 9 12 2 12 2 12 2 12
19 1 9 2 15 13 9 2 2 4 13 9 13 2 16 9 13 3 13 2
21 13 15 14 13 1 15 2 16 9 2 7 15 14 10 2 13 0 2 7 14 2
10 13 3 3 12 9 2 9 7 9 2
19 13 15 3 2 16 1 9 13 0 9 7 9 4 3 13 16 0 9 2
13 3 16 13 1 9 9 2 7 3 1 0 9 2
15 3 4 3 13 1 9 2 16 9 13 0 9 0 9 2
17 3 15 3 13 9 9 2 16 13 9 2 16 3 13 0 9 2
17 3 7 13 2 3 13 2 16 9 13 2 7 16 13 3 0 2
16 2 0 4 3 13 1 9 9 1 9 7 9 0 9 2 2
37 1 10 9 3 13 1 3 0 9 16 1 0 9 0 9 2 15 13 2 3 13 2 2 7 3 13 10 9 3 0 1 9 7 9 0 9 2
12 11 2 11 9 13 7 3 13 9 1 9 2
35 2 9 16 9 1 9 2 13 12 9 2 1 12 9 9 7 9 2 15 13 9 7 1 0 9 9 2 1 15 10 9 13 7 3 2
16 0 13 2 16 15 13 13 9 2 15 13 1 9 0 9 2
8 9 13 10 9 1 0 9 2
14 10 9 2 16 13 3 3 0 2 13 12 0 9 2
4 3 3 13 2
42 1 0 9 2 15 13 10 9 2 13 3 3 13 10 9 2 16 15 13 1 9 0 0 9 13 1 0 9 2 9 2 9 7 15 1 10 9 7 9 0 9 2
15 1 10 9 3 3 13 0 13 3 0 9 9 7 13 2
21 12 2 10 9 13 2 3 2 13 2 16 13 2 3 2 13 13 1 9 0 9
31 12 2 10 9 13 2 3 2 13 0 2 16 9 10 9 1 0 9 15 13 2 16 13 2 3 2 13 1 0 9 2
20 3 3 0 9 13 15 0 16 9 2 15 4 13 13 0 1 10 9 2 2
8 3 3 13 0 9 1 9 2
17 3 0 9 13 1 0 9 0 2 0 2 2 2 2 2 9 2
13 9 1 9 10 3 0 9 3 13 0 9 9 2
13 9 15 13 13 3 3 2 16 0 9 13 3 2
14 3 2 16 9 10 9 13 1 10 0 9 7 9 2
17 13 15 3 0 9 1 9 2 2 9 2 2 7 10 0 9 2
26 2 9 9 13 1 10 9 2 16 0 9 13 9 2 15 13 10 9 7 10 9 2 3 0 2 2
15 10 9 1 9 2 13 2 1 9 9 7 9 13 0 2
77 13 2 14 15 3 9 10 9 2 10 9 2 9 2 13 15 3 3 1 9 2 3 13 13 0 9 9 2 15 4 13 9 1 9 0 2 13 2 0 9 0 2 0 2 2 2 2 2 9 2 2 7 13 3 1 2 9 2 2 3 0 9 2 15 13 3 9 2 2 7 3 1 9 2 9 2 2
20 1 9 0 2 0 2 9 2 7 3 3 1 15 2 13 3 0 9 3 2
50 13 9 2 1 10 9 15 3 9 9 13 1 9 3 3 0 9 2 15 1 0 2 7 1 0 2 3 10 9 2 0 1 9 2 15 13 3 0 9 7 0 9 2 13 1 15 1 0 9 2
17 1 0 9 3 13 12 9 9 7 13 15 3 13 12 0 9 2
31 1 0 9 10 9 2 15 13 0 1 10 9 3 3 2 16 13 1 9 2 15 1 10 9 13 13 1 0 3 3 2
19 15 13 3 10 9 2 3 9 0 7 0 3 3 0 2 2 2 9 2
21 7 1 0 9 2 13 4 0 2 7 16 4 15 13 1 9 2 13 2 0 2
12 0 9 13 9 2 15 9 14 3 0 13 2
19 3 3 1 10 9 4 13 0 13 7 13 2 16 13 7 16 13 0 2
60 9 12 9 15 3 13 7 15 2 16 12 9 13 2 16 9 13 2 16 13 3 0 2 7 13 15 3 13 9 1 2 7 3 13 13 1 9 2 16 9 13 2 13 1 15 7 0 9 2 7 13 1 12 0 9 3 7 13 15 2
9 13 2 15 13 9 9 1 9 2
22 16 7 15 13 2 16 9 13 9 1 9 2 3 15 3 1 10 0 9 13 9 2
19 9 15 2 15 3 13 2 15 13 10 9 2 1 15 13 15 0 13 2
2 11 11
3 9 1 9
9 1 15 15 13 1 9 7 1 15
6 0 9 0 9 0 9
20 1 0 9 4 15 13 1 3 0 9 0 9 1 9 2 9 2 11 11 2
15 0 9 1 9 7 9 13 1 15 9 1 0 0 9 2
10 15 9 1 10 9 13 1 0 9 2
17 11 11 11 2 0 9 9 2 15 13 12 2 9 12 1 11 2
15 9 13 1 0 9 7 3 13 1 0 0 9 1 9 2
23 0 2 9 2 13 11 1 0 11 2 9 1 11 2 11 1 11 2 16 3 0 9 2
9 3 13 10 9 0 1 0 9 2
12 1 10 9 13 9 2 9 2 9 7 9 2
22 11 11 2 0 9 9 2 13 9 10 0 9 1 9 11 2 7 15 1 9 12 2
15 0 9 13 1 0 9 0 9 2 3 13 13 16 9 2
8 9 12 15 3 13 0 9 2
21 9 12 13 1 0 9 2 7 3 10 9 15 3 13 1 11 1 11 1 11 2
7 9 12 15 3 13 9 2
6 11 11 13 12 9 2
19 13 15 1 0 9 11 2 13 1 11 2 3 15 9 2 12 13 9 2
11 3 0 9 13 1 11 1 11 1 11 2
17 3 12 9 3 13 1 10 9 2 1 15 14 2 13 3 2 2
29 7 1 15 3 3 1 10 0 0 9 1 0 9 0 9 2 13 9 1 9 2 12 2 12 1 10 9 2 2
4 0 9 13 0
21 1 9 13 1 11 2 1 11 0 11 1 11 9 11 12 0 9 0 0 9 2
14 9 2 3 1 0 9 9 11 11 2 3 13 3 2
9 13 3 3 13 9 1 0 9 2
35 9 0 9 3 3 3 13 1 0 9 2 9 9 7 9 15 13 1 12 5 9 2 16 1 9 3 0 9 13 3 10 9 12 5 2
11 9 13 14 3 12 9 2 7 3 12 2
6 15 0 13 9 0 2
15 7 9 15 3 3 13 9 2 16 13 13 1 9 3 2
9 9 9 13 9 1 9 0 9 2
13 9 4 13 3 9 0 9 1 11 7 9 11 2
24 0 0 9 4 3 1 9 13 9 2 12 1 0 0 11 1 9 9 7 3 1 0 9 2
10 0 9 13 12 9 0 0 9 9 2
20 13 2 16 15 13 9 1 0 9 2 15 10 9 13 13 2 3 9 0 2
11 0 9 13 2 16 4 15 1 9 13 2
14 0 9 13 10 9 13 2 16 10 9 4 13 12 2
17 7 3 15 13 3 13 1 9 9 1 0 9 2 3 2 9 2
5 13 9 9 9 2
30 9 9 7 9 9 13 0 9 13 0 9 2 16 9 11 2 15 13 2 13 13 13 1 9 7 13 15 3 9 2
20 11 2 15 15 13 1 11 9 0 11 11 2 13 3 0 0 9 1 9 2
18 13 15 1 9 2 15 9 13 13 1 9 0 0 9 1 9 9 2
9 10 9 13 0 9 9 1 9 2
18 7 9 1 10 9 0 9 4 13 13 0 1 9 2 9 0 9 2
12 9 9 15 7 13 9 9 0 2 7 0 2
16 7 7 9 13 16 13 2 16 11 4 13 9 1 10 9 2
15 16 15 7 4 13 10 0 9 13 7 9 15 15 13 2
15 15 3 13 0 9 1 9 0 9 1 9 9 0 9 2
30 7 7 13 0 2 16 0 11 15 10 9 4 13 13 13 2 15 15 15 3 3 13 2 16 13 3 10 0 9 2
24 13 13 3 1 15 2 16 15 3 13 13 11 2 7 14 3 10 9 2 1 15 13 3 2
6 9 15 3 3 13 2
11 9 9 15 13 1 9 1 9 9 0 2
21 15 13 3 0 9 0 9 1 9 9 2 15 13 0 9 15 9 1 9 9 2
24 9 0 0 9 0 9 13 1 9 9 1 9 10 9 2 13 15 2 16 4 13 3 9 2
32 9 0 11 13 7 13 2 16 9 1 9 9 2 15 15 15 3 13 2 4 3 13 13 0 9 2 3 7 10 9 9 2
6 0 9 13 2 2 2
10 7 11 1 10 9 3 13 2 2 2
4 0 9 1 9
12 1 0 9 3 3 13 1 0 2 0 9 2
8 9 13 13 2 0 9 2 2
33 13 15 1 9 0 9 2 1 9 15 13 9 2 13 1 9 2 13 9 7 3 2 3 13 2 13 9 7 15 13 1 9 2
5 13 15 16 9 2
11 1 11 13 10 0 9 1 9 0 9 2
17 16 13 1 10 2 9 2 2 13 9 9 1 9 3 0 9 2
12 13 1 0 9 1 9 9 2 9 1 9 2
8 1 9 13 15 16 0 9 2
46 9 3 13 2 16 13 1 9 2 13 15 9 2 13 9 1 9 1 9 2 13 2 13 1 15 2 15 15 13 3 2 16 13 9 1 0 9 2 13 2 15 13 3 2 2 2
20 7 9 3 13 10 9 2 3 15 15 13 9 2 16 13 9 1 0 9 2
23 1 9 9 2 9 1 9 2 15 1 0 9 13 0 9 2 15 15 13 13 1 9 2
18 10 9 0 9 15 13 13 7 1 9 9 7 1 9 9 1 9 2
5 0 9 1 9 9
14 1 9 0 9 11 11 4 15 3 1 9 13 3 2
24 10 0 9 1 11 1 9 2 12 3 13 1 9 10 9 2 15 13 9 0 9 3 3 2
18 1 9 0 9 13 0 9 3 3 2 16 0 9 13 16 9 9 2
6 9 13 9 0 9 2
21 11 15 15 13 3 1 9 0 9 2 16 7 1 0 11 13 1 10 0 9 2
19 0 7 1 15 13 2 16 13 0 9 9 2 15 13 0 9 0 9 2
10 15 15 3 0 9 9 13 2 2 2
19 11 13 9 1 0 9 2 13 15 2 13 0 9 9 2 13 0 9 2
6 9 15 7 3 13 2
19 7 3 13 9 2 1 15 3 13 2 13 1 10 9 1 0 0 9 2
20 1 10 9 13 15 1 0 9 13 13 2 16 4 13 9 1 0 0 9 2
7 13 1 15 12 2 9 2
9 13 15 9 9 0 9 11 11 2
6 9 9 13 0 9 2
11 9 2 9 9 2 13 10 9 7 9 2
9 9 13 2 9 15 13 14 3 2
28 16 7 13 9 1 9 0 9 1 0 2 15 15 13 7 9 13 2 2 9 2 13 9 7 15 13 2 2
4 0 13 3 2
22 15 2 15 13 1 9 2 13 3 2 11 13 1 9 7 15 13 1 9 10 9 2
13 11 15 3 13 1 9 9 2 1 9 10 9 2
18 7 9 9 2 16 10 9 13 1 0 9 2 13 1 15 0 9 2
13 15 13 9 14 1 9 0 9 7 14 1 11 2
32 0 9 1 11 13 7 9 0 0 0 9 1 12 2 9 13 1 0 9 11 11 2 9 9 0 9 7 9 0 9 9 2
18 12 2 9 4 11 2 11 13 9 9 9 0 9 1 9 0 9 2
40 9 13 3 1 11 11 1 0 9 2 16 11 13 9 2 12 1 0 9 1 9 0 9 7 16 11 3 13 0 0 9 1 11 1 9 0 9 11 11 2
37 13 1 15 9 2 16 12 9 9 2 15 11 13 1 11 1 9 0 9 2 4 3 13 1 9 0 0 9 2 7 3 7 1 9 0 9 2
15 11 2 11 13 4 13 2 0 9 13 13 0 12 9 2
7 9 1 0 9 13 0 2
22 3 2 15 13 2 16 0 11 13 0 9 1 9 0 9 2 7 0 9 0 9 2
16 0 9 0 1 9 13 1 9 1 9 15 13 3 3 13 2
20 9 7 13 2 16 11 13 0 9 7 16 9 13 13 1 10 9 1 9 2
18 7 9 9 15 13 14 12 2 9 13 9 9 9 13 9 1 9 2
5 7 9 15 13 2
22 9 9 9 9 11 2 11 1 0 9 13 9 11 1 9 0 9 7 9 10 9 2
11 9 1 0 9 1 0 9 3 13 0 2
3 9 0 9
31 13 15 1 9 10 10 9 2 1 10 9 15 15 13 13 1 10 0 9 1 0 9 2 3 13 0 0 0 0 9 2
11 1 0 9 15 13 9 3 1 0 9 2
7 7 3 13 1 0 9 2
21 9 0 9 15 13 1 11 2 16 4 3 13 1 12 0 9 7 12 0 3 2
12 2 3 0 0 9 13 9 9 0 9 11 2
22 13 1 9 2 1 15 4 1 9 0 0 9 13 9 2 2 13 15 0 0 9 2
10 15 13 1 3 3 0 9 3 3 2
29 9 11 15 1 10 9 13 1 11 2 11 7 1 3 2 0 2 9 11 2 11 7 11 2 3 1 12 9 2
26 3 2 9 11 2 11 2 9 0 9 0 9 9 13 11 1 0 9 10 0 9 12 2 12 9 2
22 1 0 0 9 15 1 12 9 13 9 9 9 2 0 9 7 9 0 9 1 9 2
4 13 1 9 2
10 10 0 9 15 13 1 3 0 9 2
11 15 13 9 9 9 0 9 7 15 9 2
21 15 7 13 13 3 2 0 9 1 11 1 11 2 15 13 1 9 10 0 9 2
13 0 9 12 2 12 9 13 1 10 9 0 9 2
14 7 3 13 9 2 16 13 1 9 1 9 2 2 2
17 11 2 11 15 13 3 2 2 11 13 9 2 13 7 13 9 2
11 7 15 4 13 13 9 10 0 9 2 2
7 7 2 3 1 15 13 2
6 0 9 3 13 9 2
11 0 9 13 3 13 1 12 2 12 5 2
16 9 13 3 13 1 9 12 9 2 15 13 3 16 0 9 2
19 7 7 15 13 9 7 1 0 9 9 7 9 1 0 9 9 1 9 2
18 3 2 3 12 2 9 9 0 9 9 13 1 11 9 9 1 11 2
20 9 15 13 9 9 1 11 2 11 2 11 2 11 2 11 2 11 2 2 2
22 9 11 2 11 9 0 9 9 11 11 1 9 9 11 11 13 13 9 9 13 9 2
10 7 3 0 9 9 13 0 9 9 2
21 16 13 0 9 0 0 9 2 9 2 12 13 11 13 12 0 7 12 0 9 2
11 13 15 13 3 12 0 7 12 0 9 2
11 13 15 1 12 9 1 11 9 2 12 2
18 0 9 9 9 13 2 1 0 12 9 15 13 13 0 9 1 9 2
11 12 0 9 3 1 0 9 13 1 0 2
21 11 13 1 9 15 2 3 2 11 15 13 13 1 0 9 14 12 5 0 9 2
14 1 0 9 13 13 9 3 1 9 0 9 1 11 2
15 9 1 0 0 9 2 11 2 11 7 0 11 3 13 2
21 7 3 0 12 9 9 1 9 12 9 13 3 0 9 1 9 0 0 9 11 2
7 9 9 2 0 2 1 9
2 0 9
10 0 9 1 9 13 3 11 7 11 2
13 13 10 9 2 16 4 1 0 9 13 0 9 2
12 7 13 7 9 2 9 7 9 7 0 9 2
30 9 1 11 4 13 1 0 9 12 9 7 7 15 10 9 13 1 0 9 0 9 1 9 9 10 9 2 0 9 2
26 9 13 0 9 2 11 1 11 2 0 0 9 1 11 7 0 0 9 1 10 9 1 12 9 9 2
13 13 15 9 0 7 0 9 0 1 9 9 9 2
5 9 9 2 0 9
13 9 9 1 0 9 13 0 9 0 9 1 11 2
19 0 9 15 13 3 1 0 9 1 9 0 9 7 1 9 9 0 9 2
5 9 13 3 0 2
12 0 0 9 15 13 2 7 13 7 0 9 2
16 9 15 1 0 9 3 13 7 0 9 9 7 9 15 13 2
36 9 7 13 3 13 2 10 9 15 1 0 15 9 9 13 15 0 9 9 7 3 15 3 13 9 0 9 9 7 15 0 2 0 2 9 2
17 0 9 7 1 9 0 11 3 3 14 13 9 9 0 0 9 2
6 0 9 1 0 9 9
19 9 15 13 1 12 1 9 2 15 3 13 1 9 10 9 9 0 9 2
21 0 7 0 9 3 13 9 9 9 9 1 10 9 1 9 9 12 2 9 12 2
13 13 1 15 9 9 1 12 0 9 1 0 9 2
13 9 13 2 16 9 9 9 1 9 15 3 13 2
29 1 9 4 1 0 9 13 1 15 2 16 4 9 9 1 9 9 13 13 9 9 2 12 7 3 3 4 13 2
30 9 7 3 13 2 10 9 15 1 0 9 13 0 9 7 0 9 2 15 3 13 1 0 15 9 9 9 10 9 2
11 1 0 9 13 15 9 9 9 0 9 2
5 13 9 1 11 2
18 1 0 9 0 9 13 9 1 0 9 1 0 9 1 11 1 11 2
9 13 1 9 9 1 9 12 9 2
32 0 9 9 0 9 1 15 3 13 2 16 9 13 3 13 3 2 16 3 13 3 9 13 0 9 7 9 1 3 0 9 2
29 11 15 3 13 13 13 1 15 10 9 7 13 15 1 9 9 9 2 3 3 14 12 0 2 13 3 1 9 2
36 7 0 9 13 2 16 9 9 1 11 7 3 1 0 9 13 10 9 1 9 0 9 2 16 4 3 9 0 9 13 9 10 9 2 2 2
7 16 9 1 9 4 13 2
6 13 4 15 12 9 2
22 13 4 0 10 9 13 3 3 1 9 1 9 0 9 2 2 13 15 3 0 9 2
3 9 13 9
16 1 9 4 3 13 1 0 7 0 9 1 11 1 9 12 2
11 1 3 0 0 9 13 0 9 3 9 2
14 7 13 15 2 16 0 9 13 3 9 16 15 13 2
21 1 12 9 9 13 3 0 9 2 12 9 2 11 15 10 9 3 3 13 2 2
12 10 0 9 7 3 13 1 9 1 12 9 2
24 3 15 15 13 1 10 0 9 2 3 15 3 13 1 9 9 9 7 3 3 7 0 9 2
8 13 1 9 3 3 0 9 2
13 9 13 7 13 1 9 10 0 2 3 0 9 2
11 7 3 2 9 3 13 2 13 15 9 2
9 7 7 9 9 9 15 3 13 2
17 11 11 2 9 9 3 13 13 2 7 10 0 9 13 9 9 2
12 9 15 7 13 3 9 9 9 1 0 9 2
32 9 9 13 13 0 9 0 9 2 9 13 3 9 7 9 9 2 3 2 9 7 9 2 13 0 2 7 3 13 3 9 2
20 9 2 16 13 0 2 13 0 9 1 9 15 2 16 0 9 13 3 0 2
15 7 13 3 7 0 9 2 9 13 3 9 16 15 13 2
14 11 2 3 9 13 2 13 1 9 12 9 1 9 2
22 9 9 13 10 9 2 16 16 4 13 3 1 9 2 1 9 12 9 1 9 9 2
17 13 15 3 2 16 0 9 13 0 2 16 15 13 9 3 13 2
13 15 0 4 13 13 9 1 9 0 0 10 9 2
2 11 11
46 9 2 12 13 1 0 11 1 11 12 9 2 9 7 9 1 12 9 0 9 2 9 2 15 15 13 13 0 9 0 0 9 9 2 7 16 15 3 13 2 1 0 2 0 9 2
11 13 15 13 10 9 1 0 9 7 9 2
37 3 1 10 9 0 9 13 0 9 1 0 9 2 9 0 9 11 11 9 13 9 9 10 0 9 1 0 9 2 15 4 13 1 0 0 9 2
9 9 4 13 12 9 9 12 9 2
43 11 1 10 9 11 7 0 12 9 13 1 0 9 0 9 2 11 2 7 13 15 1 12 9 2 9 9 2 9 9 9 2 0 9 2 9 9 9 7 9 0 9 2
33 13 15 1 9 9 9 2 15 13 7 13 1 10 9 0 9 0 1 9 0 9 2 12 2 9 9 1 11 11 11 2 11 2
17 1 10 9 1 9 2 12 15 11 13 3 0 9 9 16 11 2
19 9 9 13 9 1 0 9 2 1 0 9 9 7 1 9 0 9 9 2
19 0 9 9 2 0 9 0 9 7 0 0 9 13 1 9 0 9 9 2
13 15 13 0 9 2 1 15 12 9 13 9 0 2
17 1 15 13 9 0 2 16 9 9 9 9 9 7 9 0 9 2
36 11 15 13 2 16 0 9 13 0 9 13 2 7 16 13 0 13 9 9 2 12 9 1 9 2 2 13 9 7 13 1 9 0 0 9 2
18 3 15 7 13 2 16 15 10 9 4 13 0 9 1 9 9 3 2
36 3 13 0 15 13 1 0 2 0 9 9 9 2 1 15 13 11 2 11 2 9 1 0 9 2 0 11 11 2 11 2 11 2 12 2 2
17 0 9 13 1 9 9 9 2 15 13 13 3 2 1 0 9 2
20 0 9 7 9 7 1 15 0 9 0 9 13 13 1 9 7 9 9 9 2
19 1 9 13 9 9 9 1 9 2 3 4 1 11 13 0 9 0 9 2
19 11 11 7 9 1 10 9 13 1 9 2 16 15 9 13 1 9 3 2
33 10 9 2 3 2 9 9 2 13 3 0 2 0 9 2 7 2 3 13 9 9 2 3 2 9 9 9 2 7 0 9 9 2
21 1 0 9 15 7 0 9 13 3 13 2 16 9 13 9 3 0 2 3 0 2
27 1 0 9 13 0 9 1 0 9 2 3 10 0 9 2 15 15 13 1 9 1 9 9 2 12 2 2
42 10 9 13 1 9 9 9 2 0 9 1 9 2 0 11 2 0 11 2 12 2 0 9 0 9 0 9 2 0 0 2 11 2 11 2 12 2 3 1 12 9 2
24 9 2 16 10 0 7 0 9 13 0 0 9 16 9 0 7 16 15 3 13 2 13 0 2
30 0 2 15 15 15 13 2 13 11 11 11 2 12 2 12 2 2 3 0 9 2 3 9 1 9 0 9 1 11 2
36 1 10 3 0 9 9 1 0 9 1 9 16 15 13 0 0 9 1 9 2 12 2 13 2 16 9 13 3 7 9 9 14 3 1 9 2
24 15 13 3 0 9 2 16 3 2 0 9 9 1 12 2 9 13 9 9 3 1 0 9 2
38 0 9 13 15 2 3 9 2 16 1 15 13 9 1 9 0 9 2 15 4 13 1 9 9 9 2 10 9 9 11 13 7 3 13 0 9 2 2
17 11 2 11 13 2 16 11 2 13 0 9 9 3 0 9 2 2
11 7 10 9 0 9 9 1 9 13 13 2
49 7 3 2 0 9 7 0 9 11 11 2 11 3 13 13 9 9 10 9 7 13 9 9 2 7 13 9 2 16 1 9 1 9 9 1 9 9 4 9 13 0 7 0 0 9 1 0 9 2
17 3 0 9 1 9 15 13 13 1 0 9 3 1 12 12 9 2
12 1 9 13 3 3 9 7 3 0 0 9 2
61 3 13 7 0 9 1 9 0 9 2 0 3 0 9 2 3 3 2 11 2 11 2 0 9 7 0 9 2 11 2 0 11 2 12 2 2 7 0 15 1 0 0 9 2 3 3 0 9 2 7 1 3 0 9 2 3 1 9 9 2 2
16 0 9 2 0 9 0 9 2 13 0 9 2 0 7 0 2
36 0 9 13 1 0 9 9 2 7 2 1 3 0 9 2 0 9 0 9 7 9 13 1 9 0 9 9 2 15 13 13 13 0 0 9 2
10 9 15 3 13 2 16 13 9 9 2
18 1 0 9 15 13 2 16 16 15 13 15 9 2 9 13 1 9 2
28 0 9 13 9 1 9 7 1 9 0 9 2 1 0 9 13 0 9 9 2 3 13 15 0 9 7 9 2
16 9 7 13 2 3 4 13 13 2 16 11 13 15 10 9 2
33 12 1 9 13 9 16 9 0 9 2 10 9 13 1 9 2 7 13 15 2 15 4 15 13 2 16 4 1 9 9 3 13 2
17 9 2 3 15 2 13 4 15 0 9 7 9 4 13 3 3 2
11 10 0 9 13 0 2 7 7 3 0 2
28 3 3 2 0 9 13 0 9 2 16 2 3 1 0 9 2 13 1 9 2 12 1 9 0 9 9 9 2
17 7 16 4 15 0 9 9 9 13 3 2 13 4 1 9 3 2
10 9 7 13 0 9 1 0 9 9 2
34 3 13 0 9 9 2 15 3 13 2 9 3 13 9 9 2 16 13 2 16 3 10 9 13 13 1 9 2 3 13 11 1 9 2
35 3 10 9 0 9 9 7 9 4 1 9 1 9 1 9 9 2 15 13 12 1 0 9 2 0 1 9 9 9 1 9 2 13 9 2
55 3 13 11 1 9 0 2 2 0 2 9 2 11 2 11 2 11 2 11 2 11 2 11 7 11 2 11 2 1 0 9 2 9 0 9 2 9 7 0 9 2 11 9 2 11 2 12 2 10 0 9 13 1 9 2
22 3 7 9 13 13 2 16 9 9 3 14 13 3 0 2 3 13 10 0 0 9 2
10 0 9 14 3 3 13 9 1 9 2
21 7 1 9 15 9 13 13 2 3 9 13 1 12 9 9 0 9 2 0 9 2
31 1 9 13 1 9 13 0 9 2 9 1 9 9 9 2 9 9 7 9 2 9 9 2 9 9 9 1 0 9 3 2
33 1 0 9 9 11 3 13 9 9 16 0 9 2 15 15 13 1 9 1 12 9 2 13 11 0 11 9 2 12 2 12 2 2
16 9 15 13 13 1 0 9 12 2 14 3 7 9 9 3 2
17 1 9 3 0 9 9 13 3 0 9 16 10 9 1 12 9 2
14 13 15 7 9 2 15 13 3 0 7 13 1 9 2
20 3 7 13 9 2 16 0 2 9 13 3 3 1 15 2 16 15 13 9 2
4 9 2 11 9
3 0 9 12
2 11 11
2 11 11
1 11
1 11
1 9
47 0 0 9 9 13 9 2 12 0 9 1 9 9 11 11 2 11 2 2 11 0 1 11 7 11 2 11 2 7 11 2 11 2 11 2 1 9 7 9 9 9 2 3 0 0 9 2
29 0 11 13 1 9 9 2 16 13 0 12 9 1 9 9 2 7 7 13 3 9 1 9 0 9 1 9 13 2
14 1 0 9 13 0 9 7 2 3 2 16 9 2 2
23 9 1 9 12 9 9 14 13 1 10 0 9 1 9 2 15 13 0 9 9 1 9 2
26 9 0 9 0 9 1 9 13 1 15 0 7 13 10 0 9 2 9 2 9 2 9 7 0 9 2
23 10 9 4 1 15 13 3 1 9 2 3 4 15 1 15 1 3 16 12 9 3 13 2
17 13 15 1 15 2 7 1 0 9 0 9 1 11 2 1 11 2
27 13 3 15 9 3 1 0 0 9 1 9 1 9 0 9 2 7 16 15 3 13 2 1 9 0 9 2
33 9 0 9 15 3 3 13 10 9 16 3 0 7 3 0 9 9 2 15 13 3 1 10 9 7 9 1 10 0 3 0 9 2
21 3 15 7 13 9 2 1 15 13 0 3 0 9 2 15 9 10 9 3 13 2
8 9 1 10 9 13 3 0 2
22 0 9 15 3 13 13 14 1 9 2 15 15 13 0 3 13 1 9 0 9 9 2
35 13 7 0 2 16 3 10 0 9 2 15 15 13 9 1 0 9 3 0 0 9 2 13 10 0 9 2 0 9 0 9 10 10 9 2
22 12 1 10 0 9 13 3 9 0 9 2 7 16 15 15 13 1 9 2 0 9 2
16 7 9 0 9 0 9 1 9 11 2 11 13 15 0 9 2
26 16 0 2 0 9 2 0 0 9 2 13 13 14 10 9 2 10 0 9 13 1 0 9 0 9 2
47 11 2 11 13 0 1 9 9 0 9 1 9 0 9 2 15 3 16 15 13 10 9 14 1 0 9 1 10 9 2 7 7 1 9 0 9 7 9 7 1 10 9 1 0 9 9 2
24 16 0 9 15 13 0 9 9 0 9 2 15 10 9 13 1 9 9 0 1 10 0 9 2
25 7 9 2 12 13 11 2 11 2 11 2 11 0 9 1 9 0 9 2 15 13 9 0 9 2
14 4 13 11 2 11 2 11 1 9 0 9 2 9 2
12 1 10 9 15 4 13 0 9 9 2 12 2
31 1 0 9 10 9 7 10 9 1 9 1 9 0 9 7 0 9 13 0 9 9 2 12 11 2 11 2 11 2 11 2
27 1 0 7 0 9 4 13 0 9 1 9 9 0 9 2 0 0 9 2 1 15 4 9 13 10 9 2
26 1 9 10 9 7 9 9 2 9 1 10 9 13 0 9 1 9 9 2 12 11 2 11 2 11 2
18 1 0 9 0 9 15 9 0 9 13 1 0 9 1 9 9 9 2
37 1 0 9 13 0 9 1 9 9 0 9 0 2 0 9 2 1 15 4 9 9 13 0 9 2 15 15 13 1 0 9 1 9 10 0 9 2
15 15 15 3 13 7 1 0 9 13 7 13 1 0 9 2
44 1 9 10 9 13 0 9 1 9 9 2 12 11 2 11 2 11 7 1 10 0 9 7 9 2 15 13 9 0 9 3 0 0 9 2 9 2 12 11 2 11 2 11 2
44 1 10 9 13 3 0 9 0 9 9 9 0 9 2 0 0 9 2 0 3 11 2 11 1 11 2 9 0 9 2 3 0 0 9 1 9 0 9 1 0 9 1 11 2
28 1 10 9 1 11 13 11 2 11 1 11 1 0 0 9 0 9 1 9 9 0 1 9 9 1 0 9 2
29 1 11 2 3 13 9 2 12 2 13 3 1 9 2 15 13 0 0 9 9 7 3 15 13 9 0 9 9 2
21 13 15 3 1 9 1 9 7 13 15 3 9 9 0 9 1 0 9 0 9 2
18 9 1 9 9 1 9 9 1 0 1 0 9 13 1 9 0 9 2
24 9 9 1 0 9 13 13 9 1 9 2 15 1 15 13 2 7 13 7 9 9 10 9 2
24 10 9 13 1 9 3 0 2 16 15 13 1 9 3 7 3 16 3 0 2 16 9 0 2
16 13 3 0 9 2 3 10 9 1 0 1 9 13 7 13 2
24 13 4 0 13 2 13 7 13 9 9 1 0 9 2 3 13 9 13 9 2 15 15 13 2
20 0 9 13 10 9 13 2 7 0 9 13 3 3 3 0 7 0 1 9 2
10 0 9 13 9 9 3 3 7 3 2
32 1 15 13 0 0 9 13 3 1 0 9 7 13 10 0 9 3 1 0 9 2 7 7 1 9 7 9 9 1 0 9 2
8 15 13 0 9 11 2 11 2
12 13 15 13 0 9 2 0 9 2 0 9 2
33 0 0 9 13 2 3 16 0 2 0 9 2 1 0 9 0 1 9 9 0 16 9 7 9 1 9 1 12 9 0 16 9 2
25 10 0 9 13 13 9 7 9 9 2 1 15 0 3 0 9 13 1 10 9 9 9 7 9 2
34 13 2 14 1 9 7 9 0 9 1 9 9 2 13 0 9 2 15 13 9 1 9 9 1 9 7 9 0 9 2 1 9 9 2
14 0 9 15 9 1 0 9 13 7 15 9 9 13 2
23 1 9 9 13 9 3 0 2 16 13 9 9 0 1 9 0 9 9 0 9 1 9 2
31 7 13 0 9 2 1 15 4 9 9 13 9 1 9 2 3 15 15 13 0 9 2 15 13 0 3 3 13 7 13 2
24 9 9 9 9 13 7 1 0 0 9 3 0 7 13 3 9 9 2 7 2 1 12 9 2
12 1 9 0 9 0 9 15 13 3 0 9 2
25 13 4 7 0 2 7 4 13 1 9 9 9 9 0 9 13 10 9 1 10 0 9 1 15 2
46 11 2 11 3 13 0 0 9 2 13 1 9 9 7 9 13 1 15 0 9 0 2 1 12 9 2 7 1 9 9 2 7 3 2 1 15 2 1 9 3 0 9 1 10 9 2
36 7 13 9 9 0 0 9 2 13 1 0 9 0 2 3 0 0 9 1 12 9 2 15 13 1 12 9 13 0 9 1 9 1 12 9 2
17 0 9 13 14 14 12 9 0 7 13 1 15 13 1 0 9 2
34 3 11 2 11 13 13 2 16 13 10 9 2 15 13 1 12 9 2 3 13 7 16 9 4 13 16 9 0 0 9 0 1 15 2
8 1 0 9 15 3 13 0 2
21 9 10 10 0 0 9 3 1 15 13 11 13 9 9 1 9 0 16 12 9 2
21 3 1 0 9 10 9 13 2 16 13 13 2 3 0 9 2 9 9 1 9 2
20 0 9 1 0 0 9 13 9 9 2 16 0 0 9 13 13 0 9 9 2
30 9 0 9 7 13 13 15 9 9 3 2 16 1 9 11 2 11 2 1 10 0 9 13 15 0 9 1 9 2 2
13 3 15 13 0 13 3 1 9 7 13 10 9 2
14 1 0 9 9 13 11 2 11 1 9 10 0 9 2
35 12 1 15 13 9 0 9 2 1 15 15 13 9 9 9 9 0 9 1 9 2 15 13 13 9 9 9 9 1 9 14 1 12 9 2
48 1 0 9 15 13 11 2 11 9 9 10 9 1 9 9 0 9 2 3 1 9 7 9 2 3 2 1 9 9 1 0 9 2 3 1 9 0 9 1 0 9 13 1 3 0 9 9 2
19 15 13 0 9 1 9 0 9 2 3 2 1 9 9 2 0 9 3 2
16 9 1 10 9 13 11 2 11 7 1 9 1 9 1 11 2
13 1 15 13 1 11 1 9 0 9 1 9 9 2
11 10 0 9 3 13 1 9 0 0 9 2
18 0 9 15 13 3 1 0 9 2 3 15 13 9 9 1 0 9 2
32 11 2 11 15 15 2 16 13 2 13 2 16 2 0 9 1 9 9 0 9 15 13 15 3 3 13 9 1 10 9 2 2
13 3 0 9 10 9 13 3 1 9 9 0 9 2
62 10 0 9 13 3 3 15 9 10 9 1 0 2 16 13 3 2 1 0 9 9 1 11 2 9 1 0 11 11 1 11 2 3 15 3 13 10 9 1 9 9 12 2 2 1 11 0 9 1 11 2 14 1 15 2 15 13 1 0 9 9 2
37 1 0 9 13 9 10 12 9 2 1 0 2 9 2 14 1 15 2 15 13 9 0 9 1 0 9 2 3 15 1 9 13 0 7 0 9 2
41 9 2 12 15 13 11 2 11 7 11 2 11 2 11 2 11 2 15 13 0 9 1 9 1 9 0 9 7 9 2 12 11 2 11 7 11 2 11 0 11 2
10 3 15 1 15 13 1 9 7 0 2
31 15 11 13 10 9 0 9 11 2 15 15 1 12 9 13 0 9 7 3 13 14 3 2 16 4 3 1 10 9 13 2
33 13 2 16 14 0 9 0 9 2 7 7 0 0 9 2 15 1 9 11 13 2 13 15 3 1 0 9 2 0 0 0 9 2
23 13 0 2 16 7 11 2 15 13 0 9 11 1 9 2 12 2 4 13 10 9 13 2
11 11 11 13 14 0 9 2 7 7 9 2
19 13 15 1 0 9 7 1 11 11 2 15 15 13 1 10 9 3 9 2
18 10 0 9 15 13 13 9 7 1 10 0 2 3 14 3 0 9 2
17 13 1 0 9 2 3 4 1 15 13 1 9 0 9 7 9 2
15 1 9 13 9 2 3 3 0 2 7 3 0 7 0 2
10 13 15 7 9 1 9 1 9 0 2
6 13 4 1 15 9 2
12 11 15 13 2 16 1 15 13 0 0 9 2
12 13 4 13 7 10 0 9 1 10 0 9 2
10 3 2 16 15 3 13 1 10 9 2
2 11 11
3 9 7 9
21 0 0 9 1 9 4 13 0 9 11 2 11 2 11 7 11 2 11 2 11 2
13 13 15 1 9 10 9 7 1 0 9 0 9 2
45 1 0 9 2 12 9 1 9 0 7 0 0 9 1 9 9 0 2 15 13 11 7 11 9 9 2 3 15 2 1 15 0 9 4 3 3 13 1 9 0 2 11 7 0 2
16 1 0 9 15 13 13 2 16 13 14 1 9 3 0 9 2
31 11 13 10 9 1 9 10 9 0 9 1 9 0 2 12 2 2 16 13 9 0 2 13 9 12 2 12 2 12 2 2
8 3 13 9 9 10 0 9 2
21 3 1 11 3 9 2 12 13 10 0 9 2 1 15 15 13 3 0 0 9 2
5 0 9 9 9 9
23 1 9 9 2 9 7 9 0 9 16 10 0 9 2 4 0 9 13 3 3 1 15 2
12 9 0 15 3 3 13 13 1 9 10 9 2
30 1 15 13 2 16 0 9 9 1 0 2 7 3 1 0 9 9 15 13 9 0 9 9 2 3 9 0 9 15 2
30 9 2 3 1 9 2 15 13 9 1 0 9 2 13 0 9 0 9 9 2 15 13 0 9 7 9 1 0 9 2
30 3 3 13 0 13 2 15 13 9 10 9 9 2 15 1 3 3 0 0 9 1 9 0 9 13 14 3 9 0 2
9 0 9 13 15 1 15 15 0 2
10 13 14 9 1 9 7 9 1 9 2
25 3 13 0 9 10 9 9 1 9 3 0 2 16 10 9 13 9 14 16 9 9 7 9 9 2
24 3 1 9 10 0 9 13 0 0 9 0 9 0 9 0 0 0 9 9 1 0 9 9 2
23 9 3 13 3 9 9 1 9 0 9 2 7 9 10 9 1 0 9 9 7 10 9 2
14 0 2 0 2 9 4 3 13 1 3 3 0 9 2
21 15 13 13 1 9 2 3 1 9 2 3 15 13 0 9 7 13 9 9 9 2
25 3 9 9 9 9 13 14 16 9 0 9 2 15 13 9 9 2 9 9 2 9 7 9 9 2
22 3 1 9 0 9 7 9 13 9 1 9 2 9 7 9 1 0 9 1 9 9 2
12 1 0 9 7 13 0 9 9 1 10 9 2
58 11 7 11 13 9 2 15 15 13 1 0 9 9 9 2 0 2 9 9 9 2 7 4 1 10 9 13 0 9 2 9 2 15 3 3 13 1 12 0 9 2 7 15 1 9 10 9 2 0 11 2 11 2 11 2 12 2 2
18 13 3 1 0 0 9 9 0 1 12 9 2 12 0 7 12 0 2
27 13 15 3 1 9 9 9 9 0 9 1 0 9 2 15 15 15 1 9 13 2 7 13 7 0 9 2
11 0 9 1 9 9 10 9 13 9 9 2
29 1 12 0 0 9 9 0 1 9 2 9 2 9 7 9 2 13 10 9 2 0 3 9 9 2 3 1 9 2
29 13 0 7 0 9 2 0 15 1 12 0 9 0 1 12 9 0 9 2 3 2 9 2 1 0 9 9 2 2
14 3 3 13 9 14 1 9 12 9 7 10 0 9 2
24 9 0 9 12 0 9 0 9 7 13 1 15 2 16 13 0 9 9 0 7 0 0 9 2
6 3 13 9 0 9 2
41 13 2 16 9 9 13 0 9 1 9 9 1 0 9 2 1 0 9 2 3 10 0 9 3 13 2 2 1 0 9 2 1 9 9 0 2 7 1 9 9 2
6 15 3 13 0 9 2
30 16 0 0 9 0 9 13 1 15 2 15 3 13 0 9 2 12 9 13 10 0 9 1 3 3 2 0 2 9 2
38 3 13 0 9 12 1 9 2 15 15 3 2 13 3 9 2 7 9 9 13 12 1 3 0 9 0 2 0 9 9 2 10 9 1 0 0 9 2
15 13 1 9 12 0 9 2 15 12 1 0 13 3 0 2
2 11 11
1 9
7 0 9 1 9 7 1 9
3 11 9 12
3 9 1 9
3 11 11 12
4 0 9 12 12
2 9 0
3 11 11 12
3 9 7 11
3 11 11 12
4 9 9 16 9
3 11 11 12
6 13 0 9 1 0 9
4 9 0 0 9
3 11 11 12
3 13 7 13
3 11 11 12
5 9 2 9 0 9
6 11 11 2 11 9 12
4 1 9 9 12
3 9 7 9
4 9 0 9 12
4 9 13 9 12
3 9 1 9
13 11 2 2 11 2 11 2 0 0 9 0 9 12
7 11 2 11 2 9 9 12
1 9
9 1 9 2 1 9 1 9 2 12
1 9
4 13 9 9 12
4 9 0 9 12
4 9 1 9 12
5 13 4 1 9 12
2 9 12
5 0 9 0 9 2
3 0 9 2
4 9 1 9 2
7 9 0 0 9 1 11 2
9 9 2 3 14 9 1 9 2 2
9 9 1 2 0 9 2 1 9 2
3 3 13 2
5 11 13 9 9 2
7 0 9 2 0 9 9 2
5 9 9 1 9 2
4 11 0 0 9
2 0 9
8 15 1 15 2 15 2 15 12
2 0 9
9 11 11 2 0 7 0 9 9 12
6 11 11 2 9 12 2
1 12
4 11 1 11 12
3 9 0 9
2 11 11
10 13 0 9 15 2 16 0 13 9 2
5 15 15 3 13 2
7 13 3 0 9 15 15 2
9 7 3 2 13 15 13 10 9 2
48 9 15 3 13 0 9 7 15 13 9 1 15 2 16 4 15 3 13 1 0 9 7 3 15 1 15 13 0 9 2 1 15 15 13 2 16 4 13 10 9 7 4 15 13 13 0 9 2
24 15 15 13 1 0 9 9 2 15 13 9 7 13 0 9 13 1 0 7 3 0 9 3 2
33 3 1 9 9 13 15 2 1 15 4 9 7 13 9 7 15 15 9 3 13 2 3 0 9 2 9 13 15 2 15 13 13 2
42 7 13 15 2 15 15 13 13 3 7 3 3 7 13 0 9 2 9 15 13 7 0 10 0 9 13 0 9 2 15 15 3 3 1 11 13 1 11 13 9 9 2
20 1 11 4 9 13 9 15 0 2 15 13 14 14 13 2 7 7 7 13 2
12 12 1 15 13 7 9 1 9 7 10 9 2
13 9 2 1 9 13 2 16 13 9 1 15 15 2
12 13 15 11 11 10 0 9 1 10 0 9 2
26 7 3 15 11 11 13 1 10 0 7 0 9 7 9 2 1 0 9 11 4 15 13 1 0 9 2
23 7 7 10 3 0 9 11 13 3 10 9 2 7 9 13 3 3 3 16 10 0 9 2
5 15 15 13 3 2
30 13 3 9 10 0 9 10 0 9 9 3 7 3 0 0 7 0 9 3 0 1 15 2 16 4 15 1 15 13 2
13 13 3 13 9 1 9 9 1 10 0 9 9 2
21 1 10 0 9 15 3 7 9 13 13 9 1 15 0 9 7 3 0 0 9 2
13 7 9 13 1 9 10 10 9 1 9 1 9 2
17 14 13 2 16 1 10 9 13 15 0 2 15 1 15 13 9 2
25 1 10 9 9 13 11 3 3 2 2 15 13 3 0 9 9 2 13 13 15 2 15 13 13 2
26 10 9 9 13 1 9 0 2 7 15 1 9 7 0 9 2 15 10 9 3 3 13 14 15 15 2
8 16 1 0 9 15 13 13 2
22 2 15 3 13 10 0 0 9 2 15 13 9 13 1 9 7 13 9 13 1 9 2
6 9 15 3 13 0 2
8 7 3 13 10 10 9 13 2
13 7 10 9 9 15 13 13 9 0 9 0 9 2
22 13 0 9 1 0 9 1 0 9 1 9 0 9 2 15 15 13 2 3 10 9 2
27 9 7 1 15 0 9 3 9 3 13 2 16 15 1 15 13 2 7 3 15 13 13 1 10 0 9 2
38 1 15 7 11 13 2 2 1 9 4 15 13 13 15 0 2 16 9 13 9 9 7 9 3 2 15 9 13 2 13 15 9 1 9 2 0 9 2
12 7 0 9 0 9 13 3 13 10 0 9 2
18 2 7 15 13 2 1 15 3 13 2 7 9 13 3 13 15 15 2
32 7 16 15 9 3 13 3 13 1 10 9 7 13 15 3 0 9 1 15 2 3 3 3 13 1 9 7 1 10 0 9 2
7 15 3 13 13 7 13 2
14 13 3 0 9 15 2 16 2 1 9 0 13 0 2
27 0 3 0 2 15 13 13 7 1 9 9 7 7 1 9 9 2 16 12 0 9 4 13 1 9 9 2
22 10 9 15 3 9 13 2 16 15 13 10 9 15 2 16 2 1 9 0 13 0 2
10 0 13 3 9 7 1 10 9 13 2
31 7 15 13 9 9 7 1 10 9 13 0 13 15 10 9 7 15 2 16 13 13 7 13 15 15 2 15 3 3 13 2
29 13 2 1 9 15 13 2 7 10 9 13 9 1 10 0 9 1 9 1 15 2 16 4 15 1 15 15 13 2
17 3 14 9 9 9 1 9 13 2 16 9 1 9 13 3 0 2
26 13 9 9 1 9 7 1 10 0 2 7 3 14 0 9 13 13 2 16 15 3 0 15 13 13 2
38 16 10 9 4 3 9 3 13 2 7 7 9 13 14 13 15 10 9 7 0 9 2 0 9 15 3 13 1 9 0 15 9 7 9 0 9 9 2
38 0 9 9 7 9 7 9 10 9 1 9 9 7 13 3 14 1 9 1 9 7 1 10 9 15 3 7 9 13 13 1 9 9 14 1 0 9 2
26 7 15 1 9 1 9 3 13 9 16 9 9 7 9 15 3 13 13 1 9 9 1 10 9 9 2
36 10 9 7 1 15 13 9 9 0 7 0 9 2 15 15 3 13 1 0 0 9 9 2 15 4 13 3 14 9 0 9 3 15 0 9 2
17 0 9 15 3 13 13 0 9 9 7 10 9 13 3 9 9 2
8 0 9 10 9 13 0 9 2
32 16 9 13 9 1 9 10 9 13 0 2 0 7 13 13 2 16 4 15 1 9 3 3 13 13 2 3 13 13 15 15 2
21 7 0 9 1 9 3 13 15 2 16 7 15 15 13 1 10 9 1 9 9 2
8 9 0 9 3 13 13 15 2
39 15 3 2 16 9 15 14 3 15 2 9 0 2 7 0 9 13 2 13 10 9 1 9 7 1 15 2 16 9 4 1 9 1 15 13 13 15 15 2
30 7 3 9 10 9 13 1 15 7 10 9 15 3 3 13 1 9 1 9 0 9 2 9 13 15 2 15 13 13 2
8 13 9 15 13 14 10 9 2
27 2 13 1 9 9 11 2 11 2 2 9 1 9 11 11 2 12 9 2 9 0 9 11 2 11 12 2
6 9 0 0 9 1 11
38 9 1 9 7 9 11 13 1 0 12 9 3 12 9 9 2 7 2 12 9 9 2 1 9 9 0 1 0 9 1 0 9 0 16 12 9 9 2
34 9 2 15 13 9 0 0 9 2 4 13 13 1 10 9 1 0 0 9 9 14 1 9 12 5 9 1 9 2 3 7 12 9 2
25 10 0 9 13 4 13 1 12 9 9 2 16 15 1 9 13 12 0 9 7 3 12 0 9 2
64 9 1 9 7 9 11 11 13 2 16 10 9 13 9 3 1 9 0 9 0 1 9 9 1 0 9 2 9 0 9 1 9 9 2 0 9 0 1 9 0 9 2 0 9 2 0 9 0 9 0 9 2 9 0 9 16 9 1 0 9 1 0 9 2
31 7 3 3 13 2 16 4 13 7 9 1 9 0 9 2 0 0 11 12 2 12 2 9 2 12 2 9 2 12 2 2
2 11 11
3 12 2 12
4 2 9 0 2
6 9 1 0 9 0 11
2 11 11
48 13 3 0 2 16 0 0 9 15 1 10 9 1 10 9 1 12 2 9 1 11 2 13 1 15 9 13 10 0 7 16 1 9 12 2 9 2 3 3 1 9 9 2 13 13 0 9 2
22 10 7 13 10 9 9 1 9 7 0 9 1 9 1 0 9 0 9 2 3 13 2
50 9 1 9 0 0 9 2 1 15 3 9 1 9 7 2 0 9 9 2 13 2 3 16 1 9 0 2 12 1 0 9 2 13 3 1 0 2 7 1 9 0 2 9 2 15 15 9 13 13 2
42 16 4 9 9 1 10 9 3 13 1 0 9 7 15 7 1 9 7 9 9 2 13 4 3 0 13 2 16 1 0 0 9 0 9 13 10 9 1 0 9 0 2
29 3 13 2 13 9 1 9 9 2 3 1 9 7 0 9 2 14 0 9 0 9 2 0 9 3 0 0 9 2
27 1 10 9 13 1 0 9 0 3 13 7 10 9 2 9 1 9 2 7 3 1 0 9 7 13 13 2
14 1 0 9 13 7 10 9 1 0 9 2 0 2 2
14 1 9 15 7 13 0 9 0 0 0 9 2 9 2
7 7 3 14 13 3 13 2
21 16 15 10 0 9 13 1 0 13 2 13 9 1 3 0 9 9 9 3 0 2
28 1 0 9 15 13 1 10 2 0 9 2 0 9 0 0 9 2 1 1 10 9 13 3 0 9 0 9 2
15 1 10 9 4 15 3 3 13 13 0 9 1 0 9 2
17 13 15 7 3 0 9 2 16 10 0 9 4 3 13 0 9 2
36 1 10 9 13 13 2 16 0 0 9 2 3 9 2 13 1 0 2 3 7 3 0 9 0 7 0 9 2 3 1 9 0 7 0 11 2
21 16 13 0 9 3 10 0 9 2 3 14 13 9 9 1 9 9 1 0 9 2
10 13 15 3 9 7 9 9 0 9 2
18 0 9 13 3 3 1 12 2 9 1 0 9 11 7 1 0 11 2
19 1 9 9 2 1 0 9 9 2 15 10 9 13 14 1 12 2 9 2
18 9 3 13 1 0 9 2 1 10 0 9 2 1 9 9 9 3 2
41 1 0 9 15 3 0 9 13 3 1 0 7 0 11 7 1 0 9 11 7 1 0 9 13 13 1 0 9 12 2 2 12 2 2 12 2 2 12 2 9 2
21 13 15 3 1 3 3 0 9 2 1 12 14 1 12 9 2 2 0 2 9 2
30 3 1 9 0 9 13 0 9 2 10 9 15 13 1 12 1 12 9 7 9 1 10 9 9 1 3 16 12 9 2
27 1 0 9 13 1 0 9 0 9 2 1 10 9 13 7 0 2 16 3 3 13 1 9 0 9 9 2
24 14 2 9 3 13 2 9 2 2 7 14 3 0 9 2 16 13 10 0 9 0 1 9 2
13 13 15 9 9 1 9 9 9 7 1 0 9 2
16 1 9 1 9 9 0 9 7 9 13 3 9 3 0 9 2
56 7 13 2 14 15 2 16 13 1 0 2 9 2 2 7 16 0 9 9 13 9 2 13 0 2 16 14 9 0 0 7 0 9 2 7 7 9 0 9 9 2 0 9 7 9 9 13 13 0 7 13 10 0 0 9 2
7 15 3 13 10 9 9 2
12 3 13 1 0 9 1 10 0 7 0 9 2
32 1 9 1 10 0 0 9 2 3 15 3 13 13 9 0 9 3 1 9 2 13 3 7 3 1 10 9 1 9 0 13 2
9 0 9 4 1 9 0 9 13 2
25 0 13 2 16 15 15 1 9 13 3 3 10 2 12 0 9 4 3 13 14 10 9 0 9 2
18 0 3 13 2 16 7 1 3 0 2 9 2 13 13 0 9 9 2
28 3 4 0 9 13 1 9 2 3 2 1 0 0 9 0 9 1 9 2 15 13 2 16 13 3 1 9 2
22 1 0 9 3 13 9 9 3 1 0 9 2 10 9 4 3 3 13 1 9 9 2
15 3 0 13 7 0 9 0 9 3 2 3 12 2 9 2
14 13 10 0 9 0 2 7 15 9 9 13 14 9 2
38 3 3 13 2 15 15 13 1 0 1 9 9 2 7 13 7 3 13 1 9 2 16 13 3 1 3 0 9 2 16 0 9 10 9 13 0 9 2
16 1 9 9 4 1 9 13 14 9 2 7 14 7 9 9 2
16 3 3 13 3 13 9 9 0 0 9 1 3 0 0 9 2
22 1 1 15 2 16 9 13 13 0 9 2 13 3 1 9 9 3 2 1 9 9 2
7 9 7 13 3 1 9 2
32 1 9 2 1 0 9 9 2 13 0 7 0 0 9 2 15 13 3 13 1 0 9 2 1 2 9 2 9 1 9 9 2
16 0 9 1 9 13 7 1 9 9 13 1 0 2 9 2 2
20 13 15 15 1 14 0 0 9 0 1 0 0 9 2 1 2 9 0 2 2
22 10 0 9 13 14 3 0 9 9 7 9 2 3 0 13 10 9 2 10 0 9 2
25 9 9 13 3 13 0 2 0 9 2 9 9 13 9 9 7 10 9 2 3 0 2 0 9 2
18 1 10 9 13 1 0 9 1 0 9 0 9 2 0 0 9 9 2
8 3 13 15 7 1 0 9 2
23 3 0 9 0 9 2 7 13 15 15 3 9 1 0 9 2 13 10 3 0 0 9 2
24 4 13 0 9 2 3 7 0 0 9 0 1 0 7 0 9 1 9 9 12 2 12 9 2
12 9 3 13 0 2 3 13 7 0 12 9 2
14 1 0 9 13 9 13 2 3 13 7 14 3 13 2
20 1 0 9 15 1 10 9 13 9 2 0 9 2 2 15 7 13 3 0 2
11 1 9 1 0 9 10 9 13 12 9 2
5 10 0 13 9 2
18 1 0 9 13 9 3 13 9 9 7 13 3 0 9 16 0 9 2
11 1 9 9 4 9 9 13 1 9 9 2
28 15 9 9 15 7 1 0 9 2 15 9 13 0 2 7 3 0 16 9 2 15 3 13 9 2 13 13 2
11 3 0 9 1 9 0 9 13 7 9 2
9 14 2 1 9 9 4 9 13 2
8 13 1 15 1 9 9 9 2
16 0 0 9 15 7 2 1 9 9 2 13 3 1 0 9 2
13 0 9 0 9 1 3 0 9 4 3 15 13 2
26 13 15 3 13 2 16 13 3 1 2 9 2 3 0 9 2 1 2 9 2 2 1 0 9 0 2
25 7 3 16 9 7 3 7 9 7 9 0 13 1 0 9 2 13 9 7 3 0 2 9 2 2
21 13 7 2 16 15 15 13 1 9 9 2 13 0 1 10 0 9 1 10 9 2
24 3 1 9 9 4 1 0 9 1 0 9 0 2 9 2 2 1 7 3 2 13 0 9 2
23 0 13 2 16 9 9 7 9 2 9 2 15 13 7 10 9 1 9 1 9 0 9 2
22 2 9 2 3 13 7 1 10 0 9 2 3 1 9 1 0 9 0 7 0 9 2
13 13 7 3 3 0 9 7 1 0 9 3 13 2
20 1 3 0 9 15 3 3 2 3 14 16 0 9 2 13 0 9 0 9 2
10 15 9 13 2 13 4 0 9 13 2
11 1 10 9 13 7 0 9 2 0 9 2
8 9 15 3 13 2 7 13 2
28 9 2 0 2 9 9 9 2 7 15 3 3 2 9 2 1 2 10 9 2 2 13 3 3 0 0 9 2
32 13 3 1 9 9 0 7 0 9 9 9 7 9 9 2 15 15 1 0 9 13 16 9 0 9 1 12 9 1 12 9 2
9 1 9 9 4 9 3 3 13 2
42 3 0 0 9 1 0 9 15 9 9 13 9 9 1 12 9 7 1 9 10 9 2 10 9 1 9 2 9 2 2 13 15 3 1 9 2 7 1 0 9 9 2
15 13 7 1 2 9 2 9 1 9 1 0 9 10 9 2
21 3 9 10 9 4 13 1 0 9 2 9 9 3 3 13 7 13 9 10 9 2
42 1 0 9 2 16 13 3 0 9 2 0 2 9 2 7 0 9 2 13 1 0 9 14 3 0 9 2 3 9 0 0 9 7 0 2 0 2 2 0 9 9 2
11 9 10 9 13 7 3 0 16 15 15 2
54 0 9 0 1 2 0 2 9 0 9 0 9 15 13 2 1 0 9 2 13 0 9 2 13 2 14 9 10 9 1 10 9 7 10 9 13 9 9 2 13 1 15 7 9 2 9 2 3 15 2 15 13 13 2
43 1 3 0 7 3 0 0 2 9 2 13 3 13 2 16 13 1 9 0 9 2 0 9 2 7 3 1 9 2 3 2 2 1 9 2 15 13 13 7 9 0 9 2
14 1 9 2 11 9 1 9 2 3 13 9 11 12 2
18 9 11 11 2 11 2 13 1 0 9 0 11 11 7 0 2 0 11
1 12
15 11 9 1 9 2 0 9 1 0 9 1 9 9 12 2
14 9 11 11 2 11 2 13 1 0 9 0 2 0 11
1 12
8 0 9 9 9 12 1 11 2
19 3 13 13 2 9 2 2 11 2 3 9 2 10 12 9 13 9 9 2
12 9 11 11 2 11 2 13 1 0 9 0 11
22 9 9 2 0 1 9 0 0 9 2 1 15 4 13 1 9 9 9 0 1 9 2
19 9 13 13 1 9 9 2 9 7 9 12 0 0 9 1 0 9 9 2
7 2 11 0 11 2 12 2
1 12
24 9 1 0 9 2 0 1 9 0 0 9 2 1 15 4 13 1 9 9 9 0 1 9 2
20 9 13 13 3 1 9 9 2 9 7 9 12 0 0 9 1 0 9 9 2
29 13 0 15 13 2 16 9 13 3 9 2 7 3 9 9 2 7 16 0 9 2 15 13 2 13 9 0 9 2
40 9 0 9 1 0 12 13 0 9 0 9 2 1 0 0 9 15 15 3 0 9 13 1 9 9 2 10 0 0 9 13 13 0 2 16 13 9 0 9 2
22 3 7 1 0 9 0 9 1 0 11 13 13 2 16 10 9 0 9 13 3 0 2
7 2 11 0 11 2 12 2
14 0 9 9 0 2 9 9 2 2 0 9 1 12 9
1 12
11 0 9 9 0 2 9 9 2 1 11 2
21 1 9 15 13 13 1 9 2 3 3 13 1 9 0 9 2 0 9 1 12 9
1 12
16 9 0 9 9 0 2 9 9 2 2 0 9 1 12 9 2
3 9 11 11
31 1 0 9 13 13 9 1 9 2 0 2 12 1 0 9 1 0 9 10 9 1 9 9 2 12 2 12 2 12 2 12
2 12 2
13 0 9 9 7 9 9 9 0 2 9 9 2 2
32 1 0 9 9 2 3 2 13 13 9 2 16 13 13 0 0 9 2 12 2 2 1 15 13 1 9 9 1 9 9 9 2
9 0 9 4 1 9 13 0 9 2
14 9 9 13 13 0 9 0 12 9 9 2 12 2 2
31 0 9 13 13 0 9 2 12 2 7 1 10 9 13 9 9 2 12 2 2 0 9 2 1 15 15 13 9 7 9 2
15 1 0 0 9 13 0 9 9 2 12 2 2 9 12 5
1 12
2 12 2
13 9 0 9 9 9 9 9 0 2 9 9 2 2
22 9 0 9 2 12 2 13 1 0 9 0 1 9 2 9 2 9 2 3 10 9 2
12 9 2 12 2 13 0 9 16 1 0 9 2
21 9 2 15 13 13 1 3 0 0 9 2 15 13 1 9 0 0 7 0 9 2
8 0 9 9 13 0 0 9 2
3 9 12 5
2 12 2
29 9 15 13 0 9 2 1 0 9 2 12 2 13 9 2 12 2 2 15 13 0 9 2 9 0 2 9 12 5
1 12
2 12 2
5 9 0 9 9 2
9 0 9 13 13 9 2 12 2 2
18 9 9 2 12 2 13 12 9 7 0 9 2 9 0 2 9 12 5
3 9 11 11
2 12 2
8 9 9 9 0 1 9 9 2
10 1 9 13 9 0 9 2 9 12 5
1 12
2 12 2
13 0 9 9 9 9 0 1 9 9 2 9 12 5
2 12 2
9 9 9 9 9 0 1 9 9 2
14 1 9 13 0 12 1 9 9 0 9 2 9 12 5
1 12
2 12 2
15 9 2 9 2 0 9 4 13 9 2 15 15 13 13 2
16 1 0 9 1 9 15 13 0 9 2 9 0 2 9 12 5
3 9 11 11
11 0 9 1 9 9 9 0 1 9 9 2
14 9 13 10 0 9 9 2 0 9 9 13 1 12 9
1 12
10 0 9 9 9 0 2 9 9 2 2
17 1 9 13 9 1 9 1 0 9 2 0 9 9 13 1 12 9
1 12
17 9 0 0 9 9 0 2 9 9 2 2 10 9 15 3 13 2
17 12 1 15 13 1 9 3 3 2 0 9 9 13 14 12 9 2
3 9 11 11
3 12 2 12
2 11 11
9 9 12 2 12 2 12 5 12 9
7 9 2 11 7 9 1 9
1 12
2 11 11
10 11 1 11 2 12 2 12 5 12 9
3 11 1 9
22 9 0 9 2 15 12 2 12 2 12 13 11 11 1 9 14 12 2 1 9 1 9
1 12
3 9 11 11
1 12
3 9 11 11
1 12
3 9 11 11
1 12
13 11 11 2 13 1 11 1 11 12 2 9 12 2
7 12 7 12 0 9 11 2
6 0 9 13 1 11 2
6 0 9 9 2 12 2
8 1 9 13 1 11 7 11 2
10 9 1 0 9 0 9 13 9 9 2
11 12 7 12 9 1 0 0 9 1 11 2
10 12 9 9 1 11 1 11 2 11 2
14 1 9 2 12 1 11 2 0 9 1 9 0 9 2
16 12 2 11 2 11 2 9 1 0 9 9 7 9 9 11 2
6 0 9 9 1 11 2
9 1 9 2 12 9 0 9 9 2
21 1 0 0 0 9 13 0 9 0 0 9 2 9 1 0 9 7 9 9 2 2
9 9 2 12 9 1 11 11 11 2
11 12 9 2 9 11 7 11 2 9 11 2
18 3 0 9 13 3 3 3 0 2 13 0 9 7 9 7 1 9 9
1 12
2 11 11
1 12
2 11 11
1 12
2 11 11
1 12
24 11 1 11 2 9 11 2 2 0 2 9 1 0 9 9 7 0 0 9 10 9 7 9 2
34 9 2 9 9 2 9 2 9 0 2 9 2 2 9 2 0 9 2 9 2 0 9 12 3 0 9 2 9 2 0 9 9 7 9
1 12
10 11 1 11 2 0 0 0 9 1 11
1 12
9 2 9 0 2 1 9 1 0 9
1 12
2 12 2
8 0 9 0 9 1 0 9 2
23 0 9 2 7 2 14 12 5 0 9 2 13 9 12 2 1 15 13 9 7 9 9 2
51 16 4 1 9 13 0 9 2 0 9 4 15 3 13 2 0 9 4 13 12 5 9 9 7 15 0 9 4 15 2 13 2 1 0 12 5 2 11 2 11 2 11 7 0 2 12 2 11 0 11 2
1 12
2 12 2
10 0 9 9 0 1 9 12 2 12 2
14 14 1 9 2 12 13 0 2 0 9 9 9 0 2
16 1 9 2 12 13 1 3 0 9 9 9 0 3 1 9 2
42 0 9 1 12 2 9 15 13 0 9 9 2 11 11 2 11 2 7 11 11 2 11 2 12 2 0 0 9 7 0 0 0 9 2 0 2 0 2 11 1 11 2
1 12
2 12 2
30 0 9 9 9 0 1 9 0 9 3 9 11 13 2 16 1 0 12 12 9 13 1 0 9 9 9 0 1 9 2
11 0 9 9 0 15 13 1 0 9 9 2
25 9 4 3 13 16 0 9 9 0 9 2 0 9 9 0 1 9 13 0 9 7 15 13 9 2
51 3 15 13 3 2 9 9 0 3 2 9 0 9 13 9 7 13 1 15 0 9 9 0 2 15 3 13 1 9 9 2 11 2 11 2 11 7 0 2 12 2 11 12 9 2 9 2 12 2 12 2
1 12
3 9 11 11
1 12
2 12 2
8 9 1 0 9 0 0 9 2
8 9 9 13 9 2 9 9 2
12 1 9 9 0 7 10 9 13 0 0 9 2
16 13 0 9 7 10 9 9 1 0 9 9 2 15 13 13 2
29 9 2 0 7 0 1 9 1 9 2 0 13 13 0 7 0 2 2 0 2 2 0 9 2 3 16 9 2 2
8 13 15 1 9 0 0 9 2
14 9 2 0 15 1 15 13 1 9 9 1 0 9 2
25 9 15 13 3 1 9 0 9 0 2 7 12 2 9 1 9 0 7 0 9 1 9 0 0 9
1 12
2 12 2
7 0 9 9 0 0 9 2
22 0 9 9 12 9 2 3 2 13 9 9 0 9 9 1 0 0 9 0 0 9 2
13 1 0 9 9 12 9 2 3 2 13 15 3 2
11 1 9 13 1 9 9 0 9 0 9 2
13 1 0 9 9 3 13 9 1 0 9 0 9 2
16 0 0 9 7 13 0 9 1 0 9 0 9 0 7 0 9
1 12
30 0 0 9 1 9 2 12 13 0 0 9 1 9 9 2 0 16 9 12 2 0 16 9 12 7 0 16 9 12 2
25 10 0 9 13 0 2 13 15 1 0 7 0 9 9 10 9 7 3 3 13 0 1 0 9 2
12 1 9 13 3 0 9 12 2 9 1 9 2
11 12 7 12 13 1 0 0 9 3 0 2
39 0 9 13 2 16 0 0 9 13 3 0 9 2 1 9 9 9 9 15 4 13 12 2 13 3 3 0 2 16 0 9 15 13 7 1 9 0 2 2
32 0 9 13 9 0 0 9 9 9 2 1 0 2 2 9 12 0 9 15 13 16 9 12 2 9 12 16 9 12 2 3 2
5 13 9 2 12 9
1 12
31 0 9 12 0 0 9 1 9 9 9 7 10 0 9 2 11 11 2 2 11 11 2 2 11 12 2 12 2 12 2 2
9 9 0 9 13 0 1 0 9 2
9 1 9 4 13 0 7 0 9 2
18 9 13 9 0 1 0 0 9 9 2 9 13 9 0 1 9 0 2
13 12 9 13 0 0 9 7 13 0 9 0 9 2
24 16 13 1 9 0 1 9 9 1 0 9 3 2 3 4 13 9 2 2 4 1 15 13 2
4 0 13 0 2
3 0 0 2
11 9 2 9 13 9 1 0 9 9 9 2
11 9 7 9 13 0 0 9 7 10 9 2
11 9 9 13 13 1 9 9 9 1 9 0
1 12
3 9 11 11
1 12
2 12 2
18 0 9 1 0 9 0 0 9 0 0 9 7 9 9 0 7 0 2
43 12 2 9 13 0 9 2 12 2 9 13 9 0 2 12 2 9 0 2 12 2 9 0 2 12 2 9 0 2 12 2 9 0 2 0 9 2 13 2 9 2 12 2
14 1 9 1 9 9 0 12 2 12 7 12 13 9 2
15 16 13 10 9 0 3 14 3 2 13 9 3 0 9 2
12 1 9 9 0 12 7 12 13 9 0 9 2
1 12
3 9 9 2
8 3 0 2 3 0 9 9 2
1 12
3 9 9 9
1 12
2 9 0
1 12
11 11 11 2 0 2 12 2 12 2 12 2
18 13 1 0 9 0 2 9 2 1 9 2 11 2 9 2 12 2 2
4 13 1 11 2
4 13 9 2 9
2 11 11
41 0 9 3 3 13 1 9 1 9 0 9 2 7 9 12 1 15 2 2 2 13 9 2 9 2 3 13 13 7 3 13 2 2 2 15 1 15 3 3 13 2
52 9 15 13 1 0 10 0 9 3 13 7 13 0 9 2 15 1 9 2 9 9 2 13 0 9 0 2 9 2 9 9 2 2 3 12 2 0 9 9 2 15 13 2 9 2 9 2 9 7 9 2 2
9 9 13 1 0 9 0 9 9 2
19 7 9 2 16 0 9 4 13 9 2 3 1 15 9 13 0 7 0 2
21 13 1 9 16 9 0 0 9 2 0 1 0 9 0 1 2 0 0 9 2 2
9 9 13 7 2 16 3 2 0 2
7 0 9 13 3 0 9 2
21 2 9 15 3 13 1 9 2 0 2 9 2 0 7 9 2 0 2 2 2 2
10 7 0 9 13 3 3 0 9 9 2
12 13 1 10 9 2 7 1 10 2 9 2 2
30 11 11 1 10 9 9 2 11 11 12 2 2 0 0 9 1 9 9 2 13 2 16 3 7 1 9 13 0 9 2
18 9 7 9 13 9 1 9 0 9 14 0 2 7 7 0 7 0 2
10 12 9 13 3 2 0 9 7 9 2
29 4 13 0 9 2 0 0 0 9 2 15 13 9 3 13 1 9 9 7 13 15 9 9 2 7 3 10 9 2
32 0 9 10 9 13 15 0 16 0 9 11 1 11 2 13 11 11 2 9 0 9 2 9 12 2 12 2 12 2 12 2 2
16 10 9 9 13 1 15 0 9 3 2 3 1 9 13 9 2
14 13 15 9 7 13 0 9 0 9 1 10 0 9 2
29 1 10 9 13 1 11 0 0 9 2 13 15 2 16 0 0 9 13 0 9 2 3 0 9 13 13 0 9 2
25 9 1 2 9 0 9 2 2 1 15 4 13 0 9 0 9 2 13 3 14 2 1 9 2 2
31 7 9 1 15 2 15 3 13 13 2 1 15 3 13 14 0 9 1 9 0 9 1 9 16 2 9 7 9 9 2 2
24 1 11 15 13 2 16 1 3 0 9 4 0 1 0 9 13 0 9 0 1 9 0 9 2
40 2 0 9 2 9 3 4 1 9 0 9 13 9 2 16 4 1 0 9 7 1 0 9 13 0 9 7 13 9 0 9 2 7 7 13 9 9 0 9 2
27 2 13 2 13 1 0 9 0 9 0 1 10 0 2 0 9 7 3 1 9 0 9 0 9 0 9 2
15 2 7 1 11 13 9 9 2 2 2 2 2 13 11 2
13 2 13 13 2 3 15 10 0 2 0 9 13 2
12 10 9 15 3 1 0 9 0 9 13 3 2
9 9 13 9 1 9 1 0 9 2
12 15 13 2 3 0 13 10 9 2 2 2 2
10 12 9 15 7 1 10 9 3 13 2
9 13 3 9 7 3 15 13 9 2
23 13 9 1 3 0 9 2 15 13 0 2 0 2 0 7 0 2 15 0 0 9 13 2
14 10 9 15 13 11 11 2 9 2 9 0 9 2 2
12 14 16 15 13 7 13 2 7 13 0 9 2
14 9 2 0 9 2 13 1 15 7 13 15 1 15 2
34 2 0 9 9 2 0 9 15 1 0 9 13 3 2 12 0 9 13 11 13 9 10 0 9 3 2 16 3 15 3 13 0 9 2
33 7 16 4 15 13 13 13 0 1 9 2 3 15 15 13 3 3 2 13 15 3 14 1 9 7 13 1 9 9 0 0 9 2
18 13 15 3 13 7 13 15 1 9 2 16 4 13 1 9 0 9 2
45 16 15 13 2 13 2 9 0 9 9 13 3 1 9 1 9 0 1 0 9 2 3 15 7 13 2 3 3 3 2 13 2 16 3 13 0 9 2 9 0 9 2 3 0 2
20 11 3 13 2 16 0 9 13 10 0 9 2 16 4 3 13 15 1 9 2
8 3 7 13 2 15 15 13 2
9 9 13 1 12 0 9 2 12 2
10 11 3 7 3 13 16 9 3 12 2
26 13 7 3 7 0 9 2 13 9 13 0 9 9 16 9 2 9 2 7 9 9 1 9 7 9 2
10 10 9 7 9 13 1 9 3 0 2
11 7 9 3 0 9 13 3 1 10 9 2
30 9 2 15 13 2 13 2 16 15 13 2 10 9 2 16 9 9 2 15 13 2 13 3 0 1 0 9 0 9 2
11 3 10 9 13 0 9 3 1 0 9 2
21 11 3 13 0 9 10 9 2 9 0 9 7 9 0 9 1 9 9 1 9 2
23 9 2 16 15 3 13 0 9 2 15 3 13 14 14 13 0 9 9 2 15 13 0 2
21 3 1 10 9 15 7 13 0 9 9 7 1 15 0 9 9 7 9 1 9 2
21 9 3 13 1 0 9 0 9 7 1 9 0 9 2 15 15 0 9 13 13 2
12 9 13 1 0 0 9 2 0 0 9 9 2
18 1 15 3 3 13 11 2 11 2 7 15 15 13 7 15 13 13 2
23 11 11 7 13 2 7 7 15 13 12 1 9 9 0 9 2 9 3 0 9 0 9 2
19 3 1 0 9 4 9 0 0 9 3 13 1 0 7 0 9 0 9 2
18 1 0 9 13 7 13 7 10 0 9 7 9 0 9 2 3 0 2
14 3 3 15 13 0 9 11 11 7 15 0 0 9 2
16 1 0 9 3 13 1 9 9 1 9 9 0 7 0 9 2
18 1 11 4 13 9 11 12 2 3 15 9 9 13 1 2 9 2 2
20 16 9 11 11 13 12 9 1 9 2 15 0 15 13 13 1 10 9 12 2
14 2 1 10 9 9 9 9 11 13 3 3 1 9 2
13 3 9 7 9 9 9 1 9 9 13 15 9 2
8 15 9 0 1 11 13 13 2
8 7 3 9 7 9 13 2 2
6 15 13 13 0 9 2
17 10 3 0 7 0 9 13 11 2 3 1 9 2 1 0 9 2
23 13 7 0 0 0 9 2 1 15 11 3 13 0 9 2 2 15 3 13 10 0 9 2
9 10 9 7 13 13 1 0 9 2
12 3 2 9 11 13 7 9 7 9 15 13 2
12 13 7 14 1 0 9 2 7 1 0 9 2
6 1 15 13 0 9 2
28 16 11 11 13 9 9 1 9 9 2 13 15 12 1 1 0 9 2 2 13 1 9 2 7 1 9 2 2
6 2 2 9 2 15 2
23 7 11 13 14 14 15 13 2 16 3 13 0 9 13 9 2 13 13 2 1 10 9 2
22 3 3 16 13 0 9 3 0 9 9 3 3 13 9 2 7 13 2 1 10 9 2
19 1 9 0 0 9 0 9 2 0 9 0 9 2 13 1 15 3 13 2
11 0 9 1 0 9 9 13 3 10 9 2
29 9 2 1 15 15 13 11 2 3 13 9 9 9 2 16 4 3 9 3 13 2 7 3 16 13 3 15 13 2
6 7 9 15 3 13 2
10 14 7 9 10 0 9 1 0 9 2
13 15 3 13 0 9 14 3 13 2 3 3 13 2
12 9 15 7 13 2 7 15 13 10 9 9 2
31 13 15 0 9 9 2 15 3 13 0 2 0 9 2 0 9 1 0 9 2 9 0 0 0 9 2 3 7 0 9 2
12 9 9 7 9 2 3 0 9 7 0 9 2
42 1 3 0 9 15 7 0 0 9 2 15 13 13 15 9 1 9 2 0 7 0 2 0 7 0 2 0 7 0 2 7 13 15 0 0 9 2 13 0 2 0 2
22 7 15 13 12 1 0 16 9 1 9 3 1 0 9 9 2 1 15 10 9 13 2
12 7 1 15 13 3 3 7 9 1 9 9 2
5 13 3 7 9 2
16 9 9 1 9 10 9 13 1 9 7 9 2 7 0 9 2
12 13 15 7 9 2 15 3 13 0 9 13 2
94 2 2 2 2 10 9 15 13 2 16 13 0 13 9 1 9 3 0 7 16 1 10 0 9 2 15 15 13 1 9 2 0 13 0 2 0 2 15 9 13 9 7 9 9 2 9 2 9 7 9 7 15 0 9 15 0 2 3 3 2 16 13 0 9 10 9 2 13 4 15 10 13 0 9 1 15 9 2 1 15 15 15 13 2 7 13 15 7 3 9 7 9 9 2
54 7 15 13 0 3 1 9 0 9 2 0 1 15 2 16 4 13 1 15 9 9 9 7 15 9 2 15 1 15 13 2 7 13 15 3 0 1 9 9 2 15 13 3 0 9 7 9 15 0 9 10 9 2 2
1 2
5 11 2 9 1 9
3 0 9 2
17 2 10 9 4 13 1 0 9 9 1 0 0 9 1 0 9 2
20 1 15 4 13 15 0 2 7 9 7 9 4 13 1 10 9 0 0 2 2
5 2 11 11 11 2
4 9 9 1 9
31 16 9 1 9 4 13 3 16 9 9 1 0 2 13 15 2 16 0 0 13 9 15 2 9 12 2 12 2 12 2 2
22 1 12 9 1 0 9 12 9 2 1 0 9 7 9 2 4 9 9 13 1 12 2
12 14 12 5 1 15 12 13 1 9 9 9 2
26 7 14 3 2 9 2 15 9 13 13 1 9 16 9 9 9 2 13 1 9 9 9 2 3 3 2
20 1 9 9 13 1 9 3 9 9 1 0 9 2 7 3 9 13 3 3 2
17 13 15 7 2 16 4 9 4 13 7 1 9 1 9 1 9 2
2 11 11
3 12 2 12
5 11 2 0 0 9
44 0 2 0 2 0 2 0 2 15 13 0 0 9 7 10 9 1 0 9 2 7 3 1 9 2 13 9 9 2 3 1 9 1 0 0 9 0 9 2 11 2 0 11 2
43 3 15 13 2 16 9 2 9 0 9 2 3 1 9 2 13 13 9 9 2 0 9 2 7 3 15 13 9 9 2 9 0 9 2 9 0 2 2 2 9 7 9 2
12 7 15 13 2 16 0 9 13 3 3 3 2
52 16 3 13 9 2 7 1 9 2 1 0 9 9 2 16 13 9 1 0 9 7 7 1 9 2 1 0 13 2 1 0 9 2 2 3 15 10 0 7 0 9 13 0 9 9 2 15 13 0 9 2 2
11 10 9 13 9 2 9 2 9 2 9 2
17 3 13 2 16 9 15 0 9 2 9 2 9 2 13 9 0 2
7 11 13 0 9 0 9 2
7 13 15 13 7 0 9 2
2 11 11
3 12 2 12
4 13 4 1 9
1 11
1 11
6 9 9 7 9 0 9
20 0 9 9 9 9 1 9 9 2 0 0 0 9 2 13 1 9 0 9 2
24 1 9 2 3 15 9 13 13 9 9 9 0 0 9 9 2 13 15 10 9 0 9 9 2
15 0 9 13 9 2 16 4 1 9 9 13 13 9 9 2
16 0 9 2 15 13 9 9 1 9 2 13 7 1 0 9 2
12 1 9 9 9 13 0 0 9 9 7 9 2
30 9 13 0 9 9 9 1 12 9 2 2 2 2 10 9 13 1 15 2 16 0 9 9 9 15 13 1 12 9 2
28 7 16 9 9 9 1 9 13 3 0 2 13 15 2 16 9 13 13 7 3 7 3 2 3 13 10 9 2
3 7 9 2
18 0 3 13 13 1 9 9 9 7 1 15 13 9 9 9 1 9 2
6 11 12 2 12 2 12
5 15 13 15 9 2
36 10 9 13 0 9 0 9 0 9 9 2 9 2 0 0 0 2 9 2 2 15 13 9 9 7 0 9 3 3 16 0 9 1 9 9 2
21 9 13 3 2 1 15 2 16 4 15 9 9 13 1 12 9 1 12 2 9 2
8 3 3 15 13 9 0 9 2
67 4 13 12 0 9 1 0 9 2 9 9 2 9 0 7 0 9 1 9 0 9 2 9 9 1 9 9 2 12 2 9 9 2 2 2 2 7 3 15 2 15 9 13 9 2 15 13 0 9 16 3 2 9 9 1 9 2 15 4 13 9 9 0 1 0 9 2
38 9 12 9 13 1 0 9 2 0 9 1 9 0 4 13 13 9 3 13 0 9 2 16 9 0 9 9 7 9 9 4 13 1 9 0 0 9 2
8 11 12 2 12 2 12 2 12
4 0 9 0 9
28 0 0 9 11 13 9 2 12 9 2 16 13 9 0 2 16 0 9 4 13 13 9 1 9 7 0 9 2
27 0 9 9 0 0 9 1 0 9 7 9 9 13 1 9 2 16 0 9 2 13 1 9 9 9 2 2
42 2 10 9 13 1 9 0 9 1 0 2 0 0 7 0 9 2 0 0 0 11 2 12 2 0 0 0 9 2 9 2 9 2 12 2 12 2 12 2 12 2 2
8 9 13 9 14 12 0 9 2
15 9 15 13 1 9 2 7 3 3 13 3 15 15 13 2
6 11 12 2 12 2 12
7 15 15 2 13 2 9 2
52 9 9 2 11 2 11 1 0 9 2 9 12 2 12 2 12 2 12 2 13 1 9 2 16 1 0 9 15 13 3 0 0 9 2 3 2 2 2 15 4 13 1 9 11 12 2 2 2 2 2 12 2
19 1 0 9 1 0 9 2 9 9 1 9 1 12 9 2 13 9 9 2
24 16 0 0 9 15 1 11 1 11 13 12 2 2 2 9 1 12 2 0 9 9 1 9 2
53 15 15 15 1 10 9 13 2 13 3 3 0 7 1 9 2 7 1 9 1 9 1 0 9 2 9 12 2 12 2 12 2 12 2 12 2 15 13 1 2 9 1 0 9 2 2 15 13 1 10 0 9 2
20 3 15 13 0 9 2 15 13 0 9 1 0 9 2 15 4 13 1 9 2
19 9 10 9 13 13 1 15 2 16 1 9 0 9 13 9 2 9 2 2
21 10 9 13 13 0 9 1 2 9 2 2 15 13 9 3 0 9 1 0 9 2
18 16 4 0 9 13 2 13 3 13 10 9 2 15 13 9 10 9 2
18 13 15 2 16 4 13 2 9 2 2 15 13 9 9 1 0 9 2
10 0 0 9 2 9 2 13 3 0 2
6 0 9 13 7 9 2
6 11 12 2 12 2 12
6 2 0 9 2 1 9
47 16 0 9 13 9 0 9 9 2 0 9 13 3 3 13 9 1 9 0 1 9 2 9 2 2 13 9 12 2 2 2 2 2 12 2 9 12 2 2 2 2 2 12 2 12 2 2
11 13 3 3 0 1 9 0 9 2 9 2
21 16 13 0 9 9 0 3 1 9 0 2 13 9 0 9 2 3 10 9 13 2
23 9 9 0 0 11 15 13 9 12 0 9 2 15 3 13 9 9 2 13 9 2 2 2
13 9 11 11 13 2 16 12 9 9 13 0 9 2
17 0 9 13 9 7 9 9 2 16 0 9 13 0 9 1 9 2
24 12 1 9 9 13 2 16 0 9 2 0 9 2 7 3 7 0 9 13 1 0 9 9 2
10 16 9 15 3 13 13 9 2 2 2
6 11 12 2 12 2 12
4 0 9 2 2
26 9 0 9 4 13 7 0 9 2 7 0 9 2 15 15 13 9 9 9 1 0 9 1 0 9 2
17 0 0 9 13 9 9 2 1 0 9 7 0 9 13 0 9 2
34 0 9 13 0 9 1 12 0 9 1 9 12 9 9 1 11 2 1 3 0 11 7 1 0 9 2 3 13 9 0 9 3 0 2
12 1 10 9 15 3 13 9 9 0 7 0 2
20 1 9 9 4 13 0 9 2 3 1 0 0 0 9 0 1 0 9 2 2
24 16 13 13 0 9 10 0 9 2 13 13 0 13 0 9 9 3 3 2 16 15 9 13 2
13 13 4 13 3 0 2 16 0 0 9 2 2 2
12 11 12 2 12 2 12 2 12 2 12 2 12
3 9 1 9
14 0 9 13 9 1 0 9 1 0 9 7 0 9 2
22 13 15 16 0 9 1 9 0 9 7 9 9 2 16 1 0 9 3 16 0 9 2
18 0 9 10 9 1 12 7 12 9 0 9 13 9 1 9 12 9 2
15 0 13 2 16 1 0 0 9 4 10 10 0 9 13 2
21 16 7 4 13 9 1 9 12 2 12 13 15 0 9 13 3 0 9 10 9 2
12 13 15 7 0 0 9 1 12 9 2 2 2
8 11 12 2 12 2 12 2 12
4 13 4 1 9
1 11
1 11
6 9 9 7 9 0 9
20 0 9 9 9 9 1 9 9 2 0 0 0 9 2 13 1 9 0 9 2
24 1 9 2 3 15 9 13 13 9 9 9 0 0 9 9 2 13 15 10 9 0 9 9 2
15 0 9 13 9 2 16 4 1 9 9 13 13 9 9 2
20 3 15 13 0 9 2 15 13 0 9 1 0 9 2 15 13 13 1 9 2
5 13 0 9 13 2
12 10 9 1 0 9 13 10 9 0 15 9 2
10 3 1 10 9 3 13 2 16 13 2
35 9 15 13 3 3 2 16 4 15 13 13 9 1 9 10 9 9 0 0 9 0 9 0 9 2 13 3 9 12 2 12 2 12 2 2
9 10 9 13 0 9 1 0 9 2
30 3 7 0 0 9 13 10 9 1 9 9 2 10 9 13 9 10 9 2 16 3 9 2 9 7 9 0 9 2 2
16 1 0 9 15 12 5 9 1 12 9 0 13 9 0 9 2
27 7 16 9 13 2 16 3 1 0 9 13 3 15 9 0 2 15 2 15 3 13 13 2 13 0 9 2
31 1 10 9 4 13 2 16 9 7 9 13 9 13 10 0 9 2 9 2 1 15 15 13 2 16 15 10 0 9 13 2
10 3 15 3 13 2 3 0 9 13 2
13 0 13 2 16 13 0 13 1 0 9 1 9 2
40 1 9 10 9 13 9 2 12 0 9 0 9 0 9 11 2 11 2 0 9 0 9 0 9 13 1 12 0 9 2 16 1 0 9 15 15 13 1 12 2
7 13 15 3 13 7 3 2
22 1 9 12 2 9 15 13 2 16 9 9 0 9 0 9 15 13 14 1 0 9 2
20 9 12 13 11 2 11 1 0 9 13 2 16 0 0 9 13 9 0 9 2
10 3 13 9 9 3 1 9 0 9 2
27 1 12 9 9 7 13 0 9 7 9 13 14 1 12 9 7 3 15 13 2 16 9 13 3 3 0 2
34 3 13 9 11 2 11 7 9 11 2 11 1 0 9 2 16 0 9 9 2 15 4 13 0 9 9 2 9 2 2 15 3 13 2
10 2 12 9 4 13 9 2 12 2 2
5 9 3 4 13 2
14 9 1 0 9 15 13 2 16 3 13 1 9 0 2
11 13 7 0 9 2 16 0 9 13 13 2
7 13 0 13 9 10 9 2
15 15 13 0 9 2 9 0 15 3 1 0 0 9 2 2
16 10 0 9 7 10 0 9 13 7 13 2 16 15 13 13 2
15 13 13 0 9 3 0 2 7 13 13 15 1 0 9 2
24 15 13 14 15 1 3 0 9 2 3 1 15 0 2 1 10 9 13 10 9 13 1 9 2
6 9 1 9 3 13 2
25 11 7 10 0 9 11 2 11 3 2 13 9 0 7 13 2 16 15 13 3 0 9 16 3 2
12 13 3 14 1 15 2 13 9 0 0 9 2
13 0 0 0 9 15 13 3 13 0 9 1 9 2
8 11 12 2 12 2 12 2 12
25 9 0 9 4 13 7 0 9 2 7 0 9 2 15 15 13 9 9 9 1 0 9 0 9 2
12 11 12 2 12 2 12 2 12 2 12 2 12
3 9 1 9
4 9 1 11 2
16 12 1 0 9 13 0 0 11 2 9 0 9 1 9 9 2
13 3 10 9 13 3 0 9 1 0 0 9 9 2
10 9 13 1 15 12 9 9 0 9 2
18 9 2 15 4 13 1 11 2 4 1 9 0 9 13 7 9 9 2
13 16 9 13 0 2 13 9 9 2 3 1 12 2
6 11 12 2 12 2 12
3 9 16 9
2 11 11
24 9 13 9 0 2 0 7 0 2 7 10 9 13 1 15 15 3 0 2 10 0 9 9 2
18 1 9 0 9 13 9 0 0 9 1 0 9 9 2 1 0 9 2
32 3 4 0 0 9 13 14 3 1 11 2 16 13 2 14 13 1 9 3 15 0 2 13 15 13 1 10 0 7 0 9 2
14 9 13 3 3 0 2 7 16 13 15 3 9 0 2
21 9 13 9 0 9 7 15 13 0 9 2 13 0 9 0 2 0 7 0 9 2
19 16 9 3 13 2 16 3 9 7 9 2 7 15 13 2 13 13 9 2
12 3 2 16 1 15 13 2 14 9 15 13 2
12 3 13 7 9 3 0 1 10 9 7 9 2
20 14 13 13 1 9 2 13 13 13 1 10 9 7 7 1 0 9 15 13 2
10 1 10 9 3 13 0 9 10 9 2
22 10 9 13 13 10 0 9 1 10 9 2 15 13 13 7 1 9 10 9 0 9 2
14 9 0 2 0 9 9 2 0 9 2 9 1 9 2
23 9 13 9 9 9 9 2 9 2 9 1 15 0 2 9 9 1 10 0 9 7 9 2
5 9 13 9 9 2
9 9 1 9 2 10 9 13 9 2
27 7 10 9 3 2 9 0 9 7 0 9 2 0 9 9 0 3 0 9 9 7 9 7 9 0 9 2
15 9 13 0 9 3 0 9 2 10 9 15 13 13 0 2
20 9 1 0 7 0 2 15 13 0 13 7 1 3 0 7 0 9 7 9 2
8 9 13 0 0 9 3 3 2
16 9 13 7 12 1 9 9 2 1 15 9 13 1 0 9 2
10 9 9 7 9 0 9 1 9 0 2
9 9 9 1 9 7 9 1 0 2
27 9 13 9 11 0 2 9 7 9 2 2 9 2 2 2 0 9 9 2 9 0 11 2 0 1 9 2
9 0 9 9 0 15 9 7 9 2
10 9 2 7 14 9 1 9 7 9 2
6 9 0 9 1 9 2
6 0 9 9 1 9 2
29 0 9 2 10 9 13 9 9 2 9 7 9 2 7 15 15 10 9 13 2 13 15 2 13 15 2 13 15 2
19 11 13 1 9 9 9 9 9 7 9 7 1 15 9 1 12 9 9 2
20 3 9 13 9 9 2 9 2 15 13 7 13 9 15 2 7 15 13 0 2
10 9 13 9 0 7 0 9 2 11 2
17 9 0 0 9 2 9 0 9 2 7 7 3 0 9 9 11 2
18 9 13 9 0 9 7 9 2 15 13 9 3 13 0 9 0 9 2
33 9 7 9 2 15 9 9 13 1 9 2 3 3 11 9 2 3 1 11 2 2 7 4 3 13 1 0 9 0 9 0 9 2
5 9 2 9 0 9
2 11 11
2 11 9
17 9 1 15 13 9 16 0 7 0 9 2 15 13 3 15 13 2
17 3 15 3 13 9 9 10 0 7 0 9 2 3 3 0 9 2
20 3 13 1 9 3 0 2 10 9 4 15 3 13 13 15 1 9 9 3 2
18 9 0 1 9 13 0 9 9 2 15 15 3 13 1 10 0 9 2
18 0 9 9 4 13 3 1 9 0 9 7 3 15 3 13 0 9 2
11 7 15 1 10 9 3 13 0 9 9 2
23 0 9 1 0 9 4 7 13 2 16 0 9 9 13 10 9 0 9 2 0 0 9 2
36 1 9 1 0 0 9 2 7 3 7 9 0 2 13 7 9 9 2 1 15 15 9 13 2 9 9 1 9 1 9 7 0 9 10 9 2
31 16 0 9 0 2 0 1 12 9 9 2 13 9 12 9 7 9 0 3 14 12 9 2 0 9 13 9 14 12 9 2
20 1 0 9 13 0 9 10 9 2 3 4 1 0 9 13 10 9 7 9 2
20 16 13 1 0 9 2 13 0 0 9 1 9 2 14 2 14 14 1 9 2
15 0 0 0 9 4 13 14 1 0 9 2 0 9 2 2
51 1 1 15 2 16 3 13 1 0 9 2 9 2 9 2 0 9 0 9 9 2 16 3 0 9 9 2 9 2 9 7 0 9 2 13 0 2 16 9 13 1 0 9 0 9 2 16 15 3 13 2
22 1 0 9 13 3 1 9 9 0 9 1 0 9 9 9 2 15 13 3 10 9 2
18 10 0 9 13 9 14 12 9 7 13 1 9 9 3 1 0 9 2
28 9 13 14 1 0 9 9 2 7 7 1 0 9 9 2 9 0 0 9 1 9 7 9 0 9 1 9 2
23 10 9 9 2 16 3 9 2 4 13 9 1 9 1 9 2 1 15 13 13 0 9 2
19 1 9 10 9 13 10 9 9 3 1 0 2 3 0 0 9 0 9 2
20 3 0 0 9 9 13 1 9 2 3 10 2 9 15 2 13 1 10 9 2
19 9 4 15 13 13 1 9 7 9 0 2 0 7 3 0 7 0 9 2
24 9 13 1 10 9 0 7 0 9 1 0 9 2 0 9 2 9 2 9 7 10 0 9 2
8 0 13 9 1 0 9 9 2
17 0 9 2 1 0 2 13 0 9 7 9 1 9 1 10 9 2
17 0 9 9 2 0 9 2 13 13 0 9 0 9 7 0 9 2
40 3 0 9 9 9 9 1 0 9 2 3 0 9 9 7 0 9 2 15 13 14 12 5 9 1 9 2 13 1 15 2 16 13 7 3 16 9 1 9 2
11 9 9 1 0 0 9 13 1 0 9 2
9 15 13 9 0 1 0 0 9 2
18 9 13 1 0 9 0 9 2 0 9 7 9 1 9 1 0 9 2
20 9 0 9 0 9 7 9 0 9 13 9 9 9 2 0 9 9 1 9 2
27 9 9 13 0 13 0 9 7 9 0 9 1 9 1 9 10 9 1 9 2 7 3 13 9 1 9 2
18 1 9 9 0 13 0 9 7 9 9 2 0 12 5 10 0 9 2
18 0 9 13 3 1 15 2 16 1 10 0 9 13 9 1 0 9 2
24 13 9 9 2 16 7 3 9 1 9 13 0 0 9 2 1 15 15 13 0 9 7 9 2
29 15 13 1 0 9 1 3 0 9 0 9 2 15 7 13 0 2 9 2 2 0 3 2 1 9 0 0 9 2
11 15 13 0 9 7 9 9 1 0 9 2
9 3 0 13 9 7 9 0 9 2
14 12 9 9 2 0 7 0 2 15 13 9 7 9 2
19 1 12 13 3 10 9 9 0 0 9 2 15 3 13 0 0 9 9 2
22 16 0 9 13 3 0 0 9 2 0 15 13 0 9 7 13 15 3 9 1 9 2
25 9 0 1 0 9 13 2 16 10 9 3 13 9 9 0 9 1 9 0 9 7 13 0 9 2
19 1 9 0 9 4 3 1 10 9 13 1 9 0 9 9 9 10 9 2
13 0 9 13 13 1 0 9 9 2 1 9 2 2
11 0 9 4 13 7 1 9 7 1 9 2
12 0 9 2 0 1 9 2 13 13 3 9 2
22 0 2 0 9 13 9 9 2 0 1 9 9 2 3 1 0 9 7 9 0 9 2
24 13 16 0 9 2 13 2 9 2 9 7 3 9 13 9 9 2 15 4 13 0 0 9 2
21 3 1 0 9 15 0 9 13 3 9 0 0 9 1 0 12 9 15 0 9 2
26 1 9 9 0 1 9 9 13 11 2 16 0 9 13 12 9 9 9 2 0 2 0 7 0 9 2
16 1 9 9 9 9 2 9 2 13 0 9 9 1 15 9 2
30 0 9 2 3 9 7 9 2 15 13 3 1 0 9 1 0 9 0 9 9 2 15 13 3 9 12 9 0 9 2
21 9 9 15 13 0 9 2 1 15 15 13 0 9 1 9 0 1 9 0 9 2
24 9 13 0 0 9 2 15 15 1 15 9 3 13 7 13 7 9 1 0 9 15 0 9 2
15 1 15 9 13 0 0 9 9 7 9 0 9 1 9 2
24 9 13 0 2 9 15 13 1 3 0 9 0 9 7 1 0 9 7 1 9 0 9 9 2
15 9 13 3 0 2 13 15 1 9 1 12 1 12 9 2
22 1 2 0 2 9 1 3 9 13 1 0 9 1 9 9 2 15 13 9 9 9 2
15 1 10 0 9 4 13 3 9 2 7 2 9 0 9 2
17 1 9 13 9 9 1 9 7 3 1 9 9 13 1 0 9 2
21 3 0 9 4 13 2 16 9 13 9 1 10 9 9 9 7 3 7 0 9 2
14 16 13 9 13 13 1 10 9 1 9 9 2 13 2
10 1 10 9 13 9 1 9 7 3 2
19 13 15 1 9 9 7 1 9 3 2 16 13 3 1 9 3 0 9 2
17 3 13 13 0 9 2 15 13 9 1 0 9 10 2 9 2 2
23 0 9 9 9 13 9 0 7 0 9 1 0 9 2 1 9 0 9 13 0 0 9 2
24 9 4 13 3 1 9 2 7 7 1 9 2 16 0 9 13 9 10 0 9 1 0 9 2
9 13 3 1 9 0 0 0 9 2
18 9 4 13 0 0 9 2 15 13 1 0 9 7 9 1 0 9 2
25 13 14 13 2 16 3 13 0 9 0 9 0 9 2 1 15 13 9 9 0 9 0 9 9 2
2 0 9
11 0 9 11 13 0 9 9 9 10 9 2
13 0 9 13 9 1 9 0 9 1 15 0 9 2
8 13 9 3 0 9 0 9 2
12 13 0 2 0 7 1 0 9 15 3 13 2
14 9 3 13 1 9 0 9 1 9 1 9 0 9 2
18 13 15 2 16 3 12 0 9 13 1 9 12 7 12 9 1 9 2
77 9 0 9 13 0 13 3 9 2 15 13 9 9 7 9 1 0 9 2 9 2 9 2 15 13 1 0 9 0 9 9 2 9 7 9 2 3 3 9 9 0 0 9 2 9 13 9 1 9 0 9 0 1 0 0 9 2 2 9 0 9 2 7 7 9 0 9 2 9 13 1 0 9 3 0 9 2
48 0 9 2 0 2 11 2 11 2 12 2 12 2 12 2 0 2 11 2 11 2 12 2 12 2 12 2 13 2 16 15 1 9 0 9 7 9 2 9 2 1 9 0 13 12 9 9 2
28 0 1 15 13 10 9 0 9 2 0 9 0 9 2 11 9 7 0 9 2 2 0 1 2 9 2 9 2
30 0 13 9 0 9 2 3 0 2 3 0 9 1 9 9 2 0 15 1 10 0 9 1 9 0 9 0 2 0 2
16 10 9 9 13 0 1 9 9 2 15 13 9 9 9 9 2
22 0 9 13 0 9 0 0 9 2 15 13 9 2 15 15 0 13 13 9 10 9 2
19 1 15 12 9 13 0 0 9 0 15 13 0 9 0 9 7 10 9 2
2 11 11
3 12 2 12
4 13 2 7 13
6 9 0 9 13 0 9
2 11 11
35 0 9 1 11 2 15 13 0 0 0 9 2 13 2 16 3 13 9 10 0 2 3 0 9 2 13 2 14 15 1 15 1 0 9 2
19 3 13 1 0 9 1 9 7 13 15 0 9 2 15 15 1 15 13 2
12 2 15 13 10 10 0 9 2 2 13 9 2
9 2 10 0 9 2 2 13 9 2
7 2 1 9 9 11 11 2
21 0 9 1 11 13 9 2 0 9 2 1 15 0 13 9 9 2 15 3 13 2
14 13 1 9 0 3 9 2 12 11 2 11 2 11 2
15 13 3 9 0 0 9 0 9 1 9 0 7 0 9 2
35 14 3 13 9 2 0 2 2 3 15 13 0 9 2 3 2 9 9 13 7 13 2 0 9 1 9 7 9 13 9 2 9 2 12 2
38 9 4 13 13 1 0 9 2 1 15 15 9 13 3 3 1 9 2 1 9 2 12 2 12 4 13 3 12 3 3 0 7 3 3 0 9 2 2
23 7 16 15 3 1 0 9 13 2 13 15 9 1 9 0 3 1 9 2 7 1 9 2
16 9 15 13 3 1 0 9 2 3 3 13 15 2 15 13 2
26 7 16 9 2 15 4 3 13 7 13 15 13 2 1 0 9 13 2 1 10 9 9 15 3 13 2
41 1 9 9 2 7 9 2 15 15 13 13 9 9 1 15 0 9 2 0 3 16 0 7 3 0 7 1 15 15 9 13 2 2 7 1 9 9 2 3 9 2
40 13 15 2 16 13 9 1 0 9 7 13 9 7 3 2 13 3 13 0 0 7 0 9 7 13 9 1 9 10 9 2 15 3 13 3 2 1 9 2 2
2 3 2
31 7 3 13 10 9 3 0 2 16 3 13 14 10 9 9 2 3 0 9 9 7 9 2 16 10 0 9 13 1 9 2
15 13 1 0 9 15 16 9 3 2 3 7 3 0 9 2
30 1 10 9 4 9 9 1 9 7 9 9 1 10 9 13 13 9 0 0 9 2 13 2 14 2 9 9 2 2 2
4 13 9 9 2
4 3 3 13 2
8 3 15 13 2 3 15 13 2
20 0 9 13 9 7 9 9 2 0 9 0 15 12 9 1 0 9 0 9 2
25 1 0 9 13 3 12 9 9 0 9 0 9 7 12 9 9 0 10 0 0 9 2 3 9 2
27 1 9 7 9 13 1 9 2 9 9 10 9 0 9 2 15 9 7 9 13 13 2 1 9 0 9 2
47 9 7 9 15 13 0 9 0 9 9 2 15 13 1 0 0 9 12 2 7 0 9 13 2 16 3 0 9 13 0 9 0 9 2 16 1 0 9 13 0 9 9 3 10 9 9 2
34 0 9 9 2 15 13 14 9 2 16 0 13 9 2 3 2 12 12 9 7 12 9 2 2 13 0 9 0 9 2 0 9 2 2
40 12 9 10 9 15 1 15 2 3 2 13 9 1 0 9 0 9 2 1 0 9 2 9 2 9 7 10 9 2 7 15 13 10 9 2 15 13 3 9 2
23 9 0 0 9 13 3 0 2 15 13 2 16 10 9 13 0 9 0 9 1 0 9 2
18 9 0 9 15 3 13 7 13 9 0 9 9 1 0 7 0 9 2
22 3 15 0 9 7 9 9 13 0 0 9 1 15 9 0 9 2 9 2 12 2 2
15 15 0 9 9 1 0 9 7 9 13 0 9 0 9 2
17 0 9 0 9 3 1 0 9 7 9 13 0 9 0 0 9 2
44 3 15 3 0 9 13 1 0 0 9 2 0 2 0 7 0 0 9 2 15 15 3 13 0 0 0 9 2 9 2 12 2 7 15 4 1 9 1 9 9 9 13 12 2
48 9 9 0 9 0 9 0 9 13 16 9 0 9 0 9 2 0 3 3 1 0 9 1 9 0 2 9 2 0 9 2 0 0 9 2 0 0 0 9 2 2 16 15 9 9 3 13 2
40 0 9 0 0 9 13 0 9 2 3 9 2 9 7 0 9 9 2 3 0 9 0 9 2 3 3 15 1 9 13 9 7 3 9 10 9 13 0 9 2
14 0 9 0 9 13 10 0 9 14 3 0 9 13 2
48 9 0 1 9 0 1 0 0 9 13 2 16 1 0 0 9 13 0 9 1 0 9 0 9 2 7 1 0 2 0 0 9 13 13 1 3 16 12 9 9 2 3 13 1 10 0 9 2
48 16 3 1 0 0 9 13 9 9 9 14 1 0 9 0 9 7 1 10 0 0 9 2 3 1 10 0 9 2 1 0 0 0 9 1 10 0 9 9 3 13 2 16 13 1 10 9 2
19 7 3 0 7 0 9 2 16 13 0 9 2 13 9 0 0 0 9 2
29 0 0 0 9 15 3 3 2 13 2 1 0 0 2 3 7 15 3 0 9 2 15 13 1 0 9 0 9 2
9 7 3 15 3 13 13 1 9 2
3 9 13 9
51 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 7 0 0 13 2 13 9 2 12 2 9 9 0 2 16 1 0 9 0 9 13 9 3 0 9 9 1 0 7 0 9 2
17 15 1 15 3 3 13 14 1 0 9 7 1 0 9 10 9 2
22 11 2 11 2 11 7 11 2 11 2 11 13 3 15 0 9 1 0 9 9 0 2
16 13 2 16 1 0 9 13 0 9 3 1 9 9 1 9 2
17 10 9 13 1 9 9 1 9 2 16 13 9 0 2 13 3 2
13 0 9 13 3 1 9 9 2 15 0 9 13 2
14 10 9 13 1 9 9 2 0 9 7 0 0 9 2
24 11 2 11 2 11 1 0 13 9 9 0 9 0 9 3 0 1 9 9 1 9 0 9 2
34 13 2 16 10 9 13 1 0 2 0 2 9 2 16 13 9 2 9 2 7 7 1 0 0 9 2 16 13 3 2 9 2 9 2
25 0 13 9 2 16 0 9 13 0 1 9 0 9 2 3 1 0 9 7 1 9 9 7 9 2
33 1 15 13 2 16 9 2 0 9 2 13 13 3 9 9 2 3 9 0 9 7 0 0 9 2 15 1 9 13 9 7 9 2
44 11 2 11 2 11 2 11 2 11 2 11 7 11 2 11 2 11 13 2 16 2 0 9 2 0 9 0 9 13 0 9 9 1 9 9 1 9 1 9 10 9 1 9 2
24 3 13 0 7 1 9 10 0 9 2 13 2 16 9 2 13 2 7 13 2 3 9 2 2
11 3 13 7 1 9 2 9 7 9 9 2
19 14 1 9 3 0 9 2 9 7 9 0 9 13 9 1 0 9 9 2
5 9 0 7 9 0
23 1 9 0 9 15 13 9 9 0 9 7 3 1 12 7 12 9 3 10 9 2 9 2
41 1 0 7 0 9 9 2 9 0 9 2 0 9 7 0 0 9 13 2 16 0 0 9 1 0 9 13 1 9 2 1 15 2 2 3 7 3 15 3 13 2
46 1 0 9 7 1 3 0 9 15 0 9 2 9 2 9 7 10 0 9 1 0 0 7 0 9 0 9 2 13 2 7 2 13 2 9 2 0 1 15 2 2 13 1 15 9 2
20 10 9 0 9 3 13 1 9 9 9 2 3 1 9 2 0 1 9 9 2
42 10 9 13 13 1 9 2 15 13 9 2 2 0 2 16 3 9 9 0 9 13 1 0 9 9 2 0 9 2 2 13 1 0 9 2 16 4 9 10 9 13 2
57 0 9 3 13 3 1 9 0 2 15 13 0 9 0 1 15 2 16 1 9 0 2 15 13 3 0 0 9 1 0 9 7 10 9 2 2 10 9 9 2 9 2 9 2 9 0 9 2 3 2 2 2 13 9 2 2 2
32 10 9 2 0 2 9 13 9 9 1 0 9 1 9 2 0 1 10 9 2 0 1 9 7 1 9 7 9 9 9 3 2
12 4 13 9 9 3 0 1 0 7 0 9 2
26 9 0 1 9 1 0 9 13 0 14 1 9 1 9 1 9 2 16 13 0 9 9 0 2 13 2
14 11 2 11 2 11 1 0 13 0 0 9 1 9 2
28 13 9 0 9 0 9 9 1 9 2 1 15 15 13 2 16 13 0 9 3 2 16 13 15 1 0 9 2
31 9 2 15 4 13 1 0 9 1 0 9 7 1 0 9 2 13 9 9 2 10 0 0 9 2 7 7 0 0 9 2
22 2 15 4 3 13 1 9 9 2 15 15 3 13 2 7 15 13 0 0 9 2 2
38 14 12 12 9 7 10 0 9 1 12 0 9 13 9 9 1 9 9 2 9 9 13 1 9 10 0 9 2 12 5 0 9 13 0 1 0 9 2
26 13 3 3 0 2 16 1 0 9 13 9 9 2 10 9 13 9 9 3 2 16 13 15 1 9 2
2 9 9
30 11 2 11 2 11 7 11 2 11 13 2 16 3 12 0 2 0 2 9 13 9 9 14 1 9 9 12 1 15 2
6 1 9 0 9 13 2
30 9 0 9 2 0 2 9 13 1 9 0 9 2 9 2 9 1 9 3 7 1 9 1 0 7 0 9 14 3 2
19 9 9 1 9 1 0 9 0 9 13 0 16 1 9 1 9 9 0 2
13 1 0 9 4 13 9 0 1 0 9 0 9 2
7 1 9 10 9 0 13 2
4 9 9 1 9
10 9 9 1 9 13 3 0 13 9 2
19 9 13 1 12 9 1 9 13 9 10 0 0 9 2 3 2 9 9 2
30 13 0 9 1 9 3 13 9 9 2 15 1 15 13 2 7 3 13 9 0 16 9 2 13 0 2 15 3 13 2
19 10 9 1 0 9 13 0 0 9 9 2 1 0 9 1 9 1 9 2
12 9 0 0 9 9 13 3 3 0 7 0 2
22 9 0 9 11 13 1 0 9 0 0 9 1 9 9 0 11 2 15 13 1 9 2
23 11 1 0 9 13 0 9 1 9 9 9 11 2 16 12 9 13 9 1 10 0 9 2
10 9 0 9 1 9 13 1 9 0 2
23 1 9 0 3 16 12 9 1 12 9 15 13 9 13 14 12 12 1 12 12 0 9 2
13 15 13 9 2 15 1 10 9 13 0 0 9 2
14 15 4 13 0 0 9 9 1 9 7 10 0 9 2
16 10 9 1 0 9 2 3 2 1 0 9 2 13 3 0 2
29 0 9 7 10 0 9 13 2 16 15 1 9 9 1 9 13 0 9 0 9 9 2 1 9 0 7 0 9 2
24 13 15 9 1 15 2 16 13 1 9 9 0 12 9 2 7 16 13 0 9 14 9 0 2
12 1 12 9 13 3 9 2 9 2 12 2 2
9 0 9 13 7 9 0 0 9 2
40 11 2 11 2 11 2 11 7 11 2 11 13 10 3 0 2 0 7 0 0 9 2 0 13 9 0 9 2 1 9 9 2 10 9 0 9 9 13 9 2
18 9 10 9 13 0 9 0 9 9 0 9 12 9 1 0 9 9 2
24 3 2 3 15 0 9 13 2 13 9 2 7 3 7 0 9 2 15 15 13 13 7 13 2
12 0 9 4 13 0 9 2 0 9 7 9 2
20 9 1 15 2 3 4 13 0 9 0 9 2 13 9 0 9 7 0 9 2
23 9 2 16 13 0 9 0 7 0 2 13 0 9 0 1 0 0 9 1 0 9 9 2
26 9 9 9 13 0 0 9 9 0 2 15 13 0 9 1 0 7 0 9 2 0 1 0 0 9 2
20 3 7 13 9 0 9 0 9 12 0 9 2 7 0 0 9 1 10 9 2
19 15 13 9 9 0 15 1 0 9 7 3 7 9 0 9 1 0 9 2
30 1 9 9 2 15 13 9 7 0 9 2 15 13 0 9 1 9 0 7 0 9 0 0 9 2 9 2 12 2 2
18 0 9 3 13 7 13 9 0 1 10 9 9 0 2 0 7 0 2
5 11 2 11 2 12
31 9 9 9 2 1 9 2 13 13 13 15 2 16 13 13 7 13 0 9 9 1 9 1 0 9 2 7 13 13 9 2
35 11 2 11 3 9 2 12 7 13 12 9 9 9 2 9 2 0 1 9 0 9 2 15 13 0 2 0 1 0 9 2 15 13 0 2
37 0 9 9 9 0 1 9 11 2 11 7 11 2 11 2 11 15 13 2 16 1 9 10 9 2 3 0 9 2 15 13 0 9 9 0 3 2
6 10 0 9 13 9 2
62 1 9 13 0 9 9 0 1 0 0 9 2 9 2 9 2 9 7 9 2 1 15 3 0 9 9 2 13 2 1 0 9 9 0 2 9 2 2 2 9 2 7 3 2 7 1 9 9 13 9 7 10 0 9 0 2 16 13 1 9 0 2
18 9 0 9 13 1 0 9 2 9 9 9 1 0 9 13 9 0 2
41 9 10 9 2 0 9 2 7 2 0 9 2 2 13 9 2 16 9 2 15 13 9 0 9 2 3 10 9 3 13 1 9 0 9 2 3 9 7 7 9 2
33 1 15 15 13 2 16 13 9 10 0 9 3 0 2 0 9 7 0 9 13 7 13 2 16 15 13 2 16 15 1 15 13 2
16 9 2 0 2 9 3 13 15 2 15 4 15 13 9 9 2
40 3 4 15 13 13 1 9 1 9 2 1 9 2 15 13 3 0 9 0 9 12 0 9 2 7 13 0 9 0 9 0 9 0 2 1 10 9 3 0 2
22 7 9 2 15 13 0 9 3 2 13 13 2 1 15 13 2 1 9 9 10 9 2
24 3 16 3 0 9 9 9 9 13 9 0 9 2 3 13 9 13 1 9 9 9 2 9 2
29 13 0 2 16 9 10 9 2 3 0 9 2 13 13 0 0 9 9 9 9 0 9 1 9 0 7 0 9 2
35 10 9 13 13 9 1 0 9 2 7 7 9 10 9 2 3 15 9 3 13 2 3 13 0 9 2 3 0 9 0 9 0 9 2 2
4 9 2 2 2
7 0 9 13 1 0 9 2
22 15 13 2 15 9 13 2 3 1 9 13 7 3 13 9 3 10 9 2 15 13 2
52 15 4 13 3 0 9 2 16 4 9 3 13 2 16 10 9 1 0 13 3 16 9 9 2 16 13 0 15 1 10 9 13 16 9 1 9 9 2 1 15 4 15 13 13 2 16 13 15 0 14 9 2
9 13 13 9 1 9 0 0 9 2
42 13 15 2 3 13 3 3 0 9 1 9 1 9 7 1 9 1 9 1 9 9 1 9 7 9 2 7 16 10 9 0 0 9 1 9 13 0 7 3 3 0 2
11 7 13 13 2 3 3 13 2 14 3 2
2 0 9
2 11 2
1 11
9 1 9 0 9 9 13 10 9 2
33 0 9 13 9 16 0 2 0 2 3 15 0 9 2 16 15 1 9 0 9 1 0 2 0 15 7 3 3 0 2 0 9 2
27 3 13 2 9 1 9 0 9 13 0 2 15 2 2 13 0 1 15 13 16 1 9 0 2 0 9 2
38 3 7 16 1 9 13 0 7 12 0 9 2 7 12 0 9 2 9 2 13 0 7 0 9 0 9 2 15 13 0 13 7 1 0 0 9 2 2
37 13 15 2 16 0 9 9 15 3 13 1 0 9 0 0 9 2 1 15 12 13 13 9 2 12 0 9 11 11 2 1 15 13 3 13 2 2
17 1 0 9 9 9 0 9 3 13 2 13 3 1 9 0 9 2
12 1 9 0 9 14 1 9 0 9 7 9 2
14 13 15 1 10 0 9 2 1 15 13 0 9 9 2
17 9 12 11 13 12 0 0 0 0 2 0 2 9 0 1 9 2
20 16 9 13 3 9 2 9 2 2 0 9 0 9 0 1 9 13 13 0 2
15 7 15 13 2 13 11 2 16 0 9 13 13 3 13 2
7 10 9 13 3 3 0 2
6 3 0 13 7 3 2
41 7 16 13 9 9 9 1 0 9 1 9 2 15 13 10 9 1 9 9 0 9 2 3 0 9 2 2 2 2 13 10 0 9 9 2 15 13 13 1 9 2
17 10 9 13 0 7 15 1 9 9 13 2 16 9 15 3 13 2
37 9 10 0 9 2 0 0 7 0 2 13 1 15 2 16 13 7 1 9 9 2 7 1 9 2 7 1 0 0 9 2 15 9 13 0 9 2
7 13 13 3 9 1 9 2
38 0 9 13 2 1 9 0 9 10 9 2 16 10 0 9 2 7 1 12 9 2 1 9 2 12 2 4 0 9 13 3 3 3 2 3 13 9 2
15 3 13 11 0 9 13 15 13 9 0 9 0 9 9 2
13 7 9 13 0 9 7 10 0 9 15 3 13 2
11 13 15 3 0 9 2 15 13 10 9 2
6 10 0 9 7 13 2
14 0 9 9 13 0 2 15 13 9 0 7 3 0 2
18 2 3 15 13 2 16 9 0 9 13 1 9 0 9 3 0 2 2
34 0 9 7 9 13 14 1 0 9 2 7 7 1 3 0 9 2 7 2 1 10 9 2 15 13 13 1 0 9 3 0 0 9 2
16 3 2 1 0 9 1 0 9 13 2 16 1 9 9 14 2
29 3 15 13 9 2 3 0 9 13 0 9 1 12 1 3 0 9 1 9 9 2 16 13 9 0 2 7 0 2
16 0 9 2 15 13 13 1 0 0 9 9 2 13 12 9 2
43 16 13 0 9 9 1 9 0 16 0 9 12 2 12 9 2 9 12 2 13 9 10 9 0 9 0 9 2 16 13 0 9 9 0 0 2 3 13 1 0 0 9 2
13 1 9 3 0 0 9 9 13 3 10 9 0 2
20 16 0 9 13 0 9 2 3 15 9 9 13 9 9 7 10 9 13 0 2
14 13 4 15 2 16 0 9 9 9 4 3 3 13 2
6 7 9 13 3 0 2
25 0 9 9 1 9 13 0 3 3 7 10 9 15 3 13 1 0 7 13 7 0 2 10 9 2
38 1 15 2 16 13 10 9 0 15 9 9 2 0 9 0 9 15 3 3 3 13 1 10 0 9 2 7 7 13 3 1 15 13 9 1 9 9 2
19 10 9 13 2 16 0 9 15 13 1 9 9 7 13 4 13 0 9 2
12 7 3 3 13 0 9 1 9 0 9 9 2
27 13 2 14 3 1 0 7 1 0 9 2 3 0 9 13 2 7 16 13 1 0 2 3 15 13 13 2
33 0 0 9 9 13 3 0 2 7 3 13 0 15 1 0 9 13 2 1 10 9 13 0 9 9 7 3 13 9 9 2 9 2
42 16 15 3 13 2 0 9 13 0 9 7 1 0 9 9 2 3 2 1 9 9 9 2 7 1 0 2 9 9 2 11 2 11 2 11 7 11 2 11 2 11 2
21 3 3 16 12 9 13 9 0 9 1 9 1 9 9 2 7 2 3 0 9 2
39 1 9 9 0 9 2 0 9 2 13 0 15 1 9 13 16 1 2 9 2 1 9 2 0 2 9 2 9 2 2 2 3 15 13 13 9 7 9 2
22 0 9 0 9 9 7 9 13 1 0 9 9 2 15 13 1 12 5 10 0 9 2
21 9 0 9 13 0 3 13 1 9 9 9 2 9 9 7 10 0 3 0 9 2
15 12 0 9 0 9 15 13 1 0 9 9 11 2 11 2
21 1 10 9 13 2 0 2 9 10 9 0 16 12 2 13 12 2 12 7 12 2
40 7 0 9 2 1 15 12 2 12 0 7 12 0 2 15 13 7 2 3 15 13 2 13 1 3 0 9 2 9 12 2 12 9 2 7 7 15 3 13 2
10 7 3 10 9 0 9 13 0 9 2
45 7 3 0 9 15 13 16 3 0 1 9 0 7 3 0 9 0 1 9 0 0 0 9 2 9 9 7 9 2 0 9 2 9 2 9 2 9 1 9 12 7 15 0 2 2
24 10 9 13 13 7 1 0 9 2 7 13 0 2 13 13 0 9 9 7 3 1 15 13 2
15 7 3 10 9 13 1 9 0 7 1 9 3 0 9 2
20 13 7 13 2 16 1 0 9 15 0 9 13 0 9 1 9 0 0 9 2
1 9
33 11 2 11 2 11 2 11 2 11 2 11 2 9 11 7 9 9 11 0 9 12 2 9 2 12 2 12 2 2 9 12 2 12
19 11 2 11 2 11 2 11 2 11 2 11 2 9 9 1 9 7 9 2
3 11 11 12
19 2 1 9 9 7 11 12 2 12 2 9 2 12 2 12 13 11 11 2
5 9 0 9 1 9
2 11 11
22 13 15 2 16 13 9 0 9 7 1 15 9 12 9 2 15 15 1 10 9 13 2
16 0 13 13 10 9 3 15 2 16 13 0 9 10 0 9 2
29 13 15 3 9 2 1 10 9 4 10 9 13 1 9 0 9 0 9 2 15 13 13 0 9 1 10 0 9 2
24 1 10 9 13 13 0 9 0 9 2 16 13 13 0 9 9 0 0 9 0 1 0 9 2
37 0 9 4 1 10 9 13 0 9 0 0 9 1 9 10 0 9 12 9 2 15 13 13 2 15 13 12 12 2 7 2 14 12 12 0 9 2
14 1 15 13 13 15 2 15 15 1 0 9 13 3 2
5 9 9 13 15 2
17 3 13 1 9 9 15 12 12 0 9 0 9 0 9 0 9 2
19 3 13 1 15 9 0 9 1 0 9 1 15 2 1 15 15 9 13 2
20 9 0 9 1 0 9 13 1 9 7 1 0 9 3 13 0 9 0 9 2
27 3 3 0 9 13 3 3 2 16 15 1 9 13 14 9 0 9 0 10 9 2 15 0 9 3 13 2
29 0 9 4 3 3 13 2 11 12 2 12 2 12 2 1 9 2 16 1 0 14 12 12 4 13 14 12 9 2
37 10 9 13 2 16 12 9 13 3 0 1 9 0 15 1 9 0 9 2 16 15 0 2 0 0 9 3 3 2 15 1 0 9 3 3 13 2
8 10 9 13 0 1 12 9 2
25 1 0 13 2 16 9 2 1 15 4 0 9 1 9 13 2 13 3 10 0 9 1 0 9 2
58 1 0 15 13 0 9 2 16 3 0 9 0 9 2 16 13 3 2 0 9 1 0 9 2 4 13 1 15 3 3 0 9 2 16 12 9 0 15 3 14 0 9 13 13 10 9 3 0 16 9 0 15 1 0 9 3 3 2
28 0 9 13 9 2 3 0 0 9 2 16 0 3 0 0 9 1 0 9 2 15 1 9 1 0 9 13 2
42 0 9 13 15 2 16 1 0 9 4 0 9 13 14 1 9 9 10 0 9 1 0 9 2 7 3 3 1 9 0 9 2 15 13 7 15 10 0 9 3 13 2
14 3 0 9 4 3 1 9 13 7 1 9 0 9 2
30 4 13 9 9 2 11 12 2 12 2 12 2 7 3 9 2 11 12 2 12 2 12 2 2 15 3 13 0 9 2
29 3 4 10 9 13 9 9 0 0 9 9 12 2 3 7 0 9 0 9 2 11 11 12 2 12 2 12 2 2
53 13 15 13 9 3 0 9 2 11 12 2 12 2 12 2 2 9 9 0 12 7 9 9 0 9 9 9 9 0 9 2 11 12 2 12 2 12 2 7 9 0 9 0 9 2 11 12 2 12 2 12 2 2
22 3 0 9 13 13 1 9 1 9 2 15 15 13 9 9 0 9 9 7 0 9 2
28 0 9 1 10 9 13 3 0 2 3 13 13 0 0 9 7 1 9 9 0 9 0 9 13 0 7 13 2
18 0 9 15 3 3 13 1 9 2 13 3 0 7 10 9 13 0 2
32 15 13 2 16 4 15 10 9 2 15 10 9 13 9 2 13 3 0 9 14 1 9 0 9 2 7 3 1 10 0 9 2
4 1 9 0 9
62 0 13 2 16 3 0 0 9 13 1 9 0 2 0 7 0 9 2 7 13 15 3 9 9 7 9 0 9 0 9 0 9 2 15 13 0 0 9 0 9 1 9 0 9 0 0 9 0 9 11 11 2 11 2 11 7 9 2 2 12 2 2
46 0 9 9 0 9 0 9 2 3 9 2 15 13 13 16 9 1 0 9 9 10 9 2 1 15 1 10 9 13 1 9 1 0 0 9 0 9 9 0 9 2 0 1 9 11 2
2 12 2
10 9 9 13 7 3 13 9 10 9 2
26 3 1 9 9 1 0 9 1 0 2 0 9 15 3 3 13 9 1 9 9 1 0 7 0 9 2
28 0 10 9 3 3 13 1 9 2 9 7 1 10 9 1 9 9 2 11 2 11 7 9 2 2 12 2 2
2 12 2
26 12 1 0 9 9 13 2 16 2 3 0 9 3 3 0 9 13 0 1 15 13 9 3 0 9 2
16 10 0 9 9 13 0 9 9 9 2 2 11 2 12 2 2
40 0 9 13 3 0 16 0 0 9 1 0 9 9 7 13 13 14 1 0 9 2 0 9 9 3 0 9 9 7 10 2 0 0 2 9 2 9 2 9 2
30 2 1 10 9 15 7 16 0 13 9 0 0 0 0 9 11 2 11 2 3 9 9 0 0 9 1 9 9 9 2
29 13 2 16 9 0 9 1 3 3 0 9 13 13 3 9 1 0 2 0 9 2 7 3 3 14 10 0 9 2
30 10 0 9 13 13 9 2 9 1 9 9 2 9 9 3 2 7 1 9 15 13 0 9 0 9 2 9 7 9 2
2 12 2
38 14 3 0 9 13 9 3 0 9 0 9 9 2 1 9 1 0 0 9 2 3 1 9 0 9 2 9 0 2 0 7 0 9 7 10 0 9 2
41 3 13 0 13 2 16 4 15 0 9 2 9 16 9 2 13 7 13 0 2 9 2 2 7 3 16 4 1 0 9 9 13 1 9 7 9 0 0 0 9 2
2 12 2
12 3 3 13 0 0 9 3 0 0 9 9 2
19 7 3 2 3 0 9 9 2 15 4 3 13 0 9 2 13 12 9 2
18 0 0 9 3 2 1 9 12 9 13 3 1 9 9 1 9 13 2
34 1 10 9 4 13 13 2 16 0 0 9 0 7 0 9 0 9 1 0 11 13 3 3 1 9 2 9 9 9 2 1 0 9 2
55 15 7 13 1 9 9 0 0 9 7 0 2 0 9 1 0 9 0 9 2 0 9 2 0 9 2 0 9 2 9 2 9 1 0 9 2 9 2 0 9 2 9 2 9 2 9 7 9 1 0 9 3 2 2 2
19 0 9 0 1 0 9 9 1 0 9 0 9 13 1 10 0 9 9 2
60 1 0 9 0 9 0 9 1 9 9 15 3 13 7 3 0 0 9 3 9 2 16 3 0 0 9 2 0 9 2 1 0 0 9 2 0 9 9 9 7 9 9 9 2 9 0 9 2 9 2 9 7 0 0 9 7 9 0 9 2
2 12 2
31 1 0 9 1 9 3 0 9 15 13 2 16 1 9 0 9 4 13 1 11 0 13 3 12 7 12 12 9 0 9 2
39 1 9 1 0 9 0 9 7 9 13 1 9 3 13 2 16 15 13 0 0 0 9 1 0 9 14 1 9 12 9 1 0 9 2 11 2 12 2 2
2 12 2
9 0 9 0 9 4 13 0 9 2
34 1 9 0 1 9 11 9 13 1 0 9 2 1 0 9 9 2 12 2 13 9 1 12 9 12 0 15 1 12 14 1 12 9 2
15 1 9 13 13 0 2 0 2 0 7 0 9 7 9 2
47 1 9 9 0 9 13 10 0 0 9 3 7 3 1 15 1 0 9 7 10 9 0 0 9 2 9 2 2 1 11 2 2 9 2 2 1 11 2 7 2 9 2 2 1 11 2 2
2 12 2
49 0 2 0 9 2 9 2 13 3 3 13 1 0 0 9 9 2 0 9 9 7 0 0 9 0 9 2 13 9 2 12 2 2 7 2 0 2 0 9 2 9 2 12 2 12 2 12 2 2
24 11 2 11 2 12 2 15 1 9 2 13 1 0 9 1 9 9 9 2 2 3 13 3 2
18 2 1 0 9 13 9 2 9 1 0 0 9 1 9 9 10 9 2
19 3 13 13 2 16 13 9 9 2 16 4 3 13 0 9 1 9 2 2
2 12 2
36 0 9 10 0 2 0 2 0 9 13 2 1 0 3 0 9 2 0 9 1 0 2 0 0 9 7 9 3 0 9 0 2 3 0 9 2
25 1 9 9 1 0 9 13 3 0 9 2 9 9 9 7 0 9 7 9 1 0 9 0 9 2
25 12 1 9 13 2 16 0 12 5 0 9 4 1 15 3 13 0 9 7 0 12 5 9 0 2
17 3 7 9 9 1 0 9 0 9 9 13 1 9 9 10 9 2
32 1 0 0 0 9 15 9 0 0 9 13 1 0 9 13 3 1 0 0 9 7 9 2 7 15 1 0 9 7 9 2 2
15 9 0 0 9 13 1 9 13 3 1 9 7 0 9 2
27 3 15 13 0 13 2 16 0 9 9 0 9 1 0 0 3 0 0 9 13 1 0 9 3 3 9 2
2 12 2
63 3 0 9 9 0 9 7 9 9 0 9 3 3 13 9 0 9 1 9 1 0 2 0 7 0 9 2 9 1 0 7 0 9 0 9 2 9 1 0 9 9 2 0 9 2 9 0 1 9 9 9 7 0 0 2 0 7 3 0 9 7 9 2
20 0 2 3 0 2 1 9 15 0 9 13 9 0 2 0 7 0 0 9 2
15 13 4 3 0 9 2 15 13 3 3 3 0 9 9 2
25 3 1 9 11 1 9 2 12 13 12 9 0 9 0 0 9 2 15 13 12 5 0 0 9 2
2 12 2
23 0 0 9 9 15 3 13 1 0 9 1 0 9 0 9 2 0 2 0 9 9 9 2
29 13 7 13 2 16 15 13 3 0 0 9 1 9 7 0 0 9 2 15 13 2 0 9 2 9 0 0 9 2
10 13 15 7 1 1 9 0 0 9 2
65 1 0 9 2 15 4 13 9 0 9 2 7 15 1 9 9 13 13 9 1 0 9 2 7 1 0 9 1 0 9 0 7 0 9 13 13 3 9 7 9 9 3 0 9 2 9 10 0 9 2 3 16 0 9 0 0 9 2 3 7 0 7 0 9 2
52 13 0 9 2 16 9 9 13 0 16 9 7 9 10 2 7 2 9 2 9 2 3 9 0 9 7 9 2 0 9 1 0 9 2 15 15 1 9 9 0 9 1 9 0 9 13 2 16 13 3 9 2
23 10 9 9 9 9 1 0 9 1 10 9 13 2 16 9 13 9 0 7 0 9 9 2
15 1 9 1 3 0 9 13 13 2 16 9 2 0 2 2
66 13 15 7 9 2 16 9 13 3 10 0 11 2 7 7 11 2 15 15 2 1 0 1 9 1 0 9 7 0 9 2 13 1 0 0 9 9 2 1 9 9 1 9 2 13 9 9 3 1 10 0 9 9 9 2 12 2 12 9 2 1 9 9 7 9 2
34 3 0 9 2 1 0 2 9 0 9 7 9 1 9 7 0 9 2 15 15 1 9 13 1 0 11 2 13 1 10 9 13 0 2
43 0 0 9 13 1 10 0 9 9 9 2 12 2 12 9 2 2 15 13 2 16 10 3 0 7 0 0 9 4 3 10 9 1 9 9 13 0 0 9 2 0 9 2
11 11 11 2 11 11 2 11 11 2 11 11
13 13 4 1 9 11 11 9 1 0 9 2 2 2
32 13 4 13 2 16 4 0 9 9 9 13 9 10 0 9 7 16 4 15 0 9 13 15 2 15 4 13 0 9 2 2 2
19 9 13 9 2 16 10 0 9 2 2 2 3 3 13 9 0 0 9 2
15 11 11 13 2 3 15 13 2 1 10 9 3 14 3 2
19 1 9 0 9 7 0 9 4 15 13 13 10 9 2 7 13 10 9 2
16 9 0 9 13 0 9 0 9 1 10 0 9 9 2 2 2
11 11 11 2 0 9 2 12 2 12 2 12
4 9 1 0 9
20 9 2 0 9 13 1 9 1 9 0 7 0 11 3 0 2 0 7 0 2
7 0 9 13 0 9 9 2
7 0 11 13 12 9 9 2
16 15 3 7 1 11 2 11 7 0 9 13 3 12 9 9 2
15 11 2 11 2 11 7 11 15 7 13 3 3 7 3 2
11 13 15 0 9 1 0 0 9 1 9 2
10 7 7 0 9 15 13 0 9 13 2
14 7 7 13 1 9 15 13 1 9 10 9 1 9 2
23 0 9 15 12 0 0 9 15 3 13 1 12 9 0 9 2 15 13 1 0 9 0 2
19 0 13 0 9 2 15 13 13 0 9 2 16 13 0 9 13 7 13 2
21 0 9 13 3 0 0 9 1 0 9 9 2 3 0 2 16 2 9 2 9 2
22 2 11 10 9 1 9 2 0 9 2 1 9 2 0 9 2 13 3 3 0 2 2
14 9 9 3 13 9 7 9 15 3 13 7 0 9 2
8 9 4 13 13 1 9 9 2
14 12 1 9 1 10 9 13 9 9 1 9 1 9 2
17 0 9 13 9 0 2 9 1 9 2 2 3 13 0 9 2 2
10 3 0 13 10 9 2 15 3 13 2
10 7 3 3 9 13 1 0 9 9 2
36 0 2 7 3 1 10 9 7 0 2 9 13 3 3 3 9 11 2 3 11 2 11 1 0 9 9 13 2 2 13 15 0 9 1 9 2
6 3 3 13 2 2 2
8 0 9 15 13 1 10 9 2
12 1 0 12 9 13 0 9 16 10 9 11 2
8 7 7 3 15 9 13 13 2
25 0 9 2 7 0 9 1 9 2 0 0 9 3 13 11 16 9 2 15 13 3 13 0 9 2
13 0 9 13 1 12 5 9 7 13 7 9 9 2
17 3 1 12 9 9 1 9 13 2 1 0 12 9 15 13 2 2
14 13 3 9 14 0 15 2 9 9 9 7 0 9 2
15 11 15 13 1 10 0 9 7 13 15 1 0 0 9 2
5 13 15 0 9 2
13 2 11 13 9 11 7 13 1 9 1 11 2 2
8 11 12 2 12 2 12 2 12
3 9 13 9
26 10 9 13 7 0 2 7 2 2 2 13 1 15 0 9 2 1 0 9 3 1 9 9 2 2 2
10 3 15 10 3 0 9 13 3 0 2
22 9 0 9 13 0 9 2 9 1 0 9 7 0 0 9 13 3 3 1 9 9 2
39 13 10 0 7 0 0 9 2 16 4 15 13 2 16 10 0 9 13 3 9 9 2 7 16 4 15 13 9 1 9 0 2 7 3 0 2 16 3 2
26 13 1 3 0 9 1 0 9 7 1 0 9 13 1 0 0 9 2 16 0 9 2 15 3 13 2
12 11 11 2 11 12 2 12 2 12 11 1 9
30 1 11 15 9 9 12 13 1 9 9 2 3 9 3 16 12 9 2 9 7 9 2 15 15 13 1 11 7 9 2
13 9 13 1 12 9 9 0 9 11 11 1 11 2
3 7 9 2
18 0 9 1 9 0 9 2 1 9 9 2 4 13 1 12 9 9 2
35 9 1 9 9 2 1 9 9 2 13 1 12 9 7 1 0 9 4 13 7 9 1 0 9 10 9 2 9 13 12 7 12 9 2 2
17 9 13 7 9 0 9 2 13 3 2 9 2 1 0 9 2 2
6 11 12 2 12 2 12
4 9 13 9 11
25 1 12 9 15 13 11 2 11 2 11 7 11 2 11 9 3 3 13 9 1 9 3 3 13 2
42 3 3 13 2 11 12 2 12 2 12 2 12 2 2 16 1 0 9 9 9 0 13 0 0 9 3 0 2 0 9 13 9 2 13 9 9 7 13 9 9 0 2
42 1 10 9 13 9 9 0 1 9 12 9 2 15 13 9 12 9 2 15 13 9 10 0 9 13 0 2 0 9 2 7 2 1 0 9 2 1 0 12 9 9 2
9 15 15 13 1 9 9 16 15 2
74 11 2 11 7 11 2 11 2 11 1 0 9 13 0 9 3 0 0 9 2 15 3 13 1 9 2 16 9 12 9 2 15 13 9 2 10 0 9 13 0 2 0 2 0 9 2 7 2 1 0 9 2 13 3 3 2 9 7 10 0 9 2 13 13 7 1 9 9 0 0 16 12 9 2
37 10 9 13 2 16 9 0 1 9 12 9 13 13 0 12 7 12 9 9 1 9 1 15 2 16 1 0 9 13 0 9 9 7 9 9 0 2
12 1 0 9 9 4 9 13 13 15 10 9 2
13 9 4 15 3 1 12 9 9 13 13 0 9 2
26 9 10 9 13 2 16 3 2 16 4 9 13 15 9 2 13 4 15 9 0 3 13 13 1 9 2
23 10 9 13 9 14 1 9 10 9 2 7 7 1 9 9 3 0 9 1 9 0 9 2
15 3 15 15 4 10 9 7 9 2 15 15 13 2 13 2
26 1 3 0 0 9 13 0 9 0 2 7 13 15 3 2 3 9 2 3 4 13 13 13 10 9 2
24 16 4 15 7 13 2 3 15 3 13 2 13 4 15 13 10 9 3 2 13 0 0 9 2
4 9 15 13 2
9 9 1 9 13 15 0 2 2 2
23 0 9 9 0 2 16 13 1 11 2 1 11 7 1 11 2 13 3 0 9 10 9 2
25 0 9 13 1 9 0 9 2 13 15 0 9 7 0 9 2 1 15 13 9 1 9 0 9 2
20 13 12 3 16 0 0 9 9 2 13 15 0 9 9 3 7 3 0 9 2
13 7 3 3 13 15 15 9 1 9 0 9 0 2
33 9 2 15 3 13 10 9 9 0 9 2 9 7 9 2 13 1 9 0 7 0 9 2 13 13 9 0 15 9 1 9 9 2
10 15 2 15 13 9 2 13 9 9 2
30 1 0 1 15 13 15 15 1 0 9 2 13 0 9 16 3 3 9 7 13 15 13 10 9 9 3 7 3 0 2
10 2 13 9 2 2 1 15 13 15 2
102 13 0 9 2 15 3 3 13 1 0 2 13 10 9 0 9 9 2 13 9 2 13 9 9 2 15 3 13 2 13 3 2 13 9 9 7 9 2 13 9 2 13 3 2 13 9 9 7 9 7 13 9 9 1 0 9 2 16 4 1 15 7 9 13 2 13 9 1 0 9 3 0 2 13 1 9 10 13 9 7 13 15 9 0 3 2 16 4 13 0 9 14 1 0 9 7 2 13 3 9 2 2
10 15 13 3 14 9 1 9 7 9 2
20 9 2 9 2 9 2 9 2 9 7 9 13 9 2 15 15 9 3 13 2
49 10 9 0 9 2 10 0 9 2 10 9 2 9 1 9 2 9 9 2 9 7 9 2 9 1 9 2 10 9 1 9 7 9 9 13 15 1 0 9 0 16 0 1 9 7 0 1 9 2
14 9 4 3 13 0 9 2 1 15 15 3 3 13 2
5 11 11 2 9 9
2 9 2
6 11 2 11 2 11 12
14 9 7 13 13 2 7 3 3 13 0 9 0 9 2
15 10 9 1 2 0 2 7 2 0 2 15 3 13 13 2
23 3 15 13 2 16 13 0 9 1 9 7 9 2 15 2 3 15 13 2 13 0 9 2
12 14 13 15 13 2 16 13 0 9 9 3 2
17 1 0 9 13 3 12 9 0 2 16 9 0 9 2 7 9 2
50 7 13 3 0 2 16 4 3 3 13 0 0 9 2 15 4 15 13 13 0 9 0 9 1 10 0 9 2 16 0 9 15 13 7 12 1 0 13 7 13 1 10 9 0 0 9 0 0 9 2
50 13 14 13 2 15 13 10 9 9 13 0 9 2 16 15 13 2 7 15 13 1 15 2 16 0 9 15 13 14 3 0 9 2 7 1 10 3 0 9 13 9 7 9 1 0 9 7 1 9 2
55 9 2 10 0 9 1 0 9 9 2 1 15 4 13 9 7 9 0 9 2 13 1 9 2 15 13 9 2 13 1 3 0 9 10 9 2 7 16 10 9 13 15 2 15 13 2 13 10 9 3 13 1 10 9 2
20 11 11 1 9 9 9 1 0 9 2 0 9 11 2 11 12 2 9 2 12
9 1 0 9 13 1 9 9 9 2
27 9 13 16 0 15 2 15 15 13 7 15 3 13 1 15 2 3 15 15 2 1 15 13 3 1 9 2
16 0 9 13 3 10 9 2 15 13 3 0 1 10 0 9 2
19 13 3 1 9 7 13 13 1 0 9 2 9 7 9 10 9 2 2 2
10 3 1 10 9 4 13 3 1 11 2
12 3 3 13 9 1 11 7 9 13 1 9 2
13 1 9 9 15 9 13 2 16 9 1 15 13 2
9 7 9 13 13 3 1 9 9 2
20 0 9 9 13 9 1 0 9 9 2 10 9 13 3 7 4 13 9 0 2
37 1 10 0 9 13 9 7 9 9 11 10 9 2 16 3 3 1 9 9 3 13 9 0 7 4 13 0 9 2 15 15 3 13 1 0 11 2
27 12 9 13 15 3 0 2 7 3 13 1 15 2 16 12 9 13 2 1 9 9 9 9 2 9 0 2
22 3 4 3 13 2 16 9 2 15 13 1 9 2 3 13 9 0 2 7 15 0 2
7 7 9 15 13 9 3 2
22 7 7 3 13 10 9 7 13 15 9 3 2 15 3 13 0 9 7 9 0 9 2
25 11 11 1 9 11 11 13 9 2 9 1 11 11 2 2 9 2 11 12 2 9 2 12 2 12
12 7 9 1 9 4 3 1 0 9 13 3 2
73 0 9 9 15 13 9 2 3 3 10 9 2 15 13 1 9 0 2 0 2 0 7 0 9 2 13 3 3 0 1 9 7 9 0 9 1 9 2 9 2 9 7 9 2 16 10 9 13 0 9 1 9 2 15 13 1 9 2 1 3 0 9 2 7 1 0 9 9 3 13 1 9 2
20 11 11 1 9 9 9 1 0 9 2 0 9 11 2 11 12 2 9 2 12
2 0 9
2 11 2
1 11
9 1 9 0 9 9 13 10 9 2
18 9 1 9 7 9 9 1 9 1 9 13 3 11 12 9 1 11 2
30 7 7 1 0 9 15 13 1 0 9 9 7 9 7 3 15 9 10 9 13 3 2 11 12 2 12 2 12 2 2
39 7 16 9 7 0 9 13 1 9 3 3 10 0 9 2 13 1 15 9 2 2 9 13 0 2 16 3 13 0 9 1 9 2 1 15 15 9 13 2
17 7 10 9 2 1 10 9 7 1 10 9 2 13 3 9 9 2
15 3 0 9 9 1 0 15 0 9 15 3 3 13 13 2
2 11 11
1 9
10 14 9 2 7 7 9 13 10 9 2
35 1 0 9 15 13 1 15 2 16 10 9 15 13 0 2 13 15 2 3 1 9 0 2 2 7 0 3 13 2 3 2 13 1 9 2
16 7 13 15 13 3 14 9 3 0 1 0 9 0 7 0 2
14 1 10 0 7 0 9 15 1 0 9 13 9 9 2
28 2 1 1 10 0 9 2 3 1 0 7 0 9 2 13 4 15 3 13 1 2 9 2 2 3 9 2 2
53 13 3 1 9 0 9 2 13 14 1 9 13 2 13 0 9 2 2 7 1 0 9 2 3 0 2 3 2 0 13 3 3 2 3 2 15 13 3 1 11 2 7 15 1 9 2 9 7 9 0 9 2 2
17 2 10 9 3 13 2 15 13 0 10 0 9 1 9 13 2 2
26 1 10 9 13 9 9 7 3 2 3 1 0 0 9 15 3 13 1 9 0 0 9 3 2 2 2
66 7 10 9 15 3 13 7 1 9 0 2 1 9 10 0 9 2 3 3 9 1 9 0 7 0 2 13 7 13 3 2 16 1 9 0 9 13 9 1 9 2 3 2 16 13 1 0 9 2 3 13 2 13 13 9 2 7 2 9 7 9 2 7 0 9 2
31 7 9 9 15 13 7 1 0 9 16 2 10 9 0 9 13 9 2 7 2 0 9 10 9 15 3 13 1 9 2 2
32 10 9 13 1 15 14 3 1 15 2 16 9 9 0 9 13 1 0 9 2 7 15 9 3 13 2 13 1 10 0 9 2
51 13 4 13 2 16 3 13 3 0 7 0 9 1 10 0 9 2 9 9 7 9 7 2 0 9 2 2 7 1 1 9 9 9 2 3 1 15 3 13 1 9 11 2 11 2 3 10 9 13 2 2
20 3 0 9 13 10 9 2 2 0 9 15 3 13 16 2 0 9 2 2 2
39 10 9 13 9 9 1 2 9 2 13 2 16 15 3 13 7 13 3 15 3 13 2 7 2 2 9 2 2 3 13 15 13 7 1 9 0 9 2 2
37 14 0 9 2 1 0 9 2 15 3 13 1 9 10 2 1 15 3 3 0 2 9 9 2 7 13 1 2 2 9 2 7 2 2 9 2 2
37 3 15 13 2 16 1 9 1 10 9 2 16 3 2 0 2 9 2 0 2 0 2 7 3 9 2 0 2 13 7 13 3 3 2 9 2 2
22 1 9 15 3 13 3 3 9 13 9 2 2 9 2 2 16 2 2 9 2 2 2
20 13 15 14 2 16 4 13 3 13 7 0 9 9 2 2 3 2 9 2 2
19 15 7 3 13 9 1 15 2 16 3 13 1 9 9 2 7 9 9 2
18 13 7 0 3 13 2 16 1 0 9 9 13 7 9 0 2 9 2
21 9 1 15 15 7 13 3 1 12 2 9 2 1 0 13 12 9 9 3 0 2
16 9 9 15 13 3 16 9 0 1 9 2 9 2 9 2 2
12 15 15 13 9 2 3 10 0 9 10 9 2
8 9 7 9 13 3 3 10 2
23 3 13 15 9 9 0 0 9 9 2 15 13 9 15 2 9 0 0 9 2 3 9 2
26 3 7 10 0 3 0 9 2 16 3 2 0 2 9 2 9 2 9 1 9 2 13 1 10 9 2
26 10 0 9 3 13 3 7 0 9 2 0 9 10 0 9 7 3 3 7 9 0 9 2 3 9 2
9 7 3 3 15 1 9 9 13 2
30 3 1 15 4 7 3 13 13 1 9 3 3 0 9 9 2 9 7 10 0 9 2 3 15 13 7 1 0 9 2
5 1 9 9 1 11
2 11 11
2 11 11
15 15 0 9 13 1 10 0 9 9 9 1 9 15 9 2
17 1 9 0 9 9 13 0 9 1 10 9 7 9 1 0 9 2
24 9 0 9 1 9 9 13 0 9 0 0 9 2 11 2 2 9 1 15 1 9 12 2 2
29 10 9 13 2 16 4 15 9 1 9 13 1 9 12 10 9 9 2 15 4 15 13 13 3 7 3 0 9 2
17 9 10 9 0 13 0 9 2 15 3 13 9 9 1 0 9 2
65 9 13 13 1 12 0 9 2 3 2 9 0 9 9 1 9 1 12 9 3 1 12 9 2 9 9 1 9 0 12 9 2 3 9 9 1 9 0 9 7 9 3 1 12 5 7 12 5 2 7 9 9 9 0 9 1 9 7 3 9 3 1 12 5 2
14 9 0 2 3 2 0 9 15 13 13 3 10 9 2
59 12 1 9 1 10 9 2 7 7 1 9 1 9 0 3 0 9 0 14 1 9 2 7 3 1 9 0 9 1 9 9 0 9 2 13 3 0 9 0 9 7 9 9 11 2 12 2 0 9 11 11 2 0 9 1 0 9 2 2
32 1 10 9 2 0 9 9 2 4 9 9 13 14 0 9 0 9 9 11 2 7 3 10 0 9 2 0 1 0 9 11 2
28 10 9 15 7 13 1 9 13 0 0 9 1 0 9 1 0 9 7 1 0 9 1 0 9 9 1 11 2
64 10 0 9 3 13 1 9 3 1 9 0 2 11 11 2 2 0 9 9 1 11 2 9 12 2 12 2 12 2 11 11 2 2 11 11 2 2 9 7 0 9 2 9 12 2 12 2 12 2 7 13 15 1 9 1 0 9 1 9 9 7 1 9 2
1 9
32 0 9 1 9 13 1 11 13 1 9 9 1 0 1 9 2 15 13 0 0 9 2 1 15 0 9 9 1 0 3 13 2
28 9 9 1 9 9 1 9 9 4 13 1 9 12 2 12 9 0 9 2 1 9 4 13 0 0 9 11 2
19 1 1 9 9 9 9 1 11 13 9 3 13 9 0 9 1 9 9 2
42 1 9 1 9 9 4 13 0 12 9 10 9 2 9 0 9 2 9 12 2 2 9 2 9 12 2 2 9 0 9 2 9 12 2 7 9 7 9 2 12 2 2
36 9 9 3 13 1 12 9 3 12 12 15 9 2 12 5 9 0 9 2 12 5 9 2 12 5 9 7 9 7 12 5 9 0 9 2 2
17 0 9 7 9 0 9 4 13 1 9 0 9 7 9 1 11 2
8 0 9 1 9 9 1 9 9
41 7 3 2 16 12 1 0 9 0 9 0 9 13 9 0 2 0 7 0 9 9 15 9 2 13 1 0 9 9 1 9 9 2 7 3 7 1 9 9 9 2
11 0 0 9 3 3 13 0 9 0 9 2
26 3 15 13 0 2 3 0 9 0 7 0 9 2 7 3 13 7 9 2 15 10 9 0 9 13 2
3 9 0 9
11 9 0 9 13 0 9 9 1 0 9 2
23 10 9 9 15 3 3 13 1 0 9 11 1 0 0 9 2 3 9 9 9 0 9 2
27 1 10 9 9 13 3 12 0 9 9 2 0 9 0 2 12 5 2 7 0 9 9 2 12 5 2 2
44 9 2 3 2 9 9 11 2 1 12 9 11 2 1 9 9 9 0 9 1 12 1 12 9 2 0 1 9 2 12 2 13 3 1 0 9 1 9 9 9 12 10 9 2
36 16 3 9 9 11 13 1 9 0 9 0 9 2 12 9 11 13 1 12 2 9 2 2 1 11 15 1 10 9 13 3 0 9 2 11 2
73 13 2 14 9 1 0 9 1 9 9 2 13 13 2 16 1 9 0 9 9 2 12 2 9 2 13 3 12 5 9 1 9 11 2 3 0 9 1 0 9 9 2 11 2 11 2 11 2 11 2 7 1 9 1 0 9 2 12 2 9 2 0 12 5 2 3 3 0 9 1 11 2 2
53 1 9 1 9 9 1 9 1 9 12 2 12 7 12 15 9 1 9 0 9 3 13 1 9 0 9 1 9 2 0 11 2 11 2 11 7 11 2 3 0 9 4 13 1 11 9 7 1 9 11 2 9 2
23 1 11 15 1 0 9 10 9 13 9 2 3 12 9 15 15 13 2 11 7 0 11 2
26 1 0 9 9 1 0 7 0 9 13 9 2 7 15 3 1 0 7 0 9 2 0 0 0 9 2
20 9 1 11 3 13 1 9 0 9 9 9 1 0 9 0 7 0 9 9 2
2 0 9
24 9 9 1 9 13 2 1 9 0 9 2 0 9 14 1 11 2 7 7 1 0 0 9 2
22 1 0 9 1 15 13 1 11 3 12 1 9 0 2 7 1 11 15 1 12 12 2
17 9 9 9 9 1 9 13 1 0 9 13 0 0 9 12 9 2
23 9 1 0 9 2 16 0 0 9 9 9 2 15 13 1 0 11 3 1 0 9 11 2
30 13 2 3 3 16 1 9 0 9 2 16 9 9 15 3 13 1 9 9 9 1 9 1 9 2 9 2 12 2 2
46 1 9 0 1 9 0 9 9 1 0 9 13 12 2 12 9 11 2 1 3 16 12 5 15 13 9 11 2 3 9 12 2 13 1 12 5 13 1 9 11 2 9 2 12 2 2
38 0 9 1 9 1 0 9 3 13 1 9 0 1 0 9 9 1 9 2 0 9 9 2 9 7 9 2 2 12 5 1 9 0 1 0 9 2 2
35 1 9 11 4 0 9 9 1 0 9 2 0 9 9 2 1 0 9 9 13 0 9 9 1 9 0 9 2 0 7 0 9 9 2 2
43 1 9 1 9 1 9 2 12 7 12 15 10 9 11 7 11 1 9 2 12 2 13 2 9 2 3 12 0 7 12 0 15 15 3 13 2 0 11 7 0 0 9 2
3 9 7 9
31 0 9 9 1 9 0 9 9 2 12 2 2 9 7 9 2 13 1 9 1 0 9 9 1 9 0 9 7 1 9 2
30 1 9 2 12 15 13 12 9 0 9 9 1 0 9 2 9 0 9 0 7 0 9 7 0 9 0 9 9 11 2
37 0 9 2 0 3 0 9 1 11 2 9 11 2 2 13 3 3 0 9 9 2 0 9 9 0 9 2 3 2 9 11 3 16 12 5 2 2
14 13 13 2 16 9 11 3 3 13 0 9 1 9 2
30 0 9 1 9 7 9 0 9 2 9 11 2 13 1 0 0 9 2 0 9 2 9 2 9 2 0 9 3 2 2
3 9 0 9
23 1 9 2 12 13 13 12 9 1 0 9 9 1 9 0 9 2 0 11 7 0 11 2
23 1 0 9 11 7 3 1 12 9 11 2 11 7 11 2 13 9 9 1 10 9 0 2
33 0 9 9 1 9 0 9 4 13 1 9 1 0 9 2 9 9 2 7 3 7 9 2 9 1 0 9 9 1 9 9 2 2
30 1 0 9 9 1 9 13 3 3 2 9 9 9 1 9 9 2 0 7 0 2 7 1 9 1 9 11 7 11 2
11 9 0 9 1 9 9 13 10 0 9 2
52 16 0 9 9 1 9 0 9 9 13 3 0 9 0 7 0 2 3 0 13 1 11 2 7 3 1 11 2 11 2 1 9 12 7 12 2 7 11 2 1 9 1 9 13 9 0 9 3 1 9 0 2
12 9 13 0 9 9 9 9 1 9 0 9 2
38 1 0 9 11 2 11 2 11 2 1 1 10 0 9 13 9 1 0 9 3 0 2 7 3 0 13 1 9 0 11 2 11 2 11 7 0 11 2
5 9 1 0 9 9
5 1 9 9 1 9
23 1 9 0 7 0 9 9 1 9 9 9 7 9 4 1 12 9 13 0 9 1 9 2
28 0 9 0 9 13 1 9 1 9 0 9 2 0 9 12 2 3 1 9 2 12 2 7 9 0 9 12 2
16 1 1 0 9 9 4 13 7 13 3 9 0 9 9 9 2
36 0 9 13 0 9 1 9 9 9 1 9 7 9 2 3 2 9 0 9 9 1 9 7 9 2 2 13 9 2 12 7 9 2 12 2 2
41 16 1 9 15 13 12 9 0 9 9 9 1 10 9 2 0 1 0 11 7 0 1 11 2 2 1 9 2 1 9 11 2 13 1 9 0 9 3 9 11 2
26 9 9 2 16 12 1 9 0 9 9 2 13 1 0 11 0 2 1 9 10 9 15 13 3 3 2
18 0 9 9 13 1 9 2 11 2 11 2 11 9 7 11 1 11 2
4 0 9 0 9
5 1 9 1 9 9
44 1 9 11 15 3 13 0 9 1 9 16 1 9 9 1 3 0 9 9 2 3 2 3 4 3 3 13 2 9 1 9 2 9 12 2 12 2 12 2 12 2 12 2 2
16 3 13 9 2 12 2 9 0 1 9 9 15 13 1 9 2
35 9 1 0 9 2 9 7 9 2 13 0 9 1 9 0 1 0 9 2 1 0 9 13 9 9 1 9 2 7 3 1 9 0 9 2
47 1 1 15 2 16 1 0 0 9 2 1 9 12 9 2 13 0 9 1 0 9 7 1 9 12 9 3 3 1 0 9 2 13 15 9 0 7 0 9 1 9 9 9 1 9 9 2
22 1 9 9 9 1 0 9 13 13 1 0 1 11 12 9 2 0 11 7 0 11 2
63 16 0 9 2 0 11 2 1 0 9 9 7 9 2 7 3 3 1 0 9 9 0 9 2 13 0 9 9 1 15 0 9 2 0 9 2 0 0 11 2 1 0 9 9 2 3 2 0 9 2 4 13 0 9 1 9 0 9 7 9 7 9 2
1 9
24 9 0 9 1 0 12 9 13 3 1 10 0 9 2 3 15 13 13 9 1 9 0 9 2
64 3 3 2 16 13 1 0 9 13 0 9 1 9 11 1 9 9 0 9 2 1 12 9 13 9 0 9 1 0 9 2 1 9 0 0 0 9 2 3 13 13 1 9 9 1 9 9 2 3 2 3 9 9 9 1 9 0 9 2 9 2 12 2 2
63 13 2 14 9 1 0 7 0 11 7 1 0 0 9 2 13 1 9 9 0 7 0 2 0 9 2 0 9 2 9 0 0 9 2 9 0 0 9 3 2 2 2 13 3 13 9 1 9 0 9 9 14 1 9 11 2 7 7 1 0 0 9 2
3 0 0 9
31 13 2 0 9 2 1 9 0 9 3 13 7 13 0 9 2 7 16 1 10 9 13 9 9 9 2 13 3 3 9 2
29 1 12 2 9 9 9 2 12 15 13 3 1 12 2 9 2 0 2 0 9 2 15 13 9 10 2 9 2 2
2 12 2
16 16 4 13 3 15 0 16 0 9 2 13 9 9 0 9 2
54 9 2 16 0 9 0 1 9 2 13 15 15 2 2 13 11 2 11 3 2 2 0 9 2 7 13 2 1 9 11 2 11 2 2 2 9 15 13 2 16 10 9 13 10 0 9 2 0 1 9 9 2 2 2
16 3 13 2 16 15 2 15 4 13 9 2 13 14 0 9 2
18 2 16 4 9 13 1 0 9 2 13 15 15 1 0 2 0 9 2
7 3 0 0 9 13 3 2
23 9 13 1 9 0 2 12 2 0 9 1 9 2 0 9 1 9 13 0 9 0 2 2
14 13 7 1 9 0 9 7 4 13 3 1 0 9 2
24 0 9 13 3 15 2 13 0 0 9 3 0 2 16 4 1 15 13 4 13 9 0 9 2
29 1 0 10 9 4 3 13 0 9 2 15 4 0 13 2 7 7 2 1 0 9 2 7 13 2 9 10 9 2
19 0 9 13 3 13 1 9 9 7 9 2 3 1 9 0 7 0 9 2
17 10 9 13 3 2 1 15 2 16 13 0 9 1 9 0 9 2
30 0 9 10 9 3 13 0 9 2 9 2 1 0 9 2 2 9 2 2 7 13 3 1 0 9 1 9 0 9 2
2 12 2
41 1 0 9 1 11 2 11 2 9 12 2 12 2 12 2 15 11 2 11 13 0 9 0 9 2 2 2 11 2 13 3 2 16 0 9 13 3 1 9 0 2
33 2 10 9 2 15 13 2 16 13 1 9 2 15 13 9 9 9 2 7 10 9 16 9 13 1 11 13 2 13 1 0 9 2
19 1 11 2 11 13 0 9 1 0 9 1 0 9 2 16 13 0 9 2
34 16 9 13 1 0 9 2 13 1 11 2 11 9 0 9 15 2 16 13 2 14 2 3 0 2 0 9 0 2 3 3 13 9 2
21 0 9 15 3 13 15 2 16 13 9 0 9 1 0 0 9 0 9 0 9 2
5 15 3 3 14 2
4 9 2 11 11
5 0 9 1 0 11
27 1 0 9 1 0 11 4 13 10 9 1 9 1 12 9 2 15 13 0 9 9 7 0 9 0 9 2
35 10 9 2 0 0 2 15 3 13 1 0 9 2 15 13 3 0 7 13 3 9 2 9 7 0 9 0 9 2 0 3 9 0 9 2
13 0 9 13 14 0 9 2 3 1 3 0 9 2
8 9 9 4 13 1 0 11 2
16 1 0 9 0 15 13 1 0 9 0 9 1 0 9 11 2
40 3 0 0 9 13 9 0 7 2 0 9 7 9 9 2 1 14 12 5 9 14 12 9 3 1 9 2 3 13 1 9 9 2 9 9 7 9 0 9 2
7 12 0 0 9 4 13 2
9 9 12 2 2 2 12 9 1 9
21 3 13 0 2 7 16 13 15 0 2 16 1 0 9 9 13 7 1 0 9 2
30 16 15 13 0 9 9 2 13 0 13 0 9 9 2 16 3 4 3 13 9 2 1 15 12 9 13 12 9 0 2
18 0 9 13 2 16 14 1 0 9 0 13 3 3 1 0 9 9 2
22 3 13 0 13 7 10 0 9 2 9 0 9 1 0 9 11 2 11 7 0 9 2
18 13 13 2 16 13 1 0 0 9 2 7 14 1 0 9 0 9 2
2 11 11
8 9 9 1 9 0 9 1 9
29 1 0 9 0 1 9 9 7 1 9 1 9 0 9 1 9 13 0 9 1 0 9 7 9 2 9 0 2 2
17 3 15 13 1 0 1 9 14 9 2 15 7 13 10 9 9 2
36 9 1 10 9 1 9 9 13 0 9 1 9 7 3 1 9 1 9 15 1 15 13 9 9 9 2 9 0 9 2 9 2 9 1 9 2
22 10 9 13 13 0 9 7 13 9 0 9 9 2 0 11 12 2 12 2 12 2 2
2 11 0
5 11 11 2 9 9
25 1 12 9 1 9 2 12 2 0 11 11 1 10 9 2 13 1 9 1 0 9 0 9 9 2
21 13 15 9 2 1 10 9 11 13 9 1 9 9 15 2 16 9 7 16 9 2
56 1 9 2 7 9 1 9 2 1 9 7 9 2 1 9 2 3 3 9 9 2 0 0 9 1 0 9 2 13 15 9 9 2 15 9 3 13 7 13 3 2 16 9 13 3 16 9 0 0 9 0 15 1 0 9 2
19 11 13 15 1 9 3 0 1 9 2 7 7 15 15 7 9 13 3 2
28 0 0 2 9 2 13 0 9 2 7 9 16 9 0 0 9 9 7 3 2 3 15 0 1 9 0 9 2
21 7 13 15 7 10 9 1 0 0 9 7 0 9 2 15 1 11 13 9 0 2
33 0 0 9 13 9 2 0 9 2 7 3 1 15 9 2 3 1 9 0 9 2 15 1 9 9 3 13 1 9 9 0 9 2
32 7 3 15 1 9 0 9 1 9 13 13 9 2 1 10 9 15 3 3 13 0 9 9 0 2 1 15 13 0 0 9 2
23 7 3 13 0 0 9 2 7 7 0 9 9 0 2 0 9 7 9 1 9 2 2 2
43 9 16 9 15 11 13 13 14 9 2 12 2 3 1 0 11 3 13 9 2 7 3 15 1 15 13 3 7 3 2 16 1 11 2 1 11 2 1 11 7 1 11 2
31 15 2 15 15 1 10 9 13 1 10 9 2 9 7 3 7 9 2 13 3 0 2 9 13 3 3 1 9 1 9 2
41 3 13 9 3 1 10 9 0 9 2 9 7 3 0 7 0 9 7 9 2 3 15 11 3 3 13 11 11 2 9 15 3 0 2 7 3 0 9 0 9 2
25 1 10 9 7 11 13 3 0 9 2 9 9 2 15 15 9 13 2 7 15 3 13 7 9 2
49 1 9 2 3 1 15 9 9 13 3 3 0 2 11 3 16 4 13 2 16 12 1 0 9 12 2 9 13 1 9 9 0 7 15 3 0 9 2 9 7 1 15 13 3 9 16 0 9 2
19 3 15 2 3 1 9 9 1 9 10 9 2 13 11 1 10 0 9 2
17 0 9 0 0 9 1 9 0 9 13 10 9 1 9 3 0 2
68 3 3 13 15 1 9 0 2 13 15 10 9 2 7 15 13 2 13 3 3 7 3 15 13 2 7 7 15 13 2 16 11 11 2 0 9 7 9 2 15 13 9 16 15 0 2 13 15 3 2 7 1 9 3 3 0 2 7 13 15 13 2 15 13 1 15 0 2
2 11 11
2 13 3
50 0 9 9 7 7 9 0 0 9 0 0 9 13 1 15 2 16 0 11 13 0 9 2 9 9 2 9 1 9 9 1 0 9 2 9 2 9 7 9 9 2 15 15 13 1 9 0 9 9 2
6 13 15 3 9 9 2
24 3 15 3 13 2 16 13 9 1 9 2 1 15 4 13 13 1 9 14 12 9 9 9 2
20 7 7 13 3 0 2 3 0 3 2 0 2 9 2 3 0 0 0 9 2
52 9 9 13 9 2 4 13 0 9 1 0 0 9 2 13 1 9 9 2 15 1 15 13 9 2 13 10 0 9 2 9 2 13 15 1 0 9 9 7 13 15 15 0 14 16 4 13 9 0 0 9 2
38 7 16 0 9 13 3 0 2 9 9 0 9 2 9 1 9 0 7 0 9 2 3 3 1 10 9 3 13 9 9 1 3 0 7 7 0 9 2
17 9 9 13 15 0 2 16 9 0 0 9 1 0 9 13 0 2
32 16 0 9 13 3 0 1 15 0 9 10 9 2 1 9 2 15 13 2 13 1 0 9 2 9 0 9 13 3 1 15 2
41 3 13 1 0 9 2 1 9 1 9 12 9 15 9 13 3 1 9 9 2 1 9 0 3 1 9 12 9 7 1 9 1 9 12 9 3 1 12 9 9 2
19 0 9 1 0 9 13 1 0 9 0 2 9 13 3 3 9 0 9 2
44 14 16 4 9 1 12 13 16 1 9 0 9 13 1 9 9 1 0 9 2 7 1 15 0 0 9 7 9 0 9 13 9 1 0 9 1 9 2 16 13 0 9 9 2
21 0 9 1 9 7 0 2 2 9 2 3 0 9 13 3 9 3 0 7 0 2
25 0 9 9 7 9 2 3 9 1 15 13 0 9 2 7 10 0 9 2 13 3 9 3 0 2
6 1 9 15 13 9 2
20 3 9 9 7 9 9 13 2 9 2 1 15 0 2 3 13 0 9 9 2
50 7 13 15 9 3 0 2 16 13 14 3 13 2 16 1 15 4 13 0 9 2 7 16 3 2 1 9 9 13 9 0 9 3 0 0 9 1 0 9 2 3 16 13 15 1 9 9 2 9 2
22 9 7 9 2 10 2 1 9 9 1 0 9 13 10 9 2 3 3 1 0 9 2
9 13 0 9 2 15 13 1 9 2
23 9 3 13 1 15 2 16 9 0 9 9 13 1 9 1 9 1 9 9 1 10 9 2
44 16 13 1 9 0 7 0 9 0 9 9 2 1 15 9 13 2 0 7 13 3 9 2 3 14 13 9 2 10 15 13 14 9 2 1 15 4 15 9 13 7 13 13 2
16 13 9 9 0 15 1 11 7 11 13 0 9 10 0 9 2
23 7 16 13 1 0 9 11 1 15 0 2 13 2 16 1 9 9 13 11 10 9 9 2
36 3 3 13 9 0 1 0 9 7 0 9 7 2 9 2 2 15 13 1 0 9 0 9 1 9 0 9 2 7 13 3 7 9 9 0 2
50 1 0 9 13 0 2 16 1 9 9 13 0 9 9 7 9 7 9 15 13 2 3 3 3 2 13 1 9 2 9 2 15 13 1 9 2 9 2 7 9 1 9 9 2 9 2 10 0 9 2
36 7 9 13 0 7 0 9 2 1 15 13 9 0 9 2 9 1 15 15 1 0 9 13 9 7 9 9 2 10 9 2 9 7 7 9 2
23 7 16 4 13 0 9 2 9 9 2 9 2 9 7 9 13 10 2 0 2 9 13 2
33 16 3 1 0 9 14 13 2 13 15 13 0 9 7 7 15 2 9 2 3 3 2 14 3 16 9 0 0 9 11 2 13 2
10 3 15 10 9 2 1 0 2 13 2
27 7 3 2 13 2 14 9 1 0 9 0 2 13 15 1 10 9 2 15 13 2 13 15 1 10 9 2
17 7 9 15 13 2 16 4 13 15 7 16 15 9 13 3 0 2
31 14 15 13 0 9 1 9 0 12 9 9 2 0 15 1 9 9 0 10 9 2 12 9 1 9 3 12 9 1 9 2
6 13 15 3 15 13 2
26 4 2 14 13 13 10 9 1 0 9 0 1 9 2 13 15 15 2 16 13 1 9 1 0 9 2
36 7 10 9 15 0 3 13 2 13 9 11 11 2 7 1 0 9 2 12 2 11 15 1 0 9 13 11 11 2 11 7 11 11 2 11 2
23 11 13 9 2 15 3 1 12 9 9 13 1 9 9 2 9 2 0 9 7 0 9 2
63 9 1 9 2 9 7 9 9 0 9 2 3 13 12 9 2 13 2 3 2 9 7 9 0 9 2 1 9 1 9 7 3 2 9 7 9 2 3 14 9 9 1 0 9 13 9 2 13 15 1 0 9 2 7 15 13 9 2 15 9 13 9 2
54 3 2 16 1 9 2 16 13 1 9 10 9 7 1 9 2 16 15 4 13 1 9 0 9 1 9 1 9 9 2 3 13 13 9 1 9 9 7 9 9 7 2 13 2 15 1 9 9 12 9 9 2 12 2
12 13 2 14 9 3 14 0 13 0 0 9 2
17 7 3 15 13 12 9 2 9 1 9 9 7 3 1 10 9 2
28 11 7 11 13 7 0 9 10 9 7 13 2 16 1 9 1 9 12 9 13 3 9 1 9 12 12 9 2
21 15 2 3 13 0 2 13 0 9 9 15 9 2 0 3 16 9 0 9 0 2
19 1 15 9 13 0 9 2 16 0 9 13 9 9 2 15 13 13 3 2
29 13 3 13 9 9 1 15 4 1 9 2 9 7 3 13 1 9 2 13 2 7 3 1 0 9 13 10 9 2
37 3 15 15 13 2 1 0 9 9 2 1 9 9 0 9 9 2 9 7 0 0 9 1 0 9 7 13 15 9 7 9 9 1 9 0 9 2
9 13 4 15 0 1 9 9 13 2
45 9 2 16 9 13 1 0 9 3 0 7 16 1 0 12 9 13 9 0 9 2 7 13 15 2 16 7 1 0 9 9 1 10 9 13 3 2 4 15 13 1 9 3 13 2
16 7 7 9 0 9 1 9 9 1 10 0 9 4 13 9 2
11 3 2 16 4 13 3 9 13 3 3 2
17 16 13 1 15 2 15 15 1 9 13 3 0 9 2 4 13 2
33 11 2 15 13 1 0 9 9 2 13 2 16 9 3 2 9 2 9 9 7 9 13 3 1 10 9 2 3 1 10 9 13 2
49 16 13 2 7 13 15 1 10 9 7 3 7 3 13 9 13 2 16 13 1 15 12 2 12 7 12 9 9 3 0 2 16 4 15 15 13 9 7 3 9 1 15 16 4 10 0 9 13 2
2 11 11
1 9
10 9 16 9 7 3 15 13 2 13 9
2 11 11
12 11 2 11 2 11 7 9 2 9 9 9 2
10 11 11 12 2 12 9 2 12 9 2
28 1 9 13 9 2 11 11 2 9 9 2 7 2 9 1 9 2 9 0 9 2 2 13 9 2 11 11 2
22 9 13 1 0 9 9 9 9 9 7 9 10 0 9 2 15 13 0 9 0 2 2
18 1 0 9 0 9 13 7 9 9 7 0 2 9 2 2 3 9 2
7 10 9 15 13 0 9 2
38 1 9 13 9 2 1 9 0 9 7 0 9 2 7 1 0 9 15 13 1 9 15 2 16 15 13 10 9 2 9 2 7 10 9 2 9 2 2
14 1 9 9 7 9 9 1 0 9 9 13 9 9 2
18 13 9 2 13 3 2 3 13 11 2 11 2 16 15 13 9 11 2
23 0 0 9 13 9 1 9 9 1 10 9 7 1 9 2 15 15 13 7 13 10 9 2
36 9 9 13 13 9 9 0 9 2 1 0 0 9 15 13 0 9 2 0 9 1 9 11 15 13 1 0 2 0 2 9 1 9 11 2 2
11 13 15 3 2 0 2 0 9 9 9 2
65 16 9 13 9 10 9 7 10 9 13 1 9 3 0 9 2 16 13 9 0 9 2 9 9 1 9 2 13 9 9 2 9 3 2 2 16 9 9 13 13 0 0 9 2 13 9 9 0 9 2 9 2 3 13 1 9 1 9 2 15 15 1 9 13 2
40 3 2 3 9 13 9 1 9 1 0 9 2 9 2 9 2 2 1 15 13 9 1 9 7 0 9 1 9 2 13 15 0 7 0 9 0 2 9 2 2
41 13 15 1 9 2 1 0 9 2 2 15 13 14 0 9 1 9 9 7 9 7 1 9 2 15 15 7 3 13 1 9 2 7 9 2 1 0 2 9 2 2
19 7 15 13 3 9 0 9 7 3 7 15 2 15 15 1 10 9 13 2
28 13 15 3 15 2 7 9 0 16 0 9 2 0 9 9 0 9 2 0 1 9 0 9 0 9 0 9 2
27 9 9 15 1 10 9 13 2 13 1 9 0 0 9 2 7 15 1 10 9 2 1 15 1 9 13 2
15 15 3 16 0 9 13 9 0 9 14 9 0 10 9 2
19 13 3 1 9 0 9 2 7 3 10 9 13 14 0 9 1 10 9 2
13 0 0 0 9 15 13 10 9 2 9 2 9 2
15 15 13 3 0 2 16 0 15 9 13 1 9 0 9 2
21 13 7 2 16 1 9 13 3 1 0 0 9 9 9 2 0 0 2 9 2 2
38 3 3 13 13 2 16 13 9 2 1 15 9 13 10 0 9 2 7 13 15 14 1 15 2 15 13 0 9 2 7 3 3 13 3 16 15 15 2
34 16 13 9 13 1 9 7 9 13 0 2 3 13 15 3 9 9 1 9 0 9 2 16 4 13 13 2 16 9 9 13 3 0 2
12 3 13 0 9 7 9 16 0 9 7 9 2
31 3 4 13 1 15 9 2 15 4 13 2 13 7 13 2 9 2 15 1 0 9 1 15 2 1 15 13 2 3 13 2
9 3 2 16 15 10 9 7 13 2
14 15 4 13 3 1 9 2 16 4 13 1 9 0 2
31 7 16 4 15 13 2 16 9 13 13 0 9 2 13 15 9 0 9 14 0 9 2 7 7 9 7 3 7 9 9 2
10 13 3 1 9 13 12 0 0 9 2
34 12 7 15 15 13 2 13 15 2 0 3 2 2 0 9 2 7 0 9 2 7 3 7 0 9 15 2 3 14 0 0 9 13 2
16 16 9 0 9 1 15 10 13 2 13 10 9 13 0 9 2
47 7 3 3 13 1 10 0 9 0 2 13 15 1 0 9 9 0 2 0 7 0 2 16 0 9 2 15 4 3 2 7 15 3 9 0 9 2 13 16 2 0 2 2 0 9 2 2
13 3 15 1 0 7 0 9 13 9 9 2 11 2
23 13 9 15 2 15 4 13 2 15 15 1 0 9 13 7 15 15 1 15 13 9 15 2
58 13 9 0 2 11 7 0 2 2 13 3 13 1 9 2 16 7 1 10 0 9 2 1 15 4 3 2 1 0 7 0 0 9 2 7 3 7 3 2 13 9 0 7 3 2 7 15 14 1 9 0 2 15 15 13 13 2 2
24 13 15 15 7 9 7 9 1 0 0 9 2 3 15 2 15 13 13 16 2 0 2 9 2
33 13 1 9 9 2 16 3 9 1 9 9 7 1 0 9 13 1 9 3 10 1 9 1 15 2 15 13 13 1 0 9 9 2
17 10 9 15 13 0 9 2 9 9 0 9 7 0 9 0 9 2
45 0 9 10 0 9 13 9 2 16 0 9 2 9 2 7 3 7 9 4 3 13 9 2 15 15 1 0 0 9 3 13 1 3 0 2 3 0 2 9 2 11 2 11 2 2
37 16 15 3 13 1 9 15 2 1 15 15 13 2 12 0 9 2 1 9 10 9 2 7 3 15 13 9 9 10 9 2 13 15 13 9 9 2
15 4 13 1 9 9 2 16 1 10 9 1 10 9 13 2
59 1 9 2 3 0 9 13 0 2 3 3 0 9 1 9 9 2 7 15 3 7 2 16 9 1 10 9 3 13 2 0 9 9 13 3 0 7 16 9 15 1 3 0 9 3 3 13 2 13 0 15 13 9 2 0 9 2 11 2
8 13 15 3 10 0 9 9 2
6 13 15 2 16 14 2
37 13 4 15 3 13 1 15 2 15 13 0 9 2 1 15 13 0 9 2 15 15 13 1 0 9 2 7 3 1 0 9 13 4 13 0 9 2
40 3 16 9 9 2 9 7 9 2 13 0 0 9 2 15 13 1 9 9 2 0 9 2 7 3 3 9 9 2 1 3 0 2 7 7 13 9 0 9 2
41 9 13 15 0 2 0 0 9 1 0 9 7 1 9 3 2 0 9 0 0 9 7 3 7 0 9 0 9 2 15 1 0 9 10 9 13 3 3 0 9 2
17 9 9 13 0 2 15 13 0 0 9 7 13 0 9 2 0 2
8 1 9 0 15 10 9 13 2
16 3 13 15 3 1 9 1 0 9 2 0 9 1 0 9 2
17 1 9 13 9 1 2 0 9 2 2 2 3 0 9 2 3 2
13 13 15 0 15 2 16 15 15 3 1 9 13 2
22 7 3 11 2 16 13 15 9 1 0 9 0 0 9 2 15 13 3 0 0 9 2
14 3 13 15 14 9 1 9 0 9 7 0 9 9 2
111 13 2 14 7 9 1 9 3 2 9 0 9 2 9 2 15 4 3 13 1 9 0 9 2 3 13 1 0 9 2 7 1 0 9 2 15 4 13 1 9 2 15 15 13 7 13 13 13 1 0 9 2 1 9 9 0 7 0 2 1 9 3 9 0 2 2 3 7 3 7 7 2 16 4 13 10 0 9 1 9 2 16 13 2 16 1 9 9 13 9 9 7 9 3 0 16 9 9 2 7 3 2 1 9 2 10 9 0 9 9 2
24 13 2 14 9 2 1 15 13 3 9 2 9 2 3 2 2 13 3 3 14 15 1 9 2
2 9 2
49 9 10 9 13 3 0 2 16 1 10 0 9 10 0 9 13 0 0 9 2 7 7 0 9 4 13 1 10 0 9 2 15 13 7 9 0 2 7 9 0 2 14 7 9 3 7 3 0 2
32 16 4 13 10 9 1 9 0 2 1 15 13 9 0 9 1 15 1 12 9 0 2 13 4 15 2 16 4 15 9 13 2
55 9 0 13 14 13 2 16 4 15 9 13 2 16 1 9 15 0 13 7 14 3 13 2 7 3 15 13 13 2 16 15 2 15 15 13 3 1 0 9 2 13 7 15 2 1 15 13 9 2 7 0 9 0 9 2
26 15 2 16 9 13 0 9 2 14 13 1 9 2 16 10 0 9 2 3 2 9 2 4 13 9 2
11 9 2 9 2 2 9 4 1 9 13 2
6 0 9 7 0 9 9
37 0 9 0 7 0 0 9 13 0 1 9 2 12 2 3 11 2 11 13 9 9 2 15 13 13 7 1 15 13 9 0 9 0 0 9 3 2
11 1 0 9 3 15 0 9 10 9 13 2
39 1 9 13 0 2 16 12 9 0 9 3 3 13 2 7 0 13 13 3 2 1 0 9 7 9 2 0 1 9 7 9 9 2 9 9 7 0 9 2
7 13 15 7 1 0 9 2
43 13 2 14 15 9 1 9 0 9 0 0 9 1 0 0 9 2 3 2 2 13 9 2 2 13 1 15 9 1 0 9 3 0 9 16 9 1 0 9 1 9 0 2
22 1 0 0 9 9 1 9 15 13 1 9 2 12 2 7 9 13 1 0 0 9 2
13 10 9 7 13 3 1 0 9 2 0 1 0 2
34 1 9 0 9 0 9 0 9 1 9 13 10 9 1 9 9 2 9 7 9 2 0 2 11 2 11 2 12 2 12 2 12 2 2
17 1 0 9 10 0 9 15 13 3 1 0 0 9 2 3 9 2
2 11 11
3 12 2 12
6 13 0 0 9 1 9
12 1 0 9 13 9 1 9 1 3 0 9 2
16 13 15 1 9 2 0 2 9 2 0 9 7 9 0 9 2
21 3 2 9 1 0 9 13 1 0 9 1 9 12 2 12 2 12 12 0 9 2
35 1 1 15 2 16 0 0 9 0 0 0 9 13 9 0 0 9 1 9 1 0 0 9 2 7 9 7 9 13 9 13 10 0 9 2
30 1 0 9 7 10 9 1 9 1 9 12 4 13 9 9 7 3 15 13 2 16 10 0 9 4 13 1 0 9 2
10 9 13 9 0 3 0 0 9 9 2
30 10 9 15 13 1 9 7 9 1 9 1 9 12 9 7 1 12 9 7 13 3 1 9 0 0 9 1 0 9 2
20 0 9 13 1 0 0 9 2 13 1 9 0 9 0 9 1 9 1 9 2
13 0 9 0 9 10 0 9 13 7 9 7 9 2
10 3 15 13 1 2 0 2 0 9 2
44 13 0 2 16 16 13 1 9 1 0 9 0 0 9 0 9 0 9 9 2 13 14 1 0 9 0 12 0 9 2 7 7 1 9 9 0 2 3 1 9 0 0 9 2
34 10 0 9 13 0 9 1 9 9 1 9 1 0 9 1 9 2 7 15 14 1 9 9 1 10 9 2 7 7 1 9 0 9 2
14 4 3 13 9 9 3 0 9 0 0 9 1 9 2
16 4 13 9 1 9 9 1 0 9 2 9 2 9 7 9 2
37 13 3 7 1 9 1 9 9 0 0 9 2 15 9 0 9 3 3 13 2 7 3 1 11 7 11 15 13 3 1 3 16 12 9 7 13 2
2 11 11
41 2 2 2 1 9 4 15 1 10 0 9 7 1 10 9 13 1 0 9 11 2 15 13 9 2 0 2 9 2 3 2 0 9 2 7 0 1 10 9 9 2
43 13 14 15 0 9 2 7 1 10 9 9 9 13 2 16 9 2 13 2 14 15 1 0 9 2 13 7 13 7 16 4 13 0 9 2 3 9 10 0 9 3 13 2
6 3 15 10 9 13 2
26 0 4 15 7 1 0 9 13 3 2 7 3 7 1 0 9 2 15 13 3 0 9 9 2 2 2
4 11 11 2 11
11 9 2 9 13 3 0 3 16 0 9 2
8 0 9 9 13 11 7 11 2
13 9 9 7 9 9 0 9 13 11 9 2 12 2
8 0 9 13 0 9 0 9 2
12 13 15 0 0 9 1 9 9 0 1 9 2
27 10 9 13 9 0 2 9 2 9 2 7 0 0 9 2 9 0 2 0 0 9 2 9 2 1 9 2
16 9 9 0 9 13 0 9 2 0 9 13 3 0 9 2 2
44 0 9 13 3 2 1 0 9 9 7 9 2 7 7 1 0 9 9 2 9 2 9 2 9 2 9 2 9 2 7 7 9 2 13 9 12 2 12 2 12 2 12 2 2
9 1 9 13 14 12 9 9 3 2
37 0 9 0 9 2 0 9 4 13 2 0 0 9 2 0 3 9 2 4 13 7 13 16 9 7 16 9 1 9 0 9 2 0 2 0 9 2
11 3 0 0 9 15 13 16 9 0 9 2
7 9 2 11 11 2 9 2
4 0 9 13 2
2 11 11
24 3 9 9 13 9 2 16 9 13 12 0 0 9 2 15 13 9 2 3 9 1 9 9 2
17 9 0 9 15 3 13 1 9 12 0 9 2 0 0 9 9 2
19 3 4 3 3 13 0 12 0 9 2 16 15 0 9 15 13 1 12 2
37 10 0 7 0 9 13 10 9 2 14 1 9 2 3 9 0 9 7 0 9 0 9 13 2 16 3 0 2 2 0 2 0 9 13 3 12 2
13 0 9 2 3 2 0 2 0 9 13 3 12 2
35 3 15 13 3 2 16 0 9 2 9 2 3 13 1 12 12 9 7 13 3 3 13 0 9 2 9 2 2 15 13 14 12 12 9 2
21 0 9 0 13 9 7 9 0 9 2 9 9 7 0 9 13 1 15 3 13 2
17 0 2 0 9 0 9 3 3 13 1 0 7 0 9 1 9 2
5 13 15 13 9 2
16 3 13 2 16 9 0 9 13 13 9 1 12 0 9 9 2
19 12 2 1 0 9 0 9 1 0 12 12 9 13 13 0 2 0 9 2
22 13 13 1 12 0 9 2 0 0 9 9 1 9 2 0 15 9 0 9 7 9 2
21 15 10 12 9 13 0 9 2 9 2 0 9 2 15 13 3 0 9 0 9 2
31 0 9 13 1 0 9 2 13 2 14 9 9 0 1 9 7 0 1 9 2 13 0 9 7 9 11 13 13 0 9 2
17 13 2 14 3 0 9 1 0 9 2 9 13 7 13 9 0 2
19 12 2 1 9 2 3 1 9 13 9 2 13 15 0 0 9 0 9 2
8 9 13 14 12 5 0 9 2
21 15 0 13 9 0 9 2 15 3 9 15 13 3 1 9 7 15 0 13 9 2
20 13 3 0 9 9 0 9 7 9 7 3 15 0 0 9 13 9 9 0 2
28 12 2 3 13 0 9 3 0 0 9 2 16 13 0 13 0 0 9 0 3 2 9 0 9 7 0 9 2
17 0 7 13 2 16 4 9 13 7 0 9 9 13 0 9 9 2
20 16 4 9 13 3 0 2 13 4 14 12 9 9 9 1 0 9 7 9 2
27 3 13 2 1 9 0 0 9 13 10 0 9 2 15 4 3 13 2 7 3 3 13 7 10 0 9 2
16 9 1 0 9 13 13 9 0 9 2 15 13 0 0 9 2
44 1 0 9 4 3 0 9 0 9 3 13 2 13 0 9 7 0 0 9 13 13 9 2 7 2 9 0 9 2 15 3 16 10 9 13 0 9 7 13 3 0 0 9 2
7 2 9 13 9 9 2 2
28 1 10 9 15 13 0 9 13 10 9 9 2 15 4 13 0 9 2 7 4 13 0 9 7 9 0 9 2
21 9 0 9 13 9 0 9 1 9 12 9 2 15 13 9 1 0 12 9 9 2
17 1 0 11 2 3 0 11 2 15 13 0 9 0 2 9 11 2
11 0 9 1 9 0 9 4 13 0 9 2
11 9 1 0 0 9 13 9 10 0 9 2
16 1 0 9 15 13 13 3 0 12 9 0 9 11 2 12 2
26 4 1 15 13 1 9 12 9 3 12 9 2 15 4 13 7 1 15 4 13 0 9 9 7 9 2
15 0 9 0 9 4 1 0 7 0 9 1 12 9 13 2
33 0 0 9 4 13 1 9 9 7 0 9 0 1 0 9 2 9 2 7 1 9 1 0 9 2 11 2 2 13 9 2 12 2
18 0 0 9 1 9 0 11 2 11 2 12 2 13 10 3 0 9 2
27 2 0 9 9 13 3 0 1 9 0 1 0 9 7 1 9 1 0 9 2 7 13 15 1 0 9 2
18 2 0 9 13 0 7 13 1 0 0 9 2 15 13 12 12 9 2
29 3 2 1 0 9 12 7 12 13 3 12 12 9 2 16 1 9 12 7 12 13 12 12 9 12 2 12 2 2
11 0 9 15 1 0 12 9 9 3 13 2
50 2 0 12 0 9 13 3 0 2 13 0 9 1 9 11 2 12 2 2 7 9 2 9 1 15 13 2 13 1 12 2 12 9 9 0 16 0 9 2 9 2 13 9 12 2 12 2 12 2 2
8 2 9 13 3 12 12 9 2
25 2 0 9 0 9 13 3 0 7 1 9 0 0 9 2 0 9 4 13 1 0 9 0 9 2
25 9 1 0 9 1 0 11 13 0 9 1 0 9 0 7 0 9 2 7 15 13 13 0 9 2
31 0 9 9 0 0 9 13 1 9 14 12 9 7 9 0 1 9 15 13 3 10 12 9 2 16 13 1 9 9 9 2
23 7 3 15 15 13 3 0 15 2 10 0 9 15 1 10 0 9 13 1 0 9 13 2
1 9
22 11 2 11 2 11 7 9 2 2 0 12 0 0 9 1 9 1 0 11 2 11 2
8 11 12 2 12 2 12 2 12
7 1 0 7 0 9 9 9
2 11 11
32 0 9 2 9 2 4 13 1 9 3 9 2 12 11 7 11 7 0 9 13 14 9 2 12 1 0 9 0 1 9 11 2
25 10 9 13 13 1 0 9 2 0 2 2 0 2 2 15 13 7 1 9 2 9 2 0 9 2
12 0 9 13 3 9 3 16 2 9 2 9 2
33 0 9 1 9 2 2 9 2 2 13 13 9 2 9 1 3 0 2 0 2 9 9 15 7 13 3 1 9 14 1 10 9 2
34 0 9 7 0 9 4 1 0 9 13 1 0 9 9 7 13 3 0 9 2 16 3 1 0 9 2 7 1 9 2 9 7 9 2
28 13 15 14 13 1 0 9 1 9 0 2 9 7 9 1 9 2 9 2 9 9 7 9 2 0 9 0 2
16 9 16 9 9 2 9 7 9 13 1 9 1 0 9 9 2
28 0 9 13 9 10 0 9 1 0 9 0 9 7 1 10 0 9 2 3 0 3 1 0 9 12 2 9 2
37 3 3 13 9 7 9 9 7 9 3 0 2 16 14 0 9 9 7 9 2 0 0 9 2 13 9 2 13 3 0 9 7 13 15 0 9 2
19 0 9 9 13 3 9 10 3 0 9 7 0 9 1 3 0 0 9 2
26 1 0 9 9 9 9 1 9 13 2 7 10 9 13 1 10 0 9 0 9 7 1 9 9 9 2
17 3 0 13 9 9 7 9 1 9 2 9 7 9 1 9 3 2
32 0 13 1 10 9 7 0 9 0 9 1 9 7 9 1 9 2 3 16 3 0 9 3 0 7 3 0 9 0 0 9 2
35 3 1 0 9 4 0 9 0 9 2 3 2 0 9 2 13 1 0 7 10 9 15 13 3 2 9 9 9 16 15 0 1 9 2 2
44 1 10 9 4 3 13 2 16 1 10 9 13 10 0 9 1 9 1 0 0 9 2 9 9 9 2 9 9 9 2 2 16 1 15 13 10 0 0 9 2 3 0 9 2
45 9 7 9 0 9 13 3 4 1 12 2 9 13 1 0 9 9 1 9 2 3 15 14 1 9 9 3 13 11 2 11 2 9 0 9 2 7 3 16 9 2 16 0 9 2
19 12 2 9 15 3 13 0 9 7 9 1 0 9 2 3 2 9 2 2
13 3 4 3 11 7 11 9 2 9 2 3 13 2
44 1 0 9 9 2 3 0 9 2 4 3 1 0 9 12 2 9 3 13 9 3 0 9 2 15 13 3 0 9 7 0 9 2 7 16 9 15 10 9 13 3 3 0 2
35 3 11 13 10 9 3 0 9 2 7 3 9 1 0 9 1 0 9 2 15 13 2 9 2 2 3 2 0 9 0 2 0 9 9 2
1 9
6 11 2 11 2 11 2
4 2 12 2 2
10 9 1 0 0 9 1 0 0 9 2
4 9 2 9 2
2 11 2
2 11 2
9 11 2 11 2 2 11 2 11 2
8 2 12 2 0 9 1 9 2
7 1 9 9 7 0 9 11
29 2 11 11 3 1 9 2 16 15 13 9 2 7 14 0 13 9 10 9 2 13 2 16 9 13 0 16 9 2
17 7 3 9 0 9 3 13 10 9 7 13 15 3 1 10 9 2
14 9 9 13 1 0 9 9 7 9 7 13 15 9 2
13 0 9 13 0 9 9 0 9 7 9 0 9 2
31 15 0 13 2 15 15 13 1 9 2 15 15 13 0 9 2 15 0 13 15 1 0 9 0 1 9 13 0 9 9 2
12 9 13 9 2 7 9 7 3 9 13 9 2
28 9 9 0 2 13 15 2 1 9 9 2 15 3 14 13 1 9 9 0 9 0 11 7 0 9 1 0 2
3 11 11 2
15 15 13 10 11 1 10 9 7 15 15 13 13 1 15 2
18 2 3 13 9 0 9 2 15 13 0 9 7 13 13 1 0 9 2
16 13 7 3 9 0 2 13 2 14 10 9 0 9 0 9 2
29 1 0 9 13 3 13 9 2 3 9 0 13 1 9 13 1 9 0 9 2 7 10 0 9 13 1 9 11 2
23 13 13 0 9 9 2 1 9 13 9 0 9 9 2 15 1 10 9 13 3 16 3 2
19 1 9 9 13 3 9 9 0 14 1 9 2 9 9 2 3 9 0 2
34 3 13 0 15 13 2 16 9 2 0 2 3 13 1 9 2 0 2 2 16 0 13 15 2 15 13 9 7 9 1 0 9 9 2
14 15 13 0 9 2 15 13 1 10 9 9 0 9 2
35 0 9 1 10 9 9 7 9 13 1 9 9 3 3 16 10 0 0 9 2 7 13 1 10 9 0 9 3 13 13 0 9 16 9 2
19 16 4 1 9 1 10 9 13 9 9 2 13 4 3 13 14 9 9 2
13 2 12 0 9 0 9 4 3 13 13 0 9 2
17 13 15 9 1 0 9 0 1 9 1 9 7 9 1 0 9 2
19 10 9 13 3 2 16 15 9 13 3 13 1 10 9 16 1 15 0 2
15 0 9 13 1 10 9 13 3 1 11 7 3 1 15 2
15 13 15 7 1 9 7 3 15 3 13 1 0 0 0 2
11 1 9 11 11 13 10 0 9 12 11 2
5 12 13 9 9 2
25 11 11 15 13 1 9 0 7 13 1 9 2 10 9 11 11 15 13 1 9 7 13 1 9 2
29 0 0 9 15 13 1 9 0 2 14 7 2 16 4 12 9 4 13 0 2 7 16 1 9 9 12 11 13 2
17 9 0 13 9 11 7 0 9 2 7 13 9 1 9 3 13 2
16 13 9 2 0 2 0 9 1 9 0 11 7 13 0 9 2
13 1 9 0 15 13 0 9 0 0 9 0 9 2
21 3 13 1 9 13 2 16 0 1 0 9 0 9 13 1 9 2 3 1 9 2
17 2 1 9 11 11 13 11 3 2 16 15 13 0 13 1 9 2
16 9 13 9 7 9 9 2 16 9 0 3 9 13 0 9 2
13 1 0 9 15 11 13 9 9 7 9 1 9 2
11 13 3 0 9 1 0 9 0 0 9 2
31 1 0 9 4 9 13 9 7 9 9 2 15 13 7 13 0 9 9 7 3 13 0 9 0 1 9 10 9 10 9 2
7 1 9 13 0 16 9 2
27 11 13 10 9 1 9 2 7 3 7 1 9 2 9 9 2 15 15 2 13 2 3 13 1 0 9 2
29 0 9 3 13 10 9 2 7 2 3 1 9 0 2 0 9 9 3 13 1 3 0 7 3 0 0 9 2 2
10 2 15 13 1 15 0 9 11 3 2
25 9 0 7 0 2 15 13 0 9 2 9 9 9 7 0 11 2 15 15 3 13 1 0 9 2
39 3 0 9 1 10 9 15 1 9 12 2 9 10 9 13 0 9 2 7 3 15 13 1 9 2 15 15 13 9 2 12 2 14 12 9 1 0 9 2
23 9 0 9 4 3 13 10 9 0 1 0 0 9 2 16 15 15 9 0 13 1 9 2
24 13 9 2 1 15 13 1 0 9 0 0 9 2 1 15 12 9 15 13 14 0 9 9 2
10 9 4 3 0 9 3 13 1 9 2
32 1 9 9 13 1 0 9 3 9 7 1 9 0 0 0 0 9 15 9 12 0 1 0 9 13 16 0 2 3 0 9 2
13 7 12 9 9 7 9 15 1 15 3 13 13 2
28 7 7 13 2 14 15 13 1 10 9 7 3 3 9 1 0 9 2 13 4 15 13 1 0 9 0 9 2
20 13 2 14 15 3 9 9 7 9 2 13 15 3 3 9 9 7 9 9 2
2 11 11
4 0 9 0 2
2 11 11
5 1 12 2 9 9
2 11 9
21 11 1 11 15 13 1 9 11 2 3 11 2 1 0 11 1 0 9 0 9 2
9 9 9 15 13 1 9 1 9 2
28 3 1 10 9 13 9 0 2 11 2 1 10 9 15 1 9 0 2 11 11 13 9 2 3 13 10 9 2
10 10 9 15 13 1 9 12 2 12 2
21 0 9 11 1 11 13 9 1 0 9 7 1 9 12 2 12 13 7 9 9 2
14 9 13 11 2 7 1 9 11 2 3 0 1 11 2
16 11 15 15 13 16 0 1 11 2 11 9 11 1 11 2 2
9 14 1 10 9 15 13 9 11 2
12 1 9 11 1 11 15 13 14 9 2 12 2
17 3 13 0 9 2 16 9 2 12 13 9 0 9 0 9 0 2
2 11 2
29 13 12 2 12 2 12 7 3 15 13 0 9 1 9 2 1 10 9 11 1 11 13 7 3 15 3 14 13 2
7 9 11 1 11 1 9 9
18 9 9 0 1 0 9 7 10 9 13 1 9 9 2 12 0 9 2
18 9 11 1 11 1 9 9 7 9 0 9 4 13 7 13 9 0 2
16 9 13 1 0 9 0 9 1 9 0 9 2 9 11 11 2
22 11 13 9 2 16 4 13 1 0 9 15 0 9 7 13 0 9 1 11 1 11 2
10 13 3 9 0 9 7 13 0 9 2
27 1 10 9 13 9 0 9 7 11 1 11 13 3 9 1 9 0 9 2 15 0 9 11 1 11 13 2
16 0 9 10 9 13 7 9 13 1 9 9 1 9 10 9 2
19 0 9 3 13 0 9 1 3 0 9 0 2 1 0 9 11 1 11 2
28 9 2 15 13 1 10 9 1 10 9 1 11 2 4 13 9 2 16 4 15 13 1 11 7 13 0 9 2
25 9 12 2 12 2 12 13 1 0 9 1 0 9 1 9 11 1 11 2 11 11 7 9 11 2
10 0 9 15 13 1 9 1 12 9 2
14 9 12 2 12 2 12 13 0 9 13 9 7 9 2
28 3 1 9 9 7 11 12 2 13 9 7 13 13 11 11 2 11 1 11 2 0 9 11 11 7 9 11 2
13 9 4 7 1 9 10 9 13 7 13 1 11 2
16 0 4 13 1 0 9 1 0 9 2 3 15 13 0 9 2
22 3 13 7 1 9 11 13 1 9 9 1 9 9 7 9 0 2 9 2 12 2 2
12 3 4 3 13 7 13 1 9 14 1 9 2
16 3 15 13 1 9 2 1 9 7 9 0 2 7 13 9 2
5 9 0 15 13 2
8 13 11 1 11 7 11 11 2
33 9 0 9 7 9 13 14 3 2 3 4 2 13 2 7 13 1 9 2 7 2 13 1 0 9 1 9 7 13 1 9 9 2
16 3 4 13 9 1 9 2 3 2 16 4 0 9 13 2 2
7 3 4 13 1 0 9 2
15 1 11 4 13 7 9 2 15 4 13 9 9 7 9 2
30 9 0 9 9 13 7 13 13 0 2 1 9 2 2 7 2 3 13 1 9 7 9 0 2 16 15 13 9 0 2
14 9 13 0 13 9 7 1 9 15 13 13 15 13 2
30 7 15 13 9 2 14 1 11 1 11 2 13 13 9 0 2 1 0 9 2 16 15 13 2 3 4 13 7 13 2
4 3 4 13 2
10 1 9 11 1 11 13 3 7 9 2
12 0 9 13 15 7 0 11 14 13 9 0 2
25 11 1 11 4 1 9 13 1 0 9 1 9 11 9 12 2 12 2 12 1 12 2 9 0 2
14 0 9 7 1 9 9 4 13 1 0 9 0 9 2
39 1 9 9 12 7 12 2 12 9 9 2 0 3 0 0 9 9 1 9 0 9 1 11 4 13 2 16 11 11 13 12 2 2 9 2 10 0 9 2
45 1 12 9 2 9 12 2 12 2 12 2 3 12 2 12 2 12 2 13 9 11 1 11 1 0 0 9 2 3 1 0 9 1 9 9 1 9 0 0 9 0 2 9 0 2
18 1 15 13 12 1 0 9 1 0 2 9 0 1 9 12 2 9 2
21 9 13 2 16 9 11 2 13 13 1 9 1 9 9 2 12 2 9 2 2 2
14 10 9 13 1 9 1 0 9 9 1 9 2 12 2
37 3 15 13 3 2 2 16 1 9 0 2 9 2 7 2 12 2 9 2 15 13 1 10 9 0 0 9 1 11 11 2 15 9 11 13 13 2
15 11 1 11 4 13 1 9 1 9 9 1 0 0 9 2
11 9 0 2 9 0 4 9 2 12 13 2
20 3 3 1 9 12 2 9 12 4 9 13 1 0 9 2 0 15 9 9 2
11 10 9 13 0 13 1 0 9 0 9 2
24 9 0 9 13 7 9 9 1 11 0 9 0 9 11 7 0 9 11 1 12 2 9 12 2
18 0 9 13 14 9 9 0 9 7 0 9 2 7 7 0 9 0 2
13 9 15 13 3 13 9 15 0 9 11 1 11 2
21 1 9 0 9 1 9 0 2 3 13 11 1 11 9 2 13 9 0 12 9 2
7 0 9 1 9 11 1 11
31 0 9 1 0 9 13 1 9 11 1 11 7 4 13 1 9 1 9 2 15 11 1 9 9 2 12 13 9 11 12 2
17 10 9 4 13 1 0 9 9 2 12 1 0 9 9 2 12 2
25 1 0 9 13 2 16 10 0 9 4 13 7 2 16 13 10 0 9 7 13 15 3 0 9 2
11 0 9 13 0 9 11 11 1 9 0 2
16 9 2 12 13 1 11 3 16 1 9 2 7 9 9 13 2
15 0 9 13 1 9 7 9 1 0 9 15 13 14 3 2
16 0 9 13 16 0 9 2 7 7 9 9 1 11 1 11 2
40 0 9 1 9 11 1 11 13 0 9 11 2 15 13 2 16 9 11 12 2 13 13 0 9 9 7 9 9 11 3 7 2 16 15 13 13 0 0 9 2
15 7 15 13 14 9 0 9 11 1 11 16 9 0 9 2
25 0 0 9 11 1 11 1 12 2 9 12 2 9 1 9 1 0 9 13 7 9 11 1 11 2
10 1 9 13 0 9 9 7 0 9 2
19 16 9 9 13 9 2 12 2 3 1 12 9 3 2 16 15 9 13 2
22 10 9 7 13 1 11 1 11 2 7 1 11 1 11 2 15 13 14 1 0 9 2
8 9 9 13 13 7 9 9 2
24 1 0 9 0 9 12 4 1 10 0 9 13 1 0 9 9 9 2 7 7 13 9 12 2
29 3 3 1 9 9 11 1 11 13 9 9 2 11 2 7 9 9 2 11 2 0 9 2 11 9 2 11 2 2
8 0 0 9 13 9 0 9 2
25 10 9 2 16 3 15 13 9 2 7 9 2 13 0 0 9 0 9 11 1 11 1 12 9 2
17 1 9 12 2 9 4 10 0 9 13 1 0 0 9 0 9 2
41 11 11 1 11 2 15 1 10 9 13 10 9 0 2 13 0 9 12 13 1 9 1 9 9 11 1 11 9 2 12 3 2 16 16 1 10 9 13 11 12 2
26 11 1 11 0 9 2 12 1 9 0 9 7 11 1 11 0 9 2 12 1 9 0 9 1 9 2
29 3 15 13 2 16 9 1 9 0 9 4 13 9 11 0 9 2 12 7 10 0 9 9 4 3 13 16 9 2
24 0 0 9 11 1 11 2 0 9 11 1 11 2 0 1 9 9 2 12 2 4 9 13 2
5 9 9 11 1 11
14 9 9 13 9 1 9 11 1 11 2 9 0 9 2
19 3 9 2 12 13 9 0 9 1 9 11 1 11 2 3 9 2 12 2
17 7 4 1 9 9 13 12 2 12 2 12 9 1 9 10 9 2
16 13 9 13 0 3 9 0 2 9 9 11 11 7 0 9 2
20 1 9 0 15 13 9 11 11 1 9 2 0 9 2 9 11 11 1 11 2
51 1 9 13 0 9 2 11 11 1 11 2 0 9 0 9 1 0 9 0 2 0 9 0 9 7 9 9 11 12 2 2 9 2 11 11 2 9 2 11 11 11 2 9 11 11 11 7 9 11 11 2
22 9 13 9 7 9 13 2 16 3 13 2 16 1 9 0 9 4 13 11 1 11 2
40 1 9 0 9 4 13 9 9 7 1 9 1 12 9 2 14 12 9 2 4 13 9 0 9 2 0 10 9 0 7 0 9 7 0 9 0 9 1 9 2
26 1 9 13 9 2 11 7 13 3 9 1 0 9 1 9 0 1 0 9 7 1 9 0 1 9 2
9 0 13 2 16 9 3 4 13 2
25 9 1 0 9 13 0 9 2 9 0 9 13 13 2 0 9 13 7 3 1 9 13 0 9 2
4 9 13 13 2
15 9 2 11 13 9 1 0 9 7 13 1 9 0 9 2
9 9 15 13 1 9 0 0 9 2
16 1 9 0 9 13 1 9 3 1 9 7 0 9 0 9 2
26 9 2 11 7 9 11 13 9 10 9 1 12 9 7 13 0 9 2 10 9 1 9 13 3 3 2
40 9 2 11 1 11 16 0 9 13 2 16 9 13 15 7 16 9 2 15 13 1 9 2 2 1 10 9 2 9 2 9 2 9 7 0 9 2 13 9 2
27 13 2 16 9 2 15 3 1 9 13 9 2 15 13 13 1 10 9 9 7 9 9 0 2 7 0 2
8 3 13 7 0 9 7 9 2
23 1 9 9 4 9 13 1 0 9 7 9 2 9 2 1 0 9 7 3 13 1 9 2
20 9 7 9 4 13 9 0 7 9 9 2 11 7 9 4 13 3 1 9 2
26 1 12 9 2 12 2 12 2 12 2 4 9 3 13 7 1 9 12 9 7 0 0 9 3 13 2
26 9 11 1 11 4 3 13 7 9 12 2 12 2 12 3 13 1 0 9 7 13 3 1 0 9 2
16 15 4 13 3 1 0 9 2 15 4 13 7 13 1 9 2
8 15 4 13 7 13 0 9 2
14 3 2 9 2 4 13 3 1 9 1 9 9 0 2
2 11 2
28 9 2 12 4 9 2 9 2 13 1 0 9 9 12 9 12 9 7 10 9 13 1 9 7 1 15 13 2
17 12 2 12 2 12 4 11 1 11 13 9 11 12 2 1 0 2
10 0 9 15 13 9 11 1 11 3 2
7 0 9 4 13 0 9 2
18 9 12 2 12 2 12 4 9 3 13 7 4 13 2 16 4 13 2
14 9 12 2 12 2 12 4 3 13 7 2 9 2 2
25 16 4 13 1 9 2 13 0 2 0 9 2 7 1 12 5 12 9 13 7 1 12 9 13 2
10 3 4 2 9 2 13 14 12 9 2
14 9 10 0 9 1 9 9 2 12 4 13 16 9 2
10 3 12 2 12 12 13 9 9 12 2
6 11 1 11 1 0 2
19 1 9 9 11 12 2 4 13 0 9 1 9 0 9 1 9 9 0 2
3 11 11 2
16 1 0 9 2 12 2 12 2 4 13 0 9 9 7 9 2
31 0 9 4 13 7 13 1 0 9 2 3 13 2 0 9 13 7 13 1 0 9 2 15 4 13 1 0 9 1 9 2
17 1 0 9 4 9 1 9 15 13 7 4 13 9 9 16 9 2
20 3 7 9 2 9 2 4 9 2 12 13 9 9 2 9 2 11 2 11 2
56 1 0 9 0 9 7 9 0 2 11 11 4 9 12 2 12 2 12 1 9 9 9 9 2 11 11 2 0 9 0 2 9 1 9 13 2 9 9 13 7 0 9 9 13 0 9 0 9 1 11 1 9 7 0 9 2
15 9 12 2 12 12 4 0 9 13 0 9 9 7 9 2
17 12 2 12 2 12 4 9 3 13 1 0 9 0 9 7 13 2
5 0 9 11 1 11
5 13 3 0 9 2
17 0 0 9 1 12 2 9 12 2 9 4 13 1 0 0 9 2
10 10 9 4 13 14 1 0 9 9 2
29 9 4 13 0 9 2 9 0 9 2 9 2 7 9 7 4 13 7 13 1 0 9 1 9 1 0 9 2 2
12 1 0 9 4 13 9 1 0 9 0 9 2
20 1 0 0 9 4 13 0 9 2 9 7 0 9 0 0 7 0 0 9 2
18 0 9 11 1 11 13 0 0 9 2 12 9 0 2 7 0 9 2
21 0 9 13 3 0 2 0 2 0 7 13 0 9 9 2 14 12 9 12 2 2
37 1 9 13 1 9 9 2 15 13 0 1 9 9 2 7 9 0 9 1 0 9 0 9 2 0 0 9 0 9 7 10 9 4 13 3 3 2
11 7 13 9 0 13 9 1 0 0 9 2
6 9 9 13 3 0 2
10 9 13 0 1 0 7 3 0 9 2
11 1 0 7 0 9 4 3 13 0 9 2
20 9 13 3 0 2 3 0 2 9 0 7 0 7 0 9 4 14 3 13 2
14 12 9 13 3 0 7 3 0 0 9 13 0 9 2
9 0 9 13 9 9 11 1 11 2
51 10 9 4 13 2 1 9 9 0 0 9 2 1 9 9 0 9 12 9 2 1 9 9 9 2 1 9 9 0 9 1 9 0 7 0 7 1 3 0 9 0 1 9 2 1 9 12 2 12 9 2
19 15 13 2 16 9 9 11 1 11 13 0 13 1 9 1 9 2 12 2
6 10 0 9 13 0 2
15 1 9 4 13 14 9 3 0 1 9 1 9 0 9 2
25 9 13 0 14 1 0 9 1 9 3 1 0 9 7 12 0 9 3 2 1 15 13 1 0 2
4 9 11 1 11
15 9 9 11 1 11 13 3 0 9 9 2 3 0 9 2
32 9 9 13 1 9 7 3 1 9 14 1 9 9 9 2 7 7 9 0 2 1 9 1 0 7 0 9 0 7 1 9 2
19 10 9 13 13 9 0 2 13 7 13 7 9 0 9 9 0 1 9 2
21 9 11 1 11 4 13 1 11 7 13 14 1 12 9 1 12 9 1 0 9 2
18 1 15 13 1 9 3 0 13 2 16 1 9 4 13 3 0 9 2
18 1 9 13 0 0 9 2 15 13 9 1 12 7 12 9 1 9 2
36 1 9 2 16 9 13 3 0 2 16 1 9 7 0 2 1 15 13 9 1 9 9 2 0 9 9 0 1 9 13 9 1 9 3 3 2
3 9 0 9
31 9 0 1 3 16 12 9 4 3 13 9 9 7 0 9 2 15 1 0 9 13 7 13 15 1 0 9 2 1 9 2
25 13 3 13 7 2 16 1 9 9 7 9 9 13 11 1 11 9 0 9 1 9 7 9 9 2
9 13 7 2 16 9 1 9 13 2
16 1 9 1 9 7 3 1 9 9 4 9 13 10 0 9 2
5 2 9 2 0 2
2 11 11
28 1 0 2 0 9 0 9 11 1 11 4 12 2 12 2 12 13 13 7 13 7 9 0 2 2 9 0 2
11 11 11 2 0 1 0 9 1 0 9 2
61 9 0 1 9 4 12 2 12 2 12 3 13 7 9 13 9 2 9 2 9 2 11 2 11 2 9 2 2 9 9 2 11 2 11 2 9 2 2 9 2 9 2 11 2 11 2 9 2 2 9 2 9 2 9 2 11 2 11 7 9 2
19 1 9 4 9 9 13 1 0 9 7 13 4 15 1 0 9 7 9 2
42 0 9 4 13 1 9 9 9 11 1 11 9 2 11 7 9 2 11 2 11 2 0 7 0 9 1 9 1 0 9 9 11 1 11 9 2 9 2 11 2 11 2
21 0 0 9 1 9 9 11 4 13 12 2 12 2 12 2 16 4 13 9 9 2
30 9 12 2 12 2 12 4 0 7 0 9 9 13 3 9 0 9 7 13 3 1 0 9 7 15 13 1 12 9 2
42 9 9 9 1 0 9 11 1 11 13 0 9 0 0 9 7 0 1 9 9 7 1 0 9 0 0 1 9 9 1 9 1 9 7 0 1 0 9 11 1 11 2
14 9 0 0 9 1 9 11 1 11 13 13 0 9 2
8 1 10 9 13 1 0 9 2
24 1 9 7 9 2 3 9 0 13 13 1 0 9 7 1 3 0 9 2 13 15 9 0 2
35 13 3 13 2 16 1 9 0 9 11 1 11 15 13 0 9 2 0 9 0 9 9 2 7 2 9 9 2 10 9 2 9 7 9 2
11 9 7 9 0 7 0 9 0 9 0 2
34 11 11 13 9 12 2 9 9 9 12 1 10 9 11 9 11 2 9 0 2 1 9 12 2 9 9 9 15 0 9 11 11 12 2
1 9
5 13 1 0 9 12
7 11 11 2 2 11 11 12
9 9 1 9 9 1 11 7 1 11
6 11 11 2 11 11 12
6 9 2 9 9 7 9
3 11 11 12
3 0 9 13
3 11 11 12
1 9
3 11 11 12
7 9 2 0 9 7 9 9
3 11 11 12
4 9 0 0 9
3 11 11 12
2 0 9
3 11 11 12
4 0 9 0 2
2 11 11
3 11 9 12
4 1 0 9 9
3 11 11 12
4 1 9 9 12
3 9 7 9
8 1 0 7 0 9 9 9 12
3 1 9 9
5 7 0 9 11 12
1 9
4 1 9 0 9
12 11 2 11 2 11 2 11 2 11 2 11 2
4 11 2 11 12
3 9 1 9
1 9
4 9 0 9 12
3 9 9 12
5 9 10 9 12 2
1 12
4 9 1 9 12
5 13 4 1 9 12
1 9
6 9 13 9 1 9 2
8 3 0 0 9 1 0 11 2
6 0 9 1 0 11 2
7 1 0 9 1 0 9 2
6 0 9 1 9 9 2
7 0 9 7 0 9 9 2
6 9 0 0 9 13 9
2 0 9
2 9 12
2 0 9
2 11 11
3 9 9 12
2 9 12
1 12
3 11 11 2
6 11 11 2 9 9 12
7 3 0 0 9 1 0 11
22 0 0 0 9 13 1 9 12 1 0 11 7 4 13 1 9 12 2 12 9 9 2
15 9 0 9 1 9 1 12 9 9 7 3 13 9 9 2
21 1 0 9 11 13 10 0 9 1 3 0 9 1 9 1 12 7 12 9 9 2
50 13 3 3 9 11 1 11 2 9 9 1 0 11 2 1 0 11 2 1 11 7 3 7 0 9 1 11 2 3 11 2 11 13 0 9 1 9 0 1 9 11 2 11 2 3 0 16 12 9 2
44 11 2 11 2 11 1 10 9 13 9 12 0 9 1 9 9 11 9 2 1 11 1 0 11 2 15 1 9 0 0 9 13 1 0 9 2 7 2 14 1 12 9 9 2
24 9 3 13 13 0 0 9 2 7 3 15 13 2 0 11 12 2 12 2 12 2 12 2 2
2 11 11
7 9 13 9 1 9 9 9
55 0 9 9 11 2 11 7 11 11 11 2 11 9 2 11 2 1 9 1 9 1 9 0 9 13 7 1 9 1 9 13 0 9 2 15 13 0 13 9 1 9 9 9 2 9 9 2 11 12 2 12 2 12 2 2
22 13 1 0 9 2 15 15 3 13 1 0 9 9 12 0 9 12 9 9 9 9 2
24 3 3 4 13 2 16 9 9 12 2 9 0 12 9 2 13 9 3 0 9 0 9 9 2
27 9 2 15 4 10 9 13 7 1 15 1 12 9 3 13 9 9 9 9 2 13 13 1 9 10 9 2
20 1 9 4 13 3 9 2 15 0 9 13 12 9 1 9 9 9 9 9 2
29 16 13 10 9 0 14 1 0 9 9 9 2 9 13 2 16 13 13 9 9 1 9 9 12 1 0 0 9 2
8 15 4 13 9 9 1 9 2
51 9 15 13 2 16 0 9 1 9 9 12 4 13 4 13 3 2 9 7 0 0 9 2 1 15 13 1 9 9 9 2 0 2 7 0 2 11 2 12 2 12 2 9 2 12 2 9 2 12 2 2
2 11 11
4 1 0 9 9
2 11 11
21 9 2 0 9 0 9 2 15 15 3 3 13 2 15 3 13 7 15 1 15 2
11 9 10 9 13 0 9 1 9 0 9 2
50 0 15 13 10 3 0 9 2 16 9 13 0 14 3 2 13 2 14 0 2 9 12 2 12 2 12 2 12 2 9 12 2 12 2 12 2 12 2 9 12 2 12 2 12 2 12 0 2 2 2
63 9 9 13 12 1 0 9 9 12 2 9 2 0 9 0 2 0 9 2 0 9 9 2 1 9 2 12 2 7 11 11 2 11 2 0 2 12 2 12 2 12 1 11 2 2 1 9 2 12 9 1 0 11 1 11 2 13 12 1 10 0 9 2
27 16 0 9 13 3 3 3 7 3 2 13 0 0 9 2 0 2 0 9 2 13 1 9 1 0 9 2
42 0 0 9 13 13 1 9 2 9 9 2 2 12 2 2 1 2 0 9 7 10 9 2 2 12 2 2 2 9 9 2 12 2 1 2 0 9 2 2 12 2 2
46 1 9 9 2 15 13 9 2 7 13 3 0 2 13 1 9 9 2 13 15 13 7 13 2 13 3 0 2 7 1 9 1 9 9 2 0 15 0 9 7 9 13 15 1 9 2
18 13 0 2 16 1 11 15 9 9 13 9 1 9 0 9 0 9 2
10 7 15 13 3 0 9 12 2 9 2
20 11 13 0 9 2 16 9 13 0 2 4 2 14 13 16 3 0 2 0 2
18 13 9 9 2 7 2 9 0 0 9 2 16 0 9 9 0 9 2
28 0 15 13 10 9 2 2 1 9 1 15 2 10 0 9 4 13 13 0 9 2 16 15 9 13 0 2 2
20 13 2 14 7 0 9 0 9 0 9 2 9 3 2 2 0 9 3 13 2
7 3 13 0 9 9 0 2
7 1 0 9 13 0 9 2
5 3 4 13 9 2
6 0 9 9 13 9 2
12 0 9 13 13 1 0 2 3 0 0 9 2
18 3 15 1 9 13 9 2 15 12 9 13 2 13 2 14 15 3 2
17 3 10 0 9 7 13 0 2 9 2 2 16 13 0 9 9 2
26 1 9 9 16 0 9 2 3 13 0 9 3 2 16 15 0 9 13 0 2 13 11 9 0 9 2
40 13 2 14 1 9 9 0 10 9 2 15 13 9 2 0 0 9 2 2 3 1 11 0 9 13 13 9 2 15 15 13 13 1 9 1 9 2 9 2 2
22 3 10 9 0 9 2 13 0 7 0 2 13 0 9 0 2 0 2 0 2 9 2
14 13 15 3 9 0 9 7 9 9 0 9 7 9 2
29 15 15 13 1 0 9 2 1 0 9 13 11 7 9 9 2 16 13 0 2 1 0 9 13 13 0 9 2 2
26 9 7 9 15 3 1 0 9 13 0 2 0 9 13 13 1 10 0 9 2 7 0 9 13 13 2
16 13 3 0 2 16 0 13 14 9 2 14 2 0 2 9 2
7 15 13 10 0 9 9 2
15 9 15 3 13 9 2 0 9 9 1 0 9 10 9 2
24 3 15 13 11 2 16 13 2 2 0 9 0 9 16 4 15 13 1 9 16 9 1 9 2
38 9 13 13 3 3 1 9 2 14 7 14 1 10 0 7 3 0 9 2 9 2 9 2 3 15 10 9 13 0 9 2 1 9 1 9 0 2 2
22 7 13 2 14 15 13 10 9 1 0 9 2 3 14 7 2 16 4 13 0 9 2
23 3 13 2 13 2 14 15 2 16 13 3 0 2 16 4 13 9 3 1 0 9 2 2
15 0 14 13 2 3 13 9 2 13 2 14 9 9 13 2
12 1 11 13 0 9 2 3 13 1 0 9 2
32 13 15 1 9 0 2 13 0 9 2 3 13 3 0 9 2 2 1 9 16 2 0 9 2 7 2 0 9 2 0 9 2
31 3 7 1 9 2 12 11 11 2 11 11 7 11 11 13 3 3 2 0 2 9 2 11 2 12 2 9 2 12 2 2
17 3 11 7 11 3 3 13 9 2 9 12 2 12 2 12 2 2
42 11 11 2 11 1 0 9 1 0 11 13 1 9 2 16 3 15 0 9 15 13 3 16 3 2 3 7 3 7 3 2 11 2 12 2 9 2 12 2 2 2 2
9 13 9 0 9 7 13 10 9 2
18 16 4 15 13 10 9 2 4 9 13 0 0 9 2 7 13 13 2
8 3 13 0 15 13 9 0 2
24 15 4 3 3 13 1 15 2 16 4 13 0 9 1 10 0 9 2 1 15 10 9 13 2
7 13 15 7 9 9 9 2
18 1 0 9 15 3 9 0 9 12 9 2 9 7 9 2 3 13 2
35 0 0 0 2 1 0 9 2 9 13 13 10 0 9 1 9 0 0 2 0 2 9 2 15 13 9 2 2 7 15 1 0 0 9 2
29 3 1 10 9 15 0 9 13 2 7 15 13 9 2 2 3 2 1 0 2 0 2 9 1 0 9 2 3 2
27 11 3 13 10 9 0 9 9 2 15 13 9 1 9 2 7 9 2 0 9 9 1 9 9 0 9 2
25 0 13 0 9 9 2 3 13 1 9 2 3 1 9 2 0 9 9 2 15 13 9 0 9 2
11 15 13 0 9 15 2 3 15 13 9 2
52 0 1 0 9 13 3 9 7 9 13 15 1 0 2 0 2 0 9 1 9 7 9 7 13 15 1 15 3 2 7 1 9 0 2 0 7 0 9 2 3 3 13 10 2 9 2 1 0 0 9 2 2
24 10 3 0 9 13 0 2 3 2 9 2 9 13 2 2 7 13 3 1 11 1 9 0 2
60 13 2 14 15 2 16 2 9 13 0 9 2 2 13 10 9 13 2 7 3 1 9 13 1 0 9 2 13 2 14 15 3 9 9 2 13 2 2 3 2 3 2 16 2 9 13 9 1 9 2 7 16 15 2 13 1 0 9 2 2
29 0 9 15 2 16 13 2 16 9 3 13 2 3 13 2 7 1 0 9 1 0 9 13 2 13 0 9 9 2
15 3 13 13 9 2 16 9 13 9 0 9 9 2 3 2
20 15 15 13 9 0 2 0 2 3 16 9 2 7 13 3 1 9 0 9 2
15 0 9 7 13 0 9 9 2 7 13 1 15 0 9 2
9 9 16 9 7 9 13 0 9 2
29 13 0 2 16 7 1 9 0 9 13 9 7 9 2 15 15 13 1 0 9 13 0 2 3 13 7 7 13 2
9 13 13 3 14 9 2 3 9 2
25 13 9 9 1 0 9 0 9 13 3 0 16 13 0 9 7 2 16 1 15 13 13 0 9 2
60 3 2 7 1 0 9 1 9 2 15 13 0 9 2 15 15 13 16 0 2 10 9 7 7 13 0 2 9 14 13 9 0 7 3 15 14 13 1 0 9 3 2 2 7 15 3 13 7 13 2 16 4 15 2 1 0 2 13 9 2
7 9 15 13 2 7 13 2
32 10 9 13 3 0 2 1 10 9 7 13 13 9 0 9 15 2 16 15 13 16 0 2 16 15 1 9 13 0 0 9 2
10 0 9 10 9 13 0 2 0 9 2
25 9 9 7 9 1 9 7 13 0 1 0 9 2 15 13 1 9 0 13 0 10 9 1 9 2
36 1 9 9 1 10 9 2 1 10 9 1 10 4 13 2 16 15 13 0 7 0 2 16 15 15 13 0 9 2 3 13 0 9 7 9 2
46 15 11 13 1 9 2 16 13 2 2 0 9 13 0 1 9 1 9 3 0 9 2 2 2 9 2 15 13 3 0 1 9 9 2 7 13 7 2 1 0 9 2 2 0 2 2
14 9 0 9 1 9 7 10 9 4 3 13 0 9 2
29 0 9 15 13 13 1 15 2 16 13 2 14 0 9 13 9 2 13 0 9 2 16 4 1 15 13 0 9 2
8 1 10 9 13 13 3 3 2
19 1 0 9 13 2 0 2 9 2 15 13 9 0 1 10 9 0 9 2
17 7 3 1 9 9 15 13 13 9 2 7 16 15 13 13 9 2
12 9 1 9 0 9 14 13 0 9 0 9 2
18 1 15 3 13 10 9 0 9 1 9 7 9 2 9 2 9 2 2
8 7 1 10 9 1 0 9 2
23 9 13 3 0 7 0 9 1 15 2 16 4 15 10 9 13 13 0 2 1 0 9 2
10 0 0 9 13 1 9 0 9 0 2
21 9 9 13 2 3 3 0 9 13 13 3 0 1 0 9 1 9 12 2 9 2
1 9
11 11 11 2 11 2 2 9 1 0 9 2
9 0 9 2 12 9 2 2 12 2
9 11 11 2 11 2 2 0 9 2
9 0 9 2 12 9 2 2 12 2
12 11 11 2 11 2 2 0 9 1 0 9 2
7 11 2 11 2 12 9 2
16 2 0 9 0 9 9 0 9 2 11 2 12 2 2 12 2
10 11 11 2 11 2 2 0 9 9 2
8 9 2 12 9 2 2 12 2
17 0 9 12 2 0 9 9 0 13 16 9 9 1 9 10 9 2
30 2 11 11 2 11 12 2 12 2 9 2 2 1 0 0 9 2 9 12 2 2 9 0 9 7 9 9 1 9 2
27 2 11 11 2 11 12 2 12 2 9 2 2 1 0 0 9 2 9 12 2 7 1 9 0 0 9 2
27 2 11 11 2 0 11 2 12 2 9 2 2 1 0 0 9 2 9 12 2 7 0 0 9 1 9 9
27 2 11 11 2 11 2 12 2 9 2 2 1 0 0 9 2 9 12 2 7 0 0 9 1 9 9 2
7 1 0 9 13 16 9 2
40 2 11 11 2 11 12 2 12 2 9 2 2 1 0 0 9 2 9 2 12 2 7 0 0 9 1 12 2 0 9 2 9 9 9 7 9 1 9 2 2
39 2 11 11 2 11 1 11 2 12 2 9 2 2 1 0 0 9 2 9 12 2 7 0 0 9 1 9 9 2 9 0 2 0 9 1 0 9 2 2
41 2 11 11 2 11 2 12 2 9 2 2 1 3 0 9 2 9 12 2 2 0 9 1 0 9 2 0 9 9 1 11 7 1 0 9 1 0 7 0 9 2
44 2 11 11 2 0 11 2 12 2 9 2 2 1 0 0 9 2 9 12 2 2 9 1 12 2 0 9 2 1 0 9 9 1 11 7 1 9 9 1 0 7 0 9 2
45 2 11 11 2 0 11 2 12 2 9 2 1 0 0 9 2 9 12 2 2 9 1 9 0 9 2 0 9 1 9 2 0 9 7 9 9 2 7 1 0 9 1 0 9 2
55 2 11 11 2 11 12 2 12 2 9 2 2 1 0 0 9 2 9 12 2 2 9 1 0 9 2 9 1 9 0 9 2 2 1 0 9 1 0 9 2 0 9 9 1 11 7 1 0 9 1 0 7 0 9 2
9 9 2 9 2 11 11 2 9 2
2 9 9
2 11 11
25 11 2 11 7 0 9 15 13 1 0 2 9 2 7 9 0 9 9 7 9 1 9 0 9 2
40 13 1 15 3 0 9 7 9 9 2 9 2 9 1 9 7 0 9 0 2 0 9 1 9 1 2 0 2 9 0 2 0 0 9 2 9 2 9 2 2
19 3 0 0 9 0 9 13 9 9 1 9 0 1 0 9 2 3 9 2
27 14 3 15 7 10 9 9 13 1 0 9 1 9 7 0 9 1 0 9 0 9 1 0 9 2 9 2
17 0 2 9 2 13 7 3 0 9 2 3 9 0 2 0 2 2
42 0 7 0 9 16 9 10 9 9 2 15 1 0 9 0 9 3 13 0 9 2 13 9 2 3 1 10 9 2 1 15 15 9 9 13 0 0 9 2 13 13 2
35 10 9 7 9 15 13 16 9 1 9 2 3 13 10 2 0 9 2 0 9 9 2 0 9 2 2 3 3 15 13 9 9 2 13 2
32 3 1 12 9 13 0 9 7 9 1 10 9 7 0 9 1 10 9 0 9 1 3 10 9 9 2 15 13 0 0 9 2
20 0 9 3 10 9 13 7 13 3 0 9 1 0 9 0 3 14 1 0 2
52 16 3 3 0 9 13 13 7 9 2 7 0 2 2 0 9 2 2 7 2 0 9 9 2 0 10 9 2 10 9 2 3 13 0 9 2 0 9 1 0 9 1 11 2 11 12 2 12 2 12 2 2
22 9 15 9 9 13 2 3 13 1 0 1 0 7 1 15 1 9 7 0 0 9 2
45 7 15 3 1 0 9 9 2 3 9 7 9 13 1 9 2 9 9 13 7 15 15 13 9 9 1 0 9 2 3 0 9 2 1 16 4 15 13 1 9 2 0 7 0 2
39 0 9 15 3 9 7 9 0 9 13 9 16 0 13 2 16 4 15 13 9 0 0 9 2 0 1 0 0 7 0 9 2 3 7 1 0 0 9 2
69 16 1 0 0 9 2 3 3 2 13 3 0 9 7 9 0 9 7 10 9 7 3 0 9 9 13 13 1 0 9 3 3 1 0 9 2 0 9 16 10 0 9 13 9 3 0 2 2 13 15 0 9 10 0 9 1 0 9 16 0 9 7 13 0 9 1 10 9 2
25 9 0 9 7 9 3 3 13 0 9 7 0 9 15 13 2 16 4 13 1 0 9 0 9 2
17 13 0 9 0 9 2 3 3 9 1 9 13 2 15 13 15 2
47 0 15 14 13 0 9 2 15 15 1 0 13 13 1 0 9 0 9 2 3 9 13 1 10 0 9 0 9 7 10 0 9 2 16 9 7 9 0 2 15 13 3 1 9 0 9 2
4 9 2 9 2
13 13 7 0 2 16 9 9 13 13 1 9 9 2
6 9 2 9 9 7 9
2 11 11
34 9 2 9 2 9 2 13 12 1 0 9 1 9 2 1 9 13 15 12 5 2 1 9 0 12 5 2 1 9 0 9 12 5 2
13 3 1 9 7 9 13 12 5 9 9 0 9 2
23 9 2 0 9 0 9 2 3 13 14 12 5 7 9 2 0 9 9 2 14 12 5 2
28 0 9 9 13 11 11 11 2 12 2 12 2 2 9 9 0 2 0 1 11 2 3 7 9 0 0 9 2
21 3 15 13 2 16 9 13 15 0 1 9 2 7 16 1 10 10 9 15 13 2
74 7 3 10 0 7 0 2 7 3 7 0 2 3 15 13 13 9 2 3 9 2 9 13 1 0 9 0 2 7 2 0 2 0 2 16 9 0 2 13 7 1 9 9 9 2 0 5 9 1 0 9 2 7 1 0 9 2 9 13 9 9 2 15 13 1 0 0 9 2 3 2 0 9 2
14 0 9 10 9 2 0 13 2 0 2 0 2 2 2
23 9 4 3 13 1 0 9 1 9 9 2 7 0 2 2 9 2 2 9 2 0 2 2
20 14 10 9 2 3 3 9 2 7 13 1 9 9 9 2 13 2 0 2 2
25 16 9 9 2 11 13 3 2 13 1 9 2 13 4 15 2 7 3 7 9 9 2 13 3 2
11 9 13 9 9 9 0 1 9 0 9 2
41 15 7 2 16 1 10 9 13 9 2 9 2 2 15 13 9 2 1 15 7 1 9 0 9 9 13 9 2 9 2 2 7 15 1 15 13 9 2 9 2 2
11 1 12 9 13 9 9 0 1 0 9 2
44 1 0 9 2 9 2 1 9 9 2 15 1 0 9 13 9 7 15 13 9 2 9 2 15 15 13 0 9 2 4 13 2 1 9 13 9 3 9 9 2 9 9 2 2
21 16 2 3 0 13 2 9 3 13 9 2 9 2 13 15 3 1 9 1 9 2
7 9 2 0 9 2 0 9
34 7 16 11 11 14 13 9 9 2 16 13 0 9 1 9 2 9 12 2 12 2 12 2 2 13 9 9 0 9 9 2 1 0 2
10 9 9 1 9 1 0 9 13 9 2
22 1 9 15 0 9 13 1 9 2 0 9 1 0 9 2 7 4 3 13 1 9 2
22 9 13 2 13 15 1 9 9 7 1 9 13 9 2 9 2 0 2 9 10 9 2
5 15 15 13 9 2
16 3 0 0 9 2 1 9 0 2 13 1 2 0 9 2 2
7 9 7 1 10 9 3 2
30 16 13 9 1 9 10 2 16 13 9 1 0 9 2 1 0 9 2 13 2 13 15 13 3 9 7 7 0 9 2
22 7 13 9 0 1 0 9 2 3 2 1 11 2 1 9 3 0 9 16 9 9 2
33 7 15 3 9 1 0 9 13 2 10 9 3 13 3 0 9 7 3 9 7 13 0 1 9 13 3 9 7 13 3 0 9 2
36 7 15 7 9 13 7 1 0 0 9 2 10 9 1 9 15 13 13 9 7 13 15 15 2 3 2 10 0 9 15 15 13 2 1 9 2
22 1 9 0 9 9 15 10 9 0 9 13 2 16 9 13 9 0 9 1 0 9 2
48 16 15 3 13 10 2 0 2 9 1 9 13 1 9 2 9 2 2 13 1 0 9 2 10 9 13 0 13 3 9 7 13 15 0 9 2 16 15 13 13 15 0 2 15 0 9 13 2
29 1 0 9 0 9 3 9 13 7 13 0 9 1 11 2 7 1 11 2 2 7 15 13 13 9 10 13 9 2
49 13 2 16 15 13 13 9 9 7 0 9 3 13 3 0 9 2 1 9 13 3 9 2 9 13 13 3 9 3 2 2 16 1 9 13 13 2 7 3 13 13 2 16 15 15 1 15 13 2
19 3 0 9 1 9 9 7 9 13 13 0 9 9 9 7 13 9 9 2
22 9 15 15 13 1 0 9 2 9 7 9 2 2 3 16 15 13 0 9 7 9 2
10 9 7 13 2 16 9 9 13 13 2
13 9 0 9 7 0 9 9 13 13 9 7 9 2
6 3 15 13 2 16 7
6 9 0 9 13 13 2
37 0 9 9 2 9 2 3 13 7 13 4 13 9 9 2 7 12 1 0 9 0 9 13 15 2 16 13 3 0 2 3 10 9 13 3 0 2
30 0 9 13 0 9 2 9 2 0 9 0 1 9 2 15 3 13 13 1 9 7 9 1 0 9 3 1 12 9 2
14 3 13 0 13 9 2 7 15 13 13 9 7 9 2
28 9 7 2 16 9 9 1 9 9 13 9 9 1 9 9 2 9 15 13 3 13 2 16 4 9 9 13 2
33 15 13 12 1 0 7 0 9 9 1 9 2 13 0 9 2 16 13 0 13 1 9 9 1 0 9 2 16 13 1 9 0 2
15 7 9 9 9 1 0 9 13 13 1 9 7 1 0 2
11 3 13 15 1 9 9 7 1 0 9 2
37 3 1 9 3 0 1 0 9 2 9 7 9 0 9 9 2 2 1 3 0 0 9 2 15 1 9 9 9 13 13 9 2 15 9 3 13 2
3 13 15 1
12 2 0 9 2 2 0 0 9 2 0 9 2
28 1 9 2 1 15 13 13 9 9 1 9 10 9 2 15 13 0 9 9 2 0 9 2 9 12 2 2 2
8 13 15 9 9 0 9 9 2
27 13 0 0 9 2 3 13 1 0 9 7 13 1 0 9 9 7 1 10 9 2 1 2 0 9 2 2
24 0 0 9 13 0 9 2 2 2 3 0 9 9 1 9 10 9 2 9 2 1 0 9 2
20 9 9 2 15 0 9 1 9 13 2 7 3 0 7 0 9 13 0 9 2
27 1 0 9 13 9 7 2 9 7 9 2 9 0 9 15 13 1 9 9 2 9 1 15 2 1 9 2
23 1 10 9 1 9 3 13 11 2 11 2 9 12 2 2 2 2 2 2 12 2 2 2
27 13 15 3 0 9 2 3 3 13 0 2 16 9 0 9 13 0 1 9 1 0 9 9 7 1 9 2
15 9 1 0 9 9 9 1 0 9 9 13 7 3 0 2
26 13 9 2 16 4 15 10 2 0 9 2 13 13 9 2 1 15 13 0 9 0 9 0 0 9 2
22 9 9 4 15 13 3 13 9 9 9 9 7 0 9 2 16 3 7 0 0 9 2
9 0 9 15 14 13 7 1 9 0
37 3 1 9 9 1 9 2 1 9 2 13 9 0 9 1 0 9 14 9 7 12 1 9 0 9 2 16 13 9 2 9 9 7 3 7 9 2
10 3 3 13 9 2 0 9 9 0 2
17 3 3 15 13 1 9 2 16 13 0 9 4 13 0 9 9 2
37 15 4 7 13 13 9 1 9 7 13 15 1 0 9 2 3 13 9 9 2 0 9 2 15 15 9 13 2 1 15 0 16 1 0 0 9 2
29 0 9 2 0 0 9 2 0 9 1 9 7 0 9 2 0 9 2 9 1 9 2 15 3 13 16 0 9 2
5 13 15 3 3 2
24 0 9 1 9 3 3 13 9 1 9 9 1 9 2 15 4 13 9 0 9 3 0 9 2
20 10 2 9 2 9 4 3 13 13 0 9 1 9 9 9 7 9 9 9 2
52 13 13 2 16 1 9 2 15 1 0 9 13 0 9 0 9 2 15 1 9 1 0 9 2 9 2 9 2 9 2 9 1 9 2 13 7 0 2 9 1 9 7 9 2 7 0 9 2 0 1 9 2
14 13 15 2 3 3 15 13 2 0 2 9 16 15 2
17 15 13 13 9 9 0 9 2 9 2 9 2 9 3 2 2 2
21 13 15 7 0 9 2 3 4 9 0 9 2 9 2 1 9 13 13 13 0 2
10 3 0 13 2 16 0 9 13 0 2
33 4 15 13 13 1 0 9 2 13 9 9 0 9 2 2 7 0 9 2 13 15 1 15 9 9 1 9 9 1 9 2 2 2
13 15 13 1 15 2 16 9 1 12 9 13 0 2
6 9 15 13 1 0 9
29 13 4 1 9 2 16 4 0 9 13 10 0 9 7 16 4 15 0 9 2 16 3 15 13 9 2 13 13 2
22 3 13 0 2 16 10 0 9 13 9 1 9 0 9 15 2 16 15 1 9 13 2
16 16 9 3 13 3 14 1 9 2 7 7 1 9 1 9 2
23 16 3 7 2 1 9 1 0 9 2 3 9 0 9 13 2 13 1 9 3 0 9 2
13 13 15 9 0 0 9 2 3 2 9 2 9 2
40 1 9 1 0 9 7 0 9 0 0 9 13 13 14 9 1 9 0 9 2 7 7 9 1 0 7 3 2 0 9 7 9 3 2 15 13 9 0 9 2
10 3 3 15 13 9 2 3 15 13 2
18 2 2 0 14 13 2 16 9 0 2 9 13 2 0 2 9 2 2
6 15 13 7 10 9 2
23 13 1 0 9 9 2 9 1 0 9 2 7 10 9 7 1 9 2 9 2 9 2 2
9 9 10 9 12 12 2 2 0 9
2 11 11
26 13 14 1 9 2 16 10 9 13 3 3 3 10 9 9 3 0 9 10 9 7 9 1 0 9 2
20 10 9 13 0 9 9 0 9 2 15 15 10 9 13 1 9 12 2 12 2
39 1 0 9 4 13 15 0 2 0 2 0 2 0 2 0 7 0 9 2 15 4 13 1 0 9 13 1 9 1 9 2 2 3 1 15 3 9 2 2
11 1 9 0 0 9 4 13 1 9 9 2
19 1 9 9 0 9 2 0 7 0 9 4 13 0 9 0 9 1 9 2
33 9 0 9 4 3 13 2 16 3 10 9 4 10 9 13 3 3 2 16 4 15 3 2 13 1 9 0 9 2 3 0 9 2
15 3 0 9 13 2 16 3 0 9 13 9 1 0 9 2
47 0 9 9 2 15 4 13 2 7 15 0 9 3 0 9 13 12 9 2 1 9 14 1 9 2 0 9 0 9 2 0 9 9 1 12 2 12 9 9 9 1 9 2 7 0 9 2
17 10 9 13 2 16 0 9 0 9 1 9 13 9 0 0 9 2
20 0 9 4 13 7 1 0 9 2 7 1 0 9 1 0 9 2 9 2 2
30 3 0 9 4 13 9 2 16 1 0 9 0 9 9 1 9 1 10 9 2 13 15 1 0 9 0 0 9 13 2
19 7 4 13 3 0 9 0 9 12 0 9 2 11 11 2 7 11 11 2
18 9 0 0 9 13 2 16 0 0 9 3 13 1 0 9 10 9 2
33 1 0 9 15 15 13 3 11 2 11 2 15 9 12 1 10 9 2 9 2 1 9 9 9 0 0 9 13 2 2 2 2 2
8 11 3 13 9 2 2 2 2
27 2 1 12 1 10 0 0 9 10 9 13 10 9 13 3 2 2 11 13 0 1 9 2 2 2 2 2
33 12 2 16 4 0 9 13 1 9 9 0 2 13 15 1 10 9 0 9 2 9 0 0 9 12 2 2 12 2 9 1 15 2
20 9 9 9 1 9 9 7 10 0 9 10 9 13 3 2 3 13 0 9 2
21 15 1 9 0 9 2 11 1 0 9 9 13 13 0 9 2 12 5 2 2 2
30 1 15 12 1 12 9 0 1 9 9 0 9 0 3 0 9 1 9 12 2 12 0 9 13 2 12 5 2 2 2
33 3 15 9 9 7 0 9 1 9 1 15 1 15 2 1 9 2 13 1 9 3 0 1 9 9 1 9 13 1 9 10 9 2
16 3 4 15 13 13 0 9 1 9 11 2 11 2 9 2 2
1 9
20 0 9 13 1 15 0 9 2 3 1 0 9 0 0 9 10 9 1 9 2
30 1 9 9 1 9 15 3 13 9 9 0 9 2 11 3 11 2 11 7 11 2 15 15 13 13 13 3 0 9 2
31 9 2 15 15 1 0 9 13 1 9 10 0 9 7 9 9 7 3 13 0 9 3 0 9 2 15 13 4 13 3 2
24 1 0 9 1 9 13 9 2 11 2 11 2 9 2 2 10 0 9 1 9 2 9 2 2
10 11 11 15 1 15 13 13 10 9 2
19 1 11 2 11 2 13 15 7 10 0 0 9 9 2 11 0 2 9 2
36 2 2 12 2 2 15 13 0 2 0 9 0 9 1 11 7 13 1 0 9 11 11 1 11 2 3 15 13 0 9 9 1 0 0 9 2
25 12 2 9 12 7 12 10 9 13 7 13 4 13 1 9 2 10 9 3 13 0 9 10 9 2
11 12 2 13 4 9 0 0 9 10 9 2
27 1 9 9 9 1 0 2 0 9 1 0 9 2 9 2 13 9 2 2 1 9 1 10 0 9 2 2
36 9 2 16 4 15 9 1 10 9 13 13 0 9 1 3 0 9 2 3 2 0 2 9 0 1 9 2 9 1 0 9 2 10 9 13 2
4 13 4 1 9
1 11
1 11
4 9 1 0 9
3 2 2 2
31 13 4 13 2 16 4 0 9 9 9 13 9 10 0 9 7 4 15 0 9 13 15 2 15 4 13 0 9 2 2 2
16 9 0 9 13 0 9 0 9 1 10 0 9 9 2 2 2
11 11 11 2 0 9 2 12 2 12 2 12
4 9 1 0 9
16 15 3 7 1 11 2 11 7 0 9 13 3 12 9 9 2
9 7 7 0 9 15 13 0 9 2
23 0 9 15 12 0 0 9 15 3 13 1 12 9 0 9 2 15 13 1 0 9 0 2
21 0 9 13 3 0 0 9 1 0 9 9 2 3 0 2 16 2 9 2 9 2
20 11 10 9 1 9 2 0 9 2 1 9 2 0 9 2 13 3 3 0 2
1 11
20 0 9 2 7 0 9 1 9 2 0 0 9 3 13 11 16 9 2 2 2
15 3 1 12 9 9 13 2 1 0 12 9 15 13 2 2
3 9 13 9
26 10 9 13 7 0 2 7 2 2 2 13 1 15 0 9 2 1 0 9 3 1 9 9 2 2 2
13 2 2 2 3 15 10 3 0 9 13 3 0 2
26 13 1 3 0 9 1 0 9 7 1 0 9 13 1 0 0 9 2 16 0 9 2 15 3 13 2
9 11 11 2 11 12 2 12 2 12
2 9 2
6 9 1 2 9 9 2
2 11 11
5 13 1 0 9 12
1 7
4 15 13 0 2
2 11 11
37 1 9 12 4 13 0 9 2 9 12 2 12 2 12 2 1 9 2 15 13 9 3 13 1 9 9 1 0 9 0 9 2 9 7 9 9 2
37 1 10 9 13 10 9 3 1 0 9 2 11 2 11 2 11 2 11 2 2 7 1 9 9 9 7 9 13 3 9 1 0 9 9 1 9 2
23 13 15 0 2 16 1 0 10 9 13 9 1 9 3 0 9 2 16 1 10 9 13 2
29 13 15 13 7 3 0 9 1 9 2 3 13 9 0 9 2 15 13 9 0 9 1 0 9 10 0 0 9 2
30 16 9 13 3 3 7 13 15 1 9 3 1 12 9 9 2 13 3 0 2 16 0 9 15 13 13 3 1 9 2
28 9 1 15 3 13 3 16 1 9 0 9 7 3 1 0 9 15 2 0 9 2 9 1 10 9 3 13 2
19 1 0 9 3 13 0 9 1 9 1 15 3 2 15 13 9 0 9 2
31 9 2 14 1 9 12 2 9 3 13 2 9 2 1 2 9 2 2 7 1 9 15 0 9 13 13 16 9 0 9 2
25 3 1 9 2 3 0 9 13 1 9 9 0 9 2 13 7 3 2 9 1 9 13 0 9 2
25 9 0 9 13 3 13 2 16 1 9 0 9 0 9 13 0 9 9 9 14 3 0 16 3 2
13 9 9 9 13 1 9 1 12 7 12 9 9 2
11 1 10 9 14 3 13 0 9 3 0 2
11 7 13 1 9 0 0 9 13 3 0 2
25 9 0 7 0 9 16 7 0 9 9 9 3 3 13 2 16 3 1 12 9 9 9 3 13 2
26 3 9 2 12 9 1 0 9 13 9 2 15 13 9 9 1 9 14 12 9 1 0 12 9 9 2
39 15 15 13 0 9 11 2 11 0 2 2 0 3 9 2 12 2 16 1 9 9 7 9 13 1 9 1 0 9 1 9 9 9 14 12 9 2 9 2
15 11 0 2 13 1 9 0 9 9 1 10 9 1 9 2
16 9 13 3 1 0 9 3 0 2 7 1 9 13 3 0 2
20 11 0 2 13 2 16 9 9 13 9 10 9 9 7 9 2 1 0 9 2
26 9 13 10 9 1 9 7 3 1 9 2 7 9 15 1 9 3 0 13 2 13 3 1 0 9 2
11 1 9 2 0 2 9 15 3 13 9 2
53 1 0 9 1 9 0 11 1 11 13 3 9 2 12 9 11 11 0 9 1 9 0 0 9 7 13 3 0 7 3 1 9 0 9 11 2 1 9 2 0 9 2 2 1 9 14 12 9 7 9 12 9 2
37 9 7 4 13 1 0 9 14 1 12 9 3 7 3 3 9 13 2 16 15 9 13 1 0 9 2 1 0 9 9 3 13 14 9 2 12 2
33 9 9 12 9 9 13 1 0 9 1 9 9 2 0 9 2 1 0 9 11 7 13 15 3 1 9 0 0 9 1 0 9 2
21 1 9 9 13 13 1 9 0 1 9 2 9 12 9 9 11 2 12 12 9 2
12 1 2 9 2 9 13 3 12 12 9 2 2
8 9 4 13 13 0 9 3 2
24 3 13 9 1 9 1 9 1 12 2 12 9 1 12 12 9 2 15 15 13 0 0 9 2
50 3 3 0 9 13 1 9 1 9 1 12 1 12 9 2 15 13 1 9 13 3 0 9 2 13 9 0 9 12 2 9 12 2 0 9 1 0 9 1 9 3 12 9 1 9 12 9 2 9 2
14 0 9 1 12 9 11 13 9 1 9 12 9 12 2
26 3 11 2 11 13 0 0 9 9 9 1 9 1 12 9 9 2 7 9 10 2 9 2 15 13 2
31 1 0 9 13 14 12 14 3 0 9 1 9 9 9 7 12 0 0 9 0 9 9 9 2 12 1 9 11 1 11 2
13 3 3 4 13 7 13 9 9 2 9 2 9 2
20 3 1 15 13 0 9 3 10 2 16 10 0 9 1 0 9 13 3 0 2
13 1 0 9 7 1 0 0 9 3 14 13 13 2
38 9 13 16 1 9 1 9 1 12 9 2 7 1 9 9 2 15 13 3 0 7 0 2 13 7 9 7 10 9 2 7 3 3 0 9 1 9 2
34 1 9 1 9 2 15 3 13 1 9 1 10 9 16 9 2 15 9 13 1 0 9 1 0 9 2 3 7 3 1 2 9 2 2
43 16 0 9 9 1 9 3 14 3 13 12 9 2 9 2 9 9 15 13 13 7 9 14 12 9 2 9 2 7 2 1 0 9 14 12 7 0 2 1 0 9 2 2
10 0 9 9 0 9 13 11 2 11 2
28 1 15 15 13 9 1 9 9 1 9 3 1 12 9 9 7 1 9 1 9 1 12 9 3 1 9 9 2
15 15 13 3 0 9 2 16 4 15 1 15 13 15 13 2
56 1 12 2 0 9 0 0 9 1 9 12 1 0 11 13 13 0 0 9 1 2 9 1 9 2 2 11 2 2 15 13 12 0 9 2 3 3 13 9 16 3 0 9 0 9 7 1 0 13 0 9 9 1 0 9 2
10 12 10 9 13 3 7 3 3 0 2
29 0 9 9 9 7 9 15 13 1 9 9 0 0 9 2 15 13 1 10 0 9 1 9 1 0 0 0 9 2
33 1 0 9 10 9 13 0 9 1 11 1 0 11 2 3 4 1 0 9 3 9 11 2 11 13 10 9 9 7 3 10 9 2
49 13 3 0 2 16 7 1 0 9 13 3 13 14 0 9 9 1 9 9 2 7 15 3 1 9 7 9 9 2 13 2 14 1 9 9 9 2 0 9 3 2 13 2 9 10 0 9 2 2
8 1 9 15 3 13 13 3 2
22 3 3 0 9 15 1 13 0 9 3 13 1 0 9 2 15 15 9 9 3 13 2
24 9 13 3 3 0 9 2 0 7 0 14 10 9 0 0 9 2 16 3 13 2 0 2 2
94 3 9 9 13 0 2 3 9 13 0 9 9 0 0 9 9 2 12 2 7 3 15 9 3 14 13 15 2 16 3 1 9 12 9 9 1 9 2 7 2 9 9 9 2 9 2 15 9 0 9 13 1 9 9 13 9 7 13 9 2 15 1 9 13 0 9 2 15 2 15 13 2 2 7 15 15 3 13 9 9 2 3 9 0 9 13 9 2 9 1 0 0 9 2
35 0 9 11 11 13 2 16 0 9 13 15 12 9 1 9 1 12 9 7 1 10 0 9 4 13 3 13 1 0 9 9 3 9 9 2
8 3 13 10 9 0 14 12 2
22 1 15 15 1 9 3 13 9 11 1 0 9 12 2 0 0 9 9 9 2 12 2
23 9 12 2 9 12 13 1 9 12 9 9 1 9 2 3 3 1 9 9 9 2 9 2
11 1 0 9 9 13 10 9 3 12 9 2
26 13 3 1 9 9 3 0 2 7 1 9 1 9 1 0 9 15 1 2 0 9 2 1 9 13 2
25 3 15 0 9 1 9 13 10 9 3 2 16 1 0 9 13 1 9 3 3 16 9 2 12 2
5 13 15 3 3 2
31 16 15 10 9 3 13 1 9 2 3 15 13 13 0 2 16 15 3 3 3 13 2 7 0 9 9 15 3 13 3 2
13 9 3 13 3 1 9 2 15 4 3 3 13 2
24 3 0 2 9 13 1 0 0 9 2 15 13 3 3 0 2 7 1 0 9 1 9 9 2
30 3 15 13 2 16 1 9 15 13 13 7 9 1 3 0 9 7 9 9 9 2 3 0 9 1 0 2 0 9 2
44 3 3 13 3 2 16 3 9 2 12 1 9 0 9 13 11 0 9 9 7 0 9 1 11 1 9 11 2 3 15 13 1 10 9 16 1 12 2 0 9 1 0 11 2
25 0 9 3 13 2 16 4 15 1 9 0 9 13 13 0 9 2 7 3 1 15 13 0 9 2
26 0 9 13 7 3 3 15 13 9 1 9 9 9 0 9 1 9 7 10 9 1 0 9 1 9 2
59 9 7 13 7 3 13 0 9 1 9 0 9 2 15 3 9 2 15 3 9 2 15 13 3 9 9 0 9 1 9 0 0 9 2 9 2 2 3 9 13 9 9 7 3 3 0 9 2 7 10 9 13 3 3 13 1 0 9 2
33 3 9 2 12 13 11 11 1 0 0 9 1 11 0 9 2 1 15 13 0 9 0 9 2 15 13 1 3 0 9 1 9 2
25 1 15 4 13 0 13 1 0 9 9 1 0 9 2 15 4 13 1 9 7 13 1 10 9 2
36 9 2 12 13 0 9 11 2 16 4 15 9 9 9 1 0 9 13 0 9 2 7 9 10 9 13 0 9 1 9 7 2 0 9 2 2
21 1 9 0 9 15 3 0 9 3 13 9 2 16 9 0 9 13 16 1 9 2
31 1 9 9 13 3 13 0 9 1 0 9 1 9 2 15 4 3 2 13 2 0 9 14 1 9 12 9 9 1 9 2
19 0 9 9 13 3 3 0 16 0 0 9 2 7 0 9 13 0 9 2
48 16 15 3 13 0 9 0 1 9 2 13 14 12 9 1 0 9 2 7 0 9 13 1 9 12 9 11 2 3 0 0 9 13 0 9 2 10 0 9 13 2 14 2 12 9 11 2 2
11 0 13 3 2 13 2 3 3 1 9 2
44 1 9 12 9 9 2 9 9 9 2 9 2 13 1 9 0 0 9 9 14 12 9 11 2 7 1 15 13 0 13 0 0 9 0 1 9 9 7 9 9 1 12 9 2
23 13 2 14 3 0 9 1 3 9 2 13 9 2 16 10 2 9 2 3 13 1 9 2
16 1 2 9 2 0 9 1 9 9 13 9 3 0 0 9 2
25 7 15 3 13 9 0 9 2 0 9 13 2 1 9 2 1 9 1 9 14 9 9 1 9 2
41 13 13 1 0 2 0 9 1 0 9 9 2 15 13 9 9 1 0 9 9 2 15 13 0 9 2 15 13 9 9 2 9 2 2 7 15 0 9 13 9 2
31 9 13 9 9 9 1 3 9 2 7 3 13 0 9 2 9 2 9 3 1 12 9 2 7 13 3 1 12 9 11 2
59 9 1 9 0 9 15 13 1 9 9 9 2 9 9 3 4 13 9 9 9 7 0 0 9 9 9 9 2 15 13 7 3 3 2 16 9 2 15 4 13 0 0 9 1 9 1 9 1 12 9 2 15 4 13 1 0 9 9 2
36 9 0 0 9 11 11 15 3 13 13 2 16 4 15 13 13 0 9 1 9 9 9 2 2 2 2 11 2 15 13 9 1 9 7 9 2
29 11 15 13 0 9 2 2 0 9 15 13 3 13 1 0 9 2 13 15 3 2 16 13 13 1 9 9 2 2
63 1 3 0 3 0 9 15 3 9 13 9 0 9 2 3 15 1 9 13 2 0 0 9 2 2 13 15 1 9 2 13 15 0 0 9 2 2 16 0 9 13 0 9 2 3 13 0 0 9 1 12 2 9 2 7 3 1 0 9 9 15 9 2
29 9 3 13 2 16 1 9 9 1 12 9 9 4 3 1 9 13 12 0 9 7 0 2 0 4 13 0 2 2
18 7 13 0 13 2 16 9 10 3 0 9 1 0 9 13 3 0 2
17 1 0 9 0 0 9 15 13 3 3 9 2 15 13 16 0 2
