118 17
24 11 2 12 2 13 16 9 0 9 2 0 9 0 9 7 0 9 2 15 13 9 12 9 2
8 9 13 7 16 0 0 9 2
13 15 13 15 12 9 9 2 15 13 15 9 3 2
30 16 11 12 9 9 11 1 13 2 3 13 9 9 0 11 9 7 13 11 15 9 1 2 13 2 15 9 11 13 2
5 0 9 13 9 9
9 9 3 13 2 16 12 9 13 2
12 11 3 9 11 11 13 9 11 0 9 11 2
26 2 15 4 13 2 15 2 11 9 9 9 2 13 2 3 11 11 11 7 11 2 2 13 11 3 2
21 11 13 3 13 2 16 11 13 3 12 9 9 7 13 11 0 9 1 9 13 2
2 11 9
16 2 3 13 15 15 9 2 15 4 13 2 2 13 11 3 2
7 15 9 13 3 0 9 2
11 1 12 9 4 4 9 13 12 9 9 2
6 11 4 9 3 13 2
21 15 9 2 15 9 13 9 2 4 3 0 13 2 7 0 13 15 3 3 13 2
9 0 11 13 11 9 15 9 9 2
5 11 13 9 9 2
7 11 13 9 1 9 1 2
5 11 13 9 1 2
6 7 0 13 9 3 2
6 11 13 1 0 9 2
11 0 9 9 1 13 12 12 0 9 9 2
8 9 1 13 15 15 0 9 2
8 0 9 4 3 9 3 13 2
5 11 13 11 3 2
9 9 12 12 13 9 1 9 3 2
5 9 13 3 0 2
10 15 9 13 0 9 1 3 1 9 2
6 9 13 15 9 13 2
6 9 1 13 0 9 2
5 13 9 15 9 2
6 11 13 15 3 9 2
8 0 9 13 11 0 0 9 2
5 11 13 9 3 2
4 9 13 9 2
7 9 1 13 15 9 9 2
6 15 9 13 15 1 2
8 15 9 13 15 9 1 3 2
9 15 13 11 9 1 15 1 9 2
5 9 13 9 13 2
6 9 13 16 0 9 2
6 12 9 13 9 9 2
6 0 9 13 0 9 2
6 9 13 9 1 9 2
4 13 9 3 2
6 11 13 9 0 9 2
5 15 13 15 3 2
4 13 9 9 2
5 11 13 9 1 2
4 13 9 9 2
11 15 4 9 1 13 9 12 7 12 8 2
9 15 0 9 13 3 0 9 9 2
8 3 13 9 7 9 15 3 2
5 13 1 9 9 2
5 13 9 9 9 2
6 9 13 0 9 3 2
4 13 9 9 2
5 0 9 13 9 2
5 15 13 15 0 2
8 15 4 3 3 9 9 13 2
7 15 13 15 9 1 3 2
4 15 13 3 2
3 13 9 2
6 15 13 0 9 9 2
7 9 13 9 9 9 1 2
5 15 4 13 9 2
9 3 13 1 9 15 9 0 9 2
7 13 15 9 3 1 9 2
5 13 3 15 9 2
5 13 11 9 1 2
5 13 0 9 3 2
6 9 13 11 0 9 2
4 9 13 3 2
5 13 0 9 9 2
4 9 13 9 2
6 13 9 1 9 9 2
7 9 13 3 3 9 9 2
8 3 9 1 13 15 15 3 2
5 9 13 9 3 2
6 11 13 3 3 3 2
4 9 13 9 2
7 11 13 9 9 9 1 2
9 9 13 9 1 9 1 9 9 2
5 9 13 9 9 2
5 9 7 9 13 2
6 9 13 9 9 15 2
7 11 13 9 9 9 13 2
5 9 13 0 9 2
8 9 13 9 9 1 9 9 2
5 11 13 9 9 2
4 9 13 0 2
5 9 13 9 9 2
6 9 13 15 9 15 2
7 9 13 9 9 9 13 2
6 9 13 1 12 9 2
8 9 13 9 9 1 9 9 2
6 9 13 9 9 9 2
6 9 13 1 9 9 2
6 9 13 9 3 9 2
5 9 13 9 9 2
6 11 13 9 9 1 2
4 13 0 9 2
6 9 13 9 3 9 2
6 11 13 9 3 0 2
7 9 13 1 9 9 1 2
5 9 13 9 9 2
7 9 9 13 3 9 9 2
5 9 13 1 9 2
6 11 13 11 0 9 2
6 9 13 9 9 1 2
3 13 9 2
7 11 13 9 9 1 13 2
8 9 13 9 1 9 9 13 2
7 9 13 9 9 1 9 2
6 11 13 9 1 9 2
9 9 13 9 1 9 7 9 1 2
4 15 13 9 1
14 9 14 13 3 16 14 12 13 15 16 15 13 16 2
