10148 11
5 9 2 13 4 13
3 1 9 9
13 3 13 1 9 2 16 9 7 9 13 0 9 2
11 9 9 13 1 15 2 16 9 9 13 2
3 13 9 2
5 11 9 2 0 9
22 0 9 9 2 15 3 13 2 1 10 9 15 9 7 0 9 13 13 2 3 13 2
41 1 9 1 12 2 12 2 12 4 13 9 0 9 0 9 1 9 2 9 12 12 2 2 0 9 0 2 9 12 12 2 7 0 9 0 2 9 12 12 2 2
12 1 15 13 9 9 13 9 9 9 1 9 2
14 9 9 0 9 13 3 0 7 1 9 13 9 0 2
12 9 13 9 9 1 0 9 7 1 0 9 2
10 1 0 9 13 13 9 13 1 9 2
36 9 2 16 9 2 7 9 2 9 13 15 2 15 4 13 9 2 4 13 9 13 1 9 2 0 9 13 2 7 1 15 1 9 13 9 2
6 9 13 0 0 9 2
7 9 9 9 0 9 1 5
5 0 12 2 12 5
4 12 2 12 5
5 0 12 2 12 5
4 12 2 12 5
5 0 9 0 7 0
9 9 1 12 9 9 12 2 12 5
4 12 2 12 5
8 1 12 9 9 12 2 12 5
4 12 2 12 5
9 2 0 9 9 1 9 13 2 2
21 9 4 13 4 1 9 0 0 9 0 9 13 2 9 2 9 2 0 9 2 2
31 1 0 9 15 9 9 1 9 13 2 15 13 1 9 1 9 9 2 12 2 12 9 2 1 9 9 2 3 1 9 2
21 9 12 2 15 13 9 13 9 1 0 9 2 9 7 9 7 13 9 10 9 2
22 9 12 2 0 9 9 9 0 2 0 2 0 2 2 2 3 2 9 1 9 9 2
16 9 12 2 1 15 13 0 0 9 3 13 1 9 0 9 2
50 9 9 15 13 3 9 12 0 9 2 9 9 12 2 12 9 2 2 2 3 15 13 2 16 0 9 13 13 0 2 2 2 9 2 9 2 9 7 9 2 13 13 1 9 7 13 0 0 9 2
12 0 13 9 2 16 4 9 4 1 15 13 2
7 9 10 9 13 13 9 2
5 11 11 2 9 11
3 9 2 12
7 9 2 9 2 11 11 12
4 9 9 2 9
10 0 9 2 2 11 12 2 9 2 12
10 9 2 2 9 2 12 5 12 5 12
6 9 2 2 9 2 12
2 9 2
4 9 1 9 2
8 9 7 9 3 13 0 9 2
10 9 0 9 14 12 0 12 0 9 2
10 0 9 0 9 7 9 1 0 9 2
3 9 9 2
11 9 0 9 9 1 0 9 2 9 2 2
3 0 9 2
5 9 9 16 9 2
5 9 9 0 9 2
5 0 9 0 9 2
2 9 2
12 0 9 9 13 1 9 1 10 9 3 0 2
22 10 9 13 3 9 2 15 13 3 2 7 1 9 1 9 7 3 13 0 0 9 2
1 9
4 9 1 0 9
20 9 11 15 13 0 9 12 0 9 0 9 1 0 9 9 1 0 9 11 2
26 0 9 4 1 9 9 1 0 9 13 1 12 9 2 1 0 9 15 13 7 0 9 7 0 9 2
3 11 1 11
18 1 0 9 11 2 15 13 1 9 0 9 2 13 0 9 11 11 2
19 3 15 13 9 12 0 9 11 12 11 2 3 13 4 13 0 12 9 2
16 9 9 11 13 1 11 3 0 9 1 0 9 11 12 11 2
12 1 9 9 13 3 11 3 1 9 1 11 2
17 12 9 3 4 13 4 13 7 1 0 9 0 9 11 11 12 2
17 0 9 11 13 9 11 2 7 16 9 13 1 12 1 12 9 2
2 0 9
12 3 1 10 9 13 0 9 11 11 13 9 2
19 3 4 13 9 13 1 0 7 0 9 12 12 9 0 9 1 0 9 2
17 9 9 13 2 16 15 0 9 13 1 12 9 13 1 0 9 2
16 7 13 3 13 3 1 9 9 7 0 0 9 1 0 9 2
13 0 15 3 13 1 9 0 0 9 1 0 9 2
15 0 9 4 13 0 9 11 11 2 0 10 9 1 11 2
4 9 2 0 9
3 9 1 9
20 7 1 15 13 9 1 9 9 1 9 2 7 15 1 15 0 9 1 9 2
14 0 9 2 15 15 13 13 0 9 2 13 13 9 2
24 9 2 15 15 13 1 0 9 9 2 13 9 0 9 0 9 7 9 3 1 0 9 3 2
18 9 15 13 13 7 3 7 15 13 0 9 9 1 0 9 1 11 2
19 7 16 15 13 9 7 1 0 9 2 13 13 0 9 3 15 9 13 2
7 12 1 15 13 0 9 2
11 1 0 9 1 12 9 13 0 0 9 2
23 13 15 1 9 7 16 15 13 12 1 9 12 9 2 13 15 15 10 9 1 0 9 2
25 0 0 9 7 0 9 9 2 7 7 0 9 2 13 2 16 15 13 1 15 0 2 1 9 2
10 3 1 9 9 13 10 9 0 9 2
19 1 9 3 2 16 4 13 10 9 2 1 0 9 4 15 13 0 9 2
7 9 9 15 13 3 0 2
19 3 12 2 9 13 1 9 9 2 0 9 2 10 9 9 7 0 9 2
13 13 15 3 12 2 14 0 9 1 9 9 13 2
7 0 13 0 7 0 9 2
4 11 11 2 11
14 0 9 0 1 10 9 13 1 0 9 7 0 9 2
11 4 3 12 3 13 1 9 1 12 9 2
27 13 14 9 2 15 4 13 1 10 0 9 2 7 7 15 2 1 15 15 9 2 9 2 13 16 9 2
3 1 0 9
10 0 11 13 1 0 9 14 12 9 2
8 15 13 9 0 7 15 0 2
5 3 3 13 11 2
5 1 9 7 9 2
22 15 13 9 2 15 9 13 15 0 2 0 9 11 11 2 15 13 3 1 9 9 2
16 9 1 10 7 0 9 13 1 0 7 3 0 9 0 9 2
13 9 9 13 1 10 9 3 10 0 9 9 9 2
12 10 0 9 3 13 9 2 3 13 3 0 2
15 1 0 9 0 9 15 13 7 15 2 15 13 9 9 2
20 0 9 1 15 2 15 1 9 9 13 2 4 13 13 9 15 1 7 1 2
19 1 15 13 2 16 13 1 9 9 2 1 0 7 0 9 9 12 9 2
4 9 1 9 2
12 3 13 0 2 0 9 2 1 0 0 9 2
18 10 3 13 0 9 2 13 2 9 2 16 4 13 13 1 10 9 2
12 1 9 1 0 9 0 9 15 13 0 9 2
3 11 11 2
5 9 2 7 9 2
8 0 9 13 9 0 16 9 9
9 1 9 13 0 9 1 0 9 2
48 1 9 2 3 4 1 15 13 1 9 9 2 12 2 12 0 9 2 13 10 9 9 12 9 9 2 13 0 0 9 2 9 13 2 9 9 15 13 1 0 3 16 12 1 3 16 12 2
27 1 0 9 15 7 13 1 9 0 9 1 9 1 11 11 2 15 15 13 13 1 12 9 1 9 11 2
2 11 11
17 9 1 0 9 2 15 15 13 1 9 2 7 13 3 3 0 2
2 9 9
26 9 1 9 1 9 9 9 9 7 9 0 9 2 15 4 13 9 1 9 2 15 13 1 9 3 2
16 15 15 13 7 9 2 9 13 3 9 9 1 12 9 9 2
16 0 9 1 0 9 12 0 9 15 3 13 1 12 7 3 2
22 3 11 13 1 9 12 3 12 0 9 7 3 1 9 1 0 9 13 14 12 9 2
12 0 9 1 0 9 13 0 9 12 9 9 2
13 3 13 9 9 2 15 7 13 0 9 3 3 2
25 16 0 0 9 13 13 3 14 9 11 1 9 9 7 0 9 1 0 9 1 9 11 2 11 2
11 3 15 13 9 2 16 11 15 3 13 2
10 3 15 13 9 2 16 11 13 9 2
3 9 1 9
6 3 13 15 1 9 2
12 0 9 13 0 9 2 15 13 13 3 9 2
20 3 3 13 3 1 9 9 2 16 15 9 13 7 13 15 13 1 0 9 2
13 13 15 9 11 2 7 13 15 9 1 0 9 2
19 1 9 4 15 13 1 11 7 1 9 1 0 9 4 13 3 11 11 2
8 13 1 9 2 12 2 12 2
6 11 1 11 1 12 9
5 9 0 0 9 11
3 9 1 9
2 0 9
3 12 2 9
3 12 2 9
4 2 0 9 2
4 13 15 9 2
6 13 2 15 3 13 2
10 13 15 15 2 16 0 9 13 3 2
8 13 15 0 10 9 0 9 2
9 13 3 1 15 13 9 0 9 2
7 10 9 13 1 10 9 2
3 9 7 9
18 13 1 9 0 9 2 10 9 13 1 9 0 9 1 11 0 9 2
19 1 9 12 4 13 1 9 9 2 9 2 0 2 9 1 0 9 9 2
22 15 9 13 9 9 1 9 2 0 9 1 9 13 1 15 14 0 9 10 0 9 2
7 15 9 9 1 9 13 2
48 9 1 9 9 12 9 2 12 13 2 16 9 2 15 13 0 9 3 1 9 9 1 9 2 13 0 15 13 16 9 9 2 16 0 9 10 9 1 9 9 7 1 15 13 9 0 9 2
32 15 7 13 2 16 4 9 9 13 12 9 1 12 9 2 7 16 4 10 9 1 9 9 7 0 9 10 9 13 0 9 2
21 1 15 9 9 2 1 1 15 2 16 15 4 13 1 0 9 2 4 13 9 2
23 13 0 1 0 9 2 3 3 3 2 16 4 15 13 1 0 9 2 13 15 9 9 2
4 11 11 2 11
2 3 2
19 9 3 13 2 7 7 13 2 9 2 15 15 1 9 9 1 9 13 2
10 7 1 0 4 3 13 9 9 0 2
31 1 0 9 4 15 3 13 1 15 9 2 15 1 9 9 13 3 2 13 2 16 0 1 15 4 13 0 13 1 9 2
2 11 11
20 9 2 0 12 2 12 12 11 12 2 9 2 2 2 12 2 12 12 12 2
4 0 9 13 9
5 13 15 1 9 2
4 9 13 0 9
5 13 13 0 9 2
7 3 0 0 9 13 9 2
6 12 12 9 13 9 2
11 9 12 7 12 9 1 9 13 1 9 2
12 9 9 2 0 9 2 9 7 9 13 0 2
2 11 11
8 1 9 9 13 3 1 0 2
9 9 7 9 9 15 13 1 9 2
7 15 15 13 13 1 9 2
13 13 1 9 2 1 15 15 13 10 9 1 9 2
3 13 15 9
14 3 0 0 9 13 10 9 9 0 9 3 0 9 2
25 3 3 13 3 3 2 3 15 3 1 9 9 13 2 7 15 13 10 0 9 2 13 10 9 2
9 16 13 13 7 1 11 7 11 2
15 1 9 1 9 11 11 1 11 9 13 12 7 3 9 2
13 1 11 12 2 12 9 2 1 11 1 9 3 2
10 9 9 9 1 9 7 9 13 0 2
13 1 9 9 11 15 0 9 1 9 0 9 13 2
13 1 0 9 9 7 9 15 3 13 9 0 9 2
7 9 13 1 9 0 11 2
4 9 13 0 2
8 1 11 13 10 9 3 0 2
23 11 11 2 9 0 9 9 7 9 2 13 9 1 0 9 9 9 1 11 10 0 9 2
7 7 1 11 15 3 13 2
4 15 7 9 2
12 9 15 3 13 1 9 2 16 15 3 13 2
15 7 15 7 1 0 9 2 15 10 9 13 2 0 13 2
2 13 15
9 1 9 13 9 9 7 9 3 2
7 6 2 3 9 0 11 2
4 14 3 9 2
3 13 9 2
7 10 9 13 12 12 9 2
21 2 7 13 13 7 12 12 2 1 11 15 9 13 1 12 1 12 12 9 2 2
7 7 9 15 13 1 9 2
12 9 9 2 0 9 2 13 9 7 9 9 2
6 13 0 9 7 14 2
4 13 7 13 2
11 3 15 13 2 1 10 9 9 13 3 2
9 9 13 0 9 2 13 13 9 2
18 3 13 2 13 9 2 7 3 12 9 1 9 15 13 0 2 9 2
12 10 9 13 9 7 9 9 2 13 9 11 2
20 13 3 2 16 13 0 13 9 12 9 0 7 0 9 1 9 1 12 9 2
4 13 15 9 2
8 9 9 13 3 13 1 9 2
16 10 9 13 9 2 1 15 13 9 0 13 2 0 2 9 2
12 3 15 13 1 9 9 2 15 13 1 9 2
10 9 2 9 2 9 2 9 2 9 2
15 9 15 13 3 1 9 9 7 13 0 9 7 0 9 2
12 13 15 0 9 7 3 13 15 3 0 9 2
14 9 9 13 13 1 9 3 0 7 9 13 3 13 2
4 13 3 13 2
14 10 0 9 13 13 3 3 9 7 13 0 9 9 2
3 9 15 13
4 13 13 9 2
13 1 10 12 9 13 3 0 2 15 13 1 9 2
9 13 15 3 13 7 9 3 13 2
10 3 15 3 13 9 2 3 1 11 2
14 13 3 0 2 1 0 9 2 1 0 9 1 9 2
10 9 12 9 13 3 14 1 12 9 2
5 3 13 15 0 2
14 0 9 2 14 12 9 1 9 2 13 13 3 0 2
5 9 13 12 9 2
15 16 15 13 9 13 9 7 13 9 9 2 13 12 12 2
6 1 15 13 9 9 2
9 7 13 0 9 9 7 9 9 2
9 3 4 13 1 10 9 1 9 2
18 9 1 11 2 11 7 0 9 13 9 1 9 7 13 15 1 9 2
7 13 1 9 1 12 9 2
13 1 15 15 9 13 1 9 7 1 9 13 9 2
7 13 1 9 1 12 9 2
4 9 13 3 2
21 10 9 2 1 15 9 13 2 13 9 1 9 1 12 9 1 9 12 12 9 2
10 9 13 0 2 13 3 1 9 9 2
25 1 9 15 3 13 9 2 13 0 9 2 12 2 9 1 9 2 12 2 2 12 9 1 2 2
11 15 13 3 2 15 13 1 9 7 9 2
3 9 1 9
12 9 13 2 16 12 2 12 5 9 13 9 2
8 1 9 13 9 13 15 9 2
8 15 13 1 9 2 16 13 2
37 9 13 1 12 12 2 9 1 9 15 13 1 12 2 12 5 9 2 2 0 9 9 1 12 12 2 9 12 12 2 12 9 7 9 12 12 2
11 9 9 13 13 14 12 5 1 0 9 2
34 13 15 0 9 0 1 9 9 2 0 9 2 9 9 1 9 2 0 9 1 9 2 9 0 9 9 2 9 1 9 7 0 9 2
8 9 15 1 0 9 9 13 2
6 13 0 2 16 13 2
2 13 13
7 9 1 11 13 12 9 2
8 13 15 1 9 12 12 9 2
3 13 9 2
12 1 0 11 13 9 2 7 10 9 3 13 2
9 1 9 9 13 3 9 13 9 2
7 9 1 9 9 13 0 2
6 1 0 9 9 13 2
17 7 0 9 13 0 9 7 9 9 2 15 3 3 15 0 13 2
13 1 9 0 9 13 1 9 3 9 0 1 9 2
4 15 13 11 2
19 1 11 13 13 9 0 9 13 1 12 9 2 15 13 14 12 9 9 2
10 9 11 13 13 3 16 12 9 9 2
12 0 9 4 13 1 9 15 9 12 9 9 2
18 16 4 9 1 9 13 2 13 4 13 12 9 1 9 9 12 9 2
19 16 15 1 0 9 13 12 9 2 13 15 1 9 9 3 1 12 9 2
4 13 9 13 2
6 13 10 9 3 0 2
4 3 3 14 2
6 0 9 13 3 9 2
20 3 15 3 1 9 13 12 2 12 5 9 1 9 1 9 0 9 9 9 2
9 1 9 9 13 3 13 12 9 2
2 0 11
10 1 10 9 15 13 1 3 0 9 2
27 0 9 2 9 9 2 0 9 9 2 9 9 1 9 2 13 15 0 9 7 3 0 0 9 2 3 2
12 9 13 12 9 2 3 4 15 13 3 9 2
8 9 12 9 13 12 9 9 2
16 1 9 9 13 9 12 9 9 2 15 4 13 9 0 9 2
6 3 13 10 9 0 2
11 9 2 11 11 2 0 11 2 12 1 11
3 9 9 9
5 15 15 9 13 2
4 15 13 0 9
22 1 9 9 1 9 9 1 0 9 9 13 2 1 9 1 0 0 9 9 2 9 2
13 13 4 1 15 3 1 9 9 2 12 2 12 2
20 1 15 0 2 15 1 9 10 0 9 13 2 13 13 9 9 9 0 9 2
132 9 9 2 12 2 12 9 2 2 1 9 1 9 9 1 12 9 2 12 1 9 2 0 9 0 1 0 9 2 15 13 9 1 0 9 1 12 10 9 7 9 1 0 9 7 1 0 0 9 1 12 9 2 12 9 9 2 12 2 12 9 2 2 15 13 0 9 16 10 0 9 2 9 13 0 7 0 9 2 13 0 0 7 0 9 9 3 3 0 7 10 9 0 0 9 1 10 9 13 10 0 0 9 2 12 2 9 2 12 9 2 7 3 1 9 2 15 13 0 7 0 9 2 13 9 9 9 9 1 9 9 2
35 9 0 9 13 1 0 9 9 0 9 1 9 9 2 12 2 12 9 2 12 5 9 2 1 0 12 5 7 1 0 9 12 5 9 2
1 9
59 0 9 1 9 1 9 0 9 1 9 9 13 7 9 9 13 1 9 2 1 15 9 13 3 1 9 0 12 9 0 1 9 2 1 15 15 13 9 1 9 9 7 3 9 13 1 10 9 9 1 9 0 9 1 9 0 0 9 2
28 9 0 9 15 13 3 9 0 7 0 0 9 2 3 0 9 2 2 0 0 7 0 9 2 3 9 2 2
21 0 9 1 9 9 13 0 13 1 9 9 2 9 2 1 9 2 3 1 9 2
1 9
40 9 9 9 9 1 9 9 13 1 12 2 9 12 2 3 13 9 9 9 2 12 2 12 9 2 2 1 9 1 9 2 15 13 9 1 9 1 9 9 2
114 9 12 9 2 12 0 9 9 2 12 2 12 9 2 13 2 16 9 9 2 12 2 12 9 2 15 13 7 1 9 9 9 9 2 12 2 12 9 2 1 9 9 9 0 1 12 9 2 12 9 9 2 12 2 12 9 2 2 15 13 0 13 1 10 9 2 16 9 2 15 9 13 2 13 0 13 12 3 0 9 7 15 7 1 9 2 3 3 13 1 9 9 9 2 12 2 12 9 2 2 1 9 1 9 9 2 16 4 4 13 1 9 9 2
1 13
70 16 3 9 13 1 9 12 9 9 1 9 9 1 9 12 5 2 16 15 13 1 0 9 9 10 0 9 1 9 9 2 12 2 12 9 2 7 9 13 16 10 0 9 2 13 3 9 1 0 9 2 1 9 12 7 12 2 9 13 2 7 13 9 1 9 9 1 9 12 2
29 1 9 2 16 1 12 2 12 2 12 4 13 1 0 9 7 13 1 9 10 9 9 0 9 2 4 9 13 2
6 11 11 2 9 9 11
4 9 1 9 2
5 9 9 1 9 2
15 1 9 9 1 9 9 13 3 0 2 16 13 0 9 2
5 13 9 9 2 12
23 2 3 1 0 9 13 0 2 7 16 15 13 2 13 15 3 2 2 13 9 11 11 2
11 13 15 9 1 12 2 9 13 0 9 2
7 3 13 9 11 3 0 2
10 2 9 9 15 13 1 9 9 0 2
15 1 9 0 11 2 9 0 9 2 15 13 1 9 9 2
8 13 9 11 13 0 0 9 2
9 2 1 0 9 15 13 0 9 2
7 9 1 11 1 9 9 2
15 1 15 2 15 15 13 13 10 9 9 2 13 11 11 2
4 9 11 11 2
2 9 9
22 9 0 1 9 1 9 9 9 2 9 1 0 9 11 13 1 9 9 1 0 9 2
14 1 0 9 13 1 0 9 0 11 0 9 11 11 2
2 11 11
6 2 15 13 9 13 2
14 9 13 3 1 9 9 9 2 9 2 9 0 9 2
13 13 9 9 1 0 0 9 7 9 1 0 9 2
14 0 11 13 0 9 7 9 10 0 9 13 3 13 2
7 9 13 1 0 0 9 2
10 2 3 13 9 9 2 15 9 13 2
14 9 1 15 9 9 13 0 2 13 9 15 3 13 2
8 13 15 7 9 1 0 9 2
26 13 15 2 16 9 9 9 13 14 0 9 0 9 9 1 9 1 9 2 7 0 9 1 0 9 2
14 3 13 9 2 16 0 9 1 9 13 3 0 9 2
22 13 15 3 9 9 2 15 13 9 2 7 9 9 2 9 2 9 2 11 2 11 2
17 13 2 16 9 9 1 9 11 7 11 1 0 9 3 15 13 2
12 2 13 0 9 1 9 0 7 0 0 9 2
20 0 9 13 3 0 7 0 9 1 10 0 9 2 1 15 15 13 3 13 2
8 0 9 13 9 13 9 9 2
15 1 10 9 15 13 13 0 9 1 9 9 2 15 13 2
22 13 15 3 1 9 9 2 3 13 0 2 16 0 9 4 1 11 13 1 12 9 2
17 3 13 0 13 2 16 10 0 9 13 0 9 0 9 7 9 2
11 2 7 10 9 1 0 9 1 9 9 2
21 1 0 9 13 3 9 0 9 15 9 7 15 13 1 9 9 0 11 0 9 2
11 7 13 0 13 1 9 7 0 9 9 2
16 3 0 9 3 3 13 9 7 9 0 9 7 9 15 13 2
26 1 15 15 3 13 7 1 9 1 0 9 15 13 3 0 9 2 14 3 0 7 0 1 0 9 2
16 1 11 15 3 13 9 9 1 0 9 2 0 0 0 9 2
18 13 1 9 2 9 0 9 7 9 9 2 15 13 3 0 7 0 2
11 13 2 3 0 9 13 3 9 0 9 2
39 9 2 0 11 2 9 2 9 2 0 2 2 12 2 9 12 2 12 12 11 12 2 9 2 2 2 12 2 12 12 2 9 2 2 12 2 12 12 12
1 9
40 9 1 9 11 11 1 11 12 2 3 7 7 0 9 2 15 13 0 9 11 2 12 7 11 2 9 2 9 0 0 9 11 0 2 2 1 9 1 9 2
22 1 0 9 13 9 0 13 0 9 2 10 9 13 7 9 2 1 10 9 1 9 2
19 3 15 1 9 13 1 0 9 7 0 9 2 16 3 9 11 2 12 2
44 7 16 9 3 1 9 13 2 3 15 13 2 13 9 9 3 7 3 15 13 3 10 9 2 16 13 9 7 0 0 9 2 3 9 7 7 9 13 1 9 0 9 2 2
1 11
27 9 9 2 1 0 9 0 0 9 11 1 9 0 9 0 9 0 9 12 2 0 9 0 9 1 11 2
8 10 9 3 13 9 0 9 2
8 9 0 9 13 3 12 9 2
23 9 2 9 9 2 11 12 2 12 12 11 12 2 9 2 5 9 2 2 12 2 12 2
5 9 13 2 15 13
10 13 15 2 16 1 0 9 13 9 2
18 13 3 1 10 9 7 13 15 2 15 13 15 2 15 13 1 9 2
19 13 11 11 2 15 4 12 2 9 12 1 0 9 3 13 9 0 11 2
2 11 11
20 2 1 9 2 15 3 3 13 9 1 9 9 9 1 0 9 2 13 9 2
10 15 13 13 2 16 4 15 13 3 2
20 1 9 15 0 9 1 9 14 1 9 13 0 3 13 1 9 1 12 9 2
15 3 4 13 4 13 10 0 9 2 15 13 9 9 13 2
19 13 3 13 0 9 2 15 4 13 13 0 0 9 9 2 15 3 13 2
19 10 9 1 0 9 13 0 9 1 10 2 15 15 13 13 3 0 9 2
19 2 15 2 15 13 1 9 1 10 9 2 3 13 2 16 15 13 9 2
15 16 13 3 16 0 9 2 16 13 0 2 0 2 0 2
10 10 9 15 1 0 12 9 13 3 2
7 1 10 9 13 0 9 2
13 13 0 9 0 9 7 3 9 2 0 9 2 2
15 0 9 3 1 9 13 2 7 1 0 9 1 0 9 2
8 3 3 13 15 1 0 9 2
16 10 9 13 13 3 2 13 0 7 1 9 9 3 13 3 2
34 10 9 13 0 2 0 2 13 9 0 9 1 10 0 9 7 1 0 12 9 15 13 2 16 15 13 7 10 9 1 9 1 9 2
12 15 13 2 13 0 2 0 9 1 0 9 2
15 2 1 10 9 13 10 0 9 2 16 3 13 0 9 2
19 3 15 13 13 1 9 2 3 13 9 0 9 3 12 9 3 1 9 2
6 9 9 3 13 0 2
9 1 9 7 9 13 15 3 0 2
15 3 0 9 15 13 9 1 9 7 7 7 1 9 9 2
18 0 9 13 1 9 13 3 15 2 16 15 13 13 9 1 0 9 2
6 13 15 7 0 9 2
16 0 9 4 15 13 3 13 10 9 7 14 15 0 9 13 2
8 2 1 9 13 9 9 9 2
10 9 15 13 13 10 9 2 13 9 2
5 9 7 4 13 2
5 13 15 1 15 2
5 3 13 9 0 2
10 1 10 9 15 7 3 9 9 13 2
10 1 0 0 9 9 13 1 12 9 2
14 7 13 0 9 0 2 7 9 13 9 15 9 13 2
12 0 9 13 1 9 9 1 0 7 0 9 2
8 9 4 3 13 1 0 9 2
5 9 15 13 13 2
34 1 9 9 13 9 1 9 0 7 9 9 1 9 2 0 9 13 9 2 10 0 9 2 0 9 2 13 13 1 9 1 0 9 2
11 9 2 0 9 2 9 2 0 9 2 9
6 0 9 2 9 2 9
4 13 9 11 2
5 1 9 15 9 13
3 0 9 0
15 10 9 13 1 9 9 1 9 2 15 15 13 16 0 2
19 1 12 9 3 13 1 9 9 9 2 7 1 9 9 15 13 10 9 2
12 3 13 1 0 9 1 9 1 12 12 9 2
23 1 1 10 0 9 4 3 1 9 13 1 10 9 9 1 9 1 3 16 9 9 9 2
5 7 3 13 9 2
21 9 1 9 9 9 1 9 13 9 1 9 2 15 7 13 0 9 1 10 9 2
24 9 1 9 13 3 0 2 16 4 13 3 0 2 9 2 9 10 0 9 2 3 10 9 2
13 3 2 1 9 9 2 4 1 9 9 13 3 2
15 1 10 9 9 3 13 2 14 1 10 9 13 0 9 2
6 15 7 13 3 0 2
17 1 10 9 15 13 2 14 1 9 0 9 15 13 0 9 9 2
15 13 2 16 10 9 13 0 9 2 7 3 13 0 13 2
13 1 9 2 1 15 4 15 13 2 9 3 13 2
5 13 4 0 9 2
27 3 15 13 0 9 0 9 7 13 2 16 4 13 9 2 16 9 4 3 13 2 16 13 1 9 9 2
24 4 2 14 13 2 13 15 13 2 16 10 9 13 2 7 3 13 1 9 1 9 7 9 2
17 1 10 9 13 3 10 9 2 7 9 0 9 15 13 3 13 2
14 3 14 1 9 1 0 9 4 13 1 12 12 9 2
13 16 4 13 1 9 13 2 13 4 15 13 9 2
10 16 13 0 9 3 2 13 15 9 2
2 9 2
11 2 1 0 9 13 1 9 9 9 3 2
25 2 9 2 15 13 0 13 10 0 9 2 7 14 0 2 9 2 9 2 3 16 0 9 13 2
9 16 3 14 2 3 1 0 9 2
20 2 13 1 0 9 2 15 1 15 9 13 7 13 15 13 1 15 15 3 2
7 11 2 11 2 2 0 11
22 9 0 1 10 9 2 0 1 0 9 9 2 13 3 13 7 3 13 9 12 9 2
10 4 3 13 1 0 9 1 12 9 2
19 13 15 1 15 2 10 9 4 15 1 9 13 7 10 1 15 13 9 2
5 9 2 10 0 9
1 11
20 0 9 1 0 9 7 11 13 1 9 1 9 1 0 3 0 9 1 0 2
24 3 0 9 1 11 15 13 1 12 9 9 3 2 7 1 0 12 2 12 9 15 3 13 2
14 3 13 0 9 12 9 9 2 16 0 9 13 9 2
12 0 9 0 9 13 9 2 9 7 0 9 2
12 1 0 9 15 13 3 9 2 9 7 9 2
16 1 9 1 0 13 0 9 1 0 12 2 12 9 0 9 2
1 9
12 0 9 13 1 11 3 13 1 9 0 9 2
12 3 4 13 3 16 9 2 3 0 0 9 2
9 0 9 15 13 1 12 9 9 2
11 0 13 3 11 11 1 9 7 9 9 2
23 0 9 15 13 1 9 9 2 1 9 7 9 0 9 7 1 9 9 2 3 0 9 2
19 1 9 15 13 3 2 0 9 1 0 9 1 9 13 0 0 0 9 2
1 9
11 0 9 0 9 13 9 0 9 7 9 2
22 1 15 13 9 3 0 9 2 15 13 0 9 1 9 1 11 2 7 1 0 9 2
21 13 3 9 1 0 9 1 9 9 2 15 13 3 2 9 1 9 9 1 11 2
15 9 3 13 9 1 9 0 9 1 9 0 9 1 11 2
29 1 9 2 16 9 13 2 16 13 9 1 0 9 9 2 13 1 15 1 0 9 2 15 4 13 12 0 9 2
29 1 11 3 13 9 1 9 9 9 1 11 7 9 11 2 15 13 1 9 0 7 0 9 1 10 3 0 9 2
1 9
13 1 0 9 11 13 9 11 0 0 9 7 9 2
17 9 1 9 0 9 13 9 0 9 1 15 2 16 0 9 13 2
8 1 0 9 13 9 1 9 2
15 9 13 3 3 0 2 16 9 9 1 11 13 12 5 2
35 9 2 0 9 2 0 9 2 1 11 12 2 12 12 11 12 2 9 2 2 2 12 2 12 12 2 9 2 2 12 2 12 12 12 2
7 9 9 2 9 2 12 2
13 9 7 0 9 0 9 2 15 13 3 0 9 2
8 15 13 2 1 15 13 0 2
4 13 15 0 2
5 2 9 2 12 2
17 9 13 0 2 9 1 9 2 9 2 15 13 3 1 0 9 2
6 13 1 9 9 13 2
2 9 11
18 9 0 9 0 2 11 13 1 0 9 1 11 7 11 9 1 9 2
2 9 9
3 9 1 9
8 9 2 3 9 9 1 9 2
5 9 16 9 9 2
2 9 9
2 0 9
4 10 9 13 2
4 9 1 9 2
4 9 0 9 2
4 9 1 9 2
2 9 13
17 1 9 0 9 13 9 3 1 9 11 9 1 0 9 0 9 2
16 13 1 15 13 2 10 9 9 13 10 0 9 1 0 9 2
20 3 15 13 1 9 0 9 2 0 9 13 2 16 12 9 9 13 1 9 2
21 16 4 15 13 10 9 2 13 4 1 0 9 0 9 7 0 9 1 10 9 2
6 13 3 9 10 9 2
53 1 0 9 2 3 15 13 1 12 9 9 7 15 4 13 15 2 16 10 9 13 1 9 1 12 2 9 2 3 13 12 10 9 2 11 2 11 1 11 2 11 2 11 1 0 9 7 11 2 11 1 11 2
15 10 12 9 15 3 13 1 12 9 7 0 13 12 9 2
52 1 0 9 2 15 4 13 12 2 9 2 3 13 12 10 9 2 11 2 11 1 9 2 11 2 11 1 0 9 2 13 1 12 9 9 0 9 2 2 11 2 11 1 0 11 7 11 2 11 1 11 2
9 12 9 15 3 13 1 12 9 2
6 1 0 13 12 9 2
11 15 13 7 13 2 16 13 10 0 9 2
4 9 13 0 9
5 0 9 0 9 2
4 0 9 13 9
7 13 9 15 13 13 0 2
15 7 15 2 15 3 13 1 9 2 13 13 9 1 9 2
6 0 9 13 10 9 2
19 9 2 15 1 9 2 13 2 2 13 1 9 3 0 9 2 7 3 2
2 11 11
14 1 9 9 1 9 11 1 11 15 13 3 10 9 2
17 16 15 13 2 16 15 13 16 1 9 2 3 15 3 9 13 2
14 0 9 9 2 11 11 2 4 15 13 1 10 9 2
8 13 9 9 2 9 13 13 2
9 1 10 14 0 9 13 12 9 2
13 1 9 13 3 14 3 0 9 16 1 0 9 2
12 9 15 13 0 9 2 7 9 9 15 13 2
14 16 15 13 1 9 2 13 15 13 7 1 0 9 2
31 9 7 9 13 0 2 9 7 9 15 13 9 7 1 9 13 14 1 12 9 0 9 2 13 15 10 0 9 11 11 2
5 0 9 13 9 2
22 3 13 13 1 12 1 12 9 2 7 3 15 13 2 16 13 13 3 1 9 0 2
9 2 13 15 15 13 13 1 9 2
22 13 3 12 9 9 2 13 15 3 2 16 16 4 4 13 2 7 9 4 13 3 2
10 13 3 14 1 10 9 7 10 9 2
11 2 13 4 1 11 2 3 13 1 9 2
6 13 1 15 10 9 2
19 1 11 13 1 3 0 9 0 9 2 9 0 9 2 0 9 7 3 2
5 3 13 0 9 2
12 13 3 3 0 9 7 15 13 9 0 9 2
5 0 9 13 0 2
8 13 0 9 2 3 15 13 2
24 1 11 15 3 13 10 7 0 9 1 9 12 1 12 2 1 9 15 0 13 14 0 0 2
12 1 9 4 13 1 9 2 0 9 7 9 2
11 13 4 2 16 15 13 0 1 10 9 2
12 9 15 7 13 14 3 3 2 3 16 9 2
11 2 13 2 16 13 0 9 1 0 9 2
7 3 15 13 1 0 9 2
20 9 15 9 13 2 16 4 13 3 1 9 0 9 16 1 9 1 0 9 2
5 13 3 9 13 2
26 16 13 0 9 2 13 1 0 11 7 13 15 13 2 13 2 14 15 0 2 1 9 2 9 3 2
5 13 15 7 3 2
14 9 13 2 16 3 13 13 14 0 9 16 1 11 2
13 2 3 3 13 9 7 9 2 1 15 9 13 2
6 1 9 13 15 11 2
6 9 13 1 0 9 2
25 13 15 13 3 3 2 7 13 1 0 0 9 2 3 13 3 10 9 7 15 7 3 0 9 2
14 1 12 9 3 13 15 1 9 1 0 9 7 9 2
8 7 0 9 1 11 7 9 2
10 1 11 13 3 0 13 15 9 13 2
20 1 15 4 13 3 2 7 0 9 4 13 13 9 1 12 7 12 9 9 2
11 13 3 0 9 2 13 13 10 9 3 2
5 13 15 3 15 2
8 2 13 15 15 13 1 9 2
12 9 7 9 4 13 7 13 14 12 9 9 2
11 0 12 9 2 7 13 4 15 13 3 2
8 1 9 13 3 0 9 9 2
16 16 1 15 13 2 13 4 15 0 9 2 13 4 15 15 2
18 1 9 13 0 9 1 9 11 2 15 13 0 9 1 11 7 11 2
16 1 10 0 9 3 13 1 12 9 9 1 12 9 9 9 2
7 3 11 13 0 9 9 2
15 9 2 0 9 2 11 11 2 11 12 2 9 12 12 2
3 9 2 12
3 9 2 11
7 9 2 11 2 11 2 11
5 0 9 2 9 11
5 9 1 9 2 12
7 9 12 2 12 9 2 12
5 9 2 9 1 9
6 9 2 9 1 11 2
16 1 9 0 9 13 0 9 1 9 7 1 0 9 1 9 2
24 9 2 9 11 13 1 9 0 0 9 1 0 9 12 9 1 2 9 2 12 9 1 11 2
11 13 1 3 0 9 11 2 1 0 9 2
8 9 13 0 1 9 7 9 2
7 9 13 13 1 9 9 2
11 9 13 0 1 9 0 9 11 1 9 2
9 9 1 0 9 1 9 7 9 2
10 1 9 13 9 0 9 7 0 9 2
5 1 9 13 9 2
9 13 0 15 13 9 7 0 9 2
5 0 9 1 9 2
7 9 13 1 9 3 9 2
3 9 1 9
4 13 3 13 2
5 13 9 7 13 2
10 10 3 0 9 13 13 13 9 9 2
24 1 9 2 16 15 13 1 9 2 13 9 1 0 7 0 9 7 10 9 13 1 0 9 2
9 0 9 13 0 3 1 10 9 2
2 0 9
23 13 4 10 9 1 9 0 9 2 16 4 15 13 3 1 0 2 3 7 1 0 9 2
23 13 4 15 2 16 15 15 13 1 9 9 1 9 9 1 9 9 12 5 0 9 9 2
39 13 15 2 16 16 4 13 1 10 9 0 9 7 9 15 13 1 0 9 2 3 4 13 0 2 16 4 13 9 1 9 9 1 9 12 5 0 9 2
5 13 10 9 13 2
6 11 2 11 2 2 11
35 1 9 2 16 13 1 9 9 2 1 15 15 13 9 1 0 9 0 2 16 13 12 5 0 9 1 9 2 13 3 1 9 0 9 2
25 9 1 0 9 10 9 7 0 9 9 13 0 9 9 7 15 4 0 7 10 9 13 1 9 2
25 0 13 13 1 9 9 2 12 0 9 1 9 12 1 9 0 9 9 9 1 0 7 0 9 2
6 9 2 9 2 11 11
24 9 2 0 7 3 0 9 2 0 12 2 11 12 2 9 2 5 9 2 2 12 2 12 12
4 15 13 9 2
11 1 9 0 2 9 9 2 13 7 0 9
7 1 9 15 15 13 9 2
4 1 9 9 2
3 9 9 2
12 7 10 9 13 3 0 2 3 4 13 9 2
11 13 15 9 7 9 0 9 1 0 9 2
17 1 9 2 15 15 13 13 10 9 2 15 13 13 3 0 9 2
6 7 13 4 15 13 2
13 7 0 9 1 0 9 0 9 9 10 9 13 2
29 1 9 2 3 15 0 7 0 9 13 9 0 0 9 13 9 2 15 1 15 13 9 13 1 15 3 0 9 2
5 7 3 15 13 2
17 1 3 0 9 0 9 1 0 0 9 13 1 9 3 9 9 2
9 3 3 0 2 1 0 9 0 2
2 9 11
16 0 9 15 13 1 0 0 0 9 2 13 3 13 10 9 2
14 13 1 9 0 9 2 13 1 0 9 0 9 9 2
28 0 9 13 3 1 9 0 9 2 15 13 13 1 9 0 0 9 7 13 3 1 10 9 7 0 9 9 2
11 3 7 13 13 9 9 9 7 0 9 2
21 16 0 9 3 13 9 2 0 9 1 9 9 2 9 2 15 1 0 9 13 2
29 9 2 15 1 15 13 2 3 14 13 0 9 2 16 0 9 13 9 9 7 13 1 15 0 2 15 9 13 2
7 15 15 3 13 1 9 2
28 9 2 15 1 9 9 12 13 0 0 9 9 2 15 3 7 1 3 12 9 3 13 2 3 14 9 3 2
34 9 11 0 2 7 9 2 11 15 13 1 9 0 9 2 9 2 12 2 12 9 9 1 11 2 1 0 11 12 2 12 9 9 2
20 1 11 11 13 9 12 2 12 9 9 2 9 12 9 2 15 1 9 9 2
19 11 11 13 12 2 12 9 9 1 9 2 12 2 12 9 9 1 9 2
32 0 1 0 0 9 2 11 2 13 9 1 9 12 5 1 10 0 0 9 2 16 4 13 1 9 2 12 5 1 0 9 2
25 9 9 1 10 9 13 1 12 5 10 0 0 9 1 11 2 1 0 11 13 0 9 12 9 2
19 1 0 9 3 13 11 9 2 11 2 15 1 0 11 13 9 1 11 2
11 10 9 1 9 2 12 2 12 9 9 2
34 1 10 9 1 11 13 1 0 9 7 9 11 2 11 2 15 15 13 12 2 12 9 9 1 9 9 7 12 2 12 9 1 9 2
16 1 0 9 0 0 9 13 1 10 9 13 7 0 0 9 2
19 3 15 9 13 7 1 0 9 2 1 0 9 15 13 3 3 3 0 2
19 9 10 0 0 9 13 3 15 2 16 13 13 9 0 2 9 9 2 2
8 3 10 9 13 3 14 0 2
4 13 2 15 13
16 15 4 15 9 2 15 13 13 9 1 9 9 2 13 13 2
14 3 14 15 2 16 9 1 15 1 10 9 13 9 2
25 13 0 9 2 13 3 13 2 10 9 1 10 9 9 13 2 7 16 13 15 13 13 3 9 2
20 3 13 0 15 13 2 16 13 1 0 9 2 7 16 4 13 9 1 9 2
7 10 9 15 3 3 13 2
17 0 9 4 13 9 2 15 10 9 7 9 3 3 13 0 9 2
13 0 9 4 13 3 1 9 10 0 9 2 9 2
10 1 9 15 13 0 9 9 0 9 2
14 13 3 12 9 13 2 7 13 1 15 2 15 13 2
12 1 9 0 9 15 14 9 9 4 13 3 2
16 9 13 1 0 9 13 9 7 0 9 0 10 9 7 9 2
17 0 9 4 7 13 13 3 9 9 2 15 9 13 1 10 9 2
2 11 11
4 9 1 9 2
6 2 13 2 15 0 2
22 9 13 13 9 7 9 0 9 7 13 9 15 2 15 1 0 9 9 13 0 9 2
1 11
3 1 0 9
13 9 11 1 9 9 1 0 9 7 9 10 9 2
9 7 1 9 9 13 14 0 9 2
16 9 2 11 2 12 12 11 12 2 9 2 2 2 12 2 12
5 9 2 9 7 15
3 9 0 9
7 13 16 0 9 1 9 2
9 1 12 2 12 2 12 13 9 2
8 13 1 10 9 13 0 9 2
6 11 2 11 2 2 11
19 0 9 13 9 0 9 2 15 13 9 9 0 0 9 1 9 9 0 2
40 1 9 12 9 2 12 2 9 9 2 0 9 15 1 0 9 0 0 9 13 9 2 1 15 15 0 9 13 2 13 2 14 0 9 9 9 1 9 0 2
40 16 4 3 13 9 10 9 2 10 0 9 9 0 9 13 7 0 9 15 1 9 12 9 2 12 13 9 13 0 9 1 0 9 0 9 2 15 15 13 2
23 16 1 10 0 9 13 13 9 2 1 15 15 0 9 13 2 13 15 1 9 9 13 2
29 1 9 12 9 2 12 0 9 4 13 9 2 1 15 13 0 9 2 15 0 9 13 2 13 7 13 0 9 2
23 12 1 10 9 13 9 2 16 9 13 13 9 1 9 0 16 12 9 1 9 0 9 2
21 3 4 3 13 13 1 9 0 9 2 16 4 9 1 9 9 13 9 12 9 2
17 1 10 9 4 15 13 9 0 9 13 0 9 2 15 15 13 2
2 9 9
12 13 1 0 9 2 3 3 9 0 9 13 2
7 10 9 13 3 12 9 2
29 10 9 13 13 9 2 16 15 1 0 7 1 0 9 13 2 1 9 9 14 1 9 2 16 13 1 9 9 2
6 11 2 11 2 2 9
39 1 9 2 16 0 9 9 13 9 2 15 13 0 13 9 9 2 7 16 9 10 9 13 2 16 4 9 1 10 9 13 2 13 9 1 9 12 9 2
29 2 1 12 0 9 13 9 2 1 0 9 9 1 9 2 15 1 0 9 13 7 13 1 9 9 3 0 9 2
9 10 9 13 0 13 1 0 9 2
17 9 1 9 9 13 2 4 2 14 13 1 12 9 1 9 9 2
30 2 16 9 13 9 7 13 2 14 3 7 9 2 13 9 1 12 0 9 9 1 9 9 2 16 9 10 9 13 2
40 16 4 1 0 9 9 0 9 13 0 9 2 13 3 13 9 0 9 1 9 7 3 13 10 9 13 1 9 7 3 2 3 13 9 0 9 3 0 9 2
8 9 9 13 1 9 9 9 2
23 13 4 9 9 7 0 9 4 1 10 9 13 0 9 0 9 1 12 9 1 0 9 2
22 3 4 7 13 13 9 1 9 2 16 13 15 1 9 1 10 9 7 0 9 0 2
4 3 13 13 2
6 13 13 3 1 9 2
7 11 2 11 2 2 0 11
19 0 0 9 9 2 15 15 13 0 9 2 13 9 9 7 9 10 9 2
20 1 10 9 13 9 0 9 9 0 9 1 0 9 2 15 9 13 10 9 2
33 9 10 9 4 3 13 0 9 9 2 15 13 16 9 1 0 9 13 2 7 15 3 3 15 15 2 3 3 3 1 9 9 2
28 13 4 13 7 0 9 0 1 10 9 0 9 2 16 3 9 9 1 9 2 9 2 9 2 9 7 3 2
29 16 13 10 9 0 1 0 9 1 9 0 9 13 2 13 0 3 13 1 9 1 9 9 3 9 1 0 9 2
17 10 9 13 0 9 0 9 15 2 16 0 9 0 9 13 0 2
19 3 3 13 9 10 9 13 2 16 3 3 13 3 12 1 0 12 9 2
17 1 9 4 13 13 2 16 3 3 13 0 9 13 9 0 9 2
58 1 9 1 9 9 2 12 2 12 9 2 2 1 9 0 7 0 0 9 1 9 2 13 9 0 0 9 9 9 1 9 9 2 7 15 1 9 0 9 0 0 9 1 9 10 9 1 9 1 9 9 9 1 9 0 0 9 2
2 11 11
29 9 13 0 9 11 2 0 2 0 12 9 2 12 12 11 12 2 11 2 9 2 2 2 12 2 12 12 12 2
7 9 1 9 2 9 11 2
33 9 9 2 13 13 1 9 0 9 2 9 2 9 2 9 7 9 2 9 1 9 1 9 7 9 9 2 16 13 9 2 2 2
6 11 15 13 1 0 9
8 9 13 1 0 9 9 11 2
5 1 0 9 15 13
14 9 11 13 9 2 16 9 13 13 3 3 1 9 2
9 1 11 13 3 16 12 9 3 2
8 7 15 13 13 3 3 9 2
10 13 13 14 9 9 0 9 0 9 2
8 1 9 0 9 15 13 11 2
12 2 2 2 2 2 2 2 2 2 2 2 2
2 11 9
11 2 2 2 2 2 2 2 2 2 2 2
18 11 13 1 11 1 9 0 9 11 14 1 0 9 9 9 9 12 2
12 10 9 1 11 1 9 11 13 9 3 9 2
19 9 9 4 13 1 0 9 7 0 9 9 7 9 4 13 1 9 9 2
2 9 9
12 1 9 9 13 11 1 0 9 9 0 9 2
17 1 11 15 3 13 3 12 9 9 2 1 15 3 12 1 11 2
14 0 9 13 0 9 1 9 9 2 9 7 0 9 2
26 13 0 3 2 16 1 15 9 9 1 11 9 13 1 15 2 16 12 5 9 13 0 7 0 9 2
13 1 0 9 15 13 13 10 9 14 1 12 5 2
18 3 12 5 9 15 3 13 3 1 11 2 9 13 1 0 9 11 2
10 0 13 3 0 9 1 10 10 9 2
36 0 9 9 11 15 3 13 1 12 9 0 2 15 13 3 1 12 5 3 16 13 9 1 0 9 2 3 13 0 9 1 10 9 1 9 2
11 3 9 0 9 1 11 3 13 9 9 2
19 13 15 9 2 16 3 1 9 9 13 0 9 9 3 1 9 0 9 2
23 0 13 3 0 9 9 1 12 0 7 0 9 2 16 11 13 9 3 1 12 9 9 2
17 13 15 15 13 3 2 16 13 1 0 9 0 9 1 9 9 2
24 0 9 4 13 3 7 1 0 9 0 9 0 9 2 15 13 13 9 7 9 9 1 9 2
24 1 0 9 1 15 13 9 1 9 2 10 9 13 12 0 9 1 11 7 12 1 0 11 2
3 9 13 9
8 1 11 13 0 9 11 9 2
18 9 7 9 15 2 15 15 13 2 13 3 16 12 9 1 9 9 2
27 13 15 15 1 12 9 2 1 15 4 13 0 12 9 2 13 11 11 0 9 11 11 2 1 9 2 2
21 9 10 9 13 2 0 9 2 1 0 9 2 15 3 13 15 9 11 1 9 2
12 0 0 9 0 9 13 12 9 7 12 9 2
14 9 13 0 9 2 1 15 9 9 13 1 0 9 2
22 1 9 9 1 9 9 1 9 2 0 9 7 9 1 9 13 13 12 9 0 9 2
11 0 9 15 13 9 13 3 1 0 9 2
14 9 15 13 9 0 1 9 14 1 9 9 0 9 2
3 9 13 9
8 1 9 1 11 3 13 9 2
11 13 15 7 13 2 16 4 9 13 3 2
8 9 13 1 9 0 0 9 2
22 9 15 13 3 13 3 3 0 9 1 12 5 9 2 15 13 0 1 9 0 9 2
17 0 0 9 13 0 9 9 2 15 15 13 1 9 9 7 9 2
13 16 3 4 13 12 9 2 3 15 13 3 9 2
17 1 0 9 15 13 1 9 12 9 2 15 15 13 13 9 9 2
11 0 9 15 13 0 9 1 0 0 9 2
25 1 9 13 9 2 16 9 0 0 9 15 13 13 1 0 9 0 9 2 15 13 12 0 9 2
10 9 1 9 4 3 13 1 0 9 2
7 15 4 13 0 0 9 2
8 3 0 9 13 1 0 9 2
16 15 2 15 1 0 9 13 2 13 0 9 9 1 0 9 2
13 1 9 9 1 9 3 13 7 0 9 1 9 2
20 13 15 15 3 1 9 13 0 9 3 2 16 4 3 3 13 0 0 9 2
27 1 0 9 13 1 0 0 13 9 1 9 2 3 13 9 10 0 9 2 3 13 13 9 1 0 9 2
8 9 15 3 13 13 0 9 2
8 1 9 9 15 3 13 9 2
10 9 15 13 1 0 9 2 7 9 2
14 0 9 15 13 3 2 0 15 13 9 1 0 9 2
27 11 13 9 2 16 15 9 7 10 9 13 2 16 13 9 0 9 7 13 1 9 0 9 15 9 9 2
19 1 9 9 15 13 9 9 2 3 9 1 15 2 15 13 9 0 9 2
9 9 1 9 2 0 9 1 11 2
13 15 9 13 1 0 9 7 1 9 13 0 9 2
2 10 9
4 14 3 10 9
8 2 9 9 2 12 2 12 2
25 16 9 0 9 15 4 3 16 10 9 9 7 9 1 10 9 13 3 0 9 1 9 0 9 2
14 9 0 9 13 1 9 13 2 14 9 0 9 9 2
29 9 11 3 13 1 10 9 1 0 9 2 13 15 9 7 13 2 16 13 15 1 9 9 9 1 0 0 9 2
50 16 9 9 4 7 15 1 9 1 9 11 2 15 13 2 16 0 9 13 0 9 1 9 2 13 3 0 9 2 7 1 9 2 16 0 9 9 2 3 3 0 1 9 2 13 9 0 9 9 2
22 1 10 9 3 15 11 1 9 0 9 13 3 0 9 2 7 7 13 1 10 9 2
27 1 9 9 2 15 4 3 13 2 15 3 0 9 13 1 9 10 9 9 1 3 0 9 1 9 9 2
26 7 0 9 1 9 3 13 13 1 10 9 9 7 9 9 2 3 16 13 10 3 0 9 1 9 2
4 11 11 2 11
2 9 9
8 2 9 9 2 12 2 12 2
10 16 9 13 1 9 0 9 0 9 2
18 9 7 13 9 2 1 15 4 15 13 1 9 13 9 1 0 9 2
17 0 9 9 7 0 9 1 9 13 9 9 9 7 3 7 9 2
14 13 15 1 10 9 2 16 4 13 13 9 0 9 2
9 13 4 15 0 7 3 0 9 2
29 9 4 13 9 16 13 9 2 0 2 0 7 0 9 2 15 13 9 1 10 9 7 9 1 9 3 0 9 2
9 13 4 3 9 9 1 0 9 2
7 9 4 0 9 13 3 2
15 13 4 9 1 9 9 7 13 15 3 13 2 15 13 2
4 11 11 2 11
2 9 9
8 2 9 9 2 12 2 12 2
10 13 9 9 2 15 1 15 15 13 2
19 14 13 1 9 7 9 9 9 2 15 13 3 3 13 1 9 1 9 2
14 3 13 0 9 0 0 9 2 9 7 0 0 9 2
30 3 0 2 0 9 13 9 9 1 9 7 9 2 7 15 13 1 9 0 9 9 7 10 9 1 9 0 12 9 2
16 1 9 13 3 2 16 15 10 9 9 1 9 10 9 13 2
24 0 9 13 9 10 0 2 15 3 1 0 9 1 0 9 2 13 2 3 9 0 0 9 2
9 3 4 1 11 13 0 0 9 2
22 3 4 15 13 2 16 10 9 9 3 13 2 9 15 3 13 0 1 9 0 9 2
35 0 0 9 9 13 13 2 9 2 9 7 16 3 9 13 9 9 2 9 9 9 3 13 7 3 1 9 13 9 9 1 12 5 9 2
10 1 15 3 3 13 1 9 0 9 2
4 11 11 2 11
2 9 9
18 1 9 12 13 11 11 1 11 16 0 1 9 0 0 9 1 11 2
14 13 13 0 9 9 2 15 13 0 0 9 0 9 2
20 1 15 2 3 15 11 13 13 10 0 9 2 4 13 1 0 9 11 11 2
17 2 1 9 9 4 13 9 9 1 3 16 12 9 0 0 9 2
9 3 0 9 4 1 15 3 13 2
11 3 13 7 13 12 7 12 12 0 9 2
13 0 0 9 2 15 0 9 13 2 13 10 9 2
14 13 15 2 16 4 15 16 9 3 1 0 9 13 2
12 2 10 0 9 13 3 9 7 13 15 3 2
17 13 9 2 16 15 13 13 14 12 9 1 0 9 9 0 9 2
21 7 10 0 9 13 3 0 9 7 13 13 2 16 1 11 13 1 10 0 9 2
14 9 3 13 2 16 10 9 1 9 13 0 0 9 2
28 16 1 9 13 9 1 11 9 3 12 9 2 1 9 12 15 13 12 9 7 1 9 0 9 14 12 9 2
8 3 15 7 13 13 0 9 2
11 13 1 15 2 16 10 9 13 9 9 2
18 7 4 13 0 9 9 1 12 0 9 2 1 15 15 13 0 9 2
17 9 13 0 9 7 15 13 9 9 13 7 3 3 13 0 9 2
6 9 9 13 9 9 2
8 2 13 9 13 7 0 9 2
9 1 9 1 0 9 13 0 9 2
8 1 9 12 9 13 9 3 2
7 9 13 9 9 7 9 2
29 13 1 10 9 2 16 13 9 0 7 0 9 11 7 9 0 9 9 2 15 4 13 0 9 9 7 10 9 2
9 2 13 15 7 9 1 9 9 2
20 13 0 0 9 7 0 0 9 2 7 13 0 9 13 10 9 16 3 0 2
6 3 4 13 0 9 2
14 0 9 10 11 9 3 13 2 16 13 3 16 0 2
4 2 9 13 2
2 0 9
15 9 9 11 9 11 13 12 0 9 2 1 11 7 9 2
13 15 15 13 1 0 9 1 9 7 9 10 9 2
2 11 11
22 1 11 15 13 1 9 1 0 9 13 9 1 9 9 7 0 9 3 1 10 9 2
21 0 9 0 9 13 9 0 9 1 0 9 1 9 12 1 12 9 1 9 0 2
16 3 0 9 13 15 2 1 15 15 3 9 13 1 0 9 2
13 3 0 9 1 0 9 9 15 13 1 12 9 2
16 0 13 3 9 0 9 9 2 1 15 13 9 9 0 9 2
22 3 0 13 9 9 1 9 9 1 9 0 7 9 0 0 9 2 15 15 13 9 2
14 9 9 9 1 9 13 3 9 9 1 9 7 9 2
15 13 0 7 3 2 13 9 2 9 2 9 2 0 9 2
17 0 9 1 11 1 9 9 9 11 9 11 11 11 1 9 13 2
8 1 9 9 0 9 7 13 2
16 15 13 9 9 1 0 9 2 15 13 0 9 13 0 9 2
3 0 7 0
11 9 9 2 9 7 9 13 0 7 0 9
19 1 10 9 15 13 0 9 0 9 2 15 13 1 12 2 9 0 9 2
16 9 9 2 9 7 9 15 13 1 0 9 11 3 12 9 2
10 9 13 0 0 9 7 0 0 9 2
3 0 0 9
14 1 0 9 13 9 0 9 2 15 13 12 0 9 2
13 13 1 3 0 0 9 7 0 9 1 0 9 2
27 1 0 9 13 9 0 9 2 0 9 2 0 7 0 9 2 0 9 1 0 7 0 9 7 0 9 2
10 0 0 9 13 9 0 7 0 9 2
8 12 1 0 9 13 0 9 2
25 1 9 1 9 0 9 4 0 2 0 7 0 9 1 3 0 9 3 13 0 9 7 0 9 2
10 0 9 13 3 0 16 1 0 9 2
22 0 0 9 13 0 9 7 3 0 0 9 2 15 13 3 3 0 1 9 1 11 2
11 10 9 10 9 13 14 12 5 10 9 2
25 9 1 9 9 9 7 13 3 1 9 2 16 9 9 0 0 9 13 0 16 0 9 0 9 2
2 0 9
24 1 0 9 4 9 9 9 9 13 3 1 9 7 9 2 13 7 0 9 7 13 9 9 2
17 1 9 13 9 0 9 2 15 3 7 3 3 13 9 0 9 2
11 9 9 13 3 10 0 9 9 7 9 2
33 1 0 9 0 9 4 13 9 1 0 9 3 12 9 9 7 1 0 9 1 0 12 9 2 15 13 3 12 9 1 0 9 2
25 13 1 9 0 9 2 9 11 2 11 7 10 9 1 0 9 2 3 9 9 2 9 7 0 2
14 9 7 9 9 15 13 1 0 9 7 0 9 9 2
16 1 0 9 15 13 0 9 2 15 13 1 0 9 3 0 2
20 1 0 9 15 13 13 0 9 7 1 0 9 0 9 1 3 0 0 9 2
17 13 15 13 0 0 9 0 9 2 9 0 9 7 9 13 9 2
5 11 11 2 11 11
32 9 2 0 0 9 2 11 12 2 12 12 11 12 2 9 2 2 2 12 2 12 12 2 9 2 2 12 2 12 12 12 2
4 9 1 0 9
7 13 3 13 10 0 9 2
27 1 0 9 1 12 2 9 13 12 5 15 2 13 2 3 12 9 2 9 2 1 9 1 9 0 9 2
7 4 13 9 3 12 9 2
19 1 0 9 4 13 12 9 2 0 9 12 9 4 13 7 1 9 0 2
10 0 9 13 1 10 9 1 0 9 2
24 1 9 0 9 11 15 13 3 12 5 2 1 9 12 5 2 7 3 12 5 1 9 9 2
24 10 9 1 0 9 13 0 0 9 2 9 1 0 9 13 7 7 1 0 9 1 9 0 2
11 1 9 1 9 13 1 9 9 7 9 2
5 9 3 2 9 3
27 9 13 9 9 0 9 0 0 9 0 0 2 0 7 0 9 2 1 15 13 9 9 0 9 3 0 2
11 1 0 9 13 15 9 10 9 7 9 2
25 1 0 9 13 9 0 7 1 15 0 0 9 2 9 13 0 9 0 1 9 1 9 0 11 2
22 15 2 3 1 3 0 7 3 0 0 9 2 13 0 9 9 7 15 13 0 9 2
33 0 9 4 13 0 9 9 1 0 9 0 9 1 0 9 0 7 0 9 2 14 1 3 0 9 1 9 0 9 7 0 9 2
3 9 1 9
29 1 9 13 0 0 9 13 16 0 9 2 13 15 0 9 2 10 0 9 7 9 1 9 1 9 15 3 13 2
24 0 2 0 9 13 0 9 10 9 2 13 15 1 0 7 3 0 9 0 1 3 0 9 2
22 1 0 9 1 0 9 9 11 7 9 11 13 10 0 9 2 9 13 7 3 13 2
20 9 9 13 13 1 3 0 2 13 7 0 13 1 9 2 9 7 0 9 2
21 1 0 0 7 0 9 3 13 0 0 9 2 9 9 2 0 9 7 9 9 2
15 9 0 12 9 13 0 1 9 9 3 3 0 0 9 2
16 0 9 13 0 3 1 0 9 2 15 13 0 9 0 9 2
3 9 0 9
40 0 0 9 9 2 15 13 1 10 9 0 9 2 13 0 9 2 15 13 9 9 2 9 2 9 2 9 2 0 9 2 9 7 9 7 0 9 7 9 2
47 10 9 13 13 1 0 9 2 9 11 2 11 11 2 11 11 2 11 11 2 0 0 9 11 2 9 1 0 7 0 9 11 1 2 11 2 2 11 11 2 11 0 11 7 9 11 2
14 10 9 13 13 3 1 0 9 1 0 9 0 9 2
22 9 9 15 3 13 1 9 0 9 7 9 10 9 13 1 0 9 7 9 0 9 2
3 0 9 9
12 0 9 13 13 1 9 9 7 0 0 9 2
21 1 10 9 4 1 0 9 13 13 1 0 9 0 9 9 2 3 0 0 9 2
15 10 9 15 13 0 9 9 0 9 7 0 9 0 9 2
43 13 15 1 9 0 9 7 9 2 9 2 9 2 9 2 9 2 0 9 2 9 2 0 9 2 0 9 2 0 0 9 2 0 9 7 0 9 2 9 7 0 9 2
27 0 9 13 13 3 0 9 2 7 15 13 1 0 9 2 1 15 1 0 12 9 13 1 0 9 9 2
21 1 9 1 0 9 13 10 9 1 0 9 2 13 15 3 1 0 7 0 9 2
21 1 9 9 1 0 9 13 0 13 1 9 9 2 0 0 9 2 2 9 2 2
21 9 9 4 13 9 0 9 2 3 3 9 0 9 0 7 0 9 1 0 9 2
13 9 9 0 9 13 0 0 9 2 0 10 9 2
23 0 9 0 9 13 1 9 9 9 9 2 7 4 3 3 13 9 9 1 0 0 9 2
2 11 0
28 1 9 9 1 9 0 9 11 1 9 12 13 0 9 9 0 9 12 9 2 1 0 9 15 9 12 9 2
17 1 0 9 9 9 0 9 3 13 2 9 13 13 12 2 12 2
11 9 9 7 9 10 9 13 9 0 9 2
20 1 12 2 12 13 0 9 15 9 12 9 2 0 9 9 0 9 12 9 2
17 0 9 13 0 9 11 12 9 2 0 9 11 7 0 9 11 2
3 11 11 2
2 11 11
14 9 2 0 0 9 2 0 2 9 2 2 11 12 2
21 12 12 11 12 2 9 2 2 12 2 12 12 2 9 2 2 12 2 12 12 12
3 9 2 9
15 0 9 11 1 11 2 1 10 0 9 13 0 15 13 2
7 3 1 9 1 0 9 2
26 16 15 9 1 15 1 9 0 9 0 1 0 9 13 2 13 15 15 14 9 2 16 13 1 9 2
14 1 0 9 3 13 9 7 15 2 16 4 15 13 2
11 1 0 9 9 13 11 9 3 1 9 2
1 11
3 1 0 9
18 9 11 2 11 1 0 9 9 7 9 2 15 13 0 9 9 11 2
19 0 9 10 9 15 13 1 9 1 9 2 0 9 7 7 1 9 9 2
14 9 9 3 13 0 9 9 2 16 13 0 9 9 2
24 9 2 11 2 11 2 0 12 2 12 12 11 2 11 2 9 2 9 2 2 12 2 12 12
19 9 11 1 9 7 9 0 9 7 0 9 1 9 2 0 7 0 9 2
14 1 0 9 15 13 13 1 0 2 0 7 0 9 2
9 1 9 9 13 9 7 0 9 2
21 9 2 11 2 0 12 2 12 12 0 11 2 9 2 9 2 2 12 2 12 2
3 0 7 0
21 1 12 12 9 13 1 15 9 0 0 7 0 9 2 11 2 0 9 0 9 2
14 10 3 0 9 2 0 9 2 13 9 7 13 9 2
15 1 0 9 13 9 0 9 7 3 13 0 9 0 9 2
13 13 4 1 15 1 0 9 0 9 11 11 11 2
14 2 3 4 13 1 9 2 16 15 9 13 1 9 2
23 3 1 9 12 4 13 1 0 9 9 1 12 9 9 2 1 9 3 13 1 12 9 2
19 13 15 0 2 16 13 13 0 7 3 0 9 2 16 13 3 1 9 2
18 13 4 2 16 9 9 13 0 7 1 9 3 13 9 1 10 9 2
20 7 4 3 13 0 9 1 9 2 7 0 0 9 4 13 13 7 3 13 2
10 2 15 13 13 1 0 9 0 9 2
21 13 4 1 9 0 9 9 12 2 15 13 9 1 0 9 14 12 9 1 9 2
11 10 9 13 7 0 9 1 3 0 9 2
12 13 9 1 0 9 12 12 9 1 0 11 2
17 15 1 10 9 15 13 2 7 13 15 1 9 16 0 0 9 2
22 9 9 12 13 3 1 9 7 10 9 13 13 9 7 0 9 1 9 0 0 9 2
14 13 7 0 9 2 3 0 0 9 1 9 0 9 2
10 2 13 4 1 9 3 1 0 9 2
10 13 4 15 1 0 0 9 3 9 2
23 13 4 3 0 9 2 13 0 0 9 2 9 2 7 3 4 13 0 2 0 9 9 2
9 1 0 12 0 9 13 12 12 2
12 0 9 4 3 13 0 9 9 7 0 9 2
5 1 9 7 1 9
12 9 1 0 9 7 9 13 16 9 2 0 3
7 9 2 0 9 0 9 2
10 13 4 15 1 12 9 2 0 9 2
23 1 0 9 0 9 0 9 15 10 9 13 1 3 0 9 12 9 1 9 9 0 9 2
41 15 2 15 3 1 10 3 0 9 13 0 0 9 2 3 13 13 1 9 2 16 1 0 9 2 0 1 12 2 9 2 13 9 1 9 0 9 1 0 9 2
2 11 11
18 13 3 2 1 9 2 1 9 12 9 0 9 2 15 13 0 9 2
18 7 15 13 15 9 13 2 9 1 9 2 2 13 9 1 12 9 2
28 13 7 9 2 16 9 9 0 9 2 3 2 16 13 0 0 9 0 0 9 2 3 3 1 9 9 13 2
50 1 15 2 3 15 7 1 3 0 9 2 1 15 15 3 13 2 14 1 9 2 0 0 9 2 9 3 13 1 3 12 9 0 9 7 10 13 0 9 2 4 13 1 11 11 2 10 0 9 2
24 2 13 0 9 9 3 15 2 16 1 9 13 0 9 1 9 3 1 9 0 9 0 11 2
30 1 9 9 0 9 13 15 3 0 9 1 15 2 15 13 1 9 13 1 9 9 2 0 0 7 0 9 0 9 2
19 3 4 7 15 13 9 1 9 2 16 15 15 1 10 9 13 1 9 2
13 15 13 9 0 9 9 12 10 0 9 1 11 2
16 2 1 0 9 15 13 0 9 2 7 9 1 9 10 9 2
15 9 1 9 3 13 3 9 2 7 15 13 3 3 3 2
7 13 15 9 16 0 0 2
18 13 1 15 2 16 4 9 1 0 9 13 9 7 9 9 3 0 2
9 7 10 9 15 1 0 9 13 2
6 2 15 13 0 9 2
19 13 15 7 2 16 9 13 7 0 9 1 0 9 9 9 1 10 9 2
26 9 9 1 10 9 15 13 1 2 0 2 9 0 9 14 1 0 9 9 9 3 3 1 9 12 2
34 1 0 9 9 9 4 3 9 9 12 7 12 13 13 9 0 9 9 2 16 3 1 9 12 4 13 13 1 0 9 7 9 9 2
9 7 15 15 13 0 9 16 15 2
24 7 15 13 14 9 7 9 9 2 7 2 1 9 1 0 9 9 2 3 7 9 0 9 2
11 2 13 1 9 9 0 2 0 9 2 2
16 9 2 15 3 3 13 13 2 3 13 1 9 3 0 9 2
35 16 7 1 9 2 16 13 11 1 0 9 2 16 15 1 15 13 15 1 12 9 13 9 9 2 13 1 0 9 9 9 14 1 9 2
17 7 13 15 1 9 9 1 9 1 3 0 9 1 0 12 9 2
11 2 15 13 3 3 2 16 13 0 9 2
21 15 13 9 2 16 3 13 9 9 2 15 3 3 13 0 9 7 3 13 13 2
8 3 3 15 13 1 10 9 2
5 2 13 9 9 2
3 3 9 2
19 15 13 2 16 3 2 3 13 1 0 9 2 13 10 9 3 0 9 2
24 0 9 10 9 2 16 15 15 13 2 15 1 9 13 2 7 9 14 3 13 2 3 13 2
14 7 9 15 13 13 0 9 7 3 13 1 0 9 2
27 2 1 9 1 0 9 4 3 13 10 0 9 2 16 1 0 9 0 9 0 9 13 3 16 0 9 2
27 16 15 13 1 0 9 13 1 3 0 9 2 13 15 10 0 7 0 9 13 7 1 9 9 0 9 2
14 2 15 13 3 0 1 9 0 9 13 9 0 9 2
4 7 3 14 2
22 15 9 13 7 1 0 9 2 3 1 9 9 10 9 1 0 2 16 0 9 9 2
27 7 3 2 1 15 15 13 7 9 0 9 1 9 0 9 2 9 1 9 9 2 9 7 9 0 9 2
8 2 9 13 3 0 0 9 2
5 13 1 15 9 2
15 0 9 0 9 13 9 0 9 14 9 2 3 0 9 2
23 13 1 15 2 16 9 0 9 9 1 0 0 9 13 13 0 9 1 0 0 0 9 2
12 7 4 13 9 0 9 1 10 9 0 9 2
29 3 4 13 9 9 0 9 3 1 10 0 9 2 3 7 9 9 7 0 9 1 10 0 9 2 1 0 9 2
8 2 3 7 9 9 3 13 2
13 14 3 13 3 16 0 7 0 9 1 0 9 2
36 13 4 15 0 9 2 9 0 9 9 1 15 2 16 1 9 13 9 0 9 7 4 13 0 9 3 1 0 9 2 3 1 9 0 9 2
17 1 15 15 13 13 3 2 1 11 2 3 1 9 0 0 9 2
19 1 0 9 3 13 1 0 9 9 2 7 15 1 9 7 9 0 9 2
18 9 2 3 9 13 2 13 1 9 0 9 1 9 9 0 9 9 2
14 2 13 13 2 16 15 9 15 4 13 9 1 9 2
4 7 3 14 2
18 3 1 9 10 9 4 3 13 9 9 3 16 9 2 3 9 9 2
33 0 9 9 1 0 9 7 1 9 3 1 9 9 2 0 9 0 7 0 9 4 13 1 0 9 2 14 0 2 7 7 0 2
18 7 14 15 2 3 15 13 7 0 0 9 1 9 3 0 0 9 2
18 7 13 3 0 1 9 9 9 7 9 7 13 3 9 2 7 13 2
7 3 7 9 13 3 3 2
8 2 13 15 15 7 0 9 2
8 3 2 16 13 3 3 0 2
29 3 14 10 0 9 3 13 9 9 1 0 9 14 1 12 9 9 2 7 13 1 9 13 3 12 1 12 9 2
2 9 2
14 9 2 15 13 1 12 9 3 0 9 2 3 13 3
7 9 1 9 13 9 9 9
2 11 11
18 9 1 9 9 7 9 1 0 9 1 0 9 4 13 1 9 9 2
17 0 0 9 15 13 13 9 0 9 9 2 15 13 9 0 9 2
16 9 0 9 11 11 13 0 9 13 2 7 1 15 3 13 2
23 3 4 15 13 3 12 9 9 9 2 1 15 4 0 9 13 9 1 9 9 9 9 2
23 1 0 9 10 9 0 10 9 13 2 16 9 1 0 9 12 10 0 9 13 3 0 2
34 1 11 11 7 11 11 3 13 0 9 2 3 15 13 1 9 2 16 1 9 1 9 9 12 1 9 12 1 15 13 12 0 9 2
43 1 0 9 10 9 15 3 13 2 0 7 0 9 2 2 2 2 13 13 14 9 1 10 9 3 0 2 16 13 9 3 9 2 9 2 7 15 0 9 2 2 2 2
21 1 0 9 3 13 2 16 9 15 13 13 7 3 7 13 1 9 0 9 9 2
12 15 13 1 0 13 7 1 0 9 0 9 2
47 16 0 9 9 9 13 10 9 13 2 15 1 15 15 1 10 9 3 13 2 2 13 9 9 1 9 3 0 0 9 3 0 0 9 9 2 3 0 0 9 9 0 9 1 0 9 2
35 1 0 9 15 4 13 12 12 9 13 1 10 9 2 16 4 7 3 13 1 15 13 12 9 2 1 10 9 4 13 3 9 7 9 2
18 3 15 1 9 9 13 9 0 0 9 2 15 4 13 0 0 9 2
33 13 2 16 3 1 9 9 10 9 0 9 13 2 0 9 3 13 9 9 7 15 13 0 9 2 15 4 13 1 3 0 9 2
9 0 0 9 15 13 1 0 9 2
17 13 0 15 13 2 10 9 4 9 9 9 7 0 9 13 13 2
16 1 0 9 4 13 1 9 1 9 0 9 13 0 0 9 2
8 2 1 1 9 0 9 2 2
16 1 9 0 4 9 13 13 0 0 9 0 1 9 0 9 2
19 7 13 9 1 9 0 0 9 10 7 15 9 4 13 3 0 0 9 2
31 13 9 9 3 2 16 4 15 13 9 1 0 9 9 9 2 13 9 2 1 15 4 1 10 0 9 3 13 13 9 2
38 1 0 0 9 1 9 7 0 9 2 15 1 10 9 13 9 3 1 9 2 3 9 13 0 0 9 9 9 2 15 1 9 1 9 10 9 13 2
7 13 4 4 13 1 9 2
3 9 13 9
5 11 2 0 11 2
26 9 0 9 11 3 13 0 9 0 9 1 9 11 3 2 16 15 1 15 13 9 0 1 0 11 2
16 9 9 11 2 11 13 2 16 9 9 13 12 9 0 9 2
29 9 4 10 9 2 15 13 1 9 1 0 9 1 9 7 11 1 9 9 9 1 11 2 13 3 1 0 9 2
15 11 7 11 13 9 9 9 1 9 9 1 11 7 11 2
14 3 13 2 16 9 11 14 13 2 7 13 3 13 2
14 1 9 11 15 3 13 0 9 1 11 11 2 11 2
29 1 11 1 9 1 0 9 0 9 13 14 9 2 15 9 9 11 13 2 7 3 0 9 2 15 11 3 13 2
5 11 1 11 1 9
9 0 9 11 1 11 11 11 2 11
7 11 13 9 2 2 2 2
12 10 12 9 3 10 9 13 1 9 0 9 2
18 9 0 9 13 9 0 9 2 9 7 9 2 0 1 9 0 9 2
7 3 15 4 13 1 11 2
38 3 7 14 3 2 16 4 0 0 9 13 1 15 0 16 10 9 1 0 9 2 7 3 3 2 16 15 11 13 10 9 1 9 1 10 0 9 2
14 0 9 13 1 9 1 11 7 13 1 9 1 11 2
22 3 16 1 0 9 7 3 9 13 2 16 9 13 1 9 0 1 9 1 0 9 2
5 0 9 13 9 2
36 13 10 0 9 0 9 2 0 9 11 11 2 1 11 2 16 4 15 3 13 13 9 0 0 7 0 9 1 9 1 0 9 1 0 9 2
14 11 3 3 13 7 11 3 13 0 0 7 0 9 2
12 3 7 13 0 9 3 1 11 3 0 9 2
16 11 14 13 15 0 9 7 13 9 1 15 9 1 0 9 2
14 14 12 13 13 2 16 4 0 9 13 13 1 11 2
19 3 13 2 3 15 13 2 15 3 1 9 7 13 0 9 9 7 9 2
9 11 2 3 0 2 0 13 9 2
7 0 13 7 7 0 9 2
30 9 0 9 13 3 9 10 0 0 9 2 9 3 13 2 2 15 13 13 9 1 11 7 11 2 13 0 0 9 2
32 3 0 13 0 9 2 16 3 11 3 13 9 1 11 2 16 4 15 3 13 3 13 3 1 11 7 13 1 15 0 9 2
15 10 15 3 13 13 9 11 7 9 0 0 9 0 9 2
29 11 7 3 13 2 16 10 0 9 7 9 13 0 7 1 9 13 2 16 13 12 9 0 9 1 0 0 9 2
16 13 0 2 16 0 9 1 0 9 13 11 3 16 0 9 2
17 13 7 3 0 2 16 11 13 1 0 9 1 10 9 3 9 2
22 16 15 7 13 0 2 13 0 9 9 1 0 9 2 1 15 15 13 1 0 9 2
19 9 10 0 9 2 16 7 3 0 0 9 13 13 7 0 9 0 9 2
10 1 11 10 9 13 15 13 0 9 2
24 7 3 7 0 9 16 0 0 11 13 0 9 0 9 9 11 7 13 15 3 1 9 9 2
24 3 15 3 13 9 9 9 11 11 2 15 13 9 0 9 1 9 1 0 9 1 0 9 2
15 1 0 9 7 9 13 3 0 13 9 1 9 7 9 2
34 9 7 13 2 16 10 9 13 0 2 7 15 1 15 0 9 2 13 0 9 7 13 0 7 16 0 0 9 1 9 9 0 9 2
15 9 1 0 9 11 11 2 11 11 2 13 9 14 1 9
5 9 11 2 9 9
10 0 9 2 11 12 2 12 2 12 2
21 1 9 4 13 9 2 0 1 9 0 9 2 15 13 1 9 1 9 9 9 2
15 13 0 13 10 9 1 9 2 7 13 15 1 9 9 2
5 0 9 3 13 2
7 13 15 9 1 0 9 2
14 15 13 0 9 7 9 1 9 13 0 9 0 9 2
11 0 9 9 9 3 13 7 9 15 13 2
16 9 9 9 2 16 0 9 13 7 13 0 9 2 13 0 2
6 13 3 1 0 9 2
22 10 9 9 13 2 13 4 13 0 9 2 1 0 9 4 13 9 13 9 0 9 2
22 16 4 9 9 13 2 16 0 9 9 13 9 1 11 2 3 13 9 10 9 3 2
8 1 9 9 2 11 11 2 11
6 1 0 9 13 0 9
19 9 0 9 2 13 0 9 1 0 9 2 13 9 2 7 13 9 1 9
4 11 11 2 11
25 13 2 14 9 9 11 1 12 9 9 11 1 11 11 2 3 9 1 9 9 15 11 3 13 2
12 9 13 15 0 7 3 0 1 0 0 9 2
38 11 3 13 0 9 10 0 0 9 2 16 13 0 9 2 7 10 0 9 1 9 0 9 13 13 1 9 0 9 0 9 0 9 1 9 0 9 2
34 3 16 11 13 11 11 7 11 0 2 11 11 11 7 9 11 2 11 11 11 7 11 11 2 7 11 11 11 2 13 0 9 11 2
5 0 9 1 0 9
36 16 1 9 11 13 1 12 2 9 11 11 11 7 9 1 9 9 15 3 13 0 11 11 2 3 13 1 9 2 15 1 11 9 3 13 2
23 9 2 11 13 0 0 9 2 0 1 0 9 2 7 15 10 0 0 9 1 11 13 2
10 13 0 9 9 2 10 9 7 9 2
7 1 10 15 13 11 3 2
21 3 0 9 1 11 7 0 9 12 2 12 1 11 13 2 16 15 1 11 13 2
18 13 0 9 1 9 1 11 2 15 0 3 13 1 9 12 2 12 2
27 3 3 13 9 9 2 9 2 11 2 0 1 9 3 1 11 2 15 15 13 1 9 2 13 1 9 2
21 1 0 9 13 0 9 11 9 9 7 13 15 1 9 9 2 3 13 9 11 2
25 0 9 11 2 11 13 9 1 11 7 3 3 15 13 1 0 9 1 11 2 12 2 12 2 2
14 7 1 12 9 3 13 2 16 9 13 9 2 2 2
26 9 9 1 12 9 1 0 9 7 9 13 1 9 13 11 9 14 1 12 2 9 2 3 13 9 2
17 1 10 9 4 0 9 12 9 13 2 3 0 13 1 0 9 2
28 3 4 13 13 2 7 3 15 15 13 2 16 9 3 13 1 15 2 15 13 9 2 13 1 9 9 11 2
15 0 9 3 13 2 16 0 9 13 11 3 1 0 9 2
30 9 1 0 0 9 13 3 0 7 13 1 15 13 14 1 9 2 16 13 9 0 9 2 9 7 0 9 1 9 2
22 15 13 0 9 11 2 15 1 9 9 13 9 0 9 7 1 9 15 3 14 13 2
17 13 7 0 9 11 2 7 3 15 13 1 9 9 15 1 15 2
11 1 9 9 0 9 13 3 9 0 9 2
19 1 9 13 11 12 2 12 3 1 0 11 2 15 3 13 3 1 11 2
29 1 0 9 1 9 1 0 11 13 11 3 1 10 9 2 3 13 1 9 11 7 13 15 0 9 12 2 12 2
6 13 9 9 7 9 2
16 9 0 9 13 7 3 1 15 0 2 1 0 9 9 9 2
19 9 11 11 11 15 1 0 9 13 9 2 16 13 13 1 9 0 9 2
15 15 15 1 15 13 2 7 9 9 15 1 10 9 13 2
14 0 3 9 9 3 13 2 7 10 9 3 15 13 2
23 13 0 9 9 2 11 13 1 11 12 2 11 1 11 13 1 11 2 11 13 1 11 2
31 3 1 15 0 9 2 7 15 0 2 13 11 9 7 15 13 3 3 2 16 0 9 13 1 9 10 9 1 0 9 2
13 3 15 13 1 0 9 13 15 0 9 0 9 2
14 7 3 1 0 9 2 16 9 9 0 9 3 13 2
15 7 7 1 9 13 2 16 15 3 13 2 3 7 13 2
32 16 11 13 1 9 1 9 9 3 12 9 9 2 13 4 15 15 7 3 13 2 9 1 12 2 9 9 11 13 0 9 2
17 16 11 13 15 1 12 10 9 2 13 15 1 10 0 9 13 2
6 10 9 13 3 0 2
26 16 4 13 9 2 3 3 1 9 2 16 1 15 4 0 9 3 13 2 13 1 0 9 11 11 2
26 3 15 0 9 3 13 2 16 1 0 9 9 2 16 15 1 9 13 13 3 0 2 15 9 13 2
21 13 15 7 2 16 4 0 9 11 13 0 9 2 9 10 9 7 7 15 0 2
4 3 0 9 2
12 3 4 15 15 13 13 1 9 0 9 9 2
2 0 9
24 16 13 1 0 9 0 9 11 11 2 12 2 3 0 2 13 15 1 9 0 9 0 9 2
16 0 0 9 2 12 2 13 0 9 1 9 7 9 0 9 2
16 13 1 12 9 2 9 1 9 2 15 15 1 9 3 13 2
24 9 3 13 9 9 1 9 9 14 1 9 9 2 9 9 7 0 0 9 1 9 0 9 2
9 2 11 2 2 11 12 2 12 2
3 9 11 11
20 16 15 13 13 2 3 15 3 13 2 1 9 13 1 9 9 11 2 2 2
4 0 9 9 11
2 11 2
19 9 0 0 9 15 12 0 9 11 11 9 0 1 10 9 4 3 13 2
19 1 15 9 13 1 9 9 3 2 16 4 15 13 1 9 1 0 9 2
39 1 9 7 1 9 15 1 11 13 0 0 9 9 9 11 9 2 11 9 2 11 0 9 2 11 11 2 11 11 2 11 11 2 11 9 7 11 9 2
16 9 15 9 4 13 13 0 0 9 1 9 1 9 0 9 2
10 13 3 1 0 9 1 9 9 9 2
44 0 9 11 11 15 13 0 9 0 9 2 9 11 11 11 2 9 11 9 0 9 0 9 9 11 11 11 7 9 11 9 11 11 2 3 0 9 1 9 9 7 9 9 2
1 3
19 0 9 1 0 11 13 1 9 1 12 9 7 1 0 9 1 12 9 2
42 9 0 2 9 2 11 13 9 3 13 9 9 11 2 11 2 11 7 11 2 1 9 3 2 16 10 0 9 9 7 0 9 11 11 4 13 9 0 9 0 11 2
11 9 4 13 4 13 12 2 9 1 11 2
4 1 0 0 9
14 11 11 2 0 9 2 9 11 2 12 9 2 2 2
17 9 13 0 9 9 2 9 2 9 2 9 7 9 9 0 9 2
29 13 13 15 0 9 1 9 9 7 0 9 2 13 1 9 9 9 0 9 7 13 13 9 1 9 1 0 9 2
16 0 13 7 9 0 9 9 7 9 9 0 0 9 1 9 2
33 11 11 2 11 11 2 11 2 9 2 1 0 1 11 2 9 9 11 2 11 12 2 12 9 2 5 12 9 2 0 9 2 2
23 0 0 9 0 9 7 0 9 2 3 0 9 9 11 2 7 3 0 9 0 0 9 2
40 9 13 1 9 0 9 1 9 0 2 11 7 11 2 2 1 10 9 1 0 0 9 1 9 0 9 2 15 13 9 3 0 9 1 9 0 9 2 11 2
25 13 7 10 9 9 0 9 11 2 0 9 0 11 2 9 9 11 11 11 3 9 2 15 9 2
23 7 15 3 13 2 16 13 0 9 9 10 9 2 15 13 1 9 0 9 1 15 0 2
21 9 13 14 9 1 9 0 9 7 9 0 9 7 9 1 0 0 7 0 9 2
49 9 9 11 7 10 0 9 2 0 9 1 0 9 2 9 9 7 9 3 0 9 2 16 13 11 2 7 11 2 3 9 13 1 0 2 1 15 0 9 0 9 4 13 16 0 0 9 9 2
8 0 13 3 2 3 3 1 15
2 11 11
8 13 13 2 13 3 10 9 2
24 9 7 9 13 13 3 2 13 1 9 9 12 1 0 9 3 0 11 11 1 11 1 11 2
4 9 9 13 2
21 1 0 9 10 9 15 0 9 0 11 9 13 7 15 3 1 10 9 13 13 2
6 3 1 15 13 3 2
10 9 9 11 13 0 9 9 0 9 2
9 1 0 9 1 9 12 4 13 2
13 1 9 12 15 13 9 13 7 15 15 13 13 2
7 1 9 3 3 13 9 2
18 3 1 9 0 9 4 13 13 1 9 3 2 13 1 9 0 9 2
22 16 15 1 9 13 2 16 15 1 11 4 13 13 2 1 9 12 14 3 9 13 2
5 7 3 2 2 2
7 9 12 15 13 1 11 2
7 13 1 9 1 9 9 2
16 16 15 13 13 1 9 2 13 7 9 7 13 1 0 11 2
17 3 4 13 1 9 2 3 3 13 1 15 2 13 15 14 3 2
17 1 9 0 9 13 3 3 2 16 4 1 9 13 9 1 9 2
6 13 3 3 0 9 2
18 9 3 1 11 13 9 10 0 9 7 3 15 7 15 13 1 11 2
27 15 0 9 2 9 0 1 9 2 9 2 9 0 11 7 0 9 2 13 1 9 9 7 0 0 9 2
13 13 3 3 0 9 7 13 0 9 1 9 9 2
10 3 13 9 2 9 7 9 1 9 2
4 13 9 0 2
8 1 9 9 13 1 0 9 2
18 3 1 9 13 12 9 2 12 1 9 2 12 1 15 7 0 9 2
8 15 9 13 14 12 9 9 2
9 9 3 3 13 16 1 12 9 2
12 0 9 2 0 0 9 2 0 9 2 9 2
11 7 15 13 13 12 9 0 9 0 9 2
7 9 7 9 13 0 3 2
9 1 9 3 13 12 9 0 9 2
12 9 1 15 13 0 2 0 13 13 1 9 2
14 1 9 13 3 9 2 3 3 9 2 9 7 9 2
12 3 4 15 13 2 9 15 14 3 3 13 2
10 1 9 13 12 9 7 12 0 9 2
11 3 12 7 12 10 9 13 1 0 9 2
9 1 0 9 13 12 9 0 9 2
3 9 13 2
22 1 9 13 9 2 1 0 13 2 7 9 13 3 1 9 0 9 2 13 9 11 2
25 3 13 2 7 16 13 15 3 3 0 7 0 2 13 15 1 9 13 10 9 2 15 13 9 2
10 3 0 9 13 3 0 9 0 9 2
9 9 1 9 7 9 13 9 11 2
7 9 15 13 3 1 9 2
4 13 12 9 2
21 13 9 2 15 4 15 1 10 9 13 13 16 1 15 2 13 3 0 2 13 2
13 1 0 9 1 9 13 7 9 2 3 1 9 2
13 3 14 9 11 2 11 9 11 11 1 0 9 2
17 13 3 7 3 2 16 3 13 1 9 10 9 1 0 0 9 2
13 1 15 10 9 13 0 0 9 1 0 9 9 2
31 9 4 14 13 2 16 4 3 1 9 3 4 13 0 9 0 0 9 2 3 9 2 16 4 13 2 1 15 4 13 2
8 13 3 0 1 9 0 9 2
14 1 3 0 9 13 9 2 16 13 13 0 0 9 2
15 0 7 0 9 15 1 15 14 3 13 0 0 0 9 2
24 15 15 3 13 2 13 0 0 9 2 15 13 3 1 9 7 15 1 15 13 3 1 9 2
6 7 15 0 9 9 2
16 13 15 2 16 4 3 13 13 3 3 0 9 2 0 9 2
15 9 0 9 13 13 3 0 9 0 9 7 0 0 9 2
20 13 3 13 9 2 16 15 13 2 3 3 15 9 13 2 13 11 2 11 2
15 9 0 10 9 13 16 9 7 9 2 15 15 3 13 2
6 14 15 7 3 13 2
11 13 4 9 3 13 2 16 4 13 3 2
5 13 15 13 9 2
5 14 13 3 9 2
26 9 11 3 13 1 0 9 2 15 15 1 9 13 1 9 7 3 2 16 1 0 9 13 0 9 2
7 9 9 4 13 0 9 2
7 15 15 13 13 2 13 2
11 15 15 4 13 1 15 2 13 15 9 2
14 9 14 3 2 13 1 11 10 9 1 9 0 9 2
13 13 2 16 3 9 2 15 3 13 0 9 0 2
17 1 0 9 15 14 9 13 13 3 2 16 4 0 9 3 13 2
5 0 9 13 0 9
10 9 1 3 16 12 9 13 1 9 9
5 11 2 11 2 2
26 9 0 9 13 1 0 9 10 9 3 0 7 3 1 9 9 7 9 0 9 13 9 0 9 9 2
17 13 15 1 0 9 9 0 9 0 9 2 15 13 0 0 9 2
25 1 9 2 15 13 1 9 9 7 9 2 13 12 0 9 2 10 9 9 13 12 5 0 9 2
13 1 0 9 1 9 13 12 9 0 12 5 9 2
24 10 0 9 13 1 9 9 7 9 1 0 9 2 15 13 3 16 12 5 9 1 0 9 2
18 14 12 5 13 10 9 16 0 7 9 1 12 5 9 9 16 0 2
15 1 9 0 9 13 0 9 0 1 9 0 12 5 9 2
18 3 13 3 9 2 15 13 3 2 9 2 0 9 2 9 7 9 2
14 16 0 13 10 9 9 0 2 0 7 15 0 9 2
16 9 10 0 9 13 9 1 12 5 9 2 9 1 12 5 2
16 9 1 12 5 9 1 9 10 0 9 1 0 12 9 13 2
15 1 0 12 9 13 9 0 9 9 1 12 5 9 9 2
7 1 9 15 13 12 5 2
10 9 1 3 16 12 9 13 9 9 2
8 3 13 3 1 0 9 9 2
23 1 9 0 9 1 0 9 13 1 9 7 9 9 10 0 9 9 1 12 5 0 9 2
12 9 0 9 15 13 9 0 12 5 0 9 2
20 9 1 12 12 9 0 9 13 2 16 10 0 9 13 1 0 12 9 0 2
20 1 12 5 13 13 0 7 1 9 3 16 0 2 15 15 13 3 0 9 2
3 15 13 9
2 11 11
11 1 0 9 15 9 13 9 7 13 9 2
3 15 13 2
18 1 9 0 9 10 0 0 9 14 9 7 0 9 1 0 9 13 2
28 3 15 13 9 0 9 0 2 9 3 3 15 0 2 16 15 3 13 13 2 3 14 13 11 2 7 0 2
16 13 2 14 0 2 13 9 9 7 9 9 1 15 13 9 2
29 13 14 9 9 2 16 1 10 9 13 3 15 2 15 1 0 9 0 7 0 9 9 13 3 16 15 0 9 2
12 13 1 15 2 16 15 13 10 0 9 9 2
5 15 13 3 0 2
14 13 7 14 1 15 12 0 2 13 1 15 1 15 2
17 13 2 14 3 0 0 9 1 9 2 13 15 9 9 1 9 2
16 15 4 13 14 7 1 0 9 2 15 3 7 1 15 15 2
11 13 15 3 3 2 16 15 9 13 9 2
3 3 0 2
23 3 13 9 13 0 9 2 16 15 13 2 16 9 13 0 1 15 13 1 9 1 9 2
37 9 13 13 9 9 2 16 15 13 1 15 2 16 10 9 13 13 2 16 9 13 15 13 2 16 15 9 13 1 9 1 9 7 9 13 9 2
14 0 9 13 3 3 9 2 15 4 7 13 13 0 2
22 1 10 9 2 3 13 9 3 1 9 0 2 13 9 1 9 3 9 7 2 9 2
10 3 0 9 15 4 3 1 9 13 2
32 15 13 3 11 2 13 2 14 9 0 9 1 10 0 7 13 2 14 15 9 1 9 2 13 9 15 0 9 1 9 9 2
20 3 7 13 9 2 15 4 0 13 13 2 1 15 7 9 13 3 7 9 2
5 3 1 11 2 2
12 10 9 3 13 14 1 9 2 13 3 0 2
30 0 9 10 9 1 0 9 15 13 1 3 0 0 9 9 2 9 9 13 9 0 9 13 7 13 1 9 1 9 2
12 15 7 13 7 15 13 1 10 0 9 9 2
27 15 0 2 14 7 14 0 9 13 2 16 9 2 15 1 10 9 7 1 10 9 3 13 2 13 3 2
5 13 15 9 9 2
5 11 2 11 2 2
31 0 9 11 2 0 10 9 9 2 9 7 0 9 2 15 13 13 9 2 16 0 9 1 15 3 13 9 1 0 9 2
24 9 9 1 0 9 13 3 1 9 2 1 0 9 1 0 9 1 9 11 13 11 9 9 2
24 0 9 9 2 13 3 1 9 2 1 9 15 13 9 0 9 2 4 13 13 0 9 9 2
26 11 1 15 1 9 0 9 1 0 9 13 13 9 1 0 7 0 9 2 15 13 7 9 3 0 2
20 0 9 0 9 11 11 13 9 2 16 9 1 9 1 11 1 10 9 13 2
22 1 1 0 9 1 0 9 1 0 9 7 9 0 11 1 0 9 13 1 3 0 2
13 15 9 1 9 13 7 1 0 9 10 0 9 2
27 1 1 0 9 1 9 4 3 13 13 1 0 9 9 1 9 2 7 3 1 10 0 9 1 10 9 2
17 0 9 4 3 9 13 1 10 9 9 9 2 13 11 1 11 2
5 9 1 9 11 13
5 11 2 11 2 2
27 1 9 2 16 4 7 3 4 9 13 9 9 11 11 1 0 0 9 2 13 11 0 9 1 10 9 2
12 1 9 1 9 11 15 13 9 11 11 11 2
20 1 11 15 9 1 0 9 3 13 11 2 7 13 1 0 9 1 9 9 2
25 9 13 9 2 16 9 0 9 13 0 9 7 16 1 9 2 15 15 13 15 2 13 13 9 2
22 10 9 14 13 11 1 0 7 13 9 2 16 13 9 0 9 7 0 9 1 9 2
28 9 0 9 15 1 11 3 3 13 15 2 1 11 7 14 13 0 9 2 1 15 13 13 14 1 0 9 2
13 7 14 13 10 9 10 9 7 1 9 0 9 2
25 1 9 11 2 3 14 13 11 0 13 1 9 9 11 2 9 9 13 2 13 1 9 0 9 2
22 3 13 0 15 1 9 3 13 2 13 7 2 16 4 10 9 13 0 9 1 9 2
16 13 2 16 13 0 1 9 0 9 13 0 9 9 7 9 2
22 9 9 3 9 9 0 9 3 13 2 13 15 3 2 16 4 4 13 10 0 9 2
3 9 1 9
5 11 2 11 2 2
15 9 9 0 13 0 0 9 11 11 2 1 11 1 11 2
27 1 9 1 0 9 13 1 0 9 0 9 11 11 2 13 10 0 9 7 13 15 1 0 9 1 9 2
12 0 0 9 0 9 13 2 9 9 13 9 2
2 0 9
9 9 0 9 9 2 9 2 12 9
6 11 2 11 2 2 12
6 11 2 11 2 2 12
8 11 2 11 2 12 2 12 2
4 9 2 12 2
5 11 2 11 2 2
5 11 2 11 2 2
4 9 2 12 2
5 11 2 11 2 2
5 11 2 11 2 2
7 11 2 11 2 2 12 2
2 9 2
7 12 2 11 2 11 2 2
5 11 2 11 2 2
7 11 2 11 2 2 12 2
2 9 2
9 12 2 11 2 11 2 2 12 2
5 9 2 12 9 2
8 12 2 11 2 11 2 2 12
6 11 2 11 2 2 12
7 11 2 11 2 2 12 2
3 12 9 2
7 12 2 11 2 11 2 2
5 11 2 11 2 2
5 12 9 9 2 2
8 12 2 11 2 11 2 2 12
6 11 2 11 2 2 12
7 11 2 11 2 2 12 2
5 12 9 9 2 2
8 12 2 11 2 11 2 2 12
8 11 2 12 11 2 2 12 2
2 9 2
11 12 2 11 2 0 2 11 2 2 12 2
2 9 2
7 12 2 11 2 11 2 2
5 11 2 11 2 2
5 11 2 11 2 2
5 11 2 11 2 2
7 11 2 0 2 11 2 2
2 9 2
7 12 2 11 2 11 2 2
7 11 2 11 2 2 12 2
2 9 2
7 12 2 11 2 11 2 2
5 11 2 11 2 2
9 11 2 11 2 11 2 2 12 2
1 2
1 2
1 2
1 2
12 9 1 0 11 2 9 2 12 9 2 12 2
14 9 9 0 9 9 1 11 2 9 9 12 2 12 2
17 0 9 1 0 9 1 11 2 11 2 9 2 9 12 2 12 2
1 2
14 9 11 1 9 1 9 1 0 9 1 11 2 12 2
12 9 0 9 9 9 2 12 2 9 2 12 2
3 13 4 2
4 2 1 9 2
14 9 9 1 9 13 9 0 9 1 0 9 0 0 9
5 9 9 2 11 11
2 9 9
2 11 2
16 9 11 9 7 0 9 11 11 13 1 9 1 0 9 11 2
28 0 9 15 13 1 0 12 9 1 0 11 2 1 0 9 10 9 13 1 9 7 1 9 13 11 0 9 2
12 0 9 13 3 13 2 0 12 13 1 9 2
7 11 11 9 9 11 1 11
7 11 1 11 2 11 2 2
22 9 11 11 3 3 13 1 10 0 9 0 9 1 11 11 11 1 0 7 0 9 2
20 9 11 13 1 0 9 1 11 2 3 15 1 9 13 9 12 2 9 11 2
46 1 9 0 0 9 13 1 15 2 15 9 13 9 1 9 2 4 9 9 9 9 7 0 11 2 0 9 11 1 11 7 9 9 9 9 9 2 15 15 13 13 0 9 1 9 2
15 11 11 1 10 9 13 9 2 15 9 13 1 0 9 2
15 9 11 1 9 13 9 0 0 9 11 1 0 9 9 2
38 1 9 11 2 16 11 13 13 9 2 15 1 15 9 3 13 2 11 2 11 13 2 13 2 16 14 2 13 15 7 0 0 0 9 13 0 9 2
22 1 9 11 0 9 3 1 11 13 7 13 0 9 2 7 13 15 1 9 0 9 2
11 11 13 1 15 0 9 2 3 15 13 2
8 11 7 0 0 9 13 9 2
6 13 15 0 9 9 2
33 13 15 3 1 9 11 7 11 1 9 9 2 7 13 3 1 9 0 9 7 1 15 2 16 9 9 13 3 13 0 9 9 2
22 16 13 1 0 9 9 9 2 13 2 16 4 15 13 13 1 12 2 9 9 11 2
17 11 11 2 15 15 13 1 11 2 13 3 1 9 1 0 9 2
29 1 3 0 9 13 9 1 9 0 9 1 9 0 9 11 2 13 11 9 11 2 15 3 13 9 0 9 9 2
10 9 11 13 1 11 9 1 0 9 2
14 3 13 1 0 13 1 9 11 7 9 11 7 11 2
18 0 9 13 3 2 16 4 13 1 11 2 11 7 11 7 1 11 2
4 0 11 13 9
2 11 11
8 9 9 13 3 13 10 9 2
28 15 13 9 1 0 9 2 0 3 0 1 9 3 2 16 13 10 0 0 9 2 7 16 3 7 1 9 2
29 1 15 2 15 13 10 9 2 15 13 7 9 0 9 0 11 2 15 13 9 9 1 9 0 1 0 2 9 2
25 16 13 1 0 0 9 2 9 15 13 2 15 13 0 13 2 16 4 1 15 9 9 3 13 2
18 1 10 9 15 13 13 1 9 2 7 0 11 15 13 9 1 9 2
5 9 13 3 0 2
11 1 9 13 9 9 9 0 16 1 9 2
21 13 2 14 1 11 2 13 15 9 10 9 1 11 12 2 3 15 13 0 9 2
19 15 15 13 13 1 9 7 1 10 9 13 1 15 13 9 1 9 9 2
9 1 12 9 1 9 9 13 9 2
14 15 13 1 9 7 10 9 13 9 2 13 13 15 2
17 16 4 13 9 1 9 2 13 2 1 0 9 2 9 12 9 2
12 9 1 9 13 13 1 9 1 9 0 9 2
7 10 9 4 3 3 13 2
28 9 13 3 0 2 16 15 13 1 9 10 9 10 9 0 9 3 7 3 2 13 1 15 3 3 10 9 2
20 13 13 7 1 0 9 2 15 10 9 13 15 2 16 3 13 9 7 9 2
8 9 10 9 15 13 0 9 2
9 7 13 13 0 9 1 9 3 2
12 13 15 13 3 1 9 7 1 9 1 9 2
9 1 15 13 9 0 7 0 9 2
4 11 13 0 9
8 11 11 1 0 9 0 9 13
9 11 2 11 2 11 2 11 2 2
28 9 11 11 11 1 9 0 9 0 9 11 13 2 16 10 9 3 13 13 9 0 9 1 3 0 0 9 2
20 11 2 11 13 2 16 1 9 10 9 13 11 12 9 2 0 7 3 0 2
13 13 0 9 13 9 1 9 2 13 11 2 11 2
18 11 1 10 9 4 9 1 0 9 13 1 3 0 9 1 0 9 2
12 9 10 9 1 0 9 11 11 2 11 13 2
40 16 4 15 13 1 9 9 0 2 16 13 15 0 9 2 0 9 15 13 2 16 14 1 9 9 2 7 3 1 12 9 15 13 0 9 2 13 9 11 2
24 9 11 11 2 11 1 9 13 2 16 9 13 0 9 1 3 0 9 4 13 13 0 9 2
25 9 0 9 11 11 11 13 9 16 0 9 2 15 1 1 9 9 1 9 13 9 13 0 9 2
21 11 11 13 2 16 11 13 9 0 9 1 10 9 7 1 9 2 7 1 9 2
14 1 11 15 9 11 13 0 9 0 9 11 1 9 2
15 1 10 9 0 9 15 13 9 11 7 9 9 11 11 2
27 1 0 9 9 11 12 7 12 9 3 13 2 16 1 0 9 15 13 13 7 16 9 2 7 16 9 2
28 1 0 9 1 15 13 1 10 9 0 9 2 1 15 10 9 13 9 2 16 15 1 9 2 1 9 13 2
19 9 2 16 15 10 9 13 1 9 0 9 11 2 11 13 1 9 9 2
19 3 13 1 15 0 0 9 9 9 2 3 16 1 3 0 2 0 9 2
6 9 7 9 1 9 12
7 0 9 0 9 9 0 9
3 9 9 9
1 11
1 11
1 11
1 11
2 9 9
4 4 13 1 9
5 11 2 11 2 2
9 0 9 13 3 13 9 9 9 2
17 9 15 13 3 12 7 10 9 15 13 1 3 16 9 9 9 2
19 1 0 9 11 4 13 12 9 2 1 15 13 12 0 2 9 1 9 2
18 13 1 9 1 9 1 12 9 0 1 0 9 2 0 9 7 9 2
7 3 0 13 3 0 9 2
8 13 15 13 0 9 7 9 2
22 1 9 9 9 9 2 11 11 0 9 9 7 3 0 9 4 3 13 9 9 9 2
8 11 11 4 13 9 0 9 11
5 11 2 11 2 2
25 11 11 4 13 1 9 9 2 15 4 13 1 12 2 9 13 9 1 12 0 9 11 1 11 2
13 13 1 15 9 0 0 9 11 1 11 1 11 2
15 1 9 11 11 2 11 4 13 12 9 1 9 12 9 2
21 13 15 1 0 9 13 2 16 11 11 13 16 9 9 0 9 2 13 11 11 2
15 1 0 9 11 11 2 11 13 9 1 11 1 11 0 2
22 13 2 16 9 1 10 9 11 13 13 0 9 10 9 1 11 1 0 15 0 9 2
27 16 15 1 15 10 9 1 10 0 9 11 13 2 13 9 10 9 13 1 0 9 1 0 9 3 13 2
3 9 0 9
3 9 11 11
8 0 9 13 1 0 9 9 2
18 13 1 15 7 15 2 3 13 1 0 9 9 1 9 0 0 9 2
11 3 4 1 15 13 0 9 1 9 12 2
25 9 13 2 16 3 1 9 12 13 1 12 9 7 1 9 12 4 9 1 9 13 12 9 11 2
8 10 9 13 14 1 0 9 2
18 1 9 10 9 15 4 13 0 9 2 7 1 9 13 3 0 9 2
17 13 3 0 9 0 9 7 0 0 9 13 12 1 10 0 9 2
10 1 10 9 15 7 13 1 0 9 2
36 15 9 9 7 0 9 11 11 15 3 13 2 16 9 9 13 3 0 2 7 3 0 9 7 16 9 7 10 9 10 0 9 4 15 13 2
9 7 4 10 9 1 9 3 13 2
11 3 15 11 13 2 16 9 4 3 13 2
11 3 3 2 7 10 9 13 1 15 0 2
18 0 9 1 10 0 9 3 3 13 9 0 9 7 3 1 0 9 2
14 3 1 12 9 4 13 4 13 0 9 1 0 9 2
14 3 13 1 15 1 9 9 7 3 13 3 0 9 2
16 13 4 13 7 7 9 2 15 4 0 13 1 0 0 9 2
34 13 4 15 13 9 1 9 9 10 2 15 13 1 9 3 7 1 0 12 9 2 7 9 0 9 9 2 15 3 3 13 0 9 2
20 9 9 15 3 3 13 1 0 2 0 9 2 15 3 13 1 0 0 9 2
20 1 15 9 0 9 13 0 9 7 9 2 15 9 13 1 0 9 10 9 2
17 1 12 9 9 13 2 16 15 3 13 9 9 7 13 0 9 2
25 1 10 9 13 9 1 0 9 2 0 2 1 15 13 9 9 9 1 0 9 7 9 9 0 2
23 0 9 4 13 13 0 1 15 7 10 0 9 4 13 1 0 9 2 3 1 0 9 2
25 0 7 13 2 16 1 9 2 3 13 0 9 2 13 3 0 0 9 1 9 0 1 9 9 2
13 1 15 15 0 0 9 2 3 0 2 3 13 2
8 3 15 13 2 13 3 9 2
20 9 11 13 2 16 3 13 1 15 2 13 9 9 9 0 1 15 10 9 2
23 15 4 1 0 9 0 9 3 3 3 13 7 13 13 0 9 2 15 0 9 9 13 2
8 12 13 7 1 11 3 0 2
10 13 15 9 13 0 9 9 1 9 2
13 15 9 13 2 16 13 15 1 1 0 9 0 2
4 0 9 4 13
2 11 2
39 0 9 1 11 2 1 15 9 13 1 9 0 15 1 0 9 9 0 9 2 9 0 0 9 7 9 0 9 2 4 3 1 0 9 9 13 1 0 2
16 0 0 9 13 2 16 10 0 9 13 14 12 5 0 9 2
20 16 4 13 9 0 2 13 4 15 15 13 3 16 12 9 1 12 9 9 2
12 9 13 0 9 0 0 0 9 11 11 11 2
6 11 15 13 2 9 0
2 11 2
20 0 9 1 0 9 13 11 2 16 13 1 9 0 9 0 9 1 10 9 2
39 9 0 9 0 9 1 11 13 0 9 2 16 4 13 10 9 13 0 9 1 11 2 7 13 15 1 0 9 2 16 4 15 13 13 1 9 1 11 2
27 1 9 4 10 9 3 13 3 2 16 4 0 1 9 9 3 13 7 16 4 15 3 13 4 13 9 2
7 0 0 9 7 0 0 9
4 11 11 2 9
9 1 9 1 15 13 1 0 9 2
31 13 15 9 2 13 15 0 7 0 9 2 3 15 9 13 2 15 1 15 3 13 2 3 15 13 7 3 15 3 13 2
56 9 13 1 0 9 3 7 13 9 2 16 16 4 15 0 9 3 3 13 2 7 4 15 15 15 3 13 2 3 1 10 0 9 9 2 15 4 13 13 1 0 9 7 13 2 15 4 13 3 2 3 3 3 2 13 2
39 3 15 3 1 9 9 13 2 16 10 0 9 9 13 1 10 9 0 0 9 2 0 1 9 0 9 2 3 12 9 13 0 2 7 15 1 0 9 2
16 1 10 0 9 13 12 0 9 12 0 9 2 9 7 9 2
7 12 3 0 9 9 9 2
27 16 1 9 0 9 14 12 9 4 3 13 9 0 9 2 3 4 13 4 1 9 0 9 1 9 9 2
20 7 3 4 10 9 13 0 2 12 1 12 13 0 9 1 0 9 15 9 2
19 13 1 15 2 16 13 0 9 3 0 0 9 13 9 14 1 0 9 2
15 3 13 9 2 0 15 9 9 9 2 9 9 11 11 2
9 12 9 1 12 13 3 0 9 2
7 9 1 9 0 9 2 2
29 10 9 7 3 1 9 10 9 13 3 0 2 7 1 9 2 15 3 1 9 9 13 15 0 2 3 13 9 2
16 9 7 9 13 1 15 2 16 4 0 9 13 1 10 9 2
11 3 2 9 13 1 9 10 9 7 9 2
12 9 0 10 0 9 2 10 9 13 4 13 2
25 2 10 9 7 9 0 9 2 15 4 13 13 0 9 7 1 0 9 1 0 7 3 0 9 2
15 1 9 15 13 12 9 2 12 9 9 2 0 9 9 2
39 7 13 1 0 9 2 9 9 13 1 9 2 9 9 1 9 2 7 13 15 1 9 14 12 2 9 1 9 3 13 2 3 15 1 9 13 7 13 2
44 13 2 3 4 13 9 2 16 9 9 13 1 0 0 9 2 16 4 3 3 13 13 1 9 9 9 2 7 9 9 15 3 13 1 0 9 2 7 15 1 9 1 9 2
45 13 9 2 16 15 0 13 1 0 9 15 0 9 10 9 2 7 13 7 1 0 0 9 9 2 16 0 9 13 9 9 9 0 9 2 15 3 2 9 9 1 15 2 13 2
20 9 0 1 10 12 9 2 15 13 13 1 9 9 11 11 2 13 9 11 2
14 9 1 9 15 9 10 9 13 3 3 7 3 9 2
18 9 11 15 13 13 2 13 15 16 9 0 9 2 7 15 13 13 2
31 0 9 13 1 10 9 3 0 2 7 3 1 15 15 13 10 0 9 2 16 4 15 3 13 3 0 9 2 3 9 2
29 3 1 0 12 9 9 9 9 13 12 2 15 13 1 0 9 9 1 0 9 2 9 0 9 2 0 1 9 2
55 2 16 4 15 9 11 13 13 7 13 3 13 14 3 0 9 9 7 3 0 2 7 3 0 0 9 2 13 4 1 0 0 9 0 9 2 16 7 0 7 0 9 10 9 3 2 16 4 15 1 10 9 13 13 2
24 0 11 3 13 2 7 3 3 2 10 0 9 2 16 9 13 14 1 11 1 9 1 11 2
5 9 13 1 0 9
26 0 0 9 2 15 3 13 10 9 2 13 3 1 9 9 9 7 3 10 9 1 9 10 0 9 2
22 1 0 9 1 15 13 3 0 9 0 2 15 13 0 9 7 12 1 12 0 9 2
38 9 11 2 15 15 3 13 16 9 0 9 2 13 16 0 9 9 0 9 11 11 3 4 13 9 2 7 15 1 9 7 9 10 0 9 11 11 2
35 1 9 11 2 15 15 13 1 9 9 9 2 15 13 9 9 11 11 7 1 9 13 9 0 3 1 9 9 2 9 11 2 11 2 2
28 1 15 15 13 13 3 0 11 1 9 0 0 9 9 11 11 2 10 9 15 13 1 9 1 9 11 2 2
26 0 9 9 13 7 3 11 11 2 15 16 0 9 9 13 0 9 0 11 7 11 2 0 12 9 2
18 0 9 0 9 0 11 11 15 13 1 10 0 9 9 9 1 11 2
20 3 1 15 13 1 9 7 10 9 2 3 11 11 2 11 11 7 11 11 2
27 0 9 2 0 9 9 12 9 1 9 11 11 7 0 9 11 11 2 4 1 10 9 13 14 1 9 2
28 1 0 1 0 9 13 11 11 2 0 0 9 1 9 11 13 11 11 2 11 11 2 11 11 7 11 11 2
51 0 9 1 0 9 11 13 11 9 12 9 1 9 9 9 11 11 2 1 0 9 15 16 0 9 13 1 0 9 11 11 11 2 3 1 9 11 11 2 7 1 11 9 11 11 1 0 9 11 11 2
11 1 9 13 7 1 9 7 9 0 9 2
39 3 9 0 9 11 7 0 11 13 12 0 9 2 0 9 11 7 0 9 0 11 2 15 16 10 0 0 9 13 0 11 7 11 2 9 11 11 2 2
14 1 0 9 11 11 13 1 9 9 0 9 1 11 2
25 1 9 0 9 11 2 11 2 11 4 1 0 9 3 13 9 11 7 11 0 7 9 11 11 2
29 0 9 11 11 15 13 0 9 9 0 9 1 11 2 10 0 9 13 0 11 1 11 7 9 1 9 11 11 2
3 2 11 2
5 1 9 2 2 2
8 2 11 12 2 12 2 12 2
14 1 9 7 0 9 1 9 4 13 9 11 2 13 2
22 14 1 0 9 15 13 13 2 16 13 13 9 2 7 7 0 9 13 1 0 9 2
5 0 2 16 0 2
11 13 7 9 2 16 0 9 13 3 0 2
14 13 15 2 16 0 9 15 13 2 16 4 13 3 2
7 3 15 13 1 0 9 2
12 7 15 3 9 0 9 13 0 9 0 9 2
10 1 10 9 4 13 1 9 13 9 2
29 13 4 0 2 16 4 15 15 13 14 9 11 2 7 7 9 11 12 2 15 15 3 1 9 0 9 13 13 2
7 11 12 13 3 0 9 2
11 13 15 2 16 9 1 9 15 9 13 2
32 3 4 15 13 7 9 1 0 7 0 9 2 16 4 13 2 13 15 2 3 0 0 0 9 1 9 11 2 11 7 15 2
14 9 0 9 9 7 9 4 15 13 3 13 15 0 2
7 1 9 11 11 2 0 11
5 11 0 11 13 11
11 0 11 7 11 13 0 9 14 1 0 9
5 11 2 11 2 2
23 12 0 9 0 0 0 9 13 14 1 12 2 9 10 9 0 9 1 10 0 0 9 2
14 1 0 2 11 3 12 9 7 1 11 3 12 9 2
19 9 9 1 12 9 1 9 13 0 9 2 11 1 11 7 11 1 11 2
12 11 13 0 9 9 2 16 9 14 13 9 2
35 0 9 1 9 9 1 11 10 9 3 13 2 16 10 0 9 1 11 2 15 13 0 9 0 0 9 2 13 1 0 9 16 0 9 2
23 11 13 10 0 9 1 0 9 7 13 2 12 2 12 2 2 15 15 13 1 9 9 2
32 9 15 13 9 2 16 0 2 11 2 15 3 13 10 0 9 7 13 1 9 1 11 2 12 2 12 2 2 9 3 13 2
26 1 0 9 3 13 1 9 0 9 2 1 0 9 1 11 3 13 9 9 0 9 1 9 7 9 2
14 0 9 13 1 11 9 2 16 10 9 13 0 9 2
20 7 1 11 13 0 2 11 0 9 7 14 9 3 13 9 11 1 0 9 2
14 0 9 9 13 0 11 2 15 3 1 11 3 13 2
10 0 9 0 9 13 1 11 0 9 2
5 9 1 9 14 13
7 9 0 9 1 0 9 13
2 11 2
23 0 0 9 1 3 0 9 4 13 3 7 3 3 1 0 9 13 1 9 0 9 9 2
15 9 4 15 13 3 13 7 9 4 13 13 7 0 9 2
7 0 9 13 9 0 9 2
26 3 15 13 9 1 12 9 2 7 0 9 15 13 9 1 12 2 7 13 13 9 7 3 0 9 2
15 9 9 2 15 9 1 0 9 13 2 13 3 0 9 2
35 3 4 13 13 1 12 9 0 16 3 2 7 1 0 9 4 13 13 3 1 10 9 2 7 9 15 4 14 13 1 3 0 0 9 2
29 1 0 12 0 9 9 9 2 0 9 9 1 11 7 3 0 9 2 3 10 9 13 1 9 9 7 9 9 2
47 3 15 13 1 0 7 0 9 1 0 9 9 2 15 4 1 0 9 2 0 9 0 1 12 9 2 13 13 1 9 12 1 9 9 1 12 0 16 3 2 3 12 9 1 9 2 2
19 9 9 4 13 9 9 1 11 7 9 9 9 1 11 2 11 7 11 2
26 0 9 9 1 12 9 13 0 9 1 0 9 9 1 9 9 7 1 0 9 9 1 3 12 9 2
17 9 9 3 3 13 1 12 1 0 9 1 11 7 0 9 11 2
20 15 2 3 1 9 1 11 7 1 11 2 3 13 1 9 9 1 12 9 2
23 4 13 0 9 7 9 3 13 1 3 12 9 2 16 0 9 4 0 9 3 3 13 2
13 9 1 0 9 12 3 13 2 13 3 11 2 2
15 3 9 1 0 11 15 3 13 7 13 15 3 10 9 2
18 1 9 9 7 9 4 13 9 9 0 15 9 7 9 1 9 9 2
16 16 15 9 13 2 13 0 9 0 7 0 9 15 3 13 2
10 0 9 0 9 9 9 4 13 9 2
16 0 0 9 3 13 9 1 0 15 9 7 1 0 9 11 2
17 9 0 9 3 13 13 9 2 7 1 9 13 3 0 0 9 2
23 0 0 9 13 9 7 9 2 16 3 4 13 13 9 9 0 2 0 9 7 3 0 2
11 3 9 9 13 3 7 3 9 7 9 2
23 1 9 9 12 15 13 9 2 1 0 9 15 7 13 0 9 7 9 1 0 15 9 2
28 1 9 0 9 9 1 12 9 0 9 15 3 3 13 9 1 3 12 9 7 1 9 12 1 0 12 9 2
10 9 9 15 13 1 9 7 9 9 2
32 0 9 13 9 0 9 2 16 9 4 3 3 13 2 7 0 9 9 9 4 15 0 9 13 13 7 1 0 9 9 9 2
17 9 3 3 13 0 0 9 2 1 9 1 12 9 1 9 2 2
19 0 9 1 11 13 10 9 2 16 9 3 3 1 9 13 1 12 9 2
25 10 9 4 2 3 1 9 9 2 3 13 1 0 9 7 3 3 0 9 2 16 11 9 13 2
4 9 4 13 3
9 11 2 11 2 11 2 11 2 2
12 1 10 9 0 9 4 9 13 1 0 9 2
9 3 4 2 11 2 11 2 13 2
37 1 11 4 13 0 9 1 9 9 3 2 13 10 9 9 0 12 9 2 13 4 13 4 7 1 9 9 2 0 9 2 9 9 7 0 9 2
22 3 2 3 4 9 13 9 2 15 13 13 9 0 9 2 13 3 2 1 9 9 2
11 1 11 13 9 14 0 9 7 9 9 2
8 9 13 1 15 13 14 3 2
16 3 1 15 13 9 9 0 9 0 9 7 15 15 3 13 2
32 1 0 9 0 9 9 13 14 9 1 0 9 2 15 13 12 9 2 14 12 9 2 7 13 3 1 9 9 1 10 9 2
15 1 11 0 0 9 13 2 3 7 3 13 0 9 13 2
9 9 3 13 9 1 9 10 9 2
14 0 9 13 14 1 9 1 9 9 7 1 10 9 2
8 0 13 13 0 0 9 0 2
6 0 13 3 10 9 2
13 0 9 1 9 12 13 0 9 7 13 9 9 2
6 9 13 1 9 9 2
26 0 13 14 9 2 15 1 9 13 2 13 1 15 2 13 1 15 9 7 9 7 15 10 9 13 2
6 9 11 1 11 7 11
2 11 2
38 0 9 1 9 12 9 9 13 9 1 0 9 7 0 9 9 0 2 11 2 1 9 1 0 9 11 11 2 11 2 7 0 0 9 2 11 2 2
21 3 3 13 9 9 11 2 11 11 11 2 13 15 15 0 9 1 0 9 11 2
5 3 13 13 9 9
11 9 0 0 7 0 9 1 11 3 3 13
2 11 11
17 1 0 9 0 9 3 3 13 9 0 0 7 0 9 1 11 2
21 13 15 15 3 9 2 9 2 0 9 2 9 2 9 2 9 2 9 7 9 2
18 1 15 9 0 9 1 0 9 13 3 1 0 9 16 1 9 0 2
14 13 15 1 0 9 2 15 15 13 9 9 0 9 2
19 3 1 0 9 13 9 1 10 0 9 7 9 1 11 3 12 2 12 2
15 3 15 7 10 9 13 3 2 16 3 13 3 16 13 2
38 3 4 1 0 9 9 0 9 13 12 9 2 0 12 0 0 9 2 12 0 9 0 9 1 9 1 9 0 9 7 3 0 9 0 9 1 11 2
12 0 9 15 13 10 9 1 9 0 0 9 2
21 3 3 13 9 9 11 11 1 0 9 9 9 11 2 0 9 1 0 9 2 2
27 10 0 9 11 11 1 15 13 2 16 1 9 1 9 0 9 9 4 3 13 14 1 0 9 1 11 2
29 1 9 0 9 9 4 1 12 2 9 1 0 0 7 0 9 13 3 12 9 1 9 9 1 0 9 1 11 2
16 12 9 4 3 13 2 12 13 7 12 9 1 9 3 13 2
11 3 3 4 0 0 9 13 9 0 9 2
38 9 10 9 13 1 12 9 2 16 1 12 2 9 12 4 1 11 13 10 9 1 12 9 2 9 2 3 1 0 9 14 1 12 9 2 9 2 2
9 3 13 1 15 7 9 0 9 2
40 9 9 15 3 13 1 12 9 2 9 1 12 9 2 0 9 1 12 9 2 9 1 12 9 2 9 1 12 9 2 9 1 12 9 2 9 1 12 9 2
12 9 9 2 9 7 0 9 13 14 1 9 2
38 1 1 0 9 1 9 9 7 1 1 15 2 16 0 9 13 13 14 1 9 0 9 2 9 10 0 9 1 0 9 0 9 11 7 11 3 13 2
25 0 9 2 1 9 2 9 2 1 11 7 11 1 12 2 9 9 12 1 9 1 0 9 9 12
11 0 9 0 11 13 1 9 9 11 1 11
2 11 2
26 0 0 9 2 11 2 2 15 13 12 9 0 9 1 9 0 11 1 0 11 2 13 3 3 9 2
20 13 15 3 0 9 0 11 2 15 7 13 2 16 13 1 9 0 7 0 2
48 9 1 9 9 2 15 15 1 9 12 13 9 14 12 9 2 13 1 0 9 9 0 9 11 11 11 11 11 1 9 9 0 9 7 9 2 11 2 11 11 2 15 13 3 9 0 9 2
19 12 9 13 2 16 1 0 9 1 9 0 9 13 1 0 9 0 9 2
22 9 13 2 16 0 9 4 9 1 9 13 9 3 9 9 12 0 9 1 0 11 2
19 0 9 13 0 9 0 9 1 15 2 16 4 13 1 9 11 0 9 2
35 1 10 9 1 9 13 0 9 2 10 9 11 11 3 13 2 16 13 0 13 2 3 9 11 11 13 10 9 9 7 13 15 13 11 2
4 9 1 9 12
6 9 13 1 9 1 9
9 0 9 9 1 0 11 13 9 9
5 11 2 11 2 2
35 9 1 0 9 0 9 9 1 0 11 9 2 11 11 2 2 0 1 9 0 9 2 13 4 1 0 0 9 11 11 13 9 10 9 2
15 4 2 14 13 0 2 13 15 9 1 12 1 12 9 2
39 1 9 9 13 0 9 3 1 12 9 1 0 9 13 1 9 9 1 12 0 9 2 15 1 0 11 13 0 9 2 1 15 12 9 11 3 3 13 2
19 9 12 2 9 13 9 9 9 2 11 11 2 7 13 9 1 0 9 2
14 9 3 13 12 9 1 0 9 7 1 9 13 9 2
12 15 7 13 1 0 7 13 15 9 1 9 2
11 1 9 7 13 9 9 1 12 12 9 2
16 9 2 11 11 2 15 13 2 16 0 9 13 7 9 13 2
16 13 3 0 9 10 9 2 1 15 4 13 9 3 1 11 2
28 9 0 9 1 11 9 2 11 11 0 9 13 2 16 9 9 1 9 13 2 7 13 1 9 9 10 9 2
25 1 15 13 7 0 2 16 9 13 0 9 2 7 7 15 4 1 9 1 0 11 13 0 9 2
19 1 11 13 9 0 9 1 9 9 2 15 1 11 13 9 9 0 9 2
23 9 9 4 7 13 2 16 4 15 9 13 7 9 4 13 2 16 13 15 1 0 9 2
7 9 9 9 0 9 13 9
2 11 2
38 3 9 1 9 9 9 0 9 3 13 2 3 15 9 1 0 0 9 4 13 2 3 2 1 10 9 2 7 15 4 1 9 13 7 0 9 13 2
12 13 15 11 11 1 9 9 0 9 0 9 2
18 11 13 2 16 3 13 0 13 1 9 9 7 13 15 1 0 9 2
17 1 9 9 13 12 2 9 9 9 7 1 0 9 4 13 9 2
27 1 0 9 4 0 9 0 0 9 7 9 7 9 1 15 13 4 13 9 12 9 1 0 9 9 0 2
25 0 9 4 13 4 13 9 11 1 9 1 15 2 16 3 13 0 9 1 11 2 7 1 9 2
15 13 7 13 1 9 2 15 3 4 13 1 9 0 9 2
5 9 0 9 1 9
2 0 9
6 11 11 2 11 2 2
27 0 9 1 9 11 11 2 0 1 0 9 9 9 2 9 7 9 2 13 3 1 0 9 1 11 11 2
50 9 1 11 2 11 13 0 9 1 0 9 2 16 3 0 1 0 9 9 12 13 1 0 9 1 11 11 9 2 1 15 13 0 9 2 1 0 1 9 0 9 1 11 2 7 9 13 1 9 2
16 9 13 11 1 9 2 16 10 9 13 1 9 0 9 9 2
22 1 0 0 9 13 12 9 2 9 2 15 13 3 1 0 9 1 0 0 9 9 2
18 1 15 13 2 16 0 13 10 0 9 7 13 0 13 9 10 9 2
29 9 2 11 11 1 9 3 13 2 16 0 13 0 9 1 0 9 1 10 9 7 1 0 9 13 7 9 9 2
37 11 2 11 13 1 0 9 1 3 0 9 11 12 2 15 1 9 13 3 12 9 0 9 11 11 2 7 9 4 13 9 13 2 11 13 9 2
48 3 4 15 13 2 16 4 15 13 2 7 13 0 9 1 0 3 16 9 7 9 2 13 1 0 9 1 9 0 2 15 9 13 9 2 16 4 4 13 0 9 1 10 9 1 0 9 2
23 9 4 13 1 9 1 9 2 16 0 9 13 9 1 0 9 9 1 9 1 12 9 2
5 9 11 1 11 13
2 11 2
22 9 9 0 0 0 0 9 2 11 2 11 11 1 0 9 3 3 13 0 0 9 2
21 0 9 1 11 2 3 15 11 13 0 9 1 9 12 2 15 13 1 0 9 2
22 9 0 0 9 13 2 16 0 9 13 13 1 9 0 9 2 7 1 9 0 9 2
3 11 13 9
13 0 9 0 9 13 1 0 9 11 11 1 11 2
27 3 1 11 13 11 11 1 9 0 9 11 2 0 9 13 13 1 15 10 9 14 1 9 9 0 9 2
14 1 12 2 9 4 0 9 11 13 1 0 0 9 2
11 9 3 0 9 13 13 3 1 12 9 2
16 9 9 4 15 13 1 11 2 11 0 9 13 1 12 9 2
10 0 9 0 9 9 13 12 9 9 2
6 9 4 13 1 9 2
38 16 4 0 0 9 1 9 13 9 2 16 0 9 9 13 13 3 9 9 1 9 2 13 11 1 9 11 2 11 13 9 3 0 9 1 9 13 2
12 1 0 9 9 13 1 9 0 9 0 9 2
24 3 11 2 11 13 2 13 1 10 9 1 9 9 1 9 9 1 0 0 9 9 9 9 2
18 0 9 7 13 13 0 9 3 1 9 10 9 1 0 9 2 13 2
15 11 3 13 0 9 1 9 0 9 1 9 12 9 9 2
10 1 0 9 4 9 11 1 9 13 2
21 9 3 1 9 13 0 2 0 9 2 15 13 13 0 9 10 9 1 9 9 2
13 1 9 4 15 13 13 1 9 13 3 9 9 2
3 2 11 2
5 11 15 13 0 9
4 11 11 2 11
12 0 9 1 11 13 2 16 11 3 13 9 2
24 12 1 0 9 13 7 10 9 2 16 9 3 0 9 13 10 9 1 0 9 1 0 11 2
20 11 3 3 13 0 7 16 4 15 3 9 13 2 13 4 13 1 0 9 2
25 7 16 4 2 15 13 3 0 2 10 0 9 2 0 9 2 3 13 0 9 7 13 13 9 2
31 13 15 7 0 0 9 1 9 9 9 7 9 2 0 1 9 1 9 0 9 1 0 9 11 2 11 2 11 7 11 2
30 1 9 0 9 11 15 11 1 9 9 13 3 10 9 2 15 13 3 7 3 13 2 16 15 9 1 9 9 13 2
23 16 3 9 3 0 9 2 15 13 1 0 9 7 0 9 2 0 9 7 3 0 9 2
37 15 7 13 2 16 0 0 9 2 16 9 9 2 11 2 9 2 9 2 9 2 11 2 0 9 0 13 7 9 2 11 13 7 13 0 9 2
17 3 2 15 4 3 13 7 13 1 0 9 1 9 1 0 9 2
43 0 9 3 13 10 9 9 1 10 9 13 2 3 7 3 2 16 9 9 13 14 9 11 7 16 15 7 13 3 13 0 9 9 7 13 15 0 9 1 9 0 9 2
18 11 1 0 12 9 13 3 9 9 2 3 0 9 1 3 0 9 2
15 13 7 2 16 13 3 12 0 0 9 2 3 0 9 2
8 13 15 15 9 1 0 9 2
11 9 13 3 1 11 2 1 9 9 11 2
19 13 15 1 9 3 12 9 2 15 1 9 0 9 3 13 1 0 11 2
19 9 15 13 13 12 1 15 2 11 11 2 7 15 13 9 1 9 0 2
16 12 9 9 1 9 11 14 13 13 0 11 11 11 0 9 2
18 16 11 13 1 9 0 9 1 10 9 2 3 14 13 0 9 9 2
21 13 7 2 16 3 3 13 1 9 0 9 2 7 16 9 10 0 9 7 9 2
44 0 13 2 16 10 9 13 1 9 0 0 9 2 15 13 9 0 9 7 0 9 3 13 2 7 3 3 13 3 2 16 3 15 13 3 7 16 11 3 3 13 10 9 2
30 16 3 4 11 1 9 10 0 9 9 11 11 13 1 0 9 1 9 0 11 2 3 1 0 9 13 1 0 9 2
20 9 2 16 1 9 13 9 13 7 13 0 9 9 2 3 13 15 0 9 2
24 1 9 0 9 13 1 9 9 7 1 9 1 0 11 9 2 15 15 13 1 9 0 9 2
18 11 11 7 11 0 1 11 13 2 11 11 15 13 1 9 1 11 2
15 0 0 11 13 11 11 2 15 3 13 3 10 0 9 2
22 0 12 9 13 9 0 0 9 1 11 7 1 11 15 13 3 9 1 9 7 9 2
19 16 1 9 13 0 9 2 1 0 9 9 9 13 1 9 9 0 9 2
13 11 11 1 9 2 1 9 2 13 3 0 9 2
7 9 13 1 12 2 9 2
6 2 11 2 9 11 11
4 11 1 12 9
1 9
17 9 2 0 0 9 11 11 3 13 9 1 0 9 0 0 9 2
35 3 9 9 2 1 9 2 9 2 0 9 2 2 2 2 2 3 0 9 13 1 10 9 15 15 2 13 3 3 1 10 9 0 9 2
15 1 9 15 1 15 3 13 0 9 1 0 9 12 9 2
23 11 15 3 13 2 16 13 10 9 13 3 2 16 4 9 1 10 9 13 9 0 9 2
53 0 9 15 13 3 2 0 9 13 3 0 2 9 1 9 9 13 3 0 9 1 9 14 0 2 15 15 13 1 0 2 3 0 9 2 13 13 9 0 9 2 9 2 15 13 1 15 1 0 9 2 2 2
8 13 15 1 15 13 1 9 2
45 9 13 12 0 9 2 16 12 9 13 13 3 1 0 9 9 2 11 13 9 3 16 0 0 9 2 2 0 9 1 0 9 2 9 7 9 13 0 9 3 13 1 10 9 2
28 12 9 7 12 9 13 0 9 9 2 16 0 9 9 1 10 0 9 13 9 9 9 2 0 7 3 0 2
20 0 9 2 0 10 9 2 13 1 9 0 9 15 0 2 14 7 3 0 2
34 16 0 1 10 9 11 13 13 1 0 0 9 2 9 1 0 2 0 7 0 9 13 3 1 9 0 9 7 10 9 11 1 11 2
28 16 9 13 1 12 9 3 16 1 0 9 2 13 1 9 3 0 2 9 0 9 15 3 14 3 3 13 2
34 3 13 0 9 1 10 9 0 9 9 2 10 0 9 4 15 9 3 13 2 13 7 1 9 2 16 10 0 9 3 11 3 13 2
13 0 0 9 0 9 15 13 7 1 9 0 9 2
26 0 9 13 3 1 12 9 2 3 0 9 15 13 14 9 7 10 9 2 7 7 0 7 0 9 2
41 13 15 3 2 16 1 9 2 3 11 13 15 12 9 2 15 13 9 11 2 1 11 3 13 1 9 11 2 11 11 9 2 13 9 9 7 11 11 13 9 2
68 1 0 9 13 15 7 15 2 14 2 11 11 2 3 1 10 9 13 11 11 9 1 9 2 13 13 0 9 2 11 1 11 2 9 13 9 9 2 9 7 13 1 15 9 7 11 11 15 13 1 9 2 1 9 13 9 0 9 2 16 16 15 12 9 13 2 2 2
2 11 11
13 11 11 2 12 9 2 9 2 9 1 0 9 2
16 13 11 11 7 11 2 0 11 11 7 11 1 11 2 9 2
15 9 2 13 0 11 2 9 11 2 2 12 2 13 11 2
33 11 11 2 11 2 7 11 11 2 11 2 1 9 0 12 9 2 1 15 15 9 1 11 3 13 0 9 0 9 9 1 0 11
2 9 9
4 0 11 7 11
6 0 0 9 9 11 11
2 11 2
30 0 0 9 1 12 9 9 11 11 13 7 1 0 9 0 9 0 9 7 13 15 12 9 9 1 9 12 9 9 2
31 1 9 1 11 2 11 7 11 13 10 9 7 1 12 2 9 9 11 1 11 7 10 9 13 0 0 0 9 12 9 2
14 0 9 0 9 13 0 9 1 9 11 11 1 11 2
21 0 9 9 13 0 9 12 9 7 13 3 16 0 9 0 9 1 9 0 9 2
31 1 0 9 9 1 12 9 15 13 9 9 11 1 11 2 12 2 2 15 13 0 9 11 1 11 7 9 11 11 11 2
23 0 0 9 11 11 15 13 9 9 12 9 2 7 12 9 1 0 9 12 9 0 13 2
18 11 11 15 13 3 3 1 0 9 9 9 9 7 11 11 1 11 2
17 3 15 7 13 13 1 0 9 2 16 0 9 13 0 9 11 2
15 0 9 1 0 9 15 13 0 9 1 9 9 11 11 2
23 13 15 13 2 3 16 1 9 1 11 2 1 0 9 2 16 10 0 9 13 12 9 2
20 3 15 3 13 11 11 2 12 2 2 15 3 3 11 13 1 9 1 11 2
14 0 0 9 1 12 9 12 13 1 11 11 11 11 2
16 1 9 1 12 9 13 11 11 0 9 1 11 11 1 11 2
2 0 9
2 11 2
4 9 2 11 2
2 11 2
1 9
15 9 9 9 1 11 2 11 11 2 11 11 12 2 12 2
18 9 9 0 9 11 11 11 13 1 9 0 9 11 11 11 7 11 2
22 0 9 13 3 1 11 1 9 9 9 11 11 11 1 0 9 0 9 9 11 11 2
27 9 9 2 10 9 13 9 11 11 2 15 13 3 0 9 11 11 7 9 0 2 0 7 0 0 9 2
5 9 11 11 2 11
6 11 2 9 1 0 9
1 11
4 11 11 2 11
36 10 9 13 3 1 12 2 9 2 13 9 1 0 9 11 2 9 2 15 4 3 13 16 0 9 2 7 3 13 3 7 9 0 9 9 2
19 13 15 1 9 2 16 1 12 9 1 9 4 1 9 13 14 0 9 2
17 9 13 1 9 3 3 9 2 16 16 4 13 9 1 9 9 2
30 9 1 0 0 9 15 7 1 0 0 9 2 15 13 1 9 1 0 9 0 9 13 9 1 9 2 13 9 9 2
18 0 9 9 2 15 15 3 13 1 0 12 9 2 13 3 0 9 2
18 13 15 2 16 9 15 14 3 13 9 2 7 3 15 13 1 0 2
18 9 0 9 13 0 9 2 9 9 7 13 0 9 9 9 1 9 2
9 1 9 13 0 2 3 0 9 2
7 9 13 3 0 7 0 2
31 16 0 9 1 11 13 3 12 12 9 2 1 0 9 2 3 13 0 9 3 0 9 2 15 13 1 12 7 12 9 2
14 9 13 7 2 3 1 9 7 9 2 3 0 9 2
34 9 1 9 15 1 0 12 9 0 9 13 1 12 9 9 2 1 0 12 9 2 2 2 7 9 9 2 9 7 0 9 3 13 2
14 9 13 9 9 0 9 9 1 9 7 0 9 9 2
6 9 0 9 13 0 2
14 1 0 9 4 13 9 0 7 13 7 12 0 9 2
14 1 9 13 12 9 9 2 15 13 9 1 0 9 2
21 0 9 7 13 2 16 1 9 0 0 9 1 0 0 9 13 9 3 12 9 2
18 1 0 9 1 0 9 13 0 9 1 9 1 9 7 0 0 9 2
9 13 0 9 0 9 9 7 9 2
7 0 9 13 1 0 9 2
13 9 1 9 9 9 1 9 7 9 13 0 9 2
14 1 0 9 0 9 1 15 13 13 3 1 9 12 2
17 9 7 4 3 13 7 9 7 10 9 13 1 9 1 0 9 2
16 9 3 13 2 16 4 3 1 9 13 3 0 9 1 9 2
12 9 3 13 0 13 9 0 9 1 9 9 2
14 13 9 9 2 3 3 16 0 0 9 0 9 9 2
19 4 3 13 2 10 9 13 9 2 7 15 2 1 15 15 4 3 13 2
6 9 3 13 3 9 2
11 1 9 9 15 1 12 9 13 12 9 2
32 3 0 1 15 15 13 1 9 0 9 9 2 7 16 9 13 3 0 9 2 13 15 10 9 1 15 9 13 15 3 3 2
20 14 3 15 9 11 11 13 13 9 0 0 9 7 13 0 9 1 0 9 2
20 13 9 11 2 1 0 9 2 15 13 1 9 0 11 2 7 3 7 11 2
18 0 0 9 4 13 4 13 1 9 3 1 9 2 3 1 0 9 2
11 0 9 1 9 9 11 13 1 9 9 12
2 11 2
24 9 11 0 9 1 0 7 0 11 7 9 0 0 9 4 1 0 9 13 1 9 9 12 2
24 1 0 9 1 0 9 9 7 9 11 11 15 13 9 9 11 1 0 7 0 11 11 11 2
22 9 11 1 9 13 2 16 0 9 13 0 9 0 0 9 2 1 15 9 11 13 2
22 13 15 3 2 16 0 9 13 0 9 3 3 2 16 10 9 3 3 13 3 0 2
19 1 9 1 0 9 16 3 11 2 11 2 7 7 11 2 13 11 11 2
17 9 7 1 10 9 13 3 1 0 9 1 11 7 3 7 11 2
29 9 9 11 13 16 9 1 9 9 7 9 3 2 0 9 0 9 11 2 11 11 2 9 11 7 0 9 11 2
34 0 9 0 9 11 1 11 13 1 0 9 9 9 1 9 9 1 0 9 1 0 9 2 7 15 7 1 0 9 7 1 0 9 2
30 1 9 11 1 0 7 0 11 4 13 3 12 9 9 2 1 15 7 3 0 9 4 13 1 9 9 1 0 9 2
4 0 9 1 9
3 0 11 2
20 16 0 1 0 11 13 9 9 11 1 11 0 9 1 9 2 15 13 9 2
25 9 9 11 11 3 1 9 9 9 13 2 16 9 10 9 13 1 12 9 1 9 9 0 9 2
11 0 9 9 15 13 1 12 9 9 3 2
7 9 11 13 3 12 9 2
18 3 9 10 0 9 13 1 9 2 3 1 11 7 1 9 0 11 2
8 9 13 10 9 1 9 9 2
12 3 10 9 1 9 13 1 9 3 9 9 2
31 1 12 2 9 13 9 1 0 9 0 0 9 10 9 2 3 0 9 2 16 13 0 9 2 9 2 9 7 9 9 2
9 10 9 3 13 0 9 9 9 2
9 10 0 9 13 7 9 7 9 2
12 0 9 9 9 15 13 1 12 7 12 9 2
23 3 9 9 1 10 9 13 9 0 9 1 9 7 0 9 13 1 9 2 3 1 11 2
6 9 9 1 9 15 13
30 0 9 2 3 1 0 11 2 7 0 9 9 1 11 7 11 13 2 16 9 9 2 9 2 1 9 13 13 9 2
21 9 10 9 2 15 15 13 3 1 9 7 3 1 0 1 9 2 3 3 13 2
42 16 13 10 9 0 9 0 11 2 1 11 15 9 0 9 2 9 2 7 0 9 1 9 13 13 9 3 3 1 10 9 2 13 3 0 9 0 9 9 1 12 2
23 3 1 0 9 15 1 11 13 9 1 10 9 1 9 1 0 9 0 9 1 12 9 2
8 9 4 13 7 1 0 11 2
17 0 9 13 1 9 1 9 10 9 1 12 1 12 9 1 9 2
11 9 1 11 15 13 1 0 9 1 9 2
27 9 1 9 4 13 7 0 9 10 9 1 9 2 12 1 0 9 1 9 9 2 1 11 7 1 11 2
14 13 4 3 12 9 9 11 1 0 11 1 0 11 2
9 0 9 9 1 11 13 0 9 2
13 9 0 9 1 9 11 13 1 9 2 7 13 9
9 11 2 11 2 11 2 11 2 2
21 0 9 15 13 13 9 0 9 1 0 9 2 15 1 0 9 13 0 9 11 2
46 13 15 1 15 2 9 0 9 2 0 15 10 9 1 0 7 0 9 9 11 2 13 13 2 16 9 0 9 13 0 9 9 1 9 0 0 9 2 15 13 0 9 0 9 9 2
86 1 1 15 2 16 0 9 0 9 13 1 9 7 9 1 9 9 7 7 9 0 9 9 1 0 9 2 15 9 0 9 13 0 15 13 3 16 9 2 15 9 0 9 13 1 0 0 9 0 9 0 9 2 0 9 0 9 15 13 7 13 3 2 16 4 1 0 0 9 9 0 9 1 9 9 7 9 9 0 9 13 0 9 0 9 2
16 13 1 9 3 0 9 13 1 0 9 9 7 11 11 11 2
13 7 3 1 0 9 11 11 10 9 0 9 13 2
19 1 11 3 13 2 16 13 3 9 0 9 2 7 3 13 1 9 9 2
28 3 3 16 0 13 15 3 14 0 9 1 9 2 13 7 13 2 16 10 9 13 0 7 3 3 13 0 2
47 9 11 11 2 11 2 11 13 2 16 16 13 1 9 0 9 11 1 0 9 1 9 9 2 13 15 3 1 1 15 2 16 13 1 0 9 0 9 3 16 9 1 9 9 16 9 2
4 3 1 9 12
6 11 13 13 9 1 9
5 11 2 11 2 2
12 0 9 13 9 0 9 2 0 1 0 9 2
24 9 13 3 13 1 9 2 0 9 11 2 15 9 13 2 15 7 13 1 9 9 11 13 2
15 0 9 7 1 9 3 15 13 2 15 1 15 13 9 2
17 11 15 13 1 9 14 1 9 2 3 4 9 9 13 0 9 2
32 9 9 9 2 11 2 11 13 9 1 15 2 16 0 9 13 4 1 0 9 1 9 0 9 1 9 1 9 1 9 13 2
25 16 11 13 9 2 11 1 0 9 9 2 9 4 1 9 9 1 0 9 13 14 1 12 9 2
8 11 11 3 13 7 1 11 11
2 9 11
4 9 1 0 9
19 9 1 9 9 1 0 9 0 9 13 1 9 0 9 13 1 0 9 2
15 9 4 13 1 0 9 16 0 9 9 3 12 9 9 2
21 1 0 11 11 15 7 13 2 16 9 10 9 13 0 7 9 1 9 13 0 2
11 9 9 4 15 3 13 14 12 9 9 2
19 9 4 7 1 9 13 1 12 9 9 0 9 2 15 15 4 3 13 2
36 9 0 9 3 13 2 16 4 9 9 10 0 9 13 1 12 9 9 2 7 15 13 2 16 9 4 13 13 1 0 9 9 10 0 9 2
16 1 11 2 11 4 15 0 9 13 13 1 9 12 0 9 2
3 2 11 2
4 9 13 0 9
5 11 2 11 2 2
9 0 9 4 13 1 11 1 11 2
21 9 1 9 12 7 12 9 15 9 13 12 9 2 9 1 0 9 7 9 11 2
13 9 13 0 9 9 1 12 9 2 3 15 13 2
22 0 1 12 9 4 1 9 3 3 3 13 2 7 7 4 3 1 9 13 1 9 2
7 10 9 4 13 1 9 2
3 9 1 0
1 9
2 11 11
19 1 3 12 12 0 2 15 15 1 0 9 13 10 9 2 0 9 13 2
7 15 9 2 15 13 9 2
22 10 9 3 13 9 2 7 14 14 3 0 9 1 15 13 9 2 7 3 3 9 2
33 0 0 9 2 15 13 2 3 13 2 3 13 0 9 0 13 9 2 1 15 12 9 1 0 9 13 1 12 7 12 9 3 2
5 3 13 0 9 2
41 7 16 13 3 7 3 0 13 9 0 9 2 15 13 3 0 9 9 2 1 15 7 3 9 13 0 7 0 9 9 2 13 3 9 2 3 4 0 13 13 2
6 15 0 3 4 13 2
42 0 0 9 3 13 1 15 2 16 0 9 1 9 1 9 4 3 13 3 13 1 10 0 9 2 16 0 9 3 3 0 13 3 3 0 9 13 15 1 0 9 2
8 13 7 3 3 1 9 0 2
21 1 0 9 2 1 0 9 14 3 0 2 13 15 9 0 2 15 0 0 11 2
8 1 9 9 13 9 3 0 2
25 13 3 1 12 9 0 9 9 2 3 0 9 2 1 15 13 0 9 14 0 0 9 1 9 2
23 13 3 7 3 9 0 0 9 2 3 9 2 15 15 13 7 13 3 14 1 0 9 2
19 13 3 9 2 15 15 13 0 9 1 9 2 1 0 9 0 9 9 2
12 7 13 3 3 0 9 1 0 9 0 9 2
30 10 9 0 2 7 3 0 9 1 15 2 15 13 9 9 1 0 9 2 16 13 3 9 2 16 10 9 13 0 2
32 13 10 9 9 7 1 15 9 9 2 0 3 3 7 9 13 15 10 9 2 15 13 10 9 2 15 4 15 0 13 13 2
8 15 15 3 1 9 9 13 2
19 1 0 9 13 0 9 3 3 0 9 2 1 15 13 0 13 0 9 2
33 1 9 7 3 13 9 7 3 0 9 2 15 4 13 15 7 10 9 13 3 9 2 7 13 3 16 9 7 9 7 9 9 2
21 0 13 3 1 10 0 9 12 9 2 0 9 7 0 9 15 13 1 0 9 2
12 13 9 1 0 13 3 3 9 0 0 9 2
16 1 10 0 14 2 9 13 15 7 9 1 9 7 1 9 2
17 13 0 14 13 15 1 0 9 7 13 15 1 9 1 0 9 2
7 11 2 11 1 0 9 9
2 11 2
26 0 9 0 9 11 2 9 2 0 1 0 9 11 0 0 9 13 3 0 9 9 9 11 11 11 2
14 13 15 0 9 1 11 7 0 0 9 1 9 11 2
14 9 11 2 11 1 0 9 13 1 10 9 3 0 2
33 13 2 10 9 13 9 1 11 1 9 0 0 0 9 2 7 13 2 16 15 1 0 9 13 16 1 9 0 0 9 0 9 2
3 1 9 9
1 9
24 9 2 13 15 1 11 11 2 3 3 3 13 1 0 9 11 2 0 9 11 9 11 11 2
5 0 13 9 9 2
6 9 9 0 7 0 2
16 7 9 0 0 9 2 13 1 9 16 9 9 7 10 9 2
11 0 0 9 11 11 10 9 9 3 13 2
20 13 15 0 9 10 9 1 12 0 9 2 15 16 9 9 3 13 1 9 2
27 11 11 2 11 11 7 11 11 13 0 0 9 7 0 1 15 1 0 9 13 7 0 7 0 9 9 2
15 16 15 15 3 3 13 2 3 15 3 3 13 1 9 2
20 3 4 13 13 9 9 9 2 7 1 9 1 0 0 9 1 9 13 13 2
17 0 12 0 9 2 9 11 11 7 11 11 2 13 9 3 3 2
54 11 11 10 0 9 9 13 1 9 9 11 11 2 12 2 12 2 2 7 13 7 9 9 11 11 2 12 2 12 2 2 11 11 2 12 2 12 2 2 7 3 1 9 9 0 9 11 11 2 0 2 12 2 2
30 11 13 9 1 9 7 10 9 2 1 15 13 9 7 9 11 11 7 9 11 11 2 1 0 9 13 16 0 9 2
40 0 2 3 0 9 2 7 3 0 9 11 11 11 13 1 9 9 11 2 15 13 1 9 9 0 7 0 2 16 4 1 9 1 10 9 13 3 3 3 2
15 3 3 11 13 9 9 11 11 11 11 7 0 0 11 2
11 10 3 0 9 7 13 1 9 1 9 2
14 9 0 0 9 0 9 13 10 9 0 9 12 9 2
5 13 0 9 11 11
9 3 3 13 0 0 9 11 11 2
15 1 10 9 13 0 9 0 9 1 9 10 9 1 11 2
20 13 15 3 9 9 3 2 16 10 0 9 13 9 0 0 9 1 0 9 2
48 13 15 12 2 9 12 1 11 2 13 1 11 7 1 0 9 15 1 9 9 13 0 9 2 13 3 1 9 11 7 11 2 1 15 1 9 3 13 2 16 15 1 1 0 9 13 13 2
35 0 0 9 10 0 9 2 12 2 15 13 1 9 9 0 9 2 15 2 3 16 3 0 0 9 2 13 3 1 0 0 9 7 9 2
41 1 9 0 9 0 9 2 12 2 13 1 11 0 9 11 11 2 1 15 3 13 7 1 9 11 2 2 2 2 2 12 2 1 9 7 9 1 12 0 9 2
31 1 0 9 0 15 9 2 2 12 2 3 13 3 0 9 0 9 7 0 9 2 0 0 9 2 0 9 7 0 9 2
37 0 9 9 15 13 7 1 10 0 9 0 9 2 12 2 2 15 0 9 11 11 2 1 9 11 11 2 13 1 0 12 9 1 10 0 9 2
32 0 9 15 13 0 9 1 9 2 0 9 7 0 9 2 15 13 7 1 9 1 0 9 2 3 15 3 3 13 1 9 2
48 9 1 0 0 9 7 10 0 9 13 0 9 11 2 9 2 11 2 12 2 2 15 1 0 0 9 13 11 11 7 11 11 7 15 9 3 13 0 9 0 1 9 9 1 0 0 9 2
23 11 11 13 1 9 2 15 15 1 9 0 9 13 0 9 2 0 9 7 3 0 9 2
28 13 0 9 7 0 9 2 7 3 13 1 0 9 2 9 10 9 4 1 1 0 9 9 3 3 3 13 2
3 2 11 2
5 0 0 2 2 2
8 2 11 12 2 12 2 12 2
13 11 2 11 13 2 16 9 14 13 3 0 9 2
11 3 15 7 3 13 2 13 15 9 0 2
19 9 9 9 2 12 2 12 9 2 1 0 0 9 1 9 12 13 0 2
9 9 13 9 1 9 9 1 11 2
28 9 13 14 9 15 2 15 13 9 9 9 7 9 1 15 1 0 9 2 1 15 15 13 13 9 9 9 2
6 1 9 11 11 2 11
2 0 9
1 9
18 9 0 9 2 11 11 2 11 11 12 2 12 2 12 2 12 2 2
3 13 4 2
4 2 1 9 2
7 1 11 13 7 9 1 9
16 9 9 1 9 0 11 15 1 11 11 13 1 9 12 9 9
2 11 11
37 0 9 1 9 9 1 12 2 9 9 0 9 1 11 1 11 1 9 11 2 12 2 11 11 2 9 11 2 11 2 13 1 0 9 11 11 2
18 13 15 1 9 16 0 9 7 9 1 10 9 1 9 0 9 9 2
17 3 0 2 0 9 15 13 3 1 9 9 0 9 1 15 13 2
14 9 10 9 13 1 9 9 9 0 11 3 1 11 2
10 9 13 2 0 2 1 0 12 9 2
26 13 15 12 9 2 9 11 7 9 11 11 2 15 3 13 13 0 0 9 1 0 9 1 0 9 2
8 15 13 15 1 12 12 9 2
11 13 15 1 9 0 9 1 9 7 13 2
9 15 0 13 3 9 1 0 9 2
20 11 11 13 1 9 12 1 0 11 7 3 13 3 9 11 2 13 7 11 2
20 3 13 0 9 11 2 3 3 3 2 16 4 13 7 13 2 16 15 13 2
15 11 1 11 13 10 9 1 11 7 13 15 3 0 9 2
16 11 13 9 9 1 11 7 1 11 2 13 1 11 7 11 2
12 1 15 7 15 1 15 3 13 1 9 9 2
19 3 4 13 9 0 0 9 2 7 1 15 3 0 9 1 9 0 9 2
20 0 9 15 15 13 7 13 15 3 13 0 9 2 16 0 9 13 15 0 2
19 0 11 13 0 3 3 1 10 9 2 16 9 3 13 1 12 12 9 2
13 1 15 1 15 13 2 13 15 9 9 7 9 2
12 16 13 14 0 2 16 10 9 13 0 9 2
17 13 2 16 13 15 3 3 0 9 2 7 3 15 1 15 13 2
24 3 13 9 3 1 9 1 9 7 3 3 7 13 10 0 9 1 9 2 1 9 10 9 2
8 3 3 15 13 1 0 9 2
18 13 9 11 7 11 7 13 15 1 9 13 2 3 3 3 13 13 2
6 13 3 3 0 9 2
9 0 9 13 3 12 2 12 9 2
9 9 9 7 9 2 9 3 0 2
24 3 13 13 0 9 2 7 10 9 13 3 0 7 3 13 7 13 2 16 15 1 15 13 2
12 3 13 14 9 2 7 7 9 7 9 9 2
7 3 15 13 1 9 9 2
19 9 4 13 0 9 11 11 11 11 2 15 4 13 1 12 9 1 11 2
13 15 13 2 13 9 9 7 13 9 1 0 9 2
18 9 2 9 7 9 2 0 9 2 0 9 2 0 9 2 0 9 2
12 13 1 15 14 9 1 9 7 0 0 9 2
7 9 13 0 13 12 9 2
10 1 0 13 1 0 9 3 12 9 2
9 1 10 9 3 3 13 10 9 2
7 15 4 13 10 0 9 2
5 13 13 9 15 2
12 9 13 10 0 9 7 13 9 2 15 13 2
7 13 9 7 3 13 0 2
21 1 9 1 9 4 3 13 1 9 15 2 16 0 9 12 9 12 12 13 0 2
19 1 9 9 9 3 13 11 11 2 0 9 11 7 11 2 0 2 9 2
11 13 4 15 13 2 16 15 13 15 0 2
6 1 11 13 0 9 2
8 14 1 15 13 7 10 9 2
8 1 11 4 13 9 1 9 2
27 13 15 7 13 12 9 1 9 7 13 9 2 16 1 1 0 9 9 7 9 3 3 15 15 3 13 2
6 13 3 10 9 9 2
7 15 4 13 13 1 9 2
12 3 15 2 7 13 9 2 16 9 15 13 2
20 9 13 3 0 2 16 16 13 10 0 9 9 2 7 4 15 15 13 13 2
9 1 12 9 13 0 9 1 11 2
10 16 4 13 9 2 13 4 1 15 2
5 1 11 3 13 2
8 13 4 15 1 10 9 3 2
6 3 15 15 15 13 2
11 13 4 3 0 9 16 3 11 7 9 2
16 13 2 16 13 3 0 9 13 2 16 4 13 14 9 9 2
6 13 3 3 0 9 2
10 11 2 11 2 11 1 11 7 11 2
11 12 13 3 7 13 15 9 1 0 9 2
16 15 3 13 1 9 9 2 7 1 9 2 16 13 15 0 2
7 16 4 15 9 3 13 2
23 16 13 12 9 2 11 7 11 2 15 13 0 9 12 0 9 2 7 3 13 10 9 2
15 13 15 0 9 11 2 1 10 0 9 13 3 10 11 2
18 3 13 15 13 2 13 15 0 2 16 4 15 15 13 13 0 9 2
9 11 1 9 13 3 3 0 9 2
9 1 0 9 1 11 13 0 9 2
10 15 15 13 1 9 9 3 1 9 2
13 9 13 12 1 9 2 15 15 3 13 13 9 2
32 13 15 3 2 16 13 15 9 1 9 9 2 7 3 1 9 1 11 13 9 11 2 1 9 1 9 2 3 4 13 15 2
21 15 2 16 9 11 9 13 9 1 9 11 2 13 0 9 3 15 13 0 9 2
9 3 3 3 13 1 0 9 9 2
6 15 13 0 0 9 2
4 3 15 13 2
11 13 15 9 9 1 0 9 7 0 9 2
23 0 9 13 9 3 9 7 1 0 9 3 13 9 2 15 13 1 11 7 0 0 9 2
15 13 15 3 1 15 3 0 9 2 16 16 4 13 0 2
13 3 13 0 2 16 0 11 1 9 11 13 9 2
13 13 1 15 9 2 14 13 15 0 9 1 0 2
10 3 4 13 2 7 3 15 3 13 2
18 13 4 15 2 16 16 3 13 10 9 2 3 1 15 3 3 13 2
12 7 1 11 9 13 9 2 9 13 1 9 2
7 9 2 9 2 7 0 9
9 0 9 9 3 13 13 1 0 9
2 11 11
11 14 9 10 9 13 3 1 9 0 9 2
13 1 0 9 13 9 2 16 9 9 13 3 0 2
4 13 15 3 2
13 3 13 13 2 16 4 9 1 10 9 13 0 2
15 9 1 0 9 13 3 0 2 13 3 7 3 3 0 2
15 9 1 15 2 7 1 0 11 2 15 13 1 12 9 2
13 13 15 3 3 1 0 0 9 15 10 0 9 2
18 9 7 3 13 3 0 0 9 0 9 2 10 9 13 3 0 2 2
25 1 15 0 9 11 4 7 9 13 1 0 0 9 2 3 9 15 13 9 1 0 0 9 2 2
8 14 1 15 15 3 3 13 2
7 9 9 16 9 3 13 2
14 9 7 13 2 16 3 7 3 1 15 13 13 13 2
7 10 9 9 13 13 9 2
7 9 1 10 9 13 0 2
12 13 3 13 1 9 9 2 7 3 1 9 2
21 11 11 2 9 9 9 0 9 1 9 9 13 2 16 15 13 13 3 12 9 2
9 16 9 13 0 9 9 2 13 2
28 3 0 3 13 2 16 9 9 13 1 10 9 3 13 15 0 9 9 2 1 0 9 14 1 0 0 9 2
14 13 15 0 3 2 16 4 10 9 13 0 2 0 2
17 13 7 0 15 13 2 16 10 9 13 1 10 9 3 3 13 2
12 15 9 4 3 13 0 9 2 0 0 9 2
7 15 15 9 9 3 13 2
12 9 13 10 9 13 7 3 15 1 9 13 2
9 1 9 13 3 0 13 0 9 2
8 13 15 1 15 3 0 9 2
35 16 3 1 0 9 1 12 9 0 0 9 13 13 14 12 12 9 2 3 12 12 9 1 10 13 13 1 9 2 9 7 9 0 9 2
26 9 13 3 1 12 9 0 2 13 15 2 16 9 1 9 0 9 13 0 16 0 9 1 9 2 2
10 3 1 12 9 9 15 9 9 13 2
12 1 15 2 16 13 7 13 13 3 9 9 2
14 1 0 9 13 3 0 2 7 9 9 1 9 13 2
15 9 13 2 16 9 1 0 9 3 13 2 16 15 13 2
8 0 9 4 13 1 0 11 2
22 9 13 3 0 9 1 11 1 9 12 7 12 2 15 3 13 9 9 7 9 9 2
17 1 9 9 1 9 12 7 1 9 12 13 1 0 11 9 9 2
8 1 0 9 15 9 3 13 2
11 1 9 4 9 1 0 9 13 7 3 2
13 3 1 15 15 1 0 9 13 10 0 9 9 2
15 13 15 13 7 0 9 0 9 2 15 13 0 9 9 2
24 1 11 7 9 9 9 13 3 3 12 9 7 9 1 10 9 13 13 3 0 9 10 9 2
6 13 4 15 7 13 2
15 15 1 15 3 3 13 2 16 13 9 1 0 0 9 2
15 1 0 9 4 1 0 9 1 0 9 13 12 9 9 2
11 1 10 9 4 1 10 9 13 14 12 2
24 0 9 13 13 1 9 0 9 1 9 2 9 9 2 9 2 9 9 1 9 2 9 2 2
8 9 1 10 9 13 9 3 2
7 9 9 13 0 0 9 2
12 9 1 9 13 0 13 1 0 9 9 9 2
14 16 4 9 13 13 0 9 2 13 0 13 15 0 2
16 9 1 9 3 13 15 2 15 1 0 0 9 9 13 9 2
12 1 9 0 9 3 9 0 9 0 9 13 2
10 9 0 9 1 11 11 13 0 1 9
2 11 2
23 9 0 9 1 9 0 0 9 9 1 9 0 9 11 11 4 13 1 9 12 2 9 2
13 13 1 0 1 0 9 1 0 9 1 9 11 2
12 1 0 0 9 15 13 0 9 9 11 11 2
22 13 4 3 12 9 2 1 9 11 11 9 2 9 2 0 2 7 1 0 9 9 2
16 0 0 9 13 12 9 2 0 9 13 1 10 9 9 0 2
14 3 13 3 1 9 9 13 0 9 1 9 10 9 2
19 1 0 9 13 0 9 1 12 9 9 2 1 0 9 1 12 9 9 2
20 16 13 2 13 9 0 0 9 9 0 9 2 7 3 13 2 13 9 11 2
16 0 9 11 11 13 0 0 9 11 2 15 3 13 0 9 2
28 1 0 9 1 0 9 13 1 12 9 9 1 9 2 3 1 0 9 2 11 2 0 11 2 7 1 11 2
36 1 9 9 13 7 15 2 16 9 11 13 0 0 9 0 9 2 3 2 9 11 7 9 1 11 2 9 11 1 11 7 9 11 1 11 2
17 9 13 1 0 9 9 12 9 9 2 9 9 13 12 9 9 2
27 1 0 12 9 12 13 9 3 16 12 9 9 9 2 1 0 0 9 4 15 13 13 3 12 9 9 2
28 9 9 13 1 9 9 1 9 13 1 9 12 9 14 1 12 9 9 2 0 9 1 9 3 12 9 9 2
11 9 4 13 13 1 0 12 1 12 9 2
13 9 4 1 9 0 12 9 13 13 12 9 9 2
28 9 10 9 13 0 9 1 9 1 9 2 16 9 4 15 13 1 0 9 9 1 9 12 13 3 12 9 2
17 9 15 13 7 1 0 9 2 3 2 1 0 9 2 11 0 2
11 1 9 11 15 9 13 13 9 1 9 2
39 1 0 9 13 9 1 12 9 9 1 12 9 9 2 7 15 3 9 0 9 3 1 9 0 9 2 0 0 9 0 9 2 0 9 2 0 9 2 2
43 0 9 9 13 13 3 9 1 9 0 9 2 3 13 12 7 12 9 2 2 15 13 3 13 3 0 0 0 9 0 9 2 3 11 2 1 0 9 11 2 11 2 2
30 0 0 9 0 2 9 2 11 11 13 9 0 9 2 9 0 9 7 0 9 2 3 0 7 0 9 2 9 3 2
5 9 9 1 11 13
5 11 2 11 2 2
12 9 0 9 1 0 9 1 11 1 9 13 2
31 16 13 11 9 0 0 9 11 11 2 13 1 12 2 9 12 9 2 0 9 2 15 13 1 9 3 12 9 2 9 2
31 1 9 9 2 15 13 1 0 2 0 9 2 13 11 0 0 9 1 12 9 2 0 9 2 14 12 9 2 9 2 2
13 10 9 13 0 9 1 0 9 1 3 0 9 2
12 0 9 11 15 1 9 1 11 13 1 9 2
12 0 9 11 3 13 1 9 0 9 1 11 2
11 11 3 13 0 9 9 9 7 0 9 2
5 9 0 9 11 13
2 11 2
41 0 9 1 11 12 13 3 9 9 9 1 9 1 0 9 0 9 9 0 11 7 1 9 11 2 1 15 9 13 9 1 9 2 16 0 9 0 9 13 9 2
32 9 15 13 1 9 1 9 10 0 9 0 9 7 9 7 9 0 1 9 12 2 15 9 13 2 10 9 4 0 9 13 2
9 9 0 0 9 13 1 9 13 2
12 9 13 15 2 16 0 9 13 9 3 0 2
10 3 0 9 4 1 9 12 13 9 2
5 9 3 4 13 2
6 9 0 9 13 9 9
5 11 2 11 2 2
39 9 9 2 15 13 1 0 9 9 0 9 2 11 2 1 9 2 15 3 13 12 9 1 9 9 1 11 2 3 13 9 1 0 2 9 7 1 9 2
13 0 9 15 3 13 0 9 0 2 9 11 11 2
14 13 7 9 9 2 15 4 9 13 0 2 0 9 2
24 1 12 0 9 2 15 15 10 9 13 2 13 3 9 0 0 9 2 9 9 7 10 9 2
7 11 7 13 1 0 9 2
22 1 15 13 3 9 13 9 9 15 9 2 15 13 9 2 9 1 0 9 10 9 2
13 10 9 15 3 2 13 15 9 0 9 0 9 2
12 1 9 13 15 9 1 12 9 1 9 9 2
21 16 13 7 9 9 1 9 3 7 9 13 10 9 2 0 9 3 10 9 13 2
11 0 9 9 3 9 13 1 9 9 9 2
16 16 13 1 9 0 3 2 9 1 10 9 15 3 4 13 2
9 0 9 1 0 9 13 9 9 13
5 11 2 11 2 2
16 3 2 3 7 1 10 9 13 9 13 1 0 9 1 9 2
32 1 10 9 15 13 9 11 11 2 11 2 1 9 11 11 7 11 11 1 9 2 1 15 15 13 1 0 9 0 0 9 2
13 10 9 13 1 9 9 11 7 13 3 12 9 2
13 1 0 0 9 15 3 13 1 0 9 0 9 2
17 1 12 2 9 12 9 0 9 13 7 9 1 9 0 9 13 2
28 13 13 15 1 9 9 9 11 11 2 1 15 4 15 13 9 0 1 11 13 1 0 9 1 0 0 9 2
26 9 11 1 10 9 13 2 16 1 12 9 13 0 10 9 1 0 9 13 2 1 1 10 0 9 2
21 13 13 2 16 0 9 2 10 0 9 9 9 7 10 0 9 2 4 13 3 2
24 13 15 7 2 16 0 9 4 13 3 13 1 10 0 9 7 1 9 13 0 9 0 9 2
22 9 4 1 10 9 13 3 13 2 10 9 7 1 10 9 13 11 1 0 9 13 2
5 0 9 13 11 11
7 11 2 11 2 11 2 2
35 0 9 11 11 7 0 9 9 11 1 9 1 11 11 11 13 3 1 9 9 0 9 1 0 11 0 9 1 10 0 9 1 0 9 2
12 1 0 9 1 11 12 0 3 13 0 9 2
24 9 9 1 12 0 13 1 9 0 9 1 11 2 7 15 12 2 9 13 1 12 9 9 2
40 3 4 1 11 13 2 11 11 2 11 11 7 0 9 9 2 0 11 11 2 4 9 0 9 9 1 11 13 1 0 9 9 1 9 1 12 1 12 9 2
36 9 9 12 3 3 13 1 0 9 1 11 13 0 9 1 9 11 2 9 11 2 11 2 2 16 4 13 9 0 9 1 9 12 9 9 2
19 9 15 13 13 9 3 2 16 9 13 7 13 15 1 9 0 9 9 2
18 0 9 3 1 9 13 0 9 2 9 7 1 9 13 14 9 9 2
19 3 15 11 2 11 2 13 2 16 11 11 7 11 11 4 13 1 11 2
11 12 0 13 0 7 1 0 9 1 11 2
29 9 9 3 0 11 2 11 2 9 13 9 1 12 9 2 7 15 13 13 9 0 9 2 1 15 13 0 9 2
27 0 9 9 1 11 15 3 13 9 9 1 0 9 2 15 15 13 13 11 11 3 1 0 12 9 9 2
15 12 9 3 13 9 2 16 4 13 11 11 1 0 9 2
26 9 11 13 3 1 9 0 9 9 1 11 2 7 0 9 0 9 9 1 0 9 9 13 12 9 2
23 1 0 9 9 2 15 15 9 13 2 13 1 9 1 9 0 9 2 7 1 0 9 2
14 1 10 9 4 11 11 7 11 11 3 13 1 11 2
16 11 11 13 1 10 9 9 9 1 0 9 1 11 2 11 2
5 0 15 3 13 9
7 0 0 9 13 0 9 9
4 11 11 2 11
28 9 9 0 0 9 2 11 2 2 0 3 3 2 13 2 1 1 0 0 9 15 11 13 13 0 0 9 2
12 15 13 9 9 1 9 1 9 12 2 9 2
8 9 13 0 9 15 0 9 2
42 1 9 15 3 13 2 13 15 2 16 13 1 0 9 2 1 15 15 13 0 9 2 7 3 13 2 16 9 1 0 11 13 9 7 7 10 9 4 16 9 13 2
8 1 9 13 3 1 0 9 2
18 3 13 9 0 2 1 0 9 0 9 2 16 4 15 13 10 9 2
29 13 3 13 1 9 10 9 2 15 4 15 13 2 7 13 0 2 16 4 15 1 0 9 13 1 9 7 9 2
33 9 1 0 9 9 2 3 0 2 16 9 13 4 3 13 2 4 13 3 2 16 4 13 13 16 0 9 1 0 0 0 9 2
5 11 13 0 9 2
38 9 11 13 9 2 16 4 11 11 2 0 9 11 2 15 1 9 0 9 13 1 10 9 2 7 11 11 2 9 11 11 2 13 9 1 0 9 2
12 3 13 13 9 0 9 11 9 1 0 9 2
10 9 1 9 4 3 13 1 0 9 2
16 3 4 13 0 9 11 11 2 15 1 9 3 13 0 9 2
17 11 11 13 2 16 15 13 0 9 2 15 13 1 0 12 9 2
30 9 9 11 11 2 0 9 11 2 11 11 7 13 11 2 16 4 15 13 9 7 13 10 0 9 1 9 0 9 2
7 9 0 9 3 0 13 2
29 9 4 13 13 9 9 9 1 11 11 2 9 10 9 1 9 1 0 9 1 9 0 11 7 7 10 0 9 2
11 9 1 11 3 13 1 0 9 1 11 2
22 0 9 13 13 1 10 9 0 2 16 15 3 13 2 3 4 1 9 13 0 9 2
44 15 3 3 13 2 16 13 14 9 0 2 7 0 1 9 11 2 7 1 10 9 15 13 13 2 16 9 0 9 13 3 0 2 7 13 15 1 9 0 9 1 9 0 2
14 13 0 9 2 16 1 0 9 0 9 15 3 13 2
35 13 9 2 16 9 15 4 13 13 10 9 14 1 10 9 2 16 11 13 9 2 16 4 4 3 13 1 9 7 11 4 13 9 9 2
14 1 0 9 11 15 3 1 9 9 13 0 9 9 2
25 16 9 9 13 0 2 0 7 0 9 1 0 9 2 13 0 9 1 9 0 11 1 0 9 2
32 9 9 7 0 9 13 3 0 9 2 7 3 13 0 2 15 3 4 13 1 9 9 2 15 4 13 7 15 3 13 4 2
4 11 13 0 9
4 11 2 11 2
28 11 3 13 12 1 0 9 12 9 2 15 4 1 0 9 13 16 9 1 11 0 0 9 9 2 11 2 2
14 9 13 2 16 0 4 13 1 0 0 9 11 11 2
28 0 12 0 9 11 13 3 1 11 7 13 3 1 9 2 15 13 9 0 9 2 13 15 1 9 9 9 2
24 0 9 11 11 15 13 1 9 1 0 11 1 9 0 0 9 11 11 1 0 9 11 11 2
25 1 11 7 11 13 0 9 2 16 11 13 11 2 16 13 9 11 1 10 0 9 1 9 9 2
9 9 1 9 12 9 13 3 0 2
6 13 15 2 9 0 9
11 11 11 2 9 2 13 16 9 0 9 9
44 9 1 0 11 11 1 12 2 9 0 9 1 9 13 15 10 9 13 0 9 2 13 15 2 0 2 0 2 0 9 1 0 9 9 2 0 9 0 9 7 0 9 9 2
23 3 15 13 0 9 0 9 7 9 13 10 9 1 9 0 9 1 9 7 9 1 9 2
20 9 1 9 2 0 9 7 9 13 10 9 0 1 9 3 1 0 0 9 2
10 10 9 13 2 3 2 13 9 9 2
35 9 10 9 1 9 0 9 0 9 2 15 1 10 9 9 1 9 7 9 13 11 11 2 11 2 12 2 12 2 12 2 3 13 0 2
41 3 7 13 1 9 13 15 1 15 2 3 0 9 9 1 9 12 2 9 13 9 1 9 1 0 9 7 1 15 13 0 9 0 9 7 10 0 9 1 9 2
49 16 15 3 13 1 0 9 1 0 11 11 2 3 3 15 13 9 1 12 9 1 11 2 1 12 1 0 2 9 0 9 1 0 11 2 0 11 0 11 1 11 7 11 1 0 11 1 11 2
35 15 13 3 9 1 15 2 16 4 15 9 0 9 1 9 3 3 0 9 13 1 9 1 9 2 15 4 13 13 0 7 3 0 9 2
26 3 1 0 9 0 9 13 3 3 9 2 7 7 0 9 2 15 7 13 0 9 2 15 9 13 2
24 9 13 9 11 11 2 9 11 9 1 0 11 2 15 13 2 16 12 9 9 13 9 9 2
23 3 0 9 1 11 13 10 9 7 15 2 3 13 1 9 11 11 2 3 7 1 9 2
32 1 9 1 11 2 3 15 10 9 13 0 9 2 15 1 10 9 13 0 9 2 7 3 13 9 7 0 9 1 10 9 2
36 9 2 15 0 0 7 3 0 9 0 9 13 2 13 1 15 0 2 16 15 4 13 1 9 3 3 3 0 7 3 0 16 10 0 9 2
21 3 9 9 0 9 1 0 0 9 2 0 9 2 15 15 13 0 9 2 13 2
35 3 16 9 0 9 13 3 9 0 9 9 13 1 9 9 9 9 9 1 9 15 2 15 4 1 15 13 0 9 7 13 10 0 9 2
34 15 15 13 9 0 9 2 15 13 3 10 9 3 3 13 0 9 2 3 0 9 7 13 15 1 15 3 10 0 9 9 0 9 2
41 11 2 11 7 1 10 9 1 9 0 9 13 3 3 2 16 13 2 16 4 13 9 1 9 0 2 13 9 7 13 0 0 9 1 0 9 3 0 7 0 2
32 9 2 15 15 3 13 2 13 2 3 10 0 9 13 9 9 7 0 9 2 1 15 4 13 3 15 2 15 15 3 13 2
30 9 3 0 13 3 9 2 1 15 15 0 9 13 3 2 16 15 10 9 9 3 7 0 1 10 9 13 10 9 2
20 15 13 16 0 9 0 9 2 13 9 2 15 15 13 1 9 3 11 11 2
17 16 3 15 15 13 15 2 13 0 13 10 9 3 1 10 9 2
36 3 3 13 13 9 2 7 15 3 3 0 2 7 9 0 2 7 15 1 9 0 9 9 2 1 15 0 1 10 9 13 3 3 0 9 2
42 9 1 9 10 9 13 9 2 16 4 13 13 10 9 1 9 9 9 2 7 2 0 9 0 9 2 9 9 0 0 9 2 9 0 9 7 9 0 9 7 9 2
23 3 13 16 13 2 16 1 15 0 9 2 15 13 3 1 9 2 9 13 10 0 9 2
8 9 0 9 9 11 9 9 2
13 1 9 9 11 15 13 1 12 12 3 0 9 2
8 1 9 9 13 9 11 11 2
1 9
6 9 15 13 1 0 9
12 0 9 1 9 9 2 9 13 1 9 9 9
2 11 11
11 0 12 2 9 13 0 9 3 0 9 2
22 9 9 13 3 3 0 12 9 2 9 7 9 0 9 13 9 12 9 7 12 9 2
17 13 7 9 0 9 9 12 2 1 12 5 2 1 0 12 9 2
28 9 15 13 1 9 9 12 0 9 2 1 15 12 13 2 12 13 7 9 3 12 1 9 1 0 9 13 2
21 0 9 13 0 9 2 15 3 13 9 12 9 7 1 9 13 12 9 0 9 2
27 0 9 2 15 13 1 10 9 2 13 0 9 1 0 9 0 12 5 2 15 15 13 1 3 12 9 2
11 16 13 1 0 9 2 13 15 13 3 2
11 9 11 13 1 0 9 1 9 12 9 2
20 10 9 0 9 3 3 13 2 16 9 7 9 9 13 7 9 15 13 13 2
24 9 0 9 1 0 9 3 13 0 9 9 1 9 2 10 0 0 9 3 13 9 0 9 2
9 9 10 9 3 13 3 12 9 2
30 9 9 9 0 9 1 9 0 15 3 3 1 9 1 0 9 13 1 12 1 12 2 7 16 13 3 0 12 9 2
16 13 15 2 11 0 2 0 11 2 11 0 7 11 0 9 2
11 15 13 0 0 9 3 12 9 2 9 2
20 7 3 1 9 1 15 15 13 9 11 1 9 9 1 12 5 1 12 9 2
17 9 9 11 0 2 0 9 2 13 3 1 12 5 1 12 9 2
11 9 9 13 1 0 9 3 12 9 9 2
15 1 0 9 1 12 9 12 13 2 12 13 7 12 13 2
22 12 9 2 11 11 7 11 15 13 3 2 10 9 13 1 12 2 3 2 12 5 2
18 1 0 9 15 3 13 0 9 7 12 2 9 1 15 3 13 11 2
16 10 9 13 1 0 9 9 0 11 11 7 9 0 0 9 2
6 13 12 9 0 9 2
2 0 9
4 15 4 13 2
39 11 2 1 12 2 7 12 2 9 13 9 2 1 12 2 13 12 9 12 9 2 1 12 2 13 12 9 12 9 7 1 12 2 13 12 9 12 9 2
9 3 4 13 12 9 1 12 9 2
7 0 9 13 0 2 0 9
5 11 2 11 2 2
14 1 9 9 9 11 13 3 1 11 0 9 11 11 2
30 9 2 15 13 1 9 2 15 13 2 16 4 13 1 0 9 1 9 9 10 12 9 7 10 9 1 9 9 11 2
15 0 9 2 15 15 1 9 13 1 0 9 2 7 13 2
14 1 11 7 11 3 13 9 1 0 9 0 9 2 2
19 9 11 11 13 1 0 9 12 9 2 16 13 1 11 1 0 0 9 2
14 3 13 9 2 15 13 3 1 15 9 3 0 9 2
13 1 9 11 11 15 7 9 3 13 13 1 11 2
29 9 1 9 2 12 7 12 9 2 13 3 1 15 2 16 9 13 9 2 13 10 0 9 7 3 13 1 15 2
24 13 1 9 9 7 3 13 2 0 2 15 15 13 2 13 9 2 16 15 15 1 9 13 2
14 12 9 15 13 2 16 13 2 3 15 10 9 13 2
34 16 15 3 13 2 13 15 2 16 13 9 1 9 7 3 13 9 1 9 3 0 0 9 2 1 15 9 4 15 13 4 13 9 2
20 10 9 3 13 2 9 9 11 2 1 15 15 13 11 2 11 2 3 14 2
16 13 2 16 9 9 15 13 9 0 15 0 9 7 13 9 2
36 9 2 15 13 1 0 9 9 2 9 2 11 2 15 13 2 16 9 1 11 12 2 15 9 13 2 4 13 13 9 0 9 3 1 9 2
5 0 11 2 0 11
2 11 2
18 1 12 9 1 12 9 1 9 13 1 10 9 9 9 11 11 11 2
13 9 9 11 13 1 12 9 1 12 9 2 9 2
13 3 1 12 9 3 13 3 10 9 9 9 11 2
27 1 0 9 0 9 11 11 11 13 1 9 1 9 1 9 1 0 9 11 3 1 0 9 9 0 9 2
14 1 10 9 15 4 9 9 7 9 13 1 0 9 2
18 3 13 1 12 9 7 3 3 1 12 9 13 2 13 11 2 11 2
10 0 9 13 3 14 1 0 0 9 9
2 11 2
45 9 3 12 9 9 3 13 0 9 0 9 7 0 9 2 11 2 2 15 13 9 7 9 0 9 1 3 16 12 9 7 13 15 1 0 9 1 9 0 9 11 2 1 11 2
14 13 1 0 9 2 15 13 9 3 1 9 10 9 2
17 3 13 3 10 9 2 11 13 3 3 12 9 9 12 0 9 2
20 1 12 9 1 15 4 13 1 0 9 0 9 2 0 9 1 12 0 9 2
14 1 0 9 13 1 9 12 9 12 0 9 1 9 2
19 1 15 13 9 1 9 12 9 0 9 7 1 12 9 0 0 0 9 2
23 13 3 1 12 9 0 9 2 12 9 2 12 0 9 2 12 9 7 12 0 0 9 2
14 1 9 12 13 0 9 1 9 9 1 0 9 9 2
8 1 0 9 13 12 9 9 2
21 3 15 9 0 9 11 13 3 0 0 9 1 9 12 9 9 1 9 0 9 2
9 0 9 13 9 13 1 0 9 2
24 9 1 9 13 3 12 9 1 9 12 1 9 1 0 9 7 1 9 12 9 2 9 12 2
20 1 1 15 2 16 15 13 9 9 2 13 4 15 10 9 1 9 3 13 2
14 1 9 12 15 13 9 12 9 1 9 12 0 9 2
11 9 7 13 13 0 9 1 9 7 9 2
12 13 3 1 0 9 2 15 13 1 0 9 2
13 1 9 10 9 4 13 0 12 7 12 9 9 2
18 1 9 4 13 4 13 9 9 0 9 2 15 13 13 1 12 9 2
11 9 1 10 9 4 13 13 12 9 9 2
6 9 13 13 11 11 2
10 1 9 9 15 1 9 13 10 9 2
5 9 13 0 9 2
6 9 1 9 9 9 12
5 11 2 11 2 2
25 9 9 9 3 3 13 9 9 7 9 11 11 9 9 11 11 1 11 1 9 1 11 1 11 2
37 10 12 9 0 9 13 9 1 12 9 9 2 12 9 2 13 11 2 12 9 2 12 0 9 2 12 9 13 1 0 9 2 9 13 9 2 2
13 9 15 1 0 9 13 0 2 9 2 0 9 2
10 0 9 9 3 13 3 9 9 12 2
20 9 11 13 2 16 9 1 9 9 13 1 0 9 7 0 9 2 7 11 2
13 1 15 13 0 1 9 9 13 10 0 0 9 2
19 0 9 3 13 0 13 0 9 2 1 12 9 2 1 9 12 9 9 2
15 9 2 0 0 9 11 2 7 13 9 9 1 0 9 2
8 11 2 9 1 11 1 0 9
2 11 2
23 0 9 2 7 7 11 13 0 9 13 3 0 9 10 9 1 11 1 0 9 0 9 2
10 10 9 4 13 4 1 9 3 13 2
19 7 13 0 1 0 9 13 1 9 0 9 2 1 9 1 3 0 9 2
9 13 15 3 9 9 11 11 11 2
14 13 2 16 13 0 15 1 9 13 0 9 0 9 2
16 13 13 0 9 1 9 1 0 9 9 9 0 9 1 11 2
21 1 9 0 9 0 9 1 0 9 1 11 2 11 13 3 3 9 9 11 11 2
21 1 10 9 13 1 10 0 9 1 9 2 13 4 15 7 13 15 2 3 3 2
5 7 3 15 13 2
17 16 14 13 9 10 0 9 2 13 1 0 9 9 0 9 3 2
5 9 11 2 11 11
11 9 13 9 13 2 7 13 4 0 9 13
9 11 2 11 2 11 2 11 2 2
11 0 9 13 1 9 1 0 9 1 11 2
19 16 0 0 9 13 1 9 12 9 9 2 3 15 1 9 9 13 12 2
21 13 7 9 2 3 2 0 9 7 0 9 11 2 3 15 13 3 0 0 9 2
29 13 9 1 0 9 13 2 13 3 11 9 11 11 2 11 2 2 15 3 1 10 0 9 13 0 9 1 9 2
34 1 9 4 15 1 15 13 10 9 9 13 7 13 15 7 1 10 0 9 2 7 2 9 9 2 1 15 4 15 9 13 9 13 2
26 16 4 9 13 7 3 15 12 1 9 3 13 2 7 1 12 9 9 0 9 3 13 2 13 11 2
18 1 0 9 14 13 9 9 0 2 7 10 9 15 1 15 9 13 2
34 1 0 13 9 9 1 0 11 2 3 12 9 13 13 2 1 11 15 7 3 1 12 2 9 13 13 0 9 2 16 9 13 0 2
27 7 16 4 13 12 5 9 0 2 7 13 0 2 16 4 9 13 0 2 16 9 13 9 2 13 11 2
24 1 9 0 9 11 11 11 13 9 3 3 9 10 0 9 2 16 15 13 13 7 3 13 2
12 16 0 9 13 2 7 9 9 9 2 13 2
28 0 9 1 15 13 9 2 16 0 9 1 12 2 12 9 13 1 15 0 9 2 15 13 1 15 3 3 2
14 11 13 2 16 0 9 1 0 9 4 9 9 13 2
38 9 0 9 13 1 15 13 7 13 2 7 13 9 4 13 0 2 16 4 15 13 0 9 2 15 15 1 12 9 13 0 9 2 13 11 2 11 2
12 1 9 9 13 9 13 0 9 11 11 11 2
27 16 1 9 9 4 1 0 9 13 2 1 9 9 13 2 16 9 13 1 9 3 0 9 2 3 9 2
12 13 1 0 9 2 15 13 0 1 0 9 2
34 16 4 15 1 9 13 2 15 4 13 3 1 9 2 13 4 3 0 9 7 0 9 2 15 4 16 9 2 3 0 9 2 13 2
27 1 11 13 3 0 13 1 9 9 7 0 9 2 7 15 13 2 16 13 0 13 15 9 1 9 0 2
9 1 10 9 13 1 9 0 9 2
20 13 0 2 16 4 0 9 0 9 9 13 7 15 3 13 2 13 15 11 2
3 9 11 11
1 9
2 11 11
24 0 9 11 11 2 11 2 15 13 2 16 13 2 16 0 9 9 13 9 0 9 0 9 2
14 0 0 9 13 3 0 9 9 9 0 9 0 9 2
13 13 15 3 1 10 0 9 2 7 1 9 9 2
26 3 4 9 11 13 1 2 16 4 7 3 1 15 13 0 9 7 1 9 10 0 9 13 9 3 2
9 10 9 13 2 1 15 14 2 2
26 13 3 0 13 3 2 16 1 11 2 16 15 13 10 9 1 0 9 7 9 15 3 13 1 9 2
17 16 11 13 2 16 9 9 13 14 1 12 9 2 3 13 9 2
16 13 15 3 1 12 9 2 3 1 15 2 15 13 0 9 2
12 13 9 15 13 2 16 9 13 15 1 9 2
14 1 9 15 9 1 15 13 13 3 2 16 13 0 2
15 4 15 13 2 3 3 16 3 9 9 2 13 0 9 2
12 0 13 9 2 16 4 15 0 9 3 13 2
23 16 13 11 1 9 9 9 2 13 3 3 1 9 9 1 9 9 7 13 7 0 9 2
13 9 9 15 1 9 11 13 1 12 7 12 9 2
13 1 10 9 14 13 13 0 9 9 9 2 2 2
17 13 4 0 15 13 2 16 1 12 9 13 13 9 0 16 3 2
17 13 7 3 0 2 16 4 3 3 1 9 13 1 0 0 9 2
13 13 4 15 1 9 0 9 2 1 15 3 13 2
12 3 13 0 1 9 13 9 1 11 7 11 2
13 9 15 13 2 16 4 10 9 13 0 9 3 2
6 13 15 1 12 9 2
14 1 9 4 0 0 9 0 9 13 13 3 10 9 2
6 0 9 15 13 1 9
2 11 11
20 9 7 9 1 11 13 3 1 0 0 9 9 12 1 0 9 3 0 9 2
20 13 15 0 2 0 9 2 3 9 9 1 0 9 7 3 1 0 0 11 2
16 10 9 15 1 0 9 13 2 7 0 9 0 9 3 13 2
12 0 9 7 9 9 15 3 13 0 9 11 2
15 0 0 9 13 9 11 0 1 12 1 10 0 0 9 2
9 13 14 1 0 9 9 7 9 2
19 12 9 15 15 3 13 13 1 9 2 1 9 1 11 13 12 0 9 2
16 9 9 7 9 2 15 15 1 0 9 3 13 2 13 0 2
12 0 0 9 13 2 1 9 1 11 2 3 2
18 9 9 11 12 2 13 2 16 0 9 13 0 9 7 13 9 9 2
8 11 7 13 7 0 9 9 2
18 0 9 13 13 7 0 9 0 0 9 9 11 11 13 1 0 9 2
25 1 0 9 15 9 10 9 13 1 14 3 16 9 9 2 1 0 9 0 9 3 9 3 0 2
15 9 11 13 0 7 11 3 13 1 9 1 0 9 9 2
33 0 9 2 15 13 1 9 0 9 2 13 0 9 16 9 2 7 10 9 13 14 0 9 1 11 2 7 3 13 15 0 9 2
18 3 15 7 13 1 12 9 1 10 0 9 0 9 9 2 11 2 2
21 15 0 9 3 13 7 13 0 9 1 9 9 2 4 2 14 1 11 3 13 2
17 1 10 9 9 15 13 2 16 15 9 1 12 9 3 3 13 2
24 3 13 0 9 9 0 9 1 9 11 2 15 13 0 9 1 9 0 0 0 11 1 11 2
12 9 1 9 4 0 9 1 9 1 9 13 2
21 15 15 4 7 3 13 13 2 7 13 2 1 9 11 2 16 15 0 9 13 2
10 0 13 13 9 1 3 9 0 11 2
17 13 3 0 9 9 9 11 12 2 2 10 9 4 9 9 13 2
16 0 9 9 11 11 13 1 9 0 9 14 2 11 0 9 2
15 9 9 13 7 1 9 2 1 9 2 7 1 0 9 2
29 1 9 9 13 7 9 1 9 11 11 2 11 2 1 9 7 9 1 9 2 13 11 2 16 4 13 0 9 2
41 0 9 13 3 3 10 9 9 1 9 2 3 13 9 7 9 1 0 9 2 7 9 9 9 1 0 0 9 1 11 13 2 16 9 13 0 7 1 10 9 2
17 1 0 9 0 9 1 11 4 11 13 3 3 13 1 0 9 2
5 1 9 11 2 11
4 11 11 13 11
2 11 11
19 1 0 9 2 3 4 13 9 2 4 15 13 1 12 9 0 0 9 2
38 0 1 15 13 0 9 2 0 9 3 0 9 1 0 9 2 13 9 0 9 7 0 0 9 9 11 11 0 9 2 1 15 13 13 0 0 9 2
12 9 11 13 10 9 11 1 9 9 11 2 2
14 0 9 11 2 3 16 0 9 2 13 9 1 11 2
17 1 0 9 13 0 2 0 9 1 3 0 9 16 0 2 0 2
6 3 15 13 10 9 2
8 1 11 13 0 10 0 9 2
42 1 1 15 2 16 10 9 13 1 0 9 11 2 11 7 0 0 9 0 9 2 11 7 11 2 2 13 1 10 9 13 9 1 11 3 3 7 1 3 0 9 2
17 0 9 2 1 9 0 11 2 1 3 0 9 13 2 7 13 2
18 9 0 2 0 9 15 7 3 13 1 9 0 0 2 0 9 2 2
19 11 15 13 3 1 0 9 0 9 1 9 9 0 9 1 9 0 9 2
22 3 15 3 13 9 10 9 1 9 9 10 9 1 3 0 9 1 0 9 7 11 2
9 0 9 15 9 0 9 13 11 2
5 9 13 13 15 2
21 9 1 0 9 13 3 1 0 9 2 7 3 2 0 9 9 15 9 3 13 2
15 1 9 2 1 15 11 13 1 10 9 2 3 13 2 2
20 10 9 10 9 3 13 2 16 15 11 13 0 0 9 2 15 13 1 11 2
9 10 9 13 1 15 3 3 13 2
5 13 1 10 9 2
19 1 0 9 13 0 13 2 15 1 9 0 9 4 0 13 13 1 11 2
12 1 11 13 9 1 9 13 7 10 0 9 2
7 15 13 13 1 11 0 2
27 7 10 9 4 15 13 13 1 9 2 3 4 13 9 9 2 3 1 9 12 2 3 4 9 13 9 2
13 10 9 13 13 2 13 9 10 0 9 1 9 2
13 13 2 16 11 13 9 2 15 13 1 9 0 2
9 1 11 7 10 9 3 13 15 2
16 13 13 7 9 9 2 15 1 1 0 9 13 3 0 2 2
17 15 1 9 0 9 13 1 10 9 0 9 13 16 0 1 11 2
4 15 13 13 2
8 13 2 15 4 15 13 13 2
5 9 3 7 13 2
13 7 1 9 9 13 0 9 2 13 10 9 3 2
13 15 15 3 13 1 11 2 11 2 11 7 11 2
8 1 10 9 13 3 0 9 2
6 1 9 7 13 3 2
17 15 15 3 13 7 1 9 0 9 2 11 2 11 7 11 2 2
11 15 15 13 1 9 1 0 9 7 11 2
9 10 9 13 1 10 12 9 0 2
5 10 9 13 0 2
9 13 4 7 13 3 0 7 0 2
8 1 9 0 7 1 15 0 2
11 10 9 4 13 1 9 1 9 3 13 2
6 0 9 0 9 1 11
5 11 11 2 9 11
10 9 13 3 13 0 0 9 10 9 2
26 10 9 1 10 9 15 7 9 13 1 15 2 16 4 13 1 3 0 9 2 16 0 10 9 13 2
13 1 0 0 9 13 9 1 9 9 1 0 9 2
32 0 0 9 15 13 13 1 11 0 9 2 0 0 9 0 9 2 1 15 13 13 3 16 12 9 2 1 15 15 1 9 2
19 9 9 7 9 9 15 13 1 0 9 2 16 4 15 13 0 0 9 2
13 1 15 15 1 0 9 13 2 16 15 9 13 2
8 1 0 9 9 4 9 13 2
41 14 0 9 13 9 2 7 15 13 9 2 0 9 13 2 16 15 9 1 15 13 2 0 3 2 16 15 9 13 13 9 1 9 9 7 1 15 15 9 13 2
10 1 0 9 13 1 0 9 1 11 2
16 1 9 1 9 1 11 1 10 9 3 13 2 15 15 13 2
6 9 13 3 3 0 2
24 0 0 9 1 12 9 15 3 13 7 13 0 9 2 0 11 11 2 9 7 9 0 9 2
6 9 15 13 10 9 2
13 0 9 13 11 0 1 9 9 3 1 10 9 2
14 1 9 2 15 15 13 9 2 4 9 1 9 13 2
4 15 4 13 2
24 1 9 2 3 15 13 2 3 3 13 0 9 2 1 9 0 2 1 9 0 0 9 9 2
13 1 9 13 0 0 9 2 1 15 13 1 9 2
6 1 9 13 10 9 2
4 3 15 13 2
29 13 1 9 2 15 1 15 15 3 13 2 7 1 0 15 9 9 13 2 16 13 0 0 9 9 1 10 9 2
7 3 15 15 13 1 9 2
31 7 16 4 13 10 9 2 3 4 3 9 13 13 1 9 2 0 9 13 12 9 7 13 15 9 10 12 9 2 2 2
13 0 9 1 11 4 13 1 9 1 9 1 11 2
10 3 13 9 7 15 13 3 1 9 2
8 1 9 15 13 14 0 9 2
20 11 4 15 15 15 3 13 2 13 3 7 3 2 13 3 0 7 13 9 2
23 13 4 1 12 9 1 9 0 9 2 1 15 0 9 13 0 9 7 14 15 15 13 2
12 14 7 3 15 13 2 16 13 10 0 9 2
25 13 1 15 9 2 15 15 13 1 11 2 7 1 0 9 15 13 9 7 15 13 10 0 9 2
13 9 4 15 13 2 1 15 15 13 13 2 13 2
10 13 15 7 9 12 9 1 9 11 2
26 11 9 3 15 13 2 13 15 16 0 11 11 2 9 9 11 11 2 9 2 15 0 9 13 10 2
11 11 4 13 1 10 9 2 3 13 9 2
14 10 9 15 3 13 2 13 1 10 9 3 0 9 2
19 13 4 15 2 16 15 13 0 9 1 9 0 9 7 10 9 4 13 2
7 10 9 13 13 3 9 2
12 11 13 1 9 3 3 2 7 3 13 9 2
8 13 13 9 2 13 7 12 2
12 0 9 15 13 16 9 9 2 15 4 13 2
17 13 9 2 16 3 13 2 15 10 9 13 2 13 15 11 11 2
32 0 9 15 3 13 2 13 0 2 0 7 14 13 2 16 4 15 15 13 2 13 15 13 15 1 9 2 15 3 13 3 2
18 13 4 2 15 15 13 2 14 1 9 15 13 2 16 15 15 13 2
13 3 15 13 2 16 3 15 13 7 15 15 13 2
25 13 2 16 13 1 15 10 9 2 7 16 16 15 13 9 2 7 13 15 7 9 2 13 9 2
17 11 11 2 3 15 13 2 16 15 10 9 13 1 15 1 9 2
20 13 10 9 2 15 4 3 13 7 3 16 15 13 13 2 13 15 12 9 2
14 1 15 13 2 3 15 13 7 3 13 15 15 12 2
11 3 15 13 13 3 1 9 7 13 15 2
15 15 4 15 13 9 2 1 15 4 15 15 13 10 9 2
28 7 16 13 9 9 7 15 10 9 13 2 13 2 16 4 9 3 13 14 1 9 2 16 3 13 15 13 2
5 1 10 9 13 2
20 7 16 15 9 13 2 16 13 13 9 1 0 9 2 3 15 9 13 9 2
26 13 15 13 2 3 0 13 15 3 13 2 16 15 13 13 2 7 13 9 2 16 4 15 9 13 2
40 9 2 3 1 9 15 13 1 10 9 2 13 0 0 2 13 15 2 16 13 1 12 9 3 15 13 9 9 9 2 7 16 15 13 1 15 7 1 9 2
21 13 9 2 16 3 13 3 2 16 15 13 15 13 2 13 7 13 15 1 15 2
4 3 13 9 2
11 15 13 1 9 3 1 9 2 3 13 2
21 9 13 2 3 15 13 0 9 1 15 9 2 1 9 2 1 0 9 7 9 2
13 11 11 2 1 10 9 7 0 9 11 15 13 2
27 15 10 9 13 3 2 16 15 15 13 3 3 7 3 2 16 3 0 9 13 9 10 9 9 9 3 2
5 13 10 0 9 2
21 14 13 2 3 15 15 13 3 1 9 2 16 7 1 0 9 13 10 9 13 2
17 1 9 15 3 9 13 2 16 10 9 13 11 13 7 15 13 2
9 1 15 13 9 9 1 0 9 2
9 15 7 13 0 0 9 1 9 2
18 13 15 9 1 3 0 9 2 7 15 13 7 13 15 9 9 9 2
10 3 4 3 13 9 9 1 0 9 2
5 14 1 0 3 2
6 9 1 9 11 13 2
4 0 9 13 11
17 0 9 0 9 1 0 0 9 13 12 2 9 9 9 11 11 2
21 10 0 9 13 3 13 9 2 15 0 9 13 1 9 1 0 9 1 9 9 2
37 3 1 9 4 1 0 9 9 13 3 9 11 11 2 1 9 9 2 2 11 11 2 1 11 2 7 11 11 2 1 11 7 9 0 9 2 2
15 1 0 0 9 15 13 11 11 2 11 11 7 11 11 2
27 1 9 9 0 9 13 9 11 11 0 9 1 11 7 13 3 9 10 0 9 2 3 0 11 1 11 2
16 1 9 9 9 15 13 9 2 9 2 0 9 7 0 0 2
23 1 9 1 0 9 15 1 9 13 9 0 0 9 1 11 2 15 9 13 11 11 11 2
3 2 11 2
4 0 9 13 0
14 11 13 1 10 9 3 0 2 16 4 9 13 10 9
2 11 11
19 16 13 11 11 0 9 2 7 15 15 9 3 13 2 13 11 11 11 2
26 16 7 13 9 13 9 1 0 9 1 12 9 9 2 12 2 15 13 1 11 3 0 2 4 13 2
25 11 13 9 13 9 9 9 11 2 16 4 1 9 9 1 9 9 1 9 2 12 13 0 11 2
13 13 14 2 16 0 9 13 13 0 9 1 9 2
15 13 15 14 9 11 7 10 9 2 15 13 13 9 9 2
34 0 9 11 1 11 2 1 15 11 13 0 9 7 13 15 7 0 9 2 13 14 1 9 11 1 9 9 1 9 2 12 15 0 2
42 1 9 15 13 13 3 0 9 0 9 2 0 15 13 9 11 2 2 9 1 11 13 7 9 9 1 0 9 11 2 16 14 13 13 0 9 1 11 1 0 9 2
7 15 13 13 7 0 9 2
22 14 15 14 13 3 13 9 9 1 3 0 0 9 2 15 9 2 12 1 11 13 2
23 9 9 2 15 9 13 9 1 9 2 15 9 11 13 3 2 16 13 1 9 0 9 2
14 9 2 16 0 9 13 9 9 2 13 1 0 9 2
13 9 2 12 13 1 9 7 13 15 2 13 11 2
25 11 4 13 0 2 16 13 1 0 9 7 15 13 13 9 9 2 16 4 15 13 13 1 9 2
18 13 9 10 9 9 7 16 13 11 2 13 15 12 9 1 9 11 2
25 1 0 9 15 7 13 9 2 16 13 1 9 2 15 15 11 13 2 3 1 9 9 0 9 2
24 11 14 3 13 1 9 0 9 7 9 2 12 13 9 14 1 0 2 7 7 15 0 9 2
16 13 3 0 2 16 4 10 9 13 9 11 2 13 10 9 2
2 9 11
2 0 9
2 11 11
20 9 11 16 4 15 1 12 1 10 9 13 13 1 9 3 0 9 0 9 2
20 1 0 11 7 0 11 13 3 1 0 9 1 0 9 0 0 9 2 11 2
24 13 1 9 12 7 12 2 1 9 1 0 0 3 2 0 9 2 9 2 0 1 9 12 2
57 7 2 3 3 13 9 0 9 1 0 9 11 11 2 13 15 3 1 0 0 9 2 13 0 0 9 2 12 2 2 11 11 2 12 2 2 11 11 7 11 2 12 2 2 0 10 9 2 12 2 7 0 11 2 12 2 2
33 3 1 9 2 3 3 13 9 11 2 3 13 0 9 0 9 2 7 3 0 9 0 9 13 3 13 0 7 0 9 11 11 2
21 1 9 7 0 11 1 0 0 9 2 13 2 14 0 9 1 9 12 2 13 2
30 13 10 9 0 9 16 9 2 7 7 16 9 7 9 7 11 2 7 3 0 13 1 15 14 9 11 1 0 9 2
45 15 7 13 2 16 1 15 13 10 3 0 9 7 16 4 1 10 9 13 1 9 9 2 3 4 15 0 9 11 13 1 10 0 9 1 0 9 1 9 11 11 7 10 9 2
28 9 11 13 1 0 9 2 13 0 7 13 1 9 12 2 3 1 9 2 3 7 0 9 13 9 0 9 2
44 0 9 13 3 3 0 2 0 9 11 11 2 9 9 16 4 13 0 9 1 10 0 0 0 9 2 2 10 9 11 13 3 0 11 11 2 3 1 0 9 10 0 9 2
45 0 9 9 3 13 1 11 11 11 2 7 13 3 7 0 9 0 9 2 3 11 11 1 9 9 11 7 3 0 2 3 0 11 11 1 12 1 10 10 0 9 2 9 11 2
29 7 0 9 13 3 13 7 13 1 9 9 7 9 0 9 1 11 0 0 9 2 3 1 0 9 0 11 11 2
25 0 9 9 13 1 0 0 9 3 0 2 3 0 13 14 9 3 15 0 0 9 0 0 9 2
16 3 13 7 1 9 2 15 4 10 0 9 13 13 1 9 2
4 9 9 13 9
15 9 0 9 13 9 9 9 2 13 0 2 0 2 0 2
7 11 2 11 2 11 2 2
32 9 9 13 0 9 0 9 2 15 13 0 9 0 9 9 11 2 11 2 2 16 4 13 9 0 9 0 9 1 0 9 2
30 1 0 9 9 9 9 1 9 0 2 0 2 0 2 2 15 13 0 9 0 9 2 15 13 9 0 9 11 11 2
34 1 15 2 16 4 9 13 13 0 9 2 15 15 13 13 0 0 0 0 9 2 13 1 9 9 0 2 0 2 0 2 11 11 2
8 0 9 1 9 10 9 13 2
33 13 3 1 9 0 9 1 9 9 11 11 7 9 9 11 11 2 15 1 9 13 2 16 9 9 1 9 13 3 9 0 9 2
20 9 0 9 13 9 9 0 2 0 2 0 2 1 9 9 1 0 0 9 2
10 10 9 4 9 13 1 9 9 9 2
18 1 10 9 9 4 13 9 0 9 1 9 9 13 9 0 9 11 2
13 1 10 9 4 0 9 9 13 1 9 0 9 2
10 11 2 11 10 9 3 1 11 13 2
16 1 15 13 9 2 16 0 9 0 9 13 0 16 9 11 2
17 3 1 10 9 7 13 0 2 16 15 0 0 9 13 3 9 2
7 0 0 9 15 13 9 9
5 11 2 11 2 2
12 1 0 9 9 1 12 2 9 4 3 13 2
47 1 1 15 2 16 10 9 13 0 9 7 1 9 9 7 0 9 13 3 0 9 2 3 3 4 13 0 0 9 2 13 2 0 9 4 13 4 13 1 12 9 7 0 9 12 9 2
28 9 4 3 13 1 9 12 9 1 9 0 0 9 2 7 10 9 15 13 13 7 13 15 3 9 0 9 2
15 13 15 3 1 0 0 9 9 9 7 0 9 11 11 2
34 1 15 3 13 2 16 1 9 0 9 4 0 9 2 15 13 0 0 9 13 2 13 4 1 9 10 9 1 9 12 9 3 13 2
28 9 9 7 0 9 11 11 3 13 1 15 2 16 13 9 2 15 4 15 13 13 9 9 0 7 0 9 2
16 13 15 1 9 9 2 16 4 0 9 13 7 1 10 9 2
4 0 7 0 9
1 9
2 11 11
13 0 9 7 0 9 0 9 13 3 7 0 9 2
16 1 9 13 3 3 0 9 7 9 13 9 9 9 0 9 2
12 9 13 9 2 1 0 9 13 9 1 9 2
26 9 2 3 15 9 13 13 9 2 13 9 9 1 9 7 9 2 1 15 3 3 13 2 9 13 2
21 15 15 13 2 16 9 9 13 2 0 13 0 9 0 9 7 0 9 0 9 2
7 9 13 1 0 9 9 2
7 13 15 2 15 15 13 2
46 9 13 0 9 2 13 2 16 9 9 15 3 13 16 9 7 1 9 9 7 9 13 10 0 0 9 2 16 3 13 15 9 0 2 0 1 9 2 7 0 2 0 1 10 9 2
28 13 4 1 9 0 9 1 15 2 16 9 10 9 13 7 13 10 9 0 2 16 0 9 2 7 9 10 2
14 13 4 2 16 9 9 0 9 13 1 10 9 9 2
10 13 4 2 16 13 9 1 10 9 2
3 15 13 2
29 13 15 2 16 1 0 9 1 9 0 9 13 0 13 9 1 0 9 0 9 3 2 3 13 2 1 9 0 2
27 13 1 9 7 1 10 9 13 3 9 0 2 0 2 0 2 0 2 1 15 15 0 9 13 3 3 2
19 0 9 3 9 13 1 10 9 2 15 15 15 13 7 13 2 7 13 2
28 13 2 14 3 9 2 13 3 9 7 14 9 13 13 2 16 15 1 9 1 9 4 13 3 16 0 9 2
38 9 1 0 9 13 15 2 15 4 1 0 9 13 9 16 9 13 7 13 1 15 10 9 0 9 2 15 13 1 9 13 0 9 2 16 13 9 2
5 9 0 9 13 2
13 15 3 3 13 2 16 3 1 9 13 10 9 2
9 15 0 2 13 15 15 0 9 2
11 0 15 13 9 1 0 9 7 0 9 2
8 1 10 9 4 7 3 13 2
11 10 9 13 13 2 13 15 1 15 13 2
17 15 10 0 9 7 0 9 13 16 15 2 13 15 10 0 9 2
8 3 13 0 9 10 0 9 2
5 11 15 13 9 11
2 11 2
24 11 15 3 1 9 12 13 9 9 9 0 9 2 11 2 2 15 15 13 9 9 1 11 2
12 13 15 3 9 11 1 9 1 0 0 9 2
19 11 1 9 12 13 1 0 9 9 7 9 9 9 15 1 10 9 13 2
17 13 3 1 9 1 0 9 0 9 1 9 0 9 1 0 11 2
29 0 9 15 13 13 2 16 0 9 0 9 9 11 11 1 9 1 11 13 0 9 9 1 0 9 11 1 9 2
11 1 0 9 2 11 12 2 12 2 12 2
16 9 11 1 10 9 13 2 2 2 2 0 9 11 13 13 2
61 13 15 7 3 9 13 2 16 9 0 9 9 11 1 9 11 2 15 9 1 15 13 9 0 9 1 11 9 2 12 2 3 15 10 9 13 0 9 1 0 9 1 9 9 11 0 2 0 3 0 9 2 2 3 1 10 9 13 10 9 2
34 1 9 12 13 3 3 1 11 2 16 15 3 1 9 13 13 1 3 0 9 9 11 0 2 0 9 1 9 0 1 12 9 3 2
14 3 0 9 2 7 16 3 14 15 2 11 13 13 2
4 11 11 2 11
2 13 9
2 11 2
30 1 9 15 13 0 9 9 9 2 15 15 13 9 1 11 2 11 2 11 7 11 2 1 0 9 4 13 0 9 2
10 0 9 13 1 12 2 9 10 9 2
4 11 13 0 9
16 1 11 1 0 9 0 0 1 0 11 13 0 9 2 0 9
8 0 9 11 1 0 11 11 11
53 3 13 0 9 11 11 2 12 2 9 11 2 1 12 2 9 0 0 0 0 9 11 11 2 3 1 10 9 9 12 1 0 11 13 0 0 11 11 12 2 12 2 12 2 12 2 12 2 12 1 12 9 2
21 0 9 0 9 13 9 11 11 11 2 15 15 13 2 16 0 9 2 0 9 2
35 9 1 9 0 0 11 7 0 0 13 1 12 2 9 11 11 11 2 12 2 9 11 2 12 2 12 2 12 2 12 2 12 2 12 2
28 1 9 15 3 13 7 0 0 11 2 11 2 11 2 15 13 10 0 9 11 12 2 12 2 12 2 12 2
55 1 9 3 13 9 11 1 2 0 9 15 16 1 9 2 13 15 0 9 7 15 4 9 1 0 0 2 9 2 13 2 7 3 15 13 2 16 4 13 0 9 2 13 11 3 2 16 1 11 11 13 7 11 11 2
32 13 4 15 16 9 2 1 15 4 13 2 13 1 9 2 11 13 0 3 13 2 13 15 11 2 10 0 9 13 11 11 2
21 0 9 13 2 16 15 4 13 0 9 2 3 1 0 9 1 11 13 1 11 2
17 3 4 13 0 2 16 4 3 13 12 9 2 3 13 1 9 2
4 14 13 0 2
13 13 0 1 9 2 7 1 9 2 15 4 13 2
14 3 15 13 10 9 2 13 15 15 15 1 9 11 2
13 1 12 0 9 1 11 13 3 1 0 9 15 2
23 1 0 9 4 13 2 9 15 15 13 9 9 2 15 3 13 9 2 13 15 13 11 2
14 10 9 11 1 9 13 2 16 1 11 13 0 9 2
5 7 3 9 13 2
36 3 15 15 13 15 13 16 3 11 1 0 9 2 13 3 0 0 11 2 15 15 3 13 0 0 9 1 9 2 15 1 12 9 13 13 2
41 1 9 15 1 9 0 9 2 0 0 11 11 2 13 1 12 2 9 11 11 2 12 2 2 2 7 16 3 13 12 2 12 2 12 2 12 2 12 2 12 2
18 13 2 15 15 13 13 1 11 7 11 2 16 9 9 15 3 13 2
9 13 0 2 13 13 1 3 3 2
12 9 2 15 13 2 13 1 9 0 0 11 2
17 11 3 13 0 9 2 1 0 9 15 1 15 3 13 7 9 2
20 1 9 13 9 0 9 2 15 15 13 7 1 9 12 2 12 1 0 9 2
31 7 3 13 7 0 9 2 15 15 15 11 13 13 2 16 3 13 11 9 2 13 15 11 13 9 1 9 1 9 3 2
4 11 13 9 13
5 11 2 11 2 2
32 9 0 9 11 11 11 11 11 3 13 1 9 13 10 9 1 0 9 2 16 15 1 9 1 11 13 10 9 11 2 11 2
19 0 9 15 3 1 0 9 0 9 11 2 11 13 1 9 11 2 11 2
26 16 13 9 13 1 9 9 2 15 1 0 9 13 1 0 1 0 9 2 13 4 2 13 3 11 2
20 9 9 1 9 7 11 13 3 0 9 1 9 9 7 0 0 2 0 9 2
20 9 9 13 2 16 1 0 9 9 7 9 1 9 4 15 9 13 3 13 2
6 1 10 9 7 13 2
16 0 9 7 14 3 13 1 12 2 9 2 3 13 0 9 2
18 15 3 2 13 7 9 9 0 9 2 15 9 9 13 1 9 12 2
4 0 9 0 9
8 1 11 11 11 13 3 11 11
2 11 11
24 13 9 2 0 9 10 9 2 7 1 9 1 0 9 13 9 2 15 1 0 9 13 9 2
7 13 15 0 9 11 11 2
10 1 0 0 9 11 11 15 13 9 2
13 3 16 9 13 1 11 11 2 0 9 1 11 2
7 9 11 13 0 9 9 2
11 1 0 9 15 13 1 9 0 0 9 2
73 0 0 9 2 9 1 9 9 2 15 13 9 11 1 9 2 15 1 0 9 2 0 1 11 11 2 13 13 2 16 16 0 9 0 13 3 0 9 2 10 9 0 13 1 9 11 11 11 2 2 2 2 2 13 0 9 2 3 15 11 11 1 10 9 0 9 13 2 13 7 3 13 2
9 12 9 1 0 3 11 11 13 2
13 9 0 15 13 1 9 9 2 9 3 9 9 2
20 9 9 13 1 0 9 3 2 14 3 3 13 15 3 2 16 13 13 0 2
10 11 11 13 1 15 7 14 15 13 2
15 0 9 15 13 11 11 1 9 11 2 15 3 13 13 2
12 13 13 2 15 1 15 13 9 1 10 9 2
22 13 0 2 16 1 15 15 13 2 15 13 0 9 1 9 11 2 13 9 9 11 2
12 13 15 3 0 9 1 9 2 13 9 11 2
6 13 2 13 11 11 2
10 13 15 3 2 16 3 10 9 13 2
7 13 2 13 15 9 11 2
9 3 15 15 13 13 1 9 9 2
17 0 0 9 15 13 13 9 0 0 9 7 0 9 15 13 3 2
11 7 3 15 14 13 7 13 15 9 9 2
3 11 11 2
17 13 2 16 13 0 9 10 9 2 16 1 15 13 3 10 9 2
24 13 15 15 2 16 0 9 13 1 9 0 9 2 9 7 9 2 15 3 9 13 0 13 2
25 15 13 3 2 15 3 9 13 1 9 2 7 11 13 1 15 2 15 13 2 16 4 3 13 2
23 16 15 13 2 3 0 9 13 11 11 2 13 2 16 13 3 12 1 0 9 1 9 2
22 2 2 2 12 9 1 0 9 2 13 9 0 9 0 9 0 0 9 1 9 12 2
18 1 0 9 13 9 0 9 11 11 7 9 11 11 1 12 9 11 2
33 13 15 3 3 2 3 1 0 9 0 9 13 9 0 0 9 0 3 10 9 2 0 1 0 9 2 0 1 9 9 0 9 2
44 7 13 3 16 0 2 16 15 13 9 0 1 9 9 2 0 9 2 0 7 0 9 2 15 15 13 13 0 9 2 0 9 2 15 1 9 7 9 3 9 9 9 13 2
47 15 16 0 9 0 3 13 2 16 9 1 11 11 1 11 13 0 0 9 1 0 9 2 9 0 9 0 9 1 11 2 0 2 0 2 2 11 11 2 0 16 11 11 11 1 11 2
50 15 2 7 0 9 0 2 3 13 2 16 1 15 2 16 4 0 9 1 12 9 9 9 12 13 12 0 9 2 15 1 0 13 12 0 9 2 12 0 9 9 7 12 0 0 9 0 0 9 2
3 11 11 2
25 15 2 13 15 9 11 11 2 15 13 3 1 0 1 11 2 3 4 15 3 13 2 13 9 2
17 16 13 13 0 11 2 13 4 15 1 11 2 16 4 15 13 2
10 13 3 0 9 2 13 1 15 13 2
46 1 0 9 4 15 3 13 2 16 4 15 13 9 1 11 7 1 15 15 13 7 9 1 11 2 1 9 9 15 0 3 13 2 16 13 9 0 9 2 13 15 11 11 13 3 2
27 3 15 13 7 3 2 13 9 9 11 1 10 0 9 1 11 2 13 9 1 11 11 11 10 0 9 2
19 3 13 3 2 16 13 1 11 2 7 3 1 15 13 2 15 13 0 2
13 11 3 13 13 2 16 13 1 11 2 3 0 2
52 16 13 9 11 1 11 2 13 3 2 16 0 9 13 0 9 2 15 13 12 9 1 0 9 2 7 15 13 0 2 15 15 13 1 9 13 2 7 15 13 13 3 9 2 16 4 15 3 13 2 2 2
19 2 2 2 11 11 15 13 16 0 1 12 9 1 9 0 9 11 11 2
5 13 9 11 11 2
58 7 2 16 15 15 9 13 3 16 9 2 1 0 2 3 4 15 13 2 13 1 11 3 0 9 2 2 13 15 11 11 2 1 0 9 13 0 9 11 11 2 9 2 9 2 2 2 11 1 9 2 7 7 15 13 13 11 2
37 13 15 3 7 1 11 2 3 4 13 1 9 2 7 16 4 15 1 12 9 13 3 1 9 1 11 2 13 4 15 2 3 10 9 3 13 2
15 7 15 15 10 9 3 13 2 15 15 3 13 11 11 2
13 15 15 14 15 13 2 7 7 15 15 13 11 2
18 3 13 9 0 9 0 9 1 9 3 3 11 11 11 1 9 12 2
39 10 9 2 15 13 1 9 0 9 1 0 9 7 1 9 13 3 2 9 1 11 2 13 1 9 12 1 0 9 11 2 0 9 11 1 11 7 11 2
20 1 9 12 13 1 0 0 9 1 0 9 1 0 9 1 15 7 10 9 2
15 15 2 16 13 1 11 1 0 11 2 13 3 0 9 2
22 0 15 7 3 3 13 1 9 1 11 2 3 15 11 11 13 9 9 1 0 9 2
7 1 9 12 13 0 9 2
26 1 15 2 16 13 2 13 11 11 7 0 9 0 9 2 3 2 0 9 7 11 12 2 9 2 2
45 13 15 15 2 15 11 13 1 15 2 16 4 13 0 9 7 0 9 1 0 0 11 2 12 1 0 0 0 9 2 7 15 15 13 1 9 9 0 9 2 9 10 0 9 2
14 9 15 13 11 1 0 0 11 7 13 1 11 11 2
35 2 9 0 9 2 9 2 13 1 0 9 9 2 15 3 13 9 0 9 2 7 1 9 14 13 2 7 3 15 7 16 9 13 2 2
15 13 4 0 9 7 3 15 15 13 13 13 1 9 9 2
11 3 3 15 13 2 3 13 0 0 9 2
19 7 3 4 13 1 9 2 3 1 0 2 3 4 13 9 1 0 11 2
16 3 4 15 3 13 1 10 0 9 11 11 2 15 13 9 2
41 9 9 1 9 4 15 13 7 13 4 1 11 2 3 9 13 13 1 0 11 7 15 2 3 1 15 0 9 1 0 9 2 4 15 13 9 0 0 0 9 2
8 7 3 3 10 0 9 13 2
18 3 4 13 1 9 1 0 9 7 15 15 15 13 2 15 13 13 2
6 9 2 13 4 15 2
51 7 15 13 0 2 13 15 2 16 1 10 9 13 13 2 16 3 1 15 13 10 9 2 15 13 1 9 1 9 2 7 1 0 3 14 2 16 15 13 3 9 7 15 4 15 1 9 15 3 13 2
11 14 16 4 15 13 10 0 9 2 0 2
14 7 15 13 3 0 2 16 4 15 13 7 13 15 2
26 15 13 2 9 0 9 2 3 0 2 1 9 2 3 9 13 2 15 15 9 13 2 16 13 13 2
6 13 4 15 15 0 2
21 13 3 14 0 2 16 1 15 2 15 13 2 13 0 2 16 16 4 13 9 2
8 15 15 0 13 3 0 9 2
44 1 0 9 2 3 15 15 13 3 12 9 2 9 7 3 3 0 2 15 1 9 2 15 13 13 1 0 9 11 2 13 1 0 9 2 3 1 0 11 2 3 1 11 2
14 1 0 9 1 11 11 13 13 9 1 9 1 11 2
12 0 9 3 13 1 9 0 9 1 9 12 2
14 3 13 2 16 9 13 15 0 2 15 1 9 13 2
7 13 15 14 1 9 12 2
20 0 9 13 1 12 0 2 13 15 1 12 9 2 3 13 9 1 9 9 2
24 3 15 3 13 1 9 0 9 11 11 2 15 15 13 13 15 1 9 9 7 9 0 9 2
16 16 15 11 3 13 2 16 15 13 1 11 2 13 4 15 2
10 13 3 3 2 13 4 15 9 0 2
23 3 4 13 14 1 10 9 2 7 16 4 13 3 1 11 2 13 4 15 1 15 13 2
15 3 4 3 13 0 9 1 11 2 7 3 15 15 13 2
10 14 1 9 12 1 9 1 0 9 2
16 7 3 3 3 13 0 0 11 7 13 2 16 13 1 9 2
31 3 4 13 1 11 7 13 15 2 3 13 13 2 7 15 13 2 13 3 9 2 15 13 15 2 15 15 1 15 13 2
15 14 7 3 4 15 13 2 7 15 3 13 3 0 9 2
11 1 9 9 15 9 11 13 13 0 9 2
30 3 13 1 0 9 0 0 9 11 11 2 3 1 0 9 2 3 13 1 0 9 10 0 9 11 1 0 0 9 2
8 1 0 9 15 1 9 13 2
27 13 15 1 15 9 2 13 1 10 9 3 1 12 9 1 0 11 2 1 3 16 0 9 15 13 13 2
10 10 9 3 11 7 9 13 0 9 2
24 0 9 10 9 3 11 11 13 1 9 7 1 9 9 1 0 9 2 11 1 0 11 2 2
22 9 13 9 2 15 15 3 13 2 13 3 9 9 9 2 15 0 9 13 10 9 2
10 15 7 10 9 1 9 13 3 3 2
10 13 2 16 13 0 9 1 0 9 2
22 9 15 3 13 0 2 7 15 13 0 9 2 16 3 0 13 7 0 13 0 9 2
15 7 0 9 3 13 13 9 9 9 9 7 9 0 9 2
4 15 13 9 2
21 1 0 9 2 1 15 2 16 4 13 1 9 2 4 15 13 9 2 14 9 2
40 11 11 1 9 9 11 2 15 3 13 1 10 9 1 11 7 13 9 15 1 9 11 13 3 2 9 2 16 15 13 1 0 2 7 0 9 2 7 13 2
30 16 15 10 9 13 13 2 9 13 13 14 1 9 2 16 15 0 7 0 13 1 9 7 15 0 7 0 1 9 2
24 7 3 10 9 2 15 3 1 9 10 9 1 9 13 2 3 1 9 13 3 10 0 9 2
26 9 1 9 9 7 0 9 13 2 13 15 2 1 11 11 3 0 7 13 1 15 13 0 7 0 2
49 1 9 12 13 1 9 11 11 10 9 1 9 9 11 11 2 1 12 9 3 13 11 2 1 0 9 12 13 3 3 10 0 0 9 2 16 9 9 1 0 9 13 13 1 9 3 0 2 2
20 16 4 11 13 9 2 4 13 9 1 11 2 16 10 9 4 13 1 0 2
13 11 3 13 13 9 9 11 2 7 3 9 11 2
10 10 9 13 3 11 11 1 9 11 2
12 13 15 7 1 0 2 3 0 9 0 9 2
9 3 13 9 0 7 11 1 15 2
5 7 13 7 0 2
68 11 11 2 15 9 9 3 13 1 0 9 2 7 1 0 9 1 11 2 12 2 12 2 13 3 2 16 3 11 2 11 3 13 7 13 15 15 2 10 9 1 11 3 13 2 2 2 2 1 9 1 15 13 2 9 11 2 3 0 1 15 2 15 13 1 11 13 2
21 13 15 3 2 16 15 3 4 1 10 9 13 2 15 3 4 1 10 9 13 2
28 0 9 7 0 9 11 13 1 11 11 3 16 15 0 9 1 9 9 3 2 16 4 3 13 0 9 9 2
15 13 3 2 16 0 9 13 3 1 0 9 10 0 9 2
23 9 13 9 9 2 1 15 4 13 13 11 1 11 7 13 4 3 13 7 0 9 9 2
40 13 7 3 9 7 16 13 1 0 9 9 0 0 9 1 9 0 9 2 0 1 0 9 2 3 9 9 9 0 9 11 11 2 2 13 1 15 3 0 2
23 15 15 3 2 1 15 2 16 4 13 1 11 2 13 3 2 16 4 15 13 1 9 2
11 13 15 15 12 9 1 9 1 12 9 2
23 1 0 7 0 13 0 9 2 15 10 0 9 13 1 15 2 16 4 13 1 9 13 2
21 13 13 1 10 9 9 2 7 13 2 16 15 4 13 1 9 9 0 9 3 2
26 1 0 13 0 9 2 15 4 15 13 13 9 0 9 2 1 15 0 9 2 7 13 3 3 9 2
6 13 15 7 13 3 2
24 1 0 9 13 9 2 15 3 13 1 0 2 7 3 4 13 9 0 9 13 2 13 9 2
12 1 0 3 13 9 2 15 13 16 9 13 2
9 15 13 3 11 2 11 2 11 2
13 3 2 16 1 0 9 2 14 15 1 15 13 2
43 3 11 2 1 12 9 9 2 15 13 9 1 0 9 2 0 9 1 15 7 3 14 13 7 10 9 13 0 2 3 13 1 10 0 9 2 3 16 4 15 13 9 2
32 1 10 0 0 9 13 9 11 9 9 9 9 9 12 2 15 13 0 0 9 1 11 1 9 3 0 9 11 1 0 9 2
24 13 15 3 0 2 13 9 2 16 4 0 9 13 13 1 0 9 2 1 9 15 0 9 2
30 13 4 9 2 16 15 13 0 16 13 9 1 9 9 1 0 9 2 7 13 2 16 15 13 3 14 15 3 0 2
36 1 0 9 13 1 0 9 2 9 1 0 9 2 0 9 15 13 2 7 15 13 9 3 0 9 1 9 2 3 15 3 3 3 15 13 2
7 13 15 0 2 7 0 2
12 9 1 0 9 13 1 11 11 3 0 9 2
29 3 3 13 0 9 13 0 9 2 13 2 16 13 13 1 0 0 9 2 16 0 9 4 13 13 3 0 9 2
11 13 4 3 2 16 9 4 13 13 3 2
43 16 9 13 1 9 2 13 7 15 9 7 1 15 2 15 4 13 1 9 2 15 13 9 7 1 15 9 13 2 13 0 9 0 7 9 13 13 3 9 7 9 0 2
10 13 4 15 2 16 4 13 3 9 2
33 10 9 3 3 13 2 16 0 9 1 0 9 9 1 0 9 15 1 15 13 0 9 2 1 15 15 13 10 0 9 0 9 2
43 3 13 0 9 0 9 11 2 1 15 4 0 9 13 9 3 9 0 9 2 7 3 10 0 7 0 9 2 13 3 13 1 9 9 0 9 10 9 13 3 7 3 2
18 13 9 1 10 9 2 16 4 13 2 10 13 9 2 13 1 15 2
10 13 1 9 0 9 7 13 13 3 2
39 11 11 1 9 1 3 0 0 9 1 0 0 9 0 0 11 1 12 2 9 12 3 13 2 16 11 11 15 13 16 0 7 0 9 0 3 0 9 2
16 13 0 9 9 9 11 7 0 9 9 1 0 9 11 11 2
9 13 13 3 0 2 7 15 13 2
38 13 15 9 2 15 15 13 2 15 13 13 2 15 13 13 0 7 3 3 3 13 1 0 9 2 15 13 0 1 9 7 10 9 2 13 11 11 2
12 2 2 2 13 9 3 2 13 15 1 0 2
36 9 0 9 1 11 11 11 2 9 11 15 13 16 9 1 10 0 9 1 9 1 0 9 0 7 0 11 2 3 13 1 9 7 13 15 2
25 0 9 15 13 1 10 9 9 2 3 0 2 1 9 9 2 1 9 0 9 2 1 9 9 2
19 3 13 0 9 11 7 0 9 1 0 9 2 3 11 2 11 2 11 2
11 1 12 9 15 13 1 9 9 11 11 2
12 15 4 15 13 9 2 11 2 13 15 3 2
26 0 9 15 3 3 13 1 3 3 0 9 9 2 15 13 3 16 0 9 2 7 15 15 3 13 2
10 11 11 15 3 2 14 9 2 13 2
7 13 9 7 13 4 3 2
15 9 15 15 3 13 2 15 13 9 1 0 7 0 9 2
28 13 4 15 2 16 9 13 2 16 9 13 13 1 10 9 2 16 9 13 2 16 15 13 9 13 1 9 2
17 13 2 16 9 13 9 2 15 9 13 13 15 2 15 13 15 2
6 14 0 13 15 15 2
9 0 2 0 7 9 9 9 13 2
17 9 13 10 0 9 2 15 13 13 15 2 15 15 15 13 13 2
5 9 11 11 2 11
3 0 9 13
7 1 12 9 2 9 1 11
17 0 9 13 14 12 0 9 0 1 11 1 12 9 1 12 9 2
21 1 9 3 13 15 1 0 9 1 9 11 7 13 16 9 1 0 3 0 9 2
21 9 14 13 9 2 1 15 7 13 15 0 9 2 1 15 13 9 3 0 9 2
22 16 7 11 13 2 16 13 0 9 2 13 9 1 11 9 2 16 4 13 10 9 2
10 16 4 13 9 2 13 11 1 0 2
20 3 1 11 13 15 12 9 7 0 9 13 11 7 13 15 1 9 1 11 2
8 4 13 12 9 7 12 9 2
13 9 7 10 9 13 1 9 7 9 1 0 9 2
17 1 9 3 1 0 0 9 13 4 11 1 9 1 0 2 11 2
20 2 0 9 12 2 12 2 9 2 12 2 9 2 12 2 9 12 2 9 2
6 1 12 9 2 11 13
18 1 10 9 13 0 9 0 9 2 16 4 0 0 9 13 1 9 2
15 9 12 2 9 13 2 16 3 0 0 9 4 13 9 2
20 15 15 13 1 0 9 9 2 15 13 9 12 2 9 1 9 11 7 11 2
24 1 9 2 0 1 9 2 13 3 9 1 9 2 13 0 9 2 16 15 13 9 0 9 2
21 0 7 0 1 9 13 10 9 1 15 14 15 2 15 13 13 1 9 7 9 2
21 9 2 15 1 0 9 4 4 13 3 13 0 7 0 9 2 13 3 1 9 2
23 1 9 10 9 15 13 9 7 0 9 1 15 2 15 13 7 15 4 13 11 7 11 2
42 0 9 11 2 15 13 15 0 1 9 0 0 9 2 13 13 9 1 0 9 2 15 13 1 0 9 10 0 9 1 11 7 1 11 2 15 11 13 1 10 9 2
6 11 13 14 12 9 2
31 13 15 0 9 1 10 9 2 15 13 0 9 1 11 2 11 7 11 7 15 13 1 9 7 9 0 2 0 0 9 2
20 2 0 9 12 2 12 2 9 2 12 2 9 2 12 2 9 12 2 9 2
7 1 12 9 2 9 0 9
17 13 1 9 9 2 15 13 1 0 9 1 0 9 12 2 9 2
15 13 4 15 1 9 0 15 9 0 9 7 0 9 9 2
22 16 15 0 9 4 13 2 16 13 0 10 0 9 13 1 3 0 9 9 2 2 2
30 13 15 2 16 1 9 2 3 13 7 9 9 9 0 9 9 9 2 13 9 3 13 10 0 9 7 9 1 9 2
10 3 7 13 1 0 9 10 9 13 2
49 10 0 9 13 7 0 2 0 7 0 9 9 7 9 0 9 2 0 1 0 9 1 9 2 3 3 3 0 2 9 10 9 2 15 0 9 3 13 10 0 9 0 9 9 2 12 9 11 2
7 7 15 1 10 9 13 2
15 10 9 15 13 1 0 7 0 9 2 15 1 15 13 2
5 2 13 12 9 2
14 2 0 0 9 2 9 12 2 9 12 2 9 12 2
6 13 11 11 7 11 11
28 0 9 2 9 7 9 9 11 3 2 9 3 2 11 11 15 13 9 12 1 3 0 0 9 16 11 11 2
18 13 1 9 11 2 3 13 0 9 2 9 13 0 9 1 9 2 2
21 1 9 12 2 12 13 9 7 9 1 0 9 2 1 9 12 13 1 0 9 2
24 1 9 0 0 2 0 9 15 13 3 1 0 2 0 2 0 9 1 0 9 2 12 2 2
9 13 3 0 9 0 9 10 9 2
8 13 0 9 1 9 1 11 2
9 1 9 13 0 9 1 9 12 2
75 0 9 0 9 2 12 2 2 3 3 3 2 12 2 2 10 11 2 12 2 2 13 15 9 2 13 15 9 2 12 2 2 1 9 0 2 12 2 2 0 9 2 12 2 3 0 9 12 2 2 13 9 2 12 2 7 0 9 2 12 2 4 13 1 12 9 7 13 1 0 9 12 9 9 2
27 9 13 9 10 0 0 9 2 1 15 3 13 0 9 0 9 2 0 15 1 0 0 9 1 9 12 2
5 9 11 11 2 11
3 9 1 11
5 11 2 11 2 2
18 0 9 13 3 1 9 1 0 11 0 9 11 2 0 0 0 9 2
32 9 13 11 11 9 11 7 9 9 2 11 11 11 2 15 3 3 1 9 13 9 7 1 0 9 13 1 0 9 0 9 2
32 11 11 1 9 1 10 9 11 2 11 15 13 0 9 1 9 7 15 3 14 3 13 1 10 0 9 1 11 11 0 11 2
23 0 9 2 11 11 2 11 11 2 11 2 11 2 11 2 11 11 2 11 11 2 11 2
15 0 11 11 9 11 2 11 13 0 0 9 12 2 12 2
6 0 0 9 13 1 11
8 11 11 2 9 0 9 9 0
1 9
25 15 0 3 13 2 16 0 9 15 13 1 9 15 3 2 15 3 0 9 15 13 1 10 9 2
22 0 9 13 3 9 13 15 1 9 1 10 0 9 7 13 10 0 9 1 0 9 2
23 9 0 0 9 1 9 1 3 0 0 9 13 3 16 0 9 0 0 9 1 0 9 2
14 13 3 1 9 0 9 0 9 0 0 9 1 9 2
49 9 2 1 15 15 0 9 13 9 0 0 9 1 9 2 13 9 0 9 2 15 1 9 0 9 13 2 16 0 9 13 9 2 7 9 2 0 0 0 9 2 13 9 9 2 3 15 13 2
16 11 11 11 13 10 0 9 9 2 9 7 9 1 9 12 2
26 0 0 9 13 0 9 0 0 9 2 1 15 9 3 13 10 9 7 15 13 13 2 3 13 9 2
25 0 9 7 3 0 9 13 2 16 0 9 9 7 9 13 13 1 10 0 9 1 3 0 9 2
27 7 2 13 11 2 4 13 9 13 1 9 7 0 9 13 9 2 15 4 13 0 9 1 10 0 9 2
11 11 15 3 13 1 0 0 9 0 9 2
15 3 0 0 9 13 1 15 3 3 0 16 1 0 9 2
15 0 9 13 4 1 11 13 3 3 2 7 1 0 9 2
26 1 9 2 3 15 9 13 1 0 9 2 13 4 9 13 1 10 9 7 13 15 0 9 0 9 2
18 1 9 0 9 4 9 13 13 1 0 9 7 13 1 0 0 9 2
11 9 13 4 13 2 3 13 1 0 9 2
17 7 9 13 3 16 9 14 9 7 0 9 13 14 1 9 9 2
13 1 9 1 0 9 15 13 13 1 0 9 3 2
7 9 1 15 13 3 13 2
33 0 9 9 0 9 7 9 9 15 3 1 0 0 9 7 0 9 9 13 1 0 9 12 2 9 2 0 9 7 9 0 9 2
8 9 14 13 2 7 3 13 2
12 1 0 9 15 1 9 13 3 9 0 9 2
19 3 1 0 11 2 1 9 0 9 2 13 9 0 9 7 0 0 9 2
13 1 0 9 3 13 0 9 2 3 0 0 9 2
28 3 15 13 14 0 9 2 15 13 9 9 13 9 2 15 1 0 9 0 9 13 9 12 5 9 0 9 2
12 0 9 0 0 9 13 9 1 0 0 9 2
18 0 7 0 9 1 0 9 13 7 3 13 16 9 10 9 1 9 2
16 9 13 7 0 2 16 16 4 15 13 13 1 12 0 9 2
34 13 2 14 3 12 0 9 13 0 2 14 15 3 13 9 0 9 2 7 3 9 9 14 0 9 1 9 9 7 0 9 0 9 2
4 11 3 9 9
1 9
2 11 2
11 11 11 11 4 12 9 13 0 9 9 2
23 9 11 11 13 1 0 9 1 0 9 3 2 1 11 2 11 2 7 11 2 11 2 2
31 11 13 12 9 7 13 15 1 0 12 9 1 12 2 9 2 11 2 12 11 2 13 12 7 11 2 11 2 12 9 2
5 0 9 13 0 9
10 0 9 13 2 16 3 13 0 9 2
16 1 10 9 15 13 9 9 9 2 15 1 9 13 1 0 2
8 7 12 1 15 13 7 11 2
14 9 11 3 13 1 9 1 9 1 9 1 9 12 2
27 1 9 1 9 10 0 9 13 12 9 2 1 9 12 9 2 12 9 2 12 9 7 9 12 2 12 2
26 0 9 1 9 13 1 9 12 2 7 15 1 11 1 9 3 12 2 12 2 16 11 11 13 9 2
29 1 9 1 9 12 3 13 1 11 7 1 12 9 3 13 0 7 3 0 9 2 11 13 0 9 9 1 11 2
9 3 0 13 11 1 9 1 9 2
22 15 15 13 1 12 9 3 1 9 2 12 2 12 2 12 2 12 2 12 2 12 2
20 0 9 13 1 9 12 1 11 2 1 12 9 3 11 3 12 2 12 13 2
9 1 0 9 13 1 11 7 11 2
7 11 3 13 3 0 9 2
21 3 1 10 9 13 1 9 1 9 13 2 3 13 1 9 1 0 9 1 9 2
21 13 1 10 9 7 10 0 9 1 10 12 0 9 2 16 13 11 12 2 12 2
13 7 9 1 11 2 12 2 12 2 13 10 9 2
12 7 9 0 9 13 9 12 2 12 1 11 2
20 1 0 9 13 0 9 12 0 11 11 11 2 15 3 1 12 13 9 11 2
15 1 9 3 13 14 12 9 1 0 0 9 11 0 11 2
14 0 9 13 0 0 9 11 1 11 7 11 11 11 2
3 2 11 2
9 15 13 1 9 2 13 9 1 9
5 11 2 11 2 2
27 9 2 7 9 2 13 15 9 2 7 7 11 2 15 1 0 9 13 3 3 0 9 0 9 0 9 2
21 9 9 11 11 7 11 11 13 1 15 7 9 2 7 9 1 9 1 12 9 2
7 13 4 14 9 2 13 2
9 1 9 9 15 13 14 9 9 2
19 3 10 11 13 1 15 3 3 2 16 4 15 13 9 7 13 0 9 2
16 14 9 1 9 13 12 0 9 1 0 9 12 12 1 9 2
19 3 12 12 13 1 9 9 7 13 2 16 15 15 9 1 12 9 13 2
27 3 16 4 13 3 13 1 3 0 7 0 9 2 15 13 0 9 2 3 13 3 13 3 12 12 9 2
36 14 2 0 9 2 15 15 1 15 13 2 13 1 15 2 16 15 9 9 0 9 7 0 9 9 1 0 9 13 13 2 13 11 2 11 2
18 1 10 9 4 15 13 13 3 1 0 9 11 12 7 13 0 9 2
17 9 0 9 13 9 2 15 13 9 1 0 9 2 12 9 3 2
16 1 15 13 14 7 0 9 2 13 1 0 9 11 2 11 2
24 0 9 13 9 1 9 7 1 9 9 7 13 15 1 9 2 15 3 13 9 1 0 9 2
4 9 9 0 9
6 11 11 2 9 0 9
22 1 0 9 15 1 0 9 13 13 9 1 9 0 9 1 9 0 9 1 0 9 2
27 9 1 0 9 1 3 0 9 15 13 0 9 9 7 0 9 2 15 15 13 13 1 9 0 11 11 2
11 1 9 13 1 0 1 10 9 13 3 2
51 1 1 9 7 9 0 9 0 9 2 1 9 13 0 0 9 9 7 1 9 1 15 2 16 9 4 13 1 9 0 0 9 2 13 9 0 9 1 9 13 1 9 9 2 15 13 0 9 9 9 2
17 13 3 9 13 9 9 1 9 0 9 1 0 9 9 0 9 2
43 0 9 13 13 9 2 9 2 9 7 9 9 9 1 9 1 0 9 1 0 9 7 1 9 1 3 0 9 9 1 0 9 2 0 0 9 9 7 9 1 10 9 2
18 10 9 13 13 3 2 7 9 9 1 9 0 9 7 9 0 9 2
15 1 0 0 9 9 13 7 13 0 9 9 0 9 9 2
44 1 9 0 9 13 3 9 0 9 9 7 3 3 13 0 9 9 3 2 16 4 4 1 9 1 0 9 7 1 9 0 1 9 13 1 0 9 7 1 3 0 0 9 2
25 9 13 7 9 10 9 1 0 9 3 13 9 0 9 7 3 7 9 7 0 9 0 9 9 2
27 9 3 13 0 0 9 7 13 9 0 9 9 2 13 9 7 9 9 7 0 2 0 7 0 9 9 2
32 0 9 0 9 9 2 0 16 0 9 2 9 1 9 2 0 9 3 2 2 13 0 1 9 1 9 0 9 3 3 13 2
26 9 2 0 9 10 1 9 3 0 9 2 7 0 1 9 7 9 1 9 1 9 13 1 15 0 2
19 3 2 9 1 0 9 4 13 13 0 9 2 16 4 13 16 0 9 2
18 9 13 3 1 9 9 1 9 7 2 15 7 9 7 9 0 9 2
24 3 3 4 1 0 9 13 9 0 0 9 1 9 15 2 16 13 3 9 1 15 7 15 2
33 9 0 9 3 13 7 13 13 9 9 9 2 16 9 15 9 13 2 3 15 13 2 1 9 10 9 2 1 0 9 1 9 2
1 9
7 9 11 2 11 1 9 12
3 9 0 9
2 9 11
4 9 9 4 13
6 0 11 13 1 0 9
2 11 11
12 9 11 13 1 0 11 7 1 9 1 0 2
19 13 0 9 1 11 7 0 1 9 2 7 9 1 0 9 10 9 13 2
20 3 13 9 10 9 2 1 15 4 13 1 0 9 11 11 9 2 11 11 2
23 12 1 9 13 0 7 1 10 9 3 0 9 1 3 2 1 9 12 2 3 0 9 2
13 0 9 15 13 3 7 13 7 0 9 1 9 2
16 15 15 13 7 3 0 9 9 9 2 7 7 9 0 9 2
14 1 9 12 4 13 1 9 12 9 7 11 3 12 2
16 1 15 4 4 0 9 13 1 9 1 0 0 7 0 9 2
8 2 15 7 13 13 0 9 2
15 11 13 3 0 9 9 16 15 7 10 9 13 1 0 2
11 0 9 13 3 0 9 16 15 1 9 2
12 3 15 13 13 9 7 9 2 3 3 9 2
11 11 13 1 9 0 10 9 1 0 9 2
4 9 2 9 2
14 7 15 3 0 9 2 15 3 13 10 9 2 13 2
27 1 15 3 3 13 9 7 3 0 9 2 16 10 1 15 0 9 13 3 1 9 16 3 3 0 11 2
6 0 13 7 9 9 2
20 9 13 3 9 15 1 9 13 2 16 15 13 1 9 1 9 7 1 9 2
14 9 10 9 13 13 11 11 2 0 1 9 9 12 2
39 16 15 13 1 0 0 9 1 0 0 7 0 9 2 15 3 9 13 2 16 4 15 13 1 9 9 2 1 15 13 0 7 9 13 0 10 10 9 2
23 9 13 0 9 2 7 3 1 11 2 3 15 9 13 1 0 9 2 15 13 3 9 2
7 2 9 9 15 13 13 2
8 13 0 9 2 3 13 9 2
9 13 0 0 9 2 13 0 9 2
25 1 9 0 9 13 9 1 12 2 1 0 9 0 9 3 1 12 1 12 0 9 7 12 9 2
18 13 0 9 11 2 1 15 13 1 9 9 1 9 3 1 12 9 2
18 1 0 9 13 9 1 9 9 11 11 2 15 13 3 0 1 11 2
8 3 15 3 13 12 12 9 2
10 3 13 7 9 2 15 4 3 13 2
10 1 9 0 9 13 10 9 9 9 9
5 9 11 11 2 11
10 11 2 11 2 3 1 9 7 1 11
3 1 0 9
5 11 2 11 2 2
30 0 9 2 11 2 13 13 2 16 9 0 9 1 0 0 9 4 13 1 9 0 9 2 3 15 3 7 9 13 2
20 13 1 15 2 16 1 10 9 15 13 13 0 9 2 7 15 9 7 9 2
23 11 2 11 2 13 0 9 2 3 7 1 11 2 3 13 1 0 9 1 9 0 9 2
19 1 0 9 4 13 3 2 0 9 1 11 13 3 0 0 9 11 11 2
5 11 11 13 9 11
2 11 2
37 9 11 7 15 13 2 16 15 13 0 2 0 9 13 0 9 9 2 13 0 9 11 11 2 15 3 13 1 11 1 9 11 1 9 7 9 2
15 13 9 2 16 9 9 13 9 2 3 3 13 9 9 2
12 13 3 1 9 9 1 11 7 10 0 9 2
16 15 13 2 16 9 9 13 1 9 1 10 0 7 0 9 2
11 11 13 1 9 1 11 9 1 0 9 2
8 3 13 10 9 9 3 13 2
5 1 11 11 3 13
2 11 2
12 11 3 13 9 13 0 9 1 0 0 9 2
11 13 15 3 1 0 11 9 11 11 11 2
16 15 13 1 9 1 9 10 9 2 7 1 0 9 15 13 2
16 11 13 2 16 15 15 13 13 9 7 1 9 0 9 9 2
6 0 11 3 14 1 11
8 11 11 2 9 0 9 1 11
15 9 0 9 0 1 11 13 3 0 9 9 9 0 9 2
27 13 15 9 2 16 1 0 9 15 13 3 2 16 15 13 1 0 9 2 7 13 1 9 0 0 9 2
25 9 13 3 1 9 9 9 11 7 0 11 1 11 1 11 2 7 1 0 9 1 0 9 9 2
20 0 9 9 11 13 3 1 12 9 13 1 9 1 9 7 9 0 9 11 2
20 1 0 9 13 13 2 16 15 2 15 15 13 2 13 0 2 3 0 9 2
37 0 9 3 13 10 0 9 1 11 2 3 13 1 11 0 0 9 7 9 2 7 13 3 3 2 16 13 0 0 9 7 9 1 9 0 11 2
58 15 13 1 0 9 3 0 3 1 9 1 0 9 2 15 4 3 13 7 1 1 15 15 0 9 13 0 9 2 15 15 2 0 9 2 3 13 13 2 16 15 0 9 2 1 0 9 10 9 2 13 0 9 13 1 10 9 2
8 3 13 9 2 0 10 9 2
8 1 0 9 9 1 9 14 13
21 9 9 1 0 9 13 0 9 9 1 9 9 11 1 11 1 9 9 1 11 2
12 11 15 13 11 11 2 9 9 9 0 9 2
7 1 10 9 13 0 9 2
17 13 9 1 11 2 0 11 7 11 2 13 15 3 0 0 9 2
22 1 11 4 9 9 13 9 13 1 9 9 7 9 4 13 9 9 13 3 10 9 2
36 1 9 11 1 11 2 3 1 0 13 11 11 11 7 3 3 13 9 10 9 2 13 3 1 9 7 0 9 3 9 1 0 9 9 9 2
16 15 13 9 9 13 1 9 9 12 7 9 13 1 9 12 2
11 1 10 9 13 0 13 1 9 0 9 2
13 13 0 2 16 4 3 13 2 4 15 3 13 2
17 7 1 9 3 13 13 0 9 7 9 13 9 2 13 11 11 2
14 9 1 0 9 13 3 1 11 3 1 9 0 9 2
12 4 3 3 13 9 12 9 2 0 7 0 2
21 1 9 1 9 9 7 10 9 1 0 9 15 13 9 13 1 0 9 12 9 2
15 13 4 1 15 1 9 9 13 2 7 13 15 0 9 2
24 13 15 1 11 13 1 0 9 7 3 15 9 13 2 13 11 11 11 2 9 9 0 9 2
3 2 11 2
6 1 0 9 3 1 9
25 1 11 7 1 11 13 9 3 0 9 1 9 2 7 1 3 2 0 2 9 2 9 14 13 9
2 11 11
17 0 0 9 13 1 15 12 9 1 9 0 0 9 11 2 11 2
11 9 2 12 9 2 12 9 2 10 9 2
24 1 9 0 9 13 1 15 7 0 9 9 0 11 2 15 15 13 1 9 1 9 1 11 2
65 1 0 9 2 15 9 11 13 1 12 0 9 1 11 2 12 2 12 7 12 2 12 2 2 1 0 11 2 1 11 1 11 12 2 12 2 7 1 0 11 2 1 11 12 2 12 2 1 11 12 2 12 7 1 11 12 2 12 2 13 9 9 3 3 2
26 9 1 3 3 0 9 2 15 15 4 13 13 1 10 0 9 2 0 10 0 9 7 11 3 13 2
25 15 0 1 10 0 9 3 14 13 2 3 13 9 9 1 11 2 3 1 0 9 13 12 9 2
30 3 9 1 12 11 13 3 0 1 12 9 15 3 2 16 9 11 1 9 13 2 16 1 9 10 9 13 3 0 2
27 13 4 15 13 1 9 1 9 2 15 1 15 13 3 7 1 9 12 1 12 3 16 15 2 13 11 2
18 9 2 15 9 13 2 4 15 13 13 13 9 2 15 15 3 13 2
8 1 0 3 4 13 10 9 2
24 11 3 13 1 0 2 16 9 0 9 1 11 2 15 13 1 9 1 9 2 13 0 9 2
17 9 1 0 7 0 9 15 3 13 7 13 9 13 1 15 9 2
33 16 9 3 15 0 0 9 13 2 3 15 13 13 1 9 2 15 15 4 3 1 0 9 1 11 7 1 0 9 1 11 13 2
18 9 13 3 1 9 0 1 0 9 7 1 9 4 15 13 13 3 2
32 9 1 9 1 11 7 9 1 0 9 0 0 9 1 0 0 9 2 0 9 7 0 9 13 7 1 9 13 7 0 9 2
26 9 0 9 0 9 11 11 7 9 3 3 13 1 14 12 9 0 11 2 3 13 1 9 0 9 2
11 13 9 7 9 16 0 9 9 15 13 2
19 16 13 3 12 1 9 0 9 2 13 13 9 13 7 9 1 10 9 2
11 9 7 3 13 10 0 0 9 1 9 2
23 16 15 13 11 11 2 13 15 3 1 0 9 1 9 9 9 2 16 10 9 13 15 2
21 1 9 12 1 9 15 14 11 11 13 7 13 2 15 13 0 2 9 13 0 2
15 0 9 0 9 13 12 9 1 0 9 7 12 1 0 2
46 3 12 1 15 4 3 13 13 1 15 2 16 4 0 9 13 7 1 0 9 0 9 16 0 9 1 9 7 16 4 15 9 2 16 3 9 13 13 2 13 1 0 9 3 13 2
6 1 11 15 3 13 2
18 1 3 2 0 2 9 2 9 7 14 13 1 12 9 9 2 2 2
31 7 11 2 15 3 13 0 9 9 0 11 2 12 1 0 0 9 2 13 2 16 15 9 13 2 1 0 9 3 0 2
14 1 9 1 11 13 14 3 13 10 9 0 9 11 2
21 9 1 9 7 4 1 0 9 13 0 9 2 15 15 1 0 9 1 11 13 2
38 1 0 12 9 2 3 13 0 9 9 7 0 9 11 2 13 7 9 9 1 9 0 9 7 9 9 1 9 9 2 1 15 15 1 9 3 13 2
37 1 12 0 9 2 15 13 1 0 9 1 9 11 0 9 2 15 1 10 9 0 11 13 0 9 1 0 0 9 2 7 1 0 9 7 9 2
22 9 0 9 11 1 9 7 9 2 15 3 13 1 11 2 15 13 9 1 9 0 9
4 9 11 2 11
8 0 9 4 13 13 9 7 9
5 11 2 11 2 2
14 0 9 13 9 9 9 1 9 12 2 12 9 9 2
16 9 9 13 2 16 4 10 9 4 13 1 9 1 0 9 2
21 1 15 2 3 4 13 4 0 9 13 2 15 1 0 9 13 9 10 0 9 2
22 9 11 11 11 15 13 2 16 9 13 2 16 4 15 0 9 3 10 9 13 9 2
18 9 11 11 11 13 13 2 16 9 3 13 0 2 7 13 3 0 2
12 3 3 9 15 2 16 13 1 9 0 9 2
10 13 1 9 0 7 0 9 2 13 2
21 16 4 13 0 12 9 3 3 13 2 3 1 11 1 9 2 15 13 9 9 2
10 9 11 11 11 13 10 9 1 0 2
37 1 1 15 2 16 1 10 9 11 13 9 9 2 9 7 9 2 13 1 11 13 2 16 4 11 13 2 16 4 0 9 13 3 1 10 9 2
32 9 0 9 11 2 11 11 11 15 13 2 16 16 9 9 1 10 9 13 2 15 15 13 0 0 9 2 13 15 3 9 2
22 9 1 15 4 15 13 0 9 2 7 16 1 0 9 13 12 9 1 9 0 9 2
11 0 9 4 13 1 9 9 1 9 9 2
15 9 11 3 13 2 16 15 1 10 9 13 1 0 9 2
17 13 2 16 4 1 0 9 13 13 0 9 1 15 1 0 9 2
20 13 4 15 1 9 9 2 16 4 15 1 9 13 1 9 0 9 2 13 2
8 9 1 11 11 2 9 11 2
26 1 11 4 13 2 16 0 9 9 11 1 9 2 3 13 1 0 9 2 4 13 13 0 2 9 2
11 1 10 9 13 7 10 4 13 9 9 2
15 1 9 1 0 9 13 0 0 9 0 9 13 10 9 2
9 9 13 2 15 13 10 9 13 2
17 13 15 7 13 9 2 15 10 9 13 2 16 9 13 3 0 2
16 1 0 7 0 9 11 2 3 13 9 2 15 9 13 15 2
23 7 3 2 3 13 0 9 2 3 1 11 7 1 11 2 9 0 9 13 0 9 11 2
25 13 1 9 2 15 15 13 1 9 2 13 0 9 1 0 11 7 13 0 13 1 9 0 9 2
27 13 2 16 15 1 9 0 0 0 9 13 2 16 16 15 10 9 1 9 13 2 13 4 13 1 0 2
3 2 11 2
1 9
14 9 13 12 9 2 16 13 1 0 9 1 9 9 2
9 13 3 12 9 11 7 0 9 2
4 0 4 13 0
2 11 11
11 0 9 13 1 0 2 15 13 0 9 2
9 13 0 2 15 15 3 13 0 9
11 1 9 12 7 12 13 1 12 0 9 2
9 0 0 9 13 1 12 10 9 2
21 3 13 14 12 0 0 9 2 15 13 1 0 0 9 7 9 1 12 12 9 2
13 3 13 2 1 1 0 9 2 1 12 0 9 2
28 1 0 9 1 9 9 9 10 9 0 9 13 9 0 9 2 7 15 1 9 12 9 1 0 0 9 9 2
23 3 13 9 7 9 2 10 9 13 1 0 9 7 4 13 2 3 9 1 9 12 9 2
9 0 9 15 4 13 1 12 9 9
31 11 13 9 12 9 7 1 9 9 1 9 0 12 2 9 12 1 11 2 7 1 9 0 9 0 1 9 9 7 9 2
39 9 11 15 3 13 13 9 1 9 12 9 0 9 9 9 1 9 0 11 7 0 7 0 11 2 15 3 13 1 11 2 11 7 11 7 13 9 9 2
12 11 3 13 0 9 1 9 0 9 0 9 2
20 9 2 16 9 0 11 13 3 13 1 9 0 9 2 13 1 0 9 3 2
24 3 1 9 12 13 0 9 0 9 9 1 9 2 10 9 9 13 1 12 2 12 2 12 2
10 0 0 9 11 7 9 10 9 13 2
13 15 9 9 1 10 0 9 4 1 0 9 13 2
22 0 9 1 9 13 1 9 2 16 11 13 14 1 9 12 1 0 9 11 0 9 2
8 9 11 13 14 9 0 9 2
7 11 13 9 12 9 9 2
24 9 2 11 11 2 9 0 9 9 1 9 4 15 13 2 13 15 1 9 3 1 9 12 2
44 1 9 12 4 13 2 16 4 15 15 13 13 3 7 1 0 9 7 9 11 11 2 15 13 0 2 0 9 2 13 2 2 13 10 0 9 2 16 4 15 15 3 13 2
13 3 4 13 2 15 15 13 7 15 1 15 13 2
8 15 4 3 13 7 0 9 2
7 11 1 15 4 3 0 2
14 3 1 9 12 13 9 11 2 16 13 3 0 9 2
7 1 10 9 0 9 13 2
19 13 3 0 9 1 9 1 15 2 16 15 13 2 10 9 7 15 13 2
7 9 4 13 1 9 2 2
6 13 15 15 1 9 2
9 3 15 13 13 1 9 2 12 2
16 9 4 13 13 7 15 2 16 11 1 15 4 13 0 9 2
20 9 1 0 9 13 2 1 9 1 11 2 15 15 1 9 0 9 15 13 2
20 0 9 13 0 13 12 0 7 12 0 9 16 0 9 1 9 12 9 9 2
13 1 9 13 2 1 0 15 9 4 9 9 13 2
17 1 0 9 9 11 3 13 15 0 2 16 16 13 9 0 9 2
5 9 9 15 13 2
18 13 15 2 13 10 9 13 1 12 9 9 2 15 13 0 9 2 2
13 15 13 1 15 2 15 13 1 9 7 15 14 2
10 9 0 9 2 7 13 15 3 3 2
6 3 15 13 7 0 2
20 3 1 9 12 13 1 0 9 10 11 2 15 15 1 11 3 13 1 9 2
10 4 3 13 7 7 0 9 13 0 2
12 7 15 13 10 9 7 11 15 13 1 9 2
5 13 3 12 9 2
13 3 3 10 9 13 2 16 3 13 0 9 2 2
16 3 13 13 2 16 0 9 13 9 0 1 0 7 0 9 2
11 13 9 9 2 15 13 1 9 12 9 2
5 13 3 1 9 2
15 15 10 9 13 7 3 15 13 9 2 16 13 0 9 2
19 13 3 13 2 15 13 9 2 15 13 9 7 15 15 1 9 14 13 2
2 14 2
12 13 9 2 15 13 9 2 16 13 3 9 2
5 13 15 0 9 2
13 16 13 2 16 15 13 13 2 7 13 15 9 2
11 16 15 13 3 2 7 15 13 0 9 2
18 9 13 2 16 11 13 3 0 1 9 9 2 1 15 4 9 13 2
10 0 3 3 13 1 0 0 0 9 2
9 1 0 15 15 7 13 13 2 2
14 13 15 3 9 2 16 9 4 13 1 9 0 9 2
2 14 2
13 13 2 16 3 13 9 1 12 7 12 9 11 2
13 3 13 2 16 9 13 4 13 3 1 9 12 2
4 13 4 15 2
9 13 7 2 16 0 9 13 11 2
63 0 9 7 9 9 2 16 3 1 9 9 11 16 0 9 0 0 9 2 7 3 1 9 9 0 9 1 9 12 2 7 7 1 10 9 2 14 16 13 1 10 0 9 2 7 10 9 13 1 15 9 9 0 7 0 2 9 9 9 1 9 2 2
7 3 4 13 9 10 9 2
4 11 1 0 9
3 0 11 2
22 3 16 12 9 9 7 0 9 13 1 10 9 0 0 9 11 2 0 9 7 9 2
33 9 7 9 9 11 11 13 2 16 11 1 12 9 13 1 9 11 11 2 0 9 9 2 0 0 0 9 1 10 9 1 11 2
25 3 1 10 9 13 9 0 9 9 0 9 2 15 4 13 10 9 13 1 0 9 2 13 11 2
8 13 15 13 1 10 0 9 2
26 9 9 13 13 2 16 13 1 15 13 7 3 2 1 0 9 2 1 9 7 1 0 9 2 13 2
15 0 9 1 15 13 3 0 9 2 0 1 9 0 9 2
12 3 15 11 13 12 2 10 9 7 3 13 2
20 9 2 1 15 3 13 2 13 0 9 2 0 9 2 0 9 7 0 9 2
20 3 0 9 9 3 13 2 7 13 1 15 9 9 7 9 9 2 13 11 2
26 0 9 2 3 3 13 0 9 9 2 13 9 11 11 3 13 9 2 15 11 13 1 0 0 9 2
14 13 3 1 0 9 7 3 15 15 13 12 12 9 2
20 13 4 0 9 0 9 9 1 0 9 2 1 10 9 15 13 2 13 11 2
1 3
24 0 7 0 9 1 9 9 1 11 11 1 0 9 15 1 9 9 13 1 0 9 1 11 2
20 1 9 15 13 1 12 2 1 12 2 9 7 1 12 2 1 12 2 9 2
12 9 13 1 9 1 9 1 12 1 12 9 2
23 9 0 0 9 4 3 1 9 12 9 9 2 9 9 7 9 13 1 11 1 0 9 2
12 9 1 12 9 13 1 9 9 16 9 9 2
34 1 9 9 13 1 9 1 0 9 9 9 9 9 9 0 9 7 9 0 9 0 9 1 11 1 11 2 15 13 14 1 9 9 2
25 1 9 9 11 4 1 9 1 0 9 0 9 9 7 9 13 9 1 9 0 0 9 11 11 2
54 3 9 9 2 9 7 9 13 11 2 15 13 1 9 12 1 0 9 2 16 9 9 1 0 9 2 9 9 7 9 2 3 1 0 9 2 7 3 10 9 1 11 2 3 1 9 12 13 1 9 0 9 11 2
10 0 9 8 2 8 2 8 2 8 2
1 9
2 11 11
9 0 9 13 7 13 3 0 9 2
11 12 13 0 7 16 13 2 13 3 13 2
33 1 0 9 2 9 1 0 9 8 2 8 2 8 2 8 2 2 15 0 9 15 1 0 9 13 3 3 3 13 1 9 11 2
21 8 2 8 2 8 2 8 2 13 9 9 0 0 9 3 1 9 1 0 9 2
25 9 11 11 1 15 1 9 12 13 0 0 9 2 15 13 0 9 7 13 10 9 7 9 9 2
12 0 9 13 1 9 2 9 7 9 1 9 2
23 3 13 0 0 9 2 3 1 11 2 7 9 9 13 15 2 16 13 13 0 9 0 2
14 0 9 1 0 9 2 3 9 13 9 7 9 0 2
9 0 9 1 9 7 1 0 9 2
17 11 15 13 14 13 9 1 0 9 1 0 0 9 1 0 9 2
12 15 9 2 15 12 0 9 2 0 7 3 2
29 12 0 9 2 9 0 11 11 7 11 11 2 13 15 0 2 14 14 10 0 0 2 1 10 9 0 0 9 2
13 13 1 3 0 9 7 13 1 15 9 1 9 2
21 1 15 7 13 7 12 0 0 9 2 1 0 0 9 2 9 7 9 0 9 2
22 1 12 0 9 3 13 9 0 0 9 7 3 13 13 0 9 10 0 9 11 11 2
10 15 9 13 0 9 2 13 0 9 2
25 16 3 13 10 9 3 0 7 0 2 3 15 13 10 9 2 0 1 11 1 9 12 7 12 2
10 13 0 9 13 1 12 9 1 9 2
9 7 15 1 9 3 13 1 9 2
7 13 0 9 0 1 9 2
10 3 13 2 16 7 15 13 0 9 2
4 13 0 9 2
37 13 9 2 1 15 1 0 9 0 0 9 1 0 9 0 9 1 0 0 9 13 0 9 1 3 0 9 2 15 9 13 11 7 9 0 11 2
6 9 15 13 13 3 2
9 1 0 9 2 7 0 0 9 2
3 3 1 9
15 9 2 9 0 9 2 12 1 9 1 9 2 12 9 2
3 0 9 2
5 9 11 13 9 11
5 11 2 11 2 2
28 9 11 11 11 11 13 1 0 9 11 1 0 11 0 0 9 2 16 4 1 10 9 13 9 0 9 9 2
29 9 15 1 15 13 0 9 3 0 9 0 0 9 0 9 2 4 15 13 9 7 4 13 1 9 1 0 9 2
22 1 0 9 13 0 9 1 15 3 13 7 1 9 15 13 14 1 0 9 1 11 2
32 1 9 2 3 15 3 13 1 10 9 2 13 2 3 13 2 3 15 1 10 9 9 13 2 7 3 15 15 14 3 13 2
23 13 15 16 15 0 2 3 16 4 15 1 0 9 13 15 9 2 1 15 4 13 9 2
20 1 9 0 9 15 9 2 11 1 0 9 13 0 9 2 7 15 13 0 2
7 3 9 13 1 9 3 2
38 13 4 9 11 2 15 13 0 9 2 7 13 4 1 15 2 10 13 9 2 16 13 0 2 16 15 9 1 9 13 13 7 0 9 16 0 9 2
26 13 4 9 7 1 15 13 10 9 1 9 2 7 1 0 9 2 15 4 13 2 15 15 13 2 2
5 3 13 10 9 2
14 13 9 1 10 9 13 7 1 0 9 15 13 13 2
18 13 15 9 2 16 1 11 13 13 7 16 0 13 13 9 1 9 2
13 13 15 0 9 1 9 12 0 9 0 9 0 2
6 9 11 2 11 2 11
2 9 9
26 13 2 16 1 10 9 13 7 15 2 10 0 9 15 13 13 9 7 10 9 2 15 13 9 9 2
12 10 10 9 13 13 7 13 15 1 9 9 2
18 14 2 0 9 9 9 15 3 13 0 9 9 2 16 0 9 9 2
35 13 2 14 1 10 9 2 16 1 0 9 13 9 9 0 9 2 13 15 7 13 9 1 9 9 7 15 15 13 9 9 0 15 9 2
16 10 9 13 0 13 3 9 9 2 15 13 3 0 9 9 2
14 1 0 9 7 13 2 16 10 9 9 9 3 13 2
24 16 0 9 13 2 7 13 1 0 9 2 13 2 14 2 10 9 2 3 15 9 9 13 2
9 7 13 2 16 4 15 11 13 2
24 9 1 9 13 3 1 9 1 9 9 11 1 9 2 11 2 9 2 9 11 12 12 11 12
7 1 11 15 9 0 9 13
5 11 2 11 2 2
11 9 0 9 0 11 11 15 1 9 13 2
31 1 0 9 13 4 9 2 15 9 13 12 9 9 2 13 1 9 12 2 9 2 3 10 9 2 3 1 11 13 11 2
23 0 13 2 16 4 10 9 13 16 1 11 2 3 15 13 13 3 3 7 9 15 13 2
33 13 2 16 4 15 3 0 9 3 13 1 0 9 2 7 1 0 9 13 1 0 9 2 13 9 11 7 3 0 9 11 11 2
19 0 9 15 1 11 13 1 12 2 9 1 9 12 2 9 1 0 11 2
32 13 3 3 12 9 2 16 1 0 9 9 11 13 1 11 2 7 4 13 12 2 9 13 1 11 11 2 13 11 2 11 2
6 13 15 11 1 11 2
6 9 9 13 9 0 9
4 9 9 0 9
5 11 2 11 2 2
26 3 4 3 13 13 1 0 9 9 7 13 1 15 13 2 13 0 9 11 9 11 10 9 11 11 2
17 1 15 13 9 3 13 7 12 2 9 13 1 9 13 0 9 2
23 9 9 11 2 11 2 7 11 2 11 2 4 13 13 13 1 0 9 9 11 2 11 2
26 9 1 11 11 2 13 15 1 11 2 13 9 9 1 11 2 7 3 15 13 1 11 11 1 11 2
28 0 9 11 1 0 9 13 9 2 15 1 9 11 11 1 9 1 11 2 0 9 11 2 3 13 1 9 2
16 0 9 4 13 13 7 11 11 1 11 2 9 0 0 9 2
26 1 9 9 13 11 3 9 9 9 11 11 1 11 2 15 4 13 9 3 13 1 0 9 9 14 2
30 9 9 11 11 13 2 16 1 9 9 9 1 9 3 13 13 2 0 0 9 15 13 13 9 14 1 12 2 9 2
19 1 10 9 13 2 16 4 15 1 11 13 1 12 9 3 13 9 11 2
17 1 11 15 13 9 7 1 10 9 15 3 13 13 14 1 9 2
15 16 15 3 13 2 3 13 9 1 10 9 2 13 11 2
38 11 13 2 16 0 2 1 11 11 11 2 3 0 11 15 3 13 1 0 9 11 7 13 1 0 2 11 2 3 15 1 0 9 3 13 0 9 2
9 3 15 13 13 0 9 3 13 2
10 11 11 15 7 1 0 9 13 13 2
9 9 13 2 16 4 15 0 13 2
1 3
13 9 0 9 1 11 4 13 3 13 9 12 9 2
20 13 15 1 9 0 0 9 2 15 13 3 12 9 1 9 9 9 9 11 2
22 11 4 1 0 9 1 0 9 11 11 13 1 12 9 13 9 9 9 1 0 9 2
4 0 11 13 9
12 16 15 9 13 13 1 9 2 4 13 16 9
3 11 11 2
17 1 0 9 11 11 11 13 10 9 1 0 0 0 0 9 9 2
23 0 0 9 2 0 3 1 9 2 13 0 2 7 13 0 9 0 3 12 9 9 9 2
34 0 0 9 15 13 1 9 9 0 0 9 9 1 9 2 15 13 0 9 1 9 12 7 1 15 15 9 13 1 9 0 9 9 2
29 16 13 9 9 11 11 2 9 13 1 9 9 9 7 9 11 1 9 2 16 13 0 13 1 0 0 9 9 2
8 3 15 9 13 13 1 9 2
18 16 15 15 15 13 2 4 13 3 16 0 9 0 9 10 0 9 2
9 13 1 10 9 13 7 9 11 2
19 1 9 0 9 1 9 13 9 1 9 2 1 15 0 9 13 7 9 2
27 11 2 15 13 1 9 0 9 10 0 9 1 12 0 9 2 1 0 9 13 12 9 7 13 10 9 2
14 13 3 13 10 9 2 15 9 9 7 9 3 13 2
19 3 9 9 13 9 2 1 10 9 15 7 1 15 13 13 2 13 11 2
33 10 9 2 1 15 13 1 12 9 9 3 9 2 13 11 13 9 0 1 9 9 7 9 9 10 0 9 2 15 15 13 9 2
18 11 2 10 0 9 13 12 9 9 2 4 13 1 0 9 0 9 2
19 3 12 9 9 13 0 9 2 12 7 9 9 11 7 9 13 0 9 2
8 3 13 0 9 12 9 9 2
4 9 13 1 11
2 11 2
20 16 4 13 0 0 9 2 13 9 11 11 12 2 9 11 0 1 10 9 2
25 11 13 2 16 9 3 13 2 16 13 13 0 9 1 9 2 1 15 4 15 13 1 11 13 2
8 9 13 9 1 0 0 9 2
10 9 11 11 11 13 1 9 11 9 2
13 1 10 9 13 9 9 11 11 2 0 1 9 2
24 1 9 11 4 1 0 9 13 12 9 11 1 0 9 2 3 13 1 9 13 9 1 9 2
2 9 2
2 11 11
27 9 12 13 0 7 0 9 14 0 7 0 11 2 7 7 15 2 15 15 0 0 9 12 9 3 13 2
25 9 12 13 0 7 0 9 7 0 9 2 15 13 3 7 3 7 1 0 0 9 13 10 9 2
13 15 13 15 3 9 11 7 15 15 1 15 13 2
21 0 9 13 1 10 0 9 1 0 9 0 9 2 0 11 7 9 1 0 9 2
6 15 13 0 0 9 2
3 10 9 2
3 10 9 2
14 15 4 1 0 11 13 9 9 2 15 9 0 9 2
24 0 11 2 9 0 2 0 9 1 9 0 9 2 15 13 9 2 15 13 0 9 0 9 2
10 13 1 15 9 11 7 0 9 11 2
53 1 9 0 9 15 13 12 2 12 7 3 12 9 2 15 13 13 2 0 4 0 13 1 9 2 15 7 13 14 12 0 2 13 0 9 9 0 9 7 9 2 15 7 0 0 9 1 12 9 1 15 13 2
15 9 1 9 13 7 1 10 9 13 7 0 2 7 0 2
14 9 13 13 9 1 9 7 13 1 10 0 9 9 2
37 13 15 9 2 9 13 2 9 3 13 1 0 7 1 10 9 13 0 2 0 2 3 14 0 9 3 7 3 0 2 15 4 13 9 0 9 2
27 13 15 16 1 10 9 2 9 13 9 2 13 3 1 9 7 6 2 1 9 13 0 9 7 0 9 2
5 9 15 14 13 2
14 15 0 13 0 9 9 2 15 3 15 13 9 0 2
40 1 9 15 3 13 0 9 0 9 2 13 3 10 3 0 9 7 0 9 9 15 4 3 13 1 0 9 2 3 15 14 0 13 0 7 0 9 9 9 2
16 15 13 9 0 9 2 0 0 9 2 9 2 9 7 9 2
12 13 7 9 0 2 0 2 1 0 9 9 2
8 13 7 9 1 9 0 9 2
17 1 15 3 15 15 13 0 2 9 13 0 7 9 12 13 9 2
6 9 13 7 3 0 2
9 9 13 0 0 9 7 0 9 2
19 1 10 9 15 13 2 0 9 3 1 11 13 9 2 0 0 9 9 2
9 10 9 13 13 2 9 1 9 2
7 9 11 13 7 10 9 2
3 7 3 2
12 9 1 0 9 2 1 15 13 13 9 9 11
5 9 11 11 2 11
22 0 9 0 9 11 11 3 13 1 9 11 1 11 7 0 9 1 9 9 11 11 2
22 11 13 2 16 7 0 9 13 1 9 1 9 7 11 3 13 7 13 13 0 9 2
20 1 9 15 13 3 1 9 9 11 11 7 13 1 15 9 1 9 7 9 2
5 9 11 11 2 11
5 0 9 1 11 2
3 1 0 9
5 11 2 11 2 2
37 3 2 3 2 3 2 3 13 0 9 9 0 9 2 15 13 1 0 9 1 11 7 13 12 0 9 2 11 2 11 2 11 2 11 7 11 2
14 13 15 1 0 0 9 9 0 9 0 9 0 9 2
30 9 9 11 11 13 9 2 16 4 15 10 9 13 13 9 1 9 0 0 0 9 7 3 9 9 1 0 9 12 2
28 0 9 11 1 9 13 2 16 9 10 0 9 15 14 3 13 0 9 12 5 12 2 15 1 9 13 11 2
1 9
16 12 9 4 13 1 9 0 2 11 1 0 9 1 11 12 2
18 1 0 9 9 13 11 2 15 15 13 13 0 9 1 9 12 9 2
10 9 4 13 1 9 7 13 1 9 2
19 0 9 2 0 11 2 4 13 2 16 15 13 3 0 9 1 12 9 2
7 7 15 13 1 0 9 2
1 3
17 0 9 9 9 12 9 0 9 7 9 0 9 13 3 1 11 2
9 9 15 13 1 9 0 0 9 2
14 11 13 13 9 9 2 9 7 0 9 1 9 11 2
36 0 9 1 9 1 9 0 9 2 9 7 9 9 13 3 1 11 0 9 11 11 7 0 9 11 11 2 11 2 15 13 1 9 1 11 2
38 0 9 13 3 1 11 2 7 16 4 13 0 9 2 7 2 16 10 9 13 15 2 13 9 2 13 3 0 9 1 11 2 1 2 11 11 11 2
16 1 12 12 0 9 13 1 9 1 0 9 11 9 7 9 2
10 11 13 9 0 9 9 11 11 11 2
17 13 3 13 2 16 4 13 14 1 9 1 9 9 12 2 9 2
39 1 0 0 9 1 11 13 1 9 1 9 1 9 11 2 3 4 13 0 9 11 11 2 12 2 2 15 13 0 0 9 1 0 9 0 1 9 9 2
12 1 9 1 9 1 11 7 11 15 13 11 2
30 11 13 2 16 4 11 9 1 9 0 9 13 9 1 0 9 7 1 0 9 7 16 4 10 9 13 1 0 11 2
10 10 9 3 13 9 0 9 11 11 2
14 13 13 0 9 1 0 9 7 13 9 1 0 9 2
29 1 0 0 9 11 15 10 9 3 13 9 0 0 9 2 15 3 13 12 9 9 2 3 12 9 0 9 2 2
15 1 0 9 15 3 3 15 13 13 0 0 9 2 9 2
9 9 1 9 9 0 9 2 12 2
95 11 13 9 0 9 7 13 15 1 10 9 2 2 15 13 9 1 9 9 1 10 9 2 2 1 10 9 13 0 9 2 2 1 10 9 13 0 9 2 2 1 15 15 13 13 9 2 1 9 2 7 0 9 2 2 15 13 0 9 2 9 1 9 12 2 2 2 9 9 9 7 0 9 2 2 9 9 2 15 15 13 2 7 15 15 13 2 3 2 0 9 1 10 9 2
11 11 2 0 9 2 11 2 9 2 11 11
24 1 9 11 2 1 0 9 11 2 9 0 9 2 9 7 9 2 13 9 1 9 16 3 2
34 9 13 9 3 0 9 9 2 3 9 1 9 9 1 9 2 9 0 9 2 3 3 0 0 9 0 9 7 0 9 0 9 9 2
24 9 1 9 13 0 0 9 2 15 13 1 10 9 9 2 7 1 9 3 1 12 12 9 2
25 1 11 15 3 13 3 9 2 15 3 13 2 3 9 1 11 2 11 2 0 11 7 0 11 2
28 0 9 13 3 1 9 1 0 9 1 9 1 9 2 1 0 9 7 3 13 0 9 9 1 3 0 9 2
32 1 15 0 9 13 1 9 2 0 9 2 9 2 9 1 0 9 2 1 0 9 2 9 2 9 1 9 7 9 1 9 2
12 9 9 1 11 15 3 13 1 9 7 9 2
6 13 3 1 0 9 2
10 1 0 9 3 13 0 12 9 9 2
38 1 9 12 5 12 15 9 13 3 1 12 1 12 12 2 1 9 12 5 12 1 12 1 12 12 7 1 9 12 5 12 1 12 1 12 12 9 2
13 0 9 1 9 11 13 14 1 12 12 9 0 2
23 0 9 15 1 11 13 3 1 12 9 0 9 2 1 9 1 9 12 2 12 9 9 2
10 15 15 13 1 9 1 12 12 9 2
26 0 9 13 0 0 9 2 3 1 0 9 2 1 9 1 12 1 12 9 9 2 15 13 3 0 2
14 16 15 13 2 7 1 9 1 12 7 12 12 9 2
37 3 15 13 0 9 2 3 1 0 9 2 3 9 0 0 9 1 0 9 13 14 1 12 9 2 1 0 9 7 9 13 1 12 7 12 9 2
52 9 9 9 1 9 9 2 3 3 13 2 3 1 0 9 2 15 13 1 12 1 12 9 2 9 12 2 1 0 9 3 1 12 1 12 9 2 9 12 2 16 1 0 9 13 9 1 9 0 3 3 2
14 10 0 9 13 9 9 0 9 11 2 11 7 11 2
15 1 9 15 13 9 1 9 12 2 12 9 0 9 9 2
12 10 9 13 0 9 9 7 10 9 1 11 2
17 0 13 3 15 2 16 15 7 13 9 0 9 1 10 9 9 2
9 0 9 13 3 1 9 0 9 2
24 0 9 11 3 13 1 0 0 9 7 1 11 2 7 13 7 0 9 13 0 9 7 9 2
8 10 9 13 9 0 0 9 2
30 16 13 9 0 15 13 2 13 9 13 3 3 7 1 9 1 0 9 0 9 1 9 2 15 15 13 0 9 9 2
7 11 11 2 0 9 2 12
5 9 11 11 2 11
10 9 11 9 13 0 9 9 12 2 12
23 9 11 11 1 10 0 9 13 1 9 12 2 9 1 9 1 9 9 12 2 12 11 2
23 10 0 9 11 2 13 15 11 2 13 0 3 0 7 0 9 7 9 7 0 0 9 2
13 1 9 13 10 0 9 3 0 2 0 7 0 2
16 0 9 15 13 7 9 11 9 2 0 0 2 0 9 11 2
19 10 9 13 13 1 3 0 9 0 9 2 3 0 9 7 0 0 9 2
29 1 0 9 2 15 13 3 2 9 1 0 9 2 15 7 11 13 0 2 3 0 9 7 9 0 7 0 9 2
19 3 7 9 9 7 9 11 11 2 15 10 9 13 9 9 3 0 9 2
10 0 9 0 0 3 1 15 13 11 2
14 9 11 11 7 11 0 9 12 2 12 11 3 13 2
24 16 3 13 11 9 9 11 11 2 1 12 2 9 13 1 0 9 13 9 0 0 9 11 2
22 1 9 1 9 9 9 13 12 2 7 12 2 9 9 11 11 2 9 0 0 11 2
26 1 9 9 1 9 9 13 0 9 11 2 9 2 15 15 0 9 11 13 9 0 0 9 1 9 2
18 16 0 9 2 12 2 9 2 13 12 2 12 11 9 0 0 11 2
23 0 13 3 9 0 2 0 2 0 2 2 15 15 13 1 0 9 12 2 9 0 9 2
11 13 15 0 0 9 11 2 11 2 11 2
3 2 11 2
11 15 13 1 11 9 2 13 13 1 9 2
14 13 1 15 3 9 0 9 2 7 9 13 0 9 2
6 9 11 2 11 2 11
5 0 9 14 1 9
5 11 2 11 2 2
40 14 1 9 13 13 0 0 0 9 0 0 9 11 2 12 5 2 7 12 0 9 2 12 5 2 2 15 3 1 0 12 13 1 9 0 9 1 9 9 2
14 3 13 3 9 9 2 10 0 9 13 12 9 9 2
30 9 4 13 10 9 0 9 2 0 9 1 0 9 2 0 9 1 9 2 0 9 7 1 0 9 9 7 0 9 2
40 9 9 2 3 13 10 9 2 13 0 9 9 2 3 0 0 9 9 9 1 9 1 0 9 2 0 9 1 9 9 9 2 0 0 9 7 9 9 9 2
17 1 9 9 4 13 0 9 2 1 15 13 3 3 12 12 9 2
5 9 9 13 3 13
2 11 2
15 0 9 9 15 1 0 9 1 9 13 1 0 0 9 2
19 0 9 1 9 0 9 13 9 0 9 1 9 9 3 1 12 9 9 2
18 0 9 3 3 13 9 9 0 9 1 12 9 1 12 9 1 9 2
12 13 15 3 14 9 1 0 0 9 12 9 2
22 0 9 13 3 13 9 9 0 1 9 7 1 0 9 2 16 4 3 13 0 9 2
23 1 9 0 9 9 9 13 2 16 1 1 9 1 9 9 1 10 9 13 13 1 9 2
26 1 0 0 9 11 4 9 0 0 9 13 0 0 9 2 15 13 0 9 9 9 2 13 9 11 2
19 0 0 9 0 11 13 1 10 0 9 0 9 2 10 9 13 3 0 9
5 9 11 11 2 11
8 11 15 13 1 11 11 2 12
2 11 2
28 0 9 11 4 13 1 0 9 11 11 2 12 2 15 15 13 1 12 2 12 2 1 12 2 12 2 12 2
23 0 9 15 13 1 9 9 9 2 3 4 13 10 9 0 12 9 2 1 15 12 0 2
21 16 3 13 0 9 0 9 11 11 2 9 13 0 9 1 9 7 9 10 9 2
14 11 4 13 1 11 3 1 9 12 9 0 0 9 2
16 0 9 1 9 2 9 7 9 9 4 9 13 1 12 9 2
15 9 13 13 0 9 11 16 0 0 9 1 9 0 9 2
16 13 4 3 13 9 0 0 9 7 13 9 1 0 9 9 2
14 1 9 13 9 0 9 11 2 0 9 1 0 9 2
5 1 0 9 3 13
5 11 2 11 2 2
30 16 9 0 9 13 3 14 3 1 9 2 3 13 1 9 1 15 2 1 15 13 9 1 3 0 9 9 0 9 2
33 9 11 11 1 10 9 13 2 16 9 9 9 2 15 13 1 9 9 12 2 12 2 15 1 9 9 1 0 9 13 3 13 2
30 9 0 9 3 1 9 13 9 0 9 2 1 15 1 9 1 9 0 9 13 9 9 0 9 1 9 0 11 11 2
11 10 9 7 13 9 11 7 12 9 9 2
8 9 13 9 9 0 9 1 9
5 11 2 11 2 2
19 0 9 13 3 13 9 0 9 7 9 9 2 15 9 1 9 13 9 2
33 0 9 2 1 15 13 13 12 9 2 9 0 9 7 9 10 0 9 2 15 1 0 9 13 1 0 12 9 3 16 0 9 2
10 9 1 0 9 9 13 0 0 9 2
15 13 3 2 16 12 9 15 0 9 13 9 1 12 9 2
21 3 15 9 9 13 1 0 9 12 12 9 7 12 12 15 15 3 13 1 9 2
11 9 9 1 11 13 12 1 0 1 9 2
9 13 15 9 1 9 9 9 0 2
7 13 15 9 7 0 9 2
5 13 15 0 9 2
15 0 3 0 9 4 13 1 9 0 2 0 7 1 11 2
13 9 15 1 10 9 13 9 10 9 7 13 9 2
27 9 13 3 15 2 16 0 9 1 9 9 7 10 9 13 1 15 9 2 7 16 9 9 13 1 9 2
11 9 13 2 16 0 9 9 13 0 9 2
26 9 3 13 3 2 16 9 13 0 2 9 9 1 9 7 1 9 9 15 13 9 1 0 9 2 2
20 9 7 13 9 0 9 1 9 9 2 0 1 9 9 1 11 7 0 11 2
9 10 9 15 13 13 3 1 9 2
20 9 13 13 9 3 0 9 7 13 9 1 0 7 9 1 10 9 1 9 2
10 9 9 4 15 13 13 1 9 12 2
5 9 15 13 1 9
5 11 2 11 2 2
27 0 9 2 9 2 9 7 0 9 13 1 0 9 0 9 1 11 12 9 0 9 1 9 1 12 9 2
18 1 9 13 1 9 1 12 2 9 3 2 16 1 9 13 0 9 2
18 0 9 15 9 13 1 10 9 1 15 2 16 15 15 13 1 9 2
20 15 12 9 4 13 1 0 9 9 2 9 15 0 9 4 13 1 12 9 2
5 9 2 0 0 9
2 11 11
38 9 13 15 0 2 13 15 13 2 0 9 2 15 13 13 1 0 9 2 3 11 2 3 11 2 2 13 1 9 13 14 3 0 9 10 0 9 2
21 0 9 15 3 9 7 13 7 10 9 13 9 3 9 16 0 12 9 10 9 2
25 1 0 9 7 3 4 13 0 9 0 9 1 9 10 9 9 2 15 9 1 11 4 13 13 2
21 16 13 0 9 2 16 3 3 0 13 2 13 9 0 2 15 15 9 3 13 2
18 0 9 11 11 15 1 15 13 3 2 9 9 15 13 0 9 9 2
6 10 9 13 0 9 2
14 7 15 15 9 13 3 0 9 10 9 1 0 9 2
28 3 1 0 11 2 3 4 15 13 15 13 7 13 0 9 0 9 2 7 1 11 2 1 10 0 9 11 2
65 0 9 7 9 0 9 11 11 13 1 9 9 9 2 9 9 2 3 0 9 2 9 9 13 12 1 3 0 9 0 9 2 2 2 13 15 1 0 9 9 0 9 2 2 2 7 3 3 2 16 15 7 10 9 13 2 7 14 9 2 15 13 0 9 2
45 9 13 3 2 3 15 13 1 9 7 9 9 2 10 9 3 4 13 1 9 2 7 3 9 2 10 9 1 9 13 0 7 15 13 3 7 3 3 9 1 9 13 1 9 2
21 9 9 2 9 2 9 7 0 9 2 3 2 11 13 0 9 2 13 9 9 2
34 3 13 15 7 11 11 2 16 13 2 16 9 2 9 7 9 0 0 9 13 13 0 2 16 4 13 1 10 9 2 7 3 0 2
28 3 13 0 9 0 2 3 3 0 2 1 10 9 13 0 0 9 2 13 9 0 1 3 0 7 0 9 2
5 13 0 9 0 2
12 15 15 13 9 2 9 7 9 2 3 3 2
12 15 13 7 14 0 2 7 14 0 9 9 2
28 0 9 2 0 2 14 0 9 10 9 7 10 9 15 13 1 10 9 7 3 1 10 9 3 1 15 13 2
8 0 9 9 13 0 7 3 2
12 0 9 2 9 7 9 13 9 0 7 3 2
18 3 9 0 9 13 1 0 9 2 1 15 1 0 9 13 10 9 2
13 14 1 0 0 9 13 3 0 14 12 12 9 2
15 1 0 0 9 3 14 12 9 2 15 2 0 2 0 2
11 7 3 13 1 11 0 3 14 11 15 2
6 15 0 2 0 15 2
27 9 9 2 1 15 15 0 13 13 9 9 1 10 9 7 13 15 16 9 9 2 15 13 13 3 3 2
13 1 10 9 13 9 9 15 9 9 0 9 3 2
13 13 3 13 0 9 2 1 10 9 15 13 9 2
8 3 0 2 15 15 13 13 2
10 13 7 15 0 2 15 1 9 13 2
7 9 1 9 7 1 9 2
32 1 0 9 7 13 0 9 1 9 11 3 0 9 2 15 13 1 0 9 11 2 9 9 11 2 2 15 13 1 9 11 2
19 15 13 13 9 2 0 12 9 0 9 2 15 13 13 9 2 0 11 2
5 16 15 13 11 2
14 16 4 15 13 12 9 2 15 4 14 3 13 13 2
4 9 13 0 9
9 1 0 9 1 0 9 13 0 9
2 11 11
4 13 10 9 2
25 15 10 9 13 2 13 2 9 13 2 13 1 0 9 0 9 9 7 9 3 0 9 11 11 2
10 0 9 1 9 7 3 3 0 13 2
16 1 9 13 0 9 0 0 9 2 15 1 9 3 13 9 2
20 9 13 16 9 2 0 9 3 1 0 9 13 1 0 9 7 9 0 9 2
6 11 13 16 13 9 2
2 3 2
5 9 13 1 9 2
28 9 10 0 0 9 3 13 9 3 0 0 9 11 11 11 2 9 1 0 3 2 0 9 1 0 0 9 2
16 0 9 9 9 2 15 1 0 9 3 13 1 9 2 13 2
16 1 0 0 9 1 11 15 13 9 1 0 9 13 3 3 2
24 11 3 1 11 2 15 13 9 0 9 9 14 1 9 12 2 13 3 1 9 0 0 9 2
30 9 0 9 2 9 2 15 13 3 0 9 16 0 9 2 15 15 13 13 0 9 1 0 12 9 1 0 12 9 2
13 0 9 11 3 13 7 0 9 15 13 1 12 2
26 1 9 0 9 13 1 12 9 9 9 1 10 0 9 11 11 1 11 1 9 9 2 12 9 2 2
17 13 15 2 16 0 9 15 13 12 2 9 13 1 3 0 9 2
9 9 9 15 7 9 3 13 13 2
21 16 1 10 9 13 12 9 2 13 15 11 2 0 9 0 9 2 1 9 9 2
7 0 9 13 13 1 9 2
11 11 13 10 9 9 9 7 13 9 13 2
19 3 15 13 9 1 9 2 10 9 12 1 9 3 3 13 0 0 9 2
12 13 1 15 2 16 15 9 1 9 15 13 2
16 3 3 2 1 9 1 0 9 9 13 9 14 0 9 9 2
5 1 0 9 13 2
22 9 13 13 7 0 0 9 11 11 2 3 9 0 9 2 2 16 0 9 3 13 2
19 9 3 1 9 9 13 2 16 1 0 9 13 9 7 0 9 15 0 2
16 0 9 1 11 2 0 9 9 2 3 10 0 9 13 13 2
13 3 13 2 16 4 0 9 0 9 1 9 13 2
17 16 15 15 10 9 3 3 13 13 2 0 9 9 3 3 13 2
11 9 9 2 15 13 1 9 2 13 9 2
22 1 0 9 0 9 1 11 13 13 10 9 2 15 13 3 9 16 15 10 9 3 2
14 1 11 4 1 9 0 9 0 9 13 12 9 9 2
18 10 9 4 13 1 12 9 3 9 2 16 4 13 15 0 9 3 2
6 1 11 13 0 9 2
37 1 10 9 13 3 14 12 9 9 9 2 16 7 1 0 9 11 13 1 0 12 9 9 2 13 15 0 9 9 2 1 15 13 14 12 0 2
10 1 0 9 4 15 13 12 2 9 2
24 13 1 9 0 9 2 4 1 9 13 3 7 13 7 1 0 9 1 0 12 9 13 15 2
7 0 11 15 10 9 13 2
31 13 14 0 9 10 9 2 3 13 7 0 9 2 15 11 3 1 9 12 2 3 13 0 9 9 2 13 9 1 9 2
14 9 1 9 9 1 15 13 7 9 9 1 0 9 2
17 9 11 1 9 0 1 0 0 9 2 9 1 12 2 9 12 2
5 9 9 2 9 9
12 0 0 7 0 9 13 9 2 13 9 11 11
2 11 11
53 0 9 9 1 0 9 2 15 3 3 3 13 9 9 7 15 0 9 3 13 2 15 13 3 0 9 7 9 11 11 2 9 0 9 1 0 9 2 0 9 2 9 7 9 10 10 9 1 0 9 0 9 2
30 1 0 9 13 11 11 2 0 1 9 12 2 1 0 10 0 0 9 1 0 9 2 3 9 9 1 0 9 0 2
8 10 0 9 13 0 2 13 2
4 9 1 9 13
48 1 10 9 1 11 2 11 2 11 2 11 2 11 2 11 7 0 2 3 1 11 7 11 1 11 2 13 10 0 0 9 0 0 9 2 3 15 13 0 9 11 11 2 3 9 0 9 2
30 0 4 15 1 15 13 2 0 9 1 9 15 3 1 11 1 15 13 9 10 9 9 7 9 11 11 2 12 2 2
35 13 9 0 9 2 15 4 15 13 13 0 9 2 13 11 2 7 1 15 15 3 13 3 0 9 9 7 9 2 15 15 13 7 9 2
18 7 16 9 0 9 3 15 1 15 13 7 10 0 9 3 15 13 2
17 13 7 0 9 2 16 15 13 1 0 0 9 2 13 3 0 2
20 1 9 13 13 9 1 9 11 11 2 1 15 15 11 13 1 9 0 9 2
16 9 15 13 3 1 9 12 2 1 9 9 1 0 9 13 2
23 1 12 9 11 13 7 1 9 1 9 7 13 14 1 15 2 16 4 9 13 3 9 2
9 7 3 15 15 7 13 3 13 2
4 11 11 7 0
11 11 11 13 1 9 0 9 1 9 11 2
31 3 1 15 1 12 9 9 0 9 13 7 9 1 0 2 3 15 15 13 2 9 11 2 2 2 9 1 0 0 9 2
13 3 15 3 1 9 12 1 0 9 13 9 11 2
19 1 9 11 11 2 15 3 13 1 10 0 9 2 4 7 13 1 9 2
19 15 7 0 9 1 10 9 13 2 9 1 10 9 13 9 12 2 13 2
17 16 4 3 13 1 11 2 13 4 9 13 15 7 1 0 9 2
30 13 4 1 9 11 11 2 15 13 9 0 9 7 3 15 3 15 0 13 1 9 2 14 1 9 2 7 13 15 2
19 13 4 1 9 11 11 7 13 4 1 10 0 9 15 1 15 15 13 2
24 9 3 0 2 3 0 9 11 11 2 11 11 2 11 11 7 0 13 1 11 3 14 3 2
12 3 0 13 15 1 10 9 0 9 11 11 2
4 9 7 9 13
13 1 9 12 9 1 0 9 7 0 9 14 13 2
22 13 14 9 2 7 7 9 2 13 11 2 10 9 11 11 13 0 9 1 0 9 2
27 1 10 9 2 15 4 3 13 13 7 15 4 3 13 1 9 2 13 2 16 15 10 9 13 15 10 2
21 13 3 0 9 2 1 0 0 9 2 3 15 15 3 13 2 15 15 3 13 2
22 0 9 15 3 1 11 13 1 9 9 0 9 2 13 4 13 10 0 0 0 9 2
9 1 0 12 9 15 13 0 9 2
8 3 15 10 9 13 1 9 2
11 3 15 7 13 2 16 15 15 0 13 2
26 0 13 1 11 3 9 9 2 0 7 0 1 9 16 0 9 9 12 2 7 9 7 9 0 9 2
8 13 15 9 2 13 15 9 2
11 10 9 9 2 9 7 9 13 10 9 2
33 0 9 13 7 13 9 9 16 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 12 3 0 3 13 1 0 0 9 2
10 9 10 9 13 11 11 2 13 11 2
19 10 9 15 3 3 3 13 2 9 7 9 3 10 9 12 9 3 13 2
4 0 9 13 9
20 3 1 9 1 0 0 7 0 9 13 0 9 1 0 9 0 0 0 9 2
29 1 10 9 13 0 3 9 9 9 11 11 2 15 3 1 0 9 7 9 0 11 1 9 0 9 13 1 9 2
16 0 0 1 0 9 13 0 9 1 9 0 9 2 13 11 2
14 13 3 9 1 9 11 1 9 7 9 3 16 11 2
21 0 9 15 13 1 9 2 16 11 13 10 0 9 7 0 9 15 1 15 13 2
18 11 1 15 13 2 16 11 13 0 9 2 7 3 1 9 10 9 2
14 3 1 0 9 3 16 0 0 9 13 9 2 9 2
9 3 15 7 13 13 10 0 9 2
3 9 1 9
27 9 9 1 0 0 9 13 1 11 7 9 0 9 2 0 9 16 11 11 2 11 11 2 9 11 11 2
14 9 1 15 13 7 0 0 0 9 11 2 11 11 2
9 13 7 13 10 9 2 13 11 2
16 0 9 14 13 1 9 0 9 2 1 9 0 9 1 0 2
20 1 10 9 13 0 9 0 9 11 11 2 0 1 0 9 16 0 0 9 2
16 15 9 13 9 2 9 3 13 3 10 9 2 3 9 9 2
19 13 15 1 15 2 16 13 9 9 2 16 15 9 15 13 1 9 9 2
21 13 15 13 1 10 9 2 14 3 1 12 1 12 12 9 2 3 0 9 12 2
3 9 1 9
2 11 2
16 1 0 9 9 13 1 9 9 9 11 11 11 12 2 12 2
19 0 9 13 9 0 9 11 13 15 1 0 11 11 3 14 1 9 11 2
33 1 9 12 2 12 7 9 14 12 9 15 15 13 0 2 7 9 11 11 13 2 2 1 11 4 13 3 0 9 16 1 11 2
24 13 15 7 15 2 16 9 13 13 0 9 12 2 12 2 1 0 9 13 12 9 7 13 2
6 3 15 13 10 9 2
20 1 9 15 13 1 0 0 9 2 13 7 13 13 3 3 1 0 9 2 2
5 9 13 1 12 2
6 1 11 14 12 0 9
2 11 2
23 0 9 4 13 13 1 0 9 0 11 14 12 9 7 3 14 12 2 3 15 3 13 2
53 2 9 11 3 9 1 15 9 13 2 13 7 3 3 0 2 16 1 9 13 10 9 9 2 16 1 9 0 9 1 11 4 13 0 9 11 2 7 15 13 1 15 3 0 2 2 13 11 11 2 9 11 2
6 16 13 9 7 13 9
28 2 11 12 2 12 2 12 2 9 9 1 10 9 13 3 2 7 13 4 0 9 2 16 3 15 15 13 2
40 9 13 12 9 2 16 4 15 3 2 13 2 16 2 2 13 2 13 15 13 2 7 1 0 9 3 13 13 2 16 4 9 3 13 1 9 0 0 9 2
31 1 10 9 13 13 9 9 1 9 10 7 15 9 2 16 4 15 7 13 1 9 2 15 4 13 1 9 9 2 2 2
31 4 2 14 13 9 2 15 4 13 0 1 12 9 2 13 10 0 9 2 16 4 15 9 13 10 9 1 0 9 2 2
23 16 9 3 2 13 1 15 2 16 9 9 9 13 1 9 0 2 7 15 15 13 13 2
19 1 9 1 9 2 13 2 14 3 15 2 15 14 4 13 10 9 13 2
8 9 7 9 2 7 3 1 11
12 11 13 1 15 3 16 9 9 7 0 9 2
28 3 15 3 13 13 12 1 0 0 9 2 9 11 11 1 9 0 9 10 9 9 7 9 2 0 1 9 2
9 3 9 7 11 3 1 11 13 2
15 1 0 0 9 15 15 7 9 0 11 13 1 10 9 2
25 1 10 9 7 13 3 13 0 9 11 11 2 10 9 15 1 0 11 13 1 9 0 9 9 2
22 9 9 7 9 2 0 9 2 2 0 0 0 9 2 13 3 0 9 0 0 9 2
25 9 1 0 0 9 1 1 10 9 9 7 9 13 3 3 2 3 7 13 3 3 7 3 3 2
13 0 9 15 3 13 0 7 0 0 9 9 9 2
35 9 11 11 1 15 1 9 13 0 9 0 9 1 0 9 11 11 2 9 9 2 0 0 9 7 0 9 13 1 0 9 0 0 9 2
19 9 13 1 9 0 9 0 9 1 9 11 11 7 13 0 9 11 9 2
15 0 9 13 3 0 0 9 0 2 9 7 0 0 9 2
8 12 13 0 9 0 0 9 2
16 3 13 1 9 9 2 0 0 9 2 7 9 0 0 9 2
36 3 0 13 7 0 0 9 2 3 0 0 9 0 11 7 11 1 0 11 2 1 9 1 9 9 2 11 2 11 2 9 2 11 11 2 2
16 3 1 0 9 0 11 3 13 3 0 9 1 0 0 9 2
28 1 15 13 9 9 11 2 1 15 0 0 9 11 11 2 11 13 0 9 7 10 0 9 1 9 9 9 2
19 1 0 9 0 9 13 0 0 0 9 9 11 2 9 2 11 11 2 2
36 3 16 1 15 0 0 9 9 11 2 9 9 2 7 9 1 2 0 9 2 15 13 13 12 1 0 9 9 2 15 13 0 7 0 9 2
7 9 1 0 9 1 0 9
11 1 0 9 11 13 0 9 1 9 11 2
20 1 0 9 13 13 2 16 15 3 13 7 0 0 9 2 14 0 0 11 2
7 0 9 13 3 3 0 2
36 0 0 9 13 11 9 1 9 9 2 7 10 9 13 1 9 12 1 9 0 9 0 9 2 13 1 15 3 0 9 1 9 11 1 11 2
16 0 9 9 2 11 2 13 12 9 2 7 1 15 0 9 2
14 11 3 13 9 12 9 11 11 7 3 15 13 9 2
16 1 9 15 13 3 9 7 1 0 0 9 0 13 9 9 2
14 9 9 13 9 2 11 11 2 9 9 9 7 9 2
13 13 7 9 0 9 2 13 0 7 3 15 13 2
18 9 9 9 2 9 2 11 11 13 9 7 9 7 1 11 3 13 2
17 9 13 0 0 9 1 9 11 2 11 2 11 1 11 1 11 2
29 9 1 11 13 9 2 3 0 9 2 11 9 7 1 9 0 9 0 13 1 9 0 9 9 10 9 1 9 2
15 1 9 15 13 0 0 9 2 15 13 0 0 0 9 2
19 3 15 1 9 13 0 0 9 0 9 2 9 0 2 1 10 11 11 2
12 0 0 0 9 11 13 0 9 0 9 11 2
27 9 7 9 13 9 0 0 9 7 9 3 13 3 1 11 2 1 0 0 11 2 1 11 7 1 11 2
8 9 13 0 9 9 0 11 2
16 9 13 9 1 9 7 0 15 3 13 7 1 10 9 13 2
25 9 1 0 0 0 0 9 13 9 9 2 1 15 15 3 13 2 7 1 11 0 1 15 13 2
13 1 0 9 0 1 11 4 13 1 9 7 9 2
22 0 9 1 10 9 13 9 2 16 1 11 4 13 0 9 0 11 2 0 9 2 2
25 1 9 13 1 11 0 9 0 0 9 2 0 0 9 2 7 0 0 0 9 1 15 3 13 2
61 0 9 0 11 13 3 9 0 0 9 1 11 9 2 9 2 11 11 2 2 0 2 0 9 1 9 0 2 7 9 0 9 9 2 9 2 11 11 1 11 1 11 2 0 9 1 11 2 2 7 3 0 9 9 11 11 2 15 13 2 2
26 9 13 9 11 0 1 0 9 2 7 3 13 9 2 16 13 1 15 9 0 9 10 9 1 15 2
23 1 9 13 0 9 9 2 9 2 11 11 7 9 13 0 11 7 1 11 7 1 11 2
21 0 2 0 0 9 13 1 9 3 3 13 1 0 9 0 0 9 1 12 9 2
16 3 10 9 13 9 0 9 2 7 3 13 7 13 9 13 2
17 1 11 7 1 15 13 0 9 2 15 1 9 1 9 3 13 2
23 3 13 1 15 2 16 4 13 13 10 9 2 15 13 0 9 7 9 9 1 0 11 2
7 0 9 9 1 11 1 11
15 16 4 9 13 13 3 0 9 2 13 9 1 15 9 0
25 1 9 11 2 9 2 2 12 2 12 2 2 13 9 1 9 9 12 1 0 9 0 1 9 2
10 10 9 13 7 13 7 1 0 9 2
21 1 9 0 9 11 2 11 13 12 2 9 9 9 1 3 0 9 2 11 2 2
24 1 9 11 2 11 2 3 13 10 0 9 1 0 11 2 13 0 0 9 0 7 0 9 2
19 1 9 1 9 11 11 13 0 13 0 0 9 7 13 0 0 0 9 2
23 9 9 12 4 13 1 9 1 11 7 0 9 1 9 2 11 2 11 7 11 2 11 2
19 0 9 9 12 2 15 13 1 0 0 9 2 13 7 0 13 1 9 2
18 1 9 1 0 9 0 9 13 9 9 9 14 1 3 0 0 9 2
37 3 2 1 9 1 9 0 9 7 0 9 1 9 9 7 0 9 2 1 9 12 13 0 9 1 9 9 12 1 9 1 0 9 12 1 9 2
48 0 9 3 1 9 12 13 1 0 0 9 0 9 1 11 2 15 13 1 9 9 9 11 7 10 0 9 3 0 7 1 10 9 13 9 13 3 7 3 2 10 9 9 7 10 9 13 2
34 7 16 9 9 0 9 9 12 1 0 9 3 13 2 9 9 9 3 13 0 9 9 9 12 0 3 2 1 0 0 9 0 9 2
34 9 10 9 15 9 3 13 1 9 1 9 9 2 12 2 12 9 2 1 9 9 7 9 2 15 1 0 9 9 9 9 3 13 2
51 0 9 9 9 12 3 13 0 9 3 1 10 9 2 16 0 9 0 9 9 7 0 0 9 2 15 13 13 0 9 0 1 9 12 2 13 0 9 9 1 0 9 1 9 9 2 12 2 12 9 2
30 1 9 0 9 0 9 9 12 4 1 9 12 2 12 13 0 9 9 7 1 0 9 2 15 3 13 0 9 9 2
34 9 13 2 16 0 9 0 1 0 9 9 12 4 1 10 0 9 4 13 1 0 9 11 2 0 9 0 11 7 0 9 0 9 2
42 9 11 2 11 1 9 0 9 3 13 9 0 0 2 0 0 9 1 9 12 2 15 1 9 13 1 0 9 7 0 9 0 9 1 9 3 0 7 0 0 9 2
30 1 9 1 9 0 1 9 13 0 0 9 9 9 0 9 0 9 11 2 11 2 15 13 0 9 1 0 0 9 2
99 9 2 0 1 9 12 0 9 1 11 2 11 7 11 2 13 1 15 2 16 9 1 9 1 11 2 0 0 9 1 0 9 9 2 4 13 1 0 9 2 1 9 0 9 9 12 4 3 13 0 9 14 1 0 9 7 1 0 9 4 13 0 9 2 16 0 9 1 11 13 1 11 2 3 13 1 0 7 0 9 12 2 9 7 9 11 2 11 13 9 0 9 11 2 11 1 2 11 2
31 16 9 1 10 9 2 16 3 13 2 13 0 2 9 9 13 0 9 11 2 11 7 11 9 9 12 3 3 0 9 2
27 9 1 3 0 9 2 11 2 13 0 9 0 9 1 3 0 7 13 9 7 9 2 15 9 9 13 2
45 0 9 11 2 11 4 13 0 0 9 9 1 9 2 3 9 9 9 9 9 7 0 9 13 3 3 1 0 1 0 0 9 2 1 0 9 0 9 9 2 11 1 2 11 2
19 0 9 9 12 13 3 0 7 3 13 9 1 9 3 0 9 0 11 2
25 10 3 0 0 9 13 9 14 1 0 9 2 7 7 1 0 9 0 9 1 0 9 9 12 2
37 11 15 13 1 9 9 0 2 0 0 9 2 16 9 16 9 0 7 0 9 2 3 16 4 13 13 3 0 9 2 13 9 1 15 9 0 2
39 13 15 1 0 7 15 7 3 0 9 2 1 0 7 0 9 3 7 3 0 0 0 9 2 15 13 1 15 0 2 16 15 13 3 0 2 0 9 2
26 13 4 9 1 12 10 9 2 16 4 10 0 9 4 3 13 9 3 0 9 2 16 13 1 11 2
59 11 15 7 13 1 9 9 9 7 13 9 9 7 9 11 2 16 4 1 9 0 9 11 2 11 3 13 10 0 9 1 9 3 0 0 9 7 13 3 0 0 7 0 9 2 15 13 0 9 0 9 14 15 2 7 3 0 9 2
16 0 9 1 11 13 2 16 9 0 0 9 11 9 9 13 2
4 0 9 1 11
2 11 2
25 9 0 9 1 0 11 13 1 9 0 0 9 1 9 1 12 9 0 16 1 0 9 0 9 2
10 9 0 9 9 13 1 9 12 9 2
19 0 9 13 9 9 1 11 2 3 13 1 9 9 1 12 9 1 12 2
13 1 11 13 9 0 9 1 12 9 1 12 9 2
24 1 15 1 11 9 13 1 12 9 1 12 9 7 1 11 15 13 1 12 9 1 12 9 2
27 0 9 1 9 0 9 15 1 11 13 9 11 1 12 9 9 2 7 16 13 1 12 9 1 9 12 2
13 9 0 9 9 9 11 13 1 12 5 1 12 2
19 10 9 1 9 13 1 12 1 12 9 11 7 1 12 1 12 9 11 2
11 1 12 0 9 1 12 9 13 9 11 2
20 9 11 13 1 12 1 12 9 7 9 0 9 15 13 1 12 1 12 9 2
21 0 0 9 9 13 11 2 1 10 9 13 1 9 9 9 1 12 9 1 12 2
12 9 11 1 9 3 13 1 12 1 12 9 2
7 11 1 9 1 11 14 13
2 11 2
37 0 11 3 13 2 16 13 1 0 9 1 9 10 0 9 2 15 13 1 0 9 2 16 15 4 11 13 2 16 4 13 0 9 1 0 11 2
20 9 0 9 9 1 9 0 9 11 13 2 16 9 9 10 9 13 15 13 2
46 11 2 0 11 7 11 13 0 9 2 15 4 13 11 1 0 9 1 11 7 11 2 0 3 1 9 1 11 2 13 0 0 9 9 1 15 2 1 15 11 13 10 0 0 9 2
6 0 9 15 13 1 9
2 11 2
28 1 0 0 9 15 9 13 9 1 10 9 1 0 9 7 9 9 13 0 9 9 3 1 9 0 0 9 2
40 1 9 4 1 0 9 2 3 15 0 0 9 1 9 13 1 9 9 1 0 16 0 0 9 1 11 2 16 9 13 2 13 13 0 9 1 0 0 9 2
11 0 9 13 13 0 9 7 13 9 9 2
24 16 7 13 0 2 13 15 15 0 9 9 2 16 9 13 2 13 0 9 11 0 11 11 2
17 3 1 9 13 9 0 9 10 0 0 9 1 12 5 12 9 2
23 1 0 0 9 12 9 15 9 13 1 9 1 9 1 9 0 9 1 9 9 9 11 2
6 11 13 1 0 0 9
2 11 2
16 0 9 13 0 9 9 1 0 9 2 15 13 9 9 9 2
28 11 13 2 16 4 15 1 9 2 15 15 13 9 1 9 2 4 3 13 3 2 1 9 1 9 9 9 2
20 9 1 9 4 1 0 9 13 13 3 9 2 10 9 13 12 9 0 9 2
23 11 13 1 10 9 9 10 9 2 15 15 1 15 13 3 0 2 7 0 7 0 9 2
5 0 9 1 9 12
2 11 2
13 0 0 9 4 3 13 1 9 1 9 0 9 2
8 9 15 13 0 9 11 11 2
24 10 9 13 1 10 9 3 0 2 0 9 7 13 1 15 2 16 4 3 13 15 0 9 2
28 9 4 1 11 13 12 9 9 2 1 0 9 4 7 3 13 3 1 12 9 2 15 13 9 1 0 9 2
39 9 13 2 16 9 9 11 12 7 12 2 1 10 9 9 13 2 13 9 1 0 0 9 0 9 2 16 4 9 13 3 2 16 15 13 0 0 9 2
26 9 4 13 13 0 0 9 1 0 9 7 1 0 9 7 13 9 12 9 2 9 9 7 9 3 2
3 9 13 9
18 1 12 3 9 1 0 9 13 0 0 9 1 0 9 9 0 9 2
5 9 13 15 0 2
17 0 9 13 7 0 9 2 1 11 7 11 7 13 3 1 9 2
12 9 9 9 13 3 9 3 1 9 0 9 2
18 3 1 9 13 7 9 3 0 2 16 15 13 0 9 7 0 9 2
5 9 13 1 9 2
31 9 11 3 13 9 9 1 0 0 7 0 9 7 3 9 0 9 0 0 9 1 9 10 9 7 0 9 0 9 9 2
24 9 2 15 13 3 3 1 9 2 13 0 13 3 2 1 10 9 7 0 9 13 3 0 2
13 11 3 3 13 1 9 0 1 0 2 0 9 2
17 1 15 13 15 3 0 9 9 2 15 13 3 9 1 10 9 2
16 11 13 1 9 1 0 9 3 0 9 10 2 0 9 2 2
35 13 3 0 2 16 1 10 9 15 13 9 10 9 11 1 0 9 2 0 9 13 15 1 15 7 3 0 9 13 15 13 1 10 9 2
24 0 9 0 9 2 3 9 13 9 2 15 13 9 3 3 13 3 1 9 2 16 13 15 2
18 1 15 3 4 9 9 13 13 9 11 2 7 14 15 2 1 9 2
18 13 9 0 9 1 9 2 16 10 9 13 1 9 2 15 13 13 2
17 3 2 9 1 9 7 9 10 9 4 13 13 12 1 9 9 2
13 0 9 2 15 13 9 13 10 9 2 13 9 2
26 0 9 3 13 2 16 10 9 13 9 2 1 15 15 13 13 9 2 7 16 15 13 13 7 13 2
7 9 0 9 9 13 13 2
16 0 9 3 13 13 7 1 9 9 0 9 3 1 9 9 2
25 0 9 4 7 13 13 1 9 1 9 0 9 9 2 1 15 2 13 15 2 13 15 1 9 2
9 0 9 4 13 13 9 1 9 2
17 3 1 12 9 13 9 11 9 1 0 9 9 9 7 0 9 2
21 16 11 7 3 13 9 13 9 9 1 15 2 13 15 0 9 13 1 0 9 2
7 9 0 9 9 13 9 3
5 14 2 0 9 2
2 11 2
25 1 9 0 9 0 9 11 11 2 11 2 11 2 13 0 0 9 9 0 9 9 9 9 11 2
12 1 10 9 13 14 0 13 9 9 0 9 2
24 1 15 13 7 9 0 9 9 2 16 4 9 1 3 0 9 13 9 13 9 0 9 9 2
14 10 9 4 15 1 0 9 13 3 9 9 9 11 2
7 13 4 15 7 9 9 2
12 9 0 9 11 11 11 13 0 9 1 0 2
19 2 13 2 14 13 9 0 9 2 13 13 0 9 9 13 2 2 13 2
29 9 1 9 11 13 1 0 9 2 2 3 13 2 16 13 9 1 9 13 3 9 2 15 13 1 0 9 2 2
30 1 9 11 11 11 13 13 9 9 1 15 2 16 4 1 9 2 3 9 13 0 15 13 2 13 9 1 9 9 2
19 9 11 11 2 11 2 13 2 16 1 9 9 9 13 3 0 13 3 2
12 13 7 9 2 3 4 13 4 3 13 9 2
16 15 2 16 4 9 13 15 13 9 1 9 9 2 15 13 2
17 3 9 11 11 9 15 13 1 2 9 9 9 1 9 9 2 2
30 9 0 9 11 11 2 11 2 13 2 16 16 4 15 13 13 0 9 2 3 4 13 1 0 9 1 10 0 9 2
14 1 9 12 14 1 15 9 9 1 9 9 3 13 2
21 2 13 2 16 11 16 0 9 13 3 13 2 16 4 13 10 9 2 2 13 2
33 11 11 2 11 2 13 1 9 0 9 1 0 9 2 3 7 1 15 2 16 4 1 9 2 3 9 13 13 2 9 13 9 2
4 13 9 9 9
5 14 2 0 9 2
4 9 9 15 13
2 11 2
20 9 9 0 0 0 9 4 0 9 13 1 9 9 7 3 3 13 9 11 2
8 1 11 15 3 13 9 9 2
26 1 0 9 0 9 9 13 1 0 9 1 9 9 9 1 9 0 9 9 1 0 9 1 0 9 2
11 3 13 4 9 13 1 0 9 9 11 2
25 15 13 0 9 9 7 9 11 2 0 9 11 2 0 11 2 11 2 11 7 0 7 0 9 2
19 0 9 7 13 0 13 11 9 1 9 9 7 3 9 13 0 9 9 2
19 7 9 9 0 9 13 2 16 0 9 7 9 9 15 13 0 9 9 2
15 0 9 1 11 11 13 0 9 9 1 12 9 9 3 2
19 9 1 9 13 13 12 9 9 2 16 0 9 4 13 12 9 15 9 2
9 0 9 13 1 0 9 0 9 9
8 11 11 3 1 9 9 1 11
5 9 13 9 1 9
14 1 3 0 9 9 15 13 13 0 9 1 12 9 2
21 0 2 15 13 9 9 2 7 0 2 9 9 1 0 9 2 15 10 9 13 2
20 7 3 13 0 9 1 0 9 1 9 7 0 9 13 0 0 9 12 9 2
3 3 0 2
12 16 13 9 2 13 15 1 9 3 0 9 2
10 16 4 15 3 13 2 13 13 3 2
21 1 0 9 3 13 3 3 9 9 2 7 0 12 0 9 1 12 7 12 9 2
11 3 3 13 1 9 3 12 0 9 3 2
14 15 13 0 9 2 7 9 2 0 15 9 3 9 2
22 3 1 10 0 9 15 10 0 9 13 12 9 7 13 3 0 13 0 9 0 9 2
10 13 1 9 9 7 9 13 9 9 2
8 1 9 9 13 12 9 3 2
16 9 13 15 3 3 13 9 2 15 13 1 9 1 0 9 2
23 13 3 1 10 9 0 7 0 9 2 16 4 3 0 7 0 9 9 4 3 3 13 2
21 13 0 9 2 7 0 9 2 3 9 2 9 7 9 13 1 0 9 9 9 2
8 13 7 13 9 9 13 9 2
16 13 9 9 7 15 13 0 15 13 1 15 0 9 16 0 2
16 0 9 13 1 9 9 2 7 1 15 0 0 9 10 9 2
3 0 0 9
2 9 2
35 3 16 1 0 0 9 0 0 9 10 9 1 15 2 12 2 13 7 1 10 9 11 1 0 9 3 0 9 2 0 1 0 0 9 2
35 0 0 9 11 11 4 3 13 2 16 4 13 9 1 9 0 9 7 15 2 13 13 14 3 7 9 2 15 13 13 1 9 1 9 2
30 1 10 9 11 3 13 2 7 0 9 13 16 9 1 9 0 0 9 2 15 13 1 2 0 2 9 1 0 9 2
23 0 0 9 3 13 3 0 9 9 11 11 2 15 9 15 0 9 13 1 9 14 0 2
15 0 9 2 0 9 7 3 0 9 13 0 9 0 9 2
59 0 7 0 9 2 15 13 0 9 1 0 9 2 1 13 1 0 9 2 0 9 7 9 1 11 2 9 1 9 2 3 13 0 2 0 0 9 2 0 10 0 9 0 9 2 15 13 2 14 16 15 13 2 14 7 14 13 2 2
21 0 7 3 3 0 9 13 9 0 9 2 0 13 9 1 0 9 7 0 9 2
15 11 11 2 11 11 2 9 11 2 0 0 0 9 2 2
6 9 12 2 12 9 2
4 13 2 11 2
7 9 1 11 2 11 11 2
23 1 9 0 9 11 11 1 9 11 11 11 13 1 9 9 0 9 1 9 9 1 11 2
8 11 13 1 11 1 9 9 2
20 1 9 9 1 11 3 13 2 16 11 3 13 9 1 9 11 7 0 9 11
7 9 1 9 11 13 0 9
5 14 2 0 9 2
4 11 2 11 2
26 11 11 7 11 11 1 0 9 7 11 0 1 0 9 0 9 13 3 0 9 9 1 9 11 11 2
14 1 0 9 9 13 3 9 12 7 9 1 0 9 2
24 2 13 2 16 4 9 9 13 10 0 9 7 3 13 0 9 1 11 11 2 2 13 11 2
12 2 9 11 13 1 0 9 9 0 9 2 2
26 0 0 9 11 11 7 11 11 3 13 2 16 4 3 13 1 9 9 9 1 11 1 9 11 11 2
15 1 11 13 9 9 11 11 16 0 1 9 0 9 13 2
46 11 11 2 12 2 4 3 1 9 13 1 0 9 9 1 0 9 1 9 9 0 9 1 11 11 11 7 0 0 9 11 11 2 15 1 9 1 9 12 13 2 9 7 9 2 2
17 11 4 1 9 13 7 13 1 9 2 16 15 3 13 0 9 2
16 1 9 15 13 13 9 7 15 1 15 3 13 0 0 9 2
16 11 13 9 0 9 11 11 2 15 1 9 12 13 1 9 2
11 11 2 11 3 13 3 11 1 9 11 2
5 15 13 1 9 2
28 15 13 10 9 1 15 2 16 9 0 9 4 13 4 13 9 2 7 0 9 9 11 1 0 7 0 9 2
15 11 11 2 9 0 2 0 2 11 2 2 9 9 13 2
14 3 1 0 9 13 9 3 7 13 9 4 13 3 2
13 7 9 1 15 2 10 9 13 13 2 13 0 2
5 9 13 0 9 2
7 1 9 14 1 0 9 2
21 3 13 1 15 9 2 15 13 14 9 2 7 3 15 2 15 13 7 0 9 2
11 9 9 0 9 13 1 15 0 3 0 2
9 16 9 13 1 10 9 2 13 2
11 11 11 2 9 11 2 9 13 1 0 2
19 16 9 13 9 2 13 2 16 1 11 13 9 3 7 3 15 4 13 2
10 1 10 9 13 2 13 0 3 13 2
18 9 1 9 9 13 3 7 13 0 7 0 9 2 15 13 1 9 2
11 11 11 2 9 9 2 13 1 0 9 2
7 12 9 13 1 11 3 2
8 15 4 3 3 13 1 9 2
16 0 9 4 13 2 16 4 13 14 15 2 15 15 13 15 2
19 1 0 9 4 15 13 3 9 2 15 4 15 2 15 13 2 3 13 2
30 11 11 2 9 11 2 1 0 9 13 16 0 9 2 7 7 9 3 13 0 9 3 2 3 9 3 13 3 3 2
26 9 15 9 2 3 0 7 0 2 1 0 9 0 0 9 1 11 7 3 1 11 3 13 7 13 2
29 13 0 9 9 7 13 14 1 10 9 7 9 2 7 7 9 7 9 1 0 2 16 3 0 2 0 2 9 2
4 9 1 9 12
8 0 0 9 13 9 0 1 9
2 11 2
26 12 0 9 13 1 9 9 0 1 0 9 1 11 1 9 9 7 1 15 3 1 12 0 0 9 2
14 13 3 9 0 0 9 11 2 15 3 3 13 9 2
17 13 12 1 0 9 0 9 1 9 2 0 0 9 2 9 2 2
21 11 1 0 9 13 3 0 0 7 3 0 9 1 9 9 1 0 7 0 11 2
13 13 3 7 1 0 9 13 9 2 9 7 9 2
13 1 12 9 3 13 13 16 0 9 2 7 9 2
20 9 13 13 1 0 0 9 1 0 9 2 3 16 1 0 0 0 9 9 2
34 11 1 0 13 2 16 4 0 9 13 3 2 12 9 1 9 2 7 3 13 1 0 9 0 9 2 0 1 9 0 9 9 0 2
6 11 1 11 3 1 9
2 11 2
13 0 9 11 11 4 3 1 9 13 13 0 9 2
27 2 9 1 0 9 11 2 15 3 7 3 13 15 0 9 2 3 13 2 2 13 0 9 11 11 11 2
29 2 13 4 0 2 15 1 0 9 9 9 11 1 0 9 3 13 1 9 9 11 11 1 0 9 2 2 13 2
10 9 0 9 13 11 3 1 0 9 2
8 9 4 13 3 1 12 9 2
4 0 13 1 9
2 11 2
21 0 1 11 13 3 0 9 1 0 9 2 15 3 13 9 0 9 0 0 11 2
15 9 10 9 13 0 0 0 9 7 13 1 15 9 9 2
8 13 1 15 3 0 9 9 2
15 16 13 2 9 13 0 9 0 9 9 0 9 1 0 2
10 13 0 9 1 9 9 0 0 9 2
14 9 7 9 9 4 0 9 1 0 13 0 9 9 2
4 11 13 12 9
5 14 2 0 9 2
2 11 2
25 0 9 1 0 9 12 9 0 0 9 9 13 3 11 1 0 9 2 11 2 1 9 9 11 2
11 13 15 3 1 11 0 9 9 7 9 2
28 0 9 9 11 11 11 13 2 16 0 9 1 10 9 2 12 9 9 2 4 13 1 9 7 9 9 9 2
17 0 12 9 4 13 1 9 0 9 7 12 9 1 9 0 9 2
18 1 9 9 2 3 1 9 9 0 9 11 2 4 13 12 9 9 2
1 3
14 0 9 13 1 9 12 9 1 0 9 12 9 9 2
24 1 0 9 1 0 9 11 13 11 11 2 12 2 1 10 0 9 0 9 1 0 9 1 11
20 11 2 3 2 13 9 2 7 1 9 15 1 9 12 2 12 1 11 13 11
6 9 1 11 1 0 9
2 11 2
15 9 0 9 1 9 1 11 13 0 1 9 0 0 9 2
29 0 9 9 1 11 13 2 16 9 1 0 11 4 13 1 11 12 2 9 12 7 1 12 9 13 12 12 9 2
6 9 1 11 13 9 9
3 0 11 2
25 9 0 0 9 13 9 2 16 4 1 9 11 13 9 2 1 15 4 9 1 9 13 9 9 2
16 9 0 9 11 11 13 2 16 12 7 12 9 4 13 0 2
23 1 11 13 10 9 13 3 0 9 7 3 13 13 1 0 9 2 15 13 1 9 9 2
14 9 15 13 9 0 9 1 0 9 0 1 9 9 2
28 7 16 9 3 13 0 9 2 1 9 0 2 0 9 2 3 9 2 13 0 9 9 0 9 1 10 9 2
3 10 9 9
13 13 15 15 3 9 9 0 1 9 13 3 0 2
37 11 11 2 11 12 2 9 12 2 13 2 9 2 0 9 2 0 9 9 1 9 2 0 14 2 9 2 7 3 2 9 2 1 10 0 9 2
56 1 9 2 3 1 11 2 7 2 10 9 13 11 2 15 3 16 9 0 0 9 13 2 10 0 2 9 11 1 2 0 2 0 2 0 11 1 9 7 3 15 1 15 2 3 1 12 9 2 13 0 9 1 0 9 2
33 13 15 0 9 0 9 2 1 0 11 7 0 11 2 2 1 0 9 9 2 7 1 15 0 9 2 1 9 0 1 0 9 2
26 0 0 9 13 0 2 0 9 7 2 16 13 0 2 16 13 9 0 9 7 0 9 1 0 9 2
13 13 3 0 2 10 9 7 0 9 13 1 9 2
16 3 4 13 1 11 13 0 2 0 7 0 9 16 1 11 2
18 9 7 3 13 2 13 15 9 2 7 15 15 3 13 2 0 2 2
24 9 1 10 9 13 1 0 9 7 1 9 2 13 15 7 3 1 0 9 0 9 7 9 2
20 2 7 3 14 13 0 2 3 2 0 0 9 2 13 7 3 1 9 2 2
29 3 13 9 2 0 3 2 3 9 3 13 9 2 3 14 0 9 2 3 3 7 3 3 2 0 2 7 0 2
14 0 2 0 11 7 3 2 0 11 13 3 3 9 2
23 0 9 13 7 13 10 0 0 9 3 2 3 0 9 2 0 9 15 13 1 9 9 2
20 1 9 0 9 15 3 13 9 12 9 2 3 3 2 3 15 13 11 11 2
19 12 10 9 9 13 0 9 2 12 1 10 2 15 13 10 9 7 9 2
14 13 15 14 3 3 3 14 7 2 16 13 3 3 2
13 0 9 13 2 9 15 13 2 7 7 9 13 2
5 13 15 7 15 2
10 14 9 13 2 7 16 0 16 0 2
26 2 4 13 2 16 13 3 9 2 7 3 0 2 16 10 2 15 13 13 9 2 7 10 0 2 2
14 9 15 3 3 13 7 13 1 9 2 7 1 9 2
12 13 2 7 15 1 0 9 3 13 1 9 2
34 13 15 1 15 3 3 0 9 2 7 16 0 9 9 3 1 9 0 0 9 13 1 9 2 13 15 9 3 0 9 9 0 9 2
19 0 9 0 9 7 9 2 3 1 0 0 9 2 3 13 0 9 9 2
20 1 9 9 13 0 9 2 0 7 0 1 15 2 14 9 2 7 3 9 2
10 0 9 3 13 7 1 9 1 9 2
13 0 9 3 2 3 0 2 9 13 7 3 13 2
41 13 15 15 1 9 2 7 0 7 0 2 2 3 7 0 0 9 2 0 1 0 9 7 14 1 0 9 9 7 9 7 1 9 2 1 0 0 9 3 13 2
17 7 1 10 9 13 2 3 1 9 1 10 10 9 2 3 3 2
19 0 9 11 4 15 2 3 3 13 2 13 0 0 9 7 9 11 0 2
21 13 1 15 15 2 7 3 2 3 1 9 12 2 13 10 9 1 9 3 0 2
19 13 4 15 7 13 3 7 3 9 2 0 9 10 9 13 1 15 9 2
12 13 15 0 9 1 9 7 3 15 15 13 2
10 13 1 15 15 3 10 0 0 9 2
19 3 3 14 2 9 1 9 13 3 2 16 1 15 3 13 9 0 9 2
22 13 3 2 3 7 13 3 0 2 13 1 10 0 9 7 15 13 9 10 0 9 2
17 7 15 3 1 2 9 2 9 13 3 7 3 0 9 10 9 2
22 3 16 1 9 9 2 1 0 11 7 0 11 2 15 3 13 7 3 3 13 4 2
36 13 15 10 9 2 13 2 3 2 15 2 15 13 3 7 14 15 2 15 15 13 11 2 11 7 0 7 15 4 15 13 13 10 0 9 2
23 16 15 15 3 9 9 9 0 13 13 0 2 13 1 15 2 0 9 2 3 0 9 2
10 9 1 9 11 11 1 0 2 0 9
2 11 2
30 13 15 13 0 9 2 13 0 9 9 2 11 11 1 9 2 3 13 9 0 2 0 9 0 1 9 9 11 11 2
35 1 9 2 3 13 1 10 9 9 0 9 15 0 9 2 0 9 13 2 16 1 10 9 15 9 11 13 3 0 9 0 2 0 9 2
31 9 13 0 9 0 2 0 9 3 1 9 11 1 0 9 13 1 9 9 11 2 11 0 9 9 11 1 9 11 11 2
35 1 9 2 16 15 15 13 0 0 9 2 13 2 16 1 9 0 9 13 3 1 9 0 0 2 0 9 7 9 3 0 7 0 9 2
26 9 9 11 11 11 1 9 11 2 11 13 2 16 9 0 1 9 13 3 0 1 0 2 0 9 2
21 1 10 9 7 13 13 0 9 7 13 15 0 2 3 9 1 0 9 7 9 2
8 1 11 15 13 11 2 9 0
3 11 11 2
21 3 13 9 9 11 11 9 13 9 1 9 1 9 9 11 2 9 1 10 9 2
20 3 13 0 9 0 9 11 11 2 9 13 3 9 2 15 1 11 11 13 2
10 1 9 13 9 0 9 9 1 9 2
28 3 3 9 13 9 1 0 9 3 1 9 9 2 7 1 9 13 1 9 9 2 15 13 9 1 9 9 2
26 3 1 9 13 9 13 9 0 9 2 1 15 15 1 9 9 11 2 9 3 13 3 12 9 9 2
5 12 9 11 4 13
2 11 2
27 1 12 9 1 0 9 1 0 9 12 0 9 0 11 1 9 12 13 0 9 9 0 9 3 0 9 2
9 13 1 15 3 9 9 11 11 2
28 1 15 12 9 15 9 11 11 11 13 1 0 9 1 9 2 16 4 13 0 9 0 9 1 9 10 9 2
16 1 12 9 4 13 9 0 9 7 12 9 4 3 3 13 2
6 1 9 15 14 13 13
55 9 1 0 9 2 15 13 1 12 12 9 2 9 3 0 1 9 0 7 0 0 9 2 3 1 0 9 1 0 0 9 1 12 9 2 7 10 9 13 1 9 1 0 9 9 2 12 2 15 3 13 1 0 9 2
25 2 9 13 3 0 13 15 2 1 9 14 1 3 0 9 2 2 13 9 9 0 9 11 0 2
22 2 9 9 7 3 13 13 1 15 2 16 9 13 14 1 9 2 7 13 7 3 2
27 9 13 0 13 15 9 1 12 9 2 0 9 2 15 13 1 9 0 9 2 7 13 1 0 9 2 2
11 7 1 9 14 13 2 16 9 13 9 2
21 0 9 0 1 9 13 9 7 9 2 16 4 3 13 2 9 15 7 13 13 2
22 1 0 15 13 13 2 16 3 16 1 9 13 9 1 9 2 1 9 2 1 9 2
16 3 13 13 7 9 0 9 2 10 0 9 13 9 1 9 2
11 9 2 3 1 0 9 2 13 0 9 2
18 9 15 3 3 13 16 0 2 13 1 0 9 7 13 0 1 9 2
15 9 1 12 9 15 9 13 1 12 9 2 9 1 12 2
8 7 15 15 3 1 9 13 2
15 9 15 13 1 15 2 16 11 13 1 9 9 3 0 2
11 3 7 1 9 13 0 9 7 0 9 2
12 9 0 9 13 7 9 2 3 9 0 9 2
26 1 9 9 3 13 7 0 12 9 0 0 9 0 9 11 2 11 2 0 1 11 1 12 0 9 2
15 1 9 15 7 9 13 3 1 9 2 1 12 9 9 2
12 3 16 3 0 0 7 0 9 13 9 9 2
18 0 9 3 13 13 7 15 2 15 1 9 1 0 9 13 7 13 2
4 11 0 9 11
4 11 13 1 9
23 0 9 0 9 13 0 0 9 11 11 11 2 15 13 12 9 7 1 12 15 13 9 2
23 0 9 13 13 1 9 1 0 9 9 2 16 15 13 9 1 0 9 1 0 11 11 2
17 3 0 9 3 13 0 0 9 2 3 15 9 13 1 0 9 2
9 3 7 10 9 9 1 9 13 2
22 9 0 15 13 15 2 16 11 13 1 15 0 0 9 2 2 1 9 13 3 3 2
14 3 15 13 3 7 2 16 1 15 13 3 13 2 2
26 2 13 15 15 7 13 4 9 2 16 15 9 13 0 9 2 2 13 3 11 2 15 13 0 9 2
15 2 1 9 4 13 1 9 10 9 2 16 13 1 9 2
18 1 11 3 13 3 12 12 9 2 7 16 1 15 13 0 9 2 2
19 11 13 1 0 9 7 10 9 0 9 2 0 13 1 0 9 7 9 2
24 13 13 7 1 10 0 9 2 15 13 2 9 2 2 2 13 4 1 11 13 3 0 9 2
27 1 9 9 15 13 1 9 2 7 16 4 1 11 13 7 1 9 2 13 2 16 13 13 3 3 2 2
31 0 2 15 11 13 2 13 9 9 0 9 1 10 9 2 2 13 2 3 15 15 15 13 2 15 3 13 0 9 13 2
10 1 11 15 7 1 9 13 1 9 2
12 9 13 9 1 11 7 15 15 1 11 2 2
5 0 9 13 1 11
16 3 9 9 11 3 13 1 11 9 13 9 9 0 0 9 2
16 1 0 9 3 13 11 11 2 11 11 7 0 0 9 11 2
49 0 9 0 9 2 15 13 9 7 0 9 2 13 9 11 1 9 9 12 0 9 1 0 9 11 1 9 7 1 9 0 0 9 2 1 15 4 4 1 0 9 13 9 9 7 0 9 11 2
13 9 15 3 13 2 16 0 0 9 13 9 9 2
22 1 11 13 7 0 9 9 11 11 7 13 15 13 10 3 0 9 1 9 0 9 2
20 9 15 13 7 11 13 0 9 9 7 9 0 9 2 3 13 15 3 2 2
20 1 0 9 11 9 2 11 13 15 7 9 3 2 15 11 13 1 10 9 2
4 11 2 0 9
20 9 0 0 9 9 1 11 13 9 9 2 1 15 15 0 9 3 3 13 2
10 1 9 0 9 13 1 9 11 9 2
14 1 9 13 9 2 15 13 3 1 0 9 1 9 2
14 1 0 9 4 13 10 0 9 2 13 1 0 9 2
14 1 9 13 0 9 2 15 13 1 9 1 10 9 2
6 10 9 13 3 0 2
25 13 7 1 11 9 2 15 4 15 13 2 3 3 2 3 3 2 16 10 9 13 1 9 9 2
26 3 1 9 0 1 9 9 1 9 9 2 3 0 9 11 11 13 12 12 9 7 3 4 15 13 2
19 0 9 1 9 2 9 9 2 13 9 2 1 0 9 13 9 1 9 2
21 1 11 7 1 0 9 0 9 13 9 9 2 9 9 2 9 9 7 0 9 2
10 1 9 3 13 9 9 1 0 9 2
14 9 9 9 13 2 16 4 15 13 9 1 0 9 2
9 1 12 1 9 9 4 13 9 2
5 13 14 0 9 2
13 9 13 9 2 16 4 9 13 1 9 1 9 2
22 0 9 0 9 0 9 13 2 13 7 7 15 2 15 4 1 11 11 0 13 9 2
17 12 1 9 13 2 2 1 9 0 1 15 13 0 11 11 2 2
24 13 2 14 12 2 13 3 7 0 9 2 1 2 0 2 9 13 11 10 9 12 2 9 2
16 15 9 2 15 9 1 0 9 2 15 13 1 9 0 9 2
14 9 14 13 13 0 9 7 15 13 1 9 0 9 2
7 7 9 13 3 0 13 2
37 9 1 0 9 15 1 11 13 9 9 2 0 9 2 1 0 9 2 11 2 11 2 11 7 11 2 16 4 15 13 13 1 0 9 1 9 2
16 9 13 15 9 11 2 16 4 15 13 9 7 13 10 9 2
21 0 9 2 0 1 9 2 13 0 0 9 2 0 9 15 9 13 1 10 9 2
6 9 15 13 1 9 2
11 3 1 15 13 9 7 13 15 1 9 2
7 9 13 1 9 7 15 2
20 0 9 2 15 13 1 9 2 15 13 2 2 3 13 13 1 9 12 2 2
13 9 1 15 2 2 7 15 13 9 2 2 2 2
22 0 9 9 11 11 1 11 13 2 16 9 1 9 0 9 13 0 14 1 9 9 2
3 13 9 2
20 0 9 11 11 13 2 16 9 13 0 13 14 1 9 9 1 9 0 9 2
6 7 15 13 3 9 2
6 9 11 3 9 13 2
19 13 2 16 13 13 1 15 2 16 4 9 13 10 9 2 9 0 9 2
6 7 15 13 7 9 2
17 9 13 3 2 3 13 0 9 15 0 9 0 1 9 0 9 2
11 15 13 10 0 9 2 15 13 0 13 2
9 3 7 13 1 9 10 11 0 2
5 11 13 11 7 11
2 11 2
40 0 9 11 11 13 1 9 1 0 9 9 11 11 9 0 9 2 16 4 0 0 9 3 13 11 7 11 1 0 9 9 1 9 0 9 0 1 10 9 2
9 13 15 3 3 9 9 11 11 2
34 11 2 13 0 13 9 2 15 15 13 2 16 0 9 2 16 4 13 0 9 9 0 10 0 7 0 9 1 11 2 2 13 11 2
16 13 2 16 0 9 13 9 11 2 15 7 13 13 13 15 2
9 11 11 13 1 11 1 9 1 11
5 14 2 0 9 2
2 11 2
32 0 9 15 1 0 9 13 0 9 2 16 9 1 11 13 15 13 7 16 13 3 1 15 2 3 7 3 13 9 0 9 2
19 1 0 9 0 0 9 1 11 15 13 9 0 9 11 11 2 11 2 2
15 1 9 9 13 12 9 1 0 9 1 9 0 9 11 2
20 1 11 13 0 11 3 13 2 16 2 0 1 9 13 1 10 0 9 2 2
25 9 9 14 1 9 13 2 16 0 9 2 15 15 13 12 0 9 2 13 9 9 9 1 9 2
58 1 0 9 0 9 9 11 11 7 9 9 9 9 11 11 1 9 9 2 15 3 2 13 9 9 2 11 2 11 2 11 2 11 2 7 9 10 9 1 11 2 12 2 9 12 2 11 13 2 16 13 1 9 1 0 0 9 2
23 2 9 9 7 0 9 12 9 1 10 9 3 13 9 2 15 4 15 15 13 3 13 2
13 13 15 14 9 13 9 3 0 9 2 2 13 2
28 11 13 2 16 0 9 0 9 11 11 9 11 2 1 15 13 0 9 1 9 9 2 4 13 14 12 9 2
40 2 15 4 15 1 11 3 15 13 2 16 4 13 2 16 13 0 9 1 10 9 2 7 13 4 15 7 10 9 10 9 9 0 7 3 0 2 2 13 2
23 11 13 3 0 2 16 11 7 1 9 0 9 13 0 9 7 13 12 1 0 0 9 2
21 2 13 2 16 15 15 1 11 7 1 10 9 13 13 0 9 2 2 13 11 2
27 9 0 7 0 9 11 11 2 11 2 13 2 16 3 1 9 13 13 9 11 1 0 9 9 1 9 2
15 9 9 12 15 14 9 13 7 3 4 3 13 0 9 2
21 2 15 13 1 15 0 2 13 13 2 16 13 9 0 1 0 2 2 13 11 2
1 3
16 0 9 1 9 1 0 9 1 11 13 9 1 3 0 9 2
14 1 0 0 9 4 1 0 9 9 13 7 9 0 2
21 1 9 13 10 9 0 7 13 15 2 16 15 13 13 0 0 0 9 1 9 2
16 9 1 9 0 9 1 9 13 11 11 1 11 1 0 11 2
21 9 0 9 0 9 2 12 9 0 9 1 11 2 15 13 1 12 9 12 12 2
3 11 13 11
5 14 2 0 9 2
3 0 11 2
22 16 0 9 9 9 13 9 0 0 9 1 0 2 3 13 1 9 9 9 11 11 2
40 2 0 9 13 1 0 2 10 0 9 1 9 13 13 2 2 13 9 9 11 11 1 9 0 9 11 2 15 15 13 1 9 1 0 11 1 0 2 11 2
32 11 13 2 16 0 9 13 0 9 9 1 9 9 9 2 3 1 9 0 9 7 9 0 9 1 9 0 9 7 0 9 2
22 9 4 3 13 3 3 13 0 9 9 7 0 9 9 7 13 9 9 1 0 9 2
27 1 11 13 9 9 13 2 3 7 3 2 3 15 4 13 9 1 0 9 9 7 0 9 7 9 2 2
20 11 13 2 16 9 15 13 7 9 9 0 9 2 15 13 9 9 11 9 2
21 1 9 11 13 2 16 9 13 2 9 3 3 0 2 7 16 9 10 9 13 2
8 3 1 0 9 11 1 9 12
4 0 9 1 9
7 0 9 15 13 7 0 9
20 7 0 9 0 9 13 9 13 9 2 7 7 13 10 9 1 3 0 9 2
13 13 1 15 7 9 1 0 9 2 11 7 11 2
41 3 15 9 13 1 11 2 11 7 11 2 7 9 15 13 7 1 3 0 9 2 15 13 3 11 7 13 15 2 16 7 0 9 3 3 13 15 2 15 13 2
13 10 9 7 13 0 2 1 0 3 11 7 11 2
13 1 9 11 3 1 9 12 13 7 12 0 9 2
21 3 13 15 3 12 7 1 0 9 12 0 9 0 1 10 9 15 13 12 9 2
13 1 11 13 9 12 9 2 12 1 9 0 9 2
15 0 9 9 1 12 9 13 12 5 2 7 9 13 15 2
31 3 0 13 7 0 0 9 9 2 15 13 0 0 9 2 15 13 1 9 0 9 1 11 2 15 13 0 10 0 9 2
16 1 9 9 13 9 1 11 2 7 9 0 13 13 1 9 2
17 9 1 9 1 0 9 1 0 0 9 13 9 13 1 0 9 2
8 7 13 1 9 0 0 9 2
14 15 7 13 13 2 16 4 15 1 9 0 9 13 2
6 0 9 13 4 13 2
28 9 11 3 3 13 15 2 16 1 10 9 13 9 11 11 2 7 15 9 2 15 13 1 0 9 10 9 2
8 0 9 15 13 7 0 11 2
12 11 7 11 13 3 9 2 9 15 15 13 2
25 10 9 15 13 15 2 16 13 9 1 9 0 9 3 0 11 1 11 7 11 11 2 9 2 2
18 12 9 9 0 1 12 9 1 0 9 13 1 12 0 0 0 9 2
11 0 9 13 10 9 7 9 1 0 9 2
10 1 9 1 9 15 7 13 13 9 2
7 3 4 15 15 13 13 2
6 9 9 13 3 1 9
15 2 13 9 2 3 15 13 12 2 2 13 9 11 11 11
21 9 1 0 9 0 0 9 13 1 11 1 11 12 1 0 9 9 1 0 9 2
18 1 9 2 15 0 9 1 9 11 13 2 7 0 0 9 3 13 2
25 16 9 9 13 2 9 11 11 3 13 9 1 0 9 7 3 15 1 15 13 12 9 1 9 2
26 1 9 9 2 15 1 0 12 9 3 13 2 7 3 15 13 13 9 2 4 15 13 1 9 11 2
42 2 1 1 0 9 2 15 1 9 13 2 4 13 13 13 0 9 2 7 7 9 9 10 9 2 16 4 13 13 2 14 2 13 13 7 13 9 13 1 0 9 2
10 1 9 13 0 9 2 11 1 11 2
34 1 9 4 13 13 11 2 7 1 1 9 9 2 15 13 2 13 11 7 1 12 9 13 2 7 7 1 11 13 0 0 9 2 2
15 11 11 13 16 0 9 2 7 3 0 9 13 1 9 2
16 1 9 1 0 9 1 9 13 2 1 0 9 15 3 13 2
12 2 13 2 1 9 13 2 14 13 0 9 2
13 1 9 3 13 7 0 9 2 3 3 13 13 2
15 11 13 9 0 9 2 1 9 15 13 0 9 0 9 2
12 10 9 2 9 2 9 7 9 13 0 2 2
5 13 15 3 3 2
3 2 13 2
10 7 13 9 2 16 15 15 13 9 2
18 3 4 1 9 13 13 0 10 9 2 7 15 1 10 9 13 13 2
14 9 13 2 15 13 0 13 7 15 1 15 13 13 2
22 13 2 16 13 9 2 7 13 2 16 11 13 0 0 9 2 7 13 1 15 13 2
18 3 16 15 13 7 1 9 13 0 9 2 3 13 11 0 15 13 2
6 7 9 15 13 2 2
17 1 9 15 3 13 1 10 9 1 9 9 11 2 1 15 13 2
15 2 13 1 10 9 2 7 3 15 13 1 9 1 9 2
11 13 15 2 16 13 0 9 1 9 9 2
15 13 15 13 9 0 9 1 9 7 13 15 1 0 9 2
13 13 1 10 9 15 13 2 3 15 3 13 2 2
18 13 1 9 9 11 2 11 2 9 2 15 1 15 13 9 1 11 2
8 2 13 4 2 16 4 13 2
13 16 4 13 1 0 9 2 3 4 13 0 9 2
20 13 11 2 11 2 9 2 11 7 11 7 9 3 13 2 13 15 10 9 2
18 12 15 3 13 7 15 13 13 9 2 15 13 1 3 0 9 0 2
14 0 13 2 16 4 1 0 9 13 1 9 13 9 2
20 1 9 13 12 12 9 1 11 2 7 13 9 2 3 15 13 14 12 2 2
11 13 2 16 3 10 9 1 9 9 13 2
32 2 9 13 3 2 7 13 15 13 1 15 2 16 15 13 13 2 16 1 0 9 13 9 2 15 1 15 13 0 0 9 2
15 15 15 7 13 2 0 9 4 13 2 16 4 13 11 2
30 1 9 1 0 9 4 13 1 9 2 16 4 13 1 9 7 13 4 13 3 9 2 15 1 0 9 13 0 9 2
33 3 15 13 2 16 4 1 0 9 13 13 12 9 2 15 4 1 9 13 2 11 1 0 11 7 11 2 15 3 13 1 11 2
15 11 13 3 11 12 9 7 15 4 13 12 2 12 2 2
23 15 15 13 2 16 1 3 0 9 2 15 13 11 1 11 2 13 9 9 1 9 9 2
8 2 0 9 13 1 0 9 2
13 15 13 2 16 15 13 15 1 9 13 2 2 2
6 13 2 13 14 13 2
10 0 9 15 9 13 13 7 7 13 2
7 13 9 2 3 15 13 2
18 16 15 13 9 2 15 13 10 0 9 2 3 15 3 15 4 13 2
34 1 11 4 13 1 9 11 11 2 9 13 0 9 2 16 4 15 3 9 13 2 13 15 13 2 7 9 1 9 9 13 13 2 2
6 15 13 1 0 9 2
26 2 3 2 16 15 1 9 13 1 0 9 2 3 0 9 13 1 9 2 16 15 13 9 1 9 2
9 9 13 9 7 13 15 13 13 2
16 9 15 9 3 13 2 0 15 13 7 13 4 15 3 13 2
8 15 15 13 2 9 13 0 2
11 11 2 11 7 11 4 13 1 10 9 2
13 1 0 9 15 13 2 15 1 9 13 16 9 2
27 9 0 9 13 1 15 0 2 7 9 1 0 9 13 3 0 7 15 15 13 2 16 13 14 0 9 2
9 1 9 4 13 1 0 9 3 2
19 1 0 9 4 13 7 9 2 15 13 14 1 9 2 7 1 0 9 2
12 13 2 16 15 4 13 9 2 15 13 9 2
12 9 7 13 0 2 13 2 16 4 3 13 2
11 13 0 2 16 13 0 9 1 15 2 2
3 9 13 3
2 11 2
22 9 0 9 15 13 1 9 1 0 9 1 12 5 7 0 9 13 14 1 12 5 2
11 13 15 1 9 0 0 9 1 0 9 2
11 0 0 9 9 13 9 9 3 0 9 2
21 3 1 0 7 0 9 9 13 1 12 5 2 9 7 9 9 13 1 12 5 2
10 3 13 0 7 0 9 1 0 9 2
23 9 0 9 9 1 0 9 3 13 2 16 9 13 1 12 9 7 0 9 1 12 5 2
11 9 0 9 13 1 0 9 1 12 5 2
4 9 4 13 13
2 11 2
25 1 0 9 9 1 0 9 13 9 0 0 9 11 11 3 2 9 0 9 1 15 7 9 11 2
27 9 1 0 0 9 9 11 4 13 1 9 9 1 12 5 7 1 9 4 9 13 1 0 9 0 9 2
22 9 0 9 4 13 9 1 9 7 4 15 13 13 9 1 9 9 3 1 9 9 2
17 1 9 3 0 1 0 9 3 10 0 9 13 7 1 0 9 2
34 2 13 2 16 15 9 2 15 13 1 9 1 9 1 9 0 9 2 4 13 2 2 13 1 9 1 9 9 0 0 9 11 11 2
5 9 1 12 2 9
2 11 2
20 0 9 15 1 15 0 0 9 1 15 4 13 1 12 2 9 0 1 9 2
14 0 9 4 13 3 2 16 4 4 9 13 9 9 2
24 1 0 9 1 9 1 0 9 7 1 9 1 9 11 15 13 1 10 0 9 0 9 11 2
3 11 13 13
2 11 2
9 9 11 11 1 0 9 15 13 2
25 9 0 9 7 9 11 2 15 3 12 9 13 9 9 2 3 13 10 9 1 0 9 1 11 2
10 2 13 4 3 0 2 2 13 3 2
16 0 9 9 13 11 1 9 1 11 11 2 12 2 9 2 2
23 7 1 10 9 7 9 3 13 1 0 0 9 1 9 12 2 16 9 13 1 0 9 2
5 9 9 1 0 9
37 3 9 9 0 1 0 9 2 15 1 9 9 2 9 13 3 2 12 9 2 2 9 11 12 2 13 9 2 9 7 9 1 0 15 0 9 2
37 9 11 11 2 12 2 1 15 1 0 0 9 13 9 9 1 12 0 9 10 9 2 1 11 2 11 7 1 11 1 11 1 0 2 0 9 2
32 9 0 9 13 11 11 2 1 15 13 9 9 2 9 2 0 9 2 9 11 2 9 1 9 11 7 13 1 9 0 9 2
22 2 9 1 9 2 3 4 13 2 13 3 0 2 16 4 13 2 2 13 11 11 2
10 2 1 11 15 0 9 14 3 13 2
17 3 4 15 3 13 2 16 0 9 3 13 1 9 1 0 9 2
32 1 11 13 9 0 0 9 1 11 2 7 3 13 3 0 2 16 1 11 15 9 1 0 9 13 0 7 1 0 15 13 2
9 9 15 3 3 13 13 0 9 2
18 3 9 13 15 13 2 16 1 11 13 10 9 9 2 2 13 9 2
18 9 0 1 0 9 1 11 13 15 3 0 7 13 15 7 10 9 2
20 2 16 13 3 1 3 0 9 2 3 15 15 1 15 13 13 7 0 9 2
15 15 3 3 3 13 2 3 0 13 10 9 1 0 9 2
21 9 9 15 3 13 2 16 13 2 14 0 9 2 15 0 15 3 13 1 0 2
15 7 1 9 4 15 3 13 2 16 3 3 15 13 2 2
38 1 9 11 2 11 13 11 11 3 9 9 1 12 9 2 1 11 0 2 9 2 9 9 9 9 1 9 11 11 7 1 0 9 9 9 11 11 2
28 1 2 0 2 9 9 13 13 9 1 9 9 2 9 7 9 0 9 2 1 15 13 1 9 9 9 0 2
27 2 9 13 13 1 9 9 2 15 1 9 13 12 9 2 13 15 1 10 9 3 3 7 3 9 13 2
16 1 9 1 10 9 15 13 7 0 9 9 2 2 13 11 2
21 0 9 15 13 9 13 7 1 0 0 9 2 1 9 2 9 2 1 0 9 2
23 2 13 15 1 15 13 1 9 2 3 15 10 9 3 3 2 9 0 9 2 13 13 2
16 3 4 13 13 2 15 1 10 9 13 9 2 2 13 9 2
15 1 0 11 13 11 0 9 1 9 7 9 10 0 9 2
25 2 12 13 11 11 2 0 13 11 2 0 11 2 16 15 0 15 13 1 11 7 1 0 9 2
9 9 10 9 4 13 13 0 9 2
29 1 15 15 3 3 13 7 13 1 9 1 9 2 15 15 0 1 9 13 2 7 9 2 1 15 1 9 13 2
26 9 13 9 1 9 0 2 0 7 0 7 9 2 15 13 1 9 9 3 2 2 13 9 11 11 2
7 11 11 4 13 1 9 9
9 11 11 13 1 9 0 0 9 9
17 14 0 0 9 0 0 9 0 9 13 1 9 1 9 0 9 2
22 1 0 9 13 0 9 7 11 11 2 12 2 1 0 9 11 11 1 11 1 11 2
9 0 0 9 13 1 9 0 9 2
28 1 9 11 11 1 9 12 13 1 0 9 9 9 0 9 2 0 9 9 2 10 9 15 13 7 11 11 2
35 9 3 1 0 9 2 3 13 3 11 9 2 11 11 7 11 11 2 1 10 9 13 0 9 7 13 9 2 15 13 9 1 0 9 2
20 10 0 9 1 9 9 1 0 9 1 9 15 3 13 7 9 1 0 9 2
25 9 13 12 7 12 9 3 2 3 1 9 1 9 7 9 1 0 9 2 1 9 9 0 2 2
8 1 0 9 13 0 9 9 2
10 10 0 9 13 9 7 0 0 9 2
23 1 0 9 13 1 9 9 11 11 2 1 0 9 13 3 9 9 1 0 9 0 9 2
2 0 9
19 0 9 15 3 13 1 9 9 7 3 1 15 7 0 9 1 10 9 2
17 1 0 9 4 15 13 13 2 16 10 9 14 13 3 0 9 2
30 16 4 7 0 9 13 3 9 0 7 16 4 3 13 9 9 9 2 13 0 2 16 4 4 13 9 15 0 9 2
6 3 7 15 9 13 2
13 9 0 9 1 9 13 14 0 9 9 0 9 2
24 9 9 1 9 1 9 13 3 0 7 2 16 13 7 13 9 2 7 7 2 16 13 9 2
21 1 9 0 9 15 1 9 13 11 2 11 2 15 3 13 9 1 0 0 9 2
10 1 9 9 3 10 9 13 1 9 2
19 12 1 9 10 0 9 13 3 9 3 0 9 2 15 15 1 11 13 2
15 11 2 11 4 3 13 1 9 7 1 10 9 0 9 2
30 13 7 13 4 2 16 9 0 13 0 9 3 0 7 3 0 2 16 0 9 3 13 13 3 1 3 15 0 9 2
21 3 4 13 2 16 3 13 1 0 9 2 7 3 1 1 9 0 9 0 9 2
23 16 15 3 1 9 0 0 9 13 7 0 0 9 2 13 15 0 9 1 0 9 9 2
35 7 16 2 16 4 10 9 1 9 1 0 9 1 9 3 12 9 3 1 15 13 1 9 1 10 9 2 13 3 3 13 9 9 0 2
15 1 10 0 9 2 15 9 13 2 4 0 13 3 15 2
22 1 0 9 13 1 9 9 7 9 3 9 0 9 2 15 3 13 9 9 7 9 2
22 0 9 0 9 9 9 9 1 9 1 9 13 1 10 9 0 9 1 9 0 9 2
12 13 0 0 9 7 13 13 9 0 9 9 2
11 13 7 1 0 9 9 1 9 1 9 2
13 0 9 13 3 1 9 12 13 9 1 0 9 2
7 13 1 15 3 10 9 2
23 9 9 4 13 1 0 9 7 13 0 9 9 2 7 7 13 1 0 9 1 9 9 2
10 9 13 9 0 9 2 15 9 13 2
14 0 0 9 13 0 14 1 10 9 2 15 9 13 2
21 13 3 0 2 16 4 9 2 1 10 13 9 9 2 1 15 13 1 9 3 2
25 13 7 3 0 13 12 9 2 1 15 9 13 2 16 4 10 9 1 9 13 3 14 1 9 2
10 9 9 13 1 9 9 1 9 9 2
16 9 9 1 0 9 7 13 9 7 1 9 2 7 1 9 2
24 1 9 12 15 13 13 2 16 0 9 9 0 9 13 7 9 9 13 1 0 9 0 9 2
28 1 10 10 9 15 3 13 2 16 0 9 9 1 0 9 13 9 1 9 12 2 12 9 1 9 0 9 2
17 9 13 7 1 15 2 16 1 10 9 15 9 0 9 3 13 2
29 16 15 1 15 3 13 3 9 0 9 9 2 15 4 13 9 9 13 2 13 10 9 0 3 1 3 0 9 2
10 1 9 1 0 9 13 1 9 9 2
29 9 10 9 7 13 13 3 10 9 0 9 2 15 13 0 7 0 9 9 2 7 2 9 1 9 14 3 0 2
11 7 13 1 0 13 1 10 9 0 9 2
15 13 3 3 13 9 9 9 9 2 15 13 13 3 0 2
10 1 15 10 9 13 0 1 9 13 2
20 0 9 13 3 0 9 7 13 1 15 13 16 1 0 9 12 9 1 0 2
17 13 15 13 0 9 0 9 2 7 14 3 2 13 2 14 0 2
11 13 2 14 2 13 15 0 9 1 9 2
4 0 9 13 9
2 11 2
39 3 3 12 9 0 9 15 1 0 9 13 1 0 9 9 9 2 9 11 11 11 2 1 15 13 1 9 13 0 9 11 11 11 2 3 1 0 9 2
23 0 9 13 0 9 1 3 0 7 13 2 16 13 1 9 9 0 13 10 9 0 9 2
25 9 9 13 7 10 0 9 2 15 13 11 2 16 4 13 1 10 9 2 7 15 13 0 9 2
15 9 9 11 7 9 10 9 13 7 0 9 13 1 0 2
3 3 0 9
1 9
10 9 15 1 9 3 13 1 0 9 2
10 3 15 13 1 9 1 9 9 9 2
15 1 9 1 11 15 7 13 2 16 15 3 13 0 9 2
4 13 10 9 2
32 16 9 1 9 3 13 2 9 13 3 3 1 9 7 0 9 2 0 9 15 3 3 13 1 9 7 9 9 15 3 13 2
22 9 13 2 16 16 9 9 13 7 0 9 15 13 2 9 9 15 13 7 3 13 2
23 1 15 9 3 13 13 0 3 1 9 7 13 3 0 9 9 2 3 9 1 9 9 2
24 9 13 3 13 7 9 13 9 2 13 0 9 9 7 13 3 10 9 1 9 9 0 9 2
15 16 13 15 2 9 13 13 1 0 2 13 0 2 9 2
11 13 7 15 2 15 4 15 3 13 9 2
12 1 10 9 13 13 2 16 13 3 1 15 2
7 1 0 9 13 15 9 2
20 1 0 9 13 0 13 2 16 0 9 0 9 13 3 3 9 16 0 9 2
27 3 3 0 0 9 1 0 9 1 9 2 9 12 9 1 9 9 1 0 9 0 9 7 9 1 9 2
6 15 1 15 15 13 2
28 15 13 13 15 2 15 15 15 13 2 16 13 3 1 0 2 7 0 9 9 2 1 10 9 3 13 3 2
11 9 11 13 9 3 9 3 1 0 9 2
10 9 2 3 15 13 13 2 13 0 2
24 9 13 2 16 13 0 13 0 9 9 2 13 9 9 7 3 13 2 15 1 15 4 13 2
23 10 9 7 13 9 3 3 3 7 13 15 2 16 3 4 15 13 13 1 9 15 13 2
11 9 13 1 9 1 0 9 0 9 11 2
15 15 15 7 13 7 3 11 15 2 16 10 9 1 9 2
11 13 1 15 2 16 15 9 13 3 13 2
11 9 0 9 11 7 9 15 1 9 9 13
1 9
2 11 2
27 1 9 0 9 2 15 9 9 13 9 1 9 0 9 2 11 2 2 13 3 0 9 11 2 12 5 2
13 11 4 1 10 9 13 12 5 7 11 12 5 2
11 11 2 11 7 11 4 13 3 12 5 2
10 0 9 4 13 3 16 12 5 0 2
9 9 11 13 0 9 0 9 11 2
17 0 0 9 0 9 2 9 0 9 2 9 2 2 10 9 13 2
9 1 9 9 13 9 11 0 9 2
21 11 13 3 0 9 9 11 7 0 9 9 11 2 11 12 2 12 2 12 2 2
22 1 11 13 11 1 0 9 12 9 2 11 0 9 1 9 0 9 1 10 9 13 2
25 0 9 9 13 0 9 9 0 9 2 1 12 5 1 9 0 9 1 12 5 1 9 0 2 2
15 1 9 11 15 11 13 3 0 9 2 1 12 5 2 2
12 0 9 12 9 15 3 13 7 1 9 11 2
21 1 11 4 10 9 13 1 9 12 5 7 1 11 1 15 3 16 12 5 0 2
33 1 9 13 7 0 9 2 3 11 13 1 9 7 9 0 9 1 0 9 11 2 2 11 2 16 0 9 13 9 12 7 0 2
2 0 9
2 11 2
10 3 1 12 12 9 13 0 9 11 2
14 10 0 9 0 9 1 9 9 4 13 1 0 9 2
36 1 10 9 2 9 0 9 11 11 11 13 1 0 0 9 2 15 4 15 13 1 9 13 9 9 2 7 7 9 7 9 1 9 0 9 2
13 1 9 1 15 13 9 2 7 7 9 7 9 2
30 2 13 4 13 1 10 9 1 0 9 2 2 13 9 2 11 7 13 2 16 0 9 0 9 11 13 3 12 9 2
14 3 13 0 9 2 1 9 12 2 2 0 13 0 2
13 1 11 2 11 7 11 13 0 9 1 10 9 2
25 1 0 9 13 0 9 11 3 12 9 2 1 15 13 3 9 11 2 7 7 9 0 9 11 2
19 2 13 2 16 4 4 16 0 3 13 16 0 9 2 7 3 7 9 2
18 13 1 0 9 2 7 3 1 9 1 9 2 2 13 11 2 11 2
14 1 10 9 15 0 9 13 10 9 1 9 3 13 2
1 3
25 0 0 9 15 13 13 1 0 9 2 9 7 0 2 15 13 0 9 0 2 9 7 0 9 2
19 13 7 1 9 1 0 9 13 3 3 12 7 12 0 9 1 0 9 2
10 0 10 9 13 9 3 9 0 9 2
15 1 10 0 9 12 0 9 13 12 9 7 13 12 9 2
5 0 9 13 1 9
9 9 3 13 9 1 0 7 0 9
3 0 11 2
20 0 9 13 1 0 9 0 9 2 0 2 2 13 3 10 0 9 11 11 2
9 1 15 15 9 13 13 0 9 2
19 3 4 13 1 10 9 1 0 7 0 9 2 15 4 9 13 0 9 2
15 15 9 13 14 0 9 2 7 3 13 15 1 0 9 2
9 0 9 1 9 0 9 13 9 2
8 9 9 3 13 9 0 9 2
12 9 3 13 0 9 1 9 1 9 7 9 2
17 3 13 9 1 9 7 13 9 2 16 13 13 1 9 15 9 2
9 1 0 13 11 2 11 9 0 2
13 7 13 0 9 9 13 9 7 9 9 0 9 2
13 1 10 9 15 3 13 13 0 9 9 7 9 2
17 9 3 13 13 3 12 9 9 0 9 1 3 16 0 9 9 2
26 0 9 4 11 13 1 12 9 1 11 11 2 9 2 9 2 0 2 2 15 13 12 9 9 11 2
19 15 3 3 13 3 12 12 9 0 9 1 9 2 1 12 3 16 3 2
24 1 9 13 3 0 9 0 9 0 9 3 0 1 12 9 2 15 15 13 14 12 9 9 2
19 1 10 12 9 9 13 1 9 9 1 0 9 11 1 0 11 1 11 2
6 0 11 13 3 0 9
2 11 2
29 0 0 9 11 0 0 2 12 1 9 9 11 2 13 1 0 9 9 12 9 9 2 9 2 2 12 9 9 2
14 9 13 0 16 0 12 9 9 9 1 3 0 9 2
24 9 9 7 9 9 7 13 3 13 10 9 1 0 9 2 13 1 9 11 1 9 0 9 2
20 1 9 12 13 9 9 11 1 12 9 9 1 9 9 12 1 12 9 9 2
11 0 9 1 11 13 15 1 9 9 13 2
15 9 1 9 1 0 9 0 11 13 4 13 1 9 9 2
19 9 1 11 7 13 2 16 1 1 9 9 9 4 13 4 9 3 13 2
7 9 11 2 11 1 9 9
2 11 2
29 0 9 11 11 13 0 9 1 9 0 0 9 2 15 13 13 9 1 9 7 9 9 1 9 1 9 7 9 2
19 13 15 3 1 9 9 2 15 13 9 1 9 0 9 9 9 7 9 2
36 0 9 9 4 1 0 9 13 0 0 9 1 0 9 2 7 9 13 0 2 9 9 1 9 2 15 4 13 9 1 0 9 7 0 9 2
11 9 0 9 13 10 9 9 0 9 13 2
17 9 15 13 1 9 0 9 2 15 13 1 9 11 13 9 3 2
4 11 1 9 13
11 1 11 13 1 0 9 0 9 7 12 9
2 11 2
23 1 0 9 1 11 13 0 9 7 12 9 2 0 9 0 9 7 0 9 0 9 13 2
18 9 9 11 11 11 11 13 9 1 0 9 3 0 2 13 0 9 2
28 13 4 15 1 15 13 7 0 9 2 3 11 11 7 11 7 9 11 2 1 15 11 3 13 1 0 9 2
25 2 1 9 9 4 13 1 11 7 11 2 7 11 15 13 9 7 1 0 9 9 13 12 9 2
14 3 15 13 7 11 2 7 15 15 1 0 9 13 2
37 1 12 9 1 9 13 9 11 2 11 7 11 2 2 13 11 7 13 3 3 3 2 16 13 13 0 9 0 9 2 15 4 13 1 0 9 2
19 2 13 4 1 0 9 2 1 15 7 13 13 0 9 9 7 9 2 2
13 1 9 2 15 1 11 13 2 13 9 3 11 2
35 2 9 13 7 0 11 2 11 4 3 13 7 1 11 4 1 0 9 13 2 16 13 2 7 4 1 15 3 13 2 2 13 11 11 2
7 2 9 1 0 9 13 2
23 3 1 0 9 4 9 13 2 16 1 15 13 15 13 2 15 15 13 7 13 1 15 2
22 15 13 13 9 2 2 13 0 9 7 13 2 16 0 9 13 1 0 9 1 9 2
25 0 9 11 2 12 2 9 2 12 9 2 12 9 2 12 9 2 9 12 2 12 2 12 9 2
38 13 2 11 2 11 2 12 9 1 11 2 2 11 2 11 2 2 11 2 11 2 13 1 11 2 2 11 2 11 2 12 1 9 9 1 11 2 2
42 13 2 11 2 11 2 2 11 2 11 11 2 2 2 11 2 11 2 2 11 2 9 9 1 11 2 2 11 2 11 2 2 2 11 2 9 9 1 11 11 2 2
3 11 13 9
10 11 13 1 9 9 2 12 9 9 2
2 11 2
21 11 2 0 9 0 0 9 0 0 9 2 13 10 0 9 11 1 9 0 9 2
33 11 2 15 13 0 0 9 1 9 12 2 15 1 15 13 0 9 7 13 0 9 1 9 2 16 15 13 10 9 1 0 9 2
19 2 13 12 9 0 9 2 2 13 3 11 11 2 0 9 0 0 9 2
23 0 9 4 0 12 9 13 0 9 1 9 1 9 2 9 2 9 2 9 7 0 9 2
10 2 1 10 0 9 13 11 3 0 2
25 9 10 9 13 13 1 0 11 0 0 9 2 15 4 15 13 14 1 9 12 2 2 13 11 2
26 2 11 13 1 0 9 10 9 7 13 3 0 9 2 16 9 13 0 1 12 9 2 2 13 11 2
11 1 0 9 12 1 11 13 11 12 9 2
18 1 9 0 9 15 13 0 9 2 12 0 9 2 1 15 12 0 2
27 1 9 0 9 13 11 9 1 10 9 9 7 9 2 1 9 9 2 0 9 2 0 9 7 0 9 2
3 3 0 11
1 9
23 9 2 0 9 11 15 9 0 9 11 2 11 2 11 13 1 0 9 1 9 0 9 2
22 1 9 0 9 9 13 0 9 9 2 9 11 11 7 9 11 11 1 9 11 11 2
20 0 0 9 0 1 0 9 2 3 7 9 2 13 9 9 1 3 0 9 2
7 9 15 13 1 0 9 2
23 9 3 3 13 1 9 10 9 2 7 13 3 9 0 9 2 10 0 9 1 0 9 2
19 3 13 7 0 9 2 3 13 9 0 9 1 0 9 7 0 0 9 2
18 3 15 7 9 13 1 9 0 9 0 0 9 2 3 0 0 9 2
20 9 4 13 0 9 0 9 2 15 15 3 13 7 13 2 0 13 0 9 2
13 7 9 10 9 3 13 7 13 14 1 0 9 2
15 0 9 9 13 0 9 1 0 9 7 0 9 10 9 2
18 9 13 13 16 1 0 9 9 2 7 1 3 0 7 0 9 9 2
13 9 13 0 0 9 2 13 15 1 0 9 9 2
23 9 15 13 1 9 0 9 11 2 11 7 11 2 16 11 7 11 3 13 13 0 9 2
47 0 9 2 0 1 9 9 2 13 9 9 7 9 2 3 9 11 7 11 2 1 0 9 2 1 0 9 15 13 1 0 9 0 2 1 9 13 0 9 7 14 9 15 3 13 9 2
24 0 9 2 1 15 15 7 13 9 0 2 13 9 3 0 9 1 9 11 2 11 11 2 2
13 1 15 13 3 9 0 0 9 1 11 3 0 2
33 0 11 13 3 3 0 2 1 0 0 9 2 7 3 1 15 13 0 9 2 13 9 2 13 11 2 11 11 2 7 13 15 2
15 10 0 9 7 13 15 9 7 13 14 1 9 0 9 2
37 1 10 9 13 0 7 0 9 0 9 2 3 15 1 9 13 0 9 0 9 2 1 0 9 15 13 9 2 13 9 7 0 11 13 0 9 2
35 0 0 9 13 9 11 7 11 2 11 11 2 2 15 3 3 13 0 9 2 9 1 9 2 2 7 1 9 15 13 3 0 9 9 2
30 11 11 15 7 1 9 11 13 13 0 9 2 13 15 1 14 0 9 2 13 15 0 9 2 15 13 1 0 9 2
12 3 13 15 7 15 7 3 3 13 0 9 2
17 10 0 9 13 3 0 9 7 9 1 11 2 15 3 7 13 2
2 11 11
15 9 11 2 11 2 11 1 11 2 11 2 11 2 11 2
8 9 12 2 7 12 2 9 2
3 9 0 9
1 9
2 9 2
24 1 0 9 1 9 13 0 9 11 11 2 9 2 7 11 11 2 9 2 9 3 0 9 2
33 0 9 13 3 1 9 1 10 0 0 0 9 7 10 0 9 2 0 9 1 9 2 0 2 3 0 9 15 13 9 0 11 2
34 11 11 13 10 9 9 0 0 9 2 0 0 2 0 9 2 7 13 15 16 9 0 9 2 9 7 9 2 0 0 7 0 9 2
24 11 11 2 15 13 9 0 0 9 1 0 9 1 11 2 15 3 13 9 16 9 0 9 2
27 10 0 7 0 2 0 7 0 9 13 12 9 1 0 9 2 13 9 9 9 3 2 3 15 13 15 2
39 13 1 15 9 9 1 9 2 9 1 9 7 9 2 15 9 7 9 15 3 13 16 9 1 9 2 3 0 0 0 9 1 0 9 1 11 11 2 2
23 0 9 9 13 9 3 0 0 9 2 1 0 15 12 13 1 9 2 15 15 13 9 2
17 9 11 11 13 0 9 2 15 13 0 9 7 9 1 0 9 2
45 10 0 9 11 2 0 9 2 0 9 2 9 2 15 1 9 13 2 0 9 2 0 9 1 9 2 9 2 2 7 0 0 0 9 2 0 0 0 9 2 13 10 0 9 2
7 11 9 15 13 7 13 2
12 11 9 7 0 0 0 9 13 3 1 15 2
12 9 9 7 9 9 13 1 9 9 1 9 2
29 9 9 4 13 13 9 11 11 0 1 9 1 9 2 2 13 0 9 9 2 13 9 2 3 9 0 3 2 2
6 1 11 13 9 1 9
2 11 2
25 1 0 9 1 0 11 13 3 1 0 0 9 9 1 9 2 15 13 0 1 9 9 11 11 2
17 11 13 16 0 9 1 0 9 7 13 0 16 0 9 0 9 2
29 9 15 3 2 3 16 9 2 13 9 0 9 7 2 9 15 9 2 11 11 2 1 10 9 4 9 11 13 2
29 11 2 15 13 1 9 12 1 0 9 1 9 0 0 9 2 13 9 1 0 9 2 15 15 13 1 0 9 2
3 3 9 13
1 9
53 1 9 1 9 11 15 9 10 0 9 2 3 11 7 11 2 13 13 2 16 13 3 14 0 2 16 4 9 7 9 0 0 9 13 9 7 0 9 1 0 9 2 16 9 0 1 9 13 0 7 13 15 2
29 3 3 11 7 11 13 0 9 1 15 2 16 4 1 9 0 9 2 3 7 9 2 0 9 16 9 13 9 2
12 13 4 3 9 1 9 9 7 3 1 9 2
12 3 4 13 0 9 13 1 0 9 1 9 2
15 13 4 9 3 0 9 13 2 16 4 13 1 0 9 2
6 0 9 13 3 9 2
29 9 3 1 9 0 9 11 11 13 2 7 16 4 15 0 9 3 13 2 13 15 1 9 9 1 9 0 9 2
21 0 9 15 13 15 2 3 3 2 16 1 15 1 0 9 15 1 0 9 13 2
10 3 0 0 9 3 13 13 1 9 2
8 1 0 9 0 9 13 13 2
33 1 11 1 9 12 9 1 9 0 0 9 0 0 9 13 0 9 7 1 9 0 0 9 0 0 0 9 15 13 0 0 9 2
10 0 9 1 11 13 10 9 9 9 2
28 13 3 0 2 16 4 15 9 2 15 3 1 9 12 1 9 13 0 9 1 9 12 2 13 13 10 9 2
12 0 9 10 9 13 7 13 1 15 0 9 2
10 9 1 11 11 2 11 2 2 9 9
23 9 9 9 0 11 1 9 9 7 10 9 4 1 9 1 0 9 1 9 13 1 0 2
14 3 13 1 15 0 9 1 3 0 9 1 9 11 2
21 1 12 9 13 3 9 1 9 2 1 9 11 13 12 9 2 1 11 14 12 2
13 0 9 13 3 1 9 10 0 9 0 0 9 2
16 10 9 15 15 13 7 0 9 2 1 9 2 0 9 3 2
9 15 15 3 3 13 1 9 12 2
20 1 1 9 9 7 0 9 9 13 1 0 9 3 0 9 13 1 9 11 2
20 7 7 15 3 3 13 1 15 2 16 9 13 1 9 7 16 13 3 13 2
19 9 11 3 13 10 9 2 3 15 3 3 13 7 13 15 9 10 9 2
17 9 2 16 13 3 15 3 1 9 9 2 13 0 9 10 9 2
26 1 9 0 9 15 3 3 1 9 11 13 9 9 7 9 2 15 13 1 9 1 10 9 13 3 2
14 0 9 13 7 10 9 13 3 0 9 1 0 9 2
1 3
36 2 0 9 1 9 2 13 9 9 2 15 1 9 7 9 3 13 0 9 11 12 2 9 9 11 7 9 1 9 7 9 0 7 0 9 2
33 9 2 0 9 2 7 0 0 9 13 1 11 9 1 11 3 1 12 2 9 2 3 1 9 9 9 11 11 12 2 1 11 2
8 10 9 13 9 11 1 9 2
24 15 13 2 16 0 9 10 9 13 2 7 15 13 1 9 1 0 9 9 1 9 7 9 2
24 9 9 12 0 1 9 12 2 2 12 2 9 1 0 9 4 13 13 1 9 0 0 9 2
16 1 3 16 12 9 9 3 13 9 9 9 2 9 7 9 2
10 4 3 3 13 0 2 0 0 9 2
9 0 9 13 10 9 1 0 9 2
23 3 9 3 1 12 2 9 13 1 9 12 0 7 12 0 9 1 11 2 11 7 11 2
7 0 9 1 11 1 11 2
2 11 2
19 0 9 15 13 9 2 16 0 9 13 1 0 9 7 9 0 0 9 2
11 0 9 3 1 9 3 13 9 7 9 2
13 10 9 13 1 3 0 9 1 0 9 7 9 2
7 1 9 9 10 9 13 2
19 13 15 15 13 15 0 2 3 16 15 1 15 10 9 13 13 0 9 2
19 0 9 9 11 11 13 3 3 1 12 1 9 11 1 9 1 0 9 2
14 1 11 13 10 9 11 11 2 12 9 13 1 9 2
22 11 13 0 9 1 0 9 2 15 13 0 9 1 9 0 7 0 9 1 0 9 11
5 9 13 7 13 9
2 11 2
28 9 13 9 1 9 9 7 9 2 15 13 9 1 9 11 13 2 10 9 13 13 1 9 9 1 10 9 2
20 1 10 0 9 11 11 15 3 13 2 16 9 13 10 9 1 9 0 9 2
17 1 0 9 15 9 9 13 9 11 2 15 13 1 0 9 11 2
18 13 3 3 12 9 7 9 13 1 10 9 9 12 9 9 0 9 2
27 9 9 13 14 13 9 2 7 3 15 13 7 1 0 9 2 9 7 0 9 0 1 9 1 10 9 2
9 1 9 15 13 1 9 9 12 2
11 1 9 0 9 15 13 0 9 0 9 2
28 1 9 13 9 1 9 9 0 15 2 16 1 0 9 9 9 13 3 3 3 9 7 13 15 9 0 9 2
12 0 9 13 7 0 9 0 9 1 9 9 2
34 0 9 10 9 9 13 7 15 15 13 2 16 1 0 0 9 15 13 9 1 0 7 0 9 2 15 3 13 0 9 7 9 9 2
12 9 1 9 0 9 13 1 0 9 0 9 2
17 1 9 0 9 1 9 9 13 9 13 0 9 1 9 0 9 2
12 9 3 13 9 1 9 2 0 15 10 9 2
13 3 13 9 13 14 0 9 9 9 1 9 9 2
17 9 10 9 13 3 0 0 9 2 7 16 4 13 1 12 9 2
9 11 4 3 13 9 1 12 9 9
2 11 2
21 1 9 9 9 0 0 9 4 13 11 2 13 2 9 9 3 1 12 9 9 2
8 13 15 3 9 9 11 11 2
15 1 9 1 12 9 4 13 0 9 3 13 1 9 9 2
13 0 9 1 0 12 9 9 13 1 0 9 9 2
20 3 2 16 9 13 0 9 7 13 0 9 2 4 10 9 13 1 0 9 2
11 9 15 13 0 9 2 0 9 7 9 2
27 9 7 13 0 0 9 1 9 9 1 12 2 9 1 9 2 15 3 3 14 12 9 7 12 9 13 2
14 1 15 4 13 11 1 0 9 9 1 12 9 9 2
23 2 1 10 9 4 13 9 2 3 1 15 4 9 3 13 10 0 9 2 2 13 11 2
28 7 2 7 3 1 9 9 7 9 2 4 9 13 7 1 9 12 2 3 13 10 0 9 2 3 0 9 2
4 0 9 1 9
2 11 2
17 9 13 1 12 7 9 9 9 7 3 3 0 9 13 10 9 2
22 9 9 0 0 9 1 0 11 13 1 0 9 1 15 2 16 15 10 9 13 13 2
13 9 0 9 0 0 9 11 11 15 13 1 0 2
9 13 2 16 9 1 10 13 9 2
16 1 9 13 1 15 0 13 9 2 1 16 4 15 3 13 2
9 9 4 3 1 9 0 9 13 2
18 9 15 1 11 11 13 1 0 9 3 3 2 16 13 1 0 9 2
24 13 3 3 16 0 0 9 15 0 0 9 2 9 2 0 9 2 0 9 7 0 9 2 2
17 9 1 9 13 1 9 11 0 9 2 7 9 9 1 10 9 2
9 16 15 13 2 13 9 9 9 2
36 1 0 9 0 9 13 1 9 7 15 2 16 9 9 13 13 3 1 9 0 9 1 9 1 9 3 1 9 2 3 15 9 1 9 13 2
27 2 9 13 7 0 13 1 10 9 2 16 14 0 9 1 9 2 0 9 7 0 9 2 2 13 11 2
23 16 1 9 13 1 11 0 9 9 12 9 2 13 15 10 9 2 16 15 1 15 13 2
20 1 11 15 3 13 1 9 2 15 3 13 9 15 9 2 15 15 13 9 2
13 2 1 15 4 10 9 14 13 2 2 13 11 2
16 13 2 16 13 9 13 3 0 9 2 13 15 3 10 9 2
15 15 15 1 9 13 13 0 9 2 13 0 7 0 9 2
5 11 2 9 9 9
6 9 11 15 13 9 11
2 11 2
15 7 0 9 1 0 11 13 0 11 1 9 13 0 9 2
10 2 13 2 16 13 15 1 10 9 2
30 9 9 15 1 10 9 3 1 9 3 13 2 3 15 9 13 14 1 9 2 2 13 9 1 11 0 9 11 11 2
34 3 0 9 1 0 9 13 1 11 9 1 0 9 2 13 1 15 12 9 2 2 0 9 1 11 2 7 3 3 0 9 13 11 2
28 2 1 9 13 1 15 9 2 7 16 3 4 13 9 9 2 2 13 9 11 11 0 9 9 1 12 9 2
19 9 11 15 13 0 9 11 7 3 11 2 15 13 0 0 9 12 9 2
18 2 0 9 13 1 0 9 11 2 16 3 13 9 2 2 13 11 2
16 1 0 0 9 13 1 9 11 1 11 2 15 13 0 9 2
24 3 0 9 11 13 0 9 3 1 12 2 9 2 16 9 15 13 1 9 14 1 9 9 2
18 9 13 3 12 9 0 1 9 2 1 15 0 9 11 13 9 11 2
15 1 15 13 9 11 0 9 2 16 13 9 9 9 12 2
9 1 9 13 11 3 12 9 9 2
17 12 12 1 10 9 13 9 11 2 0 3 11 11 7 11 11 2
11 11 13 11 3 3 12 9 1 0 9 2
13 0 9 13 11 2 9 2 2 0 11 7 11 2
27 1 9 0 9 11 13 9 3 13 2 12 9 1 0 9 2 12 9 1 0 7 12 9 1 0 2 2
15 2 13 10 9 7 9 2 15 1 0 9 1 9 13 2
16 13 13 0 9 1 9 9 2 2 13 0 9 9 11 11 2
26 0 9 11 2 12 2 9 2 12 9 2 12 9 2 12 9 2 9 2 12 2 12 2 12 9 2
16 13 2 11 2 11 2 11 2 11 2 13 1 9 9 2 2
28 13 2 9 2 11 2 2 11 2 9 1 11 2 2 11 2 9 1 11 2 2 11 2 9 1 11 2 2
7 1 9 1 0 9 1 9
2 11 2
19 1 9 0 9 1 9 7 1 9 13 1 0 9 0 9 0 9 11 2
28 16 15 4 9 13 15 9 2 9 7 9 2 13 3 0 9 0 9 11 11 2 11 2 15 15 13 3 2
12 3 0 9 0 9 3 9 13 1 9 0 2
31 0 9 4 13 7 9 11 2 11 2 12 2 9 2 2 11 2 11 2 12 2 2 7 11 2 11 2 12 2 2 2
10 9 1 0 0 9 15 13 1 9 2
9 2 13 4 0 3 1 12 9 2
13 15 4 3 13 2 2 13 9 0 9 11 11 2
20 1 9 2 15 4 13 1 0 11 2 13 3 1 10 9 1 9 0 9 2
4 0 9 13 2
15 0 0 9 13 1 12 2 9 2 15 13 9 9 11 2
18 16 4 1 15 13 11 2 13 4 0 0 9 1 9 11 2 11 2
18 1 9 13 3 0 9 1 9 11 2 11 1 9 12 2 9 3 2
24 16 0 9 13 1 0 9 1 0 2 1 9 1 9 9 13 12 9 3 2 12 2 9 2
23 2 13 4 2 16 4 0 1 0 9 13 3 0 0 9 2 2 13 9 9 11 11 2
38 0 9 11 11 13 1 0 9 9 16 0 9 1 9 11 2 1 15 13 13 9 14 9 0 9 2 3 9 0 2 15 1 9 13 9 0 9 2
23 2 1 9 11 13 9 2 16 9 13 0 2 2 13 11 1 9 0 9 9 9 12 2
12 1 9 1 0 0 9 15 13 9 0 9 2
16 2 9 13 3 1 0 9 3 9 2 16 9 13 10 9 2
14 0 9 13 13 0 9 2 2 13 9 11 11 0 2
6 9 1 0 0 9 2
20 12 2 9 2 12 2 12 2 2 2 11 2 11 1 1 12 14 1 12 2
3 9 0 9
9 0 11 1 9 0 9 7 0 9
21 0 0 9 11 2 15 13 1 9 9 9 2 3 3 1 0 13 0 0 9 2
7 13 7 1 9 3 0 2
14 9 0 9 0 2 3 0 2 9 13 3 3 0 2
19 3 13 0 9 0 2 11 2 11 2 11 2 2 7 7 0 9 0 2
34 13 15 9 0 9 2 9 0 0 9 11 11 2 11 2 11 11 2 11 1 11 2 3 9 0 0 9 9 11 11 7 11 11 2
18 11 3 13 2 16 3 0 7 0 13 3 0 0 9 7 9 0 2
2 0 9
7 0 9 13 3 9 0 2
27 13 1 15 7 9 2 16 13 1 9 3 12 9 7 12 1 15 13 0 9 2 0 9 2 9 2 2
12 9 0 2 0 9 2 7 13 7 9 0 2
18 12 1 0 9 0 9 15 3 13 0 0 9 9 11 11 2 11 2
29 0 0 9 1 0 9 3 3 13 1 9 1 9 7 9 2 0 2 9 2 1 10 9 1 9 0 7 0 2
36 0 2 0 9 2 9 0 9 9 2 0 9 2 1 9 7 9 9 2 7 0 9 13 1 10 0 0 2 9 9 3 0 7 3 0 2
26 1 11 13 7 11 11 2 9 0 0 9 9 2 9 2 7 9 1 9 2 9 1 0 9 2 2
32 12 9 3 13 0 0 9 2 1 10 0 9 2 1 0 9 11 11 2 11 1 11 2 9 0 7 0 2 3 13 9 2
2 0 11
11 9 11 3 13 0 9 9 0 7 0 2
19 1 9 13 0 11 11 10 0 9 0 0 9 0 9 2 0 9 2 2
29 1 9 9 15 7 1 15 2 7 1 0 11 11 2 13 4 15 1 0 9 2 1 9 0 0 9 2 13 2
25 1 9 4 13 7 0 0 9 11 11 11 1 9 9 2 9 2 2 0 1 0 9 0 0 2
19 1 9 11 13 3 0 9 0 9 2 15 16 10 0 9 13 11 11 2
46 0 9 0 9 2 0 9 11 1 11 2 9 0 9 11 2 13 1 0 9 10 0 0 9 9 2 0 9 2 3 13 1 0 0 9 2 10 9 1 9 13 12 9 9 2 2
18 0 9 15 13 1 9 2 10 0 9 0 0 9 13 1 0 9 2
12 9 13 3 0 9 7 3 13 10 0 9 2
23 13 15 1 9 0 0 9 2 15 13 13 1 0 9 7 10 9 15 13 13 0 9 2
25 9 13 0 2 0 9 2 1 9 1 9 9 1 0 9 7 9 2 3 0 9 13 0 9 2
17 15 7 13 1 0 0 9 0 3 14 1 0 9 9 0 11 2
19 9 4 15 13 13 1 9 0 0 9 2 3 15 13 13 3 0 9 2
4 0 9 0 9
17 12 1 0 9 0 9 13 9 7 0 9 0 0 9 7 9 2
24 0 13 15 1 0 9 2 3 0 9 13 13 9 3 0 2 15 3 3 3 13 0 9 2
21 3 15 7 1 0 9 13 3 9 1 0 9 2 15 4 0 9 11 3 13 2
9 3 7 9 13 0 9 0 9 2
22 0 9 10 9 13 0 9 16 13 9 2 16 9 13 0 2 9 2 11 11 2 2
22 13 9 0 9 1 0 0 9 7 0 9 1 0 9 2 15 13 3 1 9 2 2
18 1 0 2 3 2 16 3 0 0 0 9 13 3 1 0 0 9 2
14 1 11 4 3 13 2 16 9 15 13 1 15 13 2
6 7 0 9 3 3 2
3 9 0 9
43 16 13 1 9 9 0 0 9 13 10 0 0 9 2 13 4 15 13 1 9 0 9 2 9 1 0 7 0 9 2 7 0 9 0 2 0 9 2 0 1 0 9 2
38 1 11 3 3 3 13 0 2 0 2 0 7 3 0 9 1 2 0 9 2 2 0 9 9 2 0 0 2 9 2 0 0 9 2 3 2 2 2
22 9 15 1 15 13 1 0 9 7 9 9 2 9 7 1 0 9 9 0 7 0 2
17 3 13 0 9 0 9 7 0 9 2 0 0 0 7 0 9 2
18 9 13 3 0 2 3 0 7 0 9 1 0 2 3 0 9 9 2
23 13 9 0 9 16 9 1 9 7 9 0 9 2 9 9 0 9 2 9 9 7 9 2
6 13 0 7 13 9 2
16 9 11 11 7 9 11 11 1 9 9 15 13 1 0 9 2
3 9 1 11
2 11 2
25 9 12 0 0 9 3 13 9 1 9 9 1 0 0 9 11 7 1 9 9 1 9 9 11 2
31 9 4 13 1 11 11 11 7 0 9 11 11 11 2 1 15 0 14 3 13 9 9 2 11 13 9 7 11 9 11 2
16 12 9 15 13 1 9 9 1 9 9 7 1 9 9 9 2
9 3 13 9 1 9 0 0 9 2
5 0 9 1 15 9
36 1 0 9 1 9 9 1 0 9 13 0 13 1 9 2 16 0 9 2 15 15 13 0 0 9 2 13 1 0 7 0 9 12 1 0 2
24 10 9 4 13 1 0 9 13 3 0 9 2 15 13 1 0 13 1 9 0 9 0 9 2
26 9 15 13 13 2 0 9 13 0 9 1 0 9 7 13 15 0 9 0 7 0 9 10 0 9 2
30 1 9 0 9 0 9 9 3 7 13 1 9 13 7 13 0 9 2 15 2 15 13 13 9 9 0 9 0 9 2
22 1 0 9 13 9 13 0 9 0 9 1 0 9 1 0 9 2 15 13 9 0 2
24 10 9 4 13 9 9 2 0 9 1 0 9 2 7 2 0 9 1 9 15 0 9 2 2
8 1 0 9 4 13 3 3 2
10 3 4 13 13 10 9 1 0 9 2
11 9 13 3 0 7 9 13 13 15 13 2
7 0 13 7 9 0 9 2
28 9 3 13 9 2 3 0 7 0 9 13 9 1 0 9 1 9 2 16 9 0 9 1 10 9 0 13 2
34 3 13 1 15 2 16 0 9 13 13 9 1 9 2 7 13 3 3 9 1 10 9 2 7 16 15 1 9 9 13 0 0 9 2
23 15 3 13 9 10 9 2 9 9 7 9 9 2 9 2 15 15 1 0 9 3 13 2
19 9 1 9 0 9 2 2 9 15 9 1 0 9 2 2 15 3 13 2
11 3 0 9 13 1 0 9 13 12 9 2
37 12 1 15 13 13 9 0 9 9 1 15 9 2 0 9 2 2 3 7 13 13 7 0 9 2 15 13 3 13 7 0 9 0 9 13 9 2
17 15 4 7 13 2 16 0 0 9 13 1 15 3 0 7 0 2
31 16 3 13 7 0 7 0 9 1 9 3 0 2 3 13 9 7 9 9 2 15 13 10 9 1 9 3 0 7 0 2
11 13 4 4 3 13 7 1 9 0 9 2
21 3 4 15 13 9 9 0 0 9 2 16 9 9 4 1 0 9 3 3 13 2
20 0 0 9 0 9 4 13 0 9 2 3 2 3 13 15 1 9 1 9 2
27 9 1 9 0 0 7 0 9 13 1 3 0 2 1 0 3 2 16 3 13 0 0 9 0 0 9 2
41 16 13 0 9 9 9 9 1 9 0 9 2 13 3 1 15 2 16 4 4 0 9 13 7 1 0 9 2 3 13 1 0 9 7 3 9 13 3 0 9 2
12 13 7 0 9 2 15 13 13 3 0 9 2
17 9 0 9 13 0 9 7 1 9 13 4 13 0 9 0 9 2
48 3 15 4 13 12 0 9 1 0 9 2 10 9 4 13 9 1 0 0 9 2 0 9 9 1 0 9 7 9 0 9 9 7 9 9 2 7 15 16 0 9 2 7 7 9 9 9 2
32 0 9 13 2 16 4 10 9 13 16 0 9 7 13 0 9 1 9 1 0 9 1 9 12 9 2 13 3 9 0 2 2
24 10 9 4 13 13 7 1 9 2 3 7 1 9 0 9 2 0 9 1 9 16 9 0 2
48 0 9 1 0 9 10 9 2 3 0 1 9 0 0 9 7 0 9 0 9 7 0 9 9 2 13 13 9 3 2 3 7 3 2 1 9 2 7 1 9 0 7 0 0 9 1 9 2
7 11 2 9 1 9 13 0
3 1 0 9
2 11 2
19 9 3 3 13 9 2 13 15 9 9 7 13 10 9 13 9 0 9 2
18 13 15 15 1 0 9 11 7 0 9 0 9 2 0 7 0 9 2
19 9 11 11 11 1 15 3 13 2 16 9 10 9 1 0 9 13 0 2
15 9 11 15 3 3 13 1 9 9 9 7 0 9 9 2
16 1 11 13 9 9 1 9 9 9 1 9 0 9 0 9 2
1 3
16 9 11 11 13 1 9 1 9 11 1 11 1 12 9 9 2
17 0 9 11 11 13 2 16 12 1 0 13 3 9 11 11 11 2
17 11 7 3 13 2 16 9 13 15 0 7 13 15 14 0 9 2
18 9 2 15 13 9 1 9 1 9 1 9 7 9 9 2 13 0 2
11 1 9 9 7 4 13 3 14 1 9 2
6 3 13 0 9 13 2
16 9 9 13 13 13 12 9 0 1 10 9 9 3 1 9 2
9 0 9 4 9 3 13 9 9 2
21 13 15 9 9 2 15 10 9 13 1 9 1 9 9 2 15 15 13 1 9 2
14 11 11 15 1 11 13 3 9 10 9 9 1 9 2
8 10 9 13 1 10 0 9 2
1 3
11 1 11 0 9 13 3 3 0 16 0 2
35 16 9 9 0 9 1 9 13 1 0 9 3 12 9 2 3 12 9 2 2 0 9 9 1 11 13 1 12 9 2 3 12 9 2 2
14 11 2 11 2 11 2 11 7 11 2 11 1 9 9
5 9 2 9 2 9
2 0 9
4 13 15 3 2
7 9 13 3 0 16 9 2
4 16 13 9 2
48 9 13 9 0 2 3 0 7 3 0 2 9 7 9 1 0 7 0 2 7 3 3 3 9 1 9 1 9 2 9 9 9 1 9 2 9 1 9 2 7 3 3 9 9 1 0 9 2
19 13 15 3 0 2 16 7 1 3 0 9 15 13 9 14 3 0 2 2
17 3 2 3 4 9 7 0 9 7 9 13 0 9 13 13 9 2
42 3 2 16 0 0 9 1 9 13 2 9 2 3 2 10 9 2 13 2 0 9 2 2 3 1 9 7 1 9 10 0 9 13 9 1 9 1 9 1 11 9 2
2 9 2
12 9 13 1 0 9 9 2 7 0 0 9 2
47 15 3 0 9 13 1 10 0 0 9 9 7 9 2 16 15 0 13 13 0 2 0 9 2 16 15 0 13 3 9 13 2 7 15 3 1 0 9 1 9 2 9 2 9 2 9 2
24 7 9 0 9 1 0 9 13 14 0 0 2 9 9 7 9 2 2 7 0 7 0 9 2
9 1 10 9 9 13 1 9 9 2
23 9 9 13 4 13 7 13 1 15 9 0 9 10 10 9 2 13 15 13 1 0 9 2
23 16 13 13 9 3 3 0 9 7 0 9 2 7 3 9 9 16 9 2 3 7 9 2
11 7 3 7 9 13 0 9 7 0 9 2
19 3 2 13 1 15 7 9 9 2 16 13 13 0 2 9 13 9 2 2
15 1 9 4 15 9 13 16 9 0 2 0 2 3 3 2
11 13 15 7 2 0 2 9 1 0 9 2
38 7 13 1 10 0 9 0 9 13 13 15 9 1 9 0 2 16 9 13 14 15 2 15 3 13 2 7 7 15 15 13 7 13 13 13 9 0 2
15 9 1 0 9 13 13 2 13 4 12 1 0 0 9 2
30 13 15 2 16 4 9 13 13 0 10 9 0 2 0 2 9 7 9 0 9 2 3 13 15 3 2 1 11 2 2
41 13 4 7 13 2 1 9 2 3 1 9 9 0 7 0 2 7 13 0 9 9 2 7 3 13 9 9 1 9 12 1 0 9 0 9 2 3 1 9 0 2
32 0 9 2 10 0 7 0 2 13 7 13 0 9 0 2 0 9 16 9 9 7 9 2 7 15 1 10 0 0 0 9 2
37 13 9 1 0 9 2 3 1 9 0 0 9 13 0 9 2 0 10 9 2 7 1 9 0 2 0 14 7 14 3 2 7 2 3 7 3 2
25 14 2 7 9 13 4 13 1 10 0 2 0 9 2 3 16 9 0 9 2 16 9 3 0 2
21 3 13 7 9 2 3 9 9 13 10 9 1 0 2 0 9 1 9 9 0 2
9 1 3 0 9 13 10 0 9 2
28 9 2 0 7 0 2 4 3 13 1 0 9 2 7 15 14 3 2 7 7 3 2 3 3 13 10 9 2
11 9 13 2 13 9 7 9 0 0 9 2
4 0 11 3 13
2 11 2
35 1 0 0 9 13 11 11 1 11 11 12 2 12 1 9 2 16 9 12 2 12 1 9 0 9 13 1 9 11 11 1 9 11 11 2
32 11 11 1 9 11 13 12 9 9 0 11 11 2 7 11 7 1 0 9 1 15 13 7 13 15 13 1 9 12 2 12 2
29 3 3 15 7 13 1 9 13 0 9 7 9 11 11 11 2 15 1 9 12 2 12 13 1 0 9 12 9 2
15 0 9 13 0 9 1 9 12 2 3 15 13 9 9 2
8 11 11 1 9 1 9 1 11
6 13 1 9 7 13 9
14 13 15 3 3 2 3 1 0 0 9 13 9 9 2
12 1 9 13 1 0 2 2 9 2 9 2 2
23 16 9 4 15 13 15 2 16 4 1 0 9 13 3 3 2 9 13 2 9 13 2 2
27 13 4 15 1 10 9 1 9 2 3 10 9 13 2 16 9 4 13 1 0 9 2 7 1 10 9 2
25 7 13 4 15 15 2 9 2 16 13 1 9 7 1 9 13 1 0 2 2 9 2 9 2 2
8 9 10 9 1 15 15 13 2
4 15 13 9 2
8 1 0 9 15 7 3 13 2
19 16 0 13 9 3 1 0 9 2 9 13 14 1 0 9 3 1 9 2
9 13 1 15 16 0 2 0 9 2
10 0 9 0 9 10 9 13 1 9 2
6 9 7 13 3 3 2
9 13 9 13 7 1 9 10 9 2
8 14 4 0 9 13 3 0 2
3 7 3 2
14 0 9 0 9 4 14 13 13 1 12 9 3 3 2
6 9 2 9 2 9 2
7 14 2 15 15 13 0 2
9 13 4 15 0 9 9 2 2 2
37 9 10 9 13 15 2 16 1 9 9 4 3 7 3 0 9 9 1 10 9 13 2 1 9 15 13 3 14 15 2 15 15 1 9 9 13 2
15 7 2 13 3 7 3 7 3 3 13 0 9 1 9 2
6 13 15 7 1 9 2
5 3 4 9 13 2
14 9 2 9 2 13 15 2 16 4 15 9 3 13 2
16 13 2 7 15 4 15 3 3 13 1 0 9 7 0 9 2
17 11 13 1 9 9 15 9 2 16 4 13 1 0 9 15 0 2
15 13 10 9 2 13 4 7 15 15 0 1 0 0 9 2
15 13 15 2 16 4 15 9 13 3 3 2 3 0 9 2
14 1 15 4 1 9 13 3 2 9 3 14 13 9 2
16 7 3 13 1 9 7 13 1 9 2 9 2 9 2 2 2
4 13 9 11 11
26 0 9 7 9 11 11 2 15 15 13 0 9 9 1 0 9 2 13 1 9 3 1 9 12 9 2
20 10 9 1 9 9 11 12 2 7 9 9 11 11 4 3 13 1 9 12 2
14 1 12 9 3 4 9 13 7 11 13 11 1 9 2
35 11 1 0 9 3 13 1 0 9 11 11 7 13 15 1 10 0 9 9 11 1 11 2 9 11 2 1 15 3 13 11 2 7 11 2
24 11 2 15 7 0 9 1 0 9 13 1 9 2 3 1 9 13 0 9 1 0 11 11 2
10 13 15 0 9 1 9 9 1 0 2
23 9 9 2 12 9 0 9 1 9 12 13 0 9 13 10 9 7 2 0 9 1 9 2
36 0 9 0 9 2 15 15 0 13 9 1 9 1 9 0 9 2 1 9 13 2 16 0 9 3 15 1 9 13 2 7 10 9 13 9 2
53 9 0 9 1 9 13 3 0 9 2 15 13 9 10 9 0 1 9 9 9 9 0 2 0 7 10 9 1 9 1 10 9 1 3 0 2 15 13 9 1 9 1 9 9 9 1 10 12 2 9 0 9 2
31 9 13 9 1 15 2 16 15 1 9 9 13 9 10 9 7 9 0 2 0 9 0 7 9 9 1 9 1 9 9 2
42 1 0 9 15 13 0 2 15 1 10 0 0 9 13 12 0 9 9 7 13 0 9 2 15 4 13 9 1 10 9 2 12 2 13 7 13 9 9 3 0 9 2
21 12 2 13 15 9 3 0 9 2 9 7 9 9 9 7 9 9 1 0 9 2
9 12 2 9 9 7 9 0 9 2
23 3 16 13 0 13 9 7 9 2 13 0 13 0 9 7 9 9 1 9 1 3 0 2
30 13 13 3 1 9 7 9 1 10 9 2 7 9 0 0 9 13 9 9 1 9 1 9 9 1 0 9 1 9 2
7 2 9 2 1 2 9 2
18 10 9 13 9 0 1 10 9 2 3 15 13 0 9 1 9 0 2
28 9 9 1 11 13 9 1 11 9 12 2 9 0 15 3 13 1 15 2 16 0 9 13 15 0 7 0 2
32 13 15 1 0 9 1 9 2 15 15 13 9 2 16 0 13 13 2 15 13 3 2 15 3 2 15 13 3 2 13 0 2
32 0 9 4 13 1 0 9 16 0 9 2 4 13 1 15 2 15 0 13 7 13 1 0 9 7 13 10 9 15 1 15 2
14 0 9 0 9 13 10 9 1 9 9 1 9 0 2
38 1 10 9 9 15 0 13 13 9 1 10 9 7 13 15 16 0 9 2 15 13 10 9 2 3 7 15 2 16 9 10 9 1 15 13 1 9 2
9 14 0 9 0 13 3 0 9 2
20 0 9 3 13 2 16 13 2 16 4 9 13 0 16 15 2 16 4 13 2
20 1 9 0 13 3 0 13 2 16 0 9 13 0 9 9 9 1 9 9 2
16 2 9 15 15 13 13 1 9 2 13 10 0 9 9 2 2
14 15 0 13 3 0 13 2 16 0 13 15 15 15 2
4 9 1 9 2
12 9 0 1 0 9 1 15 13 3 10 9 2
14 9 9 1 15 13 13 0 9 2 15 13 0 9 2
25 3 1 11 13 0 9 2 3 0 9 15 13 16 0 7 9 16 0 0 9 2 1 12 9 2
36 1 9 12 13 1 0 9 0 9 16 0 9 2 16 15 13 3 3 2 3 15 13 13 2 16 15 4 1 10 9 3 13 0 9 2 2
7 1 9 13 3 0 9 2
29 13 0 9 13 1 9 1 9 2 3 3 13 9 1 9 2 16 4 1 9 13 3 9 2 15 13 0 9 2
34 9 4 3 13 13 0 9 3 2 16 4 15 1 15 13 14 0 13 1 10 9 2 7 16 4 10 9 13 13 9 2 13 9 2
28 7 3 13 3 0 9 2 3 15 0 9 13 7 3 13 10 0 9 2 16 13 9 2 15 4 9 13 2
42 0 9 13 0 13 1 9 0 1 9 0 2 9 0 15 13 1 9 0 9 1 0 9 2 11 2 11 2 11 2 7 3 4 15 3 13 0 9 13 10 9 2
41 16 15 13 0 9 1 9 2 13 9 15 13 2 13 9 2 13 9 9 9 2 15 13 3 2 9 9 0 9 2 15 13 0 9 1 9 0 9 11 11 2
12 16 4 9 13 10 2 14 15 0 13 3 2
23 0 1 9 13 3 13 2 9 9 1 9 2 7 13 9 9 0 7 9 1 9 9 2
12 9 4 13 13 9 1 9 9 1 0 9 2
16 15 3 13 2 16 0 9 7 9 4 3 7 3 13 3 2
24 9 9 4 13 3 13 9 2 16 4 15 13 2 1 9 1 9 2 13 2 10 9 13 2
10 16 9 15 13 2 1 9 15 13 2
21 13 1 0 0 9 2 15 13 7 13 9 13 2 1 15 15 13 7 0 9 2
48 10 9 13 13 9 2 9 7 9 9 2 15 4 9 13 13 2 3 13 9 2 9 2 9 1 10 9 2 3 13 10 9 2 15 13 13 0 9 2 3 0 0 9 2 1 10 9 2
16 9 16 1 9 2 13 15 2 1 10 9 15 13 9 9 2
26 1 9 9 1 9 4 13 13 9 0 0 9 1 10 0 9 1 9 9 2 15 15 13 1 9 2
3 0 9 9
16 12 13 0 9 7 0 9 0 2 13 15 3 2 15 3 2
21 0 9 1 9 13 13 3 1 9 7 10 9 13 0 9 3 12 9 1 9 2
20 0 9 2 1 15 15 13 9 1 0 0 9 2 13 3 3 1 0 11 2
20 0 9 15 3 13 15 12 9 2 15 3 13 10 9 13 15 9 0 9 2
29 16 9 13 14 1 9 2 13 15 10 9 0 9 2 13 15 1 15 0 9 7 13 15 3 16 0 0 9 2
18 1 0 9 4 13 9 9 7 9 9 1 9 1 9 0 0 9 2
17 9 0 9 2 16 1 15 3 13 2 15 7 13 1 0 9 2
20 0 13 12 9 2 0 9 11 11 2 0 9 11 11 7 9 11 11 11 2
6 15 15 9 13 3 2
23 0 9 11 11 13 9 1 0 9 7 1 9 13 0 9 1 3 0 2 7 0 9 2
28 9 11 11 2 0 1 9 0 9 0 9 15 1 9 13 14 3 2 16 16 0 1 9 13 9 1 9 2
8 0 9 3 1 0 9 13 2
36 1 9 7 13 12 3 0 9 9 2 0 9 0 9 11 11 2 1 9 1 12 9 14 3 1 11 2 7 9 0 11 11 11 2 11 2
10 11 15 3 3 1 0 0 9 13 2
19 3 2 3 16 9 11 2 13 2 16 15 9 13 1 15 7 13 9 2
9 10 9 7 1 15 13 0 9 2
29 16 0 9 13 1 9 2 3 3 15 15 3 13 0 9 2 15 15 1 9 1 9 13 13 9 1 0 9 2
16 16 7 4 13 0 9 16 10 9 2 13 9 1 9 0 2
7 1 11 13 10 0 9 2
21 10 9 2 7 13 15 1 10 9 3 10 2 13 0 9 9 0 9 0 9 2
11 13 0 2 16 1 10 0 9 13 9 2
25 9 2 15 1 10 9 13 2 13 1 10 0 9 9 1 9 0 9 2 1 15 3 3 13 2
36 13 15 2 16 9 10 2 9 2 13 2 15 15 13 2 3 3 2 16 4 1 0 9 13 3 0 2 0 2 9 0 9 1 0 9 2
8 9 11 13 3 13 1 9 2
34 16 13 1 9 9 9 2 11 1 9 2 0 9 2 2 1 9 9 9 2 13 9 1 0 9 2 3 15 15 15 3 3 13 2
14 3 15 13 1 0 9 13 3 13 2 15 13 0 2
26 16 4 11 11 3 3 13 7 3 2 13 3 0 9 2 15 1 0 9 13 1 9 12 0 9 2
6 2 9 13 1 9 2
10 0 0 9 11 2 11 1 9 9 11
15 2 9 1 9 9 0 9 11 11 1 11 13 1 9 2
31 0 9 0 0 9 2 3 11 11 2 3 13 0 9 2 3 3 0 9 13 13 2 2 13 9 11 1 9 1 11 2
33 9 0 9 0 9 13 2 16 15 3 1 0 9 3 13 9 1 0 9 7 11 2 7 10 0 9 1 0 9 10 9 13 2
18 2 11 3 3 13 2 16 13 2 14 1 9 2 13 15 1 9 2
35 3 3 15 13 0 9 0 0 9 2 15 3 13 1 9 1 0 11 2 7 13 1 11 0 9 2 16 1 9 13 2 2 13 9 2
42 1 0 9 10 0 9 2 16 0 9 0 0 9 2 3 0 2 4 13 1 0 9 2 7 7 13 0 3 13 10 9 7 3 7 13 9 12 9 2 13 9 2
22 2 9 1 0 9 13 14 3 0 7 7 15 13 13 10 0 0 9 9 10 9 2
40 3 0 9 13 9 2 16 10 9 13 14 14 15 13 0 0 9 2 7 3 1 9 1 10 9 13 3 0 1 0 9 2 2 13 0 9 9 1 9 2
9 0 9 3 13 7 1 0 9 2
14 2 1 11 13 9 13 9 0 9 7 1 0 9 2
36 14 2 1 10 9 15 13 9 1 9 15 0 9 1 11 2 2 13 11 7 13 2 16 2 1 11 4 14 13 1 12 9 12 9 2 2
30 2 3 3 13 1 3 0 9 2 15 13 9 3 13 2 2 13 1 0 0 9 11 1 9 12 9 9 1 11 2
18 1 10 9 10 9 13 9 0 9 1 9 7 9 7 11 1 11 2
33 2 0 9 3 13 3 1 2 7 1 10 0 9 15 13 13 0 9 2 3 1 9 11 2 2 13 10 9 1 9 0 9 2
22 2 3 13 1 0 0 9 2 16 4 2 14 9 11 13 11 2 13 15 1 11 2
24 3 15 13 13 1 9 9 7 1 15 2 16 4 13 3 0 1 0 9 9 7 9 2 2
19 0 13 1 0 9 7 9 9 2 16 3 1 0 9 15 13 0 9 2
25 11 13 7 13 9 2 16 9 1 9 0 9 13 13 0 9 1 9 12 9 0 9 1 11 2
52 1 10 9 2 0 13 13 2 0 9 2 16 9 1 0 9 1 11 15 13 16 0 2 16 13 0 15 13 2 16 11 13 13 1 9 0 9 7 9 7 9 1 0 9 2 15 13 0 13 0 9 2
15 9 13 11 0 2 13 15 7 9 1 12 1 12 9 9
2 11 2
22 0 9 1 11 3 13 1 0 9 9 11 11 1 12 9 1 0 12 9 9 9 2
28 13 15 0 2 16 3 1 9 12 7 3 1 9 12 13 12 0 9 7 13 15 3 14 1 12 12 9 2
22 9 11 11 3 1 9 9 13 2 2 10 9 13 9 9 2 7 7 13 9 2 2
11 11 13 2 16 9 13 1 9 0 9 2
11 11 15 1 9 9 13 2 16 13 0 2
10 9 13 16 9 0 1 0 0 9 2
13 9 13 0 9 1 9 9 0 1 9 12 9 2
17 1 9 13 7 0 9 0 7 16 0 9 2 14 16 9 0 2
25 9 3 10 9 13 3 2 16 13 1 0 9 1 9 7 1 15 2 16 15 13 2 15 13 2
13 16 2 13 9 2 1 15 13 2 0 9 2 2
11 1 0 9 13 1 11 16 9 9 9 2
6 7 10 9 13 0 2
30 16 0 9 1 9 13 2 16 15 13 0 2 16 13 9 2 0 15 3 13 1 9 2 7 3 1 9 1 9 2
22 9 15 3 0 9 3 1 9 13 2 1 16 4 15 13 7 3 13 1 9 9 2
23 16 10 9 3 13 2 3 13 1 9 12 0 9 9 2 13 10 9 9 1 9 0 2
23 1 9 11 13 3 15 2 16 1 9 1 9 2 3 1 9 13 2 4 13 10 9 2
27 9 3 13 2 3 4 13 1 10 9 3 9 11 2 3 13 15 9 2 7 13 15 3 1 9 9 2
10 13 4 1 9 9 9 9 1 9 2
10 0 9 13 9 11 11 2 1 9 2
2 11 2
22 0 9 9 0 7 0 9 15 3 13 1 9 2 15 13 9 11 11 2 11 2 2
13 13 15 1 15 2 16 4 15 13 1 9 9 2
19 11 3 1 9 9 1 9 13 7 3 1 15 15 2 13 2 9 9 2
50 3 13 10 9 9 13 9 2 15 4 13 9 11 2 16 4 13 2 16 9 13 9 1 9 11 1 0 9 1 10 0 0 9 1 9 9 7 1 9 9 2 16 15 1 9 10 9 3 13 2
33 1 10 9 15 7 13 0 9 11 11 7 11 11 7 11 11 2 11 2 1 15 2 16 4 15 1 15 13 14 1 0 9 2
28 1 9 11 13 2 16 4 9 9 0 11 11 1 11 3 13 2 7 3 3 15 13 2 16 1 15 13 2
5 9 13 3 1 9
2 11 2
16 1 0 13 9 9 9 1 9 9 9 1 9 9 0 9 2
21 1 9 0 9 7 9 9 13 2 16 9 0 9 13 1 9 9 3 0 9 2
9 13 14 15 9 2 3 15 13 2
19 2 1 0 9 9 1 0 9 14 1 9 9 2 2 13 15 1 9 2
23 0 9 2 9 2 15 1 9 9 13 13 9 2 13 15 9 1 9 7 13 15 9 2
7 9 9 0 0 9 11 13
2 11 2
11 0 9 11 13 1 12 9 2 9 11 2
23 0 0 9 1 11 13 12 9 9 2 1 11 7 11 12 9 7 1 11 12 9 9 2
12 1 9 11 7 11 9 3 15 1 9 13 2
8 13 15 1 9 0 0 9 2
24 1 9 9 7 11 10 0 9 13 9 0 0 9 2 3 13 7 0 15 13 1 0 9 2
10 0 9 13 0 11 13 1 9 12 2
12 1 9 0 9 13 9 0 9 0 0 9 2
20 1 9 12 7 12 13 0 9 9 2 7 10 0 0 9 3 13 0 9 2
12 1 9 12 3 13 0 0 9 0 0 9 2
22 1 9 0 9 13 1 0 9 10 9 3 0 9 9 2 15 4 13 1 9 12 2
5 3 9 2 9 12
3 9 9 13
2 11 2
27 9 9 9 11 1 9 1 9 13 9 10 9 1 0 9 12 9 1 9 2 15 13 10 0 0 9 2
23 13 15 3 9 1 9 1 11 7 10 0 9 1 9 0 9 1 9 1 9 0 9 2
14 1 0 12 9 9 9 1 11 13 1 0 12 5 2
16 3 13 7 3 1 9 9 0 16 3 2 3 13 0 9 2
17 3 1 15 13 9 1 9 1 11 2 15 13 0 0 9 9 2
5 9 13 3 1 9
16 1 0 9 13 0 9 7 10 9 15 7 13 7 3 3 13
29 9 9 7 0 9 2 15 1 10 9 13 1 12 9 2 1 15 1 9 1 9 13 10 3 1 9 0 9 2
19 9 1 0 9 1 0 15 1 0 13 9 3 0 9 7 0 9 0 2
15 12 1 0 9 2 15 15 3 13 0 9 2 13 9 2
17 9 13 0 9 2 0 15 9 7 9 0 9 1 0 9 9 2
13 9 0 9 13 0 9 1 9 0 7 0 9 2
17 0 0 9 1 11 13 1 10 9 0 9 10 9 1 0 9 2
16 1 0 12 9 13 1 10 9 1 3 0 0 9 0 9 2
26 1 0 9 0 9 13 0 0 9 0 9 1 0 0 7 0 9 2 15 13 3 3 7 3 0 2
21 7 1 1 0 9 9 1 0 9 9 11 13 1 10 9 0 7 0 0 9 2
28 9 13 16 0 9 13 1 0 2 0 9 9 0 7 1 3 0 9 9 7 9 1 0 9 0 1 11 2
9 0 9 9 1 11 13 12 9 2
12 0 2 0 9 2 13 13 3 1 0 9 2
26 9 15 1 9 10 9 13 0 7 0 9 1 9 9 2 9 2 0 9 2 9 9 7 9 9 2
6 3 13 0 0 9 2
14 0 0 9 13 9 0 9 7 13 2 0 2 9 2
22 0 9 2 15 3 13 0 9 2 13 1 9 3 13 1 0 9 0 9 1 11 2
19 0 2 0 9 2 13 13 7 1 9 9 9 2 3 2 2 7 3 2
20 1 0 9 9 9 1 0 9 9 7 9 0 9 0 13 3 3 12 9 2
13 1 0 9 15 13 1 9 0 3 12 9 9 2
17 1 0 9 13 0 9 7 10 9 15 7 13 7 3 3 13 2
28 13 9 1 0 0 9 2 9 2 9 2 0 9 2 1 0 0 9 7 3 1 9 0 15 9 0 9 2
6 9 13 0 9 1 11
2 11 2
21 0 9 11 13 1 9 12 2 7 12 2 9 0 7 0 9 1 11 7 11 2
24 2 0 9 13 0 9 0 9 1 10 0 9 2 2 13 3 9 9 0 9 9 11 11 2
17 9 13 9 9 7 9 9 7 9 2 15 13 9 12 0 9 2
16 0 0 9 13 3 11 11 2 11 11 7 0 7 0 9 2
22 9 11 3 1 9 13 1 11 9 1 9 0 9 1 9 12 1 9 12 9 9 2
24 0 0 9 13 2 16 1 9 13 3 0 0 9 7 9 13 7 12 0 0 9 0 9 2
21 11 11 0 2 12 13 0 9 2 0 9 7 9 2 9 0 9 9 0 11 2
5 13 10 0 9 2
4 9 1 9 9
23 13 15 9 12 2 16 15 12 2 9 13 1 11 1 11 0 0 9 11 11 9 11 2
10 1 9 1 0 9 15 13 0 9 2
29 9 9 3 3 13 11 0 9 0 9 2 7 7 15 13 2 16 4 3 0 9 0 9 13 10 0 0 9 2
25 10 9 13 9 1 9 2 12 2 9 12 13 1 11 11 11 2 9 1 11 2 9 7 9 2
13 3 10 3 0 9 13 9 10 0 9 3 0 2
19 9 9 7 9 15 3 13 1 10 9 7 9 2 16 4 10 9 13 2
24 10 9 13 3 9 9 1 0 7 0 9 9 0 9 2 0 1 0 9 0 0 0 9 2
33 3 2 16 0 0 9 13 1 0 9 9 2 7 7 1 0 9 13 0 2 16 9 10 0 9 13 13 9 7 9 0 9 2
32 13 3 0 2 7 13 15 3 1 9 9 0 9 9 2 2 16 3 16 0 9 10 9 13 0 9 2 15 3 13 13 2
9 15 13 7 1 9 9 11 11 2
20 10 0 9 13 3 9 9 2 3 15 15 1 10 9 13 3 10 0 9 2
27 3 15 2 16 10 9 13 1 9 0 0 9 2 15 13 9 2 0 13 0 9 9 2 0 0 9 2
27 13 0 2 16 1 0 9 2 15 13 10 9 9 16 9 9 0 0 9 2 13 0 0 0 9 9 2
19 15 2 15 3 13 1 11 9 7 0 9 2 13 3 9 9 0 9 2
12 13 2 16 16 9 0 9 13 14 0 9 2
12 1 12 9 15 13 1 9 0 9 7 9 2
14 13 3 12 9 2 12 1 15 13 3 1 0 9 2
30 11 11 15 13 13 0 9 2 7 3 1 9 12 15 13 13 9 2 15 13 1 0 9 2 7 13 1 0 9 2
17 1 0 9 4 13 1 9 2 1 15 4 13 3 1 9 12 2
17 0 9 13 1 10 0 9 13 15 9 2 15 4 13 10 9 2
7 13 9 2 9 7 9 2
20 1 9 15 13 1 9 12 7 1 9 12 3 13 9 1 0 9 10 9 2
18 3 13 13 3 1 0 9 2 1 9 12 13 10 9 1 0 11 2
13 13 3 2 12 0 9 7 13 7 10 9 0 2
41 1 0 9 15 13 9 11 2 12 2 12 2 2 11 2 12 2 12 2 2 11 2 12 2 12 2 7 11 2 12 2 12 2 2 15 15 3 16 9 13 2
17 1 9 12 3 9 13 3 15 7 1 12 1 10 9 3 13 2
11 10 0 9 13 0 9 11 11 14 3 2
28 7 3 13 3 0 9 1 0 0 9 2 15 0 9 9 1 9 12 13 13 15 1 9 1 9 0 9 2
26 15 3 13 0 9 1 15 2 16 15 15 13 0 9 2 7 16 15 15 13 13 1 0 0 9 2
19 1 11 9 7 0 9 1 0 9 13 0 9 2 16 13 3 10 9 2
38 1 9 2 3 15 11 13 0 9 13 3 2 13 1 11 3 0 0 9 2 11 2 11 2 11 2 11 7 0 2 2 15 3 3 1 0 9 2
26 14 1 0 9 0 9 15 1 10 2 1 10 9 0 2 9 9 13 9 0 9 13 3 11 9 2
15 13 15 13 0 9 2 15 13 1 3 0 9 0 11 2
31 15 4 3 13 3 0 9 9 7 9 11 11 1 9 9 11 1 9 12 2 15 9 13 1 0 9 2 7 13 9 2
24 1 9 9 4 0 9 13 1 9 0 9 2 9 2 3 15 13 0 2 3 0 0 9 2
17 9 2 15 15 1 11 11 13 0 0 9 2 13 3 3 0 2
36 11 11 13 0 13 16 12 1 9 0 9 9 0 9 2 16 13 10 0 9 1 0 9 0 9 1 9 1 9 0 9 0 9 0 9 2
34 0 9 10 0 9 13 1 15 2 16 1 0 9 0 9 13 3 0 9 0 9 7 3 10 9 7 0 9 13 9 0 9 9 2
25 10 0 9 13 0 9 1 0 9 0 9 2 3 9 10 9 13 9 9 9 9 7 0 9 2
19 1 0 9 10 9 13 10 9 9 7 9 11 11 0 0 7 0 9 2
18 10 9 11 9 13 1 9 2 7 7 13 0 9 9 0 0 9 2
21 3 15 13 3 13 2 16 15 3 4 13 9 1 15 2 15 0 9 13 13 2
11 1 15 15 13 3 1 0 0 0 9 2
26 1 10 0 9 2 1 9 10 9 2 7 1 9 2 15 15 13 13 10 9 1 9 7 13 15 2
15 3 13 13 2 16 3 9 11 11 15 9 13 3 3 2
26 3 1 9 9 13 10 9 0 0 9 9 2 9 7 9 0 0 9 9 0 2 12 2 12 2 2
35 12 3 0 9 10 9 2 11 11 2 12 2 2 9 7 9 0 9 2 7 10 9 11 2 12 2 2 13 1 0 9 0 0 9 2
7 11 11 2 12 2 12 2
9 0 9 2 9 2 9 7 9 2
11 1 12 9 13 1 15 1 0 9 9 2
17 3 1 0 9 15 13 1 0 9 7 13 15 0 1 9 9 2
7 0 9 13 0 10 9 2
24 16 9 13 1 11 2 11 2 11 7 1 11 2 3 15 13 3 1 11 11 7 11 11 2
45 1 10 9 7 0 9 13 1 9 7 0 2 0 9 2 16 15 11 11 13 0 9 2 2 13 15 1 10 9 9 0 9 7 0 9 3 1 9 2 1 9 10 9 2 2
35 1 0 9 4 3 13 9 9 9 2 12 2 2 12 0 9 2 12 2 2 9 1 12 9 2 12 2 2 12 9 9 2 12 2 2
15 1 9 9 9 11 2 12 2 2 0 9 2 12 2 2
4 9 13 16 11
4 9 1 9 12
5 9 13 9 0 2
25 13 4 1 0 9 1 9 11 11 2 12 9 1 9 2 1 9 0 9 2 16 15 3 13 2
24 1 0 2 0 0 9 0 0 9 7 3 0 2 7 0 9 9 7 9 9 15 13 11 2
17 9 3 13 2 14 0 9 13 9 2 16 13 13 9 10 11 2
10 10 11 15 3 13 2 13 4 15 2
10 3 15 1 15 15 13 9 0 9 2
7 0 9 15 13 3 15 2
16 1 9 1 11 2 1 0 9 2 15 4 13 3 7 11 2
30 16 15 0 9 3 13 7 13 2 0 9 3 13 7 0 9 13 0 9 2 3 0 9 9 13 1 0 0 9 2
10 3 3 0 2 3 0 9 13 9 2
22 13 2 13 11 2 9 7 9 10 9 2 3 0 2 0 2 3 9 2 3 9 2
8 16 15 9 13 2 13 3 2
12 16 4 13 9 2 13 15 2 13 2 2 2
19 3 15 13 1 0 9 1 11 2 3 3 1 0 9 9 13 1 9 2
12 7 9 9 12 3 13 9 9 3 1 11 2
10 3 1 0 9 15 13 3 0 9 2
9 13 1 9 0 7 9 1 11 2
18 1 12 2 9 1 11 2 13 9 1 11 2 11 2 11 7 11 2
17 1 0 9 11 14 11 13 9 2 15 13 3 10 0 0 9 2
4 15 15 13 2
7 13 3 9 0 1 9 2
18 9 0 2 0 2 0 0 9 1 9 1 9 13 7 13 1 9 2
10 13 1 9 2 16 4 13 10 9 2
6 1 0 9 12 9 2
9 1 9 15 12 9 13 1 9 2
22 9 1 9 0 1 9 13 9 2 14 2 9 2 0 9 2 9 2 13 15 3 2
4 13 15 0 2
8 3 2 3 13 3 7 3 2
6 14 2 14 2 14 2
4 0 9 13 2
11 9 11 11 2 11 11 2 15 3 13 2
3 0 0 9
8 3 13 9 1 11 1 11 2
4 0 0 9 2
26 1 9 13 0 9 1 9 2 0 9 1 0 9 13 9 1 9 1 9 2 0 11 2 0 11 2
7 1 9 2 3 0 9 2
5 0 2 3 0 2
19 9 0 2 0 2 1 9 13 0 0 9 7 0 9 11 11 11 11 2
11 9 0 2 3 0 9 15 13 1 9 2
4 9 3 13 2
7 1 12 9 13 12 9 2
7 1 0 9 13 1 9 2
9 13 9 13 0 9 1 12 9 2
7 1 12 9 3 13 11 2
9 3 15 13 9 2 3 13 9 2
13 3 2 1 9 12 2 3 13 0 9 0 9 2
11 9 0 9 2 10 0 9 13 3 3 2
6 13 3 9 0 9 2
10 9 15 0 9 13 3 1 12 9 2
11 10 9 14 1 9 13 9 1 9 11 2
17 1 9 15 13 3 9 2 11 15 15 13 2 13 0 2 0 2
18 1 10 9 13 1 11 0 0 9 2 12 12 2 2 3 1 9 2
4 3 3 0 2
6 1 9 11 13 3 2
24 11 2 15 13 1 15 2 16 3 13 15 13 1 9 2 3 13 0 0 9 1 0 9 2
20 11 15 13 1 9 2 3 2 13 9 2 7 3 15 0 12 9 15 13 2
12 9 1 9 13 9 7 9 1 0 0 9 2
37 1 15 13 15 14 0 0 9 2 0 9 2 9 2 9 2 1 12 9 2 2 2 9 2 9 2 1 10 0 9 15 13 13 9 2 2 2
4 1 9 9 2
9 9 13 3 2 3 1 12 9 2
21 16 13 3 2 13 15 1 12 7 13 3 2 14 2 9 2 9 13 15 13 2
8 1 9 13 0 9 1 9 2
7 15 13 9 2 15 9 2
10 13 3 2 1 9 1 11 0 9 2
5 9 1 0 9 2
13 3 13 0 0 9 2 9 11 3 1 0 9 2
5 0 9 13 9 2
15 16 1 11 3 13 0 9 2 3 9 2 13 1 9 2
6 13 15 7 3 13 2
10 0 9 2 0 9 2 13 0 9 2
6 9 13 0 0 9 2
7 3 3 0 9 0 9 2
9 9 1 9 2 13 7 13 9 2
12 0 9 9 1 0 9 2 0 1 0 9 2
9 0 9 2 9 3 1 0 9 2
17 9 0 9 2 3 15 13 9 2 10 0 9 2 0 0 9 2
10 10 15 13 9 2 15 13 0 9 2
3 0 9 2
5 9 1 11 11 2
5 3 3 0 9 2
10 15 10 12 0 9 13 3 3 13 2
13 9 2 13 1 11 0 9 3 0 9 1 9 2
6 3 13 3 0 9 2
8 15 13 0 2 13 13 15 2
2 9 9
5 1 9 11 13 2
9 14 4 13 1 11 1 0 9 2
4 13 7 9 2
10 9 1 0 9 13 0 9 9 11 2
15 13 3 9 1 9 1 11 7 11 2 1 15 13 13 2
7 9 15 3 13 9 9 2
12 12 1 11 15 1 10 3 0 9 13 9 2
11 3 13 3 0 0 2 3 3 0 9 2
4 9 1 9 2
10 9 11 1 9 1 0 0 0 9 2
9 0 9 0 0 9 1 9 9 2
8 0 2 0 2 1 9 9 2
37 11 3 13 11 9 3 2 7 13 15 0 9 2 0 2 7 3 3 0 9 1 0 9 11 7 0 9 0 11 11 13 1 9 14 15 0 2
16 13 0 2 1 9 2 0 9 15 3 3 13 1 9 9 2
11 1 15 0 13 3 9 16 9 1 9 2
19 9 2 3 1 9 0 9 2 15 3 13 13 9 2 1 10 9 13 2
10 13 15 1 15 2 15 13 3 0 2
15 9 13 0 2 0 9 1 9 1 9 7 9 0 9 2
22 11 13 10 9 1 0 9 2 9 13 9 1 12 9 2 7 1 9 1 10 9 2
21 2 12 9 13 12 7 12 12 0 9 2 9 1 9 9 1 9 13 12 9 2
7 9 13 3 2 9 9 2
23 9 13 13 12 9 2 0 2 16 13 9 2 13 13 10 9 2 15 13 2 1 9 2
7 0 9 15 13 13 0 2
8 0 9 13 9 2 9 9 2
9 7 15 13 13 9 9 10 9 2
4 13 9 9 2
3 9 9 11
7 3 3 14 13 1 11 2
9 1 9 0 11 13 14 7 11 2
12 3 3 13 13 2 1 0 3 13 3 9 2
6 1 0 9 0 9 2
10 13 15 7 13 3 2 14 2 9 2
12 0 9 15 13 0 9 2 11 2 9 9 2
8 9 1 15 13 7 13 9 2
18 3 3 13 9 0 9 7 3 3 9 1 11 7 0 9 11 11 2
20 3 13 1 9 9 7 1 15 9 1 9 13 9 2 13 15 2 2 11 2
13 1 9 4 13 1 11 2 3 15 15 3 13 2
4 13 1 15 2
5 2 11 2 11 2
8 3 3 13 15 1 15 11 2
9 9 1 9 1 9 11 1 11 2
23 13 4 15 2 7 1 0 9 13 3 9 2 7 3 13 11 9 2 2 13 3 3 2
23 9 11 7 11 13 1 12 9 11 16 9 1 0 0 9 9 1 12 0 9 1 9 2
6 12 9 1 12 11 2
10 1 9 3 0 13 7 9 3 13 2
18 0 9 2 12 9 9 2 2 9 1 9 0 9 2 15 13 15 2
44 9 11 2 15 13 1 9 1 9 12 1 0 11 11 2 0 9 0 9 2 15 7 1 9 13 2 7 1 9 12 13 1 9 9 0 0 0 7 0 9 1 12 9 2
6 0 3 13 16 9 2
43 3 11 2 9 1 0 9 2 1 0 9 2 0 11 11 1 0 9 7 0 9 2 15 13 1 9 3 1 9 1 11 2 13 0 2 2 3 11 2 11 7 11 2
54 10 0 9 1 0 9 1 0 9 2 9 11 13 1 11 11 1 12 7 9 0 9 1 0 9 2 16 3 0 9 1 0 9 13 0 2 11 15 13 9 1 9 7 13 15 13 2 11 13 2 1 15 13 2
14 7 3 4 15 15 1 9 13 2 13 11 1 11 2
14 11 2 13 15 15 2 14 13 9 2 13 15 11 2
4 1 9 7 9
29 13 1 9 9 11 1 0 0 9 11 11 2 11 13 3 3 1 9 2 9 16 9 1 9 3 13 1 9 2
37 11 13 1 9 7 9 2 1 11 2 3 1 0 9 2 13 1 9 9 9 2 12 12 9 2 12 12 9 2 12 9 9 2 12 9 9 2
14 10 9 13 0 2 0 9 2 0 9 2 9 11 2
16 9 13 0 2 13 0 2 3 15 3 3 13 2 13 11 2
16 13 3 12 9 2 13 15 2 3 2 1 9 13 12 9 2
13 12 13 0 2 0 1 9 0 9 13 1 9 2
11 9 13 16 11 2 0 2 13 9 9 2
39 7 1 9 9 2 1 9 9 1 9 9 7 1 9 9 1 9 9 2 13 13 3 1 9 2 13 13 3 1 9 2 3 3 9 13 9 1 9 2
13 13 15 1 0 9 2 3 13 0 13 1 9 2
15 1 9 9 1 9 9 2 13 4 15 3 2 13 11 2
10 3 13 15 0 2 3 1 0 9 2
7 9 13 0 9 2 9 2
44 1 9 12 13 7 10 9 1 0 9 3 13 2 0 9 1 9 7 9 9 13 1 9 9 2 12 9 9 13 0 2 15 13 13 2 16 13 2 7 13 1 15 9 2
15 1 0 9 13 9 7 13 2 15 15 3 13 3 3 2
8 11 13 0 9 9 0 9 2
10 9 13 0 7 0 2 13 3 11 2
8 0 9 3 10 0 9 13 2
7 9 9 13 9 1 9 2
6 9 0 9 1 9 2
13 13 3 2 3 3 13 1 0 9 7 0 9 2
5 9 13 11 0 2
21 13 9 7 3 0 2 0 9 2 15 13 1 10 0 9 2 13 14 15 3 2
8 13 15 2 7 15 13 15 2
11 3 13 1 11 1 9 1 12 9 9 2
7 3 1 12 7 12 9 2
19 15 3 13 13 9 2 16 14 1 0 9 7 3 1 11 15 13 3 2
19 3 15 13 15 0 2 1 12 9 13 9 2 9 2 9 2 0 9 2
4 13 15 11 2
7 9 1 12 9 13 9 2
11 13 15 7 13 15 1 15 14 12 9 2
8 7 16 9 13 11 9 9 2
25 7 1 9 12 2 3 13 2 11 13 1 11 1 9 11 7 3 9 7 1 15 0 0 9 2
16 9 13 1 9 2 16 9 13 9 7 3 13 0 9 9 2
9 13 15 1 0 0 9 0 9 2
19 14 15 13 3 1 12 9 2 3 13 11 2 15 9 3 13 1 9 2
23 16 13 15 3 2 3 13 1 12 9 0 9 1 9 2 15 15 13 0 9 1 9 2
12 9 13 3 0 7 0 9 15 13 3 0 2
12 3 7 1 12 9 9 10 9 1 9 13 2
3 9 13 2
8 1 9 9 13 0 0 9 2
2 9 2
8 3 13 7 13 15 1 9 2
30 13 1 11 11 2 10 0 9 1 11 1 0 9 2 9 2 9 1 0 9 2 0 9 1 10 0 9 7 11 2
4 9 1 11 2
3 9 1 9
13 0 9 9 15 13 1 9 0 9 1 0 9 2
5 13 1 0 9 2
5 0 9 13 0 2
14 9 0 2 13 11 2 16 15 1 9 13 0 9 2
8 9 2 0 0 9 2 9 2
4 9 2 9 2
4 1 15 9 2
3 0 9 2
10 1 9 13 3 1 9 12 9 11 2
6 9 13 1 10 9 2
13 3 7 3 13 0 9 9 7 13 0 0 9 2
7 7 3 10 9 0 9 2
5 1 9 1 9 2
14 11 15 3 13 13 2 13 2 16 15 15 13 9 2
7 7 1 9 2 3 14 2
4 13 10 9 2
26 13 9 7 1 9 3 9 0 0 9 1 9 2 0 9 2 9 1 0 0 9 15 13 0 9 2
12 9 13 3 0 9 2 0 9 2 0 9 2
4 9 3 13 2
4 9 16 9 2
14 10 9 9 13 2 9 7 13 0 9 7 0 9 2
8 1 15 0 9 7 0 9 2
26 0 9 3 13 2 1 12 9 1 0 9 2 2 16 9 15 13 11 1 9 2 7 16 13 9 2
10 13 2 14 12 9 2 13 15 9 2
6 9 15 13 9 12 2
8 3 1 9 11 11 13 9 2
14 0 9 1 0 9 13 1 11 11 3 1 9 12 2
14 1 9 3 13 3 9 2 16 3 13 9 7 11 2
8 3 13 0 9 2 3 11 2
12 13 1 9 9 1 9 2 13 0 0 9 2
6 1 9 15 13 11 2
15 11 2 9 11 11 2 3 1 11 3 13 3 12 9 2
5 13 1 0 9 2
10 9 13 1 0 0 9 7 1 15 2
25 0 9 13 9 2 13 11 2 13 11 0 9 2 9 2 9 2 9 2 9 2 9 2 2 2
20 1 0 11 7 11 2 15 13 1 0 9 9 2 13 1 15 11 3 3 2
11 9 1 9 0 9 0 1 9 0 9 2
33 9 13 0 9 9 2 3 12 9 2 2 0 9 2 14 12 9 2 2 0 9 0 0 9 2 9 7 9 2 2 0 9 2
8 13 15 3 2 3 16 13 2
6 9 13 16 0 9 2
5 11 13 1 9 2
8 11 2 11 7 11 15 13 2
3 13 3 2
11 11 13 10 0 0 9 2 9 13 0 2
2 9 9
7 9 9 11 13 11 11 2
1 9
6 15 0 7 3 0 2
15 3 4 15 15 13 2 13 2 16 13 2 2 3 6 2
16 9 9 13 16 0 9 2 16 9 2 16 10 10 9 2 2
3 13 9 2
18 3 3 2 16 9 13 0 2 1 9 1 0 9 2 3 2 2 2
7 1 10 9 15 13 9 2
18 13 15 13 15 10 9 2 9 7 9 10 9 2 15 13 15 9 2
44 13 2 2 3 16 15 1 10 9 7 3 2 2 13 15 15 2 2 1 9 1 15 3 2 2 9 13 16 2 0 9 2 2 16 7 3 3 7 3 15 13 1 9 2
5 13 13 1 9 2
22 13 9 0 1 9 9 11 2 9 0 0 9 2 7 15 0 2 0 1 0 11 2
8 13 15 1 9 2 13 4 2
15 9 15 13 2 16 4 10 9 13 2 15 15 3 13 2
9 16 9 4 13 2 16 9 13 2
56 16 13 3 1 15 2 7 1 11 11 3 1 9 2 7 16 3 1 0 9 13 2 16 1 15 13 9 2 15 15 3 13 2 7 1 11 11 1 12 2 9 2 2 16 13 9 0 10 9 9 2 15 4 15 13 2
16 3 1 15 13 0 9 2 16 15 15 2 0 2 13 3 2
9 7 3 16 15 3 0 3 13 2
3 7 3 2
12 15 15 13 2 16 3 1 9 10 9 13 2
14 7 15 15 13 13 2 3 13 7 3 1 9 13 2
25 3 1 9 7 9 4 15 13 16 3 0 2 7 0 9 2 16 9 13 9 0 16 0 9 2
7 10 0 9 4 13 13 2
29 16 7 13 0 9 3 0 2 7 16 15 13 3 0 7 0 2 7 14 3 2 16 4 15 3 13 1 11 2
11 13 15 0 9 2 0 1 9 1 9 2
15 13 4 2 16 15 1 9 13 1 9 7 9 9 11 2
3 3 13 2
25 1 0 9 15 15 1 9 13 2 16 13 10 0 9 2 7 3 15 13 2 1 9 3 13 2
31 16 15 3 9 13 2 16 9 13 15 1 9 9 2 16 9 2 13 9 2 4 15 13 2 13 4 1 9 3 9 2
17 13 4 15 2 2 9 13 15 2 15 9 7 9 13 1 9 2
37 7 16 3 9 13 1 15 2 13 15 9 2 13 9 7 13 15 14 0 0 9 2 3 16 13 1 9 2 13 13 2 16 4 15 13 9 2
7 16 9 13 9 7 9 2
7 13 0 9 7 13 3 2
16 7 15 4 3 13 16 9 2 15 13 9 0 9 1 9 2
13 3 3 13 2 15 15 13 2 16 15 13 9 2
22 3 3 4 10 9 2 1 9 2 1 9 1 0 9 2 13 7 3 13 2 2 2
14 14 7 1 10 0 9 4 3 1 9 10 9 13 2
25 13 4 2 16 0 9 3 13 9 2 7 15 13 10 9 2 1 15 13 7 10 0 9 0 2
6 7 7 15 3 13 2
6 1 9 3 7 13 2
4 1 10 9 2
5 15 1 15 3 13
5 15 1 15 3 13
23 9 11 13 3 1 9 1 9 0 9 11 13 15 1 11 7 13 15 15 9 1 9 2
19 13 9 2 16 11 15 13 1 12 9 1 15 3 16 1 0 12 9 2
26 3 7 10 0 9 13 3 0 0 9 7 13 15 2 16 16 4 13 2 13 4 9 1 0 9 2
23 15 7 13 2 16 0 9 3 13 1 9 10 0 9 2 16 13 15 2 13 13 13 2
31 0 9 0 0 9 13 3 3 9 9 7 0 9 15 2 15 3 3 3 13 2 7 3 15 2 15 4 13 3 13 2
30 16 4 0 11 3 13 0 9 10 9 7 13 15 15 16 0 9 2 15 15 15 1 9 13 7 13 0 1 0 2
2 0 9
17 0 9 10 9 13 9 2 15 0 9 13 9 10 3 0 9 2
18 16 4 3 1 9 13 2 13 15 13 0 9 1 0 9 0 9 2
28 16 0 2 9 9 14 1 12 1 9 13 15 9 0 0 9 11 7 3 15 13 2 3 14 13 9 0 2
11 0 9 13 7 10 0 2 16 0 9 2
23 13 15 13 0 9 9 7 9 2 3 12 0 9 9 2 15 13 0 12 9 1 15 2
12 10 0 9 13 3 0 2 7 16 3 0 2
24 0 9 13 3 13 3 1 9 2 15 13 9 10 9 1 9 2 15 13 9 12 0 9 2
40 10 0 2 0 9 2 3 15 13 12 10 9 2 15 13 1 0 9 3 16 0 7 0 9 2 15 3 13 0 9 2 7 3 13 2 15 13 10 9 2
2 0 9
25 15 13 0 9 2 15 3 3 1 11 13 9 0 9 2 7 15 3 13 9 2 13 1 9 2
18 9 0 9 13 2 15 4 0 13 2 16 4 15 15 10 9 13 2
32 0 9 2 10 0 9 15 2 15 3 13 11 2 15 13 0 2 7 13 9 2 16 9 9 13 1 9 2 3 13 9 2
21 0 9 15 3 13 13 16 11 2 7 3 15 13 9 7 3 13 3 0 9 2
18 0 9 4 3 13 13 15 0 2 16 13 2 3 9 1 10 9 2
30 9 0 9 13 10 0 9 2 9 13 15 3 1 0 9 13 10 9 3 2 16 9 0 9 13 15 1 9 9 2
18 11 13 9 0 9 1 0 9 7 10 9 4 13 3 10 9 13 2
7 7 13 1 9 13 0 2
9 7 13 15 9 7 9 0 9 2
15 1 0 9 15 13 13 2 16 0 9 4 13 1 9 2
26 13 15 0 2 16 9 11 13 14 0 0 9 2 15 10 9 13 2 7 16 13 15 3 9 9 2
19 11 11 3 13 2 16 1 9 10 9 13 9 13 1 10 9 7 9 2
25 10 9 13 0 9 2 7 1 15 0 9 2 7 13 7 1 9 2 16 15 4 3 13 9 2
9 9 9 13 1 11 3 1 9 2
31 0 9 13 0 14 1 10 9 2 16 3 13 9 10 9 2 13 13 1 0 9 1 9 7 9 2 13 10 0 9 2
13 1 9 1 10 9 3 13 2 16 13 3 0 2
31 1 0 9 4 15 3 3 13 13 2 16 1 11 13 1 9 13 2 16 13 1 15 0 16 1 9 1 9 7 9 2
24 13 13 2 16 0 9 1 10 9 2 15 1 11 13 3 10 9 2 13 3 14 0 9 2
39 10 9 15 3 3 13 10 9 1 9 9 2 3 0 12 9 2 9 1 0 0 9 2 7 13 15 14 3 0 9 15 2 15 13 7 3 3 13 2
19 0 9 4 13 3 1 9 9 9 2 16 3 13 1 9 7 0 9 2
15 0 9 2 15 15 13 1 11 2 13 3 14 10 9 2
3 9 1 9
50 7 3 2 3 3 2 16 4 10 9 13 3 3 2 13 0 2 1 10 9 15 9 9 2 9 2 9 0 9 7 10 9 2 15 15 13 3 15 2 16 13 0 9 2 13 1 9 10 9 2
14 16 13 1 11 0 9 2 10 9 1 15 3 13 2
5 9 11 11 2 11
5 7 9 1 0 11
8 0 9 13 9 9 11 2 11
4 11 2 11 2
26 13 15 1 9 13 9 11 11 2 15 1 0 0 9 13 1 0 9 2 7 3 13 1 9 0 2
11 1 9 1 0 0 15 9 11 3 13 2
24 9 13 9 0 9 11 1 11 2 15 9 11 11 13 1 9 0 9 2 11 7 11 11 2
26 11 13 1 0 2 0 9 11 13 12 9 2 7 0 9 2 13 14 1 0 9 7 9 9 9 2
22 2 9 4 1 10 9 3 13 14 1 11 11 2 16 4 15 13 1 0 9 11 2
16 16 7 0 9 13 2 1 11 1 15 13 2 2 13 11 2
54 1 9 9 11 0 13 2 15 13 7 15 2 16 15 15 13 13 1 0 0 9 11 2 15 13 1 0 9 9 2 2 1 12 9 4 13 1 11 1 9 11 2 1 9 4 13 12 9 7 15 15 3 13 2
24 3 4 15 13 2 16 15 1 9 0 11 13 3 1 9 13 2 2 13 15 1 9 11 2
25 0 9 11 2 12 2 9 2 12 9 2 12 9 2 12 9 2 9 12 2 12 2 12 9 2
26 13 2 11 2 11 2 2 11 2 9 1 9 1 11 2 2 11 2 11 2 12 13 1 9 2 2
26 13 2 11 2 11 2 12 9 1 11 2 2 0 2 9 1 11 2 2 11 2 9 1 11 2 2
4 9 11 7 11
9 11 13 11 9 1 9 1 0 11
3 0 11 2
31 1 9 1 0 9 0 9 0 11 13 11 3 1 11 12 2 12 2 16 0 9 9 13 1 9 11 1 12 2 9 2
27 1 0 9 15 1 9 13 12 0 9 11 11 1 11 1 9 1 11 2 1 12 9 13 1 0 11 2
18 3 1 12 2 9 15 13 9 1 0 9 7 10 9 11 11 11 2
22 9 9 7 13 11 11 2 15 13 10 0 0 9 2 7 7 15 13 11 1 9 2
14 1 11 15 0 9 13 3 1 11 11 12 2 12 2
12 1 0 9 13 11 11 10 0 9 1 9 2
29 1 9 1 0 11 12 2 12 1 11 15 13 11 11 2 1 15 1 12 2 9 13 1 12 2 12 11 11 2
6 9 11 15 13 1 9
2 11 2
41 0 9 13 3 9 12 2 9 7 16 1 9 0 9 13 1 9 14 12 9 2 13 9 13 3 1 9 9 2 15 3 13 1 9 1 0 9 1 9 14 2
48 11 3 13 2 3 1 9 2 1 9 1 11 7 3 15 3 13 9 2 3 16 15 1 0 9 13 9 1 11 2 15 3 13 1 9 0 11 7 13 15 3 3 1 9 1 9 14 2
9 11 13 11 7 13 15 0 9 2
6 11 2 11 12 2 12
24 1 2 0 2 0 12 15 13 0 9 1 0 9 1 12 2 9 2 3 11 13 0 9 2
18 11 15 13 13 9 1 12 9 3 2 7 11 13 14 9 0 9 2
15 9 13 14 1 9 12 2 12 2 3 15 9 3 13 2
17 1 12 2 9 3 13 11 0 0 9 7 11 13 12 2 12 2
9 0 9 13 3 1 9 12 11 2
7 3 13 0 9 0 11 2
33 1 0 9 11 1 9 11 13 11 1 12 2 9 3 13 9 11 2 7 1 0 12 9 15 10 9 13 7 13 3 12 9 2
13 1 9 3 15 13 3 12 2 12 1 9 11 2
9 14 3 15 13 0 7 11 13 2
25 0 11 3 3 13 9 11 1 12 9 2 7 3 1 9 10 9 9 0 1 11 7 11 13 2
17 1 9 0 9 9 3 13 0 9 2 0 13 14 13 9 11 2
12 0 15 13 1 12 2 9 13 1 9 11 2
9 7 9 1 0 12 13 3 0 2
14 1 12 2 9 15 3 13 1 9 1 0 9 11 2
8 3 1 9 13 9 0 11 2
12 1 12 2 9 13 0 11 1 9 12 9 2
14 11 7 11 3 7 12 0 9 13 1 9 0 9 2
13 1 0 12 9 13 1 9 0 9 1 9 11 2
12 0 9 9 7 13 12 9 1 9 0 11 2
6 11 2 11 12 2 12
11 3 1 12 2 9 13 0 9 1 9 2
24 15 15 7 13 14 12 9 2 3 1 9 11 11 7 1 9 3 11 13 9 1 9 11 2
20 9 1 0 12 13 3 3 0 2 16 1 12 2 9 13 9 1 9 11 2
17 1 12 2 9 13 0 9 11 11 2 11 7 13 1 9 11 2
10 1 9 12 13 9 1 9 9 11 2
17 9 1 9 3 9 15 9 13 1 12 2 9 2 3 11 13 2
13 0 13 3 9 2 16 1 0 9 13 9 11 2
6 11 2 11 12 2 12
15 0 13 1 9 10 0 9 2 7 10 9 15 13 13 2
11 15 13 0 11 7 1 0 9 13 9 2
14 1 0 12 15 13 13 1 0 9 2 7 9 13 2
23 7 1 0 12 15 9 13 1 12 9 2 13 7 3 0 1 9 11 2 12 2 12 2
11 0 11 3 1 9 3 3 13 9 0 2
6 11 2 11 12 2 12
17 0 9 9 13 1 12 2 9 2 3 15 0 11 13 11 9 2
19 1 0 9 13 2 13 2 3 0 11 13 0 9 2 13 11 0 9 2
7 9 11 13 11 0 9 2
8 9 0 12 15 13 3 9 2
16 15 13 1 0 9 9 7 12 9 1 0 12 9 13 9 2
3 9 1 11
25 9 1 9 13 0 9 1 9 1 9 0 0 9 11 11 11 2 15 3 13 9 1 9 11 2
17 1 0 0 9 9 4 1 9 13 7 13 1 9 1 0 9 2
18 9 9 9 1 11 1 11 3 13 9 0 9 1 9 11 11 11 2
18 3 3 2 16 13 9 0 9 2 3 13 9 0 9 1 0 9 2
23 1 9 9 0 9 2 15 3 9 3 13 9 1 0 9 2 15 3 7 3 13 0 2
9 9 13 7 0 9 1 9 9 2
17 1 15 2 16 10 9 13 7 10 9 13 3 9 2 9 13 2
5 11 2 9 13 9
2 11 2
19 2 1 9 0 9 1 0 9 4 15 1 9 11 11 13 13 1 9 2
27 13 7 2 3 13 9 9 13 2 16 15 9 0 9 13 2 2 13 1 0 0 9 9 11 11 11 2
30 1 12 9 2 0 13 0 9 7 11 2 4 1 0 9 3 13 3 9 11 2 2 16 13 0 9 0 9 2 2
19 9 15 14 13 10 9 2 16 0 9 9 13 13 0 12 9 1 9 2
15 2 0 9 3 13 14 1 9 0 2 7 7 0 9 2
14 15 7 13 1 1 9 9 3 13 2 2 13 11 2
6 9 1 9 3 13 9
2 11 2
33 0 9 3 1 10 9 13 13 9 1 9 1 0 9 0 7 1 9 2 15 1 15 1 9 1 9 0 9 13 0 9 9 2
9 13 15 3 9 9 9 11 11 2
35 16 0 9 9 2 9 0 2 0 2 11 2 2 13 1 9 1 9 9 1 12 2 9 12 9 2 13 2 7 9 13 2 13 3 2
38 11 14 12 2 9 0 2 0 2 11 2 13 2 16 13 13 0 0 9 2 1 15 13 9 13 9 0 9 9 1 9 12 9 9 16 12 9 2
25 2 16 4 15 13 13 9 9 2 3 4 15 13 0 9 2 2 13 9 9 9 1 9 9 2
12 1 9 1 9 3 13 7 9 11 7 11 2
2 9 9
28 0 9 13 9 2 16 12 2 9 13 0 9 2 3 13 13 0 9 9 1 9 0 9 0 9 1 9 2
5 0 9 13 0 9
2 11 2
34 2 9 15 13 2 2 13 3 9 0 9 0 11 11 11 1 9 9 2 1 15 3 13 1 12 9 1 12 0 9 9 7 9 2
13 0 9 2 3 15 13 13 2 13 9 1 9 2
10 9 9 13 1 11 2 11 7 11 2
15 9 13 9 13 9 9 1 12 5 1 12 9 9 9 2
14 9 1 11 7 11 2 11 13 3 1 0 0 9 2
15 0 9 9 11 11 13 2 16 10 9 13 9 0 9 2
22 1 0 11 13 3 1 10 9 1 9 1 0 9 7 9 2 15 13 13 1 9 2
7 1 9 15 7 9 13 2
4 9 1 9 12
3 0 0 9
2 11 2
22 11 2 12 1 0 0 7 0 9 1 0 9 0 2 13 0 0 9 0 0 9 2
24 0 9 1 0 9 13 9 11 2 1 0 9 13 9 11 7 0 9 13 9 0 2 11 2
16 0 7 3 0 0 9 0 9 13 3 12 9 1 12 9 2
22 9 2 0 1 3 9 2 4 13 1 0 9 3 1 9 2 15 15 13 0 9 2
59 0 9 13 3 16 12 12 0 0 9 2 9 7 0 9 1 12 0 9 2 9 9 2 9 9 7 9 2 9 2 9 0 9 2 0 9 2 9 13 2 13 7 13 15 0 9 2 9 1 9 7 0 9 7 0 9 0 9 2
5 14 0 13 0 9
2 11 2
23 3 12 1 0 9 12 9 13 3 1 9 0 9 0 9 2 15 13 1 14 0 9 2
11 1 9 9 12 4 13 3 12 0 9 2
16 1 12 9 2 15 1 9 13 9 2 7 1 9 3 13 2
23 13 15 3 0 9 9 2 15 15 13 10 9 0 9 1 0 9 7 9 7 9 9 2
11 9 0 9 13 0 1 15 9 1 9 2
8 10 9 13 1 9 9 9 2
15 1 9 0 9 13 3 13 3 12 9 1 0 9 9 2
14 0 9 0 9 1 10 9 13 9 3 1 12 9 2
7 0 0 9 13 3 0 9
2 11 2
21 9 1 12 12 9 13 1 9 1 0 9 2 3 4 1 9 13 0 0 9 2
26 9 7 9 1 9 13 0 0 9 2 13 13 12 9 2 9 2 9 2 9 2 9 2 0 9 2
16 0 0 9 7 0 0 9 1 9 13 14 1 12 2 9 2
22 0 12 9 13 1 1 0 9 13 3 2 3 7 1 9 2 1 12 1 12 9 2
16 9 13 12 9 2 9 1 12 9 9 1 9 13 9 3 2
23 12 9 4 16 0 9 13 3 0 9 2 15 4 13 12 2 9 0 9 1 15 9 2
8 0 9 13 1 11 0 9 2
17 0 0 9 1 15 13 1 9 12 2 16 4 3 13 13 0 2
7 2 11 2 11 3 1 9
9 9 9 11 2 11 0 13 0 9
2 11 2
19 1 0 2 0 7 0 0 9 13 3 0 9 3 1 10 9 1 9 2
2 11 2
16 11 11 2 11 1 9 11 11 2 15 13 9 1 0 9 2
24 1 9 0 9 1 11 11 13 12 9 10 9 7 13 15 13 9 1 9 1 0 9 11 2
15 11 13 13 1 9 9 1 9 1 11 11 9 11 11 2
23 9 13 1 12 2 9 12 2 12 2 1 12 9 3 11 10 0 9 1 0 9 13 2
26 11 11 13 3 12 2 12 3 0 9 11 7 13 3 0 9 1 0 9 0 9 9 1 11 11 2
2 11 2
19 3 12 2 12 13 0 0 9 11 11 1 9 12 2 9 9 1 11 2
37 15 13 15 2 16 15 4 13 0 9 11 12 2 12 1 0 9 1 9 11 2 0 7 3 9 11 7 0 9 11 13 1 0 12 2 12 2
18 7 12 2 11 11 1 2 11 2 13 0 11 10 0 9 1 9 2
16 13 12 2 12 7 0 9 1 9 15 7 13 1 12 9 2
21 1 9 9 15 13 11 2 10 9 14 13 9 9 1 11 2 12 2 12 2 2
24 11 11 2 15 13 0 1 9 12 9 2 15 13 9 1 11 9 11 2 15 15 13 3 2
21 1 0 13 1 12 2 12 11 11 2 11 13 9 10 0 9 1 12 2 9 2
2 11 2
35 0 9 0 0 9 11 11 3 14 13 1 0 9 9 11 11 2 12 2 12 2 2 7 10 9 1 0 11 0 3 13 1 12 9 2
21 0 0 9 11 1 9 1 9 3 13 1 11 1 10 9 2 12 2 12 2 2
28 1 11 15 13 3 0 9 1 9 11 0 1 0 9 1 3 16 12 9 2 1 9 3 3 0 0 9 2
12 9 13 1 0 9 1 0 9 1 0 9 2
12 11 11 13 11 11 1 10 9 12 2 12 2
16 1 9 13 1 12 2 9 11 11 7 9 13 12 9 11 2
2 11 2
28 11 11 13 1 12 2 9 0 9 13 1 9 11 9 11 7 11 7 13 15 2 16 13 9 1 0 9 2
21 1 0 9 13 1 10 9 3 14 1 12 2 9 13 11 1 0 12 2 12 2
11 9 13 9 1 0 9 1 0 9 9 2
13 1 0 9 3 13 0 11 2 15 13 1 11 2
28 0 9 15 1 0 9 13 11 11 2 15 13 1 9 11 12 2 12 2 16 10 9 13 0 9 9 11 2
8 11 11 2 2 9 15 13 2
17 0 0 9 13 9 1 15 2 16 4 13 1 9 3 1 15 9
19 9 9 9 1 9 9 13 11 11 1 0 9 1 0 9 1 0 9 2
31 11 1 11 1 11 2 10 0 9 4 13 13 9 2 13 1 0 9 3 1 9 1 9 1 11 3 1 10 0 9 2
40 9 2 9 2 13 11 1 9 11 11 2 11 0 9 2 15 13 0 9 0 9 9 0 0 2 12 9 7 12 9 2 2 9 7 9 0 0 1 9 2
32 2 1 9 15 13 0 2 16 1 9 13 11 1 0 9 2 15 9 13 2 7 13 2 3 15 4 13 2 15 3 13 2
24 13 0 3 1 9 2 7 7 13 3 2 16 11 13 2 16 1 15 13 2 2 13 9 2
27 10 9 2 0 9 9 11 2 13 1 12 2 9 1 11 0 11 11 7 13 14 1 11 1 0 9 2
6 2 9 13 13 0 2
16 13 4 1 0 9 7 9 2 7 9 1 11 13 3 0 2
12 13 4 2 16 3 15 13 2 2 13 11 2
41 1 9 1 11 2 13 3 2 11 2 7 1 11 2 11 1 0 9 2 3 13 1 9 7 16 3 1 9 1 11 13 7 11 2 13 15 0 9 0 9 2
9 1 9 13 12 2 1 9 11 2
43 2 3 4 15 13 3 13 2 16 4 9 13 2 16 9 1 11 13 14 9 2 7 15 15 1 15 13 7 13 16 9 0 9 2 16 13 9 9 2 2 13 9 2
35 3 3 11 3 13 2 16 1 0 9 13 2 2 13 15 1 10 9 2 1 11 15 1 9 13 2 3 3 2 14 16 4 13 2 2
40 15 3 3 13 1 15 2 16 4 0 3 13 2 15 14 13 1 9 9 2 7 10 9 15 13 1 2 14 2 2 14 16 9 1 15 13 7 13 9 2
20 9 9 0 1 9 7 1 13 14 11 11 2 15 11 1 11 13 1 9 2
27 2 15 15 13 11 13 2 13 15 2 15 13 0 2 1 15 13 2 2 13 9 7 9 1 12 9 2
19 3 9 1 0 9 1 0 9 1 15 13 2 16 9 13 9 3 13 2
26 2 7 15 15 13 9 2 13 2 15 15 1 15 1 9 13 2 7 3 9 1 9 15 13 2 2
22 11 13 2 16 10 9 13 2 2 16 13 1 9 13 3 2 13 15 3 3 13 2
15 1 0 9 4 15 13 7 13 15 13 2 16 13 0 2
22 16 4 13 9 2 0 3 9 13 2 15 9 13 2 3 4 13 7 1 9 2 2
23 0 9 0 1 9 13 7 9 2 1 15 15 13 13 10 0 9 2 3 0 9 11 2
25 0 9 11 1 9 3 13 1 9 2 7 15 7 1 9 1 0 9 2 16 3 13 1 9 2
24 9 1 0 2 0 9 3 9 13 1 9 2 2 16 4 13 3 7 13 15 1 15 2 2
60 15 13 13 1 9 2 10 0 0 9 13 1 12 9 9 1 9 1 0 9 2 9 0 9 2 7 9 15 13 1 9 2 2 16 15 11 15 13 2 13 4 15 10 9 2 3 9 2 15 2 1 15 13 2 15 4 15 13 9 2
38 13 4 15 1 15 2 16 4 3 13 1 9 1 15 9 2 16 16 15 9 13 2 16 15 3 1 9 9 15 13 2 3 13 10 9 0 2 2
9 0 0 9 9 0 9 3 13 2
21 2 13 16 0 9 2 1 9 3 13 2 7 14 16 13 15 10 9 7 15 2
16 3 15 3 1 11 14 13 2 1 9 3 4 13 9 2 2
37 1 0 11 2 3 13 2 4 13 13 9 0 9 1 3 0 9 0 9 2 1 15 15 13 13 3 0 9 7 3 11 1 15 13 0 9 2
14 1 0 0 9 7 13 9 2 10 1 11 15 13 2
36 2 13 4 15 0 9 7 3 13 9 1 9 2 9 2 2 13 9 2 15 1 11 13 10 9 7 3 13 0 9 0 9 1 9 9 2
29 11 11 13 1 10 0 9 0 9 1 11 7 11 2 1 0 9 1 0 9 0 9 13 0 1 9 11 11 2
55 0 9 3 15 14 3 1 9 13 2 1 9 2 3 0 13 1 10 9 1 9 2 15 15 15 13 2 2 15 4 1 9 9 3 13 2 14 3 2 15 15 13 14 12 2 4 15 13 1 11 1 9 11 2 2
32 1 9 15 7 13 1 9 2 2 11 11 3 13 2 2 15 13 3 7 16 3 13 2 3 13 2 16 15 9 13 2 2
26 15 13 0 2 0 3 13 15 3 2 16 4 15 13 3 2 16 14 3 13 2 16 15 9 13 2
12 11 15 15 13 2 16 15 12 9 13 2 2
18 9 1 9 1 9 1 0 9 13 11 1 9 1 9 1 0 9 2
32 7 3 9 9 1 11 2 15 15 13 0 9 2 1 15 3 13 2 2 15 15 10 13 2 3 13 3 3 1 9 2 2
36 9 1 15 3 13 9 0 0 9 1 0 9 9 11 2 15 1 0 2 11 13 9 7 13 1 9 1 9 2 7 9 1 9 9 11 2
11 0 9 15 13 2 3 13 9 1 9 2
23 2 15 15 13 2 16 11 13 13 3 2 3 13 2 15 13 10 9 2 2 13 9 2
17 9 0 9 2 13 0 9 1 3 0 9 1 9 2 7 13 2
17 2 13 13 15 3 2 13 0 7 13 2 16 0 7 13 2 2
5 11 13 9 1 9
2 11 2
31 0 9 0 0 9 2 11 2 13 9 1 9 0 9 9 1 0 9 11 11 2 15 15 1 9 12 13 13 0 9 2
15 9 13 9 2 15 11 13 1 9 0 9 0 9 11 2
10 15 15 9 13 1 9 1 11 11 2
7 1 9 1 9 13 9 9
13 0 9 9 1 9 3 13 0 9 0 9 9 2
23 10 9 13 12 9 0 9 9 11 11 2 15 13 1 0 9 9 9 2 9 2 9 2
24 1 9 7 1 9 2 3 1 12 2 13 9 1 9 0 9 9 11 11 1 9 0 9 2
35 0 9 9 2 15 13 3 13 1 0 9 2 13 3 1 9 12 7 13 9 3 3 0 9 0 9 7 9 0 9 0 9 1 9 2
11 0 9 0 9 13 1 0 9 9 3 2
24 1 9 7 1 9 4 1 9 9 9 13 9 11 1 9 9 1 9 0 0 9 11 11 2
13 3 3 0 9 13 1 9 9 3 1 9 12 2
23 9 1 9 7 0 9 13 0 9 9 0 9 0 1 9 2 0 2 9 2 11 11 2
27 9 13 10 9 1 9 12 2 10 0 9 3 13 1 11 13 0 0 9 0 0 9 1 9 11 11 2
3 2 11 2
3 0 9 9
30 0 9 13 1 9 1 12 2 9 9 0 0 9 12 9 9 7 9 9 1 9 2 15 15 13 9 1 0 9 2
32 1 0 13 0 9 11 11 2 0 9 11 11 2 0 9 11 11 7 3 0 9 11 11 2 15 3 13 2 16 9 13 2
26 9 1 9 9 2 10 0 9 9 1 0 9 3 13 2 15 13 1 9 0 2 11 1 0 11 2
12 1 15 4 13 0 9 1 9 9 0 11 2
27 0 9 15 13 3 10 9 2 15 4 13 9 2 3 9 2 15 4 15 13 13 0 9 0 9 9 2
12 11 13 0 9 12 2 9 9 0 0 9 2
19 0 9 11 11 13 1 12 2 9 1 11 1 12 0 9 1 0 9 2
26 1 0 9 12 2 9 9 9 1 0 11 15 12 2 9 13 9 1 0 9 7 9 11 7 11 2
28 0 9 13 9 9 9 12 2 9 2 3 9 1 9 0 9 1 11 2 1 9 1 0 9 11 1 9 2
35 0 9 1 11 13 1 11 1 0 9 9 2 15 13 13 12 2 9 1 11 2 13 12 2 9 1 11 7 13 12 2 9 1 11 2
12 11 15 13 1 12 2 9 9 9 0 9 2
23 16 9 2 3 9 13 2 1 15 13 3 3 2 16 4 10 9 3 13 9 1 9 2
34 11 3 13 2 16 4 10 0 9 13 1 9 1 9 1 9 2 7 3 1 9 13 2 16 15 10 10 9 13 0 0 9 13 2
24 1 11 15 12 2 9 3 13 1 9 0 9 0 9 2 1 15 13 0 9 9 11 11 2
30 3 13 1 9 9 10 9 11 1 11 2 15 13 1 9 12 2 9 1 9 12 9 9 1 2 9 2 1 11 2
17 13 15 7 1 9 1 9 2 15 13 10 9 16 2 9 2 2
20 13 3 9 2 15 13 0 9 2 13 1 11 1 9 3 0 9 11 11 2
10 1 0 9 7 0 0 9 13 1 2
23 1 0 9 4 15 9 11 11 13 13 9 12 2 9 1 11 7 12 2 9 1 11 2
31 0 12 2 9 9 0 0 9 4 1 11 1 9 9 13 9 0 7 0 9 2 7 0 9 0 0 9 4 3 13 2
18 11 1 9 13 9 12 9 7 1 9 13 2 15 13 9 0 9 2
16 1 0 9 15 13 1 15 2 3 9 0 9 13 11 11 2
48 0 9 13 1 0 9 13 12 2 9 0 9 2 15 4 13 1 12 9 2 1 0 9 1 11 4 13 0 9 2 16 0 9 1 9 13 1 9 1 0 9 1 0 9 1 9 9 2
21 9 4 12 2 9 13 0 9 1 11 2 1 15 13 13 11 11 7 9 9 2
22 0 0 9 2 3 9 9 2 9 7 9 2 0 9 9 9 0 0 9 3 13 2
29 13 3 3 13 2 10 0 9 4 13 2 10 0 0 9 15 15 13 7 10 0 9 7 1 10 9 4 13 2
21 9 9 15 3 1 11 13 12 2 9 2 3 4 13 11 7 13 0 0 9 2
4 13 1 12 9
2 11 2
20 0 9 2 0 1 9 1 3 16 12 9 1 0 0 9 2 13 0 9 2
35 9 0 0 9 4 13 3 16 12 9 1 0 11 2 3 15 1 9 12 13 0 0 9 12 2 0 9 1 0 9 7 9 0 9 2
16 1 0 9 4 13 9 2 9 2 9 1 9 7 3 9 2
4 10 9 1 9
21 3 13 4 1 9 1 0 9 3 13 3 3 2 16 0 9 1 9 13 9 2
23 0 4 15 13 1 9 9 7 13 4 2 16 1 15 0 9 4 13 9 15 7 15 2
45 0 9 13 15 2 16 3 1 9 9 13 3 13 14 0 7 0 9 9 2 16 13 3 0 2 16 9 9 3 13 2 7 16 14 2 16 15 13 3 3 1 0 0 9 2
26 0 9 1 12 9 11 1 11 2 3 3 9 1 9 9 13 2 13 2 16 0 9 15 9 13 2
17 7 3 3 13 2 16 3 3 15 13 2 7 13 13 0 9 2
22 13 2 14 2 16 9 9 15 3 13 3 1 12 9 2 13 1 0 9 3 9 2
20 4 2 14 3 9 13 2 13 14 0 9 9 1 0 9 2 3 13 9 2
13 3 0 13 9 9 9 1 0 9 0 0 9 2
14 12 9 13 2 0 9 2 2 0 3 9 0 9 2
4 13 15 13 2
13 15 0 3 13 7 15 2 15 15 9 3 13 2
1 3
10 10 0 9 13 3 0 11 2 11 2
24 1 0 9 1 11 1 0 9 9 9 9 11 11 13 2 16 9 9 13 13 15 0 9 2
22 11 2 11 15 14 13 0 9 9 7 15 13 2 16 4 15 13 9 12 9 9 2
12 1 0 13 11 1 9 12 9 12 9 9 2
24 2 0 4 13 1 12 7 12 9 2 7 4 15 13 13 1 15 1 10 9 2 2 13 2
10 0 9 9 0 9 0 9 1 11 13
4 11 1 11 2
31 2 0 0 9 2 2 15 13 13 9 0 9 1 9 1 12 2 9 1 12 2 9 1 0 9 2 0 0 9 13 2
31 9 0 9 13 1 10 9 13 15 9 2 3 7 0 2 1 12 2 9 12 2 3 1 0 9 0 11 13 0 9 2
10 9 15 13 9 0 9 9 11 11 2
11 9 4 1 11 13 0 9 9 1 9 2
17 10 9 13 11 1 0 9 2 16 1 9 13 13 3 0 9 2
12 2 1 0 9 15 13 1 9 2 2 13 2
24 13 15 3 1 15 2 16 9 13 1 0 9 16 9 0 9 11 11 1 9 1 0 9 2
16 9 11 9 13 2 16 1 2 0 9 2 15 13 9 11 2
13 7 15 14 13 1 9 1 9 1 9 9 9 2
13 9 0 9 13 1 11 10 9 13 9 0 11 2
25 15 1 0 9 3 10 9 13 9 15 0 2 15 13 1 0 9 1 9 0 9 1 0 11 2
11 9 0 9 13 16 0 9 1 9 12 2
27 13 2 16 4 0 9 13 9 10 0 9 2 13 9 9 0 2 0 9 7 9 9 9 11 0 11 2
6 9 1 11 13 9 9
2 11 2
25 9 0 0 9 0 11 11 11 3 13 9 2 16 0 9 1 9 7 9 1 9 9 13 0 2
20 13 2 16 9 13 9 2 16 15 9 13 1 9 1 9 2 3 15 13 2
22 0 9 13 1 9 13 1 9 9 0 9 9 7 9 0 9 1 12 1 12 9 2
9 9 13 12 9 12 9 1 11 2
9 1 9 4 15 3 9 13 13 2
33 9 9 9 1 9 7 9 2 11 2 11 2 11 11 13 15 9 10 9 2 16 9 1 9 1 0 11 1 10 0 9 13 2
5 9 13 2 9 13
37 14 10 9 1 9 9 0 9 2 1 12 9 1 9 12 2 9 2 15 11 7 11 1 9 13 7 13 1 0 9 9 1 9 9 0 9 2
30 0 9 1 15 13 9 2 16 11 13 9 12 0 0 9 2 15 3 13 0 9 7 9 2 7 12 0 9 13 2
9 1 0 9 7 13 12 0 9 2
28 0 9 13 2 16 9 9 0 9 0 9 1 9 0 9 2 9 7 9 13 0 9 3 3 1 9 9 2
29 11 15 3 13 2 16 13 2 14 9 1 11 0 2 13 1 15 9 1 10 9 0 9 12 9 9 0 9 2
10 1 0 0 9 4 3 13 7 11 2
29 0 9 13 1 0 9 0 9 11 1 0 9 2 15 13 0 9 1 9 1 9 12 9 9 1 0 0 9 2
15 13 15 0 9 2 7 1 9 4 13 9 11 1 11 2
25 9 3 13 1 0 9 11 7 13 3 13 2 16 9 13 0 2 13 0 9 9 9 11 11 2
29 0 9 13 3 1 9 13 12 9 9 2 9 12 9 7 9 12 9 9 2 7 2 12 9 0 0 9 11 2
29 0 9 9 9 13 7 13 2 16 9 9 3 1 9 9 11 9 9 1 0 9 13 0 9 1 9 1 11 2
29 11 1 9 13 9 2 1 15 15 0 9 3 16 13 2 15 4 11 13 0 12 9 9 2 12 9 9 2 2
21 1 9 0 9 13 11 2 3 9 1 11 2 3 0 9 2 7 15 13 9 2
11 0 9 9 13 0 9 1 9 0 9 2
32 1 11 1 9 10 9 1 9 13 1 0 9 1 12 9 2 12 9 2 7 1 9 1 12 2 12 0 9 2 12 9 2
40 12 1 9 2 15 9 1 0 9 13 2 13 9 9 0 0 9 11 11 2 15 13 2 16 0 9 11 15 3 13 3 7 16 0 9 4 13 13 0 2
9 9 1 10 9 13 0 9 9 2
27 1 9 9 1 0 9 1 9 13 1 12 9 7 1 12 9 2 16 1 9 1 12 9 7 12 9 2
21 0 9 0 9 13 0 9 2 15 13 3 0 2 7 16 3 0 9 9 9 2
28 0 9 9 13 1 9 2 16 0 0 9 4 13 2 0 9 3 13 1 9 9 11 1 0 9 1 11 2
29 0 9 9 9 2 3 1 0 9 2 13 0 0 9 0 0 9 2 0 0 9 1 11 7 0 9 1 11 2
14 0 9 9 9 13 2 16 10 9 1 9 13 0 2
22 9 15 13 1 0 9 1 0 2 0 7 0 9 2 13 1 0 9 7 0 9 2
7 1 9 4 10 9 13 2
35 9 1 9 0 9 3 13 1 0 9 2 15 13 0 9 2 7 9 1 9 0 0 9 1 9 1 0 9 1 0 9 9 3 13 2
23 1 9 9 15 1 0 9 1 9 13 9 1 9 12 9 1 9 1 9 1 0 9 2
27 3 15 7 13 2 16 9 3 3 13 14 14 13 3 1 9 2 15 4 9 2 13 2 1 0 9 2
13 9 3 13 9 1 9 2 7 13 15 0 9 2
23 15 15 13 13 0 9 9 10 0 9 7 7 15 9 14 1 0 9 13 3 3 9 2
24 9 7 1 9 13 2 7 16 15 1 9 13 0 0 9 9 2 0 9 9 15 14 13 2
25 1 11 9 13 9 1 12 9 1 0 9 2 16 1 9 12 2 12 2 15 13 1 12 9 2
6 11 13 2 9 1 11
2 11 2
16 3 1 10 9 13 11 1 9 9 11 7 9 1 0 11 2
12 3 15 13 0 9 1 11 13 1 12 9 2
16 0 9 1 9 13 1 0 9 11 2 11 9 11 7 11 2
15 1 0 9 1 0 9 12 9 12 4 13 3 12 9 2
2 0 2
21 9 0 15 13 9 1 2 0 9 2 2 0 16 15 0 7 0 16 15 3 2
17 1 0 10 9 7 0 9 7 0 9 13 9 1 0 9 9 2
10 16 4 3 15 3 13 13 2 2 2
19 13 15 1 9 2 7 1 12 9 9 1 9 9 15 1 15 13 15 2
23 16 2 3 15 13 2 13 2 16 4 13 0 13 1 0 9 2 16 15 13 0 9 2
25 1 9 0 9 9 2 0 1 11 11 2 13 9 11 1 10 9 1 0 9 0 9 1 11 2
37 9 1 15 2 12 5 2 1 0 12 9 13 1 9 2 12 5 2 7 15 2 15 13 0 9 7 1 0 2 7 1 0 2 12 5 2 2
39 1 9 1 15 11 2 11 2 11 2 11 2 15 13 13 15 0 2 7 3 7 3 3 3 1 9 12 9 9 9 11 2 15 13 14 1 15 0 2
24 7 3 13 15 7 15 2 16 11 13 3 3 0 9 2 16 15 7 13 13 0 2 2 2
29 13 13 2 16 9 2 15 4 3 13 2 3 3 13 3 9 3 0 9 16 0 9 0 9 7 3 0 9 2
34 3 3 13 7 10 9 0 13 16 9 0 9 2 15 1 0 9 13 0 2 9 9 2 1 2 3 0 2 0 9 0 0 9 2
18 13 4 15 1 15 3 13 7 13 1 15 2 16 15 7 13 4 2
17 0 9 7 13 10 0 9 2 16 14 1 15 1 0 9 13 2
21 7 15 13 9 2 3 3 13 3 3 0 9 1 0 9 7 3 3 0 9 2
24 16 3 1 15 15 13 14 3 0 9 1 15 2 15 13 13 2 7 3 3 13 2 2 2
2 11 11
1 11
2 9 11
2 11 2
17 0 9 11 13 1 9 1 9 9 0 0 9 1 9 0 9 2
19 13 1 15 0 9 2 15 9 11 13 1 0 1 9 0 9 1 11 2
6 0 9 1 9 12 2
4 9 0 1 9
2 0 9
7 11 2 11 2 11 2 2
12 0 9 11 13 1 0 9 0 9 0 9 2
24 3 13 10 9 13 12 0 9 2 9 12 2 11 5 12 0 2 7 0 9 1 9 9 2
34 1 9 12 9 3 1 0 9 9 11 9 13 9 1 12 0 9 2 12 0 7 0 9 2 1 15 9 13 13 10 9 3 3 2
16 1 11 3 13 13 9 0 2 9 2 0 9 12 13 9 2
15 0 9 1 9 1 9 9 11 13 3 0 0 0 9 2
4 0 9 9 2
4 1 11 1 11
5 11 2 11 2 2
32 2 13 9 0 2 0 7 0 2 2 13 1 9 0 0 9 0 9 9 2 11 2 9 10 0 0 9 9 2 11 11 2
58 9 11 7 0 15 1 10 9 13 15 2 15 13 13 0 9 10 9 2 7 2 0 9 0 9 2 9 9 1 9 2 9 13 15 1 0 9 2 0 0 9 2 2 2 2 2 9 2 0 9 2 9 9 2 9 7 9 2
4 15 11 13 2
27 1 0 9 13 2 16 9 2 9 7 9 2 2 13 13 1 15 0 9 7 3 0 9 1 9 11 2
9 13 0 2 0 7 0 9 2 2
24 1 9 15 1 9 2 13 13 3 1 3 0 9 7 0 9 4 13 13 0 9 0 9 2
33 13 3 0 13 15 0 2 3 13 0 13 15 0 2 15 4 1 10 9 13 2 7 1 10 0 9 2 13 1 0 9 2 2
45 16 9 2 11 1 9 2 10 9 11 13 1 10 0 9 2 13 3 2 2 3 3 7 3 2 2 2 0 9 1 0 9 13 3 2 11 2 11 2 11 7 11 2 11 2
2 9 9
14 1 0 9 1 0 9 15 3 13 9 1 0 9 2
16 1 9 0 9 13 12 0 9 1 9 7 9 11 7 11 2
15 9 12 9 9 1 3 0 9 15 13 13 10 0 9 2
8 1 9 13 10 9 0 9 2
29 9 1 0 9 9 13 0 2 14 11 2 11 7 11 2 10 9 13 1 9 1 9 2 13 7 13 0 2 2
3 2 11 2
10 0 9 12 9 0 9 2 12 2 2
6 12 2 7 12 9 2
43 9 9 0 9 2 9 0 9 0 9 11 2 13 9 12 9 0 9 11 2 0 15 9 7 9 9 2 9 0 2 2 9 2 9 0 2 7 9 2 9 0 2 2
34 15 12 9 13 3 13 1 9 2 1 15 0 13 1 9 0 9 7 0 9 7 0 1 9 9 0 2 0 1 0 9 7 9 2
10 1 10 9 15 13 1 0 9 9 2
34 16 13 1 0 0 9 2 1 9 0 1 12 0 0 9 2 3 15 13 9 11 2 4 13 13 0 7 1 12 2 7 12 9 2
38 13 2 14 9 0 9 2 1 15 15 3 13 9 0 9 11 2 2 0 9 4 13 12 9 7 4 13 1 11 2 9 1 12 9 13 1 11 2
21 0 9 2 12 4 4 13 1 11 7 12 1 11 2 13 13 0 16 12 9 2
17 9 11 13 13 3 9 9 2 9 0 9 11 7 11 7 9 2
22 0 13 9 9 0 9 1 9 9 9 2 13 15 12 9 7 3 13 2 15 13 2
27 9 0 9 4 1 9 13 1 9 7 13 0 9 7 0 9 1 9 0 2 0 2 0 7 0 9 2
30 0 13 1 10 9 3 0 9 0 9 2 2 13 2 16 4 1 9 9 9 15 3 7 3 13 7 13 10 9 2
57 13 2 16 13 0 0 7 0 0 9 2 4 13 10 9 7 0 9 2 13 1 9 9 1 15 10 9 7 9 3 7 3 2 15 4 13 9 10 9 2 7 4 13 10 9 3 7 1 10 9 2 1 9 0 9 2 2
16 12 1 0 9 1 0 9 13 9 2 9 7 9 9 11 2
16 1 10 12 0 9 15 0 13 16 1 9 7 3 15 13 2
13 9 13 1 12 9 0 9 0 1 9 0 9 2
35 4 2 14 13 9 2 7 1 10 9 13 9 3 0 2 0 1 9 0 9 0 9 2 7 3 0 9 0 9 9 0 1 12 9 2
14 3 4 1 9 13 9 2 3 9 11 13 9 9 2
51 13 2 14 15 0 9 1 0 9 2 4 13 13 2 16 1 9 13 9 12 9 12 2 1 15 9 11 1 10 9 13 13 7 13 9 7 10 9 2 7 16 10 9 13 7 9 9 10 9 13 2
11 1 9 1 9 4 10 9 13 10 9 2
39 1 12 9 13 9 9 13 1 9 7 1 9 0 9 11 7 1 10 9 2 7 15 1 9 2 16 15 0 9 13 10 2 15 2 9 2 7 2 2
20 4 2 14 13 0 9 7 9 2 13 15 1 10 9 1 10 9 0 9 2
32 13 3 9 13 0 9 2 15 15 7 13 13 7 13 0 9 2 13 15 1 9 11 7 13 7 13 9 1 9 1 11 2
2 11 11
6 1 11 15 13 11 2
4 11 15 13 3
4 9 0 1 9
7 11 2 11 2 0 11 2
16 1 0 9 13 1 0 11 1 9 1 9 1 12 0 9 2
10 9 13 13 13 9 1 9 10 9 2
9 11 13 0 9 0 1 0 9 2
21 13 12 9 3 11 1 9 12 1 9 0 9 2 1 15 15 13 9 0 9 2
16 0 9 3 13 2 16 0 9 11 13 0 9 7 0 9 2
18 1 0 9 13 9 0 0 9 3 9 1 9 11 7 0 9 11 2
15 1 11 13 1 9 3 12 9 7 0 12 9 4 13 2
22 11 0 0 9 11 3 3 13 1 9 2 10 9 4 13 4 13 2 0 2 11 2
33 1 9 11 15 0 9 11 2 9 9 7 9 12 3 0 0 9 1 9 13 2 16 0 9 15 13 3 12 2 9 1 11 2
15 13 4 9 15 0 9 2 15 2 13 1 9 11 2 2
38 9 9 11 11 11 0 9 13 2 16 2 0 2 11 4 13 13 11 2 0 9 7 3 9 11 2 11 7 11 2 1 15 0 0 9 13 9 2
16 0 9 1 11 13 0 9 0 1 0 9 1 12 9 9 2
13 3 13 9 9 2 10 9 13 0 7 0 9 2
13 1 0 9 13 0 9 9 3 0 9 1 9 2
17 15 7 3 2 1 1 9 9 2 13 4 13 2 13 0 9 2
26 9 0 9 13 11 2 16 1 10 9 13 0 9 9 1 0 9 1 0 9 7 9 0 9 11 2
19 0 9 9 3 13 0 0 0 9 2 15 13 2 16 11 3 13 11 2
19 10 9 9 3 13 2 16 2 0 9 4 13 1 0 9 0 9 2 2
22 11 1 10 9 2 13 2 16 4 0 9 13 1 0 9 1 9 0 0 9 2 2
27 0 9 0 9 11 11 11 15 1 9 13 1 11 2 16 4 15 3 3 13 13 9 1 9 9 11 2
10 13 15 3 1 9 9 1 0 11 2
11 3 7 13 10 9 2 16 13 1 9 2
23 1 9 2 16 10 9 13 1 0 9 2 13 3 2 7 13 2 16 15 15 13 3 2
13 13 3 2 16 0 9 11 7 11 0 9 13 2
27 1 9 11 11 1 9 13 1 11 2 15 1 12 2 9 13 0 9 2 7 1 9 3 13 1 11 2
3 9 11 11
40 9 11 11 2 16 9 14 3 3 0 2 13 1 0 9 1 10 12 2 7 12 2 9 7 0 9 1 9 11 11 2 9 11 11 7 9 11 11 2 2
43 9 9 11 0 11 1 2 2 2 2 15 13 1 10 9 2 9 7 9 3 0 3 1 9 0 9 2 3 9 13 12 9 2 2 15 13 0 9 7 1 9 9 2
20 3 4 13 12 0 9 2 0 11 2 11 2 11 7 11 11 2 9 2 2
26 3 0 0 9 10 9 11 11 13 9 0 0 9 0 9 1 0 9 9 11 11 0 11 11 2 2
43 12 1 0 9 3 0 11 2 1 15 13 9 1 9 7 9 11 2 11 7 11 2 11 2 9 11 11 2 2 15 13 2 3 1 11 2 0 9 1 0 11 2 2
19 1 0 9 1 0 9 10 9 15 3 13 7 12 1 9 9 10 9 2
30 3 16 9 0 0 9 13 9 9 11 11 11 0 7 11 11 2 15 13 10 9 1 9 2 3 2 9 9 2 2
25 0 9 11 11 2 0 1 11 16 9 0 9 0 9 2 13 1 9 12 9 1 10 0 9 2
17 1 9 12 13 1 11 2 3 1 9 11 13 3 15 0 9 2
21 1 9 12 1 15 11 13 0 0 9 1 11 0 7 0 2 0 0 9 2 2
30 11 3 13 3 12 9 1 10 9 0 3 0 2 2 2 0 9 0 2 0 2 0 9 7 0 9 12 2 9 2
2 11 11
2 1 9
23 1 12 9 13 9 9 11 2 11 7 11 1 12 9 2 2 9 11 13 0 1 9 2
3 9 1 9
3 11 11 2
40 0 0 9 0 11 11 11 15 1 10 9 13 1 10 0 0 9 1 11 1 11 2 2 1 11 4 13 12 9 7 3 15 7 13 2 16 4 15 13 2
12 13 4 10 9 2 13 4 15 16 10 9 2
17 16 1 15 13 9 1 11 2 13 4 2 16 13 1 9 9 2
12 13 4 3 13 2 16 13 15 3 0 9 2
18 15 7 13 1 0 9 3 0 9 3 7 15 4 13 13 9 2 2
30 1 9 9 2 15 11 11 13 9 1 11 11 2 1 9 2 7 7 9 9 13 2 2 0 9 13 9 9 9 2
10 0 9 15 9 13 1 9 0 9 2
16 3 15 1 15 13 16 1 9 11 11 2 15 13 3 9 2
6 3 13 3 0 9 2
10 15 3 3 15 13 1 11 11 2 2
5 3 13 0 9 2
6 13 9 9 3 15 2
8 9 9 13 2 7 2 2 2
9 3 13 1 15 9 9 1 9 2
22 10 9 4 13 1 9 2 3 15 3 13 1 9 2 9 0 9 1 9 11 11 2
22 9 13 3 0 16 1 9 2 3 4 13 13 2 16 4 13 1 9 9 1 9 2
33 3 4 13 1 10 3 0 9 12 9 2 1 9 15 3 13 12 2 16 13 13 2 15 13 9 2 7 13 9 7 0 9 2
10 14 7 0 2 16 0 9 13 9 2
20 13 15 2 16 15 3 3 13 9 2 15 13 7 3 13 9 13 1 0 2
7 3 15 13 0 9 15 2
16 3 13 15 0 1 15 3 3 12 9 2 9 15 13 9 2
3 3 9 2
15 9 3 13 2 16 15 4 13 2 13 1 9 9 13 2
10 13 9 1 0 9 3 13 3 0 2
9 15 3 13 0 9 1 9 9 2
9 12 9 15 13 9 1 12 9 2
24 3 4 7 13 0 2 15 15 13 1 9 2 7 1 15 0 12 13 13 3 3 0 9 2
9 10 9 13 3 2 16 0 9 2
20 1 12 9 15 13 9 14 12 9 3 2 3 13 3 13 7 10 0 9 2
5 13 15 3 0 2
2 3 2
18 16 13 3 0 9 9 1 0 9 9 0 2 10 0 9 13 12 2
41 0 9 13 1 12 9 0 0 9 2 15 13 3 3 3 9 2 15 15 13 1 0 9 2 7 15 15 3 13 0 9 3 16 0 9 2 3 10 9 13 2
25 13 15 3 3 2 16 1 0 9 2 16 13 3 9 2 9 2 0 9 2 9 13 12 9 2
40 1 15 1 12 0 9 2 1 15 2 3 15 13 3 7 0 9 2 13 10 0 9 2 15 4 13 13 1 0 9 0 9 1 9 2 3 0 1 9 2
11 15 13 3 0 9 2 3 0 9 13 2
53 12 3 0 9 4 13 13 1 9 9 2 13 3 3 0 9 2 2 0 12 1 9 9 9 2 13 15 3 15 9 3 2 2 2 7 0 12 4 15 9 13 1 10 9 2 16 13 0 0 9 7 9 2
5 13 9 1 9 2
12 1 0 9 14 2 1 0 13 10 9 0 2
9 15 13 2 13 15 3 0 9 2
10 7 15 2 15 15 13 2 13 9 2
10 1 0 9 4 1 15 15 13 9 2
30 16 15 4 13 2 13 13 2 16 15 12 9 9 4 3 13 1 15 12 9 2 7 14 3 2 3 15 9 13 2
30 13 4 1 15 2 16 4 9 13 13 13 14 1 15 2 15 13 3 2 7 12 1 0 9 4 15 13 9 9 2
9 13 7 13 9 1 9 1 0 2
15 14 15 13 13 7 13 15 13 9 1 9 0 9 9 2
7 7 1 15 15 14 13 2
2 11 11
8 9 12 9 13 9 1 0 9
3 9 0 9
6 11 2 11 2 11 2
23 0 9 12 9 0 11 2 15 15 3 13 1 9 1 0 11 2 13 9 1 0 9 2
15 13 15 1 0 9 1 9 9 9 0 0 9 11 11 2
18 1 0 9 13 0 2 16 9 9 1 0 9 4 13 3 10 9 2
19 0 0 9 13 9 1 9 2 0 0 0 9 2 2 15 15 13 11 2
15 11 2 11 7 11 3 3 13 2 16 13 1 10 9 2
14 9 0 9 3 13 9 9 1 0 9 9 0 9 2
19 14 0 9 13 2 16 1 0 9 9 12 9 15 4 13 13 7 11 2
22 1 11 13 14 9 1 0 0 9 2 1 15 15 9 3 13 13 11 11 1 9 2
40 0 9 15 13 1 9 2 15 4 3 3 13 2 3 13 7 3 1 0 9 2 16 15 13 1 9 14 3 0 1 15 2 15 3 13 9 9 0 9 2
20 9 13 1 11 3 9 0 9 7 15 13 2 3 1 0 9 2 3 0 2
28 13 15 2 16 9 13 9 1 9 0 0 9 3 1 9 12 2 1 0 9 1 0 2 3 0 2 9 2
39 13 0 2 3 15 10 0 9 13 1 9 11 7 11 2 15 13 13 3 3 0 0 9 7 11 3 7 0 9 2 16 15 13 0 9 1 0 9 2
13 9 15 3 1 9 2 16 13 9 2 13 9 2
24 1 0 12 9 2 3 13 4 13 1 0 9 0 12 9 2 15 13 1 9 1 0 9 2
32 13 15 7 2 16 13 0 9 13 0 9 2 1 11 7 1 11 3 2 9 9 0 2 0 9 2 15 3 13 1 11 2
18 0 9 0 0 9 13 4 13 9 9 2 0 0 9 9 0 9 2
13 9 0 0 9 3 13 2 3 4 13 9 0 2
10 3 15 3 13 13 9 11 7 11 2
24 3 2 1 9 2 15 13 9 0 9 1 0 9 2 7 11 11 13 9 11 1 0 9 2
18 0 9 1 9 11 13 1 9 1 0 9 2 15 15 13 2 13 2
15 11 13 9 9 16 0 9 1 0 2 9 2 1 9 2
36 9 0 9 2 15 3 9 13 3 0 9 2 13 13 0 9 2 7 13 0 15 2 3 3 16 3 2 13 2 3 0 2 0 2 9 2
6 15 9 12 13 7 13
4 3 4 13 9
21 1 0 9 12 2 9 12 13 11 11 2 2 0 13 3 9 2 15 3 13 2
20 1 0 13 2 16 4 1 0 9 2 16 4 13 3 0 2 13 9 2 2
3 13 4 2
16 1 0 2 0 9 2 15 13 13 7 0 2 0 9 2 2
8 1 9 15 13 13 0 9 2
15 3 2 16 13 1 0 9 2 13 15 3 3 13 9 2
14 1 9 15 13 9 7 7 10 9 1 9 9 13 2
13 11 13 13 0 10 0 9 1 0 7 0 9 2
25 12 2 9 15 9 1 9 13 1 0 9 2 16 15 3 12 0 9 13 1 9 3 0 2 2
8 12 2 9 3 13 0 9 2
11 12 2 9 4 13 9 1 0 9 11 2
17 13 15 2 7 1 0 9 15 3 13 2 1 9 0 0 9 2
29 1 9 1 11 2 1 11 7 3 7 1 11 15 3 13 9 2 16 4 15 3 13 2 16 2 13 11 2 2
23 3 1 9 9 13 1 0 9 0 9 11 11 7 13 9 2 0 1 9 0 0 9 2
15 2 0 2 9 7 3 13 0 2 0 0 9 1 9 2
13 15 12 3 0 9 9 9 1 9 9 3 13 2
20 12 2 9 13 9 11 11 11 1 9 0 9 2 1 15 3 13 11 11 2
24 1 9 11 9 13 2 0 9 2 7 13 9 11 11 7 9 11 2 15 13 13 0 9 2
9 9 13 9 9 1 9 11 2 2
13 1 10 9 3 0 9 11 11 13 1 9 9 2
24 16 9 13 1 9 9 2 15 13 13 13 10 9 2 4 1 9 13 0 9 1 9 9 2
19 16 9 1 9 13 9 3 1 9 2 13 15 9 10 3 0 9 11 2
17 15 2 15 3 9 1 9 13 3 2 13 3 13 10 0 9 2
23 12 9 1 10 9 9 13 1 15 2 15 13 3 7 3 1 9 2 3 13 1 15 2
10 12 2 9 13 0 9 0 0 9 2
19 13 3 3 12 9 2 16 16 3 13 16 0 2 13 3 3 13 9 2
17 9 11 15 3 13 2 13 15 2 13 2 7 3 13 0 9 2
12 1 9 9 13 9 1 9 9 11 11 9 2
19 0 9 13 1 10 9 1 11 7 10 0 9 3 1 11 13 15 0 2
10 11 11 15 3 13 3 2 1 11 2
10 4 3 13 9 7 9 7 11 11 2
14 0 0 9 1 15 3 13 9 1 9 1 0 9 2
11 15 0 0 9 9 13 2 15 1 9 2
6 9 9 13 9 9 2
26 15 2 15 3 3 13 13 0 7 0 9 1 11 7 11 2 13 15 15 3 0 9 7 0 9 2
8 3 15 13 9 0 9 2 2
12 1 9 13 0 9 3 0 0 9 11 11 2
10 12 2 9 9 13 0 2 0 9 2
11 9 15 13 13 15 2 15 15 0 13 2
10 3 1 15 2 13 15 2 13 9 2
9 3 9 13 10 9 2 13 0 2
9 15 1 15 13 3 10 9 2 2
5 13 0 9 2 2
17 9 9 13 9 1 11 1 9 9 9 7 0 0 9 0 9 2
32 12 2 9 2 3 1 9 0 2 13 11 11 1 9 1 9 2 15 15 0 9 13 3 0 9 2 16 15 9 9 13 2
9 3 0 9 2 3 9 1 9 2
12 7 13 3 1 10 9 13 14 15 2 2 2
8 0 9 1 9 13 3 3 2
20 0 9 2 15 10 9 2 3 0 9 2 13 3 1 9 2 15 3 13 2
8 9 13 2 1 9 2 13 2
2 11 11
3 11 2 11
3 13 4 0
2 11 2
17 2 16 0 0 9 1 9 4 3 13 9 11 7 11 1 9 2
58 3 16 0 4 13 9 9 0 9 2 2 13 3 9 9 0 9 7 13 2 2 1 9 2 3 4 13 9 10 9 2 9 0 9 9 13 9 1 9 0 2 0 7 0 9 2 15 15 3 13 3 16 9 1 9 9 2 2
40 1 9 0 9 15 10 9 13 1 9 7 9 0 7 0 9 2 16 10 0 9 4 7 13 9 13 7 13 11 1 2 0 9 0 9 0 1 9 2 2
37 11 2 11 13 0 1 9 0 7 0 9 2 2 9 0 7 0 9 1 9 13 2 16 9 13 0 9 3 13 1 9 0 9 1 9 2 2
8 1 0 0 9 11 11 1 11
4 0 9 11 2
30 0 0 9 11 2 15 13 14 12 9 3 1 11 2 13 1 9 1 9 9 0 0 9 9 0 9 7 0 9 2
14 13 1 15 0 9 1 15 2 16 0 9 9 13 2
11 1 10 9 9 9 1 0 9 3 13 2
10 1 9 0 9 7 3 13 10 9 2
18 0 9 3 13 2 16 9 11 2 10 0 9 7 9 13 0 9 2
29 9 0 9 1 9 11 13 2 16 1 9 11 13 13 0 9 2 15 15 13 1 9 1 0 9 11 0 9 2
20 0 9 3 13 2 16 1 0 9 13 11 2 11 2 11 7 0 0 9 2
32 1 0 9 13 0 9 0 9 12 0 9 2 10 9 9 7 12 0 9 0 9 11 2 12 2 15 11 13 1 0 9 2
19 1 10 9 0 9 3 13 9 0 9 2 15 13 1 9 1 0 11 2
18 9 0 9 13 9 1 0 9 1 0 9 9 11 9 9 2 9 2
11 0 9 7 1 9 3 13 0 0 9 2
24 9 9 1 0 9 13 1 9 2 3 15 1 11 13 0 9 0 9 0 9 11 11 11 2
25 0 9 9 11 2 15 4 13 1 9 9 9 0 9 0 9 1 11 2 4 13 3 13 1 11
22 9 11 7 11 11 11 13 2 16 1 0 9 15 13 9 1 0 9 7 10 9 2
20 1 11 13 0 1 0 9 13 15 2 15 15 13 1 2 9 2 0 9 2
6 0 9 2 9 7 9
6 9 0 7 0 0 9
11 9 9 9 1 0 0 9 15 3 13 2
27 9 9 7 9 1 9 13 9 1 0 9 2 15 13 0 13 15 7 3 2 14 16 15 15 13 9 2
17 13 9 0 9 2 15 4 13 3 13 1 3 0 9 0 9 2
42 1 10 0 9 13 13 2 16 13 10 0 9 2 16 9 0 9 0 1 9 0 9 7 9 9 9 1 0 9 0 15 1 9 2 0 9 7 9 3 7 3 2
26 1 9 1 0 9 13 2 16 9 0 9 13 1 9 0 7 13 0 15 3 13 2 7 3 13 2
30 1 0 9 0 9 0 9 13 14 1 15 2 16 1 10 9 13 0 0 9 2 10 9 4 13 0 9 9 13 2
14 9 13 7 1 10 9 3 0 2 16 0 9 13 2
4 9 13 1 9
12 3 13 1 0 2 16 13 1 0 9 9 2
27 0 9 9 4 1 0 9 13 0 9 7 13 4 0 0 9 1 9 2 3 15 0 9 9 3 13 2
21 9 0 9 9 4 13 9 3 7 13 4 14 1 0 9 9 7 9 0 9 2
26 13 1 0 2 16 13 1 9 9 9 1 9 2 1 0 9 9 7 1 10 9 1 9 0 9 2
28 9 9 0 9 13 1 0 0 9 1 9 11 2 15 3 13 9 0 9 2 3 0 9 10 9 7 9 2
27 13 0 2 16 0 9 13 13 1 9 0 9 2 13 7 13 2 16 10 9 13 3 0 16 13 9 2
30 0 9 9 13 13 7 7 10 0 9 2 1 15 9 1 2 0 2 9 7 2 0 2 0 9 13 14 0 9 2
35 0 9 7 9 13 3 13 14 3 0 0 9 1 9 0 9 7 3 13 9 0 9 1 9 0 9 7 1 9 9 0 9 7 9 2
11 13 0 2 16 4 3 13 1 9 9 2
17 7 0 9 4 3 13 0 9 7 13 4 15 9 0 9 9 2
31 15 4 9 3 13 9 13 1 15 2 15 15 13 7 15 15 13 13 7 1 15 2 10 9 15 13 13 3 16 0 2
18 0 9 4 13 0 9 9 2 9 0 9 7 3 0 9 0 9 2
17 9 1 9 9 13 3 1 0 9 9 7 3 1 10 0 9 2
20 14 0 9 13 13 9 7 9 2 15 13 0 9 0 7 0 9 0 9 2
8 9 1 10 9 13 15 9 2
22 1 12 2 9 12 15 0 0 9 13 14 1 9 2 7 0 9 9 15 3 13 2
14 15 13 2 16 13 1 0 9 9 14 1 12 12 2
16 13 1 9 9 12 13 0 9 14 14 12 9 1 12 9 2
16 1 9 0 9 9 13 0 9 3 0 9 0 9 7 9 2
18 1 0 9 15 4 3 13 1 3 0 9 2 7 9 13 1 0 2
16 15 14 13 9 0 9 1 0 9 0 9 7 9 1 9 2
25 1 9 9 12 15 13 2 16 1 0 9 11 13 12 9 9 1 12 9 9 1 10 0 9 2
32 15 7 13 0 7 3 0 0 9 2 15 13 2 16 14 9 3 0 9 15 13 1 0 9 0 7 0 9 1 9 0 2
22 13 3 0 2 16 0 0 9 0 1 9 9 12 13 3 3 16 12 9 1 9 2
28 9 9 9 2 9 2 0 9 9 7 9 1 9 9 13 3 3 3 0 9 7 3 9 0 9 1 9 2
23 13 1 0 7 15 2 16 4 13 0 7 0 9 2 15 3 1 10 9 13 0 9 2
11 0 9 13 13 1 0 0 7 0 9 2
45 7 16 13 0 9 0 9 1 0 9 0 9 0 2 0 9 1 0 9 9 1 9 2 3 9 3 13 13 7 3 13 10 9 2 4 13 3 1 9 9 16 1 9 9 2
21 3 3 3 13 1 0 2 16 15 1 0 9 13 9 7 9 9 1 9 9 2
15 1 0 9 0 9 13 0 13 0 7 9 0 0 9 2
41 13 2 16 13 0 3 13 9 9 1 0 9 2 13 2 16 13 0 9 9 13 0 9 7 13 3 3 13 2 16 9 0 9 13 1 9 9 0 0 9 2
27 0 9 13 3 0 9 2 3 3 13 0 9 1 9 7 10 0 9 2 15 13 3 0 0 0 9 2
25 3 13 1 0 2 16 9 13 9 0 2 0 9 0 1 2 0 2 9 7 2 0 9 2 2
12 0 9 3 13 2 16 4 0 9 13 9 2
25 9 0 2 3 2 0 9 4 3 3 13 2 16 15 13 2 16 13 0 13 10 0 0 9 2
2 13 9
11 0 9 15 7 13 3 7 3 0 9 2
23 15 1 10 9 15 9 3 13 2 7 3 13 2 13 3 0 9 2 3 1 0 9 2
13 1 0 13 15 1 10 9 2 15 13 1 0 2
24 0 0 9 13 1 15 2 16 9 3 13 3 0 9 7 9 3 0 0 7 0 0 9 2
27 1 11 15 3 3 13 2 16 13 15 0 7 0 9 2 9 0 3 1 9 2 15 13 9 0 9 2
12 10 9 4 1 15 13 3 1 9 1 9 2
15 9 0 9 13 3 7 3 1 9 9 9 0 0 9 2
19 15 13 7 1 0 0 9 0 2 16 0 0 9 13 13 14 0 9 2
17 9 9 0 9 3 13 7 9 9 4 13 7 9 9 0 9 2
29 13 2 16 15 3 0 9 3 7 12 0 9 3 13 0 9 0 9 0 7 0 0 9 7 13 1 0 9 2
19 13 14 9 2 3 3 13 0 13 14 9 0 2 7 3 9 0 9 2
34 0 9 2 3 0 1 0 2 13 2 16 1 12 9 1 0 9 4 1 0 11 0 9 13 3 14 12 12 0 9 0 0 9 2
26 1 9 15 13 0 9 0 13 0 9 1 9 0 0 9 7 0 0 9 7 13 3 9 0 9 2
36 1 0 9 13 0 9 7 0 13 3 1 9 0 9 2 15 4 13 9 1 0 9 9 7 15 4 3 13 9 1 9 9 9 7 9 2
40 9 0 9 13 13 7 9 0 9 2 15 4 1 9 9 13 9 1 9 9 9 2 13 9 9 2 13 9 9 1 0 9 7 13 9 13 9 9 9 2
9 9 7 9 9 0 9 13 9 2
28 0 9 13 9 9 0 9 2 16 15 13 9 9 9 2 13 9 0 9 7 3 13 9 9 1 9 9 2
18 10 2 16 7 3 0 2 9 13 0 9 2 15 3 13 1 15 2
38 3 0 9 13 3 13 2 16 13 3 2 15 13 0 1 9 2 16 9 15 7 16 15 7 13 1 0 9 2 13 2 7 13 15 15 10 9 2
19 13 2 14 15 0 9 0 9 2 13 15 9 14 0 2 7 7 0 2
19 3 3 13 0 2 16 9 9 9 2 16 3 0 7 0 2 3 13 2
24 13 7 9 0 9 2 15 14 3 13 9 0 9 0 9 7 13 9 1 9 0 0 9 2
19 13 15 9 2 15 1 9 2 13 2 9 2 7 15 15 13 9 9 2
23 10 9 9 2 7 9 1 9 13 0 9 2 16 9 10 0 9 13 0 16 0 9 2
15 13 15 9 9 2 7 3 9 2 15 13 13 0 9 2
29 13 3 0 2 16 9 13 0 2 9 2 1 9 9 2 16 13 1 12 0 9 9 9 9 7 9 9 9 2
26 0 1 15 13 9 2 15 3 2 16 4 15 1 10 0 9 13 2 13 0 9 0 1 0 9 2
23 9 7 9 10 9 15 3 9 9 7 9 3 13 1 0 9 7 13 7 10 9 9 2
27 13 15 3 9 2 7 3 3 0 9 7 9 9 2 15 13 9 0 9 9 7 9 2 0 2 9 2
2 0 9
15 1 0 9 13 0 9 9 2 9 7 9 1 0 9 2
33 1 12 9 15 3 13 2 16 9 0 9 1 9 10 0 9 4 13 3 15 2 16 13 1 0 9 0 0 9 7 0 9 2
28 1 0 9 15 7 3 13 9 1 0 2 7 3 1 0 0 9 2 16 4 10 0 9 13 13 10 9 2
15 10 1 9 0 9 1 0 9 15 3 13 1 9 0 2
27 15 15 13 3 1 9 1 9 0 2 15 13 1 9 0 0 9 2 1 15 13 1 11 13 0 9 2
20 0 9 13 15 13 2 15 13 0 14 1 0 9 2 7 7 1 0 9 2
22 1 15 9 1 15 4 13 14 0 9 7 9 0 9 2 7 10 0 3 0 9 2
33 0 9 13 0 0 9 1 0 9 2 13 9 1 0 9 2 13 10 9 0 9 1 9 7 13 1 0 9 0 9 7 9 2
14 15 13 3 0 2 10 0 9 13 0 9 13 3 2
19 1 15 0 9 0 9 13 3 13 0 9 7 15 13 1 9 9 9 2
28 9 2 16 1 0 9 7 0 9 4 1 0 9 0 9 13 0 0 0 9 1 12 9 2 13 3 0 2
36 1 15 2 16 15 1 15 0 9 13 3 3 2 3 15 13 2 13 2 16 7 1 0 9 13 0 9 1 0 9 3 0 16 9 3 2
9 0 9 13 1 15 3 0 9 2
23 7 3 3 14 15 15 2 15 15 1 11 13 1 9 2 15 16 9 13 9 1 9 2
19 13 7 2 16 4 0 9 3 13 13 3 15 7 16 4 13 10 9 2
5 15 4 15 13 2
20 0 9 4 13 13 0 9 2 9 7 9 7 13 9 1 9 10 0 9 2
36 3 3 4 14 13 2 16 4 4 13 15 9 2 13 9 7 3 13 9 2 13 15 12 9 15 9 2 9 2 9 7 0 9 0 9 2
12 3 4 15 13 13 3 2 16 1 12 9 2
30 7 3 1 10 9 4 0 9 13 13 1 0 9 2 16 4 13 0 9 0 9 1 0 9 0 9 7 9 9 2
19 10 9 4 13 14 3 3 2 16 4 9 9 13 0 9 1 11 0 2
55 13 7 1 3 0 2 16 15 1 0 9 13 9 2 16 3 9 0 9 1 0 9 0 9 2 9 0 9 1 0 9 10 0 9 2 0 2 0 9 2 2 9 9 1 9 9 7 3 9 9 0 9 1 11 2
27 1 0 9 2 3 13 0 9 1 0 0 9 3 0 7 3 0 2 13 0 15 3 3 13 7 13 2
14 0 9 10 9 13 3 0 0 9 1 9 0 9 2
3 9 0 9
18 1 0 9 0 0 9 13 0 9 9 0 2 0 7 3 0 9 2
51 9 2 9 2 9 0 9 2 9 0 9 2 9 0 9 2 9 0 7 0 9 2 9 2 9 9 7 0 0 9 9 2 15 15 13 2 16 4 0 9 13 0 13 0 9 0 9 1 0 9 2
17 0 9 0 9 3 13 2 16 4 0 9 10 9 13 3 0 2
25 3 0 0 9 2 15 3 1 0 2 9 13 2 13 0 9 0 9 2 9 2 9 7 9 2
15 1 9 10 0 9 4 13 3 0 13 1 10 0 9 2
13 11 13 3 0 9 13 15 3 1 0 0 9 2
13 13 7 12 2 10 0 9 15 1 10 9 13 2
39 0 9 13 10 0 9 10 9 2 13 7 13 1 15 2 16 4 15 0 9 9 7 9 0 9 13 1 0 9 7 13 3 3 0 0 9 0 9 2
18 9 10 9 13 2 16 4 15 13 9 1 9 9 0 9 1 11 2
21 9 2 1 15 4 1 0 9 13 1 0 0 9 2 0 0 9 7 0 9 2
28 10 9 13 15 0 13 3 0 9 9 0 10 0 9 2 9 7 0 9 7 13 1 15 10 0 0 9 2
10 1 9 15 13 0 9 0 0 9 2
4 9 1 9 9
19 9 15 13 2 16 13 1 9 9 3 3 2 16 0 9 3 15 13 2
25 9 0 9 15 13 2 16 16 15 13 9 15 13 1 9 2 15 2 12 9 1 9 2 3 2
32 15 2 15 13 13 1 0 9 1 9 2 15 13 3 7 13 15 10 0 9 2 15 0 13 2 16 9 15 13 3 3 2
6 13 15 13 15 0 2
3 1 9 2
16 9 12 13 3 10 9 1 9 0 2 3 15 15 3 13 2
5 13 1 9 9 2
8 15 1 9 3 2 0 1 9
27 12 2 9 13 0 0 9 9 9 9 2 12 1 9 12 7 1 9 3 9 1 0 0 9 7 9 2
9 0 9 0 9 13 15 1 9 2
14 2 9 2 4 13 1 9 2 16 13 15 14 9 2
7 3 7 13 9 1 9 2
16 0 7 0 0 9 1 15 4 13 2 16 15 13 3 0 2
9 0 12 0 9 13 11 3 3 2
36 3 13 2 16 15 13 9 9 10 0 9 2 7 0 0 9 1 9 9 1 0 9 7 9 11 2 15 13 9 1 9 3 1 0 9 2
26 13 15 1 0 9 2 16 13 15 2 16 2 0 2 0 9 13 3 3 13 1 9 9 0 9 2
26 9 13 3 0 9 2 3 13 9 9 2 13 0 9 0 9 7 13 0 0 9 3 13 7 13 2
8 15 15 13 13 12 2 9 2
17 1 0 9 1 9 15 7 9 13 9 1 9 9 1 9 9 2
39 1 0 9 2 1 9 3 0 9 9 7 0 9 2 1 0 9 13 3 0 9 9 2 0 2 9 2 2 2 1 9 0 9 2 7 0 9 9 2
8 9 4 9 13 0 0 9 2
12 15 13 15 2 15 13 0 1 0 9 9 2
14 0 9 2 15 15 13 0 0 9 2 13 0 9 2
44 10 9 13 1 15 9 2 1 0 9 3 13 1 0 0 9 7 10 9 0 3 9 0 7 0 2 0 1 15 2 16 0 9 15 4 13 13 3 1 9 9 1 9 2
13 3 2 0 9 4 13 3 3 0 9 0 9 2
18 0 0 9 2 15 13 1 9 9 3 0 2 4 13 1 0 9 2
79 3 15 4 13 7 1 9 9 2 15 13 4 13 1 12 9 2 12 2 0 9 4 3 13 9 2 12 2 9 0 1 9 0 9 7 0 15 1 3 0 9 4 13 14 1 0 0 9 2 12 2 9 2 15 13 1 0 9 2 7 13 1 10 9 0 2 4 9 3 13 15 2 12 2 9 0 3 9 2
25 1 0 9 3 13 1 9 1 9 2 9 9 1 0 0 9 7 3 7 1 9 1 0 9 2
14 1 0 9 4 10 9 13 3 9 0 9 1 9 2
26 1 9 12 1 9 0 9 15 13 1 12 5 9 1 9 1 0 9 2 16 0 12 5 13 9 2
34 10 9 13 3 0 2 16 13 10 0 0 9 1 0 9 2 1 0 9 13 3 13 2 16 15 2 15 13 2 13 3 1 9 2
20 1 9 2 0 2 9 0 9 2 9 1 0 9 7 9 13 0 9 9 2
4 9 13 0 2
21 9 2 13 0 9 1 9 9 1 10 2 15 13 0 9 2 3 3 0 9 2
9 13 13 7 9 0 3 15 13 2
58 9 2 1 15 9 15 13 9 2 9 2 3 1 0 9 9 2 15 4 3 13 3 0 7 13 13 2 16 4 15 13 0 9 13 1 0 2 1 11 13 0 0 9 9 0 9 2 16 1 0 9 15 13 12 5 9 2 2
16 0 9 3 13 9 9 2 3 2 0 2 13 2 0 2 2
27 1 9 13 2 16 9 4 1 9 13 3 1 0 2 3 1 0 0 9 2 15 4 13 9 1 9 2
19 1 15 4 13 9 0 9 2 15 10 9 13 7 4 13 3 1 0 2
10 13 15 2 16 15 13 1 12 5 2
48 10 9 4 13 3 0 9 2 15 15 4 3 13 7 9 1 0 0 9 2 15 13 3 2 1 0 7 3 0 9 2 16 15 1 10 9 13 2 13 4 7 13 1 0 0 9 2 2
30 0 9 15 13 2 1 0 9 13 10 9 14 0 1 9 1 0 9 1 0 9 9 2 9 2 9 2 9 3 2
6 9 9 7 0 9 9
8 9 13 14 0 9 9 9 2
9 0 9 3 3 13 1 0 9 2
45 9 9 9 1 9 0 9 1 0 0 9 3 11 13 7 16 4 9 1 9 0 9 13 2 13 0 0 9 2 1 9 9 1 0 9 7 9 1 0 9 2 3 1 9 2
11 11 3 13 13 9 0 9 1 10 9 2
21 9 0 9 13 3 3 0 9 1 0 9 1 9 2 9 1 9 1 9 2 2
6 3 13 10 10 9 2
28 9 9 0 9 3 2 3 15 13 9 2 13 3 0 7 13 15 1 9 1 12 1 12 9 12 0 9 2
26 1 0 9 13 7 0 2 16 9 9 13 1 9 1 0 9 3 1 15 2 3 1 9 0 9 2
20 1 0 0 9 13 1 3 0 9 3 1 9 2 9 0 9 2 0 9 2
15 0 9 13 3 3 10 9 3 1 9 2 9 7 9 2
36 12 5 9 7 12 5 0 0 9 2 9 2 13 1 9 0 9 9 1 9 2 7 12 5 2 12 5 9 2 9 0 9 0 9 13 2
17 12 5 9 7 12 5 9 13 3 9 9 9 1 0 0 9 2
19 3 12 12 9 13 2 3 0 13 0 9 1 0 9 9 1 0 9 2
16 9 7 9 15 3 3 13 1 0 9 2 16 13 9 9 2
12 14 9 7 9 15 13 2 16 13 3 13 2
21 3 13 2 16 15 0 9 2 15 0 9 1 9 7 15 3 0 9 9 9 2
5 0 13 0 9 2
13 3 15 1 9 0 9 13 9 2 12 5 2 2
26 1 12 9 15 3 13 9 9 1 9 7 9 2 1 0 9 7 0 9 1 9 1 9 1 9 2
49 3 0 13 9 2 16 9 13 0 9 1 0 9 9 2 12 5 2 2 1 0 9 0 9 2 12 5 2 2 1 9 15 9 2 12 5 2 7 1 9 3 13 9 9 2 12 5 2 2
38 0 9 9 7 0 9 9 13 1 0 2 16 4 15 2 15 1 15 13 2 15 13 13 0 0 9 7 16 4 13 0 3 13 1 0 0 9 2
12 3 13 0 9 1 9 1 9 16 1 9 2
8 0 9 1 9 13 3 0 2
12 9 13 3 9 1 9 2 9 7 0 9 2
11 3 1 9 9 13 9 2 12 5 2 2
12 1 0 9 13 12 5 9 7 12 5 9 2
23 9 13 15 0 9 2 1 0 3 9 2 3 9 2 15 7 3 13 9 0 9 2 2
20 3 15 13 7 0 7 0 9 13 13 3 1 9 12 9 3 16 0 9 2
15 12 5 13 2 16 4 13 1 0 2 1 9 1 9 2
34 0 9 15 13 9 13 7 3 13 2 3 9 13 0 9 13 9 7 0 9 2 12 5 15 13 2 16 10 9 13 1 0 9 2
15 9 13 1 9 1 9 3 0 7 13 7 9 1 9 2
11 13 1 9 2 7 9 3 4 13 0 9
18 11 11 2 0 9 9 9 11 2 2 0 9 0 9 13 13 9 2
24 9 9 2 3 16 0 9 7 0 9 2 13 13 9 7 3 13 7 13 1 9 9 9 2
28 0 9 0 9 1 10 9 15 7 13 2 16 1 0 9 2 1 9 7 9 2 1 9 0 9 0 9 2
18 4 13 9 2 13 11 2 0 0 9 13 1 9 2 3 3 9 2
49 3 15 13 2 16 4 9 13 1 9 1 9 2 3 4 15 13 9 2 3 15 13 9 1 9 2 3 13 9 2 7 2 13 9 7 13 3 2 2 16 15 0 13 1 10 0 9 0 2
9 9 9 13 7 1 0 9 13 2
28 1 0 7 0 9 4 13 9 12 0 9 1 12 9 1 0 9 7 13 15 9 9 1 12 2 12 5 2
30 0 9 9 4 15 13 13 1 0 12 9 1 12 9 1 0 9 2 15 13 4 13 14 1 12 9 1 0 9 2
10 1 0 9 4 9 13 9 0 9 2
14 9 1 0 9 13 0 2 7 11 15 4 13 2 2
24 11 11 2 9 0 9 0 9 7 9 11 2 2 9 4 7 1 9 12 13 1 0 9 2
25 1 15 13 0 9 9 9 0 9 0 1 9 2 15 15 3 13 1 9 1 0 7 0 9 2
19 9 12 13 1 9 0 9 9 0 2 3 15 9 13 1 10 0 9 2
21 9 3 4 13 1 0 9 0 9 16 3 2 15 7 0 9 13 1 0 9 2
18 13 15 9 0 0 9 1 0 9 9 2 15 4 9 3 3 13 2
18 1 0 9 13 9 0 9 9 1 9 9 1 9 0 9 7 9 2
10 13 15 1 15 9 2 9 15 2 2
18 10 15 13 9 1 9 7 13 1 9 0 7 0 9 1 0 9 2
10 3 9 13 0 9 2 7 0 9 2
20 1 9 0 7 0 9 7 1 9 9 7 9 13 9 1 0 9 13 2 2
30 11 11 2 9 9 1 0 9 7 9 11 2 2 0 11 1 9 11 13 1 10 9 7 1 9 3 13 10 9 2
28 13 15 2 16 12 9 0 9 1 15 13 0 9 2 7 3 13 10 0 9 1 0 9 0 9 13 0 2
39 13 14 9 0 0 7 0 9 0 7 0 9 2 7 15 3 0 9 1 0 9 2 13 7 0 9 9 9 7 9 2 16 15 0 13 13 14 3 2
24 9 13 3 10 2 0 9 13 0 2 9 13 0 2 1 9 13 13 0 0 9 7 0 2
22 9 4 1 0 9 13 1 0 9 9 2 0 9 2 1 0 9 2 1 0 9 2
17 3 15 15 9 13 2 16 1 9 1 9 9 4 13 9 3 2
6 14 2 15 15 13 2
13 10 9 3 0 13 7 13 4 14 0 9 2 2
2 11 11
17 9 13 15 9 11 1 12 12 9 2 9 7 9 7 15 9 2
15 13 2 13 2 0 15 2 10 9 15 1 0 9 13 2
27 1 0 9 12 13 15 9 7 9 11 3 9 2 9 1 9 2 0 9 1 9 2 9 7 0 9 2
5 9 13 14 0 12
2 3 3
2 11 2
15 9 9 9 9 7 13 1 9 1 9 9 12 2 9 2
12 14 1 0 9 15 0 2 9 13 0 9 2
17 7 1 9 0 9 13 9 3 1 9 7 9 13 14 0 12 2
6 11 2 11 12 2 12
21 3 1 0 9 15 1 9 1 0 9 13 15 12 9 2 11 2 11 7 11 2
12 7 0 9 13 1 9 0 9 2 14 0 2
14 1 0 9 15 13 3 12 2 7 0 9 3 13 2
21 1 12 9 15 0 9 13 3 0 9 1 9 11 2 1 9 1 11 7 11 2
17 3 0 9 13 0 9 9 7 13 15 10 9 2 15 13 9 2
45 3 15 1 15 13 7 0 9 2 7 3 0 9 9 11 1 9 0 9 1 11 7 0 9 1 11 3 13 14 9 2 16 1 0 9 15 0 2 0 9 13 3 0 9 2
16 13 1 9 2 16 1 9 13 12 9 2 11 7 11 2 2
15 3 15 3 13 3 9 11 2 15 13 3 9 1 11 2
2 11 2
15 1 0 0 12 15 9 13 1 9 7 13 15 0 9 2
3 11 1 11
26 2 9 15 1 0 9 11 1 11 1 11 13 2 7 1 11 3 13 9 2 0 15 0 0 9 2
9 13 14 1 9 2 3 15 13 2
17 13 15 7 1 9 1 9 10 9 1 11 2 3 3 9 13 2
23 3 3 13 9 9 7 0 9 13 2 2 13 15 3 3 1 9 9 0 9 11 11 2
14 0 9 12 9 13 2 13 15 7 1 12 9 9 2
21 7 16 9 0 11 2 11 13 2 2 9 13 1 15 0 2 16 12 9 2 2
10 3 15 3 13 1 0 9 2 2 2
26 11 15 3 13 1 9 11 1 11 2 1 9 1 11 15 13 9 11 2 16 1 11 3 13 11 2
18 9 11 13 3 12 0 9 2 11 7 13 1 10 9 7 1 9 2
3 2 11 2
3 15 1 9
2 11 2
26 9 2 15 1 9 13 0 9 2 4 13 9 0 9 2 9 0 15 0 9 1 0 16 0 9 2
30 0 0 9 2 13 15 2 16 15 13 1 9 2 4 13 3 16 9 9 0 9 11 7 13 4 9 9 7 9 2
29 9 0 9 4 15 13 13 15 9 7 9 2 15 0 9 13 1 10 9 2 7 2 9 2 9 2 9 3 2
2 0 9
5 11 2 11 2 2
19 1 0 9 9 7 9 15 1 0 2 0 9 2 3 13 0 0 9 2
29 3 2 0 9 2 2 9 12 9 11 1 9 0 7 0 1 0 9 2 13 13 2 16 15 13 15 0 9 2
18 0 9 15 13 1 12 9 2 1 0 13 9 1 12 1 12 9 2
24 9 15 13 1 9 9 2 0 9 11 2 11 1 2 0 9 2 2 9 9 1 0 9 2
10 0 9 1 15 13 0 9 12 9 2
17 0 9 13 9 0 9 11 2 15 0 9 13 1 12 9 9 2
15 3 1 9 11 1 0 9 9 13 0 9 2 12 9 2
17 12 9 1 11 7 3 13 9 0 9 1 9 9 2 13 12 2
6 9 0 1 9 1 9
4 11 2 11 2
28 9 0 0 9 2 11 2 11 11 3 13 2 16 13 9 2 3 13 0 0 9 1 11 1 0 7 0 2
30 10 9 13 1 9 1 9 11 1 11 7 9 0 0 9 2 11 2 11 11 2 15 13 1 9 9 1 12 9 2
22 1 9 1 10 0 9 2 0 0 9 2 13 0 9 3 0 2 13 3 9 11 2
25 1 9 2 3 1 0 9 1 0 12 9 13 12 9 2 9 9 0 9 1 9 13 14 12 2
4 9 1 0 9
5 9 9 3 3 13
5 11 2 11 2 2
26 9 1 0 9 0 9 11 2 11 4 3 13 0 9 1 11 7 11 2 16 13 0 13 0 9 2
14 0 9 15 3 1 9 9 1 11 14 13 1 9 2
19 13 15 3 9 9 1 11 11 11 1 15 2 16 9 13 3 14 9 2
25 2 13 15 7 3 2 16 9 1 0 9 9 13 1 9 11 1 10 0 9 2 2 13 11 2
32 13 15 1 9 9 2 16 3 13 0 9 9 2 16 4 3 13 9 11 9 0 11 9 2 7 13 1 10 0 9 9 2
19 2 1 15 15 13 13 2 16 1 10 9 7 9 9 13 15 1 9 2
17 13 15 13 2 1 10 0 9 4 13 9 13 2 2 13 11 2
16 9 13 9 9 14 1 15 2 16 1 10 9 3 13 9 2
24 3 15 7 1 11 1 0 9 13 9 1 9 0 9 2 16 11 14 0 9 16 0 13 2
7 1 9 14 9 9 1 9
2 11 2
37 16 4 9 9 13 13 1 0 9 1 0 9 11 7 11 7 10 9 1 9 13 9 9 2 4 13 1 0 9 13 0 9 12 9 1 9 2
33 3 15 13 9 9 0 9 11 9 1 15 2 16 10 1 15 0 9 13 0 9 2 3 7 9 2 1 0 9 1 9 9 2
17 9 3 13 2 16 1 9 13 3 0 9 9 1 0 0 9 2
32 1 0 9 9 0 9 9 11 11 13 2 16 1 0 9 4 9 1 0 9 1 0 0 9 1 9 0 9 13 0 9 2
7 15 9 13 9 9 9 2
11 9 2 15 13 1 0 9 2 4 13 2
17 16 15 9 13 7 13 15 0 9 2 13 15 0 9 13 3 2
11 9 4 13 1 9 10 7 0 9 1 9
5 11 2 11 2 2
25 9 0 9 15 4 13 9 1 11 7 1 10 9 4 13 9 9 0 9 0 9 3 1 15 2
11 9 4 13 1 10 9 3 13 0 9 2
12 13 15 9 2 15 3 1 9 9 13 9 2
26 1 9 15 1 9 0 12 9 13 9 0 9 13 1 9 3 12 9 7 1 0 9 1 12 9 2
35 1 9 11 13 9 1 9 0 0 9 13 12 9 2 0 9 0 9 13 13 0 16 12 9 1 12 9 2 1 10 9 7 12 9 2
20 9 13 1 15 2 16 0 9 13 13 3 1 9 1 9 9 9 1 9 2
23 9 11 11 2 11 13 2 16 9 13 9 9 2 15 13 9 9 1 9 1 9 9 2
36 9 9 1 9 1 9 9 11 2 11 2 11 2 11 2 13 2 16 2 9 13 14 1 15 9 2 16 4 13 4 13 1 9 9 2 2
13 0 9 13 13 16 9 0 9 7 9 0 9 2
15 7 3 7 9 4 13 1 9 10 9 1 0 0 9 2
3 11 13 9
5 11 2 11 2 2
16 0 7 0 9 2 11 2 13 15 9 1 9 12 0 9 2
12 1 12 0 9 11 3 1 9 13 12 9 2
8 13 1 15 0 0 9 9 2
25 9 1 9 13 9 2 15 13 9 9 11 9 12 2 12 2 12 2 9 4 13 12 2 9 2
9 0 9 11 13 3 12 9 9 2
15 0 9 9 13 12 9 9 2 1 15 12 13 0 9 2
8 0 9 1 9 13 12 9 2
22 0 9 3 3 2 13 9 12 0 9 2 0 2 0 9 2 1 9 9 0 9 2
12 0 9 13 9 9 3 12 9 1 10 9 2
26 10 9 13 1 0 9 13 12 9 0 9 2 13 0 0 9 7 9 9 1 9 1 0 9 9 2
5 11 1 9 0 9
4 11 2 11 2
35 0 0 9 3 13 2 16 9 13 0 9 2 16 4 13 9 1 0 0 9 1 0 7 0 11 2 1 15 1 0 9 13 9 9 2
15 9 9 9 9 13 2 16 9 0 9 13 9 0 9 2
30 9 1 0 9 0 9 11 11 11 7 0 9 0 10 9 11 11 11 13 1 9 3 3 1 11 3 0 9 11 2
21 9 11 3 13 1 9 9 7 13 9 2 16 4 15 2 13 13 1 9 2 2
30 9 0 0 0 9 2 1 9 2 7 0 0 0 0 9 2 1 9 2 15 1 9 12 9 1 9 12 3 13 2
8 13 13 3 0 7 0 9 2
28 0 9 11 11 2 15 9 0 9 13 1 11 11 9 16 0 9 7 1 11 2 13 1 9 1 0 9 2
22 3 13 0 9 2 7 13 3 0 9 7 9 0 9 2 15 13 10 0 0 9 2
8 9 13 1 9 9 7 9 2
12 3 13 2 0 4 1 11 13 1 0 9 2
3 2 11 2
5 9 11 11 2 11
6 1 11 13 1 9 9
11 9 9 7 0 9 1 0 9 15 13 0
37 16 4 15 10 9 13 13 9 2 3 4 0 9 1 9 9 1 11 1 0 9 1 11 1 11 1 11 2 9 1 12 9 2 3 13 9 2
9 0 9 11 1 11 1 11 11 11
8 15 13 3 1 9 1 9 2
16 9 13 9 9 1 9 0 9 0 11 11 11 1 0 11 2
16 0 9 15 13 1 9 2 1 15 1 15 9 11 3 13 2
15 9 1 0 9 3 13 3 13 9 11 2 11 7 11 2
21 1 0 9 15 3 13 0 9 9 11 7 1 10 9 1 11 15 13 0 9 2
28 1 11 1 11 15 13 0 9 1 11 9 1 11 11 2 1 0 9 15 1 9 1 11 4 13 11 11 2
6 9 9 2 11 11 2
13 9 9 13 3 1 9 1 0 9 7 11 11 2
16 1 15 4 15 1 9 9 1 12 0 9 13 12 0 9 2
28 11 7 11 13 9 1 0 9 1 9 1 11 2 1 15 4 13 1 9 12 9 1 9 1 0 9 9 2
13 11 11 7 3 11 2 13 2 1 9 1 11 2
20 11 11 3 3 13 1 9 0 9 9 14 11 2 16 4 13 13 0 9 2
14 3 13 2 16 11 1 9 2 13 2 9 1 11 2
25 16 13 9 1 9 0 2 13 9 10 9 1 9 11 2 15 4 13 9 0 9 1 0 9 2
9 3 15 13 13 0 9 12 9 2
14 2 16 11 4 13 13 2 13 1 12 9 1 11 2
11 1 9 3 3 13 13 0 11 1 11 2
12 1 9 3 11 1 11 2 7 11 1 11 2
18 0 13 3 13 9 1 12 9 16 1 12 9 2 2 13 11 11 2
44 3 1 11 3 4 10 9 13 1 12 0 9 1 15 2 16 9 13 1 9 7 11 11 7 12 0 9 2 11 2 11 2 11 2 4 1 12 12 3 13 1 12 9 2
25 11 13 3 1 0 9 0 9 1 11 2 12 2 12 2 2 16 9 12 9 13 0 11 11 2
20 1 12 9 1 9 0 9 4 13 0 9 7 3 13 1 11 9 11 11 2
6 13 0 9 2 9 2
22 0 9 13 2 16 15 13 1 10 0 9 2 1 15 15 9 13 2 13 9 2 2
29 9 13 7 15 2 16 9 15 1 15 13 3 1 0 0 9 2 7 10 9 13 9 7 10 9 3 13 9 2
22 11 13 1 0 9 1 11 1 0 9 2 15 15 1 0 9 13 9 7 13 9 2
9 0 9 7 3 13 1 0 9 2
21 11 13 1 10 9 0 9 9 2 9 11 11 2 12 2 9 13 12 9 2 2
13 9 1 11 1 15 13 1 9 1 11 0 9 2
14 1 9 9 4 3 13 13 9 10 9 1 9 9 2
32 1 0 9 9 15 3 13 11 2 12 1 9 9 7 0 0 9 4 3 1 0 9 13 1 9 14 1 10 9 3 11 2
4 9 11 16 11
9 0 9 1 11 13 1 11 1 11
2 9 9
40 3 0 9 13 9 9 11 11 2 11 11 7 11 11 2 16 3 3 1 9 13 1 9 13 1 11 1 11 2 15 15 13 0 9 10 9 1 9 9 2
6 11 11 2 11 1 11
34 1 0 9 2 3 13 13 12 1 9 1 9 2 13 1 9 11 11 2 15 15 13 1 9 1 11 13 2 16 15 9 13 9 2
14 2 9 2 15 13 13 9 0 9 0 9 11 11 2
18 16 13 1 0 11 2 13 2 2 13 0 2 16 13 1 9 2 2
23 9 9 4 3 1 10 9 13 0 9 11 11 1 11 7 3 13 1 0 2 0 9 2
7 13 3 3 0 9 9 2
25 0 9 11 15 3 3 3 13 0 9 2 7 3 15 3 13 13 9 1 9 1 0 0 9 2
27 3 2 16 15 3 11 13 9 1 11 2 13 15 1 9 9 13 7 12 9 15 1 9 13 2 2 2
15 11 11 3 1 0 9 13 9 2 7 3 13 0 9 2
23 9 2 1 15 15 13 9 9 1 9 0 9 11 1 11 0 9 11 2 13 1 9 2
15 3 3 4 13 11 13 1 9 1 11 9 1 9 12 2
17 13 15 10 0 9 2 7 9 15 3 13 1 0 9 9 12 2
13 1 11 11 13 9 2 1 11 9 2 12 2 2
19 11 15 1 11 13 1 9 2 10 0 9 13 9 0 9 11 14 3 2
17 2 1 15 15 13 15 0 2 15 3 1 11 2 2 13 11 2
20 1 0 9 3 13 2 2 15 13 15 0 2 15 15 13 1 9 14 2 2
17 11 11 15 13 2 2 15 4 15 13 3 2 7 13 4 15 2
21 2 14 4 13 13 9 2 16 4 15 13 1 9 15 13 2 2 13 3 11 2
22 9 9 11 2 15 1 9 12 7 12 13 11 11 2 13 12 3 1 0 9 9 2
7 2 9 9 1 11 13 2
27 1 0 9 13 3 3 0 9 7 9 15 13 2 16 4 15 1 15 13 13 2 14 16 13 1 9 2
14 15 15 3 9 13 4 2 13 0 2 2 13 12 2
22 11 11 3 13 1 0 9 11 1 0 9 1 0 9 2 12 9 5 12 9 2 2
15 2 3 4 13 13 9 12 9 2 10 0 9 2 2 2
18 1 0 9 4 15 13 2 13 12 9 7 13 3 12 9 1 9 2
4 13 15 15 2
9 13 4 10 9 1 9 12 9 2
8 1 9 7 13 2 2 2 2
21 3 11 11 15 1 0 9 0 1 9 13 2 12 9 7 12 9 13 0 9 2
6 2 9 15 13 9 2
25 13 4 15 13 2 16 16 15 15 12 9 13 2 3 15 1 0 13 1 9 2 2 13 11 2
19 1 9 4 15 13 2 16 13 2 3 15 9 11 2 13 2 1 9 2
12 2 13 2 16 4 13 3 2 2 13 11 2
18 2 15 13 2 16 14 2 2 13 11 7 12 15 0 13 1 9 2
2 11 11
2 9 9
4 12 9 0 9
5 11 2 11 2 2
28 3 13 4 3 1 0 9 0 9 9 1 12 2 9 9 0 9 1 9 7 9 0 9 1 9 0 11 2
19 9 9 13 9 2 16 0 0 9 2 13 0 9 2 13 3 13 15 2
13 10 0 9 1 9 9 3 13 13 13 3 3 2
7 3 1 9 9 9 0 13
3 9 9 12
5 9 1 9 3 13
6 0 11 2 11 2 2
33 1 12 9 13 9 0 9 1 0 2 11 0 9 2 15 15 1 0 9 13 1 0 9 7 1 9 4 13 4 13 1 9 2
45 1 9 9 9 9 2 11 11 13 3 1 11 1 9 7 1 9 9 3 12 7 12 0 9 7 0 9 2 15 13 0 1 0 11 2 1 10 12 9 3 10 9 3 13 2
27 9 9 14 13 1 9 0 9 1 9 7 0 9 3 13 10 0 9 2 15 4 13 1 10 9 0 2
14 13 15 3 1 9 0 9 0 9 1 11 1 11 2
24 9 15 7 9 10 9 1 10 9 13 2 15 1 9 2 11 13 3 7 1 0 0 9 2
24 9 9 1 0 9 11 13 3 3 1 9 0 1 11 2 15 13 3 12 9 1 0 9 2
24 9 2 15 3 13 3 3 1 0 9 7 13 0 9 2 15 13 1 9 14 1 12 9 2
5 9 11 2 11 11
5 11 11 13 9 11
5 11 2 11 2 2
30 9 9 11 15 13 9 2 15 4 1 9 13 1 9 1 2 9 9 2 1 9 9 0 9 11 11 2 11 2 2
10 15 7 3 13 13 1 9 10 9 2
10 13 15 1 9 9 11 11 2 11 2
17 3 7 13 2 16 2 11 1 10 9 4 13 10 0 9 2 2
36 1 15 15 16 0 9 11 13 13 0 9 11 11 2 15 9 1 11 13 2 16 15 13 1 9 2 3 15 13 9 9 9 2 9 11 2
13 11 3 13 13 1 10 9 9 1 9 16 15 2
15 2 1 9 11 11 13 15 13 2 2 13 3 11 11 2
4 15 13 11 2
2 11 2
58 1 9 0 9 13 2 16 12 0 0 0 9 2 0 9 2 11 2 2 3 0 9 9 2 11 2 2 3 0 0 9 1 9 7 9 2 11 2 7 3 0 9 12 2 9 12 2 2 13 1 0 0 9 3 0 0 9 2
20 9 13 2 16 0 9 4 0 1 10 9 13 1 0 9 3 12 0 9 2
36 9 0 9 11 7 11 13 1 15 1 15 3 2 7 0 9 4 1 0 13 1 9 14 12 5 9 2 15 15 3 13 2 15 4 13 2
15 1 0 9 13 0 9 0 9 11 2 11 7 9 12 2
5 11 15 13 0 9
6 11 2 11 2 11 2
22 9 0 9 15 13 0 9 12 0 0 9 1 9 0 9 7 13 3 13 0 9 2
14 2 13 9 2 16 15 12 9 13 1 10 9 9 2
20 13 3 13 7 13 1 0 9 1 10 9 13 0 9 2 2 13 9 11 2
19 9 0 11 13 1 9 1 9 1 9 15 0 0 9 11 1 9 11 2
24 13 15 0 2 0 2 9 2 1 15 1 9 13 12 0 9 7 0 12 0 9 4 13 2
13 11 13 13 2 16 0 9 15 13 3 0 9 2
21 13 9 2 16 16 9 1 11 7 11 13 15 9 2 3 15 13 1 9 11 2
22 1 11 7 11 15 13 1 9 2 16 15 9 0 9 13 2 16 13 15 0 13 2
24 1 11 1 9 0 9 2 15 13 0 0 9 11 2 15 3 13 0 9 1 11 11 11 2
3 0 0 9
2 9 9
2 11 11
3 9 7 9
9 0 9 13 1 0 11 9 9 2
22 12 2 9 13 9 1 0 9 1 0 11 2 12 2 9 0 9 1 11 2 11 2
75 12 2 9 4 11 13 0 0 9 2 12 2 9 13 0 9 1 0 9 7 3 0 9 1 12 0 9 2 12 2 9 9 1 0 9 1 11 7 11 2 12 2 9 1 0 9 1 11 2 1 9 9 1 0 9 1 11 2 11 7 0 11 2 11 2 12 2 9 13 9 1 0 0 9 2
53 10 12 9 13 0 9 1 11 3 3 0 7 13 0 2 16 0 0 9 2 1 15 15 13 0 9 11 2 13 13 9 1 9 9 2 9 0 0 9 2 3 11 2 7 16 3 13 9 15 0 9 13 2
10 12 1 10 9 4 13 13 3 3 2
75 1 9 11 11 7 11 11 1 9 9 9 9 11 11 2 0 9 1 0 11 2 2 15 1 9 0 0 9 1 9 13 9 0 9 11 11 2 4 12 2 12 2 12 13 1 9 3 0 0 11 13 2 2 9 9 11 11 13 3 9 0 9 2 15 11 3 13 2 2 2 2 2 2 2 2
28 12 9 3 3 3 13 9 10 9 1 0 0 9 2 2 2 2 2 9 0 11 13 7 9 0 2 2 2
15 9 0 9 4 13 13 1 9 1 0 0 9 2 2 2
10 0 0 9 13 3 9 7 0 9 2
17 9 9 1 0 11 4 13 13 9 9 1 9 0 9 9 12 2
12 1 0 9 3 13 1 0 0 9 0 9 2
24 9 9 1 9 4 3 13 1 9 9 1 10 0 9 2 16 13 9 12 2 12 7 12 2
66 2 3 3 3 4 13 9 10 9 1 0 9 2 7 15 12 9 13 2 16 0 0 9 4 0 9 2 15 13 2 13 13 2 16 4 13 9 0 9 1 0 0 9 2 2 0 9 13 1 0 0 9 1 11 3 0 2 7 13 9 11 1 3 0 9 2
36 16 13 1 0 9 2 13 15 14 0 9 2 7 3 0 9 0 9 2 7 13 3 13 10 9 1 11 2 1 15 13 0 11 0 9 2
47 16 11 3 13 0 9 13 1 9 10 9 2 13 3 10 9 13 2 7 3 13 13 0 9 15 2 1 15 0 9 13 0 7 15 13 13 9 2 16 1 15 9 4 13 10 9 2
28 15 0 2 15 4 0 0 9 13 1 9 13 2 13 9 0 9 2 3 3 10 9 2 15 13 11 11 2
24 7 10 9 4 13 9 11 13 15 0 9 7 13 4 0 9 9 11 1 0 9 2 2 2
33 16 4 0 0 9 4 15 13 9 1 0 9 2 4 4 14 13 0 0 9 2 7 3 15 13 15 13 9 10 9 2 2 2
27 16 4 9 1 10 9 13 2 4 13 3 3 16 0 9 0 9 2 7 3 16 9 0 9 3 2 2
7 0 9 2 9 7 9 2
7 13 9 11 7 9 12 2
54 1 0 0 9 13 3 0 9 13 1 15 2 16 4 0 9 9 2 3 1 0 9 2 9 10 0 0 9 2 7 9 2 0 9 2 2 15 13 3 0 9 9 12 2 2 3 3 7 3 13 0 0 9 2
10 9 9 2 1 15 13 2 15 13 2
10 13 15 12 2 9 7 12 2 9 2
55 1 1 15 2 16 0 0 9 1 0 9 13 12 7 12 5 0 9 7 3 9 0 9 7 15 11 4 13 9 9 0 0 9 1 9 2 3 9 11 13 16 0 0 0 9 2 13 7 1 11 11 3 13 11 2
27 16 15 13 2 16 12 0 0 9 13 0 9 13 0 0 9 2 13 4 1 0 9 3 1 15 13 2
61 15 3 2 16 9 9 9 15 3 13 9 9 0 0 9 11 7 9 0 0 9 1 11 2 10 0 9 1 9 1 10 9 13 9 2 16 16 9 0 9 13 1 9 9 1 9 0 9 1 11 7 11 7 1 9 1 0 9 1 11 2
1 9
9 0 9 13 1 0 11 9 9 2
13 9 12 9 13 1 9 9 7 13 1 9 9 2
16 13 15 2 16 12 0 0 9 13 0 9 13 0 0 9 2
4 9 1 9 13
5 11 2 11 2 2
22 0 0 9 15 1 9 13 1 0 9 3 1 12 5 7 0 9 13 1 12 5 2
9 13 15 1 0 9 0 0 9 2
19 0 9 1 0 0 9 13 7 3 3 1 12 5 1 9 0 9 3 2
11 9 1 10 9 3 13 9 1 12 5 2
31 0 9 1 0 9 1 12 7 3 9 15 13 1 9 1 12 5 1 12 9 7 1 0 9 1 12 5 1 12 9 2
12 0 9 2 9 2 9 12 2 12 9 2 2
23 3 15 15 3 13 2 7 3 3 3 15 9 13 2 16 1 9 13 12 3 0 9 2
28 7 15 3 1 9 13 2 16 15 0 9 2 3 13 0 13 9 1 9 2 13 3 3 0 7 3 0 2
19 1 10 9 3 15 13 15 2 16 4 15 13 9 0 9 7 0 9 2
17 13 15 3 0 0 9 2 15 15 1 9 13 13 1 10 9 2
13 7 9 15 13 2 16 9 3 10 9 13 9 2
3 15 3 2
11 9 13 0 2 7 0 9 1 15 13 2
23 7 1 9 2 3 15 13 13 2 3 13 2 16 9 13 10 0 9 1 10 0 9 2
36 0 9 13 9 13 1 9 9 10 0 9 2 7 15 3 1 0 9 2 16 9 13 1 10 9 2 13 1 15 2 15 15 13 9 9 2
13 13 15 15 2 10 9 2 7 10 9 2 2 2
8 13 13 3 1 9 1 9 2
22 15 15 7 3 13 2 16 15 1 15 13 1 9 7 9 7 2 3 15 15 13 2
17 1 9 2 3 1 15 13 9 2 13 13 0 9 7 3 13 2
11 13 10 9 7 9 15 13 3 0 9 2
16 16 1 10 9 13 7 9 1 9 13 2 4 1 9 13 2
11 10 9 13 9 9 9 13 3 3 0 2
20 13 2 14 1 9 3 10 9 2 3 13 2 15 15 1 10 0 9 13 2
20 13 15 15 9 1 9 1 9 2 1 10 9 13 0 9 9 7 9 2 2
22 13 2 15 13 10 11 3 0 2 7 13 15 2 3 15 3 13 7 3 15 13 2
6 3 4 15 15 13 2
32 13 4 3 7 1 10 0 9 2 13 4 3 14 9 1 9 2 3 1 9 1 9 2 1 15 15 13 10 0 9 11 2
13 3 15 13 2 13 1 9 7 13 1 9 2 2
10 13 3 2 13 15 2 13 15 9 2
20 9 15 15 3 13 2 3 15 13 1 0 7 0 9 15 15 13 1 9 2
19 13 4 15 1 9 1 9 3 12 9 2 16 4 1 15 13 13 2 2
13 3 15 13 2 15 15 13 2 13 0 9 2 2
13 16 4 15 15 10 9 13 2 3 4 15 13 2
16 7 3 4 13 2 3 13 2 0 9 15 13 1 9 2 2
13 14 3 2 11 2 13 1 9 2 13 15 9 2
20 3 10 0 9 3 3 13 10 0 2 1 10 9 3 0 9 7 13 15 2
14 3 9 13 2 13 1 9 7 13 15 1 9 2 2
18 6 2 13 4 7 13 15 15 2 16 9 10 9 13 1 15 0 2
79 10 11 13 3 10 9 1 0 9 2 7 13 2 16 4 15 3 1 15 13 0 9 1 11 2 11 7 0 11 2 15 15 1 0 9 3 13 9 1 9 1 9 2 0 1 15 10 0 9 2 0 9 7 0 9 2 15 1 10 9 1 15 13 0 9 7 0 9 2 15 11 3 13 16 9 1 0 9 2
34 16 15 13 3 10 9 2 13 15 2 16 11 2 9 0 9 2 13 3 3 0 0 9 2 1 15 15 1 10 9 13 0 9 2
2 11 11
3 0 9 12
22 12 2 0 9 2 11 11 7 9 11 11 12 1 9 9 1 9 11 0 2 11 2
24 12 2 0 7 3 0 9 2 11 11 1 9 11 2 11 2 11 2 9 11 2 11 11 2
25 12 2 0 9 2 11 11 7 0 9 1 9 1 9 9 11 2 11 2 11 7 11 2 11 2
15 12 2 9 9 2 11 11 1 9 0 0 9 2 11 2
25 12 2 0 9 2 11 11 2 11 1 11 2 11 11 1 9 11 2 11 11 2 2 11 11 2
21 12 2 9 9 9 7 9 0 9 2 11 11 1 12 9 0 9 2 11 11 2
6 1 9 1 9 0 9
6 0 0 9 9 0 9
2 9 9
2 11 11
46 9 2 0 9 2 0 9 2 0 9 2 9 0 9 7 0 9 9 1 9 2 3 15 9 13 1 10 9 2 10 13 9 0 9 9 0 9 2 11 2 2 0 9 7 9 2
30 2 16 13 2 3 13 2 2 2 2 13 9 2 0 1 0 9 0 9 1 9 12 0 9 2 1 11 1 11 2
9 2 9 10 9 13 1 11 2 2
21 2 9 2 7 2 9 2 0 9 13 9 0 9 2 0 1 0 9 0 9 2
16 15 13 1 9 1 9 9 2 15 13 3 16 9 1 9 2
36 4 1 15 13 3 9 1 9 11 2 11 2 11 7 0 9 11 2 11 2 11 7 1 12 9 9 15 13 0 9 0 1 0 10 9 2
16 9 7 9 13 15 9 13 15 1 10 9 2 1 0 13 2
14 7 1 0 2 13 1 0 0 9 0 9 0 9 2
36 0 9 1 9 9 16 4 13 3 1 0 0 9 2 7 14 1 10 9 2 16 1 9 13 15 2 15 1 9 13 0 0 2 0 9 2
27 2 1 10 9 15 3 13 9 1 0 9 13 2 2 13 12 1 9 9 2 9 0 9 0 11 11 2
23 2 0 0 9 10 9 13 9 0 9 1 9 12 2 1 0 9 3 15 0 13 2 2
13 1 9 9 2 0 9 9 2 4 11 13 13 2
10 3 3 13 1 9 7 9 10 9 2
9 9 2 1 0 9 13 9 0 9
5 9 11 11 2 11
5 9 9 1 11 11
7 11 2 11 2 11 2 2
42 12 9 1 12 9 2 0 0 9 7 9 1 9 2 3 16 9 3 13 0 9 13 0 9 11 11 2 3 1 9 0 9 2 9 9 9 9 1 9 9 11 2
18 11 13 0 9 1 15 2 16 10 0 9 13 3 1 9 1 9 2
26 0 9 2 11 2 3 13 0 9 1 11 2 10 9 13 11 2 7 11 13 1 2 0 9 2 2
11 2 13 3 11 13 2 2 13 3 11 2
2 9 9
3 9 1 9
14 11 11 2 9 9 11 2 2 1 11 13 9 13 2
11 10 0 9 15 1 9 1 11 13 9 2
34 2 11 11 2 9 11 2 2 9 9 15 13 1 9 2 16 15 9 13 1 9 1 9 11 11 2 15 13 9 1 9 1 11 2
9 11 13 3 0 9 1 9 2 2
7 9 1 0 9 9 11 13
5 11 2 11 2 2
18 11 13 1 9 1 11 2 12 2 12 2 1 0 9 7 13 9 2
6 2 9 0 15 13 2
14 0 9 13 13 3 2 2 13 1 9 9 9 11 2
15 2 13 4 3 16 1 0 9 2 2 13 0 9 11 2
9 9 10 9 13 0 9 9 9 2
22 2 16 15 1 10 0 9 11 2 11 2 11 2 11 15 3 13 2 13 3 3 2
7 3 13 1 15 7 9 2
19 1 0 9 9 3 13 9 2 2 13 11 2 15 12 1 0 9 13 2
16 2 11 4 13 3 3 3 2 7 11 9 3 3 13 2 2
29 0 9 11 2 1 15 2 3 16 1 0 11 7 11 2 13 9 9 1 0 9 11 1 11 2 3 9 13 2
14 0 13 3 12 7 0 9 13 1 0 3 1 9 2
6 0 9 13 1 0 9
5 11 2 11 2 2
28 9 1 9 9 7 0 0 0 9 2 11 2 1 9 0 9 4 1 0 9 3 13 2 12 2 9 2 2
26 9 11 11 11 4 3 1 10 9 1 9 11 1 11 13 1 9 2 2 3 1 0 9 15 13 2
29 13 7 0 13 2 16 9 3 11 2 9 0 9 2 13 3 9 1 9 2 3 11 2 13 3 1 9 12 2
7 0 9 15 10 9 13 2
28 1 9 0 9 4 13 13 2 16 9 1 9 13 1 9 9 12 16 9 0 9 1 11 2 9 7 11 2
28 9 1 9 13 13 1 0 7 3 2 16 10 0 9 3 13 3 0 9 2 3 9 9 3 1 9 9 2
37 9 11 1 0 9 4 0 9 2 7 3 7 9 9 13 7 13 4 15 9 1 9 0 9 0 2 1 15 0 9 9 3 10 9 13 2 2
9 9 9 15 14 1 9 13 3 3
5 11 2 11 2 2
25 1 9 2 16 4 0 9 9 13 0 9 7 9 13 3 9 11 1 9 11 11 2 12 2 2
22 9 11 13 1 9 0 9 16 0 1 9 12 2 0 1 9 7 0 1 9 12 2
23 1 0 7 0 0 9 15 1 0 9 13 12 9 7 0 9 1 9 13 3 12 9 2
23 0 9 13 0 9 11 11 2 15 4 13 12 2 9 12 7 13 12 2 9 10 9 2
11 3 0 13 11 11 2 12 2 12 2 2
24 1 9 2 15 13 9 9 11 2 11 13 0 9 2 7 15 11 11 2 12 2 12 2 2
24 1 9 2 0 9 2 13 11 2 12 9 9 13 7 9 2 12 0 9 7 12 0 9 2
26 11 15 3 3 13 2 15 4 13 0 9 0 9 2 1 0 9 4 7 13 13 1 9 1 11 2
14 1 9 13 9 9 0 9 2 15 13 0 9 9 2
33 1 9 2 1 3 13 1 9 9 1 0 9 2 13 2 16 9 0 1 9 3 0 4 13 4 13 1 0 9 12 2 12 2
2 11 11
25 1 9 9 13 3 3 12 7 9 9 7 11 15 3 13 13 0 0 9 2 15 4 15 13 2
3 3 3 2
30 9 0 7 0 2 1 0 9 15 3 13 15 7 15 2 13 7 1 0 9 2 16 15 7 9 13 0 15 9 2
7 7 16 13 3 0 9 2
40 1 9 0 9 15 3 9 13 13 2 3 1 9 9 11 11 2 16 0 9 13 3 0 9 2 0 9 2 15 4 13 9 7 3 13 9 7 0 9 2
23 13 7 9 0 2 0 9 1 9 9 13 3 13 7 0 9 15 7 3 13 1 9 2
17 9 9 9 2 3 0 9 9 2 13 3 12 1 9 10 9 2
17 3 13 2 0 9 1 0 9 3 13 1 11 13 1 15 0 2
32 0 9 13 7 9 9 9 1 9 2 11 2 11 2 2 7 7 9 9 2 11 2 11 2 7 9 2 11 2 11 2 2
17 0 11 2 9 2 1 10 9 13 16 13 9 1 9 0 9 2
32 14 3 13 9 0 0 9 3 0 2 0 13 15 2 1 11 3 13 2 13 2 9 2 10 0 9 13 1 0 9 9 2
16 0 9 13 1 10 9 0 3 2 16 15 15 13 7 3 2
34 1 9 3 4 13 9 2 7 9 2 4 13 12 9 1 0 2 3 3 2 16 15 15 0 9 1 10 9 13 2 7 3 13 2
16 13 7 9 10 9 2 3 9 9 7 9 9 2 11 0 2
16 9 10 9 13 3 2 13 3 0 9 2 7 7 15 13 2
7 7 16 14 2 3 3 2
30 9 9 13 1 9 2 7 11 1 15 13 2 16 1 9 0 0 9 3 13 3 2 16 3 3 2 16 0 11 2
9 0 9 13 2 3 2 13 9 2
20 15 1 15 7 0 0 9 2 15 1 0 9 13 2 16 0 9 13 0 2
8 9 3 13 2 13 15 15 2
1 12
9 1 11 15 13 9 1 0 9 11
5 11 2 11 2 2
19 1 11 7 11 2 11 15 3 13 0 9 0 9 1 9 0 0 9 2
11 9 9 11 13 3 0 9 0 9 11 2
15 1 0 9 15 3 13 14 12 9 9 1 11 7 11 2
11 13 1 9 2 14 3 15 13 0 9 2
8 0 9 13 3 3 1 9 2
32 1 12 9 9 1 0 9 9 3 13 12 7 12 9 9 7 16 13 9 0 9 1 11 11 11 2 9 15 3 3 13 2
22 9 0 9 11 11 15 1 9 1 0 0 9 13 2 1 10 9 9 1 11 13 2
30 3 15 9 1 11 13 3 2 1 9 7 9 1 9 11 7 11 2 15 13 3 1 9 0 9 12 9 1 11 2
20 16 13 1 0 9 2 9 15 7 1 12 9 13 7 13 3 9 7 9 2
16 16 13 9 2 1 9 12 1 0 9 3 13 9 0 9 2
29 11 11 1 11 11 13 2 16 12 9 9 2 15 13 1 0 9 1 11 2 13 0 0 9 7 0 13 9 2
25 1 3 0 9 2 3 3 13 3 12 9 9 2 13 9 9 1 9 7 9 9 1 0 9 2
13 9 13 2 16 7 0 9 13 1 9 0 9 2
11 9 2 1 11 13 9 11 3 0 9 2
12 3 4 13 1 11 13 7 9 1 0 9 2
5 9 11 11 2 11
2 11 13
2 11 2
10 1 0 9 13 1 0 9 9 9 2
18 1 12 0 9 4 13 12 9 2 1 12 3 16 1 12 9 2 2
24 1 0 3 2 0 0 9 1 9 7 9 2 12 2 7 9 0 9 9 12 2 12 2 2
4 13 15 0 9
8 11 13 9 9 11 1 3 0
5 11 2 11 2 2
15 13 1 9 0 9 13 9 2 3 3 0 7 0 2 2
33 13 15 3 9 11 11 11 1 9 11 2 3 10 9 1 0 9 1 0 9 13 11 2 11 2 11 7 11 3 1 10 9 2
31 2 13 3 13 2 16 13 1 0 9 9 2 16 15 9 1 10 9 13 2 13 15 15 2 13 7 3 15 13 2 2
23 3 4 13 1 15 13 0 9 0 9 11 2 2 13 15 9 7 9 2 13 15 2 2
26 0 9 13 1 11 3 0 9 2 16 1 10 9 13 13 1 0 9 1 0 9 1 9 0 9 2
58 1 9 1 0 9 9 11 11 11 11 2 16 9 9 1 0 9 13 0 9 9 1 10 9 2 9 11 13 2 16 2 16 15 0 0 9 13 13 2 16 4 3 4 0 9 13 2 13 0 2 16 1 15 13 10 9 2 2
22 0 0 9 9 7 9 13 13 1 11 0 9 9 2 7 2 9 2 9 7 9 2
20 2 9 13 0 9 2 13 15 15 7 3 3 13 1 9 2 2 13 9 2
21 11 1 15 13 2 16 9 3 1 10 9 2 13 13 13 0 9 0 9 2 2
20 9 7 13 1 0 9 0 2 0 9 2 15 13 13 0 2 0 7 0 2
14 0 9 1 0 9 9 11 11 4 13 3 9 13 9
2 9 9
2 11 9
57 3 16 0 0 9 3 3 13 0 9 7 16 0 9 1 9 1 9 13 9 0 9 2 13 0 12 0 9 2 1 0 2 16 15 1 0 0 9 13 10 9 9 2 16 4 13 12 0 9 7 15 7 9 13 13 9 2
23 3 1 9 15 13 1 0 2 16 0 9 13 2 16 3 13 1 11 9 2 9 0 2
14 1 0 2 0 9 9 13 10 0 9 1 0 9 2
26 1 0 9 0 9 13 7 0 2 16 1 9 10 7 15 9 3 13 9 3 10 2 0 2 9 2
34 1 0 2 16 9 0 0 9 7 0 0 9 15 9 11 11 2 1 9 9 0 12 9 2 15 1 0 9 1 0 9 4 13 2
10 1 0 2 3 1 11 13 0 9 2
27 16 10 9 13 3 3 2 1 11 2 0 1 13 9 3 3 16 1 9 0 9 2 13 15 9 0 2
10 0 9 1 9 13 7 15 1 9 2
15 1 9 11 13 1 9 9 1 0 0 9 3 0 9 2
43 16 9 9 7 0 9 13 10 9 0 0 0 9 2 11 2 13 1 0 9 3 7 1 0 0 9 1 9 7 9 2 11 2 2 7 1 0 9 9 2 11 2 2
20 0 9 0 9 11 13 9 0 9 3 1 9 2 3 0 9 13 0 9 2
45 16 9 0 9 13 13 1 11 9 2 13 3 1 9 0 9 2 16 10 0 9 13 13 2 13 15 13 1 9 1 13 9 2 1 9 1 15 2 16 13 0 7 0 9 2
10 9 1 0 9 3 3 11 4 13 2
8 10 9 15 1 15 7 13 2
10 9 1 9 13 3 1 0 0 9 2
15 1 12 9 11 15 3 9 13 9 1 9 7 0 9 2
24 0 9 4 13 9 13 0 2 7 0 9 2 9 1 0 9 7 9 1 9 15 13 13 2
9 14 3 13 13 0 9 0 9 2
13 3 0 11 4 9 10 9 3 13 7 13 15 2
20 16 15 13 13 9 9 0 9 1 11 11 2 16 13 13 2 13 3 0 2
43 0 7 13 15 2 15 3 13 15 9 0 9 2 9 2 15 13 13 1 0 0 9 2 13 0 16 10 2 15 13 1 9 9 1 9 12 2 3 11 13 1 9 2
6 1 9 9 1 0 9
30 1 11 4 3 13 4 13 0 9 1 11 7 9 1 9 11 2 11 2 1 0 0 9 1 9 11 7 1 11 2
4 15 9 13 2
21 12 2 12 2 12 2 0 9 1 11 7 11 1 0 0 9 7 1 0 9 2
18 12 2 12 2 12 2 1 11 7 1 0 9 11 13 9 0 9 2
30 10 9 15 13 3 9 0 9 2 9 0 9 0 1 11 2 9 0 9 1 0 9 1 0 2 9 0 9 3 2
7 9 3 13 9 1 11 2
29 12 2 2 12 2 12 2 12 2 11 11 7 11 11 1 9 1 11 13 0 0 9 1 0 9 0 0 9 2
21 12 2 12 2 12 2 0 9 2 0 9 11 11 13 1 9 12 9 9 2 2
18 12 2 12 2 12 2 11 7 11 13 1 11 9 1 0 0 9 2
8 13 9 1 0 9 1 11 2
10 11 13 9 0 0 9 1 0 9 2
27 12 2 12 2 12 2 11 7 11 15 13 2 16 12 2 9 13 1 11 0 9 1 9 0 0 9 2
17 12 2 12 2 12 2 0 9 13 9 11 0 1 9 0 9 2
9 9 1 9 13 7 0 9 11 2
20 12 2 12 2 12 2 11 2 11 7 11 2 11 13 1 11 1 0 0 9
3 2 11 2
6 1 15 13 1 0 9
10 0 0 9 2 1 10 9 15 9 13
2 9 9
18 9 2 0 0 9 2 11 2 13 9 0 9 1 0 9 0 9 2
9 13 0 9 1 9 1 0 9 2
9 9 3 13 1 3 0 9 9 2
15 10 10 9 7 1 15 3 3 13 16 1 12 1 9 2
18 0 9 9 11 7 3 0 0 9 2 11 2 15 13 1 0 9 2
21 3 0 0 9 11 15 13 1 9 9 1 9 1 9 2 9 2 9 7 9 2
18 11 13 2 0 2 0 9 2 15 4 13 9 2 9 7 0 9 2
30 0 9 2 3 3 13 12 0 0 9 9 13 0 9 7 13 9 0 9 2 15 3 13 3 0 9 1 0 9 2
9 0 2 0 2 9 13 7 11 2
21 11 13 0 9 9 0 9 2 15 4 0 9 13 1 9 2 9 7 0 9 2
16 13 9 2 15 4 1 0 9 13 9 7 9 12 9 9 2
17 9 9 2 9 9 9 7 0 9 13 1 0 0 9 0 9 2
32 11 13 7 1 10 9 0 9 1 2 0 0 9 2 7 0 7 0 9 2 15 4 13 9 7 13 9 0 9 1 15 2
22 9 2 15 9 13 13 1 3 0 9 2 15 13 1 12 9 9 9 12 0 9 2
17 11 13 10 9 0 0 9 2 15 4 15 13 0 1 0 9 2
14 3 4 10 9 13 13 0 0 9 2 1 15 13 2
19 13 3 0 9 1 9 0 9 2 16 4 15 13 13 9 9 1 9 2
15 11 13 9 0 9 7 9 7 9 9 1 0 0 9 2
28 0 9 11 13 2 9 0 0 9 2 1 15 13 15 13 1 0 9 7 13 10 9 1 9 7 9 2 2
17 0 0 9 13 1 9 1 10 9 1 0 9 9 9 9 9 2
8 9 2 11 13 0 0 9 2
21 11 2 0 9 7 0 9 15 13 1 0 9 1 0 9 0 7 0 0 9 2
11 0 9 13 0 0 9 2 2 9 2 2
23 11 3 0 7 3 0 9 0 9 2 1 15 4 13 3 9 9 7 9 0 0 9 2
14 0 9 7 10 0 9 2 11 12 2 12 2 12 2
16 0 0 9 1 11 4 1 9 9 11 13 3 1 9 9 2
13 11 15 3 3 13 7 14 1 12 9 3 13 2
19 13 9 1 9 2 12 7 1 0 9 11 3 1 9 2 12 1 12 2
21 9 2 1 9 9 9 2 1 9 1 9 9 2 16 13 11 2 13 0 9 2
24 1 10 9 4 1 9 12 9 1 9 7 12 9 1 9 13 0 3 13 9 1 12 9 2
28 0 9 13 9 0 9 2 3 1 9 13 1 9 2 7 1 9 9 1 9 2 10 9 7 9 0 9 2
6 13 1 15 10 9 2
10 1 0 9 4 13 9 1 9 9 2
17 16 4 13 13 9 1 12 9 7 13 1 12 13 13 9 13 2
8 0 13 9 13 9 1 9 2
19 13 9 0 9 7 9 3 13 1 9 1 0 11 1 9 1 0 9 2
25 1 3 0 9 0 9 1 9 4 15 13 9 13 3 2 3 16 15 13 3 2 1 0 11 2
14 1 0 9 9 7 9 13 7 9 9 7 10 9 2
20 15 13 12 9 1 9 1 0 7 0 9 2 16 13 1 9 9 1 9 2
11 14 13 2 16 15 1 15 4 15 13 2
42 10 9 1 9 1 9 2 12 2 3 15 9 7 10 9 13 9 7 9 9 1 11 7 1 11 2 7 1 9 2 12 2 3 3 13 1 10 9 7 9 9 2
6 1 9 11 11 2 11
3 0 9 9
6 9 11 13 1 0 9
3 0 11 2
13 0 9 13 1 0 9 9 0 9 9 0 11 2
32 9 13 1 9 11 13 7 1 0 9 1 11 2 3 13 12 2 12 2 16 0 9 13 12 2 12 1 9 9 11 11 2
23 15 13 3 1 11 11 7 0 9 11 2 15 13 12 9 0 9 2 0 9 0 9 2
22 11 3 13 9 1 12 2 9 1 11 11 7 1 0 9 13 7 1 9 1 11 2
18 0 9 15 13 13 1 10 9 7 1 9 9 3 13 12 2 12 2
41 1 0 9 15 15 13 3 13 1 12 2 12 2 7 9 11 1 11 12 2 12 1 9 3 13 9 1 9 7 15 13 1 0 9 12 9 1 0 9 11 2
2 0 9
2 11 2
26 0 0 9 9 0 9 1 9 0 9 0 0 11 11 12 13 10 9 0 9 1 0 9 1 11 2
18 0 9 13 0 7 0 9 7 1 0 9 15 13 9 1 12 9 2
21 12 9 9 15 13 1 0 9 2 0 9 1 9 1 11 7 12 1 0 11 2
16 13 15 1 9 1 12 9 2 12 9 2 9 12 7 9 2
38 9 4 13 13 9 0 9 9 1 9 1 12 9 11 11 2 15 15 3 13 1 0 0 9 1 11 7 1 0 9 13 13 7 1 0 0 9 2
5 9 2 11 0 9
2 11 2
5 11 15 13 13 11
9 9 1 11 13 1 11 9 0 9
2 9 9
7 11 2 11 2 11 2 2
25 1 9 1 11 3 1 0 9 3 13 9 11 7 0 11 2 16 4 15 13 1 9 9 9 2
22 3 1 9 1 0 0 9 1 9 12 15 3 1 9 0 9 13 0 7 0 9 2
15 9 13 9 11 11 2 15 9 13 1 9 9 1 9 2
11 16 3 11 13 2 13 16 0 9 11 2
36 9 11 11 13 1 15 1 9 15 9 2 1 0 9 1 11 11 13 13 7 1 9 11 7 0 9 11 2 1 9 15 3 13 11 11 2
23 0 9 11 11 15 3 13 1 0 9 2 13 13 11 2 11 11 2 11 7 9 11 2
24 3 11 13 2 2 15 13 13 2 16 11 13 3 0 3 2 16 15 15 1 15 13 2 2
29 1 9 1 9 9 13 3 9 1 11 0 9 13 1 0 9 3 0 9 7 1 9 15 4 13 12 12 9 2
27 11 2 10 9 13 1 0 9 1 12 9 9 2 13 3 1 12 2 9 1 9 0 9 1 9 11 2
27 9 1 0 0 9 11 13 1 12 9 2 13 11 12 2 7 13 15 9 0 9 11 2 11 2 11 2
12 9 13 9 11 2 11 1 9 7 11 2 11
5 11 2 11 2 2
33 0 9 1 11 3 13 9 1 9 9 0 9 0 0 9 11 11 1 0 0 9 2 9 2 7 1 0 9 0 9 11 11 2
19 11 13 9 9 11 0 7 0 0 9 9 9 11 2 11 1 0 9 2
35 0 15 13 13 1 15 2 16 13 9 1 9 9 11 2 11 2 15 3 2 1 11 2 13 9 11 9 11 2 16 9 13 3 0 2
15 11 4 13 1 0 9 9 1 0 0 9 1 9 12 2
42 11 13 1 9 2 16 4 15 0 9 2 13 2 13 1 15 2 16 13 9 9 7 13 10 9 2 7 15 15 2 16 13 1 9 2 16 9 0 9 13 0 2
23 11 15 13 13 1 10 9 2 0 9 11 11 2 2 11 2 12 2 12 2 12 2 2
29 1 9 13 10 9 7 0 9 9 7 13 9 9 2 2 16 9 13 2 16 0 9 0 9 9 13 13 2 2
27 9 13 9 1 9 7 2 16 15 1 9 13 9 9 9 1 9 9 7 9 1 9 9 1 0 9 2
16 9 1 11 13 7 2 16 1 9 9 13 9 2 7 9 2
25 11 7 0 9 9 15 2 1 0 9 2 3 13 15 2 16 9 13 9 1 9 1 9 9 2
15 11 2 11 1 9 9 9 13 9 0 0 9 1 11 2
5 9 1 11 1 9
5 11 2 11 2 2
21 10 9 4 13 9 9 11 2 11 2 13 1 0 0 9 2 11 2 1 9 2
9 13 1 15 9 9 11 11 11 2
24 9 11 15 13 9 0 9 2 0 9 2 0 9 15 12 9 7 9 0 1 9 9 11 2
18 9 1 9 13 9 11 13 3 1 9 11 3 1 12 2 9 12 2
5 9 9 1 9 12
2 0 11
5 11 2 11 2 2
13 0 9 11 1 9 0 9 13 3 3 3 13 2
14 13 15 9 0 7 0 9 9 11 11 2 11 2 2
8 11 1 9 9 9 9 9 13
2 11 2
24 0 9 9 13 1 9 9 1 9 0 0 9 7 1 2 9 1 9 2 1 10 0 9 2
16 9 9 13 10 9 2 16 4 1 0 9 13 9 9 9 2
20 0 9 9 11 11 13 0 9 1 9 1 9 0 9 7 0 9 1 9 2
16 13 15 1 9 1 2 9 2 2 15 13 9 1 0 9 2
5 11 2 11 2 2
33 9 11 1 11 1 0 7 0 9 7 1 0 9 1 0 9 0 1 9 11 13 3 11 11 9 0 9 0 1 11 11 11 2
23 11 11 13 1 0 9 7 0 9 9 9 0 9 7 9 11 1 9 0 7 0 11 2
21 12 9 13 9 9 0 9 1 11 2 3 13 16 0 9 1 0 9 1 11 2
16 9 11 1 11 1 0 9 13 9 10 9 10 9 0 9 2
16 9 2 9 0 11 11 11 2 9 11 11 7 9 11 11 11
5 9 11 11 2 11
4 11 15 13 11
15 9 11 13 13 9 7 13 1 9 1 0 9 7 16 0
2 9 9
28 0 0 9 13 1 12 2 9 9 1 11 9 2 15 13 1 0 9 1 0 9 2 7 3 15 13 9 2
32 3 1 12 9 13 1 11 1 15 2 16 10 9 0 9 1 15 13 0 9 9 7 13 1 9 1 9 3 0 0 9 2
24 3 0 9 13 9 11 11 2 2 15 13 1 12 9 7 3 13 1 15 13 15 0 2 2
7 0 9 11 1 11 11 11
30 11 1 9 13 9 7 1 11 2 7 1 9 0 0 9 13 0 2 16 11 15 1 0 9 13 9 12 2 12 2
18 9 11 3 1 9 13 2 16 13 1 10 9 0 11 2 7 11 2
19 9 11 2 11 7 0 9 2 11 15 13 3 2 15 11 3 13 9 2
31 10 9 7 3 1 0 12 13 12 2 12 7 15 13 2 16 4 0 9 13 1 9 1 0 12 9 11 1 9 11 2
11 11 13 12 12 2 12 7 13 15 3 2
18 2 3 4 1 15 13 13 2 2 13 3 9 0 11 11 11 11 2
18 7 7 11 13 3 13 1 15 2 16 15 0 9 13 1 10 9 2
32 12 1 9 9 11 11 11 11 13 1 11 1 11 1 11 13 0 9 7 13 15 13 2 2 9 9 13 3 0 16 7 2
52 1 10 9 13 15 12 2 1 15 4 13 2 7 9 13 3 1 15 2 16 16 11 13 1 9 2 13 3 0 2 2 13 0 0 9 9 1 0 9 2 1 15 15 10 10 9 1 11 1 11 13 2
18 0 9 13 1 9 9 2 10 9 1 9 1 11 13 3 12 9 2
29 13 1 15 10 0 9 2 16 9 11 7 9 11 2 12 11 2 2 11 2 0 11 2 2 11 2 11 2 2
16 3 7 13 11 11 2 2 11 13 9 3 3 16 9 2 2
29 2 3 13 1 9 2 2 13 9 0 9 11 11 1 0 9 10 9 2 3 15 13 3 9 7 9 1 9 2
12 2 3 15 13 2 2 13 15 9 11 11 2
16 2 9 13 0 2 16 9 1 9 13 0 9 1 9 2 2
19 3 15 7 13 2 16 4 9 13 12 9 1 0 9 10 9 11 11 2
24 11 11 3 13 2 1 15 13 0 9 10 9 2 2 11 4 13 3 0 9 16 3 11 2
9 13 4 15 3 13 3 0 9 2
12 13 15 7 0 9 1 0 9 7 1 9 2
18 9 4 13 13 9 0 9 9 7 3 3 15 9 13 3 13 2 2
25 1 9 10 9 13 11 2 1 11 11 2 15 1 0 9 0 9 13 13 2 4 13 13 11 2
19 1 9 15 4 13 12 9 1 15 2 16 16 0 0 9 13 13 11 2
15 2 1 0 12 15 13 2 15 3 2 2 13 11 11 2
22 9 11 11 2 2 13 13 10 9 2 15 13 0 2 15 4 16 9 1 9 13 2
12 15 3 13 1 9 13 1 9 1 0 9 2
3 0 9 9
3 0 11 2
18 9 0 11 13 7 3 1 0 9 1 12 2 9 9 14 1 11 2
8 9 13 13 9 1 9 9 2
16 0 11 13 3 3 3 11 11 2 7 16 3 14 1 9 2
23 0 3 13 12 2 12 2 16 1 12 1 9 13 11 2 7 9 13 1 12 2 12 2
21 9 15 3 13 12 9 1 9 11 2 7 1 10 0 9 13 1 9 9 11 2
21 4 13 0 7 0 2 1 11 7 1 11 3 0 9 12 7 12 9 5 9 2
2 0 9
2 11 11
12 1 12 0 9 13 0 9 1 9 0 9 2
14 13 15 1 11 12 2 9 12 2 0 9 0 9 2
13 9 13 0 0 9 7 13 15 15 9 7 9 2
22 15 15 13 2 15 1 15 13 2 4 13 10 9 3 1 0 0 9 1 9 11 2
15 13 15 3 9 0 2 13 0 9 9 9 1 9 0 2
15 0 9 0 9 13 1 11 3 14 9 0 9 0 9 2
19 1 0 9 15 13 9 3 9 9 2 1 12 9 9 15 3 13 3 2
42 3 13 2 16 11 13 13 2 7 9 9 2 3 13 2 16 0 9 13 13 2 1 9 13 10 9 7 1 15 11 3 13 10 9 2 15 13 2 1 9 2 2
20 3 15 7 3 13 1 15 2 16 9 2 1 15 15 9 13 2 0 13 2
8 10 9 15 13 0 0 9 2
7 11 15 1 11 13 13 2
7 9 7 13 10 0 9 2
21 15 9 1 9 1 11 13 13 7 13 7 15 1 9 4 15 1 15 13 13 2
7 9 11 7 10 9 13 2
9 13 15 13 9 2 15 13 9 2
4 13 14 9 2
7 0 9 1 0 9 13 2
16 0 11 13 1 9 0 0 9 2 15 13 1 9 0 9 2
15 16 0 9 13 2 1 11 3 9 13 1 9 0 9 2
9 0 9 1 11 3 13 10 9 2
10 1 12 9 9 13 1 12 9 9 2
9 12 9 0 0 9 13 12 9 2
11 15 13 1 9 7 9 9 1 0 9 2
10 9 9 7 3 9 1 11 13 13 2
32 4 1 15 13 3 7 3 2 1 9 12 1 9 9 1 0 9 7 1 9 9 12 1 9 0 7 0 9 3 1 11 2
19 2 13 15 13 2 2 13 9 9 0 9 2 16 13 3 13 9 9 2
10 13 4 3 3 3 7 3 1 11 2
11 12 2 9 15 1 0 9 13 0 9 2
11 0 9 13 0 2 9 0 9 15 13 2
46 16 1 9 0 9 11 11 2 1 12 9 3 13 1 11 13 1 9 2 13 10 9 9 11 2 2 3 10 9 13 1 11 1 9 0 9 3 7 1 0 9 9 0 9 2 2
26 13 15 1 9 13 2 3 7 16 3 4 0 0 9 2 0 9 11 1 9 11 2 13 10 9 2
10 13 7 9 2 15 15 13 2 13 2
15 1 11 15 12 2 9 12 13 14 9 7 0 0 9 2
10 3 13 2 16 14 1 12 0 9 2
11 0 9 13 3 0 9 14 1 9 0 9
15 1 12 2 9 13 1 0 9 12 0 7 12 0 9 2
30 1 0 9 13 0 0 9 2 12 2 7 0 0 9 2 12 2 2 16 9 13 14 12 7 9 0 3 14 12 2
36 9 7 13 1 9 0 9 2 9 2 16 4 0 9 13 0 9 9 2 15 1 9 13 1 15 1 9 2 2 4 15 13 3 12 9 2
8 15 15 13 0 9 0 9 2
24 13 4 15 9 0 0 9 2 9 2 11 11 2 9 0 0 0 9 1 11 12 2 11 2
12 2 9 13 3 0 2 0 9 15 15 13 2
21 3 3 9 9 13 1 10 9 9 1 9 9 0 9 2 16 0 9 3 13 2
14 15 13 7 1 9 1 9 2 15 9 3 13 2 2
12 16 9 9 9 7 9 0 9 1 9 13 2
32 2 9 13 2 16 10 9 3 13 7 13 2 7 13 2 16 13 15 2 15 13 1 0 2 13 1 0 9 9 7 9 2
27 1 9 0 7 0 9 15 13 13 3 16 13 9 1 0 9 7 0 9 1 9 2 15 13 3 0 2
13 13 13 1 0 9 0 9 2 16 13 9 0 2
8 9 13 9 9 1 9 2 2
11 15 3 3 13 0 9 0 9 2 2 2
7 2 13 7 0 0 9 2
29 1 0 9 4 13 4 13 9 9 2 3 4 4 13 9 1 0 9 2 13 9 2 13 9 7 0 9 3 2
32 9 7 13 1 10 9 13 2 13 13 9 9 2 7 3 15 13 13 2 16 13 15 15 2 15 13 1 9 7 9 9 2
13 1 9 13 9 9 1 15 9 0 7 0 2 2
7 13 2 16 15 4 13 2
26 2 3 1 11 15 1 12 0 9 1 0 9 13 9 9 2 16 0 9 1 0 9 15 7 13 2
12 9 13 1 15 2 16 4 15 13 9 2 2
7 9 1 0 9 3 13 2
27 1 9 9 2 11 15 3 13 0 9 9 16 3 2 12 2 2 16 3 1 11 13 0 12 0 9 2
29 0 9 3 13 0 0 9 2 15 3 13 0 9 7 9 2 16 13 13 1 0 9 1 9 9 1 0 9 2
11 13 7 13 9 0 0 9 7 0 9 2
22 9 15 3 13 2 7 16 15 13 13 9 1 0 9 2 13 9 7 9 3 3 2
11 1 10 9 3 0 0 9 13 1 9 2
30 1 3 0 9 9 0 9 1 9 7 9 9 9 0 0 7 0 9 2 15 13 1 9 9 9 2 3 3 13 2
2 11 11
4 9 2 11 11
6 15 3 3 13 9 9
19 9 7 9 13 1 0 9 0 0 9 2 12 7 12 9 1 9 0 2
26 1 9 3 13 0 9 9 1 9 1 9 2 9 7 9 2 1 15 3 4 13 0 7 0 9 2
22 3 1 9 13 1 9 1 0 9 9 1 10 9 2 3 1 9 9 13 0 9 2
14 1 0 9 13 13 1 0 9 1 0 0 0 9 2
3 0 9 2
26 1 9 1 0 9 13 9 9 7 0 9 3 0 0 9 2 10 0 9 13 9 0 9 11 9 2
34 1 0 9 1 0 9 15 13 3 3 12 9 9 2 16 4 13 13 1 12 9 9 0 9 2 3 13 0 9 9 7 0 9 2
23 9 0 0 9 2 15 13 1 9 0 9 13 0 9 2 13 1 9 1 9 11 11 2
32 13 7 9 2 15 2 13 9 9 0 9 2 13 3 3 13 9 1 9 7 9 1 9 3 3 0 2 14 3 1 9 2
56 16 9 1 9 11 7 11 1 0 9 13 9 9 1 10 0 9 2 13 15 3 9 0 9 2 15 10 0 2 0 9 0 9 13 13 9 0 0 9 3 2 16 4 15 10 9 3 13 2 7 12 9 10 9 13 2
23 1 9 0 9 13 7 1 10 9 9 0 9 0 9 2 15 3 13 9 9 11 9 2
20 7 15 15 3 13 1 9 12 9 2 10 9 4 9 2 9 13 2 13 2
40 1 0 0 9 2 3 4 3 9 1 0 9 13 0 9 9 7 9 0 9 0 9 9 2 13 9 3 1 0 9 2 1 9 2 3 3 0 9 13 2
30 13 4 0 15 13 2 16 1 9 1 0 0 9 13 3 0 9 1 0 9 9 0 9 13 1 0 9 12 9 2
14 9 1 11 7 11 3 13 0 9 0 9 1 9 2
30 1 9 7 13 13 11 9 1 9 2 9 15 4 3 13 2 16 3 1 0 9 1 9 9 13 9 1 15 0 2
24 7 16 4 7 9 13 0 2 1 0 9 13 0 0 9 2 13 9 0 9 9 3 13 2
16 9 0 0 9 4 3 9 13 1 0 9 3 0 0 9 2
3 3 13 2
25 9 2 3 13 1 11 3 7 3 2 3 9 2 1 9 3 7 3 3 3 0 9 1 9 2
23 0 9 1 11 12 7 12 9 2 9 2 1 11 7 1 11 12 7 12 9 2 9 2
16 0 12 7 12 9 2 9 2 1 12 9 12 9 2 9 2
23 0 9 12 7 12 9 2 9 2 1 9 1 9 9 3 1 9 1 12 9 2 9 2
20 2 1 11 3 3 0 9 2 1 9 9 9 7 9 2 3 1 9 2 2
17 9 13 1 9 1 12 2 12 9 7 13 1 12 2 12 9 2
17 9 13 1 9 1 12 2 12 9 7 13 1 12 2 12 9 2
23 9 9 2 0 12 9 2 9 1 9 2 12 2 0 12 9 2 9 1 9 2 12 2
11 0 9 2 0 9 0 2 0 9 0 2
5 0 9 2 11 2
4 12 9 1 11
5 11 2 11 2 2
20 1 9 1 9 0 9 0 0 9 1 0 9 11 11 4 13 0 9 9 2
27 1 0 9 9 1 9 2 9 7 9 0 9 4 3 1 0 9 13 12 9 2 3 9 11 11 9 2
18 12 9 0 9 4 13 1 9 2 11 9 3 1 0 0 1 9 2
10 1 9 1 15 4 13 9 1 9 2
4 0 9 9 13
8 1 11 13 9 9 11 2 11
34 0 0 0 9 0 11 2 0 1 9 9 0 11 2 15 3 14 13 13 9 0 2 9 9 2 1 11 11 11 7 9 11 11 2
31 7 9 9 1 9 7 9 9 0 9 1 11 7 0 9 13 9 9 1 9 9 9 12 2 15 3 1 11 13 11 2
9 7 1 9 13 9 12 9 9 2
12 3 4 9 3 13 2 3 15 13 1 9 2
25 10 9 13 2 16 15 4 13 1 9 1 0 9 2 7 1 9 11 15 3 13 13 1 9 2
12 1 12 9 13 11 2 12 2 10 0 9 2
8 1 9 9 13 11 0 9 2
19 3 15 13 10 0 9 2 7 0 9 2 0 9 1 0 9 7 0 2
12 13 1 9 2 3 10 9 13 9 0 9 2
30 1 9 9 11 11 13 11 2 3 0 9 2 7 14 13 0 9 1 15 2 16 4 9 13 13 0 0 9 9 2
17 0 9 7 3 13 0 9 2 0 11 11 11 2 0 0 9 2
12 13 15 2 16 13 1 15 1 11 3 3 2
29 10 9 13 2 3 15 11 13 13 1 9 2 0 9 3 13 0 9 3 2 16 15 13 1 9 2 9 2 2
11 11 1 11 1 0 9 13 16 0 9 2
13 10 9 7 13 13 9 2 15 13 11 10 9 2
6 13 0 9 0 9 2
18 13 15 9 9 1 0 9 2 16 10 9 4 13 13 1 0 9 2
29 9 2 15 15 13 13 13 2 13 2 16 11 13 3 13 0 9 7 9 2 13 1 9 2 13 7 13 9 2
7 7 3 15 14 13 0 2
11 1 9 11 2 11 3 0 9 13 9 2
9 1 0 9 13 9 12 0 9 2
13 16 12 9 13 12 9 2 3 13 1 0 9 2
10 9 3 13 4 13 7 13 0 9 2
21 9 4 13 1 9 0 3 2 12 9 1 9 2 7 0 15 13 13 1 9 2
16 0 9 9 13 13 1 0 0 9 2 1 3 0 9 9 2
16 14 12 9 4 13 13 1 9 12 9 2 1 0 9 9 2
7 9 4 13 0 0 9 2
10 9 13 9 0 9 1 0 0 9 2
19 15 13 13 1 9 2 16 4 9 1 0 9 9 13 4 3 13 9 2
10 11 7 13 9 2 15 13 0 9 2
9 3 2 9 13 9 1 12 9 2
18 16 7 13 3 1 15 12 9 2 13 13 9 12 9 1 0 12 2
22 1 9 9 15 3 3 13 9 1 9 11 2 11 7 3 0 9 11 2 9 9 2
22 12 0 9 13 0 9 2 1 15 15 11 0 1 0 11 3 1 9 13 1 11 2
4 13 15 9 2
10 3 1 11 2 11 2 11 2 12 2
23 9 9 9 9 1 9 9 1 12 9 11 2 11 13 3 9 1 9 1 11 1 11 2
28 10 0 9 3 1 9 9 11 3 1 9 1 0 9 13 2 13 3 1 0 9 1 11 2 11 7 11 2
35 3 13 7 9 0 2 1 9 11 13 12 0 9 0 9 2 1 15 9 11 1 11 7 9 11 1 11 11 3 3 13 1 9 7 2
41 9 0 2 2 13 14 1 0 9 2 13 4 3 13 1 9 1 0 9 2 7 7 1 9 0 9 1 9 2 9 9 13 9 15 1 0 9 9 9 13 2
8 7 4 13 9 3 0 2 2
69 0 9 2 11 2 0 2 11 2 2 9 2 11 2 2 11 2 11 2 2 11 2 11 2 2 11 2 11 2 2 11 2 11 2 7 11 2 11 11 2 2 2 11 2 11 2 2 11 2 11 2 2 11 2 11 11 2 2 2 11 2 11 2 2 11 2 11 2 2
18 16 4 13 11 1 9 1 11 2 13 4 1 9 11 2 11 2 2
10 9 1 12 2 13 11 2 11 2 2
2 0 9
23 9 7 9 9 1 0 9 1 11 7 11 13 11 1 0 2 13 1 0 0 9 11 2
26 9 11 11 11 13 2 16 2 16 15 13 9 2 13 13 10 9 2 7 1 0 9 4 13 2 2
25 1 9 11 11 2 11 1 0 2 9 9 9 0 11 11 13 2 16 15 10 9 3 13 0 2
19 0 0 9 1 9 0 9 2 11 2 4 12 2 9 13 9 9 11 2
31 0 9 10 9 11 11 13 2 16 11 15 4 3 13 16 9 0 9 2 7 15 13 13 9 1 15 1 9 0 9 2
14 1 10 9 15 11 13 1 9 0 0 2 9 0 2
21 1 10 9 15 1 0 9 13 3 12 7 12 12 9 2 7 15 3 1 11 2
10 9 11 13 11 11 2 9 11 0 2
13 9 0 9 11 7 11 13 2 9 0 9 2 2
39 1 10 9 15 9 3 13 2 0 9 2 2 3 11 10 9 3 13 2 16 4 9 9 13 9 2 13 15 1 9 0 9 11 2 0 3 1 11 2
20 1 9 9 11 15 1 15 13 2 16 13 3 13 11 2 7 1 15 13 2
23 0 9 9 11 1 9 0 9 1 0 11 11 13 13 16 9 9 11 13 0 0 9 2
3 2 11 2
23 9 9 9 11 15 15 13 1 9 1 0 0 9 2 13 3 9 0 9 11 11 11 2
13 11 13 13 2 16 1 0 9 3 13 0 9 2
18 9 11 11 11 13 9 0 0 9 2 7 15 7 1 9 9 11 2
17 11 11 1 15 13 2 16 11 4 13 9 1 9 1 0 9 2
3 2 11 2
5 12 9 1 9 9
28 13 12 2 12 2 12 4 14 12 9 1 9 13 9 11 9 7 0 9 3 12 12 9 1 9 1 11 2
15 9 15 13 3 1 9 7 1 9 7 1 12 0 9 2
10 1 15 13 2 15 13 1 0 9 2
20 9 9 11 11 11 13 2 2 1 0 9 12 15 0 9 13 12 9 9 2
11 15 13 1 9 7 1 9 2 3 13 2
7 13 15 9 1 9 9 2
12 1 9 9 9 13 2 16 13 15 13 2 2
11 0 9 13 1 12 2 9 12 1 9 2
17 9 11 11 13 2 2 3 4 13 9 1 12 9 12 12 9 2
9 10 0 9 13 3 12 9 9 2
16 1 12 9 13 9 1 10 9 3 1 0 12 9 0 9 2
14 13 3 1 9 2 1 15 15 13 3 1 0 9 2
22 3 12 9 13 9 1 9 1 9 2 0 1 9 12 7 9 12 7 10 0 9 2
11 13 9 1 0 9 7 0 9 13 13 2
21 9 1 9 1 9 7 0 9 4 15 13 13 3 1 12 2 12 2 12 2 2
17 1 9 1 0 9 13 3 1 0 9 7 1 9 13 0 9 2
2 11 12
6 12 9 2 9 2 9
4 12 9 2 9
3 12 9 9
3 12 0 9
6 12 11 2 11 2 9
3 12 0 9
2 12 11
3 12 9 9
5 9 1 12 1 12
3 12 9 9
7 12 11 2 11 2 0 9
3 12 9 9
2 12 9
6 12 9 2 9 2 9
6 12 13 2 13 2 13
4 12 13 2 13
2 12 9
4 12 9 0 9
3 12 9 11
5 12 9 2 9 9
2 12 9
2 12 9
4 12 9 2 9
3 12 9 11
2 12 9
1 11
2 12 9
4 12 9 1 9
2 12 9
3 12 11 11
5 9 1 12 1 12
3 12 0 9
4 12 9 1 0
4 12 13 1 2
3 12 0 9
4 12 14 1 11
3 12 15 2
3 12 9 11
2 12 11
4 12 9 0 9
5 12 0 9 2 9
3 12 9 11
3 12 9 11
3 12 9 11
8 12 12 12 9 2 12 2 2
5 12 9 7 9 2
5 12 1 9 1 9
2 12 9
3 12 9 11
2 12 9
4 12 1 0 9
3 12 9 9
2 9 12
3 12 9 11
2 12 9
3 12 9 11
3 12 0 0
6 12 3 13 2 13 9
3 12 11 9
3 12 9 11
2 12 11
3 12 9 11
3 12 0 0
2 12 11
4 12 0 9 11
3 12 9 11
2 12 11
4 12 0 9 11
3 12 9 9
5 12 11 2 9 2
3 12 9 11
4 12 11 9 9
2 12 11
5 12 9 0 1 9
5 12 9 1 0 11
2 12 9
2 12 9
3 12 9 11
3 12 11 9
3 12 9 9
6 12 9 2 12 2 2
2 12 11
6 12 9 2 9 7 9
3 12 9 11
3 12 11 11
4 12 11 2 11
4 12 0 9 11
3 12 0 0
4 12 0 0 3
3 12 9 11
11 1 11 15 13 3 2 7 9 13 3 13
1 9
17 1 11 15 13 3 2 7 9 13 3 13 0 9 1 11 1 11
24 0 9 1 15 2 16 4 11 13 13 10 9 3 1 11 3 1 9 0 9 2 3 13 2
20 14 3 11 13 2 16 13 13 9 1 9 0 16 12 2 7 3 12 9 2
31 13 3 1 9 2 9 9 2 15 13 4 13 2 2 1 9 0 9 11 1 0 9 11 2 15 15 13 13 1 9 2
24 11 13 1 9 0 9 2 15 13 2 16 4 15 9 0 0 9 13 13 2 16 2 2 2
32 7 9 0 9 0 9 1 0 9 2 3 1 11 2 1 11 7 1 11 2 13 3 0 2 16 15 3 7 1 9 13 2
33 1 12 9 13 3 1 0 7 0 9 2 16 9 12 9 2 11 2 13 10 9 1 3 0 9 7 13 3 1 10 0 9 2
15 0 9 9 13 9 2 16 11 3 13 2 15 1 15 2
39 11 13 3 13 9 1 0 11 2 1 11 2 1 11 7 1 0 9 2 3 15 1 9 13 1 0 2 7 3 3 0 2 9 1 2 0 9 2 2
25 1 0 9 7 11 3 11 13 2 16 9 3 3 13 2 7 15 13 7 0 9 11 7 11 2
10 7 9 13 2 16 13 14 1 9 2
28 9 0 9 4 3 11 13 13 1 9 2 7 13 3 0 2 3 13 9 9 1 9 1 9 12 0 9 2
7 0 9 13 3 12 9 2
23 7 13 0 7 3 7 0 9 1 0 9 9 2 7 15 13 1 9 9 1 0 9 2
12 13 0 2 15 1 12 9 13 1 15 0 2
9 1 9 9 15 13 3 9 0 9
2 11 2
21 1 0 9 0 9 1 11 15 9 9 13 1 0 0 9 1 0 7 0 11 2
21 1 0 9 11 13 1 9 14 12 9 9 7 0 9 1 0 9 9 1 9 2
19 9 9 13 7 1 0 9 1 9 4 13 12 9 0 9 7 12 9 2
12 3 1 11 13 12 9 9 7 9 9 9 2
23 1 11 15 9 0 9 15 13 13 9 0 0 9 2 1 15 13 3 13 1 12 9 2
14 9 13 14 1 0 9 7 4 13 14 9 9 9 2
14 0 9 13 1 0 9 0 9 0 9 7 0 9 2
33 16 3 1 10 9 4 13 1 3 0 9 1 0 9 1 11 2 3 15 13 9 9 9 1 10 9 1 0 0 9 1 11 2
18 1 10 0 2 7 0 9 15 9 0 9 13 1 0 9 7 9 2
23 0 9 0 9 1 10 0 0 9 1 11 13 1 0 9 1 0 15 0 9 1 11 2
23 9 9 7 9 1 9 4 1 9 13 7 1 11 2 11 2 11 2 11 7 0 9 2
19 12 1 9 0 0 9 2 15 3 11 13 2 7 13 3 9 0 9 2
10 15 13 13 1 9 9 1 0 9 2
3 9 3 0
5 11 2 11 2 2
16 1 12 9 1 9 0 13 1 9 9 9 0 9 7 9 2
20 1 10 9 9 11 13 1 10 9 7 9 9 9 3 1 9 9 9 9 2
26 9 10 9 2 16 15 9 13 0 9 7 1 0 12 0 9 2 13 3 11 11 2 0 9 11 2
27 2 10 9 4 13 3 1 12 9 9 9 3 7 14 1 10 9 4 10 9 13 9 1 0 9 2 2
4 0 9 1 11
12 9 1 11 13 0 7 0 2 16 15 13 2
23 0 0 9 3 13 1 0 9 0 0 9 1 12 9 2 1 0 9 13 0 9 2 2
16 0 12 0 9 15 13 1 0 9 13 1 12 7 12 9 2
17 9 9 4 13 7 1 9 1 12 7 12 9 1 0 12 9 2
18 9 9 9 13 1 0 9 9 9 1 9 2 15 3 13 1 9 2
15 1 0 0 9 13 0 9 9 2 3 12 9 9 2 2
21 0 9 1 9 7 9 0 1 9 13 0 9 2 15 13 9 0 0 0 9 2
3 3 0 9
39 9 11 3 13 11 11 2 11 2 2 16 4 16 9 9 13 1 0 9 0 9 0 2 0 9 2 3 15 13 1 9 0 9 11 0 9 1 11 2
35 9 9 13 7 9 7 9 0 0 9 2 7 9 9 9 0 9 12 2 9 2 12 9 9 2 0 9 1 9 0 9 2 9 2 2
24 9 9 11 11 1 9 13 2 16 1 3 0 9 9 13 0 2 16 9 9 9 13 9 2
27 1 11 2 11 2 4 9 0 16 9 7 13 16 9 2 7 13 1 9 2 3 3 13 1 9 2 2
2 9 9
2 11 2
26 3 3 16 12 9 2 15 13 9 1 12 12 9 2 4 13 1 0 9 1 9 9 1 0 11 2
19 3 13 9 0 9 1 9 9 11 11 2 1 10 9 4 13 0 9 2
15 0 3 0 9 4 13 7 1 9 0 9 4 13 3 2
4 0 9 1 9
5 11 2 11 2 2
35 12 0 0 7 12 0 9 1 9 2 9 7 9 2 1 15 7 9 13 13 12 2 3 2 12 9 2 13 3 1 0 9 0 9 2
13 1 0 9 9 13 1 9 1 9 13 10 0 2
19 1 9 13 7 0 9 1 12 1 12 9 7 9 9 1 0 0 9 2
24 3 15 13 11 11 2 9 9 9 0 7 0 9 9 9 11 2 13 10 9 9 10 9 2
30 2 1 9 0 9 4 7 13 13 0 9 1 0 9 2 16 4 13 1 9 9 1 0 9 2 2 13 11 11 2
9 2 13 9 0 9 9 2 12 2
2 9 11
20 0 9 11 13 0 9 1 9 9 11 2 15 15 13 3 16 12 9 9 2
10 9 13 1 0 9 9 0 9 11 2
23 1 9 0 0 9 13 3 12 9 7 0 9 1 0 9 1 0 0 2 0 2 0 2
20 0 2 11 2 2 13 13 9 11 2 10 0 9 4 1 10 9 13 13 2
11 13 15 9 2 7 4 13 7 9 13 2
9 4 13 3 2 9 15 3 13 2
15 16 13 1 9 2 9 15 15 13 2 13 7 13 2 2
30 11 2 11 2 2 13 4 1 9 2 13 4 2 16 4 13 1 9 1 0 9 2 7 1 10 9 3 13 9 2
11 13 4 9 2 7 1 9 13 9 2 2
7 1 11 2 2 13 9 2
12 0 9 2 0 9 2 7 15 13 1 11 2
17 11 1 11 2 11 2 2 0 0 9 12 2 13 3 0 9 2
19 0 9 11 15 1 15 13 2 16 13 15 3 3 0 2 0 0 9 2
7 7 9 1 9 3 0 2
17 13 4 15 3 13 12 9 16 1 0 9 1 11 1 9 12 2
11 2 13 15 3 0 9 2 1 0 9 2
19 7 16 4 15 15 13 13 12 9 2 13 4 15 1 0 9 9 2 2
14 15 3 15 7 10 9 13 1 9 1 10 0 9 2
13 2 12 9 13 1 0 2 15 2 11 7 11 2
7 11 13 9 0 9 2 2
9 15 1 0 9 13 1 15 0 2
4 2 11 2 2
18 13 4 1 9 9 11 1 9 9 1 11 2 3 13 1 9 11 2
7 15 13 1 15 12 9 2
17 2 13 1 15 10 3 0 9 2 13 0 9 7 9 9 2 2
20 13 2 16 13 13 1 15 2 16 15 11 13 1 11 1 0 9 0 9 2
11 15 15 1 10 9 2 13 2 1 15 2
14 2 3 4 13 2 16 13 1 9 12 7 12 9 2
9 0 13 2 16 4 13 15 2 2
11 15 3 13 2 0 9 2 11 7 11 2
21 2 1 9 2 3 15 13 12 9 2 13 2 7 12 13 1 11 16 9 2 2
15 4 13 1 11 1 9 2 7 15 4 3 13 13 12 2
14 2 12 9 4 15 13 3 2 12 4 13 9 2 2
8 3 4 15 1 15 3 13 2
8 13 4 15 9 1 10 9 2
3 2 3 2
13 13 9 10 9 2 13 3 7 10 0 9 2 2
10 2 1 10 9 1 11 3 13 2 2
13 1 0 9 15 13 9 2 16 13 9 1 11 2
4 13 15 9 2
13 2 13 15 0 9 2 15 13 9 1 0 11 2
15 13 9 1 0 9 2 7 15 13 9 1 0 9 2 2
8 4 4 3 13 0 9 11 2
16 3 1 15 2 16 4 13 9 2 7 1 0 9 10 9 2
13 2 4 4 13 9 11 1 9 9 1 9 9 2
13 1 0 9 2 1 15 13 9 2 7 13 11 2
16 16 13 1 15 2 13 2 16 15 13 9 10 0 0 9 2
7 13 9 2 13 3 9 2
27 1 11 7 1 11 13 0 14 15 2 16 13 0 9 2 7 7 15 2 16 13 1 9 9 9 9 2
9 15 13 9 9 0 2 7 0 2
9 2 0 3 13 7 0 13 0 2
7 7 3 14 1 9 2 2
9 11 2 0 2 9 2 2 1 9
2 11 2
16 9 1 9 1 9 0 9 9 11 13 3 1 0 0 9 2
44 13 2 16 9 10 0 2 9 2 7 9 0 9 9 11 1 10 9 13 9 0 9 9 9 2 9 7 9 11 7 9 9 7 9 11 1 9 1 9 0 9 0 9 2
40 9 7 13 9 9 11 11 11 2 0 9 11 11 2 16 4 1 0 9 9 2 15 13 2 16 1 10 9 13 13 3 13 9 9 9 11 2 13 9 2
4 0 9 1 9
5 0 9 0 9 13
19 11 11 1 0 9 13 14 9 1 12 9 2 15 15 13 1 10 9 2
16 3 13 9 9 0 15 0 7 0 9 7 9 0 9 11 2
14 13 12 9 7 13 0 9 2 1 10 9 13 9 2
38 10 0 9 13 1 9 9 1 0 9 1 0 9 2 13 15 2 16 13 9 7 13 0 9 1 0 9 0 0 9 2 1 15 13 1 12 9 2
15 16 9 9 9 7 9 13 2 16 0 13 0 13 0 2
8 11 11 0 13 7 13 13 2
23 1 9 1 0 9 15 13 2 16 1 9 13 9 1 9 9 2 3 1 9 0 9 2
6 13 15 9 0 9 2
25 2 13 3 3 2 7 16 15 10 9 0 13 2 2 13 10 9 1 9 9 0 9 11 11 2
10 2 9 7 9 13 3 13 9 9 2
7 1 9 13 3 3 3 2
13 13 9 1 11 2 7 13 15 7 9 9 2 2
11 1 0 9 4 3 13 0 9 11 11 2
13 15 13 9 12 9 9 1 9 0 1 9 9 2
8 0 13 7 9 9 10 9 2
19 2 11 11 13 2 15 13 2 2 13 9 0 9 1 0 9 11 11 2
8 2 10 0 9 13 9 9 2
12 1 0 9 13 3 1 9 12 9 0 9 2
24 13 9 2 16 13 1 0 0 9 14 12 9 2 3 9 2 15 4 13 1 0 9 9 2
12 0 9 4 15 13 9 12 7 12 9 9 2
17 11 11 15 1 9 9 13 1 9 1 9 1 9 12 9 9 2
15 7 15 3 13 3 1 9 9 2 16 9 10 9 13 2
15 3 4 13 13 9 3 2 7 13 15 13 1 0 9 2
22 13 3 9 2 16 7 15 12 13 9 3 2 1 1 9 0 9 1 0 9 2 2
12 13 15 9 1 15 2 16 11 11 13 9 2
17 2 13 15 2 16 11 11 13 9 3 2 16 13 1 15 9 2
16 9 13 2 16 13 1 10 9 7 1 9 3 10 9 2 2
23 11 11 15 13 1 9 2 15 0 9 13 1 0 9 11 2 1 15 13 1 12 11 2
16 9 11 11 11 13 13 2 16 15 13 1 9 9 0 9 2
13 7 3 1 9 10 9 13 11 11 9 1 11 2
25 15 7 3 3 13 0 9 13 3 2 16 1 12 9 2 3 9 0 9 13 13 1 9 9 2
7 11 11 13 14 3 0 2
2 9 2
22 1 9 9 2 16 15 13 0 9 2 13 12 11 2 16 4 15 3 3 12 13 2
4 13 0 9 2
14 1 11 3 15 13 3 0 2 3 9 0 9 13 2
5 1 0 9 14 2
9 0 9 13 0 9 1 9 9 2
15 13 15 13 1 15 2 16 9 13 9 0 1 11 11 2
11 15 15 7 7 1 10 0 9 9 13 2
3 13 9 9
6 0 11 2 11 2 2
27 9 9 0 1 9 0 2 9 4 3 1 9 0 9 1 12 0 9 13 1 0 0 9 1 0 11 2
38 3 1 15 9 13 0 0 9 9 7 9 11 11 7 11 11 2 13 1 0 9 1 9 2 3 1 9 9 4 9 9 13 9 0 9 7 9 2
16 9 9 13 11 2 11 13 12 1 12 9 2 15 15 13 2
57 9 1 0 0 9 1 11 2 0 1 9 12 1 11 2 15 13 1 9 3 12 2 9 2 13 2 16 0 2 9 13 13 3 12 9 2 12 0 9 2 12 9 2 9 7 0 0 9 2 12 0 9 7 12 0 9 2
3 9 11 11
4 9 9 15 13
1 11
4 9 9 15 13
2 11 2
17 0 9 13 0 9 1 0 9 1 9 1 2 9 9 9 2 2
20 10 9 0 7 0 9 0 1 11 13 9 2 1 15 13 1 9 9 9 2
12 1 11 3 4 13 9 1 9 7 0 9 2
8 9 0 9 13 9 1 9 2
16 0 9 13 9 0 9 7 9 2 15 13 3 9 1 9 2
24 9 11 13 9 1 9 9 2 15 15 13 9 0 9 2 7 4 15 13 13 0 9 9 2
5 11 7 11 13 3
4 13 7 0 9
2 11 2
9 1 9 1 11 3 13 0 9 2
26 0 9 9 13 2 16 0 9 15 13 13 3 0 9 7 0 9 1 9 11 3 0 0 9 11 2
14 0 9 3 13 2 16 0 9 15 13 0 9 13 2
45 0 9 11 11 13 2 16 0 9 13 1 0 9 2 7 4 3 13 2 16 4 13 0 9 0 11 7 11 1 11 2 15 4 13 2 3 2 0 9 9 0 9 11 2 2
21 11 15 13 9 9 0 9 7 0 9 2 13 11 2 7 9 13 10 9 13 2
21 10 11 4 3 13 1 0 9 2 15 13 0 0 9 3 1 11 1 0 9 2
10 0 9 1 0 11 13 1 9 1 9
4 9 13 1 9
2 11 2
16 1 0 0 11 13 1 9 1 9 9 1 9 9 1 9 2
15 3 0 9 13 1 9 1 9 9 9 1 11 1 11 2
11 9 13 1 9 9 7 13 12 0 9 2
5 3 4 15 13 2
10 1 9 0 9 13 0 7 9 9 2
34 1 0 9 13 3 9 1 9 1 11 2 15 15 1 11 13 1 9 3 2 16 0 9 13 10 0 9 1 11 2 3 1 11 2
21 0 9 15 13 13 3 1 0 9 1 11 2 0 9 7 0 9 1 9 13 2
5 12 9 9 13 2
29 3 1 0 11 15 13 1 0 12 9 13 0 9 0 9 1 0 9 9 14 1 0 7 0 9 9 1 9 2
26 9 15 13 1 12 9 2 13 15 7 2 16 1 9 1 0 9 13 1 12 0 9 1 0 11 2
14 1 11 4 1 9 1 9 13 3 9 9 1 11 2
19 1 11 13 9 14 12 9 7 1 9 13 9 13 9 1 0 0 9 2
15 11 1 15 13 9 0 9 9 2 15 13 14 12 9 2
14 3 0 9 2 3 9 13 10 0 0 9 0 9 2
27 0 9 0 9 0 9 2 16 4 4 13 0 0 0 9 2 15 7 1 0 9 13 3 1 0 9 2
22 13 4 15 3 1 9 1 9 2 7 10 2 0 9 2 4 13 1 9 0 9 2
11 9 1 0 9 2 9 7 9 1 0 9
5 11 2 11 2 2
32 1 9 9 1 0 9 1 9 11 13 13 1 0 9 1 0 9 7 9 1 9 9 7 12 9 9 0 9 1 0 9 2
9 13 1 9 3 0 1 9 12 2
15 1 0 9 13 0 1 9 9 0 1 10 9 0 9 2
28 3 13 1 9 3 0 7 0 9 0 9 2 15 1 9 1 11 7 11 13 1 11 0 9 11 11 11 2
15 1 9 13 9 0 9 2 9 11 7 9 11 7 11 2
14 9 15 13 1 12 7 12 9 9 1 0 12 12 2
23 2 9 2 0 0 9 7 0 9 15 13 3 1 15 2 16 9 2 2 13 15 9 2
20 1 0 9 13 0 9 9 2 1 15 13 2 16 4 10 9 13 1 9 2
20 3 15 1 9 13 2 16 9 13 13 7 13 9 1 0 9 0 1 9 2
19 9 13 2 16 0 9 7 9 9 10 9 13 0 1 9 0 0 9 2
14 11 11 0 9 0 9 2 2 13 15 1 9 0 2
23 10 9 13 13 1 9 9 1 9 7 9 2 15 1 9 9 13 9 2 9 0 0 2
9 13 4 1 15 1 0 0 9 2
18 1 9 1 0 9 15 13 1 9 15 0 9 1 9 12 9 2 2
2 0 11
13 0 0 0 9 11 15 13 13 7 1 0 9 2
22 3 13 0 9 1 0 9 9 2 15 15 1 0 13 9 0 9 2 1 9 12 2
21 1 10 0 0 9 13 9 12 9 11 9 12 2 15 15 13 1 12 9 9 2
21 9 11 13 9 9 2 16 9 13 0 13 9 1 0 9 1 9 12 9 9 2
13 9 2 0 12 9 2 3 13 9 12 9 9 2
12 1 0 12 9 15 10 9 13 1 12 9 2
21 11 15 1 0 9 13 9 9 11 9 0 1 0 9 1 9 9 1 0 9 2
11 9 11 13 0 10 0 7 3 0 9 2
43 0 9 0 9 2 15 15 13 13 1 0 9 0 11 1 11 2 13 3 9 1 0 0 9 1 0 9 2 0 0 9 1 0 9 1 0 11 7 9 0 9 11 2
22 2 1 0 9 3 1 9 13 9 0 15 9 7 9 7 9 1 9 0 9 2 2
30 0 9 1 9 2 12 9 9 3 2 15 3 13 2 1 0 9 0 9 11 13 1 12 9 7 13 12 9 9 2
8 11 13 1 9 9 12 9 2
25 9 7 13 9 1 0 9 2 3 1 12 9 1 12 2 9 9 0 9 13 14 1 12 9 2
17 1 11 1 11 7 9 1 11 9 1 9 9 9 11 7 11 2
39 2 0 0 9 1 11 13 3 1 9 1 15 2 2 13 1 0 2 3 0 2 9 1 11 1 11 11 7 10 0 0 9 9 0 0 9 11 11 2
15 13 12 9 0 2 0 2 0 9 0 9 1 9 9 2
24 3 3 9 13 0 9 9 2 0 1 0 9 11 7 11 2 15 13 9 1 9 9 9 2
27 7 3 13 9 13 15 1 0 9 15 2 15 15 3 13 1 0 9 9 1 0 9 3 3 0 11 2
13 11 2 12 2 12 2 12 2 2 0 9 1 9
16 1 0 0 9 15 3 15 13 0 9 13 12 0 1 9 2
30 0 9 15 7 13 11 2 15 13 1 11 13 2 16 9 11 13 0 9 7 0 9 13 13 13 10 9 0 9 2
34 0 9 15 13 1 9 11 1 3 0 9 3 0 11 2 3 4 15 9 0 9 13 1 9 9 2 7 13 14 1 9 7 9 2
16 0 2 1 15 0 9 13 13 2 13 0 9 0 0 9 2
29 11 13 13 2 3 0 0 9 0 9 2 13 11 0 0 9 0 9 0 9 2 9 7 1 0 9 7 9 2
12 1 0 9 3 13 13 9 1 0 0 9 2
25 1 11 15 13 13 14 0 9 0 9 2 9 0 9 4 13 13 0 9 9 2 7 3 3 2
14 15 10 9 13 1 15 3 1 15 9 9 1 11 2
46 16 3 11 11 7 11 11 13 1 12 9 2 9 0 9 1 0 9 13 0 9 3 0 9 0 2 0 9 2 15 3 3 13 9 11 11 11 16 9 1 0 11 1 0 9 2
41 13 4 3 1 2 0 9 2 2 10 9 0 9 2 1 12 0 9 1 0 9 2 1 12 0 9 1 0 9 2 1 12 3 0 9 7 1 10 0 9 2
11 10 15 13 13 0 9 11 2 1 9 2
26 1 9 9 11 2 16 13 1 3 0 9 7 0 9 3 2 13 9 11 2 13 15 7 1 9 2
28 9 10 9 4 13 7 11 11 2 16 15 1 11 11 13 1 9 9 7 13 15 2 1 15 13 3 9 2
14 12 0 9 3 13 1 3 0 9 0 2 0 9 2
13 3 7 3 13 1 0 9 1 9 11 7 11 2
16 11 11 13 9 1 9 7 13 9 1 11 2 15 13 9 2
37 11 11 15 1 0 9 3 13 7 1 15 1 0 9 3 13 9 2 16 0 9 1 0 2 0 9 13 1 9 10 9 1 3 0 9 3 2
32 7 3 2 16 1 9 0 9 13 12 9 1 9 7 0 9 2 13 9 11 9 1 9 2 16 1 10 0 9 13 9 2
26 11 3 3 13 9 1 0 9 2 7 15 3 15 3 13 0 2 16 11 1 9 13 1 0 9 2
18 1 9 0 2 1 15 15 12 9 13 2 13 2 16 9 13 13 2
12 11 2 12 2 12 2 2 2 9 2 9 0
19 1 12 9 3 13 9 11 1 0 9 1 0 9 11 13 9 7 9 2
22 1 10 9 4 9 12 9 13 2 0 0 9 7 13 1 0 9 9 10 0 9 2
34 13 15 2 3 1 11 13 10 9 2 3 1 9 13 0 9 0 9 2 16 4 13 0 9 11 2 1 15 1 11 3 13 9 2
31 16 15 13 1 9 0 0 9 2 15 13 9 0 9 2 11 11 15 3 13 1 10 9 0 9 1 9 12 0 9 2
19 13 3 9 11 11 2 16 10 9 4 14 13 9 9 7 3 0 9 2
15 3 7 10 9 13 7 3 15 1 0 9 13 11 11 2
14 0 9 2 9 0 9 2 1 0 9 13 14 3 2
19 15 15 13 1 9 1 9 0 9 2 9 2 9 2 9 2 0 9 2
25 10 9 15 3 13 1 0 9 1 9 9 1 12 9 2 13 1 9 2 0 9 2 0 9 2
24 0 4 1 9 11 13 3 3 2 11 13 3 0 9 1 0 9 1 11 7 0 0 9 2
5 9 9 13 0 2
41 2 1 12 9 13 9 7 3 0 9 2 0 1 0 9 11 2 13 1 12 1 9 11 11 2 16 15 13 9 2 13 15 3 9 7 13 3 1 9 2 2
29 0 9 13 2 16 9 0 0 9 11 7 2 9 2 0 0 9 1 0 9 13 9 0 2 1 15 13 13 2
26 3 11 11 13 2 13 15 2 16 1 15 13 2 15 15 13 2 7 10 9 15 13 1 15 13 2
17 1 0 9 15 9 11 3 13 16 4 9 13 3 10 9 13 2
28 1 12 9 3 11 11 13 0 9 1 9 10 9 2 1 15 15 13 9 1 9 7 0 9 12 0 9 2
27 1 9 2 15 9 11 3 13 1 9 2 13 1 0 9 0 9 7 3 3 9 1 0 9 1 9 2
33 0 10 9 13 9 11 9 2 16 16 4 10 9 13 2 13 11 1 12 9 0 9 7 0 9 13 1 11 13 3 16 3 2
9 0 7 0 13 7 9 0 9 2
30 11 11 15 13 1 9 11 1 9 9 7 1 1 9 1 11 11 2 3 4 13 3 1 9 11 2 13 1 11 2
23 0 9 3 13 10 0 9 2 15 13 3 3 1 11 2 11 11 11 13 1 10 9 2
42 14 1 10 12 9 2 7 7 1 0 9 2 1 15 3 13 9 2 7 3 9 11 13 3 1 9 2 16 13 10 0 0 9 1 9 9 2 15 13 0 9 2
31 1 12 1 9 3 11 11 13 3 9 2 16 13 13 2 16 0 9 13 1 10 9 7 10 9 13 1 9 2 2 2
23 7 16 4 13 10 9 2 13 2 13 2 9 9 2 16 15 4 15 1 10 9 13 2
11 11 2 12 2 12 2 2 2 2 2 2
3 7 9 13
11 9 1 0 0 9 13 9 0 0 9 2
43 9 11 1 15 13 13 13 0 9 2 16 4 13 9 2 7 13 0 9 1 0 2 0 11 2 7 13 0 9 1 3 0 9 2 15 13 9 9 1 12 0 9 2
24 3 15 1 9 13 1 10 0 9 2 1 15 13 0 9 9 7 10 9 1 0 0 9 2
20 16 4 0 9 3 13 10 0 9 2 13 11 13 9 1 9 0 9 13 2
32 11 11 9 11 13 2 16 4 12 13 1 0 9 2 7 15 13 9 3 3 2 16 12 9 3 1 9 13 1 0 9 2
9 10 9 4 1 9 11 3 13 2
14 11 11 3 3 13 2 16 11 11 13 9 0 9 2
19 1 0 9 1 9 0 9 3 3 7 3 13 9 11 1 0 0 9 2
25 7 15 3 3 2 16 10 0 9 11 11 13 9 13 2 16 9 0 11 13 1 0 9 11 2
29 11 11 1 12 9 13 2 16 0 9 13 9 1 0 9 2 7 13 15 9 11 2 13 0 9 2 7 13 2
12 3 3 13 11 11 0 9 2 0 1 15 2
25 3 15 1 10 9 7 13 2 16 10 9 15 10 3 0 9 13 2 12 9 13 12 0 9 2
15 3 3 15 11 11 13 13 9 11 7 13 15 0 9 2
17 9 1 9 9 1 11 7 11 1 0 9 3 3 13 3 0 2
19 3 15 13 1 9 2 7 0 9 1 9 13 0 9 1 9 9 9 2
17 3 0 1 9 11 13 0 9 1 9 9 9 9 11 0 9 2
13 2 13 15 3 0 0 9 1 9 9 9 2 2
22 3 3 13 3 11 11 13 9 2 16 4 3 3 13 1 0 9 9 0 0 11 2
34 7 3 0 9 1 9 9 2 1 10 9 3 3 11 0 3 13 2 16 13 3 0 2 7 0 16 10 0 2 13 13 9 11 2
20 3 1 0 9 1 9 0 9 13 10 9 0 9 13 2 13 4 11 3 2
22 13 11 11 1 0 9 0 1 9 0 9 0 9 3 13 0 0 9 10 9 2 2
32 1 0 9 1 0 0 9 13 9 11 1 15 2 16 0 9 4 13 13 3 7 0 9 2 15 13 3 0 9 11 11 2
3 11 11 2
2 11 11
4 9 2 11 2
2 11 11
2 9 11
2 0 11
15 9 0 15 9 9 13 9 1 3 0 9 1 9 9 2
9 13 7 13 11 11 1 9 1 11
7 9 2 2 12 2 12 12
6 9 2 12 2 12 12
3 0 9 9
9 11 2 9 2 1 9 2 0 2
3 13 9 2
3 3 13 2
9 9 2 1 11 13 3 7 3 2
11 0 9 12 7 12 2 0 12 7 12 2
9 2 1 11 13 13 3 7 3 2
12 0 9 12 7 12 2 0 12 7 12 2 2
29 1 9 13 9 12 2 12 7 13 1 12 2 12 2 9 13 1 9 1 12 2 12 7 13 1 12 2 12 2
20 9 9 2 0 9 12 9 11 13 1 9 12 2 0 12 9 1 9 12 2
8 0 0 9 13 12 9 11 2
12 0 9 2 0 9 0 2 0 9 3 0 2
2 0 9
15 0 9 2 1 10 9 1 15 4 13 0 9 1 9 2
9 7 0 9 4 13 13 3 0 2
16 13 15 3 0 9 2 3 7 1 9 9 9 2 3 9 2
11 0 9 12 7 12 2 0 12 7 12 2
2 0 11
28 1 9 1 9 0 9 1 0 11 13 0 2 9 11 11 2 12 2 12 2 12 2 1 9 9 0 9 2
30 9 1 12 9 0 9 13 11 1 11 2 12 2 12 2 12 2 7 0 13 11 11 2 12 2 12 2 12 2 2
43 0 9 2 9 9 2 12 9 2 2 12 2 11 2 11 2 12 2 12 9 2 12 2 11 2 12 11 2 12 2 12 2 12 2 11 2 11 2 2 12 2 12 2
3 11 13 9
2 1 9
2 11 2
14 9 1 9 2 9 2 11 2 11 2 2 2 2 2
8 12 2 11 2 9 2 11 2
9 9 2 11 2 11 2 2 2 2
17 12 2 11 2 11 2 12 2 12 2 12 2 9 2 11 2 2
4 0 11 15 13
28 11 11 2 12 2 11 11 2 13 1 0 9 9 1 11 2 12 2 12 2 9 7 13 1 12 2 9 2
25 3 3 7 0 9 1 11 13 7 3 15 13 1 9 0 2 9 1 11 1 9 1 0 9 2
5 15 15 3 13 2
18 2 1 0 9 4 13 3 1 9 9 12 1 9 7 13 15 9 2
24 13 9 7 13 15 3 2 7 3 1 9 2 3 13 0 9 2 15 9 9 13 12 9 2
32 13 15 2 16 4 13 13 13 2 7 9 13 0 9 2 3 13 0 1 0 9 2 7 1 15 3 7 1 15 1 11 2
8 16 15 3 13 1 11 2 2
4 0 9 11 2
31 9 11 1 10 9 13 2 16 0 9 11 1 11 13 12 0 9 2 15 15 4 3 13 9 9 0 0 9 9 11 2
21 11 11 13 2 16 9 10 9 13 0 1 9 9 7 16 9 13 0 9 11 2
8 1 9 3 13 1 0 9 2
20 11 16 0 0 0 9 1 11 13 2 3 1 9 1 11 2 9 1 9 2
27 10 0 2 9 2 0 9 1 11 3 0 0 9 1 11 13 1 9 2 16 4 13 0 13 9 9 2
20 9 11 11 2 16 16 13 13 9 9 9 2 13 13 9 2 3 15 13 2
15 3 15 13 7 3 0 2 13 2 14 1 9 9 11 2
21 15 0 2 16 14 15 7 10 9 2 4 13 13 1 9 0 9 1 9 9 2
21 16 15 0 0 9 1 9 13 13 2 0 9 2 2 3 15 3 0 9 13 2
26 7 13 3 3 12 9 2 15 3 13 1 9 11 11 2 7 3 2 16 11 13 13 3 3 13 2
3 9 13 9
6 0 11 2 11 2 2
31 9 1 9 0 0 9 9 9 7 9 1 9 11 1 0 9 7 9 13 11 11 2 9 0 9 7 9 9 9 0 2
26 9 9 7 1 0 9 1 9 2 15 4 13 9 9 9 2 15 13 3 9 2 13 0 0 9 2
23 0 9 0 9 9 2 0 1 9 9 9 7 9 2 13 1 0 9 0 0 9 9 2
9 15 4 15 3 0 9 13 9 2
35 2 13 1 15 2 16 4 9 9 9 13 15 2 15 10 9 1 9 9 9 13 1 0 9 1 0 9 2 2 13 3 11 2 11 2
24 1 10 9 4 9 13 13 1 9 7 9 1 9 9 0 9 2 7 15 7 0 9 9 2
3 0 9 14
14 11 11 2 11 2 2 13 13 9 2 15 15 3 13
18 16 9 0 9 4 13 9 9 1 9 9 9 3 1 15 0 9 2
10 13 3 7 9 7 9 0 0 9 2
5 10 13 9 9 2
15 2 1 9 2 15 13 1 0 9 2 15 13 3 3 2
24 7 3 2 1 9 10 9 2 7 1 10 9 2 3 15 9 13 13 3 0 2 4 13 2
25 1 9 15 7 13 0 9 2 1 9 3 9 10 0 9 13 0 9 2 15 7 0 9 13 2
28 2 3 15 13 2 16 15 9 2 14 1 9 2 4 13 1 15 2 16 4 15 13 0 9 9 0 9 2
26 15 3 13 1 15 2 16 4 15 13 9 2 16 4 15 13 0 9 2 15 13 3 1 9 2 2
13 13 7 13 7 1 15 2 16 9 9 9 13 2
8 2 13 4 15 1 9 9 2
24 13 15 9 2 16 13 13 1 9 0 11 2 1 0 9 2 15 13 3 7 1 9 0 2
13 3 13 13 10 9 2 15 3 15 3 13 2 2
5 15 4 3 13 2
8 2 13 4 15 0 9 2 2
14 15 3 7 13 9 9 3 9 0 9 16 9 11 2
7 2 13 15 1 0 9 2
8 0 9 13 0 1 3 9 2
16 1 0 9 13 0 9 2 16 4 4 13 0 9 1 9 2
22 1 0 7 3 2 16 0 9 1 9 9 9 13 9 9 9 16 12 1 12 9 2
18 7 0 9 1 9 13 1 9 9 2 14 2 1 9 9 9 2 2
9 7 9 0 9 13 3 3 13 2
8 15 4 15 13 0 9 15 2
12 2 13 0 3 13 15 0 9 1 0 9 2
10 3 4 15 13 1 10 9 7 3 2
16 0 9 4 13 3 13 10 3 0 9 1 9 10 9 2 2
38 1 9 7 10 9 13 2 16 9 1 9 9 9 13 0 2 16 0 9 1 9 12 13 2 16 11 13 13 1 0 9 2 7 10 9 13 13 2
14 2 9 9 1 9 9 3 9 11 13 1 9 13 2
19 10 9 0 9 9 13 0 2 16 15 13 3 1 9 0 9 1 9 2
7 11 7 1 9 13 2 2
15 16 4 3 4 13 9 0 9 2 13 4 9 0 9 2
4 2 3 2 2
28 7 16 4 9 1 10 9 13 2 14 2 2 13 15 2 16 13 9 9 9 13 3 1 9 10 0 9 2
18 2 13 4 1 0 9 2 16 9 9 4 4 13 3 9 9 2 2
18 3 4 7 13 4 13 0 0 9 2 15 3 13 9 7 13 9 2
18 15 13 2 16 1 9 9 0 9 9 4 9 13 1 10 0 9 2
7 2 11 13 9 1 9 2
21 3 9 3 0 9 2 14 3 2 3 13 0 1 9 7 1 9 9 7 9 2
32 13 9 9 2 15 4 13 9 9 7 1 0 9 2 1 15 2 16 13 3 13 2 13 1 11 1 9 2 15 15 13 2
21 13 9 2 16 4 3 13 0 9 1 10 12 9 2 16 4 3 13 0 9 2
35 14 2 10 0 9 13 3 1 9 2 7 13 15 13 10 0 9 2 16 15 13 3 2 16 4 9 13 1 9 12 7 0 9 2 2
37 13 7 9 2 16 1 9 0 9 15 9 13 9 0 9 7 0 9 9 11 15 13 1 10 9 2 9 2 16 11 3 13 9 1 9 9 2
8 2 0 9 1 9 15 13 2
6 0 9 13 0 2 2
4 13 15 11 11
4 9 2 11 2
2 11 11
4 0 9 1 11
4 9 0 0 9
2 11 2
21 3 0 0 0 9 2 11 2 13 1 11 10 0 9 2 15 13 1 0 9 2
19 1 9 0 9 11 13 9 9 9 1 9 9 7 1 9 9 1 9 2
32 3 13 9 11 11 11 2 13 10 9 1 2 0 9 0 11 2 7 1 0 9 11 13 4 0 0 9 13 0 0 9 2
27 9 0 9 1 9 9 11 11 13 2 16 10 9 3 13 3 16 12 0 9 1 0 7 0 0 9 2
18 1 0 9 9 3 0 9 1 9 13 1 10 9 9 1 11 13 2
6 1 9 0 9 15 13
8 11 2 1 10 0 9 2 2
29 0 9 13 0 9 2 1 9 0 9 1 9 2 1 10 9 0 0 9 1 9 1 9 9 0 9 11 11 2
8 15 9 0 9 14 3 13 2
15 10 9 2 1 0 9 7 9 2 15 14 13 0 9 2
62 2 13 3 3 13 2 16 1 0 7 3 1 0 11 4 9 9 1 9 0 9 13 0 9 2 7 9 0 9 2 10 9 4 13 2 7 9 9 0 9 2 0 9 7 9 9 7 9 1 9 0 9 2 15 4 13 0 9 2 2 13 2
18 10 11 11 3 13 9 0 9 11 1 2 0 9 1 0 9 2 2
44 9 0 9 1 11 3 13 2 3 1 10 9 13 2 2 14 0 9 1 9 2 7 7 1 15 0 9 9 1 11 13 1 9 0 9 2 13 1 0 9 0 9 2 2
41 1 10 9 13 3 0 7 0 9 0 1 9 10 11 2 15 1 9 13 1 9 2 15 13 10 9 2 2 13 1 15 13 3 1 9 11 2 3 0 11 2
11 1 9 0 9 15 3 3 3 13 2 2
46 0 9 9 11 11 11 3 13 1 11 10 9 2 16 0 0 2 14 2 4 4 4 2 13 1 9 9 2 1 0 0 9 11 2 3 15 3 13 9 2 3 13 0 9 2 2
28 3 15 13 2 16 1 11 2 9 11 2 11 2 3 13 0 0 9 2 13 0 9 9 1 9 12 9 2
11 10 9 10 9 13 1 0 2 14 2 2
17 13 4 1 15 1 9 3 7 1 9 9 11 1 0 9 11 2
44 3 0 1 15 3 13 2 3 13 2 14 2 2 7 13 15 1 0 9 12 9 2 2 2 13 2 16 4 15 3 3 3 13 9 1 9 1 12 9 9 7 0 9 2
14 1 11 15 3 13 7 1 0 9 3 16 3 3 2
13 7 15 13 7 1 10 9 1 11 2 11 2 2
47 7 3 15 1 11 2 11 13 15 2 15 1 0 9 11 3 13 2 0 9 3 1 9 9 7 9 0 9 13 2 9 1 14 2 2 1 10 9 15 13 0 9 0 9 11 11 2
24 3 9 9 7 1 15 3 0 9 7 9 13 9 1 9 2 15 13 1 2 0 11 2 2
27 15 7 16 9 10 0 9 1 9 13 0 9 2 1 0 0 9 2 15 4 15 3 13 13 1 9 2
20 0 9 0 9 2 1 15 13 12 2 9 12 11 2 3 13 0 0 9 2
31 16 4 3 13 1 15 2 16 4 15 0 9 13 1 9 3 1 12 2 9 12 2 1 15 13 7 1 11 0 9 2
24 0 0 9 15 3 13 2 16 0 9 11 11 13 1 0 9 1 0 9 10 3 0 9 2
3 11 1 9
2 11 2
24 2 1 9 2 16 4 13 1 9 9 2 4 15 1 9 0 9 10 9 13 3 12 9 2
28 10 9 13 3 0 1 15 2 16 4 13 1 9 9 2 2 13 3 1 11 9 0 9 9 11 11 11 2
14 0 9 13 9 0 9 7 9 15 13 2 9 13 13
30 0 9 0 9 3 0 9 9 13 9 2 15 13 0 9 1 9 9 9 1 9 7 9 2 7 9 1 9 2 2
34 3 15 3 13 9 3 15 0 9 13 9 10 9 7 3 3 13 1 0 9 9 9 12 2 12 9 2 1 9 12 2 9 12 2
33 1 10 9 15 3 13 9 2 3 3 9 7 9 13 0 1 9 0 3 1 9 2 15 0 9 10 3 0 9 3 15 13 2
21 3 1 9 14 12 9 2 1 15 4 1 0 9 13 9 1 9 1 10 9 2
37 9 13 3 0 2 9 15 0 9 15 3 13 13 3 1 15 2 7 1 9 9 9 2 15 4 13 1 0 9 9 2 13 3 15 1 15 2
20 9 13 3 7 1 10 9 3 0 9 2 9 9 13 13 10 0 9 2 2
29 9 7 1 10 0 9 13 3 0 9 1 9 9 2 3 9 2 9 9 13 1 0 9 10 9 1 9 9 2
7 7 3 13 1 15 13 2
27 1 0 0 9 0 9 13 3 12 9 0 0 9 7 3 1 9 0 9 2 16 13 9 1 0 9 2
6 15 0 15 9 13 2
13 7 13 15 15 3 7 9 9 1 9 7 9 2
30 0 9 0 9 9 4 13 1 12 9 9 2 15 13 9 14 12 12 0 9 9 0 9 7 9 1 10 9 0 2
14 9 9 7 13 2 16 1 3 0 9 13 13 9 2
34 3 7 7 0 9 13 3 3 1 9 2 16 3 0 9 9 9 1 9 3 12 9 9 0 9 9 0 9 13 0 7 0 9 2
18 2 3 15 10 9 13 2 2 13 3 0 0 9 1 9 0 9 2
21 1 0 9 0 9 9 1 9 13 3 0 2 1 15 15 3 13 3 15 0 2
29 3 0 9 1 10 9 13 14 3 2 3 15 2 15 13 1 9 3 0 9 9 2 13 1 9 9 1 9 2
30 16 9 13 9 9 7 9 9 1 9 9 2 15 4 1 9 13 1 0 9 9 2 13 10 9 1 0 9 9 2
26 10 9 15 1 9 13 9 7 7 10 9 2 15 3 13 0 9 9 2 4 13 16 0 1 9 2
34 1 0 9 9 7 9 13 2 16 15 3 13 9 1 9 0 1 9 9 9 7 1 9 10 0 9 2 0 15 1 0 0 9 2
25 0 9 9 1 9 13 9 9 7 10 9 3 2 16 4 4 13 9 9 3 2 7 3 3 2
15 1 9 2 15 4 13 9 2 15 3 3 13 0 9 2
23 1 9 0 9 9 7 0 9 4 3 3 13 0 9 9 14 12 12 9 14 1 11 2
22 0 9 13 1 15 2 16 0 9 9 1 0 9 4 1 10 9 13 3 9 9 2
12 3 3 13 9 0 1 0 9 9 0 9 2
26 0 9 9 1 9 1 9 13 14 3 2 0 9 3 13 9 2 15 3 13 0 9 0 0 9 2
48 15 7 13 0 9 14 10 9 1 0 9 12 2 9 2 9 13 1 12 9 2 2 10 9 15 7 13 10 2 0 2 9 2 15 9 9 1 12 2 9 14 1 9 9 13 1 0 2
30 7 9 2 3 3 0 2 13 0 9 2 13 0 9 10 9 9 1 9 7 9 2 15 4 13 1 9 12 9 2
18 1 11 1 11 7 9 1 11 9 1 9 9 9 11 7 11 2 12
23 1 0 9 4 15 13 13 2 15 15 3 13 1 0 12 9 0 9 1 11 7 11 2
18 7 1 15 13 3 3 0 2 16 15 12 9 9 13 13 0 9 2
24 13 11 11 0 1 0 9 13 0 0 9 0 9 2 15 4 13 10 9 1 9 9 9 2
15 15 13 15 2 16 1 12 9 15 3 13 9 0 9 2
26 0 1 0 3 13 13 2 16 0 9 11 7 11 13 1 0 9 0 1 9 0 9 1 12 9 2
22 3 1 9 15 11 11 13 9 11 11 2 15 1 9 11 1 15 16 0 9 13 2
23 0 11 15 7 3 3 13 2 16 1 9 4 13 1 9 11 13 1 9 0 0 9 2
27 7 3 1 9 10 9 15 3 13 9 15 2 16 11 11 13 14 1 3 0 11 11 16 0 1 0 2
33 9 11 10 9 13 1 0 7 15 2 16 13 0 13 1 0 9 3 0 0 9 2 7 15 3 3 7 1 9 0 0 9 2
12 11 2 12 2 12 2 12 2 2 11 13 9
21 10 9 2 0 3 0 0 9 2 15 3 13 1 9 3 2 16 4 3 13 2
10 7 15 3 1 0 0 9 11 11 2
14 15 7 13 2 16 1 9 11 3 13 1 0 9 2
31 1 12 1 10 0 3 11 11 13 2 16 16 4 13 9 9 9 11 7 10 9 0 9 2 13 11 1 0 0 9 2
29 10 9 1 11 13 3 0 9 9 1 12 9 2 15 3 12 7 9 9 13 1 9 9 11 11 7 11 11 2
21 0 9 3 7 3 13 10 9 7 15 15 3 13 9 1 9 2 16 13 9 2
22 3 1 9 9 11 2 16 3 9 13 0 0 9 9 2 15 15 13 1 9 9 2
12 3 10 0 9 11 1 12 14 3 0 9 2
21 3 0 9 7 9 1 10 9 13 9 11 3 1 9 0 9 0 9 11 11 2
29 15 0 9 7 9 2 15 11 11 13 1 15 12 9 9 1 11 2 13 2 16 12 10 9 13 0 0 9 2
34 11 11 13 3 13 2 16 15 11 3 1 0 9 13 7 13 1 15 0 9 3 1 9 12 2 3 1 9 10 9 1 0 9 2
25 3 1 10 0 9 1 3 0 9 1 15 7 0 11 13 0 9 1 11 7 3 7 0 9 2
19 13 3 9 2 16 9 1 11 11 3 13 2 7 3 1 9 11 11 2
39 3 7 1 0 9 1 11 11 11 13 1 9 10 0 3 0 9 2 3 13 1 9 9 11 7 13 9 9 11 11 0 1 9 9 9 0 2 9 2
15 3 13 9 11 13 2 15 15 15 3 1 10 9 13 2
32 3 1 9 1 3 12 0 9 4 13 9 9 2 15 4 1 9 0 9 1 9 13 13 1 0 9 9 1 9 10 9 2
32 1 0 9 13 7 9 0 0 9 2 15 4 13 3 3 2 16 15 12 9 13 3 13 2 1 15 15 1 15 4 13 2
31 1 15 0 13 1 11 9 2 1 15 11 11 2 16 15 1 15 15 13 2 13 9 0 9 11 2 12 2 9 12 2
31 3 9 2 16 9 11 3 13 1 0 9 1 0 9 2 13 11 2 16 0 9 3 13 1 9 7 3 7 13 13 2
32 7 3 13 9 11 11 11 1 10 3 0 9 1 9 11 3 13 2 2 0 0 9 1 11 13 3 1 9 1 15 2 2
2 0 9
31 16 13 9 1 0 9 0 9 2 13 1 0 9 2 3 14 1 12 2 9 13 9 12 9 0 2 0 9 0 9 2
32 1 9 13 9 11 11 2 11 11 2 11 11 7 11 11 2 3 15 0 1 9 2 15 15 3 13 13 1 9 0 9 2
24 15 9 15 3 3 13 1 0 9 2 7 3 13 1 0 9 0 9 2 13 3 3 13 2
18 15 15 9 13 2 7 13 15 3 3 0 9 2 15 0 9 13 2
13 15 3 2 15 3 2 13 15 0 2 0 9 2
18 1 10 0 9 13 1 15 1 10 9 9 12 3 3 3 0 11 2
17 16 3 13 1 9 2 9 7 11 2 9 13 3 0 0 9 2
10 13 15 7 9 3 0 1 10 9 2
7 10 9 13 0 9 9 2
31 13 13 0 9 1 0 9 16 0 0 9 2 0 9 15 13 1 0 9 2 3 13 9 1 0 13 13 9 2 2 2
7 14 2 13 15 0 9 2
20 0 9 9 1 11 3 13 7 11 11 2 10 0 9 15 13 1 9 0 2
5 13 0 2 0 2
5 7 3 3 0 2
7 3 0 11 11 13 9 2
34 10 0 9 9 2 13 15 2 11 2 13 15 13 0 14 9 2 15 4 15 3 1 0 9 13 2 7 0 9 2 15 3 3 2
4 0 9 0 9
47 9 0 2 15 1 0 9 13 3 1 12 12 15 9 9 9 1 10 9 9 0 0 7 0 9 2 11 2 2 15 1 9 9 13 1 0 9 2 1 15 15 13 1 9 3 0 2
15 10 0 9 15 13 3 1 10 0 9 1 9 0 9 2
45 2 10 0 9 15 1 9 0 13 2 7 1 9 0 9 7 9 1 9 13 2 16 9 1 12 9 1 9 9 4 13 4 13 2 2 13 15 3 9 0 9 11 11 11 2
22 2 9 0 13 1 10 0 9 3 3 13 2 16 4 3 1 15 13 13 3 15 2
18 9 1 3 0 9 15 13 1 9 13 3 1 10 0 9 1 9 2
9 9 0 13 0 1 9 7 9 2
27 1 0 9 4 13 9 14 1 9 1 12 0 9 1 9 2 7 3 4 13 2 16 13 1 0 9 2
17 3 13 9 7 1 0 0 9 2 10 9 15 13 3 13 2 2
22 9 13 9 9 0 9 2 2 3 13 2 13 15 15 13 2 2 13 9 11 11 2
13 2 9 13 13 9 2 9 7 0 2 0 9 2
28 1 9 1 9 2 3 4 1 9 1 9 13 9 13 1 0 9 9 7 0 9 2 1 0 15 13 2 2
5 13 0 0 9 2
12 9 3 13 1 12 1 12 9 9 1 9 2
22 2 9 13 12 9 2 16 16 13 9 13 2 15 13 2 13 4 15 3 13 3 2
10 3 1 0 9 13 9 1 9 2 2
36 1 0 9 0 9 13 11 11 2 2 1 9 13 13 11 2 7 13 13 2 16 9 4 13 3 1 15 2 16 15 3 10 9 3 13 2
23 13 9 3 2 3 9 13 1 9 0 9 7 9 13 9 0 9 12 7 9 0 9 2
22 1 9 13 0 9 9 2 3 15 9 13 3 1 0 9 2 3 13 1 0 9 2
15 13 1 9 2 7 9 13 0 2 9 13 1 9 2 2
3 12 0 9
12 3 1 11 9 1 9 12 2 11 2 0 9
29 16 0 0 9 13 3 1 11 1 10 0 0 9 1 9 12 1 9 9 2 0 9 2 13 10 9 3 0 2
10 1 0 9 15 3 3 13 13 9 2
19 7 3 0 2 16 15 13 13 2 13 0 9 1 3 0 9 0 9 2
11 9 13 1 12 9 7 13 15 11 11 2
8 15 3 2 16 9 13 9 2
25 9 0 9 11 2 12 2 2 2 13 0 9 16 0 9 1 9 2 16 9 13 0 3 3 2
12 7 15 14 3 2 16 10 9 3 3 13 2
11 13 15 1 15 0 9 2 13 1 9 2
28 7 0 9 13 1 15 0 0 9 9 2 9 15 1 15 3 13 7 13 13 2 16 3 4 13 3 3 2
15 13 3 9 2 7 1 0 9 13 1 9 1 9 2 2
14 9 11 10 9 13 2 13 15 12 3 0 9 9 2
16 16 13 10 9 2 3 15 1 3 0 9 13 1 0 9 2
17 1 10 9 3 0 9 13 13 2 1 10 9 14 13 1 9 2
14 15 9 9 9 15 14 13 13 9 14 1 0 9 2
22 10 9 11 2 1 9 1 9 1 11 2 3 13 2 10 2 0 9 9 0 9 2
32 1 9 13 9 2 1 0 9 14 1 0 9 2 7 3 2 16 1 10 3 0 9 13 13 9 0 9 2 2 2 2 2
9 10 9 9 4 13 11 1 11 2
10 9 1 9 3 13 0 0 9 11 2
19 13 2 16 15 4 9 0 9 13 3 2 16 15 13 1 9 1 11 2
9 13 15 3 9 1 11 7 0 2
30 1 9 9 11 1 0 13 9 2 15 15 13 1 10 0 9 2 16 3 1 9 1 11 13 1 0 9 11 9 2
18 1 9 11 3 2 16 1 10 9 13 2 13 9 11 2 16 3 2
8 9 11 2 11 2 12 2 2
50 11 2 12 2 2 11 2 12 2 2 11 2 12 2 2 11 2 12 2 2 9 2 12 2 2 11 2 12 2 2 11 2 12 2 2 11 2 12 2 2 0 2 12 2 2 11 2 12 2 2
27 9 2 9 2 12 2 2 11 2 12 2 2 11 2 12 2 2 11 2 12 2 2 11 2 12 2 2
3 9 1 11
19 0 9 13 1 0 9 11 2 11 2 1 10 0 9 9 0 9 11 2
30 9 1 9 2 12 2 12 9 2 9 2 4 13 3 1 9 9 2 16 16 4 4 13 14 1 0 9 1 9 2
10 1 0 9 15 3 13 0 9 9 2
24 3 4 1 9 1 0 9 13 1 0 9 0 9 1 9 9 2 15 13 12 9 2 9 2
15 0 9 11 7 13 13 9 9 1 9 0 9 12 9 2
16 16 0 0 9 13 3 3 9 2 1 9 15 13 9 9 2
15 1 9 11 11 2 11 11 7 11 11 2 15 1 11 2
2 0 9
5 11 2 11 2 2
49 9 13 3 9 1 0 9 7 1 9 9 15 7 1 9 13 9 0 9 0 0 9 2 15 13 9 7 0 9 2 13 3 1 11 1 9 0 9 2 9 7 9 9 2 9 2 11 11 2
21 9 15 13 2 16 1 0 9 13 14 0 9 9 9 2 9 7 0 9 9 2
3 9 1 9
6 0 11 2 11 2 2
20 3 12 2 9 0 0 9 9 7 9 0 9 11 13 3 1 0 9 11 2
36 1 9 13 0 9 7 9 12 0 9 1 12 9 9 2 16 0 9 13 3 12 9 1 12 9 2 9 1 12 9 7 9 1 12 9 2
18 3 15 1 9 13 10 0 9 2 3 11 2 11 2 11 7 11 2
6 10 9 13 3 0 2
3 11 11 2
5 1 9 9 1 9
19 0 9 13 9 9 0 1 0 9 11 0 9 2 0 1 9 9 0 9
4 9 13 1 9
5 1 11 13 11 9
4 11 2 11 2
46 0 0 0 9 1 9 1 9 9 1 0 9 1 11 3 13 0 9 9 11 1 0 9 7 13 2 16 13 0 15 13 1 9 9 7 1 9 2 1 15 9 0 9 9 13 2
17 1 0 9 13 0 9 9 0 0 9 1 9 0 9 1 11 2
25 9 11 13 2 16 11 13 12 9 10 0 9 1 9 11 2 7 7 10 0 9 13 9 13 2
20 0 11 13 0 13 16 9 2 3 16 9 2 3 13 3 3 13 0 9 2
26 0 9 1 10 9 13 0 9 1 0 9 7 4 13 0 9 2 16 4 13 0 9 1 0 9 2
8 9 15 4 13 7 9 11 2
13 0 9 4 13 1 9 9 13 1 0 9 9 2
3 0 9 13
5 9 13 1 9 9
2 11 2
35 9 0 9 1 0 9 1 0 9 1 11 11 11 1 9 13 2 16 1 9 1 11 2 13 10 9 2 2 13 7 9 1 9 13 2
34 9 0 9 11 1 0 9 13 2 16 2 15 13 10 0 9 2 15 13 9 2 16 4 13 4 13 0 9 3 1 9 9 2 2
15 3 1 9 15 1 9 13 13 0 9 0 7 0 9 2
19 1 12 9 1 0 12 13 1 9 0 9 0 9 0 9 1 0 9 2
19 1 0 9 13 1 2 9 0 9 2 1 11 1 9 0 9 1 11 2
19 0 9 15 13 3 1 11 1 0 9 2 15 4 13 1 9 0 9 2
3 9 1 11
21 0 9 2 0 9 7 3 0 9 13 1 0 9 9 9 11 11 9 11 11 2
15 2 9 13 2 16 1 0 9 13 13 3 1 0 9 2
8 13 13 7 9 7 9 9 2
14 0 9 13 9 10 0 9 11 2 0 11 1 11 2
27 13 15 2 16 7 1 0 0 9 7 0 9 13 0 1 0 9 3 13 15 9 1 10 0 9 2 2
15 9 9 15 13 0 9 11 2 15 13 9 1 9 9 2
7 9 9 13 1 12 9 2
37 1 9 13 7 0 3 12 9 2 7 3 9 11 2 15 13 0 9 0 9 1 9 2 3 13 2 2 14 13 1 11 3 10 0 9 2 2
17 1 9 2 15 13 1 9 2 13 9 11 13 1 0 9 9 2
3 9 0 9
3 0 0 9
6 0 9 11 2 9 11
6 9 1 15 0 9 2
2 9 9
4 10 9 7 11
5 11 2 11 2 2
11 9 0 9 11 2 11 1 9 3 13 2
29 11 13 1 10 9 2 16 13 9 10 9 10 0 9 1 11 2 11 7 11 1 0 0 9 1 9 10 9 2
19 0 9 13 1 9 9 2 15 13 10 9 9 2 0 9 7 0 9 2
15 0 9 0 0 9 0 0 9 13 0 9 1 10 9 2
11 9 13 3 3 2 1 10 9 3 13 2
31 15 7 13 2 16 0 9 1 0 9 13 0 2 3 11 7 0 9 13 3 1 15 2 0 2 2 16 3 11 11 2
22 3 1 9 9 13 10 0 9 1 0 9 0 9 2 3 15 13 1 9 7 9 2
12 3 13 0 9 1 15 0 2 16 0 9 2
2 0 9
8 9 4 15 13 13 3 3 2
5 13 14 1 9 2
13 12 16 13 1 9 7 1 9 2 13 15 3 2
12 9 3 13 2 7 3 15 1 10 9 13 2
4 15 15 13 2
18 7 10 0 9 13 13 10 9 16 0 9 2 15 15 13 13 9 2
24 13 15 7 0 9 2 0 1 9 1 9 9 1 0 9 1 0 9 1 11 1 11 12 2
36 9 0 9 1 9 4 13 3 13 9 10 9 1 0 9 11 2 3 4 1 12 9 13 14 9 9 7 9 2 7 13 4 7 0 9 2
15 13 4 15 9 9 11 11 2 9 9 0 9 1 11 2
31 13 15 9 9 2 15 4 13 1 9 2 9 15 13 3 13 14 9 2 1 11 3 12 2 9 2 1 15 1 9 2
23 2 1 9 4 13 1 0 9 9 2 1 15 7 3 13 2 7 15 13 1 0 9 2
21 0 0 9 2 0 9 1 11 15 7 13 3 2 7 1 0 9 4 9 13 2
7 7 13 4 13 10 9 2
17 16 13 1 9 7 9 9 2 7 9 2 1 9 1 0 9 2
17 0 9 13 0 9 2 13 3 0 9 7 4 13 9 9 9 2
8 13 15 1 9 1 9 9 2
21 9 2 15 13 1 9 9 2 4 1 9 9 9 13 7 9 13 0 0 9 2
14 1 9 10 0 9 4 13 1 0 9 9 9 2 2
17 0 9 2 15 0 9 0 9 1 9 13 1 9 1 11 12 2
27 0 15 0 2 9 2 9 13 9 9 11 11 11 11 1 0 9 2 15 4 11 13 1 9 0 11 2
4 9 3 1 11
5 11 2 11 2 2
26 15 12 9 11 2 12 0 9 2 15 15 13 0 9 9 11 13 1 11 2 4 13 3 1 11 2
17 13 15 1 0 9 9 0 9 9 2 0 9 7 0 0 9 2
44 2 1 9 9 7 9 0 0 9 13 0 0 9 13 1 0 7 13 9 13 0 9 1 0 9 2 1 10 9 1 11 2 2 13 15 3 0 9 0 0 9 11 11 2
37 16 0 9 0 9 11 11 13 1 15 2 16 1 0 9 13 1 0 2 0 7 0 9 9 2 0 9 9 3 13 2 16 13 1 0 9 2
36 9 12 9 9 4 13 9 13 14 3 2 16 13 1 0 9 0 9 1 9 2 7 7 3 2 16 13 9 1 10 9 1 9 1 9 2
12 0 9 13 3 1 12 2 9 12 9 9 2
37 0 9 1 0 9 11 1 11 11 9 13 3 2 16 13 2 16 0 9 11 2 15 9 13 16 9 2 13 9 3 1 9 3 1 10 9 2
3 9 1 11
22 1 9 9 13 0 9 9 0 9 11 11 2 12 2 7 9 11 11 2 12 2 2
17 12 15 13 13 1 11 11 2 10 9 2 16 1 11 13 9 2
9 11 1 9 12 2 11 1 12 2
17 2 9 4 3 13 13 2 2 13 9 9 11 9 2 11 11 2
22 2 15 1 9 10 0 9 13 2 16 10 9 13 2 7 10 0 9 15 15 13 2
19 12 1 9 13 1 11 1 10 0 9 2 14 1 10 9 3 13 13 2
12 2 13 9 2 16 11 13 9 9 0 9 2
16 2 14 4 1 11 13 1 11 12 9 9 2 2 13 11 2
17 2 15 13 9 2 16 9 13 13 2 3 3 13 1 10 9 2
10 3 2 11 15 13 1 12 12 9 2
14 9 13 2 3 15 13 0 9 2 7 15 15 13 2
14 13 3 2 16 16 10 9 13 1 11 2 13 15 2
18 3 7 13 2 16 1 9 1 11 13 7 1 10 9 15 15 13 2
24 3 13 1 11 7 13 13 1 11 2 3 15 9 0 9 9 2 9 13 9 9 7 9 2
8 1 0 9 4 9 13 2 2
4 9 1 0 9
10 11 7 0 12 9 1 0 9 13 9
21 3 1 9 15 10 0 9 3 13 9 2 3 3 1 9 1 11 13 11 2 2
18 1 9 9 1 0 9 1 9 1 9 12 13 14 1 0 9 9 2
20 3 3 13 11 7 12 9 1 9 2 1 9 1 0 9 2 13 0 9 2
19 9 13 10 9 1 12 9 1 0 9 2 11 1 9 13 11 1 11 2
7 9 13 1 9 0 9 2
20 11 3 13 7 1 12 2 3 13 0 11 2 7 10 9 10 0 9 13 2
13 1 9 9 7 1 0 9 1 9 7 3 3 2
18 3 1 12 2 9 2 13 11 1 2 15 1 9 3 13 9 11 2
20 1 12 2 9 2 13 0 9 11 2 3 13 11 7 15 3 13 9 11 2
20 1 9 3 15 3 1 9 11 13 0 0 9 1 9 11 2 12 2 12 2
11 3 3 15 13 0 9 1 9 9 13 2
35 9 1 0 9 11 13 1 0 9 2 3 0 3 13 11 2 15 15 9 2 13 2 1 9 14 1 11 2 7 13 15 3 1 15 2
5 3 3 0 9 2
7 9 13 9 2 9 9 2
25 1 10 9 9 13 3 9 1 0 9 7 13 15 1 9 3 2 1 9 9 0 9 7 9 2
21 13 14 1 9 2 16 0 9 13 3 0 2 16 9 13 15 3 1 15 13 2
15 1 3 0 9 15 15 0 9 3 13 13 7 1 9 2
13 9 3 13 2 7 0 9 1 0 9 9 13 2
18 1 9 13 3 9 11 1 12 2 9 2 7 9 11 10 9 13 2
10 1 9 13 9 11 13 0 7 13 2
14 11 2 15 3 13 1 9 1 11 2 13 10 9 2
16 3 15 13 9 7 11 2 15 13 12 9 1 9 9 9 2
15 9 9 13 0 0 9 1 9 0 1 9 11 2 11 2
10 0 9 10 9 13 0 7 0 11 2
10 14 2 14 3 13 9 1 10 9 2
3 9 12 2
7 11 2 12 2 7 12 2
4 11 2 12 2
6 0 2 1 9 2 2
6 9 11 2 11 2 2
3 9 12 2
5 15 11 1 11 13
7 9 1 0 11 13 0 9
11 2 13 15 3 0 2 3 4 15 13 2
5 13 4 0 9 2
31 1 12 9 3 1 9 7 3 3 13 1 9 2 2 2 2 2 13 9 3 3 1 0 11 0 9 11 11 11 11 2
30 9 9 12 3 1 11 2 9 7 9 3 2 0 1 11 2 2 7 1 15 0 9 1 9 7 1 9 1 9 2
29 9 11 2 3 13 0 9 11 2 11 2 9 7 11 2 1 9 0 9 11 9 2 13 0 9 1 0 9 2
16 10 0 9 13 12 9 1 12 2 9 15 15 13 12 9 2
11 3 1 11 15 13 1 0 0 9 11 2
29 0 9 13 0 9 7 9 0 9 15 0 9 13 13 9 2 16 3 3 13 9 2 0 1 9 3 1 9 2
8 13 15 13 0 9 2 2 2
24 7 2 9 11 12 2 12 15 13 1 12 2 12 2 0 11 3 13 2 7 9 3 13 2
18 9 15 13 1 12 2 16 15 13 0 9 2 1 15 9 9 13 2
20 11 11 14 3 13 1 9 2 2 9 9 2 1 9 15 15 15 13 2 2
12 0 13 2 16 3 15 13 13 1 11 9 2
9 16 15 13 2 13 11 3 13 2
5 15 1 11 13 2
6 0 9 13 1 9 11
24 9 9 1 0 9 0 9 1 9 9 11 3 13 9 11 0 9 2 0 2 11 7 11 2
8 9 13 12 9 0 9 11 2
47 13 1 0 9 11 2 1 9 11 7 11 2 1 9 9 0 1 9 0 9 11 7 0 9 11 7 0 9 11 7 1 9 0 9 7 0 9 1 11 3 3 0 9 11 7 11 2
17 1 9 1 0 9 9 4 13 0 9 0 0 7 0 9 9 2
3 9 1 11
6 0 11 2 11 2 2
21 1 12 2 9 4 13 4 13 0 9 1 9 0 0 9 1 0 9 0 9 2
24 1 0 11 7 11 2 3 9 1 0 9 3 9 13 2 1 9 13 3 12 0 0 9 2
18 3 4 15 13 13 0 10 0 9 2 16 0 9 13 1 12 9 2
24 9 1 9 2 0 9 7 9 4 13 12 9 9 7 0 9 4 13 4 13 1 9 12 2
8 9 0 9 13 1 0 9 0
36 11 7 11 13 1 9 1 11 1 9 2 9 2 0 9 2 7 1 9 13 9 1 15 2 16 15 11 13 3 2 3 7 13 15 9 2
20 9 15 3 13 1 0 2 16 13 0 9 13 2 16 4 15 13 10 9 2
10 0 9 15 9 13 1 0 9 0 2
23 1 9 12 15 13 9 10 9 2 16 15 9 13 1 0 9 2 15 13 7 9 9 2
28 3 2 16 9 13 9 13 9 9 10 0 9 2 13 3 0 9 2 16 13 9 2 15 13 1 9 0 2
5 11 1 9 1 11
23 15 3 13 0 9 2 15 13 2 16 3 11 7 10 9 13 9 9 1 11 7 11 2
15 0 9 13 11 11 2 16 4 10 9 1 9 13 9 2
29 9 1 9 11 13 1 9 9 1 0 9 0 9 9 11 11 9 0 9 9 2 15 15 1 9 13 16 9 2
29 11 13 2 16 9 13 1 9 15 9 0 0 11 2 16 0 9 13 1 9 1 11 3 1 9 0 11 13 2
9 11 13 2 16 9 13 13 9 2
17 9 1 9 0 9 1 0 9 13 9 11 2 11 7 0 9 2
18 13 2 16 9 7 9 9 9 1 10 9 13 1 9 1 9 11 2
20 9 13 1 9 1 11 2 11 7 11 2 11 2 11 2 11 7 0 9 2
17 0 9 13 0 9 2 16 9 13 15 0 0 9 1 0 9 2
33 0 9 3 13 1 9 2 7 13 9 2 16 9 13 1 9 1 9 2 16 15 13 1 12 9 0 9 0 0 9 11 11 2
29 1 15 1 9 2 16 1 9 9 13 10 3 0 9 2 15 4 13 4 3 13 1 9 2 0 9 13 13 2
50 9 9 2 3 13 3 11 7 11 2 7 1 9 13 9 1 9 2 16 11 13 0 9 0 9 1 9 12 0 0 9 2 15 15 3 13 1 9 9 1 9 2 1 15 11 13 14 12 9 2
21 11 2 1 11 15 13 1 9 2 9 0 9 2 11 1 10 9 1 0 9 2
36 1 9 9 0 1 9 9 4 0 11 2 15 15 13 3 1 11 7 0 9 2 13 1 9 2 15 15 13 1 11 13 9 1 0 9 2
31 9 0 9 4 11 4 3 13 1 9 2 16 4 13 3 13 0 9 2 13 0 9 1 10 0 9 7 13 10 9 2
5 11 13 13 0 9
2 11 2
2 11 2
5 11 13 13 0 9
2 11 2
11 11 13 1 11 7 11 13 12 0 9 2
37 13 15 3 1 0 9 1 11 0 9 7 9 0 9 1 0 9 11 11 2 15 15 1 0 9 13 0 9 0 9 1 0 9 2 11 2 2
18 1 10 9 7 1 9 3 4 13 10 9 7 15 13 1 9 9 2
11 0 9 13 0 9 0 9 0 9 9 2
3 10 9 9
28 0 9 9 11 11 3 13 2 16 16 4 2 9 2 13 9 11 2 3 13 13 7 0 9 1 0 9 2
13 0 9 15 13 2 16 3 12 9 3 15 13 2
19 9 0 9 11 11 3 13 2 16 11 11 13 9 1 9 9 1 11 2
17 9 13 3 3 0 7 13 15 2 16 9 1 12 9 13 0 2
22 12 9 13 15 0 2 0 9 15 1 9 13 3 1 9 2 1 15 13 9 9 2
35 16 15 15 0 13 0 9 1 9 9 2 13 15 3 3 13 2 0 9 13 9 9 0 9 7 9 15 13 13 2 16 15 9 13 2
26 16 15 7 1 9 13 0 9 7 13 15 2 15 13 1 9 7 9 1 9 2 13 15 1 9 2
9 1 9 11 11 7 14 1 9 2
27 9 1 11 7 0 9 13 0 15 1 15 7 9 0 9 9 0 1 9 9 0 9 13 0 7 0 2
26 13 3 9 1 9 3 0 7 13 7 9 0 9 1 9 2 15 13 3 0 2 13 14 0 9 2
17 9 9 7 0 9 0 9 11 11 13 3 0 2 7 3 0 2
23 9 9 13 1 9 0 9 7 0 9 7 0 9 0 9 1 9 15 1 15 14 13 2
39 3 1 0 9 9 9 15 3 1 9 13 0 9 2 0 0 9 13 9 0 7 0 9 2 15 3 13 1 9 10 0 9 3 0 9 0 0 9 2
14 9 13 1 9 10 9 13 7 13 15 14 1 9 2
7 1 15 13 9 3 0 2
19 0 9 13 9 7 13 9 2 3 16 15 13 13 15 0 16 0 9 2
9 0 9 4 15 15 13 3 13 2
26 1 9 9 9 9 1 9 13 9 9 9 0 15 0 9 0 9 2 15 4 13 0 9 7 9 2
21 9 9 11 11 3 13 2 16 9 13 13 1 10 9 2 0 9 1 9 2 2
2 9 13
10 11 11 2 9 0 9 9 1 9 2
22 10 9 1 0 12 1 11 12 2 15 4 13 1 9 2 15 13 1 0 10 9 2
18 13 3 7 13 1 9 9 7 9 3 9 9 0 0 7 0 9 2
20 13 3 9 9 1 0 9 1 11 7 9 7 9 3 0 9 1 9 9 2
31 0 4 13 2 16 9 0 9 2 7 16 15 15 10 9 13 2 7 3 13 13 15 2 13 3 0 16 9 3 0 2
24 3 13 3 3 0 2 7 10 9 15 3 13 13 3 14 9 7 10 0 9 13 3 0 2
17 13 13 9 2 15 0 9 3 13 7 13 15 13 15 1 9 2
4 9 9 3 0
6 0 11 2 11 2 2
24 7 0 9 9 0 9 1 0 0 9 1 9 0 9 0 11 7 11 13 1 10 9 9 2
11 9 13 1 10 0 9 2 9 13 9 2
26 9 13 1 15 9 1 0 9 11 2 3 9 3 1 9 13 1 9 0 9 2 15 15 13 9 2
23 9 9 3 0 0 9 3 3 13 1 12 9 9 1 15 2 16 1 15 13 0 9 2
32 0 9 2 16 0 9 13 0 9 2 15 13 9 2 7 16 9 7 9 9 15 9 13 2 4 1 10 9 3 13 9 2
25 9 9 15 13 2 16 9 0 12 9 2 1 15 13 3 13 0 9 2 15 0 9 4 13 2
25 13 7 9 10 9 13 7 13 15 9 1 3 0 0 9 0 0 9 2 15 4 13 9 9 2
27 2 9 9 13 12 1 0 9 2 15 4 13 1 9 0 0 9 2 2 13 0 9 10 9 1 9 2
20 15 9 1 9 7 9 1 10 9 13 1 9 1 9 0 9 7 10 9 2
19 15 4 13 3 13 2 16 0 9 1 0 11 15 4 1 9 3 13 2
2 9 13
9 1 0 9 9 9 13 1 9 2
22 9 9 9 11 15 13 13 1 0 9 11 7 11 2 15 1 9 9 13 1 11 2
11 1 0 9 15 13 3 7 11 1 11 2
25 11 1 0 12 9 13 1 11 11 2 12 9 0 9 2 7 12 9 0 9 11 1 11 11 2
23 0 9 11 11 4 13 11 2 13 1 11 2 7 11 11 7 11 2 0 13 3 11 2
15 11 11 11 15 13 1 0 9 11 7 0 0 9 11 2
10 0 9 4 13 1 9 9 0 11 2
21 1 11 11 7 11 3 13 7 11 1 11 7 11 2 11 11 7 11 1 11 2
10 0 13 3 0 9 11 7 11 11 2
18 3 1 9 13 0 0 9 11 11 7 0 11 11 2 3 11 2 2
16 1 0 11 13 0 9 12 0 9 9 12 2 12 11 11 2
2 1 9
40 0 9 1 12 2 9 0 0 9 2 11 13 1 11 2 12 2 9 2 12 2 12 7 13 13 2 13 15 9 0 1 9 0 9 2 11 2 11 0 2
7 0 9 0 9 13 11 2
9 13 1 9 11 11 12 2 12 2
6 9 11 13 11 11 2
14 11 2 11 7 11 13 1 0 9 1 9 9 12 2
21 9 11 13 11 0 2 11 9 12 9 1 0 9 9 9 1 9 1 11 11 2
18 1 9 13 11 1 11 2 12 12 9 2 2 2 1 9 14 11 2
3 13 11 2
3 3 1 9
24 0 9 15 3 13 0 0 9 7 13 9 2 13 11 0 0 9 7 1 9 1 0 11 2
16 9 13 3 9 11 1 11 2 15 3 14 13 1 0 9 2
6 9 2 7 9 9 2
5 11 2 11 2 2
31 9 11 3 13 9 11 11 2 11 2 2 16 4 4 0 9 9 1 0 9 2 0 9 2 13 1 9 0 9 9 2
42 16 1 15 13 9 0 7 0 9 2 9 9 11 2 10 9 11 7 0 0 9 0 0 9 2 7 13 1 10 9 9 9 2 13 15 0 9 7 0 9 11 2
24 9 12 9 13 1 9 0 9 2 15 13 9 9 13 9 9 2 16 1 15 0 9 13 2
15 14 9 11 11 2 11 2 15 13 1 9 13 9 9 2
30 3 2 10 9 2 3 1 11 7 11 2 0 9 13 16 9 9 2 15 9 13 2 1 9 1 9 9 7 9 2
37 9 9 11 11 2 11 2 15 3 1 10 0 9 13 2 2 13 15 2 16 0 9 2 15 9 3 1 9 13 2 4 10 0 9 13 13 2
34 7 1 9 2 3 9 13 12 9 1 9 7 10 9 13 3 3 13 2 3 2 16 15 13 3 1 9 2 13 4 13 9 9 2
9 0 9 13 3 1 15 1 9 2
34 15 15 15 3 13 2 16 1 9 2 15 4 13 2 4 13 9 7 13 1 9 2 15 13 3 0 9 9 2 16 13 0 2 2
5 9 13 3 0 9
13 3 0 9 3 13 9 9 9 1 11 1 11 2
15 9 13 1 9 3 7 3 15 13 14 1 9 12 9 2
34 3 15 13 9 9 0 9 9 0 9 1 11 1 11 9 2 11 11 2 1 9 15 1 15 13 9 2 15 13 1 9 12 9 2
7 13 0 7 0 9 9 2
10 9 15 13 1 0 0 9 0 9 2
13 9 3 13 13 2 14 9 1 9 13 1 9 2
47 1 9 9 15 0 12 9 13 14 12 9 2 1 0 9 9 0 9 1 11 1 11 2 9 2 0 9 0 9 2 11 7 9 1 11 7 10 0 0 9 1 0 9 1 0 11 2
24 1 0 9 1 9 4 13 7 9 2 15 1 9 13 12 9 9 2 7 13 9 15 13 2
7 3 15 9 13 14 9 2
16 0 9 3 1 9 0 9 3 13 2 16 1 9 13 9 2
10 9 0 9 9 11 13 9 0 9 2
1 9
2 11 12
6 12 9 2 9 2 9
4 12 9 2 9
3 12 9 9
2 12 9
12 12 1 9 1 9 2 11 11 2 11 11 2
2 12 9
2 12 9
3 12 9 9
5 9 1 12 1 12
3 12 9 9
5 12 9 9 11 12
2 12 11
4 12 9 2 12
3 12 9 9
2 12 11
7 12 11 13 2 13 2 13
3 12 0 9
5 12 14 11 2 12
4 12 9 2 9
6 12 11 2 12 2 2
2 12 9
2 12 9
3 12 9 9
4 12 13 9 9
7 12 9 0 2 12 2 2
5 9 1 12 1 12
3 12 9 11
2 12 9
3 12 9 12
4 12 9 0 9
7 12 9 0 2 12 2 2
7 12 9 1 11 2 11 11
3 12 0 9
5 12 9 1 9 11
3 12 0 9
6 12 11 11 5 11 11
3 12 0 9
3 12 9 9
4 12 11 0 11
6 12 9 2 12 2 2
4 12 9 1 9
3 12 9 11
4 12 11 2 11
5 12 11 2 0 9
2 12 11
5 12 9 9 2 12
3 12 9 11
7 12 9 1 9 7 1 9
6 12 13 2 2 2 2
2 13 2
4 12 9 2 12
4 12 11 1 11
4 12 13 9 9
2 12 9
3 12 9 11
4 12 0 9 11
12 1 9 11 15 1 9 3 13 13 0 9 11
2 11 2
19 13 4 3 2 16 4 13 2 13 1 10 9 1 11 0 9 11 11 2
21 1 2 0 9 2 3 13 10 9 1 9 0 9 12 0 0 9 9 9 11 2
16 13 2 16 0 9 1 9 11 11 3 3 13 10 0 9 2
30 9 15 1 9 1 9 13 0 9 11 11 2 16 13 2 16 13 0 7 0 2 15 15 15 1 15 1 9 13 2
12 3 15 13 7 1 0 9 1 11 11 11 2
10 13 2 7 13 11 9 9 0 9 2
6 10 9 3 1 0 11
3 0 11 2
27 0 9 1 0 9 3 3 13 1 9 9 0 9 2 15 15 1 9 13 13 11 9 13 1 0 9 2
11 1 10 9 13 3 3 1 11 0 9 2
54 1 0 0 9 2 1 15 13 9 15 1 9 7 3 3 13 7 3 3 0 9 13 9 15 9 1 11 1 9 9 2 3 1 9 13 9 2 16 11 13 7 3 9 11 7 16 9 0 9 13 3 3 12 2
10 13 15 15 3 0 0 9 1 11 2
8 11 7 9 13 0 9 1 9
2 11 2
30 9 11 2 11 11 11 7 0 7 0 9 3 13 9 9 7 9 11 11 11 0 15 0 9 2 0 1 0 9 2
36 1 9 9 11 3 2 13 2 2 0 9 13 13 9 2 15 13 3 0 10 9 7 0 0 9 1 11 13 10 0 9 1 0 9 2 2
24 11 13 2 16 13 9 2 3 15 13 9 16 12 1 9 3 0 0 9 7 3 15 13 2
27 2 3 3 13 9 2 3 15 3 13 0 13 2 3 3 13 0 13 9 15 3 0 2 2 13 9 2
9 0 9 13 11 1 0 7 0 2
14 13 2 16 0 9 13 13 3 16 16 9 0 9 2
23 2 9 16 2 0 9 2 7 2 13 0 13 9 15 3 0 2 2 15 13 9 9 2
24 9 13 0 9 7 13 9 1 9 7 0 2 15 3 3 1 9 15 13 2 2 13 11 2
33 2 9 2 16 4 15 13 9 7 4 13 1 15 2 16 15 7 15 13 0 9 10 9 2 13 1 15 3 0 2 2 13 2
10 0 7 0 9 13 1 0 9 9 2
34 2 10 9 1 10 9 4 13 10 9 2 7 3 3 9 10 9 0 9 2 2 13 9 1 9 0 9 0 7 9 0 11 11 2
20 2 13 15 15 0 1 9 0 9 13 13 2 15 9 13 2 7 13 13 2
17 13 7 9 1 15 2 16 15 16 9 13 3 2 2 13 9 2
12 13 2 16 13 0 13 1 9 9 1 9 2
11 1 9 9 9 13 3 9 11 11 11 2
10 3 13 13 0 9 16 0 9 9 2
14 0 11 11 13 10 9 1 9 2 15 13 9 13 9
5 9 9 1 9 12
5 11 2 11 2 2
20 9 2 9 7 9 9 0 9 13 1 0 9 3 13 1 12 2 9 12 2
17 3 1 9 0 9 13 13 9 9 2 1 15 13 10 9 13 2
18 9 9 2 0 9 2 13 13 9 9 9 9 2 15 3 13 9 2
19 0 1 9 0 0 9 2 0 2 9 2 13 13 1 12 2 9 12 2
21 9 0 9 4 1 9 13 4 3 13 9 2 9 13 9 0 0 9 9 2 2
16 9 7 9 13 3 0 13 1 0 9 9 0 9 12 9 2
10 9 1 9 9 13 12 7 12 9 2
13 9 9 11 11 13 9 1 9 9 1 10 9 2
23 13 2 16 1 9 9 13 1 9 1 12 12 0 9 1 9 1 12 7 12 9 9 2
9 1 9 13 12 9 1 0 9 2
8 1 9 13 11 13 0 9 2
5 0 9 13 1 9
7 11 2 11 2 11 2 2
21 9 14 10 10 9 15 1 0 9 0 2 9 13 1 9 1 0 9 0 9 2
13 10 9 13 9 9 16 0 9 1 9 7 9 2
33 13 15 2 16 3 1 9 11 13 9 0 2 9 0 13 1 9 3 1 9 12 7 12 9 1 9 1 0 9 12 9 9 2
14 13 15 9 1 12 9 10 9 1 9 12 12 9 2
19 15 13 2 16 0 0 9 9 9 13 12 9 2 3 0 9 0 9 2
41 3 1 9 9 11 0 11 2 15 13 0 9 12 7 12 12 9 2 7 13 15 3 0 9 1 9 0 9 2 4 13 0 9 2 7 15 1 0 9 9 2
23 9 0 9 15 13 1 0 9 0 9 2 15 13 9 2 16 13 1 0 9 3 0 2
37 1 0 9 4 13 9 9 12 9 9 1 9 12 9 2 1 0 9 12 9 9 1 9 9 12 9 7 1 0 9 12 12 9 1 0 9 2
28 9 0 9 4 13 1 12 9 9 1 9 12 9 2 15 13 9 1 12 9 0 2 16 13 9 0 9 2
20 3 3 1 9 9 0 9 15 13 1 0 9 0 9 2 3 1 12 9 2
13 3 13 9 12 9 1 0 9 1 12 12 9 2
33 9 11 4 3 13 1 0 9 2 10 9 15 3 3 13 1 9 0 9 7 13 3 0 9 9 9 1 0 9 0 2 9 2
33 16 15 13 2 1 0 9 0 9 4 13 3 9 0 9 11 2 12 9 2 2 15 15 1 9 9 13 0 9 13 3 0 2
25 3 9 9 7 9 11 1 11 2 12 9 2 7 11 11 2 12 9 2 13 0 9 0 9 2
17 12 9 1 9 0 9 15 13 1 9 11 11 2 12 9 2 2
7 9 9 13 12 9 9 2
23 13 15 3 9 2 16 1 9 10 9 13 3 0 9 2 16 4 1 0 9 3 13 2
29 9 0 9 11 2 15 4 13 1 3 0 2 4 13 1 0 9 0 9 2 12 9 2 1 9 12 12 9 2
22 1 12 9 9 15 13 9 0 9 2 11 7 15 3 1 0 0 9 2 12 9 2
22 3 15 13 1 9 9 11 2 15 13 3 9 1 9 7 1 0 9 15 13 9 2
15 13 15 15 1 12 9 1 9 12 9 2 0 9 2 2
13 9 0 9 7 0 0 9 9 13 1 0 9 2
4 9 9 3 13
2 11 2
17 12 1 0 9 9 13 1 9 9 1 0 9 3 9 0 9 2
19 1 0 1 15 13 9 2 9 2 2 15 9 13 1 9 0 9 9 2
28 9 2 15 15 9 13 1 0 0 9 2 15 13 1 9 9 9 3 13 1 0 9 0 1 3 0 9 2
9 9 1 9 13 1 9 12 9 2
21 9 4 13 13 0 9 9 2 1 15 13 13 2 16 9 9 13 3 0 9 2
31 1 0 9 13 3 0 9 3 9 0 2 0 2 0 2 9 2 1 15 13 13 2 16 9 9 13 1 15 3 0 2
16 1 12 2 9 13 13 0 9 1 10 9 9 0 9 11 2
14 10 0 9 13 12 12 9 7 0 0 9 12 9 2
20 9 9 2 16 13 1 0 9 2 13 12 9 2 1 12 2 9 12 2 2
28 9 15 13 9 1 0 9 13 1 0 12 2 9 2 3 13 0 9 13 3 1 9 3 0 1 0 9 2
16 3 0 9 13 12 2 9 9 3 0 9 1 0 9 9 2
9 10 0 9 13 3 12 12 9 2
24 0 9 13 1 0 9 13 0 9 12 9 7 1 0 9 3 2 1 9 0 9 7 9 2
7 0 9 15 3 13 13 2
26 9 1 0 9 3 13 2 3 16 1 0 9 15 9 13 9 13 1 15 9 0 9 1 0 9 2
10 9 15 1 10 9 13 3 1 9 2
27 9 1 0 9 12 2 12 2 12 7 12 12 9 0 12 2 9 12 13 1 9 12 3 9 11 11 2
16 13 0 9 12 9 7 0 9 14 12 9 1 0 0 9 2
7 9 9 15 13 12 3 2
11 15 0 9 13 0 1 9 0 9 11 2
14 1 9 13 9 9 1 9 1 9 0 9 0 9 2
3 0 0 9
2 11 2
32 12 0 9 7 9 2 11 11 11 2 11 11 11 2 11 11 11 2 11 2 11 11 11 2 11 11 11 7 11 11 11 2
25 9 2 12 0 9 2 9 0 1 9 7 1 9 9 11 11 2 3 13 0 0 9 0 9 2
36 0 9 13 1 9 9 1 0 11 11 2 1 9 15 13 1 9 0 11 7 0 9 0 9 9 15 13 1 9 1 9 0 9 1 11 2
25 13 15 4 0 9 14 1 9 9 2 1 9 13 1 0 9 2 15 13 9 1 9 1 11 2
33 0 9 1 0 9 13 11 1 12 9 2 16 13 9 1 11 11 2 2 13 4 1 12 9 7 13 1 15 9 1 0 9 2
20 0 9 13 7 3 0 2 13 4 15 9 2 16 10 9 4 13 0 9 2
12 3 13 1 9 0 9 7 9 12 9 2 2
14 9 2 16 13 2 14 2 9 2 9 9 3 13 2
23 9 13 9 12 0 9 2 9 9 13 14 9 1 9 2 15 13 12 2 0 9 2 2
30 9 9 2 9 11 11 2 15 13 9 9 2 9 2 1 15 13 9 1 10 9 0 16 1 0 2 0 2 9 2
11 3 3 13 7 9 2 3 3 7 3 2
33 10 9 7 3 13 1 0 9 2 3 16 15 9 13 9 9 9 2 11 1 9 2 16 4 1 15 13 1 0 9 2 2 2
30 1 9 9 15 1 11 11 1 0 11 1 11 11 13 0 11 2 7 3 0 9 0 9 1 9 9 1 11 11 2
32 2 13 13 0 9 1 0 9 2 1 0 9 7 9 2 1 15 15 13 1 0 9 9 2 2 13 1 9 9 11 11 2
6 2 13 15 16 9 2
9 13 9 2 15 4 15 13 13 2
17 9 9 15 3 13 9 2 16 4 1 15 13 2 15 13 2 2
5 0 9 9 7 11
23 0 9 2 16 0 0 9 13 1 0 9 9 7 9 1 10 9 15 13 2 15 13 2
13 11 11 3 13 14 9 9 2 7 7 10 9 2
28 9 9 11 11 11 1 9 1 11 0 7 4 13 12 1 9 9 2 3 9 9 0 9 1 10 0 9 2
21 2 13 15 13 9 9 2 16 3 13 10 9 2 2 13 3 1 9 11 11 2
20 0 9 2 1 15 4 15 9 13 0 13 2 15 7 1 15 9 13 13 2
8 13 3 9 11 11 0 9 2
9 3 9 1 9 13 2 16 13 2
31 1 0 9 9 13 9 14 11 7 11 7 1 9 1 0 7 11 2 11 2 7 3 0 9 11 2 11 7 0 9 2
20 9 2 3 9 9 13 9 1 9 0 9 2 13 3 2 12 13 3 0 2
17 3 13 15 3 9 2 15 13 9 2 16 4 9 1 9 13 2
14 15 13 1 9 2 16 4 13 7 9 2 7 9 2
27 0 9 13 9 11 11 2 15 15 3 1 0 9 13 0 9 7 9 9 14 0 9 2 7 7 9 2
11 13 0 0 9 9 11 1 0 0 9 2
24 13 0 2 16 0 9 3 13 0 9 1 0 9 2 7 3 3 10 9 13 0 9 9 2
29 7 11 13 0 9 0 9 9 7 1 10 9 2 16 15 9 13 2 4 15 13 2 16 4 0 9 9 13 2
32 12 9 4 13 9 1 9 2 16 9 1 11 2 3 14 9 9 2 4 13 15 2 10 9 15 2 10 2 9 13 13 2
4 9 13 9 11
5 11 2 11 2 2
14 0 9 1 0 9 7 11 4 13 13 9 9 11 2
17 10 9 0 0 9 1 9 0 11 7 0 11 1 10 9 13 2
14 3 15 1 15 1 11 13 0 0 2 0 0 9 2
24 1 9 9 13 7 12 9 1 10 9 2 16 9 1 9 13 13 1 9 9 9 1 9 2
10 0 9 4 13 4 13 1 9 12 2
3 9 1 9
5 1 9 1 11 2
17 1 9 12 9 1 12 1 12 1 9 11 1 11 2 0 9 2
5 9 1 9 11 2
18 9 2 3 1 11 2 12 9 1 11 2 9 2 12 7 12 9 2
4 9 9 9 2
15 12 2 12 2 12 9 1 9 1 11 12 7 12 9 2
6 0 9 13 9 1 9
10 9 11 2 13 1 9 16 1 9 2
5 11 2 11 2 2
23 0 9 0 9 4 13 13 1 10 0 9 1 9 12 9 9 7 0 12 9 10 9 2
18 13 15 3 0 9 0 9 1 9 2 15 15 13 1 15 0 9 2
32 13 1 15 2 16 1 9 0 9 11 4 9 13 9 13 15 0 9 2 15 15 3 4 3 13 14 1 9 10 0 9 2
14 0 9 7 10 0 9 13 13 2 13 15 1 9 2
32 9 1 10 9 13 3 9 11 11 2 1 0 9 7 9 9 9 2 0 10 9 11 11 2 13 9 2 9 2 14 9 2
26 2 13 1 9 16 1 9 2 7 14 16 1 9 2 2 13 1 10 9 9 9 0 9 11 11 2
25 2 14 2 16 3 13 9 2 3 0 9 13 1 0 9 9 2 15 0 9 9 3 13 2 2
23 9 11 13 2 16 10 9 13 13 3 9 1 9 7 9 2 7 10 10 9 4 13 2
20 11 11 2 9 0 9 11 11 2 13 2 16 10 9 3 10 9 9 13 2
14 2 16 9 15 13 2 14 13 9 9 2 2 13 2
16 2 10 9 13 1 0 9 2 2 13 0 9 9 11 11 2
18 2 0 9 13 1 9 0 9 2 7 9 0 9 13 15 1 9 2
8 13 15 9 1 0 9 2 2
39 9 3 3 13 1 0 9 9 7 13 15 3 1 10 9 9 2 1 15 15 13 1 15 2 16 2 9 13 0 9 0 7 3 0 9 0 9 2 2
28 2 14 16 4 3 15 1 9 0 9 9 13 1 10 3 0 9 1 10 9 2 2 13 0 9 9 11 2
27 1 9 15 13 7 1 15 2 16 9 1 0 9 13 10 9 7 16 2 14 3 15 10 9 13 2 2
19 2 15 13 0 9 2 2 13 9 11 2 2 1 10 9 9 3 13 2
12 0 9 1 10 9 13 3 1 3 0 2 2
7 9 0 9 13 0 0 9
26 9 9 9 9 11 11 1 10 9 2 16 13 13 0 9 9 11 2 13 2 16 10 9 9 13 2
15 0 9 4 9 13 1 0 9 7 15 15 13 10 9 2
21 9 15 13 3 1 9 9 9 2 9 9 15 1 9 9 3 0 9 13 9 2
38 9 11 2 15 3 13 1 11 2 15 1 0 9 10 0 9 13 2 13 7 2 16 3 13 1 10 9 1 9 9 11 9 1 9 12 2 9 2
12 0 9 14 3 13 13 2 13 13 0 9 2
5 2 13 0 9 2
25 3 1 15 13 9 9 2 7 13 4 15 3 2 16 13 0 9 2 16 4 13 0 9 3 2
5 3 4 15 13 2
34 0 4 1 12 9 9 1 0 9 7 1 11 9 13 1 10 9 2 7 4 15 9 0 9 13 1 9 2 2 13 11 2 11 2
10 0 0 9 4 15 13 13 9 9 2
15 9 0 9 1 0 13 11 11 2 11 11 7 11 11 2
3 13 0 9
5 11 2 11 2 2
24 1 9 12 4 13 13 1 0 9 9 9 1 11 1 0 12 9 1 12 7 12 9 3 2
10 13 15 3 9 9 0 9 11 11 2
26 16 3 13 2 9 0 9 0 0 9 3 13 1 0 9 9 10 9 2 7 3 13 10 0 9 2
27 10 9 4 13 13 1 10 9 2 16 9 4 15 13 3 0 2 3 2 1 9 9 9 1 0 9 2
25 9 9 7 9 13 1 10 9 1 9 13 9 9 2 15 13 1 9 9 13 2 1 9 9 2
5 11 4 14 13 9
5 11 2 11 2 2
12 0 9 15 7 1 9 13 13 0 0 9 2
11 9 9 7 13 9 0 9 1 9 9 2
16 9 3 13 1 9 9 2 3 9 0 9 13 0 0 9 2
24 1 0 9 9 11 11 4 0 9 1 12 9 13 3 12 9 9 2 3 3 4 13 9 2
7 0 9 9 9 1 9 9
5 11 2 11 2 2
32 1 11 1 0 9 11 13 3 0 1 12 9 2 1 15 15 13 2 16 15 13 9 9 1 9 2 1 15 13 9 9 2
17 9 11 11 2 12 2 13 9 3 2 16 13 12 0 11 11 2
11 0 9 13 1 9 12 12 0 11 11 2
31 9 11 11 1 0 11 1 11 13 1 9 12 2 16 13 13 9 9 2 7 1 9 3 15 1 15 13 9 9 9 2
15 3 7 13 1 0 9 3 14 1 10 9 1 9 12 2
5 1 9 11 13 9
2 11 2
30 0 9 13 1 9 1 0 9 1 0 0 9 11 2 15 9 9 11 13 1 12 1 12 0 2 2 0 9 2 2
7 13 1 15 3 0 9 2
28 0 9 2 15 13 0 11 0 9 0 9 2 3 4 13 7 1 9 11 13 1 0 0 9 0 9 13 2
16 0 0 2 0 9 2 11 13 1 0 9 1 9 9 9 2
18 0 9 11 3 13 2 16 0 0 9 13 1 11 1 0 9 9 2
21 1 0 0 9 0 7 0 9 1 0 11 7 3 11 3 1 11 13 0 9 2
28 0 0 9 11 13 3 3 0 9 2 15 1 0 9 13 3 10 9 7 0 9 1 0 9 1 9 9 2
29 12 0 2 12 0 7 12 0 9 13 1 9 1 9 1 0 11 12 9 9 0 9 1 9 1 9 9 11 2
16 15 12 9 15 1 9 1 9 13 1 9 1 11 1 11 2
22 1 9 4 3 13 9 0 0 9 1 0 11 1 11 2 15 4 13 12 2 9 2
16 1 0 0 0 9 13 12 9 9 2 12 11 12 9 9 2
1 11
4 15 13 10 9
1 11
26 12 9 1 11 4 13 13 9 10 9 2 15 15 3 13 1 9 9 2 1 0 2 9 2 2 2
29 13 3 2 16 13 7 9 9 7 16 1 9 9 2 7 9 2 4 13 9 11 2 9 2 2 11 7 11 2
24 3 4 13 9 10 9 3 13 2 7 3 15 13 1 9 2 15 4 13 1 0 0 9 2
27 13 0 2 16 15 9 11 13 1 9 9 2 7 1 9 2 9 2 1 15 15 13 9 2 9 2 2
15 13 2 14 9 9 2 13 15 3 1 9 0 9 11 2
35 9 2 1 0 9 15 9 13 3 3 16 1 9 0 2 9 15 13 1 9 0 2 2 7 1 0 9 13 3 1 9 1 9 0 2
5 3 13 9 11 2
17 9 0 0 9 11 2 15 13 0 9 0 9 11 2 7 2 2
22 9 13 10 9 1 9 2 7 15 15 15 13 1 9 2 11 2 3 2 11 2 2
28 1 9 2 11 2 11 13 0 9 2 15 15 13 1 0 9 16 9 0 2 3 2 10 9 13 9 2 2
26 9 12 2 15 13 0 9 9 2 13 3 2 12 2 2 7 1 0 9 13 9 1 10 0 9 2
4 13 9 11 11
2 11 2
23 0 0 9 7 0 9 11 11 13 10 9 1 9 12 9 1 9 12 2 9 1 11 2
14 13 13 3 7 1 0 9 15 13 0 9 0 9 2
15 13 3 1 10 9 1 0 9 7 13 0 9 9 9 2
9 1 9 13 9 10 0 9 0 2
30 0 12 9 13 2 3 15 13 2 13 0 9 2 9 9 1 11 2 9 2 9 1 0 9 2 9 7 3 13 2
31 13 1 0 0 9 7 15 13 0 9 2 0 9 2 15 13 0 0 9 7 1 0 9 13 1 9 12 9 11 11 2
14 1 0 9 13 1 9 10 9 7 0 9 9 9 2
10 0 9 15 3 13 16 10 0 9 2
48 4 13 16 0 0 9 2 3 13 1 0 2 11 2 7 1 9 1 0 11 2 13 9 3 3 0 0 9 2 13 0 9 1 0 9 2 13 1 0 9 2 9 2 9 7 0 9 2
25 13 0 9 10 9 2 9 9 2 12 2 7 13 0 0 9 16 3 0 9 1 11 1 9 2
3 3 0 11
2 11 2
28 11 11 11 3 1 9 13 10 0 9 9 12 2 0 9 11 2 7 1 9 1 9 9 3 3 0 13 2
46 2 3 4 15 0 9 13 2 0 4 13 1 0 9 2 2 13 11 1 15 2 16 10 0 9 11 11 11 13 13 12 9 1 9 1 12 2 9 1 0 9 1 10 9 11 2
17 2 11 14 13 9 2 7 3 1 9 13 9 2 2 13 11 2
17 0 9 11 15 3 3 13 9 9 2 7 0 9 11 3 13 2
16 11 9 13 1 11 1 0 9 1 10 0 9 1 9 12 2
13 16 13 2 13 0 9 9 1 12 9 2 9 2
36 2 13 0 15 3 2 16 15 13 13 10 9 2 3 3 13 2 7 3 15 13 15 2 15 13 13 2 2 13 11 0 9 9 1 9 2
8 13 7 15 2 15 13 9 2
19 11 11 13 3 1 11 1 0 9 11 2 7 1 0 9 15 13 9 2
17 11 11 3 3 13 7 0 9 2 16 3 1 9 13 1 9 2
24 1 9 9 9 12 13 3 12 9 2 1 0 12 13 11 12 7 13 1 11 1 12 9 2
5 9 1 9 11 11
5 11 2 11 2 2
30 3 1 0 9 0 15 3 9 12 1 9 9 11 11 1 11 13 9 2 15 13 3 0 9 2 0 12 1 9 2
33 10 9 13 3 13 0 12 9 2 15 15 1 10 9 1 9 13 2 7 9 0 9 1 9 1 9 13 9 9 1 0 9 2
24 9 1 0 9 13 10 9 2 16 9 0 3 0 9 1 9 9 3 13 12 9 7 9 2
13 1 9 4 0 3 13 1 9 0 9 1 11 2
9 13 0 9 1 9 2 13 11 11
14 1 9 9 4 3 13 2 16 0 9 1 9 13 2
19 3 7 13 1 9 9 2 16 4 3 13 9 2 12 1 0 0 9 2
12 2 13 1 15 2 15 15 13 1 9 9 2
31 16 15 13 0 0 9 1 9 9 9 2 9 0 9 7 9 10 9 2 3 13 3 13 2 16 0 11 4 13 2 2
10 1 15 3 3 1 15 13 0 9 2
26 2 9 13 9 2 3 15 1 9 13 0 9 0 9 2 1 15 15 13 0 7 0 9 1 0 2
8 10 9 3 4 7 3 13 2
18 3 10 9 13 3 3 0 2 13 15 2 0 9 2 7 0 9 2
16 7 13 10 0 9 3 13 7 13 7 13 0 9 0 9 2
7 7 15 3 13 9 2 2
14 1 0 9 13 3 1 9 7 0 0 9 7 9 2
13 1 9 1 0 9 4 15 7 1 11 3 13 2
18 2 9 9 3 1 9 13 2 3 16 1 9 9 13 9 0 9 2
18 1 15 13 13 7 15 3 15 13 9 0 9 1 15 2 15 3 2
22 9 13 1 15 2 16 13 3 0 9 9 9 13 3 10 9 2 0 7 0 9 2
22 0 1 15 13 10 9 2 0 13 1 9 10 9 7 13 15 10 9 1 9 13 2
10 9 3 13 1 9 2 15 3 13 2
18 15 13 7 9 0 7 9 0 2 15 0 9 3 13 1 0 9 2
17 9 1 9 9 3 13 3 1 9 9 7 3 1 9 3 2 2
18 7 12 1 0 9 2 0 1 0 9 2 13 1 0 9 3 9 2
23 15 4 3 13 1 15 9 7 0 9 9 2 16 0 9 13 13 0 9 1 10 9 2
9 9 9 11 13 10 9 1 0 2
7 13 3 1 9 0 9 2
8 2 0 9 1 9 3 13 2
7 9 13 3 1 9 0 2
21 9 9 11 15 13 13 1 15 2 16 9 10 3 0 9 13 15 2 10 13 2
10 15 15 2 13 2 13 1 0 9 2
8 15 3 0 4 1 9 13 2
50 3 4 13 2 16 15 13 1 0 9 9 10 9 2 3 3 13 0 2 16 4 15 2 15 13 1 0 9 15 0 2 13 16 0 9 13 15 0 0 9 7 13 1 0 9 1 9 15 0 2
26 7 15 3 3 2 16 4 1 0 9 13 0 9 1 9 0 9 2 1 15 3 9 3 13 2 2
27 13 2 14 7 9 0 9 9 1 11 1 2 0 9 2 2 13 15 3 16 4 9 13 9 1 9 2
9 2 3 3 13 1 9 1 9 2
61 3 13 1 15 2 16 11 11 13 1 0 9 2 13 3 9 13 9 7 13 9 2 7 16 15 1 15 9 13 9 9 2 3 15 13 2 6 2 15 13 3 10 9 2 3 4 15 3 13 2 16 15 13 1 10 0 2 0 9 2 2
10 0 9 7 13 7 9 9 1 9 2
10 2 15 3 15 3 13 2 15 3 2
12 13 7 9 2 16 9 1 9 14 3 13 2
15 10 10 0 9 2 10 9 7 9 13 1 0 3 0 2
8 7 15 13 14 9 9 2 2
9 3 4 3 13 10 9 1 11 2
18 2 13 4 2 16 7 3 15 13 1 0 9 0 9 1 9 2 2
16 13 1 0 2 16 15 1 0 9 13 3 1 15 3 13 2
6 2 15 13 0 9 2
21 15 4 15 1 0 12 9 13 1 0 9 1 3 3 9 16 1 0 9 3 2
33 10 9 13 0 9 2 3 9 1 11 13 15 3 0 7 15 4 13 0 13 15 1 9 9 9 1 10 9 1 0 9 9 2
21 3 13 3 7 12 0 9 2 15 16 15 1 15 13 2 13 15 10 0 9 2
26 1 11 4 15 13 3 1 9 11 2 1 11 13 1 9 1 9 0 9 1 10 9 1 0 9 2
10 7 0 0 9 3 3 13 4 2 2
16 7 9 13 15 1 0 9 13 9 0 9 16 9 9 9 2
29 2 10 9 4 13 9 1 15 2 16 9 15 13 1 0 9 2 1 15 0 13 10 9 7 15 4 13 0 2
15 1 10 9 13 3 13 9 9 2 16 9 11 13 0 2
22 7 15 1 10 0 9 13 1 11 1 9 2 3 15 13 15 13 7 13 0 9 2
8 13 3 9 9 7 0 9 2
12 0 9 3 13 7 13 9 15 3 13 2 2
35 13 13 2 16 0 9 4 13 2 16 4 11 13 9 11 1 9 11 2 13 10 9 1 10 9 1 9 2 16 4 13 3 0 9 2
8 2 9 1 15 10 3 13 2
18 0 9 13 3 1 9 9 2 15 4 13 1 9 9 7 0 9 2
29 13 1 9 2 15 4 13 9 1 15 1 15 2 15 15 15 3 13 13 3 1 9 9 9 7 3 0 9 2
21 3 4 13 9 2 16 15 2 9 14 2 4 13 13 1 0 9 1 15 0 2
10 7 13 2 13 15 14 0 9 2 2
29 13 15 3 1 10 9 0 0 9 2 3 1 12 0 9 13 9 2 1 0 9 7 3 1 15 13 9 9 2
4 13 15 10 2
4 2 3 14 2
23 9 2 9 9 7 15 3 13 9 2 13 9 9 7 15 10 9 3 13 13 3 0 2
41 15 1 15 13 3 12 9 2 0 0 2 15 15 13 13 1 0 7 0 9 2 0 3 13 0 2 0 9 2 15 13 0 14 15 2 16 15 15 15 13 2
37 16 15 3 15 1 9 2 0 9 9 9 13 9 1 9 1 11 2 15 13 1 9 0 0 9 2 3 15 3 13 1 9 7 13 15 4 2
20 15 13 2 16 4 9 9 9 9 2 9 9 7 15 3 13 0 9 2 2
17 13 9 2 16 15 1 0 9 13 9 9 11 0 9 1 9 2
7 2 15 13 0 9 2 2
25 0 9 1 9 7 9 9 15 13 3 1 10 9 2 16 9 13 13 9 1 9 1 0 11 2
15 9 10 9 14 10 9 1 0 9 13 9 11 1 9 2
12 2 13 9 9 9 2 7 1 9 15 13 2
16 13 2 16 9 9 1 3 0 9 13 10 9 13 3 0 2
8 7 0 9 13 0 7 0 2
19 7 10 9 1 0 9 4 13 3 9 11 2 3 0 15 9 1 11 2
25 3 1 10 9 13 1 0 0 13 2 16 13 13 3 0 9 10 9 2 15 3 4 13 13 2
7 15 13 1 15 13 2 2
36 13 7 9 9 2 16 9 13 10 9 13 1 0 9 9 1 0 11 2 3 1 15 11 13 7 15 9 3 13 2 16 0 9 13 0 2
6 2 10 9 3 13 2
17 10 9 13 1 3 15 0 0 9 2 1 15 13 10 9 13 2
16 16 13 3 2 3 15 13 9 2 16 13 2 3 13 9 2
15 10 0 9 1 0 11 13 0 2 7 13 1 0 9 2
9 3 3 15 13 9 2 3 9 2
10 15 13 2 16 13 1 9 10 9 2
24 15 7 1 0 11 2 16 9 9 2 13 13 9 2 7 3 14 15 2 15 13 10 9 2
14 13 13 9 2 15 4 13 3 1 12 10 9 2 2
9 13 15 13 0 9 1 9 11 2
3 2 3 2
9 11 13 3 12 1 0 9 2 2
13 0 9 9 9 15 1 9 9 9 13 11 11 2
16 4 4 13 1 9 10 9 2 1 15 4 13 1 10 9 2
7 15 13 0 9 10 9 2
12 2 0 9 4 13 3 7 14 0 9 9 2
26 1 3 0 2 0 9 10 9 9 11 4 13 0 9 1 15 2 16 3 13 1 9 13 9 11 2
4 15 13 9 2
17 9 7 9 1 0 9 7 13 9 2 3 13 0 10 9 13 2
12 1 9 1 9 4 3 1 11 13 0 9 2
22 13 13 2 7 0 9 9 0 9 15 14 13 2 16 9 11 11 13 0 9 2 2
20 0 9 11 15 0 9 13 13 0 9 1 9 7 13 9 9 9 11 11 2
24 13 7 9 9 9 1 15 2 16 9 13 13 10 9 2 10 9 0 9 9 1 9 9 2
7 2 15 15 1 15 13 2
35 16 4 13 13 0 9 2 13 4 1 15 3 9 15 2 16 13 1 9 0 9 2 16 9 9 15 13 3 13 7 13 10 0 9 2
16 1 10 9 4 13 2 16 0 9 13 0 7 0 9 2 2
17 9 7 13 13 9 1 9 2 13 9 2 13 13 7 0 9 2
13 3 3 9 13 2 16 0 1 9 13 9 11 2
27 2 10 9 2 15 13 13 2 13 11 7 0 9 2 15 4 13 3 2 16 4 0 9 13 3 9 2
27 1 0 9 13 2 16 9 9 9 13 3 9 1 9 2 3 13 1 9 9 7 0 9 3 9 2 2
13 13 15 9 10 0 9 1 0 9 7 0 9 2
6 2 10 9 13 0 2
15 3 4 13 15 1 15 2 16 4 9 13 0 7 0 2
17 7 1 0 9 1 15 7 9 9 13 13 1 0 9 0 9 2
16 16 13 2 16 9 1 9 4 3 13 2 4 13 0 2 2
3 13 11 11
10 0 2 0 9 2 0 15 10 9 13
5 11 2 11 2 2
25 16 1 9 12 13 0 9 1 11 1 0 9 9 12 9 9 2 3 3 13 15 1 12 9 2
16 13 15 3 9 9 11 11 1 9 1 10 0 9 11 11 2
21 2 9 11 2 3 7 11 2 15 1 9 1 9 13 16 1 9 10 0 9 2
17 15 15 13 16 9 9 7 9 13 15 1 11 2 2 13 11 2
15 1 9 0 9 13 0 9 9 0 9 2 7 0 9 2
13 2 0 9 13 3 0 2 7 13 7 10 9 2
19 13 10 9 2 15 13 3 0 9 2 13 15 9 2 9 7 0 9 2
17 1 9 15 13 13 1 0 9 7 13 0 9 2 2 13 11 2
17 0 9 13 2 16 3 9 9 11 1 11 4 13 0 0 9 2
6 0 9 9 3 13 9
5 11 2 11 2 2
18 14 1 0 9 15 13 1 9 9 9 1 11 1 9 0 0 9 2
18 3 13 4 0 9 1 9 13 2 7 1 1 0 9 4 9 13 2
21 1 9 9 1 0 9 15 7 4 13 9 2 16 15 13 1 0 9 9 11 2
14 9 15 13 1 12 9 7 13 0 9 12 9 9 2
17 1 0 9 13 9 9 2 15 13 7 1 12 2 9 1 9 2
14 9 11 2 15 4 9 13 2 13 1 9 0 9 2
11 15 7 13 4 13 2 7 13 0 9 2
15 3 13 1 12 9 9 2 1 15 15 13 9 9 11 2
15 16 4 4 13 0 9 2 13 9 11 9 1 9 9 2
24 1 12 9 15 13 9 11 2 15 16 0 13 0 1 12 9 13 9 1 9 12 9 9 2
18 2 9 4 15 13 1 12 0 9 2 2 13 9 9 11 11 11 2
19 2 13 13 2 16 7 1 9 9 4 13 13 1 9 9 3 9 9 2
8 3 3 13 9 9 10 9 2
21 13 15 2 16 9 4 13 4 1 9 13 2 7 13 4 1 15 13 0 9 2
18 13 15 14 9 9 2 7 13 7 9 2 15 4 13 1 0 11 2
18 9 15 13 1 9 9 7 12 9 9 1 15 13 9 0 9 2 2
16 1 11 11 1 9 11 13 0 9 1 9 0 9 9 9 2
6 9 1 9 13 9 9
5 11 2 11 2 2
34 9 9 2 15 4 13 4 1 9 9 1 9 0 9 7 9 1 15 13 1 0 9 0 1 0 9 2 13 3 0 16 10 9 2
19 13 3 1 9 2 10 9 4 3 2 1 2 0 2 9 2 4 13 2
26 9 9 7 9 11 11 3 13 9 1 9 0 9 2 16 2 13 15 0 9 11 1 12 9 2 2
17 9 11 13 2 16 9 1 10 0 9 2 13 3 0 9 2 2
13 3 7 11 13 2 16 13 3 2 16 9 13 2
31 1 10 9 10 9 2 15 1 10 9 13 2 15 3 4 13 1 0 9 13 9 2 2 1 10 9 13 10 9 2 2
46 0 9 1 9 7 9 9 1 0 9 1 9 9 12 7 12 2 0 1 0 9 2 3 13 1 12 12 9 2 1 15 4 15 13 13 9 0 9 1 0 9 0 1 0 9 2
18 9 9 11 11 15 13 2 16 1 9 15 13 13 3 12 1 15 2
6 2 9 13 3 0 2
26 16 13 1 9 9 1 0 9 2 15 15 13 13 2 13 0 2 2 13 15 9 0 9 11 11 2
5 9 1 9 2 12
3 9 1 11
2 11 2
27 9 9 0 2 9 2 11 1 11 2 3 13 9 7 0 9 0 9 2 3 13 9 1 9 11 11 2
25 1 12 9 1 9 11 13 0 9 11 2 1 15 13 1 11 11 11 13 9 10 9 1 11 2
3 9 1 11
5 11 2 11 2 2
9 0 9 0 9 15 13 11 11 2
16 1 9 0 9 13 1 9 0 9 10 9 9 11 11 12 2
2 9 9
5 11 2 11 2 2
13 9 9 0 9 0 1 11 13 3 0 0 9 2
12 13 15 15 12 9 2 1 12 1 12 9 2
17 9 13 3 9 1 9 2 9 9 2 9 1 0 9 7 3 2
7 9 13 0 9 1 9 9
6 0 11 2 11 2 2
18 1 12 9 11 3 13 12 7 12 12 9 1 0 9 1 9 9 2
28 10 9 13 1 9 0 0 9 1 9 0 9 2 15 13 1 9 12 2 12 0 9 7 9 2 3 0 2
16 1 10 0 9 13 9 7 0 9 13 7 0 9 0 9 2
12 3 0 9 13 1 9 1 9 9 2 9 2
17 9 13 7 3 0 1 9 1 0 9 7 1 9 1 0 9 2
16 0 9 9 13 1 0 0 9 1 0 9 0 7 0 9 2
6 9 1 9 1 0 9
9 1 0 9 11 15 1 9 13 9
2 11 2
8 1 9 9 15 3 9 13 2
12 3 4 10 9 3 13 1 9 0 11 11 2
21 1 9 11 2 15 13 1 10 9 1 11 2 3 13 11 9 9 9 12 9 2
18 16 1 9 9 1 12 9 9 3 13 9 2 9 1 9 10 9 2
7 9 3 13 7 1 9 2
24 1 15 15 13 9 10 9 1 0 9 9 11 11 2 15 1 9 13 3 2 11 7 11 2
12 0 0 9 13 0 9 11 11 2 12 2 2
20 15 7 3 1 9 13 0 9 1 9 0 0 9 11 11 2 3 12 2 2
23 1 15 13 0 0 9 9 1 0 9 1 11 2 3 13 1 9 14 1 12 2 9 2
19 3 7 13 1 9 12 0 9 9 7 10 0 9 1 9 9 1 11 2
8 3 1 15 15 3 13 9 2
20 9 13 11 11 13 1 11 2 3 13 1 0 11 7 13 9 1 11 11 2
28 14 1 0 9 13 2 0 2 0 9 11 9 12 9 2 9 0 2 15 13 3 11 2 13 9 12 9 2
19 1 0 0 9 1 0 9 1 11 7 13 11 3 12 9 1 0 9 2
11 3 13 12 9 2 12 9 7 12 9 2
42 0 9 13 0 2 0 2 0 9 2 0 13 0 0 9 7 3 0 0 9 11 2 3 1 9 12 9 2 7 3 0 9 3 0 9 2 15 3 0 9 13 2
20 1 12 9 15 11 2 13 2 3 9 9 1 9 9 1 11 1 2 11 2
24 3 3 13 1 15 2 3 13 1 9 2 2 3 15 13 2 13 4 2 16 1 15 13 2
19 13 4 9 12 9 2 3 3 3 2 7 15 3 13 3 0 9 2 2
19 1 9 1 9 7 9 1 9 11 13 2 2 10 12 9 15 13 13 2
5 9 13 3 0 2
10 3 15 2 16 13 1 12 0 9 2
9 1 9 13 0 15 13 9 2 2
11 3 1 9 13 7 11 11 3 1 9 2
19 2 16 15 13 3 3 2 2 13 9 11 2 2 13 13 7 12 9 2
15 13 2 16 4 9 13 3 2 16 4 15 9 13 2 2
15 1 9 0 0 9 4 7 7 0 12 9 14 15 13 2
17 7 2 3 3 13 14 9 2 3 4 7 9 13 12 9 2 2
3 13 9 9
13 3 13 3 0 2 16 1 0 9 13 9 9 2
25 1 0 0 9 1 9 2 3 15 13 1 12 9 9 9 1 0 9 2 13 9 0 9 3 2
27 1 0 9 0 2 9 15 13 1 9 1 12 9 9 7 15 13 3 9 2 15 13 0 13 1 9 2
16 3 15 3 13 13 2 7 13 1 0 1 0 9 9 9 2
21 13 9 0 9 1 9 1 0 2 15 4 14 3 3 13 9 7 0 0 9 2
11 3 15 13 10 9 1 15 9 1 9 2
14 13 15 9 9 2 0 9 7 9 7 3 0 9 2
21 13 15 3 3 10 9 2 15 1 0 9 13 1 9 3 13 7 13 0 9 2
29 4 13 1 9 9 9 2 1 9 7 9 9 0 1 0 0 9 2 15 2 3 13 10 9 2 7 3 3 2
8 15 13 15 0 7 0 9 2
10 13 15 13 13 15 1 9 0 9 2
26 13 0 9 0 9 2 3 13 0 9 2 0 9 2 0 9 2 1 0 9 3 9 7 3 3 2
18 1 0 9 15 3 13 3 3 16 9 9 2 15 13 3 3 0 2
8 13 15 0 2 7 0 9 2
18 0 9 13 3 0 9 0 9 0 9 2 1 15 3 13 3 9 2
46 1 9 9 1 9 7 1 0 9 3 13 3 9 2 3 15 1 0 9 3 3 13 12 1 0 9 0 9 2 9 13 1 10 9 3 3 2 16 4 15 13 9 7 9 9 2
4 9 9 3 13
5 11 2 11 2 2
29 1 9 7 9 4 13 3 12 9 1 9 0 9 2 0 2 9 2 1 9 2 1 12 9 9 1 15 13 2
9 13 1 15 3 9 9 11 11 2
14 1 0 9 13 12 0 7 12 1 0 0 9 9 2
16 14 1 9 9 1 9 0 9 7 10 9 4 13 12 9 2
3 9 1 11
5 11 2 11 2 2
21 0 0 9 1 15 7 3 7 0 0 9 13 1 0 9 1 11 0 9 9 2
45 1 0 9 1 9 3 12 9 0 7 0 9 9 1 9 2 9 1 9 2 0 9 1 9 0 9 7 0 9 15 9 9 11 11 13 0 9 1 9 12 7 12 9 9 2
13 9 9 13 7 0 9 0 0 9 9 0 9 2
4 9 9 1 11
2 11 2
32 0 9 9 11 11 11 7 10 0 9 1 9 11 11 11 4 3 13 0 11 1 9 0 0 9 0 9 1 0 9 11 2
33 11 7 0 0 9 11 2 12 13 2 16 1 15 12 4 1 9 13 3 0 9 11 11 2 1 15 11 13 2 16 13 13 2
11 3 13 13 3 0 9 2 0 9 11 11
2 11 2
24 0 9 11 11 11 4 3 13 1 9 2 16 15 13 13 1 9 9 2 15 13 0 9 2
11 1 3 0 9 13 0 12 0 9 13 2
14 1 9 13 14 3 0 9 7 9 0 7 0 9 2
30 9 0 9 1 0 9 11 2 3 4 1 12 9 13 12 0 9 0 9 11 2 3 13 12 9 9 11 7 9 2
23 0 9 9 7 1 0 9 3 13 9 0 0 9 2 15 4 13 10 9 1 0 9 2
9 9 13 3 9 0 9 11 11 2
26 0 9 13 3 2 16 15 9 0 9 1 11 13 13 2 16 1 0 9 11 15 13 0 0 9 2
35 11 11 11 4 1 10 9 13 2 16 16 1 9 1 0 9 11 1 11 13 1 9 10 9 2 13 0 0 9 1 9 10 9 9 2
19 0 9 11 11 13 2 16 1 0 9 13 13 12 11 7 0 12 13 2
36 1 10 9 7 11 13 7 13 2 7 13 1 9 1 9 2 3 15 13 9 0 9 11 2 0 0 9 2 11 2 9 2 1 10 9 2
10 10 9 7 13 0 13 1 0 9 2
15 1 0 9 13 0 9 11 9 12 9 7 9 0 12 2
8 1 12 9 13 9 7 9 2
10 0 0 9 0 9 15 13 7 1 11
2 11 2
26 9 9 7 9 1 10 0 9 4 13 1 9 7 9 1 0 9 4 3 13 1 0 7 0 9 2
12 13 15 3 1 9 1 0 7 0 0 9 2
12 11 13 0 9 9 2 3 1 11 7 11 2
32 0 9 13 1 9 0 0 9 7 0 11 2 0 9 4 13 1 11 2 11 2 11 2 11 2 11 2 11 7 0 11 2
4 9 9 7 9
26 13 3 3 2 16 15 2 0 9 2 13 13 9 1 0 9 3 9 9 2 1 0 9 3 9 2
34 0 12 9 2 7 0 9 0 0 9 2 3 15 1 15 3 7 3 13 2 13 3 0 2 1 0 0 9 7 14 3 3 0 2
14 3 15 13 3 1 9 16 1 9 0 7 0 9 2
19 7 1 0 9 15 9 0 13 1 9 7 2 3 1 9 2 1 9 2
21 2 3 2 13 15 2 3 15 1 0 9 9 13 3 16 1 0 9 2 2 2
14 9 10 9 13 9 2 1 15 13 0 9 7 9 2
27 13 7 9 9 1 0 0 9 2 3 2 1 9 1 15 13 0 0 9 3 0 9 16 9 7 9 2
44 1 0 9 10 9 13 3 0 9 9 2 0 9 2 15 15 9 10 9 3 13 1 9 2 13 10 0 9 2 13 1 9 7 9 2 13 15 3 0 9 7 13 9 2
62 0 9 13 2 16 15 13 1 9 1 0 9 2 0 9 2 0 9 1 9 2 1 11 2 11 2 11 2 1 0 9 9 2 1 0 9 16 13 0 9 7 0 9 2 1 9 2 9 2 9 2 9 2 9 14 2 9 2 7 1 9 2
28 9 2 2 1 0 2 0 0 9 2 2 15 13 2 2 2 9 2 2 2 10 9 2 16 4 13 9 2
26 9 2 2 0 9 2 2 13 1 9 0 9 10 0 9 2 15 3 13 1 10 0 2 9 2 2
23 14 15 9 3 3 13 3 2 0 4 15 13 9 9 2 16 9 7 9 13 10 9 2
42 13 15 2 16 15 2 9 2 9 13 3 0 9 2 16 15 13 0 7 0 2 16 15 7 13 1 2 0 2 9 0 9 7 9 13 0 9 10 9 3 0 2
26 16 13 1 9 2 13 15 2 16 13 1 3 0 9 2 9 13 2 14 0 0 9 13 3 0 2
20 0 9 11 11 13 9 9 2 15 4 10 0 9 1 10 9 13 0 9 2
21 9 13 3 0 13 0 9 9 7 9 2 10 9 15 3 13 13 9 10 0 2
15 2 9 13 2 16 15 13 15 2 3 1 9 9 2 2
21 10 9 4 13 2 9 9 2 1 10 9 1 0 0 9 2 3 9 1 9 2
58 3 4 9 13 3 0 0 9 2 2 13 2 4 15 2 15 15 13 13 0 9 14 15 3 7 3 13 9 2 13 2 9 2 13 2 2 3 14 15 3 2 9 10 9 2 15 0 4 13 14 0 2 0 7 3 0 9 2
36 10 0 9 4 13 1 9 7 9 2 7 13 4 10 0 0 9 2 0 9 9 2 9 2 15 4 15 13 7 1 10 0 9 7 9 2
25 7 15 15 4 13 3 3 16 10 0 9 2 16 16 9 1 15 2 3 2 7 2 3 2 2
24 9 15 2 15 2 4 13 7 3 0 2 0 2 0 2 2 16 3 0 2 0 2 0 2
18 0 9 0 9 15 13 13 2 16 9 9 15 13 1 10 0 9 2
8 1 15 15 1 10 9 13 2
33 3 1 15 3 16 1 9 2 3 3 4 13 1 12 0 9 9 2 0 1 10 9 2 15 15 9 2 3 3 3 2 13 2
32 13 15 7 9 2 3 0 13 13 2 13 2 14 1 2 0 2 9 7 3 15 13 3 10 9 9 2 15 13 15 0 2
39 9 13 3 0 2 9 0 9 2 0 9 2 7 14 9 2 16 9 1 0 9 9 2 7 9 0 2 0 3 16 0 9 2 9 2 9 9 2 2
13 9 3 13 9 2 1 15 1 15 15 3 13 2
4 11 11 2 11
4 9 1 0 9
7 1 15 13 0 9 0 2
2 11 11
29 9 9 2 7 2 9 9 3 2 16 4 13 0 14 9 0 2 2 9 2 2 2 13 0 2 0 7 0 2
16 0 3 3 3 14 1 9 2 7 3 1 9 9 1 9 2
16 13 15 3 13 1 12 0 9 9 2 0 1 9 0 9 2
25 13 1 9 0 9 2 15 3 13 2 16 3 13 2 0 2 7 14 3 0 2 9 0 9 2
3 9 0 9
21 13 13 9 0 9 2 1 15 3 13 14 15 2 16 13 0 16 13 12 9 2
20 1 9 4 13 2 16 9 4 13 3 2 7 2 1 12 9 12 7 12 2
22 2 16 15 1 9 13 1 0 9 2 13 15 13 1 0 9 9 1 0 9 2 2
26 9 9 12 7 12 2 3 1 9 7 9 1 0 9 2 13 15 2 16 15 13 13 1 0 9 2
22 12 5 12 5 12 2 12 5 12 5 12 5 12 5 12 2 12 5 12 5 12 2
42 3 13 2 3 4 0 9 13 2 7 13 15 13 15 2 16 1 15 7 9 13 0 9 2 7 2 0 9 9 7 9 1 9 12 9 2 13 9 2 12 2 2
27 0 9 13 13 3 2 3 2 16 13 9 7 13 12 5 9 7 12 5 9 15 2 3 0 9 13 2
13 15 7 9 4 3 13 9 2 15 3 3 13 2
29 1 9 2 3 13 1 9 0 0 9 2 13 15 9 0 9 2 13 9 2 12 2 7 3 15 3 3 13 2
21 13 2 14 9 0 16 12 9 2 3 3 13 14 10 0 9 7 9 9 13 2
16 9 2 15 15 13 0 9 2 7 13 9 2 15 13 15 2
19 13 2 14 9 3 3 0 9 9 7 9 2 13 7 0 9 3 0 2
6 9 1 15 3 13 2
31 7 15 13 1 0 9 9 2 7 15 13 0 9 2 16 13 2 14 3 15 2 13 0 9 2 13 2 9 2 12 2
22 2 13 15 2 16 13 14 12 5 12 5 12 2 7 3 12 5 12 5 12 2 2
15 9 10 9 13 0 9 9 2 16 15 13 3 13 9 2
6 13 7 7 10 9 2
17 13 2 14 1 9 9 0 16 12 9 2 13 9 3 1 9 2
17 13 3 9 13 3 1 9 2 7 1 15 3 13 9 15 13 2
14 3 0 9 2 3 3 0 2 9 13 13 3 0 2
3 9 0 9
35 9 2 12 13 11 2 11 11 2 11 2 11 7 11 2 11 2 11 9 2 1 15 15 0 9 13 2 7 3 15 9 1 9 13 2
15 9 4 13 1 0 9 0 9 2 13 0 9 0 9 2
28 15 13 3 0 2 7 13 1 12 1 0 0 9 2 15 15 3 9 13 2 0 9 13 1 9 9 9 2
25 3 1 12 0 9 2 15 13 9 12 9 2 13 10 9 7 0 9 3 16 1 9 9 9 2
13 13 4 2 16 13 0 9 2 3 13 3 0 2
19 7 16 13 1 9 3 0 2 13 15 2 16 1 9 4 0 9 13 2
30 1 0 9 7 13 0 9 9 1 9 9 1 12 7 0 0 9 13 14 14 2 13 2 1 0 9 10 10 9 2
21 13 10 9 7 1 9 0 9 15 3 2 2 2 12 13 2 13 9 7 9 2
21 10 9 3 13 2 7 13 10 9 9 5 9 2 9 2 15 13 1 12 9 2
22 9 2 16 7 1 9 9 9 13 9 13 9 9 7 9 2 13 1 0 0 9 2
25 16 9 10 9 13 10 0 9 9 2 3 9 5 12 2 3 9 5 12 7 9 5 12 2 2
16 15 3 15 13 2 7 4 1 10 0 9 13 0 9 9 2
22 13 2 16 9 4 13 1 9 12 2 12 2 12 2 2 2 2 2 9 2 12 2
12 2 13 2 14 13 1 0 9 2 13 15 2
27 3 2 1 9 5 12 9 0 1 0 9 13 1 9 0 2 7 9 13 10 9 1 9 2 3 2 2
27 1 9 9 2 0 2 7 9 2 9 2 0 2 13 3 12 0 9 9 2 3 16 4 13 0 16 9
16 9 2 9 2 5 2 9 2 12 2 2 2 9 2 12 2
18 7 16 4 12 9 9 2 12 7 9 2 12 13 1 9 7 0 2
48 2 3 2 13 2 14 9 5 12 2 13 9 12 9 9 9 2 16 9 2 12 2 5 12 2 12 5 12 2 13 13 1 9 12 2 12 2 12 2 12 2 12 2 12 2 12 2 2
44 1 9 9 13 0 2 16 1 0 10 9 9 9 13 3 12 9 9 0 16 9 2 9 2 2 1 15 13 2 16 9 9 2 9 2 12 13 0 9 9 2 9 2 2
20 2 3 2 13 2 14 9 5 12 7 9 5 12 2 13 9 5 12 2 2
29 9 9 13 0 2 7 13 15 3 13 2 9 9 13 0 2 7 15 13 2 16 4 15 15 13 13 0 9 2
31 16 13 9 9 3 0 0 9 7 2 13 4 1 9 9 9 2 9 2 2 13 2 1 9 9 9 7 9 2 13 2
25 13 2 14 9 9 7 9 2 13 13 2 9 0 9 13 1 9 2 10 7 9 13 9 9 2
11 9 1 10 9 13 0 9 7 15 13 2
24 13 2 14 3 9 9 2 13 3 13 2 0 9 13 1 9 2 10 7 9 13 9 9 2
9 9 1 10 9 13 0 0 9 2
10 0 10 9 4 13 1 9 2 12 2
7 9 0 9 13 0 9 2
20 13 13 7 0 9 2 7 3 9 2 16 14 12 9 9 2 9 7 9 2
6 9 13 3 3 0 2
45 13 2 14 3 12 9 9 7 9 1 12 9 7 0 9 9 2 13 2 0 2 9 13 2 16 13 0 9 9 9 5 9 2 9 2 7 15 15 15 13 1 0 9 2 2
25 0 9 13 15 2 16 13 13 15 2 16 1 0 9 13 9 13 7 16 0 9 9 9 2 2
29 0 9 2 15 10 9 13 2 13 9 0 9 1 0 9 2 9 7 9 2 2 15 15 1 9 7 9 13 2
9 7 13 1 9 3 3 0 9 2
2 9 2
10 11 2 11 2 9 2 11 11 12 2
4 3 9 13 2
18 1 11 15 9 13 13 3 1 9 9 2 16 9 13 3 0 9 2
20 1 9 7 9 1 0 9 13 3 12 9 9 7 3 0 13 7 0 9 2
22 12 1 0 9 9 13 9 2 3 15 16 3 3 13 9 7 16 15 13 14 3 2
24 7 14 0 9 9 9 7 9 9 13 13 9 0 9 7 3 10 9 14 1 10 9 9 2
12 3 12 9 15 1 0 10 9 9 13 3 2
25 9 13 0 9 3 1 12 2 12 5 7 3 0 9 13 0 9 2 0 9 4 13 3 9 2
5 9 13 14 3 2
39 13 15 2 16 0 9 9 9 13 1 9 0 9 0 9 2 9 12 2 12 2 12 2 12 2 2 15 7 3 13 13 1 9 2 3 9 3 13 2
29 13 15 2 16 13 13 10 0 0 9 2 2 0 2 11 2 15 9 13 1 0 0 9 3 1 12 9 9 2
31 11 2 11 7 11 2 11 2 11 1 9 1 11 2 11 2 11 13 10 9 1 9 1 0 7 0 9 0 1 9 2
35 9 0 1 0 9 0 13 0 9 0 9 7 15 9 13 1 9 2 16 0 9 0 13 1 9 9 0 9 7 15 15 13 1 9 2
12 11 12 2 12 2 12 2 12 2 12 2 12
4 9 0 9 9
38 0 0 9 2 15 13 9 9 0 1 9 2 13 0 9 2 15 13 9 0 0 1 0 9 1 0 9 0 9 7 15 13 3 0 9 0 9 2
29 0 9 7 1 9 10 9 13 3 9 2 3 12 9 9 1 12 9 9 2 2 9 7 1 0 9 3 9 2
33 11 2 11 2 11 1 10 9 13 2 16 3 0 9 0 0 9 1 0 9 13 9 0 9 2 15 3 13 0 9 9 0 2
36 0 9 13 2 16 4 4 1 0 9 2 15 13 9 0 9 12 2 13 9 0 9 9 2 15 9 4 13 9 9 12 0 9 0 9 2
24 1 0 9 13 3 0 9 2 15 3 13 11 2 11 11 1 10 9 9 1 9 0 9 2
22 7 1 3 0 9 2 16 13 9 9 1 10 9 2 13 2 10 9 13 9 9 2
20 9 1 10 9 13 1 9 0 9 2 15 13 0 7 0 9 3 0 9 2
8 13 9 10 9 13 3 0 2
30 0 9 13 1 0 9 7 1 0 0 9 1 0 9 9 9 12 9 7 9 12 9 0 1 0 9 1 9 12 2
20 3 9 0 0 1 0 9 7 0 15 3 9 3 13 9 9 0 9 9 2
31 10 9 13 7 2 14 2 3 0 2 16 4 0 9 13 13 1 9 3 10 9 9 2 16 4 15 13 3 0 9 2
10 0 0 9 12 2 12 2 12 2 12
10 9 0 0 9 2 12 2 12 2 12
5 0 9 7 9 9
26 0 9 9 13 2 16 9 13 12 9 9 2 7 16 0 9 4 13 14 1 9 1 12 9 9 2
20 0 9 11 2 11 11 7 11 2 11 7 13 0 0 9 1 12 9 9 2
33 13 15 1 0 9 9 2 15 13 3 0 14 12 9 0 0 9 2 15 1 10 9 13 3 12 2 12 5 0 0 9 9 2
18 9 13 0 9 2 16 3 13 1 12 1 0 9 9 0 0 9 2
15 10 0 9 15 13 1 0 9 0 9 7 0 0 9 2
19 13 3 0 0 9 9 7 4 1 15 13 3 2 1 11 7 0 11 2
45 0 9 9 13 2 16 0 0 9 13 1 10 9 15 9 0 1 9 7 3 1 9 0 9 12 5 1 9 12 5 13 13 1 9 9 9 1 9 7 15 1 9 0 9 2
31 9 9 9 7 0 9 9 0 9 13 9 3 0 9 1 0 12 9 9 1 9 7 13 7 0 9 1 0 0 9 2
12 11 12 2 12 2 12 2 12 2 12 2 12
11 9 9 1 9 9 1 0 12 9 9 2
11 9 2 9 2 13 0 9 0 9 9 2
14 13 15 0 9 1 9 9 1 12 7 12 9 9 2
19 0 9 13 9 1 9 9 2 0 9 13 9 9 9 1 1 0 9 2
12 0 9 0 9 13 9 0 9 9 0 0 9
5 9 9 1 0 9
27 0 9 13 0 9 9 9 0 1 9 7 9 9 2 15 13 16 0 9 0 9 7 13 1 9 9 2
25 7 15 3 13 2 3 0 9 13 1 9 9 0 9 2 12 2 12 9 2 0 9 0 9 2
23 9 14 1 12 5 15 13 1 0 9 2 3 1 9 0 1 9 2 13 2 0 9 2
12 0 9 0 9 1 0 9 13 3 3 0 2
26 9 0 9 13 1 9 10 9 7 9 0 9 13 0 1 9 2 15 15 13 13 7 1 10 9 2
12 9 3 13 1 9 2 7 4 13 0 9 2
21 0 9 3 13 9 9 7 0 9 3 0 0 0 9 2 15 13 9 0 9 2
19 13 3 9 2 16 9 1 0 9 0 9 11 15 13 3 9 9 9 2
6 0 9 13 3 0 2
25 0 9 9 9 12 5 12 12 9 1 9 9 0 9 3 13 3 10 9 0 0 9 0 9 2
8 11 12 2 12 2 12 2 12
7 15 15 0 0 2 2 2
27 1 9 2 12 11 11 13 1 9 11 2 11 1 9 10 9 2 11 12 2 12 2 12 2 12 2 2
39 0 9 11 2 11 7 11 2 11 13 1 9 9 10 9 2 16 3 0 9 1 9 9 0 9 9 0 13 0 9 2 3 15 9 13 9 9 9 2
16 9 1 0 0 0 9 1 9 9 13 1 0 9 3 0 2
14 2 9 4 14 13 0 13 0 2 0 9 2 2 2
13 12 9 13 9 9 3 9 1 9 1 0 9 2
35 1 9 10 9 13 9 0 9 9 0 2 15 15 1 0 9 13 9 1 0 9 16 10 3 0 9 9 0 2 9 0 7 9 0 2
13 7 9 2 15 13 9 13 2 13 1 3 0 2
21 3 13 2 16 0 9 13 14 12 5 9 2 1 15 15 13 9 2 1 9 2
23 13 3 3 2 16 0 9 9 0 9 9 9 13 7 1 9 2 7 1 0 9 9 2
6 11 12 2 12 2 12
8 2 2 2 7 15 3 3 0
14 1 10 9 11 13 0 9 3 0 2 0 2 9 2
19 1 15 13 9 3 9 9 0 1 0 9 2 15 13 9 12 9 9 2
34 13 15 2 16 9 4 13 1 9 1 12 9 9 7 16 1 12 9 9 13 13 10 0 9 2 7 13 14 14 13 0 0 9 2
15 3 9 10 0 9 0 13 13 9 9 0 9 9 9 2
18 13 7 1 9 0 9 9 9 2 15 3 3 13 3 3 0 9 2
8 11 12 2 12 2 12 2 12
6 9 2 0 2 9 2
17 9 1 0 9 0 9 1 9 1 12 9 13 13 9 0 9 2
27 16 0 9 4 13 1 3 16 12 9 2 9 9 15 13 3 1 9 2 16 3 15 13 0 10 9 2
17 3 15 13 9 2 16 15 13 9 1 9 2 16 13 1 9 2
19 9 9 1 15 13 3 0 2 0 9 13 12 2 12 9 1 0 9 2
17 1 0 0 9 0 9 2 12 7 12 9 2 13 7 3 0 2
21 1 9 1 12 9 4 9 1 9 3 13 9 1 0 9 1 9 0 0 9 2
17 1 9 1 12 9 4 9 3 13 7 9 9 4 13 1 9 2
42 11 2 11 2 11 2 11 2 11 2 11 13 1 9 2 12 1 9 2 12 9 0 9 7 13 2 16 9 10 9 13 1 9 1 12 9 2 3 9 2 3 2
7 9 15 13 9 0 9 2
26 1 9 9 0 9 1 12 9 2 1 9 12 2 12 2 13 3 2 13 9 0 9 1 12 9 2
6 11 12 2 12 2 12
6 11 13 9 1 0 9
18 1 1 0 0 9 9 1 0 9 4 13 9 1 9 9 0 9 2
14 3 9 1 0 9 16 12 1 12 13 13 0 9 2
24 0 9 0 9 3 13 2 16 10 9 4 13 13 9 9 2 7 3 0 9 2 9 2 2
29 9 13 9 2 2 15 13 3 0 1 9 2 3 10 9 16 11 2 11 7 11 13 9 9 0 0 9 2 2
6 11 12 2 12 2 12
9 3 13 9 0 9 1 0 9 2
41 1 12 2 0 9 0 9 0 9 2 11 2 1 9 2 0 9 1 0 0 9 2 15 1 9 12 13 1 11 12 9 7 9 0 9 1 12 9 15 9 2
47 1 9 0 7 0 9 15 9 0 9 2 9 12 2 12 2 12 2 13 3 3 2 16 4 15 9 7 0 0 9 13 10 0 7 0 9 2 10 9 1 10 9 15 13 1 0 2
39 0 9 13 3 1 12 2 12 9 9 7 0 9 9 2 14 9 2 0 9 0 9 7 0 9 2 1 15 9 3 2 13 9 1 0 7 0 9 2
22 13 15 15 3 9 2 9 7 9 1 0 7 0 2 0 7 0 2 9 0 9 2
25 1 9 15 13 2 16 13 3 13 14 1 9 9 2 7 7 0 9 1 0 9 13 3 9 2
14 9 13 13 9 2 7 13 15 9 3 0 0 9 2
42 1 10 9 9 13 7 9 0 9 7 9 9 2 3 13 2 16 15 10 9 9 9 13 1 9 2 0 9 4 1 15 3 3 7 3 13 7 1 9 0 2 2
28 0 13 0 9 2 15 13 0 9 1 0 9 2 3 9 9 1 9 1 9 7 9 2 1 0 9 2 2
11 9 13 3 13 2 16 1 0 13 9 2
32 9 0 9 1 9 0 9 13 2 16 1 0 9 0 9 9 13 1 3 7 3 0 0 13 15 9 2 1 0 9 2 2
42 1 9 1 0 0 7 0 9 2 3 9 7 9 0 9 13 9 15 0 0 9 2 4 1 9 3 3 0 9 2 7 3 2 9 0 9 2 13 3 0 9 2
16 9 7 0 9 9 15 3 13 3 0 9 0 9 7 9 2
39 15 0 2 7 2 9 0 2 0 2 0 2 9 1 9 7 9 2 13 3 3 12 0 9 2 3 9 1 0 9 2 15 13 1 9 3 16 9 2
19 3 0 13 10 9 2 15 13 13 3 2 1 0 2 0 7 0 9 2
55 10 9 15 3 13 7 2 1 0 9 2 2 0 9 9 9 13 1 11 12 9 2 7 1 0 9 14 13 0 9 9 1 9 2 15 13 0 13 7 1 12 9 5 9 2 10 9 15 3 13 0 0 9 2 2
28 13 2 14 9 0 9 3 1 0 9 2 13 9 0 2 13 12 2 12 9 1 12 9 3 10 0 9 2
14 0 9 9 13 13 9 14 1 12 9 1 12 9 2
46 3 15 3 4 3 13 7 9 9 1 11 7 10 9 4 3 3 13 2 16 13 15 1 0 9 9 2 0 9 13 0 7 0 9 1 10 9 9 3 1 12 1 0 9 2 2
2 11 11
42 14 10 9 9 2 15 13 0 9 2 13 10 0 9 2 7 14 15 13 0 2 15 13 0 2 3 15 2 15 13 1 10 9 9 2 1 15 4 15 13 9 2
33 1 15 2 15 13 1 9 2 15 13 14 1 9 2 3 3 2 3 1 15 2 15 15 3 13 13 2 16 3 3 7 3 2
11 1 9 13 9 9 2 1 9 9 9 2
13 9 15 13 14 15 2 15 13 0 2 2 2 2
6 11 11 2 9 1 9
8 11 2 11 12 2 9 2 12
3 9 1 9
21 11 11 2 11 2 0 9 7 0 9 1 0 9 9 9 12 9 2 0 11 12
19 0 9 2 9 1 9 2 13 9 1 0 9 2 15 13 1 15 13 2
28 9 9 13 13 2 16 10 0 9 2 15 13 1 15 2 16 4 1 15 13 2 13 13 7 1 0 9 2
7 9 4 13 1 12 9 2
56 1 0 12 15 11 13 0 9 7 9 2 9 7 9 2 2 15 13 3 7 9 0 9 2 2 0 0 7 0 9 7 9 2 11 15 13 2 0 9 2 2 9 2 15 1 15 1 10 9 13 10 9 1 0 9 2
41 1 10 9 13 0 0 9 2 16 9 13 9 0 9 2 13 3 15 3 13 7 14 15 13 1 9 0 7 0 9 2 2 15 13 7 13 10 9 0 9 2
31 1 10 9 13 11 1 9 3 0 9 2 3 1 9 10 9 13 2 16 15 13 1 0 9 2 15 13 1 15 13 2
17 15 13 2 16 13 13 0 9 0 9 2 15 0 9 13 13 2
23 0 9 3 13 1 15 2 16 13 2 16 15 13 3 0 9 2 15 4 15 13 13 2
8 9 9 13 9 12 7 12 2
32 1 0 9 2 9 0 9 9 2 15 13 9 13 9 2 13 2 15 13 15 9 2 9 2 15 13 9 7 15 13 9 2
24 13 1 9 2 16 1 10 9 13 0 2 16 15 3 13 13 2 7 16 13 10 9 13 2
17 2 3 4 13 13 0 9 3 0 2 2 2 9 2 12 2 2
23 0 13 2 16 4 1 10 9 4 13 9 1 9 2 1 0 9 15 1 15 3 13 2
39 11 7 13 14 12 9 2 9 0 7 0 2 7 13 2 16 13 1 9 3 12 2 16 4 10 10 9 13 3 2 13 2 2 7 3 2 3 2 2
12 0 9 15 13 2 13 4 13 3 2 2 2
19 10 0 9 13 2 16 9 10 0 9 13 0 2 7 3 0 7 0 2
34 9 15 4 1 0 9 3 13 3 3 2 3 1 15 2 16 13 0 9 2 7 3 2 16 1 0 9 15 15 10 9 13 0 2
17 1 11 13 9 0 9 2 9 2 1 9 2 15 13 10 9 2
32 13 0 9 2 15 9 2 9 13 1 0 2 13 15 3 9 2 2 7 13 15 13 3 2 16 4 10 9 13 3 0 2
22 11 3 13 2 16 9 13 9 2 13 9 2 16 3 3 4 13 2 3 15 13 2
6 10 9 15 13 13 2
12 15 3 4 13 2 13 2 2 15 3 13 2
14 15 13 15 2 15 11 13 2 9 0 9 9 2 2
28 0 7 0 9 2 3 13 0 9 2 2 15 13 3 0 7 0 9 0 9 2 3 9 0 9 7 9 2
25 11 13 0 9 1 9 2 15 0 9 13 1 15 2 16 4 10 9 13 1 9 7 9 9 2
30 1 15 13 2 16 9 2 9 2 9 2 13 13 10 0 9 2 15 1 11 13 2 9 16 9 0 9 1 9 2
18 9 3 13 1 10 9 9 2 10 9 13 1 0 9 2 0 2 2
16 1 10 9 13 0 9 9 0 9 1 0 9 12 0 9 2
9 2 13 1 0 9 13 0 9 2
17 3 7 3 1 9 1 0 9 13 9 0 1 0 7 0 9 2
20 13 9 2 1 9 2 9 7 9 2 1 0 9 2 3 13 13 10 9 2
18 4 13 2 16 9 13 9 2 16 13 0 9 2 13 0 9 3 2
22 13 9 2 2 3 13 10 9 2 2 13 11 2 2 7 16 13 15 0 9 2 2
17 13 2 13 2 0 9 2 2 13 3 9 2 2 4 11 13 2
19 2 7 16 10 9 4 15 13 2 13 15 1 0 9 2 13 13 0 2
9 13 15 3 0 9 1 0 9 2
7 9 2 9 2 9 2 2
12 2 13 1 0 9 9 13 1 12 0 9 2
24 0 2 13 2 2 3 16 0 2 13 2 2 13 12 3 0 9 2 15 15 7 3 13 2
19 2 13 7 13 13 3 7 0 9 2 7 15 1 10 9 13 0 2 2
30 2 13 2 13 13 7 2 13 15 0 2 13 15 0 9 1 9 9 2 7 2 13 15 3 2 1 9 0 2 2
11 0 9 4 13 9 0 2 16 0 0 2
15 13 13 9 2 12 2 5 12 2 3 4 15 13 2 2
5 15 13 9 0 2
25 1 15 1 15 4 3 9 9 13 2 16 13 2 13 0 2 16 4 9 2 9 2 2 12 2
5 15 13 9 0 2
19 0 9 1 9 9 3 13 3 3 14 0 9 13 3 2 3 14 0 2
49 11 15 15 10 9 13 1 9 12 7 0 2 7 13 1 9 2 16 0 9 2 15 13 1 15 16 9 0 2 13 9 0 2 3 0 2 0 13 15 2 1 15 13 2 16 13 15 0 2
46 4 2 14 13 0 9 2 13 15 3 13 2 16 9 2 9 2 13 13 0 16 12 2 7 4 2 14 13 3 9 0 2 4 13 2 16 15 15 13 13 9 11 7 11 11 2
22 10 9 13 1 9 1 9 0 9 2 0 13 1 15 15 2 15 13 1 15 0 2
32 9 2 9 4 13 0 0 9 2 3 12 9 9 13 9 1 9 2 7 13 15 13 0 2 15 15 1 9 0 9 13 2
13 16 13 3 3 0 2 13 9 0 7 0 9 2
2 11 11
4 1 9 1 15
17 12 1 0 0 9 2 11 11 2 13 13 1 9 9 2 12 2
46 1 9 1 0 9 2 3 1 9 13 12 1 10 0 9 2 9 2 13 11 11 2 0 9 11 7 11 0 2 9 10 9 2 0 9 7 3 0 9 2 12 2 1 0 9 2
43 13 3 7 1 9 2 13 14 1 0 9 2 7 1 9 9 2 9 9 7 9 9 2 3 9 0 7 0 2 9 9 12 4 13 3 0 9 1 0 9 0 11 2
14 11 13 3 1 9 7 9 7 3 1 9 0 9 2
32 7 3 1 9 0 9 2 15 13 13 1 9 15 9 1 9 2 12 0 14 0 9 9 2 9 2 15 3 13 1 9 2
29 0 0 9 13 3 0 2 13 15 0 9 1 0 0 9 0 9 2 1 15 13 12 0 9 0 1 0 9 2
9 12 9 13 9 2 9 9 2 2
9 0 9 15 1 0 9 3 13 2
37 9 13 1 9 2 13 15 1 9 1 0 9 9 2 0 0 9 2 9 7 0 9 4 13 0 9 2 9 2 9 2 0 0 9 10 9 2
17 3 9 4 13 1 9 2 7 9 13 3 2 3 3 2 0 2
11 16 16 4 7 15 13 9 7 9 9 2
42 7 9 9 13 3 0 7 0 2 9 2 9 12 2 9 2 9 9 2 9 2 9 9 2 2 2 2 9 9 3 13 2 9 9 2 9 2 9 2 0 9 2
20 15 4 13 16 9 9 2 9 2 0 9 2 9 2 9 7 0 0 9 2
13 15 15 13 13 9 2 7 3 15 13 15 13 2
23 3 9 2 9 2 9 13 13 0 9 10 9 2 3 3 3 2 16 10 9 4 13 2
19 7 15 10 9 13 9 9 9 2 10 9 7 9 9 2 9 7 9 2
21 0 9 2 9 7 9 1 15 13 15 2 7 3 3 0 9 2 9 7 9 2
66 13 15 15 3 2 16 0 9 11 11 13 12 0 9 3 2 9 2 15 4 3 13 2 1 9 1 15 2 2 9 1 3 3 0 7 0 9 2 0 15 1 9 2 1 9 2 0 14 1 0 9 2 0 1 9 2 0 2 0 9 2 7 15 3 9 2
18 15 3 13 9 2 9 2 15 3 13 15 15 2 15 0 1 15 2
9 13 9 2 16 0 9 13 13 2
27 3 14 3 16 1 15 15 2 15 13 7 15 15 2 15 0 1 15 2 13 13 9 1 9 0 9 2
20 7 3 13 1 0 9 1 9 9 2 9 7 9 2 7 1 9 7 9 2
2 11 11
6 13 15 2 13 0 2
2 11 11
19 3 3 15 13 2 16 9 2 9 7 9 13 9 2 14 16 3 13 2
24 3 3 7 4 3 13 7 0 9 10 9 2 0 9 2 9 7 9 13 13 7 13 9 2
21 9 2 15 13 2 13 10 0 9 7 13 13 15 0 2 3 3 13 1 9 2
6 3 13 3 0 9 2
4 3 13 9 2
11 13 15 13 9 2 13 9 7 13 9 2
23 9 3 3 13 1 9 2 10 9 13 9 0 0 9 7 13 9 9 13 1 15 9 2
16 1 12 1 0 9 0 9 9 7 9 15 13 9 0 9 2
17 9 13 3 3 13 9 1 9 7 1 9 0 9 1 0 9 2
40 9 7 9 9 13 9 7 1 0 9 9 0 2 0 9 2 1 15 15 13 2 16 4 13 3 2 7 4 3 13 0 0 9 2 13 10 0 0 9 2
48 1 12 2 0 9 0 0 9 2 15 15 13 3 9 9 1 11 2 13 3 3 1 9 10 9 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 7 0 2 1 11 2
22 10 0 0 9 13 0 9 13 12 0 9 0 9 2 1 15 15 3 7 3 13 2
17 9 9 13 2 16 1 9 10 9 15 3 13 0 9 0 9 2
30 13 15 9 0 9 9 2 1 15 7 15 2 15 15 13 0 9 7 10 9 13 13 0 9 2 15 13 1 9 2
10 3 13 3 0 13 9 1 0 9 2
14 9 1 15 0 13 3 0 9 7 13 3 3 0 2
26 13 2 14 15 2 16 9 0 9 1 9 13 0 9 16 9 9 2 4 15 13 0 9 1 9 2
16 13 3 9 2 15 3 13 9 2 9 7 0 9 1 9 2
20 10 9 15 3 13 3 13 7 13 15 0 9 7 9 1 9 1 0 9 2
11 13 1 9 4 13 13 0 16 13 9 2
11 4 7 0 9 13 9 1 9 0 9 2
11 13 0 9 7 0 9 7 9 1 9 2
25 13 1 15 13 15 7 1 0 9 2 13 3 3 12 9 2 16 0 9 1 0 9 13 9 2
14 3 3 3 13 15 13 2 16 9 7 9 9 13 2
14 0 9 2 13 15 2 16 15 10 9 13 0 9 2
16 0 0 9 15 3 2 1 0 9 2 15 13 1 0 9 2
23 3 1 10 9 13 2 7 16 15 3 13 9 2 13 4 7 3 15 1 0 9 13 2
22 7 3 12 0 9 2 1 9 2 3 4 13 1 9 9 2 15 15 9 13 0 2
9 15 10 9 13 1 0 9 9 2
4 11 11 2 11
5 0 9 7 0 9
39 3 3 15 13 2 16 0 0 9 1 11 13 9 0 9 2 15 1 0 9 2 11 7 1 9 1 11 7 11 13 1 11 3 7 3 0 0 9 2
13 1 9 4 10 9 13 9 16 2 0 9 2 2
19 3 1 9 0 9 15 11 2 11 2 11 13 13 9 2 0 9 2 2
14 3 13 1 12 9 2 15 15 13 1 9 2 12 2
17 3 1 10 9 4 0 9 3 13 14 1 9 12 9 2 12 2
15 3 15 13 1 9 1 9 2 3 15 13 16 0 9 2
13 13 3 0 11 2 11 2 11 7 9 1 11 2
35 0 3 0 9 9 0 1 9 2 12 13 12 9 2 9 12 2 7 13 2 16 9 2 12 1 11 13 10 9 2 16 13 0 9 2
18 1 10 9 13 0 9 9 3 0 1 3 0 9 7 9 0 9 2
22 3 0 0 9 13 11 1 9 12 1 11 7 12 1 11 7 1 9 12 2 12 2
10 9 2 0 9 2 15 13 1 10 9
31 2 13 15 13 9 0 9 7 10 9 2 3 13 0 2 16 0 9 15 13 1 9 9 9 7 0 1 9 0 9 2
23 2 3 0 9 13 1 10 9 3 14 0 9 0 9 7 3 13 9 9 1 0 9 2
19 2 11 2 11 2 0 9 2 0 9 2 9 12 2 12 2 12 2 2
2 11 11
3 12 2 12
4 13 4 1 9
1 11
1 11
3 0 11 2
5 12 9 9 1 9
54 1 10 9 2 16 11 11 13 9 10 9 2 16 0 0 9 3 13 0 9 11 2 13 9 9 7 10 9 2 9 9 7 9 9 0 7 0 3 16 9 9 0 9 0 0 2 16 0 2 9 9 1 9 2
14 1 0 12 9 13 9 9 13 15 1 10 9 3 2
21 0 9 7 0 9 4 13 9 0 9 7 1 9 15 13 1 9 9 1 9 2
39 4 13 0 0 9 1 15 2 16 9 9 0 13 1 0 9 0 9 9 1 9 2 7 15 0 9 1 9 0 9 2 2 7 9 9 13 3 0 2
26 1 11 2 14 12 9 1 0 11 2 15 13 0 11 2 0 9 0 1 0 9 0 9 11 11 2
11 1 9 9 15 1 0 9 13 0 9 2
35 9 13 1 12 9 12 9 0 9 9 2 15 13 9 1 9 9 1 0 12 9 2 9 9 4 13 9 1 9 9 12 7 12 2 2
36 0 9 13 0 9 2 7 1 10 9 13 0 9 0 13 14 1 12 9 1 9 0 1 9 9 0 9 7 7 13 1 9 1 0 9 2
26 11 2 11 2 11 1 0 2 11 0 9 1 11 2 1 11 2 10 9 13 9 2 2 13 13 2
15 9 1 15 13 2 16 9 0 11 13 0 2 15 13 2
26 7 9 1 15 3 13 2 16 9 1 0 0 9 7 0 9 13 3 0 2 16 4 15 13 2 2
9 7 14 1 9 13 3 3 13 2
8 11 12 2 12 2 12 2 12
8 11 12 2 12 2 12 2 12
29 9 9 0 9 1 12 2 9 0 2 9 2 2 9 0 9 1 9 0 9 7 9 0 9 9 1 0 11 2
16 2 9 1 0 11 13 13 1 0 9 2 3 1 9 2 2
20 1 9 1 0 11 13 0 9 0 3 3 3 3 16 13 9 1 0 9 2
12 9 3 13 9 2 1 15 4 13 9 9 2
12 9 3 13 0 9 9 0 1 0 9 0 2
8 0 9 4 13 1 12 9 2
31 15 13 9 2 15 4 13 1 10 9 13 9 1 9 2 1 15 9 1 9 13 1 9 9 1 9 1 9 9 9 2
12 13 15 2 16 9 1 0 11 13 0 9 2
5 9 2 9 7 11
38 9 7 9 15 13 1 15 2 16 0 0 9 9 0 2 9 9 2 9 7 9 2 15 1 11 13 14 1 12 2 9 2 1 0 9 1 11 2
41 0 9 7 13 1 0 9 1 9 0 9 9 9 10 9 1 0 9 11 2 0 11 1 11 2 2 15 10 9 13 1 9 12 2 12 2 3 1 0 9 2
26 3 9 9 2 0 4 1 11 13 1 11 2 7 1 11 13 1 9 9 2 1 12 9 9 2 2
17 10 9 1 9 11 13 2 16 4 3 13 3 2 16 15 13 2
18 13 3 13 11 2 11 11 13 11 1 9 2 12 10 2 9 2 2
6 11 12 2 12 2 12
10 0 9 7 0 9 7 13 9 13 2
40 13 15 2 16 0 3 0 9 13 1 9 9 0 9 2 7 2 9 0 3 2 0 9 7 1 0 9 10 9 2 10 9 4 3 13 9 0 9 2 2
24 9 2 16 0 0 9 13 9 9 2 13 0 2 7 9 9 16 0 9 13 0 0 9 2
24 10 9 1 9 1 0 9 0 9 13 13 0 2 9 10 9 9 4 9 13 3 3 13 2
20 0 9 13 7 13 1 0 9 16 9 2 13 9 9 1 10 9 2 2 2
8 11 12 2 12 2 12 2 12
6 9 2 9 2 9 9
15 9 0 9 13 1 9 2 16 9 9 13 0 9 0 2
13 9 2 1 15 4 9 13 2 13 7 3 0 2
23 0 9 7 13 0 9 0 9 2 7 10 9 0 1 9 9 2 2 10 9 13 4 2
20 1 10 0 9 13 3 2 0 9 2 15 15 9 15 13 1 9 7 9 2
19 1 12 0 9 2 15 15 13 1 0 9 2 15 4 3 13 3 12 2
21 9 13 9 13 15 16 1 9 3 1 3 0 9 2 16 0 9 13 3 0 2
30 13 15 2 16 0 11 3 13 12 9 0 9 2 12 9 0 9 2 1 9 1 0 9 12 9 9 0 9 2 2
17 3 15 13 2 16 9 15 13 1 0 9 9 7 1 0 3 2
14 12 1 9 0 9 2 15 13 9 13 2 13 9 2
30 1 3 16 9 9 2 15 13 1 9 9 13 2 4 9 13 3 1 12 2 1 15 12 13 0 3 1 12 9 2
15 3 13 10 12 9 12 9 1 9 0 9 1 9 9 2
7 0 11 13 12 9 3 2
25 1 9 2 15 13 9 9 3 2 13 2 16 0 0 9 4 1 9 0 1 0 9 3 13 2
16 1 9 3 3 2 13 2 16 4 9 9 13 0 0 9 2
18 9 9 13 2 16 13 0 3 13 9 2 10 9 13 9 9 9 2
24 0 9 9 0 1 9 9 1 9 2 12 1 9 2 13 13 0 7 13 13 0 0 9 2
36 1 9 0 9 15 3 2 13 2 16 9 13 7 0 9 10 9 1 9 15 13 0 7 3 13 1 9 9 9 2 15 3 9 9 13 2
8 11 12 2 12 2 12 2 12
4 0 9 7 9
5 0 9 16 0 9
24 1 9 9 1 9 0 16 12 9 13 10 0 9 2 13 0 9 7 13 15 1 0 9 2
31 10 0 9 0 9 13 9 0 9 10 9 2 7 14 12 9 10 9 2 3 3 9 9 2 7 9 0 3 9 9 2
23 3 3 12 9 15 13 2 16 3 0 9 13 9 7 13 15 2 9 3 2 13 2 2
12 1 9 9 4 3 0 9 13 16 0 9 2
20 0 9 7 13 1 0 9 2 0 9 15 13 3 16 15 3 13 1 15 2
22 10 0 9 7 3 13 1 0 9 9 0 9 2 15 4 13 1 9 0 9 2 2
11 3 0 9 13 7 3 0 1 0 9 2
9 3 12 9 1 0 7 0 9 2
10 11 12 2 12 7 12 2 12 2 12
12 0 9 9 2 9 2 13 13 9 2 12 9
26 0 9 9 13 0 9 9 2 15 15 13 1 0 9 9 2 13 3 9 12 2 12 2 12 2 2
15 3 9 9 2 15 13 1 9 9 13 3 1 9 9 2
13 0 0 9 2 15 13 0 0 9 2 13 0 2
30 4 13 9 10 9 1 9 9 2 3 9 0 9 2 7 2 9 10 9 2 15 13 9 9 0 1 0 9 9 2
41 1 10 9 13 0 0 9 2 1 9 2 16 9 9 2 12 2 3 16 9 9 2 12 2 13 9 9 1 0 9 2 13 9 9 2 12 1 0 0 9 2
29 16 3 1 9 9 4 13 13 0 9 7 9 7 9 9 9 9 2 12 4 13 13 9 1 9 10 0 9 2
8 11 12 2 12 2 12 2 12
5 13 9 9 9 2
23 15 13 9 9 2 13 3 9 2 7 0 9 10 9 13 1 12 0 9 2 0 9 2
14 9 9 4 15 13 1 9 2 9 9 3 1 9 2
39 1 0 9 7 3 12 7 12 9 13 9 2 15 13 0 9 1 9 1 10 9 0 2 13 3 11 2 11 2 9 12 2 12 2 12 2 12 2 2
14 10 9 4 13 3 2 1 9 7 10 0 0 9 2
22 0 9 11 11 1 0 0 9 13 1 0 9 2 16 10 9 13 13 0 9 9 2
25 0 9 11 11 15 10 9 13 3 1 9 2 12 7 13 2 16 0 0 9 13 9 9 9 2
8 11 12 2 12 2 12 2 12
8 11 2 9 7 9 0 0 9
24 11 13 13 9 16 9 1 0 9 1 9 1 9 2 7 13 13 1 0 9 1 9 9 2
50 1 1 15 2 16 0 9 13 0 9 1 15 9 1 0 9 2 13 9 0 0 0 11 2 15 13 0 9 1 0 9 1 9 7 9 2 2 16 11 4 13 13 10 0 0 9 1 0 9 2
13 3 15 9 13 1 0 0 9 9 1 9 0 2
8 0 9 4 13 7 3 13 2
13 9 4 3 3 13 2 16 15 13 3 0 9 2
16 9 10 9 13 3 0 9 3 1 9 2 3 1 0 9 2
28 11 13 9 2 1 15 4 10 9 13 4 13 2 16 4 4 13 1 9 0 9 9 9 1 9 7 9 2
18 15 4 0 9 13 9 0 9 2 1 9 9 7 9 3 0 9 2
8 11 12 2 12 2 12 2 12
3 9 2 9
5 7 9 9 9 2
5 15 13 15 9 2
25 3 3 13 13 15 9 3 0 0 7 0 9 1 0 9 2 15 15 9 13 13 1 10 9 2
20 16 1 0 9 13 9 13 2 0 2 0 9 13 13 0 9 7 9 9 2
15 9 13 0 9 2 0 9 15 13 13 10 0 9 9 2
3 14 15 2
32 16 0 9 13 0 7 0 2 14 1 9 9 1 9 2 2 13 9 10 9 2 0 2 2 0 2 9 9 15 13 13 2
10 12 1 9 9 15 13 9 1 9 2
41 9 3 13 0 9 2 3 15 13 13 2 7 0 9 13 2 13 2 3 13 0 0 9 2 0 9 2 0 9 3 2 16 4 15 13 2 13 0 7 0 2
13 9 9 13 9 2 15 3 9 13 1 0 9 2
18 3 13 4 9 2 9 2 13 2 13 2 13 1 9 7 9 9 2
21 3 15 1 15 13 2 16 4 15 13 9 2 16 9 7 13 10 0 9 2 2
31 9 15 13 13 9 0 0 9 0 2 0 7 0 9 2 7 2 13 13 1 9 0 2 0 15 0 2 9 2 9 2
16 9 2 9 2 2 0 9 4 13 9 9 1 9 7 9 2
18 13 7 9 0 9 2 0 9 2 2 0 9 4 13 13 1 9 2
8 9 7 9 4 13 0 9 2
6 9 16 9 4 13 2
17 9 15 13 3 0 13 1 9 9 0 9 7 0 9 10 9 2
29 10 9 15 13 9 11 2 11 2 11 2 11 11 11 2 0 9 2 0 9 2 9 2 7 0 9 1 9 2
15 11 15 13 1 0 9 16 1 9 9 2 9 0 9 2
7 9 13 13 16 9 9 2
19 11 13 1 9 7 9 2 7 9 1 9 2 7 9 9 1 9 9 2
31 0 9 1 0 0 9 4 15 13 13 1 0 9 1 9 16 15 13 1 0 0 0 9 1 0 2 0 2 0 9 2
1 3
3 9 0 9
2 11 11
47 16 9 3 13 1 9 3 3 0 9 2 1 0 9 3 9 0 9 7 9 5 9 9 2 1 3 0 3 0 9 15 1 0 9 2 2 3 14 15 3 13 1 3 0 9 9 2
21 3 1 11 2 0 9 1 9 9 2 7 1 11 2 0 9 1 9 11 2 2
12 3 3 15 1 0 9 13 1 12 0 9 2
12 9 10 0 9 9 13 7 3 3 3 0 2
22 15 3 3 13 2 16 10 9 13 3 1 9 2 7 15 14 3 2 7 7 3 2
40 13 3 7 7 10 9 2 16 13 11 2 9 11 2 2 0 1 9 2 11 2 9 11 2 2 9 1 9 2 7 11 2 9 11 2 2 0 1 9 2
24 0 13 2 16 0 9 3 3 13 9 16 9 2 7 3 15 13 16 0 0 9 0 9 2
17 7 15 14 1 9 2 7 7 1 9 0 9 7 1 0 9 2
22 3 1 9 9 1 9 0 9 13 1 9 1 0 9 7 1 9 0 9 7 9 2
27 1 9 4 13 0 9 2 1 15 1 0 13 0 11 2 15 9 13 7 9 0 12 9 1 12 9 2
42 1 2 0 2 2 3 3 0 0 9 2 3 2 11 2 13 9 0 2 0 9 9 9 1 11 1 9 2 3 2 11 2 11 2 7 3 3 2 0 2 11 2
22 1 0 9 9 9 13 0 9 2 15 15 1 10 0 9 13 2 3 11 7 11 2
14 13 1 9 0 3 1 11 2 7 15 1 0 9 2
24 0 9 13 1 9 0 9 9 0 9 1 11 1 12 2 7 12 2 9 2 3 1 11 2
27 10 14 0 9 2 7 7 3 2 0 9 2 4 1 9 13 1 0 9 2 3 9 2 9 7 9 2
13 3 1 12 2 9 4 13 9 0 9 0 9 2
12 1 9 0 9 15 7 13 3 7 0 9 2
15 3 13 10 0 9 9 3 9 9 7 0 9 1 9 2
9 0 9 13 3 0 9 9 9 2
25 7 3 0 13 3 9 1 9 2 9 1 9 9 2 0 10 0 9 1 9 9 7 0 9 2
11 7 7 1 15 3 13 9 0 0 9 2
1 9
17 1 9 7 1 0 9 15 13 3 1 9 7 9 7 1 9 2
10 3 3 9 1 0 9 13 2 13 2
10 1 9 9 15 13 7 13 9 9 2
14 1 9 9 1 9 1 0 9 15 0 9 13 9 2
27 3 9 3 13 14 9 9 1 9 2 15 4 15 13 13 1 0 2 3 14 0 2 9 2 9 2 2
37 10 9 13 3 0 9 2 9 1 9 13 9 1 9 2 3 3 15 9 13 1 9 1 0 9 7 9 15 3 13 1 0 9 1 9 0 2
24 9 7 9 13 3 9 7 9 12 9 0 9 2 0 2 3 2 0 9 2 3 0 9 2
28 3 13 13 9 3 3 2 16 1 15 0 9 0 3 9 13 9 2 1 0 9 15 13 9 7 9 2 2
23 1 1 0 9 2 3 2 9 2 13 1 9 2 9 13 3 9 2 7 10 9 13 2
16 0 9 13 3 3 0 2 3 10 2 15 13 1 0 9 2
33 3 3 9 2 1 9 9 9 0 9 1 0 9 0 9 16 9 0 9 2 1 15 15 3 16 9 13 9 7 9 0 9 2
9 10 9 15 7 13 1 10 9 2
18 1 9 3 0 9 13 0 13 9 3 0 2 15 13 3 3 13 2
17 13 15 13 2 16 1 9 15 3 13 9 2 3 9 0 9 2
17 15 15 3 3 13 2 3 1 0 9 1 0 9 9 7 9 2
17 0 0 9 13 7 15 2 1 15 15 1 0 9 13 3 9 2
28 9 9 0 9 3 13 2 16 4 15 13 1 9 3 0 2 13 15 3 9 0 9 4 14 13 0 9 2
10 15 15 13 1 9 1 9 9 9 2
22 13 15 9 3 10 2 0 2 9 2 3 2 9 2 9 2 7 9 2 15 13 2
34 1 10 0 9 15 3 13 7 1 9 0 9 2 16 13 3 9 2 3 10 9 2 7 1 0 9 15 0 9 13 1 9 0 2
25 3 0 0 9 13 0 2 9 0 2 3 3 13 12 9 0 0 9 2 7 0 15 3 9 2
6 10 9 13 3 2 9
32 16 13 9 9 0 7 9 0 2 13 15 10 9 1 9 0 9 9 12 5 7 0 9 9 12 5 7 3 1 0 9 2
20 15 4 13 2 3 15 15 13 13 2 12 9 9 9 4 3 13 1 15 2
16 13 2 0 9 4 3 13 0 7 15 15 4 13 1 0 2
23 9 10 9 13 13 2 13 2 14 12 9 9 3 0 2 1 0 9 13 13 9 2 2
41 16 9 0 9 13 9 0 9 0 1 0 9 2 3 2 1 12 9 9 2 7 1 0 0 9 2 3 2 1 12 9 9 2 2 15 15 13 1 0 9 2
52 9 9 13 3 0 2 7 7 3 0 9 13 1 0 9 1 9 2 3 9 9 9 2 2 0 13 9 2 0 9 0 9 2 7 0 9 7 9 9 2 9 1 0 9 2 3 2 1 0 9 2 2
24 0 9 0 9 1 9 11 11 11 15 3 13 0 0 9 3 1 0 9 2 7 1 9 2
8 3 13 3 0 0 9 1 9
18 9 12 5 2 9 2 5 9 2 9 2 5 9 12 5 2 9 2
11 3 9 2 9 2 13 9 1 0 9 2
34 0 1 9 9 10 9 13 9 2 16 9 1 9 13 3 2 0 2 2 7 16 13 13 0 9 9 2 15 13 0 2 0 9 2
47 10 0 9 13 13 3 2 7 2 9 10 9 13 3 2 1 9 0 9 2 15 13 0 0 9 2 16 1 9 0 9 2 12 9 15 3 13 14 9 2 7 7 9 10 0 9 2
37 9 9 7 13 2 16 4 1 15 13 14 1 9 9 9 0 1 0 9 2 14 7 1 9 9 9 2 15 15 13 2 0 2 0 9 2 2
22 1 10 9 4 7 13 9 12 9 2 1 0 9 2 0 7 9 4 13 3 13 2
13 12 0 9 7 13 9 1 9 9 7 1 15 2
19 1 10 9 15 12 0 9 13 13 1 0 9 1 2 0 2 9 9 2
20 1 10 9 13 9 9 0 2 7 0 13 3 2 16 13 3 3 0 9 2
31 9 1 9 1 0 9 0 9 7 1 9 0 9 9 15 13 9 9 2 16 13 9 9 0 1 9 7 9 0 9 2
14 3 10 9 13 9 0 9 2 15 13 9 0 9 2
24 0 9 13 3 1 9 9 2 7 7 11 13 13 9 9 1 0 0 9 7 13 10 9 2
19 13 15 9 9 3 1 0 9 2 7 15 3 9 0 2 7 9 0 2
80 1 0 9 15 11 13 1 9 0 1 9 2 3 2 1 9 9 9 9 2 15 13 3 0 9 1 0 9 0 9 2 1 9 9 1 9 12 0 9 2 13 4 0 9 2 16 3 10 9 2 15 4 15 13 1 0 9 9 2 13 1 10 9 1 11 9 2 12 1 9 0 9 2 3 15 10 9 13 2 2
9 10 9 11 3 13 1 9 9 2
21 3 9 9 9 9 1 9 3 13 0 9 2 9 13 3 3 0 1 9 9 2
35 3 10 9 9 2 11 2 11 2 9 2 11 2 11 7 9 2 11 2 11 13 2 16 0 9 9 13 9 0 9 0 1 0 9 2
31 3 13 1 0 9 9 2 7 0 9 13 1 9 7 0 9 2 9 2 2 1 15 9 13 3 3 16 1 10 9 2
10 10 9 7 3 13 1 9 0 9 2
5 3 1 0 9 2
11 13 15 12 2 9 12 1 11 1 11 2
17 13 1 0 0 11 11 2 3 3 13 9 9 1 9 2 12 2
15 1 9 12 2 12 13 9 0 11 11 1 11 1 11 2
17 0 9 13 1 9 12 1 0 11 2 3 15 13 3 0 9 2
23 3 13 1 0 0 11 1 11 2 3 15 3 13 1 9 9 0 9 1 10 0 9 2
12 1 11 13 9 2 12 1 9 0 0 9 2
2 11 11
36 3 13 13 9 9 1 0 0 11 2 1 11 2 2 12 2 12 2 12 2 2 1 15 9 9 13 9 0 9 1 9 0 9 1 11 2
25 1 10 0 9 3 13 1 10 9 16 9 2 16 15 13 9 0 9 0 1 15 2 3 13 2
17 2 14 3 3 13 3 16 9 7 3 7 12 7 3 9 2 2
27 9 13 7 3 13 9 2 15 13 0 9 1 0 9 2 3 13 0 9 2 1 15 4 9 9 13 2
42 10 9 2 15 13 1 9 2 7 3 1 9 2 13 13 9 0 9 10 9 2 16 15 3 13 3 9 2 16 3 13 0 2 9 0 9 2 1 0 9 13 2
2 11 11
3 12 2 12
5 0 9 7 0 9
51 3 15 2 15 13 1 9 7 1 9 0 7 7 0 2 13 12 0 2 13 15 1 0 9 9 7 9 2 15 1 15 3 13 2 3 15 13 2 13 7 13 2 7 15 3 13 2 13 7 13 2
12 13 15 13 9 9 2 9 9 2 9 9 2
15 13 15 13 9 9 2 9 9 2 9 9 2 9 9 2
7 7 9 9 2 9 9 2
15 13 15 13 7 0 9 9 2 9 9 2 9 0 9 2
12 9 0 0 9 2 9 0 9 2 9 0 9
34 1 0 9 0 9 2 9 2 9 7 0 0 9 3 4 13 7 13 10 0 9 2 15 4 15 13 0 9 1 0 9 0 9 2
23 13 15 7 13 9 2 16 10 9 13 13 7 16 2 16 4 13 2 13 15 10 9 2
11 7 13 2 16 1 15 7 4 3 13 2
42 14 3 13 1 10 9 0 9 2 15 3 1 0 9 9 11 11 7 10 9 13 0 9 0 13 1 9 9 16 1 0 2 0 9 10 9 2 9 7 9 2 2
55 0 9 2 16 15 0 9 0 9 13 13 1 9 0 9 9 2 7 9 2 13 13 0 9 0 0 9 2 2 2 13 2 13 13 2 13 15 2 3 2 2 7 13 2 16 4 3 0 9 9 13 1 12 9 2
29 13 2 14 15 0 9 2 3 14 15 13 2 9 3 3 15 13 2 2 7 13 1 0 3 7 0 9 9 2
52 13 15 3 2 10 9 2 13 2 14 15 9 2 3 2 0 9 9 1 0 9 10 9 2 3 0 2 3 1 9 13 0 15 2 15 13 3 3 0 9 9 2 13 2 16 10 9 13 0 9 2 2
24 3 15 15 15 4 13 16 0 9 9 1 10 0 9 2 7 3 13 2 16 9 9 9 2
28 0 9 2 3 0 9 9 1 0 9 2 2 16 3 0 2 13 3 0 2 3 16 4 13 9 0 9 2
34 9 9 1 1 9 13 3 13 16 10 0 9 9 2 0 13 3 3 7 1 15 2 3 1 15 2 3 4 15 1 9 13 9 2
16 3 0 9 1 0 9 13 9 0 9 9 2 0 0 9 2
18 1 10 9 13 1 15 3 0 9 1 11 11 2 9 2 12 2 2
51 0 9 13 0 9 2 0 2 9 2 13 3 1 0 9 0 9 10 9 2 13 15 13 14 9 7 9 2 13 15 13 2 3 15 1 9 13 2 7 0 9 2 0 9 2 0 9 7 0 9 2
25 3 15 9 9 13 1 9 9 2 13 1 0 1 15 2 10 9 13 0 9 7 9 1 9 2
24 0 9 13 2 16 0 9 2 13 2 9 14 10 10 9 7 1 15 3 13 10 0 9 2
16 1 9 1 9 3 13 13 3 3 2 1 9 3 0 9 2
12 0 9 13 3 2 0 2 9 9 12 9 2
18 13 2 14 15 3 2 16 1 0 9 1 0 2 13 9 3 0 2
22 16 4 9 1 11 9 13 0 2 13 4 7 1 0 9 9 9 1 9 1 9 2
24 3 2 16 15 1 15 15 13 7 1 9 0 2 3 4 15 15 13 1 0 0 9 2 2
14 9 9 13 9 3 0 9 9 2 15 3 3 13 2
38 13 4 3 0 9 13 0 9 1 9 2 9 9 9 2 7 10 9 2 16 3 13 9 2 15 13 9 9 2 7 15 4 13 3 14 0 9 2
20 13 3 2 16 1 9 13 3 3 0 9 9 2 0 15 13 2 0 3 2
29 13 2 14 10 0 9 16 1 9 2 3 15 1 15 13 1 3 0 9 2 2 13 15 0 0 9 3 0 2
33 9 15 3 13 13 15 2 1 15 10 9 13 13 7 3 2 10 0 0 9 13 13 3 1 0 9 2 0 9 7 0 9 2
4 11 11 2 11
7 9 2 11 11 2 9 2
23 2 2 12 2 13 9 1 0 9 0 9 1 11 7 9 1 0 2 0 9 9 0 2
11 13 15 0 9 1 0 9 9 7 9 2
15 9 2 11 11 2 2 12 2 13 0 9 11 1 11 2
21 1 9 0 7 0 9 10 9 15 13 9 0 9 9 7 9 9 7 0 9 2
18 9 2 11 11 2 2 12 2 13 0 9 1 0 9 11 1 11 2
10 1 0 9 11 15 13 9 7 9 2
7 9 2 11 11 2 9 2
10 2 2 2 13 1 0 9 9 0 2
21 1 9 1 9 7 9 1 12 2 0 9 9 0 9 1 11 15 13 3 9 2
7 9 2 11 11 2 9 2
12 2 2 12 2 13 9 1 0 9 9 0 2
10 1 0 9 11 11 15 13 9 9 2
6 9 2 11 11 9 2
16 2 2 12 2 13 1 0 9 9 0 7 1 0 0 9 2
4 13 15 9 2
28 1 0 9 13 7 9 0 0 9 2 3 2 9 7 9 2 0 9 12 2 9 9 2 0 9 12 2 2
6 13 1 0 9 11 2
9 9 2 9 2 11 11 2 9 2
12 2 2 12 2 13 0 2 0 9 9 0 2
19 1 9 0 9 7 1 9 0 9 15 13 0 0 9 7 9 0 9 2
13 10 9 13 16 0 9 1 11 1 11 2 11 2
9 9 2 9 2 11 11 2 9 2
15 2 2 12 2 13 0 9 11 7 9 1 0 9 11 2
15 13 15 9 9 9 7 0 2 0 9 0 9 0 9 2
2 0 9
2 11 11
23 0 9 0 9 13 9 9 2 16 9 13 2 10 9 2 3 2 9 2 15 3 13 2
12 1 10 0 9 13 7 1 9 0 0 9 2
10 9 0 9 15 7 13 14 1 9 2
30 1 0 9 15 13 1 9 0 9 2 1 9 9 0 9 9 7 9 9 1 9 2 1 9 9 9 2 2 2 2
13 1 9 15 1 9 9 1 9 13 0 9 9 2
11 9 4 15 0 1 9 13 9 1 0 9
15 3 3 15 15 15 13 2 9 13 3 0 7 13 15 2
23 3 15 7 13 2 13 0 7 0 9 2 16 12 9 9 10 9 1 0 15 9 13 2
21 0 9 4 9 1 9 13 3 2 7 16 13 0 13 2 16 15 13 3 3 2
11 13 15 9 13 2 16 10 9 3 13 2
15 7 13 3 9 2 16 1 15 13 0 9 16 1 9 2
17 15 9 13 3 3 3 3 13 7 13 2 16 13 15 3 3 2
52 13 2 14 2 16 9 0 9 3 0 1 9 13 0 9 0 7 13 3 3 2 13 3 0 9 9 1 9 9 0 15 9 0 9 2 3 0 2 9 2 0 9 2 2 3 4 9 13 1 9 2 2
27 13 15 3 1 9 0 9 2 13 4 14 13 9 0 9 2 15 13 1 9 2 3 15 10 9 13 2
13 3 16 1 0 9 2 15 3 3 13 9 9 2
19 9 9 3 13 1 0 0 9 2 16 15 3 3 13 0 9 0 9 2
11 13 3 1 0 9 7 1 0 0 9 2
36 14 0 9 1 12 9 2 9 9 9 7 10 9 2 13 1 9 7 9 9 1 0 0 9 9 3 2 3 15 1 9 13 10 10 9 2
9 7 15 13 1 9 13 0 9 2
14 14 16 13 1 0 9 2 3 15 13 1 0 9 2
8 0 9 13 9 9 9 9 2
23 16 9 13 2 13 14 0 9 9 2 1 3 0 9 2 1 9 1 0 1 0 9 2
14 3 1 9 15 0 9 13 1 9 0 2 9 2 2
15 13 1 0 9 10 9 2 15 1 15 13 3 0 9 2
25 0 9 12 9 2 3 9 2 13 1 0 9 9 9 2 9 15 1 0 9 13 1 0 9 2
21 1 9 9 9 1 9 13 9 9 2 1 9 9 9 1 9 13 0 1 9 2
7 3 13 1 3 0 9 2
10 1 9 12 0 9 15 15 0 13 2
18 7 2 3 3 0 9 2 9 2 13 2 3 13 1 0 9 9 2
12 13 0 2 16 9 15 13 1 0 9 9 2
20 13 4 0 13 2 16 15 9 0 3 14 12 9 13 1 9 0 7 0 2
12 1 9 9 13 1 0 0 7 3 0 9 2
19 3 1 15 13 15 9 10 9 2 16 0 9 15 13 1 0 9 9 2
23 13 15 3 3 3 7 3 13 2 3 15 9 1 0 9 0 9 13 3 0 9 9 2
15 3 13 0 13 2 16 15 1 0 9 13 3 15 0 2
14 9 13 1 9 1 0 9 7 13 15 1 9 9 2
30 13 2 14 1 9 1 0 9 9 2 7 0 0 9 2 2 13 1 9 14 9 10 10 9 2 7 7 10 9 2
19 3 13 2 13 7 1 15 2 10 0 0 9 1 10 3 0 9 13 2
24 13 0 14 2 10 9 13 9 1 0 9 2 7 7 2 10 9 1 15 13 1 9 2 2
15 13 2 14 9 1 9 12 2 9 2 13 3 12 9 2
24 1 0 9 2 9 2 13 9 9 1 0 9 0 9 3 2 16 4 0 9 13 3 0 2
12 7 3 2 9 14 3 13 1 10 0 9 2
42 1 9 0 2 7 3 3 1 9 0 2 13 9 13 3 2 10 0 9 13 0 2 7 4 13 1 3 0 9 2 2 7 1 15 13 3 3 9 0 0 9 2
20 2 13 10 9 3 13 9 1 0 9 2 7 14 12 9 3 15 13 2 2
18 3 15 15 13 13 2 16 9 0 1 12 9 2 13 9 2 2 2
12 12 1 15 13 0 7 0 7 13 9 0 2
10 0 13 0 7 0 7 13 9 0 2
18 12 2 1 0 9 13 0 9 1 9 0 7 9 15 13 14 3 2
14 1 10 9 15 13 16 9 15 13 0 9 2 9 2
20 13 2 14 15 9 2 9 15 13 3 7 2 13 3 3 9 1 9 2 2
9 7 15 9 13 0 2 0 9 2
31 13 0 9 2 1 9 13 15 2 1 0 9 2 12 9 9 2 2 1 15 12 9 13 1 0 2 13 1 0 9 2
21 0 9 1 12 9 9 2 0 2 0 7 0 2 12 2 7 9 3 13 13 2
27 3 0 9 13 13 0 9 2 0 9 2 1 9 1 9 2 9 3 2 2 13 13 1 0 0 9 2
13 1 9 1 9 9 7 9 13 9 3 1 9 2
8 13 3 1 2 0 9 2 2
10 9 3 13 0 2 9 2 0 9 2
24 9 1 0 9 2 1 15 13 1 0 9 0 9 3 16 1 9 9 2 3 13 0 9 2
35 7 0 9 2 15 13 1 0 9 7 9 3 1 9 9 0 9 2 13 1 0 9 1 9 0 1 0 2 1 0 7 1 0 9 2
27 9 0 9 3 0 9 13 0 2 9 9 1 0 9 2 15 1 0 9 9 2 9 13 1 0 9 2
24 13 1 9 0 15 0 9 2 0 15 3 1 0 9 2 2 15 13 0 9 0 9 9 2
17 15 7 13 15 10 0 9 0 1 9 9 2 1 15 4 13 2
13 9 3 13 1 3 12 9 2 0 9 1 9 2
32 9 1 0 9 0 0 9 15 13 13 16 0 9 2 15 13 13 13 14 12 0 2 3 0 9 2 13 9 2 12 2 2
28 0 9 13 9 13 15 0 9 7 7 1 0 9 13 12 9 7 9 13 0 0 9 7 1 0 0 9 2
37 1 0 9 7 2 3 16 13 15 1 9 9 2 0 9 13 10 9 3 2 16 0 9 4 13 1 9 3 3 3 2 0 9 9 13 0 2
19 1 9 12 2 1 10 12 9 13 1 0 2 0 2 0 2 9 9 2
26 3 16 1 9 0 9 13 3 1 9 9 1 9 1 0 2 0 2 9 1 9 0 2 0 2 2
9 15 15 7 13 2 0 9 2 2
16 1 0 9 4 3 3 2 1 9 2 3 15 9 13 3 2
7 3 3 13 9 3 0 2
25 13 1 9 2 12 13 1 0 9 1 0 1 9 9 3 2 16 13 14 9 0 9 0 3 2
5 13 15 15 15 2
10 3 7 3 13 1 9 9 0 3 2
16 13 2 14 15 1 15 1 9 0 3 2 13 10 9 3 2
21 0 9 15 13 13 15 2 16 13 0 9 0 14 9 12 9 7 0 0 9 2
8 7 15 3 3 13 0 9 2
17 9 9 3 13 0 9 2 1 15 1 0 9 10 9 3 13 2
27 1 9 0 16 9 13 9 1 0 9 13 3 3 2 16 7 1 12 9 9 13 0 9 0 0 9 2
40 3 2 7 16 15 9 1 9 0 0 9 3 3 13 2 13 1 9 1 0 9 2 1 15 13 0 0 9 9 2 1 9 2 1 15 13 15 9 0 2
21 7 13 15 10 9 2 15 15 13 1 3 0 9 2 9 13 7 0 7 0 2
23 9 1 9 9 7 9 2 7 3 0 9 2 13 0 2 16 4 15 1 0 9 13 2
11 1 9 15 12 13 13 16 9 9 9 2
11 9 10 9 1 10 0 9 13 1 9 2
7 9 3 13 2 9 2 2
43 13 2 14 3 9 9 1 9 2 12 16 9 2 15 13 1 9 9 0 7 1 9 12 2 9 0 2 3 13 1 15 2 1 10 9 9 4 9 0 9 9 13 2
6 15 13 14 0 9 2
15 0 9 4 3 2 13 1 9 9 0 1 9 9 9 2
24 1 0 9 2 3 15 9 3 13 1 9 2 15 3 13 14 14 12 2 12 5 0 9 2
22 1 0 9 2 3 15 13 13 14 12 5 0 9 2 4 9 13 9 0 1 9 2
14 15 13 1 15 2 10 9 13 13 1 9 0 9 2
22 7 3 1 9 15 2 15 15 13 1 9 9 9 2 13 0 9 0 9 0 9 2
32 0 9 1 0 9 13 2 13 2 14 9 16 0 9 2 3 0 9 13 3 13 1 9 9 7 13 1 9 12 2 9 2
24 13 2 14 9 9 1 0 7 0 9 9 2 13 2 16 1 9 2 9 15 9 13 0 2
9 0 9 13 0 9 0 0 9 2
10 0 9 13 3 1 0 1 0 9 2
8 3 0 9 13 13 0 9 2
19 13 15 9 13 16 0 9 1 12 0 0 9 1 15 13 13 9 9 2
24 13 2 14 3 1 9 3 3 0 9 2 13 1 10 0 9 1 9 7 9 15 13 0 2
2 12 2
11 3 2 1 0 9 13 1 0 0 9 2
32 9 9 0 9 13 1 9 9 3 0 2 15 13 9 9 2 7 0 0 9 13 0 13 3 2 16 4 13 7 10 9 2
35 3 0 9 0 9 13 2 13 2 14 15 9 9 0 9 1 9 2 7 3 2 1 1 9 9 2 1 9 2 2 15 15 13 9 2
13 9 15 2 16 9 13 1 0 9 2 13 9 2
21 2 13 1 15 2 3 3 13 9 13 2 3 13 0 2 15 13 9 3 2 2
11 1 9 9 2 9 15 9 13 3 3 2
21 13 2 14 9 2 9 2 9 13 1 15 2 16 13 2 14 2 0 9 9 2
13 3 0 9 7 13 2 13 2 14 7 9 9 2
17 0 9 9 2 9 2 1 9 9 10 9 13 9 0 12 9 2
19 2 9 2 9 2 5 12 2 13 2 14 9 9 13 2 0 2 9 2
20 2 9 2 9 2 5 12 2 12 2 13 2 14 13 9 2 15 3 13 7
19 2 9 2 9 2 5 12 2 16 9 1 9 9 3 2 3 2 13 2
18 1 9 0 9 2 3 1 12 9 2 13 0 9 9 2 9 2 2
48 2 1 0 9 2 1 15 9 2 9 2 5 12 2 4 9 2 9 2 5 12 2 12 1 9 9 2 16 15 1 10 9 9 13 1 9 9 2 9 2 5 12 2 12 2 13 2 2
16 2 16 15 1 0 9 13 2 13 9 2 9 2 5 12 2
27 2 9 2 1 15 9 2 9 2 5 12 2 12 2 13 1 9 2 9 2 5 12 2 9 13 2 7
22 2 9 2 1 15 9 2 9 2 5 12 2 13 13 2 9 2 9 2 5 12 2
53 9 10 9 2 13 13 1 9 0 2 0 0 9 2 13 0 3 13 1 9 7 3 15 13 2 16 1 9 0 16 0 9 9 15 9 1 12 0 9 4 3 13 2 16 1 9 2 9 1 0 9 13 2
12 1 1 9 9 13 13 1 9 10 0 9 2
18 3 13 13 14 1 9 0 9 2 3 0 9 1 9 13 0 9 2
11 0 9 4 13 3 7 1 9 9 9 2
14 0 9 1 10 9 4 1 10 9 13 12 9 9 2
23 13 2 14 9 9 14 1 9 0 16 9 2 13 9 14 3 2 13 2 1 9 9 2
33 7 3 0 9 2 3 1 9 9 9 9 1 9 2 3 15 15 1 9 13 1 0 11 2 13 1 0 9 1 9 9 9 2
25 1 9 10 9 1 9 9 9 1 9 13 0 13 1 9 7 9 9 9 2 3 2 9 2 2
45 15 15 13 3 2 15 2 16 7 13 9 7 1 0 9 9 2 7 9 1 9 3 3 13 2 9 2 9 2 3 13 13 9 9 9 2 7 0 9 9 1 0 9 2 2
25 0 9 4 13 9 9 1 9 2 9 2 5 12 2 0 1 9 2 9 2 5 12 5 12 2
24 9 9 2 9 2 5 12 3 13 2 16 9 9 13 13 9 2 15 9 13 7 13 0 2
30 9 13 0 13 3 2 16 1 0 9 13 9 2 9 2 5 12 3 1 9 2 9 2 5 12 2 9 15 13 2
12 7 1 15 10 9 15 0 9 13 10 9 2
30 1 9 9 9 13 14 0 9 9 9 2 3 2 7 9 9 2 9 2 2 9 9 2 1 0 9 1 9 9 2
11 7 9 9 15 1 9 13 13 0 9 2
29 9 1 9 9 0 1 9 7 2 9 2 2 2 2 13 9 9 2 9 2 5 7 2 9 2 2 2 2 2
24 9 9 3 13 15 2 3 9 9 13 10 9 1 9 1 9 0 9 7 1 0 0 9 2
38 7 3 2 7 0 9 2 3 3 2 0 9 13 10 9 3 2 16 4 13 1 0 9 1 9 1 0 9 1 10 0 9 2 13 1 0 9 2
20 9 10 9 1 0 9 0 9 1 0 9 13 3 0 2 7 3 3 0 2
21 13 2 14 1 9 2 7 1 9 13 9 9 2 1 15 13 9 9 0 9 2
13 13 1 9 0 15 1 0 9 0 7 0 9 2
7 9 9 13 13 0 9 2
15 7 1 0 9 0 9 13 0 9 2 13 2 3 3 2
15 15 3 13 1 0 9 10 9 9 1 9 1 0 9 2
10 12 2 13 3 1 14 3 0 9 2
14 9 9 13 9 15 9 2 1 15 15 10 9 13 2
13 12 2 7 12 2 13 2 14 1 9 7 9 2
34 12 2 1 9 13 2 16 16 9 13 9 0 2 0 9 0 9 2 3 13 1 0 9 0 9 2 7 3 2 1 0 0 9 2
18 12 2 13 14 1 0 9 7 13 9 2 16 4 15 15 13 13 2
5 12 2 3 13 2
11 0 4 13 13 9 0 1 9 10 9 2
35 16 13 1 9 7 0 0 9 1 0 9 2 3 9 2 13 13 0 0 9 2 10 9 13 1 15 2 1 10 9 13 0 0 9 2
3 9 1 9
9 1 15 15 13 1 9 7 1 15
3 11 1 9
34 0 0 9 2 15 13 9 2 12 13 9 11 2 15 3 13 0 9 1 9 7 9 7 3 3 13 13 1 0 9 10 0 9 2
28 3 4 1 10 9 13 2 16 0 9 2 15 13 13 9 9 0 1 0 9 2 13 2 13 15 15 13 2
28 9 0 9 15 9 11 13 9 13 15 2 16 9 13 1 9 3 2 16 4 15 9 3 13 7 3 13 2
3 7 3 2
22 3 11 13 1 9 2 15 4 13 9 13 2 13 15 1 15 1 9 2 13 2 2
13 7 1 10 9 3 2 9 7 13 1 9 13 2
31 11 13 1 9 0 9 3 0 2 0 0 9 13 7 14 0 2 0 2 9 2 13 13 1 11 3 12 9 1 9 2
15 16 3 2 1 12 9 4 13 0 13 3 12 2 12 2
17 9 1 0 9 9 7 1 9 0 9 1 9 7 9 3 13 2
24 12 2 9 15 11 13 7 15 2 16 13 9 9 1 9 0 9 2 1 0 9 1 0 2
8 13 15 9 0 9 0 9 2
5 9 11 13 12 2
30 1 12 9 11 11 1 0 0 11 1 11 13 9 9 11 7 13 2 16 13 3 13 12 0 9 2 15 15 13 2
37 1 9 15 9 2 11 13 1 0 9 0 9 2 3 3 0 11 2 1 15 15 3 3 13 2 16 15 13 1 15 13 2 13 0 9 2 2
20 9 9 11 13 0 7 14 13 0 1 9 13 1 15 9 0 16 12 9 2
19 13 15 2 16 7 10 9 13 13 12 9 1 9 12 9 7 12 9 2
20 3 15 13 7 13 15 3 3 7 13 1 0 9 3 1 12 2 12 9 2
19 13 15 14 3 2 16 14 0 0 9 13 10 9 2 13 9 2 11 2
14 13 3 2 16 1 9 0 9 15 12 9 9 13 2
11 9 13 0 0 9 2 16 13 10 9 2
14 7 9 11 2 15 13 9 11 2 13 3 0 9 2
4 11 13 13 9
15 13 4 3 1 9 0 0 9 1 9 2 0 9 11 2
16 2 0 0 9 13 9 9 0 11 11 2 3 15 13 2 2
19 13 10 9 2 16 0 9 9 13 2 16 4 13 13 10 0 9 9 2
40 9 15 13 1 9 11 11 2 9 9 14 7 14 3 1 9 1 10 0 9 2 7 7 2 16 9 9 3 13 9 9 10 0 9 1 9 9 7 9 2
23 13 3 2 16 13 1 9 0 9 1 9 2 9 1 9 2 15 13 13 9 1 9 2
8 9 0 11 11 13 3 0 2
23 0 9 1 9 9 3 13 2 16 9 4 13 0 7 0 13 1 3 0 9 7 9 2
6 9 3 13 3 3 2
13 9 3 13 2 1 10 9 13 9 1 9 13 2
22 0 9 10 9 13 2 9 1 0 9 1 11 3 13 10 0 9 1 9 1 9 2
4 9 9 9 12
8 1 9 15 13 1 9 12 2
18 13 7 1 0 0 9 7 9 9 2 16 15 15 13 0 9 9 2
27 0 9 1 0 0 9 13 9 2 3 13 9 9 9 12 2 1 15 15 9 13 1 9 9 0 9 2
22 9 10 9 15 13 13 0 7 0 9 9 15 3 13 13 3 3 3 1 0 9 2
17 0 9 4 13 2 16 4 9 13 13 1 0 9 10 0 9 2
26 9 13 3 1 9 2 3 15 9 13 13 0 9 9 9 2 16 4 1 15 13 13 1 0 9 2
3 9 1 9
18 1 10 9 4 3 13 7 1 0 9 13 0 9 1 0 9 12 2
20 1 9 9 1 9 4 15 13 1 15 2 16 12 9 13 9 7 9 9 2
9 1 9 15 10 9 3 3 13 2
22 9 9 1 9 0 0 9 13 0 9 2 9 13 4 3 13 7 3 4 13 9 2
19 9 13 2 3 13 13 0 9 1 0 9 1 0 9 9 9 1 9 2
31 9 9 3 3 13 9 2 1 15 13 3 12 5 9 2 7 3 16 12 5 2 15 13 9 1 9 1 9 12 9 2
9 1 9 13 3 9 13 9 9 2
17 9 1 0 9 15 3 13 9 9 2 9 7 9 9 2 2 2
4 7 9 13 9
28 0 0 9 1 9 9 1 9 13 9 9 2 11 11 1 0 9 9 9 9 1 9 1 9 0 0 11 2
28 16 1 12 9 15 3 1 9 13 9 9 3 3 2 3 1 10 0 9 13 9 2 11 14 12 9 3 2
25 9 9 9 13 3 1 0 9 2 9 2 9 7 15 3 1 10 2 15 13 1 3 0 11 2
16 11 15 3 3 12 9 13 0 9 2 13 2 13 2 13 2
22 15 13 13 12 9 2 1 9 15 13 2 13 1 9 9 7 13 0 9 1 9 2
10 7 15 3 13 13 7 1 0 9 2
22 9 4 15 13 13 1 9 1 9 2 9 4 13 13 1 0 9 7 9 1 9 2
10 3 10 9 13 15 9 7 1 15 2
18 7 1 9 9 13 3 1 0 9 1 9 0 15 9 9 2 2 2
5 10 9 15 3 13
39 0 0 9 13 2 16 15 9 1 0 12 9 9 12 13 1 9 2 12 1 12 9 7 1 12 9 1 9 2 12 2 15 13 0 9 1 0 9 2
25 9 13 13 3 0 9 9 0 9 2 12 9 11 11 1 0 9 7 3 7 9 9 0 11 2
21 7 0 9 13 13 14 0 9 3 0 0 9 9 9 0 9 1 0 12 9 2
5 0 9 1 0 9
26 1 9 13 12 0 9 2 11 2 11 2 11 2 11 2 11 7 11 9 1 9 0 9 1 11 2
9 9 13 13 9 1 9 7 9 2
22 9 9 13 3 1 9 7 13 4 13 13 9 2 12 2 3 1 9 0 9 9 2
12 13 4 1 0 9 3 7 3 1 0 9 2
30 9 3 0 9 13 0 9 2 1 10 9 0 3 3 9 10 9 13 0 9 13 3 1 9 2 3 1 0 9 2
13 0 9 2 13 2 0 9 0 0 9 0 9 2
17 9 13 13 0 9 1 9 2 0 9 2 9 7 9 0 9 2
18 7 15 7 3 13 9 0 9 2 15 13 3 3 13 7 10 9 2
30 7 9 1 12 2 9 12 2 10 9 1 9 0 9 13 0 13 14 1 11 2 13 0 9 1 0 9 0 11 2
4 0 9 1 9
14 0 0 9 13 13 0 9 2 13 3 1 0 11 2
11 0 9 3 13 12 5 9 1 10 9 2
20 0 7 0 0 0 9 15 13 3 3 13 0 9 1 11 2 15 13 9 2
10 3 3 13 12 5 15 0 0 9 2
21 11 2 11 3 13 2 16 4 11 13 1 11 13 15 9 2 9 7 0 9 2
19 9 9 0 0 9 15 13 16 0 2 16 10 9 13 13 1 9 9 2
7 3 13 3 3 1 9 2
18 9 9 13 2 16 1 0 9 15 9 13 3 7 3 1 0 9 2
12 13 11 1 0 0 9 4 13 10 9 9 2
9 7 1 11 7 13 15 1 9 2
8 13 13 12 9 3 1 11 2
10 1 9 9 11 13 3 3 13 9 2
14 1 11 13 9 0 9 7 0 9 3 13 1 9 2
13 3 1 15 13 9 0 9 2 15 13 3 0 2
15 1 11 11 13 3 1 10 9 1 12 9 9 2 2 2
24 13 16 0 9 13 2 16 4 0 9 13 3 7 16 4 0 9 13 1 3 3 0 9 2
16 9 3 13 0 9 3 13 1 10 2 3 3 3 0 9 2
6 11 13 12 0 9 2
22 1 15 1 9 13 1 9 9 11 2 16 9 1 15 13 0 9 15 1 7 1 2
7 1 0 9 13 7 11 2
15 9 9 0 9 13 9 9 0 0 9 1 9 2 12 2
13 11 3 13 0 9 9 2 13 15 3 0 9 2
26 9 0 0 9 1 11 13 2 11 13 10 9 7 0 9 13 1 9 2 16 4 13 0 0 9 2
10 7 15 15 13 0 9 2 0 9 2
13 1 11 3 3 12 9 13 12 5 0 9 9 2
20 9 0 9 0 9 13 3 13 9 10 0 9 2 15 4 13 1 9 9 2
13 3 13 12 2 12 9 9 9 1 9 12 9 2
13 12 1 15 13 13 13 1 11 1 11 1 9 2
16 0 9 9 11 2 0 0 2 13 13 13 1 0 0 9 2
7 0 9 1 10 9 13 2
19 9 13 3 13 12 9 1 9 12 2 12 9 7 12 1 9 3 0 2
18 13 1 9 9 0 3 1 0 9 2 15 0 9 13 1 3 0 2
34 9 13 7 12 0 9 2 1 15 12 1 11 1 11 2 3 9 13 9 2 12 2 7 4 1 12 9 3 13 1 9 0 9 2
11 1 9 0 9 13 9 9 1 0 9 2
22 13 15 2 16 4 11 13 13 3 0 9 1 0 9 2 15 4 13 4 13 3 3
5 0 0 9 9 11
13 11 11 15 3 13 10 9 1 9 9 7 9 2
38 16 9 9 11 2 11 13 0 9 7 3 2 16 4 13 0 9 2 9 0 9 1 0 9 2 0 9 15 9 13 2 13 3 1 9 0 9 2
42 11 11 3 13 16 0 9 1 0 0 0 11 1 11 2 13 7 12 9 1 11 1 11 2 13 0 9 2 7 1 9 2 12 13 16 9 0 11 1 0 11 2
25 13 3 0 10 0 0 9 2 7 9 1 9 0 9 1 9 2 9 0 9 7 0 0 9 2
44 9 15 1 10 9 13 0 9 0 9 9 1 0 9 3 2 1 2 0 9 2 2 3 0 0 9 2 0 9 0 9 2 9 9 0 3 0 9 7 9 0 0 9 2
23 9 13 2 16 10 0 9 13 3 9 2 7 9 2 16 3 12 9 13 1 0 9 2
9 0 0 9 2 9 9 7 9 2
17 11 15 13 15 15 13 2 7 15 7 1 9 10 9 7 9 2
33 0 9 11 11 2 15 13 12 9 2 13 10 9 1 9 1 15 2 16 11 13 0 9 9 3 0 0 9 7 10 0 9 2
14 1 9 13 9 9 7 9 1 0 9 1 10 9 2
4 9 3 13 2
22 15 2 15 13 1 0 9 2 1 15 2 2 7 3 13 7 13 14 1 0 9 2
19 7 1 15 2 15 3 13 1 9 0 9 0 9 2 13 3 9 9 2
22 11 2 11 2 11 13 10 0 9 16 12 1 0 9 1 0 9 1 11 2 11 2
26 0 9 15 13 1 0 9 2 0 9 1 9 15 13 13 1 10 9 2 13 13 1 9 2 2 2
6 3 15 15 3 13 2
16 13 9 0 9 3 0 0 9 2 15 15 13 13 0 9 2
14 11 13 2 16 3 3 15 13 1 0 7 0 9 2
16 16 1 11 13 1 0 0 9 0 9 0 9 2 9 13 2
24 13 2 16 11 2 11 7 11 2 11 1 9 12 2 12 13 9 9 0 0 9 9 9 2
10 3 3 13 13 9 0 9 7 9 2
17 11 2 11 7 11 2 11 10 0 9 13 0 9 9 2 2 2
28 9 2 12 13 0 9 0 9 11 2 11 1 0 9 2 16 4 4 13 9 1 0 9 2 7 1 9 2
17 9 2 12 13 15 1 10 9 11 2 11 2 11 11 2 11 2
9 0 0 9 7 13 10 9 9 2
12 7 3 3 1 11 13 9 0 9 11 11 2
25 1 0 9 13 1 9 1 0 11 7 9 2 12 4 13 1 11 1 9 1 9 0 0 9 2
26 16 13 2 16 9 4 13 1 0 9 2 9 1 9 2 13 9 9 9 11 1 0 9 1 11 2
25 9 1 11 3 13 9 2 15 13 1 3 3 0 9 2 3 13 9 11 2 3 13 10 9 2
32 1 11 2 11 15 11 13 3 1 9 10 9 13 0 9 1 9 0 9 2 15 9 15 13 1 9 11 2 11 11 11 2
18 9 13 15 0 1 11 11 2 7 13 9 9 9 2 12 9 9 2
18 9 2 12 15 13 1 9 2 15 15 3 13 0 0 9 0 9 2
9 9 2 12 3 4 13 0 9 2
9 4 13 9 1 9 7 9 9 2
11 1 11 13 3 0 0 9 1 9 11 2
11 13 3 1 11 2 9 13 7 0 9 2
13 1 11 0 9 13 0 9 3 13 1 9 9 2
18 1 11 3 2 13 1 0 9 0 9 7 0 9 0 0 0 9 2
11 1 9 7 4 13 9 9 7 9 9 2
11 13 3 13 2 16 0 9 13 3 9 2
13 10 9 13 2 16 4 1 11 13 3 0 9 2
34 3 13 3 0 13 0 0 9 2 2 1 0 9 2 15 13 0 9 11 2 11 2 13 15 13 15 0 9 3 0 2 2 2 2
17 7 11 3 13 11 2 11 2 16 4 11 3 3 13 2 2 2
12 1 0 9 4 15 13 13 1 11 3 3 2
11 9 0 9 13 11 2 11 9 2 12 2
17 9 2 12 3 4 13 2 16 13 1 15 2 3 10 9 13 2
10 3 2 16 7 10 9 13 1 11 2
21 9 2 12 15 7 1 11 13 2 16 13 1 0 9 2 16 0 9 13 0 2
17 11 13 1 0 9 1 11 7 1 9 2 16 15 13 1 11 2
13 10 9 7 9 7 13 10 9 0 9 1 11 2
16 11 4 9 2 12 13 1 12 9 7 1 9 13 1 11 2
19 9 0 9 15 3 3 13 7 9 14 13 13 1 0 0 9 0 9 2
10 16 9 13 9 0 0 9 15 13 2
20 1 11 13 9 2 16 10 9 13 9 9 9 9 1 9 1 9 0 9 2
18 11 13 2 16 1 10 0 9 15 3 0 9 13 0 13 2 2 2
29 0 9 13 13 3 3 0 0 9 7 9 11 2 11 1 0 9 11 2 11 2 11 2 11 7 11 2 11 2
25 11 11 2 15 13 1 11 2 11 1 9 2 0 9 13 2 0 9 13 3 13 9 0 9 2
27 0 9 13 1 11 11 2 0 9 10 9 2 3 15 0 1 9 13 9 3 0 2 7 0 0 9 2
23 15 9 7 9 0 0 9 4 13 2 0 7 0 9 2 2 16 0 13 3 0 9 2
8 1 11 15 3 13 0 9 2
30 16 11 13 9 9 0 9 12 2 9 12 7 13 2 3 15 2 14 2 13 9 9 2 13 9 2 16 13 13 2
19 11 13 2 16 10 9 13 1 9 7 16 11 13 13 9 1 10 9 2
20 15 15 13 0 9 2 2 0 9 13 4 13 2 16 4 15 13 15 2 2
16 9 0 0 9 13 3 1 11 2 11 2 11 7 15 15 2
28 7 0 2 0 2 9 4 1 9 0 9 13 14 14 1 0 9 2 7 1 9 0 9 13 9 3 3 2
10 9 11 9 1 11 13 13 3 0 2
5 9 0 11 13 2
30 9 0 9 11 11 13 0 9 1 9 2 15 2 2 15 4 13 13 9 1 9 12 2 12 9 7 9 12 9 2
21 0 1 15 13 15 2 16 9 13 12 9 3 1 9 2 1 15 13 0 11 2
10 0 9 13 3 0 9 9 0 9 2
31 16 1 15 13 1 12 2 9 1 11 2 9 4 3 13 13 1 10 9 2 3 15 13 9 12 2 12 9 1 11 2
10 9 9 4 13 0 9 9 10 9 2
13 3 13 10 9 0 2 3 13 0 9 0 9 2
29 9 13 3 9 3 9 11 2 3 4 3 13 13 9 13 2 3 1 9 13 0 9 11 2 0 9 2 2 2
2 11 11
12 13 1 0 9 0 9 1 11 2 9 11 11
10 3 2 9 0 2 11 11 1 0 9
13 3 2 0 9 0 2 11 11 2 9 11 2 11
26 1 9 9 9 0 2 11 1 0 9 15 9 2 12 13 7 1 9 9 7 9 0 2 11 11 2
21 13 15 9 1 0 9 0 9 9 7 9 13 7 13 0 9 1 11 1 11 2
22 13 1 9 0 9 1 9 0 9 2 15 14 13 13 0 0 9 7 13 0 9 2
33 13 15 3 2 16 9 0 13 14 0 9 0 9 2 0 15 3 1 0 2 7 16 1 15 13 7 9 3 0 2 13 11 2
16 13 2 16 7 10 9 13 2 7 13 2 16 1 9 0 2
16 0 9 9 0 13 1 11 7 0 9 15 2 15 13 3 2
30 2 2 2 9 9 13 0 0 9 1 9 11 2 16 15 13 3 15 2 15 13 2 16 9 13 3 13 9 0 2
31 1 9 2 1 15 15 0 0 11 9 11 1 11 13 2 13 3 2 2 2 9 0 9 2 0 7 3 0 2 2 2
21 2 11 9 2 12 9 1 9 1 0 2 11 11 2 9 9 2 11 12 2 2
32 0 9 7 9 1 9 1 9 0 9 11 1 11 13 3 1 9 0 2 0 9 0 0 9 10 9 0 9 7 0 9 2
41 9 7 9 11 12 2 13 10 9 2 0 9 11 12 2 2 12 2 12 2 2 3 0 9 2 13 15 0 9 7 1 0 9 9 15 13 0 9 7 9 2
13 12 1 10 9 13 7 0 0 9 11 1 11 2
18 13 1 9 0 9 2 15 13 9 2 12 1 0 9 9 11 12 2
20 13 9 0 9 2 13 13 0 9 9 2 13 9 0 9 7 13 10 9 2
7 10 0 9 13 0 9 2
8 13 9 1 0 7 0 9 2
14 9 11 1 11 7 13 0 7 10 9 15 13 3 2
20 1 9 9 2 12 15 13 1 0 9 0 9 2 0 0 9 11 1 11 2
25 10 9 1 12 9 13 9 9 0 7 1 9 0 13 10 9 13 1 9 0 9 1 0 9 2
9 1 9 11 2 11 1 9 2 12
12 0 9 1 0 0 9 0 9 1 9 0 11
4 11 2 11 2
17 9 1 0 9 1 9 1 0 9 2 0 13 0 0 0 9 2
15 9 2 3 15 1 9 12 7 12 13 11 2 0 9 2
12 1 10 9 4 3 12 2 9 12 13 9 11
17 0 9 1 0 0 9 2 15 15 13 1 9 1 0 9 11 2
4 9 11 2 11
6 12 2 12 13 1 9
2 11 2
6 9 1 2 9 9 2
27 0 12 9 3 1 11 1 9 12 9 1 2 9 2 15 1 0 0 9 13 14 12 9 0 0 9 2
15 1 10 9 15 13 9 9 1 9 0 12 9 12 9 2
19 10 0 9 2 15 13 1 9 9 2 13 1 12 1 0 0 9 9 2
23 13 15 3 3 3 12 9 2 16 15 11 11 13 1 0 0 9 1 0 9 1 11 2
15 13 15 3 12 9 2 13 9 9 7 13 10 0 9 2
12 3 13 1 0 9 0 0 9 0 0 9 2
8 13 9 0 9 1 9 9 2
22 9 13 14 9 2 12 2 3 15 1 0 9 1 11 13 11 9 11 2 9 9 2
22 3 13 0 9 1 10 9 2 3 15 9 13 13 15 15 7 14 13 9 0 9 2
16 0 12 9 0 9 13 1 0 9 1 9 12 9 12 9 2
15 1 10 9 13 0 13 10 9 0 9 1 9 12 9 2
12 9 13 0 9 0 1 0 0 9 1 9 2
18 9 9 13 13 0 0 9 2 15 13 9 3 0 9 1 9 9 2
13 9 9 7 13 12 2 12 9 0 9 0 9 2
17 11 13 0 9 10 9 2 15 15 13 13 15 9 1 9 9 2
19 0 9 13 1 9 9 1 0 9 9 2 7 4 13 3 0 0 9 2
21 3 1 10 9 13 7 9 2 7 3 3 0 0 9 2 15 13 0 9 9 2
10 15 13 7 3 0 9 1 0 9 2
32 9 10 9 13 1 9 0 9 0 0 9 2 16 9 9 2 0 3 0 0 9 2 10 13 0 7 0 9 2 13 9 2
51 1 9 1 9 0 9 15 13 2 16 15 13 13 1 0 9 0 9 2 3 3 15 13 1 9 0 9 2 0 9 0 9 2 9 7 0 9 2 0 0 11 11 2 9 12 2 11 2 11 2 2
2 11 11
23 9 1 9 9 1 9 11 2 15 4 9 2 12 13 0 0 0 0 9 11 1 9 9
9 1 11 13 1 12 9 0 9 2
37 1 9 1 9 12 7 9 12 13 1 0 9 9 0 9 2 1 9 14 12 9 2 9 11 1 9 12 9 2 0 1 12 9 1 0 9 2
2 9 2
3 11 2 11
8 9 1 9 2 9 2 0 2
4 11 1 11 2
6 9 1 9 11 2 11
10 9 0 2 11 11 1 0 0 9 2
4 9 11 2 11
1 12
20 3 3 9 9 1 0 0 9 1 9 9 9 7 9 1 0 9 0 9 2
10 10 9 13 9 0 9 1 9 0 2
9 11 1 11 7 13 1 10 9 2
2 9 2
3 11 2 11
1 12
13 9 0 9 1 0 9 16 9 2 9 2 0 2
4 9 11 2 11
2 9 9
7 0 9 13 9 10 9 2
14 0 9 13 3 13 1 9 0 9 7 1 9 9 2
8 3 13 13 7 0 9 0 2
13 1 0 9 0 9 0 9 13 0 9 0 9 2
8 3 0 9 4 13 9 9 2
11 0 9 13 9 7 15 13 1 0 9 2
12 1 9 13 13 1 9 9 0 9 1 9 2
38 9 9 13 9 9 0 9 12 7 12 2 15 13 10 9 0 9 2 0 0 9 1 9 0 9 7 0 9 0 9 2 9 2 9 3 2 2 2
16 3 13 9 2 3 1 9 1 9 4 13 9 11 1 11 2
6 3 3 13 0 13 2
22 0 9 0 9 0 9 1 9 0 1 0 9 13 13 1 9 9 9 0 1 9 2
32 1 0 9 13 10 9 13 1 9 1 0 7 0 9 1 0 9 2 0 1 9 0 1 0 9 1 9 1 0 2 9 2
9 3 3 2 9 1 0 9 1 9
10 3 3 2 0 9 1 9 1 9 2
5 0 9 13 0 9
15 3 3 2 0 0 9 1 9 9 11 2 5 12 2 2
4 9 1 9 9
8 2 9 2 0 2 11 1 11
31 9 13 9 4 1 12 2 9 13 1 10 9 1 9 9 1 9 1 9 12 5 12 9 7 1 9 12 7 12 9 2
20 4 13 0 9 0 7 3 3 0 9 2 13 0 2 3 0 2 0 9 2
12 4 13 9 9 2 9 9 7 9 9 9 2
17 1 0 0 9 13 3 1 0 9 0 9 2 0 0 9 9 2
16 1 9 13 1 9 12 0 9 9 2 9 0 9 0 9 2
10 9 4 3 3 13 9 7 0 9 2
36 1 9 15 1 3 3 0 9 13 0 7 3 0 9 2 15 13 1 0 9 9 2 16 1 0 9 13 0 9 13 1 0 9 0 9 2
13 1 0 9 9 15 13 1 0 7 0 9 9 2
11 0 7 0 9 13 2 16 2 9 0 2
8 11 11 2 13 3 0 9 2
31 9 0 0 9 13 10 3 0 9 2 13 7 0 7 1 0 9 1 0 9 4 13 0 9 2 0 9 7 0 9 2
30 9 13 0 0 0 9 2 15 13 13 1 0 7 0 9 1 9 9 1 9 9 9 11 7 9 1 12 2 9 2
35 10 9 13 0 9 1 0 9 9 2 15 7 13 0 9 0 9 2 0 1 9 0 9 9 2 7 15 13 1 9 9 0 1 9 2
10 10 0 0 9 13 0 9 9 0 2
12 9 9 13 1 10 9 7 1 9 10 9 2
19 16 1 9 9 11 1 11 13 1 9 14 10 0 9 1 0 9 0 2
14 7 10 9 13 13 1 9 9 0 9 0 1 9 2
17 0 9 13 9 9 2 15 15 1 9 13 1 9 0 9 0 2
20 1 9 9 9 2 12 13 10 0 9 3 0 7 0 2 1 9 0 9 2
19 7 1 9 1 0 9 13 2 3 13 9 1 0 9 9 9 2 12 2
18 9 0 0 9 13 1 9 10 0 0 9 7 7 1 0 9 9 2
3 12 2 12
7 11 11 2 9 9 2 12
9 9 2 9 2 12 9 12 9 2
4 13 1 0 9
4 0 9 1 11
3 9 11 11
16 11 11 2 9 2 12 2 9 2 9 2 12 9 12 9 2
16 13 1 0 9 0 9 0 9 1 11 1 11 2 9 11 11
18 9 9 9 0 9 1 9 1 9 1 9 9 9 2 9 1 9 2
14 9 13 13 1 9 9 1 9 2 9 5 12 2 2
1 12
2 12 2
7 9 0 0 9 1 9 2
12 3 4 13 1 12 9 1 9 14 12 9 2
21 0 9 9 1 9 13 13 0 9 2 3 0 0 9 0 9 7 0 9 9 2
20 9 9 4 3 1 0 9 3 13 9 9 9 2 9 2 9 7 0 9 2
11 3 15 3 13 13 0 9 1 9 9 2
1 12
2 12 2
40 9 0 9 2 3 2 1 0 9 0 9 1 12 2 9 12 15 10 9 3 13 1 9 1 10 9 2 1 15 4 13 9 12 0 0 9 0 15 9 2
11 0 9 10 9 13 3 1 12 9 0 2
1 12
2 12 2
9 2 0 0 9 2 1 0 9 2
20 3 13 13 9 2 15 15 9 9 13 1 9 7 3 15 1 15 13 13 2
19 1 3 0 9 4 13 9 1 9 12 2 0 0 9 2 0 9 2 2
11 3 13 3 13 9 0 9 1 9 9 2
26 9 0 9 9 15 13 9 9 9 7 15 13 0 9 2 15 9 9 2 13 9 2 9 9 9 2
12 9 10 9 1 0 9 9 9 3 9 13 2
1 12
4 9 11 2 11
1 12
8 0 1 9 9 2 9 2 12
1 12
4 9 11 2 11
1 12
16 9 9 9 1 9 0 9 1 9 12 7 12 2 11 2 9
1 12
4 9 11 2 11
3 13 15 2
11 15 13 13 9 7 13 15 1 0 9 2
5 13 9 2 13 2
21 13 2 3 3 13 11 11 2 11 2 16 15 15 13 13 1 9 3 9 2 2
1 12
37 9 9 0 9 12 1 0 9 7 1 9 9 12 9 2 0 9 9 1 9 1 0 9 2 11 2 7 9 9 1 12 2 9 9 2 9 2
9 0 0 9 13 3 9 0 9 2
9 9 1 15 13 9 1 0 9 0
1 12
7 0 9 11 11 7 0 11
1 12
3 9 11 11
1 12
20 9 1 0 9 15 13 13 16 0 9 2 15 13 4 13 14 12 3 0 9
1 12
1 12
3 9 0 2
9 11 1 11 1 9 9 7 9 2
4 9 11 2 11
1 12
7 0 9 9 1 0 9 2
28 13 10 3 0 9 2 13 7 0 2 13 0 0 9 2 3 0 9 7 0 9 2 15 13 0 0 9 2
11 3 1 9 12 7 2 3 12 12 7 2
4 9 11 2 11
1 12
3 9 11 11
1 12
22 2 16 0 9 15 13 13 2 16 15 3 9 13 2 16 3 13 9 9 9 2 2
3 9 11 11
15 9 0 11 2 1 15 4 3 13 0 9 9 0 9 2
7 9 13 9 9 0 9 2
12 0 0 9 13 0 9 9 1 0 9 0 2
12 0 9 13 0 7 0 9 0 9 0 9 2
15 0 9 13 13 9 2 1 15 3 13 1 9 15 9 2
14 0 9 13 3 13 9 2 3 1 9 9 3 13 2
1 9
6 11 2 11 2 11 2
2 11 2
15 11 2 11 7 9 2 2 11 12 2 12 2 12 2 12
1 12
23 11 11 2 12 2 2 2 12 2 2 2 13 1 9 2 9 2 9 3 1 12 9 2
1 12
5 0 9 1 0 9
4 9 0 0 9
10 2 0 9 1 9 2 12 2 9 2
2 11 11
76 1 0 15 3 7 15 4 13 1 9 2 16 13 2 14 9 9 7 13 2 14 1 15 9 9 9 9 2 3 13 9 9 2 7 3 7 1 9 2 16 13 2 14 9 9 9 9 7 13 2 14 9 9 2 3 13 7 9 9 2 7 9 9 2 16 4 13 0 9 2 16 15 13 15 0 2
16 13 9 10 9 0 1 9 9 2 15 13 0 1 9 9 2
7 9 9 13 1 12 9 2
22 0 1 15 13 0 9 9 0 1 10 9 2 10 9 1 9 9 3 13 9 9 2
20 0 9 13 0 9 9 0 1 10 9 2 10 9 1 9 9 13 9 9 2
32 13 2 14 9 9 1 0 1 10 9 7 13 2 14 9 9 1 9 9 2 3 3 7 9 9 13 1 0 1 10 9 2
33 3 13 2 14 9 9 1 0 1 10 9 7 13 2 14 9 9 1 9 9 2 3 3 7 9 9 13 1 0 1 10 9 2
13 9 9 9 1 10 12 9 13 3 3 10 9 2
16 13 9 9 1 15 1 10 9 13 2 13 9 2 12 2 2
7 9 9 3 13 9 9 2
42 16 4 15 3 13 1 10 9 9 2 3 3 9 9 2 3 9 9 13 1 9 9 1 9 9 2 13 9 9 2 7 3 7 9 9 1 10 10 0 9 9 2
33 7 0 9 9 9 13 1 0 3 0 9 2 1 15 4 13 9 9 2 7 3 9 9 9 13 13 9 9 2 15 13 9 2
24 1 15 9 2 15 13 9 9 7 13 9 9 2 13 3 9 9 0 9 1 9 9 9 2
10 9 9 13 9 9 9 1 9 9 2
19 0 9 9 9 1 9 9 13 3 9 0 1 9 9 1 9 9 9 2
22 9 1 9 9 1 9 9 1 9 9 13 9 9 9 9 1 9 9 1 9 9 2
11 9 9 13 9 9 9 9 1 9 9 2
7 3 10 9 13 3 0 2
3 9 12 2
16 13 9 9 9 1 9 9 2 13 9 9 0 1 9 9 2
27 3 9 9 13 9 9 9 1 9 9 7 10 9 9 1 9 9 13 1 9 9 15 16 1 9 9 2
2 9 2
16 13 9 2 9 9 9 0 1 9 9 2 9 1 9 9 2
31 13 9 9 9 9 1 9 9 2 10 9 9 13 1 9 9 1 10 9 0 9 9 16 9 9 9 9 1 9 9 2
10 13 2 16 9 9 2 9 13 0 2
45 1 9 9 13 9 9 0 1 9 9 3 2 16 4 9 1 9 9 1 9 9 13 1 10 9 0 9 9 16 9 1 9 9 1 9 9 2 13 9 2 12 2 12 2 2
29 9 9 13 1 9 9 9 9 0 2 16 13 9 9 9 9 1 9 9 2 7 13 3 9 9 1 9 9 2
17 3 13 0 2 16 9 9 13 9 9 9 9 2 15 13 9 2
32 16 4 13 10 9 2 13 3 13 2 1 10 10 9 13 9 9 9 9 9 7 1 10 9 13 13 9 9 1 9 9 2
3 9 12 2
34 2 9 2 13 9 2 9 0 9 2 13 9 9 0 9 9 1 9 9 7 9 9 1 9 9 2 3 9 2 9 13 0 9 2
24 14 9 0 9 2 15 13 9 9 2 9 1 9 9 1 10 12 9 13 0 12 9 0 2
10 3 13 13 0 9 9 9 2 9 2
9 2 9 2 13 9 9 9 9 2
11 3 9 9 2 9 13 13 10 0 9 2
2 9 2
51 2 9 2 13 9 9 9 2 9 2 13 9 9 2 15 13 9 9 0 1 9 9 1 9 9 2 13 9 9 0 1 9 9 1 0 9 9 9 16 9 9 2 16 9 9 2 9 13 3 0 2
16 16 9 9 2 9 13 3 0 2 13 9 9 2 9 0 2
9 9 9 13 3 0 1 9 9 2
20 16 3 9 9 2 9 13 3 0 2 13 9 9 2 9 2 9 1 9 2
17 9 9 13 3 0 9 9 9 2 9 2 13 9 2 12 2 2
23 2 9 2 13 9 9 0 1 9 9 2 13 9 9 9 0 1 9 9 1 9 9 2
10 14 9 9 13 0 1 9 9 9 2
31 16 9 13 9 9 9 2 13 10 9 7 1 9 9 2 7 3 9 9 9 9 1 9 9 13 0 2 15 13 9 2
25 9 9 9 1 9 9 13 9 9 9 9 2 3 9 13 9 9 0 1 9 9 1 9 9 2
36 1 15 9 0 1 9 9 13 9 9 0 9 1 9 9 2 15 3 13 2 13 2 14 15 2 16 1 0 9 13 9 0 16 10 9 2
23 15 13 3 0 9 9 2 1 15 1 9 1 0 9 13 0 9 2 15 13 0 9 2
12 14 9 9 1 9 9 13 0 16 9 9 2
24 13 9 9 1 9 9 10 2 16 9 9 13 3 0 16 9 9 2 13 9 2 12 2 2
16 9 9 13 0 2 7 3 9 9 13 3 0 16 9 9 2
24 9 9 13 0 16 9 9 7 1 9 12 1 0 9 1 9 13 9 9 0 16 9 9 2
3 9 12 2
6 13 9 9 9 9 2
11 13 9 2 9 0 9 0 1 9 9 2
17 14 9 1 9 9 1 9 9 13 9 9 9 9 1 9 9 2
13 3 9 9 13 1 9 9 0 9 16 9 9 2
2 9 2
16 13 9 2 9 9 9 0 1 9 9 2 9 1 9 9 2
11 13 2 16 9 9 13 0 16 9 9 2
25 13 9 9 1 9 9 10 2 16 9 9 13 3 0 16 9 9 2 13 2 9 2 12 2 2
33 3 9 13 11 9 7 1 9 1 9 10 9 13 9 9 0 1 9 9 2 3 9 13 9 9 9 7 9 13 9 9 9 2
15 1 9 12 1 0 9 0 9 9 9 3 13 9 9 2
35 13 2 14 9 9 0 1 9 9 2 3 9 9 13 1 9 9 9 0 9 2 16 13 9 9 9 9 1 9 9 2 15 13 9 2
33 13 2 14 9 5 9 2 3 9 9 13 1 9 9 7 9 9 13 0 9 9 9 2 9 2 15 13 1 9 1 9 12 2
30 13 4 3 2 16 4 2 14 15 9 9 13 1 9 9 9 9 1 9 9 2 4 15 10 9 1 9 9 13 2
19 4 2 14 15 7 13 1 0 9 2 4 15 10 9 1 9 9 13 2
48 3 13 13 2 16 13 2 14 3 10 9 2 13 15 0 2 3 4 2 14 15 9 9 13 1 9 9 9 9 1 9 9 1 9 2 10 9 1 9 9 3 13 1 10 3 0 9 2
39 3 13 13 2 16 13 2 14 3 10 9 2 3 4 2 14 15 9 9 13 1 10 9 1 9 1 9 0 2 10 9 1 9 9 3 13 10 9 2
35 10 9 7 3 13 4 2 15 13 9 2 16 4 15 13 2 16 13 3 0 13 9 0 9 1 10 0 9 2 16 3 0 9 13 2
3 9 12 2
16 14 9 9 13 1 9 9 0 9 16 9 9 1 9 9 2
6 14 10 9 13 0 2
20 3 9 9 9 9 1 9 9 13 3 0 16 9 9 9 9 1 9 9 2
8 9 13 3 1 9 0 9 2
3 9 12 2
16 14 9 9 13 1 9 9 0 9 16 9 9 1 9 9 2
6 14 10 9 13 0 2
19 3 9 9 9 9 1 9 9 13 0 16 9 9 9 9 1 9 9 2
2 9 2
38 1 0 9 13 3 13 2 16 9 9 2 9 13 0 7 16 9 9 13 0 9 9 9 9 2 3 9 13 9 9 0 1 9 9 1 9 9 2
15 13 9 9 9 9 0 9 9 2 13 9 2 12 2 2
23 13 9 9 0 1 10 9 0 9 9 9 2 1 15 13 9 9 9 9 1 9 9 2
15 14 9 9 13 3 0 16 9 9 9 9 1 9 9 2
29 9 9 2 9 13 1 9 9 1 12 10 9 0 9 2 10 9 13 0 12 9 0 2 7 7 15 3 13 2
10 1 9 12 9 9 13 9 9 9 2
17 13 9 9 0 1 9 9 10 2 16 9 9 13 9 9 9 2
12 9 9 13 9 9 2 7 3 7 9 9 2
30 15 13 2 16 9 9 9 0 9 9 13 1 9 9 9 9 3 10 16 9 9 2 7 3 0 16 9 9 9 2
3 9 12 2
7 14 9 13 9 9 9 2
7 3 9 13 9 9 9 2
2 9 2
20 13 9 9 0 1 9 9 2 13 9 9 9 0 1 9 9 1 9 9 2
39 13 2 16 9 9 13 9 9 9 0 9 9 2 7 3 1 9 2 15 13 1 10 9 0 9 9 9 16 9 9 9 9 1 9 9 1 9 9 2
7 13 2 16 15 3 13 2
37 3 13 1 10 9 13 9 9 10 2 16 9 9 13 1 9 1 9 9 1 9 9 9 9 9 7 9 9 13 0 2 13 9 2 12 2 2
13 13 9 9 9 0 1 9 9 1 9 9 9 2
10 3 9 9 13 0 9 9 9 9 2
34 1 9 12 13 9 9 9 9 1 9 9 0 16 9 9 9 9 1 9 9 2 7 7 9 9 2 9 15 13 1 10 9 9 2
27 9 9 9 13 9 9 9 13 7 13 9 9 2 7 9 9 13 1 9 9 2 15 13 1 9 9 2
22 15 7 13 2 16 9 9 9 13 9 6 2 7 3 7 9 9 2 15 13 9 2
24 13 2 14 3 2 16 9 9 2 9 13 9 2 3 3 13 0 13 2 15 13 9 15 2
3 9 12 2
22 13 9 2 9 2 9 0 9 7 14 9 9 13 1 10 9 9 9 9 2 9 2
8 3 9 9 2 9 13 9 2
2 9 2
17 14 3 9 9 13 1 9 9 2 9 2 13 9 2 12 2 2
20 13 9 9 0 1 9 9 2 13 9 9 9 0 1 9 9 1 9 9 2
25 13 9 9 9 9 0 9 9 2 10 9 9 13 1 10 9 0 9 9 16 9 9 9 9 2
7 14 9 2 9 13 0 2
19 3 7 9 9 13 9 9 1 10 9 9 2 7 9 13 9 9 9 2
22 16 9 9 13 9 9 9 1 9 9 2 13 9 9 3 9 9 2 15 13 9 2
18 14 3 3 9 9 13 1 9 9 2 9 2 13 9 2 12 2 2
29 13 9 9 0 1 9 9 2 13 9 9 9 0 1 9 9 1 9 9 2 13 9 9 9 9 1 9 9 2
8 9 9 2 9 15 3 13 2
44 16 4 15 3 13 1 10 9 9 2 3 4 10 9 13 13 1 10 9 0 9 9 2 1 15 13 9 9 9 9 2 7 9 13 0 9 9 1 9 9 16 9 9 2
35 16 7 9 13 9 9 9 1 9 9 2 13 4 9 9 13 9 9 2 7 1 9 9 13 1 9 1 9 9 9 0 16 9 9 2
11 14 9 13 0 9 9 9 0 9 9 2
10 13 2 16 9 9 2 9 13 0 2
17 16 9 9 13 9 9 9 1 9 9 2 13 9 9 9 9 2
12 1 9 15 13 7 9 9 2 15 13 9 2
17 9 9 2 9 2 15 15 3 13 7 13 9 2 15 13 9 2
22 9 9 2 15 13 1 9 9 2 13 3 13 3 12 9 9 9 7 3 10 9 2
18 0 9 0 9 13 1 11 11 2 7 13 15 3 0 9 10 9 2
3 9 12 2
6 13 9 2 9 9 2
13 3 13 13 9 2 15 13 0 1 12 10 9 2
2 9 2
22 13 9 2 9 2 9 0 9 0 1 9 9 10 2 16 9 9 13 1 9 9 2
20 13 9 2 9 2 9 9 9 0 1 9 9 2 9 2 9 1 9 9 2
35 13 2 14 9 9 2 9 3 0 2 13 9 11 9 7 1 9 1 9 10 9 13 9 9 9 9 2 9 0 1 9 9 2 9 2
12 14 3 3 9 9 13 0 9 16 9 9 2
24 13 9 9 0 1 9 9 10 2 16 9 9 2 9 13 0 9 2 13 9 2 12 2 2
30 13 9 9 10 2 16 9 9 13 3 0 16 9 9 2 3 9 13 9 0 1 10 9 0 9 9 16 9 9 2
27 13 9 9 9 9 2 16 9 9 10 9 13 9 1 9 9 1 9 9 7 1 9 9 1 9 9 2
27 13 9 10 9 2 16 9 9 2 9 13 3 0 7 9 9 13 1 10 9 0 9 9 16 9 9 2
10 1 9 12 13 9 9 2 9 9 2
50 9 9 2 9 15 13 1 10 9 9 2 7 1 0 9 4 9 9 9 0 9 9 13 1 9 9 0 9 16 9 9 2 15 13 3 10 9 2 15 1 9 9 13 9 9 9 0 9 9 2
16 13 9 9 0 1 10 9 9 9 0 9 9 16 9 9 2
9 14 9 9 2 9 13 0 9 2
16 13 9 2 9 9 9 0 1 9 9 2 9 1 9 9 2
22 3 13 3 0 2 9 11 2 9 13 0 2 7 3 9 11 2 9 13 0 9 2
27 3 13 2 16 9 9 13 11 9 2 7 3 9 0 9 9 9 2 9 13 0 1 9 9 2 9 2
31 13 15 2 16 10 12 0 9 13 13 12 0 0 9 2 7 4 15 13 9 2 1 15 13 9 9 0 12 9 0 2
36 1 0 9 13 2 16 12 0 15 9 9 2 9 13 9 3 3 2 16 13 10 0 9 2 7 9 3 3 2 16 13 3 12 0 9 2
3 9 12 2
6 13 9 2 9 9 2
27 13 9 9 2 9 9 0 3 1 9 9 2 9 10 2 16 9 9 13 0 1 12 9 9 2 9 2
18 13 9 2 9 9 0 1 9 9 2 16 9 9 13 1 9 9 2
13 3 9 9 13 0 9 1 9 9 16 9 9 2
2 9 2
22 13 9 2 9 9 9 0 1 9 9 2 9 1 9 9 2 13 9 2 12 2 2
26 16 9 9 1 9 13 0 16 12 9 0 2 13 9 9 0 2 7 1 9 15 9 9 13 0 2
34 16 4 9 12 2 9 13 0 9 2 13 4 9 11 9 2 7 3 9 9 9 9 2 9 4 13 0 0 9 9 9 2 9 2
12 14 3 9 9 9 13 0 9 16 9 9 2
19 13 9 9 0 1 9 9 9 10 2 16 9 9 2 9 13 3 0 2
18 3 9 13 11 9 2 7 3 1 9 1 11 9 13 9 9 0 2
27 1 9 12 1 9 1 9 13 9 9 0 16 9 9 2 7 3 7 9 9 13 0 2 15 13 9 2
35 4 2 14 15 3 9 9 13 1 12 1 12 9 1 10 0 9 2 16 3 1 12 7 0 9 2 4 15 10 9 1 0 9 13 2
33 3 1 10 9 13 13 2 16 4 2 14 15 13 1 9 2 3 16 3 13 10 9 2 3 10 9 1 0 9 10 9 13 2
29 3 9 0 9 2 15 1 10 9 13 2 13 1 11 2 7 14 3 7 2 16 4 15 13 0 9 0 9 2
8 1 0 9 13 3 0 9 2
3 9 12 2
23 13 9 9 2 9 9 2 15 1 15 13 2 9 9 9 0 1 9 9 1 9 9 2
26 13 9 9 0 1 9 9 2 0 1 10 9 0 9 9 16 9 9 2 7 14 9 9 13 0 2
12 13 9 9 0 1 9 9 1 9 9 9 2
16 13 9 2 9 9 9 0 1 9 9 2 9 1 9 9 2
21 13 9 9 9 9 0 9 9 2 16 9 1 9 9 1 9 9 13 9 9 2
11 14 9 9 9 13 9 9 6 2 9 2
16 3 9 9 13 9 9 6 2 9 2 13 9 2 12 2 2
2 9 2
12 13 9 9 0 1 9 7 1 9 9 9 2
7 3 9 13 9 9 6 2
22 13 9 2 9 9 9 6 1 9 1 9 9 1 9 9 2 0 9 9 2 9 2
11 14 3 12 1 15 13 0 1 9 9 2
24 13 9 9 9 0 1 9 9 1 9 6 2 13 9 9 9 0 1 9 9 1 9 9 2
17 16 3 9 9 13 9 9 9 2 9 13 9 11 2 9 0 2
14 1 9 15 9 9 2 9 13 1 9 9 0 9 2
9 1 9 12 13 9 2 9 9 2
12 1 9 12 13 15 7 9 2 15 13 9 2
21 9 9 2 9 13 3 0 1 9 9 2 1 9 15 13 9 9 9 9 6 2
11 3 13 2 16 9 9 13 9 9 9 2
3 9 12 2
4 13 0 9 2
21 3 13 13 9 9 7 9 9 10 2 16 9 9 9 9 1 9 9 13 9 2
2 9 2
31 13 9 2 9 2 9 0 9 10 2 16 9 6 2 9 13 3 0 7 9 9 13 9 12 2 13 9 2 12 2 2
17 13 9 9 9 9 1 9 1 9 9 1 9 9 0 9 9 2
13 13 9 9 0 1 9 7 1 9 9 9 9 2
14 3 9 13 9 9 6 1 9 9 9 1 9 9 2
23 13 9 9 2 15 13 9 9 7 13 10 9 9 6 2 7 2 1 15 13 9 9 2
11 13 9 9 0 1 9 9 1 9 9 2
11 3 9 9 13 0 9 9 9 2 9 2
32 9 9 2 9 13 1 10 9 9 6 2 1 15 13 9 9 2 1 9 6 0 9 2 10 9 13 0 16 12 9 0 2
37 3 3 13 2 16 9 9 2 9 13 1 10 9 9 9 2 1 15 13 9 9 2 1 9 9 0 9 2 10 9 13 0 16 12 0 9 2
23 16 15 3 9 9 2 9 13 2 3 1 10 9 0 9 9 2 1 15 13 9 9 2
22 16 9 9 2 9 13 9 2 3 10 9 9 13 1 9 9 2 9 1 10 9 2
17 16 9 9 2 9 13 9 2 3 10 0 9 13 1 10 9 2
10 13 2 16 9 9 2 9 13 9 2
39 16 15 4 13 2 3 0 9 9 13 10 0 9 2 7 1 0 9 13 10 9 9 9 6 2 9 2 7 3 9 9 9 9 1 10 9 13 9 2
17 13 2 3 3 2 16 9 9 2 9 15 13 1 10 9 9 2
16 3 9 9 13 1 9 9 7 9 11 2 9 13 0 9 2
19 13 9 9 9 6 1 9 1 9 9 1 9 9 2 15 13 9 9 2
11 1 9 12 13 3 9 9 2 9 9 2
66 16 9 2 15 13 9 9 1 9 9 6 0 9 9 2 1 15 13 9 9 2 7 9 2 15 13 9 9 1 9 9 9 0 9 9 7 10 9 9 1 9 6 2 13 0 9 2 13 9 9 9 9 1 9 6 3 0 16 9 9 9 9 1 9 9 2
32 1 9 15 13 9 9 9 0 9 9 7 9 9 1 9 6 2 9 3 0 9 3 1 9 9 2 3 7 1 9 9 2
13 0 1 10 9 13 7 3 0 2 15 13 9 2
11 13 3 2 16 9 9 2 9 13 9 2
8 13 9 9 9 9 2 9 2
13 10 9 15 13 2 7 9 6 13 9 9 9 2
28 9 9 13 1 9 9 2 7 1 0 9 4 13 7 1 9 9 2 15 13 1 9 9 0 1 9 9 2
9 9 9 2 9 4 15 3 13 2
16 13 7 2 16 9 14 2 9 13 3 0 2 15 13 9 2
25 14 3 9 2 13 9 0 1 9 9 2 0 1 9 9 7 9 14 2 9 2 13 3 0 2
11 13 9 2 9 9 9 0 9 9 2 2
44 9 2 15 13 9 9 2 1 9 9 0 9 9 7 9 9 1 9 9 2 13 3 0 16 9 2 15 13 9 14 1 9 9 9 0 9 9 7 9 9 1 9 6 2
33 1 9 15 13 9 9 2 9 9 0 9 9 2 13 1 9 9 2 9 3 0 9 16 9 9 9 0 9 9 1 9 9 2
23 0 1 10 9 13 7 3 0 16 9 2 15 13 9 9 9 0 9 9 1 9 9 2
24 9 9 2 2 9 3 13 1 9 9 1 12 9 0 9 2 10 9 13 0 12 9 0 2
11 1 9 12 13 9 9 2 2 9 9 2
14 9 9 13 7 10 0 9 2 7 3 1 10 9 2
11 1 9 12 13 3 9 2 2 9 9 2
30 13 2 14 15 10 0 9 3 0 9 2 9 15 13 1 0 1 15 2 15 4 14 3 1 10 0 0 9 13 2
23 3 3 16 13 3 0 9 2 3 3 1 10 9 13 13 9 2 15 3 13 10 9 2
42 13 3 13 9 0 1 9 10 9 1 9 1 9 2 15 13 3 0 2 7 0 16 9 9 9 1 9 9 2 10 9 9 1 9 9 13 0 9 10 0 9 2
43 13 2 14 0 0 9 1 3 0 9 2 3 9 10 9 13 3 13 9 9 2 3 9 13 9 9 9 1 9 9 2 10 9 9 1 10 9 13 0 9 9 0 2
38 13 2 14 12 0 9 9 2 9 0 15 1 9 9 7 13 3 1 0 9 1 9 9 9 0 1 10 9 2 4 3 13 9 1 3 0 9 2
28 16 7 10 9 13 3 0 9 9 2 13 9 10 9 1 9 2 7 3 10 2 0 2 9 15 3 13 2
2 0 9
16 1 9 1 9 11 13 4 1 0 9 13 11 11 2 11 2
27 10 9 4 7 3 13 9 9 7 13 1 15 9 9 2 15 13 0 1 0 7 0 9 3 0 9 2
29 13 7 1 9 10 0 0 9 10 9 2 1 15 4 13 13 2 16 13 3 0 1 15 2 15 3 13 11 2
19 13 15 7 0 9 2 15 11 13 2 16 15 13 3 13 13 1 9 2
11 10 9 13 9 1 9 9 7 9 9 2
44 4 15 13 9 10 9 1 9 9 7 9 9 2 15 15 13 11 2 7 3 15 13 1 15 2 15 4 3 13 9 2 7 1 10 9 4 15 1 0 9 13 15 0 2
11 3 0 9 12 7 12 10 9 3 13 2
28 13 2 14 10 9 9 2 3 10 9 13 9 9 9 9 9 1 9 9 2 1 15 13 9 9 9 9 2
13 3 0 9 9 13 1 10 9 3 12 0 9 2
20 1 9 12 3 13 2 16 3 3 2 0 9 0 9 13 3 12 9 9 2
23 4 2 14 1 0 13 1 9 1 9 9 7 9 9 2 4 13 1 9 9 3 0 2
14 9 10 9 2 16 3 9 0 7 3 2 13 0 2
16 15 13 2 16 15 13 9 2 3 4 13 1 0 9 9 2
23 1 0 9 15 13 9 0 2 7 9 0 9 2 9 0 9 7 3 2 13 9 0 2
32 13 2 14 0 9 2 1 15 4 13 0 9 2 3 15 15 14 13 3 13 10 9 2 7 0 9 15 15 3 13 13 2
26 1 10 0 0 9 13 7 0 7 10 9 9 2 3 15 2 15 1 3 0 9 13 0 9 9 2
51 15 13 7 0 13 3 2 16 16 4 15 15 1 0 0 9 13 10 9 2 7 14 0 9 2 3 16 15 3 0 7 0 2 3 15 15 13 10 9 2 3 4 1 15 7 10 9 9 13 0 2
25 16 4 0 9 13 0 1 9 10 0 0 9 2 3 4 1 15 13 3 0 9 1 0 9 2
50 13 4 1 15 3 13 10 0 9 2 7 3 4 13 13 13 15 1 10 9 2 7 7 16 4 13 15 0 9 2 15 13 10 9 2 13 4 15 3 13 2 3 16 13 3 3 13 0 9 2
27 1 0 7 0 9 1 10 0 0 9 13 13 3 10 9 2 15 1 3 0 9 13 9 9 0 9 2
9 10 9 4 13 9 10 0 9 2
24 1 0 9 13 0 2 16 9 13 0 1 15 9 9 2 15 13 13 9 10 0 0 9 2
48 13 15 3 0 9 10 2 16 13 2 14 12 3 0 9 9 2 9 0 15 1 9 9 2 3 9 0 1 10 9 1 9 9 3 1 9 9 2 9 15 13 2 13 9 2 12 2 2
35 9 2 0 1 9 1 9 9 7 9 9 2 15 13 0 11 2 11 2 11 2 15 15 3 1 9 12 13 1 0 9 10 0 9 2
55 13 1 9 3 2 16 13 0 2 16 4 0 9 13 1 9 0 0 9 2 1 9 15 13 0 2 16 4 3 1 10 9 13 0 13 0 0 9 2 15 9 13 10 9 2 7 1 10 0 9 15 3 0 13 2
25 15 15 7 13 0 9 15 2 3 3 13 1 9 0 9 1 3 3 15 1 9 0 0 9 2
7 9 1 9 0 9 0 9
48 13 2 14 15 15 13 10 0 0 9 1 0 9 2 15 15 13 2 14 1 15 13 9 2 15 4 15 13 13 15 15 16 0 1 9 2 13 3 3 9 13 15 1 9 9 0 9 2
15 10 9 7 13 7 2 16 4 13 0 9 1 9 0 2
39 1 10 9 13 2 7 13 3 10 9 1 0 9 13 1 9 0 2 7 14 3 2 16 15 1 0 9 13 2 16 3 10 7 15 9 13 7 13 2
30 16 0 0 9 2 15 15 13 9 2 15 4 13 13 2 13 9 2 13 15 3 13 2 15 13 9 1 0 9 2
18 0 9 1 0 9 7 9 0 15 13 1 9 1 0 9 0 9 2
28 16 4 15 13 9 2 1 15 13 2 4 7 15 13 0 9 16 9 2 16 10 9 4 3 13 1 0 2
13 13 2 14 1 3 0 9 2 3 13 0 9 2
26 9 10 0 9 13 13 3 0 2 16 9 10 9 15 13 1 9 0 0 9 9 9 1 0 9 2
31 3 3 10 9 13 13 0 16 12 9 2 7 13 9 2 16 4 13 13 0 0 9 2 10 9 13 0 16 12 9 2
18 16 4 15 1 15 13 2 13 13 9 0 0 9 0 1 9 12 2
27 3 10 9 13 13 0 16 12 9 2 7 9 0 0 9 1 9 0 16 12 9 15 3 4 13 9 2
22 7 14 15 2 1 10 0 9 13 13 10 9 3 0 16 9 9 2 3 13 11 2
50 3 2 16 4 10 9 13 0 3 9 9 2 3 13 1 9 2 13 4 9 9 2 0 1 9 9 7 0 13 15 1 12 9 2 13 1 12 9 3 1 9 7 13 4 13 1 12 9 3 2
15 0 12 9 4 13 0 1 9 2 13 9 2 12 2 2
14 3 13 2 1 0 9 4 13 3 12 9 10 9 2
9 1 9 7 13 3 9 10 9 2
25 3 0 9 4 3 13 9 10 0 9 14 3 1 0 9 2 7 13 15 3 15 15 3 13 2
26 7 7 10 9 4 1 15 13 13 9 2 16 9 2 1 15 4 15 13 2 15 13 1 0 9 2
8 13 4 3 13 3 0 9 2
13 13 15 2 16 9 13 10 0 9 2 3 15 2
17 13 9 9 7 9 9 2 15 15 1 15 13 1 9 0 9 2
19 1 9 9 0 9 9 7 9 9 13 9 9 9 9 2 9 9 9 2
9 3 9 9 2 9 13 3 0 2
41 13 15 3 1 9 9 1 9 0 1 10 9 1 9 9 3 3 2 16 4 1 10 9 13 9 9 7 9 9 2 9 2 9 3 13 2 16 1 9 2 2
16 3 16 3 1 9 13 0 13 0 9 1 9 11 7 11 2
17 9 9 9 2 9 15 15 4 7 1 10 9 13 16 9 0 2
29 1 10 9 7 3 3 13 9 9 2 9 3 2 16 4 13 9 9 2 7 9 9 15 15 13 13 1 9 2
14 10 9 13 7 0 7 9 9 1 15 0 13 0 2
20 16 4 15 3 3 13 13 0 9 16 9 2 3 15 13 10 9 13 3 2
16 7 9 0 1 10 9 13 3 13 9 9 10 0 0 9 2
21 13 4 10 9 13 1 9 2 16 4 13 1 10 9 13 9 0 9 0 9 2
30 16 4 13 9 9 7 9 9 2 9 2 9 1 15 16 1 9 2 13 15 13 1 9 9 1 9 0 16 9 2
50 15 7 13 2 16 9 9 13 3 10 9 0 1 10 9 2 15 13 1 0 9 2 15 0 9 13 1 9 1 9 9 9 3 0 16 9 9 9 2 1 15 15 13 10 9 2 1 9 9 2
27 13 2 14 15 1 9 2 15 13 1 10 9 2 3 15 1 9 9 13 2 7 10 9 9 9 13 2
10 0 9 9 15 15 3 13 16 9 2
13 15 13 1 10 9 2 15 3 1 9 9 13 2
14 15 0 9 9 2 9 13 9 9 1 9 10 9 2
33 15 2 15 13 1 10 9 2 13 14 0 9 2 7 9 0 10 9 1 10 2 9 2 9 9 13 2 13 9 2 12 2 2
16 0 7 13 2 16 1 10 9 4 13 0 13 0 0 9 2
25 9 0 9 3 13 13 9 0 0 9 2 7 15 4 13 9 2 16 0 9 13 0 0 9 2
24 16 4 10 9 13 0 2 13 4 13 1 9 9 2 16 0 9 13 9 10 0 0 9 2
31 9 9 1 0 9 2 7 1 9 9 0 2 15 3 13 1 9 2 16 10 2 9 2 9 13 0 9 1 10 9 2
45 1 9 9 10 0 0 9 1 3 0 7 0 9 13 13 3 10 9 13 3 0 7 0 9 2 7 13 15 13 7 9 10 9 13 3 7 9 9 2 7 9 15 0 9 2
20 9 0 9 9 9 13 3 3 3 3 13 1 9 0 15 9 9 1 9 2
60 13 2 14 2 16 9 9 1 10 9 2 10 9 9 7 9 9 4 13 2 15 13 1 12 9 0 1 10 9 2 15 13 0 16 0 9 9 2 15 4 15 1 10 9 13 13 2 3 3 3 13 13 2 3 3 13 13 9 0 2
23 9 2 15 15 13 13 2 4 3 13 2 7 0 9 3 4 13 9 10 10 9 13 2
20 16 7 9 9 2 7 9 9 3 3 13 2 4 13 3 1 10 9 13 2
30 0 9 2 3 4 13 3 3 2 16 4 13 1 0 9 13 2 16 1 10 9 13 9 9 0 3 12 9 0 2
23 3 3 3 13 7 9 2 7 7 15 13 13 10 9 3 2 15 4 3 0 9 13 2
12 1 9 1 15 13 3 1 9 13 3 3 2
13 9 1 9 10 0 0 9 9 0 3 3 13 2
73 16 4 3 13 9 13 3 3 9 0 9 7 9 2 16 4 15 13 3 0 9 0 9 2 13 15 15 13 9 0 0 9 3 13 1 3 0 7 0 9 2 7 3 13 13 15 2 16 15 0 9 13 1 9 3 0 2 7 1 10 9 15 13 10 9 2 15 4 13 13 9 9 2
20 3 9 2 15 4 13 2 13 0 2 7 13 1 9 2 13 13 0 9 2
30 9 9 9 1 0 9 3 13 10 0 0 9 2 7 13 13 2 16 4 15 15 10 9 13 13 13 0 0 9 2
40 1 15 4 13 3 2 16 4 1 9 9 1 10 9 13 2 16 9 10 9 1 12 9 0 13 0 16 0 9 9 2 15 4 15 1 10 9 13 13 2
28 1 10 9 4 3 9 9 1 10 9 13 0 12 9 0 2 15 13 1 9 1 9 0 1 0 0 9 2
16 9 10 9 13 11 1 9 9 1 9 11 2 11 2 11 2
20 9 9 9 1 12 0 2 15 1 10 9 13 2 13 7 1 9 0 9 2
13 7 10 0 9 13 0 9 0 9 1 9 0 2
25 3 14 1 9 0 9 2 7 15 9 3 15 9 13 2 7 1 9 9 2 1 15 4 13 2
56 15 0 9 4 13 1 9 7 2 16 4 13 9 2 15 4 3 3 13 0 0 9 2 7 13 3 9 10 9 1 9 2 7 16 4 13 9 2 15 13 0 1 0 9 0 9 13 1 9 2 3 14 13 1 9 2
47 1 15 0 9 4 13 9 1 3 3 0 9 0 0 9 2 7 3 4 13 7 2 16 4 10 9 13 2 15 15 1 15 3 13 13 2 7 16 4 13 2 16 10 9 13 0 2
47 9 2 16 4 13 3 0 9 13 0 0 9 2 15 13 1 9 1 15 2 16 9 2 16 1 0 9 13 9 9 1 9 0 12 9 0 2 4 3 13 1 9 9 0 0 9 2
33 0 9 2 16 4 1 10 9 13 13 13 9 15 2 15 4 1 9 13 1 9 0 2 7 1 15 13 1 15 9 0 9 2
9 1 15 10 4 13 13 7 13 2
13 13 4 15 1 15 0 9 2 14 7 0 9 2
47 16 4 13 7 3 13 1 9 2 16 0 9 13 0 1 9 0 2 15 15 13 13 0 9 16 9 1 0 9 2 3 1 10 9 4 13 0 9 13 2 7 1 15 3 13 0 2
49 1 15 9 2 16 1 0 9 13 9 9 1 9 0 12 9 0 2 15 15 3 13 1 9 0 9 16 9 2 15 3 13 0 0 9 3 13 2 7 7 15 13 13 1 0 9 10 9 2
21 10 9 4 13 9 1 0 0 9 2 7 0 9 4 15 3 13 0 9 13 2
28 9 4 15 13 3 1 9 2 16 0 9 13 0 1 0 0 9 7 16 3 9 10 9 4 15 13 9 2
42 3 7 0 9 4 15 1 0 9 13 1 9 0 9 2 7 16 4 15 13 14 0 9 0 9 7 13 3 0 9 1 9 2 3 4 15 0 9 13 0 9 2
24 3 13 2 9 1 0 0 7 0 9 13 9 1 10 9 2 14 7 9 1 15 1 15 2
25 10 9 13 13 9 2 1 15 4 10 9 13 2 3 9 0 9 16 9 0 1 0 0 9 2
8 15 1 10 9 7 13 13 2
26 16 4 15 10 9 13 2 3 4 7 0 0 9 13 13 10 0 9 1 0 9 10 0 0 9 2
12 3 3 15 7 13 7 1 10 0 0 9 2
31 10 9 1 9 10 9 7 9 0 2 1 15 3 13 3 7 9 2 3 4 15 13 13 2 13 13 10 0 0 9 2
11 9 13 0 0 9 9 0 3 13 3 2
22 9 2 15 15 4 13 2 7 13 9 2 15 15 13 9 0 9 1 0 0 9 2
14 3 2 3 13 9 2 16 9 10 9 13 1 9 2
