2837 11
70 9 9 9 1 12 9 2 0 4 13 4 16 4 16 9 1 9 1 9 1 13 16 4 9 9 9 9 1 9 1 13 4 9 2 9 1 9 1 13 9 0 12 12 12 9 1 9 9 1 2 3 9 9 1 9 1 9 9 1 9 1 13 4 9 1 0 4 13 4 2
32 9 1 13 9 9 9 1 9 1 1 9 9 14 1 9 1 12 12 12 12 2 9 1 1 12 12 12 9 1 1 13 2
42 9 11 9 1 9 9 1 9 1 13 4 14 2 9 1 9 1 13 16 9 1 9 1 13 16 2 15 14 9 1 9 9 1 15 1 13 4 16 4 4 4 2
22 9 1 9 1 0 9 1 13 9 2 9 9 9 9 9 9 1 13 4 16 4 2
8 9 1 9 9 9 1 13 2
42 11 1 1 9 9 2 9 9 9 2 9 9 2 9 2 9 1 9 2 9 9 1 9 9 14 1 9 1 13 2 9 9 1 3 12 12 12 9 1 13 4 2
54 9 9 1 2 9 1 9 1 13 9 2 9 2 9 2 9 1 9 1 0 9 1 13 2 9 9 9 9 1 9 9 7 9 9 2 9 12 9 9 1 9 9 1 9 9 9 1 9 1 13 16 13 4 2
34 11 1 9 9 1 9 9 1 13 16 13 4 2 12 12 12 12 9 9 1 9 1 11 1 9 12 12 12 9 9 1 13 4 2
30 9 9 1 13 16 1 2 15 14 11 9 1 9 14 1 13 4 4 16 4 4 16 2 9 9 1 13 4 4 2
48 9 1 1 2 3 9 9 4 9 9 9 1 9 9 1 9 9 1 12 12 9 1 12 12 12 12 9 1 13 1 13 4 16 4 16 2 9 9 1 13 4 4 9 1 3 0 4 2
26 9 1 9 9 1 9 12 9 1 9 1 0 4 2 9 1 13 16 9 1 9 1 13 4 4 2
26 11 1 1 9 9 2 11 9 1 9 2 9 9 1 12 12 12 12 12 9 1 9 1 13 4 2
30 9 9 1 9 9 1 0 13 4 16 4 16 2 9 1 9 1 13 4 16 4 4 9 9 1 0 16 1 9 2
17 11 1 9 9 1 9 1 9 1 13 16 13 4 16 4 4 2
78 9 1 13 4 11 9 1 2 9 1 0 9 1 13 4 4 9 1 9 9 1 9 2 9 1 9 7 9 1 0 4 13 2 9 9 14 4 4 2 9 9 7 9 9 1 9 9 4 9 9 1 13 16 13 4 4 2 1 13 4 2 9 1 12 9 9 1 9 9 1 13 9 1 13 4 16 4 2
30 9 7 9 9 14 2 9 1 9 9 1 9 1 13 16 2 9 2 9 2 9 14 1 9 1 13 4 0 9 2
29 13 9 1 9 1 13 4 9 9 7 2 9 1 9 1 9 1 13 4 9 1 13 4 9 9 1 9 9 2
32 12 12 12 12 9 1 3 13 2 9 1 1 9 14 4 4 9 2 9 14 14 9 1 13 4 4 9 1 13 16 4 2
17 9 9 1 9 12 9 1 12 12 12 9 1 1 9 1 0 2
38 11 9 1 12 9 2 9 1 9 11 9 1 13 16 4 4 11 9 9 1 9 1 2 9 4 9 1 9 1 13 4 16 4 1 13 4 4 2
14 7 2 11 9 1 9 9 1 13 16 4 1 13 2
25 7 2 9 1 9 1 9 4 16 14 2 9 9 1 13 4 9 9 4 16 14 1 0 4 2
46 9 9 1 13 16 2 11 9 9 1 9 9 1 12 9 9 2 11 1 11 9 9 9 1 13 2 9 1 9 1 13 16 11 9 1 13 9 1 13 9 1 13 4 1 13 2
27 11 9 9 1 12 9 2 2 11 9 1 9 0 1 12 9 1 9 1 13 4 2 1 13 4 4 2
44 12 9 9 12 12 9 12 9 9 2 11 9 11 9 11 12 2 9 11 5 11 11 9 1 11 9 1 9 12 12 9 2 0 9 12 12 9 1 13 16 9 1 13 2
43 9 9 1 13 4 9 1 13 16 2 11 9 11 9 1 2 9 9 1 9 2 1 12 9 9 14 11 9 1 12 9 2 9 12 9 1 13 4 4 1 13 4 2
29 9 11 9 14 1 13 4 4 16 2 9 9 2 9 1 10 9 1 9 1 13 2 12 9 1 9 1 9 2
18 12 9 1 9 1 9 9 1 9 1 9 11 1 9 9 4 4 2
29 9 9 1 1 2 9 9 9 9 14 9 12 12 9 1 13 4 4 16 2 9 12 9 2 9 1 13 4 2
10 12 9 9 1 9 1 13 4 9 2
17 11 9 9 1 12 9 1 14 9 13 2 12 9 1 9 9 2
29 2 9 9 1 9 2 1 9 1 12 9 9 2 9 9 1 12 9 13 2 12 9 1 13 4 9 4 4 2
44 10 9 2 9 12 9 9 9 9 1 9 1 12 9 1 13 4 16 1 13 4 9 2 11 9 9 2 11 9 14 13 4 16 2 12 9 1 13 4 16 4 4 4 2
29 7 2 9 1 12 9 1 9 1 9 9 1 13 4 4 4 16 1 2 9 11 1 9 9 1 13 4 4 2
12 9 1 9 1 9 12 5 12 12 12 9 2
30 12 9 1 9 9 1 9 12 12 12 9 1 9 1 12 12 9 9 0 2 9 1 9 9 1 13 16 4 4 2
36 11 1 11 9 1 12 9 2 12 9 9 12 9 1 13 16 2 9 1 9 11 1 1 9 1 13 4 4 13 9 9 1 13 4 4 2
83 9 1 11 11 9 9 9 5 9 1 12 9 2 11 9 1 13 2 9 1 9 9 1 13 16 2 9 7 9 1 13 4 16 4 12 12 12 9 9 1 1 9 1 9 9 1 13 4 4 4 2 9 9 1 9 2 9 1 13 4 2 1 13 2 9 9 1 1 0 9 9 1 13 4 4 4 1 1 9 1 13 4 2
38 7 2 9 1 13 16 2 11 1 12 12 9 9 1 1 13 2 9 13 4 16 2 9 1 13 16 4 2 1 13 2 9 9 1 13 4 4 2
39 11 11 9 1 12 9 1 9 9 1 9 1 9 3 13 4 16 2 9 1 9 9 14 1 9 1 13 2 9 9 1 3 0 4 9 1 13 4 2
47 2 12 9 1 1 9 1 13 9 1 13 4 2 4 4 16 2 9 1 9 9 9 9 1 1 9 1 9 9 2 3 13 4 16 4 4 9 1 9 9 1 13 4 4 9 4 2
15 9 9 1 9 1 12 12 9 1 3 13 9 1 13 2
31 11 11 9 9 9 1 2 0 4 9 4 1 4 2 1 13 2 9 9 14 1 1 13 4 4 9 1 13 4 4 2
45 9 1 12 9 1 9 1 9 9 14 1 9 1 13 16 4 16 2 9 1 13 9 1 13 9 1 9 9 13 16 4 2 9 1 13 16 1 10 9 1 13 4 1 13 2
21 9 1 9 9 1 12 12 12 12 9 1 11 11 9 9 2 9 1 9 9 2
35 9 9 1 12 12 9 1 11 11 9 9 4 16 2 10 9 1 9 9 1 9 1 9 9 1 9 1 0 1 13 4 16 4 4 2
15 2 9 1 9 1 2 9 1 9 9 3 2 1 13 2
70 9 1 11 11 9 9 1 12 9 2 11 5 11 1 9 9 1 13 4 4 9 9 9 1 13 4 2 9 9 7 9 1 9 9 1 13 16 2 3 9 4 4 9 1 9 1 9 1 13 4 14 4 2 12 9 9 2 9 9 4 9 1 13 4 2 1 13 4 4 2
18 7 2 11 9 1 9 1 9 1 0 4 13 16 4 2 1 13 2
25 2 9 1 13 4 9 2 1 1 9 1 13 4 4 4 9 1 9 9 9 9 9 9 9 2
21 7 9 9 9 1 2 9 1 9 4 13 2 1 13 9 1 3 12 12 9 2
41 2 9 1 0 9 1 13 2 2 0 9 1 13 2 2 9 1 1 9 1 13 2 14 9 1 13 4 1 13 16 4 9 1 9 12 12 9 1 13 4 2
21 9 9 4 1 2 9 4 13 2 1 9 1 3 0 16 1 9 1 12 9 2
13 9 4 0 4 4 16 1 9 1 12 12 9 2
21 7 9 9 9 1 13 16 4 16 2 9 9 1 0 9 9 1 12 12 9 2
36 9 1 9 9 9 2 0 2 9 9 9 2 1 13 4 9 7 9 1 2 3 0 9 1 13 16 4 1 13 0 4 9 1 13 4 2
24 11 2 9 1 2 9 1 1 9 1 13 2 1 1 9 1 9 12 12 2 12 12 9 2
24 10 9 1 13 9 2 9 4 9 9 1 13 16 4 4 16 14 3 14 2 9 1 13 2
39 9 1 12 9 1 9 13 1 13 2 11 11 9 9 9 1 13 9 9 9 9 1 13 2 2 9 9 9 9 2 9 1 13 9 9 1 13 4 2
55 9 12 12 9 1 9 9 9 9 1 0 1 9 9 1 9 1 13 2 9 9 9 2 1 12 2 12 1 9 1 9 1 13 2 9 9 14 1 9 1 13 9 1 13 16 4 2 9 9 1 0 9 1 13 2
17 11 11 9 9 1 12 9 2 11 11 9 1 1 9 1 13 2
66 9 1 9 9 9 1 13 16 2 11 11 9 1 0 9 1 13 9 1 9 1 0 2 7 2 9 1 13 2 9 1 9 1 13 16 9 1 0 13 16 1 0 4 2 13 4 3 13 4 4 16 2 0 9 1 13 16 4 2 1 1 9 1 13 4 2
10 9 1 13 4 16 13 4 16 4 2
24 11 1 1 9 1 13 9 1 1 4 16 2 12 12 9 9 1 9 1 9 1 13 4 2
9 15 1 13 4 4 4 9 4 2
15 7 9 1 13 4 1 13 1 1 0 9 1 9 4 2
40 9 2 13 4 4 9 7 9 1 9 12 9 1 2 9 1 0 9 2 9 1 0 9 1 13 9 14 1 1 13 4 4 4 2 1 13 16 4 4 2
28 12 12 12 12 9 1 3 12 9 1 13 16 4 4 11 1 4 4 9 9 1 9 9 1 13 16 4 2
29 11 1 1 9 9 1 0 13 4 4 16 2 3 9 1 9 1 13 4 9 1 9 1 9 1 13 4 4 2
16 11 1 1 9 1 0 9 1 13 4 9 1 13 16 4 2
20 9 9 9 9 1 1 9 9 4 12 12 9 9 13 4 4 16 4 4 2
12 9 2 9 9 2 9 14 1 1 0 4 2
22 9 9 1 12 12 9 9 13 16 2 10 9 9 1 13 16 4 4 16 4 4 2
6 9 1 9 1 13 2
5 9 12 12 9 2
9 9 9 1 13 4 16 4 4 2
18 7 2 9 9 2 1 2 9 14 1 1 13 4 4 16 4 4 2
10 11 1 13 4 16 4 4 9 4 2
12 9 9 1 1 2 9 9 7 9 9 4 2
17 9 9 9 9 1 9 9 1 15 14 1 9 1 13 14 4 2
27 0 9 1 13 16 4 16 2 10 9 1 9 1 9 1 9 9 2 9 9 1 13 16 4 4 16 2
30 9 1 13 16 4 9 1 1 2 0 9 9 1 13 4 16 2 0 0 9 1 9 1 13 16 9 9 1 13 2
8 11 1 1 15 1 3 0 2
6 9 9 1 0 4 2
13 15 1 9 9 1 9 14 13 4 0 1 13 2
21 11 9 9 1 2 11 9 9 9 2 13 4 4 16 1 12 12 9 9 4 2
8 7 9 9 13 16 0 4 2
20 9 13 9 13 4 9 1 2 9 1 9 1 13 4 0 13 14 3 14 2
20 7 2 9 9 9 9 1 9 9 1 9 9 1 9 4 13 14 13 4 2
6 3 13 4 0 4 2
18 9 9 1 9 1 13 0 9 1 2 3 13 4 9 1 0 4 2
51 9 9 1 9 14 1 2 9 1 0 4 13 9 1 13 16 2 9 9 9 1 12 9 1 13 9 2 9 9 9 1 13 14 1 13 9 1 2 9 2 9 9 7 9 1 9 1 9 1 13 2
23 15 1 3 13 4 4 2 3 9 1 13 2 9 1 13 16 4 16 1 0 9 4 2
14 9 9 9 1 9 9 1 13 9 1 0 9 4 2
31 3 13 4 9 1 9 13 1 13 9 1 1 4 16 2 9 9 9 9 1 13 9 1 3 13 4 16 4 4 4 2
41 3 9 9 9 1 1 13 4 16 2 9 1 13 4 9 1 13 16 4 4 9 1 13 16 4 1 4 2 13 9 1 13 16 1 4 16 4 1 4 14 2
26 7 9 9 9 1 1 3 0 9 1 13 16 1 2 15 1 9 9 1 13 4 1 13 4 4 2
11 0 9 1 12 12 9 9 1 3 13 2
21 9 9 1 9 1 13 16 1 2 3 13 4 3 0 4 9 1 1 13 4 2
18 9 9 9 9 9 9 9 1 13 16 1 9 1 1 0 1 13 2
26 9 9 1 9 1 9 9 0 4 4 9 9 1 13 16 4 9 1 0 16 4 1 4 14 14 2
15 10 9 1 13 9 9 1 13 16 9 9 1 0 4 2
22 11 9 1 9 9 1 13 4 4 9 2 9 1 9 9 1 13 9 1 13 4 2
7 9 1 9 1 13 4 2
19 9 9 1 1 0 9 9 1 13 4 16 2 9 1 9 1 1 4 2
10 9 9 1 13 4 9 1 0 4 2
17 9 9 1 9 1 9 1 13 9 1 13 4 16 1 4 4 2
25 9 9 1 9 1 13 16 0 1 13 16 0 1 13 16 2 0 13 0 9 1 9 1 0 2
20 15 1 9 9 9 1 13 4 4 16 1 9 9 1 9 1 13 4 16 2
9 15 1 9 1 13 13 4 4 2
32 3 1 9 1 13 4 16 2 9 1 9 9 9 1 9 9 9 9 1 13 4 9 1 14 2 9 1 13 9 1 13 2
17 9 9 9 9 1 9 4 4 16 2 13 4 4 9 1 13 2
13 9 9 1 0 1 13 4 15 14 13 4 4 2
19 9 9 9 1 9 9 1 13 16 9 1 13 9 1 13 4 16 4 2
6 9 4 9 1 13 2
8 9 1 13 4 16 1 9 2
7 15 14 0 9 1 13 2
33 9 1 9 1 13 14 13 4 16 2 9 1 0 4 9 9 13 9 1 0 16 1 9 14 13 16 13 4 16 4 4 4 2
19 9 1 10 9 1 9 1 9 1 0 4 9 1 13 16 4 1 13 2
11 9 9 1 9 1 0 13 4 16 4 2
14 2 9 9 2 1 13 16 4 4 1 13 16 4 2
17 9 9 1 9 9 1 13 4 16 4 16 13 9 1 1 4 2
36 9 1 12 9 14 1 2 12 12 12 12 9 1 1 0 4 9 9 9 9 9 9 1 13 16 1 9 9 1 1 9 9 1 13 4 2
32 7 2 9 9 1 9 9 1 13 2 9 9 1 9 9 1 9 1 13 9 2 9 9 9 1 9 9 1 13 4 9 2
41 9 1 11 9 9 1 2 9 9 9 13 9 9 7 9 9 9 1 0 9 2 9 14 9 9 9 9 1 9 12 12 12 12 12 12 12 12 12 12 9 2
50 11 9 1 2 0 9 9 1 9 9 2 1 9 9 1 13 4 4 1 13 4 1 13 16 4 16 2 9 9 1 12 9 9 1 11 9 1 13 4 16 4 2 9 1 9 2 1 1 9 2
25 9 9 1 1 9 1 13 2 9 9 9 1 9 9 1 1 13 4 4 9 1 13 16 4 2
60 9 9 9 1 2 11 9 1 9 9 1 9 1 13 14 1 0 13 4 16 4 16 2 11 9 1 2 9 1 9 1 1 13 4 2 1 9 1 13 9 2 9 9 14 1 9 9 9 1 2 0 4 13 4 9 1 13 16 4 2
83 11 9 1 9 1 1 9 9 9 9 1 9 9 9 1 9 9 1 9 1 0 4 16 2 11 1 11 1 0 13 16 4 9 7 2 9 1 0 4 1 4 1 1 9 1 13 16 0 4 13 4 9 4 16 2 9 9 1 1 2 9 9 1 9 9 1 9 1 13 4 2 1 1 11 1 13 2 7 9 1 0 4 2
47 11 9 1 9 9 1 9 1 9 1 13 16 4 16 1 2 0 9 9 1 13 2 13 4 4 9 9 1 9 1 12 12 9 1 9 9 1 9 9 12 12 12 9 9 1 13 2
22 10 9 12 12 12 9 1 0 9 9 1 13 1 13 0 9 1 13 4 4 9 2
44 9 9 9 9 1 0 13 16 2 9 1 9 9 1 13 1 13 9 1 9 1 0 2 9 1 13 2 9 9 1 0 9 1 0 9 1 13 16 4 16 1 9 4 2
41 9 1 3 9 9 1 13 4 4 11 11 9 1 9 1 13 16 11 11 9 9 5 9 1 12 9 2 11 9 11 9 1 13 2 9 9 1 13 4 4 2
11 11 11 9 9 12 9 1 13 4 4 2
25 11 9 1 9 9 1 2 9 1 1 9 1 0 2 9 1 0 4 1 13 2 1 13 4 2
24 9 9 1 9 9 9 9 1 13 16 9 9 9 1 9 9 1 0 9 1 13 16 4 2
51 0 9 1 2 9 9 9 2 1 13 16 2 9 9 9 9 1 13 2 9 9 1 9 1 9 1 13 4 9 2 9 9 1 9 9 9 1 13 2 9 9 2 9 1 9 1 13 4 16 4 2
20 9 9 1 9 1 13 9 1 1 2 9 9 1 9 7 9 1 13 4 2
28 9 1 13 4 16 2 15 1 13 16 9 1 13 4 2 1 13 16 1 0 16 11 1 2 9 2 4 2
28 3 2 9 9 9 7 9 9 9 1 13 9 9 1 9 1 9 1 9 1 13 4 1 13 4 5 5 2
35 9 9 1 9 9 9 1 1 9 1 9 9 9 1 13 16 9 9 9 1 2 9 2 1 9 1 13 4 9 1 9 1 13 4 2
25 15 1 9 9 1 1 2 9 1 9 9 9 9 7 9 9 9 1 1 13 4 4 16 4 2
46 9 1 9 9 9 1 9 1 13 9 9 14 1 2 9 1 13 16 2 9 9 1 9 1 13 4 2 7 15 1 9 13 2 7 9 2 13 16 12 9 9 1 9 1 13 2
27 7 2 9 2 9 1 9 9 9 7 9 9 1 12 9 9 1 9 14 12 12 9 9 1 9 4 2
36 9 1 1 9 1 2 9 9 1 1 9 9 1 13 4 9 2 9 9 1 9 9 9 1 13 16 0 9 1 13 16 1 9 9 4 2
49 9 9 9 14 13 4 4 9 1 13 9 1 13 4 9 1 2 0 4 9 9 1 9 1 2 9 9 9 2 9 9 9 1 13 9 1 13 2 14 13 9 1 13 16 4 14 13 4 2
46 11 1 11 11 9 1 12 9 2 9 1 9 9 1 9 9 9 9 1 13 2 12 12 12 12 9 1 9 9 1 13 4 4 2 9 1 9 1 13 9 1 0 4 13 4 2
55 7 2 12 12 9 1 13 16 1 2 9 9 9 1 0 2 1 13 16 9 1 13 4 16 2 3 9 9 1 9 1 13 4 16 1 9 9 2 1 9 1 13 4 9 1 9 9 1 13 16 4 1 13 4 2
40 11 1 12 12 9 1 9 1 13 16 4 2 12 12 9 1 9 9 1 9 12 12 9 13 4 16 9 2 12 9 9 1 9 9 1 13 9 1 13 2
15 9 12 12 12 9 1 11 9 9 9 1 0 9 13 2
32 9 11 1 11 1 11 11 9 1 9 1 13 16 13 4 16 4 4 9 9 9 9 1 12 9 2 9 1 9 1 13 2
14 11 1 1 9 1 13 4 2 9 9 1 13 9 2
37 9 11 1 13 4 9 1 13 16 2 9 1 9 9 9 1 9 9 9 14 13 16 12 9 13 16 9 9 1 13 2 9 9 13 4 4 2
25 12 9 1 9 9 1 13 2 11 2 11 9 1 12 9 9 2 11 9 9 1 13 4 9 2
21 9 1 9 9 1 13 4 4 4 12 9 1 2 12 12 9 9 4 13 4 2
20 9 1 9 9 9 9 1 13 16 4 2 9 1 9 1 9 12 9 9 2
54 11 9 9 9 9 1 2 9 9 1 13 9 1 2 9 1 0 9 9 1 0 4 4 2 11 9 9 9 1 9 1 1 13 9 9 14 2 11 9 9 1 13 4 9 1 9 1 13 4 2 1 13 4 2
17 11 1 9 1 9 9 9 1 13 4 4 2 11 9 1 13 2
25 9 9 1 13 4 4 4 9 9 1 9 1 13 4 2 9 9 1 9 9 1 13 16 4 2
27 9 1 2 9 12 12 9 2 9 9 9 1 2 9 9 2 1 13 16 15 1 13 14 1 13 4 2
48 9 1 2 9 9 2 12 12 9 4 2 12 9 9 1 2 9 9 2 12 12 9 2 2 9 9 5 9 5 11 2 9 2 2 9 9 9 2 12 12 9 1 12 9 13 4 4 2
23 2 9 9 2 1 13 4 9 1 12 12 9 4 2 9 1 12 12 9 1 0 4 2
28 9 9 4 16 2 12 12 9 1 12 12 9 1 9 1 0 13 14 2 7 9 9 14 13 9 1 13 2
43 2 9 9 2 1 12 9 2 2 9 9 5 9 5 11 2 1 12 12 9 9 1 9 1 9 1 0 2 2 9 9 9 2 1 9 1 9 1 12 9 4 4 2
72 7 2 2 9 9 2 1 13 9 9 1 9 1 11 9 1 9 1 13 16 1 15 1 9 1 13 16 14 1 13 9 1 1 2 2 13 4 4 9 9 2 1 9 1 12 12 9 2 2 9 9 13 9 1 9 2 1 12 12 9 2 2 11 9 9 2 1 12 9 4 4 2
12 2 13 4 2 1 12 12 9 1 13 4 2
24 2 13 4 4 9 9 2 1 9 1 12 12 9 1 13 2 9 1 12 12 9 4 4 2
28 9 9 4 16 2 12 12 9 1 12 12 9 1 9 1 0 13 14 2 7 9 9 14 13 9 1 13 2
22 7 9 9 14 0 2 3 9 9 1 12 12 9 1 9 1 12 12 9 9 0 2
33 9 1 9 12 9 1 12 9 2 9 1 9 12 12 9 1 9 1 2 9 9 1 13 16 13 4 16 4 13 9 1 13 2
7 9 9 1 12 12 9 2
48 9 9 2 9 2 9 1 9 9 9 1 2 11 9 9 9 1 9 9 2 11 9 1 9 1 9 2 9 7 9 9 9 9 9 12 12 12 9 1 9 9 13 16 9 1 13 4 2
54 9 9 9 5 9 1 13 9 9 1 9 1 9 1 13 4 14 1 2 9 12 12 9 1 9 7 9 9 1 9 1 13 2 10 9 1 2 12 12 9 1 13 9 9 1 9 9 9 9 1 13 4 4 2
10 3 0 9 1 9 9 9 4 4 2
19 9 9 1 2 9 1 9 1 9 1 1 2 9 9 2 1 13 4 2
26 9 13 9 1 2 2 3 9 1 0 9 4 4 2 3 9 1 13 16 4 4 4 4 2 4 2
13 7 2 15 1 15 1 13 4 9 1 13 4 2
25 0 4 9 9 1 13 4 9 1 2 13 4 16 4 4 3 1 2 9 2 1 13 16 4 2
40 2 9 9 2 1 9 1 9 1 2 9 1 13 16 4 4 9 1 13 2 9 1 9 9 4 13 4 1 13 4 9 1 1 4 2 1 13 9 4 2
33 9 1 9 1 2 0 4 9 1 13 9 1 13 4 2 9 9 1 9 1 9 1 9 1 13 4 1 13 16 1 9 4 2
32 9 9 1 9 1 13 16 2 9 9 1 13 2 9 1 13 4 4 2 9 9 2 1 0 2 9 9 1 13 4 4 2
18 9 9 1 9 1 9 1 9 1 13 4 1 13 9 1 3 4 2
6 9 1 9 14 13 2
14 7 2 9 1 9 1 13 4 4 9 4 4 14 2
33 3 0 4 13 16 2 9 9 1 9 9 2 9 9 2 1 2 9 9 1 0 9 1 13 16 9 1 9 1 13 9 4 2
17 9 9 1 0 4 9 1 9 4 2 2 9 9 2 4 4 2
39 3 9 1 13 2 7 13 1 1 9 9 1 13 4 9 1 9 1 2 3 2 9 2 1 13 9 1 13 16 2 9 9 1 9 9 1 13 4 2
12 3 1 2 9 9 1 13 4 4 4 4 2
17 9 1 9 14 1 13 16 9 1 9 9 7 9 9 1 0 2
21 12 12 12 12 9 1 9 1 13 4 4 2 9 9 1 9 1 13 4 4 2
46 10 9 1 13 4 2 9 9 2 1 2 9 1 13 4 2 9 1 9 1 13 4 11 1 9 9 1 2 9 9 1 9 1 11 9 1 13 16 4 4 1 13 9 4 4 2
23 9 2 9 9 9 9 9 9 1 9 1 13 16 4 9 9 9 1 9 1 9 4 2
17 9 9 1 9 1 2 9 9 1 9 7 9 1 13 4 4 2
28 9 1 13 4 4 4 9 1 13 4 16 1 2 9 9 9 1 14 13 4 4 2 9 9 2 4 4 2
24 9 9 1 9 0 4 9 9 1 2 9 9 1 9 7 9 1 9 9 1 13 4 4 2
43 10 12 9 9 1 2 9 9 2 1 1 2 9 9 7 0 9 14 1 9 1 9 9 9 1 2 9 9 9 1 13 2 9 9 1 9 1 9 9 1 13 4 2
25 9 1 9 1 9 1 13 4 9 2 9 2 7 9 9 9 1 2 10 9 9 1 13 4 2
19 9 2 9 1 13 4 4 9 1 9 1 2 9 2 7 2 9 2 2
10 3 9 2 13 4 9 9 4 4 2
23 2 9 9 2 1 9 12 1 2 9 9 1 9 1 13 4 4 2 1 13 9 4 2
36 9 1 9 1 9 1 13 4 12 12 9 9 2 2 9 9 1 9 9 1 13 2 1 1 9 1 13 2 9 9 9 1 13 4 4 2
6 9 9 9 1 13 2
40 12 9 9 1 11 12 9 1 13 4 2 9 9 1 9 9 1 13 4 16 2 9 12 9 9 1 9 1 3 1 9 9 1 13 16 4 4 1 13 2
21 9 9 1 1 13 9 9 1 13 4 4 16 4 16 2 9 9 1 13 4 2
12 3 2 9 7 9 1 9 1 13 16 4 2
11 10 9 1 2 13 4 16 4 4 14 2
18 15 9 9 9 1 2 9 13 4 4 4 9 1 9 1 13 4 2
12 2 9 2 2 13 2 2 9 2 5 5 2
25 9 1 0 4 16 2 13 4 16 4 4 16 1 2 2 9 1 9 2 1 0 9 4 4 2
19 15 1 1 2 2 15 1 9 9 1 12 9 2 1 9 1 3 0 2
53 9 9 13 4 4 0 9 1 2 9 9 2 9 9 7 9 9 2 9 9 9 9 9 12 12 12 9 1 13 4 2 9 1 1 9 1 9 1 13 4 2 9 9 9 9 2 1 13 4 16 4 4 2
41 2 10 9 1 2 9 1 9 1 9 14 9 1 0 4 2 9 9 1 13 16 3 2 6 2 9 1 3 13 16 14 14 1 13 4 2 1 2 13 4 2
35 9 9 1 9 12 9 13 16 4 4 16 2 13 4 16 1 9 1 9 9 1 12 12 12 12 12 9 1 13 4 9 14 1 13 2
5 7 2 13 14 2
22 9 1 9 1 2 0 3 9 9 1 13 4 1 13 9 1 13 16 4 4 14 2
32 15 1 9 2 13 16 4 4 9 9 1 9 1 2 9 1 9 1 12 12 12 12 12 9 1 13 16 4 4 9 4 2
38 3 9 9 13 4 4 9 1 9 9 1 2 9 9 1 15 4 16 14 13 4 9 2 13 4 16 4 4 2 1 2 9 9 9 1 13 4 2
21 7 2 0 1 9 4 16 2 2 13 4 4 2 1 2 9 9 1 13 4 2
23 9 9 1 9 1 9 2 9 1 2 0 4 9 9 1 13 4 1 1 9 1 13 2
26 7 2 9 1 9 1 1 3 2 9 9 1 9 9 1 13 9 1 9 1 13 4 9 1 13 2
20 7 2 10 9 4 4 9 1 13 9 1 2 9 9 1 9 9 4 4 2
12 0 9 1 2 9 1 9 1 9 1 13 2
30 9 9 9 9 9 9 1 13 16 2 9 1 9 9 1 12 12 9 1 2 9 9 9 9 1 13 4 16 4 2
38 2 15 1 9 9 1 12 9 2 1 13 4 2 0 4 9 1 13 4 16 2 9 1 9 1 9 9 1 13 4 4 4 1 13 9 4 4 2
24 2 9 1 9 1 9 1 0 4 2 2 9 9 1 13 4 4 2 1 2 13 4 4 2
8 9 1 9 9 1 13 4 2
10 10 9 9 9 1 13 4 12 9 2
35 9 1 9 9 1 12 12 12 12 12 9 2 12 12 12 12 12 9 1 9 9 1 13 4 4 12 12 12 9 1 9 1 9 4 2
19 9 9 1 0 9 1 13 4 9 1 2 9 9 9 1 9 1 13 2
34 2 12 12 12 12 9 14 1 9 9 1 13 4 2 11 1 0 4 1 13 4 16 4 16 2 9 1 0 2 11 1 10 9 2
18 10 12 9 2 9 9 1 9 9 4 13 16 4 4 9 1 13 2
21 9 1 1 9 9 4 12 12 12 9 9 2 9 9 9 9 1 0 4 13 2
28 2 10 9 1 13 4 4 2 11 1 9 9 4 2 9 3 13 9 1 13 16 1 2 9 4 16 4 2
23 9 13 4 16 4 9 9 12 12 12 12 12 9 1 9 9 1 12 12 12 9 9 2
19 2 9 9 9 1 9 9 1 13 16 4 4 16 2 9 1 0 4 2
18 9 1 11 9 12 9 1 9 2 9 2 9 1 9 9 9 4 2
29 2 9 1 9 4 16 2 9 9 1 9 1 3 13 4 2 7 2 9 9 4 4 16 2 9 1 9 1 2
17 9 9 1 12 9 9 1 13 2 9 1 13 9 1 13 4 2
37 2 9 1 9 1 13 4 16 2 3 3 9 4 13 4 16 2 9 1 13 16 4 4 4 16 2 9 1 9 4 14 2 1 0 4 13 2
22 9 1 13 2 9 1 9 1 13 9 2 9 1 9 1 11 1 9 1 3 13 2
19 9 1 9 1 9 1 2 9 9 1 2 12 9 9 1 9 1 9 2
32 9 9 1 9 9 9 9 1 13 4 16 2 12 9 1 9 1 9 9 1 13 4 9 7 9 1 9 11 1 13 4 2
26 9 1 9 1 2 12 12 12 12 9 9 1 13 4 4 9 9 1 13 2 9 9 9 2 9 2
27 7 9 9 12 12 12 9 1 1 2 9 12 12 12 12 9 1 9 1 13 16 9 1 13 4 4 2
26 11 9 1 12 9 1 2 9 1 13 9 1 9 1 13 2 9 5 9 1 13 4 14 9 9 2
23 9 9 1 1 2 2 0 9 9 1 13 4 4 2 1 1 0 9 1 13 16 4 2
24 12 12 9 9 2 11 9 9 9 1 9 9 1 1 2 9 1 9 1 9 1 13 4 2
12 9 12 12 12 9 2 9 12 12 12 9 2
31 0 4 4 9 1 13 4 9 1 13 16 14 2 9 1 9 1 9 1 13 4 14 2 9 9 9 1 0 1 0 2
23 2 10 9 1 3 2 9 9 1 1 13 4 4 16 14 2 1 13 9 1 0 4 2
31 11 9 1 13 9 1 1 9 9 1 9 9 13 9 2 11 9 1 1 0 4 9 1 13 4 9 1 13 16 4 2
25 15 14 1 9 1 13 9 1 12 12 9 1 13 1 13 4 2 9 9 1 13 16 0 9 2
37 9 1 12 9 1 9 9 9 1 13 11 9 1 9 1 2 12 12 12 12 9 9 1 9 1 9 9 2 9 1 11 9 1 13 16 4 2
64 11 9 1 9 9 1 13 4 4 9 9 9 1 2 9 1 12 12 12 12 12 12 12 12 12 12 12 12 12 9 2 9 1 12 12 12 12 12 12 12 12 12 12 12 12 12 9 4 2 12 12 12 12 12 12 12 12 12 12 9 1 9 9 2
32 9 9 1 9 1 13 4 9 9 9 1 9 12 12 12 9 1 13 2 9 9 1 13 9 9 9 1 9 1 3 9 2
32 7 2 9 9 1 9 9 9 1 9 14 1 13 4 9 1 1 13 4 4 16 4 4 2 10 9 1 13 9 1 0 2
29 11 9 1 13 16 11 1 1 9 9 1 13 4 9 1 2 9 9 1 12 9 14 1 9 12 12 12 9 2
26 9 1 12 9 1 13 4 9 9 1 9 1 2 12 12 12 12 12 9 1 13 4 9 1 13 2
46 7 2 9 9 14 4 4 2 9 1 13 4 4 4 9 9 9 1 9 9 7 2 9 1 13 4 4 9 1 9 1 13 16 2 10 12 9 1 1 9 1 13 9 1 13 2
18 7 0 9 1 13 16 4 16 1 2 9 1 9 9 1 9 9 2
40 9 1 2 9 9 1 9 4 4 9 9 1 9 1 9 9 13 2 9 9 1 9 1 13 9 1 2 9 1 9 9 1 0 4 9 1 13 16 4 2
36 7 2 11 9 9 1 1 9 9 1 1 9 9 1 13 9 14 1 2 10 9 1 1 9 1 0 2 9 9 1 13 4 16 4 4 2
72 9 9 2 9 5 9 2 1 11 1 11 9 2 11 1 9 9 1 13 4 2 11 14 11 1 9 1 9 7 9 7 1 9 9 1 13 4 4 14 13 4 16 2 11 1 9 1 1 13 2 1 2 9 1 9 1 9 1 13 4 2 9 9 1 9 9 1 13 4 16 4 2
20 11 2 11 9 9 1 12 9 2 11 1 9 9 9 9 1 13 4 4 2
19 9 1 9 2 9 9 1 9 9 2 9 9 1 9 14 1 13 4 2
19 11 1 9 2 11 9 1 11 1 13 4 2 11 5 9 9 1 13 2
26 9 9 9 1 9 9 4 4 11 1 1 9 0 9 1 13 16 4 2 9 9 9 1 10 9 2
40 11 1 11 9 9 2 9 2 1 12 9 13 4 9 1 13 16 2 11 11 9 9 9 1 9 1 2 9 11 9 9 9 9 2 1 13 4 4 4 2
17 9 9 9 1 9 1 11 9 1 9 1 13 4 16 1 13 2
23 9 1 13 16 2 9 9 9 9 1 11 9 9 1 9 9 1 13 16 4 1 13 2
67 11 1 1 9 1 13 16 2 11 1 9 9 9 1 13 16 4 9 9 9 5 9 9 9 9 1 12 9 2 11 9 1 9 9 11 9 9 1 9 1 13 2 12 12 12 9 1 12 12 12 9 14 11 1 9 9 1 9 9 9 1 13 4 13 4 4 2
27 9 9 1 11 9 9 1 13 9 12 9 9 9 1 9 1 13 16 1 2 13 4 1 13 16 4 2
71 12 9 9 1 2 9 2 1 13 16 2 9 9 1 13 4 9 9 9 9 9 1 9 9 9 9 9 1 9 9 1 2 11 9 1 9 9 9 9 1 9 9 1 13 4 16 4 4 9 9 1 13 2 9 1 1 9 9 1 13 4 0 9 1 11 9 1 13 4 4 2
59 9 1 13 4 4 11 9 9 9 1 9 1 13 16 2 11 1 9 9 1 9 9 2 9 9 1 13 16 11 9 1 9 9 9 1 9 9 9 1 13 0 9 1 13 4 2 11 9 1 9 1 1 9 1 13 4 4 13 2
42 11 9 1 2 11 9 1 11 9 9 1 9 9 1 13 9 9 9 9 1 13 16 9 1 13 4 4 4 2 1 13 9 9 1 9 9 1 13 4 1 13 2
29 9 9 1 9 1 2 11 1 13 4 16 9 1 13 9 1 13 4 9 1 2 11 9 1 1 9 1 13 2
40 11 1 11 9 1 12 9 2 9 1 9 9 1 2 9 1 11 9 1 13 16 2 9 9 9 11 1 1 9 1 9 9 1 0 4 1 13 4 4 2
84 11 1 11 9 9 1 9 1 2 12 9 1 11 1 13 4 11 9 1 1 9 1 13 9 9 1 13 4 9 4 2 9 9 1 2 11 1 9 1 9 1 2 11 1 1 9 1 13 4 1 13 9 1 9 1 2 3 3 13 4 4 2 9 1 9 1 13 16 4 14 1 1 2 9 1 1 13 4 2 1 13 4 4 2
58 11 1 9 9 0 9 2 9 5 9 2 1 12 9 2 9 11 9 1 13 4 11 9 9 9 9 12 12 12 12 9 1 9 2 9 9 7 9 1 9 1 13 16 4 4 9 12 12 9 1 13 4 4 4 1 13 4 2
18 11 9 9 1 13 4 11 9 9 1 9 9 1 0 4 13 4 2
14 9 1 13 16 2 9 9 1 9 1 9 1 9 2
22 9 9 9 1 9 9 1 9 1 2 9 9 1 9 1 9 1 13 16 4 4 2
15 9 9 1 0 9 1 13 16 4 4 9 1 13 4 2
24 9 9 1 2 9 9 4 9 9 1 2 9 9 1 9 1 13 4 16 4 2 1 13 2
15 9 9 1 9 9 9 1 3 0 4 11 1 13 4 2
40 12 9 1 11 9 2 9 9 2 1 2 11 9 9 9 1 9 1 13 16 2 11 9 1 9 9 9 9 12 9 1 11 1 13 4 4 1 13 4 2
11 9 12 12 12 12 12 12 12 9 9 2
19 11 9 1 11 9 1 9 9 9 1 9 9 13 9 1 13 1 13 2
22 9 1 9 1 12 12 9 2 9 1 13 16 1 3 0 13 4 9 11 1 9 2
33 9 9 1 9 3 9 9 1 0 16 2 9 1 9 1 15 1 13 2 9 2 1 9 1 2 9 1 9 1 13 16 4 2
39 12 12 12 9 9 2 9 7 9 1 1 2 13 7 13 1 9 9 9 1 13 4 16 2 15 1 9 9 7 9 9 2 3 9 9 9 1 9 2
20 2 9 1 11 9 1 9 2 1 13 4 14 9 2 9 1 13 4 4 2
10 9 12 9 2 9 9 1 9 9 2
21 9 1 13 16 4 9 9 1 2 9 2 1 2 13 4 4 13 16 4 4 2
24 9 1 3 9 7 9 1 9 1 1 9 1 1 2 15 1 2 9 2 9 2 11 2 2
25 9 1 9 1 9 1 0 2 0 4 9 9 9 1 9 9 1 1 2 12 12 9 1 9 2
13 9 1 9 1 9 1 1 9 1 2 9 2 2
17 15 14 13 9 1 1 4 9 9 2 9 2 9 2 11 2 2
22 13 16 9 1 13 9 2 9 0 4 9 1 13 9 2 9 1 9 1 13 9 2
45 11 1 1 9 1 13 16 2 11 1 9 9 9 1 12 9 2 9 11 1 9 1 13 9 1 9 12 9 1 13 4 2 9 9 1 11 9 1 13 9 1 13 4 4 2
18 9 11 9 1 13 16 2 12 9 1 11 9 1 9 7 10 9 2
21 9 9 12 12 12 9 9 1 9 1 13 9 2 0 9 1 13 4 4 4 2
19 9 1 11 1 13 4 4 16 4 4 9 2 13 1 13 4 1 13 2
31 12 9 1 9 2 11 1 13 4 13 4 4 16 2 9 1 13 4 16 9 1 13 4 4 2 9 1 13 4 4 2
32 11 9 1 9 1 2 11 1 1 9 9 1 13 4 16 4 11 1 2 11 5 11 9 1 9 9 1 9 1 13 4 2
45 9 9 1 9 9 9 9 1 11 9 1 9 1 13 16 4 16 2 11 9 1 2 11 7 9 9 7 1 9 9 1 2 3 13 4 4 4 4 9 1 13 16 4 4 2
53 11 1 9 9 1 12 9 2 9 1 13 2 11 1 13 9 9 9 1 11 1 9 1 13 4 4 16 1 4 4 2 9 1 11 2 11 9 1 9 1 2 9 9 4 13 4 4 4 2 1 13 4 2
25 9 1 9 1 1 9 9 1 9 1 2 9 1 9 9 1 1 0 9 1 13 1 13 4 2
26 11 1 12 9 2 9 9 1 13 16 1 3 11 1 9 1 9 9 13 9 1 0 4 13 4 2
38 11 9 1 11 9 9 1 9 9 9 1 9 1 13 16 4 2 9 1 1 9 9 1 9 9 9 1 13 16 4 11 9 9 1 9 1 13 2
35 9 9 1 9 9 7 9 9 1 0 4 16 2 11 1 12 12 9 9 1 13 4 2 9 9 12 12 9 1 13 4 4 9 4 2
31 9 1 11 9 9 1 13 2 9 1 9 1 1 9 1 13 4 16 2 11 1 1 9 1 13 16 4 4 1 13 2
34 11 1 9 9 1 9 12 12 12 5 12 12 12 12 9 1 2 9 1 12 12 12 9 9 14 13 4 1 13 4 4 16 4 2
40 11 1 11 9 9 1 9 2 9 14 1 13 4 9 9 9 1 13 4 16 4 4 16 2 9 1 9 1 13 9 1 9 9 1 13 9 1 13 4 2
31 12 12 12 12 9 9 1 1 9 9 9 9 9 9 9 1 13 4 4 9 1 13 2 9 9 1 9 1 9 9 2
16 12 12 9 1 9 9 9 1 13 16 1 9 9 1 13 2
58 9 1 11 11 9 1 2 9 1 9 1 13 9 1 1 2 9 14 2 9 9 4 9 4 4 16 4 4 9 1 13 2 9 1 9 1 13 9 0 9 1 13 4 2 1 9 1 9 9 1 13 16 9 1 13 4 4 2
47 2 9 1 9 9 1 13 4 9 1 9 1 13 2 9 9 7 9 9 1 13 2 9 9 1 12 9 2 9 9 1 10 0 4 9 9 9 1 9 1 13 4 1 13 4 4 2
38 9 9 1 9 9 1 9 1 9 1 9 9 1 0 9 7 0 9 1 9 9 1 9 5 9 13 2 10 9 1 9 14 9 14 14 1 13 2
25 9 1 12 9 9 4 2 9 1 9 7 9 9 14 1 13 4 2 9 1 9 1 13 4 2
11 12 12 9 9 1 1 9 9 13 9 2
43 9 1 12 9 2 11 5 11 1 13 4 9 12 12 12 9 9 1 13 9 9 2 9 9 9 2 1 13 16 2 11 9 1 9 1 13 4 4 1 13 4 4 2
16 11 1 9 9 1 11 1 9 9 1 13 4 16 1 3 2
18 9 2 9 1 0 1 9 1 13 16 4 2 9 13 4 4 9 2
67 9 9 1 9 1 13 4 12 9 1 11 9 9 9 1 9 9 1 2 9 9 1 9 9 9 1 9 9 1 13 4 9 1 13 16 9 9 1 13 4 2 9 9 12 12 9 9 2 12 9 9 9 1 12 9 5 12 12 12 9 9 1 9 1 13 4 2
42 9 12 9 9 2 9 12 12 9 9 12 9 1 13 12 9 12 12 9 9 9 12 9 9 1 12 9 5 12 12 12 9 12 12 9 1 13 4 4 16 4 2
18 9 12 9 14 1 9 1 12 12 12 12 12 12 12 12 12 9 2
55 9 1 12 9 2 9 1 9 1 13 9 5 9 9 14 9 9 12 12 9 1 9 9 9 12 12 9 1 9 1 9 9 9 9 1 9 9 1 9 1 9 1 9 12 12 12 5 12 12 12 9 1 13 4 2
33 9 1 9 1 13 9 2 9 9 2 9 9 1 13 4 16 1 9 4 2 9 9 1 9 9 1 3 9 1 13 4 4 2
33 13 4 16 1 2 9 9 9 12 12 12 9 2 9 9 12 9 1 9 1 9 1 0 9 9 9 1 2 9 5 9 2 2
42 9 1 9 1 13 16 1 2 9 1 9 9 9 12 12 9 1 9 2 9 1 9 14 9 9 1 13 9 12 12 9 1 13 4 12 12 9 9 1 9 9 2
36 9 1 9 9 1 9 9 1 9 12 12 12 12 9 4 4 16 2 9 5 9 1 9 9 1 13 4 2 9 1 9 12 12 12 9 2
33 7 2 9 9 1 9 9 1 9 9 1 9 1 9 1 2 9 1 3 12 12 12 9 13 2 12 12 12 9 1 13 4 2
39 9 1 9 9 1 13 4 4 9 9 9 9 9 1 13 2 9 1 9 2 11 5 11 1 9 9 9 1 9 9 9 9 9 1 13 4 16 4 2
18 9 9 1 2 9 9 9 1 12 9 12 1 13 4 9 1 9 2
43 9 9 1 10 9 9 1 2 9 9 1 9 2 9 9 9 7 9 5 9 9 9 1 13 4 9 2 9 9 9 7 9 1 9 9 9 1 9 9 9 1 13 2
20 9 12 9 9 2 9 9 9 12 12 12 9 4 2 9 1 13 4 9 2
42 11 9 9 9 1 12 9 2 12 12 12 12 9 1 9 9 9 9 1 9 9 12 12 9 9 1 12 12 12 12 12 12 12 9 1 13 4 1 13 4 4 2
10 11 7 11 9 1 3 0 4 4 2
33 15 1 13 2 9 1 9 9 9 1 9 12 12 12 9 9 1 12 12 12 12 12 9 1 2 9 9 1 12 12 12 9 2
43 9 1 12 9 2 9 1 1 9 9 1 2 9 9 2 1 9 1 13 9 9 9 1 9 2 11 9 2 1 9 9 2 11 1 13 4 9 1 0 4 13 4 2
12 2 9 9 2 1 9 1 9 1 1 3 2
28 9 5 9 5 9 1 9 1 1 2 9 9 2 1 9 1 0 2 11 2 11 1 9 9 9 1 9 2
15 9 9 1 9 9 9 1 2 9 9 1 12 9 0 2
23 3 13 9 9 12 12 9 1 9 1 9 1 9 1 9 1 1 3 0 4 9 4 2
44 9 1 2 9 9 1 9 5 9 7 11 1 9 1 13 16 9 9 1 13 9 4 2 9 1 0 13 14 2 3 0 4 9 9 1 9 1 1 9 1 0 4 13 2
42 11 11 9 9 1 12 9 2 9 9 9 9 9 1 9 5 9 9 9 1 9 1 2 9 9 1 13 4 9 1 9 9 9 1 13 4 4 1 13 4 4 2
29 9 9 1 9 7 2 9 1 9 1 13 9 9 1 9 1 2 9 1 9 1 13 4 2 9 1 13 4 2
27 7 9 9 9 1 9 1 2 9 9 9 12 12 12 9 1 13 9 1 1 4 2 1 13 4 4 2
54 9 9 1 9 9 1 11 1 9 9 9 1 12 12 12 9 1 13 4 16 9 2 13 4 16 4 4 16 2 9 1 13 16 1 11 9 1 13 16 4 4 9 1 9 9 1 13 4 4 9 1 13 4 2
97 9 5 9 9 9 9 1 9 1 13 4 9 1 13 16 2 11 9 9 9 1 11 11 9 1 12 9 2 2 9 9 1 9 7 2 9 1 9 9 1 9 1 9 1 9 1 13 4 1 13 9 1 0 4 13 4 4 9 1 1 9 4 4 9 1 13 4 4 2 9 9 14 2 9 9 1 13 4 4 9 1 13 16 9 9 1 13 4 2 1 1 9 1 13 4 4 2
27 11 9 9 9 1 12 9 2 9 9 1 9 9 9 9 1 9 1 13 4 9 1 0 4 13 4 2
22 11 11 9 9 1 12 5 12 12 9 1 9 1 2 11 2 11 9 1 13 4 2
26 11 1 1 9 9 1 9 1 9 4 2 11 5 11 9 2 11 5 11 9 9 1 13 1 9 2
12 9 9 9 1 9 1 13 4 16 1 3 2
34 11 1 12 12 12 12 9 1 11 9 1 9 9 2 9 9 1 9 9 13 4 2 9 9 1 9 1 0 13 9 1 9 9 2
27 11 1 11 9 9 1 9 9 9 9 1 13 2 9 1 1 9 9 9 1 9 9 4 13 16 4 2
27 9 9 1 2 9 2 1 9 9 1 2 9 9 1 2 12 12 9 1 9 1 9 2 1 13 4 2
37 9 9 1 9 12 9 1 9 1 9 1 9 4 16 2 9 1 0 9 1 9 14 1 2 9 9 1 0 9 1 13 4 16 4 4 4 2
7 12 12 9 5 10 9 1
9 12 12 9 5 12 12 9 1 9
7 12 12 9 5 9 9 11
7 12 12 9 5 9 12 9
8 12 12 9 9 5 9 1 9
11 3 9 1 13 4 16 1 12 12 9 2
21 9 1 0 9 13 16 4 9 7 2 9 9 1 9 4 9 1 9 1 4 2
31 12 12 9 2 12 12 9 1 9 12 1 9 1 13 16 4 2 9 1 13 16 0 13 4 16 4 16 1 13 4 2
92 2 9 1 9 2 11 1 9 4 4 16 2 9 1 15 2 11 1 9 1 13 4 4 2 9 9 12 12 9 13 4 9 1 13 16 4 9 1 9 4 2 3 1 9 1 1 13 4 4 2 7 2 9 14 9 9 1 9 1 13 16 9 1 13 16 4 2 9 1 9 7 9 9 1 9 9 1 13 16 4 2 9 1 9 1 1 15 1 13 4 4 2
51 2 9 9 1 2 9 7 9 1 3 13 16 2 9 9 2 9 9 1 1 9 2 11 2 9 14 1 13 4 1 2 15 2 0 16 14 2 9 1 12 9 9 2 9 1 13 16 4 4 4 2
61 2 9 1 0 2 12 12 9 14 1 9 1 13 4 9 1 9 1 13 2 9 9 1 13 2 9 1 2 9 7 9 2 9 2 9 2 9 14 2 9 1 9 1 13 16 4 2 15 1 9 1 9 1 2 13 16 4 4 16 4 2
103 2 9 1 9 9 1 9 2 1 13 16 4 4 2 9 12 12 9 1 13 16 2 15 1 11 9 9 1 11 5 11 1 9 1 13 4 9 7 9 2 9 12 9 2 9 12 9 1 12 9 1 9 1 9 1 13 4 2 9 2 11 9 2 9 1 9 2 9 2 9 9 9 1 13 16 4 2 9 1 0 9 7 9 9 2 9 1 0 9 1 9 1 2 9 1 13 4 9 1 13 16 4 2
57 2 0 9 13 4 12 12 9 7 15 1 9 7 9 1 2 15 1 9 1 13 4 14 2 13 4 4 2 10 9 1 9 4 13 16 1 4 4 2 9 1 13 4 9 9 1 9 1 9 1 9 4 2 1 13 4 2
61 2 11 9 1 9 9 5 9 1 13 4 2 9 7 11 5 9 9 9 9 14 2 9 9 16 1 13 16 2 9 9 16 1 0 2 10 9 1 2 9 1 11 11 9 7 9 14 1 13 4 9 1 2 9 1 13 16 4 4 4 2
53 2 9 9 1 1 2 9 1 0 4 2 2 11 9 9 2 1 14 9 1 13 16 2 0 9 7 9 1 13 4 16 4 2 1 13 2 9 1 13 16 9 1 13 2 9 1 13 4 16 1 13 4 2
66 2 9 1 9 1 9 1 2 3 2 11 9 2 1 14 13 9 1 13 9 4 2 9 1 9 9 7 9 1 13 4 9 1 13 2 7 2 9 9 1 13 16 4 9 1 2 13 16 4 4 2 1 13 9 1 13 4 2 3 0 9 1 13 4 4 2
9 9 9 1 9 12 9 1 13 2
21 9 9 1 13 16 9 1 13 2 12 12 9 1 9 9 11 11 9 1 13 2
20 12 12 9 1 9 1 13 2 2 9 1 9 1 0 9 2 14 1 13 2
6 11 11 9 1 9 2
13 10 12 9 2 12 9 9 1 9 1 13 4 2
8 9 1 12 12 9 1 13 2
8 9 9 14 9 12 12 9 2
13 10 9 1 4 1 13 16 2 9 12 12 9 2
30 9 9 1 9 1 12 12 1 13 4 4 1 13 16 2 15 14 13 4 16 4 0 4 16 14 9 2 1 13 2
45 3 9 1 13 4 9 1 13 9 1 2 0 9 1 9 1 9 1 9 1 13 4 1 13 2 9 9 9 1 13 2 9 9 1 9 1 13 4 9 1 13 4 16 4 2
20 9 1 9 1 13 14 4 16 2 13 16 1 3 13 4 1 1 13 4 2
35 12 9 9 1 13 13 4 9 1 9 1 2 9 9 1 13 4 9 4 16 2 9 14 9 1 13 9 1 1 13 4 4 4 4 2
9 9 1 9 1 9 1 13 4 2
15 12 9 14 13 16 0 13 16 2 10 9 9 1 13 2
30 9 2 15 1 9 1 13 16 1 12 12 12 9 9 1 13 4 9 1 13 16 4 4 9 1 13 16 4 4 2
28 12 9 4 3 9 9 1 13 4 9 4 16 2 15 1 9 1 0 9 1 13 4 4 9 14 13 4 2
26 9 1 13 4 2 13 2 9 1 9 1 13 4 4 2 1 13 4 4 4 9 1 13 16 4 2
23 7 9 1 9 1 13 16 2 9 1 9 1 13 2 0 4 9 1 13 16 4 4 2
18 9 9 1 12 9 2 0 9 1 13 16 2 10 9 1 13 4 2
25 9 9 1 13 4 4 4 11 9 1 2 9 9 2 1 2 9 9 9 9 13 4 4 4 2
36 12 9 1 2 11 9 9 2 1 2 10 9 1 13 4 16 1 2 9 9 1 15 1 13 4 16 14 2 0 4 9 1 13 16 4 2
27 9 9 4 9 1 13 4 9 2 9 9 9 1 9 9 2 9 9 1 0 4 9 1 13 4 4 2
57 9 1 13 16 2 9 1 11 11 9 9 2 9 9 1 9 9 12 9 1 9 9 1 13 2 3 9 12 12 9 1 1 9 1 9 4 4 9 2 11 9 9 9 9 12 9 1 11 1 9 9 1 9 9 13 4 2
26 9 9 1 2 9 1 13 4 9 1 9 9 1 13 16 4 2 9 9 1 9 1 9 1 9 2
28 7 2 9 1 9 1 0 1 13 1 2 3 0 4 9 2 1 2 9 1 9 1 13 4 4 1 13 2
44 13 4 11 11 5 11 9 9 9 9 9 9 9 9 9 9 9 1 9 9 1 13 4 16 2 9 1 13 4 2 11 9 9 1 9 12 12 9 1 11 1 13 4 2
31 9 1 9 1 9 1 13 2 9 9 1 2 9 9 9 2 1 2 11 9 9 9 9 2 1 13 9 1 13 4 2
34 9 9 5 9 9 9 9 1 2 9 9 1 9 1 13 4 9 1 13 16 2 9 1 11 1 13 16 4 4 14 2 1 13 2
41 11 9 9 1 2 9 9 1 13 4 4 2 1 13 2 12 12 12 9 1 2 9 1 9 9 9 1 2 9 9 1 9 1 13 4 2 1 13 4 4 2
40 9 1 12 9 2 11 5 9 9 9 1 9 9 9 1 13 2 9 9 5 9 1 9 9 1 9 1 2 11 9 1 11 9 1 9 1 13 4 4 2
28 9 9 1 12 9 9 2 9 9 12 9 7 9 2 9 1 9 12 9 1 9 1 11 9 1 13 4 2
58 9 9 9 1 9 9 9 1 12 9 13 4 4 2 9 9 1 13 16 12 12 9 9 1 13 4 4 11 9 1 9 2 11 9 5 11 1 9 9 1 12 9 1 13 2 12 12 9 9 12 9 1 9 9 1 13 4 2
18 9 11 9 1 1 9 9 12 12 9 9 1 13 16 9 1 13 2
19 12 9 13 4 9 1 9 1 13 4 16 2 9 1 0 9 1 0 2
36 9 9 1 9 1 1 2 9 9 1 9 9 1 13 14 1 2 9 1 13 16 9 1 13 4 4 4 2 1 9 1 13 4 14 4 2
41 3 9 1 13 4 4 7 0 9 1 0 16 1 2 9 9 1 9 1 9 1 2 9 1 13 4 9 1 2 9 9 2 1 3 13 16 4 16 4 4 2
20 7 13 16 9 9 1 0 9 1 2 9 1 0 4 13 16 4 9 4 2
30 11 9 1 9 9 1 9 9 4 13 2 9 1 9 9 9 1 9 1 2 9 1 0 9 1 13 16 4 4 2
31 9 2 9 2 9 2 9 14 1 1 13 4 1 1 2 13 1 9 1 9 9 1 9 1 9 1 13 9 1 3 2
45 9 9 1 12 12 9 1 13 4 9 9 1 9 1 13 4 9 4 2 2 9 1 0 16 2 9 1 0 2 9 1 13 4 16 2 13 4 14 2 1 9 1 0 4 2
28 9 9 1 2 9 1 13 4 1 9 1 13 9 4 9 4 2 9 13 1 9 1 13 4 9 1 13 2
29 9 1 1 9 7 11 14 2 9 1 13 9 1 13 9 1 9 1 13 16 2 10 9 1 3 9 1 13 2
30 9 1 11 9 1 2 9 1 13 16 2 3 13 4 2 9 1 13 1 13 16 4 16 5 5 2 1 9 9 2
26 9 5 9 1 1 9 9 9 1 12 9 12 12 9 1 13 4 9 1 9 1 2 15 1 13 2
31 9 1 13 2 3 9 1 13 1 1 2 0 9 1 9 1 13 2 3 9 1 13 9 1 13 4 9 1 0 4 2
25 9 9 1 11 1 2 9 1 12 12 9 9 1 9 9 5 11 1 1 9 1 13 4 4 2
20 11 1 11 1 9 1 13 4 4 9 1 13 16 2 9 1 3 0 13 2
23 12 12 12 12 9 9 9 9 9 9 1 2 12 9 1 1 11 5 9 1 13 4 2
43 9 2 12 9 9 9 9 1 13 4 11 5 9 1 9 2 11 5 11 2 9 5 11 2 11 5 11 2 9 5 11 9 1 9 1 13 4 9 1 13 4 4 2
21 12 12 12 9 1 9 1 9 9 1 9 2 9 1 9 9 1 9 12 9 2
26 12 12 9 1 12 9 9 1 12 9 2 9 9 1 12 9 1 2 9 9 9 2 1 13 4 2
20 9 9 1 12 9 4 4 16 2 9 9 7 9 9 1 13 4 16 4 2
9 9 1 9 1 13 4 4 4 2
24 12 12 12 9 1 9 2 12 12 12 9 1 11 1 2 9 9 1 12 9 1 1 9 2
27 12 12 12 9 2 12 12 9 1 13 4 9 1 11 1 9 1 0 9 1 9 13 4 9 1 13 2
22 12 9 1 13 9 1 13 4 11 1 9 9 1 13 4 9 9 1 0 4 4 2
10 11 1 9 1 9 1 9 9 9 2
10 9 9 1 1 9 9 1 13 4 2
12 9 9 1 3 13 4 16 4 16 1 11 2
27 12 12 9 9 12 9 1 9 9 1 9 4 4 9 1 9 12 12 12 9 9 1 9 9 12 9 2
21 9 9 1 1 12 9 1 13 4 16 2 9 9 1 13 4 0 9 1 0 2
10 9 9 1 9 1 9 9 1 13 2
29 9 1 13 4 4 9 1 1 2 12 12 9 9 9 1 11 5 11 7 9 1 9 5 11 1 9 1 13 2
24 9 1 12 9 9 9 1 13 4 11 1 9 1 11 5 9 1 13 4 2 9 1 13 2
13 9 1 11 9 1 0 4 9 1 13 4 4 2
23 11 1 9 9 1 13 16 2 9 1 9 1 9 1 13 2 0 4 9 1 13 4 2
19 2 9 1 9 2 1 13 4 9 9 14 1 2 9 9 13 4 4 2
10 9 9 1 13 9 1 1 11 9 2
24 9 1 1 9 1 0 9 1 13 11 11 1 9 4 15 14 13 4 14 1 9 1 9 2
15 9 1 9 9 1 12 9 1 11 1 9 11 1 13 2
25 9 13 16 1 9 9 1 9 2 11 2 11 2 11 2 11 2 11 7 9 11 1 12 9 2
21 11 11 9 13 9 11 9 1 9 9 1 13 16 2 9 1 15 1 9 9 2
27 12 12 12 12 9 1 11 9 1 9 9 9 1 13 11 1 2 9 1 9 1 15 14 13 4 14 2
13 9 9 1 12 9 1 13 2 9 9 1 13 2
17 12 9 9 1 9 2 12 9 9 1 12 9 9 9 1 13 2
18 11 1 9 9 1 2 12 9 1 11 2 12 9 1 11 1 9 2
8 9 1 15 1 9 12 9 2
28 9 1 11 1 9 1 9 12 2 9 12 2 9 12 14 9 12 2 9 12 2 9 12 1 13 4 4 2
41 12 9 1 13 4 16 1 2 9 1 9 9 1 13 4 16 4 9 1 13 2 2 9 9 1 9 2 9 1 1 9 1 9 1 13 4 2 1 13 9 2
16 9 1 1 9 1 12 9 13 2 9 9 1 9 1 13 2
22 9 1 13 4 4 9 1 13 1 11 1 9 9 1 9 1 13 4 9 1 13 2
19 9 1 11 1 9 1 9 9 2 11 1 9 9 9 1 9 1 13 2
24 9 1 9 9 1 11 1 9 9 1 13 2 9 7 9 1 13 2 9 1 9 1 0 2
19 11 1 9 1 9 9 12 9 1 13 4 4 9 2 9 9 1 13 2
15 9 1 13 4 9 1 9 1 0 4 9 1 13 4 2
34 3 9 1 13 4 4 4 9 2 9 9 1 14 9 9 1 13 4 16 4 4 9 1 13 16 2 9 1 13 4 4 1 13 2
9 9 1 9 9 1 9 1 9 2
13 9 9 4 13 16 2 11 1 9 1 13 4 2
23 11 1 9 2 11 1 9 1 13 2 11 9 1 13 9 9 1 15 14 13 4 14 2
23 9 1 13 16 2 9 9 1 13 2 9 1 13 9 1 0 13 9 1 13 14 4 2
33 11 1 11 9 9 1 9 9 9 1 13 2 9 1 9 2 11 9 1 12 9 2 11 1 9 9 1 0 4 13 4 4 2
60 11 9 1 2 9 1 13 4 16 1 2 15 1 13 16 4 4 11 1 9 1 13 9 4 2 1 13 2 12 12 12 12 9 9 1 11 1 1 9 2 12 12 12 12 9 1 9 9 9 1 13 16 4 9 1 0 4 13 4 2
27 9 1 9 9 9 1 13 16 2 11 9 9 1 13 4 4 9 9 1 9 12 12 12 12 12 9 2
35 9 9 1 11 9 1 13 4 16 1 2 2 9 9 4 9 1 13 2 9 1 13 16 9 1 3 13 16 4 2 9 1 4 4 2
51 9 1 9 9 9 9 9 9 12 9 1 12 9 2 11 9 1 12 9 1 13 2 11 1 11 1 12 5 12 1 13 16 9 9 9 1 13 2 9 9 1 12 9 12 9 12 9 1 13 4 2
23 9 12 12 12 9 9 9 9 9 1 9 12 1 13 2 12 9 1 9 9 1 13 2
30 9 9 1 9 1 12 9 4 2 9 9 1 9 1 12 9 1 9 1 13 2 9 9 1 9 1 13 16 4 2
32 12 9 1 9 2 11 9 2 11 9 2 11 9 2 9 9 1 11 9 1 12 9 1 9 1 9 9 9 1 13 4 2
26 15 1 13 9 1 4 4 16 2 0 9 7 9 9 1 13 2 9 1 9 1 13 16 4 4 2
15 9 9 1 9 1 1 2 9 5 9 1 13 4 4 2
19 9 1 9 9 9 9 2 9 1 9 12 9 1 9 9 9 1 9 2
15 12 9 1 9 1 13 9 1 2 9 1 9 1 0 2
24 9 1 13 4 9 1 1 9 1 0 2 9 1 9 12 9 1 13 9 1 0 9 4 2
14 9 1 9 2 9 9 2 9 9 1 9 1 13 2
32 9 1 9 9 1 13 4 16 2 9 9 1 13 16 9 11 1 11 9 9 1 12 9 1 13 14 9 9 1 13 4 2
18 9 9 1 13 4 4 11 9 1 11 9 1 9 1 13 16 4 2
12 11 9 7 11 9 1 2 3 9 1 13 2
24 9 1 13 4 4 11 9 1 9 1 9 9 1 0 4 11 9 1 3 13 14 1 9 2
27 12 9 1 12 12 9 1 9 9 1 13 4 9 1 2 9 11 11 1 9 1 0 4 9 1 13 2
18 11 11 1 12 9 9 9 1 9 9 1 13 2 9 1 13 4 2
42 11 9 9 1 13 16 9 1 12 9 9 1 13 4 11 9 1 2 9 1 13 4 11 9 1 13 2 0 4 9 1 13 16 13 9 9 1 9 1 13 14 2
33 12 9 1 9 9 9 2 9 9 9 9 1 9 9 1 9 2 9 1 9 9 12 9 1 9 9 1 13 16 4 4 4 2
10 0 1 11 2 11 2 11 4 4 2
7 13 4 16 13 4 4 2
17 11 11 2 11 1 9 1 9 1 3 9 1 9 1 13 4 2
15 9 1 9 1 1 9 9 1 11 9 1 13 16 9 2
31 9 1 13 4 16 12 9 1 13 4 16 2 9 5 11 11 1 9 7 9 1 9 9 1 9 1 9 1 13 4 2
36 11 11 1 9 1 12 9 9 12 12 9 2 12 9 9 1 12 12 9 1 2 9 1 13 16 4 4 9 1 3 9 13 16 4 4 2
42 11 9 1 12 12 9 2 12 12 9 1 13 16 3 13 4 2 9 2 9 1 11 9 1 9 1 9 9 1 13 16 12 12 9 1 13 16 9 1 13 4 2
25 11 11 1 13 16 1 2 9 1 9 9 1 9 9 13 16 1 9 9 1 11 9 9 4 2
36 9 1 9 9 1 13 2 12 9 12 9 1 0 9 1 9 1 13 9 1 9 9 9 1 1 11 1 12 9 1 0 9 1 13 4 2
70 7 2 11 11 1 2 9 12 9 1 13 16 1 9 4 4 2 9 9 1 13 4 4 2 3 9 1 13 4 2 11 1 13 16 4 16 2 15 1 9 1 9 4 1 13 16 2 9 1 13 16 1 9 1 0 13 16 4 16 4 2 1 9 9 1 13 4 4 4 2
33 9 1 0 4 15 14 9 1 13 16 4 4 11 1 2 9 1 13 4 9 1 2 9 1 13 4 4 2 1 9 1 13 2
18 9 2 11 11 2 11 11 1 13 16 9 9 1 13 4 4 4 2
24 2 0 4 2 9 1 3 4 4 2 9 1 1 3 13 16 4 4 2 1 0 4 9 2
30 13 9 1 13 4 16 14 2 9 9 7 9 9 9 9 1 9 1 13 4 2 9 9 1 9 1 0 13 4 2
20 11 11 5 11 11 1 13 9 1 13 16 1 11 1 9 1 13 11 9 2
17 11 9 1 11 11 1 13 4 2 9 9 1 9 9 1 13 2
16 9 1 9 4 16 9 1 13 9 1 1 9 9 1 1 2
9 2 9 2 9 2 2 9 2 9
9 2 9 1 13 9 14 1 9 2
5 9 12 12 9 9
15 11 12 12 9 2 9 1 9 1 9 1 13 4 11 2
20 9 9 1 13 9 1 2 0 4 9 1 9 1 9 1 3 1 13 4 2
24 9 9 1 13 4 11 11 9 2 9 1 13 9 2 1 11 11 9 1 9 1 13 4 2
15 9 1 11 9 1 13 4 16 1 12 12 12 12 9 2
47 2 13 4 1 13 16 4 4 4 16 2 3 12 12 9 9 1 13 16 4 4 2 15 1 9 12 9 1 9 9 1 13 4 9 4 4 4 2 13 16 4 9 13 4 4 14 2
11 11 9 1 0 4 9 1 9 1 9 2
7 9 1 9 1 13 4 2
59 11 9 1 13 16 9 2 0 9 2 9 1 0 16 2 15 14 1 9 1 9 7 9 1 13 2 9 9 1 13 4 16 2 11 9 1 13 16 4 4 0 9 1 13 4 4 4 4 2 1 13 9 1 13 4 9 1 13 2
5 15 1 13 4 2
40 2 9 1 13 16 1 2 9 1 9 9 1 13 4 16 2 13 4 16 4 16 4 14 14 2 9 1 15 1 13 16 14 2 1 13 4 16 13 7 2
35 2 9 1 13 9 2 1 1 2 9 7 9 9 1 13 16 13 4 2 9 9 1 9 1 13 16 4 9 1 9 1 9 1 13 2
24 2 0 4 9 1 13 9 1 13 9 1 13 9 2 1 11 9 1 3 13 4 9 4 2
23 9 9 1 11 11 9 9 9 1 11 11 14 2 11 9 2 1 9 2 9 1 13 2
18 9 1 9 1 9 2 9 9 1 13 11 1 9 14 9 0 4 2
15 2 0 9 1 13 4 16 2 13 4 16 0 2 4 2
20 9 1 11 9 1 9 1 1 9 1 4 4 9 14 1 9 1 13 4 2
11 9 1 9 1 11 9 9 1 13 4 2
17 11 9 1 0 4 4 14 4 4 2 0 9 14 13 16 4 2
33 11 9 9 2 9 2 1 2 9 9 1 9 1 11 9 1 2 9 2 1 13 4 4 9 1 9 1 13 16 4 16 4 2
33 9 9 1 13 16 3 9 1 13 4 11 9 1 2 9 1 13 16 9 1 13 4 4 9 1 2 11 9 1 1 3 13 2
54 2 9 1 9 1 12 9 14 1 9 1 13 16 2 9 1 3 1 13 4 9 1 0 2 9 4 2 13 4 16 1 13 4 16 1 2 13 16 1 9 14 2 0 9 1 11 9 1 13 4 16 4 4 2
10 10 9 1 11 9 9 1 0 4 2
31 12 12 9 1 13 16 1 9 2 9 1 13 2 2 12 12 12 12 9 9 9 11 2 1 11 11 9 1 13 4 2
25 11 1 9 1 9 9 9 1 13 16 4 4 11 11 9 1 2 6 2 1 13 16 4 4 2
43 2 9 2 11 1 3 0 9 1 13 16 4 2 15 1 13 4 4 16 4 14 2 15 1 12 12 9 1 13 16 2 0 9 1 9 1 13 16 4 16 0 4 2
15 9 9 1 1 9 1 2 9 9 2 1 13 4 4 2
13 9 9 1 11 9 1 9 9 9 1 9 4 2
25 9 1 9 9 14 9 9 1 9 14 4 4 16 2 9 9 2 1 9 1 0 4 13 4 2
30 9 1 9 1 1 2 9 9 1 13 4 3 1 2 3 1 13 16 4 9 9 9 12 9 1 9 1 13 4 2
35 11 1 13 4 9 2 9 1 13 4 9 12 9 2 11 9 9 9 2 1 12 9 9 12 9 1 11 9 1 11 9 1 13 4 2
39 9 1 11 2 11 2 11 14 12 9 12 12 12 9 1 9 9 1 9 1 11 1 12 9 2 9 1 12 9 1 13 4 4 2 9 1 13 4 2
17 3 13 4 4 16 1 11 1 9 9 1 2 9 14 13 2 2
32 9 1 13 9 1 13 16 13 16 4 4 9 1 2 9 1 9 1 13 1 13 9 1 2 11 9 9 1 9 1 13 2
46 11 9 1 1 2 9 1 9 0 4 9 9 1 13 0 9 1 13 4 11 9 2 9 1 9 1 9 9 11 9 1 9 5 11 2 14 1 0 9 1 9 1 13 16 4 2
51 9 11 5 11 9 1 12 9 9 2 9 1 11 9 1 9 9 12 9 5 12 9 1 9 1 13 4 4 1 13 4 9 1 2 9 9 1 1 9 9 1 13 9 9 9 1 13 4 4 4 2
14 9 1 9 1 9 1 9 9 1 9 9 4 4 2
37 10 9 1 9 9 9 1 2 9 1 9 1 9 1 9 1 9 12 9 4 16 2 9 1 13 2 9 1 13 4 16 9 1 12 9 9 2
92 9 1 9 9 2 9 11 1 13 4 11 9 11 9 1 9 2 11 11 9 1 2 11 9 1 9 1 13 2 9 12 12 9 9 2 9 1 9 1 13 16 12 12 9 9 1 12 9 1 13 16 4 16 1 13 4 2 12 12 9 12 9 9 2 9 1 13 16 4 16 2 12 9 1 9 1 13 4 4 4 2 1 9 1 9 1 9 1 0 13 4 2
127 11 9 9 1 13 16 2 9 9 1 13 11 9 9 1 1 9 12 12 12 9 1 2 9 9 1 1 9 12 12 9 1 9 9 1 13 4 4 16 4 4 16 2 2 9 9 1 9 2 1 9 1 2 9 1 9 1 12 9 0 13 4 0 4 4 9 9 11 9 11 2 9 9 2 11 9 9 1 2 9 1 13 16 4 16 1 13 4 4 2 9 1 3 4 16 2 9 1 11 9 1 9 4 16 9 1 13 16 4 4 4 2 9 1 13 1 1 3 13 4 4 2 1 13 16 4 2
40 9 1 1 9 1 9 9 7 9 1 9 9 9 1 13 16 2 9 9 1 9 9 1 13 4 1 13 16 4 16 2 9 1 9 1 9 9 1 13 2
72 9 1 13 4 16 4 9 11 9 9 9 9 1 11 11 9 9 1 2 9 1 9 1 11 12 12 9 14 1 1 13 16 9 1 9 12 9 14 0 2 9 1 9 9 1 9 1 9 1 13 16 4 4 4 4 2 1 9 1 0 9 4 4 4 9 1 13 4 16 4 4 2
23 9 9 1 13 4 11 11 9 1 9 9 12 12 9 2 9 9 12 12 9 1 9 2
18 9 9 9 12 12 9 1 13 4 11 9 9 1 13 16 4 4 2
23 13 4 4 1 13 4 12 9 1 9 7 9 1 0 9 1 9 1 9 1 13 4 2
31 2 9 9 1 9 2 1 9 2 9 9 9 9 1 1 2 9 1 11 9 9 1 9 1 9 1 9 1 13 4 2
38 9 1 13 16 13 4 9 1 9 1 2 11 9 1 9 1 1 13 16 4 9 1 9 2 3 0 4 13 16 4 9 2 1 13 16 4 4 2
46 11 9 11 1 9 1 13 1 9 9 2 11 11 9 1 9 11 9 1 2 9 1 12 9 14 9 1 13 16 4 4 2 9 9 4 1 13 16 4 4 16 2 1 13 4 2
50 9 1 9 1 9 1 9 1 9 1 1 13 4 4 4 9 9 2 11 11 9 1 13 16 2 9 9 1 12 12 12 9 13 16 4 9 9 9 1 9 1 2 9 1 9 12 12 12 9 2
24 9 9 1 11 9 9 1 2 11 9 9 1 12 9 9 1 9 9 1 11 1 9 9 2
20 12 2 12 9 1 9 9 1 13 4 2 12 9 1 13 4 9 4 4 2
68 11 9 1 2 12 9 1 9 11 1 3 4 4 16 1 11 9 14 1 11 9 1 9 1 0 2 15 1 13 16 1 3 9 1 13 16 4 4 2 3 13 4 9 1 13 4 16 9 2 9 1 13 16 9 1 13 2 9 1 9 1 13 4 2 1 13 4 2
29 9 9 1 11 9 9 1 11 11 9 1 13 4 4 1 13 4 11 11 9 1 11 9 11 1 9 1 13 2
53 9 1 9 1 2 15 1 9 9 1 12 9 9 13 2 9 9 1 11 11 1 1 13 16 4 4 2 15 1 13 1 9 14 9 9 1 9 1 13 14 3 13 4 9 4 16 2 1 13 16 4 4 2
20 9 7 9 9 9 1 9 9 2 9 9 2 1 2 9 1 12 9 14 2
11 9 12 9 1 9 12 9 14 13 4 2
15 9 1 12 12 12 12 12 12 12 12 12 12 12 12 2
65 9 9 9 1 0 9 9 1 13 4 4 4 11 9 11 9 1 9 1 13 9 9 2 9 2 1 9 12 12 9 1 12 9 2 9 14 1 9 1 13 4 4 4 1 13 16 2 9 9 1 9 9 9 1 9 9 9 1 11 9 1 13 4 4 2
44 11 9 11 9 1 2 9 9 2 9 1 9 9 2 9 1 1 9 9 1 13 2 9 9 1 2 9 1 9 1 9 1 13 16 4 4 2 1 13 4 16 4 4 2
51 9 9 1 9 9 7 9 9 1 13 16 2 9 9 9 1 9 9 9 1 9 1 13 2 9 1 13 16 2 9 14 1 9 9 1 13 2 9 1 13 16 9 9 1 13 4 4 1 13 9 2
53 13 4 4 4 9 9 9 1 2 9 1 9 1 1 9 1 13 4 9 1 0 4 16 2 13 4 4 4 9 1 3 9 1 13 4 2 15 1 9 1 13 4 4 9 1 13 4 2 1 13 16 4 2
20 2 9 13 4 2 1 13 9 1 11 9 1 9 14 1 13 13 16 4 2
31 2 9 1 0 13 2 1 1 13 4 9 1 13 4 2 13 4 9 1 9 1 9 1 13 4 1 13 16 4 4 2
39 9 1 1 9 9 7 9 14 9 1 9 9 1 9 1 13 4 16 1 9 1 2 9 9 1 2 9 9 2 0 4 9 2 1 13 4 16 4 2
29 9 9 1 13 16 2 10 9 1 9 1 9 9 9 9 1 2 11 9 9 1 9 14 1 0 13 4 4 2
31 9 9 1 2 13 4 4 4 9 9 1 9 1 9 2 13 4 4 4 9 4 2 9 1 13 4 9 1 13 4 2
49 2 12 12 9 1 9 9 2 1 13 10 9 1 2 12 12 9 14 13 16 2 15 14 12 9 1 9 1 13 2 12 9 1 13 4 16 2 9 9 4 9 1 0 2 1 13 4 4 2
49 7 2 0 1 9 1 13 16 4 9 1 9 1 9 1 13 9 2 9 9 1 9 9 1 13 16 2 13 16 1 15 1 9 4 16 2 0 9 1 13 4 2 1 9 1 13 4 4 2
52 9 9 1 13 4 9 9 1 13 9 2 11 9 9 9 9 2 1 11 9 9 1 2 9 0 9 2 9 9 1 9 9 1 13 9 9 14 1 9 14 13 4 4 9 1 13 2 1 13 16 4 2
55 12 9 9 12 9 12 12 12 9 9 2 11 9 5 9 1 9 9 12 12 9 1 9 4 2 11 9 1 9 9 2 11 5 9 2 1 2 13 4 4 2 1 1 9 1 9 12 9 9 9 9 1 13 4 2
42 9 9 9 9 12 12 12 9 1 9 1 13 4 2 9 1 9 9 1 11 9 1 9 9 1 12 9 1 13 4 16 2 12 9 1 9 1 13 4 9 9 2
13 13 12 12 9 1 9 11 1 13 4 16 4 2
31 9 9 2 11 2 1 9 1 9 9 1 13 16 4 16 2 9 9 1 11 9 1 2 9 1 9 14 1 9 9 2
57 9 1 13 4 9 9 1 9 1 13 2 9 11 1 9 9 9 9 1 9 1 9 9 1 9 7 9 1 9 9 13 4 2 9 1 9 9 1 9 1 9 1 13 2 13 4 4 9 1 12 9 2 0 4 13 4 2
34 9 9 1 9 9 1 13 16 3 9 9 1 0 9 1 13 16 1 15 14 13 4 4 4 9 1 0 2 9 1 9 1 13 2
26 11 9 1 1 9 9 1 9 9 1 14 13 4 2 9 9 1 13 9 1 13 4 16 4 4 2
40 10 9 2 9 1 13 9 9 1 11 1 9 1 9 2 9 15 14 1 9 1 13 2 9 9 1 9 1 13 4 2 9 1 13 9 1 13 16 4 2
18 7 2 9 2 9 9 1 9 1 13 4 9 1 15 14 0 4 2
21 9 9 1 13 16 2 13 4 4 16 1 11 9 1 13 12 12 9 1 9 2
27 9 1 9 9 1 9 1 0 9 1 3 0 1 13 4 4 2 9 1 9 1 13 9 1 13 4 2
34 9 1 9 9 1 11 9 9 1 9 9 9 1 13 16 9 9 1 9 1 13 2 11 1 13 2 9 1 9 1 13 1 13 2
21 12 9 9 12 9 12 12 12 9 9 2 11 9 1 9 1 9 1 13 4 2
23 9 1 9 1 13 16 2 9 9 1 11 9 9 1 9 1 0 9 1 12 12 9 2
8 9 1 9 1 9 1 9 2
39 11 9 11 9 11 1 9 2 9 9 11 11 2 9 1 9 1 2 9 14 9 12 12 12 9 1 13 4 16 4 4 9 1 12 9 2 13 4 2
33 3 13 4 4 9 2 9 1 13 16 13 4 4 1 13 4 2 11 9 9 9 1 0 4 9 1 13 16 13 4 16 4 2
35 9 9 9 7 11 9 1 13 16 2 12 9 9 12 9 9 2 11 9 1 2 9 1 9 1 13 16 4 2 1 9 1 13 4 2
28 13 4 9 2 9 1 9 12 9 9 1 9 14 1 9 9 1 9 1 9 14 1 13 4 16 4 4 2
18 13 4 4 9 1 3 2 9 9 1 9 1 13 4 9 4 4 2
13 9 1 12 9 1 9 1 9 12 9 1 13 2
30 9 1 13 4 12 9 9 1 1 13 16 4 9 1 2 3 13 4 4 4 9 1 13 16 13 4 1 13 4 2
24 13 4 16 4 4 9 1 2 9 14 1 0 4 9 2 12 9 9 1 3 13 4 4 2
33 11 9 9 1 1 2 9 1 1 9 9 12 12 9 1 9 1 13 16 4 4 1 13 9 1 13 2 9 1 13 16 4 2
16 9 1 9 1 2 9 9 9 9 2 1 9 1 13 4 2
13 9 2 9 12 12 9 9 12 12 9 9 2 2
33 9 1 9 12 2 12 2 12 2 12 2 12 12 2 12 12 2 12 12 2 12 12 2 12 12 2 12 12 2 12 12 9 2
6 9 1 13 16 4 2
18 9 1 2 9 9 2 1 13 16 4 16 2 9 1 9 1 13 2
18 9 1 9 1 2 9 2 1 13 16 2 13 9 2 1 13 4 2
102 2 9 1 9 9 9 1 9 1 9 2 14 1 13 16 9 12 12 9 9 1 9 1 13 4 4 2 9 9 9 1 13 16 4 11 9 11 9 2 9 9 9 9 9 2 11 11 9 1 12 9 2 2 9 1 13 16 1 13 4 16 9 1 13 4 2 9 1 9 9 1 9 1 9 1 13 9 4 2 1 13 2 9 9 1 13 9 9 9 1 9 1 9 1 2 9 9 2 1 13 4 2
55 9 9 9 9 9 1 9 9 1 9 1 13 4 7 9 9 1 9 1 13 14 1 2 9 2 9 1 2 9 9 1 2 9 1 13 16 4 1 13 4 16 4 16 2 9 1 13 4 4 2 1 13 16 4 2
23 9 9 9 9 1 2 9 1 13 16 9 5 9 1 9 9 1 13 9 1 9 9 2
27 9 9 1 9 9 1 13 2 9 1 9 9 13 9 9 9 12 9 1 9 1 13 16 13 16 4 2
25 11 9 1 12 12 12 12 9 1 13 4 2 9 1 0 13 9 1 9 12 12 9 1 13 2
19 12 12 9 9 2 9 9 1 9 9 1 0 4 9 9 1 13 4 2
54 9 9 1 9 9 1 13 4 12 12 9 9 9 2 11 9 1 9 9 1 13 4 16 2 2 11 9 1 9 9 1 1 9 1 1 9 9 1 9 2 1 9 1 13 4 9 12 12 9 2 13 4 4 2
61 11 9 1 10 9 9 12 9 9 1 9 9 1 13 11 11 5 9 9 9 9 9 9 1 13 2 2 9 9 14 1 9 1 9 1 13 2 9 9 1 9 1 13 4 2 9 7 9 1 9 1 0 2 1 9 1 9 1 13 4 2
53 11 9 1 2 9 1 1 9 5 9 1 9 1 13 13 7 13 7 13 16 9 1 9 1 13 9 1 9 2 7 2 9 1 1 9 9 1 9 1 9 9 9 1 9 1 13 4 4 2 1 13 4 2
28 11 9 1 9 9 9 1 2 9 9 2 1 13 2 9 9 1 13 9 1 13 9 1 13 4 16 4 2
42 9 9 9 9 9 9 1 13 16 2 9 1 0 4 13 9 9 1 13 16 1 2 9 1 9 1 9 9 1 13 9 9 1 9 9 1 13 4 4 1 13 2
76 9 9 1 0 11 11 5 9 9 9 1 2 9 9 14 9 1 0 4 9 1 13 4 3 2 9 9 9 1 9 1 13 16 2 9 1 13 16 9 1 13 4 4 4 2 9 1 13 4 9 1 2 9 9 1 13 9 1 13 4 9 9 9 1 0 16 4 1 4 14 2 1 13 16 4 2
50 12 9 9 12 12 9 9 2 11 9 11 9 11 9 2 9 9 9 9 2 11 11 9 9 9 12 9 1 13 4 9 7 9 1 13 16 4 16 1 11 9 1 13 2 11 9 1 13 4 2
25 9 1 1 2 9 1 11 11 9 2 9 2 14 1 9 9 12 12 9 7 2 9 12 9 2
21 9 9 14 1 9 1 9 1 9 1 4 4 9 1 13 4 4 16 4 4 2
30 11 9 1 9 9 1 13 4 9 12 12 12 9 9 12 9 9 1 9 9 14 1 9 1 2 13 4 4 4 2
16 9 9 1 11 9 1 9 9 13 16 4 4 9 4 4 2
38 11 9 1 9 1 9 9 1 9 9 9 9 1 13 4 9 12 12 12 12 12 12 12 9 9 1 9 9 9 9 1 12 9 2 13 4 4 2
34 15 1 13 16 2 9 9 9 1 9 1 2 9 1 9 9 1 9 1 0 2 9 9 1 9 1 1 9 1 9 9 4 4 2
40 9 1 9 1 9 9 1 9 1 13 2 9 1 9 1 13 16 12 12 12 9 9 1 9 14 1 9 1 13 2 9 9 1 13 4 4 16 4 4 2
33 9 1 13 4 4 2 9 9 9 9 9 2 1 1 12 12 12 9 1 9 1 9 13 4 2 9 9 1 9 1 13 4 2
36 9 9 1 13 16 2 9 9 9 1 9 1 12 9 9 2 9 12 12 12 12 12 12 12 9 1 9 1 13 4 4 2 9 9 2 2
19 3 9 9 1 9 9 1 2 9 1 9 9 9 9 1 3 4 4 2
21 9 1 9 1 9 9 1 13 4 16 1 12 12 12 12 9 9 12 12 9 2
23 9 12 12 9 1 9 1 2 9 9 1 1 2 9 9 9 2 1 13 4 16 4 2
17 7 2 9 1 9 9 1 12 9 9 1 12 12 9 4 4 2
62 9 1 2 9 1 9 9 2 9 9 1 13 16 9 1 13 4 9 2 1 2 9 1 13 2 1 9 1 13 16 4 16 2 9 1 2 9 9 2 1 13 9 2 2 9 9 1 9 9 2 1 13 2 9 1 9 1 13 4 1 13 2
55 11 11 5 9 9 1 2 9 9 1 9 1 9 9 1 0 2 9 1 9 9 1 9 9 14 13 4 9 1 0 2 9 1 9 1 13 4 2 9 1 9 1 13 4 16 1 1 9 1 13 2 1 13 4 2
33 9 9 9 1 9 9 1 12 12 9 1 9 12 9 1 13 2 9 1 9 1 12 9 9 1 2 3 1 9 1 13 4 2
39 9 9 1 9 9 9 9 2 11 11 9 1 2 11 1 9 9 1 13 9 1 13 16 4 4 11 1 9 1 13 4 9 2 1 9 1 13 4 2
25 7 2 11 9 1 1 9 1 9 9 1 2 9 9 9 9 9 9 2 1 13 16 4 4 2
40 9 9 1 2 9 1 13 4 9 1 0 2 1 13 16 2 9 9 1 9 1 13 4 4 9 9 9 1 2 9 1 9 9 1 13 4 2 1 13 2
32 11 1 9 9 9 1 2 11 9 1 9 1 13 16 4 1 13 2 9 9 1 13 4 16 13 4 4 2 1 13 4 2
33 11 9 1 2 9 1 0 2 15 1 13 4 4 16 13 4 4 4 1 13 9 1 9 1 0 2 1 9 1 13 4 4 2
13 0 4 9 1 9 1 1 13 4 4 16 4 2
6 9 9 12 12 9 2
33 11 5 11 1 9 9 4 2 9 1 9 7 13 4 14 3 14 1 13 4 9 9 1 9 9 9 9 9 1 13 4 4 2
35 9 9 9 1 2 11 9 9 9 1 9 9 9 2 11 5 11 1 9 2 12 12 9 2 1 0 4 13 4 4 16 13 4 4 2
24 9 1 9 2 9 9 2 9 2 11 11 9 9 1 2 9 9 1 9 9 1 13 4 2
23 2 12 12 9 2 7 2 11 9 1 11 5 11 1 2 9 2 1 9 1 13 4 2
33 2 9 2 1 12 12 12 12 12 9 1 9 9 2 2 12 12 9 2 1 12 12 12 9 1 9 9 1 13 4 4 4 2
23 9 9 4 12 12 12 12 12 12 9 1 2 12 12 9 2 14 1 9 1 13 4 2
26 7 9 2 2 9 9 1 9 9 1 9 2 14 1 13 2 9 2 1 9 9 9 1 13 4 2
12 9 1 9 1 9 2 9 9 1 13 4 2
39 9 1 9 9 1 9 1 2 2 9 1 2 9 1 9 1 13 2 1 9 1 13 4 16 4 4 9 2 1 9 9 1 9 1 13 4 4 4 2
56 7 9 11 5 9 9 9 1 2 9 1 13 16 4 4 2 1 13 2 11 9 1 2 9 1 2 9 1 13 4 16 2 15 1 13 16 2 1 9 1 13 2 13 4 9 1 9 13 16 13 4 2 1 13 4 2
67 9 1 9 5 9 1 13 9 9 1 12 9 1 2 9 9 1 10 12 9 9 1 12 12 12 12 12 9 9 1 9 1 13 4 4 14 2 12 9 1 9 1 2 9 9 9 4 1 9 1 13 2 15 9 1 10 9 1 13 16 4 4 2 1 13 4 2
27 9 1 9 9 1 2 9 2 3 9 1 9 1 13 16 1 9 4 1 9 1 13 4 2 1 13 2
36 11 9 1 2 15 1 9 14 1 13 4 16 2 0 4 9 4 4 2 9 9 1 13 4 4 16 9 9 1 13 4 2 1 13 4 2
5 9 9 1 13 2
54 2 12 12 9 9 14 2 9 9 1 9 9 1 13 4 2 15 9 12 12 9 9 1 9 1 12 12 12 12 9 1 9 1 13 4 4 4 2 9 9 1 9 3 4 13 16 4 2 9 9 1 0 4 2
19 9 1 9 9 1 9 1 13 16 2 9 9 9 1 9 1 13 4 2
22 7 2 9 1 0 9 1 13 4 9 9 1 9 7 9 1 1 9 9 1 13 2
39 9 9 12 12 12 12 12 9 2 9 9 9 12 12 12 12 9 1 0 4 9 1 13 2 3 13 4 11 9 9 9 1 9 1 1 9 1 13 2
13 9 9 1 13 9 9 2 9 1 9 13 4 2
15 9 1 12 12 12 12 12 12 12 12 12 12 12 12 2
55 11 11 5 9 9 9 1 12 9 2 9 9 1 3 12 9 13 9 1 9 9 1 13 16 2 9 9 1 9 7 9 1 13 2 9 9 1 11 9 1 13 9 9 9 9 1 13 4 9 1 0 4 13 4 2
13 11 9 9 1 9 1 9 1 9 1 13 4 2
40 9 9 9 1 11 9 1 13 4 9 1 13 4 9 4 2 10 9 1 9 1 13 9 12 9 9 9 12 9 9 1 1 0 9 1 13 1 13 4 2
65 11 9 1 2 9 9 1 0 9 1 9 9 1 1 2 12 9 9 1 0 2 9 1 2 9 7 9 1 9 9 1 13 16 9 9 13 9 1 13 16 4 2 9 1 9 1 11 9 1 13 4 2 9 0 4 9 1 15 14 0 2 1 13 4 2
50 7 11 9 1 13 16 2 9 7 11 9 1 9 1 13 4 2 11 1 9 1 13 16 2 3 13 2 11 1 13 16 4 2 1 9 9 9 1 9 1 9 9 1 13 4 4 1 13 4 2
39 11 11 5 11 9 9 9 9 9 1 2 9 14 1 9 1 0 4 9 9 1 9 1 13 9 7 9 1 9 9 9 1 0 9 1 13 4 4 2
33 9 9 9 1 9 1 9 13 9 4 2 9 9 7 9 1 9 1 0 13 2 9 9 9 1 9 1 13 1 13 4 4 2
25 9 9 1 9 7 9 1 9 1 9 1 13 4 16 4 9 1 13 4 9 1 13 4 4 2
20 9 1 1 9 2 9 2 9 2 9 2 9 2 9 14 1 9 1 13 2
20 15 1 9 9 1 0 4 0 9 1 13 2 9 9 1 0 13 16 4 2
34 9 1 12 9 1 9 9 9 1 13 4 16 12 9 9 1 9 7 9 1 9 9 1 13 16 9 1 13 9 1 13 16 4 2
28 7 2 9 1 12 9 14 13 9 9 1 9 7 9 1 9 1 9 9 1 3 0 4 13 4 4 4 2
46 9 7 9 9 9 9 1 12 12 9 9 1 12 9 9 1 9 1 9 1 0 2 9 9 2 1 13 9 1 13 4 4 16 2 12 9 9 1 9 1 13 4 4 1 13 2
14 9 9 9 1 2 9 1 9 9 1 9 1 0 2
21 9 1 3 9 7 9 1 9 1 9 1 9 1 13 16 9 9 14 1 13 2
25 9 7 9 1 9 1 13 14 13 4 9 1 9 9 9 1 13 2 9 1 9 9 1 13 2
29 7 2 0 1 9 1 9 1 9 14 1 1 13 2 9 1 9 1 9 0 4 2 9 1 0 9 1 13 2
9 9 1 12 2 12 9 1 0 2
17 9 1 9 9 1 3 4 9 1 2 9 1 9 1 13 4 2
26 3 1 2 9 9 1 13 4 9 9 9 1 9 1 2 12 12 9 9 12 9 13 4 1 13 2
59 11 9 1 2 12 9 9 1 9 1 0 9 9 1 13 4 16 2 9 9 9 1 9 1 13 2 9 1 9 9 1 13 4 9 2 9 1 2 9 1 9 1 12 12 9 14 13 16 2 9 9 1 13 2 1 13 16 4 2
28 11 9 1 0 9 1 13 4 9 9 1 9 1 9 12 12 9 1 9 11 2 11 1 3 13 4 4 2
54 9 1 9 1 13 16 4 9 9 9 9 9 1 2 9 1 0 9 1 13 16 4 2 9 9 1 9 9 1 13 9 2 9 1 9 1 2 9 1 0 4 9 1 9 1 13 16 4 2 1 13 16 4 2
18 9 9 1 13 16 1 11 9 11 9 1 9 9 2 11 11 9 2
32 11 9 1 12 12 12 12 9 2 9 1 9 11 1 13 2 9 1 3 9 11 9 1 13 16 11 1 13 4 4 4 2
12 12 12 9 9 1 9 14 9 9 1 13 2
40 9 2 9 9 1 9 2 9 1 9 1 9 1 13 2 9 1 0 9 9 7 9 9 1 13 4 9 14 12 12 12 12 9 1 13 4 4 16 4 2
22 12 12 9 9 1 2 11 14 9 12 9 1 9 9 1 13 2 9 1 13 4 2
43 9 9 2 9 9 9 9 9 1 13 4 13 4 4 11 9 9 9 9 9 9 9 9 1 11 5 11 9 1 11 9 1 13 2 2 9 1 13 9 2 1 13 2
46 9 9 9 1 11 9 1 2 9 11 1 1 2 11 9 1 9 1 13 4 4 4 2 9 11 1 1 9 9 1 2 1 13 4 2 11 9 1 12 9 1 9 1 13 4 2
83 11 9 1 9 1 13 4 9 9 1 9 1 13 11 9 1 2 9 1 9 1 9 1 13 16 2 9 1 9 1 9 7 0 9 1 13 16 4 4 2 9 1 9 7 9 1 9 1 13 16 2 9 1 13 16 4 4 2 11 1 9 1 1 2 11 1 9 1 1 2 9 1 9 1 13 16 4 2 1 13 16 4 2
43 12 9 9 12 9 12 9 9 2 9 9 9 9 1 2 9 9 9 1 9 1 13 9 9 1 9 9 9 2 9 2 1 2 9 1 13 4 4 9 1 3 9 2
24 9 1 13 4 2 9 9 9 12 12 12 9 1 9 12 12 9 2 9 9 1 13 4 2
20 9 9 1 9 9 1 13 4 2 9 1 0 9 1 9 1 13 4 4 2
58 9 1 13 4 9 9 1 2 9 1 9 1 9 9 1 9 1 13 4 9 2 9 1 13 4 4 4 9 2 9 1 0 9 1 13 4 9 9 1 13 2 9 9 1 13 4 4 12 9 1 9 1 9 1 13 16 4 2
14 9 9 2 9 9 1 9 1 13 4 16 1 3 2
26 9 13 16 4 11 9 1 1 9 1 1 2 9 1 9 1 3 0 9 1 13 4 16 4 4 2
31 9 1 13 16 9 1 1 2 3 9 9 13 4 9 9 9 1 9 9 1 13 9 1 13 4 16 4 1 1 9 2
17 9 1 9 1 13 4 4 9 1 13 4 9 1 0 9 1 2
22 2 9 1 9 1 13 16 0 4 9 1 13 16 4 2 1 11 9 1 9 9 2
12 9 9 1 1 2 9 13 9 1 2 1 2
4 9 1 9 2
11 10 9 2 9 1 1 9 1 0 1 2
26 11 9 1 9 1 13 9 9 2 9 13 2 1 12 9 2 11 9 11 9 1 9 4 13 4 2
32 9 1 9 2 12 9 9 1 9 1 2 9 2 9 1 13 4 4 5 9 2 9 9 1 0 4 9 9 1 13 4 2
62 9 1 11 9 1 11 1 13 4 4 1 13 4 2 9 2 9 9 1 9 9 9 1 9 1 12 9 12 9 1 9 1 13 2 2 6 2 2 6 2 2 6 2 1 9 9 2 9 9 12 9 1 0 9 9 1 9 1 13 13 4 2
31 11 12 9 12 9 1 9 1 9 9 9 1 9 9 9 9 4 4 9 1 12 9 2 9 9 1 9 1 13 4 2
41 9 1 9 9 1 13 4 4 9 9 9 1 9 12 9 1 13 16 4 2 9 1 2 9 9 2 1 9 9 2 11 1 3 0 4 9 1 13 4 4 2
34 9 1 13 16 2 11 1 9 1 9 9 9 1 12 12 12 12 9 1 2 12 12 12 12 9 1 12 12 12 12 9 1 13 2
12 12 12 12 12 9 1 9 9 9 2 9 2
15 11 7 11 1 9 9 4 4 12 12 9 1 13 4 2
34 11 9 11 9 9 1 12 9 9 2 11 9 9 9 2 9 2 11 11 9 9 1 9 9 9 9 9 1 9 1 13 4 4 2
34 9 1 1 2 11 9 9 1 9 2 11 9 1 9 9 9 9 1 13 2 9 12 12 9 1 1 3 9 1 13 4 4 4 2
20 7 2 11 9 9 1 9 1 1 13 4 2 9 9 1 13 4 1 13 2
28 10 9 2 11 9 1 12 9 9 2 9 1 9 1 9 1 9 9 1 13 9 9 9 1 13 4 4 2
15 11 9 9 1 11 9 1 12 9 1 13 16 4 4 2
25 12 9 9 2 11 9 9 1 2 9 1 13 16 4 2 1 9 1 11 9 9 1 13 4 2
32 9 1 13 2 13 4 4 1 13 4 16 13 16 13 4 9 2 9 1 13 2 0 13 4 2 1 13 16 4 1 13 2
75 11 9 9 9 12 1 9 9 2 11 11 9 9 1 9 9 2 9 11 9 1 9 9 1 13 4 9 1 9 1 13 4 9 1 13 4 9 1 2 9 9 1 12 9 2 13 4 16 4 4 9 9 9 1 9 9 9 2 9 9 9 2 11 11 9 9 1 9 9 9 1 13 4 4 2
11 9 1 1 2 11 9 9 1 11 9 2
34 9 9 1 9 9 12 12 9 2 11 5 11 1 13 2 9 12 12 9 1 11 1 13 2 9 14 1 13 16 4 4 1 13 2
53 11 11 9 9 1 12 9 2 9 5 11 9 1 9 9 1 13 4 2 9 1 11 11 9 9 9 1 9 1 13 4 9 9 1 13 16 2 13 4 4 9 2 9 9 1 13 4 4 2 1 13 4 2
50 11 11 9 1 12 9 9 2 9 9 1 13 4 4 9 9 1 9 9 1 13 4 2 2 9 9 1 9 1 13 16 2 9 1 9 1 13 16 13 16 4 2 1 2 9 1 9 1 13 2
65 7 2 11 11 9 9 1 9 1 13 16 13 16 4 9 1 9 9 4 13 4 2 1 13 2 9 9 5 9 9 1 9 1 13 16 9 9 1 13 9 1 1 9 1 3 13 2 9 1 9 9 9 1 13 16 1 9 1 9 9 9 1 13 4 2
68 11 9 7 11 9 1 9 1 9 1 13 16 13 4 4 16 4 11 11 9 9 9 9 1 13 16 2 9 1 13 11 9 1 9 1 13 4 2 9 9 9 9 9 9 2 1 12 9 2 9 9 1 11 9 4 12 9 9 13 9 1 9 9 4 13 4 4 2
56 7 2 11 9 1 9 1 0 9 1 1 4 9 1 2 9 9 9 1 11 9 1 9 1 13 4 2 9 1 9 1 9 9 1 9 9 1 9 1 13 16 2 12 9 1 9 1 11 9 9 1 0 9 1 13 2
32 9 1 12 12 9 1 9 1 11 9 1 9 1 13 4 4 9 1 2 0 4 9 9 13 14 13 4 14 1 13 4 2
36 11 9 1 11 2 11 1 13 4 9 9 1 13 16 1 2 9 2 1 13 16 4 2 9 9 9 1 9 9 1 13 14 3 14 0 2
70 11 9 11 9 1 9 11 5 11 11 9 1 11 9 1 12 9 13 4 4 9 4 2 11 9 1 12 9 12 9 1 13 4 9 9 4 13 4 9 1 2 11 9 1 12 9 9 12 9 12 12 12 9 1 2 11 9 7 9 9 9 9 12 12 9 1 9 1 13 2
63 9 12 12 9 9 2 9 9 1 9 12 12 9 2 0 9 12 9 1 9 1 9 1 11 9 11 9 9 12 2 9 9 2 11 11 9 7 2 13 4 16 4 4 11 9 11 9 11 12 2 9 9 2 11 11 9 1 9 1 13 4 4 2
46 10 9 1 9 1 2 9 9 1 2 9 11 2 1 9 9 1 9 2 11 11 9 1 2 9 1 13 4 12 9 1 13 4 4 11 9 9 1 9 1 9 1 13 4 4 2
29 9 1 9 9 1 9 1 13 2 12 9 1 13 4 9 1 9 1 9 1 9 1 13 16 1 0 4 9 2
21 9 1 9 9 1 13 4 9 1 2 11 9 9 12 9 1 13 16 13 4 2
46 10 9 2 9 1 9 1 13 4 2 9 9 1 9 2 1 11 9 11 9 11 12 2 9 9 2 9 9 9 9 1 12 9 1 9 1 9 1 13 16 4 1 13 16 4 2
18 7 2 9 9 1 9 1 9 1 0 2 9 1 13 4 16 4 2
35 11 9 1 2 9 1 9 11 5 11 9 1 13 4 4 9 1 9 1 2 12 9 9 13 4 9 1 13 9 9 1 13 16 4 2
29 9 9 1 2 9 9 2 9 9 1 9 1 13 16 13 9 9 1 0 9 1 0 2 1 13 4 16 4 2
30 2 9 1 11 9 1 13 16 1 9 9 1 9 2 7 2 9 2 9 9 9 1 9 9 4 9 1 9 2 2
22 9 9 9 1 11 9 9 1 13 16 2 9 9 9 9 1 10 9 1 13 4 2
26 12 9 14 1 9 1 13 4 4 2 9 9 9 1 9 9 1 13 16 2 1 0 4 13 4 2
18 15 1 13 16 2 9 9 9 1 9 9 1 9 1 13 16 4 2
44 7 2 9 1 9 1 0 9 1 13 4 9 1 9 9 9 1 13 9 9 1 9 1 9 2 1 2 3 9 9 9 1 13 9 1 1 4 9 1 13 4 16 4 2
28 9 5 9 9 9 1 11 9 9 1 9 1 9 1 3 9 9 4 13 9 4 2 9 1 13 4 4 2
22 9 1 9 1 13 4 2 9 9 2 1 10 12 9 14 9 9 1 13 16 13 2
15 9 9 1 9 9 1 0 4 9 9 1 13 16 4 2
34 7 9 11 1 13 4 16 4 11 1 9 9 9 9 1 9 2 12 9 9 1 9 12 12 12 12 12 12 9 1 13 4 4 2
15 2 9 9 4 1 4 16 9 9 1 9 2 1 13 2
22 0 9 1 2 9 1 9 9 1 9 9 2 9 9 9 1 13 16 9 1 13 2
56 9 9 9 1 2 12 2 9 1 3 9 2 12 2 9 9 9 9 9 2 9 2 1 13 2 11 9 1 3 13 2 12 2 9 1 9 2 9 2 13 2 9 9 1 13 2 13 9 14 1 9 1 13 16 13 2
21 2 9 9 9 1 9 9 1 13 16 2 1 13 4 9 9 1 13 4 4 2
22 15 1 13 16 2 9 9 4 15 1 9 1 9 9 9 1 9 1 13 4 4 2
53 9 9 12 12 9 2 9 1 9 1 13 4 9 1 13 4 9 1 9 9 1 9 2 2 9 9 9 9 12 9 2 9 9 1 9 9 1 13 4 9 2 9 9 7 9 9 1 13 2 1 9 4 2
17 7 2 9 9 1 9 1 9 9 1 3 13 4 16 4 4 2
19 7 9 1 13 9 1 9 9 14 1 13 4 16 4 4 16 1 9 2
48 9 9 1 1 2 2 9 9 1 1 9 5 9 1 9 9 1 13 2 11 1 9 2 9 9 9 9 1 9 2 9 1 0 9 9 1 13 4 2 9 1 9 1 9 1 13 4 2
74 10 9 1 13 16 11 1 2 9 9 1 9 9 1 9 1 13 16 1 12 9 4 16 2 9 9 1 13 16 1 9 9 1 13 1 1 9 1 13 16 4 2 1 13 16 1 2 7 9 9 1 3 13 4 9 1 2 9 2 9 9 4 9 1 13 16 4 4 2 1 13 16 4 2
13 11 1 9 1 0 2 15 1 3 13 16 4 2
10 11 1 4 4 9 1 13 4 4 2
18 11 1 1 3 9 1 13 9 9 1 9 9 1 9 4 16 4 2
27 11 1 9 1 13 16 1 2 9 9 1 13 4 2 0 9 1 9 14 4 2 1 13 9 4 4 2
34 7 9 2 12 9 1 9 1 2 9 9 1 0 9 1 1 9 9 4 2 11 9 1 9 9 1 9 7 9 1 9 4 4 2
25 9 12 9 9 1 3 13 4 16 4 4 11 1 1 0 4 9 4 4 9 1 13 1 4 2
17 7 2 10 9 9 1 9 1 9 14 9 14 1 9 1 13 2
32 9 1 2 9 9 1 13 2 9 9 1 13 16 1 2 3 9 1 13 4 2 1 9 9 1 9 1 9 1 0 4 2
31 3 9 1 9 12 12 12 9 1 9 9 1 9 1 13 2 0 9 1 2 9 1 9 2 1 13 9 1 13 4 2
32 11 1 1 2 9 7 9 1 9 1 13 2 1 3 13 4 16 2 9 1 2 9 1 9 1 13 2 1 13 9 4 2
12 9 9 1 9 1 9 4 16 14 13 4 2
47 11 9 1 13 16 9 2 12 12 9 9 1 9 9 12 9 1 9 1 9 1 13 4 9 2 2 9 1 9 1 0 4 2 1 13 4 4 9 1 12 12 9 1 1 13 4 2
20 3 12 12 9 1 2 9 9 1 9 5 9 1 2 1 13 4 1 13 2
31 9 1 9 2 9 9 1 0 9 1 13 2 1 13 4 16 4 16 2 9 1 9 5 9 1 13 4 4 9 4 2
15 7 9 9 13 4 4 16 1 9 9 1 9 9 4 2
64 0 4 9 4 16 2 0 9 9 1 2 9 1 9 9 14 1 13 16 4 9 1 9 1 9 4 2 1 13 16 12 9 1 13 16 4 16 14 2 9 1 2 9 1 13 16 2 9 9 2 1 13 16 2 13 4 16 4 2 1 9 9 4 2
16 7 9 2 9 9 1 9 1 13 4 9 9 1 13 4 2
26 9 9 1 9 9 13 2 9 12 9 9 1 11 5 11 9 1 2 12 12 9 13 9 1 9 2
29 9 9 1 9 1 13 16 9 7 9 1 9 1 13 4 2 9 1 9 1 13 16 1 9 1 13 16 4 2
26 9 9 1 2 9 9 2 1 9 9 1 0 9 1 13 16 14 2 3 0 9 1 0 4 4 2
27 9 1 9 2 9 9 1 9 1 13 4 2 12 9 1 12 12 9 1 9 1 13 4 2 9 2 2
17 9 9 14 13 16 2 9 1 0 4 9 1 13 4 4 4 2
16 9 1 9 1 13 4 16 1 2 9 9 1 9 1 9 2
29 10 9 1 9 9 1 9 1 13 2 2 9 1 13 4 9 9 9 1 2 9 1 13 16 4 4 1 13 2
21 13 4 16 9 1 1 13 4 9 14 1 2 9 1 1 9 1 3 13 4 2
25 9 1 9 9 1 9 1 13 16 2 9 9 1 1 2 9 2 1 9 9 1 13 16 4 2
11 9 1 9 9 1 3 13 4 9 9 2
26 10 9 9 1 0 4 13 2 9 1 13 4 4 4 9 1 13 4 16 4 16 1 9 1 13 2
27 9 1 12 9 1 9 9 14 1 2 3 9 1 13 16 1 13 4 1 13 9 1 0 2 4 4 2
4 9 1 9 2
20 7 2 2 12 12 9 9 1 9 1 9 1 9 1 13 4 4 14 2 2
39 9 1 13 4 9 2 9 1 13 9 5 5 6 2 1 13 4 4 9 1 9 2 2 9 9 2 2 9 9 9 2 1 13 9 1 13 4 4 2
22 0 9 1 13 16 9 9 1 13 9 1 9 0 2 9 1 10 9 1 13 4 2
19 7 2 9 12 9 5 9 1 13 2 13 2 2 1 13 16 4 4 2
10 13 9 4 9 1 9 1 13 4 2
34 13 16 4 9 1 13 4 9 1 1 4 2 9 1 13 16 2 9 9 1 9 9 9 1 13 16 9 1 3 4 13 16 4 2
21 9 1 2 9 9 2 1 2 13 4 4 16 1 9 9 1 9 9 9 9 2
33 11 9 9 1 9 1 13 9 2 9 0 1 9 9 1 13 9 1 13 16 4 2 9 1 14 9 1 3 1 1 13 0 2
34 9 1 13 16 1 13 9 1 0 2 9 1 2 13 16 4 16 13 9 1 13 2 1 13 9 1 9 9 1 13 4 1 13 2
10 13 9 1 13 16 2 13 9 1 2
19 9 9 9 1 11 5 9 11 1 13 4 4 2 9 1 13 9 2 2
32 3 9 1 9 4 16 4 16 2 9 1 13 16 9 1 9 1 13 9 1 9 2 13 16 3 2 9 9 2 1 13 2
27 9 1 9 12 12 9 9 1 9 9 1 2 9 1 9 2 9 1 9 1 13 4 4 2 1 13 2
22 13 16 1 13 4 9 2 9 9 2 1 9 9 1 13 16 1 9 9 1 11 2
19 15 14 0 9 1 9 9 1 1 2 15 14 1 13 16 9 4 4 2
29 10 9 2 9 1 12 12 9 13 4 4 9 2 9 1 13 4 9 9 1 9 9 1 9 1 13 1 13 2
60 9 1 2 2 9 9 2 1 9 2 9 1 9 9 1 13 2 2 9 9 5 9 9 1 13 2 1 9 1 13 4 9 2 9 9 12 2 2 9 9 7 9 9 1 13 4 4 9 2 9 9 2 1 9 9 9 1 9 9 2
19 9 9 1 1 9 9 4 4 9 9 9 1 9 1 9 9 1 13 2
28 9 9 1 1 2 11 9 9 1 2 9 1 9 9 2 9 1 9 2 1 9 1 9 9 1 13 4 2
14 9 1 9 1 9 1 13 16 4 16 2 3 0 2
25 9 1 9 1 9 9 1 13 16 1 9 4 16 2 2 9 9 1 9 2 9 1 13 4 2
15 11 9 11 9 11 1 1 9 1 13 4 9 1 13 2
19 9 11 9 9 1 9 9 1 9 1 13 0 9 12 12 9 1 9 2
18 9 1 13 4 2 9 9 9 9 9 9 14 13 4 4 16 4 2
7 7 2 9 9 1 0 2
35 1 13 16 1 2 2 9 1 9 4 4 2 9 9 1 9 2 4 16 4 2 9 1 13 16 2 9 2 9 2 9 14 1 13 2
16 9 13 9 11 9 9 9 1 12 9 1 9 1 13 4 2
23 9 9 1 9 9 1 2 13 4 9 1 13 16 12 12 12 12 12 9 9 1 13 2
8 9 9 1 9 9 1 13 2
14 9 1 13 4 16 4 9 5 9 12 12 12 9 2
21 9 9 1 1 13 4 2 9 1 9 9 12 12 9 9 1 9 1 13 4 2
24 9 1 2 9 1 9 1 13 16 4 16 0 16 2 3 4 4 16 9 1 9 1 0 2
18 7 9 1 13 9 2 9 9 1 9 14 1 13 0 9 1 13 2
23 2 0 9 1 0 4 2 9 9 1 13 9 1 13 4 9 1 1 13 2 1 9 2
39 0 9 1 13 16 1 2 6 2 1 9 4 16 2 9 9 1 13 9 1 2 10 9 1 9 9 1 9 1 13 4 9 1 13 16 4 4 4 2
73 12 9 9 1 9 9 9 9 11 5 9 1 13 16 2 9 11 9 9 1 10 9 13 4 11 1 9 9 1 13 9 9 1 9 1 2 11 9 1 0 9 9 1 9 1 9 1 13 4 4 1 9 2 9 9 1 0 9 1 13 9 1 13 4 0 9 1 13 1 13 16 4 2
53 9 1 13 16 2 9 9 1 2 11 9 1 9 9 1 13 4 16 4 4 2 1 13 2 9 9 1 0 9 9 1 2 9 9 2 1 13 2 9 1 11 1 1 9 1 13 4 4 1 13 16 4 2
12 11 9 9 9 9 1 9 1 13 16 4 2
54 9 9 1 9 9 1 12 9 2 13 4 4 9 1 11 9 1 2 11 5 11 9 9 1 3 2 9 2 1 13 4 9 1 2 9 1 9 1 9 1 9 1 0 4 13 2 7 9 9 1 13 4 4 2
65 7 2 10 9 1 9 1 2 15 14 1 9 1 13 16 13 16 4 2 1 13 9 1 13 16 2 9 2 13 4 9 4 2 11 9 1 2 9 1 13 4 9 2 9 1 13 4 16 1 0 4 9 2 1 9 4 9 1 9 1 13 4 16 4 2
38 15 1 2 11 9 1 9 9 9 2 11 5 11 9 1 2 11 9 1 9 11 9 1 9 1 12 9 1 13 16 13 4 4 9 1 14 9 2
21 9 1 12 9 1 9 4 16 2 11 1 12 9 2 9 9 1 13 4 4 2
37 15 1 13 16 2 11 9 1 9 9 1 3 13 4 16 4 4 14 13 4 4 11 9 1 2 11 9 1 9 2 13 4 4 2 1 13 2
39 11 9 1 2 15 14 1 9 4 3 13 16 4 4 4 14 2 1 13 16 13 16 2 15 1 9 4 2 1 13 16 4 4 14 2 1 13 4 2
20 15 1 13 4 11 1 2 0 4 9 4 2 13 4 16 4 2 1 13 2
64 0 9 1 2 15 14 1 9 4 2 1 13 16 1 9 4 13 16 4 1 13 9 4 2 0 4 9 1 2 9 13 4 16 4 4 15 1 9 1 0 13 9 1 13 16 1 0 4 1 4 14 2 1 13 2 11 9 1 9 1 13 16 4 2
32 15 1 13 2 11 9 1 2 10 9 1 13 16 1 0 4 1 4 1 13 2 1 13 16 2 9 9 13 4 9 4 2
44 9 1 12 12 9 9 1 9 9 1 13 4 4 9 9 12 12 12 9 1 12 9 2 13 4 2 9 1 1 9 1 9 5 11 9 1 0 4 9 1 13 4 4 2
47 9 1 9 9 9 1 9 2 9 9 9 1 9 9 14 2 9 1 9 1 9 9 9 1 9 1 13 2 9 1 9 1 13 13 16 4 4 9 1 9 9 1 0 9 1 13 2
20 9 9 1 9 9 1 13 4 9 9 1 9 9 9 9 1 0 13 4 2
72 11 9 9 1 12 12 12 12 9 9 2 1 13 9 1 1 9 1 13 4 4 9 1 2 9 9 1 9 9 1 9 1 12 12 12 9 1 2 9 9 12 9 1 13 9 1 3 1 13 4 4 2 1 13 9 9 2 9 1 2 9 14 1 13 9 1 9 5 9 1 13 2
16 9 9 1 13 4 4 9 1 9 9 1 9 1 13 4 2
66 0 4 9 9 1 2 12 9 9 9 7 12 12 12 9 9 9 1 9 7 2 9 9 1 12 9 12 9 2 9 9 9 1 9 12 9 9 9 2 9 9 1 9 2 9 9 9 1 1 15 14 1 9 1 12 9 12 1 9 1 9 1 13 9 14 2
31 7 2 9 9 1 13 16 4 9 9 9 14 9 9 9 1 9 1 9 9 1 9 1 1 13 4 9 1 13 4 2
77 11 9 9 1 9 9 1 2 9 1 11 1 9 9 1 13 16 4 4 0 4 9 9 9 1 9 9 4 4 2 10 9 1 9 9 1 13 4 16 1 9 1 9 9 4 4 2 9 1 9 1 9 1 9 1 13 4 4 2 1 13 2 12 12 9 1 9 1 9 1 9 1 9 1 13 4 2
53 7 2 10 9 1 9 9 1 12 12 9 1 2 11 9 2 1 9 1 3 13 9 9 1 13 2 15 1 11 1 2 9 9 1 13 9 1 9 1 9 1 13 9 1 13 4 16 4 4 2 1 13 2
14 9 9 1 9 9 1 9 1 0 9 1 13 4 2
27 7 2 9 1 9 9 4 9 1 13 4 9 9 9 9 1 11 5 9 9 9 9 1 13 4 4 2
10 9 1 9 9 1 12 12 9 9 2
13 11 9 1 2 9 1 9 9 9 9 4 4 2
19 9 9 1 9 9 1 2 9 1 9 12 12 12 2 9 12 12 12 2
22 9 1 9 12 12 12 12 2 9 12 12 12 2 9 9 1 12 1 13 16 4 2
46 11 9 9 1 9 11 1 9 1 13 4 4 9 1 9 1 13 16 4 4 11 9 1 2 11 9 1 9 1 13 16 12 9 9 12 9 1 9 9 1 13 4 4 9 4 2
8 9 1 1 9 9 1 0 2
49 9 9 9 1 13 16 2 9 9 1 12 9 2 9 1 9 9 2 9 9 1 11 9 1 9 1 13 4 9 2 9 9 1 9 1 13 4 9 1 13 4 16 13 4 4 4 1 13 2
55 9 9 1 9 12 12 12 9 2 0 9 1 9 9 1 9 1 13 4 4 16 2 9 1 0 9 1 13 4 2 3 9 1 9 1 13 16 1 9 9 9 1 1 11 9 1 13 9 1 9 9 1 13 4 2
39 11 9 9 9 9 1 12 9 1 9 1 2 11 5 9 1 9 9 1 13 2 9 9 9 9 1 0 9 1 13 4 9 1 9 1 13 4 4 2
30 11 1 9 1 1 11 9 1 1 9 1 0 4 9 2 9 9 1 9 1 13 4 9 1 13 16 4 1 13 2
49 9 9 9 1 13 16 2 9 9 1 13 4 16 9 9 9 9 1 13 16 4 11 9 1 2 9 12 9 1 13 16 1 2 9 12 12 12 9 9 1 9 9 1 13 4 16 4 4 2
49 9 1 13 4 16 1 2 11 2 11 9 2 11 2 11 1 12 9 1 2 9 9 9 9 12 12 12 9 1 9 9 9 9 2 9 5 9 5 11 14 1 13 4 4 13 4 16 4 2
37 9 9 1 12 9 2 11 9 9 1 12 9 1 12 12 9 14 11 2 11 2 11 2 11 1 12 9 1 13 4 9 1 0 4 13 4 2
23 9 9 9 1 11 2 11 9 9 1 2 12 12 12 12 9 1 11 9 9 1 13 2
23 11 2 11 9 1 1 9 9 1 9 1 1 9 9 9 5 9 9 1 13 9 4 2
48 11 9 1 11 9 1 13 16 11 9 1 9 1 2 11 9 1 9 9 7 11 1 13 4 16 4 9 9 9 9 1 9 1 13 16 9 1 9 9 1 13 9 1 13 16 4 4 2
20 9 9 9 9 9 1 11 7 9 1 9 1 3 9 9 13 9 1 13 2
39 9 9 9 1 13 16 2 11 9 1 9 9 4 4 11 1 11 9 1 12 9 2 9 9 1 13 16 11 1 11 1 13 4 9 1 13 4 4 2
62 10 9 1 13 16 2 11 1 11 9 9 1 13 4 4 9 1 1 2 9 9 1 1 9 9 1 9 1 13 4 2 9 1 13 9 5 9 9 1 9 9 2 1 13 16 4 9 2 11 1 11 1 9 1 13 4 9 1 13 4 4 2
73 9 9 1 12 9 2 12 12 12 12 9 1 9 9 9 9 1 2 9 1 1 12 12 12 12 9 13 4 16 9 9 1 12 12 12 12 12 12 9 1 13 2 9 9 1 12 9 9 9 1 2 9 9 1 12 12 12 12 12 12 9 1 9 1 13 1 1 9 1 13 4 4 2
31 10 9 2 9 9 9 1 13 9 9 1 9 1 12 12 9 1 12 12 9 1 12 12 9 1 1 13 4 1 13 2
81 11 9 9 9 9 9 1 12 9 2 9 9 9 9 9 1 9 9 9 9 1 13 16 9 9 13 2 9 9 1 9 9 1 9 13 16 4 4 2 15 1 9 13 9 1 13 4 16 4 2 1 13 16 1 2 9 9 1 9 1 9 9 12 12 12 9 1 13 9 1 1 4 1 1 9 1 0 4 13 4 2
25 11 9 1 9 9 1 13 2 9 9 1 13 9 1 13 4 9 1 9 1 13 16 4 4 2
46 11 9 1 7 2 9 9 9 9 1 13 2 2 9 9 2 11 5 9 9 9 9 2 9 9 14 1 9 1 13 2 9 9 1 3 9 1 9 1 13 4 2 1 13 4 2
16 9 11 9 2 9 9 9 9 9 2 1 13 4 4 4 2
30 2 9 2 1 12 12 12 12 9 9 2 9 9 1 9 9 1 9 1 11 9 9 1 13 4 16 13 4 4 2
39 9 0 9 1 1 12 12 12 9 0 9 7 10 9 9 1 13 4 2 11 11 9 9 9 9 12 9 13 12 12 9 1 9 1 13 4 4 4 2
38 9 1 11 1 13 4 9 2 12 12 9 1 11 9 9 1 13 2 12 12 9 1 13 4 4 4 9 1 9 1 9 9 14 1 13 16 4 2
49 10 2 9 2 1 2 9 2 1 9 1 9 9 2 9 7 9 14 9 9 1 9 2 9 1 1 9 2 9 1 9 14 1 13 16 2 13 9 9 4 9 1 13 16 13 4 16 4 2
21 9 13 4 4 16 4 4 9 1 9 7 9 14 1 0 4 13 4 16 4 2
12 9 1 1 9 7 9 9 1 13 16 4 2
39 9 1 9 9 1 9 1 13 16 13 4 16 4 4 9 9 2 11 9 9 2 1 10 9 13 4 4 4 9 12 12 12 9 1 9 1 13 4 2
35 12 12 12 12 9 1 13 4 4 4 9 1 2 9 5 9 1 9 9 1 13 4 2 9 9 9 14 1 13 4 4 16 4 4 2
33 9 2 9 1 9 9 9 1 13 4 4 16 4 16 2 9 1 0 4 9 1 1 4 4 16 2 10 9 1 13 16 4 2
16 9 1 0 9 1 0 4 14 1 9 1 13 9 1 0 2
10 9 1 2 9 9 4 9 1 13 2
62 9 1 13 4 9 1 1 2 11 9 1 0 4 9 9 1 13 2 9 1 9 1 3 1 0 9 1 13 4 16 4 4 2 9 1 13 4 16 1 2 9 9 5 9 9 9 2 1 13 14 0 1 9 1 13 16 4 4 2 1 13 2
19 9 9 1 2 9 11 2 1 1 2 9 1 4 4 13 4 16 4 2
79 2 9 9 1 13 9 2 11 12 9 1 13 4 1 13 16 4 2 10 9 1 3 2 11 9 9 2 9 9 1 9 1 13 4 2 9 1 13 16 1 2 0 9 1 9 1 13 9 1 2 0 9 1 1 13 2 3 0 9 4 4 4 2 3 9 1 13 4 9 9 1 0 9 1 13 4 4 4 2
29 2 9 12 9 9 5 9 2 1 2 9 12 9 1 12 12 9 14 2 9 1 9 2 11 1 13 4 4 2
66 9 9 1 2 11 11 9 9 2 1 9 2 2 9 1 9 9 2 2 2 9 2 14 9 1 1 3 9 9 1 9 7 2 11 9 2 11 2 11 2 11 14 9 1 9 1 9 1 2 9 1 9 1 13 4 4 0 9 1 9 1 13 4 16 4 2
29 7 2 9 1 12 9 1 12 9 13 4 2 9 9 2 1 13 2 11 1 9 9 9 1 10 9 1 13 2
17 9 1 9 9 1 13 4 4 9 5 9 1 9 9 1 9 2
10 11 9 11 1 9 1 13 4 4 2
32 9 9 1 13 4 9 1 13 4 4 2 3 0 4 1 9 1 13 4 16 4 4 16 2 9 9 1 11 9 1 13 2
36 10 9 2 9 1 9 4 2 13 4 9 1 1 12 12 5 12 12 9 2 9 1 13 16 12 9 2 12 9 1 9 9 13 16 4 2
12 13 16 1 12 2 12 9 1 9 9 14 2
45 9 9 1 13 4 4 12 12 9 1 9 1 2 9 0 13 4 2 7 9 1 0 4 9 14 2 9 1 13 9 1 13 9 9 1 13 4 2 9 1 13 4 9 4 2
30 9 1 1 2 12 12 9 9 1 9 1 13 4 16 4 2 9 1 9 1 1 9 13 4 2 1 13 16 4 2
8 9 1 9 1 4 4 9 2
10 9 1 9 1 3 0 9 1 9 2
23 9 1 9 7 9 1 13 2 9 1 13 2 13 13 4 9 1 13 16 9 1 13 2
9 9 1 11 9 1 11 9 9 2
18 11 1 12 12 5 12 12 12 9 1 9 2 9 1 12 9 9 2
29 9 1 3 2 9 9 1 13 16 4 16 2 9 1 3 14 2 9 1 12 12 12 9 14 1 9 1 13 2
18 9 12 9 1 9 1 13 2 10 9 14 13 16 2 0 4 13 2
29 9 1 2 9 9 1 13 2 9 1 13 4 16 13 16 4 16 2 15 1 1 2 3 13 4 9 1 0 2
21 9 9 1 3 2 9 13 4 2 13 4 1 2 14 9 13 16 1 3 13 2
22 9 1 11 9 1 2 9 2 9 12 12 12 12 12 12 12 12 12 12 12 12 2
25 9 12 9 9 12 12 12 12 9 2 12 9 12 12 12 12 9 2 9 9 12 12 12 9 2
8 11 1 13 16 2 11 9 2
48 10 9 1 9 1 9 1 13 4 4 16 2 9 9 5 9 1 11 9 1 2 11 1 0 1 9 9 1 13 4 16 4 4 9 9 9 1 2 11 9 9 9 2 1 13 4 4 2
21 9 9 9 1 9 1 9 12 9 9 1 9 1 13 2 3 9 1 13 4 2
38 9 1 1 11 9 2 9 2 9 2 9 11 9 14 1 13 4 2 9 1 9 2 9 9 1 9 2 9 9 9 1 13 4 12 9 1 13 2
17 9 1 9 1 13 2 9 1 9 1 13 4 0 9 1 0 2
18 9 9 9 7 9 9 14 1 9 9 1 9 13 4 16 4 4 2
22 9 9 12 9 13 12 12 12 12 9 2 0 9 12 9 13 12 12 12 12 9 2
14 9 12 12 12 12 12 12 12 12 12 12 12 12 2
26 11 1 9 11 1 9 9 1 13 4 9 9 1 9 2 9 1 9 2 1 1 13 4 16 4 2
29 10 9 1 13 9 1 0 9 11 1 11 1 13 16 2 12 12 1 1 9 9 1 13 4 16 4 16 4 2
39 9 1 13 4 4 2 9 2 1 13 16 4 2 9 1 9 1 13 16 4 4 4 9 9 1 9 1 9 9 1 9 9 7 2 9 9 1 13 2
44 10 9 1 9 1 9 1 0 4 13 4 16 1 2 12 12 9 1 9 2 9 5 11 9 1 9 9 1 9 1 2 11 1 11 1 9 9 1 13 4 9 1 13 2
32 0 1 13 4 9 1 9 1 2 9 1 13 9 1 9 1 13 0 4 9 1 13 16 2 9 9 1 9 1 13 4 2
29 0 9 9 1 9 1 2 2 11 2 2 11 2 2 9 2 1 13 4 9 1 3 9 1 13 4 16 4 2
10 11 1 12 12 12 12 9 1 9 2
33 9 9 1 11 1 13 4 11 9 9 9 1 9 9 1 1 2 11 9 1 9 1 12 12 12 12 9 1 13 4 16 4 2
26 10 9 1 13 4 4 11 5 11 9 1 9 2 11 1 1 2 9 1 12 9 1 9 1 13 2
41 10 9 12 9 1 12 12 9 1 13 4 14 4 16 2 9 1 11 2 11 1 13 4 9 9 1 9 1 13 4 14 2 9 1 13 4 4 9 9 14 2
29 11 1 9 2 9 1 9 1 1 9 1 9 13 1 13 4 2 9 9 1 9 9 1 13 4 9 1 13 2
33 13 4 9 1 13 1 2 9 9 14 2 0 4 9 1 9 1 13 16 4 9 1 2 15 14 13 16 4 16 1 13 4 2
39 11 1 1 2 9 7 9 1 9 1 13 16 4 2 9 1 9 1 9 1 9 1 9 1 13 7 2 13 4 14 1 9 1 0 4 9 1 13 2
40 9 1 3 1 2 3 1 13 4 9 9 1 9 1 1 9 9 1 9 1 13 4 9 7 2 9 1 13 9 9 1 9 1 9 1 13 4 16 4 2
31 9 9 1 9 9 2 9 2 9 9 14 2 9 1 13 4 9 1 13 4 1 13 9 1 3 9 1 13 16 4 2
18 12 12 12 12 9 1 13 4 4 4 11 1 2 11 9 1 9 2
17 12 12 9 1 13 9 9 1 2 9 2 9 1 13 16 4 2
23 10 9 1 1 15 14 1 9 1 9 9 1 13 2 0 4 9 1 13 4 16 4 2
44 9 9 1 9 1 13 4 9 9 1 13 14 2 9 9 9 9 0 1 9 1 13 16 4 2 9 1 9 1 2 9 9 1 1 13 9 1 13 16 4 16 1 0 2
45 2 9 1 9 2 1 13 1 1 2 11 1 11 1 13 9 1 13 16 2 9 9 13 16 1 0 16 2 9 1 9 1 13 16 9 1 13 4 9 1 0 14 13 4 2
24 0 9 1 13 16 1 9 1 13 4 16 2 9 1 9 9 1 13 16 4 16 1 0 2
16 11 1 11 14 1 9 1 9 12 9 9 1 9 1 13 2
38 9 12 12 9 9 9 2 9 2 1 1 2 0 4 9 1 9 1 9 9 7 9 1 13 4 9 9 1 9 9 9 2 9 9 2 1 13 2
9 12 12 9 5 12 12 9 9 2
28 9 2 9 1 9 1 9 9 7 9 9 9 1 9 9 9 2 9 12 9 9 9 9 14 1 9 1 2
18 9 12 12 12 12 12 12 12 12 12 12 12 12 5 9 9 9 2
15 0 4 9 5 9 1 9 1 9 9 1 9 1 13 2
7 3 9 1 2 11 2 2
15 9 5 9 1 9 1 1 9 1 9 1 13 11 9 2
10 9 1 9 1 13 9 1 13 4 2
19 9 1 11 11 2 11 11 9 1 9 2 11 11 9 1 9 1 13 2
7 9 1 9 1 11 11 2
11 11 9 9 1 9 9 1 2 11 2 2
18 9 2 9 1 9 9 4 11 1 13 2 3 9 9 1 13 4 2
43 12 9 9 1 9 1 2 12 12 12 12 9 1 9 9 13 4 9 5 9 1 2 12 12 9 1 13 4 4 4 11 11 1 9 9 9 13 16 1 9 5 9 2
19 11 9 1 9 1 2 12 12 9 1 9 1 2 11 2 1 11 9 2
15 11 7 11 1 1 9 1 13 4 9 1 13 9 4 2
25 12 12 9 1 11 9 1 1 2 0 4 9 7 0 4 9 1 13 9 1 9 1 13 4 2
29 11 9 1 11 1 9 9 1 11 5 9 7 11 11 2 9 9 1 11 1 11 5 9 7 11 11 1 9 2
6 9 9 1 11 9 2
5 9 1 11 11 2
11 7 9 1 1 11 9 9 1 13 4 2
37 12 12 12 12 9 1 13 4 4 2 11 1 2 11 5 11 2 1 13 2 11 9 1 9 1 13 4 4 9 1 13 9 1 9 9 4 2
25 9 1 10 2 11 5 11 2 7 2 3 10 9 1 9 9 1 13 4 2 11 1 9 2 2
26 9 9 4 0 4 9 1 13 9 1 1 4 16 2 9 1 9 1 13 16 4 14 1 13 4 2
5 9 9 11 9 2
17 9 9 1 9 1 13 16 12 12 12 9 9 1 9 6 4 2
49 9 1 9 9 11 11 9 1 9 1 2 9 0 9 2 9 9 2 9 1 9 7 10 9 1 11 2 9 1 11 1 9 1 13 7 2 7 9 1 13 7 1 9 1 13 16 4 4 2
15 11 9 1 9 1 9 1 2 9 1 13 16 4 4 2
23 11 9 1 9 1 13 9 1 0 4 9 1 13 16 4 16 1 2 3 1 9 4 2
36 9 1 9 9 9 1 9 1 9 1 9 1 13 2 15 1 9 1 13 4 4 16 2 15 1 13 1 13 4 9 1 9 1 13 4 2
26 11 1 13 16 4 4 9 1 13 4 4 11 9 1 2 11 1 11 1 9 1 9 1 13 4 2
18 7 11 9 1 9 1 13 4 9 1 9 1 13 4 1 13 4 2
21 3 0 13 4 11 9 4 16 2 9 9 14 1 9 9 13 4 7 13 4 2
15 9 1 13 4 4 4 11 9 14 2 1 13 9 4 2
7 7 2 3 4 4 14 2
22 11 9 9 1 9 1 2 11 9 1 9 13 16 13 4 14 1 1 4 4 4 2
13 9 1 2 3 9 0 4 4 9 1 9 4 2
11 7 2 9 1 13 4 4 16 4 4 2
25 9 4 4 11 1 2 9 1 9 1 13 4 2 11 1 9 1 9 1 13 16 9 13 4 2
23 10 9 14 1 9 1 13 16 4 4 11 1 2 3 9 1 13 7 13 16 4 4 2
40 15 1 2 3 9 9 1 11 9 7 11 1 13 16 4 4 4 13 16 2 2 6 2 3 3 13 4 16 14 2 1 13 9 1 13 16 4 16 4 2
23 11 9 1 0 9 1 2 15 1 13 9 4 2 0 4 9 1 13 16 4 9 4 2
27 11 9 1 11 1 9 1 9 1 13 4 9 1 2 9 1 9 1 13 16 4 4 9 1 13 4 2
21 10 9 1 11 11 1 9 1 13 16 2 15 14 1 3 1 13 16 4 4 2
17 9 14 11 1 0 9 1 9 1 9 1 13 16 1 13 4 2
15 11 9 1 9 1 13 16 1 13 4 16 4 4 14 2
20 9 1 9 1 13 4 2 11 1 13 4 16 9 1 13 14 13 16 4 2
25 11 2 11 2 11 1 2 9 1 1 9 1 0 4 9 1 9 2 9 9 13 4 4 9 2
21 9 9 2 13 13 2 1 0 4 2 10 9 0 4 9 1 13 16 4 4 2
38 9 1 2 9 9 1 3 9 5 9 13 4 2 9 13 4 4 11 9 2 9 5 9 2 1 9 5 9 9 1 9 1 9 1 13 4 4 2
41 2 9 1 9 2 9 9 1 2 3 2 9 2 1 13 4 4 2 9 2 9 12 9 2 2 12 9 2 1 13 16 4 4 2 1 9 1 3 0 4 2
39 2 9 9 1 9 2 1 13 4 9 1 9 1 2 9 14 1 12 12 9 2 12 12 12 9 1 13 2 9 9 1 10 9 9 1 13 4 4 2
63 2 11 1 0 9 1 13 4 16 1 9 1 9 1 9 1 13 16 4 2 7 2 9 9 1 11 1 13 16 9 1 3 0 9 1 13 4 4 2 1 13 9 1 9 1 2 9 1 9 9 1 2 9 1 9 7 9 1 0 4 13 4 2
22 11 1 1 2 11 5 11 4 1 12 9 14 13 4 4 9 1 12 9 1 9 2
28 9 9 1 2 9 9 9 1 9 1 13 16 4 4 9 1 2 9 1 9 1 13 16 9 1 13 4 2
19 9 9 1 3 2 9 1 13 4 4 9 1 9 1 9 14 13 4 2
19 11 1 1 2 9 1 9 1 9 1 13 2 9 9 1 13 4 14 2
60 2 9 1 9 1 0 9 1 9 1 13 16 13 4 16 2 9 9 2 0 9 1 13 4 2 1 13 9 1 2 9 9 1 13 16 2 9 1 9 9 13 4 16 4 16 2 9 14 1 9 9 13 9 1 2 9 9 4 4 2
19 10 9 1 2 3 9 9 4 13 4 16 1 2 9 1 9 9 4 2
64 2 9 5 9 9 2 9 9 1 3 1 9 4 4 16 2 9 7 9 1 13 16 1 2 9 1 3 13 1 13 4 4 2 7 2 3 9 1 9 1 13 16 13 4 9 1 1 4 2 1 9 9 2 9 5 9 2 1 9 9 13 4 11 2
16 9 1 2 3 9 9 4 9 1 13 4 4 9 5 9 2
9 9 1 3 9 1 13 9 4 2
75 9 9 1 11 5 11 1 13 16 2 15 14 11 1 9 1 9 1 3 13 16 4 4 16 2 9 1 9 1 13 16 3 9 1 13 4 9 4 1 13 4 2 13 4 4 9 9 1 9 1 13 4 9 2 13 4 9 1 9 4 4 16 4 2 9 1 13 4 4 2 1 9 1 13 2
37 9 1 9 1 0 4 9 1 2 9 2 12 9 1 13 4 16 2 9 1 13 16 1 9 1 9 2 9 1 9 1 13 16 4 9 4 2
42 9 1 2 9 9 1 2 9 1 9 1 13 16 4 9 5 11 1 9 1 13 2 11 1 2 9 1 9 5 9 2 9 9 1 1 9 1 13 4 16 4 2
35 2 9 1 13 16 2 9 9 1 13 9 1 9 1 13 9 4 9 1 9 1 13 16 2 9 1 0 9 9 1 13 9 1 13 2
28 3 9 9 1 13 2 13 4 4 9 1 2 9 1 9 9 2 11 1 9 1 9 1 13 9 1 13 2
30 9 1 13 16 1 9 1 0 9 2 9 1 0 9 7 9 1 0 9 1 2 0 9 1 13 16 14 13 4 2
7 9 1 9 0 13 4 2
7 2 9 1 3 13 4 2
29 11 1 9 1 9 11 11 1 12 12 12 12 9 1 10 9 9 1 11 11 1 9 1 13 16 13 4 4 2
5 11 9 1 9 2
4 9 11 11 2
35 12 12 12 12 9 9 9 9 9 1 9 12 9 1 13 2 12 12 9 1 9 1 2 11 2 1 11 1 13 16 13 4 4 4 2
20 13 16 11 1 2 9 1 9 2 1 9 1 13 2 3 9 1 13 4 2
30 9 9 1 13 9 9 4 9 1 9 1 13 2 9 1 9 1 13 4 16 12 9 1 13 4 9 4 4 4 2
28 11 1 12 12 9 9 1 11 9 1 13 2 10 12 9 9 2 11 2 1 9 9 1 9 1 13 4 2
25 2 9 12 12 12 9 9 9 9 9 9 9 9 2 1 12 9 2 11 5 9 1 13 4 4
25 9 12 9 1 9 1 13 4 4 9 9 1 12 12 9 14 9 12 12 12 12 9 1 9 2
33 11 5 11 1 9 9 1 9 12 2 12 9 12 12 9 7 9 9 9 1 9 1 13 4 2 9 0 4 9 1 13 4 2
19 9 1 2 9 9 2 7 2 0 9 2 14 9 9 1 12 12 9 2
22 0 9 1 9 12 12 12 2 12 12 12 1 9 2 9 9 9 1 13 4 4 2
32 12 9 9 12 9 12 12 12 9 9 2 11 9 11 9 11 9 1 9 11 11 9 9 9 12 9 1 9 9 13 4 2
19 11 1 13 16 2 9 9 9 1 9 9 1 13 2 9 9 1 9 2
21 9 9 1 9 14 1 13 16 4 16 2 9 9 9 1 9 1 0 1 13 2
19 9 1 9 9 1 9 1 13 4 9 1 2 9 1 9 9 1 13 2
9 9 1 9 1 13 4 4 4 2
12 12 9 1 9 9 9 9 1 13 4 14 2
35 11 9 11 9 11 9 1 9 1 9 1 1 3 2 9 1 9 2 9 14 1 9 9 9 9 2 9 9 9 2 1 9 13 4 2
39 9 1 2 11 11 9 9 1 2 9 9 2 1 9 9 1 9 1 13 4 16 4 16 1 9 1 2 9 9 9 2 11 9 9 2 1 9 9 2
21 9 9 1 9 1 9 1 2 9 1 1 9 9 1 9 9 1 9 1 13 2
23 9 9 1 13 9 12 12 9 9 1 9 1 9 1 2 9 1 9 1 13 16 13 2
25 2 9 9 2 1 2 9 1 13 9 1 9 1 9 1 12 12 12 12 9 1 9 9 9 2
34 9 9 1 2 9 1 9 9 7 9 1 1 9 1 9 9 4 9 1 13 2 9 1 9 1 9 1 1 9 1 13 16 4 2
26 7 2 9 1 9 1 12 12 9 1 1 12 12 12 12 9 1 13 16 4 4 16 1 9 9 2
38 2 9 1 9 9 2 1 13 4 9 1 12 12 12 9 1 13 2 9 12 12 12 12 9 1 9 9 9 2 11 9 9 2 9 1 13 4 2
14 9 1 2 9 9 1 9 1 12 2 12 9 9 2
41 9 9 9 9 1 13 9 12 12 9 1 13 4 16 4 16 2 3 1 9 9 4 2 9 2 9 9 2 9 9 2 9 2 9 2 9 14 0 4 9 2
52 11 1 12 9 9 2 9 9 9 1 13 4 4 4 9 1 2 9 13 4 4 4 11 9 1 11 5 9 9 9 1 9 9 1 9 1 9 1 13 16 13 4 16 4 4 9 1 12 9 13 4 2
33 9 1 13 16 2 9 9 9 1 9 9 2 9 1 13 9 1 9 9 1 9 1 9 1 13 16 9 1 13 4 1 13 2
63 12 9 9 12 9 12 9 9 2 11 9 11 9 11 1 9 1 13 16 4 4 9 9 2 9 2 11 9 9 1 2 9 1 13 4 9 9 11 9 11 9 11 2 11 11 9 1 9 9 9 1 13 4 2 9 1 0 13 16 13 4 4 2
25 11 9 9 1 9 1 1 2 9 9 1 9 1 9 1 9 1 9 12 9 14 0 4 4 2
9 11 9 1 9 1 9 4 4 2
30 9 1 1 9 1 9 9 1 9 1 13 16 2 9 1 9 1 9 1 13 16 13 4 16 1 2 9 9 2 2
44 9 9 1 1 9 1 13 4 4 16 4 16 2 9 9 9 1 1 10 9 1 0 2 0 9 1 2 9 2 1 13 4 9 4 2 0 13 4 16 4 2 1 13 2
62 9 9 1 13 4 9 9 9 9 9 9 9 9 9 1 13 4 4 9 9 1 1 9 9 1 13 16 2 9 1 9 1 9 9 1 9 1 0 4 9 14 1 9 1 13 4 4 9 1 9 9 1 13 2 1 13 16 13 4 16 4 2
79 7 2 9 9 9 1 2 12 12 12 12 2 12 12 9 1 2 11 7 9 14 1 9 9 9 1 13 9 9 1 13 16 13 4 4 4 9 1 2 9 9 2 12 12 9 1 13 4 11 9 9 9 9 9 9 1 13 4 9 7 0 4 9 1 9 14 2 9 1 9 1 13 4 9 9 1 13 4 2
22 7 2 10 9 1 9 9 1 13 4 2 9 9 2 1 13 16 1 9 1 0 2
34 7 9 9 9 1 2 3 9 1 9 1 13 16 4 16 1 2 9 7 9 9 1 13 4 4 2 0 4 2 1 13 16 4 2
31 9 9 1 13 16 9 9 9 1 9 9 1 9 1 9 1 13 9 1 1 2 9 9 1 9 9 1 13 1 13 2
43 0 9 9 1 2 9 9 1 13 4 4 16 2 9 9 1 0 16 2 9 9 1 9 1 1 9 9 1 9 1 9 9 1 13 9 1 0 2 1 13 16 4 2
20 12 9 9 12 9 9 2 11 9 11 9 9 12 2 11 9 9 1 13 2
28 9 9 9 1 9 9 1 9 9 1 9 9 12 9 9 9 9 9 9 12 12 12 9 1 13 4 4 2
23 9 1 11 9 1 9 1 13 4 9 2 11 9 1 9 11 9 1 9 1 0 9 2
27 12 9 9 12 9 12 12 9 9 2 11 9 11 9 11 9 11 1 9 2 11 9 2 9 1 13 2
15 9 12 9 9 9 9 12 12 12 9 1 13 4 4 2
26 9 12 9 1 9 9 9 9 1 9 1 2 9 9 1 11 11 9 1 13 4 9 1 13 4 2
27 11 9 1 2 12 9 9 9 1 13 4 4 16 4 1 4 14 1 13 16 2 9 1 13 16 4 2
34 9 1 9 1 1 9 2 11 9 1 9 1 9 1 13 4 9 4 4 9 2 12 9 1 9 9 1 9 9 1 13 4 4 2
11 9 9 1 12 12 12 12 9 1 9 2
16 12 9 1 12 9 2 12 9 1 9 7 9 1 13 4 2
82 12 9 9 2 9 12 9 9 9 9 1 13 4 9 1 13 16 2 9 9 5 9 1 9 9 12 12 9 1 9 1 9 2 9 1 13 4 11 9 1 9 9 2 11 5 9 2 1 9 9 12 9 1 12 9 9 12 9 12 9 9 2 9 9 1 9 11 1 9 9 2 11 2 1 9 9 1 13 4 4 4 2
14 9 1 13 9 2 12 9 1 9 1 13 9 9 2
18 9 11 1 1 12 12 9 1 13 16 4 2 13 12 9 1 9 2
19 9 1 12 9 1 2 9 1 9 9 1 9 9 1 13 4 4 4 2
17 9 1 12 9 9 2 9 1 9 9 9 1 9 1 13 4 2
48 9 1 9 1 13 16 2 9 12 9 12 12 9 9 1 11 9 11 9 12 12 12 9 1 9 12 9 12 12 12 9 9 1 11 9 9 12 12 12 9 1 9 1 9 9 1 13 2
20 10 9 2 9 12 12 9 2 9 1 9 1 9 1 13 16 13 4 4 2
23 2 9 9 1 0 4 13 16 4 4 2 10 9 1 9 1 13 4 1 1 2 9 2
16 11 9 1 9 11 5 11 9 1 12 9 13 4 4 9 2
56 13 4 4 2 9 9 1 9 2 1 12 9 14 13 2 9 1 9 1 12 9 13 4 2 9 1 13 4 11 9 11 9 11 1 11 9 9 1 13 4 11 9 1 2 12 9 1 2 13 4 4 2 1 13 4 2
27 11 9 1 13 4 4 12 9 9 14 1 2 9 1 0 2 9 1 13 16 1 9 4 4 1 13 2
39 2 9 1 9 2 9 11 1 0 4 9 1 3 13 4 2 9 1 9 9 9 14 2 9 14 1 9 0 2 1 13 4 16 4 4 2 1 13 2
39 9 9 1 0 4 2 9 1 9 9 9 9 1 9 9 4 4 11 9 1 2 15 12 12 9 14 2 9 1 1 3 11 11 1 13 16 4 4 2
32 11 9 1 13 16 2 9 1 12 9 1 9 1 14 9 13 2 10 9 1 9 9 1 9 1 9 1 13 16 13 4 2
8 11 9 1 2 9 1 9 2
28 2 13 4 4 9 4 4 2 1 11 9 1 13 4 4 2 10 9 1 9 1 9 1 13 4 1 13 2
14 11 9 9 1 12 9 9 9 1 11 11 1 13 2
15 9 9 1 9 9 1 13 2 9 1 9 1 13 4 2
34 11 9 1 2 12 9 1 13 16 9 1 13 2 9 1 0 16 9 9 1 13 4 1 13 16 4 4 16 4 16 5 5 2 2
40 9 1 13 16 2 11 9 1 9 9 9 9 1 13 4 16 2 12 9 9 12 12 9 9 2 2 12 9 9 1 13 2 1 9 1 9 1 13 4 2
48 9 9 1 2 9 2 1 9 1 13 9 4 9 1 9 1 2 11 9 9 9 1 11 11 9 9 9 7 9 1 11 11 9 9 1 9 1 13 4 9 9 1 3 0 4 13 4 2
34 9 2 9 1 9 1 13 9 9 4 9 1 13 4 4 16 2 9 9 1 9 9 7 9 9 1 9 14 0 13 4 4 4 2
22 11 9 9 9 9 1 2 12 9 9 1 9 1 13 4 9 1 12 12 9 9 2
56 9 9 1 9 12 9 2 9 9 1 9 9 9 1 9 9 1 13 4 2 12 12 12 9 1 9 9 1 9 1 13 2 9 9 14 1 1 9 9 1 9 1 2 9 12 12 9 14 1 9 1 9 1 13 4 2
8 10 9 1 9 1 9 9 2
16 9 9 1 9 1 9 2 9 9 9 1 9 1 13 4 2
24 9 1 9 1 2 9 9 1 9 14 1 9 1 9 1 9 1 13 4 4 16 4 4 2
24 7 2 9 1 9 1 13 16 2 9 7 9 1 9 1 9 9 1 9 1 13 4 4 2
31 9 1 1 9 9 1 2 9 9 12 12 9 2 9 12 12 9 1 9 9 1 9 9 9 1 9 1 13 4 4 2
53 9 1 2 0 9 1 9 1 9 9 1 13 9 1 9 9 1 1 13 9 2 9 1 9 1 9 1 2 9 9 9 1 13 9 1 2 9 1 9 1 9 9 1 13 9 1 9 1 13 4 16 4 2
21 9 1 9 1 9 1 13 0 9 9 1 13 4 9 9 1 9 1 13 4 2
39 9 9 5 11 1 2 9 9 13 9 2 1 12 9 9 2 11 9 11 9 1 11 9 1 13 4 2 9 9 1 9 12 12 12 9 1 13 4 4
27 9 13 9 1 2 12 9 1 9 9 1 13 9 9 1 9 1 2 11 9 1 13 4 1 13 4 2
59 9 12 9 2 0 4 9 9 1 9 12 12 12 9 1 9 9 1 13 4 4 9 2 9 9 1 11 9 1 9 9 9 1 2 9 1 9 1 9 2 9 9 2 9 14 0 4 9 9 1 13 2 3 1 9 1 13 4 2
27 9 1 11 9 9 1 2 13 9 2 1 9 9 1 2 9 9 7 9 2 9 1 13 16 13 4 2
35 9 9 1 2 9 1 13 9 9 2 9 1 13 16 4 4 4 13 16 2 10 9 2 9 9 1 0 1 13 9 1 9 1 13 2
21 10 9 9 1 2 10 9 4 2 9 11 1 9 1 0 9 7 9 1 13 2
19 9 1 0 4 9 1 13 4 4 16 9 1 15 1 0 2 9 2 2
38 3 13 4 9 9 1 9 1 9 1 13 2 9 1 13 16 2 9 9 1 9 1 9 1 13 16 4 4 2 1 9 9 9 1 13 16 4 2
23 9 1 2 9 7 15 1 9 1 9 1 13 12 9 1 9 9 1 9 1 13 16 4
13 3 1 3 9 1 2 9 9 1 9 1 11 2
25 9 1 12 9 1 9 9 1 11 1 9 1 13 4 2 0 2 9 9 2 1 13 16 4 2
17 15 1 9 1 3 13 4 9 1 9 9 9 1 13 16 9 2
37 9 1 12 12 9 9 1 11 5 11 4 2 10 9 9 9 1 13 16 4 16 2 0 4 16 1 2 9 1 9 9 1 13 11 5 9 2
53 2 9 3 2 10 9 1 13 4 4 2 11 9 1 2 9 1 9 1 9 1 9 1 0 2 15 14 9 9 1 13 16 4 9 1 3 0 4 2 9 13 4 2 1 13 16 1 0 4 9 4 4 2
105 2 12 12 9 9 2 9 1 9 1 13 3 9 2 11 9 1 13 9 4 4 14 2 11 9 1 9 1 9 1 13 4 1 2 9 1 13 4 16 4 2 9 1 9 1 2 1 13 4 16 2 9 11 11 2 1 13 4 2 15 1 13 16 2 0 9 2 1 13 9 1 13 16 4 1 13 4 2 15 14 1 13 4 2 9 1 9 9 4 4 11 11 9 1 2 11 1 13 4 9 13 16 4 4 2
48 2 9 1 13 4 4 4 16 2 9 1 13 16 2 12 9 1 13 16 3 13 9 1 13 4 4 2 3 9 4 16 2 1 9 9 1 13 4 16 2 9 4 13 16 13 4 4 2
73 2 13 16 1 0 4 14 2 11 1 13 9 1 2 3 9 13 4 16 1 13 4 2 0 9 1 11 1 9 4 2 3 9 5 1 9 4 16 4 14 2 9 9 1 9 1 13 4 4 16 2 9 1 9 1 13 4 16 1 9 14 4 2 9 1 9 9 9 4 13 4 4 2
73 2 9 1 9 9 1 2 9 1 9 4 4 2 9 1 9 1 9 9 4 1 1 2 9 1 12 9 1 13 4 4 2 9 1 2 9 4 13 16 4 4 4 2 1 13 4 4 4 4 2 9 12 9 2 13 4 4 2 10 9 1 1 2 0 4 9 1 13 4 4 4 14 2
86 2 11 1 9 9 1 9 9 1 2 11 1 9 1 2 11 12 12 9 4 4 2 9 1 0 9 1 13 16 2 0 9 4 4 2 9 1 9 1 13 14 2 9 1 2 9 1 13 9 1 13 4 9 1 13 4 1 2 9 1 13 4 4 2 10 9 1 13 16 1 2 9 1 9 1 13 4 16 2 13 16 1 4 4 4 2
34 11 12 9 2 9 1 9 9 2 9 1 0 1 9 9 1 13 16 13 4 2 11 1 9 1 9 1 13 16 1 12 12 9 2
65 15 1 13 4 16 11 1 9 9 4 9 7 2 9 9 1 9 2 11 11 9 9 9 1 9 9 1 9 1 13 4 2 2 11 2 7 2 11 2 5 11 1 9 9 2 1 12 9 1 12 12 9 14 11 9 11 9 1 11 9 9 1 13 4 2
26 9 1 2 11 1 11 9 9 9 9 1 9 1 12 9 14 0 1 13 11 1 9 14 1 13 2
43 11 1 9 2 11 11 2 11 11 2 11 11 9 1 9 1 13 9 12 12 12 9 1 13 4 2 11 9 1 9 9 2 9 11 11 1 9 1 13 4 16 4 2
13 9 2 11 1 9 1 9 1 9 4 4 9 2
44 10 9 9 1 9 1 0 4 9 1 13 2 9 1 3 13 4 2 3 12 9 1 9 1 12 12 12 12 1 1 9 1 13 16 2 3 9 1 13 4 11 1 9 2
31 11 9 1 13 16 10 11 1 9 9 1 9 13 4 2 3 11 1 9 1 4 4 11 1 9 1 9 1 13 4 2
24 12 9 5 12 12 9 12 12 9 5 12 12 9 2 9 1 12 12 9 14 2 11 9 9
13 9 9 1 9 7 12 12 9 9 1 9 9 2
14 12 9 12 12 9 2 9 9 12 12 9 9 9 2
11 2 11 7 11 1 9 2 11 11 9 2
82 12 9 9 12 9 12 12 9 9 2 11 9 11 9 11 9 1 11 9 9 9 5 9 9 2 11 11 9 5 4 2 9 9 1 13 16 4 4 9 9 2 9 2 11 11 9 9 1 2 9 9 1 13 4 11 9 1 9 1 13 2 2 12 12 9 14 13 16 4 2 12 9 9 1 1 13 2 1 9 1 13 2
24 11 9 1 13 4 2 9 1 13 4 16 2 11 9 9 1 15 1 13 4 1 13 4 2
28 9 1 13 4 9 11 9 1 9 9 12 12 9 1 11 9 9 9 9 1 9 1 11 9 9 1 13 2
26 9 9 13 4 9 2 2 9 1 13 4 2 1 13 4 9 2 9 9 9 1 9 9 13 4 2
22 9 2 9 1 9 1 13 4 2 11 9 7 9 9 12 9 1 9 1 0 4 2
52 9 13 9 1 9 1 13 9 12 9 13 4 4 4 11 9 9 1 2 9 1 9 9 1 13 11 5 9 1 9 9 7 9 9 1 9 9 1 3 13 2 9 1 13 16 13 0 9 1 13 4 2
15 9 9 4 9 9 9 1 9 1 13 9 1 9 9 2
22 9 9 1 9 1 9 9 1 9 1 13 4 9 2 9 1 9 9 9 1 13 2
13 15 14 9 1 9 9 1 13 4 16 4 4 2
51 9 2 9 9 1 0 9 9 7 9 9 1 9 9 9 1 9 1 9 1 13 16 2 9 9 9 1 9 9 1 13 2 9 1 9 9 9 1 2 1 1 9 1 9 1 11 9 1 13 4 2
32 10 9 2 11 9 1 13 4 4 11 9 9 9 1 1 2 9 1 9 2 1 13 16 9 9 1 9 9 9 1 13 2
26 11 9 1 9 1 11 9 1 13 9 7 9 9 1 9 1 2 9 1 1 9 1 9 9 4 2
51 11 11 9 1 9 1 9 1 11 9 9 1 13 4 16 2 9 11 1 9 9 1 11 1 9 1 13 16 4 16 1 13 16 2 9 1 1 12 9 1 13 4 4 2 1 9 9 1 13 4 2
27 11 9 1 1 11 11 5 9 9 1 9 9 1 13 4 16 4 16 2 9 1 1 0 4 9 1 2
75 9 9 1 13 9 9 2 9 1 9 1 13 9 2 9 9 1 11 11 9 1 2 0 4 13 0 9 2 10 9 1 2 9 9 1 9 9 4 13 4 4 9 1 1 4 2 9 9 1 13 4 9 2 9 9 4 9 1 0 2 9 9 1 9 1 9 1 13 16 4 4 2 1 13 2
51 9 9 9 1 12 9 2 9 1 13 4 4 9 12 12 9 1 9 1 9 1 13 16 13 9 9 1 2 9 9 2 1 13 2 9 9 9 1 9 7 9 1 13 9 1 2 9 1 13 4 2
16 9 1 13 4 4 11 9 1 9 9 1 13 16 4 9 2
48 9 9 1 9 9 1 13 4 9 9 12 9 2 0 9 9 12 12 9 1 9 9 1 9 12 12 12 12 9 1 9 9 1 9 1 13 2 9 1 13 9 12 12 9 1 13 4 2
16 12 9 14 9 9 12 12 9 1 9 12 9 1 13 4 2
24 9 1 9 9 1 9 9 1 12 9 2 9 12 9 1 12 12 12 12 9 1 13 4 2
10 9 9 1 9 1 12 9 1 0 2
27 12 12 12 12 9 9 1 9 9 1 11 9 11 9 11 2 9 9 9 9 12 9 2 11 11 9 2
22 9 1 11 9 11 9 1 9 1 9 13 2 9 12 9 1 9 9 1 13 4 2
22 9 9 1 2 9 9 1 11 11 9 1 9 9 1 13 2 9 1 13 4 4 2
14 9 9 1 9 9 9 1 12 2 12 9 1 13 2
47 9 9 1 9 12 12 12 9 1 2 11 9 1 12 12 9 1 13 16 2 9 9 1 9 9 9 1 9 13 2 9 9 1 12 9 9 2 12 12 12 12 9 1 13 16 4 2
18 9 2 9 1 9 9 1 9 1 13 4 4 9 1 0 4 4 2
33 9 1 0 9 7 9 1 9 9 1 9 1 1 2 9 1 13 16 2 9 1 9 7 9 14 1 13 9 1 13 16 4 2
5 9 1 0 4 2
28 15 1 15 1 0 4 16 2 9 3 1 9 1 13 4 4 2 13 9 1 13 4 16 1 13 9 4 2
25 9 9 9 1 11 11 9 1 9 2 11 1 9 2 1 9 1 13 4 16 4 9 1 13 2
30 13 4 9 4 4 11 11 9 1 2 0 9 2 9 1 9 1 13 16 4 16 2 9 14 9 1 13 4 4 2
25 3 4 4 1 13 16 13 16 2 2 15 1 2 13 4 16 4 14 2 1 13 4 1 13 2
19 9 7 9 1 13 4 9 2 9 1 9 1 14 13 4 9 1 13 2
5 15 1 0 4 2
31 9 9 1 9 11 9 1 9 1 0 4 4 16 2 3 13 4 9 1 13 4 9 1 9 9 1 13 16 4 4 2
32 9 1 9 11 11 1 13 16 11 9 1 2 0 9 1 9 9 1 9 1 9 9 1 0 2 1 13 4 16 4 4 2
22 9 1 9 9 1 2 9 1 13 4 9 1 3 13 4 16 4 4 16 4 4 2
32 9 14 0 4 9 4 9 1 9 1 13 4 2 9 4 13 4 9 1 9 1 13 4 2 14 13 9 1 0 4 4 2
3 11 11 9
24 9 9 9 1 9 1 13 4 9 1 2 9 1 0 1 11 9 1 13 4 4 16 4 2
43 11 9 1 13 4 4 4 9 12 9 9 2 12 9 5 12 12 9 2 9 1 12 9 2 0 9 1 9 9 12 9 1 0 4 13 2 9 12 9 1 13 4 2
49 11 9 1 9 1 1 2 9 11 9 1 9 9 9 1 9 9 12 12 12 9 2 9 11 9 1 13 4 4 9 1 12 9 4 2 9 9 1 2 11 12 12 12 12 12 12 9 2 2
19 9 9 1 11 9 1 9 9 9 1 13 4 4 9 1 9 4 4 2
18 9 9 1 9 4 2 9 9 1 2 9 9 2 1 13 16 4 2
9 11 9 9 1 13 9 1 13 2
28 9 9 1 13 9 9 4 13 2 9 9 1 0 4 13 4 4 9 9 9 1 13 4 16 4 9 4 2
37 11 9 9 1 9 1 9 12 9 1 0 4 2 11 14 1 9 1 9 1 13 16 1 12 12 9 1 2 9 12 12 9 1 13 16 4 2
30 9 9 1 9 9 1 9 1 9 9 1 13 1 13 16 0 9 4 16 2 9 1 3 9 9 1 13 4 4 2
21 11 9 14 1 13 16 2 11 9 1 9 9 1 9 12 12 12 12 12 9 2
15 9 12 12 12 12 9 4 4 11 9 1 9 1 9 2
10 10 9 9 1 11 9 14 3 13 2
65 9 9 1 0 4 13 9 9 9 1 13 4 4 16 1 9 9 1 4 2 9 9 9 1 2 11 5 9 2 1 1 2 9 12 9 5 9 12 12 12 9 9 1 11 9 9 9 1 11 9 1 9 1 12 12 12 12 9 0 12 12 9 1 13 2
43 2 9 5 9 2 1 9 12 9 5 12 12 12 9 9 1 9 1 13 16 1 2 11 0 9 9 1 1 9 1 12 12 12 12 9 0 12 12 12 12 9 1 2
25 2 9 2 1 2 11 9 1 12 12 12 12 9 0 12 12 12 12 9 1 13 4 16 4 2
54 9 9 1 9 9 1 9 1 9 9 1 9 1 13 2 9 1 9 9 1 9 1 9 9 1 13 16 9 9 1 9 9 9 1 13 16 4 2 10 9 1 9 9 1 9 1 13 4 9 1 13 16 4 2
11 10 9 1 1 9 9 1 9 1 13 2
38 11 9 1 9 2 11 9 7 11 14 12 9 1 13 16 4 16 2 11 9 1 11 9 9 1 9 12 9 1 2 9 12 12 9 1 13 4 2
15 9 1 9 9 9 1 9 12 9 13 4 4 1 13 2
40 9 1 2 13 4 4 16 2 15 1 13 14 9 1 13 4 2 9 9 9 1 9 9 1 13 4 2 9 1 13 0 9 1 9 2 1 13 16 4 2
47 0 9 9 1 13 16 11 5 9 1 2 9 9 1 13 9 9 1 13 2 9 9 1 9 9 2 0 9 1 3 13 4 4 16 2 3 10 9 1 13 16 4 1 2 1 13 2
40 15 1 13 9 9 9 9 1 2 9 1 9 9 14 13 4 16 2 9 9 1 9 9 9 2 9 9 4 13 16 9 1 13 4 2 1 13 16 4 2
30 9 9 1 9 9 4 13 9 1 9 1 13 4 9 9 9 9 1 9 9 13 4 2 9 1 13 4 4 4 2
25 13 4 16 4 4 9 9 1 9 1 3 13 4 9 1 13 4 9 4 2 10 9 1 0 2
47 11 9 1 2 9 9 9 9 1 13 9 1 9 9 1 9 1 13 2 9 1 9 9 9 4 9 9 9 14 1 1 0 4 9 1 13 4 4 4 9 1 15 9 1 13 4 2
39 9 7 9 1 9 9 1 9 7 9 9 9 1 1 9 1 9 1 13 4 9 4 4 2 9 9 1 13 16 0 4 9 1 1 4 4 4 14 2
48 9 9 9 9 1 9 2 9 1 9 1 13 4 16 1 2 9 1 9 9 1 13 4 9 1 9 9 9 4 4 2 9 9 9 2 1 2 0 9 1 9 1 13 4 14 4 4 2
35 9 9 2 9 9 9 14 9 12 9 7 9 9 9 9 1 2 9 9 9 1 0 9 1 13 4 4 2 1 13 16 13 4 4 2
41 7 2 9 1 9 9 1 13 4 2 9 9 1 13 9 9 2 1 1 2 9 9 9 1 9 1 9 1 13 4 1 1 9 1 0 9 1 13 4 4 2
17 9 9 9 1 3 13 14 1 2 10 9 1 9 9 4 4 2
21 15 9 1 2 9 1 9 14 9 1 13 16 4 1 9 1 13 16 4 4 2
19 9 9 4 1 2 9 9 9 1 9 1 3 13 4 9 1 13 4 2
39 9 9 4 1 3 2 9 9 1 9 9 9 1 13 9 1 9 9 4 9 1 9 1 13 4 2 9 9 1 13 4 16 9 1 13 4 4 4 2
40 7 2 0 9 7 9 1 9 1 9 1 13 4 9 2 9 9 1 9 9 7 9 1 9 9 1 13 4 7 2 9 1 13 9 1 0 4 13 4 2
19 15 1 9 4 9 4 4 2 9 1 9 1 13 4 9 1 13 4 2
30 11 11 9 1 2 9 9 1 2 9 9 2 9 9 2 9 9 1 13 9 1 9 0 9 1 13 16 4 4 2
38 9 9 1 1 2 9 9 9 9 1 9 9 1 13 16 4 4 16 2 9 9 14 9 9 1 9 1 13 4 7 4 16 9 1 13 4 4 2
17 9 9 1 9 7 9 1 13 4 1 13 4 4 16 4 4 2
17 1 1 13 2 15 1 3 9 9 1 13 1 1 13 4 4 2
7 13 4 4 9 1 0 2
16 10 9 1 2 9 9 9 1 9 12 9 1 9 4 4 2
19 0 9 9 1 13 4 14 1 2 9 1 9 1 13 4 4 16 4 2
40 9 9 1 1 9 9 1 2 13 1 13 9 1 0 16 2 9 1 1 9 1 9 9 4 9 1 13 9 9 7 9 9 9 1 0 13 4 4 4 2
10 9 9 9 1 13 14 13 16 4 2
19 3 9 1 2 9 1 3 9 9 13 16 4 14 1 0 4 9 4 2
31 9 9 9 14 1 9 1 2 3 13 4 16 4 16 14 13 16 2 9 1 9 9 9 7 9 1 9 1 13 4 2
19 10 9 1 1 9 1 13 4 4 16 2 3 9 1 9 1 14 4 2
25 9 9 1 13 16 9 7 9 9 1 2 3 0 9 1 9 7 9 9 1 13 4 16 4 2
21 9 9 1 13 16 2 0 4 9 9 9 1 13 16 4 9 1 13 4 4 2
9 9 1 1 13 4 9 1 13 2
46 9 9 1 1 2 9 1 9 1 13 16 4 1 13 16 4 1 4 2 2 9 9 2 1 13 16 4 1 13 14 1 9 1 13 2 9 1 1 9 1 3 13 4 4 4 2
48 9 9 1 12 12 12 9 13 4 4 2 9 9 9 2 1 2 11 1 0 4 9 9 1 13 16 4 1 13 4 2 12 12 9 9 1 9 9 1 11 9 9 1 0 4 13 4 2
35 9 1 2 11 9 1 0 11 9 1 13 1 1 2 11 9 9 1 9 1 13 9 9 7 11 9 1 0 4 13 4 9 4 4 2
54 11 1 9 9 2 9 9 9 7 11 9 9 9 1 9 1 13 9 9 1 9 1 13 4 9 9 1 9 1 13 2 11 1 1 9 9 1 9 9 1 3 0 4 16 14 1 2 9 1 13 13 16 4 2
44 7 2 9 1 1 11 9 1 13 4 16 14 2 11 1 3 9 1 9 1 13 4 2 9 9 1 9 7 11 9 9 9 1 13 4 16 4 14 1 13 4 16 4 2
23 9 9 1 9 1 13 4 2 9 9 1 9 9 1 13 4 9 1 1 13 16 4 2
29 9 1 2 11 1 9 7 9 9 1 9 9 1 2 11 1 1 9 4 9 1 13 4 4 9 1 13 4 2
22 7 2 11 9 9 1 4 4 9 9 1 2 13 4 0 9 1 13 4 16 4 2
49 0 9 9 1 2 11 1 11 1 1 9 9 9 1 13 4 16 2 2 9 1 9 1 2 11 7 9 9 1 9 9 4 9 1 13 4 9 1 13 16 13 0 9 1 13 2 1 9 2
18 7 2 9 1 13 2 9 9 9 2 1 1 9 1 13 16 4 2
28 11 9 1 2 9 9 9 1 13 11 1 9 9 1 2 9 1 9 1 9 9 9 1 13 16 4 4 2
54 15 1 13 9 1 2 11 1 9 9 1 13 16 1 2 9 9 1 11 1 9 1 13 1 13 4 4 9 1 2 11 1 9 9 1 2 9 9 7 9 1 9 0 1 1 13 4 4 1 13 4 16 4 2
35 9 9 1 13 4 16 1 2 11 1 9 9 1 0 4 13 1 1 9 1 0 4 13 4 9 4 2 3 9 9 4 9 1 13 2
59 11 1 1 9 1 13 16 1 2 2 11 14 0 4 12 9 9 9 1 0 2 1 13 2 9 9 9 1 2 11 1 9 9 9 1 9 1 13 2 1 0 13 4 2 11 1 9 1 0 11 9 9 1 9 1 13 16 4 2
27 9 1 7 2 9 9 9 1 9 9 14 1 13 4 9 9 7 2 9 1 13 9 1 9 1 13 2
27 9 11 1 9 9 7 9 9 9 1 9 1 2 9 11 9 9 9 9 1 9 1 13 4 16 4 2
37 9 1 9 1 2 11 1 9 1 2 9 2 13 4 2 15 14 1 0 0 4 9 9 7 11 9 1 13 4 9 1 13 16 13 4 4 2
28 7 2 11 1 9 1 9 1 3 13 4 4 16 4 9 1 1 2 9 1 13 4 9 1 1 13 4 2
35 11 1 9 9 1 9 1 13 9 1 13 16 1 4 16 2 11 1 9 1 9 1 13 16 3 0 4 9 9 4 9 1 0 4 2
36 9 9 9 1 9 9 9 7 2 11 7 11 1 9 1 13 4 16 4 9 1 2 9 9 1 9 1 9 9 1 13 4 9 4 4 2
34 9 1 9 1 1 2 11 1 9 1 13 4 4 16 4 16 2 9 1 9 9 7 9 1 3 13 1 1 13 4 4 4 4 2
38 9 9 9 1 9 9 1 1 9 9 1 13 4 14 3 14 1 13 4 4 9 1 2 9 1 10 0 9 1 9 1 13 9 9 1 13 4 2
18 9 9 9 1 9 9 1 9 1 0 13 4 4 9 1 13 4 2
32 9 11 9 12 9 9 1 9 9 1 13 4 4 16 2 3 9 9 4 9 1 13 16 1 0 13 4 9 1 13 4 2
61 7 2 2 9 1 9 9 9 1 9 9 1 13 4 9 1 13 9 1 9 9 2 13 4 4 16 4 4 2 1 13 9 2 2 10 4 4 9 1 13 4 16 1 13 16 9 1 9 1 13 9 4 1 4 2 1 1 13 16 4 2
15 9 1 9 9 1 3 9 1 13 4 4 9 4 4 2
16 9 1 0 4 13 2 9 1 13 4 4 4 16 4 4 2
31 9 9 1 13 16 1 9 9 2 9 9 1 9 2 4 4 2 9 1 9 9 9 1 9 9 1 13 16 4 4 2
77 9 9 9 1 13 16 1 2 9 1 13 4 2 1 9 1 13 4 16 4 2 2 9 2 1 9 1 13 9 1 1 4 4 16 2 9 1 2 9 1 9 9 1 0 4 13 4 9 9 1 10 9 1 9 1 9 1 13 13 4 4 2 1 13 9 1 9 9 1 9 1 13 9 1 13 4 2
13 9 9 1 9 1 13 4 9 1 13 16 4 2
29 9 1 9 2 9 9 1 9 9 1 13 4 9 1 1 3 0 9 1 13 2 1 13 9 1 13 16 4 2
8 0 4 9 1 9 1 13 2
53 9 2 2 9 1 9 1 9 9 1 13 4 16 4 2 9 9 1 9 1 13 4 9 1 13 4 16 1 2 9 9 1 9 1 13 4 4 2 1 2 9 9 9 1 13 4 9 1 13 16 4 4 2
81 9 9 1 1 2 9 1 13 4 16 2 9 1 9 9 1 9 9 1 9 9 1 9 1 13 4 16 4 1 1 11 1 13 2 2 7 2 9 9 1 0 4 9 9 4 4 9 9 9 1 9 1 9 1 13 4 4 9 1 0 1 13 11 1 13 2 1 9 1 9 1 9 1 13 9 1 13 16 4 4 2
22 0 9 1 9 1 9 9 1 13 4 4 9 4 2 9 1 9 1 1 13 4 2
19 9 9 9 1 9 9 9 1 13 9 1 15 12 9 13 16 4 4 2
45 2 9 1 13 9 1 13 4 16 0 4 9 1 1 13 4 4 2 1 13 9 1 9 1 13 9 1 9 9 1 9 14 4 4 2 9 1 9 9 1 1 13 16 4 2
50 12 12 12 12 9 9 1 11 9 1 11 9 1 9 9 1 1 9 9 1 9 1 13 9 9 1 13 4 4 16 1 9 1 2 9 1 9 9 1 9 9 7 9 1 9 1 13 16 4 2
14 9 1 1 9 9 9 1 9 9 1 13 16 4 2
42 7 2 9 1 9 9 9 1 9 1 9 9 9 1 13 4 2 9 9 9 1 9 1 1 9 9 1 13 9 1 1 9 9 9 1 13 4 4 16 4 4 2
29 2 9 1 9 1 9 9 1 13 9 1 9 9 1 13 2 1 9 9 4 1 13 4 9 1 9 1 13 2
24 2 3 9 1 13 9 9 1 13 16 1 9 9 1 13 4 4 2 1 13 9 1 13 2
49 9 1 9 9 9 1 9 1 9 1 2 9 1 9 9 9 1 9 9 7 9 9 1 12 12 9 1 1 9 9 9 2 9 9 9 1 9 9 9 9 1 13 4 1 13 4 16 4 2
12 9 1 9 1 9 1 9 9 1 13 4 2
15 0 9 1 13 4 9 9 1 13 9 1 13 16 4 2
29 9 9 1 9 1 13 4 16 4 4 9 1 9 9 11 9 1 2 3 3 1 0 4 13 4 4 16 14 2
27 3 12 12 12 9 1 9 1 2 9 1 12 12 9 9 1 9 1 13 4 9 1 13 4 16 14 2
8 3 13 4 4 9 4 4 2
21 9 9 1 3 3 13 16 4 4 9 2 3 1 9 1 13 9 1 13 4 2
16 7 2 10 9 1 9 1 2 11 1 9 1 1 13 4 2
29 9 1 9 1 3 13 2 9 9 1 9 1 13 16 11 1 9 2 9 2 9 9 1 9 1 13 16 4 2
21 3 2 9 1 9 1 13 16 1 2 9 1 9 1 13 4 9 9 4 4 2
38 9 9 1 9 2 9 1 13 4 9 2 9 14 1 9 9 9 1 13 4 9 1 13 4 9 1 13 16 2 9 9 1 9 4 13 16 4 2
38 9 1 9 2 9 14 1 9 9 1 13 2 9 9 1 13 9 1 9 1 13 9 2 0 9 1 0 9 1 13 2 9 9 4 9 1 13 2
31 7 2 9 1 9 9 9 1 9 13 4 4 4 9 9 9 1 9 1 9 2 9 9 1 9 1 9 1 0 4 2
29 7 2 11 1 1 10 9 1 13 2 9 1 9 9 2 9 9 9 1 1 0 4 9 9 1 13 16 4 2
27 9 9 2 9 1 9 9 1 9 1 9 2 9 9 1 9 1 9 9 14 2 9 9 1 0 4 2
21 11 9 1 9 1 2 3 9 9 1 9 4 9 1 9 1 13 4 9 4 2
12 9 1 3 9 9 1 13 4 4 16 14 2
12 9 1 9 9 14 1 2 10 9 1 0 2
21 11 1 1 11 9 1 10 9 4 12 12 12 12 12 9 1 9 1 13 4 2
33 9 11 9 9 9 1 1 2 9 9 1 9 1 9 1 9 1 13 4 2 9 5 9 14 0 9 1 9 1 13 16 4 2
33 11 1 9 1 9 1 9 1 13 2 9 1 9 9 1 13 16 4 2 10 9 9 9 1 13 4 4 9 1 13 16 4 2
22 7 9 1 3 1 0 4 9 1 13 16 1 2 9 9 1 13 16 4 16 4 2
17 7 2 9 1 9 9 1 13 16 4 2 9 1 13 4 4 2
30 9 9 1 0 4 9 9 9 1 1 2 9 9 1 9 2 9 9 1 9 1 13 16 4 1 13 9 1 13 2
21 7 2 9 9 1 13 9 9 1 0 9 1 2 13 16 13 4 16 4 4 2
25 12 9 1 9 1 13 16 1 2 9 1 4 4 2 9 5 9 9 1 9 1 13 16 4 2
29 9 9 9 1 9 1 1 2 15 14 1 9 9 1 9 2 9 1 9 1 13 9 1 13 4 16 4 4 2
22 9 1 9 1 9 1 13 14 1 2 9 9 7 9 1 9 1 13 11 1 0 2
29 7 2 9 5 9 9 1 9 1 13 4 9 1 1 2 9 9 7 9 9 1 9 1 0 9 13 4 4 2
33 9 9 1 9 9 1 13 4 4 16 2 9 9 1 13 2 9 1 9 9 1 1 9 1 13 9 1 13 4 4 16 4 2
13 9 9 1 15 9 1 9 1 1 4 9 4 2
24 10 9 1 2 13 4 9 9 1 1 2 3 9 1 13 9 1 13 4 4 16 4 4 2
15 15 1 9 1 15 14 1 9 1 13 4 1 13 4 2
19 9 1 9 1 13 2 2 15 1 12 9 1 9 1 13 16 4 2 2
16 0 4 16 1 9 1 1 4 2 9 4 16 4 5 5 2
26 9 1 12 9 1 9 1 13 16 2 9 9 9 1 9 1 9 1 9 1 13 9 4 1 13 2
13 13 16 12 9 9 1 13 4 4 1 1 13 2
21 3 13 16 2 0 4 9 9 1 0 4 13 9 1 0 2 4 16 1 13 2
28 15 1 0 4 9 4 16 14 0 4 16 2 3 9 1 9 7 9 1 9 1 9 1 13 4 4 4 2
29 9 1 13 16 1 3 0 4 9 14 2 9 1 13 16 4 16 14 2 3 0 4 9 1 13 9 4 4 2
15 3 9 12 1 2 10 9 1 13 4 9 9 4 4 2
35 2 9 9 9 1 9 9 9 9 2 1 9 9 9 1 0 9 9 4 4 4 2 12 12 9 1 9 1 9 9 1 13 4 4 2
28 9 1 9 9 9 1 13 4 4 1 13 16 2 9 1 9 1 9 9 2 10 9 2 9 9 4 4 2
10 7 13 4 9 1 3 1 12 9 2
21 9 9 1 1 9 4 2 9 1 9 1 9 1 13 4 16 1 9 1 0 2
10 9 12 1 9 1 0 4 9 4 2
12 7 9 9 9 1 9 1 0 4 1 13 2
13 9 1 13 16 9 9 1 13 16 4 4 4 2
16 9 1 9 0 9 9 1 9 9 1 13 16 13 16 4 2
18 9 1 3 9 1 9 9 1 9 9 9 9 9 1 9 9 4 2
17 9 9 1 13 9 1 9 9 1 13 9 1 0 9 1 13 2
29 9 1 9 9 14 2 9 9 14 1 13 4 16 2 9 1 13 4 9 1 9 1 0 4 13 4 16 4 2
31 9 12 1 2 7 15 1 3 0 4 9 4 16 2 9 9 7 2 10 0 1 9 1 13 9 9 1 9 4 4 2
35 9 9 1 9 1 2 9 1 9 1 9 13 4 4 9 2 1 9 1 13 16 4 16 2 3 13 4 14 1 13 4 16 4 4 2
29 11 9 11 9 1 9 1 9 9 9 1 9 1 9 9 1 13 4 16 4 4 9 1 9 2 13 4 4 2
18 9 1 9 1 0 9 1 0 16 2 3 9 1 13 16 4 4 2
8 3 9 9 1 13 4 4 2
15 9 1 13 16 1 2 10 9 1 9 9 4 16 4 2
12 9 1 15 1 2 13 4 9 4 1 4 2
14 7 9 1 9 1 9 1 13 4 4 1 13 4 2
19 9 9 9 1 9 1 13 9 9 1 13 16 3 12 12 9 9 13 2
22 9 9 9 1 9 1 3 9 1 9 9 9 1 9 9 1 13 4 16 4 4 2
21 11 9 1 0 4 13 4 16 4 16 2 9 1 3 13 16 13 16 4 4 2
11 9 1 0 13 4 16 4 16 4 4 2
10 9 9 1 1 9 1 9 1 13 2
35 9 1 9 1 13 9 1 0 4 13 9 2 3 1 9 1 9 1 9 1 3 13 4 4 16 4 14 1 13 4 9 2 4 4 2
25 9 9 9 1 13 16 2 9 1 9 1 13 9 1 9 1 13 4 9 1 13 9 4 4 2
14 7 10 9 1 9 2 3 9 9 13 4 16 4 2
23 9 9 9 1 9 1 1 13 4 16 2 9 1 9 1 9 1 13 4 4 1 13 2
15 10 9 13 4 9 1 9 9 1 13 4 4 4 14 2
39 2 9 1 0 4 4 2 9 1 13 4 4 2 9 1 9 4 4 2 1 13 16 1 11 5 11 1 13 4 9 9 1 9 1 1 9 4 4 2
17 9 1 9 9 1 13 16 4 4 4 4 2 10 9 1 13 2
15 2 9 4 16 14 13 4 9 2 9 3 13 16 2 2
30 9 9 1 9 9 1 2 3 1 0 9 1 13 4 9 9 9 1 2 9 9 1 9 9 1 13 4 9 4 2
17 9 1 13 9 9 9 1 9 1 2 0 4 13 4 16 4 2
13 9 1 9 1 9 1 9 0 9 1 13 4 2
12 9 1 3 0 13 4 4 4 16 4 4 2
17 7 9 9 1 9 9 13 9 2 9 1 9 1 13 9 4 2
25 9 1 9 9 1 13 4 9 1 9 1 2 9 9 1 1 13 9 7 9 1 3 13 4 2
22 11 9 1 1 9 9 2 9 12 9 12 12 9 1 9 9 1 13 16 4 4 2
19 9 11 5 11 9 14 9 9 9 1 2 9 7 9 1 9 1 0 2
21 7 9 9 1 13 4 9 9 9 1 9 12 12 9 13 4 1 13 4 4 2
25 9 1 13 4 2 9 7 9 1 13 4 16 2 9 1 3 0 4 13 4 4 16 4 4 2
11 9 1 0 2 9 9 1 9 1 13 2
6 9 1 13 4 4 2
21 9 7 9 9 1 13 2 9 1 13 4 4 9 9 1 9 1 13 16 4 2
14 9 1 9 1 9 4 9 9 1 9 1 1 4 2
13 9 13 4 9 1 9 1 13 16 1 9 0 2
37 9 9 1 2 13 4 4 9 9 1 13 9 1 9 7 9 13 1 13 16 4 16 2 9 5 9 1 9 9 4 9 1 1 13 4 4 2
35 9 9 1 9 2 9 1 9 2 9 9 1 9 2 9 9 1 9 1 13 9 9 14 2 15 1 9 1 13 4 9 1 13 4 2
34 7 2 9 9 1 9 9 4 4 9 9 1 1 2 9 14 1 9 1 1 9 7 9 1 13 4 2 1 1 9 1 13 4 2
6 9 1 9 1 13 2
11 9 0 4 9 9 1 13 4 4 4 2
30 9 9 1 1 9 9 14 1 2 9 1 9 9 1 12 9 1 13 4 4 1 13 4 0 4 13 4 16 4 2
15 9 9 9 9 1 2 3 0 9 1 13 4 16 4 2
15 9 1 9 9 1 13 4 4 16 4 1 13 16 4 2
27 11 14 1 9 1 13 9 1 9 1 9 4 16 2 9 9 1 9 1 13 4 16 13 9 1 0 2
11 9 9 1 0 4 16 1 10 9 4 2
24 10 9 2 9 1 9 1 9 1 13 16 4 9 9 1 9 1 13 16 1 9 4 4 2
11 9 1 9 1 13 4 9 1 13 4 2
16 9 9 1 0 9 9 9 1 9 1 0 4 13 16 4 2
21 12 9 9 1 9 9 1 9 9 1 13 4 4 2 9 9 9 1 9 4 2
23 3 2 9 9 1 13 4 2 1 1 9 1 9 9 1 9 9 1 13 4 16 4 2
26 9 7 9 1 13 16 1 2 9 9 9 1 13 9 1 9 9 9 1 13 4 4 13 16 4 2
10 9 9 9 1 13 4 9 1 13 2
27 0 9 9 1 9 7 9 9 1 9 1 13 4 4 2 9 1 13 4 4 9 1 13 4 4 4 2
26 9 9 9 1 9 9 1 9 1 9 1 0 9 4 16 2 9 1 1 0 13 4 9 1 13 2
30 9 9 9 1 9 9 2 9 9 1 0 4 9 9 2 9 9 1 9 14 2 0 4 9 1 0 4 13 4 2
29 9 9 9 1 3 2 9 9 9 9 1 9 9 1 2 9 1 9 1 13 16 3 9 1 13 9 4 4 2
16 9 1 9 1 1 2 9 1 13 4 13 1 13 16 4 2
23 9 1 9 0 9 1 9 1 2 9 9 1 13 4 4 4 9 1 9 1 13 4 2
33 11 9 1 9 9 1 13 9 7 9 2 9 9 7 9 1 9 1 13 16 2 15 1 0 9 1 13 16 4 1 1 13 2
43 10 9 2 9 9 7 9 9 1 9 9 14 1 13 16 12 12 9 1 13 4 16 4 4 2 11 5 11 9 9 2 1 2 9 1 2 7 0 9 1 13 4 2
22 11 9 5 9 1 13 9 9 7 9 9 1 9 9 1 2 7 0 4 13 4 2
21 9 1 9 1 1 2 9 1 9 1 0 9 1 13 4 1 13 4 16 4 2
35 9 9 1 13 11 9 11 9 1 2 9 1 3 0 9 1 13 2 9 7 9 14 9 9 1 13 4 9 1 3 2 0 4 4 2
26 2 10 9 1 13 16 4 9 1 1 4 2 1 1 9 1 2 9 3 0 13 4 16 4 4 2
32 9 9 1 9 9 1 3 13 2 9 9 9 1 9 1 13 9 1 0 4 13 4 16 1 13 4 4 9 1 13 4 2
38 9 9 1 2 9 9 1 9 12 9 1 13 12 12 12 9 1 2 9 9 2 4 4 2 9 9 1 9 7 9 9 1 9 1 13 1 13 2
11 0 9 14 13 4 9 4 9 4 4 2
9 9 1 9 1 3 13 4 4 2
12 7 2 0 4 9 1 13 4 1 13 4 2
21 9 9 1 13 4 4 9 9 1 12 9 9 1 13 2 1 13 4 14 4 2
14 10 9 9 1 1 13 13 4 9 1 13 4 4 2
43 7 2 9 1 1 2 9 9 9 1 9 9 9 1 13 4 2 9 1 1 9 9 7 9 9 7 1 9 9 1 13 14 2 9 9 1 9 1 0 4 13 4 2
17 9 9 1 2 9 1 9 2 1 13 9 1 0 14 1 13 2
35 9 9 9 1 2 9 1 0 4 9 1 13 4 4 9 1 1 2 9 9 1 13 9 1 9 9 1 1 9 9 1 9 1 13 2
34 11 11 2 11 12 9 2 11 2 9 1 12 9 9 1 2 15 1 9 1 9 9 9 1 13 2 9 1 13 16 4 16 4 2
37 9 1 9 1 9 1 9 9 1 2 3 2 9 9 1 9 1 13 9 1 1 9 1 13 9 4 2 0 9 1 13 16 4 9 4 4 2
18 7 1 2 0 9 1 13 4 4 4 9 1 2 3 0 4 4 2
42 9 9 1 1 9 9 1 13 16 2 9 9 9 1 9 1 13 4 16 4 9 9 9 9 1 9 7 11 9 9 1 2 9 1 13 16 4 4 9 4 4 2
28 11 1 9 1 3 2 9 9 1 13 4 9 9 9 1 2 9 9 9 1 13 9 1 0 4 0 4 2
11 9 1 10 9 1 9 1 9 4 4 2
20 9 9 1 1 9 9 1 2 11 11 7 11 9 9 1 1 13 16 4 2
50 9 9 1 9 9 9 1 13 4 4 9 12 12 9 9 1 11 9 9 1 2 9 1 9 1 1 9 9 1 13 4 2 9 1 9 2 1 14 13 4 4 9 1 13 4 4 9 1 13 2
25 9 7 11 9 9 1 2 3 2 9 0 2 1 1 13 4 4 9 1 0 13 4 16 4 2
22 3 2 9 9 1 13 9 9 4 9 5 9 9 1 9 1 9 1 0 13 4 2
44 11 1 9 9 1 2 9 9 1 9 1 13 4 4 9 1 9 9 1 1 2 9 9 1 9 1 13 2 9 1 9 1 13 4 2 1 1 9 1 13 4 16 4 2
26 9 9 7 9 9 1 3 9 1 9 1 13 9 1 1 2 10 4 4 9 1 9 1 0 4 2
23 11 9 1 9 9 1 1 2 3 2 15 1 13 4 16 4 9 1 9 1 13 4 2
37 11 9 1 11 9 2 9 1 9 9 1 9 9 1 9 1 13 16 1 9 9 1 13 4 4 9 4 2 9 1 9 1 13 4 4 4 2
16 7 9 1 9 9 1 13 16 2 9 1 9 1 13 4 2
21 3 2 9 9 1 13 9 2 11 9 1 9 9 1 0 4 13 4 4 4 2
14 7 2 9 4 9 1 0 4 13 9 1 13 4 2
20 3 13 4 16 4 9 1 2 9 9 1 13 9 1 9 1 13 14 4 2
14 9 9 1 9 1 2 9 1 9 1 13 4 4 2
34 9 9 1 9 1 13 9 9 1 1 2 9 13 9 1 13 16 2 15 1 9 9 1 13 4 16 2 9 1 13 4 4 4 2
33 9 12 1 2 9 9 1 9 1 13 4 14 4 1 4 2 9 9 1 9 1 13 4 9 1 9 1 13 16 4 9 4 2
23 11 1 0 9 9 1 9 1 3 9 13 9 2 9 9 9 1 13 4 4 4 4 2
39 9 12 1 2 9 9 1 4 4 9 9 1 13 16 1 13 4 4 2 9 9 9 1 13 4 4 1 13 9 9 1 9 1 13 4 16 4 4 2
19 9 9 1 9 9 1 9 1 0 9 1 13 9 1 9 9 1 13 2
43 10 9 1 9 1 2 9 1 1 12 12 12 9 14 14 13 4 4 9 1 9 1 3 13 4 16 2 11 1 4 4 9 1 9 1 10 9 2 13 4 9 4 2
37 0 4 9 1 2 9 9 1 1 3 9 9 9 1 9 1 9 1 13 16 4 2 9 9 1 9 9 1 9 1 13 9 1 0 9 4 2
56 9 9 9 1 9 2 9 9 1 9 1 9 1 13 1 13 16 1 2 0 9 1 13 4 9 9 9 1 13 16 1 2 0 4 0 9 9 1 9 1 13 1 13 4 9 1 9 9 1 13 4 4 4 4 14 2
52 11 9 1 13 4 9 9 9 1 1 2 11 9 7 11 9 7 1 9 9 9 1 9 1 9 1 13 2 9 9 9 1 0 4 9 9 9 9 14 1 9 1 13 4 4 2 9 1 13 4 4 2
37 9 1 2 9 9 1 9 9 7 9 9 1 1 9 1 13 4 9 1 9 7 2 0 4 9 9 1 9 7 1 13 4 4 16 4 4 2
11 9 1 9 9 9 1 9 9 4 4 2
33 9 1 9 9 1 9 1 2 9 1 13 16 13 16 9 9 1 13 4 9 1 13 4 4 2 0 1 9 1 0 4 4 2
64 13 16 2 11 1 13 4 4 9 9 9 1 9 2 13 4 4 16 2 10 9 1 13 9 9 2 9 7 2 9 1 9 9 1 9 1 13 1 13 2 9 5 11 1 3 15 1 13 16 4 4 16 14 2 1 1 9 1 13 4 1 13 4 2
21 9 9 9 1 9 9 1 0 4 4 9 2 9 1 13 16 4 4 16 14 2
22 7 2 9 9 1 13 4 9 9 1 9 1 13 9 1 1 15 4 4 16 14 2
13 9 1 13 16 2 15 1 13 4 9 1 0 2
49 12 12 12 12 9 2 11 1 9 7 9 7 1 9 9 1 13 4 16 9 2 9 9 1 9 1 9 4 13 2 9 1 9 1 2 9 7 9 9 1 13 16 11 1 13 4 16 4 2
23 9 9 9 1 1 2 9 1 9 11 1 2 9 1 13 2 9 4 4 4 16 14 2
15 9 4 2 9 1 9 1 13 9 1 13 16 1 13 2
14 9 9 1 11 11 9 1 0 9 1 13 16 4 2
21 12 9 9 2 2 9 9 1 9 1 13 9 2 1 13 4 9 1 9 4 2
41 2 9 1 13 4 4 16 2 0 1 9 1 3 9 1 14 1 13 4 2 11 9 14 4 4 2 3 9 1 9 9 1 13 4 1 13 16 4 9 4 2
25 11 9 1 9 9 9 7 9 9 1 13 2 9 9 9 9 9 2 1 0 9 1 12 9 2
23 9 9 1 13 16 1 9 1 0 4 9 1 0 4 13 16 4 16 4 1 4 14 2
36 0 4 9 9 1 2 13 16 1 13 9 1 4 4 2 0 9 1 13 16 4 4 2 1 13 4 16 1 9 1 0 9 1 13 4 2
16 9 1 13 16 9 1 13 4 1 13 4 4 16 4 4 2
18 11 12 12 9 1 13 16 2 9 9 1 9 1 9 1 13 4 2
26 11 12 12 12 9 2 11 11 9 1 2 11 1 9 9 9 2 1 13 4 16 9 1 13 4 2
20 11 1 9 1 2 9 14 9 9 1 13 4 4 2 1 13 9 4 4 2
18 10 9 9 1 13 4 4 9 4 2 0 4 9 9 1 13 4 2
41 10 9 1 1 3 9 1 0 4 4 9 1 2 9 1 9 9 2 11 11 9 9 1 13 4 2 9 1 13 4 2 9 9 2 1 1 9 9 4 4 2
50 9 12 9 1 9 2 9 2 9 1 9 9 1 13 2 9 12 9 1 9 2 9 9 1 13 2 9 9 1 12 12 12 12 12 9 1 13 9 1 13 16 1 0 4 9 1 9 4 4 2
40 9 9 4 12 12 9 1 13 1 13 9 1 9 1 13 4 2 9 1 9 1 0 9 13 4 16 2 11 9 1 9 1 3 9 1 13 16 4 4 2
47 9 9 1 9 9 9 13 4 1 13 4 16 14 2 9 1 11 12 12 12 9 1 9 2 12 12 12 9 1 11 1 9 7 9 9 1 9 9 2 1 13 9 1 13 16 4 2
34 12 9 9 2 12 9 1 9 1 13 4 16 2 10 9 1 13 4 4 4 16 1 2 9 9 1 2 9 9 9 2 4 4 2
22 10 9 1 0 4 4 4 16 1 2 9 11 9 9 1 13 16 4 9 4 4 2
56 9 1 9 9 9 1 1 3 9 4 9 1 9 1 13 4 9 1 11 9 9 7 11 1 1 9 1 13 4 4 1 13 9 1 2 0 4 15 14 1 9 9 1 12 9 9 1 13 4 9 1 13 4 4 4 2
15 10 9 14 1 9 9 1 1 9 14 1 9 1 13 2
20 9 1 9 1 1 3 9 9 9 1 13 16 2 15 1 9 1 13 4 2
13 9 9 9 1 13 2 9 2 9 1 13 4 2
32 9 1 0 4 13 4 16 1 0 16 2 9 9 1 9 9 1 13 4 4 2 9 1 9 9 13 4 9 1 13 4 2
24 11 12 12 9 1 12 12 9 1 13 16 2 9 9 1 13 9 1 9 4 3 13 4 2
21 10 9 1 2 11 1 1 9 9 1 3 13 2 9 1 14 13 16 4 4 2
33 9 5 9 9 1 0 9 13 2 9 9 9 14 0 9 1 9 1 13 4 2 9 1 9 1 13 4 1 13 9 4 4 2
13 15 1 13 16 9 9 1 3 9 1 13 13 2
35 9 9 1 1 2 11 12 9 9 2 9 9 12 9 1 9 1 2 9 9 1 9 2 9 7 9 9 1 9 2 1 13 4 4 2
31 15 1 13 16 11 12 9 9 2 9 9 1 0 9 9 4 4 2 9 9 9 9 9 2 1 9 9 1 13 4 2
32 9 1 9 9 1 2 9 9 1 9 1 13 9 2 1 13 4 4 2 9 9 9 9 9 1 9 1 13 4 4 4 2
12 9 9 1 9 11 1 9 9 1 13 4 2
49 10 9 1 1 2 11 9 9 1 9 14 4 4 2 15 9 2 11 1 9 2 1 13 11 9 1 9 9 1 9 1 1 2 9 9 1 0 4 1 13 16 4 16 1 0 9 4 4 2
32 15 14 1 9 9 1 9 1 13 16 4 16 2 11 12 12 9 14 1 2 9 1 3 2 9 9 13 4 2 4 4 2
20 10 9 2 9 9 9 1 2 9 9 9 2 1 9 1 13 16 4 4 2
24 9 9 1 1 9 9 1 9 12 9 9 9 1 13 2 9 14 1 9 1 13 9 4 2
14 10 9 2 3 9 9 1 9 1 13 9 1 13 2
35 9 1 11 9 1 9 1 1 9 1 0 9 1 13 4 2 10 9 9 4 13 16 4 4 9 9 9 1 3 0 4 13 16 4 2
11 3 9 9 1 9 9 1 13 4 4 2
44 9 9 2 9 1 13 4 2 9 9 1 9 1 13 9 9 2 1 2 2 9 9 9 1 9 2 1 13 16 3 0 4 9 1 2 9 1 9 9 1 9 4 4 2
29 7 2 9 5 9 9 7 9 9 1 9 1 2 9 9 13 16 1 0 4 9 1 13 2 1 13 9 4 2
29 15 9 1 15 14 1 13 4 16 4 4 4 4 2 9 9 1 1 3 0 1 0 4 9 1 9 1 13 2
25 9 9 7 2 9 4 9 1 13 16 1 2 3 1 15 14 1 9 1 9 1 13 16 4 2
29 10 9 1 13 16 2 3 9 9 1 13 16 4 4 11 11 5 9 9 9 9 1 9 1 9 1 1 4 2
19 9 9 9 1 9 1 9 1 2 9 14 9 1 13 4 16 4 4 2
15 15 1 11 9 1 3 13 14 2 1 13 9 4 4 2
45 9 9 1 9 9 1 3 13 4 4 9 1 2 11 9 9 2 11 9 9 1 13 0 9 1 9 1 13 9 1 2 11 1 9 1 13 16 1 3 14 1 13 9 4 2
17 9 1 13 4 16 2 11 1 9 1 9 9 1 13 16 14 2
22 9 1 9 1 13 14 3 14 13 4 16 2 9 1 13 16 4 9 1 0 4 2
24 9 1 13 2 9 1 13 4 9 9 4 4 16 1 9 1 9 1 0 0 9 1 13 2
27 9 1 9 1 9 1 13 4 4 2 12 12 12 12 9 9 1 0 9 1 13 4 4 9 1 0 2
25 9 12 12 9 1 11 1 13 4 11 9 1 13 9 2 12 9 1 9 9 1 13 4 4 2
14 9 9 9 1 11 11 5 9 9 9 9 4 4 2
8 3 12 12 9 1 13 4 2
40 11 9 9 9 1 12 12 12 12 9 2 9 12 9 1 11 9 1 9 1 13 4 4 9 1 13 2 9 9 9 9 0 9 9 1 9 1 13 4 2
18 11 9 1 9 12 12 9 9 1 13 4 1 9 1 13 16 4 2
15 9 9 1 1 2 9 9 1 9 2 1 13 4 4 2
24 2 9 9 1 13 4 2 1 13 9 1 13 2 9 9 1 13 9 1 9 1 13 4 2
17 2 9 9 1 13 14 1 1 9 2 1 13 9 9 4 4 2
49 9 1 2 11 9 1 9 1 9 1 13 16 9 9 1 13 9 9 1 13 16 4 0 4 9 9 2 1 13 4 11 9 1 2 13 4 4 9 1 9 1 9 1 13 4 2 1 13 2
34 9 1 9 1 13 4 16 2 9 9 13 4 9 1 9 1 12 9 1 13 4 9 9 9 2 0 9 14 1 3 1 13 4 2
10 11 1 13 9 9 1 13 4 4 2
17 12 12 9 1 9 1 1 12 12 12 9 9 1 13 4 4 2
45 12 12 9 1 12 12 9 14 1 11 2 9 9 2 11 2 9 2 11 9 1 9 12 9 9 1 9 1 9 13 4 4 16 2 9 9 1 9 3 13 4 4 4 4 2
14 9 2 9 9 1 9 9 13 4 4 4 13 4 2
18 10 9 1 11 9 1 0 9 1 13 2 9 9 1 13 4 4 2
23 9 9 9 1 9 1 13 4 2 9 9 2 9 2 9 9 9 14 1 13 4 4 2
16 2 9 9 1 9 9 1 9 2 1 13 9 1 13 4 2
24 9 1 13 2 9 1 9 1 13 4 9 1 13 9 1 0 4 9 4 13 16 4 4 2
57 9 9 9 9 9 1 11 11 5 11 9 1 9 1 9 1 2 11 9 9 2 11 9 1 9 9 1 13 4 9 1 1 4 2 12 12 9 1 11 9 9 9 14 9 1 9 1 13 4 16 1 13 4 1 13 4 2
21 9 9 4 0 4 9 1 9 13 4 9 1 1 0 9 1 13 4 4 4 2
33 11 9 9 1 9 7 9 1 13 4 9 9 1 13 4 2 9 1 1 9 1 13 4 16 2 9 9 1 9 1 13 4 2
25 9 9 9 1 9 9 9 1 15 13 16 1 0 4 16 2 9 1 0 4 13 4 4 4 2
24 9 7 9 1 9 1 1 2 3 9 1 13 16 1 3 14 2 1 13 9 1 0 4 2
26 11 9 1 2 9 9 1 9 2 1 13 4 9 1 2 0 4 2 1 13 4 9 1 13 4 2
22 3 14 2 11 1 1 9 9 1 13 4 2 1 13 9 9 4 9 1 13 4 2
17 10 9 1 9 9 9 1 13 13 4 4 11 9 1 13 4 2
20 9 7 9 9 1 0 4 9 1 13 4 1 9 9 1 9 1 13 4 2
18 9 1 13 4 9 1 2 9 1 13 4 9 1 9 1 13 4 2
25 9 9 9 4 9 1 13 4 11 1 11 9 1 0 9 1 13 4 9 1 9 1 13 4 2
21 0 9 9 1 13 2 9 1 1 9 1 9 1 13 4 9 4 16 5 5 2
12 9 4 9 9 1 9 1 9 1 13 4 2
7 3 9 1 13 4 4 2
26 9 1 9 9 9 1 9 9 1 9 1 13 16 9 1 9 9 1 13 4 1 13 11 1 13 2
40 9 1 1 13 4 11 9 1 11 9 9 1 9 1 13 2 9 9 1 1 13 9 9 9 9 9 1 13 4 1 13 16 1 11 9 1 9 4 4 2
9 3 9 1 13 16 1 4 4 2
13 9 1 0 9 9 1 0 4 13 9 1 13 2
23 9 1 9 7 0 9 1 13 9 1 9 9 1 0 4 9 1 11 9 1 13 4 2
21 9 1 9 1 9 9 1 9 1 13 4 11 9 1 9 1 9 1 13 4 2
15 9 1 13 4 1 1 0 4 9 9 7 9 1 13 2
12 7 3 13 9 9 9 1 13 4 4 4 2
52 9 1 9 9 1 13 4 4 9 9 1 9 1 13 4 16 9 1 9 9 14 9 2 15 1 9 9 1 13 16 4 14 14 1 9 1 13 2 9 9 1 9 7 9 9 1 13 1 13 9 4 2
54 15 1 13 11 9 1 2 11 7 11 5 9 14 1 1 9 1 13 4 2 11 9 1 9 1 13 2 9 9 9 1 9 1 13 4 14 9 9 1 13 4 9 9 9 1 3 13 9 1 0 4 1 13 2
12 9 9 1 9 1 1 3 9 1 13 4 2
40 12 12 5 12 12 9 1 11 9 5 11 9 9 1 9 2 9 1 9 1 2 9 9 0 16 1 9 1 9 4 2 1 13 9 1 9 1 1 13 2
33 9 9 7 9 9 1 9 1 13 9 9 7 2 9 1 9 9 1 9 1 13 9 9 1 9 1 9 1 13 9 1 13 2
61 11 11 5 11 9 9 1 2 15 14 9 2 9 2 9 9 2 9 14 1 9 9 1 9 1 9 0 1 0 4 9 1 13 16 4 4 9 1 2 9 1 9 1 0 13 4 9 1 9 1 1 4 14 2 1 9 1 13 16 13 2
25 9 1 0 9 1 13 2 9 9 1 13 4 4 9 1 9 1 13 9 1 9 1 1 13 2
29 11 9 1 4 4 9 13 9 1 13 4 9 1 13 9 2 9 9 1 3 13 4 9 1 13 16 4 4 2
22 9 9 9 9 1 9 9 12 9 1 0 4 9 9 9 9 1 9 9 13 4 2
58 9 1 13 9 9 1 2 12 12 12 12 9 1 9 9 9 9 12 9 9 2 12 12 9 1 9 1 13 16 9 1 9 9 9 1 9 1 13 16 9 9 1 9 9 4 13 9 1 13 4 16 9 12 9 9 4 4 2
33 12 9 1 9 9 1 9 9 9 1 9 9 9 1 9 1 13 2 9 1 13 16 9 9 1 13 4 16 4 4 1 13 2
33 9 1 3 9 1 13 4 16 4 4 1 13 4 4 16 2 9 1 9 1 0 4 12 12 9 9 1 13 16 13 4 4 2
36 9 1 13 9 9 1 2 9 9 1 9 9 1 0 4 9 1 13 2 7 9 1 13 4 1 13 4 0 4 9 1 13 16 13 4 2
22 10 9 1 13 16 1 9 1 9 1 3 0 4 4 2 9 9 1 9 4 13 2
29 9 1 1 2 11 1 9 9 1 13 2 9 9 4 1 9 1 13 4 4 9 9 1 9 1 13 16 4 2
19 9 0 9 1 2 9 9 4 1 9 9 4 1 0 9 9 1 13 2
21 0 9 1 9 1 9 9 1 13 4 9 1 2 0 13 4 4 16 4 4 2
34 9 1 3 12 12 9 9 1 13 4 16 4 4 1 13 16 2 11 1 9 9 9 1 12 12 9 1 9 1 0 13 4 4 2
35 9 9 1 9 1 13 4 2 9 9 1 13 9 9 7 9 9 1 13 4 4 2 9 13 4 4 4 9 9 1 13 4 4 4 2
23 15 1 13 2 2 9 2 1 13 16 1 9 7 9 1 1 9 1 13 4 9 4 2
29 0 9 4 2 3 9 1 13 16 4 4 9 1 2 0 9 9 1 13 9 4 4 1 13 4 1 13 4 2
46 9 4 9 1 2 9 9 4 4 9 9 9 9 1 9 1 13 4 7 2 9 1 9 9 7 9 9 9 1 9 9 1 13 4 7 4 16 4 4 9 1 0 4 9 4 2
16 9 1 9 1 13 4 9 1 13 16 13 4 9 4 4 2
21 9 1 2 9 9 1 15 1 13 4 14 1 9 1 9 1 13 4 16 4 2
29 15 9 1 2 11 1 9 9 4 9 1 13 16 10 4 4 9 9 1 13 4 4 9 1 3 0 4 13 2
20 10 9 1 11 1 9 9 1 9 9 1 3 0 9 14 1 13 16 4 2
45 9 9 9 1 13 16 13 4 16 1 9 1 9 1 13 4 9 9 1 1 9 1 9 1 0 13 4 16 4 1 9 4 1 1 9 1 2 0 16 13 9 1 13 4 2
24 0 9 1 13 4 9 1 1 2 9 1 1 9 9 1 3 13 4 9 1 0 4 4 2
58 9 9 1 9 1 13 4 16 12 12 9 1 13 4 16 2 11 1 12 12 9 1 13 16 0 2 7 11 1 1 9 9 12 12 9 1 1 9 9 1 13 4 16 4 16 2 11 1 1 12 9 1 12 9 1 13 4 2
23 9 9 1 0 9 1 9 9 2 3 9 1 9 1 9 9 4 13 4 9 4 4 2
17 7 2 3 0 4 16 1 2 9 9 9 1 9 9 4 4 2
36 9 1 9 1 2 9 1 9 4 4 2 0 4 0 4 9 2 1 13 9 1 11 1 9 9 1 1 2 3 13 4 9 1 13 4 2
36 9 9 1 15 1 1 9 9 9 1 9 4 4 2 9 1 9 1 13 4 9 1 9 9 1 9 1 9 1 0 4 13 4 4 4 2
43 3 2 11 1 9 9 9 1 9 1 9 1 9 9 4 0 13 2 9 9 1 9 4 4 2 0 4 0 4 9 2 1 13 16 2 3 9 1 13 4 13 4 2
35 12 12 12 1 9 2 12 12 12 1 9 1 13 11 1 9 2 9 11 11 9 2 1 13 9 0 4 9 1 9 1 13 16 4 2
66 12 9 13 4 4 11 9 9 9 9 1 1 9 9 9 1 2 10 9 0 4 9 1 9 1 2 9 9 9 2 11 11 9 9 2 9 12 9 2 9 9 1 15 14 9 1 9 4 9 1 13 4 4 1 13 16 4 9 1 13 4 9 1 13 4 2
35 9 1 13 9 1 2 3 9 9 9 2 11 11 9 1 13 4 16 4 4 4 4 0 4 9 9 9 7 0 9 9 1 1 4 2
54 9 1 9 2 9 9 2 9 2 9 1 9 14 3 13 4 16 4 9 9 1 9 1 9 1 13 2 9 1 1 9 1 13 2 3 0 4 9 2 3 9 1 13 4 9 9 1 13 4 1 13 16 4 2
38 11 9 1 9 12 9 9 1 12 12 9 9 1 0 9 1 13 2 9 1 13 2 9 9 9 1 12 12 12 12 9 1 9 9 4 13 4 2
8 9 1 9 1 9 9 4 2
50 11 11 9 1 9 1 9 9 9 1 12 5 12 9 1 9 1 9 1 9 4 13 2 9 9 9 1 13 16 1 12 12 9 1 9 0 4 9 1 13 4 9 1 9 4 9 1 13 4 2
51 9 9 9 9 9 1 13 16 1 2 9 9 14 1 9 9 4 13 4 9 1 13 4 4 16 2 3 15 1 0 4 9 1 13 1 1 3 12 2 12 12 9 1 13 1 9 9 1 9 4 2
27 13 4 2 3 2 11 1 9 1 1 13 4 9 9 9 1 13 4 2 13 4 4 1 13 9 4 2
22 9 9 1 13 16 1 9 9 1 9 4 4 2 9 1 0 9 1 3 13 4 2
25 9 1 9 1 9 9 13 4 4 16 4 4 9 9 1 9 1 13 4 1 1 13 16 4 2
42 9 1 9 9 1 9 9 9 1 13 16 1 2 9 1 13 9 9 9 14 0 9 1 13 4 1 13 16 4 16 2 3 9 1 12 9 9 1 13 1 13 2
31 9 1 9 1 1 0 4 2 9 9 9 1 9 2 1 13 4 16 4 16 1 9 9 1 13 4 16 14 13 4 2
20 3 1 1 9 4 16 9 9 1 9 9 13 9 1 13 16 4 16 4 2
42 15 14 1 9 9 9 9 1 9 9 9 1 13 0 9 9 9 1 13 4 4 14 1 2 9 9 1 9 1 11 9 1 0 4 9 1 9 1 13 4 4 2
15 9 9 1 13 16 9 9 1 1 9 1 9 1 13 2
53 10 9 9 9 1 1 9 9 9 1 1 9 1 9 1 13 9 2 9 1 13 4 4 9 2 9 9 9 1 1 9 1 13 4 9 1 3 0 13 4 16 4 2 9 9 1 9 1 0 4 13 4 2
26 11 11 9 1 2 9 1 9 1 9 2 9 1 0 4 13 2 9 1 9 9 1 9 1 13 2
45 12 12 12 9 14 1 9 12 9 2 11 1 2 9 11 11 9 2 1 9 1 0 4 13 2 0 4 9 13 16 13 4 16 4 9 1 2 9 9 1 13 16 1 0 2
24 10 9 1 1 11 11 9 1 13 9 9 2 9 9 9 1 9 9 4 13 4 16 4 2
10 7 9 9 1 0 9 1 1 4 2
15 9 1 13 9 9 1 9 1 3 13 4 4 9 4 2
10 9 1 9 1 1 0 4 9 4 2
35 11 7 11 14 9 9 1 9 9 1 13 11 9 9 1 9 1 13 16 4 16 4 1 13 16 9 1 13 4 9 1 13 14 4 2
27 11 1 3 1 9 4 4 2 9 9 5 9 9 2 1 9 9 1 13 16 9 9 1 13 4 4 2
36 9 5 11 1 2 9 1 9 2 9 4 13 4 2 3 9 1 1 2 9 1 13 0 0 13 9 1 9 9 2 4 16 4 4 14 2
63 9 1 13 4 9 9 9 9 1 9 1 11 5 11 9 9 9 4 16 2 10 9 9 9 1 13 4 9 1 9 1 9 1 9 1 13 4 9 2 9 2 7 2 9 9 9 2 9 1 13 16 4 4 1 14 13 9 1 0 16 4 4 2
51 11 9 1 1 11 11 9 9 9 9 1 9 14 9 9 1 9 9 1 13 16 13 4 9 1 3 9 2 11 9 1 1 9 9 9 9 1 9 1 13 4 9 1 9 1 13 16 4 16 4 2
26 9 1 1 13 9 9 9 1 1 3 0 9 9 1 13 9 1 13 0 1 13 4 16 4 4 2
47 7 1 11 9 1 9 1 9 9 1 9 1 9 9 1 13 16 4 16 4 2 11 9 1 4 4 9 9 1 9 1 13 0 9 1 9 1 9 1 13 1 13 9 1 9 13 2
48 7 2 3 9 9 9 1 13 4 9 4 1 4 16 2 3 14 9 9 1 0 4 9 1 13 4 4 16 1 9 1 13 4 16 9 1 13 9 1 1 9 9 1 1 14 13 4 2
83 11 9 1 9 2 3 1 9 9 13 4 16 1 9 9 1 11 11 5 11 9 9 4 4 16 2 9 2 11 11 5 11 9 1 9 9 2 11 11 5 11 9 11 9 9 9 2 11 11 9 9 9 2 11 11 9 9 9 1 3 1 9 1 13 2 9 1 11 11 5 9 9 1 9 9 1 9 14 13 16 4 4 2
37 12 12 9 13 14 1 9 4 16 2 9 9 1 9 9 1 1 9 9 1 9 1 1 9 4 13 4 4 1 1 9 14 1 13 4 4 2
58 3 11 1 13 9 9 12 9 1 9 1 2 9 2 9 14 12 9 1 9 1 13 4 9 2 0 9 9 1 13 4 9 1 1 9 1 9 1 2 13 9 2 9 1 13 2 9 9 1 15 1 13 4 4 4 4 4 2
24 7 1 11 9 1 1 2 3 0 4 2 9 9 9 9 2 9 1 9 1 13 4 4 2
24 3 9 1 9 1 11 11 9 1 13 4 4 16 2 9 9 1 9 13 9 13 1 9 2
39 13 4 16 9 9 9 1 9 9 1 11 11 9 9 1 9 1 9 14 13 4 16 2 9 9 1 9 1 14 13 4 4 4 9 1 13 16 4 2
17 2 9 9 0 2 1 2 9 9 12 9 2 1 13 16 0 2
69 9 1 13 9 1 9 1 9 1 9 1 13 16 0 4 13 4 9 1 2 12 9 9 1 11 9 9 1 2 9 11 9 2 1 13 4 4 11 11 9 1 9 9 12 9 9 9 1 13 4 9 1 9 1 2 9 9 9 14 13 1 9 1 9 1 0 14 4 2
55 12 9 9 1 9 1 11 1 2 3 9 9 1 13 16 2 9 9 1 1 13 4 14 13 4 2 1 1 9 1 2 9 13 4 9 1 9 1 13 4 4 4 16 2 10 9 1 0 4 16 4 1 4 14 2
27 15 1 9 14 1 9 1 9 14 1 2 0 1 9 9 1 1 9 1 9 1 9 1 13 4 4 2
33 9 13 9 1 0 16 2 0 9 9 9 1 1 9 2 9 1 9 1 9 13 4 16 4 2 9 9 1 9 1 9 4 2
28 2 13 9 2 2 9 13 9 2 13 1 2 9 12 9 1 9 7 9 1 9 1 0 4 4 9 4 2
13 10 9 1 9 1 9 14 13 4 16 1 0 2
17 3 3 9 9 1 13 1 13 4 16 2 3 9 1 13 4 2
18 9 1 1 3 9 9 1 13 2 9 9 9 1 13 4 16 4 2
26 9 9 1 1 4 2 2 9 9 9 4 2 2 9 1 9 9 4 2 1 13 16 1 13 4 2
31 9 9 12 9 9 5 9 9 1 15 1 9 13 16 14 1 13 16 2 3 11 1 9 1 13 16 4 9 4 4 2
9 11 1 9 9 1 13 16 4 2
31 11 1 9 1 9 9 1 9 1 2 9 1 2 9 9 2 1 13 16 1 2 9 9 1 9 9 1 9 1 13 2
29 12 12 9 0 9 9 1 9 9 1 9 9 1 13 4 16 2 9 9 1 9 1 13 9 1 13 4 4 2
31 15 1 10 9 4 2 9 9 1 13 16 2 12 9 1 9 9 1 9 1 9 1 9 1 12 12 9 1 1 13 2
30 9 9 1 12 9 1 12 12 9 2 12 12 12 9 9 1 9 1 13 16 1 2 9 1 13 4 9 1 0 2
34 9 1 9 1 0 1 13 16 2 9 9 9 1 9 9 14 0 16 2 11 1 11 9 9 1 9 1 9 1 13 16 1 0 2
9 11 1 9 1 13 9 1 0 2
20 9 2 11 1 9 9 9 1 2 9 13 9 9 9 4 9 4 4 4 2
29 7 2 9 9 1 9 1 1 2 9 9 1 9 1 13 2 13 4 16 4 16 1 9 1 1 11 1 13 2
20 9 1 13 1 1 2 11 1 9 9 2 9 9 1 13 4 16 4 4 2
12 7 2 9 9 1 13 4 4 16 4 4 2
17 7 2 9 9 1 9 4 2 3 13 16 1 13 4 1 4 2
27 12 12 12 9 9 1 9 7 9 7 1 9 9 1 13 4 16 9 2 9 1 9 9 1 13 4 2
27 9 9 1 13 16 9 1 13 4 16 9 1 9 1 13 16 4 9 2 9 1 9 1 9 4 4 2
38 12 9 9 1 9 1 11 9 1 9 9 13 4 9 2 9 9 1 9 1 9 1 9 1 13 2 9 9 1 9 1 9 1 9 4 13 4 2
25 9 9 1 9 2 9 2 9 1 13 4 9 2 11 9 1 9 1 9 1 13 4 9 4 2
35 7 2 9 1 9 1 13 4 2 15 1 9 14 1 2 9 9 1 9 9 13 2 9 9 1 13 9 1 13 9 4 16 4 4 2
23 9 9 1 9 1 2 3 11 1 9 1 13 16 4 2 11 1 1 9 1 13 4 2
30 12 9 9 1 9 9 1 9 1 2 12 9 5 12 12 12 9 4 4 9 9 1 2 12 12 9 14 13 4 2
28 7 2 10 9 2 9 9 9 1 3 13 4 2 9 1 0 9 1 0 9 1 9 1 13 16 4 4 2
13 10 9 1 9 2 9 9 9 13 16 1 13 2
19 9 1 13 9 0 2 9 9 9 1 9 1 9 14 1 13 16 4 2
15 9 9 2 9 9 1 11 1 9 1 0 4 4 13 2
54 7 2 12 12 12 12 9 9 1 9 9 1 13 16 2 11 9 1 0 9 9 2 9 9 1 9 1 2 9 1 12 12 9 9 1 13 4 2 9 1 9 9 13 16 2 9 9 1 13 4 9 1 13 2
31 2 9 9 1 9 2 1 13 16 2 13 4 4 16 7 2 9 9 4 9 9 1 13 4 4 9 4 16 4 4 2
42 11 1 10 9 2 9 1 13 4 9 2 9 9 1 9 1 2 11 2 11 1 9 1 13 4 2 9 1 13 4 4 9 9 9 1 9 1 13 4 16 4 2
24 11 1 9 9 1 13 4 16 2 12 12 12 9 1 1 2 9 1 13 4 9 13 4 2
8 9 1 10 9 9 1 13 2
30 11 7 11 2 11 1 12 9 1 12 9 2 9 1 9 9 1 13 4 9 9 9 9 1 0 4 13 4 4 2
39 9 9 1 13 4 9 9 1 9 9 9 1 2 11 1 5 5 9 9 1 1 9 7 9 1 9 9 9 9 1 13 4 2 1 13 4 16 4 2
13 9 9 1 2 10 9 1 13 13 4 4 4 2
20 9 9 9 1 0 4 9 1 13 16 2 9 9 1 9 1 13 4 4 2
32 9 9 9 1 1 2 9 9 9 1 9 12 12 12 9 14 1 2 13 4 4 4 13 4 2 1 2 13 4 16 4 2
32 10 9 11 1 9 1 13 4 2 11 1 9 9 9 1 13 4 16 4 4 16 2 9 1 1 9 1 13 4 1 0 2
37 15 1 2 11 9 1 9 9 9 1 9 1 13 4 9 1 2 9 9 4 9 9 1 13 4 4 16 4 4 2 11 1 9 1 13 4 2
43 9 1 9 1 13 16 1 2 2 11 9 2 1 13 4 9 9 9 11 1 13 2 11 1 2 11 9 1 9 9 1 9 1 13 2 1 13 16 13 4 16 4 2
26 7 2 11 1 9 1 9 1 13 4 9 2 9 9 4 1 2 11 1 11 9 1 13 9 4 2
31 7 2 9 9 9 14 1 9 1 13 9 1 9 1 13 16 2 13 4 16 4 1 13 4 1 13 16 4 4 4 2
20 7 2 9 9 9 1 9 9 9 1 13 1 1 2 7 9 1 13 4 2
12 9 9 9 14 9 1 13 4 14 13 4 2
29 11 1 2 9 14 1 9 1 13 4 16 2 9 9 1 9 9 5 9 9 14 1 13 4 16 4 4 4 2
17 11 1 9 1 2 9 9 9 1 9 1 13 4 9 4 4 2
16 7 2 11 9 1 9 1 9 1 0 4 9 1 1 4 2
17 7 3 13 4 4 16 4 4 9 1 2 0 4 13 16 4 2
21 3 2 9 9 9 1 9 1 2 11 7 11 1 13 4 9 1 13 16 4 2
14 3 11 1 9 9 1 9 1 13 4 4 16 14 2
16 11 9 1 11 1 9 9 1 13 4 4 16 4 4 14 2
22 9 9 9 1 1 11 1 9 9 1 2 12 12 12 9 9 1 13 4 16 4 2
6 0 4 9 4 4 2
23 10 9 1 2 11 1 1 9 4 16 14 9 9 4 16 14 1 3 0 4 1 4 2
25 15 1 13 16 1 2 2 11 1 9 9 1 9 1 9 2 1 13 4 4 16 4 14 4 2
36 11 1 2 9 9 1 13 4 9 9 1 9 1 13 16 9 1 0 1 13 16 4 2 11 1 13 1 13 4 9 9 1 9 4 4 2
14 10 9 9 1 1 13 4 4 4 1 4 4 14 2
44 11 1 11 9 9 1 2 11 1 1 9 9 1 13 16 2 9 1 13 9 9 1 13 9 1 9 9 1 1 13 4 2 9 1 13 4 4 9 1 13 4 16 4 2
41 9 1 2 9 11 1 9 9 7 9 1 13 4 9 11 9 1 0 4 13 2 11 9 1 0 4 4 13 4 16 14 2 9 1 3 13 4 4 4 4 2
22 0 9 1 13 2 9 1 13 2 9 1 13 16 9 1 9 7 9 1 13 4 2
16 15 1 9 9 1 9 1 9 1 9 1 13 9 4 4 2
25 11 1 9 11 1 11 1 9 9 1 2 9 9 9 2 1 9 1 15 9 1 0 13 4 2
40 9 12 12 12 9 1 9 9 1 13 9 9 1 12 9 1 2 9 2 1 2 9 9 2 1 9 1 13 2 12 12 9 1 9 9 1 13 4 4 2
35 11 11 9 1 2 3 13 4 2 9 1 0 9 2 1 0 4 4 9 9 1 13 9 14 1 2 9 9 1 0 4 13 16 4 2
39 9 9 1 9 9 1 13 4 4 9 9 9 1 2 9 1 1 9 1 11 1 9 1 13 16 2 0 9 1 9 9 1 0 4 13 16 4 4 2
42 9 9 1 1 9 1 9 1 13 2 9 1 9 1 13 2 9 9 4 9 1 9 1 13 4 16 4 13 1 0 2 9 1 9 4 9 1 13 9 4 4 2
34 9 9 1 9 7 9 1 9 1 13 2 0 9 2 9 9 2 9 1 9 9 1 1 9 1 9 9 1 1 13 4 16 4 2
68 9 9 1 9 4 13 4 16 4 4 9 9 7 9 2 9 14 1 9 1 13 4 4 12 12 12 12 9 1 2 9 9 9 2 2 12 12 9 1 2 9 9 2 2 12 12 9 1 2 9 9 9 2 7 2 9 9 9 2 1 0 9 1 9 9 4 4 2
30 9 1 9 1 2 9 1 9 4 9 12 1 9 9 1 13 4 9 9 1 9 2 1 13 16 4 16 1 13 2
22 7 2 9 1 12 12 12 12 12 9 1 13 4 2 12 12 9 1 9 1 13 2
15 9 4 9 1 0 2 9 1 9 1 0 4 1 4 2
39 2 9 2 9 1 3 9 2 9 2 9 1 9 1 13 4 16 4 16 1 9 2 9 1 13 2 9 1 9 1 13 16 4 9 4 4 16 4 2
43 9 9 1 9 1 13 16 2 9 1 9 9 7 9 14 9 9 9 1 2 9 9 1 9 9 2 9 9 2 9 14 9 1 9 9 1 13 4 4 13 16 4 2
47 10 9 1 13 16 2 9 9 1 12 12 9 12 12 9 2 2 7 9 9 9 9 1 12 12 9 7 9 1 12 12 9 1 9 9 1 13 4 16 13 2 1 13 4 16 4 2
39 9 1 9 9 1 13 4 2 12 9 9 9 1 3 4 12 9 1 9 9 1 13 4 16 4 9 1 2 3 13 16 4 14 1 13 4 16 4 2
27 9 7 9 9 14 9 9 1 1 9 1 13 9 4 11 1 9 1 9 1 13 4 9 1 13 4 2
12 9 1 9 1 9 9 1 9 9 4 4 2
34 2 9 2 1 9 9 1 2 9 1 13 4 9 9 4 9 1 13 2 9 1 9 4 13 2 9 9 1 13 4 13 16 4 2
12 3 15 9 1 9 1 13 4 16 4 4 2
22 2 9 2 1 9 9 9 1 13 9 9 1 9 1 1 9 1 13 4 16 4 2
36 9 9 9 2 11 1 13 9 1 9 9 9 1 2 9 9 1 13 9 9 7 9 9 1 13 9 9 1 9 1 9 1 13 16 4 2
26 10 9 9 9 4 9 7 9 9 1 9 9 9 1 9 2 9 14 1 13 1 1 9 4 4 2
24 11 1 13 11 2 9 1 9 9 1 13 16 11 1 9 9 1 13 4 16 1 4 4 2
19 9 1 9 1 13 1 1 2 0 4 9 1 13 4 16 1 4 4 2
28 9 1 13 4 2 9 1 13 4 9 1 13 4 16 13 4 2 9 9 1 9 4 13 4 16 4 4 2
64 9 9 1 13 4 4 11 9 2 9 1 9 9 1 13 4 11 9 9 9 9 1 1 9 9 1 12 9 2 9 9 9 9 1 13 4 4 16 2 9 1 13 16 9 2 9 9 1 0 0 14 1 9 1 3 13 4 16 1 3 0 4 4 2
44 9 13 9 1 0 1 9 1 13 4 9 2 9 1 0 2 9 9 7 9 9 1 13 9 1 9 1 9 1 13 16 4 1 2 0 9 1 13 16 1 9 4 4 2
29 0 4 9 9 4 4 2 0 2 9 9 2 1 9 14 13 4 9 9 4 16 9 9 1 9 1 13 4 2
82 9 1 2 9 9 1 13 16 9 12 12 12 12 9 1 1 13 1 13 2 9 9 1 13 4 9 9 1 13 4 9 1 9 1 12 12 12 9 1 13 4 2 11 9 1 12 12 12 9 1 9 9 13 2 7 9 2 9 1 9 1 9 9 1 9 1 13 4 9 1 9 13 1 13 4 2 1 13 9 4 4 2
54 9 1 9 1 9 1 2 9 1 9 9 1 9 9 1 13 4 16 2 9 7 11 1 9 1 9 1 13 4 2 9 1 1 9 9 1 13 4 16 11 9 9 9 1 9 9 1 13 9 9 1 4 4 2
68 7 9 1 9 9 1 13 9 1 3 0 4 4 2 9 9 1 9 1 9 9 1 9 1 13 16 2 3 9 9 1 9 9 1 0 9 1 13 4 16 4 4 16 14 2 9 9 1 9 2 9 9 9 1 9 14 1 13 16 9 1 13 4 9 1 13 4 2
18 9 1 15 1 13 4 2 13 4 4 16 2 0 4 13 4 4 2
39 9 9 9 1 9 9 1 0 13 4 4 16 4 9 2 11 1 13 9 2 9 9 9 1 1 9 1 13 4 4 9 9 1 9 1 13 16 4 2
37 7 2 9 1 9 1 1 11 9 9 1 9 9 9 2 11 11 9 1 1 0 9 9 1 9 1 13 4 16 4 9 1 9 9 1 13 2
42 9 1 9 1 9 1 13 9 9 2 9 9 9 1 13 2 9 1 9 9 1 9 9 9 9 1 9 1 13 4 16 4 2 1 13 16 9 4 9 4 4 2
64 3 9 1 0 9 9 1 1 4 4 16 2 9 9 1 9 9 1 9 1 9 9 4 1 4 16 0 4 13 4 16 2 11 9 7 9 9 2 9 7 1 9 9 1 13 4 9 9 2 9 9 1 9 4 9 1 9 1 0 4 13 4 4 2
51 7 2 9 9 1 9 9 1 13 4 9 1 3 0 4 9 1 13 4 16 14 2 9 1 1 9 9 1 13 16 0 4 9 1 13 4 9 1 9 9 14 9 1 3 13 4 2 1 13 4 2
60 12 12 9 1 1 9 9 9 1 11 11 5 9 11 9 2 11 11 11 9 1 13 9 9 9 1 13 4 4 16 4 16 2 9 1 13 9 1 9 1 13 9 1 1 9 1 1 13 4 4 9 9 1 9 1 13 16 4 4 2
17 9 9 1 9 1 9 9 1 13 16 1 13 4 16 4 4 2
19 9 9 1 9 9 4 4 4 7 9 1 9 9 1 9 9 4 4 2
66 15 9 1 3 9 1 13 9 1 13 2 9 1 13 16 9 9 1 0 4 9 9 1 13 9 1 1 9 9 1 9 9 1 13 4 4 13 4 16 4 4 16 2 9 7 9 1 2 9 1 9 9 2 14 1 13 16 9 1 9 13 4 16 4 4 2
26 9 1 9 1 9 9 1 13 4 4 0 4 9 9 1 9 1 13 4 2 9 1 13 4 4 2
19 11 9 1 9 9 1 1 9 9 1 12 12 12 12 9 1 13 4 2
10 9 9 1 13 16 1 9 9 4 2
12 9 1 1 0 9 1 9 1 9 4 4 2
13 7 2 9 9 1 1 9 9 1 13 16 4 2
22 9 9 1 9 9 1 2 9 7 9 9 1 13 16 4 16 1 0 4 9 4 2
24 2 9 1 9 1 9 2 1 13 9 1 13 9 1 13 16 2 13 4 4 9 4 4 2
29 9 12 9 9 1 2 9 5 9 9 9 7 9 1 9 5 9 1 9 12 12 9 1 9 13 4 16 4 2
54 11 9 1 9 11 2 11 1 11 9 2 9 9 9 2 9 9 14 12 12 12 9 1 13 4 9 9 9 9 1 9 1 13 2 11 9 1 13 9 9 1 9 1 3 9 12 12 12 9 1 13 4 4 2
20 9 1 2 9 9 9 1 13 4 4 9 9 1 9 1 13 16 13 4 2
21 9 9 9 1 2 9 9 2 1 13 4 4 4 9 9 1 1 9 9 4 2
30 9 9 1 0 13 4 2 11 9 14 1 1 2 9 9 1 13 4 9 12 9 9 1 9 1 13 16 4 4 2
28 10 9 2 9 9 9 1 13 12 12 12 9 9 1 13 16 9 12 9 9 1 9 1 13 4 16 4 2
12 3 1 9 1 9 1 13 16 4 9 4 2
26 15 1 9 1 13 4 4 16 4 4 2 9 9 1 9 1 13 16 13 9 1 9 9 13 4 2
26 9 9 1 0 9 7 2 9 7 9 9 1 9 2 9 1 1 9 1 13 4 9 1 13 4 2
19 0 9 1 9 1 2 9 1 9 1 1 9 1 13 4 9 1 13 2
31 7 2 0 9 4 16 9 1 13 13 9 1 13 4 1 13 4 2 9 9 1 9 1 13 4 16 1 3 4 4 2
32 9 9 9 1 2 9 14 4 4 2 9 1 9 9 9 7 9 9 1 13 2 7 9 5 9 1 9 9 1 1 13 2
19 9 9 1 1 9 9 1 9 1 13 4 9 4 9 9 1 13 4 2
14 1 1 13 2 9 1 9 1 13 16 1 4 4 2
27 12 9 9 1 13 16 4 9 1 9 13 4 16 14 2 0 4 9 9 1 9 1 13 4 4 4 2
14 9 9 9 1 13 9 1 0 4 9 1 1 4 2
29 7 2 9 1 1 9 9 9 1 13 4 4 9 1 9 2 9 9 1 9 13 4 4 9 1 9 1 13 2
36 10 9 1 13 4 4 4 16 2 9 1 9 1 13 2 9 9 9 1 12 9 9 13 4 9 1 9 9 13 9 1 9 1 13 4 2
20 2 9 1 13 16 2 9 1 9 1 13 16 0 4 2 1 1 9 4 2
14 9 9 1 9 1 13 4 0 4 9 1 13 4 2
24 9 9 9 1 2 9 9 12 9 9 1 13 16 13 2 9 9 7 9 1 0 4 13 2
9 7 2 9 9 1 13 16 4 2
11 9 9 1 9 1 3 13 16 4 4 2
22 9 9 1 9 2 9 1 9 9 1 1 9 9 1 13 4 16 1 3 4 4 2
16 9 9 1 0 9 9 7 9 9 9 1 1 9 1 0 2
11 9 1 9 1 9 12 12 9 14 13 2
17 9 1 9 1 3 13 2 9 12 9 9 1 13 4 4 4 2
29 7 2 9 9 1 9 1 0 4 2 11 5 9 7 11 5 9 9 9 1 4 4 9 9 1 3 0 4 2
28 3 2 12 9 4 1 9 1 9 9 1 9 1 9 1 13 4 4 9 1 9 1 13 4 16 4 4 2
41 9 1 9 1 9 9 9 1 2 9 9 1 0 16 9 9 1 13 16 4 2 1 13 16 2 11 9 1 9 7 9 9 1 9 9 1 13 16 13 4 2
30 12 12 12 12 9 9 1 9 1 13 4 16 4 4 9 1 9 1 0 1 9 9 1 13 4 4 4 16 4 2
31 9 1 1 9 7 9 2 9 2 9 14 9 1 9 1 0 4 16 2 9 9 1 9 1 9 1 13 4 4 4 2
37 3 9 9 1 13 0 4 9 4 4 9 9 9 9 7 9 9 9 1 9 2 9 9 9 1 9 9 12 9 2 12 9 9 1 13 4 2
23 7 9 9 9 1 9 9 9 9 1 9 12 9 9 1 13 0 9 1 13 4 4 2
32 15 1 2 13 4 4 4 9 1 13 16 13 16 4 4 4 2 1 13 9 9 1 9 9 4 13 4 9 1 13 4 2
23 10 9 1 13 16 9 1 13 16 4 4 9 9 1 9 1 13 9 1 13 4 4 2
12 7 9 1 9 1 13 9 1 13 4 4 2
22 9 1 9 9 1 9 1 9 12 12 9 2 9 1 9 12 9 1 13 16 4 2
24 9 1 9 1 9 1 13 9 1 13 16 2 9 1 3 9 13 16 13 4 4 16 4 2
27 9 1 9 1 9 1 9 1 9 1 13 4 4 9 4 2 9 9 9 1 9 1 13 9 1 13 2
28 7 1 9 1 9 9 1 13 16 1 2 11 9 1 9 1 9 1 9 1 13 16 4 4 1 13 4 2
25 15 1 3 9 1 9 9 4 4 9 9 1 13 16 13 4 4 4 11 9 1 13 4 4 2
33 12 9 5 12 12 9 1 13 4 9 9 1 9 1 0 2 9 9 9 1 9 1 13 16 4 16 1 9 1 9 4 4 2
32 9 9 1 1 13 4 9 1 10 9 1 2 9 9 2 1 13 1 13 16 4 16 2 3 1 0 4 9 4 16 4 2
27 13 4 16 4 16 2 9 9 1 13 14 14 2 9 9 1 4 4 0 9 9 1 13 9 14 13 2
7 7 3 13 16 4 14 2
9 0 16 2 9 1 9 1 0 2
30 9 9 1 15 14 13 14 1 9 9 1 9 1 9 4 4 2 9 1 9 1 9 1 13 2 1 1 13 4 2
26 9 9 1 9 9 4 1 9 1 9 9 4 4 2 11 14 1 9 1 13 4 9 4 1 4 2
8 9 1 3 0 16 4 4 2
14 7 2 0 9 1 13 16 4 9 1 1 13 4 2
13 13 4 9 1 9 1 0 4 13 9 1 13 2
13 10 9 2 0 4 9 1 9 1 13 9 4 2
17 9 7 9 1 13 16 3 4 9 1 13 16 1 9 1 0 2
33 9 9 1 9 1 13 16 1 9 9 1 3 13 4 2 9 9 1 13 9 9 14 9 9 1 13 4 4 4 4 1 13 2
37 15 9 1 9 9 1 12 12 9 9 1 13 9 1 9 1 13 2 9 9 1 13 9 1 13 4 16 4 4 16 2 3 1 13 4 4 2
39 9 1 1 9 1 9 1 13 16 2 12 12 9 9 1 9 9 9 1 9 2 9 9 1 12 9 14 1 13 2 9 9 1 13 4 13 4 4 2
21 9 9 1 1 9 1 9 1 9 1 9 9 1 9 1 13 4 4 4 4 2
11 9 1 9 1 13 9 1 13 4 4 2
18 9 1 13 16 13 14 9 1 0 13 9 1 3 13 4 16 4 2
28 9 1 9 1 9 9 1 9 1 13 14 9 9 1 13 2 11 9 1 9 9 1 3 9 1 13 4 2
24 10 4 4 9 9 1 3 9 9 13 4 16 2 9 9 9 1 9 0 4 9 1 13 2
22 9 9 9 9 9 1 9 1 9 9 1 9 9 1 9 9 13 4 4 16 4 2
17 9 9 1 9 1 9 1 13 4 4 9 1 1 9 4 4 2
20 9 9 1 9 1 9 1 13 9 1 9 13 16 1 3 9 9 4 0 2
48 10 9 9 1 1 3 9 14 1 13 4 9 7 9 9 9 14 9 1 9 9 9 1 13 2 9 1 9 1 9 9 13 2 9 1 13 9 1 9 1 13 1 13 9 1 13 4 2
25 15 14 1 0 9 9 1 9 1 13 9 1 9 2 9 1 9 9 9 1 13 16 4 4 2
27 15 1 1 9 1 0 13 16 1 13 9 9 7 2 9 1 12 9 9 1 13 9 9 9 1 13 2
16 15 1 9 1 13 4 4 16 9 9 1 13 9 1 0 2
18 9 1 9 1 13 16 0 9 1 2 9 9 4 1 9 1 13 2
12 9 9 1 9 9 9 1 9 9 1 13 2
36 9 9 9 1 13 4 4 9 1 2 9 1 13 4 16 9 1 0 16 9 1 13 16 1 0 4 16 4 2 1 9 1 13 16 4 2
32 9 9 1 9 1 2 9 13 9 1 13 4 1 13 9 1 13 16 4 2 9 1 13 16 9 1 9 1 9 1 0 2
7 9 1 1 13 4 4 2
10 7 9 9 1 0 4 9 1 13 2
8 9 1 9 9 1 9 4 2
50 9 1 12 5 12 9 1 13 4 4 9 1 12 2 12 9 1 9 1 13 16 9 1 13 4 2 9 4 9 1 9 1 9 1 13 16 2 9 1 13 7 4 4 14 1 13 9 1 13 2
52 9 1 1 9 9 1 9 9 9 1 9 12 9 13 2 9 9 1 1 9 9 1 13 4 4 1 9 9 1 13 4 16 2 9 1 13 4 16 1 9 0 4 1 13 9 1 1 13 16 4 4 2
15 9 4 16 13 4 16 4 1 13 9 1 1 13 4 2
40 9 1 9 1 13 9 1 9 9 4 13 4 9 1 9 1 9 1 13 16 2 9 9 9 1 13 9 1 9 7 9 1 13 1 13 4 9 1 0 2
30 7 9 9 1 9 1 13 9 9 1 13 9 9 9 1 0 2 9 7 9 1 9 1 1 9 1 9 1 13 2
18 9 1 9 14 1 13 9 1 1 9 1 9 1 9 1 13 0 2
44 0 4 9 1 13 9 1 9 9 1 9 9 9 1 9 1 13 9 1 13 9 1 13 16 11 9 9 9 1 13 16 4 2 9 9 1 9 4 1 13 9 1 13 2
33 7 2 9 9 1 10 9 13 4 9 2 9 1 3 13 0 9 1 13 2 9 1 9 1 9 13 4 16 4 9 1 13 2
36 9 9 9 1 12 9 9 9 1 13 16 13 4 4 16 2 9 1 9 7 9 9 1 9 14 1 9 1 0 4 4 1 1 13 4 2
32 9 9 1 1 9 9 4 9 1 13 4 9 1 9 9 1 13 16 1 13 4 4 9 9 1 13 16 4 9 9 4 2
25 9 7 9 9 9 14 1 9 9 1 9 1 13 9 1 13 16 1 4 16 4 1 4 14 2
14 9 9 1 13 16 1 9 1 9 1 3 13 4 2
24 9 9 9 1 13 1 1 0 9 1 2 12 9 1 9 14 1 13 9 1 1 13 4 2
14 9 1 9 1 9 9 1 1 9 1 13 16 4 2
16 2 9 9 2 1 9 13 12 9 1 9 1 9 1 13 2
35 9 2 9 9 1 13 4 4 0 9 9 9 1 2 9 1 1 9 1 2 9 3 2 2 9 9 2 1 13 9 1 13 16 4 2
31 9 1 9 1 13 4 16 3 9 1 9 1 13 2 9 1 13 4 14 2 9 9 9 2 1 13 4 4 16 4 2
89 7 2 9 9 1 15 14 9 7 9 14 1 0 4 9 1 13 4 16 4 4 9 1 9 9 4 13 16 2 3 0 1 9 2 3 13 4 9 9 1 13 4 16 4 4 1 13 9 4 2 1 9 1 13 2 12 12 12 9 1 13 4 9 1 13 16 2 9 9 1 9 1 1 9 1 9 9 4 13 2 14 9 1 9 1 13 16 4 2
35 9 9 13 16 2 12 12 9 9 13 9 1 3 1 13 2 11 1 9 9 9 1 9 1 13 16 4 1 2 1 13 14 4 4 2
24 10 9 1 9 7 12 9 13 4 4 4 9 9 1 9 9 1 14 9 1 13 9 14 2
24 9 9 1 9 9 1 1 4 1 13 9 1 13 4 16 1 9 1 13 4 9 9 4 2
20 0 9 1 9 1 1 13 4 4 2 1 13 16 1 9 1 1 4 4 2
69 2 9 9 1 1 9 9 9 9 1 9 9 1 9 2 2 9 9 1 9 9 1 9 9 1 1 9 2 2 9 1 9 9 9 1 9 2 2 9 9 1 9 9 1 9 2 14 9 1 13 4 16 4 4 9 1 9 1 2 9 9 2 1 3 13 4 16 4 2
34 7 2 9 1 13 9 1 9 2 2 9 9 9 9 9 1 13 9 9 2 14 1 9 1 2 9 9 2 1 13 4 4 4 2
30 9 9 4 13 4 2 9 9 2 1 12 12 9 1 13 4 16 2 9 1 3 9 9 14 1 9 9 1 9 2
28 0 13 4 4 9 1 9 1 13 16 1 2 11 9 9 7 9 1 9 9 1 13 9 9 9 4 4 2
32 7 13 4 4 16 4 4 9 1 9 9 1 9 9 9 1 9 1 13 4 14 4 2 9 9 1 9 1 13 16 4 2
21 7 9 9 1 9 1 13 9 1 9 9 1 13 16 13 4 4 16 4 4 2
20 9 9 1 9 1 13 4 9 1 9 9 1 9 1 13 9 1 13 4 2
41 15 1 9 9 1 2 9 9 2 2 9 9 2 2 9 9 2 1 12 9 13 4 9 1 13 9 1 9 4 9 9 1 13 16 4 9 1 0 16 4 2
30 9 1 1 9 9 1 13 9 9 1 9 1 13 4 4 16 4 9 9 1 13 16 2 9 9 1 0 4 13 2
29 9 1 9 9 13 16 9 1 13 2 9 1 9 9 1 13 4 9 1 13 2 9 9 4 9 1 3 13 2
10 15 1 13 4 9 4 16 4 4 2
16 10 9 7 9 1 9 1 13 16 1 9 9 14 13 4 2
28 9 1 9 9 4 4 15 9 1 9 1 13 2 9 9 1 13 14 9 1 13 4 9 4 16 4 4 2
47 9 9 1 12 12 9 2 9 9 1 9 9 9 1 13 2 9 1 13 4 9 1 0 4 9 1 13 2 9 1 2 9 9 12 9 9 2 1 13 16 9 9 13 9 1 13 2
30 11 9 1 9 9 7 0 9 1 9 1 9 9 1 9 1 9 2 9 1 9 1 13 2 1 13 4 16 4 2
19 13 4 4 9 1 0 4 16 9 1 9 1 9 1 13 4 16 4 2
37 2 12 12 9 1 9 2 12 12 12 9 1 9 2 12 12 9 1 9 1 13 4 16 9 1 13 16 4 2 9 1 9 1 13 16 4 2
44 2 12 12 12 9 1 9 1 13 4 16 4 16 2 9 1 12 12 12 9 2 15 1 12 12 12 9 1 3 9 9 2 15 1 13 16 1 0 4 1 4 9 4 2
29 11 9 9 9 9 9 1 2 9 9 7 9 9 1 13 4 9 9 9 1 2 0 9 1 9 1 13 4 2
24 9 12 12 12 9 1 9 1 2 3 9 9 1 13 16 2 9 1 0 9 2 1 13 2
25 9 9 1 9 2 0 9 9 9 14 1 9 2 9 1 9 1 13 4 16 12 12 12 9 2
18 9 9 1 13 16 1 9 9 1 12 9 7 9 1 12 9 4 2
21 10 9 1 9 7 9 9 1 13 9 1 13 9 1 15 14 13 4 4 14 2
26 9 1 12 12 12 9 13 9 0 13 2 7 9 1 13 16 1 4 4 0 4 9 9 4 4 2
20 10 9 9 7 9 9 1 13 14 2 9 1 15 1 13 2 3 13 14 2
12 9 9 4 9 1 13 4 16 4 16 4 2
12 9 1 9 9 9 1 2 10 9 1 13 2
50 2 9 1 13 4 16 1 11 9 2 2 9 9 4 4 15 9 1 9 4 16 2 9 9 1 13 4 16 13 4 2 9 1 13 16 1 9 1 13 2 9 1 9 1 13 16 4 4 16 2
71 2 9 1 9 12 9 1 9 12 9 1 1 3 13 4 2 2 9 9 1 9 1 13 16 1 9 9 7 9 9 1 13 4 2 2 9 9 1 3 9 12 9 1 13 16 4 2 2 12 9 9 7 12 9 9 1 0 1 9 1 13 2 9 9 1 12 12 9 1 0 2
76 2 9 9 1 9 9 1 9 9 1 0 2 2 9 1 9 1 12 9 2 9 1 13 2 15 1 9 1 13 2 9 9 9 1 13 9 1 13 16 1 9 0 2 2 9 1 13 4 9 1 9 1 9 1 0 4 16 2 9 1 0 2 3 0 4 9 1 9 4 9 1 0 2 5 5 2
5 13 9 9 4 2
30 9 9 1 9 1 2 3 2 9 1 9 2 1 13 2 10 9 1 9 1 9 9 1 3 0 4 9 4 4 2
44 9 1 9 14 9 1 9 1 12 9 13 2 9 9 1 13 4 0 13 9 9 1 2 9 9 1 13 4 4 9 4 2 13 4 16 12 9 9 1 1 13 4 4 2
71 9 9 1 9 1 9 1 9 9 4 13 4 16 4 9 14 1 2 0 4 9 1 13 16 2 9 9 1 9 7 9 1 11 9 1 9 9 9 9 1 13 4 2 9 9 1 9 9 4 13 1 13 9 9 1 9 1 9 12 12 12 12 12 12 12 9 1 13 16 4 2
34 9 1 2 12 9 1 13 9 9 9 1 9 12 9 1 0 13 4 4 16 9 9 9 1 13 4 4 9 13 4 16 4 4 2
66 9 1 9 2 15 14 1 0 9 9 4 9 1 13 16 4 9 1 1 2 12 12 12 12 9 9 1 9 12 9 9 1 9 9 9 1 13 9 9 4 9 7 2 9 9 1 9 9 1 9 9 1 13 4 16 4 9 2 7 9 9 1 9 1 13 2
49 7 2 9 1 9 9 1 13 4 9 9 7 9 9 1 3 9 1 9 1 14 4 2 9 9 1 13 16 13 4 4 9 9 9 1 9 9 1 13 16 13 4 4 16 4 14 4 4 2
44 9 1 1 9 9 1 13 16 1 9 9 1 12 12 12 12 9 1 13 4 4 16 2 9 9 14 1 9 1 12 9 9 1 13 4 4 4 2 0 4 9 1 13 2
35 7 9 9 1 9 9 1 9 1 13 2 9 1 0 9 1 13 4 16 1 13 9 1 13 9 1 13 14 2 1 1 9 1 13 2
49 9 9 1 13 4 9 1 13 1 13 16 2 9 9 1 9 1 1 4 2 3 9 9 1 1 13 4 15 9 9 1 9 1 9 2 9 1 13 9 1 13 4 2 1 13 9 4 4 2
24 9 1 13 4 4 16 1 2 9 7 9 1 9 4 13 4 9 1 13 9 1 1 4 2
49 7 9 9 1 9 9 1 13 9 9 1 13 4 4 7 2 9 1 9 9 1 13 16 13 16 2 9 9 1 9 1 13 16 2 3 1 9 9 1 9 1 1 13 16 4 1 4 14 2
40 9 9 1 0 9 4 9 9 1 3 13 9 1 9 9 1 9 1 13 4 14 2 9 4 9 1 13 12 9 1 9 1 9 9 4 13 9 1 13 2
41 7 2 9 1 13 4 4 9 1 1 3 9 1 13 4 2 9 9 1 3 13 4 16 4 4 4 9 4 9 9 1 13 16 2 9 1 9 1 0 13 2
28 10 9 1 13 9 7 9 9 1 0 4 0 9 1 13 9 9 1 13 4 16 4 4 16 1 4 4 2
10 9 1 13 0 1 9 1 0 4 2
48 3 13 16 4 16 2 9 9 1 1 2 9 7 9 1 13 4 16 4 16 1 9 4 4 9 2 9 1 9 9 1 9 1 9 9 1 9 14 1 13 12 9 1 2 3 0 4 2
20 9 1 9 1 9 1 9 1 13 9 14 1 9 4 9 1 1 4 14 2
28 7 2 9 1 9 1 13 9 2 7 12 9 14 1 9 1 13 4 16 1 9 1 2 10 9 4 4 2
9 9 1 1 2 7 13 4 4 2
17 12 9 1 9 1 13 16 2 9 1 1 9 1 12 9 13 2
40 9 1 13 4 16 9 9 4 13 4 9 2 9 1 1 9 1 9 7 9 14 1 13 4 16 1 2 9 9 4 9 1 13 16 1 2 3 0 4 2
5 0 9 4 4 2
25 0 9 1 9 5 9 9 1 2 9 9 9 1 9 1 13 4 4 16 12 9 1 13 4 2
17 7 9 1 9 2 9 9 14 13 4 4 9 1 3 4 4 2
16 7 2 9 9 9 9 1 1 2 15 1 13 16 4 4 2
20 2 9 1 0 16 1 0 9 2 14 1 2 13 16 4 9 1 1 4 2
27 9 9 1 13 16 2 0 9 1 9 1 2 11 9 1 9 1 13 4 0 9 1 13 4 4 4 2
20 9 1 9 9 1 2 11 9 1 13 9 9 1 9 1 9 1 13 4 2
24 9 1 12 9 1 9 9 1 1 13 1 13 16 2 3 9 1 9 1 13 1 9 4 2
7 3 9 1 0 16 4 2
12 3 2 15 9 1 9 1 13 16 4 4 2
20 12 12 13 9 9 9 1 9 2 9 9 1 9 9 9 1 13 16 4 2
20 9 1 9 1 13 4 16 2 9 1 9 13 9 1 0 4 9 1 13 2
32 0 9 1 9 1 13 16 13 4 4 4 4 2 0 9 1 9 1 13 4 4 9 2 0 4 9 9 13 4 4 4 2
24 7 9 1 0 9 1 2 9 1 9 1 9 1 13 16 2 9 9 1 13 4 4 4 2
28 3 2 9 9 9 14 13 16 2 9 1 9 1 9 1 9 1 13 16 4 9 1 13 16 1 3 4 2
22 9 13 9 1 2 9 9 1 9 1 2 9 9 9 14 3 14 1 13 16 4 2
18 9 1 13 4 9 1 2 2 9 2 7 2 9 2 1 13 4 2
42 3 9 9 4 2 9 1 13 4 4 9 9 1 1 13 4 4 9 2 7 11 1 13 16 1 13 4 4 16 2 9 1 1 9 9 13 4 9 14 1 13 2
27 7 2 9 1 3 4 4 16 1 2 3 9 9 9 1 1 9 0 4 13 16 4 9 1 0 4 2
22 3 15 1 13 4 16 4 16 2 10 9 9 9 1 9 1 9 1 13 4 4 2
23 3 0 9 9 1 9 1 9 1 13 2 9 9 1 9 1 13 9 1 13 16 4 2
11 9 7 9 14 1 15 1 13 4 4 2
33 11 1 12 12 12 12 9 1 2 9 9 2 1 9 1 13 4 4 4 16 2 10 9 1 9 1 3 9 1 13 4 4 2
19 7 3 9 1 0 9 1 14 2 9 1 13 9 1 0 4 4 4 2
27 7 2 9 1 2 9 9 1 9 1 9 1 0 13 4 9 1 1 2 10 9 1 13 4 4 4 2
27 9 9 1 13 14 2 7 9 9 9 9 9 1 13 4 14 9 9 1 13 4 4 4 1 4 14 2
30 10 9 2 2 9 2 1 13 16 1 9 1 9 1 13 9 1 13 4 4 16 4 9 1 0 9 1 1 4 2
24 9 1 9 1 2 9 7 9 9 9 9 1 13 9 9 9 1 1 9 1 13 16 4 2
21 9 1 15 1 13 16 1 10 9 1 9 1 2 9 9 1 13 4 16 4 2
22 7 2 9 1 9 9 1 13 16 2 9 1 9 1 0 16 2 9 1 1 0 2
24 3 9 9 9 1 2 9 2 9 1 13 16 2 9 9 9 1 13 4 16 4 1 13 2
13 3 13 16 2 13 4 4 9 1 3 4 4 2
21 9 7 9 1 2 0 4 9 9 4 9 1 13 9 1 0 4 13 4 4 2
16 9 1 9 1 9 9 1 9 1 13 9 1 13 4 4 2
7 3 1 9 4 4 4 2
17 7 2 15 14 1 9 1 9 1 3 13 4 9 1 1 4 2
25 9 1 13 9 1 3 0 9 1 1 9 1 0 4 2 9 1 1 0 9 1 13 4 4 2
36 9 1 9 9 1 2 9 9 1 13 4 4 11 9 9 1 11 11 9 9 9 1 9 9 1 11 1 1 9 9 1 13 4 1 13 2
17 9 1 1 15 1 13 9 7 9 9 1 13 4 16 4 4 2
5 3 9 4 4 2
29 9 1 9 9 1 2 9 9 1 9 1 13 16 4 4 14 1 2 9 9 1 9 1 1 9 1 13 4 2
15 9 9 1 1 9 1 2 9 1 1 9 1 13 4 2
23 0 9 9 1 9 1 2 9 9 1 9 7 9 1 13 4 9 1 3 0 4 4 2
39 9 9 2 9 9 9 1 0 16 1 9 1 0 16 2 9 9 1 2 0 9 1 9 1 13 4 2 9 9 1 13 9 1 0 13 4 1 13 2
24 7 2 9 9 9 1 13 4 16 9 1 13 4 9 9 1 9 13 9 1 13 16 4 2
16 9 1 9 9 1 1 2 0 9 1 3 13 1 13 4 2
22 7 2 9 9 1 9 14 4 4 2 9 1 1 13 16 4 16 4 1 4 14 2
22 10 9 2 9 1 9 9 7 9 9 2 9 1 13 16 2 9 1 13 4 4 2
22 9 2 9 1 12 9 9 4 4 9 1 9 1 2 9 1 13 4 16 4 4 2
41 9 1 9 1 2 9 9 7 9 1 9 1 13 4 9 1 9 9 1 13 4 16 2 9 9 1 9 1 13 4 16 4 4 1 13 9 1 13 4 4 2
64 7 2 12 12 9 9 1 9 7 9 1 9 1 9 1 2 9 1 9 1 2 15 1 0 9 14 1 13 1 1 2 2 9 1 9 1 13 2 1 13 4 4 2 9 1 13 4 9 9 7 9 9 1 9 1 13 16 4 16 4 1 4 14 2
24 7 2 9 1 9 9 4 4 2 10 9 2 9 9 1 0 4 4 9 1 13 16 4 2
29 7 9 7 9 1 13 9 1 2 9 9 1 9 1 13 1 13 13 4 9 1 9 9 1 13 16 4 4 2
42 3 13 16 2 15 1 13 16 4 16 14 2 0 16 14 1 9 1 0 2 9 1 13 2 9 1 9 1 13 0 9 14 1 13 4 16 4 4 16 4 4 2
47 0 9 9 1 2 9 14 13 4 16 4 9 1 1 4 16 4 16 2 9 1 9 1 9 14 13 16 4 4 4 14 2 15 1 1 13 9 1 9 1 3 13 9 2 1 13 2
20 0 4 2 9 9 1 2 9 9 1 0 4 4 16 2 9 1 3 13 2
27 9 2 9 1 13 1 2 9 2 9 9 1 9 9 1 13 16 2 9 1 13 9 16 13 9 4 2
26 11 9 9 9 1 4 4 2 9 9 1 13 2 9 9 1 13 4 4 13 4 9 1 3 13 2
27 9 2 9 1 13 4 16 1 2 9 1 12 2 12 9 1 13 9 14 1 2 9 1 13 4 4 2
26 9 2 9 2 9 2 9 2 9 9 1 9 14 9 1 9 1 13 16 4 9 1 9 1 0 2
33 9 1 9 2 9 9 1 9 9 4 13 2 0 4 13 4 16 2 9 1 9 1 13 16 9 1 13 4 4 9 1 13 2
17 9 9 4 1 9 1 9 1 1 13 16 2 9 1 3 0 2
17 2 9 1 9 1 13 9 1 0 9 1 13 0 9 1 13 2
63 11 11 9 1 11 1 13 4 4 11 1 11 11 9 1 2 9 12 12 9 1 13 9 1 13 2 9 1 9 1 13 4 9 5 9 1 9 1 9 1 13 4 1 13 9 1 1 2 9 9 2 9 1 13 16 2 10 9 1 13 4 4 2
56 11 9 1 2 10 9 1 13 4 4 16 1 3 1 9 4 16 2 10 9 1 2 3 11 1 9 9 1 9 1 13 7 13 16 2 9 9 9 14 4 4 11 9 1 9 1 13 4 4 9 1 13 4 16 4 2
43 9 2 9 1 9 1 12 9 1 0 2 9 1 9 1 13 4 4 4 9 1 13 2 11 9 1 9 1 13 2 9 1 13 4 1 13 9 1 13 16 4 4 2
42 9 9 9 1 13 16 1 2 11 9 1 11 11 9 2 11 9 1 1 11 9 9 9 1 9 9 1 1 4 4 1 13 9 1 9 1 13 16 13 4 4 2
37 9 1 9 1 9 4 13 4 2 15 1 3 9 1 13 4 9 1 13 16 4 4 14 1 2 9 1 13 16 1 0 2 0 9 4 4 2
26 9 9 4 4 4 16 1 3 2 9 9 4 1 4 4 9 1 13 4 16 4 4 16 4 4 2
16 7 13 16 13 4 9 4 4 9 1 7 9 4 4 4 2
72 15 9 1 2 9 1 9 1 13 16 9 9 1 13 16 1 9 9 1 13 4 9 1 9 4 13 4 9 4 4 2 10 9 1 1 9 9 7 9 9 9 1 1 9 5 9 2 9 1 13 4 9 5 9 1 13 14 1 9 1 13 4 9 9 1 9 1 13 16 4 4 2
51 9 9 1 9 9 9 9 1 2 11 11 9 9 1 2 15 9 1 9 1 13 16 9 4 9 1 13 4 4 11 1 9 9 1 1 9 1 9 1 9 3 13 4 16 4 4 2 1 13 4 2
6 0 4 9 4 4 2
47 2 9 9 2 1 2 11 1 11 1 9 1 13 16 9 1 9 9 1 9 1 13 4 9 1 13 4 2 11 9 1 1 9 1 9 1 9 1 13 9 1 13 9 4 1 13 2
59 9 11 1 13 4 4 9 9 9 1 12 9 9 1 9 1 2 9 12 12 9 1 9 1 2 9 1 9 1 13 4 2 9 1 9 1 1 9 1 13 4 9 9 1 9 14 1 9 9 4 13 2 9 1 13 4 16 4 2
33 9 1 11 11 9 7 11 11 9 9 2 11 11 2 9 1 9 2 9 9 9 9 1 9 1 9 9 1 13 4 16 4 2
12 9 1 0 9 7 9 9 1 13 16 4 2
59 7 13 16 2 9 9 1 0 4 4 2 3 1 9 9 1 13 4 4 4 16 2 3 1 9 2 9 9 9 1 9 9 1 9 1 9 9 9 1 13 2 9 1 9 1 13 4 9 14 13 4 16 4 16 1 9 4 4 2
13 11 9 1 2 10 9 1 13 4 4 9 4 2
43 9 1 9 9 1 9 1 13 4 4 1 13 16 9 1 9 9 4 16 2 9 9 9 1 9 1 13 16 4 2 9 9 9 9 1 13 4 4 4 9 4 4 2
20 9 1 1 2 3 13 4 16 9 9 9 1 1 1 9 1 13 16 4 2
49 11 2 9 9 9 9 2 13 4 4 1 13 16 9 1 9 1 13 4 4 16 13 4 16 4 16 4 4 16 2 10 9 1 13 4 9 1 13 4 4 16 4 1 4 14 1 13 4 2
15 10 9 2 11 1 13 9 1 9 1 13 16 4 4 2
27 9 9 9 1 1 9 9 1 13 2 9 3 0 9 7 9 2 9 9 1 13 16 4 9 4 4 2
33 2 9 1 13 2 9 1 9 1 13 4 2 1 1 11 11 9 9 5 9 1 9 1 9 9 1 13 16 13 4 4 4 2
27 9 1 12 12 9 13 4 4 9 9 12 12 9 1 9 9 9 9 9 9 9 1 1 9 4 4 2
15 15 9 1 9 1 9 1 2 10 9 1 13 1 13 2
11 9 1 2 9 2 1 13 9 4 4 2
36 10 9 1 1 11 9 9 12 12 9 2 9 9 9 12 12 9 1 13 4 2 13 16 12 12 12 12 9 1 13 9 9 1 13 4 2
13 9 1 9 1 2 11 9 1 3 13 4 4 2
14 10 9 1 13 4 9 1 13 1 1 2 3 0 2
12 9 9 1 9 9 1 9 9 4 9 4 2
9 9 1 13 16 12 12 9 9 2
29 9 9 1 2 9 4 9 2 2 13 4 9 2 7 2 9 1 13 2 1 13 4 9 4 9 1 13 14 2
30 9 1 1 9 1 13 4 4 9 1 13 1 13 4 4 16 2 10 9 1 9 1 3 1 13 16 4 4 4 2
36 9 12 12 9 1 9 1 13 16 2 9 9 1 9 1 13 9 1 3 13 16 14 2 9 1 3 9 1 13 16 4 9 1 13 4 2
17 9 9 1 9 9 9 1 13 16 4 4 16 1 10 12 9 2
40 9 1 9 1 11 1 1 9 9 1 2 12 12 12 2 1 13 4 14 4 2 10 9 1 9 9 1 13 4 4 1 13 9 1 13 16 4 9 4 2
23 9 1 13 4 16 1 2 9 9 1 9 4 13 16 1 2 9 0 16 14 13 4 2
35 9 1 9 1 9 9 4 4 4 9 14 1 13 4 2 9 9 4 4 4 9 1 13 4 1 13 16 4 2 1 3 13 4 4 2
23 9 9 1 1 9 9 1 13 11 9 1 9 1 1 2 9 9 1 9 1 13 4 2
40 9 1 10 9 11 1 2 11 9 1 1 2 9 9 2 9 1 13 4 2 9 7 9 1 13 4 11 1 9 1 9 9 13 2 1 13 4 1 13 2
39 10 9 1 9 1 0 4 4 16 2 11 1 3 9 1 13 16 4 4 1 1 9 1 2 11 1 13 4 9 1 9 1 13 16 4 1 4 14 2
24 2 9 4 2 13 4 2 1 13 4 16 13 14 2 1 1 9 1 9 1 0 14 13 2
26 10 9 1 13 4 16 3 9 1 13 4 16 1 2 9 1 13 4 4 9 1 13 4 4 4 2
27 7 2 9 1 9 1 13 9 1 0 1 13 4 4 10 9 1 2 9 1 3 0 4 4 4 14 2
11 9 1 9 1 3 0 4 4 4 14 2
26 10 9 14 9 1 13 4 16 2 3 9 9 1 3 1 13 2 10 9 1 13 4 16 4 4 2
16 10 9 1 7 2 9 9 1 13 9 1 1 4 16 4 2
34 2 11 1 1 9 1 13 4 2 7 2 11 14 1 1 9 1 2 3 9 9 9 9 1 9 4 4 2 1 1 9 1 13 2
24 12 12 9 9 9 1 9 1 13 2 9 7 13 4 16 9 1 9 1 13 4 16 4 2
15 7 2 11 9 1 0 16 9 1 0 4 9 4 4 2
21 9 1 13 4 4 9 9 1 13 16 2 9 14 1 9 4 1 4 4 4 2
23 15 1 9 1 0 9 1 13 16 2 9 12 12 9 1 13 9 1 13 9 1 13 2
44 10 9 1 9 1 13 4 16 4 1 4 2 0 4 2 9 9 4 9 1 13 4 1 13 16 2 3 9 1 9 7 9 7 2 7 9 1 13 9 1 13 4 4 2
16 9 1 13 16 1 2 9 1 14 13 9 1 13 4 4 2
11 9 1 1 9 1 13 9 1 13 4 2
18 9 9 9 9 1 9 9 1 2 9 5 9 1 9 1 13 4 2
22 9 7 9 9 9 9 1 2 12 9 9 1 9 1 13 4 1 13 16 4 4 2
31 0 9 1 9 1 9 1 13 16 2 0 9 1 13 16 13 4 9 9 4 9 1 1 13 4 4 4 9 4 4 2
31 9 9 4 4 11 11 9 7 11 11 9 9 1 2 9 1 2 9 9 1 9 13 2 1 10 9 1 13 16 4 2
11 9 1 13 16 1 3 0 1 4 14 2
28 7 9 1 9 1 13 16 0 9 1 9 1 13 4 4 16 1 2 9 9 1 1 4 11 9 4 4 2
32 9 9 1 12 9 1 13 9 1 13 4 4 9 2 9 1 13 4 9 1 2 9 1 13 4 1 13 9 4 4 4 2
28 3 0 9 1 9 14 4 2 9 1 9 1 13 16 1 0 4 1 13 9 1 2 9 1 13 16 4 2
24 13 16 4 16 2 10 9 1 3 1 13 9 1 13 16 13 4 16 4 4 16 4 4 2
10 9 1 13 4 16 1 9 9 0 2
23 3 9 9 9 1 0 1 0 4 4 2 9 1 13 9 1 9 1 0 9 4 4 2
27 13 4 4 4 4 0 4 2 9 9 1 9 13 2 13 2 9 9 1 9 9 13 4 14 13 4 2
20 7 2 10 9 1 9 1 2 0 4 13 14 1 9 1 1 4 16 4 2
10 15 1 13 16 2 9 1 3 13 2
20 3 2 9 9 1 13 4 9 9 9 9 1 2 9 1 9 1 13 4 2
43 7 2 9 9 7 9 1 9 1 13 16 2 9 9 1 9 9 1 13 4 4 2 1 1 9 1 9 9 4 13 4 9 2 12 12 12 12 9 1 13 4 4 2
6 3 1 9 4 4 2
17 9 1 9 1 9 1 13 16 1 2 14 9 2 4 16 4 2
13 15 1 13 1 9 1 3 9 1 13 4 4 2
33 11 9 1 13 16 2 9 7 9 9 1 9 9 1 0 9 1 13 16 2 13 4 4 9 9 9 1 13 4 2 4 4 2
42 7 2 9 5 9 1 9 9 1 1 3 2 12 9 9 1 9 14 1 2 9 9 9 9 14 1 9 9 2 9 9 1 9 1 13 4 13 2 1 13 4 2
28 2 9 1 9 9 2 1 9 1 2 9 9 4 9 1 13 1 13 9 7 9 1 15 14 1 9 14 2
25 9 5 9 1 9 9 1 2 10 9 7 13 4 9 1 3 13 16 4 16 1 3 4 4 2
19 10 9 1 13 16 2 13 9 1 3 0 14 2 1 3 13 4 4 2
15 15 1 9 1 13 4 2 0 9 9 13 9 1 0 2
6 9 4 9 1 13 2
33 9 2 9 5 9 1 9 1 13 16 4 4 9 7 2 9 9 9 2 9 9 9 14 1 2 3 9 1 13 16 4 4 2
21 10 9 1 2 9 9 9 9 1 9 2 9 1 9 9 14 13 16 4 4 2
30 11 14 1 9 9 1 9 9 1 0 9 1 15 1 0 16 9 1 13 4 4 2 1 13 9 1 13 16 4 2
12 9 4 1 13 4 0 9 4 1 4 14 2
28 9 1 13 0 9 1 13 9 1 1 2 0 9 1 9 1 13 4 16 13 4 4 11 9 1 13 4 2
22 10 9 2 9 9 1 9 1 13 4 9 9 1 9 9 1 13 9 1 0 4 2
15 9 9 1 13 9 1 9 9 1 13 4 16 4 4 2
21 9 1 9 1 2 9 9 1 13 9 1 9 1 9 1 12 9 1 13 4 2
29 9 1 2 9 1 9 1 13 9 1 13 4 2 1 13 2 9 1 13 9 9 1 9 9 1 13 4 4 2
33 10 9 2 9 1 13 4 16 2 9 1 2 13 4 14 13 2 2 9 1 2 9 1 13 16 1 9 2 1 3 13 4 2
17 11 9 5 11 9 9 1 1 2 9 9 9 1 13 4 4 2
30 12 9 1 0 9 1 13 4 2 9 7 9 1 13 4 9 1 9 9 1 13 16 9 9 1 9 1 13 4 2
19 2 9 7 9 2 1 13 4 4 4 9 9 9 9 1 9 4 4 2
37 9 12 9 1 9 9 1 9 9 1 13 16 2 9 9 2 9 9 2 9 1 13 4 16 9 1 13 4 9 9 1 13 4 2 1 13 2
26 9 1 9 1 13 4 4 9 1 13 9 9 9 1 9 1 13 4 9 9 1 9 1 13 4 2
9 9 1 9 1 9 9 13 4 2
10 10 9 1 13 4 0 9 1 13 2
36 2 9 9 1 9 1 13 4 4 9 1 9 1 13 16 4 4 2 2 9 1 9 9 1 13 9 1 9 1 13 16 4 2 5 5 2
13 10 3 1 13 9 1 2 3 13 4 16 4 2
16 9 9 1 9 1 2 9 9 5 9 1 13 4 9 4 2
64 9 12 12 12 12 9 1 9 9 1 9 9 9 9 2 9 5 9 9 2 9 9 1 12 9 9 1 13 9 1 2 9 1 13 16 1 9 1 9 1 1 4 16 2 12 9 9 0 2 3 9 9 1 13 9 1 13 16 1 4 4 9 4 2
22 9 9 1 13 12 12 9 1 11 9 9 1 2 7 2 10 0 9 1 13 4 2
39 9 1 9 1 2 9 12 9 1 9 9 9 1 9 9 1 13 16 4 4 16 2 9 9 1 2 9 2 1 13 2 9 9 9 1 13 4 4 2
15 9 12 9 1 2 0 4 9 2 1 9 1 13 4 2
32 9 1 2 9 1 9 1 2 9 1 13 2 1 2 3 13 4 4 16 2 9 9 9 1 9 1 9 9 1 13 4 2
80 9 1 13 9 1 9 9 9 14 1 9 1 13 4 16 2 2 9 9 9 1 12 12 9 9 1 13 2 9 1 9 9 9 1 13 4 4 9 1 12 9 9 13 4 2 2 9 9 9 1 9 1 9 9 1 13 4 16 4 16 2 9 1 1 9 9 4 3 0 4 9 1 13 2 1 13 4 16 4 2
11 9 1 9 1 0 4 4 16 4 4 2
17 3 2 10 9 7 9 1 13 2 13 9 4 4 16 4 4 2
25 9 1 9 1 13 4 7 2 9 1 13 9 1 2 9 1 9 9 1 9 7 9 1 13 2
66 12 12 12 12 9 9 1 1 2 9 1 13 16 9 9 9 1 13 2 13 4 4 9 4 9 1 9 9 9 1 13 16 2 11 9 1 2 9 4 9 7 9 1 13 14 1 9 4 4 9 2 9 9 9 1 1 9 1 13 4 2 1 13 4 4 2
20 10 0 4 9 1 13 4 2 13 4 16 1 9 1 9 4 4 9 4 2
39 9 1 13 4 9 12 9 1 9 9 1 13 9 1 2 9 1 13 4 4 9 7 9 1 9 9 7 1 1 2 9 7 9 14 1 13 4 4 2
23 11 9 2 9 1 12 9 9 1 13 9 1 2 9 9 4 9 1 9 1 13 4 2
37 9 12 1 2 9 2 11 9 9 1 9 1 13 9 9 1 9 9 4 4 2 9 12 1 9 9 1 9 9 2 7 9 1 9 4 4 2
25 12 12 9 1 9 9 9 9 1 9 9 9 1 2 3 9 1 9 1 9 1 13 16 4 2
36 7 2 13 16 4 4 16 1 2 0 4 9 9 1 9 9 1 9 2 13 4 4 2 0 4 4 13 4 4 14 2 1 13 9 4 2
39 9 9 1 9 1 11 11 9 1 2 9 5 9 5 9 5 9 2 1 13 9 9 1 13 16 2 2 0 4 9 1 13 4 2 1 13 4 4 2
34 9 1 13 9 1 1 4 16 2 9 1 9 9 1 9 1 9 7 9 1 3 13 16 4 14 2 13 16 4 16 4 4 14 2
41 9 9 1 9 1 2 9 9 1 1 9 1 13 16 13 4 1 13 9 1 9 1 13 2 9 7 9 2 9 1 13 16 13 4 1 13 9 1 13 4 2
14 10 9 1 9 1 9 2 9 1 13 4 16 4 2
16 2 9 1 13 4 4 2 1 1 9 1 13 4 16 4 2
25 11 1 9 5 9 5 9 1 9 9 1 9 9 1 13 4 16 4 2 10 9 1 3 0 2
31 9 9 1 13 16 1 2 9 1 9 14 1 13 16 4 4 1 1 9 1 2 10 9 1 0 13 9 4 1 4 2
17 10 9 1 13 4 9 1 2 9 1 13 9 1 13 4 4 2
14 9 9 1 2 9 1 13 9 1 13 4 16 4 2
56 9 9 1 9 1 9 1 2 9 9 1 9 9 1 9 1 13 4 16 2 10 9 1 9 9 2 9 9 1 13 9 9 4 9 1 13 1 2 9 7 9 9 9 7 1 9 1 9 9 1 9 1 13 4 4 2
20 7 2 9 9 1 9 1 9 1 2 9 1 0 4 9 1 13 16 4 2
32 9 1 9 9 4 9 9 1 9 1 13 16 2 9 1 13 2 9 1 9 1 2 9 9 1 9 1 13 4 16 4 2
6 15 1 9 1 0 2
23 9 9 1 9 1 9 1 2 9 7 9 1 9 1 13 9 1 13 16 4 16 4 2
22 0 9 1 2 12 12 12 12 9 1 1 11 9 9 1 9 1 1 13 4 4 2
25 9 1 11 9 7 11 9 7 1 9 1 2 9 7 9 1 13 4 4 16 4 4 16 4 2
19 7 2 9 0 4 16 1 2 9 9 9 1 1 9 1 9 4 4 2
22 9 9 1 9 7 13 14 1 1 2 9 9 1 13 4 4 9 1 13 4 4 2
42 10 9 1 1 2 3 9 1 13 2 9 0 4 2 9 1 13 9 9 1 2 9 1 13 4 2 15 1 9 9 1 9 9 1 9 1 9 1 13 9 4 2
14 13 4 16 2 9 1 13 4 1 1 15 14 4 2
24 9 13 9 9 9 1 2 9 1 0 2 9 1 9 1 1 13 4 4 14 0 4 4 2
30 9 9 13 4 9 1 9 9 1 3 13 14 1 2 9 1 1 2 9 1 1 2 11 1 9 1 1 13 4 2
20 9 1 9 1 2 15 14 1 15 14 13 16 4 4 4 1 13 16 4 2
14 7 2 3 1 1 9 1 1 15 9 9 1 4 2
25 9 1 9 1 13 16 4 16 2 2 9 9 2 1 0 9 2 13 16 4 4 9 1 0 2
15 9 9 9 1 9 9 1 9 1 13 16 1 4 4 2
6 11 9 1 12 9 2
26 9 1 9 9 13 4 0 4 9 9 1 2 9 7 9 7 1 9 1 9 1 13 16 4 4 2
30 9 9 9 7 9 9 1 9 1 0 9 1 13 4 1 13 9 9 9 1 9 1 13 13 4 9 9 4 4 2
20 0 4 9 9 1 13 4 4 16 2 9 9 1 9 2 1 9 1 13 2
26 9 9 9 1 2 12 12 9 14 1 11 9 7 9 9 1 9 9 9 9 1 13 4 4 4 2
11 12 12 9 1 1 9 1 13 4 4 2
44 11 9 14 12 9 9 9 1 9 1 0 4 4 12 12 9 9 12 12 12 9 1 9 1 2 9 1 9 9 13 16 0 9 7 9 1 13 9 9 4 9 9 4 2
46 9 9 1 13 16 1 2 9 7 9 9 1 9 9 1 13 4 9 4 4 2 9 1 13 16 1 9 1 13 4 2 9 9 1 9 9 14 1 13 4 4 0 9 4 4 2
26 9 1 13 16 9 9 1 9 1 13 16 2 9 1 2 9 9 1 9 9 2 1 13 4 4 2
55 0 4 2 9 9 1 9 9 9 5 9 9 1 12 9 9 1 9 1 9 9 9 2 9 9 9 9 2 9 1 13 0 9 1 2 9 1 13 9 1 13 4 4 9 1 13 1 13 4 16 1 9 1 0 2
26 9 9 1 9 1 13 4 4 2 0 1 13 4 4 9 1 9 9 1 1 9 1 0 4 4 2
21 9 9 1 9 1 13 9 1 13 4 16 2 0 4 13 4 9 1 0 4 2
23 9 9 1 9 1 1 9 1 13 4 9 1 13 16 4 4 1 13 4 1 13 4 2
23 11 9 1 9 9 1 1 2 9 1 13 9 9 7 9 9 1 9 9 1 13 4 2
12 15 1 9 1 9 9 1 9 4 4 14 2
16 2 9 1 13 16 14 2 1 1 9 9 1 13 4 4 2
38 9 9 1 9 1 9 9 7 2 0 9 1 13 16 1 2 9 4 9 1 13 2 9 9 4 9 1 13 9 2 1 2 13 9 1 13 4 2
51 12 9 1 13 9 9 9 1 9 9 9 9 1 13 4 1 1 2 9 9 9 9 1 9 1 13 16 2 9 1 9 1 13 4 1 9 1 13 16 2 3 9 1 13 4 4 2 1 1 13 2
10 9 1 9 1 13 16 9 1 13 2
35 7 2 9 1 9 1 9 2 2 9 1 13 16 2 12 12 9 2 12 9 13 2 14 2 9 9 1 9 1 9 9 1 13 4 2
21 0 4 9 9 1 9 1 13 2 11 9 2 1 1 9 1 13 16 4 4 2
10 9 9 1 13 16 4 9 1 13 2
18 2 9 9 2 1 13 4 4 9 9 1 9 1 9 9 1 13 2
25 9 9 1 9 1 1 2 9 1 9 1 13 13 4 16 4 1 4 14 2 1 9 1 13 2
21 3 9 1 9 1 1 2 9 9 9 1 9 1 13 9 1 9 9 1 13 2
27 9 9 1 2 3 9 1 13 4 14 4 2 9 9 4 9 9 1 3 13 4 2 1 13 16 4 2
28 7 9 1 2 13 4 4 9 1 9 1 13 9 1 13 2 9 9 9 1 9 9 1 13 4 4 4 2
21 9 1 13 9 9 1 2 9 7 9 1 9 1 9 1 13 4 9 1 13 2
15 7 2 15 14 1 9 9 1 13 9 1 13 4 4 2
22 9 9 9 1 9 9 1 13 2 9 9 1 13 9 1 9 9 1 13 4 4 2
8 0 4 13 4 4 13 4 2
17 9 1 2 9 1 13 2 3 3 9 1 13 9 1 13 4 2
8 9 9 1 9 1 0 4 2
31 7 2 9 9 1 9 1 9 13 9 1 13 9 2 9 9 1 9 1 13 4 16 9 1 13 4 4 13 4 4 2
22 11 9 1 9 1 9 1 12 1 13 4 4 9 1 9 9 1 13 16 4 4 2
13 10 9 9 1 13 4 1 1 9 1 13 0 2
42 9 1 12 9 1 12 12 9 1 13 16 4 4 9 9 1 13 16 2 9 1 9 9 1 12 9 1 9 1 12 9 13 16 9 9 1 0 9 1 13 4 2
55 3 9 2 9 9 9 9 1 9 4 13 9 1 12 12 12 9 9 9 1 9 9 9 9 1 12 12 9 9 1 12 12 12 12 12 9 4 2 9 1 12 12 12 12 9 0 2 15 7 9 9 1 13 4 2
20 9 1 9 1 1 9 9 1 1 13 4 2 9 9 9 1 13 16 4 2
11 9 1 3 0 9 1 9 9 1 13 2
20 7 2 9 4 9 1 9 1 0 13 4 4 9 9 1 13 16 4 4 2
25 9 9 4 9 9 1 0 9 1 13 4 16 9 1 13 4 16 4 16 4 16 14 13 4 2
44 7 2 9 7 9 9 1 9 1 13 4 2 9 1 13 16 4 9 1 9 1 13 2 9 9 1 9 1 13 16 4 9 1 9 1 9 1 0 13 4 9 1 13 2
28 9 1 9 2 2 12 12 9 9 2 9 7 9 9 1 13 2 9 9 2 1 9 1 9 1 13 4 2
66 2 12 12 9 9 2 9 1 2 9 1 9 1 9 9 9 4 4 2 9 9 2 1 13 9 1 13 16 2 9 9 1 9 9 9 1 13 4 4 4 9 9 1 9 9 13 4 0 4 9 9 4 16 2 3 9 1 9 1 13 16 1 9 1 13 2
62 9 1 13 16 9 1 9 9 9 1 13 16 0 9 9 1 13 9 9 1 13 4 4 2 2 9 9 2 1 9 1 13 2 9 1 13 4 9 9 2 9 9 1 13 4 16 4 9 14 1 2 9 1 13 4 4 16 13 4 4 4 2
80 7 2 2 12 12 9 9 2 9 1 9 1 13 4 0 1 9 9 1 13 16 2 2 9 9 2 1 1 2 9 9 9 1 9 2 1 13 4 16 4 16 2 9 9 1 13 9 9 4 9 2 0 4 4 9 2 9 1 13 4 16 4 16 14 14 1 3 0 4 2 0 2 9 9 2 1 13 16 4 2
38 15 1 1 2 9 13 16 9 13 4 2 1 2 15 1 9 1 13 4 4 2 2 12 12 9 9 2 9 14 9 4 9 9 1 13 16 4 2
57 2 9 9 2 1 13 4 4 9 9 9 9 9 1 9 1 9 1 9 9 1 9 9 4 9 2 11 11 9 9 9 1 13 4 16 4 2 9 14 1 2 9 9 2 1 13 16 1 9 1 9 1 13 16 4 4 2
53 3 2 9 1 9 9 9 1 13 9 1 2 11 11 9 9 9 9 9 9 1 9 9 4 9 1 9 1 13 16 13 1 13 4 9 9 1 9 1 13 3 9 9 9 1 0 2 9 9 2 4 4 2
37 15 1 13 16 1 2 9 9 1 9 14 4 2 9 9 1 13 16 0 9 1 13 16 4 4 1 13 2 9 2 1 2 9 2 1 0 2
38 11 9 1 11 1 9 9 9 1 13 4 2 9 1 9 1 13 14 4 4 2 9 3 0 9 1 13 4 16 4 4 2 1 9 1 0 13 2
26 9 9 9 1 1 9 1 9 1 9 2 1 1 9 1 9 9 1 14 3 1 13 4 16 4 2
14 9 1 3 13 16 14 2 9 1 3 13 16 14 2
19 15 1 1 9 1 2 10 9 14 13 4 16 4 4 16 4 4 14 2
29 11 1 11 9 1 12 12 9 1 12 9 2 9 1 13 16 11 1 13 2 11 11 9 9 1 13 4 4 2
27 9 9 1 11 5 11 9 1 13 11 9 1 9 1 2 9 1 11 9 1 0 4 9 1 13 4 2
8 11 1 11 1 9 4 4 2
44 12 12 12 12 9 1 9 9 1 13 16 9 12 12 9 2 11 9 1 13 16 3 11 1 1 9 1 13 2 9 1 11 9 1 9 1 13 4 9 1 9 1 0 2
35 10 9 9 1 2 11 1 9 2 1 13 4 1 13 16 11 9 1 9 9 9 1 13 4 4 2 11 1 11 9 1 13 4 4 2
39 7 2 11 9 9 1 13 4 11 9 1 9 1 2 12 12 9 9 1 1 11 9 1 9 1 9 2 12 12 9 1 1 11 9 1 13 4 4 2
16 11 9 1 13 4 16 1 2 12 12 9 1 9 9 4 2
26 11 9 1 9 11 9 1 13 4 16 9 9 1 13 4 9 2 9 9 1 1 9 1 13 4 2
39 9 9 9 1 11 9 1 11 9 9 1 9 1 13 4 2 11 7 11 9 9 1 9 9 9 2 11 5 11 9 9 14 1 9 1 13 4 4 2
24 7 2 9 1 9 1 13 11 7 11 1 9 1 2 11 9 9 1 9 1 13 16 4 2
32 0 9 1 9 1 11 1 2 15 14 0 4 4 9 1 9 1 13 4 2 9 9 1 9 1 13 4 1 13 16 4 2
16 11 9 9 1 9 1 2 10 9 1 9 1 13 16 4 2
21 9 9 1 11 1 9 1 13 2 11 9 9 9 1 10 9 1 13 4 4 2
48 11 1 13 2 11 1 1 9 1 11 1 9 1 9 1 13 4 9 1 9 9 1 13 4 9 1 13 4 16 2 9 3 11 9 1 13 4 9 1 13 4 16 4 9 1 9 4 2
21 10 9 2 9 1 13 16 1 11 1 9 1 1 9 1 13 4 4 4 4 2
44 11 1 9 9 1 9 9 9 1 12 12 9 2 9 9 1 13 4 9 1 13 16 9 1 12 12 9 9 1 13 2 15 1 13 1 9 9 1 9 1 13 4 4 2
22 9 1 9 1 2 11 9 1 9 1 9 9 1 13 4 4 9 1 13 4 4 2
26 9 1 1 9 9 13 4 11 9 9 9 1 1 9 9 9 2 9 9 1 13 16 1 4 4 2
17 11 9 9 9 1 9 1 2 11 1 1 9 9 9 1 13 2
35 11 9 1 1 9 9 4 9 7 9 1 9 1 9 1 13 9 1 9 1 9 1 2 9 9 9 1 13 9 1 13 4 16 4 2
13 11 1 9 1 11 9 1 9 1 13 4 4 2
29 11 9 1 9 1 13 4 9 1 1 2 9 1 9 9 4 9 1 13 16 11 1 9 1 13 4 4 4 2
70 7 2 9 9 9 9 1 9 9 1 9 1 13 16 2 11 9 1 9 1 9 9 1 13 4 13 4 4 16 9 2 11 9 1 2 11 1 9 1 13 4 4 9 2 9 9 1 13 16 4 2 1 13 2 9 1 1 9 9 1 1 13 4 9 1 0 4 13 4 2
39 11 1 9 2 11 12 9 9 9 1 13 16 11 1 9 9 9 1 13 9 1 13 4 14 2 10 9 1 11 9 1 0 9 9 1 13 16 4 2
20 11 1 11 1 13 4 16 2 11 1 9 9 1 13 9 1 13 4 4 2
14 9 1 13 9 1 2 9 1 9 1 1 13 4 2
10 3 9 7 2 9 1 13 16 4 2
16 9 1 9 1 9 1 13 4 9 1 13 16 4 16 4 2
48 9 1 9 2 9 9 9 12 9 1 13 4 9 9 1 13 2 9 9 1 11 1 1 9 1 9 7 9 1 9 1 13 4 4 16 2 9 1 3 9 4 13 16 4 9 1 13 2
37 7 2 9 7 11 1 0 9 1 13 16 1 9 7 9 0 1 2 9 1 1 9 9 1 9 1 3 2 9 1 1 9 1 13 4 4 2
35 10 9 1 1 2 12 12 12 12 9 1 11 11 5 9 9 9 9 1 13 2 9 9 1 2 9 1 13 2 9 1 9 1 0 2
23 9 1 2 9 12 9 1 13 9 9 9 1 9 9 1 13 2 9 1 13 16 4 2
38 9 9 1 2 9 9 9 9 1 9 1 13 4 4 1 13 16 2 3 9 9 9 9 1 2 9 1 9 1 13 4 4 16 4 4 16 14 2
13 9 9 1 0 4 4 2 9 9 1 13 4 2
16 7 11 1 14 2 3 9 9 9 1 9 9 4 16 14 2
25 9 9 9 9 9 1 15 13 4 2 0 4 4 9 1 13 14 1 9 9 1 9 4 4 2
22 9 9 1 2 9 7 9 1 13 9 0 9 9 1 13 4 4 4 1 4 14 2
23 9 9 9 9 9 1 2 11 9 9 1 12 9 9 9 1 13 16 13 4 4 4 2
24 10 9 2 11 1 12 9 9 1 13 4 4 4 2 9 1 13 2 1 13 4 16 4 2
22 9 9 9 1 12 9 9 9 1 13 4 1 13 16 1 2 11 1 9 4 4 2
11 11 1 9 1 13 16 3 4 4 4 2
32 9 1 2 9 9 1 13 4 16 9 9 1 9 1 13 1 1 9 9 1 0 4 11 1 9 9 1 0 9 4 4 2
39 7 2 9 9 1 13 4 16 4 4 9 9 1 9 9 9 9 9 9 1 13 16 2 9 9 9 1 0 9 1 13 9 1 1 9 1 0 4 2
18 0 9 1 2 9 1 9 9 9 1 13 9 1 0 4 4 14 2
37 13 4 4 16 4 9 9 1 1 2 9 9 9 9 1 9 1 13 4 4 16 4 16 2 9 1 13 2 9 9 1 9 1 0 1 13 2
12 9 9 1 9 1 9 9 1 9 4 4 2
9 9 1 13 9 4 1 4 4 2
27 11 9 9 1 2 9 9 1 9 1 9 1 9 1 13 9 1 0 9 1 9 1 13 16 13 4 2
10 7 2 9 1 13 9 1 13 4 2
24 9 1 9 9 9 1 1 2 9 9 7 9 1 1 9 1 13 16 1 4 4 16 14 2
17 7 2 9 9 1 13 9 9 1 9 1 0 16 4 4 14 2
19 9 9 7 9 9 9 1 2 11 1 1 9 1 13 16 1 4 4 2
35 9 9 9 1 13 14 1 9 9 9 1 13 4 16 4 2 9 1 9 9 1 9 1 9 1 13 4 16 1 9 1 1 4 14 2
22 9 9 1 2 9 9 9 9 9 1 9 9 1 0 13 4 1 1 9 1 13 2
8 3 9 4 9 4 4 4 2
26 11 1 2 9 9 9 1 9 1 13 4 9 9 1 1 9 9 9 9 1 9 1 13 16 4 2
35 7 11 9 1 1 2 9 9 1 9 9 9 1 13 4 4 4 16 9 9 9 1 13 4 4 9 1 1 2 9 1 9 1 13 2
12 3 9 9 9 4 4 16 4 4 16 14 2
16 9 7 9 9 2 9 9 1 9 1 0 4 13 16 4 2
12 9 1 9 1 9 1 1 9 1 13 4 2
19 9 5 9 9 1 9 1 13 16 1 9 4 9 1 13 4 16 4 2
20 7 2 9 9 1 9 9 5 9 1 9 1 1 2 3 0 9 1 13 2
7 9 9 1 9 4 4 2
30 9 9 1 12 9 1 9 12 12 9 1 9 9 1 13 4 2 10 12 12 9 1 9 9 1 13 4 16 4 2
22 9 9 1 9 1 13 16 2 9 9 1 9 9 12 9 1 9 9 1 1 4 2
51 7 2 9 9 7 9 9 9 1 9 1 9 9 1 13 2 9 9 1 12 12 9 9 1 9 9 4 4 2 11 1 9 9 9 1 1 4 9 2 9 2 9 2 9 2 9 1 13 16 4 2
19 9 1 9 1 13 16 2 9 1 9 9 1 9 1 13 9 1 13 2
35 2 9 9 1 9 2 1 9 1 9 2 11 1 13 4 4 9 9 1 2 10 9 1 13 9 1 0 4 9 1 13 16 4 4 2
25 3 13 4 4 1 2 9 1 9 1 9 9 1 0 4 9 1 13 16 1 4 4 9 4 2
29 9 1 9 1 9 9 9 1 2 9 9 1 12 12 12 12 9 9 1 12 9 12 9 1 13 4 16 4 2
32 9 11 1 9 1 13 4 9 1 11 7 11 1 1 9 9 1 13 2 11 1 9 1 13 4 9 1 0 13 16 4 2
27 15 1 9 9 4 2 0 4 9 9 1 13 16 4 11 1 2 9 9 9 1 9 1 13 16 4 2
31 12 12 9 9 14 1 9 1 9 9 1 12 12 9 9 4 4 16 1 2 9 1 12 12 9 9 1 13 4 4 2
26 9 9 1 1 12 9 1 13 4 16 2 10 9 1 11 1 9 9 1 13 16 4 4 16 4 2
13 3 9 9 1 9 9 1 9 1 13 16 4 2
30 9 9 1 13 4 4 9 2 9 1 9 9 1 2 9 9 1 13 4 9 1 1 9 1 9 1 13 16 4 2
10 0 9 1 11 1 13 16 1 13 2
38 11 1 9 11 9 1 9 9 7 9 9 1 11 1 0 4 13 4 16 1 2 11 1 9 1 11 1 9 9 1 13 16 4 12 9 4 4 2
16 0 9 1 2 9 9 1 9 9 1 9 9 1 13 4 2
21 9 1 0 9 1 13 4 2 9 9 7 9 9 1 9 1 9 1 0 4 2
32 3 11 1 9 9 7 9 9 9 1 9 1 2 9 9 2 9 2 9 2 9 9 14 9 13 4 9 1 13 16 4 2
15 9 9 1 13 9 9 1 9 1 1 0 9 1 13 2
22 7 2 9 9 1 9 1 13 16 4 4 11 1 9 9 4 9 1 13 4 4 2
24 12 12 9 1 13 4 11 1 1 9 9 1 9 9 1 9 1 2 9 1 9 4 4 2
46 9 1 9 1 9 9 1 0 9 1 13 2 9 9 1 9 9 4 9 1 13 9 4 16 2 9 9 1 1 9 9 2 9 2 9 14 1 9 9 1 13 4 16 4 4 2
20 9 11 1 9 9 9 1 1 9 9 1 9 1 9 9 1 13 16 4 2
26 9 9 1 13 4 9 9 9 1 9 9 1 13 4 9 2 9 9 1 9 7 9 9 1 0 2
16 9 9 1 9 9 1 13 16 2 9 12 1 9 1 0 2
42 9 9 9 1 9 9 9 4 4 11 1 2 9 7 9 9 9 1 13 4 2 11 1 9 9 1 9 9 1 9 12 1 13 9 1 13 4 4 1 4 14 2
37 15 1 13 16 2 11 9 1 1 9 1 13 2 11 5 9 9 1 13 9 9 7 9 9 1 9 9 1 1 9 1 13 16 4 1 13 2
27 15 1 9 14 2 6 2 0 9 1 2 13 1 9 4 4 16 14 2 1 2 13 16 4 4 14 2
18 15 12 9 2 9 1 9 1 13 4 2 1 13 4 16 4 4 2
21 7 2 9 12 12 9 1 9 1 2 3 9 1 13 4 16 4 1 4 14 2
10 9 1 9 1 11 9 1 13 4 2
12 10 9 1 2 0 4 9 9 1 13 4 2
26 15 4 4 16 2 9 14 13 4 4 9 0 9 9 2 9 1 9 9 2 9 1 13 9 9 2
19 3 9 1 12 9 1 13 4 9 13 2 10 9 1 9 9 1 13 2
16 7 2 9 1 9 9 1 9 1 9 1 13 9 1 0 2
15 9 9 1 13 9 9 1 9 1 2 13 4 16 4 2
28 11 1 9 9 9 1 9 1 13 9 9 9 9 2 9 1 9 9 1 13 9 9 9 1 9 9 4 2
13 9 1 9 9 9 1 13 4 1 13 16 4 2
12 9 9 1 9 1 9 9 1 9 1 13 2
14 9 9 1 9 1 13 4 11 1 9 9 1 13 2
17 11 1 9 9 1 9 9 1 12 12 12 12 9 1 13 4 2
37 10 12 12 9 9 1 13 11 9 9 9 9 9 1 2 9 9 12 9 9 1 9 1 9 9 1 12 12 12 9 14 13 4 16 4 4 2
24 9 9 9 9 1 9 1 13 16 1 9 9 1 10 9 1 13 16 9 9 1 13 0 2
26 9 9 1 9 1 9 1 13 4 4 2 9 9 4 4 9 9 9 9 1 13 4 4 9 4 2
14 9 9 1 9 9 1 2 9 9 9 1 3 13 2
18 3 9 9 1 13 9 1 9 1 2 9 9 1 15 1 13 4 2
7 7 9 9 1 9 4 2
23 9 9 9 2 9 9 1 13 9 9 1 2 9 9 1 9 9 13 4 9 1 13 2
26 0 4 9 1 9 1 2 2 9 1 9 1 9 1 1 2 13 9 1 9 9 1 1 9 2 2
7 10 9 14 13 16 4 2
9 11 1 9 9 9 1 3 0 2
6 12 12 12 12 9 2
11 12 9 9 1 12 12 12 12 9 4 2
20 11 1 0 9 9 1 13 4 11 0 9 1 2 9 9 1 13 16 4 2
4 9 9 4 2
10 9 9 1 9 1 13 9 4 9 2
32 15 9 1 13 4 4 9 1 0 9 9 9 2 9 9 2 9 9 1 2 0 13 4 1 13 9 1 13 11 4 4 2
14 9 9 1 0 9 1 13 16 4 16 4 4 14 2
23 11 1 9 9 1 9 1 9 1 13 4 16 1 2 0 9 9 1 0 9 4 4 2
36 0 9 1 15 14 1 9 1 13 4 14 1 13 4 9 9 9 1 1 2 12 9 5 12 12 12 9 9 1 9 1 13 4 16 4 2
9 9 1 9 1 9 1 12 9 2
33 9 9 2 9 2 9 9 1 9 1 2 9 1 9 9 1 0 9 1 1 0 4 2 9 9 1 9 9 0 9 1 13 2
8 9 1 9 9 9 1 0 2
23 7 9 9 1 0 9 1 2 9 9 9 9 1 13 4 2 9 1 13 9 1 13 2
18 0 4 13 9 1 9 9 1 9 9 1 9 9 1 13 16 4 2
20 10 9 1 13 4 9 1 9 1 2 7 9 9 1 13 4 16 4 4 2
17 9 9 1 3 1 0 9 2 9 9 1 9 1 13 4 4 2
23 9 9 1 9 1 9 1 9 1 13 4 9 9 1 2 9 2 9 9 1 13 4 2
18 9 1 13 9 9 1 1 4 9 9 1 13 9 9 1 13 4 2
20 9 12 12 9 2 9 12 1 9 1 9 1 12 12 12 12 9 4 4 2
17 10 9 2 9 9 1 12 12 9 1 13 9 1 13 4 4 2
18 9 9 1 9 9 1 0 4 13 4 2 9 9 1 13 4 4 2
37 7 2 15 1 1 11 9 1 9 1 9 1 13 16 9 9 1 13 4 16 1 2 9 4 4 4 16 2 3 9 9 9 1 9 4 4 2
18 9 7 9 1 13 13 4 16 1 2 11 1 9 12 12 9 9 2
8 11 9 9 9 1 13 4 2
14 9 1 9 1 1 13 12 12 9 9 1 13 4 2
9 11 9 1 9 9 1 13 4 2
12 10 9 1 1 13 4 4 9 4 4 4 2
31 0 9 1 9 2 9 9 9 9 9 9 9 1 9 9 1 13 4 0 4 9 9 2 9 9 9 1 13 4 4 2
18 9 1 9 1 9 9 9 9 1 13 16 4 9 1 1 4 4 2
30 3 2 9 9 1 1 12 12 9 9 2 3 0 2 9 2 16 14 4 9 1 13 4 16 4 1 4 4 14 2
26 2 9 1 13 2 1 13 4 4 9 1 1 2 3 9 9 1 0 9 1 9 9 1 3 13 2
11 7 9 9 1 13 4 9 1 13 4 2
17 3 0 4 9 1 13 4 9 1 9 9 1 13 9 1 13 2
14 9 1 9 1 9 9 1 9 1 13 16 4 4 2
41 9 1 2 9 9 7 9 9 2 9 9 1 13 4 16 4 9 9 1 9 1 2 13 9 1 9 1 13 4 1 13 4 9 9 1 13 4 16 4 4 2
31 9 1 9 9 1 13 4 2 9 9 9 9 9 2 9 1 2 10 9 1 9 1 13 4 16 2 9 1 0 4 2
6 9 1 9 1 9 2
15 9 1 15 14 1 9 9 4 4 16 4 9 1 0 2
17 9 9 9 1 2 9 1 0 16 4 1 13 9 4 1 4 2
43 9 1 3 2 9 9 1 9 1 3 0 4 13 9 1 9 2 7 9 9 7 9 9 1 13 16 1 9 1 13 4 9 9 9 2 9 9 1 9 1 3 13 2
17 10 9 1 13 16 1 0 4 16 1 9 1 9 4 9 4 2
18 15 1 13 4 4 9 1 9 4 4 4 13 4 16 1 4 4 2
13 9 9 1 9 9 9 1 1 10 9 1 13 2
8 9 9 1 13 4 16 14 2
27 9 9 9 1 2 9 2 1 13 4 9 9 1 9 9 9 4 13 2 9 1 9 9 1 13 4 2
8 9 1 0 13 9 4 4 2
11 15 1 10 9 1 10 9 4 9 1 2
10 9 9 1 1 0 4 9 1 13 2
10 12 12 9 9 1 9 9 4 4 2
29 11 9 1 13 9 5 9 2 9 1 9 7 9 9 1 9 9 1 13 2 9 1 9 1 3 1 13 4 2
11 13 4 4 9 1 9 1 13 16 4 2
5 9 1 0 4 2
39 9 1 2 9 9 9 1 9 2 9 1 0 9 1 0 2 1 13 4 2 9 9 9 9 9 9 9 9 2 1 13 4 9 9 1 13 4 4 2
47 9 1 9 12 9 9 9 9 1 11 1 13 4 4 9 9 4 4 2 12 9 1 12 9 1 13 4 9 1 12 12 9 13 4 14 1 9 1 9 1 9 1 13 2 1 13 2
17 9 1 13 4 9 9 1 9 1 13 4 1 13 9 1 13 2
41 9 1 13 2 9 1 0 9 1 0 9 1 13 4 4 9 4 4 2 15 1 9 1 9 1 13 4 1 13 4 9 1 13 9 1 13 4 1 13 4 2
44 9 1 13 16 2 9 11 1 12 9 1 9 2 12 12 9 9 1 14 9 1 13 4 11 9 11 9 1 9 9 9 1 1 9 9 1 2 9 2 1 13 16 4 2
30 10 9 2 11 9 1 9 1 13 4 4 9 9 1 1 9 1 13 4 9 9 9 9 1 13 4 4 16 4 2
5 15 1 0 4 2
39 7 2 9 1 9 1 13 4 9 7 9 9 1 13 4 1 13 9 9 1 13 16 2 9 9 1 1 9 1 13 16 3 12 9 13 4 16 4 2
37 9 5 11 9 1 9 9 9 1 1 9 1 9 1 13 2 11 9 1 9 9 1 9 9 1 1 9 9 1 13 1 13 9 1 13 4 2
22 9 2 9 1 9 9 1 9 9 1 13 2 9 9 1 9 1 13 4 4 4 2
13 9 1 1 2 9 9 2 1 9 1 13 4 2
14 7 2 9 1 9 1 0 13 2 9 2 1 9 2
37 0 4 9 1 11 1 9 1 13 2 9 4 9 2 1 13 4 4 9 1 9 1 9 1 13 4 16 4 2 1 13 16 9 4 4 4 2
12 3 2 11 1 3 13 16 4 4 16 14 2
19 9 1 2 9 1 9 9 1 13 9 9 2 1 9 13 4 16 4 2
47 9 1 9 9 1 13 16 2 2 9 1 13 9 2 1 13 9 1 2 9 1 0 9 2 1 13 4 9 1 12 12 12 12 9 2 9 9 1 13 16 12 12 9 1 13 4 2
34 2 11 1 0 4 4 9 1 13 16 4 14 2 1 9 1 1 2 0 9 2 1 13 4 9 1 12 12 12 12 9 13 4 2
27 9 9 1 9 1 2 9 1 13 16 4 4 9 1 13 9 1 9 1 13 4 4 16 4 4 4 2
17 0 9 1 9 9 1 0 4 13 4 16 4 16 4 4 14 2
12 0 16 2 9 2 1 13 4 1 13 4 2
20 9 9 9 14 2 0 4 0 9 1 3 13 16 9 9 1 3 0 4 2
26 11 9 1 9 9 9 1 1 12 9 1 13 16 2 9 1 13 16 4 1 13 9 1 13 4 2
21 9 1 9 1 13 2 9 1 9 9 1 13 16 3 13 4 9 4 16 14 2
12 9 1 9 1 13 9 1 13 4 4 4 2
16 2 9 1 13 9 9 1 0 2 1 13 4 1 4 14 2
14 9 1 9 1 3 13 4 4 4 16 1 4 4 2
4 7 13 4 2
25 3 2 9 9 1 9 1 13 4 4 9 1 13 16 2 9 9 1 9 1 9 1 13 4 2
32 9 9 1 11 9 2 9 1 12 9 1 13 4 11 9 9 1 9 1 13 4 2 12 9 1 9 9 1 13 4 4 2
25 9 9 1 1 13 2 15 14 13 4 9 1 9 9 1 9 1 3 0 9 13 4 4 4 2
15 9 1 13 4 16 2 3 9 9 1 13 16 4 4 2
11 9 9 1 13 9 1 0 9 1 13 2
15 9 9 1 13 9 9 1 9 1 9 1 13 1 13 2
38 12 9 1 13 4 9 1 9 1 13 4 16 2 9 1 9 1 0 4 13 9 1 9 9 9 1 13 9 1 9 1 0 13 4 16 4 4 2
21 9 1 9 9 1 15 9 13 4 16 2 11 9 1 1 9 1 13 13 4 2
24 11 11 2 11 11 9 9 9 9 1 9 9 1 13 4 4 16 1 2 3 9 1 0 2
17 7 2 9 9 1 9 9 1 3 9 9 1 13 4 16 4 2
12 9 9 1 1 9 9 1 10 9 0 4 2
15 9 9 1 13 16 1 9 1 13 16 4 1 13 4 2
32 9 1 0 9 1 1 13 2 12 12 12 9 9 1 9 9 1 13 14 1 2 10 9 1 9 1 13 16 1 0 4 2
19 7 2 9 9 1 9 9 1 9 1 13 4 14 1 1 13 4 4 2
23 2 9 5 9 9 2 2 9 9 2 1 9 9 4 4 2 9 1 0 9 4 4 2
10 9 4 16 9 1 9 1 13 4 2
8 7 2 3 1 13 4 4 2
42 3 9 1 2 9 9 9 9 9 9 2 1 13 9 4 4 2 9 9 7 9 9 1 9 9 2 9 9 1 9 1 9 1 13 9 9 1 9 9 4 4 2
34 9 5 9 1 9 2 9 9 1 13 4 2 9 9 9 1 1 9 7 12 9 9 1 9 9 1 13 16 1 0 9 1 13 2
12 12 9 1 0 9 1 13 16 4 4 4 2
42 15 14 14 2 9 1 9 9 9 1 9 1 9 1 13 2 9 9 7 9 9 9 2 9 9 14 2 0 4 9 1 13 4 4 9 9 1 13 16 4 4 2
63 12 9 1 9 9 9 1 9 9 1 2 9 9 1 13 16 1 2 9 9 1 9 2 1 13 4 2 9 9 1 13 16 1 2 11 9 1 1 13 4 16 4 4 2 2 9 1 9 9 1 13 4 2 1 9 9 1 13 9 1 13 4 2
34 7 2 9 1 9 9 1 9 4 1 13 16 1 9 1 13 16 2 9 9 0 9 1 0 0 9 2 1 13 9 9 1 13 2
42 9 9 1 9 1 9 1 9 9 4 16 2 9 1 9 9 1 9 9 1 13 16 4 16 2 9 1 9 9 1 13 4 0 9 1 0 1 13 16 4 4 2
50 2 0 9 9 1 13 4 4 9 1 13 4 4 2 1 11 11 9 1 13 4 4 4 16 2 9 2 9 1 9 9 5 9 1 13 16 9 9 1 9 1 13 4 9 1 3 13 4 4 2
7 9 1 9 1 1 4 2
28 9 9 1 13 16 2 9 9 7 9 1 9 1 13 4 16 1 2 15 14 9 1 13 4 4 1 13 2
22 9 9 1 13 4 16 9 9 2 7 1 9 9 1 9 1 14 13 16 4 4 2
16 3 2 9 1 9 9 1 9 1 13 9 1 13 4 4 2
11 9 1 9 1 13 9 1 1 13 4 2
38 9 9 1 13 9 7 9 2 7 1 11 9 9 9 1 9 9 1 9 4 4 11 14 1 13 4 16 9 1 13 4 2 9 1 13 4 4 2
34 9 9 1 1 9 1 13 4 9 1 1 2 9 9 5 9 1 3 13 16 4 4 15 14 1 9 1 1 9 1 3 13 4 2
26 9 9 9 9 1 9 12 9 4 4 12 12 9 9 9 1 9 12 12 12 9 1 13 4 4 2
23 13 16 12 12 12 9 9 9 7 12 9 9 9 1 12 12 12 9 1 13 4 4 2
9 15 1 9 12 9 1 9 9 2
27 9 1 9 9 9 2 9 9 2 9 9 2 9 9 9 1 9 12 12 12 9 1 9 9 4 4 2
28 9 9 9 1 9 12 12 9 9 1 1 13 16 3 2 9 2 1 9 1 13 4 4 16 4 16 4 2
41 3 9 9 1 9 9 9 12 9 9 1 13 4 2 9 9 9 1 13 16 13 9 1 11 2 11 2 11 2 11 2 11 1 13 16 1 9 1 13 4 2
49 7 2 7 12 9 1 9 12 12 12 12 1 1 9 9 9 1 9 12 9 9 1 9 12 12 12 12 1 9 1 9 1 13 4 9 4 2 11 9 1 9 9 1 13 4 9 1 13 2
60 9 9 1 3 13 4 4 16 4 4 16 1 2 9 9 1 1 13 12 12 9 9 9 9 9 1 9 9 1 9 4 4 2 9 1 9 9 2 7 3 0 4 9 1 13 4 1 13 4 9 9 1 13 16 13 4 9 4 4 2
42 9 9 1 9 2 9 9 1 13 16 1 9 9 1 2 9 9 9 2 9 7 2 15 1 9 1 9 9 13 16 4 9 9 1 1 2 9 2 9 4 4 2
64 10 9 3 1 9 9 9 1 9 9 1 9 9 1 13 16 13 4 2 7 11 12 12 9 1 9 9 1 9 1 9 1 4 4 13 16 2 13 16 9 9 1 9 9 9 1 13 4 14 9 9 7 9 9 1 9 1 13 4 4 16 4 4 2
14 15 1 9 1 13 16 4 16 4 16 1 9 4 2
79 15 1 9 9 1 9 9 9 1 9 9 1 9 9 13 4 16 4 4 9 1 1 13 2 3 9 9 1 9 9 1 13 9 1 9 9 13 16 4 4 9 2 9 9 14 9 9 1 13 4 2 7 9 1 1 9 9 4 9 9 7 9 1 1 15 1 0 4 1 9 9 13 4 9 1 9 4 4 2
51 7 2 7 9 9 1 9 9 9 1 3 2 9 1 0 9 9 1 13 4 2 1 13 9 1 9 1 9 1 13 4 4 2 9 1 15 1 13 4 4 4 16 4 14 1 1 4 4 4 14 2
18 3 9 9 1 9 9 1 13 4 2 9 9 1 9 9 1 0 2
31 9 9 1 1 9 9 1 9 9 4 9 9 9 1 9 1 9 1 13 2 3 9 9 1 9 1 13 4 16 4 2
24 9 1 2 9 1 0 2 13 4 9 2 1 9 1 1 9 1 13 9 1 1 4 14 2
24 9 9 1 9 9 13 9 1 9 9 1 9 9 1 1 9 1 13 9 1 9 0 4 2
31 9 1 9 7 9 1 13 4 4 9 1 13 16 4 9 1 9 9 1 13 16 0 4 9 1 13 4 4 4 4 2
38 10 9 1 9 9 9 1 0 9 1 13 16 4 9 1 2 9 9 1 1 9 7 9 9 1 13 16 4 9 9 9 9 4 9 4 4 4 2
27 9 1 9 1 3 9 13 4 4 4 16 1 2 11 9 1 9 1 0 9 1 13 4 9 4 4 2
59 11 9 1 9 1 9 9 1 9 9 9 1 9 1 13 4 9 2 9 14 9 9 1 0 9 9 1 9 1 0 9 1 13 16 4 2 9 9 9 1 1 9 7 9 9 9 1 13 0 9 1 13 4 9 1 13 4 4 2
50 11 9 1 13 4 9 13 9 1 9 9 9 1 9 9 1 13 16 4 4 16 1 9 1 9 1 9 4 16 2 15 1 13 9 1 12 9 1 13 9 1 9 1 0 9 4 16 4 4 2
34 11 9 11 9 1 9 9 9 9 1 13 4 4 4 9 1 2 9 9 1 9 9 9 5 9 1 9 9 1 9 9 13 4 2
34 9 9 9 1 13 4 4 9 1 13 1 13 9 1 2 9 9 1 9 9 9 1 12 9 1 9 9 1 13 16 4 1 13 2
27 12 12 12 12 9 1 9 9 2 9 9 1 13 4 16 4 2 15 1 3 13 4 9 1 13 4 2
21 9 9 1 2 9 4 9 9 4 4 2 9 9 4 2 1 13 4 16 4 2
9 9 1 3 13 4 16 4 4 2
20 7 2 9 9 1 1 0 4 9 1 9 1 0 0 4 13 16 4 4 2
34 9 1 9 1 9 1 13 4 16 1 2 9 9 1 9 1 9 9 9 9 7 9 9 9 1 9 9 1 9 13 4 9 4 2
9 15 1 9 1 13 4 9 4 2
19 7 9 9 9 1 9 9 1 1 9 1 13 4 4 2 1 1 13 2
17 9 1 9 1 9 9 1 0 4 9 1 13 4 16 4 4 2
28 11 9 1 9 9 1 9 1 1 9 9 1 9 9 1 13 2 9 9 9 9 1 13 4 4 16 4 2
20 9 9 1 1 9 1 9 4 4 2 9 1 9 2 1 13 4 4 4 2
38 9 1 1 2 12 12 9 1 2 9 9 9 2 1 9 1 13 4 4 4 9 9 1 9 1 9 1 13 4 4 4 2 1 13 9 1 13 2
18 10 9 9 1 2 9 9 2 1 13 16 15 14 0 4 13 4 2
22 3 4 4 16 1 2 10 9 1 1 12 12 9 9 1 9 9 1 13 16 4 2
21 9 1 9 1 13 9 1 9 5 9 1 9 1 9 1 13 16 13 16 4 2
20 9 9 1 9 1 9 1 0 4 3 13 4 4 16 4 4 4 4 4 2
20 9 1 9 4 4 9 9 1 9 12 12 12 9 2 11 9 1 13 4 2
26 3 9 1 0 9 12 9 9 2 9 9 1 9 9 1 12 2 12 9 1 9 1 13 4 4 2
32 2 13 16 2 1 13 3 1 9 1 1 13 4 2 0 12 9 14 1 9 1 9 9 1 13 4 16 9 1 13 4 2
23 9 1 9 9 1 9 1 9 1 13 4 9 4 2 0 9 1 13 4 9 4 4 2
21 9 9 1 9 1 9 1 9 1 9 1 13 16 9 1 13 4 2 1 13 2
24 9 9 1 9 9 1 13 4 4 9 4 2 9 9 1 1 9 9 1 13 16 4 4 2
28 9 1 13 16 2 12 12 12 12 9 9 1 11 9 1 13 4 9 9 12 9 9 9 1 9 1 0 2
10 10 9 1 3 9 1 0 1 13 2
12 15 1 15 1 9 1 13 4 4 16 14 2
7 10 9 1 13 4 4 2
13 7 9 1 11 1 1 9 4 9 1 0 4 2
22 9 9 9 9 7 0 9 2 9 9 14 9 9 1 13 4 4 4 9 1 13 2
14 10 9 1 9 1 9 1 13 4 16 4 1 0 2
13 9 9 1 15 1 13 1 13 16 4 4 14 2
12 3 9 1 13 4 4 14 1 1 4 14 2
14 9 1 9 9 1 13 4 9 1 3 0 4 4 2
13 7 2 15 1 13 4 4 9 1 3 0 4 2
12 9 2 15 1 13 4 16 9 1 13 4 2
20 9 1 9 2 0 9 1 9 9 1 13 1 9 1 13 16 4 4 4 2
20 11 5 9 9 9 1 9 1 9 4 9 2 9 1 13 16 13 4 4 2
10 9 9 1 13 16 1 9 4 4 2
34 10 9 2 9 1 2 9 2 1 13 4 9 1 13 11 4 16 2 9 9 1 1 2 9 9 2 1 9 1 3 13 16 4 2
12 10 11 1 9 1 9 4 13 4 16 4 2
5 0 4 4 4 2
16 9 1 9 1 9 2 13 4 4 1 13 4 16 4 4 2
17 9 9 1 9 1 9 1 3 4 13 16 4 4 16 4 4 2
25 10 9 1 2 9 1 12 12 12 9 0 11 1 9 1 13 4 9 9 9 9 1 13 4 2
16 9 9 1 2 9 1 13 4 9 1 13 4 9 4 4 2
34 12 12 12 9 2 9 1 9 1 13 4 9 1 9 2 9 14 0 9 9 9 1 9 1 2 9 9 1 9 9 1 13 4 2
8 3 2 3 13 4 16 14 2
13 9 1 2 9 1 0 4 4 1 13 9 0 2
28 9 12 12 9 1 9 2 9 9 1 13 11 9 9 9 9 9 1 2 9 9 1 9 1 0 13 4 2
17 9 9 1 13 16 9 9 1 9 9 1 13 4 16 4 4 2
20 9 1 9 1 13 2 9 9 1 9 1 0 4 9 1 13 16 1 0 2
7 3 13 4 16 4 4 2
16 3 9 9 9 4 4 9 1 13 4 4 9 4 4 4 2
28 3 9 1 13 16 1 2 0 9 1 13 9 1 2 9 1 9 1 9 1 13 4 9 9 9 1 13 2
11 15 1 9 1 9 9 1 9 4 4 2
14 3 2 9 1 9 1 9 1 13 4 1 13 4 2
13 9 1 12 12 9 9 1 13 4 9 1 9 2
22 9 1 9 9 1 9 1 9 1 13 2 15 1 9 1 13 4 4 9 1 13 2
33 9 1 9 1 9 2 9 12 12 2 12 12 9 1 9 2 9 2 11 1 9 9 1 9 1 9 1 13 4 1 13 4 2
13 10 9 9 1 9 4 9 1 13 4 4 4 2
7 9 1 3 4 4 14 2
10 9 2 9 1 9 9 1 13 4 2
26 11 1 9 5 11 1 9 12 9 1 0 12 12 12 12 9 2 12 12 12 9 1 13 4 4 2
17 11 9 1 9 1 0 2 9 9 1 13 16 9 1 13 4 2
8 15 1 9 1 9 4 4 2
11 9 1 11 9 9 1 13 4 16 4 2
26 9 9 1 9 1 2 9 1 13 4 4 4 2 1 13 9 1 13 4 2 1 13 4 16 4 2
36 9 1 9 1 13 9 9 1 13 4 4 16 1 2 0 9 9 1 9 1 13 4 4 4 2 13 4 16 2 1 13 9 1 13 4 2
26 0 4 9 4 16 1 2 9 1 9 9 9 1 2 10 11 9 9 1 2 13 4 9 1 13 2
26 9 9 14 1 9 1 2 9 9 14 13 4 16 2 9 9 1 1 12 9 1 13 4 4 4 2
17 15 1 1 9 9 1 9 13 2 1 13 4 4 1 13 4 2
13 9 1 9 1 13 4 9 1 1 4 16 14 2
15 9 9 1 9 1 9 1 13 4 4 4 4 16 14 2
16 0 4 9 1 9 9 1 13 4 1 13 16 1 4 4 2
25 9 9 1 1 4 9 9 1 13 9 9 2 7 9 9 9 9 9 9 1 10 9 4 4 2
14 7 2 9 9 9 1 9 9 1 13 4 16 4 2
18 9 1 13 4 1 1 2 9 9 14 1 13 4 16 1 0 4 2
21 9 1 9 9 1 13 4 14 1 9 9 2 9 9 1 0 4 16 4 4 2
31 9 1 9 1 13 2 9 1 9 9 9 1 1 13 4 16 4 2 9 1 10 9 1 9 1 13 4 16 4 4 2
17 9 1 9 9 1 0 16 1 2 15 1 9 9 1 13 4 2
16 12 9 9 1 13 4 2 9 1 9 4 9 1 13 4 2
24 0 9 9 2 9 9 1 9 1 13 9 1 9 4 16 2 9 1 9 1 13 16 4 2
26 15 1 2 9 1 9 9 7 9 9 1 9 1 1 2 9 1 13 16 13 4 4 9 4 4 2
13 3 9 1 2 9 1 3 1 9 2 4 4 2
11 9 1 9 1 0 2 9 1 3 0 2
11 2 9 9 2 1 7 13 4 4 4 2
4 9 1 13 2
17 2 9 1 9 9 2 4 4 2 9 1 9 1 0 13 9 2
29 9 1 9 12 9 9 1 13 4 4 9 9 1 1 2 9 1 13 9 9 1 9 9 1 9 1 13 4 2
11 15 1 9 1 12 9 9 9 4 4 2
15 9 9 1 13 16 13 16 2 9 9 1 0 13 4 2
24 10 9 2 9 1 9 4 4 9 9 1 2 9 9 1 12 9 1 0 9 1 13 4 2
12 3 11 9 9 1 12 9 1 9 4 4 2
14 9 1 13 16 1 3 9 1 9 1 13 16 4 2
26 9 9 9 9 1 9 4 4 9 1 2 9 1 3 9 9 1 13 1 13 16 4 1 4 14 2
40 0 9 9 1 9 1 13 4 16 2 9 9 1 9 1 9 9 1 9 9 1 9 1 12 12 12 9 1 12 12 12 9 1 1 3 16 13 4 4 2
28 9 1 9 9 1 9 9 9 9 1 9 1 13 4 4 9 4 16 2 9 9 1 12 12 9 1 0 2
20 15 1 12 12 9 1 13 4 16 2 9 9 1 12 12 12 9 1 13 2
23 13 9 1 13 16 2 3 3 0 13 16 4 2 1 13 16 1 9 4 9 4 4 2
41 12 9 9 9 9 1 9 9 1 12 9 9 1 2 1 13 9 1 13 16 2 12 12 12 9 9 1 9 1 13 9 1 9 1 13 16 4 1 4 14 2
18 10 9 1 13 1 1 2 3 9 1 9 14 1 9 1 1 4 2
22 9 1 9 9 1 9 2 3 9 7 9 1 13 9 9 1 9 4 13 16 4 2
23 9 1 0 9 1 13 9 9 1 2 9 1 9 9 1 13 2 15 1 9 1 13 2
31 9 9 9 1 9 1 2 9 9 1 13 16 9 9 1 9 9 1 0 9 1 13 9 1 3 13 4 16 4 4 2
39 12 12 12 12 9 1 9 1 13 4 11 9 1 9 9 1 2 9 12 12 12 9 14 13 4 16 2 9 1 12 12 12 12 9 14 13 4 4 2
11 15 1 3 9 9 1 9 1 0 4 2
19 7 9 1 3 0 4 9 1 13 16 4 4 2 1 13 9 1 13 2
19 0 4 2 15 14 1 9 1 13 16 0 11 1 13 4 9 1 13 2
29 7 2 9 9 1 12 12 9 9 1 9 9 1 3 9 9 4 9 1 13 16 4 4 1 13 16 3 14 2
31 7 2 9 9 1 9 9 1 0 9 1 13 9 9 2 9 4 9 1 13 4 14 2 1 13 4 9 1 13 4 2
19 3 9 9 7 9 9 1 9 1 13 4 4 2 1 1 9 1 13 2
15 15 1 13 16 1 2 9 1 9 1 3 13 16 4 2
20 9 12 1 2 9 9 4 13 16 2 11 1 9 1 9 1 13 16 0 2
17 11 1 9 12 9 2 11 1 9 12 9 1 13 0 9 4 2
17 15 1 3 2 11 1 13 9 9 1 9 9 1 13 16 4 2
26 9 12 1 2 10 9 1 9 1 9 1 0 13 4 16 4 4 2 9 9 2 1 9 4 4 2
30 9 7 9 1 9 9 1 9 1 13 16 2 9 9 1 9 1 9 9 1 9 1 13 4 16 4 4 9 4 2
33 7 2 9 1 9 1 9 1 2 9 1 11 9 1 9 1 13 16 4 4 9 1 13 16 4 1 13 16 3 4 4 14 2
13 2 9 1 9 2 1 9 1 2 3 0 13 2
5 9 1 3 0 2
42 11 9 9 9 9 12 9 1 9 9 1 2 12 9 12 9 9 1 12 12 12 12 9 9 1 13 16 4 16 2 15 1 9 1 9 9 1 13 4 16 4 2
13 15 1 9 9 12 9 9 1 9 1 13 4 2
17 11 9 1 1 9 2 12 9 5 12 12 9 9 14 13 4 2
21 9 9 1 9 7 9 9 1 9 1 13 2 9 1 1 9 1 13 16 4 2
25 9 1 9 1 13 9 1 1 2 9 1 13 16 9 0 9 1 9 9 1 9 1 0 4 2
31 7 2 9 9 1 11 9 9 9 1 9 9 1 9 1 13 4 4 4 2 9 9 9 9 1 9 1 13 16 4 2
11 7 2 9 9 1 9 1 15 1 13 2
21 9 9 1 9 9 1 13 1 13 16 4 9 1 9 1 13 4 4 16 4 2
14 15 1 9 9 1 9 1 9 1 3 0 13 4 2
42 9 11 9 2 9 1 12 9 1 9 9 1 13 9 1 2 9 1 9 9 1 1 9 1 9 1 13 2 9 9 1 9 9 1 9 1 9 1 13 16 4 2
29 9 1 9 7 9 9 1 9 1 13 13 9 1 9 1 13 2 9 1 9 1 13 2 9 9 1 13 4 2
21 9 1 9 1 13 4 16 4 16 2 3 1 9 9 9 1 13 4 16 4 2
28 9 1 9 9 1 12 12 12 12 9 9 14 13 4 12 12 12 12 9 9 1 13 2 3 0 4 4 2
10 7 2 15 1 13 4 4 16 14 2
22 9 1 9 9 1 0 9 1 13 4 4 2 9 1 9 1 3 3 1 13 4 2
14 7 2 9 9 4 0 9 1 0 9 1 13 4 2
20 9 9 1 13 16 1 2 12 12 9 1 9 9 9 1 9 9 1 13 2
13 9 1 13 2 9 9 1 1 9 1 13 4 2
28 7 2 12 12 9 9 1 9 9 9 1 13 2 9 9 1 12 9 9 1 9 1 9 1 13 9 4 2
29 9 2 9 9 7 9 9 1 13 9 7 9 1 9 1 13 2 9 1 9 1 0 13 16 4 9 1 13 2
13 9 9 1 2 9 1 3 0 13 4 9 4 2
9 15 1 1 9 9 1 13 4 2
44 9 1 9 9 1 9 9 9 1 9 1 13 4 16 2 9 9 1 13 9 1 13 16 2 9 9 1 13 4 16 2 9 9 9 9 1 9 9 1 13 16 1 0 2
17 3 2 9 9 1 1 9 1 9 1 9 1 13 16 4 4 2
35 9 1 12 12 12 12 9 1 9 9 4 9 9 1 13 2 15 9 13 16 2 15 1 9 1 14 9 1 9 1 13 9 1 13 2
41 7 2 9 9 9 1 13 4 11 1 2 11 2 11 9 9 9 1 9 9 1 9 12 12 9 13 16 4 9 9 1 13 16 2 9 9 1 3 3 0 2
31 13 4 16 2 9 9 1 11 1 9 1 9 1 9 1 13 16 2 9 9 1 9 1 13 9 1 13 14 13 4 2
21 9 9 2 9 9 1 9 1 13 4 4 16 2 13 4 9 1 0 4 4 2
18 7 2 9 9 1 13 16 1 2 9 1 9 5 9 1 0 4 2
20 9 1 9 9 14 9 9 1 9 1 9 1 0 9 1 13 4 4 4 2
29 9 1 9 9 1 1 9 1 13 16 2 9 9 5 9 1 9 1 2 9 1 11 9 1 9 1 13 4 2
23 9 9 9 9 1 9 1 13 9 1 9 14 2 9 9 9 1 9 0 9 4 4 2
28 2 13 4 4 2 1 9 1 2 9 13 4 9 12 12 12 9 9 9 9 9 1 11 9 9 1 13 2
23 11 1 10 9 1 9 1 9 9 1 13 4 4 16 1 2 11 9 1 9 4 4 2
29 2 9 9 1 13 2 9 1 9 9 1 13 4 2 1 9 9 1 13 9 4 16 2 3 9 1 9 4 2
26 13 4 4 9 1 13 16 2 12 12 12 9 1 9 9 1 2 9 1 13 4 9 9 1 13 2
24 0 9 7 9 1 9 1 3 2 13 4 16 2 9 7 13 1 9 1 13 14 4 4 2
21 9 9 1 12 9 4 16 2 9 9 1 12 12 9 1 1 13 16 1 0 2
19 9 9 1 13 1 9 2 12 12 9 9 1 9 14 0 9 1 13 2
6 9 9 1 9 4 2
28 3 9 1 0 16 1 2 9 9 1 9 1 13 4 9 2 9 2 9 9 1 12 9 1 9 9 4 2
10 9 1 9 1 9 1 13 4 4 2
28 9 1 9 9 9 1 2 3 13 4 16 14 2 9 9 1 15 14 13 4 4 16 4 4 14 2 1 2
12 12 9 1 9 9 9 1 0 4 13 4 2
15 11 1 12 9 2 9 1 12 9 1 9 1 13 4 2
10 9 1 9 1 9 1 9 9 4 2
18 9 1 13 2 9 9 7 9 9 1 9 1 13 4 9 1 0 2
12 3 1 9 14 4 1 4 4 1 9 4 2
10 7 2 9 9 1 9 1 0 4 2
23 9 9 1 13 2 9 9 9 1 9 1 9 7 9 1 9 1 9 9 1 13 4 2
20 9 9 1 13 4 9 1 0 9 1 9 1 11 11 9 1 13 16 4 2
32 2 9 1 13 16 2 13 9 1 9 1 0 9 1 13 4 4 2 9 1 11 9 1 9 1 13 4 9 1 13 4 2
15 0 9 1 13 4 4 4 2 9 1 9 4 4 4 2
25 9 1 1 9 1 13 16 2 9 9 1 1 13 4 2 1 9 9 1 9 1 13 16 4 2
11 9 9 1 13 9 1 9 13 4 4 2
20 10 9 1 2 9 1 13 4 9 1 2 13 4 9 1 3 1 13 4 2
15 9 9 1 13 4 9 1 9 1 13 1 13 9 4 2
19 13 16 2 9 1 1 9 9 1 9 1 9 1 9 1 13 16 4 2
8 9 1 9 9 1 3 0 2
10 9 9 1 1 9 1 13 16 4 2
28 9 1 9 1 2 9 9 1 13 15 1 1 3 9 9 1 1 4 1 13 4 9 1 0 4 16 4 2
27 9 9 1 9 14 9 9 1 9 1 13 4 9 9 1 2 9 9 1 9 9 1 9 1 1 4 2
35 9 9 1 9 1 2 9 9 9 1 0 9 1 9 9 1 13 16 9 5 11 9 1 9 12 9 1 9 9 1 13 16 13 4 2
17 9 1 9 12 9 1 2 9 9 1 9 1 9 9 1 13 2
6 11 9 1 9 4 2
15 9 1 9 1 13 2 10 9 1 13 4 9 4 4 2
20 7 2 9 1 9 1 9 9 1 13 4 1 1 9 1 1 9 1 13 2
29 9 1 13 4 10 4 4 9 1 9 1 1 2 9 9 7 9 9 1 1 0 4 9 1 13 1 13 4 2
13 9 9 1 9 9 9 1 13 4 4 16 0 2
35 9 1 9 1 13 16 1 9 1 13 9 1 2 12 9 1 9 1 13 9 1 1 2 9 9 1 9 9 1 13 9 1 1 4 2
16 0 4 2 13 4 2 9 1 9 9 1 1 4 4 14 2
18 9 9 1 9 1 9 0 4 9 1 13 2 9 1 9 4 4 2
73 2 0 9 9 1 3 9 9 1 13 4 16 14 2 9 7 15 1 9 9 4 16 2 13 4 4 9 2 3 2 3 1 13 4 16 9 4 9 1 13 16 4 16 13 4 2 7 0 16 9 1 9 1 13 14 0 2 9 9 1 13 9 1 15 9 1 9 1 0 4 9 4 2
35 9 1 9 9 1 9 1 9 9 9 1 13 16 4 4 11 11 9 1 0 9 1 9 1 13 16 2 9 1 0 4 13 16 4 2
17 11 9 7 9 9 7 1 9 1 12 12 12 12 9 1 13 2
58 9 9 1 9 9 1 9 1 9 1 9 9 1 9 4 13 4 4 16 1 9 12 12 9 1 13 4 4 4 2 9 1 9 1 9 2 1 13 2 1 2 9 9 2 1 9 1 13 4 9 1 2 9 2 1 13 4 2
40 9 2 9 12 12 9 1 9 1 13 16 13 4 16 13 4 16 4 4 9 1 2 12 9 1 9 2 1 13 16 1 2 9 1 9 2 4 4 4 2
18 12 12 9 1 1 3 9 1 2 9 9 9 9 2 1 13 4 2
24 2 9 9 2 1 9 9 9 1 9 1 13 4 16 4 4 9 1 0 9 1 13 4 2
35 9 9 1 9 1 13 4 9 1 2 9 1 13 4 4 9 9 1 9 9 1 13 16 9 9 9 1 1 9 1 0 13 4 4 2
92 9 1 9 12 9 9 9 9 9 1 9 1 9 1 9 9 9 9 1 9 9 9 1 13 4 4 9 9 9 9 9 9 9 1 9 1 9 1 13 4 9 2 11 9 1 9 1 9 9 1 9 1 13 9 2 9 9 2 9 1 13 16 2 9 9 1 13 9 9 9 9 2 1 13 2 2 9 9 2 9 1 9 1 13 2 9 2 9 1 13 4 2
34 9 1 9 1 12 12 9 1 9 1 9 1 13 9 14 9 12 12 9 1 13 16 9 9 9 9 1 13 4 4 16 4 4 2
46 10 9 2 9 1 12 12 9 1 9 9 2 11 2 11 2 11 2 11 1 12 9 1 9 9 9 9 9 1 9 1 13 4 16 2 15 1 9 1 0 9 1 9 1 13 2
38 12 12 9 2 9 1 13 4 16 13 4 4 4 9 11 1 11 9 1 9 1 2 9 9 2 1 9 1 13 4 4 1 13 9 1 13 4 2
64 11 9 9 2 9 1 9 9 9 9 1 13 4 16 1 2 2 9 9 2 1 13 4 9 1 13 4 16 2 9 4 9 1 9 9 1 9 1 13 16 9 9 1 9 9 9 1 13 9 1 13 4 9 9 1 9 1 13 4 4 9 4 4 2
67 9 9 1 9 9 9 1 13 9 9 1 9 9 1 13 1 13 4 9 9 9 9 1 13 2 12 9 12 9 9 1 9 9 9 9 1 9 1 13 4 2 9 9 1 13 4 9 9 4 2 1 13 16 1 9 9 9 9 9 1 0 4 9 4 4 4 2
72 7 2 9 9 9 9 1 9 1 13 4 2 9 9 2 1 9 1 13 4 16 1 10 12 9 12 9 1 9 1 9 1 13 16 2 0 9 9 1 9 1 9 1 9 1 9 9 1 13 4 4 16 14 3 14 2 3 0 13 16 4 16 4 16 1 9 1 1 4 4 14 2
49 9 9 9 9 9 1 9 1 13 4 9 9 9 1 2 9 9 9 1 9 9 9 1 9 1 13 4 9 9 9 9 1 9 1 0 13 2 9 1 9 1 9 1 13 4 4 16 4 2
29 9 1 1 9 9 1 9 9 1 13 16 0 1 9 3 1 0 9 1 9 1 13 4 4 16 4 1 13 2
50 9 9 2 9 9 1 9 1 2 9 2 9 1 9 1 9 1 13 16 1 9 9 7 9 9 1 13 4 9 1 2 9 9 1 9 9 1 13 4 2 9 1 9 9 1 13 4 9 4 2
42 12 9 9 1 1 9 1 2 9 12 9 1 9 9 1 1 13 16 2 9 4 0 9 1 9 1 13 11 9 9 9 1 9 9 9 1 9 1 13 16 4 2
58 15 1 1 0 16 1 2 9 9 9 9 9 1 9 2 9 2 9 9 1 9 1 9 9 9 9 1 14 13 16 9 1 9 4 4 9 1 0 4 13 2 9 9 1 13 4 16 9 9 1 9 1 13 16 4 9 4 2
33 9 1 9 13 4 4 9 9 1 1 2 2 9 9 0 2 1 12 12 9 1 13 2 9 9 3 12 12 9 1 13 4 2
37 9 1 9 9 1 13 2 12 9 9 1 9 1 13 16 13 4 9 9 1 9 1 2 3 0 9 9 1 9 1 1 9 1 9 4 4 2
19 13 4 4 2 9 9 9 2 1 3 13 16 9 9 1 13 16 13 2
28 2 9 9 0 2 1 1 13 9 2 9 1 9 9 1 9 4 4 2 9 1 9 9 1 9 4 4 2
36 9 1 9 1 13 9 1 13 4 4 9 1 0 4 13 4 16 2 9 9 9 1 9 9 9 1 9 1 13 9 9 0 1 13 4 2
16 9 9 1 9 1 9 1 13 4 4 0 4 9 4 4 2
22 9 1 13 16 3 13 9 1 9 1 13 4 4 16 4 4 16 1 3 4 4 2
31 3 9 1 9 1 2 9 2 1 0 13 4 2 9 1 0 4 9 1 9 1 13 16 0 4 13 4 4 4 4 2
36 9 9 9 9 1 9 1 13 4 4 2 2 9 9 9 2 1 13 4 9 1 2 9 12 12 9 9 1 9 9 9 1 13 4 4 2
54 9 9 2 9 9 1 13 16 0 4 9 1 13 9 4 4 9 4 16 2 9 2 9 2 9 2 9 2 9 9 5 5 14 2 9 2 1 9 1 13 9 1 13 4 16 4 16 1 0 9 4 4 14 2
14 9 9 1 9 9 9 1 12 9 1 13 16 4 2
45 9 1 9 9 1 1 2 10 9 9 1 9 1 13 4 9 1 9 1 2 9 1 1 9 1 9 14 1 2 9 1 13 2 9 9 9 2 1 9 1 3 13 16 4 2
51 9 1 2 9 1 9 1 9 1 13 9 1 1 13 4 2 2 9 1 9 1 13 4 16 2 14 1 13 4 16 2 9 1 9 1 9 9 9 1 2 9 1 3 9 1 9 1 13 16 4 2
5 10 9 1 0 2
59 12 12 12 9 9 9 1 12 12 12 9 1 13 4 4 16 2 9 1 9 1 1 2 9 9 9 1 9 1 9 9 1 13 9 9 1 9 9 4 2 9 1 12 9 9 1 9 9 1 13 9 1 0 13 16 4 1 13 2
58 9 1 9 9 1 13 2 0 4 9 1 9 1 13 16 2 9 1 9 1 13 9 9 1 13 16 4 4 16 2 9 9 9 1 9 9 1 13 16 13 14 9 1 9 1 13 2 9 1 13 16 9 9 1 9 1 13 2
18 9 2 9 9 9 1 9 9 1 9 1 13 9 1 13 16 4 2
29 3 13 16 4 16 2 9 9 9 1 13 9 1 1 9 9 1 13 16 4 16 4 1 13 4 1 13 4 2
27 9 1 2 9 7 9 2 1 13 9 1 13 2 9 9 1 13 4 4 4 16 1 0 4 4 4 2
23 9 9 1 9 9 1 9 7 9 1 9 1 9 1 13 4 9 1 13 4 4 4 2
37 9 1 9 9 1 3 13 14 1 13 16 1 2 12 12 12 12 9 1 9 9 9 9 9 7 9 9 7 1 9 1 9 9 1 13 4 2
85 9 9 1 9 9 1 1 9 1 2 9 1 9 1 9 7 9 1 3 5 9 9 1 13 4 4 1 13 4 4 16 9 2 9 1 2 9 9 1 9 1 13 16 3 9 9 4 9 1 13 16 4 4 2 7 9 1 9 9 4 9 1 13 16 0 4 9 9 13 4 4 9 9 1 9 9 1 13 4 4 2 16 4 4 2
39 9 9 4 9 9 9 1 13 16 1 2 9 2 9 1 9 9 9 7 2 9 1 9 7 9 1 9 1 13 9 1 13 9 9 14 1 13 4 2
26 9 2 9 9 9 1 13 4 4 4 12 12 9 9 1 9 12 9 9 9 9 1 13 4 4 2
22 13 4 4 16 1 9 1 9 1 13 2 9 1 9 1 13 1 13 9 4 4 2
7 15 1 12 12 12 9 2
33 9 9 1 9 9 1 9 1 0 9 1 13 4 4 16 2 9 9 9 1 9 1 9 9 4 9 1 3 13 16 4 4 2
51 13 4 16 4 1 13 16 2 15 14 4 16 2 9 1 13 16 2 9 9 9 1 9 1 13 4 9 1 9 9 9 1 9 1 9 1 9 1 13 9 1 13 16 4 1 1 9 1 0 13 2
36 10 9 9 9 9 1 2 9 9 2 7 2 9 1 9 9 9 1 12 12 9 1 9 12 12 9 9 9 9 9 1 9 9 4 4 2
41 9 1 13 16 2 9 9 1 9 2 1 13 4 2 10 9 1 9 9 13 16 9 9 1 13 9 1 1 9 4 16 2 9 1 13 9 4 13 16 4 2
49 9 9 9 1 1 9 9 9 1 9 9 1 13 16 9 1 9 2 2 9 9 1 13 16 2 9 9 1 1 9 9 1 13 4 16 1 9 1 13 4 2 1 1 9 1 3 13 4 2
33 9 9 4 1 11 9 1 3 9 9 9 1 13 2 11 9 9 9 9 1 1 9 9 9 1 9 9 1 13 4 16 4 2
46 9 1 1 9 1 9 9 2 9 1 9 9 9 9 1 9 1 9 9 1 13 4 4 1 1 9 9 1 13 4 9 9 1 13 2 3 12 12 12 12 9 1 13 16 4 2
27 10 9 1 11 1 9 9 7 2 9 1 13 4 16 4 9 1 1 9 9 9 9 13 4 16 4 2
17 13 4 16 9 9 1 13 9 1 13 9 1 13 9 4 4 2
19 9 2 9 1 9 9 1 13 0 4 9 9 1 13 4 4 4 4 2
32 10 9 9 9 1 3 9 9 4 4 9 1 0 1 1 9 1 2 9 9 9 1 13 4 4 4 1 1 9 1 13 2
29 9 9 1 9 9 1 9 2 13 4 9 4 16 2 9 1 9 9 1 13 16 1 9 1 13 9 4 4 2
15 3 9 1 13 14 4 16 4 1 13 9 4 1 4 2
22 7 9 9 1 13 16 9 1 9 1 9 7 9 1 9 1 13 9 1 0 4 2
36 9 1 9 7 9 1 9 1 13 2 9 7 9 1 9 9 1 13 9 1 9 1 13 4 9 9 1 13 4 4 1 13 9 4 4 2
32 9 9 1 13 9 1 13 9 1 13 2 9 9 1 13 4 4 2 9 9 4 13 16 4 9 1 13 4 16 4 4 2
24 11 9 11 9 1 13 9 1 9 1 13 9 1 2 9 9 1 9 9 9 1 13 4 2
19 9 1 9 1 0 4 9 1 13 4 9 1 13 1 13 16 4 4 2
13 15 14 1 9 1 9 1 9 1 13 16 4 2
28 10 9 1 12 12 1 12 12 9 1 1 13 2 9 9 5 9 1 9 9 1 13 16 4 4 1 13 2
11 0 4 9 9 1 13 16 4 4 4 2
15 9 9 1 0 4 4 13 4 1 13 16 4 4 14 2
50 9 9 1 3 13 4 2 9 1 9 2 2 9 9 1 13 9 2 2 9 9 1 9 9 1 13 16 4 2 14 1 13 4 16 4 1 13 16 2 9 9 1 0 1 13 4 1 13 4 2
24 9 9 9 1 2 9 1 13 9 1 9 7 9 14 1 13 4 4 9 1 13 4 4 2
27 9 1 9 1 1 2 9 1 9 9 9 1 9 1 13 4 4 1 13 9 9 1 13 16 4 4 2
40 7 2 9 9 9 1 9 1 0 9 9 1 9 1 0 9 1 13 4 4 9 2 13 4 4 1 13 9 4 2 9 9 9 1 1 9 1 13 4 2
18 9 1 9 4 4 2 9 2 9 9 1 9 9 1 13 4 4 2
8 9 1 13 9 1 3 13 2
22 9 2 9 9 2 9 14 1 9 1 9 1 9 1 9 1 9 1 13 16 4 2
9 9 1 9 1 13 9 1 13 2
14 9 9 4 4 16 1 9 9 1 9 1 13 4 2
22 9 9 1 13 4 9 1 13 16 0 4 9 1 13 4 4 4 16 1 4 4 2
6 15 14 1 1 4 2
20 9 9 9 9 1 9 9 1 1 2 3 9 1 9 1 13 16 4 4 2
19 11 9 9 7 9 9 9 1 13 0 9 1 9 9 1 9 4 4 2
16 9 9 1 9 1 0 4 0 4 13 4 16 1 4 4 2
14 9 4 13 4 16 4 9 1 9 1 15 1 13 2
33 7 2 13 4 4 16 1 9 9 5 9 1 0 9 4 4 2 12 9 9 2 1 9 1 9 4 13 4 1 13 9 4 2
32 9 9 1 2 9 1 9 2 1 1 13 4 2 3 9 1 9 1 9 1 12 12 9 1 2 3 0 9 9 1 13 2
33 12 12 9 14 9 1 11 1 13 4 4 4 16 2 9 12 9 9 9 1 1 9 1 13 4 4 1 1 13 4 16 4 2
35 9 1 9 1 12 9 9 1 3 9 1 13 4 4 1 13 4 16 2 12 12 12 9 9 1 1 9 9 1 13 4 4 4 4 2
11 13 4 4 14 1 9 1 9 1 13 2
29 9 9 4 13 4 4 2 12 9 9 1 2 9 1 13 9 1 13 2 1 13 9 1 13 1 4 4 14 2
23 9 1 13 9 9 1 9 9 9 9 1 9 1 9 1 13 4 4 9 1 13 4 2
17 15 1 2 9 9 2 1 0 9 1 9 1 9 1 13 4 2
15 9 7 9 9 1 9 1 1 4 4 16 2 9 0 2
29 9 9 9 1 13 4 16 9 14 9 9 9 1 9 2 9 1 13 4 9 1 9 9 1 13 4 9 4 2
30 3 0 4 9 4 16 2 15 14 1 1 9 9 9 1 9 9 1 13 16 1 3 9 1 13 4 16 4 4 2
12 0 4 16 1 2 10 9 1 1 9 4 2
38 9 9 1 0 4 4 2 12 9 9 14 9 1 9 9 1 13 9 1 9 1 9 5 9 13 2 3 0 9 1 13 4 16 4 1 4 14 2
15 9 1 9 9 1 9 9 4 0 9 1 13 16 4 2
17 9 1 13 4 16 2 9 9 1 9 9 1 3 13 4 4 2
30 9 0 9 1 9 1 13 4 14 12 12 12 9 1 9 12 9 14 11 1 9 1 2 9 9 2 1 13 4 2
36 12 12 12 12 9 1 9 9 1 13 4 4 4 2 9 9 9 9 2 1 1 12 12 12 12 9 1 13 2 9 9 1 13 4 4 2
48 9 1 9 9 1 2 9 7 9 1 13 16 13 4 9 1 9 9 9 9 1 2 12 12 12 12 9 1 9 7 15 9 1 12 12 12 12 9 1 9 1 13 4 2 13 16 4 2
36 9 9 1 9 11 2 11 14 9 9 12 12 9 1 9 2 9 14 0 9 9 1 0 4 4 9 1 13 14 9 9 1 13 4 4 2
28 3 9 9 4 2 11 1 12 12 12 12 9 1 12 12 9 1 1 12 9 14 9 9 1 13 9 4 2
28 7 2 9 1 0 9 9 1 9 9 1 9 1 13 9 9 9 1 9 13 9 0 1 9 1 13 4 2
38 11 9 1 12 12 9 1 9 9 1 9 1 2 9 9 9 1 15 9 1 9 9 1 12 12 9 2 9 9 1 1 12 12 9 1 13 4 2
32 9 1 9 9 1 9 12 12 9 1 13 16 2 9 1 9 9 1 9 9 1 12 12 12 9 1 13 16 4 9 4 2
35 11 12 12 12 12 9 2 9 11 12 12 12 12 9 2 11 1 12 12 12 12 9 1 13 2 11 1 9 9 1 0 9 1 13 2
29 15 1 9 1 2 11 1 3 13 4 9 1 13 4 2 1 9 1 9 1 9 9 4 9 1 9 9 4 2
13 7 2 9 9 4 13 4 9 1 1 4 4 2
35 9 1 9 9 9 1 13 9 1 9 11 1 12 9 2 9 11 1 12 12 12 9 1 13 11 12 9 1 12 12 12 9 1 13 2
20 9 9 1 9 12 9 1 9 1 9 9 1 13 16 1 3 0 4 4 2
24 0 9 1 9 1 13 4 4 2 9 1 13 4 16 4 9 1 0 4 9 1 13 4 2
24 9 9 4 9 9 1 10 12 12 9 1 11 1 13 4 4 9 1 9 1 0 4 4 2
22 9 9 1 13 4 16 4 9 1 3 9 1 12 12 9 1 1 9 9 1 13 2
36 9 9 1 9 1 13 4 4 16 2 11 1 9 1 9 9 9 1 12 12 9 2 9 9 12 12 9 1 9 1 13 4 16 4 4 2
11 10 9 1 9 1 13 16 1 3 4 2
41 11 9 1 13 11 7 9 1 9 9 9 1 2 9 9 1 9 9 1 9 1 13 9 1 13 14 9 1 13 16 1 9 2 1 13 16 4 16 1 13 2
39 11 1 0 9 9 1 9 4 1 13 9 1 13 16 2 9 1 9 1 13 4 16 4 4 2 9 9 5 11 2 1 9 1 13 4 9 4 4 2
13 10 9 1 9 1 0 4 9 1 13 16 4 2
61 11 14 12 12 12 1 9 9 9 1 0 9 1 13 9 9 1 9 1 2 9 2 13 9 1 13 1 13 16 2 9 9 1 2 12 12 12 12 9 14 1 9 1 9 9 1 12 12 9 9 1 12 12 9 13 4 2 13 16 4 2
50 7 11 1 9 1 2 9 9 1 9 7 9 14 9 0 4 9 1 13 2 3 9 9 1 13 2 12 12 12 12 9 9 1 9 1 9 9 1 9 9 13 9 1 9 9 9 1 13 4 2
50 12 12 9 1 13 9 1 9 9 1 13 4 2 9 9 1 13 9 9 9 2 1 0 9 9 1 13 2 9 1 0 0 9 1 1 9 9 1 13 4 2 9 1 9 9 1 13 4 4 2
34 9 4 9 9 9 1 13 13 16 2 9 5 9 9 1 9 1 13 9 9 1 2 3 9 9 9 1 1 13 16 4 16 4 2
27 11 1 13 4 16 4 9 9 1 13 2 9 1 13 4 9 9 1 9 9 1 13 4 16 4 4 2
19 12 9 1 9 1 13 4 9 7 9 7 1 9 1 9 1 13 4 2
29 9 1 9 1 13 16 1 2 9 2 11 9 1 13 4 16 9 11 9 1 13 4 16 9 1 9 1 13 2
29 9 2 9 1 11 11 9 1 2 9 1 13 4 4 2 9 13 9 1 0 4 2 1 13 4 16 4 4 2
17 9 1 9 1 2 9 9 1 13 16 9 13 9 4 4 4 2
18 9 1 13 3 9 1 0 9 14 4 4 2 0 4 9 1 13 2
36 3 9 1 9 1 9 1 13 4 9 4 2 9 9 1 9 9 1 0 4 16 2 9 1 1 9 1 9 9 1 13 4 9 1 13 2
22 11 1 9 9 7 11 1 9 9 1 13 4 9 9 1 9 9 1 13 4 4 2
27 9 1 9 1 13 16 14 13 4 16 2 15 1 13 16 9 9 9 1 13 4 9 5 9 1 13 2
21 9 9 1 9 3 13 16 2 9 1 9 1 13 4 4 16 1 9 4 4 2
16 9 1 9 9 2 9 1 9 9 1 9 1 13 16 4 2
17 11 1 9 9 9 1 13 9 1 1 12 9 1 9 1 13 2
59 9 1 9 5 9 9 7 1 9 4 2 11 1 13 4 4 9 9 0 9 1 9 4 2 9 9 1 9 1 13 4 16 2 9 1 0 4 0 1 9 9 1 13 4 16 2 9 9 7 9 1 9 1 9 1 9 1 13 2
28 13 4 4 16 1 2 9 1 9 9 1 10 9 1 13 4 4 16 2 0 4 4 9 1 13 14 4 2
18 9 9 1 13 4 16 2 9 9 1 9 9 1 3 13 16 4 2
26 7 2 15 14 1 9 1 9 9 1 9 1 13 16 2 9 1 9 1 13 9 1 0 4 4 2
44 9 1 9 4 2 9 9 9 1 9 9 9 1 13 16 4 2 10 9 11 1 9 1 9 1 13 16 9 1 9 1 13 2 9 1 9 1 0 9 1 13 16 4 2
23 15 1 9 1 13 16 2 3 9 9 13 2 9 1 0 4 13 9 1 13 4 4 2
21 9 9 1 9 1 9 1 9 1 13 9 2 9 9 1 13 4 16 4 4 2
16 9 9 1 13 16 2 9 7 9 1 1 9 9 1 13 2
15 3 1 9 16 2 3 9 9 9 1 9 1 13 4 2
24 7 2 9 1 9 1 9 9 1 9 1 13 2 9 9 1 9 9 4 13 4 4 4 2
13 9 1 1 0 4 9 1 3 13 4 4 4 2
26 3 2 9 9 1 9 1 1 2 9 4 9 1 9 1 13 4 2 9 1 13 4 16 4 4 2
20 9 9 1 12 9 1 9 1 9 1 9 1 13 2 9 1 13 16 4 2
34 9 1 0 9 13 4 12 12 12 12 9 9 1 9 1 2 9 9 4 9 1 13 16 2 3 9 1 13 16 4 4 4 4 2
23 9 1 4 4 9 1 9 9 1 13 16 4 4 4 16 2 9 9 1 3 13 4 2
29 9 9 1 9 9 1 3 1 9 9 9 1 2 9 1 9 9 1 9 1 12 9 12 9 14 13 16 4 2
24 15 1 3 9 9 13 4 2 9 1 9 1 9 9 13 16 4 14 1 9 1 9 4 2
25 11 2 9 1 0 4 9 1 2 11 1 9 9 7 9 1 9 9 1 13 9 1 13 4 2
37 9 1 1 9 9 1 2 9 7 9 1 3 0 9 1 13 16 1 2 9 9 9 9 1 11 9 9 9 1 13 4 9 4 4 1 13 2
30 9 9 9 1 13 16 2 11 1 9 1 9 1 3 13 4 4 9 1 13 2 9 1 9 1 13 9 1 13 2
11 7 2 9 9 1 3 0 9 1 13 2
49 11 1 11 1 13 4 16 4 4 9 9 1 9 9 1 13 9 9 1 2 9 1 9 1 13 16 12 12 12 9 13 4 4 16 1 2 11 1 0 9 9 1 13 4 9 4 4 4 2
31 11 1 2 9 9 1 9 12 12 12 9 14 1 9 9 1 13 4 9 1 9 9 1 13 4 1 13 4 16 4 2
22 9 1 13 4 16 4 16 1 2 2 11 9 9 2 1 9 1 13 9 4 4 2
17 9 9 9 11 1 2 11 9 2 9 1 11 1 13 16 4 2
19 7 2 11 1 2 11 9 1 13 9 1 0 2 1 13 4 16 4 2
17 9 9 9 1 9 1 2 9 9 1 9 9 9 9 1 13 2
26 9 9 1 1 2 13 4 4 9 1 9 7 9 1 13 16 9 9 4 9 1 13 4 4 4 2
15 11 1 2 10 2 9 2 1 0 13 16 4 9 4 2
41 9 9 9 9 1 13 16 2 11 9 9 1 9 1 13 9 1 13 14 2 9 9 1 13 4 4 9 4 4 16 2 11 9 1 9 1 13 4 1 13 2
27 9 1 2 9 9 1 9 9 9 1 9 1 9 9 4 9 1 9 1 13 16 4 4 16 4 4 2
21 9 9 1 9 1 9 4 4 9 2 11 1 9 1 3 0 1 1 13 4 2
27 11 1 2 11 9 2 1 13 16 2 11 1 9 9 13 4 16 1 3 13 4 4 9 4 4 4 2
38 3 9 9 9 11 1 2 2 11 9 2 9 1 13 16 13 14 2 11 1 0 4 2 9 9 2 1 13 1 13 9 4 9 1 13 16 4 2
37 9 1 1 2 9 2 1 13 4 4 9 1 9 9 1 13 16 2 2 11 9 2 1 13 2 9 1 9 2 1 9 1 0 4 1 4 2
19 9 9 7 9 9 0 1 1 2 9 1 9 1 13 4 4 16 4 2
20 11 1 2 9 9 1 13 4 9 1 10 9 1 13 4 9 4 4 4 2
36 11 1 2 3 11 1 9 9 9 1 13 4 4 4 9 1 13 16 2 11 9 1 1 9 1 13 1 1 9 1 0 4 13 16 4 2
19 10 9 1 1 2 9 9 7 9 9 1 13 0 9 1 9 1 13 2
15 11 1 2 11 1 9 1 9 1 9 13 4 4 4 2
35 11 11 9 9 9 5 9 1 9 1 13 9 12 9 9 9 1 2 12 12 12 9 1 9 9 9 9 9 9 9 1 13 4 4 2
46 7 9 9 9 1 13 4 2 9 9 1 9 1 13 4 9 9 1 1 9 9 9 9 9 1 2 9 9 9 1 9 1 13 4 16 4 9 1 13 4 16 4 4 4 4 2
39 9 9 9 9 9 9 1 9 1 13 16 1 2 9 9 1 9 7 9 9 9 1 9 1 0 9 1 13 4 4 4 2 9 4 9 1 13 4 2
68 9 1 13 9 1 9 1 2 9 9 9 9 1 1 9 9 1 9 1 0 4 13 4 9 1 9 1 13 16 4 16 2 11 9 9 7 11 11 5 9 12 9 9 1 13 9 9 9 9 1 13 4 2 9 1 9 9 4 9 7 9 1 9 1 13 16 4 2
18 2 9 1 13 9 1 1 2 9 1 9 9 1 13 4 4 4 2
15 11 9 1 11 11 9 1 9 9 1 13 4 9 4 2
37 9 2 11 9 1 9 9 1 1 2 9 1 13 4 4 16 2 9 1 9 7 9 1 9 9 1 13 9 1 3 12 12 9 9 1 13 2
15 9 9 2 9 9 1 9 9 9 1 9 9 4 4 2
14 9 9 1 0 4 9 1 2 9 1 9 4 4 2
29 9 9 1 3 13 4 16 1 2 9 1 9 1 9 1 13 4 4 9 1 1 2 9 1 9 1 13 4 2
16 9 2 9 1 2 9 9 12 2 1 1 9 1 13 4 2
38 9 9 1 9 9 1 2 9 12 9 9 1 13 16 2 12 12 9 1 9 1 9 1 4 4 9 1 13 16 4 16 1 9 4 9 4 4 2
22 9 9 9 1 13 4 2 9 1 9 2 1 0 4 4 1 13 4 1 13 4 2
21 9 1 13 16 2 9 4 9 9 1 9 7 9 1 9 14 9 12 12 9 2
13 15 14 1 9 9 1 13 4 4 4 14 4 2
17 9 9 1 9 7 9 9 7 9 9 1 9 1 9 1 13 2
9 9 1 0 9 1 13 4 4 2
40 9 1 13 16 1 2 9 9 1 1 9 9 1 9 1 9 5 9 9 1 13 4 2 9 9 1 13 4 4 16 1 9 1 0 9 9 1 13 4 2
17 9 1 13 14 1 9 1 13 14 2 0 4 9 1 13 4 2
14 13 4 16 13 4 4 9 1 12 12 9 9 13 2
18 9 1 0 9 9 1 13 16 13 16 4 16 2 3 4 16 14 2
47 2 0 16 9 1 9 1 0 2 13 4 9 7 9 1 9 1 13 4 2 2 9 9 1 9 1 2 9 7 9 1 9 1 1 3 0 4 9 14 2 14 1 9 9 1 13 2
13 9 9 1 9 1 9 1 13 9 1 13 4 2
15 10 9 9 1 9 1 2 9 2 1 13 9 1 0 2
13 0 4 9 13 16 1 9 9 1 9 4 4 2
39 11 9 11 9 1 1 9 1 9 9 1 12 12 9 9 14 13 4 4 2 3 12 12 9 1 13 9 9 1 0 1 1 9 1 13 4 16 4 2
48 9 9 1 2 9 9 1 3 9 9 1 2 9 9 1 9 7 9 14 1 13 4 16 9 12 12 9 1 9 1 0 2 1 2 9 1 13 9 9 1 13 16 9 1 13 4 4 2
25 9 9 7 9 9 1 0 9 9 4 4 2 0 9 1 0 13 4 9 1 0 4 9 4 2
34 9 9 7 9 9 1 9 1 1 2 9 1 9 9 1 13 2 9 1 1 9 1 13 4 9 9 9 9 1 13 9 1 0 2
19 9 1 9 7 0 9 1 2 9 9 9 1 0 13 4 9 1 13 2
36 9 9 4 9 7 9 9 2 9 9 4 9 1 1 9 9 14 2 9 9 12 2 1 9 1 1 9 9 4 9 1 13 4 16 4 2
19 9 9 1 9 9 1 9 1 0 0 4 9 1 13 9 1 0 4 2
25 9 1 13 16 14 13 4 16 0 4 16 14 2 0 9 7 9 9 1 13 4 4 16 14 2
14 13 13 16 9 9 9 1 13 9 1 13 16 4 2
17 12 9 1 13 9 9 1 2 9 1 1 9 1 13 4 4 2
11 9 9 1 13 4 9 9 1 0 4 2
23 9 1 9 1 13 2 9 1 9 9 1 9 14 1 9 9 9 1 13 9 1 13 2
6 9 1 13 14 4 2
48 11 9 1 9 2 9 9 9 1 9 1 9 13 2 9 1 13 4 16 2 3 9 1 13 4 9 9 14 1 1 2 9 1 9 1 9 9 1 13 4 4 16 4 9 1 13 4 2
10 9 9 1 9 1 13 4 4 4 2
18 9 9 9 1 1 2 7 1 9 5 9 9 1 1 13 4 4 2
13 2 9 9 2 1 9 1 13 4 0 9 4 2
7 0 4 9 9 1 13 2
17 3 4 4 16 2 0 2 0 9 1 9 2 9 1 13 4 2
36 11 11 5 9 9 1 9 1 12 12 9 9 2 9 1 9 9 9 1 13 4 9 1 2 9 1 12 9 13 4 2 9 1 13 4 2
17 13 4 9 1 13 4 1 13 9 1 13 2 9 1 13 4 2
19 9 1 13 4 9 1 13 16 4 4 16 2 9 9 1 13 4 4 2
7 9 1 9 1 13 4 2
37 9 9 9 1 1 2 9 1 13 9 9 1 13 11 5 11 1 2 9 2 1 13 11 1 13 2 9 9 9 1 9 9 4 4 1 13 2
27 7 2 3 3 1 0 4 13 4 16 4 4 16 14 2 1 13 16 1 9 9 1 13 4 9 4 2
26 9 9 1 1 9 1 9 9 4 4 2 10 9 1 9 9 1 9 9 1 10 9 1 13 4 2
15 9 1 0 1 13 9 1 13 4 4 1 1 13 4 2
17 7 2 9 1 9 9 2 9 9 1 1 9 1 13 4 4 2
6 9 1 13 4 4 2
12 9 9 1 9 1 9 1 13 4 16 4 2
20 11 9 1 9 7 9 9 1 13 9 1 9 9 4 13 4 16 4 4 2
18 9 9 9 1 1 9 1 9 9 1 13 2 0 4 13 16 4 2
35 7 2 9 1 1 9 9 9 7 11 9 9 2 7 1 9 9 1 9 1 1 9 1 9 9 9 1 13 16 13 4 16 4 4 2
25 0 7 9 4 9 1 9 1 13 9 1 9 1 9 1 13 9 7 9 1 0 1 4 4 2
19 9 1 9 1 3 13 4 14 1 2 9 1 9 1 1 3 0 4 2
19 7 9 9 1 1 4 2 9 1 1 9 1 13 4 9 1 13 4 2
26 11 4 4 9 2 9 9 1 2 9 2 1 13 9 1 0 2 3 9 1 1 13 9 1 13 2
17 7 2 3 1 13 4 4 2 9 2 1 13 4 4 4 13 2
16 15 1 13 4 16 4 16 1 9 1 9 1 1 4 14 2
15 9 1 9 9 2 9 9 1 10 9 1 1 4 14 2
24 2 9 1 9 4 9 2 1 2 9 1 9 4 9 2 1 13 4 4 14 1 4 4 2
15 3 1 15 1 13 14 2 15 1 1 9 1 13 4 2
8 7 9 1 9 1 13 4 2
10 9 1 9 9 4 13 4 9 4 2
18 2 3 2 1 1 4 13 16 9 9 1 10 9 1 13 16 4 2
7 9 9 1 1 13 4 2
11 15 14 1 2 1 13 16 4 1 4 2
18 9 12 9 2 9 1 13 0 9 1 13 4 4 14 1 9 4 2
8 9 9 1 13 14 13 4 2
8 9 1 0 13 14 13 4 2
23 15 1 13 4 16 4 4 14 2 11 1 9 1 13 16 4 16 4 1 4 4 14 2
6 9 1 13 16 4 2
30 9 12 12 9 2 9 9 4 1 0 9 1 13 16 2 9 9 2 1 13 4 16 4 4 4 13 16 4 4 2
8 9 9 1 9 14 4 4 2
12 9 1 1 2 9 1 9 1 1 13 4 2
15 15 1 7 2 9 9 1 9 1 13 9 1 13 4 2
11 10 9 1 9 1 1 9 1 1 13 2
12 7 2 9 9 1 13 4 16 1 4 4 2
31 3 2 9 1 1 2 13 16 13 4 9 2 1 9 0 9 2 9 9 1 3 9 1 0 4 13 16 4 16 4 2
25 2 9 4 11 2 1 13 9 1 9 9 2 15 1 13 14 1 0 4 13 4 16 4 4 2
24 2 9 1 13 4 4 16 1 13 16 2 10 9 1 9 1 13 4 16 1 4 4 2 2
14 11 9 1 12 12 9 2 3 0 4 13 4 4 2
16 9 1 13 9 9 1 13 16 1 2 9 1 9 4 4 2
15 9 1 9 1 9 2 9 1 0 9 1 13 4 4 2
10 9 4 9 4 4 1 13 4 4 2
20 3 2 9 9 1 9 1 9 1 3 1 13 14 3 14 1 13 4 4 2
32 9 1 11 9 1 9 9 9 1 13 9 3 2 9 1 9 9 9 9 1 13 4 4 12 12 12 9 1 9 4 4 2
26 9 1 9 1 13 9 1 2 12 12 12 12 9 9 2 13 4 4 9 2 9 9 1 13 4 2
23 10 9 2 9 1 13 4 9 1 9 9 9 1 13 4 4 2 9 9 1 13 4 2
17 13 4 4 9 1 2 9 9 9 9 1 9 1 13 4 4 2
23 9 9 1 9 9 1 9 9 1 13 4 4 2 9 1 1 9 9 1 13 4 4 2
16 10 9 2 9 1 1 9 1 9 1 13 4 16 4 4 2
17 9 9 1 9 9 1 13 4 9 2 3 9 9 1 13 4 2
28 15 1 2 9 9 1 9 1 13 4 9 4 4 16 1 0 2 1 2 9 1 9 1 9 1 13 4 2
17 9 9 7 9 9 2 9 9 1 9 1 13 4 16 4 4 2
11 9 1 9 9 4 9 1 9 13 4 2
17 9 1 2 9 9 9 4 16 9 1 13 4 4 16 14 2 2
14 9 1 2 9 1 9 1 13 4 4 16 14 2 2
25 9 9 1 9 9 1 9 1 9 1 13 2 9 9 1 1 9 1 13 4 1 13 4 4 2
25 7 2 11 9 1 15 1 13 16 1 2 9 9 1 9 1 9 9 4 13 4 16 4 4 2
15 9 9 9 7 2 9 2 9 1 9 1 3 13 14 2
12 7 9 9 2 9 1 9 1 13 16 4 2
26 15 1 1 2 9 1 13 4 16 4 9 9 1 9 1 9 1 13 4 2 1 13 4 16 4 2
23 7 2 2 9 9 1 9 1 13 9 1 9 9 9 2 1 9 9 1 13 16 4 2
11 9 1 9 9 1 1 13 4 16 4 2
30 9 2 9 9 1 13 9 9 2 13 4 4 9 1 9 4 4 2 9 9 1 13 9 4 4 1 13 16 4 2
29 9 1 15 14 0 4 13 4 9 1 1 2 9 1 13 4 4 14 1 1 9 9 1 2 9 1 13 4 2
20 9 2 9 9 1 9 9 9 1 1 12 9 9 1 9 1 13 4 4 2
30 13 4 4 9 7 2 9 1 13 4 9 7 1 2 3 13 9 4 16 4 16 2 13 4 4 4 16 4 4 2
9 7 7 2 9 1 3 1 13 2
24 9 9 9 1 13 4 16 1 2 15 9 1 9 1 9 9 1 9 1 0 4 13 2 2
23 9 9 1 13 4 16 4 14 1 12 12 9 9 1 9 9 2 9 9 9 1 13 2
19 9 9 9 9 9 9 1 9 1 2 0 9 1 13 9 9 1 0 2
35 9 1 9 1 3 4 4 2 9 2 3 9 1 13 9 1 13 4 4 16 2 9 9 2 9 1 9 1 9 9 13 16 1 0 2
13 7 2 9 9 1 9 1 3 0 4 1 4 2
27 9 9 2 9 1 12 12 12 12 12 9 1 9 9 9 9 9 1 9 1 13 4 9 9 1 13 2
45 15 1 1 9 1 9 9 1 13 4 9 2 9 1 13 9 1 13 16 2 13 4 2 9 9 2 9 9 2 13 16 13 2 1 13 16 2 12 12 9 9 1 13 4 2
21 11 9 1 9 1 2 9 9 2 9 1 9 1 9 1 9 1 13 4 4 2
3 3 13 2
5 15 1 0 4 2
