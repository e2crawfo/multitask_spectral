704 17
8 9 8 13 9 1 9 9 9
41 8 12 2 12 2 8 8 2 2 13 9 9 0 7 9 9 9 9 9 8 8 9 9 1 8 9 1 9 9 9 15 13 15 9 9 1 0 0 1 9 2
26 7 13 8 1 9 7 2 9 0 0 7 9 9 9 2 0 2 13 9 1 9 12 1 9 2 2
27 7 13 9 1 0 9 1 9 9 9 1 9 9 2 13 1 9 9 13 15 9 1 9 2 9 0 2
26 7 1 12 9 2 9 13 9 9 8 12 9 9 9 9 1 15 1 1 13 9 0 1 12 9 2
23 7 13 8 2 14 13 1 9 9 15 9 2 2 1 9 1 0 15 14 13 0 9 2
21 2 8 8 2 14 13 2 8 2 1 2 8 2 1 9 12 12 9 2 9 2
58 8 12 2 12 2 8 8 2 2 13 1 9 9 2 8 8 2 7 2 8 8 8 2 1 9 9 9 7 9 0 2 8 8 2 14 13 9 0 2 8 2 1 9 0 0 1 9 9 0 2 8 2 1 9 12 12 9 2
56 7 1 1 9 2 8 8 2 1 9 2 7 14 13 9 9 2 8 2 9 1 9 1 9 9 15 13 7 13 15 9 15 12 12 9 1 9 1 10 9 0 15 14 13 9 9 15 1 9 15 0 0 1 9 0 2
50 7 1 9 9 9 2 14 13 2 8 8 2 1 9 9 2 8 2 1 2 8 2 9 7 9 7 9 1 9 1 9 12 12 9 1 9 9 1 9 0 1 9 9 2 8 8 2 1 9 2
43 7 14 13 9 2 8 2 1 9 10 9 1 15 1 12 1 12 5 1 9 0 15 14 13 1 9 9 2 8 8 2 7 2 8 2 1 1 9 2 8 8 2 2
22 7 1 0 7 13 9 9 2 8 8 2 9 10 9 1 1 2 8 8 8 2 2
9 7 1 0 7 13 1 9 9 2
30 7 13 2 8 2 9 9 0 2 8 2 8 2 7 9 2 8 8 2 0 7 9 0 0 2 8 8 8 2 2
49 7 13 3 9 9 1 2 8 2 7 2 8 2 7 2 8 8 2 7 3 9 0 9 1 9 9 2 8 8 2 7 2 8 2 7 1 9 9 1 9 0 2 8 2 7 2 8 2 2
11 9 0 0 0 1 9 12 12 9 1 9
43 9 12 2 12 2 8 8 2 2 13 9 2 9 2 0 9 9 7 9 0 7 0 13 9 9 0 2 0 2 1 9 12 12 9 1 9 9 0 0 1 9 0 2
38 7 1 1 9 7 14 9 13 9 1 9 9 0 1 9 12 9 7 13 9 9 1 9 8 8 1 9 7 9 1 9 7 9 1 9 7 9 2
38 7 13 2 9 2 7 9 0 8 9 0 1 9 2 0 2 7 9 2 11 8 2 0 8 13 0 1 9 0 1 9 1 9 0 8 8 8 2
29 7 13 9 1 9 9 9 12 9 0 9 9 0 1 9 1 9 12 12 9 7 13 1 9 9 0 1 8 2
34 7 9 0 0 15 8 1 9 15 1 9 8 8 9 9 1 9 0 0 9 1 9 15 8 8 15 13 1 0 1 9 2 9 2
8 9 9 9 0 0 1 9 0
48 9 12 2 12 2 8 8 8 2 2 13 9 0 7 9 0 1 9 1 9 0 0 1 9 2 8 2 9 9 13 9 1 9 1 9 9 1 9 1 9 9 9 13 9 9 1 9 2
41 7 13 8 8 7 11 8 1 9 1 9 12 9 0 1 9 9 15 0 1 8 9 9 13 9 1 9 0 8 8 1 9 9 7 9 9 1 9 9 9 2
23 7 14 13 0 9 0 1 9 9 9 1 9 9 10 9 15 13 1 9 9 1 9 2
29 7 13 7 8 15 8 9 0 0 8 8 8 0 1 9 8 8 7 9 1 9 2 9 9 0 1 9 2 2
44 7 13 8 1 9 9 9 1 9 7 15 9 9 8 8 8 9 0 15 13 1 9 0 2 9 12 1 9 9 13 1 15 9 1 9 9 9 1 9 9 0 13 9 2
54 7 13 8 8 7 15 9 1 9 9 2 9 8 0 15 13 9 0 1 9 7 0 0 2 1 9 9 13 9 9 1 15 7 15 8 2 9 9 0 1 9 1 8 8 8 2 1 1 9 0 1 9 0 2
19 7 13 9 7 8 13 7 9 8 2 1 9 9 2 1 9 9 9 2
32 7 13 2 1 1 9 9 15 7 2 12 1 12 1 9 15 13 9 1 15 0 7 13 9 1 9 1 8 8 8 2 2
20 7 13 8 1 9 2 9 9 0 1 9 2 0 7 2 9 1 9 2 2
37 7 13 9 7 8 8 8 13 9 1 9 8 10 2 9 0 2 1 8 8 1 12 9 2 9 7 1 8 8 2 1 12 9 2 9 2 2
34 7 13 9 7 2 8 13 14 15 13 1 9 1 15 13 1 15 7 7 9 10 9 13 1 9 1 8 7 1 9 10 0 2 2
30 7 13 7 8 8 9 9 0 1 9 2 8 8 8 2 0 9 1 9 9 13 3 1 9 9 8 7 9 15 2
61 7 1 9 8 8 8 8 8 2 13 1 9 9 15 12 9 15 8 8 8 13 9 9 0 1 9 9 8 8 8 8 8 9 1 9 9 9 0 8 8 8 8 8 8 8 8 8 8 8 8 8 2 15 14 13 0 9 1 9 15 2
7 9 1 9 9 0 1 8
46 8 2 8 2 12 2 12 2 8 8 2 2 13 9 7 9 13 9 9 9 1 8 2 9 2 1 1 12 9 1 9 0 13 13 1 9 9 7 1 1 12 9 1 9 0 2
33 7 13 9 7 9 9 0 13 9 0 1 9 7 9 7 9 7 13 9 9 1 9 1 9 8 1 9 9 0 7 9 9 2
8 9 0 0 13 1 9 0 0
57 9 12 2 12 2 8 8 2 2 13 9 0 0 0 9 9 9 7 9 13 7 9 14 13 1 9 1 9 0 1 9 0 9 1 9 12 7 14 13 1 9 15 9 9 0 1 9 13 15 9 1 9 1 9 12 9 2
46 7 13 9 1 9 0 9 9 1 9 15 2 7 9 14 13 1 9 1 9 0 0 9 12 7 14 13 1 9 12 9 1 13 9 0 13 9 15 1 9 0 1 9 9 2 2
36 7 13 9 1 10 9 1 9 9 9 9 9 15 2 1 9 2 9 0 1 9 9 2 9 2 8 12 2 15 13 9 15 1 12 9 2
19 7 13 9 2 14 9 13 1 9 15 9 9 0 1 1 9 8 2 2
46 7 13 9 1 9 1 9 9 7 9 9 9 2 9 2 8 12 2 13 9 0 7 7 15 13 8 8 8 7 12 9 2 9 15 13 1 15 1 9 1 9 0 1 9 2 2
25 7 13 9 7 8 13 1 9 15 1 9 1 8 0 13 8 13 9 15 9 1 9 8 0 2
35 7 13 9 1 7 9 13 2 1 0 9 9 9 2 0 7 2 9 0 1 9 0 0 7 14 3 1 9 0 7 0 13 9 2 2
32 7 13 9 1 9 0 7 2 9 8 14 13 8 1 9 7 7 8 8 14 13 12 8 1 9 8 14 1 10 9 2 2
38 7 13 9 9 9 9 8 8 9 9 7 9 2 14 13 15 13 9 0 2 1 9 9 2 9 2 8 12 2 0 15 13 8 8 1 12 9 2
27 7 13 8 1 9 0 2 7 9 14 13 9 15 1 9 9 0 1 10 9 2 1 1 9 1 9 2
25 7 13 9 0 9 9 7 15 13 2 1 9 2 9 0 1 9 9 2 9 2 8 12 2 2
32 7 13 9 1 9 9 0 1 9 9 7 2 9 0 5 8 12 5 13 1 9 0 1 9 1 9 15 1 9 0 2 2
27 7 13 13 1 9 2 9 12 1 9 0 9 1 10 9 15 13 7 13 9 9 9 7 1 15 9 2
4 9 8 2 9
121 8 12 2 12 2 8 8 8 2 2 1 9 0 1 9 8 0 0 1 9 9 13 9 8 8 1 9 8 8 12 2 12 7 12 2 12 2 7 9 8 8 1 9 8 8 12 2 12 7 12 2 12 2 7 9 8 8 1 9 8 8 12 2 12 7 12 2 12 7 12 2 12 2 7 9 8 8 1 9 8 8 12 2 12 7 12 2 12 7 2 12 2 12 2 2 7 9 8 8 1 0 8 8 8 12 2 12 2 12 2 12 2 7 12 2 8 7 12 2 12 2
178 7 13 0 8 8 1 9 8 8 12 2 12 7 12 2 12 2 7 9 8 8 1 9 8 8 12 2 12 7 12 2 12 2 7 9 8 8 1 9 8 8 12 2 12 7 12 2 12 2 7 9 8 8 1 9 15 8 8 12 2 12 7 12 2 12 7 12 2 12 2 7 0 8 8 1 9 8 8 12 2 12 7 12 2 12 7 12 2 12 2 7 9 8 8 1 9 8 8 12 2 8 7 12 2 12 2 7 0 8 8 1 9 8 8 12 2 12 7 12 2 12 2 7 9 8 8 1 9 8 8 12 2 12 7 12 2 12 2 12 2 12 2 12 2 12 2 7 9 8 8 1 0 8 8 12 2 12 7 12 2 12 2 7 9 8 8 1 9 8 8 12 2 12 7 12 2 8 2
5 9 8 1 8 0
40 8 12 2 12 2 8 8 8 2 2 13 9 9 9 1 9 9 8 8 9 13 1 9 15 1 9 8 0 1 9 0 1 9 12 9 1 12 12 9 2
38 7 13 9 8 8 8 2 8 0 1 9 9 1 9 8 2 14 15 9 0 13 15 9 0 1 9 8 8 0 7 15 8 8 8 9 0 2 2
33 7 13 8 9 0 0 15 13 1 8 2 7 15 13 13 9 1 8 7 9 1 9 0 1 7 13 1 9 1 9 8 8 2
84 7 13 8 2 12 9 2 13 1 8 8 9 9 0 1 9 1 9 0 7 13 1 9 9 15 1 9 0 8 8 2 9 8 8 0 2 7 15 14 13 9 15 0 1 9 9 7 13 9 0 1 9 1 9 9 1 8 2 7 15 13 9 9 9 8 8 1 9 0 7 13 9 15 9 1 9 7 13 1 9 0 1 9 2
30 7 13 8 7 1 9 0 15 13 15 13 8 2 9 9 8 8 1 9 1 8 7 9 15 1 9 1 9 2 2
35 7 13 7 15 13 1 9 0 1 9 15 7 7 9 15 2 8 2 14 13 1 9 0 1 9 0 7 13 9 15 0 1 8 0 2
55 7 13 8 9 0 1 8 7 13 9 15 0 2 8 7 13 1 9 0 7 15 14 13 1 9 9 15 0 1 9 9 8 2 13 15 1 8 8 0 7 15 14 13 9 1 0 7 15 14 13 9 1 9 15 2
39 7 13 8 2 8 1 9 1 8 1 9 9 1 9 1 8 8 0 1 8 8 2 2 0 2 8 8 1 9 1 8 1 9 8 8 1 9 2 2
36 7 13 2 8 0 9 1 9 0 3 1 7 8 1 8 2 2 7 13 2 14 15 9 8 1 15 0 7 8 8 8 13 1 8 2 2
9 9 2 0 2 1 9 0 9 0
45 8 12 2 12 2 8 8 2 2 13 9 0 0 7 9 13 2 0 2 1 9 0 0 1 12 9 2 9 0 7 7 9 9 7 9 13 9 9 0 0 1 9 9 15 2
27 7 13 9 1 9 0 0 8 8 7 2 9 0 1 9 7 7 9 9 1 9 9 1 9 9 2 2
62 1 9 15 2 13 9 9 0 1 8 2 9 8 0 0 1 9 2 1 9 15 0 7 9 9 13 12 1 9 9 1 8 7 13 9 15 2 7 13 7 0 8 1 8 9 2 7 7 9 15 13 1 8 2 7 13 9 2 1 9 0 2
33 7 13 9 0 7 9 13 9 7 9 9 15 1 9 0 1 9 7 7 15 2 13 9 9 1 9 0 15 13 9 9 2 2
52 7 13 9 9 8 2 8 1 9 0 7 9 9 13 9 1 9 9 15 1 9 0 1 9 9 9 2 7 13 7 9 9 2 8 2 13 9 15 1 9 9 9 0 9 1 8 7 9 1 9 0 2
17 7 8 13 7 9 0 0 14 13 9 2 9 0 2 1 9 2
41 7 14 13 0 9 0 1 9 9 15 1 8 2 9 9 0 2 2 7 14 13 9 1 12 9 0 2 9 0 1 9 0 0 1 9 9 0 1 9 0 2
20 7 13 9 0 0 9 12 12 9 1 9 1 15 12 1 12 1 9 9 2
54 7 13 9 9 0 0 8 8 8 7 12 9 9 14 13 1 9 1 15 12 9 0 1 9 9 0 1 9 2 7 13 2 14 9 1 7 9 9 14 13 0 2 2 0 7 9 14 13 2 9 1 9 2 2
46 7 13 9 9 0 0 8 8 7 9 9 13 9 1 9 7 15 14 13 2 9 9 15 9 2 2 0 1 7 12 12 9 3 13 1 9 0 15 13 1 12 9 2 9 0 2
32 7 14 13 10 9 0 9 9 1 9 0 0 7 1 9 9 9 15 14 13 1 9 1 9 9 1 12 9 2 9 0 2
26 7 13 0 1 9 9 7 9 9 9 7 9 9 9 1 9 1 9 9 1 9 0 1 9 0 2
52 7 13 9 9 8 8 8 7 15 13 1 9 0 1 9 9 2 7 9 9 13 1 9 9 0 7 13 8 9 9 0 2 7 15 14 13 1 9 1 15 7 13 15 9 7 13 15 1 9 9 0 2
6 9 8 1 9 2 9
46 8 12 2 12 2 8 8 8 2 2 13 9 9 1 8 9 9 9 8 0 1 9 9 1 9 2 1 12 9 2 15 13 15 8 1 12 1 12 9 2 9 0 1 9 8 2
43 7 13 9 12 0 1 9 13 8 8 7 9 7 9 8 8 8 2 7 0 2 15 13 1 15 9 2 9 9 2 2 8 7 9 7 9 0 9 7 9 8 8 2
9 9 0 13 1 12 9 0 2 9
51 9 12 2 12 2 8 8 8 2 2 13 9 0 1 9 9 1 9 12 2 12 1 12 9 0 2 9 0 1 9 12 9 15 8 8 8 8 8 8 8 8 8 8 8 8 8 8 8 8 8 2
20 7 13 9 9 1 12 9 0 2 9 1 1 14 13 1 1 9 9 9 2
42 7 13 9 0 1 9 9 0 15 13 1 9 9 7 13 1 12 9 2 9 0 2 13 15 9 9 8 0 1 0 1 9 0 2 9 7 13 1 12 1 15 2
64 1 15 2 14 13 9 9 1 9 9 8 15 13 15 9 1 12 1 12 9 0 2 9 2 7 13 9 0 0 1 9 9 12 1 9 0 0 7 15 14 13 9 1 12 1 12 9 2 9 0 1 8 8 7 9 1 12 1 12 1 15 1 9 2
11 8 8 0 1 9 9 9 1 9 7 9
42 9 12 2 12 2 8 8 2 2 13 9 9 9 0 1 9 9 0 8 8 9 9 1 8 1 9 15 1 9 9 1 9 1 9 7 9 1 2 9 2 0 2
38 7 13 8 8 13 9 15 9 9 8 0 1 9 9 1 9 9 8 8 8 2 8 0 1 9 1 9 9 2 1 9 0 2 7 9 0 2 2
17 7 13 9 0 2 13 9 9 1 9 7 9 1 9 0 2 2
43 7 13 8 9 1 9 15 1 9 0 9 9 9 8 8 2 7 13 1 9 0 7 13 9 9 0 1 9 8 8 1 9 7 9 15 13 1 9 9 1 9 9 2
13 7 13 8 8 1 9 15 1 8 0 1 9 2
30 7 13 8 1 9 8 8 9 0 8 8 7 9 9 0 1 9 8 11 8 1 9 9 0 1 9 9 9 9 2
11 9 13 1 9 9 8 2 8 2 1 9
51 9 12 2 12 2 8 8 2 2 13 9 9 0 0 7 9 13 9 9 1 9 9 9 8 0 15 8 1 9 0 2 1 9 9 2 1 9 0 2 1 9 9 9 8 1 0 15 0 1 9 2
22 7 13 9 1 9 0 9 15 7 9 8 1 9 13 9 9 1 0 1 9 0 2
54 7 13 8 7 9 1 9 0 2 9 12 9 13 9 1 9 15 1 9 9 7 8 12 12 8 1 9 2 7 13 12 5 1 9 9 1 8 1 9 2 7 1 9 10 9 13 9 8 0 12 9 1 9 2
29 7 13 9 8 8 1 8 8 0 7 0 0 9 0 1 9 9 1 9 9 9 1 9 9 7 9 15 0 2
31 7 1 9 0 13 9 1 9 8 1 9 9 9 0 7 9 1 10 9 7 14 3 1 9 1 9 0 1 9 9 2
12 9 9 8 0 1 9 1 8 1 9 9 8
44 8 12 2 12 2 8 8 2 2 13 9 1 9 9 9 0 1 8 7 9 9 8 8 14 13 1 9 1 9 9 9 0 1 8 2 8 2 1 8 1 9 8 8 2
36 7 13 9 1 9 1 9 8 8 7 2 9 14 13 1 1 9 9 0 9 9 0 1 9 15 14 13 1 15 1 10 1 15 8 2 2
36 7 1 1 9 2 7 14 9 0 1 9 1 9 13 9 0 2 7 13 9 1 9 7 2 9 9 0 1 9 9 0 1 8 8 2 2
69 7 1 9 15 13 15 9 8 8 0 0 1 12 9 2 9 0 0 8 8 8 2 12 9 2 8 13 9 7 8 8 2 12 9 2 8 13 9 0 1 9 0 1 9 9 2 7 15 9 1 9 9 0 15 13 1 9 8 0 1 12 9 2 9 1 9 9 0 2
11 9 9 0 9 0 1 9 0 1 9 0
58 8 12 2 12 2 8 8 2 2 13 9 1 0 1 9 2 9 1 9 9 1 8 2 9 8 0 2 0 1 9 0 9 0 13 1 9 14 1 0 1 9 0 1 9 0 2 7 13 9 9 1 9 8 11 8 9 9 2
35 7 13 9 1 9 7 9 14 13 1 9 12 9 7 14 13 9 9 0 1 9 0 7 3 1 9 2 9 2 0 9 1 9 9 2
31 7 13 9 8 7 9 2 14 13 1 9 8 7 9 9 9 9 14 13 1 9 1 9 9 9 0 1 8 8 2 2
44 7 14 13 9 9 15 13 1 15 9 2 8 2 2 8 8 8 8 2 1 9 12 9 2 9 1 9 9 8 2 8 15 13 0 1 8 8 1 8 2 9 0 2 2
35 7 14 13 9 15 13 1 15 9 0 2 9 12 1 9 7 14 13 1 9 9 1 9 1 8 7 8 7 9 0 7 8 7 8 2
12 11 8 13 1 9 1 9 0 7 0 1 9
47 9 12 2 12 2 8 8 2 2 13 9 9 0 1 9 8 11 8 9 9 1 9 15 1 9 1 9 9 0 1 9 1 9 9 2 9 7 9 9 2 9 13 1 9 9 0 2
55 7 13 11 8 1 9 0 1 9 9 2 7 15 13 1 9 2 1 9 0 1 9 0 1 9 9 9 2 9 7 9 9 2 9 1 9 15 13 9 1 15 1 8 8 2 7 15 14 13 1 9 9 0 2 2
50 7 13 11 8 7 2 9 0 1 9 9 0 1 9 1 9 13 1 15 9 9 9 0 1 9 9 0 15 13 1 15 8 2 9 0 2 7 9 2 2 1 9 1 9 9 9 9 9 0 2
50 7 13 11 8 7 2 1 9 9 1 9 9 1 12 9 5 9 1 9 9 8 8 2 9 5 9 12 2 2 8 8 8 14 8 8 1 15 7 15 14 13 1 9 0 8 9 9 0 2 2
41 7 13 8 1 9 9 8 8 1 12 9 5 9 1 9 13 15 1 0 1 12 9 2 7 14 13 1 9 1 9 0 1 9 9 0 1 0 8 9 0 2
51 7 1 1 11 8 2 7 14 9 7 9 14 13 1 8 8 1 9 1 9 9 9 0 0 7 9 9 0 7 9 7 9 1 9 0 1 9 9 9 15 13 1 9 9 0 0 1 9 1 9 2
50 7 13 7 9 13 13 1 7 2 13 12 9 0 1 9 0 1 9 15 7 7 13 10 9 1 9 0 1 9 0 7 9 8 8 8 8 8 2 2 1 1 7 13 9 9 9 9 9 0 2
31 7 13 11 8 1 9 0 7 9 13 2 7 15 14 13 7 13 1 9 15 1 9 8 2 1 9 7 13 9 0 2
41 7 13 9 7 9 9 15 13 9 9 15 1 9 1 12 5 1 9 1 9 0 2 14 13 9 9 8 7 8 8 7 9 0 1 9 1 9 9 0 2 2
34 7 14 13 11 8 14 1 9 9 9 7 14 1 9 0 15 13 1 15 9 1 9 7 9 9 2 9 9 0 1 0 7 9 2
29 7 13 7 9 15 9 7 9 0 1 9 0 1 9 0 13 1 12 1 9 0 2 14 13 2 9 0 2 2
33 7 0 2 13 11 8 1 9 1 7 14 13 9 9 9 0 1 9 9 0 1 12 9 5 9 1 9 2 9 1 9 2 2
11 9 9 0 2 9 9 1 9 12 2 12
62 9 12 2 12 2 8 8 8 2 2 13 9 9 0 1 9 12 2 12 2 9 12 2 12 7 12 2 12 7 12 2 12 7 12 2 12 7 12 2 12 2 7 13 1 9 0 1 9 0 0 1 9 0 15 13 15 9 7 13 9 9 2
21 7 13 9 9 15 1 12 9 13 15 9 12 9 7 9 7 1 15 12 9 2
40 7 1 9 0 2 13 9 9 15 0 7 13 1 9 9 9 12 2 12 2 12 2 12 7 12 2 12 7 12 2 12 7 12 2 12 7 12 2 12 2
28 7 13 9 9 1 9 2 7 1 9 9 0 14 13 9 2 1 1 13 9 9 1 9 0 1 9 0 2
10 0 13 9 12 0 9 1 9 1 9
53 8 2 8 2 12 2 12 2 8 8 2 2 13 0 9 2 1 9 13 15 9 0 1 9 8 8 7 13 9 8 8 9 1 15 9 9 2 7 15 2 13 9 9 2 1 12 0 9 1 9 9 0 2
44 7 13 9 7 2 12 12 9 13 1 9 9 8 2 15 13 15 8 2 13 1 9 2 1 15 12 1 0 9 2 2 9 1 9 13 15 9 8 1 9 9 1 8 2
17 7 13 9 7 2 10 9 13 15 9 0 0 7 9 0 2 2
45 7 14 13 9 1 0 9 1 8 1 9 8 2 7 13 9 9 9 0 1 9 7 12 1 15 13 1 9 9 1 9 9 0 7 13 9 1 9 7 13 9 1 9 15 2
55 1 9 0 2 13 9 9 1 9 0 9 9 1 9 1 9 9 1 9 8 13 9 2 7 13 7 2 10 9 14 13 9 1 9 15 1 9 0 2 7 14 13 9 0 1 9 1 9 15 7 13 9 15 2 2
10 9 9 8 0 14 13 9 0 1 9
54 8 12 2 12 2 8 8 2 2 13 8 8 15 13 9 1 9 8 1 9 12 7 12 7 15 14 13 1 9 0 2 9 9 1 9 9 0 14 13 2 0 7 0 2 7 4 0 1 9 7 13 9 0 2
37 7 13 8 15 13 9 3 1 9 8 1 9 2 7 9 13 1 15 1 0 1 9 7 14 3 1 9 15 13 9 15 1 9 9 1 12 2
29 7 13 8 1 9 15 7 13 8 1 9 0 14 13 15 1 15 0 2 7 15 13 9 15 1 9 1 9 2
35 7 1 9 13 9 9 13 8 7 9 15 14 13 8 9 15 13 1 9 9 1 12 9 2 9 12 1 8 1 9 9 15 8 8 2
38 7 13 9 2 1 9 15 8 1 9 15 14 8 1 15 15 13 1 15 7 9 15 9 0 7 9 15 13 1 15 13 1 9 1 9 15 2 2
24 7 13 1 7 2 9 9 0 7 0 7 13 1 9 8 0 8 8 13 1 9 15 2 2
28 7 10 9 14 13 1 0 9 8 7 9 8 0 15 14 13 9 3 9 13 1 15 1 9 15 9 9 2
33 7 13 8 7 15 13 9 15 13 9 1 8 1 9 9 9 9 15 0 2 8 1 9 7 15 14 13 2 7 14 13 9 2
8 8 2 9 0 0 13 12 9
36 8 2 9 9 2 2 13 9 0 8 8 9 0 0 13 1 9 15 9 9 0 7 9 1 9 15 1 1 13 8 8 8 9 1 9 2
36 7 13 9 7 8 8 8 9 9 9 9 9 7 0 9 13 9 9 9 9 8 8 8 7 13 9 8 8 9 9 9 0 9 9 0 2
17 7 13 9 9 0 7 9 13 12 9 1 15 9 0 7 9 2
20 7 13 8 8 8 13 9 1 9 9 0 9 1 0 9 1 9 8 8 2
17 7 13 8 1 15 9 9 9 7 9 1 9 0 0 1 9 2
7 7 1 15 13 9 9 0
9 9 9 9 8 8 2 9 1 9
8 9 9 8 8 2 9 1 9
9 9 9 8 8 8 2 9 1 9
8 9 9 8 8 2 9 1 0
11 9 9 8 8 8 2 9 1 9 7 9
9 9 9 8 8 8 2 9 1 9
7 9 8 8 2 9 1 9
12 9 9 8 8 8 2 9 1 9 0 7 9
38 7 13 9 15 13 1 0 1 9 1 9 9 8 1 2 9 2 1 9 9 2 9 9 9 7 9 7 9 7 9 7 9 0 7 9 7 9 2
29 7 13 9 1 9 13 1 15 9 1 9 0 0 1 8 7 1 9 0 7 0 1 9 15 1 9 7 9 2
7 1 9 9 1 9 9 9
9 8 7 8 13 9 9 0 1 9
59 8 2 9 9 2 2 13 9 8 8 3 7 9 9 0 8 8 13 1 0 0 9 9 9 0 1 9 1 9 9 1 9 15 1 9 9 9 2 7 13 9 1 9 0 7 0 9 15 7 9 0 1 9 14 13 9 9 0 2
42 7 1 9 0 13 8 7 8 7 8 1 9 1 9 13 9 1 9 15 1 9 9 9 0 7 15 9 14 13 1 9 9 1 9 9 9 7 1 9 9 0 2
86 7 14 13 9 1 0 9 1 9 9 7 15 14 13 9 9 7 13 1 9 0 9 9 0 1 15 2 7 13 9 1 8 8 7 9 8 14 13 9 9 0 9 14 7 15 14 13 9 0 12 1 9 15 1 9 9 1 9 13 7 13 15 8 1 9 0 9 0 1 9 9 7 1 0 9 9 0 1 9 1 9 0 1 10 9 2
71 7 13 9 0 7 9 0 9 0 1 9 9 9 1 9 1 15 7 10 9 14 13 9 0 14 13 9 0 0 9 1 8 8 2 9 1 15 14 13 1 9 9 0 1 15 13 9 7 13 9 0 1 9 0 8 8 14 13 9 8 8 1 9 9 1 9 0 1 9 0 2
77 7 13 8 14 15 7 13 9 1 9 0 7 14 13 9 13 9 9 0 1 9 0 9 1 9 0 7 14 13 1 9 9 9 7 13 9 2 7 13 9 7 9 0 9 15 14 13 1 9 9 9 1 9 0 15 13 9 15 1 8 7 14 13 9 15 13 9 1 9 9 9 1 9 15 0 0 2
9 9 1 9 0 1 9 0 1 9
44 1 9 0 13 9 0 0 3 7 9 0 1 9 0 1 9 0 13 1 9 1 9 9 1 9 15 14 13 15 9 0 1 9 8 8 1 12 9 1 9 9 1 9 2
16 7 13 9 12 9 7 13 15 9 9 0 1 9 8 8 2
15 7 14 13 9 9 1 9 1 7 13 1 15 1 9 2
9 9 11 8 13 9 1 9 9 0
30 8 2 8 2 13 9 9 7 9 9 15 1 9 0 9 9 9 8 8 11 8 9 3 1 9 8 8 9 0 2
26 7 13 9 9 1 10 9 9 1 9 13 1 9 9 0 1 9 9 0 0 1 9 7 9 0 2
39 7 13 10 9 15 13 9 9 0 13 9 9 0 1 9 9 0 7 9 15 1 9 13 7 9 0 8 1 9 9 0 1 9 9 0 1 9 0 2
48 7 13 9 9 15 13 15 1 9 1 9 9 9 7 9 0 1 10 9 1 15 13 1 9 9 0 13 1 15 9 0 9 1 9 7 9 7 9 8 8 1 15 9 9 7 9 0 2
55 7 1 9 0 13 9 9 9 1 9 9 1 9 0 1 10 9 1 9 9 9 0 0 1 9 9 9 7 9 9 8 0 14 3 1 9 9 0 1 9 9 0 7 9 9 0 1 9 0 7 9 15 9 0 2
73 7 13 9 9 15 13 15 1 9 0 1 9 9 1 9 9 9 1 9 1 0 9 7 9 9 8 1 9 1 0 9 0 7 1 9 9 7 9 7 9 9 0 9 1 9 8 7 9 9 1 9 8 8 1 9 9 1 9 9 9 0 7 9 1 9 15 13 9 15 1 10 9 2
25 7 13 9 9 1 9 9 15 9 9 9 9 9 0 1 9 9 9 9 7 9 1 9 0 2
4 1 9 8 2
9 14 13 9 0 7 0 1 9 2
37 9 2 9 9 2 2 13 9 3 7 9 9 9 0 8 8 15 13 1 1 8 1 9 9 9 0 14 13 1 9 9 0 7 0 1 9 2
27 7 13 9 8 7 9 9 0 9 1 9 0 1 9 9 9 9 8 8 0 9 1 9 9 1 9 2
25 7 13 9 0 1 9 7 9 8 9 13 9 1 9 1 9 7 13 7 13 9 0 9 0 2
34 7 13 0 0 13 1 9 9 0 0 1 9 8 8 7 2 9 8 1 9 0 15 15 13 9 0 1 9 0 1 9 9 2 2
34 7 13 7 2 9 13 1 9 10 14 13 8 0 1 9 15 1 9 9 0 9 2 9 1 15 9 13 9 0 0 1 9 0 2
55 7 13 10 0 2 9 1 9 8 14 13 0 9 0 1 9 9 0 9 9 2 0 1 15 1 9 15 13 1 15 9 9 0 1 9 0 1 8 7 9 0 0 15 13 9 15 9 0 1 9 1 9 9 15 2
19 7 13 9 1 9 9 0 13 12 12 9 7 13 8 9 9 0 0 2
46 7 13 9 8 7 13 9 7 9 0 9 1 15 8 8 9 9 9 1 9 9 9 0 13 1 9 9 9 7 13 9 0 2 1 9 9 2 1 9 9 1 9 9 9 12 2
51 7 13 9 0 1 9 0 8 8 13 1 9 13 1 0 1 9 7 9 14 13 9 9 12 15 13 15 9 1 0 1 9 7 13 1 9 1 12 12 9 0 0 1 9 7 9 9 9 1 9 2
40 9 1 15 13 9 7 9 0 8 8 9 9 9 9 15 0 15 13 12 9 9 1 10 9 0 7 9 9 9 8 1 9 9 9 8 1 0 1 9 2
40 7 13 9 15 13 0 9 7 9 0 7 0 13 9 15 1 8 13 1 7 13 9 9 0 1 9 15 0 1 8 9 0 13 1 9 9 8 12 9 2
20 7 13 12 9 1 15 9 1 9 8 1 9 12 13 9 9 1 9 0 2
15 7 13 12 9 7 13 1 9 7 13 9 1 9 0 2
24 7 14 13 8 9 1 2 9 9 0 2 1 9 9 8 8 8 13 9 9 12 15 13 2
6 9 9 9 1 9 0
2 8 8
33 13 9 1 9 0 1 9 9 9 0 9 9 8 9 1 9 1 9 0 0 1 9 9 15 1 9 1 9 9 1 9 9 2
99 7 13 9 12 9 1 15 9 8 8 2 12 9 2 15 13 1 2 9 2 7 9 14 13 9 1 9 0 2 8 8 2 7 15 9 1 12 8 0 14 13 9 15 1 9 1 9 13 1 12 9 7 12 9 2 7 13 7 9 0 14 13 1 9 8 9 1 9 9 13 0 7 9 1 9 7 9 1 1 9 0 2 0 1 7 10 9 12 13 1 9 9 0 7 9 0 1 9 2
64 7 13 7 9 9 15 9 0 1 9 9 0 1 9 9 7 13 9 0 1 9 9 1 10 9 2 7 13 9 9 15 14 13 1 12 12 9 1 9 2 7 1 9 15 14 13 9 9 0 7 9 0 7 9 0 2 9 1 9 0 1 9 2 2
28 9 0 13 9 12 9 1 9 9 2 9 2 8 8 2 0 0 1 9 9 1 9 9 7 9 15 1 9
2 8 8
37 13 9 0 13 1 9 9 9 9 0 1 9 0 2 7 13 7 9 15 1 9 0 13 1 9 9 7 0 0 15 13 15 9 1 9 0 2
62 7 13 9 9 0 1 9 2 8 8 2 8 8 1 2 9 2 7 9 15 13 9 9 9 9 1 8 8 1 9 0 2 1 9 9 9 8 0 1 9 9 0 1 9 9 7 9 9 0 1 15 7 15 14 13 9 0 1 12 12 9 2
90 7 13 2 8 8 2 2 15 13 1 8 9 1 15 2 9 9 12 0 1 9 1 9 9 2 7 15 13 2 7 13 1 9 2 12 9 1 9 7 8 7 9 9 0 7 9 13 0 9 15 1 12 12 9 1 9 7 12 12 9 0 1 9 9 0 2 1 9 1 12 9 13 0 12 12 9 9 1 12 9 9 7 9 2 12 1 15 1 9 2
58 7 13 9 9 0 1 9 9 1 9 9 0 1 9 12 1 12 7 13 1 12 12 9 9 12 1 12 12 9 9 0 2 7 13 9 15 0 1 9 9 15 1 9 13 12 1 12 0 2 1 12 12 9 1 12 12 9 2
76 7 13 8 2 8 13 1 9 0 1 9 8 15 13 9 0 9 12 2 2 8 1 9 9 8 1 9 8 8 0 7 9 7 9 2 7 13 9 9 9 9 0 1 9 9 0 9 9 0 2 7 13 9 9 15 8 1 15 1 10 9 1 9 9 8 8 1 9 0 13 1 9 9 0 2 2
170 7 13 9 9 15 13 1 15 2 8 8 2 9 12 1 12 1 9 2 8 2 0 2 7 12 1 12 1 9 2 8 2 0 2 7 9 9 0 13 12 1 12 1 9 2 8 2 0 13 15 2 8 8 2 1 2 8 2 0 8 13 0 0 9 1 9 1 9 9 2 7 9 9 2 8 2 0 0 1 9 1 9 14 13 12 12 9 2 2 7 15 9 0 9 7 14 13 12 9 9 8 0 2 2 7 13 2 2 8 8 2 1 9 1 9 2 1 9 2 1 2 8 2 0 2 8 13 0 9 1 9 9 1 9 2 7 13 9 8 8 1 12 1 12 1 9 0 13 1 9 0 12 1 12 1 2 9 8 8 1 9 2 1 9 9 15 12 12 9 2
53 7 13 9 1 2 8 8 2 8 13 1 12 12 9 1 9 1 9 13 15 1 9 9 9 1 9 8 8 8 2 9 1 9 8 8 0 1 2 9 8 8 1 9 2 7 15 13 1 12 8 9 0 2
70 7 13 8 2 2 9 8 8 13 12 12 9 1 9 0 2 7 13 9 15 9 12 7 13 9 8 9 0 15 13 1 15 9 9 1 9 9 2 7 13 1 9 15 9 7 15 1 9 1 9 7 8 1 15 1 9 9 13 1 9 8 8 12 1 12 1 9 0 2 2
34 7 13 2 2 9 8 8 0 7 0 8 8 0 8 8 8 1 10 9 1 9 0 7 1 15 0 1 9 0 1 9 9 2 2
131 7 13 7 9 0 0 1 9 7 13 2 2 9 0 1 9 13 1 9 0 2 7 9 9 9 0 1 9 1 9 0 14 13 1 9 15 1 9 0 7 9 9 0 1 1 9 0 2 7 3 0 15 13 9 1 15 1 9 7 1 0 14 13 9 9 0 1 9 9 2 2 7 13 9 9 9 9 1 9 1 12 12 9 2 7 13 9 13 9 0 1 9 0 14 7 9 9 1 9 9 0 13 1 9 0 1 9 2 1 9 13 1 15 9 9 7 9 9 0 1 9 9 9 1 9 9 9 1 9 0 2
88 7 13 8 2 2 9 9 13 7 3 9 1 9 1 10 14 13 1 9 0 14 9 1 9 15 1 15 2 7 7 0 9 9 0 1 9 13 9 8 9 0 1 9 7 9 15 1 9 1 9 9 9 9 2 8 8 13 7 3 9 1 9 9 1 9 8 7 3 1 9 9 9 0 7 0 2 7 1 0 14 13 9 1 9 9 0 2 2
40 7 13 2 2 13 9 1 9 1 9 7 14 13 1 9 9 9 15 9 1 9 0 1 9 2 7 15 9 15 13 9 0 1 9 9 1 9 9 2 2
187 7 13 2 2 7 8 1 9 14 13 3 0 1 9 0 1 9 2 7 13 9 13 8 2 7 1 0 9 7 13 1 9 14 13 1 15 0 1 9 15 1 9 2 2 7 13 8 2 2 3 7 13 9 1 9 9 1 9 15 14 13 9 0 2 14 7 9 13 9 0 1 9 2 2 7 13 9 9 9 8 8 12 9 2 7 13 8 2 2 13 9 9 0 1 9 12 12 9 2 1 12 12 9 2 2 8 8 9 9 1 12 12 9 9 12 2 8 8 8 0 1 9 9 7 9 9 2 7 8 8 8 1 9 1 9 9 9 1 8 8 8 2 2 7 13 2 2 8 8 0 1 12 9 1 9 1 9 2 14 7 9 13 1 9 7 3 9 9 1 12 9 1 12 9 2 7 8 1 15 9 0 1 0 1 9 2 2
70 7 13 1 7 9 15 13 1 9 1 9 0 7 9 9 1 15 2 7 13 7 9 0 1 9 8 8 8 9 15 1 9 2 7 13 2 2 9 0 13 9 9 1 12 1 9 9 9 2 7 15 9 1 9 9 9 1 9 2 7 13 7 8 15 14 13 1 9 2 2
39 7 13 7 9 9 15 1 9 0 0 2 7 13 2 2 8 8 0 1 9 1 1 2 14 7 9 13 1 9 9 0 14 7 13 1 9 9 2 2
60 7 13 2 8 8 2 9 0 1 9 9 1 9 1 9 2 8 2 2 14 7 15 13 15 9 7 13 9 15 1 9 1 9 2 7 13 9 1 9 0 1 13 2 8 2 0 2 8 2 7 13 15 1 9 15 0 1 9 9 2
11 13 1 9 0 7 13 1 9 15 1 8
36 8 2 8 2 13 8 8 8 8 9 8 2 7 13 15 8 8 7 13 8 8 0 2 7 13 8 1 9 15 1 8 1 9 12 8 2
155 7 13 9 1 9 8 8 0 1 8 8 8 2 7 15 9 1 9 8 2 9 15 1 9 9 7 15 13 8 8 0 7 15 13 1 9 15 0 1 8 8 1 9 8 2 7 7 14 13 1 9 15 9 1 9 9 0 2 7 13 8 8 2 12 9 2 8 8 9 2 8 2 2 2 8 9 9 8 1 9 13 7 8 8 7 14 8 8 8 8 14 1 8 8 8 8 8 2 2 7 13 9 15 15 13 9 1 9 1 8 1 15 13 8 1 9 15 2 7 13 8 8 0 0 1 9 0 1 9 1 9 0 1 15 9 15 2 7 13 8 8 2 7 13 8 8 1 9 1 12 9 1 8 9 2
55 7 15 13 9 0 15 13 1 15 9 13 9 1 9 1 9 13 1 15 12 9 7 13 9 2 7 1 9 2 9 2 13 9 1 9 9 1 9 15 1 9 2 1 15 13 1 15 9 2 1 9 1 9 0 2
6 9 0 1 8 7 8
3 8 8 9
38 9 0 1 9 0 9 9 9 0 9 1 9 0 2 14 13 0 9 15 14 13 15 9 0 8 8 1 9 15 0 8 8 1 8 9 9 0 2
24 7 14 13 8 9 8 1 9 9 7 9 9 0 2 7 13 9 1 9 9 9 8 0 2
65 0 15 9 0 15 13 9 15 1 9 15 2 9 1 9 9 2 9 15 13 7 15 14 13 1 9 0 9 15 13 1 9 9 15 8 8 7 9 9 15 8 8 2 7 13 7 9 0 13 15 15 9 0 1 9 9 1 9 7 9 2 1 9 8 2
54 7 8 9 13 9 1 9 15 8 8 8 8 2 8 1 9 0 2 15 13 9 15 2 7 9 1 9 15 0 1 9 2 3 1 9 1 9 9 15 8 8 15 13 9 15 13 9 1 9 1 9 9 0 2
38 7 8 13 1 9 9 0 1 9 15 1 7 15 13 1 9 15 9 1 10 9 2 7 15 1 15 13 8 8 1 9 0 8 8 8 1 9 2
51 9 9 0 8 1 10 9 0 7 1 9 15 9 0 0 2 15 13 0 2 7 8 8 9 8 8 9 8 8 7 1 9 9 9 15 1 9 0 2 1 9 15 1 9 0 8 8 8 1 15 2
35 7 9 0 14 13 8 9 8 1 9 9 1 9 9 2 7 9 0 1 9 7 9 0 1 10 9 0 2 7 13 9 15 1 9 2
56 7 9 0 1 9 9 0 13 15 9 9 9 8 8 8 15 13 9 7 9 0 1 12 9 2 9 2 0 2 1 9 9 9 0 7 0 1 7 9 1 9 1 0 9 2 9 15 0 1 9 9 7 9 9 9 2
24 7 13 9 0 9 9 9 7 9 15 2 7 13 9 9 0 7 9 9 0 1 9 9 2
30 7 9 15 7 13 9 0 7 9 15 9 0 2 7 15 13 15 0 1 9 0 2 1 9 9 9 15 1 9 2
5 2 9 1 8 2
105 9 15 13 15 9 0 1 9 1 9 0 7 15 13 15 1 8 8 8 2 13 1 9 9 0 1 0 8 8 2 13 3 9 9 0 7 0 0 2 7 13 9 2 8 8 8 2 9 1 9 2 9 1 8 2 2 7 13 9 9 2 8 8 2 1 9 8 2 7 15 9 0 1 9 15 13 8 9 2 1 9 1 1 9 1 9 2 1 9 1 9 9 9 0 2 9 15 1 9 2 9 9 8 2 2
46 14 9 9 2 8 8 2 7 13 9 1 9 0 1 9 2 9 13 9 9 0 8 8 13 9 1 8 2 2 13 15 8 8 9 9 13 9 1 9 7 13 9 9 8 8 2
47 7 13 8 3 1 9 9 0 0 2 7 13 9 2 8 2 1 2 8 0 2 1 9 2 9 0 13 1 9 1 12 9 1 0 2 2 7 13 9 1 9 9 0 7 15 13 2
62 14 9 2 8 2 7 13 9 15 9 0 2 2 9 0 1 9 9 2 2 7 3 9 2 8 8 2 13 9 15 1 9 8 8 0 8 8 0 1 9 2 9 0 8 1 9 0 2 8 8 9 2 0 2 13 1 9 9 9 1 8 2
32 7 1 8 2 13 9 0 8 8 1 8 1 9 2 7 13 9 2 8 8 2 1 9 2 12 9 1 9 9 0 2 2
13 9 2 8 9 0 8 8 8 13 9 9 9 9
3 9 8 8
45 13 9 2 8 1 9 2 7 9 15 8 0 15 13 1 9 12 12 9 2 12 12 9 2 13 1 9 1 9 9 9 0 0 1 9 7 9 9 13 1 9 1 9 0 2
104 7 13 9 9 2 8 2 1 9 0 0 1 2 8 1 9 2 8 8 1 2 9 2 7 9 9 9 9 0 2 0 1 9 8 8 0 9 0 8 13 15 9 0 1 9 15 1 9 9 1 9 1 8 8 2 2 7 13 7 9 15 13 1 9 9 1 12 8 8 1 1 15 12 9 0 1 8 8 2 7 1 9 9 13 8 8 1 9 1 15 13 8 8 1 9 1 8 8 1 9 0 1 9 2
67 7 1 9 15 13 9 15 0 9 9 9 9 1 9 0 1 9 7 9 1 9 0 7 9 0 0 2 1 9 13 9 9 0 9 9 9 15 9 1 9 1 9 9 0 1 9 9 15 2 7 13 9 1 9 9 0 7 9 0 1 9 9 13 9 15 0 2
50 7 13 8 7 9 0 1 9 14 13 1 9 1 9 9 9 7 9 9 9 8 2 1 9 7 9 8 1 9 9 9 0 0 2 7 13 9 9 0 1 9 1 9 0 1 12 12 9 0 2
57 7 13 2 8 2 7 8 9 0 8 8 8 8 8 8 13 8 8 8 8 14 9 1 15 13 9 1 9 9 1 9 2 7 13 9 9 9 0 9 8 8 1 9 8 1 9 9 0 0 1 9 7 9 1 9 15 2
95 7 13 8 7 9 8 9 0 1 9 13 12 12 9 9 0 2 7 9 9 9 9 0 8 8 1 9 9 8 8 13 9 9 1 8 9 0 1 12 1 12 2 2 7 9 1 8 8 8 9 9 0 1 10 9 1 9 9 0 2 13 9 9 9 1 9 0 8 9 0 1 9 15 8 8 1 9 9 9 9 0 15 8 8 7 9 9 9 15 13 1 9 9 2 2
32 7 13 9 8 9 0 1 9 8 8 12 1 9 12 12 9 2 12 12 9 2 1 12 9 12 1 9 9 12 1 12 2
19 9 1 9 0 1 9 8 8 8 2 9 0 2 0 1 9 9 0 2
2 8 8
84 13 2 9 0 1 9 0 2 1 9 7 8 9 0 1 9 8 8 13 1 9 1 9 15 1 8 12 1 9 9 9 0 2 7 13 9 0 1 9 0 1 2 9 2 7 8 8 8 13 1 9 1 2 9 9 0 2 1 9 9 2 7 13 9 15 2 7 13 7 9 0 13 9 1 9 0 1 9 9 8 1 9 8 2
38 7 13 1 7 9 13 9 1 9 9 9 15 13 9 15 7 13 9 0 7 9 2 9 9 7 9 8 8 8 0 9 0 1 0 9 13 2 2
137 7 1 9 0 13 15 2 9 2 1 8 3 13 9 9 0 1 9 0 0 8 8 7 2 9 9 15 13 1 15 8 8 8 15 9 9 0 1 9 9 7 9 15 7 9 9 0 1 0 2 7 9 9 0 7 0 1 9 0 1 9 9 0 1 8 2 2 7 13 1 7 8 14 13 2 9 9 0 2 15 13 15 8 7 8 1 9 9 0 2 7 13 2 2 9 9 8 8 8 8 7 15 13 9 0 1 9 2 7 13 7 8 14 13 9 0 2 7 15 0 1 9 0 15 13 13 15 1 9 15 7 14 13 9 0 2 2
33 7 13 7 2 9 10 9 15 9 1 9 0 2 0 7 9 13 15 2 0 7 13 9 0 7 1 15 9 0 7 0 2 2
114 7 1 9 9 0 2 0 13 9 9 0 1 9 0 15 13 15 8 8 7 15 2 13 9 9 9 0 1 9 2 7 13 9 15 1 9 9 8 2 8 2 7 15 13 1 0 0 2 0 2 0 1 1 9 9 2 8 8 13 15 9 1 12 1 9 9 2 9 8 2 7 0 13 15 9 2 9 2 1 9 2 9 9 8 2 7 1 9 9 9 13 9 0 2 2 7 13 7 9 0 2 13 0 9 7 9 1 9 0 1 9 9 2 2
54 7 13 1 7 9 9 2 14 13 10 9 1 9 15 2 7 9 9 9 7 9 2 8 8 9 8 8 8 8 2 2 7 13 9 1 9 13 1 9 1 9 0 0 1 9 9 9 1 9 0 1 9 0 2
5 2 9 9 2 8
92 1 15 2 13 9 9 2 9 0 2 2 1 9 8 8 8 2 1 8 9 8 8 1 2 9 2 7 8 13 1 12 9 0 2 9 2 0 1 2 9 0 1 9 15 13 15 12 1 9 9 9 0 8 9 8 8 8 7 9 8 8 2 2 7 13 8 8 13 7 13 1 9 0 2 0 8 8 13 7 13 1 9 9 15 15 13 13 15 1 9 15 2
19 9 13 1 0 1 9 9 9 7 9 2 9 13 9 9 9 1 9 9
2 8 8
65 13 9 9 1 8 9 8 7 13 15 9 2 7 13 9 9 0 1 9 0 13 15 1 9 9 8 1 8 9 9 0 1 10 9 2 14 7 10 9 13 9 7 9 0 9 15 9 15 13 15 9 0 7 1 9 0 2 1 9 9 1 0 9 0 2
63 13 9 0 0 9 13 1 9 9 9 9 1 9 2 15 7 15 13 1 9 9 9 9 0 1 9 0 7 13 1 9 9 9 1 9 9 7 9 15 9 1 10 9 1 9 0 15 13 1 9 9 1 9 7 9 9 1 9 9 9 9 15 2
96 7 13 9 9 0 9 8 8 8 1 2 9 2 7 9 9 1 9 13 9 2 1 9 10 13 1 9 0 0 14 13 1 15 9 1 9 15 13 1 15 9 9 0 1 9 0 0 7 9 0 0 1 9 0 1 9 9 9 1 9 0 7 9 0 7 0 0 2 7 13 7 10 9 13 9 0 9 1 9 15 1 9 8 0 2 7 13 9 7 13 9 1 9 9 9 2
75 7 15 13 1 7 9 10 9 13 1 9 0 8 13 15 9 9 1 9 9 8 8 13 12 9 13 9 15 1 9 9 1 9 15 2 7 13 10 9 8 9 1 9 9 2 7 13 10 9 7 13 9 9 0 0 7 14 8 1 9 10 9 7 13 9 1 9 9 1 9 0 1 9 0 2
69 7 7 13 9 9 9 1 9 1 0 1 9 13 9 1 15 9 9 9 15 1 9 9 0 13 1 15 9 2 9 15 13 1 9 0 9 1 9 10 9 1 9 9 0 0 2 7 13 8 8 9 1 9 10 9 1 9 14 8 1 15 1 9 10 9 7 9 15 2
77 7 13 9 2 8 8 8 2 1 8 8 8 2 7 8 8 8 13 0 12 9 1 9 13 1 15 1 9 15 0 1 9 7 9 0 7 0 7 0 7 15 13 1 9 1 2 9 2 9 9 2 7 13 7 15 14 9 1 9 9 1 10 9 2 7 9 9 1 0 9 1 9 10 0 1 9 2
55 7 13 1 9 9 1 9 0 15 13 15 10 9 7 15 13 9 1 9 9 9 9 0 1 9 9 15 1 9 1 9 7 9 7 9 9 0 2 7 9 9 7 9 15 1 9 15 13 9 0 13 1 9 0 2
105 7 13 9 9 9 9 2 8 1 9 2 9 8 8 9 9 8 13 9 15 1 0 9 0 8 8 13 1 9 0 1 0 1 12 9 1 9 0 2 1 9 7 15 13 15 9 9 15 1 8 14 13 12 9 2 7 1 9 10 9 0 14 13 9 9 15 13 1 9 12 7 1 12 9 0 2 8 8 1 9 12 12 9 13 9 9 9 0 0 1 9 1 9 7 9 15 13 15 13 9 0 1 9 0 2
39 7 13 8 7 9 9 13 9 9 0 2 7 13 9 15 1 9 9 2 9 1 9 8 1 9 15 9 9 1 9 9 1 9 7 1 9 9 15 2
40 7 1 9 9 12 1 9 8 13 9 9 2 8 1 9 2 9 9 9 0 1 1 9 0 15 13 15 1 9 9 7 13 15 9 9 9 9 1 9 2
10 2 9 0 2 0 1 9 15 9 0
45 1 2 8 2 9 10 1 12 9 2 7 9 0 13 9 2 9 8 2 0 1 9 0 2 7 14 13 2 1 15 13 9 9 9 1 9 0 2 15 9 0 0 1 15 2
79 8 9 7 2 8 8 2 13 1 9 15 0 2 8 8 9 8 9 0 2 2 2 9 0 2 14 9 9 0 2 2 2 8 8 9 9 0 2 2 2 7 15 8 9 1 9 2 2 2 1 7 13 2 1 9 0 2 14 13 8 8 9 9 7 9 9 15 0 1 9 2 8 2 1 9 0 2 2 2
13 14 3 1 15 2 8 2 9 8 0 1 9 2
80 8 1 9 14 2 7 14 13 13 9 1 8 8 8 1 7 15 0 9 0 2 2 2 7 7 15 2 7 8 0 8 2 7 13 2 8 8 9 15 9 8 0 2 7 7 7 15 13 1 2 9 9 15 2 3 1 8 8 8 8 13 1 15 1 9 2 8 8 8 0 2 7 1 9 2 8 8 8 0 2
42 8 3 9 0 1 9 2 2 2 7 2 8 2 8 0 0 0 1 8 9 2 2 2 7 1 9 15 9 15 13 2 8 2 1 9 0 1 9 2 2 2 12
49 7 1 9 1 9 0 7 0 0 1 9 2 7 9 2 1 9 0 1 2 9 0 2 7 7 9 9 3 13 7 12 9 13 9 0 0 2 7 9 15 1 9 2 14 0 0 1 15 2
4 9 8 8 2
15 7 9 9 1 9 0 2 2 2 7 2 9 2 0 2
72 10 9 8 2 0 2 9 0 1 9 9 0 8 8 8 8 1 9 8 0 7 0 8 1 15 1 9 0 8 7 0 2 9 1 15 1 9 0 0 2 2 2 7 15 8 9 15 13 1 8 9 2 7 9 15 13 1 9 2 7 1 9 2 1 9 1 9 0 1 10 9 2
155 14 13 9 8 0 1 9 1 2 9 0 2 0 9 0 8 8 2 7 13 3 9 0 0 2 7 13 9 0 9 9 0 2 2 2 7 2 8 2 0 2 1 15 15 9 7 9 9 0 0 1 9 0 9 8 0 2 9 7 9 7 9 2 8 8 9 2 13 1 0 1 8 7 14 13 8 1 9 10 15 8 1 9 0 2 2 2 7 7 15 8 1 9 9 2 7 10 9 8 0 3 7 13 13 9 7 9 0 2 8 8 13 2 8 2 8 1 0 8 2 9 2 0 9 2 2 2 3 2 8 2 2 2 2 8 8 8 13 15 7 13 1 9 15 8 0 1 9 0 1 8 8 8 8 2
49 7 15 9 9 0 8 1 2 9 0 2 14 13 3 1 9 8 0 8 13 8 1 15 1 8 8 8 2 8 2 2 13 9 0 1 9 2 13 1 9 15 8 9 9 1 2 8 2 2
71 13 1 9 7 8 1 10 9 7 8 8 10 9 0 8 15 8 8 1 8 9 1 9 0 0 2 8 8 13 7 13 10 9 1 9 1 9 12 2 2 2 1 15 13 9 7 3 9 8 1 9 14 8 8 0 1 9 0 0 2 2 2 8 8 8 8 13 13 9 0 2
62 9 0 2 0 2 15 9 8 2 9 0 2 1 9 8 8 1 15 1 15 9 15 0 1 9 0 1 9 15 0 0 2 1 15 15 1 9 15 8 2 9 9 1 9 10 15 0 2 3 9 10 15 2 8 2 1 9 0 0 1 9 2
54 8 13 8 0 7 0 8 8 1 9 9 2 9 0 2 8 8 8 1 2 9 0 2 3 7 15 13 9 0 1 9 2 9 2 8 2 9 1 10 9 0 1 9 0 8 8 8 0 1 9 0 2 0 2
76 7 7 13 9 15 13 15 8 0 0 1 9 0 1 9 9 2 9 2 15 9 0 8 8 0 8 2 7 14 2 9 2 8 7 7 8 8 8 1 9 9 0 0 1 12 1 8 9 0 2 14 13 7 13 8 0 1 9 1 9 8 2 8 2 2 7 7 13 10 9 14 13 1 9 15 2
162 10 9 0 1 9 15 0 2 9 1 2 9 2 0 7 3 0 7 13 9 9 0 1 9 9 9 10 1 12 9 2 1 9 9 1 9 0 1 9 0 2 2 2 10 9 0 13 0 1 9 1 9 0 0 7 0 1 2 9 0 2 1 9 15 1 9 1 9 2 7 9 9 9 0 2 7 9 0 9 1 2 9 0 2 0 7 15 0 0 1 9 0 2 1 15 14 13 2 9 0 2 2 1 15 15 9 7 9 9 0 1 9 0 2 1 9 9 2 7 13 9 1 2 9 2 1 9 2 2 2 0 1 15 15 2 9 2 9 1 15 13 13 2 9 0 0 2 1 9 2 9 2 0 1 9 1 9 9 8 1 9 2
42 14 14 13 2 9 0 2 0 1 9 1 9 15 0 1 9 9 8 1 8 0 8 2 2 2 7 13 0 9 9 0 1 15 15 0 1 9 8 8 8 8 2
19 9 9 14 12 1 9 0 0 0 8 2 1 8 8 13 8 9 9 9
142 13 9 0 0 1 9 0 0 0 9 15 0 12 1 9 2 8 1 9 0 1 8 9 0 7 9 1 9 2 2 3 1 9 8 2 1 9 9 0 0 9 8 8 2 8 8 8 8 2 8 8 9 9 9 9 8 2 7 9 9 9 8 8 8 9 8 8 2 8 8 8 8 8 2 8 8 9 9 9 0 8 8 9 0 0 1 9 8 8 2 8 8 9 0 0 8 8 2 8 8 8 9 9 9 1 9 0 8 8 2 8 8 9 0 1 9 7 9 9 0 7 0 8 8 7 0 2 7 9 0 7 0 1 8 7 8 8 8 8 7 8 2
109 1 9 9 1 8 9 9 0 7 0 1 9 0 0 8 8 2 13 8 8 1 8 9 9 1 9 7 1 15 1 9 0 2 2 8 8 7 15 8 8 8 9 0 1 9 7 1 9 15 0 1 0 9 9 2 7 0 15 7 9 9 15 13 1 15 8 9 8 8 9 1 9 9 13 1 8 8 8 8 8 8 8 8 8 2 8 8 7 9 0 1 9 7 9 13 7 13 7 13 7 13 9 8 8 1 9 0 2 2
53 7 13 8 1 9 9 8 8 8 8 1 9 12 9 9 1 9 9 2 7 13 9 9 9 0 1 9 0 8 8 8 8 8 8 8 8 1 9 0 8 1 8 9 0 7 9 8 8 7 9 9 2 2
72 7 1 9 15 2 13 8 8 1 9 15 1 9 9 1 9 9 1 9 1 9 15 8 8 1 0 8 9 2 7 13 1 0 0 7 9 8 0 1 9 1 8 8 8 8 7 8 7 8 15 13 15 8 1 9 2 1 9 1 9 9 1 9 9 1 9 2 9 1 12 9 2
71 7 13 2 2 14 9 1 7 8 8 8 1 10 9 15 15 9 15 8 1 15 2 7 6 8 13 1 15 9 1 8 8 8 2 7 1 0 9 8 2 7 14 8 9 7 9 15 14 13 1 15 8 8 8 1 9 8 8 7 9 8 8 8 8 8 9 0 7 0 2 2
45 7 13 8 8 7 9 13 9 1 9 9 0 1 9 1 9 15 1 9 9 9 9 7 1 9 15 1 9 9 0 8 8 9 1 9 8 8 8 8 8 9 0 1 9 2
50 7 13 2 2 7 9 15 9 9 0 1 9 0 7 0 7 0 7 0 2 7 7 15 13 9 9 9 9 1 9 9 9 15 8 9 9 7 9 0 8 8 8 8 15 13 15 9 0 2 2
102 8 8 13 15 8 8 8 13 2 2 8 8 8 9 2 8 8 8 13 7 8 8 1 9 9 9 8 8 8 7 8 8 1 9 2 8 8 1 8 9 9 0 7 9 0 7 1 8 9 9 0 15 8 9 9 8 8 9 2 7 1 9 1 8 7 9 15 8 8 8 2 8 8 8 1 9 8 15 13 9 1 9 7 9 7 13 1 9 2 7 9 0 15 8 8 2 7 1 15 8 2 2
49 7 13 1 15 13 1 15 8 0 1 9 0 8 8 9 12 1 7 13 9 9 9 12 1 12 1 9 2 7 7 13 1 9 9 9 8 8 1 9 1 15 1 15 9 9 7 9 9 2
98 7 1 9 2 13 9 9 13 9 8 2 7 1 9 9 1 9 9 1 9 8 7 9 10 9 8 8 8 1 9 2 9 9 2 9 9 2 9 9 7 9 0 1 15 2 8 8 9 9 7 9 9 2 9 1 9 7 9 1 9 7 9 7 9 1 9 9 2 9 9 1 9 7 9 9 1 9 0 2 7 9 1 8 9 0 8 8 9 1 9 9 8 8 0 8 8 9 2
29 7 1 9 9 2 13 1 9 9 0 1 8 8 1 9 9 7 9 7 9 0 7 9 7 9 0 7 0 2
10 9 7 9 8 13 9 9 1 9 9
47 13 9 0 1 9 9 9 9 9 7 9 9 0 0 9 8 11 8 8 7 9 9 1 9 8 8 8 8 2 1 9 13 15 9 12 2 12 0 1 9 2 9 9 1 9 9 2
16 7 13 9 9 0 13 1 9 0 1 9 14 13 1 15 2
32 7 14 13 9 9 9 7 13 9 8 1 9 0 8 1 2 9 1 9 9 1 9 7 13 9 0 13 1 9 9 2 2
43 7 13 8 7 9 2 13 0 1 9 7 9 2 7 15 13 7 15 2 1 9 15 13 15 13 1 9 2 7 13 7 2 9 0 1 9 14 13 9 1 9 2 2
47 7 13 9 9 8 1 9 8 8 8 9 1 7 15 2 0 13 9 0 1 9 1 9 2 7 13 7 13 2 9 1 9 1 9 0 4 1 9 0 7 3 2 7 1 9 9 2
43 7 13 8 1 9 1 2 9 2 1 7 2 9 0 9 7 9 0 2 7 13 7 2 0 1 9 9 1 9 14 13 0 1 9 9 9 1 9 7 9 15 2 2
12 7 13 9 9 15 1 9 9 15 1 9 2
48 7 13 9 9 0 1 7 9 9 13 1 9 13 9 1 9 2 9 0 2 0 1 7 2 9 0 1 15 13 8 0 7 13 1 9 12 9 9 0 1 12 12 9 1 10 9 2 2
17 7 13 1 7 9 15 13 12 1 12 1 9 15 0 1 9 2
50 7 13 9 8 8 13 9 0 1 7 13 8 8 1 9 0 9 8 11 8 11 8 8 9 9 9 7 9 1 9 0 2 7 9 8 8 8 9 9 9 2 7 9 9 0 7 0 7 0 2
9 9 2 0 2 1 9 0 13 9
59 13 9 2 0 2 1 9 0 9 0 1 9 9 15 1 9 1 9 1 9 7 9 9 9 9 1 9 15 0 15 13 1 9 9 8 8 7 9 15 0 1 15 7 15 13 0 1 9 15 1 9 0 1 9 0 1 9 0 2
114 0 7 0 9 9 15 13 9 12 2 12 0 1 12 9 9 7 15 13 1 9 15 2 7 9 15 13 15 9 15 0 1 9 0 0 2 9 1 9 9 0 7 0 7 0 2 13 1 9 0 13 15 13 0 9 15 1 9 1 9 1 9 9 15 2 14 3 7 7 9 9 2 9 2 1 0 9 0 7 9 1 15 13 1 9 2 9 2 1 15 13 1 12 7 12 9 13 1 15 9 0 2 1 9 15 0 1 9 9 2 1 9 9 2
68 0 7 9 0 1 9 0 13 9 0 1 9 1 9 0 15 13 9 9 1 9 9 0 9 1 15 13 9 15 1 9 9 0 1 9 0 1 9 0 7 0 2 7 14 13 1 9 9 0 1 9 1 0 7 9 1 15 7 9 1 9 9 1 9 1 1 9 2
26 7 14 14 10 9 13 1 9 9 1 9 1 10 1 15 1 9 9 9 1 9 0 1 9 0 2
71 7 13 7 9 1 9 9 2 0 2 13 0 1 9 9 0 1 9 9 0 1 9 1 9 9 0 1 9 9 7 9 0 1 9 9 0 1 9 9 1 15 1 9 9 10 13 9 1 15 7 9 15 1 9 9 0 1 9 9 0 9 0 1 9 15 1 9 9 0 0 2
127 7 1 10 9 13 9 9 1 2 9 1 9 15 13 9 1 15 2 2 7 13 9 0 1 9 9 8 8 2 9 0 1 9 9 1 9 15 14 13 9 9 2 1 9 9 2 8 2 15 13 9 2 12 2 12 2 12 2 7 15 2 1 9 9 8 8 9 0 1 1 10 9 8 8 8 8 1 9 9 1 15 2 2 0 1 7 2 0 9 13 7 14 13 1 9 0 7 7 13 1 9 1 9 9 9 0 1 9 9 7 13 1 15 9 9 1 9 0 9 15 7 13 9 9 1 9 2
8 12 12 9 9 0 1 9 0
47 13 9 8 8 9 9 7 9 0 7 9 12 14 13 9 9 12 9 0 0 1 9 0 0 13 9 15 12 12 9 7 13 9 15 12 12 9 0 13 1 9 12 8 1 9 9 2
73 7 13 8 2 8 7 10 9 13 12 9 0 2 7 12 1 9 7 9 7 9 0 12 1 9 7 9 15 2 7 12 1 9 7 9 15 7 9 7 9 7 12 9 1 9 0 2 7 12 1 9 0 7 0 7 12 9 1 9 0 7 0 7 1 9 9 7 9 7 0 7 9 2
64 7 13 7 9 0 13 1 9 0 1 7 9 2 7 13 9 9 1 12 12 9 13 12 5 1 9 9 0 1 10 9 2 7 13 1 15 9 9 7 9 1 9 12 5 2 7 0 1 9 12 5 2 7 9 9 0 7 9 15 1 9 12 5 2
94 7 13 9 8 8 8 9 9 9 0 1 9 7 9 0 13 9 9 0 0 2 7 1 15 12 9 1 9 12 9 2 7 12 8 8 0 7 12 1 9 9 0 7 12 1 9 2 7 12 1 0 1 9 7 12 1 9 9 0 7 12 1 9 9 8 8 8 8 2 7 1 15 1 9 9 1 9 2 7 9 1 9 1 8 1 9 0 8 7 9 0 1 9 2
41 7 13 10 9 12 9 1 9 8 8 0 12 1 9 8 0 12 8 8 7 9 1 9 8 0 7 9 1 9 0 8 8 8 2 7 12 9 1 9 8 2
77 7 13 8 2 0 7 9 9 0 0 9 9 15 1 9 12 13 3 9 0 0 1 9 9 0 1 9 2 13 9 15 12 9 1 9 9 9 9 7 9 1 9 7 1 9 9 9 1 9 9 9 1 0 2 7 9 0 1 9 9 1 9 9 0 1 9 1 9 1 9 0 0 7 9 9 0 2
15 7 9 9 0 1 9 9 7 9 7 9 7 9 0 2
52 7 13 1 7 15 14 13 9 9 1 9 9 0 0 15 13 1 9 9 1 9 1 9 12 9 8 8 12 8 2 8 8 1 9 1 9 12 9 8 8 1 9 9 0 1 1 9 0 1 10 9 2
7 12 12 9 9 9 9 0
42 13 9 9 0 1 9 9 0 15 13 9 15 1 9 9 0 9 1 15 13 9 15 1 9 9 1 9 12 12 7 12 12 9 2 2 15 13 12 12 9 2 2
48 7 13 0 9 1 9 0 0 7 9 9 15 13 9 15 1 9 9 0 13 12 12 7 12 12 9 2 12 12 9 2 1 12 12 7 12 12 9 2 12 12 9 2 1 9 9 0 2
30 7 13 9 7 9 9 9 0 1 9 12 9 13 12 12 7 12 12 9 1 12 12 7 12 12 9 1 9 9 2
35 7 1 15 13 1 9 0 1 9 12 9 7 14 13 1 9 9 0 12 12 7 12 12 9 1 12 12 7 12 12 9 1 9 9 2
29 7 13 9 1 7 9 9 9 0 1 9 12 9 13 1 9 9 15 15 13 1 1 12 12 7 12 12 9 2
16 0 0 13 1 9 9 9 9 1 9 0 0 1 9 9 0
77 13 0 0 7 9 1 9 1 9 9 9 9 0 0 1 9 9 9 1 9 9 12 5 1 9 9 9 9 9 0 7 9 9 10 9 7 9 1 15 2 7 13 9 1 7 9 10 9 1 9 15 9 9 9 9 0 7 9 9 1 9 0 7 3 9 1 9 0 15 13 1 9 9 1 9 0 2
67 7 13 9 7 10 9 14 13 9 1 9 7 13 1 9 9 0 1 9 7 14 13 1 9 9 9 1 9 15 1 9 7 9 10 9 0 9 1 9 15 2 7 13 1 7 9 10 9 0 14 13 9 1 9 0 7 13 1 9 15 9 0 13 9 1 9 2
119 7 13 9 9 9 0 9 8 8 7 9 1 9 10 9 0 0 15 9 9 0 0 7 13 9 9 1 9 9 1 9 0 2 0 7 9 9 9 0 13 9 15 1 9 9 7 13 9 9 0 1 9 2 8 8 9 1 9 9 9 9 9 9 0 7 9 1 9 9 0 1 9 9 9 0 1 9 2 7 13 7 9 14 13 1 12 9 7 14 13 0 7 7 9 9 7 9 14 13 1 15 9 7 14 13 9 0 9 9 9 15 0 1 9 0 0 1 9 2
148 7 1 9 15 2 13 9 9 9 9 9 0 8 8 7 9 10 9 0 0 1 9 12 5 14 13 1 9 0 13 9 9 9 1 9 9 9 0 7 13 9 1 9 9 7 9 15 9 1 9 15 1 9 2 7 7 10 9 14 13 9 0 1 9 1 9 9 0 1 9 9 1 9 7 9 9 15 1 9 0 2 7 13 7 0 9 15 9 9 9 1 9 1 9 9 9 0 1 9 15 1 9 0 2 0 7 9 9 0 1 9 0 9 7 14 13 9 15 7 9 15 2 7 13 1 9 9 1 9 1 9 8 7 9 1 9 0 7 9 9 9 7 9 9 1 9 0 2
85 7 13 9 9 9 0 0 8 8 8 7 15 1 9 0 9 9 0 1 9 7 1 9 13 12 5 7 13 9 1 9 1 9 0 1 9 0 0 7 10 9 14 13 1 9 9 7 13 9 9 0 15 13 15 9 1 9 13 12 5 1 9 15 13 1 15 9 1 9 1 0 1 12 5 9 15 13 9 0 1 12 12 9 0 2
39 7 13 7 9 0 13 1 9 0 1 10 9 0 7 9 13 1 9 9 15 1 9 9 0 2 7 7 15 13 9 0 1 9 1 9 9 12 0 2
97 7 13 9 0 9 8 8 1 7 0 9 1 9 9 9 1 9 1 9 0 14 13 1 9 1 9 1 9 1 9 2 0 7 9 1 9 9 13 7 13 1 9 9 7 9 0 0 7 9 9 1 9 9 8 1 9 0 1 9 9 0 1 9 1 9 9 2 7 13 7 9 9 9 14 13 7 13 1 9 9 0 1 9 9 7 9 9 0 7 9 9 1 9 1 9 0 2
55 7 13 8 1 7 8 10 9 1 9 9 9 9 9 0 1 9 2 7 13 1 7 8 1 9 9 9 9 0 1 9 7 9 9 15 1 9 7 8 1 9 0 1 10 9 7 13 1 9 9 9 9 0 0 2
10 9 0 1 9 1 9 9 2 0 2
78 1 0 9 0 1 9 9 0 8 8 15 13 15 1 9 7 13 1 15 7 9 15 14 13 9 0 1 9 9 0 1 9 9 1 15 13 9 9 9 9 0 1 9 13 1 15 9 9 9 13 1 9 9 12 12 9 0 1 9 8 9 15 13 15 8 8 8 8 8 9 1 9 9 0 0 1 9 2
92 7 1 1 9 0 7 0 0 7 14 9 0 14 13 15 8 0 1 9 1 9 9 9 9 0 2 7 15 1 9 9 0 1 9 9 2 7 1 1 15 9 15 13 1 15 9 0 9 1 9 15 0 2 9 14 15 1 9 10 13 15 1 9 9 1 9 2 9 15 13 9 0 1 9 0 1 9 7 9 9 2 7 13 1 9 9 9 0 0 1 9 2
4 1 15 2 2
44 7 1 9 9 0 0 1 9 7 9 0 2 13 1 9 0 0 9 9 13 9 0 1 9 9 9 0 15 13 1 9 0 1 9 0 7 9 15 13 15 1 0 2 2
23 7 13 9 7 9 0 13 9 1 9 9 15 13 1 15 9 1 9 9 1 9 0 2
54 7 1 1 9 7 14 9 2 9 0 2 7 2 8 2 7 15 13 1 9 0 9 8 8 8 15 13 1 10 9 0 7 0 1 8 8 8 13 9 9 15 9 10 9 1 9 1 9 1 0 9 1 15 2
112 7 1 9 1 7 0 1 9 8 13 14 13 9 9 10 9 1 9 7 9 15 9 9 0 0 1 9 0 2 7 7 9 1 15 14 13 9 7 0 1 9 0 0 2 8 7 9 0 13 9 9 8 1 9 10 13 15 1 9 9 0 1 9 0 1 9 0 2 0 9 7 9 0 2 7 7 10 9 13 1 9 9 0 7 9 15 13 9 1 15 1 9 9 9 0 2 7 7 9 9 1 9 9 15 9 1 9 1 9 9 0 2
65 7 13 10 9 0 7 3 9 0 1 9 1 9 13 1 9 0 0 2 7 15 13 9 0 1 9 0 2 8 7 3 9 9 0 1 9 7 9 0 1 9 9 0 2 7 9 8 1 9 2 7 7 10 9 13 9 0 0 1 9 9 15 1 9 2
16 9 0 1 9 9 13 9 0 12 9 7 9 1 9 9 8
57 13 9 0 2 7 9 9 1 9 9 8 14 13 9 13 1 9 1 9 0 0 1 9 9 13 9 15 1 0 9 2 9 2 2 7 7 15 13 9 9 9 7 13 15 9 0 2 9 1 15 13 15 8 0 1 3 2
25 7 13 9 0 0 15 13 15 9 0 1 9 0 7 9 15 13 9 9 0 1 1 12 9 2
50 7 10 9 0 1 9 9 9 0 7 9 7 9 9 2 14 7 9 13 7 0 1 9 8 1 15 1 15 9 7 8 7 9 7 8 2 14 13 1 15 9 0 13 15 1 9 9 1 15 2
33 7 13 9 9 1 9 0 7 9 0 1 15 1 15 9 9 7 9 15 14 13 1 9 0 14 13 1 15 1 9 9 0 2
55 7 13 9 13 9 9 1 9 1 9 0 7 8 1 15 13 1 9 1 9 1 8 2 1 9 9 15 7 14 0 1 9 15 13 9 1 15 14 13 1 9 0 2 1 7 9 15 13 9 9 9 7 13 9 2
43 7 13 9 0 1 9 9 0 1 1 9 0 0 1 9 9 12 9 2 9 2 9 7 13 9 9 1 9 2 9 0 2 7 9 0 1 9 9 0 1 9 15 2
35 7 13 9 0 1 9 9 9 1 9 9 7 9 1 9 9 13 1 9 9 0 7 9 0 1 9 1 9 9 1 9 7 9 0 2
38 7 13 9 2 7 9 8 15 13 1 9 12 9 9 0 14 13 1 9 1 9 9 0 15 13 15 9 0 1 9 2 9 0 2 1 9 12 2
36 7 13 9 0 7 9 0 9 1 9 0 1 9 13 9 9 1 9 15 1 9 0 1 9 2 14 7 15 14 13 9 0 1 9 9 2
24 7 13 9 7 9 13 9 0 1 9 1 9 0 2 7 15 14 13 9 13 1 9 15 2
13 14 9 7 14 15 1 9 9 9 1 9 9 2
18 7 8 15 13 1 9 9 0 1 9 0 13 0 0 1 10 9 2
26 7 13 9 0 13 9 9 1 9 9 9 8 1 10 13 1 9 0 7 2 8 14 13 9 2 2
33 7 4 3 9 0 1 9 9 9 0 1 8 1 9 7 9 7 9 7 8 7 9 0 0 0 1 9 1 1 8 1 8 2
15 9 13 9 9 9 9 1 8 1 9 12 12 9 1 9
46 13 9 1 9 9 0 3 7 15 13 9 9 9 1 9 9 9 15 13 1 9 9 1 9 9 1 9 8 0 1 9 0 1 0 1 9 2 9 2 0 1 9 13 9 9 2
38 7 13 9 0 1 9 1 8 2 13 9 9 1 9 1 9 0 9 9 7 13 1 9 12 12 9 0 1 9 2 7 1 12 12 9 1 9 2
26 7 13 9 2 13 1 15 12 9 1 9 7 9 13 1 15 12 12 9 7 15 13 9 9 2 2
38 7 13 9 14 13 12 12 9 1 9 1 9 13 15 9 0 1 9 9 9 9 1 9 1 9 9 0 2 7 13 9 9 12 12 9 1 9 2
75 7 13 9 9 14 13 1 9 9 0 1 7 15 13 15 0 15 12 12 9 1 9 9 1 9 1 9 1 9 15 1 7 13 1 9 0 1 9 9 2 9 2 9 0 7 13 9 9 9 15 1 7 15 1 9 1 9 1 9 9 1 9 0 15 13 15 9 9 0 7 0 1 12 9 2
35 7 13 9 9 1 9 1 12 9 1 7 13 9 1 9 9 9 1 8 9 0 0 1 9 0 1 9 13 12 1 12 12 9 0 2
34 7 13 9 9 0 1 9 1 9 9 1 9 10 0 15 12 12 9 7 15 9 15 13 13 15 1 9 9 0 1 0 1 9 2
33 7 1 9 0 13 8 8 9 9 1 9 9 0 7 9 9 9 1 9 9 13 1 9 13 1 12 12 7 12 12 9 0 2
8 9 9 13 1 9 9 9 9
62 1 9 9 0 1 9 0 9 9 1 9 2 7 7 9 0 1 9 8 8 13 0 1 9 15 13 1 15 0 2 1 9 9 1 9 9 9 15 1 9 0 7 9 15 1 9 1 9 9 15 2 3 9 7 9 9 9 1 9 13 0 2
39 7 1 9 7 9 0 13 9 9 9 1 9 9 9 7 9 15 1 9 9 15 2 7 7 9 9 9 1 9 9 9 13 13 9 7 9 9 3 2
41 7 13 9 1 7 13 9 9 9 2 9 2 9 9 1 9 0 1 9 12 9 13 1 15 9 9 1 9 9 1 9 9 9 1 9 9 15 1 9 0 2
18 7 13 9 9 1 9 10 9 7 9 9 9 0 1 0 1 9 2
39 7 1 9 7 9 13 1 7 8 8 9 9 0 15 0 9 1 9 1 9 9 15 2 7 7 9 0 13 8 8 14 1 9 9 9 15 1 9 2
16 7 13 9 1 9 0 15 13 15 9 0 1 9 0 0 2
39 7 13 9 13 1 9 15 1 9 0 9 0 1 9 9 7 13 7 15 13 9 1 9 1 9 7 13 12 1 15 2 7 15 14 13 9 1 9 2
28 7 13 9 1 9 9 1 9 15 7 13 9 9 1 9 0 1 9 0 0 9 0 7 13 9 9 15 2
55 7 1 0 1 9 1 9 15 13 1 9 7 9 13 1 2 9 0 1 9 2 7 7 15 13 8 0 1 9 1 9 7 7 8 13 9 9 1 9 7 7 13 0 1 9 15 9 1 9 7 9 1 9 15 2
37 7 1 9 9 15 13 15 9 15 1 9 9 0 7 9 1 9 7 9 0 2 7 7 8 8 13 1 9 0 7 13 9 9 0 1 9 2
28 7 7 9 15 9 9 0 1 9 9 9 0 1 9 13 1 15 9 1 9 1 9 13 1 15 9 0 2
50 7 3 15 13 7 9 9 9 1 8 8 1 9 9 15 1 9 0 1 7 13 1 15 9 9 9 1 15 1 15 9 7 9 7 9 2 7 13 9 15 7 13 9 9 7 13 1 9 15 2
62 14 9 0 15 13 7 14 15 14 13 1 9 1 15 9 1 9 0 1 9 9 8 8 8 7 9 9 8 8 15 13 13 9 9 0 2 7 0 9 9 9 8 8 15 13 1 9 0 13 15 1 9 12 0 1 1 9 15 1 9 0 2
61 7 8 13 1 9 1 9 0 7 1 9 14 13 9 9 15 2 7 15 13 1 9 9 15 1 9 0 3 2 7 15 9 9 0 1 9 9 15 15 13 1 15 8 2 15 13 7 9 12 13 12 2 15 13 1 9 9 15 9 0 2
65 7 1 9 2 3 1 9 9 13 1 9 0 1 9 9 9 8 8 2 7 13 9 9 8 8 8 8 7 9 9 8 8 8 7 9 9 0 8 8 2 12 13 9 15 0 7 9 15 1 9 1 9 9 0 2 7 1 2 9 0 2 1 9 0 2
12 7 13 0 1 7 9 15 0 15 1 9 2
19 7 7 9 15 1 9 8 13 7 13 8 8 0 1 9 9 9 0 2
29 7 13 0 1 9 12 15 13 1 15 8 1 9 9 7 13 1 9 7 8 13 9 9 7 0 9 1 9 2
11 9 9 0 13 8 7 13 1 9 0 0
39 13 9 9 0 2 8 8 2 9 12 2 12 0 1 8 2 9 0 9 0 1 9 0 2 8 8 2 7 13 15 1 9 9 15 1 9 0 0 2
95 7 1 0 7 13 8 1 9 7 2 9 0 2 14 13 9 9 15 7 7 13 9 1 9 0 2 7 1 15 7 15 13 1 9 0 1 9 9 9 2 7 14 13 1 15 7 13 1 9 10 9 0 1 9 0 1 9 9 9 0 1 9 0 15 14 13 9 1 8 1 9 9 0 2 7 14 13 1 15 1 9 9 1 9 15 0 1 9 7 9 15 1 9 3 2
83 7 13 9 8 1 8 7 9 15 1 9 9 1 9 2 7 13 9 9 0 9 1 9 9 0 1 9 0 1 9 9 0 2 7 7 2 9 0 1 15 14 13 1 9 9 0 0 1 9 9 15 2 2 7 15 14 13 15 9 1 0 9 1 9 9 7 15 13 1 9 15 9 1 9 9 9 15 13 1 9 1 9 2
36 7 13 9 1 9 9 1 10 9 7 13 2 2 14 9 15 13 1 9 9 2 1 9 2 15 14 13 1 15 7 13 9 10 9 2 2
33 7 14 13 1 15 1 9 2 8 2 2 9 0 0 2 15 13 7 13 1 9 15 9 9 0 1 9 1 9 15 9 0 2
38 7 14 13 9 1 9 9 7 1 8 1 10 9 1 9 14 13 9 9 8 8 2 1 9 9 0 1 9 13 1 9 7 13 9 1 8 8 2
10 9 0 1 9 9 0 1 9 7 9
49 13 9 0 0 0 9 9 9 0 1 9 9 0 1 9 7 9 1 9 0 1 9 0 0 1 7 9 10 9 14 13 9 9 15 14 13 1 15 9 0 0 1 9 1 9 1 9 0 2
55 7 13 8 8 9 9 0 1 9 0 1 9 1 9 0 1 2 9 9 2 9 9 1 9 9 1 9 10 9 0 7 15 1 0 7 13 9 1 15 9 9 9 1 9 0 15 13 9 15 1 9 0 1 9 2
64 13 9 0 1 9 15 1 9 15 13 1 15 9 1 9 1 9 0 7 13 7 9 13 9 0 1 9 10 9 7 13 9 9 1 9 9 1 9 9 0 1 15 1 7 9 0 7 0 13 1 9 9 1 9 9 9 7 9 0 9 0 7 0 2
47 7 13 8 8 7 9 0 0 13 9 0 13 1 15 9 9 1 9 13 1 9 7 9 9 8 8 1 9 0 7 1 9 9 13 9 1 9 7 13 9 9 0 12 1 10 9 2
28 7 13 9 0 7 13 9 0 1 9 0 1 9 0 7 13 9 0 1 9 9 1 9 9 0 1 9 2
5 9 1 9 9 9
16 13 9 9 9 1 9 0 1 9 0 0 12 2 12 2 2
23 1 12 12 9 1 12 12 9 1 9 12 5 1 9 0 1 9 0 0 12 2 12 2
24 13 9 13 15 9 8 8 8 9 9 1 9 9 9 9 1 9 9 1 12 12 9 2 2
16 1 12 12 9 1 9 9 15 1 9 0 1 9 12 5 2
28 13 9 7 9 9 9 13 1 9 0 1 9 0 0 1 12 12 9 1 12 12 9 1 9 12 5 2 2
20 1 9 15 13 9 9 1 9 9 15 1 12 12 9 1 12 12 9 1 9
8 12 5 9 1 9 9 1 8
39 13 8 8 9 9 9 0 7 9 9 1 9 13 1 9 9 9 0 1 9 1 8 1 12 5 7 13 1 12 9 1 9 12 1 12 9 9 12 2
69 13 7 15 13 9 1 9 0 1 9 9 0 1 9 7 9 7 9 1 8 13 7 9 13 1 9 12 5 7 13 1 12 9 1 12 9 1 9 12 8 8 9 1 9 9 9 9 8 1 9 1 9 12 7 15 13 8 0 1 9 0 0 1 9 1 9 9 3 2
31 7 13 7 9 0 13 1 9 9 0 1 9 12 9 1 9 12 7 3 9 9 15 14 13 1 9 9 9 10 9 2
7 9 13 9 9 0 1 9
23 13 9 12 2 12 0 8 8 9 9 0 1 9 9 0 1 9 1 9 9 0 0 2
41 13 8 1 9 9 9 12 2 12 0 13 9 9 1 9 0 2 9 9 1 9 2 8 8 2 0 15 13 1 9 1 9 9 7 13 9 1 9 9 0 2
23 13 8 9 9 1 9 9 1 9 7 9 1 9 9 1 9 9 15 0 1 9 0 2
26 7 13 8 8 9 0 1 9 0 7 8 8 9 9 8 13 1 8 9 9 9 1 9 8 8 2
14 7 13 8 1 9 9 1 9 9 9 9 1 9 2
22 7 13 2 8 2 2 2 8 14 8 9 1 9 7 14 8 9 1 9 2 2 2
26 7 13 9 0 0 0 1 8 8 9 9 0 1 9 9 8 15 13 15 1 9 9 9 1 9 2
18 7 13 9 0 1 9 15 1 9 8 1 9 9 0 1 9 0 2
16 7 13 8 8 9 9 0 0 1 9 15 9 9 1 9 2
22 7 13 9 8 8 0 1 9 1 7 9 9 15 13 9 1 9 9 9 1 9 2
33 7 13 9 1 9 7 9 1 9 0 7 0 14 13 1 9 10 9 7 7 9 9 14 13 0 1 9 9 1 9 9 9 2
28 7 13 9 9 0 1 9 1 9 1 9 1 9 8 8 0 2 0 15 13 9 9 1 9 1 9 0 2
12 7 13 9 14 13 1 9 9 9 1 9 2
12 7 13 9 0 0 9 9 9 9 1 9 2
27 7 2 9 2 13 9 0 15 9 1 10 9 0 9 12 2 12 0 1 9 9 1 9 9 0 2 2
5 9 9 9 9 0
31 13 2 9 2 1 9 9 0 1 9 9 8 8 8 9 9 0 9 12 2 12 0 7 9 9 8 8 9 1 15 2
17 13 9 8 8 0 9 1 9 0 1 9 9 9 1 9 0 2
16 7 13 2 9 2 14 13 1 10 9 1 9 1 9 15 2
18 14 13 8 8 1 9 1 9 15 7 13 0 9 9 1 9 0 2
26 13 9 0 1 2 9 2 7 1 9 8 8 9 9 1 9 9 7 9 7 9 0 7 9 15 2
36 7 13 9 8 8 8 1 9 9 9 15 1 0 15 13 15 1 15 9 0 7 15 13 7 13 1 9 9 0 1 9 0 7 3 0 2
29 13 8 8 1 9 0 1 15 1 9 0 8 8 8 1 9 15 2 7 13 9 9 15 0 1 9 9 2 2
16 7 13 9 9 0 1 9 9 15 1 9 0 7 9 15 2
52 7 13 1 10 9 7 9 0 1 9 9 13 1 9 9 8 9 0 1 9 0 2 7 13 15 8 8 8 13 9 9 0 13 1 15 9 0 7 13 9 1 9 9 7 9 1 9 7 9 13 9 2
26 7 13 9 9 9 1 12 9 0 2 7 15 9 13 15 9 7 13 1 9 9 15 1 9 0 2
14 7 13 9 1 9 9 9 1 0 9 7 9 0 2
19 13 9 8 8 8 8 2 9 9 9 1 9 1 9 9 0 1 9 2
18 7 13 8 8 9 9 9 9 0 1 9 7 9 15 1 9 0 2
23 7 13 1 9 1 9 9 9 0 2 7 9 1 9 9 9 9 1 9 9 9 8 2
12 7 13 9 0 1 9 1 9 0 0 2 2
30 7 13 9 1 9 10 1 9 8 8 9 9 8 8 8 8 2 7 13 9 9 8 1 9 9 9 9 9 0 2
18 7 13 9 9 9 1 9 9 2 1 9 9 9 1 9 1 15 2
33 7 13 2 8 2 1 10 9 1 7 15 14 13 9 9 9 7 13 9 7 9 7 9 0 2 1 9 1 9 9 9 9 2
31 7 13 9 1 7 9 0 14 13 9 15 9 1 9 9 1 9 9 9 1 9 9 0 1 9 0 1 9 0 2 2
9 7 14 13 9 9 9 1 15 2
12 7 13 9 9 9 9 0 1 9 10 9 2
30 7 14 13 9 9 1 9 9 9 7 9 9 0 1 15 2 7 13 1 9 9 9 9 1 9 0 1 10 9 2
11 7 13 0 9 15 1 2 9 0 2 2
30 7 13 9 9 0 1 8 8 8 8 7 9 9 9 15 1 9 1 9 9 1 9 15 1 13 9 9 8 8 2
8 9 9 9 0 13 1 9 0
30 13 9 9 7 9 9 1 9 9 9 9 9 9 0 7 0 7 0 9 15 1 9 9 1 9 0 7 9 9 2
16 13 9 1 7 9 13 9 1 9 13 9 0 1 9 15 2
50 13 8 1 9 9 9 9 0 1 9 0 7 15 13 15 9 9 8 8 1 9 0 1 9 9 2 7 13 15 9 8 8 8 9 9 9 0 2 7 9 8 8 8 9 0 9 0 7 9 2
37 13 9 8 8 8 8 9 9 9 9 9 0 1 9 9 0 2 7 13 0 1 9 0 1 9 0 1 9 7 9 1 15 13 1 9 0 2
36 7 13 7 9 9 0 7 0 13 12 7 12 12 9 2 7 13 1 1 12 5 1 9 9 0 15 13 15 9 0 2 7 13 9 9 2
24 13 8 7 9 1 15 0 1 12 9 1 9 9 0 7 14 13 1 15 1 12 5 3 2
9 7 13 9 1 9 13 12 5 2
18 7 13 7 9 0 13 12 12 9 13 9 15 1 9 0 1 9 2
47 7 13 9 9 9 1 9 9 0 1 10 14 13 12 5 3 7 13 2 8 2 1 9 9 0 1 9 9 0 1 1 9 7 9 7 9 9 8 8 13 0 1 9 1 9 9 2
28 7 13 9 8 8 8 9 0 9 0 1 9 9 9 0 1 9 1 9 9 1 9 9 9 1 9 0 2
50 7 13 9 8 8 8 9 9 9 0 7 9 0 13 9 9 1 9 7 13 9 9 1 9 0 0 15 13 1 9 2 7 13 7 10 9 15 9 8 0 7 9 9 9 1 9 1 9 9 2
11 9 2 9 0 2 1 8 7 9 9 0
70 13 8 8 8 9 0 1 8 9 9 9 9 9 0 1 8 7 1 9 9 8 8 13 9 1 9 9 0 0 7 9 9 0 1 1 9 9 1 9 0 1 9 7 9 15 0 14 15 1 9 10 9 14 13 0 1 9 0 1 9 0 0 7 13 9 15 1 9 0 2
76 7 13 9 9 1 9 13 15 1 9 9 0 1 9 9 0 1 9 0 1 9 1 9 1 9 0 1 9 9 9 0 0 15 14 13 1 9 12 1 9 1 9 9 1 9 0 1 9 0 7 14 15 1 9 0 7 13 9 0 9 10 9 15 13 7 9 1 9 13 1 9 0 1 9 9 2
85 7 13 9 9 0 9 1 9 9 0 0 7 1 9 8 9 0 8 1 9 9 0 7 7 13 1 9 9 1 15 1 9 8 1 9 0 1 9 9 0 1 8 7 9 0 0 1 7 13 1 15 1 9 9 0 0 13 1 8 1 7 13 1 9 9 0 1 9 15 7 1 9 1 9 0 7 13 9 10 9 7 9 9 15 2
104 7 13 8 8 8 1 9 9 0 1 8 13 1 9 1 9 0 1 8 7 9 0 9 0 1 9 0 7 9 9 9 9 0 7 9 9 1 9 9 0 1 8 1 9 15 9 9 9 1 9 0 7 9 9 0 1 9 0 7 15 13 13 1 9 9 9 9 1 8 14 13 0 7 9 9 1 9 9 15 13 0 1 9 9 0 7 9 0 1 9 7 9 0 1 9 9 1 9 0 1 9 1 9 2
8 9 1 9 7 9 1 9 9
102 13 9 1 9 0 9 8 2 1 9 15 12 9 1 9 9 1 9 9 2 9 9 2 1 9 13 1 15 1 9 12 9 1 9 15 1 9 9 15 9 9 0 1 9 1 9 0 7 9 1 15 2 1 9 0 1 9 7 9 0 2 1 9 9 8 1 9 1 9 0 15 13 1 15 1 9 1 15 1 7 15 13 1 9 9 1 9 9 1 9 9 7 9 15 13 1 15 1 9 1 15 2
62 7 13 9 1 9 9 0 1 9 2 7 1 9 15 9 9 0 9 8 8 2 14 13 9 12 2 12 0 9 9 0 1 9 8 8 9 9 0 8 8 8 9 0 7 9 8 8 8 9 9 1 9 9 9 1 9 9 9 7 9 9 2
33 7 13 9 1 9 9 1 9 9 12 0 1 9 12 0 9 9 1 9 9 8 1 9 10 13 1 15 7 1 15 9 8 2
21 7 13 9 1 9 9 9 1 9 9 13 1 9 1 9 1 15 1 9 9 2
12 9 1 9 12 9 0 0 1 8 0 1 9
12 1 10 9 13 9 2 9 0 2 9 0 2
69 13 9 8 8 1 9 0 13 15 1 9 9 15 13 15 15 1 0 7 13 9 1 9 7 13 15 13 15 2 9 0 2 15 13 9 9 7 13 9 0 0 1 9 0 9 7 13 8 1 9 15 0 1 12 12 9 1 9 9 15 1 9 0 7 9 9 9 15 2
86 13 8 1 0 15 1 9 9 1 9 1 1 9 9 15 7 9 9 9 1 9 15 2 9 2 9 2 8 8 2 9 9 2 1 9 0 0 2 2 7 13 9 15 1 9 15 1 2 9 2 0 2 8 8 2 1 9 8 2 7 13 1 15 9 0 1 9 1 9 12 9 0 1 9 7 1 9 1 9 2 9 1 9 9 2 2
120 7 13 8 14 13 9 0 1 9 15 8 8 7 15 13 15 1 1 2 8 2 7 15 9 0 13 9 9 9 2 2 1 9 7 8 9 15 14 13 9 8 8 7 13 1 9 15 1 9 10 9 2 7 1 9 7 15 13 9 1 9 0 15 13 2 2 15 13 9 13 15 2 2 7 7 13 15 13 9 0 0 2 7 15 13 9 9 2 1 9 8 1 9 0 1 9 10 9 0 1 8 9 15 0 15 13 15 1 9 15 15 13 3 3 1 9 0 1 9 2
106 7 8 14 9 1 9 15 2 7 14 15 13 8 1 7 13 2 9 0 2 1 0 0 8 1 9 15 7 15 13 9 1 1 9 2 7 7 13 9 0 2 8 8 2 1 9 1 9 9 0 1 0 8 0 1 9 14 13 15 13 1 9 9 9 2 1 9 9 1 9 2 7 13 0 7 0 1 10 9 0 15 0 8 2 7 13 7 15 14 13 9 8 1 9 0 1 15 12 9 1 12 9 13 15 8 2
62 7 13 9 1 9 15 14 13 15 7 9 9 9 9 14 13 1 9 9 0 2 7 15 15 9 9 7 13 9 0 0 1 9 2 7 15 9 9 9 15 13 9 1 9 0 2 7 15 13 1 9 15 1 9 0 2 9 1 9 9 2 2
45 7 13 8 8 2 9 9 8 8 1 12 9 0 9 9 1 9 9 0 8 2 7 13 7 15 7 13 9 0 8 1 9 12 14 13 12 9 13 9 15 1 12 9 12 2
28 7 13 8 8 2 8 8 2 1 12 9 0 7 13 1 2 9 0 7 15 13 9 0 1 9 2 2 2
109 7 13 8 1 9 9 7 1 9 8 2 7 13 9 9 0 0 2 8 8 2 7 13 1 9 9 15 13 15 9 1 0 8 2 7 13 2 7 1 9 0 8 9 0 2 14 8 7 15 8 8 14 9 9 15 13 1 0 9 1 9 9 13 0 7 9 2 7 8 8 13 1 9 2 7 13 8 8 2 9 1 9 9 0 1 9 9 0 1 9 1 9 15 13 9 0 7 9 15 0 9 1 9 0 1 9 1 9 2
68 7 1 7 9 0 0 7 13 15 9 9 9 15 7 14 13 8 0 8 8 8 2 0 2 2 7 9 9 0 13 1 9 0 2 7 1 9 15 8 8 8 0 9 9 1 9 9 1 9 0 2 7 9 9 1 9 9 7 13 7 0 13 9 1 1 9 0 2
84 7 9 9 9 9 1 9 9 2 13 1 9 15 13 1 15 8 7 13 9 15 9 9 1 15 2 7 13 1 9 9 2 2 13 7 13 15 1 9 7 13 9 1 9 9 2 7 13 7 13 9 15 1 1 0 9 1 9 13 1 9 8 2 7 13 7 14 13 9 9 1 9 0 2 7 13 9 15 1 0 9 2 2 2
9 9 8 12 2 12 2 12 2 2
59 7 14 13 9 1 9 1 9 1 9 9 9 2 7 7 13 9 0 8 13 1 9 9 1 9 15 1 9 1 9 10 13 15 7 13 9 15 2 1 9 15 13 1 15 9 9 1 7 15 13 1 9 9 0 7 13 9 9 2
43 7 9 9 0 13 0 2 7 1 9 12 13 9 12 0 2 13 9 15 1 12 9 1 9 12 2 8 8 9 1 9 13 1 15 8 8 7 13 9 1 9 2 2
69 7 9 1 9 15 13 15 8 9 12 13 9 9 0 0 9 1 9 0 12 9 7 13 1 15 7 9 15 1 9 9 0 1 0 2 8 1 9 2 1 9 0 1 9 9 9 0 1 9 0 2 9 2 8 2 9 2 9 2 7 9 1 7 13 9 7 13 0 2
115 7 7 13 8 7 13 9 9 9 0 2 13 9 15 1 9 9 9 0 2 7 13 1 15 2 9 0 7 0 2 14 13 9 15 1 0 9 0 2 7 13 1 9 0 2 2 13 1 9 0 7 13 9 8 7 1 15 9 9 1 9 15 9 9 0 2 8 8 0 1 9 7 1 9 0 7 0 1 9 15 9 15 13 0 9 1 9 2 7 14 8 7 9 15 1 9 14 13 9 2 7 14 13 1 7 15 9 1 9 0 1 9 9 0 2
60 7 8 7 9 15 1 0 9 9 1 9 9 15 0 14 13 7 15 14 13 9 10 9 1 9 15 1 9 15 7 13 7 15 13 1 7 13 9 15 1 9 7 13 9 0 15 13 1 15 2 7 13 1 15 9 15 13 7 13 2
13 9 13 9 0 1 9 0 0 9 1 9 9 0
43 13 9 0 7 9 9 0 0 1 9 9 1 9 9 0 0 15 13 15 9 8 8 14 13 1 9 1 9 0 1 9 9 9 9 7 9 0 7 9 0 1 9 2
19 7 7 15 13 0 0 1 9 0 1 15 13 9 9 9 1 9 0 2
48 7 13 9 8 8 9 9 9 0 7 9 9 9 9 0 7 9 0 0 1 9 9 0 13 1 9 0 1 9 0 9 1 9 9 15 7 9 9 15 1 15 14 13 1 0 9 0 2
59 7 13 1 7 9 0 13 0 1 9 15 13 9 7 9 0 1 9 9 0 0 1 9 0 1 9 0 1 9 9 0 1 9 9 0 7 9 9 0 9 1 9 7 9 9 0 7 0 7 0 1 15 13 1 9 0 1 9 2
39 7 13 8 7 9 0 1 9 9 0 13 0 1 9 1 9 0 7 13 15 0 9 7 13 1 9 9 7 13 9 1 15 7 14 13 9 1 15 2
50 7 13 7 9 0 13 9 0 1 9 7 13 15 1 9 3 15 9 0 7 0 9 1 9 9 0 1 1 9 7 14 9 1 15 14 1 9 9 7 13 3 9 0 7 0 7 0 7 0 2
40 7 13 9 0 1 9 0 7 9 0 0 1 9 9 13 0 9 0 1 9 0 7 13 0 9 1 1 9 7 9 0 9 0 1 9 9 7 9 0 2
41 7 13 7 9 0 9 7 15 13 13 1 0 9 0 14 7 15 13 13 9 9 0 1 9 9 7 15 15 13 13 1 9 15 0 7 9 0 13 10 9 2
38 7 13 9 0 1 9 0 7 9 0 13 9 0 1 9 9 0 1 9 7 7 9 15 13 13 13 13 1 1 9 9 0 7 9 9 9 0 2
33 7 13 7 9 0 13 9 7 9 1 0 1 9 9 0 7 13 1 9 0 1 9 9 7 13 9 1 9 0 1 9 0 2
35 7 13 1 7 9 9 9 9 13 0 1 9 9 9 0 1 9 0 0 7 9 0 13 9 0 1 9 9 0 7 9 9 0 0 2
49 7 13 7 9 0 13 13 1 9 0 9 9 0 1 9 1 9 9 0 1 9 7 9 1 15 7 7 14 13 9 0 1 9 10 7 13 15 9 9 0 7 15 15 13 15 9 0 0 2
59 7 13 1 7 9 9 9 0 1 12 9 2 0 1 12 12 9 2 1 9 0 13 1 9 9 1 9 0 1 9 0 1 9 9 9 1 9 9 15 9 7 9 14 13 1 9 1 9 7 7 9 9 0 1 9 13 9 0 2
43 1 9 15 13 8 8 8 9 9 9 7 9 0 0 1 9 9 0 13 9 9 9 1 9 9 7 9 1 9 0 9 9 7 9 0 7 9 1 9 9 9 0 2
10 1 9 9 2 9 12 12 9 1 9
79 13 9 9 9 13 1 9 9 7 13 9 0 1 9 0 1 9 1 9 9 9 1 9 0 0 1 12 5 1 9 12 2 12 1 12 5 12 2 12 1 9 9 15 13 15 9 9 1 9 9 9 1 9 9 9 13 1 9 15 1 9 7 1 9 9 0 1 9 9 1 9 7 9 1 9 9 1 9 2
37 9 0 13 1 9 9 1 0 9 0 0 7 9 9 1 9 9 0 3 7 13 9 1 9 0 12 9 1 9 12 1 15 13 13 1 12 2
24 13 9 7 15 13 8 8 9 0 7 9 0 13 1 9 0 1 15 13 1 15 9 0 2
65 13 9 9 9 7 9 8 8 8 13 1 9 2 7 9 15 13 15 9 13 7 9 15 13 15 9 9 0 7 9 0 9 1 0 7 1 9 2 7 7 9 15 13 14 13 1 2 8 2 0 7 9 2 8 2 13 8 1 9 9 0 1 9 0 2
56 13 9 9 7 9 0 1 9 9 1 9 1 9 0 0 1 12 5 9 12 2 12 1 12 5 3 9 12 2 12 7 13 9 0 9 7 0 0 13 7 0 1 12 12 9 1 9 9 0 0 1 12 12 9 3 2
80 9 1 9 1 9 13 9 15 9 9 7 13 9 0 1 9 9 0 1 9 12 5 9 12 2 12 1 12 5 8 9 8 8 9 9 1 9 9 9 8 8 13 7 9 13 1 9 9 0 7 13 15 1 9 1 9 9 9 7 9 9 7 9 9 9 0 7 9 1 9 1 9 1 9 9 9 7 9 0 2
75 7 13 1 7 9 0 13 1 9 1 9 9 7 13 1 9 9 7 9 1 9 9 1 9 0 2 7 1 0 13 9 9 1 9 8 13 15 9 7 15 15 13 1 9 9 0 1 9 9 7 13 9 9 7 9 0 0 1 7 13 1 15 1 9 9 7 1 9 7 13 1 2 8 2 2
77 7 1 9 9 9 7 9 9 0 8 8 13 1 9 9 9 7 9 9 7 9 9 0 15 13 15 9 1 9 15 1 9 9 14 7 9 9 0 1 9 9 0 14 13 1 12 5 1 9 12 2 12 1 12 5 1 9 12 2 12 1 9 9 1 9 9 1 12 12 1 12 12 9 1 9 9 2
40 9 9 7 15 13 9 13 1 9 9 13 7 9 10 13 15 9 1 9 9 7 9 14 13 1 9 1 9 9 7 7 15 14 13 14 9 1 9 2 2
44 7 14 13 9 13 9 9 9 0 1 12 5 1 9 0 0 7 13 1 12 5 7 15 10 13 13 7 13 9 9 1 12 5 0 7 15 14 13 9 7 13 1 9 2
41 7 13 9 1 7 9 1 9 9 0 1 15 7 9 9 13 7 1 9 7 13 9 1 9 0 1 12 9 12 2 12 1 12 12 9 1 9 12 2 12 2
47 9 1 9 15 7 1 15 13 9 13 13 1 9 0 7 0 0 1 9 9 7 1 1 9 1 9 13 9 1 9 9 7 9 0 9 1 9 1 9 7 1 9 0 15 9 9 2
23 9 13 3 7 9 9 13 9 0 7 9 0 7 0 13 15 13 15 0 9 1 9 2
46 7 1 9 1 9 0 7 0 7 1 9 10 9 7 14 13 1 9 9 1 12 12 9 1 9 12 5 1 9 9 1 12 5 1 9 9 7 1 9 12 5 1 9 0 0 2
39 9 13 3 7 15 13 9 12 12 9 1 9 0 1 9 7 9 9 9 1 9 15 1 9 9 7 9 15 13 15 1 9 7 9 7 9 9 2 2
28 7 13 9 1 1 9 15 15 13 1 9 0 1 9 0 9 0 1 9 12 12 9 0 1 8 7 8 2
42 7 13 9 0 1 9 1 9 9 9 0 1 9 9 7 15 14 13 12 8 9 1 9 12 1 9 13 1 12 8 9 7 13 9 1 9 0 1 12 8 9 2
29 7 9 7 9 13 9 0 7 15 13 9 15 12 7 12 12 9 2 7 1 9 13 1 12 5 1 9 9 2
74 9 9 0 13 1 9 15 13 1 15 9 0 7 0 1 9 9 15 12 9 1 9 1 9 12 7 1 12 7 1 15 9 1 12 1 12 12 9 2 8 0 1 12 1 12 8 2 9 2 8 1 12 1 12 8 9 2 8 8 1 12 1 12 8 9 7 9 1 12 1 12 8 9 2
25 7 13 9 7 9 9 9 0 14 13 1 10 9 12 5 1 12 5 1 0 9 1 9 0 2
32 7 13 9 9 9 1 9 0 1 7 15 13 9 0 1 9 9 0 0 7 3 13 9 0 1 9 1 9 9 9 0 2
33 7 13 9 1 7 9 0 1 9 1 9 0 13 3 1 9 9 0 1 9 0 7 13 1 12 1 12 12 9 1 8 9 2
21 9 10 9 7 13 9 15 7 9 1 9 9 7 9 9 0 1 9 10 9 2
20 7 13 7 9 10 9 13 1 9 1 0 1 9 7 8 9 1 9 0 2
15 9 15 13 1 15 9 15 9 9 1 9 9 9 9 2
31 7 10 13 15 1 9 1 9 9 0 1 9 7 10 9 14 13 9 0 1 9 0 2 7 1 0 9 9 9 0 2
73 7 13 9 7 9 9 9 7 7 13 9 15 1 9 9 9 8 7 9 9 14 13 7 13 9 9 1 9 9 8 8 1 9 0 3 14 7 15 14 13 9 1 15 1 9 1 9 9 1 9 0 9 1 7 9 14 13 1 9 9 0 1 9 9 1 9 15 1 0 9 15 0 2
33 7 1 15 13 15 9 1 9 15 13 9 9 9 0 1 10 13 9 9 9 0 1 9 1 9 0 7 9 0 7 9 0 2
20 14 7 15 1 9 14 13 1 9 9 0 1 9 9 0 15 13 1 9 2
6 9 13 1 9 9 0
17 13 9 0 0 1 9 9 9 9 0 0 1 9 1 9 0 2
17 13 9 2 9 9 9 0 1 9 0 1 9 13 1 12 5 2
31 13 9 9 9 9 9 9 0 0 1 9 0 1 15 1 12 12 9 9 12 2 12 1 12 12 9 9 12 2 12 2
11 7 13 1 12 12 9 9 12 2 12 2
30 7 13 9 0 0 1 9 9 1 12 8 9 1 12 8 9 7 1 12 8 9 9 12 2 12 1 9 12 5 2
27 7 13 9 0 1 7 9 9 0 0 1 9 9 2 13 9 1 9 1 9 9 9 0 1 9 0 2
34 7 13 9 9 1 9 9 1 12 12 9 9 12 2 12 7 13 1 12 12 9 9 12 2 12 7 1 12 12 9 1 9 0 2
25 13 9 0 1 9 9 9 1 9 9 0 9 1 9 12 1 9 12 7 9 12 1 9 12 2
22 13 9 12 9 1 8 0 1 9 0 12 2 12 1 9 0 9 15 12 12 9 2
16 7 13 9 1 12 9 1 9 0 12 12 9 1 9 0 2
41 7 13 9 9 9 0 9 1 9 9 7 9 9 1 12 9 1 9 12 12 9 7 13 1 12 9 1 9 12 12 9 1 9 0 1 9 0 12 2 12 2
17 7 13 9 9 9 1 9 9 9 1 9 0 9 0 7 0 2
24 13 9 1 9 9 1 9 9 9 0 1 9 9 1 9 9 2 8 2 1 9 12 5 2
18 7 13 9 9 1 9 1 9 9 0 2 7 9 9 7 9 9 2
26 7 13 9 9 8 9 9 9 7 9 0 7 9 8 9 9 9 0 13 1 9 9 0 1 9 2
9 12 12 9 9 0 7 0 1 9
71 13 0 9 0 9 9 0 7 0 15 13 9 9 0 0 1 9 9 7 9 0 1 9 15 7 15 1 9 0 7 0 7 1 15 13 9 9 15 13 9 15 1 9 9 9 0 1 0 1 9 9 0 7 1 9 1 12 12 9 13 9 15 1 9 0 0 7 8 7 8 2
29 13 7 9 0 1 9 13 9 9 0 1 9 0 7 15 1 9 9 0 1 9 0 1 9 7 9 7 9 2
10 9 0 1 9 9 0 1 9 8 8
52 13 9 0 8 1 9 1 9 9 8 8 9 9 9 9 2 1 9 9 0 1 9 9 1 9 9 9 0 1 9 1 12 9 2 7 15 13 1 9 9 9 9 1 9 9 9 0 8 8 1 9 2
14 7 13 9 1 9 0 15 13 0 1 9 8 8 2
51 7 13 9 9 0 1 9 1 9 9 8 8 9 9 9 9 14 13 1 9 15 15 13 15 0 0 2 1 7 9 9 9 1 9 8 8 1 9 2 13 9 1 9 0 7 9 1 9 0 0 2
33 7 13 9 7 15 13 15 0 1 9 14 13 9 15 1 9 9 7 15 13 13 1 9 9 7 9 9 7 13 9 9 9 2
19 7 13 9 7 0 13 9 7 13 1 15 12 9 7 13 1 8 8 2
36 7 7 10 9 14 13 7 13 9 2 9 1 7 9 0 13 7 15 13 1 9 9 9 7 9 7 13 15 8 0 1 9 9 1 9 2
27 7 13 9 7 9 9 9 13 9 1 9 12 2 7 10 13 9 0 7 0 9 9 9 9 15 0 2
53 7 13 9 1 7 9 0 1 9 1 9 13 1 15 9 1 9 7 9 7 9 13 9 9 7 9 1 9 7 13 1 15 1 9 0 7 14 13 1 9 0 2 7 15 15 13 15 9 0 0 1 9 2
8 9 0 13 9 0 1 9 0
35 13 9 0 1 9 7 9 1 9 15 9 0 1 9 1 9 0 1 9 0 1 9 0 0 13 1 12 12 9 7 13 1 9 0 2
57 7 13 9 9 0 1 9 8 8 7 9 1 0 9 15 1 9 0 7 15 13 1 9 9 0 8 8 7 9 8 7 9 0 1 9 1 9 9 1 9 9 15 13 1 12 12 9 7 13 1 9 0 7 1 9 9 2
43 7 13 8 1 9 1 15 13 9 12 2 12 0 7 9 9 13 1 9 15 0 0 7 9 0 1 0 9 13 9 1 9 15 1 9 1 9 7 9 7 9 0 2
40 7 13 2 7 9 9 0 0 0 1 9 13 12 12 9 2 12 9 2 0 1 0 1 9 2 1 1 13 9 2 8 2 12 12 9 2 12 9 2 2
32 14 9 7 14 9 13 15 9 9 0 8 0 2 0 1 2 7 15 14 13 1 9 9 9 0 1 0 1 9 0 2 2
13 9 2 8 13 9 9 0 0 13 9 9 7 9
67 13 2 8 8 2 7 9 0 9 8 8 1 9 9 9 0 1 9 9 9 7 9 1 9 0 0 1 9 15 13 15 9 0 0 7 15 9 9 0 1 9 10 9 1 9 0 1 9 9 9 7 9 1 9 0 1 9 9 0 15 13 1 15 8 9 12 2
78 7 13 9 0 0 0 9 13 1 9 15 1 9 0 9 2 7 9 0 1 9 9 9 0 1 9 9 0 1 9 9 0 9 13 9 1 9 0 7 0 1 8 1 9 15 1 9 9 9 15 0 1 9 0 7 9 0 2 7 9 9 9 1 9 12 1 9 8 0 9 15 9 1 9 9 9 0 2
70 7 13 9 7 10 9 14 13 9 1 9 9 0 1 9 9 9 0 2 15 13 9 0 1 9 0 15 13 15 9 9 12 2 7 9 12 1 9 0 1 15 1 9 15 13 1 9 15 0 1 9 9 7 9 9 9 1 9 15 0 1 9 0 7 0 15 13 1 9 2
33 7 13 9 0 0 1 8 9 1 0 1 9 9 0 15 13 1 9 0 15 13 15 1 9 8 9 8 13 1 9 9 0 2
65 7 13 9 0 0 1 2 8 8 2 7 8 1 9 9 1 9 9 0 1 9 0 2 7 15 13 1 9 9 1 7 8 14 13 9 1 9 1 9 9 0 1 9 0 7 9 9 0 15 13 1 9 0 9 9 9 15 1 9 15 1 1 9 0 2
46 7 13 1 9 15 1 7 13 10 9 0 9 9 9 7 9 0 9 0 1 9 9 7 9 1 9 0 2 0 7 9 15 13 15 8 9 9 9 0 13 1 9 1 10 9 2
41 7 13 1 7 9 1 8 0 1 9 9 0 1 9 9 1 9 1 1 9 2 9 7 14 13 8 8 0 1 9 7 9 1 9 9 0 1 9 9 15 2
45 7 13 9 9 0 1 9 2 0 7 9 0 15 13 9 0 0 13 0 9 0 7 13 9 9 1 9 15 7 9 15 1 9 1 9 9 7 1 1 9 1 0 8 0 2
87 7 9 1 9 0 1 2 8 8 2 7 14 9 0 1 8 13 0 1 9 9 1 9 9 15 13 7 13 1 9 8 1 9 9 9 0 9 1 9 15 1 9 0 1 9 9 0 15 13 15 8 9 0 1 9 9 1 10 9 7 9 15 1 9 9 15 0 7 9 1 9 9 0 1 9 9 0 1 9 1 9 0 1 9 9 0 2
108 7 13 9 1 9 9 12 2 12 0 1 9 1 2 9 0 9 7 9 10 9 2 8 7 9 0 9 0 13 9 1 7 9 13 1 9 9 9 15 13 15 0 9 0 0 9 9 1 9 9 15 7 9 15 2 0 1 7 9 0 1 9 0 1 9 0 1 9 9 0 1 9 7 9 1 9 9 9 0 7 1 9 15 9 9 1 9 9 0 1 9 1 9 0 7 9 0 0 1 9 9 9 1 1 9 9 0 2
50 7 13 10 9 1 9 9 2 8 8 2 9 1 9 9 9 0 2 15 13 9 0 1 9 0 0 1 15 1 8 1 9 12 2 9 9 0 1 9 9 1 9 0 0 7 1 9 9 15 2
44 7 1 9 2 9 0 1 9 0 2 13 9 0 1 9 1 15 9 12 2 12 0 2 7 9 9 7 9 0 2 9 0 0 2 13 1 9 9 15 13 1 9 9 2
61 7 13 9 15 13 1 9 0 0 2 1 9 9 1 9 15 13 1 9 9 0 7 0 7 9 9 0 1 9 0 7 1 9 9 1 9 0 2 9 9 9 7 9 7 9 9 1 9 0 1 9 9 1 9 9 9 7 9 7 9 2
74 7 13 9 0 7 9 0 1 15 13 15 1 9 7 9 9 0 1 0 9 9 0 1 9 7 1 15 7 1 9 0 0 1 9 7 9 0 2 9 0 0 2 1 9 0 7 9 9 15 7 9 9 0 13 10 9 2 7 13 9 1 9 9 9 9 1 9 10 9 9 7 1 9 2
51 7 13 7 8 8 14 13 0 1 7 15 13 9 9 13 1 15 9 9 0 8 14 13 15 7 13 9 1 9 7 9 9 15 2 1 9 9 0 1 1 9 9 0 1 9 8 8 1 9 0 2
84 7 13 9 9 0 1 9 0 7 15 14 13 0 9 1 9 9 9 1 9 0 2 7 13 1 9 9 1 9 9 9 7 9 9 9 7 9 9 9 1 9 2 15 13 9 0 0 1 9 9 9 9 0 15 13 1 15 9 0 1 9 1 9 1 9 7 9 9 7 9 0 1 9 7 9 9 10 9 7 9 9 1 15 2
10 9 9 9 0 13 9 9 0 1 9
38 9 9 9 0 13 9 9 0 1 9 8 12 9 2 8 2 13 9 0 9 9 9 0 1 9 1 9 9 0 15 13 15 9 1 9 9 0 2
45 7 1 9 9 0 1 9 9 9 1 9 8 0 9 2 13 9 9 0 8 8 15 13 9 9 1 9 0 7 15 13 9 10 9 2 1 9 1 7 8 2 1 9 9 2
25 7 13 9 0 0 8 8 1 2 9 1 9 9 1 9 9 0 1 9 1 0 9 0 2 2
25 7 7 15 14 13 1 15 7 13 9 9 14 13 9 0 1 9 0 13 1 9 0 1 9 2
15 12 9 1 9 8 8 1 9 0 2 9 0 7 0 2
3 12 2 12
64 12 9 1 9 8 8 1 9 0 2 9 0 7 0 2 7 13 9 0 1 8 8 7 15 14 13 9 1 9 9 7 14 13 9 9 15 1 9 0 1 10 9 2 7 13 1 7 15 14 13 3 1 9 0 15 14 13 1 8 8 1 9 0 2
113 7 13 9 1 9 9 1 9 9 0 0 2 7 9 14 13 9 0 0 0 9 1 10 9 1 9 9 1 9 8 2 7 1 15 13 15 7 15 14 13 0 9 8 1 9 2 7 7 9 0 0 1 10 9 14 13 3 1 9 0 2 1 7 14 13 9 0 1 8 8 0 9 9 7 9 1 9 2 2 7 13 9 7 10 9 13 9 0 1 9 0 7 0 1 8 8 2 7 13 9 1 9 9 8 8 7 13 9 1 9 8 8 2
10 8 2 8 1 15 9 1 9 9 0
6 9 12 9 12 2 12
25 13 8 8 9 9 0 1 9 0 8 8 7 8 13 9 1 9 9 0 0 7 0 1 9 2
45 7 13 7 9 9 13 9 1 9 7 7 13 9 8 9 7 15 13 9 1 9 13 1 9 9 8 8 8 0 1 2 8 8 8 7 9 9 9 15 1 9 9 9 2 2
45 7 13 9 9 0 9 7 2 9 9 8 8 8 8 8 8 8 8 9 15 14 13 15 7 7 9 8 8 0 14 13 9 7 9 2 0 1 7 8 14 13 0 1 15 2
92 7 13 8 1 9 0 1 9 2 2 8 8 2 2 0 1 9 9 9 9 7 15 13 10 9 9 7 9 8 13 1 7 15 13 1 9 9 0 9 1 9 0 1 9 0 7 7 3 9 13 15 9 7 9 13 15 9 0 7 7 9 0 0 13 9 9 0 13 9 1 9 1 7 13 1 9 9 7 9 7 13 9 7 9 15 9 9 1 9 9 9 2
25 7 13 7 8 13 9 1 9 9 0 0 7 0 1 9 2 7 3 0 1 9 0 1 9 2
24 7 13 8 1 9 15 1 7 13 9 9 9 7 0 13 1 9 9 9 8 1 9 9 2
96 7 13 9 0 7 9 13 1 15 9 1 9 0 1 0 15 13 1 9 0 7 9 9 9 0 7 9 9 9 1 9 2 7 7 13 9 9 0 7 13 9 0 14 13 1 9 9 9 15 1 9 12 9 12 2 9 10 1 9 2 7 7 15 1 0 9 7 13 9 1 9 1 9 9 9 9 1 9 0 2 7 1 0 3 7 13 9 0 1 9 1 9 1 10 9 2
13 8 13 1 9 1 9 1 9 0 1 9 9 9
6 8 12 9 12 2 12
25 13 9 9 0 8 8 9 9 7 9 15 14 13 9 0 1 9 9 1 9 1 9 9 9 2
61 7 13 8 1 9 0 13 15 1 15 9 9 0 2 8 2 1 8 0 2 8 1 9 1 9 7 9 9 0 7 9 15 1 9 15 7 8 8 1 10 9 2 2 13 9 1 7 8 13 1 9 9 0 8 8 1 9 1 9 0 2
24 7 13 8 7 8 13 1 9 7 9 1 9 0 1 9 9 9 0 1 9 9 9 9 2
29 7 13 7 9 9 9 2 7 15 9 1 9 9 0 15 13 15 9 0 2 14 13 9 9 1 15 0 9 2
28 13 7 9 14 13 1 9 7 13 9 0 0 1 9 9 0 7 13 1 9 9 0 7 9 15 1 8 2
26 7 13 9 9 8 8 8 8 7 9 0 8 8 8 8 9 12 9 0 1 9 9 1 9 9 2
32 13 7 8 13 7 13 9 0 1 9 9 9 1 9 1 8 9 9 0 1 9 8 1 9 9 1 9 0 0 1 9 2
47 0 1 9 7 8 13 0 9 0 1 9 7 9 1 9 7 13 9 9 15 0 1 12 9 1 9 7 13 9 0 1 1 12 1 12 1 9 13 9 9 15 1 9 0 7 8 2
26 15 7 14 13 8 1 15 13 1 12 9 0 1 9 0 1 9 0 1 9 9 15 1 9 9 2
8 9 13 9 0 0 1 9 8
3 9 12 9
43 13 9 0 1 9 9 9 9 7 9 15 13 15 9 0 1 9 8 7 13 9 15 12 9 1 9 7 9 13 9 0 0 1 9 9 0 1 9 8 9 1 9 2
74 7 13 8 8 9 9 0 8 1 9 9 1 9 9 2 7 8 8 13 1 9 8 15 9 1 9 0 1 9 1 7 15 14 13 9 0 7 0 2 2 0 1 7 2 9 13 1 9 0 15 13 15 9 0 7 13 1 9 15 0 1 9 1 9 0 2 7 9 9 9 9 9 2 2
26 7 13 8 9 1 7 15 2 9 0 8 8 9 9 8 8 7 8 8 7 9 9 1 15 2 2
52 7 9 1 9 1 9 9 0 9 8 0 1 9 0 1 15 1 15 9 9 13 8 2 7 9 15 9 0 1 9 1 8 8 2 7 13 7 13 9 1 9 9 8 8 13 9 9 8 8 0 2 2
28 7 13 7 9 8 13 9 9 8 8 0 1 9 9 2 8 8 9 7 9 7 9 9 0 0 9 2 2
48 7 13 2 7 9 13 8 8 9 0 7 9 0 8 1 15 1 9 0 2 2 9 7 2 8 8 13 8 7 14 13 7 13 1 15 1 9 7 15 13 9 1 9 1 10 9 2 2
12 9 0 1 9 0 0 13 1 9 9 1 9
3 9 12 9
45 13 9 0 1 9 9 0 1 9 9 9 1 9 9 9 1 9 1 9 9 1 9 1 9 9 9 0 8 8 1 12 9 0 1 9 15 13 15 9 0 7 0 1 15 2
56 7 13 9 9 9 0 1 7 13 0 9 9 0 1 9 7 9 9 7 0 7 9 7 9 0 1 9 9 1 9 1 9 9 0 0 13 1 9 9 0 13 1 9 9 7 9 7 9 1 9 9 7 9 9 0 2
8 9 0 13 9 9 1 9 0
3 9 12 9
25 13 9 9 9 9 0 1 9 9 1 9 0 7 13 9 7 9 15 0 1 9 15 13 9 2
42 7 7 13 8 1 9 1 9 9 1 9 15 13 15 9 9 0 1 9 9 13 8 13 15 7 3 8 8 1 8 9 0 1 9 13 0 1 9 1 9 9 2
58 7 10 9 7 9 13 9 9 14 13 7 13 9 15 1 15 1 15 9 9 0 8 8 8 8 8 8 7 9 15 13 9 1 9 15 1 7 13 9 1 9 1 9 0 1 9 8 8 9 9 0 8 8 1 12 9 0 2
35 7 13 9 9 9 10 9 7 13 8 1 9 8 8 8 7 15 14 13 8 9 15 9 1 8 7 13 9 1 9 9 1 9 0 2
37 9 7 9 0 1 9 15 13 1 9 1 9 7 9 0 13 9 9 8 9 9 15 13 9 9 8 8 8 8 13 8 8 9 1 9 0 2
39 7 1 9 15 13 9 9 7 9 14 13 8 8 0 7 14 13 15 13 8 8 9 8 0 1 9 12 9 1 9 9 13 1 9 15 8 8 9 2
47 7 9 0 0 15 13 9 13 9 9 15 13 9 15 1 9 15 2 7 1 9 8 9 0 8 9 9 13 1 9 1 9 9 1 9 15 15 14 13 10 9 0 1 9 9 15 2
13 9 0 0 13 9 2 9 9 0 7 0 0 2
3 9 12 9
23 13 9 9 0 8 1 9 8 8 3 9 9 1 9 9 2 9 0 7 0 0 2 2
58 7 13 8 1 9 0 13 15 1 9 9 1 9 9 0 8 8 2 7 8 8 8 8 7 9 13 1 9 9 0 7 0 0 8 8 9 0 8 8 13 1 15 0 9 1 9 8 8 7 13 1 15 9 8 1 9 2 2
28 7 13 9 15 13 9 0 9 1 9 1 7 15 2 9 0 9 14 13 1 15 9 0 9 0 9 2 2
51 7 13 2 7 15 7 13 9 7 9 0 0 7 14 8 1 9 9 0 1 9 9 8 8 7 8 1 9 1 9 9 7 7 8 1 9 1 9 1 8 7 8 7 8 7 9 0 8 8 2 2
21 7 13 9 1 2 7 0 15 9 0 7 4 9 1 9 9 9 0 0 2 2
34 7 13 9 0 0 1 9 7 0 9 9 1 9 1 9 0 2 0 1 9 15 2 1 9 9 1 9 0 7 0 7 0 2 2
36 7 13 9 1 7 13 3 9 0 1 9 0 1 9 9 1 9 0 2 0 1 2 9 9 9 9 1 9 9 9 15 13 1 9 2 2
26 7 1 9 0 13 9 0 0 7 15 14 13 1 9 1 8 1 9 0 1 9 9 15 0 0 2
42 7 13 8 2 7 15 1 9 1 9 9 8 1 9 9 1 9 0 1 9 9 0 14 7 8 13 9 8 0 8 8 7 13 7 13 8 8 0 1 9 2 2
7 8 13 9 12 12 8 0
3 8 12 9
42 13 9 8 8 0 0 0 0 9 7 9 0 14 13 9 0 1 12 12 8 0 13 0 1 9 8 1 9 8 0 1 9 9 9 8 8 9 9 1 9 0 2
49 7 13 1 8 8 0 8 8 9 8 8 9 9 9 15 7 15 13 9 9 8 8 9 9 15 13 1 9 8 13 15 9 1 9 15 1 8 2 8 8 8 8 0 1 9 1 9 0 2
23 7 13 8 3 7 2 3 9 8 8 9 9 0 1 8 1 9 9 7 12 9 2 2
33 13 8 9 13 9 1 9 0 1 9 9 7 9 1 9 0 7 9 1 9 8 9 8 8 9 1 9 9 0 1 9 9 2
20 7 13 9 8 8 8 9 8 0 7 12 8 14 13 1 9 1 9 9 2
38 13 9 14 13 9 8 8 8 8 8 0 1 3 15 14 13 9 9 9 1 15 7 1 9 8 8 8 8 8 13 1 15 0 1 12 12 0 2
13 7 13 9 3 9 9 8 8 8 1 9 8 2
26 14 7 9 13 7 9 9 9 9 0 2 7 15 15 13 15 9 9 0 7 9 0 8 8 0 2
23 7 7 8 13 7 15 14 13 9 9 9 0 1 9 1 8 1 9 1 9 9 9 2
34 7 14 13 8 8 1 9 9 1 9 12 12 9 1 8 1 9 9 9 9 7 9 9 12 12 12 8 0 1 8 1 9 9 2
15 9 0 2 9 9 0 1 8 0 13 7 13 8 8 0
66 9 0 2 9 9 0 1 8 0 13 7 13 8 8 0 11 12 9 2 8 2 13 9 8 8 9 9 7 9 7 9 0 0 3 9 7 9 0 1 8 0 14 13 9 15 0 1 1 9 0 1 9 0 7 9 7 9 7 8 1 9 9 9 8 8 2
55 7 13 9 0 15 13 9 9 0 7 9 0 1 9 8 0 15 7 15 14 13 9 1 9 0 1 9 7 7 10 9 13 9 15 1 9 7 9 0 0 1 7 15 14 9 1 8 0 1 9 1 9 9 0 2
72 7 13 9 0 15 13 13 1 9 1 9 8 1 9 7 9 15 13 1 9 9 9 0 1 11 1 7 9 8 0 13 7 9 8 8 8 9 0 1 9 9 1 0 0 7 9 15 0 9 1 9 0 15 14 13 9 9 8 0 7 9 0 1 9 1 1 9 1 9 8 0 2
64 7 13 1 9 9 9 1 0 7 13 9 9 7 9 3 1 9 0 7 9 15 0 1 7 13 1 9 7 13 15 1 9 9 9 9 1 10 9 1 7 9 9 9 1 9 7 9 15 0 1 9 0 1 9 13 9 0 1 9 9 0 1 0 2
46 7 1 9 15 13 1 8 0 7 9 13 9 0 7 15 9 0 7 7 15 14 13 1 9 0 8 8 7 7 13 9 9 0 7 0 7 9 15 0 10 9 1 7 15 0 2
41 7 13 1 7 9 9 0 1 9 0 7 13 8 0 1 9 9 0 7 0 7 13 1 15 9 7 9 0 0 1 9 15 1 9 9 0 15 13 15 9 2
44 7 1 9 9 0 1 8 0 8 8 13 8 7 8 0 7 9 9 13 8 8 8 8 0 0 1 9 0 2 7 13 9 9 0 8 8 1 9 0 1 12 12 9 2
52 7 13 9 0 7 9 15 0 0 9 0 1 9 9 7 7 9 13 9 0 1 9 0 1 8 0 0 7 9 15 13 1 9 1 9 0 1 9 0 4 3 1 9 9 7 7 3 1 9 1 9 2
9 8 9 1 9 9 8 9 1 9
4 9 0 12 9
23 13 9 0 7 8 9 1 9 9 13 9 9 8 8 9 0 0 1 12 9 1 9 2
39 8 8 8 13 8 9 15 13 1 9 9 2 2 13 9 0 7 8 1 9 9 9 0 7 9 15 13 1 9 1 9 15 9 2 1 9 9 9 2
38 2 13 9 0 7 8 8 8 8 1 9 9 2 13 3 1 9 2 9 2 2 9 1 9 0 2 7 13 1 0 0 1 9 8 8 1 9 2
50 2 13 9 9 1 9 2 9 9 0 2 1 9 1 9 0 1 9 9 2 7 9 9 2 7 9 9 0 2 7 9 9 0 0 2 7 13 9 9 0 1 9 9 7 9 0 1 10 9 2
24 2 13 9 9 2 8 1 9 9 2 2 7 1 9 1 9 0 8 7 1 9 9 0 2
45 2 13 9 9 9 9 0 0 2 13 1 15 9 1 9 0 2 7 9 9 0 2 7 9 0 2 7 13 1 9 9 15 9 0 0 13 15 9 0 2 1 9 9 9 2
3 2 13 2
9 8 8 8 1 9 8 8 12 9
3 8 12 9
42 13 12 9 0 8 8 7 13 8 1 8 9 9 1 15 13 8 8 13 8 2 7 15 1 9 8 2 12 8 8 1 9 9 2 9 1 15 13 15 9 8 2
20 7 13 9 7 9 0 13 1 7 9 9 13 9 7 13 1 9 9 0 2
32 7 13 8 9 8 13 9 9 9 15 7 15 13 7 9 13 8 8 9 1 7 13 1 9 9 1 9 1 9 8 0 2
6 0 9 8 13 1 9
3 8 12 9
29 13 9 0 3 7 15 1 0 7 13 8 8 0 9 8 8 1 8 3 9 9 0 1 8 1 9 9 3 2
54 13 7 8 12 9 2 0 9 9 8 9 8 8 8 2 13 1 15 9 9 8 8 8 1 8 2 7 14 13 1 8 8 0 0 1 8 1 9 8 0 0 1 9 8 0 15 13 1 15 9 1 9 9 2
28 13 0 9 14 13 1 8 1 9 9 2 1 9 9 9 12 9 9 9 9 1 9 15 13 1 9 0 2
39 7 13 9 0 7 15 13 9 1 9 2 1 7 9 8 8 13 1 9 0 1 9 2 7 7 15 1 9 1 9 7 9 1 9 9 0 1 8 2
12 8 8 13 0 9 1 9 8 1 9 9 0
3 8 12 9
45 13 9 9 9 0 9 9 7 9 9 1 9 0 0 0 2 8 2 1 8 8 13 9 12 7 12 1 12 1 9 1 9 9 15 13 9 1 15 1 9 9 0 1 9 2
61 7 13 8 8 9 9 9 9 8 0 1 9 9 7 15 1 9 8 13 9 0 1 8 7 8 0 8 8 1 0 9 1 10 9 1 9 0 2 7 13 7 15 13 9 12 1 12 1 9 9 8 1 9 0 1 9 12 0 9 15 2
26 7 13 1 7 9 9 8 1 12 9 1 15 8 8 8 13 1 9 9 1 9 15 13 1 15 2
