705 17
18 0 3 15 13 16 13 12 9 15 7 3 15 9 15 13 13 1 9
28 15 3 13 15 3 13 15 3 7 9 16 9 13 0 7 9 16 9 13 9 15 7 11 16 9 13 0 9
13 7 16 15 13 15 1 9 9 12 13 1 15 12
8 16 3 13 13 15 15 9 13
3 13 9 15
5 3 13 15 3 15
12 16 3 13 9 9 15 13 3 15 9 15 0
9 3 3 13 9 15 3 3 9 15
17 3 13 15 9 15 15 13 7 15 13 7 9 15 1 15 13 15
18 16 3 9 0 3 13 7 3 1 9 13 9 3 13 3 3 15 0
4 13 9 9 15
3 13 7 13
9 3 0 9 7 0 9 13 1 9
13 3 13 9 0 9 0 13 7 9 0 9 0 13
20 0 3 15 13 9 15 0 7 13 15 13 15 9 0 15 13 9 15 1 9
11 13 3 15 1 9 1 9 15 13 9 0
17 15 3 13 7 13 13 15 9 7 13 9 15 13 11 1 9 15
6 7 13 0 13 7 13
4 7 13 11 9
23 3 3 13 13 1 15 0 0 7 13 9 9 7 15 0 13 16 13 15 13 9 11 13
9 9 13 15 3 13 7 13 9 15
3 7 13 15
9 13 3 3 1 15 9 9 0 13
11 7 13 1 9 11 13 7 13 1 15 9
11 15 3 13 0 13 13 15 9 15 7 13
20 7 13 15 13 1 9 7 6 0 9 7 9 13 13 1 11 7 1 9 15
14 1 15 15 7 9 13 15 3 7 9 15 3 13 15
13 3 13 15 1 15 6 9 13 13 15 15 13 16
7 7 13 13 9 1 9 0
13 13 3 15 1 9 13 1 15 9 7 13 15 11
8 0 3 13 6 13 9 0 0
6 9 3 0 7 9 3
9 13 3 13 13 16 13 15 9 0
14 1 15 3 9 7 1 9 13 13 15 1 15 0 13
4 13 3 1 9
10 3 3 13 15 1 9 0 13 1 0
11 7 3 13 15 13 9 7 9 3 13 13
8 3 13 16 13 13 9 1 9
11 7 13 3 13 11 13 12 1 12 9 15
5 15 13 13 1 9
7 0 3 13 1 15 13 13
12 0 13 9 13 1 9 15 13 9 15 7 13
6 6 15 11 6 15 11
8 6 9 16 3 13 9 1 15
10 6 9 15 13 15 3 13 13 1 9
8 7 6 9 13 3 9 13 0
7 7 13 15 0 3 3 0
15 9 13 3 13 7 9 13 15 3 13 16 13 1 9 9
10 7 16 9 9 13 1 15 13 15 13
11 7 15 3 13 9 1 9 0 13 15 15
8 3 13 15 1 9 7 9 13
6 7 13 13 0 13 13
6 6 9 15 7 9 15
11 7 0 13 1 9 7 13 9 7 13 15
11 7 15 3 13 3 15 13 13 15 1 15
17 0 15 13 9 9 7 3 13 13 3 9 7 13 13 1 9 15
14 13 3 9 13 9 15 7 13 9 1 9 9 7 13
3 0 3 13
16 0 13 9 0 9 15 13 9 13 1 9 12 9 16 13 15
5 7 9 13 15 9
13 3 0 13 9 0 9 13 1 9 15 13 9 13
3 13 15 11
6 3 0 3 13 0 9
12 1 9 0 13 11 9 9 0 7 13 9 15
14 0 3 13 9 15 13 15 13 3 1 9 9 11 9
3 0 13 9
4 13 15 15 3
12 1 0 3 9 9 13 1 15 11 13 1 9
3 0 3 13
7 7 13 15 1 9 13 9
5 0 3 13 13 15
18 13 15 15 9 0 9 15 7 9 13 15 7 9 15 3 13 1 15
2 13 15
12 1 9 3 13 9 0 9 9 9 9 9 9
7 13 15 16 13 1 9 15
5 3 13 11 13 15
14 13 1 9 16 3 12 9 13 15 7 3 13 15 13
13 7 13 15 7 13 15 7 13 9 9 12 9 0
3 9 0 0
4 0 3 13 13
12 13 15 3 1 9 0 7 1 9 0 7 0
5 13 3 11 11 13
8 7 13 15 11 13 13 15 13
9 7 15 13 9 15 15 1 13 15
6 9 0 13 15 3 13
10 13 3 9 15 3 13 15 3 11 12
9 3 13 9 16 1 11 9 13 15
14 7 13 15 11 7 13 1 15 9 7 13 9 0 9
5 7 15 0 13 15
5 15 15 15 13 11
8 1 0 9 13 9 1 11 13
5 9 3 13 13 9
4 15 15 15 13
3 6 13 15
18 0 1 13 15 13 9 0 9 9 15 13 13 15 1 9 1 9 15
7 13 1 15 7 15 13 15
10 7 1 15 13 9 0 7 13 15 3
8 15 3 9 13 9 3 3 13
4 0 3 13 15
7 7 13 1 15 9 13 3
4 11 3 13 15
6 11 3 13 1 9 15
4 15 3 13 15
6 13 3 15 1 9 15
2 13 15
6 13 3 13 1 9 13
7 3 13 0 0 7 0 0
18 13 16 13 0 9 15 12 1 0 15 7 12 1 0 15 1 9 15
13 7 10 13 1 0 7 1 0 15 13 15 0 13
10 7 13 15 1 11 1 15 13 9 0
6 9 16 13 15 15 9
3 13 9 0
4 9 3 13 16
4 11 3 13 15
4 3 3 13 9
10 9 0 3 13 1 9 3 7 1 9
5 15 3 15 13 15
4 0 3 13 13
7 9 3 7 9 13 15 9
8 9 3 3 13 9 13 1 15
6 13 3 13 3 1 9
5 3 13 15 9 13
4 9 3 0 13
12 13 15 9 7 9 13 15 7 13 1 9 0
8 0 3 13 13 9 9 7 3
3 3 13 15
8 1 9 3 15 1 12 13 9
17 9 3 13 16 13 9 13 15 3 7 13 1 15 9 13 15 13
6 15 15 15 13 1 11
7 7 15 3 13 13 15 9
9 15 3 9 15 13 16 13 13 9
9 7 13 15 9 16 9 15 12 13
5 6 15 9 0 13
11 13 15 3 9 13 15 15 7 13 1 15
9 3 3 15 3 3 13 15 9 0
25 3 13 1 15 0 9 0 13 1 9 1 9 11 0 1 9 11 9 0 15 13 1 9 7 9
5 0 3 13 13 15
7 0 3 13 1 9 15 13
5 15 3 0 9 9
12 13 3 15 16 3 13 9 15 9 7 1 9
3 3 13 9
12 6 13 15 16 3 13 9 0 16 15 0 13
7 12 13 15 7 12 13 15
14 3 13 15 9 0 12 9 15 13 9 15 13 3 9
3 0 13 0
3 6 13 15
6 9 12 9 15 13 13
4 13 15 9 15
15 0 9 7 0 13 16 13 3 3 13 7 13 3 3 13
7 3 13 9 13 1 0 15
5 3 13 15 9 13
7 3 13 7 13 1 0 15
4 3 13 15 13
23 11 3 13 1 11 1 9 11 0 13 1 15 9 13 9 9 0 7 13 1 9 15 13
12 13 3 0 9 0 1 9 15 1 9 15 13
3 0 3 13
9 7 13 3 13 13 15 12 15 15
2 13 15
4 13 1 15 15
5 13 3 11 13 15
7 13 3 16 13 13 15 3
9 3 3 3 13 12 9 13 1 15
3 7 13 15
2 13 15
6 13 9 15 1 15 9
14 0 3 13 11 13 1 11 9 3 9 7 9 13 15
3 11 3 13
4 15 3 13 9
6 11 3 3 13 1 9
8 3 1 0 3 13 13 13 11
15 9 3 13 9 13 15 9 7 9 0 1 11 16 13 15
10 0 13 13 15 1 9 16 9 9 13
4 11 3 13 15
12 15 13 1 12 13 15 11 3 7 11 13 11
1 11
18 13 3 11 16 15 3 13 7 3 9 13 13 9 13 9 1 9 13
4 13 15 9 0
4 0 13 9 0
3 13 1 9
8 9 15 9 15 3 15 13 13
17 9 3 7 15 13 1 15 13 11 13 9 7 13 13 15 3 13
16 1 0 3 9 15 13 1 9 13 15 9 7 9 1 11 13
3 13 3 13
6 13 3 16 11 13 13
14 7 13 3 1 9 1 9 7 9 0 13 13 9 15
4 7 13 15 9
6 7 13 11 13 15 13
12 13 11 13 1 9 7 13 9 9 1 9 9
5 7 13 9 1 9
4 7 13 15 11
10 7 13 1 9 9 0 9 7 13 13
12 7 13 15 9 0 7 13 9 0 13 1 15
13 3 3 13 3 13 9 13 1 15 15 0 7 0
12 7 13 13 1 9 15 1 15 11 7 9 13
4 15 15 3 13
12 13 3 15 1 9 3 13 7 13 1 9 15
13 7 13 1 15 16 13 15 15 7 13 9 13 16
3 13 3 0
4 7 13 15 11
17 7 13 13 15 11 1 9 1 9 7 13 9 15 9 13 13 9
12 7 13 3 1 9 7 13 3 9 0 9 13
2 7 13
13 7 13 1 9 7 13 15 15 13 7 13 1 15
16 7 9 13 1 11 13 16 11 13 7 16 1 9 9 13 9
6 3 13 16 9 0 13
15 15 3 3 13 9 0 0 9 15 7 9 15 7 9 13
10 9 3 13 13 7 16 3 13 9 13
3 7 13 15
24 7 0 13 13 1 0 9 15 13 9 7 13 15 7 13 15 1 12 12 7 12 12 7 12
7 15 3 3 13 13 15 15
35 3 0 9 15 3 13 13 1 9 0 15 9 0 7 3 13 13 13 7 13 0 15 9 7 13 9 0 16 13 1 9 15 9 0 13
8 7 13 15 1 9 1 9 13
4 15 3 0 13
3 3 13 15
6 7 13 15 15 9 13
8 11 3 3 13 15 7 13 15
43 7 9 15 13 1 9 9 9 12 1 12 7 3 13 1 0 9 7 13 15 15 7 3 12 9 13 7 3 1 0 13 13 1 11 13 1 9 1 3 13 15 9 15
6 7 13 15 13 13 0
8 11 3 3 13 9 13 13 9
7 7 13 1 9 9 13 15
13 7 13 9 13 1 9 13 7 0 13 13 15 13
6 7 13 15 1 9 15
26 7 13 9 11 9 0 3 13 9 15 7 13 16 11 13 13 1 0 7 0 1 9 13 15 1 15
24 11 3 13 15 11 13 15 9 0 7 0 7 13 15 7 13 15 3 13 7 1 9 15 13
9 7 13 3 1 9 1 9 13 13
10 13 15 0 1 0 9 12 7 13 3
5 0 3 13 13 15
11 7 13 15 13 15 9 1 9 1 9 0
22 7 13 15 13 1 9 13 3 0 9 15 7 1 0 9 0 13 1 15 1 9 13
9 7 13 1 15 1 9 7 13 9
39 9 3 7 15 9 16 3 13 9 13 3 13 13 9 9 7 1 9 16 3 13 15 3 13 7 15 0 13 15 13 13 9 9 7 9 7 9 7 9
9 3 13 15 9 0 16 9 15 13
11 15 13 15 1 9 13 1 15 13 13 15
8 15 0 0 3 13 7 13 9
9 3 3 9 1 9 13 1 9 0
15 7 3 13 15 9 15 7 13 15 9 9 15 7 13 3
6 0 3 15 3 13 13
5 7 13 3 9 3
5 15 9 0 9 13
3 9 3 13
3 0 3 13
5 9 3 9 13 13
4 7 0 13 15
14 13 1 15 9 16 3 13 15 13 0 7 15 13 0
41 7 1 12 9 13 11 11 7 11 7 11 7 13 15 1 9 0 12 7 13 15 1 15 7 13 9 15 13 15 0 3 3 9 15 3 13 9 1 9 3 13
12 7 3 13 15 3 13 3 7 11 12 1 15
16 7 13 15 16 11 13 7 13 15 15 13 3 13 13 1 15
5 0 3 13 15 13
2 1 9
17 0 7 0 9 15 15 13 13 1 15 7 1 0 3 13 1 15
25 13 3 9 15 7 13 15 16 9 0 13 13 1 9 0 7 13 15 7 13 13 1 0 9 13
11 15 3 12 0 9 13 1 9 15 15 13
27 7 15 3 13 12 1 0 0 13 1 15 0 15 13 3 16 13 9 0 1 9 15 7 13 15 1 9
9 16 3 3 9 3 0 13 15 13
11 7 1 9 9 9 7 9 13 15 13 9
4 9 3 13 13
8 9 0 15 13 16 9 0 13
2 3 13
6 7 13 11 13 9 15
7 1 9 3 0 7 1 9
32 6 13 1 11 7 9 0 13 13 9 7 9 7 13 15 1 9 7 13 15 9 7 13 15 15 7 13 15 7 0 9 13
15 13 3 13 9 15 15 13 7 9 15 15 13 15 13 15
13 13 16 13 15 13 9 13 15 7 0 15 13 15
4 0 3 3 13
5 15 13 16 13 15
3 13 15 13
8 7 13 7 1 9 13 13 13
5 7 13 11 13 15
12 13 3 15 15 16 15 9 13 15 1 9 15
4 0 1 13 15
16 13 3 15 15 12 9 7 13 15 7 13 15 15 9 0 13
2 3 13
6 15 0 0 13 0 13
5 15 3 13 9 9
14 7 13 1 15 15 1 9 7 9 16 15 13 13 9
6 0 3 13 7 13 15
4 13 3 12 9
11 3 0 3 1 13 3 13 9 7 9 0
4 0 9 13 15
13 3 9 1 9 13 16 12 13 7 13 15 1 15
11 13 1 0 15 16 13 9 15 9 9 15
6 7 13 9 15 13 15
15 13 15 3 0 13 7 15 13 9 3 13 13 15 15 0
5 13 3 15 1 9
8 6 3 0 7 13 1 0 9
30 7 1 0 9 1 9 0 9 13 15 7 9 3 13 9 15 7 9 13 13 1 9 7 9 15 13 1 9 13 15
5 13 15 7 13 15
2 13 3
3 11 3 13
14 11 0 12 1 12 1 12 13 1 9 16 15 13 15
8 7 3 3 13 13 9 9 16
12 0 3 13 13 7 13 7 13 15 12 1 15
8 7 13 15 13 11 9 13 13
5 7 13 15 11 16
16 15 3 1 0 9 3 16 3 9 3 13 12 9 13 15 15
19 7 13 3 13 1 9 7 13 15 16 16 0 13 13 1 15 9 7 13
8 7 3 13 13 15 0 9 13
1 13
3 7 13 15
8 0 3 13 9 0 13 1 15
4 3 13 3 15
4 15 3 13 9
5 0 3 13 15 13
5 7 9 15 13 15
5 0 3 13 13 15
13 13 3 13 11 1 15 9 13 15 1 9 9 13
2 13 15
4 13 15 9 0
7 13 3 9 0 7 13 15
6 3 13 1 15 13 15
13 13 3 15 13 9 9 7 13 1 9 13 15 13
5 13 9 16 3 13
4 13 3 0 3
10 13 9 15 7 11 16 13 15 1 11
5 3 0 3 9 13
1 6
21 3 13 15 11 16 13 13 9 15 7 9 15 11 13 9 15 7 13 9 15 11
24 7 6 13 13 7 3 13 13 1 15 9 13 0 16 3 13 9 15 15 13 15 1 9 15
6 7 13 1 15 9 13
13 7 6 13 1 9 7 13 9 7 13 9 15 11
3 13 3 11
11 7 3 0 15 16 13 9 9 15 1 15
4 13 9 9 15
5 7 13 9 15 13
26 7 13 1 15 9 13 3 15 7 1 15 9 0 13 13 15 9 0 7 13 15 13 1 9 15 13
8 0 9 0 13 13 11 7 11
4 7 0 15 9
10 11 3 13 15 9 0 13 1 9 15
12 7 13 11 7 9 15 13 15 1 13 1 15
16 9 3 13 7 13 15 9 13 15 9 7 9 0 13 1 15
4 7 13 1 15
4 9 13 1 9
3 9 13 11
6 13 3 3 9 13 15
19 13 3 9 7 13 15 1 9 15 1 11 3 0 13 11 13 11 15 13
91 7 0 13 11 16 12 12 9 13 9 13 16 13 13 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0
18 15 13 9 0 15 7 9 15 16 15 13 13 7 15 3 13 13 15
8 7 13 11 13 15 16 13 13
19 13 15 13 13 9 13 9 9 7 0 9 13 13 1 9 13 9 0 0
4 9 13 15 0
13 7 13 11 1 11 1 9 0 7 13 13 1 9
1 13
5 3 3 13 13 15
13 3 0 9 13 15 13 9 0 16 1 0 13 13
6 1 9 3 15 13 9
4 3 9 13 13
7 7 0 13 15 15 3 13
7 7 13 13 9 7 9 13
10 13 7 13 9 15 7 13 1 9 15
12 7 13 9 0 9 7 15 15 13 1 15 13
12 3 13 9 0 16 9 13 1 15 13 13 15
2 13 3
10 7 13 9 3 7 9 0 15 13 0
7 7 13 1 15 15 13 15
9 7 0 13 9 15 1 9 15 13
6 6 15 13 16 13 15
14 13 15 1 9 13 0 7 13 15 9 3 9 3 13
13 3 13 9 15 7 13 7 1 9 13 15 3 13
4 13 3 9 15
8 0 3 9 1 9 15 13 15
18 7 13 7 3 13 0 13 9 13 9 1 9 1 9 15 13 15 9
5 11 3 13 1 15
7 7 9 15 13 0 7 13
3 3 13 15
8 7 13 11 9 15 1 15 0
10 7 0 13 15 3 3 13 15 1 15
3 6 13 15
10 15 3 13 9 9 0 7 15 13 0
7 7 13 15 9 1 9 15
2 9 13
7 7 13 15 1 9 13 11
8 13 15 15 9 0 16 13 3
58 13 3 1 0 7 0 13 1 9 7 9 13 7 13 9 0 7 12 1 12 1 15 7 9 15 15 13 13 1 9 0 7 9 11 13 9 1 15 13 12 9 7 11 9 0 9 0 7 11 7 15 0 15 13 15 1 9 15
6 13 3 15 9 15 13
22 7 13 1 9 0 13 13 7 1 9 7 9 0 13 13 15 7 3 1 9 9 13
6 0 3 13 13 1 15
2 9 13
31 13 3 15 1 9 13 15 9 15 1 9 15 13 9 1 9 0 7 1 9 3 13 15 7 1 9 3 13 7 1 9
4 15 15 9 13
9 13 3 15 3 13 3 13 15 13
15 7 6 13 9 1 11 15 13 9 11 7 0 9 9 13
5 15 13 13 15 15
10 3 15 13 13 12 1 9 13 15 16
3 0 3 13
30 13 3 11 12 1 12 13 15 9 7 9 1 15 9 7 9 13 7 13 15 13 9 0 7 13 13 7 13 1 15
9 15 3 13 0 1 15 15 13 0
4 13 15 15 13
15 7 13 3 13 15 12 1 15 13 9 15 7 13 15 13
4 13 3 1 15
14 7 13 3 13 15 9 9 15 15 7 9 15 13 15
2 0 13
4 13 3 11 13
6 0 3 3 13 9 0
2 3 13
5 7 13 1 15 9
4 13 3 15 11
4 13 3 1 15
7 16 3 3 1 15 13 15
13 13 3 15 16 9 3 13 1 0 9 3 9 0
3 13 3 15
28 15 15 13 13 1 9 15 7 15 3 13 15 13 9 3 9 7 15 13 9 3 9 7 15 3 13 9 13
4 0 3 13 13
12 1 9 3 9 15 13 9 0 7 13 15 13
4 13 9 1 15
6 13 3 15 16 15 13
5 3 13 15 9 15
7 9 13 15 1 9 12 9
5 13 7 13 15 15
6 13 3 9 13 13 0
12 16 3 15 1 11 13 9 9 15 1 15 13
19 3 13 7 13 0 0 12 9 7 13 13 3 7 13 0 9 0 0 0
12 9 0 13 1 9 1 9 9 0 7 13 15
22 16 3 9 15 15 0 13 3 13 9 12 0 13 0 15 3 6 3 9 9 13 15
8 0 3 13 13 7 0 3 13
6 0 1 7 9 0 13
14 15 3 13 13 15 3 13 15 7 0 15 3 13 15
9 7 3 12 1 15 13 13 1 9
20 3 3 13 15 1 9 7 9 7 9 3 13 15 3 7 15 13 7 15 13
6 9 15 0 13 15 9
1 13
4 13 1 9 15
5 3 13 15 7 13
18 13 15 9 3 13 9 3 13 1 9 3 9 3 13 15 7 9 13
14 3 15 3 13 0 16 1 15 9 3 13 9 0 13
10 3 13 3 13 3 0 9 13 13 3
4 13 3 3 9
5 7 13 11 13 15
9 7 13 13 9 1 15 7 3 13
10 13 3 13 11 1 15 1 9 1 9
6 13 1 15 9 7 13
2 3 13
17 3 3 13 9 9 7 13 9 7 13 3 13 7 13 1 9 13
6 13 1 15 15 9 9
19 3 13 15 3 7 3 7 1 0 9 13 16 3 0 13 9 13 3 11
3 0 3 13
16 7 3 13 13 13 13 1 0 9 16 3 13 13 15 13 15
7 0 15 13 9 1 9 0
3 7 0 13
17 13 3 1 9 7 9 9 7 0 7 0 7 0 7 0 13 3
16 7 15 3 13 9 15 7 1 9 15 13 3 13 13 15 9
3 3 13 15
22 7 15 9 13 12 9 16 13 9 12 3 13 3 9 7 13 9 7 13 3 16 13
20 7 3 1 0 9 13 15 0 9 13 1 9 3 7 3 13 9 15 13 3
7 9 13 1 9 7 1 15
16 13 9 0 7 13 15 7 13 9 1 9 15 7 9 1 9
7 13 3 15 7 3 13 13
17 9 15 13 0 15 13 9 7 0 13 13 1 15 3 13 9 15
15 13 15 13 16 3 13 13 1 9 9 13 15 1 9 15
5 15 3 15 0 13
17 0 1 0 3 1 0 0 13 7 0 1 0 3 1 0 0 13
5 9 3 13 9 15
11 13 3 13 0 7 13 13 9 1 9 0
27 7 1 15 0 1 15 7 15 9 0 13 15 16 3 13 13 3 1 15 3 13 7 15 3 1 15 13
15 16 11 7 9 3 13 3 16 15 1 0 13 3 13 9
3 13 15 9
8 3 13 9 9 0 16 13 13
6 7 13 13 15 13 15
13 13 3 13 1 9 3 13 9 0 13 15 7 13
2 3 11
1 13
5 12 13 7 0 13
16 13 3 7 9 1 15 3 13 3 13 15 7 3 13 15 13
19 7 9 3 13 3 13 9 13 15 13 1 15 9 7 9 7 13 1 15
5 9 13 9 15 13
5 11 3 13 15 13
6 15 13 0 3 12 9
6 13 3 0 11 13 15
5 3 15 13 13 13
13 6 13 1 11 7 13 15 15 13 9 1 9 0
6 7 13 13 15 16 13
1 13
4 7 13 1 15
8 13 3 9 0 13 7 13 13
23 7 13 3 15 13 13 9 7 13 16 13 15 9 0 15 13 9 16 13 15 9 13 13
4 7 0 13 13
3 7 13 13
18 13 1 0 9 1 15 13 13 9 13 1 15 15 3 1 9 3 13
7 13 3 15 13 9 1 9
13 3 13 13 1 9 0 15 3 15 15 1 9 15
6 7 3 13 15 13 15
5 1 15 3 13 15
13 7 1 9 13 1 9 9 16 1 9 9 13 15
5 3 0 13 13 15
3 3 3 13
4 7 13 15 13
5 0 3 13 1 15
7 1 9 3 15 15 13 9
5 15 3 0 0 13
10 11 15 3 9 13 3 3 15 13 9
20 15 3 0 1 9 15 13 1 9 0 7 0 1 9 15 15 9 15 13 13
6 15 13 7 9 13 15
6 13 3 15 15 1 9
32 13 3 9 0 1 9 7 9 1 9 0 7 13 1 9 9 7 13 13 1 9 15 7 11 13 13 9 16 13 15 9 9
12 6 13 15 16 3 13 13 9 10 16 15 13
13 13 3 9 1 11 13 11 13 1 9 12 1 12
12 6 13 15 1 9 13 15 9 1 9 9 13
4 7 13 1 15
5 0 13 1 15 9
15 15 3 3 3 7 0 15 3 13 3 0 7 0 3 13
8 7 15 3 13 15 13 9 15
1 15
4 0 3 13 15
8 3 3 15 9 7 15 3 13
6 0 3 13 9 13 15
7 7 13 1 9 15 13 15
5 3 0 13 1 15
3 3 9 13
4 13 3 15 13
3 13 3 15
15 0 13 13 9 15 7 13 13 9 9 13 15 11 9 13
7 11 3 13 11 0 13 3
7 13 15 9 0 3 13 9
13 15 13 1 15 9 13 1 9 7 9 13 1 9
15 0 3 13 9 0 13 15 1 9 7 13 9 15 7 0
4 3 13 13 9
6 3 13 3 15 15 13
4 0 13 9 0
8 13 15 9 3 13 1 9 15
7 13 3 9 13 13 9 13
7 13 3 15 13 9 7 9
15 13 9 0 13 13 1 9 9 9 13 13 7 0 9 13
11 15 13 9 0 1 15 13 15 1 15 13
13 7 3 1 15 0 0 6 9 13 3 3 0 13
4 7 13 15 13
15 7 0 13 15 13 1 9 7 16 15 13 15 1 9 9
3 15 13 13
3 0 13 15
13 7 13 3 13 15 13 1 15 7 13 15 1 9
9 1 9 3 15 13 15 15 3 13
7 13 9 13 3 9 1 9
12 13 3 15 11 7 13 15 1 15 13 13 15
6 13 0 3 9 15 11
3 13 1 15
4 7 13 1 15
5 13 11 7 13 15
3 9 3 13
5 7 13 15 1 9
10 7 1 13 9 0 7 13 11 1 11
8 13 9 0 7 12 9 13 15
5 0 13 1 15 9
11 3 13 3 1 9 13 9 15 7 13 15
5 13 11 7 13 15
21 3 3 9 13 9 16 9 15 0 13 16 0 13 1 15 3 13 7 13 9 0
17 1 0 13 11 7 9 15 1 0 9 7 3 13 1 15 7 13
8 13 15 11 7 13 13 1 15
7 15 3 13 9 9 0 13
10 11 3 13 15 1 9 13 3 1 9
5 13 11 7 13 15
8 0 13 1 9 0 13 15 3
3 13 15 11
3 13 15 11
6 3 0 13 13 15 15
8 13 3 1 9 7 13 1 15
12 3 15 3 13 16 3 12 9 13 7 9 13
13 3 3 13 9 1 15 13 15 16 13 13 1 15
6 3 0 3 13 1 9
4 13 1 15 11
4 9 15 0 13
4 13 3 0 13
4 13 3 9 13
8 11 3 13 15 9 13 1 9
23 0 3 1 13 3 9 15 13 16 3 3 13 9 7 3 9 15 13 9 0 15 13 9
27 6 6 13 15 16 13 9 15 7 9 13 13 15 13 9 0 7 1 9 3 13 7 13 1 9 1 9
8 15 13 1 11 7 13 1 9
10 13 9 16 15 13 1 15 13 9 0
11 16 3 13 9 13 11 9 13 13 3 15
5 0 3 13 13 15
6 13 3 9 0 1 9
20 7 16 3 13 13 9 15 1 9 7 13 1 9 13 1 0 9 9 1 11
14 7 15 13 9 1 11 1 9 3 13 9 9 13 9
4 13 3 1 15
3 13 15 11
10 7 13 15 16 7 13 15 7 3 13
3 1 9 13
3 0 13 9
7 13 3 15 9 1 15 13
14 0 13 9 13 1 9 3 3 13 9 15 9 7 13
4 9 13 15 13
5 3 3 15 13 13
11 0 3 13 13 15 12 13 1 12 1 12
4 13 3 15 11
2 7 13
7 3 0 9 13 3 13 15
4 13 9 7 13
7 3 0 3 13 15 13 13
18 13 3 13 15 7 15 3 13 9 1 15 16 3 3 13 13 9 15
9 3 1 9 0 13 13 7 13 9
5 0 13 1 9 9
5 1 15 3 13 15
4 13 7 13 15
9 7 1 9 15 11 13 0 9 13
6 13 3 15 11 13 15
4 15 13 9 9
4 15 3 13 15
9 0 9 13 11 1 9 13 1 9
4 15 1 0 13
5 9 3 3 13 15
8 13 3 11 1 13 1 15 9
6 0 13 9 9 13 9
3 13 15 11
9 16 9 9 15 13 13 13 15 13
9 15 3 16 9 13 3 13 9 15
9 7 13 9 15 7 15 3 13 15
9 3 15 0 13 9 15 11 15 13
7 7 13 15 7 9 15 13
8 7 13 11 13 9 0 1 9
1 13
5 3 15 15 13 9
2 3 13
7 3 13 9 0 0 9 13
11 13 16 0 13 9 15 7 16 0 15 13
2 0 13
4 3 13 9 15
5 13 9 7 13 15
6 15 13 3 1 9 0
15 1 9 15 1 9 0 13 16 3 13 13 7 13 0 13
14 3 13 9 1 9 0 7 13 3 0 9 13 7 9
4 15 13 9 9
11 7 9 13 16 9 13 7 3 13 1 9
5 13 3 0 1 15
7 13 3 15 9 7 13 15
18 9 15 15 13 15 0 15 13 7 15 3 13 13 15 1 9 9 15
7 13 3 13 1 9 15 16
8 11 3 9 3 13 3 12 3
9 13 3 11 11 7 9 15 7 11
12 16 3 15 13 9 13 15 16 13 9 1 15
14 11 13 7 13 15 15 1 16 9 13 16 3 13 3
5 13 3 11 1 11
6 13 1 15 16 13 13
29 9 3 13 1 15 1 9 7 13 15 13 11 16 3 13 7 13 1 15 13 13 16 13 1 9 16 13 15 3
4 7 13 15 11
5 13 15 9 13 11
13 7 9 1 13 3 13 16 9 13 16 15 15 13
10 13 3 9 7 9 9 1 11 7 13
12 7 13 3 11 7 13 3 1 15 1 9 13
13 13 3 12 1 9 15 11 0 0 15 15 13 13
23 1 0 3 9 9 0 13 1 9 13 16 11 13 1 11 13 9 1 9 7 13 1 15
5 9 3 13 1 15
5 11 3 13 15 13
6 9 13 15 1 9 0
4 13 11 7 13
5 15 0 13 9 0
6 7 9 0 15 13 15
14 15 9 1 9 13 16 0 13 1 15 1 9 3 13
43 7 9 13 9 3 13 1 9 11 0 0 16 15 13 13 11 16 15 13 15 9 1 9 7 16 1 9 13 7 1 9 13 13 1 9 7 13 9 7 13 9 13 15
6 3 13 9 15 1 9
4 13 3 13 15
4 6 6 13 15
13 13 3 15 13 15 13 7 13 15 13 13 7 15
2 13 11
3 13 3 9
13 1 0 13 15 16 15 9 13 16 9 13 1 15
6 9 3 15 1 15 13
3 13 15 11
7 9 13 15 9 7 13 15
11 9 13 15 16 15 1 9 7 9 1 15
8 15 3 13 15 16 1 15 13
5 13 15 11 3 0
4 9 15 13 15
14 7 3 13 9 16 13 9 7 3 13 15 9 3 13
2 15 9
11 0 13 9 15 16 13 15 15 3 13 15
10 16 1 9 13 13 9 3 15 13 13
6 13 15 3 9 15 13
13 7 13 9 16 0 15 13 15 13 15 9 13 9
10 16 3 3 13 15 9 3 13 1 15
10 0 15 13 16 1 15 13 7 13 15
2 1 0
7 3 15 3 3 3 0 13
16 0 3 9 13 15 16 15 15 13 7 13 16 15 1 9 13
12 6 13 9 7 3 13 16 13 15 15 1 15
5 15 13 15 1 9
13 7 15 15 15 13 7 15 15 7 13 15 1 15
4 9 15 9 13
20 7 13 15 9 15 7 13 16 9 15 15 13 13 1 15 13 7 15 1 15
2 15 13
7 16 15 13 3 13 0 13
9 9 3 7 9 7 9 0 13 11
4 13 3 15 9
7 9 15 7 9 13 15 15
6 15 13 16 9 13 15
4 13 3 15 13
15 6 13 15 15 3 16 13 16 1 15 9 3 13 3 12
7 15 3 3 13 1 15 9
2 13 11
4 9 13 3 0
2 13 9
15 0 3 9 0 13 1 9 16 1 13 9 9 3 13 11
4 13 3 1 15
4 9 6 9 15
2 13 15
5 13 1 15 15 13
14 13 3 7 13 1 11 11 7 1 0 9 15 13 11
14 3 3 13 3 0 9 13 3 1 9 7 13 7 13
9 13 9 15 7 3 13 3 13 15
1 9
7 7 13 1 9 7 13 15
6 15 13 9 13 15 15
4 1 0 13 11
22 0 3 13 13 16 9 13 16 11 13 11 9 0 7 16 13 9 0 13 1 9 15
8 9 3 3 13 13 11 1 9
7 13 3 9 15 13 11 11
7 3 0 13 3 13 15 9
2 13 15
3 13 9 15
