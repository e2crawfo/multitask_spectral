11699 17
2 11 2
5 9 1 10 9 2
2 11 2
7 0 9 1 10 11 11 2
28 10 9 4 4 4 13 1 10 9 1 9 0 1 10 9 0 1 9 15 13 2 10 9 1 10 9 2 2
37 13 10 9 1 9 1 15 1 10 9 0 15 13 10 9 2 10 9 4 13 13 10 0 9 1 9 7 1 12 9 10 9 4 13 10 9 2
9 10 9 13 1 10 0 11 11 2
31 13 2 11 1 11 2 2 13 10 9 1 10 9 7 1 10 9 13 9 2 15 13 1 10 9 15 4 13 1 9 2
11 11 11 4 13 1 10 12 1 12 9 2
8 0 10 9 13 9 0 0 2
17 9 1 11 1 10 12 9 1 9 7 1 11 11 1 10 9 2
9 0 9 2 9 0 1 10 9 2
60 4 13 11 11 2 0 1 11 11 2 1 10 9 1 10 12 9 1 9 2 11 11 2 0 2 4 4 3 13 2 2 4 13 10 0 11 11 2 0 3 0 9 1 10 9 1 10 9 9 11 11 2 1 10 9 1 10 9 0 2
37 11 11 1 10 9 1 12 2 3 13 1 12 2 4 13 3 1 9 1 10 9 15 4 13 10 0 9 1 10 0 9 2 10 9 11 11 2
26 13 2 11 11 4 13 2 1 10 11 2 1 10 9 13 1 9 13 10 9 1 10 10 0 9 2
11 2 6 11 2 15 4 13 10 9 2 2
2 11 2
13 9 1 9 1 10 9 13 7 13 1 12 9 2
24 11 2 10 9 4 4 13 1 10 9 1 10 9 7 13 1 9 1 10 9 2 1 11 2
52 9 2 11 11 2 12 9 2 0 2 15 3 3 1 10 12 1 3 9 15 13 1 10 9 1 10 9 11 11 2 12 9 2 9 1 9 1 9 2 1 10 9 1 10 9 3 1 10 9 1 11 2
27 10 9 4 4 13 1 10 9 7 13 1 12 9 13 1 9 2 3 12 9 1 10 11 1 10 11 2
26 1 10 10 9 10 9 4 13 9 1 9 2 1 15 10 12 9 1 10 9 3 4 13 10 9 2
9 9 15 4 4 13 1 10 9 2
7 10 12 13 15 9 0 2
12 15 1 15 4 3 4 13 1 10 12 9 2
6 3 15 13 10 9 2
33 11 7 11 2 15 15 13 1 3 12 9 2 4 13 1 9 1 10 12 1 9 7 15 4 13 3 1 10 9 1 10 9 2
22 1 10 9 2 11 11 4 13 1 10 9 1 10 9 3 0 7 4 13 10 9 2
20 10 9 1 11 4 13 1 10 10 9 2 1 9 2 9 1 9 7 9 2
37 10 9 2 9 1 10 9 1 10 9 3 13 1 10 9 2 4 13 1 9 1 10 12 2 1 9 1 9 2 16 4 4 13 1 10 9 2
11 9 1 10 9 1 10 9 1 10 11 2
11 10 9 13 1 12 1 12 9 1 9 2
10 9 1 9 3 10 9 1 10 9 2
6 9 1 10 11 0 2
36 11 2 1 10 9 1 10 9 1 10 9 1 10 9 15 4 13 10 9 0 1 10 9 1 10 11 1 11 2 3 10 9 1 10 9 2
20 1 10 9 13 3 13 15 9 1 10 9 1 9 1 10 9 1 10 11 2
40 1 10 9 2 0 2 1 15 1 10 9 1 9 1 10 11 1 10 11 4 4 13 10 9 1 0 9 1 10 9 1 11 11 11 7 1 10 9 11 2
21 1 15 1 10 9 13 1 10 2 12 2 4 4 3 13 10 9 1 10 9 2
15 10 9 4 4 13 7 10 10 9 13 2 0 9 2 2
16 1 10 9 10 9 0 1 10 9 11 11 4 13 10 9 2
30 15 13 1 10 9 1 9 1 10 9 1 10 9 1 10 11 2 15 13 1 10 12 1 10 12 9 1 9 0 2
8 10 9 4 13 10 0 9 2
25 10 0 9 4 13 1 13 1 9 10 9 1 9 7 10 9 1 10 9 1 10 15 4 13 2
10 10 9 1 10 9 4 4 3 13 2
30 10 0 9 4 4 13 1 10 11 1 10 11 2 3 10 9 4 13 1 10 9 1 10 9 1 9 1 10 11 2
6 10 9 4 4 13 2
28 1 9 4 13 3 1 10 9 16 3 13 13 15 1 9 7 16 1 15 15 4 13 1 10 2 9 2 2
6 9 0 1 12 9 2
17 11 2 10 9 4 13 3 12 9 1 10 11 2 1 11 11 2
10 13 0 7 10 9 4 13 15 0 2
30 16 4 4 13 1 10 9 1 10 9 2 4 13 1 10 9 2 1 9 7 9 1 9 2 13 15 1 10 9 2
17 10 0 9 1 9 4 13 9 3 1 10 9 7 1 10 9 2
25 12 9 4 13 2 15 13 10 9 1 10 9 2 7 10 15 4 13 10 9 13 1 10 9 2
11 1 10 9 3 9 7 12 9 1 9 2
6 13 1 9 1 11 2
12 13 1 9 7 13 1 9 1 13 10 9 2
7 9 1 9 1 10 11 2
14 12 9 7 12 9 0 13 1 10 9 1 10 9 2
44 11 2 12 9 2 12 9 0 7 12 10 9 2 4 4 13 7 3 13 1 10 9 1 9 1 10 9 1 10 9 0 1 11 2 10 9 1 10 9 2 0 1 9 2
45 10 12 13 1 10 11 1 9 1 2 11 11 2 2 10 9 3 0 1 10 9 1 9 1 11 2 1 10 9 1 10 9 7 1 10 9 0 1 11 2 1 10 9 11 2
66 10 9 13 10 9 11 11 2 12 9 2 1 11 11 2 11 2 2 10 10 9 11 2 12 9 2 7 11 2 12 2 10 9 11 11 2 12 9 2 1 11 2 11 2 2 10 9 11 11 2 12 2 1 11 2 10 9 11 11 2 12 9 2 1 11 2
14 13 7 1 9 1 9 10 9 0 1 11 2 11 2
2 13 2
12 2 4 13 1 9 0 3 1 10 9 2 2
46 10 9 4 13 9 9 2 7 10 9 4 13 1 11 3 3 2 1 10 9 15 13 1 10 9 1 11 2 15 1 10 3 0 7 0 9 0 1 10 9 2 13 1 10 12 2
22 1 13 10 9 1 10 9 4 13 10 9 1 9 1 9 0 7 1 10 9 0 2
29 10 11 4 13 1 9 15 1 10 9 3 0 1 10 10 11 2 13 1 9 2 9 1 10 11 2 9 0 2
12 3 13 16 10 9 1 10 9 4 13 9 2
22 13 1 11 3 15 13 10 9 9 1 2 11 11 2 2 4 13 10 9 3 0 2
25 1 10 12 1 10 0 9 4 4 13 10 9 11 11 2 15 15 13 1 10 9 1 10 9 2
10 11 2 11 11 1 9 12 11 1 9
5 12 9 1 9 2
8 2 10 11 3 13 3 2 2
14 11 2 0 9 0 1 10 11 13 1 10 9 0 2
26 1 10 9 1 10 11 0 15 4 13 10 9 0 12 9 1 9 1 9 2 1 9 7 1 9 2
14 3 9 4 13 1 10 9 2 1 9 7 1 9 2
15 1 10 11 13 12 12 10 9 1 9 2 9 11 2 2
13 10 9 0 4 3 13 16 10 9 13 3 0 2
3 1 9 2
6 13 13 1 10 9 2
53 11 1 11 2 11 2 2 10 0 9 2 11 11 1 12 9 2 1 9 1 10 9 2 11 2 1 11 1 11 1 10 11 2 4 13 9 1 10 9 0 16 13 10 9 1 10 9 15 13 1 10 9 2
27 3 13 1 10 9 7 1 10 9 0 1 10 9 2 10 9 4 13 9 1 10 9 1 11 1 11 2
19 10 9 2 0 1 11 3 16 1 9 0 2 4 13 10 9 1 9 2
15 1 10 9 1 10 9 10 11 1 11 4 13 10 9 2
3 10 9 2
21 11 2 10 9 2 3 13 9 9 9 1 10 9 2 4 4 13 1 10 12 2
20 1 3 10 3 12 9 15 13 1 10 9 0 7 1 10 9 1 10 11 2
15 1 15 3 1 10 0 9 4 13 1 9 7 9 0 2
28 1 10 12 11 11 13 10 9 1 10 9 13 15 1 9 9 9 2 1 9 1 10 9 7 1 10 9 2
15 10 9 13 10 9 7 11 11 11 4 13 10 0 9 2
2 9 2
7 9 1 9 1 10 11 2
39 11 2 11 2 2 10 9 2 15 15 4 13 1 9 0 2 4 3 13 1 11 2 11 2 2 10 9 1 9 1 11 11 2 0 1 10 10 9 2
10 10 9 1 10 11 3 13 1 9 2
11 4 13 10 9 0 1 0 11 1 11 2
15 10 9 13 13 13 1 10 9 1 10 9 1 10 11 2
15 1 13 10 9 2 10 9 1 10 9 4 13 1 11 2
19 1 10 9 4 13 3 10 9 1 10 9 1 11 2 15 4 13 9 2
9 1 10 9 3 4 13 13 9 2
2 9 2
7 10 9 11 13 1 11 2
36 11 2 10 9 15 13 11 11 2 10 0 9 1 10 11 11 2 13 10 0 12 9 1 10 9 1 9 1 9 2 15 13 3 1 11 2
52 10 9 0 2 13 1 9 1 10 9 1 11 2 4 13 10 9 2 9 2 2 10 11 11 11 2 1 9 0 1 11 2 15 4 13 9 0 1 9 1 10 9 0 11 11 1 3 12 9 1 9 2
23 9 1 10 9 4 4 13 1 11 11 1 2 13 2 10 9 1 10 9 1 9 0 2
11 13 0 13 15 2 7 15 0 15 13 2
12 10 10 9 0 13 9 3 13 2 3 13 2
32 10 9 1 10 0 9 2 13 1 0 9 2 13 1 10 0 9 2 4 13 10 0 9 2 10 0 9 2 10 0 9 2
10 10 0 9 4 13 15 10 0 9 2
9 1 15 13 0 7 13 1 13 2
21 1 15 2 10 9 13 0 2 16 15 13 9 16 10 9 4 13 0 1 15 2
21 1 15 13 0 16 13 16 15 2 15 15 13 1 10 10 0 9 2 15 13 2
42 15 13 1 9 10 10 0 9 15 2 13 10 9 1 10 0 9 0 2 1 11 11 1 11 2 1 11 2 1 11 2 13 16 4 13 0 1 13 15 3 15 2
10 1 10 9 16 10 9 13 3 3 2
11 1 9 2 10 9 13 10 9 1 9 2
27 15 3 13 3 3 0 2 3 0 2 3 0 1 10 15 2 7 13 3 10 9 1 9 0 7 0 2
14 1 11 2 16 13 16 10 9 4 13 1 9 0 2
30 3 2 1 10 9 2 10 9 3 13 3 2 16 10 9 4 13 1 15 2 15 13 16 4 3 4 13 15 15 2
5 3 3 13 0 2
22 3 1 10 9 2 3 2 10 9 1 10 0 9 13 0 16 13 13 3 1 15 2
5 3 3 13 0 2
12 16 15 13 10 9 13 3 2 13 1 9 2
14 7 16 10 9 1 10 9 13 9 15 15 3 13 2
18 13 13 10 9 2 13 1 10 9 2 13 10 0 2 13 10 9 2
8 13 13 0 2 13 2 13 2
11 13 10 9 0 2 10 9 1 10 9 2
3 15 3 2
34 3 1 10 9 0 2 10 9 1 10 9 0 13 3 0 1 13 1 15 2 1 13 10 10 0 9 2 7 13 1 4 15 13 2
12 3 15 4 13 7 13 10 9 1 10 9 2
10 1 1 15 2 15 3 13 3 3 2
20 13 0 1 10 9 0 1 10 9 2 1 15 10 9 13 16 10 9 13 2
6 15 13 3 10 3 2
28 7 1 10 0 9 2 1 10 0 9 2 9 2 9 2 10 9 2 10 9 4 13 10 9 1 15 3 2
11 13 11 11 2 10 10 9 13 1 9 2
12 13 11 10 11 2 13 10 9 1 10 11 2
14 7 3 13 10 9 1 13 3 1 10 0 9 0 2
34 3 1 10 10 9 0 15 13 10 9 1 15 13 10 9 1 10 10 9 2 10 9 1 10 10 9 2 10 9 1 10 10 9 2
7 7 15 3 4 13 15 2
22 3 15 13 9 1 10 9 0 2 1 10 9 1 9 2 1 9 15 13 1 15 2
11 10 9 4 13 1 10 9 10 9 0 2
7 11 11 11 1 10 12 2
8 2 11 0 1 10 9 2 2
2 11 2
12 15 13 13 10 9 1 13 12 9 1 11 2
16 2 13 10 9 7 9 1 9 1 10 9 1 10 9 2 2
14 11 2 9 1 11 1 9 0 7 9 1 9 0 2
35 11 11 2 10 2 9 2 1 10 0 9 2 4 13 1 10 9 1 4 13 10 9 0 1 13 10 9 1 12 9 0 13 1 11 2
29 9 1 10 9 13 15 1 13 10 9 1 10 11 1 10 9 0 0 2 10 11 2 13 1 10 9 1 11 2
15 15 13 1 10 9 3 0 13 1 10 9 1 11 0 2
19 1 12 9 10 9 1 11 15 4 13 1 13 9 1 10 9 13 11 2
5 1 10 9 13 2
8 2 15 13 10 9 13 2 2
11 3 1 10 0 11 4 4 13 0 9 2
20 7 3 1 10 0 9 3 1 10 0 9 11 11 2 11 4 13 10 9 2
35 2 1 10 9 4 13 10 9 7 9 1 9 0 1 10 9 1 10 9 0 1 10 9 1 12 9 2 9 0 1 13 10 11 2 2
16 10 9 0 15 4 13 1 11 2 11 7 11 1 10 12 2
29 11 2 0 9 0 1 10 11 2 13 0 9 1 10 3 0 9 0 7 4 13 10 9 0 1 10 9 0 2
28 1 10 9 4 13 3 9 0 1 10 9 7 1 10 11 11 11 2 13 2 0 1 10 9 1 11 2 2
36 1 10 10 9 15 13 16 1 10 12 10 9 1 11 13 0 1 13 1 11 12 9 1 10 9 1 10 9 0 0 11 7 1 10 11 2
26 10 9 3 13 1 9 2 3 1 9 1 10 9 1 11 1 11 7 1 10 9 11 1 10 11 2
53 10 9 1 10 9 0 4 13 0 1 10 12 2 16 1 13 10 9 11 11 15 4 4 13 1 10 9 1 12 9 0 1 10 11 11 2 11 11 7 11 11 2 13 10 12 9 12 1 10 9 1 11 2
32 1 10 9 10 9 4 13 1 10 9 0 0 2 3 3 4 13 10 9 1 10 9 1 11 11 2 10 3 0 9 0 2
30 10 11 4 4 3 9 13 1 13 9 1 10 9 1 11 11 2 7 1 10 9 11 13 10 15 1 13 10 9 2
13 7 1 10 9 9 2 9 7 9 13 1 9 2
11 3 1 10 9 15 15 13 1 10 9 2
40 2 10 11 2 4 13 11 1 15 1 10 0 9 1 10 9 0 1 11 11 2 13 1 10 0 9 1 10 9 0 0 1 10 9 12 1 10 9 0 2
18 13 10 9 0 1 9 15 13 1 10 9 1 13 1 10 9 0 2
17 10 11 2 13 1 10 9 11 2 9 2 13 0 1 10 9 2
31 1 10 9 10 9 4 3 13 1 13 10 9 1 9 1 10 9 1 10 11 16 1 10 0 4 13 10 9 0 2 2
19 10 12 9 0 4 13 1 11 3 3 2 1 10 9 1 10 9 12 2
21 3 4 3 13 10 9 4 13 0 1 10 9 7 15 13 1 9 1 10 9 2
14 3 1 13 10 9 1 10 9 11 4 13 12 9 2
13 15 4 13 3 1 10 9 1 10 12 9 0 2
17 1 10 9 1 10 9 11 11 4 13 3 10 9 1 10 9 2
10 1 10 10 9 10 9 0 3 13 2
26 7 3 10 9 0 4 13 10 9 1 10 0 9 1 10 9 1 10 9 15 4 13 10 10 9 2
30 1 10 9 1 9 3 10 9 1 11 15 4 13 12 9 1 10 9 1 10 11 2 13 1 12 12 9 1 9 2
14 7 10 9 1 10 9 11 13 10 12 9 3 0 2
17 2 3 12 12 9 4 13 1 13 1 10 9 0 10 9 0 2
3 7 3 2
22 10 9 0 13 1 13 10 9 1 9 0 13 10 9 1 11 2 0 1 0 11 2
17 10 9 1 10 9 13 1 13 0 10 9 0 3 1 11 2 2
21 10 0 9 13 0 0 2 3 10 9 1 10 9 1 11 13 1 10 0 9 2
26 2 1 10 9 13 12 9 1 11 2 9 1 11 11 2 7 12 1 10 9 1 10 11 2 11 2
24 9 1 10 10 9 13 10 9 1 9 1 10 11 1 9 1 10 9 1 10 11 11 11 2
9 11 13 10 9 1 9 1 9 2
21 10 9 4 13 1 10 11 1 12 9 1 10 9 15 11 11 13 1 11 2 2
9 1 9 1 10 9 11 1 11 2
13 2 13 9 16 10 9 1 10 9 4 13 2 2
3 10 11 2
11 2 10 9 13 9 1 10 9 0 2 2
2 11 2
9 16 10 9 13 10 11 13 0 2
3 10 11 2
7 9 0 1 10 0 9 2
12 11 2 15 13 9 7 9 2 9 7 9 2
29 15 4 13 11 1 9 2 1 10 9 1 10 2 11 2 2 13 1 10 0 9 11 1 11 1 10 9 0 2
61 10 11 13 10 2 0 9 2 1 10 0 9 1 10 9 1 9 0 2 13 2 0 9 2 1 15 2 13 10 9 11 1 0 9 2 7 3 13 2 10 9 3 3 0 1 10 9 3 3 1 0 2 7 3 1 9 2 1 9 0 2
21 2 13 9 16 10 9 1 9 4 3 13 2 2 13 2 7 13 10 9 0 2
14 2 10 9 13 3 1 3 9 1 10 9 0 2 2
6 13 0 2 9 2 2
22 7 10 11 13 1 10 9 1 10 0 9 0 3 13 1 10 9 2 9 9 2 2
10 10 9 11 11 3 13 10 0 9 2
46 2 13 3 16 11 13 1 2 13 15 1 9 2 1 9 1 10 9 1 11 2 13 2 7 16 4 15 13 10 9 1 10 9 15 13 1 10 0 1 10 9 1 10 9 2 2
12 3 2 7 3 2 1 11 2 13 10 9 2
34 2 16 1 13 10 9 1 10 9 0 13 13 1 10 11 2 3 1 10 0 0 9 2 16 15 13 1 10 13 3 10 9 0 2
20 16 2 13 15 2 1 9 1 10 11 2 11 13 10 9 1 10 9 2 2
14 7 10 9 16 11 4 2 13 1 9 2 1 11 2
11 2 3 10 9 3 15 13 2 13 2 2
15 11 1 10 9 1 11 4 13 3 10 9 1 9 2 2
29 3 2 11 13 0 1 10 13 10 9 1 10 0 9 2 3 13 16 2 10 9 0 4 4 13 1 9 2 2
15 2 13 10 3 1 13 1 10 9 10 9 1 13 9 2
19 13 3 2 7 15 13 15 16 3 1 10 9 15 15 13 10 9 2 2
15 1 10 10 9 13 3 10 9 1 10 9 11 11 11 2
23 2 10 11 4 13 10 0 9 1 9 2 3 3 1 10 2 9 9 2 2 13 2 2
23 1 10 9 13 10 11 1 10 9 1 10 9 2 7 15 13 3 3 1 10 9 0 2
22 3 3 13 1 9 3 0 2 3 16 15 4 13 15 1 10 9 9 1 10 9 2
35 10 15 13 10 0 9 3 1 10 9 1 10 9 1 10 9 2 13 16 13 10 9 1 10 9 2 7 0 1 10 9 1 10 9 2
22 6 2 11 3 15 4 3 13 13 3 2 7 15 15 13 13 10 9 1 11 2 2
12 10 9 13 3 1 10 9 1 10 9 11 2
6 13 2 13 0 9 2
12 1 10 9 9 7 9 1 9 1 10 9 2
8 10 9 4 13 10 9 3 2
3 10 9 2
10 9 1 10 9 1 10 9 1 11 2
38 11 2 1 10 9 1 10 9 1 10 9 1 10 9 15 4 4 13 1 9 1 10 9 1 11 2 1 10 11 13 10 2 9 2 1 10 9 2
18 1 10 9 1 10 9 1 10 11 13 4 15 13 10 9 1 9 2
38 15 4 3 13 16 13 15 1 10 9 13 1 10 9 1 10 9 10 9 1 10 9 1 0 9 0 15 13 1 9 10 0 11 7 10 9 11 2
33 3 0 1 10 9 2 10 9 4 13 3 10 9 1 10 9 2 13 1 10 9 0 1 13 13 1 9 10 9 1 10 11 2
12 10 9 4 13 1 10 9 1 10 0 9 2
24 3 1 10 9 1 10 9 1 10 9 4 13 9 1 10 15 15 13 3 11 7 10 9 2
17 10 9 4 3 13 1 9 10 9 1 13 10 9 1 10 9 2
7 10 9 3 4 4 13 2
30 10 9 1 13 1 3 13 3 16 13 15 1 0 15 4 13 1 9 16 4 4 13 10 9 1 10 15 4 13 2
7 13 10 9 1 10 9 2
44 4 13 0 13 10 9 1 9 1 10 2 9 2 7 4 3 13 0 16 10 9 0 1 10 9 1 10 9 13 3 15 15 4 1 0 13 1 10 0 11 7 10 9 2
20 13 16 15 1 10 9 4 4 13 1 10 9 16 13 1 9 1 10 11 2
9 15 15 13 3 1 13 10 9 2
15 1 9 10 0 9 4 4 13 1 10 9 1 10 11 2
23 1 9 1 9 15 4 13 16 10 9 13 1 9 1 10 9 0 7 4 4 13 11 2
40 10 15 13 1 10 9 2 15 3 1 9 1 10 9 1 10 9 1 10 11 2 15 13 9 0 1 10 9 1 12 1 10 9 1 12 9 1 9 0 2
32 1 13 3 10 9 2 11 4 13 10 9 1 13 1 10 9 1 10 11 7 10 0 9 4 13 1 9 1 10 0 9 2
17 10 9 13 3 10 9 7 3 1 10 9 15 13 1 10 15 2
34 1 10 9 0 10 0 9 4 13 7 3 10 9 2 13 7 3 13 1 10 9 2 4 13 1 13 10 9 1 10 2 9 2 2
18 1 10 9 2 1 10 9 2 13 3 0 10 9 0 1 10 9 2
6 11 2 13 7 13 2
6 2 13 10 9 2 2
7 0 10 9 13 9 11 2
17 11 2 10 9 1 10 0 15 13 1 10 0 9 1 9 0 2
31 1 10 9 10 9 11 11 2 12 9 2 0 9 0 1 10 11 2 13 10 9 3 3 0 2 7 13 10 9 0 2
14 10 9 15 4 13 10 9 1 9 1 10 9 0 2
36 1 10 10 9 3 4 4 13 10 9 2 3 16 3 15 1 13 1 9 1 10 9 1 10 9 1 9 11 7 1 10 9 0 1 9 2
20 3 1 10 9 0 2 4 13 2 3 1 9 0 2 1 10 9 1 3 2
2 9 2
16 2 1 9 13 1 9 2 1 15 13 10 9 1 10 9 2
16 10 9 13 10 10 9 2 13 10 9 11 2 12 9 2 2
11 13 9 1 13 2 3 4 13 1 15 2
8 15 4 13 1 9 1 9 2
6 10 9 15 4 13 2
5 3 0 2 2 2
12 15 13 10 9 2 0 2 11 11 2 0 2
17 2 15 13 1 10 9 0 1 11 0 1 9 1 10 11 2 2
30 13 1 11 2 3 1 10 9 1 11 11 7 3 1 10 9 1 11 2 10 9 4 13 10 9 0 10 12 9 2
26 3 1 13 13 1 10 9 11 16 1 10 11 13 10 0 11 2 3 3 13 1 15 2 0 2 2
6 10 9 13 1 11 2
34 13 0 16 10 9 1 11 2 1 10 15 3 1 10 9 13 10 9 1 9 10 12 9 2 4 13 10 9 1 10 9 1 11 2
31 13 0 16 10 9 1 11 7 1 11 2 15 3 0 2 15 13 1 10 9 16 11 13 3 7 13 3 1 13 15 2
41 3 10 9 3 3 0 13 10 0 9 0 1 10 12 1 10 0 9 0 1 3 2 13 10 9 0 1 10 11 11 1 10 0 9 1 10 9 1 3 11 2
23 3 3 16 12 9 1 9 0 0 4 13 10 9 15 15 13 10 9 1 11 7 11 2
21 3 3 16 3 1 3 10 9 13 0 2 15 13 3 1 9 2 9 7 9 2
35 7 3 3 16 1 10 0 9 1 11 4 13 9 1 9 2 16 12 9 3 10 9 1 10 12 9 0 13 9 1 10 9 1 11 2
79 10 9 1 11 11 13 3 2 13 1 10 9 1 10 10 0 9 15 1 0 9 4 13 0 10 9 1 11 2 13 1 10 9 1 10 9 1 9 0 15 10 9 13 2 9 1 10 9 2 7 15 4 13 10 10 9 0 3 3 1 10 10 9 2 13 15 2 3 2 1 13 1 10 9 1 10 3 9 2
3 1 3 2
34 1 10 0 9 6 2 16 13 7 13 1 10 9 0 10 9 1 10 9 0 2 16 10 9 1 10 9 0 13 13 10 10 9 2
72 7 4 13 10 9 1 13 3 1 3 10 9 1 11 2 7 4 13 3 10 9 1 12 9 15 3 1 15 15 4 13 2 15 4 13 10 9 1 10 9 1 9 0 16 13 10 15 0 7 10 15 0 2 15 13 10 9 1 10 9 1 10 9 13 9 7 9 1 10 9 13 2
9 10 9 3 4 13 10 9 0 2
7 3 13 15 10 10 9 2
55 7 16 10 9 0 15 4 13 13 10 2 9 2 13 1 9 1 11 2 4 13 10 9 1 10 9 0 2 13 1 9 0 3 7 3 1 3 7 0 3 1 10 9 0 15 10 12 11 0 4 13 1 12 9 2
13 15 4 13 3 1 3 10 9 1 11 4 13 2
18 16 4 13 1 10 11 1 10 9 1 10 9 0 2 0 2 0 2
40 7 3 10 9 4 13 1 10 10 9 13 1 10 9 0 2 3 1 10 9 4 13 1 10 10 9 10 9 0 2 3 4 13 10 10 9 13 10 9 2
15 15 13 2 3 2 9 1 0 2 9 1 10 9 2 2
32 10 11 2 10 11 2 10 9 0 2 3 13 3 2 3 1 10 9 1 10 12 0 9 2 1 10 9 1 10 9 0 2
30 7 1 0 9 10 9 4 13 1 11 2 1 10 9 1 10 9 1 10 12 11 2 3 3 11 4 4 13 15 2
5 3 15 4 13 2
56 10 9 15 10 9 0 4 13 1 10 9 15 13 3 0 2 13 1 10 10 9 16 10 9 1 11 11 15 13 1 3 10 0 9 2 16 10 9 0 2 13 10 9 1 10 9 2 13 10 9 1 10 9 1 11 2
18 15 13 10 9 15 15 13 1 10 9 1 10 1 3 1 10 9 2
13 10 9 13 2 7 10 9 11 4 13 1 9 2
36 10 9 3 3 13 13 15 2 16 13 3 11 11 2 16 13 10 9 1 13 10 9 2 7 3 10 9 2 16 13 2 1 10 9 11 2
23 7 3 16 15 4 13 9 1 10 9 0 2 1 10 10 9 15 15 13 7 15 13 2
62 10 9 15 10 9 13 1 9 2 15 9 7 9 3 1 15 2 13 10 9 1 10 2 9 9 2 1 9 0 1 13 10 9 1 10 0 11 2 10 9 1 10 0 9 0 2 10 9 1 10 9 15 10 9 1 11 3 13 3 1 13 2
30 1 10 9 4 13 1 10 11 7 9 15 9 1 11 11 15 3 4 13 13 1 10 0 0 9 1 10 3 9 2
2 11 2
8 1 10 12 13 12 10 9 2
66 10 12 9 12 2 12 1 10 12 2 11 12 2 1 10 12 11 13 1 10 11 11 1 10 11 1 10 2 9 0 2 1 9 1 10 9 0 7 1 10 9 1 10 11 2 13 1 10 9 1 11 1 10 9 1 9 1 9 1 10 9 0 1 10 11 2
33 10 9 0 13 1 9 16 12 9 1 9 1 10 2 11 11 11 2 2 0 2 13 9 1 10 9 7 15 13 1 9 0 2
10 15 13 7 13 1 10 9 1 11 2
10 3 3 15 13 3 1 10 9 0 2
21 10 9 4 13 1 10 9 2 15 13 1 9 7 13 1 10 9 1 10 9 2
2 11 2
7 13 7 13 12 9 11 2
8 10 9 4 13 10 0 9 2
22 1 10 9 1 10 9 1 10 9 2 10 0 9 0 4 13 1 13 1 10 9 2
38 13 16 10 12 2 13 3 7 13 1 0 9 2 2 10 9 1 10 11 11 2 1 13 0 9 2 4 13 16 10 9 4 13 1 9 1 9 2
25 10 0 9 1 10 11 11 4 13 16 10 9 4 13 1 12 9 7 16 15 1 15 4 13 2
28 3 10 9 1 9 1 15 1 10 9 4 4 13 1 10 9 1 10 9 1 10 15 4 4 13 10 9 2
25 12 9 0 7 12 1 10 10 9 4 4 13 7 13 1 10 9 1 10 9 1 10 9 0 2
10 11 2 9 1 10 9 1 10 9 2
8 10 9 9 1 10 9 0 2
7 4 4 13 3 1 12 2
9 2 4 13 9 3 1 10 9 2
9 13 9 0 7 10 9 0 2 2
14 11 2 15 4 13 2 0 1 10 9 1 12 9 2
42 10 9 1 11 11 2 1 10 10 9 11 2 12 9 2 7 11 2 12 2 1 11 11 2 1 11 11 2 1 11 11 4 4 13 1 10 9 1 10 10 9 2
43 10 9 4 13 9 9 2 7 10 9 4 13 1 11 3 3 2 1 15 1 10 9 0 3 0 1 10 9 2 15 1 11 2 1 11 2 0 1 10 9 1 9 2
31 10 12 9 13 0 1 10 11 11 11 7 1 11 2 1 10 9 1 10 11 2 4 13 10 9 0 1 10 9 9 2
17 1 10 9 4 13 10 9 0 12 9 1 9 1 10 10 9 2
66 3 1 10 12 9 4 13 9 1 10 9 3 10 9 0 1 11 2 11 11 2 13 11 2 2 13 0 3 3 7 3 13 1 10 9 1 11 2 10 0 9 2 11 11 2 3 0 2 7 3 1 0 9 1 9 2 7 10 9 0 1 10 9 7 9 2
10 1 10 9 1 10 9 15 13 3 2
29 10 9 4 3 13 10 9 1 9 1 10 9 2 10 9 3 13 2 16 4 4 13 1 10 9 1 9 0 2
57 10 0 9 1 10 9 2 11 11 2 4 13 16 1 13 15 4 13 9 2 15 13 9 0 7 13 10 9 13 7 15 2 4 13 1 9 0 3 1 10 9 15 4 13 1 13 1 10 9 7 3 1 10 0 9 2 2
41 2 4 4 13 7 3 13 2 2 4 13 1 10 9 1 10 9 1 11 11 1 11 10 9 2 11 11 2 15 3 4 13 1 3 13 1 9 1 0 9 2
11 10 9 3 4 4 13 7 13 1 11 2
27 10 9 4 13 1 11 2 10 9 1 10 9 15 4 13 3 7 15 13 3 3 9 1 10 9 0 2
8 13 0 16 3 15 13 9 2
17 15 4 13 1 10 9 1 13 1 15 3 10 12 9 3 0 2
30 10 9 1 11 2 1 9 1 10 9 1 10 11 2 1 10 11 7 1 10 11 2 13 10 3 0 1 10 11 2
28 13 1 10 12 4 3 3 13 1 10 9 13 1 10 9 0 2 3 1 9 0 2 7 1 10 9 0 2
26 3 15 13 3 10 0 7 0 9 1 9 16 13 10 9 11 11 2 13 1 9 0 1 10 12 2
24 10 9 1 10 9 13 3 15 13 3 1 10 9 1 11 7 1 10 9 1 10 11 0 2
25 15 2 13 10 9 2 13 10 10 9 2 7 15 13 7 13 15 1 13 10 9 1 9 0 2
58 1 10 9 2 16 13 0 2 16 4 13 1 10 11 10 9 1 10 9 1 11 2 11 11 2 16 10 9 13 1 10 9 1 9 13 9 4 13 0 2 13 3 0 16 10 11 13 15 1 10 9 3 0 1 10 10 11 2
44 1 9 10 9 0 2 1 9 0 2 1 9 7 1 9 2 15 15 13 1 9 7 1 9 2 3 9 7 9 4 13 1 10 9 1 9 1 10 9 7 13 10 9 2
22 3 13 0 13 15 1 10 9 1 9 0 15 15 4 13 3 13 10 2 9 2 2
13 13 1 10 9 1 11 13 10 0 7 0 9 2
38 13 13 15 3 1 10 13 10 10 9 1 10 9 1 9 15 3 13 10 9 1 13 15 13 7 13 15 13 3 1 10 9 1 12 9 1 9 2
21 10 9 13 3 10 9 7 1 9 0 13 13 10 9 1 10 9 1 10 9 2
27 9 1 11 1 10 9 1 11 11 2 10 9 1 10 15 10 9 13 10 9 1 10 9 1 10 11 2
8 2 9 4 13 10 11 2 2
18 10 9 11 4 13 1 3 1 11 2 11 3 4 13 1 12 9 2
13 11 2 10 9 1 9 4 13 0 10 9 3 2
13 2 13 15 0 1 13 1 10 9 1 9 2 2
22 1 10 0 9 11 11 2 11 2 2 13 1 10 9 0 2 4 13 10 9 0 2
24 11 11 4 13 1 13 1 3 1 10 11 2 7 9 0 2 1 10 0 9 2 4 13 2
17 2 11 13 15 2 15 2 11 2 10 9 2 13 11 2 2 2
36 3 2 1 10 9 0 1 11 11 2 9 1 12 9 1 10 9 0 2 1 11 11 3 4 13 10 0 9 2 2 10 9 4 13 2 2
43 2 15 4 13 1 10 12 2 15 1 10 11 11 11 2 15 4 13 16 9 11 4 4 13 1 10 9 2 2 2 13 10 9 15 1 10 9 2 11 2 12 9 2
13 11 11 2 12 9 2 13 10 9 0 1 11 2
24 12 9 3 4 13 1 13 1 10 11 2 15 4 13 1 10 9 0 1 13 1 12 9 2
7 9 2 2 9 2 9 2
17 3 4 13 3 10 9 2 1 10 9 11 11 2 1 15 11 2
13 1 10 12 15 4 13 1 11 7 15 4 13 2
33 2 1 15 10 9 1 10 11 13 15 2 13 11 2 2 7 16 4 13 11 7 11 4 13 16 3 4 4 13 3 1 3 2
19 10 9 4 13 10 9 0 2 1 10 9 9 11 4 13 13 1 11 2
11 10 9 4 13 2 3 13 10 9 2 2
2 9 2
20 2 7 6 2 10 9 0 4 13 1 11 1 0 9 7 3 4 13 15 2
12 15 13 1 13 16 13 3 10 9 2 2 2
18 13 0 3 15 2 13 1 9 2 1 10 0 9 1 10 10 9 2
6 2 4 4 13 15 2
24 1 9 15 4 13 2 2 2 13 11 2 1 10 9 10 9 9 1 10 9 13 1 11 2
20 3 9 11 2 10 9 2 15 1 11 11 13 10 9 1 9 7 10 9 2
31 2 6 2 13 10 9 1 9 2 13 11 11 2 9 1 10 9 2 2 1 10 9 1 10 15 2 3 1 3 2 2
10 9 3 3 0 2 1 10 0 9 2
9 11 11 2 12 9 2 9 0 2
26 1 10 11 4 13 1 10 0 9 9 0 2 3 1 10 9 9 11 11 2 12 9 2 1 11 2
33 13 15 1 10 9 2 11 11 2 1 11 2 13 1 9 2 4 4 13 10 9 13 1 11 11 2 9 1 10 9 1 9 2
8 2 13 0 2 13 1 11 2
21 3 11 11 2 12 9 2 0 1 11 2 9 1 9 2 3 13 3 10 9 2
45 2 10 9 15 4 13 1 10 9 1 10 11 2 13 11 11 2 9 1 11 11 2 15 1 12 9 15 13 1 9 1 10 11 2 2 7 3 15 4 13 9 1 0 9 2
10 15 3 13 16 10 9 3 15 13 2
25 3 1 10 0 12 9 2 1 9 1 9 4 13 12 1 9 7 9 2 7 12 13 0 2 2
6 2 10 9 13 3 2
10 13 10 10 9 2 2 13 10 9 2
12 15 2 1 10 9 2 13 3 1 10 9 2
29 2 10 9 11 11 15 4 13 1 9 2 13 11 2 2 7 1 10 11 10 9 1 10 9 4 13 0 2 2
8 10 3 0 9 0 1 11 2
10 11 2 9 1 10 9 1 10 9 2
48 11 2 10 9 1 10 11 2 9 1 10 9 2 4 13 1 10 10 9 9 1 10 9 1 11 11 2 10 9 0 15 4 13 10 9 1 10 9 1 13 10 9 1 9 1 10 9 2
24 10 9 4 4 13 3 1 10 9 2 1 10 9 2 11 1 10 9 2 13 1 11 11 2
34 1 10 9 1 10 9 1 10 11 2 15 3 1 4 15 13 13 12 9 1 10 9 0 2 15 13 10 0 9 1 10 9 0 2
39 11 11 13 1 10 9 1 13 10 9 1 10 9 13 1 13 1 10 9 2 3 3 1 12 9 2 15 15 13 7 13 10 0 9 1 15 7 15 2
5 13 1 10 9 2
16 10 9 1 10 11 4 13 3 0 1 10 9 1 10 9 2
12 7 10 9 4 13 1 10 9 1 10 9 2
20 10 9 1 11 2 11 7 11 13 10 9 15 13 1 10 9 1 9 0 2
25 3 3 1 3 10 9 1 9 0 3 4 13 2 1 10 12 2 9 1 9 0 1 10 9 2
26 1 3 10 9 4 13 1 9 1 9 2 9 7 3 1 9 15 13 10 9 1 13 9 1 9 2
25 10 9 1 11 11 2 15 1 10 10 9 4 13 10 0 9 2 4 3 13 1 10 9 0 2
8 9 1 15 2 9 1 15 2
33 13 1 13 1 13 10 9 1 9 1 9 2 13 9 7 0 9 2 7 1 10 9 4 13 1 9 10 9 1 10 11 12 2
27 4 3 13 1 13 1 10 9 1 9 0 2 13 1 10 10 10 9 10 9 1 9 0 7 10 9 2
57 1 0 2 1 9 2 15 13 1 10 9 13 3 10 9 1 9 1 10 9 15 3 13 1 10 9 2 3 13 1 9 1 10 9 0 2 13 10 9 1 10 9 1 9 1 10 9 2 9 1 13 2 9 1 13 2 2
25 3 2 1 10 9 1 9 1 10 10 9 2 10 10 9 15 4 3 13 1 9 1 10 9 2
18 10 9 1 10 11 4 13 9 0 2 3 4 13 13 15 1 9 2
30 10 9 1 10 9 2 15 1 10 10 9 1 11 4 13 10 9 1 9 2 15 4 13 10 9 1 10 0 9 2
23 9 15 13 9 1 10 9 1 9 2 0 9 4 13 1 3 10 9 1 9 7 9 2
11 0 3 10 9 1 10 9 1 9 0 2
42 10 9 11 2 10 3 0 9 0 1 11 2 13 1 10 12 7 13 1 3 12 9 2 4 3 13 1 0 9 1 9 7 9 0 3 1 10 0 9 1 9 2
12 2 1 10 9 15 13 7 3 15 13 2 2
18 3 3 15 3 2 1 9 10 9 1 10 9 15 3 13 1 13 2
5 10 9 13 0 2
18 15 13 3 12 12 9 15 13 1 9 0 7 13 9 1 10 11 2
27 15 13 12 9 1 10 9 2 3 1 13 2 16 10 10 9 1 10 11 13 3 3 1 13 2 2 2
34 13 10 9 1 10 0 9 1 11 11 2 15 1 10 9 13 3 1 11 2 13 1 10 9 11 7 1 10 9 11 12 9 3 2
25 11 13 15 1 10 9 1 2 9 2 0 15 13 1 11 2 3 1 10 9 1 10 9 0 2
40 13 1 3 12 1 10 12 9 3 0 13 1 10 11 2 7 3 1 10 9 1 0 9 2 10 10 9 15 13 1 11 2 11 2 11 2 11 7 11 2
26 7 13 3 1 10 9 2 13 2 0 2 1 10 9 1 9 0 2 16 15 4 3 13 0 9 2
44 2 1 10 11 2 3 2 3 1 3 2 3 15 4 3 13 9 1 10 0 9 1 10 9 1 9 2 13 11 11 2 9 1 10 11 0 1 10 9 1 10 9 2 2
11 3 2 10 9 13 1 0 9 7 9 2
30 15 13 1 10 9 0 7 10 9 15 15 13 1 13 1 10 9 1 11 2 7 1 15 3 4 3 13 9 0 2
25 3 1 10 9 3 4 4 13 2 3 1 9 2 9 7 9 1 10 11 13 3 3 13 15 2
21 3 13 16 10 9 13 9 1 9 7 9 2 7 9 3 15 15 13 3 2 2
74 11 2 15 4 13 1 11 10 0 9 7 4 13 11 2 13 16 1 10 9 2 3 1 10 9 7 10 9 1 9 1 10 11 2 10 9 15 4 13 2 7 16 10 9 0 4 13 10 9 7 13 10 9 2 2 13 10 9 0 15 4 13 10 9 2 2 2 15 0 13 1 10 9 2
35 3 1 11 11 2 15 4 13 9 7 9 0 2 10 11 0 13 10 9 0 1 10 10 11 1 11 2 15 13 0 1 10 11 11 2
23 10 11 2 11 0 2 2 9 0 1 11 2 15 13 1 10 9 0 1 10 9 0 2
13 11 11 2 9 0 1 11 2 13 10 9 0 2
22 3 15 13 10 11 1 11 2 11 2 2 10 11 1 11 7 10 9 0 7 0 2
20 13 3 15 0 15 2 1 10 11 0 2 4 13 10 9 1 9 3 0 2
22 1 9 11 11 2 0 2 13 1 10 9 12 1 10 9 0 1 15 13 10 9 2
27 7 9 11 11 2 0 2 13 1 0 12 9 1 10 9 1 10 11 2 9 11 2 1 10 9 12 2
41 7 11 11 2 0 2 12 9 2 13 3 1 10 12 1 10 9 1 9 7 15 1 10 9 16 13 1 13 10 9 1 10 2 10 2 9 0 2 1 11 2
5 11 1 10 11 2
19 11 2 3 1 10 0 11 11 11 15 13 1 15 1 10 10 9 0 2
43 7 13 1 10 9 1 10 11 1 11 11 11 11 1 9 2 1 9 2 1 10 9 0 15 13 10 9 1 10 9 0 7 15 0 2 13 1 9 15 2 11 11 2
23 7 10 0 9 1 9 15 10 9 1 10 11 4 13 1 10 9 1 10 11 1 11 2
47 2 4 13 10 9 0 2 7 13 15 1 11 7 13 9 1 9 1 10 9 1 10 9 0 2 4 13 10 9 0 2 4 13 13 9 1 10 9 11 2 15 13 10 9 0 2 2
33 16 2 13 10 9 1 10 11 11 2 2 13 13 10 9 1 10 9 0 7 10 9 0 2 15 13 1 2 13 10 9 2 2
21 10 9 2 15 2 15 1 11 4 13 1 9 0 2 1 10 9 2 11 11 2
31 2 1 10 9 2 4 13 2 15 13 10 9 1 9 7 1 11 10 10 9 4 13 1 10 9 0 1 10 9 2 2
20 10 9 1 11 7 10 9 1 10 11 13 9 0 1 10 9 9 1 9 2
28 2 1 10 9 0 2 4 13 2 13 1 9 1 9 9 0 7 1 10 9 1 11 2 1 3 10 11 2
12 7 1 10 9 1 10 11 15 13 11 2 2
12 7 15 2 13 2 13 0 1 13 10 9 2
24 2 15 4 13 1 11 16 3 10 9 3 0 4 4 13 13 10 9 1 10 9 0 2 2
19 11 4 13 16 10 11 3 4 13 10 9 1 11 1 10 10 9 11 2
5 10 9 11 0 2
26 10 9 3 13 0 2 10 9 1 10 9 13 2 0 2 2 7 10 9 3 4 13 15 1 13 2
2 11 2
8 2 11 1 10 9 0 2 2
16 2 3 3 1 13 13 13 10 11 7 13 10 9 12 2 2
12 2 10 9 15 4 13 2 7 15 13 0 2
9 3 10 9 1 10 9 4 13 2
9 3 3 13 10 9 13 9 2 2
12 2 16 10 9 3 15 13 1 13 2 2 2
27 10 11 4 13 10 9 1 10 9 2 10 9 13 2 10 9 13 2 15 13 1 13 2 1 10 9 2
31 7 3 15 2 11 11 2 15 1 10 0 9 3 4 3 13 1 10 10 9 0 7 1 9 9 0 2 3 13 0 2
8 10 9 3 13 3 3 0 2
14 16 10 9 2 3 2 2 3 15 13 1 13 2 2
19 15 1 10 9 11 13 1 3 10 9 0 1 10 0 9 1 10 9 2
12 13 1 9 1 9 7 1 10 2 9 2 2
20 1 11 11 2 3 11 15 13 3 1 10 13 16 2 10 9 4 13 2 2
2 3 2
12 10 9 2 1 10 10 9 2 3 4 13 2
9 2 10 11 4 13 9 3 0 2
19 3 2 13 15 15 4 13 2 10 10 11 4 13 1 10 9 0 2 2
8 15 13 10 9 1 13 3 2
37 2 3 15 4 2 13 11 2 13 1 13 1 3 4 13 10 11 2 7 1 4 13 3 10 9 2 1 10 9 1 10 9 12 1 10 11 2
12 15 13 10 9 2 13 15 13 10 9 2 2
5 13 9 2 3 2
5 3 2 3 13 2
18 7 3 10 11 12 3 4 3 13 7 3 15 4 13 10 0 9 2
23 11 11 15 4 13 3 9 1 10 9 0 1 10 9 0 1 13 15 1 9 10 9 2
6 15 13 3 10 9 2
12 10 9 13 13 10 9 1 10 9 1 9 2
51 3 10 0 9 15 4 13 1 13 10 10 2 9 1 10 9 2 1 10 9 7 10 9 1 10 9 0 15 13 1 10 9 1 10 9 1 10 9 7 1 15 3 0 1 10 9 9 3 9 3 2
16 1 10 15 4 13 2 0 2 3 10 9 1 10 9 11 2
41 10 9 13 10 9 1 10 11 1 10 0 9 1 10 9 0 7 13 16 10 0 11 13 2 10 0 9 1 9 7 1 9 1 10 11 7 1 10 11 2 2
12 13 3 10 0 9 1 10 9 1 10 9 2
18 1 10 9 10 9 1 10 9 1 10 9 1 9 13 1 10 9 2
8 11 13 10 9 1 10 11 2
18 13 3 16 13 10 9 0 1 10 9 1 10 9 2 13 11 11 2
24 11 11 13 16 11 13 10 9 1 10 10 9 1 2 10 0 9 1 9 1 10 9 2 2
32 1 10 9 1 9 2 3 2 13 13 10 9 1 13 3 10 2 9 2 2 13 1 13 10 9 1 10 11 2 1 9 2
19 16 9 15 13 2 15 15 4 13 1 10 9 1 10 9 2 1 11 2
8 7 13 3 16 13 10 9 2
19 16 1 10 11 10 9 1 10 9 4 13 10 9 1 15 1 10 9 2
15 3 3 16 10 9 11 13 4 15 13 1 10 9 0 2
21 11 2 3 2 3 13 10 0 1 13 1 10 9 10 9 1 9 1 10 9 2
31 11 11 4 13 3 9 3 3 1 10 10 9 3 0 1 10 9 1 10 9 2 1 10 15 11 13 3 10 10 9 2
11 11 11 13 1 10 0 9 10 9 0 2
11 15 13 3 1 9 0 7 1 9 0 2
18 1 11 2 16 10 9 4 13 1 12 1 10 9 13 3 0 2 2
14 16 10 9 1 10 9 13 10 9 1 9 1 15 2
22 10 9 1 10 9 0 4 13 13 10 9 7 4 13 10 9 1 10 9 1 9 2
7 3 4 13 10 9 0 2
12 2 3 10 9 1 10 9 4 3 13 2 2
11 16 2 10 9 3 15 13 1 13 2 2
3 10 9 2
11 1 10 9 0 1 10 9 1 10 11 2
5 3 1 10 9 2
10 1 15 7 11 9 0 7 0 9 2
15 11 11 4 13 12 0 9 2 1 13 10 10 0 9 2
52 10 9 0 15 15 4 13 11 11 2 9 0 1 11 2 10 15 2 3 2 3 15 4 3 13 1 10 0 9 2 0 9 1 11 2 0 0 7 0 0 15 13 2 13 1 9 1 9 2 10 11 2
9 10 9 2 3 2 3 13 9 2
33 11 13 10 9 3 2 1 10 9 1 10 9 2 1 11 2 9 1 9 3 1 11 2 3 13 10 9 1 10 9 1 11 2
21 15 15 4 13 15 13 0 2 0 2 1 9 0 2 0 9 1 10 0 11 2
12 15 13 3 3 2 1 11 1 10 9 12 2
32 13 2 1 10 0 9 2 1 4 13 1 10 9 0 9 15 11 4 13 1 2 13 10 9 1 9 1 10 12 9 2 2
37 1 9 11 15 13 7 15 13 2 1 10 9 16 2 1 4 13 10 9 1 10 9 2 13 1 10 13 10 9 1 10 11 1 10 9 12 2
13 10 11 11 2 9 0 2 4 3 13 10 9 2
53 15 13 3 11 11 1 11 2 9 1 11 7 11 2 16 1 10 12 13 1 10 0 9 10 9 1 9 7 9 1 10 9 13 1 13 15 1 10 9 1 10 9 1 13 10 9 1 10 11 7 10 9 2
15 1 10 12 11 11 13 10 0 10 9 0 13 11 11 2
41 1 3 10 9 1 11 7 10 11 4 13 3 1 15 2 10 11 7 11 2 9 1 9 0 7 0 13 1 10 9 0 2 9 1 10 2 9 2 3 0 2
12 15 13 1 10 15 7 1 10 0 11 11 2
5 7 15 13 3 2
6 10 9 13 3 11 2
19 13 15 15 15 10 9 15 4 13 7 13 1 9 10 9 3 3 0 2
22 10 9 1 11 11 15 15 13 1 10 11 11 1 10 10 0 9 7 3 9 11 2
14 9 7 9 0 3 4 3 13 1 10 9 1 11 2
44 1 10 12 3 0 3 13 10 9 0 7 10 9 0 13 1 10 0 11 11 2 13 1 9 7 13 10 9 0 1 11 11 2 9 0 9 0 2 2 3 13 1 11 2
14 15 13 3 3 10 9 0 15 13 1 0 12 9 2
9 10 9 0 15 13 9 7 9 2
23 10 11 0 15 13 10 0 9 0 1 10 15 15 13 1 10 12 1 10 9 1 9 2
46 1 10 12 13 9 10 2 9 1 10 9 2 13 1 12 9 1 9 7 1 9 2 1 9 2 1 11 11 2 9 1 10 11 11 1 10 11 1 10 11 7 9 0 1 11 2
62 15 13 1 13 10 9 1 10 9 7 1 10 9 2 1 10 9 1 10 0 0 9 1 9 0 2 3 9 1 10 9 16 2 3 9 1 10 9 0 2 4 3 13 15 1 13 10 9 0 1 10 11 2 1 10 11 2 1 10 11 11 2
11 9 2 3 2 13 3 9 0 7 0 2
13 1 10 12 2 12 2 10 0 9 13 10 9 2
21 10 9 1 9 13 10 11 1 10 9 1 2 11 0 2 2 3 10 11 0 2
21 13 1 10 9 2 13 1 12 9 1 9 2 11 13 1 9 0 10 10 9 2
23 7 15 13 1 10 0 9 1 9 0 2 1 10 9 1 13 10 9 7 10 9 0 2
37 13 1 13 10 9 0 1 10 0 9 2 1 9 2 9 7 9 2 13 1 10 0 11 11 1 10 11 1 11 2 10 10 9 0 4 13 2
26 1 3 1 13 10 11 8 8 10 9 13 0 7 11 2 3 13 10 9 0 2 15 13 1 13 2
28 1 10 12 13 10 9 13 2 10 9 1 10 9 0 2 15 13 10 9 1 9 0 0 2 0 7 0 2
15 3 2 1 13 10 9 0 13 1 10 0 9 1 9 2
14 3 2 1 10 0 9 1 10 9 13 10 9 0 2
29 13 10 11 11 11 2 10 9 0 15 15 2 1 13 15 0 1 10 9 2 13 0 1 10 11 1 11 11 2
22 10 11 7 10 11 13 3 1 15 2 1 11 2 1 10 9 2 1 10 9 0 2
48 10 12 9 12 13 16 10 9 1 10 0 11 4 13 2 7 10 10 9 0 4 4 13 1 10 9 2 0 7 0 2 1 10 11 2 3 15 13 1 11 1 10 9 1 10 11 11 2
11 3 10 10 9 4 13 3 1 10 9 2
18 3 2 13 1 11 10 9 15 13 1 9 1 10 0 9 1 11 2
9 10 9 13 0 7 0 10 9 2
11 10 9 13 16 11 4 3 13 1 9 2
28 3 1 13 10 9 4 13 1 3 2 0 1 10 9 0 1 10 11 7 4 13 10 9 1 10 11 11 2
20 1 10 9 4 4 13 3 2 4 3 13 10 9 0 13 15 10 9 0 2
14 2 11 11 2 2 13 10 9 10 9 1 10 9 2
17 7 13 10 9 3 1 4 13 2 13 2 13 10 9 1 11 2
32 10 9 1 13 15 10 9 1 11 11 3 15 4 3 13 2 3 2 15 4 13 1 11 7 3 4 13 10 9 1 9 2
49 7 10 9 1 10 9 0 15 13 1 13 15 3 7 16 10 10 0 9 15 15 13 2 16 13 11 11 2 9 0 15 4 13 10 0 9 1 10 11 3 13 2 3 16 3 0 0 2 2
8 11 2 13 9 7 13 9 2
35 16 13 1 9 7 1 9 2 1 0 9 7 1 0 9 2 11 11 15 13 3 10 9 1 9 2 1 9 2 1 9 1 9 0 2
64 10 0 9 2 13 10 9 3 1 10 9 1 10 9 2 15 4 3 13 10 9 1 9 2 1 10 9 0 1 10 11 7 9 11 11 1 11 2 7 10 9 1 9 1 2 9 2 9 7 9 1 13 2 1 9 1 11 11 2 0 9 1 11 2
6 15 4 13 10 11 2
19 1 15 13 1 10 9 1 11 2 1 9 3 0 4 13 1 10 15 2
17 2 16 13 16 15 4 13 11 2 13 0 2 13 9 7 9 2
5 1 15 3 13 2
28 1 10 9 0 2 16 13 0 2 10 11 13 1 9 1 13 15 2 15 4 3 13 10 9 1 10 11 2
20 11 11 2 0 9 1 11 2 13 3 15 15 15 1 10 9 13 3 0 2
6 7 3 13 10 9 2
12 2 10 9 0 2 13 15 2 13 1 11 2
15 1 11 10 0 9 0 13 15 1 10 9 0 2 2 2
9 11 3 3 13 10 9 1 13 2
22 2 15 13 0 2 15 13 2 7 13 10 9 1 9 0 7 1 9 1 10 9 2
9 11 4 13 9 0 1 10 9 2
8 9 2 9 2 9 1 13 2
16 3 10 9 4 13 10 9 0 2 15 4 13 3 1 15 2
8 3 15 4 3 13 10 15 2
10 10 9 15 1 10 11 4 13 0 2
39 1 10 0 2 0 9 1 10 9 0 1 10 9 16 10 11 13 10 9 7 2 3 2 10 9 2 4 3 13 1 10 9 1 9 1 10 9 0 2
14 9 0 2 15 4 13 3 1 10 9 1 10 9 2
31 3 16 10 11 15 15 4 13 3 1 15 2 1 13 10 9 2 16 4 13 1 13 13 15 2 10 9 1 11 2 2
13 7 11 1 10 9 13 0 2 7 13 0 9 2
41 2 3 13 0 2 15 13 10 9 1 10 9 11 2 16 11 13 3 0 2 16 4 13 9 7 9 7 3 15 15 13 1 13 0 9 15 13 10 9 0 2
13 4 13 3 15 1 10 9 16 13 1 10 9 2
22 1 9 1 10 9 9 1 11 15 11 4 13 1 10 10 9 1 2 9 0 2 2
26 11 3 1 10 9 2 1 10 9 1 9 2 1 10 9 1 10 9 2 3 2 3 15 13 3 2
12 1 15 10 9 13 15 2 7 3 2 0 2
14 1 10 9 2 3 13 10 0 9 16 13 10 9 2
22 3 2 16 13 1 9 2 16 10 9 15 13 15 4 3 13 1 13 10 9 2 2
29 7 16 1 11 11 13 10 9 1 9 0 0 1 13 7 1 13 2 10 9 0 2 1 10 9 2 15 13 2
6 2 15 13 1 11 2
17 2 3 15 15 13 1 15 2 7 1 15 15 13 3 2 2 2
3 7 13 2
35 2 3 3 0 3 13 10 9 1 10 9 2 15 3 13 9 3 1 10 9 1 11 16 10 10 9 13 1 10 9 1 10 11 2 2
12 13 15 2 3 2 11 13 1 9 10 9 2
9 2 9 1 10 9 1 10 9 2
18 16 13 10 9 1 2 11 2 2 2 7 1 15 2 6 2 2 2
26 3 2 3 11 3 13 3 1 9 2 10 9 1 10 11 4 13 2 15 13 16 15 13 2 2 2
19 2 13 3 1 13 15 13 1 10 9 11 2 3 15 4 13 2 2 2
8 2 10 11 13 10 11 2 2
5 11 11 13 0 2
14 2 15 13 9 3 16 15 13 1 10 0 9 2 2
30 11 2 15 15 13 10 11 2 7 3 13 16 13 3 0 13 0 7 0 10 0 11 11 7 10 0 11 11 11 2
18 3 11 11 15 13 3 2 3 13 1 10 9 12 9 1 9 0 2
38 6 2 3 13 3 9 1 9 2 3 10 9 0 9 1 10 9 11 13 1 9 2 1 9 1 10 9 15 13 0 2 0 7 2 3 2 0 2
26 13 11 11 2 13 1 11 7 9 16 4 13 12 9 0 1 11 2 1 10 9 0 1 10 9 2
41 11 11 1 10 9 1 10 11 4 13 1 15 2 2 0 2 0 2 0 1 11 2 2 7 3 10 11 13 1 9 2 16 13 10 11 2 1 13 10 11 2
51 15 2 3 2 13 10 9 1 9 13 7 3 16 10 9 11 13 2 16 3 15 13 2 16 13 10 9 2 3 2 2 2 16 12 9 15 13 1 9 2 15 13 3 1 10 9 1 10 12 2 2
14 4 13 11 11 1 10 11 11 1 10 9 1 11 2
21 10 11 2 10 11 11 11 7 10 10 0 11 15 4 13 16 4 13 15 15 2
14 15 4 13 2 10 11 4 13 1 10 9 2 2 2
6 3 13 3 10 9 2
16 15 3 15 4 3 13 16 10 11 3 15 4 13 1 11 2
11 15 4 13 3 1 15 2 13 16 13 2
17 16 13 15 13 10 9 1 9 1 10 9 1 9 9 2 2 2
3 15 13 2
9 2 15 13 9 1 10 9 11 2
14 13 1 15 13 10 9 1 10 9 1 10 9 0 2
14 1 3 4 13 9 2 15 4 13 1 10 10 9 2
18 15 4 3 13 10 9 2 7 15 4 13 10 9 1 10 10 9 2
30 13 10 9 1 11 2 3 13 1 15 7 15 13 2 13 1 10 9 1 10 9 2 13 9 0 3 1 15 2 2
10 1 10 9 15 4 13 1 11 11 2
12 1 10 15 2 4 13 10 9 1 10 9 2
24 15 10 11 3 15 13 2 7 3 13 3 11 11 2 15 3 15 4 13 3 1 10 9 2
3 15 13 2
11 2 15 15 13 3 0 2 10 9 2 2
7 3 4 13 10 11 2 2
5 15 4 13 0 2
20 3 15 13 2 15 13 16 1 10 9 10 11 4 13 1 13 15 1 15 2
9 2 0 11 2 13 3 0 2 2
30 3 2 1 10 9 7 10 15 2 10 9 1 10 9 3 13 3 0 7 10 9 0 13 1 10 9 1 11 3 2
14 2 3 13 0 2 15 13 10 0 9 1 10 11 2
5 10 9 15 13 2
32 3 13 9 10 16 2 1 13 13 10 0 9 15 13 1 9 2 10 9 1 10 9 0 2 15 4 13 1 10 9 2 2
40 13 2 11 2 1 11 13 15 2 10 9 15 13 3 16 13 1 10 11 2 13 1 13 10 9 7 13 0 2 10 11 0 15 4 13 3 10 9 2 2
7 3 13 3 13 1 9 2
13 2 1 10 9 3 3 2 15 4 13 3 0 2
34 10 9 1 10 9 4 13 1 10 9 3 16 13 0 2 15 13 10 9 1 9 0 15 13 3 10 3 2 10 9 13 3 0 2
14 1 15 1 9 13 3 1 9 1 9 1 10 11 2
10 6 2 3 16 11 13 10 0 9 2
17 10 0 9 2 1 10 10 9 0 2 15 4 13 15 2 2 2
2 3 2
9 2 15 15 4 13 1 10 9 2
33 2 1 9 0 7 0 15 13 10 0 9 1 1 10 9 15 13 3 1 10 9 7 15 15 13 1 9 1 10 10 9 2 2
15 15 15 4 13 3 7 15 4 13 1 13 15 10 9 2
5 15 15 4 13 2
11 2 3 3 15 13 2 2 15 4 13 2
23 3 2 1 13 1 10 9 7 1 10 9 1 13 9 2 13 16 11 11 13 3 9 2
27 10 9 13 10 9 1 10 9 1 9 3 0 7 3 3 0 2 16 13 1 10 13 15 1 1 15 2
8 3 13 11 11 7 11 2 2
9 3 15 13 9 2 15 4 13 2
18 6 2 10 9 1 10 11 1 10 11 3 13 10 9 1 10 9 2
5 0 11 2 2 2
7 2 15 15 4 3 13 2
14 3 2 16 15 13 1 13 10 0 9 3 15 13 2
27 15 13 16 13 2 13 13 10 9 2 3 16 13 10 0 9 1 13 15 1 9 1 9 1 10 11 2
11 3 15 3 13 3 9 1 10 9 11 2
2 6 2
31 13 16 1 11 10 11 13 1 13 15 13 9 7 2 16 13 1 13 10 9 2 13 10 9 1 13 3 10 11 2 2
15 7 10 11 13 1 9 10 10 9 1 10 11 11 2 2
10 2 1 10 9 1 10 11 3 13 2
12 4 13 1 9 10 1 10 9 1 10 9 2
6 3 15 4 13 2 2
20 9 1 10 9 1 10 9 9 2 13 2 2 10 9 15 13 1 11 12 2
2 11 2
2 13 2
39 11 2 9 2 13 2 1 9 2 0 2 11 11 15 13 7 13 0 1 13 7 13 10 2 9 2 3 3 1 10 9 0 7 3 3 1 9 0 2
26 9 1 10 9 2 10 9 1 10 11 12 1 10 15 4 4 13 2 1 9 0 0 2 11 11 2
28 10 15 2 13 11 2 13 3 0 2 7 1 2 9 2 2 1 10 9 16 4 13 9 1 10 11 0 2
31 10 9 13 1 10 9 16 10 11 12 3 4 13 10 2 9 2 2 3 10 9 15 13 10 2 9 2 1 10 9 2
12 7 3 2 3 2 13 2 3 10 9 9 2
28 13 15 3 10 9 2 3 0 2 3 0 2 1 9 15 15 4 13 7 15 4 3 13 1 10 9 0 2
8 1 11 3 15 13 9 10 2
24 2 9 2 3 2 3 16 10 9 0 1 10 9 1 9 4 2 13 2 1 10 9 0 2
3 10 9 2
2 0 2
3 13 0 2
47 2 6 2 7 3 10 10 9 16 13 10 9 1 11 11 2 0 9 0 1 10 9 11 2 9 2 3 4 13 15 2 2 15 13 2 0 2 11 11 2 9 1 10 11 12 2 2
9 3 2 0 9 1 10 11 2 2
32 10 9 1 10 13 9 3 13 3 15 1 2 13 2 10 9 2 3 16 2 15 13 2 4 13 1 15 15 13 3 2 2
17 10 9 13 16 10 9 13 1 13 0 2 10 9 11 13 0 2
22 3 2 10 9 4 4 13 3 2 7 13 1 15 16 15 13 0 9 1 10 9 2
23 7 3 3 15 13 3 9 2 0 2 2 3 15 13 3 15 15 13 3 0 1 15 2
9 15 4 13 3 1 10 0 9 2
23 7 16 3 13 1 13 10 9 2 13 3 12 9 1 10 0 9 2 7 13 1 9 2
22 3 2 16 13 13 10 9 9 1 9 2 3 4 13 1 13 3 15 1 9 2 2
16 3 2 1 10 9 2 13 1 9 7 10 9 15 13 2 2
12 11 11 2 9 1 10 11 12 2 15 13 2
2 13 2
14 2 1 10 9 15 13 3 0 2 13 3 13 2 2
10 13 10 9 1 10 10 9 11 11 2
5 15 3 13 9 2
13 2 10 11 12 13 2 10 2 9 2 15 13 2
6 16 13 0 2 3 2
11 11 11 2 9 11 12 2 3 15 13 2
10 2 7 16 4 15 13 2 3 13 2
7 13 13 0 1 10 9 2
22 7 15 1 10 11 12 15 13 1 13 10 9 2 16 15 13 3 3 13 2 2 2
10 13 1 10 9 0 1 13 10 9 2
10 15 13 9 1 9 1 10 9 0 2
3 11 13 2
5 2 11 0 2 2
15 9 1 9 0 1 9 2 13 2 10 9 1 10 11 2
31 1 10 0 9 11 2 15 4 13 1 13 1 9 2 13 15 10 9 1 13 1 10 9 1 9 0 13 1 10 9 2
16 15 15 4 13 1 9 1 10 9 1 9 13 1 10 9 2
57 10 9 4 13 1 9 7 9 10 9 1 9 0 1 9 1 9 1 9 3 1 10 0 9 1 9 2 1 10 9 3 1 10 9 7 10 9 13 1 10 9 1 10 9 15 13 1 10 10 9 0 1 9 0 7 0 2
9 2 4 13 10 10 9 1 15 2
33 13 10 9 2 2 13 11 11 2 12 9 2 15 1 10 12 4 13 10 0 9 1 9 2 13 1 10 9 1 10 9 0 2
8 2 13 10 0 9 1 9 2
17 3 4 4 13 2 7 10 3 3 4 13 1 13 10 10 9 2
10 7 3 16 13 1 9 15 4 13 2
30 3 3 13 1 11 2 2 13 11 11 2 10 9 1 10 9 0 2 10 9 1 9 7 10 9 13 1 10 9 2
22 1 11 10 9 15 4 13 11 11 2 1 15 1 10 9 1 10 9 1 10 11 2
44 7 3 9 1 2 13 15 2 1 15 1 11 2 10 0 0 9 1 10 11 7 0 9 0 2 4 13 10 9 1 10 9 2 0 1 13 1 9 10 9 1 10 9 2
13 7 15 0 1 13 1 3 12 9 3 4 13 2
93 10 9 3 16 10 9 0 4 13 10 0 9 0 2 7 16 1 9 13 3 10 9 2 0 2 15 13 10 9 0 1 10 9 0 2 10 0 9 1 0 9 1 11 4 13 1 13 15 3 1 10 0 9 2 1 9 1 9 0 1 10 9 3 13 1 10 9 2 1 9 0 1 9 15 13 1 13 10 0 9 7 1 9 1 9 15 13 15 13 3 10 9 2
24 2 15 13 9 13 2 15 13 10 9 1 11 3 3 1 3 9 15 3 4 3 13 9 2
21 13 0 2 13 0 2 2 13 11 2 15 13 1 9 10 0 9 0 0 0 2
14 10 9 13 1 9 0 2 7 10 9 13 3 0 2
22 7 10 9 1 11 4 13 1 10 9 1 13 1 11 7 1 10 0 9 3 13 2
33 2 3 4 3 13 10 10 9 16 10 9 15 4 13 1 0 9 15 15 4 13 1 10 9 2 2 4 13 10 9 11 11 2
46 7 3 1 10 9 1 10 9 2 1 13 10 11 13 3 10 9 1 9 4 13 1 10 9 0 2 3 10 9 13 0 2 10 9 1 10 9 9 2 10 9 1 15 13 0 2
31 13 10 9 0 2 10 11 2 0 7 0 2 1 10 9 11 11 15 4 13 1 10 9 1 10 9 1 10 0 9 2
51 7 3 10 0 9 1 9 0 2 1 9 1 10 9 15 13 1 13 9 1 10 9 1 0 9 1 9 7 13 3 1 9 1 4 13 2 13 1 10 9 1 9 1 13 3 1 10 9 1 11 2
14 13 10 9 0 2 3 3 10 9 4 13 1 13 2
18 10 9 4 13 1 9 2 1 10 9 0 15 13 10 9 1 9 2
16 2 3 4 13 0 10 9 0 7 3 4 13 10 0 9 2
23 1 10 10 9 0 1 9 0 1 10 11 4 13 10 9 7 10 9 1 10 10 9 2
38 16 3 4 13 9 1 9 4 13 2 2 13 10 9 11 2 15 13 1 0 9 10 9 13 1 10 9 1 10 9 0 3 13 1 0 12 9 2
12 2 10 11 3 13 3 2 2 13 10 9 2
16 1 3 1 10 9 10 9 13 1 13 10 0 9 1 9 2
15 3 9 4 4 13 3 11 2 1 10 9 1 10 11 2
27 10 9 0 1 10 9 1 11 2 15 1 10 2 9 2 0 13 1 10 11 2 4 13 1 9 0 2
13 7 10 9 11 2 15 4 13 11 2 4 13 2
15 2 3 13 3 13 10 9 1 10 11 0 7 0 2 2
9 1 10 9 15 13 10 0 9 2
28 10 9 13 2 10 9 1 9 0 15 13 1 10 9 7 13 2 1 10 9 1 10 9 15 13 10 9 2
30 7 1 10 9 15 13 1 11 2 1 10 3 0 11 2 9 1 9 4 13 1 10 9 1 10 9 1 10 9 2
23 13 10 9 0 1 10 9 15 4 4 13 10 3 9 1 3 10 12 9 3 4 13 2
15 2 15 13 10 9 1 10 9 2 2 13 10 9 0 2
29 7 3 10 0 11 2 10 9 1 11 2 4 13 3 1 13 1 0 10 0 2 9 2 1 11 7 1 11 2
21 10 9 13 3 16 10 9 3 4 13 2 7 3 4 13 2 13 10 9 0 2
14 10 0 9 1 10 9 1 11 4 13 10 9 0 2
13 2 10 0 9 1 11 15 4 13 1 10 9 2
10 3 13 3 1 11 2 2 13 11 2
28 2 3 4 3 13 1 13 15 1 9 2 2 13 10 9 15 4 13 3 1 11 1 10 9 1 10 9 2
11 10 10 9 4 3 13 1 9 10 9 2
9 10 0 9 15 13 10 9 0 2
12 2 13 1 10 9 1 10 9 2 2 13 2
6 10 9 1 10 9 2
9 1 9 7 9 10 9 1 11 2
8 2 3 13 1 13 11 2 2
56 1 10 0 9 11 2 10 9 13 10 9 7 13 10 9 1 9 2 1 10 9 13 10 9 0 7 1 10 9 10 9 13 1 10 9 1 11 2 13 1 10 9 7 13 1 10 9 3 13 1 12 9 1 10 9 2
29 15 13 16 15 13 7 10 9 3 0 1 10 9 2 1 9 2 1 9 13 13 1 9 7 3 1 10 9 2
45 3 11 2 12 9 2 15 1 10 9 15 4 13 1 10 0 9 1 2 0 2 9 0 1 10 9 0 2 4 13 1 13 15 1 10 0 9 1 11 2 7 4 13 3 2
11 2 4 13 3 1 10 12 2 13 2 2
3 13 0 2
15 0 13 16 13 10 9 1 9 1 3 4 13 1 13 2
37 4 4 13 15 3 3 1 0 2 1 10 10 9 2 13 15 3 1 11 16 10 9 15 13 1 11 2 10 10 9 2 1 12 9 1 11 2
3 7 13 2
15 15 4 3 13 10 9 0 0 1 10 0 2 9 2 2
5 10 9 1 11 2
10 13 3 1 10 9 2 1 10 9 2
21 13 0 2 3 2 7 1 9 10 15 13 10 0 9 16 13 3 1 10 9 2
14 13 3 0 2 13 10 9 1 9 2 3 1 9 2
8 7 15 15 13 3 1 9 2
19 15 2 1 9 2 13 1 10 9 15 13 2 16 15 13 1 13 3 2
5 15 3 2 2 2
19 10 9 1 10 9 13 1 11 1 13 10 9 0 0 1 11 7 11 2
18 7 2 3 2 1 13 1 10 0 9 1 10 9 10 0 9 0 2
14 2 4 13 15 3 2 13 11 2 3 15 4 13 2
10 10 9 1 11 2 10 15 1 11 2
28 15 4 13 1 13 1 13 10 10 9 2 11 2 7 16 15 4 13 4 13 1 11 1 13 10 10 9 2
17 2 9 2 9 2 15 4 13 11 2 3 4 13 1 9 2 2
8 10 15 4 13 1 9 2 2
5 15 13 2 11 2
11 13 10 9 7 13 10 9 2 1 9 2
9 2 13 15 13 10 9 2 2 2
12 3 16 15 13 2 11 11 2 11 10 11 2
3 2 9 2
14 6 2 6 2 6 2 13 11 2 6 2 3 9 2
6 10 9 13 10 9 2
14 4 13 15 2 10 0 9 2 16 13 16 15 13 2
11 13 1 9 2 7 15 3 15 4 13 2
9 1 15 4 13 0 16 13 3 2
9 7 13 0 16 3 13 3 2 2
36 10 9 1 9 1 9 1 9 1 10 9 0 2 10 9 1 3 2 11 13 10 9 1 10 15 15 15 13 1 13 15 3 3 1 9 2
15 13 15 15 1 9 1 9 4 13 15 1 13 10 9 2
28 16 13 10 9 0 2 1 13 16 13 1 13 9 1 10 9 2 13 10 9 0 1 13 1 0 10 9 2
21 2 6 2 6 2 6 2 13 3 11 2 16 3 13 3 3 4 13 1 9 2
27 7 10 9 2 3 15 0 2 13 16 15 13 1 13 1 10 9 7 1 10 9 2 7 3 2 2 2
26 3 16 16 15 13 1 15 2 1 10 9 13 1 9 2 13 1 10 9 0 1 10 11 11 2 2
10 3 2 15 3 13 10 9 1 11 2
31 6 2 15 1 9 1 15 4 13 11 7 11 16 1 12 9 3 15 4 4 13 2 7 3 3 13 13 15 10 9 2
11 7 3 15 13 10 9 0 1 10 9 2
5 15 13 10 9 2
14 13 15 13 10 10 9 0 16 13 1 10 9 0 2
6 13 1 10 9 0 2
11 1 11 2 10 11 2 7 3 10 11 2
2 3 2
3 10 11 2
6 6 2 3 10 11 2
17 13 1 10 10 9 1 11 7 13 15 2 6 2 6 6 2 2
19 13 10 9 1 10 9 1 11 2 13 3 11 2 1 13 15 13 3 2
24 10 0 9 15 15 4 13 13 2 1 0 9 2 10 9 1 9 2 0 2 1 10 9 2
3 1 13 2
12 1 13 2 3 1 10 9 2 3 10 9 2
27 2 1 9 2 15 13 1 10 9 10 9 11 2 15 4 13 10 11 1 13 15 1 2 13 15 2 2
10 15 13 10 9 1 4 13 1 15 2
9 15 1 11 7 11 7 11 2 2
6 6 2 13 1 11 2
8 3 15 13 0 9 2 2 2
8 12 9 13 13 1 10 9 2
6 9 1 10 11 0 2
8 2 3 13 1 13 15 2 2
8 9 2 9 0 1 10 9 2
6 10 11 13 10 9 2
12 2 11 0 13 1 9 0 1 10 9 2 2
32 1 10 0 9 11 2 10 2 9 1 9 0 2 4 13 3 10 9 2 13 10 10 9 1 10 10 9 1 10 0 11 2
16 0 9 1 9 1 9 15 4 13 1 10 9 1 10 9 2
34 7 1 10 9 0 1 10 11 10 0 9 1 10 9 1 10 12 13 3 10 9 2 0 1 13 1 11 7 1 11 2 0 2 2
18 7 13 10 0 9 1 10 9 15 10 9 13 1 3 10 9 0 2
33 1 10 9 0 1 10 11 11 13 12 12 10 9 1 9 1 10 9 1 10 11 0 2 3 1 10 2 9 2 0 11 11 2
20 10 9 1 11 2 3 2 13 16 13 2 3 2 12 12 10 9 1 9 2
15 1 11 10 9 0 13 16 10 9 13 1 12 12 9 2
20 10 0 9 1 10 11 1 10 0 9 0 2 7 13 1 15 10 9 0 2
29 15 13 10 9 1 9 2 10 9 0 13 16 4 4 13 7 13 3 10 9 1 9 0 1 10 9 3 13 2
12 2 4 13 1 10 10 9 1 11 1 13 2
10 4 13 15 10 9 1 10 10 9 2
18 10 9 4 13 3 10 10 9 2 2 13 10 9 1 10 11 0 2
39 2 3 4 13 1 13 3 1 15 15 13 10 9 1 9 7 3 4 13 9 1 10 9 13 1 10 9 1 9 1 10 9 0 2 2 13 3 11 2
27 1 10 9 3 15 13 9 1 9 13 1 10 9 13 1 11 7 1 11 12 9 3 1 13 10 11 2
11 13 10 11 1 4 13 10 9 3 0 2
30 9 0 0 4 4 13 1 10 9 1 10 9 1 9 0 7 13 1 0 9 1 9 0 1 9 1 10 9 0 2
24 10 9 1 11 13 3 7 13 1 2 13 10 9 2 16 4 13 1 10 9 1 10 9 2
14 10 9 1 10 11 1 11 2 11 11 2 3 13 2
14 2 4 13 12 9 1 10 9 1 10 0 9 2 2
28 10 0 9 1 10 11 1 10 9 2 11 2 13 1 2 0 9 0 2 1 9 1 10 9 1 10 9 2
6 2 13 16 13 9 2
35 10 9 4 13 3 0 16 15 13 1 10 10 9 7 4 13 10 9 0 2 2 13 11 11 1 10 9 1 11 11 1 10 11 11 2
19 13 10 9 0 2 3 16 10 9 4 4 13 1 9 1 10 9 0 2
18 3 13 15 1 15 2 2 13 11 11 2 9 1 10 11 1 11 2
33 1 10 9 2 1 10 9 1 10 0 11 7 10 11 0 15 4 13 10 9 1 12 9 1 9 2 15 1 9 15 1 9 2
8 1 1 15 15 13 10 9 2
10 3 1 11 11 4 13 12 12 9 2
21 1 1 15 15 13 9 1 9 2 9 7 0 9 0 1 10 9 1 10 9 2
13 10 12 12 9 4 13 3 11 2 1 10 11 2
18 10 11 13 1 4 13 12 9 1 9 15 10 9 4 13 1 9 2
14 7 3 13 3 15 15 13 1 10 9 1 10 9 2
19 10 11 0 13 10 9 0 7 3 10 9 1 13 10 0 9 1 9 2
14 7 3 10 11 11 3 13 10 9 1 13 10 9 2
12 1 10 9 0 10 9 13 15 1 9 0 2
42 3 1 10 11 0 2 13 0 1 10 9 7 3 1 9 0 2 15 4 13 10 9 1 10 0 9 1 10 9 7 10 9 15 4 3 13 1 9 1 10 11 2
13 1 11 13 10 9 1 3 1 10 9 3 0 2
29 10 9 1 10 11 0 2 3 2 4 13 1 13 3 9 7 9 7 1 13 1 9 7 9 1 13 10 9 2
21 2 3 3 13 3 3 0 2 16 15 13 10 9 4 13 15 2 2 13 11 2
10 10 9 0 1 10 9 4 13 0 2
32 3 1 11 11 4 13 12 9 7 12 9 2 7 3 10 12 12 2 9 0 2 1 10 11 0 4 4 13 10 10 9 2
8 1 15 3 15 13 3 9 2
8 11 13 2 13 10 9 2 2
33 11 2 11 0 1 11 4 13 1 13 10 9 1 10 9 11 1 11 7 10 9 1 9 11 11 11 13 1 10 9 1 3 2
38 2 1 0 9 1 9 1 10 10 9 7 10 9 13 1 10 0 9 1 10 9 1 10 0 11 13 1 10 0 9 1 10 11 1 10 9 2 2
70 15 2 4 13 1 10 9 1 11 2 2 3 13 13 9 1 15 1 10 9 1 9 2 7 13 10 0 9 1 9 1 10 9 15 13 3 10 9 0 2 1 15 2 1 9 1 9 2 0 9 4 13 1 10 9 1 10 0 9 0 1 15 1 10 9 1 9 2 2 2
65 15 13 3 0 2 13 10 9 2 16 1 10 9 0 0 13 3 1 9 3 1 0 9 2 7 3 1 13 10 10 9 2 16 10 10 9 1 10 9 2 10 9 7 10 9 0 2 3 1 13 10 0 9 2 4 13 9 0 2 13 9 7 9 2 2
3 10 9 2
8 7 11 15 13 1 10 9 2
10 2 4 13 15 2 7 4 13 2 2
37 1 10 0 9 11 2 10 9 13 0 1 10 9 1 10 9 0 2 15 4 13 3 1 3 2 1 12 9 2 10 9 0 1 10 9 0 2
36 9 0 13 1 11 1 11 2 2 9 2 1 10 0 9 2 3 10 10 9 2 11 2 4 13 1 10 9 15 13 10 9 2 0 2 2
41 3 13 0 10 9 1 13 15 2 10 9 3 2 1 10 9 2 3 16 10 9 3 4 13 1 10 9 11 7 10 9 13 3 1 9 1 10 9 1 9 2
56 9 9 4 13 10 9 1 9 1 10 9 0 2 10 9 1 9 11 13 0 2 10 9 7 10 9 13 11 1 10 9 3 7 1 9 1 10 9 2 16 4 13 3 1 12 9 2 15 13 2 2 0 1 10 9 2
11 13 16 4 15 13 2 1 10 9 0 2
9 15 13 13 1 10 9 7 13 2
6 2 3 15 13 2 2
3 13 9 2
12 2 6 2 9 2 15 13 10 9 11 2 2
9 4 13 0 10 9 1 10 11 2
6 2 13 3 1 3 2
14 10 9 1 10 9 2 10 9 0 2 13 10 9 2
10 10 9 4 13 1 11 1 10 9 2
31 2 10 9 2 13 10 9 0 2 13 1 10 9 3 1 10 9 1 9 1 9 2 2 15 13 1 11 1 10 9 2
25 10 10 9 13 0 2 7 15 13 3 10 9 7 10 9 2 1 10 9 3 15 15 13 15 2
18 10 9 1 11 3 13 1 9 1 10 9 7 1 10 11 0 0 2
14 13 16 13 10 10 9 2 7 15 3 15 15 13 2
8 3 10 9 15 4 13 2 2
8 4 13 11 2 4 13 11 2
11 10 9 0 13 1 9 2 10 9 0 2
27 9 3 13 0 10 9 2 9 1 9 2 1 9 1 11 7 11 1 10 9 0 0 1 11 7 11 2
22 3 15 13 9 1 9 1 9 1 11 11 1 10 9 7 1 10 9 1 10 11 2
21 9 2 10 15 7 10 15 2 1 9 0 13 1 9 1 10 9 1 10 9 2
22 10 9 7 10 9 1 10 9 11 13 1 9 3 1 10 12 2 16 13 10 9 2
34 7 10 9 13 0 7 15 13 10 9 3 0 2 10 9 0 1 9 2 10 9 1 9 7 10 9 16 4 13 1 13 10 9 2
3 9 0 2
34 10 9 1 9 9 2 12 9 7 12 9 2 9 0 7 0 2 15 13 1 0 7 1 0 2 1 10 9 7 10 9 3 0 2
21 11 2 10 9 0 3 0 15 4 13 10 9 1 10 9 1 11 2 13 0 2
15 13 1 10 10 9 2 3 1 10 11 11 1 9 0 2
14 9 2 1 10 11 11 2 13 10 9 1 10 9 2
14 7 10 9 2 1 9 1 9 0 2 13 10 9 2
26 15 13 10 9 13 0 1 13 16 3 13 10 9 1 4 13 1 11 10 0 2 0 9 1 9 2
33 15 15 13 16 10 9 0 3 4 3 13 1 10 0 9 0 1 10 9 1 13 10 9 15 13 10 9 1 9 1 10 9 2
31 10 9 4 13 3 10 9 0 7 0 2 16 13 1 10 9 1 13 0 1 13 15 10 9 1 10 9 1 10 9 2
51 10 9 1 9 0 15 15 4 13 2 1 10 0 9 2 10 2 11 12 2 2 10 9 1 9 0 13 1 10 9 1 10 9 2 15 4 4 13 10 0 2 2 0 2 9 1 10 9 1 11 2
24 15 13 9 12 9 1 10 11 1 10 11 2 12 9 0 2 9 2 9 2 9 2 9 2
28 10 9 13 1 10 9 1 11 3 12 9 0 4 13 10 9 0 1 11 7 13 10 9 1 10 9 0 2
19 15 1 10 9 15 13 0 1 10 2 9 2 1 10 9 0 1 11 2
26 2 15 13 3 2 13 2 16 15 1 15 15 13 1 9 7 15 13 9 1 11 11 1 11 2 2
20 3 10 9 15 13 1 10 9 0 2 15 2 1 9 0 2 4 4 13 2
38 4 13 9 1 10 9 11 2 15 1 10 10 9 0 13 3 10 9 1 10 9 1 10 11 11 2 11 11 2 7 10 9 1 10 9 2 11 2
27 2 15 13 10 11 0 2 13 15 1 10 2 11 12 2 2 2 3 13 10 9 1 10 9 0 2 2
22 15 13 1 9 2 15 4 13 1 10 11 2 13 1 10 9 2 10 9 3 0 2
32 1 10 15 3 15 4 13 10 9 1 10 9 1 10 9 2 1 9 0 2 1 10 9 2 7 13 15 1 10 9 0 2
13 2 10 9 2 13 13 2 13 10 9 0 2 2
21 13 0 13 16 10 9 2 13 3 3 2 13 15 15 13 1 9 1 10 9 2
15 10 0 2 0 9 2 7 10 0 9 1 10 9 0 2
7 10 9 13 3 2 0 2
7 10 9 1 11 1 11 2
8 7 10 9 13 1 10 9 2
6 11 2 9 1 9 2
12 7 11 2 13 2 10 9 1 10 9 0 2
13 9 1 10 0 9 1 10 9 1 10 0 9 2
10 10 11 0 1 2 9 1 9 2 2
12 1 10 9 0 13 10 9 1 10 0 9 2
34 1 11 2 2 9 2 1 10 9 1 11 2 10 2 9 2 11 11 7 10 9 11 11 15 4 13 1 10 9 1 10 0 9 2
7 10 9 1 3 13 0 2
51 10 9 1 9 15 4 13 1 11 2 16 10 2 9 2 1 11 13 1 11 2 15 9 4 13 1 15 10 9 0 1 10 9 0 0 2 13 11 1 10 2 9 2 1 10 9 1 11 7 11 2
25 10 9 0 1 9 0 16 15 13 16 10 11 13 3 0 2 13 1 10 9 1 10 9 0 2
13 7 3 12 9 1 10 9 0 15 4 13 9 2
63 13 1 11 11 2 1 10 11 1 10 11 2 10 12 9 4 13 10 9 1 10 9 15 13 2 10 9 2 1 11 2 10 9 0 1 10 9 1 10 9 1 10 10 9 2 1 10 10 9 2 1 10 10 9 7 1 10 10 9 1 13 2 2
9 7 1 13 10 0 9 1 11 2
13 2 15 13 3 10 9 1 10 10 9 11 2 2
17 7 3 9 10 9 0 4 2 13 1 9 2 10 9 1 11 2
23 1 9 1 10 0 9 1 11 7 1 10 10 9 2 11 4 13 1 13 10 9 0 2
9 2 13 16 13 10 9 0 2 2
52 7 10 10 9 13 16 1 11 4 13 1 10 9 1 10 9 11 11 2 10 9 1 11 0 9 1 10 2 9 0 2 7 3 13 1 13 10 9 0 15 13 1 9 1 11 10 9 1 10 9 0 2
32 13 10 9 1 11 2 10 9 0 15 3 4 13 13 10 0 9 1 10 11 11 2 3 11 13 10 9 1 13 15 15 2
37 15 13 16 11 4 3 13 1 13 9 0 1 11 1 11 1 9 1 10 11 0 2 10 9 0 1 10 9 1 10 11 0 1 10 9 0 2
15 7 3 9 10 11 0 4 13 2 10 9 1 9 2 2
37 3 10 0 9 11 11 2 9 1 11 2 4 13 1 10 11 11 11 16 2 10 0 9 1 9 13 10 9 1 11 1 10 9 1 9 2 2
24 7 4 4 13 3 10 9 1 11 11 2 2 9 2 1 10 0 9 0 0 2 10 11 2
24 10 9 0 4 13 9 1 15 11 4 4 13 16 13 1 13 7 3 15 4 13 10 9 2
8 3 11 13 3 0 1 11 2
16 10 9 1 10 9 2 3 13 2 13 10 9 1 10 9 2
10 13 10 9 10 9 13 1 10 9 2
34 11 2 1 10 12 0 1 10 9 0 1 11 13 3 3 1 12 10 9 13 1 10 9 1 10 11 1 9 1 10 9 0 0 2
25 1 15 2 13 1 10 9 2 15 13 10 9 1 11 11 2 10 9 1 10 9 0 1 11 2
47 11 11 2 9 1 10 11 11 2 15 13 10 9 7 1 11 2 7 1 11 2 4 13 10 9 1 15 10 9 9 1 10 9 1 11 4 13 1 10 9 3 10 9 1 9 0 2
29 11 13 10 0 9 1 10 9 2 15 2 1 10 9 2 13 1 13 1 0 9 7 9 10 9 1 10 9 2
16 10 0 9 0 0 15 13 1 12 10 9 0 1 10 11 2
42 10 9 2 1 9 1 10 9 0 2 1 10 9 1 11 11 2 15 13 10 9 1 10 10 9 3 1 11 7 3 3 1 10 9 2 10 11 1 10 11 2 2
16 10 9 1 9 1 10 9 0 1 15 13 10 10 9 0 2
44 10 9 1 15 12 9 3 10 9 0 1 10 9 11 13 1 9 10 9 1 11 11 13 1 10 0 9 2 13 1 10 9 1 10 9 2 10 9 1 10 9 1 11 2
44 1 9 10 0 9 0 0 0 1 10 9 1 9 13 1 10 9 2 10 0 9 1 9 13 10 9 13 1 10 9 1 10 3 16 10 9 4 13 10 9 1 10 9 2
57 1 10 0 9 13 10 9 0 2 15 3 3 13 10 9 9 1 10 9 12 2 13 3 0 7 13 1 13 1 11 7 3 1 11 1 10 11 2 13 10 9 0 1 11 2 11 2 2 11 2 11 7 11 2 11 2 2
64 13 3 0 2 0 7 0 1 10 11 2 13 16 10 9 3 3 2 15 1 11 11 1 10 11 9 0 2 13 12 9 1 11 7 16 9 1 11 2 1 15 10 9 13 1 10 9 1 12 10 9 11 11 1 11 7 11 2 13 3 1 9 0 2
37 10 9 1 10 9 0 0 0 1 11 13 1 12 9 2 1 11 11 2 3 10 9 1 9 1 9 1 9 1 10 11 2 11 11 7 11 2
62 10 9 3 0 1 10 9 15 3 13 1 11 1 10 9 13 10 9 0 7 1 10 11 2 15 13 9 7 10 9 2 7 1 10 9 10 9 2 1 10 10 9 1 9 2 9 1 9 7 9 1 10 9 4 3 13 10 9 1 10 9 2
7 10 0 9 13 1 11 2
8 11 2 10 9 1 10 9 2
15 2 10 10 0 9 13 10 0 9 1 10 9 0 2 2
34 11 2 10 11 11 4 13 1 10 0 9 1 9 0 2 15 15 13 3 0 1 3 2 1 10 9 13 1 11 11 1 10 9 2
48 4 13 10 0 9 10 9 0 2 9 1 10 9 2 15 4 13 10 0 9 1 10 9 1 10 9 1 10 9 1 9 11 11 2 13 9 1 10 9 1 10 1 15 0 9 11 11 2
33 10 9 1 11 11 2 0 7 0 2 13 10 0 9 7 10 9 2 16 10 9 13 3 13 2 10 9 0 13 0 1 3 2
30 10 0 7 0 11 0 4 13 10 9 11 2 13 10 9 3 2 13 1 11 10 9 1 10 0 9 13 1 9 2
53 3 2 1 9 2 15 2 15 13 12 9 2 13 13 1 10 9 16 10 9 2 3 3 3 13 3 0 2 7 3 16 3 13 1 10 9 10 10 9 7 10 9 2 16 3 13 10 2 9 1 9 2 2
6 7 10 9 4 13 2
58 13 16 10 9 15 4 13 7 3 2 16 10 12 9 15 4 3 13 1 10 9 1 11 3 15 15 13 1 13 15 1 9 2 16 13 10 9 2 7 16 13 0 16 1 10 9 15 15 13 2 9 2 7 15 2 9 2 2
57 13 0 3 16 1 9 13 13 15 1 10 9 1 10 12 9 1 10 9 2 16 15 13 1 13 15 9 3 2 12 9 1 10 9 2 7 16 3 1 10 9 4 13 3 1 9 10 2 3 1 9 2 16 13 1 15 2
12 10 9 1 10 12 13 4 13 1 0 9 2
31 15 13 1 15 10 9 9 1 10 9 0 7 15 13 1 15 10 9 1 10 9 15 13 10 9 1 10 9 1 9 2
8 11 2 10 9 3 13 9 2
8 9 2 9 7 9 1 9 2
66 11 2 0 9 1 9 0 1 9 7 9 1 11 2 10 9 1 10 11 11 2 3 1 9 9 4 13 3 12 0 9 1 10 10 11 2 1 13 10 2 9 1 10 9 2 2 10 9 15 1 10 12 15 13 3 10 10 9 1 10 0 0 9 1 9 2
68 1 10 9 1 12 9 7 12 9 1 9 2 15 4 13 1 9 7 9 10 9 1 10 9 1 11 2 10 9 2 3 3 0 2 13 1 12 9 0 2 1 15 12 2 12 3 2 1 10 9 0 1 9 2 3 3 3 0 1 15 1 10 9 2 1 10 9 2
51 10 9 1 10 9 2 15 1 10 9 1 10 2 9 1 10 9 2 2 10 0 7 0 2 9 2 13 2 4 13 1 9 12 9 2 4 13 3 12 9 2 1 15 10 9 13 3 1 10 9 2
49 10 0 9 1 9 15 4 13 9 9 2 16 9 1 9 15 4 3 13 1 10 9 1 10 0 9 0 2 13 10 0 9 1 9 7 9 9 1 10 9 2 15 4 13 1 9 7 9 2
31 10 9 2 13 1 9 1 9 1 10 2 9 9 0 2 2 15 13 9 1 9 2 4 13 13 1 10 9 10 9 2
24 3 3 12 9 4 13 10 9 2 7 10 9 3 13 16 4 13 15 10 0 9 1 9 2
11 10 9 1 11 13 10 9 1 10 9 2
27 9 7 9 0 13 2 9 1 10 9 13 7 13 2 9 1 10 9 1 9 2 9 7 9 0 13 2
13 10 0 9 1 9 0 1 0 9 4 4 13 2
10 9 1 10 9 1 10 11 1 11 2
18 10 9 1 10 9 13 13 10 9 0 2 15 9 3 15 13 2 2
54 11 2 10 11 2 13 1 10 0 9 1 9 1 10 9 1 10 11 11 11 7 10 9 2 4 13 1 9 3 10 9 0 1 10 11 1 11 2 10 3 0 9 1 10 9 7 10 9 1 9 1 10 9 2
27 10 9 1 10 2 11 1 9 2 4 13 2 1 11 2 11 11 11 2 10 9 12 1 10 0 11 2
31 2 4 13 3 10 10 9 2 4 13 10 9 15 4 13 10 9 2 2 7 13 1 15 10 10 9 1 9 0 2 2
14 10 9 4 13 16 10 9 13 2 13 3 3 2 2
17 10 9 1 10 9 15 13 1 10 9 1 10 9 1 10 9 2
53 2 15 3 4 13 9 1 10 9 11 2 16 15 13 10 9 0 2 15 15 13 13 10 9 2 2 4 13 2 13 10 9 1 10 0 9 1 10 9 0 1 10 9 15 4 13 1 10 9 1 10 9 2
5 10 9 1 11 2
6 9 9 1 10 11 2
8 11 2 15 1 9 1 9 2
15 1 10 9 0 3 4 13 10 9 1 10 9 1 11 2
36 2 3 4 13 15 1 10 9 1 10 9 1 10 9 1 15 3 13 1 10 9 1 13 10 9 1 10 9 7 1 13 1 13 15 15 2
20 10 9 4 13 10 0 9 1 9 3 1 10 9 1 10 10 9 0 2 2
50 10 9 0 1 11 2 13 1 10 9 13 1 11 2 16 1 10 3 0 2 3 13 1 9 1 10 0 9 0 7 1 10 0 9 0 1 10 0 9 2 10 11 2 9 1 11 2 10 11 2
39 7 3 15 4 13 16 10 9 3 4 13 1 10 9 10 0 9 1 10 9 0 2 3 1 9 0 9 2 13 15 15 3 0 2 3 13 1 9 2
38 7 10 12 9 1 10 11 11 3 15 4 4 13 2 16 1 9 15 1 13 10 11 4 13 1 2 13 2 10 9 0 1 9 1 10 9 0 2
18 15 3 4 4 13 10 9 1 10 9 1 10 0 9 1 10 9 2
31 10 11 4 13 1 13 1 10 9 1 9 15 7 12 10 9 13 3 1 10 9 1 11 11 2 11 11 7 11 11 2
45 10 0 13 16 10 10 9 2 10 2 11 7 11 2 2 13 1 10 2 11 11 2 2 2 4 13 10 9 1 9 1 10 10 9 2 1 9 1 10 9 1 10 9 0 2
9 1 10 2 9 2 4 4 13 2
7 9 2 9 9 2 9 2
5 3 11 1 11 2
19 13 0 1 2 10 9 1 10 9 2 2 7 3 10 9 13 12 9 2
21 7 1 10 9 10 9 1 11 13 10 9 1 0 9 13 1 10 9 1 11 2
18 1 10 0 9 11 2 13 1 10 9 7 3 13 1 10 10 9 2
35 10 9 0 1 9 1 10 9 1 9 2 3 1 10 9 9 13 1 10 9 2 9 0 2 9 2 2 9 2 7 9 0 1 9 2
14 13 10 9 0 1 10 9 13 1 9 1 10 9 2
20 2 11 11 2 2 2 11 11 2 2 2 11 11 2 2 2 11 11 2 2
12 1 10 9 13 1 0 9 10 2 11 2 2
22 2 10 9 1 13 0 9 0 2 2 1 10 9 12 9 1 9 7 12 1 9 2
33 10 9 1 10 9 7 10 9 0 13 3 1 13 10 9 0 1 10 0 9 1 10 9 9 7 13 10 0 9 1 9 0 2
2 0 2
31 10 9 13 10 9 1 9 2 15 15 13 1 13 10 9 2 15 13 10 9 1 9 1 10 9 0 1 10 9 0 2
47 7 15 4 13 1 10 10 9 1 10 9 2 12 9 1 12 13 1 9 2 2 10 9 0 1 10 9 1 10 9 1 16 2 1 10 9 12 2 11 4 13 10 9 1 10 9 2
7 1 9 13 3 1 3 2
15 15 13 10 9 7 10 9 1 9 2 2 13 10 9 2
9 3 1 11 10 9 4 3 13 2
43 13 10 9 1 10 9 9 2 10 9 3 1 10 9 13 9 2 7 3 10 9 15 13 1 10 11 2 10 9 1 10 9 7 10 9 0 1 10 9 1 10 9 2
10 7 3 1 10 9 15 13 3 9 2
13 1 0 9 10 9 1 10 9 7 10 9 0 2
22 2 3 12 9 0 1 9 1 10 9 13 12 9 2 3 12 9 7 12 9 2 2
42 7 13 3 3 0 13 16 15 13 15 13 0 1 13 2 2 13 11 11 11 2 10 9 15 13 10 9 1 9 1 10 9 0 13 1 10 9 1 10 11 11 2
22 3 3 4 3 13 12 9 1 9 1 10 9 1 10 9 1 11 2 10 9 0 2
23 3 12 9 1 9 1 10 9 3 0 2 13 1 9 2 9 0 7 13 1 9 13 2
29 3 15 13 9 1 10 0 9 9 1 2 11 2 2 3 3 10 3 0 9 1 9 3 13 3 10 12 9 2
15 1 11 10 9 0 1 10 9 1 9 13 1 12 9 2
5 15 13 10 9 2
31 2 15 2 10 9 15 13 1 10 11 1 10 11 2 2 13 11 11 11 2 10 9 13 1 13 10 9 1 10 9 2
27 2 13 12 9 16 13 1 10 11 1 10 9 1 13 3 10 9 0 15 15 13 1 13 1 9 2 2
33 10 0 9 1 10 9 13 1 10 3 12 9 1 10 11 13 1 10 9 1 10 9 2 15 15 13 10 9 0 15 15 13 2
34 1 15 15 13 15 4 13 10 0 9 2 10 9 7 10 9 1 11 2 1 11 2 7 3 13 13 15 1 10 9 0 1 11 2
32 13 16 3 10 9 13 9 2 15 13 1 13 1 11 2 11 7 11 2 3 15 13 16 10 9 0 13 3 2 0 2 2
13 7 10 9 1 10 9 0 13 10 9 3 0 2
11 7 3 1 11 15 13 15 15 15 13 2
52 9 1 9 1 10 9 0 1 10 9 1 10 11 13 10 0 2 11 11 2 2 3 15 15 13 1 13 1 9 2 13 0 9 13 1 10 9 1 11 7 3 13 15 9 1 10 9 0 1 9 0 2
23 13 15 10 0 9 1 10 3 12 12 9 13 1 11 7 3 9 0 1 10 9 0 2
19 10 9 0 2 3 1 13 13 10 9 1 10 9 1 10 9 1 11 2
23 16 12 9 3 10 9 1 9 4 13 3 1 12 12 9 2 3 3 13 10 12 12 2
9 11 4 3 13 10 9 1 11 2
11 10 0 9 10 10 12 9 4 15 0 2
9 10 9 15 4 13 11 1 9 2
45 10 9 1 10 9 0 2 10 9 1 9 0 2 10 9 1 10 9 3 1 10 9 0 0 1 10 9 7 10 9 1 10 9 1 10 9 0 1 13 10 9 1 10 9 2
42 3 10 9 1 2 11 2 4 13 10 9 1 10 9 1 10 10 9 2 11 11 2 3 13 10 9 1 13 1 10 0 16 3 12 9 13 2 0 1 11 2 2
8 3 13 1 15 1 13 9 2
20 2 1 10 9 10 9 1 11 13 1 10 9 0 2 2 13 10 9 0 2
50 3 16 10 9 1 9 0 1 11 11 2 15 1 10 9 1 10 11 1 10 9 0 1 11 2 4 13 1 13 10 9 0 1 13 10 9 9 1 11 2 1 10 9 1 10 9 1 10 9 2
33 7 2 16 10 9 1 10 9 13 0 2 15 4 13 2 9 1 10 9 11 2 2 1 10 9 1 10 9 3 13 1 11 2
21 1 10 9 0 10 9 1 9 7 2 3 3 2 9 0 15 16 1 0 9 2
14 10 9 1 10 9 0 1 10 9 1 9 1 9 2
9 7 1 10 9 15 13 10 9 2
18 1 12 9 1 10 0 9 2 10 9 1 10 9 13 1 10 9 2
11 11 1 9 1 10 9 1 10 9 0 2
55 11 2 1 10 9 1 10 15 2 1 11 1 11 7 1 11 1 10 11 7 1 10 9 0 2 10 0 9 1 11 11 13 3 1 15 1 11 11 7 11 11 11 2 10 9 1 10 9 0 13 2 11 11 2 2
15 1 10 9 1 10 9 1 11 15 3 13 1 10 9 2
14 10 9 13 10 9 3 16 10 12 9 13 10 9 2
38 10 9 1 12 9 3 15 13 10 9 1 10 9 9 11 1 13 10 9 1 10 11 7 10 9 0 15 2 3 2 3 13 1 10 9 1 11 2
11 1 10 9 2 15 13 1 12 1 12 2
25 11 11 4 4 3 13 1 9 1 10 9 0 1 11 7 13 2 0 2 1 13 10 0 9 2
72 1 9 2 11 13 1 10 9 1 10 9 10 3 3 2 3 1 11 2 1 10 9 1 10 15 4 4 13 10 0 9 0 2 1 11 2 1 11 2 1 11 2 1 11 3 2 3 1 11 11 2 9 1 10 9 1 11 2 4 4 13 9 1 9 1 13 10 0 9 1 11 2
17 7 3 1 10 11 3 10 9 0 11 4 13 3 13 1 11 2
7 2 10 9 0 4 13 2
25 3 15 13 10 9 1 13 1 10 0 9 12 7 10 0 9 1 10 9 1 10 9 1 11 2
44 11 11 2 9 0 1 10 11 0 0 2 13 2 3 2 10 9 1 4 13 2 3 2 1 10 9 0 0 2 1 15 7 1 15 0 1 15 1 9 1 9 1 11 2
14 2 10 9 0 13 10 11 2 2 13 1 13 11 2
29 3 2 1 10 9 0 7 0 10 9 1 9 0 13 11 1 10 12 9 1 11 7 1 10 12 9 1 11 2
35 13 3 2 0 2 1 10 9 2 15 1 9 13 10 9 0 1 10 9 0 2 2 13 10 9 2 1 3 11 13 9 1 9 0 2
34 1 11 10 9 1 9 2 13 1 10 9 1 15 10 12 5 1 10 9 13 1 10 9 1 13 1 10 10 9 2 13 10 9 2
10 2 11 2 13 15 1 11 7 11 2
6 10 9 4 13 15 2
8 15 4 13 2 13 15 2 2
19 3 1 10 9 13 1 10 9 1 10 11 1 10 11 4 13 12 9 2
24 7 3 1 10 9 0 11 11 15 4 3 13 1 10 9 1 2 9 2 1 10 9 0 2
14 0 2 11 11 15 4 13 3 1 10 9 0 0 2
7 2 10 9 11 4 13 2
17 4 13 10 9 1 13 10 9 13 1 10 11 2 2 4 13 2
29 10 11 3 13 10 9 0 2 3 1 4 13 1 9 2 1 2 9 2 2 10 9 1 10 11 1 10 12 2
21 7 10 0 9 1 11 13 3 10 15 1 0 1 10 9 13 3 1 10 9 2
31 10 9 2 11 11 2 10 2 9 2 1 12 9 2 15 13 1 10 10 9 10 9 1 10 9 0 2 4 13 2 2
13 15 3 13 16 10 9 1 3 13 10 10 9 2
5 13 7 13 0 2
12 10 11 3 15 4 3 13 1 10 10 9 2
14 3 4 13 15 10 9 1 15 13 10 9 0 2 2
18 2 10 9 1 10 9 0 1 10 11 13 10 9 1 10 9 0 2
6 11 4 13 15 2 2
15 10 9 0 0 13 10 9 1 9 0 1 10 0 9 2
7 2 11 9 2 13 2 2
11 10 9 13 10 9 1 10 9 1 11 2
17 1 10 0 9 11 2 7 16 10 9 0 13 1 13 11 11 2
22 3 13 10 9 0 1 10 9 0 2 7 10 9 3 0 13 1 10 9 0 0 2
42 10 9 13 10 9 2 3 3 10 9 4 13 1 10 9 2 13 10 9 1 10 9 1 9 1 10 9 7 10 9 9 4 3 13 1 10 9 1 10 0 9 2
44 10 9 11 13 16 4 4 13 10 9 1 9 3 1 11 2 1 10 9 1 9 0 11 2 1 10 9 1 10 11 11 2 1 15 1 10 11 11 7 1 10 11 11 2
40 10 0 9 1 10 9 1 9 1 10 9 0 1 10 11 2 3 1 10 9 1 15 15 4 13 1 9 10 9 1 10 9 1 10 11 0 1 10 11 2
9 3 11 13 1 13 15 1 11 2
18 0 9 1 10 3 12 9 0 0 1 10 9 15 13 13 2 13 2
10 13 10 9 1 10 9 1 10 9 2
13 2 3 1 3 10 9 1 9 4 13 3 0 2
14 10 9 1 10 11 1 11 7 11 4 13 9 0 2
28 7 3 15 4 13 10 9 1 10 9 1 10 11 2 3 15 13 15 1 10 9 3 0 1 10 9 0 2
15 15 13 3 3 0 2 2 13 10 0 9 1 10 9 2
51 3 1 13 10 9 4 13 10 9 1 10 2 11 11 11 2 2 1 15 10 9 13 10 9 1 10 0 7 0 11 2 1 9 1 10 9 1 10 0 9 0 7 1 10 9 1 10 12 0 2 2
39 10 9 1 10 9 1 13 1 13 1 10 9 1 10 9 1 10 9 0 1 11 2 3 4 13 10 12 9 2 7 13 10 9 1 13 10 9 0 2
14 10 9 0 4 1 10 9 13 10 9 1 10 9 2
24 3 10 9 1 10 9 7 10 9 1 10 9 1 10 9 0 4 13 10 13 1 10 9 2
13 7 1 10 9 13 10 2 9 1 10 9 2 2
8 9 1 10 2 11 11 2 2
9 11 9 0 1 10 2 9 2 2
17 1 10 2 9 2 0 10 9 1 9 13 0 1 9 1 9 2
16 11 2 10 9 0 3 13 10 9 1 10 2 9 2 0 2
38 1 10 0 9 3 11 13 10 2 9 1 9 2 7 10 9 15 13 13 1 9 2 0 2 2 0 1 13 10 10 9 1 10 2 0 9 2 2
28 15 15 13 1 10 9 13 1 10 9 0 2 11 11 2 1 10 9 1 10 9 1 9 1 10 9 0 2
38 10 9 4 13 16 10 9 0 10 9 3 4 13 10 9 0 1 13 10 9 0 15 12 9 2 13 1 10 9 1 10 9 1 11 2 4 13 2
48 16 4 13 12 0 9 2 1 3 13 1 9 1 10 9 2 1 12 9 2 10 2 9 2 1 11 15 4 13 10 0 9 3 1 15 2 1 10 9 2 1 11 2 11 7 11 11 2
40 16 1 11 1 9 15 13 3 9 2 13 10 9 2 15 13 15 15 3 3 13 1 9 3 2 2 3 13 16 10 9 13 0 1 0 9 1 9 2 2
35 10 9 0 2 15 13 2 3 13 3 3 1 10 9 7 13 2 13 13 2 7 13 15 1 10 9 13 10 2 9 1 10 9 2 2
14 10 9 1 10 9 3 13 7 15 13 3 15 13 2
6 2 15 13 2 2 2
43 15 13 3 15 2 13 10 9 13 9 13 1 11 11 2 13 1 10 9 1 13 15 1 2 13 15 10 9 2 7 15 13 1 10 9 2 3 3 2 2 1 11 2
30 13 3 2 3 3 1 10 11 2 15 13 10 9 13 15 1 9 0 2 3 13 9 1 9 1 9 1 10 9 2
34 13 1 10 9 1 10 9 1 11 11 2 10 9 1 10 9 11 11 13 16 9 2 1 10 9 0 2 15 4 13 15 10 9 2
28 1 9 10 9 1 10 9 15 4 13 1 9 13 15 1 13 10 9 2 1 9 13 1 13 1 10 9 2
10 3 13 10 15 2 15 13 10 9 2
9 2 13 1 9 1 9 2 13 2
21 1 1 15 2 3 2 10 15 4 13 10 9 2 0 2 3 3 3 0 2 2
21 1 9 2 13 10 9 2 15 13 3 15 13 3 13 10 0 9 1 10 9 2
10 2 13 1 10 9 1 10 11 2 2
21 7 1 0 2 13 2 10 9 4 13 10 2 9 0 1 10 9 1 13 2 2
2 9 2
23 10 2 9 2 13 3 1 10 0 9 1 10 2 11 2 1 10 9 0 1 10 11 2
8 2 10 9 15 3 15 13 2
32 10 9 2 3 15 0 2 13 11 11 2 12 9 2 9 0 2 2 13 10 9 7 15 1 15 15 13 0 3 13 0 2
14 13 10 9 0 15 1 10 10 9 3 15 13 2 2
7 2 3 10 9 13 0 2
16 10 9 3 15 13 10 9 1 9 7 13 1 10 9 2 2
15 3 11 2 12 9 10 0 9 13 3 1 10 9 0 2
10 2 13 15 0 2 13 3 1 9 2
18 7 1 10 9 10 9 13 3 0 16 3 15 13 1 10 9 2 2
25 3 2 16 13 2 15 13 1 9 7 1 9 2 13 3 10 0 9 1 10 9 1 10 11 2
12 10 0 9 1 9 1 10 0 9 1 9 2
8 9 7 0 9 1 10 9 2
5 9 1 10 9 2
8 9 0 2 9 1 10 9 2
15 9 1 9 15 1 10 9 2 10 15 13 10 9 13 2
17 11 2 0 0 9 1 9 1 10 9 7 1 10 9 1 11 2
22 12 0 9 13 2 10 15 15 4 13 10 9 1 10 9 7 12 9 1 10 9 2
12 13 10 0 9 1 10 9 13 3 10 9 2
14 7 3 9 0 1 9 15 4 13 3 10 12 9 2
14 1 10 9 10 9 15 4 13 10 9 1 10 9 2
27 15 1 10 12 9 13 1 10 9 1 11 11 13 10 0 9 1 10 9 7 1 10 11 9 1 11 2
6 11 11 2 12 9 2
10 4 1 3 13 1 10 11 1 11 2
30 10 10 9 2 3 1 15 1 10 9 11 11 2 12 2 1 11 2 4 4 13 3 2 1 9 7 9 1 9 2
9 10 12 4 13 13 1 10 9 2
27 3 10 9 7 3 3 10 9 1 13 1 13 3 1 10 9 0 10 9 1 10 9 1 10 12 9 2
24 15 13 15 13 16 15 4 13 1 10 9 1 11 1 13 10 9 0 13 1 10 9 13 2
13 3 1 10 9 1 11 10 9 9 1 10 9 2
25 11 11 2 12 9 2 1 11 2 4 4 13 1 10 9 1 10 9 1 12 9 16 4 13 2
8 10 9 15 4 13 10 9 2
17 4 4 13 1 10 11 11 1 11 2 7 10 10 9 13 0 2
30 1 10 9 1 10 11 1 11 7 1 10 9 0 4 13 2 3 2 11 11 2 12 9 1 11 11 2 11 2 2
42 9 0 3 1 12 9 2 1 10 12 7 10 12 9 2 13 1 9 9 1 10 9 1 10 11 11 2 1 0 9 2 3 16 10 10 9 13 9 1 10 9 2
25 9 1 10 9 2 1 10 9 7 10 9 1 3 9 1 9 0 0 2 12 1 3 10 9 2
42 10 9 3 0 4 13 1 11 11 11 2 11 2 3 4 13 10 9 12 9 1 15 10 9 7 10 9 1 12 9 16 10 0 9 1 12 13 1 9 1 9 2
19 9 2 10 9 1 9 13 1 10 11 5 11 2 10 9 1 10 11 2
21 1 11 11 7 11 2 1 10 11 2 10 0 9 1 9 4 13 10 12 9 2
38 10 0 9 13 1 12 9 1 9 2 3 1 10 11 2 1 11 7 11 7 15 1 10 9 1 10 11 5 11 7 10 11 5 11 1 10 11 2
32 9 2 4 13 3 1 12 9 1 13 15 1 11 11 11 2 9 11 2 1 9 1 10 2 9 2 1 9 1 10 11 2
5 9 3 1 11 2
19 10 9 1 12 12 9 7 12 12 9 1 13 4 13 0 7 3 0 2
8 1 10 11 2 1 11 11 2
8 9 1 10 9 13 12 9 2
13 4 13 1 3 1 12 9 13 15 1 10 9 2
5 9 13 10 9 2
51 11 2 12 9 4 13 3 9 1 10 11 2 1 11 11 2 1 10 9 1 10 11 2 13 1 10 9 15 15 4 13 13 1 3 12 9 3 1 13 15 1 10 9 1 10 9 1 10 9 11 2
34 10 9 13 11 11 11 2 1 11 11 2 11 2 2 11 11 2 1 11 11 2 11 2 2 7 11 11 2 1 11 2 11 2 2
31 10 9 15 4 13 1 10 0 9 3 1 10 11 7 4 13 10 9 2 3 1 10 9 1 11 11 2 1 11 11 2
7 15 3 13 1 0 9 2
5 9 3 1 11 2
10 10 9 1 12 9 4 4 3 13 2
5 13 0 1 11 2
10 10 12 9 1 10 11 13 0 9 2
9 10 9 15 4 13 1 10 9 2
10 10 9 1 9 1 9 4 13 0 2
32 16 10 9 15 4 13 10 9 3 2 16 13 3 1 9 7 3 13 1 15 2 3 15 4 13 13 3 3 1 10 9 2
34 10 9 4 4 13 3 3 1 10 9 1 10 9 1 10 9 7 4 4 13 1 10 11 2 10 9 1 9 0 1 10 11 11 2
24 7 4 4 3 13 10 9 1 11 11 11 2 10 0 9 15 13 0 1 10 9 1 9 2
23 10 9 1 10 12 9 4 4 13 7 13 3 1 10 9 1 11 11 2 1 11 11 2
28 3 1 3 4 4 13 1 10 9 0 1 11 11 3 4 13 10 0 7 0 9 1 9 1 10 12 9 2
12 3 1 0 9 4 13 0 13 10 0 9 2
24 13 7 13 1 9 3 10 12 9 13 1 9 9 1 10 0 9 1 10 11 2 1 11 2
7 4 2 3 2 13 9 2
14 9 0 13 1 9 1 10 9 1 10 10 9 0 2
12 11 2 2 15 10 9 3 15 4 13 2 2
38 3 4 4 13 10 0 9 1 10 9 1 10 15 9 9 10 9 0 11 11 2 1 10 9 11 11 2 4 13 1 4 13 1 9 1 10 9 2
22 4 13 1 10 9 1 10 9 2 11 11 2 2 1 9 11 2 1 10 9 11 2
19 11 2 13 1 10 9 7 1 10 9 2 15 13 13 1 10 9 11 2
15 1 10 9 1 10 9 10 9 13 3 9 1 11 11 2
32 10 9 1 10 9 1 15 4 13 11 4 13 10 9 1 10 12 3 1 13 1 10 9 2 10 0 9 2 10 9 0 2
28 7 1 10 0 9 2 11 11 4 13 10 9 7 13 1 10 9 1 10 9 2 13 15 3 1 10 9 2
20 10 9 1 10 9 1 10 9 1 10 11 1 11 2 10 9 1 10 9 2
7 13 1 10 9 7 13 2
13 10 9 1 10 9 1 10 9 2 13 12 9 2
14 11 2 13 1 10 9 1 10 9 7 13 1 9 2
21 10 9 1 11 11 2 12 9 2 4 13 1 10 9 10 9 1 10 10 11 2
33 12 9 2 3 0 2 13 1 9 15 4 3 13 1 10 9 1 10 9 2 1 10 9 1 10 9 3 1 10 9 1 11 2
11 7 1 10 9 15 4 13 1 1 15 2
26 10 9 4 4 13 1 12 9 7 15 4 13 1 9 0 2 1 10 9 1 10 9 1 10 9 2
8 9 2 9 1 9 2 9 2
29 10 9 4 13 9 1 9 7 1 10 9 4 13 10 9 1 10 9 1 10 11 1 10 11 15 4 4 13 2
9 7 4 13 15 1 10 12 9 2
40 10 9 1 11 7 1 10 10 9 2 11 11 2 12 9 2 9 1 9 1 9 2 4 13 3 3 1 3 1 12 9 1 10 9 1 10 9 1 11 2
8 10 10 9 13 1 9 9 2
16 11 13 1 10 9 7 10 9 1 12 9 3 1 10 11 2
13 9 7 9 13 9 1 10 9 3 10 9 13 2
8 10 9 3 3 13 10 9 2
23 12 9 3 4 13 11 2 9 1 9 1 10 9 2 13 1 9 1 10 9 1 11 2
15 10 9 13 1 10 0 9 2 13 3 1 10 9 11 2
14 10 12 13 10 0 9 1 10 9 1 10 10 9 2
20 10 9 2 10 9 1 10 9 2 10 9 1 9 15 13 3 1 10 9 2
14 3 11 7 11 15 13 3 9 9 2 1 10 12 2
8 13 15 3 2 1 10 9 2
13 3 13 10 9 2 16 10 9 3 13 10 9 2
30 10 9 3 13 1 13 13 10 11 11 1 11 2 1 10 9 1 10 9 2 1 10 9 1 10 9 1 10 11 2
14 10 9 13 10 9 1 10 9 15 3 13 1 9 2
19 7 2 1 10 9 2 1 10 0 9 15 3 4 13 15 10 0 9 2
17 15 13 10 9 0 1 9 1 11 2 10 9 2 10 9 9 2
11 10 12 9 13 1 13 3 1 10 9 2
13 16 13 2 15 13 10 9 1 10 9 1 9 2
16 15 13 1 9 1 10 9 3 15 13 10 9 1 10 9 2
16 13 10 9 1 10 9 7 15 13 1 10 0 9 1 9 2
20 3 1 10 12 10 9 1 9 1 10 0 9 1 11 13 13 10 9 13 2
8 13 11 2 15 13 1 9 2
8 15 4 13 13 1 10 0 2
15 15 15 4 13 3 2 7 10 15 4 13 3 10 9 2
9 15 4 13 7 4 13 3 11 2
21 4 13 1 13 12 9 2 3 4 13 13 10 9 7 15 4 13 13 3 2 2
16 10 9 15 13 13 10 9 7 13 1 10 9 1 10 9 2
15 10 9 1 10 9 1 9 1 9 1 9 4 3 13 2
12 10 9 1 11 3 13 3 1 9 1 9 2
11 1 9 15 13 3 10 9 2 15 13 2
13 2 6 2 11 3 9 4 13 1 10 10 9 2
11 7 13 2 13 9 1 10 10 9 2 2
13 10 9 4 13 1 10 9 2 1 9 1 9 2
12 3 1 10 9 1 11 4 13 13 10 9 2
25 10 9 15 13 10 9 2 10 9 11 11 11 2 13 13 10 9 15 13 1 11 7 1 11 2
14 7 13 10 9 1 13 10 9 1 9 13 1 9 2
10 16 11 4 3 13 10 9 3 0 2
19 2 1 15 2 13 10 9 2 1 10 9 2 10 12 13 0 7 0 2
7 3 13 1 10 11 2 2
10 1 10 11 0 3 3 15 13 9 2
8 1 10 12 10 9 1 9 2
8 11 13 1 10 9 1 9 2
9 3 13 0 2 3 3 13 15 2
5 7 13 3 0 2
9 2 15 4 13 2 13 13 2 2
8 15 4 13 13 1 10 9 2
18 3 15 4 13 1 10 9 7 15 4 13 13 2 3 1 9 2 2
21 10 9 13 16 15 13 2 3 15 13 1 10 9 11 3 10 9 13 10 9 2
6 10 9 3 15 13 2
17 1 9 10 9 13 1 9 12 9 15 13 10 9 1 10 11 2
6 7 15 13 3 3 2
8 10 9 13 3 1 12 9 2
17 15 13 0 1 10 11 1 10 11 1 9 7 1 9 1 9 2
9 10 12 4 13 1 10 12 9 2
15 15 4 4 13 2 7 1 10 9 10 9 3 13 9 2
7 1 4 13 1 10 9 2
11 3 10 9 1 10 9 4 3 4 13 2
14 10 9 1 10 9 1 11 2 13 1 10 12 9 2
13 12 1 15 13 10 9 15 4 13 7 13 11 2
6 1 10 11 1 11 2
8 11 13 13 12 9 1 11 2
14 10 9 0 4 13 1 10 9 2 11 11 11 2 2
8 11 2 9 1 10 0 9 2
26 4 13 1 11 10 12 9 1 10 0 9 1 10 11 11 1 11 11 7 1 10 11 1 10 11 2
34 10 9 1 9 1 10 9 0 1 10 9 13 1 10 10 0 9 2 11 2 1 10 9 11 11 1 10 3 0 2 11 2 0 2
10 10 0 9 15 4 13 1 10 9 2
14 1 10 9 2 3 2 10 9 15 13 1 10 9 2
9 3 11 4 4 13 1 10 9 2
29 10 9 13 10 9 1 10 9 9 11 12 13 1 10 9 2 11 11 11 2 1 11 11 2 9 1 11 11 2
9 10 9 2 3 2 13 3 0 2
17 10 9 2 3 2 4 4 4 13 3 1 10 9 1 10 9 2
18 3 3 2 1 10 9 0 1 10 9 2 15 15 4 13 1 3 2
24 15 1 10 11 2 10 0 9 3 0 2 15 4 13 1 9 13 1 11 2 11 7 11 2
11 3 10 9 1 10 9 0 2 0 9 2
20 12 9 11 12 13 1 11 7 13 1 10 9 2 11 11 11 2 0 9 2
124 12 9 11 12 13 1 11 13 12 9 11 12 13 1 11 11 12 13 1 11 13 12 9 11 12 13 1 11 11 12 13 1 11 13 12 9 11 12 13 1 11 11 12 13 1 11 11 12 13 1 11 11 11 2 11 2 11 12 13 1 11 11 12 13 1 11 11 12 13 1 11 11 12 13 1 11 2 11 2 11 12 13 1 11 11 12 13 1 11 11 12 13 1 11 11 11 12 13 1 11 11 12 13 1 11 2 11 2 11 12 13 1 11 11 11 12 13 1 11 11 12 13 1 11
23 4 13 10 9 1 10 9 11 1 13 10 9 1 10 9 1 10 9 1 10 0 9 2
9 9 1 10 9 2 13 3 9 2
2 11 2
7 2 9 0 1 13 2 2
2 11 2
8 2 15 13 3 10 9 2 2
12 11 2 10 9 13 3 10 9 1 10 9 2
24 13 1 10 9 1 10 2 9 2 1 10 9 1 10 9 1 15 3 4 9 0 7 0 2
57 1 10 9 1 10 11 1 10 9 1 10 11 11 11 11 2 15 4 13 10 9 1 10 9 1 10 9 13 1 10 9 1 13 2 13 10 9 1 10 9 2 12 1 10 9 2 1 2 13 13 10 10 9 1 9 2 2
41 10 9 2 1 10 9 4 13 2 4 13 11 2 13 13 10 0 9 1 10 9 2 0 1 15 1 10 9 1 10 11 11 15 15 4 13 1 10 9 2 2
2 3 2
32 1 10 9 4 13 10 9 1 10 9 1 9 2 13 1 10 11 2 1 13 10 9 1 10 9 1 10 0 9 1 9 2
62 10 9 1 10 0 9 1 9 4 13 15 10 9 2 9 15 1 10 15 13 1 10 9 1 9 0 1 10 9 0 2 3 3 16 13 3 0 13 0 7 3 2 1 13 9 15 4 13 10 9 1 10 9 1 10 9 1 13 1 13 2 2
27 1 10 9 0 1 2 13 10 9 1 10 0 9 15 13 10 9 1 10 9 7 1 10 10 9 2 2
11 1 3 3 1 12 9 1 15 10 9 2
39 10 9 15 4 13 15 1 2 13 0 9 1 9 2 1 10 9 15 2 3 13 15 1 0 2 1 10 9 0 2 1 10 9 0 1 10 9 2 2
14 2 13 1 9 1 10 9 7 10 9 13 15 2 2
39 11 2 2 16 10 9 1 10 11 15 4 13 1 13 10 9 2 1 10 9 1 10 10 9 1 10 11 2 4 13 16 10 9 1 10 9 13 0 2
7 3 1 15 15 4 13 2
11 13 16 10 0 9 0 13 10 9 2 2
21 11 11 2 0 9 1 10 11 2 10 9 1 10 9 1 10 9 15 13 3 2
13 3 13 10 9 1 11 2 3 13 10 0 9 2
7 9 2 13 3 3 0 2
12 2 6 2 13 0 2 10 9 15 4 13 2
17 16 4 13 10 9 1 10 11 15 13 1 13 3 1 12 9 2
14 11 4 3 13 10 9 1 10 9 1 10 9 0 2
3 10 9 2
5 2 13 1 9 2
12 15 15 15 13 13 10 9 1 13 10 9 2
10 13 13 15 13 1 10 9 1 9 2
39 1 9 10 9 2 10 9 13 1 9 10 10 9 1 13 1 10 9 2 4 2 13 2 2 13 10 0 9 2 7 15 15 13 1 9 1 10 9 2
23 1 13 10 0 9 1 9 2 1 9 2 13 9 2 9 7 9 1 13 2 9 2 2
8 3 2 10 9 0 0 2 2
36 2 15 3 13 1 15 15 13 10 9 0 1 10 10 9 2 7 2 1 15 13 10 9 1 10 9 2 3 15 13 9 0 3 0 2 2
6 13 1 10 11 11 2
27 2 4 13 10 9 1 13 2 3 1 15 13 10 9 15 2 16 13 3 2 13 3 0 7 0 2 2
17 10 9 1 9 4 13 10 0 9 1 10 9 1 10 9 0 2
13 10 9 13 16 10 9 13 3 0 1 10 9 2
21 3 13 16 15 13 1 9 15 2 3 1 13 15 2 13 10 9 0 3 0 2
11 3 2 13 10 9 1 13 0 2 0 2
20 13 0 16 13 1 13 10 3 0 1 10 9 10 9 2 13 10 9 2 2
7 10 9 3 4 13 15 2
5 2 1 10 9 2
14 13 0 13 10 0 9 0 1 10 9 13 9 2 2
10 15 13 1 10 9 2 0 2 2 2
8 2 6 2 1 10 9 0 2
8 1 11 3 13 1 3 2 2
12 3 13 10 9 15 13 1 13 3 10 9 2
44 2 3 1 16 10 9 3 13 16 13 1 10 9 3 4 13 13 10 9 7 16 13 15 13 3 13 10 9 1 2 1 9 2 13 15 1 10 0 9 1 10 9 2 2
23 11 2 10 9 1 10 9 7 1 10 10 9 2 10 9 2 0 2 1 10 9 0 2
33 11 11 2 0 9 11 1 10 11 7 0 9 1 10 11 11 2 3 13 15 1 0 1 10 9 1 10 9 1 10 11 11 2
19 2 13 10 9 1 13 10 9 1 10 9 1 10 9 0 2 2 13 2
20 16 10 9 13 9 2 4 3 13 10 2 9 2 1 10 9 1 10 11 2
5 2 13 1 3 2
10 3 1 10 9 10 9 15 4 13 2
19 4 13 3 10 9 13 1 10 9 2 10 9 15 13 3 1 10 12 2
16 10 9 1 15 3 15 13 10 9 1 9 1 11 7 9 2
13 3 2 1 10 9 13 3 2 10 9 4 13 2
18 3 3 1 10 9 1 2 9 2 1 10 9 1 10 9 1 9 2
25 3 15 13 13 0 13 1 9 0 3 1 10 2 9 2 1 10 9 1 10 9 1 9 2 2
17 1 9 13 10 9 15 4 13 7 13 1 9 10 11 11 2 2
11 2 3 2 3 16 1 15 13 3 0 2
14 10 11 11 13 10 9 0 2 15 4 13 3 13 2
21 15 1 10 9 4 13 10 9 3 1 10 1 3 1 10 9 1 10 9 0 2
15 13 9 15 13 1 9 1 9 2 0 2 9 0 2 2
10 3 15 13 2 1 10 9 1 11 2
13 13 10 9 1 9 2 4 13 1 10 9 0 2
9 3 16 10 9 3 13 3 0 2
37 16 1 11 2 3 1 10 9 3 0 2 15 4 13 10 9 1 10 9 2 15 13 3 9 1 9 0 2 3 0 1 10 9 1 3 15 2
24 15 13 3 10 9 0 1 11 2 3 10 9 0 4 13 1 10 9 1 13 10 9 2 2
3 0 9 2
16 10 9 9 1 2 11 2 1 10 9 1 2 11 11 2 2
8 2 11 3 0 7 0 2 2
3 0 11 2
14 2 3 15 13 10 10 4 13 3 2 3 0 2 2
20 13 10 10 9 1 10 0 9 1 10 9 7 1 10 0 9 1 10 9 2
7 13 10 9 1 9 0 2
27 7 13 10 10 9 1 10 9 2 10 15 15 3 10 11 11 7 10 11 4 13 1 10 9 0 2 2
11 11 11 3 13 9 15 13 10 0 9 2
15 7 13 3 13 9 1 13 3 10 10 9 1 11 11 2
13 3 2 1 9 1 13 2 3 13 3 11 11 2
23 3 10 10 2 0 9 2 13 15 0 2 3 16 1 13 2 0 2 15 13 3 0 2
28 11 4 3 13 10 2 0 9 2 2 15 4 13 3 3 2 13 1 9 2 0 1 15 2 0 2 2 2
12 3 2 1 3 13 10 2 9 2 13 0 2
6 13 1 10 0 9 2
17 2 13 16 11 13 10 9 1 13 15 1 13 1 10 9 2 2
45 7 11 13 1 2 9 0 2 7 3 0 0 2 2 1 10 2 9 3 3 0 15 1 10 9 13 10 9 1 10 0 9 1 10 9 7 1 10 0 9 1 10 9 2 2
5 7 13 1 9 2
34 1 13 10 9 1 10 0 9 1 11 2 15 13 10 10 9 0 1 10 12 2 1 10 12 2 2 2 1 10 9 11 7 9 2
30 9 2 3 2 13 3 13 1 11 2 15 13 1 13 1 10 9 0 1 10 9 1 11 11 1 2 3 9 2 2
12 3 2 11 2 10 9 13 2 3 9 2 2
25 2 3 1 11 0 10 9 1 11 15 13 3 0 1 9 2 1 9 2 7 3 1 9 0 2
19 13 0 1 10 9 1 9 15 15 13 1 3 7 15 15 13 9 9 2
25 1 13 15 2 11 4 13 10 10 9 7 3 13 3 1 10 9 7 9 0 1 10 11 11 2
42 3 16 3 4 13 1 10 0 12 9 1 10 9 2 13 1 10 9 1 10 9 9 2 3 13 16 2 1 11 2 11 13 10 9 1 3 3 3 1 11 2 2
2 9 2
12 13 10 9 15 13 1 15 13 1 10 9 2
33 2 3 1 11 0 2 11 3 13 10 9 1 9 0 2 3 13 1 10 9 0 1 10 9 2 1 10 9 2 1 10 9 2
7 7 13 9 13 3 15 2
9 13 10 9 15 13 1 10 9 2
39 7 11 3 4 3 13 0 9 0 1 10 11 7 1 10 11 2 10 10 9 13 3 0 1 10 10 9 2 2 10 10 9 4 13 1 9 3 0 2
44 3 2 13 16 10 0 9 0 2 7 1 15 0 2 1 10 9 1 11 11 13 10 9 1 11 11 2 1 15 15 13 10 0 9 1 15 0 2 10 0 9 1 9 2
20 7 13 0 10 10 4 13 3 2 3 0 2 2 10 10 9 1 13 15 2
19 3 16 3 2 1 9 2 10 9 9 15 13 3 0 1 15 2 2 2
22 3 15 4 13 1 13 15 1 10 9 15 1 3 4 13 1 13 1 9 15 0 2
17 2 3 2 15 13 10 9 1 9 15 13 1 13 10 0 9 2
24 15 1 0 1 10 9 16 11 13 10 9 1 15 0 2 13 15 0 10 9 15 13 3 2
9 3 2 10 9 13 10 9 0 2
11 3 13 2 1 10 9 2 10 9 0 2
33 15 13 3 10 9 1 10 9 0 0 2 10 9 15 13 3 0 7 15 13 3 1 15 1 9 10 3 0 2 3 0 2 2
9 7 1 11 0 2 10 9 13 2
26 2 11 1 9 2 3 1 10 13 10 0 9 2 13 3 0 2 10 9 1 10 9 0 7 0 2
27 1 11 0 15 13 3 10 9 1 10 9 9 2 1 10 9 1 9 1 10 10 9 4 13 10 9 2
36 7 1 11 11 2 15 4 13 3 10 0 9 2 3 1 10 0 9 11 4 13 15 0 1 10 9 1 9 1 10 9 0 1 0 9 2
18 13 3 16 10 10 9 4 13 3 1 10 9 1 10 9 7 3 2
43 0 9 13 10 10 9 3 0 2 3 13 1 9 1 9 2 1 13 1 10 9 7 1 10 9 2 7 10 0 9 1 15 10 9 1 9 4 3 13 13 10 9 2
6 13 10 9 1 11 2
40 1 10 9 1 10 0 9 15 13 2 13 2 10 9 0 1 11 2 13 10 10 9 3 0 7 9 15 13 2 3 3 1 11 2 10 11 4 13 2 2
14 11 13 10 9 1 10 0 9 0 1 10 10 9 2
18 2 7 10 9 1 9 3 13 10 9 2 13 3 10 9 0 2 2
17 3 2 11 13 1 13 16 3 16 10 9 11 13 10 0 9 2
17 2 11 13 10 9 15 15 4 13 2 13 10 0 10 9 2 2
28 16 15 13 3 1 10 9 16 10 3 1 10 9 13 3 15 15 15 13 3 2 15 13 1 10 9 0 2
12 7 10 9 1 11 13 0 1 10 9 0 2
8 1 9 2 15 4 13 9 2
3 13 11 2
35 13 0 3 16 3 15 15 13 3 1 10 9 0 0 15 4 13 1 10 9 0 2 0 2 0 2 3 0 2 1 10 9 0 2 2
19 13 10 9 1 13 2 10 9 1 9 1 13 9 1 10 9 1 11 2
10 13 2 9 2 10 9 9 1 11 2
53 2 4 3 13 10 15 2 13 2 13 2 13 15 15 4 13 1 10 9 2 1 10 9 2 1 10 9 2 1 10 9 2 1 10 9 2 1 10 9 2 13 9 7 13 10 9 2 9 2 9 2 9 2
50 13 10 9 15 13 1 10 9 1 11 1 13 9 2 3 13 3 1 10 10 9 10 9 13 1 10 9 2 15 13 3 10 9 0 15 13 3 15 10 9 13 1 10 9 2 1 0 9 0 2
40 10 15 13 10 9 0 7 3 0 7 0 2 10 0 9 13 3 0 2 7 13 1 13 3 10 10 9 3 16 13 1 13 10 10 9 2 10 10 9 2
20 11 3 15 13 1 9 3 1 9 2 13 15 0 3 16 15 13 3 2 2
5 13 10 9 0 2
29 2 13 16 11 4 13 15 1 10 15 2 1 11 2 10 9 11 7 10 11 2 1 13 1 3 13 1 11 2
15 10 9 1 13 3 10 10 2 9 2 7 10 10 9 2
28 10 9 1 10 2 9 2 2 15 13 10 0 9 1 10 0 9 2 13 3 1 13 15 1 9 3 0 2
15 10 9 2 2 0 2 2 13 1 10 10 9 1 11 2
14 2 3 2 1 10 9 1 15 3 2 3 1 3 2
29 13 16 11 13 1 13 15 2 7 16 13 1 10 10 9 13 15 10 9 1 10 11 13 3 1 3 13 15 2
46 3 13 3 0 1 11 11 2 7 0 1 9 7 1 9 2 3 16 10 0 11 4 13 2 1 10 9 1 9 4 13 10 2 0 2 9 0 1 10 9 0 0 7 0 2 2
13 1 13 10 9 1 10 11 9 2 0 1 11 2
29 2 1 10 11 11 4 13 10 10 10 9 1 9 0 0 1 13 15 15 15 13 2 10 0 9 1 10 9 2
25 10 9 3 13 3 10 15 2 7 13 16 13 1 11 16 11 15 13 2 9 15 3 3 13 2
35 13 16 13 0 3 16 0 2 3 16 10 0 9 0 0 4 13 11 7 10 0 11 4 13 1 9 7 1 0 9 3 1 11 2 2
22 7 1 9 1 11 2 13 1 10 9 0 2 1 10 2 9 2 1 10 11 9 2
8 7 1 10 2 0 9 2 2
18 2 11 13 10 9 1 13 15 2 3 13 2 1 13 1 10 9 2
45 13 16 4 3 13 10 10 9 1 9 0 2 13 10 10 9 1 10 9 2 10 15 15 3 10 11 11 7 10 11 13 1 10 9 0 3 16 3 1 10 9 0 0 0 2
27 7 13 15 2 11 2 15 13 2 1 10 10 0 13 15 2 10 9 0 1 9 15 13 1 4 13 2
38 7 1 9 2 3 1 10 0 9 13 1 10 2 9 9 2 1 11 11 2 13 3 10 9 2 1 10 10 0 9 7 9 2 1 10 10 9 2
17 13 3 0 16 10 9 1 11 4 3 13 1 10 10 9 0 2
12 10 10 9 3 4 13 0 1 10 0 9 2
37 15 4 3 13 1 11 10 9 15 15 0 3 4 3 13 2 3 13 16 10 10 9 13 3 10 9 1 10 9 0 1 10 2 9 2 0 2
19 10 9 3 3 13 3 15 2 10 9 0 1 13 1 13 2 1 13 2
24 11 13 10 9 1 10 9 7 10 9 0 1 13 10 9 0 7 3 3 0 9 0 2 2
7 15 1 9 2 1 9 2
16 13 2 1 11 2 10 9 1 10 9 1 10 2 13 2 2
6 2 13 10 9 11 2
33 3 1 13 15 1 13 1 10 9 1 10 9 1 9 2 11 2 9 7 9 2 15 4 13 9 1 9 1 9 7 9 0 2
5 3 16 2 2 2
3 3 16 2
27 2 3 16 3 10 9 13 1 9 0 2 3 0 7 0 1 15 2 3 2 7 3 3 0 7 0 2
26 1 12 9 2 15 13 2 1 9 3 4 3 13 1 10 9 3 0 1 10 0 9 0 1 9 2
22 13 15 2 13 10 9 15 13 1 11 2 1 11 1 10 11 1 11 11 1 11 2
18 3 2 13 1 10 11 9 10 3 10 15 15 13 1 10 10 9 2
16 9 3 7 3 3 2 3 2 1 10 9 1 9 0 2 2
69 13 15 2 11 13 0 3 1 13 10 9 1 11 2 1 13 10 10 9 1 10 13 10 9 1 10 9 0 0 1 10 9 9 3 16 2 13 11 2 2 1 10 13 10 9 2 3 10 9 9 4 13 10 0 9 1 9 0 1 9 2 9 9 2 7 1 9 2 2
9 3 2 3 1 9 2 10 9 2
10 2 3 1 10 9 1 11 2 2 2
9 7 10 9 2 3 2 3 13 2
41 2 1 10 9 9 11 4 13 1 9 7 1 15 15 13 2 1 9 1 10 3 13 10 9 3 0 1 10 9 1 9 1 10 9 1 10 0 9 11 11 2
36 1 9 4 13 1 13 15 13 1 10 0 9 0 2 4 13 16 15 4 13 15 0 1 15 15 3 13 7 1 10 9 15 3 13 2 2
78 7 1 10 9 15 13 3 1 13 1 9 2 1 10 2 0 9 0 15 15 13 7 15 13 2 1 15 2 7 3 1 15 2 1 10 10 10 9 7 1 10 10 9 15 6 7 1 9 13 3 3 0 1 10 15 15 2 1 13 10 10 9 7 1 13 3 1 13 2 3 1 15 0 8 1 11 2 2
10 12 9 3 0 1 9 1 10 9 2
5 9 2 0 9 2
12 12 9 3 0 2 15 1 11 7 1 11 2
21 3 2 1 10 9 1 10 9 7 1 10 9 2 12 7 12 9 1 10 9 2
15 10 9 1 10 9 0 7 1 10 2 0 9 2 0 2
16 10 9 1 9 2 11 11 2 13 1 13 2 12 9 0 2
8 10 9 7 10 11 1 11 2
20 3 13 1 9 2 13 9 0 2 15 13 1 11 1 10 9 0 1 11 2
20 10 9 13 9 0 2 10 9 1 11 2 10 9 1 11 2 11 2 11 2
8 11 13 1 11 1 10 12 2
37 0 13 10 0 9 1 11 12 2 16 10 10 0 9 2 15 13 10 9 2 1 10 12 2 13 10 0 9 7 4 13 1 10 11 1 11 2
40 1 10 12 2 11 11 7 3 2 1 9 2 11 1 9 2 12 2 2 11 2 12 2 2 10 11 4 13 2 12 2 15 13 10 11 1 9 1 11 2
27 1 10 12 2 11 0 7 3 11 11 1 10 12 2 9 1 15 10 11 1 11 15 13 10 9 0 2
34 1 10 12 2 13 9 2 11 11 7 11 11 1 11 11 2 7 1 10 12 9 1 9 1 10 9 0 1 11 2 10 11 11 2
2 11 2
6 1 13 10 9 11 2
9 2 15 13 10 9 1 9 2 2
42 11 11 11 3 4 13 9 2 3 1 10 9 1 11 11 3 9 9 10 9 13 3 3 0 1 10 9 1 9 13 3 1 10 9 2 3 0 1 10 9 0 2
55 10 11 2 9 1 10 9 0 3 0 2 4 13 13 13 15 2 11 11 11 7 2 3 2 11 2 10 9 0 1 2 11 1 9 2 10 9 15 10 9 4 13 10 0 9 11 2 10 0 1 10 9 0 11 2
26 4 13 10 9 11 11 1 13 9 1 10 9 1 10 11 11 2 13 12 9 3 1 10 10 9 2
60 7 1 10 11 10 9 1 10 11 0 1 11 2 11 11 2 2 1 10 9 15 4 13 15 7 13 10 9 11 10 11 2 15 3 16 4 13 1 10 9 1 10 9 1 11 11 11 15 4 13 1 4 15 13 1 9 3 3 0 2
68 1 13 10 9 7 1 13 10 10 9 1 11 11 15 13 3 11 11 2 11 11 7 3 10 9 2 11 11 11 2 15 1 10 9 1 11 4 13 1 10 10 9 1 2 11 13 11 2 2 10 11 1 10 9 1 10 9 1 9 15 4 13 3 1 10 9 11 2
26 1 13 9 7 9 1 10 10 9 11 11 11 13 3 10 10 9 2 13 10 3 1 10 10 11 2
32 2 13 10 9 15 4 13 1 11 2 2 4 13 2 13 3 10 9 16 10 9 1 10 9 13 3 1 9 1 10 9 2
2 9 2
22 1 11 10 9 1 10 0 9 0 2 0 7 0 2 15 13 10 9 1 10 9 2
14 10 9 1 13 10 9 1 9 9 3 1 10 9 2
27 13 1 10 9 1 11 7 1 10 9 0 2 13 3 1 9 1 10 9 13 1 10 10 9 1 13 2
19 11 10 11 1 11 15 13 0 1 10 9 15 13 1 9 1 11 11 2
22 10 9 0 2 13 3 1 10 9 0 2 4 3 13 3 1 10 9 1 10 11 2
34 13 15 1 10 9 15 13 1 10 9 2 3 3 15 13 9 1 9 13 1 10 9 1 10 9 2 15 13 3 10 9 1 9 2
26 15 15 13 3 1 9 0 2 0 2 13 0 3 1 10 0 9 15 13 1 10 9 15 15 13 2
43 1 10 9 0 7 1 10 9 4 13 10 9 1 11 11 11 2 12 2 12 2 2 13 1 10 9 1 10 11 1 11 7 13 3 16 13 10 9 1 10 0 9 2
45 10 9 13 10 9 1 10 11 1 10 11 7 1 10 12 2 9 3 1 10 0 9 1 11 11 2 15 4 13 9 1 10 9 3 1 10 9 0 1 10 9 1 10 9 2
34 10 15 2 1 15 1 10 11 1 11 11 2 13 10 9 3 0 3 16 13 9 7 9 2 10 9 0 13 1 9 7 9 0 2
23 1 9 1 10 9 2 10 9 2 10 9 1 10 9 0 15 13 1 9 10 9 0 2
41 1 10 12 9 7 1 10 12 9 1 9 15 13 10 9 0 1 10 11 1 10 11 3 4 4 13 10 9 13 1 9 0 7 13 1 9 3 1 10 9 2
46 10 9 3 13 1 15 0 16 15 4 13 10 9 1 9 1 10 9 1 10 9 13 3 3 0 1 4 13 1 10 2 9 1 10 9 0 2 10 0 12 9 1 10 10 9 2
37 9 0 7 0 1 10 10 9 0 2 1 10 9 15 3 13 10 10 9 1 9 1 10 9 1 10 9 2 1 9 0 1 11 7 1 11 2
50 3 11 1 10 9 0 1 11 1 10 0 9 12 3 15 13 10 0 9 7 1 10 9 15 15 13 1 11 12 9 3 2 13 10 9 1 10 9 1 10 9 7 1 10 0 9 1 10 9 2
29 10 15 13 10 9 0 1 10 9 1 10 11 2 1 10 9 15 13 3 1 15 2 1 2 3 2 10 9 2
48 10 9 15 11 13 3 3 2 7 1 10 15 13 9 2 1 3 13 2 1 9 7 1 10 15 15 13 3 16 4 13 11 1 10 11 2 10 11 2 10 11 2 10 11 2 3 11 2
61 16 15 13 15 15 13 13 10 9 1 10 10 9 2 0 1 9 2 7 3 1 9 0 15 15 13 3 1 9 7 15 13 1 10 9 1 0 9 1 9 1 10 9 0 1 10 10 9 1 13 2 1 10 10 9 7 1 10 10 9 2
30 10 9 3 13 1 10 9 1 11 11 1 11 2 1 10 15 13 13 10 9 1 13 10 9 15 13 0 7 0 2
54 10 9 2 8 8 10 10 9 1 10 9 0 2 10 9 2 10 9 1 10 9 2 10 9 1 13 10 9 1 9 2 1 9 3 13 3 1 0 2 13 1 15 10 9 0 2 10 9 1 11 8 8 8 2
48 7 1 11 7 3 1 11 7 1 11 11 13 10 9 1 10 10 0 9 7 10 9 2 0 2 15 13 1 10 9 1 11 2 3 3 13 10 9 1 11 7 10 9 0 1 11 11 2
49 10 9 13 3 1 11 11 2 1 11 11 2 11 11 7 11 11 1 9 1 11 1 10 11 7 1 10 11 1 10 11 0 7 0 13 10 9 3 0 15 3 15 4 13 1 10 9 0 2
42 1 10 9 15 13 10 9 2 11 10 11 2 10 9 13 3 10 9 1 9 0 7 0 2 13 1 10 9 11 2 11 7 11 7 1 9 1 10 10 9 11 2
8 15 9 1 10 0 9 0 2
45 7 1 9 2 1 13 1 10 9 1 10 10 9 2 10 9 13 9 0 1 10 9 0 1 15 15 13 9 1 10 9 1 10 0 11 11 2 1 15 13 0 13 10 15 2
14 10 10 9 13 0 2 0 1 10 9 7 3 0 2
28 1 13 10 9 1 10 9 2 3 3 0 2 13 16 13 10 9 3 0 1 10 10 9 7 10 3 0 2
22 3 3 0 10 9 1 15 10 9 15 13 1 9 2 3 3 0 2 1 10 9 2
19 1 10 0 9 2 3 12 5 12 9 2 13 10 9 11 1 11 0 2
52 15 13 10 9 1 9 1 10 9 1 10 9 0 1 10 9 2 1 10 9 10 13 0 2 0 2 0 1 10 9 1 10 9 1 10 9 2 3 10 9 0 1 10 11 15 15 13 1 13 10 9 2
10 1 10 9 10 9 1 10 9 0 2
26 9 13 1 10 9 15 13 1 10 9 2 1 10 9 0 15 3 13 1 11 1 11 1 10 9 2
22 1 10 0 9 10 9 7 10 9 15 4 13 0 7 10 9 1 9 13 10 9 2
44 10 9 1 10 0 9 15 13 16 11 13 10 9 0 2 1 10 9 0 15 13 13 9 3 0 1 9 15 4 3 1 10 9 4 13 1 10 9 0 1 10 9 0 2
49 13 10 9 3 13 1 10 10 9 2 10 10 9 0 13 10 10 9 2 10 10 9 15 13 1 9 7 1 9 2 10 9 1 10 9 13 13 1 10 9 13 1 3 10 9 1 11 11 2
31 7 3 1 10 0 9 15 13 1 10 10 9 3 1 10 11 1 11 15 13 10 9 7 10 9 1 9 7 9 0 2
26 10 0 9 15 13 1 9 1 9 1 10 9 2 11 11 11 11 2 3 13 1 10 11 10 11 2
27 10 9 1 9 15 13 2 9 15 13 2 9 2 9 2 9 2 10 9 0 15 15 13 1 10 9 2
11 13 0 1 10 10 9 1 10 0 11 2
15 10 9 0 7 0 13 11 2 3 0 2 7 3 0 2
3 9 0 2
9 10 0 9 4 13 1 10 9 2
20 11 11 4 13 1 0 9 10 9 0 0 1 9 2 9 2 9 1 9 2
55 16 3 13 2 10 0 2 9 2 1 10 9 1 9 2 15 10 9 9 1 10 0 9 15 13 1 9 0 1 10 2 9 1 10 9 2 2 13 4 15 13 1 9 1 13 10 10 9 0 7 0 1 10 9 2
25 3 13 2 1 10 9 2 9 0 2 9 1 9 0 2 9 0 13 1 0 2 9 2 0 2
12 7 10 9 13 1 0 9 10 9 1 9 2
29 10 9 11 11 2 15 4 13 1 9 1 9 10 9 0 2 13 10 9 1 10 0 9 1 10 2 9 2 2
35 1 15 13 10 9 1 11 2 10 9 1 9 11 2 10 9 0 1 10 9 11 7 1 10 10 9 3 13 2 1 10 9 0 2 2
22 16 3 15 13 1 13 1 10 9 1 10 9 0 7 0 10 9 3 0 1 11 2
8 10 9 1 10 9 4 13 2
50 11 2 15 1 10 9 4 13 10 9 3 1 10 9 1 10 9 2 4 13 3 10 10 1 10 9 1 9 2 11 9 2 9 12 2 9 12 2 1 10 9 0 1 10 9 2 1 10 9 2
56 9 1 10 0 9 2 13 1 3 4 3 13 2 1 9 2 13 10 9 1 10 15 7 15 1 10 9 13 3 1 1 13 10 0 9 1 10 3 0 9 0 2 2 11 13 16 13 10 0 9 1 10 9 1 9 2
21 2 10 9 15 13 1 10 9 1 10 9 2 2 13 15 1 10 10 9 0 2
15 1 10 9 2 10 9 2 10 0 9 13 10 0 9 2
42 10 10 0 9 2 10 9 2 11 11 2 9 1 10 11 0 2 9 1 11 11 2 4 13 1 10 9 2 1 9 2 13 15 1 10 9 1 10 9 0 2 2
3 10 9 2
15 11 2 1 10 9 1 11 11 2 4 13 1 13 15 2
3 10 9 2
27 3 1 10 9 11 2 1 9 3 3 0 2 4 13 9 1 2 9 2 0 10 12 9 1 10 9 2
27 11 2 1 10 0 9 2 4 13 1 13 9 0 1 13 1 10 9 1 10 3 0 2 9 0 2 2
8 7 10 0 9 4 3 13 2
23 11 11 2 10 9 1 11 11 2 13 2 3 1 4 1 10 9 13 2 9 3 0 2
22 1 11 2 15 1 10 9 13 1 10 9 3 0 1 15 2 13 1 10 13 3 2
15 2 11 2 15 13 1 9 2 1 10 10 9 2 3 2
10 13 3 2 1 10 10 9 2 2 2
15 13 3 1 10 9 1 10 9 2 13 2 1 0 9 2
16 3 4 13 2 3 1 15 2 10 0 12 9 1 11 11 2
32 1 10 9 1 10 0 9 2 15 4 13 9 3 1 10 9 1 11 2 13 15 15 11 13 2 10 9 1 10 9 2 2
13 13 15 10 9 13 13 10 0 9 1 10 9 2
2 11 2
8 9 7 9 1 10 9 0 2
12 10 2 11 2 15 11 4 13 2 11 2 2
17 10 9 1 10 9 1 10 9 13 3 9 1 9 1 10 9 2
28 15 13 9 15 3 13 1 13 10 9 2 3 3 13 1 10 10 9 2 16 3 3 4 13 16 13 15 2
36 15 13 3 1 10 9 1 10 9 2 7 13 3 16 10 0 9 1 10 9 13 10 9 2 7 3 13 9 1 10 9 7 1 10 9 2
5 15 7 10 15 2
6 3 0 7 3 0 2
6 10 0 9 13 0 2
28 7 3 10 9 1 9 13 10 9 15 13 10 9 0 2 9 1 10 10 0 9 1 10 9 1 10 9 2
14 3 13 9 2 3 16 10 9 13 0 7 3 0 2
46 7 15 13 0 2 1 13 10 9 13 1 10 9 1 10 12 2 3 13 1 10 0 9 1 11 2 1 11 2 1 11 2 1 11 2 1 11 2 1 11 2 1 11 11 2 2
14 10 9 13 3 10 9 1 9 2 10 9 1 9 2
68 1 9 2 15 13 3 13 1 10 9 15 13 1 13 15 1 13 10 9 1 9 0 1 10 9 0 7 10 10 9 2 1 10 9 1 9 1 15 10 9 15 13 1 10 9 7 10 2 9 2 2 1 13 10 9 1 10 9 0 2 15 1 10 9 13 7 13 2
16 10 9 0 15 4 13 0 1 13 10 9 0 1 10 9 2
48 12 9 3 2 1 10 9 1 10 12 2 2 11 11 13 1 11 10 0 9 1 10 11 1 9 1 11 11 2 15 1 10 9 0 1 10 9 0 2 7 3 3 0 2 1 10 12 2
42 10 9 1 10 0 9 4 13 3 1 10 12 9 1 10 9 1 10 9 1 10 2 11 2 2 10 9 1 15 11 13 1 13 10 13 1 10 9 1 10 9 2
40 7 15 4 13 12 9 1 9 2 13 10 9 3 0 2 3 1 0 2 1 10 9 0 1 10 0 11 2 2 0 2 0 2 1 10 9 3 0 2 2
11 10 9 13 1 12 9 7 13 12 9 2
6 15 4 13 12 9 2
12 11 13 0 1 10 9 7 3 13 10 9 2
15 15 13 2 3 2 1 13 13 12 9 1 9 7 9 2
21 3 1 10 0 9 2 2 11 2 2 13 0 10 9 1 10 9 1 10 9 2
19 6 3 13 2 1 10 9 1 9 1 10 9 2 13 1 3 1 3 2
16 2 13 2 10 9 0 7 10 9 2 13 1 10 9 2 2
6 13 1 10 10 9 2
25 11 1 9 13 1 9 1 9 15 1 10 9 3 13 2 3 13 2 3 0 1 10 10 9 2
18 1 10 9 7 1 10 9 15 13 0 13 15 3 1 10 0 9 2
3 15 13 2
27 10 9 1 10 11 2 10 9 1 10 11 2 10 9 7 10 9 1 10 11 2 10 9 1 10 11 2
73 7 3 1 0 2 1 10 0 9 1 9 13 1 10 9 0 2 4 4 3 9 13 1 10 9 0 10 12 0 9 1 10 9 2 15 3 3 4 13 15 2 2 15 15 3 13 2 15 15 3 13 2 2 1 10 0 9 1 10 9 2 16 13 2 16 13 10 11 1 10 11 2 2
40 16 2 1 10 9 1 10 0 9 0 2 11 11 2 12 2 12 2 2 11 4 3 13 1 10 9 0 1 11 1 9 2 13 1 10 0 2 0 9 2
2 11 2
33 3 4 13 10 9 15 3 15 13 1 13 9 1 9 0 7 0 2 7 3 3 9 13 7 13 1 10 9 7 1 10 9 2
38 10 15 15 13 0 1 10 2 0 9 2 2 10 9 13 1 11 11 2 1 10 11 15 13 10 0 9 1 10 9 1 10 12 7 10 12 9 2
6 3 10 9 13 15 2
39 16 11 4 13 1 10 10 0 9 2 16 10 10 0 9 1 9 15 4 13 11 7 3 11 1 9 2 10 9 2 10 9 3 0 4 13 10 15 2
27 10 9 1 10 9 2 10 9 1 10 9 2 10 9 7 10 9 1 10 9 2 10 9 1 10 9 2
17 10 9 15 13 3 10 2 3 2 2 3 4 13 10 0 9 2
11 7 3 1 10 9 15 4 13 9 2 2
9 10 15 3 15 13 1 10 9 2
14 15 13 1 10 1 3 1 10 9 0 1 10 9 2
28 10 11 13 10 10 0 9 3 12 9 3 2 10 12 9 12 2 16 1 11 4 13 1 11 10 9 11 2
53 10 9 11 11 2 1 10 9 0 2 13 10 0 9 7 13 16 2 10 9 0 1 11 4 13 10 9 0 15 13 13 1 10 0 9 1 10 9 0 2 1 10 9 0 15 15 13 1 9 1 9 2 2
31 1 15 2 3 0 1 9 2 13 16 10 0 9 0 1 11 1 9 4 4 13 1 10 9 1 10 9 1 10 9 2
12 7 3 13 10 9 1 10 9 1 10 9 2
12 2 11 2 1 11 1 10 9 15 15 13 2
26 11 2 3 11 11 11 4 13 10 9 11 11 1 10 9 0 1 11 2 1 10 9 1 10 9 2
29 11 11 2 11 11 2 11 11 2 0 9 1 9 0 2 11 11 2 11 11 7 11 11 2 13 1 11 11 2
36 2 7 10 9 13 1 15 15 15 4 13 2 3 1 15 15 4 13 13 2 2 13 1 11 11 11 2 3 11 11 15 13 1 12 9 2
25 7 1 9 1 10 9 2 10 9 4 13 10 2 3 2 9 1 9 1 11 7 9 1 9 2
21 10 9 1 10 9 1 2 11 2 2 1 10 15 4 4 13 3 10 9 11 2
7 10 9 1 10 9 0 2
51 2 7 13 3 16 15 13 16 10 11 2 3 11 2 13 10 11 0 2 2 13 11 11 2 9 7 9 1 9 0 1 9 2 15 1 10 9 13 10 9 1 9 7 10 9 1 11 1 10 12 2
2 11 11
2 9 2
6 9 1 10 9 0 2
6 11 2 11 13 11 2
12 0 9 1 10 11 3 1 10 9 1 9 2
6 10 9 1 10 9 2
31 11 2 0 9 1 11 11 9 1 10 9 0 1 2 11 2 2 1 10 15 10 2 11 2 13 1 9 0 3 2 2
20 0 3 10 9 1 10 0 11 11 2 15 1 9 9 15 4 13 10 9 2
9 1 10 9 15 13 10 9 0 2
11 13 10 9 0 1 10 9 0 1 11 2
40 3 3 1 10 9 3 15 13 16 10 9 0 11 11 2 13 15 1 10 9 0 2 4 4 13 1 10 9 1 10 9 11 2 16 1 10 9 4 13 2
19 10 9 1 9 13 1 0 9 7 4 4 13 1 10 9 1 9 13 2
13 10 9 1 9 2 3 12 9 1 9 7 9 2
26 10 11 4 13 10 9 15 1 10 9 15 13 13 1 10 10 9 0 7 0 7 10 10 9 0 2
21 9 3 1 11 11 2 11 11 2 7 11 11 2 10 9 2 2 13 1 9 2
14 10 11 11 13 1 11 4 13 10 0 9 1 9 2
19 2 11 2 4 13 10 12 9 2 10 0 9 4 13 10 12 9 2 2
30 1 9 9 15 13 1 10 11 11 1 11 2 15 15 4 13 3 1 10 11 0 2 10 9 2 10 12 9 2 2
5 11 11 4 13 2
9 3 13 0 16 13 10 9 0 2
11 13 10 9 0 2 1 10 0 9 2 2
6 9 1 9 11 11 2
31 1 10 9 0 11 11 2 10 9 11 11 7 11 11 13 10 2 9 2 16 1 11 2 11 13 10 2 9 0 2 2
38 1 10 9 1 9 15 4 13 3 10 9 0 13 9 1 10 9 1 11 1 10 9 1 11 13 1 10 9 10 9 3 1 10 2 11 11 2 2
39 3 11 2 16 4 15 13 10 2 11 11 2 1 10 0 9 2 13 16 11 11 13 10 9 7 16 11 2 1 11 7 10 0 11 11 13 10 9 2
8 9 1 9 1 10 9 0 2
30 9 1 9 13 1 9 2 1 11 11 2 13 10 9 10 9 1 9 1 9 15 13 9 0 1 10 9 1 9 2
49 13 10 9 9 2 7 3 2 10 9 1 10 9 2 1 10 9 1 0 9 13 2 8 8 8 8 2 7 13 1 10 9 11 11 1 10 11 11 2 10 9 1 10 9 3 0 1 11 2
2 9 2
24 1 11 2 1 10 9 15 13 13 10 10 9 1 10 9 2 10 9 13 10 10 0 9 2
10 10 10 9 1 10 9 0 1 11 2
3 11 11 2
14 2 15 15 13 2 1 12 9 4 3 13 15 2 2
19 2 1 12 9 1 10 9 2 11 3 13 10 9 7 13 1 9 2 2
6 2 10 9 1 11 2
5 13 15 1 0 2
6 3 4 13 15 2 2
14 2 10 9 15 13 13 1 10 9 1 12 9 2 2
23 11 2 13 3 3 1 9 2 10 9 4 13 10 9 1 12 9 2 3 1 10 9 2
21 15 7 11 2 12 9 3 2 4 13 10 9 0 0 2 15 4 13 1 9 2
27 15 13 12 9 1 10 9 2 13 3 10 10 10 9 2 7 10 9 13 10 9 1 10 0 9 2 2
17 10 3 9 0 7 10 9 2 15 1 11 11 2 15 13 3 2
21 2 1 10 9 1 11 15 4 13 3 2 1 10 10 9 2 13 10 11 2 2
17 7 15 15 13 2 13 3 2 3 4 13 16 4 13 3 0 2
10 3 13 10 9 2 13 1 9 2 2
74 10 9 1 9 1 10 9 2 1 11 1 11 2 13 0 7 13 1 10 9 2 9 0 1 9 2 9 15 13 1 10 9 2 1 10 9 1 10 9 2 9 0 1 0 2 10 0 9 1 9 15 13 10 9 0 2 0 2 1 10 9 2 10 9 0 7 10 9 0 1 13 10 9 2
14 3 2 10 9 3 3 0 7 10 9 0 1 9 2
36 2 13 10 9 3 0 2 13 10 9 2 2 1 12 9 4 13 1 9 1 10 9 0 7 10 9 2 10 9 2 10 9 1 10 9 2
9 15 13 3 11 1 13 10 9 2
21 10 0 9 15 13 10 9 2 13 10 9 1 10 9 2 10 9 2 10 9 2
10 10 9 1 9 16 11 13 10 15 2
14 3 15 13 10 10 9 0 1 13 15 13 1 9 2
19 7 3 15 13 10 9 2 15 4 13 3 10 9 1 10 9 1 12 2
9 2 15 13 10 0 9 2 2 2
46 16 11 2 12 9 2 3 4 13 10 9 1 9 2 15 15 4 13 1 9 12 9 3 2 10 9 15 4 13 1 13 10 12 9 15 1 9 4 13 1 9 1 10 11 11 2
16 2 11 11 1 10 9 1 10 11 2 1 15 2 2 9 2
9 6 2 3 1 13 2 1 15 2
18 7 3 3 15 15 13 3 15 2 10 9 1 9 3 4 13 3 2
13 2 13 1 0 2 2 10 11 13 10 9 2 2
15 15 15 4 3 13 2 7 3 13 2 3 4 13 15 2
8 6 2 3 15 15 13 2 2
48 10 9 3 2 1 10 9 1 9 3 1 11 2 1 13 3 10 10 2 9 1 9 2 2 3 13 1 0 11 2 2 1 9 1 10 11 11 2 11 3 4 4 13 15 15 1 9 2
18 10 9 4 13 2 13 2 15 4 13 9 2 15 15 4 13 0 2
19 1 10 9 13 15 15 15 4 4 13 10 9 1 10 11 2 1 9 2
52 3 2 10 9 1 9 2 15 15 4 13 2 11 0 13 1 9 2 2 4 13 9 1 10 9 2 13 10 12 9 1 13 2 10 9 1 10 9 0 15 4 13 1 10 9 0 1 10 9 0 2 2
5 10 11 15 13 2
17 2 7 3 15 13 1 13 10 9 16 10 9 13 13 1 15 2
3 10 9 2
31 7 13 16 16 4 13 10 9 1 13 1 9 10 9 15 13 1 9 2 9 1 15 10 9 13 0 2 11 15 13 2
8 2 3 4 13 9 2 9 2
10 2 13 10 9 1 13 2 13 2 2
11 16 15 13 1 9 3 15 13 15 2 2
23 1 10 9 0 7 10 9 1 9 1 9 9 2 11 11 2 12 9 2 13 3 0 2
2 13 2
48 2 13 10 9 15 4 13 2 13 1 9 10 10 9 2 1 13 1 9 1 10 9 10 9 7 10 9 13 15 3 0 1 10 9 2 13 15 10 9 2 13 10 9 1 10 10 9 2
11 15 15 13 1 15 2 3 1 10 9 2
6 4 13 1 10 9 2
21 10 9 1 10 10 9 13 0 3 13 1 10 9 2 1 10 9 1 12 9 2
7 3 15 0 7 0 2 2
24 13 10 9 1 11 7 3 3 10 9 1 9 2 7 10 11 3 13 3 0 1 10 9 2
22 9 0 2 9 0 2 10 1 11 2 2 15 15 15 13 16 13 1 13 10 9 2
10 13 3 0 3 10 9 3 2 2 2
5 15 15 13 13 2
10 2 10 9 13 1 10 9 1 3 2
35 16 15 4 13 15 2 16 10 9 13 10 9 2 16 4 13 0 1 3 13 15 13 1 10 9 1 10 2 13 12 2 13 12 2 2
17 1 9 13 3 15 15 15 13 1 9 1 13 10 10 9 2 2
2 13 2
18 2 3 13 1 9 2 4 13 10 0 11 11 2 3 15 4 13 2
3 13 3 2
16 3 2 13 3 9 2 13 13 10 9 3 0 1 10 9 2
10 15 12 13 1 13 10 10 9 2 2
18 11 11 3 15 4 13 2 13 1 10 9 2 13 1 10 0 9 2
14 3 13 1 10 9 0 2 3 13 10 10 10 9 2
2 9 2
3 2 11 2
3 10 9 2
3 11 11 2
3 0 2 2
2 11 2
5 13 0 13 0 2
5 10 9 1 11 2
13 2 13 3 9 2 7 10 9 15 4 13 2 2
10 13 1 11 1 10 9 10 9 13 2
15 2 15 13 9 0 2 7 15 13 11 1 11 11 2 2
6 7 13 1 13 0 2
20 11 2 3 16 13 3 0 2 2 13 10 9 13 15 1 10 9 11 11 2
10 2 6 2 2 15 13 13 10 9 2
18 7 3 2 3 16 13 10 9 2 2 4 13 3 11 11 12 2 2
18 15 2 13 1 10 9 1 9 0 2 15 13 1 13 9 1 9 2
17 1 10 0 9 1 11 1 10 9 1 9 1 2 11 0 2 2
8 10 9 0 1 10 10 9 2
3 1 12 2
29 16 11 10 9 2 16 16 10 12 9 13 0 2 13 10 0 9 1 9 0 2 7 0 2 1 12 9 3 2
25 4 13 1 9 10 9 1 2 11 10 9 2 1 10 10 9 15 13 1 15 2 1 11 11 2
19 1 9 1 13 3 1 12 9 2 13 3 9 1 9 0 1 0 9 2
18 1 10 9 1 10 9 7 10 9 1 10 9 15 15 13 3 0 2
7 13 0 7 2 0 2 2
8 13 10 0 9 1 11 11 2
20 13 3 10 9 2 11 13 10 9 0 1 9 1 9 2 9 0 7 11 2
20 7 13 1 10 9 1 10 10 9 1 9 1 10 9 0 3 0 1 13 2
24 2 11 11 11 2 1 11 11 11 2 1 15 13 10 9 0 7 0 1 10 9 11 11 2
21 2 15 13 1 13 9 3 16 13 2 13 16 10 9 15 13 1 10 9 0 2
37 7 3 13 0 2 2 13 10 9 11 2 9 0 2 9 1 10 0 9 13 1 10 9 3 1 13 10 0 2 9 1 10 9 2 0 2 2
8 2 1 10 9 13 10 9 2
16 15 13 9 0 2 1 9 1 9 0 2 9 0 1 9 2
34 3 13 0 1 10 9 1 10 9 2 7 13 13 1 9 0 1 11 2 11 11 2 15 15 13 13 2 9 2 1 9 1 9 2
17 10 9 1 15 15 15 4 13 15 1 11 11 3 13 3 2 2
9 13 3 1 9 4 13 10 9 2
8 2 13 10 9 1 0 9 2
15 13 15 2 7 9 16 10 9 15 13 1 10 0 9 2
9 13 15 15 13 2 1 11 11 2
23 4 13 1 13 10 0 9 9 3 2 11 1 11 11 2 9 2 3 16 15 13 15 2
21 15 4 13 1 10 2 9 2 1 10 11 11 2 11 15 4 13 10 9 2 2
7 15 13 10 9 1 9 2
5 3 15 4 13 2
6 2 15 13 16 13 2
7 15 13 3 1 10 9 2
13 7 3 1 11 2 16 13 1 13 15 13 3 2
9 15 13 3 9 1 15 9 2 2
17 2 15 13 3 2 13 0 2 13 2 3 2 1 10 9 2 2
10 13 3 0 1 15 15 13 10 9 2
19 1 9 4 13 10 3 0 2 7 3 13 2 9 2 1 10 10 9 2
15 13 9 0 16 15 13 1 10 3 1 10 9 2 2 2
15 13 0 16 4 13 15 10 9 1 11 11 1 11 11 2
8 2 6 2 15 13 11 2 2
12 1 11 13 1 0 9 2 3 4 13 11 2
13 10 10 9 13 10 9 3 1 10 15 2 6 2
20 4 13 15 2 2 13 0 2 13 10 9 1 9 1 10 9 1 9 0 2
8 3 16 13 10 9 1 11 2
7 9 1 9 1 10 9 2
5 9 13 10 9 2
40 1 10 10 9 15 4 3 13 1 10 9 1 12 2 0 7 0 2 7 1 9 1 9 7 10 9 1 9 1 9 4 13 1 13 0 9 1 10 9 2
9 4 3 13 3 9 10 3 13 2
9 9 0 2 9 1 10 0 9 2
12 10 9 0 4 13 1 0 10 9 1 9 2
3 9 0 2
10 3 15 13 1 13 10 10 9 3 2
22 11 11 2 11 2 2 15 13 10 9 2 15 13 2 16 15 4 13 10 0 9 2
24 4 13 3 1 10 9 13 1 13 13 1 10 9 1 10 9 1 9 0 1 13 10 9 2
15 3 2 1 9 1 9 2 13 3 3 13 10 10 9 2
35 3 16 15 13 15 2 7 3 13 16 10 9 9 2 13 10 9 0 2 13 10 10 9 7 1 9 13 1 13 1 0 10 10 9 2
6 1 10 9 13 0 2
21 13 10 9 1 9 7 1 10 9 4 13 16 13 13 9 0 1 9 0 2 2
28 9 1 10 9 2 0 9 2 3 16 3 4 3 13 1 15 13 10 9 7 2 3 2 13 13 10 9 2
27 7 3 3 13 13 16 10 10 9 13 3 0 7 3 0 1 15 2 1 9 1 10 0 9 1 9 2
49 13 15 2 13 16 4 13 15 1 13 1 10 9 16 2 16 4 3 13 15 2 1 3 16 10 10 9 2 7 15 13 3 3 0 2 15 13 1 10 9 2 15 13 0 13 1 13 15 2
19 10 2 9 2 3 13 3 9 0 1 9 0 7 1 0 9 1 9 2
11 10 9 4 13 10 9 0 1 0 0 2
50 15 13 10 9 16 15 13 1 13 1 0 9 0 2 9 2 9 2 9 7 9 3 13 1 15 1 9 2 1 10 10 9 9 0 4 13 1 13 9 2 9 2 9 1 10 9 3 3 0 2
7 10 11 11 1 11 11 2
3 9 0 2
3 13 13 2
16 1 9 0 1 0 9 1 9 15 13 9 1 10 9 0 2
26 13 13 1 10 9 1 9 1 10 9 0 1 9 1 10 11 0 11 11 2 3 1 10 9 0 2
10 7 15 1 10 9 15 3 3 13 2
28 12 2 1 10 9 1 13 10 9 1 10 9 1 10 3 0 7 3 3 0 9 15 13 9 7 9 0 2
60 12 2 1 10 0 7 0 9 1 9 15 13 10 9 1 9 2 16 1 10 9 1 9 1 10 9 1 10 12 5 1 10 9 1 9 13 10 9 3 0 1 10 11 2 7 16 10 9 1 9 15 3 4 13 13 3 10 9 0 2
40 10 9 13 1 10 9 16 2 3 2 2 15 4 13 1 3 1 12 9 1 10 9 0 0 1 10 0 9 2 3 1 10 4 13 7 3 10 9 2 2
42 13 3 10 9 1 13 16 10 9 1 10 9 0 3 13 10 9 1 13 7 13 2 7 16 10 0 9 2 7 0 7 0 2 13 10 0 9 1 0 9 0 2
16 9 2 16 10 0 9 1 9 4 13 13 1 10 9 0 2
42 9 2 16 2 13 10 9 0 1 12 9 2 0 7 0 2 4 13 10 9 0 7 13 1 10 0 9 1 10 9 2 9 3 2 7 3 0 9 1 9 2 2
15 9 2 16 4 13 1 9 10 9 1 10 9 1 9 2
27 9 2 16 2 1 9 0 2 10 9 0 3 4 13 1 9 0 1 10 0 9 1 10 11 1 9 2
39 10 9 15 1 11 13 1 10 11 1 10 11 4 3 3 13 1 10 9 0 15 13 1 10 9 10 9 3 0 1 13 10 11 2 3 12 9 2 2
39 13 3 0 2 3 1 10 9 1 10 11 1 10 9 2 13 10 9 0 0 2 10 9 13 10 9 16 1 3 12 9 1 11 15 13 10 11 2 2
18 3 15 1 10 15 2 1 10 11 10 9 4 13 15 1 10 12 2
12 10 9 0 13 3 13 7 10 0 9 0 2
17 13 1 10 11 16 3 13 0 13 15 1 10 9 1 10 12 2
3 11 11 2
2 11 2
3 9 0 2
5 9 1 10 9 2
13 10 0 9 1 9 13 1 13 9 1 10 9 2
22 1 0 9 2 13 10 11 2 13 1 11 11 2 9 11 11 11 9 1 10 11 2
21 3 15 4 13 2 7 15 4 3 13 2 15 15 4 13 1 10 9 1 11 2
25 0 9 2 0 9 2 0 9 2 7 4 13 12 9 1 3 16 1 10 9 2 3 9 12 2
20 1 10 10 9 1 9 10 9 15 4 13 10 9 1 10 0 7 10 0 2
3 11 11 2
9 10 9 1 11 9 1 10 11 2
9 1 10 9 0 15 13 10 9 2
35 3 13 9 13 15 1 9 7 13 15 1 10 0 9 15 2 1 9 2 9 7 9 2 3 13 15 1 13 1 15 3 13 1 11 2
31 15 13 11 0 1 11 1 10 10 11 1 11 7 15 2 9 0 13 1 10 9 0 2 15 13 0 7 0 16 13 2
12 1 10 9 13 1 0 7 10 9 3 0 2
20 13 10 10 9 3 13 1 9 7 9 1 9 2 1 9 7 9 1 9 2
15 13 10 9 7 10 9 3 13 1 9 7 1 9 0 2
11 13 10 9 10 9 0 15 15 13 11 2
16 12 9 1 9 13 1 9 0 2 3 1 10 9 3 0 2
20 15 1 16 13 1 10 9 1 10 9 9 0 2 0 1 9 7 1 9 2
18 10 9 15 15 13 3 1 10 11 15 15 3 3 13 1 9 0 2
5 11 11 2 11 2
3 9 9 2
6 9 1 10 9 0 2
67 10 9 9 1 10 2 9 0 2 1 10 9 2 1 15 1 9 9 10 9 4 13 10 2 9 2 2 3 1 9 12 9 7 12 12 9 2 1 10 9 1 9 7 1 10 9 1 9 2 13 1 9 10 9 0 1 10 2 9 9 2 2 13 10 10 9 2
47 1 10 9 16 15 4 13 1 9 10 0 9 1 10 2 9 2 1 10 0 9 0 2 13 0 1 10 9 13 15 3 10 9 1 10 0 9 2 1 10 15 10 9 4 13 3 2
21 3 2 3 1 3 4 13 10 9 0 2 10 9 13 1 13 3 1 12 9 2
2 0 2
95 16 13 1 9 10 9 0 1 10 9 1 9 2 13 16 10 9 13 3 2 1 10 9 1 13 9 3 3 0 1 9 1 9 7 9 2 3 3 1 10 9 7 10 15 2 7 1 15 1 10 11 7 15 1 10 11 2 13 13 10 9 1 10 2 9 2 1 11 2 1 11 7 1 11 2 2 2 3 13 3 13 13 10 10 9 1 10 9 2 3 1 10 10 9 2
62 7 1 9 2 10 0 2 9 2 3 13 1 13 2 7 3 1 2 13 2 1 10 9 0 10 9 3 0 2 3 16 3 13 10 0 2 0 2 9 1 10 9 1 10 9 2 1 9 1 15 15 10 0 9 0 13 2 0 7 0 2 2
2 11 2
64 3 13 16 3 15 13 0 9 1 10 2 9 9 2 2 10 9 3 15 3 10 9 11 15 13 1 13 3 9 2 16 4 13 1 0 9 2 2 10 9 2 10 9 13 16 10 9 1 9 7 9 13 3 10 9 1 10 9 1 10 10 9 0 2
57 3 13 15 1 10 9 2 7 13 10 9 1 13 10 9 0 13 1 10 9 1 10 9 7 1 10 9 2 1 3 13 1 10 9 2 3 0 1 13 10 9 13 2 15 13 10 0 9 3 1 10 9 1 10 9 2 2
9 15 13 3 1 13 10 9 0 2
34 10 2 9 9 2 3 4 2 7 4 2 13 15 1 10 9 3 10 9 15 4 13 1 13 15 1 10 9 1 10 9 7 9 2
20 13 10 9 1 13 2 16 15 13 16 2 3 9 2 13 2 0 9 2 2
3 10 9 2
8 3 15 13 1 10 0 9 2
8 16 13 11 11 2 15 13 2
8 2 3 15 13 1 9 0 2
43 1 10 10 9 2 3 1 10 15 2 13 1 10 9 2 3 1 10 9 1 9 2 4 13 1 9 10 9 0 7 0 1 9 7 15 13 9 16 15 3 4 13 2
40 10 9 1 10 9 15 15 13 1 9 1 13 1 0 9 13 10 9 0 2 1 15 13 9 1 13 2 7 2 15 13 2 3 4 13 3 1 10 9 2
23 3 2 13 15 0 1 10 0 9 1 10 9 0 2 4 13 10 9 1 10 10 9 2
30 2 10 0 9 13 16 2 1 10 9 0 2 15 4 13 1 10 0 9 2 15 3 10 9 4 13 10 10 9 2
26 3 16 1 3 1 9 15 15 15 13 3 3 7 3 1 10 10 9 2 0 1 10 1 13 15 2
10 2 13 2 13 7 13 10 9 2 2
12 3 3 0 1 10 9 0 15 13 15 0 2
32 3 13 3 0 13 13 15 2 3 16 1 10 9 2 6 2 10 9 13 1 13 2 10 9 0 15 13 1 10 10 9 2
32 7 13 10 0 9 15 10 9 13 2 1 9 16 15 13 1 10 9 2 1 10 9 2 1 0 9 2 1 10 9 0 2
46 13 3 0 16 10 9 1 10 9 15 13 1 13 1 10 9 1 10 9 10 9 1 10 0 9 2 3 13 1 10 9 1 10 9 2 7 1 10 0 9 10 0 9 1 9 2
18 2 4 13 16 13 1 10 10 9 2 7 16 13 0 10 10 9 2
15 13 2 3 2 16 10 9 1 9 1 10 9 13 0 2
38 15 13 10 9 0 2 10 15 13 1 13 16 10 11 1 10 11 15 13 10 10 9 2 1 13 13 13 10 15 15 15 13 4 13 1 10 9 2
22 7 3 13 16 3 13 2 1 9 1 10 9 2 10 0 9 7 9 1 10 9 2
58 16 15 15 13 1 10 9 1 10 9 7 1 10 9 2 3 15 13 9 16 10 10 9 3 13 2 16 10 10 9 4 13 2 3 2 1 9 2 10 11 1 10 11 13 10 9 2 1 9 2 15 1 13 15 16 13 9 2
12 3 13 10 9 2 7 13 16 3 4 13 2
21 2 1 10 9 0 9 7 9 4 13 10 10 9 3 1 15 1 10 9 11 2
5 3 15 13 0 2
31 10 9 1 11 13 15 1 10 0 9 1 9 2 7 10 10 0 9 13 1 10 13 2 16 3 15 4 13 2 0 2
14 7 3 15 9 2 3 0 3 0 2 15 13 13 2
59 3 10 10 9 2 0 11 2 13 1 10 9 10 9 0 2 15 13 10 9 1 10 9 3 0 2 1 10 15 10 9 0 13 1 10 10 10 9 2 7 1 9 13 1 13 3 1 10 9 1 10 9 15 15 13 1 1 15 2
13 13 16 15 13 1 13 10 3 10 10 0 9 2
17 10 9 13 10 9 1 10 9 15 3 13 1 11 1 10 11 2
7 11 11 2 9 1 9 2
16 2 11 3 13 3 10 9 1 11 2 3 13 10 9 2 2
21 1 10 0 9 11 2 3 1 9 1 10 11 13 10 9 0 1 10 9 0 2
34 11 13 1 13 10 9 1 10 9 13 2 3 3 1 4 15 13 2 10 9 1 10 12 9 2 2 3 15 15 13 3 2 2 2
20 2 13 3 3 0 1 12 9 3 2 13 10 9 2 2 13 10 9 0 2
3 10 9 2
14 15 13 15 2 10 11 2 10 11 7 10 11 2 2
32 9 1 9 0 1 9 1 13 1 9 10 9 0 7 0 2 13 1 10 15 1 13 1 0 9 10 9 1 10 9 0 2
20 7 3 1 10 9 2 10 11 4 4 13 9 1 10 0 2 9 2 0 2
3 11 11 2
60 3 1 13 10 9 3 13 10 9 15 2 3 2 13 9 1 10 0 9 2 13 9 1 0 9 2 2 15 13 3 3 1 10 0 9 2 15 13 0 2 4 13 1 10 0 1 10 15 1 13 15 15 13 2 15 13 1 13 2 2
34 3 1 13 1 9 13 11 11 2 9 0 2 0 9 0 1 11 11 1 10 9 0 1 10 9 9 2 15 1 11 13 10 9 2
18 1 11 1 0 13 2 15 10 9 2 10 9 4 13 9 1 11 2
46 7 13 16 10 9 1 11 7 11 1 10 9 13 0 2 1 10 9 1 9 1 11 7 10 0 9 0 0 2 3 16 10 0 9 4 13 15 1 10 0 9 0 1 10 9 2
19 13 3 1 10 9 1 11 16 12 9 3 11 7 11 13 10 9 0 2
10 4 13 10 10 9 2 13 11 2 2
29 10 9 13 1 10 0 9 1 10 9 1 10 11 2 11 2 10 15 4 13 1 15 1 10 9 1 10 9 2
10 15 13 16 15 13 1 10 9 11 2
18 15 13 1 9 1 10 9 13 1 10 9 2 7 13 1 10 9 2
14 11 1 11 3 13 10 9 7 3 10 9 13 12 2
17 7 13 9 10 9 7 10 9 15 15 4 13 1 10 11 2 2
10 1 10 11 15 13 3 1 9 0 2
7 1 10 12 10 9 9 2
8 11 12 9 9 1 10 9 2
21 11 11 1 11 2 12 9 12 2 13 10 9 1 10 0 9 1 10 9 12 2
44 10 11 15 13 1 10 9 1 11 7 11 13 15 10 9 1 12 9 2 9 0 1 10 9 2 13 10 9 15 13 10 9 0 2 0 1 10 9 2 1 11 1 11 2
13 1 10 9 13 3 1 9 10 9 1 10 9 2
13 1 10 9 12 11 13 3 13 1 10 0 9 2
9 10 9 7 10 9 1 10 9 2
16 11 9 1 10 12 9 2 10 11 13 10 9 1 10 9 2
6 11 0 1 10 9 2
7 11 9 0 2 13 11 2
10 1 10 0 9 11 2 10 9 0 2
34 15 13 1 13 2 15 13 1 13 2 16 10 9 13 3 1 9 2 7 10 9 7 10 9 2 15 13 2 13 10 10 0 9 2
38 3 13 12 9 1 9 2 12 9 0 15 3 13 10 11 1 9 1 10 9 2 7 15 13 10 3 13 1 13 10 9 15 13 1 11 7 11 2
30 11 15 3 3 15 13 7 11 15 15 13 10 9 7 3 13 10 9 0 1 10 9 2 16 13 1 10 9 0 2
12 6 2 13 10 9 10 0 2 4 13 11 2
10 9 0 1 9 2 13 1 10 9 2
41 10 9 0 15 13 1 13 15 2 16 11 11 13 12 9 7 10 9 3 13 9 1 9 2 16 11 11 13 1 10 0 9 7 15 13 3 10 10 9 3 2
28 1 13 2 3 2 16 15 13 11 1 9 2 16 10 9 1 9 4 13 10 9 1 9 2 9 2 9 2
40 15 15 13 13 1 9 2 3 10 11 7 10 11 11 13 12 9 1 9 1 12 2 1 10 11 7 10 11 2 7 11 3 13 3 10 9 1 10 9 2
50 3 15 15 13 2 13 3 1 9 2 1 11 11 2 10 9 0 15 15 13 1 10 9 2 9 1 10 9 13 3 1 10 9 1 10 9 7 10 9 1 10 10 9 0 15 13 10 0 9 2
27 16 10 0 9 15 15 13 2 3 3 15 15 13 10 15 0 1 13 15 2 1 10 9 1 10 9 2
62 3 1 10 9 2 13 15 0 1 15 13 1 11 7 11 1 10 12 2 7 13 0 9 1 10 9 0 2 10 9 0 1 10 11 2 2 10 9 1 10 9 15 13 13 1 10 13 15 2 13 1 13 10 9 1 10 9 1 10 10 9 2
17 7 3 11 2 13 10 10 12 9 1 10 9 2 13 10 9 2
9 1 9 15 15 15 13 1 9 2
15 1 9 2 9 2 9 15 13 13 7 15 13 10 9 2
10 10 9 0 3 3 0 1 10 11 2
13 11 2 10 9 1 9 1 10 9 1 10 11 2
27 10 9 15 13 10 0 11 3 4 13 10 9 1 10 0 9 1 10 11 0 4 4 13 1 10 9 2
7 10 9 0 1 11 11 2
49 10 9 0 0 2 15 13 10 9 1 10 9 1 9 1 13 10 9 1 10 9 1 9 1 11 7 13 15 3 1 9 1 10 9 2 4 13 3 10 0 9 1 10 9 0 1 10 11 2
11 7 3 4 13 10 9 3 1 10 11 2
42 11 11 15 4 2 13 2 1 13 1 12 10 0 11 2 1 12 10 0 11 7 1 12 10 0 11 2 15 13 10 0 9 1 9 7 1 10 9 1 3 12 2
41 1 10 11 2 3 1 10 0 9 1 9 2 1 11 7 3 1 11 2 10 0 9 2 0 9 0 2 4 13 1 13 10 9 1 3 3 1 10 10 9 2
18 10 9 1 9 15 4 13 1 13 15 15 0 2 1 13 10 9 2
46 3 3 10 9 4 13 1 13 1 10 11 2 3 13 10 9 1 9 2 11 15 4 13 1 9 1 10 9 1 13 10 9 7 2 15 1 10 15 2 15 4 13 10 10 9 2
30 0 1 13 10 10 9 0 2 4 13 10 9 1 12 9 1 3 12 1 9 2 12 9 2 12 9 2 10 9 2
65 7 0 1 13 15 1 15 1 10 9 1 9 2 16 1 11 4 13 10 0 9 1 10 9 1 13 10 9 13 1 10 9 0 2 1 10 9 1 10 9 13 3 15 1 10 9 2 1 9 0 2 1 10 9 1 9 7 9 15 15 13 1 10 9 2
30 11 11 1 11 11 2 9 1 11 2 4 13 10 11 13 1 10 9 1 9 3 3 0 1 3 4 13 11 11 2
37 10 15 4 13 9 1 9 2 10 0 0 11 4 13 13 10 10 9 1 9 3 1 10 11 1 11 2 7 3 4 3 13 10 9 3 0 2
22 10 9 1 13 10 9 0 1 11 11 11 2 1 11 2 9 0 2 13 3 0 2
41 3 3 15 13 10 0 9 1 10 9 3 1 11 2 9 12 2 7 10 0 9 11 11 3 1 10 11 15 4 13 4 13 1 3 13 10 9 1 10 9 2
15 1 9 1 11 11 15 15 15 4 13 1 10 10 9 2
42 10 0 11 13 3 10 0 9 1 11 11 2 10 2 11 1 9 2 15 12 9 3 13 2 3 1 10 11 2 13 13 1 9 7 9 10 9 1 10 9 0 2
11 9 15 15 13 3 13 1 10 0 9 2
12 7 11 2 1 9 11 2 15 4 3 13 2
6 11 2 10 9 0 2
12 11 1 10 9 1 13 15 15 4 3 13 2
18 4 13 11 1 9 2 13 15 3 1 9 1 0 9 7 0 9 2
16 4 13 16 15 13 2 3 2 10 10 0 9 1 10 9 2
27 15 4 13 12 9 0 2 1 15 11 15 11 4 13 1 9 13 2 3 2 1 13 15 10 10 9 2
32 10 0 9 0 4 4 13 1 9 1 4 13 13 1 10 9 0 1 11 2 0 9 1 10 11 7 9 0 1 10 9 2
17 10 15 3 13 9 1 13 15 3 3 13 15 7 10 10 9 2
36 16 4 13 1 13 15 16 3 13 1 13 2 11 4 13 3 1 11 10 9 1 9 0 2 11 2 10 9 7 9 2 1 3 13 15 2
7 9 13 1 9 1 11 2
13 1 11 10 0 9 1 9 13 12 9 1 9 2
9 16 13 10 9 2 3 4 13 2
26 1 13 11 4 13 3 11 1 13 15 1 9 16 4 4 13 1 13 1 10 9 0 1 10 11 2
5 10 9 13 0 2
12 11 4 4 13 10 9 7 10 9 1 11 2
18 10 3 1 13 15 1 13 3 0 7 1 13 15 1 13 10 9 2
8 9 1 10 15 15 13 11 2
16 15 13 10 0 9 16 11 4 4 13 10 9 1 10 9 2
25 13 0 2 10 9 13 15 10 9 2 4 13 3 3 11 2 16 15 13 10 9 13 1 15 2
30 15 13 1 13 7 2 13 16 13 1 10 9 0 7 13 16 11 4 13 10 9 1 10 9 2 10 9 13 0 2
15 3 16 10 9 1 11 13 3 0 1 3 13 0 9 2
17 4 13 1 10 9 10 10 9 2 10 10 9 2 10 10 9 2
50 10 9 0 4 13 10 9 2 13 10 9 0 2 3 13 16 15 13 10 9 3 4 3 13 10 9 1 13 15 1 9 0 2 16 10 10 9 4 13 15 1 13 10 9 2 3 1 13 15 2
14 3 7 15 13 0 9 1 10 9 7 15 15 13 2
14 3 13 9 1 9 2 3 15 4 13 15 1 9 2
25 9 16 10 9 15 15 13 3 10 9 0 15 4 13 1 10 9 7 13 15 3 1 0 9 2
11 13 10 9 1 10 9 10 9 1 9 2
8 11 13 16 3 13 10 9 2
36 3 2 13 3 16 7 15 7 10 9 11 13 2 16 13 10 9 0 2 1 13 1 10 9 1 10 9 10 9 1 11 7 10 9 0 2
34 1 10 9 0 2 1 12 7 12 9 1 9 1 10 9 2 10 9 7 10 9 1 10 11 4 13 1 10 1 3 1 10 9 2
16 7 15 13 1 9 10 9 1 10 9 4 13 1 0 9 2
15 16 10 9 0 13 13 1 3 13 15 15 3 13 0 2
30 3 1 10 9 3 0 15 13 1 10 9 10 10 9 1 10 9 4 3 13 1 10 9 16 1 0 9 4 13 2
22 1 10 1 3 1 10 9 7 1 10 9 0 2 3 15 4 13 16 15 13 3 2
32 10 0 9 13 1 13 15 11 2 0 9 1 11 2 1 13 15 10 9 7 15 13 1 13 10 9 1 9 1 10 9 2
17 11 13 3 0 1 13 2 13 16 15 4 13 1 9 12 9 2
17 10 9 3 13 1 10 0 9 1 10 10 9 3 1 10 9 2
12 15 13 7 13 1 13 15 0 10 3 0 2
20 11 13 0 9 2 13 15 13 3 3 1 12 9 1 9 3 0 7 0 2
14 3 13 10 9 1 13 10 0 9 1 10 9 0 2
13 3 2 7 11 13 0 9 1 11 7 15 13 2
6 10 9 0 3 13 2
5 9 1 10 9 2
5 9 1 10 11 2
29 9 11 2 16 13 0 16 10 9 1 10 10 9 3 13 10 9 7 10 9 2 10 9 13 9 1 10 9 2
31 15 13 1 10 9 1 13 11 2 13 12 9 2 4 13 13 10 9 15 3 15 13 2 15 3 13 7 3 13 3 2
30 3 16 10 9 1 10 9 2 10 9 1 10 0 9 1 11 11 7 11 11 2 13 3 10 0 9 1 10 9 2
20 3 16 10 9 1 10 9 3 4 13 1 10 9 10 9 2 9 2 9 2
8 3 16 10 9 15 13 0 2
48 3 11 11 2 1 10 9 2 2 10 9 0 1 10 9 1 11 7 0 1 11 2 4 13 1 9 10 10 9 1 10 12 7 4 13 3 2 1 10 9 1 10 0 9 1 10 9 2
30 1 3 10 0 9 2 0 9 0 1 13 10 9 0 2 3 13 3 1 10 9 9 2 4 13 1 9 1 9 2
20 4 13 1 10 0 9 2 10 9 7 10 9 1 10 10 9 15 4 13 2
26 4 13 10 0 9 2 3 9 11 4 13 9 1 10 9 1 10 9 2 2 3 0 1 10 9 2
29 13 1 9 2 16 10 11 2 10 9 0 1 10 9 0 2 3 4 13 16 10 9 13 0 1 13 10 9 2
8 7 3 0 1 13 10 9 2
6 3 10 12 9 9 2
18 11 2 3 10 9 1 11 2 7 10 9 0 3 4 13 1 13 2
39 10 11 3 15 13 2 7 10 11 13 3 13 2 1 13 1 11 11 2 1 10 9 2 2 9 0 1 11 1 10 12 7 15 1 10 11 1 11 2
7 10 11 3 13 13 9 2
30 2 15 13 16 10 9 13 3 0 2 13 10 9 0 2 3 16 13 10 3 9 1 10 9 1 9 1 10 9 2
18 9 1 9 2 10 9 13 10 12 9 1 10 9 1 3 13 11 2
8 11 2 0 9 1 11 11 2
9 2 7 3 4 13 10 9 2 2
7 11 11 13 13 10 9 2
9 4 13 15 1 10 12 9 0 2
23 11 2 10 12 9 1 9 4 13 10 9 3 7 3 0 2 13 0 1 10 0 9 2
41 10 9 13 1 10 9 11 4 13 1 12 9 1 10 9 2 10 0 9 15 10 9 4 13 10 9 1 13 1 13 3 1 9 2 9 1 10 10 9 0 2
22 10 9 0 2 9 1 10 9 0 0 1 10 9 1 12 9 7 12 1 12 9 2
47 11 15 13 10 9 1 9 1 9 7 3 4 13 2 1 9 1 12 1 10 12 9 2 12 1 10 12 9 7 3 10 0 9 1 9 3 1 10 12 9 13 1 10 9 1 12 2
28 1 3 4 13 10 9 0 1 10 9 15 4 13 1 12 13 10 9 3 0 1 10 12 9 0 1 12 2
28 11 4 13 1 10 9 12 9 13 10 9 0 1 9 2 1 10 1 3 1 10 10 12 9 7 12 9 2
42 1 10 9 1 13 0 10 9 2 1 9 9 1 13 15 1 10 9 1 10 12 2 3 1 9 1 10 0 9 13 1 10 12 9 7 9 7 13 1 10 9 2
39 3 3 10 9 4 4 13 1 10 9 2 3 3 0 3 3 0 1 10 9 2 13 11 2 2 16 3 1 10 9 16 4 13 1 10 10 11 11 2
30 10 9 1 10 9 4 4 3 1 9 13 1 9 1 10 0 9 1 9 2 15 13 13 1 10 9 1 9 0 2
30 3 16 10 9 13 13 2 13 15 10 9 0 1 13 10 9 1 10 9 1 10 0 9 13 1 9 3 3 3 2
27 1 10 0 9 11 2 0 9 0 2 0 7 0 1 10 9 1 9 2 1 10 9 15 13 13 15 2
22 4 13 11 11 10 0 9 1 10 9 1 10 9 1 10 9 0 2 1 11 12 2
39 7 1 3 13 10 9 2 1 10 9 15 2 13 2 1 15 2 15 13 10 13 2 10 9 2 10 9 0 15 15 13 3 3 3 10 9 13 13 2
16 13 12 9 11 11 2 10 0 9 1 9 0 1 10 11 2
9 7 10 9 0 2 9 1 9 2
24 7 3 15 15 15 13 3 16 13 1 4 15 13 2 3 1 13 1 10 9 1 10 9 2
7 13 4 13 2 13 2 2
26 3 1 15 13 13 15 1 10 9 2 16 10 9 13 15 1 10 9 2 16 10 9 15 13 3 2
7 7 15 11 13 1 13 2
12 2 4 3 13 3 2 1 10 9 1 9 2
21 4 13 1 10 9 1 11 1 11 11 2 15 13 2 3 13 1 13 0 2 2
7 7 15 3 13 1 13 2
31 2 10 9 1 10 9 1 11 11 7 10 2 9 2 1 10 10 9 2 1 11 11 15 15 4 13 3 1 3 2 2
14 11 11 13 10 9 0 1 10 9 1 9 1 9 2
40 9 1 10 10 9 2 9 1 11 2 11 11 13 1 0 9 1 13 15 3 10 9 1 9 0 7 10 9 0 1 10 9 13 1 10 9 1 10 9 2
38 13 15 10 9 0 15 15 13 9 0 2 15 13 1 9 0 2 7 3 1 9 7 9 13 2 13 2 13 2 13 9 0 2 3 0 1 9 2
28 10 9 1 11 1 10 9 1 10 11 13 9 0 2 10 9 1 10 9 1 10 11 7 1 9 1 9 2
19 10 9 13 1 10 9 1 10 9 1 11 2 1 15 1 11 7 11 2
14 3 2 1 10 9 4 13 10 9 2 13 11 11 2
12 10 9 1 10 9 13 3 10 9 1 9 2
31 7 11 11 3 13 10 10 9 1 9 2 13 15 10 9 16 15 15 13 10 9 2 2 16 3 1 15 13 1 13 2
13 7 4 3 13 2 16 3 15 15 13 3 15 2
19 13 1 13 15 2 15 13 1 11 2 13 1 10 9 2 13 10 9 2
5 7 13 3 0 2
14 3 13 16 15 13 10 10 9 2 7 4 13 3 2
13 11 13 7 15 13 10 9 1 10 10 9 2 2
23 11 13 7 11 11 13 10 9 2 13 3 1 10 9 2 7 3 13 16 15 4 13 2
23 11 13 0 2 7 15 3 13 10 9 2 13 10 9 0 2 13 15 3 7 3 2 2
24 0 16 10 9 0 3 4 13 15 1 10 9 7 16 10 9 13 1 13 15 9 1 9 2
37 0 9 0 15 1 10 9 2 10 9 1 9 15 13 1 10 9 2 13 1 10 9 1 10 9 15 13 0 1 10 9 7 3 1 10 9 2
9 10 11 2 15 3 13 1 9 2
30 11 11 2 3 13 1 9 1 10 9 2 1 10 9 13 16 13 10 9 1 10 9 7 13 15 15 13 3 2 2
11 11 7 11 2 13 1 10 9 1 11 2
5 9 1 11 11 2
14 1 3 13 15 1 9 2 1 3 13 15 1 9 2
9 1 13 15 10 9 10 10 9 2
51 3 15 4 13 1 9 11 11 2 7 6 16 13 1 16 13 12 9 7 9 2 16 10 9 2 15 3 13 1 11 2 1 11 2 15 13 1 9 7 15 13 1 15 2 16 13 10 9 1 9 2
22 11 15 13 3 1 10 11 11 2 13 3 10 9 7 13 16 4 13 10 12 9 2
55 3 16 10 9 13 9 1 10 9 2 10 9 15 13 1 10 9 0 2 10 9 13 1 13 15 13 9 2 1 11 2 1 12 9 1 9 2 2 7 10 10 9 15 3 15 4 3 13 2 7 3 10 10 9 2
14 13 1 10 9 3 16 13 10 11 15 15 13 0 2
5 3 15 13 3 2
25 13 3 15 13 15 15 15 13 1 13 2 10 9 0 11 2 7 15 13 1 10 0 9 2 2
6 9 0 2 1 9 2
22 10 9 2 9 2 13 1 10 11 11 1 11 2 3 15 13 10 0 9 1 11 2
9 2 10 9 15 15 4 13 13 2
5 7 3 13 2 2
68 3 4 13 10 0 11 7 10 0 11 2 9 12 1 10 9 1 3 2 1 10 9 1 15 4 13 1 9 2 1 15 3 4 3 13 9 2 1 15 13 10 10 9 2 15 13 0 2 15 13 3 2 15 13 1 10 9 7 3 13 0 16 13 0 7 0 2 2
14 1 15 13 10 9 1 13 15 15 13 2 1 9 2
17 11 11 2 11 2 11 2 10 10 9 15 1 3 13 10 15 2
13 15 1 9 2 3 1 10 11 1 11 0 0 2
7 10 9 1 10 11 11 2
9 10 9 2 10 11 13 10 9 2
8 3 13 10 9 1 11 12 2
16 10 9 1 9 1 10 9 0 13 10 9 1 9 3 0 2
31 10 11 4 3 13 10 9 1 11 12 2 16 10 9 15 13 1 11 2 12 9 2 7 11 2 12 9 1 9 2 2
8 1 11 12 2 10 9 0 2
42 10 9 0 0 2 3 1 11 7 11 2 4 4 13 1 11 2 12 2 1 10 12 2 2 11 7 11 1 10 12 2 11 2 12 9 1 9 2 1 10 12 2
29 11 11 13 10 0 9 1 13 10 9 0 7 13 10 0 9 1 13 10 9 1 9 2 13 0 3 10 11 2
34 3 1 15 2 4 13 10 9 0 11 11 2 12 9 2 12 2 2 11 11 2 9 2 12 2 7 11 11 2 12 2 12 2 2
21 10 9 1 11 3 0 1 12 9 2 12 9 2 13 13 10 9 1 10 9 2
20 1 10 12 2 10 9 1 11 2 13 1 11 2 13 3 0 1 12 9 2
34 1 10 11 1 10 12 2 11 13 1 9 0 10 9 1 10 12 9 2 13 1 11 2 1 13 15 16 4 4 13 10 0 9 2
35 1 10 11 12 2 1 10 12 2 10 9 4 13 1 12 9 1 10 9 1 11 7 11 2 1 9 1 10 9 2 13 10 9 2 2
6 11 9 1 10 12 9
5 13 1 9 11 0
5 13 3 12 9 2
3 12 9 2
2 12 2
8 10 11 0 2 10 11 13 2
6 9 0 1 10 12 2
6 13 11 10 0 11 2
20 1 10 0 9 11 2 10 0 9 1 10 9 1 10 11 15 15 4 13 2
17 9 1 9 2 13 11 2 13 11 2 2 0 9 1 9 2 2
39 10 12 9 13 1 0 10 9 0 2 9 0 1 9 3 3 13 2 3 11 11 13 10 9 1 10 11 1 13 1 10 9 16 13 15 10 0 9 2
35 3 2 1 9 15 13 3 12 2 15 1 10 12 9 15 13 11 11 2 9 2 2 1 10 9 1 9 7 15 13 13 1 10 9 2
11 2 15 4 13 13 15 1 10 9 2 2
34 1 10 9 12 9 15 10 9 1 10 9 0 3 4 3 13 1 9 10 2 16 3 11 11 2 9 2 13 10 9 1 9 9 2
21 1 10 9 10 9 0 7 10 9 15 13 15 7 3 15 4 13 9 1 15 2
20 10 0 9 16 10 9 1 9 13 1 9 15 13 1 11 2 12 9 3 2
8 0 11 11 2 11 2 12 2
12 1 0 10 9 9 2 10 0 9 1 11 2
9 10 9 15 13 15 13 3 3 2
3 13 11 2
10 2 13 10 9 2 4 13 10 9 2
6 3 13 3 10 9 2
7 7 3 13 1 11 2 2
8 13 13 10 0 9 1 13 2
16 11 13 10 9 13 1 10 9 2 9 2 7 1 10 9 2
49 10 10 9 1 0 9 7 0 9 15 13 1 10 9 1 10 9 2 9 1 10 9 1 10 9 2 15 13 10 15 1 10 9 1 9 2 16 3 15 4 3 13 1 12 9 1 10 9 2
44 13 1 9 1 10 9 2 16 10 10 9 2 12 2 0 2 13 16 10 10 9 13 1 10 9 2 3 1 15 4 3 13 16 2 11 11 4 13 10 9 15 13 2 2
26 1 9 16 11 11 2 7 6 2 1 11 11 2 10 9 1 10 9 0 2 13 10 0 9 0 2
35 2 11 7 15 13 1 10 0 9 2 9 0 2 3 10 10 9 15 4 13 1 13 15 1 10 0 9 15 13 9 2 10 0 2 2
14 1 9 16 10 11 1 10 11 13 10 9 1 9 2
16 11 13 1 11 2 11 2 2 11 1 11 7 11 1 11 2
26 2 16 15 13 13 1 10 9 1 15 2 13 9 2 13 10 9 1 10 9 2 13 10 0 9 2
9 3 1 10 9 10 11 1 11 2
19 3 10 11 15 4 13 15 10 9 16 11 13 3 1 9 1 10 9 2
27 10 9 3 0 1 10 12 1 13 2 9 1 9 15 13 0 2 13 3 3 3 2 7 13 3 15 2
21 10 9 1 11 13 1 10 9 0 1 11 11 2 1 10 10 9 1 0 9 2
15 2 4 13 3 2 7 15 15 4 13 2 3 13 13 2
11 3 1 10 12 9 15 13 7 3 3 2
15 3 1 11 2 10 10 9 13 10 9 2 10 15 3 2
13 15 4 13 1 13 16 4 13 16 13 1 9 2
20 4 4 13 1 9 2 13 3 3 16 11 2 10 9 2 15 4 13 2 2
7 3 13 1 13 15 13 2
13 12 10 9 1 10 9 1 10 9 1 10 12 2
12 3 13 2 1 9 0 2 1 3 12 9 2
18 9 1 9 2 1 10 11 2 9 1 10 9 11 2 9 1 9 2
10 11 2 10 9 13 10 9 1 9 2
6 9 0 1 10 12 2
11 10 11 1 9 13 10 9 1 9 9 2
11 2 6 11 2 15 4 13 10 9 2 2
27 11 2 13 10 12 1 9 12 9 7 1 10 9 11 1 11 13 3 1 11 11 10 9 1 10 9 2
19 1 10 9 13 3 9 0 1 9 1 9 2 10 9 0 1 10 11 2
27 10 9 1 9 0 2 0 1 9 2 13 1 10 9 2 3 13 10 9 1 13 1 13 10 9 11 2
28 10 9 11 11 2 10 9 0 15 15 4 13 12 9 3 13 15 1 13 10 9 0 2 3 3 15 13 2
12 4 13 3 13 1 11 1 3 13 10 9 2
24 7 10 11 2 9 1 10 9 0 2 13 1 10 12 9 1 13 0 1 10 9 3 0 2
13 11 4 13 0 9 2 11 2 13 15 2 11 2
7 0 2 0 2 9 2 2
8 7 15 2 3 2 15 13 2
8 2 11 2 6 2 11 2 2
17 2 13 3 9 3 2 13 3 1 9 2 15 13 2 13 11 2
35 2 8 8 8 8 2 13 1 9 10 11 15 1 9 2 9 1 9 7 10 9 1 10 9 1 10 11 11 11 13 9 1 13 15 2
7 2 3 15 13 10 9 2
11 2 6 11 2 15 4 13 10 9 2 2
29 10 0 9 1 10 9 13 11 1 10 15 1 9 0 2 1 10 9 1 10 9 1 9 1 10 9 1 11 2
10 11 4 13 1 10 9 1 10 9 2
32 7 10 9 1 9 4 13 16 10 9 2 15 4 4 13 10 9 1 9 1 11 2 15 4 13 13 15 10 9 1 11 2
8 15 3 15 4 13 1 9 2
25 2 3 2 1 15 3 4 13 1 13 10 15 15 13 3 2 13 3 10 9 1 10 9 2 2
18 15 4 13 13 15 15 1 9 16 13 1 13 15 13 10 9 2 2
14 1 9 15 4 9 2 16 11 4 13 1 10 9 2
17 2 13 1 3 7 4 15 13 3 1 9 13 16 10 15 13 2
5 3 15 13 13 2
19 3 4 3 13 1 10 0 7 4 13 0 1 10 9 3 1 9 13 2
8 6 2 3 10 9 3 2 2
24 3 4 4 13 1 10 12 13 1 10 9 7 15 3 13 3 10 10 9 0 2 12 2 2
31 3 13 9 16 13 3 7 1 10 9 15 4 13 16 10 9 2 0 7 0 2 13 10 9 1 9 1 13 10 9 2
13 3 1 9 2 3 2 4 13 10 9 11 11 2
22 13 10 9 1 10 9 13 3 1 10 9 0 2 16 13 10 10 0 9 1 12 2
28 3 1 10 0 11 11 2 3 15 4 3 13 1 10 9 3 13 1 13 3 10 0 2 9 2 1 9 2
25 10 9 15 4 13 1 10 11 1 11 1 10 9 7 10 10 0 9 2 10 9 0 11 11 2
39 10 9 3 13 1 10 9 1 10 9 2 13 16 10 9 3 9 2 3 1 10 9 2 4 13 3 9 0 7 3 4 13 10 9 0 1 10 9 2
27 3 10 0 9 11 2 3 0 1 10 9 1 10 9 1 10 12 9 1 9 2 4 13 3 1 9 2
39 3 15 4 13 16 1 11 10 9 4 3 13 2 1 10 9 0 1 10 0 11 2 15 1 12 13 10 0 9 1 9 1 10 0 11 2 12 2 2
21 0 10 0 9 2 10 11 2 12 2 2 15 11 11 2 0 1 10 10 12 2
26 1 10 9 10 9 0 4 13 3 1 9 9 2 7 3 3 1 10 9 3 15 4 13 1 3 2
21 11 11 4 13 11 11 1 10 12 1 11 1 10 9 0 9 2 15 15 13 2
18 13 10 9 15 10 11 11 13 1 0 7 15 10 11 3 3 13 2
6 11 11 1 10 11 2
6 11 13 10 11 9 2
11 12 9 1 10 11 2 1 9 3 11 2
8 11 11 2 10 9 1 11 2
6 15 13 10 9 0 2
17 10 11 13 10 11 9 9 1 10 9 0 7 13 10 11 9 2
45 1 10 9 1 10 11 13 3 15 1 10 11 11 2 12 12 2 9 1 12 9 7 1 10 0 9 1 10 9 1 10 9 1 10 9 1 10 9 0 1 10 12 1 9 2
24 0 7 0 11 4 13 1 9 1 10 12 1 10 0 9 13 1 10 9 10 9 11 11 2
63 10 11 2 13 3 1 10 12 12 12 13 1 10 9 0 1 11 2 11 2 11 7 11 2 1 9 11 11 2 11 7 11 7 9 13 1 11 1 9 11 7 11 2 15 4 13 1 9 9 1 11 9 1 10 9 1 9 1 9 0 1 11 2
30 10 0 9 13 10 11 15 13 10 9 7 3 13 9 1 10 9 13 1 10 9 1 10 9 1 11 13 1 9 2
34 1 10 9 1 10 0 9 10 11 13 1 10 9 0 1 13 10 9 1 10 9 1 10 11 11 2 12 2 15 13 1 0 9 2
41 3 15 13 1 0 11 1 13 10 9 1 10 12 12 1 10 9 15 13 10 9 0 1 10 9 1 9 0 1 11 2 12 2 13 1 10 9 1 10 9 2
12 10 9 13 9 7 9 1 9 1 10 9 2
5 13 11 7 11 2
2 15 2
35 9 0 1 10 11 1 11 2 1 11 2 3 10 9 1 11 11 4 4 13 1 12 12 1 10 11 11 2 9 1 10 9 11 0 2
11 12 10 9 13 7 12 13 1 10 9 2
20 1 10 12 1 10 0 9 9 0 1 11 1 9 1 9 1 9 1 11 2
12 1 10 12 1 10 9 9 1 10 11 11 2
8 9 1 9 1 11 3 13 2
12 9 0 1 10 11 1 10 9 1 10 11 2
7 12 12 1 9 1 11 2
16 1 11 10 9 1 10 9 0 4 13 10 11 1 12 12 2
18 9 1 11 7 11 11 1 10 9 7 1 11 1 10 9 1 11 2
9 1 10 11 10 11 11 1 9 2
24 11 2 13 1 13 10 11 0 1 10 9 15 11 11 4 13 1 9 1 10 11 1 11 2
31 10 0 11 4 13 10 9 2 11 11 2 13 10 11 1 12 12 2 12 12 2 12 12 2 12 12 2 12 12 2 2
43 1 0 9 2 15 10 9 4 13 1 10 9 2 11 2 1 3 1 9 0 1 10 0 12 9 2 10 9 0 11 11 2 15 4 13 1 10 9 0 1 10 9 2
31 3 10 11 13 1 11 1 11 3 4 13 10 0 9 3 1 10 9 11 1 9 1 11 1 10 12 1 10 12 9 2
21 10 9 2 13 10 9 1 10 9 1 11 2 1 9 1 10 9 1 10 9 2
9 9 2 13 10 9 1 10 9 2
6 9 11 7 9 0 2
8 10 9 13 1 10 9 11 2
7 13 10 9 1 10 9 2
45 3 10 9 1 10 9 1 9 11 7 11 2 11 2 11 2 11 2 11 2 11 2 7 10 9 1 10 9 2 11 2 11 7 11 2 13 10 9 1 10 11 2 11 11 2
73 10 9 9 4 3 9 13 10 9 1 3 2 13 1 13 9 7 13 10 10 9 1 10 9 1 11 1 9 2 7 2 1 10 9 0 2 13 1 9 1 11 1 10 12 7 1 9 1 9 7 13 0 13 16 15 13 1 10 9 3 3 1 10 9 2 3 1 10 9 11 1 11 2
51 15 13 10 9 2 0 0 2 1 12 9 2 13 1 10 9 2 1 13 7 1 13 3 7 10 9 3 4 13 1 13 3 2 1 10 9 1 12 9 2 15 15 4 13 1 10 12 1 9 9 2
12 11 4 13 1 13 10 9 1 10 10 9 2
7 1 11 15 4 13 3 2
29 2 10 9 4 13 1 10 9 12 9 2 13 10 9 0 2 16 15 13 0 1 12 2 12 9 0 1 9 2
17 15 13 9 15 13 13 9 0 7 3 10 9 13 3 0 2 2
48 1 9 1 10 9 1 11 2 1 9 1 10 9 1 11 2 2 13 1 3 2 4 3 13 10 9 1 10 9 2 2 10 9 4 13 10 9 1 9 2 3 4 13 9 1 9 0 2
35 7 1 10 9 2 10 9 1 10 9 13 10 9 1 10 0 9 1 9 1 10 9 1 10 9 1 9 10 9 1 9 11 7 11 2
26 10 9 13 3 0 2 3 10 9 4 13 13 15 1 9 3 0 7 0 1 10 9 1 10 11 2
15 7 10 9 11 13 16 3 1 10 9 10 11 13 0 2
8 13 3 10 9 1 10 9 2
10 11 11 13 11 15 1 10 9 0 2
6 9 11 13 10 11 2
35 10 9 1 11 11 2 10 0 9 1 10 13 3 1 9 1 11 2 13 1 13 10 2 11 11 2 2 1 9 1 11 11 9 12 2
17 13 10 9 15 1 10 12 13 10 9 1 11 2 13 1 11 2
27 11 2 3 2 4 4 13 0 1 10 9 13 1 10 2 11 2 7 10 2 11 2 7 4 4 13 2
22 3 11 11 2 10 9 7 9 2 4 4 13 1 13 10 9 1 9 1 10 9 2
29 3 15 13 1 10 9 7 3 15 13 0 9 3 16 10 9 0 13 10 10 0 9 2 7 15 13 10 9 2
26 3 2 1 9 3 13 1 10 9 2 15 13 10 9 1 10 0 9 1 10 9 2 10 0 9 2
9 7 3 2 15 13 10 9 9 2
3 10 12 2
9 1 10 12 2 12 2 12 9 2
9 1 10 12 2 12 2 12 9 2
8 1 10 12 2 12 2 12 2
7 10 9 13 1 12 9 2
5 11 1 10 11 2
7 9 0 1 10 11 11 2
7 9 2 11 0 1 11 2
29 13 10 9 1 10 9 1 9 0 2 15 13 1 10 11 11 2 1 10 11 1 11 13 3 1 10 0 11 2
13 11 11 2 0 1 11 2 13 1 10 0 9 2
6 1 10 9 11 11 2
2 9 2
16 9 13 1 11 11 2 10 9 0 13 1 10 9 1 9 2
12 4 4 13 1 10 9 1 10 9 1 9 2
9 9 2 1 11 9 1 11 11 2
7 13 11 2 9 1 11 2
45 9 11 2 10 9 1 11 2 7 3 10 9 1 9 0 2 4 13 10 9 1 10 0 9 1 10 11 11 13 1 10 9 0 10 11 11 11 2 9 1 11 1 10 9 2
25 11 11 2 13 1 11 12 9 3 13 1 9 0 15 13 10 9 2 4 3 13 10 0 9 2
38 1 9 4 13 3 10 9 0 2 3 10 9 0 4 13 1 13 15 1 15 0 3 10 9 1 10 9 1 9 13 3 3 0 1 1 9 10 2
48 3 13 1 10 9 0 2 13 16 10 9 13 1 11 1 10 9 2 7 1 11 4 13 15 2 1 10 9 1 9 1 11 7 11 1 15 13 10 10 9 1 10 9 13 1 11 11 2
10 10 9 12 1 9 15 4 13 9 2
7 4 13 11 1 10 9 2
18 2 4 13 1 10 9 1 10 9 2 16 3 13 3 3 1 13 2
13 13 10 12 9 1 10 9 7 3 10 0 9 2
6 3 3 15 13 3 2
10 1 12 9 1 9 4 13 1 13 2
30 1 10 9 15 13 1 10 9 13 16 13 1 10 9 0 1 10 9 7 9 1 9 4 13 10 0 9 1 9 2
16 4 13 10 10 9 1 9 11 15 15 4 13 1 15 2 2
19 1 9 1 11 2 11 4 4 13 1 11 15 4 3 13 1 13 0 2
33 11 15 4 13 10 0 9 1 12 16 11 1 12 4 13 1 10 9 10 0 11 15 13 10 9 1 10 9 7 10 0 11 2
10 9 1 10 9 2 1 12 9 2 2
2 12 2
9 11 2 11 2 9 12 2 12 2
16 9 1 9 2 10 9 0 13 10 9 1 10 9 1 11 2
5 11 13 10 11 2
6 2 11 1 9 2 2
17 2 4 13 10 9 2 10 9 13 13 1 9 1 10 11 2 2
31 11 2 10 9 1 10 11 7 10 9 1 11 15 13 9 1 11 11 2 10 15 15 13 10 9 0 2 13 7 13 2
27 2 13 0 1 10 9 0 1 10 11 2 15 13 16 10 10 9 4 13 1 10 9 3 0 7 0 2
14 7 3 13 16 15 15 13 2 13 16 4 13 2 2
24 15 13 1 10 9 13 1 15 4 13 9 1 10 9 1 10 12 9 3 13 1 10 11 2
11 3 0 7 0 2 1 10 9 1 11 2
9 2 13 16 10 9 4 3 13 2
16 13 1 13 10 9 3 0 2 2 13 3 11 13 10 9 2
17 7 10 9 0 3 13 3 1 10 9 1 10 9 1 10 11 2
23 10 10 9 13 3 0 7 10 9 13 3 1 10 9 13 1 10 11 1 10 0 9 2
24 2 16 10 9 13 10 0 9 4 13 0 2 3 10 9 15 4 13 10 3 3 13 2 2
28 3 11 3 4 13 10 9 1 10 10 0 9 0 1 10 11 1 10 12 2 13 1 11 12 1 11 11 2
25 7 3 13 16 10 0 9 1 11 7 11 4 13 3 10 9 1 10 9 1 10 9 1 11 2
10 10 9 13 16 10 9 13 10 9 2
21 10 9 7 10 9 13 1 10 0 9 13 0 9 1 12 9 13 1 10 9 2
18 10 9 2 3 2 4 13 10 9 7 4 4 13 3 2 1 9 2
5 15 13 9 2 2
16 3 10 11 3 15 13 3 2 3 1 10 9 1 11 11 2
17 3 15 13 1 10 9 10 9 1 10 9 1 10 11 2 3 2
26 2 4 3 13 3 15 4 13 11 2 3 15 13 3 1 13 1 10 9 0 15 15 15 4 13 2
31 13 16 15 4 13 1 9 10 10 9 7 10 10 9 2 15 13 3 0 13 3 1 10 9 0 16 15 13 9 0 2
11 13 10 15 16 1 9 13 10 11 2 2
26 10 9 1 10 9 1 10 9 0 4 13 2 1 11 2 2 1 10 9 1 9 1 10 9 2 2
8 10 9 1 10 11 13 3 2
23 2 12 9 3 13 10 10 9 1 9 1 11 11 7 3 1 15 13 3 1 10 9 2
15 3 15 13 9 1 10 9 7 1 10 11 15 13 9 2
14 7 9 7 9 4 13 13 10 0 0 9 1 9 2
13 13 0 15 1 10 9 1 9 1 10 9 2 2
46 7 2 16 13 0 16 15 13 1 10 9 1 9 2 13 3 0 16 10 9 3 4 4 13 1 10 11 13 16 11 2 3 4 13 15 1 10 9 1 10 9 2 3 13 3 2
19 2 10 9 3 4 13 10 0 9 2 0 2 1 12 9 1 9 2 2
28 1 15 13 10 10 9 3 1 10 9 1 10 9 15 4 13 10 9 1 9 0 7 3 3 1 10 11 2
28 2 3 13 16 13 1 9 10 9 13 10 9 1 11 7 3 3 2 1 9 1 12 9 2 13 11 2 2
21 15 2 16 13 9 7 3 9 1 10 9 2 13 10 15 15 13 0 1 13 2
13 3 2 9 1 10 9 2 13 3 10 9 2 2
38 13 1 9 10 9 0 2 3 10 11 13 1 11 2 13 1 9 10 9 11 11 2 7 13 0 10 9 1 11 11 1 10 0 9 1 10 11 2
25 7 15 1 15 4 13 1 10 9 0 2 3 10 9 7 10 9 0 2 1 13 10 9 2 2
21 10 11 13 1 10 11 7 13 3 11 11 13 1 12 2 11 13 1 10 9 2
29 1 10 0 9 11 2 3 13 1 10 9 1 10 9 7 3 13 1 10 9 2 1 10 11 11 9 1 9 2
17 3 13 9 10 0 11 2 7 15 4 13 1 13 10 10 9 2
15 7 2 16 13 1 10 9 7 10 9 2 4 13 3 2
34 0 9 7 0 9 2 7 15 1 11 2 12 12 2 1 9 1 11 7 1 11 2 13 3 0 1 10 9 2 1 11 7 11 2
22 10 9 1 10 9 2 1 9 11 2 7 3 10 9 1 10 9 3 0 7 0 2
29 11 1 10 0 9 1 10 9 2 13 1 10 9 0 2 3 11 2 11 2 11 2 7 3 0 1 10 15 2
23 11 11 3 13 10 9 3 13 7 3 13 10 9 1 13 15 10 3 1 10 10 9 2
13 11 2 1 0 9 2 15 4 13 3 1 9 2
29 9 1 12 2 1 11 0 1 13 15 3 7 11 11 11 1 9 1 9 1 13 15 1 10 12 0 9 0 2
22 9 13 1 11 2 1 11 7 11 1 13 15 3 10 9 1 10 9 1 10 9 2
14 11 1 9 1 10 9 0 7 0 2 1 0 9 2
14 11 7 11 1 9 2 0 1 13 10 10 9 0 2
3 10 9 2
12 10 0 9 1 10 9 3 13 9 1 9 2
20 10 9 4 13 10 9 1 10 9 1 11 2 1 10 10 9 15 4 13 2
13 4 13 1 10 11 3 12 9 1 11 7 11 2
7 0 2 7 1 3 9 2
22 10 9 13 3 3 1 11 2 10 11 11 0 9 1 9 7 3 0 1 9 13 2
14 10 9 4 13 1 10 10 0 9 10 9 3 0 2
32 10 12 9 4 13 1 9 7 11 15 4 13 10 15 2 1 9 1 11 2 13 1 11 1 10 9 1 9 13 7 13 2
45 10 11 4 13 1 12 9 0 2 13 10 9 0 1 10 12 12 12 15 11 4 13 1 11 11 2 1 13 15 3 10 9 2 11 7 11 13 2 11 3 0 1 9 2 2
43 12 9 1 10 9 1 10 9 2 1 10 9 1 10 9 9 2 13 1 0 9 1 11 1 10 12 2 9 1 11 2 7 1 11 1 10 12 2 9 1 11 2 2
16 9 1 9 0 2 16 10 0 9 15 13 13 1 10 9 2
99 4 13 10 9 1 13 11 7 11 2 1 10 0 9 2 2 13 3 10 9 1 9 1 11 7 11 2 13 10 9 0 2 9 1 11 7 11 13 1 10 9 1 11 2 2 16 10 9 15 4 3 13 10 9 11 15 13 13 3 1 10 9 7 3 1 10 0 9 1 9 1 11 2 2 0 2 1 4 13 2 10 12 9 2 1 10 11 2 3 10 9 1 10 0 9 1 10 11 2
27 3 13 1 9 12 9 0 2 1 10 11 1 10 0 11 1 11 7 1 10 11 11 1 11 1 11 2
15 12 9 1 13 1 9 1 0 9 10 0 9 13 3 2
32 11 4 13 3 11 2 15 13 11 1 9 4 13 10 9 1 11 11 2 10 9 15 3 4 13 10 9 1 10 9 0 2
16 7 4 13 1 10 11 1 10 9 0 1 9 0 1 11 2
10 15 4 13 1 13 15 3 1 11 2
3 10 9 2
9 0 9 1 9 2 11 1 9 2
19 10 9 1 10 11 7 10 9 1 10 9 13 1 9 0 3 1 9 2
12 9 0 1 15 7 3 0 1 10 0 9 2
55 3 1 10 11 10 9 3 10 9 1 10 9 1 10 9 2 11 2 2 0 1 9 1 10 9 1 10 9 2 15 4 13 10 9 1 12 9 0 1 10 9 1 10 11 2 1 0 9 0 1 10 9 1 11 2
32 10 0 9 13 11 11 7 11 11 11 2 13 1 10 9 1 10 9 1 9 1 10 9 1 11 2 3 13 9 1 9 2
22 1 10 9 13 9 11 11 2 13 1 10 9 11 11 2 11 11 11 7 11 11 2
44 11 11 11 2 12 9 2 9 0 2 10 9 0 1 10 9 0 2 4 3 13 10 12 9 1 10 0 9 1 11 2 13 1 10 9 0 0 1 11 2 10 9 0 2
26 10 0 9 2 13 1 10 0 9 2 10 9 3 1 4 13 3 1 10 9 0 4 13 10 9 2
15 2 13 1 0 9 2 10 9 13 15 4 13 2 2 2
38 10 12 9 1 12 9 3 2 11 11 11 2 12 9 2 1 11 2 9 1 11 2 4 3 13 1 10 9 15 13 1 10 9 1 15 15 13 2
14 10 9 13 12 9 7 13 9 12 9 1 10 9 2
17 4 13 1 10 9 0 7 1 10 9 3 15 13 15 1 13 2
25 10 9 1 10 9 1 10 9 3 13 3 9 13 1 10 9 2 1 10 9 2 1 10 9 2
13 15 4 13 1 10 9 1 9 7 3 1 9 2
47 10 12 9 12 11 11 2 1 11 2 7 11 11 11 2 1 11 2 13 1 10 12 9 13 1 10 0 9 1 10 2 11 2 2 15 1 10 9 1 9 1 10 9 1 10 11 2
16 10 9 4 13 1 10 9 1 9 13 1 10 9 1 9 2
13 10 9 1 10 9 4 13 16 13 1 10 9 2
40 10 0 9 0 1 10 9 0 3 1 10 9 13 15 13 1 10 11 12 13 1 10 9 1 10 12 1 10 0 9 1 11 11 7 13 1 10 9 11 2
18 9 7 9 1 9 15 13 1 10 0 9 1 10 9 1 10 9 2
10 0 10 9 0 2 1 9 15 0 2
30 12 10 9 13 1 10 9 1 11 1 10 11 3 4 13 10 9 0 13 1 10 15 3 1 10 9 11 11 11 2
53 2 12 9 1 10 9 0 2 2 13 3 10 11 1 10 11 1 10 9 1 10 12 9 12 2 1 9 1 10 9 1 10 9 13 10 9 3 2 7 1 10 9 0 1 9 2 1 10 9 1 10 11 2
23 1 15 9 1 9 1 9 2 9 2 9 1 9 7 3 10 9 1 10 9 11 11 2
56 9 7 1 10 0 9 1 10 12 9 0 10 9 3 1 11 1 10 9 1 10 9 7 0 1 10 9 1 10 9 1 10 9 0 7 1 10 9 1 9 2 13 2 1 10 9 1 11 2 13 7 13 1 9 0 2
17 1 10 9 1 11 7 11 10 9 1 10 11 13 1 10 9 2
9 2 13 9 1 9 7 9 2 2
14 11 11 13 10 9 1 11 1 10 11 7 11 0 2
65 16 10 9 1 10 11 2 11 11 2 7 10 9 0 1 10 11 2 11 11 2 13 9 1 9 1 9 7 9 2 10 9 1 10 11 2 11 11 2 13 1 10 9 1 10 9 15 2 3 1 9 0 2 13 1 9 7 9 1 9 11 10 0 9 2
8 11 1 10 11 7 11 0 2
39 11 4 13 10 0 9 0 1 11 7 2 13 1 10 9 16 9 7 9 1 15 7 1 10 0 9 3 15 13 2 13 1 10 11 4 4 13 15 2
18 2 10 9 13 2 13 2 13 16 10 11 4 13 1 10 0 11 2
27 1 9 2 1 0 2 3 10 9 1 10 11 4 13 10 9 1 9 0 7 0 7 10 9 0 2 2
13 10 9 1 9 13 10 9 1 9 13 1 11 2
22 2 10 9 0 2 13 11 2 13 1 10 15 15 13 0 10 9 1 10 9 2 2
12 10 9 1 13 13 10 9 1 10 9 0 2
30 2 3 9 2 13 10 9 2 1 10 9 11 11 15 4 13 9 16 10 11 13 1 13 15 1 3 3 13 2 2
48 10 0 9 1 10 9 1 10 11 1 10 11 7 1 10 11 0 4 13 10 9 1 10 9 1 9 15 13 10 9 1 9 7 9 7 15 13 1 13 1 10 9 10 9 1 10 9 2
14 3 2 1 9 1 10 11 15 4 13 10 9 0 2
18 2 3 2 13 11 2 13 0 3 10 9 15 13 1 10 11 0 2
24 13 3 16 1 10 9 2 10 11 13 3 0 1 10 0 9 1 10 9 7 1 10 9 2
28 16 15 13 16 13 7 16 10 10 9 0 13 1 9 1 9 2 10 0 9 15 13 3 10 0 9 2 2
5 2 15 13 2 2
6 7 15 0 13 9 2
29 13 1 10 9 10 9 4 13 10 9 3 16 2 1 10 9 2 10 9 15 4 13 10 9 1 13 10 9 2
29 11 11 2 12 9 2 0 1 10 11 2 16 4 13 10 9 1 9 4 4 13 1 10 9 1 10 9 11 2
14 10 9 1 10 9 15 4 13 1 10 12 10 9 2
20 10 9 4 13 16 1 10 9 0 2 11 15 4 13 13 1 4 13 9 2
22 10 9 1 10 9 2 11 11 2 4 13 1 10 9 1 10 9 1 10 0 9 2
10 10 9 4 4 13 1 10 11 11 2
14 4 13 1 10 9 2 10 9 1 9 15 4 13 2
8 9 13 0 3 1 10 9 2
9 13 0 1 10 9 1 10 9 2
18 11 11 11 2 10 9 0 0 1 11 11 2 4 13 1 9 0 2
37 13 7 13 1 9 1 9 16 2 1 10 0 9 1 9 2 4 13 1 10 9 0 1 10 9 15 4 13 1 10 9 1 9 1 10 9 2
68 11 2 3 15 13 10 9 2 13 10 9 1 10 11 11 1 10 9 11 1 11 7 9 2 16 13 3 1 10 0 9 2 4 13 1 10 9 0 1 13 2 3 1 10 9 2 10 9 7 10 9 1 10 9 1 10 10 0 9 0 2 1 10 9 1 11 11 2
49 11 11 11 2 9 1 10 2 11 2 2 10 9 1 9 3 13 1 10 9 1 10 9 2 15 4 13 1 10 9 1 10 9 0 15 10 9 1 10 10 0 9 4 13 1 10 9 0 2
18 3 4 13 10 9 1 10 9 1 10 15 4 4 13 10 9 0 2
18 11 11 11 4 13 13 1 10 9 1 10 9 0 1 9 7 9 2
28 3 16 4 15 13 13 2 11 15 4 13 1 10 9 7 4 13 1 13 1 9 0 2 13 7 13 9 2
30 10 9 1 10 9 1 11 11 2 13 1 10 9 2 15 4 13 0 16 13 3 10 9 1 10 9 1 10 9 2
49 3 1 13 10 9 3 0 1 9 2 10 9 4 4 13 1 12 9 1 9 7 1 12 9 1 13 1 13 1 10 9 9 1 0 9 2 15 15 4 13 10 12 1 10 9 1 9 2 2
9 11 11 11 4 4 13 1 9 2
16 13 10 9 0 13 1 12 9 3 16 3 4 13 1 9 2
18 1 13 10 9 1 9 4 4 13 3 10 9 1 10 9 1 11 2
18 3 10 9 0 1 10 9 0 13 0 1 13 10 9 1 10 9 2
22 7 3 2 13 16 1 10 9 3 15 13 3 15 1 13 2 4 4 13 10 9 2
30 10 0 9 11 11 2 9 1 9 1 10 9 0 1 11 2 3 4 13 0 13 10 9 7 10 9 1 10 9 2
10 13 3 0 10 9 13 1 10 9 2
19 11 2 3 1 10 9 13 3 1 10 9 2 10 0 9 1 9 0 2
12 10 0 9 0 1 10 2 0 2 9 0 2
6 3 2 3 1 9 2
22 10 0 9 2 13 1 12 9 0 1 12 9 15 2 13 0 1 10 9 1 11 2
11 11 11 2 10 9 2 13 1 10 9 2
16 10 9 13 0 2 3 15 13 10 0 9 2 0 7 0 2
35 1 10 0 2 1 10 9 1 10 9 1 11 11 2 1 12 9 1 10 9 1 11 2 10 9 13 1 10 9 2 10 9 13 13 2
10 11 13 3 10 9 2 13 1 9 2
15 15 13 1 10 9 2 7 10 9 1 10 9 15 13 2
17 10 2 11 2 4 13 10 9 2 10 9 15 4 13 10 9 2
18 1 10 9 15 4 13 7 4 13 2 7 1 10 9 13 10 12 2
25 13 10 9 2 10 9 2 15 13 11 11 2 13 12 9 2 4 13 1 0 1 10 11 11 2
18 15 4 13 1 10 9 1 11 11 1 10 9 2 3 1 10 9 2
17 15 4 3 13 1 9 2 16 15 4 13 3 10 9 1 9 2
31 1 2 13 15 2 4 13 10 9 15 13 1 10 9 1 10 9 2 7 11 11 10 9 13 1 3 4 15 3 13 2
11 3 11 11 13 1 13 2 3 16 13 2
18 10 9 1 10 9 15 13 1 9 1 10 9 10 9 1 10 9 2
7 15 13 0 2 1 3 2
6 3 3 0 7 0 2
24 3 10 0 9 0 13 16 10 9 3 13 3 2 0 2 16 4 13 1 10 9 1 9 2
10 7 10 0 9 13 3 1 13 15 2
6 9 2 9 2 9 2
22 10 9 1 10 9 0 4 13 9 2 1 10 9 1 10 9 0 1 10 9 0 2
42 0 9 2 10 12 9 0 2 4 13 10 9 0 1 11 2 11 11 2 12 9 2 13 13 1 10 9 1 10 9 1 10 9 1 10 9 2 11 1 9 2 2
32 10 9 2 4 13 3 10 9 2 4 4 13 1 10 9 1 10 15 10 9 15 4 13 2 13 3 1 13 1 13 9 2
27 10 12 9 2 1 11 2 13 10 9 1 10 0 9 0 2 11 11 2 12 9 2 13 1 10 11 2
35 10 9 10 9 4 13 7 11 2 15 4 13 1 10 9 1 9 1 10 9 2 4 13 1 9 13 10 9 1 15 1 10 9 0 2
34 9 0 3 1 11 11 2 10 9 0 1 12 9 2 13 10 12 9 1 11 11 1 10 9 1 10 9 1 10 9 1 10 9 2
9 10 9 4 4 13 1 10 9 2
8 10 12 9 10 0 9 0 2
38 10 9 1 12 9 2 11 11 2 7 10 10 9 0 2 11 11 2 13 1 10 9 1 10 9 1 10 9 1 10 9 2 10 9 2 1 11 2
43 10 9 3 3 13 1 11 11 2 10 9 1 12 9 1 11 2 1 9 1 11 1 10 9 2 15 13 1 10 9 1 9 0 10 9 16 16 15 15 13 1 15 2
10 11 2 10 9 0 13 1 13 13 2
8 1 9 15 13 1 9 0 2
7 1 10 11 2 10 9 2
16 10 9 1 10 9 0 3 1 10 9 3 4 13 10 9 2
24 1 10 0 9 11 2 10 9 1 10 9 13 10 9 0 2 1 10 9 0 1 10 9 2
37 9 13 1 9 2 1 10 9 10 9 13 15 13 10 9 1 11 2 10 9 3 10 9 1 11 4 13 9 1 9 1 10 9 1 10 11 2
10 10 9 1 10 9 3 13 16 9 2
10 10 9 2 3 9 0 1 13 15 2
8 7 3 3 10 9 1 11 2
23 10 9 13 1 4 15 13 13 15 1 10 9 2 13 1 10 9 0 1 10 9 0 2
7 4 1 3 13 10 9 2
44 10 9 0 4 3 13 10 12 7 1 10 9 4 4 13 10 9 0 1 10 9 13 1 13 10 9 1 10 9 11 7 2 6 2 3 1 13 15 9 1 10 9 0 2
24 1 9 2 1 10 9 2 10 9 1 9 11 2 1 15 0 2 1 3 13 10 9 0 2
13 3 10 9 0 2 12 9 0 2 13 1 9 2
8 7 3 10 9 2 9 9 2
22 10 0 9 15 4 13 9 2 1 10 0 9 1 10 0 9 1 10 9 1 9 2
40 10 9 1 10 9 13 1 11 11 11 15 4 13 1 10 9 2 3 1 10 9 2 13 1 10 9 10 9 1 10 9 1 10 9 1 9 1 10 9 2
31 2 13 10 9 1 9 2 2 4 13 10 9 13 10 10 9 1 10 9 1 10 9 7 1 10 9 1 10 0 9 2
16 10 9 15 13 2 13 10 9 2 13 9 1 10 10 9 2
15 3 3 15 13 1 13 16 1 10 9 3 15 13 3 2
11 10 9 3 4 13 10 0 7 0 9 2
7 2 3 15 4 13 9 2
23 3 15 13 9 2 2 13 11 11 15 10 9 1 0 7 0 4 13 10 0 1 13 2
5 3 10 9 13 2
11 3 3 13 9 16 1 11 13 9 0 2
19 7 15 1 9 2 13 10 9 2 15 4 3 13 2 7 1 9 12 2
15 10 9 1 11 13 9 15 13 1 10 9 1 10 0 2
14 4 13 9 1 9 13 1 13 15 10 9 1 9 2
22 3 2 10 0 9 2 13 3 3 7 3 16 13 1 0 9 10 9 1 10 9 2
35 15 13 1 10 9 1 10 9 1 12 2 12 9 15 13 1 10 9 11 2 3 10 9 15 13 10 9 1 9 2 7 13 10 9 2
7 3 10 9 0 15 13 2
10 7 10 9 0 3 4 4 3 13 2
30 13 10 0 9 11 1 13 1 9 10 9 1 10 9 1 11 16 15 13 1 13 1 9 10 9 1 10 0 9 2
16 2 10 11 3 4 13 9 1 10 9 1 10 9 0 2 2
27 10 9 3 10 9 0 4 13 1 10 9 1 10 9 1 10 9 13 1 10 9 1 11 2 11 11 2
32 15 13 9 13 1 9 10 11 2 3 15 13 10 9 0 7 3 15 13 1 13 10 11 2 10 10 9 4 13 1 9 2
24 13 3 10 9 15 13 1 10 9 1 11 11 2 3 10 9 13 10 9 1 3 10 9 2
17 10 9 9 11 11 11 13 0 7 0 1 10 0 9 1 9 2
8 2 9 1 9 1 10 9 2
38 3 15 13 2 3 15 13 3 1 15 2 13 13 10 9 1 10 9 1 3 10 9 0 2 10 9 15 4 13 2 10 9 13 10 9 1 9 2
30 6 2 13 0 2 1 11 15 13 10 9 2 7 3 3 1 15 15 15 13 1 10 9 2 1 11 2 1 9 2
10 13 16 1 10 9 13 3 0 2 2
9 9 1 10 9 2 9 1 9 2
3 10 9 2
29 9 2 9 2 9 2 9 0 7 3 2 1 10 9 1 10 2 11 15 13 2 2 3 10 9 1 10 9 2
9 10 9 1 10 9 2 15 13 2
5 9 15 13 3 2
13 1 3 10 9 1 15 15 4 13 3 1 3 2
9 10 0 0 9 15 13 1 11 2
5 15 1 0 11 2
26 10 9 13 1 10 0 9 1 10 9 1 10 9 15 4 13 9 13 13 15 1 9 1 10 9 2
11 9 2 9 0 2 9 2 9 1 9 2
7 3 10 9 13 3 0 2
16 3 1 10 9 1 9 1 10 9 9 4 13 9 7 9 2
16 3 13 0 16 10 0 9 1 9 13 10 9 1 10 9 2
13 1 10 9 15 13 3 1 10 9 13 10 9 2
26 3 3 2 1 10 9 2 10 9 2 16 3 15 13 1 13 10 9 2 4 13 1 10 9 11 2
9 10 9 13 1 10 9 1 9 2
28 3 10 0 9 1 10 2 11 11 2 7 15 1 10 9 0 1 9 2 4 3 13 10 9 1 10 9 2
27 3 0 2 10 9 1 10 9 0 1 10 11 4 13 10 9 1 13 10 9 1 10 9 1 10 9 2
3 15 0 2
9 10 9 3 13 9 1 10 9 2
7 7 1 3 13 10 9 2
10 3 1 10 9 0 2 13 1 11 2
19 10 9 1 0 9 2 1 10 9 15 13 1 11 7 10 0 9 0 2
7 0 9 2 15 1 11 2
28 13 3 2 3 3 2 1 10 9 1 10 9 1 9 0 2 7 1 9 15 15 4 13 1 10 10 9 2
29 1 10 9 1 10 12 9 2 7 3 3 2 13 1 4 13 9 0 1 12 0 1 12 2 12 7 12 9 2
13 9 1 0 1 10 9 1 9 3 13 1 15 2
26 7 15 15 13 1 9 10 9 1 15 1 10 9 15 4 13 1 9 15 1 10 9 1 10 9 2
29 7 10 0 9 1 10 9 13 3 1 0 1 13 7 3 1 13 1 10 9 0 1 10 9 7 10 10 9 2
5 9 7 3 3 2
24 3 1 10 9 1 10 0 9 1 10 11 0 1 13 10 9 0 1 15 1 10 10 9 2
21 13 10 9 13 2 1 13 10 9 1 10 9 0 2 1 10 9 0 11 11 2
9 2 3 10 9 13 10 9 0 2
14 13 10 9 1 10 9 15 3 13 3 0 1 3 2
16 11 4 13 1 10 0 9 13 1 10 0 7 1 10 9 2
13 1 13 10 9 0 15 13 10 9 1 9 2 2
17 10 9 16 10 0 9 13 4 13 1 10 2 9 1 9 2 2
6 10 9 1 10 11 2
19 10 9 1 10 9 1 11 2 9 1 11 1 13 10 9 1 10 9 2
9 2 15 4 13 10 0 9 2 2
9 0 9 1 10 9 1 11 11 2
6 15 4 13 10 9 2
12 2 3 15 4 13 3 10 9 1 11 2 2
43 11 11 2 10 9 1 12 9 13 3 1 10 11 2 4 13 2 7 3 3 2 1 10 10 9 1 10 9 0 10 9 3 1 13 2 1 10 9 1 10 9 0 2
57 3 2 1 10 11 3 1 9 4 13 1 13 10 10 9 0 1 10 9 0 2 9 4 4 13 3 1 10 12 9 1 10 9 11 11 2 11 11 2 11 11 7 11 11 7 1 10 12 9 1 10 9 2 11 7 11 2
16 3 9 4 13 11 2 10 9 1 11 2 1 13 10 9 2
61 1 10 12 2 16 10 9 4 4 13 1 9 1 10 9 1 11 11 2 7 1 10 10 9 10 9 1 11 15 4 13 1 10 9 1 10 9 1 11 3 13 11 2 10 9 0 1 11 2 10 9 11 2 10 10 12 9 11 7 11 2
18 10 9 0 4 13 1 10 9 1 10 0 9 2 13 10 9 3 2
22 7 1 10 0 9 1 10 9 1 12 9 13 2 1 10 10 9 1 11 2 11 2
34 4 13 9 1 10 12 2 16 10 9 15 4 13 3 10 9 11 2 7 4 13 1 13 3 1 10 9 15 4 13 1 10 9 2
10 3 11 2 12 9 2 13 1 11 2
11 10 9 2 3 2 3 3 15 4 13 2
23 13 2 13 1 10 0 9 3 13 2 3 1 10 10 9 2 1 9 7 1 0 11 2
24 10 9 15 15 4 13 1 13 7 15 4 13 3 4 13 15 3 1 10 9 1 10 11 2
23 2 13 12 1 12 2 7 15 3 13 2 13 1 10 9 1 15 1 10 0 9 13 2
6 3 3 15 13 9 2
12 3 10 9 9 1 11 11 7 3 3 0 2
12 11 13 2 3 2 10 9 16 15 13 0 2
13 2 10 12 9 2 3 2 13 10 9 11 2 2
9 10 9 4 13 3 12 9 3 2
10 13 1 10 9 1 9 1 10 11 2
7 1 10 9 3 3 0 2
19 13 10 9 1 10 9 11 2 9 1 10 11 2 1 10 9 1 9 2
22 2 1 9 13 10 9 1 13 15 2 16 11 4 13 13 15 10 9 2 13 15 2
5 13 10 9 11 2
15 10 9 3 4 13 10 9 2 3 15 13 1 10 9 2
24 2 13 9 1 13 3 1 10 9 1 10 9 0 2 1 9 2 15 13 3 1 10 9 2
11 7 3 15 13 10 9 15 3 13 0 2
16 2 4 13 16 1 10 9 15 4 13 9 1 13 1 13 2
7 13 15 15 13 10 9 2
16 1 10 9 1 9 11 11 10 9 4 13 13 3 1 3 2
29 2 10 9 1 11 2 15 4 13 0 9 2 4 13 1 10 12 1 10 9 11 11 2 10 9 1 11 11 2
20 1 10 9 1 11 2 10 9 2 10 9 2 10 9 4 13 0 2 0 2
7 3 0 16 3 15 13 2
7 13 9 11 2 10 9 2
21 11 15 13 13 10 9 2 10 9 1 10 9 7 15 1 10 9 2 10 9 2
18 2 10 11 2 3 15 13 2 3 15 4 13 2 13 10 9 2 2
18 4 13 1 13 15 1 12 2 12 9 2 16 4 13 1 9 2 2
8 0 9 2 3 1 9 0 2
20 3 4 13 9 1 10 9 2 3 1 10 9 9 1 15 13 10 0 9 2
24 11 11 2 10 9 1 15 13 2 4 3 13 1 11 7 1 11 2 3 13 10 10 9 2
16 10 9 1 9 4 3 13 1 10 9 0 10 9 1 11 2
37 10 9 13 3 9 1 10 9 0 1 11 2 13 10 9 1 2 9 2 1 10 9 3 0 1 10 0 9 7 1 10 9 1 10 9 13 2
5 9 2 0 9 2
14 10 9 11 15 13 3 3 1 10 9 1 10 11 2
18 2 9 1 10 9 2 0 9 7 10 0 9 13 1 9 2 2 2
26 10 9 1 11 2 15 13 10 9 1 10 9 1 9 1 11 11 2 13 3 10 9 1 10 11 2
25 13 0 10 9 1 10 9 0 13 1 10 2 9 2 1 13 10 3 3 10 9 1 10 9 2
10 10 9 13 1 10 9 1 10 11 2
44 1 15 2 1 10 10 9 1 10 9 2 4 13 1 10 9 11 1 10 9 1 13 10 9 0 1 10 9 7 10 0 9 1 10 9 1 9 1 10 9 1 10 9 2
11 7 3 9 1 9 1 10 9 1 9 2
21 10 9 15 10 9 13 13 10 9 1 10 9 13 1 13 15 1 10 9 0 2
23 1 10 9 3 13 1 10 2 9 2 1 10 9 0 15 13 9 11 11 7 9 11 2
31 10 9 1 10 0 9 1 9 1 11 4 13 3 9 0 1 10 9 1 10 9 11 2 1 10 0 9 1 10 9 2
10 7 10 9 3 13 3 10 9 0 2
8 13 3 10 9 1 10 11 2
10 2 15 13 16 15 13 10 9 0 2
5 3 13 10 9 2
12 13 13 1 10 9 10 9 1 9 0 2 2
24 1 10 9 1 10 12 0 2 1 9 1 10 12 2 15 13 10 9 11 11 2 12 9 2
10 2 13 16 13 10 9 1 10 9 2
18 9 11 13 0 0 7 16 10 9 13 10 9 0 13 10 0 9 2
17 7 10 3 0 2 13 3 10 0 9 0 2 13 3 10 9 2
30 2 13 10 9 2 13 1 0 9 11 11 2 10 9 15 1 12 9 13 10 12 1 9 11 1 10 9 0 2 2
36 16 13 1 9 0 13 13 1 10 9 2 7 16 15 3 15 15 13 1 9 1 9 7 3 15 13 13 1 13 10 9 1 10 9 2 2
16 7 13 3 0 13 1 10 9 9 0 1 10 9 1 9 2
18 4 13 1 10 11 11 7 15 4 13 1 10 9 1 10 9 0 2
41 2 10 10 9 2 3 15 0 2 3 4 13 1 3 1 12 9 0 2 13 11 11 11 2 12 9 2 15 1 10 12 9 13 1 10 9 1 9 0 2 2
24 1 10 0 9 15 13 3 1 13 1 10 9 16 10 9 3 13 3 7 10 9 15 13 2
17 1 10 9 1 9 15 13 3 10 9 2 7 3 3 13 15 2
11 13 1 15 1 13 10 9 10 3 3 2
19 7 10 9 1 10 9 0 13 3 16 10 0 1 13 15 13 15 2 2
5 15 13 10 0 2
12 1 10 0 9 1 10 9 3 1 0 9 2
24 2 16 15 15 13 3 2 13 10 9 11 2 1 10 12 9 1 9 4 13 1 10 9 2
9 7 13 10 9 1 10 9 2 2
11 11 11 2 12 9 2 3 13 10 9 2
11 2 3 4 3 13 10 9 1 10 9 2
5 3 10 9 13 2
23 13 16 10 9 13 3 2 7 1 9 13 0 9 1 10 9 7 1 10 0 9 2 2
35 3 1 13 1 10 9 1 10 9 1 9 1 10 9 2 10 9 3 0 13 10 10 9 1 10 9 2 1 9 1 10 9 1 9 2
16 2 10 9 3 13 3 1 10 9 2 7 3 1 10 9 2
5 10 9 13 0 2
21 1 9 13 10 9 3 4 13 10 9 2 16 16 13 1 10 9 4 13 2 2
14 10 9 1 9 1 11 4 13 10 9 1 10 9 2
8 11 2 10 9 1 11 11 2
18 7 11 11 1 10 0 2 0 2 9 1 9 15 4 13 10 9 2
22 1 10 9 2 1 9 1 10 0 9 1 9 13 1 11 1 10 11 1 9 0 2
42 1 10 0 9 2 9 1 10 9 0 1 10 10 9 9 2 10 9 15 4 13 1 9 10 9 1 9 0 2 1 11 2 13 1 9 1 9 2 9 7 9 2
52 10 9 3 15 13 1 13 10 10 9 0 2 11 11 2 12 9 2 9 1 9 0 2 9 0 1 11 2 15 1 10 9 2 12 9 7 12 9 15 4 13 10 9 1 11 1 10 12 9 1 9 2
50 10 9 1 9 0 1 9 11 11 0 2 1 12 9 1 10 0 9 11 2 4 3 13 1 10 9 2 7 13 10 9 1 10 9 7 10 9 1 10 9 1 13 13 3 7 3 9 7 9 2
26 2 10 9 4 13 3 2 13 13 1 9 1 10 9 7 1 9 2 3 15 13 10 0 9 2 2
34 1 9 11 2 12 0 9 1 10 9 9 2 15 13 3 10 9 1 10 9 2 11 2 12 9 2 15 13 1 10 9 1 11 2
39 13 13 1 10 9 16 13 10 9 0 7 11 2 10 3 9 1 10 9 2 10 9 2 11 1 12 9 13 1 11 2 13 1 10 9 1 10 9 2
47 2 3 15 13 3 2 13 2 2 16 1 10 9 2 1 10 0 9 2 4 13 10 9 1 9 7 13 1 2 13 15 2 15 4 13 0 2 7 3 15 4 13 13 1 9 2 2
19 10 9 1 10 9 13 1 11 2 1 9 1 11 2 7 4 3 13 2
38 9 11 2 9 2 12 9 2 0 9 1 11 2 7 9 11 2 9 0 1 10 9 1 9 2 13 3 1 13 1 10 0 9 10 9 1 11 2
36 3 9 7 9 1 9 15 13 1 13 16 4 13 10 9 1 10 9 1 10 9 0 13 1 0 15 13 3 2 10 11 1 11 11 2 2
55 10 9 11 2 3 0 7 3 0 1 9 2 1 3 13 1 11 11 2 10 9 4 15 13 3 1 10 9 1 10 9 1 10 9 1 9 7 3 3 10 9 13 0 1 10 0 9 1 9 13 1 10 0 11 2
24 9 2 9 2 9 2 9 0 2 9 2 9 2 9 7 9 2 10 9 13 1 10 11 2
16 1 9 15 13 12 12 9 2 1 9 15 13 1 12 12 2
25 1 10 9 2 10 9 4 13 1 13 10 9 1 10 9 0 2 1 3 10 10 9 0 0 2
31 15 13 10 9 3 1 9 2 7 3 15 13 10 9 2 1 10 9 0 2 13 3 0 15 15 3 4 13 1 9 2
15 10 9 2 3 2 3 13 0 3 1 10 9 3 0 2
10 7 1 15 13 2 13 15 10 9 2
3 12 12 2
38 1 3 10 9 13 1 9 2 7 3 13 1 10 9 1 9 2 13 2 1 10 11 2 3 12 12 2 1 10 9 1 12 9 7 12 12 9 2
45 1 10 0 9 2 10 9 15 13 3 2 3 1 13 10 9 1 12 12 1 11 2 1 10 9 1 9 1 10 9 7 1 0 9 2 3 1 10 12 5 1 9 0 2 2
15 1 9 9 7 3 15 4 13 10 0 9 1 10 9 2
24 12 12 9 4 13 3 1 10 9 1 11 7 11 2 3 10 10 9 0 13 1 10 9 2
3 9 0 2
8 11 2 11 2 11 7 11 2
39 1 15 15 4 13 1 9 1 9 2 16 3 4 13 9 9 2 15 4 13 10 9 1 10 9 0 2 15 10 9 15 13 0 7 3 3 3 3 2
36 3 1 10 9 15 4 13 9 1 10 9 1 9 1 10 11 1 11 2 3 16 1 9 0 2 10 9 7 9 2 3 1 12 9 3 2
12 3 10 9 4 13 7 10 9 15 4 13 2
17 1 10 9 1 3 2 3 2 10 9 9 13 13 1 10 9 2
20 1 10 9 1 10 11 10 9 4 4 13 1 10 9 1 9 1 10 11 2
14 1 15 13 1 9 2 15 13 10 9 1 10 9 2
10 9 1 10 9 1 10 11 1 11 2
35 1 10 9 0 11 11 2 10 9 0 2 13 1 3 3 1 11 11 2 1 12 9 1 10 9 1 9 11 2 7 13 10 9 0 2
50 0 13 16 10 9 1 10 10 9 13 10 9 2 15 10 11 10 9 4 13 1 13 1 10 9 1 10 0 9 13 1 10 9 0 7 1 10 9 1 10 10 9 1 9 2 10 9 11 11 2
33 11 2 13 1 9 2 4 13 10 0 9 10 9 1 11 1 10 0 9 1 10 9 2 1 10 12 9 13 1 11 1 11 2
43 1 10 9 0 10 11 13 3 1 10 12 9 2 10 9 3 13 10 9 1 10 9 0 2 1 3 13 11 2 3 10 12 4 13 1 10 9 1 11 1 10 11 2
17 1 10 9 0 2 3 2 10 9 3 0 1 10 9 1 9 2
41 10 9 1 11 11 2 1 15 3 0 9 1 10 9 0 1 9 2 7 3 4 13 1 9 2 11 11 2 3 1 10 9 11 2 15 1 3 13 12 9 2
30 11 2 3 2 4 13 1 10 9 1 13 15 13 1 9 7 9 2 15 4 13 9 1 10 9 3 0 1 11 2
27 3 9 10 0 9 15 4 13 1 10 10 9 7 1 10 9 10 9 4 13 1 9 7 1 9 0 2
22 3 10 0 9 0 3 4 13 10 9 0 2 15 3 1 9 4 13 1 9 11 2
14 13 3 3 12 10 9 15 4 13 10 9 1 11 2
28 1 10 9 0 2 3 2 10 9 1 11 15 4 13 12 9 1 9 1 10 12 9 1 9 13 1 11 2
24 9 9 10 9 4 13 10 9 1 11 2 12 12 2 7 3 4 4 13 0 1 10 9 2
22 9 3 13 11 7 11 2 3 1 9 1 10 9 1 10 9 11 1 10 0 9 2
23 3 13 10 9 1 10 12 9 7 11 1 9 1 10 0 13 1 10 0 9 1 9 2
31 1 15 13 10 9 13 1 11 2 10 9 11 13 1 13 10 9 2 11 7 11 10 9 3 13 2 1 13 10 9 2
10 13 1 10 9 15 13 1 10 9 2
3 9 11 2
6 0 9 1 9 11 2
18 12 9 4 13 1 9 2 1 9 1 9 3 0 2 10 0 9 2
27 10 9 15 4 13 16 13 9 16 15 13 1 13 9 1 10 9 1 10 9 7 15 4 13 13 15 2
34 11 11 2 12 9 2 4 4 13 1 10 9 1 10 0 9 1 10 11 2 1 10 11 11 2 15 15 4 13 0 1 12 9 2
8 1 10 9 4 13 10 9 2
5 4 13 9 9 2
40 11 11 4 13 16 4 13 1 13 15 13 15 1 10 9 1 10 9 1 11 11 1 10 11 2 16 4 13 10 9 1 9 15 13 7 13 1 9 0 2
28 2 15 4 13 1 10 9 1 3 15 13 15 2 4 13 10 9 2 7 13 0 1 13 15 1 0 2 2
12 3 11 4 13 1 13 15 1 13 3 9 2
11 2 13 15 13 2 13 3 1 3 2 2
47 3 3 2 12 1 10 9 2 15 0 7 10 15 0 1 10 9 1 10 9 2 15 4 13 1 10 9 15 13 1 4 13 2 4 13 10 9 1 9 7 15 4 13 1 10 9 2
20 3 4 13 10 10 9 2 15 3 15 4 13 1 10 9 2 7 4 13 2
11 12 9 3 10 9 2 3 11 1 11 2
3 9 11 2
12 3 13 10 0 9 1 10 9 1 11 11 2
20 1 10 9 10 9 13 13 10 11 7 10 9 1 10 9 4 13 3 0 2
44 10 9 1 10 9 13 10 12 9 1 10 12 1 12 9 1 9 1 9 11 3 13 10 9 7 3 1 10 9 1 15 3 0 4 4 13 10 9 3 4 13 10 11 2
38 3 3 10 9 11 11 2 9 1 10 0 11 2 13 10 9 3 1 10 11 1 10 9 1 4 13 11 2 9 2 4 13 1 13 1 10 9 2
47 2 10 9 4 4 13 1 10 0 9 2 3 0 2 16 3 15 4 13 10 9 0 7 3 15 15 4 13 1 9 2 1 15 15 13 10 9 11 1 10 9 1 10 9 0 2 2
34 11 2 1 9 1 15 1 10 9 1 10 9 2 11 11 2 4 13 16 2 10 9 4 13 2 13 0 15 15 4 4 13 2 2
16 2 4 13 1 10 9 15 13 1 10 9 1 9 3 0 2
23 9 15 3 3 15 4 3 13 1 13 15 1 9 7 1 13 1 10 10 9 10 9 2
20 10 9 13 9 1 13 15 9 7 3 15 4 13 3 10 9 1 9 2 2
13 9 1 9 7 9 1 10 9 1 10 9 9 2
3 11 11 2
23 12 10 9 13 1 10 9 16 13 0 1 13 1 9 15 13 9 1 10 9 1 9 2
17 3 1 15 2 4 4 13 10 12 9 15 13 10 9 1 9 2
12 12 9 1 9 3 1 10 9 1 10 9 2
23 10 9 11 4 1 9 13 3 10 9 1 9 1 10 9 1 9 7 1 10 9 0 2
16 12 9 1 10 9 3 0 7 15 13 9 1 10 0 9 2
16 10 9 1 9 4 13 10 9 1 9 7 9 2 3 0 2
28 7 3 16 4 13 1 9 11 11 11 2 12 9 2 0 2 13 16 13 10 9 1 9 1 10 0 9 2
17 13 9 7 9 16 10 9 1 10 9 4 4 13 1 10 11 2
21 10 9 0 2 7 1 9 1 10 9 1 9 2 15 4 13 1 10 9 11 2
19 7 1 10 9 10 9 2 11 2 12 9 2 4 4 13 1 9 0 2
18 13 10 11 1 9 0 7 10 10 9 15 13 0 1 10 9 0 2
18 9 1 9 2 11 11 2 0 1 12 9 2 13 15 13 10 9 2
8 2 3 13 1 10 11 2 2
15 1 9 7 9 2 9 7 9 1 9 1 13 10 9 2
17 13 10 9 1 11 11 2 1 10 11 2 2 10 0 9 0 2
16 10 9 0 2 13 2 15 3 13 9 16 3 15 4 13 2
11 3 13 3 10 9 1 15 3 13 9 2
36 10 9 3 4 13 1 10 9 1 10 3 0 7 0 9 0 1 10 9 15 15 13 1 13 1 10 9 1 9 10 10 12 9 1 9 2
10 11 11 13 12 9 7 15 13 3 2
22 7 16 13 10 9 0 1 9 0 2 10 9 7 10 9 0 13 0 1 10 9 2
24 9 1 10 9 1 11 2 13 1 10 9 1 9 1 9 7 1 9 1 10 9 1 9 2
12 13 10 9 1 10 9 1 3 1 12 9 2
10 10 0 1 9 3 15 4 13 0 2
12 10 9 15 13 1 10 9 1 10 9 0 2
5 4 13 1 15 2
22 10 10 9 1 9 13 1 10 9 1 11 11 1 10 12 1 10 12 1 10 9 2
14 10 9 1 9 1 11 11 13 10 9 1 10 9 2
16 15 13 9 2 15 13 9 1 10 9 2 10 9 3 13 2
26 2 3 13 0 13 3 1 13 1 15 7 3 1 13 10 9 2 13 1 15 2 2 13 11 2 2
32 1 10 9 1 10 11 1 9 2 1 10 9 1 9 0 2 4 13 13 9 3 0 16 10 9 13 1 10 10 9 2 2
20 10 9 13 0 1 9 1 10 12 7 10 12 9 2 1 9 7 1 9 2
22 10 0 12 9 2 1 9 1 10 2 11 2 2 13 9 1 4 15 13 1 9 2
11 10 12 9 0 13 0 1 10 10 9 2
20 10 0 12 9 13 0 2 7 3 16 13 9 7 3 15 13 9 1 13 2
9 2 10 9 2 6 6 10 9 2
29 13 1 13 10 2 9 2 15 3 13 10 12 9 1 9 2 7 4 13 3 0 2 2 2 13 10 0 9 2
56 2 6 2 3 16 15 13 10 0 7 3 13 1 9 1 10 9 1 9 1 10 9 2 1 9 7 12 9 1 10 9 1 10 9 2 13 1 13 15 13 1 9 16 3 1 10 9 4 4 13 1 9 1 10 9 2
26 3 2 15 13 1 13 2 13 10 9 0 16 1 15 13 1 9 1 13 10 9 3 1 10 9 2
19 3 1 10 9 3 10 9 1 10 9 3 0 4 13 10 2 11 2 2
39 10 9 1 9 1 9 1 10 15 10 9 2 13 1 9 2 4 13 15 1 13 1 9 10 9 13 0 2 1 13 15 10 9 0 1 9 1 9 2
20 9 1 9 7 9 0 7 10 0 9 1 9 13 3 1 9 1 10 9 2
17 1 9 2 0 1 10 0 9 15 13 3 9 2 9 7 9 2
8 10 9 4 13 1 10 9 2
16 2 13 1 9 1 10 0 9 16 13 3 0 13 10 9 2
16 1 9 15 13 3 10 9 1 10 9 2 2 13 11 2 2
27 1 9 1 10 9 1 9 7 1 9 2 9 2 9 2 9 0 2 13 1 9 1 10 9 0 2 2
33 2 15 13 9 1 9 1 13 3 10 9 1 10 11 1 11 7 10 9 1 10 9 1 10 11 1 10 11 15 3 13 3 2
18 15 1 15 15 4 13 10 9 1 13 15 13 10 9 1 10 9 2
8 15 13 3 15 13 10 9 2
23 13 1 13 10 12 9 15 15 13 0 2 16 10 9 13 1 13 1 9 0 10 9 2
16 16 15 13 4 13 10 9 0 1 13 15 1 10 9 2 2
9 2 7 15 13 3 9 3 0 2
26 1 9 2 16 10 9 1 10 11 13 0 15 4 13 13 7 15 4 13 2 13 2 13 1 9 2
22 15 13 10 9 7 13 1 11 2 10 10 9 2 15 13 10 9 0 1 11 2 2
19 2 10 9 1 9 1 10 9 7 1 10 9 1 10 9 13 0 9 2
13 10 11 11 15 13 3 2 3 1 10 9 2 2
11 10 9 10 9 13 13 1 0 7 0 2
28 13 10 9 1 13 10 9 1 10 9 2 1 9 1 0 9 0 0 0 15 1 13 1 9 0 7 0 2
49 3 9 7 9 13 13 2 1 9 1 10 0 7 0 9 15 1 9 4 13 10 9 1 10 2 9 2 1 10 9 2 16 13 10 9 1 10 9 1 10 9 11 1 10 9 1 10 9 2
3 10 9 2
47 10 11 1 10 11 11 4 13 1 10 12 2 1 10 9 1 10 0 9 0 1 10 11 0 7 13 10 10 9 3 0 1 9 1 10 9 1 9 1 10 9 1 11 1 10 12 2
19 12 9 2 9 2 13 1 10 12 1 10 9 1 10 9 11 11 11 2
26 10 10 9 13 2 1 10 13 9 7 9 1 10 9 0 1 10 11 11 7 1 10 10 9 2 2
13 4 13 3 1 12 9 7 10 9 0 1 12 2
15 10 9 0 4 13 1 10 9 0 1 10 0 9 0 2
5 1 9 1 11 2
10 11 2 3 13 2 10 0 11 2 2
19 10 9 0 1 10 9 0 2 9 1 10 9 2 10 9 2 10 9 2
25 10 10 9 7 10 10 9 2 13 1 10 0 9 1 10 9 0 2 4 13 10 9 1 9 2
27 1 9 12 2 1 10 9 2 10 9 1 9 2 0 13 15 3 15 1 10 10 9 11 0 1 13 2
8 1 9 12 2 10 0 9 2
8 1 10 9 10 9 1 9 2
17 1 10 9 3 2 10 9 1 10 9 2 12 9 2 10 9 2
22 1 10 9 10 9 15 3 4 13 3 10 0 2 0 2 0 9 1 10 9 11 2
14 1 10 9 2 12 0 9 1 9 1 9 1 9 2
10 1 10 15 13 13 10 9 1 9 2
23 1 9 2 9 7 9 3 0 0 11 2 3 10 9 11 13 3 1 13 10 0 9 2
14 1 10 9 0 2 0 9 1 9 1 9 1 9 2
31 10 10 9 1 11 11 15 13 10 9 4 13 1 10 0 9 2 11 2 1 11 11 2 3 13 1 11 1 11 11 2
8 10 9 13 13 1 9 0 2
5 9 1 11 11 2
11 9 11 11 5 11 11 11 2 11 11 2
30 10 9 1 10 9 0 2 15 4 4 13 1 11 2 7 3 13 2 1 13 0 1 11 11 2 13 1 10 9 2
37 10 9 1 9 0 9 2 1 15 13 13 15 10 9 1 11 2 7 1 10 15 10 0 9 4 13 13 12 9 1 9 2 2 13 1 9 2
21 10 9 13 10 9 3 1 10 9 1 10 0 9 1 10 11 0 1 10 11 2
21 3 0 1 10 9 15 3 13 1 10 9 2 1 13 10 9 15 15 4 13 2
13 15 13 1 10 9 1 9 2 0 1 10 9 2
30 11 11 2 9 7 9 0 1 9 0 2 9 1 10 9 2 15 13 16 10 9 13 10 9 1 9 7 1 9 2
20 1 10 9 4 13 3 10 9 0 2 1 10 9 2 1 0 9 1 9 2
28 13 15 10 9 1 9 2 0 13 1 0 9 1 9 2 15 13 1 10 9 13 1 10 9 1 10 9 2
13 11 13 16 3 13 10 2 9 2 1 10 9 2
26 10 9 1 13 13 13 1 10 9 10 2 9 0 2 0 2 2 1 10 9 2 0 2 0 2 2
23 1 9 0 2 15 13 1 10 9 0 2 15 13 10 9 2 3 0 1 10 0 9 2
21 7 10 0 9 0 4 13 1 10 0 9 1 10 9 15 13 1 10 0 9 2
3 10 9 2
11 10 9 13 10 9 1 10 9 9 11 2
39 15 13 1 10 9 7 1 10 9 9 1 9 1 9 2 13 1 10 9 0 1 10 11 1 11 2 7 15 13 10 9 13 1 10 9 1 10 12 2
29 10 9 2 0 1 13 10 9 1 9 2 3 15 13 1 10 9 1 13 15 7 13 9 0 1 10 9 0 2
10 10 9 13 10 9 1 10 9 11 2
17 3 10 12 9 13 1 10 9 2 1 13 10 9 1 10 9 2
38 1 10 9 0 2 2 10 9 1 11 2 7 15 13 1 11 7 10 0 9 0 2 3 13 1 11 2 3 15 13 2 10 9 1 9 0 2 2
28 1 3 10 9 1 9 2 1 10 9 0 1 10 9 2 11 15 4 13 1 13 10 9 0 1 10 11 2
15 13 3 0 13 12 9 1 10 9 1 10 2 9 2 2
42 1 13 1 10 12 2 15 13 1 12 9 1 11 1 10 9 0 15 13 1 9 10 9 0 0 1 10 9 12 2 12 2 1 10 11 1 11 1 10 9 2 2
29 15 13 1 10 9 0 2 13 1 10 11 11 2 13 1 11 2 13 1 10 0 9 0 1 10 9 1 11 2
17 10 9 0 7 0 1 10 9 2 1 10 9 2 1 10 9 2
21 10 11 0 15 13 10 9 0 7 15 15 4 3 13 1 10 10 10 9 0 2
6 10 9 15 13 11 2
3 3 13 2
25 13 10 9 1 10 0 0 9 2 15 13 10 0 9 2 1 0 9 2 15 3 13 1 13 2
22 10 9 13 1 13 2 10 9 13 10 9 1 10 9 7 13 3 3 10 9 0 2
57 10 9 13 1 0 9 7 13 10 9 1 10 9 1 10 9 1 10 9 2 7 1 0 9 1 10 9 0 2 10 9 13 3 0 2 15 13 1 3 2 3 1 13 2 1 10 0 9 1 9 2 3 10 0 9 0 2
31 10 9 13 9 1 10 9 3 0 7 0 7 4 13 1 10 9 2 1 10 15 3 15 13 10 9 0 1 10 9 2
22 10 9 10 9 1 12 9 13 3 0 7 15 1 10 10 9 4 13 1 10 9 2
26 10 9 2 1 10 9 1 10 0 9 2 10 9 13 10 9 2 13 15 7 13 1 10 9 0 2
31 10 9 13 13 16 15 13 10 0 9 0 2 13 1 9 1 9 1 9 13 7 10 0 9 2 15 13 10 0 9 2
15 1 10 9 2 10 9 13 13 7 4 13 1 10 0 2
29 15 13 13 10 9 1 10 9 7 2 13 10 9 1 10 9 2 15 15 13 1 13 10 9 1 13 15 3 2
10 7 3 10 9 0 2 1 9 0 2
14 3 10 2 9 2 2 1 10 9 7 10 9 13 2
22 1 10 9 11 13 10 0 9 1 10 9 0 2 7 3 13 1 9 7 9 0 2
19 3 2 1 10 9 1 9 2 10 9 13 1 9 7 3 1 9 0 2
13 10 9 1 10 9 7 1 10 9 13 3 0 2
21 7 13 3 13 15 3 9 1 9 3 13 1 9 2 16 10 9 15 13 3 2
32 10 0 9 3 0 13 10 9 2 15 2 13 15 2 13 10 9 13 1 10 9 1 10 9 7 2 10 9 2 10 9 2
23 0 13 10 9 1 9 2 1 9 0 7 0 2 1 4 3 13 7 13 10 0 9 2
16 1 0 2 10 10 9 13 3 0 7 13 1 9 7 9 2
43 1 10 9 15 13 2 1 10 9 0 1 10 9 0 2 9 7 9 2 1 9 2 15 13 1 9 1 10 0 9 1 10 9 2 2 15 1 10 0 9 1 9 2
8 9 2 9 2 9 1 11 2
10 7 1 11 3 9 2 9 2 9 2
20 3 4 13 16 10 9 11 3 13 10 9 1 9 2 1 9 1 10 9 2
17 3 3 13 3 10 9 1 10 11 7 10 9 1 10 11 11 2
17 1 10 9 15 13 1 9 2 1 10 9 2 10 0 9 0 2
22 10 9 10 9 15 13 3 0 2 3 1 10 0 9 2 1 9 2 1 10 9 2
22 10 9 3 0 2 1 15 13 9 10 9 1 0 2 3 13 3 1 10 0 9 2
13 0 13 10 9 1 10 9 2 1 10 9 11 2
12 1 10 9 2 3 1 10 9 13 10 9 2
27 10 9 0 13 0 7 0 13 10 0 9 2 15 13 2 1 10 9 2 1 13 10 9 1 10 9 2
32 16 3 15 13 9 0 2 1 9 1 9 2 13 9 15 15 13 1 10 9 1 10 0 2 1 10 0 9 1 9 0 2
31 7 10 9 3 13 16 10 9 13 0 7 3 13 2 16 10 9 1 9 13 13 1 9 7 16 10 9 13 10 9 2
29 7 15 1 10 9 13 3 10 0 9 1 10 9 2 15 13 13 1 10 0 9 1 10 10 9 1 10 9 2
29 1 10 9 1 9 0 2 1 11 2 10 0 9 13 13 1 10 9 1 9 11 3 15 4 13 10 10 9 2
31 13 3 16 13 0 13 2 1 10 9 0 2 10 0 0 9 2 13 1 10 9 2 1 9 1 9 13 1 0 9 2
73 7 2 1 10 9 1 9 1 9 7 9 2 3 4 13 10 9 1 9 1 9 2 2 10 9 1 9 2 10 9 1 9 13 2 10 9 13 2 1 9 0 1 10 9 2 13 1 13 13 10 9 13 1 10 9 1 11 2 1 11 2 1 11 11 2 7 13 15 10 10 9 0 2
22 10 9 1 9 2 13 3 1 9 2 7 3 1 10 9 1 10 9 7 10 9 2
20 10 11 3 13 3 10 9 2 7 3 10 9 1 9 13 1 9 7 9 2
35 10 0 9 1 10 11 13 10 15 15 13 1 10 9 1 10 12 2 16 11 4 13 2 1 10 11 0 2 1 10 9 1 10 11 2
52 15 13 10 9 2 0 2 1 10 10 9 2 1 13 1 9 2 13 10 9 0 2 10 9 0 2 10 0 9 2 10 0 9 1 10 9 2 0 2 15 4 13 15 3 2 1 10 9 1 10 9 2
32 9 7 9 3 3 0 15 13 1 10 9 0 2 1 10 9 0 2 1 10 9 1 9 2 1 10 0 9 1 9 0 2
25 3 2 1 10 9 1 9 2 3 16 9 7 9 15 13 3 9 0 7 2 3 2 9 0 2
18 13 10 11 2 3 13 1 9 2 10 9 2 2 3 10 9 0 2
27 1 9 2 3 2 1 10 0 9 1 10 9 15 4 13 15 2 3 1 10 9 1 11 1 10 9 2
34 13 3 16 2 3 1 10 9 1 9 0 2 1 10 10 0 9 1 9 7 3 1 9 2 13 3 10 9 1 10 0 9 11 2
21 16 13 10 9 1 10 9 11 2 13 1 4 13 10 0 9 1 10 10 9 2
25 7 13 3 16 13 10 10 0 9 1 10 9 1 10 0 9 2 13 15 1 9 1 11 0 2
9 0 9 4 13 1 10 9 0 2
29 3 10 9 4 13 1 9 2 1 10 9 15 13 10 9 2 7 13 9 1 9 2 9 1 10 0 9 0 2
33 1 10 9 0 7 0 2 13 9 1 15 10 9 1 9 3 13 2 1 15 10 9 1 9 13 13 3 9 2 1 9 2 2
20 4 4 13 9 1 10 9 1 9 0 2 1 15 10 9 4 13 0 9 2
19 15 13 9 1 10 9 1 10 9 1 9 1 9 2 7 1 10 9 2
30 4 13 10 9 13 1 9 1 15 15 13 1 10 9 10 0 9 11 11 2 3 13 3 1 10 11 16 0 2 2
9 10 9 13 3 13 1 10 9 2
25 15 4 13 16 4 13 2 1 0 9 2 1 9 0 15 13 1 10 9 2 9 1 9 0 2
22 7 3 15 13 16 13 10 9 2 10 9 1 10 9 9 7 1 10 9 1 9 2
19 7 3 2 1 10 0 9 2 15 13 1 10 9 0 2 1 10 9 2
12 1 10 9 0 1 11 1 10 9 1 11 2
74 7 16 15 13 1 10 0 9 2 3 4 4 13 10 9 1 10 12 7 10 9 15 15 13 9 7 9 2 15 13 3 10 10 9 0 1 11 2 15 1 9 2 1 10 15 2 3 13 3 10 9 1 9 2 7 1 10 10 0 9 13 4 13 3 12 9 1 11 2 11 7 11 2 2
31 7 10 9 3 0 13 10 2 8 2 8 2 8 2 2 1 15 2 1 0 9 2 15 4 13 10 9 0 1 11 2
16 3 1 13 10 9 1 3 16 3 3 10 9 13 0 0 2
17 1 9 1 11 10 9 0 1 10 9 0 10 9 10 9 10 9
28 10 0 9 1 10 9 1 10 9 13 10 9 7 10 9 0 2 7 3 15 13 10 0 9 1 10 9 2
8 0 2 0 2 0 1 13 2
5 0 1 10 9 2
23 3 1 0 9 0 1 9 2 1 15 1 11 2 13 0 9 2 3 3 0 7 0 2
25 2 11 2 2 1 11 2 13 10 9 1 9 0 2 9 12 2 1 0 9 2 12 9 2 2
22 9 1 10 9 0 10 9 13 10 9 0 2 13 1 9 13 1 10 9 1 9 2
19 13 1 9 2 13 1 9 12 1 9 12 10 9 1 10 9 1 9 2
8 10 9 1 11 13 1 11 2
27 10 0 9 1 10 9 0 2 2 11 2 13 3 0 1 9 1 9 0 13 1 9 1 10 0 9 2
6 10 9 13 9 12 2
12 13 1 11 11 2 13 3 9 12 10 9 2
24 10 9 7 10 9 1 9 2 1 11 11 2 13 1 9 1 11 2 1 10 9 1 9 2
2 12 2
9 12 9 2 9 12 7 9 12 2
11 1 10 12 1 10 12 9 1 10 9 2
2 12 2
24 2 11 13 2 2 9 13 13 1 9 7 13 3 2 1 10 9 2 11 2 1 11 11 2
13 10 9 2 11 2 13 1 9 9 1 9 0 2
11 9 1 9 12 2 12 2 12 2 12 2
2 12 2
2 12 2
16 3 1 11 11 3 2 11 2 2 1 9 1 9 1 9 2
19 10 12 9 3 0 13 3 9 1 2 11 2 2 13 1 9 7 9 2
2 12 2
26 2 11 2 2 1 11 2 1 10 9 2 11 1 11 2 2 2 11 11 2 7 2 11 11 2 2
10 9 1 10 12 1 10 12 10 9 2
2 12 2
2 12 2
21 1 11 9 1 9 0 2 9 2 11 2 2 1 9 12 1 9 12 10 9 2
12 9 1 9 0 2 13 1 9 1 0 9 2
13 1 11 2 13 1 9 12 1 9 12 10 9 2
2 12 2
24 2 11 2 2 0 7 0 2 7 2 11 11 2 2 0 9 1 11 2 13 1 11 11 2
10 9 12 2 9 12 7 12 10 9 2
2 12 2
14 9 13 7 13 1 9 1 11 11 2 9 11 2 2
12 10 9 1 9 13 3 9 12 13 10 9 2
2 12 2
16 1 11 11 2 9 13 1 9 1 9 0 9 2 11 2 2
18 9 12 10 9 2 1 0 2 7 9 12 10 9 2 1 0 2 2
18 2 11 2 7 2 11 2 2 1 9 0 2 13 9 12 10 9 2
2 12 2
15 11 11 1 11 2 9 11 2 13 1 12 9 1 9 2
18 9 1 9 0 0 7 0 2 13 1 9 12 1 9 12 10 9 2
2 12 2
20 1 11 11 2 9 11 2 9 1 0 9 2 12 9 2 2 13 1 9 2
5 9 12 10 9 2
5 9 1 11 11 2
5 9 1 11 11 2
44 1 10 0 9 1 11 2 13 1 9 1 9 2 9 7 11 2 4 13 1 13 0 9 3 1 9 1 9 2 10 9 0 2 15 3 4 13 1 10 9 1 10 9 2
8 13 10 9 1 10 9 0 2
32 10 9 3 13 3 1 10 9 13 2 3 1 10 9 1 10 9 7 1 10 9 16 10 9 0 3 13 9 1 9 0 2
14 10 9 2 3 2 13 10 0 9 7 13 3 0 2
19 3 3 1 10 0 9 0 1 9 2 7 1 9 2 16 13 3 3 2
41 10 0 0 9 2 15 13 1 13 10 9 1 9 16 4 13 1 9 0 1 15 13 1 10 9 2 0 2 2 1 10 9 2 13 10 0 9 1 10 9 2
70 10 9 2 13 1 9 1 10 9 1 10 9 0 11 2 13 2 1 9 0 2 1 13 1 10 9 9 0 2 12 9 2 7 1 0 9 2 1 13 7 13 10 9 2 13 15 3 1 10 0 9 1 9 1 9 15 15 13 1 13 15 10 9 2 13 10 11 11 2 2
21 13 0 3 13 9 15 13 9 0 1 10 9 13 1 10 9 7 1 10 9 2
8 3 1 9 12 7 9 12 2
27 15 13 9 3 0 16 10 0 9 13 10 9 1 10 9 3 0 1 4 13 2 13 7 13 1 9 2
5 7 3 13 15 2
61 1 0 9 1 9 2 10 11 13 9 1 0 9 13 9 2 0 2 1 15 3 2 13 10 10 9 1 9 2 13 10 9 1 9 7 9 0 2 13 1 10 9 0 0 9 2 1 10 9 13 7 10 9 1 10 9 2 9 11 2 2
24 13 9 1 0 9 2 1 0 9 2 1 9 7 9 13 1 12 15 3 1 10 9 0 2
60 10 9 1 9 7 15 1 9 1 9 2 13 2 3 2 1 9 0 2 10 9 0 1 10 9 2 13 0 2 3 1 0 9 2 3 10 9 0 7 0 2 15 15 2 3 2 13 3 0 7 0 1 9 1 10 3 0 9 0 2
17 3 1 10 9 1 9 13 3 0 13 1 10 2 0 9 2 2
24 10 9 1 10 9 13 3 0 1 10 9 2 3 1 15 1 15 3 1 3 4 13 0 2
27 9 7 0 9 13 2 13 3 9 2 0 9 1 9 2 3 1 0 9 7 1 0 9 1 10 9 2
18 3 3 4 3 13 10 9 1 10 9 7 3 15 1 10 0 9 2
47 16 4 13 10 9 1 13 9 1 9 2 10 11 4 13 3 10 9 1 13 15 1 0 9 1 9 1 13 15 0 3 1 10 9 0 2 1 10 9 0 2 1 9 7 1 9 2
9 7 1 15 13 1 10 0 9 2
16 10 11 11 2 3 2 15 13 9 13 1 10 9 1 9 2
35 10 0 9 13 13 7 13 2 13 10 9 1 12 9 2 7 10 9 13 1 9 1 9 2 7 1 9 16 10 9 0 13 3 0 2
31 3 1 10 9 2 13 1 10 0 9 1 10 9 2 15 4 13 9 0 7 13 3 9 2 9 0 2 9 7 9 2
19 10 9 0 3 0 13 1 13 9 7 9 0 7 1 9 1 10 9 2
30 13 1 9 2 13 1 10 0 9 2 13 1 9 13 13 1 9 9 2 12 2 12 1 12 2 7 3 13 3 2
55 15 13 1 10 2 11 2 2 13 1 11 11 2 15 2 3 1 9 15 13 15 1 10 9 2 3 1 9 1 9 2 2 13 9 0 0 2 1 10 9 2 10 9 2 10 9 0 2 10 9 7 9 3 0 2
16 1 10 9 1 10 9 2 4 13 1 9 9 1 10 9 2
52 10 9 4 3 13 9 1 10 9 1 0 9 1 10 9 7 1 10 9 2 7 3 2 7 15 13 10 9 1 9 2 1 10 9 1 9 0 2 1 9 2 1 9 1 9 2 1 9 1 0 9 2
27 13 0 3 1 10 9 16 10 9 0 2 9 12 2 12 2 12 2 12 2 13 10 9 1 0 9 2
5 0 3 10 9 2
12 1 10 0 9 12 3 1 10 0 9 12 2
37 1 10 9 1 10 9 2 10 9 2 0 2 7 0 1 9 15 2 0 2 4 13 0 9 1 10 11 7 1 10 0 9 1 10 10 9 2
40 10 10 9 0 13 3 0 7 15 13 10 9 1 13 9 1 10 9 2 7 4 13 10 9 1 3 13 15 10 9 2 13 16 13 0 13 15 1 9 2
20 9 0 1 10 9 2 9 0 7 9 0 2 1 9 0 2 0 2 0 2
22 3 15 1 15 13 3 2 1 10 0 9 2 10 0 9 15 13 10 9 1 13 2
7 13 10 9 0 7 0 2
21 3 15 13 3 15 13 9 1 9 1 10 0 9 7 10 0 9 1 10 9 2
21 13 10 11 1 11 15 13 1 9 3 12 9 2 13 1 0 9 1 10 9 2
38 10 9 4 13 1 9 2 15 1 15 2 13 9 0 3 4 13 10 9 0 1 9 0 13 1 15 15 13 10 9 2 9 7 9 1 9 2 2
13 15 13 2 15 13 1 10 0 9 7 15 13 2
21 1 13 10 9 2 10 0 9 1 9 4 13 2 9 1 9 2 1 10 9 2
24 3 1 10 0 2 7 0 2 9 15 4 13 9 0 7 9 2 1 13 9 7 9 9 2
35 15 13 1 9 1 9 7 9 7 15 13 1 9 7 9 1 11 2 13 15 3 3 0 1 9 1 13 3 9 16 13 1 10 9 2
16 7 3 15 1 10 9 2 10 9 3 3 13 1 10 9 2
18 13 1 9 1 9 13 1 9 2 1 9 0 7 0 7 0 9 2
37 10 9 1 9 1 10 9 13 3 10 9 2 1 10 15 4 13 10 9 1 9 0 3 4 3 13 10 9 1 9 0 1 9 1 9 0 2
7 15 13 3 1 10 9 2
56 3 2 10 9 1 9 4 3 4 13 1 9 0 2 0 12 7 12 9 7 2 1 13 10 9 7 13 10 9 1 0 9 2 0 9 1 10 9 0 15 13 1 9 13 1 9 7 3 0 2 7 1 9 0 2 2
23 10 9 0 13 3 10 9 13 1 9 2 1 10 9 2 7 10 9 13 3 10 15 2
12 9 9 2 9 9 2 9 2 9 2 9 2
14 9 0 2 0 15 13 7 15 13 1 10 9 0 2
38 15 15 13 3 0 1 10 9 1 10 9 4 13 1 10 9 1 2 13 2 10 9 2 3 13 10 9 0 2 7 13 10 3 0 9 1 9 2
15 10 9 13 1 10 9 0 7 1 9 3 1 15 0 2
18 3 1 10 9 0 7 1 10 9 15 13 9 1 9 13 1 9 2
23 1 10 9 0 10 9 13 3 0 2 16 10 9 2 16 13 0 2 3 13 1 9 2
7 1 9 15 13 10 9 2
21 13 15 10 9 15 13 1 10 9 2 9 2 0 13 1 10 9 1 10 9 2
33 3 1 10 10 9 0 10 9 13 1 9 2 1 9 13 1 9 2 1 10 11 11 1 11 15 13 1 10 9 0 1 9 2
28 15 13 1 10 9 3 10 9 1 10 9 2 11 11 2 1 11 1 10 11 2 13 1 11 1 11 2 2
30 13 7 13 3 1 9 2 10 9 13 1 10 9 1 9 2 1 10 9 0 2 1 10 9 0 2 10 10 9 2
27 0 2 0 2 0 2 0 2 1 9 2 1 9 2 1 9 2 10 9 13 9 0 2 1 10 9 2
38 3 10 11 11 13 1 10 9 1 9 10 9 0 15 13 1 9 9 13 1 10 9 0 2 1 9 0 2 3 1 9 0 2 7 0 1 9 2
27 3 15 4 13 10 9 0 1 9 13 1 9 0 1 9 0 2 3 4 3 13 10 9 1 10 9 2
18 0 10 9 1 9 7 1 9 1 0 7 0 1 13 1 9 0 2
39 1 10 9 1 10 9 4 4 13 10 0 7 0 9 3 10 2 9 2 9 13 10 9 0 1 9 15 2 1 10 9 2 4 13 1 10 10 9 2
22 1 13 10 10 9 13 10 9 1 9 15 1 10 10 9 15 13 1 10 0 9 2
30 15 13 2 11 11 2 2 13 1 11 7 13 1 11 1 11 2 7 13 1 10 0 9 1 9 0 13 1 9 2
30 4 4 13 7 13 2 3 3 9 7 2 1 10 10 0 9 2 4 13 1 10 9 7 3 1 15 1 0 9 2
18 12 9 1 13 15 2 12 9 1 13 15 2 12 9 1 13 15 2
3 9 9 2
31 13 10 9 1 10 9 1 13 10 9 0 2 10 9 13 13 1 9 15 12 9 9 15 15 13 10 9 1 0 9 2
12 3 3 2 3 2 3 2 1 9 1 9 2
3 9 0 2
2 9 2
3 9 13 2
5 9 1 10 9 2
2 9 2
17 7 3 3 15 13 10 9 1 3 13 7 15 15 13 10 9 2
14 1 13 1 10 9 2 3 15 13 1 10 9 0 2
8 0 1 13 7 3 1 13 2
13 7 1 10 0 9 2 10 0 9 3 15 13 2
3 15 13 2
17 1 0 9 2 12 9 1 10 9 2 13 10 9 1 15 0 2
8 13 12 9 1 13 15 3 2
6 7 4 13 9 0 2
2 3 2
17 16 13 16 10 0 9 13 3 0 13 1 9 10 9 7 13 2
10 10 9 1 9 7 10 9 1 9 2
15 10 9 13 10 9 1 10 9 1 9 2 9 2 9 2
16 13 3 0 13 3 1 10 9 1 10 9 1 10 9 0 2
20 13 3 3 13 10 9 1 9 0 15 13 1 9 1 9 0 7 9 0 2
2 3 2
13 3 2 7 3 16 1 10 9 0 7 3 13 2
29 13 3 2 3 16 10 9 13 13 1 10 9 1 10 9 7 10 9 2 1 10 9 3 2 15 15 13 2 2
2 3 2
13 1 10 9 0 15 13 3 12 9 1 9 9 2
9 3 10 9 1 13 7 13 3 2
2 11 2
16 15 13 3 3 15 16 10 9 0 13 9 1 10 9 13 2
14 13 1 13 15 13 15 1 10 0 9 1 10 9 2
10 10 9 13 0 7 15 4 13 3 2
17 13 10 9 0 2 3 2 13 1 13 3 16 13 10 9 0 2
7 10 9 4 13 12 9 2
3 9 0 2
8 13 1 13 3 1 10 9 2
15 13 1 13 10 9 7 13 16 10 9 15 13 1 9 2
14 16 15 13 15 0 3 13 15 7 13 1 13 15 2
11 13 3 7 13 3 10 9 2 13 2 2
12 13 10 10 9 7 13 10 9 0 7 0 2
21 0 2 15 13 1 10 9 1 10 9 0 1 10 9 7 10 9 1 10 9 2
13 10 9 4 13 10 9 7 3 12 9 7 12 2
20 16 13 2 13 10 10 9 2 9 7 13 1 10 9 1 9 1 10 9 2
2 9 2
5 15 13 10 9 2
10 10 3 0 13 10 9 1 10 9 2
13 13 10 9 2 13 3 7 3 2 7 1 9 2
7 3 13 1 13 10 9 2
6 0 2 0 7 0 2
17 13 15 15 1 10 9 3 16 13 10 2 9 2 15 13 0 2
10 3 13 1 10 0 13 1 13 3 2
12 3 13 1 10 9 2 10 9 7 10 9 2
14 13 1 10 9 16 3 13 1 2 13 15 2 3 2
8 13 10 9 7 13 10 9 2
19 1 10 9 13 10 9 1 9 0 0 7 10 9 1 4 15 3 13 2
8 12 9 1 13 15 1 3 2
32 11 11 2 16 13 7 13 10 9 2 11 1 9 7 1 9 2 11 11 11 11 11 11 2 16 13 15 2 11 11 11 2
10 2 7 10 9 1 13 1 10 9 2
18 15 13 1 10 9 1 10 12 7 15 13 10 9 1 10 0 9 2
20 10 9 1 9 0 11 12 15 13 10 9 1 10 9 7 13 1 9 0 2
3 12 9 2
10 9 7 9 1 9 13 1 0 9 2
14 7 1 12 9 15 13 16 13 9 2 9 2 9 2
11 10 9 13 1 9 12 13 12 9 0 2
10 1 10 11 2 11 11 1 11 11 2
6 9 0 9 1 13 15
3 9 9 2
14 9 2 9 2 9 2 9 2 9 2 9 2 9 2
10 3 10 0 9 7 10 9 3 0 2
3 13 3 2
16 10 0 13 10 11 11 11 2 3 10 9 1 10 9 0 2
11 13 3 10 9 7 13 3 15 15 13 2
8 9 2 9 2 9 2 9 2
11 15 13 1 15 2 7 3 13 10 0 2
27 10 9 13 9 0 2 13 7 13 10 9 2 13 9 1 10 9 7 2 10 9 15 13 10 9 0 2
13 7 1 13 3 1 9 13 0 10 9 1 9 2
15 13 13 15 1 9 2 1 9 2 1 10 9 1 9 2
11 3 3 15 4 13 10 9 0 7 0 2
14 10 9 2 3 2 10 9 7 10 9 1 0 9 2
10 16 13 1 9 3 13 3 3 0 2
5 13 15 10 9 2
21 2 16 3 13 0 1 15 2 3 13 15 2 7 13 10 9 13 15 1 9 2
3 2 0 2
36 2 16 13 10 9 1 9 1 15 2 1 10 11 11 2 11 11 12 2 11 2 9 12 2 15 13 1 10 0 9 1 13 15 10 9 2
13 2 16 10 9 13 10 9 2 13 10 9 0 2
5 10 9 13 0 2
30 10 9 0 4 13 1 10 9 0 2 10 9 15 13 1 10 9 7 4 13 1 13 1 10 9 10 9 15 13 2
2 9 2
3 10 9 2
2 9 2
3 12 9 2
2 3 2
13 1 11 2 11 9 12 2 11 2 9 12 2 2
19 2 16 4 2 13 15 10 9 2 2 10 9 3 0 13 1 10 11 2
8 15 13 11 7 13 0 9 2
17 12 9 1 9 1 12 9 4 13 9 1 9 7 9 1 9 2
5 13 1 10 9 2
15 13 10 9 1 10 9 1 9 7 9 1 9 1 9 2
22 13 10 9 2 9 2 2 7 10 0 9 1 13 10 9 1 10 9 0 2 0 2
12 13 10 10 10 9 1 9 7 9 1 9 2
3 13 0 2
16 10 9 0 4 3 13 15 0 7 13 1 9 9 7 9 2
4 13 13 15 2
17 10 9 13 10 9 1 10 9 2 10 9 13 1 9 1 9 2
6 1 9 2 13 9 2
2 9 2
16 16 10 15 13 2 0 2 1 9 2 13 3 0 7 0 2
12 10 9 2 16 13 1 10 9 2 13 0 2
20 16 2 3 2 3 13 1 0 9 15 13 7 15 13 2 13 15 10 9 2
3 10 9 2
13 10 9 2 9 0 2 9 2 9 7 9 0 2
20 16 13 3 0 2 13 16 4 3 13 10 9 0 7 1 9 1 9 11 2
23 16 15 13 3 3 4 13 15 1 10 9 13 1 10 9 2 10 9 15 13 10 9 2
7 1 10 9 13 10 9 2
4 13 15 3 2
11 16 13 0 2 13 15 1 3 12 9 2
10 16 13 0 7 1 9 3 12 9 2
8 9 7 9 0 7 9 0 2
34 0 10 9 0 13 1 0 9 13 0 11 2 15 15 13 16 4 13 10 9 1 10 9 1 10 9 1 9 2 15 1 11 2 2
2 9 2
13 16 10 15 13 2 0 4 13 10 9 1 9 2
11 16 13 0 2 3 13 9 1 10 9 2
18 1 13 1 10 9 1 10 9 13 10 10 9 4 13 10 10 9 2
13 10 9 1 10 9 13 10 0 9 1 0 9 2
11 13 9 0 1 9 1 9 7 10 9 2
14 16 10 9 15 13 3 4 13 15 9 1 9 9 2
4 13 15 3 2
3 3 13 2
15 16 13 1 0 10 9 2 1 9 2 4 13 10 9 2
7 13 15 2 7 3 3 2
22 16 13 1 13 0 2 10 9 0 13 1 10 9 3 0 2 13 2 3 1 3 2
16 13 10 9 3 12 9 1 10 9 1 9 0 7 3 0 2
13 10 9 10 9 0 1 10 9 0 13 10 9 2
11 13 3 10 9 13 3 7 3 13 15 2
10 10 9 3 0 1 10 9 3 13 2
16 16 2 3 2 13 0 2 13 16 9 7 9 15 13 3 2
18 10 9 2 3 2 13 10 9 1 10 0 2 9 7 13 10 9 2
20 13 1 10 0 2 9 1 9 7 9 10 10 9 7 1 10 9 1 9 2
2 9 2
21 16 10 15 13 2 10 3 0 3 16 13 1 10 12 13 10 9 0 1 9 2
12 4 13 15 1 9 0 7 2 3 2 13 2
16 16 10 9 13 3 0 2 9 1 10 9 0 15 15 13 2
8 4 13 15 1 10 9 0 2
7 8 8 8 2 10 9 2
5 13 15 16 13 2
16 1 15 2 13 10 9 2 9 1 3 7 9 1 3 2 2
7 13 15 3 1 9 0 2
13 9 0 1 13 10 9 10 9 16 13 10 9 2
17 9 3 7 3 2 3 16 13 1 10 9 1 10 0 2 0 2
12 1 9 3 10 9 16 11 13 10 10 9 2
13 1 10 9 0 7 0 10 9 1 9 13 9 2
25 1 13 10 9 0 2 11 9 9 2 1 11 2 9 0 1 13 1 10 9 1 10 9 11 2
22 1 9 2 11 11 11 2 1 11 11 1 13 1 10 9 10 9 1 9 7 9 2
30 1 10 0 9 0 2 11 11 1 10 9 2 1 11 15 13 1 13 10 9 1 10 9 13 15 10 9 7 9 2
13 0 3 2 11 11 1 10 9 2 1 11 11 2
16 7 1 10 9 2 9 13 11 2 12 7 12 9 10 9 2
2 9 2
11 3 15 15 13 2 0 2 0 2 0 2
9 15 10 9 0 16 15 3 13 2
14 0 10 9 0 2 9 2 9 1 9 0 7 0 2
11 7 4 13 15 3 1 9 0 7 9 2
4 13 15 3 2
16 16 10 9 13 0 2 10 0 9 0 13 13 15 1 9 2
28 16 10 9 13 0 2 13 3 9 1 10 9 0 2 9 13 2 7 1 10 9 1 10 9 2 13 2 2
42 13 1 13 0 2 13 10 9 1 10 9 1 10 9 7 13 10 9 2 7 1 13 10 9 2 10 9 16 13 2 3 1 10 9 7 1 10 9 1 10 9 2
6 15 13 1 9 0 2
3 9 13 2
18 2 11 11 11 2 1 11 2 13 10 9 0 7 13 10 9 0 2
22 2 11 9 0 1 10 9 2 1 11 2 15 13 10 9 9 13 9 1 10 9 2
2 9 2
19 16 10 15 13 2 1 10 9 1 9 1 9 4 13 16 13 10 9 2
27 9 13 2 9 0 7 0 13 10 9 2 0 2 1 0 9 0 2 9 0 2 9 0 1 10 9 2
4 13 15 3 2
27 1 10 9 2 1 9 9 0 7 9 1 9 10 9 15 13 10 9 2 1 10 9 13 1 9 12 2
32 1 10 9 1 10 9 2 13 13 1 10 9 3 12 9 1 10 9 7 13 10 9 16 4 13 1 13 1 9 1 0 2
32 0 3 10 0 2 9 1 10 9 8 8 2 9 2 9 1 10 9 2 1 11 1 13 1 9 1 9 1 10 9 0 2
21 9 0 7 0 1 10 0 9 2 11 2 1 11 11 7 10 9 2 11 2 2
17 13 10 0 2 9 0 0 2 13 10 9 7 13 10 10 9 2
29 13 15 3 1 9 2 9 10 9 15 15 13 0 2 13 15 1 10 9 2 10 9 7 10 9 1 10 9 2
2 9 2
23 16 15 13 2 11 2 1 9 0 7 0 2 0 2 13 10 10 9 16 15 3 13 2
27 4 13 15 1 0 9 2 1 9 0 2 1 9 0 3 16 2 10 9 2 1 9 3 2 13 2 2
10 10 0 9 13 0 2 10 9 0 2
4 13 15 3 2
11 1 10 9 9 7 9 15 13 7 13 2
16 10 9 0 2 9 9 2 13 10 9 7 13 10 9 0 2
7 13 9 2 9 7 9 2
13 3 2 13 1 10 9 10 9 0 1 10 9 2
2 13 2
16 16 4 13 1 9 7 9 1 13 3 13 3 13 10 9 2
18 1 9 2 13 1 10 9 0 2 13 2 3 15 4 13 10 9 2
6 13 3 9 0 0 2
9 13 15 16 10 9 13 9 13 2
16 10 0 9 0 1 13 1 10 0 9 1 10 9 1 3 2
9 13 13 10 9 1 10 9 0 2
18 10 9 4 4 13 1 10 9 1 10 9 1 10 9 1 10 9 2
21 7 1 9 1 9 1 10 0 9 1 10 9 13 10 9 0 1 9 2 9 2
14 11 11 1 11 2 15 13 1 10 0 7 0 9 2
9 13 15 11 2 7 1 9 2 2
6 10 9 1 10 9 2
2 0 2
15 1 15 0 1 15 0 2 1 10 9 0 1 10 9 2
3 10 9 2
6 15 7 3 15 0 2
24 10 0 9 2 10 9 2 0 2 2 3 13 7 13 3 16 3 15 13 1 10 9 0 2
20 1 13 10 9 1 9 13 13 2 1 0 2 13 15 10 0 9 1 9 2
10 1 10 9 9 2 9 7 9 0 2
7 12 2 13 15 1 9 2
6 13 13 10 9 9 2
25 13 1 10 9 10 9 1 9 16 10 9 1 10 9 13 1 0 2 9 1 9 2 15 13 2
19 12 2 1 10 9 0 13 1 10 9 1 9 2 0 7 0 1 9 2
7 12 2 13 1 10 9 2
6 13 9 1 9 0 2
13 10 9 13 15 1 9 2 9 7 9 1 9 2
15 12 2 13 10 9 2 3 10 9 7 9 1 10 9 2
16 12 2 13 15 10 9 1 12 9 3 1 9 1 9 0 2
5 9 1 10 9 2
8 15 0 15 13 1 10 9 2
19 12 2 13 9 0 7 9 3 0 15 15 13 1 10 9 1 10 9 2
7 12 2 9 1 10 9 2
6 4 13 10 9 0 2
12 15 15 10 9 3 13 2 15 15 13 15 2
13 13 10 11 11 11 2 7 9 1 10 9 0 2
46 13 1 10 9 7 13 1 3 12 9 15 2 13 15 1 10 9 2 10 15 1 10 9 15 13 16 10 10 9 1 9 13 9 7 16 10 9 1 9 0 7 9 0 13 0 2
9 10 9 13 10 9 7 13 0 2
12 2 10 9 0 15 13 3 16 13 10 9 2
10 3 4 13 1 9 2 9 2 9 2
11 15 15 13 0 13 10 9 1 10 9 2
56 15 4 3 13 9 3 0 2 7 0 1 9 0 7 3 2 2 13 1 10 11 1 10 11 1 10 11 2 13 1 10 9 1 10 11 11 1 11 7 15 1 11 1 13 10 9 2 9 1 10 0 11 11 1 11 2
55 10 9 13 10 9 1 9 0 7 0 2 10 9 13 10 9 0 1 10 9 0 1 13 2 15 13 10 9 1 13 1 10 9 7 3 10 9 1 9 1 9 2 9 2 9 9 9 2 7 10 9 1 9 0 2
13 10 9 1 10 11 1 10 11 1 10 11 13 2
14 11 11 2 9 1 11 2 12 2 11 2 9 12 2
9 13 15 13 10 0 0 2 9 2
10 9 0 2 9 0 2 9 1 9 2
3 9 0 2
20 0 2 3 2 13 1 10 9 2 3 3 16 10 9 4 13 1 10 9 2
15 15 13 9 3 2 15 3 13 10 9 1 13 1 9 2
13 13 15 7 2 16 13 13 0 1 10 10 9 2
7 9 9 15 13 7 13 2
6 9 1 9 7 9 2
2 9 2
3 9 0 2
7 0 9 1 10 9 0 2
2 9 2
8 13 10 0 9 1 15 0 2
9 7 16 15 13 3 1 10 9 2
2 9 2
10 15 13 0 7 3 13 10 10 9 2
18 3 1 13 1 10 9 13 1 13 10 0 9 3 1 2 15 2 2
5 3 10 0 9 2
15 2 13 10 9 1 10 9 15 3 15 13 7 13 15 2
5 13 3 10 9 2
26 2 13 10 9 7 10 9 1 9 0 2 9 10 9 11 11 2 1 10 11 1 11 2 1 11 2
17 2 13 1 9 10 9 0 7 9 7 13 10 9 2 3 0 2
13 2 16 1 13 15 1 10 9 2 13 10 9 2
16 2 13 15 13 0 13 7 15 2 3 2 13 0 7 0 2
14 2 3 13 1 10 9 2 7 13 3 1 10 9 2
23 2 3 2 13 16 3 13 10 9 1 13 10 9 2 7 10 10 9 1 0 2 9 2
27 0 9 7 9 1 13 15 1 9 9 9 9 1 9 9 1 9 9 2 9 13 11 2 1 11 11 2
2 9 2
2 0 2
2 9 2
3 12 9 2
14 2 11 13 1 10 9 0 1 10 9 2 1 11 2
2 9 2
2 0 2
2 9 2
3 12 9 2
7 2 11 0 2 1 11 2
2 9 2
5 15 13 1 13 2
2 9 2
3 12 9 2
2 9 2
8 12 2 12 9 1 10 9 2
12 2 11 0 2 9 9 9 2 1 11 0 2
2 9 2
10 1 10 0 9 2 12 9 10 9 2
9 9 2 11 11 12 2 1 11 2
2 9 2
2 0 2
2 9 2
3 12 9 2
2 9 2
17 15 13 10 9 1 9 1 13 10 9 1 10 9 1 10 9 2
7 2 11 11 2 1 11 2
2 9 2
9 10 10 9 2 1 9 7 9 2
2 9 2
3 12 9 2
2 9 2
6 4 13 3 1 9 2
11 9 13 9 2 11 11 11 2 1 11 2
2 9 2
2 0 2
2 9 2
3 12 9 2
13 9 9 2 11 9 9 0 2 0 2 1 11 2
2 9 2
2 9 2
8 12 9 2 12 9 10 9 2
10 9 2 0 2 9 11 2 1 11 2
2 9 2
2 0 2
2 9 2
3 12 9 2
10 9 2 11 11 11 2 1 11 11 2
2 9 2
2 0 2
8 10 9 15 13 1 0 9 2
9 1 9 2 11 11 2 1 11 2
3 9 13 2
2 12 2
5 9 1 10 9 2
2 3 2
6 1 10 9 13 11 2
15 2 9 0 2 12 9 1 10 9 2 1 9 7 9 2
23 2 11 2 1 13 1 10 9 13 1 10 9 12 9 3 1 10 9 7 1 10 9 2
19 9 9 2 15 13 1 10 9 0 1 10 9 1 4 13 10 0 9 2
16 10 9 13 1 2 11 2 13 10 9 1 10 11 1 11 2
2 9 2
26 10 9 0 2 10 9 1 10 9 2 10 9 13 1 10 9 2 10 9 9 0 7 10 9 0 2
5 3 10 10 9 2
16 11 11 1 10 12 2 9 1 10 9 0 1 10 9 11 2
12 1 9 2 11 11 2 10 9 7 10 9 2
3 1 11 11
25 10 9 1 11 2 3 1 12 9 1 10 10 0 9 2 13 1 13 15 3 1 10 9 0 2
24 3 13 3 3 0 10 9 1 10 9 9 2 3 13 1 10 12 1 10 9 1 11 0 2
29 15 4 13 1 9 10 2 9 13 2 1 11 2 1 13 10 9 1 10 0 7 0 9 15 13 10 9 11 2
42 15 13 13 10 0 9 1 11 1 10 9 15 10 9 11 11 4 13 1 10 11 2 9 1 10 9 0 1 11 11 2 7 15 10 10 9 4 13 12 9 3 2
62 0 3 16 15 15 1 11 7 1 11 4 4 13 1 10 0 9 0 1 10 9 3 3 0 2 13 0 1 12 9 1 10 10 0 7 0 9 2 1 11 4 13 2 16 4 13 10 9 1 3 2 10 0 7 0 9 0 2 10 9 0 2
7 13 3 10 0 9 0 2
14 13 10 9 1 13 15 1 3 2 16 13 10 9 2
17 10 0 9 1 10 2 11 2 13 2 16 15 13 2 11 11 2
17 4 13 15 10 0 9 1 11 2 1 3 3 16 11 13 9 2
55 16 10 9 0 2 11 11 2 13 1 10 9 0 7 4 13 3 1 10 9 1 9 2 11 1 10 11 13 1 10 0 9 1 11 7 13 1 10 9 3 1 10 9 0 1 10 9 2 13 3 1 10 0 9 2
18 13 11 15 1 10 0 9 15 1 10 0 12 9 12 13 0 11 2
19 13 11 15 15 15 4 13 0 1 10 9 1 9 10 9 1 10 9 2
6 1 3 12 9 13 2
23 2 3 15 4 13 10 9 2 16 4 13 11 11 1 10 0 9 10 9 1 10 9 2
5 11 15 4 13 2
16 15 4 13 1 10 9 1 10 0 9 15 15 4 13 11 2
11 3 13 16 3 15 4 13 10 9 2 2
9 7 1 12 9 15 15 13 9 2
2 9 2
2 9 2
20 15 13 15 13 16 2 13 10 9 2 10 11 4 13 1 13 15 10 9 2
10 15 2 16 10 9 15 4 4 13 2
54 11 11 13 10 9 1 9 0 2 9 1 10 9 11 2 13 1 0 2 13 1 11 7 10 11 0 2 13 9 0 1 11 11 11 1 15 4 13 3 10 0 9 0 2 11 2 7 3 10 0 9 2 11 2
41 3 15 2 1 11 2 4 13 15 1 10 0 0 9 1 13 1 9 16 10 9 15 4 4 13 1 11 1 10 9 7 10 10 9 0 3 13 1 10 9 2
16 15 13 1 10 9 7 2 4 13 2 13 10 9 1 15 2
52 2 4 13 10 9 1 10 11 2 2 15 13 11 3 2 1 10 9 2 1 9 2 2 1 10 9 1 15 3 15 4 13 9 13 1 10 9 1 11 15 3 4 13 1 13 15 9 2 9 2 9 2
16 7 1 10 11 7 1 10 10 9 15 4 3 13 10 9 2
2 3 2
10 3 4 13 10 9 2 10 9 0 2
10 15 4 13 10 9 1 10 0 9 2
18 7 3 2 1 10 15 15 4 13 2 3 13 16 15 13 3 2 2
2 3 2
6 1 11 2 15 0 2
46 10 0 9 1 10 9 0 15 3 13 9 1 13 12 9 1 10 9 1 11 11 7 1 10 0 9 1 10 9 0 2 15 4 13 3 1 10 13 3 3 10 9 1 10 9 2
34 7 12 9 3 16 11 4 13 1 11 2 1 11 1 10 11 10 0 9 1 10 9 2 11 11 2 13 3 10 9 1 0 9 2
24 7 10 9 3 15 13 3 2 3 1 0 9 2 13 10 9 7 10 9 1 10 9 0 2
26 1 10 0 9 15 15 13 10 10 0 9 2 13 15 1 0 2 1 9 7 9 2 1 0 9 2
14 3 3 15 0 1 10 9 11 7 1 10 11 0 2
12 7 3 15 1 10 9 7 3 1 10 9 2
34 3 1 12 9 1 10 9 1 10 2 9 2 2 10 12 9 10 9 1 11 2 11 11 2 4 13 1 10 0 9 1 0 9 2
7 2 10 9 15 13 2 2
3 10 9 2
23 10 9 0 3 3 13 3 15 13 11 11 2 15 1 12 9 3 4 3 13 1 9 2
13 1 9 0 15 9 3 10 11 2 13 1 9 2
39 3 3 2 1 10 9 15 13 1 11 2 3 13 10 9 1 10 9 1 11 11 2 2 3 4 13 10 0 9 2 3 10 9 2 2 2 3 13 2
13 2 15 4 13 1 4 13 10 9 2 13 15 2
10 2 15 4 13 2 2 13 10 15 2
6 7 15 15 4 13 2
12 13 16 13 0 2 3 3 15 13 3 3 2
17 7 13 0 16 3 10 11 13 1 13 9 2 4 13 1 11 2
24 2 3 4 3 13 10 9 1 10 9 11 11 2 15 15 4 13 15 7 15 4 3 13 2
45 10 9 15 15 13 13 0 7 3 13 10 9 1 10 10 9 2 2 13 3 1 10 11 10 0 9 1 2 0 9 2 7 10 9 3 1 11 1 15 4 13 10 9 13 2
3 9 0 2
9 7 3 16 13 2 9 0 2 2
16 15 13 3 3 3 10 0 11 2 3 1 10 9 0 11 2
26 7 3 1 12 9 10 9 1 11 1 9 1 10 9 4 13 10 2 9 1 11 2 1 10 9 2
29 10 9 0 15 2 1 10 0 9 2 15 13 1 3 13 15 1 10 9 0 2 13 3 0 1 10 9 13 2
44 15 13 1 11 11 2 10 9 1 11 11 2 15 3 13 3 10 3 0 9 0 2 7 3 10 3 0 7 13 9 1 9 1 10 9 0 1 10 9 1 10 9 11 2
19 15 4 13 1 10 9 15 1 10 0 9 1 10 10 9 2 11 11 2
28 2 13 3 16 3 4 13 10 9 16 11 15 4 13 15 15 4 13 3 9 1 11 2 2 15 13 11 2
8 2 3 7 3 15 13 15 2
8 1 10 9 2 13 10 9 2
18 3 16 15 4 13 1 15 1 3 13 15 13 1 10 2 9 2 2
33 1 10 9 0 2 6 2 13 3 10 9 16 15 13 9 0 1 10 2 9 2 2 7 15 3 13 13 1 10 2 9 2 2
5 7 3 2 15 2
16 2 4 3 13 10 9 0 1 10 9 1 11 7 10 11 2
33 13 3 1 15 1 10 9 16 1 10 9 10 9 11 11 13 1 11 1 13 10 9 1 10 9 1 9 1 9 7 9 0 2
28 7 15 13 1 10 9 1 11 2 1 10 9 3 15 3 15 4 13 1 15 3 1 9 1 10 9 0 2
23 7 3 2 10 9 1 9 4 13 1 9 15 1 10 9 15 3 13 10 9 1 3 2
22 15 4 13 6 1 10 9 2 1 10 9 2 1 10 9 1 10 9 15 13 11 2
21 3 16 3 3 13 10 2 9 1 10 9 2 1 13 15 2 7 10 0 11 2
16 7 3 4 13 10 9 1 10 9 1 11 7 1 11 11 2
36 1 9 2 10 9 16 11 11 2 3 1 10 9 0 2 13 1 9 1 9 2 7 11 11 15 4 13 10 9 2 16 11 13 3 9 2
26 7 1 3 10 9 2 1 3 13 10 9 1 15 10 11 4 13 1 10 11 1 10 10 0 9 2
19 10 9 1 11 1 10 0 9 1 15 13 1 9 0 1 10 10 11 2
28 10 9 1 10 2 9 1 9 1 10 11 11 2 1 13 10 9 2 16 1 10 9 10 9 0 4 13 2
21 10 9 1 10 9 1 10 9 0 13 1 10 9 3 13 1 10 9 1 11 2
26 10 9 1 15 1 11 2 3 1 10 9 7 1 10 9 2 7 16 3 13 0 1 10 11 2 2
23 7 3 2 1 10 0 9 1 10 9 1 11 11 2 10 0 9 1 10 9 0 2 2
26 2 13 13 1 11 16 3 11 11 2 1 10 9 1 11 1 10 9 1 10 12 2 13 10 9 2
11 7 3 2 13 2 3 4 13 10 9 2
42 2 1 10 9 1 0 9 1 9 2 16 4 13 10 9 11 11 1 10 0 9 11 11 2 10 0 9 13 1 10 0 9 1 10 9 0 1 10 9 3 0 2
14 7 10 9 3 0 4 13 15 1 10 9 11 2 2
6 2 10 9 15 13 2
9 4 13 10 0 9 15 13 11 2
18 10 9 7 15 1 10 9 4 4 10 9 13 7 1 0 1 9 2
31 16 13 1 13 15 2 9 3 2 1 10 10 9 2 13 3 1 4 13 10 0 9 1 11 1 10 9 1 10 9 2
3 7 3 2
5 2 13 1 11 2
2 13 2
35 2 11 4 13 10 0 9 1 10 9 15 4 3 13 2 1 9 1 10 9 1 10 11 2 16 2 3 13 13 15 1 13 10 9 2
15 3 1 16 13 1 11 10 9 1 10 9 1 10 11 2
81 2 1 9 2 2 13 11 2 2 15 13 3 2 10 9 1 10 9 2 10 9 1 11 11 2 9 1 10 2 9 1 10 3 1 10 9 1 10 12 2 2 7 1 11 11 2 9 1 11 2 7 10 9 1 9 0 13 1 11 1 10 9 11 11 1 10 11 0 4 3 13 10 11 1 10 0 9 1 10 9 2
22 7 3 1 10 9 1 10 3 0 2 15 2 4 13 2 3 13 3 15 13 11 2
22 7 1 10 9 1 10 9 1 12 2 12 9 10 9 1 10 11 13 1 13 13 2
20 3 1 10 9 1 2 9 2 15 15 15 13 10 9 15 15 13 1 11 2
8 10 15 2 13 2 13 0 2
18 16 13 0 16 10 11 13 2 1 10 0 9 2 10 9 1 11 2
24 13 3 1 11 1 10 9 0 11 11 15 13 10 9 1 11 11 11 2 10 9 0 0 2
9 3 13 3 16 13 1 13 2 2
2 11 2
31 12 9 2 15 1 9 2 15 0 2 13 1 9 1 9 2 1 10 9 1 9 2 1 10 9 1 10 9 1 11 2
14 10 9 15 13 1 10 9 7 13 2 9 1 9 2
17 7 3 10 9 13 16 10 9 4 13 1 9 0 7 9 0 2
16 1 10 9 1 10 9 10 2 9 2 13 13 1 10 9 2
61 12 9 2 13 1 9 2 13 1 10 9 2 13 3 1 10 9 1 10 9 4 4 13 2 10 9 3 2 1 10 9 1 11 2 1 11 2 15 9 7 9 0 1 10 0 9 1 9 15 4 13 1 13 10 11 1 10 9 1 9 2
10 10 12 13 3 3 10 12 4 13 2
8 1 9 1 9 7 1 9 2
33 7 15 2 15 3 13 10 11 2 13 1 13 10 9 1 10 9 15 3 13 10 11 2 16 16 15 13 3 9 2 7 9 2
40 15 4 3 13 13 10 9 1 10 9 10 9 0 10 9 1 11 11 15 13 1 10 9 1 10 9 7 12 9 13 1 10 9 1 10 9 1 9 0 2
40 15 4 3 13 16 10 9 1 9 3 2 1 10 11 2 10 9 13 1 10 9 1 9 15 13 1 13 12 9 0 2 13 3 3 10 9 1 10 9 2
37 7 1 10 3 0 13 10 9 15 13 3 9 1 9 0 1 13 10 9 2 1 13 15 1 10 9 1 10 9 7 13 1 9 1 10 9 2
12 10 9 2 16 3 0 3 2 3 3 0 2
23 9 1 9 2 13 1 9 2 1 9 2 1 9 4 13 1 13 10 9 1 10 9 2
43 15 13 10 0 9 0 1 10 9 0 2 3 10 9 1 9 0 13 7 3 13 13 10 9 1 10 9 1 10 9 1 10 9 7 15 13 1 13 15 1 10 9 2
8 15 13 10 9 0 2 0 2
32 15 13 10 9 1 10 9 2 10 9 0 7 13 1 10 11 11 2 1 10 10 9 3 13 7 13 10 9 1 10 9 2
39 3 3 2 15 13 16 10 15 2 10 0 9 1 10 15 15 13 9 1 9 1 10 11 3 13 10 9 1 10 9 15 13 1 13 1 10 9 0 2
19 16 15 13 3 9 1 9 1 10 9 1 11 2 15 13 3 9 13 2
19 7 10 9 1 10 9 2 0 2 3 13 3 15 7 13 0 13 15 2
27 10 9 1 9 15 13 1 15 2 7 3 13 10 9 1 13 10 9 1 9 2 1 10 11 7 3 2
21 3 15 13 10 9 0 7 0 1 10 9 1 10 9 1 9 0 1 9 9 2
25 7 10 0 2 9 2 4 13 3 1 0 9 2 9 7 9 2 1 1 9 1 10 11 11 2
11 3 10 10 11 4 13 1 10 11 11 2
24 15 15 13 0 2 0 2 10 9 0 13 3 3 10 9 1 9 2 10 10 2 9 2 2
23 1 15 2 1 11 2 10 9 13 1 13 15 1 9 1 9 0 2 1 10 9 0 2
38 10 9 1 10 9 7 1 10 10 9 2 13 1 10 0 9 1 10 9 1 10 11 2 7 1 10 10 9 13 0 1 13 15 1 10 9 0 2
46 3 10 9 15 13 1 13 10 9 1 10 9 2 3 2 13 10 9 1 13 10 10 9 1 9 0 1 10 9 1 10 9 2 7 1 9 0 2 1 10 9 7 10 9 9 2
29 6 2 10 9 3 13 1 10 9 2 9 1 11 2 13 10 10 9 2 10 10 9 2 4 13 10 10 9 2
83 1 10 9 15 13 12 9 2 1 10 9 1 10 9 2 1 10 3 12 9 1 9 10 9 2 10 9 15 13 1 11 15 13 1 10 9 2 1 10 9 0 1 10 11 2 1 10 9 16 10 9 3 13 9 1 9 0 7 1 9 0 1 13 15 2 7 13 10 9 0 1 10 9 0 7 3 1 10 9 1 10 9 2
49 13 10 0 2 0 9 1 11 11 1 10 2 9 1 10 9 2 15 4 13 3 2 1 10 10 9 1 9 2 3 1 10 0 9 0 2 3 16 13 10 9 13 7 13 10 11 1 9 2
17 15 13 1 13 10 9 7 15 13 2 1 10 9 2 10 9 2
8 1 9 15 13 10 9 9 2
10 1 10 9 1 10 9 13 10 9 2
17 1 10 9 7 10 9 1 0 7 0 9 15 13 10 9 0 2
3 10 9 2
13 9 2 9 2 9 7 9 13 10 9 1 13 2
7 1 9 3 1 10 9 2
23 11 11 2 9 1 9 1 10 11 9 1 11 2 13 1 10 10 9 3 1 10 9 2
17 10 9 0 0 15 4 13 3 1 10 9 7 1 10 9 0 2
3 1 11 11
23 10 9 0 10 9 1 9 4 13 10 9 1 12 9 1 9 1 3 12 12 9 13 2
23 10 9 0 10 9 13 3 3 16 13 1 10 9 0 1 12 9 1 12 12 9 13 2
49 1 11 13 3 12 12 10 9 0 0 7 1 9 7 3 1 12 12 10 9 3 1 9 15 13 9 2 9 9 2 9 0 2 9 2 9 7 10 9 0 7 0 1 9 1 9 1 9 2
82 1 10 9 10 9 1 9 7 9 9 1 10 10 0 9 4 13 10 9 1 10 9 1 10 9 0 0 7 16 3 15 13 10 0 9 1 10 9 1 10 9 1 10 9 2 13 1 10 9 2 7 15 1 10 9 0 2 3 13 1 10 9 2 2 3 10 9 4 13 1 10 9 16 10 0 13 3 3 9 1 9 2
47 13 0 3 16 10 9 1 10 9 1 10 9 9 2 0 9 7 9 1 9 2 7 1 10 0 2 9 7 9 2 0 1 13 9 1 9 4 13 10 9 3 3 1 10 9 9 2
53 7 1 10 9 0 7 0 2 7 1 10 9 1 0 7 0 9 15 15 13 1 9 0 1 10 9 1 0 9 2 1 13 1 9 7 9 2 10 9 1 10 9 0 13 3 3 0 2 11 9 12 2 2
48 1 10 10 0 7 0 9 15 13 9 0 7 0 2 1 9 7 9 2 13 3 3 9 1 10 9 9 2 10 9 0 15 13 3 1 10 9 1 13 10 9 0 2 11 9 12 2 2
52 1 16 4 13 1 13 15 1 10 9 0 2 13 1 9 11 11 2 9 1 10 3 0 2 0 2 9 1 10 11 2 11 0 1 10 9 1 9 2 2 10 10 9 3 1 13 3 0 13 3 0 2
15 7 10 0 9 1 10 9 1 15 4 13 13 10 9 2
55 13 10 9 3 0 1 15 4 13 10 9 1 10 9 9 7 10 0 9 0 2 1 10 9 1 10 9 1 9 2 15 13 3 9 7 9 2 13 10 9 1 13 3 0 10 10 9 2 3 16 13 3 3 0 2
25 1 9 3 1 10 9 10 0 9 1 10 9 1 10 9 0 15 4 13 10 9 1 10 9 2
54 16 13 1 10 9 10 9 1 0 9 3 0 1 10 9 1 9 2 1 12 9 2 1 10 0 11 12 12 2 7 1 12 9 2 10 9 1 9 4 13 1 10 9 3 0 1 10 12 9 1 9 3 0 2
34 1 10 0 9 1 9 15 13 9 3 7 3 0 1 10 9 2 7 15 13 1 10 9 3 9 0 15 4 13 0 10 9 0 2
46 10 0 9 1 9 2 1 9 1 12 9 2 4 13 1 9 10 3 13 1 10 9 1 9 2 3 15 0 1 9 1 9 7 9 2 2 9 1 9 7 9 1 10 9 0 2
21 13 3 10 9 1 10 9 1 10 9 7 10 9 3 0 9 1 10 9 0 2
16 1 11 15 13 3 12 9 13 1 9 1 12 9 1 9 2
33 10 9 1 9 13 1 12 12 9 2 11 12 13 1 10 11 2 1 12 9 2 11 11 11 5 11 11 13 1 10 11 2 2
41 12 9 13 10 9 1 10 9 2 15 13 1 12 9 1 10 11 11 12 12 1 12 9 1 10 11 11 12 2 9 0 13 1 11 1 10 11 11 11 2 2
37 10 11 3 4 13 1 9 3 10 9 1 12 9 2 10 11 11 11 2 13 1 10 0 9 1 9 3 1 10 0 9 1 15 1 12 9 2
64 3 16 10 0 9 2 1 11 2 11 12 11 7 11 11 12 13 9 0 1 15 0 15 4 3 13 10 9 2 10 9 1 9 1 9 15 13 3 1 10 9 1 0 9 15 13 1 10 9 1 10 9 13 7 15 3 13 9 1 0 9 1 9 2
40 1 9 1 9 13 1 9 1 12 7 12 9 1 9 2 10 0 9 9 3 13 10 9 0 7 13 1 3 10 9 1 13 9 0 2 13 1 9 2 2
26 3 0 7 0 1 13 1 10 15 13 3 10 9 9 2 10 10 9 1 9 0 13 3 3 0 2
21 10 10 9 3 1 10 9 1 10 10 9 15 13 3 1 10 9 1 10 9 2
9 1 9 13 0 10 9 1 9 2
37 4 13 1 0 1 12 9 1 10 9 2 7 10 9 13 15 3 16 10 9 13 3 9 2 16 1 9 0 10 9 1 9 13 3 1 10 2
41 10 0 9 15 13 1 9 10 9 4 13 1 10 9 1 13 3 9 1 10 9 11 12 2 15 13 3 1 10 9 2 3 16 3 0 1 10 9 0 2 2
9 10 9 1 13 13 10 9 0 2
20 10 9 0 1 3 12 9 1 9 13 3 0 1 15 13 1 10 0 9 2
85 1 9 1 10 9 1 10 9 2 10 9 0 1 10 9 0 13 3 12 2 13 1 12 9 2 1 15 13 3 10 9 3 0 1 10 9 1 11 2 15 13 10 9 3 0 2 13 1 12 9 1 9 2 2 11 2 11 11 2 11 2 11 7 11 1 10 9 3 13 2 3 11 2 11 2 11 11 2 11 12 7 11 12 2 2
62 10 9 1 10 9 9 13 3 3 3 13 1 10 9 1 10 9 2 1 10 9 1 10 9 2 10 9 9 11 12 4 4 13 3 1 9 2 7 1 10 9 3 0 2 11 7 11 11 13 0 11 9 1 10 9 1 12 9 1 9 2 2
8 9 1 10 11 0 11 9 2
7 3 10 9 13 9 0 2
2 10 9
11 9 7 9 1 10 0 9 1 10 9 2
32 10 9 1 11 15 13 10 9 1 9 13 10 12 5 10 12 5 13 1 9 7 9 16 4 13 10 9 13 1 10 9 2
41 1 12 9 1 10 12 7 12 9 2 13 2 1 10 9 11 3 10 12 1 12 13 10 9 1 10 9 7 3 10 12 1 12 13 1 9 0 7 1 9 2
79 10 9 13 2 13 1 10 10 9 1 11 7 13 1 10 9 0 7 1 10 3 0 9 0 2 1 10 9 1 10 9 2 1 10 9 1 10 9 2 4 13 1 13 1 10 9 3 1 10 12 1 12 1 10 9 1 15 13 9 0 0 2 10 15 13 1 10 12 1 12 1 10 9 2 1 10 9 2 2
42 10 9 13 4 13 1 10 9 9 0 1 10 12 1 12 1 10 9 2 0 1 10 12 2 0 1 10 12 2 0 7 0 3 1 10 12 1 12 1 10 9 2
34 1 10 12 1 12 1 10 12 9 10 9 9 13 15 7 1 10 12 1 12 13 0 10 9 1 10 9 1 10 9 1 9 0 2
22 3 10 9 13 0 1 10 9 2 3 7 3 2 3 1 10 15 1 10 9 13 2
14 1 10 9 1 9 0 10 9 13 10 12 1 12 2
24 10 9 15 13 1 13 1 10 9 16 13 10 10 9 13 1 10 12 1 10 12 1 12 2
29 1 9 1 9 13 0 13 10 9 1 10 9 13 1 10 9 9 1 10 9 0 1 9 1 10 12 1 3 2
38 10 9 1 9 11 11 4 13 16 10 9 9 13 3 1 10 12 1 12 1 10 9 2 16 1 10 9 0 13 10 12 1 12 1 10 9 0 2
29 10 9 0 1 10 9 4 13 1 10 9 12 2 12 2 9 1 10 15 4 13 10 9 1 9 7 1 9 2
17 10 9 0 13 3 15 1 10 9 7 10 9 1 9 1 0 2
35 1 10 0 9 1 10 9 10 9 13 2 10 9 0 3 1 10 9 2 1 10 9 2 1 10 9 2 1 10 9 2 1 10 9 2
8 1 12 9 3 12 13 13 2
22 1 9 1 15 3 10 9 1 10 9 9 1 10 9 1 10 9 1 10 0 9 2
45 12 9 1 15 12 9 2 12 9 2 12 9 2 12 9 2 12 9 2 12 9 2 10 9 2 10 9 2 12 9 0 7 12 9 4 13 13 1 10 9 1 12 9 0 2
6 10 9 1 10 9 2
15 12 9 1 10 11 2 3 2 10 9 1 11 11 2 2
33 10 0 9 1 11 11 13 3 10 9 1 11 11 11 11 2 16 13 1 11 11 2 13 3 2 1 10 0 9 1 10 11 2
10 1 15 2 3 11 11 13 9 3 2
7 7 10 9 4 13 0 2
26 9 2 9 2 9 2 9 2 9 1 10 9 2 9 2 9 2 9 7 9 2 9 1 10 9 2
35 10 10 11 0 4 13 2 13 2 13 2 13 2 13 9 0 1 10 3 0 9 1 10 11 2 15 1 10 9 3 0 1 10 9 2
18 10 9 11 11 2 13 1 10 11 3 3 15 13 3 2 4 13 2
8 15 13 10 9 1 10 9 2
28 13 1 10 9 1 11 2 13 3 1 10 9 1 12 9 1 9 2 10 11 13 3 0 2 7 3 0 2
33 3 2 13 0 13 16 15 13 1 11 11 4 13 15 15 1 10 9 1 3 0 1 15 0 1 13 1 10 9 1 9 0 2
27 7 3 3 3 13 10 9 1 10 11 2 3 1 10 9 15 13 10 9 1 10 9 7 1 10 9 2
67 13 2 1 9 2 10 9 0 13 1 11 11 2 11 2 9 2 3 1 10 12 9 2 10 9 1 12 9 2 12 9 1 11 11 2 13 2 1 11 2 10 9 7 12 12 9 1 9 0 1 9 7 9 1 9 1 9 7 9 1 10 9 11 2 0 2 2
15 13 10 11 2 10 9 13 1 12 9 7 12 12 9 2
13 1 10 9 3 0 2 15 13 3 10 9 9 2
65 12 9 2 12 9 1 10 11 11 2 1 9 0 1 9 11 2 9 1 11 11 1 9 0 1 9 2 9 1 10 9 3 1 9 2 9 1 9 3 1 11 1 9 1 9 1 9 2 9 1 9 1 10 9 7 10 9 1 10 0 9 1 11 11 2
3 10 9 2
7 12 9 7 12 12 9 2
2 9 2
11 9 12 9 1 11 11 1 10 9 0 2
19 12 9 2 0 2 11 11 13 10 2 13 2 3 1 9 1 10 9 2
25 1 3 1 12 9 1 10 0 9 4 13 1 10 9 1 11 2 3 4 13 1 9 1 9 2
20 1 10 9 0 2 11 11 2 1 10 9 0 7 0 2 3 1 10 9 2
22 3 1 9 2 10 9 1 10 9 0 1 0 9 1 9 1 10 9 1 11 11 2
15 11 11 1 10 9 1 10 11 1 10 9 1 11 11 2
19 1 10 10 9 13 11 11 2 9 1 10 9 7 9 1 10 9 0 2
14 2 4 4 13 10 9 1 9 1 10 10 9 2 2
5 9 1 11 11 2
15 3 10 9 1 13 10 9 13 1 11 1 10 9 0 2
21 3 3 11 2 9 0 2 10 0 2 9 2 1 10 9 2 13 10 0 9 2
28 10 10 9 3 4 13 1 10 9 1 13 1 9 10 12 9 7 12 9 15 13 10 9 1 9 1 11 2
41 3 4 13 3 10 9 0 1 11 11 2 1 10 9 12 9 2 12 9 2 10 9 0 3 1 12 9 3 2 1 10 0 9 1 10 0 9 1 11 11 2
32 12 9 2 9 1 11 11 2 1 9 1 11 2 11 4 13 1 10 9 1 11 3 1 10 9 1 11 11 1 0 9 2
26 13 10 0 9 0 1 10 0 9 4 13 10 9 13 3 1 10 1 3 1 10 9 1 9 0 2
33 12 9 2 12 9 7 12 9 10 9 2 0 9 1 2 9 2 2 10 0 4 4 13 1 10 9 1 11 1 10 9 2 2
3 3 3 2
86 13 10 9 0 1 10 9 2 13 16 15 13 0 1 10 10 9 1 10 0 9 1 10 9 1 11 2 11 11 15 15 4 13 1 10 9 1 13 7 10 9 0 2 1 12 9 1 9 7 12 1 9 1 13 1 11 11 2 16 10 9 15 15 4 13 1 10 10 9 13 9 1 10 10 9 2 15 15 15 13 3 1 13 1 9 2
52 2 4 13 10 9 0 2 2 13 11 2 9 7 9 0 2 9 0 2 0 2 3 0 10 9 2 2 1 10 10 9 4 4 13 1 10 9 1 10 9 0 7 0 2 15 15 4 13 1 10 9 2
52 1 10 9 2 1 10 9 1 10 9 11 7 1 10 9 11 2 12 9 2 10 10 0 9 4 13 1 11 2 10 9 0 13 1 10 9 0 2 15 15 4 13 10 9 7 13 10 9 1 13 3 2
6 10 9 1 10 9 2
54 2 6 2 16 10 10 9 4 13 10 9 2 13 3 15 1 13 1 10 10 9 2 7 1 10 2 9 2 1 9 2 16 10 9 13 7 4 13 3 0 2 0 2 0 2 3 1 15 13 0 1 10 9 2
14 15 2 1 10 9 2 3 3 4 13 1 12 9 2
22 13 1 9 2 4 13 1 13 2 13 1 15 2 13 10 9 2 13 10 10 9 2
57 7 1 10 15 4 13 9 1 10 9 1 15 4 4 13 1 10 9 1 9 1 11 11 2 13 1 10 9 11 11 2 10 9 15 15 13 3 10 9 7 1 10 15 4 13 10 9 1 13 1 10 9 1 11 11 2 2
32 0 2 0 2 0 1 9 7 1 9 2 11 11 4 13 10 2 13 2 3 1 9 1 10 9 3 9 1 10 10 9 2
10 15 15 4 13 1 10 9 3 0 2
14 2 10 0 9 15 13 16 13 1 10 9 1 9 2
19 13 10 12 2 2 13 11 2 2 13 1 13 7 13 1 9 1 9 2
7 10 9 1 10 0 9 2
13 10 9 2 10 9 2 10 9 0 2 10 9 2
10 3 10 9 13 1 13 15 12 9 2
20 4 13 1 10 9 1 9 1 10 9 1 11 1 10 9 1 10 9 11 2
8 1 10 0 9 10 9 13 2
11 7 15 13 3 3 2 15 13 1 15 2
10 1 10 12 10 0 9 0 2 0 2
8 2 10 10 9 13 3 0 2
7 10 0 9 13 10 9 2
9 13 1 11 7 13 10 0 9 2
8 13 12 9 2 0 2 0 2
8 3 10 9 16 13 15 0 2
17 13 1 9 0 1 10 9 1 10 9 1 10 12 1 10 9 2
12 10 9 15 13 3 1 10 12 1 10 9 2
8 16 13 10 9 15 13 0 2
27 13 0 1 10 9 1 13 3 1 15 10 9 15 3 1 10 9 3 4 13 1 10 9 1 10 15 2
7 13 12 9 1 9 0 2
11 10 9 3 13 0 1 10 9 1 9 2
13 1 12 9 7 9 2 3 2 10 9 1 9 2
14 3 13 1 11 1 10 9 10 12 2 12 9 2 2
24 1 10 9 0 1 10 9 1 9 1 10 12 9 1 10 9 1 11 11 10 9 13 0 2
29 2 13 0 1 15 1 15 2 3 1 10 9 2 13 0 1 4 13 10 9 1 9 2 2 13 3 11 11 2
14 2 10 9 9 4 13 1 10 9 1 10 9 0 2
9 15 3 4 3 13 1 9 10 2
10 3 1 9 4 13 10 3 1 9 2
14 1 9 4 13 1 11 11 1 12 9 1 10 9 2
54 1 10 10 9 2 1 10 9 7 1 10 9 1 10 9 2 15 4 13 3 10 9 11 11 2 9 7 9 1 10 9 1 11 11 2 15 15 4 3 13 2 13 2 13 7 15 4 13 3 10 9 3 0 2
30 13 15 1 13 12 9 1 9 2 1 10 0 9 1 15 10 0 9 2 3 0 3 16 13 10 12 9 2 2 2
7 10 9 1 10 10 9 2
14 2 1 11 13 10 9 12 9 7 12 0 9 0 2
22 1 15 3 12 13 10 0 9 1 15 1 10 12 9 0 1 9 1 10 9 0 2
5 3 3 15 2 2
27 1 13 13 10 9 11 11 2 9 1 10 9 1 9 1 11 11 2 9 1 10 9 0 1 11 11 2
23 2 10 9 2 15 4 13 2 4 13 10 2 13 2 1 13 10 12 9 1 10 9 2
17 7 3 13 1 9 1 13 3 10 9 1 10 9 1 10 9 2
21 7 13 0 16 10 9 1 10 11 4 13 10 9 1 10 3 0 9 1 9 2
27 3 15 15 13 10 9 0 13 16 10 10 9 2 1 10 9 1 3 2 4 13 1 3 13 3 9 2
21 13 10 9 16 10 12 1 12 1 10 9 13 13 7 4 13 9 1 10 9 2
12 16 10 12 1 12 4 13 3 10 9 0 2
10 16 3 15 13 10 9 1 9 0 2
6 10 15 3 13 9 2
27 3 3 15 13 16 1 10 10 9 13 3 3 0 10 9 1 9 1 10 9 1 10 12 2 12 9 2
5 9 1 9 12 2
29 7 1 10 9 13 10 9 1 10 9 0 1 10 9 15 4 10 3 13 1 11 10 9 1 10 9 0 2 2
23 9 11 2 3 4 10 9 2 13 2 1 10 9 13 10 9 1 15 1 13 10 9 2
14 2 13 0 2 10 9 1 10 2 9 2 13 13 2
21 1 15 10 9 1 15 15 13 3 4 13 3 0 7 0 2 7 0 7 0 2
49 1 0 9 3 1 10 0 2 3 10 9 2 13 2 4 13 1 10 9 1 10 9 7 15 1 10 9 0 2 1 9 1 9 13 1 10 9 0 7 13 1 10 9 0 1 10 9 0 2
17 10 9 1 11 11 13 1 3 13 3 10 12 9 1 10 9 2
17 3 1 10 12 9 1 9 2 4 13 12 9 1 10 9 2 2
5 15 13 10 9 2
9 2 10 9 13 3 1 9 12 2
11 10 9 4 13 3 1 10 9 1 11 2
21 4 13 0 9 9 7 10 12 4 4 13 1 10 9 1 9 1 0 9 2 2
13 10 9 1 10 9 4 13 10 9 1 11 11 2
27 2 10 0 9 4 13 16 10 9 1 10 9 4 13 3 2 1 15 13 10 9 0 1 10 9 0 2
31 11 4 13 1 10 9 1 9 0 7 13 13 1 10 9 3 10 0 9 13 1 10 9 0 1 10 9 0 2 9 2
17 9 7 9 13 0 1 10 9 3 16 13 1 9 0 7 0 2
19 13 1 10 9 0 7 0 2 13 10 9 2 13 10 9 1 10 9 2
25 10 9 0 2 9 13 10 9 1 9 1 10 9 0 7 10 13 13 3 13 1 9 2 9 2
13 7 3 1 10 9 11 4 13 3 10 9 2 2
13 9 1 11 11 10 9 15 4 13 1 10 9 0
2 9 2
7 10 9 0 1 10 9 2
39 11 2 1 10 11 2 13 10 9 1 12 12 9 15 13 7 13 3 1 9 1 10 9 3 0 1 10 9 7 1 10 9 0 15 3 1 15 13 2
28 3 2 1 10 9 1 10 11 2 13 12 12 9 1 10 9 2 13 2 1 12 9 7 1 12 12 9 2
3 10 9 2
12 10 9 3 0 1 10 9 15 15 4 13 2
14 11 11 11 15 1 10 12 9 13 1 10 11 11 2
15 11 11 13 3 16 15 13 10 9 3 0 1 10 9 2
9 11 11 3 4 13 10 10 9 2
47 11 11 11 11 9 1 9 7 9 1 10 9 11 7 11 11 11 10 9 1 11 11 11 11 10 0 9 13 1 10 11 11 1 10 9 2 10 0 9 15 13 3 1 10 9 11 2
25 11 2 10 9 1 10 11 2 11 2 3 13 10 0 9 2 13 3 1 9 1 10 11 11 2
17 1 10 9 1 9 2 1 3 2 10 9 15 13 10 9 11 2
40 1 3 2 11 11 11 2 10 9 1 10 9 9 16 13 10 9 1 15 10 9 11 2 1 10 9 1 10 9 2 13 10 9 0 1 10 10 0 9 2
26 3 3 2 15 1 10 9 1 9 1 15 10 9 1 10 9 13 3 1 4 13 1 10 9 0 2
33 1 10 12 9 0 1 10 9 1 9 2 10 11 11 11 10 9 0 1 13 10 9 1 12 9 1 10 9 1 10 10 9 2
18 3 3 2 3 16 13 10 9 1 10 9 2 13 2 1 10 11 2
28 10 9 13 0 1 10 9 2 4 13 12 9 1 9 7 4 4 13 1 9 1 10 9 1 10 9 11 2
11 1 10 12 9 0 1 10 9 1 9 2
26 1 9 2 10 9 0 15 13 10 9 1 10 9 1 9 0 15 10 9 4 4 13 1 10 9 2
14 7 1 10 9 11 3 15 4 13 1 10 9 0 2
14 3 3 2 10 9 13 1 9 0 10 9 1 9 2
35 9 1 11 11 9 0 2 11 11 1 10 0 9 1 11 2 15 13 12 9 0 1 13 1 10 9 3 13 1 9 10 9 1 11 2
18 10 0 9 1 9 3 13 7 13 1 9 0 15 13 10 0 9 2
15 9 1 9 16 15 13 3 15 13 10 9 3 3 0 2
5 3 15 13 9 2
8 10 10 9 13 10 9 11 2
25 15 10 9 1 9 2 7 13 15 3 13 9 7 9 2 7 9 3 0 7 1 9 1 13 2
9 13 10 9 1 9 2 1 11 2
17 15 15 13 1 13 15 2 13 15 2 13 3 0 3 13 15 2
33 10 9 11 2 1 3 2 13 1 9 1 10 10 9 10 0 9 1 9 10 10 9 13 13 9 1 9 1 10 9 1 9 2
23 11 13 10 9 0 2 10 9 1 9 1 15 13 1 9 10 0 9 13 1 9 0 2
9 1 10 0 13 1 10 9 11 2
16 10 9 2 10 9 2 10 9 2 10 9 2 15 13 11 2
18 10 9 2 13 1 10 9 1 10 9 2 3 13 15 1 1 15 2
10 3 15 13 11 2 11 2 7 11 2
11 12 12 9 15 13 1 7 9 1 15 2
14 10 9 3 0 1 10 9 4 13 1 9 1 9 2
17 10 9 13 3 2 7 3 15 13 3 15 15 13 1 10 9 2
5 10 9 13 0 2
12 11 13 10 0 9 10 10 9 13 1 11 2
9 10 9 0 1 10 9 13 0 2
7 3 13 3 10 9 11 2
7 15 3 13 0 2 0 2
20 12 12 9 2 12 9 7 12 12 9 10 9 13 1 10 9 1 10 9 2
3 1 13 2
3 3 3 2
20 10 9 11 2 1 9 1 9 2 3 13 15 1 16 13 1 10 9 0 2
11 15 13 1 10 0 9 2 13 1 11 2
8 9 1 9 13 1 12 9 2
32 1 3 10 9 3 13 13 16 3 13 3 1 13 9 7 1 10 9 1 15 2 12 9 1 12 2 15 13 1 10 9 2
18 10 9 1 9 0 13 10 9 1 13 1 10 9 1 10 9 11 2
7 3 15 4 13 1 15 2
6 9 2 9 2 9 2
5 1 9 10 9 2
14 4 13 10 0 1 10 11 1 13 15 1 10 11 2
13 11 11 11 2 13 15 1 10 9 1 10 11 2
30 13 9 1 10 0 9 1 10 11 2 10 2 0 9 2 13 1 11 2 3 15 0 1 10 9 2 1 10 12 2
28 15 13 2 15 13 2 13 1 13 10 10 9 7 1 10 12 13 10 9 2 13 1 10 0 9 0 2 2
8 11 7 11 13 3 15 9 2
13 11 2 10 9 2 13 1 9 10 9 1 9 2
19 9 1 10 9 3 1 10 9 2 13 10 10 9 1 13 15 10 9 2
17 10 9 4 4 13 7 4 3 13 1 10 9 1 10 9 0 2
22 1 10 9 1 10 12 9 2 1 10 12 2 10 9 11 13 3 15 15 13 3 2
6 10 9 1 10 9 2
35 11 15 13 3 7 2 1 3 9 2 10 9 1 9 2 3 1 13 10 9 2 9 2 13 1 13 10 0 2 9 1 9 11 2 2
24 1 13 10 9 13 9 1 10 9 2 9 7 9 15 15 13 9 1 9 1 10 9 0 2
17 13 10 9 3 1 10 9 1 9 2 10 9 3 1 10 9 2
5 15 13 1 9 2
7 15 13 3 1 4 13 2
19 16 10 9 13 0 10 9 13 10 9 2 16 3 4 13 3 12 9 2
20 1 10 9 4 13 10 9 2 15 15 13 12 15 13 1 9 12 9 2 2
7 7 15 13 3 1 3 2
12 15 15 13 1 10 9 0 1 10 10 9 2
19 1 10 9 2 1 9 0 10 9 1 9 15 15 4 1 10 9 13 2
10 1 10 12 15 13 1 10 0 9 2
20 15 13 10 9 3 0 2 10 2 11 11 11 2 13 10 10 9 1 9 2
10 1 10 9 13 10 0 7 0 9 2
13 1 10 9 3 0 2 10 0 9 1 10 9 2
26 13 15 15 2 1 10 9 1 12 15 1 9 2 13 15 15 4 13 10 2 9 1 10 9 2 2
9 10 9 1 12 9 1 9 0 2
13 10 9 1 10 9 13 0 2 7 3 3 13 2
16 1 10 0 9 15 13 3 12 3 0 7 15 13 3 13 2
9 10 0 9 15 15 4 13 13 2
7 2 4 13 9 2 2 2
21 10 9 0 16 10 9 13 4 13 3 10 10 9 1 10 0 9 1 10 9 2
24 13 15 15 2 1 10 9 1 10 9 2 13 7 13 1 10 9 10 9 7 13 10 9 2
38 16 15 4 13 1 11 11 2 9 1 10 2 11 11 11 2 2 10 9 15 13 12 12 9 2 2 10 9 1 9 7 9 13 3 1 0 9 2
24 2 13 1 12 9 16 13 15 13 10 9 1 10 9 1 10 11 7 3 3 15 15 13 2
11 10 9 3 13 9 2 10 9 13 0 2
7 10 9 3 13 3 9 2
14 10 9 3 13 3 3 1 12 9 1 10 9 2 2
11 1 10 12 1 10 12 10 9 15 13 2
28 1 10 12 9 2 0 9 2 2 3 10 9 1 10 9 7 15 15 10 9 4 13 1 10 2 9 2 2
21 10 9 0 2 0 1 10 9 1 10 9 2 13 1 10 9 0 15 13 11 2
11 13 10 9 1 10 9 15 13 1 15 2
18 12 12 9 1 9 13 10 9 1 10 12 9 1 10 0 9 0 2
16 10 9 13 3 1 10 9 1 10 9 13 1 10 10 9 2
19 10 9 2 3 13 1 10 10 9 2 4 13 1 10 9 1 10 15 2
21 10 9 1 10 9 13 1 12 9 7 10 9 0 7 13 1 0 9 1 9 2
17 13 1 10 9 2 0 9 1 9 7 9 0 2 9 1 9 2
11 10 9 1 10 9 13 1 12 12 9 2
64 1 10 9 1 10 9 10 9 13 1 10 0 9 3 10 9 1 9 1 9 13 10 9 15 1 12 12 0 9 15 13 1 13 10 0 9 1 9 2 15 4 13 10 9 1 10 9 11 2 10 9 1 15 15 13 10 9 7 10 9 13 3 2 2
31 11 11 11 2 9 1 10 9 1 9 2 15 13 10 9 1 13 10 9 1 10 15 1 10 9 13 1 10 9 11 2
11 0 9 3 15 4 13 7 13 1 9 2
47 10 9 11 2 9 1 10 9 2 3 4 4 13 1 9 10 0 9 13 2 13 10 10 9 1 10 12 1 3 2 16 16 10 9 13 10 9 13 13 15 15 4 13 10 9 2 2
16 1 9 13 15 4 13 10 9 3 1 10 2 9 9 2 2
21 13 15 3 15 13 3 10 9 15 13 1 13 1 10 9 10 10 9 1 11 2
5 13 13 15 15 2
11 10 9 1 10 9 13 1 10 9 13 2
9 10 9 1 9 13 3 12 9 2
8 12 16 15 4 13 10 9 2
9 12 16 10 9 4 13 3 0 2
24 2 13 3 0 1 10 9 1 10 9 2 2 13 11 11 2 10 0 9 1 10 9 0 2
16 2 10 9 1 10 9 11 13 15 1 13 10 9 1 9 2
6 15 15 4 13 2 2
19 1 3 13 1 10 9 0 2 11 11 13 3 10 9 0 1 10 9 2
18 15 13 16 13 10 0 9 1 10 9 16 13 10 9 1 10 11 2
15 1 10 9 10 9 4 13 1 10 9 1 10 0 9 2
14 15 13 16 3 13 0 1 11 13 10 9 1 9 2
39 3 2 3 2 10 9 13 1 10 9 1 10 9 7 11 4 3 13 9 1 10 9 0 2 1 9 2 3 2 16 10 9 4 13 1 10 9 2 2
12 2 11 7 9 2 2 10 9 1 11 11 2
14 1 10 12 4 4 13 1 10 9 12 9 1 9 2
21 2 4 13 0 9 1 9 1 9 2 7 13 1 10 0 9 1 10 10 9 2
15 15 13 9 2 3 2 15 1 11 3 4 4 13 2 2
9 10 9 10 9 1 3 12 9 2
7 10 2 9 1 9 2 2
3 10 9 2
20 1 10 12 10 9 11 13 10 9 1 9 1 9 1 10 11 1 10 11 2
12 1 10 12 10 9 13 10 10 9 1 9 2
54 10 9 12 9 15 13 1 10 2 11 11 11 1 11 2 2 1 10 2 11 11 11 2 2 1 10 2 11 11 1 11 11 11 2 2 1 10 9 1 12 9 15 13 10 3 0 9 1 9 1 10 9 0 2
26 2 3 2 10 9 0 1 11 13 0 2 10 9 15 13 12 12 9 10 9 2 2 13 11 11 2
15 2 1 15 13 3 1 3 9 1 10 9 1 10 9 2
13 9 15 3 1 10 12 15 4 13 1 13 2 2
13 7 10 11 11 13 1 15 3 0 1 10 9 2
8 1 12 9 13 10 9 0 2
12 2 13 10 9 15 13 1 10 10 9 2 2
36 10 11 11 4 13 1 9 1 11 2 11 2 1 10 9 1 10 12 7 10 15 4 4 13 1 11 2 11 2 1 10 9 1 10 12 2
7 10 9 13 1 10 12 2
12 1 10 9 15 13 1 10 9 10 0 9 2
36 9 0 1 10 9 2 9 0 1 10 9 1 10 9 2 2 3 16 13 15 1 11 15 3 15 13 2 7 9 0 1 0 9 7 9 2
10 7 1 10 12 10 9 13 3 0 2
23 2 15 13 3 1 10 12 1 9 1 10 9 1 10 9 3 2 2 15 13 10 9 2
10 6 3 15 3 13 13 10 9 11 2
21 13 10 9 15 4 13 10 9 0 2 10 9 1 9 2 10 9 2 10 9 2
14 10 9 15 13 7 10 9 3 13 9 1 10 9 2
7 15 13 10 9 0 0 2
15 10 0 9 13 4 13 10 9 2 0 2 1 10 9 2
14 3 1 10 12 15 13 1 0 9 1 10 10 9 2
20 3 4 3 13 10 9 16 3 10 9 4 13 1 10 9 7 1 10 9 2
8 7 3 15 13 15 1 13 2
10 15 13 2 1 9 1 10 9 2 2
6 1 10 9 10 9 2
5 13 15 1 15 2
3 15 13 2
2 9 2
9 1 3 13 10 9 1 10 11 2
3 10 9 2
33 11 11 2 9 1 11 2 9 1 10 11 1 10 12 1 10 12 7 1 9 9 1 10 11 2 1 10 9 0 13 3 0 2
49 10 9 13 13 1 11 10 12 9 1 10 9 1 10 11 13 16 11 11 2 1 10 9 1 10 9 13 10 12 9 12 2 4 13 2 1 10 9 13 15 1 11 2 10 9 1 12 9 2
20 13 1 9 0 2 12 9 1 9 1 10 9 13 1 3 12 9 1 3 2
14 10 9 11 13 9 1 9 1 9 1 10 11 11 2
28 1 13 10 9 2 11 13 10 0 9 1 11 1 15 13 3 15 2 1 10 9 2 15 4 13 10 9 2
16 12 2 12 0 1 10 9 0 1 10 9 10 11 1 11 2
7 12 2 11 0 3 13 2
48 13 0 13 11 2 16 10 9 2 3 0 1 10 0 9 1 10 9 0 2 4 1 10 0 9 1 11 11 13 3 1 0 9 1 10 9 2 16 1 10 0 9 1 10 9 3 0 2
45 10 0 11 2 1 10 9 1 11 2 13 10 9 0 3 1 10 9 2 3 0 2 1 3 12 9 2 1 13 1 10 9 15 2 1 10 10 9 2 13 10 9 3 0 2
12 7 12 9 1 10 12 3 13 10 9 0 2
9 13 1 3 12 9 1 9 0 2
17 3 2 15 13 10 9 2 1 10 9 1 11 7 11 1 11 2
20 3 10 9 13 1 11 13 1 9 11 11 2 13 15 10 9 10 3 0 2
19 13 16 13 1 10 10 9 2 15 11 4 13 1 10 0 9 1 9 2
17 10 9 13 10 0 9 1 10 9 1 11 2 3 13 1 9 2
6 10 9 3 13 9 2
19 1 10 12 10 9 1 11 13 10 9 0 1 10 9 1 10 9 11 2
5 10 9 13 9 2
6 10 9 13 1 11 2
27 10 12 9 12 10 11 13 16 3 13 9 0 7 0 13 1 10 9 1 10 9 2 1 13 10 9 2
42 1 10 11 2 3 13 9 0 16 11 11 13 0 1 10 9 13 1 10 9 12 2 3 1 4 13 1 9 0 1 10 9 7 1 10 9 1 10 9 0 2 2
28 15 13 2 13 0 2 2 13 10 11 2 2 10 9 1 15 0 2 15 13 10 9 1 0 9 3 13 2
19 7 13 0 16 10 9 3 13 10 9 0 2 10 10 9 13 3 0 2
17 3 2 1 9 1 10 9 1 10 9 0 2 10 9 4 13 2
2 9 2
11 7 15 13 10 9 1 10 9 1 11 2
6 11 2 10 3 0 2
36 13 1 10 9 11 2 4 13 1 9 1 10 11 0 1 10 9 1 10 9 1 10 9 1 3 0 9 13 1 11 1 10 9 1 11 2
20 10 11 13 1 11 1 4 13 10 9 1 12 9 1 10 12 7 10 12 2
36 11 13 1 9 1 10 9 7 13 2 1 13 15 2 16 10 9 3 13 1 10 9 4 13 1 10 9 9 0 1 10 10 9 1 9 2
20 10 9 13 0 2 7 11 13 1 10 9 1 10 9 7 10 9 4 13 2
20 1 10 12 10 9 1 11 13 10 9 0 1 10 9 11 15 4 3 13 2
86 10 9 1 11 1 9 11 2 10 9 1 11 2 10 9 1 11 1 9 11 11 1 10 11 2 10 9 1 10 9 1 10 9 0 11 11 2 10 0 9 1 10 9 10 11 11 2 12 9 1 9 1 10 9 7 9 2 12 9 1 9 2 12 9 1 9 2 9 0 1 12 9 7 9 1 9 1 10 9 1 9 1 10 11 11 2
13 10 9 2 10 9 7 10 9 13 1 10 9 2
20 10 9 13 1 1 10 9 1 11 2 7 10 12 9 12 4 13 10 9 2
62 1 13 0 1 10 9 13 1 10 9 12 1 10 9 12 2 13 10 11 2 15 13 10 9 3 3 0 1 10 9 0 0 1 10 9 12 2 12 1 10 9 7 1 10 9 2 7 1 9 3 13 1 10 9 1 10 9 7 1 10 9 2
22 1 10 11 2 15 3 13 10 9 1 11 2 15 13 0 2 3 2 1 9 0 2
5 10 9 4 13 2
73 4 3 13 16 10 9 1 11 2 10 9 1 10 9 2 10 0 0 9 0 2 16 13 13 15 2 2 15 15 1 9 1 10 9 4 13 10 9 13 15 1 10 9 1 13 10 9 1 9 1 13 15 13 9 1 10 9 13 1 10 9 11 2 10 9 3 4 13 10 9 3 0 2
7 12 2 9 1 10 9 2
53 10 9 13 9 1 13 2 12 2 7 13 2 12 2 1 10 9 1 9 0 2 12 2 7 0 2 12 2 2 1 10 9 7 1 10 9 1 10 9 13 1 10 9 0 2 9 12 2 12 2 12 2 2
16 2 12 2 10 9 4 13 16 2 16 7 16 13 10 9 2
28 3 10 3 9 13 10 9 1 13 1 10 9 1 9 0 2 3 10 9 1 9 3 15 13 1 3 9 2
27 2 12 2 10 9 4 13 10 9 1 9 1 10 9 2 4 3 13 15 2 13 15 1 9 2 3 2
16 2 12 2 10 9 4 13 7 13 1 10 9 1 10 9 2
20 9 13 1 10 9 1 10 9 0 2 9 13 1 10 9 1 10 9 0 2
10 10 10 9 1 9 13 10 9 0 2
40 10 9 2 1 3 13 10 9 1 10 9 3 1 10 15 2 3 15 1 10 9 15 13 1 10 9 1 10 15 1 10 0 9 2 13 12 2 12 2 2
3 10 9 2
22 10 9 0 1 10 9 1 9 3 13 3 1 10 9 2 7 13 3 1 10 9 2
15 9 2 13 0 1 10 9 2 10 9 3 4 13 0 2
32 1 13 10 9 1 10 9 13 1 10 9 0 13 13 16 10 9 2 1 10 9 12 2 13 1 10 9 3 10 9 0 2
17 10 9 1 10 9 4 4 3 7 3 13 1 13 10 9 0 2
19 10 9 2 7 10 9 0 2 13 10 9 1 10 15 13 10 9 0 2
5 1 9 15 13 2
45 10 9 1 0 9 2 13 12 2 2 10 9 2 2 13 12 2 10 9 2 10 9 1 10 9 0 2 13 12 2 12 2 2 10 9 1 10 9 0 2 13 12 0 2 2
49 10 9 13 1 10 9 0 2 3 2 13 10 9 1 9 0 2 7 10 9 13 1 10 0 9 1 9 1 10 9 2 9 1 9 2 13 12 2 12 2 2 9 2 13 12 2 12 2 2
8 9 2 13 12 2 12 2 2
55 1 13 0 16 10 9 13 1 10 9 0 3 4 13 1 10 9 2 15 13 3 10 0 9 1 9 0 15 15 13 1 10 9 13 1 10 9 1 13 10 9 1 10 0 9 13 1 10 0 9 2 13 12 2 2
6 12 2 9 1 9 2
25 10 9 3 4 13 9 10 15 3 13 0 9 1 15 1 13 7 13 9 1 15 2 12 2 2
25 9 1 10 9 4 13 16 10 9 12 13 10 9 15 4 3 13 10 9 1 10 9 1 9 2
33 13 15 10 9 0 15 13 10 9 1 15 10 9 0 13 1 13 9 16 4 13 1 10 1 3 1 10 9 13 1 10 9 2
7 12 2 9 1 0 9 2
35 15 4 4 13 1 15 7 1 9 1 10 9 1 10 9 16 3 1 9 1 0 9 2 3 13 2 7 1 10 9 1 10 0 9 2
5 10 10 9 13 2
18 9 1 0 9 2 9 1 10 9 1 13 2 9 1 10 0 9 2
27 1 9 1 10 9 1 10 9 1 10 9 1 9 15 4 13 0 9 1 10 9 7 1 10 9 0 2
42 10 0 4 2 3 2 13 16 10 9 1 9 13 1 9 1 9 4 13 10 0 9 1 10 9 13 1 10 9 2 7 16 3 4 13 10 9 3 0 7 0 2
24 16 13 0 7 0 9 0 2 0 7 0 2 4 4 13 10 9 1 10 9 0 7 0 2
9 1 10 9 4 13 10 0 9 2
12 10 9 0 1 10 9 4 13 1 9 0 2
7 12 2 9 7 9 0 2
44 1 10 9 13 1 10 9 0 10 9 0 2 1 10 9 7 1 10 9 13 1 9 0 2 4 13 1 0 9 7 9 2 9 12 2 1 9 0 10 9 0 7 0 2
46 10 9 1 10 9 15 13 13 16 10 9 1 10 12 4 4 13 10 9 2 1 9 1 9 2 1 4 13 1 10 9 0 7 0 9 1 10 9 7 9 1 10 9 1 13 2
8 10 9 3 4 3 13 9 2
25 1 10 9 1 13 10 9 1 10 9 0 7 0 1 10 9 1 10 9 0 4 13 10 9 2
20 10 9 1 10 9 1 10 9 1 10 9 13 0 1 9 0 2 12 2 2
16 12 2 9 1 9 15 13 10 9 0 7 1 0 9 0 2
92 0 10 9 1 10 9 0 2 9 12 2 7 1 9 2 7 10 9 1 10 9 0 2 2 12 2 7 10 9 0 13 9 0 2 16 10 9 13 10 9 2 10 9 7 10 9 1 9 15 13 10 9 0 2 1 9 1 13 3 1 10 9 1 10 9 0 2 4 13 15 9 1 10 9 1 10 9 1 9 1 10 9 0 2 13 10 9 1 10 0 9 2
25 10 9 1 10 9 0 3 4 13 10 9 2 7 10 9 1 10 9 0 4 13 15 3 0 2
46 16 1 9 1 9 0 1 10 15 7 1 10 0 9 15 13 0 10 9 1 10 9 0 1 10 9 2 4 13 10 9 1 10 9 1 10 9 1 15 10 9 0 4 13 9 2
20 10 9 13 10 9 0 1 10 9 2 13 1 10 9 0 2 13 12 2 2
27 3 0 10 9 13 1 10 0 9 2 15 13 9 1 10 9 0 1 10 9 1 13 10 0 9 0 2
40 10 0 9 15 13 16 10 9 1 10 9 13 1 9 1 13 3 1 10 9 1 10 9 7 1 10 9 1 10 9 2 1 10 9 7 1 10 9 0 2
22 10 9 1 10 9 13 1 13 16 10 9 1 10 9 13 10 9 1 10 9 0 2
10 3 13 16 10 9 4 4 3 13 2
9 12 2 9 1 9 0 7 0 2
40 10 9 1 9 0 2 0 7 0 2 15 13 9 0 2 0 2 0 7 0 2 12 2 2 9 12 2 4 13 1 10 9 1 10 9 0 2 12 2 2
10 12 2 9 7 9 13 1 10 9 2
39 10 9 1 10 9 15 13 1 10 9 2 1 10 15 15 15 15 13 2 12 2 2 7 10 9 4 13 10 9 7 9 15 3 13 9 1 10 9 2
26 10 9 3 15 13 1 15 13 9 1 10 9 1 10 9 2 9 7 9 2 12 2 2 12 2 2
42 13 1 10 9 0 10 9 13 1 10 9 1 10 9 7 0 9 2 12 2 2 1 10 9 2 12 2 2 1 10 9 0 7 1 0 9 0 2 9 12 2 2
43 10 9 1 10 9 3 4 13 15 1 9 1 15 15 15 13 1 10 9 1 10 9 7 1 10 9 1 10 9 13 2 12 2 2 16 15 3 13 9 1 13 15 2
7 12 2 9 1 10 9 2
16 10 9 4 13 2 12 2 1 10 9 10 9 2 12 2 2
20 10 9 1 13 10 9 13 15 1 10 9 1 10 9 1 10 9 1 9 2
16 10 9 15 13 1 13 7 13 15 3 13 1 10 9 12 2
6 12 2 9 7 9 2
53 10 9 1 10 9 3 4 13 16 15 15 13 1 10 9 1 10 9 2 1 3 16 10 9 4 13 2 12 2 2 1 10 9 13 1 10 9 1 10 9 2 12 2 7 15 13 9 1 9 0 1 9 2
16 1 10 9 1 10 9 13 10 9 1 10 9 1 10 9 2
7 12 2 9 1 10 9 2
50 10 9 4 13 10 9 2 12 2 7 10 9 1 10 10 9 2 3 16 15 4 13 10 9 2 12 2 2 1 10 9 1 13 7 13 10 9 7 10 9 10 1 10 9 7 0 2 12 2 2
12 16 10 9 13 9 2 4 13 10 0 9 2
32 10 9 4 3 13 10 9 1 15 4 13 10 9 10 15 15 15 13 3 7 10 9 15 15 15 4 13 13 1 10 9 2
16 10 9 4 13 10 9 13 10 9 7 10 9 2 12 2 2
22 1 10 13 10 9 10 9 0 4 13 10 9 1 10 9 1 10 9 1 10 9 2
14 4 13 9 1 10 9 1 10 0 9 2 12 2 2
25 10 9 13 9 1 9 0 2 7 13 3 0 3 1 10 9 2 7 1 15 13 1 10 9 2
59 3 13 2 3 2 15 13 16 10 9 12 2 3 4 13 1 10 9 1 13 10 9 0 2 4 13 0 9 1 9 1 10 9 2 1 10 9 1 10 9 12 9 2 0 3 1 10 9 2 15 13 1 10 9 2 13 9 13 2
8 10 9 13 2 3 2 0 2
19 1 13 13 10 9 0 10 9 4 13 1 10 9 13 1 10 9 12 2
19 16 1 10 9 13 0 13 3 10 9 2 10 9 4 13 10 9 12 2
10 12 2 9 0 1 9 1 0 9 2
37 10 9 0 13 0 1 9 0 1 10 9 1 9 1 0 9 1 10 9 13 1 10 9 0 2 12 2 7 1 10 9 13 1 10 9 0 2
25 10 9 15 13 1 13 15 13 1 10 9 2 9 12 0 2 7 1 13 1 10 9 12 0 2
6 12 2 0 9 0 2
59 1 10 9 1 9 2 1 10 9 7 1 10 9 1 10 9 2 13 1 9 9 13 1 9 7 0 1 9 2 7 1 10 9 7 1 10 9 1 9 0 1 10 9 0 3 4 13 15 9 1 9 15 3 13 10 0 9 0 2
47 15 13 1 0 9 0 10 9 1 9 0 7 0 1 10 9 1 10 9 0 7 2 16 3 15 13 1 9 0 2 12 2 2 1 13 10 0 9 1 10 9 1 10 0 9 0 2
33 10 9 13 10 9 1 10 9 1 9 1 10 9 2 13 12 2 1 10 9 1 10 9 0 2 3 2 1 13 10 9 0 2
17 10 9 13 10 9 1 10 9 1 9 0 1 13 10 0 9 2
29 10 9 3 13 3 10 9 1 9 1 10 9 1 10 9 0 2 7 3 10 9 1 9 1 9 0 1 9 2
9 12 2 9 1 10 0 9 0 2
49 10 9 1 10 0 9 0 4 13 3 1 9 2 13 9 1 10 9 0 7 1 10 9 0 0 2 1 9 1 10 9 0 2 12 2 2 2 1 13 15 13 10 9 0 2 2 12 2 2
40 10 0 9 1 10 9 1 9 1 10 0 9 0 4 1 10 15 13 2 13 0 2 10 0 9 1 10 9 1 10 9 0 13 1 10 9 1 10 12 2
7 12 2 9 1 10 9 2
25 10 9 13 1 10 9 1 10 9 12 4 4 13 1 10 9 0 2 1 9 1 10 0 9 2
16 10 9 15 13 1 12 9 1 10 9 1 9 1 10 9 2
9 12 2 9 0 1 0 9 0 2
66 3 1 10 9 1 10 9 13 1 10 9 0 2 10 9 1 9 1 10 15 4 13 9 13 1 15 2 1 9 0 1 10 0 9 0 2 4 13 16 15 4 13 10 9 1 10 15 2 13 15 10 9 2 1 10 9 1 13 10 0 9 1 10 9 0 2
29 1 9 1 9 13 10 9 0 2 13 10 9 0 2 12 2 1 10 9 1 10 9 15 13 10 9 1 9 2
25 1 13 10 0 9 7 9 1 10 9 0 10 9 4 13 10 9 1 10 9 1 10 9 0 2
50 10 9 13 10 9 0 1 13 1 10 0 9 2 7 1 10 9 2 1 10 9 13 1 10 9 12 2 10 9 1 10 9 1 9 0 1 10 0 9 0 13 1 15 15 4 13 1 10 15 2
25 10 0 9 1 10 9 1 10 0 9 0 4 13 10 9 2 1 10 15 2 1 10 15 0 2
9 12 2 9 1 9 1 9 0 2
64 16 10 9 0 7 0 1 10 0 9 0 13 1 10 9 2 4 2 1 9 1 15 1 10 13 7 1 9 1 10 9 0 2 4 13 10 9 2 12 2 1 10 0 9 2 1 10 9 1 13 1 10 9 0 0 1 10 0 9 1 10 9 0 2
17 1 10 9 1 10 9 15 13 10 9 13 1 10 9 1 9 2
40 10 9 1 10 9 4 4 13 1 10 9 3 1 9 1 9 2 13 12 2 2 9 0 2 13 12 2 2 9 0 1 10 9 2 13 12 2 12 2 2
5 12 2 9 0 2
14 10 9 13 1 10 9 0 4 13 10 9 1 9 2
18 1 10 0 9 1 10 9 0 4 13 15 1 9 7 1 9 0 2
14 4 3 13 15 1 9 1 9 7 1 9 1 9 2
8 12 2 9 13 1 10 9 2
12 1 10 9 0 13 1 10 9 0 4 13 2
13 12 2 10 9 13 1 9 1 9 0 7 0 2
15 12 2 10 9 0 1 10 9 7 13 9 1 10 15 2
11 12 2 10 9 2 10 9 2 10 9 2
17 12 2 10 9 0 1 9 7 9 1 9 1 9 0 7 0 2
16 12 2 10 9 0 1 9 2 1 9 7 1 0 0 9 2
25 12 2 10 9 15 1 10 10 0 9 2 9 7 9 1 9 13 9 1 0 9 2 12 2 2
8 12 2 9 1 10 9 0 2
29 1 10 9 0 2 12 2 10 9 0 4 13 2 13 7 13 1 9 1 10 9 1 10 0 9 2 12 2 2
54 10 0 9 0 1 9 4 13 1 10 9 13 1 9 7 2 16 3 4 13 1 10 10 9 1 10 0 9 2 4 13 3 1 10 9 0 1 10 9 13 1 9 2 15 13 1 9 1 10 9 1 15 13 2
36 10 9 15 3 4 13 1 10 10 9 1 10 0 9 4 13 1 10 9 1 0 9 1 10 9 13 1 9 1 10 9 1 15 4 13 2
50 1 9 1 9 13 1 10 9 13 1 9 1 10 9 2 10 9 4 13 1 9 7 10 9 4 13 2 1 10 9 1 10 9 2 1 10 9 1 10 9 13 1 10 9 0 1 10 9 0 2
11 12 2 9 7 9 1 10 9 1 9 2
37 10 9 1 9 4 4 3 13 1 9 1 10 13 2 7 3 1 15 4 13 9 1 9 0 2 1 10 9 7 1 10 9 13 1 9 0 2
31 10 9 0 1 9 0 1 10 9 4 4 13 1 10 9 1 10 9 0 1 10 10 9 4 13 10 9 2 12 2 2
12 12 2 9 1 10 9 1 10 9 1 9 2
27 1 10 9 1 10 9 1 9 2 12 2 15 13 10 9 1 9 7 1 10 0 9 0 2 12 2 2
16 4 3 13 10 9 13 1 10 9 0 2 12 2 12 2 2
8 12 2 9 1 10 9 0 2
29 1 10 9 13 1 10 9 12 7 0 13 0 10 9 1 10 9 0 0 1 10 9 1 10 9 1 10 13 2
36 10 9 0 3 4 3 1 10 10 9 13 10 9 1 10 9 1 9 2 7 4 13 1 10 9 7 9 1 9 1 10 9 1 15 13 2
7 12 2 9 0 1 9 2
85 1 10 9 1 9 0 2 0 2 0 7 1 0 9 0 4 4 13 0 1 9 10 9 15 15 13 1 10 9 2 1 15 13 9 2 9 2 9 7 9 0 2 7 13 1 9 0 13 1 10 9 0 7 0 2 7 1 9 3 13 1 0 9 1 9 0 7 0 2 10 15 13 0 1 10 0 9 1 10 9 0 2 12 2 2
48 10 9 0 1 10 9 0 4 13 1 10 9 1 10 9 0 2 12 9 12 2 9 12 2 10 9 2 1 10 9 2 15 13 1 13 10 9 3 13 1 15 7 1 10 0 9 0 2
31 10 9 0 1 10 9 0 13 1 15 0 1 10 9 7 9 2 7 13 3 1 9 1 10 9 2 13 9 12 2 2
26 10 9 1 9 7 10 9 0 1 10 9 7 1 9 0 4 13 7 13 1 9 1 10 9 0 2
9 12 2 9 1 9 1 10 9 2
23 10 9 0 13 1 10 9 0 13 10 9 1 9 13 1 9 1 10 9 2 12 2 2
10 12 2 9 1 10 9 1 10 9 2
46 10 9 1 10 9 13 1 10 9 1 10 9 4 13 1 13 1 10 9 0 2 12 2 1 10 9 2 10 9 7 10 9 1 10 9 1 9 1 10 9 15 13 1 10 9 2
9 12 2 9 1 9 1 10 9 2
54 10 9 1 10 9 13 1 10 9 0 4 13 1 13 2 1 9 1 10 9 0 1 9 7 1 10 13 9 1 9 0 2 10 9 1 9 0 15 13 1 9 0 1 10 9 7 1 9 0 1 15 1 15 2
6 12 2 9 1 9 2
28 1 10 9 2 1 10 9 7 1 10 9 1 10 9 1 9 4 13 15 1 9 1 9 1 10 9 0 2
34 1 10 9 4 4 3 13 10 9 2 10 9 7 10 9 1 10 0 9 1 9 0 1 10 9 7 1 9 0 1 15 1 15 2
28 10 9 4 13 1 9 1 10 9 1 10 9 7 2 1 9 1 10 9 0 2 4 4 13 3 1 9 2
19 15 13 9 0 0 7 13 10 10 9 1 10 9 13 1 10 9 0 2
7 12 2 9 1 9 0 2
42 1 10 9 13 1 10 9 1 9 4 4 13 3 9 1 10 9 2 10 9 7 10 9 1 10 9 1 9 0 0 1 10 9 7 0 1 10 9 0 1 9 2
6 15 13 9 0 0 2
48 4 3 13 10 9 1 9 0 0 16 2 1 10 10 0 9 0 7 1 10 0 9 1 10 10 9 1 10 9 1 10 9 1 10 9 2 4 13 1 9 0 1 9 1 10 9 0 2
5 12 2 9 0 2
40 10 9 1 10 9 1 10 9 1 9 2 9 7 9 1 10 9 1 9 7 1 9 0 13 0 1 10 9 7 10 9 13 1 10 9 0 2 12 2 2
9 12 2 9 1 9 1 10 9 2
54 16 10 9 1 10 9 13 1 10 9 2 12 2 12 2 13 0 1 13 10 9 1 10 9 1 9 2 4 13 15 9 1 10 9 0 7 0 1 10 9 13 1 10 9 0 2 13 10 9 1 10 9 0 2
37 10 9 13 9 1 9 1 10 9 2 16 15 15 13 9 2 7 2 1 9 2 1 9 1 10 9 15 15 13 1 13 10 9 13 0 9 2
11 12 2 9 1 9 0 7 1 0 9 2
63 3 3 1 10 9 1 9 2 12 2 12 2 2 10 9 1 10 9 7 9 4 4 13 1 9 0 2 13 10 9 7 10 9 13 1 10 9 0 2 1 10 9 1 13 16 4 1 9 0 13 9 2 13 10 9 7 13 10 9 1 10 9 2
45 10 9 1 10 9 7 10 0 10 9 2 10 9 1 10 9 2 10 9 1 10 9 7 1 10 9 4 13 2 1 9 1 10 9 2 1 10 9 13 1 10 9 1 9 2
64 3 2 1 9 1 10 9 0 2 4 4 13 1 9 1 10 10 9 10 9 15 1 10 10 0 9 13 9 7 9 1 10 9 1 9 2 1 10 9 1 10 9 2 1 10 9 7 1 10 9 1 10 9 2 7 15 13 0 1 10 9 0 0 2
18 10 9 0 13 10 9 1 0 9 0 1 15 0 2 1 15 13 2
38 8 2 10 9 1 9 1 9 0 13 1 10 9 12 9 9 12 1 10 12 2 15 13 10 9 1 15 15 13 0 10 9 1 9 1 9 0 2
39 8 2 9 0 13 1 10 9 12 2 12 2 12 2 9 12 2 0 9 11 2 15 4 13 10 9 1 9 1 10 9 1 10 9 1 0 9 0 2
46 1 10 9 1 10 9 7 1 10 9 10 9 13 4 4 13 1 9 2 1 9 0 7 1 9 1 10 9 1 10 9 2 1 10 9 7 1 10 9 13 1 10 9 1 9 2
10 12 2 9 0 1 10 9 1 9 2
65 10 9 1 9 13 1 9 1 9 1 9 15 13 7 13 9 1 10 9 2 1 9 7 1 9 1 9 0 4 13 2 3 3 1 10 9 1 9 2 1 13 1 10 9 1 10 9 0 1 10 9 1 10 9 1 9 1 10 9 13 1 10 9 0 2
5 12 2 9 0 2
37 10 9 1 9 1 10 9 3 4 13 9 0 2 12 2 4 13 10 9 1 10 9 0 1 10 9 7 1 10 9 7 9 1 10 9 13 2
50 16 4 13 10 9 1 9 2 12 2 2 13 9 0 1 0 9 1 9 7 1 9 2 10 13 9 1 10 9 13 1 10 9 4 13 10 10 0 9 1 9 1 13 0 10 9 1 10 9 2
13 4 3 13 15 1 9 1 10 9 1 10 9 2
19 1 9 1 9 2 4 13 15 1 10 9 1 9 1 10 9 1 9 2
10 12 2 9 1 9 7 1 9 0 2
21 10 9 1 13 15 1 10 9 4 13 1 10 9 0 7 1 10 9 0 0 2
18 10 9 0 13 3 10 9 1 13 15 1 10 9 1 10 9 0 2
9 12 2 9 1 10 9 1 9 2
49 15 15 1 9 1 10 9 4 13 9 4 4 15 13 2 0 10 9 1 13 10 9 1 9 2 12 2 16 15 13 1 10 9 1 10 9 0 1 10 9 0 7 1 15 13 2 12 2 2
7 12 2 9 1 10 9 2
30 10 9 1 9 0 2 16 3 4 13 7 0 2 4 4 13 2 12 2 1 9 3 0 1 12 9 2 12 2 2
14 1 10 9 0 4 4 13 10 9 0 2 12 2 2
17 10 9 1 10 9 13 10 9 1 10 9 0 1 10 9 0 2
10 15 15 13 3 1 10 9 3 0 2
29 10 9 1 10 9 13 1 13 16 15 13 9 0 2 7 1 13 9 0 1 9 2 9 7 9 1 10 9 2
12 1 10 9 0 10 9 0 13 1 12 9 2
11 12 2 9 0 1 10 9 1 10 9 2
41 10 9 1 10 9 0 1 10 9 10 4 13 15 10 9 2 12 2 2 1 10 10 9 7 1 9 1 15 2 16 15 13 1 10 10 9 1 10 10 9 2
43 1 13 10 9 4 13 2 12 2 10 9 1 10 9 1 10 9 2 7 1 10 9 1 9 13 0 2 7 10 9 1 10 9 1 10 9 1 15 10 9 4 13 2
14 12 2 9 0 1 10 9 15 3 13 1 10 9 2
98 16 10 9 15 13 1 10 9 1 10 9 0 1 10 9 7 9 7 1 9 0 1 10 9 1 15 13 1 10 9 0 2 10 9 4 13 10 9 1 10 9 2 12 2 12 2 3 1 10 9 1 13 2 12 2 1 10 9 0 2 13 2 1 10 9 1 10 9 1 10 9 2 10 9 1 10 9 1 13 1 10 0 9 2 3 16 10 9 13 13 10 10 9 3 1 10 9 2
29 10 9 15 13 13 10 9 4 13 3 10 9 16 13 1 13 10 9 1 10 9 7 1 13 1 10 10 9 2
35 15 4 13 10 10 9 1 10 9 1 9 12 7 4 13 1 10 9 7 1 10 9 1 12 9 1 10 9 1 15 4 13 10 9 2
10 12 2 9 1 10 9 1 10 9 2
21 10 9 12 13 1 15 13 1 10 9 12 7 10 9 1 10 9 13 3 0 2
34 10 9 4 13 16 10 9 4 13 1 13 10 9 0 1 10 0 9 15 13 1 10 9 16 15 13 0 3 10 9 1 10 15 2
6 12 2 9 1 9 2
40 10 9 2 1 13 10 9 1 10 9 2 12 2 13 1 10 9 2 4 13 1 10 9 0 1 9 2 7 1 13 2 12 2 10 10 9 1 15 0 2
14 10 9 15 13 3 1 10 9 13 1 10 9 12 2
14 10 9 1 10 9 4 13 3 10 9 1 10 9 2
6 12 2 9 1 9 2
37 10 9 1 9 7 10 0 9 0 15 3 13 10 9 0 1 10 12 9 3 4 13 1 10 9 1 10 9 13 1 10 9 12 2 12 2 2
39 15 2 16 4 13 1 10 9 2 4 4 13 0 3 1 9 1 9 2 16 3 13 1 10 1 3 10 9 1 9 0 1 10 12 9 2 12 2 2
16 12 2 9 3 0 1 10 9 1 10 9 7 1 9 0 2
47 1 10 9 0 3 13 0 10 9 13 1 10 9 0 7 15 0 1 10 0 9 2 12 2 2 7 10 9 15 4 13 1 9 0 2 0 7 0 2 1 9 1 10 9 1 9 2
15 10 9 3 4 3 13 1 10 9 13 1 10 9 12 2
38 1 10 9 15 15 13 1 9 1 10 9 7 10 9 0 3 15 13 10 9 0 1 10 9 2 7 4 13 15 10 9 7 10 9 15 15 13 2
22 10 9 1 10 9 1 10 9 0 7 1 10 9 3 13 10 9 0 0 7 0 2
33 13 13 16 16 10 9 3 4 13 10 9 0 1 10 9 0 2 10 9 4 13 10 9 1 10 9 0 1 9 1 10 9 2
22 10 9 13 9 1 10 9 1 13 10 9 1 10 9 0 15 10 9 0 4 13 2
10 12 2 9 1 9 1 10 9 0 2
46 10 9 15 13 1 9 1 9 15 13 0 2 12 2 1 1 10 10 9 7 2 1 9 1 9 0 2 1 1 10 9 1 15 15 1 10 9 13 1 13 3 0 2 12 2 2
29 15 13 3 0 10 9 15 13 1 9 1 9 2 9 7 9 7 1 9 1 10 9 2 12 2 2 12 2 2
11 12 2 9 1 9 0 1 10 9 0 2
39 15 13 2 12 2 16 10 9 0 1 10 9 2 9 2 9 7 9 13 1 10 9 1 10 9 1 10 15 13 10 9 7 1 9 1 10 9 0 2
69 16 13 9 2 1 9 2 9 7 0 2 7 9 15 15 13 1 10 9 1 10 9 1 10 9 2 7 10 15 7 10 15 13 13 1 10 9 0 2 15 13 16 15 13 1 10 9 1 10 10 9 10 9 7 10 9 15 13 2 3 16 15 13 3 15 1 10 9 2
26 16 15 7 15 1 15 13 1 10 9 2 7 15 7 15 1 10 9 0 2 10 9 4 13 0 2
8 12 2 9 1 10 9 0 2
51 10 9 7 10 9 0 2 12 2 1 10 9 0 13 1 9 1 10 15 15 15 13 9 7 1 9 1 10 9 1 15 2 3 16 10 9 4 4 13 1 10 9 1 15 1 10 9 2 12 2 2
48 10 9 1 10 9 0 4 13 15 1 10 9 1 13 1 10 9 1 9 7 9 2 13 1 10 9 1 9 2 16 10 9 0 3 13 10 9 1 10 9 2 12 2 12 9 12 2 2
11 12 2 9 1 9 13 1 10 9 0 2
42 10 9 15 4 13 10 9 13 1 10 9 0 4 13 1 10 9 1 15 2 7 4 13 15 10 9 7 10 9 15 10 9 13 0 1 13 10 9 1 10 9 2
14 12 2 9 7 9 1 9 7 9 1 10 9 0 2
80 10 9 1 10 9 0 4 13 13 15 2 12 2 10 10 9 7 4 13 15 9 2 16 15 13 1 9 1 12 9 1 10 9 0 2 0 10 9 1 10 0 9 1 13 13 10 9 1 1 10 9 1 10 9 2 1 10 9 1 15 15 4 13 10 9 1 10 0 9 2 13 15 10 9 7 13 15 10 9 2
20 10 9 4 3 13 10 9 0 1 9 7 9 1 9 2 13 10 0 9 2
16 15 4 13 1 10 9 1 13 10 9 13 1 10 9 13 2
27 3 4 13 9 1 10 9 0 2 7 13 15 10 9 15 15 13 10 9 7 15 1 0 9 15 13 2
28 9 3 0 2 1 16 2 13 10 9 1 9 1 10 9 0 2 13 1 10 9 1 10 9 12 2 12 2
41 10 9 1 10 9 1 10 9 2 13 12 2 12 2 13 1 10 9 16 15 4 13 10 9 13 1 10 9 3 4 13 10 9 1 10 0 9 1 10 9 2
8 12 2 9 1 10 9 0 2
16 3 15 4 1 10 9 4 13 0 1 9 1 10 9 12 2
28 16 10 9 3 13 0 1 13 10 9 2 15 15 15 13 4 13 1 13 15 7 1 13 15 1 10 9 2
32 1 10 0 9 15 13 0 2 10 9 4 4 13 1 10 9 10 2 3 16 9 0 13 1 13 15 1 15 1 10 9 2
31 1 10 10 9 10 9 13 7 13 13 1 9 0 2 7 10 9 4 4 13 1 10 9 13 1 10 9 1 10 9 2
25 1 10 0 9 10 9 13 9 1 13 3 10 9 1 10 9 1 10 9 13 1 10 0 9 2
40 16 10 9 4 13 10 9 1 10 9 13 1 10 9 2 15 13 9 2 1 10 13 10 9 1 15 2 3 1 10 9 13 1 10 9 7 1 10 9 2
12 10 9 13 10 9 1 10 9 1 10 9 2
29 3 15 1 10 9 4 2 1 13 10 9 1 10 9 2 13 10 9 0 2 13 3 9 0 1 10 9 13 2
9 12 2 9 1 10 9 1 9 2
43 15 4 13 10 9 1 13 1 9 1 10 9 2 12 2 1 9 1 9 1 9 2 12 2 15 13 10 0 9 2 10 9 7 10 9 13 1 10 9 2 12 2 2
25 10 9 1 15 2 16 3 4 3 13 1 10 9 0 7 1 10 9 2 4 13 1 12 9 2
9 12 2 9 1 9 1 10 9 2
64 16 1 12 9 13 1 10 9 15 13 0 7 10 15 0 2 12 2 2 10 9 1 10 9 0 4 13 1 9 10 9 1 9 7 9 1 10 9 1 10 9 1 10 9 1 10 10 9 2 12 2 2 7 10 10 9 4 13 1 10 10 13 9 2
25 10 9 4 4 13 1 9 1 10 9 1 10 9 0 7 1 9 1 10 9 1 10 9 0 2
10 12 2 9 1 10 9 1 10 9 2
46 10 9 15 4 13 1 10 13 1 10 9 1 9 1 10 9 1 9 7 0 2 13 2 12 2 2 1 9 1 9 2 10 9 1 10 9 1 15 10 9 1 9 4 4 13 2
55 1 10 9 10 9 13 1 9 1 15 15 15 4 13 2 0 10 9 1 10 9 1 13 15 0 1 10 9 1 10 9 12 2 1 10 9 3 1 13 10 9 1 10 9 1 10 9 1 15 10 9 4 4 13 2
55 15 4 13 9 2 9 2 12 2 2 9 1 9 7 1 9 1 10 9 2 3 16 1 15 15 13 10 9 0 2 4 13 10 9 1 3 12 9 1 10 9 7 10 9 3 0 1 10 9 0 1 10 9 13 2
31 1 10 9 1 9 0 7 0 2 1 15 1 9 7 0 7 10 9 4 13 15 10 9 1 3 10 9 1 10 9 2
12 13 0 1 10 9 10 9 1 10 9 0 2
40 10 9 4 13 1 0 9 1 9 7 9 1 10 9 16 15 13 16 10 9 2 16 13 1 10 9 0 1 15 13 1 10 9 2 13 0 1 10 9 2
9 10 9 13 0 2 13 12 2 2
10 3 4 13 2 3 2 10 9 0 2
11 12 2 9 1 9 7 9 0 7 0 2
98 15 1 10 9 2 3 16 1 15 15 13 10 9 0 2 4 13 9 2 9 2 9 1 9 2 12 2 2 9 7 0 2 12 2 2 7 4 13 9 0 7 13 7 1 0 9 0 2 7 13 9 2 1 10 15 4 13 9 1 9 2 4 13 10 9 13 1 10 9 2 12 2 7 2 1 9 2 15 0 1 13 10 9 0 1 10 9 1 10 9 2 9 7 9 2 12 2 2
8 12 2 9 1 9 7 9 2
40 15 4 13 9 7 9 2 12 2 1 10 9 2 16 3 13 1 9 0 10 9 0 2 4 13 10 9 0 1 10 9 1 10 9 7 9 2 12 2 2
33 10 9 15 13 1 10 9 1 10 9 1 10 9 3 0 2 10 15 4 13 1 9 0 2 12 2 7 0 1 9 1 9 2
38 16 10 9 15 13 1 10 9 0 7 1 10 9 0 2 10 9 15 13 1 9 1 9 7 1 10 9 1 10 9 0 1 10 9 2 12 2 2
23 10 9 13 10 9 0 1 9 2 1 10 9 7 9 13 1 10 9 0 1 15 0 2
15 10 9 0 2 3 2 4 13 10 9 1 9 7 9 2
19 16 10 15 7 10 15 3 13 2 4 4 13 10 0 9 1 10 9 2
58 3 1 10 9 2 15 13 9 1 0 9 15 10 10 9 2 0 7 13 1 9 2 13 1 9 0 2 16 13 10 9 2 10 9 2 10 9 2 10 9 2 10 9 2 10 9 2 10 9 2 10 9 7 9 2 12 2 2
14 12 2 10 9 7 9 1 10 9 1 3 0 9 2
22 4 13 15 15 10 10 9 2 13 1 9 3 0 1 12 9 2 15 13 1 9 2
29 12 2 0 9 1 10 9 2 10 9 2 10 9 0 2 10 9 1 9 1 9 3 0 1 12 9 7 9 2
42 10 9 4 13 3 1 10 9 2 16 10 9 13 1 9 2 1 9 7 1 0 9 0 15 15 13 3 3 1 10 9 2 7 1 12 9 1 10 9 1 9 2
41 10 9 15 13 1 10 9 1 10 9 1 10 9 0 1 10 9 1 10 9 1 10 9 1 10 9 2 7 1 10 9 0 1 10 9 3 4 13 10 9 2
36 10 9 0 3 15 4 13 16 1 10 9 13 10 9 0 2 10 7 0 2 16 10 9 4 13 1 9 15 3 13 10 9 1 10 9 2
31 10 0 9 1 10 9 1 10 9 2 13 1 13 10 9 1 10 9 1 10 10 9 1 9 2 13 12 2 7 9 2
17 10 9 13 10 9 15 15 13 7 3 15 3 13 1 10 9 2
20 10 9 4 2 3 2 13 1 10 9 13 1 10 9 7 1 10 9 0 2
14 12 2 9 1 9 2 9 7 1 10 9 1 9 2
57 1 10 9 15 13 7 15 13 1 10 9 2 1 10 9 1 9 3 0 2 7 1 10 9 7 10 9 1 10 9 2 15 13 2 13 15 1 9 2 9 7 9 1 9 0 2 10 9 7 2 1 9 2 10 9 0 2
19 16 10 15 7 10 15 3 13 2 15 13 10 9 13 1 10 9 0 2
8 12 2 9 1 9 3 0 2
31 10 9 4 13 16 15 13 10 9 7 10 9 15 4 13 7 13 1 9 0 1 15 13 1 10 9 0 2 12 2 2
11 12 2 9 1 13 9 1 9 3 0 2
44 16 15 4 13 10 9 1 13 9 1 9 0 1 15 3 13 2 7 10 9 13 7 4 13 7 13 2 10 9 3 4 13 15 2 16 3 13 10 9 0 2 12 2 2
17 10 9 3 15 13 16 10 9 13 9 1 9 13 1 10 9 2
10 12 2 9 1 9 13 7 1 9 2
56 15 1 10 10 9 15 13 10 9 1 10 9 1 10 9 2 12 2 4 1 10 9 13 15 1 13 15 2 7 4 15 0 13 10 9 15 15 13 1 10 10 9 2 0 3 1 10 10 9 10 9 7 10 9 0 2
37 16 10 9 0 3 13 3 2 10 9 3 13 1 10 9 13 1 10 9 1 10 9 13 1 10 9 1 10 9 1 15 4 13 2 12 2 2
31 16 1 9 1 10 9 0 10 9 13 1 10 9 1 10 9 2 1 10 9 1 15 15 13 10 9 1 10 9 12 2
6 12 2 9 1 9 2
51 15 13 16 10 9 13 1 10 9 15 15 15 13 1 10 9 1 10 10 9 2 7 1 10 9 1 10 9 1 10 10 9 13 10 9 1 10 9 7 10 9 13 15 1 3 12 9 2 12 2 2
26 16 15 7 15 1 10 9 13 1 10 9 7 15 7 15 1 10 9 0 2 10 9 15 13 0 2
6 12 2 9 1 9 2
28 10 9 1 12 9 15 13 0 7 4 13 1 9 0 2 3 16 15 13 9 1 9 7 10 9 1 9 2
44 16 15 0 1 10 9 4 13 2 15 13 16 10 9 13 1 10 9 1 10 9 13 2 7 1 15 1 10 10 9 15 13 10 9 0 1 9 1 10 9 1 9 13 2
6 12 2 9 1 9 2
10 10 9 13 1 10 9 0 13 0 2
19 10 9 13 1 10 9 1 9 15 13 0 2 0 9 7 9 1 9 2
41 10 9 15 13 1 9 7 15 15 13 1 10 9 0 3 4 4 13 2 16 3 1 0 9 7 3 16 10 9 0 4 13 10 9 7 10 9 1 10 9 2
6 12 2 9 1 9 2
16 10 9 7 0 9 1 10 9 1 10 9 13 1 12 9 2
26 9 2 16 13 9 1 10 9 7 1 10 9 2 7 3 13 1 13 15 1 10 9 1 10 9 2
17 10 9 1 10 9 4 13 3 1 10 9 13 1 10 9 12 2
33 3 13 10 0 9 1 9 2 16 10 9 15 3 13 0 1 9 4 13 9 0 2 13 12 2 7 4 13 1 10 9 12 2
13 10 9 15 15 13 1 10 9 1 10 9 13 2
39 12 2 4 13 1 10 9 2 12 2 0 1 13 10 9 1 10 9 7 1 10 9 2 12 2 0 1 9 10 10 9 3 13 0 1 12 9 0 2
57 12 2 13 10 9 0 1 10 9 3 0 1 12 9 7 9 1 10 9 7 1 10 9 1 10 9 1 10 15 15 4 13 9 7 9 2 16 15 13 1 10 9 0 2 7 3 0 1 12 9 16 13 1 10 9 0 2
64 12 2 13 10 9 0 1 10 9 3 0 1 12 9 7 9 1 10 9 1 10 9 0 2 1 3 16 15 13 1 9 15 13 1 15 7 1 9 1 9 0 1 10 9 1 10 9 7 10 9 1 10 9 3 13 1 13 10 9 0 2 12 2 2
12 12 2 9 0 1 10 9 13 1 10 9 2
31 10 9 15 3 13 10 9 1 9 7 1 9 4 13 1 9 2 3 16 3 4 4 13 10 9 13 1 10 9 12 2
21 10 9 13 3 10 9 1 13 16 15 4 13 0 1 10 9 1 10 9 13 2
13 12 2 9 1 10 9 10 7 1 10 9 0 2
20 10 9 4 4 13 1 10 9 1 10 9 2 12 2 0 1 10 9 10 2
26 16 10 9 13 0 2 12 2 2 15 1 10 9 4 13 9 1 10 9 2 12 2 1 10 15 2
26 7 15 4 13 10 9 0 4 13 15 1 10 0 9 1 15 10 9 3 4 4 13 2 12 2 2
8 12 2 9 1 13 10 9 2
29 10 9 1 9 1 10 9 3 13 1 10 9 1 13 10 9 1 10 9 2 12 2 0 7 1 13 1 9 2
24 15 13 10 9 1 10 9 3 4 13 10 9 16 1 15 3 13 10 10 9 2 12 2 2
12 12 2 9 1 10 9 1 9 0 7 9 2
56 3 15 4 13 9 0 1 10 9 0 7 3 0 7 3 1 10 9 1 10 9 2 16 1 10 9 1 15 7 10 9 0 1 10 9 1 15 15 13 10 9 0 3 15 13 10 9 1 10 9 7 9 2 12 2 2
54 3 15 4 3 13 9 7 0 9 2 9 2 9 0 7 0 2 0 1 9 15 13 1 13 15 1 10 9 1 10 9 2 16 3 15 13 10 9 1 10 9 7 0 1 10 9 7 10 9 0 1 0 9 2
21 10 9 13 16 1 10 12 9 0 15 13 10 9 0 2 12 2 2 12 2 2
18 10 9 1 10 9 13 15 1 13 10 9 7 10 9 1 10 9 2
12 12 2 9 1 10 9 1 9 0 7 0 2
44 3 15 4 13 9 0 7 0 1 10 9 1 10 9 16 3 15 13 10 9 1 12 9 2 10 15 4 13 15 1 10 3 0 9 1 10 9 7 1 10 3 0 9 2
43 16 15 4 13 10 9 2 12 2 1 13 9 0 1 10 9 0 2 10 9 1 15 3 4 13 2 12 2 1 9 0 1 12 9 2 13 1 9 1 10 9 12 2
32 16 10 9 0 13 3 9 0 2 10 9 1 12 9 4 3 13 15 1 10 9 1 10 9 1 15 10 9 0 15 13 2
33 16 15 4 13 10 0 9 1 10 9 1 15 13 10 0 9 0 7 0 2 15 4 13 15 3 1 12 9 1 10 10 9 2
46 10 9 0 2 0 1 10 9 1 9 13 1 10 9 12 4 13 1 10 9 16 10 9 1 10 9 1 10 9 1 10 9 1 10 9 13 0 1 10 9 1 10 9 1 13 2
16 10 9 13 10 0 9 1 10 9 12 2 7 13 9 0 2
30 3 10 9 12 2 13 10 9 2 4 13 10 9 1 9 0 2 7 10 9 12 4 13 1 13 10 9 1 9 2
12 10 9 1 15 13 4 13 1 10 0 9 2
38 10 9 1 9 4 13 1 10 9 1 10 9 2 13 12 2 13 1 10 9 12 2 7 3 4 13 1 10 9 1 10 9 13 1 10 9 12 2
8 12 2 9 1 10 9 0 2
30 10 9 4 13 10 9 1 9 16 10 9 0 13 1 10 10 9 7 3 4 13 15 13 1 10 9 1 10 9 2
19 16 13 0 9 2 4 13 16 10 9 0 15 4 13 1 9 7 9 2
16 15 13 1 10 9 10 9 0 7 10 9 1 10 9 0 2
17 10 9 12 13 10 9 1 10 9 1 9 13 1 10 9 12 2
28 10 9 4 3 4 13 1 10 9 15 4 13 10 9 2 13 12 2 1 9 2 9 2 13 12 2 2 2
11 12 2 9 1 10 9 13 1 10 9 2
41 10 9 1 10 9 13 9 1 13 10 9 1 15 13 2 12 2 2 0 10 9 1 10 9 0 1 10 9 0 2 12 2 7 1 10 9 0 2 12 2 2
18 15 4 3 13 15 1 9 1 15 2 16 3 13 10 9 1 15 2
20 7 2 16 4 15 13 1 10 9 2 3 4 13 15 1 9 1 0 9 2
21 13 4 10 9 1 10 9 1 10 9 1 10 9 1 10 9 0 1 15 13 2
38 15 13 16 10 9 13 1 10 9 13 1 10 9 0 2 13 12 2 1 10 9 2 7 16 4 13 1 9 0 7 0 1 10 9 1 10 9 2
29 10 9 4 13 1 10 9 0 1 10 9 1 10 9 2 15 13 16 10 9 13 10 9 1 9 1 10 9 2
41 16 10 9 1 10 9 13 9 1 10 9 13 0 13 16 15 13 10 9 1 9 1 3 10 9 4 3 13 1 10 9 1 10 9 1 9 2 13 12 2 2
26 15 13 16 10 9 1 10 9 13 9 1 10 9 3 0 15 1 15 13 1 9 1 10 9 12 2
20 1 9 10 9 13 10 9 0 3 1 10 9 2 7 15 13 10 9 0 2
23 3 10 9 13 10 9 1 9 7 9 3 0 16 13 1 10 15 0 1 10 9 9 2
38 1 15 13 10 9 0 15 13 16 13 10 9 0 2 9 1 10 9 0 11 12 2 12 2 12 2 9 12 2 0 1 10 9 13 10 9 0 2
13 12 2 9 1 10 9 15 13 7 13 10 9 2
14 13 4 10 9 1 10 9 1 10 9 1 10 9 2
2 3 2
52 8 2 3 13 10 9 1 9 1 10 9 1 10 9 13 7 13 1 10 9 2 1 3 10 9 1 10 0 9 3 4 13 1 10 9 0 2 3 10 9 1 10 9 4 13 1 9 2 13 12 2 2
24 8 2 3 13 10 9 1 9 0 2 1 3 10 9 1 9 4 13 1 13 3 10 9 2
30 15 13 16 10 9 1 15 1 10 9 12 4 13 1 10 9 0 2 15 13 1 13 1 10 9 10 0 9 0 2
10 12 2 9 1 0 9 7 0 9 2
118 15 4 13 9 2 12 2 2 13 9 7 9 1 9 7 1 9 13 9 1 13 9 1 10 9 7 13 9 7 9 2 7 13 15 2 13 15 7 13 15 10 9 2 13 15 7 13 15 10 9 7 13 15 10 9 2 12 2 2 4 2 1 10 9 13 1 10 9 12 2 13 10 0 9 7 13 10 9 15 13 0 1 3 13 9 1 10 9 10 2 9 2 9 7 9 1 9 2 9 7 9 0 7 13 1 10 9 1 10 9 7 1 10 9 0 7 0 2
39 10 9 13 16 10 9 4 13 1 10 9 0 1 3 13 10 9 1 10 9 0 2 7 1 13 16 10 9 13 0 10 9 1 10 9 0 3 13 2
7 12 2 9 1 0 9 2
66 16 13 9 2 12 2 1 10 9 1 15 10 9 3 0 4 13 0 2 10 9 0 4 13 10 9 1 10 0 9 1 10 10 9 7 3 1 10 9 15 4 13 1 10 9 7 1 10 9 1 10 9 1 15 10 9 4 13 7 15 4 13 2 12 2 2
21 10 9 0 4 13 10 9 1 10 9 15 13 9 1 10 10 9 2 12 2 2
21 1 10 10 9 4 13 15 10 9 1 10 9 1 10 9 7 1 10 9 0 2
31 10 9 0 13 0 1 13 10 9 15 1 10 9 3 0 13 3 2 1 16 4 13 10 9 1 10 9 2 12 2 2
25 10 9 1 10 9 0 3 4 13 10 9 2 7 10 9 1 10 9 0 4 13 15 3 0 2
27 3 0 10 9 13 1 10 0 9 2 15 13 9 1 10 9 0 1 10 9 1 13 10 0 9 0 2
34 15 13 3 1 10 9 10 9 3 0 1 10 9 1 10 9 15 1 10 9 1 10 9 13 15 1 10 9 0 1 10 10 9 2
22 1 13 16 10 9 1 10 9 1 10 9 1 10 9 4 13 3 1 10 9 0 2
11 12 2 9 1 13 10 9 1 10 9 2
20 15 13 1 10 9 10 9 1 10 15 7 1 10 0 9 1 10 9 12 2
35 10 9 2 15 13 1 10 9 0 13 1 10 9 12 2 13 13 10 9 1 10 9 1 9 1 10 9 0 1 10 9 1 10 9 2
8 12 2 9 1 9 7 9 2
95 16 10 9 7 10 9 15 13 1 9 1 10 9 4 4 1 15 7 1 9 13 7 13 2 7 1 10 0 9 1 10 9 1 10 9 15 13 0 13 0 9 7 9 2 7 10 9 1 10 9 3 13 3 1 13 15 7 1 13 15 2 15 1 10 9 15 4 13 7 4 13 9 4 13 15 2 0 9 1 10 9 2 12 2 2 15 13 1 9 1 9 2 12 2 2
37 10 9 4 4 13 1 9 16 10 9 1 10 9 2 1 15 15 15 13 2 3 15 13 9 2 1 15 0 13 1 10 9 1 10 9 0 2
7 12 2 9 1 10 9 2
61 10 9 1 10 9 0 15 13 3 16 15 13 1 13 10 9 13 15 1 10 9 1 10 9 7 1 10 9 2 9 2 9 7 0 9 2 1 9 1 9 1 15 13 2 1 9 16 10 9 13 7 13 1 13 10 9 0 2 12 2 2
45 10 9 12 7 12 13 10 0 9 0 1 10 9 2 13 12 2 2 9 15 15 13 1 10 9 1 10 9 1 13 1 9 1 10 9 0 16 4 13 10 9 1 10 9 2
11 12 2 9 1 10 9 2 9 7 9 2
39 10 10 9 2 1 10 15 13 0 16 10 9 7 10 9 4 13 7 13 7 10 9 13 2 4 13 1 10 9 1 9 1 10 9 15 15 15 13 2
59 3 2 16 10 9 1 10 9 2 10 9 1 10 9 7 10 9 1 10 10 9 13 1 9 1 15 1 10 9 2 10 9 1 9 2 1 9 7 1 9 13 3 1 1 15 2 0 1 10 9 10 9 1 10 9 2 12 2 2
20 16 13 0 13 10 0 9 13 1 10 9 2 10 9 15 13 1 9 0 2
5 12 2 9 0 2
31 4 13 15 1 9 10 9 1 9 0 15 4 13 7 13 1 9 10 9 13 1 10 0 9 1 9 7 1 9 0 2
24 10 9 1 10 0 7 10 9 1 10 9 4 13 1 9 13 2 12 9 12 2 12 2 2
25 10 9 1 10 9 4 13 1 10 9 13 1 9 1 10 9 1 10 9 1 15 13 10 9 2
7 12 2 9 1 10 9 2
42 10 9 1 10 9 3 13 9 16 3 16 4 13 1 10 9 13 10 12 9 2 7 16 2 4 15 10 9 13 1 0 9 2 15 4 13 1 15 1 10 0 2
5 12 2 9 0 2
24 1 15 4 13 1 10 9 0 2 15 13 1 10 9 0 3 13 10 9 13 1 10 9 2
49 13 10 0 9 1 10 9 13 1 10 9 12 3 13 0 7 10 9 12 2 1 3 10 9 1 9 1 10 9 4 13 1 9 1 10 9 1 10 9 15 13 10 9 2 7 10 9 12 2
5 12 2 9 0 2
38 1 10 9 13 1 10 9 12 2 10 9 4 3 4 13 1 9 1 10 9 0 2 1 10 9 1 13 1 10 0 9 1 10 9 2 12 2 2
20 1 10 9 1 9 7 10 9 15 13 10 9 13 1 10 9 1 9 0 2
20 10 9 4 3 13 1 10 9 1 10 0 9 1 10 9 1 10 13 9 2
6 12 2 9 1 9 2
72 10 9 15 13 1 9 2 12 2 2 1 9 2 12 2 2 1 9 2 12 2 2 1 9 2 12 2 2 1 9 7 9 2 12 2 2 1 9 2 12 2 2 1 9 1 9 2 12 2 2 1 9 1 9 1 9 2 12 2 7 1 10 0 9 13 1 10 9 2 12 2 2
24 10 9 0 2 12 2 2 12 2 15 3 13 9 2 12 2 1 15 15 13 1 10 9 2
20 0 13 10 9 0 7 10 9 15 13 9 1 9 2 12 2 7 1 9 2
6 12 2 9 1 9 2
30 10 9 1 9 1 9 13 9 1 13 15 1 10 9 2 12 2 10 2 7 13 9 1 10 9 13 1 10 9 2
30 16 3 15 4 13 1 12 9 7 4 13 1 12 9 1 13 15 2 4 13 15 7 13 15 10 9 1 10 9 2
29 10 9 0 4 4 13 1 10 9 1 10 9 10 2 0 10 9 1 10 9 1 10 9 1 9 1 10 9 2
30 15 13 1 15 15 15 4 13 2 16 3 4 13 1 12 9 1 16 10 9 4 13 9 1 10 9 3 15 13 2
10 12 2 9 1 9 2 9 7 9 2
32 10 9 7 9 15 13 1 10 0 9 7 9 15 13 1 10 9 1 15 2 16 3 15 4 4 13 1 9 7 1 9 2
28 10 0 9 15 13 1 10 9 15 13 1 0 9 2 0 10 0 9 1 9 1 10 9 0 2 12 2 2
34 10 9 2 16 13 1 10 9 13 1 10 9 7 1 10 9 2 13 1 9 10 9 1 9 1 10 9 1 9 2 13 12 2 2
5 12 2 9 13 2
55 15 13 10 9 0 4 13 15 1 10 9 2 12 2 2 7 2 16 3 15 13 2 4 13 15 2 12 2 1 9 1 10 9 2 12 2 1 10 9 1 15 15 4 13 2 13 10 9 1 10 9 2 12 2 2
7 12 2 9 1 10 9 2
10 12 2 9 1 9 1 10 9 13 2
40 13 10 9 1 10 0 9 1 10 9 1 16 15 13 10 9 2 10 9 7 10 10 9 2 16 10 9 15 4 13 10 9 2 13 1 15 15 4 13 2
24 3 10 9 1 10 9 2 13 10 9 7 13 10 9 2 4 13 10 9 13 2 12 2 2
20 10 0 9 1 10 9 1 9 13 3 1 13 10 9 15 4 13 10 9 2
13 1 9 4 3 13 10 9 1 10 9 1 9 2
40 15 13 16 15 13 1 10 9 1 9 2 13 12 2 2 10 10 9 0 15 13 3 16 4 13 10 9 1 10 9 2 16 3 10 9 15 13 8 8 2
16 1 15 10 9 13 9 1 10 9 0 0 13 1 12 9 2
8 12 2 9 13 1 10 9 2
34 10 9 4 13 1 9 1 9 2 12 2 1 10 9 2 16 15 15 13 2 10 9 1 10 9 7 1 10 9 1 10 9 13 2
24 16 10 9 7 9 13 10 12 2 12 2 9 2 10 9 1 10 9 13 3 1 10 15 2
27 16 10 9 3 13 9 0 2 12 2 2 10 9 1 10 9 4 13 1 10 9 1 10 10 0 9 2
12 12 2 9 1 10 9 7 9 1 10 9 2
30 1 10 9 1 10 9 0 1 10 9 12 7 0 2 1 10 9 4 13 2 1 10 9 2 10 9 7 10 9 2
33 1 13 15 4 13 10 9 2 10 9 13 16 15 4 13 15 3 1 15 15 4 13 1 4 13 16 15 13 7 3 10 9 2
24 9 13 10 9 0 1 9 2 12 2 2 13 7 13 2 1 15 15 4 13 1 13 9 2
17 10 9 13 1 10 9 1 10 9 2 12 2 1 15 15 13 2
43 16 10 9 4 13 1 10 9 10 2 16 4 4 13 1 0 9 1 10 9 2 12 2 2 13 1 9 1 10 9 1 10 9 7 1 9 1 10 9 2 12 2 2
19 10 0 9 15 13 16 10 9 4 13 1 10 9 0 10 2 12 2 2
32 1 10 9 1 10 9 1 9 0 2 0 2 0 2 0 7 0 15 13 10 9 1 10 9 0 2 12 2 2 12 2 2
10 12 2 9 13 1 7 1 10 9 2
52 10 9 2 9 7 9 13 1 7 1 10 9 13 1 10 9 1 15 2 1 15 4 13 1 10 9 12 2 12 2 12 7 12 7 3 16 13 3 1 10 9 2 12 2 7 1 10 9 2 12 2 2
28 1 10 9 4 13 10 9 1 10 9 2 9 2 9 7 10 9 2 1 10 9 0 1 9 7 10 9 2
31 1 10 9 13 10 9 15 4 13 9 0 7 10 15 15 15 13 1 15 4 13 9 1 10 9 0 2 8 8 2 2
14 12 2 9 13 1 10 9 1 10 9 1 9 10 2
57 10 9 1 10 9 15 4 13 9 2 9 7 9 1 9 10 4 13 15 10 9 2 16 10 9 3 4 13 1 10 9 1 10 9 2 7 3 4 13 15 1 16 15 13 0 9 1 10 9 13 7 1 16 13 10 9 2
28 13 3 2 3 1 10 9 16 15 13 10 9 2 10 9 1 10 9 2 16 13 1 9 0 2 12 2 2
31 1 10 9 10 9 1 10 9 3 4 13 13 12 9 2 12 2 1 10 9 1 15 10 9 4 13 9 1 10 9 2
35 10 0 9 13 1 10 9 12 13 1 13 16 10 0 9 1 10 9 1 10 15 9 1 10 9 13 2 13 1 10 9 1 10 9 2
11 12 2 9 13 1 10 15 1 9 10 2
42 16 10 9 2 9 7 9 4 4 13 1 10 15 2 12 2 1 10 9 2 10 9 1 10 9 13 9 1 13 15 7 1 13 15 15 15 4 13 1 13 15 2
39 16 10 9 13 1 13 15 2 4 13 1 10 9 10 9 1 10 9 7 10 9 1 10 9 1 9 7 10 9 1 9 13 1 10 9 2 12 2 2
24 16 10 9 1 10 9 13 16 4 13 2 15 4 13 15 1 9 1 15 15 15 4 13 2
12 15 4 3 4 13 1 10 9 1 10 9 2
41 10 9 3 4 13 10 15 1 13 10 9 2 9 7 9 2 16 4 4 13 1 10 9 7 1 9 7 16 4 4 13 1 10 15 1 0 9 2 12 2 2
26 10 9 3 4 4 13 13 12 9 2 12 2 1 10 9 1 15 10 9 4 13 9 1 10 9 2
16 10 9 13 1 10 9 13 1 13 10 9 0 1 10 9 2
27 1 9 15 4 13 16 1 10 9 13 9 0 3 0 1 10 9 1 10 9 2 1 9 1 10 15 2
22 10 9 2 3 2 15 13 1 10 9 15 13 10 0 9 2 13 12 2 12 2 2
11 12 2 9 13 1 10 15 1 9 10 2
51 16 10 9 2 9 7 0 9 4 4 13 1 10 15 1 9 10 2 10 9 1 15 4 13 15 2 0 9 1 9 1 10 15 2 16 10 9 4 13 15 1 0 9 1 10 9 7 1 10 9 2
25 10 9 3 4 13 13 12 9 1 10 9 1 15 10 9 4 13 9 1 10 9 2 12 2 2
59 1 10 9 16 10 9 1 10 9 3 4 13 7 16 10 9 13 0 2 10 0 15 15 4 13 9 7 10 9 1 10 9 15 4 13 1 9 2 12 2 4 13 1 9 1 10 9 1 10 9 0 1 10 9 1 10 9 0 2
33 10 9 1 10 9 4 3 13 10 9 1 10 9 1 10 9 2 3 1 0 9 2 3 1 10 9 15 1 15 4 3 13 2
47 4 3 13 10 9 1 10 9 2 3 1 10 9 1 10 15 15 15 4 13 9 1 10 10 9 2 7 1 10 9 1 10 9 1 10 9 15 1 9 4 13 10 9 2 12 2 2
9 12 2 9 1 9 1 9 0 2
78 16 1 10 9 1 10 9 15 13 1 0 9 2 12 2 10 9 2 12 2 1 10 9 0 2 7 10 9 1 15 3 13 9 1 12 9 2 12 2 1 10 9 1 15 13 9 10 9 2 10 9 0 2 13 9 1 10 9 2 4 13 1 10 9 10 9 1 10 9 7 1 10 9 13 2 12 2 2
32 10 9 4 13 1 13 1 10 9 1 10 9 10 9 1 10 9 1 10 9 13 2 1 10 9 1 10 9 2 12 2 2
8 10 9 13 10 0 9 0 2
37 16 1 10 9 1 9 13 10 9 1 10 9 16 13 9 1 10 15 15 15 13 1 15 2 1 10 9 1 10 9 0 15 13 10 9 0 2
21 1 13 16 10 9 15 13 3 7 3 16 10 9 1 9 4 13 1 10 9 2
17 10 9 0 13 3 10 9 1 9 3 3 0 3 1 10 9 2
13 10 9 1 10 0 9 1 10 9 13 3 0 2
27 10 9 12 13 10 9 1 9 1 10 9 2 10 10 9 0 4 13 1 10 9 0 2 13 12 2 2
6 12 2 9 7 9 2
50 16 10 9 13 1 10 9 4 4 13 2 12 2 7 13 2 12 2 1 9 1 13 10 0 15 2 7 13 0 1 0 9 2 15 13 10 9 1 10 9 10 7 13 9 1 13 15 10 9 2
24 1 9 0 2 10 9 15 13 0 1 9 1 10 9 1 10 9 13 1 15 2 12 2 2
46 16 3 15 1 10 9 15 4 13 1 0 7 13 1 3 0 1 9 2 12 2 2 16 13 1 10 15 1 9 2 12 2 2 10 9 1 10 9 0 13 10 9 1 10 9 2
51 7 16 10 9 7 10 9 4 13 1 10 10 9 1 9 1 10 9 1 10 9 0 2 15 3 4 13 1 13 16 10 9 0 1 10 9 1 9 13 1 10 9 0 7 10 9 1 10 9 0 2
17 4 3 13 10 9 1 10 9 1 9 1 9 0 2 12 2 2
22 10 0 9 1 10 9 13 10 9 2 13 12 2 1 10 9 0 1 0 9 0 2
36 13 1 13 0 16 16 10 9 7 10 9 13 1 9 1 10 9 7 1 9 1 15 13 1 13 15 10 9 0 2 15 13 10 9 12 2
30 3 1 15 13 1 10 9 12 2 3 15 13 9 1 9 16 13 10 9 15 13 10 9 1 10 9 1 10 9 2
24 4 13 0 3 3 10 9 15 13 10 9 0 0 2 7 3 15 15 13 10 9 0 0 2
61 16 15 4 13 10 9 15 3 15 13 1 13 10 0 9 2 12 2 2 4 7 3 4 10 9 13 10 10 0 9 2 15 13 10 9 13 1 10 9 10 9 1 10 9 2 3 16 10 9 1 10 9 13 3 15 1 10 9 1 9 2
26 1 10 0 9 10 9 13 1 10 9 1 10 9 2 10 15 4 13 10 9 1 10 9 1 9 2
41 10 9 12 13 10 9 1 9 1 10 9 0 3 1 15 13 1 10 9 0 2 7 1 10 9 3 4 13 10 9 1 12 9 7 10 9 1 9 7 9 2
55 16 1 10 0 9 10 9 4 1 9 13 1 9 1 10 9 1 10 9 2 10 9 12 2 3 2 13 10 9 13 1 9 0 10 9 1 10 9 2 3 16 15 13 10 9 0 0 1 13 1 15 10 9 13 2
47 10 9 1 9 7 10 9 2 15 15 13 3 7 3 2 12 2 1 10 9 13 1 10 9 1 10 9 7 9 2 13 1 10 9 1 10 9 2 1 15 4 13 1 10 9 0 2
9 12 2 9 13 1 10 9 0 2
49 2 12 2 10 9 13 1 10 9 0 2 15 3 2 12 2 15 13 1 15 1 10 9 13 15 1 10 15 2 13 1 10 9 0 2 1 16 10 9 1 10 9 0 4 13 10 9 13 2
30 1 10 9 1 10 0 9 2 15 13 1 9 0 10 9 2 10 9 7 10 0 9 13 0 1 10 9 1 9 2
33 15 13 1 10 0 9 13 3 1 10 9 13 1 10 9 2 1 10 9 2 1 10 9 7 1 10 9 13 1 10 9 0 2
6 12 2 9 7 9 2
44 10 9 15 10 9 13 16 15 13 1 10 9 1 10 9 1 10 9 7 1 10 9 13 1 10 9 1 10 9 7 1 10 9 2 16 10 9 1 10 9 13 1 13 2
23 10 9 3 13 10 9 1 10 9 1 10 9 15 10 9 13 1 10 9 1 9 0 2
51 9 7 9 15 13 1 10 9 13 1 10 9 12 7 0 2 16 10 9 1 10 9 7 1 10 9 13 9 3 1 10 9 13 1 10 9 7 10 0 9 1 10 9 3 4 13 1 10 9 13 2
57 16 10 9 7 9 13 1 9 0 2 12 2 10 9 0 7 0 1 10 9 0 1 10 10 9 7 15 13 1 10 9 0 7 1 10 0 9 2 10 9 1 10 9 1 10 15 15 4 13 10 9 13 15 13 10 9 2
24 4 3 13 1 10 0 9 10 9 1 10 9 1 10 0 9 13 1 10 9 1 10 9 2
8 12 2 9 7 9 1 9 2
53 10 9 7 9 1 9 15 15 13 1 10 9 1 10 9 7 9 13 1 10 9 0 2 16 10 9 15 4 13 1 9 2 12 2 2 10 9 1 10 9 2 1 15 4 13 10 9 2 15 13 10 9 2
41 10 0 9 15 13 16 10 9 7 10 9 2 13 10 0 9 2 13 7 13 10 9 7 9 1 10 9 1 10 9 13 2 13 15 10 9 2 2 12 2 2
8 12 2 9 0 2 12 2 2
30 16 10 9 7 10 9 15 13 10 0 9 2 13 10 0 2 10 9 0 13 13 1 10 9 0 1 10 9 0 2
43 10 9 1 10 9 12 2 12 7 12 15 13 1 10 9 3 13 7 1 9 1 9 0 7 1 9 0 13 1 10 9 0 3 13 3 10 9 0 1 9 1 9 2
19 1 10 9 4 13 10 9 0 1 10 9 1 10 9 0 2 12 2 2
6 12 2 9 1 9 2
48 10 9 2 12 2 4 13 10 9 1 15 15 13 7 13 7 4 13 10 9 1 10 9 3 16 15 2 1 10 9 2 4 13 2 1 9 10 2 1 13 7 13 10 9 2 12 2 2
39 1 10 9 10 9 4 13 1 13 15 1 10 9 1 10 9 2 7 2 1 9 2 1 13 15 15 10 9 2 3 1 13 15 10 9 2 12 2 2
36 10 9 2 16 13 3 1 10 0 9 7 9 10 9 1 10 9 2 4 13 1 13 1 10 0 9 7 9 10 9 13 1 9 1 15 2
24 10 9 1 9 3 15 13 2 0 10 9 1 10 9 1 10 9 1 9 1 15 1 9 2
57 3 3 4 3 13 1 10 9 0 2 15 13 16 10 9 4 3 13 10 0 9 1 9 1 10 9 2 1 10 15 13 3 1 13 13 1 10 9 10 10 9 2 1 13 1 10 9 3 10 9 1 10 9 1 10 9 2
5 12 2 9 0 2
29 10 9 4 13 1 13 13 10 9 1 9 13 1 15 1 10 9 2 16 13 9 1 13 15 9 2 12 2 2
32 16 13 3 9 7 9 2 10 9 4 13 16 15 15 13 10 9 2 1 10 9 1 10 9 1 10 9 2 9 12 2 2
8 12 2 9 1 9 1 9 2
23 16 10 9 1 12 9 13 0 2 15 1 10 9 2 12 2 4 13 16 4 13 3 2
7 10 9 1 9 4 13 2
22 1 9 1 0 9 2 10 9 15 13 1 10 9 13 1 10 9 0 2 12 2 2
8 12 2 9 1 9 1 9 2
33 16 10 9 1 9 0 13 7 4 13 0 2 12 2 2 15 1 10 9 13 9 1 13 16 15 4 13 7 13 1 9 0 2
9 12 2 9 1 10 9 1 9 2
55 13 3 10 9 13 1 9 0 2 9 2 9 7 9 2 2 10 9 1 9 13 10 9 1 10 9 0 1 10 9 0 2 13 12 2 2 1 10 15 10 15 15 13 1 10 9 13 1 10 9 1 10 9 0 2
32 1 0 9 2 9 7 9 0 1 10 9 1 9 13 15 1 13 10 13 15 1 10 9 1 9 1 9 1 10 8 8 2
51 1 9 1 10 10 9 2 10 9 4 13 10 9 1 9 0 2 13 12 0 2 3 1 2 16 13 10 9 1 10 9 2 13 12 0 2 2 3 10 9 1 9 1 10 9 2 13 12 0 2 2
67 15 13 2 3 2 16 10 9 8 8 2 1 15 13 10 9 1 13 7 13 10 9 1 10 1 3 1 10 9 10 2 4 2 1 10 9 2 13 10 9 0 1 10 9 0 7 13 10 9 1 10 9 0 1 9 1 9 0 0 1 10 0 9 1 10 13 2
31 1 13 16 15 15 13 3 1 10 9 1 9 7 1 10 9 0 1 9 2 13 13 9 1 10 0 9 1 10 9 2
7 12 2 9 1 9 0 2
27 10 9 1 10 9 1 9 1 9 1 10 9 2 12 2 13 10 9 1 10 9 0 13 1 10 9 2
29 10 9 13 1 10 9 15 13 1 10 9 2 0 2 1 10 9 2 10 9 1 10 0 9 1 10 9 12 2
29 10 9 1 9 2 15 13 1 9 10 9 2 3 13 2 16 3 1 10 9 1 9 1 10 9 1 10 9 2
34 10 9 1 13 10 9 1 10 9 10 15 13 1 9 1 9 1 10 3 9 13 1 12 9 2 12 2 2 12 2 2 12 2 2
10 12 2 9 1 10 3 1 10 9 2
31 10 9 0 15 13 3 1 10 9 1 15 4 13 10 9 1 13 7 13 9 1 10 3 1 10 9 10 2 12 2 2
10 12 2 9 1 9 0 1 10 9 2
25 3 4 4 13 7 13 10 9 1 10 9 3 1 10 9 1 10 9 2 12 2 2 12 2 2
5 12 2 9 0 2
24 10 9 2 3 16 10 9 13 3 2 4 13 1 10 9 13 1 10 9 0 2 12 2 2
43 10 9 2 12 2 12 2 12 2 3 4 3 13 1 10 9 0 1 10 9 12 2 0 9 2 12 2 0 9 2 12 2 12 2 12 2 12 7 12 2 12 2 2
13 13 10 9 13 16 4 13 1 10 0 9 0 2
32 15 13 1 10 9 10 9 1 9 0 2 1 10 9 1 10 9 1 0 9 2 7 9 0 2 3 13 1 10 9 2 2
12 10 9 4 13 0 7 1 9 2 12 2 2
16 10 9 0 3 4 4 13 1 10 9 0 1 10 12 9 2
7 12 2 9 1 10 9 2
49 10 9 13 10 0 9 15 13 10 9 1 10 9 1 10 9 2 12 7 0 2 2 1 10 9 2 12 2 7 3 1 10 9 1 10 9 1 9 1 10 9 1 10 9 0 2 12 2 2
22 10 9 1 10 9 15 13 1 10 9 2 12 7 0 2 12 7 0 2 12 2 2
7 12 2 9 1 10 9 2
19 10 9 13 10 9 1 13 10 9 7 1 13 1 10 13 10 9 0 2
17 15 4 13 1 10 9 1 9 7 1 10 9 0 1 9 0 2
23 10 9 3 4 13 9 7 9 1 10 9 1 10 0 9 1 10 9 7 9 1 9 2
7 12 2 9 1 10 9 2
36 10 9 1 10 9 1 10 9 2 12 2 12 2 13 3 2 12 7 0 2 1 10 10 9 7 1 10 9 1 10 9 16 13 10 9 2
40 1 10 9 1 15 13 10 9 7 10 9 4 13 3 1 10 9 7 1 10 9 2 15 13 1 10 9 0 1 10 9 3 1 10 9 1 10 10 9 2
10 12 2 9 1 10 9 2 13 2 2
10 12 2 9 0 7 0 1 10 9 2
12 16 10 9 0 13 3 2 10 9 15 13 2
69 16 4 13 10 9 0 1 10 9 7 10 9 13 0 1 10 9 1 10 9 0 2 10 9 2 1 10 9 2 4 13 10 0 9 1 10 9 2 7 13 1 10 10 9 2 13 10 9 1 10 13 2 0 10 9 1 10 9 1 10 9 1 10 9 0 2 12 2 2
38 16 10 9 4 13 7 10 9 4 13 3 1 10 9 1 10 13 2 10 9 4 13 1 10 13 7 10 9 1 9 1 10 9 1 10 0 9 2
23 1 10 9 1 9 1 0 9 2 12 2 2 10 9 15 13 1 9 1 10 9 0 2
7 12 2 9 7 0 9 2
26 10 9 7 10 0 9 15 13 1 10 9 13 1 9 1 10 9 2 0 10 9 1 10 9 0 2
25 16 1 9 1 10 9 0 13 1 9 1 10 13 2 10 9 3 4 13 10 9 1 10 9 2
10 12 2 9 1 10 9 1 10 9 2
38 10 9 4 13 1 10 10 9 2 7 1 9 1 9 2 12 9 12 2 12 9 12 2 12 2 2 7 1 9 1 0 9 2 12 2 12 2 2
22 1 10 9 1 10 9 1 10 9 3 4 13 10 9 1 10 13 2 9 12 2 2
40 1 10 9 0 4 4 13 1 10 9 1 13 1 9 1 9 2 1 15 7 1 9 2 1 10 10 9 2 1 10 9 3 0 1 12 9 2 12 2 2
40 1 10 9 1 9 13 1 10 9 2 10 9 3 4 13 1 10 10 9 2 12 2 1 10 13 7 4 13 1 15 3 2 12 7 0 2 1 10 9 2
12 12 2 9 1 9 1 10 13 2 13 2 2
17 12 2 9 7 9 1 10 9 7 1 10 13 1 9 1 9 2
28 1 9 1 9 2 10 0 9 4 13 3 2 12 7 0 2 1 10 0 1 10 9 1 10 9 3 13 2
24 10 0 9 3 4 13 1 10 10 9 2 3 16 4 4 13 10 9 1 9 1 10 13 2
37 1 9 1 9 1 10 9 1 10 13 2 10 9 3 4 13 10 9 1 10 9 1 10 9 3 16 1 15 4 4 13 10 9 2 12 2 2
6 10 9 3 4 13 2
34 10 13 4 13 10 9 1 10 10 9 1 15 15 13 1 10 9 1 10 9 0 10 9 3 1 10 9 1 10 9 2 12 2 2
15 1 9 1 9 3 4 13 10 9 2 12 2 12 2 2
12 10 9 1 10 9 13 1 9 1 10 13 2
10 12 2 9 1 10 9 1 10 9 2
23 16 15 13 10 9 2 10 9 4 13 15 3 1 15 0 1 15 2 7 1 10 9 2
34 1 10 9 10 13 13 2 12 2 1 10 9 1 10 13 1 10 0 9 2 0 2 1 9 1 15 2 10 9 0 1 10 9 2
20 16 15 13 10 13 2 10 9 4 13 15 1 10 9 15 13 1 10 13 2
32 10 9 15 13 1 10 9 1 10 9 2 12 2 13 1 10 9 1 10 9 0 1 10 9 1 10 9 0 2 12 2 2
12 10 9 4 13 1 9 0 2 9 12 2 2
17 10 9 4 13 10 9 1 10 9 0 2 12 2 9 12 2 2
18 12 2 16 10 9 13 10 9 7 3 13 1 10 9 1 13 15 2
20 12 2 16 10 9 13 1 9 1 10 9 1 12 9 1 9 2 12 2 2
43 10 9 3 13 9 16 10 9 4 13 10 9 1 10 9 13 3 16 4 13 1 10 9 9 2 12 2 2 3 1 0 9 2 15 4 13 10 9 2 9 12 2 2
25 10 9 1 9 3 13 1 10 9 10 9 1 13 2 3 16 13 10 9 13 1 10 9 12 2
6 12 2 9 0 0 2
26 10 9 1 10 13 1 13 15 1 10 9 0 0 2 12 2 3 13 10 9 1 10 9 1 9 2
10 12 2 9 1 10 9 1 10 9 2
38 10 9 1 10 9 4 13 1 10 9 1 9 1 13 10 10 9 2 12 2 2 13 15 1 10 9 3 1 10 9 1 9 15 13 1 10 9 2
21 4 13 10 9 1 10 9 7 13 9 2 12 2 1 10 9 2 9 12 2 2
52 10 9 2 15 4 13 9 1 10 9 3 1 10 9 1 10 9 1 9 7 1 10 15 15 3 4 4 13 1 9 0 1 4 13 2 13 10 9 1 9 3 1 13 10 9 2 12 2 9 12 2 2
6 12 2 9 7 9 2
42 16 13 10 9 1 10 9 13 10 9 1 10 9 1 10 9 1 10 9 1 9 13 1 10 9 1 9 1 10 9 0 2 15 4 13 1 10 9 1 10 9 2
36 16 1 9 4 4 13 10 9 1 10 9 1 9 1 10 9 2 1 10 9 13 10 9 1 10 9 3 1 16 3 4 13 10 10 9 2
38 1 10 9 13 1 10 9 2 16 4 4 13 1 9 1 10 9 2 10 13 2 16 4 13 15 2 4 13 15 10 9 1 10 9 1 10 9 2
28 16 10 9 3 13 0 1 9 7 13 9 2 15 13 10 9 1 10 0 9 1 10 9 2 9 12 2 2
8 12 2 9 13 1 10 9 2
16 1 10 9 13 1 10 9 15 13 10 9 1 10 9 12 2
29 10 9 13 1 10 9 0 15 13 3 1 10 9 13 1 10 9 0 2 3 16 4 13 3 1 10 9 0 2
12 1 10 9 2 1 10 9 7 1 10 9 2
4 1 10 9 2
3 9 0 2
41 10 9 4 13 1 10 9 2 12 2 12 7 0 2 12 2 12 2 7 1 10 9 1 10 9 2 12 2 12 9 12 2 12 2 12 9 12 2 12 2 2
12 4 3 13 15 1 9 2 12 7 0 2 2
25 10 9 1 10 9 3 4 13 10 9 1 10 9 2 12 2 12 2 12 2 12 2 12 2 2
22 10 9 13 1 9 1 10 9 0 3 4 13 15 1 12 9 2 12 2 12 2 2
7 12 2 9 1 10 9 2
41 10 9 4 13 10 10 9 1 10 0 9 7 1 10 10 10 9 2 16 15 3 4 13 1 10 9 0 2 12 2 12 9 12 2 12 9 12 2 12 2 2
9 10 9 4 4 13 1 10 9 2
21 16 3 4 4 13 2 10 9 4 3 13 1 10 9 1 10 9 2 12 2 2
3 9 0 2
8 1 10 9 13 1 10 9 2
9 12 2 9 1 10 9 1 9 2
18 10 9 13 9 1 13 1 10 9 2 7 4 13 15 10 9 0 2
7 12 2 9 1 10 9 2
21 10 9 15 13 1 10 10 9 1 10 9 2 12 7 0 2 12 7 0 2 2
42 16 10 9 1 10 9 1 10 9 2 1 10 9 1 10 9 2 4 13 1 10 9 9 7 9 2 10 9 4 13 1 13 10 9 2 12 2 1 10 9 13 2
24 10 9 15 13 3 1 10 9 1 15 10 9 7 9 4 4 13 1 9 1 10 0 9 2
23 10 9 0 7 10 9 0 13 1 10 9 1 10 9 1 10 10 9 2 12 0 2 2
64 16 10 9 7 10 9 15 13 1 10 9 1 10 9 1 10 9 0 7 1 10 9 1 10 9 0 1 0 9 2 10 9 1 10 10 9 15 13 1 10 15 7 10 15 1 9 1 10 9 1 10 0 9 1 10 9 0 2 12 2 9 12 2 2
40 10 9 1 10 9 7 10 9 13 1 9 1 10 9 7 1 10 9 1 10 9 13 1 10 9 0 7 1 10 9 1 10 9 1 10 9 2 12 2 2
30 10 9 15 4 13 1 10 0 9 1 10 9 1 10 9 7 10 9 1 9 13 1 10 9 1 9 1 10 9 2
42 10 9 0 2 13 9 1 10 9 2 4 13 16 10 9 1 10 9 13 1 10 9 0 4 13 3 2 13 1 10 9 0 9 2 12 2 9 9 0 12 2 2
15 10 9 4 13 9 15 3 13 10 9 0 1 10 9 2
34 15 13 9 1 13 15 1 10 9 1 10 9 2 16 15 4 13 15 1 9 1 10 9 2 3 16 10 9 13 13 10 9 0 2
35 1 10 9 4 4 13 1 10 9 10 9 0 1 10 0 9 1 10 9 1 10 9 7 10 9 1 10 9 1 10 9 1 10 9 2
23 10 9 13 1 10 9 7 9 2 12 2 3 0 7 1 9 1 10 9 1 10 9 2
14 3 13 9 1 13 15 15 1 10 9 1 10 9 2
34 1 10 9 7 10 9 0 2 1 15 4 13 10 9 2 10 9 4 13 10 9 1 10 9 15 4 13 1 10 9 1 10 9 2
33 16 10 9 4 4 13 1 10 9 7 1 10 15 2 15 13 1 10 9 10 9 13 1 10 13 9 1 10 9 1 10 9 2
31 10 9 1 10 9 3 15 13 1 10 9 15 15 13 1 10 9 2 0 10 9 15 15 4 13 1 9 2 12 2 2
12 12 2 9 2 9 7 9 13 1 0 9 2
58 16 1 10 9 4 13 9 7 9 0 7 9 7 9 1 0 9 13 1 10 9 1 9 2 10 9 4 13 1 10 9 0 2 13 10 9 1 10 0 9 1 10 9 7 1 10 9 7 13 2 16 13 2 1 10 10 9 2
43 1 10 9 2 10 9 2 10 9 7 10 9 1 10 9 2 10 9 4 13 1 13 15 2 3 16 1 10 9 7 1 10 9 0 2 1 10 9 0 1 10 9 2
21 10 0 9 15 13 1 10 9 1 0 9 13 1 10 9 2 13 1 4 13 2
12 12 2 9 1 0 9 13 2 13 7 13 2
17 10 9 1 0 9 13 2 13 7 13 1 9 13 1 10 9 2
5 12 2 9 0 2
27 10 9 0 15 13 7 15 13 7 13 1 9 13 1 10 9 2 7 15 13 10 9 1 13 15 15 2
10 12 2 9 1 9 7 1 0 9 2
31 10 9 4 13 1 10 9 10 9 13 1 10 9 7 1 10 0 9 15 15 13 2 13 3 10 9 0 1 10 9 2
38 10 9 4 13 15 1 10 9 1 10 9 2 7 4 13 10 9 0 1 10 9 1 10 9 7 10 9 1 10 9 7 1 10 9 1 10 9 2
11 12 2 9 1 10 9 7 1 10 9 2
48 16 10 9 4 13 1 10 9 7 10 9 2 10 9 4 13 1 13 10 9 13 2 1 1 10 13 9 1 10 0 2 3 16 10 9 7 10 9 4 13 1 13 13 1 10 9 0 2
36 16 10 9 7 10 9 13 3 1 9 3 0 1 10 9 2 15 3 4 13 1 10 9 16 1 13 9 1 10 9 7 1 10 10 9 2
5 12 2 9 0 2
38 16 10 9 13 9 0 2 12 2 2 10 9 13 9 1 13 15 15 7 13 10 9 1 13 15 10 9 1 10 9 1 10 9 1 10 9 13 2
41 13 10 9 2 13 1 9 1 10 9 1 13 10 9 1 10 9 15 13 1 10 9 1 15 13 10 9 7 1 13 15 15 1 0 9 7 9 2 12 2 2
5 12 2 9 0 2
59 16 10 9 13 9 15 2 1 13 15 1 10 9 2 15 13 1 3 1 3 2 10 9 13 9 1 13 15 15 1 10 9 1 10 15 4 13 2 7 1 10 9 1 10 9 4 3 13 1 13 15 1 10 9 1 15 15 13 2
8 12 2 9 2 9 7 9 2
45 16 10 9 13 9 2 9 7 9 15 13 10 9 0 2 10 9 4 13 1 13 7 1 13 1 10 9 10 9 15 15 13 2 1 9 1 13 10 0 9 1 10 9 0 2
39 16 10 9 4 13 9 15 13 15 1 10 0 9 2 12 2 2 10 9 2 1 10 9 1 10 9 2 4 13 1 13 15 10 0 9 2 12 2 2
7 12 2 9 0 7 0 2
17 10 9 0 7 0 1 10 9 4 4 13 1 0 9 7 9 2
24 10 9 7 10 9 1 15 4 4 13 1 9 2 1 10 10 9 1 10 9 1 10 9 2
8 12 2 9 13 1 10 9 2
60 10 9 13 1 10 9 2 1 9 1 10 9 1 10 9 1 10 9 2 16 13 1 9 0 2 12 2 7 1 9 0 1 9 0 2 12 2 0 2 13 1 10 9 13 2 12 2 2 7 3 1 10 9 1 10 9 1 10 9 2
70 16 10 9 1 10 9 13 1 10 9 1 10 9 13 2 10 9 3 13 1 10 9 16 3 1 10 9 7 2 13 15 1 9 0 1 10 15 10 0 9 13 0 7 0 2 16 3 1 10 9 7 9 15 15 13 1 9 1 10 9 1 15 13 10 9 2 9 12 2 2
6 12 2 9 1 9 2
31 1 10 9 1 9 15 13 10 9 13 1 9 2 12 2 2 13 0 10 9 1 10 9 1 10 9 7 1 10 9 2
34 10 9 13 1 15 0 1 15 3 13 0 1 10 15 2 0 1 10 9 10 9 0 1 10 9 1 10 9 2 12 7 0 2 2
18 10 9 13 4 4 13 1 9 0 7 1 1 15 15 13 10 9 2
21 16 10 9 3 13 1 9 1 10 9 1 9 2 13 10 9 0 2 12 2 2
3 9 0 2
8 1 10 9 13 1 10 9 2
6 12 2 9 1 9 2
5 9 1 10 9 2
21 1 10 9 1 10 9 15 4 13 10 9 1 10 0 9 1 9 2 12 2 2
6 12 2 9 7 9 2
16 10 9 13 10 9 1 10 9 1 15 15 13 2 12 2 2
26 15 4 13 1 13 1 10 9 10 9 1 10 9 2 0 9 1 10 9 2 9 9 0 12 2 2
22 16 10 9 4 13 1 10 13 10 9 2 15 4 4 13 1 10 9 1 10 9 2
27 1 10 9 1 10 9 4 13 10 9 15 13 10 9 0 1 10 9 1 10 10 9 0 2 12 2 2
16 4 3 13 10 9 7 10 13 1 9 1 9 2 12 2 2
16 7 2 16 15 13 10 9 2 10 9 4 13 1 13 9 2
22 10 9 3 4 13 10 9 1 10 9 2 12 2 3 1 4 13 10 9 3 13 2
9 12 2 9 7 9 1 10 9 2
18 16 10 9 3 13 10 9 1 15 4 13 2 15 13 10 9 0 2
29 10 9 4 13 7 13 1 9 2 0 10 9 1 10 9 1 13 15 13 1 10 9 10 9 13 1 10 9 2
46 10 9 4 13 2 1 10 9 1 10 9 2 1 10 9 7 3 1 10 15 13 1 0 9 1 9 7 9 7 2 1 9 1 10 9 2 13 1 10 9 0 2 9 12 2 2
12 10 9 4 13 1 9 2 12 2 12 2 2
57 10 9 1 10 9 15 13 1 0 1 9 1 10 9 1 10 9 1 10 9 2 7 15 13 1 10 0 9 2 13 1 10 9 2 7 1 10 9 1 9 2 10 10 9 2 1 9 1 9 2 4 13 1 10 9 0 2
19 10 9 4 13 7 10 10 9 4 3 13 1 9 2 12 2 12 2 2
22 1 10 9 13 1 10 9 10 9 1 10 9 2 10 9 2 10 9 7 10 9 2
32 16 15 13 1 9 10 15 15 13 1 10 9 2 10 9 4 13 16 4 13 7 15 4 13 10 9 1 15 1 10 9 2
17 10 9 4 3 13 16 15 4 13 10 9 0 1 10 10 9 2
9 12 2 9 1 9 1 10 9 2
28 10 9 7 2 1 9 2 10 9 0 1 10 9 2 9 7 9 0 1 10 9 13 1 9 1 10 9 2
20 13 3 1 10 9 10 9 0 13 0 1 10 9 1 10 9 1 0 9 2
5 12 2 9 0 2
10 10 9 0 13 1 9 1 10 9 2
54 9 0 13 15 0 1 13 10 9 1 10 9 0 7 1 10 9 2 10 9 1 10 9 2 10 9 2 1 9 7 1 10 9 0 2 1 10 9 2 9 2 9 2 9 2 9 2 9 1 9 7 1 9 2
26 10 9 4 13 1 10 9 2 1 10 9 2 10 9 2 12 2 1 10 9 13 1 10 9 0 2
10 12 2 9 1 10 9 1 10 9 2
35 16 10 9 13 1 13 10 9 13 1 10 9 7 15 13 10 9 1 0 9 2 13 1 9 1 10 9 1 13 15 13 1 10 9 2
14 10 9 4 4 13 1 10 9 1 10 9 1 9 2
21 1 9 1 10 9 10 9 13 9 1 13 10 9 13 2 12 2 9 12 2 2
8 12 2 9 0 1 9 0 2
39 10 9 1 10 12 9 0 15 13 3 1 10 9 1 15 2 1 9 7 9 0 2 13 3 1 9 10 9 15 13 9 0 1 10 9 0 1 9 2
12 12 2 9 7 0 9 1 9 1 10 9 2
37 10 9 4 13 1 10 9 1 10 10 9 2 1 10 9 0 2 1 10 9 2 10 9 2 10 9 0 7 10 0 9 15 13 1 10 9 2
38 1 10 9 1 9 1 10 9 7 1 10 9 1 10 9 10 9 15 13 1 10 9 7 10 9 1 9 1 10 9 1 10 0 9 2 12 2 2
12 12 2 9 7 0 9 1 9 1 10 9 2
41 1 10 9 1 10 9 13 1 10 9 1 10 9 2 1 0 9 1 9 2 4 13 10 9 2 7 10 9 15 4 13 10 9 2 12 2 1 10 9 13 2
23 16 10 9 15 13 10 9 2 13 9 1 4 13 1 10 9 1 10 9 1 10 9 2
9 12 2 9 13 1 9 1 9 2
48 1 10 9 1 10 9 1 10 9 7 1 10 9 2 15 15 13 0 1 10 9 2 13 1 9 1 10 9 1 13 10 9 13 2 15 15 4 4 13 1 9 1 10 9 1 10 9 2
57 16 10 9 3 4 7 3 4 13 10 9 2 10 9 4 13 10 9 2 1 10 15 10 9 4 13 15 10 9 2 12 2 1 10 9 2 7 4 13 10 9 1 10 9 0 1 10 9 1 1 10 9 1 10 9 13 2
37 16 1 10 9 1 10 9 15 13 0 10 9 1 10 9 2 15 4 13 1 9 1 9 7 9 2 1 9 1 10 9 0 1 9 1 9 2
8 10 9 13 4 13 1 15 2
8 12 2 9 1 10 9 13 2
51 1 10 9 13 1 10 0 9 1 10 9 12 7 1 10 0 9 1 10 9 12 2 10 9 13 9 1 9 1 10 9 15 13 1 10 9 1 1 10 9 1 10 9 1 15 13 2 9 12 2 2
47 16 1 10 9 10 0 13 9 1 10 9 7 3 13 10 9 1 10 9 2 10 9 4 13 1 13 15 15 9 7 2 13 15 2 13 0 1 10 9 15 3 4 13 1 10 9 2
39 10 9 4 13 13 2 12 2 10 9 1 10 9 1 9 1 10 9 2 12 2 7 10 9 1 15 15 15 13 1 13 1 10 9 0 2 12 2 2
17 15 4 1 10 9 13 1 9 10 9 2 9 9 0 12 2 2
7 12 2 9 1 10 9 2
29 10 9 1 10 9 15 13 3 10 9 1 10 9 4 13 1 10 9 7 1 10 9 1 9 1 10 0 9 2
3 9 0 2
7 9 7 9 1 10 9 2
7 12 2 9 1 10 9 2
17 1 15 4 13 1 10 9 12 2 12 2 2 10 9 15 13 2
20 12 2 1 9 1 9 1 10 3 9 13 1 12 9 2 12 7 0 2 2
20 12 2 1 10 9 1 10 9 7 1 10 9 1 10 0 9 2 12 2 2
19 12 2 1 10 0 9 1 10 9 1 15 4 13 2 12 7 0 2 2
42 10 9 4 3 13 1 10 9 2 12 2 12 2 15 13 10 9 1 10 10 9 13 10 9 7 13 15 7 13 15 13 1 9 1 9 1 0 9 2 12 2 2
62 10 9 0 4 2 1 10 9 2 13 16 10 9 13 9 2 16 15 13 0 2 7 16 10 9 4 13 7 13 1 9 1 9 1 15 2 7 3 13 1 9 1 10 9 1 10 9 1 13 3 1 10 9 2 1 10 9 2 10 9 0 2
32 10 9 1 10 9 4 13 1 10 9 1 13 10 10 9 2 13 10 9 1 10 9 7 13 9 1 10 9 2 12 2 2
8 12 2 9 0 1 10 9 2
22 16 10 0 9 1 10 9 0 1 10 9 13 2 10 9 15 13 1 15 15 13 2
13 12 2 9 1 10 9 1 9 7 9 1 15 2
28 16 10 9 1 10 9 3 13 9 1 9 0 2 10 9 15 13 1 10 9 13 1 10 9 1 10 9 2
7 12 2 9 1 10 9 2
40 16 10 9 4 13 1 10 9 2 1 10 15 13 9 10 9 2 7 15 13 1 10 9 1 13 2 10 9 13 9 1 13 1 10 9 7 1 10 9 2
60 1 10 9 2 3 2 10 9 2 16 13 13 10 0 9 2 13 10 9 1 13 10 9 7 1 13 15 1 10 9 2 13 1 10 9 2 1 10 9 2 10 9 2 12 2 1 10 9 0 1 10 9 1 10 9 7 1 10 9 2
36 16 10 9 4 13 1 10 9 1 10 9 7 1 10 9 1 10 9 1 10 9 3 13 2 10 9 15 13 1 10 9 13 1 10 9 2
12 10 9 1 10 9 15 13 1 10 9 13 2
33 16 3 10 9 13 1 10 9 13 0 1 15 13 1 9 2 10 9 1 10 9 1 10 0 9 4 13 1 9 1 10 15 2
6 12 2 9 7 9 2
3 9 0 2
8 1 10 9 7 1 10 9 2
48 15 13 10 9 1 9 1 10 9 2 4 13 15 1 15 7 2 16 13 0 2 4 13 10 9 2 12 2 1 15 13 1 10 9 10 7 1 10 10 9 2 12 7 0 2 12 2 2
16 10 9 15 4 13 1 10 9 0 1 10 9 1 10 9 2
23 15 13 10 9 1 9 1 10 9 4 13 15 3 1 10 9 10 7 1 10 10 9 2
7 12 2 9 1 10 9 2
38 1 10 9 15 13 3 10 9 13 3 16 4 13 10 9 1 9 7 1 9 2 16 1 10 9 1 15 10 9 4 13 10 9 3 4 13 9 2
30 15 13 3 10 9 15 13 1 10 9 1 10 9 1 13 1 15 7 1 10 10 9 10 10 9 2 9 12 2 2
6 12 2 9 1 9 2
19 10 9 1 9 7 1 9 3 15 4 13 2 12 2 7 13 1 9 2
12 12 2 9 0 1 10 9 7 1 10 9 2
53 15 13 10 9 1 10 9 7 15 13 10 10 9 7 15 13 10 9 1 9 7 13 10 10 9 4 13 1 10 9 1 9 2 1 10 9 0 7 1 10 9 1 10 9 1 10 9 2 12 7 0 2 2
27 16 3 13 16 10 9 1 10 9 7 3 13 16 10 9 1 10 9 2 13 1 9 1 15 15 13 2
10 12 2 9 1 10 9 1 10 9 2
26 10 9 0 1 10 9 2 12 7 0 2 15 13 2 1 3 0 2 1 10 9 7 1 10 9 2
3 9 0 2
3 9 0 2
3 9 0 2
7 12 2 9 1 10 9 2
16 10 9 4 13 3 1 10 0 9 7 9 1 10 9 13 2
19 4 1 10 9 13 0 1 10 9 0 1 10 9 2 12 7 0 2 2
7 12 2 9 1 9 0 2
16 4 13 10 9 1 10 9 1 13 1 10 9 10 9 0 2
49 4 13 3 1 9 7 1 9 1 10 9 1 13 7 1 10 9 1 13 2 7 1 10 9 10 9 3 13 9 16 3 1 10 9 1 15 10 9 4 13 7 10 9 4 13 2 12 2 2
5 12 2 9 0 2
46 10 9 1 10 9 13 3 4 13 1 13 10 9 1 13 0 10 9 1 10 9 1 9 1 10 9 2 3 16 10 9 7 10 9 13 3 2 12 7 0 2 12 7 0 2 2
7 12 2 9 1 10 9 2
22 10 9 0 4 4 13 3 2 12 2 12 7 0 2 7 3 2 12 7 0 2 2
20 4 3 4 13 1 9 7 1 9 1 10 9 1 9 2 12 7 0 2 2
5 1 10 9 0 2
6 12 2 9 1 9 2
52 16 2 1 9 1 9 2 10 9 1 10 9 13 9 1 13 1 9 1 10 9 1 10 0 9 10 9 1 10 9 2 15 2 1 9 1 9 2 4 13 1 9 2 12 2 12 9 12 2 12 2 2
24 4 3 4 13 1 9 1 10 9 0 1 10 9 3 13 1 10 9 2 12 7 0 2 2
14 10 9 13 10 9 1 10 9 7 13 10 9 13 2
23 3 1 10 9 1 10 9 10 9 1 10 9 13 4 13 15 1 10 9 1 10 9 2
9 1 10 9 7 1 10 9 0 2
10 12 2 9 1 13 9 1 10 9 2
49 10 9 4 13 1 13 9 1 10 10 9 1 10 9 1 10 9 15 15 4 13 1 9 1 15 13 2 3 3 3 2 10 9 1 13 15 1 10 9 1 10 9 7 1 9 0 7 0 2
20 13 0 1 10 9 10 9 2 10 9 2 10 9 7 10 9 1 15 0 2
7 12 2 9 1 0 9 2
37 15 13 9 1 13 9 1 10 9 10 4 13 10 0 9 2 7 3 4 13 13 10 9 1 10 9 3 13 7 13 1 10 9 1 0 9 2
38 10 9 1 10 9 0 1 10 9 4 3 13 10 9 2 13 10 9 1 10 10 9 3 13 2 16 15 3 13 0 9 1 10 9 15 15 13 2
51 1 10 9 1 10 9 1 10 9 4 13 10 9 1 13 15 13 9 1 10 9 15 15 13 2 1 10 9 1 10 9 2 1 10 9 15 15 13 0 1 10 0 9 7 1 10 0 9 1 9 2
25 10 9 13 1 10 9 0 3 4 13 1 10 9 1 10 9 13 1 10 9 1 10 0 9 2
6 12 2 9 1 9 2
55 15 4 13 10 9 1 10 9 10 4 13 1 10 1 3 7 1 10 1 3 10 9 0 2 13 15 1 10 9 1 10 9 7 1 15 2 16 13 10 9 0 1 13 10 9 7 9 1 10 9 0 2 12 2 2
9 12 2 9 1 9 7 1 9 2
32 16 1 10 9 1 10 9 13 13 9 0 7 0 1 9 0 2 15 13 10 9 7 10 9 1 10 9 7 1 10 9 2
27 15 4 13 13 10 9 1 10 9 10 4 13 16 4 13 1 10 9 1 10 9 1 15 13 10 9 2
15 16 10 15 13 0 1 10 9 1 10 15 15 4 13 2
49 16 10 9 13 13 10 3 0 7 10 3 0 1 10 9 13 2 13 9 1 10 9 1 10 9 0 2 1 10 9 7 1 10 0 9 1 10 9 2 1 10 9 7 10 9 1 10 9 2
76 3 1 13 10 9 1 10 9 2 15 4 13 9 1 10 9 10 4 13 10 9 2 1 10 9 2 1 10 9 1 13 2 1 9 1 10 9 7 1 10 0 9 0 1 10 9 2 1 10 9 1 10 9 2 3 13 15 13 1 10 9 1 12 7 10 9 7 1 0 9 1 10 9 1 13 2
52 1 10 9 2 3 2 15 4 13 3 1 10 9 1 10 9 13 7 1 10 9 1 10 9 3 15 4 13 16 10 9 1 10 9 1 10 9 2 7 3 1 9 1 10 9 7 1 10 0 9 0 2
56 16 10 9 1 10 9 4 13 1 10 9 3 0 1 12 9 2 10 9 1 10 9 7 1 10 9 13 1 10 9 0 4 13 1 10 0 9 2 7 1 10 9 2 13 10 9 2 1 13 10 9 1 10 0 9 2
39 10 9 0 4 4 13 0 3 1 10 9 1 10 9 1 10 9 1 10 0 9 1 10 9 0 2 12 2 1 10 9 1 15 10 9 4 4 13 2
20 13 10 9 2 3 15 13 3 9 1 15 15 4 4 13 1 10 9 0 2
7 12 2 9 1 10 9 2
34 15 13 10 9 1 10 9 10 3 4 13 15 0 9 1 9 2 16 10 9 3 15 13 0 7 15 4 13 9 1 10 9 13 2
55 16 10 9 1 10 0 9 1 9 13 0 9 2 15 3 4 13 15 2 16 3 3 15 15 13 10 9 7 10 9 7 3 15 13 10 9 13 1 10 9 1 13 7 1 10 9 1 10 9 13 1 10 9 12 2
24 10 0 9 15 13 3 16 1 10 9 1 10 9 13 13 10 9 1 10 9 9 7 3 2
7 12 2 9 1 10 9 2
34 13 3 1 9 1 10 9 1 10 9 13 1 13 13 3 10 9 1 10 9 1 10 9 1 9 7 9 1 13 15 1 9 0 2
29 16 3 1 10 9 15 3 4 13 9 1 10 9 1 10 9 1 10 9 2 4 13 10 9 1 10 9 13 2
14 12 2 9 0 1 10 9 1 9 0 1 9 10 2
105 16 10 9 1 9 13 1 10 9 1 10 9 0 10 9 1 10 15 2 7 10 9 1 10 9 7 1 10 9 1 10 9 2 15 15 15 13 1 10 9 4 13 2 1 9 1 10 9 15 15 13 2 1 13 7 1 13 10 9 7 10 10 9 0 1 10 0 7 0 9 2 1 3 10 9 0 2 10 9 2 9 7 0 9 0 1 13 10 9 7 10 9 2 0 10 9 13 1 10 9 7 1 10 9 2
5 12 2 9 0 2
40 10 9 13 1 10 9 0 1 10 9 1 10 9 15 13 3 16 10 9 4 13 1 10 9 1 13 9 13 15 10 9 3 13 1 13 1 10 10 9 2
23 10 9 4 4 3 13 1 9 0 2 16 4 13 10 9 0 1 13 10 9 7 9 2
79 0 10 9 1 10 9 1 10 9 7 1 10 9 0 2 10 9 15 13 13 7 13 10 10 9 1 9 2 1 9 7 0 9 13 9 2 13 10 9 1 10 9 7 1 10 0 9 0 2 1 13 1 9 7 1 9 10 9 1 9 1 10 9 15 13 10 10 9 1 10 9 1 9 7 1 10 0 9 2
67 16 10 9 13 1 9 1 10 9 1 15 15 13 10 9 13 1 10 9 0 2 7 16 10 0 9 3 15 4 13 1 0 9 15 13 10 9 0 1 10 9 2 10 9 0 13 10 9 1 13 10 9 0 2 13 1 10 9 9 1 10 9 0 1 10 9 2
24 16 15 13 9 1 10 9 2 4 4 13 10 0 9 1 15 15 1 10 9 15 4 13 2
10 12 2 9 1 9 7 1 9 10 2
108 10 9 1 10 9 13 1 9 7 1 9 10 2 7 15 3 4 13 1 10 9 13 1 9 1 10 9 0 2 13 9 1 13 15 15 1 13 10 10 9 2 1 9 16 3 15 13 9 1 10 9 3 13 7 16 15 13 10 0 9 13 1 13 10 9 3 13 2 16 15 13 1 9 1 13 3 1 10 9 13 2 7 3 13 10 9 0 1 10 9 3 13 7 1 15 13 1 10 9 1 10 9 2 10 15 13 0 2
10 12 2 9 1 10 9 1 10 9 2
31 1 10 9 1 10 9 13 1 10 9 0 13 0 10 9 1 10 0 9 1 10 9 12 7 1 10 9 12 7 12 2
3 9 0 2
7 12 2 9 1 10 9 2
7 12 2 9 1 10 9 2
49 1 10 9 7 1 10 9 1 10 9 1 9 1 10 0 9 2 4 13 15 1 10 9 0 7 10 0 10 0 9 15 4 13 1 10 9 2 1 10 9 7 1 10 9 1 10 9 0 2
3 9 0 2
14 1 10 9 0 1 9 1 10 9 7 1 10 9 2
9 12 2 9 1 9 1 10 9 2
67 16 1 10 9 7 1 10 10 9 13 10 9 0 1 10 9 1 10 9 7 1 10 9 7 1 10 0 9 0 2 7 3 13 0 13 15 1 0 9 2 10 9 1 10 9 0 4 2 12 2 13 16 4 13 10 9 1 9 1 10 9 0 1 10 9 0 2
27 3 16 4 13 10 9 2 4 13 15 10 9 1 10 9 2 15 15 13 1 13 2 13 1 10 9 2
16 15 4 3 13 10 10 9 1 10 9 1 9 7 1 9 2
14 15 13 3 10 9 1 10 0 9 1 10 9 12 2
23 1 9 1 9 2 10 9 13 10 9 1 10 9 7 10 9 13 2 12 2 12 2 2
9 12 2 9 1 9 1 10 9 2
45 10 9 13 1 10 9 0 15 13 3 16 10 9 1 10 9 3 13 9 1 13 15 2 16 10 9 1 10 9 0 13 10 0 9 2 1 13 10 9 0 2 0 7 0 2
28 10 9 1 10 9 7 1 10 9 3 15 13 1 10 9 1 15 1 10 9 15 13 1 9 1 9 0 2
3 9 0 2
5 1 10 9 0 2
5 12 2 9 0 2
57 10 9 2 10 10 9 4 13 1 9 10 2 7 15 3 13 9 1 10 9 0 7 4 13 15 15 1 0 9 7 9 2 13 9 2 12 2 1 13 10 9 1 10 9 0 1 10 9 7 10 0 9 1 10 10 9 2
36 10 9 15 4 13 2 12 2 1 10 9 1 15 10 9 1 10 9 0 13 3 0 7 13 1 0 9 1 10 9 1 10 15 4 13 2
31 15 4 4 13 3 1 9 2 16 15 13 0 2 13 9 1 10 9 1 10 9 13 7 1 10 9 1 10 9 13 2
40 10 0 9 15 13 1 10 9 1 15 15 2 13 10 9 1 10 9 10 2 13 9 1 10 9 0 1 13 15 1 10 9 1 10 9 3 1 9 0 2
11 12 2 9 0 1 9 1 9 3 0 2
42 10 9 1 10 9 0 15 4 13 3 16 10 9 1 10 9 13 10 9 1 10 9 0 2 7 15 13 0 7 0 1 10 9 1 10 9 7 3 4 4 13 2
31 10 9 4 4 13 1 10 9 0 2 12 2 3 16 15 13 16 10 9 13 1 10 9 1 10 9 7 1 10 9 2
22 1 10 9 13 1 10 12 9 0 4 13 10 9 0 1 10 9 13 1 10 9 2
61 16 2 1 13 10 9 2 13 0 13 1 9 0 7 13 0 10 9 1 10 9 13 2 10 9 15 15 13 4 2 3 1 13 10 9 7 1 13 10 9 2 13 10 9 1 10 9 13 1 10 9 13 1 10 0 9 1 10 9 12 2
11 12 2 9 1 9 1 9 7 1 9 2
37 16 10 9 4 13 1 10 9 0 1 9 1 9 1 9 0 2 10 9 13 9 1 13 1 10 0 9 10 9 1 10 9 2 9 12 2 2
13 10 0 9 15 13 1 9 1 9 2 12 2 2
7 12 2 9 1 10 9 2
29 16 10 9 13 1 13 0 2 4 4 13 1 10 9 1 9 1 10 9 1 10 9 13 7 1 10 9 13 2
8 10 0 4 13 10 9 13 2
3 9 0 2
13 1 10 9 0 7 1 10 9 0 1 9 0 2
7 12 2 9 1 9 0 2
27 10 9 4 13 2 12 2 1 13 9 1 10 10 9 1 10 9 0 2 1 9 1 10 9 1 9 2
7 12 2 9 1 9 0 2
50 10 9 4 3 13 1 13 13 1 10 10 9 10 9 1 9 0 0 1 9 0 7 0 7 1 13 1 10 9 10 9 2 10 9 7 10 9 0 1 10 9 2 1 9 1 10 9 1 9 2
3 9 0 2
5 1 10 9 0 2
6 12 2 9 1 9 2
32 10 9 0 4 4 13 1 9 2 12 2 12 2 12 9 12 2 12 9 12 2 7 1 9 2 12 7 0 2 12 2 2
10 12 2 9 13 1 15 1 10 9 2
32 10 9 13 1 15 1 10 9 1 10 9 0 3 4 13 16 3 16 10 15 15 4 3 15 13 3 7 3 2 12 2 2
40 10 9 2 3 2 13 1 15 1 10 9 2 3 1 10 15 2 13 10 13 2 7 10 10 9 7 13 9 1 3 13 9 1 10 9 1 10 9 13 2
9 12 2 9 13 1 10 0 9 2
30 10 9 4 2 1 10 9 1 10 9 2 13 1 10 9 10 9 15 3 13 10 9 1 9 2 12 2 12 2 2
3 9 0 2
15 1 10 9 13 1 9 7 1 9 1 10 9 1 9 2
6 12 2 9 3 0 2
28 10 9 3 0 3 4 13 15 1 9 2 12 2 9 12 2 7 1 9 1 10 9 1 9 2 12 2 2
19 3 0 13 10 9 16 3 15 13 9 0 7 0 13 1 10 10 9 2
9 12 2 9 1 10 9 1 9 2
57 10 9 1 10 9 1 9 13 9 16 13 2 1 10 9 1 9 2 12 7 0 2 2 16 12 9 2 3 13 2 4 4 13 1 10 0 9 2 7 16 15 4 13 7 13 10 9 1 10 9 1 10 15 13 10 9 2
37 16 10 12 9 13 1 13 1 10 0 9 2 1 10 9 0 1 10 9 2 15 15 13 13 3 7 3 1 9 7 1 15 1 10 9 0 2
3 9 0 2
7 1 10 9 1 10 9 2
23 10 9 7 10 9 1 10 9 4 13 1 10 9 7 2 1 9 2 1 10 9 0 2
9 12 2 9 1 10 9 1 9 2
14 10 9 1 9 13 10 15 15 13 0 1 13 15 2
36 16 10 9 4 13 2 12 2 2 10 9 4 13 15 0 7 0 10 9 1 15 13 10 9 1 9 15 13 0 10 9 1 10 9 0 2
12 12 2 9 0 1 10 9 7 1 10 9 2
25 15 15 13 10 9 1 9 3 4 13 15 16 3 1 9 1 10 10 9 7 1 10 10 9 2
7 12 2 9 1 10 9 2
44 1 10 9 1 9 1 10 9 15 13 9 1 10 9 1 10 9 0 7 2 16 15 13 1 9 13 1 9 0 1 10 9 2 15 13 9 1 10 9 1 10 0 9 2
13 12 2 9 1 13 7 13 10 9 1 10 9 2
21 10 9 1 10 9 13 3 4 13 9 15 13 3 0 10 9 1 10 9 13 2
27 10 9 1 10 9 13 3 4 13 10 9 15 13 1 13 10 9 1 10 9 7 1 13 15 3 0 2
10 12 2 9 1 10 9 1 9 0 2
27 10 9 1 10 9 13 3 4 13 10 9 1 10 9 1 9 0 1 15 1 10 15 4 4 13 3 2
64 3 2 16 10 0 9 4 13 3 0 1 10 9 13 7 16 13 1 13 9 2 9 7 9 2 10 9 1 10 9 13 4 13 1 10 9 1 10 0 9 10 9 3 0 1 10 9 1 10 10 9 2 7 15 3 4 13 15 2 12 2 12 2 2
53 10 9 1 9 1 10 9 1 10 9 15 4 1 10 9 13 1 9 2 9 9 0 12 2 1 10 9 1 10 9 13 2 16 15 13 16 10 9 13 1 15 1 0 9 7 3 13 9 1 10 9 13 2
45 10 9 0 4 3 13 16 10 9 4 13 1 0 9 1 10 9 1 10 9 13 7 1 10 15 15 15 13 2 16 10 9 1 15 13 3 0 1 10 9 1 10 9 13 2
8 12 2 9 1 10 9 13 2
39 10 9 1 10 9 13 2 1 10 13 10 9 0 1 13 10 9 2 4 13 10 9 7 10 9 15 13 1 13 0 9 1 10 9 1 10 9 13 2
25 15 4 13 10 9 1 10 9 2 3 16 4 3 13 1 10 9 7 1 10 9 2 12 2 2
22 16 3 10 9 13 3 1 10 9 13 2 10 9 4 13 1 9 1 10 0 9 2
8 12 2 9 1 10 9 13 2
66 10 9 1 10 9 13 2 16 4 13 1 9 1 10 9 7 1 10 9 1 10 9 0 1 10 9 7 1 10 9 1 10 9 2 12 2 2 4 3 13 15 15 2 13 1 10 9 1 10 9 13 1 9 1 10 9 1 10 9 13 2 12 2 12 2 2
29 1 10 9 1 15 10 9 1 10 9 4 13 1 10 9 1 10 9 2 10 9 4 13 15 1 10 9 0 2
13 12 2 9 1 10 9 13 7 1 10 9 13 2
29 16 10 9 13 4 13 2 10 9 4 13 1 10 9 2 1 16 3 15 13 3 0 10 9 1 10 9 13 2
25 16 10 9 13 4 13 7 10 9 13 1 10 9 0 1 10 9 0 2 10 0 9 4 13 2
3 9 0 2
7 1 10 9 1 10 9 2
6 12 2 9 1 9 2
6 12 2 9 1 9 2
20 10 9 15 13 1 9 16 3 15 15 13 1 12 9 2 12 7 0 2 2
44 7 2 16 15 13 1 9 0 7 1 9 1 10 10 9 3 13 0 10 9 1 10 9 2 10 9 13 1 10 9 1 15 15 4 13 10 9 15 15 4 13 10 9 2
31 1 10 9 15 15 13 1 9 2 10 9 13 1 10 9 1 15 10 9 15 4 4 13 7 3 15 4 13 10 9 2
24 1 10 9 1 10 9 15 13 3 10 9 1 10 15 10 9 3 4 13 1 10 0 9 2
28 16 10 9 13 13 1 10 9 1 9 2 10 9 1 10 9 13 1 15 1 15 13 10 9 3 1 15 2
26 10 9 7 10 9 1 10 9 2 12 7 0 2 1 9 1 15 1 10 9 13 3 1 10 15 2
10 12 2 9 1 9 7 9 1 9 2
37 10 9 1 9 1 13 1 10 9 7 10 13 3 1 10 9 1 10 15 3 13 13 10 9 2 16 3 4 13 10 9 13 1 10 9 0 2
26 10 9 13 1 9 1 13 15 10 9 0 1 15 13 1 10 9 15 13 1 9 2 9 12 2 2
14 9 1 10 9 3 0 1 10 9 7 1 10 9 2
26 10 9 1 10 9 1 9 0 1 15 13 1 10 9 7 1 10 9 3 15 13 10 9 1 9 2
7 9 13 1 10 9 0 2
14 9 13 1 9 1 10 9 0 2 0 7 1 9 2
22 10 9 13 1 10 9 1 9 1 10 9 0 3 13 1 10 13 15 1 10 9 2
9 1 10 9 1 9 1 10 9 2
10 9 1 10 9 7 0 9 1 9 2
37 10 9 1 10 9 4 13 15 13 1 9 10 9 1 15 15 13 10 9 2 12 2 7 4 13 13 10 0 9 7 9 2 12 7 0 2 2
21 4 3 13 10 9 1 10 9 1 9 2 1 10 9 1 10 9 2 12 2 2
8 1 10 9 1 9 1 9 2
15 10 9 1 10 9 1 9 0 15 4 13 1 10 9 2
26 1 10 9 1 15 4 13 7 13 10 0 9 1 9 2 10 9 4 13 15 1 9 1 10 9 2
29 15 13 10 9 1 9 15 13 1 10 0 9 1 12 9 1 10 9 0 7 15 13 1 9 2 9 7 9 2
10 9 1 10 9 7 1 10 9 0 2
38 16 2 1 10 9 1 10 0 7 0 9 1 9 0 2 4 4 13 10 9 1 10 9 7 1 10 9 0 2 10 9 3 4 13 15 10 9 2
37 16 10 9 3 4 4 13 2 7 10 9 7 10 9 0 4 4 13 7 13 1 12 9 2 3 4 3 13 1 10 9 10 9 1 10 9 2
17 1 9 1 9 7 1 9 2 10 9 4 13 1 10 9 0 2
32 16 10 9 1 9 3 4 4 13 2 7 10 9 4 4 13 1 10 0 9 2 15 13 13 10 9 0 1 10 9 0 2
35 1 10 9 1 10 9 1 9 1 9 2 16 3 13 10 9 7 3 13 0 13 15 1 10 9 2 12 2 2 15 13 10 9 0 2
15 1 9 1 10 9 15 13 10 9 1 10 12 9 0 2
25 10 9 1 10 9 1 9 15 13 2 1 10 9 0 2 1 10 9 1 9 1 15 1 9 2
20 10 9 1 9 1 9 7 1 9 15 13 1 10 9 7 1 10 9 0 2
35 10 9 1 10 9 1 10 9 0 4 13 1 10 9 1 9 13 1 10 9 1 15 10 9 4 13 7 1 15 15 4 13 1 13 2
42 1 10 9 1 9 10 9 15 13 10 9 1 13 1 10 9 1 9 1 10 9 15 13 1 10 9 2 7 10 9 1 10 9 13 1 15 1 15 13 10 9 2
42 1 10 9 0 1 9 1 9 10 9 13 7 13 2 7 13 1 10 9 1 10 9 2 3 4 13 15 7 13 15 1 10 9 16 1 10 9 1 10 10 9 2
25 10 9 1 10 0 9 4 13 7 13 1 15 10 9 2 16 10 9 3 13 9 1 10 15 2
30 15 13 9 1 13 15 1 10 9 1 9 0 3 4 2 1 0 9 1 10 9 2 13 15 7 13 15 10 9 2
14 9 1 10 13 1 1 10 9 1 9 1 10 9 2
29 10 9 1 10 9 4 4 13 1 15 13 9 1 13 15 7 1 13 15 1 10 9 1 15 10 9 15 13 2
30 10 13 1 10 9 4 13 1 10 0 9 1 10 9 1 10 9 1 10 9 13 15 1 9 0 7 1 9 10 2
16 1 10 9 4 13 10 0 9 1 10 9 1 10 9 13 2
9 9 1 10 9 0 1 10 9 2
27 15 13 9 0 10 9 1 10 9 1 9 13 7 13 1 10 9 1 10 9 1 15 10 9 4 13 2
9 9 1 10 9 1 10 9 13 2
46 10 9 1 10 9 3 13 1 10 9 1 10 9 13 10 9 1 13 3 1 10 9 1 9 1 10 10 9 2 1 13 10 9 1 15 7 1 13 1 15 7 1 9 10 9 2
43 16 10 9 4 13 2 13 7 13 2 12 2 1 10 0 9 2 1 9 1 10 13 7 1 15 1 15 15 15 13 2 10 9 3 4 13 15 1 9 1 10 9 2
42 10 9 1 10 9 0 1 10 9 1 10 9 7 1 10 9 1 9 4 3 13 15 1 10 9 1 10 9 7 10 9 1 10 9 13 1 10 9 1 9 0 2
12 10 9 1 10 9 1 10 9 15 13 0 2
26 10 9 1 10 9 2 3 1 10 9 3 1 10 9 1 10 9 2 13 1 9 1 10 0 9 2
33 10 9 4 13 15 1 10 9 0 2 16 3 15 13 10 9 7 3 13 1 10 0 9 1 13 15 3 9 1 10 10 9 2
19 1 10 9 4 13 1 10 9 10 9 0 1 10 0 9 1 10 9 2
36 10 9 3 4 13 10 10 9 1 10 9 0 1 9 1 10 0 9 2 16 3 13 0 0 1 13 10 9 1 10 10 9 2 12 2 2
25 10 9 4 13 1 10 10 9 7 13 1 15 10 9 1 10 9 1 10 9 1 10 10 9 2
30 1 10 9 13 1 15 1 10 9 15 13 10 9 0 1 10 9 0 1 10 9 0 1 10 9 0 2 12 2 2
34 10 9 4 13 1 10 9 0 1 10 9 7 1 10 9 1 10 9 0 7 1 10 9 13 1 10 9 1 9 1 10 9 0 2
15 10 9 3 13 1 10 9 15 4 3 3 13 10 9 2
31 10 9 2 12 2 1 10 9 4 13 1 9 2 12 7 0 2 1 10 13 1 13 10 9 1 15 13 7 3 13 2
18 10 10 9 13 9 1 13 1 10 9 1 10 9 0 2 12 2 2
31 1 10 9 1 0 9 10 9 1 10 9 1 10 9 2 13 1 10 9 1 10 10 9 2 13 0 1 10 9 0 2
26 1 10 9 1 10 9 1 10 9 15 13 16 10 10 9 4 4 3 13 1 10 9 1 10 9 2
39 16 3 15 13 10 9 0 1 10 9 1 10 9 0 7 3 15 13 10 9 2 7 16 10 9 13 3 4 13 2 10 9 4 13 1 10 9 0 2
16 15 13 1 9 1 9 7 4 3 13 10 9 2 12 2 2
9 9 1 10 9 7 9 1 9 2
32 1 10 9 13 1 10 9 13 1 10 9 0 2 4 4 13 10 9 1 10 0 9 7 1 10 0 9 1 10 9 0 2
32 1 10 0 9 10 9 4 4 13 1 15 7 10 9 2 7 3 1 10 9 2 13 15 10 9 7 10 9 1 10 9 2
31 15 1 10 9 0 4 13 3 1 10 9 0 10 9 1 10 9 1 12 9 2 12 2 1 10 9 15 15 4 13 2
15 10 9 0 13 1 0 9 1 10 9 13 2 12 2 2
32 13 10 9 13 1 10 9 0 1 16 10 9 4 4 13 2 15 13 9 3 1 10 9 7 10 13 9 1 10 0 9 2
9 9 7 0 9 13 10 0 9 2
46 1 9 1 10 9 1 10 9 15 13 3 12 9 1 10 9 0 1 10 9 0 2 15 4 13 10 10 9 0 1 10 9 1 10 9 7 1 13 15 3 0 7 0 10 9 2
29 1 10 0 9 15 4 13 10 0 9 13 10 0 9 2 3 16 3 13 0 1 10 9 1 15 1 10 9 2
34 13 0 10 9 1 10 10 9 1 10 9 1 9 7 1 9 1 9 0 1 10 9 0 7 1 10 9 1 9 0 1 12 9 2
39 10 9 4 4 3 13 1 10 9 13 1 10 0 9 2 16 13 10 9 1 13 10 9 1 10 9 13 1 10 9 7 1 10 9 1 10 9 0 2
20 15 1 10 9 10 9 0 4 13 3 1 10 9 0 10 9 1 10 9 2
23 10 9 4 4 13 2 1 9 1 9 2 12 7 0 2 2 1 12 9 1 10 9 2
5 9 1 10 9 2
18 1 9 1 10 9 2 10 9 0 4 13 10 9 1 10 9 13 2
16 15 1 10 9 4 3 13 10 9 1 10 9 2 12 2 2
33 10 9 0 4 13 10 0 9 2 1 10 9 3 0 1 12 9 2 16 10 0 9 4 13 10 9 1 10 15 2 12 2 2
28 10 9 1 13 1 9 1 10 9 3 0 1 12 9 13 0 7 13 9 3 1 10 13 9 1 10 9 2
16 16 4 4 13 1 10 9 0 1 15 15 13 1 12 9 2
22 16 0 9 15 13 2 10 9 0 4 13 10 9 1 10 9 3 1 10 9 13 2
30 10 9 1 10 9 3 4 4 13 16 15 13 1 9 15 2 16 13 2 13 1 13 1 10 9 1 15 4 13 2
35 10 9 7 10 13 9 1 10 9 4 13 1 10 9 1 10 9 2 7 3 4 13 10 9 3 13 2 1 3 16 4 13 10 9 2
29 10 9 13 9 1 9 2 16 10 9 4 4 3 13 1 9 13 1 10 9 1 10 9 2 12 7 0 2 2
35 10 9 4 13 16 4 13 10 9 1 9 2 12 2 13 1 10 9 0 2 10 15 4 13 7 13 1 10 9 1 10 9 1 9 2
32 10 9 15 4 13 10 9 1 9 7 3 4 13 9 13 1 10 9 1 10 0 9 13 1 10 10 9 1 10 0 13 2
38 1 10 9 1 10 9 0 15 13 10 9 1 10 9 1 10 9 2 12 7 0 2 12 7 0 2 2 1 3 3 13 1 9 1 15 3 13 2
29 13 9 1 9 0 1 10 9 1 10 10 9 7 9 1 9 1 10 9 2 16 10 9 3 13 1 10 9 2
9 9 1 10 9 1 10 9 0 2
36 10 9 1 10 9 1 10 9 13 1 10 9 0 13 0 1 10 9 1 10 9 7 9 1 9 15 15 13 2 16 10 9 3 13 3 2
30 10 9 3 4 2 13 1 10 9 1 10 9 0 2 13 15 1 10 9 1 10 9 1 10 10 9 2 12 2 2
33 10 9 0 1 10 9 3 13 0 1 9 2 1 3 16 10 9 4 13 15 1 13 3 0 10 9 1 10 9 1 10 9 2
44 10 9 2 1 10 9 13 1 10 0 9 1 10 9 12 2 4 13 10 10 9 0 1 10 9 7 1 10 9 3 0 7 1 10 0 9 1 10 9 0 2 12 2 2
43 4 13 10 9 15 4 13 9 1 10 9 7 1 10 9 1 10 9 2 15 15 13 10 9 0 7 15 13 10 9 0 1 10 9 0 1 10 9 7 1 10 9 2
34 16 10 9 0 3 13 0 2 10 9 3 4 13 2 3 16 10 9 1 10 9 15 15 4 13 7 13 13 13 15 3 10 9 2
45 1 10 9 13 1 10 0 9 10 9 7 10 10 9 7 13 9 4 3 2 1 10 9 2 13 1 10 9 1 10 9 2 13 1 10 9 1 9 7 1 9 1 10 9 2
11 9 1 10 9 1 10 9 1 9 0 2
29 10 9 2 1 10 9 7 9 1 9 1 10 9 2 3 4 13 9 15 13 9 1 10 9 0 1 10 9 2
17 10 9 4 13 7 13 1 10 9 1 10 10 9 1 15 13 2
43 1 10 9 1 10 9 1 10 9 1 10 9 2 15 4 13 1 9 1 10 9 2 15 13 1 9 10 9 2 10 9 0 2 10 9 7 9 1 9 7 10 9 2
28 10 9 0 2 13 0 9 1 10 9 2 4 13 10 9 1 10 9 2 7 13 15 2 13 10 0 9 2
17 10 9 0 2 16 15 13 10 9 13 0 9 1 10 9 0 2
29 10 9 13 1 9 2 1 9 0 2 7 1 10 0 9 2 7 9 0 1 13 15 1 9 1 10 9 0 2
26 10 9 7 10 9 4 13 15 1 10 9 1 10 9 2 1 9 1 10 9 1 10 9 0 2 2
30 1 10 9 1 10 9 0 1 10 9 1 10 9 0 2 10 9 4 13 15 1 9 1 10 9 1 10 9 13 2
17 10 9 1 13 10 9 0 13 15 1 13 15 3 1 10 9 2
29 16 10 9 13 1 9 10 9 1 9 13 3 1 10 9 2 10 9 4 13 9 1 9 3 0 1 10 9 2
36 15 4 13 1 13 10 9 2 1 16 15 4 13 10 9 7 10 9 2 4 13 1 10 9 10 0 9 0 7 0 2 7 10 0 9 2
31 10 9 4 4 13 1 10 15 2 3 1 10 9 1 10 9 2 16 15 3 13 9 1 16 10 9 13 3 10 9 2
23 3 10 9 4 13 10 9 13 15 1 10 15 2 16 10 9 15 4 13 10 10 9 2
24 10 9 4 13 10 9 0 3 16 10 9 13 0 2 3 16 10 9 7 10 9 13 3 2
44 16 10 9 1 10 15 10 9 4 4 13 3 4 13 1 10 9 7 1 10 9 7 3 4 13 15 1 10 9 1 10 9 7 1 0 9 2 15 13 10 9 15 13 2
27 10 9 1 13 10 9 0 7 0 4 4 13 1 10 9 1 15 15 13 10 9 16 10 9 4 13 2
26 10 9 13 1 9 10 9 1 9 4 4 13 1 10 9 15 10 9 13 1 10 9 1 10 9 2
44 16 10 9 13 15 1 15 15 10 9 13 16 4 13 10 9 7 15 13 3 0 10 9 2 10 9 2 0 9 1 10 9 2 13 9 1 13 10 9 1 10 10 9 2
23 1 10 0 9 10 9 4 4 13 1 10 9 15 10 9 13 1 10 9 1 10 9 2
21 16 3 4 13 10 9 1 15 10 9 4 4 13 2 10 9 4 13 15 3 2
47 16 3 2 1 9 1 10 9 7 1 10 9 1 10 9 7 1 10 9 7 10 9 1 10 9 2 13 0 10 9 2 15 2 1 9 1 9 1 10 9 2 4 13 1 10 9 2
27 16 10 9 1 10 9 4 13 1 10 9 1 10 9 2 13 3 1 10 9 1 13 15 1 10 9 2
25 16 4 13 1 10 9 1 10 9 2 10 9 4 4 13 1 9 1 10 9 15 13 13 15 2
31 16 1 10 9 4 13 10 9 2 15 15 13 1 9 1 10 9 2 16 3 13 13 1 9 1 10 9 7 1 15 2
23 10 9 3 4 13 10 9 1 1 10 9 2 3 16 10 9 4 13 3 1 10 9 2
19 10 9 13 1 10 9 1 10 9 4 13 1 10 9 1 10 9 12 2
23 10 9 0 1 10 9 1 10 9 15 13 1 9 0 15 13 16 3 15 13 9 0 2
9 13 0 1 10 9 10 0 9 2
34 10 9 4 4 13 1 10 9 7 1 10 10 9 7 1 10 9 13 1 10 9 7 13 1 10 9 7 1 10 9 1 13 15 2
26 10 9 13 1 15 3 4 13 1 13 15 13 10 9 2 16 10 9 15 13 7 16 15 4 13 2
30 10 9 15 13 10 9 1 15 13 13 1 13 15 1 9 1 9 0 2 4 13 16 13 1 4 13 1 0 9 2
33 10 9 13 1 10 9 0 1 13 15 3 13 10 9 2 16 15 3 13 16 15 15 4 13 4 4 13 1 9 1 10 0 2
20 10 9 15 4 13 10 9 13 3 4 13 10 9 1 9 1 10 10 9 2
31 10 9 3 4 13 10 9 13 1 9 1 15 3 4 13 2 3 16 13 1 13 10 9 13 1 9 1 15 4 13 2
24 10 9 15 4 13 10 9 1 0 9 4 13 15 2 0 10 9 1 10 9 1 10 9 2
23 15 13 10 9 1 10 0 9 1 10 0 9 4 13 2 16 13 2 10 9 13 13 2
16 1 9 1 10 9 2 10 9 4 4 13 1 10 9 13 2
28 10 9 3 4 13 10 9 1 10 9 2 3 1 1 10 9 7 1 10 9 2 1 10 9 1 10 9 2
18 10 9 13 1 9 1 9 7 1 9 4 4 13 3 1 10 9 2
12 10 9 1 10 9 13 1 9 1 10 9 2
28 10 9 3 4 13 15 13 10 9 0 1 15 13 2 3 16 1 9 0 7 0 2 3 16 10 9 13 2
12 1 10 9 3 13 10 9 13 1 10 15 2
32 16 1 9 1 10 9 4 13 10 9 2 10 9 15 13 1 10 9 1 10 9 2 16 3 13 10 0 9 1 10 9 2
14 13 0 15 4 13 1 10 0 9 1 10 9 12 2
36 10 9 15 13 10 9 4 2 1 9 7 1 9 1 10 9 2 13 9 7 13 15 9 1 10 9 2 16 15 3 4 13 1 10 9 2
16 10 9 1 10 9 1 10 9 13 13 10 9 1 10 9 2
34 10 9 15 4 13 10 9 4 13 10 9 1 10 9 1 10 9 0 13 1 10 9 7 1 10 0 9 15 3 15 13 10 9 2
19 10 9 2 13 10 9 1 10 15 2 4 2 13 15 1 10 10 9 2
21 10 9 13 1 10 0 9 13 9 3 1 10 15 15 4 13 9 1 10 9 2
21 16 10 9 4 13 1 9 2 15 13 10 9 1 10 0 9 1 10 9 12 2
31 16 10 9 13 0 2 10 0 13 7 10 9 13 1 10 9 1 10 9 1 9 1 15 4 15 13 2 0 9 0 2
25 16 10 9 13 1 9 2 13 1 10 9 10 9 1 10 9 13 1 9 3 0 1 10 9 2
21 3 4 3 13 10 9 7 10 9 1 10 9 15 3 4 4 13 1 10 9 2
30 10 9 4 3 13 1 13 10 9 13 1 10 10 9 7 1 13 10 9 1 10 9 7 10 9 1 10 9 13 2
33 10 9 1 10 9 15 13 1 10 9 1 10 9 2 16 15 4 3 13 0 1 9 13 1 9 7 16 4 13 1 10 9 2
32 10 9 4 13 10 9 1 10 9 1 10 9 0 1 13 10 9 1 10 9 0 7 1 0 9 15 3 15 13 10 9 2
28 16 10 9 13 1 9 9 9 1 9 7 9 0 1 13 1 10 9 1 10 9 2 10 9 4 13 0 2
42 16 15 13 3 1 9 0 1 13 1 9 0 2 10 9 13 1 10 9 1 10 9 1 13 15 2 13 1 9 1 15 13 1 10 9 13 1 10 9 1 9 2
29 16 10 9 13 1 13 10 9 0 7 3 15 13 1 13 10 9 13 15 1 9 2 10 9 4 13 10 9 2
36 13 10 9 2 16 15 4 13 1 10 9 7 4 13 0 1 9 13 1 9 2 10 9 3 4 3 13 15 7 4 13 1 10 10 9 2
31 10 9 3 13 9 16 10 9 15 13 3 16 4 4 13 1 10 9 7 3 16 4 4 13 0 1 9 13 1 9 2
20 16 10 9 0 7 10 9 13 0 2 10 9 13 13 1 9 1 10 9 2
21 16 4 4 13 10 9 2 10 9 13 1 10 9 1 10 9 1 13 15 9 2
18 10 9 4 4 13 1 10 9 13 1 10 0 9 1 10 9 12 2
20 10 9 1 10 9 1 10 9 2 4 13 1 10 9 10 9 1 10 9 2
20 1 10 9 15 4 13 1 10 9 1 15 4 13 1 10 9 10 9 13 2
37 16 10 9 13 1 10 13 2 10 9 4 13 1 9 1 10 9 1 13 10 9 7 1 13 10 9 15 13 1 9 10 0 1 13 15 0 2
11 10 9 4 4 13 1 10 9 1 9 2
43 10 9 15 3 13 3 10 9 13 4 13 1 10 9 1 10 9 2 16 3 13 16 10 9 7 10 9 4 4 13 1 9 1 10 9 13 1 9 1 15 3 0 2
14 10 9 4 13 1 9 1 9 7 9 13 1 9 2
39 16 10 9 13 1 10 9 1 10 9 2 10 9 3 4 13 1 9 15 1 9 7 9 13 1 9 2 7 13 12 9 1 10 9 7 1 10 9 2
47 10 9 3 4 4 13 1 9 2 16 3 4 13 9 1 10 9 13 2 3 1 13 10 9 13 1 10 9 0 1 10 0 9 2 1 3 16 10 9 15 4 13 1 10 9 0 2
40 10 9 15 13 1 9 3 4 13 1 10 13 9 1 10 9 13 1 9 1 15 3 0 2 16 3 13 16 10 9 1 10 9 4 3 13 1 10 9 2
31 1 10 9 4 13 7 13 10 9 3 13 2 10 9 1 15 3 13 15 15 4 13 1 10 9 1 13 15 10 9 2
15 10 9 1 10 9 3 15 13 1 10 9 1 3 13 2
13 10 9 13 1 9 1 15 13 1 1 15 9 2
35 10 9 1 10 9 1 10 9 7 1 10 9 4 13 3 10 9 13 1 10 9 1 10 0 9 2 1 3 15 13 9 0 7 0 2
25 16 1 1 10 9 4 13 9 1 9 0 1 15 0 2 10 9 0 4 13 1 10 0 9 2
16 1 10 9 15 13 1 13 13 10 9 0 13 10 0 9 2
15 15 3 4 13 16 4 4 13 10 9 1 10 9 0 2
35 16 10 9 7 10 9 3 13 1 9 1 10 9 2 10 9 4 13 1 10 9 15 4 13 15 1 10 9 1 15 4 13 10 9 2
22 16 10 9 3 4 4 13 1 10 10 0 9 2 4 13 1 10 9 1 9 0 2
35 16 10 9 0 1 10 9 4 13 1 13 10 9 2 10 9 4 13 1 10 9 1 10 9 7 10 9 1 10 9 15 15 4 13 2
19 10 9 3 4 13 1 10 9 15 10 9 4 4 13 13 10 0 9 2
21 13 0 10 9 15 13 7 13 3 10 9 1 10 9 1 9 7 1 9 0 2
39 13 0 3 10 9 0 1 9 7 1 9 1 9 1 10 9 1 15 10 9 1 10 9 7 1 10 10 9 13 9 1 9 13 1 9 1 9 0 2
21 10 9 15 13 16 10 9 13 1 10 9 0 10 0 9 1 9 7 9 0 2
14 10 9 1 13 10 9 0 4 13 1 9 3 0 2
30 10 9 1 10 9 7 10 10 9 2 10 9 7 10 9 1 10 9 7 10 0 9 0 1 10 9 3 13 9 2
30 10 9 2 10 9 7 10 9 2 1 10 9 0 15 13 2 16 10 9 3 13 3 1 13 15 1 10 0 9 2
13 10 9 13 1 9 2 16 3 13 10 9 0 2
31 16 10 9 0 13 1 10 9 0 2 10 9 13 0 16 10 9 4 13 3 10 0 9 13 10 9 1 10 9 0 2
26 16 10 0 9 4 13 1 15 0 15 4 13 2 15 13 10 9 0 1 10 9 0 1 10 9 2
33 10 9 1 10 9 1 13 10 9 13 10 9 16 4 13 1 10 9 2 3 16 15 13 1 10 0 9 1 3 4 15 13 2
31 16 10 9 1 10 9 13 1 9 0 2 10 9 0 1 10 9 13 1 9 0 13 13 10 9 2 0 10 9 0 2
17 10 9 1 10 9 1 10 9 3 13 13 10 9 1 10 9 2
11 10 9 13 1 10 9 0 13 10 9 2
21 10 9 13 1 15 1 10 9 3 13 10 15 16 1 10 9 1 10 9 13 2
45 10 9 15 4 13 2 1 9 2 1 10 9 13 1 10 15 4 13 1 10 9 0 15 4 13 2 1 9 1 10 9 7 1 15 15 4 13 9 1 10 9 1 10 9 2
14 10 9 13 10 12 9 1 10 9 1 10 10 9 2
9 10 9 3 4 13 15 1 9 2
22 10 9 3 13 10 9 2 16 3 4 13 16 15 4 13 10 9 1 10 12 9 2
15 10 9 13 3 1 10 9 3 13 1 9 1 10 9 2
27 16 10 12 9 3 13 0 1 10 0 9 2 15 4 13 10 9 1 10 9 1 10 9 1 10 9 2
17 10 9 4 13 1 9 10 9 15 10 9 13 1 10 9 0 2
16 10 0 9 13 1 10 15 15 4 13 10 9 7 10 9 2
25 10 9 3 13 1 10 9 2 7 1 15 13 2 13 10 9 1 10 9 13 3 1 10 9 2
27 16 10 9 13 1 10 15 10 9 0 2 15 13 1 10 9 10 9 1 10 0 9 1 10 9 12 2
21 1 9 1 10 9 4 13 9 9 3 16 3 13 10 9 13 1 10 9 0 2
12 10 9 4 3 13 3 10 9 1 10 9 2
33 16 10 9 1 9 7 1 9 15 13 1 10 0 9 2 10 9 15 13 2 7 10 0 15 4 13 9 1 10 9 4 13 2
22 10 9 3 13 1 9 1 10 15 15 4 13 9 1 9 7 1 9 1 10 9 2
29 16 1 10 0 9 15 13 10 9 1 9 7 1 9 0 2 10 9 13 1 9 2 16 10 9 15 13 9 2
20 10 9 15 13 16 2 1 10 9 3 0 1 10 9 2 10 9 13 0 2
24 16 10 9 13 3 0 2 10 9 2 16 15 13 2 3 13 0 1 10 9 1 10 9 2
28 10 9 15 13 1 9 10 9 0 15 13 13 0 3 16 10 9 4 13 1 16 4 4 15 13 10 9 2
28 16 10 9 4 13 0 3 1 9 2 10 9 15 13 1 10 9 13 10 9 1 10 9 15 4 13 0 2
39 10 9 4 13 1 9 0 7 0 10 10 9 2 3 1 10 9 1 10 9 2 16 10 9 3 13 9 3 0 7 10 9 3 4 13 1 10 9 2
10 10 9 4 13 10 9 1 10 9 2
25 7 10 9 3 13 0 1 10 9 2 16 3 15 13 16 15 15 13 1 10 9 1 10 9 2
36 10 9 1 10 9 0 3 15 13 1 10 9 1 9 0 1 9 2 7 1 15 13 1 9 1 9 7 1 9 1 9 13 1 10 9 2
29 1 9 1 10 9 2 10 9 4 13 1 10 9 1 10 9 2 1 10 9 0 7 0 7 1 10 0 9 2
12 0 9 0 2 10 9 3 13 10 9 13 2
23 10 9 13 9 1 10 9 1 10 9 13 16 15 15 4 13 7 16 15 4 4 13 2
19 10 0 9 15 13 16 10 9 4 13 9 1 9 1 9 7 1 9 2
36 16 10 9 13 1 9 0 2 10 9 4 13 3 1 10 9 7 1 10 9 1 15 10 9 13 1 9 1 10 13 10 9 1 10 9 2
13 1 10 9 15 13 1 10 9 1 15 4 13 2
28 4 3 13 10 9 2 13 10 9 1 10 9 7 15 15 10 9 4 13 1 13 10 9 7 13 10 9 2
40 16 10 9 13 1 10 9 10 0 9 2 10 15 15 13 1 10 9 2 10 9 0 3 4 13 1 10 10 9 2 3 16 10 9 13 3 1 13 15 2
30 3 10 9 15 4 13 10 9 1 10 15 3 4 13 15 1 10 13 2 16 3 3 4 13 1 10 9 10 9 2
28 16 10 9 1 13 10 9 4 13 10 15 2 15 4 13 15 1 10 9 2 3 16 10 9 15 4 13 2
22 10 15 13 1 13 10 9 3 4 13 1 13 10 9 2 16 13 9 1 10 13 2
33 10 13 4 13 10 9 2 3 1 16 10 9 3 4 13 10 9 1 9 1 10 9 7 3 4 13 10 9 1 9 1 15 2
27 10 9 4 13 10 9 7 13 10 9 1 9 1 10 9 3 1 10 9 7 10 0 9 1 10 13 2
17 10 9 4 13 1 10 9 10 9 0 1 10 10 9 1 15 2
30 10 9 3 4 3 13 10 9 0 1 10 9 1 10 13 7 10 9 2 16 1 15 10 9 3 4 13 0 9 2
27 16 3 15 4 13 3 2 10 0 3 4 13 1 10 9 10 9 0 1 10 10 9 1 10 9 0 2
34 4 13 15 3 10 9 15 1 10 9 4 4 13 10 9 0 2 16 3 13 0 1 10 15 7 3 13 1 9 0 1 10 9 2
23 3 4 13 15 10 9 15 4 4 13 10 9 0 2 16 15 4 13 1 1 10 9 2
6 10 9 1 10 9 0
2 9 0
3 9 12 2
12 10 11 13 10 9 0 2 0 1 10 9 2
21 10 9 13 1 10 9 2 15 15 13 1 10 9 7 1 10 9 1 10 9 2
3 9 12 2
43 10 9 13 7 13 10 9 0 1 10 9 2 7 1 9 7 1 10 9 0 3 15 13 10 10 9 2 7 13 10 9 1 10 9 0 1 9 0 2 0 7 0 2
3 9 12 2
39 10 10 9 13 0 9 0 7 13 0 3 1 10 9 2 1 9 1 9 2 1 9 2 1 9 2 1 9 2 1 9 0 2 1 9 0 7 0 2
56 13 9 1 10 9 13 10 9 1 9 0 7 0 2 15 2 13 1 9 10 9 7 10 9 1 10 9 2 13 10 0 9 1 10 9 0 7 10 0 9 1 10 10 9 1 10 9 0 2 0 7 0 1 10 9 2
3 9 12 2
22 10 9 13 1 10 10 9 10 9 1 10 9 7 13 10 9 15 13 0 10 9 2
34 10 9 13 10 9 1 13 2 1 10 10 9 7 10 10 9 2 10 9 7 10 9 15 13 1 10 9 0 7 0 1 10 9 2
3 9 12 2
14 10 9 2 0 7 0 2 13 7 13 10 9 0 2
15 13 1 10 9 15 13 1 10 9 10 3 0 9 0 2
21 13 10 9 7 10 9 1 10 10 9 1 10 9 1 10 9 7 1 10 9 2
3 9 12 2
10 10 9 13 1 0 9 10 9 0 2
3 9 12 2
18 10 9 7 10 9 0 13 2 15 1 10 10 9 2 0 7 0 2
10 10 10 9 4 13 1 10 9 0 2
18 10 9 1 10 9 13 1 10 12 9 2 3 13 9 1 9 0 2
3 9 12 2
12 10 10 9 0 13 3 0 3 1 10 9 2
27 10 9 0 0 1 10 0 13 9 1 13 15 1 10 10 9 2 1 3 3 13 1 10 9 0 0 2
20 10 10 9 1 10 9 4 13 1 9 1 10 9 1 9 1 10 0 9 2
3 9 12 2
15 10 9 13 10 9 1 10 9 7 10 9 0 7 0 2
13 13 10 9 7 10 9 0 7 0 1 10 9 2
3 9 12 2
22 10 9 0 1 10 9 4 13 1 10 9 1 9 1 10 9 7 1 10 9 0 2
43 10 9 2 1 10 15 4 13 1 10 10 9 10 0 9 1 10 9 0 13 1 10 9 0 2 13 9 1 9 1 10 9 1 10 9 1 10 9 13 1 10 9 2
12 3 4 13 10 9 1 10 9 1 9 0 2
3 9 12 2
26 10 11 13 10 9 1 9 1 9 1 10 9 1 10 0 9 7 1 9 1 9 1 10 9 0 2
31 13 2 1 9 1 9 1 10 0 9 2 1 10 9 1 9 0 1 10 9 15 13 10 9 7 10 9 1 10 9 2
11 13 7 13 10 9 0 13 1 10 9 2
3 9 12 2
24 10 9 1 10 9 13 10 9 0 2 0 2 0 7 0 2 1 12 9 0 1 0 9 2
2 9 0
7 9 7 9 1 10 9 2
2 9 0
2 9 0
3 9 12 2
6 10 9 0 13 0 2
44 3 4 13 9 10 1 9 2 1 9 7 9 0 2 7 10 0 9 1 10 9 0 2 16 3 1 9 0 1 10 9 0 7 1 10 0 9 7 9 13 1 10 9 2
58 1 9 0 1 9 7 9 2 13 3 1 10 9 2 10 9 1 0 9 4 13 9 0 2 15 4 4 13 1 12 9 1 10 9 0 7 2 16 15 3 15 13 1 10 0 12 9 2 15 13 13 7 13 0 1 10 9 2
17 4 13 10 9 0 7 0 1 10 9 3 13 1 9 1 9 2
11 10 9 13 10 9 0 1 10 9 0 2
3 9 12 2
5 10 9 13 0 2
34 3 15 15 4 13 9 7 9 7 9 2 16 3 1 10 9 7 9 13 1 10 9 1 10 9 13 1 10 9 1 10 9 0 2
3 9 12 2
18 10 9 7 10 9 1 10 9 7 1 10 0 9 1 9 13 0 2
21 10 10 9 4 13 3 1 9 0 1 10 9 0 1 10 9 13 1 10 9 2
3 9 12 2
33 10 9 4 13 7 13 3 1 10 9 1 10 9 0 2 1 10 9 15 10 9 13 1 9 0 1 9 1 9 7 1 9 2
9 10 9 4 4 13 1 9 0 2
23 10 9 13 0 1 13 1 10 9 1 10 9 7 1 13 15 2 1 10 9 1 9 2
3 9 12 2
12 10 9 13 9 1 13 15 3 7 1 9 2
17 1 10 9 2 3 1 9 0 1 10 9 2 3 4 13 9 2
29 1 10 9 1 9 0 4 4 13 9 1 10 9 2 15 4 13 15 3 1 13 9 1 9 7 1 9 0 2
3 9 12 2
26 10 9 13 9 1 13 15 3 2 1 9 2 1 9 15 3 4 13 1 10 9 1 10 9 0 2
21 4 13 10 9 0 7 15 15 13 2 3 3 2 9 0 1 9 1 9 0 2
3 9 12 2
46 15 13 9 1 13 3 10 10 9 0 1 10 9 2 0 7 13 2 1 13 15 9 7 1 13 15 1 9 7 1 9 10 9 2 16 3 15 13 1 9 0 1 10 0 9 2
3 9 12 2
43 10 9 0 7 10 9 1 9 7 1 9 1 10 9 7 9 3 4 13 9 1 0 9 0 2 7 1 0 9 0 1 10 10 9 2 9 0 7 10 9 1 9 2
3 9 12 2
22 15 13 9 1 13 3 10 10 9 1 10 9 2 10 9 7 10 0 9 1 9 2
11 10 9 3 4 13 0 1 9 7 9 2
54 1 10 9 2 16 15 13 0 9 7 3 13 0 10 0 9 1 10 9 0 2 10 9 1 10 9 0 4 4 13 1 9 1 9 0 2 15 4 3 2 7 3 3 1 12 9 2 13 9 1 10 9 0 2
22 16 15 3 15 13 1 10 12 9 0 2 10 9 15 13 13 7 0 1 10 9 2
24 10 9 4 13 2 1 9 1 9 0 2 16 4 13 0 10 9 1 9 1 10 9 0 2
20 4 13 10 9 1 9 2 10 9 7 10 10 0 9 0 1 10 0 9 2
13 10 9 13 9 0 1 13 7 1 13 10 9 2
3 9 12 2
22 15 4 4 13 2 1 9 0 2 1 10 9 0 2 1 10 9 2 1 10 9 2
3 9 12 2
16 10 9 0 7 0 4 4 13 16 3 1 9 1 10 9 2
3 9 12 2
16 15 4 13 1 9 1 10 9 1 10 10 9 7 9 0 2
23 4 13 1 10 3 0 2 1 0 9 2 10 9 1 13 7 13 15 3 1 10 9 2
16 10 9 13 10 9 7 10 9 1 10 9 1 10 9 0 2
3 9 12 2
12 15 4 4 13 1 10 9 0 13 1 9 2
22 15 4 4 13 16 3 1 9 1 10 9 15 4 13 1 9 3 1 10 9 13 2
18 15 4 4 13 1 9 1 9 16 3 1 10 9 13 1 10 9 2
3 9 12 2
18 10 9 1 10 9 4 4 13 3 16 4 3 13 1 10 9 0 2
11 3 4 1 10 9 4 13 1 9 0 2
3 9 12 2
6 10 9 0 13 0 2
23 10 9 3 4 13 1 9 0 1 10 9 1 9 7 4 13 1 10 9 1 10 9 2
8 3 4 13 10 9 1 9 2
3 9 12 2
35 10 9 7 10 9 1 10 9 7 1 10 9 0 13 3 0 2 1 10 9 0 2 0 7 0 2 1 10 9 13 1 9 1 9 2
17 1 10 9 10 9 0 15 13 1 10 9 7 1 10 9 0 2
2 9 0
3 9 12 2
16 10 9 13 10 9 1 10 9 1 9 0 0 1 10 9 2
28 10 9 4 13 1 10 9 0 7 0 1 10 9 2 1 10 9 13 1 10 9 1 9 1 10 9 0 2
3 9 12 2
23 13 9 7 9 1 10 9 13 2 13 7 13 10 9 2 3 16 13 3 1 10 9 2
20 1 10 9 1 9 1 10 9 2 10 9 13 1 16 4 13 10 10 9 2
29 10 9 13 1 10 9 13 3 1 10 9 10 9 0 7 0 2 0 1 10 9 1 10 9 1 10 9 0 2
15 10 9 13 10 9 7 10 9 1 10 9 1 10 9 2
3 9 12 2
3 9 12 2
25 10 9 13 10 9 1 0 9 1 10 9 7 9 1 10 9 2 7 13 9 0 1 10 0 2
16 15 4 4 13 1 10 0 9 0 16 3 1 9 1 9 2
19 10 9 3 4 1 10 9 13 10 9 13 1 10 9 1 10 9 0 2
3 9 12 2
14 10 9 7 10 9 13 0 7 0 15 13 10 9 2
20 10 9 13 10 9 0 1 10 9 7 13 9 0 1 10 10 9 7 9 2
45 10 9 2 1 10 13 10 9 7 10 9 1 10 9 3 0 15 13 10 9 2 4 13 1 15 0 9 7 1 10 10 9 10 9 0 0 1 15 1 10 9 1 9 0 2
32 4 13 10 9 1 9 1 10 9 1 10 0 9 7 9 1 9 7 1 10 9 1 15 7 1 10 9 1 10 9 0 2
29 10 9 1 0 9 2 9 7 9 2 13 10 9 1 13 15 9 0 1 10 9 13 1 10 9 1 10 9 2
3 9 12 2
7 10 9 13 0 1 15 2
15 10 9 0 2 13 1 3 12 9 2 13 0 7 0 2
23 10 0 7 0 2 3 16 0 1 9 2 13 9 1 13 10 9 3 0 1 10 9 2
26 10 9 13 0 10 9 1 9 1 9 2 9 1 10 9 7 0 9 2 15 4 4 13 1 9 2
2 9 0
2 9 0
3 9 12 2
13 10 9 13 10 9 1 10 10 10 9 7 9 2
11 13 10 9 7 10 9 0 1 10 9 2
27 13 10 9 1 9 2 1 10 9 13 1 10 9 1 10 9 0 2 7 13 10 9 0 1 10 9 2
3 9 12 2
36 10 9 13 9 1 10 9 0 1 10 9 7 9 1 10 10 9 7 1 10 9 0 1 13 1 15 7 1 10 9 10 9 0 7 0 2
13 10 9 0 1 10 9 0 4 13 1 10 9 2
20 10 9 13 9 1 10 9 0 7 1 9 0 13 2 7 3 4 13 15 2
3 9 12 2
23 10 9 0 13 10 0 9 7 2 1 9 1 9 2 10 0 9 15 13 1 10 9 2
28 10 9 1 9 4 13 10 9 1 10 10 0 9 0 7 13 1 10 9 7 1 10 9 10 0 0 9 2
13 10 9 13 10 9 0 1 9 1 10 9 0 2
29 10 9 13 10 9 1 10 9 1 0 9 7 13 1 15 2 1 9 1 9 2 10 9 1 10 9 1 9 2
3 9 12 2
25 10 9 0 1 10 9 7 0 1 10 9 0 1 13 13 9 1 10 9 7 1 10 9 0 2
31 10 9 13 9 16 4 13 7 13 9 0 1 10 10 9 1 9 1 9 1 9 2 9 2 9 7 9 2 9 0 2
18 1 10 9 13 1 10 9 13 9 7 9 13 7 13 1 10 9 2
6 10 9 0 13 0 2
3 9 12 2
6 10 9 0 13 0 2
26 1 10 9 3 4 4 13 0 9 16 3 10 10 9 1 9 0 7 0 2 1 10 9 1 9 2
19 13 9 1 10 9 16 10 9 1 10 9 13 10 9 0 1 9 0 2
7 10 9 13 13 9 0 2
34 4 2 13 3 1 9 1 10 10 9 2 13 9 0 1 9 1 9 0 1 10 10 13 1 10 9 1 10 15 10 9 15 13 2
3 9 12 2
16 10 9 1 9 15 13 1 10 9 1 10 9 15 15 13 2
3 9 12 2
7 10 9 0 0 13 0 2
29 3 4 13 15 1 9 1 10 9 0 7 1 9 1 13 9 1 10 9 2 1 10 9 2 1 10 9 0 2
25 10 9 13 10 9 7 10 9 0 16 10 9 0 0 7 0 4 4 13 7 13 1 9 0 2
3 9 12 2
7 10 9 13 0 7 0 2
14 10 9 0 13 1 10 9 2 1 9 7 1 9 2
41 10 9 0 4 13 7 13 1 10 9 2 15 15 13 10 9 1 9 2 1 9 7 10 9 1 10 9 1 13 15 10 9 0 7 1 13 15 0 1 15 2
25 10 9 0 4 4 2 1 10 9 13 1 10 9 2 7 1 9 2 13 1 9 1 9 0 2
24 10 9 13 10 9 7 10 9 1 10 9 0 7 0 7 10 9 1 10 9 1 10 9 2
3 9 12 2
66 1 9 1 9 0 10 9 4 13 3 7 13 2 1 9 7 1 9 2 1 10 9 2 1 9 0 7 1 9 1 9 7 1 9 10 9 7 9 1 9 2 15 15 13 1 9 0 0 7 1 9 1 9 7 1 9 1 9 7 13 9 1 0 9 0 2
3 9 12 2
66 1 10 9 1 13 10 0 9 1 10 9 7 1 13 0 9 0 2 10 9 13 9 7 9 1 10 9 0 0 2 13 9 1 10 10 9 1 10 9 7 10 9 0 2 13 7 13 10 9 1 10 9 2 10 9 1 10 9 7 10 9 1 10 9 0 2
11 10 9 13 9 1 9 1 10 9 0 2
3 9 12 2
20 10 9 13 10 9 0 1 10 9 1 9 1 9 7 1 9 1 9 0 2
28 10 9 15 13 7 13 10 9 1 10 9 3 0 7 15 13 2 1 10 0 9 2 10 9 7 10 9 2
14 10 9 13 1 10 9 7 1 10 9 1 10 9 2
3 9 12 2
51 1 10 9 1 10 9 0 7 0 1 10 9 1 9 1 10 9 1 10 9 2 10 9 13 10 9 1 10 9 1 13 2 1 10 9 7 1 10 9 13 1 10 9 2 1 10 9 1 10 9 2
3 9 12 2
13 10 9 13 7 13 10 9 1 10 10 10 9 2
11 13 2 13 7 13 10 9 1 10 9 2
36 13 10 9 1 10 9 0 1 10 9 1 10 9 2 1 10 9 0 0 7 1 10 0 7 0 9 0 1 10 0 9 0 1 10 9 2
2 9 0
2 9 0
3 9 12 2
17 13 9 10 10 9 2 9 7 9 2 15 4 13 10 0 9 2
11 10 9 13 0 7 0 2 0 7 0 2
7 10 10 9 13 9 0 2
27 10 9 13 9 7 9 1 10 9 1 10 9 1 9 1 10 9 0 1 10 9 7 15 13 10 9 2
36 1 10 9 4 13 10 9 11 1 10 9 1 10 9 2 1 10 15 4 13 9 1 10 9 13 1 9 0 7 1 9 13 1 10 9 2
3 9 12 2
22 10 10 9 13 9 1 13 15 3 1 9 1 13 1 9 0 1 13 10 9 0 2
3 9 12 2
18 10 10 9 4 13 9 1 10 9 1 13 9 0 7 13 0 9 2
3 9 12 2
35 10 10 9 1 10 15 7 1 10 0 9 4 13 1 10 9 0 7 1 10 9 0 1 9 1 9 2 1 10 9 13 1 10 9 2
17 1 10 9 10 9 13 1 0 9 10 0 9 1 9 7 9 2
29 10 9 4 2 1 10 9 1 10 0 9 7 1 10 9 0 2 13 1 10 9 10 9 3 13 1 10 9 2
28 15 4 13 1 9 0 0 13 9 1 13 1 10 9 0 1 10 10 9 7 1 13 10 10 9 1 9 2
3 9 12 2
12 10 9 1 10 9 13 0 9 1 10 9 2
15 10 9 0 13 0 1 10 9 7 9 13 1 10 9 2
21 10 10 9 3 13 10 9 1 9 1 10 9 2 7 10 9 1 10 9 0 2
16 10 9 1 10 9 0 15 13 1 10 9 0 1 10 9 2
3 9 12 2
17 15 4 13 1 13 1 10 9 0 1 9 1 10 10 9 0 2
10 10 9 0 4 13 1 9 1 9 2
3 9 12 2
22 10 10 9 13 10 9 1 13 0 1 10 9 7 1 13 15 10 9 7 10 9 2
28 10 9 15 4 13 9 0 13 10 9 1 13 15 1 9 7 9 2 13 9 1 10 9 13 1 10 9 2
2 9 0
4 9 1 10 9
2 9 0
2 10 9
2 9 0
2 10 9
3 9 12 2
18 10 9 15 13 1 10 9 1 10 9 7 1 10 9 1 10 9 2
23 10 9 15 13 1 9 0 1 10 9 1 10 12 9 1 10 0 9 13 1 10 9 2
3 9 12 2
13 10 9 1 10 9 4 13 1 9 0 7 0 2
19 10 9 1 10 9 13 1 12 2 12 1 10 15 13 1 10 9 11 2
74 10 9 1 10 9 1 10 9 2 13 0 10 9 1 10 9 13 1 10 9 11 2 15 13 13 10 9 1 10 9 1 10 9 2 15 13 1 10 0 9 0 1 10 9 2 1 12 7 13 10 9 1 9 1 10 9 1 10 9 2 1 10 9 1 10 9 0 7 1 10 3 0 9 2
3 9 12 2
20 10 9 1 10 9 4 13 1 9 0 2 0 10 9 13 1 10 9 11 2
20 10 9 1 10 9 0 13 1 12 2 12 1 10 15 13 1 10 9 11 2
12 10 9 4 13 10 9 1 9 0 1 12 2
12 10 11 15 13 12 2 10 11 1 11 12 2
65 10 9 1 10 9 1 10 9 2 13 0 10 9 1 10 9 13 1 10 9 11 2 0 9 1 10 9 1 10 0 9 2 15 13 1 9 1 10 9 1 10 9 2 15 13 1 10 0 9 0 2 1 10 9 1 10 9 0 7 1 10 3 0 9 2
3 9 12 2
21 10 9 4 13 1 9 0 7 0 1 10 9 15 4 13 10 0 9 1 9 2
13 13 0 1 9 10 9 15 4 13 10 0 9 2
3 9 12 2
19 13 9 1 9 7 1 9 2 1 9 2 15 4 13 9 1 10 9 2
31 10 9 1 10 9 4 13 9 1 9 12 9 15 4 13 10 9 1 0 9 1 10 9 0 2 0 2 0 7 0 2
3 9 12 2
17 10 9 1 10 9 7 10 9 1 10 9 4 13 1 12 9 2
20 10 9 1 10 9 3 4 4 13 16 3 1 9 7 3 1 9 1 9 2
3 9 12 2
18 10 9 1 10 0 9 13 9 1 12 9 1 10 9 1 10 0 2
14 10 0 9 13 9 3 1 10 0 9 1 10 9 2
15 16 3 4 13 10 0 9 4 13 10 9 1 10 0 2
3 9 12 2
17 10 9 15 13 1 9 10 0 9 3 0 1 9 7 1 9 2
30 10 11 4 4 13 1 9 0 1 9 1 10 10 9 7 1 10 9 1 10 9 7 1 10 15 1 10 10 9 2
17 16 15 13 1 9 0 10 11 2 4 13 1 9 3 10 15 2
3 9 12 2
15 10 11 13 1 10 10 9 10 9 7 10 9 1 9 2
25 16 10 9 15 13 1 9 0 2 10 9 7 10 9 1 9 13 15 1 10 9 1 10 9 2
3 9 12 2
14 10 9 13 10 10 9 1 9 0 1 10 10 9 2
5 10 9 13 0 2
21 3 15 1 10 12 9 7 10 9 1 9 13 4 13 1 13 15 1 9 0 2
43 10 9 1 10 9 7 1 10 9 3 13 0 16 3 13 0 10 9 1 10 10 9 2 7 16 3 4 13 1 9 1 10 9 2 3 16 10 9 13 10 9 0 2
29 10 9 1 10 9 2 3 16 3 13 9 1 10 9 2 13 9 2 7 16 13 9 2 1 13 1 10 9 2
9 4 4 13 10 9 16 15 13 2
3 9 12 2
18 10 9 13 10 9 1 9 7 9 1 10 9 1 9 7 1 9 2
9 15 4 13 3 1 10 12 9 2
3 9 12 2
23 10 9 13 1 10 9 1 9 1 10 10 9 7 1 10 9 13 1 9 7 1 9 2
3 9 12 2
18 10 9 1 10 9 13 10 9 7 13 10 10 9 1 9 1 9 2
3 9 12 2
28 10 9 1 10 9 3 4 4 13 1 13 1 10 9 13 7 1 10 9 13 1 10 9 1 10 10 9 2
74 1 9 1 10 9 1 10 15 13 2 10 9 1 10 9 4 4 13 1 9 0 7 0 2 7 4 4 13 7 3 13 1 10 9 0 2 7 13 1 9 2 3 16 1 9 1 10 9 0 1 9 2 7 16 4 13 1 10 9 1 13 10 9 1 10 15 4 13 10 9 0 1 9 2
28 0 9 4 13 1 13 10 9 1 10 9 1 9 2 1 10 9 2 1 9 7 9 7 1 9 1 9 2
3 9 12 2
13 10 9 1 10 9 13 10 9 13 1 10 9 2
2 9 0
5 10 9 1 10 9
3 9 12 2
11 10 9 0 4 13 3 1 10 12 9 2
3 9 12 2
31 10 9 1 10 9 13 1 10 9 2 1 10 9 1 10 9 7 1 10 9 7 9 1 10 15 4 13 1 9 0 2
27 10 9 13 10 9 1 10 9 2 1 10 9 2 1 9 1 3 12 9 2 1 10 9 13 1 9 2
3 9 12 2
41 10 9 1 9 2 13 1 10 9 4 2 1 10 9 1 10 10 9 2 13 1 10 9 7 3 1 10 9 0 2 15 15 13 9 1 9 7 1 9 0 2
18 10 9 13 9 0 1 10 9 1 9 1 10 15 4 13 10 9 2
38 4 3 13 1 10 9 7 9 10 9 7 10 9 1 10 9 1 9 4 13 1 9 2 3 0 2 13 1 9 1 13 10 9 1 10 9 0 2
68 3 1 10 9 2 3 1 10 9 1 10 10 9 0 2 10 9 1 9 4 13 1 10 9 2 16 10 9 7 10 15 1 10 9 1 10 11 7 10 15 1 10 9 13 16 4 13 7 13 1 10 9 0 7 16 4 13 1 10 10 9 0 1 0 9 1 9 2
14 10 9 13 10 9 1 9 1 10 9 1 10 9 2
48 10 9 0 1 9 7 1 9 0 1 9 1 10 9 4 3 13 1 10 9 1 9 1 9 0 7 0 7 1 15 1 9 0 2 1 9 1 13 9 0 2 1 9 1 9 7 9 2
3 9 12 2
17 10 9 4 13 1 10 9 1 10 9 1 10 9 1 10 9 2
29 16 10 9 2 15 1 9 0 1 10 10 9 2 15 13 10 9 2 10 9 4 13 1 10 9 1 15 13 2
31 10 9 4 13 3 1 10 9 7 13 1 9 10 0 9 0 1 10 10 9 2 3 16 10 9 0 13 10 9 0 2
3 9 12 2
24 10 9 1 10 9 2 3 1 13 10 9 2 4 1 9 0 1 10 9 13 10 0 9 2
13 16 10 9 13 3 10 9 2 15 4 4 13 2
3 9 12 2
35 4 13 9 0 1 13 10 9 2 0 7 0 2 1 10 9 7 1 10 9 13 9 1 9 2 16 15 13 12 9 7 12 9 0 2
26 3 4 13 10 9 1 10 9 0 7 1 9 2 1 9 7 1 9 2 1 9 1 13 9 0 2
19 13 9 1 13 1 10 9 10 10 9 13 1 13 10 9 1 10 9 2
32 10 9 0 1 9 4 13 16 4 13 1 10 9 10 9 1 10 13 9 2 7 16 4 13 10 9 1 10 9 3 13 2
11 10 9 13 10 9 1 9 1 10 9 2
3 9 12 2
32 10 9 1 10 9 0 3 4 4 13 1 10 9 16 3 1 9 1 9 7 9 0 7 3 1 9 13 7 1 9 13 2
3 9 12 2
20 10 9 3 4 2 1 9 1 10 9 2 13 9 15 13 9 1 9 0 2
55 16 2 1 9 0 1 9 7 1 9 2 10 9 13 2 1 10 10 9 2 9 0 1 9 1 9 2 4 10 9 0 13 15 1 10 9 1 10 9 15 2 3 16 13 2 4 3 13 7 15 13 1 12 9 2
23 10 9 13 9 3 1 10 9 2 16 3 4 13 1 9 1 12 9 1 10 10 9 2
20 10 9 4 3 13 1 9 10 9 0 13 1 10 9 1 10 9 3 13 2
3 9 12 2
16 10 9 13 10 9 1 9 7 13 1 10 9 10 9 0 2
3 9 12 2
33 10 9 7 10 9 4 13 1 9 13 1 9 1 10 12 9 1 10 9 1 10 11 2 1 10 10 9 7 1 10 9 0 2
17 10 9 15 13 10 9 7 10 9 13 10 9 1 10 10 9 2
26 1 10 9 10 9 7 10 9 3 4 13 15 1 10 9 13 3 1 10 9 1 10 9 1 9 2
3 9 12 2
40 10 9 13 1 9 10 9 1 10 9 0 15 13 1 9 0 2 7 13 9 7 9 0 2 7 13 9 1 10 9 7 9 1 10 9 7 9 1 9 2
3 9 12 2
16 10 9 13 10 9 10 9 7 10 9 0 13 1 10 9 2
24 10 9 0 1 10 9 3 4 4 13 16 3 1 9 7 1 9 3 0 3 1 12 9 2
18 10 0 9 15 13 0 7 0 9 4 13 10 9 1 13 15 9 2
3 9 12 2
11 10 11 4 13 9 1 9 1 0 9 2
22 1 10 9 13 1 10 10 9 10 9 13 1 9 1 13 10 9 1 10 0 9 2
25 10 9 1 9 13 1 10 9 7 1 10 9 1 10 0 9 7 10 0 9 1 10 9 0 2
2 9 0
5 10 9 1 10 9
3 9 12 2
18 10 9 1 10 9 4 13 1 10 9 1 9 0 1 10 10 9 2
25 1 10 9 13 12 9 1 10 9 13 1 10 9 0 1 9 16 4 13 10 9 1 10 9 2
9 10 11 1 11 13 10 0 9 2
22 10 9 1 10 9 1 10 9 13 9 1 9 0 1 9 1 12 9 1 10 9 2
10 1 10 0 9 13 0 10 9 0 2
3 9 12 2
25 4 4 13 9 1 10 9 10 9 15 4 13 12 9 1 9 7 13 1 10 9 0 7 0 2
14 10 9 1 9 1 10 9 13 0 1 10 0 9 2
13 10 9 7 10 9 1 10 9 4 13 1 9 2
3 9 12 2
11 10 9 1 10 9 4 13 1 12 9 2
36 12 9 3 16 13 10 9 2 10 9 1 10 9 1 10 9 13 1 9 0 10 9 7 10 9 0 2 1 13 10 0 9 1 10 9 2
32 16 10 9 4 13 2 7 13 15 1 12 9 1 10 10 9 2 10 9 13 9 1 12 9 1 10 9 1 10 9 0 2
13 1 10 9 4 13 10 9 1 10 9 1 9 2
3 9 12 2
28 10 9 1 10 9 1 10 9 2 1 10 9 15 15 3 4 13 15 2 4 13 1 10 9 1 10 9 2
61 1 9 1 9 0 7 1 9 7 1 9 1 10 9 1 10 9 2 10 9 1 10 9 1 10 9 13 10 9 1 10 0 9 1 10 9 1 12 9 2 1 10 0 9 13 16 10 9 4 13 7 13 15 1 12 9 1 10 10 9 2
3 9 12 2
17 10 9 1 10 9 13 10 9 1 10 9 7 13 10 9 0 2
7 4 13 9 1 10 9 2
14 13 10 9 1 10 0 9 7 15 13 10 0 9 2
17 13 10 9 1 10 9 1 10 9 1 9 1 9 1 10 9 2
15 13 10 9 7 13 10 9 13 9 1 9 7 10 9 2
12 13 10 9 0 1 10 9 13 1 10 9 2
16 13 2 1 10 9 13 1 10 9 2 10 9 1 10 9 2
23 13 7 13 10 9 0 2 13 10 9 0 2 0 2 16 13 2 10 9 1 10 9 2
29 13 10 9 1 10 9 0 2 13 10 9 0 1 9 13 1 10 9 2 13 10 9 1 9 13 1 10 9 2
8 13 10 9 0 1 10 9 2
8 4 13 9 7 13 10 9 2
7 13 10 9 1 10 9 2
3 9 12 2
22 10 9 1 10 9 4 2 13 10 10 9 2 13 10 9 7 3 15 0 1 15 2
33 3 4 13 10 9 1 10 0 12 9 1 10 10 9 2 3 16 15 13 1 15 7 1 9 1 10 0 12 9 1 10 9 2
3 9 12 2
25 10 9 1 10 9 1 10 9 13 0 16 3 4 13 1 10 9 13 2 15 15 13 10 9 2
3 9 12 2
32 10 9 1 10 9 3 13 0 1 10 9 13 1 10 9 1 10 10 9 2 1 16 1 0 9 7 1 9 1 10 9 2
24 1 10 9 4 13 1 9 1 9 1 10 9 1 9 0 2 1 9 0 1 10 10 9 2
3 9 12 2
2 9 0
2 10 9
2 9 0
5 10 9 1 10 9
3 9 12 2
27 10 9 1 10 9 4 13 1 10 9 1 10 9 7 1 10 9 2 15 13 3 10 9 1 10 9 2
3 9 12 2
3 9 12 2
11 10 9 4 13 10 9 1 10 12 9 2
16 10 11 13 7 13 10 9 1 9 13 7 13 1 9 0 2
20 1 12 9 1 10 10 9 10 9 15 13 1 10 9 1 13 15 10 9 2
22 10 9 0 1 15 7 1 10 10 9 1 10 9 1 10 9 3 13 9 1 9 2
33 10 9 1 9 4 4 13 1 3 10 15 1 10 9 1 10 9 7 3 4 4 13 1 9 3 1 12 9 1 10 10 9 2
3 9 12 2
20 10 9 1 10 9 1 10 9 13 10 9 0 1 10 9 7 15 13 0 2
18 13 10 9 1 9 0 7 0 2 13 7 13 10 9 1 10 9 2
25 10 9 13 0 3 1 10 9 1 10 9 1 10 9 2 7 3 1 10 9 1 10 10 9 2
3 9 12 2
63 10 9 1 10 9 1 10 9 7 10 9 2 3 16 13 1 10 9 2 4 13 2 1 10 9 13 1 10 9 1 10 10 9 2 1 10 9 0 2 0 9 1 10 9 1 10 9 7 1 10 9 1 10 9 2 1 10 9 13 1 9 0 2
2 9 0
3 10 0 9
3 9 12 2
25 10 0 9 4 13 1 9 1 9 2 1 9 16 4 13 10 0 9 7 10 9 1 10 9 2
20 1 10 9 1 10 0 9 15 13 1 9 2 1 10 9 13 1 10 9 2
3 9 12 2
12 10 0 9 13 1 10 9 0 1 10 9 2
16 16 13 9 1 10 9 2 3 4 13 9 16 3 1 9 2
44 15 4 1 9 13 9 1 10 9 1 13 15 1 10 9 0 1 10 9 2 10 9 1 9 1 9 0 2 10 9 7 9 1 9 2 10 9 0 7 0 1 10 9 2
2 9 0
3 10 9 0
3 9 12 2
44 10 9 0 1 10 9 7 1 10 9 4 13 2 1 10 9 13 1 10 9 2 1 9 7 1 9 1 10 9 0 2 1 9 15 13 9 1 10 10 9 0 7 0 2
26 13 9 1 9 1 10 9 7 1 10 9 1 10 9 7 1 10 9 15 15 4 13 1 10 9 2
28 13 10 9 0 7 4 13 1 10 9 1 10 9 0 7 0 1 10 9 7 1 10 9 13 1 10 9 2
3 9 12 2
21 10 9 1 9 13 9 1 9 0 2 0 7 1 9 1 10 9 1 10 9 2
32 10 9 1 10 9 13 10 9 0 1 9 1 10 9 1 10 9 2 7 3 15 0 1 10 9 1 10 9 1 10 9 2
33 13 2 1 10 9 7 1 10 9 13 1 10 9 2 1 10 9 1 10 9 0 1 10 9 1 15 10 9 13 1 9 0 2
13 13 3 1 10 9 1 10 9 1 10 9 13 2
20 10 9 13 10 9 1 10 12 9 7 1 10 10 9 1 9 1 10 9 2
2 9 0
2 10 9
2 9 0
2 9 0
3 9 12 2
9 10 9 13 0 3 1 10 9 2
3 9 12 2
19 10 9 0 4 13 1 9 0 13 7 13 1 10 9 1 10 9 0 2
10 3 4 4 13 9 0 7 9 0 2
27 4 3 13 15 1 10 9 0 0 9 0 1 10 9 2 3 1 10 9 1 9 0 0 1 10 9 2
22 10 9 13 10 9 7 10 9 1 10 9 0 1 10 9 1 10 9 1 10 9 2
3 9 12 2
22 10 9 1 10 9 13 9 1 10 9 1 9 0 7 1 10 15 13 1 10 9 2
15 10 9 0 1 9 1 9 13 10 9 13 1 10 9 2
19 1 9 1 9 13 9 3 1 10 9 0 13 1 13 1 10 9 0 2
3 9 12 2
13 10 9 13 10 9 0 7 0 1 10 0 9 2
15 10 9 0 1 10 9 4 13 1 10 9 1 10 9 2
18 15 13 9 1 9 10 0 9 7 10 9 0 1 10 9 1 9 2
47 10 0 9 4 13 1 12 9 1 10 10 9 0 1 10 13 1 10 0 9 2 7 1 10 15 1 10 9 1 9 0 1 9 0 1 9 1 9 0 7 9 1 12 9 1 9 2
14 10 9 13 10 0 9 1 10 9 13 1 10 9 2
17 10 9 0 1 10 9 13 1 9 12 9 7 3 13 3 0 2
27 3 4 2 16 13 1 9 2 4 13 1 10 9 0 2 7 13 9 1 10 9 7 1 10 9 0 2
3 9 12 2
39 13 1 10 9 0 1 10 9 2 1 10 9 1 10 9 0 2 10 9 2 10 9 7 10 9 2 10 9 7 10 9 0 1 10 9 1 10 9 2
3 9 12 2
10 10 9 1 10 9 13 9 1 9 2
26 10 9 1 10 9 0 4 13 10 9 2 3 0 2 1 9 0 1 10 10 9 13 1 9 0 2
51 1 9 1 10 9 0 1 10 9 4 4 13 1 10 9 1 9 1 9 2 1 9 0 2 9 0 1 9 1 9 0 7 9 15 13 12 9 1 9 7 4 13 1 10 9 0 1 10 9 0 2
3 9 12 2
52 3 4 4 13 7 13 1 10 9 7 13 1 0 9 7 9 16 3 1 9 1 9 1 10 9 0 1 10 9 2 13 7 1 10 9 7 1 10 9 1 9 13 1 10 9 0 7 1 10 10 9 2
13 10 9 1 10 9 13 9 1 13 10 9 0 2
12 10 9 15 13 1 15 3 1 9 1 9 2
20 10 0 9 13 1 10 9 13 1 10 10 9 1 10 9 1 10 9 0 2
3 9 12 2
15 10 9 1 10 9 0 7 1 10 9 4 13 1 9 2
34 10 9 13 10 9 1 10 9 1 10 9 0 2 1 10 0 9 3 1 15 2 7 1 10 9 15 13 1 10 9 1 10 9 2
3 9 12 2
10 10 9 0 13 3 1 10 9 0 2
3 9 12 2
31 0 10 9 1 10 9 0 1 10 9 2 13 1 10 9 1 10 9 10 9 7 10 9 1 10 9 0 1 10 9 2
2 9 0
4 9 1 10 9
3 9 12 2
13 10 9 15 13 1 10 0 9 13 1 10 9 2
23 10 9 15 13 1 10 9 1 10 9 2 1 9 1 9 2 3 1 9 0 7 0 2
41 1 10 9 0 2 10 9 13 16 10 9 13 1 10 9 4 2 1 10 3 0 9 0 2 13 3 1 10 9 7 1 10 9 1 10 9 13 1 10 9 2
15 13 1 10 9 7 1 10 9 0 1 13 10 10 9 2
56 13 10 9 2 3 1 10 9 2 1 13 7 1 13 13 10 9 15 13 9 1 10 9 2 1 13 10 9 7 10 9 1 9 1 10 9 1 10 0 9 1 10 9 7 10 9 1 10 0 9 1 9 1 10 9 2
18 4 13 1 10 9 16 3 13 7 3 13 10 9 13 1 10 9 2
18 10 9 0 4 13 1 10 9 1 10 9 1 10 9 1 10 9 2
37 10 9 13 10 9 1 15 10 9 1 10 9 3 13 9 1 9 1 9 1 10 9 7 1 13 9 1 9 0 7 1 9 1 13 9 0 2
8 10 10 9 0 4 4 13 2
32 1 10 9 7 1 10 9 1 10 9 0 2 13 1 10 9 0 0 7 0 2 4 3 13 9 1 9 1 9 1 9 2
19 15 4 13 1 10 9 3 1 10 9 1 10 9 0 1 9 1 9 2
30 1 10 9 1 10 9 1 9 7 1 10 9 1 10 9 10 9 1 9 4 13 1 10 0 9 0 1 10 9 2
3 9 12 2
12 10 0 9 13 10 9 1 13 10 9 0 2
3 9 12 2
31 1 10 9 1 10 0 9 4 3 13 10 9 0 1 10 9 7 1 10 9 0 3 1 10 9 1 9 0 7 0 2
21 10 9 0 3 4 4 13 7 13 1 0 9 1 9 7 1 10 9 1 9 2
28 10 9 13 10 9 1 9 4 13 10 9 1 10 0 9 1 10 9 7 1 10 9 13 1 10 9 0 2
2 9 0
8 10 9 2 10 9 2 10 9
3 9 12 2
25 10 9 4 13 1 10 9 2 1 10 9 2 1 10 9 0 2 1 10 9 7 1 10 9 2
30 10 9 2 10 9 2 10 9 0 7 10 9 13 9 0 1 10 9 2 9 7 9 1 10 9 13 1 10 9 2
8 11 13 10 9 1 10 9 2
10 10 9 1 10 9 13 10 10 9 2
3 9 12 2
3 2 13 2
3 9 12 2
47 10 11 2 11 11 2 10 11 2 10 11 2 10 11 2 11 11 5 11 7 10 11 1 11 5 11 1 11 13 1 9 7 9 0 1 9 2 1 10 0 9 0 13 1 9 0 2
20 10 9 11 2 11 11 5 11 4 13 1 10 9 0 1 11 7 1 11 2
93 0 9 7 9 0 1 9 2 13 10 9 1 15 1 10 0 9 1 10 9 12 7 10 9 13 1 10 0 9 1 10 0 9 1 10 9 8 2 2 3 1 10 9 1 10 9 1 9 2 8 2 7 8 2 2 4 4 13 1 0 9 2 1 9 1 10 9 2 1 9 1 10 9 0 2 13 10 9 0 2 1 10 9 1 10 9 1 15 1 10 9 12 2
27 10 9 4 13 1 10 9 1 9 0 1 10 9 2 1 10 9 1 9 1 10 9 7 10 9 0 2
3 9 12 2
34 10 9 0 4 13 1 10 9 7 1 10 9 1 10 9 1 10 9 2 7 1 10 9 13 1 10 9 0 7 1 10 9 0 2
310 10 9 13 9 0 1 10 0 9 2 8 2 9 0 7 9 0 1 10 9 2 9 1 10 9 1 10 9 0 2 9 1 9 7 9 0 1 10 9 1 9 3 13 1 10 9 0 2 8 2 9 2 8 2 9 1 10 9 7 10 9 0 2 8 2 9 7 11 0 2 9 1 10 9 2 9 2 9 7 9 2 8 2 9 2 9 1 10 9 7 9 0 2 9 1 10 9 2 9 0 2 9 0 7 0 1 10 9 2 9 1 10 9 0 2 8 2 9 1 10 9 7 0 9 0 2 9 0 2 9 1 10 9 0 2 8 2 9 7 9 0 1 10 9 7 1 10 9 0 0 2 8 2 9 0 7 9 2 1 9 1 10 9 0 0 2 8 2 9 2 9 0 7 9 2 8 2 9 7 9 0 2 9 0 7 0 2 13 0 2 8 2 9 1 10 9 0 1 10 9 13 10 9 0 7 0 15 4 4 13 1 10 10 9 0 2 8 2 9 0 1 10 9 2 8 2 9 0 2 8 2 9 0 2 9 1 9 7 9 0 1 11 2 9 7 11 0 2 8 2 9 2 9 1 10 9 0 7 9 0 2 8 2 9 2 9 7 9 1 10 9 2 9 0 0 7 0 1 10 9 1 10 9 0 2 0 7 0 2 9 1 10 9 2 8 2 9 1 10 9 2 1 10 9 7 1 10 9 0 2
176 13 9 1 9 13 15 0 1 2 9 0 7 1 10 9 0 1 10 9 2 9 1 10 9 2 9 7 9 1 10 9 2 9 2 0 10 9 1 10 9 0 7 1 9 1 10 9 7 1 10 9 0 2 9 2 9 0 7 0 7 9 1 10 9 1 10 9 0 2 9 1 10 9 2 9 2 9 0 2 9 0 2 9 1 10 9 2 9 7 9 0 2 0 9 1 9 7 1 9 2 9 1 10 9 2 9 2 9 7 9 0 1 10 9 2 9 0 7 0 2 9 1 10 9 0 7 9 1 10 9 0 7 1 10 9 0 2 9 1 10 9 0 7 0 7 9 7 9 1 9 0 2 9 1 9 2 9 0 2 9 1 9 1 9 0 2 9 1 9 0 7 0 1 9 0 2
32 1 10 9 1 9 0 13 1 10 9 10 9 0 2 3 16 1 10 9 1 10 9 0 2 13 1 10 9 1 10 9 2
22 13 1 10 9 10 9 0 1 9 1 10 9 3 3 13 1 10 9 1 10 9 2
84 10 9 7 10 9 0 1 11 7 1 11 2 1 10 9 1 10 9 2 13 1 10 9 0 1 10 9 1 10 9 0 0 7 13 1 10 9 7 1 10 9 1 10 9 0 7 1 10 9 1 10 9 0 2 1 10 9 1 10 9 1 9 13 1 9 1 10 9 2 15 13 10 9 1 9 1 10 9 0 1 9 1 9 2
20 10 9 0 13 1 10 9 1 10 9 1 9 0 2 0 9 1 10 9 2
12 10 9 0 13 1 10 9 1 10 0 9 2
30 10 9 2 10 9 7 10 9 0 13 9 0 1 9 1 10 9 1 10 9 7 1 10 9 1 10 9 15 13 2
41 10 9 0 13 10 9 15 13 10 0 9 1 10 9 7 1 10 9 1 10 9 0 2 0 7 0 7 13 10 9 1 9 1 9 7 9 1 10 9 0 2
28 10 9 0 13 10 9 1 10 9 1 0 9 1 10 0 9 1 10 10 9 2 3 1 9 1 9 0 2
37 1 10 9 1 10 9 10 9 4 13 9 1 9 7 9 1 9 0 0 1 0 9 2 1 10 9 7 1 10 9 13 1 9 1 10 9 2
3 9 12 2
43 10 9 0 4 13 1 10 9 3 16 2 1 13 15 10 9 0 2 4 13 1 9 2 9 0 2 9 7 9 2 1 10 9 1 10 9 1 9 2 9 7 9 2
30 10 9 2 10 9 7 10 9 0 13 0 1 9 0 10 7 1 15 13 1 9 0 7 0 2 1 10 0 9 2
52 10 9 0 13 9 1 9 1 9 7 9 1 10 9 1 15 1 10 9 8 2 7 8 2 1 10 0 9 1 10 9 12 2 7 13 3 9 1 9 7 9 1 10 9 1 10 9 1 10 9 0 2
40 9 2 9 2 11 0 2 9 7 11 13 10 0 9 1 10 9 2 0 7 0 2 1 10 9 1 9 1 9 0 2 1 10 9 1 10 9 1 9 2
3 9 12 2
21 10 9 2 10 9 2 10 9 0 7 10 9 13 9 0 1 9 7 1 9 2
16 10 9 2 10 9 2 10 9 0 7 10 9 13 9 0 2
29 13 7 13 9 7 9 10 2 1 9 1 10 9 7 1 10 9 1 9 1 10 9 0 7 1 10 9 0 2
15 13 1 9 1 10 9 1 9 0 0 1 10 10 9 2
25 10 9 1 10 9 13 10 9 0 2 1 9 1 9 2 1 10 9 1 0 9 0 1 9 2
38 10 9 13 1 10 9 1 15 1 10 9 0 13 1 10 9 2 1 10 9 2 1 10 9 0 7 1 10 9 1 13 3 10 9 0 15 13 2
70 1 13 10 9 0 2 10 9 7 10 9 0 2 1 13 10 9 0 7 0 2 1 13 10 0 9 1 10 9 1 10 9 2 7 1 13 1 9 0 1 10 0 9 1 10 10 9 2 10 9 13 9 0 7 13 9 0 1 9 1 10 9 2 9 2 9 0 7 9 2
30 10 9 2 10 9 2 10 9 0 7 10 9 13 10 10 9 2 13 1 10 9 0 13 1 10 9 1 10 9 2
12 4 13 1 10 9 3 1 13 9 1 9 2
15 4 13 10 9 1 10 9 1 10 9 1 10 0 13 2
3 9 12 2
56 10 9 3 4 13 9 1 9 7 9 7 9 1 10 9 2 7 13 9 15 13 1 10 9 10 0 9 1 10 9 7 1 10 9 1 10 9 2 7 13 10 9 1 10 9 1 10 9 1 10 9 1 10 9 0 2
95 10 9 4 13 15 1 9 1 10 9 2 1 10 9 0 2 1 10 9 7 1 10 9 1 10 9 1 0 9 1 9 7 9 0 7 1 10 9 0 7 1 9 0 1 10 9 7 10 9 0 2 7 16 15 13 10 9 1 10 9 0 7 1 10 9 0 7 1 9 10 9 1 10 9 0 1 10 9 13 10 9 0 7 0 2 13 1 10 9 0 1 10 9 0 2
30 10 9 13 10 9 0 1 13 16 10 9 0 4 13 1 10 9 1 10 9 1 9 7 1 10 9 1 0 9 2
3 9 12 2
17 13 9 1 10 9 2 10 9 0 2 10 9 7 10 10 9 2
25 10 9 0 13 10 9 0 13 1 10 9 7 10 0 9 13 15 1 10 9 7 1 10 9 2
9 4 13 9 1 9 1 10 9 2
11 10 9 0 13 10 9 0 1 10 9 2
9 10 9 1 10 9 13 10 9 2
11 13 10 9 1 10 9 7 15 13 0 2
9 13 10 9 7 13 10 9 0 2
24 13 10 9 0 13 1 10 9 1 10 9 2 13 15 1 10 9 1 10 9 1 10 9 2
3 9 12 2
60 10 9 1 9 7 10 9 1 9 7 1 9 1 10 9 7 1 10 0 9 1 10 9 0 7 1 10 9 0 4 13 1 9 1 10 9 1 10 9 1 10 9 0 13 1 9 1 10 9 2 15 13 3 10 9 1 10 9 0 2
38 15 4 13 3 1 10 9 7 1 10 9 0 7 1 15 1 10 9 1 10 9 2 1 10 0 9 7 1 0 9 0 2 7 1 10 9 0 2
15 10 9 13 1 10 10 9 10 9 7 10 9 1 9 2
26 10 9 0 3 4 4 13 1 13 1 10 9 13 7 1 10 9 13 1 10 9 1 10 10 9 2
23 10 9 1 10 9 0 2 3 16 10 9 0 13 3 2 4 13 1 9 0 7 0 2
3 9 12 2
28 10 9 13 10 9 15 2 1 9 1 10 9 2 15 13 10 9 1 9 7 10 9 0 1 9 7 9 2
34 10 9 13 10 9 1 10 9 1 9 7 1 10 9 1 9 7 9 0 1 10 9 7 10 9 1 10 9 7 1 10 9 0 2
34 10 9 4 13 7 13 1 10 9 0 1 9 13 1 9 0 1 10 10 9 2 1 12 9 0 13 1 9 3 0 1 12 9 2
20 1 10 9 3 4 13 10 9 1 10 9 1 9 1 10 9 1 10 9 2
36 10 9 4 13 1 9 0 16 1 12 9 1 10 10 9 15 13 9 10 0 1 10 9 1 10 9 7 10 15 1 10 9 10 9 0 2
20 10 9 13 1 9 3 4 13 16 3 4 13 1 10 9 1 10 9 0 2
26 1 10 9 2 10 9 13 10 9 1 10 9 0 2 1 9 1 9 1 10 9 7 10 9 0 2
3 9 12 2
3 2 13 2
3 9 12 2
23 1 10 9 4 13 9 1 9 0 1 0 9 2 1 10 9 13 1 9 1 10 9 2
14 4 13 15 9 1 9 0 1 10 9 1 10 9 2
3 9 12 2
40 1 9 13 1 10 9 1 10 9 4 13 10 9 1 10 9 0 7 10 9 1 10 9 1 10 9 15 4 13 9 0 1 10 9 7 0 9 1 9 2
15 10 9 7 10 9 4 3 4 13 1 9 1 9 0 2
28 10 9 4 13 13 10 9 1 9 7 9 13 2 1 10 9 0 2 1 10 9 13 1 9 1 10 9 2
41 10 9 0 4 13 10 9 1 10 9 1 10 9 1 10 9 1 9 0 2 13 1 3 10 15 1 10 10 9 7 13 1 9 0 1 9 0 1 10 9 2
16 10 9 3 4 4 13 1 9 3 1 12 9 1 10 9 2
53 10 9 1 10 9 1 9 1 10 9 1 10 9 1 10 9 13 1 9 0 7 0 2 7 10 9 2 10 9 0 2 10 9 7 10 9 0 1 10 15 13 10 9 1 10 9 7 10 9 1 10 9 2
20 1 10 9 10 0 9 13 1 10 9 0 1 10 9 1 10 9 10 9 2
3 9 12 2
36 10 9 2 16 13 16 10 9 0 13 10 9 1 10 9 2 4 13 10 9 1 9 0 3 1 10 9 0 1 12 9 1 10 10 9 2
3 9 12 2
3 2 13 2
3 9 12 2
3 2 13 2
3 9 12 2
3 2 13 2
3 9 12 2
56 4 13 10 0 9 2 11 2 11 1 11 2 11 2 11 2 11 11 2 11 2 11 2 11 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2
3 9 12 2
65 15 4 2 1 9 0 2 13 10 9 0 2 13 10 9 1 9 13 7 10 9 1 0 9 1 10 9 1 10 9 1 9 2 16 15 13 9 10 9 0 15 13 3 10 15 1 10 9 0 2 7 10 9 4 13 1 9 1 10 9 1 10 9 0 2
66 15 4 2 1 10 9 1 10 9 1 10 9 1 10 9 7 1 10 9 0 7 1 10 9 7 1 10 9 0 13 1 9 7 1 9 1 10 9 2 13 10 9 0 2 13 16 9 7 9 2 15 15 13 9 2 4 13 1 10 9 7 13 1 10 15 2
3 9 12 2
37 10 9 1 10 9 0 7 10 9 1 0 9 1 10 9 1 10 9 4 13 1 9 1 10 9 2 1 9 1 10 9 2 13 10 0 9 2
27 10 9 2 13 10 9 0 2 4 1 10 9 13 1 10 10 9 0 9 7 13 10 10 9 7 9 2
2 9 0
2 9 0
2 9 0
3 10 9 0
3 9 12 2
77 10 9 0 13 2 1 10 9 0 1 10 9 0 1 10 9 7 1 10 9 2 13 9 1 9 2 1 10 9 7 1 10 9 2 1 10 9 1 9 1 10 9 1 10 9 7 1 15 1 10 9 7 10 9 2 7 1 10 9 2 1 10 9 13 1 10 9 1 10 9 2 1 9 1 10 11 2
3 9 12 2
40 10 9 0 4 13 1 12 9 13 1 10 15 1 10 9 1 10 9 2 1 10 15 1 10 9 1 9 0 7 1 10 15 1 10 0 9 0 7 0 2
39 10 9 1 10 9 0 4 13 1 10 9 3 1 9 1 10 9 0 0 7 0 2 10 9 0 1 9 1 9 0 7 10 9 1 12 9 1 9 2
31 10 9 1 10 9 0 4 13 1 12 9 2 13 1 15 1 15 1 10 9 1 10 9 2 7 3 4 4 3 13 2
21 1 10 9 1 10 9 10 9 0 13 1 10 9 7 1 10 9 1 10 9 2
45 10 9 13 1 10 10 9 2 1 10 9 13 1 10 9 2 10 9 2 15 13 1 9 1 10 9 2 7 13 0 2 0 1 10 9 10 9 1 9 1 10 9 1 9 2
41 10 9 1 9 1 10 9 13 0 1 15 1 9 1 10 9 2 1 10 9 0 2 1 10 9 1 10 9 1 9 7 1 10 9 7 9 13 1 10 9 2
63 1 10 9 1 9 1 10 9 1 10 9 2 13 2 1 10 9 0 1 10 9 2 12 9 13 1 9 1 10 9 1 9 13 10 9 1 10 9 1 9 2 15 10 9 13 10 12 9 1 9 1 10 0 9 13 1 10 9 1 10 9 0 2
3 9 12 2
37 16 10 9 13 10 9 0 1 10 9 1 9 7 1 9 13 9 1 9 2 10 9 13 1 13 9 1 10 9 0 1 10 9 1 10 9 2
32 10 9 1 10 9 4 13 7 13 1 10 9 7 1 10 9 0 0 2 16 2 16 15 13 0 2 13 1 10 9 0 2
3 9 12 2
13 1 10 9 1 10 9 0 3 4 13 10 9 2
2 9 0
4 9 1 10 9
2 9 0
3 9 12 2
46 10 9 1 9 1 10 9 7 10 0 9 0 4 13 1 10 9 1 12 0 9 1 9 3 0 1 12 9 2 7 4 13 1 9 0 1 10 9 1 10 9 1 10 0 9 2
37 10 9 0 4 13 1 9 0 16 2 1 12 9 1 10 10 9 2 15 13 9 10 0 1 10 9 1 10 9 7 12 9 7 12 9 0 2
21 10 9 13 1 9 3 4 13 2 16 3 4 13 1 10 9 1 10 9 0 2
31 3 15 13 9 1 9 16 10 9 4 4 13 1 10 0 9 1 15 1 10 9 1 9 1 12 9 1 10 10 9 2
3 9 12 2
11 10 9 0 3 4 13 9 1 9 0 2
1 0
28 1 10 9 1 9 1 10 9 10 9 0 1 10 9 13 10 9 1 9 1 10 9 7 15 13 10 9 2
1 0
33 16 1 10 9 1 10 9 1 10 9 1 10 9 3 4 13 10 10 9 0 2 13 1 10 9 3 10 9 1 10 12 9 2
1 0
128 1 10 0 9 1 10 11 1 10 9 4 13 9 2 1 9 1 10 9 1 10 9 2 10 9 1 10 9 0 15 13 10 9 1 9 1 13 9 7 15 2 2 4 13 9 1 10 9 1 10 9 7 1 9 0 2 2 4 13 9 1 10 13 11 2 2 4 13 3 12 9 2 0 15 1 10 9 0 2 2 4 4 13 13 1 10 9 1 10 11 1 10 9 1 10 12 9 12 2 2 4 13 10 9 1 10 9 3 0 1 12 9 1 9 1 9 1 10 9 0 0 1 10 9 1 10 9 2
29 4 13 3 9 2 1 9 1 10 9 1 10 9 2 10 9 1 10 13 9 15 4 13 9 1 10 9 0 2
20 1 10 9 1 4 13 9 15 4 13 3 1 10 9 1 10 9 1 9 2
19 10 9 1 10 9 1 10 9 0 13 9 1 10 9 1 9 1 9 2
1 0
33 1 10 0 9 1 10 9 10 11 4 13 1 9 1 15 0 2 1 10 9 1 10 9 15 15 13 1 9 1 10 10 9 2
1 0
38 10 9 1 10 9 12 1 10 9 2 1 15 13 10 9 0 15 13 9 1 10 9 7 9 1 9 2 13 9 1 10 9 1 9 1 10 9 2
1 0
46 1 12 9 1 10 9 1 9 1 10 9 15 13 1 10 9 1 10 9 0 1 9 3 13 2 1 10 9 1 10 9 1 9 2 1 10 9 1 10 9 7 1 10 9 0 2
26 1 10 9 1 10 0 9 15 13 1 9 1 10 9 1 10 9 0 0 1 9 1 10 9 12 2
1 0
30 3 1 16 3 4 13 10 0 9 1 10 9 0 1 9 1 10 9 2 13 1 13 15 10 9 1 10 9 13 2
1 0
29 10 9 1 10 9 0 7 1 10 9 0 1 10 9 0 4 13 1 10 9 1 10 9 1 9 1 10 9 2
23 9 1 10 9 13 1 10 9 1 10 0 9 10 9 1 10 9 0 13 1 10 9 2
46 3 1 16 3 4 13 1 10 9 7 1 10 9 1 10 9 0 1 10 9 0 13 1 10 9 7 1 10 9 10 9 15 13 3 7 10 15 1 15 10 9 13 15 10 9 2
33 9 1 10 9 13 10 9 1 10 9 1 9 7 9 1 10 9 2 3 1 10 9 0 2 15 4 13 0 1 10 0 9 2
33 1 10 9 1 10 10 9 10 9 4 2 1 16 1 9 1 9 2 13 10 10 9 1 15 1 10 9 7 1 10 9 0 2
1 0
36 10 9 2 1 12 9 1 10 9 1 9 1 10 9 2 13 10 10 9 1 10 9 1 10 9 0 7 1 10 9 0 13 1 10 9 2
1 0
1 0
63 3 1 12 9 1 10 9 1 9 1 10 9 15 4 2 1 9 0 2 13 0 9 2 1 9 1 10 9 1 15 1 10 9 12 2 3 1 10 9 1 10 9 13 1 10 0 9 1 10 9 12 2 0 13 3 10 9 1 13 10 9 0 2
1 0
15 4 13 10 9 2 1 10 9 2 1 10 13 9 0 2
1 0
34 10 9 2 13 1 10 9 0 2 1 10 0 9 1 9 11 2 1 10 10 9 7 1 10 10 9 0 2 4 13 1 10 9 2
25 10 9 7 10 9 1 9 0 1 10 9 0 15 15 4 13 1 10 12 9 12 2 13 0 2
1 0
7 10 9 0 3 4 13 2
18 10 9 1 15 13 3 1 10 12 9 12 13 1 9 1 10 9 2
18 10 9 0 4 13 1 9 0 7 13 1 10 9 13 1 10 9 2
10 10 9 13 10 9 1 10 9 0 2
1 0
1 0
37 1 10 9 1 10 9 1 9 1 10 9 15 13 1 10 9 7 1 10 9 1 15 1 10 0 9 0 15 3 4 13 3 3 7 3 13 2
1 0
44 10 9 0 4 13 1 10 10 9 1 13 2 1 10 12 9 12 2 1 10 9 1 10 9 1 10 9 1 10 9 2 1 10 9 0 0 7 1 10 9 1 10 9 2
10 1 10 9 10 9 0 13 1 9 2
23 15 0 13 1 10 9 10 9 1 9 2 1 15 13 2 1 0 9 7 9 1 9 2
14 10 9 4 13 1 10 9 9 1 9 1 9 13 2
36 10 9 0 2 1 10 9 1 15 1 10 0 9 1 10 0 9 2 4 13 1 10 10 9 1 9 0 1 10 9 7 1 3 12 9 2
1 0
35 10 0 9 4 13 1 10 9 0 1 10 9 1 12 9 1 10 10 9 1 9 1 10 9 0 2 7 13 1 9 10 0 9 12 2
36 10 9 1 10 9 4 13 1 10 9 0 1 10 9 1 10 9 1 13 15 0 2 1 10 10 9 12 2 16 10 9 4 13 15 9 2
28 10 9 2 13 1 10 9 1 10 9 2 4 13 1 10 9 0 1 10 9 7 1 10 9 1 10 9 2
8 9 1 11 2 9 12 9 12
3 11 11 11
21 13 2 10 9 1 10 9 0 11 11 10 9 1 10 9 1 10 9 11 11 11
5 13 2 10 9 11
79 9 12 5 12 5 11 1 10 9 0 7 1 10 9 1 10 12 9 12 0 1 10 9 1 10 9 1 10 9 1 9 1 10 9 0 1 10 9 15 13 9 7 13 9 1 10 9 12 5 12 5 11 1 10 9 7 1 10 9 12 5 12 5 11 7 12 5 12 5 11 1 10 9 0 7 1 10 9 2
68 10 9 0 7 10 9 1 10 11 11 2 13 10 9 15 13 10 9 0 2 1 9 10 9 12 2 13 10 9 1 10 9 2 13 10 9 1 10 9 0 7 0 0 2 12 2 2 13 1 10 9 1 15 1 10 9 12 1 10 9 2 12 2 2 13 15 13 2
62 2 12 2 10 9 13 1 10 9 7 10 9 0 13 1 10 9 9 1 9 1 10 9 0 1 10 9 15 13 9 4 13 9 1 10 9 7 13 10 9 1 10 9 7 4 3 13 10 9 0 1 10 9 7 1 10 9 1 10 9 0 2
22 10 9 1 10 9 0 13 10 0 9 1 13 10 9 1 10 9 7 10 9 0 2
27 2 12 2 1 10 9 15 13 9 13 0 10 9 0 1 10 9 1 9 0 7 1 9 1 10 9 2
11 15 13 3 10 0 9 0 1 0 9 2
31 1 10 0 9 1 10 9 1 9 0 1 10 9 0 15 4 13 9 3 0 1 9 0 16 10 10 9 0 13 0 2
48 1 10 9 1 10 9 0 2 4 4 13 10 0 9 1 10 9 0 0 1 10 9 2 1 9 13 10 0 9 1 9 0 0 7 13 10 9 1 10 9 16 10 9 3 13 9 0 2
25 2 12 2 10 9 0 1 10 9 13 10 9 0 1 10 9 0 1 10 9 0 1 10 9 2
42 1 9 0 13 1 10 9 1 10 9 0 1 10 9 13 3 10 10 9 1 9 2 15 13 0 7 0 9 1 10 9 2 10 9 7 10 9 1 10 10 9 2
50 2 12 2 10 9 1 10 9 0 2 15 1 10 10 9 0 13 10 9 3 0 1 10 9 2 4 13 10 9 0 1 10 9 1 10 9 1 9 1 10 9 1 9 1 9 9 1 10 9 2
46 10 9 1 9 13 15 15 13 10 0 9 1 10 9 1 9 0 1 9 7 15 13 16 15 13 1 10 0 12 2 12 9 2 1 9 1 10 9 0 15 15 13 1 10 9 2
29 10 0 9 1 10 9 1 9 2 16 13 1 10 9 1 10 9 0 1 10 9 0 2 11 2 2 13 0 2
39 10 9 0 13 15 1 10 9 1 10 0 9 1 9 1 10 9 2 13 1 9 9 12 5 12 5 11 1 10 9 0 7 1 10 9 2 12 2 2
33 10 9 0 13 15 1 10 9 3 0 2 1 10 9 1 10 9 2 1 13 10 9 1 10 9 7 13 10 9 1 10 9 2
15 4 3 4 13 9 7 9 0 1 10 9 1 10 9 2
52 2 12 2 13 0 13 1 10 9 0 1 10 9 15 13 9 2 16 4 13 16 13 1 10 9 16 15 13 10 9 13 1 10 9 1 9 1 10 9 7 13 3 16 15 13 10 0 9 1 10 9 2
50 2 12 2 13 13 10 9 0 1 10 9 1 10 9 0 1 10 9 0 1 10 9 15 13 9 1 10 9 1 13 10 0 9 1 10 9 15 13 1 10 9 7 1 13 15 10 9 0 0 2
17 10 9 0 4 13 10 9 1 10 9 0 7 1 10 9 0 2
49 2 12 2 10 9 1 10 9 0 4 4 13 13 9 1 10 9 7 1 10 9 1 10 0 9 0 1 9 1 9 0 2 13 2 16 0 2 10 9 0 1 10 0 9 0 1 10 9 2
45 2 12 2 10 0 9 4 13 1 13 10 0 9 1 9 13 10 9 0 0 1 10 9 15 13 9 2 10 15 15 13 1 0 1 10 9 1 10 9 7 10 0 9 0 2
21 10 9 0 13 3 10 0 9 1 10 9 0 2 0 7 0 1 10 9 13 2
37 10 9 1 10 9 0 1 10 9 13 1 13 10 9 1 10 9 0 2 15 15 13 10 9 0 1 10 0 9 0 7 3 1 10 9 0 2
105 2 12 2 10 9 9 15 13 0 13 9 0 1 9 1 9 0 1 9 1 9 1 10 9 2 7 13 0 9 0 1 0 9 0 13 1 10 9 1 10 9 1 9 1 10 9 0 1 10 9 9 13 1 10 9 1 10 9 1 9 0 2 4 13 15 1 10 9 1 10 9 13 1 10 9 12 2 9 12 2 12 7 12 2 1 10 9 2 15 13 10 9 0 1 10 9 7 10 9 1 9 1 10 15 2
53 2 12 2 1 13 10 9 0 13 1 10 9 1 10 9 2 4 13 0 13 10 9 1 9 1 10 9 7 1 10 9 0 1 10 9 15 13 9 7 13 15 9 1 10 9 1 10 9 0 1 10 9 2
56 2 12 2 10 9 13 1 10 9 0 1 10 9 0 0 1 10 9 2 15 13 10 0 9 1 10 0 9 0 1 9 1 9 1 9 2 13 0 1 13 10 9 0 1 10 9 1 10 9 1 10 0 9 1 9 2
37 13 1 9 2 1 10 9 1 10 9 2 10 9 0 15 10 9 13 1 10 0 9 1 10 10 9 4 13 3 1 10 9 7 1 10 9 2
28 13 0 9 1 13 16 10 9 4 13 1 10 9 1 10 9 3 13 9 1 10 9 0 2 0 7 0 2
47 2 12 2 16 13 0 10 9 0 1 10 9 0 2 10 9 1 10 9 1 9 9 1 10 9 1 10 9 0 4 4 13 10 9 0 0 1 9 1 10 9 1 10 9 1 9 2
41 2 12 2 4 13 0 7 0 13 0 9 0 1 10 9 0 1 10 9 7 9 0 1 15 0 1 10 9 1 13 16 10 10 9 0 4 13 1 10 9 2
72 13 10 0 9 1 13 1 10 9 1 10 9 13 1 10 9 1 10 9 1 11 13 1 10 9 9 1 10 11 11 1 10 9 0 2 7 13 0 10 9 0 13 1 10 0 9 2 13 13 9 1 10 9 15 13 10 0 9 1 9 1 10 9 1 9 1 9 9 1 0 9 2
47 10 9 4 13 3 1 13 10 9 0 1 10 9 7 13 10 0 9 1 10 9 0 1 9 1 10 9 7 10 9 0 13 1 10 9 0 1 10 9 0 1 11 1 10 9 12 2
48 2 12 2 16 13 13 1 9 10 9 7 10 9 3 0 0 1 10 9 2 13 10 9 0 2 10 9 1 10 9 1 10 9 0 4 4 13 1 10 9 1 9 0 2 0 7 0 2
18 10 9 0 1 9 1 10 9 4 13 10 0 9 1 10 9 0 2
13 10 9 0 4 4 13 7 13 3 1 10 9 2
14 10 9 1 9 0 13 10 0 9 1 10 9 0 2
20 10 9 4 13 1 9 10 9 1 10 9 1 9 0 7 1 9 1 9 2
33 10 9 1 9 0 13 10 9 1 10 9 2 13 1 13 10 9 1 9 1 10 9 7 13 10 9 1 0 9 1 10 13 2
37 2 12 2 13 13 10 9 1 9 0 1 10 9 1 9 1 10 9 16 15 13 1 13 10 9 1 9 3 0 7 3 0 1 1 9 13 2
24 9 0 4 13 15 0 16 10 9 1 9 3 15 13 1 10 0 9 7 1 10 9 0 2
59 2 12 2 10 9 2 13 10 9 0 1 10 9 0 1 9 1 10 9 2 4 13 0 9 1 9 1 10 9 0 7 0 1 10 9 1 9 1 10 9 7 13 10 9 0 7 0 1 10 9 0 7 1 10 9 1 10 9 2
38 2 12 2 1 10 9 1 10 9 1 9 0 7 1 0 9 1 9 13 1 9 1 10 9 1 9 2 4 4 13 10 9 3 1 10 0 9 2
38 9 0 2 9 0 2 9 2 9 13 7 13 2 9 1 10 9 0 2 9 7 9 2 9 9 5 9 1 10 9 1 10 9 1 9 2 9 2
63 2 12 2 1 9 1 9 1 10 9 1 9 1 9 1 10 9 1 10 9 1 10 0 9 2 10 9 12 1 10 9 1 10 9 1 10 9 0 1 9 1 9 1 10 9 1 10 9 1 9 2 13 7 13 10 9 2 4 13 1 9 0 2
33 2 12 2 10 0 9 4 3 13 10 9 1 10 9 1 9 0 1 9 1 10 0 7 0 9 2 11 2 7 1 10 9 2
28 10 9 4 4 13 1 10 0 9 1 9 1 10 9 1 10 10 9 7 1 10 9 1 9 1 10 15 2
28 10 9 0 1 10 9 1 9 13 0 1 13 10 9 0 1 10 9 15 13 9 13 7 13 10 9 0 2
74 2 12 2 1 10 9 1 10 9 1 9 7 1 10 9 1 9 2 10 9 4 13 10 9 1 10 9 9 7 10 0 9 0 1 10 9 1 9 2 1 10 9 2 13 11 7 9 2 10 9 2 10 9 2 10 9 2 10 9 2 10 9 1 10 9 1 10 9 7 10 9 1 9 2
61 2 12 2 1 9 1 9 1 10 9 1 9 2 10 9 4 3 13 1 10 0 9 10 13 9 0 1 9 1 9 2 13 1 9 10 9 0 2 15 10 9 9 4 13 1 13 0 13 1 13 10 0 9 0 1 9 1 10 9 9 2
85 2 12 2 13 13 9 1 10 9 7 1 10 9 1 13 1 10 9 1 9 0 1 15 1 10 9 12 5 12 5 11 1 10 9 2 1 10 12 9 12 2 13 10 9 0 1 10 10 9 1 10 9 1 9 1 10 9 7 10 9 1 10 9 7 10 9 1 10 9 11 1 9 2 1 13 1 10 9 1 9 0 2 12 2 2
35 2 12 2 10 9 13 1 10 9 4 13 15 9 1 10 9 13 1 10 9 1 10 0 9 1 10 9 1 13 10 9 1 10 9 2
19 10 9 4 13 15 10 3 0 1 9 0 1 9 7 1 0 9 0 2
28 4 4 13 10 9 1 9 1 10 9 1 10 9 0 1 10 9 1 9 7 1 10 9 1 9 1 9 2
35 10 9 7 10 9 1 10 9 1 10 9 13 1 10 9 1 9 0 1 10 9 13 15 1 10 9 0 1 9 0 1 10 0 9 2
53 2 12 2 10 9 0 13 1 9 10 9 0 7 0 2 13 1 10 9 0 2 15 13 10 0 9 1 9 7 9 1 9 0 1 13 10 9 1 10 9 1 15 13 10 10 9 1 10 9 1 9 0 2
33 2 12 2 13 9 1 10 9 1 13 10 3 9 2 10 9 9 4 13 16 13 0 10 9 0 1 10 0 9 1 10 9 2
33 2 12 2 1 15 13 10 9 7 10 9 1 10 0 7 0 9 1 9 1 9 0 2 4 13 0 13 1 9 9 1 9 2
22 2 12 2 13 1 10 9 1 10 9 1 10 9 0 13 1 9 13 1 9 0 2
58 10 9 13 10 9 1 10 9 1 10 9 0 1 10 11 11 2 10 9 1 15 4 13 10 9 1 9 1 10 0 9 13 1 10 9 1 9 13 1 10 9 1 10 0 9 2 3 16 4 4 13 0 9 1 13 10 9 2
33 2 12 2 15 1 10 9 0 1 10 9 13 4 13 1 10 13 10 9 1 13 10 9 1 9 13 1 9 1 10 0 9 2
19 10 9 4 13 1 9 0 1 10 9 1 10 9 1 9 7 1 9 2
41 1 10 9 1 9 0 1 9 0 2 10 9 13 4 13 3 1 13 10 9 1 10 9 1 10 9 0 1 10 10 9 1 10 9 1 10 9 1 9 0 2
17 10 9 4 13 3 10 9 1 10 10 9 7 10 9 1 9 2
17 10 9 13 3 4 13 10 9 1 13 9 3 1 10 9 0 2
26 2 12 2 1 10 9 13 1 10 0 9 2 13 0 13 15 1 10 0 9 0 2 1 11 12 2
61 2 12 2 10 0 9 13 0 1 10 9 1 10 9 1 10 0 9 13 1 10 9 1 10 9 2 1 10 12 9 12 2 0 1 10 0 9 1 9 1 9 0 7 9 2 12 2 2 7 1 10 9 1 13 9 1 10 9 0 13 2
57 10 9 1 10 9 1 10 12 9 12 1 10 9 1 10 9 1 11 2 12 2 13 1 10 9 1 13 16 10 9 1 10 0 9 4 4 13 1 9 3 3 13 1 9 2 1 9 1 13 7 13 10 3 0 10 9 2
290 2 12 2 10 0 9 13 0 1 10 13 9 0 2 1 10 9 12 5 12 5 11 1 10 9 2 1 10 12 9 12 2 13 10 9 1 10 9 1 9 7 1 0 9 1 10 9 0 2 1 10 9 7 9 0 0 1 10 9 2 12 2 2 10 9 2 11 2 9 12 5 12 1 10 9 0 7 1 10 9 2 1 10 12 9 12 2 0 1 10 9 0 2 13 2 1 9 1 10 9 1 9 0 2 12 2 2 10 9 2 11 2 9 12 5 12 1 10 9 0 7 1 10 9 2 1 10 12 9 12 2 13 10 9 0 1 9 0 1 10 9 0 1 10 9 1 10 9 1 9 2 12 2 2 10 9 12 5 12 5 11 1 10 9 0 7 1 10 9 2 1 10 12 9 12 2 1 10 9 1 9 0 7 0 2 11 2 2 12 2 2 10 9 12 5 12 5 11 1 10 9 0 7 1 10 9 2 1 10 12 9 12 2 1 10 9 1 10 9 1 10 9 0 1 10 9 0 7 0 2 12 2 2 7 10 9 12 5 12 5 11 1 10 9 2 1 10 12 9 12 2 13 10 9 1 10 9 0 2 0 7 0 1 10 9 9 0 1 10 9 1 9 1 9 1 10 9 7 1 9 1 10 9 7 9 0 2 12 2 2
30 10 9 1 10 0 9 7 10 9 0 13 4 13 1 13 10 0 9 7 1 13 9 0 1 13 13 1 10 9 2
147 2 12 2 10 9 12 5 12 5 11 1 10 9 2 1 10 12 9 12 2 13 10 9 1 9 1 10 0 9 1 9 0 13 1 9 0 7 0 2 12 2 2 10 9 12 5 12 5 11 1 10 9 0 7 1 10 9 2 1 10 12 9 12 2 1 10 9 1 9 0 1 9 2 9 7 10 9 1 9 0 2 12 2 2 7 10 9 12 5 12 5 11 1 10 9 0 7 1 10 9 2 1 10 12 9 12 2 1 10 9 1 9 0 1 10 9 1 9 0 2 12 2 2 15 3 13 9 1 9 1 10 9 1 10 9 1 9 0 2 4 4 13 1 10 0 9 2
31 2 12 2 10 9 12 5 12 5 11 13 10 9 1 9 1 10 9 1 9 1 10 10 9 0 1 10 9 1 9 2
35 16 10 9 9 7 10 9 4 13 16 0 9 3 4 13 10 9 13 2 10 9 12 5 12 5 11 4 4 13 1 13 9 3 0 2
167 2 12 2 10 9 1 10 9 12 5 12 5 11 1 10 9 2 1 10 12 9 12 2 13 10 9 1 10 9 1 9 13 1 10 9 1 9 7 10 9 1 9 0 1 10 9 3 0 0 7 3 13 2 7 10 9 1 10 9 1 10 9 7 1 9 0 1 9 0 1 10 0 9 3 0 2 12 2 2 4 4 13 1 10 9 1 10 9 12 5 12 5 11 2 1 10 9 12 5 12 5 11 1 10 9 2 1 10 12 9 12 2 13 10 9 1 10 9 1 10 9 9 1 9 1 9 1 9 2 12 2 2 7 1 10 9 12 5 12 5 11 1 10 9 0 7 1 10 9 2 1 10 12 9 12 2 1 10 9 0 1 10 9 2 12 2 2
12 10 9 12 5 12 5 11 4 3 4 13 2
33 9 1 10 9 1 10 9 0 7 1 10 9 1 10 9 7 9 1 10 9 11 0 1 10 9 1 10 9 1 10 9 0 2
52 9 1 9 1 10 9 15 13 7 13 10 9 1 10 9 1 10 12 9 12 2 15 13 10 9 1 9 1 9 1 9 2 9 7 9 1 10 9 1 10 9 1 10 9 0 2 9 2 11 2 2 2
80 11 2 10 9 0 0 1 10 9 2 1 10 9 7 1 10 9 1 10 9 1 10 9 1 10 9 0 2 4 4 13 1 10 9 9 12 5 12 5 11 1 10 9 2 1 10 12 9 12 2 7 4 13 1 13 7 13 10 9 13 1 10 9 9 7 13 1 9 13 1 10 9 1 10 9 1 10 9 0 2
34 0 9 13 10 9 1 9 2 9 2 9 2 9 7 9 2 2 10 9 7 10 9 1 9 2 7 10 9 0 2 0 7 0 2
27 10 9 12 1 10 9 11 13 16 10 9 1 9 13 9 10 0 9 12 7 15 13 10 12 9 12 2
26 10 9 12 1 10 0 9 13 1 10 9 1 10 9 10 9 1 9 0 0 1 12 9 1 11 2
31 10 9 12 2 9 12 2 1 10 9 11 13 16 10 9 13 1 10 9 0 7 1 10 9 2 1 10 12 9 12 2
28 2 10 9 1 9 0 1 1 10 9 1 10 9 1 10 9 2 10 9 7 10 9 1 10 9 2 7 2
19 2 10 9 1 10 9 1 13 7 13 10 9 2 13 1 10 9 0 2
16 10 9 1 9 1 10 9 11 4 4 13 10 12 9 12 2
39 10 0 9 13 9 1 10 9 7 9 1 10 9 1 9 2 13 9 1 10 9 1 10 9 7 4 13 1 10 9 1 9 7 9 1 10 9 0 2
27 1 10 9 1 10 9 12 2 10 9 9 13 13 16 13 1 9 15 4 13 1 12 9 1 10 9 2
40 10 9 13 0 1 10 9 0 10 9 1 10 9 2 0 1 1 10 9 0 1 10 9 0 7 3 0 1 9 1 10 12 9 1 9 9 0 1 9 2
31 1 10 0 9 15 13 10 0 9 1 10 9 1 9 13 2 15 4 13 1 10 9 13 0 13 10 9 13 1 9 2
35 10 9 1 9 4 3 13 1 9 1 9 10 9 1 9 2 13 9 0 7 13 0 9 1 9 7 9 13 3 16 4 13 1 9 2
20 10 9 12 8 7 12 8 13 10 9 1 10 9 1 9 7 9 1 9 2
31 10 9 3 0 13 10 9 1 10 0 9 1 9 7 0 7 0 7 13 10 0 9 1 9 13 1 9 0 7 0 2
26 10 9 4 13 10 9 0 0 1 10 9 1 10 9 1 10 9 13 3 1 10 12 2 12 2 2
69 10 9 4 3 13 1 10 12 10 9 1 9 2 12 2 2 15 13 10 9 0 1 10 9 1 9 2 7 15 4 4 13 1 10 9 9 1 10 9 2 12 2 2 13 1 10 12 2 1 15 10 9 1 10 9 1 9 1 9 0 4 13 7 2 1 9 2 13 2
25 1 10 12 2 3 2 10 9 1 11 4 4 13 1 10 9 1 10 9 1 9 2 12 2 2
25 1 9 1 10 9 0 2 10 9 4 13 12 9 2 12 2 1 10 9 1 10 0 9 9 2
10 10 9 1 9 15 15 13 13 0 2
38 1 10 9 1 13 10 0 9 1 10 9 1 10 9 0 2 10 0 9 7 10 0 9 1 9 2 4 4 13 9 0 0 1 10 10 9 9 2
14 1 10 11 7 11 13 0 9 9 7 9 1 9 2
36 4 4 3 13 0 9 1 10 9 0 1 10 9 13 1 10 9 9 2 1 10 11 2 1 10 9 2 7 10 9 2 1 10 9 2 2
49 10 9 11 13 10 9 1 9 1 10 9 1 10 9 0 1 10 9 1 10 9 1 10 9 7 1 10 9 1 10 9 1 9 1 9 0 2 9 1 10 9 1 9 7 1 10 13 9 2
33 10 9 0 13 0 1 13 10 9 13 1 10 9 1 10 9 1 10 9 1 10 9 7 13 15 9 1 13 1 10 9 0 2
21 10 9 7 10 9 0 13 3 0 1 10 9 7 13 3 0 13 10 9 11 2
48 3 1 10 9 12 1 10 9 11 2 10 9 1 10 9 11 4 4 13 1 10 9 0 1 10 9 0 1 10 9 0 2 11 2 2 15 4 13 10 0 9 1 9 10 12 9 12 2
35 10 9 4 13 10 9 0 1 12 1 10 9 1 10 9 11 13 3 1 10 9 12 2 1 9 1 10 0 9 9 7 1 10 9 2
32 13 15 1 10 9 15 4 13 9 7 9 7 1 10 9 1 10 13 2 10 9 4 13 1 10 0 9 0 2 12 2 2
17 2 10 9 4 13 1 13 10 9 1 10 9 0 1 10 9 2
37 15 13 3 10 0 9 2 1 9 1 10 9 2 1 10 9 7 1 10 9 13 2 1 9 1 10 0 9 0 7 1 10 3 0 9 0 2
34 2 1 15 13 10 9 1 10 9 1 9 7 10 9 5 10 9 2 4 13 1 10 0 9 13 1 10 10 9 2 9 7 9 2
12 2 10 9 1 10 9 4 4 13 3 3 2
44 15 4 13 3 10 0 9 1 9 1 0 9 2 16 10 9 1 10 9 1 10 9 0 2 9 0 2 7 1 10 9 1 9 7 15 1 10 9 0 4 13 3 0 2
18 2 10 9 13 4 4 13 0 7 0 1 10 9 0 1 10 9 2
21 2 1 15 13 10 9 2 10 9 4 13 3 0 10 9 2 13 15 9 0 2
9 10 9 4 13 10 0 9 0 2
8 1 12 9 13 10 0 9 2
49 2 10 9 4 13 1 9 1 10 10 9 9 7 4 13 10 9 2 1 0 9 2 1 10 9 15 4 13 3 1 10 9 7 3 4 13 9 1 10 0 9 2 7 1 10 0 9 9 2
11 2 13 0 13 10 9 1 10 9 0 2
20 10 9 4 13 1 10 9 1 9 7 1 10 9 0 2 13 9 1 9 2
11 10 9 13 3 10 0 9 9 2 9 2
55 2 4 13 10 9 1 10 9 5 10 9 0 5 0 2 9 5 11 2 11 7 11 2 1 13 9 1 9 0 7 13 3 10 9 1 10 0 9 2 9 1 9 2 9 2 9 2 1 10 9 1 10 9 0 2
51 2 1 9 1 10 9 1 10 9 1 10 9 1 10 9 1 0 9 1 9 2 3 4 13 0 13 1 10 9 1 3 3 13 0 0 9 1 10 9 1 10 9 0 7 10 9 1 10 9 11 2
53 2 1 13 10 9 1 10 9 1 10 9 2 1 10 15 3 1 9 1 10 9 1 10 9 1 0 9 1 9 2 10 9 13 10 9 1 10 9 0 1 13 3 1 10 9 1 9 1 10 0 9 11 2
27 10 9 1 10 9 4 13 3 0 2 1 9 3 1 10 9 16 10 9 4 4 13 1 10 9 12 2
50 10 0 9 1 10 9 11 4 4 3 13 3 1 10 9 12 7 10 9 13 1 10 12 4 13 1 3 0 1 10 12 5 1 10 9 0 2 10 9 4 4 13 1 10 9 1 10 9 2 2
21 3 10 9 4 13 7 10 9 4 4 3 13 7 1 10 12 7 1 10 12 2
17 1 9 1 10 9 1 10 12 2 3 10 9 0 4 3 13 2
32 1 10 9 5 9 2 10 9 0 1 10 9 1 10 9 12 2 12 13 0 1 10 12 5 1 10 9 1 9 0 0 2
17 10 0 9 1 10 9 1 10 9 11 4 13 1 10 9 12 2
14 1 10 0 12 9 1 10 9 4 4 13 12 9 2
19 1 10 12 4 13 0 12 9 2 13 1 10 9 9 7 1 10 9 2
36 1 10 12 9 0 2 12 13 1 10 9 1 10 9 0 1 10 9 9 2 16 10 13 12 4 13 1 9 1 10 9 5 1 10 11 2
20 10 0 9 1 10 9 13 13 1 9 2 9 2 9 7 9 1 9 0 2
26 1 13 3 16 10 9 1 9 4 13 3 0 9 7 4 4 3 13 1 10 9 1 10 9 11 2
29 1 9 1 10 9 13 0 16 10 9 1 10 9 1 9 13 2 3 1 10 9 1 10 9 1 10 9 11 2
27 1 10 9 1 10 0 9 4 4 13 3 10 9 0 2 15 15 13 13 1 9 3 0 1 10 12 2
20 10 9 1 10 9 11 1 9 1 10 9 1 9 4 13 1 10 9 12 2
11 1 10 0 9 4 13 9 3 12 9 2
44 1 10 0 9 10 9 13 1 10 0 9 9 1 10 9 1 9 2 1 9 1 10 9 13 1 10 9 1 3 0 9 0 1 10 9 3 0 1 10 9 1 10 9 2
40 1 10 9 2 10 9 1 9 2 9 12 7 12 2 13 16 2 3 1 10 9 12 2 10 12 5 1 10 9 4 13 3 1 9 1 10 9 1 9 2
54 1 13 1 10 12 15 13 3 10 0 9 1 10 9 0 2 7 1 10 12 2 12 15 13 10 9 1 10 9 1 9 1 10 9 0 2 9 0 1 10 9 0 2 9 0 0 2 9 0 7 9 0 2 2
12 3 10 9 13 0 1 10 9 1 10 9 2
15 4 13 1 10 9 10 9 1 10 0 9 1 9 0 2
29 1 10 9 1 10 9 15 4 13 1 13 9 1 10 9 7 10 9 1 9 4 13 16 10 9 4 4 13 2
26 1 10 9 1 9 13 16 10 9 13 1 12 9 2 16 15 13 10 9 1 9 1 10 9 9 2
21 4 4 13 10 0 9 1 10 9 2 1 10 15 15 1 10 9 1 10 9 2
22 15 4 4 13 1 9 1 9 0 3 1 0 2 7 15 4 13 1 13 10 9 2
34 10 9 13 3 0 1 15 1 10 9 1 10 9 2 1 10 11 15 13 1 9 1 10 12 5 1 10 9 0 1 10 9 13 2
19 1 10 12 3 10 0 9 9 4 13 1 13 9 0 1 10 9 11 2
68 10 9 1 9 13 3 2 9 12 2 16 10 9 1 10 9 0 1 10 9 11 4 13 10 10 9 0 1 10 9 1 10 9 2 9 1 9 2 9 0 2 0 7 0 2 2 13 1 9 10 9 1 9 1 10 15 13 1 0 9 10 9 1 10 9 1 9 2
39 1 10 9 1 10 9 11 4 13 10 9 1 10 11 2 1 10 9 2 1 11 7 2 1 10 9 2 3 1 11 2 11 7 1 10 9 0 0 2
30 1 9 1 10 9 1 10 9 1 10 9 1 9 1 10 9 9 2 4 4 3 13 10 9 1 10 0 9 0 2
18 10 9 1 10 9 11 4 1 10 9 13 1 10 9 1 10 11 2
69 15 1 15 4 4 3 13 1 10 9 0 7 1 10 9 9 1 10 9 1 13 9 1 9 0 13 1 10 9 1 10 9 2 3 1 10 9 1 10 9 13 1 11 2 1 10 10 9 1 10 11 1 10 9 2 7 1 11 2 3 1 10 0 9 1 10 11 0 2
19 4 4 3 13 10 9 0 7 0 13 1 10 9 12 1 10 9 11 2
24 10 9 4 4 13 7 1 9 1 9 0 1 10 9 7 1 9 1 10 9 1 10 9 2
31 3 1 10 9 12 1 10 9 11 2 10 9 7 10 9 1 10 9 4 13 1 0 9 1 10 9 7 10 9 9 2
68 10 9 1 10 9 1 10 9 7 1 0 9 1 9 4 13 1 10 9 1 9 1 10 9 1 10 9 2 1 15 13 9 9 1 10 10 9 9 7 1 10 9 9 7 1 15 13 9 1 11 2 1 10 11 7 1 11 2 3 1 10 0 9 1 10 9 11 2
51 10 9 11 13 3 3 10 10 9 1 10 9 7 1 10 9 9 1 9 0 1 15 13 1 10 9 1 10 9 7 4 3 13 1 0 9 10 9 1 9 0 1 10 9 2 9 1 10 9 2 2
34 10 9 0 1 9 0 1 10 9 1 10 9 1 10 9 0 4 13 1 10 9 1 0 9 0 2 1 11 7 10 9 1 9 2
51 15 13 1 9 1 9 0 1 10 0 9 7 13 10 0 9 2 3 0 3 1 10 9 1 10 9 11 2 2 15 4 3 13 1 10 9 11 1 10 9 0 1 10 9 1 9 1 10 9 9 2
36 3 1 10 10 9 1 9 7 9 2 10 9 1 10 9 11 4 13 10 9 0 7 1 0 9 7 1 10 9 9 7 1 10 9 0 2
5 1 13 15 15 2
17 1 10 9 4 4 13 9 0 0 1 10 9 1 10 9 0 2
25 12 9 11 4 13 10 9 2 1 10 9 2 1 9 1 9 1 13 10 9 1 10 9 0 2
19 4 4 13 10 9 1 9 1 10 9 0 1 10 9 7 1 10 9 2
40 3 1 10 0 9 7 1 10 9 1 10 9 1 10 9 1 10 9 11 2 10 0 9 4 13 1 10 9 0 1 10 9 7 1 10 9 1 10 9 2
86 3 1 10 9 12 1 10 9 9 12 5 12 5 11 1 10 9 2 1 10 12 9 12 2 15 13 10 9 1 9 1 9 1 9 2 9 7 9 1 10 9 1 10 9 1 10 9 0 2 9 2 11 2 2 7 1 10 9 1 10 9 1 9 1 10 9 11 1 10 12 9 12 2 15 13 16 10 9 1 10 9 4 13 7 13 2
27 10 9 1 9 13 13 1 12 9 2 7 10 9 1 9 0 13 0 1 12 9 1 11 1 10 9 2
5 10 9 13 13 2
13 10 9 1 10 9 1 9 13 1 10 9 0 2
20 10 9 1 10 9 1 10 9 1 10 9 13 1 10 9 9 7 0 9 2
28 3 10 9 1 10 9 1 10 9 0 7 0 1 10 9 0 1 10 9 1 9 2 1 10 9 1 11 2
23 3 3 1 10 9 1 10 9 1 10 9 11 2 13 0 13 10 9 13 10 9 1 2
40 2 13 10 9 0 1 13 7 13 10 0 9 1 10 9 1 10 9 1 9 7 13 10 9 1 10 9 1 10 9 1 9 15 13 10 9 1 10 9 2
38 2 13 9 5 9 1 10 9 1 0 9 7 13 10 9 3 1 10 9 15 4 3 13 1 10 9 11 2 9 0 2 0 9 7 9 0 2 2
31 2 13 9 1 10 9 0 3 1 10 9 1 10 9 1 9 1 10 0 9 2 15 4 13 1 10 9 1 10 9 2
33 2 13 3 1 10 9 7 1 10 9 0 1 10 0 9 9 2 13 10 9 1 10 9 15 1 15 13 10 9 1 9 0 2
20 9 1 10 9 1 9 1 10 9 1 10 9 12 7 12 1 10 9 11 2
12 2 9 1 10 15 10 9 3 13 9 2 2
20 10 9 0 1 10 9 13 1 12 9 1 11 2 3 12 9 1 9 2 2
25 10 9 1 10 9 1 10 9 13 9 2 1 9 1 10 9 0 2 13 0 1 10 9 5 2
50 9 1 10 9 0 13 10 9 12 5 12 2 11 1 10 9 0 7 1 10 9 2 1 10 12 9 12 2 0 1 10 9 1 9 7 1 9 1 10 9 1 10 9 2 9 7 9 1 9 2
24 2 9 0 1 10 9 1 9 0 1 10 9 1 9 0 7 0 13 11 1 10 11 2 2
66 1 9 13 10 12 9 12 2 10 9 11 11 11 2 1 9 0 1 12 9 11 11 2 11 2 12 2 11 2 2 7 11 11 11 2 1 9 0 1 11 12 2 11 2 12 2 11 2 2 4 13 10 9 0 1 12 9 1 10 9 1 9 0 7 0 2
34 10 9 2 13 2 11 11 11 11 2 2 13 10 9 1 3 12 9 0 2 13 1 10 9 1 10 9 1 10 11 2 11 2 2
10 10 9 13 1 9 13 15 1 11 2
95 10 9 0 4 13 13 9 1 10 9 1 12 9 1 13 1 10 9 1 10 0 9 2 13 10 9 13 1 10 2 9 0 1 10 9 1 9 0 1 9 1 11 2 13 1 10 9 0 1 10 9 0 9 8 12 1 10 12 9 12 2 9 12 2 7 13 1 10 9 0 12 2 12 1 10 12 9 12 0 1 10 9 0 2 11 0 1 10 11 11 1 10 12 2 2
53 9 1 10 9 2 1 10 12 9 12 2 13 10 9 1 9 1 9 0 13 1 10 9 1 10 9 1 10 9 1 9 1 11 2 1 10 9 11 2 11 11 2 1 9 1 10 9 12 1 10 9 11 2
13 2 10 9 1 9 0 13 10 0 13 9 2 2
57 1 9 12 9 12 10 9 0 4 13 1 10 9 1 10 11 11 2 1 9 1 10 9 12 1 10 9 11 2 10 9 0 1 10 9 0 1 10 9 1 9 0 13 1 10 9 1 10 9 1 10 9 1 9 1 11 2
50 1 10 9 1 10 9 7 1 10 9 0 13 1 10 9 10 12 9 12 7 13 1 10 9 1 10 11 11 10 12 9 12 2 7 16 4 13 10 9 1 9 2 10 9 4 13 10 0 9 2
26 8 2 10 9 1 10 9 7 10 9 9 3 0 2 1 10 9 10 11 2 13 1 3 12 9 2
31 8 2 1 9 0 0 2 10 9 1 9 0 7 0 3 13 1 0 9 9 10 9 1 10 9 0 1 10 9 0 2
33 10 9 0 7 10 9 1 9 3 0 2 13 1 10 9 1 9 2 4 13 1 10 9 1 9 0 7 1 10 9 7 9 2
27 15 13 1 10 9 1 10 9 13 1 10 9 1 10 9 0 1 9 2 9 12 5 12 2 11 2 2
18 13 10 9 1 10 9 0 16 10 9 0 15 4 13 1 10 9 2
7 11 1 9 1 10 9 2
11 13 1 11 10 9 1 10 9 1 9 2
8 10 9 1 11 13 1 9 2
13 13 10 9 0 10 0 9 3 1 13 1 11 2
11 10 9 1 10 9 2 1 9 11 11 2
33 15 13 3 2 9 1 15 2 2 3 2 1 10 9 15 13 10 9 1 10 9 2 15 13 9 2 9 1 9 7 9 0 2
23 11 13 1 9 1 10 9 2 3 1 10 9 2 10 9 4 13 2 13 1 10 9 2
9 10 9 1 9 13 1 10 9 2
35 11 2 11 2 11 2 10 9 1 10 10 2 9 0 2 13 2 10 9 1 10 9 7 1 10 9 1 9 2 10 9 2 10 9 2
27 15 13 10 9 0 2 13 10 9 13 1 9 1 9 13 2 9 7 9 1 9 13 1 13 10 9 2
13 13 9 7 9 2 3 1 10 9 7 10 9 2
13 1 10 9 1 10 9 3 15 13 15 7 15 2
25 3 4 13 10 0 9 1 10 9 3 0 2 10 9 0 1 10 9 0 1 10 9 11 11 2
67 7 3 10 9 13 9 0 7 15 4 13 1 10 9 1 10 9 0 2 13 1 10 9 7 10 9 2 13 1 10 9 1 10 9 11 2 15 1 15 3 1 9 1 9 7 15 13 10 0 9 1 11 11 2 9 1 10 9 12 13 1 10 9 1 11 11 2
31 10 9 4 4 13 1 10 9 2 4 13 11 11 2 10 9 1 11 7 1 10 15 13 1 10 9 1 10 10 9 2
44 11 10 9 3 15 13 1 11 7 3 1 10 9 2 3 13 1 10 9 1 9 1 10 9 2 4 13 1 15 7 1 10 10 9 10 9 1 0 13 1 10 9 13 2
3 7 3 2
55 3 15 4 13 10 2 9 2 1 3 12 9 1 9 13 1 10 9 1 10 11 3 4 13 10 9 1 10 0 9 7 3 9 1 9 1 9 0 2 1 10 9 2 1 10 9 2 1 10 9 1 10 9 0 2
18 3 4 4 13 10 9 1 10 9 0 2 7 3 3 1 15 0 2
24 10 9 1 9 13 0 7 4 3 13 7 13 1 9 2 0 9 1 10 11 2 9 0 2
33 3 10 9 1 9 3 2 16 3 15 13 3 1 9 2 11 4 13 3 10 9 1 10 9 7 3 10 10 9 1 10 9 2
16 10 0 9 1 10 9 0 15 13 10 9 13 1 10 9 2
19 3 15 13 10 9 0 1 13 3 13 1 11 10 9 1 10 9 0 2
11 10 11 11 1 11 11 1 10 11 13 2
23 10 9 1 10 9 0 1 11 13 0 2 10 9 1 10 9 0 0 1 10 10 9 2
20 13 1 10 9 1 3 13 10 9 1 9 1 10 9 1 15 1 10 9 2
16 7 11 13 3 10 9 1 10 9 0 1 10 9 1 9 2
41 10 9 1 10 9 4 13 1 11 11 2 10 9 15 1 10 12 13 1 10 0 9 10 9 0 16 10 9 1 10 9 13 3 1 10 9 1 10 9 0 2
44 1 10 12 10 9 0 2 1 10 9 0 2 4 13 1 9 2 16 1 10 0 9 0 1 10 9 0 1 10 9 1 10 11 11 15 13 10 9 1 9 1 10 9 2
58 3 15 10 9 1 10 9 1 9 1 10 9 2 10 0 9 1 9 3 15 4 13 1 9 1 10 9 1 11 11 2 13 15 10 9 1 9 1 9 13 1 10 9 0 1 10 9 0 1 12 9 2 10 9 1 10 11 2
60 3 10 9 15 4 13 1 10 9 0 1 10 9 1 10 9 1 13 15 1 10 9 1 11 11 2 10 9 1 10 9 2 13 1 10 9 0 1 10 9 0 1 11 11 7 1 9 0 2 13 3 1 10 0 9 1 10 0 9 2
48 1 3 4 13 10 9 1 10 9 15 13 10 9 0 2 13 7 13 16 3 4 13 10 9 3 1 10 9 2 15 1 10 9 1 10 9 0 4 13 10 0 9 1 10 9 1 11 2
18 1 9 11 7 10 9 2 13 10 0 11 16 13 13 15 10 9 2
28 3 3 15 13 3 10 9 1 10 9 0 15 3 1 11 4 13 10 0 9 1 10 12 5 1 10 9 2
29 3 11 11 2 0 0 0 9 2 10 9 9 1 10 9 1 9 2 13 10 9 7 15 13 1 9 1 9 2
8 10 9 3 13 3 10 9 2
8 15 13 10 9 1 10 9 2
38 7 3 13 9 0 1 10 9 1 10 0 2 9 0 2 2 15 15 1 9 1 10 0 9 15 4 13 1 10 9 7 15 3 4 13 10 9 2
26 16 13 10 9 1 10 9 2 3 10 9 1 11 2 1 11 7 1 10 9 4 13 15 1 11 2
54 10 9 13 2 3 13 1 13 10 9 1 9 13 2 15 13 3 10 9 1 10 9 16 10 9 2 15 13 1 10 11 10 9 1 9 1 10 0 9 1 10 9 1 11 0 2 13 1 10 9 0 1 9 2
13 7 1 10 9 1 10 9 15 13 9 1 9 2
7 10 9 1 11 4 13 2
7 10 9 0 13 1 11 2
23 1 10 9 1 11 15 4 13 10 15 1 10 9 15 13 10 9 1 10 9 0 0 2
19 1 13 10 9 4 13 10 9 1 10 11 1 10 9 0 1 10 9 2
49 7 10 9 2 15 13 1 9 10 0 9 1 10 9 1 9 2 4 4 13 1 10 9 0 0 2 11 11 11 2 7 1 10 9 1 10 9 0 0 2 11 2 1 10 9 2 11 11 2
40 13 9 1 10 9 1 10 9 0 1 10 9 1 10 9 0 4 13 11 2 13 16 10 11 4 3 13 9 1 9 7 4 13 3 10 9 1 10 9 2
15 1 10 9 0 3 4 13 1 13 10 9 2 4 13 2
29 11 4 13 15 13 1 10 9 1 10 9 2 13 15 1 13 16 1 10 9 0 9 13 1 9 3 1 11 2
6 3 4 13 1 3 2
34 9 3 2 4 13 10 9 1 10 11 2 3 1 11 15 13 9 15 13 10 9 1 10 12 5 0 1 15 13 15 10 10 9 2
14 3 15 13 10 9 2 15 13 3 10 9 1 9 2
14 10 9 13 3 10 9 1 13 15 1 10 9 0 2
36 0 1 10 9 7 1 10 9 1 10 11 2 1 10 9 1 9 1 9 2 13 1 10 9 0 15 15 13 1 10 0 9 1 10 9 2
15 15 13 10 9 0 15 4 13 10 9 1 10 12 9 2
12 15 9 1 15 13 10 0 9 1 10 9 2
26 15 13 13 1 10 9 1 10 12 1 11 7 11 13 1 10 9 1 10 9 2 1 9 7 9 2
25 7 3 10 9 2 3 13 10 9 0 2 15 13 16 1 10 0 9 1 10 9 13 10 9 2
45 10 9 2 7 3 1 0 9 2 1 10 2 11 11 2 13 3 16 3 1 13 4 4 13 1 9 10 9 0 1 13 3 13 10 9 2 13 1 10 9 7 1 10 9 2
7 15 13 10 10 9 0 2
49 1 10 9 1 10 9 15 3 13 10 9 13 10 9 1 10 9 0 2 10 9 1 10 9 1 9 3 0 1 10 9 2 10 9 1 15 1 11 4 13 1 10 9 1 11 1 10 12 2
23 10 11 13 7 13 10 9 1 10 9 2 10 9 7 10 9 13 1 10 9 1 9 2
10 3 10 9 4 13 1 13 10 11 2
8 10 0 9 3 4 13 0 2
29 1 10 9 1 11 10 9 4 4 13 1 10 9 0 1 10 9 1 10 11 2 9 13 1 10 0 9 0 2
39 7 10 9 15 13 3 3 1 10 9 1 10 9 13 2 1 9 1 9 0 7 3 0 2 1 10 9 15 1 12 9 1 9 15 13 1 10 9 2
15 3 1 10 9 0 2 10 11 13 3 1 13 1 11 2
12 1 10 12 1 10 12 4 4 13 12 9 2
42 3 1 13 10 9 1 10 9 0 10 9 4 13 2 1 10 0 9 1 9 2 1 13 10 9 0 2 15 0 2 1 13 0 10 9 7 10 9 11 2 11 2
7 3 4 13 10 9 0 2
44 10 9 3 13 0 7 15 13 1 12 2 12 9 1 9 2 1 3 12 12 9 0 7 15 1 10 9 7 1 10 9 1 10 12 5 1 10 9 1 10 9 0 0 2
21 10 11 13 3 9 1 0 9 1 15 15 1 13 1 13 10 9 1 10 9 2
52 15 3 4 13 13 10 9 1 1 10 15 7 13 2 3 1 10 9 0 7 1 10 9 0 2 10 9 0 7 0 0 1 13 1 10 9 1 10 2 9 2 2 13 10 9 0 7 10 0 9 0 2
13 1 10 9 13 15 4 13 10 9 0 7 0 2
42 13 10 9 11 11 1 10 9 1 10 9 7 10 9 1 10 11 2 15 13 1 10 0 9 1 10 9 2 1 13 1 9 1 10 11 15 13 1 3 12 9 2
32 16 10 11 11 2 15 4 13 3 11 16 4 15 13 1 9 2 13 10 9 2 3 10 9 0 4 13 10 9 3 0 2
23 3 2 3 1 10 9 13 1 0 2 9 2 0 2 15 13 10 0 9 1 9 0 2
23 12 9 3 11 11 2 10 2 9 2 2 13 1 10 9 16 10 10 9 0 4 13 2
13 10 9 4 13 3 2 1 10 9 1 10 11 2
23 11 13 10 2 9 2 1 11 7 13 1 13 10 9 15 1 10 9 0 3 13 15 2
32 10 9 2 13 2 13 9 1 10 12 5 1 10 9 1 10 9 13 1 10 10 9 7 13 1 13 1 15 1 13 0 2
14 2 3 1 15 2 13 2 15 13 10 9 0 2 2
33 7 10 9 2 13 0 11 2 15 15 4 13 12 12 9 15 4 13 1 10 11 2 7 3 15 15 4 13 1 9 10 9 2
52 10 9 1 10 9 4 13 10 9 1 10 9 7 16 4 13 1 10 0 15 1 0 7 0 9 2 7 1 15 3 15 13 3 10 9 1 11 2 4 3 13 1 10 9 1 10 9 0 0 7 0 2
35 1 11 7 11 2 1 9 7 1 9 0 2 13 1 10 9 1 11 7 11 9 0 1 9 2 13 1 9 7 9 1 10 9 13 2
22 1 10 9 13 16 4 13 10 9 1 9 0 2 13 1 10 9 9 15 13 0 2
8 15 13 9 0 1 10 9 2
35 10 9 2 1 9 2 13 13 9 2 9 7 0 9 1 9 2 1 10 9 0 15 1 10 9 13 12 7 1 9 3 12 9 0 2
32 9 13 15 13 10 9 1 0 9 1 9 1 10 9 1 10 15 2 1 10 9 1 10 15 2 1 10 9 1 10 15 2
26 1 10 9 3 0 1 11 7 1 10 9 3 13 1 13 1 10 9 1 10 9 2 13 9 0 2
44 1 11 4 13 9 1 9 1 12 9 1 9 7 15 4 13 2 13 10 9 1 10 9 0 2 13 1 10 9 1 9 3 0 3 1 10 9 1 10 9 1 9 0 2
28 13 0 16 1 10 9 15 4 13 9 13 2 7 3 3 13 10 9 16 10 10 9 1 9 13 1 11 2
27 15 13 11 11 2 9 1 10 9 11 2 13 3 9 1 10 9 1 10 9 0 1 10 9 11 11 2
42 1 10 9 13 1 13 10 9 0 1 11 2 13 11 2 4 4 13 10 9 15 4 13 1 13 0 9 0 2 3 10 9 1 9 0 7 10 9 0 1 9 2
5 7 13 10 9 2
11 10 9 1 10 9 3 13 0 1 13 2
15 10 9 1 11 4 13 10 9 0 1 10 9 0 0 2
10 13 15 15 15 1 9 13 1 3 2
16 15 15 13 2 13 16 13 1 10 9 7 15 15 4 13 2
31 1 10 9 1 10 2 9 2 1 9 13 1 9 1 10 9 2 1 15 13 10 9 7 13 1 10 12 5 10 9 2
21 3 2 1 10 9 1 10 12 2 4 13 1 13 9 7 9 13 15 1 15 2
16 10 9 1 10 9 0 0 13 1 10 12 1 10 12 9 2
17 3 1 3 13 10 9 13 1 10 9 2 9 2 9 2 9 2
11 12 9 1 13 10 0 9 1 10 11 2
23 1 10 9 1 11 1 10 11 1 13 10 9 2 10 9 0 4 13 1 13 10 9 2
25 1 10 12 1 12 9 4 4 13 12 9 2 10 9 0 15 10 9 1 11 3 4 3 13 2
17 10 9 1 9 2 3 15 1 12 2 4 4 1 9 13 13 2
25 1 11 2 3 3 4 4 13 10 0 9 1 9 15 4 13 12 9 2 10 9 13 3 0 2
19 7 1 9 10 9 1 9 1 10 9 1 9 4 4 13 1 10 9 2
28 10 9 1 9 15 4 13 16 15 4 13 10 9 2 0 2 16 4 4 13 10 9 3 1 10 9 0 2
21 10 9 3 4 13 2 7 4 4 13 1 9 10 9 1 10 9 1 10 9 2
9 1 10 9 10 9 3 13 3 2
28 3 4 13 3 1 10 0 10 10 9 1 13 10 9 1 10 9 0 2 1 15 1 10 9 1 10 9 2
24 15 15 3 4 13 10 10 9 1 10 9 15 4 13 9 0 1 10 9 2 9 2 9 2
18 10 3 0 4 13 1 13 10 9 1 11 2 1 9 1 10 9 2
22 9 0 2 3 10 9 15 13 10 9 1 11 11 7 3 15 1 10 9 11 11 2
23 1 10 9 2 3 1 13 1 10 2 9 1 10 9 2 2 15 13 10 9 1 11 2
31 13 10 9 2 11 4 13 1 10 9 1 13 10 9 1 9 13 1 10 9 15 1 10 9 3 1 9 1 10 9 2
23 10 0 9 2 15 1 10 9 1 9 13 12 9 10 9 1 9 1 10 9 1 9 2
28 11 1 10 9 13 10 0 9 0 1 10 9 1 10 9 1 10 9 0 2 0 7 3 9 1 12 9 2
22 3 15 13 10 9 0 1 11 11 13 1 10 9 15 13 1 10 9 10 10 9 2
22 1 10 9 0 1 11 7 11 2 1 10 9 1 10 12 11 13 1 13 15 3 2
18 7 10 9 13 1 9 7 13 10 9 1 13 15 15 13 12 9 2
30 11 13 1 13 15 3 7 3 4 13 10 9 1 11 7 1 10 9 1 10 9 2 7 3 3 11 15 4 13 2
12 15 13 3 10 9 1 10 9 11 7 11 2
23 10 9 13 13 2 1 3 2 13 9 0 2 13 13 10 9 7 13 1 13 10 9 2
6 7 10 9 13 0 2
18 3 10 9 11 15 4 13 10 0 9 1 10 0 9 1 10 11 2
29 13 0 10 9 1 11 2 16 10 11 13 10 9 1 10 9 15 13 7 15 13 9 1 9 1 10 9 0 2
51 10 9 1 10 9 2 15 4 13 1 13 1 9 10 9 1 9 2 4 13 1 10 9 0 1 13 10 10 9 1 11 1 15 13 1 9 0 2 1 10 9 1 10 9 15 4 13 1 10 9 2
16 1 10 9 1 9 0 2 3 3 10 9 13 0 1 9 2
52 1 11 10 9 4 13 0 9 13 10 9 1 0 9 2 16 15 1 10 9 1 10 9 1 10 9 2 9 4 4 13 1 10 10 0 9 1 4 13 1 10 9 0 1 15 13 9 3 9 1 9 2
14 1 11 11 10 9 4 13 1 10 9 1 10 9 2
13 10 9 1 10 9 13 1 10 9 1 10 9 2
10 10 10 9 4 3 13 1 10 9 2
13 15 13 15 3 7 3 13 1 15 1 13 15 2
5 15 13 1 15 2
36 13 1 10 9 2 16 10 9 0 15 13 1 10 9 2 16 10 9 1 11 2 11 11 13 10 0 0 9 1 12 9 1 10 9 12 2
16 3 1 10 9 0 1 9 13 1 13 10 9 1 11 11 2
33 9 2 9 1 10 9 11 11 1 10 9 0 1 15 13 9 2 11 13 3 0 1 11 2 3 13 10 9 1 10 9 13 2
28 10 9 1 10 9 3 15 13 2 7 4 13 10 9 1 15 7 10 10 0 9 1 10 9 1 10 9 2
6 15 13 10 9 0 2
33 13 15 2 1 15 10 0 9 11 11 2 13 1 10 9 1 10 9 0 2 1 9 1 15 1 11 11 2 10 2 9 2 2
6 13 10 9 3 0 2
11 4 13 10 9 1 9 7 1 10 9 2
6 0 16 13 10 9 2
19 4 13 10 9 1 10 9 1 10 9 7 3 13 16 4 13 10 9 2
10 13 1 3 16 15 13 10 9 0 2
2 15 2
42 1 11 15 4 13 10 9 1 10 9 7 10 9 15 4 13 10 10 9 0 2 1 10 9 2 1 10 9 2 1 10 9 7 1 10 9 2 15 13 10 9 2
15 10 9 1 15 1 10 9 4 13 10 9 1 10 9 2
37 7 10 9 11 4 4 13 1 9 1 11 3 16 4 13 1 13 10 9 0 2 1 10 9 1 10 9 1 10 9 1 10 9 1 10 9 2
22 10 9 4 4 13 1 13 10 9 1 13 10 9 0 3 16 4 13 0 9 0 2
9 10 9 0 7 0 3 15 13 2
22 1 9 15 4 13 1 10 9 0 15 13 1 15 7 1 10 10 9 1 15 0 2
20 16 13 0 15 15 13 2 3 15 13 3 3 1 13 9 7 10 0 9 2
13 11 13 0 2 13 11 2 13 10 9 3 0 2
16 10 10 9 0 13 15 1 13 3 10 10 9 0 7 0 2
15 7 13 16 15 13 10 9 1 10 9 1 13 10 9 2
51 1 9 1 10 9 1 10 9 7 1 9 0 15 13 10 9 1 11 2 1 11 15 13 10 9 15 4 13 1 3 13 10 9 2 16 3 15 13 2 7 1 13 1 9 10 10 9 1 10 9 2
19 13 11 11 2 9 1 10 9 2 10 9 15 13 10 9 1 10 9 2
33 11 2 9 1 11 0 2 4 13 10 9 9 1 15 4 13 1 4 13 1 15 1 10 9 13 1 10 9 0 12 12 9 2
13 9 0 2 7 3 3 1 10 9 0 1 11 2
15 3 4 13 10 9 1 10 9 7 3 13 13 10 9 2
22 4 13 3 2 1 10 9 13 2 7 11 3 15 4 13 7 4 13 10 9 0 2
17 9 13 1 10 9 2 13 15 3 7 13 1 13 1 10 9 2
44 15 13 10 9 16 1 13 10 9 1 10 9 1 11 11 0 2 10 9 15 4 13 10 9 1 9 2 3 13 7 10 9 7 0 9 7 13 3 10 9 1 9 0 2
8 9 1 12 2 12 12 9 2
43 6 1 10 9 0 2 1 0 9 2 2 12 2 12 12 9 2 2 3 16 4 13 2 1 10 9 1 9 2 10 9 1 10 9 0 1 10 9 0 1 10 12 2
21 10 9 1 10 9 12 2 1 10 9 1 10 9 2 13 3 0 7 3 0 2
16 4 13 3 1 10 11 1 11 10 0 9 1 10 11 11 2
8 3 10 0 9 1 11 11 2
20 10 9 1 11 11 11 15 4 13 1 10 9 0 1 10 9 0 9 9 2
14 0 9 1 11 11 0 1 10 9 0 1 10 9 2
19 9 0 1 10 9 1 10 9 1 10 11 1 9 1 10 9 1 9 2
21 10 9 1 10 9 13 1 13 12 9 1 13 10 9 1 11 7 1 10 11 2
12 10 9 1 10 9 4 3 13 10 0 9 2
38 1 10 11 1 11 10 9 0 1 10 9 4 13 10 9 1 10 9 1 9 7 3 1 10 9 1 9 1 10 9 9 2 3 1 10 0 9 2
7 2 9 1 9 12 2 2
9 1 9 10 9 0 13 10 9 2
10 6 13 0 2 13 10 9 0 2 2
17 10 11 4 13 10 9 0 1 10 12 5 1 10 9 0 0 2
11 15 13 3 10 9 1 9 1 10 9 2
34 9 1 10 11 2 3 10 0 9 1 10 9 1 10 9 0 1 10 9 2 10 9 1 12 9 1 9 10 9 2 13 3 13 2
7 10 9 4 13 1 3 2
21 10 9 0 0 2 0 2 0 4 13 1 13 10 9 1 10 9 0 1 9 2
38 10 9 1 10 9 11 11 4 13 3 2 1 10 0 9 9 1 10 9 2 10 9 1 10 9 2 15 3 4 13 9 1 9 0 7 1 9 2
22 13 1 11 10 9 1 10 9 11 0 1 13 10 9 1 10 9 1 10 9 9 2
26 10 9 4 4 13 1 11 11 2 9 1 11 1 10 9 0 1 10 9 1 10 9 2 11 11 2
21 10 9 1 9 2 12 2 12 9 1 9 2 13 1 13 10 9 1 10 9 2
9 10 9 0 1 9 1 10 11 2
14 10 9 1 9 3 0 1 10 11 3 4 13 9 2
66 10 9 1 10 9 2 10 9 1 10 2 9 0 1 11 2 2 10 9 3 1 10 9 15 13 1 10 9 0 1 10 9 0 2 9 7 9 1 10 9 1 10 9 1 9 7 9 0 2 13 11 1 13 1 9 1 10 9 1 10 9 7 10 9 0 2
37 1 10 9 0 4 13 10 9 1 10 9 0 1 10 9 1 13 1 9 10 9 1 9 0 7 0 13 1 13 10 9 1 10 2 9 2 2
20 10 9 4 4 13 1 10 9 1 11 1 10 9 0 7 10 0 9 9 2
41 10 9 2 13 3 1 10 11 2 4 13 1 10 11 11 15 10 12 9 1 10 9 1 10 9 1 10 9 13 1 9 1 10 9 10 9 1 10 9 0 2
31 10 9 2 1 10 10 9 10 9 11 11 2 4 13 3 1 13 10 9 1 10 9 1 10 9 3 0 1 10 9 2
52 3 15 13 3 10 9 0 1 10 9 1 10 9 7 1 10 9 1 10 9 0 15 13 1 10 9 1 12 2 12 9 1 9 2 13 3 1 13 10 9 1 10 9 0 13 1 10 9 1 10 9 2
35 10 9 1 10 9 2 1 10 0 9 4 13 10 12 5 1 10 9 2 13 10 9 0 1 13 10 0 9 1 10 9 1 10 11 2
15 7 1 9 1 9 0 3 4 13 10 0 9 1 9 2
19 9 1 0 9 13 1 10 9 0 4 13 10 9 1 9 1 10 9 2
54 10 9 13 3 3 1 10 9 2 7 3 1 9 0 7 0 1 9 1 10 2 9 2 1 9 1 9 2 9 1 10 9 1 9 2 1 10 9 2 1 10 9 2 1 10 9 2 1 10 9 1 9 0 2
16 13 10 9 2 13 13 10 9 2 13 10 9 1 10 9 2
15 4 3 13 3 15 15 4 13 9 1 12 2 12 9 2
32 11 2 13 10 9 1 10 9 11 11 2 13 9 1 10 11 11 1 10 9 1 9 13 1 13 10 9 1 9 3 0 2
12 9 1 9 7 9 1 10 9 1 13 9 2
46 11 2 13 12 9 3 1 10 9 1 10 9 1 11 2 13 3 9 1 10 9 0 15 15 4 13 1 4 13 1 10 9 1 9 2 0 1 10 9 0 1 11 7 0 11 2
30 10 9 13 1 10 0 9 2 3 13 3 10 9 7 13 0 1 10 9 0 2 13 1 11 15 15 15 13 3 2
15 1 10 9 0 13 9 2 9 2 9 7 10 9 0 2
15 10 9 13 0 2 0 3 1 10 3 0 1 10 9 2
36 3 4 13 10 9 1 9 3 0 1 10 9 2 13 3 13 1 10 9 2 1 10 9 2 15 13 10 9 0 0 1 12 9 1 9 2
45 1 10 9 2 11 13 1 10 9 1 10 9 1 10 0 11 2 13 1 10 9 7 1 9 0 1 10 9 2 4 13 10 9 1 9 1 9 1 10 0 12 2 12 9 2
36 3 10 11 3 13 3 15 7 3 9 1 10 9 2 9 0 1 9 0 15 4 13 9 7 9 1 10 9 13 1 12 9 1 9 13 2
36 7 15 4 3 13 15 1 10 9 3 0 1 10 0 9 2 16 10 10 9 0 3 4 13 1 10 9 7 15 13 1 10 10 10 9 2
18 3 15 13 10 9 2 2 0 2 16 3 13 10 10 9 1 9 2
14 10 2 9 2 4 13 10 9 1 12 9 1 9 2
19 3 15 13 1 11 2 3 1 10 2 9 2 4 4 13 10 9 0 2
23 7 3 1 11 15 13 3 15 2 16 13 10 9 0 11 11 2 15 13 3 3 0 2
53 10 11 2 15 1 10 0 9 0 13 3 0 1 11 2 4 13 3 1 13 10 9 1 10 9 1 10 9 15 15 4 13 10 10 9 7 1 13 10 9 1 10 9 1 15 4 13 3 1 12 12 9 2
21 10 0 1 4 13 2 10 9 13 3 2 13 15 15 4 13 3 1 12 9 2
32 10 9 2 13 1 11 1 10 9 1 10 9 2 11 11 2 4 13 13 10 9 1 10 9 1 10 11 1 10 9 9 2
28 10 9 13 1 10 0 9 0 7 0 2 13 1 10 10 9 10 9 1 12 9 2 9 0 7 10 9 2
25 1 15 10 9 9 1 10 9 4 13 0 2 16 4 13 10 0 9 2 0 1 9 0 0 2
30 10 9 4 13 0 7 4 13 10 0 9 1 9 1 10 0 9 10 10 9 13 1 13 13 10 9 0 1 11 2
50 1 10 0 9 10 11 4 13 10 9 0 1 13 1 13 10 9 1 9 2 13 3 10 9 1 9 7 13 1 10 9 3 10 9 2 13 3 1 10 9 1 10 12 1 10 12 5 10 9 2
49 1 10 9 1 9 4 13 1 11 10 9 0 15 4 13 10 9 1 13 11 1 10 9 1 10 9 2 7 3 13 0 16 10 9 13 3 1 10 9 11 4 13 10 0 9 1 10 9 2
35 1 10 9 1 10 9 10 9 0 4 13 10 9 1 10 9 1 10 9 1 9 13 1 10 9 1 11 1 13 10 9 1 10 9 2
32 1 16 4 13 10 9 0 1 10 9 1 10 9 0 15 13 3 10 9 2 13 1 9 2 3 2 1 10 0 9 0 2
14 10 9 0 4 13 1 11 7 13 3 16 4 13 2
45 1 15 10 9 0 1 15 4 13 3 13 11 11 2 10 9 0 1 10 9 1 11 2 9 1 10 9 0 1 10 9 2 3 10 12 5 1 10 9 0 2 12 9 2 2
11 15 13 10 9 1 10 0 2 9 2 2
57 3 13 10 9 1 1 15 2 13 1 10 9 1 11 11 10 9 11 11 2 9 1 10 0 9 1 10 11 2 7 9 1 10 0 9 2 10 9 0 2 11 2 2 15 4 13 10 9 1 10 9 0 1 10 9 0 2
66 10 9 1 10 9 3 4 4 13 1 10 9 0 2 3 13 1 13 15 1 9 0 2 13 10 9 0 1 10 9 1 11 2 11 11 2 9 1 10 9 0 2 11 2 2 0 1 10 9 0 1 11 2 7 3 1 10 9 0 15 13 3 1 10 9 2
36 1 10 9 0 10 9 1 11 11 2 3 13 1 4 13 10 9 1 11 1 13 10 9 1 10 9 0 1 11 2 13 13 9 3 0 2
19 10 9 13 12 12 2 13 2 13 1 9 0 2 1 11 7 1 11 2
23 10 9 1 10 9 13 1 10 9 0 0 1 10 11 11 7 1 10 9 0 1 11 2
5 10 9 13 0 2
30 10 9 1 9 4 13 1 10 9 1 10 9 0 7 15 3 13 3 10 0 9 16 13 10 9 1 10 9 0 2
8 15 13 10 9 1 10 11 2
29 10 9 1 10 11 1 10 9 0 2 10 10 9 0 4 13 1 10 9 0 1 10 11 2 10 9 0 2 2
21 15 3 13 1 11 7 16 13 1 13 15 7 3 15 13 13 3 15 10 9 2
14 4 13 10 10 9 0 1 10 9 1 9 0 0 2
7 11 3 15 4 13 9 2
6 3 4 13 0 9 2
8 13 10 9 2 7 10 9 2
30 4 13 10 10 9 0 2 15 15 13 1 10 9 0 1 10 9 7 3 15 15 13 3 9 1 10 9 1 11 2
19 10 10 9 4 13 10 9 1 9 0 7 10 9 13 1 10 15 0 2
25 15 13 10 9 13 1 9 2 13 2 1 9 0 7 10 15 0 2 9 1 9 7 9 0 2
10 10 9 13 9 13 1 10 9 0 2
19 15 2 1 9 2 4 13 1 10 9 0 13 1 10 11 1 10 9 2
12 4 4 13 15 16 15 4 13 1 10 9 2
21 3 4 13 1 10 12 2 4 4 13 7 3 13 1 12 9 1 9 1 11 2
15 7 13 2 10 9 4 13 1 9 15 13 10 9 10 2
18 10 9 1 10 9 1 10 9 1 11 4 4 13 1 10 9 13 2
7 10 9 13 1 10 11 2
5 3 1 10 9 2
17 13 3 0 13 13 10 9 1 10 11 1 3 1 10 9 0 2
9 15 13 16 4 13 1 9 0 2
11 10 9 13 3 1 10 9 1 10 9 2
10 15 3 4 13 9 2 13 11 2 2
41 10 10 9 13 10 9 2 10 9 0 2 10 9 1 10 11 2 10 9 0 0 2 10 2 9 2 1 11 2 10 10 9 13 0 1 10 11 11 1 11 2
10 16 11 15 13 10 9 10 9 13 2
26 10 11 2 9 1 10 9 1 10 9 1 10 9 1 10 9 12 1 10 11 2 4 13 1 11 2
59 10 9 1 10 9 7 10 9 1 10 11 4 13 13 10 15 1 10 0 9 0 2 10 9 0 2 13 10 9 3 1 9 0 1 10 0 9 2 13 1 9 0 1 10 9 1 10 9 1 10 11 7 3 3 13 1 10 9 2
58 9 0 1 10 9 11 11 2 15 3 1 15 4 13 3 1 3 10 9 0 2 4 13 15 1 13 1 10 9 0 10 9 0 1 10 9 1 10 11 7 1 10 11 2 13 15 3 3 1 10 11 1 10 9 1 10 11 2
18 7 15 13 3 16 1 11 7 1 11 11 7 11 13 3 3 0 2
40 15 4 13 10 9 1 10 9 2 13 10 9 15 13 1 10 9 0 2 1 10 12 1 10 12 5 2 1 9 1 10 9 0 2 10 9 1 10 9 2
29 1 11 12 9 4 13 7 10 9 4 13 0 1 9 1 9 1 9 1 10 0 9 1 10 9 13 3 9 2
8 0 10 9 1 10 10 11 2
32 10 3 0 9 1 9 1 10 9 1 11 4 13 3 10 0 9 1 10 0 9 1 9 0 1 10 9 1 11 1 11 2
14 9 7 9 15 4 13 1 10 9 13 1 10 9 2
9 10 11 4 13 10 9 1 9 2
40 3 10 9 11 11 4 13 1 10 9 1 10 9 1 13 10 9 0 1 10 9 1 10 9 0 2 13 1 10 9 11 1 10 9 0 7 10 9 0 2
40 11 7 11 1 10 9 0 1 10 0 9 1 10 11 1 13 10 9 1 9 1 10 9 1 11 1 10 9 2 1 10 11 2 1 3 12 9 1 9 2
48 10 9 1 10 11 11 1 10 0 9 12 4 4 13 1 10 9 1 10 12 1 10 12 5 2 1 9 1 10 9 1 10 9 1 9 2 13 1 10 12 5 10 9 1 10 0 9 2
33 13 10 9 1 10 9 11 2 1 3 0 1 12 9 1 9 16 10 9 13 1 10 9 2 16 13 1 10 9 1 10 9 2
27 1 3 9 1 10 11 3 0 1 9 0 1 10 12 5 1 10 9 9 7 1 10 9 11 7 11 2
18 10 9 4 13 1 10 9 1 10 9 0 7 10 9 1 10 9 2
37 10 9 1 10 11 2 11 11 2 4 13 10 12 5 1 10 11 2 10 9 9 1 9 1 10 9 11 7 15 13 9 1 10 9 11 11 2
26 9 0 1 10 9 1 10 9 1 10 12 9 1 9 1 10 9 1 15 10 9 4 13 10 9 2
17 9 11 11 0 13 11 1 10 12 1 10 12 1 10 0 9 2
8 9 1 9 0 1 10 11 2
29 1 12 9 1 9 1 10 9 1 10 2 9 2 0 2 10 11 4 13 1 10 9 1 10 9 1 10 9 2
21 1 11 10 9 4 13 1 9 1 10 9 7 9 1 9 1 10 9 1 9 2
38 12 9 4 4 13 2 12 13 1 10 9 1 10 10 9 13 1 10 9 2 10 15 13 1 10 9 0 2 12 9 13 1 9 1 9 1 9 2
39 9 1 9 4 13 1 9 1 10 0 9 1 10 9 2 1 11 9 7 9 15 4 13 3 1 10 9 3 1 10 12 13 10 9 1 10 9 0 2
19 3 10 0 9 11 11 4 13 10 9 1 10 9 1 10 9 11 11 2
54 9 7 9 2 15 1 9 2 7 1 10 9 0 1 10 9 0 13 10 9 0 2 13 10 9 1 10 9 1 10 9 0 13 0 1 10 9 1 10 9 0 3 4 4 13 12 9 1 9 1 9 7 9 2
50 1 11 10 9 4 13 1 10 9 0 13 1 10 9 2 1 10 0 9 2 1 9 0 15 3 13 10 9 1 9 1 9 13 15 4 13 1 10 9 1 10 9 1 10 9 1 10 9 0 2
43 1 11 10 9 1 10 9 7 10 9 1 10 11 2 10 9 0 15 4 13 10 9 1 10 0 11 2 3 4 13 1 13 10 9 1 12 9 7 10 9 13 0 2
14 10 9 13 10 9 7 13 10 9 0 2 0 2 2
43 10 11 13 3 3 0 1 10 9 0 7 15 13 1 13 2 1 10 9 7 1 10 9 2 1 10 9 2 1 10 9 2 0 1 10 9 11 11 13 3 1 9 2
17 11 13 10 9 0 1 10 9 15 13 10 0 9 1 10 9 2
17 7 3 13 10 10 0 9 2 3 13 3 10 9 1 0 9 2
13 9 1 10 9 1 11 1 13 15 9 7 9 2
13 13 1 10 0 2 9 10 9 1 10 9 0 2
8 10 9 13 3 1 10 9 2
38 10 9 1 10 9 0 2 12 9 1 9 1 9 2 3 10 9 0 1 10 9 0 1 11 2 9 0 1 3 2 9 1 9 2 9 7 9 2
26 1 10 9 1 10 11 2 1 12 9 1 10 9 0 2 10 11 13 1 10 9 1 10 9 0 2
29 1 10 9 2 1 3 3 0 7 3 0 2 1 10 0 9 0 1 10 12 9 1 9 0 13 1 11 11 2
32 7 10 9 0 2 1 10 9 7 1 10 9 2 4 4 3 13 1 10 9 1 10 9 0 1 10 9 0 1 10 12 2
41 10 9 1 10 9 0 2 13 1 10 9 7 13 3 1 10 11 11 2 10 0 9 1 11 2 4 13 10 9 0 1 10 9 15 3 4 13 1 10 9 2
35 1 9 1 10 9 1 11 15 4 13 1 10 0 9 1 9 10 9 13 1 10 0 9 2 0 7 1 10 9 1 9 1 1 9 2
18 15 4 13 9 1 10 0 9 7 10 9 1 9 1 10 9 0 2
18 7 3 1 13 1 10 9 10 11 4 13 1 9 1 10 9 0 2
51 1 10 9 10 9 1 10 0 11 7 10 9 2 1 10 9 1 9 2 1 15 0 1 10 9 2 4 13 2 3 1 10 9 1 10 9 2 10 9 1 10 9 7 13 10 9 1 10 9 0 2
24 1 10 9 1 10 11 7 10 11 1 10 9 4 13 1 15 2 1 10 9 1 10 9 2
12 11 3 15 4 13 1 10 11 1 10 11 2
36 3 13 10 9 10 9 13 1 10 0 11 15 1 10 9 4 13 3 1 10 9 1 11 10 9 1 9 1 10 9 1 9 7 1 9 2
16 10 9 7 10 0 9 4 3 13 1 10 9 1 10 9 2
42 15 1 10 9 2 9 2 1 13 0 9 2 4 13 1 10 9 1 10 9 0 15 3 1 10 9 0 1 11 11 4 13 10 9 1 9 1 10 10 9 0 2
34 10 9 1 10 9 4 13 15 15 1 15 2 9 3 1 10 9 1 10 9 7 1 10 9 1 10 11 2 4 13 1 10 9 2
35 3 13 10 9 16 3 4 13 10 0 9 13 1 13 2 1 0 9 1 9 2 9 0 7 1 13 9 0 2 1 3 3 3 0 2
40 1 10 9 0 4 13 15 0 2 9 0 2 9 2 9 2 13 3 1 10 9 15 15 4 13 2 1 10 9 1 9 2 3 10 9 1 9 1 9 2
26 10 9 0 1 10 9 1 12 9 1 9 1 10 9 1 12 9 7 10 9 0 0 1 12 9 2
27 1 10 9 1 10 9 0 7 0 10 9 0 2 7 3 3 15 2 7 10 11 4 13 10 0 9 2
39 9 7 9 15 4 13 1 10 10 9 1 10 9 7 1 10 9 0 2 1 10 9 1 9 2 7 3 1 9 2 15 4 13 3 1 10 9 3 2
10 10 9 15 4 13 1 12 9 0 2
27 1 11 7 10 0 9 1 9 1 10 0 11 15 4 13 10 9 0 1 10 9 13 1 13 10 9 2
25 10 9 0 2 15 4 13 1 9 0 9 0 2 1 15 0 2 13 1 10 9 1 2 9 2
21 10 9 1 11 2 1 9 0 2 4 4 3 13 1 13 1 13 10 9 0 2
22 9 1 9 7 9 4 13 10 9 1 10 9 1 10 9 7 10 9 1 10 9 2
18 3 15 4 13 10 9 13 1 9 1 10 9 0 1 10 9 0 2
17 10 9 1 10 9 1 10 9 7 10 10 9 4 13 10 9 2
13 1 13 10 9 2 11 3 13 1 9 12 9 2
24 10 9 1 10 0 9 11 11 7 10 10 9 1 10 9 2 1 10 9 13 3 1 9 2
34 16 13 1 13 10 9 1 10 9 2 3 13 1 9 1 13 10 9 1 10 9 0 1 13 3 10 9 1 10 9 0 1 11 2
38 7 16 4 13 1 10 9 1 10 9 1 10 9 15 15 4 13 1 10 10 9 2 3 3 10 11 3 2 0 13 9 1 10 9 1 10 11 2
43 10 2 9 1 10 9 2 1 10 9 11 11 7 10 9 1 10 9 0 4 13 1 9 3 12 9 0 7 12 1 9 0 13 1 10 9 1 10 9 0 1 11 2
37 10 9 1 9 4 13 3 12 9 7 4 4 13 1 9 0 1 10 9 2 9 7 9 1 10 9 0 13 3 1 10 9 0 1 11 11 2
15 1 11 3 10 9 1 10 9 4 13 1 10 9 0 2
50 10 9 11 2 13 3 1 12 9 1 10 9 2 4 13 2 16 4 13 10 9 2 1 13 10 9 0 1 10 9 1 10 9 2 1 9 1 11 3 13 1 9 10 9 0 1 10 9 0 2
17 10 9 1 9 1 9 0 4 4 13 1 10 9 1 9 0 2
16 10 9 1 11 4 13 10 0 9 1 10 10 9 1 9 2
49 10 9 13 0 1 10 9 1 10 9 1 10 9 1 9 0 13 1 9 1 10 9 1 11 7 11 2 3 1 10 9 13 1 10 9 13 10 9 13 1 9 1 9 7 9 0 1 9 2
2 9 2
17 15 13 1 13 3 3 2 13 15 1 10 9 1 10 9 2 2
69 10 9 1 13 10 9 1 10 9 13 1 10 9 1 10 9 2 10 0 9 1 10 9 15 13 3 1 13 1 9 7 10 9 4 3 13 10 9 1 13 1 11 2 1 9 9 1 10 9 1 11 3 1 9 1 10 9 2 1 1 10 9 10 10 9 1 10 11 2
45 10 0 9 15 4 13 11 2 1 10 9 9 0 1 10 9 0 2 4 13 10 9 1 11 11 2 10 9 1 9 0 15 4 13 3 1 13 3 10 9 1 13 10 9 2
8 1 15 3 15 13 3 9 2
19 10 10 9 0 7 1 9 4 13 1 11 11 2 9 1 10 9 0 2
44 15 13 15 1 10 9 1 10 9 1 10 9 1 9 2 3 1 10 9 2 1 10 12 1 9 1 10 12 1 10 9 2 7 1 10 9 13 3 1 10 9 1 9 2
43 10 9 1 10 0 9 0 11 11 2 13 1 10 9 0 2 0 11 11 2 4 4 13 1 10 9 1 12 0 9 13 1 9 0 1 9 0 13 1 15 1 9 2
17 10 9 15 13 1 10 9 1 10 9 7 10 10 9 4 13 2
33 13 10 9 1 10 9 1 10 9 0 7 10 9 1 11 2 11 2 2 13 10 9 11 2 16 15 13 3 1 9 13 2 2
18 4 3 13 10 9 7 10 15 15 13 1 10 0 1 10 9 0 2
12 10 9 2 3 15 0 2 13 3 1 9 2
37 10 9 2 3 10 9 1 10 0 9 1 9 1 11 2 3 15 1 10 11 1 11 2 9 0 1 10 9 1 10 9 2 15 13 3 13 2
8 10 0 9 0 1 10 11 2
30 1 11 1 10 9 1 10 2 9 2 7 10 9 1 10 9 13 1 9 10 9 1 10 9 3 3 15 13 9 2
10 3 1 10 9 0 13 4 13 0 2
24 1 3 10 10 9 2 11 13 2 3 13 3 9 16 4 4 13 10 9 1 9 1 9 2
60 1 10 0 9 2 1 11 2 10 9 0 13 1 9 3 4 13 3 10 0 9 1 10 9 0 1 10 11 16 10 9 1 11 2 15 1 10 9 1 10 9 15 4 13 3 12 12 9 7 9 1 9 2 4 13 10 10 9 0 2
23 10 9 1 10 9 0 15 4 13 3 1 13 10 9 3 1 10 9 13 9 1 9 2
38 10 9 0 1 10 9 2 0 1 10 9 1 10 9 7 13 1 10 9 0 13 1 10 9 7 1 10 9 1 9 0 2 13 1 13 10 11 2
17 3 4 13 1 9 10 9 2 13 10 9 1 10 9 11 2 2
22 1 15 10 9 15 4 13 1 10 0 9 3 3 1 11 7 3 1 11 7 11 2
22 4 13 10 9 1 10 0 12 9 16 4 13 16 4 13 15 13 10 9 1 9 2
15 7 10 9 1 11 9 4 3 13 1 12 9 1 11 2
14 16 3 4 13 1 9 10 9 3 13 1 10 9 2
6 7 3 15 10 9 2
30 1 10 9 1 11 2 12 9 13 1 9 2 3 12 9 1 9 1 9 0 1 10 9 2 13 9 0 1 9 2
10 9 1 9 1 9 1 10 9 0 2
20 4 13 1 10 9 2 10 9 1 10 9 15 4 4 3 13 1 10 9 2
15 15 13 10 9 3 0 1 10 9 11 7 10 9 0 2
16 12 12 13 1 11 3 4 4 13 1 10 9 2 0 2 2
46 13 3 12 12 10 9 15 4 3 13 1 10 9 1 11 2 1 15 15 13 10 9 1 9 7 9 1 9 1 10 11 2 10 9 0 15 1 10 9 1 11 4 13 12 9 2
31 10 0 9 2 16 4 4 13 10 9 1 9 2 10 9 15 4 13 1 9 7 4 13 10 9 1 9 1 10 9 2
21 13 3 10 11 1 13 10 2 9 0 2 2 16 7 16 10 9 13 1 11 2
31 10 10 9 13 15 1 13 9 1 9 1 13 10 9 1 10 9 2 15 1 10 9 15 4 13 10 9 1 10 9 2
29 10 9 2 11 2 3 3 13 10 9 0 7 4 13 15 1 10 9 1 9 1 9 0 3 0 1 10 11 2
46 1 10 9 0 15 13 1 10 9 0 2 10 11 4 2 13 2 1 10 0 9 1 10 12 12 1 10 12 12 9 1 9 2 9 1 9 0 7 0 3 3 0 7 3 0 2
75 13 0 16 1 10 9 1 11 15 13 10 9 1 10 9 2 9 13 1 10 0 9 0 7 2 9 2 2 7 10 9 2 3 15 13 3 1 10 9 1 10 2 9 2 2 13 0 1 10 9 7 13 3 1 10 9 0 1 9 10 10 9 3 13 1 10 9 13 1 10 9 1 10 9 2
8 1 15 13 9 3 13 0 2
25 1 11 13 16 10 0 9 0 2 9 1 9 1 10 9 1 10 10 11 2 3 4 13 3 2
40 1 10 9 2 3 2 15 13 10 9 7 10 9 13 9 2 3 16 1 9 2 1 10 9 0 0 2 3 0 2 15 13 9 1 10 9 3 1 13 2
20 1 10 9 1 10 9 10 9 0 1 11 13 3 10 9 1 13 10 9 2
8 10 9 4 13 1 10 9 2
50 10 9 1 10 9 1 11 4 13 1 10 9 1 9 0 1 10 9 0 2 16 13 10 9 16 1 10 9 13 11 11 7 10 9 1 13 10 9 1 10 9 0 15 13 3 1 10 9 0 2
10 10 9 0 1 11 13 10 0 9 2
16 15 4 13 3 13 15 9 2 9 1 10 9 0 2 9 2
27 1 10 10 0 9 2 3 0 2 10 9 1 10 9 4 13 1 10 0 12 9 10 2 0 9 2 2
38 10 9 3 10 9 1 10 9 3 13 10 12 9 1 10 9 2 10 9 1 10 9 0 4 13 1 12 9 2 10 11 13 1 10 12 1 12 2
34 1 10 12 2 16 10 11 13 10 9 1 9 1 10 9 2 4 13 3 12 9 0 2 1 9 0 15 13 10 12 9 1 9 2
21 1 10 9 15 13 1 0 9 1 10 9 0 2 0 2 0 2 0 2 0 2
75 1 10 9 3 0 1 10 9 1 9 0 2 15 1 10 9 0 11 11 2 15 4 13 1 11 10 9 1 10 9 1 10 11 2 4 13 1 12 9 0 9 1 12 9 1 9 2 7 1 10 9 0 11 2 15 4 13 1 11 10 0 9 1 10 9 1 9 1 9 13 12 9 1 9 2
36 7 13 3 0 10 9 13 1 10 0 9 0 1 0 9 2 15 13 10 9 1 10 9 0 1 10 9 1 11 2 1 10 9 1 11 2
28 10 11 2 1 12 9 1 9 1 9 7 12 1 9 1 10 12 2 13 3 10 0 9 0 1 10 11 2
20 10 9 1 9 13 1 10 9 1 9 15 13 11 1 11 2 11 7 11 2
27 1 15 3 2 1 10 10 9 0 15 15 4 13 1 10 9 1 10 9 0 2 10 9 4 13 0 2
8 9 0 7 0 1 0 9 2
8 9 1 10 9 15 1 13 2
12 0 9 1 9 0 2 0 2 0 7 0 2
6 9 1 9 0 0 2
12 15 10 0 9 15 4 4 13 10 9 0 2
57 1 13 10 9 3 0 2 10 9 1 10 9 0 7 10 13 9 15 3 1 12 9 13 10 9 0 15 3 4 13 10 10 9 1 13 1 10 11 1 10 9 7 15 3 1 9 15 15 13 3 1 10 10 9 1 11 2
27 15 4 13 1 10 9 0 2 4 13 10 9 1 10 9 15 4 13 1 10 9 7 4 13 1 11 2
25 7 15 4 13 0 1 10 9 0 2 3 13 0 1 13 15 1 9 1 10 9 1 10 9 2
33 1 11 11 2 9 1 10 9 1 10 9 0 1 11 10 9 13 9 1 10 9 0 7 13 16 10 9 13 0 2 1 15 2
41 4 13 1 10 9 1 9 10 12 9 1 9 15 2 1 10 9 2 9 13 3 12 9 7 13 1 9 0 2 4 13 1 9 1 10 9 1 11 12 9 2
8 12 9 7 12 1 9 0 2
32 10 9 4 3 13 10 9 11 15 15 13 2 1 9 1 0 9 2 1 10 9 1 10 9 0 1 1 9 10 0 9 2
13 12 11 1 10 9 0 0 13 7 13 9 0 2
16 7 4 13 12 10 9 3 0 1 11 1 10 9 1 11 2
58 10 9 13 1 10 9 1 9 1 10 11 15 13 1 12 2 12 2 10 9 1 10 10 9 15 3 15 13 1 10 2 9 1 10 9 2 2 13 3 10 0 9 0 1 10 12 9 7 9 0 15 13 10 9 1 10 11 2
37 10 9 13 3 15 0 1 11 2 11 7 11 2 3 15 13 3 13 0 9 2 3 16 13 0 10 9 1 10 11 1 3 13 15 1 11 2
8 10 9 1 9 1 9 0 2
56 15 13 16 2 1 10 0 9 1 10 9 0 2 10 0 9 4 1 0 9 13 10 9 0 1 9 2 7 1 15 13 10 9 1 10 9 0 1 10 9 7 1 10 9 0 13 1 10 9 1 10 2 9 2 0 2
45 13 0 2 1 10 11 2 16 1 10 9 1 10 9 0 2 1 10 9 3 0 2 10 0 9 13 1 10 9 0 2 9 7 9 2 1 10 9 1 9 1 13 10 9 2
58 1 10 9 1 10 9 0 15 15 13 16 4 3 13 1 9 1 10 9 0 2 10 9 1 10 9 0 0 7 1 10 9 0 1 10 9 1 9 1 10 9 0 1 0 7 0 9 15 13 1 10 9 0 0 1 10 9 2
52 3 1 9 1 10 9 3 13 9 2 10 9 11 11 4 13 13 10 9 1 10 9 1 10 9 11 11 11 2 1 9 1 10 9 15 10 11 4 13 1 10 13 10 9 0 1 13 9 1 10 9 2
72 3 4 4 13 9 1 10 10 9 1 11 1 10 9 1 10 9 1 9 11 2 1 15 4 4 13 10 9 3 1 9 1 9 2 7 1 10 9 0 0 2 11 0 0 7 11 0 2 10 10 9 0 0 3 1 10 11 2 11 2 15 4 13 1 10 9 0 3 1 11 2 2
58 1 10 9 1 10 9 1 9 1 10 11 2 9 1 10 9 7 10 9 1 11 2 2 10 9 1 10 9 0 11 11 11 2 11 4 13 16 10 11 13 10 9 1 13 1 11 2 3 1 10 9 1 10 9 1 10 9 2
38 11 3 13 13 10 9 1 11 1 10 0 2 9 3 3 10 0 9 15 4 13 7 4 13 1 4 13 1 10 9 0 7 1 10 9 0 0 2
13 10 9 1 9 0 15 11 4 13 1 0 9 2
26 10 9 1 9 1 10 9 11 11 4 13 3 1 9 15 15 10 9 13 10 9 1 2 9 2 2
37 1 9 15 4 13 1 10 0 2 9 0 2 0 7 0 2 13 1 10 0 0 9 1 10 9 7 1 9 3 0 7 1 9 1 10 9 2
25 1 15 1 10 9 1 0 7 0 9 2 16 1 10 9 15 4 13 2 15 13 10 0 9 2
36 10 9 1 10 10 9 1 9 1 15 3 3 15 13 10 9 1 9 7 10 9 1 9 1 9 0 13 1 10 9 2 9 1 10 9 2
27 10 9 1 9 3 13 9 1 10 9 1 10 0 9 0 2 7 1 10 0 9 1 10 9 1 9 2
14 10 9 3 13 3 0 2 7 10 9 4 3 13 2
36 10 11 13 1 10 9 0 10 9 0 2 9 1 9 1 9 7 1 10 0 9 1 9 1 10 9 13 1 9 1 10 9 1 11 11 2
27 10 9 1 9 4 13 0 7 13 3 0 2 13 3 3 0 1 10 0 9 1 9 0 7 9 0 2
28 10 9 0 1 11 11 2 3 3 0 1 10 9 0 2 7 1 15 0 1 9 2 4 13 10 9 0 2
46 10 9 0 1 10 12 9 12 4 4 13 1 10 9 3 0 1 9 2 9 7 9 2 1 13 10 9 0 1 10 11 2 15 3 4 3 13 1 13 10 9 1 10 9 0 2
45 15 0 2 13 15 10 0 9 1 9 2 4 4 13 1 10 0 9 1 9 2 1 15 10 9 2 7 15 4 13 3 3 2 3 1 13 13 1 10 9 0 1 10 9 2
14 10 9 0 1 10 0 9 4 3 13 13 10 9 2
14 10 11 13 3 10 9 1 10 0 7 0 9 0 2
53 10 9 1 10 9 0 13 1 10 9 1 9 1 13 10 9 1 9 2 7 3 1 13 10 9 0 7 1 13 1 9 1 10 9 10 9 1 10 9 0 2 11 11 2 3 4 3 13 1 13 10 9 2
6 10 9 0 13 0 2
17 10 11 13 3 3 3 2 1 10 9 0 1 10 10 9 0 2
30 13 3 0 16 2 3 1 10 9 2 15 13 1 10 9 1 10 0 9 7 1 10 9 1 9 1 10 0 9 2
14 10 9 13 0 2 7 4 13 3 0 16 15 13 2
53 10 9 1 10 11 1 13 10 10 9 0 1 10 11 13 1 10 15 0 7 0 2 7 13 1 13 1 9 10 9 1 10 9 1 10 12 9 15 4 4 3 13 1 10 9 1 10 9 1 10 11 11 2
32 10 9 1 11 4 3 13 15 1 10 9 0 1 10 11 2 13 1 10 9 1 9 2 7 3 1 10 9 0 1 11 2
8 10 0 0 9 1 9 0 2
30 10 0 9 1 13 1 10 9 13 13 15 1 13 0 9 0 2 1 13 15 2 10 9 2 1 10 0 9 0 2
36 7 10 0 1 4 15 15 13 4 13 10 0 9 2 1 13 1 10 9 13 10 0 9 7 3 3 3 0 2 3 1 10 9 0 2 2
16 3 1 10 9 13 3 3 0 13 1 0 9 1 9 0 2
39 16 3 10 9 4 13 7 13 15 1 0 7 0 9 0 2 3 3 15 13 10 9 1 10 9 2 16 3 15 1 13 9 0 1 10 0 9 0 2
17 10 9 1 10 0 12 9 13 1 13 1 9 10 9 1 9 2
27 1 10 9 1 10 9 2 10 9 1 11 4 13 0 9 1 10 11 2 13 15 10 9 1 10 9 2
11 3 1 10 0 12 2 11 11 4 13 2
47 7 1 10 11 0 2 3 4 13 10 9 0 2 1 10 12 4 13 10 2 9 0 2 10 10 9 4 13 1 10 9 11 11 1 10 9 1 10 9 2 10 11 1 10 9 2 2
29 13 10 0 9 0 2 10 9 0 13 10 9 1 10 9 7 10 15 13 2 1 13 1 10 12 2 15 0 2
58 1 10 12 2 1 10 9 1 11 2 10 9 11 13 10 9 1 10 11 1 10 9 1 10 11 2 7 10 9 0 2 0 1 10 9 12 2 15 13 10 9 1 11 2 4 13 3 1 10 9 7 11 13 1 10 9 0 2
45 10 0 9 13 16 10 11 15 13 1 10 9 7 10 9 0 4 13 10 9 1 10 11 1 10 9 1 10 9 2 15 13 10 12 9 12 3 1 10 9 1 10 10 9 2
18 1 10 12 10 0 11 11 13 10 9 7 12 9 3 4 13 9 2
29 1 10 9 1 9 1 10 11 13 10 10 9 1 10 11 1 15 13 10 12 9 12 10 9 1 9 7 9 2
43 10 9 2 3 2 4 13 10 9 1 9 1 10 9 1 10 9 0 1 10 0 9 1 10 9 1 9 2 1 10 0 9 1 10 9 0 1 10 9 1 11 0 2
18 3 4 13 1 10 10 9 2 4 13 11 2 7 1 10 9 13 2
40 1 13 0 9 4 4 3 13 1 10 9 10 9 1 9 1 10 9 0 2 15 4 13 10 9 1 9 7 10 9 0 1 11 3 13 3 1 0 9 2
9 1 10 9 13 10 9 3 0 2
28 1 10 9 15 13 10 9 1 11 7 1 10 9 2 1 10 15 15 13 1 13 10 9 1 9 7 9 2
30 10 0 9 15 4 13 10 0 9 1 10 9 2 15 3 3 15 13 1 9 2 7 3 15 15 13 3 10 0 2
26 1 10 2 9 2 0 7 1 10 9 15 4 13 10 9 7 10 9 1 10 9 13 3 0 9 2
9 15 2 3 2 13 3 9 0 2
14 1 9 10 9 1 10 9 0 1 9 2 11 11 2
35 1 10 0 9 2 12 9 3 2 4 13 13 1 10 10 9 9 1 12 12 9 2 10 9 13 1 9 9 15 15 4 13 3 13 2
27 3 15 1 15 15 4 13 1 10 9 4 13 10 9 1 10 9 7 13 1 13 10 10 9 1 15 2
44 10 9 0 1 10 11 11 2 15 3 4 13 10 9 2 13 16 2 3 1 10 9 1 15 13 1 13 9 0 1 10 9 1 10 9 11 2 4 13 10 9 1 9 2
6 7 15 13 10 15 2
19 1 11 13 1 15 1 13 16 10 2 9 2 3 4 13 1 10 9 2
3 10 9 2
37 11 2 11 2 11 2 15 1 9 3 3 13 1 10 9 0 16 15 2 3 13 13 7 1 10 9 13 2 4 13 3 10 9 1 0 9 2
29 15 3 13 10 9 13 10 9 11 11 15 1 10 9 11 4 13 9 1 13 10 10 9 1 10 9 1 9 2
9 11 13 3 3 10 0 9 0 2
21 10 9 1 10 9 0 2 9 1 10 9 1 9 2 1 10 9 0 1 9 2
18 7 3 13 10 9 10 9 7 10 9 1 13 1 9 10 10 9 2
13 0 2 13 11 2 4 13 9 1 9 1 9 2
25 7 3 13 0 16 13 3 10 15 1 15 4 4 13 1 10 9 2 10 10 9 13 10 9 2
28 16 10 9 4 13 2 3 10 9 1 10 9 0 7 1 10 9 0 4 13 1 9 10 10 9 1 9 2
16 16 15 13 1 11 2 3 2 13 10 10 9 1 9 0 2
18 13 0 1 10 15 15 13 9 7 9 0 2 1 13 15 1 3 2
30 7 10 9 1 10 9 7 1 10 9 13 1 10 9 1 9 1 13 10 9 15 13 10 9 0 3 0 1 11 2
57 16 10 9 15 4 13 1 9 1 13 3 1 10 9 1 10 9 1 15 1 10 2 9 2 2 13 9 16 10 9 4 13 10 9 13 1 9 7 11 0 1 13 10 12 0 9 7 10 9 1 9 13 1 9 1 9 2
31 10 9 1 10 9 4 3 13 1 9 3 3 10 9 1 10 9 7 3 10 9 1 10 9 1 11 1 10 9 0 2
19 10 9 2 4 13 2 4 4 13 1 9 7 9 1 10 13 9 0 2
15 1 10 10 9 1 9 10 9 4 13 13 3 9 0 2
37 1 10 9 1 11 4 4 13 12 9 2 15 12 1 10 9 1 11 2 10 2 9 2 1 15 4 13 15 1 10 3 0 9 1 9 0 2
23 1 10 9 4 13 10 9 1 10 9 2 1 15 3 10 9 1 10 9 0 1 11 2
65 16 1 9 9 0 7 9 0 13 10 9 1 10 2 9 2 0 1 11 2 13 1 9 10 9 1 10 9 15 13 1 0 9 7 3 1 9 1 10 9 9 1 9 1 9 2 10 0 9 15 13 10 9 1 10 9 0 2 13 15 1 10 9 13 2
45 1 11 10 9 1 10 9 2 15 13 10 9 1 2 11 2 4 13 10 9 7 10 9 1 10 9 7 10 9 1 9 1 9 3 4 13 2 3 2 1 13 9 0 0 2
30 13 1 9 1 10 9 1 10 9 0 2 4 13 1 13 1 9 10 9 15 13 9 1 10 12 5 1 10 9 2
8 3 1 10 9 1 0 9 2
10 16 10 9 15 13 2 13 10 9 2
31 11 4 13 1 13 15 1 8 8 1 13 2 0 7 0 9 0 1 10 15 4 13 1 9 2 1 10 13 2 9 2
18 3 12 12 9 2 1 15 3 9 2 9 7 9 2 15 4 13 2
19 3 10 9 3 4 13 3 10 9 15 15 4 13 3 12 9 1 9 2
11 3 1 10 11 13 10 9 1 10 9 2
28 13 1 10 9 2 4 13 3 10 9 1 9 3 11 2 7 10 9 4 13 1 11 10 9 1 10 9 2
47 10 2 9 2 13 1 11 11 13 10 9 1 9 16 13 1 13 1 10 9 1 9 10 9 11 2 15 1 10 10 2 9 0 2 15 1 10 9 1 10 9 4 13 10 9 0 2
82 10 9 1 10 9 0 0 2 13 1 9 1 9 2 13 10 9 1 9 1 10 9 3 0 1 11 7 13 1 13 10 0 9 1 10 9 1 10 0 9 11 11 7 1 10 9 2 1 10 9 3 13 1 10 9 0 2 1 10 9 11 11 2 13 1 10 9 0 1 3 4 13 1 9 1 13 10 9 1 10 9 2
46 10 9 0 15 3 13 1 9 13 15 1 10 9 7 13 1 9 10 9 1 9 7 1 10 9 1 10 9 0 2 3 13 1 13 3 1 11 7 1 11 10 9 1 10 9 2
32 10 9 1 11 2 13 3 1 10 9 0 2 7 1 10 0 9 2 4 3 13 1 3 10 0 9 1 11 1 10 9 2
34 1 11 7 11 13 1 10 0 9 2 1 11 1 10 9 1 9 2 15 1 10 15 13 1 10 9 1 10 11 1 10 9 0 2
9 7 10 9 3 4 13 1 9 2
34 3 3 1 10 9 13 0 9 1 13 9 2 1 9 11 11 1 10 9 12 13 10 9 9 1 10 11 0 1 10 9 1 11 2
24 15 1 10 0 9 13 1 10 9 7 2 1 10 9 2 1 10 9 2 10 0 9 0 2
17 1 9 2 4 4 13 10 9 0 2 13 10 9 1 10 9 2
35 3 10 9 1 9 3 2 16 3 10 9 1 9 0 13 1 13 10 9 2 10 9 2 10 9 0 2 4 13 10 9 1 10 9 2
37 10 9 2 3 13 1 10 9 1 9 2 13 1 13 1 11 9 0 7 13 9 1 9 0 3 1 13 1 10 9 1 10 2 9 0 2 2
25 3 2 10 9 4 13 10 0 9 1 13 9 2 9 2 9 2 15 15 13 1 13 10 9 2
16 10 9 1 10 9 0 1 11 13 3 10 0 9 1 9 2
41 10 9 1 11 7 0 9 0 4 13 1 10 9 1 10 2 9 1 10 9 2 2 10 9 15 3 13 3 10 9 7 3 10 0 9 13 1 10 9 0 2
53 10 9 2 1 10 15 4 13 3 10 12 5 1 10 9 0 2 13 1 10 9 7 3 11 2 15 10 9 13 10 9 0 2 4 13 1 13 10 9 16 10 9 0 4 3 13 1 10 9 1 10 9 2
20 3 1 10 9 13 10 9 2 1 15 10 11 4 13 10 3 0 9 0 2
17 1 12 9 1 10 9 13 3 1 3 10 9 0 1 10 9 2
9 10 9 0 4 13 10 9 0 2
65 13 10 9 1 10 9 1 10 9 7 10 9 1 11 2 3 10 9 0 4 13 10 9 1 10 9 1 10 9 1 9 1 12 1 10 12 9 15 4 4 13 1 10 9 1 10 9 1 9 11 1 10 0 9 1 10 9 3 13 1 10 9 1 11 2
33 10 9 0 4 3 13 1 10 9 0 10 9 1 10 9 0 15 4 13 1 10 9 0 10 9 1 11 1 10 9 1 11 2
11 7 3 10 9 1 10 9 13 10 9 2
53 1 9 1 9 2 9 9 10 9 0 0 4 13 10 9 1 10 9 1 9 1 13 16 15 13 1 10 9 15 1 12 9 4 13 10 9 1 10 9 1 10 9 0 1 10 11 11 2 10 9 1 11 2
5 10 9 10 9 2
22 10 9 0 3 4 3 13 1 9 1 10 0 9 1 10 12 7 1 10 12 9 2
18 10 9 0 11 3 13 16 11 13 3 0 1 13 10 9 1 9 2
10 7 1 10 11 13 3 10 0 9 2
73 1 10 11 3 3 15 13 1 9 1 11 7 1 10 0 2 9 0 7 0 2 7 3 1 13 1 10 9 10 9 1 10 0 2 10 9 2 9 7 10 9 0 2 0 1 10 9 1 10 0 2 3 0 16 10 9 13 3 10 9 0 1 13 9 7 9 1 10 9 0 7 0 2
19 0 9 13 1 10 9 13 1 11 2 15 3 9 4 4 13 1 9 2
14 16 4 13 13 10 9 2 10 9 4 13 10 9 2
9 9 15 13 3 1 10 0 9 2
58 1 10 9 0 1 11 2 1 11 2 1 11 2 3 3 9 1 10 9 4 13 10 9 1 9 2 2 11 2 11 2 11 2 1 10 9 1 10 9 4 13 10 9 1 10 9 0 2 11 11 2 15 4 13 10 9 2 2
28 1 9 1 9 2 10 9 0 9 4 13 2 3 1 0 9 2 10 9 2 15 1 11 15 13 10 9 2
25 10 9 0 1 11 4 13 10 9 11 1 13 15 1 0 9 1 10 9 7 1 13 10 9 2
35 10 9 1 9 2 15 4 13 1 12 0 9 0 13 9 0 2 4 13 16 3 4 4 3 13 9 0 1 13 10 9 1 10 9 2
71 13 15 1 10 3 0 9 1 10 10 9 1 16 4 13 10 0 9 1 10 12 2 10 9 1 11 11 4 13 1 13 10 9 1 10 9 2 15 13 1 13 10 9 1 10 0 9 2 13 10 9 1 9 1 9 2 13 9 0 3 1 12 9 1 10 9 7 13 10 9 2
43 1 15 1 10 9 1 10 9 4 13 10 9 2 7 10 9 4 13 10 0 1 10 9 1 10 9 1 10 9 1 4 15 13 2 16 3 9 2 1 10 9 9 2
32 7 3 10 9 1 10 9 1 10 9 4 13 13 1 10 9 10 9 2 13 16 10 9 13 1 3 13 3 10 10 9 2
19 10 9 1 9 2 13 11 11 2 9 1 11 1 10 9 0 0 2 2
23 15 13 10 10 9 2 1 9 2 1 10 9 13 1 10 9 15 13 10 11 9 0 2
38 13 10 0 2 0 11 11 1 13 1 10 11 1 11 11 10 9 0 15 1 10 11 0 1 10 9 12 4 13 2 3 13 2 10 9 1 9 2
7 15 13 10 2 11 2 2
53 15 2 13 2 10 9 7 15 15 13 1 9 10 15 2 10 0 13 13 3 10 0 9 1 13 1 10 8 8 1 10 2 9 2 0 2 3 1 16 10 3 0 13 3 1 9 2 7 15 13 10 9 2
26 1 10 9 12 11 13 9 1 9 1 10 9 15 13 1 10 0 9 1 10 9 1 10 0 9 2
10 10 0 13 2 3 2 1 10 0 2
30 15 1 0 2 1 9 2 1 10 9 1 10 2 9 1 10 9 2 2 7 10 9 1 10 9 10 9 13 0 2
22 13 10 9 1 9 13 10 9 0 7 10 12 9 1 10 9 1 10 9 1 9 2
37 10 9 1 10 9 1 10 11 11 4 4 13 1 9 7 9 1 9 15 4 13 1 11 2 11 2 11 7 11 12 9 1 9 0 1 9 2
29 1 10 9 13 9 7 9 0 2 9 1 9 2 9 7 9 1 9 7 9 1 9 1 10 9 1 10 9 2
33 10 9 13 1 10 9 1 13 13 1 10 9 0 13 7 13 1 10 11 2 9 7 9 1 9 0 13 1 0 9 7 9 2
27 10 9 0 1 10 9 1 10 11 11 13 3 1 10 9 2 1 10 9 2 13 1 12 9 1 9 2
30 10 9 2 1 10 9 2 13 10 9 0 1 10 9 7 1 10 9 1 10 9 1 15 4 13 7 13 10 9 2
12 9 7 9 1 9 4 3 13 10 9 0 2
8 15 13 10 9 1 10 9 2
24 1 9 2 3 1 10 9 1 10 9 2 10 9 13 1 10 9 1 10 9 10 10 9 2
37 2 1 15 2 13 10 9 1 10 9 2 11 11 2 10 9 4 13 1 10 9 1 10 9 3 0 2 13 1 10 9 1 10 9 13 2 2
31 11 4 13 10 9 0 1 10 11 1 10 10 9 2 7 3 4 13 10 9 1 10 9 13 1 10 9 1 10 9 2
23 1 3 10 9 1 2 10 9 3 0 7 0 16 4 13 10 9 1 10 9 0 2 2
40 3 10 11 2 1 10 9 1 10 11 2 11 11 2 13 10 9 2 16 3 4 13 3 10 11 1 13 10 9 0 2 0 2 0 1 10 10 9 2 2
30 1 10 9 10 9 1 9 4 3 13 0 2 1 10 9 15 13 15 13 10 9 3 1 10 12 2 12 9 2 2
17 1 10 9 10 9 1 10 9 9 2 13 10 9 13 1 11 2
13 10 9 1 10 11 2 3 2 4 13 1 13 2
19 7 13 0 16 13 3 10 9 1 13 10 9 1 10 9 1 10 9 2
26 10 0 9 13 1 13 10 9 1 9 1 10 0 12 1 12 1 10 0 9 1 10 12 1 12 2
37 10 13 2 1 10 9 1 10 9 2 4 13 1 13 2 3 1 10 9 0 2 10 9 1 0 9 2 0 7 0 2 2 13 1 10 9 2
35 10 9 0 4 13 3 1 13 10 9 15 1 10 0 9 1 10 12 13 10 9 0 1 10 9 1 9 1 10 0 12 9 1 12 2
29 13 10 9 15 3 2 1 12 1 3 2 13 10 9 7 1 10 9 10 12 2 7 1 10 9 10 12 9 2
23 3 1 10 12 3 13 9 7 15 13 10 9 1 15 13 1 13 1 10 9 10 9 2
15 10 9 11 13 1 10 9 1 11 2 9 1 10 12 2
19 10 0 11 2 10 0 9 1 13 10 9 1 11 2 13 3 1 11 2
14 7 3 15 13 3 10 9 1 9 0 2 1 11 2
21 10 9 0 1 10 0 9 13 1 11 10 9 0 1 10 12 5 1 10 9 2
14 13 3 10 3 9 1 9 1 10 9 1 10 9 2
17 0 13 10 12 5 13 1 10 9 0 1 10 11 2 11 11 2
29 0 2 13 10 9 1 10 9 2 11 15 4 3 13 1 10 9 1 4 13 13 2 10 0 9 2 1 11 2
14 4 3 13 9 13 3 1 15 1 10 10 9 0 2
23 1 10 9 11 2 10 10 9 1 10 12 4 1 0 9 13 9 2 9 7 0 9 2
18 15 2 10 9 2 1 3 15 4 3 13 1 10 13 9 1 9 2
14 10 10 9 11 4 3 9 0 1 10 11 1 11 2
12 15 4 13 10 9 1 10 9 1 10 9 2
37 11 2 15 3 9 4 3 13 1 11 1 13 15 2 2 15 4 13 7 15 4 13 10 10 9 1 10 0 9 2 2 4 13 10 0 9 2
37 13 1 3 12 9 7 12 9 10 0 9 1 10 9 1 10 12 9 0 13 3 1 10 9 1 11 2 11 7 11 2 13 1 10 9 0 2
30 10 0 9 4 13 1 9 10 9 1 9 1 11 2 12 9 1 9 1 11 2 13 12 9 7 13 15 0 12 2
29 10 0 9 15 4 13 13 1 10 9 1 10 9 1 11 2 1 11 2 13 3 12 9 7 13 15 0 12 2
38 10 9 4 13 3 1 10 12 2 9 0 2 1 3 1 12 9 1 10 9 0 2 10 9 13 1 10 9 3 15 13 10 9 0 7 10 9 2
12 10 0 9 1 10 9 1 10 9 1 11 2
28 10 9 13 1 9 4 4 13 1 10 9 13 1 9 1 10 9 0 2 1 10 9 0 1 10 0 9 2
21 10 9 13 1 3 10 9 7 12 9 2 10 9 4 4 13 1 10 9 0 2
40 15 4 13 9 1 10 13 10 9 1 10 12 2 12 1 10 9 1 13 1 10 9 1 9 3 10 9 1 11 2 15 4 13 10 9 13 10 9 0 2
30 13 10 9 1 9 1 10 0 9 13 1 9 2 16 15 13 10 9 1 13 10 9 7 16 3 15 15 13 3 2
9 11 3 13 3 10 9 1 9 2
8 3 15 4 13 10 0 9 2
10 10 9 1 10 9 3 15 13 3 2
43 10 11 15 13 3 10 9 1 3 4 13 10 9 1 10 9 3 0 2 1 11 11 2 7 4 13 1 9 1 10 9 1 3 13 1 9 3 1 10 0 12 9 2
9 10 9 15 4 13 15 1 9 2
15 1 10 15 2 1 10 12 2 11 15 4 13 10 9 2
47 7 4 13 10 9 1 10 9 1 13 7 3 2 10 9 3 2 3 1 10 9 1 9 1 11 2 11 13 1 9 2 11 3 1 10 9 13 7 11 13 10 9 1 10 9 0 2
20 10 11 1 10 12 9 0 15 4 13 1 13 0 10 9 1 10 0 9 2
23 7 15 13 10 9 13 1 10 9 2 15 1 16 13 1 10 9 0 1 10 9 0 2
47 16 10 11 1 9 1 13 15 2 3 1 10 9 13 7 1 11 13 1 10 0 9 0 2 16 3 13 3 2 13 10 9 1 10 0 1 10 9 13 10 9 1 10 9 0 0 2
25 10 9 13 10 9 1 16 10 0 9 10 9 13 0 2 3 13 1 11 7 1 10 9 11 2
35 16 11 13 10 9 1 10 9 0 7 0 1 11 13 10 9 1 13 1 9 1 11 2 0 9 1 10 9 2 15 13 10 9 0 2
14 10 9 13 1 10 0 9 1 10 9 0 7 0 2
13 10 9 1 10 9 1 11 1 2 11 11 2 2
25 13 9 10 0 9 1 10 9 1 10 9 15 15 13 1 10 11 1 10 12 1 10 12 9 2
17 13 10 9 10 2 9 12 2 2 9 13 3 1 10 9 0 2
17 10 2 11 2 2 7 10 9 13 1 10 9 1 10 9 0 2
30 16 4 13 11 11 2 11 11 2 2 2 13 9 13 1 15 1 12 9 2 15 3 4 4 13 0 1 11 2 2
11 3 10 9 12 13 10 9 1 10 9 2
27 13 2 11 7 9 2 2 15 13 3 2 1 9 1 9 2 2 1 13 10 9 2 2 4 13 11 2
18 10 9 1 10 9 2 0 2 13 1 9 1 10 12 9 1 11 2
31 1 13 2 7 3 13 2 10 9 1 10 9 2 4 13 10 9 2 7 13 3 0 9 1 9 2 3 1 11 2 2
16 10 9 13 10 9 12 2 12 7 12 2 15 1 11 11 2
41 10 12 4 13 10 0 9 1 10 9 1 10 9 11 2 3 15 13 10 9 1 10 9 2 1 9 3 1 10 9 11 2 1 10 11 7 1 10 11 11 2
13 10 9 13 3 10 9 3 0 1 10 0 9 2
37 1 9 1 9 4 13 10 9 1 9 2 4 13 16 11 4 13 10 9 0 2 4 13 3 11 1 10 15 7 1 10 10 9 15 4 13 2
13 0 9 2 13 10 0 9 1 10 10 12 9 2
19 10 0 9 7 4 13 1 9 2 4 13 1 11 10 9 1 0 9 2
24 11 13 3 2 3 16 11 13 1 13 15 10 9 1 10 9 1 10 9 1 3 13 3 2
33 10 11 13 2 11 13 10 11 1 9 1 9 0 2 11 13 0 1 10 11 1 10 9 2 15 10 9 13 1 9 1 9 2
11 12 9 10 9 1 10 12 1 10 11 2
6 10 9 13 10 9 2
12 10 9 2 3 2 13 1 11 1 13 11 2
12 4 13 10 9 7 15 13 3 1 10 9 2
12 13 10 9 1 10 9 2 10 9 15 13 2
19 10 0 9 13 15 1 13 1 0 9 11 2 15 3 4 13 10 9 2
43 13 10 9 1 10 9 12 2 10 9 1 10 9 13 1 0 9 7 15 13 3 1 10 9 2 9 1 9 2 10 9 3 3 15 13 1 10 9 0 1 11 2 2
21 2 10 9 15 4 13 3 10 9 7 13 1 11 3 1 9 1 10 9 2 2
39 9 11 3 13 0 2 3 13 3 1 9 2 3 13 1 10 9 1 10 9 1 10 11 7 3 1 13 10 9 1 9 15 4 13 10 9 3 0 2
6 15 13 9 1 13 2
15 10 9 12 13 10 9 1 9 3 1 13 15 1 11 2
16 9 0 2 16 1 9 10 9 13 10 0 9 1 11 11 2
8 15 13 10 12 9 1 11 2
21 11 7 11 2 1 10 9 2 13 10 9 1 10 9 7 1 9 1 10 9 2
19 3 9 1 10 9 0 1 11 2 3 7 9 9 0 7 9 1 11 2
48 15 13 3 1 10 9 2 13 10 9 2 10 9 1 10 0 9 2 10 0 9 1 10 2 9 1 9 2 2 0 9 1 10 0 13 1 10 11 2 10 9 1 10 0 9 1 11 2
36 10 9 1 10 9 0 13 10 9 1 9 15 13 10 9 1 10 12 2 7 15 13 3 1 10 9 2 10 9 13 1 10 11 1 9 2
10 13 10 9 1 10 11 2 11 11 2
24 1 10 12 2 13 1 10 9 1 2 10 9 0 2 11 11 2 13 10 9 1 10 9 2
30 11 11 11 11 2 0 9 1 10 9 9 1 10 11 1 10 9 2 13 1 10 9 0 1 9 1 10 9 0 2
42 10 9 1 10 0 4 13 1 11 11 2 1 15 13 10 9 1 9 1 10 9 2 7 1 11 11 2 9 9 1 10 11 2 1 10 9 1 9 1 10 9 2
23 1 3 10 9 13 1 10 9 7 2 1 9 2 10 9 13 10 9 0 1 10 9 2
32 10 9 13 10 9 1 10 9 0 1 9 2 10 9 1 10 9 2 3 15 15 15 13 1 13 10 9 1 9 1 9 2
27 4 13 1 9 1 13 16 2 1 10 0 9 1 15 15 13 2 13 0 1 9 1 9 0 1 9 2
17 10 9 1 10 9 0 13 12 1 9 0 7 9 1 10 9 2
27 1 9 7 9 4 13 1 11 10 9 2 10 0 9 13 12 12 2 2 1 9 1 10 9 7 3 2
38 10 9 0 1 10 9 13 10 9 13 1 10 0 2 3 15 4 13 10 9 1 10 10 9 2 9 2 9 2 9 2 9 2 9 7 9 0 2
15 10 9 13 11 11 13 1 13 15 1 10 9 13 9 2
21 13 3 10 9 11 1 10 9 1 11 1 10 9 1 10 9 1 10 9 11 2
28 1 13 15 15 13 9 3 1 0 9 2 16 10 9 4 13 0 1 15 15 13 3 1 3 13 10 9 2
46 10 9 15 13 1 13 10 9 1 10 9 4 13 2 3 16 1 10 0 9 1 10 9 1 11 2 3 1 10 9 9 2 13 1 9 1 9 1 10 9 0 1 10 9 0 2
18 10 2 9 1 9 2 4 13 1 10 0 9 1 10 11 1 11 2
15 3 15 13 3 10 9 2 3 15 15 13 3 10 9 2
27 3 11 11 2 9 1 10 9 13 2 10 9 4 13 1 9 10 9 7 4 13 10 9 1 10 9 2
25 10 0 9 2 12 1 9 1 10 9 2 4 3 13 1 9 10 9 1 11 7 1 11 11 2
38 7 1 10 0 9 1 10 9 0 2 3 10 9 1 10 9 4 4 13 1 9 1 10 9 7 4 13 10 9 1 10 9 2 10 9 11 11 2
27 7 10 9 10 9 1 10 9 1 10 9 4 13 9 1 10 9 0 1 10 9 1 11 7 1 11 2
33 1 9 11 2 1 10 9 1 9 7 9 2 4 13 3 3 12 9 0 1 3 15 1 12 9 1 9 2 1 9 1 9 2
16 11 11 2 15 15 13 1 9 1 9 0 2 3 13 9 2
19 2 11 15 1 10 0 9 2 10 9 15 4 13 10 9 1 9 2 2
11 1 10 9 2 11 11 13 1 13 0 2
22 2 15 4 13 16 4 13 1 10 9 1 10 11 7 10 9 4 13 10 9 2 2
22 1 3 16 15 3 15 4 13 10 9 1 13 9 0 2 15 15 15 13 3 0 2
22 2 4 13 9 3 1 9 1 13 3 10 9 1 10 9 2 2 13 3 10 9 2
15 10 9 13 10 9 0 7 0 2 7 3 15 13 3 2
32 2 16 15 13 1 10 9 13 1 9 1 10 9 2 15 13 10 9 16 13 3 0 7 13 9 0 7 3 10 9 2 2
17 2 13 16 4 13 1 10 3 0 10 9 1 13 0 9 2 2
14 3 16 10 9 0 3 13 10 9 1 10 9 0 2
33 2 16 15 13 1 10 0 9 13 1 9 2 4 13 16 15 4 13 7 13 1 9 1 13 2 2 13 10 9 1 10 9 2
15 3 10 9 1 10 9 13 1 4 13 1 15 10 9 2
26 3 1 9 2 1 10 9 1 11 11 2 4 13 13 10 9 13 13 11 11 2 0 9 1 11 2
17 15 13 0 2 15 13 3 2 7 10 9 13 16 4 13 3 2
12 15 13 9 10 9 1 11 11 2 11 11 2
18 2 4 3 13 13 10 9 1 10 9 1 10 9 1 10 9 2 2
28 7 1 0 9 2 4 13 10 9 1 9 1 10 10 9 1 10 9 7 1 10 9 1 9 1 10 9 2
24 13 1 10 9 3 12 9 2 3 10 9 1 10 9 1 10 9 1 10 12 9 13 0 2
46 1 11 2 11 7 11 10 9 2 9 4 3 13 10 10 9 2 16 7 10 11 2 13 1 10 9 1 10 9 2 7 10 9 1 10 9 11 4 3 13 10 10 10 0 9 2
28 10 9 1 9 1 11 13 10 9 1 11 1 10 9 1 10 9 1 10 9 2 11 11 2 1 10 11 2
47 3 7 10 9 7 10 9 4 13 13 16 3 15 13 9 1 1 15 2 16 11 11 4 13 10 9 1 10 9 1 13 10 2 9 2 1 10 9 1 15 1 10 9 1 10 9 2
43 11 11 4 13 10 9 1 11 2 1 10 15 15 13 1 10 9 1 10 11 16 2 12 9 0 4 3 3 13 16 15 13 9 1 10 9 1 9 7 1 9 2 2
10 13 10 9 1 10 9 2 11 11 2
22 15 3 4 13 13 9 1 15 7 1 15 2 15 4 13 10 10 9 0 7 0 2
15 7 1 11 10 10 9 2 11 11 2 13 1 10 9 2
29 1 10 9 1 10 12 1 12 1 10 9 15 13 1 10 11 2 1 0 9 15 13 1 10 9 1 10 9 2
42 10 11 1 11 1 10 9 4 13 10 0 9 0 2 10 12 1 12 1 10 9 2 7 3 10 9 1 10 10 9 3 13 11 11 2 10 9 0 1 11 11 2
28 10 9 0 2 1 10 9 11 11 1 9 1 9 7 11 2 13 3 1 13 15 1 10 3 0 7 0 2
26 7 3 1 11 10 9 11 2 11 7 1 11 15 11 2 11 15 13 1 10 9 1 10 0 9 2
10 15 13 1 15 12 9 1 9 0 2
22 10 9 0 1 10 9 4 13 1 13 10 0 9 7 1 13 9 13 1 10 9 2
21 1 11 1 9 15 13 1 10 9 0 1 10 9 9 13 1 10 9 1 9 2
36 13 10 9 0 11 11 16 13 1 13 10 9 0 1 9 1 9 2 15 1 12 1 10 9 2 2 1 10 9 1 10 11 1 10 9 2
8 15 13 1 15 4 13 15 2
18 15 13 9 1 9 2 9 2 9 1 10 9 1 10 0 9 0 2
18 1 9 1 10 10 0 9 2 10 0 9 4 13 1 10 15 0 2
12 7 2 1 10 9 2 4 13 3 3 0 2
23 3 3 10 9 4 13 10 9 1 10 9 0 2 1 10 9 0 7 1 10 0 9 2
16 1 1 9 0 15 4 13 1 9 1 10 0 9 1 9 2
16 7 3 4 13 2 1 15 13 2 10 0 9 1 9 0 2
36 11 4 13 3 1 11 15 15 1 9 0 4 13 9 2 7 10 9 3 4 13 10 9 0 1 10 11 2 16 4 13 10 0 9 0 2
44 3 1 9 2 10 9 0 1 10 9 4 13 1 10 9 1 9 0 7 9 2 13 9 1 9 1 10 9 1 9 15 13 1 1 10 0 9 1 10 9 2 11 11 2
16 10 15 15 4 13 2 1 0 9 2 9 1 10 0 9 2
30 11 15 4 13 1 13 15 3 2 13 1 10 0 9 15 1 3 0 2 1 15 11 7 11 4 13 10 10 9 2
33 11 11 2 1 10 11 2 15 4 13 2 9 2 2 1 0 9 1 10 9 0 1 10 9 13 1 10 9 1 12 9 3 2
22 7 2 3 2 13 0 13 1 10 10 9 15 15 13 1 10 9 1 10 0 9 2
15 15 15 13 13 11 11 11 2 1 10 9 1 11 11 2
29 7 16 13 0 16 10 9 3 13 1 15 3 15 13 3 4 13 2 0 2 1 10 9 1 15 15 13 3 2
20 15 4 13 10 9 1 12 9 7 1 9 15 10 9 3 4 3 13 3 2
68 1 10 9 0 1 10 9 2 3 3 1 3 3 15 13 10 9 1 15 1 12 9 1 10 9 0 7 3 15 15 13 1 9 2 4 13 10 2 9 2 1 9 7 9 13 1 10 9 13 1 10 10 0 9 13 1 9 10 9 1 10 9 1 11 13 1 11 2
43 1 12 9 2 12 9 2 10 9 7 10 9 2 15 9 1 0 9 7 0 9 13 1 10 9 16 4 13 10 9 2 4 13 1 13 15 1 10 9 2 1 9 2
7 3 2 0 9 1 9 2
29 10 9 10 9 1 10 0 9 11 11 2 16 4 13 10 9 1 10 9 13 1 11 2 13 10 9 1 9 2
40 10 0 9 4 13 1 10 9 1 9 1 9 2 3 10 9 0 2 11 3 13 2 16 3 13 1 10 9 1 9 1 10 9 0 2 13 10 9 2 2
45 13 10 9 3 0 1 15 0 15 4 13 16 10 2 9 1 9 2 2 1 15 10 9 13 0 1 1 15 13 10 9 1 10 9 2 4 13 3 0 7 13 3 12 9 2
37 3 10 12 1 12 1 10 9 13 1 9 0 2 7 10 12 1 12 1 10 9 15 13 1 10 9 2 13 10 9 1 10 9 2 0 2 2
24 1 10 9 7 1 10 9 2 10 9 15 15 4 13 10 9 1 9 2 13 15 1 3 2
32 3 4 3 13 2 15 9 2 16 4 13 10 9 1 11 11 5 11 13 13 1 10 9 1 10 9 1 10 9 1 11 2
44 3 13 3 16 13 10 0 9 2 9 13 7 9 13 1 10 0 9 15 13 1 10 9 1 10 9 1 10 0 9 0 2 4 15 13 1 10 11 7 13 1 10 9 2
13 3 16 16 13 10 9 2 13 16 13 10 11 2
33 1 15 2 3 2 13 1 10 9 1 9 1 10 9 13 10 0 9 15 10 9 4 13 1 10 9 1 10 9 1 0 9 2
44 15 1 10 3 15 4 13 1 10 2 9 2 1 10 9 13 1 13 3 1 10 9 1 10 10 9 2 1 10 2 9 2 0 3 7 0 2 13 16 13 3 9 0 2
47 10 9 1 11 7 1 11 2 3 2 13 1 10 10 9 1 9 0 2 9 15 1 10 9 1 11 3 4 3 13 9 0 13 10 9 13 1 10 9 1 2 13 2 1 11 11 2
14 10 9 13 10 9 1 10 9 1 10 9 1 9 2
25 9 1 9 1 10 9 1 10 9 1 10 9 1 11 7 11 1 10 9 1 9 1 10 11 2
29 3 10 9 4 13 1 13 10 9 13 2 13 16 13 10 9 1 10 9 1 10 11 1 10 9 1 10 11 2
67 1 9 0 2 10 9 13 10 9 0 1 10 9 7 3 10 9 2 15 4 13 13 1 13 1 10 0 9 1 10 9 0 13 15 2 13 10 9 13 3 9 2 1 10 9 1 9 1 10 9 1 9 0 1 15 0 2 2 7 1 9 9 7 1 9 0 2
61 2 13 0 10 9 1 10 13 9 1 10 9 1 10 11 2 4 13 10 9 0 2 9 0 1 13 10 13 15 1 10 9 0 1 9 0 1 9 0 2 0 1 13 10 0 9 15 10 0 9 0 4 3 13 1 9 1 10 12 2 2
9 3 16 1 11 15 15 13 15 2
41 2 13 10 9 3 1 10 9 2 15 13 9 1 10 9 1 15 13 10 9 1 10 9 2 7 15 13 9 1 10 9 1 10 15 2 1 10 9 10 9 2
8 13 9 1 13 9 0 3 2
16 15 13 1 10 11 3 10 9 1 9 0 1 1 9 0 2
15 15 0 1 9 1 10 9 7 15 0 1 13 10 9 2
78 3 3 2 1 9 1 9 7 1 9 2 11 11 4 13 10 9 7 10 9 1 9 1 15 13 2 1 4 15 13 1 10 9 1 10 9 0 0 3 4 4 13 2 4 13 1 11 1 11 1 9 3 9 7 4 13 1 10 0 9 1 11 3 10 9 1 10 9 1 10 9 11 13 1 9 1 9 2
31 10 9 1 9 4 4 13 1 10 9 1 10 9 0 3 9 2 3 16 4 4 13 2 1 10 0 9 1 12 9 2
63 3 2 13 15 10 9 2 15 4 13 10 9 1 10 9 1 11 1 10 9 15 13 1 11 7 13 3 3 3 10 9 1 10 9 1 10 10 9 2 7 3 10 0 9 1 13 3 10 9 0 3 13 1 10 0 9 2 1 10 9 3 0 2
7 13 10 9 7 13 15 2
35 2 13 16 16 4 13 15 1 10 9 2 2 4 13 11 2 2 15 4 13 1 9 1 10 10 9 0 2 7 3 4 4 13 2 2
31 2 10 9 2 2 4 13 11 2 13 1 10 9 2 2 13 10 9 1 10 9 2 1 10 15 4 13 10 9 2 2
18 1 10 9 9 10 9 1 10 9 1 11 13 1 0 9 1 9 2
13 2 2 1 11 13 15 2 11 13 10 9 2 2
12 10 10 9 0 4 13 10 9 3 13 3 2
24 13 3 16 13 16 1 10 10 9 13 0 9 7 9 1 10 9 2 7 13 16 13 3 2
81 10 9 0 15 1 3 10 9 4 13 1 10 9 1 10 11 10 9 3 0 1 10 9 2 13 13 10 10 9 1 12 1 12 9 1 9 2 13 3 10 9 1 10 10 9 1 10 9 2 0 2 1 11 15 13 1 10 9 0 0 10 9 1 2 9 2 7 9 2 13 1 10 0 9 1 10 10 9 9 0 2
57 13 10 0 9 0 1 15 1 10 2 9 2 0 2 7 3 1 9 7 9 7 1 9 0 2 10 9 13 1 15 15 13 9 1 0 9 1 10 9 1 10 9 2 0 1 13 15 3 1 10 9 1 10 2 9 2 2
13 10 11 1 9 16 10 9 15 13 15 4 13 2
66 11 2 11 11 2 7 3 13 7 13 2 10 9 1 11 2 10 11 2 10 9 0 2 10 0 9 2 15 2 3 1 10 9 2 4 13 7 13 1 9 7 9 15 15 13 3 1 16 13 1 10 9 1 10 9 2 1 10 9 0 7 1 10 9 0 2
42 3 2 1 10 13 10 9 11 15 13 0 9 1 10 0 9 1 10 9 0 2 1 10 15 1 10 9 1 9 1 10 9 0 0 10 9 0 13 3 15 0 2
81 1 10 9 1 10 10 0 9 2 2 10 9 4 13 2 15 13 10 9 1 9 2 2 10 9 13 1 10 9 1 10 9 1 10 11 7 13 10 9 1 10 11 1 4 13 10 9 0 2 15 13 1 9 10 9 3 1 10 9 1 10 9 2 2 3 1 13 10 9 7 13 16 13 2 3 1 13 10 9 2 2
19 16 13 2 15 13 10 9 1 13 15 15 13 16 3 13 15 1 13 2
66 15 4 2 13 2 10 9 0 2 13 16 10 9 1 9 13 10 12 5 1 10 12 7 1 10 12 4 3 13 10 12 1 12 2 3 1 10 9 1 9 1 9 9 7 0 9 13 2 10 0 9 0 2 4 3 13 7 3 13 10 12 5 1 10 9 2
7 13 10 9 1 9 13 2
63 4 4 13 1 10 9 1 10 9 1 10 11 1 10 11 2 1 10 9 0 1 10 11 2 10 9 1 11 11 2 12 9 2 10 9 1 11 13 10 12 9 1 10 0 9 7 1 10 10 9 15 4 13 3 10 9 0 2 15 15 4 13 2
22 7 3 3 13 3 7 1 10 0 9 15 13 3 15 3 13 1 10 9 10 9 2
29 1 10 15 2 1 13 1 10 9 2 13 3 13 3 1 10 9 3 13 15 0 3 0 1 9 0 7 0 2
35 10 9 4 13 1 0 10 9 1 10 11 0 2 15 3 2 3 2 4 13 13 1 9 2 7 1 0 9 2 10 9 1 10 9 2
49 10 9 15 4 13 0 1 10 0 9 1 10 9 1 10 9 0 2 7 4 13 10 9 1 10 9 1 9 1 11 1 10 9 13 1 10 9 1 2 0 9 2 2 1 0 9 10 11 2
59 2 15 4 13 16 3 1 10 9 3 4 4 13 9 3 1 10 9 1 9 0 2 13 3 11 11 2 7 15 13 1 13 9 16 1 10 9 13 3 10 9 2 10 9 1 10 10 9 7 10 9 13 3 0 7 3 0 2 2
8 15 13 3 1 10 0 9 2
30 7 15 13 16 3 2 1 10 9 0 1 9 1 10 9 1 9 2 0 1 10 9 1 9 2 15 13 1 9 2
19 15 13 3 15 15 15 13 2 13 10 9 1 9 2 13 1 10 9 2
46 10 0 9 15 15 4 13 0 1 13 1 10 0 11 11 1 10 9 2 3 11 11 4 13 10 2 11 1 11 2 1 11 1 10 9 0 2 13 10 9 0 1 10 10 9 2
21 7 3 13 10 9 1 13 15 15 13 16 1 9 15 13 1 10 9 1 9 2
20 10 9 13 1 13 9 2 3 15 13 13 10 9 1 9 2 1 9 2 2
44 10 11 11 4 13 13 1 10 11 10 9 2 15 1 0 9 1 12 9 0 13 10 9 2 11 9 0 2 13 1 13 11 1 9 1 10 12 2 0 9 1 10 9 2
11 2 15 10 9 1 10 9 1 11 2 2
23 13 3 16 15 4 13 1 9 7 4 13 1 13 10 9 1 10 9 1 9 3 0 2
15 10 9 1 9 1 15 4 13 10 9 3 13 15 0 2
33 7 3 13 3 1 13 15 1 10 11 11 2 16 2 12 9 1 10 9 16 13 10 9 10 9 3 2 13 1 10 10 9 2
23 6 2 15 4 13 13 1 9 1 10 11 11 5 11 2 7 3 4 13 15 1 0 2
12 15 4 13 1 9 3 3 1 10 10 9 2
21 2 3 10 12 1 10 9 9 15 4 13 2 7 4 4 13 1 12 9 2 2
21 9 2 10 9 1 11 13 10 9 0 2 13 3 1 13 10 9 1 10 9 2
55 7 10 9 4 13 10 9 1 10 13 9 1 9 11 2 10 15 4 3 13 15 15 0 13 1 10 9 1 10 9 1 13 16 10 9 13 0 1 13 2 1 13 10 9 0 1 10 9 1 11 2 1 12 9 2
20 11 4 4 3 13 13 1 9 1 11 15 13 10 9 1 9 10 9 0 2
11 11 7 11 15 4 13 9 1 0 9 2
26 10 9 4 4 13 3 1 11 15 3 3 4 4 13 0 9 1 9 1 10 9 1 3 1 11 2
18 15 13 10 9 1 10 9 4 13 16 3 4 13 7 13 10 9 2
8 15 1 16 13 1 10 9 2
13 7 13 3 10 0 15 13 3 13 10 10 9 2
11 1 10 9 15 4 13 10 9 1 9 2
44 13 3 10 9 1 13 3 1 3 10 9 1 10 9 1 9 2 1 13 3 16 10 9 2 13 1 15 15 13 2 13 0 2 13 3 1 10 9 10 2 1 10 9 2
25 1 10 9 1 10 9 0 2 11 4 13 10 9 0 2 13 10 10 9 2 1 13 10 9 2
32 15 13 3 2 3 2 3 10 9 1 10 9 1 9 11 1 10 9 1 10 12 7 1 11 0 9 3 15 15 4 13 2
2 13 2
38 16 13 1 10 9 1 4 13 10 0 9 15 13 10 9 0 3 4 13 1 10 2 9 0 2 15 3 13 1 1 15 10 9 1 10 0 9 2
24 13 16 13 3 0 16 10 9 2 3 2 3 13 3 3 0 1 10 1 15 3 13 9 2
69 7 13 16 2 11 11 2 2 3 16 10 9 2 10 9 0 2 10 9 0 1 10 12 1 10 9 1 9 1 10 9 1 10 9 0 2 16 4 13 1 10 0 9 1 10 9 13 3 10 9 1 9 2 15 4 13 15 3 10 9 13 1 10 9 1 9 1 9 2
35 9 0 2 1 9 1 9 1 12 9 15 13 10 9 0 2 13 10 9 1 9 1 10 9 7 10 9 1 0 9 1 10 9 0 2
65 10 9 3 15 13 1 0 9 2 10 9 2 3 16 10 9 0 7 0 15 4 13 10 9 1 10 9 1 11 2 4 13 10 9 1 15 1 10 3 0 7 0 1 10 9 1 13 9 1 10 9 1 10 2 9 0 2 16 4 13 1 10 0 9 2
80 13 10 9 10 9 2 3 16 13 1 10 9 1 10 9 1 9 1 10 9 2 11 2 1 10 11 11 2 10 9 1 11 2 10 9 1 9 1 11 2 10 12 7 10 9 1 9 1 11 11 7 10 9 1 10 9 1 11 11 2 15 13 3 3 1 13 10 9 1 10 9 0 13 1 0 9 1 10 9 2
10 2 3 13 10 9 0 10 9 0 2
20 15 1 10 12 8 2 15 13 1 10 9 1 10 11 7 13 10 9 0 2
25 3 3 2 7 10 9 1 13 15 1 9 13 10 9 1 9 2 1 15 9 0 13 3 0 2
66 1 10 0 9 1 9 2 1 9 10 9 0 15 4 13 1 9 2 7 10 9 1 11 11 4 4 13 1 10 9 1 10 9 12 2 1 9 1 10 9 1 10 9 1 11 11 2 7 1 15 1 10 0 9 0 15 13 10 9 0 2 3 0 1 11 2
9 2 13 15 15 4 13 2 2 2
45 15 15 15 4 13 2 4 13 15 10 9 1 10 9 1 3 2 10 9 11 2 15 15 4 13 9 1 10 9 11 2 15 13 10 0 9 1 9 1 9 9 1 10 9 2
26 13 1 16 13 1 13 2 11 11 2 1 11 11 2 10 0 9 15 10 9 15 13 1 10 9 2
30 4 3 13 2 10 9 1 11 11 2 1 11 11 2 10 9 7 4 4 13 15 2 7 3 3 13 10 9 3 2
29 10 11 1 3 3 13 15 1 16 13 1 10 9 13 1 10 9 7 1 10 15 10 10 9 4 4 13 3 2
19 13 16 15 13 13 1 9 2 10 0 9 2 2 9 15 15 3 13 2
13 2 11 2 1 10 9 1 10 2 9 2 2 2
16 4 13 10 9 1 11 13 3 1 10 11 1 10 10 9 2
34 7 10 10 9 1 11 11 2 1 10 10 0 9 0 2 3 13 3 0 1 13 15 4 13 2 7 13 10 3 0 9 1 9 2
36 15 13 13 7 13 10 9 1 10 10 9 0 2 15 15 1 9 13 7 13 9 1 9 7 15 4 13 1 10 9 2 13 15 1 9 2
32 10 9 2 2 10 9 2 2 1 13 10 9 1 10 9 13 1 10 9 0 2 10 0 2 2 15 15 4 13 2 2 2
37 10 11 2 11 11 2 11 11 2 10 11 11 2 11 11 11 11 2 11 11 7 11 11 13 10 9 3 1 9 1 10 9 1 10 9 0 2
46 9 12 2 1 9 2 16 4 3 13 2 13 1 11 2 1 10 11 2 11 11 2 1 15 1 10 9 3 13 1 10 9 15 15 13 1 9 9 12 7 9 12 9 1 11 2
39 10 2 9 9 2 1 10 9 13 10 9 1 10 2 11 11 2 13 1 9 1 10 9 1 10 9 1 10 9 0 15 13 9 1 10 9 10 9 2
38 10 0 12 9 15 4 13 2 3 2 2 13 16 1 10 9 0 3 13 10 9 1 9 1 10 9 2 13 3 10 9 1 10 9 1 9 0 2
20 2 1 9 9 13 3 1 9 1 9 2 13 3 1 9 1 10 9 2 2
10 2 1 12 9 3 13 10 11 2 2
8 10 9 1 10 9 3 0 2
12 9 1 10 9 1 10 9 1 11 7 11 2
7 10 9 4 13 1 9 2
11 4 13 10 9 13 7 13 10 9 13 2
25 10 9 0 2 3 10 9 2 7 15 13 10 9 1 10 9 13 1 15 15 4 13 13 15 2
36 3 3 4 13 10 10 9 1 15 15 13 2 16 3 0 9 2 1 10 9 15 13 2 10 9 1 3 2 10 9 1 3 10 9 0 2
30 16 4 13 1 9 3 1 10 0 9 1 10 9 9 1 15 4 4 13 10 9 1 10 9 0 13 3 1 11 2
13 1 11 9 1 10 9 1 10 9 1 10 9 2
10 11 11 15 15 13 1 10 9 12 2
15 9 1 9 2 9 2 9 2 9 1 9 2 9 0 2
28 15 13 13 1 10 9 1 10 9 2 1 10 9 0 7 0 1 10 11 2 0 9 13 1 9 1 9 2
20 15 13 13 1 10 9 1 10 0 9 7 3 2 1 9 2 13 1 9 2
9 3 2 15 13 7 15 15 13 2
28 15 13 9 16 15 2 1 10 12 9 1 10 11 13 1 10 11 11 2 13 15 1 15 15 13 7 13 2
13 13 13 0 13 13 3 10 0 9 1 10 9 2
38 11 2 3 2 4 13 10 10 9 2 15 15 4 1 9 13 3 1 15 2 16 15 4 13 2 1 10 9 16 10 9 0 13 3 1 9 2 2
13 2 1 3 10 9 13 15 7 3 15 2 2 2
33 7 11 13 10 9 3 13 1 10 9 0 7 0 2 0 1 10 10 9 1 9 2 9 2 9 2 9 2 9 1 9 2 2
54 0 7 3 0 2 10 9 9 13 1 10 11 13 1 13 9 0 1 10 9 0 1 10 9 2 7 10 9 1 10 9 1 12 9 13 1 10 9 11 13 1 9 10 0 9 1 10 9 1 9 0 2 0 2
27 15 13 10 9 1 13 10 9 1 11 2 11 2 1 10 0 9 11 15 4 13 10 9 1 10 9 2
60 3 2 1 1 10 11 13 1 0 9 10 9 1 9 15 13 3 9 1 10 9 0 2 10 9 13 3 1 3 13 1 10 0 12 5 1 9 1 0 9 7 9 0 1 10 9 1 10 9 1 9 1 10 9 0 1 10 9 0 2
32 13 1 13 3 10 9 15 13 1 10 9 1 10 9 1 10 9 1 10 9 13 10 9 0 1 10 9 1 9 7 9 2
56 10 11 13 1 0 9 7 16 1 11 4 13 10 10 9 1 10 9 1 10 0 9 0 2 13 1 9 0 2 1 9 1 10 12 2 10 9 1 9 1 9 0 0 15 13 10 11 11 1 10 9 1 10 9 0 2
50 13 10 9 1 13 1 10 9 1 10 9 10 9 3 16 4 4 13 1 10 10 9 0 7 16 4 13 3 1 10 9 15 2 1 10 9 1 12 9 2 4 13 13 10 10 9 1 9 0 2
46 2 13 2 13 11 11 2 16 0 1 10 9 1 10 9 13 1 10 9 10 0 7 0 9 1 9 15 10 9 2 3 2 10 9 2 15 13 13 1 10 9 1 10 9 2 2
20 3 10 10 9 13 1 13 15 13 9 3 1 9 1 10 9 1 10 9 2
70 10 15 4 4 13 2 13 1 10 9 10 9 0 1 10 9 2 15 4 13 13 3 10 9 1 10 9 2 10 9 0 0 4 13 3 1 10 9 10 9 13 1 10 12 7 2 16 15 13 9 13 9 2 11 4 1 10 9 13 3 1 10 9 10 9 1 10 12 2 2
21 3 2 1 10 9 1 9 1 10 9 2 1 10 9 7 10 9 1 10 9 2
33 7 10 9 1 10 9 15 13 3 1 10 9 13 1 10 9 1 9 1 10 9 1 10 9 15 4 13 10 9 1 10 11 2
40 1 10 9 0 2 11 4 13 1 10 9 1 10 15 4 4 13 10 9 0 1 13 1 9 10 9 0 1 9 2 13 1 10 9 1 10 9 1 9 2
34 2 11 4 13 1 11 11 1 12 9 2 3 1 13 9 2 7 3 4 3 13 11 2 13 11 11 2 15 4 13 10 9 13 2
22 13 16 10 11 13 10 9 0 7 0 2 1 9 1 10 0 9 0 1 10 12 2
19 3 16 10 9 13 0 2 4 13 15 10 9 0 1 9 1 10 12 2
10 3 2 13 1 10 12 1 12 2 2
10 2 6 2 10 9 3 15 13 2 2
39 11 2 10 9 15 3 13 10 10 12 9 2 9 1 9 2 9 2 13 1 4 13 10 9 0 2 1 10 9 1 11 2 2 11 2 1 9 0 2
14 2 13 10 0 9 2 13 2 1 10 11 0 2 2
22 2 10 11 2 15 13 10 9 2 13 1 10 9 1 9 7 1 2 9 2 2 2
11 2 13 10 9 1 10 9 0 2 2 2
31 10 9 1 13 2 13 16 10 10 9 1 9 0 4 3 13 16 10 9 1 10 9 13 2 10 9 7 10 9 2 2
10 10 9 0 1 10 10 9 1 9 2
18 7 3 15 13 1 10 9 1 9 1 10 10 9 10 9 1 11 2
6 2 15 13 13 2 2
23 1 10 0 9 2 10 9 1 9 13 1 9 11 13 1 10 0 11 7 1 11 11 2
57 13 1 15 1 10 9 15 4 13 10 9 1 13 1 11 15 1 10 9 3 0 1 10 9 1 9 1 10 9 1 10 12 2 10 9 1 15 1 15 13 15 4 13 15 2 1 10 9 1 9 1 10 9 1 9 0 2
19 1 10 9 1 9 0 13 16 10 9 15 13 1 10 9 1 9 0 2
40 9 1 9 3 1 9 9 11 2 10 9 13 10 9 0 1 0 9 2 1 11 1 11 2 1 11 1 11 2 11 2 11 2 1 9 1 10 9 9 2
18 13 10 9 10 9 13 10 9 13 10 0 2 15 13 15 2 2 2
18 10 9 4 13 10 10 0 9 1 10 0 9 15 15 4 13 9 2
13 11 15 13 10 9 15 13 16 13 0 1 13 2
34 10 9 1 11 4 13 10 0 9 15 4 13 10 9 3 0 2 9 15 1 15 3 15 13 3 1 10 3 0 9 1 9 11 2
9 3 13 15 1 13 15 1 9 2
9 10 9 1 9 1 10 9 0 2
11 10 9 13 1 9 1 9 1 10 9 2
32 10 9 1 9 1 9 2 12 9 1 9 7 9 2 12 9 13 1 10 9 0 7 0 7 10 0 9 1 10 9 0 2
37 3 1 10 9 3 1 10 9 1 10 9 0 10 9 4 13 1 10 9 0 2 3 15 15 13 3 1 9 1 10 9 15 3 13 3 0 2
31 7 2 1 10 9 12 2 10 9 13 3 0 1 10 9 1 9 13 1 10 9 2 1 10 9 0 13 1 0 9 2
14 13 16 1 11 2 10 9 0 13 0 10 0 9 2
13 2 13 16 13 7 1 10 0 9 13 11 2 2
22 7 16 15 13 1 10 9 2 13 7 16 3 4 13 10 9 7 3 15 4 13 2
36 2 3 13 15 13 9 1 10 9 2 1 15 3 3 13 15 2 3 15 1 16 13 1 15 15 4 13 12 9 3 1 11 7 11 2 2
17 3 1 10 9 1 10 11 13 13 3 13 10 10 9 1 9 2
60 11 11 11 7 11 11 11 2 1 10 13 10 9 1 10 9 13 1 10 11 11 1 11 1 10 12 2 10 9 7 10 9 2 11 2 11 2 13 10 9 1 10 9 1 10 9 1 9 1 10 10 9 2 7 1 10 10 9 0 2
37 2 16 10 9 13 1 13 15 1 10 9 16 15 4 13 10 9 2 2 3 10 9 1 10 9 1 11 12 15 4 13 1 13 10 10 9 2
91 13 3 16 13 9 11 2 2 15 4 13 2 7 4 13 10 9 1 10 9 1 10 9 0 15 15 13 1 10 9 2 2 2 13 10 9 16 10 9 2 3 1 10 13 15 1 9 1 9 1 9 13 1 9 7 9 3 7 3 0 2 13 10 9 1 15 1 10 13 1 10 0 9 2 1 10 9 1 9 0 2 10 9 13 1 10 9 15 13 0 2
19 13 10 9 7 15 13 16 10 9 2 1 9 2 3 15 13 1 9 2
23 3 15 13 1 9 3 10 9 1 10 12 9 2 15 1 9 15 13 3 16 13 9 2
26 15 1 16 13 1 10 9 1 9 2 9 2 9 7 9 15 15 13 1 13 1 9 1 10 9 2
15 3 2 9 1 10 0 1 11 3 15 15 4 3 13 2
29 4 13 10 9 1 10 11 2 7 13 1 9 1 10 10 9 13 1 9 1 13 9 2 1 13 2 13 9 2
48 13 1 13 15 10 9 3 0 13 3 0 16 10 0 9 2 3 1 0 9 0 2 3 4 4 13 1 15 7 1 15 1 10 0 9 1 9 1 10 9 2 1 9 10 9 0 2 2
48 10 9 4 13 1 10 0 9 2 15 3 0 2 3 15 13 16 1 10 9 1 10 9 10 12 9 13 13 10 9 1 12 9 7 16 4 4 13 3 15 13 1 10 9 3 3 0 2
30 7 15 13 3 10 0 9 15 13 1 10 9 1 15 15 4 13 1 11 7 1 10 9 1 10 9 1 10 9 2
13 7 1 10 9 1 9 0 10 9 13 3 0 2
31 10 9 3 13 3 1 9 10 9 2 3 16 1 10 9 1 10 9 0 10 9 15 4 13 1 11 11 7 11 11 2
21 7 10 9 4 13 15 3 13 10 0 9 1 10 9 15 13 1 10 9 0 2
47 3 2 15 4 13 2 16 1 10 9 1 11 1 10 11 7 1 11 11 2 1 10 9 1 10 9 1 10 11 2 3 1 10 9 3 13 1 15 1 13 2 13 10 9 1 11 2
15 11 4 3 3 3 13 1 10 9 2 11 11 1 9 2
28 7 15 13 3 15 13 11 9 1 10 11 2 1 9 1 11 1 11 2 15 13 9 1 10 9 1 11 2
46 1 10 13 3 1 10 9 1 9 13 1 10 11 2 10 9 1 10 0 2 1 9 2 4 4 13 3 1 3 2 2 15 13 1 13 10 2 9 2 4 13 10 9 1 9 2
9 1 9 2 15 13 3 9 0 2
48 16 15 15 15 4 13 3 1 11 11 4 13 2 1 13 15 1 10 9 1 10 9 2 2 10 9 13 7 10 9 13 2 1 3 1 10 9 1 9 2 2 10 9 15 4 3 13 2
32 10 9 15 13 13 3 1 10 0 9 1 10 9 0 2 13 15 1 10 9 1 9 1 10 9 1 9 0 1 15 0 2
51 1 10 0 9 1 9 2 10 9 13 1 9 10 0 9 1 10 9 11 2 13 1 10 9 11 11 7 15 13 10 9 1 10 9 1 10 9 1 9 1 10 9 1 10 12 5 1 10 9 0 2
15 7 15 4 13 10 9 15 13 13 15 1 9 10 9 2
8 10 9 1 11 2 11 2 2
15 9 1 9 1 9 1 10 11 2 9 1 10 9 11 2
12 13 3 10 9 1 13 7 13 10 10 9 2
32 1 9 1 10 9 2 13 3 10 0 9 1 10 9 1 9 7 10 9 1 10 0 9 1 10 9 1 10 9 0 0 2
29 0 3 13 10 0 9 15 13 10 9 1 10 9 1 13 1 15 13 10 9 1 3 2 16 1 15 15 13 2
8 13 3 16 13 15 1 9 2
6 13 1 13 10 9 2
3 13 3 2
25 13 13 10 9 0 1 10 9 7 13 15 1 10 9 1 9 1 10 0 9 2 13 9 2 2
14 7 13 16 10 2 9 2 1 10 12 4 13 15 2
21 15 13 3 10 9 0 0 15 4 13 10 0 9 0 1 9 13 1 9 0 2
11 9 13 1 10 9 1 13 11 7 11 2
64 1 13 7 13 10 9 1 10 9 1 10 2 11 2 4 13 3 12 9 1 10 9 7 2 13 2 10 9 4 13 1 10 9 1 10 9 2 15 1 11 13 3 1 10 0 9 2 13 1 10 0 9 0 2 15 15 4 13 9 1 10 0 9 2
11 9 13 2 9 0 7 10 9 1 9 2
8 3 10 0 9 1 13 9 2
22 3 15 3 2 1 10 9 13 2 10 9 0 2 10 9 1 9 2 10 9 13 2
20 10 9 15 13 7 13 9 0 7 15 13 3 10 9 3 0 10 9 0 2
19 1 10 0 9 10 9 15 3 15 13 1 10 9 1 9 13 10 11 2
14 10 0 9 1 10 9 0 13 1 13 0 10 9 2
51 10 9 1 15 10 11 13 13 10 9 1 9 7 10 11 13 1 13 15 1 10 9 1 9 2 15 13 3 15 15 13 10 9 1 10 9 0 1 10 9 7 1 10 9 1 10 9 1 10 9 2
68 13 15 10 9 1 10 9 0 1 10 11 2 11 11 2 15 13 10 12 9 2 3 13 2 16 2 3 4 3 13 1 9 10 9 13 16 13 1 13 15 10 9 2 2 7 13 16 13 10 9 0 1 10 9 0 13 10 9 0 1 9 1 10 9 1 10 9 2
32 15 3 15 4 13 10 9 1 13 10 9 1 9 7 1 13 10 9 1 9 2 7 10 9 1 10 9 3 0 1 9 2
36 11 2 15 3 13 10 9 1 10 9 0 3 1 13 1 11 2 3 4 13 10 9 1 10 9 0 13 10 0 9 1 10 11 11 11 2
18 2 10 9 13 10 9 1 10 9 1 15 3 15 13 10 9 2 2
28 2 13 16 16 4 13 15 1 10 9 2 15 4 13 1 9 1 10 10 9 0 7 3 4 4 13 2 2
79 1 10 12 9 9 2 1 10 12 1 10 9 1 10 9 2 1 10 12 13 10 9 2 1 10 12 10 11 2 9 0 0 2 1 10 11 2 1 10 12 10 9 2 1 10 12 10 9 2 1 10 12 1 10 11 2 1 10 12 1 10 11 2 1 10 12 1 9 1 10 9 2 1 10 12 1 10 9 2
38 1 10 0 9 4 13 3 10 11 1 10 9 0 7 0 2 13 1 10 9 7 0 1 13 10 9 1 10 9 1 11 7 1 10 10 9 0 2
40 11 2 0 2 4 13 9 3 1 10 10 0 9 2 15 15 4 13 2 15 4 13 1 9 7 2 13 1 10 9 0 2 4 13 2 1 9 1 9 2
25 16 13 0 2 10 9 13 10 9 0 1 9 2 7 3 0 7 0 1 10 10 9 1 9 2
16 2 1 10 10 10 9 3 4 3 13 15 1 10 9 2 2
27 1 9 1 10 9 10 9 13 1 9 2 3 7 3 2 7 3 15 13 10 9 0 1 10 9 0 2
75 2 7 3 13 13 10 9 2 10 9 1 10 9 1 11 7 15 1 10 9 7 9 3 1 11 11 1 11 2 13 13 10 9 2 10 9 2 10 9 2 10 9 7 3 1 10 9 0 15 15 13 16 10 9 3 13 10 9 0 2 10 9 0 7 1 9 0 4 13 1 10 0 9 2 2
58 10 0 9 1 11 13 9 1 11 11 2 1 15 13 1 9 2 11 2 1 11 11 2 1 10 9 15 13 10 9 1 9 1 9 1 10 9 1 10 9 2 1 10 9 1 10 9 13 10 9 1 10 9 13 1 10 9 2
79 1 11 13 10 0 9 1 10 15 4 13 1 10 9 0 15 15 4 13 13 9 1 9 2 13 15 1 10 10 3 0 9 1 11 2 2 11 2 13 2 13 1 2 11 11 2 2 13 9 1 10 9 1 2 10 9 1 11 11 2 7 1 15 1 10 0 2 11 2 2 1 10 15 4 13 3 1 9 2
10 2 2 10 9 15 13 2 13 2 2
29 1 12 9 0 2 1 10 9 1 10 9 2 2 2 11 2 13 1 9 1 10 9 15 3 15 13 10 9 2
38 13 1 11 3 1 10 0 11 11 2 13 1 11 2 10 9 13 10 9 13 1 9 12 9 1 9 13 1 10 9 0 1 15 1 9 15 13 2
40 1 10 0 9 1 9 2 10 9 13 10 9 1 9 15 13 9 10 9 7 10 9 0 2 7 10 3 0 9 0 0 2 10 11 2 1 0 9 0 2
23 13 13 2 10 0 9 15 13 13 10 9 15 13 1 10 9 2 3 15 4 3 13 2
17 3 15 4 13 1 13 10 9 1 10 12 2 13 1 10 9 2
5 3 15 4 13 2
62 10 9 15 4 13 1 11 10 9 0 2 10 9 0 2 7 10 0 9 15 13 10 9 1 11 11 1 13 10 9 2 4 13 10 9 1 0 9 2 16 11 13 1 13 10 9 1 9 1 9 2 7 16 15 15 4 13 13 1 10 9 2
15 7 15 13 1 13 16 3 15 13 3 1 9 10 9 2
31 7 3 13 3 1 15 2 15 13 1 9 2 10 9 2 7 1 10 9 15 13 1 10 9 13 0 3 15 1 15 2
34 16 15 13 13 2 0 2 1 9 1 10 9 0 2 1 10 0 9 1 10 9 2 15 13 10 9 2 16 4 13 13 10 9 2
17 7 3 3 13 13 10 9 1 10 9 1 9 2 0 7 0 2
28 11 2 15 13 3 1 15 2 15 15 13 13 13 2 15 15 13 3 2 7 15 13 3 1 13 10 9 2
10 10 9 15 15 13 3 1 13 15 2
8 1 9 15 15 13 3 3 2
22 3 16 13 1 10 9 0 2 7 15 13 13 10 9 2 13 0 7 13 1 11 2
47 7 1 10 15 11 1 9 11 3 15 4 13 13 7 1 10 9 2 7 1 10 9 2 16 15 4 13 9 1 15 1 11 2 10 15 13 10 9 7 13 12 9 1 11 1 9 2
37 3 15 13 1 11 15 13 1 10 9 1 10 9 1 10 9 2 7 1 10 13 15 2 3 15 13 7 0 7 0 16 3 4 13 9 10 2
27 1 15 2 1 9 2 13 1 13 15 3 1 10 9 0 2 7 3 13 9 1 13 15 1 0 9 2
10 15 13 1 9 16 15 13 1 15 2
31 7 10 9 15 13 1 10 9 2 1 10 9 1 10 9 1 13 13 10 10 0 9 1 9 15 15 4 13 10 9 2
17 2 13 2 16 3 4 13 3 2 3 15 13 10 9 1 13 2
27 13 11 2 3 4 13 3 16 4 13 1 10 9 11 1 10 9 11 13 1 9 1 9 1 10 9 2
26 2 10 9 2 9 11 2 13 10 9 16 3 15 13 2 7 4 13 15 1 10 9 15 13 15 2
51 7 3 1 13 3 4 13 10 10 9 15 15 4 13 1 13 15 13 2 1 10 9 1 13 10 9 2 16 10 9 15 13 2 7 16 13 0 11 15 13 1 10 9 1 3 13 13 10 10 9 2
22 3 16 4 13 10 10 9 1 10 9 2 15 13 1 13 15 3 3 1 10 9 2
18 2 4 10 9 13 15 15 13 10 9 1 13 3 2 13 11 11 2
48 1 11 11 13 10 9 1 9 2 10 15 13 10 9 1 9 2 15 15 13 12 9 1 9 1 0 9 10 15 1 10 9 2 15 15 4 13 2 7 13 1 13 10 9 1 10 9 2
23 2 13 15 3 15 15 13 10 9 2 16 15 13 2 16 13 10 9 2 13 10 9 2
38 10 9 16 15 13 3 1 10 9 2 3 15 13 3 2 3 16 3 15 4 3 13 2 7 3 11 13 10 9 1 10 9 15 4 13 10 9 2
15 11 7 11 3 15 4 3 13 1 10 9 1 10 9 2
42 11 3 15 13 10 9 2 7 13 16 4 13 1 15 2 7 15 4 13 10 9 7 15 15 4 13 1 10 9 2 16 15 15 4 3 13 1 9 16 13 0 2
13 7 15 3 15 13 3 13 15 2 15 13 0 2
27 10 9 15 13 10 9 16 15 13 13 2 0 1 10 9 2 1 10 13 0 7 0 1 10 9 0 2
75 1 10 9 1 9 7 9 2 1 15 3 15 13 1 9 9 0 2 10 9 11 13 10 0 9 0 15 15 13 13 1 10 9 2 1 10 9 0 1 10 9 2 1 10 9 0 1 10 9 0 2 15 15 13 1 10 9 2 3 3 2 1 10 11 0 2 3 10 9 15 13 1 10 9 2
42 11 13 9 7 9 2 7 1 10 9 15 13 1 9 10 9 13 1 9 7 1 9 2 1 10 9 3 15 2 16 15 13 13 1 10 9 0 7 0 10 9 2
9 3 15 15 13 13 3 2 3 2
9 15 4 13 10 9 1 10 9 2
12 16 3 15 13 13 3 1 15 7 1 15 2
32 7 4 4 13 15 10 9 1 3 13 15 1 10 11 2 15 16 15 15 13 1 10 15 15 13 13 10 9 7 10 9 2
58 10 11 15 13 13 2 0 7 0 2 1 10 9 15 13 1 10 9 2 7 3 15 13 1 10 0 9 2 3 13 10 9 2 13 1 13 15 3 2 1 10 9 0 1 9 1 9 0 2 7 13 15 15 1 10 9 0 2
18 13 10 9 1 0 9 2 7 13 13 10 9 16 13 1 10 9 2
23 16 15 15 4 13 13 1 10 10 9 2 4 13 16 3 13 0 9 1 11 11 13 2
88 3 13 16 10 9 1 10 9 15 13 1 10 9 1 10 9 15 1 10 9 1 10 9 0 2 1 10 9 2 16 10 0 9 15 13 1 10 9 2 16 13 1 10 9 2 1 10 9 1 10 9 2 13 1 9 1 13 15 10 9 2 1 15 7 1 10 9 2 1 13 15 16 11 15 4 13 1 13 1 10 9 2 7 15 15 4 13 2
49 15 13 1 10 9 1 13 15 2 7 13 1 13 1 10 9 3 16 15 4 13 10 9 2 1 13 15 3 1 10 9 2 16 3 10 9 7 10 9 15 13 0 1 10 0 1 10 9 2
32 2 13 2 2 9 9 2 2 2 15 13 2 16 15 13 10 0 9 1 9 10 2 16 13 0 9 2 15 13 10 9 2
20 15 15 13 15 1 3 16 11 15 13 13 10 9 1 10 9 0 1 9 2
88 1 10 9 15 13 10 2 0 9 0 2 13 1 10 9 11 0 2 1 11 7 1 10 9 0 1 11 2 15 15 13 1 10 11 11 2 1 10 12 9 1 10 12 9 2 7 15 13 3 3 13 1 10 9 1 10 0 9 9 13 1 10 9 1 11 7 3 1 10 9 10 9 1 10 0 9 15 13 10 0 9 1 9 1 10 9 0 2
9 10 9 13 1 10 13 10 9 2
50 10 9 2 13 15 15 13 1 9 2 7 1 9 12 9 3 1 10 0 2 13 1 0 1 13 15 2 7 4 13 15 1 9 2 1 13 15 10 9 0 2 16 15 13 10 9 1 10 9 2
78 16 13 1 15 10 0 9 1 9 2 16 10 9 4 13 1 10 9 2 16 13 1 10 9 15 3 13 15 1 13 2 7 13 10 9 1 9 1 13 15 10 9 1 10 9 0 2 7 3 16 15 13 10 9 2 16 15 3 13 1 10 9 10 15 13 13 15 13 1 9 0 1 10 9 1 10 9 2
9 3 4 13 15 15 13 1 9 2
55 10 9 2 1 9 2 16 13 10 9 2 15 1 10 9 2 13 15 10 9 1 13 2 7 10 9 15 3 13 9 3 1 13 15 2 7 10 9 10 15 13 1 10 9 1 13 10 9 1 10 9 2 4 13 2
18 2 13 1 13 16 15 3 4 13 10 9 1 15 9 15 4 13 2
56 16 10 9 13 0 1 9 2 10 10 9 13 0 2 10 9 0 2 7 10 9 0 1 10 9 2 16 10 10 9 3 15 15 13 10 9 2 7 4 13 15 3 0 9 1 9 2 3 1 13 10 9 1 10 9 2
27 15 13 16 13 9 1 10 9 1 9 2 7 13 13 1 15 15 15 13 1 9 10 9 7 10 9 2
30 10 9 1 10 0 9 1 10 15 7 10 15 1 10 15 13 10 9 1 3 10 10 9 1 11 1 10 9 0 2
31 9 0 2 3 3 1 10 10 9 2 7 3 1 10 9 1 9 0 2 13 15 15 15 13 1 10 9 1 10 9 2
8 9 0 1 10 9 1 11 2
21 7 3 15 13 1 3 13 10 9 1 9 7 15 13 13 1 3 13 10 0 2
43 1 9 2 3 10 9 1 10 15 10 9 4 3 13 13 1 13 10 9 15 4 13 15 2 3 2 1 10 9 13 7 4 3 13 1 9 7 2 3 1 9 0 2
28 10 9 1 10 0 2 1 10 9 2 1 10 9 4 4 3 13 1 15 1 0 1 10 10 9 1 9 2
34 1 10 9 1 10 9 12 2 15 13 3 10 9 1 9 15 13 1 9 10 10 9 7 1 10 9 1 9 0 7 1 15 0 2
65 3 1 10 9 2 3 2 10 9 13 3 1 13 15 2 13 2 3 9 1 10 9 15 2 1 3 13 1 10 9 0 7 3 2 0 2 2 4 13 0 9 7 10 0 9 0 2 15 13 13 15 10 9 1 10 9 11 11 7 1 10 9 11 11 2
59 10 11 2 1 9 2 15 13 1 13 1 10 0 2 9 2 15 13 3 13 10 9 1 13 10 10 9 7 2 9 3 0 2 3 13 1 13 15 10 9 2 10 9 7 10 9 0 1 10 9 7 1 10 9 1 10 0 9 2
40 1 10 9 1 9 0 2 7 1 10 9 1 10 11 11 2 0 1 10 9 0 1 10 10 9 2 10 9 1 10 9 13 10 10 9 1 13 10 9 2
18 10 9 13 3 1 10 9 0 10 9 1 10 10 0 9 1 9 2
37 2 1 10 0 9 4 4 13 10 9 0 7 15 4 13 16 15 4 13 2 3 1 9 2 1 10 9 1 10 9 1 9 1 10 9 0 2
18 15 3 2 16 13 3 2 10 9 0 1 10 9 0 3 13 0 2
26 3 1 10 11 2 10 9 0 1 10 9 1 9 0 13 9 1 10 9 1 10 9 1 0 9 2
31 1 10 9 0 13 16 10 9 7 10 9 4 13 1 10 9 1 15 10 9 0 4 13 1 10 9 0 1 10 9 2
45 1 10 0 9 15 13 3 1 10 9 1 9 2 15 4 13 2 1 10 9 15 13 3 3 2 1 10 9 2 0 2 0 1 10 0 9 1 9 0 1 9 2 9 2 2
26 10 9 1 9 13 10 9 16 13 1 9 1 9 2 13 9 2 15 4 3 13 1 2 9 2 2
49 15 4 13 9 15 3 13 1 10 9 2 13 10 9 12 2 7 9 2 0 2 15 4 4 13 1 10 9 2 3 1 9 12 2 1 15 2 9 2 13 1 10 12 9 11 7 11 2 2
75 10 9 2 1 3 10 9 0 2 2 15 13 1 3 0 1 13 7 1 10 9 1 9 7 1 15 1 9 1 9 2 4 13 10 9 2 15 13 2 11 7 15 12 2 2 11 12 2 2 1 13 10 9 1 9 0 2 13 10 9 0 15 1 9 13 10 9 1 9 2 15 13 3 2 2
15 11 4 13 10 9 1 10 9 7 1 15 13 1 9 2
13 10 9 15 13 1 10 9 7 3 3 1 3 2
22 7 1 10 9 1 9 1 9 7 1 10 9 1 9 10 9 13 3 0 1 13 2
44 10 12 9 1 9 0 4 4 13 1 9 0 2 10 0 1 10 15 13 0 1 9 1 9 2 7 10 0 13 12 7 10 9 2 7 10 9 13 2 1 9 3 0 2
60 3 2 15 13 16 1 10 0 9 1 10 9 1 10 9 1 9 2 3 9 3 0 2 1 10 9 7 10 9 2 7 10 9 1 0 9 2 4 4 13 1 10 9 2 3 13 2 2 1 13 10 9 1 9 2 15 13 3 2 2
38 1 10 9 0 1 10 9 7 1 10 9 1 10 9 0 1 10 9 2 15 13 2 3 2 11 2 11 12 8 2 7 2 11 7 15 12 2 2
56 1 10 9 1 9 1 10 9 0 2 10 9 4 13 1 9 0 2 16 0 9 4 13 1 10 9 2 7 1 9 2 16 10 9 0 4 4 13 1 10 9 1 9 0 7 2 3 2 4 4 13 1 9 0 2 2
50 10 9 4 4 13 1 10 9 0 15 13 1 13 10 9 1 10 9 2 13 15 10 9 7 10 9 2 4 4 13 1 10 9 1 10 9 1 10 9 7 13 3 10 9 0 1 10 9 0 2
27 3 2 3 16 15 13 0 1 10 9 1 9 0 2 10 10 9 4 13 1 10 9 1 4 13 3 2
32 1 9 2 1 10 9 0 2 10 9 4 4 13 1 10 9 3 0 2 15 4 1 9 13 1 13 10 0 9 1 9 2
23 1 10 9 0 4 13 10 9 1 9 2 0 2 1 9 1 9 2 10 9 1 9 2
17 1 10 9 13 16 10 9 0 7 0 4 4 13 1 10 9 2
3 12 9 2
33 10 0 9 13 10 0 9 1 13 0 10 9 15 2 1 15 2 13 0 16 10 9 4 4 13 0 1 10 9 1 9 0 2
37 10 9 4 13 1 9 1 9 13 1 9 1 10 9 9 2 9 2 1 2 1 9 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2
35 10 9 4 4 13 1 10 9 1 10 9 1 10 9 13 1 10 9 1 9 2 1 10 9 1 10 11 11 2 1 10 10 9 0 2
44 1 9 2 10 9 2 1 9 1 15 13 1 10 9 0 2 13 10 9 12 2 2 4 13 9 1 12 9 2 7 10 10 9 0 13 3 16 10 10 10 9 13 0 2
29 3 1 10 9 2 10 9 0 1 10 9 2 15 13 10 9 12 2 13 0 10 0 9 1 10 9 1 9 2
32 1 9 2 11 13 10 9 3 0 1 9 0 3 13 2 3 16 10 9 13 3 0 2 16 15 4 13 2 1 10 9 2
52 10 9 0 15 13 1 10 9 0 2 11 7 11 1 10 9 2 4 1 9 13 1 13 10 9 1 10 9 0 2 15 4 13 1 10 9 2 3 13 2 1 10 9 15 4 4 13 1 10 9 0 2
42 16 13 2 10 9 1 9 1 9 0 0 2 7 15 3 13 10 9 2 13 10 9 1 13 9 3 13 15 13 1 13 1 10 9 1 10 9 1 10 9 0 2
21 15 1 10 9 1 13 10 0 9 0 2 15 13 10 9 12 1 10 9 2 2
20 15 13 3 3 10 9 1 9 2 15 13 10 9 11 2 11 3 3 2 2
35 1 10 9 1 9 10 11 11 13 10 9 1 9 1 10 9 1 10 9 1 10 9 0 13 13 10 9 0 1 13 1 10 9 13 2
35 15 13 10 9 1 13 10 9 1 10 9 1 10 9 0 2 1 15 1 10 9 2 1 13 15 2 15 1 9 3 3 0 13 9 2
69 10 9 2 10 9 1 12 9 13 1 10 11 11 7 13 1 10 9 1 9 13 1 10 9 11 11 2 9 1 9 1 10 9 1 10 9 1 11 2 13 2 9 1 10 9 2 15 15 4 13 2 10 9 1 10 9 0 2 1 10 9 7 10 9 1 10 9 0 2
50 10 9 15 3 13 13 10 9 1 15 2 3 15 13 0 7 13 9 1 10 9 2 7 1 10 9 16 15 13 1 15 7 1 10 10 9 2 16 13 1 10 9 2 3 0 7 13 15 13 2
62 7 3 13 3 2 13 2 1 10 9 1 11 15 3 13 2 7 15 4 13 3 3 2 1 2 13 2 10 9 2 1 13 1 10 9 10 9 16 10 9 4 13 1 10 9 0 10 10 9 2 15 15 10 9 13 2 10 9 1 9 2 2
31 3 15 13 16 10 9 1 11 13 1 13 1 9 1 10 0 9 1 10 9 13 1 13 15 1 10 9 1 10 11 2
35 7 9 1 10 12 1 10 12 2 16 10 0 0 9 2 16 3 15 13 2 4 13 1 10 9 10 10 9 0 2 11 15 4 13 2
17 3 1 10 11 9 1 10 2 9 1 10 9 2 1 10 11 2
6 11 13 2 11 13 2
42 16 10 9 1 9 13 15 15 13 2 15 15 13 7 3 9 2 13 0 16 3 13 10 9 13 3 10 9 1 10 9 0 1 10 9 1 10 9 1 10 9 2
29 9 1 9 2 10 9 1 9 2 10 3 0 2 13 10 9 1 9 7 9 15 13 10 9 1 10 9 2 2
31 3 3 10 9 4 13 1 13 2 10 9 1 10 9 1 10 9 2 1 11 7 11 4 4 13 1 10 9 1 9 2
37 1 10 12 1 3 9 2 1 10 9 1 10 9 2 13 1 9 10 9 1 9 15 2 1 10 9 1 3 2 4 13 1 15 1 12 9 2
61 2 3 2 15 13 10 9 7 15 13 11 2 4 13 2 1 10 9 1 10 9 0 11 11 2 10 9 1 10 0 9 2 11 11 11 2 2 15 1 9 4 13 0 10 2 9 2 1 10 9 1 11 11 2 11 2 11 2 1 11 2
6 11 11 13 1 9 2
13 1 10 9 0 1 10 9 15 13 2 9 2 2
53 4 4 13 0 2 1 9 0 9 7 9 2 7 10 9 4 4 13 1 9 13 3 1 13 15 1 11 11 7 13 1 10 9 15 4 13 2 0 2 1 10 9 0 2 15 1 10 9 13 10 9 11 2
26 1 10 9 2 4 13 10 9 1 13 15 1 9 2 3 10 9 0 1 10 15 10 9 11 11 2
46 13 1 13 1 3 10 10 9 13 1 2 9 15 13 2 1 10 9 1 10 9 2 1 3 3 15 13 11 2 2 11 13 1 10 9 13 10 0 7 0 11 11 1 9 0 2
7 11 7 11 13 15 11 2
11 9 1 0 9 2 3 2 1 11 11 2
61 15 13 15 15 13 2 11 2 2 1 10 9 1 9 0 7 0 2 16 1 10 9 1 10 11 13 3 10 9 1 13 7 3 3 15 13 10 9 1 13 15 3 2 16 13 0 16 1 9 9 15 13 10 9 0 1 10 9 2 9 2
38 15 13 11 11 2 13 12 9 2 13 3 2 7 13 3 1 10 9 1 10 11 11 1 13 15 1 10 11 1 10 9 2 9 1 10 11 9 2
12 15 13 11 7 13 10 9 1 10 11 11 2
47 11 15 4 13 3 0 2 13 1 15 10 9 1 10 9 2 13 1 9 0 9 2 1 10 3 9 1 10 0 11 1 11 11 2 11 2 13 10 9 1 10 10 0 9 1 3 2
33 10 9 3 0 15 2 3 1 13 1 9 10 11 1 11 2 13 9 1 10 9 1 10 9 1 15 3 13 2 10 11 11 2
24 15 13 10 9 2 15 3 15 13 2 11 9 2 2 7 15 13 10 9 1 13 10 9 2
47 10 0 9 7 10 9 13 10 9 1 13 10 9 7 9 1 9 2 10 9 0 15 13 3 2 3 16 13 10 9 15 13 10 9 1 10 9 1 10 13 2 1 9 10 10 9 2
30 10 9 0 15 13 9 1 9 7 13 1 10 13 3 16 10 0 9 4 13 15 7 3 1 10 9 1 10 9 2
27 10 9 11 4 13 10 9 1 10 12 2 13 1 11 2 10 0 9 2 2 10 9 15 13 16 0 2
29 10 9 1 10 9 2 3 4 13 10 9 2 4 4 3 13 9 9 16 10 12 9 15 13 1 13 1 9 2
11 10 9 1 10 9 2 3 2 13 0 2
14 1 9 2 10 9 1 9 13 15 13 7 15 13 2
44 13 2 1 15 15 4 13 13 1 11 2 10 9 0 2 1 9 15 1 11 2 9 2 11 11 2 11 11 2 13 10 0 9 3 1 15 15 15 13 3 2 9 2 2
16 7 13 10 9 16 13 10 9 2 15 13 11 7 11 11 2
50 1 10 12 4 13 10 9 0 1 9 1 10 11 15 2 15 13 3 1 10 9 1 0 9 1 13 10 0 9 0 2 13 9 2 15 13 1 0 9 15 1 4 13 1 9 7 0 9 2 2
57 1 13 1 11 2 1 10 11 11 11 2 15 1 10 15 13 10 9 2 9 2 3 0 2 10 9 0 1 10 11 11 11 4 3 13 2 11 2 2 1 10 9 0 1 10 11 2 3 13 10 9 3 0 1 10 9 2
39 10 9 2 10 9 1 11 15 13 1 9 13 1 11 7 1 11 2 10 10 0 9 2 15 4 13 11 2 1 12 9 10 9 2 3 12 12 9 2
40 10 0 9 15 13 15 13 2 11 11 2 2 9 0 2 7 10 9 1 10 9 2 3 3 13 2 2 13 2 13 10 9 0 1 16 13 0 2 2 2
20 11 11 2 13 3 1 9 1 10 9 1 10 9 2 15 15 13 1 9 2
42 1 11 7 11 13 3 10 9 1 10 11 15 13 1 3 1 9 1 10 0 9 1 9 1 11 1 13 10 9 1 10 9 0 0 1 10 9 1 10 0 11 2
40 13 16 10 9 15 13 1 10 9 3 0 2 1 10 9 11 2 7 13 16 15 13 9 1 10 9 1 10 9 2 7 13 10 9 7 13 1 10 11 2
11 15 13 10 9 15 4 13 3 10 9 2
11 4 13 10 9 7 4 13 1 10 9 2
24 11 1 10 11 2 11 2 1 12 2 11 2 12 9 12 2 4 13 10 9 7 9 0 2
42 10 10 9 0 2 13 3 3 1 9 1 9 0 2 13 1 9 1 9 1 10 9 0 2 0 1 15 10 0 0 9 1 10 9 1 10 9 2 11 1 11 2
31 13 10 9 3 0 7 3 0 1 10 9 0 3 1 13 16 15 2 16 3 13 2 4 13 13 10 9 1 10 9 2
14 3 1 10 0 9 0 15 13 10 9 0 1 11 2
55 0 9 1 10 9 0 7 0 2 9 0 1 10 9 2 9 13 1 10 9 1 15 15 4 13 15 2 9 0 1 10 9 1 9 7 10 15 1 13 0 9 2 9 3 0 7 0 2 15 13 10 10 10 9 2
31 11 13 1 11 1 10 11 2 9 7 9 2 7 1 11 1 11 1 11 1 10 9 0 13 1 10 12 1 10 12 2
47 15 13 3 16 2 3 1 10 10 9 2 4 3 13 2 11 11 2 2 7 2 11 11 2 7 2 11 11 2 2 7 10 9 1 10 11 16 4 13 10 9 1 10 9 13 0 2
55 15 13 10 0 9 1 10 9 1 11 1 11 2 3 3 0 1 11 2 7 3 9 1 10 9 2 16 13 10 12 9 12 10 9 1 10 9 1 10 9 1 10 9 7 1 10 9 0 1 10 9 1 10 9 2
44 15 4 13 3 10 9 1 10 9 1 11 11 7 0 9 13 16 11 13 10 9 2 7 13 0 13 10 9 1 10 9 2 1 10 9 16 1 11 3 15 13 10 9 2
21 3 0 2 1 10 9 1 11 2 13 10 9 1 11 3 3 3 1 10 12 2
24 10 9 0 1 11 7 15 0 7 0 1 11 3 13 1 9 1 10 9 1 10 0 11 2
49 1 10 11 2 13 1 11 3 1 11 1 10 9 1 11 11 1 10 2 9 1 10 9 1 10 9 1 10 9 2 7 16 2 13 1 9 2 15 13 0 2 2 4 3 13 1 11 11 2
64 10 0 10 9 15 15 4 13 13 10 11 1 10 9 2 3 1 10 0 9 11 11 2 10 9 13 9 1 11 7 13 1 10 0 9 1 11 1 10 12 1 11 11 2 1 13 13 1 10 9 12 2 12 2 1 10 15 13 3 9 1 11 11 2
16 1 10 9 1 10 9 4 13 10 9 2 3 10 9 0 2
36 1 10 12 13 3 0 1 11 11 3 2 10 12 9 1 10 12 13 1 10 9 1 10 11 10 9 1 10 9 1 10 9 1 10 9 2
34 10 9 13 10 9 1 10 9 1 12 9 7 10 10 0 9 2 3 1 10 9 1 13 7 3 13 10 9 1 10 12 9 0 2
63 1 9 2 10 9 1 10 9 15 13 2 1 9 1 10 9 3 13 2 1 15 1 12 9 2 16 13 10 9 1 10 9 11 11 11 2 1 9 1 11 2 13 1 10 12 1 10 9 2 15 1 10 0 9 13 10 9 15 13 10 0 9 2
18 13 1 10 9 1 11 11 2 1 10 12 4 13 1 10 9 0 2
8 10 9 15 13 1 12 9 2
11 1 3 2 10 11 2 1 9 1 11 2
25 3 2 1 0 9 2 11 11 1 11 2 10 9 13 2 10 11 7 11 11 2 13 15 0 2
27 13 3 10 9 11 7 11 11 2 10 11 1 10 9 7 10 9 11 7 11 1 11 2 3 15 0 2
24 1 11 1 10 12 13 1 10 9 1 10 11 7 1 10 9 1 11 11 2 9 13 2 2
34 1 10 12 13 1 11 2 13 1 11 11 11 1 13 1 10 9 11 3 13 10 9 0 13 11 11 11 1 9 3 1 11 11 2
17 3 13 11 11 11 2 7 15 13 3 1 11 2 11 7 11 2
19 10 9 0 4 13 1 13 11 1 11 1 10 9 1 11 11 1 11 2
33 1 10 12 13 3 1 11 11 11 3 2 1 10 9 0 2 13 10 9 1 10 9 1 10 9 0 1 10 9 1 11 11 2
34 3 3 2 13 1 9 11 0 2 15 13 1 11 2 3 13 9 1 10 9 1 11 11 11 2 1 10 9 13 3 10 9 2 2
19 1 10 0 9 1 11 1 10 12 13 1 9 3 13 1 10 9 0 2
22 1 10 9 15 4 13 13 10 9 1 11 2 10 9 2 10 11 0 7 10 9 2
24 13 3 1 11 1 10 9 1 11 1 11 3 13 1 9 1 11 1 11 7 1 11 11 2
26 13 10 9 1 10 9 1 10 9 7 1 10 9 2 10 0 9 2 10 11 1 11 7 10 9 2
21 13 1 11 1 10 12 2 13 9 1 10 12 7 13 1 11 10 12 9 12 2
37 1 10 0 9 4 13 1 10 0 9 1 10 9 7 3 1 13 13 10 11 11 11 2 10 11 11 11 11 7 10 9 1 9 13 11 11 2
52 13 1 11 11 11 10 4 13 10 9 0 1 10 9 1 10 11 1 10 11 1 11 2 11 1 10 11 12 2 9 1 9 12 2 2 9 3 13 7 13 1 0 9 2 2 0 2 16 13 10 9 2
27 1 10 10 9 13 10 9 11 1 11 2 1 15 4 13 1 11 1 10 9 1 10 9 1 11 11 2
30 13 3 1 0 9 10 9 13 1 10 9 1 11 11 1 10 11 1 11 1 11 2 1 15 13 3 0 9 0 2
36 11 1 10 11 4 13 12 9 0 1 15 13 0 10 9 1 9 0 2 13 1 10 9 1 10 9 2 7 9 0 2 13 1 10 9 2
45 10 0 9 4 13 10 8 8 8 8 8 2 10 9 13 1 10 9 2 15 4 13 9 0 1 9 0 2 0 2 13 3 1 10 9 1 4 15 13 1 9 1 10 9 2
58 1 10 0 9 8 8 8 4 13 10 9 1 9 13 1 10 9 0 2 13 0 9 1 10 9 1 4 15 13 15 1 10 9 1 10 0 9 0 2 7 1 10 9 4 13 10 9 2 1 3 13 3 0 1 10 9 0 2
24 1 10 9 13 13 10 9 1 10 9 1 10 9 7 10 9 0 1 10 9 1 10 9 2
27 1 15 13 10 9 1 10 0 9 2 9 1 9 2 4 4 13 1 9 0 1 3 0 1 10 9 2
34 10 9 0 7 15 0 4 13 3 0 3 1 10 9 1 10 10 9 2 3 1 10 9 0 1 15 10 9 4 13 9 3 0 2
36 10 10 9 13 3 1 0 9 0 1 10 9 1 9 7 13 10 9 0 1 9 1 10 9 1 10 9 1 10 9 1 10 9 1 11 2
11 10 11 11 13 10 9 0 9 9 0 2
58 13 15 1 10 12 1 10 9 11 11 1 10 9 11 11 2 10 9 11 11 7 11 11 2 10 9 11 11 7 10 9 11 11 2 10 9 13 3 9 1 11 11 1 10 12 2 1 9 1 10 9 1 10 9 9 0 9 2
25 1 10 12 4 13 10 0 9 9 1 9 0 7 1 10 12 13 10 10 0 9 10 0 9 2
29 1 10 9 9 2 12 2 2 11 11 13 10 9 1 10 12 1 13 15 1 10 0 9 0 2 10 11 11 2
17 11 11 2 3 1 10 9 0 13 9 7 11 13 1 10 9 2
11 11 13 3 10 9 1 10 9 11 11 2
26 1 10 9 1 9 7 0 9 2 1 10 12 2 13 10 0 0 9 1 10 11 11 2 10 9 2
25 1 10 9 10 9 13 10 10 9 2 13 1 10 9 0 3 0 2 0 7 0 1 10 9 2
12 0 9 15 15 13 1 10 9 1 9 0 2
41 1 10 12 13 10 9 13 0 9 7 10 9 0 10 9 10 9 15 2 15 13 3 10 9 1 10 9 3 0 7 0 2 3 1 9 1 10 9 3 0 2
39 1 10 9 1 9 2 11 13 10 9 7 15 13 10 9 11 11 2 1 9 9 7 3 9 0 2 7 10 9 11 11 2 7 11 13 1 10 9 2
43 1 10 12 13 9 2 9 13 1 13 2 3 0 2 2 15 15 13 3 3 1 10 0 9 2 0 2 7 3 1 10 9 1 9 0 7 15 13 3 9 7 9 2
86 10 9 0 7 10 9 1 10 9 13 2 1 10 12 2 1 8 8 2 9 3 0 3 1 10 0 2 15 13 15 1 10 9 3 13 1 10 9 1 10 0 9 1 10 9 2 3 1 10 9 15 1 15 13 10 9 3 0 2 2 1 9 0 7 0 2 13 1 9 0 13 1 10 9 0 15 4 13 7 13 1 13 10 9 0 2
11 10 9 15 13 10 9 13 3 3 0 2
25 1 10 12 13 10 9 0 2 8 8 15 13 15 1 12 9 1 9 2 9 2 9 2 3 2
30 1 10 12 4 13 10 0 9 1 9 1 10 9 2 13 1 10 9 7 13 2 2 9 0 7 9 1 10 9 2
48 1 10 9 8 8 8 2 12 2 13 9 2 9 12 2 2 13 1 10 9 3 0 7 0 2 7 15 15 13 1 10 9 0 7 1 10 9 0 2 3 3 3 0 3 1 10 9 2
37 10 9 3 15 13 3 1 15 1 8 8 2 1 15 10 9 15 4 13 0 1 0 9 2 3 13 15 2 1 10 9 2 3 13 7 13 2
35 1 10 12 2 1 10 9 9 9 13 9 2 9 15 13 3 10 9 1 9 2 1 10 9 13 1 10 9 3 13 1 10 9 9 2
22 10 9 13 2 0 2 7 10 9 15 13 1 9 0 1 10 0 9 1 10 9 2
15 1 10 9 1 10 12 11 11 13 10 9 1 9 0 2
37 1 10 9 1 11 2 10 2 9 2 3 13 10 9 1 10 9 1 10 9 2 0 9 9 2 2 10 15 4 13 1 10 9 1 10 9 2
36 3 10 0 9 1 10 9 3 13 10 9 1 10 9 1 10 11 11 2 1 16 1 10 9 9 7 9 15 4 13 1 3 0 7 0 2
33 3 2 10 9 2 15 13 10 0 9 2 13 3 0 2 7 15 13 13 1 9 1 2 0 9 2 7 2 0 2 9 2 2
26 1 10 9 2 13 16 10 9 13 0 9 0 1 10 9 2 15 13 10 9 1 2 9 11 2 2
35 10 11 11 4 3 13 10 9 1 2 10 9 1 9 2 2 9 1 10 11 0 1 10 9 0 2 3 13 2 10 0 9 2 2 2
23 10 9 4 4 13 1 10 9 13 9 1 10 11 2 0 9 2 10 9 1 11 2 2
9 10 9 4 13 1 0 9 9 2
16 4 3 13 2 12 9 9 2 2 0 9 1 10 11 11 2
30 10 9 13 0 1 10 9 9 11 11 9 2 1 9 1 10 9 7 3 15 4 13 1 9 9 2 3 1 9 2
47 10 9 9 4 13 1 10 12 7 13 10 9 1 10 9 0 9 9 7 9 2 7 16 13 10 9 13 10 9 15 13 10 9 9 1 13 10 9 2 10 9 7 10 9 1 9 2
29 3 10 0 9 2 7 1 0 9 10 3 0 2 13 10 9 1 9 2 9 7 3 10 9 1 9 7 9 2
44 1 10 9 10 9 0 4 4 13 3 1 10 9 2 7 4 4 13 9 0 1 9 1 13 1 9 3 3 9 2 9 7 0 9 2 7 3 9 7 9 1 10 9 2
13 10 9 13 10 9 1 10 9 1 9 1 9 2
31 10 9 0 1 10 9 13 10 9 1 10 9 2 10 9 0 1 10 9 15 13 1 13 9 1 9 1 9 3 0 2
42 1 10 9 0 2 10 9 13 10 9 1 9 2 15 4 13 1 10 9 1 10 9 3 0 2 3 1 10 9 0 1 10 9 2 10 0 9 1 10 9 2 2
23 3 1 10 9 10 0 9 4 13 1 10 9 0 2 15 13 1 9 1 10 9 13 2
24 16 15 13 10 9 2 10 9 13 4 13 7 3 13 1 10 9 7 4 13 1 10 9 2
50 13 10 9 15 13 1 10 9 1 10 9 7 10 9 1 10 9 13 0 13 1 10 9 15 13 10 9 2 13 16 10 9 1 15 15 13 10 9 13 0 7 13 0 1 10 9 1 10 9 2
8 11 13 10 9 1 10 9 2
8 11 13 10 9 1 10 9 2
18 11 13 10 9 13 1 10 9 1 13 10 9 7 13 1 10 9 2
36 10 9 1 9 1 10 9 4 13 3 10 3 0 0 2 3 13 10 9 1 10 9 13 16 13 10 9 0 1 15 10 9 4 13 9 2
15 3 2 10 9 3 4 4 13 16 3 4 13 10 9 2
28 10 9 1 9 1 10 9 13 10 0 9 0 2 7 10 9 0 1 15 10 0 9 1 9 4 13 9 2
65 10 0 9 1 10 15 13 0 13 9 4 1 9 13 2 1 10 9 1 10 9 2 13 3 2 2 1 10 9 1 9 7 1 10 10 0 9 1 9 1 10 9 0 1 10 9 2 10 10 9 7 1 10 9 15 13 10 9 1 10 9 1 10 9 2
42 10 9 13 1 10 9 1 10 9 1 10 9 1 10 9 1 10 9 7 1 10 9 1 9 1 10 9 13 10 9 1 10 9 1 10 9 1 9 1 10 9 2
34 10 9 1 12 9 0 2 7 10 9 9 1 10 0 9 2 1 10 9 3 0 2 13 9 7 9 1 10 9 1 10 9 13 2
58 1 10 0 9 13 1 9 0 2 9 15 15 13 3 2 15 13 10 9 1 9 0 2 16 10 9 1 9 1 9 9 13 3 3 9 9 1 9 1 13 2 1 10 9 1 9 1 10 9 2 10 9 1 9 1 10 9 2
51 1 10 9 1 3 10 9 4 13 1 9 2 7 1 10 9 9 15 2 13 2 10 9 9 1 9 7 13 10 0 9 15 13 2 13 2 10 9 0 1 10 9 13 1 10 9 1 10 9 0 2
15 10 9 4 3 13 1 10 9 9 1 10 9 1 9 2
46 3 1 10 9 1 9 10 9 13 1 9 1 13 1 10 9 2 15 1 10 9 0 3 15 13 1 9 1 9 1 9 2 10 9 0 7 1 10 9 3 0 3 10 9 9 2
14 10 9 2 9 7 9 13 1 10 9 1 10 9 2
45 10 0 1 13 10 9 9 1 13 2 10 9 1 9 0 0 2 13 11 11 2 15 1 10 12 13 10 9 1 13 10 9 1 10 9 1 10 9 2 7 3 10 10 9 2
32 1 10 9 1 10 12 11 11 13 10 0 1 13 10 9 1 10 9 1 10 9 7 1 10 9 1 9 1 10 0 9 2
43 1 10 12 11 11 13 10 9 1 10 9 1 13 1 9 9 0 7 1 10 12 1 10 9 0 15 13 10 9 1 10 9 1 9 0 1 10 15 10 9 11 11 2
59 10 0 2 0 1 10 9 7 1 10 9 1 10 9 2 15 13 1 10 9 11 11 2 10 0 7 0 9 15 1 10 9 0 13 3 10 9 7 13 10 9 2 7 3 13 10 9 7 10 9 0 1 13 1 10 9 9 0 2
59 10 9 1 10 9 3 13 3 1 9 1 10 9 1 11 7 3 1 10 9 1 9 11 2 13 3 1 10 9 1 10 9 1 9 1 10 9 2 10 9 1 10 9 13 3 10 9 0 1 13 10 0 9 0 13 9 7 9 2
21 1 10 12 10 0 11 11 13 10 0 1 13 10 9 13 1 10 9 1 11 2
25 10 9 13 1 10 9 1 10 9 1 10 9 1 13 10 0 9 7 9 1 10 0 9 0 2
29 1 10 9 10 9 1 10 9 4 4 13 1 10 9 1 10 9 0 0 2 9 0 7 9 1 10 9 0 2
39 10 9 13 16 10 9 1 10 9 13 13 1 10 0 9 1 10 9 2 3 10 9 1 10 9 13 13 3 0 2 1 9 1 10 9 13 3 0 2
45 10 9 1 10 9 1 10 9 0 4 13 9 1 10 9 1 9 1 9 1 9 1 10 0 9 0 7 13 3 1 9 7 1 10 9 0 7 1 15 0 1 10 10 9 2
19 4 4 13 1 10 11 11 1 10 11 2 7 1 9 0 1 10 11 2
23 10 0 9 1 10 9 13 10 9 15 13 10 9 1 10 9 13 0 7 1 10 9 2
35 10 0 9 1 10 9 1 9 9 2 1 10 9 7 10 9 0 2 11 2 2 4 3 13 10 9 13 1 10 9 0 1 10 9 2
25 1 9 0 4 13 3 0 13 2 13 7 3 13 10 9 0 7 13 16 10 9 13 10 15 2
5 10 0 9 0 2
54 1 10 0 9 13 3 2 15 13 10 9 1 2 0 9 2 1 9 1 10 9 13 2 7 10 9 1 9 9 1 10 0 9 7 9 7 13 2 1 9 1 13 13 10 9 3 0 7 0 1 15 3 13 2
18 10 9 1 15 7 1 10 0 3 0 9 13 10 9 1 9 9 2
48 10 9 0 1 3 3 13 3 0 1 9 2 0 2 1 15 13 2 16 13 9 1 9 13 1 9 0 9 2 11 2 7 1 0 9 11 2 8 8 8 2 7 11 2 8 8 8 2
32 1 15 10 9 1 9 1 9 2 1 9 9 2 7 10 9 1 9 1 10 9 2 1 13 3 10 9 13 1 15 13 2
41 10 9 9 2 1 10 0 9 5 9 2 9 2 13 2 3 1 10 9 9 7 1 15 2 15 1 10 9 1 9 0 1 10 9 11 2 0 9 2 0 2
16 10 0 9 1 10 11 13 11 2 0 0 9 2 9 0 2
30 13 1 10 9 0 1 9 9 15 13 1 10 9 1 10 9 13 10 9 1 10 9 7 13 0 9 1 10 9 2
54 9 1 10 9 4 13 10 9 1 9 2 1 10 9 1 3 13 13 1 10 9 10 9 1 9 1 9 1 9 2 7 10 9 1 10 9 1 9 9 2 1 10 9 1 13 1 10 0 9 10 9 1 9 2
7 13 12 9 1 9 9 2
31 10 9 0 4 13 1 9 15 13 10 7 10 9 10 9 13 1 10 9 2 13 3 0 9 1 10 9 1 10 9 2
5 10 9 0 13 2
44 10 9 4 13 1 9 2 9 7 9 0 1 0 9 15 2 13 0 9 1 9 2 13 10 9 0 1 0 9 9 2 1 9 1 10 15 13 3 0 13 10 9 0 2
42 10 9 4 3 13 1 0 9 2 13 10 0 7 0 9 7 9 1 9 15 2 1 10 9 1 9 0 1 13 10 9 1 9 2 4 13 2 9 1 9 2 2
36 1 9 2 3 4 13 1 9 1 9 1 9 7 9 1 9 7 9 0 2 1 13 10 9 1 10 9 7 13 10 9 1 9 7 9 2
24 10 9 9 2 1 9 2 9 9 2 2 13 9 0 1 10 9 2 7 13 3 3 0 2
15 4 13 1 9 0 1 9 0 13 1 13 10 9 9 2
13 13 3 0 1 10 9 2 4 13 1 9 0 2
34 10 9 9 2 1 9 9 2 13 9 7 9 15 13 1 13 10 9 13 10 9 1 15 0 1 15 1 10 9 15 15 4 13 2
24 1 13 10 9 3 0 2 1 10 9 4 13 13 1 9 1 13 10 9 1 10 0 9 2
35 16 3 0 13 3 0 2 16 4 13 10 9 1 0 9 2 13 1 10 0 9 13 1 13 15 1 10 9 1 9 1 10 10 9 2
38 10 9 4 13 13 1 9 10 9 1 13 15 13 1 10 9 3 0 1 10 10 0 9 2 13 10 9 15 13 1 10 9 7 1 10 9 0 2
14 10 9 13 1 9 1 13 9 0 7 1 13 9 2
50 10 9 0 13 10 9 1 9 0 1 10 15 10 9 1 9 10 2 9 2 13 9 3 0 7 0 1 13 10 9 1 10 9 1 10 9 0 7 1 13 10 9 1 9 13 1 9 7 9 2
14 10 12 9 0 13 10 9 1 9 7 10 9 0 2
25 10 9 1 9 7 9 9 15 13 16 10 9 2 9 2 13 10 10 10 9 1 10 0 9 2
39 10 9 13 1 9 1 13 10 9 1 9 1 9 1 0 9 2 7 13 3 0 1 10 9 1 9 3 0 15 13 9 13 1 2 9 1 9 2 2
31 1 13 10 9 1 9 1 9 1 13 1 9 10 9 1 9 2 13 0 13 10 9 3 2 3 3 13 1 10 9 2
28 10 9 1 9 7 0 9 15 13 16 10 9 1 0 9 1 10 9 4 13 13 1 9 1 10 9 13 2
38 1 10 9 2 15 13 10 9 1 13 10 9 1 9 2 7 1 3 10 9 3 13 3 1 10 10 9 7 15 13 10 9 1 10 9 1 9 2
19 1 10 9 2 10 9 13 1 9 1 13 10 0 9 1 9 9 0 2
24 10 9 1 9 7 9 9 13 10 9 3 0 13 1 9 1 9 1 13 1 10 9 3 2
37 10 9 13 15 1 4 13 10 9 3 2 7 10 9 13 10 9 1 9 3 0 2 16 13 1 10 9 1 13 10 10 9 1 10 9 0 2
15 1 9 2 10 9 4 13 2 0 9 15 13 1 15 2
32 10 2 9 9 2 13 10 9 1 9 9 1 10 15 4 13 10 9 1 9 1 10 0 9 7 15 4 13 10 0 9 2
39 10 11 1 10 9 0 9 9 9 2 9 0 1 10 9 9 2 13 10 9 3 0 15 13 1 10 9 1 10 9 9 13 7 9 1 10 9 13 2
22 10 9 13 4 13 2 13 7 13 1 9 1 13 10 9 1 15 15 10 9 13 2
57 1 10 9 15 4 13 10 9 1 9 0 2 16 15 4 13 10 9 2 10 9 7 10 9 1 10 9 13 2 3 13 10 9 1 9 2 10 9 9 7 13 9 1 9 1 9 1 13 1 10 9 0 1 10 9 9 2
20 1 10 9 2 10 9 4 4 13 1 9 0 7 13 10 9 1 9 0 2
18 10 9 0 0 13 3 0 1 9 1 10 9 10 1 10 9 0 2
12 15 13 3 7 1 10 9 0 16 15 0 2
27 10 9 0 0 4 13 1 10 9 1 9 1 9 0 0 15 13 0 1 10 0 9 0 1 10 9 2
20 10 9 1 10 9 1 9 0 4 4 13 1 10 0 9 1 10 9 0 2
11 1 15 2 1 10 9 10 9 13 0 2
31 1 13 10 9 1 10 9 10 9 0 13 10 9 1 10 9 9 2 13 3 10 9 0 13 15 1 1 10 0 9 2
53 10 9 0 13 1 9 1 13 15 1 10 9 1 9 1 10 9 2 1 9 2 0 13 10 9 1 10 9 1 10 9 9 1 9 2 0 13 10 9 1 13 10 9 7 13 1 13 10 9 1 10 9 2
41 10 0 9 13 1 9 1 10 9 2 13 1 10 13 10 9 13 13 15 1 9 0 13 3 2 1 10 9 1 13 3 0 1 10 9 10 9 7 10 9 2
20 13 3 0 13 10 9 9 3 13 7 0 1 10 9 7 1 10 10 9 2
27 10 9 4 13 1 9 7 2 13 9 16 10 9 13 0 2 4 13 1 10 9 1 13 10 0 9 2
17 16 3 13 1 9 2 10 9 4 13 0 9 1 10 9 9 2
14 15 13 9 16 12 9 3 0 13 1 10 0 9 2
9 10 9 0 13 9 1 10 9 2
43 10 9 13 10 9 1 10 2 9 15 13 2 2 2 0 9 2 1 9 2 10 9 15 15 13 1 10 9 9 7 15 4 3 13 10 9 9 13 15 1 0 9 2
19 10 9 3 13 0 1 10 9 1 9 2 16 3 4 1 9 13 0 2
31 10 9 13 3 3 0 1 10 9 1 10 9 13 7 13 1 9 2 3 1 9 1 9 7 9 13 1 12 9 0 2
14 10 9 1 9 4 3 13 13 1 10 9 1 9 2
20 10 0 9 1 9 13 15 15 13 1 0 9 13 13 1 1 10 0 9 2
17 10 9 13 15 1 15 10 9 13 1 13 1 10 9 1 9 2
35 10 9 4 13 13 9 7 9 1 10 0 9 2 7 13 10 9 9 1 10 9 1 10 9 1 10 9 2 1 9 2 9 2 2 2
29 16 3 13 10 9 2 3 1 9 0 2 0 9 2 1 9 1 10 9 2 15 13 9 0 1 9 1 9 2
53 16 10 9 15 13 10 9 1 10 15 13 10 9 3 4 13 1 10 9 1 9 2 7 13 0 11 2 9 9 9 2 2 10 9 0 13 1 9 0 1 10 9 7 10 9 4 13 1 7 3 1 15 2
14 10 9 1 10 9 13 1 9 13 3 10 9 0 2
50 10 9 9 4 4 13 1 10 9 13 1 10 0 9 2 1 10 9 2 10 9 1 10 9 7 10 9 1 10 9 1 10 9 13 10 9 3 0 2 7 0 1 10 0 9 1 10 9 0 2
37 13 1 9 9 13 1 10 9 1 13 10 9 1 10 9 13 1 10 9 11 7 1 10 9 0 2 7 3 10 11 2 1 10 9 1 9 2
14 10 9 13 13 3 0 1 15 0 2 7 3 0 2
28 1 10 9 2 10 9 9 2 9 1 11 9 2 1 9 13 1 11 2 11 2 11 2 13 10 0 9 2
16 10 9 0 15 13 2 13 7 13 10 9 1 10 9 0 2
17 10 9 0 15 13 10 9 13 1 9 1 10 9 13 7 13 2
43 1 9 10 9 1 10 9 1 9 4 13 9 1 3 13 10 9 1 10 9 1 9 2 8 8 5 8 5 0 2 1 15 1 9 2 8 8 5 8 5 0 2 2
33 1 10 9 0 2 10 9 1 10 9 2 10 9 2 10 9 0 7 0 4 13 1 10 0 9 1 10 0 9 1 9 0 2
31 10 9 0 0 0 13 3 10 9 1 9 2 1 3 2 9 1 10 9 7 10 9 1 9 1 9 0 2 11 2 2
30 10 9 9 3 2 13 4 13 3 1 9 0 9 1 9 2 11 2 2 1 9 0 2 0 7 0 2 1 9 2
42 15 13 1 10 9 1 13 3 1 10 9 2 1 1 13 1 10 0 9 2 7 13 10 9 1 9 0 1 13 10 9 1 10 9 0 1 13 15 1 0 9 2
37 10 0 9 1 9 15 13 1 10 9 1 9 9 2 9 2 1 15 1 10 9 1 10 9 0 7 1 10 9 0 1 9 2 9 9 2 2
31 10 9 4 13 7 1 10 9 1 10 9 0 7 1 15 1 10 9 0 1 13 10 9 9 2 13 10 9 3 0 2
46 10 0 9 1 10 9 13 1 9 1 13 9 1 10 9 7 10 9 1 12 9 0 1 9 9 7 2 9 9 2 2 1 13 10 9 1 10 9 0 1 13 10 9 1 9 2
35 10 9 9 13 1 9 7 4 13 1 13 10 9 7 13 10 9 1 10 9 1 9 0 2 1 10 9 1 10 9 7 1 10 9 2
17 10 9 11 11 13 10 9 0 1 0 9 1 10 9 1 11 2
12 15 13 1 10 9 1 10 11 1 10 9 2
36 10 9 4 13 1 10 9 7 9 11 11 2 0 1 9 2 3 1 10 9 11 11 11 2 1 10 0 9 1 11 1 10 11 1 11 2
23 15 13 1 10 11 3 10 0 9 1 9 1 10 11 1 11 2 0 1 11 11 11 2
21 10 9 1 10 9 4 13 0 9 1 10 9 13 1 10 9 1 10 9 11 2
25 10 9 4 13 1 10 0 9 1 9 0 2 1 10 9 1 10 15 15 13 10 9 1 9 2
13 1 10 9 13 12 9 1 9 13 1 10 9 2
15 1 10 9 1 10 9 4 13 12 9 13 1 9 0 2
35 10 9 13 10 9 13 1 9 1 9 1 10 9 1 13 10 9 1 9 2 7 4 13 1 9 0 15 13 15 12 9 1 0 9 2
46 12 9 13 1 9 2 1 9 3 0 2 1 10 9 3 13 7 0 2 7 0 1 9 7 9 2 2 13 0 3 1 10 0 9 1 10 11 2 10 9 11 7 1 10 9 2
33 1 9 10 9 15 13 2 1 10 0 9 2 1 10 9 0 2 7 4 3 13 1 10 9 1 10 9 1 9 1 10 9 2
43 1 10 9 1 10 9 1 10 9 1 11 10 9 4 3 13 2 1 10 9 1 10 9 1 10 11 1 10 9 2 7 3 1 10 9 4 4 13 10 9 0 0 2
57 1 10 12 10 9 0 4 4 13 1 10 9 0 2 13 1 10 9 0 2 1 10 0 9 1 10 9 1 9 1 10 9 1 10 9 0 2 10 9 1 9 0 1 10 9 1 10 9 7 10 9 1 10 9 0 0 2
39 10 9 1 10 9 15 13 3 1 10 9 1 11 2 3 15 13 1 10 11 7 13 3 1 10 9 1 10 9 1 10 11 1 10 9 1 10 9 2
8 10 9 11 15 4 3 13 2
17 4 13 1 10 0 9 1 10 9 1 11 2 3 3 15 13 2
29 10 9 1 11 13 10 0 9 15 15 13 1 10 9 0 1 10 0 9 7 15 13 1 10 9 10 9 0 2
63 13 10 12 9 12 1 10 9 1 10 9 1 11 1 10 9 0 13 1 3 12 9 13 1 11 7 10 9 0 2 13 1 9 7 9 7 0 1 3 12 9 2 13 1 10 9 0 11 7 1 10 9 1 10 9 0 2 10 9 11 11 11 2
26 11 2 10 0 9 1 11 1 11 1 10 9 0 2 15 13 1 11 2 3 1 12 9 1 11 2
25 10 9 1 11 4 13 1 10 0 9 1 10 9 0 13 1 10 9 11 11 11 11 1 11 2
38 1 10 0 9 1 9 15 3 13 9 2 11 4 13 1 13 10 9 0 11 2 15 15 13 0 1 10 9 1 11 2 3 16 13 10 9 0 2
24 10 12 9 11 4 13 1 13 15 3 1 13 2 13 1 11 10 9 1 10 9 0 11 2
8 11 13 9 1 10 9 0 2
44 10 10 9 13 3 0 1 10 0 9 2 10 10 9 1 9 15 4 13 3 7 3 3 4 13 15 1 10 9 1 10 11 13 9 0 1 10 10 9 0 1 10 9 2
53 11 1 10 9 1 13 1 10 9 10 9 1 9 13 13 1 10 15 16 10 10 9 13 0 2 13 15 3 0 1 10 9 0 7 13 13 1 10 10 9 10 9 1 10 11 2 15 13 10 9 1 9 2
19 13 10 9 1 13 10 9 13 10 9 0 15 11 4 3 13 3 0 2
33 10 9 4 13 10 0 9 1 10 10 9 1 10 9 0 0 7 10 10 9 15 13 1 9 3 13 0 10 0 9 1 9 2
29 10 9 4 13 3 10 9 0 1 3 13 1 10 9 15 13 1 11 2 9 0 7 0 9 1 9 1 11 2
46 13 10 9 1 10 9 13 10 9 4 3 13 1 0 9 0 10 9 15 11 3 13 1 13 3 2 13 15 10 9 1 10 9 13 1 12 9 2 1 10 9 1 10 9 11 2
22 10 9 1 11 4 13 1 10 0 9 7 2 1 10 0 9 2 4 13 1 9 2
26 1 10 9 13 2 10 12 9 1 10 9 4 13 3 7 3 3 13 1 13 15 3 1 13 3 2
43 3 3 11 13 9 1 13 10 9 0 13 1 10 9 1 11 7 1 10 9 0 1 11 2 13 1 10 10 9 1 13 10 9 1 10 9 1 9 1 15 4 13 2
14 10 9 0 7 0 13 1 10 9 0 1 10 9 2
15 1 10 9 1 10 9 10 9 0 13 0 1 10 9 2
21 12 12 1 9 2 9 7 9 0 1 10 3 12 12 1 10 9 0 2 0 2
33 1 9 1 10 9 10 9 15 13 1 10 11 7 10 9 4 13 1 13 10 12 9 10 9 1 11 13 10 9 1 10 9 2
44 10 9 1 11 4 3 13 9 1 10 12 9 16 15 13 9 0 1 10 10 9 10 9 11 0 2 10 9 11 0 1 11 2 7 10 9 1 10 0 0 9 11 0 2
72 3 10 9 1 11 2 13 1 9 1 10 9 0 2 4 13 10 9 0 1 10 9 0 1 11 11 2 7 1 10 9 1 9 7 1 9 0 1 10 9 7 1 9 1 10 0 9 13 1 10 9 0 7 0 2 1 10 9 7 1 10 9 1 9 0 0 1 15 1 10 9 2
9 10 9 13 10 9 1 9 0 2
20 10 9 13 1 9 1 10 12 9 0 9 2 9 2 7 9 2 9 2 2
24 16 4 13 10 9 2 15 4 13 1 10 0 9 0 2 13 3 3 1 9 1 9 0 2
48 3 10 9 4 13 3 1 13 10 9 0 15 15 13 1 9 0 1 10 9 7 1 10 9 1 10 9 0 1 10 9 2 3 1 9 1 9 1 9 7 1 9 0 1 10 0 9 2
21 1 10 9 0 1 10 0 9 1 11 4 13 10 0 9 1 10 9 1 9 2
17 10 9 13 1 10 10 9 7 10 9 15 13 1 10 9 0 2
18 10 9 13 0 1 9 2 15 1 10 9 13 9 0 7 9 0 2
26 15 15 13 3 1 10 9 0 13 9 0 7 9 0 2 9 0 1 10 9 1 10 9 0 2 2
17 3 2 1 10 10 9 2 13 1 9 1 13 3 9 7 9 2
34 10 9 1 9 0 4 3 13 9 0 7 9 1 11 16 3 0 1 9 7 3 0 1 10 9 1 9 0 7 0 2 1 11 2
14 1 10 9 1 9 0 2 10 9 4 13 9 13 2
18 3 10 9 1 9 0 15 13 3 3 7 1 9 1 9 3 0 2
15 10 9 7 10 9 0 13 3 1 9 3 0 10 9 2
17 1 10 9 2 1 10 11 2 10 9 4 3 1 10 15 13 2
15 0 9 2 1 10 9 2 13 9 2 7 1 9 0 2
7 10 9 3 4 3 13 2
33 1 15 13 10 9 1 9 2 4 4 13 10 0 9 1 13 10 9 1 9 1 10 9 1 0 2 1 0 9 7 9 2 2
22 9 0 4 13 16 10 9 1 10 9 0 4 13 1 10 9 1 9 1 10 9 2
41 10 9 4 13 1 13 10 9 1 10 9 0 1 10 12 9 1 11 7 5 7 9 1 9 2 1 10 1 3 1 10 15 3 15 13 9 0 1 10 9 2
56 10 9 0 1 10 9 4 13 16 10 3 0 9 1 9 13 1 9 1 10 9 1 10 9 1 9 1 10 9 0 13 1 10 9 0 1 10 12 9 1 12 9 5 11 1 11 13 1 12 9 5 11 1 9 0 2
23 10 9 2 9 0 2 13 10 9 1 9 15 13 9 2 9 1 9 7 9 0 0 2
14 0 1 10 9 1 10 9 13 10 9 1 9 0 2
27 10 9 0 13 10 0 9 1 10 9 15 15 13 1 10 9 13 1 9 0 1 9 7 1 0 9 2
25 10 9 0 15 13 1 10 0 9 1 9 0 2 0 15 4 13 9 1 10 9 7 9 0 2
35 0 9 1 10 9 13 0 9 1 10 9 2 9 1 10 9 1 9 2 7 1 10 9 2 0 9 1 10 9 7 1 10 9 2 2
49 10 9 1 9 2 11 2 7 10 9 0 0 2 11 2 2 13 1 10 9 1 10 9 0 7 0 2 13 1 1 10 0 9 1 9 0 13 1 10 9 0 0 1 10 9 1 10 9 2
29 10 15 13 1 10 9 1 9 2 11 2 2 9 2 11 2 2 9 2 11 2 2 9 7 9 1 0 9 2
39 10 0 9 15 4 3 13 1 10 10 0 9 15 13 1 10 9 2 9 1 10 9 2 9 13 1 10 9 1 10 9 1 0 9 1 9 1 9 2
40 10 9 15 13 10 9 0 13 9 0 1 10 9 0 2 1 10 9 7 3 1 10 9 2 3 13 1 9 1 13 10 9 0 1 10 10 0 9 0 2
14 1 10 9 1 9 0 2 10 9 4 13 9 13 2
47 10 9 0 13 3 0 1 9 2 16 1 9 1 10 9 13 1 10 9 0 1 10 9 1 9 0 1 9 2 3 3 15 13 10 9 1 9 1 10 9 2 0 9 1 10 9 2
55 3 13 3 3 0 10 9 13 1 10 0 9 1 0 9 1 9 3 16 15 4 13 10 9 1 10 15 15 13 10 9 1 10 9 1 10 9 0 1 9 1 10 9 1 10 9 1 10 9 2 11 2 12 2 2
11 10 9 0 13 3 0 3 1 15 0 2
32 9 0 13 1 9 1 9 1 3 12 9 5 11 2 13 1 9 7 9 9 1 9 1 10 9 2 9 2 9 1 9 2
21 10 9 13 1 10 9 1 9 13 1 10 9 1 10 9 7 1 10 9 0 2
21 10 0 9 4 4 13 1 10 9 1 9 0 1 10 9 2 11 2 12 2 2
19 10 9 1 10 9 13 0 2 1 10 9 1 10 9 3 1 10 9 2
48 10 9 1 9 2 3 13 1 11 2 8 8 8 8 8 12 8 2 2 1 10 1 3 1 10 15 15 13 9 0 0 1 10 9 0 2 13 1 12 9 5 3 2 13 1 12 9 2
42 10 9 1 9 1 10 15 15 13 9 1 9 1 10 9 3 0 13 1 12 9 5 9 1 9 13 1 10 12 9 1 10 9 0 2 11 7 15 2 12 2 2
33 10 9 1 10 9 0 1 10 9 0 7 10 9 0 4 4 3 13 2 11 2 12 2 1 10 9 1 9 0 1 9 0 2
47 10 9 13 1 13 10 9 9 2 16 13 1 10 9 1 10 0 9 9 2 1 10 9 0 7 10 9 0 2 9 1 11 2 2 10 9 1 9 7 15 2 9 1 11 11 2 2
29 10 9 0 4 13 3 1 10 9 1 9 2 11 2 7 2 1 9 0 2 1 10 9 1 9 2 11 2 2
24 15 4 13 16 10 9 13 3 0 1 10 9 2 1 10 15 13 1 10 9 3 7 3 2
58 16 3 13 1 9 1 9 1 9 2 10 9 4 13 15 1 10 9 1 9 0 13 1 10 9 1 10 9 2 1 9 7 9 2 2 1 10 9 1 9 1 9 1 10 9 13 7 1 10 9 0 7 0 1 10 9 0 2
24 1 10 9 10 9 0 1 11 7 1 11 13 3 1 10 9 1 10 0 9 1 10 9 2
9 10 9 4 13 1 10 0 9 2
67 1 9 4 4 13 1 10 9 11 11 2 1 10 0 7 10 0 2 1 10 9 0 1 10 9 1 9 0 1 10 9 0 2 9 1 10 9 9 0 13 1 10 12 1 11 11 11 2 0 2 9 12 2 12 2 2 10 9 9 2 0 3 1 9 7 9 2
35 9 13 1 11 2 9 1 9 0 7 0 7 1 9 1 9 0 13 15 3 1 9 0 15 13 1 9 1 9 2 9 0 2 2 2
42 10 9 11 2 11 2 11 2 8 2 13 10 9 0 0 1 11 2 1 9 0 2 13 7 13 1 10 9 11 11 11 11 2 13 9 1 10 9 11 11 2 2
41 1 10 10 3 12 9 1 9 1 10 9 2 3 15 1 10 0 9 1 9 1 11 11 2 2 10 11 15 13 1 15 1 10 9 0 3 0 1 10 9 2
44 10 9 1 10 11 13 1 9 1 10 9 1 11 7 13 10 9 3 1 10 9 1 10 9 2 13 0 9 1 10 0 9 1 10 9 1 11 2 15 13 15 1 12 2
20 10 9 1 10 11 13 3 0 1 9 1 10 10 0 9 0 1 9 0 2
19 1 10 9 10 9 13 10 9 3 1 10 9 0 1 10 9 1 11 2
21 10 9 4 13 1 0 9 7 15 13 1 10 9 1 13 1 10 10 9 3 2
14 15 1 10 12 9 4 13 1 10 0 9 1 9 2
39 10 0 9 13 1 10 12 1 10 9 2 10 0 9 4 13 1 10 12 1 9 7 13 3 0 16 10 9 15 13 16 4 13 10 10 9 1 9 2
34 1 10 9 1 9 15 13 9 10 12 9 12 9 1 10 10 9 2 10 0 9 13 10 9 15 13 1 10 12 1 10 12 9 2
38 10 9 4 13 1 9 13 7 1 0 9 9 1 12 9 2 13 1 9 0 1 9 1 10 9 2 15 13 10 9 1 9 1 9 7 9 0 2
47 1 10 9 13 0 10 9 1 10 9 15 13 10 9 1 10 9 2 10 9 1 15 15 13 1 13 1 10 9 13 2 10 0 9 7 10 9 1 10 9 1 15 15 13 10 9 2
42 15 1 10 9 13 10 9 0 2 1 9 7 9 2 1 10 9 2 3 3 3 1 10 9 15 4 13 1 10 9 15 13 10 9 1 10 0 9 1 10 9 2
14 10 9 3 0 1 10 9 13 10 9 11 2 11 2
21 11 13 10 9 3 0 1 10 9 2 7 11 10 0 1 9 1 10 10 11 2
24 10 9 1 10 9 13 9 1 9 9 11 13 1 12 9 13 3 1 13 1 10 9 12 2
26 10 9 4 13 10 0 9 9 12 2 15 4 13 1 10 12 7 13 3 1 10 9 1 10 12 2
17 1 9 10 9 4 13 1 9 9 12 15 4 13 1 10 12 2
42 10 9 11 13 9 1 10 12 2 1 9 1 10 9 1 10 9 1 10 11 2 1 10 9 1 10 9 1 10 11 11 1 10 9 1 11 7 10 9 1 11 2
21 10 12 9 4 13 1 10 12 1 10 9 1 10 9 1 9 13 10 9 11 2
55 1 10 9 1 10 9 1 10 12 9 10 9 3 13 0 7 1 15 10 9 4 13 1 10 9 1 10 11 11 11 7 10 9 11 2 11 2 13 1 11 1 10 9 1 11 1 3 13 10 9 11 3 1 11 2
30 1 10 9 13 1 10 0 9 0 10 9 1 10 9 3 13 16 0 9 0 13 10 11 1 13 1 10 9 0 2
22 10 9 13 1 10 9 1 0 9 0 3 1 10 9 13 1 9 1 10 9 0 2
49 10 11 11 13 1 13 10 9 0 1 10 12 2 16 4 13 10 9 1 9 1 10 9 11 2 11 7 4 13 1 10 10 9 0 1 10 9 1 9 1 10 9 2 1 11 7 11 2 2
29 1 15 10 11 13 1 13 3 10 9 1 10 9 11 2 11 2 3 1 10 9 1 9 1 10 9 0 0 2
25 1 10 12 4 13 1 10 9 0 1 10 9 11 2 11 7 1 15 10 11 13 1 13 15 2
30 1 10 12 2 1 9 1 10 9 1 10 9 9 1 10 9 2 4 13 1 13 10 9 1 9 1 10 9 11 2
29 1 13 9 1 10 9 1 10 11 11 1 13 10 10 9 13 4 13 3 10 11 11 7 10 11 11 2 11 2
26 1 10 12 2 10 11 11 13 10 9 1 12 9 1 9 10 9 2 3 12 9 1 9 10 9 2
13 10 9 15 13 10 9 0 3 0 1 10 9 2
36 2 11 2 3 13 2 1 10 9 2 1 10 9 1 10 9 2 2 7 13 10 9 13 1 13 10 9 1 9 1 15 0 1 10 9 2
31 10 9 13 3 1 10 12 9 0 8 2 9 2 2 8 9 9 2 11 2 9 2 2 7 2 9 1 10 9 2 2
26 11 4 4 13 3 9 2 1 1 9 2 11 11 2 15 13 0 1 10 9 9 1 10 9 11 2
18 3 10 9 11 2 9 1 11 7 10 9 11 1 11 13 10 9 2
35 1 10 0 9 0 2 10 9 0 1 10 9 0 13 16 10 9 1 10 10 9 4 13 2 7 10 11 4 13 1 2 9 9 2 2
52 13 10 10 9 3 1 10 12 2 16 10 9 0 0 13 1 13 10 0 9 1 2 11 2 2 15 1 13 1 13 9 1 10 9 1 11 1 10 11 11 1 11 2 1 10 0 9 1 10 9 11 2
17 10 9 1 10 9 3 13 1 13 15 3 1 2 11 11 2 2
81 10 0 9 0 4 13 1 10 9 0 1 10 11 9 1 9 1 9 7 9 1 11 11 2 10 9 13 10 10 9 1 10 9 1 10 9 1 11 1 10 11 2 2 11 2 10 9 13 15 1 10 9 0 15 13 10 9 1 10 9 2 7 11 11 2 10 9 15 13 1 10 11 1 13 15 1 10 10 9 2 2
43 10 9 1 9 4 3 13 3 10 9 1 10 11 9 1 10 0 9 1 9 1 9 1 9 11 2 1 9 7 9 0 2 7 11 11 11 2 2 1 9 9 2 2
47 10 9 13 10 9 1 10 9 0 0 15 2 1 10 9 1 10 11 11 12 10 12 9 12 2 13 10 11 1 13 10 0 9 1 13 10 9 0 1 9 1 11 11 7 11 11 2
45 10 9 13 1 10 9 13 10 11 1 10 11 7 10 9 1 9 0 2 11 2 2 3 0 1 9 1 9 9 11 11 2 1 10 9 1 10 9 1 11 2 10 9 2 2
31 9 7 9 1 10 9 13 10 9 11 11 10 15 13 1 13 10 9 0 1 10 9 2 11 2 7 10 9 0 0 2
72 10 9 13 10 9 1 10 9 1 9 1 10 9 1 9 1 10 11 1 10 9 9 11 2 10 9 1 10 9 11 11 2 10 10 9 1 12 9 2 10 9 1 10 9 0 2 10 9 1 10 9 13 1 11 11 1 11 2 10 9 1 9 7 3 10 9 1 9 1 10 9 2
22 10 9 1 10 11 1 10 9 1 10 9 0 15 13 3 1 13 1 10 9 12 2
50 1 10 12 2 12 9 1 10 9 1 10 0 9 1 9 0 1 11 2 10 9 0 1 10 9 0 13 1 11 11 10 9 1 13 0 9 1 10 9 1 13 3 10 9 1 10 9 0 0 2
25 11 13 1 10 9 1 9 2 9 1 9 2 1 10 15 4 13 10 9 0 11 13 10 9 2
69 1 10 9 1 9 1 10 0 9 3 1 10 9 1 11 1 10 9 1 10 11 0 2 11 2 2 11 13 9 1 13 1 10 9 2 3 3 2 3 1 10 9 1 10 11 13 10 15 1 13 1 10 9 1 10 9 9 7 10 9 1 10 9 0 1 10 10 9 2
53 10 12 9 12 2 10 9 0 13 3 10 9 0 0 2 1 9 13 1 9 11 11 2 13 1 11 11 2 1 9 1 9 1 10 9 1 10 9 0 2 11 2 2 7 1 11 11 2 9 1 10 11 2
21 10 9 1 10 9 13 1 11 1 13 1 10 11 10 9 1 13 10 0 9 2
15 1 10 9 1 10 12 10 9 0 13 10 10 9 0 2
55 9 7 9 1 10 9 3 13 10 9 11 11 1 10 15 13 1 13 10 9 1 10 9 1 10 9 1 10 9 9 1 10 9 2 11 2 7 1 10 9 0 0 2 1 10 15 13 1 9 1 10 9 1 9 2
55 10 9 15 1 10 0 9 13 10 9 1 9 1 10 12 9 1 9 0 4 13 1 11 10 12 9 12 1 10 9 1 10 9 0 0 1 10 11 2 10 9 11 11 2 7 1 10 11 2 10 9 11 11 11 2
13 10 9 1 9 13 10 9 1 9 1 12 9 2
59 10 0 13 10 9 1 10 9 0 1 10 9 2 10 0 9 4 13 10 9 1 9 1 10 9 0 1 10 9 1 11 11 7 1 10 0 9 4 4 13 10 9 0 1 10 9 0 1 10 9 1 10 0 9 7 1 10 9 2
32 10 9 1 10 9 13 1 10 0 9 1 10 9 15 15 13 1 13 3 10 9 13 7 1 3 13 15 10 9 1 9 2
38 10 9 3 2 1 3 3 13 1 10 9 0 7 0 2 4 4 13 10 0 9 1 10 9 1 10 9 0 7 1 10 9 1 9 1 10 11 2
35 10 9 0 1 10 9 13 10 12 9 12 1 11 16 10 3 9 1 10 9 0 11 11 7 10 0 9 0 11 11 11 13 10 9 2
34 13 10 9 0 1 10 9 1 10 9 10 9 0 13 10 9 0 9 12 1 10 9 1 12 9 1 9 1 13 15 1 12 9 2
22 1 10 9 1 10 9 1 10 9 0 7 0 13 9 10 9 1 10 9 0 0 2
85 13 3 12 10 9 7 9 1 4 13 1 10 11 1 10 12 7 10 12 1 10 11 9 9 9 2 11 2 2 10 11 9 9 2 11 2 2 10 9 11 2 11 2 11 2 11 2 7 10 9 1 10 11 1 11 11 1 10 9 1 13 15 1 10 9 1 10 9 2 1 10 9 7 9 1 10 9 9 7 1 10 9 1 9 2
34 1 10 0 9 1 10 12 10 11 13 1 10 9 1 10 9 10 9 1 9 0 7 0 1 10 9 1 9 7 9 1 10 9 2
15 10 9 1 9 11 4 13 1 10 9 1 9 15 13 2
73 10 9 13 1 10 9 1 12 9 1 9 2 10 9 0 7 10 9 1 9 1 9 1 13 12 2 12 11 2 10 9 0 0 1 13 9 3 1 12 9 1 9 0 1 10 12 7 10 12 9 7 3 9 0 1 0 7 0 1 10 9 0 7 0 1 10 9 7 1 10 10 9 2
37 10 11 13 1 10 0 9 12 9 9 7 12 1 15 4 13 1 9 9 1 10 11 9 9 1 9 0 3 10 12 9 7 10 12 9 12 2
35 10 9 13 2 1 10 9 0 13 1 10 0 9 2 13 1 13 10 9 1 10 9 1 10 9 1 10 12 7 10 12 9 1 9 2
21 10 0 9 4 13 0 10 9 1 10 9 0 1 10 0 9 0 1 10 11 2
34 1 10 9 1 10 12 3 10 0 11 13 1 11 13 10 9 1 10 9 1 9 11 11 13 10 9 0 13 1 9 1 10 11 2
42 10 9 13 10 9 1 9 11 11 2 1 9 1 10 9 1 10 9 2 7 10 9 11 1 10 15 4 13 10 9 0 1 10 9 1 10 9 7 1 10 9 2
51 10 9 1 10 9 1 9 13 1 10 12 9 7 10 12 9 12 1 9 1 9 9 11 11 13 1 11 15 13 3 1 13 10 9 1 10 9 1 9 7 1 15 1 10 9 1 9 1 10 9 2
41 10 9 1 13 9 9 11 4 13 1 10 11 3 0 1 10 9 13 1 10 10 9 7 9 9 1 10 9 1 9 2 9 1 9 2 13 3 1 10 12 2
26 10 0 7 10 0 9 3 13 1 9 3 10 9 1 10 9 1 10 9 1 10 9 1 0 9 2
58 10 0 9 1 10 9 13 10 10 9 10 12 9 12 1 10 12 11 16 4 13 1 9 10 11 11 12 1 10 9 1 10 11 1 11 11 1 10 9 0 7 4 13 1 9 1 10 9 1 12 9 7 10 9 1 12 9 2
22 10 11 11 13 3 10 0 9 1 4 3 13 7 13 1 10 9 1 10 11 0 2
20 10 9 15 13 1 10 9 1 12 9 1 9 7 13 3 15 1 12 9 2
54 10 9 1 10 9 13 10 9 1 10 9 0 1 10 12 7 10 12 9 1 9 7 10 9 1 9 1 10 9 0 13 1 9 1 10 9 9 1 11 13 1 10 9 11 11 2 9 1 11 11 1 10 11 2
44 10 9 1 9 1 10 11 13 1 10 9 11 11 15 13 10 9 12 1 13 10 13 9 1 10 9 13 7 13 16 15 4 4 13 1 0 9 7 10 0 9 1 9 2
53 9 13 10 9 0 0 1 10 9 1 10 9 0 1 10 0 9 1 10 11 13 15 1 11 11 1 10 9 1 10 12 7 10 9 0 4 13 0 10 9 1 10 12 1 11 1 10 9 1 10 11 0 2
29 10 9 1 10 9 7 10 9 0 3 3 13 0 1 13 10 9 1 9 0 1 10 9 7 1 10 9 0 2
48 1 9 3 1 10 9 13 1 10 11 2 1 10 11 7 1 10 9 0 1 10 9 0 1 10 9 1 10 9 12 2 10 9 11 11 13 1 13 15 3 1 10 9 1 10 10 9 2
35 10 9 13 11 1 13 1 13 1 10 9 0 10 9 0 1 10 11 2 15 1 10 9 13 10 9 0 1 10 9 0 1 10 9 2
80 1 10 9 13 16 10 9 0 1 10 12 5 1 10 9 1 10 11 4 13 1 10 9 0 2 3 3 1 10 0 9 11 11 2 2 7 13 10 0 9 1 9 1 10 9 0 2 3 1 9 1 11 7 0 9 9 1 10 9 0 0 2 11 2 3 13 1 10 9 1 10 9 11 12 7 12 1 10 11 2
43 3 13 9 1 10 10 9 11 7 0 9 1 10 11 13 1 13 1 10 9 9 0 15 3 13 9 1 10 11 7 3 4 13 1 10 11 13 10 9 0 3 0 2
30 1 10 0 9 1 10 9 4 13 3 10 9 1 10 9 0 1 11 7 10 9 1 10 9 1 9 1 10 9 2
34 10 9 1 10 9 1 10 11 11 12 1 10 9 1 10 0 9 13 1 13 1 10 9 1 10 9 11 11 7 1 10 10 9 2
44 10 11 7 10 11 13 10 9 0 1 10 0 9 1 10 12 16 10 11 13 1 10 9 1 10 9 1 9 1 10 11 1 10 9 11 11 0 7 10 9 0 1 9 2
30 10 12 9 12 9 11 0 13 10 9 1 10 9 13 15 1 10 9 11 11 2 1 10 9 7 9 1 10 11 2
54 10 9 0 4 3 4 13 1 11 13 10 9 1 9 1 11 11 2 9 9 1 10 10 9 0 7 1 10 9 7 10 9 0 1 10 9 13 3 3 10 9 1 10 9 0 1 10 9 7 1 10 10 9 2
59 1 10 9 1 10 9 1 9 1 11 4 13 10 0 9 11 11 2 3 13 1 10 9 0 7 13 1 10 9 1 9 1 10 9 1 10 11 2 1 10 9 1 3 12 9 1 10 11 11 1 10 15 4 13 10 9 1 9 2
46 10 9 0 1 10 9 7 1 10 9 1 10 9 4 13 1 10 9 0 1 10 9 9 12 1 10 9 0 1 12 9 1 9 1 13 15 3 1 10 9 1 10 9 11 11 2
31 9 13 3 10 9 1 10 9 1 10 9 1 10 11 1 10 9 1 11 13 3 16 10 15 13 3 1 10 10 9 2
26 1 9 1 15 2 11 13 3 10 9 1 10 11 1 10 9 1 9 0 0 1 10 9 11 11 2
33 1 10 9 1 9 12 10 9 1 10 9 9 7 1 10 9 11 11 12 4 13 7 15 13 1 10 9 0 3 1 10 9 2
50 10 12 9 1 10 9 12 11 10 9 0 1 10 11 13 10 11 11 12 1 10 9 9 11 11 2 13 1 9 1 10 11 9 9 2 1 10 9 1 11 11 2 1 10 11 7 1 10 11 2
25 10 9 13 1 9 1 9 0 0 2 13 1 10 9 1 12 9 7 1 10 9 1 12 9 2
28 10 9 13 9 1 10 9 1 0 9 1 10 9 0 7 1 10 9 1 10 9 1 9 1 10 9 0 2
16 10 10 9 13 1 9 3 10 12 9 7 10 12 9 12 2
28 10 9 13 3 0 3 1 10 10 9 2 13 10 12 9 12 1 12 9 1 9 1 10 9 7 12 9 2
40 1 10 9 1 10 12 2 11 2 3 3 16 4 13 10 9 1 10 9 13 1 10 9 2 13 10 9 0 1 10 0 9 1 10 11 13 15 1 11 2
69 10 12 9 12 3 2 10 9 1 10 9 1 10 9 1 11 11 11 11 7 10 9 1 10 11 11 11 13 10 9 1 9 15 13 10 9 1 9 1 10 15 4 4 13 10 9 1 9 1 9 1 10 9 1 9 7 9 13 1 9 11 1 10 9 1 9 11 11 2
11 10 9 13 10 9 0 1 10 10 9 2
39 10 9 1 10 11 11 2 11 11 2 13 10 9 10 12 9 12 7 10 9 0 13 10 10 9 10 12 9 1 10 0 9 1 10 9 11 11 11 2
24 10 9 0 3 13 10 0 9 1 9 0 1 10 15 10 11 11 13 10 9 1 10 9 2
18 3 10 9 4 13 1 10 9 0 1 10 9 1 10 9 11 11 2
50 13 10 9 1 10 11 2 11 13 1 10 9 0 13 1 10 11 7 13 3 10 9 1 11 7 10 10 9 2 10 15 13 10 10 9 1 10 11 7 13 10 9 1 15 13 1 10 10 9 2
21 3 0 13 3 10 9 1 10 9 15 13 10 9 1 10 11 1 10 9 0 2
37 13 10 0 9 1 10 9 1 10 11 11 12 1 10 9 0 1 10 12 2 10 9 13 1 10 9 0 15 13 1 10 9 1 10 0 9 2
51 10 9 0 1 10 9 13 1 13 15 1 10 9 0 15 13 10 11 1 10 9 12 2 13 1 10 9 0 1 10 12 2 7 1 10 9 0 15 3 13 1 10 9 1 10 9 10 10 9 0 2
65 10 9 9 12 1 10 12 9 12 15 13 12 9 1 10 12 9 1 9 13 1 9 1 10 9 0 1 10 9 0 0 13 10 9 1 10 9 0 7 16 4 13 1 10 9 12 2 12 2 4 13 1 13 9 3 1 10 9 1 10 9 12 7 12 2
42 11 3 13 0 10 9 1 10 9 0 3 1 10 12 7 10 12 9 1 10 9 1 9 1 9 1 9 1 11 11 7 11 11 7 10 9 1 10 9 9 0 2
42 10 9 3 13 1 10 11 12 2 13 11 2 9 2 1 13 10 9 1 10 11 13 1 10 9 1 10 9 2 13 9 1 10 0 9 1 9 1 11 7 11 2
24 10 9 3 4 13 1 10 9 1 10 9 0 1 10 9 11 11 1 10 9 1 9 9 2
37 11 1 10 0 9 13 10 9 7 10 9 1 10 9 1 9 1 9 1 9 9 13 3 10 9 1 13 15 10 9 7 10 9 1 10 9 2
26 1 10 9 10 9 11 11 13 1 10 9 1 10 9 11 11 12 10 12 9 12 1 10 12 11 2
24 10 9 0 1 10 9 0 4 13 2 1 10 0 9 2 1 12 0 9 1 10 11 11 2
55 10 0 13 10 9 1 13 10 9 0 1 10 0 9 7 4 13 1 10 11 7 10 0 9 2 13 1 10 9 1 10 11 7 10 9 1 10 11 2 4 13 1 13 15 10 9 7 10 9 1 10 9 1 9 2
22 13 10 9 13 13 0 13 3 10 9 0 1 10 9 1 10 12 7 10 12 9 2
45 10 9 3 13 1 13 10 0 9 1 9 7 10 11 11 12 15 4 13 10 12 9 12 1 10 12 11 13 10 9 3 13 1 10 11 11 12 7 3 13 1 9 3 0 2
40 1 10 11 11 12 2 10 9 13 10 11 11 1 10 9 15 13 1 10 9 1 10 9 11 12 1 10 9 9 11 1 9 1 9 0 10 12 9 12 2
18 10 12 13 13 10 9 1 9 0 1 10 9 0 1 10 9 0 2
50 10 9 9 12 1 10 12 9 7 10 9 9 12 1 10 12 9 12 3 13 1 10 9 1 10 9 1 10 9 0 7 0 10 9 1 13 1 10 9 10 9 1 10 9 1 10 9 0 0 2
40 1 10 9 13 0 10 9 1 0 9 1 10 9 11 11 3 1 9 0 3 0 3 1 10 9 1 10 9 13 1 10 9 0 1 10 0 9 9 12 2
26 10 9 2 10 9 2 3 13 9 1 12 9 1 9 1 10 9 1 10 9 13 1 12 9 0 2
18 10 12 9 12 4 13 1 9 10 9 0 11 12 13 1 10 11 2
20 10 10 9 13 1 9 10 9 1 10 9 0 1 10 9 0 1 9 9 2
50 15 1 10 11 12 3 13 10 0 9 13 1 10 9 0 0 2 15 13 3 0 1 13 1 10 9 1 10 12 1 9 1 10 9 1 10 9 0 1 10 3 0 9 11 13 1 10 9 0 2
48 1 10 9 1 10 12 9 1 15 4 13 10 9 1 10 9 9 12 2 10 11 13 10 9 1 12 9 1 9 13 1 10 10 9 1 10 9 12 13 15 12 9 1 10 9 11 11 2
41 1 10 9 1 10 9 1 9 1 10 9 0 0 1 10 9 1 10 9 2 10 9 0 1 10 9 3 13 10 9 1 10 9 1 10 9 7 1 10 9 2
31 1 10 12 10 9 9 0 15 13 1 10 9 1 10 9 0 11 11 11 15 13 0 10 9 1 10 11 7 10 11 2
19 10 9 1 9 1 10 12 9 13 9 0 1 15 13 1 10 9 0 2
20 10 9 1 10 9 13 10 9 1 12 9 7 10 10 9 1 12 9 0 2
28 10 9 13 10 9 1 10 9 1 10 9 0 7 10 9 0 1 10 9 0 15 13 10 9 7 10 9 2
14 1 10 12 10 9 11 11 13 3 10 9 1 9 2
31 1 10 9 0 0 3 1 10 9 11 11 4 13 1 13 1 10 12 9 12 9 9 1 10 9 3 1 13 10 9 2
21 10 9 1 9 13 12 11 11 2 12 11 2 11 2 11 7 12 11 2 11 2
16 3 10 9 0 13 10 9 1 10 3 11 11 11 5 11 2
37 10 10 9 13 10 12 9 12 1 10 12 11 1 10 9 11 11 1 10 9 11 7 13 10 9 0 1 9 1 12 9 7 9 1 12 9 2
33 10 10 9 0 13 3 1 9 1 10 9 1 9 7 9 2 11 2 1 10 9 0 2 15 13 1 13 1 12 9 1 9 2
20 10 9 3 13 1 10 9 10 12 9 1 10 0 9 1 12 9 1 9 2
15 10 0 9 4 13 1 10 10 9 1 12 9 1 9 2
34 1 10 12 10 9 0 2 10 9 7 10 9 13 15 1 10 9 11 11 13 1 10 0 9 1 10 9 2 10 9 2 1 11 2
8 10 9 1 11 9 11 11 2
21 10 10 9 13 0 1 10 9 9 0 1 10 9 1 10 9 1 9 11 12 2
16 10 9 4 13 1 9 1 9 2 11 2 13 1 9 0 2
15 10 10 9 13 10 9 0 2 10 9 7 10 9 0 2
41 1 10 9 13 10 10 9 2 10 9 1 9 2 1 9 1 10 11 2 13 10 9 13 1 10 9 7 1 10 9 1 10 9 1 10 9 11 11 1 11 2
27 1 15 15 13 10 9 1 10 9 1 9 2 9 7 9 1 9 0 1 9 1 9 7 1 9 0 2
44 10 9 1 9 3 2 3 3 0 1 10 9 1 9 9 2 4 4 13 1 10 9 1 9 1 10 9 1 9 13 1 10 11 0 3 1 10 9 7 13 1 9 0 2
49 0 9 13 10 9 1 10 9 1 9 1 10 9 7 10 9 1 9 9 1 10 9 0 0 1 10 9 0 7 3 10 9 1 10 9 0 13 1 10 9 1 10 9 0 2 0 7 0 2
27 3 2 16 10 9 1 9 3 4 3 13 1 10 9 1 9 1 10 12 2 13 1 9 12 0 9 2
21 10 0 13 10 9 1 13 9 7 9 1 10 9 1 9 7 9 13 1 9 2
27 10 0 3 15 13 1 10 9 1 10 9 1 9 0 1 10 9 0 7 0 1 9 1 10 9 0 2
43 10 0 9 13 10 9 1 13 7 13 10 9 1 9 0 1 10 9 1 13 10 9 1 10 9 0 1 10 9 1 9 1 9 1 9 7 10 9 1 10 9 0 2
37 10 0 9 13 10 9 1 10 9 11 2 9 0 1 9 9 9 2 7 13 13 1 9 0 9 1 10 9 0 1 10 9 0 1 9 0 2
32 10 0 9 13 1 10 9 1 10 9 1 9 1 10 9 1 10 9 1 9 13 1 9 9 1 10 9 1 10 9 0 2
32 10 0 9 13 13 10 9 1 9 1 10 9 1 9 1 10 11 11 11 3 1 9 1 10 9 0 7 0 1 10 15 2
26 10 9 13 10 9 0 13 1 10 9 1 10 11 0 2 9 2 13 1 3 10 12 5 1 9 2
26 1 10 10 9 0 2 10 9 13 10 9 0 1 10 9 0 15 13 1 10 12 1 10 12 9 2
13 10 10 9 15 13 1 10 12 1 10 12 9 2
7 10 9 13 10 9 0 2
19 10 9 1 9 0 1 10 9 1 10 0 9 4 13 1 12 1 12 2
16 10 9 13 10 9 0 2 15 13 1 10 9 0 7 0 2
12 1 9 1 9 10 9 15 13 13 15 3 2
13 4 13 3 1 9 2 16 13 13 9 0 0 2
19 10 9 1 10 9 4 13 1 10 9 0 1 10 9 2 13 3 9 2
41 1 13 15 10 9 2 13 2 15 13 1 13 1 10 9 1 9 1 9 2 7 2 1 9 3 0 2 15 13 1 10 9 1 10 9 0 7 1 0 9 2
19 10 9 15 13 1 15 10 9 15 13 7 15 13 2 13 3 10 9 2
33 10 9 4 3 13 13 2 3 9 1 10 9 1 9 1 9 13 0 2 13 1 9 7 3 2 15 13 7 13 10 9 0 2
20 10 9 0 13 10 9 2 15 13 1 10 13 10 9 0 7 13 10 9 2
31 15 13 3 1 10 9 0 2 15 4 13 1 10 9 1 13 10 9 0 1 10 9 0 7 13 2 15 13 10 9 2
40 9 0 2 15 13 1 9 0 2 0 1 10 9 1 9 0 2 9 9 2 1 9 7 9 2 9 0 15 15 13 1 9 0 2 9 0 1 9 0 2
31 10 9 1 9 4 13 1 10 9 1 9 1 10 9 2 9 2 9 2 9 2 7 1 10 9 0 7 0 7 0 2
18 13 10 9 0 10 9 13 10 9 13 2 9 0 15 13 10 9 2
19 9 1 9 4 13 1 10 9 1 9 9 7 1 0 9 1 9 13 2
25 1 10 9 1 9 4 4 13 9 1 9 2 15 13 1 10 9 0 9 7 0 9 1 9 2
36 10 9 13 10 9 0 0 15 15 13 1 10 9 1 9 2 9 7 10 9 1 9 2 2 9 2 9 2 9 2 7 10 9 1 9 2
22 15 15 13 1 10 9 1 9 2 7 9 10 9 2 15 1 10 9 13 1 9 2
12 10 9 15 15 13 1 13 4 13 9 0 2
20 10 0 9 1 13 10 9 13 15 1 13 15 1 10 9 1 10 9 0 2
13 10 9 3 13 10 9 13 1 10 9 1 9 2
9 15 13 1 10 9 1 9 13 2
27 10 9 2 15 4 13 1 10 9 0 2 10 9 2 13 9 1 10 12 7 10 12 9 7 9 0 2
28 10 9 13 1 10 9 9 2 9 2 9 7 0 9 0 1 9 2 1 9 1 10 9 13 1 10 9 2
9 0 3 10 9 1 10 9 0 2
45 10 9 4 13 2 3 2 1 10 12 1 10 12 9 2 1 3 1 10 9 1 10 9 9 7 1 10 9 1 10 9 2 7 1 10 12 1 10 9 1 12 9 1 9 2
36 10 9 1 9 1 10 9 4 13 1 10 9 2 15 13 10 9 1 10 9 1 10 9 2 1 9 2 7 10 10 9 2 1 9 2 2
13 1 10 9 0 13 2 3 2 10 9 3 0 2
24 1 10 9 0 4 13 10 9 1 10 9 1 10 9 2 10 0 9 7 10 9 1 9 2
16 1 3 10 9 3 13 10 9 7 4 13 13 10 10 9 2
15 10 9 13 10 9 0 1 10 9 7 13 1 0 9 2
25 10 0 9 13 16 10 9 13 1 10 9 13 3 0 1 10 0 9 1 10 0 9 1 9 2
12 10 9 13 1 10 9 1 10 9 10 9 2
19 10 0 9 15 15 13 1 10 0 9 4 13 3 1 10 12 9 11 2
11 1 12 9 11 13 10 0 7 0 9 2
11 1 12 9 11 15 13 10 9 1 9 2
21 3 10 9 4 13 13 1 0 9 1 13 9 3 1 10 9 1 12 9 11 2
13 10 9 4 13 1 10 9 1 10 9 1 9 2
36 10 9 13 3 0 1 10 9 7 2 13 2 13 10 9 0 1 10 9 13 3 1 10 9 1 0 9 0 15 2 16 13 2 15 13 2
8 10 9 4 13 3 1 9 2
38 15 4 13 1 10 9 16 10 9 13 10 9 0 2 7 15 13 1 10 9 1 9 1 9 0 2 16 15 13 1 10 9 1 9 1 9 0 2
14 3 10 9 1 10 9 13 10 0 13 10 9 0 2
32 1 10 0 9 1 10 9 10 10 9 4 13 3 1 10 9 7 1 0 9 1 9 0 2 3 1 10 9 0 7 0 2
32 10 0 9 1 9 1 9 0 1 10 12 13 13 10 11 2 13 1 11 11 2 9 0 2 11 2 11 2 11 7 11 2
36 1 10 10 9 2 10 9 4 13 3 1 10 9 2 7 13 3 9 1 10 9 1 10 9 1 9 7 1 10 9 2 9 7 9 2 2
10 3 4 13 1 10 9 0 7 0 2
13 3 3 2 10 9 4 13 1 9 1 0 9 2
43 15 15 4 13 1 10 9 2 1 9 1 0 9 2 1 9 7 9 2 1 10 9 1 9 0 2 1 10 9 2 1 9 0 2 1 9 0 1 13 9 1 9 2
35 3 2 1 9 1 10 9 2 1 9 1 10 9 2 15 4 13 1 13 10 9 1 9 1 9 2 1 13 9 7 9 1 10 9 2
26 10 9 3 4 13 3 0 1 10 12 9 5 9 7 10 9 1 10 9 3 0 1 10 12 9 2
18 10 9 3 0 13 10 0 9 15 15 13 13 10 9 1 9 0 2
32 10 9 13 10 9 0 0 15 13 10 9 1 10 9 0 2 13 3 10 9 0 2 1 15 4 3 13 2 9 0 2 2
26 4 4 13 1 13 9 1 9 3 0 15 13 1 10 9 1 10 9 15 13 10 9 1 10 9 2
30 10 9 4 13 1 10 12 1 10 9 0 9 11 11 1 11 2 15 15 13 1 10 11 11 1 11 1 10 12 2
29 13 3 9 0 7 1 10 12 9 2 10 9 4 13 1 13 1 10 9 1 9 0 1 10 9 7 3 0 2
24 10 9 2 1 10 0 9 7 9 2 13 3 10 12 5 1 10 9 0 13 1 10 9 2
36 4 13 1 13 1 10 9 1 9 1 10 9 2 7 3 1 10 9 2 1 10 9 2 3 2 13 1 10 9 1 9 0 2 11 2 2
24 4 3 13 9 1 9 2 11 2 7 15 13 9 1 9 15 4 3 13 1 0 9 0 2
6 10 9 0 13 13 2
20 10 9 15 13 1 10 9 13 10 9 0 15 4 13 1 10 9 1 9 2
33 1 9 10 9 4 13 1 9 1 10 9 7 3 10 9 13 7 13 1 0 9 1 9 13 0 1 10 9 0 1 10 9 2
21 13 13 10 9 1 10 0 9 13 1 10 9 1 9 0 15 4 13 10 9 2
29 10 9 2 1 9 13 2 1 10 9 15 13 1 9 3 0 1 10 9 2 7 1 9 13 2 1 9 2 2
19 1 9 1 9 1 9 2 9 0 2 0 2 10 9 13 10 9 0 2
2 9 12
2 12 2
36 10 9 1 10 9 15 13 13 1 10 9 7 1 10 9 1 10 9 2 10 9 7 10 10 0 9 0 1 10 9 3 4 13 9 0 2
2 12 2
32 16 4 13 1 9 1 10 9 10 9 2 15 4 13 1 9 0 2 0 7 13 10 9 2 7 10 9 0 1 15 13 2
17 9 2 10 9 2 10 9 2 10 9 7 10 9 1 9 13 2
50 9 2 10 9 1 9 7 10 9 1 9 2 10 9 2 10 9 7 10 9 1 9 7 10 9 0 1 10 15 2 10 10 9 7 9 0 1 10 9 1 10 9 1 10 11 9 1 9 0 2
10 9 2 10 9 13 2 9 9 2 2
5 9 2 10 9 2
43 9 2 10 9 1 9 0 13 10 9 0 1 10 9 1 10 11 7 1 10 11 9 1 9 1 9 1 9 7 9 7 10 9 0 0 1 13 10 9 7 10 9 2
24 9 2 10 9 7 10 9 1 10 9 1 13 1 9 7 10 9 1 10 9 1 10 9 2
17 10 9 13 1 10 9 13 10 9 7 10 9 2 1 3 16 2
21 2 3 1 10 9 1 10 9 13 13 3 13 1 10 9 9 1 10 9 0 2
10 10 9 4 13 0 9 1 15 3 2
17 2 15 13 3 9 1 9 1 10 9 1 10 9 1 10 9 2
2 9 12
2 12 2
86 9 2 10 9 7 10 9 13 1 10 9 2 1 9 7 1 10 0 9 0 2 3 1 10 9 1 10 9 2 10 9 1 9 0 13 10 9 0 1 10 9 1 10 11 9 7 1 10 11 9 1 9 1 9 1 9 7 9 1 9 1 15 13 10 9 1 13 15 2 7 10 9 0 1 10 9 0 0 1 13 10 9 7 10 9 2
36 9 2 10 9 7 10 9 4 13 1 10 9 2 1 9 7 1 10 0 9 0 2 1 9 3 1 10 9 1 10 9 2 10 9 0 2
11 0 2 9 2 9 1 9 0 7 9 2
26 9 13 1 10 9 2 1 9 2 9 7 9 1 10 9 2 9 1 9 7 9 9 1 10 9 2
40 16 0 9 7 9 3 13 2 10 9 4 1 10 9 13 1 10 9 0 1 9 7 1 10 0 9 15 15 13 1 13 1 9 1 10 9 7 10 9 2
34 0 2 1 10 9 7 10 9 1 9 1 10 9 2 9 15 13 1 13 10 9 0 1 10 9 7 10 9 0 1 10 10 9 2
42 0 2 9 1 10 9 0 1 10 9 1 9 15 13 10 9 1 9 1 9 1 10 9 7 1 10 9 1 9 15 13 10 9 1 9 1 9 1 9 7 9 2
2 12 2
14 10 11 9 13 16 15 13 1 10 9 10 9 0 2
23 9 2 1 9 1 10 9 15 13 1 9 2 10 9 13 3 10 9 9 1 10 9 2
34 9 2 10 10 9 0 4 13 1 9 7 1 10 0 9 0 7 0 1 10 9 7 4 4 15 13 3 1 10 9 1 10 9 2
6 10 9 15 13 9 2
28 9 2 10 9 1 10 9 9 2 3 4 13 10 9 0 7 2 1 10 0 9 2 1 9 7 1 9 2
2 12 2
51 10 9 15 13 1 10 9 1 13 1 10 9 15 13 2 4 13 10 10 9 2 16 4 13 10 9 7 10 9 1 10 9 0 3 1 10 9 2 1 10 9 15 13 10 10 9 13 1 10 9 2
50 10 9 15 13 10 10 9 15 13 7 10 9 13 3 0 1 10 9 1 10 9 7 1 10 9 9 1 10 9 1 10 9 1 10 9 1 10 9 2 7 1 10 0 9 0 0 1 0 9 2
2 12 2
49 9 2 10 9 13 1 10 9 3 4 4 13 2 1 3 16 10 9 3 15 13 3 10 9 2 1 9 7 1 9 2 7 13 10 0 9 1 9 2 3 1 13 9 1 10 9 1 10 2
12 2 9 1 9 2 13 10 9 1 10 9 2
26 2 9 7 9 1 10 9 2 10 9 1 9 2 1 9 7 1 9 1 10 9 7 1 10 9 2
13 2 9 1 9 13 1 10 9 15 13 1 9 2
24 9 2 10 9 13 1 10 9 3 4 13 1 10 12 9 15 13 10 9 13 1 10 9 2
2 12 2
46 16 3 1 10 9 10 9 4 13 1 13 1 9 0 10 9 0 1 10 9 1 10 9 2 4 13 15 1 10 3 3 1 10 9 1 13 15 1 13 10 0 9 2 1 9 2
10 2 13 1 10 9 1 9 1 9 2
23 2 7 13 10 9 0 1 10 9 10 15 13 10 9 13 7 10 10 9 1 10 9 2
16 10 9 4 13 3 3 10 9 7 10 9 1 10 10 9 2
2 12 2
41 1 10 9 1 10 9 0 0 0 2 15 13 10 9 0 1 10 9 1 10 9 16 4 13 1 10 9 12 2 9 12 2 9 9 2 2 13 10 9 0 2
28 0 2 10 9 15 10 9 4 13 1 10 9 1 10 0 9 15 4 13 7 15 13 1 10 9 1 9 2
69 0 2 10 9 1 9 1 9 2 3 3 10 9 1 10 9 1 10 9 13 1 13 10 9 13 1 9 1 9 1 10 9 2 1 10 9 1 10 9 7 1 10 0 9 1 1 10 9 1 15 10 9 3 13 1 10 0 9 1 9 1 9 7 0 9 13 3 0 2
34 3 10 9 3 15 13 1 10 9 1 9 1 0 9 7 1 0 9 2 3 1 10 9 16 4 13 1 9 7 1 10 0 9 2
39 0 2 10 9 13 1 9 1 10 9 1 9 7 1 9 13 1 9 13 1 10 9 1 9 2 3 16 0 9 4 10 9 1 10 9 1 10 9 2
10 0 2 10 9 1 10 9 7 9 2
64 13 3 13 15 15 13 13 1 13 10 9 1 10 9 1 9 1 9 2 9 2 9 7 9 1 10 9 2 1 10 9 0 7 0 1 10 9 0 1 10 9 2 13 10 9 7 10 0 9 7 15 4 13 3 1 10 9 1 10 9 1 10 9 2
42 2 12 2 13 16 10 11 9 4 4 13 10 9 1 9 0 1 9 1 10 9 15 13 13 10 9 0 2 16 13 1 10 9 0 1 13 9 1 10 9 13 2
25 16 10 11 9 4 4 13 16 10 9 0 13 3 1 10 9 0 0 13 1 10 11 9 0 2
2 12 2
55 1 10 9 1 10 9 1 15 1 10 9 12 2 12 7 12 2 10 11 9 3 13 1 10 9 10 9 0 1 9 1 10 9 15 13 7 13 7 10 9 0 1 13 3 9 7 9 15 13 10 9 1 9 0 2
2 12 2
73 10 11 9 4 13 16 10 9 1 9 1 10 9 1 10 9 4 13 1 13 1 9 10 0 9 0 1 13 9 7 9 0 1 10 9 1 10 10 9 7 1 13 1 10 9 0 2 1 10 9 2 9 15 13 10 9 1 10 9 1 10 10 9 1 15 13 9 1 9 1 10 9 2
44 2 12 2 10 9 1 10 11 9 1 13 10 9 1 10 9 1 9 0 13 3 10 9 13 1 9 0 7 3 10 9 0 13 1 10 9 1 13 9 0 1 0 9 2
36 2 12 2 10 11 9 13 1 10 9 1 13 10 9 1 10 9 1 9 0 1 9 1 10 9 0 1 9 1 9 13 1 10 9 0 2
63 2 12 2 13 16 10 11 9 2 1 10 9 1 13 10 9 1 10 9 1 9 2 13 2 1 15 13 10 9 3 0 2 10 9 1 13 10 9 1 9 7 1 9 1 9 15 13 0 1 10 9 1 13 10 9 1 10 9 1 9 1 9 2
65 2 12 2 13 10 9 1 13 1 10 9 10 0 9 1 9 7 10 9 1 10 11 1 13 15 1 9 0 15 13 9 7 13 10 9 13 1 10 11 9 1 10 9 1 10 9 0 2 0 7 0 1 10 9 1 9 1 10 9 1 10 9 15 13 2
72 2 12 2 13 16 10 9 1 13 10 9 1 9 7 10 9 1 9 1 9 13 1 9 0 1 10 9 1 10 9 1 10 9 2 1 3 13 1 10 9 3 0 1 10 9 9 0 1 13 7 1 13 10 9 1 10 9 7 3 13 15 1 13 1 9 0 1 9 1 9 0 2
2 12 2
2 12 2
14 10 9 13 4 3 13 10 0 9 0 1 10 9 2
35 1 9 1 9 2 1 10 9 1 10 0 9 13 10 9 1 9 1 15 10 11 9 4 13 10 9 0 1 10 9 13 1 3 0 2
23 2 12 2 10 0 9 3 13 10 9 0 1 10 9 0 13 10 9 13 1 10 9 2
44 3 10 0 9 3 4 13 10 9 1 13 10 9 1 10 9 1 15 13 1 9 1 9 0 1 9 1 9 0 13 1 10 9 1 10 11 9 1 15 13 10 9 0 2
20 10 0 9 13 0 1 10 10 10 9 7 3 0 1 15 1 10 11 9 2
2 12 2
37 16 10 9 1 9 4 4 13 1 10 9 3 1 10 0 9 2 10 9 4 13 1 10 9 1 10 9 13 1 10 9 2 15 4 13 3 2
32 10 0 9 3 1 9 1 10 9 13 1 10 9 1 10 10 9 1 9 13 10 9 0 1 9 1 10 9 1 10 9 2
17 10 9 4 13 1 10 0 9 0 7 1 10 9 1 12 9 2
2 12 2
38 10 11 9 13 1 10 10 9 9 0 16 10 9 4 13 1 13 1 10 9 15 13 9 1 10 9 0 7 1 10 9 0 10 9 1 10 9 2
73 12 2 16 13 10 9 1 15 1 10 9 12 2 0 9 2 10 9 4 13 1 13 16 1 10 9 3 10 9 15 2 3 1 10 9 0 2 4 13 1 10 9 1 10 9 7 10 9 7 15 13 1 9 1 13 3 3 1 10 13 1 10 9 1 15 1 10 9 12 2 0 9 2
11 10 0 9 4 4 3 13 1 10 9 2
2 12 2
50 10 9 4 13 1 13 1 10 9 2 3 3 7 1 10 3 3 1 12 9 1 9 2 10 10 9 1 15 13 15 1 9 1 10 9 1 9 2 1 9 1 10 9 1 15 1 10 9 12 2
2 12 2
86 1 10 9 1 9 13 9 15 13 1 13 10 9 1 9 7 10 9 7 10 9 1 10 9 2 10 15 4 13 1 10 9 0 0 0 7 3 4 4 13 1 10 9 1 10 10 9 2 10 9 0 0 0 4 13 1 10 9 16 10 9 7 10 0 9 15 13 13 3 1 10 9 0 7 15 13 3 1 10 9 1 10 9 1 9 2
2 12 2
47 10 9 1 15 1 10 9 12 13 9 15 13 1 13 1 10 9 0 10 9 7 10 9 0 0 1 13 13 10 9 0 1 10 9 1 10 0 9 1 15 7 3 1 10 0 9 2
2 12 2
48 0 9 13 2 16 1 10 9 2 10 9 2 1 9 1 9 0 2 1 10 9 1 10 10 9 1 10 9 7 9 2 1 9 10 9 2 1 9 1 9 2 1 10 9 1 10 9 2
46 13 16 3 13 13 10 9 1 10 11 9 1 13 7 13 10 9 2 0 7 0 2 1 13 9 3 1 10 9 0 16 15 4 13 2 1 10 9 2 1 10 9 1 10 9 2
22 10 0 9 13 10 0 9 0 1 10 9 0 0 15 13 10 9 0 1 10 9 2
19 15 13 3 9 13 10 9 0 0 2 15 3 3 4 13 1 9 0 2
46 0 9 0 4 2 1 9 2 13 9 1 9 0 7 9 0 15 13 1 13 9 1 10 9 7 13 15 2 3 1 10 9 1 10 9 0 7 10 9 1 10 9 1 10 15 2
2 12 2
7 10 9 0 0 4 13 2
2 12 2
26 10 9 7 10 9 0 1 10 9 1 10 0 9 4 13 1 9 13 1 10 9 7 4 3 13 2
46 2 12 2 10 9 3 0 1 10 9 1 9 1 10 9 7 1 10 9 4 4 13 10 9 1 9 0 13 1 10 9 7 4 3 13 1 10 9 0 7 1 10 9 0 13 2
39 10 11 1 10 9 0 2 1 10 9 12 7 12 2 13 10 9 13 1 10 9 7 13 16 4 13 10 9 1 10 9 7 10 9 1 10 10 9 2
2 9 0
2 9 0
2 9 12
3 9 1 9
2 12 2
23 10 0 9 15 13 1 10 9 0 1 9 2 9 7 9 2 13 1 9 1 9 0 2
20 15 15 13 3 1 10 9 1 9 13 1 9 0 1 10 9 1 9 0 2
2 12 2
88 1 10 9 1 10 0 9 10 9 9 0 13 10 9 1 15 2 1 9 1 9 1 10 9 2 10 9 1 9 7 10 9 1 9 2 16 15 13 7 3 9 1 9 7 9 2 4 13 7 1 10 9 1 12 11 9 7 1 10 9 1 10 0 11 9 16 4 13 10 9 1 10 9 1 10 0 11 2 3 16 10 11 3 13 10 11 9 2
36 1 10 9 1 10 0 9 3 15 13 9 0 10 9 1 12 9 1 10 9 1 10 0 11 9 1 9 13 1 10 9 1 10 0 11 2
2 12 2
81 1 10 9 1 10 0 9 10 9 13 1 3 9 0 15 13 13 10 0 9 16 10 9 15 4 13 1 10 0 9 2 3 1 10 9 16 4 4 13 1 9 1 10 0 9 7 1 9 1 3 9 7 10 10 9 0 3 13 3 1 10 0 9 16 10 9 7 3 9 4 4 13 3 1 10 9 1 10 0 11 2
2 12 2
23 10 0 9 15 13 3 1 10 9 1 15 1 10 9 0 2 13 0 10 9 3 13 2
2 9 12
10 9 13 1 10 11 7 9 1 9 0
2 12 2
31 10 0 9 15 13 1 10 9 13 1 10 11 7 1 10 9 0 1 9 0 16 13 10 9 1 15 1 10 9 12 2
2 12 2
35 1 10 9 1 9 0 10 9 13 0 3 1 10 9 1 10 9 0 0 3 1 10 9 0 1 10 9 1 10 9 7 10 9 0 2
2 12 2
24 1 15 13 1 10 9 12 2 10 9 1 10 0 9 3 15 13 1 10 9 1 9 0 2
2 9 0
16 9 7 9 1 10 9 1 9 1 9 1 9 2 9 7 9
2 9 12
3 9 7 9
2 12 2
19 1 9 1 10 9 1 9 4 4 13 10 9 1 9 0 7 0 13 2
13 9 2 10 9 1 10 9 1 9 7 1 9 2
44 9 2 16 10 9 1 9 7 1 9 4 13 1 10 9 1 10 0 11 9 7 16 13 13 15 7 3 9 1 10 9 1 10 0 9 2 10 9 1 15 1 0 9 2
2 12 2
28 1 9 1 10 9 1 9 1 15 1 10 9 12 4 13 10 9 1 10 9 9 15 13 10 9 3 0 2
29 16 4 13 15 10 1 10 0 9 10 9 4 13 15 1 13 1 10 9 10 9 0 13 10 9 1 15 13 2
2 12 2
14 10 9 13 1 10 9 10 9 0 1 10 9 13 2
2 12 2
47 1 10 9 4 4 13 10 9 13 1 10 15 4 13 16 10 9 1 10 9 1 9 7 9 2 1 9 2 9 7 9 1 10 9 7 1 9 13 0 1 10 0 9 2 16 0 2
2 12 2
2 9 12
1 9
2 12 2
13 1 10 9 1 9 4 13 10 9 1 9 0 2
2 12 2
27 1 9 1 10 9 1 9 0 4 13 10 9 1 10 0 9 15 13 10 9 0 1 10 9 1 13 2
41 16 4 13 15 1 0 9 10 9 13 1 10 9 2 1 9 1 10 9 2 10 9 1 9 15 13 10 9 1 10 9 7 10 9 1 10 9 1 15 13 2
2 9 12
13 13 1 10 9 1 9 0 7 1 10 9 1 9
13 10 9 1 9 0 7 10 9 1 9 4 13 2
13 9 2 10 9 1 10 9 1 9 7 1 9 2
43 9 2 16 10 9 1 9 7 1 9 4 13 1 10 9 1 10 0 11 9 7 4 13 15 7 3 9 1 10 9 1 10 0 11 2 10 9 1 15 1 0 9 2
11 9 2 10 9 1 10 9 1 10 9 2
2 9 12
8 9 0 1 10 9 1 10 9
36 16 0 1 10 9 1 10 9 0 2 1 9 7 9 1 9 0 0 2 10 9 4 4 13 1 13 10 9 15 13 10 9 1 10 9 2
18 10 9 3 4 13 1 9 1 10 9 10 9 2 9 7 0 9 2
2 9 12
7 9 1 10 9 1 9 0
2 12 2
15 10 9 1 9 0 4 13 1 10 9 1 12 9 0 2
2 12 2
18 10 0 9 13 10 9 2 1 10 9 2 7 4 13 1 10 9 2
22 10 0 9 13 10 9 2 1 10 9 2 7 4 13 1 10 9 7 1 10 9 2
2 12 2
19 10 9 1 10 9 7 15 1 10 9 4 4 13 7 13 1 10 9 2
2 12 2
35 16 2 1 9 1 10 9 2 10 9 13 10 9 1 9 0 2 15 13 2 3 1 9 0 2 16 15 4 13 1 9 1 10 9 2
2 9 12
2 12 2
39 10 9 9 13 10 9 0 2 0 7 0 0 1 13 15 1 10 0 9 1 10 9 1 12 9 1 10 10 9 2 12 2 7 15 13 3 10 11 2
2 12 2
24 10 9 1 15 1 10 9 12 2 9 12 2 15 13 1 13 1 10 9 1 10 0 9 2
16 10 9 13 0 1 10 9 13 1 10 9 1 10 10 9 2
2 9 12
2 9 12
30 10 9 9 13 1 13 1 10 11 10 9 1 10 9 0 1 9 0 15 15 13 1 10 9 13 1 10 0 9 2
2 9 12
28 10 11 13 10 12 9 1 10 11 10 9 1 10 9 1 10 0 9 7 15 13 2 16 0 2 9 0 2
2 9 12
10 10 9 9 13 9 1 10 0 9 2
30 1 10 9 1 10 0 9 2 1 2 9 2 15 13 10 9 0 2 3 16 13 9 1 10 0 9 0 7 0 2
10 1 2 9 2 15 13 3 10 9 2
2 9 12
2 12 2
54 10 9 2 9 2 13 10 9 1 10 9 0 2 10 9 1 10 9 0 7 10 9 1 10 9 0 2 7 10 9 15 2 13 10 10 9 2 9 7 10 9 0 1 10 9 2 15 13 1 9 1 10 15 2
2 12 2
73 1 9 1 10 9 1 10 9 2 15 13 10 9 1 10 11 0 1 10 9 1 10 9 2 1 10 9 2 1 10 2 9 2 7 1 10 0 9 1 9 1 10 9 1 10 10 9 0 2 4 13 9 1 10 15 1 10 9 1 10 0 9 7 13 0 1 10 0 9 1 10 9 2
2 12 2
46 16 3 4 4 13 10 9 1 10 9 15 13 15 10 9 1 9 16 10 9 13 1 10 9 2 1 10 9 0 2 10 9 1 10 9 7 1 10 9 15 15 4 13 10 9 2
36 10 0 9 15 13 1 10 9 13 2 16 15 3 13 10 9 1 10 9 1 15 1 10 9 12 2 3 16 4 13 10 9 1 10 9 2
2 9 12
18 10 9 4 13 10 9 2 10 9 7 10 9 0 1 9 7 9 2
2 9 12
35 16 2 1 9 1 10 0 9 2 3 9 13 9 1 10 0 9 2 15 13 1 9 2 13 0 10 9 0 1 9 1 9 1 9 2
2 9 12
2 12 2
25 10 9 13 0 16 3 13 10 9 15 15 15 4 3 13 13 9 1 10 10 9 2 1 15 2
8 9 2 10 9 1 10 9 2
14 9 2 10 9 1 10 15 10 9 4 13 3 13 2
13 9 2 10 9 1 10 9 1 9 1 10 9 2
2 12 2
25 10 9 3 4 4 13 0 1 10 0 9 16 10 9 3 13 4 4 13 1 9 3 1 15 2
2 9 12
15 10 9 3 13 0 1 10 9 1 10 0 9 16 13 2
11 9 2 16 3 4 13 10 9 1 9 2
34 9 2 16 2 13 9 1 10 9 2 13 9 13 16 10 9 15 4 13 10 9 3 13 16 15 4 13 1 9 7 4 13 3 2
36 9 2 16 3 4 13 10 9 1 10 9 7 10 0 9 1 9 1 9 0 2 7 15 4 13 7 13 1 10 9 1 10 10 9 0 2
22 9 2 16 10 9 4 13 1 10 9 1 10 9 1 9 0 13 1 10 9 0 2
32 9 2 16 10 9 1 10 9 0 7 9 1 10 9 1 15 4 13 1 9 10 9 3 13 1 13 10 9 1 10 9 2
43 9 2 1 10 9 1 10 9 1 10 9 0 2 16 10 9 4 13 1 10 9 1 10 9 1 15 4 4 13 10 9 7 1 10 9 13 1 10 9 1 10 9 2
2 9 12
2 12 2
40 13 0 10 9 0 1 9 1 9 1 9 2 10 9 1 10 9 3 13 13 16 10 9 4 13 3 1 10 9 1 10 9 7 1 10 9 1 10 9 2
2 12 2
47 10 9 1 10 9 4 4 13 7 0 2 13 9 1 10 10 9 2 16 10 9 4 13 3 1 10 9 1 10 9 7 1 9 1 10 9 7 1 10 9 1 15 10 9 13 0 2
2 9 12
15 1 10 9 1 10 9 12 2 1 2 9 2 15 13 2
29 9 2 10 9 7 10 9 1 10 9 0 1 10 9 0 2 0 9 1 10 9 1 12 11 2 16 10 9 2
15 0 2 13 1 10 9 3 13 1 10 9 7 9 0 7
16 0 2 4 4 13 1 10 9 3 1 10 9 7 9 0 2
14 10 0 9 13 0 10 9 0 0 1 10 9 0 2
16 13 10 9 15 13 10 11 0 0 2 1 9 10 9 12 2
10 13 10 9 1 10 11 2 12 2 2
11 13 10 9 1 10 11 0 2 12 2 2
86 13 16 10 9 1 10 9 0 1 9 1 9 1 10 9 1 10 9 13 1 10 9 0 1 10 10 9 13 0 16 10 9 0 1 0 9 4 13 10 9 1 10 9 7 13 10 0 9 1 10 9 1 10 9 1 10 9 0 13 9 1 10 9 1 9 1 10 9 1 10 9 13 1 10 10 9 7 1 10 10 9 1 10 9 0 2
28 13 16 1 10 9 1 10 9 10 9 15 13 2 10 9 1 9 13 3 0 7 10 9 0 7 0 13 2
25 16 3 13 3 0 13 16 10 9 13 0 2 1 9 1 9 2 1 10 9 1 10 10 9 2
22 16 10 10 9 4 3 13 15 1 10 9 1 9 0 2 13 3 0 10 9 0 2
35 13 16 1 10 9 1 10 0 9 1 10 9 4 4 13 10 9 1 13 1 9 0 1 10 9 1 10 9 1 10 9 1 10 9 2
42 13 16 1 10 9 0 1 10 9 9 10 9 4 13 9 1 10 9 1 9 1 10 9 0 7 1 10 9 0 1 10 9 0 13 1 15 9 1 10 0 9 2
32 16 2 1 10 9 1 15 0 9 13 3 15 10 9 1 10 0 9 1 10 9 2 15 3 4 4 0 1 10 0 9 2
47 16 2 1 10 9 1 15 10 9 0 1 10 9 1 10 9 1 10 9 0 4 3 13 1 10 9 9 3 1 10 9 0 1 9 2 4 3 13 1 13 0 9 13 1 10 9 2
43 13 16 2 1 10 9 1 15 10 9 1 9 0 13 3 13 1 10 10 9 9 1 0 9 0 2 13 0 13 1 10 9 1 9 1 10 0 9 9 1 10 9 2
52 13 16 10 9 1 10 9 0 7 1 10 9 1 10 9 1 10 9 1 9 1 10 0 9 4 4 13 1 10 9 9 2 13 9 1 10 9 1 10 9 1 10 9 2 1 10 0 9 1 10 9 2
16 16 13 3 13 0 1 10 9 9 13 10 9 1 10 9 2
66 13 16 1 0 9 10 9 1 10 9 1 13 15 1 10 9 16 13 16 10 9 1 10 9 0 7 9 1 10 9 1 15 4 13 10 9 1 9 3 13 1 13 10 9 1 10 9 2 4 4 13 1 10 9 9 1 10 9 0 1 10 9 1 10 9 2
27 16 4 3 13 0 1 10 11 9 13 1 10 10 9 7 13 1 10 0 9 10 9 1 10 9 0 2
39 16 1 9 1 0 9 10 9 1 10 9 4 3 4 13 1 10 9 1 8 8 0 1 13 2 16 0 2 1 9 0 10 9 1 9 1 10 11 2
38 13 16 2 13 9 1 10 9 0 1 10 0 9 1 10 9 9 2 3 4 13 13 10 9 0 1 10 9 1 10 9 2 0 1 10 10 9 2
84 16 3 2 1 10 9 1 15 13 9 0 2 13 0 13 16 10 9 9 4 13 1 10 9 1 10 9 0 13 10 9 1 10 9 0 1 10 9 1 10 9 7 10 9 0 13 1 9 0 15 13 10 0 9 2 1 9 16 10 9 4 13 1 10 9 3 13 1 13 10 13 9 1 10 9 7 10 13 9 1 10 9 0 2
24 13 16 10 9 0 1 10 0 9 3 4 1 9 13 0 7 13 10 9 1 10 0 9 2
31 16 13 0 3 16 1 10 11 13 13 1 9 0 9 1 10 11 1 10 9 1 10 0 9 2 13 3 1 9 0 2
64 13 16 1 10 9 13 3 0 13 1 10 9 1 10 9 1 10 0 9 13 10 9 13 1 10 9 9 2 1 10 9 1 10 9 3 0 1 4 13 1 10 9 0 1 10 9 1 0 9 1 10 9 1 10 9 7 1 10 9 1 10 9 0 2
47 13 16 3 10 9 1 10 9 2 0 1 10 10 9 2 13 10 13 9 1 10 9 2 0 1 10 9 13 1 10 9 0 2 1 10 0 9 1 10 9 0 1 10 9 0 0 2
19 13 16 10 9 15 13 3 1 10 9 0 15 13 9 1 10 9 0 2
35 16 3 13 13 1 13 9 10 9 0 7 10 9 1 10 9 2 3 16 4 4 13 1 10 9 1 9 0 15 4 13 15 10 9 2
28 16 10 9 13 1 10 0 9 13 3 1 10 9 0 9 1 10 9 1 9 1 9 7 13 1 9 0 2
40 13 16 1 10 9 1 10 9 1 10 9 13 0 13 0 10 10 9 1 10 9 0 16 10 9 0 7 10 9 0 7 10 9 0 1 15 13 13 0 2
52 16 1 10 0 9 13 0 16 4 13 10 9 1 10 9 15 13 9 1 10 11 0 7 15 1 15 15 13 1 9 13 10 10 9 2 9 7 10 9 0 7 13 10 9 10 10 9 3 4 4 13 2
37 13 16 2 16 1 10 0 9 13 0 3 9 2 10 9 1 10 9 13 16 10 9 4 13 10 9 0 1 10 9 1 15 10 1 10 9 2
65 13 16 1 13 10 9 1 10 10 9 0 7 1 10 10 9 13 0 16 10 9 0 1 10 9 4 13 3 3 1 9 1 10 9 1 10 9 1 10 9 1 9 1 10 10 9 2 7 1 9 1 10 9 1 10 9 15 10 0 9 4 3 13 15 2
19 16 10 9 4 13 13 10 9 0 1 10 9 15 1 10 9 4 0 2
35 13 16 10 0 9 1 10 9 1 10 9 7 10 9 13 16 10 9 4 13 15 1 10 9 16 13 10 9 1 10 9 15 15 13 2
30 13 16 10 9 1 10 9 13 16 10 9 1 10 9 3 13 1 10 9 1 10 9 15 4 13 1 13 10 9 2
20 16 3 10 9 0 1 10 9 4 4 13 1 9 1 13 7 13 10 9 2
12 1 10 9 4 13 10 9 11 1 11 11 2
9 15 13 10 9 0 1 10 11 2
11 1 10 9 15 13 10 9 1 11 11 2
9 15 13 10 9 1 9 1 9 2
9 1 15 13 10 9 0 10 9 2
10 15 13 10 9 9 1 10 9 11 2
15 10 9 1 10 9 4 13 1 10 9 1 10 9 11 2
5 15 13 11 11 2
6 10 9 13 11 11 2
9 15 13 10 9 0 1 10 11 2
16 1 15 13 10 9 1 10 9 0 15 15 4 13 1 11 2
7 1 10 9 13 10 11 2
8 3 4 13 10 9 0 0 2
16 10 9 13 10 0 9 1 9 1 10 9 1 10 11 11 2
12 1 10 9 4 4 13 10 9 0 1 11 2
6 1 10 9 13 11 2
7 10 9 15 13 1 11 2
13 10 9 1 9 4 4 13 1 10 11 11 11 2
10 3 15 13 10 9 1 9 1 11 2
13 15 13 10 3 0 9 1 9 0 1 10 9 2
10 1 10 9 4 13 10 11 11 11 2
9 15 13 10 9 1 9 1 11 2
7 10 9 15 13 1 11 2
10 15 13 10 9 1 2 11 11 2 2
8 15 13 10 9 1 10 11 2
9 10 9 0 13 10 2 11 2 2
20 15 13 10 9 1 10 9 1 11 11 1 11 11 2 11 11 7 11 11 2
9 10 9 13 1 9 1 10 11 2
10 15 13 10 0 9 1 10 11 11 2
8 15 13 10 9 1 11 11 2
13 15 13 11 11 1 10 0 9 1 10 9 12 2
13 15 13 11 11 1 10 0 9 1 10 9 12 2
7 1 15 15 13 10 9 2
13 10 9 13 11 2 10 9 0 1 10 9 11 2
11 1 10 9 0 13 9 11 11 1 9 2
6 3 4 13 11 11 2
9 15 13 10 9 1 11 11 11 2
7 1 15 4 13 11 11 2
19 1 10 9 11 11 4 13 1 13 1 10 9 1 10 2 11 11 2 2
9 1 10 9 0 15 13 11 11 2
10 3 15 13 10 9 0 1 11 11 2
8 15 13 10 9 1 10 9 2
6 10 15 13 10 11 2
6 10 15 13 10 11 2
17 1 10 9 4 4 13 11 11 1 10 9 1 10 11 1 11 2
11 10 9 4 4 13 1 10 11 1 11 2
8 15 13 10 9 0 3 13 2
10 10 9 13 1 9 1 10 11 11 2
10 15 13 10 9 9 1 10 9 0 2
8 1 10 9 4 4 13 11 2
7 3 4 13 10 9 0 2
21 1 10 9 13 10 9 15 4 13 10 9 0 3 1 11 7 11 1 10 12 2
7 3 4 13 10 9 0 2
7 15 13 10 0 1 11 2
9 3 15 13 10 9 1 11 11 2
8 15 13 10 9 1 10 11 2
12 10 9 0 13 1 9 1 13 10 9 0 2
9 1 10 15 4 13 10 9 0 2
11 1 10 15 4 13 10 9 1 10 9 2
9 15 4 13 10 9 1 10 9 2
22 1 10 1 3 1 10 9 0 4 4 13 10 9 0 1 2 9 1 10 9 2 2
6 10 9 13 10 9 2
9 15 13 10 9 0 1 10 9 2
8 15 13 10 9 1 10 9 2
8 15 13 10 9 1 10 9 2
11 1 10 9 15 13 10 9 1 11 11 2
10 10 9 1 11 13 10 9 1 9 2
14 10 9 0 15 4 13 1 10 11 11 1 10 12 2
11 1 10 9 4 4 13 10 9 1 11 2
9 1 15 13 10 9 1 10 11 2
9 10 9 1 9 4 13 11 11 2
8 3 15 13 10 9 0 0 2
13 10 9 15 13 1 10 9 1 10 9 1 11 2
6 10 15 13 10 11 2
12 1 10 9 13 10 9 1 10 9 1 11 2
13 3 4 4 13 10 9 1 10 9 1 10 9 2
10 13 10 9 1 10 9 13 1 9 2
16 1 10 9 10 9 4 13 1 13 15 1 10 9 1 9 2
8 10 9 15 13 1 10 9 2
9 15 13 10 9 1 10 9 0 2
5 3 13 10 9 2
10 10 9 0 4 13 0 1 10 9 2
6 15 4 13 10 9 2
5 3 4 13 11 2
7 1 10 9 13 0 11 2
12 15 13 10 9 1 10 0 9 13 1 11 2
9 10 9 13 1 9 1 10 9 2
9 15 13 10 9 0 1 10 9 2
11 15 13 10 9 1 9 1 10 9 0 2
14 15 13 10 9 0 3 1 9 1 9 1 10 9 2
15 13 10 9 1 10 9 1 10 9 13 1 10 9 11 2
11 3 15 13 1 10 0 9 10 9 11 2
13 13 10 9 1 15 15 13 10 9 1 9 11 2
11 10 15 13 10 11 11 1 10 11 11 2
7 3 15 13 10 9 11 2
7 13 10 9 1 10 9 2
11 1 10 9 13 10 9 1 10 9 0 2
6 3 15 9 11 11 2
5 3 15 13 11 2
10 1 15 4 13 10 9 1 10 11 2
8 1 15 13 10 9 10 9 2
6 15 13 10 9 0 2
5 15 13 10 9 2
6 15 13 10 9 0 2
7 10 9 13 9 1 11 2
6 3 13 0 10 11 2
9 3 15 13 10 9 1 11 11 2
13 13 10 9 1 10 9 15 13 0 1 13 9 2
8 15 4 13 10 2 11 2 2
8 3 13 10 11 1 10 11 2
9 3 15 13 10 9 1 9 0 2
9 3 15 13 10 0 11 7 11 2
9 15 4 13 10 9 1 10 11 2
10 1 10 9 15 4 13 10 9 11 2
6 10 15 13 10 11 2
9 13 10 9 1 9 1 10 9 2
8 1 10 9 0 4 13 11 2
11 1 10 9 10 9 15 4 13 1 11 2
9 1 10 15 4 13 10 9 0 2
7 15 4 13 2 11 2 2
6 15 13 11 11 11 2
13 3 15 4 13 10 9 1 10 11 1 10 11 2
5 13 10 9 0 2
11 3 13 10 9 0 1 10 11 11 11 2
5 15 13 10 9 2
6 3 4 13 11 11 2
10 1 10 9 10 9 1 11 13 0 2
8 1 3 4 13 10 9 0 2
6 3 13 10 11 11 2
11 3 15 13 10 9 1 9 1 10 9 2
5 15 13 11 11 2
5 15 13 10 9 2
8 3 15 13 10 9 1 11 2
11 15 13 10 9 1 2 11 1 9 2 2
6 10 15 13 10 9 2
7 3 4 4 13 10 9 2
9 1 10 9 13 10 9 1 9 2
8 15 13 10 9 1 11 11 2
6 10 15 13 10 11 2
9 10 9 3 13 10 9 1 9 2
6 3 13 10 9 11 2
10 10 9 13 10 9 1 13 10 9 2
9 15 13 10 9 1 9 1 11 2
7 1 10 9 13 11 11 2
7 1 10 9 13 10 11 2
11 1 10 9 4 13 10 11 1 10 9 2
5 15 4 13 11 2
8 15 13 10 9 1 10 11 2
9 10 9 1 9 15 13 1 11 2
5 15 13 10 9 2
9 3 15 13 10 9 1 11 11 2
9 13 10 9 1 10 9 1 9 2
12 1 10 9 15 4 13 10 11 1 10 11 2
11 10 9 4 13 10 9 1 10 9 0 2
10 15 13 10 3 0 9 0 1 11 2
5 10 9 13 11 2
5 10 9 13 0 2
6 10 15 13 11 11 2
5 15 13 11 11 2
8 10 15 13 2 11 11 2 2
6 10 15 13 10 9 2
9 13 10 9 1 10 9 1 9 2
8 3 4 4 13 10 9 11 2
5 15 13 10 11 2
6 10 15 13 10 9 2
10 1 10 15 4 4 13 11 11 11 2
7 3 15 13 10 11 11 2
16 10 9 4 13 1 10 9 0 1 10 9 2 11 11 2 2
15 13 10 9 1 10 9 0 15 4 4 13 1 11 11 2
10 1 10 9 9 11 11 11 13 9 2
10 15 13 10 9 1 11 1 10 11 2
5 15 13 11 11 2
6 10 9 13 11 11 2
9 1 10 9 4 13 10 11 11 2
7 13 10 9 1 10 9 2
6 3 15 4 13 9 2
11 10 9 15 13 1 10 9 0 1 11 2
5 3 13 10 9 2
9 1 10 15 4 13 10 9 0 2
8 1 10 9 13 10 11 11 2
10 13 10 9 1 15 15 13 10 9 2
7 13 10 9 15 13 9 2
9 10 9 13 10 0 9 1 9 2
7 10 9 4 13 11 11 2
13 10 9 4 13 1 10 11 1 12 9 1 9 2
13 10 9 4 13 11 11 2 11 11 7 11 11 2
17 10 9 1 10 9 0 1 10 9 4 13 1 11 1 10 12 2
14 10 9 13 1 11 7 11 1 10 9 1 10 12 2
8 10 9 13 10 9 1 11 2
7 3 9 13 10 9 11 2
7 15 13 0 10 11 11 2
12 15 4 13 11 1 13 10 11 0 1 11 2
15 10 9 4 13 0 1 10 11 1 10 9 2 11 2 2
11 10 9 15 13 1 9 1 10 9 11 2
11 10 9 13 1 9 1 10 0 1 11 2
13 10 9 1 10 9 1 11 7 11 13 1 9 2
9 3 15 13 10 9 1 10 9 2
13 10 9 4 13 10 9 1 10 2 11 11 2 2
10 13 10 9 1 10 9 0 7 0 2
5 3 13 10 11 2
13 10 9 13 3 1 12 9 7 9 1 10 11 2
12 10 9 13 1 11 11 11 15 13 10 9 2
16 10 9 0 4 4 13 1 11 11 1 10 9 1 10 12 2
14 10 9 0 13 1 9 10 9 0 1 10 0 9 2
7 1 10 9 15 13 11 2
6 3 4 13 10 11 2
10 3 15 13 10 11 11 1 10 12 2
11 1 10 9 15 13 10 9 1 10 9 2
9 1 10 9 13 10 9 1 9 2
9 3 15 13 10 9 1 10 11 2
7 3 15 13 11 1 11 2
11 3 4 13 9 10 11 0 1 10 9 2
5 3 15 13 11 2
8 10 9 0 4 13 10 11 2
11 15 13 10 9 0 1 10 11 11 11 2
16 15 4 13 10 9 0 2 10 9 0 1 10 10 9 2 2
11 15 13 1 9 1 10 0 9 1 11 2
10 15 4 13 2 10 9 1 11 2 2
31 15 4 13 10 9 11 1 10 11 1 10 9 0 7 0 1 10 10 9 1 10 9 1 10 0 9 0 1 10 9 2
15 15 4 13 1 13 10 9 1 9 2 11 11 11 2 2
17 15 4 13 10 0 11 1 10 11 11 7 11 11 1 10 11 2
12 15 4 13 10 9 1 10 11 11 1 11 2
15 15 4 13 10 0 11 11 1 9 2 11 1 11 2 2
10 3 13 1 9 10 0 9 1 11 2
11 1 10 9 10 11 4 13 1 10 11 2
9 1 10 9 4 4 13 11 11 2
10 10 9 13 10 9 1 10 0 9 2
12 1 10 9 1 10 9 12 13 10 9 9 2
7 3 10 9 13 10 11 2
7 3 13 1 9 10 11 2
9 3 11 11 11 15 13 1 11 2
5 13 10 9 0 2
10 13 10 9 1 10 9 1 9 9 2
9 1 10 9 11 11 13 1 9 2
14 1 10 9 0 10 11 4 13 10 9 1 9 0 2
6 10 9 4 13 11 2
8 10 9 4 13 11 11 11 2
11 10 9 13 10 0 9 0 1 10 11 2
16 10 9 0 4 3 13 1 10 0 9 10 9 7 10 9 2
13 10 9 4 13 0 9 1 10 9 1 10 9 2
24 10 9 4 13 11 2 11 2 11 2 11 2 11 11 7 11 2 11 7 11 11 1 11 2
6 10 15 13 10 11 2
8 10 15 13 10 2 11 2 2
5 15 13 11 11 2
5 15 13 11 11 2
5 15 13 11 11 2
5 15 13 11 11 2
6 10 15 13 10 11 2
6 15 13 11 11 11 2
7 10 15 13 10 11 11 2
18 1 10 9 10 9 1 10 11 11 4 13 1 1 10 12 9 12 2
15 15 13 10 9 1 10 11 1 10 11 3 1 10 12 2
14 15 13 10 9 1 10 11 1 10 11 1 10 12 2
10 10 9 0 15 4 13 1 10 12 2
19 1 10 9 2 3 1 10 12 2 15 4 13 10 11 0 1 10 9 2
12 15 13 10 9 11 1 10 9 1 10 12 2
14 10 9 4 13 10 9 0 1 10 9 12 2 12 2
16 10 9 0 4 13 12 9 2 11 11 11 2 1 10 12 2
22 15 13 10 9 0 1 10 11 1 10 9 12 2 12 1 10 9 1 10 9 0 2
10 15 13 10 9 0 1 13 10 9 2
12 3 15 4 13 10 9 1 9 1 10 9 2
10 3 4 4 13 10 9 1 10 9 2
12 3 15 13 1 13 3 10 9 0 1 11 2
11 1 10 9 11 2 3 13 9 10 9 2
7 3 4 13 10 9 0 2
9 3 4 13 10 2 11 11 2 2
11 3 4 4 13 10 9 1 10 9 0 2
7 3 15 13 10 9 11 2
8 3 13 10 9 1 10 9 2
5 15 13 11 11 2
5 15 13 11 11 2
5 3 15 13 11 2
5 15 13 11 11 2
6 10 15 13 10 11 2
5 3 15 13 11 2
14 15 13 10 9 1 10 11 1 9 1 10 9 0 2
8 15 13 10 9 1 10 11 2
6 10 15 13 10 11 2
7 15 13 10 0 9 0 2
7 11 1 10 9 15 13 2
10 15 13 10 9 1 10 9 0 0 2
8 11 11 1 10 9 13 9 2
8 13 10 9 1 10 9 0 2
5 3 15 13 11 2
6 10 9 13 1 11 2
8 15 13 10 9 1 10 11 2
6 10 15 13 10 11 2
9 3 13 10 9 0 1 10 11 2
6 10 9 13 10 11 2
5 15 4 13 11 2
10 1 10 9 15 13 10 9 11 11 2
14 15 13 10 9 1 10 9 1 10 9 0 11 11 2
8 13 10 9 1 10 9 0 2
6 10 15 13 10 11 2
6 10 15 13 10 11 2
7 1 10 9 15 13 11 2
10 1 10 9 0 15 13 10 11 11 2
5 15 13 11 11 2
5 15 13 11 11 2
9 15 4 13 10 9 1 10 11 2
7 10 15 13 11 11 11 2
9 15 13 10 9 1 10 9 0 2
8 15 13 10 9 1 10 11 2
10 15 13 10 9 0 1 10 9 0 2
8 1 10 9 15 13 11 11 2
5 10 15 13 11 2
11 3 15 4 13 10 9 1 9 1 11 2
6 3 4 13 11 11 2
12 15 13 10 9 1 10 9 1 10 9 0 2
19 15 13 10 9 1 10 9 1 10 9 7 9 1 10 9 11 11 11 2
11 15 13 10 9 1 10 11 1 10 11 2
8 15 13 10 9 1 10 11 2
5 15 13 11 11 2
6 10 9 13 10 11 2
6 10 15 13 10 11 2
10 15 4 13 10 11 11 11 1 11 2
7 15 13 10 9 1 11 2
12 3 15 13 10 9 1 10 9 0 11 11 2
8 1 10 9 15 13 11 11 2
7 15 13 10 0 9 0 2
7 15 13 10 9 1 11 2
10 1 10 9 1 9 13 11 11 11 2
12 10 9 1 10 11 4 13 9 1 10 11 2
12 15 13 10 9 1 10 9 1 10 11 11 2
8 13 10 9 1 10 9 0 2
10 1 10 9 4 13 10 9 0 11 2
5 15 13 11 11 2
8 1 10 9 4 13 11 11 2
6 15 13 11 11 11 2
8 3 11 13 10 9 1 11 2
6 3 15 13 10 11 2
9 15 13 10 9 1 10 9 11 2
7 10 15 13 10 11 11 2
10 1 10 9 15 13 10 9 1 11 2
10 3 15 13 10 9 1 10 11 11 2
9 1 10 9 4 4 13 10 11 2
6 3 4 13 11 11 2
7 15 13 10 0 9 0 2
7 10 9 15 13 1 11 2
7 10 15 13 10 9 11 2
6 15 4 13 11 11 2
13 15 13 10 9 1 9 1 10 9 1 9 11 2
8 1 10 9 13 9 11 11 2
10 10 9 13 10 0 9 0 11 11 2
10 15 13 10 9 1 10 11 11 11 2
12 3 15 4 13 11 11 1 10 9 1 11 2
5 15 13 11 11 2
14 15 13 10 9 2 11 2 16 15 13 1 9 11 2
7 1 10 9 13 11 11 2
13 15 4 13 10 0 9 1 10 9 0 1 11 2
10 10 9 13 1 10 9 1 11 11 2
10 13 10 9 15 13 1 10 9 9 2
9 3 15 13 10 9 1 9 0 2
5 10 15 13 11 2
10 10 9 13 10 0 9 1 11 11 2
12 15 13 10 3 0 9 1 9 1 10 9 2
6 10 15 13 10 11 2
5 15 13 11 11 2
5 15 13 10 11 2
6 10 15 13 10 11 2
6 3 4 13 11 11 2
7 15 13 10 11 1 11 2
6 3 4 13 11 11 2
6 3 4 13 11 11 2
5 3 15 13 11 2
5 15 13 10 11 2
14 15 13 10 9 1 10 11 1 10 9 1 10 11 2
8 10 9 0 13 1 10 11 2
5 10 9 13 11 2
10 1 10 15 11 13 10 9 1 11 2
6 3 11 13 10 9 2
11 15 13 10 9 1 10 9 0 1 11 2
8 3 10 9 11 11 13 11 2
11 3 13 10 9 0 1 10 11 11 11 2
5 15 13 10 11 2
9 10 9 13 10 9 0 1 11 2
7 3 4 4 13 11 11 2
5 15 13 10 11 2
6 10 15 13 10 11 2
8 15 13 10 9 1 10 11 2
13 15 13 10 9 0 1 10 9 0 1 11 11 2
15 15 15 4 4 13 1 0 9 1 10 11 1 10 12 2
8 3 4 4 13 10 11 11 2
7 15 4 13 10 11 11 2
8 10 9 13 1 10 11 11 2
5 15 13 11 11 2
13 15 4 13 10 9 11 1 10 9 1 10 12 2
5 15 13 11 11 2
8 15 13 10 9 1 10 11 2
11 15 13 10 3 0 9 0 1 10 11 2
18 1 15 13 10 9 1 10 9 0 1 9 7 9 11 1 10 12 2
11 3 10 11 4 13 1 9 10 0 11 2
11 3 4 4 13 10 11 11 2 11 2 2
14 10 9 4 13 1 10 11 1 10 9 1 10 12 2
6 3 13 10 9 11 2
5 3 13 10 11 2
7 10 9 9 13 10 11 2
20 15 4 13 1 13 12 9 13 10 9 1 10 11 2 9 9 1 11 11 2
5 15 13 11 11 2
11 3 13 10 9 0 1 10 11 5 11 2
6 3 4 13 10 11 2
7 10 9 13 1 10 11 2
8 15 13 10 9 1 10 11 2
6 10 9 13 10 11 2
5 15 13 11 11 2
13 3 10 9 0 1 10 9 0 4 13 1 11 2
9 10 9 4 13 10 11 11 11 2
9 3 9 4 13 10 11 11 11 2
7 3 4 13 10 11 11 2
8 15 13 10 9 1 10 11 2
5 15 13 11 11 2
13 1 10 9 10 11 4 13 10 9 1 10 12 2
5 15 13 11 11 2
11 15 4 13 1 10 9 1 9 0 11 2
6 10 15 13 10 11 2
9 3 11 13 11 0 1 10 9 2
5 15 13 11 11 2
13 3 13 10 9 1 10 11 11 11 2 11 2 2
6 10 15 13 10 11 2
12 3 15 13 10 9 0 1 10 9 0 0 2
6 10 15 13 10 11 2
6 10 15 13 10 11 2
7 15 13 10 2 11 2 2
9 3 4 13 1 10 9 10 11 2
14 10 0 9 4 4 13 1 10 11 7 1 10 11 2
11 10 15 13 10 11 11 11 2 11 2 2
7 10 9 13 10 9 11 2
5 15 13 10 11 2
10 3 10 11 4 13 1 10 10 9 2
11 3 15 13 10 3 0 9 1 10 9 2
10 15 13 10 9 3 0 1 10 11 2
7 15 13 10 9 1 11 2
12 1 10 15 4 13 3 10 11 1 10 12 2
11 10 9 13 13 1 10 11 1 10 12 2
10 15 13 2 11 11 2 1 10 11 2
10 1 15 4 13 12 9 1 10 11 2
8 10 9 15 4 13 1 11 2
9 3 4 13 10 9 1 9 11 2
9 15 15 13 1 11 1 10 11 2
11 15 4 4 13 9 1 10 11 11 11 2
8 10 15 13 10 9 0 11 2
6 10 15 13 10 11 2
9 3 4 13 10 9 11 1 11 2
8 10 15 13 11 11 1 11 2
11 10 9 13 10 9 1 11 1 10 11 2
10 10 15 4 13 1 10 11 11 11 2
5 15 13 11 11 2
6 10 15 13 10 11 2
10 3 15 13 10 9 1 10 9 0 2
5 3 15 13 11 2
14 3 4 13 10 9 1 10 9 0 1 11 1 11 2
5 15 13 11 11 2
6 3 15 13 10 11 2
12 10 9 4 13 1 10 9 1 9 1 11 2
10 10 15 13 10 11 1 10 11 11 2
8 3 15 13 10 9 0 0 2
13 3 15 13 10 9 15 13 1 11 1 10 12 2
11 15 4 13 10 9 1 10 0 1 11 2
11 3 4 13 9 10 11 0 1 10 9 2
6 3 13 9 10 11 2
8 3 10 11 4 13 1 11 2
7 15 13 10 9 1 11 2
5 15 13 11 11 2
5 15 13 10 11 2
9 3 15 13 10 9 1 11 11 2
9 15 13 10 9 1 2 11 2 2
10 3 15 13 10 9 1 10 11 11 2
5 15 13 11 11 2
11 15 4 13 10 11 1 11 1 10 12 2
5 15 13 11 11 2
8 15 13 10 9 1 10 11 2
5 15 13 11 11 2
6 10 15 13 10 11 2
7 3 15 13 10 9 11 2
6 10 15 13 10 11 2
8 15 13 10 9 1 10 11 2
17 3 15 4 13 10 0 9 1 10 9 0 1 11 1 10 12 2
9 10 9 13 11 11 1 10 12 2
12 3 4 4 13 10 9 1 9 1 11 11 2
10 3 15 4 13 10 0 9 1 11 2
13 15 4 4 13 9 1 10 11 11 1 10 11 2
13 3 15 13 10 0 9 0 13 1 10 9 12 2
9 3 4 4 13 10 9 1 11 2
8 15 13 10 9 1 11 11 2
7 15 13 10 0 9 0 2
12 3 15 4 13 10 11 0 1 9 7 9 2
10 3 15 4 13 10 0 11 1 11 2
8 15 13 10 9 1 10 11 2
9 10 9 13 10 11 1 11 11 2
10 3 15 13 10 9 1 10 9 0 2
5 3 15 13 11 2
10 15 13 10 9 1 10 11 11 11 2
12 15 13 10 9 1 10 11 11 1 10 12 2
6 3 4 13 11 11 2
9 10 15 13 10 9 2 11 2 2
9 15 4 13 10 9 0 1 11 2
7 10 9 4 13 11 11 2
17 15 4 4 13 1 11 11 1 10 9 1 10 11 1 11 11 2
9 1 10 9 13 10 9 11 11 2
8 15 4 13 10 11 1 11 2
10 15 13 10 9 1 9 1 11 11 2
7 3 4 13 11 11 11 2
11 3 15 13 10 0 9 0 1 10 11 2
8 15 13 10 9 1 10 11 2
7 10 9 13 1 9 11 2
12 15 13 10 9 1 9 1 11 1 10 12 2
8 15 13 10 9 1 10 11 2
8 15 13 10 9 1 10 11 2
15 3 15 4 13 10 0 9 1 10 9 1 10 11 11 2
9 1 10 9 11 11 13 9 0 2
14 10 9 4 13 10 11 1 10 11 11 1 10 12 2
18 10 9 13 1 9 1 11 11 1 10 9 1 10 9 1 10 11 2
6 3 15 13 10 11 2
9 3 15 4 13 10 11 11 11 2
6 10 9 13 10 11 2
14 15 13 10 9 1 11 11 2 0 9 1 10 11 2
21 10 9 4 13 10 0 9 0 1 10 9 1 10 11 0 1 10 9 1 11 2
11 15 13 10 9 1 2 11 1 11 2 2
18 15 4 13 10 9 1 0 9 1 10 11 0 1 10 9 1 11 2
10 3 15 13 10 0 9 1 10 11 2
12 15 13 10 9 1 9 1 10 9 11 11 2
8 15 13 10 0 9 1 11 2
7 3 4 4 13 11 11 2
8 10 9 13 11 11 1 11 2
12 10 9 11 11 13 13 1 13 1 10 12 2
16 3 4 13 10 11 1 10 11 11 16 4 4 13 1 11 2
8 10 9 13 1 10 9 11 2
10 3 15 4 13 11 11 7 11 11 2
16 15 13 10 9 1 9 1 10 11 1 10 9 1 10 12 2
11 15 13 10 9 0 3 0 1 10 9 2
11 3 15 4 13 10 9 0 1 10 9 2
12 15 13 10 9 0 1 10 11 1 10 11 2
8 1 10 9 4 13 11 11 2
6 3 4 13 11 11 2
11 1 3 13 1 9 10 9 1 10 11 2
9 15 13 10 9 1 11 11 11 2
7 3 13 10 11 1 11 2
8 3 15 13 10 9 11 11 2
5 3 13 11 11 2
6 3 4 13 11 11 2
9 15 13 10 3 0 9 1 11 2
9 15 13 10 0 9 1 10 11 2
8 1 10 9 13 11 1 11 2
5 3 13 11 11 2
6 3 4 13 11 11 2
9 3 15 13 10 9 11 1 11 2
11 15 13 10 3 0 9 1 10 11 11 2
10 15 13 10 9 3 0 1 10 11 2
8 15 13 10 9 1 10 11 2
8 1 10 15 13 10 9 11 2
9 1 10 9 10 11 13 10 11 2
9 1 10 9 0 15 13 11 11 2
9 3 15 13 10 11 1 10 11 2
6 15 4 13 10 9 2
9 15 4 13 2 10 0 9 2 2
11 15 13 10 9 0 1 9 1 10 9 2
8 15 13 2 10 9 0 2 2
11 15 13 10 9 0 1 10 11 11 11 2
7 1 15 13 9 11 11 2
7 15 13 10 9 1 11 2
7 15 13 10 9 1 11 2
8 15 13 10 9 0 1 11 2
6 15 4 13 11 11 2
10 15 4 13 10 0 9 1 11 11 2
8 15 13 10 9 1 10 11 2
10 15 13 10 9 1 10 9 1 11 2
10 15 4 13 10 9 2 11 11 2 2
9 3 15 13 10 9 1 10 11 2
8 15 13 10 0 9 1 11 2
7 10 9 4 13 11 11 2
9 1 10 9 11 11 13 10 0 2
12 10 9 4 13 10 11 11 1 9 1 9 2
8 1 10 9 13 9 11 11 2
10 10 9 13 10 9 1 11 1 11 2
8 1 10 9 13 9 11 11 2
12 15 13 10 11 2 9 0 1 9 0 2 2
7 10 9 13 10 11 0 2
7 10 9 15 13 1 11 2
7 15 13 0 10 9 11 2
7 10 9 13 11 1 11 2
6 15 13 11 1 11 2
6 15 13 0 10 11 2
9 15 13 10 9 1 10 11 11 2
7 10 9 13 10 11 11 2
10 10 9 4 13 11 1 10 10 9 2
7 1 10 9 13 10 9 2
12 3 4 13 10 11 11 1 11 1 10 11 2
7 3 4 13 0 11 11 2
10 3 4 13 10 9 2 11 11 2 2
11 3 4 13 10 9 0 1 10 9 0 2
6 3 4 13 11 11 2
11 1 10 9 15 13 10 9 1 10 11 2
10 3 2 10 11 2 4 13 9 0 2
9 1 10 9 4 13 10 12 9 2
6 9 4 13 10 11 2
13 15 13 10 9 1 10 9 1 10 11 1 11 2
8 15 4 13 10 12 9 12 2
8 1 10 15 13 0 11 11 2
11 10 9 13 10 9 1 10 9 1 9 2
5 3 4 13 11 2
16 10 11 3 4 13 9 1 10 9 1 9 1 10 0 9 2
8 15 13 10 0 9 0 0 2
8 10 15 13 11 1 10 9 2
8 10 0 13 9 1 10 11 2
8 15 13 10 9 1 11 11 2
7 1 10 9 13 11 11 2
7 1 10 9 13 11 11 2
12 1 10 9 1 9 13 11 0 1 11 11 2
11 1 10 9 4 13 10 9 1 10 11 2
7 10 9 0 13 11 11 2
7 1 10 9 13 10 9 2
6 15 13 10 9 0 2
9 15 13 10 9 1 10 9 11 2
5 15 13 11 11 2
5 15 13 11 11 2
5 15 13 11 11 2
5 15 13 11 11 2
6 15 13 11 1 11 2
5 15 13 11 11 2
5 15 13 11 11 2
8 10 15 13 10 11 11 11 2
6 10 15 13 10 11 2
6 10 15 13 10 11 2
6 10 15 13 10 11 2
7 3 4 13 10 11 11 2
15 10 9 9 1 10 11 4 3 13 1 2 10 9 2 2
9 3 4 4 13 10 11 1 11 2
8 15 13 10 9 1 10 11 2
11 1 10 9 4 4 13 10 11 11 11 2
6 15 13 10 9 11 2
17 15 13 10 9 1 10 15 4 4 13 10 9 11 1 10 9 2
16 15 13 10 9 15 13 10 11 11 1 10 11 1 10 11 2
13 10 9 13 16 10 2 11 2 15 13 7 13 2
8 1 10 9 15 13 10 11 2
9 15 4 13 10 0 9 1 11 2
14 10 9 13 9 1 10 9 1 10 2 11 11 2 2
17 10 9 1 9 0 4 13 10 11 1 10 9 1 10 10 9 2
8 3 13 10 9 1 10 11 2
8 15 13 10 9 1 10 11 2
9 15 13 10 9 1 10 11 11 2
11 1 10 9 1 10 11 15 13 10 9 2
8 15 4 13 10 9 1 11 2
11 10 9 13 1 11 1 10 9 1 11 2
9 10 9 0 13 1 10 11 11 2
11 3 15 13 10 9 7 9 1 10 11 2
13 10 9 13 1 10 9 1 10 9 2 11 2 2
8 13 10 9 13 1 11 11 2
11 10 9 4 13 1 10 11 1 10 9 2
7 3 4 4 13 10 11 2
10 15 13 10 11 1 10 11 11 11 2
13 10 9 1 9 13 10 9 15 13 10 11 0 2
7 10 15 13 10 9 11 2
5 3 13 10 11 2
10 15 13 10 9 1 10 9 1 11 2
5 3 15 13 11 2
9 1 10 9 0 13 10 11 11 2
13 10 9 0 1 11 12 13 10 9 0 11 11 2
7 15 13 10 9 1 11 2
5 10 9 13 11 2
13 1 10 9 4 4 13 10 11 11 1 10 11 2
15 15 13 10 9 0 1 10 2 9 1 10 9 0 2 2
8 3 15 13 10 11 11 0 2
8 1 10 15 13 10 9 11 2
6 10 9 13 10 11 2
13 1 10 9 4 13 10 9 1 9 0 7 0 2
15 10 9 13 11 16 10 9 0 13 1 11 1 10 12 2
8 3 4 13 10 0 9 0 2
10 15 13 10 9 9 1 10 11 11 2
9 10 9 13 10 11 1 10 12 2
18 10 11 11 13 10 9 1 9 1 9 1 9 1 10 11 1 11 2
8 1 10 9 4 13 10 11 2
11 10 9 0 13 1 10 9 1 12 9 2
6 3 4 13 11 11 2
6 10 9 13 11 11 2
8 15 13 10 9 1 11 11 2
8 15 13 10 9 1 10 11 2
8 15 4 13 2 11 11 2 2
7 3 13 10 2 11 2 2
10 1 10 9 13 10 9 2 11 2 2
11 15 13 10 9 1 10 11 1 10 11 2
10 1 10 9 0 15 13 10 11 11 2
9 1 10 9 15 13 10 11 11 2
9 1 10 9 13 11 11 11 11 2
15 10 9 4 13 10 9 1 10 11 1 10 11 1 11 2
7 1 15 13 10 9 0 2
5 10 9 13 11 2
9 3 15 13 10 9 0 0 0 2
9 10 9 13 1 10 9 1 11 2
9 3 15 13 10 9 1 11 11 2
9 3 15 13 10 9 1 11 11 2
9 3 15 13 10 9 1 10 11 2
8 15 13 10 9 1 10 11 2
6 3 4 13 11 11 2
10 3 4 13 10 9 1 10 12 9 2
12 1 10 9 1 10 9 15 13 10 9 0 2
16 10 9 13 9 1 10 9 1 10 11 1 10 9 1 11 2
11 3 10 11 11 4 13 10 9 1 11 2
9 1 10 9 0 15 13 11 11 2
8 15 13 10 9 1 10 11 2
13 1 10 9 1 9 1 9 4 13 1 10 9 2
12 15 4 4 13 10 3 0 9 1 10 9 2
9 15 13 10 9 1 9 1 11 2
12 1 10 9 4 4 13 10 9 1 10 9 2
13 1 10 9 13 10 9 1 10 9 2 11 2 2
6 15 13 10 9 0 2
12 10 11 11 0 13 10 11 11 1 10 12 2
10 15 4 13 10 0 9 1 10 11 2
6 10 9 13 10 11 2
9 1 10 9 13 10 9 0 11 2
15 15 13 10 9 0 1 10 3 0 9 1 9 1 9 2
11 15 4 13 10 9 1 9 0 11 11 2
8 15 13 10 9 1 10 11 2
8 15 13 10 9 1 10 11 2
17 10 9 1 10 9 4 13 1 10 9 1 10 9 2 11 2 2
8 15 13 10 9 1 11 11 2
7 1 10 9 13 9 11 2
11 1 10 9 15 13 10 11 1 10 11 2
10 13 10 9 1 10 9 1 10 11 2
12 15 13 10 9 1 10 11 1 10 11 11 2
8 15 4 13 10 9 1 11 2
10 15 4 13 10 2 11 1 11 2 2
9 10 9 4 13 10 11 1 9 2
10 15 13 10 9 1 2 9 0 2 2
7 13 10 9 1 11 11 2
8 3 4 13 10 0 9 0 2
7 10 15 13 10 9 11 2
13 15 13 10 9 1 10 9 1 10 11 1 9 2
10 1 10 9 4 4 13 10 11 11 2
9 10 9 0 13 10 9 1 11 2
7 1 10 9 15 13 11 2
10 3 15 13 10 9 1 9 0 0 2
12 1 10 9 15 13 10 9 0 2 11 2 2
5 3 15 13 11 2
6 10 9 13 10 11 2
10 1 10 11 11 4 4 13 11 11 2
8 15 13 10 9 1 10 11 2
23 10 9 13 10 9 1 10 9 11 11 2 11 11 2 1 10 11 1 10 11 1 11 2
9 15 13 10 9 1 10 9 0 2
9 10 9 0 0 4 13 10 9 2
9 1 10 9 13 10 2 11 2 2
5 13 10 9 0 2
7 3 15 13 10 9 11 2
7 10 15 13 10 9 11 2
6 15 13 10 9 11 2
17 3 15 4 13 10 9 0 1 10 11 1 10 11 1 10 11 2
9 10 9 4 13 10 9 0 11 2
10 1 10 9 4 13 10 9 1 11 2
11 15 4 13 2 10 9 1 10 9 2 2
7 10 11 11 4 13 11 2
6 3 15 13 10 11 2
9 10 9 4 13 10 13 13 0 2
7 1 10 9 13 11 11 2
8 15 13 1 10 9 1 11 2
8 15 13 10 9 1 10 11 2
9 3 4 4 13 10 0 11 11 2
11 3 15 13 10 9 1 10 11 11 0 2
6 10 9 13 10 11 2
10 1 10 9 4 13 0 10 11 11 2
12 10 11 4 13 1 10 9 2 11 12 2 2
11 10 9 13 1 10 11 11 1 10 11 2
7 15 13 10 11 11 0 2
10 3 15 13 10 9 1 11 11 11 2
12 1 10 9 15 13 10 9 1 10 11 11 2
9 1 10 9 13 10 9 1 9 2
8 3 4 13 10 11 1 11 2
12 1 10 9 10 11 4 13 1 10 11 11 2
9 3 15 13 10 11 1 10 11 2
9 15 13 10 9 1 10 11 11 2
9 15 4 13 13 10 9 1 11 2
13 15 13 10 9 1 9 1 10 9 1 11 11 2
5 3 15 13 11 2
9 3 15 13 10 9 1 10 9 2
6 10 9 13 10 9 2
9 1 10 9 15 13 11 7 11 2
6 15 13 10 9 0 2
7 15 13 10 9 1 11 2
11 1 10 9 15 13 10 0 9 1 9 2
14 15 13 10 9 1 10 9 11 2 11 1 10 9 2
11 15 13 10 9 1 10 11 1 10 11 2
5 10 9 13 11 2
10 3 15 13 10 9 0 1 11 11 2
8 15 13 10 9 1 10 11 2
8 10 9 4 13 10 11 11 2
16 10 15 4 13 10 9 1 10 9 1 10 9 0 1 11 2
11 1 10 9 15 13 10 11 1 10 11 2
11 15 13 10 9 1 10 11 1 10 11 2
21 10 9 4 13 1 9 1 10 9 1 9 1 10 9 1 10 9 2 11 2 2
13 11 11 11 11 13 10 9 1 10 9 1 9 2
17 1 10 9 4 13 1 10 9 1 11 1 10 11 11 11 11 2
9 15 13 10 9 1 10 11 11 2
11 15 13 10 9 1 10 9 1 10 11 2
9 13 10 9 0 13 1 10 9 2
8 15 13 10 9 1 10 11 2
8 15 13 10 9 1 10 11 2
7 10 15 13 10 9 11 2
10 15 13 10 9 0 1 10 11 11 2
14 1 10 9 15 13 1 9 10 2 11 1 11 2 2
15 15 13 10 9 1 10 9 1 9 1 10 11 1 11 2
5 3 13 11 11 2
8 1 10 11 4 13 11 11 2
10 10 0 9 0 4 4 13 1 9 2
8 3 15 13 10 9 0 0 2
9 15 13 10 11 1 10 11 11 2
13 10 9 0 4 13 1 10 0 9 0 1 11 2
9 10 9 13 10 11 1 10 11 2
8 10 9 4 13 1 11 11 2
10 3 13 10 11 3 1 10 10 9 2
5 3 13 11 11 2
8 10 9 15 13 1 10 9 2
19 15 4 13 10 9 1 10 9 0 1 10 11 1 11 11 1 10 12 2
8 10 9 1 9 13 11 11 2
7 3 13 10 0 11 11 2
11 10 15 13 10 2 9 15 15 13 2 2
6 3 13 0 10 11 2
12 15 13 10 9 1 2 10 11 11 11 2 2
15 15 13 10 0 9 1 10 2 9 1 10 9 0 2 2
9 10 9 1 11 11 4 13 11 2
9 15 13 10 9 0 1 10 11 2
6 1 3 13 11 11 2
12 15 13 10 0 9 1 10 2 9 11 2 2
7 1 10 9 13 11 11 2
6 10 9 13 11 11 2
12 10 0 9 15 13 1 11 1 10 0 9 2
10 15 13 10 9 0 1 10 9 11 2
7 3 13 10 9 11 11 2
10 15 13 10 9 3 0 1 10 11 2
8 1 10 15 4 13 10 9 2
13 15 13 10 9 1 9 1 10 9 1 11 11 2
10 1 10 9 13 10 9 11 7 11 2
11 15 4 13 10 9 1 9 2 11 2 2
5 10 9 13 11 2
5 3 13 11 11 2
9 3 13 1 10 9 0 11 11 2
14 1 10 11 4 13 10 9 2 11 1 10 11 2 2
10 15 13 10 0 9 1 10 11 11 2
6 10 9 13 10 11 2
10 10 11 13 1 10 11 1 11 11 2
8 10 15 13 2 9 9 2 2
11 1 10 9 13 10 9 1 10 11 11 2
17 1 9 2 10 9 4 13 10 9 9 1 10 11 1 11 11 2
9 3 4 13 10 11 1 10 11 2
8 10 9 4 13 1 11 11 2
7 1 10 9 13 11 11 2
5 13 10 9 0 2
14 1 10 11 4 13 1 13 1 10 11 11 10 9 2
7 3 10 11 13 10 9 2
10 3 4 13 10 11 1 10 11 11 2
8 10 9 13 11 11 16 13 2
9 3 15 13 10 9 1 11 11 2
15 10 9 4 13 1 1 10 12 1 10 11 11 1 11 2
13 10 9 0 1 9 13 1 11 11 1 10 12 2
7 3 15 13 10 9 11 2
9 3 4 13 10 11 11 1 11 2
11 3 4 4 13 10 11 11 1 10 12 2
10 15 13 10 9 1 10 9 1 11 2
12 15 13 10 9 0 1 10 9 2 11 2 2
8 15 13 10 9 1 10 11 2
14 3 15 4 13 10 0 9 1 10 9 1 11 11 2
14 3 15 13 10 9 0 13 1 10 9 1 10 11 2
8 10 9 13 11 11 16 13 2
12 15 13 10 9 1 10 9 0 0 11 11 2
10 10 0 4 13 1 11 1 10 12 2
13 15 13 10 9 1 10 11 11 1 10 11 11 2
16 1 10 9 1 10 0 1 11 13 10 9 1 10 9 9 2
11 15 13 10 9 1 10 11 1 10 11 2
8 15 13 10 9 1 10 11 2
11 15 13 10 9 1 10 9 0 11 11 2
13 3 10 9 9 11 11 13 10 9 1 10 9 2
10 3 4 13 10 9 0 1 10 11 2
7 3 13 10 9 11 11 2
7 13 10 9 1 11 11 2
9 3 15 13 10 0 9 0 0 2
18 15 4 13 10 9 1 9 1 10 9 1 10 11 11 1 10 12 2
9 3 15 13 10 9 1 11 11 2
5 3 13 11 11 2
13 10 9 0 15 13 1 10 11 11 1 10 12 2
7 13 10 9 13 1 11 2
8 3 4 13 10 9 1 11 2
8 1 10 9 11 13 10 9 2
6 13 10 9 0 0 2
9 10 9 4 4 13 1 11 11 2
5 3 13 11 11 2
13 1 10 9 15 13 13 10 9 0 1 11 11 2
16 1 10 9 10 9 0 1 10 11 0 4 13 1 11 11 2
16 1 10 9 4 4 13 10 9 1 10 15 9 11 11 11 2
11 15 13 10 0 9 1 11 11 11 11 2
9 1 10 9 1 9 13 11 11 2
8 3 4 13 10 2 11 2 2
8 1 10 9 4 13 10 11 2
14 15 13 10 9 1 10 0 9 1 15 4 13 11 2
8 1 10 9 0 13 11 11 2
7 3 11 13 10 11 11 2
8 3 4 13 10 9 1 11 2
11 10 9 1 10 11 3 13 10 9 0 2
13 10 9 4 13 10 9 1 10 11 11 1 11 2
10 15 13 10 9 3 0 1 10 11 2
8 10 9 13 11 11 16 13 2
7 15 13 10 11 11 0 2
10 1 10 9 11 11 11 13 10 9 2
12 1 10 0 9 4 13 10 11 11 1 11 2
8 15 4 13 9 1 10 11 2
12 10 9 0 4 13 1 11 11 1 10 12 2
12 15 13 0 10 9 1 10 9 1 11 11 2
5 10 9 13 11 2
7 15 13 10 0 9 0 2
12 1 10 9 11 11 13 10 11 11 1 11 2
9 10 15 13 10 9 2 11 2 2
15 15 13 10 9 1 10 0 9 1 10 9 1 11 11 2
12 15 13 10 9 1 10 15 9 1 10 11 2
7 1 10 9 13 11 11 2
9 1 10 9 15 13 10 11 11 2
8 10 9 13 0 10 11 11 2
14 10 9 4 13 1 10 9 1 11 11 1 10 12 2
8 1 10 9 4 13 11 11 2
8 1 10 9 4 13 11 11 2
7 10 15 13 10 9 11 2
11 1 10 9 11 11 13 1 10 9 11 2
12 10 9 13 10 9 1 11 10 9 1 11 2
6 10 9 13 11 11 2
11 1 10 9 10 11 13 9 1 10 11 2
8 15 4 13 2 11 11 2 2
10 15 4 13 10 11 11 1 10 12 2
9 1 10 9 11 11 15 13 9 2
10 10 9 0 13 10 0 9 1 9 2
6 3 10 11 13 11 2
14 15 13 10 0 9 3 0 1 10 11 11 11 11 2
5 3 13 11 11 2
11 15 13 10 9 0 1 9 1 10 12 2
6 1 10 9 13 11 2
7 10 15 13 10 9 11 2
8 15 13 10 9 1 10 11 2
5 3 13 11 11 2
10 3 15 13 10 0 11 1 10 11 2
13 1 15 4 13 10 9 1 9 9 12 1 11 2
11 3 15 13 10 9 1 10 9 11 11 2
9 3 13 10 9 11 11 11 11 2
13 10 9 13 10 0 0 9 1 9 1 10 9 2
11 3 13 10 9 1 10 9 1 10 9 2
9 15 4 13 10 9 1 10 11 2
10 15 13 10 9 1 9 1 10 11 2
15 10 9 0 4 13 1 10 11 1 10 11 1 10 12 2
7 1 15 4 13 11 11 2
8 10 9 0 4 13 11 11 2
8 15 4 13 10 2 11 2 2
9 11 11 13 10 9 1 10 9 2
13 3 15 13 10 9 0 13 1 2 11 12 2 2
15 10 9 4 13 1 3 10 9 2 11 2 1 11 11 2
14 1 10 9 13 10 9 0 13 1 10 11 1 11 2
9 10 9 13 9 13 10 0 11 2
11 15 13 10 9 1 10 9 0 1 11 2
14 15 13 10 9 1 10 9 0 1 10 11 11 11 2
12 15 13 10 9 1 10 9 1 10 9 0 2
7 3 4 13 11 11 11 2
9 10 11 13 1 10 9 1 11 2
6 13 10 9 1 11 2
5 3 13 11 11 2
7 10 9 4 13 11 11 2
6 10 9 13 11 11 2
10 15 13 10 11 11 1 10 11 11 2
15 1 10 9 15 13 10 11 1 10 11 11 1 10 11 2
6 13 10 9 0 0 2
10 3 15 13 10 11 11 1 10 11 2
10 15 13 10 0 9 13 1 11 11 2
8 15 4 13 10 9 0 11 2
6 15 4 13 10 9 2
10 3 4 13 10 0 9 1 11 11 2
19 15 4 13 2 13 1 11 10 10 9 7 1 10 11 10 10 9 2 2
10 15 13 10 0 9 1 11 11 11 2
10 3 11 11 13 2 10 11 11 2 2
11 10 9 4 13 10 9 1 13 9 0 2
5 10 9 13 11 2
7 10 9 13 0 1 11 2
8 15 13 10 9 1 10 11 2
10 1 10 9 15 13 10 9 1 9 2
7 3 4 13 11 11 11 2
12 3 13 10 9 15 13 10 9 1 11 11 2
12 1 10 15 4 13 10 9 2 11 11 2 2
13 3 4 4 13 10 11 11 1 10 11 1 9 2
13 10 9 13 10 0 9 1 9 0 1 10 9 2
14 15 13 10 9 3 0 15 4 4 13 1 10 9 2
8 15 13 10 9 1 10 11 2
14 10 9 1 0 9 13 10 9 1 10 9 11 11 2
8 15 13 10 9 1 10 11 2
7 10 9 4 13 11 11 2
9 15 13 10 11 11 1 10 11 2
11 1 10 9 4 13 10 9 1 10 9 2
7 1 15 4 13 11 11 2
14 3 15 13 10 9 15 4 13 10 0 9 1 11 2
12 3 0 9 0 13 1 10 9 10 12 9 2
6 3 4 13 10 9 2
9 15 13 10 9 1 10 9 0 2
9 1 10 9 11 11 13 12 9 2
8 3 4 13 10 9 1 9 2
7 10 9 13 10 9 0 2
8 10 9 15 13 1 10 9 2
10 3 15 13 10 9 1 11 7 11 2
9 1 10 9 0 13 9 11 11 2
15 10 9 0 1 9 7 9 4 13 1 2 11 11 2 2
6 10 9 13 9 0 2
8 10 9 0 13 10 9 11 2
8 15 13 10 9 1 10 11 2
11 10 9 4 13 2 9 1 10 11 2 2
11 3 13 0 10 0 9 1 10 9 11 2
10 3 13 10 0 9 16 13 1 9 2
6 3 4 13 11 14 2
15 15 13 10 0 9 1 13 10 9 1 15 1 12 9 2
7 3 15 13 10 9 11 2
9 1 10 9 10 11 13 10 9 2
7 15 13 0 10 11 11 2
9 3 11 11 13 10 9 1 11 2
17 10 12 9 0 4 13 1 10 9 1 10 11 11 1 10 11 2
8 15 13 10 9 1 10 11 2
11 15 13 10 9 1 0 9 1 10 12 2
8 15 13 10 9 1 10 11 2
8 15 13 10 9 1 10 11 2
11 15 4 13 10 0 9 0 1 10 9 2
13 15 4 13 10 9 11 1 10 9 1 10 12 2
9 3 15 13 10 9 1 11 11 2
15 10 9 13 13 1 4 15 13 1 10 11 1 10 11 2
10 15 4 13 1 2 11 11 11 2 2
8 3 13 10 11 1 10 11 2
10 15 13 10 9 1 10 9 3 0 2
8 1 3 13 11 1 10 12 2
9 10 9 13 10 9 1 10 11 2
9 3 15 13 10 9 1 11 11 2
6 3 13 10 9 11 2
7 15 13 0 10 11 11 2
10 15 13 10 9 3 0 1 10 9 2
10 15 13 10 9 0 1 10 0 9 2
6 3 4 13 11 11 2
11 10 9 13 9 1 10 11 1 11 11 2
8 3 13 10 9 1 11 11 2
5 3 13 11 11 2
8 15 13 10 9 1 10 11 2
9 3 15 13 10 9 1 10 9 2
6 10 9 13 11 11 2
11 10 9 0 13 10 3 0 9 1 9 2
10 10 9 4 13 1 10 9 1 9 2
8 10 9 13 10 9 0 0 2
8 10 9 0 4 13 11 11 2
10 3 15 13 10 9 1 2 11 2 2
9 15 13 10 9 0 1 10 11 2
15 3 15 13 10 9 1 10 9 1 9 2 11 11 2 2
17 10 9 1 9 4 13 1 10 9 11 1 10 9 1 10 12 2
12 3 15 13 10 3 0 9 1 10 11 11 2
8 15 13 10 9 0 9 0 2
10 15 13 10 9 1 2 11 11 2 2
7 10 9 13 10 9 11 2
6 15 13 0 11 11 2
10 1 10 9 10 11 11 13 10 9 2
13 16 15 15 4 13 2 1 10 9 15 4 13 2
8 3 13 10 9 11 11 11 2
7 3 13 10 9 11 11 2
6 15 13 0 10 9 2
9 3 15 13 2 9 2 1 0 2
10 15 13 10 9 3 0 1 10 11 2
11 15 13 10 0 9 1 13 10 11 11 2
9 15 13 10 9 0 1 10 9 2
10 1 10 15 4 13 10 9 1 9 2
13 3 15 13 10 9 1 2 3 1 10 9 2 2
8 15 4 13 2 10 11 2 2
9 15 13 10 0 9 1 10 11 2
8 15 13 10 9 1 10 11 2
10 1 10 9 1 10 11 15 13 11 2
7 10 9 4 13 11 11 2
14 15 13 10 9 9 1 10 2 9 1 12 9 2 2
7 3 13 10 9 11 11 2
8 15 13 10 9 1 11 11 2
21 15 13 10 9 1 10 9 1 9 0 1 11 11 2 1 10 11 1 10 11 2
8 1 10 9 15 13 10 11 2
10 15 13 10 9 1 10 9 1 11 2
9 3 15 13 10 9 1 11 11 2
10 10 9 13 11 11 16 13 1 9 2
5 3 13 11 11 2
23 15 13 2 10 9 13 10 9 2 10 9 13 10 9 7 10 12 3 15 13 3 2 2
8 3 13 10 9 1 11 11 2
7 1 10 9 15 13 11 2
14 15 13 10 9 0 3 1 2 11 11 11 11 2 2
6 10 9 13 11 11 2
13 1 10 9 0 10 9 13 10 0 9 1 9 2
7 3 15 13 10 11 11 2
14 15 1 10 9 0 1 10 11 11 13 1 9 0 2
9 1 10 9 4 13 10 9 11 2
11 15 13 10 0 9 3 0 1 10 9 2
8 3 15 13 10 11 1 11 2
7 10 9 15 13 1 11 2
9 3 15 13 10 9 1 11 11 2
9 3 15 13 10 9 1 11 11 2
8 15 13 10 9 1 11 11 2
8 3 13 10 9 1 11 11 2
15 15 13 2 10 9 13 10 9 1 13 10 9 0 2 2
8 10 9 13 10 10 9 0 2
11 15 13 10 9 0 1 11 2 1 11 2
10 15 13 10 9 3 0 1 10 11 2
10 15 13 10 0 9 1 10 9 11 2
8 1 10 15 13 10 9 11 2
9 15 13 10 9 0 1 10 11 2
9 1 10 9 11 11 13 1 11 2
6 3 13 11 11 11 2
8 15 13 10 9 1 10 11 2
10 1 10 9 11 11 13 1 10 9 2
14 3 15 13 10 9 15 13 10 9 1 10 11 11 2
13 15 13 10 9 1 10 9 0 1 10 11 11 2
13 3 15 13 10 9 1 9 3 13 10 11 11 2
6 10 9 13 11 11 2
9 15 13 10 9 1 10 9 0 2
9 3 13 10 9 1 10 12 9 2
5 3 13 11 11 2
13 15 13 10 3 0 9 1 9 13 1 10 9 2
7 10 15 13 10 9 11 2
11 15 13 10 9 1 10 9 0 1 11 2
10 15 4 13 10 9 2 11 11 2 2
10 1 3 12 9 4 13 3 10 9 2
7 15 13 10 2 11 2 2
10 3 1 10 9 15 13 10 11 11 2
8 10 9 0 15 13 1 11 2
11 15 13 10 0 9 11 1 2 11 2 2
9 15 13 10 9 13 1 11 11 2
9 15 13 10 9 3 0 1 11 2
13 10 9 15 13 1 10 9 1 10 9 1 9 2
10 3 15 13 10 9 0 0 1 11 2
7 3 15 13 10 9 9 2
12 1 10 9 4 13 10 9 2 11 11 2 2
9 15 13 10 9 0 1 10 9 2
13 10 9 13 10 11 15 13 1 10 11 11 11 2
11 15 13 10 9 3 1 9 1 10 11 2
7 10 15 13 10 9 11 2
6 10 9 13 11 11 2
7 15 13 10 9 11 11 2
9 15 13 10 9 0 1 10 9 2
9 3 15 13 10 9 11 1 11 2
8 1 10 9 13 0 11 11 2
9 15 13 10 0 9 1 10 9 2
10 15 13 13 10 9 1 10 11 11 2
12 1 10 9 1 11 9 11 13 10 10 9 2
10 15 13 10 0 9 0 1 11 11 2
11 3 4 13 10 0 9 1 10 9 0 2
7 3 13 10 11 11 0 2
9 3 13 10 11 11 1 10 11 2
8 15 13 10 9 1 11 11 2
11 10 0 9 0 13 1 10 11 11 11 2
10 3 4 13 10 9 11 11 1 11 2
8 10 9 13 11 11 16 13 2
8 3 13 10 11 1 10 11 2
10 15 13 10 9 0 1 13 1 11 2
8 3 9 15 13 1 10 9 2
9 1 15 13 10 9 1 10 11 2
8 15 13 10 9 1 10 11 2
13 3 13 10 10 0 9 1 9 10 2 11 2 2
10 15 13 10 9 1 9 1 10 11 2
11 15 13 10 9 3 0 1 10 11 11 2
19 1 10 9 1 11 13 10 9 2 10 0 0 9 1 9 7 3 2 2
6 15 13 0 10 11 2
9 10 9 13 10 0 9 1 9 2
11 3 15 13 10 9 1 15 13 9 0 2
6 15 13 0 10 9 2
10 3 4 13 10 9 1 10 9 0 2
11 3 4 13 11 11 11 9 1 10 11 2
9 15 13 10 9 3 13 1 11 2
8 3 4 13 10 9 11 11 2
7 3 4 13 10 11 12 2
21 15 13 10 0 9 1 13 10 11 1 11 2 1 11 7 9 1 10 0 9 2
5 15 13 10 9 2
6 3 4 13 10 11 2
11 10 9 1 10 9 0 13 1 10 11 2
16 3 0 9 1 11 11 4 13 1 10 9 7 13 1 11 2
5 10 9 13 11 2
11 1 10 9 11 13 1 10 9 1 11 2
10 3 15 13 10 9 0 1 11 11 2
9 15 13 10 9 0 1 10 11 2
7 10 9 0 13 10 11 2
10 15 13 10 9 1 9 9 3 13 2
11 3 15 13 11 11 11 1 10 11 11 2
6 1 10 15 13 11 2
9 10 9 13 16 13 1 10 9 2
10 15 13 10 9 1 9 1 10 9 2
15 15 13 10 0 9 1 9 1 10 9 1 10 9 0 2
10 15 13 10 9 13 1 10 0 9 2
10 15 13 10 9 1 11 1 10 11 2
9 3 1 9 4 13 10 9 0 2
7 3 4 0 9 11 11 2
7 15 13 10 9 1 11 2
10 15 13 10 9 3 0 1 10 11 2
8 3 13 10 9 1 11 11 2
12 3 15 13 10 9 1 10 9 1 10 11 2
6 3 4 13 10 9 2
12 10 9 1 10 9 13 12 9 1 10 12 2
17 1 10 9 15 13 10 0 9 1 11 1 10 9 1 10 11 2
14 3 15 13 10 9 13 1 10 11 1 11 7 11 2
9 15 13 10 11 11 1 11 11 2
9 1 10 9 13 2 11 11 2 2
10 15 13 10 9 3 0 1 10 9 2
11 15 13 10 0 9 1 9 1 11 11 2
13 15 15 4 13 1 10 9 0 1 10 9 0 2
10 15 13 0 10 9 0 1 10 11 2
6 3 4 13 11 11 2
6 3 4 13 10 9 2
8 15 13 10 9 1 10 11 2
8 10 9 15 13 1 10 9 2
11 15 13 10 9 0 3 0 1 10 9 2
6 10 9 13 10 11 2
8 3 4 13 10 9 1 11 2
14 3 15 13 10 9 1 12 9 13 3 1 10 9 2
7 10 9 0 13 9 0 2
19 10 9 13 10 9 1 11 11 1 10 9 2 11 11 2 1 10 12 2
6 15 4 13 10 11 2
11 1 3 4 13 10 10 9 10 11 11 2
8 3 15 13 10 9 1 9 2
6 15 4 13 11 11 2
7 3 13 11 1 10 11 2
8 3 4 13 10 0 9 0 2
8 1 10 9 15 13 10 11 2
13 10 15 13 10 9 11 1 10 9 1 10 9 2
8 1 10 9 13 10 9 11 2
9 1 10 9 15 13 11 2 11 2
10 15 13 10 0 9 1 10 11 11 2
11 3 13 10 11 11 1 10 11 11 11 2
11 3 15 13 10 11 11 11 5 11 11 2
5 3 13 11 11 2
12 10 9 4 13 10 9 2 1 9 0 2 2
10 3 13 10 11 10 11 1 10 11 2
7 1 10 9 13 11 11 2
5 3 13 11 11 2
9 15 13 10 0 9 1 11 11 2
9 10 15 13 2 11 11 11 2 2
9 3 4 13 11 1 10 9 11 2
11 3 4 13 10 9 15 13 9 1 9 2
10 15 13 10 0 9 1 13 10 9 2
9 3 13 11 11 1 10 11 11 2
10 3 15 13 10 9 0 0 1 11 2
10 15 13 10 9 1 10 9 1 11 2
12 15 13 10 3 0 9 0 1 10 11 11 2
7 15 13 0 10 11 11 2
13 15 13 10 9 1 10 11 1 10 11 1 11 2
7 3 15 13 10 11 11 2
13 10 9 9 0 13 10 0 9 1 9 1 9 2
12 1 10 9 1 10 9 10 9 0 15 13 2
10 1 10 9 11 11 13 1 10 11 2
10 10 9 13 10 9 2 11 11 2 2
8 3 4 13 10 9 1 11 2
5 3 13 11 11 2
11 15 13 10 9 1 10 11 1 10 12 2
8 15 13 10 9 1 10 11 2
7 1 10 9 13 11 11 2
7 3 13 11 11 11 11 2
15 1 10 9 4 3 13 10 9 1 9 0 11 11 11 2
11 1 10 9 1 9 15 13 3 12 9 2
11 15 13 10 9 3 0 1 10 11 11 2
7 15 13 10 9 0 0 2
9 10 9 13 10 9 1 10 11 2
9 1 10 9 4 13 10 11 11 2
16 1 10 9 15 13 1 10 9 2 9 1 10 0 9 2 2
7 10 15 13 10 9 11 2
11 3 4 13 10 9 2 3 1 9 2 2
9 15 13 0 10 11 11 1 11 2
9 1 10 9 10 11 13 10 9 2
11 1 10 9 13 10 9 11 1 11 11 2
6 3 4 13 10 9 2
5 3 13 11 11 2
9 1 10 9 15 13 10 9 11 2
8 3 15 13 10 11 1 11 2
7 3 4 13 10 9 11 2
15 1 15 13 10 9 0 2 10 9 13 10 0 9 2 2
8 15 13 10 9 0 1 9 2
7 1 15 15 13 10 9 2
12 15 13 10 9 1 9 1 10 9 0 11 2
17 3 15 13 10 9 1 10 9 1 10 9 13 1 10 9 11 2
10 3 13 10 9 1 10 9 11 11 2
14 15 13 10 9 13 1 15 13 1 10 9 1 9 2
9 15 13 10 9 1 10 9 0 2
7 3 4 13 10 0 9 2
8 15 4 13 10 9 1 13 2
10 10 15 13 10 9 1 10 9 12 2
14 1 10 9 1 10 11 15 13 10 11 1 10 11 2
9 10 9 11 4 13 1 10 9 2
10 15 13 10 0 9 1 10 11 11 2
16 15 13 10 0 9 1 10 9 1 13 10 9 1 10 9 2
7 3 4 13 10 11 11 2
7 3 13 11 1 10 11 2
13 16 10 9 1 9 4 13 2 15 13 10 9 2
15 1 10 9 3 13 10 9 1 10 9 1 10 9 9 2
9 1 10 9 13 10 9 11 11 2
7 15 13 10 9 1 11 2
8 15 13 15 1 10 9 0 2
8 3 13 10 9 11 11 11 2
10 3 15 13 10 9 1 10 9 0 2
7 10 15 13 10 9 11 2
10 3 13 1 10 0 9 10 11 11 2
8 3 15 13 10 9 1 11 2
9 15 13 10 0 9 1 11 11 2
13 10 15 10 9 0 13 10 9 0 1 10 9 2
11 15 13 10 0 9 1 10 9 1 11 2
11 15 13 10 9 1 9 1 10 9 0 2
9 1 10 9 15 13 10 11 11 2
10 1 10 9 1 10 9 13 10 9 2
8 15 13 13 10 9 10 9 2
7 3 4 13 10 9 11 2
10 15 13 10 9 0 1 10 9 11 2
9 1 10 15 4 13 10 11 11 2
11 10 9 15 13 1 10 9 2 11 2 2
6 3 13 10 9 0 2
14 10 9 13 10 3 0 9 1 9 1 10 11 11 2
8 10 9 0 4 13 10 11 2
8 1 10 15 4 13 10 9 2
6 15 4 13 11 11 2
8 3 4 13 10 11 11 11 2
9 3 15 13 10 13 1 11 11 2
6 3 4 13 10 11 2
8 15 13 10 9 1 10 11 2
10 3 15 13 10 9 0 1 11 11 2
9 3 15 13 10 9 1 11 11 2
15 3 4 13 1 11 11 10 9 1 10 9 1 10 11 2
10 3 15 13 10 11 1 10 11 11 2
9 10 9 13 10 9 0 11 11 2
11 3 13 10 9 1 10 9 1 11 11 2
9 3 15 13 10 9 1 11 11 2
10 15 13 10 2 9 1 10 9 2 2
9 15 13 2 9 1 10 9 2 2
12 10 9 0 4 13 1 11 11 1 10 12 2
5 10 9 13 11 2
7 15 13 10 9 0 0 2
8 3 4 13 10 0 11 11 2
8 1 10 9 0 13 11 11 2
8 1 15 13 10 11 11 11 2
13 15 13 10 3 0 9 13 1 11 11 2 11 2
5 3 13 10 11 2
6 15 4 13 10 9 2
11 15 13 10 3 0 9 0 1 11 11 2
7 10 15 13 10 9 11 2
10 1 10 9 4 13 10 0 9 0 2
11 15 4 13 11 11 1 2 11 11 2 2
6 3 4 13 11 11 2
10 15 13 10 9 3 0 1 10 11 2
15 15 13 10 0 9 1 9 9 1 10 9 1 9 0 2
9 1 10 9 13 2 11 11 2 2
12 15 13 10 0 9 1 13 15 1 10 9 2
9 1 10 9 4 13 10 9 11 2
9 15 13 10 9 0 1 10 9 2
6 3 13 10 9 11 2
14 15 4 13 10 9 0 15 11 11 13 1 10 9 2
9 3 13 10 9 1 11 11 11 2
5 15 13 10 9 2
11 15 13 10 9 1 10 9 1 11 11 2
12 1 10 9 15 13 10 9 0 1 10 11 2
6 3 13 3 10 11 2
13 15 13 10 9 13 1 9 3 0 1 10 9 2
10 15 13 10 9 3 0 1 10 9 2
8 1 10 9 13 10 9 9 2
5 3 13 11 11 2
8 1 10 9 15 13 10 11 2
13 15 13 10 9 1 9 0 1 10 9 1 11 2
11 10 9 13 1 9 13 9 1 10 9 2
12 3 15 13 10 9 3 0 1 10 9 0 2
6 15 13 0 11 11 2
10 3 11 11 11 13 10 9 1 9 2
12 15 4 13 9 1 10 11 11 1 10 12 2
9 3 4 13 10 0 9 1 9 2
8 10 9 4 13 10 11 12 2
11 10 9 13 10 11 11 1 10 11 11 2
10 3 4 13 10 11 1 11 1 11 2
10 3 4 13 1 10 0 9 10 9 2
11 3 4 13 10 0 9 1 10 11 11 2
9 10 9 13 0 1 10 0 9 2
10 15 13 10 0 9 0 1 10 11 2
14 15 13 10 9 0 1 4 13 9 1 10 11 11 2
11 15 13 10 0 9 1 13 1 10 9 2
5 3 13 11 11 2
6 3 15 13 11 11 2
9 3 15 13 10 9 1 10 11 2
11 15 13 10 9 15 13 10 11 11 11 2
8 15 13 10 9 1 10 11 2
14 10 9 10 9 13 13 1 9 9 1 10 9 11 2
8 1 10 9 13 10 11 12 2
16 10 9 4 13 10 0 9 1 10 0 9 1 10 11 11 2
8 3 4 13 10 9 1 11 2
9 15 13 10 9 0 1 10 11 2
11 15 13 0 10 9 1 10 11 1 11 2
10 1 10 9 15 13 10 11 1 11 2
12 3 15 13 10 0 9 0 1 11 7 11 2
11 15 13 11 11 1 10 9 1 10 9 2
6 15 13 0 11 11 2
11 10 9 13 12 9 1 9 1 13 11 2
9 15 13 10 0 9 1 11 11 2
9 10 9 13 1 11 2 1 11 2
8 3 15 13 10 9 1 11 2
9 15 13 10 9 0 1 10 11 2
17 15 13 10 0 9 1 10 9 2 10 11 2 1 11 11 11 2
13 15 13 10 9 1 9 1 9 1 10 9 12 2
7 1 10 9 13 3 9 2
7 3 15 13 10 11 11 2
7 1 10 9 4 13 11 2
8 15 13 10 3 0 9 0 2
9 15 13 10 0 9 1 11 11 2
13 3 15 13 10 9 15 13 10 9 0 1 11 2
9 15 13 10 0 9 1 11 11 2
7 10 9 4 13 11 11 2
8 3 13 1 10 11 11 11 2
8 3 15 13 10 9 1 11 2
7 1 10 9 9 10 11 2
12 10 9 4 13 1 10 9 0 1 10 9 2
9 15 13 0 10 9 1 11 11 2
10 10 9 0 13 10 10 9 1 11 2
16 1 10 9 1 11 4 13 10 9 2 10 9 13 15 2 2
6 3 4 13 11 11 2
8 15 13 10 11 1 10 11 2
12 15 13 2 15 3 4 13 1 13 2 2 2
13 3 15 13 10 0 9 13 1 11 1 9 0 2
8 15 13 10 0 9 1 11 2
15 10 9 1 10 9 13 1 13 1 10 9 1 10 9 2
18 10 9 0 13 10 9 1 10 11 1 11 11 1 10 11 7 11 2
9 10 9 15 13 1 10 9 11 2
11 1 10 11 2 15 13 10 9 1 11 2
7 1 10 9 15 13 11 2
7 10 9 15 13 1 11 2
5 3 13 11 11 2
8 15 13 10 9 1 10 11 2
8 3 15 13 10 9 1 11 2
8 3 13 10 11 1 10 11 2
8 3 15 13 10 9 3 13 2
8 1 10 9 4 13 10 9 2
11 1 10 9 4 3 13 11 11 11 11 2
6 3 13 11 11 0 2
11 15 13 10 9 0 1 10 9 1 9 2
7 1 10 9 13 11 11 2
9 15 1 10 9 1 9 4 13 2
9 3 15 13 10 11 1 10 11 2
9 10 9 15 13 1 10 11 11 2
9 15 13 10 9 0 1 10 11 2
10 3 15 13 10 0 9 1 9 13 2
8 1 10 9 4 13 10 9 2
7 10 9 13 10 11 11 2
16 15 13 10 9 1 10 9 2 10 9 9 1 11 11 2 2
12 15 13 10 0 9 1 10 9 0 1 9 2
6 1 3 13 10 9 2
8 10 9 0 13 0 1 11 2
10 15 13 10 9 1 10 11 7 11 2
8 3 1 10 3 13 0 11 2
12 15 13 10 0 9 1 10 9 1 11 11 2
7 1 10 9 15 13 11 2
9 10 9 13 11 11 1 10 12 2
11 1 10 9 15 13 10 11 11 1 11 2
5 15 13 11 11 2
15 15 1 10 0 7 0 9 1 11 13 10 9 1 11 2
8 15 13 0 10 9 1 9 2
12 10 15 13 10 9 1 9 2 9 9 2 2
6 3 13 10 9 11 2
8 1 10 15 4 13 10 9 2
17 15 13 10 9 1 10 9 15 13 10 9 1 10 10 9 0 2
9 1 10 9 15 13 10 9 11 2
19 10 9 1 9 4 13 10 9 2 0 1 11 2 1 10 11 11 11 2
14 10 9 13 10 9 1 10 11 7 11 11 1 11 2
8 13 10 9 1 9 1 13 2
8 1 10 9 4 13 11 11 2
7 10 15 13 11 5 11 2
5 3 13 11 11 2
5 15 13 0 11 2
10 3 4 13 10 9 2 11 11 2 2
5 3 13 11 11 2
8 15 13 0 10 9 1 9 2
14 10 9 13 3 3 7 13 10 11 11 1 10 11 2
7 3 4 9 10 0 9 2
11 11 11 13 1 9 10 9 1 10 9 2
10 3 4 13 10 11 1 10 11 11 2
5 3 13 11 11 2
5 3 13 11 11 2
20 10 9 13 10 9 1 10 9 1 10 12 2 10 11 1 10 9 11 2 2
8 1 10 9 0 13 11 11 2
7 3 4 13 10 11 11 2
10 3 4 4 13 10 11 11 11 11 2
6 15 13 11 10 11 2
14 1 10 15 4 13 10 9 0 2 11 11 11 2 2
15 1 10 9 13 10 9 3 0 1 10 9 1 10 11 2
7 10 9 13 10 11 11 2
10 10 9 15 13 1 10 11 11 11 2
8 10 9 15 13 1 13 9 2
12 10 11 4 13 1 9 1 10 0 11 11 2
9 3 15 13 10 9 1 11 11 2
8 11 11 3 13 10 10 9 2
5 3 13 11 11 2
10 1 10 9 1 10 9 11 15 13 2
7 10 9 13 11 11 11 2
11 10 9 13 10 9 1 13 10 10 9 2
9 15 13 10 9 1 10 9 0 2
10 15 4 13 10 9 0 1 11 11 2
14 1 10 9 4 13 10 9 1 2 11 1 11 2 2
14 1 1 10 9 1 10 9 10 9 0 13 1 13 2
7 10 9 15 13 1 11 2
9 10 9 13 10 11 1 10 9 2
6 15 13 11 10 11 2
10 15 13 10 9 3 0 1 9 0 2
6 10 9 13 10 9 2
9 1 10 9 4 13 15 10 9 2
9 1 10 9 2 10 9 13 9 2
11 10 9 1 9 15 13 1 10 11 11 2
11 10 9 13 10 9 1 9 0 11 11 2
14 10 9 4 13 1 10 2 9 1 10 11 11 2 2
6 13 10 9 9 0 2
5 15 13 11 11 2
6 10 9 13 10 11 2
13 10 9 15 4 13 1 10 9 1 10 11 11 2
12 10 9 13 10 11 1 10 12 1 10 12 2
11 1 10 9 1 10 9 15 13 10 9 2
7 10 15 13 10 9 11 2
8 15 13 10 9 0 0 0 2
14 1 10 9 15 13 1 10 9 10 11 1 10 9 2
8 15 13 11 1 10 11 11 2
15 10 9 1 10 9 1 9 13 3 1 10 9 1 9 2
12 15 13 10 9 1 11 1 2 11 11 2 2
9 15 13 10 9 1 10 11 11 2
12 15 13 0 10 11 1 10 11 1 9 0 2
6 15 13 0 10 11 2
5 10 9 4 11 2
13 15 13 0 2 1 9 2 10 11 1 10 11 2
8 15 13 0 10 11 11 11 2
14 10 9 13 10 11 11 1 10 0 9 1 10 12 2
10 1 10 9 15 13 10 11 11 11 2
8 10 15 13 10 11 1 11 2
10 13 10 9 1 9 13 1 11 11 2
16 1 10 9 2 10 9 1 11 13 10 9 1 9 1 9 2
8 3 13 10 10 9 10 11 2
6 15 13 0 10 11 2
7 10 9 0 13 10 11 2
16 15 13 10 0 9 1 10 11 1 13 10 0 9 1 9 2
18 10 9 13 10 9 1 13 10 9 1 9 1 10 9 1 10 11 2
9 1 10 9 15 13 10 11 11 2
13 10 9 1 10 11 11 13 11 11 1 10 11 2
8 10 9 13 11 11 16 13 2
16 15 1 10 10 9 13 11 1 13 10 9 3 1 10 11 2
11 10 9 9 13 2 10 0 0 9 2 2
9 15 13 10 9 1 10 9 0 2
13 1 15 13 10 9 1 10 9 0 1 10 9 2
8 15 13 10 9 0 3 0 2
5 15 13 11 11 2
10 10 9 13 10 9 1 10 9 0 2
7 10 15 13 10 9 0 2
13 1 10 9 4 13 11 1 10 10 9 1 11 2
6 3 13 11 1 11 2
5 3 13 11 11 2
9 10 9 15 13 1 10 9 0 2
6 13 10 9 1 9 2
12 1 10 9 15 13 10 11 1 11 11 11 2
16 10 9 1 10 11 11 13 0 1 10 10 0 9 1 9 2
12 10 9 1 10 9 0 4 13 1 10 11 2
10 10 9 15 13 1 10 9 1 11 2
19 10 9 1 10 11 11 11 13 10 9 1 10 9 2 1 10 9 13 2
7 1 10 9 13 10 11 2
11 15 13 10 3 13 9 0 1 10 9 2
9 1 10 9 0 13 10 9 0 2
13 1 10 9 15 13 10 3 0 9 1 10 9 2
5 15 13 11 11 2
15 10 9 0 4 4 13 2 10 0 9 1 10 9 2 2
7 3 15 13 10 0 11 2
9 3 4 4 13 1 9 11 11 2
10 15 13 10 9 3 0 1 10 9 2
7 10 9 0 13 10 11 2
8 3 13 2 9 2 1 9 2
19 15 13 10 9 1 10 0 9 15 13 9 1 10 9 7 1 10 9 2
13 10 9 0 13 9 1 10 0 9 1 10 12 2
6 10 9 0 0 13 2
7 13 10 9 7 9 9 2
6 10 9 13 10 9 2
7 10 9 15 13 1 11 2
8 3 13 10 10 9 10 11 2
6 10 9 13 11 11 2
6 10 9 13 11 11 2
9 3 15 13 10 0 1 10 9 2
6 10 15 13 10 11 2
5 15 13 11 11 2
9 10 9 11 1 11 13 10 9 2
13 1 10 9 1 11 15 15 13 1 2 11 2 2
9 3 4 13 10 9 1 11 11 2
15 10 9 1 10 11 11 13 10 9 13 2 11 11 2 2
7 3 13 11 1 10 11 2
5 3 4 13 11 2
11 10 9 13 1 9 1 12 9 3 0 2
6 10 15 13 10 9 2
17 10 9 4 13 3 9 1 9 1 9 1 10 15 1 10 9 2
11 1 10 9 1 10 11 15 13 11 11 2
21 10 9 13 10 11 1 10 0 0 9 16 15 13 16 13 10 10 9 1 9 2
12 10 9 13 11 11 1 0 1 10 9 0 2
18 10 9 4 13 1 0 9 0 2 0 1 10 9 7 9 1 9 2
20 1 10 9 10 9 1 10 11 11 11 11 2 11 11 2 13 10 10 9 2
7 10 9 4 13 11 11 2
7 3 13 10 10 9 11 2
5 15 13 11 11 2
13 10 9 0 13 10 9 1 10 9 11 1 11 2
6 10 9 13 10 9 2
14 10 9 0 4 13 2 2 10 9 13 10 9 2 2
9 1 10 9 15 13 10 11 11 2
7 3 15 13 10 9 9 2
8 1 10 9 15 13 10 9 2
8 15 13 10 2 11 11 2 2
15 10 0 13 0 1 10 0 9 1 9 0 1 10 9 2
10 3 4 13 10 0 9 1 11 11 2
13 15 13 10 9 1 10 9 1 10 9 0 0 2
7 10 9 15 13 1 11 2
5 3 13 11 11 2
10 1 10 9 13 10 9 1 10 9 2
8 15 13 0 10 9 3 0 2
11 1 10 9 1 10 11 4 13 11 11 2
7 3 0 4 13 10 9 2
9 3 15 13 2 15 2 1 0 2
12 10 9 1 9 13 9 1 10 11 11 11 2
11 15 13 10 9 3 0 1 10 13 0 2
5 15 13 11 11 2
12 10 9 1 9 4 4 13 1 13 10 9 2
10 10 2 8 8 2 4 13 11 11 2
6 3 13 11 1 11 2
9 3 4 13 10 9 1 10 9 2
10 10 9 0 13 10 0 9 1 9 2
9 10 9 15 13 1 10 11 11 2
10 1 10 9 0 13 9 11 1 11 2
12 10 9 1 11 11 4 13 1 10 12 11 2
8 15 13 10 0 9 1 11 2
7 3 4 4 13 10 9 2
6 1 10 9 13 11 2
5 3 4 13 11 2
6 10 15 13 10 9 2
10 13 10 9 1 9 0 1 9 0 2
18 10 9 4 13 1 12 9 10 9 2 9 9 2 1 10 9 0 2
9 1 10 9 0 13 9 11 11 2
7 15 13 11 3 1 13 2
8 1 10 9 13 11 11 11 2
10 10 9 0 0 15 13 1 11 11 2
11 10 9 0 13 9 1 10 9 1 11 2
6 3 4 13 10 9 2
9 10 9 13 10 0 9 1 9 2
8 15 13 10 9 0 1 11 2
8 15 13 10 9 0 1 11 2
7 10 9 13 9 1 9 2
10 3 4 13 10 9 1 10 11 11 2
9 15 13 10 0 9 1 11 11 2
10 10 9 10 11 4 13 10 11 11 2
6 15 13 11 11 11 2
9 10 9 0 13 1 10 10 9 2
27 13 10 9 1 9 15 4 13 1 10 9 7 1 10 10 9 9 1 9 15 4 4 13 1 10 9 2
7 15 13 0 10 9 11 2
7 1 10 9 13 11 11 2
8 10 9 7 9 13 11 11 2
8 3 13 10 9 1 11 11 2
14 1 10 15 13 10 9 2 11 2 2 9 0 2 2
16 10 9 13 1 10 9 12 7 12 10 9 2 11 11 2 2
10 3 15 13 10 9 0 1 10 9 2
5 3 13 11 11 2
17 1 10 9 11 11 13 1 10 0 9 1 10 9 0 1 9 2
5 15 13 11 11 2
11 1 10 9 15 13 11 11 2 1 11 2
8 1 10 9 11 15 13 0 2
11 1 10 9 13 10 9 1 10 11 0 2
5 15 13 11 11 2
8 15 13 10 9 1 11 11 2
11 15 13 10 9 1 9 2 9 0 2 2
5 3 13 11 11 2
13 15 13 10 0 9 1 11 11 1 10 11 11 2
7 3 13 0 10 9 11 2
5 10 9 13 11 2
13 10 9 0 1 10 9 4 13 2 10 11 2 2
14 13 10 9 0 1 10 9 15 1 9 13 10 9 2
10 1 10 9 4 13 11 11 11 11 2
11 10 9 13 10 11 11 1 10 11 11 2
13 3 4 13 1 10 9 1 10 0 9 10 11 2
5 3 13 11 11 2
15 10 9 1 11 11 4 4 13 1 10 9 1 10 11 2
6 10 15 13 10 9 2
5 15 13 11 11 2
9 10 9 0 13 10 9 13 11 2
8 10 15 13 10 11 1 9 2
9 10 9 1 9 0 13 11 11 2
6 10 15 13 11 11 2
11 10 9 4 13 1 10 9 1 11 11 2
8 3 4 13 10 11 11 0 2
9 3 15 13 10 9 1 10 9 2
10 1 10 9 4 9 10 9 0 11 2
9 10 9 13 10 9 1 11 11 2
14 10 9 13 10 0 9 1 9 1 10 9 1 11 2
15 10 0 9 1 10 0 9 15 13 2 11 1 9 2 2
9 15 13 10 9 0 1 10 9 2
12 15 13 10 9 1 10 9 0 0 1 9 2
13 15 13 0 10 9 1 10 9 1 9 9 0 2
15 10 9 1 9 4 13 2 4 13 9 7 15 4 13 2
8 3 13 10 9 1 11 11 2
13 15 13 10 9 1 10 9 1 10 9 1 11 2
8 3 13 10 9 1 11 11 2
10 1 10 9 4 13 15 1 10 11 2
9 10 9 13 10 0 9 1 9 2
13 10 15 15 13 10 11 1 10 11 1 9 0 2
7 3 0 4 13 10 9 2
11 15 13 10 0 9 0 1 10 0 9 2
9 15 13 10 9 1 2 11 2 2
5 15 13 11 11 2
11 10 9 4 13 1 10 11 1 10 12 2
10 3 4 13 10 2 11 2 1 11 2
5 15 13 11 11 2
7 15 13 0 10 11 11 2
10 10 0 9 13 11 11 1 10 12 2
11 10 9 1 13 15 13 1 10 9 11 2
7 1 10 9 13 10 11 2
15 1 10 9 0 15 4 13 9 0 13 1 9 1 9 2
8 10 0 1 11 13 10 11 2
10 3 1 9 4 13 10 9 0 0 2
11 3 15 13 10 0 9 1 10 9 0 2
7 15 13 2 11 11 2 2
7 1 10 9 13 10 11 2
9 1 10 9 15 13 10 11 11 2
5 3 13 11 11 2
13 1 10 9 1 10 9 1 10 9 15 13 11 2
11 1 10 15 4 13 10 9 1 10 9 2
7 3 15 13 1 11 11 2
10 1 10 9 15 13 10 9 1 11 2
16 3 15 13 10 9 0 0 1 9 13 1 10 11 1 11 2
11 3 15 13 10 11 11 1 10 11 11 2
14 1 10 9 0 13 9 11 11 3 1 10 11 11 2
6 15 13 0 10 9 2
5 10 15 13 11 2
11 10 2 9 2 13 11 11 1 12 11 2
6 10 15 13 10 9 2
7 10 9 1 11 15 13 2
9 10 9 0 13 10 9 11 14 2
5 15 13 11 11 2
14 1 10 9 15 13 10 9 0 13 13 1 10 9 2
8 10 9 15 13 1 10 9 2
14 10 9 4 13 1 10 9 10 9 1 10 0 9 2
7 10 9 9 4 13 11 2
9 3 15 13 10 0 1 10 9 2
14 10 0 9 3 1 10 11 13 1 9 0 10 0 2
5 3 13 11 11 2
7 1 10 9 13 10 11 2
8 10 9 13 10 9 11 11 2
6 15 13 0 11 11 2
11 10 9 4 13 1 10 9 1 12 9 2
20 10 9 0 0 2 0 7 0 2 4 4 13 1 9 1 9 1 9 0 2
8 10 15 13 11 1 10 11 2
9 3 4 4 13 10 0 9 0 2
5 15 13 11 11 2
12 1 10 0 9 15 13 10 0 9 1 11 2
11 3 4 4 13 10 9 1 10 11 11 2
9 10 9 4 13 2 11 13 2 2
10 1 10 9 4 13 10 9 1 11 2
7 10 15 13 10 11 11 2
13 10 9 4 13 10 3 0 9 0 1 10 9 2
17 3 4 13 10 9 15 2 1 10 10 9 4 13 2 3 13 2
19 10 9 1 10 9 11 11 15 13 4 13 1 10 9 1 10 11 11 2
16 1 10 11 2 3 13 10 9 1 10 12 9 1 10 9 2
5 15 13 11 11 2
10 15 13 10 9 3 0 1 10 11 2
8 1 10 9 13 10 11 11 2
12 10 9 13 10 9 3 13 1 10 10 9 2
6 15 13 0 10 11 2
8 1 10 9 4 13 11 11 2
17 10 15 13 10 9 1 10 9 0 0 1 10 9 1 10 9 2
13 15 13 0 10 9 0 1 10 9 1 11 11 2
16 1 10 9 10 9 0 15 13 1 9 1 10 9 15 13 2
18 13 10 9 1 10 11 15 4 4 13 7 13 1 10 9 0 0 2
6 10 9 13 11 11 2
14 1 10 9 15 13 3 10 9 1 10 9 1 11 2
12 1 10 9 11 11 13 10 11 1 0 9 2
12 10 9 0 1 9 4 13 12 9 1 9 2
10 10 9 15 13 1 10 10 11 11 2
7 10 9 13 3 10 0 2
7 15 13 0 10 11 11 2
5 10 9 4 13 2
22 1 10 9 1 10 11 7 1 10 9 1 11 11 2 11 2 15 13 9 1 11 2
9 15 13 10 9 1 10 9 0 2
10 3 15 13 2 15 13 2 1 9 2
10 10 9 4 13 9 0 1 10 9 2
10 15 13 10 9 3 0 1 10 9 2
7 10 15 13 10 11 11 2
8 3 4 4 13 10 9 0 2
9 1 10 9 11 13 10 10 9 2
21 15 13 0 10 2 11 11 2 15 15 13 1 10 9 11 2 11 1 10 12 2
7 10 9 13 11 16 13 2
6 3 13 11 11 11 2
14 10 9 4 13 1 11 11 7 11 11 1 10 12 2
5 15 13 11 11 2
11 1 9 10 9 1 10 9 10 9 13 2
9 15 13 10 9 1 10 9 11 2
8 15 13 10 9 1 10 11 2
9 1 10 9 1 9 13 10 11 2
9 10 9 1 9 13 10 11 11 2
13 10 9 13 10 0 9 1 0 1 10 10 9 2
5 15 13 11 11 2
7 15 13 0 10 9 11 2
6 3 4 13 11 11 2
7 1 10 9 15 13 11 2
11 15 13 10 9 1 4 13 1 10 9 2
5 3 13 11 11 2
13 10 9 0 13 16 10 11 13 1 10 11 11 2
13 10 9 15 13 1 10 11 11 7 10 11 11 2
9 15 13 10 9 0 13 1 11 2
11 10 9 0 13 1 10 12 1 10 12 2
6 15 13 10 11 11 2
9 1 10 15 4 13 10 9 0 2
9 10 15 13 11 1 10 11 11 2
8 1 10 9 15 13 10 11 2
6 3 4 13 10 9 2
16 13 10 9 1 9 13 1 10 10 9 1 11 7 11 11 2
9 3 4 13 10 9 1 10 9 2
10 10 9 1 10 9 13 10 9 0 2
19 10 9 1 10 11 11 0 1 10 12 13 1 10 9 10 9 1 9 2
13 10 9 0 4 13 1 0 9 0 1 10 12 2
9 15 13 10 0 9 1 11 11 2
17 1 10 9 1 10 9 0 13 13 1 13 10 9 1 10 9 2
6 3 13 10 0 11 2
10 15 13 10 9 3 0 1 10 9 2
11 3 13 10 9 1 10 9 1 10 11 2
7 15 13 0 10 11 11 2
9 1 10 9 13 9 11 11 11 2
8 10 9 13 10 9 0 0 2
8 3 9 15 13 1 10 9 2
13 10 9 0 15 4 13 1 10 9 1 10 11 2
11 1 10 9 10 11 11 13 10 10 9 2
17 10 9 13 9 7 9 1 10 9 1 9 1 10 11 1 11 2
7 10 9 13 3 10 9 2
10 15 13 10 9 3 0 1 10 11 2
6 10 9 13 11 11 2
6 10 9 13 10 9 2
7 3 4 13 10 0 11 2
8 10 9 15 13 1 11 11 2
13 10 9 1 10 0 0 13 1 10 9 1 9 2
7 3 13 9 10 0 11 2
11 15 13 0 10 9 1 9 1 10 9 2
5 15 13 11 11 2
7 1 10 9 13 11 11 2
9 10 9 15 13 1 10 9 0 2
12 10 9 13 1 10 9 11 11 1 11 11 2
10 10 9 4 13 3 9 1 10 11 2
12 10 9 4 13 1 4 13 1 10 9 0 2
9 10 9 13 11 11 1 12 9 2
5 3 13 11 11 2
6 10 9 1 9 13 2
5 3 13 11 11 2
6 3 13 11 11 11 2
9 10 9 13 10 9 9 11 11 2
8 3 4 4 13 10 9 13 2
13 3 10 11 11 4 13 1 9 1 10 0 9 2
9 10 9 4 13 11 1 10 12 2
10 10 9 13 10 11 0 1 10 12 2
18 15 13 10 9 1 10 9 1 10 9 0 1 10 9 1 11 11 2
13 10 9 4 13 10 11 1 10 11 1 9 0 2
9 10 15 13 10 9 1 0 11 2
5 15 13 11 11 2
7 15 13 0 10 9 0 2
11 1 10 9 10 9 4 13 1 10 9 2
10 10 9 13 10 9 1 11 11 11 2
5 3 13 11 11 2
15 10 9 0 1 10 0 9 13 1 11 11 2 1 11 2
6 10 9 13 11 11 2
13 10 3 0 9 0 1 10 9 4 13 11 11 2
13 15 13 9 1 10 9 1 11 1 2 11 2 2
13 10 9 1 10 9 15 13 1 10 9 1 11 2
9 15 13 10 9 1 10 0 9 2
13 1 10 9 15 13 10 0 9 11 13 1 9 2
7 15 13 0 10 11 11 2
17 15 4 4 13 3 12 9 1 10 11 11 7 3 4 3 13 2
10 3 0 13 1 10 11 1 10 9 2
8 1 10 9 13 10 9 11 2
6 10 15 13 10 11 2
7 15 13 0 10 11 11 2
5 15 13 11 11 2
9 3 4 4 13 10 0 9 0 2
10 10 9 1 9 13 9 1 10 9 2
7 15 13 10 11 14 11 2
10 15 13 10 9 3 0 1 10 9 2
6 10 9 13 11 11 2
15 1 10 9 13 10 9 1 10 9 3 0 1 10 9 2
9 10 9 13 10 0 9 1 9 2
5 3 13 11 11 2
10 15 13 10 9 0 1 10 9 0 2
13 3 15 13 10 9 0 1 10 9 1 10 11 2
11 15 13 10 9 1 9 1 11 1 11 2
9 1 10 9 15 13 10 11 11 2
5 3 13 11 11 2
8 1 15 13 10 9 1 11 2
6 10 15 13 10 11 2
5 3 13 11 11 2
11 1 10 9 15 13 10 9 1 11 11 2
14 10 9 0 1 11 11 13 10 10 9 1 11 11 2
7 10 9 15 13 1 11 2
21 3 0 9 1 10 11 4 13 1 9 0 9 1 9 0 1 12 1 12 9 2
7 10 9 13 10 9 0 2
14 1 10 9 13 10 9 1 11 11 3 1 13 9 2
3 15 13 2
6 15 15 4 13 3 2
7 15 4 13 1 10 9 2
8 15 13 1 10 9 1 15 2
9 15 4 13 1 10 9 1 11 2
6 15 13 1 10 9 2
5 15 4 13 11 2
6 1 15 15 4 13 2
12 15 13 10 9 0 1 10 9 2 11 2 2
12 1 15 4 13 10 11 1 9 1 10 12 2
9 15 13 10 9 0 1 10 11 2
11 15 4 13 10 9 1 11 1 10 12 2
7 1 15 13 9 10 11 2
7 1 15 4 13 10 9 2
3 15 13 2
5 15 13 10 11 2
7 15 4 13 1 10 11 2
8 10 15 4 13 1 10 11 2
6 15 13 1 10 9 2
7 10 15 13 1 10 9 2
8 10 15 4 13 10 9 11 2
8 15 4 13 10 11 11 11 2
5 15 13 10 11 2
5 15 13 10 11 2
6 11 4 13 10 9 2
7 10 15 4 13 10 9 2
6 15 4 13 10 9 2
6 15 4 13 10 9 2
7 10 15 4 13 10 9 2
8 15 4 13 10 9 1 13 2
7 15 4 13 1 10 9 2
6 15 4 13 10 11 2
6 15 4 13 10 9 2
6 15 4 13 10 9 2
6 15 4 13 10 9 2
11 1 10 15 4 13 10 9 1 10 9 2
6 1 15 13 10 9 2
3 15 13 2
3 15 13 2
5 15 4 13 11 2
5 15 13 1 11 2
8 15 13 10 9 15 13 11 2
9 15 13 10 9 0 9 1 9 2
3 15 13 2
5 1 15 13 3 2
9 1 15 13 10 9 1 10 11 2
7 15 13 0 10 11 11 2
5 1 15 13 11 2
3 15 13 2
3 15 13 2
3 15 13 2
8 15 13 1 15 15 4 13 2
5 15 9 13 11 2
8 1 10 9 13 11 1 11 2
8 1 10 9 4 13 11 11 2
7 1 10 9 13 9 11 2
6 10 9 13 3 0 2
5 10 0 4 13 2
6 10 9 4 4 13 2
5 10 9 4 13 2
5 10 9 15 13 2
5 10 9 4 13 2
5 10 9 4 13 2
6 10 9 13 15 3 2
9 10 9 15 13 1 10 10 9 2
6 10 9 13 1 13 2
10 10 9 13 3 0 1 10 11 11 2
15 1 10 9 15 13 10 9 1 10 11 11 1 10 11 2
11 10 9 0 13 1 10 9 1 12 9 2
6 10 9 13 10 9 2
6 10 9 13 10 9 2
8 10 9 4 13 10 9 0 2
8 10 9 4 13 1 10 9 2
8 10 9 4 13 1 10 9 2
6 10 9 13 1 15 2
6 10 9 13 1 9 2
6 10 9 13 1 9 2
6 10 9 13 1 13 2
5 10 9 13 11 2
6 10 9 13 10 11 2
7 10 9 4 13 1 13 2
3 3 13 2
10 3 15 13 10 9 9 1 10 11 2
6 3 4 13 10 9 2
7 3 15 13 1 10 9 2
11 3 15 13 10 9 1 10 9 0 0 2
6 3 13 10 11 0 2
11 3 4 13 10 9 9 1 4 4 13 2
6 3 15 13 10 9 2
10 3 15 13 10 9 0 1 10 12 2
6 3 4 13 10 9 2
7 3 15 13 10 9 0 2
3 3 13 2
6 3 4 13 10 9 2
5 3 15 4 13 2
5 3 10 9 13 2
6 3 3 4 3 13 2
6 3 11 3 4 13 2
7 3 3 15 15 4 13 2
6 3 11 13 10 9 2
11 3 10 11 4 13 1 9 10 0 9 2
18 1 10 9 1 9 2 3 2 10 0 9 0 15 13 1 10 11 2
13 9 11 11 2 13 10 9 1 9 1 11 11 2
8 11 4 13 1 9 1 9 2
50 1 12 9 0 1 9 1 11 2 9 1 10 9 0 1 10 11 2 15 4 13 10 9 1 9 1 11 11 2 0 9 1 10 9 0 1 11 7 15 1 10 2 9 0 2 1 10 9 0 2
41 10 9 0 4 13 10 9 0 1 11 2 13 16 10 10 2 0 2 9 1 10 9 1 9 7 9 1 9 2 3 13 9 1 10 9 13 1 10 9 2 2
41 10 9 0 1 11 4 4 13 10 0 9 1 10 9 1 15 10 9 2 11 11 2 4 4 13 1 4 13 10 9 1 9 0 7 9 1 9 2 11 11 2
58 11 11 2 9 1 10 0 9 11 2 13 3 1 10 9 7 1 10 9 11 7 1 10 9 11 1 10 9 1 10 9 11 2 4 13 10 9 1 12 9 7 12 9 1 9 1 10 9 1 9 1 9 13 7 9 1 9 2
20 10 9 0 11 4 13 9 1 10 9 1 10 11 1 10 9 1 10 11 2
36 10 9 2 1 10 15 3 15 4 13 1 10 9 1 10 9 1 10 9 2 11 11 7 11 11 13 15 9 1 10 9 11 1 10 11 2
18 10 9 11 11 7 11 11 13 15 9 1 10 9 11 1 10 11 2
25 11 11 11 2 10 9 13 1 9 0 2 4 13 1 4 13 3 10 9 1 9 1 10 9 2
43 1 10 0 9 11 11 2 10 11 1 11 2 15 4 13 10 9 1 10 12 2 13 10 9 3 1 11 11 2 10 9 1 10 9 1 10 15 10 9 15 4 13 2
19 1 10 9 10 9 11 11 7 10 0 9 2 0 9 11 2 11 11 2
30 10 12 9 12 10 9 11 11 13 10 9 1 10 15 13 0 12 9 1 15 11 11 1 10 9 1 9 1 9 2
35 1 10 9 1 10 12 13 10 9 1 10 9 1 11 11 7 0 9 1 10 9 1 4 13 1 13 10 9 1 10 9 0 1 11 2
40 1 10 9 1 10 9 1 10 9 1 10 9 11 11 11 2 13 1 10 11 2 15 13 16 10 9 11 11 4 13 7 13 10 9 1 10 10 0 9 2
39 10 12 9 0 10 9 4 13 10 9 13 1 10 9 0 11 11 7 11 11 11 15 13 3 1 10 9 1 10 9 1 10 9 1 10 9 1 11 2
32 1 10 9 1 10 11 11 11 1 10 9 11 11 11 2 15 9 12 9 13 9 1 10 9 1 9 0 1 10 11 11 2
7 11 11 13 9 11 11 2
13 10 9 11 11 4 13 10 9 11 1 9 0 2
17 10 9 1 10 11 11 11 2 11 11 2 3 13 1 10 9 2
25 10 9 1 11 2 11 11 2 13 1 10 9 1 10 0 9 2 3 13 1 11 1 11 11 2
12 1 10 9 10 9 1 11 11 2 11 11 2
15 11 11 7 10 10 11 11 11 13 10 0 9 1 11 2
14 11 11 2 9 0 2 0 1 11 7 0 1 11 2
11 10 9 4 13 11 7 4 4 13 11 2
27 10 9 0 1 11 11 11 2 1 10 11 1 10 11 2 4 13 1 9 1 9 3 1 10 12 9 2
11 10 9 3 13 1 13 1 9 11 11 2
21 11 2 9 1 11 7 9 1 11 11 2 4 3 13 1 10 9 1 10 9 2
13 1 10 9 1 10 9 4 13 10 12 9 0 2
18 13 1 10 9 1 10 9 2 11 13 1 13 0 1 13 10 9 2
18 7 16 10 11 13 1 0 11 2 10 9 4 13 10 9 1 11 2
16 10 9 4 4 13 3 1 10 9 1 13 10 9 11 11 2
26 10 9 1 10 11 11 11 4 13 1 11 10 9 1 10 9 1 10 9 1 10 9 1 10 11 2
20 7 10 9 1 10 9 13 3 0 1 13 0 9 1 10 11 1 10 11 2
16 10 11 4 13 3 1 13 10 9 1 10 9 1 10 11 2
27 13 11 11 10 9 1 10 9 1 10 9 0 15 4 13 1 13 11 11 9 1 10 11 1 10 12 2
27 10 12 4 13 1 13 10 9 1 10 9 1 10 9 1 10 0 9 1 10 9 13 3 1 10 9 2
12 4 3 13 10 9 7 13 10 9 1 13 2
26 10 9 4 13 9 9 7 3 10 9 2 0 1 10 9 1 9 13 1 10 9 2 15 4 13 2
21 10 9 4 4 13 1 9 0 1 10 12 9 1 9 0 2 3 1 10 9 2
25 10 9 0 2 15 13 1 10 12 2 13 10 9 1 10 12 9 0 1 10 9 1 10 9 2
21 3 2 10 9 1 10 9 4 13 10 9 2 13 15 3 1 10 9 1 11 2
17 9 13 3 10 11 11 2 15 13 9 1 10 11 11 7 11 2
23 10 9 0 4 13 1 4 13 1 10 9 0 2 9 15 13 1 13 10 9 1 9 2
20 3 3 10 11 11 4 13 1 13 15 9 0 2 13 10 9 1 12 9 2
25 10 9 11 11 15 4 13 1 13 16 13 10 9 1 9 0 7 4 13 15 1 10 12 9 2
20 1 10 9 4 4 13 10 10 9 1 9 2 13 10 9 0 1 11 11 2
23 13 16 13 1 9 2 13 0 16 15 13 3 10 9 11 2 13 10 9 11 11 11 2
26 10 9 4 13 1 10 11 1 11 1 9 0 1 10 9 1 9 1 10 9 1 9 1 10 9 2
16 1 10 0 9 1 10 9 10 9 13 10 9 1 9 0 2
23 9 1 11 1 10 9 1 10 11 11 1 10 9 1 10 9 11 11 7 10 9 11 2
34 1 9 1 10 9 0 11 11 7 11 11 11 4 4 13 10 9 1 9 1 9 1 11 11 2 0 9 0 1 10 9 1 11 2
28 13 3 11 11 2 10 0 9 13 13 1 10 9 1 10 9 1 10 9 1 11 1 10 9 11 1 11 2
8 4 13 3 10 10 9 11 2
38 3 4 13 10 9 3 1 9 1 11 11 2 10 0 9 1 11 11 2 1 10 9 0 1 11 11 2 1 10 9 1 9 0 1 10 9 11 2
73 10 9 13 1 10 11 1 11 7 1 10 9 1 10 11 1 11 2 4 13 1 10 9 1 9 1 10 9 0 1 11 2 11 11 2 2 4 13 10 9 13 1 12 9 1 10 9 11 11 11 2 11 7 11 2 1 10 9 1 11 1 10 9 1 10 9 13 1 10 9 0 2 2
31 13 9 1 15 10 9 11 2 1 10 9 1 15 1 10 9 1 11 2 11 11 2 13 1 9 1 9 2 1 9 2
22 1 10 9 1 10 12 9 2 1 11 7 11 2 15 13 1 10 15 1 10 9 2
24 1 15 13 11 2 9 1 10 9 0 2 4 13 9 1 15 7 10 9 13 1 9 0 2
18 3 10 9 1 11 11 2 11 11 2 3 13 10 9 1 10 9 2
27 3 1 9 1 10 9 15 13 10 11 11 1 11 11 2 9 0 1 10 9 0 1 9 1 11 11 2
13 11 13 10 0 9 1 10 9 1 11 7 11 2
25 4 13 1 10 12 1 10 9 1 9 3 13 3 10 9 1 10 11 1 10 11 11 11 11 2
23 10 9 1 11 2 3 1 15 1 11 2 13 1 10 9 1 10 11 11 11 1 11 2
67 13 1 10 9 1 10 9 1 10 9 1 10 11 11 15 4 13 3 10 9 1 11 11 2 13 1 10 9 10 0 9 1 10 9 2 7 11 11 2 9 1 11 11 2 9 1 9 1 10 9 1 11 1 11 2 1 10 9 9 0 1 10 9 11 11 11 2
67 10 9 11 5 11 2 1 15 11 11 13 9 2 1 10 9 1 10 9 1 10 9 4 13 1 10 9 1 10 11 1 11 11 2 9 1 11 2 3 15 1 10 9 1 10 9 1 10 9 1 10 0 9 1 10 9 0 1 10 11 11 11 11 2 5 2 2
59 1 10 9 1 10 11 11 1 10 12 4 3 13 10 9 1 10 11 5 11 7 10 9 1 10 11 11 2 10 15 13 1 10 9 11 7 11 11 1 13 15 1 9 1 10 9 0 15 13 1 13 1 10 12 5 1 10 9 2
20 2 1 10 9 13 15 12 9 1 10 11 2 3 10 9 3 13 15 2 2
22 7 10 11 2 1 10 0 9 1 11 2 11 2 9 12 2 13 3 10 9 11 2
19 3 9 10 9 1 9 1 10 11 13 1 9 10 9 13 11 11 11 2
57 1 13 10 10 9 13 1 9 2 1 10 9 1 10 0 9 2 12 9 1 9 2 10 0 9 12 1 11 11 11 11 7 10 0 9 1 9 0 1 10 9 11 11 7 10 9 0 11 11 2 9 1 10 0 9 11 2
23 7 10 0 9 1 9 13 10 9 1 10 9 0 11 11 2 1 9 1 9 1 11 2
33 3 1 10 11 4 13 10 0 9 1 10 9 0 1 11 2 11 11 2 13 1 10 9 9 1 10 9 1 4 13 10 9 2
31 3 13 1 9 1 11 16 10 9 1 10 9 11 11 11 4 4 13 1 10 9 11 11 16 15 13 11 1 10 9 2
36 11 4 3 13 0 16 4 4 13 3 10 9 1 10 9 11 11 7 16 4 4 13 9 1 10 9 1 10 11 1 10 11 2 11 11 2
18 1 9 10 11 11 4 13 1 9 10 9 1 10 9 1 10 11 2
7 11 4 13 16 13 11 2
21 10 11 4 13 10 0 9 1 11 2 1 10 9 0 1 11 1 10 0 9 2
28 16 11 13 2 1 10 9 9 0 4 13 1 0 9 11 11 2 0 9 0 11 11 2 3 1 10 9 2
30 1 9 4 13 15 10 9 11 11 2 13 1 9 2 3 9 0 1 10 11 11 11 2 10 9 9 1 10 9 2
29 7 3 11 2 10 9 1 10 9 0 15 4 13 3 1 10 9 1 4 13 12 9 1 9 0 1 10 11 2
73 10 9 11 13 1 10 10 9 3 1 10 9 2 3 1 16 10 9 4 4 13 1 10 9 1 10 9 1 10 9 13 1 11 11 2 11 11 2 1 10 9 1 10 9 1 10 0 9 13 1 11 1 11 11 2 15 13 13 2 1 9 0 2 11 11 2 9 0 1 9 11 11 2
31 10 9 4 13 2 13 11 1 10 9 1 10 9 1 10 9 0 7 1 9 0 2 13 7 9 7 9 0 2 2 2
29 16 11 13 1 10 11 10 9 1 11 11 2 10 9 1 10 9 0 11 11 13 10 9 0 15 13 10 9 2
36 16 11 13 10 9 1 10 11 1 13 10 0 9 1 11 11 2 10 0 9 1 9 11 13 10 9 1 13 10 9 1 10 9 1 11 2
23 10 9 13 1 11 2 1 10 9 1 10 9 9 11 11 11 2 7 1 10 0 11 2
21 12 9 2 0 9 11 2 11 4 13 1 10 0 9 1 13 9 1 10 9 2
13 12 7 12 4 13 9 1 10 9 0 7 0 2
26 10 9 13 13 10 9 1 11 11 2 15 13 3 1 10 9 1 9 1 11 1 9 1 10 9 2
29 11 13 3 3 9 1 10 9 1 9 1 11 11 7 13 1 10 9 10 9 0 15 15 13 9 13 1 11 2
16 10 9 1 11 11 1 10 9 1 10 9 1 9 1 11 2
28 7 10 9 7 9 0 1 10 11 11 11 3 13 9 7 2 11 2 11 2 3 9 13 9 1 11 2 2
24 10 9 13 1 10 9 0 1 10 9 2 11 11 2 11 2 13 10 12 9 1 10 12 2
58 1 10 9 1 10 9 13 1 10 11 1 10 11 0 10 9 13 1 9 1 10 9 0 1 10 11 11 1 11 2 9 1 9 2 15 13 1 10 9 1 10 9 11 1 10 11 11 11 1 11 1 10 9 1 9 12 2 2
46 11 11 11 4 13 1 11 11 2 0 9 1 10 9 13 1 9 0 1 10 9 1 10 9 1 10 9 0 1 10 11 1 11 7 1 10 9 1 11 1 10 9 11 1 11 2
16 11 3 13 13 1 10 9 1 10 9 1 10 11 11 11 2
48 10 9 0 4 13 1 13 1 10 12 7 10 12 2 3 16 10 11 1 10 11 2 7 1 9 11 2 4 13 1 15 1 9 0 1 10 9 1 11 10 0 9 1 12 9 1 9 2
46 3 2 10 11 11 11 4 13 10 9 0 1 10 9 1 10 11 11 11 1 11 11 2 15 1 10 9 4 13 1 10 11 11 11 2 13 3 3 7 0 3 1 10 0 11 2
14 10 0 9 1 10 15 3 13 10 9 1 10 11 2
19 11 13 0 1 10 9 0 0 11 11 1 10 15 4 13 1 10 9 2
18 10 9 1 10 9 2 1 10 15 3 13 10 9 2 4 4 13 2
10 10 9 1 10 15 13 10 11 0 2
11 10 9 1 9 1 10 15 13 10 9 2
12 13 10 9 0 2 1 10 15 3 15 13 2
16 10 9 0 1 10 15 13 10 9 2 15 4 13 10 9 2
58 10 9 0 1 10 15 10 9 1 10 11 11 2 11 11 2 4 13 0 1 10 9 1 9 1 10 9 13 1 10 9 1 9 0 1 9 1 10 11 0 1 10 15 4 13 2 1 10 9 1 9 2 10 0 9 11 11 2
17 10 9 1 10 9 0 11 11 13 10 9 0 15 13 10 9 2
8 10 9 15 15 13 13 9 2
22 1 9 1 11 11 11 11 3 11 11 2 15 13 10 9 1 9 1 10 9 0 2
7 11 4 13 16 13 11 2
17 10 9 13 16 11 2 13 2 13 10 10 9 1 10 9 0 2
18 11 4 3 13 0 16 4 4 13 3 10 9 1 10 9 11 11 2
12 11 4 13 16 11 3 4 3 13 10 11 2
19 1 10 9 15 13 16 1 10 9 1 10 9 1 10 11 15 13 9 2
34 10 9 11 5 11 2 1 15 11 11 13 9 2 1 10 9 1 10 9 1 10 9 4 13 1 10 9 1 10 11 1 11 11 2
21 10 9 1 10 9 13 10 9 13 1 15 10 9 11 13 13 10 9 1 11 2
11 1 10 0 9 1 15 13 0 13 9 2
37 10 9 1 10 9 0 11 13 10 9 1 10 9 1 12 9 1 10 9 0 1 9 1 11 2 13 1 11 2 1 15 13 3 9 0 11 2
14 12 9 1 15 12 4 13 1 9 1 10 9 11 2
15 11 2 13 1 11 2 7 1 15 13 3 9 0 11 2
22 10 9 2 15 1 10 9 7 1 10 9 1 15 4 13 10 9 1 9 7 9 2
17 9 0 1 9 2 9 1 9 2 9 1 15 15 13 1 9 2
20 13 12 9 2 1 15 10 0 9 11 11 7 10 9 0 1 11 11 11 2
24 1 10 9 1 10 12 4 13 1 12 9 1 9 1 9 11 11 2 9 0 0 1 11 2
18 10 9 15 13 3 1 10 9 1 9 10 1 11 2 1 10 9 2
17 16 11 11 15 4 13 7 15 4 13 2 11 11 4 1 0 2
18 13 10 9 1 11 11 2 3 13 1 10 9 15 15 13 1 9 2
5 11 11 1 9 2
23 10 12 9 9 1 10 9 1 11 12 4 13 1 9 1 10 9 1 11 2 11 2 2
14 1 10 9 2 15 13 9 0 2 10 9 13 3 2
17 10 9 2 15 13 10 9 15 15 4 13 1 12 2 13 3 2
40 4 13 1 10 9 0 1 10 12 7 10 12 9 0 11 11 2 10 12 9 9 1 10 9 1 11 12 2 13 1 9 1 10 9 1 11 2 11 2 2
23 2 3 4 13 15 1 10 9 1 11 11 2 4 13 3 10 9 13 1 13 10 9 2
17 15 13 1 2 9 0 0 2 7 0 2 9 0 7 0 2 2
18 10 0 9 0 4 4 2 13 10 0 9 7 10 9 4 13 3 2
9 4 4 13 1 9 1 9 2 2
14 10 9 2 2 1 9 3 4 13 0 1 9 2 2
34 10 9 2 13 1 10 9 1 10 9 2 13 16 15 13 1 10 2 9 0 7 16 10 9 13 0 1 10 9 1 10 9 0 2
24 10 10 9 4 4 13 1 9 2 13 2 7 3 4 13 15 1 10 9 1 11 11 2 2
29 15 2 1 10 9 2 13 1 9 0 0 7 9 2 2 9 15 13 1 10 0 9 0 7 13 10 9 0 2
12 13 9 1 9 7 3 4 13 1 9 0 2
14 10 9 0 7 3 15 4 13 1 10 9 1 9 2
16 1 9 3 4 13 0 1 9 2 13 10 9 1 10 9 2
22 3 4 13 10 9 2 10 9 11 4 13 1 10 0 9 15 3 3 4 4 13 2
14 4 13 7 3 13 1 10 9 2 13 10 9 0 2
32 10 10 9 13 9 7 9 2 7 13 3 3 3 1 13 10 9 2 2 4 13 10 9 1 10 9 1 11 2 11 11 2
18 10 11 1 11 4 13 10 9 1 10 9 7 10 9 1 10 9 2
48 1 10 9 11 11 4 13 2 3 2 16 10 9 15 4 13 1 10 9 3 2 3 1 10 9 0 1 11 2 7 16 2 3 4 13 15 10 9 2 10 9 7 10 9 1 9 2 2
29 10 9 15 4 13 3 1 10 12 2 1 10 9 1 9 3 10 9 13 0 1 9 7 3 1 10 9 2 2
25 1 10 9 11 2 4 13 3 10 9 1 15 1 10 9 16 4 13 13 1 10 0 9 2 2
13 10 9 1 10 9 13 10 9 1 15 1 11 2
38 11 11 2 10 9 9 15 4 13 10 9 1 10 9 1 10 9 1 11 1 10 12 2 13 0 16 10 0 9 0 4 13 1 9 1 10 9 0
33 10 9 4 13 1 4 13 1 10 9 0 1 9 2 7 15 4 13 1 10 9 0 1 10 9 1 10 0 9 13 1 3 2
36 10 9 0 4 13 1 13 10 9 1 10 9 1 10 9 7 4 13 10 10 9 0 1 10 12 7 12 9 2 1 9 1 10 9 13 2
17 11 15 13 11 2 13 10 9 1 10 11 2 11 11 1 11 2
24 10 9 13 10 9 1 10 9 13 1 11 2 15 15 13 3 3 1 10 0 9 1 9 2
15 3 1 10 12 4 13 10 9 9 1 10 9 1 11 2
13 10 9 13 10 9 1 10 9 1 10 0 9 2
14 1 11 3 10 9 1 10 9 1 10 11 11 11 2
26 2 10 10 9 13 1 11 11 1 10 9 0 2 11 3 1 15 15 13 10 9 1 13 15 2 2
45 2 11 1 15 4 13 1 10 9 2 4 13 2 7 13 2 1 10 10 9 1 10 9 1 10 10 9 1 11 12 2 13 11 11 2 9 1 10 11 1 9 1 11 12 2
19 11 4 13 3 10 9 1 9 15 15 13 1 10 0 9 1 10 11 2
18 13 1 13 3 3 10 9 0 2 13 11 11 2 9 1 10 11 2
24 10 9 1 10 9 1 11 11 1 11 11 3 1 11 11 11 13 10 10 9 1 10 9 2
13 9 1 10 9 1 10 9 3 1 10 9 0 2
46 2 1 9 1 9 2 10 11 7 10 9 1 10 9 4 13 0 16 4 13 1 10 0 9 1 10 9 1 11 11 2 4 13 13 10 9 1 11 11 2 11 11 2 1 11 2
31 2 4 13 0 1 10 13 16 13 1 9 0 7 13 1 9 10 0 9 0 1 11 2 13 13 10 11 1 10 9 2
26 2 13 15 3 13 0 10 9 0 1 11 7 15 13 10 10 10 9 7 10 9 1 10 0 9 2
14 13 3 16 13 3 7 16 13 3 3 1 15 2 2
6 11 11 2 11 11 2
9 2 11 13 9 2 9 7 9 2
12 10 12 1 11 11 13 10 9 1 10 9 2
21 1 9 10 0 9 0 1 11 15 13 1 11 11 3 1 10 9 1 11 11 2
20 10 0 9 16 11 13 10 9 7 15 13 1 3 1 10 9 7 10 9 2
31 10 0 11 11 1 11 11 4 3 13 1 10 9 0 1 10 9 13 1 10 9 1 15 13 9 1 10 12 9 0 2
15 2 11 2 4 13 11 2 13 10 9 1 10 9 0 2
9 10 10 9 0 7 0 13 0 2
39 3 2 3 1 11 15 13 10 9 13 1 9 0 7 0 2 9 0 2 0 2 0 2 15 13 10 9 3 3 1 10 0 9 2 7 1 10 9 2
28 1 11 3 13 3 0 10 9 1 10 9 0 7 0 1 9 0 2 7 10 9 0 1 15 13 3 9 2
20 11 13 10 9 0 1 9 2 2 4 13 10 11 2 7 3 0 1 9 2
27 7 15 13 10 9 1 4 13 1 10 0 9 1 9 7 1 9 2 16 15 13 9 1 9 0 2 2
22 1 10 10 9 1 10 9 1 10 12 11 11 4 4 13 3 10 9 1 9 0 2
11 2 3 13 10 9 1 10 9 1 11 2
5 13 1 10 15 2
11 3 13 10 9 1 10 10 2 9 2 2
21 10 9 4 13 2 1 10 10 2 0 2 2 1 13 15 0 2 0 2 0 2
22 1 9 2 10 9 1 10 9 13 1 10 9 10 10 9 13 10 15 15 15 13 2
14 1 3 10 9 1 10 11 15 4 13 1 10 9 2
21 2 10 9 13 2 3 13 1 10 0 9 2 1 13 10 3 0 10 10 9 2
52 10 11 1 10 9 0 13 10 9 3 3 0 16 13 3 3 0 1 9 2 0 2 0 2 16 10 15 4 0 7 0 1 15 13 1 9 2 16 13 13 1 9 0 7 0 2 1 10 9 1 15 2
66 10 11 1 10 9 0 13 0 16 3 15 13 9 15 15 13 2 1 0 2 2 15 13 10 10 9 3 2 1 10 9 2 2 1 13 15 1 10 9 0 2 9 1 9 7 9 15 2 1 10 9 7 1 10 9 2 15 13 7 3 2 13 10 9 2 2
12 10 12 1 11 11 13 10 9 1 10 9 2
24 1 10 9 0 1 10 0 9 1 10 11 0 3 1 10 9 1 10 9 1 10 11 11 2
26 9 0 1 9 1 10 0 11 15 1 10 9 1 10 10 9 3 15 4 13 3 10 9 1 9 2
10 10 9 1 10 11 13 3 3 0 2
51 1 10 12 1 10 12 9 15 13 10 0 9 1 10 9 1 10 12 2 0 2 9 15 13 11 1 10 9 1 10 9 0 7 15 4 13 10 0 9 1 10 11 0 1 13 1 10 9 1 11 2
33 10 12 7 10 12 9 10 10 9 1 10 9 2 1 10 9 0 13 3 1 10 11 2 13 1 11 10 9 1 10 9 0 2
16 10 12 9 10 11 0 13 10 9 0 1 10 10 0 9 2
21 10 12 9 10 0 9 1 11 11 7 11 11 11 1 15 3 13 3 11 11 2
44 1 9 10 0 9 0 1 11 15 13 1 11 11 3 1 10 9 1 11 11 11 1 13 10 9 1 9 13 3 12 9 3 3 1 10 9 1 11 1 11 11 7 11 2
26 1 9 1 11 10 9 1 10 9 1 10 9 1 1 10 9 10 9 1 10 9 1 10 9 0 2
27 12 10 9 1 11 3 13 2 1 10 9 1 10 9 15 2 3 16 3 4 4 3 13 3 10 9 2
30 11 3 11 13 10 10 9 7 11 12 9 1 10 11 13 1 11 11 10 9 1 11 1 10 9 0 1 10 9 2
10 11 11 2 13 0 9 7 9 13 2
64 10 9 13 1 2 9 2 2 7 10 9 1 0 9 1 10 9 7 1 10 9 1 10 9 2 12 9 2 7 12 9 2 10 9 1 12 9 7 10 9 1 10 9 1 12 2 2 13 3 1 10 11 11 1 11 2 11 2 4 13 3 3 13 2
34 10 9 2 12 9 2 13 1 10 9 2 4 4 13 1 9 1 9 0 7 4 13 1 10 9 1 4 13 10 9 1 10 9 2
7 15 4 3 13 10 9 2
26 10 9 4 4 13 1 10 9 1 11 7 11 2 15 4 13 10 9 2 1 10 9 1 10 9 2
38 10 9 4 4 13 1 10 9 1 10 9 0 7 0 15 15 4 13 0 7 1 0 9 16 10 9 1 10 9 1 9 4 13 3 10 12 9 2
41 11 11 4 13 1 4 13 10 9 1 10 9 7 1 4 13 10 9 1 15 15 13 13 10 9 0 1 13 1 13 9 7 3 1 4 15 13 1 10 9 2
40 1 3 15 13 3 16 10 9 13 1 10 9 1 9 7 16 10 9 1 10 9 2 11 11 2 13 1 9 1 13 2 10 9 15 4 13 1 10 9 2
18 1 3 10 10 9 4 3 13 0 2 3 10 9 4 13 10 9 2
24 10 9 4 4 13 1 10 9 1 11 3 10 9 4 13 10 10 9 2 15 3 13 9 2
23 2 12 9 1 12 7 12 9 2 1 10 9 2 1 3 12 9 2 2 13 12 9 2
19 4 13 0 13 15 16 4 13 1 10 9 2 4 13 1 11 11 11 2
10 2 13 1 9 2 13 3 1 9 2
8 3 15 13 16 4 4 13 2
33 15 4 13 10 9 2 4 13 9 2 3 1 13 1 10 9 4 13 1 10 15 2 4 13 1 10 9 7 4 9 10 9 2
12 10 9 0 13 0 2 13 2 13 2 13 2
31 10 9 4 13 1 10 9 7 10 9 1 10 9 2 3 15 4 13 9 7 15 4 13 2 7 4 13 1 10 9 2
32 10 9 15 4 13 3 1 10 9 2 10 9 1 10 9 2 7 4 13 0 10 0 9 1 12 9 1 3 12 1 9 2
25 6 1 10 11 1 10 9 2 1 10 9 0 2 1 9 2 11 11 2 9 2 1 10 9 2
13 1 10 9 15 15 13 9 16 10 11 13 2 2
21 2 13 1 10 9 3 0 2 13 13 16 4 13 3 2 4 13 10 9 2 2
11 15 4 13 3 0 2 4 13 3 3 2
8 3 10 9 4 13 10 9 2
13 1 9 1 10 9 13 0 3 13 15 3 2 2
120 2 10 9 0 1 10 9 0 1 10 11 11 4 13 1 1 10 0 9 2 1 9 0 2 3 1 10 11 11 1 10 11 2 1 10 9 2 1 10 9 1 10 9 2 1 10 9 0 1 10 9 7 1 10 9 2 1 10 9 1 9 1 10 9 13 1 10 9 11 7 1 10 12 9 15 13 1 15 2 13 13 2 1 10 9 2 10 11 11 13 16 2 15 4 13 12 9 1 9 0 2 1 15 12 1 9 0 2 1 3 12 9 7 12 3 1 9 7 9 2
14 4 4 3 13 1 9 10 9 0 1 9 0 2 2
44 2 10 9 13 1 12 9 1 10 9 1 15 4 13 10 9 1 10 9 7 1 15 4 3 13 10 9 2 4 13 10 9 1 10 9 1 10 9 1 11 2 11 11 2
23 11 13 1 11 10 9 1 10 12 5 13 1 10 9 0 1 10 9 0 11 1 11 2
10 10 9 4 13 1 10 12 9 12 2
22 11 13 1 11 12 9 1 9 2 1 15 12 9 1 9 7 12 9 1 9 9 2
32 1 10 9 1 10 9 1 9 1 10 9 11 2 13 10 11 1 10 9 2 3 4 13 10 9 1 9 1 9 1 11 2
58 11 11 7 10 11 4 3 13 10 9 1 9 2 1 9 1 10 0 9 0 1 11 11 2 1 10 15 4 13 0 9 1 9 1 11 11 1 10 11 1 10 9 0 0 1 12 9 1 9 1 12 9 0 0 1 9 0 2
43 10 9 1 10 0 9 13 1 9 1 10 9 1 10 9 1 11 7 10 12 0 9 4 13 1 10 12 9 0 1 10 9 1 10 9 1 10 9 1 10 0 9 2
17 11 11 13 1 10 9 1 10 0 9 1 10 9 1 9 0 2
36 2 13 10 9 3 1 10 0 9 2 3 1 3 1 10 12 4 4 13 1 13 1 10 9 1 11 2 13 11 11 2 9 1 11 2 2
24 10 9 2 10 9 7 10 9 13 1 11 1 10 0 12 9 7 9 13 15 1 0 2 2
50 10 9 1 9 1 11 1 10 12 5 1 11 2 15 13 1 13 3 10 10 9 1 13 10 9 1 9 0 1 10 9 1 9 2 9 1 9 7 9 0 1 10 9 2 13 10 9 11 11 2
26 2 1 10 9 1 10 0 9 7 1 10 10 9 15 13 9 0 2 15 13 1 10 9 1 9 2
18 10 9 3 13 1 11 13 1 9 15 1 10 9 1 11 7 1 11
38 13 1 3 0 2 13 11 2 1 10 8 1 8 1 10 9 7 1 10 10 0 9 1 10 13 10 9 1 9 15 3 13 10 10 9 0 2 2
6 9 1 10 11 11 2
31 2 13 3 0 2 1 10 9 16 3 10 9 11 7 11 4 13 10 9 1 10 9 1 10 13 9 1 10 9 11 2
31 3 13 0 1 9 0 13 1 13 2 1 13 2 1 10 9 0 1 13 1 11 7 11 2 13 10 9 0 11 11 2
18 2 10 0 9 15 13 3 10 9 11 13 10 10 9 1 9 9 2
18 10 9 0 1 15 15 13 0 9 3 1 10 11 7 1 11 2 2
17 11 2 11 13 9 1 10 9 10 0 9 1 10 9 1 11 2
16 16 10 11 4 13 1 9 11 2 11 11 4 13 11 11 2
48 10 9 1 10 11 12 11 13 10 0 9 1 10 9 1 10 10 9 1 10 9 13 0 1 4 0 1 13 10 9 1 10 9 1 10 9 1 10 9 1 10 9 1 9 1 11 11 2
30 10 9 3 3 13 1 10 10 9 1 10 9 1 9 1 10 11 2 15 4 13 3 9 0 1 10 9 1 11 2
50 2 10 9 2 1 9 1 9 1 9 2 15 13 10 9 2 15 13 3 10 11 2 15 1 10 12 9 0 1 10 11 2 13 10 9 1 10 9 2 2 15 13 1 10 9 1 10 9 0 2
23 2 13 13 10 0 9 1 10 11 14 11 1 13 10 9 1 9 2 2 13 10 9 2
12 10 9 1 10 9 13 10 9 0 11 11 2
17 2 1 10 9 1 10 9 0 13 10 9 13 10 9 0 2 2
22 10 9 15 13 1 9 1 13 16 2 11 4 13 1 10 9 1 1 10 9 2 2
18 2 10 15 15 13 13 0 7 3 0 2 7 3 13 3 1 15 2
7 10 9 4 13 0 9 2
8 7 10 9 4 13 15 0 2
14 2 1 15 11 13 10 9 1 9 1 10 9 2 2
27 10 9 3 4 3 13 1 10 9 1 10 9 1 11 15 1 10 9 4 13 10 10 9 1 10 9 2
13 13 10 9 1 10 10 9 2 2 13 11 11 2
24 2 3 4 13 1 13 16 2 1 10 9 13 1 10 9 2 15 4 4 13 1 10 9 2
46 2 1 10 10 9 10 9 2 3 0 1 15 15 13 1 10 9 2 13 1 0 9 10 9 15 13 10 9 1 10 9 7 10 9 15 15 13 1 10 9 2 2 13 11 11 2
17 7 15 13 15 15 13 1 10 9 1 10 9 2 1 11 11 2
42 2 10 9 3 13 3 10 9 1 9 2 13 3 10 9 1 13 10 9 1 9 1 15 2 3 1 10 0 9 2 15 4 2 13 2 1 16 3 13 3 13 2
31 13 0 1 10 10 9 13 1 10 8 8 2 15 13 1 10 9 0 1 10 0 9 1 10 0 9 1 10 9 2 2
17 10 9 1 10 9 1 9 1 9 3 13 10 9 9 2 9 2
13 11 11 13 9 1 13 15 2 3 16 13 2 2
27 11 11 3 13 10 9 1 10 9 13 7 15 13 1 10 9 1 10 9 13 1 10 9 1 10 15 2
3 10 9 2
18 10 9 4 13 1 10 9 1 9 7 5 7 1 10 0 9 0 2
41 1 10 0 9 1 10 9 1 15 10 1 10 9 3 1 9 13 2 15 13 7 15 13 1 13 3 10 9 1 10 0 9 1 10 9 1 10 9 12 8 2
30 10 9 13 1 15 10 9 3 1 9 13 1 9 16 15 13 1 13 10 9 7 10 9 1 15 1 10 0 9 2
69 1 10 9 7 1 10 9 1 10 0 9 2 15 13 1 2 11 1 11 2 2 10 9 2 1 10 9 1 10 9 2 10 9 7 10 9 2 1 10 15 10 9 1 10 10 9 7 9 0 2 3 1 0 9 13 15 0 9 0 7 0 2 4 13 1 10 9 0 2
25 10 9 15 13 11 1 11 3 4 13 9 0 2 1 3 13 2 1 10 9 1 10 0 9 2
69 2 9 0 2 2 10 9 0 1 10 9 7 1 10 9 1 1 0 9 0 2 1 10 9 2 10 9 0 2 10 9 0 2 0 2 0 2 10 9 1 9 2 10 9 1 9 2 10 9 2 10 9 2 7 10 0 9 1 15 10 9 4 4 13 2 13 7 13 2
31 1 10 9 1 15 10 9 1 15 3 13 13 3 11 1 11 2 15 3 4 13 9 0 1 10 9 1 10 0 9 2
50 1 10 9 1 13 9 4 13 16 2 16 10 9 13 10 9 0 7 9 1 9 2 10 9 1 10 9 1 9 1 10 9 1 9 2 2 9 2 2 4 13 11 11 1 10 9 1 10 9 2
24 2 11 2 2 10 9 7 10 9 15 13 10 9 1 10 9 7 10 9 1 10 0 9 2
13 2 9 0 2 2 10 9 15 4 13 10 9 2
39 2 11 2 2 10 9 1 10 9 0 1 9 1 9 1 10 9 1 10 9 1 9 2 10 10 9 4 13 1 10 9 1 10 9 1 10 0 9 2
69 2 15 2 5 2 15 2 2 10 9 7 10 9 15 13 10 9 13 1 10 0 9 7 15 3 4 3 13 10 9 1 10 0 9 0 1 10 9 2 7 15 2 1 10 0 9 1 10 15 2 4 13 0 9 1 10 11 1 10 9 1 10 9 13 1 10 0 9 2
26 2 9 1 10 9 2 2 10 9 0 1 10 9 13 1 10 9 7 13 1 10 9 1 10 9 2
8 9 2 13 1 10 0 9 2
5 12 2 0 9 2
54 10 0 9 3 13 1 10 9 13 2 13 7 13 10 9 1 0 9 7 10 13 10 9 1 10 9 1 10 9 7 0 9 1 10 9 0 1 10 9 13 1 10 9 1 10 9 1 9 7 1 0 9 0 2
7 12 2 9 1 10 9 2
59 1 10 9 1 10 9 7 1 10 9 13 1 10 0 9 2 10 11 13 1 15 10 9 1 10 10 9 2 0 2 3 0 7 0 2 1 10 9 1 10 9 1 9 0 2 15 13 1 13 10 9 1 10 9 3 1 9 13 2
29 9 1 10 9 2 9 1 10 9 1 12 7 10 9 1 9 7 9 1 10 9 16 13 1 10 9 1 9 2
8 9 7 9 1 10 11 9 2
55 9 1 9 1 10 9 7 1 9 0 1 15 10 9 4 13 2 9 1 10 9 2 9 2 9 2 9 7 9 1 9 2 3 13 10 9 0 0 1 10 9 2 7 15 3 16 10 9 4 13 1 9 1 9 2
43 9 1 9 1 10 9 7 1 9 0 1 15 10 9 0 4 13 2 9 1 10 9 2 9 2 9 2 9 7 9 1 9 2 3 13 10 9 0 0 1 9 0 2
18 9 1 10 9 1 10 9 7 10 9 7 9 1 9 0 1 9 2
56 10 11 13 1 10 9 0 1 13 9 2 3 7 1 10 9 1 10 9 1 9 0 2 1 9 2 11 2 2 1 10 9 1 10 9 7 10 9 7 9 2 3 1 9 0 2 1 9 2 1 9 2 1 10 9 2
47 10 11 13 1 10 9 0 1 13 9 2 3 7 1 10 9 1 10 9 1 9 0 2 1 9 2 11 2 2 1 10 9 15 15 13 7 13 1 13 1 10 9 2 9 9 2 2
63 1 10 9 1 13 9 2 4 13 16 16 10 9 13 10 9 1 9 2 10 11 13 1 10 9 0 1 13 9 2 3 7 1 10 9 1 10 9 1 9 0 2 1 9 2 11 2 2 1 10 9 1 10 9 1 10 9 2 3 1 9 0 2
8 0 9 13 1 10 9 0 2
62 1 10 11 13 1 10 9 10 9 0 1 15 13 1 10 0 9 2 1 9 2 10 0 9 13 1 10 9 1 9 0 2 0 2 0 7 1 9 1 9 1 9 1 10 9 1 9 1 10 9 1 10 9 12 2 3 9 12 5 12 2 2
18 10 9 3 13 4 4 13 1 10 9 1 9 7 1 10 10 9 2
39 1 10 9 1 15 3 15 13 13 10 9 1 13 1 10 9 10 9 15 15 13 3 0 1 10 9 1 0 9 1 0 9 1 9 7 1 0 9 2
12 10 10 9 3 3 13 1 10 11 13 0 2
23 10 9 13 1 9 1 10 0 9 12 4 3 13 1 2 7 13 1 2 10 0 9 2
97 15 4 13 2 13 1 10 9 2 13 2 13 2 13 7 13 1 9 10 9 2 3 1 9 0 2 3 13 16 10 9 1 15 1 10 0 9 4 13 7 2 1 1 10 9 1 10 9 2 7 9 0 1 15 4 13 10 9 2 15 13 2 13 1 10 9 7 13 2 13 2 13 7 13 1 9 2 3 1 9 0 2 4 13 10 9 1 10 0 9 7 10 10 11 11 11 2
35 3 4 13 7 13 10 9 0 1 10 9 15 13 7 13 10 9 1 10 0 9 7 10 9 1 9 1 10 9 1 10 9 3 13 2
8 3 4 13 10 9 1 9 2
21 4 13 0 10 10 0 15 15 13 1 10 0 9 7 1 10 9 1 10 9 2
55 3 4 13 2 13 1 10 9 2 13 2 13 2 13 7 13 1 9 10 9 2 3 1 9 0 2 13 9 0 13 1 13 10 9 1 10 9 7 10 9 1 10 9 2 1 9 0 1 10 9 1 10 0 9 2
52 15 3 15 13 1 10 9 3 16 15 13 9 1 10 9 1 9 2 3 16 15 3 13 16 10 9 1 9 1 1 15 7 3 1 10 9 0 4 13 0 1 10 9 7 1 10 9 1 10 0 9 2
50 16 15 13 10 9 1 11 2 1 9 1 10 9 2 4 13 1 10 9 1 9 0 2 3 3 0 2 10 9 1 10 11 7 2 1 9 1 10 9 0 2 1 10 9 0 2 1 1 9 2
52 16 15 13 10 9 0 2 1 9 1 10 11 4 13 1 10 9 0 0 2 1 10 9 1 15 15 13 0 2 10 9 1 10 11 7 2 1 9 1 10 11 11 2 1 10 9 0 2 1 1 9 2
50 16 15 13 10 9 1 11 2 1 9 1 10 11 2 4 13 1 10 9 1 9 0 2 3 3 0 2 10 9 1 10 9 7 2 1 9 1 10 11 11 2 1 10 9 0 2 1 1 9 2
52 16 15 13 10 9 0 2 1 9 1 10 11 4 13 1 10 9 0 0 2 1 10 9 1 15 15 13 0 2 10 9 1 10 11 7 2 1 9 1 10 9 0 2 1 10 9 0 2 1 1 9 2
50 16 15 13 2 13 1 10 9 2 13 2 13 2 13 7 13 1 9 2 3 1 9 0 2 10 9 7 10 9 0 7 9 1 9 2 4 13 0 10 10 9 1 10 9 1 9 1 10 9 2
40 4 13 1 10 9 0 10 9 0 1 1 10 9 1 9 7 9 15 13 13 10 9 2 7 10 9 2 16 1 10 9 2 1 10 9 0 2 16 13 2
9 10 9 1 10 9 2 16 13 2
52 1 10 9 1 15 13 3 0 2 10 11 11 11 2 15 10 11 13 4 4 13 1 10 9 2 1 16 10 11 3 13 9 1 10 9 1 9 1 9 1 9 7 3 13 9 1 10 9 1 10 9 2
50 3 2 1 9 1 11 11 2 4 13 10 9 1 10 9 1 10 9 9 2 1 9 2 2 9 0 1 10 9 1 10 9 0 2 2 7 2 9 0 1 10 9 0 1 10 9 0 2 2 2
11 10 9 4 4 13 1 10 9 0 0 2
51 1 10 9 2 1 9 1 9 0 7 9 1 11 2 10 9 13 3 4 13 1 10 0 9 3 4 13 10 9 1 0 9 1 9 0 7 1 10 0 9 13 1 10 9 1 0 9 1 9 0 2
10 12 2 9 2 9 7 9 1 9 2
20 10 9 3 13 10 9 1 9 0 7 3 10 9 4 3 13 15 1 15 2
6 12 2 9 1 9 2
73 0 10 9 13 1 10 9 0 2 10 9 3 13 1 10 9 9 1 10 10 9 1 10 9 1 10 9 1 9 2 13 15 0 2 0 2 0 2 0 7 0 2 13 1 10 0 9 7 1 10 9 1 10 9 2 3 1 10 9 1 15 10 11 4 13 13 1 10 9 1 10 9 2
81 10 0 9 15 13 13 1 9 7 10 9 1 15 13 13 3 2 1 9 1 10 9 1 10 9 1 9 1 10 9 2 1 9 1 10 9 1 10 9 1 10 0 9 1 9 10 2 7 1 9 1 10 9 1 15 1 10 9 12 8 2 12 8 7 12 8 2 13 10 0 9 13 3 1 10 13 15 1 10 9 2
57 1 10 9 2 10 9 1 10 0 9 3 13 10 9 13 1 9 7 9 15 4 13 1 15 9 0 7 9 1 9 2 1 10 9 1 10 0 9 2 1 9 16 10 9 7 9 13 1 13 3 10 9 1 15 13 9 2
25 10 9 12 2 12 2 12 2 12 2 12 7 12 13 0 1 9 1 10 9 1 10 0 9 2
36 3 16 4 13 10 9 7 10 9 1 15 3 2 10 0 9 13 0 2 7 13 1 10 10 9 1 10 9 1 9 1 10 9 0 2 2
35 1 15 2 10 11 15 13 10 9 1 13 10 9 1 10 9 1 10 9 1 10 0 9 7 1 13 10 9 1 10 9 1 10 9 2
64 9 13 16 2 1 10 9 2 10 9 3 13 9 1 10 0 9 2 7 1 10 0 9 15 4 4 13 2 7 15 4 13 16 4 13 2 1 10 9 1 10 0 9 2 2 7 10 0 9 13 1 13 0 9 2 1 16 15 13 9 1 3 13 2
3 12 2 0
52 10 9 16 15 13 2 7 13 2 13 7 13 3 1 9 0 10 9 7 10 9 1 11 2 10 9 13 1 10 9 10 9 1 10 9 1 10 0 9 7 9 15 1 15 4 4 13 1 10 0 9 2
49 10 9 16 15 13 2 7 13 2 13 7 13 3 1 9 0 10 9 9 2 10 11 13 1 10 9 10 9 1 10 9 0 1 10 0 9 7 9 15 1 15 4 4 13 1 10 0 9 2
71 10 9 7 10 9 2 1 10 9 0 2 1 12 7 3 1 10 9 1 10 0 9 2 3 13 10 9 7 10 9 1 10 0 9 7 2 1 9 1 0 9 1 10 9 2 10 9 0 7 0 13 1 13 15 13 1 10 9 1 10 9 15 13 0 1 13 15 0 7 0 2
51 1 10 9 10 9 7 10 9 1 15 1 10 0 9 4 4 13 13 2 7 10 9 4 4 13 13 2 1 16 10 9 7 9 13 1 9 1 10 9 13 1 10 9 1 15 13 10 9 7 9 2
19 10 0 9 13 10 0 9 1 10 9 3 1 10 9 3 13 1 9 2
19 3 13 0 9 2 9 7 9 0 1 10 9 15 3 13 15 3 13 2
20 10 11 3 4 13 1 10 0 9 0 15 4 13 1 10 9 1 15 13 2
18 10 0 9 3 4 4 13 1 10 0 9 13 1 10 11 7 15 2
3 9 11 2
16 10 9 13 9 1 10 9 1 15 10 9 4 13 1 11 2
15 16 15 13 10 9 2 15 13 3 10 9 1 9 0 2
28 1 10 0 9 10 9 15 13 1 13 10 9 1 10 0 11 11 11 0 15 13 1 10 11 11 11 11 2
46 0 11 3 13 0 1 10 10 9 7 1 10 9 1 0 9 1 10 9 1 10 9 2 13 2 1 9 2 10 9 0 2 0 2 0 7 0 15 13 1 9 1 10 0 9 2
40 1 15 13 1 10 12 0 9 2 16 11 11 3 13 15 0 10 9 1 10 9 1 15 1 10 0 9 2 13 10 10 9 7 10 10 9 1 10 9 2
57 1 16 1 10 0 9 1 13 1 10 9 16 10 9 4 13 1 9 1 10 9 1 10 11 2 10 9 4 13 10 9 2 11 11 2 7 10 0 9 13 2 7 10 9 1 11 11 2 1 10 0 9 13 1 11 11 2
48 10 9 13 4 13 1 10 9 1 10 9 9 1 10 9 1 10 9 11 11 2 1 9 1 10 9 2 16 1 9 1 9 13 1 10 9 9 1 11 11 7 3 13 1 9 1 9 2
10 11 11 4 4 13 1 10 9 9 2
5 9 1 10 9 2
31 13 13 10 9 1 10 9 0 2 13 9 12 9 7 13 1 15 10 10 0 9 1 10 9 16 4 13 10 0 9 2
19 16 4 13 9 1 13 10 0 2 9 1 10 9 2 3 15 4 13 2
46 1 10 9 13 10 9 2 1 1 10 9 15 4 4 13 1 10 9 2 13 10 9 1 9 1 9 1 10 10 9 1 10 9 15 15 4 13 1 10 10 9 1 10 11 11 2
16 15 13 3 1 13 15 1 9 1 13 3 10 9 1 9 2
10 2 10 9 13 10 9 1 9 2 2
10 9 9 2 13 1 10 9 1 9 2
25 16 4 13 1 10 9 7 13 1 10 9 2 1 11 11 15 4 13 10 9 7 9 1 9 2
25 15 1 10 9 3 0 4 13 11 11 2 15 10 9 0 4 13 1 9 3 1 10 9 0 2
61 9 9 2 13 0 16 13 10 9 1 10 9 1 10 11 11 1 13 10 9 1 10 9 1 15 7 10 0 9 0 13 15 15 1 11 11 7 1 13 15 1 13 15 1 10 9 1 10 9 1 13 1 10 9 0 1 10 9 3 0 2
14 16 10 9 13 1 9 13 10 9 1 10 9 11 2
9 9 9 2 10 9 1 10 9 2
14 13 13 10 10 9 1 1 10 9 12 1 10 9 2
26 10 10 9 15 13 1 10 9 1 10 9 1 10 9 1 9 7 15 13 1 0 1 10 9 0 2
26 13 16 10 9 13 10 9 0 0 1 10 9 0 1 10 9 7 10 9 13 1 13 15 13 3 0
40 4 13 16 13 0 13 10 9 1 10 9 1 10 9 1 10 0 9 2 7 3 1 10 9 0 2 7 16 13 1 10 10 9 13 10 0 9 9 0 2
31 13 3 1 10 9 15 2 16 15 13 2 13 9 1 13 10 10 9 0 2 7 9 1 9 1 10 9 1 10 9 2
50 9 9 2 1 9 1 10 0 9 10 9 1 10 9 0 2 1 10 11 11 1 11 4 4 13 2 3 1 9 0 2 10 9 1 10 9 1 9 2 10 9 1 12 9 15 13 1 9 11 2
96 1 9 1 10 9 0 2 10 9 11 2 4 3 4 13 10 9 2 15 4 13 10 9 1 15 10 9 2 7 15 13 2 1 9 1 10 9 3 3 9 1 10 9 0 7 1 10 10 9 0 2 1 13 2 1 10 9 1 10 10 9 7 1 10 9 15 15 13 2 1 10 9 7 10 9 1 10 11 11 2 15 13 10 9 1 13 10 9 1 9 7 1 13 10 9 2
13 7 10 15 1 9 1 10 9 15 4 3 13 2
10 15 13 2 9 11 2 15 13 3 2
17 1 9 15 13 3 0 1 10 9 15 10 10 9 4 3 13 2
24 9 9 2 4 13 10 9 1 10 9 15 10 9 13 1 9 2 7 10 9 1 11 11 2
31 15 15 13 0 16 10 9 15 4 13 2 13 16 3 1 11 10 9 1 9 1 10 9 13 10 9 13 1 10 9 2
19 3 2 3 2 4 13 3 1 9 1 9 16 10 0 9 13 1 9 2
65 16 13 7 16 4 13 13 1 0 9 2 3 1 10 0 9 0 1 10 9 0 2 3 15 13 3 1 10 9 0 7 13 10 0 9 13 11 11 1 4 13 9 7 9 0 2 3 15 16 15 2 1 3 9 0 2 4 13 10 9 1 10 10 9 2
18 10 9 13 1 10 9 1 10 9 0 1 9 1 10 9 1 11 2
39 15 13 3 1 13 1 9 10 9 1 10 9 1 15 4 13 10 9 0 7 1 13 1 10 9 0 10 9 13 1 10 9 2 3 1 10 10 9 2
24 3 2 9 11 2 13 3 10 9 0 1 10 9 1 15 0 3 3 4 13 10 10 9 2
22 9 9 2 15 13 1 13 15 1 15 10 10 9 1 4 13 9 1 10 9 0 2
24 1 9 10 9 1 9 0 0 1 10 10 9 4 13 3 1 10 0 9 1 10 9 0 2
16 3 2 9 9 2 3 4 3 4 13 9 1 10 10 9 2
20 13 0 16 3 13 12 9 0 7 10 9 2 7 3 13 3 10 9 0 2
30 7 13 3 15 15 4 13 2 13 16 15 9 0 2 16 4 13 1 10 9 0 2 13 4 13 10 9 1 9 2
8 13 3 10 9 10 10 9 2
28 9 11 2 11 11 2 4 13 15 16 10 9 13 1 10 9 1 10 9 1 10 9 1 10 9 1 9 2
9 13 16 4 13 1 10 9 0 2
23 9 9 2 4 13 16 10 9 3 13 10 9 1 9 1 9 7 9 15 15 0 13 2
22 16 3 4 4 13 10 9 1 10 9 1 10 9 1 10 9 1 16 4 4 13 2
15 16 1 10 12 10 9 9 7 9 3 15 4 3 13 2
24 16 3 4 4 13 9 1 10 9 0 7 1 10 9 1 10 9 1 11 7 3 1 11 2
11 16 3 13 9 1 13 1 9 1 9 2
14 16 1 10 10 9 3 4 4 13 9 1 10 9 2
19 16 3 4 13 13 10 9 1 13 1 10 9 0 3 1 10 3 9 2
15 13 3 0 16 3 15 3 13 10 9 1 15 0 13 2
22 9 11 2 15 13 3 9 7 13 13 16 10 15 15 4 13 3 3 4 4 13 2
34 13 3 13 10 9 1 10 9 1 10 9 7 13 0 16 1 10 10 9 13 1 9 13 1 9 16 10 9 13 10 9 15 13 2
29 9 9 2 10 9 11 11 7 15 4 13 10 9 1 9 1 10 9 1 10 9 11 11 13 1 10 9 0 2
28 10 9 0 3 15 4 13 1 10 9 1 10 9 2 1 3 4 13 16 4 3 13 9 1 10 9 9 2
35 10 9 15 4 4 13 9 1 9 13 10 9 1 10 9 1 11 1 10 9 0 2 3 10 9 13 1 10 9 11 10 12 9 0 2
15 4 13 15 15 1 10 9 10 9 15 13 10 9 0 2
13 7 13 1 0 9 1 13 0 16 15 4 13 2
63 9 9 2 13 13 16 10 9 10 9 13 13 10 9 0 1 13 10 10 0 1 1 10 9 13 3 1 13 10 9 1 10 9 1 10 9 1 10 11 2 13 7 13 16 1 9 10 0 9 1 10 9 4 13 10 9 1 10 9 1 10 11 2
17 10 9 0 1 3 13 15 13 0 2 13 10 9 1 10 9 2
17 10 9 4 3 13 10 9 2 16 13 10 0 9 1 10 9 2
15 10 9 9 1 10 9 4 13 0 1 3 13 10 9 2
28 16 4 3 4 13 2 10 9 1 11 13 3 0 2 1 10 0 9 15 1 9 15 13 10 9 1 9 2
31 3 13 15 4 13 7 3 15 13 16 15 4 13 1 10 9 1 9 1 10 11 1 13 15 9 1 9 1 9 0 2
19 16 13 2 10 9 3 4 13 1 10 9 1 10 9 1 9 1 9 2
5 9 1 10 9 2
70 9 9 2 10 9 16 10 9 11 13 10 10 9 0 1 10 10 9 13 3 1 10 9 1 10 9 1 10 9 1 10 9 0 2 13 1 10 9 1 10 9 1 10 9 1 9 7 3 13 3 1 10 9 11 2 15 4 13 10 10 9 1 10 9 1 10 9 1 9 2
50 15 13 1 10 9 0 1 3 10 9 13 10 9 15 13 10 9 1 9 2 3 1 10 9 2 7 1 9 13 10 9 0 1 15 15 13 10 9 0 7 0 1 10 9 1 10 0 12 9 2
26 13 3 2 9 9 2 16 1 10 0 9 10 9 4 13 12 9 10 9 1 9 1 10 9 11 2
34 1 10 0 9 15 4 13 1 0 1 9 7 3 2 1 10 9 1 10 0 9 2 4 13 3 10 9 1 10 0 9 1 9 2
34 7 15 4 3 13 9 1 9 1 13 1 10 9 1 13 10 10 9 7 1 13 15 1 13 15 9 1 3 13 15 1 10 9 2
25 1 10 9 13 10 9 1 10 12 9 0 2 1 15 15 13 1 13 10 9 10 15 3 0 2
40 10 9 1 10 9 0 2 13 1 8 1 10 9 1 10 9 2 13 3 1 13 7 13 9 13 1 10 1 3 1 15 2 15 13 1 9 1 10 9 2
23 7 10 9 3 13 1 9 1 13 10 9 2 1 10 9 2 13 0 16 15 13 2 2
13 1 13 10 10 9 2 13 1 9 1 13 15 2
35 13 16 10 9 4 13 1 10 9 11 11 2 13 16 1 1 13 13 13 16 10 9 4 3 0 1 13 10 9 2 3 1 10 9 2
17 7 10 9 3 13 1 9 1 13 10 9 2 1 3 13 15 2
46 13 16 10 9 0 4 13 1 9 2 4 13 1 10 9 2 1 3 10 9 3 10 9 7 11 4 13 10 9 1 10 10 9 7 3 10 9 3 13 3 9 1 13 15 15 2
29 1 10 10 9 2 10 9 13 1 13 2 13 7 13 2 3 1 10 9 3 15 13 10 9 15 13 10 9 2
39 16 10 9 13 1 9 1 13 10 9 2 1 15 13 3 1 9 1 13 10 9 0 13 1 10 9 7 10 9 7 13 15 3 1 1 10 10 9 2
45 16 10 9 1 10 9 1 10 9 1 10 9 0 2 1 15 13 2 13 16 9 15 13 10 9 1 10 9 1 10 9 1 10 9 11 2 13 15 3 10 9 1 9 0 2
9 7 4 13 15 1 10 9 0 2
57 1 10 9 16 3 15 13 10 9 2 15 13 1 10 9 10 9 1 10 9 1 10 9 1 13 15 1 10 9 2 7 1 10 15 16 13 9 10 9 1 10 9 2 1 16 10 9 13 3 3 10 9 1 15 15 13 2
24 3 2 9 9 2 15 13 1 13 1 10 9 1 13 15 3 7 3 1 13 1 10 9 2
17 2 9 1 10 9 1 10 9 1 10 9 1 10 9 0 2 2
39 9 9 2 0 9 2 13 3 0 1 10 9 1 10 9 2 9 11 11 2 15 3 13 16 10 9 1 9 4 13 1 10 9 1 10 9 1 9 2
6 3 15 13 1 15 2
9 4 3 13 16 15 4 4 13 2
9 10 9 11 4 13 1 10 9 2
12 1 9 1 9 1 10 9 15 4 13 9 2
14 3 10 9 0 13 10 9 1 15 0 1 10 9 2
9 10 9 4 4 13 1 10 9 2
31 10 9 1 9 4 13 9 1 10 9 1 15 2 16 3 9 2 15 4 13 12 9 0 7 12 1 9 1 10 9 2
13 10 10 15 13 1 10 9 7 3 4 4 13 2
8 4 3 13 3 1 10 9 2
39 13 9 1 10 9 2 1 11 11 7 10 0 9 1 10 10 9 0 2 16 15 13 2 1 10 0 9 4 13 10 9 1 11 11 7 1 10 9 2
55 3 13 3 1 10 9 16 10 9 1 10 9 4 13 1 10 9 1 10 9 0 2 3 3 1 9 1 10 9 13 3 1 10 9 7 3 1 9 1 10 9 13 1 10 9 15 13 10 9 1 10 0 12 9 2
8 7 10 0 9 3 13 3 2
11 10 9 13 10 9 1 10 12 1 9 2
3 4 13 2
16 16 10 9 3 4 13 10 9 12 1 9 15 13 1 9 2
12 3 13 3 10 9 13 1 9 1 10 9 2
20 1 10 9 2 13 16 1 15 0 10 9 7 10 9 4 13 10 9 0 2
32 10 9 2 3 2 13 3 9 1 9 1 10 9 1 10 9 7 3 10 15 15 4 13 1 10 15 4 3 13 15 0 2
21 13 16 1 10 9 1 10 9 0 4 13 15 3 1 10 9 1 10 9 0 2
17 3 13 0 13 15 13 10 9 1 15 3 13 1 9 10 9 2
71 16 13 2 7 13 10 9 16 3 10 9 13 0 1 13 10 9 2 1 13 1 9 10 9 1 0 9 1 10 9 15 15 13 1 1 10 12 2 13 16 1 10 9 10 9 4 13 10 9 15 15 13 2 7 2 3 1 9 2 3 10 9 0 1 10 9 1 10 9 12 2
34 13 3 1 10 9 1 10 9 0 15 13 1 13 3 10 12 9 7 1 10 9 10 10 9 0 13 3 10 9 1 10 9 0 2
35 9 9 2 13 13 3 16 2 1 15 2 10 9 13 10 0 9 1 10 9 1 10 9 1 15 15 1 13 10 10 9 1 10 9 2
58 7 4 13 3 3 15 10 9 11 15 4 13 1 10 9 1 13 10 0 9 2 16 4 13 10 9 11 2 1 1 10 9 0 1 10 9 0 1 10 9 2 1 10 0 9 1 9 1 10 0 9 2 7 1 10 0 9 2
33 13 1 13 2 9 9 2 16 2 1 10 9 13 1 10 9 0 2 10 9 4 13 1 10 9 1 10 9 0 1 10 9 2
26 7 13 13 13 16 2 1 15 13 10 9 2 13 0 7 0 1 13 10 9 16 15 15 13 0 2
35 13 3 0 1 13 15 10 9 2 3 1 10 9 0 2 1 10 9 1 10 9 1 10 9 1 10 9 1 10 9 0 10 9 3 2
61 3 2 9 9 2 13 16 1 9 10 4 13 1 10 9 1 9 1 10 0 9 7 16 13 0 1 13 15 16 13 10 9 2 3 10 9 2 16 13 1 10 9 2 16 10 9 0 13 1 10 9 1 10 12 2 3 16 4 4 13 2
10 9 9 2 13 10 9 1 10 9 2
56 15 4 4 13 16 3 10 9 0 1 10 9 0 13 16 10 9 4 13 1 10 9 1 10 9 2 1 3 1 10 9 1 9 1 9 1 10 9 4 13 10 9 1 10 9 1 9 1 10 9 0 1 10 9 0 2
37 3 13 16 10 9 4 13 2 7 15 1 10 11 2 11 13 3 0 16 10 0 9 4 13 9 15 10 9 15 4 3 13 3 1 10 9 2
8 13 3 10 9 1 10 9 2
25 1 10 9 10 9 1 10 11 2 11 13 16 10 9 1 9 4 13 1 10 9 1 10 9 2
6 15 13 2 9 11 2
11 13 9 10 9 11 15 13 1 10 9 2
45 9 9 2 4 1 15 13 10 9 1 9 1 9 1 10 9 11 15 4 3 13 10 9 1 10 9 0 1 4 13 1 10 9 13 1 10 9 1 10 9 1 10 0 9 2
9 3 2 15 4 13 10 0 9 2
22 15 4 13 7 15 15 4 13 1 9 2 1 10 9 11 2 11 7 10 9 11 2
48 1 10 9 2 10 0 9 9 15 13 2 4 3 13 16 10 9 3 13 3 13 16 13 1 9 7 1 10 9 11 2 7 16 13 10 9 1 13 10 9 15 13 10 9 7 10 9 2
5 3 13 13 3 2
72 3 2 13 10 9 1 13 1 10 9 1 10 9 10 9 0 1 10 9 7 1 10 9 2 1 13 2 10 9 1 15 2 10 9 1 10 12 9 1 10 9 3 0 2 7 15 13 10 9 0 1 10 9 0 2 3 1 10 9 1 10 9 13 1 10 9 1 10 9 1 11 2
29 13 3 1 9 10 9 1 10 9 11 2 11 0 1 13 1 10 9 1 10 9 10 9 0 1 10 9 0 2
18 2 10 9 13 10 9 1 12 9 0 2 12 9 7 12 13 2 2
19 9 9 2 13 10 9 11 1 10 0 9 15 4 3 13 1 10 9 2
2 3 2
23 9 9 2 4 4 13 10 10 9 2 15 3 4 4 13 3 2 16 3 13 10 9 2
6 10 10 9 13 0 2
14 9 9 2 10 9 4 3 13 10 9 1 10 9 2
5 3 4 13 9 2
50 9 9 2 13 16 13 10 10 9 2 7 1 10 9 0 1 10 9 1 10 9 0 1 10 9 4 13 10 9 1 13 1 9 1 10 10 9 1 1 10 9 2 7 3 15 4 13 10 9 2
31 15 13 3 0 16 1 1 13 10 9 1 10 9 1 10 9 15 13 1 13 10 9 1 9 1 9 1 10 10 9 2
34 15 13 1 10 9 0 7 13 0 4 13 1 9 10 9 1 10 10 9 1 10 9 1 10 9 1 10 9 1 10 10 9 0 2
30 9 9 2 3 13 10 9 13 10 9 2 7 3 15 4 13 1 13 1 13 9 1 10 9 1 10 9 11 11 2
8 15 3 15 4 13 10 9 2
26 15 13 0 3 16 3 10 9 4 3 4 13 2 10 9 13 7 3 10 9 13 1 13 15 13 2
19 15 15 13 2 9 11 7 11 2 3 15 4 13 16 4 13 10 9 2
16 16 15 13 16 10 9 13 0 7 4 13 1 10 9 0 2
24 16 3 13 10 9 0 1 10 9 0 10 9 15 4 13 15 0 4 13 16 15 4 13 2
6 15 13 10 0 9 2
16 3 10 9 0 1 10 9 1 9 13 10 10 0 9 0 2
20 15 13 10 9 0 1 15 13 3 1 10 9 1 9 15 15 13 3 3 2
10 9 11 2 9 11 2 13 1 9 2
19 9 9 2 16 10 9 13 3 10 9 1 10 10 9 3 13 10 9 2
21 7 16 10 10 9 13 16 3 4 13 10 9 1 9 2 15 13 1 10 9 2
18 13 10 9 3 1 10 9 1 10 9 0 2 1 1 15 13 3 2
11 16 15 3 13 3 10 9 4 4 13 2
13 2 10 9 13 10 9 1 10 9 3 13 2 2
11 9 1 10 9 1 10 9 1 9 0 2
104 10 9 1 10 9 13 10 9 1 10 9 2 11 5 12 2 2 13 1 10 9 11 1 9 1 10 9 1 10 9 0 2 10 9 7 10 9 2 1 10 9 0 13 1 10 9 1 9 1 10 9 1 10 9 1 10 9 0 7 1 10 9 0 1 10 9 0 0 1 10 9 1 9 1 10 9 1 10 9 1 9 2 1 9 7 1 9 0 1 9 0 2 11 5 12 2 12 5 12 2 11 2 2 2
63 9 9 2 3 4 7 3 4 13 15 1 10 0 9 1 10 9 15 15 13 1 10 9 1 9 2 1 9 7 1 10 9 0 1 0 9 2 13 3 3 7 3 1 10 9 16 10 0 9 3 15 13 1 0 9 1 10 9 1 10 9 0 2
35 13 3 16 2 1 9 7 0 9 1 10 9 7 1 0 9 1 10 0 9 1 9 2 10 0 9 15 13 1 10 9 1 0 9 2
70 13 0 15 4 13 13 3 1 10 9 2 7 13 10 15 13 1 15 15 2 10 9 1 10 9 1 10 9 11 15 4 13 10 9 1 10 9 7 1 15 3 1 10 9 7 1 10 0 9 0 15 4 4 13 16 4 4 13 1 10 9 1 10 9 1 9 1 10 9 2
31 10 9 1 9 2 13 9 2 4 13 10 9 1 10 9 1 10 0 9 1 9 1 10 9 7 10 9 1 10 11 2
26 10 9 1 10 9 13 15 0 4 13 9 1 10 9 1 10 9 1 9 1 9 1 10 11 11 2
14 1 10 9 1 10 10 9 10 9 4 13 3 0 2
48 10 10 9 1 9 1 10 9 4 13 10 9 7 10 9 1 9 3 1 9 13 10 0 9 1 13 10 0 9 1 10 9 1 10 9 2 16 15 13 1 10 9 7 1 10 9 0 2
18 3 3 4 13 15 1 13 10 9 0 13 1 13 10 9 1 9 2
26 4 3 13 15 15 10 9 13 4 13 3 1 10 9 9 7 2 3 3 2 15 15 4 3 13 2
25 13 2 1 9 2 15 15 13 10 0 9 1 15 15 13 1 10 4 13 10 9 1 10 9 2
41 3 4 13 15 1 13 10 0 9 1 10 9 1 9 2 13 10 9 1 10 9 15 13 1 13 3 1 3 1 9 1 9 1 10 9 1 10 9 1 11 2
51 1 10 9 13 1 10 9 9 0 2 7 3 0 2 1 13 1 10 15 3 10 9 1 9 2 16 1 9 15 4 13 0 9 1 10 9 1 9 1 3 4 3 13 1 11 1 9 1 10 9 2
57 9 9 2 3 15 4 13 10 9 11 1 10 10 9 13 1 10 9 1 10 9 1 10 9 7 1 9 1 10 9 1 10 9 0 1 10 9 1 9 1 10 9 1 10 9 1 9 0 1 9 2 9 7 9 9 0 2
9 15 13 1 15 1 10 0 9 2
44 10 10 9 15 4 13 1 10 0 12 9 7 15 13 16 10 9 1 10 9 3 4 3 4 13 1 13 7 15 10 9 1 10 9 1 10 9 4 4 3 0 7 0 2
37 10 9 13 16 2 1 10 10 9 0 2 10 9 4 13 12 1 10 12 9 13 1 10 9 1 0 9 7 4 13 10 9 1 10 12 13 2
42 3 10 10 9 13 13 1 9 1 10 0 9 0 7 13 1 3 10 9 1 10 9 15 15 13 1 10 0 9 1 13 10 9 1 10 11 11 10 3 0 0 2
19 10 10 9 13 3 1 9 1 10 9 13 1 13 10 9 1 10 9 2
20 10 9 1 13 1 10 9 13 3 3 2 16 4 13 10 9 13 15 3 2
12 9 9 2 15 13 1 13 10 9 1 9 2
30 13 3 15 10 9 1 10 10 9 3 0 7 0 1 10 9 1 9 2 7 1 0 9 10 9 1 10 9 13 2
30 10 9 13 10 9 1 10 9 1 9 2 3 2 1 9 13 3 1 9 0 2 15 15 15 1 10 0 9 13 2
16 10 15 13 0 2 7 3 0 13 10 9 1 10 9 13 2
37 15 13 10 9 1 13 9 1 10 9 2 13 13 10 9 15 4 13 1 10 9 0 1 9 1 9 1 11 2 7 1 11 7 1 0 9 2
33 15 13 10 9 1 15 4 13 13 9 15 13 9 0 7 15 1 10 9 0 3 4 4 13 1 1 13 15 3 1 10 9 2
20 7 13 1 10 9 13 1 10 9 1 10 11 0 15 13 1 9 3 0 2
39 1 9 0 1 10 9 0 2 0 7 3 0 4 3 13 16 10 12 9 1 10 9 13 1 9 9 0 2 3 4 13 1 10 9 1 10 9 13 2
11 1 0 2 10 9 1 10 9 13 0 2
35 1 15 13 1 10 9 1 10 9 1 10 9 2 1 10 9 9 1 13 1 10 0 9 1 10 9 10 9 4 3 13 15 15 0 2
25 3 10 9 13 1 10 9 13 15 2 3 1 10 9 3 0 2 15 3 13 1 9 0 0 2
29 1 9 10 9 4 13 1 13 1 10 10 9 7 1 13 15 1 10 0 9 2 1 10 0 9 15 15 13 2
45 1 10 9 15 13 1 10 9 1 13 10 9 1 10 9 0 2 7 1 10 9 0 2 1 13 3 1 9 11 12 10 9 0 13 0 2 3 4 13 15 1 10 10 9 2
16 13 15 1 13 10 0 9 2 3 13 10 9 1 10 9 2
39 13 13 10 9 0 1 10 9 1 10 11 0 2 13 16 15 13 1 10 9 1 9 3 1 13 1 10 0 9 12 2 7 3 1 10 9 7 9 2
16 10 9 3 13 1 10 0 9 0 2 10 15 3 13 0 2
46 3 2 15 13 16 15 4 13 10 9 1 10 9 15 13 10 9 1 10 9 0 2 0 7 1 9 9 0 2 7 13 3 10 9 1 10 9 0 1 10 9 13 1 10 9 2
26 9 9 2 1 10 9 2 1 9 1 15 2 15 13 3 1 9 10 9 1 10 9 1 10 9 2
31 10 9 3 0 1 9 15 13 10 11 13 2 3 7 3 2 13 1 10 10 9 1 10 9 2 10 9 7 10 9 2
15 3 2 15 15 4 13 10 0 9 4 13 9 3 0 2
34 10 9 13 1 10 0 9 2 10 9 12 5 12 5 11 2 13 3 0 1 13 10 9 0 1 10 9 1 10 9 1 9 0 2
49 15 13 16 15 4 13 10 9 1 10 9 1 9 1 9 0 1 10 9 1 10 9 1 10 9 2 16 4 13 16 4 4 13 9 7 9 0 9 1 13 10 9 1 10 9 1 9 0 2
12 3 2 13 16 10 15 13 3 10 0 9 2
22 3 2 10 9 13 1 10 9 13 15 10 9 7 3 4 13 1 10 10 10 9 2
23 9 9 2 9 9 2 0 9 2 1 15 4 13 15 1 10 9 11 1 10 9 13 2
21 3 13 15 1 9 1 9 0 2 13 0 9 1 10 9 1 9 1 10 9 2
6 15 13 1 10 9 2
52 1 0 9 4 13 10 9 9 2 7 4 13 16 10 10 9 13 10 9 0 2 1 13 15 16 4 13 0 9 1 10 9 1 10 9 1 10 9 1 9 2 7 1 10 9 0 7 1 10 9 0 2
46 13 16 10 0 9 1 10 9 4 4 13 10 12 9 12 7 15 3 15 15 4 3 13 2 16 10 9 15 4 13 1 10 0 9 2 4 13 13 16 15 4 13 1 0 9 2
26 15 3 4 13 3 1 10 9 7 9 15 4 13 15 3 3 1 13 1 10 9 3 1 10 9 2
25 1 9 13 1 10 9 16 1 10 9 1 10 9 1 10 9 13 0 10 0 9 7 9 0 2
31 1 15 13 10 9 3 13 3 0 1 3 10 9 1 11 3 13 3 15 1 10 9 1 11 2 1 11 7 1 11 2
17 4 3 13 10 9 0 2 7 13 10 9 1 13 10 0 9 2
9 3 10 0 9 4 3 4 13 2
22 3 15 2 1 10 9 11 2 13 1 10 9 1 9 1 15 10 9 13 0 9 2
22 3 15 13 1 13 3 10 9 1 9 1 10 9 2 13 9 1 9 1 10 11 2
35 13 3 15 13 13 10 15 15 13 1 10 10 9 1 9 10 3 0 10 9 1 9 0 1 10 10 9 2 13 15 1 9 7 3 2
40 1 10 9 15 13 10 0 9 2 0 1 10 9 0 1 10 9 0 1 10 9 1 10 9 1 10 9 1 9 0 1 9 2 1 9 7 1 9 0 2
45 1 10 9 2 13 0 10 9 7 10 9 13 3 1 10 12 9 2 9 7 9 2 7 10 9 13 1 10 9 1 10 9 0 2 7 1 9 1 10 9 13 2 13 0 2
27 10 9 0 13 3 10 10 9 13 1 10 9 7 13 10 9 0 0 1 10 9 1 9 1 10 9 2
41 1 0 9 2 4 3 13 10 9 0 1 10 9 1 9 13 2 3 3 0 1 1 15 13 3 1 10 9 2 13 16 13 3 0 9 15 13 1 10 9 2
30 13 3 13 3 10 0 9 1 10 10 9 7 13 15 15 1 10 9 10 9 13 10 9 1 10 9 1 10 9 2
24 7 16 4 13 3 3 10 9 11 2 10 9 3 15 4 3 13 1 13 2 13 7 13 2
26 10 9 1 10 9 2 1 10 9 1 9 1 10 9 13 10 9 15 4 13 1 13 9 1 9 2
24 1 10 9 2 13 3 13 3 9 1 10 9 1 10 9 2 13 1 10 9 11 7 11 2
28 1 10 9 1 10 11 2 15 13 3 1 10 9 3 0 2 15 13 10 9 1 13 16 13 15 10 9 2
20 1 15 1 10 0 9 13 15 3 2 10 9 13 3 13 1 1 15 0 2
24 10 9 7 10 9 1 9 15 2 1 9 1 0 2 3 13 9 2 4 13 10 0 9 2
17 13 0 3 13 16 13 0 13 3 10 9 1 13 10 0 9 2
15 3 2 13 16 4 13 10 9 1 10 10 9 1 9 2
46 10 9 13 1 10 9 10 9 1 10 9 1 10 9 0 2 1 9 1 10 9 1 10 11 2 7 1 10 9 1 10 9 4 13 1 10 9 1 9 1 9 1 10 9 0 2
15 7 2 0 9 2 10 9 13 10 9 0 1 10 9 2
60 16 13 9 1 13 1 10 9 1 10 9 1 10 11 2 3 13 10 9 1 13 15 1 10 9 1 10 9 1 10 9 2 7 15 13 1 13 1 10 9 2 15 3 13 15 16 13 15 13 0 13 10 9 0 1 10 9 1 9 2
18 13 3 10 9 10 15 15 4 13 2 7 1 9 10 9 9 11 2
5 10 9 4 13 2
10 10 9 15 13 3 2 1 10 12 2
7 9 1 9 0 1 9 2
93 10 9 1 10 9 13 10 9 2 11 5 12 2 13 1 10 9 11 1 9 1 10 9 1 10 9 0 2 10 9 7 10 9 1 10 9 1 9 1 10 9 0 7 1 10 9 2 11 2 12 2 12 2 11 5 12 2 12 5 12 2 11 2 2 15 13 10 9 12 5 12 5 11 13 10 9 1 10 9 1 10 9 9 0 1 10 9 1 9 0 1 9 2
69 9 9 2 9 9 2 0 9 2 10 9 13 1 9 10 0 9 12 13 10 9 1 10 9 1 10 9 9 0 1 10 9 1 9 0 1 9 13 10 9 0 10 10 9 13 1 9 7 13 1 10 9 1 10 9 1 9 1 9 1 10 11 2 10 9 0 1 9 2
19 10 9 1 10 9 1 10 11 4 13 9 1 10 9 1 10 0 9 2
22 1 9 2 10 9 3 4 4 4 13 1 10 3 0 9 1 10 9 0 7 0 2
17 15 13 1 10 9 0 7 15 13 1 13 1 13 1 9 10 2
18 13 3 10 9 1 9 1 10 9 12 5 12 5 11 3 1 9 2
45 10 0 9 1 9 1 10 11 11 13 10 9 9 1 13 10 10 9 0 9 1 10 0 9 2 7 1 1 10 9 1 10 9 1 10 11 2 10 15 13 0 9 7 9 2
34 10 9 1 10 9 3 1 9 3 13 10 9 1 10 9 3 13 1 10 9 1 10 9 1 10 9 1 9 1 9 1 9 0 2
29 15 15 13 1 13 10 9 0 13 10 9 2 1 13 10 9 13 3 0 7 1 13 10 9 1 10 0 9 2
9 8 2 9 8 8 1 9 0 2
29 8 2 9 1 9 0 3 0 2 1 9 1 15 13 10 9 1 9 3 0 1 9 0 1 9 0 3 13 2
15 10 9 1 10 9 13 3 3 0 1 10 9 1 9 2
9 1 10 9 9 4 13 0 9 2
36 10 9 13 16 10 9 9 4 13 10 9 2 13 1 10 9 1 10 9 1 9 1 10 9 1 10 9 0 1 10 9 1 10 9 0 2
66 10 9 1 10 9 1 10 9 1 9 1 9 1 10 9 4 4 13 1 10 9 1 10 9 1 10 9 12 10 9 1 9 13 10 9 1 9 0 1 9 3 1 9 13 3 1 10 9 12 7 2 3 2 3 4 4 13 9 1 10 9 1 9 3 13 2
26 10 9 13 7 13 1 10 9 1 9 1 9 13 9 1 12 9 1 10 0 9 1 9 3 13 2
36 13 13 16 10 9 13 3 1 10 9 7 16 10 9 13 1 9 0 1 10 15 10 9 4 13 10 9 4 13 1 10 9 1 12 9 2
10 15 13 3 10 9 1 10 0 9 2
39 10 0 9 13 1 10 9 9 1 13 9 3 0 2 3 1 10 9 16 10 9 9 1 10 15 15 13 7 15 13 10 9 13 1 9 0 1 12 2
15 15 1 10 9 2 3 2 1 10 9 1 10 11 0 2
54 10 0 9 15 13 1 13 16 13 1 4 13 1 10 9 0 9 7 9 13 1 10 9 0 1 10 0 9 12 7 10 9 1 9 1 10 9 2 10 10 9 7 9 13 1 9 1 10 9 1 10 0 9 2
25 3 13 16 15 13 3 1 10 0 9 1 10 0 9 2 15 9 1 13 1 9 1 10 9 2
37 13 10 0 9 15 13 1 11 7 4 13 1 13 3 0 2 10 9 16 13 1 10 0 9 15 3 2 1 9 2 4 13 15 1 12 9 2
10 13 13 0 16 10 9 4 13 3 2
44 7 10 9 9 4 13 1 13 10 10 9 0 1 10 9 1 9 3 0 7 15 13 3 9 0 7 2 3 10 9 2 13 10 9 1 10 9 1 10 9 1 10 11 2
27 1 0 9 2 1 10 9 1 10 9 3 4 13 1 9 10 9 2 1 10 9 0 1 10 9 0 2
27 4 13 3 0 13 10 9 1 13 1 10 0 9 1 10 9 11 2 15 4 4 13 1 9 1 9 2
21 10 9 13 10 9 1 10 0 9 1 10 9 13 1 10 9 1 10 9 0 2
17 1 10 9 1 10 9 15 4 13 16 3 12 9 4 13 0 2
24 1 15 15 13 1 10 9 1 10 11 13 0 13 16 1 11 10 9 4 13 3 0 9 2
25 0 9 2 3 1 11 15 13 10 9 1 10 11 11 2 3 13 0 13 3 9 1 10 9 2
14 1 9 2 4 13 1 13 10 9 1 3 12 9 2
19 10 9 13 0 3 1 13 0 10 9 1 9 1 9 1 10 9 0 2
18 13 16 10 10 9 4 13 1 9 1 10 9 1 10 9 1 9 2
5 15 4 13 0 2
48 13 1 10 9 2 13 16 10 9 0 4 4 13 0 16 10 9 1 11 1 9 2 1 9 7 1 0 9 2 13 1 9 1 0 9 2 3 1 10 9 1 15 15 13 1 9 0 2
10 10 0 9 13 10 9 1 10 9 2
17 10 9 16 3 4 13 1 13 13 2 1 9 1 9 2 0 2
56 10 9 2 9 11 2 1 10 15 13 10 10 9 1 10 9 13 2 4 13 13 16 4 3 4 4 13 10 9 16 3 15 4 13 9 1 10 9 1 10 11 13 1 10 9 1 10 9 7 1 10 9 1 10 9 2
57 3 15 13 3 16 13 2 1 10 9 4 13 10 15 2 15 1 10 12 4 3 13 1 9 0 1 9 1 9 1 9 0 1 9 2 13 1 10 9 7 1 10 0 9 1 10 9 7 1 10 0 9 1 10 10 9 2
19 9 9 2 10 9 15 13 3 3 13 2 1 15 2 9 1 0 9 2
57 10 0 9 1 10 9 13 1 9 3 0 2 7 13 3 10 9 1 13 16 2 10 9 16 13 9 1 10 9 2 15 13 1 9 1 10 9 1 9 0 2 1 10 9 1 13 9 0 1 10 0 9 1 10 9 0 2
29 1 10 0 9 1 10 9 4 13 0 9 1 9 0 2 15 13 1 10 9 2 1 10 9 7 1 10 9 2
15 15 13 0 10 9 1 10 0 9 1 10 9 1 9 2
20 9 1 9 2 15 13 1 10 9 0 1 9 0 15 10 9 9 4 13 2
8 15 13 15 10 9 3 0 2
16 10 9 1 10 9 13 0 3 1 10 9 1 10 9 0 2
44 16 15 13 2 3 2 16 10 9 0 1 10 9 4 13 3 2 13 3 0 3 3 13 15 1 9 2 7 3 13 16 10 9 13 2 1 10 0 9 0 2 9 0 2
25 1 9 2 13 13 10 0 9 2 3 1 0 9 2 1 9 1 10 9 13 1 10 9 11 2
12 10 9 0 13 3 1 10 9 1 10 15 2
23 15 13 0 2 1 10 9 2 13 9 1 10 0 9 1 9 3 0 1 9 7 9 2
17 9 9 2 1 10 9 1 9 13 3 0 13 15 1 13 0 2
10 13 3 16 10 9 4 13 10 9 2
47 9 9 2 4 13 3 3 10 9 2 9 11 2 7 3 10 9 1 10 9 1 4 13 1 9 3 0 7 0 10 9 1 10 9 1 10 9 1 10 9 7 10 9 1 10 9 2
37 10 9 11 4 4 13 10 10 0 9 1 3 10 9 1 10 11 7 3 15 1 10 9 0 1 10 11 11 3 4 4 13 1 10 13 9 2
18 3 13 1 15 0 13 9 15 13 1 10 1 3 1 10 9 0 2
42 16 10 9 9 3 13 1 9 1 13 15 3 2 4 3 0 1 13 1 9 10 9 0 1 10 9 1 10 9 7 1 10 9 1 10 9 1 11 7 9 0 2
42 9 9 2 15 13 3 1 10 9 11 1 10 9 13 1 9 1 10 0 9 15 2 1 10 0 15 9 2 13 10 9 15 4 13 10 0 9 1 10 9 0 2
29 10 9 7 10 9 1 10 9 3 1 9 15 13 1 13 9 1 9 1 9 15 13 10 9 1 10 10 11 2
24 3 3 10 9 11 15 13 1 9 0 3 1 12 9 1 12 2 7 1 12 9 1 12 2
9 3 13 10 9 2 13 3 9 2
43 13 16 15 4 13 9 1 9 0 2 15 13 10 9 0 1 10 11 11 7 15 3 15 13 3 1 9 7 9 0 2 16 15 13 1 13 9 7 9 1 9 0 2
58 1 9 1 15 4 13 10 9 11 1 10 9 1 10 11 2 4 13 16 10 9 4 13 1 10 9 2 1 3 13 0 16 2 1 10 0 9 2 1 3 15 1 10 9 15 13 1 9 1 10 0 9 16 3 15 4 13 2
56 3 2 9 9 2 4 3 4 13 10 9 0 15 13 10 9 1 10 9 2 4 13 10 9 1 10 11 2 10 9 1 10 9 2 10 9 1 10 9 1 10 9 7 10 9 1 10 9 2 10 9 1 10 0 9 2
32 10 10 9 1 10 9 0 7 1 10 9 2 9 11 2 13 1 0 9 2 15 13 3 12 2 4 4 13 1 10 9 2
11 7 13 10 12 9 15 15 4 4 13 2
5 10 9 4 13 2
10 10 9 15 13 3 2 1 10 12 2
8 9 11 0 5 11 1 9 2
84 10 9 1 10 9 13 10 9 2 11 5 12 2 13 1 10 9 11 1 9 1 10 9 1 10 9 0 2 10 9 7 10 9 1 10 9 1 10 9 0 1 10 9 0 7 1 10 9 1 10 9 1 9 2 11 9 1 10 9 1 10 9 12 2 12 2 11 2 12 2 12 2 11 5 12 2 12 5 12 2 11 2 2 2
43 9 9 2 13 1 15 10 0 9 4 13 10 10 0 9 1 10 9 0 1 10 9 13 10 3 0 1 10 9 1 10 11 11 15 15 13 1 10 9 2 10 11 2
30 16 3 13 2 0 9 1 10 11 4 13 10 9 1 9 1 10 9 12 1 10 9 1 10 9 1 10 9 0 2
35 13 3 0 16 15 1 11 13 1 10 9 0 1 10 9 0 1 1 10 9 1 13 15 1 10 3 0 9 15 3 4 13 1 13 2
27 10 9 1 11 13 1 9 2 7 1 10 12 4 3 13 2 16 10 9 1 0 7 0 15 4 13 2
30 3 1 10 9 1 10 9 0 3 15 13 3 10 9 0 2 7 3 10 0 9 1 10 0 9 0 1 10 11 2
29 3 2 10 9 16 10 9 1 10 9 0 13 1 10 9 10 9 1 10 9 0 13 10 9 15 15 13 3 2
18 1 9 2 3 3 13 15 16 10 9 1 10 0 9 1 10 11 2
25 15 13 10 9 1 15 13 1 13 1 9 15 1 10 9 15 1 10 9 10 9 4 13 0 2
13 15 13 16 10 9 13 10 9 13 1 10 9 2
23 13 16 10 9 1 10 9 4 4 13 1 10 9 1 10 9 0 1 10 10 11 11 2
15 15 13 3 16 10 9 13 10 0 9 1 10 0 9 2
42 15 13 16 13 1 10 9 0 10 9 1 10 9 0 1 10 9 1 9 2 9 15 1 9 4 13 10 9 0 1 10 9 1 10 9 1 9 1 10 9 0 2
22 3 2 13 1 10 9 1 13 16 10 9 13 1 10 9 0 4 13 1 9 0 2
11 10 9 1 10 9 3 13 1 9 0 2
16 13 16 1 10 9 10 9 4 13 10 0 9 1 10 11 2
19 9 9 2 10 10 9 4 13 10 9 2 13 15 1 10 9 1 9 2
11 13 10 10 9 13 15 10 9 10 9 2
80 10 10 9 13 3 0 10 9 16 10 9 4 13 1 10 9 10 10 9 1 13 10 9 1 10 9 1 10 9 9 1 10 9 1 9 2 13 3 1 10 9 7 1 10 9 1 9 1 9 1 13 15 1 3 13 10 9 1 10 9 1 10 9 3 0 7 1 13 3 16 10 9 13 1 10 10 9 1 9 2
21 10 9 0 13 0 7 10 9 1 10 9 0 13 3 1 13 10 9 1 9 2
14 10 0 9 15 13 13 4 3 13 1 10 9 0 2
45 1 10 9 1 10 9 1 10 9 0 7 1 10 9 1 9 2 10 9 4 4 13 3 1 9 10 9 1 10 9 2 1 10 9 0 7 1 10 9 1 10 9 1 9 2
18 1 9 10 9 7 10 9 13 3 1 10 9 1 10 9 0 0 2
13 10 9 1 0 9 0 4 2 3 2 13 9 2
21 3 10 9 13 3 15 2 3 4 13 1 10 9 2 7 10 9 15 4 13 2
23 13 3 0 13 1 0 9 2 1 10 0 9 0 7 1 10 9 2 15 13 10 9 2
20 15 2 1 10 9 2 4 4 3 13 1 10 9 0 15 4 13 10 9 2
27 10 9 1 10 9 2 10 9 0 2 10 9 7 10 9 13 3 10 9 1 13 0 9 1 10 9 2
37 3 2 1 9 1 9 1 10 9 2 4 4 13 10 0 9 0 1 10 9 0 0 1 10 9 1 10 9 0 7 1 10 9 1 9 0 2
26 1 10 9 4 4 13 10 0 9 1 10 9 0 0 2 13 10 9 0 1 10 9 1 9 0 2
17 9 9 2 10 10 3 0 9 1 10 9 11 1 10 9 13 2
41 13 13 10 10 9 1 10 9 9 12 7 12 2 13 1 9 1 9 1 10 9 7 10 9 0 2 7 3 1 9 1 10 9 0 2 10 9 7 10 9 2
39 10 9 13 1 10 9 0 7 1 10 9 1 13 9 0 1 9 7 1 13 9 0 1 10 9 0 13 1 13 9 1 9 7 1 13 10 9 0 2
18 1 9 10 9 4 13 10 0 9 1 9 1 9 1 10 9 0 2
26 3 10 0 9 13 1 10 9 1 10 9 1 15 10 9 0 13 10 0 9 15 13 10 9 0 2
29 13 16 15 15 4 13 1 13 1 10 9 13 9 3 0 1 13 1 10 9 7 1 10 9 1 9 1 9 2
32 1 10 10 9 2 10 9 11 13 3 1 9 10 9 1 15 13 10 0 9 1 9 2 1 15 3 15 13 10 0 9 2
30 10 9 1 10 9 15 13 1 10 12 9 1 10 9 1 10 9 7 1 10 12 9 1 9 1 10 9 0 0 2
47 10 9 1 9 9 0 3 15 13 13 1 0 9 2 13 16 10 9 1 13 10 9 1 10 9 0 1 10 9 1 10 9 4 13 1 10 0 9 1 10 9 1 9 12 2 12 2
30 13 16 10 9 15 4 13 16 15 4 13 1 10 9 1 10 9 1 10 15 15 4 13 1 10 9 1 9 0 2
37 9 9 2 9 9 2 0 9 2 10 9 13 1 10 9 3 1 10 10 9 13 10 9 1 9 0 1 10 9 1 10 9 7 10 9 0 2
18 15 3 13 1 13 16 10 9 1 9 15 13 10 9 15 15 13 2
45 13 1 9 16 10 9 3 13 10 9 0 1 9 1 10 9 1 9 1 10 10 9 0 2 13 10 0 9 1 9 1 10 9 0 1 10 0 9 1 9 1 10 9 0 2
41 10 9 2 1 1 10 9 1 10 9 1 9 7 9 7 1 10 9 1 9 1 9 3 0 7 1 10 9 0 7 3 0 2 13 10 9 1 10 9 0 2
5 10 9 13 0 2
35 1 13 15 15 13 10 9 2 15 15 13 10 9 7 13 10 9 1 10 1 3 1 10 9 0 2 7 15 15 13 3 1 1 15 2
22 10 9 1 9 13 10 9 3 1 10 9 1 9 7 1 10 9 1 9 1 9 2
20 3 4 13 16 10 9 0 13 3 10 12 0 1 10 9 1 10 11 11 2
22 3 2 12 0 1 10 10 9 13 9 2 9 7 13 9 1 13 3 10 10 9 2
73 1 10 9 2 1 10 9 0 15 4 13 15 1 10 11 11 13 10 9 1 13 0 9 1 9 1 10 9 0 2 1 10 1 3 1 10 9 0 2 1 9 1 10 9 0 2 10 9 2 10 9 2 10 9 1 10 9 2 10 9 7 9 1 9 2 10 0 9 2 10 9 2 3
64 15 1 2 3 3 13 0 10 9 1 10 9 2 9 0 1 13 10 9 0 7 0 1 10 9 0 7 10 9 1 0 9 9 2 16 3 15 3 16 10 9 13 10 9 0 1 10 9 1 10 9 2 10 9 1 10 9 7 10 9 1 10 9 2
18 7 13 1 9 1 10 9 0 7 1 9 0 0 1 10 9 13 2
32 1 10 9 1 10 0 9 10 9 0 4 13 0 7 0 7 1 10 9 0 7 13 15 1 10 9 1 10 9 3 0 2
63 13 0 13 9 0 1 9 1 10 9 7 1 9 1 10 9 2 7 13 9 1 10 9 1 10 9 1 10 9 7 10 9 0 0 1 12 9 0 2 13 3 1 9 1 10 9 1 10 9 2 10 9 0 7 10 9 1 10 9 12 7 12 2
26 13 2 13 1 10 9 1 13 9 1 10 12 9 16 15 13 1 13 10 9 0 1 10 12 9 2
24 13 3 16 1 10 11 11 10 9 1 10 9 1 10 9 0 4 13 15 1 10 9 0 2
28 9 9 2 9 9 2 0 9 2 13 1 15 13 10 9 9 11 1 10 9 13 2 1 10 9 2 3 2
58 15 13 3 1 10 9 1 10 9 15 4 13 1 10 9 1 10 0 9 0 2 16 15 4 13 1 13 9 1 9 1 9 1 10 9 1 9 2 3 3 10 1 10 13 2 7 15 1 9 13 10 9 1 10 9 1 9 2
46 1 15 13 0 16 10 9 13 1 10 9 1 10 9 4 13 1 9 1 10 9 2 15 3 1 10 9 2 16 1 10 9 4 13 16 3 4 13 3 10 9 0 2 3 0 2
46 10 9 13 16 13 13 2 7 15 15 13 3 1 10 9 1 10 9 2 16 10 9 4 13 9 1 10 9 1 10 9 2 3 1 9 1 10 9 1 10 9 0 1 9 9 2
48 1 13 10 9 3 0 7 0 1 10 9 1 10 9 2 13 16 1 10 9 4 13 10 9 1 9 1 9 2 10 0 9 1 9 7 15 15 13 3 0 9 1 9 2 7 10 9 2
15 3 10 0 7 0 9 4 13 1 10 9 1 10 9 2
39 3 2 16 15 13 13 2 16 3 4 13 2 3 13 3 1 10 9 7 3 1 10 9 1 10 9 2 4 13 10 9 1 13 10 10 9 3 3 2
44 3 2 1 13 10 10 9 2 1 13 1 13 10 9 1 9 7 13 9 1 9 13 0 13 3 1 9 1 10 0 9 2 10 9 1 9 7 1 9 7 10 9 0 2
48 10 15 2 13 2 13 15 1 10 9 1 10 9 0 2 15 13 10 10 9 1 15 1 10 9 0 2 1 10 9 1 9 15 3 13 3 9 7 9 2 13 9 0 7 13 1 9 2
33 9 9 2 13 10 9 1 13 1 10 10 9 2 9 11 10 0 9 1 15 10 11 4 13 10 9 1 9 1 10 9 12 2
14 4 13 1 9 1 10 0 9 1 10 10 9 0 2
53 7 15 13 1 13 15 3 16 2 16 13 11 1 9 1 10 11 2 10 9 1 10 10 9 2 11 2 4 13 10 10 9 1 10 9 7 1 15 13 10 0 9 1 10 9 11 2 11 1 10 9 0 2
22 4 13 15 16 10 9 0 13 0 1 10 10 9 0 1 10 9 1 10 9 12 2
13 13 1 10 9 11 1 13 1 13 15 10 9 2
15 10 10 9 4 13 0 9 1 10 10 9 1 9 3 2
79 13 16 15 13 1 10 9 0 1 10 9 9 2 1 10 9 13 10 9 7 10 9 1 13 7 13 10 9 0 2 1 13 10 9 3 0 0 1 10 9 1 10 9 1 10 0 9 7 13 10 9 1 10 9 1 10 9 7 1 10 9 0 1 9 16 1 10 9 3 13 3 9 1 4 13 1 9 3 2
68 13 0 13 10 9 7 10 9 1 10 10 9 1 10 9 1 10 0 9 2 2 3 1 10 9 1 10 9 13 1 10 9 1 9 2 1 15 10 11 4 3 13 9 1 9 1 10 11 11 1 15 13 1 10 9 1 10 9 1 0 9 0 2 13 1 10 9 2
28 3 10 9 1 10 0 9 1 9 13 3 0 2 1 3 15 13 15 3 4 13 10 9 1 10 9 0 2
53 3 4 4 13 1 13 0 9 1 9 7 9 2 7 1 13 10 9 7 10 9 1 9 1 10 9 1 10 9 2 1 10 9 1 0 9 7 9 1 10 9 2 3 1 10 9 1 10 0 9 1 9 2
30 10 9 7 10 9 1 10 9 0 3 4 4 13 1 10 0 9 1 10 0 9 1 10 9 7 1 10 9 0 2
31 10 9 1 10 9 0 1 10 9 4 13 0 2 3 1 10 9 1 10 9 0 7 0 0 1 10 9 1 10 9 2
46 1 9 2 10 9 0 4 13 0 2 0 7 0 2 1 13 9 1 10 9 1 10 9 7 1 10 9 1 10 9 7 1 13 1 10 9 10 9 1 10 10 0 9 1 9 2
43 16 13 1 13 10 9 1 9 1 10 9 0 7 3 0 2 1 10 9 13 1 13 15 1 9 3 4 13 0 9 1 9 1 10 9 2 9 9 1 10 9 0 2
15 13 1 10 9 16 13 10 9 1 10 9 0 1 9 2
53 13 16 10 9 0 11 2 1 9 0 0 2 0 7 1 9 2 13 1 9 1 13 0 9 7 1 13 1 10 9 0 7 3 0 1 13 3 10 10 9 7 13 1 10 9 7 1 10 9 1 10 11 2
22 9 9 2 9 9 2 0 9 2 13 1 1 15 13 10 9 11 1 10 0 9 2
7 3 13 3 3 1 9 2
16 1 1 10 9 13 2 10 9 4 13 1 9 1 10 9 2
15 4 4 13 10 9 2 15 4 13 3 1 10 9 0 2
36 10 10 9 13 10 9 1 10 9 1 9 1 10 9 9 7 1 10 9 1 10 9 0 1 9 1 10 9 7 1 10 9 1 10 9 2
14 1 10 9 2 13 3 0 13 10 0 7 0 9 2
28 10 10 9 13 3 0 13 3 1 9 10 9 7 10 9 0 7 13 10 9 1 10 9 0 7 15 0 2
39 15 13 1 10 0 9 1 10 11 11 7 1 10 9 0 1 10 9 9 7 13 16 4 13 10 9 2 15 13 13 10 9 7 10 9 1 10 9 2
17 3 4 4 13 9 15 3 4 13 10 9 0 1 10 9 0 2
17 10 9 4 13 3 0 2 3 0 7 1 9 1 13 9 0 2
24 1 10 9 1 10 9 4 13 0 13 1 10 9 0 0 1 10 9 0 1 10 11 11 2
28 1 15 2 0 9 1 10 9 2 15 4 13 10 0 9 2 7 4 13 16 4 13 10 9 1 0 9 2
14 10 9 13 0 7 13 1 10 9 1 10 10 9 2
79 9 9 2 9 9 2 0 9 2 10 9 15 10 9 13 3 10 9 0 7 0 4 13 1 10 9 1 10 0 9 1 10 9 1 10 10 9 2 9 11 11 2 1 13 1 9 0 2 16 10 9 1 9 0 1 10 9 12 2 12 1 10 9 1 10 9 12 3 1 10 9 13 1 10 9 1 10 9 2
94 13 9 1 15 2 10 10 9 4 13 2 1 10 9 2 16 1 1 10 10 9 10 9 0 1 9 1 10 0 9 4 13 7 13 1 10 9 10 1 10 9 1 10 9 13 3 2 16 13 16 13 10 0 9 1 13 9 1 10 9 3 0 7 3 0 2 13 15 3 1 13 1 13 10 9 0 15 13 10 9 13 1 10 9 0 7 1 13 1 10 11 3 0 2
34 9 9 2 3 4 13 16 10 9 0 7 0 1 10 9 0 7 1 9 2 7 1 10 10 9 2 13 13 10 9 0 7 0 2
21 15 4 13 1 13 1 10 9 1 10 9 9 7 3 1 10 9 1 10 9 2
29 7 15 16 13 10 9 1 10 9 1 10 11 1 10 9 7 3 3 1 10 11 1 10 9 7 1 10 9 2
21 13 16 10 9 13 10 9 0 2 7 3 0 2 1 13 10 9 0 7 0 2
17 16 13 1 9 0 10 9 0 0 1 9 2 4 3 13 15 2
14 10 9 4 3 13 1 10 9 7 1 10 9 0 2
28 4 13 10 9 1 9 15 15 13 1 13 10 9 7 10 9 1 10 9 0 15 13 1 9 0 1 15 2
33 1 10 9 13 3 1 11 2 13 3 16 10 12 9 0 3 0 13 10 9 1 12 9 0 1 15 1 10 12 9 3 0 2
23 15 13 1 10 9 0 2 1 10 9 9 7 1 10 9 1 13 1 9 0 7 0 2
34 13 0 16 10 9 0 3 4 13 10 9 2 7 3 15 4 4 13 2 3 13 10 9 1 10 9 2 1 13 1 10 9 9 2
9 3 13 3 16 10 9 13 3 2
35 13 10 9 0 1 4 13 7 13 3 10 0 9 1 10 9 12 7 10 9 1 9 0 13 1 1 10 9 1 9 1 10 9 9 2
9 10 9 1 10 9 0 4 13 2
38 13 15 1 9 1 10 13 16 10 9 4 13 0 1 10 9 1 10 9 0 1 9 9 1 9 1 10 9 2 13 16 13 10 9 1 10 9 2
20 10 9 3 4 13 16 10 11 11 13 9 1 9 2 3 1 9 2 0 2
18 13 9 16 13 10 9 0 2 16 13 9 2 16 15 13 1 15 2
10 15 13 15 13 3 1 10 9 9 2
43 13 16 13 1 9 2 1 10 9 1 10 10 0 9 1 9 1 9 2 1 10 13 10 9 1 1 10 9 1 9 1 10 9 0 7 0 7 3 3 1 10 9 2
87 9 9 2 13 10 0 9 1 10 9 1 10 9 1 10 9 0 7 1 10 9 1 9 1 10 9 12 2 12 7 10 10 0 9 2 1 15 15 1 15 10 9 0 1 10 9 1 10 9 0 7 1 10 9 1 9 4 3 4 13 2 10 15 13 16 13 13 10 0 9 1 10 9 0 7 10 9 0 1 9 1 10 9 1 10 9 2
26 10 9 9 4 13 1 13 0 9 1 10 9 0 13 1 13 10 9 1 10 9 7 10 9 0 2
60 15 13 1 10 9 1 0 9 16 2 1 15 10 9 0 13 0 2 1 10 10 9 4 3 13 10 9 1 10 9 1 10 9 0 7 10 9 1 10 9 1 9 1 10 9 1 10 9 0 16 3 4 13 10 11 13 3 1 9 2
49 10 9 0 4 13 10 9 9 1 10 9 1 10 9 7 0 7 0 1 10 9 0 2 3 1 10 9 1 10 9 0 2 1 10 9 1 9 1 10 9 0 7 1 10 9 1 9 13 2
117 3 15 13 9 16 10 0 9 11 13 1 10 12 2 10 12 2 10 12 7 10 12 4 13 1 13 10 9 0 1 10 9 0 7 1 10 9 1 10 9 12 10 0 3 13 13 10 9 13 3 7 13 15 0 2 1 9 1 13 16 10 9 0 7 10 9 0 2 10 9 3 0 1 11 2 4 13 1 9 7 1 10 0 9 1 10 9 7 1 10 9 0 2 15 13 1 0 9 7 1 15 10 0 9 1 9 2 9 2 9 7 9 13 3 10 9 2
49 3 2 16 1 13 1 10 9 0 1 9 0 7 1 10 9 1 9 4 4 13 9 0 0 2 3 4 13 16 10 9 0 9 4 13 10 9 0 1 10 13 10 3 0 1 10 10 9 2
62 9 1 10 9 0 4 4 13 10 10 9 1 0 9 2 13 10 10 9 1 10 9 15 13 10 9 7 13 0 9 1 10 9 1 10 9 0 7 1 0 9 2 1 13 15 13 10 9 1 0 9 7 13 9 3 0 1 9 1 10 0 2
39 9 9 2 1 9 15 4 13 10 9 1 9 1 10 9 1 9 1 10 10 9 1 9 1 9 0 2 7 10 9 4 1 13 15 1 9 1 15 2
22 3 13 16 15 15 13 1 13 1 10 0 9 2 7 4 3 13 15 10 10 9 2
40 10 0 9 15 4 13 13 16 4 13 2 16 4 13 10 9 11 7 15 1 9 1 9 1 10 9 0 2 16 10 9 9 4 13 1 10 9 1 9 2
16 3 3 3 4 13 7 10 9 3 13 3 1 10 9 11 2
10 13 10 9 1 9 1 10 0 9 2
12 15 13 13 1 13 3 10 9 1 10 9 2
38 10 0 9 15 13 13 13 16 2 3 2 10 9 0 15 13 3 1 9 2 1 10 9 1 15 3 15 13 1 10 9 15 4 13 1 10 9 2
48 13 10 0 9 1 10 9 9 2 7 1 9 15 13 13 10 9 13 1 10 9 1 10 9 0 2 1 10 9 1 10 9 2 1 9 1 1 10 0 9 2 1 10 9 1 10 9 2
12 13 1 9 0 2 4 13 15 3 1 9 2
23 3 2 3 2 1 9 1 13 13 1 13 10 0 9 13 1 10 9 1 10 9 0 2
19 3 15 4 3 13 10 13 9 2 7 3 13 10 0 9 16 15 13 2
38 15 13 1 10 0 9 2 15 15 13 3 1 16 4 4 13 1 10 9 2 12 9 0 2 9 2 13 0 16 4 3 13 10 9 1 10 9 2
14 1 9 2 10 9 4 3 13 1 9 10 0 9 2
15 3 2 9 9 2 4 3 13 10 9 1 13 10 9 2
23 3 2 10 9 9 4 1 10 9 13 15 9 1 10 10 9 7 13 3 10 10 9 2
26 3 1 10 9 2 13 1 13 16 13 10 9 1 0 9 13 1 9 7 13 10 0 9 1 9 2
35 13 1 10 15 0 16 10 9 4 13 7 16 10 9 4 13 1 10 9 1 10 9 1 9 7 1 10 9 1 10 9 1 10 9 2
29 9 9 2 9 9 2 0 9 2 1 10 9 7 0 1 9 1 10 9 4 1 15 13 15 1 10 9 11 2
29 10 15 15 4 3 13 2 7 15 13 3 1 10 0 9 7 9 15 4 13 1 10 0 9 13 1 10 9 2
19 13 16 10 10 9 4 13 1 10 10 9 10 9 15 10 3 15 13 2
32 15 13 1 10 9 13 1 10 10 9 1 10 9 16 10 9 1 10 0 9 15 4 13 1 13 1 10 9 3 1 9 2
35 10 9 0 1 10 9 0 1 10 9 9 13 3 3 13 1 3 13 15 1 13 16 10 9 4 13 10 9 0 2 7 15 15 13 2
36 15 13 2 3 2 16 10 9 4 1 13 7 13 10 9 0 1 10 9 0 1 10 12 7 3 13 10 0 9 1 9 0 1 10 12 2
6 4 13 12 0 9 2
22 10 0 13 10 9 1 10 9 1 9 1 10 9 0 7 1 10 9 1 9 0 2
18 10 9 3 13 1 13 10 9 16 10 9 7 10 9 0 13 0 2
9 13 3 13 15 10 9 1 9 2
18 16 13 10 9 1 10 9 1 10 9 0 0 1 9 1 10 9 2
20 3 12 9 1 9 15 13 1 10 9 7 1 10 15 15 9 1 13 15 2
27 13 2 1 10 9 1 9 0 1 15 15 4 13 2 15 13 13 10 9 1 10 9 1 10 9 0 2
15 13 0 16 13 1 10 9 9 13 10 9 1 10 9 2
15 3 1 15 3 13 10 9 9 10 11 3 4 13 3 2
29 1 10 9 1 3 10 9 0 7 10 9 15 13 1 4 13 16 3 13 15 1 13 0 9 1 10 9 0 2
12 13 16 4 13 0 1 13 15 0 7 0 2
38 13 16 13 3 0 13 7 13 1 10 9 9 1 13 10 9 1 10 9 0 10 3 15 4 13 1 13 9 1 10 9 13 1 9 0 7 9 2
21 9 9 2 10 9 13 1 10 9 0 7 0 13 10 13 10 9 1 10 9 2
30 1 10 9 1 10 9 0 2 10 9 3 3 0 13 10 13 15 1 10 9 1 10 9 1 10 9 1 10 9 2
26 10 10 9 1 10 11 13 1 13 10 9 0 13 1 13 10 9 1 10 0 1 10 9 1 9 2
19 13 15 13 3 13 10 9 1 9 1 10 9 2 1 3 10 9 0 2
26 16 2 10 9 2 15 4 13 1 13 10 9 0 2 4 13 1 10 9 1 9 0 7 3 0 2
31 10 9 1 9 10 3 13 1 10 9 10 9 15 15 13 2 13 10 9 1 10 9 1 10 9 7 1 10 9 0 2
9 13 1 10 9 15 13 1 9 2
17 9 9 2 3 15 15 4 13 1 10 9 1 10 0 9 13 2
39 1 10 9 2 10 11 1 10 10 9 2 7 10 9 9 1 9 2 4 13 1 10 9 10 10 10 9 7 10 10 9 2 3 3 10 9 0 0 2
53 1 13 15 15 13 9 1 10 9 0 15 2 1 10 1 3 1 10 0 9 2 13 0 9 1 10 10 9 0 7 15 13 1 10 9 1 10 9 1 9 1 10 9 1 10 9 1 9 1 10 9 9 2
48 10 11 2 1 9 2 1 10 0 9 4 13 9 1 10 9 1 10 9 0 2 3 1 9 1 10 0 9 2 1 10 9 0 7 1 10 0 9 1 10 9 0 7 0 1 9 0 2
15 13 3 12 10 9 1 15 4 13 10 9 1 10 9 2
38 1 0 9 2 13 13 1 10 0 10 9 1 9 1 9 7 1 9 1 10 9 1 9 1 10 10 9 0 7 0 2 3 1 13 9 7 9 2
49 1 0 9 2 13 10 0 9 1 9 7 9 1 10 9 0 2 15 3 3 13 3 0 7 0 1 10 9 1 13 10 9 1 10 9 2 9 1 15 15 13 3 10 0 7 0 9 0 2
41 13 2 9 9 2 13 16 13 3 0 16 1 10 9 1 10 9 4 4 13 10 0 9 1 10 9 0 7 3 1 10 9 1 9 1 10 9 0 7 0 2
9 9 0 1 10 9 1 10 9 2
15 9 13 1 10 11 0 1 10 11 11 10 12 9 12 2
7 9 0 1 10 11 11 2
2 9 2
69 13 16 10 9 7 10 9 1 10 9 0 4 13 1 9 1 9 15 13 10 9 1 10 9 2 7 15 10 9 1 10 9 1 15 10 9 0 13 1 10 9 1 9 7 1 9 7 1 10 9 1 10 9 7 1 10 9 4 4 13 1 10 3 0 9 1 10 9 2
40 13 16 13 0 16 10 9 0 4 13 1 9 0 2 16 15 4 13 16 10 9 4 13 1 13 2 1 0 9 2 1 10 9 1 10 9 7 10 9 2
14 13 16 13 0 13 10 9 1 9 0 1 10 9 2
67 13 16 10 9 1 10 11 11 4 13 1 10 9 10 10 9 1 10 9 0 0 2 1 10 9 7 1 10 9 1 10 9 0 2 1 10 9 1 10 9 1 10 9 7 1 10 9 2 7 4 13 1 13 10 9 0 7 10 0 9 1 9 1 10 0 9 2
34 13 16 10 9 9 15 4 13 1 13 2 1 9 1 10 11 11 2 10 9 7 10 9 0 1 10 9 0 7 1 10 9 0 2
25 13 16 10 9 0 1 10 9 7 1 10 9 13 1 10 0 9 1 10 0 9 1 10 9 2
111 10 9 0 13 10 0 9 0 1 10 9 0 1 9 0 1 13 15 1 10 10 9 7 1 10 10 9 2 1 10 9 16 10 9 7 10 9 1 10 9 2 13 3 0 10 9 2 15 13 1 13 2 1 10 9 7 10 9 2 10 9 1 10 9 7 1 10 9 7 1 13 15 2 1 9 0 1 9 0 7 0 2 10 0 7 0 9 7 9 3 1 10 9 1 10 0 9 9 2 1 1 15 1 10 9 13 1 10 10 9 2
3 9 12 2
13 10 10 9 0 13 0 7 0 1 9 7 9 2
21 15 4 13 1 9 7 1 9 7 4 13 10 15 1 10 15 1 9 1 9 2
3 9 12 2
62 1 10 9 13 10 10 9 7 10 10 9 13 1 10 0 9 2 1 9 10 2 1 9 1 9 2 1 9 2 1 9 2 1 9 2 1 9 2 1 9 0 7 1 0 9 2 1 9 0 7 0 2 1 9 2 1 9 7 1 0 9 2
48 10 9 4 3 13 1 10 9 1 10 9 0 2 0 7 0 1 10 9 7 1 10 9 15 10 9 13 2 13 0 2 7 13 1 9 0 7 3 0 2 7 0 1 10 9 1 9 2
3 9 12 2
20 10 9 13 9 1 10 9 2 1 10 9 7 1 10 9 1 10 10 9 2
3 9 12 2
13 10 9 4 4 13 1 9 1 9 7 1 9 2
14 10 9 7 10 9 1 10 9 4 13 1 10 9 2
3 9 12 2
19 10 9 4 4 13 1 9 7 1 9 7 1 9 0 2 0 7 0 2
3 9 12 2
18 10 9 13 9 2 1 10 9 2 1 10 9 1 10 10 9 0 2
3 9 12 2
25 15 13 0 1 1 10 9 7 13 9 2 1 10 9 2 1 10 0 9 1 9 1 10 9 2
23 15 13 9 1 10 0 9 1 10 9 15 13 10 0 9 1 1 10 9 1 10 9 2
3 9 12 2
31 10 9 13 9 1 10 0 9 1 9 1 0 9 1 9 15 13 10 9 0 1 15 13 1 10 9 7 1 10 9 2
3 9 12 2
11 10 9 4 4 3 13 2 13 7 13 2
3 9 12 2
54 10 9 13 9 2 1 9 1 0 9 2 1 10 0 7 0 9 1 1 10 9 0 7 0 2 1 10 9 1 10 9 1 10 10 9 7 1 10 10 9 2 7 1 10 9 1 10 9 0 15 15 4 13 2
3 9 12 2
39 10 9 13 1 10 9 4 13 9 1 1 16 10 10 9 3 4 4 13 3 1 10 0 9 1 10 15 15 4 13 10 10 9 0 1 10 10 9 2
34 10 9 4 13 1 10 9 0 7 0 15 2 1 10 9 1 15 4 4 13 2 3 13 9 1 10 9 0 7 1 10 9 0 2
24 3 4 1 10 9 4 13 10 9 0 1 15 0 1 10 9 1 15 10 9 4 4 13 2
3 9 12 2
42 10 9 4 4 13 1 9 0 1 10 10 9 0 2 1 10 10 9 2 1 10 10 9 2 1 10 10 9 2 7 1 9 1 10 10 9 7 1 10 10 9 2
16 10 9 13 9 1 4 13 1 10 9 1 10 9 7 9 2
3 9 12 2
19 10 9 13 9 1 10 9 1 9 7 1 9 1 10 9 1 10 9 2
3 9 12 2
18 10 9 13 10 9 1 13 7 1 13 1 0 9 9 1 10 9 2
32 10 9 3 4 4 13 16 10 9 4 3 13 1 9 3 0 7 1 9 0 1 10 9 7 1 10 9 1 10 11 11 2
3 9 12 2
17 10 9 4 4 3 13 10 10 9 2 7 10 9 1 13 9 2
3 9 12 2
21 15 13 0 9 1 1 10 9 2 1 10 9 7 1 10 9 1 10 10 9 2
17 10 9 4 4 13 3 1 10 0 7 0 9 1 10 0 9 2
25 10 9 13 10 9 0 7 0 1 10 9 7 13 9 1 4 13 1 10 9 7 1 10 9 2
3 9 12 2
17 10 9 13 10 9 1 13 10 9 10 0 7 1 9 1 15 2
10 10 9 4 4 3 13 10 10 9 2
3 9 12 2
16 10 9 13 9 1 10 9 1 9 2 1 9 7 1 9 2
58 10 9 13 10 9 1 13 1 9 7 1 9 2 7 10 9 1 13 2 3 7 1 9 2 7 7 1 9 7 1 9 2 10 10 9 7 10 10 9 1 10 9 2 1 10 9 2 1 10 9 7 1 10 9 1 10 9 2
3 9 12 2
43 10 9 13 9 1 10 9 1 9 7 1 9 13 10 9 1 3 4 13 1 10 10 9 7 15 1 13 2 13 7 13 9 7 9 1 10 9 7 1 9 1 9 2
3 9 12 2
14 10 9 13 9 1 10 9 1 9 7 1 9 0 2
11 15 4 4 13 1 13 9 1 10 9 2
3 9 12 2
23 10 9 13 9 1 13 1 10 9 1 10 10 9 2 7 3 2 7 1 9 3 13 2
13 10 9 0 13 10 9 1 10 9 1 10 9 2
32 10 9 4 4 13 1 0 7 0 9 2 13 1 9 0 7 0 2 7 1 9 0 2 7 1 10 9 0 1 0 9 2
3 9 12 2
65 10 9 2 1 3 9 1 10 9 2 13 9 1 10 9 0 2 7 1 10 9 1 10 9 0 7 10 9 0 7 1 9 1 10 9 7 10 9 1 10 9 2 1 10 9 0 2 0 7 0 0 1 10 10 9 7 1 10 0 9 1 10 10 9 2
3 9 12 2
31 10 9 13 9 1 10 9 2 1 10 0 9 1 10 9 2 1 0 7 0 9 1 9 7 1 10 9 1 10 9 2
15 10 9 2 1 9 2 13 9 1 0 9 1 0 9 2
20 10 9 13 9 1 13 10 9 7 1 13 15 1 10 9 1 10 10 9 2
3 9 12 2
28 10 9 13 9 1 10 9 7 1 10 9 2 13 1 15 10 0 9 1 10 9 1 9 7 9 0 13 2
3 9 12 2
51 10 9 13 9 1 10 9 1 9 0 1 13 10 9 7 10 9 10 7 1 10 10 9 2 1 0 9 1 10 9 2 1 10 9 2 1 10 9 2 7 1 10 9 0 7 1 10 9 0 0 2
36 7 13 9 1 10 9 1 9 1 9 2 9 2 9 2 9 2 9 7 1 0 9 1 9 1 9 1 9 1 9 0 1 10 10 9 2
13 10 9 7 10 9 13 9 1 0 9 7 9 2
21 10 10 9 2 0 1 10 9 7 1 1 15 2 4 13 1 10 0 9 0 2
3 9 12 2
8 10 9 13 9 1 10 9 2
15 10 9 4 13 0 3 1 15 13 10 9 0 7 0 2
7 10 9 0 4 13 0 2
30 10 9 0 7 0 4 4 13 1 10 9 1 15 7 10 9 0 4 13 3 0 1 15 1 10 9 1 10 9 2
30 10 9 4 4 13 1 10 0 9 1 10 9 0 7 1 10 9 1 10 9 1 10 9 0 7 1 10 9 0 2
38 15 4 13 10 9 2 10 9 2 10 9 1 10 10 9 2 10 9 0 7 0 2 7 4 13 10 9 1 10 11 11 1 10 9 1 10 9 2
21 10 9 13 9 1 9 1 10 9 1 10 9 1 9 1 13 1 10 10 9 2
3 9 12 2
34 10 9 13 9 1 13 9 3 1 10 9 0 1 10 9 2 1 13 1 10 9 7 1 13 1 10 9 0 7 1 10 10 9 2
28 10 9 13 9 1 10 9 1 10 9 0 7 0 13 1 10 9 0 2 0 7 0 1 15 15 13 9 2
3 9 12 2
27 10 9 13 9 1 10 9 0 7 0 1 10 15 10 9 7 10 9 13 1 10 9 4 4 3 13 2
3 9 12 2
25 10 9 13 10 9 1 10 9 2 1 10 15 3 13 0 10 0 7 0 9 1 10 10 9 2
68 1 10 9 1 10 10 9 7 1 10 10 9 2 15 4 4 13 3 1 10 9 15 4 13 1 10 9 1 13 10 9 7 10 9 1 10 9 7 1 10 9 1 10 15 7 1 13 10 0 9 1 10 9 2 1 10 9 0 7 1 10 9 0 1 10 9 0 2
24 10 0 7 10 9 3 4 1 10 9 4 13 1 9 1 10 9 7 9 1 10 11 11 2
3 9 12 2
49 15 1 10 0 9 4 4 13 1 10 9 1 13 10 9 1 10 0 9 2 9 7 9 1 13 10 9 7 1 13 10 9 13 1 10 9 1 15 1 10 9 7 1 10 9 1 15 13 2
6 1 1 13 10 9 2
7 11 13 10 9 1 9 2
8 13 0 16 11 13 1 9 2
19 11 13 10 9 0 7 3 4 13 1 13 10 9 1 10 9 1 9 2
24 13 3 10 9 1 13 9 11 2 15 4 4 13 1 13 9 7 13 9 1 9 7 9 2
12 15 13 10 9 0 13 1 13 15 1 11 2
16 1 4 15 13 1 11 2 4 13 3 12 2 12 2 9 2
15 4 13 10 9 11 0 7 13 10 9 11 1 10 15 2
9 10 9 11 13 3 1 9 0 2
10 15 13 16 10 9 0 3 4 13 2
16 3 2 13 0 13 10 0 9 11 0 1 10 0 9 9 2
22 16 10 9 13 1 10 0 9 2 13 16 1 10 10 9 15 13 10 10 9 0 2
10 1 10 9 13 3 1 15 15 13 2
11 0 9 1 10 10 9 0 1 10 9 2
26 16 4 13 10 9 2 4 13 10 9 9 1 13 10 10 9 1 10 10 10 9 1 10 0 9 2
12 3 13 10 9 1 9 1 11 1 10 9 2
17 13 10 9 16 10 9 1 11 15 4 13 1 13 15 1 11 2
21 11 13 1 10 9 1 13 9 1 10 10 9 13 10 9 9 7 13 10 9 2
24 16 13 2 4 13 10 9 9 1 10 10 9 11 1 13 0 1 3 13 0 9 1 9 2
24 16 3 13 3 10 9 1 11 7 4 13 15 2 4 13 10 9 1 13 10 9 1 9 2
27 16 3 4 3 13 9 1 10 10 9 2 4 13 10 9 1 9 1 10 9 13 1 9 1 10 9 2
13 0 9 1 10 9 10 9 13 9 15 4 13 2
6 9 1 10 0 9 2
12 15 13 10 9 1 13 10 9 7 13 15 2
18 16 3 13 10 9 11 2 4 13 15 1 13 15 15 1 10 9 2
20 16 13 3 10 9 11 2 4 13 10 9 1 10 10 9 1 10 0 9 2
23 13 10 10 9 9 7 10 9 1 10 9 1 10 9 0 1 10 9 7 9 1 13 2
11 15 13 10 9 1 9 0 1 10 9 2
9 3 13 1 13 10 10 9 0 2
29 16 13 10 0 9 2 13 15 16 13 0 3 12 9 7 1 13 10 9 0 1 9 2 9 7 9 1 9 2
25 16 10 9 1 15 13 3 13 3 0 2 13 1 13 9 0 7 0 7 13 10 9 3 0 2
22 10 9 1 15 13 4 2 1 9 2 13 0 1 13 7 0 1 13 1 10 15 2
22 1 13 10 9 2 10 9 1 11 4 13 3 15 1 10 15 1 15 13 1 9 2
13 3 13 1 13 10 9 1 9 1 10 10 9 2
23 13 10 9 1 9 13 10 9 0 1 13 10 10 9 1 10 9 13 10 9 1 15 2
19 4 3 13 10 9 1 9 1 10 10 9 11 1 10 9 9 1 9 2
19 13 1 10 9 11 1 3 1 9 1 10 0 9 11 7 13 9 9 2
13 1 10 9 1 10 9 1 9 2 13 1 9 2
16 13 1 10 9 9 1 9 7 13 10 9 13 1 10 9 2
18 10 9 3 13 0 16 4 3 13 10 9 1 9 1 10 10 9 2
10 9 1 16 13 10 9 1 9 0 2
12 13 10 9 7 10 9 0 1 15 1 13 2
9 3 13 1 15 10 9 1 9 2
15 13 15 16 10 9 13 3 0 1 3 4 4 13 3 2
18 4 13 10 9 0 1 10 10 9 1 10 9 1 10 9 1 9 2
14 13 3 12 9 1 9 15 15 13 7 13 3 11 2
11 13 10 9 7 13 10 10 9 1 9 2
5 13 10 10 9 2
10 13 15 1 3 12 9 1 0 9 2
14 13 10 10 9 1 9 1 9 0 2 9 7 9 2
16 13 10 9 1 9 7 9 0 7 13 15 15 13 10 9 2
11 13 10 10 9 11 7 10 10 9 9 2
17 13 10 10 9 2 15 13 2 1 13 10 9 1 10 10 9 2
9 13 10 9 1 1 10 10 9 2
6 13 1 9 10 9 2
9 13 10 9 0 15 13 3 0 2
8 13 10 10 9 1 10 9 2
22 13 16 13 3 16 10 9 13 2 13 11 2 7 13 2 13 11 2 10 10 9 2
9 13 10 9 0 1 10 9 0 2
13 11 13 1 10 9 10 9 13 1 10 10 9 2
19 4 13 10 9 1 13 15 1 9 0 2 1 15 13 3 10 10 9 2
16 10 9 1 11 4 13 1 9 11 1 13 15 10 9 0 2
25 10 10 9 1 9 0 1 10 12 7 10 12 9 15 4 13 1 11 1 13 0 1 10 9 2
29 1 12 9 2 10 9 13 1 11 11 1 13 1 10 9 0 1 3 12 9 1 11 4 13 1 3 12 9 2
34 10 12 5 1 10 9 1 11 13 1 10 9 9 1 11 11 1 10 9 4 13 0 9 7 4 13 10 10 9 1 13 0 9 2
27 9 1 10 9 1 9 0 7 1 10 9 13 1 9 0 2 10 9 0 13 10 0 9 9 2 9 2
20 1 10 9 1 11 2 13 7 13 1 9 0 10 9 0 13 0 7 0 2
39 9 1 10 9 1 9 0 1 11 13 1 9 1 12 9 0 1 1 10 9 0 2 15 13 1 9 10 9 1 9 9 11 2 11 4 13 0 9 2
48 10 9 13 1 9 0 13 1 10 10 9 0 1 10 9 4 13 11 1 13 10 9 1 10 10 9 1 9 1 10 9 1 10 9 1 10 9 2 9 2 9 1 9 7 9 0 2 2
27 10 9 13 1 10 9 0 1 11 1 11 4 13 1 10 0 3 13 1 10 10 9 13 1 10 9 2
20 9 1 10 9 0 0 1 10 12 5 1 1 10 9 0 1 10 0 9 2
13 9 1 9 0 7 0 0 1 15 1 11 11 2
22 10 9 0 4 4 13 1 10 9 1 12 9 2 1 13 1 10 11 1 12 9 2
11 9 0 1 9 0 1 12 9 1 9 2
14 9 0 1 10 9 1 9 0 1 12 9 1 9 2
13 9 1 10 9 0 1 9 1 9 13 3 11 2
61 16 10 10 9 1 11 13 1 2 1 9 2 1 10 9 1 11 7 9 11 7 9 2 10 10 9 0 4 13 15 1 10 0 7 0 9 2 1 10 9 16 10 9 1 10 9 15 4 3 13 10 9 1 10 10 9 13 10 10 9 2
21 11 4 13 10 9 13 10 11 11 1 13 10 9 1 9 0 1 10 9 13 2
23 10 9 0 0 1 11 13 1 9 10 9 1 9 13 13 1 10 12 7 10 12 5 2
16 10 9 13 9 1 10 9 1 11 4 13 1 10 12 5 2
46 10 9 4 13 10 9 1 10 9 0 2 9 0 1 10 9 1 11 2 13 16 10 9 13 3 13 1 9 9 1 0 9 7 16 10 11 3 4 3 13 1 10 9 1 9 2
9 10 0 9 2 13 10 9 2 2
9 13 3 13 10 9 15 15 13 2
10 4 3 13 10 9 1 10 10 9 2
17 3 4 13 10 9 1 9 2 9 2 9 0 7 10 0 9 2
26 13 1 10 9 2 13 10 9 2 1 10 9 1 15 1 13 10 10 9 0 1 10 10 9 9 2
8 13 9 1 15 13 10 9 2
6 13 10 10 9 9 2
22 13 10 9 2 13 10 9 2 1 13 10 9 1 9 7 15 13 1 10 9 9 2
29 1 10 9 2 4 13 10 9 0 1 10 9 2 13 3 10 9 2 13 10 9 1 10 9 0 7 15 3 2
4 13 15 13 2
10 13 1 15 1 13 10 10 9 0 2
31 13 1 10 15 1 13 10 10 9 2 4 13 13 3 10 10 9 1 11 2 13 10 9 0 3 1 15 15 13 3 2
3 9 0 2
12 1 11 13 1 3 10 9 1 10 10 9 2
17 3 10 9 1 13 10 9 1 10 9 3 13 1 10 10 9 2
16 3 10 9 15 13 10 9 13 10 0 9 1 10 10 9 2
13 3 13 10 9 1 13 10 9 1 10 10 9 2
22 10 9 16 4 13 10 9 2 1 10 10 9 4 13 10 9 2 13 10 9 2 2
18 13 1 1 15 2 10 9 13 10 10 9 0 1 10 10 9 9 2
13 16 13 1 10 9 1 13 15 2 10 9 13 2
11 10 9 4 13 3 10 9 15 13 3 2
12 4 3 13 10 7 10 9 1 9 0 13 2
17 1 0 9 1 10 9 2 13 10 9 2 2 13 10 9 9 2
16 13 10 9 1 10 9 1 10 9 7 10 9 1 10 9 2
19 11 1 11 2 12 9 12 2 12 9 12 2 13 10 9 7 9 0 2
42 10 10 9 13 10 9 1 9 0 7 0 13 3 2 10 9 0 2 2 15 13 10 9 1 10 9 0 1 10 9 0 1 10 9 1 11 11 13 1 10 12 2
34 9 1 10 10 0 9 1 10 9 7 1 10 9 1 9 1 10 9 2 11 4 13 15 1 10 9 1 10 9 1 10 9 0 2
62 10 10 9 13 15 1 10 9 0 1 11 11 2 11 11 2 11 11 2 11 11 11 2 11 1 11 2 11 11 2 11 11 2 11 11 11 2 11 11 2 11 11 2 11 11 2 11 11 7 11 11 2 7 10 9 1 11 11 7 11 11 2
28 15 1 10 9 1 11 4 4 13 7 4 13 10 9 2 7 13 0 9 1 9 1 9 2 9 7 9 2
26 0 9 7 9 0 3 1 9 2 11 13 10 0 9 1 10 9 1 9 1 10 10 9 1 9 2
30 10 10 9 0 15 13 10 9 1 10 9 1 10 10 9 7 13 10 10 9 1 4 9 1 10 9 1 10 9 2
32 16 13 10 9 2 11 13 9 1 10 9 0 2 7 13 10 10 9 1 9 16 4 15 13 1 10 10 9 7 0 9 2
29 3 7 1 10 10 9 1 9 2 13 1 13 10 9 2 10 9 2 10 9 1 9 2 10 9 7 10 9 2
6 13 1 10 10 9 2
19 10 11 11 13 10 9 1 10 10 9 0 7 13 9 1 10 10 9 2
25 11 13 1 9 1 9 1 10 9 1 10 10 9 2 3 1 9 1 10 10 0 9 1 9 2
25 10 9 1 10 10 9 4 3 13 1 9 0 7 0 2 7 13 10 9 1 9 1 9 0 2
13 1 10 12 13 11 11 2 10 9 1 0 9 2
5 13 12 9 3 2
18 11 1 11 4 13 1 10 9 15 15 4 3 13 1 13 10 9 2
29 10 9 2 13 11 11 2 13 15 1 10 12 9 1 10 9 1 10 11 2 10 9 1 10 9 1 10 11 2
29 1 10 12 10 0 11 15 4 13 1 11 1 1 9 3 10 9 1 10 11 2 0 1 13 10 10 9 0 2
16 1 10 12 15 13 9 1 10 9 1 10 9 7 0 9 2
29 4 3 13 10 10 9 1 15 1 10 0 0 9 2 7 13 2 1 10 9 0 2 10 9 0 2 11 2 2
24 1 10 9 1 10 9 2 12 2 12 2 2 4 13 1 11 1 13 10 9 1 10 9 2
22 10 9 1 11 2 0 11 11 11 11 2 13 1 10 9 1 9 1 9 1 11 2
14 10 9 1 10 10 9 13 10 9 0 1 10 9 2
15 1 10 9 1 10 9 15 13 0 2 7 11 11 9 2
11 1 3 9 7 9 0 11 0 11 13 2
8 15 3 4 13 1 10 9 2
36 2 11 2 1 10 9 11 11 1 11 2 15 15 13 10 12 9 2 12 9 1 1 10 9 1 11 2 13 1 9 10 9 1 10 11 2
15 3 10 9 3 4 13 11 2 11 7 13 3 10 9 2
29 10 9 1 11 2 11 7 11 2 4 13 1 10 12 7 1 10 12 2 7 10 9 11 2 11 1 10 12 2
9 1 9 11 4 13 1 10 9 2
15 10 9 0 15 13 10 9 11 7 13 12 9 1 9 2
44 2 16 10 0 9 1 10 9 0 11 2 11 11 11 4 13 10 9 1 10 9 1 13 10 10 9 2 13 10 0 1 10 9 13 3 0 1 10 9 0 7 0 2 2
25 16 10 9 11 13 1 9 2 4 13 1 0 9 1 10 9 2 15 15 13 3 10 0 9 2
26 10 10 9 1 10 12 10 11 1 10 11 13 10 0 9 1 9 11 11 2 13 1 10 10 9 2
23 1 10 9 1 12 9 11 4 13 1 10 9 0 1 9 1 11 2 3 13 12 9 2
33 10 9 2 13 1 13 10 0 0 9 1 10 9 15 15 4 13 10 9 1 9 1 10 9 2 13 3 3 9 1 10 9 2
15 15 15 13 9 1 9 1 10 10 3 0 9 1 9 2
22 1 9 2 4 13 3 1 10 2 9 2 2 10 9 1 9 0 1 10 9 0 2
18 2 16 15 4 13 16 15 13 1 11 2 10 9 1 10 9 13 2
6 2 13 15 11 11 2
17 4 13 10 9 1 13 15 1 10 0 15 1 12 9 2 2 2
20 3 2 10 9 13 1 9 15 13 10 10 9 1 13 10 9 15 15 13 2
32 11 13 10 9 1 10 10 9 2 16 13 10 9 1 10 10 9 7 1 15 1 10 9 1 1 15 2 1 10 11 11 2
23 2 13 13 1 10 9 2 13 15 3 1 9 0 2 1 9 7 9 2 9 7 9 2
19 15 13 1 4 13 10 9 0 1 10 13 10 9 1 9 1 0 9 2
27 2 11 15 13 3 2 1 10 9 1 13 10 9 1 13 10 10 9 1 13 2 10 9 1 9 2 2
9 16 13 1 9 2 10 9 13 2
14 2 3 3 16 10 9 15 13 10 9 15 15 13 2
29 2 11 0 13 10 10 9 1 10 2 9 0 2 2 7 15 13 9 1 10 2 9 2 13 3 1 10 9 2
54 2 1 10 9 2 10 9 4 13 10 9 3 2 10 0 1 13 9 7 9 7 13 15 15 15 4 13 1 10 9 0 1 10 9 2 2 1 15 13 10 10 10 9 1 10 9 1 9 1 13 10 9 2 2
28 1 10 12 10 9 11 15 13 1 11 2 7 11 4 13 1 9 0 7 9 1 10 0 12 9 7 9 2
23 15 13 10 9 0 1 10 10 9 2 1 15 13 1 13 15 1 10 9 1 10 11 2
16 1 10 12 11 13 1 10 11 2 3 13 1 12 9 0 2
16 11 11 2 15 1 9 13 0 9 2 13 9 1 9 0 2
22 11 2 11 11 2 13 1 0 1 10 11 11 2 13 9 1 9 7 1 9 0 2
24 7 2 3 0 1 15 2 10 9 1 9 1 11 11 13 10 10 9 1 13 1 9 0 2
21 16 10 10 9 4 13 2 11 4 13 1 10 9 1 13 10 10 9 1 9 2
19 1 12 9 13 9 7 13 1 10 9 1 11 11 2 10 9 1 9 2
14 1 10 9 11 13 1 13 10 9 1 10 9 0 2
50 1 10 9 10 11 1 10 12 2 13 16 10 9 1 10 9 0 13 2 10 9 13 1 10 9 2 10 0 9 1 10 9 1 9 3 3 0 2 10 9 0 15 15 13 1 10 11 0 2 2
24 1 10 12 11 13 1 11 1 13 10 9 2 7 10 10 9 15 4 13 3 1 10 9 2
27 13 0 1 10 10 13 2 10 9 2 10 9 2 10 0 9 2 15 13 2 13 7 13 1 9 0 2
7 4 13 1 10 10 15 2
24 7 15 13 15 15 13 13 2 10 9 13 1 10 9 2 1 13 10 0 9 3 7 3 2
16 13 0 2 7 3 15 4 13 15 15 13 10 10 9 2 2
9 2 13 10 10 9 1 13 9 2
22 10 9 1 10 9 13 10 0 9 1 10 9 11 2 3 16 11 3 4 3 13 2
75 3 2 1 10 9 1 10 12 15 4 13 1 13 1 10 9 0 2 16 13 1 10 9 0 11 11 2 2 1 10 9 13 1 10 9 3 0 2 1 10 9 1 9 7 10 9 0 15 15 13 1 15 2 2 16 10 9 1 10 9 15 13 1 10 9 1 12 9 2 12 9 2 1 11 2
24 10 0 9 1 11 13 10 9 1 10 9 0 13 10 11 2 13 1 10 11 1 11 11 2
18 13 16 4 13 9 1 13 10 9 2 3 2 15 13 1 0 9 2
14 1 10 12 11 13 10 9 1 12 9 1 9 11 2
19 3 16 13 1 9 1 9 0 2 10 9 15 13 10 9 1 0 9 2
19 16 15 13 2 11 15 13 1 11 7 13 10 0 9 1 10 10 9 2
7 15 3 15 13 3 0 2
14 1 10 0 9 13 2 7 3 13 3 2 12 9 2
6 11 2 11 7 11 2
28 1 10 12 11 13 10 0 11 11 2 15 13 10 9 1 13 9 0 2 15 11 4 3 13 1 10 9 2
32 11 15 13 1 13 9 3 0 2 7 1 10 12 15 4 13 12 9 2 15 13 1 9 7 3 13 1 9 1 0 9 2
43 1 9 2 10 0 9 11 1 11 2 12 2 2 13 1 10 10 9 1 9 3 0 7 2 3 3 0 2 1 10 9 13 2 13 1 2 11 1 11 2 11 2 2
18 10 9 13 0 13 1 13 2 13 1 4 13 3 7 13 10 9 2
15 0 11 2 2 15 13 0 1 9 0 2 0 7 13 2
20 2 11 13 16 11 11 11 13 1 13 15 1 10 13 10 9 0 1 11 2
58 10 9 0 11 11 2 3 2 13 16 2 13 0 13 16 4 13 10 11 11 1 10 9 15 13 1 11 2 15 13 1 9 10 10 9 1 10 10 9 0 1 9 2 7 1 10 9 15 15 13 1 9 1 13 1 0 9 2
16 2 10 9 11 11 13 16 13 10 9 2 11 13 15 0 2
19 1 10 9 11 13 12 9 1 9 1 10 9 7 1 10 9 1 11 2
20 10 0 2 1 10 9 1 10 9 2 13 10 10 0 9 1 10 9 0 2
9 1 10 9 1 10 11 11 13 2
31 2 10 9 2 7 1 9 10 9 2 1 3 0 9 1 10 0 9 1 10 9 2 13 10 3 0 9 1 9 0 2
32 2 1 10 9 1 10 9 12 1 10 12 11 15 13 1 0 9 0 2 10 9 15 10 9 13 1 10 9 1 10 9 2
27 10 10 0 9 13 10 9 0 1 13 1 9 0 1 10 0 9 10 9 0 1 15 10 9 1 11 2
17 10 9 13 3 2 1 15 1 10 9 2 13 1 9 1 9 2
27 2 11 13 0 9 1 10 9 1 10 9 1 11 11 2 11 1 11 2 1 10 15 13 3 10 9 2
28 11 13 1 9 9 1 10 10 9 7 1 10 10 9 7 13 1 13 10 9 0 2 1 9 10 9 0 2
15 10 10 9 7 9 1 9 13 10 10 9 1 10 9 2
24 13 1 9 10 9 1 10 9 2 10 15 15 13 1 10 9 2 7 13 0 1 10 9 2
14 1 9 12 11 13 1 9 1 10 9 1 12 9 2
11 11 3 13 3 10 10 9 1 10 9 2
33 15 13 1 9 1 0 9 16 2 3 9 0 7 13 2 13 1 11 1 10 9 1 13 10 9 1 10 9 0 1 10 9 2
36 16 4 13 10 9 2 1 10 12 11 13 10 9 1 13 10 0 9 1 9 15 4 13 10 9 0 1 2 10 10 9 1 10 9 2 2
7 2 11 1 13 10 9 2
46 2 3 16 3 15 13 11 1 11 2 11 1 11 2 2 1 10 9 4 13 0 1 10 11 11 2 7 1 15 11 13 10 10 9 15 4 13 1 10 10 9 1 10 10 9 2
17 15 4 13 10 9 1 10 9 1 11 7 10 15 3 0 9 2
25 1 10 9 1 10 10 9 0 2 11 13 1 11 7 13 1 10 9 11 1 10 9 1 11 2
24 3 13 9 1 11 11 2 12 2 2 10 9 1 9 13 3 1 10 9 0 1 10 9 2
31 15 13 10 0 9 15 11 13 1 10 10 9 2 7 10 9 15 13 15 15 10 9 13 2 9 1 10 11 9 2 2
36 15 15 13 1 13 15 1 9 0 1 9 2 1 10 9 4 13 1 11 11 2 7 15 13 10 9 1 10 1 3 1 10 10 0 9 2
43 3 3 2 1 10 3 1 10 9 1 10 9 1 10 9 2 11 13 11 11 2 15 13 1 10 9 1 12 9 15 13 10 9 2 11 13 12 9 1 10 9 2 2
12 15 13 10 0 9 13 2 11 1 11 2 2
32 1 10 9 2 13 10 9 0 1 13 15 13 1 10 9 0 2 7 13 10 9 1 13 15 9 2 3 1 9 1 9 2
29 2 10 9 7 9 1 10 9 2 13 3 0 1 10 9 1 9 7 1 10 9 0 2 2 13 1 10 12 2
13 3 10 9 1 10 0 9 1 10 9 13 0 2
15 2 10 9 1 10 9 13 1 10 9 1 10 9 0 2
32 2 1 10 9 15 4 13 10 10 9 1 10 9 1 10 9 0 2 11 13 10 0 9 7 10 9 10 0 9 1 9 2
31 16 10 9 1 9 13 10 9 1 11 0 1 10 12 2 11 15 13 0 2 13 10 9 11 1 11 2 7 1 9 2
41 15 13 16 10 0 9 1 9 2 15 13 10 0 9 0 2 13 0 7 0 1 9 2 7 13 1 10 9 1 10 9 7 10 9 0 15 13 10 9 0 2
29 15 13 2 10 9 0 7 0 15 3 13 7 1 10 9 7 1 10 9 2 7 15 15 13 1 10 12 2 2
32 7 1 9 1 10 9 3 0 1 10 12 2 13 1 9 7 15 13 10 9 2 2 11 13 1 3 13 15 1 10 9 2
51 10 12 13 10 9 1 10 11 1 11 2 10 9 1 9 7 10 9 0 2 2 10 9 1 9 0 15 13 1 10 0 9 1 9 1 9 11 1 11 15 13 10 9 1 9 15 13 9 7 9 2
15 15 13 10 9 2 7 13 10 9 1 13 15 10 9 2
22 1 11 10 9 13 10 0 9 1 10 9 2 10 10 2 9 13 1 13 15 2 2
16 1 10 12 11 13 11 11 2 10 10 0 9 9 1 9 2
30 10 9 1 10 0 9 15 13 10 9 1 10 9 2 15 13 3 10 9 3 13 1 10 9 1 10 10 10 9 2
26 10 9 13 0 2 7 10 9 0 7 0 2 3 15 1 10 9 15 13 10 9 1 10 9 2 2
15 3 10 9 1 11 13 15 1 10 12 9 0 1 11 2
51 10 11 11 2 10 0 9 11 2 12 2 13 10 10 9 0 2 1 15 11 13 1 10 11 1 10 12 10 9 1 11 11 1 13 10 9 1 10 9 0 1 10 9 1 9 1 15 1 10 9 2
68 10 9 1 10 9 1 10 9 13 1 10 9 1 10 0 11 2 3 3 1 9 1 10 10 0 9 0 1 9 2 11 11 2 7 3 10 9 16 2 3 3 2 15 4 13 9 1 10 9 2 11 2 11 2 13 1 10 10 9 13 1 10 15 2 11 11 11 2
21 1 10 12 11 13 10 9 1 10 11 1 11 2 10 9 0 1 9 7 9 2
20 1 10 10 9 15 13 1 13 10 0 9 7 10 9 13 1 10 0 9 2
25 16 13 11 2 2 11 13 0 1 10 9 0 2 0 7 0 2 7 1 9 7 1 9 2 2
19 10 9 13 2 7 1 10 12 13 10 0 9 2 10 2 11 11 2 2
6 15 4 13 12 9 2
36 10 0 9 0 2 7 10 10 9 1 11 2 15 13 10 9 0 1 15 13 10 12 9 1 10 2 11 11 2 2 11 11 2 12 2 2
31 10 9 13 1 11 1 11 2 10 0 9 1 9 1 9 2 15 13 13 1 10 9 1 10 9 3 0 1 10 9 2
18 10 9 1 9 1 11 4 13 1 10 9 0 1 11 1 10 9 2
27 2 11 7 9 1 9 2 2 11 7 9 1 10 9 2 12 2 2 13 10 9 1 10 9 1 11 2
22 15 4 13 1 10 9 11 2 11 2 1 10 9 0 7 0 1 13 10 9 0 2
8 10 9 13 10 0 9 0 2
28 10 0 9 2 1 10 12 2 13 10 9 1 9 1 12 9 2 16 10 0 12 15 13 1 0 12 9 2
22 10 9 0 1 10 9 7 9 13 10 9 13 1 10 9 16 13 10 0 9 9 2
21 10 9 1 11 4 13 1 10 9 1 13 10 9 1 10 12 9 10 9 0 2
18 15 1 10 10 9 1 10 9 4 13 1 9 2 1 15 1 11 2
55 11 11 15 13 1 12 9 1 10 9 0 1 10 9 1 10 9 2 16 10 8 1 8 1 8 2 10 9 1 10 9 1 9 2 12 2 13 1 10 0 9 1 11 2 7 13 3 10 9 0 1 0 12 9 2
9 10 9 1 9 1 11 13 0 2
14 3 13 3 2 7 13 3 1 10 0 9 7 9 2
17 3 15 13 7 13 1 10 9 2 13 1 0 9 1 9 0 2
10 13 3 1 12 9 7 15 1 9 2
22 13 1 4 13 10 9 1 12 9 1 10 0 9 0 1 12 9 1 9 1 15 2
21 11 13 10 10 9 1 9 0 2 13 10 9 1 9 1 9 7 9 1 13 2
24 1 9 13 10 9 1 10 9 1 10 9 2 13 9 0 7 1 15 0 7 1 10 9 2
15 1 9 10 9 0 13 3 10 9 15 1 10 9 0 2
38 16 1 10 9 15 1 10 10 9 3 4 3 13 10 9 0 2 15 1 15 2 1 11 11 2 10 9 2 12 2 2 4 3 13 1 10 9 2
22 13 0 1 11 11 7 11 11 11 1 11 1 11 1 10 11 2 7 13 11 11 2
22 3 2 3 13 3 9 1 10 9 0 7 1 10 9 16 13 15 1 10 10 9 2
24 2 1 10 0 9 13 3 0 2 2 13 11 2 2 3 3 15 4 3 13 1 9 3 2
19 13 16 10 10 9 3 13 1 10 13 10 9 7 1 10 13 15 2 2
43 2 15 3 13 3 10 0 9 1 10 9 1 11 2 1 1 11 2 10 9 1 10 10 9 11 1 11 2 9 1 10 9 7 9 1 10 9 3 0 1 10 15 2
20 15 1 10 9 13 1 11 4 13 1 10 0 9 1 9 1 10 0 9 2
14 3 10 9 13 10 9 13 1 10 9 1 10 9 2
56 1 10 9 1 10 12 11 13 10 9 1 11 2 1 10 9 1 10 9 7 13 3 2 10 11 2 2 2 10 9 2 2 2 15 13 9 1 10 9 7 10 9 1 10 11 1 11 7 10 10 9 0 1 10 9 2
20 13 13 10 9 0 1 10 9 1 11 2 13 16 10 10 9 0 15 13 2
21 3 13 10 9 0 12 9 1 11 7 2 10 9 1 10 10 10 0 9 2 2
3 11 11 2
26 11 4 13 1 10 9 12 9 3 0 1 15 2 11 11 2 10 0 0 9 15 13 3 1 11 2
14 13 10 9 1 9 1 13 10 9 1 10 10 9 2
30 1 11 11 13 10 9 1 10 10 9 7 10 10 9 0 2 1 1 3 10 9 1 10 9 1 10 13 9 0 2
40 11 13 16 13 2 1 10 9 0 1 15 10 9 0 13 3 1 13 15 1 9 0 16 10 9 13 0 1 13 15 13 2 1 9 1 13 10 9 2 2
25 11 11 13 1 10 12 7 10 10 9 7 10 10 9 13 3 10 9 1 13 3 10 10 9 2
28 1 9 1 10 9 0 11 11 2 11 13 1 13 15 1 0 11 1 10 12 7 15 13 13 1 10 9 2
25 1 10 9 1 9 0 2 9 1 9 7 9 1 9 1 10 9 2 10 9 4 3 13 15 2
48 10 12 9 12 2 1 10 9 1 11 1 0 9 2 15 13 1 10 10 9 1 11 2 10 9 1 10 11 2 1 10 9 1 11 2 1 10 9 1 11 2 3 11 2 7 15 13 2
26 10 9 1 12 9 1 13 15 1 10 9 7 13 3 13 10 9 7 1 10 9 7 1 10 9 2
18 10 9 1 15 13 3 0 1 13 2 7 15 13 10 0 9 0 2
16 16 15 4 13 3 2 11 4 3 13 12 9 1 10 9 2
10 9 1 10 9 7 11 1 9 0 2
12 10 9 13 10 9 1 10 9 1 0 9 2
17 11 13 16 2 10 0 3 4 13 1 2 9 2 1 10 9 2
13 2 1 0 9 10 0 2 9 15 13 1 11 2
18 13 1 10 9 0 10 12 9 2 10 9 1 10 0 9 1 15 2
13 11 13 12 9 1 10 10 9 2 10 12 9 2
7 9 11 4 13 1 13 2
28 10 9 4 13 10 9 1 11 11 2 15 3 3 1 10 9 1 11 13 1 13 10 9 7 13 10 9 2
12 11 4 13 1 10 9 1 11 11 1 11 2
23 2 3 2 2 13 11 1 10 9 2 2 4 13 1 0 16 4 13 10 9 1 9 2
9 10 9 13 1 9 1 10 9 2
27 2 1 10 9 13 2 3 10 10 9 1 11 2 2 13 11 11 2 11 11 2 11 9 7 11 9 2
32 1 9 2 11 13 10 9 1 10 9 0 1 10 9 0 11 11 2 15 15 13 1 1 10 9 1 11 11 7 11 11 2
12 11 3 13 11 1 15 1 10 10 0 9 2
33 10 11 11 13 0 1 10 9 1 10 10 0 2 11 13 9 1 13 15 10 0 9 2 15 1 10 15 3 13 3 1 13 2
23 15 13 3 1 10 9 1 9 2 7 10 9 2 13 2 4 3 13 1 10 0 9 2
22 10 9 0 13 10 9 0 1 10 9 2 10 0 9 1 13 15 0 1 10 9 2
43 2 10 9 0 2 2 13 11 2 2 15 4 4 13 1 10 11 11 1 2 11 2 1 9 1 11 2 1 11 7 1 11 4 13 10 9 0 3 1 10 10 9 2
33 2 10 9 0 15 11 13 10 9 2 3 9 1 9 2 1 13 10 9 1 10 10 9 15 13 10 0 9 1 10 9 0 2
18 1 10 9 1 10 0 9 1 2 11 1 10 11 0 2 2 13 2
22 2 10 9 13 3 16 1 3 1 3 13 3 10 9 1 13 10 9 1 10 9 2
17 9 0 1 9 2 9 2 7 9 13 1 13 9 1 10 9 2
21 1 9 2 11 1 11 2 9 1 11 2 13 10 0 9 1 13 9 1 9 2
32 11 15 4 13 1 10 10 9 1 10 11 11 1 10 11 11 2 13 13 10 9 1 9 1 10 9 1 15 15 15 13 2
15 10 9 0 11 11 4 13 11 10 9 1 10 0 9 2
37 11 13 16 16 10 0 13 10 9 1 10 9 0 2 10 9 13 1 10 9 0 2 3 10 9 1 9 15 11 13 1 13 1 10 10 9 2
42 2 1 13 1 10 9 2 2 4 13 1 10 9 1 10 11 1 10 11 2 2 10 9 13 10 9 0 15 13 0 1 13 10 0 9 0 1 10 10 9 2 2
26 2 10 9 1 11 2 2 13 11 2 2 15 13 3 0 16 16 15 4 13 1 10 9 0 2 2
14 2 10 9 4 13 1 10 9 11 11 2 15 13 2
25 2 15 1 10 9 3 0 1 10 10 9 13 10 9 1 11 1 11 2 9 1 11 11 2 2
9 15 13 1 10 10 9 1 9 2
5 15 9 16 13 2
19 10 0 9 2 10 9 2 10 0 9 2 10 0 9 2 15 13 9 2
27 16 11 13 0 1 13 10 9 1 10 9 1 10 9 1 10 9 0 13 9 1 10 9 1 10 9 2
20 10 9 4 13 16 2 15 13 10 9 7 10 9 1 10 9 1 11 2 2
25 10 9 15 11 13 1 9 0 2 15 13 7 13 1 10 9 1 10 11 2 13 10 9 0 2
19 2 16 10 9 13 1 0 2 2 13 11 2 2 3 13 1 10 15 2
23 13 1 10 9 1 10 10 9 15 2 1 10 9 1 9 2 15 4 13 1 13 15 2
40 2 4 13 3 10 0 9 15 10 9 0 11 11 1 9 4 13 2 9 0 2 2 1 10 15 10 9 1 10 9 15 13 3 9 1 10 10 0 9 2
15 10 9 3 0 1 9 13 10 9 1 10 9 1 11 2
28 13 1 10 9 1 10 9 0 7 1 10 9 2 4 13 3 3 1 15 4 13 2 7 3 3 15 13 2
45 10 9 0 13 10 9 1 10 9 0 10 1 11 2 1 10 10 9 2 7 1 10 9 1 10 9 7 9 0 11 11 2 10 15 13 10 9 1 10 9 1 10 9 0 2
38 11 13 3 1 10 9 2 0 7 0 2 1 9 2 7 10 9 1 11 11 1 10 11 1 11 13 10 9 1 10 9 1 10 9 1 0 9 2
45 10 9 1 10 9 2 1 10 9 7 1 10 9 1 9 13 0 1 10 9 1 11 2 3 0 1 13 10 9 0 1 9 1 10 15 10 9 1 10 9 13 10 9 0 2
10 15 15 4 13 10 9 1 9 9 2
18 1 9 10 9 0 1 10 9 15 13 1 10 12 1 10 12 9 2
8 10 9 1 11 13 10 11 2
25 10 9 13 1 10 9 0 2 1 9 1 10 9 1 10 9 7 1 10 9 0 1 10 9 2
3 11 13 2
36 2 16 1 11 15 15 13 1 13 1 10 9 13 1 10 9 3 3 10 9 4 13 2 10 9 0 3 3 13 1 10 10 9 0 2 2
3 11 13 2
24 2 10 9 1 11 13 9 0 7 3 4 13 3 10 9 15 15 13 1 10 10 9 2 2
25 10 10 9 0 13 10 9 0 13 3 3 1 10 9 0 11 11 7 1 10 9 0 11 11 2
20 10 9 1 11 1 2 10 11 11 2 13 10 9 1 10 9 1 11 9 2
16 2 10 9 3 13 16 3 0 2 2 13 10 9 11 11 2
36 10 9 1 10 9 15 13 1 10 9 1 13 9 13 0 1 10 9 0 2 7 13 3 1 10 9 1 11 2 1 1 2 11 11 2 2
24 10 9 0 1 11 15 4 13 1 10 9 1 9 7 9 1 9 7 9 2 7 3 9 2
19 10 11 1 11 2 1 10 0 9 2 13 10 9 0 1 9 7 9 2
29 7 10 9 13 1 10 13 10 10 9 2 7 10 9 1 11 11 13 9 1 15 15 4 4 13 1 10 9 2
26 11 15 13 3 1 10 9 3 0 1 10 9 0 7 1 10 9 0 13 1 10 9 7 0 9 2
31 13 1 10 9 1 10 9 1 10 10 9 3 0 2 13 3 1 9 1 10 9 1 10 9 0 1 13 10 10 9 2
24 13 10 9 1 10 9 10 7 1 10 9 1 1 15 2 1 9 1 11 11 7 11 11 2
7 11 13 10 9 3 0 2
15 1 10 9 2 15 13 10 9 1 10 9 0 11 11 2
24 3 2 10 10 0 9 1 10 9 1 10 9 0 15 13 13 10 9 1 10 0 7 0 2
10 11 13 16 11 13 10 10 9 13 2
28 3 10 9 1 11 11 11 13 0 9 1 10 9 1 11 7 13 11 1 13 10 9 1 11 10 9 0 2
15 11 4 13 10 9 1 10 10 9 7 3 1 15 0 2
17 4 4 13 1 11 11 7 4 4 13 15 1 10 9 1 11 2
22 10 0 11 11 11 13 10 15 2 10 11 0 2 7 10 15 2 10 11 0 2 2
24 10 9 11 11 13 16 2 11 13 10 9 1 10 9 0 1 11 7 10 9 1 11 2 2
9 3 11 11 4 3 13 1 11 2
20 13 10 10 9 1 10 9 7 13 10 10 9 1 9 2 11 10 9 13 2
12 2 10 9 4 13 16 4 4 16 13 2 2
31 16 13 10 9 1 2 9 2 2 11 4 3 13 1 11 10 9 1 10 9 7 10 9 0 7 0 1 10 9 0 2
23 10 9 15 13 1 10 9 1 11 10 9 0 2 15 15 13 1 10 11 11 1 11 2
19 2 15 15 11 4 13 2 2 13 11 2 2 11 4 13 1 13 15 2
14 2 1 10 0 9 11 11 4 13 1 10 9 0 2
22 13 11 7 15 13 3 10 9 2 3 16 13 15 15 13 10 2 9 1 11 2 2
50 10 9 1 11 10 11 1 10 9 2 10 9 1 10 10 9 2 12 2 2 1 15 10 9 0 4 13 1 0 9 0 13 10 0 9 1 10 9 15 11 4 13 1 1 10 9 1 9 0 2
20 3 2 11 13 1 9 16 10 9 0 1 13 11 1 11 13 2 9 2 2
15 3 10 9 3 13 1 11 13 10 9 0 13 11 11 2
42 1 10 12 11 13 1 9 1 10 9 1 9 1 9 1 10 9 1 10 9 1 11 7 15 13 3 1 12 9 2 1 10 12 2 12 2 12 2 7 12 2 2
6 1 10 12 11 13 2
17 2 1 15 0 13 11 2 13 15 1 10 9 7 13 15 3 2
22 2 11 1 9 1 10 9 1 11 1 13 1 10 13 2 10 9 1 12 9 2 2
27 1 10 10 9 11 13 3 10 9 0 1 10 9 7 3 10 9 0 13 1 11 2 10 0 9 0 2
30 2 3 2 10 10 9 13 10 9 1 10 9 0 1 13 10 9 1 10 9 7 10 9 1 9 1 10 9 0 2
36 10 9 1 11 1 10 9 1 15 9 2 9 7 9 0 13 10 0 9 1 9 4 4 13 1 9 1 9 0 7 1 9 7 1 9 2
6 10 0 11 11 13 2
23 2 15 4 13 3 2 1 11 2 1 1 10 10 9 1 9 2 9 7 0 13 3 2
32 1 10 12 11 11 13 11 5 11 2 10 0 9 1 10 9 1 11 1 11 7 10 9 9 1 10 9 1 10 9 0 2
8 11 4 3 13 10 9 0 2
16 15 1 10 10 9 4 4 13 1 9 3 0 7 9 0 2
42 11 11 2 12 9 12 2 13 2 2 12 9 12 2 13 10 9 2 9 7 9 0 2 3 13 1 10 3 0 9 1 9 0 7 10 3 0 9 1 10 9 2
16 4 3 13 10 9 0 9 7 10 2 9 1 10 11 2 2
37 10 10 9 13 2 15 13 10 9 2 13 3 12 9 0 2 12 9 2 12 0 9 0 7 10 0 9 2 1 10 15 15 13 1 9 0 2
27 10 10 9 0 4 4 13 1 10 10 0 9 13 7 4 13 1 9 3 3 1 15 1 10 0 9 2
11 11 13 7 13 1 11 2 9 2 11 2
9 11 2 7 10 0 11 7 11 2
36 1 10 12 7 10 12 2 13 10 9 1 9 1 11 1 9 2 9 2 9 1 10 9 0 13 10 11 11 11 2 3 13 10 11 11 2
27 13 16 2 1 1 10 12 2 1 10 9 1 12 9 2 15 4 13 1 11 3 13 12 9 3 3 2
44 13 10 9 1 10 9 0 1 11 7 15 4 13 10 0 9 1 9 1 10 10 9 0 2 10 10 9 2 10 10 9 0 7 16 10 9 1 15 13 4 13 1 15 2
17 11 13 10 0 9 1 10 10 9 13 1 10 12 7 10 12 2
30 10 10 0 9 0 13 3 9 7 9 2 9 15 13 1 10 9 1 10 9 7 9 1 10 9 1 10 0 9 2
29 3 13 3 9 1 1 10 12 3 1 15 15 11 2 11 7 11 2 13 1 15 1 10 9 0 1 9 0 2
21 1 10 10 0 9 2 13 9 2 13 3 1 2 9 2 7 13 1 0 9 2
20 15 1 10 10 9 0 4 13 1 9 1 0 9 7 9 16 13 1 9 2
45 1 10 12 2 11 11 7 11 11 2 12 9 7 9 9 1 11 2 13 10 11 11 2 10 9 1 9 0 15 13 15 1 12 1 10 9 15 4 3 13 16 13 1 11 2
31 4 13 1 10 9 1 11 11 2 1 10 15 11 4 13 2 3 2 1 2 3 1 10 9 7 1 10 10 9 2 2
29 10 11 2 1 9 2 13 10 9 1 11 2 7 10 11 13 11 1 10 9 15 11 11 11 13 2 9 2 2
25 1 10 0 9 2 10 10 9 4 3 13 7 13 1 10 0 9 1 10 9 7 1 10 9 2
29 10 10 9 0 13 3 3 0 7 4 3 13 2 13 1 9 7 13 1 10 9 0 7 0 1 10 10 9 2
37 11 11 13 9 1 11 11 2 10 9 0 7 9 1 9 13 1 10 11 2 7 1 11 11 2 10 9 1 10 0 9 2 9 1 9 0 2
17 15 13 1 11 2 9 2 11 7 15 4 13 10 12 9 12 2
35 10 9 2 15 4 13 1 10 9 13 1 10 0 9 1 10 9 2 4 4 13 0 1 10 9 2 9 16 11 13 10 12 9 12 2
13 13 10 0 1 12 9 7 10 3 0 1 13 2
49 16 3 13 10 9 1 10 9 2 10 0 9 1 10 9 13 0 1 10 13 16 11 3 13 10 11 11 11 1 11 2 10 9 0 13 1 10 12 2 0 3 10 0 1 9 1 9 10 2
57 1 10 9 0 2 15 13 9 1 9 1 0 9 2 3 10 9 1 10 9 1 9 13 0 2 10 9 1 10 9 13 10 9 0 13 1 10 9 0 2 7 10 9 4 4 13 10 9 0 1 9 0 1 9 0 0 2
23 15 13 16 10 9 1 11 11 2 1 11 2 1 2 11 4 13 10 9 0 1 11 2
16 1 10 9 1 12 9 2 11 15 13 1 10 0 11 11 2
20 10 12 9 12 2 10 9 1 10 9 1 10 9 1 11 13 10 9 0 2
24 10 9 0 2 12 9 1 10 11 13 10 9 15 13 16 10 9 0 4 4 13 10 9 2
57 10 9 3 4 13 3 2 1 10 9 16 10 9 1 11 13 1 13 10 9 1 9 3 10 9 1 9 1 10 0 12 9 2 7 12 9 1 10 9 11 13 1 10 9 10 9 2 11 2 15 4 13 10 12 9 12 2
25 3 12 9 3 13 10 9 1 12 9 2 11 7 10 9 11 2 15 4 13 10 12 9 12 2
19 11 13 1 9 0 1 10 9 1 12 9 7 4 13 10 12 9 12 2
32 1 10 9 1 10 9 2 11 13 10 9 1 10 9 1 1 16 3 4 13 1 9 1 10 9 0 1 11 1 10 12 2
40 10 0 9 13 10 9 1 10 10 9 1 10 2 9 9 2 1 10 9 0 1 9 1 10 9 1 10 11 11 1 11 0 11 11 12 7 12 9 12 2
25 10 9 13 9 1 10 9 1 9 1 10 9 12 7 12 1 1 10 2 9 13 2 1 11 2
14 10 9 13 1 13 9 1 10 9 13 10 9 13 2
46 11 11 2 10 0 9 1 11 2 13 10 9 1 11 1 15 11 13 1 10 9 13 15 1 11 1 13 1 10 9 1 10 9 1 9 1 10 9 1 10 9 0 2 11 11 2
19 15 13 3 13 16 11 15 4 13 1 11 13 10 9 0 1 1 15 2
29 10 0 9 1 10 0 9 13 16 11 4 13 10 10 9 1 9 13 15 1 10 9 1 10 9 0 1 11 2
13 11 11 4 13 16 11 4 13 10 9 1 9 2
40 10 9 1 10 0 9 4 13 16 11 4 4 13 1 9 1 11 11 1 10 11 2 10 9 0 0 15 4 13 10 0 2 11 11 2 1 10 10 9 2
28 10 9 13 10 9 1 1 10 9 13 1 10 10 9 2 7 11 13 10 9 0 1 10 9 1 10 11 2
28 3 3 2 4 3 13 1 11 1 4 13 1 0 1 10 9 11 11 1 10 10 9 11 2 11 1 11 2
41 2 15 13 10 0 9 2 13 1 10 10 9 2 15 1 10 10 9 1 9 0 1 9 1 9 2 13 1 13 0 1 13 0 9 0 1 10 0 1 15 2
29 7 13 10 9 2 11 9 2 2 15 13 1 10 10 9 10 0 9 1 9 2 11 2 9 2 1 10 9 2
56 10 9 13 9 0 1 10 0 9 1 10 9 2 7 15 13 0 16 11 4 13 11 1 13 3 1 3 1 10 13 1 13 15 1 9 1 10 9 0 1 11 11 2 11 11 7 11 0 2 2 10 9 0 2 2 2
60 10 9 1 9 2 9 1 10 9 2 3 2 9 1 9 0 1 9 1 9 2 1 10 0 9 1 10 11 0 1 11 2 1 1 10 9 1 9 1 10 9 2 11 2 9 2 2 9 1 9 2 2 13 11 1 10 9 1 11 2
35 1 10 0 11 11 2 2 10 9 2 2 13 15 9 1 0 9 15 13 1 10 9 1 10 15 2 3 16 13 10 2 9 0 2 2
20 10 9 1 11 13 10 0 9 13 3 1 3 1 1 10 9 0 1 11 2
32 10 9 13 16 10 10 9 4 4 13 1 10 9 1 10 9 1 10 9 12 1 10 9 7 3 3 1 10 9 1 11 2
41 1 10 12 10 9 1 11 4 13 1 9 3 1 10 11 11 11 2 10 9 1 9 1 10 9 1 9 2 0 11 2 15 3 13 10 0 9 0 1 11 2
34 1 10 9 1 10 11 11 1 10 12 2 10 9 13 10 9 0 1 10 0 9 2 11 0 7 13 10 10 9 1 10 11 11 2
13 1 10 12 2 10 9 13 3 10 9 0 11 2
30 1 10 12 13 11 11 2 10 0 9 3 0 1 11 2 7 1 10 12 13 1 10 9 1 10 9 0 1 11 2
16 15 1 10 9 1 11 4 13 1 9 1 15 1 10 12 2
20 1 10 12 10 10 9 4 13 10 9 1 9 7 13 1 13 1 10 9 2
18 1 10 9 1 9 2 11 13 1 13 10 10 9 7 15 1 15 2
36 10 9 1 10 12 1 10 9 1 11 11 15 13 1 10 9 1 10 9 1 10 9 1 0 11 2 12 2 7 11 11 11 2 12 2 2
40 10 9 1 10 10 9 1 10 9 1 10 9 1 10 9 1 11 1 10 12 4 13 1 10 9 1 10 9 16 10 10 9 1 9 13 0 1 10 9 2
56 10 0 9 1 9 1 10 12 2 3 2 13 11 1 10 9 1 15 1 10 2 11 11 1 10 10 9 2 2 15 1 10 15 4 13 1 9 1 10 0 9 1 11 2 3 16 3 4 13 1 9 10 9 4 13 2
21 1 10 12 2 11 11 1 11 13 16 2 10 0 11 2 13 9 2 0 2 2
20 1 10 12 2 11 13 10 9 1 15 11 13 10 9 1 10 9 1 11 2
29 9 0 13 16 13 3 11 1 11 11 11 11 7 10 9 1 11 0 2 16 10 9 13 10 9 1 10 9 2
12 1 10 10 9 11 15 13 1 11 7 11 2
35 1 10 12 2 10 9 3 16 13 1 11 11 11 2 10 10 9 2 11 13 1 10 9 1 11 11 2 11 2 1 9 1 10 11 2
23 15 13 1 10 9 1 11 1 10 12 2 10 9 1 15 10 10 9 13 10 11 11 2
32 11 4 13 10 0 9 1 13 10 9 2 13 1 11 2 15 11 15 4 13 1 11 2 10 9 1 1 10 10 9 2 2
10 1 10 12 13 3 1 9 1 11 2
58 1 10 9 1 10 9 1 10 9 1 10 12 11 11 13 16 2 1 10 9 7 10 9 1 10 11 11 1 10 12 1 9 1 11 11 2 10 11 11 13 3 1 10 9 2 1 10 15 15 13 11 2 11 2 11 2 3 2
46 1 10 9 1 10 12 9 12 1 10 9 13 1 11 1 11 11 2 11 4 13 1 2 0 9 1 9 9 11 2 2 2 10 9 13 15 3 1 10 9 1 11 11 2 2 2
18 3 13 3 0 13 16 10 9 0 15 13 1 11 1 10 10 12 2
44 10 9 0 1 11 4 3 13 1 10 0 9 1 9 2 10 9 1 3 12 9 1 9 1 9 1 10 12 7 9 1 10 12 2 2 15 13 16 3 15 13 9 0 2
12 10 9 1 10 9 3 13 0 1 10 9 2
12 11 13 1 13 11 1 10 9 12 2 12 2
14 1 10 9 12 13 10 9 1 10 0 9 1 11 2
17 7 1 10 9 12 13 10 9 1 1 10 10 9 2 11 11 2
22 1 10 12 2 11 13 10 9 0 2 7 15 1 15 4 13 1 15 1 10 12 2
20 11 13 10 12 9 1 10 12 7 1 15 13 10 9 7 10 10 12 9 2
31 11 4 13 10 9 2 11 11 2 1 10 12 7 11 4 13 11 11 2 10 9 2 12 9 1 1 10 9 1 11 2
13 11 13 10 0 9 7 10 9 10 12 9 12 2
29 10 9 3 10 10 0 9 2 11 11 4 13 0 1 4 13 10 9 0 1 11 11 2 15 13 1 10 9 2
25 11 4 13 1 10 9 0 1 13 0 9 2 13 15 4 13 0 9 7 9 1 10 9 11 2
16 1 9 2 11 13 10 0 9 1 10 10 9 0 2 11 2
27 10 9 1 10 9 13 16 15 4 13 10 9 0 1 10 2 0 9 0 15 10 10 9 4 13 2 2
13 10 11 13 12 9 2 15 13 1 4 13 9 2
36 10 11 13 10 9 2 11 2 15 15 13 12 9 7 13 1 13 1 10 9 10 9 1 10 12 2 13 9 1 10 9 0 0 1 11 2
26 1 10 10 9 2 11 3 13 10 9 2 11 2 15 3 13 3 0 1 10 15 1 10 10 9 2
30 0 9 0 1 9 2 10 9 1 13 15 2 10 0 10 9 0 2 2 10 9 15 4 13 9 1 3 10 9 2
30 10 9 13 10 9 1 10 9 1 11 2 15 3 13 16 10 0 9 0 4 13 15 0 2 7 3 0 1 9 2
28 3 1 1 10 12 2 4 13 10 9 0 1 10 9 1 10 9 9 2 1 10 9 15 15 13 16 13 2
13 10 10 9 0 15 13 1 11 2 11 7 11 2
20 1 10 12 2 3 1 10 9 1 10 11 11 2 4 13 10 9 1 11 2
32 11 4 4 13 1 10 9 7 9 1 9 1 10 9 2 13 10 9 0 1 10 9 1 11 7 10 11 11 1 11 11 2
45 10 0 9 1 10 9 1 10 9 3 13 10 15 1 10 15 1 10 9 2 7 10 9 13 1 10 9 16 11 13 10 15 2 3 1 10 9 7 1 10 13 10 10 9 2
33 10 9 2 1 11 11 7 10 0 9 0 2 13 0 2 16 0 12 0 9 7 10 9 4 13 11 13 15 3 13 9 0 2
21 9 0 13 3 10 9 16 10 9 13 9 1 9 1 0 9 1 10 9 0 2
35 10 0 9 13 1 11 13 11 0 7 10 12 9 1 11 0 2 13 1 10 0 9 12 1 10 12 2 1 10 9 1 10 9 0 2
45 3 2 10 9 1 11 13 0 1 13 7 10 9 1 10 9 13 16 11 11 2 10 9 1 10 9 2 10 0 13 7 10 12 9 1 11 4 3 13 1 10 10 0 9 2
56 10 10 0 9 0 2 15 15 13 3 1 10 9 1 10 12 1 10 11 1 11 2 11 7 11 1 11 11 2 13 10 9 0 1 10 9 0 7 0 7 4 4 13 1 10 9 1 10 9 1 10 9 1 10 11 2
35 10 0 9 4 13 1 10 9 1 0 9 0 2 3 11 11 7 11 11 2 1 10 9 1 10 9 0 2 7 1 10 9 1 11 2
43 10 9 1 10 9 4 3 13 1 9 0 2 7 3 4 4 13 10 9 1 10 11 13 2 16 4 13 1 10 0 7 0 9 7 3 4 13 9 1 10 9 0 2
48 1 0 12 9 1 11 2 1 15 12 9 13 13 10 9 2 10 9 1 10 11 7 1 10 9 1 10 9 1 13 10 9 0 1 10 9 1 9 13 1 9 10 9 7 10 9 0 2
45 10 0 9 0 1 11 7 15 1 9 0 2 15 13 0 0 9 7 0 9 0 2 13 9 1 10 9 1 10 9 12 1 10 12 1 10 9 0 1 10 10 9 3 0 2
24 9 1 10 9 1 11 11 13 10 0 9 1 9 0 2 9 0 7 0 9 1 9 0 2
43 10 0 9 1 11 2 10 3 0 10 9 1 11 2 13 10 9 1 10 0 9 0 11 2 15 13 10 9 1 9 0 7 4 13 0 1 10 9 1 10 9 0 2
40 10 9 7 10 9 1 9 1 10 9 1 15 2 10 13 9 0 1 16 15 13 2 7 10 0 9 1 10 0 9 13 10 9 1 10 0 9 1 11 2
42 1 10 0 11 0 2 13 3 3 1 9 2 11 13 10 9 1 9 1 10 9 1 10 0 9 12 1 10 12 2 11 0 2 9 0 7 0 2 7 11 0 2
40 10 10 9 13 3 0 7 0 9 9 16 13 3 1 10 9 0 1 10 9 2 1 10 9 1 10 9 2 7 13 10 9 0 1 10 15 3 0 9 2
9 10 9 13 7 13 1 12 9 2
23 11 7 11 2 10 0 9 0 1 10 0 9 0 2 1 10 9 2 7 1 10 9 2
30 7 11 11 2 13 1 10 9 13 1 10 12 1 11 11 11 1 11 11 1 11 2 15 13 10 0 9 1 9 2
44 1 11 11 0 1 11 2 1 10 11 11 2 10 0 9 1 9 2 9 2 9 2 9 0 2 3 10 0 9 1 11 1 10 9 2 13 1 13 15 10 15 10 15 2
41 1 10 9 1 10 0 9 2 11 13 10 0 2 9 0 2 9 1 11 2 11 7 11 2 7 15 13 3 15 15 13 3 7 10 1 10 10 3 0 9 2
17 10 9 13 16 10 0 9 1 11 13 10 9 1 10 10 9 2
38 10 9 1 10 9 1 15 1 10 9 3 0 1 11 2 11 2 4 4 3 13 15 1 10 0 9 0 2 3 1 10 10 0 9 15 13 1 2
35 1 9 1 10 0 11 2 10 10 0 9 13 10 9 2 1 10 9 1 10 9 0 2 11 7 11 2 0 13 10 9 0 1 9 2
31 10 9 1 10 9 1 11 15 13 3 1 9 0 7 9 1 10 9 15 13 10 9 7 13 10 9 7 10 10 9 2
27 1 10 11 10 9 11 13 10 9 0 1 11 1 10 9 1 13 15 1 13 10 9 0 15 15 13 2
52 1 10 11 11 10 0 9 13 10 0 9 1 13 1 10 10 9 13 9 1 10 9 1 9 15 13 1 10 9 7 1 10 9 1 10 9 1 11 7 1 10 9 1 11 2 10 9 3 0 1 11 2
27 1 10 9 11 11 2 2 10 9 3 13 7 1 10 9 0 7 1 10 9 9 1 10 10 9 2 2
54 1 10 11 2 10 3 0 7 10 3 0 1 10 9 1 11 2 10 9 0 13 11 7 10 9 2 11 11 2 1 13 10 9 0 7 1 13 10 9 1 1 16 3 4 13 1 10 9 1 10 9 1 9 2
13 1 10 9 11 13 1 10 9 0 10 9 0 2
38 10 10 0 9 3 0 2 11 7 11 7 11 2 13 1 10 9 3 0 1 11 7 4 13 10 10 9 0 13 1 10 9 7 9 11 11 11 2
19 1 10 9 0 2 11 13 9 7 9 7 13 1 9 0 12 9 0 2
24 11 2 10 9 1 9 7 10 9 2 3 1 11 2 9 1 11 2 9 9 1 10 9 2
34 3 0 1 10 9 2 10 12 9 13 10 9 3 0 1 10 9 1 10 9 12 7 13 1 9 7 1 10 9 1 9 3 0 2
40 10 9 4 13 10 9 1 9 1 10 9 1 10 9 1 10 9 3 0 1 9 1 11 2 7 4 3 3 13 10 0 9 1 10 9 0 1 10 9 2
14 3 13 0 1 10 9 0 11 13 10 10 0 9 2
25 10 9 1 10 9 1 10 12 1 10 11 11 13 16 10 9 4 4 13 1 12 9 0 0 2
42 1 9 1 10 9 1 9 1 10 12 2 12 2 10 9 1 11 4 13 1 10 10 9 1 10 10 11 7 1 10 11 11 1 10 11 2 1 9 1 10 11 2
43 10 9 15 15 13 1 9 1 13 10 0 9 1 10 11 0 2 13 1 11 11 2 2 16 13 11 2 11 2 11 7 10 9 2 7 15 13 1 9 10 9 2 2
49 16 10 9 0 15 13 13 1 10 9 1 10 9 2 13 10 11 7 13 10 9 1 13 10 11 11 2 10 0 9 1 9 13 1 9 1 9 2 1 10 9 9 1 10 11 2 1 11 2
24 10 11 13 1 10 9 1 10 12 2 1 10 11 11 2 15 1 10 0 9 1 4 13 2
29 10 0 9 1 10 3 0 9 1 11 0 1 10 12 2 0 11 2 11 7 11 11 2 4 13 1 10 11 2
26 1 10 12 2 4 13 9 1 11 11 11 1 11 11 2 10 9 13 10 9 0 1 11 11 0 2
40 1 10 9 1 10 9 13 0 2 10 11 11 13 1 0 12 9 1 11 1 10 12 9 12 7 10 12 9 12 2 1 15 12 9 1 10 9 1 11 2
20 1 10 12 2 1 9 15 13 1 10 9 0 11 7 1 9 1 10 11 2
26 10 9 0 2 13 1 10 9 1 10 0 9 0 2 13 1 11 1 13 0 7 3 0 9 0 2
24 1 10 9 1 11 13 9 9 1 10 9 1 11 11 2 11 11 2 11 11 7 11 11 2
27 11 13 1 10 9 1 9 1 10 0 9 1 10 9 0 2 1 10 15 11 0 2 11 7 11 11 2
30 10 0 9 0 11 11 13 2 1 10 15 2 10 9 1 10 9 11 1 11 7 11 7 11 1 10 11 1 15 2
33 4 13 1 11 11 1 9 1 10 0 9 2 15 13 1 9 1 15 1 11 1 1 15 13 7 15 1 10 0 1 11 11 2
35 3 2 10 12 9 10 9 13 10 9 1 10 11 2 13 15 3 2 10 9 15 13 1 0 9 10 9 1 9 1 10 9 1 11 2
37 1 10 12 11 11 7 11 11 2 12 1 10 9 1 11 15 13 9 1 10 11 11 2 13 10 11 11 2 10 9 0 1 10 9 1 11 2
31 15 1 10 9 4 3 4 13 1 10 10 9 1 15 2 9 0 1 9 1 9 13 1 12 1 9 1 13 12 9 2
27 3 15 13 9 15 13 10 9 1 11 1 10 9 2 13 1 10 11 11 1 2 9 13 7 0 2 2
30 11 11 13 15 1 15 2 9 9 2 13 16 13 9 13 2 13 7 13 7 2 1 10 9 2 4 13 1 9 2
14 16 10 9 1 10 9 13 2 15 13 1 1 15 2
35 10 9 4 13 1 9 1 9 7 1 9 2 1 10 9 1 10 9 7 1 10 9 1 10 9 2 7 3 1 10 0 9 1 11 2
33 1 10 9 2 1 1 9 11 2 11 2 11 7 11 2 11 4 4 13 10 9 1 10 9 1 10 9 1 15 7 1 9 2
67 1 10 9 1 10 11 11 2 3 2 16 15 1 10 9 3 0 13 1 1 15 9 2 10 9 1 9 1 10 12 13 3 15 1 15 1 15 1 10 12 16 10 10 9 4 4 13 1 10 9 11 11 2 13 16 3 15 15 4 13 10 0 9 1 13 9 2
37 1 10 9 12 7 12 2 16 10 9 13 13 1 9 1 10 9 2 11 13 12 9 0 1 10 9 0 2 11 7 11 7 10 9 1 11 2
17 1 10 9 11 7 11 2 10 0 11 13 10 9 0 1 11 2
20 16 1 10 9 1 11 2 10 9 2 9 0 2 4 13 1 10 0 11 2
28 13 15 1 10 9 1 11 2 10 9 13 10 9 1 10 9 7 1 10 9 0 15 13 1 10 9 0 2
14 15 13 0 7 4 13 10 9 1 10 9 1 11 2
38 10 0 9 0 2 10 9 1 10 9 2 1 15 10 0 9 4 13 16 13 1 10 9 0 2 4 13 1 10 0 9 1 10 9 1 10 12 2
18 10 9 3 13 0 1 10 13 16 11 4 13 10 9 1 10 9 2
15 10 9 13 16 10 10 0 9 4 13 1 9 3 0 2
37 1 10 9 7 10 9 2 13 1 11 11 2 1 11 11 1 10 12 2 15 13 10 9 1 10 0 9 7 1 10 10 0 2 10 0 9 2
30 1 10 12 2 12 9 0 1 10 9 12 7 12 13 1 10 9 0 2 13 1 9 1 11 7 1 10 10 9 2
21 13 1 10 12 2 10 9 13 10 0 1 10 9 3 0 1 11 1 4 13 2
38 10 9 3 13 0 1 10 9 1 9 1 15 1 10 12 9 2 7 13 0 13 16 11 15 4 13 1 10 9 1 10 10 9 2 1 9 0 2
39 3 1 1 10 9 3 13 1 10 12 9 1 10 9 0 1 10 12 2 11 11 4 13 9 1 10 12 1 10 2 0 9 1 10 10 9 0 2 2
20 10 9 13 16 1 10 9 13 4 13 10 9 1 10 9 15 11 13 13 2
9 13 16 13 1 9 12 9 13 2
39 15 1 10 0 9 1 10 9 13 1 10 9 0 2 10 2 0 9 2 2 2 7 15 1 10 9 0 1 10 0 9 2 10 2 0 9 2 2 2
45 3 13 0 16 10 9 13 9 0 2 7 16 10 2 15 2 1 10 9 15 15 13 15 13 10 0 11 2 3 16 11 13 16 1 10 11 11 4 2 13 10 10 9 2 2
23 10 9 1 10 12 4 13 1 2 9 11 2 2 13 2 10 0 9 2 1 10 9 2
25 10 9 13 10 11 1 10 0 9 1 10 9 1 10 9 2 9 0 2 9 2 9 7 9 2
16 10 0 9 0 1 11 4 13 1 10 9 0 1 10 9 2
24 15 13 1 10 9 0 15 3 3 13 1 9 0 1 10 9 1 10 9 7 1 10 9 2
30 10 9 15 13 1 9 7 9 0 7 3 13 7 10 9 13 3 0 2 13 1 4 13 3 1 13 1 10 9 2
18 1 9 10 0 9 1 11 11 2 1 10 9 2 3 13 10 9 2
14 7 10 9 1 10 12 9 1 11 4 4 13 9 2
16 3 3 3 2 11 13 1 13 10 9 0 1 10 10 9 2
21 10 9 0 1 11 0 13 10 10 9 1 10 9 1 9 1 10 9 0 0 2
26 1 10 0 9 2 10 0 9 1 15 1 11 13 10 9 1 10 9 1 10 9 3 0 1 11 2
19 3 13 10 9 1 9 15 13 10 9 1 10 9 0 1 15 3 0 2
23 11 15 13 1 10 10 10 9 2 11 7 11 13 3 10 9 0 1 10 9 1 9 2
41 1 10 9 1 10 9 12 1 10 12 2 1 10 9 1 11 7 11 2 11 0 7 9 1 10 9 1 0 9 2 11 4 3 13 1 13 1 9 3 0 2
18 13 3 3 10 10 9 7 10 10 9 1 10 9 1 10 9 0 2
17 10 9 0 10 1 11 13 10 9 0 2 13 1 10 9 0 2
23 1 9 2 15 13 1 10 9 0 2 3 1 9 2 13 1 10 9 1 10 9 0 2
20 10 9 0 1 10 10 0 9 0 13 3 15 1 15 1 10 10 0 9 2
30 1 10 10 9 2 10 10 9 13 1 13 2 13 15 7 13 1 10 9 1 10 9 2 1 10 9 1 13 0 2
19 10 9 13 9 1 10 9 0 2 11 13 1 13 7 13 10 10 9 2
18 10 9 13 0 9 7 9 1 10 9 1 9 1 11 11 7 11 2
17 11 15 13 2 1 9 2 1 13 10 9 1 10 9 1 11 2
35 10 9 0 11 11 4 13 10 10 9 1 2 3 9 2 9 2 0 2 7 2 1 10 9 2 3 0 2 3 3 13 7 0 2 2
19 1 10 0 9 1 10 10 9 2 11 4 13 10 9 1 13 10 9 2
23 15 13 9 2 9 7 9 0 2 7 9 0 1 10 9 7 1 10 9 1 10 9 2
21 1 11 2 1 9 2 10 9 13 1 10 9 7 9 3 13 2 1 10 15 2
9 10 9 4 13 1 13 10 9 2
61 10 0 9 2 1 10 10 9 0 7 10 0 9 1 10 9 2 4 13 10 0 9 0 2 1 15 9 0 7 0 4 13 10 15 1 10 15 2 10 9 4 13 2 9 7 9 4 13 2 7 10 9 4 13 2 13 10 9 1 9 2
13 11 13 10 9 0 1 10 0 9 1 10 9 2
20 1 10 10 9 1 10 9 2 13 1 10 9 9 1 9 1 11 7 11 2
24 13 10 9 1 13 10 9 1 9 2 7 1 13 1 10 9 10 3 9 0 1 10 9 2
33 10 9 1 9 13 16 10 9 1 11 4 13 1 10 9 2 1 10 9 7 1 0 9 1 10 9 1 10 9 1 10 9 2
26 1 10 13 10 10 9 2 11 4 13 1 10 10 9 9 3 0 7 0 2 7 9 1 9 0 2
18 1 10 9 2 4 13 9 1 10 10 9 0 1 10 0 9 0 2
17 10 9 1 11 4 13 10 9 0 1 10 9 7 10 9 0 2
17 1 9 2 4 13 10 9 0 1 9 2 9 2 9 7 9 2
23 1 1 11 7 11 2 1 9 2 10 9 1 9 3 4 13 1 9 0 1 10 9 2
14 10 9 4 13 3 1 13 9 1 1 9 7 9 2
12 7 11 15 13 1 13 10 9 1 10 9 2
10 10 10 9 4 3 13 10 9 0 2
20 10 9 0 4 13 1 13 13 10 9 1 10 9 0 2 7 1 10 9 2
25 10 9 11 11 4 13 10 10 9 1 9 1 11 1 11 1 2 0 9 1 10 9 0 2 2
14 11 13 9 1 11 11 2 11 11 2 7 11 11 2
13 10 9 1 10 9 0 11 11 13 15 1 11 2
19 10 10 11 11 1 11 2 11 13 10 0 9 0 2 0 1 11 11 2
15 10 9 4 13 12 9 1 9 13 1 10 9 1 11 2
14 11 4 3 13 10 9 2 13 10 0 7 10 11 2
19 10 9 0 0 11 11 2 9 1 11 11 2 4 3 13 11 1 9 2
28 10 9 11 11 15 4 13 1 10 9 0 2 1 9 1 15 1 11 2 1 10 10 9 1 10 9 0 2
28 11 11 15 4 13 3 3 1 10 0 9 1 10 10 11 1 10 0 9 2 10 0 9 0 1 10 9 2
33 9 1 2 1 10 9 13 2 2 11 1 11 2 7 2 9 0 2 2 11 2 4 13 9 1 10 9 0 1 10 10 9 2
16 11 3 4 4 13 16 13 1 9 2 7 4 13 10 9 2
34 1 10 12 2 10 9 7 9 11 11 15 4 13 1 2 10 3 9 2 1 10 9 1 9 0 7 1 10 9 7 1 10 9 2
27 10 9 1 10 9 0 1 10 11 1 10 11 11 11 1 11 15 4 13 1 1 11 2 11 7 11 2
45 1 10 11 11 2 11 11 13 1 11 1 2 11 1 10 9 2 9 2 9 2 7 9 1 10 10 9 2 2 3 16 4 13 1 10 0 9 15 2 11 13 10 9 2 2
24 1 10 9 1 10 9 1 10 12 7 10 9 1 10 0 9 2 13 1 9 10 9 0 2
22 1 9 2 10 9 1 10 9 13 3 11 1 10 1 3 1 11 11 7 11 11 2
16 11 11 2 1 9 2 13 11 1 10 9 1 0 7 0 2
28 3 2 10 9 7 9 11 11 13 10 0 9 1 11 2 13 1 11 2 2 15 13 2 7 13 11 2 2
10 1 0 9 2 10 9 1 11 13 2
28 7 1 10 0 9 2 10 9 13 1 13 1 11 1 10 10 9 7 1 13 15 15 13 10 10 9 0 2
34 10 9 1 9 0 1 10 10 9 2 3 15 1 11 11 1 10 12 7 11 11 1 10 12 2 13 1 13 1 10 10 0 9 2
12 1 10 12 2 4 4 3 13 1 9 0 2
16 1 15 15 15 13 15 13 11 2 11 2 11 7 11 11 2
19 1 10 9 1 10 9 2 11 4 13 1 10 9 7 9 0 11 11 2
18 7 10 9 11 11 11 13 10 10 9 1 10 9 1 10 9 0 2
19 1 10 0 9 2 10 9 0 1 10 9 1 11 3 13 1 10 9 2
49 2 10 9 1 10 11 2 2 10 9 11 11 13 1 10 12 2 2 15 3 13 2 1 10 9 13 2 1 15 15 2 1 10 3 0 2 10 3 0 2 7 10 3 0 1 10 9 0 2
2 0 2
16 2 10 9 13 10 10 9 1 10 9 0 2 1 0 9 2
25 10 9 7 9 11 11 11 15 13 9 1 10 9 1 10 9 1 11 2 13 15 2 9 2 2
14 13 16 10 0 9 1 10 9 1 11 13 11 0 2
30 10 9 0 1 10 9 1 10 0 9 2 3 0 1 10 13 11 2 13 3 10 10 9 1 10 9 1 10 9 2
17 10 9 1 11 7 10 9 1 11 13 10 9 1 10 10 9 2
17 10 9 7 9 0 11 11 13 10 9 0 1 10 9 1 11 2
24 10 9 7 9 11 11 11 13 1 11 16 10 2 9 2 1 11 1 9 15 13 3 0 2
30 11 2 1 1 11 11 11 7 10 9 1 10 11 11 2 13 1 10 9 1 10 9 3 0 1 10 9 1 11 2
35 1 10 9 12 2 10 9 1 11 15 13 1 0 9 1 10 9 2 10 9 2 10 0 9 2 9 0 2 0 2 7 0 9 0 2
25 3 12 9 1 10 9 1 11 2 10 9 1 10 9 1 10 9 1 15 13 2 13 1 13 2
19 9 0 13 13 11 11 2 11 11 7 11 11 11 2 0 9 1 11 2
11 10 2 9 1 9 2 4 4 3 13 2
21 10 9 13 16 10 9 1 10 9 1 11 13 9 16 10 13 0 4 13 0 2
17 10 9 1 11 2 11 11 2 13 3 1 10 9 0 3 0 2
36 10 9 3 13 4 13 10 9 1 9 0 13 1 11 11 2 13 1 10 12 1 10 9 1 10 9 1 10 10 9 1 9 1 11 11 2
21 3 2 3 2 10 9 4 4 13 7 10 9 3 13 1 9 1 10 10 9 2
30 1 10 12 10 9 13 16 11 11 3 13 1 9 2 1 9 1 10 9 1 9 2 2 10 9 0 1 10 9 2
31 1 10 12 10 9 1 10 9 1 11 2 11 2 9 1 10 9 1 15 15 3 13 10 9 1 10 9 0 1 11 2
30 10 9 13 9 1 10 10 9 2 7 1 9 7 1 2 1 10 9 1 10 10 9 2 7 10 9 3 13 0 2
11 10 9 1 10 9 0 1 11 4 13 2
18 11 2 10 0 1 10 12 9 2 13 12 9 3 10 12 9 12 2
25 1 10 9 10 9 4 13 16 10 9 1 11 13 0 2 13 15 1 10 9 1 10 10 9 2
20 15 13 10 0 9 1 10 9 1 10 0 9 2 3 7 1 10 9 0 2
24 10 12 9 2 13 2 11 11 2 2 4 13 1 10 9 13 7 13 1 9 1 9 0 2
51 10 9 0 13 10 9 0 1 11 7 3 15 13 9 1 15 4 3 13 10 10 9 2 7 2 10 9 1 11 15 11 11 13 0 2 7 10 10 9 1 11 13 10 0 9 1 10 10 9 0 2
27 1 10 0 9 2 10 9 1 4 9 0 1 11 13 10 9 1 9 1 9 1 0 9 15 13 11 2
23 10 9 13 3 1 10 9 1 0 9 2 9 0 2 9 7 9 1 9 1 0 9 2
32 10 9 1 11 13 12 9 0 2 13 1 10 11 11 1 10 12 2 13 13 10 9 1 10 11 1 9 2 9 7 9 2
46 12 9 15 3 4 13 1 10 11 11 2 10 12 0 9 7 11 2 9 1 11 2 4 3 13 1 9 13 1 10 9 1 9 2 13 16 11 13 10 9 0 1 10 10 9 2
14 10 9 1 11 4 13 1 10 9 2 11 11 2 2
10 4 13 10 9 3 0 2 10 9 2
15 7 4 13 10 9 3 0 2 10 9 1 10 9 0 2
13 7 13 3 10 12 9 4 13 10 9 3 0 2
36 7 15 15 4 13 1 13 13 16 2 3 1 10 9 2 13 9 0 15 2 15 13 2 16 13 1 13 2 15 13 1 13 0 9 3 2
20 7 10 0 9 3 13 10 9 1 10 9 2 7 9 15 15 15 13 3 2
6 7 4 13 1 15 2
6 15 13 15 2 0 2
5 15 4 13 15 2
18 7 16 13 10 9 7 13 1 3 2 3 4 13 1 10 9 0 2
3 15 13 2
6 9 0 2 15 0 2
9 13 15 10 9 1 10 10 9 2
14 7 15 4 13 10 9 3 0 1 10 7 10 9 2
11 15 13 10 9 1 11 11 1 10 12 2
18 11 11 2 1 10 9 2 13 10 3 0 9 0 1 10 9 9 2
15 15 13 0 9 1 9 0 1 10 9 7 1 10 9 2
23 11 11 2 10 9 1 10 11 11 11 2 1 10 15 15 13 2 1 10 9 12 13 2
29 2 10 9 1 10 9 15 13 1 10 9 1 10 9 13 3 0 1 13 13 0 10 9 1 9 1 9 2 2
20 15 15 13 1 10 9 4 1 0 9 13 10 0 9 1 9 1 10 9 2
9 7 13 1 10 9 15 15 13 2
2 13 2
8 2 11 10 9 4 13 2 2
8 2 10 9 1 10 9 2 2
8 1 10 9 10 9 13 9 2
22 7 10 9 13 10 9 7 15 13 1 10 9 7 1 10 9 16 13 9 1 9 2
7 15 4 13 10 9 0 2
12 13 10 9 3 0 2 7 15 4 13 13 2
28 10 9 1 10 9 1 10 9 7 15 1 10 9 0 2 1 9 15 13 1 10 9 1 0 9 1 13 2
6 7 4 13 15 15 2
12 2 13 10 9 2 13 3 1 10 9 2 2
7 10 9 1 10 9 0 2
32 16 10 9 13 10 9 2 4 13 15 2 15 15 13 1 9 3 0 2 7 13 9 0 1 15 15 13 10 9 1 9 2
16 16 16 10 9 13 10 9 2 15 13 1 13 10 10 9 2
41 13 10 9 1 10 9 0 2 10 9 2 10 9 0 2 7 13 16 10 9 13 10 9 1 10 9 1 10 9 1 10 9 2 7 3 3 2 13 10 9 2
26 7 15 13 1 9 2 1 10 9 1 1 10 9 1 10 9 2 13 10 9 0 15 10 9 13 2
12 7 13 3 15 15 15 13 1 13 16 13 2
10 2 13 10 9 2 13 10 9 2 2
14 3 2 3 10 15 13 0 1 10 9 1 10 9 2
23 16 16 15 13 10 9 1 10 9 1 9 15 3 4 13 2 15 13 10 9 3 13 2
2 9 2
57 10 9 15 4 13 15 2 9 1 10 11 2 15 10 10 9 3 13 1 13 2 7 15 13 1 10 9 1 10 9 2 7 13 2 7 1 10 9 4 13 1 10 0 2 1 10 9 1 1 10 9 1 9 1 10 9 2
7 7 1 10 9 15 13 2
15 3 2 1 13 15 13 3 2 4 13 1 13 10 9 2
10 3 4 13 3 2 4 3 13 15 2
11 13 10 9 1 10 9 7 1 10 9 2
20 13 16 2 16 4 13 1 10 9 2 1 15 4 4 13 12 9 1 9 2
43 3 13 16 15 15 13 3 2 7 13 15 1 9 2 16 10 9 13 16 2 10 9 16 13 1 13 1 15 2 15 13 10 9 7 15 13 3 10 10 9 1 9 2
33 15 15 13 13 16 10 9 1 9 13 1 13 15 1 10 9 1 10 10 9 2 7 15 13 1 10 9 3 0 7 3 0 2
25 3 13 0 9 1 10 9 16 3 16 10 9 13 1 10 9 3 3 0 1 9 1 9 0 2
14 7 13 3 15 15 13 1 10 11 1 10 9 0 2
8 15 13 1 9 1 10 9 2
24 3 13 2 1 10 9 1 10 9 1 9 2 1 13 10 0 9 2 7 1 13 1 15 2
16 3 2 15 1 15 15 15 13 1 1 13 15 13 1 9 2
25 7 2 1 1 13 15 2 13 1 10 10 9 1 13 15 1 10 0 9 2 16 15 15 13 2
28 7 13 15 10 9 1 10 11 7 15 1 0 1 2 13 2 10 11 2 15 13 13 1 10 9 0 0 2
13 10 11 15 13 7 2 3 2 15 13 0 9 2
20 10 11 15 13 1 10 9 1 10 9 1 11 2 1 11 2 1 11 11 2
6 13 1 10 9 0 2
27 10 9 13 10 9 15 4 13 10 11 1 10 9 2 7 10 11 2 13 0 2 15 13 1 10 9 2
26 3 2 10 9 2 9 9 2 10 9 2 15 13 10 0 9 1 15 10 11 4 13 1 10 9 2
7 1 10 9 1 10 9 2
17 3 10 9 1 10 9 1 11 1 10 9 1 10 9 1 11 2
7 9 0 2 10 9 0 2
6 9 2 10 9 0 2
15 9 2 1 10 9 1 10 10 0 0 2 10 9 0 2
7 10 9 3 15 13 3 2
27 7 10 9 4 13 10 11 1 10 9 1 10 10 9 0 2 1 10 10 9 2 15 3 13 1 13 2
27 10 9 1 9 1 10 9 2 1 10 0 9 13 1 10 9 2 13 1 10 12 5 7 10 12 5 2
13 10 9 13 1 10 0 9 10 9 0 1 9 2
9 7 10 0 9 1 10 0 13 2
27 3 10 9 4 13 1 13 15 2 7 1 0 9 15 13 1 9 1 10 9 1 10 9 1 10 9 2
8 10 9 1 10 10 0 9 2
12 13 10 0 9 1 9 1 10 9 0 0 2
15 7 3 15 13 10 9 15 13 1 15 1 10 0 9 2
22 15 13 9 1 9 2 15 4 13 1 10 9 1 9 1 11 2 7 15 13 3 2
44 15 15 4 13 10 9 0 4 13 13 16 13 1 0 1 10 9 1 9 0 1 11 7 13 15 1 13 3 10 11 1 9 1 9 1 9 1 13 1 15 15 13 3 2
11 15 1 10 9 1 9 13 9 1 9 2
9 7 15 13 9 1 9 13 3 2
7 7 15 13 10 0 9 2
9 7 15 3 13 3 9 1 9 2
13 3 16 4 13 1 9 1 9 2 13 1 9 2
11 9 13 9 1 9 2 9 9 1 9 2
17 7 10 9 1 9 13 10 9 1 11 0 2 9 7 9 0 2
15 7 10 9 3 0 13 1 10 9 0 15 13 10 9 2
20 10 9 13 16 10 9 4 13 1 9 1 9 1 10 9 1 10 10 9 2
8 13 10 9 1 10 10 9 2
21 7 13 10 9 3 1 10 9 15 15 13 16 3 13 16 15 13 1 9 0 2
49 13 10 9 10 9 0 2 7 13 16 15 15 13 3 1 10 9 2 3 7 3 10 0 9 1 10 9 15 13 16 10 9 1 9 13 1 10 9 1 9 13 9 1 9 2 7 13 0 2
16 13 1 12 1 12 9 10 9 1 9 3 13 1 10 11 2
11 7 13 16 2 13 1 10 9 2 13 2
8 2 3 2 3 15 13 2 2
8 2 13 10 0 9 0 2 2
5 7 13 3 0 2
5 11 12 2 12 2
3 9 0 2
13 11 2 16 4 13 3 10 9 1 10 9 13 2
35 3 3 9 0 15 4 13 1 10 9 1 9 1 10 9 0 2 10 9 1 10 9 13 1 13 15 16 10 11 11 7 10 11 13 2
14 3 2 3 2 10 9 4 13 10 9 1 10 9 2
30 10 9 15 10 9 1 10 9 4 13 1 9 1 10 9 1 10 9 0 1 9 1 10 11 11 13 3 10 9 2
10 3 15 13 2 13 13 15 9 0 2
17 10 11 7 10 11 4 13 10 9 1 10 9 0 13 1 3 2
16 10 11 7 10 11 13 1 10 0 9 1 0 9 1 9 2
20 10 11 7 10 11 15 13 13 1 10 9 0 15 13 9 0 13 1 9 2
36 1 11 13 10 9 1 10 9 1 9 0 7 9 2 16 10 9 0 15 13 10 11 13 16 10 9 0 15 13 1 10 9 0 7 0 2
27 15 3 13 10 0 9 16 10 9 1 9 1 9 13 9 1 10 0 9 1 9 1 10 9 0 0 2
14 7 10 9 15 3 13 13 10 9 16 15 4 13 2
17 10 9 2 1 9 2 4 4 13 10 9 0 3 10 9 0 2
20 1 0 9 2 10 9 13 1 10 9 13 13 2 1 10 9 2 3 9 2
49 10 9 0 15 13 1 9 2 7 1 10 0 9 2 7 10 9 0 1 9 0 13 1 13 7 13 10 9 2 13 3 16 10 9 13 10 9 1 9 7 9 1 10 9 2 13 10 9 2
59 10 11 7 2 1 10 10 9 1 0 9 2 10 11 1 10 9 2 11 7 10 11 13 10 9 1 10 9 2 7 10 0 9 15 4 13 4 13 0 9 1 10 11 11 2 1 10 11 11 2 1 10 11 7 1 10 11 0 2
30 1 10 9 2 10 9 1 10 9 13 1 10 0 12 9 15 4 13 1 10 9 0 2 7 0 2 1 9 0 2
17 9 0 1 10 9 0 2 9 1 9 0 7 0 0 3 0 2
32 10 9 1 9 1 9 0 7 9 0 4 13 3 15 10 10 9 2 7 15 13 1 9 15 13 2 3 13 2 10 9 2
14 1 0 9 2 10 9 0 4 4 13 1 9 13 2
25 10 9 1 10 9 1 9 4 4 13 10 9 0 7 13 10 9 0 2 3 4 13 10 9 2
48 1 9 13 16 10 9 1 9 7 1 0 9 13 10 9 1 10 9 7 10 9 0 2 13 9 0 16 10 9 1 10 9 2 16 13 0 2 13 1 13 15 7 10 9 1 13 15 2
31 10 9 15 4 13 10 9 1 10 9 0 1 10 9 3 4 4 13 15 1 10 9 16 3 4 13 10 9 1 9 2
36 1 9 2 10 9 0 13 1 10 9 4 13 10 9 0 1 10 9 1 10 9 0 2 13 16 10 9 13 7 13 16 10 9 4 13 2
18 1 9 2 13 15 10 9 1 9 1 13 10 0 9 0 1 13 2
29 10 0 9 0 13 10 9 0 1 10 9 2 16 10 0 9 13 10 9 1 10 9 0 2 13 10 9 0 2
16 9 1 9 13 4 13 10 9 1 9 2 7 3 13 15 2
15 1 0 9 2 10 9 1 10 9 0 0 13 3 13 2
30 10 9 0 7 0 1 10 11 11 2 1 9 2 15 13 3 3 2 7 3 1 15 2 2 1 9 1 9 0 2
25 1 0 9 2 10 9 0 13 1 9 1 13 15 1 10 10 9 0 2 13 15 1 15 0 2
9 3 2 15 3 13 10 9 0 2
37 10 0 9 0 1 9 1 0 9 1 9 1 10 11 2 10 0 0 9 2 4 13 10 9 0 13 10 9 7 10 9 0 1 10 11 11 2
21 1 10 11 2 15 3 10 11 4 3 13 2 10 9 0 4 13 3 3 13 2
28 1 10 0 9 2 16 10 9 13 1 13 10 9 0 0 7 1 13 10 0 9 2 10 9 15 13 13 2
34 10 9 4 13 1 9 1 10 9 1 9 1 9 15 4 13 1 10 9 1 13 15 1 9 0 16 15 13 0 7 1 0 9 2
33 1 10 9 1 9 2 3 2 10 9 1 10 9 0 1 9 0 13 10 9 1 9 3 0 15 10 9 1 9 0 4 13 2
11 10 9 15 13 1 9 1 10 9 0 2
34 13 0 9 0 1 10 9 1 9 2 7 13 0 1 13 10 0 9 1 9 1 10 9 1 0 2 9 13 0 9 1 9 0 2
23 10 9 3 0 13 10 0 9 1 10 9 0 15 15 4 13 1 13 1 10 9 12 2
37 10 9 0 15 15 4 13 2 9 1 10 9 2 0 9 2 0 9 1 9 1 10 9 0 2 4 13 1 13 10 9 1 10 9 1 13 2
28 13 0 2 16 0 2 13 16 10 9 4 13 3 15 0 1 4 15 13 1 10 0 9 1 9 3 0 2
25 3 2 3 2 4 13 10 9 1 13 1 1 10 9 4 13 10 0 9 1 9 7 9 0 2
5 9 1 11 11 2
5 9 12 2 12 2
8 10 9 0 7 10 9 0 2
57 11 2 9 2 1 10 10 0 9 1 10 9 1 10 9 10 9 1 10 11 11 2 11 11 2 4 13 10 10 9 1 13 1 9 10 11 2 11 11 2 10 9 1 10 9 0 1 10 11 7 10 12 9 1 10 11 2
25 1 10 9 2 10 11 11 7 10 11 4 13 9 1 13 10 10 9 1 10 11 7 15 9 2
51 16 10 9 1 9 0 13 13 10 9 0 1 9 1 10 9 1 9 1 9 2 4 3 3 13 10 9 0 2 7 13 3 10 9 0 1 10 9 0 2 1 15 10 9 0 1 9 1 9 0 2
53 10 9 7 9 1 10 9 13 1 9 0 10 9 1 10 0 9 1 10 9 0 7 10 9 0 13 16 10 9 1 9 0 13 10 9 1 10 9 7 3 4 3 4 13 16 10 9 3 13 10 9 0 2
36 10 9 13 3 0 1 11 15 4 3 13 10 9 1 10 11 7 15 4 13 0 1 10 9 1 10 9 0 1 10 11 9 1 10 9 2
29 16 4 13 10 9 0 1 10 9 2 11 11 2 2 13 0 13 1 10 9 1 9 1 9 10 9 0 2 2
68 1 1 13 10 9 1 9 0 2 10 9 1 9 1 9 2 1 10 11 2 4 13 16 10 9 1 10 9 1 10 9 13 10 9 1 13 10 9 0 0 1 10 9 1 10 10 9 2 1 10 9 1 9 1 9 7 1 10 9 1 10 9 1 9 1 10 9 2
16 3 2 10 9 0 13 0 9 1 10 9 1 10 0 9 2
44 1 10 9 13 1 10 12 1 10 0 9 1 9 0 2 10 9 0 2 9 2 9 2 9 2 9 7 9 0 2 13 10 12 5 1 10 9 0 1 9 1 10 9 2
39 10 9 3 13 3 10 9 1 13 1 13 7 1 4 13 10 10 9 0 2 7 4 1 3 13 3 9 0 13 16 10 10 9 0 13 1 10 0 2
17 10 9 1 9 1 9 13 3 1 13 1 10 13 10 9 0 2
36 3 2 10 9 13 0 9 0 15 13 1 9 2 13 1 10 9 10 9 2 13 10 9 1 10 9 2 13 10 9 7 13 10 9 0 2
58 1 10 9 2 10 11 13 3 10 12 5 1 10 9 0 1 10 9 7 10 9 2 1 10 9 1 10 11 15 2 1 10 9 1 9 1 9 0 3 0 2 15 13 3 10 12 5 2 16 10 11 11 15 13 10 12 5 2
47 10 9 1 10 11 11 13 16 1 10 12 7 10 12 10 9 0 0 1 11 13 0 1 10 12 5 1 10 11 2 7 3 0 1 10 9 1 10 9 13 0 1 3 10 12 5 2
45 1 10 9 0 13 1 10 9 11 11 7 11 11 2 16 10 11 13 10 9 1 9 1 9 0 1 10 11 2 10 9 0 1 9 0 0 13 1 10 12 5 1 9 0 2
74 1 10 9 0 2 3 0 1 10 9 1 10 9 0 2 10 9 3 0 1 10 9 0 4 13 13 10 9 1 10 9 0 0 1 12 9 1 9 10 9 1 12 9 1 9 1 10 12 2 1 10 9 1 10 9 1 10 9 7 1 10 9 0 1 1 12 9 1 9 1 10 0 9 2
22 10 9 1 10 9 0 0 13 3 10 9 1 12 0 9 1 9 1 10 9 0 2
33 16 10 11 13 1 13 10 10 9 1 9 0 1 10 9 1 10 9 0 2 3 3 0 1 15 0 2 10 9 13 3 0 2
20 10 9 0 0 1 10 9 4 3 13 10 12 5 1 9 0 1 10 12 2
42 3 1 10 9 0 2 10 9 0 0 4 13 1 12 9 1 9 2 16 10 9 1 10 9 7 1 10 9 4 13 10 12 9 1 9 13 12 0 9 1 9 2
19 10 0 9 1 10 9 0 1 10 9 0 0 13 10 9 3 3 0 2
49 1 10 0 12 9 2 10 11 4 13 7 13 10 9 1 12 9 13 1 9 0 1 13 10 9 1 10 9 0 2 13 16 10 9 13 1 10 9 1 13 10 9 0 1 9 1 10 9 2
37 1 10 9 2 3 2 13 1 10 9 0 1 13 10 9 13 13 10 9 1 10 9 7 10 9 1 10 9 1 10 9 1 9 1 10 9 2
32 7 10 9 1 10 9 7 10 9 3 13 10 0 2 7 3 0 2 9 1 10 9 1 10 9 1 10 9 0 1 11 2
34 10 9 3 0 2 16 4 13 10 9 1 9 11 10 9 0 2 13 10 9 1 9 2 9 7 9 1 0 9 1 10 9 0 2
28 3 10 9 0 7 10 9 15 15 13 2 3 13 0 1 9 1 10 0 9 1 9 1 9 1 10 9 2
22 3 2 10 9 3 13 9 1 10 9 0 2 1 0 9 1 15 13 10 9 0 2
30 15 2 1 1 10 9 1 10 9 0 0 2 13 10 9 0 10 9 1 9 0 3 1 10 9 1 10 9 0 2
35 1 1 13 10 9 1 10 9 1 10 9 2 10 9 0 1 10 9 0 4 3 13 10 0 9 1 10 11 1 10 9 1 10 9 2
31 3 2 13 3 0 16 10 9 0 1 9 0 13 10 9 16 10 9 0 13 10 9 15 3 10 9 0 4 13 15 2
32 10 9 13 16 10 9 1 10 9 0 13 10 9 0 1 15 10 9 1 10 9 1 9 1 9 3 4 4 13 1 13 2
5 9 1 11 11 2
5 11 12 2 12 2
7 10 9 15 13 10 9 2
56 11 2 10 9 1 10 11 11 11 2 11 2 2 11 11 2 4 13 10 9 1 10 9 1 10 9 1 10 0 9 13 10 9 16 10 9 1 9 1 11 13 7 13 3 12 9 10 9 1 10 11 11 1 10 12 2
11 10 10 9 13 10 0 9 1 12 9 2
43 15 0 7 0 9 0 1 10 10 9 2 7 2 10 9 1 10 9 0 3 0 1 15 1 10 9 0 2 7 10 9 1 10 11 1 10 10 9 1 9 0 0 2
13 3 13 9 0 2 7 10 9 4 3 13 15 2
20 13 10 0 9 0 2 1 9 0 1 0 9 2 4 13 0 1 10 9 2
22 1 11 7 11 2 10 9 4 13 10 9 1 10 10 9 1 13 15 1 10 9 2
7 7 10 9 4 13 0 2
30 1 9 10 0 9 1 9 2 1 15 10 9 0 13 10 9 0 13 15 1 9 7 9 15 4 4 13 3 3 2
24 7 11 13 3 16 10 9 1 10 9 0 13 10 9 1 4 13 1 10 10 9 0 0 2
51 2 13 1 10 9 1 10 9 0 0 2 2 4 13 2 2 13 10 9 1 9 1 10 9 15 15 13 1 10 9 0 7 13 10 9 1 10 9 7 1 10 9 0 0 1 13 1 9 0 2 2
23 13 3 10 9 1 15 4 4 13 10 9 1 11 7 10 9 15 4 13 10 0 9 2
6 7 3 13 1 9 2
39 13 2 1 10 9 1 10 9 9 2 10 9 1 10 9 0 2 9 7 9 2 2 2 16 10 9 13 1 10 9 0 1 10 9 4 4 3 13 2
7 12 9 0 13 0 9 2
60 1 2 10 9 1 10 9 0 2 2 11 11 7 11 11 1 10 11 11 11 13 16 10 9 1 9 1 10 9 0 4 3 13 1 10 12 7 10 12 2 3 1 1 10 9 1 10 9 0 2 13 1 10 12 5 1 10 12 5 2
50 10 12 9 0 15 4 13 10 9 4 13 10 9 1 10 9 7 10 0 9 1 10 9 0 1 10 9 1 10 9 2 13 2 3 1 9 2 1 10 9 0 1 10 9 1 10 9 0 2 2
16 1 9 1 11 7 11 10 9 0 15 4 13 10 0 9 2
37 4 4 13 15 10 9 1 9 1 10 9 7 0 9 13 1 9 1 10 9 2 7 10 9 13 1 10 9 1 9 1 10 9 4 13 0 2
41 1 10 9 13 9 0 7 1 10 15 10 0 9 1 9 13 10 9 1 10 9 0 1 10 10 9 7 13 0 9 0 1 10 9 1 15 10 9 13 13 2
25 11 11 11 7 11 11 1 10 11 11 11 11 2 10 9 15 13 10 9 0 2 15 13 3 2
19 13 16 10 0 9 1 10 9 0 13 10 9 1 10 9 1 0 9 2
29 13 10 9 1 12 9 0 2 13 10 9 0 1 10 9 1 9 1 10 9 0 7 10 9 1 10 9 0 2
21 7 13 0 16 10 9 0 13 1 15 1 10 9 2 3 1 10 9 9 0 2
51 9 7 9 1 9 4 13 1 13 0 9 0 1 10 9 1 10 9 1 10 9 1 9 7 10 0 9 2 3 13 0 1 10 9 1 2 11 11 2 2 3 2 9 9 2 2 2 7 9 0 2
16 7 4 13 10 10 9 1 13 2 13 2 0 7 0 9 2
25 11 7 11 4 13 10 9 1 15 13 3 10 9 15 13 1 9 1 13 3 1 10 9 0 2
12 7 3 13 3 1 10 0 2 9 0 2 2
39 1 10 9 0 10 9 0 1 10 12 2 1 10 15 1 10 11 1 11 7 10 9 0 1 9 1 10 11 11 1 11 4 13 1 13 1 9 0 2
30 2 15 4 3 13 16 13 10 11 7 10 9 3 1 10 0 9 13 10 9 2 7 13 16 15 13 3 0 2 2
9 10 9 13 3 10 0 9 0 2
31 10 9 1 0 9 1 10 9 0 4 3 13 1 10 9 0 2 1 9 16 10 9 0 3 13 1 9 1 10 9 2
32 7 10 9 1 9 1 10 9 1 10 9 13 0 2 7 10 9 1 10 9 13 1 10 9 3 15 13 13 0 7 0 2
13 7 10 9 4 13 9 1 10 0 9 1 11 2
15 10 0 9 9 13 3 3 9 1 10 10 9 1 9 2
29 7 0 9 1 10 9 15 13 9 1 10 9 0 2 10 9 11 7 10 9 9 2 1 9 2 4 3 13 2
46 15 15 13 1 10 9 0 7 1 10 0 9 1 10 0 9 0 2 3 13 16 1 9 10 9 1 2 9 9 2 1 10 11 15 13 0 1 15 4 13 10 9 1 10 9 2
5 9 1 11 11 2
8 10 9 1 10 11 4 13 2
19 11 11 2 1 10 9 1 9 2 10 9 0 4 13 10 9 3 0 2
39 3 1 10 10 9 0 2 10 9 1 9 0 3 1 9 7 9 13 1 9 1 9 7 9 1 10 9 1 9 4 13 10 9 1 9 1 9 0 2
12 15 4 13 10 9 2 7 10 9 4 13 2
21 10 9 13 15 1 10 9 0 15 13 1 9 13 1 10 9 0 1 10 9 2
10 3 4 4 13 10 9 1 10 9 2
17 10 9 1 10 9 1 10 9 0 1 11 11 13 10 9 13 2
23 1 9 0 2 10 9 0 4 13 15 7 1 0 9 7 1 9 1 10 9 3 0 2
29 1 0 9 2 10 9 1 10 9 0 1 15 13 1 11 13 1 16 13 1 10 9 1 9 1 10 9 0 2
38 10 9 1 10 9 15 13 1 9 0 7 1 9 13 9 1 9 3 0 2 7 10 9 1 10 9 1 10 9 13 1 10 9 13 1 10 9 2
36 16 10 9 4 13 10 9 0 1 10 9 0 1 11 10 12 9 2 10 10 9 1 13 2 10 9 2 13 1 0 0 10 9 1 13 2
26 10 9 4 13 15 1 13 1 9 3 13 1 10 9 1 10 9 0 1 10 9 1 9 1 9 2
14 10 13 7 15 1 10 9 13 1 3 13 10 11 2
36 10 0 4 13 10 10 9 1 10 11 11 15 13 15 0 3 9 2 1 10 9 1 10 9 15 13 11 9 7 9 10 15 1 10 15 2
27 13 1 10 9 16 10 11 4 13 3 3 0 1 10 11 1 10 9 1 10 11 1 10 9 1 9 2
20 16 13 2 10 11 1 10 9 0 4 13 10 15 7 13 3 1 10 11 2
54 3 2 3 16 10 9 1 10 9 0 1 10 9 3 0 1 10 11 4 13 10 0 9 0 2 10 11 2 1 1 10 9 0 0 2 13 3 10 9 1 9 1 9 1 9 1 13 10 9 1 10 9 0 2
18 7 3 13 1 13 10 9 0 1 15 13 10 11 1 10 0 9 2
19 4 13 10 11 11 1 11 1 10 12 2 3 16 10 9 13 10 9 2
25 10 9 3 4 13 1 10 0 9 2 7 15 4 13 1 9 1 15 4 13 1 10 9 0 2
28 10 9 3 13 0 1 13 10 0 9 1 10 0 1 13 9 0 0 2 3 10 9 0 0 7 0 2 2
15 7 10 11 13 9 1 9 0 15 3 10 11 4 13 2
10 9 1 10 9 7 9 1 10 9 2
54 1 10 0 9 1 10 9 1 10 11 0 13 1 10 9 12 2 10 9 1 10 9 7 10 9 1 10 9 13 10 9 1 10 0 9 1 10 9 0 7 0 2 15 13 10 9 0 1 10 9 1 9 0 2
25 10 11 2 1 10 10 9 0 1 0 9 7 10 9 13 2 13 10 9 3 0 1 10 9 2
51 7 13 10 9 13 10 9 1 10 9 0 1 10 10 9 1 10 10 9 7 1 10 9 1 10 0 9 2 3 13 10 9 0 7 10 0 9 1 9 15 4 13 9 0 7 0 1 10 0 9 2
46 1 1 13 10 9 0 0 2 10 11 4 13 10 9 1 13 10 9 1 10 9 0 7 13 15 1 13 10 10 9 0 2 1 0 9 13 1 9 1 9 7 9 1 10 9 2
26 10 9 0 1 13 10 9 1 10 0 9 1 9 13 1 13 15 1 9 0 13 1 10 9 0 2
35 1 13 10 9 2 10 9 0 1 10 9 7 10 9 2 11 2 4 13 1 9 1 1 9 0 7 0 2 16 4 13 1 11 0 2
51 10 11 4 3 13 10 10 9 0 1 10 9 13 7 13 1 10 9 3 7 3 0 1 10 9 0 2 16 10 11 13 10 9 1 10 9 1 10 9 0 7 15 13 1 13 15 1 10 9 0 2
18 13 7 13 16 10 11 1 10 9 0 13 1 10 9 1 10 9 2
22 13 1 10 9 16 10 11 4 13 10 9 7 10 9 1 10 10 9 13 1 11 2
32 3 2 10 11 13 1 10 0 0 1 10 9 11 2 1 10 15 10 11 11 4 13 1 13 10 11 1 10 0 9 0 2
15 10 11 4 13 3 10 0 9 10 9 13 1 10 11 2
7 4 3 13 1 10 9 2
23 10 9 11 3 13 10 9 0 2 3 13 10 9 1 10 11 1 9 1 10 9 0 2
31 10 9 1 10 9 0 13 9 0 7 1 10 11 7 1 10 11 2 7 3 1 10 11 2 15 15 13 1 10 9 2
21 10 11 13 1 10 9 0 2 7 13 10 9 1 10 9 0 1 10 10 9 2
10 4 3 13 0 9 1 10 10 9 2
31 10 9 11 11 4 13 15 1 10 9 11 11 1 13 16 10 11 13 10 9 2 7 3 10 9 2 1 10 9 0 2
5 11 12 2 12 2
7 10 9 1 10 9 0 2
44 11 11 2 3 10 9 2 10 9 1 15 4 13 1 10 9 13 2 1 9 9 1 10 9 1 10 9 0 2 15 1 10 9 1 10 12 13 13 1 10 9 1 9 2
22 10 9 1 9 15 15 15 13 2 3 2 4 13 10 9 1 10 13 9 1 9 2
19 10 9 1 10 0 9 1 9 13 1 10 11 11 4 13 1 9 13 2
38 10 9 13 3 0 1 10 9 1 9 0 2 1 9 10 11 2 10 11 2 10 11 2 10 11 7 10 11 2 13 3 9 1 13 10 9 0 2
34 7 10 9 1 10 9 1 10 11 13 3 0 2 7 10 0 9 1 10 0 2 9 0 2 1 10 9 0 4 13 3 3 0 2
12 1 10 9 1 10 9 2 15 13 1 13 2
12 1 10 9 2 3 2 13 13 10 9 13 2
54 1 9 1 10 9 13 0 1 10 9 2 15 3 13 1 0 9 2 7 10 10 9 13 1 9 0 15 1 10 9 0 13 1 10 9 0 1 10 9 1 10 9 12 2 10 11 13 10 9 1 10 9 0 2
29 3 2 3 13 10 9 1 9 1 10 9 1 9 1 9 1 10 9 1 10 9 1 9 1 9 1 10 11 2
34 7 2 3 2 10 0 9 0 1 10 11 2 0 1 12 9 1 9 1 9 1 9 0 2 13 10 0 9 1 9 1 9 0 2
18 3 2 10 9 0 4 13 2 7 10 9 1 15 3 4 3 13 2
30 10 9 1 10 9 3 13 15 1 16 13 1 10 9 15 13 0 9 13 2 1 10 9 2 15 13 10 9 0 2
33 3 13 2 3 2 7 0 7 0 1 10 11 13 10 9 1 10 12 5 1 9 0 15 4 13 10 12 9 0 1 10 12 2
61 7 2 13 10 0 9 1 10 9 1 10 9 0 1 10 11 2 7 15 13 3 16 10 9 1 10 12 5 2 0 1 10 9 0 1 10 12 2 12 5 2 4 13 1 10 9 1 10 9 1 10 3 0 9 1 9 1 10 9 0 2
62 10 9 0 13 16 10 0 9 1 10 11 3 13 16 10 9 1 0 9 0 2 10 9 15 13 10 9 0 7 13 1 10 9 1 9 0 2 15 13 1 10 9 0 7 1 10 9 0 1 10 9 0 7 1 10 9 1 10 9 0 9 2
21 3 16 10 9 3 4 13 2 15 1 15 13 1 10 9 1 10 9 1 9 2
23 1 9 2 10 9 1 10 9 1 9 13 10 9 0 1 10 13 9 1 10 9 0 2
56 1 0 9 2 15 1 15 4 13 13 10 9 1 10 0 9 1 10 9 0 13 1 10 9 7 1 10 9 2 9 1 10 0 9 0 2 1 10 9 1 9 1 10 9 1 10 9 7 1 10 9 3 0 7 0 2
32 1 10 12 2 3 2 10 9 1 10 9 0 4 13 10 3 0 1 10 9 2 13 10 9 13 1 10 9 0 7 0 2
54 10 9 2 16 4 13 1 10 10 0 9 11 2 10 11 1 11 7 11 2 3 13 10 11 2 7 10 9 0 2 7 10 11 11 1 9 2 15 3 13 0 1 13 10 9 1 10 9 0 15 10 9 13 2
30 10 9 1 9 13 10 9 1 10 9 0 2 16 12 9 2 1 9 7 9 2 15 13 1 9 7 1 9 0 2
45 1 0 13 2 10 9 13 1 10 9 1 9 2 0 9 7 2 3 2 1 10 9 0 2 1 3 16 15 7 10 10 9 3 13 1 13 15 7 1 13 1 10 10 9 2
17 10 0 0 1 10 9 15 13 1 11 11 7 11 1 9 0 2
23 10 0 9 0 13 1 10 9 2 13 1 10 9 12 2 3 4 13 1 10 9 0 2
30 1 10 9 10 2 10 11 11 4 13 9 1 10 9 0 1 0 9 1 13 10 9 1 9 1 10 9 3 13 2
60 3 2 4 13 1 13 1 10 9 1 9 1 10 11 1 13 10 10 9 1 9 2 10 3 0 1 10 9 2 2 7 4 13 10 0 9 0 1 9 1 10 9 0 1 13 1 13 0 9 1 9 7 13 10 0 9 1 9 0 2
44 1 10 12 9 4 13 9 1 10 0 9 1 9 2 1 15 10 9 2 10 9 1 9 1 10 9 2 10 9 0 2 10 9 0 7 10 9 0 2 1 13 15 15 2
26 7 2 3 16 4 13 10 9 2 15 1 10 9 2 10 11 2 4 13 1 13 1 10 10 9 2
35 10 9 1 10 11 13 1 10 9 1 13 10 9 1 9 2 15 4 13 1 13 10 9 1 9 0 7 13 10 9 1 10 9 0 2
20 1 9 1 15 2 10 11 3 13 3 3 0 1 13 9 1 10 11 11 2
24 1 10 9 0 1 9 1 15 0 2 10 9 1 10 9 0 2 9 4 13 10 9 0 2
10 15 1 10 0 9 13 0 1 9 2
10 10 15 2 3 2 13 10 0 9 2
39 1 10 9 2 10 11 11 4 13 9 1 10 9 2 1 9 15 1 10 11 0 2 15 3 13 10 10 0 9 1 10 9 1 9 7 9 1 9 2
14 1 1 0 9 13 2 10 11 13 1 10 9 0 2
34 1 10 9 0 0 1 10 9 1 10 9 12 4 13 1 10 9 3 0 1 10 9 2 7 13 10 9 16 3 3 13 10 15 2
19 10 9 13 0 2 1 10 11 2 10 11 7 10 9 1 10 9 0 2
5 9 1 11 11 2
5 9 12 2 12 2
8 11 2 11 7 10 9 0 2
23 11 2 10 9 16 10 9 15 15 13 3 1 10 9 13 10 9 0 1 10 9 0 2
37 1 9 2 10 0 9 1 10 9 0 4 13 10 9 2 13 13 10 9 1 9 1 10 0 9 2 1 10 9 1 9 1 9 7 9 0 2
35 3 1 10 9 1 9 1 9 10 0 9 1 10 9 4 13 1 13 10 13 9 1 10 9 1 9 7 4 3 13 0 9 1 9 2
15 7 10 0 9 2 3 1 10 9 0 2 13 10 9 2
31 3 2 10 9 1 10 9 0 1 10 9 1 10 9 1 10 9 2 1 11 11 1 11 11 2 15 4 13 3 0 2
12 10 9 0 4 13 10 9 1 10 9 0 2
31 10 9 0 0 2 3 0 2 3 3 2 4 13 16 10 0 9 1 10 9 15 13 9 2 16 15 3 15 1 15 2
22 1 9 2 10 9 1 11 1 10 9 1 9 3 15 4 13 1 10 9 0 0 2
38 7 2 1 10 0 9 1 10 9 1 9 1 10 9 1 10 0 9 2 10 9 1 0 9 13 3 10 9 1 11 1 15 10 9 13 10 9 2
12 10 9 1 9 1 10 10 9 13 1 13 2
23 7 10 0 9 1 10 9 3 13 9 1 9 1 10 9 0 1 10 9 1 10 9 2
22 13 1 9 10 0 9 0 2 13 0 9 1 13 2 3 13 1 9 7 9 0 2
21 10 0 9 1 9 13 9 13 15 13 10 9 2 10 9 0 13 10 9 0 2
30 16 10 9 0 13 3 2 0 2 3 1 10 9 1 10 9 7 1 10 9 2 10 9 4 13 1 13 9 0 2
27 3 13 10 0 9 1 10 9 1 4 13 10 0 9 1 10 9 0 7 1 10 9 1 10 9 0 2
30 10 0 9 1 9 13 10 9 1 13 16 10 9 0 4 13 16 3 0 2 15 13 10 9 1 10 10 9 0 2
46 3 15 4 3 13 1 0 10 9 2 1 10 9 16 10 9 1 9 7 9 4 13 10 9 7 10 9 1 9 1 10 9 1 10 9 2 3 16 4 4 13 10 9 1 9 2
37 3 10 10 9 15 4 13 3 0 1 10 13 15 1 10 2 0 9 2 2 7 1 10 9 1 10 9 3 0 1 10 9 1 10 9 0 2
43 7 10 9 1 10 9 1 10 0 9 4 13 0 9 2 13 1 10 0 9 1 9 1 10 9 1 10 9 2 1 9 3 1 9 1 10 3 0 7 10 10 15 2
21 10 9 4 13 7 13 10 9 0 1 10 9 2 7 10 9 0 15 15 13 2
22 10 0 9 13 10 9 0 2 10 9 15 13 9 0 3 1 10 9 0 3 13 2
31 10 9 1 10 9 0 3 13 10 9 2 16 1 10 0 9 4 13 7 1 13 10 10 9 7 1 13 10 10 9 2
40 10 9 0 13 10 0 9 1 9 15 13 10 9 1 10 9 1 0 9 1 9 1 10 9 15 3 13 3 10 9 7 10 9 1 13 15 1 9 0 2
17 4 3 13 16 4 13 10 0 9 1 10 9 0 1 0 9 2
9 15 13 9 0 1 10 0 9 2
34 10 9 0 13 10 9 0 2 10 9 3 10 9 4 3 13 9 3 3 13 3 7 3 13 16 3 3 10 9 4 13 1 13 2
50 15 15 15 13 3 13 16 10 9 0 4 13 0 1 10 9 2 1 10 0 9 1 10 9 1 9 1 9 12 7 9 0 2 15 15 13 10 0 9 0 1 10 9 1 9 1 10 0 9 2
23 10 9 0 1 9 1 9 2 13 11 11 2 11 11 7 11 11 2 4 13 10 9 2
23 10 9 0 1 3 2 3 1 2 9 1 10 0 9 1 9 2 15 4 13 3 0 2
50 10 9 0 1 10 9 13 2 15 10 9 13 1 10 2 9 2 2 4 13 10 9 1 10 9 1 15 15 15 13 0 2 7 4 3 13 1 9 1 10 9 2 1 10 9 1 10 9 0 2
19 7 3 2 1 10 0 9 1 9 1 9 2 10 9 0 4 13 13 2
34 13 10 9 13 10 0 9 1 9 0 0 2 1 1 9 13 1 10 9 1 10 0 2 3 13 10 9 3 0 1 10 0 9 2
36 10 9 0 13 1 10 9 1 10 9 0 4 4 13 13 10 9 1 10 9 0 7 13 10 9 7 9 1 13 7 13 1 10 9 9 2
16 7 15 15 13 10 9 1 13 9 10 9 1 10 15 0 2
23 10 9 0 4 13 3 0 1 10 13 10 0 9 1 9 0 2 3 1 10 0 9 2
50 16 15 13 1 9 0 2 1 10 9 2 10 9 2 10 9 7 10 0 9 2 10 9 1 3 13 3 13 2 7 10 9 0 1 10 9 4 13 13 1 0 9 1 10 9 1 10 9 0 2
19 10 9 0 13 1 13 1 10 0 9 1 10 9 1 1 10 10 9 2
23 1 10 9 1 9 1 9 15 3 4 3 13 10 9 0 2 10 9 13 3 3 3 2
20 1 10 9 0 2 16 3 3 10 9 4 13 3 2 10 9 4 13 0 2
5 9 1 11 11 2
5 9 12 2 12 2
6 10 9 1 10 9 2
21 11 11 2 1 10 10 9 15 13 10 0 9 1 10 9 0 0 1 11 11 2
22 1 10 9 2 10 9 1 10 11 13 10 10 0 9 0 2 15 15 13 1 13 2
7 7 13 10 9 1 13 2
15 13 0 13 10 9 1 10 9 1 10 9 1 10 9 2
25 15 15 13 3 13 0 1 10 9 1 10 9 0 2 1 10 9 1 10 9 1 10 9 9 2
40 1 10 12 10 9 11 11 2 13 10 11 11 1 10 10 0 9 1 10 9 2 13 16 2 10 9 0 15 13 3 1 16 1 10 9 1 10 9 2 2
8 4 13 15 10 9 1 9 2
22 3 10 9 3 13 3 10 9 1 10 9 1 9 13 1 10 9 1 10 9 0 2
14 16 4 13 2 15 13 15 1 9 1 10 10 9 2
29 15 13 1 16 10 9 0 2 3 3 1 10 9 1 11 11 2 10 9 0 15 13 1 10 10 9 1 9 2
25 13 16 10 9 0 13 10 0 7 10 3 9 1 10 10 9 2 3 15 4 13 15 1 15 2
46 1 10 9 3 0 2 3 2 13 0 16 0 9 1 10 9 13 13 9 0 1 13 10 15 2 13 10 9 1 4 13 2 3 1 10 0 9 2 7 13 10 9 1 10 9 2
29 1 10 9 2 16 10 9 13 1 10 9 2 0 2 2 10 9 1 10 9 13 3 0 16 1 10 9 0 2
40 3 1 10 9 0 3 15 13 1 10 9 1 10 9 1 9 2 16 3 1 10 9 2 2 7 1 10 9 13 1 10 9 1 15 3 3 15 4 13 2
13 10 9 0 0 1 10 10 2 9 2 13 0 2
36 1 9 0 2 10 9 11 2 11 15 4 13 10 9 4 13 1 10 9 2 10 9 9 1 10 15 15 4 13 9 1 9 7 9 0 2
16 10 9 3 13 1 9 10 0 9 1 9 7 10 9 0 2
47 7 3 13 9 0 13 3 10 9 1 9 13 1 10 9 0 7 10 9 1 9 1 9 13 1 10 0 9 2 1 10 9 1 9 1 10 9 9 2 13 1 10 10 9 1 9 2
6 12 9 4 13 0 2
29 10 0 13 16 10 9 1 10 9 3 3 13 10 9 0 1 13 10 10 9 0 1 10 10 9 1 10 9 2
50 1 10 10 9 1 10 2 9 13 15 2 2 10 9 0 15 13 10 0 9 9 1 10 9 9 7 10 9 1 9 1 9 4 13 15 1 10 9 13 9 1 13 9 1 9 2 13 0 9 2
17 7 1 10 9 1 9 2 15 1 10 9 4 3 13 1 15 2
18 10 9 0 1 10 9 9 1 10 9 0 4 1 9 13 3 0 2
61 3 2 16 10 9 2 1 10 9 11 1 10 9 0 2 13 1 10 0 9 2 15 1 10 9 0 2 7 10 9 1 15 15 4 13 7 10 0 9 0 1 10 9 1 10 9 1 9 1 15 13 2 15 13 1 10 9 1 10 9 2
27 1 9 0 2 10 10 9 9 3 13 10 9 1 10 0 9 13 1 10 9 15 13 1 13 10 9 2
18 7 3 3 13 1 9 0 10 9 1 10 9 0 13 1 10 9 2
37 1 10 9 3 0 2 3 10 9 13 3 10 9 1 10 9 1 9 2 1 9 2 1 10 9 2 13 0 13 10 9 1 10 9 1 15 2
10 7 15 13 3 3 0 1 0 9 2
50 3 4 13 1 9 0 10 9 16 2 9 1 10 9 13 1 9 0 2 10 9 0 13 1 13 0 9 3 1 1 9 2 13 1 10 0 9 1 10 9 1 9 7 1 10 9 1 10 9 2
39 3 15 4 3 13 16 2 1 10 9 2 10 9 1 10 0 9 0 1 10 9 1 0 9 1 10 9 1 9 4 13 3 0 1 15 13 10 9 2
36 4 4 13 10 9 0 1 10 13 9 0 1 13 10 9 13 1 10 9 7 1 10 9 2 13 10 9 2 3 10 0 9 1 10 9 2
38 7 10 9 1 9 4 4 13 1 3 16 10 10 9 0 4 4 13 1 10 9 3 0 2 7 1 10 9 3 13 15 4 4 13 1 0 9 2
22 3 2 10 13 3 0 10 15 1 10 15 2 1 11 7 11 2 13 10 10 9 2
37 7 3 4 13 10 9 1 15 1 10 9 2 10 9 2 10 9 1 11 7 10 9 1 10 9 0 2 15 4 13 15 10 9 1 9 0 2
8 4 3 13 10 9 1 9 2
42 3 16 3 13 15 10 0 9 0 4 13 1 10 10 9 2 3 13 16 2 3 1 10 9 1 9 0 15 4 13 10 9 0 0 2 9 2 10 9 13 0 2
5 9 1 11 11 2
5 9 12 2 12 2
7 10 11 11 1 10 9 2
29 11 2 10 9 0 2 10 11 11 11 1 10 9 1 11 4 13 10 10 0 9 1 10 9 13 1 11 11 2
20 10 9 1 10 9 4 13 2 10 9 7 10 9 0 7 1 10 9 2 2
34 10 9 0 1 10 9 1 9 2 13 1 11 11 2 9 1 10 11 11 11 2 13 10 9 13 12 0 9 0 1 13 10 9 2
31 15 13 0 7 0 2 16 10 15 13 0 2 0 2 1 1 9 10 9 1 9 2 7 13 1 10 0 9 1 9 2
5 10 9 13 0 2
12 3 15 13 10 9 1 10 0 9 1 9 2
11 3 2 15 3 13 10 9 1 9 0 2
44 10 9 1 9 1 10 9 2 10 9 0 2 10 9 0 2 0 7 10 9 0 1 10 9 1 10 9 2 7 2 1 9 2 1 10 9 0 7 0 2 4 3 13 2
18 10 9 13 16 10 9 3 4 13 10 9 1 0 9 1 9 0 2
18 7 10 0 2 3 3 13 9 0 2 10 9 0 2 4 13 15 2
28 1 10 9 1 11 2 15 13 1 1 10 2 9 2 7 10 2 13 2 13 1 13 10 9 1 10 9 2
27 3 2 3 1 10 9 0 2 10 0 9 0 4 13 0 1 13 10 9 7 10 9 1 10 9 0 2
13 7 10 9 7 10 9 4 13 3 10 0 9 2
55 10 9 1 10 9 0 13 1 0 9 7 13 10 9 1 10 9 1 9 0 7 1 10 9 2 10 0 9 1 10 9 2 7 9 0 0 15 4 13 10 9 1 10 9 0 1 0 9 1 10 0 9 1 9 2
26 3 2 10 9 0 4 13 10 9 1 9 0 1 10 9 2 10 9 7 10 9 0 1 9 0 2
59 4 4 13 1 10 13 16 10 9 13 1 10 0 9 1 10 10 9 2 1 9 16 13 10 0 9 7 16 3 4 13 1 9 0 2 9 15 4 13 10 9 0 16 10 9 7 10 9 13 10 0 9 1 10 9 1 10 9 2
36 3 2 16 4 13 10 0 9 2 10 9 0 9 0 4 13 16 4 13 3 0 1 10 9 16 13 1 9 16 4 13 15 15 13 3 2
34 10 9 1 10 9 4 13 16 9 0 1 13 9 0 2 9 1 10 9 1 10 9 0 1 10 9 0 7 0 13 1 0 9 2
37 1 15 2 16 10 9 3 0 13 9 0 1 10 9 1 10 9 1 10 10 9 2 10 9 4 4 13 10 9 1 10 9 1 10 9 0 2
16 10 9 0 9 4 3 13 1 10 9 1 9 1 9 0 2
33 10 9 1 10 9 7 1 10 9 1 10 9 0 1 10 9 1 9 0 13 1 1 10 9 0 2 16 3 15 13 10 9 2
47 13 10 0 9 4 13 10 9 1 15 10 9 1 10 9 13 10 9 1 10 10 9 2 3 13 0 16 10 9 13 3 0 1 15 13 10 9 1 0 9 1 10 9 1 10 9 2
16 7 10 9 0 13 0 2 7 13 16 15 13 1 10 9 2
10 10 0 9 13 16 15 13 10 9 2
47 9 1 9 1 9 3 1 10 9 2 9 0 1 10 9 1 9 2 9 0 1 10 9 2 9 1 9 0 2 10 9 0 1 9 2 15 4 15 13 0 1 10 13 10 9 0 2
13 10 9 4 4 13 1 9 15 13 9 0 0 2
25 1 13 10 9 1 13 10 9 15 13 9 1 10 0 9 1 9 15 13 9 1 10 10 9 2
42 1 11 2 10 9 0 1 10 9 15 10 9 1 9 0 4 13 1 10 9 1 10 9 0 2 10 9 0 1 10 9 9 2 4 3 13 10 9 1 10 9 2
36 9 13 1 13 10 9 0 1 10 9 13 3 15 0 2 3 1 15 16 4 13 10 9 1 13 9 1 10 10 9 16 13 1 10 9 2
36 4 4 13 1 10 9 10 9 1 9 1 10 9 9 2 15 4 13 16 0 9 1 10 9 1 10 9 1 10 9 0 1 10 11 11 2
26 10 9 1 10 9 1 10 11 11 4 13 1 13 10 9 3 3 0 1 10 9 7 10 9 0 2
19 7 2 1 10 0 9 0 1 10 9 2 10 9 1 10 9 4 13 2
27 4 13 10 9 1 13 16 15 13 1 10 9 2 7 13 2 9 2 10 9 1 15 10 9 4 13 2
5 9 12 2 12 2
11 10 9 1 10 11 1 10 9 13 9 2
40 11 2 1 10 0 12 9 10 11 1 10 9 4 13 0 9 1 9 0 2 13 10 9 8 8 1 12 9 1 10 12 1 15 1 12 9 10 0 9 2
50 3 3 2 10 10 9 1 9 13 13 2 7 15 1 9 1 10 13 9 1 10 10 9 1 9 0 2 13 1 13 10 12 5 1 10 12 2 7 10 0 9 1 10 11 7 1 0 9 13 2
39 1 10 9 1 13 10 9 2 10 11 1 10 9 4 13 9 0 7 13 10 9 1 9 0 2 13 3 1 13 10 10 9 0 2 1 9 10 9 2
31 10 9 1 10 11 1 10 9 1 10 0 0 9 13 15 1 10 0 9 1 10 10 9 9 1 10 0 9 1 9 2
29 1 10 12 7 10 12 2 10 9 1 0 1 10 9 1 9 0 4 13 1 10 12 5 1 3 10 12 5 2
50 13 10 9 2 13 10 9 1 10 9 7 13 10 9 7 10 9 1 9 0 2 10 9 1 9 1 10 0 9 1 9 4 13 10 9 1 9 1 10 9 1 9 13 1 10 9 1 10 9 2
16 7 10 9 13 13 2 1 9 1 10 9 1 10 10 9 2
45 1 9 2 1 13 0 10 9 1 9 4 13 1 13 0 7 0 9 0 1 10 9 2 3 1 10 9 1 9 1 9 3 0 7 10 9 1 10 9 0 3 0 7 0 2
24 1 10 9 2 4 13 16 10 11 1 10 9 4 13 10 10 9 1 10 0 9 1 9 2
51 10 9 1 9 1 9 1 10 9 1 9 1 10 9 1 9 0 7 0 13 0 2 7 10 9 1 10 9 1 9 1 9 1 10 9 9 2 9 7 1 10 9 0 4 13 3 1 10 0 9 2
19 1 10 12 2 10 9 4 13 10 10 0 9 9 2 11 11 2 11 2
20 1 9 1 9 1 10 9 0 2 3 2 10 9 1 9 13 7 13 0 2
44 1 10 9 13 1 10 11 2 3 10 12 5 1 10 9 1 9 0 1 10 12 7 10 12 9 13 9 1 10 9 9 2 1 10 9 1 10 12 5 1 10 9 0 2
30 10 9 1 9 1 10 9 9 0 2 3 2 15 13 1 1 10 12 5 2 3 13 10 0 11 1 10 12 5 2
46 10 9 1 9 1 10 9 9 1 10 9 1 10 9 3 0 13 1 10 12 5 2 3 0 1 1 15 1 10 9 15 4 13 3 10 9 0 7 0 2 0 1 10 12 5 2
24 3 2 3 1 10 9 0 3 0 7 0 10 9 1 10 9 13 10 0 9 1 10 9 2
26 1 9 2 1 1 10 12 9 10 10 9 1 10 9 9 1 9 13 0 1 15 1 10 9 11 2
45 13 10 9 2 3 2 10 9 13 3 1 10 12 5 1 10 12 5 16 9 1 9 3 0 7 10 9 1 9 1 10 9 0 13 1 15 0 13 1 13 1 10 10 9 2
17 10 0 9 13 16 10 9 11 4 13 1 13 10 9 1 9 2
19 15 15 13 3 0 13 16 10 9 13 13 0 9 1 9 1 10 9 2
40 1 10 9 15 13 2 1 9 2 15 1 13 9 1 9 0 13 3 10 9 11 2 11 2 7 13 9 1 10 9 15 13 1 13 10 10 9 1 9 2
33 3 2 1 10 9 16 10 9 9 0 13 3 10 9 0 1 9 0 2 13 10 9 0 4 13 15 0 1 13 10 9 0 2
23 10 9 0 13 15 15 13 10 9 1 9 1 9 1 9 1 10 9 1 10 9 0 2
42 1 10 9 0 2 3 16 10 9 1 10 9 13 1 10 12 5 1 10 9 1 10 9 2 10 10 9 1 9 13 3 1 10 1 3 1 15 1 10 9 0 2
55 10 9 13 1 10 9 1 10 9 0 1 0 9 2 1 10 9 1 10 9 7 1 10 9 7 10 9 2 13 1 10 9 1 9 9 0 7 1 0 9 1 10 9 2 10 9 2 10 9 0 7 10 9 0 2
19 13 3 0 13 10 9 1 10 9 1 10 9 7 10 10 9 1 9 2
34 10 0 9 2 3 2 13 1 13 10 9 1 9 2 13 10 9 1 13 9 3 13 2 1 1 13 15 15 9 7 10 9 0 2
45 10 9 0 2 1 9 2 13 3 3 0 1 13 9 0 1 10 0 9 11 2 9 2 9 2 9 7 9 2 2 9 9 10 9 1 9 2 1 10 9 7 10 9 0 2
37 10 9 1 9 1 10 9 0 7 0 4 13 1 13 10 10 9 2 13 1 0 9 1 9 10 9 0 1 13 10 9 0 1 9 0 0 2
25 3 2 10 0 9 1 9 0 7 0 1 10 9 0 0 3 4 13 1 10 11 1 10 9 2
37 3 10 0 9 0 11 11 4 13 1 10 9 16 10 0 9 0 1 10 9 9 13 0 1 13 1 13 10 9 1 9 0 1 10 10 9 2
21 10 9 13 16 10 9 0 13 0 1 13 9 1 10 10 0 9 1 9 0 2
5 9 1 11 11 2
5 9 12 2 12 2
16 10 9 1 9 1 10 9 0 0 2 3 16 13 13 15 2
19 11 2 3 2 10 11 1 10 11 4 13 3 3 1 1 10 0 9 2
36 16 15 13 1 10 9 15 13 10 9 2 15 13 3 10 9 0 1 10 9 2 10 9 7 10 9 2 7 10 9 0 7 1 10 9 2
12 15 13 3 1 10 9 15 15 13 11 11 2
23 11 13 10 9 0 15 13 9 2 9 7 9 1 10 0 9 1 9 1 10 11 0 2
30 16 15 4 13 1 10 12 2 4 3 13 1 9 10 0 9 1 9 13 1 10 9 13 1 10 9 1 10 11 2
36 3 1 10 9 1 10 9 0 1 10 9 15 4 13 10 9 1 0 9 1 10 9 13 1 11 2 10 9 1 10 9 4 3 13 3 2
52 1 10 9 10 10 9 4 4 13 10 9 2 7 3 3 9 1 10 9 1 10 9 10 9 1 11 4 13 1 13 9 0 1 9 7 3 10 9 3 0 1 13 10 9 1 10 9 1 10 10 9 2
18 16 13 10 9 1 11 2 10 9 13 0 1 10 9 1 10 11 2
30 10 9 13 10 12 5 1 10 9 9 0 2 13 10 9 1 10 10 9 7 10 9 9 1 13 10 9 3 0 2
26 10 9 13 16 10 9 1 10 9 0 13 10 9 3 0 1 13 10 9 1 10 11 0 2 0 2
30 1 9 2 10 9 1 10 9 13 1 10 9 0 10 0 9 1 13 10 9 0 1 9 1 10 9 0 1 9 2
29 3 16 10 9 7 10 11 11 1 10 10 9 4 13 10 12 1 10 9 1 10 9 0 7 0 1 10 11 2
12 10 9 1 11 13 0 3 1 10 0 9 2
26 10 10 9 13 0 1 10 9 1 10 11 3 3 16 13 10 9 0 2 7 3 16 13 10 9 2
55 13 3 9 2 1 10 11 11 2 13 1 13 10 0 9 1 15 10 9 7 10 9 13 10 9 7 15 13 13 1 10 9 2 1 10 9 2 7 1 10 9 1 10 10 9 2 7 3 1 9 9 1 10 9 2
47 15 15 4 13 3 13 16 2 16 10 11 13 1 13 10 9 0 2 10 9 1 10 9 4 3 13 3 15 1 10 0 9 15 13 1 10 9 1 13 2 7 10 0 9 1 9 2
27 10 9 3 13 10 9 1 9 0 2 7 3 10 9 1 10 9 0 13 9 2 7 13 3 10 9 2
26 1 10 10 9 2 10 9 0 13 1 9 13 1 13 15 1 9 1 9 1 15 13 1 10 9 2
41 15 13 2 3 1 10 12 2 10 9 1 9 0 1 10 9 1 9 2 7 10 9 0 1 10 9 2 1 10 9 7 1 10 9 1 10 9 13 3 0 2
34 1 13 1 13 3 10 9 2 10 11 0 7 10 11 11 4 13 3 10 9 1 9 1 10 9 15 10 9 0 15 13 1 13 2
9 10 9 13 1 3 10 9 0 2
12 10 9 1 9 13 0 7 1 10 9 0 2
38 16 15 13 10 9 7 10 9 0 1 10 9 1 9 1 9 1 0 9 7 9 2 10 9 1 9 4 13 1 1 10 12 5 2 1 1 11 2
41 1 9 2 10 9 13 16 10 9 0 1 10 9 13 1 3 16 10 9 0 13 10 9 1 9 1 10 9 0 1 10 9 2 10 9 7 3 10 9 0 2
11 7 3 13 16 10 9 13 3 3 0 2
34 1 10 0 9 1 10 9 4 13 16 2 3 2 10 9 1 9 13 1 13 15 3 16 10 9 0 13 9 1 10 0 9 0 2
29 10 9 0 13 1 9 1 9 2 7 15 1 15 13 1 9 0 13 15 13 1 10 9 1 13 10 10 9 2
25 1 9 2 10 9 4 13 16 10 9 13 9 1 13 10 9 9 0 1 13 13 10 9 0 2
42 10 9 13 3 0 9 1 10 9 1 10 9 7 1 10 9 1 10 9 1 1 10 9 2 10 15 13 0 13 0 9 1 10 9 0 7 0 10 9 9 13 2
25 10 9 4 13 3 1 10 9 16 10 9 13 1 9 10 9 0 15 3 13 15 1 13 9 2
48 3 2 10 0 9 3 13 3 10 9 7 10 9 1 10 9 2 7 13 3 9 0 1 13 10 9 15 13 10 9 1 9 16 10 9 1 10 9 0 13 1 9 1 10 10 9 0 2
46 1 10 9 2 15 4 13 4 13 1 10 9 0 16 13 10 10 9 3 0 1 10 9 0 2 7 13 15 1 13 10 10 9 1 9 1 15 10 9 13 1 10 9 1 9 2
37 1 0 9 2 4 3 4 13 13 10 9 1 10 9 1 10 9 2 7 13 9 1 9 1 10 9 1 13 15 1 13 1 10 9 10 9 2
33 1 0 9 2 4 3 13 10 9 1 9 0 1 10 9 2 1 9 10 16 10 9 0 4 13 1 13 10 9 1 10 9 2
30 1 10 9 2 10 9 13 3 16 10 11 11 0 13 1 10 9 0 10 9 15 13 2 7 15 1 9 0 0 2
33 1 9 2 10 9 1 10 10 11 15 13 1 11 2 1 10 11 11 2 1 13 10 9 1 10 9 0 1 10 0 12 9 2
35 16 10 9 13 10 9 1 10 9 1 10 9 0 0 7 10 9 1 10 9 0 2 10 11 11 4 13 10 9 1 10 9 1 11 2
5 9 1 11 11 2
5 9 12 2 12 2
6 10 9 1 13 0 2
35 11 2 11 2 10 11 11 11 13 10 9 3 0 2 1 9 1 0 9 1 13 10 0 9 1 9 0 7 9 3 3 1 10 9 2
18 15 13 3 10 0 9 1 4 13 1 10 9 1 15 1 3 0 2
30 3 1 10 11 2 3 13 0 16 13 10 9 0 3 3 0 1 13 10 9 1 10 11 11 1 13 10 0 9 2
47 10 9 0 4 13 15 10 9 2 3 16 1 10 9 3 3 0 2 10 15 4 13 3 2 16 15 1 10 9 0 3 13 10 9 1 10 9 1 10 9 3 0 1 15 3 0 2
33 1 10 12 1 10 12 2 4 13 0 13 10 9 0 0 2 1 0 9 16 10 10 9 13 4 13 1 9 0 1 0 9 2
31 1 10 9 1 10 11 1 10 12 2 15 1 10 0 9 4 13 1 9 2 3 3 0 2 7 3 3 0 1 13 2
29 10 11 3 13 9 1 0 9 1 10 11 11 7 1 10 0 0 9 2 1 16 15 4 13 10 9 0 0 2
52 10 0 9 1 10 9 13 1 15 4 4 13 1 10 9 12 2 16 10 9 0 1 0 11 11 11 4 4 13 1 13 15 2 1 10 9 1 9 0 1 10 9 1 10 9 1 10 9 1 11 11 2
42 1 3 2 15 15 15 4 13 2 11 11 2 4 13 1 13 10 9 1 10 9 2 7 1 13 10 9 0 1 10 10 9 7 9 1 10 0 7 0 9 0 2
39 2 16 4 13 1 10 11 1 10 9 12 2 10 9 1 10 10 9 1 10 0 9 1 10 9 3 0 4 3 13 0 1 10 9 1 0 9 2 2
22 3 2 10 11 13 0 9 1 10 9 15 13 9 2 1 10 11 1 10 0 9 2
18 7 1 10 9 1 10 9 1 10 11 11 2 10 9 15 13 9 2
16 1 10 9 3 0 1 11 2 15 13 3 3 3 10 9 2
39 13 16 1 10 9 1 10 9 1 9 1 10 9 1 9 13 0 10 9 1 10 9 2 1 3 13 1 10 9 1 9 1 10 9 1 10 11 11 2
23 1 9 15 13 7 13 0 10 9 1 10 11 11 2 1 9 1 10 10 10 0 9 2
39 15 15 13 4 13 10 0 9 13 1 10 9 1 11 11 2 13 1 10 9 1 10 9 1 9 1 10 9 13 1 0 9 1 9 2 9 7 9 2
5 10 0 9 13 2
23 2 10 11 4 3 13 10 9 0 1 13 10 9 0 1 10 11 11 1 9 0 2 2
19 10 11 11 3 13 15 15 13 1 10 11 2 7 3 13 10 9 0 2
53 13 10 9 1 10 9 1 13 1 13 10 11 1 10 0 9 0 2 3 10 9 0 13 3 3 13 1 10 10 9 0 7 1 9 1 9 1 9 2 7 3 1 10 9 1 10 9 1 10 9 0 2 2
36 1 10 0 9 2 15 1 10 0 9 4 13 15 1 13 10 9 1 9 1 10 11 3 3 1 10 11 2 1 10 9 13 1 10 9 2
23 1 10 0 9 1 10 9 1 9 0 2 10 9 3 13 0 2 7 15 13 1 13 2
28 2 1 10 9 0 2 15 13 10 0 9 1 11 11 11 2 10 10 9 1 10 11 11 1 11 11 2 2
26 10 9 4 4 13 2 1 9 0 2 1 9 1 10 9 1 10 11 11 3 16 4 13 1 9 2
46 1 10 9 2 1 10 12 7 1 10 9 1 10 12 10 9 1 10 9 11 11 3 4 13 10 9 1 9 2 7 10 9 1 9 1 0 9 1 10 11 4 3 13 1 13 2
31 10 9 11 4 13 1 13 10 9 1 10 11 1 10 9 2 3 0 2 1 9 1 10 9 1 10 9 1 10 11 2
15 15 13 10 0 9 0 2 7 3 13 0 1 9 0 2
23 7 10 9 3 0 13 16 10 11 3 13 3 9 1 10 9 0 1 9 1 10 11 2
62 15 1 15 13 9 10 11 13 10 0 9 1 10 9 2 3 1 1 10 0 9 2 1 10 9 2 1 10 9 15 4 13 1 9 10 9 1 10 9 2 10 9 15 1 10 9 1 10 0 12 9 4 13 10 9 1 10 9 7 10 9 2
11 10 9 1 10 11 13 0 7 4 13 2
31 10 9 3 13 9 1 10 10 0 9 1 9 2 7 10 9 7 10 9 1 10 9 1 0 7 0 9 4 4 13 2
21 13 0 16 10 9 11 13 10 9 1 10 9 1 9 3 0 7 1 0 9 2
12 7 10 9 0 1 10 11 13 10 9 0 2
5 9 12 2 12 2
6 11 7 10 11 0 2
31 11 2 1 10 10 9 2 10 9 11 11 4 13 16 15 13 2 1 10 9 2 12 9 0 1 10 9 0 1 11 2
51 3 2 10 9 1 15 10 9 1 10 9 7 10 9 1 10 9 4 13 1 10 9 1 10 9 1 10 9 9 1 10 9 1 10 9 1 9 7 1 10 0 9 1 10 9 1 9 1 10 9 2
50 1 0 9 2 10 9 1 11 1 13 16 10 9 1 10 9 1 9 1 9 0 7 0 1 10 9 0 4 13 1 0 9 1 10 9 1 10 9 1 9 2 13 1 10 9 0 1 10 9 2
19 1 0 9 2 10 9 1 11 1 10 9 1 10 9 1 10 9 9 2
14 7 10 0 7 10 0 9 13 10 0 9 1 9 2
45 7 2 16 10 9 1 11 1 15 10 9 7 10 9 9 4 13 9 0 7 3 0 4 3 0 1 10 10 9 7 1 10 9 1 10 9 0 2 3 4 3 13 3 0 2
12 13 10 9 1 10 9 1 10 9 15 13 2
15 10 9 0 13 12 9 0 0 1 10 9 1 10 9 2
8 13 10 9 1 10 9 0 2
12 13 3 10 9 1 10 9 1 10 9 0 2
30 13 10 9 2 10 9 2 10 9 2 10 9 7 10 9 1 13 16 10 9 7 10 9 1 9 13 10 9 13 2
24 13 15 1 9 1 9 0 7 1 10 9 1 13 1 9 16 10 10 9 13 10 0 9 2
25 13 9 0 2 1 9 10 9 2 15 13 9 0 2 0 7 1 9 2 7 15 4 4 13 2
39 10 0 12 9 13 10 9 0 1 15 15 13 3 2 9 2 2 16 10 9 1 10 15 7 1 10 0 9 15 13 1 15 15 13 1 2 9 2 2
48 10 11 0 2 7 10 9 1 10 9 1 9 1 10 9 1 9 7 10 9 1 10 9 1 10 9 1 10 9 2 4 13 3 10 9 1 13 1 10 9 7 1 10 9 1 10 9 2
49 7 2 1 0 9 2 4 13 1 9 0 10 9 1 10 9 2 1 10 9 2 1 10 9 2 1 10 9 7 1 10 9 1 10 9 7 1 10 9 1 10 9 7 1 15 1 10 9 2
72 1 10 13 10 9 2 10 9 0 1 10 9 4 13 1 13 2 16 10 9 0 1 10 9 1 9 0 2 0 1 13 13 10 9 1 10 9 0 2 3 4 13 1 3 10 9 1 9 13 1 13 1 10 9 0 15 13 9 1 10 9 1 9 2 9 7 9 1 3 12 9 2
43 3 15 13 2 3 2 10 9 1 9 1 10 9 15 13 10 9 13 1 10 9 1 10 9 7 1 10 9 1 13 3 3 1 10 9 1 10 0 7 1 10 9 2
54 3 2 10 9 1 10 9 0 13 1 10 9 1 10 9 0 1 10 9 1 0 9 1 10 9 1 9 1 10 9 7 1 10 9 1 9 2 7 1 10 9 1 10 9 1 10 9 7 1 15 1 10 9 2
29 15 1 15 4 4 13 1 10 9 1 10 9 0 7 16 15 4 13 9 0 1 10 9 2 1 9 0 2 2
48 10 9 0 15 13 1 10 9 16 15 15 2 1 15 2 15 13 1 13 10 0 9 1 9 0 1 10 9 2 9 1 10 9 0 7 1 10 9 1 9 2 13 3 1 9 1 9 2
29 11 13 3 1 13 10 9 16 10 9 1 10 9 0 1 10 9 0 4 13 10 9 1 10 9 1 10 9 2
38 3 2 10 9 1 10 9 3 4 4 13 1 10 9 10 1 13 10 15 15 4 13 10 9 1 9 2 9 1 10 9 7 9 1 9 2 0 2
16 1 9 4 4 13 15 2 7 10 9 1 11 13 0 9 2
44 10 9 3 2 10 9 0 11 2 11 7 11 3 13 1 13 16 10 9 1 10 9 9 0 13 1 10 9 4 13 1 10 1 3 1 10 12 5 1 13 10 9 0 2
39 3 2 1 10 9 13 1 9 2 9 0 2 9 0 7 1 9 2 10 9 1 10 9 0 7 1 10 9 4 13 1 10 9 15 15 13 10 0 2
20 3 2 10 9 1 10 9 1 9 3 4 4 13 15 16 13 9 7 9 2
55 7 11 7 10 9 4 4 13 10 9 3 13 15 4 13 10 9 13 10 9 1 13 10 12 5 1 10 9 9 1 10 9 7 10 0 12 5 1 10 9 1 9 7 1 10 9 1 9 1 10 9 7 10 9 2
58 3 2 10 9 0 13 16 15 13 10 9 1 9 13 1 13 1 10 9 1 13 13 1 10 15 1 13 10 10 9 3 0 7 0 2 7 16 10 9 1 10 9 13 10 9 1 9 1 9 1 10 9 13 15 1 9 0 2
24 7 13 10 0 9 1 10 9 1 10 9 7 1 10 9 2 3 10 9 0 13 10 9 2
43 1 10 9 2 10 9 1 10 0 9 13 1 13 0 1 10 9 0 7 3 0 2 16 10 0 9 2 13 15 1 10 9 0 7 1 10 9 2 13 1 4 13 2
33 0 3 1 10 9 0 1 10 9 15 13 10 9 2 1 10 9 1 10 15 15 1 15 4 13 1 10 9 7 1 10 9 2
16 10 9 1 9 1 9 1 10 0 9 1 11 2 1 3 2
5 9 1 11 11 2
5 11 12 2 12 2
5 10 9 1 11 2
44 11 2 10 9 1 9 13 1 10 9 1 9 1 10 9 1 10 12 7 10 9 0 1 10 11 7 1 10 11 1 10 9 1 10 12 4 3 13 10 2 9 13 2 2
38 1 16 10 11 4 13 7 13 10 11 2 7 4 13 1 13 9 7 13 9 1 10 10 9 0 2 15 1 11 4 13 1 10 2 9 13 2 2
26 3 15 13 15 1 13 2 3 2 1 10 9 13 1 15 0 1 13 10 10 9 7 10 10 9 2
24 10 9 7 10 9 1 10 10 9 15 4 13 1 0 1 10 9 0 1 3 4 13 3 2
37 10 10 9 4 13 10 9 1 10 9 1 9 1 10 9 0 0 15 15 13 15 1 10 9 1 15 13 9 1 13 10 10 9 0 7 0 2
25 10 9 13 10 0 9 0 2 7 10 9 4 13 1 13 15 10 9 3 1 13 10 10 9 2
53 1 10 9 1 9 2 10 9 1 15 15 2 1 10 9 1 11 2 13 16 10 9 1 10 9 3 4 3 4 13 1 0 1 10 9 2 4 13 10 9 1 10 9 2 1 10 9 0 1 10 10 9 2
11 3 13 3 10 9 1 10 9 0 0 2
26 7 10 9 0 13 16 2 16 10 11 13 10 10 9 1 1 15 2 15 4 13 1 10 9 0 2
45 10 0 9 1 10 9 0 11 11 1 10 9 0 11 11 1 13 10 9 0 2 13 1 10 9 0 1 16 13 10 9 1 9 1 10 11 2 13 1 9 0 1 10 9 2
45 10 9 1 11 13 0 1 10 0 9 1 11 1 10 12 2 3 11 11 13 11 11 7 11 11 11 9 1 10 9 1 10 11 15 4 13 9 1 10 9 1 3 12 9 2
48 3 11 4 13 1 13 10 9 9 1 10 9 1 10 11 13 10 9 0 13 1 10 11 1 9 1 13 10 9 1 11 2 0 9 1 9 15 10 11 4 13 3 3 1 10 0 9 2
8 10 9 4 13 10 0 9 2
19 13 10 9 0 3 16 3 13 10 9 13 3 13 2 7 1 9 0 2
16 7 10 9 1 10 9 0 3 13 15 15 13 1 9 11 2
38 1 10 9 2 10 9 0 13 10 9 13 1 9 1 10 11 1 13 9 0 7 1 10 9 13 10 9 0 7 0 1 10 11 1 10 9 0 2
16 1 13 11 2 10 9 1 11 13 10 9 13 1 0 9 2
12 13 13 10 9 13 1 0 1 10 9 0 2
27 10 0 9 0 1 10 11 13 10 9 1 13 1 9 1 10 2 9 1 10 9 0 1 10 11 2 2
27 10 9 13 1 11 1 13 1 13 7 13 10 9 1 9 0 1 13 15 1 10 9 0 1 10 9 2
17 10 9 0 1 10 11 4 4 13 3 1 10 9 1 10 11 2
26 10 11 3 4 13 9 1 9 2 7 4 13 15 1 9 0 9 2 1 15 0 13 10 10 9 2
34 10 11 3 13 10 11 2 3 10 9 4 13 1 9 1 9 15 13 9 1 9 1 0 9 1 10 9 1 10 9 1 10 11 2
22 7 3 13 10 11 2 15 13 0 1 10 0 9 1 15 4 13 10 10 9 0 2
19 10 11 13 10 9 3 0 2 13 1 0 1 10 9 2 13 10 11 2
40 13 9 1 10 9 0 1 11 13 13 10 9 15 10 11 13 1 13 1 10 0 9 1 9 1 10 11 7 1 10 9 7 10 9 0 15 4 13 11 2
34 10 9 1 11 13 16 10 9 1 9 0 15 13 1 11 13 1 9 2 7 3 13 1 13 10 0 9 1 9 15 4 13 15 2
38 10 9 1 9 0 13 1 10 11 0 7 1 10 11 4 13 1 11 2 7 10 9 1 9 0 4 13 9 0 3 1 10 1 3 1 10 9 2
5 10 9 13 0 2
21 3 15 13 10 9 1 10 9 1 9 0 1 11 2 7 3 15 4 3 13 2
14 10 9 1 10 11 1 11 13 0 2 0 7 0 2
6 7 13 10 0 9 2
18 3 10 11 4 4 13 1 13 10 0 9 0 0 1 10 0 9 2
15 15 1 15 13 9 13 10 9 0 2 0 7 3 0 2
17 7 2 1 10 9 7 10 9 0 1 10 11 2 15 13 15 2
19 10 9 1 10 9 1 13 10 9 0 1 10 9 1 10 11 13 0 2
22 7 10 9 13 1 10 11 2 16 13 1 10 9 2 13 3 10 9 1 10 11 2
42 7 9 0 2 13 10 9 1 10 11 13 10 9 16 10 9 0 4 13 10 9 15 15 13 3 1 13 1 10 10 9 2 1 1 13 15 13 1 10 10 9 2
13 10 11 13 1 10 9 2 1 0 2 16 0 2
15 15 13 1 13 1 10 9 0 1 10 0 9 1 9 2
5 11 12 2 12 2
6 10 9 1 10 9 2
23 11 2 10 9 10 9 13 1 10 9 13 9 1 9 7 13 9 1 9 1 15 10 2
21 1 10 12 4 4 13 12 9 1 9 1 9 15 4 3 13 1 12 12 9 2
32 10 9 9 13 15 1 10 0 9 1 9 7 9 1 10 9 0 7 0 7 13 3 12 9 10 9 15 4 13 10 9 2
32 1 10 9 1 10 9 13 7 0 2 13 10 0 9 1 10 9 0 2 7 10 9 15 13 7 15 13 1 10 9 0 2
55 13 16 3 13 0 7 9 1 9 1 10 9 9 7 10 9 1 10 11 0 2 7 13 3 16 13 0 13 1 10 9 1 9 1 10 9 1 10 9 1 9 2 13 3 0 10 9 3 0 1 9 1 10 9 2
18 10 0 9 13 16 15 13 10 0 9 0 1 4 13 1 10 9 2
11 13 3 1 10 9 0 13 15 15 9 2
53 3 2 10 9 0 13 1 10 9 1 10 9 2 10 0 2 9 1 9 1 10 9 2 2 11 2 2 15 13 1 10 9 1 9 1 10 9 1 10 9 9 15 4 3 13 1 10 9 13 1 10 9 2
31 7 10 9 2 15 4 13 1 1 10 9 1 10 9 0 2 3 4 13 10 9 1 10 9 1 9 1 10 10 9 2
20 10 0 9 1 10 9 1 10 9 0 13 10 9 0 2 7 3 3 0 2
33 1 10 9 1 9 0 13 1 10 9 0 2 10 9 0 11 4 13 10 0 9 1 13 10 9 1 9 15 13 10 9 9 2
40 10 9 9 4 13 1 10 9 1 10 9 0 1 15 13 10 9 1 0 9 1 10 9 15 13 10 9 0 1 10 9 13 15 13 3 16 13 10 9 2
31 10 9 9 3 13 7 3 13 10 9 1 10 9 7 13 16 10 10 9 13 10 9 3 13 13 1 13 1 10 9 2
28 16 10 9 9 4 13 1 10 9 1 10 9 2 15 4 1 9 13 1 10 9 0 1 10 9 1 9 2
12 3 13 1 13 16 10 9 13 1 10 9 2
51 10 9 0 13 1 10 9 1 9 1 10 9 0 13 7 10 9 11 4 13 13 1 9 3 0 1 10 9 3 0 2 7 1 10 9 2 1 9 0 1 10 9 1 9 13 1 15 13 10 9 2
38 3 16 10 11 4 13 10 9 1 10 9 1 10 11 11 2 1 11 7 1 11 2 15 4 3 13 1 13 10 9 1 0 9 13 10 11 11 2
28 10 9 4 3 3 13 7 13 1 13 10 9 7 10 9 2 1 10 9 3 1 10 9 0 1 0 9 2
25 1 10 9 1 13 10 9 0 1 9 2 10 9 0 4 13 10 9 1 10 9 1 9 0 2
25 10 9 13 16 10 9 0 0 13 3 3 0 7 0 1 10 9 0 7 3 0 1 10 9 2
68 7 2 16 1 10 9 10 9 11 13 1 3 4 13 1 10 9 1 0 9 1 10 9 2 1 10 15 10 9 0 1 10 9 13 3 13 13 1 4 13 7 0 1 10 10 9 2 16 10 9 13 2 7 13 1 9 3 1 13 2 10 9 1 9 1 10 9 2
24 1 9 2 10 9 7 10 9 1 10 9 0 13 3 0 2 13 10 9 7 13 10 9 2
23 7 10 15 13 3 3 0 1 10 9 1 10 9 1 10 9 13 10 9 1 10 9 2
74 10 9 0 1 10 9 7 10 9 1 10 9 0 1 10 9 0 1 10 9 4 13 10 9 1 10 9 1 9 16 13 2 10 9 13 1 9 0 2 9 1 9 2 1 10 0 9 1 9 1 10 9 2 2 1 1 13 15 3 2 10 9 0 15 13 1 9 1 13 10 9 0 2 2
31 1 0 9 2 10 9 1 9 4 13 10 9 7 10 9 0 1 10 9 15 10 9 4 13 7 13 10 9 1 9 2
54 13 10 9 1 9 13 1 10 9 13 1 10 9 2 10 9 0 3 4 13 10 9 1 10 9 0 1 13 15 2 1 10 0 1 10 9 0 0 7 9 15 4 1 9 13 10 9 1 10 9 0 3 13 2
5 9 1 11 11 2
5 11 12 2 12 2
7 10 0 9 1 10 11 2
62 11 2 1 10 0 9 1 10 9 1 10 9 0 11 11 2 2 10 9 1 10 9 11 4 13 1 10 9 0 2 2 10 9 1 13 15 0 9 16 3 10 9 1 10 11 13 13 10 10 9 0 1 3 15 4 13 1 10 0 9 0 2
12 10 10 9 4 3 13 1 10 0 9 0 2
26 7 13 3 10 9 1 13 10 9 13 1 10 11 16 13 1 9 3 0 1 10 9 1 10 9 2
22 11 13 1 0 9 1 10 9 1 10 11 1 13 10 11 1 4 15 13 10 9 2
48 1 10 9 2 4 13 1 13 10 9 1 10 9 1 13 10 2 9 0 2 0 15 13 10 9 1 13 0 0 13 7 13 10 9 0 1 10 9 9 16 3 13 0 1 10 9 13 2
19 1 10 9 2 10 9 4 13 3 1 10 9 1 10 9 0 1 9 2
24 3 16 4 13 0 2 10 9 1 11 13 2 1 10 0 1 10 9 2 10 9 3 0 2
27 3 1 13 2 10 9 0 13 0 7 1 10 9 1 9 2 3 1 15 1 10 0 9 1 10 11 2
35 1 10 0 9 2 16 10 9 9 13 10 9 0 2 3 10 0 9 1 13 1 9 10 9 15 13 10 9 1 9 0 4 13 15 2
28 1 10 0 12 9 2 10 9 1 13 10 9 11 0 4 13 1 10 9 1 10 9 15 13 13 10 9 2
26 3 2 16 10 9 13 1 0 1 9 2 13 9 1 13 1 13 10 9 1 10 9 0 1 9 2
19 3 2 1 10 9 1 10 11 4 13 2 3 3 10 9 13 16 13 2
45 1 13 10 9 2 10 9 1 9 0 2 13 3 1 10 11 11 7 1 10 9 0 0 2 4 13 10 9 0 16 4 13 10 9 1 10 9 3 0 7 13 10 0 9 2
25 15 2 1 9 2 4 13 10 9 1 10 9 0 7 13 10 9 1 10 9 1 10 9 0 2
25 7 11 2 15 1 15 13 13 3 10 9 2 13 10 11 1 10 9 1 10 3 3 0 11 2
7 10 11 13 1 0 9 2
36 13 10 9 1 10 9 7 1 10 9 0 0 7 13 1 9 0 1 13 10 9 1 9 2 10 9 13 4 13 10 11 1 10 9 0 2
22 1 0 9 2 10 11 3 4 0 1 13 10 9 1 10 10 9 1 13 10 11 2
15 1 3 2 10 0 9 0 13 3 3 3 1 10 9 2
42 10 9 0 1 10 9 4 13 1 3 10 12 5 1 10 12 7 1 10 12 9 1 10 9 0 3 1 0 9 15 1 10 9 13 10 9 1 9 7 9 0 2
35 3 3 2 3 2 10 9 1 10 9 0 4 13 2 15 1 10 9 0 4 13 10 15 2 13 1 10 1 3 1 10 12 5 0 2
29 1 9 15 13 10 0 9 2 7 10 9 1 10 9 0 13 16 10 9 1 9 0 1 10 0 9 13 0 2
39 10 12 0 9 1 10 9 2 10 0 7 0 2 4 13 10 9 0 1 10 11 1 10 9 1 10 9 1 10 12 15 4 13 10 10 9 1 9 2
36 3 3 9 13 10 9 1 11 1 10 9 11 2 15 13 1 10 9 0 0 1 13 9 0 1 9 1 10 9 3 0 1 10 9 2 2
75 16 10 11 0 15 13 3 2 7 3 2 1 10 9 16 3 13 1 10 9 1 10 9 2 3 1 10 9 1 9 2 13 3 9 1 10 9 0 0 2 10 9 4 4 13 1 10 9 16 10 9 0 0 2 1 10 13 10 9 1 10 9 2 4 13 10 9 13 1 10 9 1 9 0 2
23 10 11 13 10 9 0 13 15 13 1 13 10 9 1 10 9 2 9 1 10 0 9 2
17 7 10 9 1 10 9 0 3 4 13 1 13 1 10 0 9 2
24 10 9 4 13 10 3 0 1 10 9 2 10 9 1 0 9 0 7 1 10 3 13 9 2
21 13 15 4 13 10 9 1 9 0 2 10 10 9 4 13 3 1 10 9 0 2
31 3 2 10 9 1 10 11 13 1 9 2 13 10 0 9 0 10 9 1 10 9 1 9 1 9 0 15 3 4 13 2
40 7 10 9 7 10 9 1 10 9 1 9 4 13 1 9 10 9 0 1 10 9 2 10 9 15 10 0 9 1 10 9 0 4 3 13 1 10 0 9 2
16 3 2 10 9 0 13 1 13 10 9 13 3 0 16 3 2
49 13 9 1 10 9 1 10 9 0 1 13 10 9 0 13 3 0 2 7 13 1 9 1 10 9 2 3 16 1 13 15 13 10 9 1 10 9 0 2 13 1 3 15 1 10 0 9 0 2
31 10 9 1 10 9 4 13 10 9 2 7 3 10 9 4 13 7 13 3 10 9 0 3 13 16 13 10 9 3 0 2
49 13 10 9 9 0 1 13 1 10 10 9 2 10 0 9 1 10 11 13 15 1 13 15 1 10 9 1 10 9 13 7 13 16 10 9 7 10 9 13 10 10 9 2 7 13 1 15 13 2
13 13 1 10 9 3 0 13 1 10 0 9 0 2
5 9 1 11 11 2
