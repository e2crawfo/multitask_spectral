727 11
6 13 4 12 9 13 2
7 9 3 13 15 13 9 2
7 9 13 15 1 0 9 2
8 13 9 7 13 15 13 9 2
4 0 9 13 2
12 2 14 13 2 3 12 9 13 3 1 15 2
36 9 0 0 9 0 13 0 9 9 1 13 8 2 9 2 9 7 13 9 7 9 1 0 13 9 1 9 0 2 0 15 13 9 9 0 2
4 2 13 9 2
5 9 13 1 9 2
25 14 13 13 0 9 7 14 13 1 15 13 1 9 1 9 9 2 16 9 4 13 14 1 15 2
4 14 13 15 2
19 2 12 9 13 4 1 9 2 16 13 9 1 0 9 2 1 0 9 2
3 14 13 2
8 13 15 2 3 13 0 9 2
10 2 12 0 9 13 2 16 4 13 2
10 9 0 9 1 9 13 9 1 0 2
9 3 13 0 9 9 7 15 9 2
9 15 9 9 14 13 16 0 9 2
9 14 1 13 14 13 15 0 9 2
30 9 13 2 16 1 0 9 13 3 14 12 9 0 7 9 1 0 9 2 0 9 13 1 9 9 13 1 13 9 2
18 2 13 0 14 0 9 0 2 0 13 1 9 1 9 1 0 9 2
4 9 13 4 2
8 2 0 9 13 3 0 9 2
11 0 9 2 13 1 9 2 13 1 9 2
37 9 2 0 9 9 0 7 9 9 9 2 7 9 2 0 9 0 9 9 2 13 15 9 9 2 4 14 13 1 13 9 7 9 8 2 9 2
10 1 0 8 2 4 1 0 9 13 2
10 14 13 4 2 16 0 9 13 3 2
23 1 9 13 2 16 13 4 15 14 1 9 13 2 16 13 1 9 9 1 9 2 2 2
18 9 13 2 16 1 9 9 9 0 9 9 0 13 9 0 7 9 2
13 3 13 9 9 2 0 9 13 0 9 9 9 2
14 13 12 9 2 1 0 13 9 0 13 1 15 0 2
13 13 9 9 0 9 0 9 7 0 9 0 8 2
11 9 13 13 1 9 1 9 9 0 9 2
13 3 9 9 9 13 0 9 1 9 9 9 9 2
9 9 13 9 9 7 9 0 9 2
18 9 9 9 0 1 9 7 9 9 13 15 1 9 9 9 9 9 2
4 9 9 13 2
7 3 7 3 9 14 13 2
10 3 3 14 13 0 9 1 9 9 2
10 9 0 3 13 15 2 14 3 13 2
17 14 13 9 9 2 13 2 16 9 0 13 13 15 3 0 9 2
6 14 4 13 0 9 2
7 13 13 15 15 0 9 2
9 14 9 1 0 9 3 13 0 2
6 13 14 9 0 9 2
23 13 14 13 2 16 1 0 9 0 9 14 1 9 14 13 2 0 1 9 14 15 13 2
13 14 9 1 9 13 14 3 13 1 3 0 9 2
8 9 13 0 9 1 9 0 2
12 9 1 13 9 9 1 0 9 13 9 9 2
14 9 9 9 13 1 15 9 1 13 1 9 9 9 2
13 13 15 9 1 9 9 9 2 0 1 9 0 2
12 14 1 9 0 9 13 15 15 13 0 9 2
5 1 0 9 13 2
18 12 9 13 1 9 9 9 9 2 13 13 9 2 13 9 7 9 2
14 9 12 2 0 9 0 9 2 4 13 1 0 8 2
23 9 2 16 4 13 1 0 9 2 14 4 13 9 9 2 16 14 13 15 9 9 0 2
13 13 4 1 15 7 3 13 4 9 1 9 0 2
10 3 13 1 9 9 9 0 1 9 2
12 0 9 13 2 16 1 9 9 13 15 9 2
7 9 13 12 9 1 13 2
10 9 13 1 0 9 14 12 9 9 2
9 0 9 0 9 13 1 9 0 2
12 9 9 13 2 16 1 9 14 13 0 9 2
8 1 15 9 9 13 0 9 2
6 3 13 15 12 8 2
12 1 0 9 9 0 13 0 0 9 15 13 2
12 0 9 13 2 16 9 13 3 0 0 9 2
18 3 7 1 9 0 7 9 9 13 0 9 1 9 2 9 7 9 2
5 9 3 13 9 2
17 9 9 0 4 1 0 9 13 2 7 14 13 13 0 9 0 2
16 16 13 1 9 2 7 9 13 13 0 9 1 0 1 9 2
4 9 13 9 2
3 13 15 2
26 4 9 13 1 9 0 13 9 7 0 9 0 2 4 13 1 14 0 9 13 15 1 9 9 0 2
5 9 13 14 9 2
8 1 9 0 13 9 0 9 2
15 13 4 1 0 9 9 2 16 13 15 13 9 13 9 2
12 1 0 9 13 12 0 9 9 7 12 0 2
5 4 3 13 9 2
5 14 13 9 9 2
5 14 13 9 9 2
9 13 9 2 16 13 9 0 9 2
14 7 9 3 13 15 3 0 7 9 14 13 15 13 2
20 1 9 0 9 13 4 1 9 9 9 0 7 0 2 13 13 9 0 9 2
7 0 1 15 13 9 9 2
18 13 9 1 0 9 9 3 4 13 1 9 1 13 9 1 0 9 2
10 13 0 9 2 16 13 1 14 9 2
8 4 13 0 9 2 0 9 2
9 9 13 3 2 16 14 13 13 2
20 9 7 15 9 13 2 16 13 9 9 2 9 1 9 9 13 15 13 9 2
19 3 13 15 1 0 9 9 1 9 0 2 9 1 9 9 9 13 9 2
13 1 0 9 13 2 16 13 9 9 1 9 9 2
17 13 15 13 2 16 13 1 15 0 9 2 7 1 9 14 13 2
14 0 7 13 15 1 9 2 0 13 9 9 9 9 2
10 9 13 2 16 13 15 13 0 9 2
21 9 13 15 1 9 1 9 7 9 9 13 15 2 16 15 0 0 9 14 13 2
22 0 9 13 1 9 13 1 9 2 16 1 9 1 9 9 14 13 13 15 1 9 2
5 13 1 15 9 2
9 1 9 13 15 0 9 9 9 2
12 3 13 9 9 2 14 13 14 9 1 9 2
3 13 3 2
4 14 13 9 2
13 13 9 1 9 2 1 9 13 13 1 9 9 2
6 14 14 13 1 9 2
12 9 13 2 16 9 2 0 13 2 4 13 2
12 14 3 2 1 12 9 2 9 13 1 9 2
6 9 9 9 13 0 2
7 1 9 9 13 14 13 2
4 13 1 9 2
6 13 14 9 1 9 2
7 12 9 13 3 1 9 2
7 13 15 1 9 1 9 2
10 13 14 2 16 15 3 13 2 2 2
13 3 3 13 15 1 3 13 0 9 1 0 9 2
9 13 0 9 2 14 13 15 3 2
7 12 9 13 15 1 9 2
6 9 13 3 7 13 2
28 9 9 0 9 9 14 13 2 16 0 1 12 9 1 9 9 0 2 0 3 13 9 2 13 1 9 0 2
9 13 12 9 2 1 0 13 9 2
6 9 9 13 3 0 2
5 7 14 4 0 2
6 9 9 13 0 9 2
7 1 9 9 13 14 4 2
14 1 0 9 9 3 13 13 0 9 7 9 15 13 2
13 13 15 9 9 0 1 0 9 7 0 9 0 2
10 1 9 0 9 9 0 13 15 9 2
12 3 13 15 9 0 9 7 13 9 1 9 2
16 3 13 4 9 9 13 13 2 3 9 13 15 3 3 13 2
9 0 9 1 9 1 9 9 13 2
7 9 1 9 13 9 9 2
13 1 9 1 0 9 9 13 14 8 2 12 8 2
7 9 9 0 13 0 9 2
13 1 9 13 15 1 9 7 9 7 13 1 9 2
11 1 9 0 0 9 13 15 13 1 9 2
15 1 0 9 13 1 9 2 7 1 15 9 13 0 9 2
5 3 13 9 9 2
26 13 9 1 0 9 9 13 2 16 9 2 9 2 9 2 0 9 0 13 15 1 9 1 9 0 2
2 13 2
4 14 13 9 2
4 13 15 15 2
11 13 1 0 9 0 9 9 13 1 9 2
4 3 14 13 2
13 1 9 13 9 9 9 9 1 3 13 1 9 2
8 9 0 13 3 13 1 9 2
7 9 9 13 12 9 9 2
19 9 1 9 9 1 9 13 15 3 3 2 7 9 4 0 14 1 9 2
29 9 1 9 9 2 0 13 1 13 9 9 0 9 2 13 0 9 0 9 2 16 13 0 9 1 9 7 9 2
14 2 1 0 9 13 4 0 9 1 13 9 1 9 2
15 0 9 14 13 15 9 2 3 0 2 15 15 9 13 2
8 14 4 3 13 1 9 9 2
6 7 15 14 13 9 2
9 1 9 13 9 3 0 1 9 2
13 1 0 13 15 13 9 2 0 13 15 1 9 2
10 9 9 13 2 16 14 13 15 9 2
17 1 9 1 9 0 7 9 9 9 9 13 15 1 9 1 9 2
14 13 13 2 1 0 9 13 14 0 0 2 0 9 2
7 1 9 13 15 14 9 2
12 14 13 14 2 14 15 0 13 15 1 9 2
9 9 1 12 0 9 13 1 0 2
9 9 14 4 14 13 1 9 0 2
8 1 9 0 13 3 0 9 2
6 13 9 1 9 9 2
5 1 9 13 9 2
6 3 4 4 0 9 2
4 13 1 9 2
3 14 13 2
11 14 0 9 13 15 3 1 9 1 9 2
11 9 9 13 3 1 9 9 9 9 9 2
16 9 13 14 9 0 9 2 13 2 16 13 15 0 9 9 2
17 16 9 9 13 1 9 9 2 7 14 13 14 12 8 1 9 2
9 14 3 9 0 9 13 0 9 2
14 9 3 13 2 16 1 9 13 15 13 14 1 9 2
6 14 2 9 13 0 2
5 14 13 4 9 2
5 13 13 9 9 2
5 13 15 1 9 2
14 1 9 9 9 13 9 9 9 7 9 8 2 9 2
11 13 14 0 9 2 13 1 0 9 9 2
19 9 9 14 13 9 0 1 13 0 2 0 9 9 2 13 1 9 0 2
22 13 2 16 1 0 0 9 2 0 9 2 9 7 13 9 9 0 13 14 3 13 2
4 14 13 15 2
14 3 9 9 9 1 9 13 15 1 0 9 9 0 2
27 9 9 2 0 9 13 9 9 9 2 13 9 9 0 1 0 8 2 7 13 12 0 9 1 0 9 2
8 15 9 4 9 14 1 15 2
5 13 1 9 0 2
14 9 13 9 0 9 2 9 13 2 16 13 13 9 2
3 9 13 2
9 2 9 13 9 1 9 1 9 2
14 3 13 9 2 0 3 13 1 15 9 2 9 9 2
18 0 1 0 9 9 0 9 13 13 0 2 14 0 2 9 9 0 2
14 14 9 9 13 1 9 7 0 9 13 15 0 9 2
4 13 0 9 2
6 0 9 4 0 9 2
14 3 13 1 9 2 13 1 9 1 9 9 1 9 2
14 1 12 9 13 4 14 9 1 9 13 0 9 0 2
10 9 7 9 14 13 1 9 0 9 2
10 7 9 9 1 9 13 9 9 0 2
4 3 15 13 2
11 3 13 9 2 7 13 14 0 9 9 2
12 3 13 9 2 4 3 13 14 1 9 9 2
20 16 1 9 13 9 9 9 7 9 9 9 2 1 9 1 9 15 14 13 2
9 9 13 2 16 0 9 13 0 2
5 14 13 1 9 2
6 14 14 13 4 9 2
7 9 4 3 9 1 9 2
8 13 15 1 9 13 1 9 2
7 13 4 1 9 0 9 2
21 9 9 14 0 15 1 0 9 13 9 1 0 9 2 16 13 4 15 0 9 2
8 0 9 4 3 13 9 9 2
4 13 1 9 2
8 0 3 13 9 13 0 9 2
14 1 9 9 0 9 2 13 15 13 14 1 9 9 2
13 1 9 13 1 0 9 0 9 9 1 9 9 2
11 13 4 0 9 1 9 7 9 1 9 2
8 1 9 9 13 15 14 13 2
12 13 2 16 9 9 9 14 3 15 14 13 2
6 14 13 15 14 15 2
11 1 9 13 9 9 2 13 13 12 9 2
7 1 9 1 9 14 13 2
22 3 2 9 0 9 0 8 2 0 9 0 13 9 9 9 0 1 9 12 9 9 2
12 1 9 0 13 9 0 9 9 0 0 9 2
14 1 15 9 0 9 13 15 9 13 13 3 9 0 2
20 16 13 13 1 9 0 9 1 9 7 9 2 1 0 9 9 13 13 12 2
4 0 13 3 2
6 13 9 0 9 0 2
14 9 3 13 14 0 7 13 14 13 1 9 0 9 2
8 9 14 13 15 9 1 9 2
7 7 9 14 13 1 9 2
24 9 9 14 13 2 16 9 3 13 9 3 13 1 0 9 7 9 14 13 1 9 0 9 2
9 1 9 13 1 0 9 1 9 2
10 1 9 9 13 1 9 1 9 0 2
8 14 13 2 9 13 9 9 2
3 14 13 2
17 1 3 13 9 9 13 1 9 0 2 12 9 1 9 1 9 2
6 1 9 13 1 9 2
15 9 0 0 13 13 1 9 0 2 1 0 13 9 9 2
4 9 13 0 2
14 9 9 13 1 9 9 7 1 9 13 13 9 9 2
16 1 9 0 9 9 9 13 9 9 9 1 13 9 9 0 2
8 9 9 13 13 9 13 9 2
5 7 13 14 0 2
9 13 9 3 13 9 7 13 9 2
13 3 14 13 2 16 13 4 15 1 9 1 15 2
13 7 1 9 13 2 13 9 7 13 15 1 9 2
10 13 9 2 14 15 9 1 9 13 2
3 7 13 2
9 16 15 3 3 1 9 14 13 2
6 13 14 9 7 9 2
17 7 13 4 14 3 13 2 16 9 14 13 1 15 7 13 15 2
9 7 3 9 9 13 1 15 9 2
11 9 9 1 9 0 9 13 3 3 9 2
7 13 1 0 0 9 9 2
4 13 13 9 2
9 13 14 9 9 0 9 7 9 2
19 13 3 9 0 3 3 9 2 1 0 13 15 8 0 1 0 9 9 2
7 13 3 2 16 14 13 2
9 13 3 2 16 0 15 14 13 2
6 13 14 9 9 9 2
11 13 1 15 9 2 9 2 9 9 9 2
8 13 0 0 9 1 9 9 2
3 13 15 2
19 14 13 14 2 16 9 3 13 15 9 9 2 13 0 9 13 9 9 2
6 13 9 9 13 9 2
19 1 9 1 9 9 7 9 13 4 9 1 0 9 2 13 1 9 9 2
15 1 9 1 9 9 9 13 9 1 0 9 1 9 0 2
18 9 9 2 9 14 13 1 9 9 0 9 0 2 13 14 9 13 2
15 3 14 13 14 2 0 9 9 13 1 15 9 9 9 2
10 13 15 15 1 9 0 0 9 0 2
7 15 13 13 1 9 0 2
6 3 0 9 4 13 2
12 0 9 13 15 1 9 9 14 1 9 9 2
16 9 1 9 9 1 0 9 9 13 0 9 2 13 12 9 2
13 9 13 15 2 3 13 9 9 13 1 0 9 2
11 9 13 9 9 1 9 8 2 12 8 2
7 1 9 13 9 1 9 2
23 1 9 1 9 3 13 9 9 9 0 9 0 1 9 0 7 1 9 9 9 4 13 2
17 1 9 1 9 0 9 13 13 9 9 1 9 2 0 13 9 2
16 3 13 4 2 16 3 13 1 9 7 13 1 9 9 9 2
8 13 4 1 15 9 1 9 2
14 13 4 2 3 3 15 13 2 14 13 15 13 9 2
13 13 4 1 0 9 2 0 13 0 2 0 9 2
13 13 4 15 9 1 15 9 7 13 15 0 9 2
10 1 9 9 13 4 15 2 16 13 2
18 13 4 2 16 9 14 13 9 2 7 14 13 4 15 1 9 9 2
11 13 15 15 2 16 13 1 9 0 9 2
13 7 3 13 15 9 0 2 3 13 4 1 15 2
11 15 13 2 7 1 9 13 4 14 12 2
17 13 4 0 0 9 7 13 4 15 2 16 15 15 13 1 9 2
12 1 9 13 0 9 2 9 13 15 1 9 2
6 13 4 15 13 9 2
10 13 14 3 2 3 13 4 0 9 2
11 13 15 1 9 2 16 15 1 15 13 2
7 13 1 9 2 1 9 2
6 13 2 3 13 0 2
4 13 3 9 2
22 3 14 13 0 2 7 3 14 15 14 13 2 9 15 15 13 2 9 13 1 9 2
11 3 13 4 15 2 3 3 15 3 13 2
2 13 2
11 3 13 4 1 9 2 9 13 1 9 2
6 13 15 1 0 9 2
15 14 1 0 9 9 13 4 2 16 4 13 9 13 3 2
7 3 13 14 9 14 13 2
16 9 9 13 1 9 7 13 2 16 3 14 13 3 13 9 2
5 13 3 0 9 2
3 9 13 2
7 13 15 13 2 16 13 2
6 9 9 13 1 9 2
7 13 13 1 13 9 9 2
7 9 0 4 13 1 9 2
6 7 14 9 3 13 2
13 7 14 13 4 2 16 14 3 13 15 0 9 2
9 12 9 1 13 1 9 9 9 2
6 0 9 9 13 9 2
8 3 13 9 1 0 0 9 2
12 9 9 13 9 2 0 9 2 9 2 9 2
6 9 9 13 15 9 2
3 13 0 2
5 14 13 12 9 2
4 9 15 13 2
7 9 3 4 13 1 9 2
5 9 13 9 9 2
14 1 0 9 2 3 3 2 13 12 9 13 1 9 2
6 13 2 3 15 13 2
7 1 9 9 13 9 0 2
8 0 9 4 13 1 0 9 2
12 1 9 9 13 1 9 2 13 3 1 9 2
5 13 15 1 9 2
4 7 9 13 2
5 9 14 13 13 2
25 9 13 9 0 9 1 9 7 13 1 0 9 9 13 9 2 13 0 9 9 2 9 9 0 2
5 3 14 13 4 2
9 1 0 9 13 1 9 1 9 2
13 0 9 13 2 7 12 3 13 15 9 0 9 2
12 0 9 3 13 1 9 9 7 15 9 0 2
6 0 9 13 15 13 2
9 1 0 9 13 15 14 9 0 2
19 1 9 0 2 13 0 9 1 9 0 9 2 0 9 13 12 0 9 2
18 13 1 9 0 9 2 1 9 0 9 13 1 9 0 12 0 9 2
6 9 13 1 9 3 2
14 13 1 9 9 9 2 9 13 1 9 13 9 9 2
10 9 13 13 2 16 13 0 9 9 2
8 0 9 13 9 1 9 9 2
12 9 13 2 16 0 9 13 9 1 9 9 2
10 0 13 9 2 9 9 13 1 9 2
10 3 9 9 9 13 15 1 9 9 2
5 9 13 9 9 2
6 9 13 1 13 9 2
7 9 13 15 1 0 9 2
13 1 9 0 13 1 9 0 9 7 9 12 9 2
15 9 15 9 4 3 13 7 9 13 1 0 9 0 9 2
8 7 13 14 9 1 0 9 2
15 13 0 2 0 9 1 0 9 7 3 13 2 0 9 2
5 9 9 15 13 2
4 13 1 9 2
8 9 13 1 9 2 13 9 2
10 1 9 13 15 9 1 9 1 9 2
7 7 15 14 13 7 13 2
7 7 13 3 14 1 9 2
6 13 14 1 9 9 2
10 13 0 9 1 0 9 7 13 9 2
8 0 0 9 13 15 14 9 2
14 9 14 1 9 1 0 9 13 7 14 13 9 9 2
12 13 15 1 9 2 3 7 13 1 0 9 2
4 13 9 0 2
5 1 9 3 13 2
12 1 9 13 15 1 9 9 0 9 9 9 2
6 1 9 13 15 9 2
5 13 3 0 9 2
17 9 13 1 9 9 2 0 13 15 15 1 0 9 9 0 9 2
7 9 1 9 13 1 15 2
7 13 1 15 9 1 9 2
4 9 13 4 2
11 0 9 2 13 4 14 13 15 0 9 2
13 13 4 1 9 2 0 3 13 9 0 0 9 2
4 14 13 4 2
7 2 7 3 13 9 0 2
8 2 7 0 0 9 13 0 2
7 1 9 9 13 12 9 2
6 13 0 0 9 9 2
5 2 3 15 13 2
9 14 9 9 14 13 13 1 9 2
5 13 0 3 9 2
7 9 9 13 15 1 9 2
6 9 3 13 0 9 2
10 2 7 13 9 1 15 1 9 9 2
10 13 1 9 7 14 13 2 9 13 2
9 2 13 1 9 2 13 9 13 2
15 13 9 1 9 7 9 13 2 16 13 15 1 9 9 2
5 13 15 7 13 2
9 2 9 13 2 16 13 1 15 2
11 2 15 14 13 9 2 16 15 3 13 2
7 14 3 13 3 1 9 2
18 9 13 15 7 13 13 0 9 2 7 9 13 1 3 13 3 9 2
8 2 7 3 13 14 0 9 2
9 2 9 13 13 9 0 0 9 2
6 9 13 15 3 0 2
6 2 7 3 13 9 2
7 2 13 2 0 13 9 2
6 2 14 3 15 13 2
7 2 9 13 15 1 9 2
6 9 14 13 0 9 2
6 7 9 13 1 9 2
7 7 9 3 13 7 13 2
6 7 9 13 0 9 2
5 15 9 14 13 2
8 2 3 2 14 13 0 2 2
7 2 14 9 0 13 2 2
7 13 15 2 13 1 9 2
5 13 2 9 9 2
9 13 1 13 9 9 9 9 9 2
10 2 13 2 9 9 2 0 9 13 2
13 13 1 9 14 9 9 2 16 4 9 3 13 2
7 1 0 9 13 4 3 2
4 13 1 9 2
6 9 13 1 15 13 2
12 1 9 1 0 9 13 1 9 9 1 9 2
8 14 9 14 13 14 15 13 2
4 14 13 9 2
3 13 9 2
6 2 13 2 9 9 2
13 14 14 4 2 9 9 2 13 1 0 9 9 2
6 13 9 2 16 13 2
28 3 13 1 13 9 1 9 2 7 9 9 9 13 1 13 1 0 9 9 2 16 9 15 13 1 0 9 2
3 13 9 2
10 13 1 0 9 1 9 9 7 9 2
5 2 13 9 9 2
9 9 7 15 9 14 13 1 9 2
6 14 9 13 0 9 2
7 9 15 1 0 9 13 2
4 2 13 15 2
13 9 2 13 1 0 9 2 13 2 16 15 13 2
20 16 13 1 9 9 7 9 9 1 9 13 1 9 9 0 2 9 13 13 2
7 2 9 2 9 15 13 2
8 13 2 7 9 9 4 13 2
5 14 13 13 9 2
2 13 2
3 13 15 2
4 13 14 13 2
14 0 9 9 9 13 1 0 2 14 3 13 1 9 2
3 9 13 2
6 1 9 13 0 9 2
21 3 2 16 9 13 1 9 12 9 1 9 2 3 9 13 9 1 9 13 9 2
17 13 15 9 1 0 9 0 2 0 9 14 13 15 1 0 9 2
9 1 12 9 9 13 13 9 9 2
6 9 13 15 14 12 2
11 13 15 9 9 0 1 9 0 2 0 2
4 13 15 9 2
5 13 4 0 9 2
5 13 9 1 9 2
8 2 13 2 14 13 9 2 2
6 3 9 13 0 0 2
11 2 3 2 9 2 14 1 15 13 2 2
5 13 9 2 2 2
12 1 0 9 13 15 0 0 9 13 15 9 2
9 13 13 0 9 13 1 0 9 2
12 13 1 0 0 9 0 1 15 9 1 9 2
11 13 2 16 9 13 15 2 16 13 9 2
22 16 14 13 0 1 13 9 9 2 14 13 9 9 7 13 15 3 3 1 0 9 2
12 13 0 1 15 2 16 9 0 15 14 13 2
6 14 4 13 9 0 2
15 3 13 14 9 2 7 0 0 9 3 13 0 0 9 2
11 9 7 0 9 13 13 1 15 0 9 2
11 13 4 1 9 9 2 0 13 1 9 2
10 13 1 15 3 2 3 9 15 13 2
9 14 3 13 3 0 1 0 9 2
18 9 13 9 2 3 13 15 9 2 16 9 13 3 13 1 0 9 2
14 9 9 2 9 9 2 13 1 15 1 3 13 9 2
6 3 13 15 1 9 2
10 1 9 13 15 7 13 15 1 9 2
5 3 13 15 9 2
9 13 15 1 9 7 13 1 9 2
3 13 9 2
7 13 9 0 9 0 9 2
10 1 0 9 13 9 1 9 0 9 2
18 12 9 13 1 9 2 16 9 13 15 9 1 0 2 0 9 9 2
4 9 13 3 2
6 2 1 9 15 13 2
7 2 7 13 14 1 9 2
10 13 9 13 1 0 13 9 9 0 2
14 9 14 13 3 2 0 9 4 3 13 1 9 9 2
14 2 3 2 3 2 13 2 13 2 16 4 14 3 2
6 2 9 15 3 13 2
3 2 13 2
4 13 2 9 2
9 1 13 9 9 13 15 13 9 2
4 9 9 13 2
4 9 13 15 2
10 2 9 14 13 1 15 1 9 9 2
2 13 2
2 13 2
24 0 2 0 9 13 0 9 0 9 2 3 13 0 9 2 13 1 0 9 0 1 13 9 2
3 3 13 2
6 9 14 13 1 9 2
6 9 13 15 13 3 2
5 9 13 0 9 2
6 13 15 1 0 9 2
6 3 13 12 0 9 2
5 9 13 15 3 2
9 13 9 0 9 2 16 13 9 2
8 13 1 9 13 0 0 9 2
13 13 13 2 3 2 14 13 14 2 13 15 9 2
9 2 9 13 9 2 9 1 9 2
2 13 2
8 13 15 9 7 13 1 9 2
3 2 13 2
7 13 15 1 9 9 0 2
3 7 13 2
12 2 9 2 15 15 13 2 16 14 13 9 2
3 13 9 2
6 3 13 1 9 9 2
6 13 2 16 13 9 2
15 1 0 9 13 1 8 2 0 1 9 2 14 14 13 2
14 14 9 15 13 0 9 2 3 13 13 0 9 9 2
5 14 13 0 9 2
7 13 15 14 9 1 9 2
18 7 16 13 1 9 7 13 1 12 9 2 9 14 13 1 0 9 2
5 14 9 13 0 2
6 9 9 15 14 13 2
20 2 1 0 9 13 4 1 9 2 16 13 1 15 12 9 13 1 9 2 2
10 3 2 9 9 9 9 0 13 9 2
4 3 13 9 2
12 9 1 9 4 13 1 9 0 9 2 9 2
8 13 14 9 1 9 1 9 2
35 13 15 14 0 9 9 9 2 9 0 9 13 1 0 8 2 2 0 9 9 9 2 9 9 1 13 1 15 9 3 9 7 13 9 2
14 9 13 15 1 9 9 2 0 13 4 9 0 9 2
7 1 3 9 9 13 9 2
7 13 14 12 9 1 9 2
11 3 0 9 13 13 1 13 9 1 9 2
10 9 1 0 9 13 0 9 0 9 2
4 3 15 13 2
8 9 0 13 0 9 9 9 2
14 14 15 14 13 15 13 2 0 13 9 1 9 9 2
8 13 14 14 9 1 0 9 2
8 9 0 9 13 3 0 9 2
14 1 9 9 3 13 9 9 2 13 9 7 13 9 2
12 13 1 9 7 9 9 9 13 15 1 9 2
9 2 7 13 1 9 0 13 9 2
7 14 13 9 9 1 9 2
9 2 14 14 0 9 15 13 4 2
18 9 13 3 3 0 2 13 0 9 2 7 13 3 13 9 14 3 2
7 14 13 2 1 9 13 2
8 2 13 15 1 15 2 9 2
4 2 13 15 2
10 9 13 2 16 14 13 9 0 9 2
6 13 0 0 0 9 2
17 9 9 13 13 1 9 1 9 0 9 2 0 13 1 9 9 2
17 9 13 15 9 13 2 13 9 1 9 2 0 13 9 1 9 2
13 3 0 13 14 9 0 9 1 9 0 0 9 2
5 3 3 9 13 2
7 3 4 13 13 1 9 2
15 14 0 9 9 13 2 16 9 13 4 13 0 9 9 2
8 13 4 1 9 13 0 9 2
7 13 4 3 9 0 9 2
10 2 1 9 14 3 14 13 9 2 2
12 13 2 13 13 9 2 13 7 13 1 0 2
10 2 13 2 13 9 1 9 2 2 2
5 13 9 0 9 2
6 13 9 0 2 0 2
7 1 9 9 13 14 3 2
4 7 13 15 2
6 1 9 3 13 4 2
6 13 4 7 13 4 2
10 0 9 15 13 2 15 13 3 3 2
16 13 4 1 15 2 16 1 9 9 13 1 9 1 9 9 2
4 9 13 9 2
17 3 14 1 9 13 4 1 12 2 16 13 4 13 1 0 9 2
6 12 9 13 0 9 2
11 9 0 9 2 9 0 13 12 8 9 2
25 9 2 0 13 0 1 9 9 9 9 0 1 9 0 2 13 1 0 9 14 0 9 9 0 2
8 0 9 13 9 9 1 12 2
2 13 2
2 13 2
5 13 15 15 9 2
8 1 9 13 1 14 12 9 2
6 9 13 1 9 3 2
10 13 1 9 7 13 1 9 9 0 2
14 9 9 13 9 1 9 13 1 0 9 0 9 9 2
8 9 13 14 0 9 7 9 2
15 9 9 13 0 2 7 9 0 13 15 1 13 0 9 2
7 0 9 13 4 1 9 2
6 9 13 9 0 9 2
20 9 0 9 1 9 0 13 9 1 9 9 1 9 9 7 13 9 0 9 2
5 9 13 1 9 2
9 9 13 9 9 1 9 7 9 2
10 9 13 2 16 13 13 1 9 9 2
10 14 2 12 1 0 9 13 15 9 2
6 1 9 13 9 9 2
13 1 9 13 15 12 0 9 2 0 13 1 9 2
5 12 9 3 13 2
7 9 9 13 1 9 9 2
10 1 9 9 13 9 1 9 0 9 2
9 3 9 13 14 12 8 2 8 2
8 1 9 1 9 13 0 9 2
10 12 9 9 13 1 13 12 8 8 2
9 13 9 9 7 9 0 9 0 2
2 13 2
12 1 8 2 9 9 13 1 9 0 0 9 2
8 1 9 0 13 0 9 9 2
18 13 2 16 3 13 1 0 2 0 9 2 13 9 2 1 9 0 2
16 9 4 13 1 9 7 13 13 9 9 9 0 9 7 9 2
7 12 13 1 9 1 9 2
12 13 14 13 9 2 0 13 1 9 9 9 2
17 3 13 14 1 9 0 9 1 9 13 9 7 13 1 15 9 2
15 13 14 12 0 9 0 2 9 13 0 1 0 9 9 2
18 7 3 14 13 9 2 0 3 3 13 15 9 2 0 9 3 13 2
4 13 9 3 2
5 7 13 14 13 2
15 9 2 1 9 13 1 9 1 9 2 1 9 13 9 2
15 9 9 13 2 16 9 9 9 14 13 1 9 1 9 2
12 0 9 13 15 2 16 3 13 13 9 9 2
10 9 13 3 0 2 0 7 0 9 2
5 13 2 16 13 2
12 9 15 13 2 16 13 15 13 7 13 9 2
14 13 15 3 7 13 1 15 9 3 0 1 15 0 2
16 16 1 0 13 9 9 7 13 1 0 9 9 2 13 3 2
11 1 0 9 3 3 13 4 15 3 0 2
10 14 9 1 9 0 13 1 15 9 2
24 3 2 1 12 9 13 2 13 1 9 13 1 9 2 9 15 1 15 13 1 0 0 9 2
31 9 9 13 3 2 16 1 0 0 9 13 9 0 9 7 1 0 13 1 13 9 2 1 0 13 13 15 14 1 9 2
6 9 13 2 16 13 2
12 0 9 13 14 0 9 9 2 9 7 9 2
7 0 9 13 15 15 13 2
10 1 0 9 13 15 9 14 12 9 2
4 13 15 9 2
4 13 13 9 2
5 13 0 13 9 2
20 3 1 8 2 0 1 9 8 2 0 12 9 13 15 1 13 1 9 9 2
4 13 1 9 2
10 0 9 14 14 13 13 0 9 9 2
6 13 1 9 0 9 2
10 1 9 0 1 9 9 13 15 9 2
8 13 2 16 13 9 1 9 2
10 3 13 15 9 1 12 9 9 9 2
7 9 13 15 1 0 9 2
10 1 9 9 14 13 2 1 0 9 2
15 14 1 0 0 9 13 4 9 9 1 0 9 1 9 2
2 13 2
5 9 1 15 13 2
5 14 9 14 13 2
11 9 13 3 3 2 7 9 13 1 9 2
9 13 2 7 14 13 1 9 9 2
10 14 13 14 2 9 15 13 1 9 2
8 14 13 2 3 15 3 13 2
5 13 15 1 9 2
6 7 9 13 1 9 2
6 9 13 9 1 9 2
9 13 0 9 13 9 1 0 9 2
11 9 13 1 9 2 15 9 14 13 9 2
22 9 13 14 15 1 12 0 9 2 7 14 9 1 9 2 13 15 9 7 9 9 2
18 1 9 13 9 0 13 1 9 0 9 9 2 9 7 0 13 9 2
6 3 14 13 1 9 2
7 1 12 9 13 1 9 2
10 7 14 13 15 13 1 13 9 9 2
5 13 1 9 9 2
16 1 0 9 1 9 9 13 2 16 0 0 9 3 15 13 2
11 9 0 13 9 9 9 1 0 9 9 2
18 13 0 9 2 16 9 0 4 15 1 15 13 9 1 9 9 0 2
21 9 9 0 13 2 16 9 13 0 9 1 9 9 2 0 13 0 9 1 9 2
8 9 4 13 1 9 1 9 2
17 9 13 1 15 9 1 0 9 9 2 0 13 1 0 9 9 2
5 3 13 9 9 2
8 9 9 9 13 14 9 9 2
10 3 13 15 1 9 9 0 1 9 2
9 9 1 9 14 13 1 9 9 2
7 0 9 13 3 0 9 2
9 13 1 15 9 2 14 13 9 2
8 14 13 2 16 9 13 0 2
9 13 2 16 3 15 1 15 13 2
12 9 3 13 15 1 9 2 13 15 1 9 2
6 13 1 15 12 9 2
7 3 15 13 1 0 9 2
11 0 9 13 14 13 0 0 9 1 9 2
8 9 13 16 4 13 1 9 2
16 0 9 13 13 0 13 9 1 0 9 2 0 13 0 9 2
17 7 1 9 13 4 2 16 13 4 2 16 13 3 0 7 0 2
7 13 4 1 9 12 9 2
5 3 15 13 4 2
10 16 14 13 9 2 14 13 9 0 2
12 3 3 1 9 1 9 13 15 3 0 9 2
19 14 13 14 9 1 9 13 1 9 2 0 14 13 1 0 9 0 9 2
9 13 3 0 7 13 1 15 9 2
5 1 0 13 9 2
10 2 0 13 0 9 9 1 0 9 2
7 2 0 13 9 9 9 2
6 0 9 13 13 9 2
3 13 9 2
9 13 0 0 9 2 9 2 2 2
14 1 15 9 13 9 9 2 13 15 1 9 2 2 2
10 7 3 13 15 9 1 0 9 13 2
7 3 13 4 13 0 9 2
10 1 9 0 9 13 15 9 2 2 2
11 14 2 13 9 13 2 16 1 15 13 2
4 13 15 9 2
8 2 3 14 13 14 3 3 2
6 2 14 13 2 9 2
11 2 7 3 14 13 14 4 15 13 3 2
8 13 14 4 15 14 1 9 2
8 15 13 1 0 9 1 9 2
7 2 13 2 9 15 13 2
6 3 14 13 0 9 2
7 15 9 13 15 14 9 2
6 9 13 1 0 9 2
3 9 13 2
5 13 1 0 9 2
8 9 13 15 1 0 0 9 2
8 9 13 15 7 13 1 15 2
16 1 0 9 14 13 0 9 7 9 2 14 0 2 0 9 2
9 1 9 13 2 9 1 9 13 2
5 13 1 15 9 2
5 13 15 0 9 2
14 2 13 13 1 0 9 2 9 2 3 15 14 13 2
5 13 13 9 9 2
2 13 2
3 13 15 2
6 13 4 13 15 9 2
7 13 4 15 9 1 9 2
5 13 4 1 15 2
12 7 13 4 15 13 2 16 14 13 0 9 2
9 0 9 1 0 9 13 3 3 2
18 0 9 13 0 0 9 1 0 0 9 2 1 0 13 15 0 9 2
16 0 9 2 0 1 0 0 9 1 9 2 13 0 13 9 2
8 13 9 2 9 13 0 9 2
11 1 9 13 4 1 0 9 0 9 9 2
21 14 1 0 9 1 9 9 0 2 9 0 13 0 0 9 0 2 0 15 13 2
8 14 13 2 14 13 13 9 2
13 3 15 13 9 1 9 9 7 0 9 1 9 2
6 3 15 3 3 13 2
