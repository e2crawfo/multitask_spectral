131 11
8 9 13 0 7 13 0 9 2
10 11 3 4 3 13 0 0 9 9 2
20 12 9 9 13 11 11 9 0 9 11 9 9 1 7 13 15 3 3 13 2
16 12 9 13 9 9 7 9 1 2 16 11 4 4 15 13 2
17 15 9 16 11 9 9 9 13 2 13 0 11 3 15 11 9 2
18 9 13 11 0 2 9 13 15 3 3 9 11 11 16 0 11 11 2
18 9 13 11 9 3 0 9 9 2 16 13 9 9 7 9 9 1 2
13 9 4 13 2 15 9 13 11 9 7 9 9 2
19 15 9 13 13 11 9 9 9 9 7 15 9 1 9 11 9 13 4 2
3 9 9 1
14 2 9 1 9 4 13 2 2 13 11 9 0 9 2
8 15 4 13 3 9 11 9 2
4 9 13 9 2
3 9 9 9
10 13 0 0 9 2 9 13 3 12 2
11 15 9 13 9 9 3 9 15 0 9 2
34 3 9 13 0 9 9 7 9 2 7 16 9 13 7 9 13 0 2 13 15 3 0 7 0 3 13 9 2 15 4 3 3 13 2
8 3 13 9 3 15 0 9 2
7 0 9 13 9 1 9 2
10 11 7 11 13 0 9 1 0 9 2
4 11 13 3 2
6 7 3 13 11 3 2
4 11 13 9 2
7 9 13 15 0 9 9 2
14 9 13 1 9 0 9 1 0 9 9 1 3 3 2
8 7 11 7 11 13 0 9 2
7 9 13 9 9 3 9 2
10 9 0 9 7 0 9 13 9 9 2
7 9 12 13 15 15 9 2
11 11 13 12 0 9 12 9 9 1 9 2
10 9 13 3 0 9 0 9 7 9 2
8 16 9 1 13 9 0 9 2
8 9 13 3 9 1 9 13 2
5 13 9 1 9 2
5 13 9 7 9 2
5 9 13 9 3 2
6 15 4 9 3 13 2
6 15 13 3 3 9 2
5 9 13 15 9 2
6 9 13 15 9 9 2
6 9 13 9 9 1 2
8 15 9 13 15 0 9 9 2
6 15 13 0 9 3 2
7 15 13 0 9 1 9 2
6 15 13 3 9 3 2
6 9 13 3 16 9 2
8 0 9 9 13 15 9 1 2
5 9 13 9 1 2
4 9 13 9 2
12 1 0 9 13 15 0 9 1 9 0 9 2
7 3 13 9 9 11 1 2
7 3 13 15 9 3 3 2
4 13 9 1 2
5 13 9 1 3 2
11 15 9 13 9 11 1 9 15 9 1 2
4 13 15 0 2
10 15 0 11 13 3 15 9 9 13 2
7 11 13 15 9 1 9 2
9 3 13 15 9 9 3 9 13 2
4 13 9 9 2
5 13 9 9 1 2
6 3 13 15 12 9 2
11 9 7 9 1 0 0 9 13 9 9 2
5 13 9 1 9 2
4 9 13 15 2
6 15 13 9 15 9 2
7 9 3 13 15 15 1 2
7 15 13 15 9 9 1 2
6 15 13 9 1 3 2
6 13 15 9 9 9 2
6 15 13 15 9 3 2
8 15 13 9 1 9 0 9 2
8 15 1 13 0 9 0 11 2
7 0 11 13 15 1 9 2
8 11 13 11 9 1 9 13 2
4 13 3 9 2
13 3 15 9 16 3 13 11 3 3 0 9 9 2
6 13 9 15 9 3 2
5 13 3 1 9 2
6 9 13 9 9 9 2
4 9 13 9 2
4 13 9 1 2
4 9 13 13 2
5 13 9 9 13 2
10 0 9 13 1 0 0 9 0 11 2
4 9 13 9 2
7 9 13 0 9 9 3 2
5 9 13 9 3 2
4 13 9 9 2
4 13 1 9 2
7 9 13 9 9 9 13 2
6 11 13 9 1 9 2
9 11 13 9 9 9 9 9 1 2
9 9 13 9 1 9 7 9 1 2
9 9 13 9 1 9 9 9 13 2
5 1 9 13 9 2
5 11 13 9 1 2
5 9 13 9 9 2
6 9 13 9 11 1 2
4 11 13 9 2
6 11 13 9 9 9 2
4 11 13 9 2
6 11 13 9 9 9 2
9 11 13 15 1 1 9 12 9 2
6 9 13 9 9 1 2
5 9 13 9 3 2
5 9 13 9 13 2
6 9 13 9 9 13 2
5 9 13 11 11 2
5 9 13 9 9 2
8 11 13 1 9 13 9 13 2
5 9 13 11 9 2
7 11 13 9 9 1 9 2
4 11 13 0 2
5 11 13 9 1 2
8 9 13 9 1 0 9 1 2
6 11 13 9 9 1 2
4 9 13 9 2
5 11 13 9 9 2
4 9 13 9 2
9 11 13 9 9 1 9 9 13 2
4 9 13 9 2
6 11 13 9 9 9 2
5 9 13 15 1 2
7 11 13 9 9 9 13 2
8 9 13 9 9 9 9 13 2
7 11 13 9 11 9 13 2
5 11 13 9 9 2
4 11 9 13 2
8 15 15 11 14 11 13 15 14
1 2
