6800 17
14 1 9 9 9 9 13 9 1 9 0 9 9 9 2
9 1 9 9 9 9 13 1 9 2
13 7 9 9 9 13 9 9 9 1 9 2 2 2
7 3 9 0 7 13 0 2
11 13 15 1 9 12 9 1 9 9 9 2
13 1 0 9 9 9 9 9 13 9 1 0 9 2
15 1 9 3 1 9 7 9 1 0 9 9 13 0 9 2
29 3 13 0 9 2 13 1 15 9 2 13 1 15 0 9 1 9 2 0 3 0 9 13 1 9 1 9 9 2
18 1 9 13 0 9 13 0 9 7 3 3 13 15 1 9 1 9 2
5 2 9 9 13 2
8 9 13 9 7 13 1 9 2
7 9 13 3 1 15 9 2
19 1 9 9 13 1 0 9 14 13 14 2 16 0 9 13 1 0 13 2
5 3 13 13 9 2
4 14 13 9 2
8 13 9 13 13 1 9 0 2
11 13 15 0 0 9 0 9 0 1 9 2
20 0 9 9 13 14 9 0 9 2 1 0 0 9 9 13 1 13 9 9 2
7 9 13 9 7 13 9 2
11 13 4 0 9 7 13 4 15 3 13 2
9 13 14 4 3 13 1 9 9 2
10 13 4 15 1 9 7 13 4 9 2
14 9 13 15 1 9 2 9 9 13 1 9 1 9 2
16 1 9 13 4 12 9 1 9 2 7 9 13 4 0 9 2
3 13 15 2
25 1 9 3 13 1 9 9 9 9 9 0 1 9 9 9 7 8 2 9 2 3 13 9 9 2
5 3 3 13 9 2
13 9 2 9 13 9 2 3 1 9 13 15 9 2
16 9 9 13 9 9 9 1 9 0 1 0 2 13 9 9 2
8 0 1 15 14 13 14 9 2
15 13 15 14 9 9 2 0 13 9 2 16 13 9 0 2
9 9 13 14 9 1 9 7 9 2
4 9 4 0 2
15 16 14 13 2 7 14 4 1 3 13 2 16 4 13 2
5 7 13 0 9 2
8 1 0 9 13 15 1 9 2
18 2 13 9 1 9 9 13 0 2 7 1 9 9 9 13 13 9 2
17 2 14 9 0 13 9 13 1 0 9 2 7 13 1 13 9 2
13 14 1 15 14 13 2 16 9 0 13 3 3 2
4 9 3 13 2
9 2 14 13 2 16 4 15 13 2
19 13 1 15 9 9 9 1 9 2 9 2 9 2 9 2 9 7 9 2
17 9 13 9 4 13 1 9 9 1 9 0 9 9 0 1 9 2
28 9 0 9 9 9 13 14 9 9 0 1 0 9 2 1 0 15 9 4 9 0 9 0 2 0 9 9 2
14 9 13 15 3 1 8 2 0 1 9 0 9 0 2
9 13 14 2 16 13 1 0 9 2
16 2 9 13 9 0 2 9 13 2 1 0 0 9 13 9 2
15 0 1 0 9 4 13 1 9 3 1 0 9 1 9 2
7 9 9 4 0 9 9 2
6 9 13 12 0 9 2
22 9 13 9 9 0 7 9 2 13 1 9 0 2 13 9 9 9 7 13 1 9 2
19 13 14 1 15 9 0 1 9 13 1 9 2 13 2 13 2 13 9 2
19 13 9 1 9 9 0 1 9 2 9 0 2 0 9 2 9 7 9 2
15 1 9 0 9 3 13 15 0 2 0 2 0 7 0 2
20 1 15 13 15 1 9 13 9 2 13 15 13 9 0 2 3 13 0 9 2
6 0 9 13 15 9 2
5 9 9 13 0 2
7 13 1 9 1 0 9 2
6 2 0 9 13 3 2
5 2 13 3 3 2
6 13 4 15 14 9 2
8 2 14 13 2 9 15 13 2
5 3 13 4 9 2
11 15 9 13 0 2 0 2 13 1 9 2
9 3 13 4 2 16 13 1 15 2
4 13 4 9 2
15 2 14 14 13 13 2 16 14 9 0 13 15 1 9 2
16 1 9 0 0 9 7 9 2 7 14 9 13 1 0 9 2
12 9 9 9 0 1 13 9 0 3 13 9 2
5 13 15 14 3 2
7 9 0 9 13 9 0 2
16 2 1 0 9 14 13 9 2 0 13 9 3 13 1 9 2
5 9 15 14 13 2
6 9 15 14 3 13 2
7 16 3 13 4 13 9 2
8 4 4 13 1 14 0 9 2
9 16 14 13 4 13 1 9 9 2
18 1 0 9 9 13 9 1 9 2 13 1 15 9 7 13 1 9 2
8 7 0 9 13 15 1 15 2
6 14 13 15 15 9 2
11 1 9 0 0 9 14 13 9 7 9 2
11 3 0 0 9 1 0 9 9 13 9 2
19 7 16 9 13 15 13 1 9 2 0 13 9 13 4 15 13 1 15 2
12 16 3 13 2 13 15 9 1 12 9 9 2
8 1 9 14 13 15 15 9 2
13 0 0 0 9 3 14 13 9 1 9 9 0 2
9 13 3 9 9 9 1 9 0 2
6 9 13 1 9 9 2
19 9 14 4 14 13 13 0 9 2 16 13 15 9 7 13 15 1 9 2
16 1 9 0 0 9 1 0 9 13 9 0 9 0 1 9 2
14 2 1 9 13 12 9 2 3 13 4 0 9 13 2
12 9 13 15 14 1 9 1 9 9 9 9 2
4 13 15 9 2
5 9 9 14 13 2
6 9 1 9 15 13 2
7 3 9 13 1 9 0 2
7 1 15 13 13 0 9 2
17 9 2 0 13 15 13 1 9 0 9 2 13 13 1 9 0 2
10 9 13 9 1 0 9 1 13 9 2
9 9 9 13 9 9 1 9 0 2
6 2 13 14 3 0 2
7 13 3 0 1 0 9 2
5 3 15 14 13 2
5 13 1 9 9 2
7 13 9 14 13 1 9 2
5 9 13 0 9 2
14 14 9 2 13 15 2 13 13 14 3 0 9 2 2
6 7 3 4 13 9 2
10 1 9 2 9 9 7 9 13 9 2
16 13 14 9 1 9 2 7 14 13 9 1 9 14 1 9 2
8 4 13 2 13 9 7 9 2
6 1 9 9 13 9 2
6 13 3 1 9 9 2
12 1 9 9 9 1 12 9 13 15 0 9 2
12 9 0 9 7 15 9 13 15 14 9 9 2
9 13 0 9 13 15 1 9 9 2
13 3 9 1 9 13 9 7 13 15 1 13 9 2
7 13 14 12 8 2 8 2
12 0 9 13 1 9 2 1 12 9 13 9 2
10 3 13 1 9 9 2 1 9 13 2
8 0 9 13 9 9 9 9 2
7 13 0 9 13 12 9 2
5 1 9 13 9 2
9 1 0 9 13 9 13 1 9 2
13 3 13 1 9 7 1 9 13 9 9 0 9 2
7 13 9 2 3 1 9 2
6 3 9 15 14 13 2
7 1 0 9 13 0 9 2
14 1 9 13 14 13 2 16 13 9 1 9 1 9 2
5 1 9 13 9 2
7 0 9 13 13 1 9 2
6 3 13 9 1 9 2
10 16 9 14 13 1 9 2 13 9 2
6 1 9 9 15 13 2
6 9 13 15 1 9 2
8 13 13 9 1 0 9 9 2
21 13 1 15 13 1 9 2 13 0 9 2 9 9 2 1 9 13 15 1 9 2
12 1 0 9 13 9 2 1 12 1 12 9 2
15 9 13 9 13 9 2 0 3 13 1 0 9 9 9 2
5 13 13 14 0 2
15 1 0 13 9 7 13 15 1 9 2 16 13 9 9 2
14 3 13 9 0 9 2 16 9 13 1 15 3 13 2
8 13 1 0 9 0 9 0 2
7 0 9 0 9 13 9 2
4 0 9 13 2
22 9 9 13 13 0 2 16 1 9 13 14 9 2 0 14 13 15 1 9 0 9 2
20 1 9 13 14 9 14 12 0 9 2 0 13 15 1 9 1 9 9 9 2
13 13 15 2 16 9 13 15 13 1 15 0 9 2
7 9 13 9 13 1 9 2
13 9 9 2 9 9 2 14 13 9 1 12 9 2
15 3 4 3 2 16 14 0 9 13 2 14 13 9 9 2
5 1 9 9 13 2
7 9 13 15 3 9 0 2
17 1 9 9 1 9 13 12 9 2 0 1 9 13 1 0 9 2
9 1 9 13 14 3 13 0 9 2
11 9 13 9 9 1 9 1 9 1 9 2
11 16 9 13 14 9 2 13 13 9 9 2
4 13 15 9 2
9 3 14 13 9 2 14 13 9 2
9 16 9 4 13 9 1 0 9 2
6 0 13 9 13 9 2
8 2 3 13 15 1 9 9 2
10 9 13 9 2 13 9 2 13 9 2
3 13 9 2
6 9 13 15 1 9 2
5 13 2 4 13 2
13 2 3 9 13 2 13 15 1 9 1 0 9 2
11 2 14 13 9 0 2 13 14 3 13 2
7 9 9 1 9 14 13 2
12 2 9 13 15 2 16 14 13 13 9 9 2
23 9 9 7 9 13 1 9 0 2 9 1 9 9 4 13 9 1 9 1 9 15 9 2
17 9 9 3 13 1 9 0 2 7 1 0 13 9 14 13 15 2
5 9 14 14 13 2
6 1 9 13 0 9 2
5 13 9 1 9 2
11 14 13 15 3 2 16 14 13 0 9 2
6 2 9 14 13 9 2
5 13 13 0 9 2
8 13 9 2 9 0 2 12 2
13 0 9 13 15 1 13 9 7 13 9 1 9 2
5 13 1 9 9 2
21 1 0 9 9 13 4 9 9 9 2 9 2 0 9 9 2 3 13 0 9 2
9 14 13 13 1 9 1 0 9 2
6 7 3 13 9 9 2
11 9 13 9 7 1 9 14 13 15 13 2
9 0 0 9 13 0 0 9 9 2
4 3 13 0 2
8 1 9 14 13 15 15 13 2
7 14 13 15 3 1 9 2
6 9 15 3 14 13 2
10 2 1 9 13 15 1 0 9 2 2
8 3 13 2 16 0 9 13 2
7 12 0 9 13 1 9 2
13 1 9 9 2 9 13 9 9 13 14 1 9 2
12 1 9 9 0 7 9 13 15 3 12 9 2
19 0 9 0 13 15 2 1 9 9 9 2 9 9 1 0 9 9 0 2
9 9 8 2 13 9 1 0 9 2
12 15 9 3 14 13 2 7 14 13 0 9 2
16 9 9 2 9 0 2 13 15 2 16 9 0 14 4 13 2
15 16 14 9 0 15 13 2 9 13 15 14 1 0 9 2
11 0 9 13 2 16 14 13 9 9 13 2
8 1 0 9 9 14 13 9 2
12 9 13 1 0 9 13 1 9 1 0 9 2
9 13 15 2 16 9 13 15 13 2
16 1 9 1 9 9 3 1 9 13 13 1 13 9 1 9 2
3 13 9 2
9 3 9 13 2 16 13 1 9 2
12 3 9 13 1 9 13 1 9 0 1 9 2
22 1 0 9 9 3 13 1 9 2 9 15 13 2 7 9 13 7 13 9 1 9 2
6 9 13 9 7 9 2
5 9 13 13 9 2
16 3 9 4 13 13 9 9 2 0 3 13 1 0 9 9 2
7 1 13 9 13 12 9 2
7 12 0 9 13 15 9 2
4 12 9 13 2
6 12 9 13 15 9 2
13 9 7 9 13 1 9 9 14 13 13 1 9 2
5 9 13 0 9 2
10 3 1 0 2 12 0 9 13 3 2
6 3 13 9 0 9 2
7 0 9 14 13 0 9 2
5 14 9 15 13 2
14 9 2 0 13 1 9 2 1 0 9 4 13 9 2
12 14 13 9 1 9 7 14 13 9 1 9 2
5 13 9 9 9 2
3 13 9 2
7 3 9 13 9 0 9 2
12 1 12 0 9 9 13 3 13 9 7 9 2
18 9 9 1 9 9 13 2 16 13 1 0 9 9 2 7 14 13 2
12 9 9 13 9 2 0 13 1 9 1 9 2
8 9 0 4 13 1 9 0 2
12 9 13 2 16 9 13 1 9 1 12 9 2
13 16 14 13 9 1 15 9 2 9 13 1 9 2
7 0 9 13 15 3 3 2
5 14 13 14 9 2
6 1 9 9 4 0 2
10 1 9 9 9 0 4 13 15 13 2
4 9 0 13 2
15 13 15 0 9 1 0 9 13 15 9 1 9 0 9 2
4 13 0 9 2
8 9 13 15 3 0 1 9 2
10 9 13 2 7 9 4 14 3 13 2
11 13 4 15 1 0 9 2 13 1 9 2
9 2 9 1 0 9 13 1 9 2
6 15 9 3 15 13 2
8 1 9 9 0 9 9 13 2
10 13 3 9 1 9 13 1 0 9 2
5 13 3 12 9 2
14 9 13 9 9 1 13 9 0 7 13 1 9 9 2
9 0 9 9 14 13 3 13 9 2
8 2 9 0 14 14 13 4 2
8 0 9 9 14 13 14 9 2
8 2 1 9 14 13 0 9 2
22 14 13 13 2 16 14 12 9 1 9 13 2 16 13 9 9 7 13 15 1 9 2
4 13 9 13 2
10 1 0 9 9 13 2 16 13 9 2
8 13 9 13 15 1 0 9 2
5 13 4 14 9 2
12 1 9 1 15 2 9 2 13 4 1 9 2
9 0 9 13 1 0 9 1 9 2
7 9 13 2 16 13 9 2
15 9 4 14 13 1 0 9 9 7 9 1 9 9 9 2
10 3 13 9 2 1 0 13 15 9 2
6 3 13 1 9 0 2
9 1 13 0 9 13 14 12 9 2
8 9 9 13 1 9 1 9 2
8 9 9 13 1 9 1 9 2
6 13 13 14 9 0 2
5 13 13 9 9 2
7 1 9 13 15 0 9 2
13 9 14 9 2 0 13 1 9 0 2 13 9 2
6 0 9 13 9 9 2
5 1 9 9 13 2
5 3 9 13 9 2
8 3 1 9 1 9 13 9 2
5 9 13 1 9 2
3 9 13 2
18 9 8 2 13 15 9 2 7 15 9 9 8 2 13 1 9 9 2
6 13 15 3 1 9 2
9 13 15 13 2 7 14 13 13 2
8 2 13 15 1 9 12 9 2
7 9 13 9 13 14 0 2
11 2 9 4 0 1 13 1 0 9 9 2
9 0 0 9 4 13 1 9 0 2
7 7 15 14 13 9 0 2
6 9 13 1 9 9 2
16 13 0 2 16 9 13 13 0 9 7 13 15 1 9 13 2
12 13 15 13 13 9 2 14 13 1 9 9 2
6 13 2 16 9 13 2
4 9 13 13 2
6 9 13 1 9 9 2
8 2 9 13 15 1 9 9 2
7 1 9 12 9 13 4 2
10 1 9 1 9 14 13 4 9 9 2
14 1 9 1 9 13 4 2 16 14 13 15 1 9 2
7 0 9 3 13 0 9 2
16 3 1 15 13 4 13 0 9 2 0 14 1 0 9 13 2
7 3 13 15 12 0 9 2
5 14 13 15 9 2
5 9 13 1 9 2
9 2 9 13 1 15 2 13 0 2
8 9 1 0 9 14 4 13 2
10 1 0 9 13 9 1 9 12 9 2
5 13 15 14 13 2
7 12 9 1 15 13 9 2
22 9 8 2 2 9 9 2 9 9 2 14 13 13 2 16 15 9 9 15 14 13 2
7 2 14 15 9 14 13 2
14 9 13 15 2 16 1 0 9 13 0 9 0 9 2
6 9 14 15 13 9 2
6 13 15 15 13 9 2
6 7 0 9 4 13 2
9 1 0 9 13 13 1 9 0 2
6 2 9 13 9 2 2
21 0 9 13 1 9 2 0 13 1 9 2 7 1 9 13 2 9 13 15 9 2
4 9 13 15 2
30 1 9 0 1 9 9 9 2 0 4 13 1 9 9 2 13 2 16 9 13 9 1 13 1 0 9 0 9 0 2
16 1 9 0 9 9 3 1 0 9 0 9 13 0 9 0 2
14 9 1 9 1 9 13 1 9 13 9 1 0 9 2
6 13 1 9 1 9 2
5 13 4 15 9 2
12 13 4 15 13 1 9 2 7 13 1 15 2
8 1 9 13 0 2 0 9 2
6 13 4 2 16 13 2
4 13 4 9 2
10 13 4 15 1 9 7 13 4 13 2
4 13 4 9 2
8 2 13 1 9 2 13 9 2
9 13 2 16 14 13 9 1 9 2
12 2 1 9 9 9 0 14 4 14 13 9 2
8 9 9 13 2 16 13 3 2
9 9 13 9 1 9 0 9 9 2
10 1 0 9 9 13 1 9 0 9 2
19 9 1 9 13 0 9 2 0 1 9 13 1 0 9 1 9 0 9 2
12 2 3 0 13 13 1 0 9 1 13 9 2
8 9 15 13 2 12 9 13 2
17 0 9 13 9 13 15 9 1 9 7 9 9 7 9 9 0 2
7 1 9 14 13 0 9 2
9 14 15 15 13 13 1 0 9 2
7 13 15 9 1 0 9 2
7 1 9 13 15 1 9 2
13 1 0 9 9 9 2 9 1 9 2 13 0 2
11 9 9 14 14 13 3 13 9 1 9 2
6 13 14 1 9 9 2
11 9 2 0 13 13 9 2 14 13 9 2
14 3 9 9 0 1 9 2 9 9 2 13 9 9 2
16 2 9 13 3 1 0 9 7 14 13 2 16 13 1 9 2
3 9 13 2
8 0 9 4 13 1 0 9 2
5 9 13 0 9 2
6 9 13 2 3 13 2
10 2 9 13 9 9 9 1 9 9 2
10 12 0 9 13 14 9 1 0 9 2
17 14 4 13 1 9 9 9 2 16 14 13 15 1 15 9 0 2
17 1 0 9 2 13 1 12 9 1 9 2 13 4 1 9 8 2
15 13 15 13 0 9 2 0 9 7 9 1 13 9 0 2
12 9 0 1 9 13 1 9 1 9 9 9 2
13 13 1 9 0 0 9 1 9 12 8 2 8 2
4 0 13 3 2
7 0 2 0 13 1 9 2
12 2 15 9 13 0 9 1 9 0 9 0 2
5 13 9 13 9 2
13 13 2 16 1 9 1 9 9 14 13 0 9 2
12 9 9 4 13 9 1 9 1 9 9 9 2
7 9 13 15 9 9 9 2
7 14 9 13 9 0 9 2
8 12 9 13 9 1 9 0 2
6 9 13 15 1 9 2
6 1 9 13 12 9 2
5 1 9 13 12 2
11 0 9 13 16 9 0 9 0 9 0 2
15 1 9 1 0 9 13 14 9 2 0 14 13 1 9 2
8 12 13 1 9 13 1 9 2
3 4 3 2
7 3 9 13 1 9 9 2
12 1 0 9 13 15 13 0 9 13 9 0 2
8 9 13 1 12 9 13 9 2
22 12 9 0 1 9 2 1 9 9 2 0 13 9 13 9 2 13 0 2 0 9 2
5 2 13 13 9 2
23 0 9 13 0 2 0 9 13 13 9 7 0 0 9 1 9 7 9 9 1 12 9 2
7 0 9 13 15 0 9 2
9 1 9 13 15 0 9 1 9 2
3 13 15 2
4 9 4 13 2
9 2 0 9 13 1 9 0 9 2
11 0 0 9 14 13 9 1 15 15 13 2
4 15 3 13 2
12 0 13 9 2 7 3 13 9 0 7 0 2
11 1 9 0 1 0 8 2 13 12 9 2
12 0 9 9 13 1 9 13 0 9 7 9 2
5 13 9 1 9 2
6 9 1 9 14 13 2
18 16 9 9 13 13 9 1 9 14 12 8 1 0 9 1 15 9 2
4 2 9 13 2
10 3 1 9 13 13 15 9 1 9 2
21 9 9 9 13 9 1 0 9 13 1 0 9 2 0 13 13 0 9 9 0 2
6 3 15 3 0 13 2
9 9 9 1 0 9 13 3 0 2
7 7 9 13 1 15 13 2
5 2 14 13 9 2
8 13 9 15 9 13 0 9 2
8 9 9 1 9 0 13 9 2
7 9 8 2 13 15 9 2
12 1 9 13 1 8 2 0 2 12 9 0 2
12 0 13 12 0 9 2 12 9 0 7 9 2
5 9 0 13 0 2
6 15 9 14 13 9 2
11 9 4 13 1 9 9 9 1 9 9 2
15 1 13 9 7 13 12 9 13 9 1 9 1 9 9 2
17 0 9 14 13 15 13 2 16 14 13 9 1 9 1 9 9 2
18 2 9 13 2 16 9 15 3 13 2 7 14 13 14 13 2 2 2
7 15 0 9 14 13 9 2
7 1 0 9 13 9 9 2
10 0 9 9 8 2 13 1 9 9 2
10 13 9 13 2 16 9 9 13 9 2
6 13 1 9 9 9 2
3 9 13 2
12 0 9 13 0 2 16 9 13 1 0 9 2
6 9 7 9 13 9 2
8 13 1 0 9 9 7 9 2
3 14 13 2
7 9 13 3 0 9 0 2
12 3 13 2 7 9 1 9 9 13 14 9 2
6 2 9 13 9 9 2
4 14 13 9 2
11 13 12 9 1 9 7 13 1 0 9 2
8 13 9 2 13 15 7 13 2
13 1 0 9 9 8 2 13 2 16 13 15 13 2
5 13 1 0 9 2
8 1 9 13 9 1 0 9 2
5 13 1 9 9 2
10 9 9 1 9 9 13 15 1 9 2
9 1 9 1 9 13 1 12 9 2
18 9 1 9 13 9 9 2 16 13 9 2 16 9 13 15 1 9 2
5 13 15 9 13 2
4 0 9 13 2
2 13 2
4 3 13 3 2
7 14 13 2 9 15 13 2
4 9 13 9 2
12 0 9 9 13 1 9 14 12 9 1 9 2
14 14 12 9 13 3 9 1 0 2 9 0 1 9 2
9 9 14 1 0 9 13 0 9 2
4 2 14 13 2
5 1 9 13 9 2
9 3 13 15 15 13 1 0 9 2
4 13 0 9 2
6 9 13 1 9 9 2
8 9 13 15 1 9 12 9 2
10 9 13 9 7 1 0 9 13 9 2
15 9 1 0 9 13 1 0 9 2 3 13 14 12 9 2
5 0 13 3 13 2
10 13 14 9 13 0 9 0 9 0 2
9 13 9 14 9 7 13 0 9 2
5 13 9 7 9 2
11 9 13 1 15 9 2 16 14 15 13 2
3 13 9 2
10 13 15 1 0 9 2 13 0 9 2
4 3 13 9 2
7 13 14 14 9 15 9 2
13 1 13 1 9 13 9 2 3 13 15 14 9 2
8 9 8 2 4 14 3 13 2
6 13 15 1 0 9 2
13 9 13 13 1 9 1 9 7 13 1 9 9 2
9 14 13 9 2 16 13 1 9 2
5 0 9 9 13 2
6 13 15 1 12 9 2
4 3 9 13 2
5 0 9 14 13 2
9 14 13 15 9 3 13 1 9 2
8 7 13 15 9 1 0 13 2
5 13 15 0 9 2
2 13 2
8 3 1 9 13 15 1 9 2
4 13 1 9 2
6 3 13 9 1 9 2
15 1 0 9 9 2 12 9 1 9 13 4 9 1 9 2
7 14 15 13 9 1 9 2
8 13 9 9 7 13 1 9 2
11 9 14 13 2 16 1 9 9 9 13 2
15 1 9 13 9 7 1 0 9 13 15 1 15 1 9 2
5 13 15 1 9 2
10 12 9 1 9 13 1 9 1 9 2
10 12 9 1 9 13 15 1 15 9 2
14 1 0 9 1 9 9 1 0 9 9 13 12 9 2
6 9 1 9 13 9 2
9 3 9 13 15 13 1 0 9 2
15 1 12 9 9 13 9 7 13 15 15 3 13 1 9 2
16 1 0 9 9 9 13 1 9 2 14 14 13 14 9 13 2
17 0 9 2 0 3 13 15 0 2 4 13 0 9 1 9 9 2
6 9 13 15 1 9 2
6 2 13 9 9 0 2
6 13 9 1 12 9 2
17 13 13 0 2 0 7 13 3 1 9 9 12 8 2 9 9 2
17 13 0 9 2 0 9 2 0 9 0 2 0 9 2 0 9 2
9 1 9 9 13 15 14 0 9 2
8 7 13 14 12 8 2 8 2
14 13 3 1 0 0 9 9 14 13 2 16 13 13 2
10 9 13 15 1 15 2 13 9 9 2
12 2 0 0 9 13 15 1 9 1 12 9 2
8 9 1 0 9 13 15 3 2
13 1 9 13 9 13 9 2 7 1 15 13 9 2
8 9 9 9 13 9 0 8 2
4 9 14 13 2
18 9 9 13 2 16 1 9 13 13 9 7 3 9 13 4 3 3 2
7 1 9 13 15 1 9 2
10 1 15 13 9 13 12 8 2 9 2
16 2 13 4 1 9 2 1 0 1 9 0 9 13 0 9 2
12 3 1 9 9 9 7 9 13 9 1 9 2
4 13 0 9 2
7 14 14 13 9 1 9 2
21 9 9 13 2 16 9 9 13 9 9 0 2 9 9 0 7 9 0 2 0 2
11 16 9 13 9 2 15 9 13 14 0 2
13 9 1 9 9 13 9 1 13 9 1 9 9 2
9 9 13 9 1 9 0 13 9 2
6 9 9 13 1 9 2
7 3 9 9 13 1 9 2
18 3 9 13 9 2 1 0 3 13 2 16 9 13 1 9 0 9 2
9 9 9 13 1 0 9 1 9 2
20 16 9 14 13 9 2 16 15 13 2 9 13 1 0 9 2 0 15 13 2
6 3 14 13 0 9 2
11 7 3 15 3 13 2 13 15 0 9 2
6 12 13 1 0 9 2
16 1 9 9 9 0 9 13 15 0 9 2 8 2 9 9 2
6 13 1 15 1 9 2
5 2 0 13 9 2
24 2 1 12 9 13 4 9 1 9 9 2 7 3 2 3 15 3 13 2 13 15 1 15 2
7 9 9 9 0 13 9 2
19 14 9 13 1 9 0 9 2 16 9 13 13 9 0 12 8 2 8 2
9 14 9 4 13 13 14 9 0 2
24 13 15 2 16 9 14 4 3 13 9 9 2 0 9 2 0 1 14 12 9 13 9 0 2
7 1 9 3 14 13 0 2
11 2 16 4 13 9 2 9 13 14 0 2
29 1 9 9 9 13 0 8 2 9 9 2 0 1 9 14 0 9 13 0 9 7 13 0 9 1 9 1 9 2
8 13 15 9 1 0 0 9 2
10 14 13 9 2 7 12 9 14 13 2
10 1 9 9 14 13 4 1 0 9 2
4 13 4 9 2
13 13 15 13 9 2 13 9 2 16 15 9 13 2
10 9 13 1 9 2 16 15 14 13 2
5 0 9 13 15 2
10 0 13 0 9 9 2 9 2 13 2
4 13 9 0 2
12 13 9 2 16 15 3 13 4 7 13 4 2
6 13 3 0 2 0 2
17 9 1 9 1 9 1 9 13 9 2 7 9 13 1 9 0 2
13 1 9 13 4 3 9 9 9 1 0 9 9 2
23 9 13 1 9 12 0 9 13 1 9 0 9 0 2 13 1 9 9 1 0 9 0 2
7 9 13 0 7 13 9 2
16 13 3 0 2 15 9 13 14 9 0 1 9 1 0 9 2
16 13 3 0 9 2 13 4 15 1 9 7 3 13 4 9 2
17 1 0 9 9 13 13 1 9 9 9 1 0 9 1 0 9 2
12 12 8 2 8 1 9 9 0 13 9 0 2
10 1 0 9 13 15 9 14 9 0 2
16 9 9 13 3 0 9 2 0 1 9 0 7 0 0 9 2
13 9 0 13 9 0 1 0 9 1 9 1 9 2
11 9 0 13 14 9 13 7 13 1 9 2
13 9 9 2 9 13 1 9 9 13 0 9 0 2
4 7 13 0 2
16 2 13 15 2 9 2 9 2 13 3 2 0 13 0 9 2
12 9 9 13 9 1 9 9 7 13 4 9 2
6 2 9 13 13 9 2
20 4 13 16 9 0 2 0 2 0 13 15 0 9 2 16 14 13 0 9 2
10 0 0 9 13 0 9 1 15 9 2
11 13 9 3 2 14 9 13 1 9 9 2
5 3 14 13 13 2
21 12 0 3 9 13 0 0 9 0 1 9 1 9 2 13 1 0 9 13 3 2
14 3 13 15 9 9 7 9 13 15 9 1 0 9 2
7 9 9 3 13 0 9 2
6 3 13 3 9 0 2
6 9 3 14 13 15 2
8 13 1 9 1 0 0 9 2
8 13 9 7 13 1 0 9 2
12 3 14 12 9 13 1 9 12 0 9 9 2
8 9 13 9 2 9 7 9 2
14 1 15 13 0 9 2 0 13 1 9 1 13 9 2
5 13 15 0 9 2
11 2 0 9 13 14 2 16 13 0 9 2
5 13 4 0 9 2
10 2 14 2 14 14 13 9 1 15 2
4 14 9 13 2
19 9 13 0 9 1 0 9 2 7 0 9 9 13 15 1 9 15 9 2
8 1 0 9 9 3 15 13 2
20 9 1 9 1 0 9 14 13 14 1 9 13 9 2 13 13 9 1 9 2
7 9 13 1 0 9 9 2
7 9 0 9 13 1 9 2
4 3 13 9 2
6 9 13 1 9 9 2
17 14 0 9 1 9 13 9 1 9 2 13 12 7 12 9 0 2
9 3 13 1 9 13 1 9 9 2
23 3 9 4 13 9 1 13 9 1 13 9 7 13 15 0 9 2 14 13 9 9 0 2
23 3 13 13 15 1 9 2 16 1 13 0 9 9 1 9 9 13 13 0 2 0 9 2
13 15 9 1 9 9 0 13 0 9 9 9 9 2
45 0 0 9 2 1 0 1 9 13 0 9 7 9 13 1 0 9 2 13 14 0 0 9 9 3 13 1 9 9 7 14 0 0 9 9 2 16 1 15 13 14 14 9 9 2
7 7 9 13 9 9 9 2
4 13 15 3 2
7 1 9 9 0 13 9 2
13 2 13 9 2 3 13 1 9 9 2 9 9 2
5 3 3 13 9 2
10 7 16 14 13 9 2 7 3 13 2
11 14 13 3 9 9 2 7 9 13 0 2
9 2 13 9 1 9 1 0 9 2
10 2 13 2 16 13 15 1 9 3 2
16 13 3 0 9 2 0 1 9 13 2 9 15 3 14 13 2
3 13 9 2
12 1 13 9 13 9 9 0 1 9 9 0 2
9 1 15 0 9 13 9 0 9 2
6 4 3 13 1 9 2
8 13 1 9 1 9 0 8 2
10 1 9 2 14 13 14 0 9 0 2
11 1 9 9 1 9 0 9 13 9 9 2
16 13 15 3 3 1 9 2 7 15 9 14 13 9 1 9 2
10 3 13 9 9 1 9 13 1 9 2
10 7 9 13 15 3 1 9 2 2 2
7 2 1 9 15 14 13 2
10 7 1 9 13 2 16 9 13 3 2
11 13 2 16 9 3 13 9 0 1 9 2
7 2 16 14 14 13 3 2
3 9 13 2
10 13 2 16 13 15 2 9 13 3 2
9 9 13 9 13 1 13 0 9 2
12 9 13 13 2 16 9 13 9 1 9 0 2
8 13 1 9 9 0 13 0 2
8 13 15 7 13 1 9 9 2
6 2 9 3 3 4 2
8 7 15 14 13 1 13 9 2
4 2 13 15 2
6 9 13 15 1 9 2
15 9 3 13 9 2 9 9 13 15 1 0 9 0 9 2
18 9 1 15 9 13 1 12 9 13 2 13 13 1 0 9 1 9 2
6 9 3 13 1 9 2
11 13 0 9 2 14 14 13 1 9 9 2
8 2 15 3 1 0 9 13 2
6 2 13 9 2 9 2
6 2 7 14 9 13 2
5 2 7 13 9 2
4 2 9 13 2
9 3 13 1 0 9 2 13 3 2
7 3 13 1 9 0 9 2
3 3 13 2
18 13 1 9 3 2 16 1 9 1 9 9 13 3 3 13 9 9 2
11 9 13 15 7 9 13 9 1 9 0 2
11 1 0 9 0 9 13 9 0 7 0 2
21 7 3 2 1 9 0 2 13 15 0 0 9 1 9 9 0 2 0 2 2 2
11 14 13 14 9 13 12 9 1 0 9 2
18 14 13 9 9 13 1 0 9 0 9 9 0 7 0 1 9 9 2
6 7 15 13 4 15 2
13 7 1 0 9 13 15 15 3 2 9 9 13 2
9 13 4 13 15 0 1 9 9 2
7 1 9 9 13 0 9 2
11 2 0 13 0 9 1 9 9 9 9 2
5 4 13 0 9 2
11 2 13 9 2 3 7 9 13 3 0 2
18 1 0 9 13 14 12 8 2 9 2 1 9 14 12 8 2 13 2
16 2 1 0 9 0 9 13 4 9 0 1 9 1 9 0 2
3 13 0 2
6 13 4 15 1 9 2
10 13 7 1 0 9 0 9 7 9 2
17 13 13 15 1 12 9 1 9 2 16 13 15 0 9 1 9 2
5 3 14 15 13 2
6 3 14 13 0 9 2
6 3 13 9 1 9 2
5 3 14 13 0 2
4 13 15 9 2
9 13 9 7 13 1 9 1 9 2
7 9 13 0 9 13 9 2
6 9 13 15 0 9 2
16 13 3 9 0 7 15 0 9 7 0 9 9 1 9 9 2
7 3 2 9 13 3 9 2
7 13 9 7 13 1 9 2
14 13 9 2 1 0 13 9 2 13 15 7 13 9 2
16 13 1 9 2 16 9 13 15 3 3 2 14 1 13 9 2
10 0 9 9 13 15 1 0 9 13 2
7 0 9 13 9 14 3 2
15 1 9 9 3 15 14 13 2 14 15 15 1 9 13 2
7 13 1 15 9 7 9 2
12 0 9 3 14 13 15 13 1 9 9 0 2
24 13 13 1 0 9 1 0 9 2 16 13 0 9 2 9 7 9 1 9 7 13 15 9 2
8 9 14 14 13 1 15 9 2
6 13 15 1 0 13 2
4 13 1 9 2
5 9 13 1 9 2
8 1 9 13 15 1 9 9 2
20 9 13 1 15 1 9 2 9 15 13 2 7 9 2 1 9 2 13 9 2
18 0 9 0 1 9 9 9 1 9 0 4 13 1 9 1 9 0 2
39 3 3 2 16 9 13 1 9 0 9 1 9 1 9 1 9 2 1 9 1 9 13 15 9 9 2 0 13 15 1 9 0 9 1 13 15 9 9 2
10 13 15 9 2 13 1 15 3 13 2
6 14 13 4 1 9 2
4 14 4 9 2
3 13 9 2
4 13 15 9 2
4 9 13 9 2
4 13 15 0 2
4 13 1 15 2
6 13 2 16 3 13 2
2 13 2
6 13 15 1 15 3 2
2 13 2
6 13 15 3 9 13 2
4 9 14 13 2
14 13 4 1 9 0 9 2 13 4 7 14 13 4 2
4 13 4 13 2
12 7 3 2 13 15 2 1 9 13 1 15 2
7 7 14 13 15 15 13 2
11 13 4 1 9 1 9 1 15 1 9 2
32 13 1 9 1 0 0 9 2 13 15 1 9 2 1 9 2 9 2 9 2 9 2 9 2 9 2 9 7 15 2 9 2
15 1 9 13 4 9 13 2 14 3 13 1 9 1 9 2
6 13 15 15 1 9 2
8 13 4 15 2 13 1 9 2
10 3 14 13 15 1 15 1 13 9 2
17 7 14 2 16 1 0 9 14 15 13 1 9 2 3 13 15 2
12 1 9 0 1 3 13 9 13 7 13 15 2
4 4 14 13 2
10 0 9 1 9 13 1 9 9 0 2
10 15 9 13 9 0 9 9 1 9 2
26 9 0 2 0 1 0 9 0 13 0 9 9 13 1 9 0 9 2 0 4 13 1 9 1 9 2
11 9 13 1 9 7 13 13 15 3 9 2
8 9 9 0 1 9 13 0 2
12 9 2 1 0 13 9 2 13 13 0 9 2
10 3 1 9 2 9 14 13 9 0 2
14 1 9 9 2 0 1 15 13 2 13 0 7 0 2
6 0 0 13 1 9 2
24 1 9 1 9 0 1 9 13 12 9 2 1 9 7 12 9 9 13 15 9 1 0 9 2
7 1 9 13 15 12 9 2
10 1 9 1 0 9 13 15 12 9 2
9 9 13 13 9 13 9 13 9 2
6 9 0 13 3 3 2
8 1 9 9 13 9 0 9 2
6 0 9 14 13 0 2
8 9 0 14 13 13 1 9 2
16 3 13 1 9 9 2 9 2 0 9 14 13 0 1 9 2
13 14 13 1 15 9 2 9 7 14 0 9 0 2
13 1 9 13 9 12 9 7 13 15 1 9 9 2
24 9 1 13 9 14 13 2 7 9 2 1 9 9 2 1 9 1 9 1 9 13 15 0 2
11 1 15 2 9 13 15 3 14 1 9 2
17 14 13 15 2 14 2 0 9 2 9 1 9 7 14 9 0 2
8 13 14 13 9 1 9 0 2
12 0 0 9 0 7 0 13 1 9 1 9 2
5 1 9 13 9 2
13 9 0 9 9 9 0 13 1 0 9 0 9 2
16 13 3 9 2 9 7 9 13 0 9 1 13 0 9 9 2
23 3 14 13 2 16 3 13 1 9 4 9 13 1 9 0 2 9 0 9 7 9 9 2
29 9 9 13 2 16 13 1 15 9 9 1 9 9 1 9 7 1 12 9 13 9 1 9 2 16 9 0 13 2
12 9 13 9 13 1 15 1 9 9 7 9 2
15 13 1 9 1 13 9 0 7 0 0 9 9 1 9 2
6 3 13 13 9 0 2
21 1 0 9 9 9 1 9 13 14 12 0 9 13 1 9 0 9 1 0 9 2
18 1 9 9 9 1 9 13 1 9 1 0 9 1 3 12 0 9 2
12 9 1 3 13 0 9 9 13 9 9 1 2
9 1 9 13 15 9 1 15 13 2
7 9 9 0 13 1 9 2
9 1 9 0 13 15 12 9 0 2
14 0 0 9 2 0 2 0 7 0 2 13 1 15 2
19 1 9 0 13 3 0 1 13 9 2 0 13 13 1 15 0 0 9 2
17 0 9 9 13 1 9 14 0 1 9 1 13 1 0 9 9 2
13 2 9 13 9 9 2 3 2 16 14 13 9 2
27 3 13 15 1 9 2 13 9 2 13 1 9 2 13 4 9 9 7 9 2 1 9 13 15 0 9 2
6 2 13 2 3 13 2
5 13 14 0 9 2
17 14 1 9 2 1 9 7 9 1 9 13 9 1 9 1 9 2
8 3 13 13 1 9 1 9 2
13 9 13 9 0 2 9 13 9 0 9 9 9 2
7 13 9 13 3 9 9 2
22 9 14 13 1 9 1 9 2 0 14 4 13 0 9 0 8 2 2 1 9 9 2
21 3 13 9 0 7 1 9 9 0 1 9 9 2 0 13 9 9 1 0 9 2
5 9 13 0 0 2
16 13 15 14 2 16 9 13 1 9 13 14 9 1 9 9 2
16 16 3 15 2 0 1 9 2 13 12 9 1 9 7 9 2
9 0 9 7 9 13 15 1 9 2
18 14 14 3 9 7 9 1 9 13 2 16 9 14 13 3 13 9 2
8 1 9 0 9 4 14 0 2
11 13 9 1 9 13 13 7 9 12 9 2
7 13 1 9 1 0 8 2
20 1 0 8 2 1 0 9 13 9 2 7 13 9 9 9 0 13 1 9 2
13 14 14 3 9 3 13 2 16 9 0 3 13 2
7 12 9 13 9 0 9 2
17 9 13 15 13 9 9 9 0 1 9 9 9 13 3 0 9 2
9 1 0 14 13 9 1 0 9 2
5 9 13 12 9 2
2 13 2
9 7 9 3 15 1 15 14 13 2
10 13 15 13 3 2 16 3 4 3 2
8 9 0 0 13 1 0 9 2
11 9 0 13 9 2 9 9 3 13 13 2
14 0 9 9 13 15 13 9 2 0 13 0 9 0 2
6 15 9 13 14 9 2
6 1 9 13 9 0 2
15 1 9 13 15 9 0 2 1 0 13 1 15 13 9 2
12 1 9 9 9 13 14 9 7 9 1 9 2
7 9 4 13 1 9 9 2
11 1 9 13 13 9 0 1 9 12 8 2
8 1 0 0 9 13 12 8 2
6 7 13 15 0 9 2
7 13 1 15 9 7 9 2
13 1 9 2 16 9 13 1 9 2 9 14 13 2
17 1 9 13 2 16 9 1 9 2 3 13 1 9 2 13 13 2
3 13 9 2
6 13 15 1 0 9 2
3 13 9 2
5 13 1 0 9 2
5 9 13 1 9 2
4 13 1 9 2
8 2 14 13 4 15 1 9 2
11 13 4 15 7 3 13 1 9 9 0 2
6 1 0 9 15 13 2
23 9 9 13 1 0 8 2 1 9 1 0 9 2 16 13 2 16 15 9 14 15 13 2
13 0 9 1 9 14 4 15 13 1 0 9 9 2
7 14 13 1 9 12 9 2
9 3 13 4 9 1 0 0 9 2
12 13 4 15 2 16 14 14 9 15 9 13 2
24 9 1 9 1 0 9 13 1 9 7 1 9 2 14 1 9 1 9 2 13 1 12 9 2
4 13 1 9 2
14 1 0 8 2 3 1 9 13 1 13 9 1 9 2
9 9 7 9 13 15 1 9 0 2
12 1 9 1 12 8 2 9 9 7 9 13 2
11 9 13 0 9 1 9 12 8 2 9 2
6 7 3 15 13 4 2
5 7 13 13 9 2
8 7 13 2 16 13 4 9 2
4 15 13 9 2
19 2 3 13 9 1 9 9 13 15 9 7 0 9 1 9 0 9 2 2
12 9 13 9 1 3 0 7 13 3 0 9 2
13 1 9 14 1 0 9 13 15 3 13 0 9 2
8 3 14 13 15 13 13 9 2
7 13 9 14 13 9 9 2
8 0 9 13 13 9 3 3 2
12 2 15 14 3 2 9 2 15 1 9 13 2
10 13 2 13 7 13 13 2 13 9 2
7 13 4 3 9 1 9 2
16 1 9 13 15 14 0 0 9 2 7 9 14 13 14 0 2
9 15 9 13 0 2 0 9 9 2
7 13 0 9 1 9 9 2
13 9 13 0 2 7 9 15 1 9 1 15 13 2
13 14 15 9 13 0 9 1 9 0 9 9 0 2
11 9 1 9 13 15 3 3 9 1 9 2
7 0 9 13 15 9 0 2
9 7 13 9 14 13 3 9 0 2
5 13 0 9 0 2
10 3 1 9 13 15 0 9 1 9 2
16 9 9 13 2 16 14 14 13 9 1 15 2 15 9 13 2
10 1 0 2 13 4 1 3 0 9 2
13 2 9 9 0 13 1 0 8 2 9 9 0 2
25 1 9 9 9 9 3 13 3 0 1 13 1 9 2 16 1 9 13 9 3 14 1 0 9 2
15 7 9 13 13 1 9 2 16 9 9 4 1 9 13 2
8 13 4 1 9 1 0 9 2
11 1 9 0 9 9 13 14 0 7 0 2
3 9 13 2
5 3 13 12 9 2
9 12 9 1 13 9 1 9 0 2
9 12 9 1 1 9 13 0 9 2
5 13 2 16 13 2
14 15 14 13 1 0 9 7 9 2 7 13 9 0 2
17 1 9 9 0 2 0 0 9 13 1 13 9 2 13 15 3 2
7 7 9 9 3 9 13 2
5 14 13 1 3 2
7 13 1 13 0 9 0 2
11 1 0 9 13 15 0 9 13 1 9 2
7 1 9 0 9 13 3 2
11 0 9 1 9 0 13 0 9 1 9 2
6 9 13 1 9 9 2
9 13 0 1 3 0 9 0 9 2
7 3 13 7 13 1 9 2
14 1 0 9 14 13 15 1 13 1 9 1 0 9 2
7 0 9 13 1 0 9 2
14 1 9 13 9 9 9 7 9 2 9 13 9 9 2
12 3 14 13 9 1 9 2 0 13 0 9 2
7 9 13 0 9 0 9 2
10 7 1 13 0 9 9 13 15 9 2
8 2 3 13 3 9 9 9 2
8 13 1 9 7 0 9 0 2
8 0 9 13 13 9 1 9 2
18 9 0 1 9 13 3 2 16 1 0 9 9 9 14 4 0 9 2
17 1 9 0 9 13 15 1 13 9 2 15 9 14 13 9 0 2
10 9 9 13 3 0 9 13 1 9 2
16 15 15 13 0 9 2 0 15 13 9 2 7 13 14 9 2
6 13 4 14 1 9 2
7 9 1 0 9 13 0 2
11 14 13 2 3 14 13 4 15 1 9 2
8 9 0 13 14 1 0 9 2
9 9 9 13 9 14 1 9 0 2
14 12 13 9 9 2 7 15 9 13 15 1 9 0 2
8 9 13 3 1 9 9 0 2
16 9 0 13 14 13 1 0 9 7 9 0 13 1 9 9 2
9 14 13 4 2 14 13 14 9 2
12 0 9 13 14 0 9 13 13 9 0 9 2
21 3 14 13 15 9 0 0 9 1 9 9 1 9 0 9 7 9 1 0 9 2
6 1 3 13 1 9 2
5 0 9 14 13 2
7 7 15 3 13 1 9 2
5 15 14 13 9 2
5 16 14 13 9 2
7 16 0 13 9 0 9 2
7 15 9 13 15 15 9 2
28 9 9 2 3 1 15 0 2 13 3 1 9 2 13 3 9 0 9 2 9 9 2 13 3 0 2 0 2
4 9 13 13 2
7 3 13 2 16 13 3 2
16 16 13 2 3 2 3 14 15 9 14 13 2 3 13 9 2
8 1 9 14 13 9 3 3 2
10 14 13 9 2 16 15 1 9 13 2
4 3 13 9 2
13 7 1 0 9 2 3 13 15 1 0 0 9 2
16 13 9 14 13 7 13 9 2 7 14 3 3 13 1 9 2
18 1 0 9 2 0 13 9 9 2 13 0 9 13 0 13 15 9 2
7 14 2 13 4 0 9 2
6 9 3 3 14 13 2
9 13 0 9 2 7 3 15 13 2
13 7 14 14 13 2 1 0 9 13 0 9 0 2
11 13 15 1 9 7 1 0 9 13 9 2
12 3 13 15 2 16 14 13 9 1 0 9 2
18 1 0 9 13 15 13 0 2 7 14 13 2 3 9 4 3 13 2
11 3 13 9 1 9 1 15 9 2 9 2
12 0 13 14 0 9 2 7 7 13 1 9 2
14 3 14 13 2 16 13 14 1 0 9 0 7 0 2
5 14 13 0 9 2
13 9 13 2 13 1 9 2 7 3 14 13 3 2
14 7 0 9 0 0 9 7 0 9 9 13 14 13 2
13 1 0 9 13 0 9 1 0 2 3 0 9 2
19 16 13 9 2 13 14 3 13 9 2 7 15 3 13 3 9 2 13 2
8 9 13 0 9 9 9 0 2
26 1 12 9 13 14 9 7 9 7 13 1 0 9 0 0 9 2 13 14 1 9 9 7 14 9 2
10 3 13 14 12 8 2 8 9 0 2
7 13 15 1 9 9 9 2
12 1 0 9 13 2 16 1 12 9 13 9 2
12 0 2 1 9 2 13 0 7 13 0 9 2
30 1 9 0 13 12 9 2 12 9 1 0 9 2 0 13 0 7 0 2 16 0 9 14 13 1 15 0 13 9 2
11 9 14 13 7 0 9 2 7 0 9 2
9 1 15 0 7 9 14 13 9 2
9 7 13 15 9 2 16 15 13 2
4 13 1 0 2
13 1 15 9 13 3 9 9 2 0 13 1 9 2
31 9 1 0 9 13 2 16 9 9 13 0 7 0 2 7 9 7 9 13 9 7 13 9 7 13 15 1 9 1 9 2
15 1 9 2 9 3 13 15 1 9 2 13 14 0 9 2
16 9 7 2 16 13 1 15 0 9 2 13 0 2 1 9 2
7 4 13 9 0 7 0 2
12 1 9 9 13 9 0 1 9 9 9 9 2
7 3 14 13 1 15 9 2
9 3 13 15 1 9 1 0 9 2
10 1 9 13 2 16 13 15 0 9 2
6 13 4 15 0 9 2
7 1 9 9 13 4 3 2
16 1 9 9 0 2 9 1 0 9 13 1 9 9 1 9 2
6 3 13 13 9 9 2
10 9 9 13 9 0 1 9 0 9 2
20 1 9 0 9 13 2 16 13 9 0 9 1 9 4 13 0 0 9 0 2
14 14 13 2 3 13 9 2 16 14 13 0 9 0 2
9 13 15 1 0 9 1 9 9 2
6 12 13 15 1 9 2
6 9 4 13 1 9 2
5 1 9 9 13 2
13 13 4 9 0 9 2 7 9 13 15 1 9 2
14 13 4 9 1 0 9 1 9 7 13 4 1 9 2
6 13 4 14 13 15 2
19 3 14 13 4 15 14 0 2 16 13 4 1 15 14 0 7 13 9 2
6 13 1 13 0 9 2
8 13 4 9 2 16 13 9 2
7 14 13 4 13 9 9 2
14 13 15 1 9 13 2 16 9 13 9 1 9 0 2
6 9 13 4 1 13 2
10 0 1 15 9 14 13 1 0 9 2
36 0 9 13 15 2 16 15 9 1 0 9 0 9 13 15 13 0 2 16 1 9 9 9 13 15 14 3 0 9 2 0 13 9 1 9 2
5 9 9 14 13 2
11 9 13 12 9 7 13 4 1 9 0 2
15 9 13 1 13 9 0 2 0 4 3 13 1 0 9 2
12 9 9 3 13 1 9 13 9 9 0 9 2
14 1 9 0 13 14 0 9 1 0 9 0 2 0 2
12 13 14 9 1 9 1 9 2 9 7 9 2
15 13 15 15 2 16 1 0 9 9 13 9 14 0 9 2
22 14 13 0 9 9 2 9 9 9 2 9 9 2 0 9 14 13 1 9 1 9 2
10 9 9 14 3 14 13 15 1 9 2
8 13 15 14 1 9 1 9 2
7 9 9 13 9 1 9 2
15 2 16 13 9 1 9 1 9 2 9 14 15 14 13 2
9 13 9 0 9 3 7 13 13 2
12 3 1 0 9 1 9 14 13 15 9 9 2
7 3 13 15 9 7 4 2
13 1 9 4 13 1 0 9 2 0 9 14 13 2
15 13 15 3 14 9 0 1 9 2 9 0 7 9 9 2
13 1 9 0 13 15 1 0 9 4 13 9 0 2
14 1 0 9 9 0 7 0 1 9 0 1 9 13 2
11 13 15 14 9 9 13 7 13 1 9 2
14 3 14 9 9 9 13 2 16 1 9 13 0 9 2
9 0 9 9 0 13 9 9 0 2
19 3 1 13 1 0 9 9 2 9 9 7 9 0 13 15 1 0 9 2
12 13 1 15 9 12 9 9 0 1 9 9 2
14 1 0 12 9 12 13 1 9 0 1 9 7 9 2
10 14 9 0 3 14 13 1 9 0 2
5 9 13 9 0 2
8 9 13 9 0 9 0 9 2
15 12 9 0 9 13 14 3 1 9 9 0 1 9 0 2
7 9 1 15 13 1 9 2
10 0 9 0 13 1 13 9 1 9 2
12 1 9 9 13 1 9 14 12 8 2 9 2
13 9 3 15 13 2 7 9 0 9 13 14 0 2
9 1 9 13 13 0 9 9 0 2
11 13 14 13 1 0 9 0 0 9 0 2
16 1 9 13 14 12 9 9 2 3 12 1 15 13 13 9 2
8 9 13 9 9 13 1 0 2
20 9 0 9 13 14 15 13 2 13 14 2 16 9 4 13 9 9 1 9 2
7 1 15 13 9 7 9 2
14 13 0 9 4 3 13 13 1 9 1 13 0 9 2
13 9 13 1 9 2 16 13 9 1 9 1 9 2
16 16 13 15 1 9 2 14 13 1 15 7 9 2 7 9 2
12 14 13 2 16 13 1 9 1 9 0 9 2
5 13 15 12 9 2
10 13 9 13 15 0 9 13 0 9 2
13 2 0 9 13 9 1 9 13 13 1 13 9 2
18 9 13 0 9 7 3 13 15 1 9 2 13 1 0 9 0 9 2
8 13 15 9 1 9 7 9 2
8 4 13 1 13 9 9 0 2
3 14 13 2
7 9 13 15 1 9 9 2
4 13 14 9 2
9 9 13 15 1 9 9 2 2 2
5 1 9 13 9 2
5 2 13 3 9 2
11 13 1 12 0 9 2 0 15 14 13 2
8 13 2 16 0 9 15 13 2
7 9 13 1 9 9 9 2
7 14 13 15 9 1 9 2
5 3 13 0 9 2
11 2 4 3 13 2 16 9 15 14 13 2
8 9 9 13 15 1 9 0 2
7 13 15 1 9 7 9 2
6 2 0 13 9 9 2
4 9 13 9 2
12 9 15 13 2 7 15 0 15 14 14 13 2
22 14 13 2 14 9 13 9 0 2 0 13 14 13 9 1 9 2 16 13 15 0 2
15 9 1 0 9 13 13 9 2 13 9 2 13 0 9 2
13 13 9 1 9 9 0 2 0 2 0 2 0 2
4 13 15 9 2
5 3 3 13 9 2
3 9 13 2
14 0 1 9 13 15 1 9 2 16 13 1 0 9 2
13 7 13 9 9 7 9 13 9 2 9 2 9 2
7 13 4 1 9 0 9 2
10 0 9 3 13 0 9 9 13 9 2
16 0 9 0 9 9 0 13 1 9 0 2 14 15 13 9 2
8 13 15 14 12 9 1 9 2
5 9 13 15 14 2
5 13 2 13 9 2
5 1 15 9 13 2
6 3 13 9 7 9 2
5 13 2 16 13 2
5 7 9 14 13 2
5 14 15 14 13 2
8 1 9 13 1 15 1 9 2
6 3 13 1 9 9 2
12 9 3 13 2 13 1 9 1 0 0 9 2
6 1 9 13 0 9 2
17 9 13 7 13 15 1 9 2 1 15 2 3 2 13 15 9 2
9 13 3 2 13 9 1 0 9 2
7 9 13 3 7 14 13 2
4 9 13 3 2
24 9 1 9 13 2 16 1 0 9 13 4 14 9 0 9 2 7 9 1 9 7 0 9 2
8 2 13 9 2 9 2 2 2
5 0 9 13 9 2
14 4 13 14 9 0 9 0 2 1 0 3 15 13 2
12 1 3 13 9 2 14 1 9 13 0 9 2
9 15 9 13 1 0 13 0 9 2
9 9 13 15 1 9 1 9 9 2
6 9 14 13 1 9 2
10 1 0 9 13 2 16 9 14 13 2
11 9 13 1 9 7 13 1 9 1 9 2
5 0 14 13 15 2
8 14 2 1 0 9 14 13 2
16 9 13 1 9 7 13 9 2 0 15 1 13 13 1 9 2
8 7 1 9 13 9 9 9 2
17 9 9 2 1 0 3 13 4 9 2 13 4 12 8 2 9 2
8 2 7 3 9 13 14 13 2
7 2 14 13 15 0 9 2
7 7 14 9 13 1 9 2
3 9 13 2
2 13 2
6 2 13 4 15 13 2
4 2 13 9 2
11 2 0 9 13 1 9 2 9 9 0 2
14 9 13 15 1 9 2 13 9 7 13 3 1 9 2
10 1 9 12 13 9 2 9 2 9 2
3 3 13 2
6 2 13 15 15 3 2
15 2 13 4 1 0 9 12 9 7 13 15 15 3 0 2
10 2 7 13 4 14 9 1 15 9 2
12 14 15 13 2 7 14 13 14 9 1 9 2
9 2 7 13 2 9 13 15 3 2
16 14 4 14 13 1 9 0 2 0 13 15 3 1 0 9 2
7 13 0 9 1 9 0 2
8 2 7 9 15 1 15 13 2
11 3 1 14 12 9 4 13 9 9 0 2
13 1 0 9 9 13 15 0 9 0 9 9 0 2
5 9 0 9 13 2
7 2 1 9 13 4 9 2
7 2 1 9 13 13 3 2
8 15 3 13 2 15 3 13 2
10 9 13 1 15 7 13 15 1 9 2
9 0 9 1 15 3 13 2 2 2
4 9 15 13 2
13 13 14 4 9 9 7 9 1 0 9 9 9 2
20 2 14 13 9 2 16 1 9 2 16 13 9 2 9 13 9 1 9 9 2
6 2 13 3 9 0 2
9 2 3 13 9 9 1 12 9 2
12 2 9 13 13 9 14 1 9 1 9 0 2
13 7 1 0 9 13 1 9 14 12 9 1 9 2
5 9 13 15 3 2
6 9 13 15 1 9 2
11 9 13 15 1 9 7 13 15 0 9 2
7 13 15 9 1 13 9 2
9 2 9 13 7 13 15 1 9 2
8 9 9 0 13 1 0 9 2
8 0 9 9 13 15 1 9 2
9 3 3 13 15 13 15 7 13 2
11 14 1 9 13 1 0 9 1 13 9 2
15 16 13 9 2 9 13 2 16 13 15 1 15 1 9 2
12 9 7 9 13 1 9 0 9 1 9 9 2
5 3 13 15 15 2
14 16 0 9 13 2 16 9 13 13 9 2 9 13 2
21 1 9 9 3 3 13 2 9 13 13 0 1 13 15 3 3 1 9 0 9 2
26 2 9 0 13 15 1 0 9 1 9 13 2 7 0 0 9 1 9 9 9 13 9 9 1 9 2
19 0 9 13 9 1 9 9 0 1 9 2 0 13 15 1 13 0 9 2
13 1 0 9 13 3 1 9 1 9 0 9 0 2
18 16 1 9 13 15 9 1 9 0 9 2 9 13 15 1 0 9 2
16 13 9 1 9 13 9 2 7 9 9 0 2 7 14 9 2
5 13 9 0 9 2
5 13 15 0 9 2
15 2 1 9 13 4 1 9 0 2 0 13 15 1 9 2
7 9 0 13 0 9 0 2
9 9 13 9 1 0 9 0 9 2
8 9 3 13 15 1 9 9 2
29 13 1 0 9 13 1 0 9 9 9 0 1 0 2 0 9 2 0 13 9 1 9 13 1 0 9 1 9 2
23 14 3 9 13 13 9 9 9 9 9 7 12 0 9 7 9 13 15 1 0 9 9 2
11 9 0 9 9 0 13 1 9 0 9 2
6 13 0 9 2 2 2
4 13 0 9 2
6 13 4 15 2 2 2
9 3 13 2 13 1 9 0 9 2
5 2 13 4 15 2
5 14 4 0 9 2
6 13 9 7 13 15 2
4 2 13 15 2
5 13 4 1 15 2
6 14 13 14 1 15 2
9 2 3 14 13 4 15 1 9 2
4 9 15 13 2
7 13 9 7 13 1 9 2
20 9 14 13 9 2 14 13 9 2 14 13 3 0 9 7 14 13 13 9 2
11 13 4 14 9 2 16 13 1 15 9 2
6 9 13 3 3 0 2
8 13 4 14 13 1 0 9 2
15 9 13 3 2 7 1 9 9 13 15 9 9 7 9 2
10 9 9 9 13 1 9 1 0 9 2
12 13 9 1 9 7 13 1 9 9 13 9 2
5 9 13 1 9 2
5 13 4 1 9 2
12 14 13 0 9 2 0 9 13 15 1 9 2
4 13 4 9 2
6 2 3 9 13 13 2
6 9 3 13 15 13 2
18 12 9 13 1 13 9 2 0 13 15 13 9 0 1 9 1 9 2
6 1 0 9 13 9 2
4 13 4 9 2
6 14 13 4 3 9 2
11 2 13 2 16 14 13 4 15 13 9 2
12 2 14 13 9 2 16 15 15 13 2 2 2
7 2 4 13 13 0 9 2
3 2 13 2
5 13 4 15 9 2
3 13 9 2
3 13 4 2
11 13 13 4 2 16 9 13 15 1 9 2
5 13 4 0 9 2
5 2 9 15 13 2
5 13 4 9 9 2
11 1 0 9 13 4 2 16 13 15 9 2
13 13 4 1 9 1 9 2 13 15 1 0 9 2
10 13 4 9 9 7 13 4 1 9 2
12 13 4 3 12 9 7 13 4 15 1 9 2
5 13 4 1 9 2
8 4 13 9 9 2 0 13 2
15 9 13 9 9 0 2 1 0 13 9 1 15 0 9 2
9 3 13 9 7 13 15 1 9 2
10 9 13 15 12 9 7 13 2 2 2
6 3 13 1 15 9 2
18 9 13 1 0 9 13 3 0 9 9 9 2 0 3 3 13 9 2
14 9 7 9 13 14 9 2 3 13 1 0 9 9 2
7 13 15 13 15 1 9 2
7 13 9 13 1 0 9 2
10 9 1 9 9 13 9 0 1 9 2
6 9 14 13 1 9 2
7 9 8 2 13 0 9 2
7 13 1 15 13 0 9 2
9 1 9 12 0 9 13 0 9 2
15 13 9 9 0 2 0 13 1 9 9 9 7 9 9 2
20 9 13 0 9 2 13 13 9 7 9 2 0 9 13 0 9 1 13 9 2
8 9 13 1 9 7 9 9 2
9 1 12 9 3 13 0 0 9 2
12 1 12 9 13 1 9 14 1 13 9 0 2
9 9 9 4 13 1 12 9 9 2
11 13 2 16 3 13 15 1 0 9 9 2
14 1 9 0 1 8 2 1 9 13 15 13 12 9 2
16 9 9 13 14 13 2 14 9 9 0 13 9 3 1 9 2
11 9 13 0 9 1 9 1 9 7 9 2
15 9 9 0 13 9 1 9 0 1 9 9 2 9 9 2
23 2 1 0 13 9 9 0 0 0 9 9 2 7 0 9 1 0 9 13 1 9 9 2
9 1 0 9 13 15 9 9 9 2
17 1 15 13 13 15 9 9 1 9 2 9 0 2 0 7 0 2
12 0 0 2 0 9 4 13 1 0 9 0 2
9 1 0 9 9 0 13 3 3 2
11 9 9 9 0 13 1 9 1 0 9 2
11 9 0 9 1 9 13 0 9 0 9 2
7 13 9 1 9 9 0 2
11 1 0 9 9 1 9 9 13 0 9 2
9 13 1 9 9 13 9 1 9 2
11 1 0 14 9 0 13 14 9 9 0 2
11 9 0 13 7 14 12 9 1 0 9 2
5 13 4 14 9 2
19 9 0 9 0 13 1 13 9 7 13 0 9 1 0 9 0 1 9 2
10 0 1 0 9 13 16 14 1 9 2
8 1 9 9 4 13 0 9 2
9 13 15 15 1 9 0 1 9 2
13 13 14 13 2 16 13 4 1 9 0 0 9 2
6 9 13 15 1 9 2
15 9 9 13 2 16 1 9 0 13 9 13 0 0 9 2
20 1 9 13 15 9 1 9 1 9 1 0 0 9 9 0 1 9 7 9 2
7 9 13 9 13 9 9 2
7 13 9 14 1 9 0 2
11 1 0 9 13 14 13 1 9 0 9 2
8 0 9 0 13 12 0 9 2
8 14 1 9 9 13 9 0 2
19 16 13 9 9 13 13 9 2 13 14 13 0 9 13 15 1 9 9 2
7 3 3 13 15 9 9 2
13 13 13 0 9 2 14 9 0 13 0 9 0 2
7 0 9 0 13 9 0 2
7 13 0 2 0 9 9 2
6 0 9 9 14 13 2
16 3 1 9 1 9 1 9 13 9 2 1 0 13 12 9 2
13 13 0 14 9 2 0 13 15 1 13 0 9 2
14 3 15 13 7 13 2 14 15 9 14 13 0 3 2
14 16 3 13 4 15 1 9 0 2 13 4 0 9 2
20 1 9 0 2 14 1 9 9 2 13 9 13 1 9 9 13 1 9 9 2
16 9 9 0 4 13 1 9 9 1 9 13 9 0 9 0 2
16 0 9 0 13 9 0 1 9 9 0 9 1 9 9 0 2
20 14 0 9 1 9 1 9 9 13 9 9 9 7 13 1 9 0 9 9 2
13 2 0 9 9 13 1 9 0 0 9 1 9 2
6 13 0 9 1 9 2
8 9 13 1 9 13 9 0 2
10 13 1 9 2 13 15 13 9 0 2
14 1 13 9 7 13 15 1 9 1 0 9 13 9 2
8 9 4 13 1 13 9 0 2
6 13 9 9 1 9 2
6 9 0 13 15 3 2
6 9 0 13 1 9 2
8 14 1 0 9 13 15 9 2
7 14 9 14 13 15 9 2
4 3 13 9 2
6 0 9 1 9 13 2
7 3 13 13 9 1 9 2
6 14 13 15 9 9 2
6 9 13 15 1 9 2
22 9 13 1 9 7 13 3 1 9 13 15 1 9 7 13 9 2 1 0 4 13 2
3 3 13 2
15 16 13 4 1 0 9 2 13 4 15 14 13 15 9 2
12 13 2 16 9 13 15 2 13 15 0 9 2
15 3 15 9 13 2 3 15 13 7 3 0 9 13 9 2
13 13 2 16 3 13 15 2 7 15 9 14 13 2
18 13 14 3 2 16 9 14 13 2 9 13 2 7 9 14 15 13 2
5 9 4 1 9 2
5 13 15 13 3 2
11 9 2 13 2 13 15 2 14 0 9 2
5 14 15 14 13 2
4 14 13 15 2
6 13 14 9 0 9 2
6 3 13 9 9 9 2
6 9 13 1 0 9 2
7 13 13 15 9 14 3 2
18 9 9 2 9 13 2 16 9 0 1 0 9 13 1 0 9 9 2
7 9 15 1 0 9 13 2
13 13 4 0 9 2 0 9 2 0 9 2 2 2
8 13 15 14 3 0 2 2 2
13 1 9 0 1 3 0 9 14 13 4 15 13 2
4 13 15 9 2
11 2 13 4 9 2 9 14 0 13 0 2
5 2 14 0 13 2
10 0 9 9 13 1 9 12 9 1 2
10 1 9 9 13 4 13 14 12 9 2
9 0 1 9 9 13 9 13 9 2
12 0 1 9 9 13 1 9 9 7 13 9 2
15 9 1 9 1 13 3 9 0 14 13 9 13 0 9 2
20 9 13 1 8 2 9 13 2 16 1 0 8 2 13 15 1 9 9 9 2
8 8 9 9 13 1 9 9 2
22 1 0 1 9 8 2 9 13 13 9 9 13 1 9 2 16 13 9 1 9 0 2
20 13 3 12 9 2 3 1 12 9 1 9 2 13 15 14 1 0 9 9 2
7 1 9 14 13 0 9 2
9 1 0 9 13 1 0 9 9 2
10 0 0 9 13 0 9 1 9 9 2
11 3 13 1 9 9 7 13 9 1 9 2
17 13 0 9 1 9 2 13 0 9 9 2 13 9 1 0 9 2
11 13 15 9 9 2 13 4 13 1 9 2
4 13 1 9 2
14 1 15 13 13 0 0 9 14 1 9 14 1 9 2
7 1 9 13 15 1 9 2
12 0 9 13 9 2 13 0 9 1 0 9 2
21 1 13 9 0 9 1 9 13 15 15 13 13 1 9 9 2 13 9 9 9 2
16 14 1 0 9 13 14 9 13 9 9 13 2 16 3 13 2
15 3 9 13 9 1 9 2 0 13 9 2 13 1 9 2
12 0 9 13 15 0 1 9 0 9 1 9 2
8 9 9 0 13 9 0 9 2
8 13 15 1 15 0 9 9 2
5 9 13 15 3 2
5 9 13 15 9 2
7 1 9 13 15 0 9 2
9 9 3 9 13 15 1 9 0 2
12 9 9 13 1 15 9 13 15 1 0 9 2
5 9 13 1 9 2
5 13 15 3 13 2
5 9 13 15 9 2
13 1 0 9 13 4 15 0 9 7 13 4 9 2
7 9 1 9 13 0 9 2
21 14 13 4 15 3 2 16 1 0 9 0 13 14 9 2 7 3 13 1 9 2
13 15 9 13 13 9 9 2 7 9 9 1 9 2
15 1 12 9 1 9 0 13 0 9 1 9 9 1 9 2
6 3 9 13 15 9 2
15 9 13 1 9 0 9 2 7 9 9 13 12 9 9 2
17 1 9 13 9 1 9 0 12 9 0 2 1 0 13 12 9 2
25 2 13 4 14 12 9 2 3 13 9 7 14 13 4 14 1 9 2 1 0 13 0 9 0 2
9 13 0 9 9 7 13 1 9 2
17 13 9 0 9 1 9 9 13 9 1 9 7 13 1 0 9 2
4 9 13 0 2
8 9 13 1 13 15 1 9 2
5 9 13 9 9 2
9 9 13 1 0 9 9 9 0 2
15 9 3 13 1 0 9 7 13 9 1 0 9 1 9 2
11 9 14 13 15 13 9 2 16 13 9 2
6 9 9 13 1 9 2
11 3 13 9 3 2 3 13 15 9 9 2
14 9 13 9 9 2 13 1 9 9 13 9 2 13 2
18 13 9 13 2 0 9 13 1 9 2 16 13 15 1 13 0 9 2
6 3 15 13 9 9 2
12 9 13 9 1 9 2 3 13 15 7 13 2
13 9 13 15 1 9 2 16 13 14 1 0 9 2
10 1 9 13 15 0 0 2 0 9 2
4 13 14 9 2
8 3 14 14 13 3 3 0 2
10 14 13 1 0 9 13 9 1 9 2
17 9 13 15 2 16 9 9 3 13 1 9 2 15 15 14 13 2
4 12 13 0 2
7 9 13 9 1 9 9 2
17 4 13 0 9 9 1 0 9 2 7 1 15 13 12 0 9 2
11 9 0 9 7 9 9 0 13 0 9 2
15 2 14 9 13 13 9 9 2 0 1 9 13 1 9 2
5 2 14 13 9 2
38 13 1 9 2 16 9 13 15 1 9 2 16 1 0 9 13 9 0 9 7 16 14 13 0 9 13 9 2 13 9 2 13 9 0 7 13 9 2
6 0 9 14 13 0 2
4 0 13 9 2
8 9 1 9 13 13 1 9 2
14 15 9 13 0 13 9 0 9 1 0 9 1 9 2
7 9 13 9 9 9 9 2
9 9 9 0 13 1 9 9 9 2
23 9 9 13 1 9 2 16 1 0 9 4 13 13 9 0 2 7 14 13 14 15 9 2
7 9 13 7 3 9 13 2
7 9 4 13 1 9 9 2
12 3 1 0 9 9 0 13 14 1 0 9 2
13 0 9 13 13 9 1 0 9 9 7 9 9 2
11 1 15 9 0 4 0 9 1 13 9 2
4 13 12 9 2
8 13 14 9 9 1 0 9 2
12 9 1 9 13 9 8 2 9 9 9 9 2
10 9 1 0 9 0 9 14 15 13 2
5 3 9 9 13 2
8 0 9 4 0 1 12 9 2
25 0 9 9 13 2 16 9 1 0 9 14 4 13 1 9 2 1 0 9 13 9 13 9 0 2
20 3 1 15 13 15 14 0 9 2 0 1 0 9 4 13 1 9 1 9 2
12 9 1 9 13 9 0 9 7 13 1 9 2
11 9 9 7 9 13 9 2 9 7 9 2
8 15 14 4 13 9 0 9 2
12 16 13 9 1 9 2 13 1 9 1 9 2
16 16 13 1 9 9 9 2 9 9 13 9 0 7 13 9 2
6 3 9 13 1 9 2
7 0 9 13 15 1 9 2
17 13 9 9 2 0 13 0 9 2 7 13 14 3 0 1 9 2
12 13 3 14 12 9 0 2 0 13 13 9 2
6 0 9 13 1 9 2
9 0 0 9 14 13 13 9 9 2
5 9 13 1 9 2
8 1 9 0 9 13 14 0 2
6 9 13 15 14 0 2
15 13 15 2 16 15 9 1 9 9 1 9 14 4 13 2
11 1 15 13 1 9 9 2 9 7 9 2
7 3 13 1 12 9 12 2
28 14 1 13 9 2 0 9 13 13 0 3 9 1 9 12 9 7 9 12 9 1 9 7 12 1 9 0 2
7 14 0 9 4 1 9 2
21 0 9 1 9 1 9 9 1 9 1 9 13 1 9 9 13 9 0 9 9 2
14 13 3 9 9 0 9 9 13 14 3 9 9 0 2
14 13 2 16 1 9 9 14 13 1 9 1 0 9 2
9 13 1 9 2 13 15 1 9 2
10 3 9 9 13 13 0 9 1 9 2
7 9 1 9 9 0 13 2
11 1 0 9 0 1 9 14 13 13 9 2
11 13 9 2 16 13 15 15 1 0 9 2
12 13 1 9 9 1 9 13 9 1 0 9 2
8 13 9 9 1 9 1 9 2
10 0 9 13 14 1 0 9 0 9 2
7 1 0 9 13 0 9 2
11 9 13 7 13 9 1 0 0 9 0 2
9 9 0 9 13 0 9 9 0 2
13 9 9 1 0 9 13 14 1 9 0 9 0 2
8 2 0 9 0 13 9 9 2
5 9 4 9 0 2
6 2 14 13 0 9 2
4 9 13 9 2
17 2 14 13 15 2 16 9 13 1 9 14 13 1 15 9 0 2
16 1 9 13 14 9 9 9 2 0 1 0 9 13 0 9 2
15 1 9 9 13 9 13 9 2 0 13 9 7 15 9 2
17 9 0 13 15 13 9 2 16 9 1 0 9 14 13 12 9 2
5 9 0 13 9 2
13 7 12 1 12 0 9 14 13 13 15 1 9 2
8 13 2 16 13 15 9 9 2
11 0 9 13 9 9 0 1 9 0 9 2
9 1 9 9 13 15 3 0 9 2
12 1 0 9 1 9 0 9 13 14 12 9 2
24 1 9 0 9 13 1 9 0 2 0 9 0 2 1 0 9 13 1 9 13 1 9 9 2
10 0 9 13 3 14 0 0 9 9 2
18 1 0 9 9 0 9 13 9 9 9 9 0 7 0 1 9 0 2
4 13 9 0 2
14 3 13 3 1 9 12 9 7 13 1 9 0 9 2
5 9 14 9 13 2
10 13 4 1 9 7 14 13 4 9 2
15 1 9 2 1 0 9 9 2 13 1 9 9 0 9 2
15 1 9 0 13 9 0 2 3 1 0 9 13 15 9 2
7 13 7 13 15 14 9 2
14 1 9 0 8 2 13 1 9 2 16 3 13 9 2
7 1 9 13 4 14 9 2
13 3 13 2 16 0 9 13 13 1 9 7 9 2
11 1 0 13 2 16 13 9 13 1 9 2
10 3 3 13 15 14 1 9 0 9 2
12 3 14 1 9 13 13 1 9 9 9 9 2
24 13 15 14 0 9 13 1 9 9 7 1 9 13 15 1 9 1 13 9 13 1 9 0 2
5 9 9 14 13 2
7 0 9 13 1 9 9 2
9 0 9 4 13 1 9 1 9 2
8 12 9 13 13 1 9 9 2
9 3 13 15 0 2 0 9 9 2
8 13 4 9 2 9 4 13 2
15 9 13 15 1 15 7 13 2 3 13 9 1 0 9 2
19 13 1 9 9 2 13 9 9 2 0 13 15 1 15 1 9 7 9 2
5 3 9 13 3 2
8 13 2 13 4 0 9 9 2
26 1 9 13 9 0 9 1 9 0 13 9 2 16 1 13 0 9 0 13 1 0 9 0 9 0 2
13 9 0 14 4 13 3 13 7 13 3 13 9 2
20 13 0 9 13 0 1 0 9 9 13 1 9 0 2 1 8 2 9 9 2
18 9 13 1 0 9 1 0 2 0 9 0 1 9 1 9 1 9 2
31 9 9 0 1 9 9 9 2 13 15 9 9 2 13 1 0 9 9 9 1 9 2 14 9 13 15 1 13 15 9 2
18 13 15 2 16 13 15 0 9 9 7 9 9 9 9 1 9 0 2
10 13 15 1 9 7 13 15 1 9 2
6 9 1 9 15 13 2
19 1 9 13 1 9 2 13 3 7 1 9 9 13 15 2 9 15 13 2
18 2 9 2 14 13 4 9 1 9 2 3 13 14 4 13 1 15 2
9 3 9 9 13 9 1 0 9 2
8 9 7 9 13 13 9 0 2
5 3 13 1 9 2
12 3 15 13 4 2 16 14 3 14 13 9 2
16 3 14 13 14 4 15 13 15 3 1 9 2 16 13 0 2
18 13 4 2 3 13 9 1 0 9 2 13 2 16 13 3 1 9 2
3 9 13 2
3 9 13 2
8 7 14 9 13 1 0 9 2
11 14 13 14 0 9 0 2 9 1 0 2
6 7 9 13 4 9 2
3 9 13 2
7 13 2 3 9 13 9 2
5 13 3 9 9 2
27 1 9 2 0 3 13 0 9 2 13 12 9 9 2 12 9 7 12 9 0 2 1 9 9 1 9 2
11 0 9 13 1 9 0 9 12 0 9 2
15 7 0 9 9 13 4 13 14 1 3 13 9 13 9 2
10 13 13 2 16 1 0 9 13 3 2
4 3 13 9 2
12 0 9 9 13 15 1 9 1 13 9 0 2
19 9 9 9 2 9 9 0 2 13 9 1 9 0 1 9 0 9 0 2
17 9 9 9 13 13 15 3 0 1 9 2 14 13 3 15 9 2
10 9 13 1 9 9 13 15 1 0 2
20 9 9 1 9 1 0 9 9 13 3 2 7 15 9 13 4 13 1 0 2
22 9 9 9 3 1 15 9 13 14 0 2 7 3 1 9 1 0 9 13 14 3 2
8 1 0 9 9 13 15 3 2
5 0 9 13 9 2
22 9 9 1 13 0 9 13 3 13 13 9 2 0 14 13 1 15 1 13 0 9 2
17 1 9 0 13 9 1 0 9 1 9 2 1 0 13 0 9 2
6 13 9 1 0 9 2
18 9 13 3 0 0 9 1 9 0 9 2 1 0 13 9 0 9 2
11 9 1 9 13 9 7 13 15 9 9 2
10 1 9 0 9 1 9 14 13 0 2
12 3 13 15 1 9 0 9 1 0 9 0 2
14 0 9 14 13 1 9 2 13 9 9 7 0 9 2
12 1 0 9 9 9 13 15 3 0 9 9 2
10 0 9 0 13 1 0 9 12 9 2
13 7 16 9 0 9 14 13 2 13 4 15 13 2
12 13 9 13 13 15 9 0 2 13 0 9 2
8 0 9 4 13 0 9 9 2
11 13 4 2 16 13 4 9 1 0 9 2
4 9 3 13 2
10 3 3 0 9 13 9 9 1 9 2
14 13 0 9 2 1 0 0 1 9 13 14 12 9 2
10 1 9 0 0 9 9 13 12 8 2
11 9 0 0 9 1 0 9 13 12 8 2
10 1 9 12 9 13 15 1 12 8 2
19 13 2 16 9 13 9 1 9 9 9 9 1 9 9 0 2 13 9 2
24 3 9 0 13 4 3 13 2 7 9 9 0 4 3 13 9 2 16 1 15 9 4 13 2
8 3 9 7 9 14 13 9 2
5 7 14 15 13 2
7 9 13 1 9 1 9 2
10 13 9 9 2 13 1 12 9 9 2
6 13 15 1 9 9 2
17 3 13 9 1 9 0 1 9 0 2 13 9 7 9 1 9 2
13 1 9 13 15 2 16 4 13 14 1 15 13 2
18 9 9 13 13 0 9 1 9 13 9 9 7 9 7 9 9 0 2
15 9 9 13 9 0 2 7 9 9 4 13 1 9 9 2
5 7 3 13 4 2
13 9 9 13 1 9 0 1 9 0 9 7 9 2
17 13 15 0 9 1 9 2 0 13 9 1 9 9 1 0 9 2
3 14 13 2
4 9 13 0 2
19 9 0 9 2 0 13 0 9 1 9 0 2 13 13 9 9 7 9 2
18 9 13 9 13 0 1 0 9 9 2 0 13 0 9 9 7 9 2
6 13 14 1 0 9 2
12 9 13 13 15 1 0 9 9 1 9 0 2
16 13 0 9 2 13 15 1 9 1 0 9 7 13 1 9 2
5 13 13 0 9 2
7 0 9 1 9 13 9 2
16 3 9 1 9 13 3 1 9 2 13 1 9 7 15 9 2
4 2 14 13 2
4 9 13 9 2
7 13 4 15 13 1 9 2
9 16 13 3 3 2 9 13 9 2
5 2 13 9 14 2
8 13 0 9 2 13 1 9 2
7 9 13 1 9 9 0 2
6 2 13 0 0 9 2
7 1 15 13 14 4 12 2
10 9 2 13 1 9 2 3 13 9 2
3 13 9 2
6 9 3 3 13 9 2
8 2 9 3 3 13 0 9 2
3 2 13 2
10 13 2 16 14 13 0 1 0 9 2
5 13 13 2 2 2
4 9 13 9 2
6 2 13 14 4 13 2
7 1 9 15 1 9 13 2
6 14 15 1 9 13 2
12 7 15 15 14 13 2 7 15 15 14 13 2
8 14 13 4 1 0 9 9 2
6 13 15 9 2 2 2
9 9 13 2 9 13 1 9 0 2
12 1 9 0 2 0 9 0 13 9 1 9 2
8 1 9 13 15 14 9 9 2
17 14 9 0 13 2 16 9 0 0 9 13 0 9 0 1 9 2
14 13 15 2 16 0 1 9 9 9 4 13 1 9 2
8 9 13 14 15 9 1 9 2
18 3 2 1 13 9 0 2 0 9 13 2 16 9 9 13 1 9 2
9 3 15 13 2 16 13 1 9 2
7 14 0 9 13 9 0 2
5 3 9 13 9 2
7 14 0 9 13 1 9 2
8 14 9 1 9 14 13 9 2
10 9 7 13 15 1 0 9 0 9 2
10 9 2 1 0 13 2 13 3 0 2
12 13 1 15 1 9 9 0 9 13 1 9 2
19 13 15 1 9 1 0 9 9 9 2 0 13 9 0 9 13 9 0 2
9 9 9 7 9 13 9 9 0 2
10 14 1 9 14 13 9 1 0 9 2
5 9 9 14 13 2
7 15 15 13 1 0 9 2
14 16 1 9 1 9 14 13 0 2 7 8 9 13 2
8 16 3 2 9 13 3 0 2
12 9 7 9 0 8 2 13 0 13 9 0 2
8 13 15 9 3 0 9 9 2
24 9 2 0 9 0 9 9 2 13 1 9 2 16 0 9 0 9 4 0 9 1 0 9 2
10 1 9 9 7 9 13 14 0 9 2
9 3 13 15 14 0 3 0 9 2
5 9 13 0 9 2
7 3 13 15 1 9 9 2
6 14 1 0 13 9 2
9 3 14 13 4 2 16 13 0 2
6 1 9 9 13 9 2
8 13 9 0 1 9 9 9 2
4 3 15 13 2
20 0 9 13 15 14 1 12 9 2 7 3 14 13 1 15 1 9 2 2 2
14 3 13 4 9 2 13 4 1 9 7 13 4 9 2
11 13 4 1 9 7 3 13 4 1 9 2
10 3 9 13 9 1 9 7 13 9 2
10 13 1 9 2 16 9 13 1 9 2
11 14 13 1 9 7 1 9 9 15 13 2
4 13 1 9 2
7 1 9 14 13 0 9 2
6 13 2 13 1 9 2
8 1 9 13 14 1 0 9 2
5 3 15 15 13 2
12 9 13 1 9 13 1 13 9 1 0 9 2
9 13 0 2 3 3 1 9 13 2
12 13 15 7 13 2 16 13 12 0 9 3 2
11 0 9 0 13 13 9 9 0 1 9 2
7 9 0 13 12 0 9 2
6 2 7 14 13 0 2
6 1 9 13 15 9 2
10 9 13 1 0 9 7 13 1 9 2
14 2 7 3 15 9 13 2 13 4 15 9 3 3 2
12 2 13 9 2 13 9 2 14 15 14 13 2
14 2 13 4 2 14 13 4 2 13 4 7 13 4 2
8 0 9 0 9 3 14 13 2
13 13 9 0 7 9 13 15 3 1 0 9 0 2
21 3 9 9 3 13 2 3 1 0 9 13 0 9 1 9 0 2 13 0 9 2
6 13 14 14 13 9 2
22 16 1 13 12 9 0 9 15 13 2 3 9 13 1 9 13 1 9 3 13 9 2
19 9 0 9 13 15 1 13 0 9 2 13 9 3 3 1 0 9 9 2
13 9 13 2 16 13 1 15 13 9 13 2 2 2
7 0 9 13 7 0 9 2
9 7 9 9 9 13 9 13 9 2
26 9 9 3 13 2 16 15 9 13 13 9 1 9 1 9 9 7 1 9 13 0 9 1 0 9 2
12 1 9 9 9 9 13 15 1 9 0 9 2
5 13 0 9 9 2
12 0 1 9 13 1 0 9 9 13 1 9 2
11 9 9 1 0 1 9 13 9 3 13 2
4 13 9 9 2
9 15 0 13 9 3 0 2 0 2
10 1 9 9 13 9 9 1 0 15 2
8 13 0 0 9 1 12 9 2
10 13 9 1 9 9 1 9 9 0 2
7 9 3 14 9 14 13 2
9 7 15 1 0 9 13 15 9 2
10 14 13 15 14 2 16 13 9 0 2
13 16 0 0 9 13 2 13 1 9 0 14 9 2
12 14 14 0 9 14 13 15 1 9 0 9 2
11 14 13 1 0 9 13 14 1 9 9 2
9 1 12 9 13 9 15 0 9 2
24 16 9 13 3 0 2 13 9 2 16 0 9 13 9 0 1 12 13 1 9 1 0 9 2
13 9 14 14 13 2 7 0 13 15 1 0 9 2
9 2 1 9 9 13 3 0 13 2
9 14 1 9 13 13 1 9 0 2
7 12 9 13 1 9 13 2
15 13 9 13 0 9 9 7 9 2 13 9 1 0 9 2
9 1 9 13 9 9 1 0 9 2
9 9 13 4 1 0 9 0 9 2
9 0 9 13 14 13 7 13 9 2
12 3 1 13 1 0 9 13 14 9 2 2 2
9 2 1 9 13 4 1 0 9 2
22 2 13 4 9 9 2 3 13 3 13 9 12 2 1 0 13 13 9 9 9 9 2
10 2 9 3 14 13 0 9 2 2 2
4 9 13 9 2
24 7 1 9 2 1 9 9 1 9 7 13 9 2 9 9 13 15 1 9 9 13 0 9 2
8 0 9 14 13 4 14 3 2
20 2 1 0 9 9 2 0 13 9 9 2 13 13 9 2 16 4 3 13 2
7 7 3 13 15 2 2 2
7 1 9 13 9 1 9 2
11 13 2 16 3 3 0 13 15 0 9 2
17 2 9 0 9 1 9 15 9 0 4 1 3 3 13 1 9 2
9 3 3 7 13 15 1 0 9 2
14 13 1 9 9 14 13 14 14 9 1 13 9 0 2
7 7 9 13 13 15 9 2
18 0 9 9 0 13 9 1 9 1 9 9 7 13 9 1 13 9 2
10 13 9 13 1 9 13 14 1 13 2
26 7 9 13 1 9 13 0 9 1 9 2 0 9 13 13 0 9 1 3 0 9 1 0 9 9 2
6 13 4 14 0 9 2
9 2 9 13 3 0 9 1 15 2
23 13 14 1 9 2 1 9 13 1 3 2 7 1 9 13 15 7 13 1 9 9 0 2
5 13 15 9 9 2
8 9 1 0 9 0 13 0 2
7 1 0 9 13 15 9 2
5 3 0 4 9 2
9 9 14 13 9 0 13 9 9 2
17 9 9 13 3 0 1 0 13 9 2 0 3 13 15 1 9 2
17 1 9 1 9 9 3 4 13 1 9 7 14 13 1 9 9 2
10 9 9 9 1 9 13 1 15 9 2
10 0 9 14 13 4 3 13 1 9 2
15 9 4 13 1 9 2 0 1 9 13 15 1 0 9 2
9 0 9 0 4 3 0 1 9 2
22 1 0 9 0 9 13 8 2 9 2 8 2 9 2 8 2 9 2 8 2 9 2
10 0 9 2 14 9 2 13 15 13 2
18 13 1 9 0 9 1 0 9 2 13 9 1 9 3 13 1 9 2
11 9 13 9 1 9 13 0 9 1 9 2
10 13 1 9 0 1 9 0 9 9 2
13 13 15 12 2 16 13 14 13 14 9 0 9 2
9 1 0 9 13 15 1 12 9 2
15 3 0 9 3 13 2 16 1 0 9 9 1 9 13 2
8 1 0 9 13 15 3 3 2
15 9 0 13 14 9 9 7 4 13 1 13 1 15 9 2
16 9 13 2 16 0 9 15 13 7 1 9 9 9 13 9 2
16 3 9 0 3 15 13 2 7 14 3 9 13 13 0 9 2
11 0 9 9 13 2 7 0 13 14 13 2
15 3 1 13 1 9 13 4 9 2 7 14 13 14 13 2
8 13 4 15 2 13 1 9 2
6 1 9 13 4 9 2
9 1 9 9 4 13 1 9 9 2
5 9 13 0 9 2
13 0 9 9 1 9 1 0 13 9 13 0 9 2
26 13 9 7 13 2 16 13 0 2 7 13 9 1 9 13 15 2 16 3 14 13 14 1 9 0 2
7 1 9 9 9 13 15 2
3 13 9 2
10 13 15 7 13 3 13 1 0 9 2
3 13 9 2
5 13 13 9 9 2
5 15 9 13 15 2
5 1 0 15 13 2
4 15 15 13 2
4 15 14 13 2
5 1 9 13 9 2
10 13 0 2 0 1 13 9 1 9 2
22 13 1 9 2 13 15 9 0 2 13 4 0 0 9 2 0 13 2 13 1 9 2
8 13 0 2 13 0 0 9 2
6 13 2 3 15 13 2
12 9 13 15 3 1 9 13 15 15 3 0 2
19 9 13 1 0 9 2 7 15 2 13 9 2 13 1 0 1 13 9 2
8 0 0 9 13 0 9 9 2
7 14 9 0 9 0 13 2
8 14 1 9 15 3 9 13 2
13 14 0 4 13 9 0 9 2 16 15 15 13 2
7 1 15 13 9 0 9 2
23 3 3 13 2 7 3 13 15 0 9 13 1 9 2 0 9 0 9 13 1 9 9 2
7 9 13 15 3 0 9 2
9 9 9 13 0 1 9 9 9 2
8 0 13 2 1 9 9 13 2
16 2 9 14 13 0 2 16 14 13 2 16 13 15 0 9 2
5 13 4 0 9 2
7 1 9 13 15 3 3 2
8 13 15 9 1 9 13 9 2
13 9 0 9 13 2 16 14 9 3 14 13 3 2
10 2 13 1 9 9 2 15 14 13 2
7 9 9 13 15 1 9 2
20 9 0 13 1 9 8 2 12 9 2 16 9 1 15 13 13 1 9 13 2
6 3 15 13 2 2 2
10 14 13 15 15 2 3 2 2 2 2
5 16 13 15 13 2
4 2 13 15 2
12 13 3 13 2 16 14 13 2 1 9 13 2
4 15 9 13 2
10 2 9 2 13 4 15 1 9 2 2
6 2 14 13 15 13 2
5 3 2 13 9 2
5 7 3 15 13 2
9 3 13 1 9 1 9 9 9 2
8 13 4 9 1 9 9 9 2
9 9 1 12 9 13 15 0 9 2
7 13 15 1 9 0 9 2
18 3 13 4 13 0 2 0 9 1 9 2 1 0 13 13 3 9 2
7 13 2 16 9 13 0 2
13 13 14 2 16 9 0 9 13 3 13 9 0 2
11 1 0 9 9 13 13 3 13 0 9 2
6 13 13 9 1 9 2
22 16 13 3 0 9 9 2 9 2 14 13 1 13 15 1 0 9 2 9 7 9 2
9 13 9 1 13 2 13 0 9 2
10 13 15 13 2 16 3 3 13 15 2
6 13 7 13 0 9 2
15 1 0 9 13 1 9 9 2 13 4 9 8 2 9 2
6 14 13 15 2 2 2
13 1 9 2 16 13 15 13 1 9 2 13 15 2
10 14 13 15 9 7 13 3 13 9 2
11 2 14 13 4 7 13 4 9 2 2 2
3 2 13 2
4 9 13 3 2
3 9 13 2
15 7 15 13 0 2 0 2 0 2 0 7 0 2 2 2
16 9 13 15 0 0 9 1 9 9 2 13 2 16 15 13 2
10 2 9 1 0 9 13 1 0 9 2
3 9 13 2
4 2 13 0 2
19 13 14 7 1 9 1 9 2 9 15 13 1 9 2 3 1 0 9 2
8 9 3 14 13 0 13 9 2
10 12 13 1 9 2 9 2 0 9 2
9 9 9 7 9 14 13 0 9 2
30 15 9 2 13 1 9 0 2 13 9 9 0 2 7 3 13 3 3 9 1 0 9 2 16 1 0 9 13 9 2
11 4 13 9 2 9 1 0 9 7 9 2
5 14 13 9 0 2
5 14 13 9 0 2
5 7 13 9 9 2
7 9 9 13 15 3 0 2
10 9 14 13 15 1 9 9 9 0 2
6 13 15 14 9 9 2
27 16 14 1 12 9 1 9 13 0 0 9 9 0 9 0 2 7 3 13 15 9 13 2 7 7 0 2
11 9 9 9 9 3 13 1 9 1 9 2
8 9 13 2 13 14 0 9 2
23 9 0 9 2 4 13 0 9 2 16 9 13 2 16 9 9 13 1 9 0 9 0 2
11 13 15 2 16 9 1 9 13 0 9 2
12 14 14 3 13 7 14 13 9 13 0 9 2
12 2 3 14 13 4 0 9 2 13 4 2 2
5 2 13 4 2 2
5 13 15 15 3 2
7 13 4 3 9 1 9 2
7 13 15 3 0 1 9 2
4 13 0 9 2
3 13 15 2
4 9 13 9 2
9 9 13 1 15 13 1 9 0 2
5 7 3 3 13 2
8 7 9 14 13 2 3 13 2
13 9 3 13 9 13 1 0 2 0 7 0 9 2
9 3 1 9 1 9 13 0 9 2
3 14 13 2
7 13 1 9 0 1 9 2
11 9 2 0 13 2 13 14 9 1 9 2
6 7 14 13 15 9 2
7 13 2 16 9 14 13 2
20 9 13 1 9 7 4 13 3 13 1 0 9 2 9 1 9 0 15 13 2
14 0 9 1 9 1 0 9 13 2 3 13 15 9 2
5 13 1 15 13 2
14 3 1 9 0 13 1 9 0 0 9 1 9 9 2
8 16 14 13 13 3 1 9 2
11 13 15 9 2 13 1 9 2 13 9 2
5 3 13 1 9 2
5 2 9 13 9 2
6 2 13 4 13 9 2
7 13 0 9 1 0 9 2
7 2 9 13 15 1 9 2
17 3 3 13 9 0 2 16 13 9 9 0 2 0 13 13 0 2
15 1 9 0 9 13 1 3 12 9 1 9 9 9 0 2
12 13 15 9 7 9 1 9 13 9 9 0 2
8 13 9 9 1 9 9 0 2
10 9 1 9 13 9 13 1 9 0 2
12 3 9 0 13 1 9 2 9 7 9 9 2
23 0 9 0 9 13 15 1 0 9 0 1 0 9 0 9 1 9 9 0 7 9 0 2
11 9 9 13 1 9 9 9 7 9 9 2
8 9 4 13 1 0 0 8 2
12 2 9 1 0 8 2 14 4 14 15 13 2
13 3 3 13 0 2 0 1 9 7 9 9 9 2
16 0 9 2 1 0 9 9 1 0 9 2 13 9 9 9 2
15 14 0 13 9 13 1 9 0 9 1 13 0 9 9 2
7 3 13 9 9 1 9 2
5 13 9 0 9 2
10 13 15 3 3 2 3 9 13 0 2
6 13 9 1 0 9 2
8 13 3 0 0 9 7 9 2
9 2 3 0 13 9 0 2 0 2
6 13 13 9 1 9 2
10 2 13 15 13 2 3 13 3 13 2
10 2 14 13 0 9 7 13 1 15 2
5 9 13 3 9 2
9 9 9 0 13 1 9 0 9 2
7 0 9 13 9 13 9 2
10 14 14 1 0 9 13 15 9 13 2
5 13 9 1 9 2
6 13 0 13 2 9 2
14 1 9 13 7 13 0 0 9 13 9 1 9 9 2
7 13 9 9 9 2 13 2
7 4 9 9 0 2 2 2
7 12 13 9 13 1 9 2
8 13 3 7 13 1 9 9 2
12 9 13 9 9 2 1 9 13 0 0 9 2
16 13 15 2 13 9 0 9 2 0 13 15 1 9 2 2 2
6 9 13 13 1 9 2
8 9 13 15 15 1 0 9 2
28 16 1 12 9 13 4 1 9 0 1 0 9 2 14 13 15 2 16 3 13 15 1 9 12 9 1 15 2
7 16 13 9 2 13 9 2
13 1 0 14 9 9 7 9 13 15 1 9 0 2
7 1 0 9 9 14 13 2
8 3 13 9 13 15 0 9 2
9 3 0 9 13 0 9 0 9 2
7 13 14 1 15 0 9 2
9 13 15 9 13 15 1 0 9 2
14 2 13 3 0 1 9 2 7 3 15 14 13 4 2
5 9 14 13 9 2
9 9 14 13 0 13 1 15 9 2
7 9 14 13 9 7 9 2
10 9 14 13 9 7 9 1 15 3 2
5 9 14 13 9 2
5 9 14 13 9 2
5 9 14 13 9 2
9 9 14 13 0 9 2 14 9 2
8 9 14 13 9 13 7 9 2
11 13 2 16 13 1 0 9 9 7 9 2
13 1 0 9 9 9 13 2 13 0 9 1 9 2
3 13 15 2
7 13 14 15 13 1 9 2
16 3 3 13 9 2 7 13 2 16 13 9 3 0 7 0 2
22 7 9 2 9 7 9 9 13 15 9 2 9 2 9 7 9 1 9 0 7 0 2
9 1 0 9 15 9 13 0 9 2
11 9 9 13 1 9 9 2 7 14 9 2
8 9 13 0 9 7 0 9 2
12 9 13 2 16 13 0 2 7 13 13 9 2
5 3 13 9 9 2
3 13 9 2
12 12 9 1 13 15 1 0 9 0 1 9 2
13 13 3 0 2 1 0 2 7 13 1 15 9 2
4 7 13 15 2
5 7 9 13 0 2
11 1 13 9 0 7 9 9 9 14 13 2
12 9 13 0 7 0 2 7 13 15 13 9 2
6 9 14 13 15 13 2
13 15 1 9 13 9 7 14 13 15 3 1 15 2
6 13 1 9 0 9 2
12 9 9 7 9 13 1 9 2 15 9 13 2
9 13 4 2 1 9 15 13 4 2
7 9 13 12 9 1 9 2
6 9 13 15 3 13 2
11 2 13 1 9 0 7 14 4 13 9 2
20 1 9 13 2 16 3 14 13 13 9 2 7 14 13 1 9 0 9 9 2
9 13 1 15 12 9 7 0 9 2
10 2 13 9 13 2 16 9 14 13 2
9 2 15 1 0 9 13 0 9 2
6 2 7 9 15 13 2
6 2 7 15 15 13 2
12 7 15 13 9 0 9 2 7 13 14 15 2
7 2 13 7 13 0 9 2
6 2 9 13 14 3 2
14 2 15 12 13 14 3 2 16 1 9 13 15 9 2
13 2 14 15 1 9 13 2 7 15 14 14 13 2
4 9 13 9 2
12 0 9 13 1 9 9 2 3 13 15 13 2
2 13 2
12 1 15 13 7 13 9 9 9 13 15 9 2
11 15 9 13 15 1 9 2 13 9 0 2
5 9 13 1 9 2
8 13 9 7 9 13 1 9 2
6 9 13 15 1 15 2
4 13 2 2 2
6 1 9 14 14 13 2
6 2 9 15 15 13 2
8 1 9 9 13 4 0 9 2
8 3 15 14 13 1 0 9 2
11 14 2 13 2 13 2 3 13 2 2 2
6 2 3 14 13 4 2
10 13 4 15 1 9 2 7 13 4 2
4 13 1 9 2
12 9 13 1 9 1 9 12 9 1 9 13 2
9 13 4 2 16 13 2 9 13 2
11 1 9 13 4 15 1 9 2 13 9 2
6 14 15 9 14 13 2
8 9 1 0 9 13 9 9 2
8 14 14 9 1 9 15 13 2
12 14 13 15 9 2 3 15 9 13 1 9 2
18 3 14 14 13 2 14 2 13 9 2 7 0 9 4 13 0 9 2
3 14 13 2
17 9 0 13 1 0 9 1 9 9 1 13 9 7 9 9 0 2
4 9 3 13 2
6 9 13 1 0 9 2
6 3 9 13 1 9 2
8 14 15 14 13 1 0 9 2
4 0 9 13 2
7 14 0 13 13 0 9 2
16 14 1 9 13 4 15 2 16 3 13 4 1 9 0 9 2
9 13 4 3 2 16 9 4 13 2
4 13 4 15 2
7 13 2 16 13 9 9 2
5 13 4 0 9 2
32 9 13 1 9 9 7 14 13 0 2 13 9 9 9 2 16 0 9 0 9 9 13 13 2 7 9 13 0 1 9 9 2
8 1 0 9 13 15 9 9 2
4 9 9 13 2
10 3 13 2 13 15 9 7 13 9 2
10 16 13 15 9 2 9 13 9 9 2
23 9 15 13 9 7 15 9 2 7 0 9 1 9 13 0 9 14 9 1 9 1 9 2
8 14 13 4 15 1 9 13 2
9 14 0 0 9 14 13 15 9 2
10 1 9 14 14 13 4 13 15 9 2
22 3 13 13 1 9 7 9 9 2 7 0 13 9 13 13 9 2 16 13 15 9 2
16 15 14 9 13 4 2 16 13 4 15 1 9 1 9 0 2
16 13 9 1 9 1 9 2 13 2 16 13 13 1 0 9 2
9 12 0 9 9 9 13 0 9 2
9 3 3 0 13 15 9 13 9 2
6 9 13 1 9 9 2
9 9 0 4 13 1 9 1 9 2
19 1 9 0 9 1 9 9 2 0 9 1 9 13 15 1 15 0 9 2
18 13 1 0 9 2 13 7 13 9 1 9 1 0 9 9 9 9 2
6 7 3 13 1 9 2
9 1 9 1 9 0 13 12 9 2
11 9 1 12 9 13 0 9 1 9 9 2
12 1 0 9 9 9 13 9 9 2 9 9 2
10 1 0 9 9 13 1 9 9 13 2
7 1 9 9 13 1 0 2
20 3 13 9 0 1 9 2 16 13 2 16 1 9 13 14 12 9 1 13 2
15 1 9 13 4 15 13 2 16 13 0 9 1 9 9 2
17 13 15 3 0 2 13 9 0 9 1 0 9 9 1 9 0 2
12 0 0 9 13 1 9 0 9 1 0 8 2
13 9 0 13 0 9 2 0 13 15 9 7 9 2
9 7 9 0 13 14 0 1 9 2
14 9 0 1 9 13 15 14 1 9 1 0 9 9 2
7 9 0 9 13 2 2 2
13 1 9 2 9 13 2 7 9 9 4 13 9 2
19 0 9 4 9 0 9 0 1 9 0 2 7 14 9 0 7 9 0 2
8 13 14 9 9 0 7 0 2
9 13 14 0 9 9 1 9 0 2
20 3 13 9 0 9 0 7 9 9 0 9 1 0 9 9 7 9 7 9 2
8 9 13 15 0 9 1 9 2
8 1 9 13 0 9 7 9 2
8 9 0 13 13 15 0 9 2
20 1 0 0 9 2 0 13 9 9 9 2 9 13 14 9 1 9 9 0 2
3 13 15 2
12 1 9 9 13 9 9 0 2 0 7 0 2
15 14 0 9 1 9 13 7 9 9 2 7 9 9 0 2
10 0 13 1 9 0 9 0 13 0 2
11 13 1 0 9 7 13 1 9 0 9 2
12 3 13 13 0 9 2 14 13 2 3 13 2
9 1 9 13 1 9 1 0 9 2
10 13 4 0 9 2 16 13 9 9 2
4 9 13 15 2
8 2 9 15 15 1 15 13 2
6 9 13 15 0 9 2
17 14 0 13 4 3 1 9 2 3 13 4 9 13 1 0 9 2
5 13 4 1 9 2
8 13 14 13 1 9 9 0 2
25 13 4 2 16 0 9 1 9 14 13 2 7 1 0 9 14 13 4 15 1 9 9 0 9 2
7 3 9 4 13 9 0 2
11 9 9 8 2 13 15 14 9 9 0 2
13 9 0 9 13 15 1 9 1 0 12 9 0 2
25 1 9 0 1 9 9 0 2 0 13 1 9 0 2 13 0 9 9 0 1 0 9 9 0 2
16 3 0 9 0 13 9 0 9 1 9 1 9 0 1 9 2
6 3 14 13 9 0 2
15 3 3 2 0 0 9 9 13 9 0 2 13 9 9 2
7 13 9 14 9 9 13 2
14 0 9 13 1 9 2 7 15 1 15 9 3 13 2
11 0 9 13 2 0 9 4 13 9 9 2
6 3 14 13 15 12 2
9 2 14 1 9 13 13 0 9 2
6 2 14 13 0 9 2
6 9 13 1 9 9 2
13 2 14 13 1 9 9 7 3 13 1 0 9 2
8 9 0 9 3 15 15 13 2
7 9 13 1 9 9 13 2
5 13 0 9 9 2
23 13 9 2 9 0 2 7 1 9 9 3 13 9 1 13 9 2 0 3 12 3 13 2
7 0 9 13 1 0 9 2
7 9 9 13 15 3 3 2
23 0 9 9 13 1 9 7 13 15 1 13 9 2 0 9 13 1 9 0 1 0 9 2
20 9 0 2 13 1 0 8 2 7 13 1 9 2 14 13 14 0 9 0 2
8 16 3 13 0 9 13 3 2
8 2 14 13 9 1 13 9 2
7 2 14 13 9 9 9 2
6 15 15 14 13 0 2
13 13 1 0 9 2 4 14 1 0 9 3 13 2
8 1 9 15 3 14 13 4 2
14 3 13 1 15 0 9 7 3 15 1 15 13 4 2
13 1 0 9 13 4 15 2 13 1 0 0 9 2
16 3 1 9 13 1 0 9 0 13 9 9 14 13 1 0 2
16 1 9 3 13 9 9 2 1 9 9 9 13 15 3 3 2
13 13 2 16 13 13 1 9 7 9 1 0 9 2
8 3 13 4 0 15 9 0 2
15 1 9 13 4 9 1 9 2 0 9 13 9 0 9 2
18 3 13 2 16 13 13 2 16 13 0 9 2 7 9 13 3 0 2
9 13 4 0 9 1 13 9 9 2
10 13 1 9 1 12 9 13 0 9 2
8 9 9 13 15 1 15 13 2
8 9 14 13 7 13 9 13 2
7 3 3 4 13 9 0 2
14 12 9 1 1 9 1 0 9 0 9 13 13 9 2
12 2 13 9 2 13 9 2 7 9 13 0 2
7 1 9 0 13 13 9 2
9 13 14 3 9 2 9 9 9 2
17 16 13 9 0 1 9 2 0 9 13 1 15 0 9 9 9 2
16 15 0 9 13 1 12 9 3 1 15 0 1 0 14 9 2
6 14 13 9 1 15 2
6 14 13 15 1 9 2
9 9 13 1 0 9 0 9 9 2
13 9 0 9 13 1 9 9 0 1 0 9 9 2
24 13 14 9 1 9 7 9 9 0 13 2 16 12 9 2 9 7 9 2 13 4 9 9 2
12 0 9 13 15 14 3 13 3 0 9 9 2
9 14 13 4 9 8 2 9 9 2
19 9 13 0 2 9 0 14 13 15 1 0 9 7 13 15 1 9 13 2
9 9 14 13 7 9 1 0 9 2
12 13 14 12 9 2 1 0 9 3 14 13 2
19 1 0 2 0 2 0 9 13 15 1 9 9 7 9 2 9 7 9 2
8 9 1 9 9 13 3 12 2
14 0 0 9 0 13 12 9 2 1 0 3 13 12 2
8 9 13 2 13 15 2 13 2
14 9 13 15 3 2 1 0 9 1 9 13 0 9 2
23 3 3 9 13 9 0 9 2 9 2 16 14 13 15 15 13 0 9 1 3 13 9 2
10 13 1 9 2 13 13 1 9 0 2
7 0 9 13 0 9 9 2
9 9 1 9 13 15 1 13 9 2
10 9 13 0 1 0 9 7 0 9 2
20 9 13 15 0 7 14 9 1 15 13 2 3 13 1 0 9 0 0 9 2
16 9 0 9 13 16 9 0 9 2 14 13 14 15 0 9 2
8 15 9 13 1 0 9 0 2
13 1 0 9 9 9 3 14 4 13 1 9 0 2
11 0 9 13 9 12 9 1 1 9 0 2
16 12 8 2 9 9 13 2 16 9 9 1 9 13 3 0 2
11 13 9 13 15 3 9 2 9 7 9 2
17 1 0 9 1 9 0 9 13 0 9 2 13 9 1 13 9 2
8 9 1 13 9 13 0 9 2
12 0 9 0 4 0 1 0 9 7 9 0 2
13 9 1 9 1 0 13 15 1 9 1 0 9 2
12 1 9 9 9 1 9 13 15 13 12 9 2
5 15 15 13 2 2
5 2 15 14 13 2
4 9 14 13 2
3 2 13 2
10 2 13 4 15 2 9 9 2 2 2
5 9 1 15 13 2
6 9 7 9 9 13 2
11 2 7 9 14 3 13 9 2 2 2 2
7 14 9 3 13 0 9 2
4 13 3 3 2
9 9 13 9 13 9 9 9 0 2
12 1 9 9 9 13 13 13 9 13 1 9 2
18 1 0 9 9 13 1 9 9 13 15 1 9 7 15 9 9 0 2
10 9 9 14 13 2 9 13 1 15 2
7 13 3 2 1 0 9 2
5 9 9 14 13 2
8 9 1 9 14 13 0 9 2
5 13 9 1 13 2
4 13 0 9 2
9 0 9 14 13 15 1 9 13 2
16 1 9 13 4 9 7 13 15 1 0 9 2 1 0 9 2
5 13 4 1 0 2
11 16 13 4 12 9 2 13 15 1 9 2
15 14 13 4 13 1 0 7 0 2 7 14 13 0 9 2
5 13 9 1 9 2
9 3 13 13 1 0 9 2 13 2
6 13 13 1 0 9 2
7 13 14 3 9 2 13 2
12 7 3 13 9 9 2 14 15 3 14 13 2
5 16 15 9 13 2
6 13 4 13 1 9 2
5 0 9 13 12 2
2 13 2
6 9 13 1 0 9 2
4 9 14 13 2
6 13 15 15 1 9 2
3 13 9 2
8 15 9 1 9 9 13 0 2
6 9 0 13 1 9 2
16 9 13 15 9 0 7 1 9 9 14 13 0 9 13 9 2
6 9 13 13 0 9 2
11 13 13 1 9 9 1 9 0 7 0 2
9 9 13 7 13 15 1 9 9 2
6 2 3 9 3 13 2
17 9 7 0 9 2 13 3 2 13 9 1 9 7 13 1 9 2
6 2 9 15 15 13 2
4 2 3 13 2
11 2 13 14 4 13 0 2 16 15 13 2
5 9 15 3 13 2
11 7 9 9 7 9 13 0 1 0 9 2
15 0 13 1 15 9 2 1 3 13 14 15 9 3 3 2
5 0 9 13 9 2
7 1 0 9 13 15 9 2
6 1 9 13 0 9 2
4 3 13 9 2
6 13 4 9 1 9 2
6 1 9 7 9 13 2
6 13 1 15 0 9 2
6 9 14 13 1 9 2
10 9 9 1 9 13 1 9 1 9 2
17 9 0 13 14 1 9 9 2 16 0 13 14 9 9 1 9 2
4 9 13 9 2
14 9 2 1 9 9 9 2 13 9 7 9 0 9 2
3 13 9 2
15 9 13 15 1 9 9 2 13 9 7 13 13 1 9 2
5 13 15 7 13 2
10 1 0 9 13 4 14 9 1 15 2
18 9 13 14 1 15 1 0 0 9 2 1 0 13 4 15 3 3 2
6 2 13 0 0 9 2
9 3 0 9 9 13 15 0 9 2
15 9 9 2 9 9 2 13 12 9 1 0 9 1 9 2
26 13 15 15 0 9 1 0 9 2 13 1 0 1 0 9 2 7 14 0 9 2 0 9 7 9 2
6 3 1 9 14 13 2
10 13 15 2 16 1 9 13 12 9 2
9 3 14 13 1 13 9 7 9 2
6 7 13 15 9 13 2
13 13 2 16 1 9 9 0 14 13 15 9 9 2
19 1 9 13 12 9 9 9 2 0 13 1 12 9 1 0 9 9 9 2
10 9 4 13 1 9 0 9 1 9 2
12 9 0 1 9 13 3 0 9 13 9 0 2
17 1 0 9 13 4 0 9 2 13 1 0 9 1 9 9 9 2
12 1 9 0 13 1 9 9 0 0 9 9 2
12 1 9 13 1 9 1 9 1 9 0 9 2
7 9 9 1 9 14 13 2
15 9 4 13 13 1 13 3 1 9 8 2 9 9 0 2
11 0 13 9 9 9 2 0 13 13 9 2
8 13 1 0 9 9 9 0 2
7 9 3 13 1 9 9 2
6 1 9 13 15 9 2
13 13 9 1 9 9 13 0 9 9 2 9 9 2
8 3 9 3 13 1 9 9 2
11 9 13 9 0 2 0 3 13 0 9 2
5 3 9 13 9 2
9 1 0 9 9 9 13 9 0 2
18 0 9 2 14 13 0 9 9 1 9 0 9 2 3 13 1 9 2
23 14 1 9 13 15 1 9 0 7 14 3 13 9 2 3 13 9 7 0 9 1 9 2
4 13 4 9 2
10 14 2 14 0 9 15 13 13 9 2
7 13 1 9 1 9 0 2
13 9 13 12 9 1 9 9 9 1 9 1 9 2
5 3 13 15 9 2
5 1 9 13 9 2
22 1 9 13 0 9 2 16 9 0 9 13 9 1 12 9 13 1 9 1 0 9 2
8 0 9 13 9 0 0 9 2
5 9 13 1 15 2
6 2 13 9 2 2 2
19 1 0 9 9 9 13 15 13 1 0 9 2 1 0 9 13 0 9 2
3 13 9 2
5 2 9 15 13 2
11 2 13 2 13 15 2 9 13 1 13 2
10 14 13 2 3 3 9 13 1 9 2
7 2 13 9 1 0 9 2
20 1 15 9 13 9 2 13 13 2 3 9 13 9 14 13 15 1 13 9 2
4 9 13 9 2
6 2 9 3 15 13 2
20 9 13 9 1 9 7 13 15 1 9 2 9 9 13 2 16 15 3 13 2
4 9 13 9 2
6 9 13 1 9 9 2
16 9 13 9 2 16 13 13 1 9 2 7 14 3 13 9 2
5 14 13 14 0 2
15 0 9 9 13 9 1 0 0 9 9 0 9 1 9 2
19 12 0 9 3 13 14 15 1 9 9 9 2 16 9 13 9 0 9 2
15 13 9 2 7 9 13 15 1 0 9 13 15 1 9 2
5 9 0 13 9 2
8 13 15 9 0 9 7 9 2
12 9 0 9 13 3 1 9 0 13 0 9 2
18 9 13 2 16 13 0 2 16 14 13 2 16 9 13 13 0 9 2
10 12 9 1 1 9 13 13 9 9 2
9 1 0 9 9 0 13 0 9 2
13 13 9 9 0 7 9 0 9 13 3 3 0 2
12 0 9 13 1 9 9 1 9 0 9 0 2
15 0 9 13 15 2 16 13 15 0 9 1 9 0 9 2
18 1 13 2 0 9 9 9 1 9 9 13 15 15 9 7 9 0 2
12 0 9 13 9 0 9 2 9 7 15 9 2
9 9 0 9 13 9 13 12 9 2
7 9 13 14 9 9 0 2
13 9 2 9 9 7 13 9 13 9 1 9 9 2
5 3 13 4 13 2
13 9 13 13 15 1 9 3 1 9 9 9 0 2
5 13 9 9 9 2
9 9 13 13 9 2 9 2 9 2
8 13 2 16 9 13 15 3 2
5 9 13 9 9 2
20 1 9 13 9 1 9 9 2 13 1 9 2 13 9 2 13 8 1 9 2
11 9 13 9 2 16 15 13 1 0 9 2
6 13 9 9 0 9 2
18 9 13 13 0 9 1 0 9 0 1 12 9 7 9 0 7 0 2
10 1 9 9 9 13 4 13 9 0 2
4 9 13 15 2
4 14 4 13 2
5 15 9 14 13 2
7 9 13 15 3 1 9 2
5 13 9 1 9 2
4 9 13 9 2
17 2 13 1 9 1 12 9 7 13 2 16 13 3 1 9 9 2
4 2 13 0 2
8 14 13 14 4 13 0 9 2
9 9 15 13 9 7 3 13 4 2
11 14 3 4 14 4 15 9 13 1 9 2
11 9 14 1 9 14 13 9 0 1 9 2
4 13 15 12 2
10 14 14 13 2 14 3 3 13 13 2
16 0 13 15 0 9 13 3 1 0 9 0 14 9 0 9 2
11 3 13 15 15 9 0 7 9 9 0 2
11 14 13 7 9 1 9 7 9 9 0 2
13 13 4 1 9 0 12 9 2 13 9 1 12 2
5 3 13 15 13 2
6 7 13 9 1 9 2
4 13 1 9 2
7 1 9 9 13 9 9 2
3 13 9 2
5 13 15 9 9 2
3 14 13 2
6 14 13 13 9 13 2
9 1 15 14 13 14 0 9 0 2
20 13 9 2 16 3 9 14 4 13 9 1 9 2 16 9 13 0 3 9 2
13 0 9 14 13 3 0 0 9 1 9 0 9 2
8 7 1 0 9 13 3 3 2
22 15 9 13 4 2 16 13 4 1 9 1 9 1 0 9 7 13 4 9 1 9 2
13 9 15 13 1 9 9 9 2 9 9 2 2 2
18 9 9 2 9 2 9 0 13 13 1 9 9 7 9 9 9 9 2
10 3 0 9 1 9 13 9 9 9 2
14 9 9 2 9 7 9 13 15 1 0 9 1 9 2
8 2 1 0 15 13 3 3 2
8 2 4 3 1 0 0 9 2
10 2 13 3 2 4 1 3 2 2 2
26 13 4 14 1 9 9 0 12 9 2 3 4 13 12 9 2 7 4 3 3 1 0 2 7 0 2
26 2 14 3 15 3 1 0 9 9 13 2 16 0 13 9 1 15 2 7 0 3 13 7 9 13 2
3 2 13 2
7 1 9 13 13 1 9 2
7 14 9 1 0 3 13 2
7 2 14 13 4 0 9 2
11 0 9 9 0 13 0 9 13 1 9 2
13 15 9 13 2 16 13 1 9 9 13 1 9 2
11 0 9 9 13 1 9 1 0 9 0 2
15 7 13 1 15 0 0 2 0 1 0 9 2 9 0 2
6 13 1 9 9 9 2
9 13 2 16 9 0 1 9 13 2
12 15 1 9 13 0 9 1 0 9 9 0 2
17 1 13 0 9 1 9 0 9 9 0 2 0 1 9 9 13 2
15 13 3 9 7 13 0 9 2 0 14 9 9 15 13 2
26 0 9 0 2 3 13 9 9 1 0 9 1 9 0 9 2 13 15 1 9 9 1 0 9 0 2
16 2 13 0 9 2 13 15 2 14 13 2 16 9 14 13 2
11 14 9 9 14 13 2 13 1 0 9 2
9 2 0 9 9 13 1 13 9 2
10 13 15 0 9 0 9 9 1 9 2
8 3 13 9 2 0 13 9 2
5 13 0 9 9 2
5 13 9 7 9 2
13 2 14 1 0 9 13 4 2 16 9 4 13 2
5 7 9 13 0 2
4 16 13 9 2
9 0 9 1 9 1 9 13 9 2
5 3 15 14 13 2
12 3 13 9 7 9 13 15 1 9 1 9 2
20 1 0 9 14 3 13 2 16 0 9 14 13 15 1 15 2 14 13 9 2
7 1 9 13 9 13 9 2
16 13 2 16 14 13 9 1 0 9 9 9 0 1 0 9 2
13 1 9 2 1 9 14 13 13 0 9 9 9 2
22 9 7 9 13 9 1 9 2 0 4 13 13 0 9 9 2 9 2 9 7 9 2
26 9 12 13 14 9 1 13 15 1 0 9 0 2 0 9 2 0 13 2 16 0 9 4 9 9 2
13 1 8 2 9 13 3 1 9 9 1 0 9 2
7 9 14 13 1 15 9 2
13 13 15 2 16 1 9 13 9 0 0 9 9 2
6 13 15 9 14 3 2
8 1 0 9 9 13 0 9 2
6 1 9 13 0 9 2
9 2 13 9 2 3 4 13 2 2
3 13 9 2
6 13 4 15 1 9 2
6 7 9 14 15 13 2
12 3 13 9 7 13 1 0 9 2 16 13 2
8 0 9 14 13 1 0 9 2
10 2 9 1 15 13 13 1 15 9 2
6 2 13 15 1 9 2
12 2 3 14 13 9 9 1 9 1 0 9 2
4 3 9 13 2
10 2 7 13 2 16 9 13 1 9 2
16 2 13 4 1 9 9 2 1 0 0 9 13 15 0 9 2
4 13 15 9 2
9 1 9 3 9 14 13 0 9 2
7 13 9 13 9 0 9 2
12 14 13 2 16 1 0 9 13 15 0 9 2
6 9 13 15 1 9 2
8 0 13 15 3 0 7 0 2
14 0 9 13 7 9 1 9 1 9 0 2 0 3 2
8 13 4 0 9 1 13 9 2
8 13 3 2 7 4 14 9 2
5 13 14 14 13 2
8 9 9 13 14 1 0 9 2
3 3 13 2
20 13 13 9 1 9 2 16 0 9 0 13 15 1 9 9 0 7 9 9 2
7 9 13 9 2 0 13 2
7 1 9 9 13 9 9 2
11 3 13 9 9 2 16 0 9 13 9 2
11 13 2 16 9 9 3 13 9 1 9 2
8 9 9 9 12 13 12 9 2
19 16 13 15 13 9 13 2 13 14 15 9 9 13 0 9 0 9 9 2
37 9 8 2 13 2 16 15 9 14 13 0 9 2 7 9 13 1 9 2 13 9 7 3 13 0 0 9 2 13 15 1 9 1 9 1 9 2
11 14 9 3 15 13 2 16 9 13 9 2
8 9 14 9 13 1 9 0 2
12 0 9 9 7 9 9 13 0 9 1 9 2
9 1 15 14 13 9 1 0 9 2
5 9 13 9 0 2
16 9 2 0 14 4 13 1 9 2 1 9 4 1 15 13 2
12 0 9 1 13 9 13 9 0 13 1 9 2
6 1 9 13 12 9 2
5 16 14 13 9 2
13 7 3 13 9 2 0 13 1 9 9 1 9 2
4 13 9 0 2
14 9 2 0 13 0 9 1 9 2 14 13 0 9 2
17 1 9 0 9 3 13 1 9 0 12 0 9 2 1 9 9 2
4 14 13 15 2
5 7 13 15 13 2
9 1 13 13 15 0 9 9 9 2
10 1 0 9 0 3 9 15 13 4 2
4 13 4 9 2
19 13 4 9 3 1 13 15 1 0 9 2 0 2 0 3 14 13 9 2
7 9 1 9 9 14 13 2
13 16 9 0 13 15 1 9 2 3 13 14 9 2
21 14 13 4 7 9 9 2 9 9 7 15 9 2 9 1 9 9 7 9 9 2
8 1 0 9 9 14 15 13 2
16 13 9 13 12 9 9 2 0 13 0 9 13 1 9 9 2
19 14 2 0 9 1 9 1 9 13 3 7 14 13 13 2 9 13 9 2
13 0 14 14 13 15 0 9 2 16 9 13 0 2
3 13 9 2
6 2 13 15 13 9 2
5 9 0 13 9 2
15 13 14 9 2 0 13 13 9 1 9 1 13 1 9 2
13 14 13 9 1 9 2 14 13 15 0 13 13 2
19 14 1 0 9 0 9 13 1 9 2 7 1 9 9 1 9 4 0 2
7 13 3 9 9 2 2 2
7 0 9 13 15 9 9 2
14 9 0 13 2 9 15 13 9 9 1 9 0 9 2
14 3 9 0 4 13 2 16 9 14 13 15 1 0 2
12 1 0 9 9 13 9 2 1 0 15 13 2
12 0 9 13 13 0 9 7 13 15 1 9 2
6 3 0 9 9 13 2
15 9 9 14 13 2 7 1 0 9 13 15 13 1 9 2
15 13 1 9 2 1 0 9 9 9 7 9 13 0 9 2
15 1 9 1 9 0 13 1 9 0 9 13 1 9 9 2
15 13 0 9 7 13 2 16 9 13 15 1 3 0 9 2
9 7 3 14 13 2 9 13 9 2
5 2 13 0 9 2
8 9 0 1 15 13 0 9 2
12 9 9 13 1 15 9 13 9 0 9 9 2
7 2 3 9 13 0 9 2
6 9 9 13 2 2 2
22 3 9 9 14 13 2 16 0 9 13 3 7 13 9 2 16 13 15 9 2 2 2
7 1 9 9 14 13 9 2
31 9 0 1 9 2 0 13 9 1 9 9 9 1 0 8 2 2 13 2 16 13 9 1 9 1 12 9 1 12 9 2
10 0 9 1 9 9 13 8 2 9 2
7 9 9 3 1 15 13 2
10 13 0 9 0 13 13 9 1 9 2
10 12 9 1 9 13 9 7 13 9 2
25 0 9 9 1 13 0 9 13 14 14 1 15 0 9 2 13 9 9 9 0 9 0 0 9 2
24 1 0 9 2 1 0 9 0 9 9 0 13 3 0 7 0 2 13 14 9 0 9 9 2
11 1 0 9 1 9 3 13 12 8 9 2
17 3 1 0 9 9 2 9 7 9 13 15 1 9 1 13 9 2
6 9 13 9 0 9 2
14 9 13 1 9 2 0 13 15 1 0 9 1 9 2
6 13 1 15 12 9 2
6 2 13 3 1 9 2
5 3 13 15 9 2
5 4 15 14 12 2
8 13 15 9 13 3 9 9 2
5 3 13 9 0 2
8 3 1 9 13 15 15 9 2
15 2 1 9 2 1 14 9 9 2 14 13 4 1 9 2
14 7 9 14 13 14 1 9 3 2 4 13 15 13 2
13 2 13 9 0 7 13 9 9 2 16 9 13 2
6 2 13 4 15 3 2
8 2 13 9 13 1 9 9 2
10 1 9 9 1 9 13 14 1 9 2
22 9 0 7 9 13 2 16 3 13 15 9 12 9 2 1 9 9 2 9 7 9 2
12 9 13 1 9 2 3 1 9 13 15 9 2
26 9 9 14 13 1 9 14 12 9 2 7 3 1 0 9 14 13 13 1 9 1 9 1 0 9 2
4 13 0 9 2
16 7 14 9 9 13 3 9 9 7 3 14 9 14 13 0 2
14 9 13 9 9 1 9 9 1 9 9 13 0 9 2
18 13 15 2 16 9 9 13 9 9 7 13 9 1 15 7 15 9 2
13 13 1 0 9 9 7 9 9 7 9 1 9 2
15 16 7 0 0 9 9 13 1 9 9 2 13 14 9 2
23 1 9 0 1 9 2 1 0 9 0 2 13 9 0 1 9 13 1 0 9 7 9 2
9 9 13 9 2 9 0 0 9 2
19 1 15 9 14 13 15 9 9 2 0 13 15 1 0 9 0 1 9 2
16 14 13 1 9 0 9 2 0 13 14 1 0 9 1 15 2
19 3 14 13 4 2 16 13 1 15 0 9 2 16 4 13 1 0 9 2
9 1 9 1 9 9 13 13 9 2
14 13 9 1 0 9 2 16 13 15 14 1 15 13 2
9 9 13 2 16 15 9 14 13 2
12 13 2 7 3 1 9 0 13 15 1 9 2
3 9 13 2
11 7 1 9 2 12 13 9 1 9 0 2
5 13 9 1 9 2
6 13 2 13 1 9 2
2 13 2
19 0 9 13 9 1 13 9 0 1 0 9 2 13 1 9 9 2 13 2
4 3 15 13 2
14 1 9 13 1 0 9 13 15 9 2 9 2 9 2
12 13 4 9 2 0 3 13 9 9 1 9 2
18 9 9 9 9 3 15 13 2 3 13 9 1 9 1 0 0 9 2
11 3 15 14 13 4 2 14 1 12 9 2
6 2 9 13 3 0 2
9 0 9 1 9 13 15 0 9 2
10 13 15 3 2 16 9 9 14 13 2
9 3 1 9 13 0 9 0 9 2
3 14 13 2
15 1 9 7 0 9 13 1 9 2 13 15 9 7 9 2
12 13 14 13 2 16 1 9 9 13 0 9 2
6 0 9 13 1 9 2
23 9 9 0 9 9 0 2 9 9 2 13 2 16 14 13 9 1 9 1 9 7 9 2
3 9 13 2
10 13 9 1 9 0 7 3 13 9 2
10 3 15 13 3 1 9 1 0 9 2
5 2 13 0 9 2
4 9 13 12 2
15 9 1 0 0 0 9 13 0 9 1 9 1 9 9 2
10 9 3 3 13 14 9 2 14 9 2
11 3 4 13 15 0 9 2 0 13 13 2
16 13 3 0 9 2 0 9 2 3 3 13 2 3 3 13 2
6 9 13 0 9 0 2
5 9 13 9 0 2
5 13 15 1 9 2
6 12 9 13 0 9 2
4 9 13 9 2
14 1 0 9 9 9 7 9 7 9 9 13 0 9 2
7 1 0 9 3 13 9 2
11 9 0 13 13 15 14 1 0 9 0 2
7 14 9 13 1 15 9 2
3 13 9 2
14 14 13 0 2 7 9 13 2 16 9 13 13 9 2
8 7 3 13 9 2 0 13 2
12 1 9 8 2 13 14 9 0 9 1 9 2
15 2 9 13 9 7 9 2 16 9 13 13 1 0 9 2
10 9 2 9 13 2 16 9 13 9 2
12 13 9 2 13 9 7 13 15 1 0 9 2
8 9 13 1 9 1 9 9 2
11 2 14 13 1 9 9 13 13 1 9 2
12 2 13 13 2 7 1 9 14 13 9 9 2
8 9 9 2 14 13 13 9 2
9 13 9 14 9 9 9 2 2 2
9 1 0 9 9 9 14 13 0 2
11 1 9 0 9 13 15 9 0 0 9 2
7 9 9 13 15 13 9 2
5 13 1 0 9 2
23 13 13 1 9 2 13 9 13 1 9 9 9 2 13 1 9 7 0 0 2 0 9 2
8 2 3 13 9 0 1 9 2
7 13 9 9 12 9 9 2
10 13 2 16 1 9 13 4 13 9 2
7 1 0 9 13 0 9 2
16 9 9 13 2 16 13 3 0 9 1 9 0 2 9 9 2
6 13 9 2 13 9 2
21 3 0 9 14 13 0 9 1 0 13 9 0 2 7 13 9 13 13 9 9 2
13 7 1 9 13 0 9 0 9 9 9 7 9 2
9 9 9 13 4 13 1 13 0 2
8 1 9 0 13 13 9 9 2
30 1 9 0 9 0 13 15 2 16 9 14 13 3 2 16 13 9 2 7 9 13 0 9 0 1 9 7 0 9 2
5 3 13 0 9 2
3 13 15 2
8 13 15 0 9 7 13 9 2
5 13 14 15 13 2
11 1 13 9 9 13 15 9 1 9 0 2
10 9 0 13 9 0 9 9 7 9 2
5 14 13 3 13 2
9 2 16 14 9 9 13 15 9 2
9 14 9 9 14 13 2 9 13 2
17 7 9 13 0 2 9 9 1 9 9 0 13 0 7 0 9 2
11 0 9 9 14 9 14 13 1 0 9 2
7 4 13 9 1 9 0 2
18 1 0 9 1 9 8 2 9 1 9 13 4 13 9 13 9 9 2
5 0 9 13 9 2
8 9 9 13 0 9 1 9 2
9 9 9 13 13 12 8 2 9 2
17 1 9 13 9 2 16 9 0 7 0 13 14 12 8 2 9 2
9 9 1 9 4 13 12 9 1 2
20 9 2 0 13 12 8 2 9 1 0 9 0 2 13 1 12 9 9 9 2
8 14 13 9 14 1 0 9 2
9 2 13 2 7 1 9 14 13 2
11 2 13 9 14 9 0 7 9 1 9 2
5 2 13 1 9 2
12 13 9 2 16 0 9 0 13 15 0 9 2
8 3 0 9 13 9 9 9 2
10 4 13 13 1 9 0 0 9 0 2
9 3 13 13 1 9 0 9 9 2
10 12 9 4 3 13 7 13 1 9 2
10 1 9 1 9 13 15 3 14 13 2
8 1 0 4 15 1 9 13 2
18 0 9 13 2 16 13 9 9 0 2 7 14 15 9 0 2 0 2
10 13 15 9 1 9 9 0 7 9 2
9 0 9 13 15 0 0 9 9 2
9 2 9 9 14 13 1 9 9 2
6 13 1 0 9 0 2
5 2 4 3 13 2
12 9 13 9 9 0 2 13 14 12 8 9 2
12 9 2 0 13 9 2 13 0 9 1 9 2
24 14 13 9 0 1 9 9 13 9 2 13 1 9 0 7 9 0 1 9 12 8 2 8 2
15 1 13 1 0 9 9 13 15 9 13 7 13 9 0 2
9 3 13 15 1 9 0 2 0 2
6 9 13 9 7 9 2
9 1 9 13 15 9 1 9 9 2
7 13 15 1 15 0 9 2
10 9 13 1 15 9 1 9 9 9 2
4 13 9 9 2
22 16 13 1 9 0 9 0 9 2 7 13 15 2 16 14 9 13 0 9 1 9 2
9 0 9 0 8 2 9 13 9 2
11 13 3 2 1 0 9 2 9 2 9 2
9 7 14 1 9 13 0 9 9 2
15 1 9 9 13 15 0 9 9 2 16 1 9 13 9 2
4 9 13 9 2
12 9 13 2 16 1 9 9 9 9 4 13 2
15 7 1 9 13 9 2 16 13 13 9 0 9 8 2 2
7 9 9 14 9 14 13 2
6 3 13 15 15 9 2
12 3 9 9 13 1 9 1 9 0 1 9 2
12 3 13 9 1 9 12 8 13 1 9 9 2
11 13 1 9 9 13 3 0 1 13 9 2
6 13 1 3 0 9 2
14 1 9 13 9 2 13 4 15 9 7 13 14 3 2
4 13 1 9 2
12 13 3 0 9 1 9 7 9 13 1 9 2
7 13 4 9 1 0 9 2
15 1 15 13 1 12 9 13 1 13 2 13 7 13 9 2
4 14 15 13 2
4 13 14 9 2
6 3 1 9 14 13 2
22 1 0 9 0 13 14 9 13 1 9 7 9 1 9 13 1 9 7 9 1 9 2
14 13 15 9 9 2 0 13 1 13 9 9 9 0 2
10 9 13 1 9 2 9 2 14 9 2
9 13 15 14 13 2 3 15 13 2
24 13 2 16 1 9 9 9 9 13 15 1 9 2 7 0 9 13 12 9 2 16 9 13 2
7 14 13 1 9 9 0 2
4 9 14 13 2
6 9 9 13 15 3 2
19 9 9 9 1 9 13 0 7 1 0 9 13 1 9 2 1 9 9 2
11 0 9 13 15 0 0 9 1 9 0 2
17 9 2 13 1 9 9 0 1 9 2 13 1 0 9 1 9 2
5 13 9 1 9 2
4 13 0 9 2
13 1 9 9 13 9 1 13 9 1 9 7 9 2
8 1 0 9 4 1 9 13 2
12 7 3 13 3 3 2 16 15 13 14 4 2
10 13 0 9 1 9 2 16 3 13 2
4 13 1 9 2
7 2 9 1 9 13 9 2
10 9 13 1 9 2 7 9 9 13 2
14 13 15 3 7 13 1 9 2 13 15 3 1 9 2
6 9 13 1 9 9 2
4 14 13 0 2
6 9 14 15 14 13 2
6 14 15 3 13 4 2
6 14 3 14 13 4 2
21 2 14 13 14 0 9 9 2 16 1 9 13 2 7 9 14 1 9 15 13 2
7 2 7 13 4 13 3 2
7 7 13 2 13 9 9 2
9 14 13 9 1 9 2 13 9 2
8 13 15 1 9 1 0 9 2
8 13 2 13 15 1 9 13 2
10 9 13 15 1 9 2 1 9 9 2
3 2 13 2
4 14 13 13 2
12 2 13 2 9 13 2 7 14 14 13 4 2
3 2 13 2
5 13 2 2 2 2
7 9 13 2 16 14 13 2
3 3 13 2
5 3 3 9 13 2
11 1 9 7 9 13 14 13 0 9 9 2
9 2 9 13 14 13 15 1 15 2
15 9 13 15 14 13 1 9 2 9 13 1 0 9 9 2
7 13 9 9 1 0 9 2
6 9 14 13 4 13 2
5 13 4 15 9 2
6 7 9 3 3 13 2
16 9 0 0 13 15 1 9 1 9 0 1 9 9 9 9 2
10 9 1 0 13 9 13 13 9 9 2
14 9 9 13 13 15 1 9 9 9 13 7 9 13 2
13 1 0 9 9 9 1 9 0 13 9 0 9 2
12 9 13 14 1 9 9 2 13 9 7 9 2
11 12 9 13 15 2 14 13 1 9 0 2
6 3 15 15 14 13 2
3 14 13 2
10 1 0 9 0 9 9 9 13 9 2
20 16 13 9 1 13 9 0 9 2 13 0 9 9 1 0 9 9 1 9 2
6 14 4 13 14 9 2
9 0 9 0 13 1 9 9 0 2
4 9 13 15 2
4 9 13 9 2
6 1 0 9 13 9 2
15 2 9 0 9 13 15 0 9 0 9 2 13 1 9 2
8 9 13 15 9 1 9 9 2
18 0 9 2 0 1 9 13 1 9 1 9 2 9 9 2 14 13 2
5 9 13 9 9 2
6 13 1 15 0 9 2
8 1 9 13 15 15 12 9 2
7 3 4 1 3 0 9 2
8 9 9 13 9 1 0 9 2
11 14 0 9 9 13 3 1 9 7 9 2
10 16 1 9 13 15 9 2 14 13 2
18 7 12 9 1 9 13 15 1 15 9 2 13 9 7 13 15 9 2
5 13 1 0 9 2
19 16 9 1 0 9 13 3 2 13 13 9 1 9 2 0 13 3 3 2
9 14 13 14 0 9 1 9 13 2
17 1 9 0 9 9 0 1 9 0 7 0 9 13 1 12 9 2
26 13 0 9 0 13 2 16 9 13 9 0 9 2 13 9 0 7 13 1 9 1 13 9 0 9 2
12 15 9 3 3 13 9 9 1 13 0 9 2
8 1 0 9 13 15 9 9 2
3 2 13 2
3 13 9 2
7 2 0 9 9 15 13 2
6 0 9 13 0 9 2
7 3 13 4 1 9 9 2
6 2 3 15 14 13 2
8 13 9 9 7 13 9 9 2
14 1 12 9 3 13 4 1 0 9 7 9 0 9 2
9 1 12 9 0 9 13 1 9 2
5 9 13 1 9 2
10 13 4 15 1 9 2 0 13 3 2
6 13 4 15 1 15 2
3 13 9 2
11 2 3 13 14 4 13 9 0 0 9 2
6 13 4 15 1 9 2
12 9 3 4 13 1 9 1 9 7 0 9 2
13 14 0 9 1 0 9 13 1 9 1 0 9 2
5 2 14 4 3 2
4 9 15 13 2
11 2 13 2 14 13 9 1 3 0 9 2
18 9 13 15 7 13 13 1 9 0 9 2 7 9 14 13 15 13 2
9 2 13 1 15 9 2 15 9 2
5 2 13 2 13 2
5 3 13 1 9 2
8 2 3 2 3 2 14 13 2
7 1 9 13 15 1 9 2
8 3 13 1 9 12 9 9 2
14 1 0 9 13 13 15 0 1 9 0 9 13 9 2
10 9 13 15 1 9 2 7 13 9 2
9 14 0 9 9 13 13 1 9 2
16 0 12 0 9 0 2 0 9 9 13 1 0 9 0 13 2
17 1 9 0 13 15 2 16 9 13 9 1 9 9 1 9 9 2
5 3 13 12 9 2
6 9 13 15 1 9 2
10 12 9 13 9 1 0 9 0 9 2
13 13 9 7 9 9 13 9 9 7 13 0 9 2
11 14 9 0 13 0 1 9 13 1 9 2
21 0 13 9 9 2 9 7 9 9 2 7 13 15 9 9 1 9 2 9 0 2
14 0 9 9 13 0 9 2 16 14 13 15 3 9 2
15 1 9 9 13 9 9 0 9 2 9 0 7 9 0 2
18 9 9 9 13 2 16 9 1 9 14 13 15 1 9 9 9 9 2
23 9 9 9 9 9 13 2 16 9 0 3 13 15 9 7 13 9 1 0 9 0 9 2
21 1 9 9 13 1 9 1 9 9 0 7 9 9 0 2 1 9 9 7 9 2
9 9 9 9 13 1 8 2 0 2
20 9 9 9 9 9 1 9 13 1 0 9 9 1 0 9 1 9 9 9 2
23 9 9 13 15 3 1 0 9 2 7 1 9 1 9 9 13 12 2 12 7 12 9 2
10 2 9 13 1 15 3 9 0 9 2
6 9 9 3 15 13 2
11 1 9 0 9 9 9 13 0 9 0 2
14 9 0 12 8 2 4 14 13 1 0 9 0 9 2
26 15 9 1 9 1 0 9 13 2 9 0 2 9 7 9 2 7 1 0 9 14 4 13 1 9 2
24 3 14 9 1 9 0 13 15 9 2 14 13 0 9 2 13 14 15 13 2 13 1 9 2
6 14 9 14 14 13 2
4 1 9 13 2
4 3 15 13 2
7 13 0 9 1 15 13 2
6 1 9 13 1 9 2
2 13 2
25 13 1 15 2 16 1 8 2 0 2 12 1 9 9 0 13 13 9 7 9 1 0 9 9 2
20 13 1 9 9 0 13 2 16 9 2 1 0 13 4 9 0 2 13 0 2
7 1 9 13 0 0 9 2
7 1 13 0 9 13 9 2
7 2 13 9 13 1 15 2
4 13 1 9 2
9 9 13 2 7 15 13 1 9 2
16 13 14 2 16 9 13 9 9 0 9 2 0 13 1 9 2
10 3 13 2 16 9 13 15 7 13 2
9 1 0 9 13 1 9 0 9 2
17 13 0 9 7 13 9 1 0 13 9 9 7 0 9 1 9 2
15 7 14 9 3 13 2 16 9 9 13 15 3 1 9 2
8 0 13 9 1 9 1 9 2
18 1 9 0 9 9 9 13 9 0 1 9 7 9 1 0 9 0 2
13 14 13 1 9 2 9 7 0 0 9 2 2 2
13 0 13 2 13 2 0 9 13 15 3 15 9 2
18 4 13 14 0 2 13 14 3 2 9 1 9 0 2 0 13 9 2
10 13 0 9 2 0 9 2 0 9 2
5 9 0 13 9 2
12 9 9 0 14 13 15 14 1 0 9 0 2
11 9 9 1 9 0 13 9 9 7 9 2
16 1 9 0 9 14 13 9 0 2 0 13 15 1 9 0 2
20 1 9 9 7 9 13 15 3 0 9 7 9 0 2 13 3 1 9 0 2
18 1 0 0 9 9 13 9 0 9 2 13 9 9 7 0 9 15 2
4 15 13 9 2
4 15 13 9 2
14 9 13 0 9 1 9 2 7 14 14 0 9 9 2
7 13 9 1 9 9 9 2
8 9 13 9 7 9 15 13 2
11 9 1 0 9 13 9 1 9 12 9 2
5 2 9 3 13 2
5 3 15 13 9 2
7 2 15 14 9 14 13 2
8 2 9 15 15 14 3 13 2
9 13 14 4 15 2 3 15 13 2
11 14 13 14 9 9 7 9 1 15 9 2
5 9 14 13 9 2
10 14 13 15 13 2 14 13 15 13 2
3 14 13 2
3 13 15 2
7 13 15 13 1 12 9 2
3 2 13 2
5 9 13 9 9 2
17 1 0 13 9 0 1 9 2 13 15 2 13 13 1 9 9 2
9 9 9 9 13 15 7 13 9 2
10 14 1 9 13 9 13 1 9 9 2
4 14 13 15 2
15 13 9 2 0 1 9 9 13 0 9 1 9 0 9 2
9 1 12 9 1 9 13 9 0 2
10 13 15 9 1 13 1 9 1 9 2
10 0 9 13 9 1 9 1 0 9 2
7 13 9 13 14 9 9 2
14 1 9 9 0 9 13 9 9 13 1 9 1 9 2
6 0 9 13 9 9 2
14 14 3 13 15 9 1 9 9 1 9 0 2 0 2
12 3 14 0 9 9 0 13 9 1 0 9 2
27 0 9 9 9 0 13 1 9 1 9 0 9 9 7 9 1 0 9 0 2 13 1 9 9 9 0 2
6 3 9 13 14 9 2
10 1 9 13 15 1 9 0 1 9 2
8 13 9 7 13 1 9 9 2
3 9 13 2
6 9 13 2 13 9 2
21 9 13 15 1 9 2 13 1 9 13 9 2 13 9 2 13 9 7 0 9 2
11 1 9 13 12 9 2 7 12 13 9 2
6 3 13 15 1 9 2
12 0 9 13 15 1 9 2 13 15 2 9 2
2 13 2
9 3 9 14 13 9 1 0 9 2
13 1 0 9 2 9 13 1 9 9 1 9 9 2
3 13 9 2
12 2 9 13 3 0 2 16 13 0 9 2 2
3 13 9 2
4 2 9 13 2
3 2 13 2
4 2 9 13 2
5 13 9 2 2 2
13 13 2 16 1 9 13 15 9 7 13 0 9 2
5 9 13 1 9 2
5 13 1 15 3 2
18 1 9 13 15 1 9 0 9 1 3 0 9 7 0 2 0 9 2
7 13 0 9 7 0 9 2
12 13 14 3 2 7 3 1 15 13 0 9 2
5 9 13 3 0 2
16 1 9 13 0 9 2 0 1 0 9 1 0 9 7 9 2
8 15 14 13 1 9 9 0 2
5 9 13 15 9 2
13 15 9 13 3 9 2 7 3 3 13 15 13 2
11 1 0 9 13 1 15 9 1 0 9 2
6 0 9 13 15 9 2
9 16 9 13 2 13 15 9 0 2
7 2 9 13 1 15 0 2
12 9 13 9 0 9 9 2 13 15 15 9 2
9 3 13 3 0 9 0 1 9 2
10 13 15 0 9 9 13 15 9 0 2
14 13 4 13 2 16 9 1 0 9 14 13 13 0 2
15 9 13 13 9 7 15 3 1 0 0 9 13 0 9 2
5 2 16 15 13 2
12 14 13 1 9 9 1 9 15 13 2 2 2
16 1 0 9 13 4 13 14 0 9 2 0 13 0 9 9 2
11 1 12 9 1 9 9 13 15 13 9 2
11 0 9 13 15 3 0 9 1 9 0 2
18 1 9 9 7 9 9 2 9 8 13 13 1 9 13 3 9 9 2
13 9 13 9 1 13 9 9 1 13 0 9 9 2
12 9 1 0 9 0 13 9 1 9 7 9 2
10 1 9 1 0 9 0 13 13 9 2
9 9 13 3 13 9 7 9 0 2
7 13 4 15 3 1 15 2
13 13 9 3 0 2 13 4 14 13 1 0 9 2
17 13 1 9 7 14 13 2 16 9 13 2 16 13 0 0 9 2
7 9 13 13 9 1 9 2
9 7 3 13 13 1 9 1 9 2
17 9 2 3 13 9 0 2 1 0 9 13 2 16 3 13 9 2
7 2 13 15 0 9 2 2
27 13 1 9 2 1 9 13 15 1 9 2 9 2 0 13 15 9 1 9 13 1 13 1 9 1 9 2
8 2 9 13 15 14 9 2 2
9 1 9 9 14 13 15 9 9 2
7 1 15 9 9 13 9 2
7 13 4 9 2 0 9 2
16 9 14 13 13 0 9 2 7 14 14 13 13 9 1 9 2
10 14 13 9 9 2 13 15 14 9 2
9 13 9 2 0 9 2 0 9 2
14 14 13 15 13 9 2 13 14 2 16 9 13 0 2
8 13 15 2 16 13 15 9 2
10 14 1 0 9 9 0 13 9 9 2
8 9 0 13 7 3 9 9 2
11 9 13 0 9 13 9 9 9 1 9 2
7 9 13 13 1 9 9 2
7 4 13 3 0 9 9 2
25 16 9 13 1 15 9 2 7 0 9 13 13 1 12 9 1 13 9 9 1 9 0 9 0 2
7 3 13 15 9 1 9 2
6 14 9 13 1 9 2
7 3 7 13 9 1 9 2
16 0 9 14 13 1 9 7 13 13 1 0 9 13 1 9 2
6 13 15 9 1 9 2
19 16 13 2 16 9 3 13 9 0 1 9 2 13 13 0 9 7 9 2
12 16 14 13 9 2 9 4 14 14 3 13 2
7 0 9 13 9 7 9 2
8 13 15 9 2 13 13 9 2
5 13 15 14 9 2
9 2 7 0 9 13 13 0 9 2
6 1 9 15 14 13 2
4 14 13 9 2
21 13 9 9 14 13 9 9 2 16 1 0 9 9 9 13 15 15 1 9 0 2
15 1 9 9 9 13 14 14 13 12 9 0 7 12 0 2
3 7 13 2
21 13 3 9 9 2 9 9 2 9 9 2 9 9 2 9 9 7 13 9 9 2
3 9 13 2
11 9 0 9 0 13 1 9 1 9 9 2
9 0 9 9 13 14 0 0 9 2
10 0 9 13 15 9 1 9 1 9 2
6 7 0 9 13 0 2
11 2 15 13 9 9 1 9 3 1 9 2
6 7 1 9 13 9 2
8 2 1 0 9 13 9 9 2
5 2 14 3 13 2
7 15 14 13 3 13 9 2
11 13 3 9 2 13 3 13 1 15 9 2
11 13 15 15 2 7 3 14 13 1 15 2
12 9 1 0 9 13 0 7 13 15 15 3 2
9 13 15 2 9 2 9 0 9 2
11 9 3 1 15 13 14 15 13 1 9 2
12 14 0 0 9 13 15 1 9 9 1 9 2
8 13 15 1 9 14 1 9 2
4 13 2 9 2
18 9 13 14 9 9 2 1 0 9 0 0 15 13 9 3 0 9 2
13 9 1 0 9 13 15 2 16 3 1 9 13 2
8 9 3 13 9 3 13 9 2
3 13 9 2
5 9 13 15 3 2
8 9 0 9 13 15 0 9 2
5 9 13 1 9 2
8 9 13 2 3 13 1 15 2
27 1 0 9 1 9 2 13 1 9 2 13 0 9 0 9 2 13 15 1 0 9 0 9 9 9 0 2
12 9 13 0 9 1 0 9 7 9 0 9 2
12 9 9 0 13 0 3 9 9 2 9 9 2
10 0 9 15 13 2 0 9 15 13 2
16 7 9 15 13 2 16 14 13 15 0 9 2 15 0 9 2
23 7 14 1 3 1 9 0 9 1 0 9 13 9 9 2 1 0 13 1 9 9 0 2
13 0 9 9 13 13 9 0 1 9 1 9 9 2
9 3 9 0 9 13 9 0 9 2
8 13 1 9 9 1 9 9 2
24 0 9 13 14 13 15 1 9 2 13 14 13 0 0 9 2 14 9 14 13 14 0 0 2
4 2 13 2 2
12 13 2 16 13 9 7 15 9 13 1 9 2
7 0 9 9 13 14 9 2
13 13 1 9 2 3 14 13 13 1 15 0 9 2
20 9 1 9 9 9 3 3 13 9 9 0 2 7 1 9 0 9 14 13 2
28 1 15 0 9 1 0 9 13 15 0 9 2 0 9 0 2 1 13 0 7 0 3 9 2 13 14 0 2
6 9 3 13 0 9 2
8 13 15 7 14 13 0 9 2
9 9 13 1 9 0 9 1 9 2
9 9 14 13 14 1 9 2 2 2
7 14 9 13 13 9 0 2
7 14 9 0 13 13 9 2
5 3 9 13 3 2
6 14 13 0 0 9 2
12 2 13 1 9 2 16 13 0 1 9 9 2
4 9 14 13 2
4 15 13 0 2
6 2 14 9 13 0 2
5 2 13 9 0 2
10 2 3 3 9 15 1 15 14 13 2
16 9 13 15 9 2 1 9 1 0 9 1 9 13 0 9 2
6 13 2 14 13 9 2
7 2 13 15 9 7 9 2
10 12 8 2 9 13 1 9 1 9 2
9 14 1 12 9 4 13 1 9 2
20 1 0 9 9 4 13 7 14 13 9 1 0 9 2 1 0 12 13 13 2
9 3 4 13 1 9 7 9 0 2
16 0 9 1 0 9 13 3 12 9 9 1 13 9 9 9 2
4 13 15 9 2
15 4 7 3 13 2 3 13 1 9 2 7 1 9 13 2
23 13 15 1 15 2 13 9 0 9 2 16 13 15 0 9 2 13 3 15 9 1 9 2
4 13 0 9 2
15 15 13 1 0 9 2 0 15 13 2 0 1 9 13 2
23 3 9 13 0 0 9 3 1 15 7 13 1 9 0 2 7 4 3 9 7 9 9 2
19 9 13 15 1 15 3 3 2 16 14 1 0 2 9 9 9 13 9 2
30 1 9 0 9 9 14 3 13 1 0 9 2 9 1 9 9 0 13 1 9 2 7 0 13 2 13 9 1 9 2
15 1 3 13 9 13 9 7 14 3 13 1 15 0 9 2
11 13 9 0 2 14 1 9 13 1 9 2
10 1 0 9 4 13 3 13 9 9 2
17 9 0 0 13 0 0 9 2 7 14 14 4 9 9 15 9 2
11 9 13 1 9 13 13 1 9 9 0 2
13 9 13 1 9 12 9 13 9 13 1 13 9 2
15 14 13 13 9 1 9 0 1 9 13 9 7 9 13 2
7 0 13 14 9 0 9 2
11 0 9 9 14 13 9 13 3 1 9 2
7 1 9 13 4 9 0 2
23 9 13 9 1 9 9 13 1 0 9 2 0 14 1 9 1 9 13 13 1 0 9 2
9 1 9 0 9 13 15 9 9 2
7 0 15 13 9 1 9 2
12 9 13 9 7 13 15 1 9 1 9 0 2
5 9 13 3 9 2
10 3 1 9 13 9 9 7 13 3 2
4 9 13 9 2
3 13 4 2
5 9 13 1 9 2
4 2 14 13 2
4 9 13 15 2
7 13 9 7 13 9 9 2
6 14 9 13 14 13 2
4 9 13 3 2
6 9 13 15 1 9 2
4 13 15 2 2
8 9 13 15 0 2 0 9 2
12 13 15 1 9 7 13 1 9 1 0 9 2
3 2 13 2
6 13 2 16 9 13 2
7 9 13 1 9 7 9 2
12 2 13 0 9 2 13 15 1 15 3 13 2
4 9 13 9 2
12 15 9 13 13 9 9 1 9 9 7 9 2
10 9 13 14 12 9 1 9 7 9 2
14 9 4 9 9 9 2 9 7 9 9 1 9 9 2
5 3 13 0 9 2
6 3 9 9 14 13 2
5 3 9 14 13 2
5 3 9 3 13 2
6 3 0 9 13 9 2
7 13 15 13 1 12 9 2
5 13 2 9 13 2
12 2 9 2 13 2 13 0 9 2 2 2 2
11 2 13 2 3 9 0 13 2 2 2 2
8 1 9 13 14 0 9 13 2
11 13 4 2 16 9 13 3 13 0 9 2
13 3 13 2 16 9 14 13 15 1 0 0 9 2
10 13 9 9 1 9 7 13 15 9 2
4 2 3 13 2
6 7 3 1 9 13 2
15 9 0 9 0 7 9 0 9 0 13 9 9 0 9 2
13 9 13 9 2 13 9 1 9 7 13 9 9 2
24 9 9 0 13 1 9 9 9 9 1 9 2 9 9 7 9 2 7 14 9 1 0 9 2
16 9 13 1 9 9 13 14 0 9 1 9 13 1 9 9 2
14 13 13 1 9 0 9 9 9 2 3 1 9 9 2
11 9 9 3 13 1 9 9 7 9 9 2
22 0 9 13 1 9 0 9 0 2 0 9 13 0 9 9 2 9 0 7 0 9 2
11 9 0 4 14 13 1 9 9 7 9 2
8 3 0 9 9 13 9 0 2
9 13 15 1 15 3 9 7 9 2
15 1 9 0 9 13 9 0 2 0 13 13 1 9 0 2
17 9 1 9 9 1 9 9 13 0 9 7 13 0 9 1 9 2
13 1 0 9 1 9 13 14 14 12 8 2 9 2
14 13 7 9 2 0 9 14 13 1 9 1 0 9 2
6 9 4 13 1 9 2
18 1 0 9 14 13 2 13 2 16 14 13 13 9 1 9 1 9 2
6 13 15 3 0 9 2
21 13 0 0 1 12 9 9 1 9 1 0 9 2 13 12 9 2 13 9 9 2
8 13 3 1 9 14 1 9 2
8 7 7 3 3 13 15 9 2
26 13 15 15 14 2 16 1 9 0 9 2 1 9 13 14 9 9 0 2 13 15 9 1 0 9 2
16 13 9 1 9 0 9 9 0 1 9 0 13 9 0 9 2
13 13 2 16 14 1 9 0 9 13 1 13 9 2
7 9 1 13 9 13 3 2
9 9 4 13 3 0 9 0 9 2
10 9 0 4 13 1 9 9 9 0 2
15 9 13 2 16 13 0 9 0 9 2 0 14 13 3 2
7 0 9 13 14 1 9 2
19 2 9 13 2 16 9 0 1 9 9 1 9 13 1 9 1 0 2 2
10 1 15 9 13 13 9 0 9 9 2
22 13 15 1 9 2 16 0 9 13 13 0 9 1 12 9 9 0 2 13 1 15 2
8 14 13 1 15 1 12 9 2
16 13 2 16 14 13 9 1 9 2 16 14 13 14 15 13 2
11 14 4 9 0 9 1 9 1 0 9 2
9 3 1 9 9 9 9 13 0 2
11 13 2 16 9 9 9 9 9 0 13 2
6 9 13 15 1 9 2
5 2 9 13 0 2
11 2 13 9 9 1 13 9 1 9 0 2
11 1 9 1 13 0 9 1 0 13 9 2
17 1 9 13 9 1 13 9 9 1 9 9 9 0 1 0 8 2
4 13 1 13 2
12 2 13 1 13 1 9 9 0 1 0 8 2
14 16 14 1 9 13 15 9 2 7 13 14 15 0 2
5 2 9 13 0 2
5 9 0 13 12 2
6 9 13 15 1 9 2
5 14 13 9 9 2
5 13 1 0 9 2
8 13 15 2 14 13 9 9 2
17 1 9 13 13 2 16 9 9 0 13 1 13 9 1 0 9 2
10 2 14 9 4 13 1 12 9 3 2
5 2 13 2 13 2
6 2 14 9 9 13 2
6 13 1 13 9 9 2
8 2 13 2 16 9 9 13 2
7 2 13 9 2 9 9 2
7 9 13 1 13 0 9 2
4 13 1 9 2
12 2 13 2 16 9 9 1 13 9 9 13 2
2 13 2
6 2 13 2 9 9 2
12 13 4 3 1 9 13 1 0 9 9 0 2
4 13 1 9 2
18 2 13 3 2 16 1 9 0 13 0 9 1 13 9 0 9 2 2
11 1 9 13 13 9 9 0 1 9 0 2
5 13 3 13 9 2
4 2 13 9 2
6 1 9 13 3 3 2
8 13 1 9 1 9 9 9 2
12 2 13 2 16 9 9 1 8 2 0 13 2
13 13 2 14 1 9 9 9 13 1 12 9 9 2
17 13 4 13 1 9 2 1 0 13 15 9 2 13 15 13 9 2
6 2 13 2 9 9 2
10 13 3 2 9 9 9 9 1 9 2
16 9 9 13 14 14 13 9 2 3 13 9 1 9 9 0 2
15 2 14 9 1 9 7 9 9 13 13 9 1 0 9 2
38 2 16 9 9 14 13 9 9 0 1 0 9 7 15 9 2 13 2 16 13 15 1 15 13 2 16 13 15 9 0 7 14 13 2 1 9 13 2
19 9 0 9 13 2 16 12 0 9 13 1 9 1 9 7 13 1 9 2
10 0 9 13 1 9 0 13 1 9 2
19 1 9 13 9 1 0 9 0 9 0 9 2 9 0 2 9 9 9 2
14 0 13 9 9 9 2 9 7 9 9 9 9 9 2
19 9 9 7 15 9 13 0 1 9 9 2 9 13 14 1 9 1 9 2
7 1 9 9 9 14 13 2
12 13 1 15 2 13 9 2 13 9 0 9 2
11 13 14 14 0 9 1 9 1 0 9 2
16 13 15 1 1 9 2 13 2 16 9 15 13 14 13 0 2
17 9 13 15 1 9 1 9 2 0 0 0 9 2 1 9 9 2
15 3 1 0 9 13 9 7 9 2 7 14 0 9 9 2
12 13 15 9 14 9 9 2 9 7 9 9 2
7 9 2 13 4 1 9 2
3 7 13 2
8 9 14 13 14 1 0 9 2
6 13 1 0 0 9 2
8 13 0 2 0 9 1 9 2
5 14 13 15 9 2
7 14 13 13 15 0 9 2
3 9 13 2
4 14 13 9 2
9 14 13 0 9 7 14 14 4 2
10 13 15 9 7 13 13 15 0 9 2
14 1 9 9 13 9 2 13 3 2 16 9 14 13 2
28 15 9 13 1 0 9 9 2 0 1 9 14 13 2 7 0 9 13 3 9 1 9 9 9 7 14 9 2
7 9 13 12 9 1 9 2
10 14 13 9 14 2 16 13 15 13 2
11 9 2 9 7 9 13 0 9 9 9 2
4 9 13 0 2
10 14 13 1 9 2 15 9 7 9 2
9 7 9 1 15 14 13 15 0 2
5 0 13 1 9 2
7 14 9 9 0 13 9 2
13 13 9 9 1 9 2 7 9 13 15 1 9 2
5 9 3 14 13 2
7 13 0 9 13 9 9 2
10 7 0 9 13 15 13 1 9 9 2
11 7 9 14 13 2 16 9 13 1 9 2
9 13 4 15 1 9 7 13 4 2
8 0 13 7 13 15 1 9 2
8 13 9 2 13 7 13 13 2
13 9 9 13 4 15 1 9 7 13 4 1 9 2
22 13 15 0 9 7 9 2 7 1 0 9 9 13 15 9 9 1 0 2 0 9 2
12 2 3 1 0 13 1 9 1 9 9 2 2
6 9 13 13 0 9 2
14 13 15 1 9 0 2 0 9 7 13 9 1 9 2
4 1 9 13 2
10 13 1 9 2 13 7 13 9 9 2
7 2 13 15 2 16 13 2
24 1 9 0 2 0 1 9 2 0 13 12 9 1 0 9 2 9 13 4 1 0 9 9 2
11 0 2 3 0 2 9 13 9 9 0 2
20 16 14 13 0 9 2 13 15 2 9 13 13 0 9 13 1 9 1 0 2
19 3 1 9 14 12 9 13 1 9 0 2 7 8 2 12 8 13 9 2
17 9 1 3 0 9 13 13 1 9 9 7 0 1 9 9 0 2
6 13 7 13 15 9 2
13 13 9 14 13 2 16 9 9 13 1 9 9 2
10 9 9 13 13 2 3 0 2 0 2
5 14 13 15 9 2
10 9 9 13 0 9 7 9 1 9 2
7 3 13 1 9 1 9 2
8 9 1 9 13 15 0 9 2
9 1 9 13 15 9 9 9 9 2
12 9 13 1 9 9 2 9 13 1 9 3 2
14 1 9 0 9 9 7 0 9 13 3 9 0 9 2
18 13 9 9 2 13 9 1 0 9 2 0 13 13 1 15 9 9 2
12 9 14 13 9 1 9 2 16 13 1 9 2
25 3 13 15 1 9 1 9 2 3 9 13 0 9 2 9 13 9 2 16 13 15 1 0 9 2
8 2 9 14 13 13 1 9 2
8 7 9 13 3 3 3 0 2
4 2 3 13 2
5 2 7 9 13 2
6 13 14 9 0 9 2
16 1 9 0 13 0 9 9 13 2 3 13 2 0 9 0 2
10 0 9 1 9 0 13 9 9 0 2
15 0 9 0 9 1 0 9 9 13 7 13 9 9 9 2
5 9 13 15 9 2
23 9 1 9 9 13 14 12 9 9 2 13 15 1 0 0 9 2 13 1 15 0 9 2
7 0 9 13 0 7 0 2
15 0 9 13 9 13 15 1 0 9 9 1 0 0 9 2
6 9 13 14 9 9 2
9 13 3 2 13 0 2 0 9 2
14 9 13 1 9 12 9 2 12 9 1 13 1 9 2
12 13 9 9 9 7 0 9 0 1 15 9 2
18 9 13 9 2 16 12 0 9 9 13 13 15 3 1 12 0 9 2
19 1 13 15 1 9 0 9 9 0 9 13 3 13 9 14 1 0 9 2
9 9 13 1 15 9 13 9 0 2
15 1 9 13 14 13 0 9 1 9 0 9 1 9 0 2
11 9 2 1 9 2 9 0 9 13 9 2
17 16 9 13 1 9 9 9 2 9 14 13 9 1 0 0 9 2
8 9 13 15 9 13 0 9 2
17 13 15 15 1 0 9 7 0 9 2 13 13 1 0 9 9 2
19 1 0 9 9 13 13 1 9 9 0 9 1 9 0 9 9 7 9 2
23 0 0 2 0 9 13 9 9 9 9 9 2 7 1 9 15 9 13 15 1 0 9 2
9 1 9 1 9 13 3 13 9 2
10 13 3 9 3 0 2 13 1 9 2
7 13 9 2 16 15 13 2
8 9 13 9 2 13 9 0 2
14 9 9 0 13 1 13 9 13 9 3 1 15 9 2
10 1 9 9 13 9 13 12 9 9 2
21 13 9 3 0 1 9 2 0 0 13 9 2 16 13 13 1 9 0 0 9 2
11 9 13 14 13 9 1 12 9 1 9 2
14 9 13 1 9 13 4 3 13 1 12 9 1 9 2
23 13 9 2 16 9 9 3 3 13 1 9 7 13 13 15 0 9 7 9 1 15 9 2
15 9 9 9 13 1 0 9 0 9 2 0 14 9 13 2
9 2 1 9 13 4 3 0 2 2
10 2 1 9 13 4 3 0 9 2 2
9 2 1 9 4 4 3 13 2 2
11 2 1 9 4 4 3 13 7 13 2 2
9 2 1 9 3 4 4 13 2 2
16 2 1 9 4 4 3 13 1 9 2 7 9 15 13 2 2
9 9 0 13 1 9 13 9 0 2
14 1 12 9 1 0 2 0 9 9 13 0 9 0 2
11 1 9 0 1 9 9 0 13 15 9 2
12 9 13 9 13 1 9 9 9 14 0 9 2
7 13 2 13 9 0 9 2
13 9 7 15 0 9 4 13 1 9 0 2 0 2
8 9 9 0 9 0 9 13 2
7 13 9 12 3 0 9 2
7 15 13 13 9 0 9 2
8 13 15 1 9 9 1 9 2
5 13 1 9 13 2
11 12 8 9 7 9 13 1 0 9 9 2
12 9 4 13 1 9 2 0 13 9 0 9 2
6 13 14 3 0 9 2
13 13 14 13 2 16 12 9 13 15 1 0 9 2
5 0 13 9 9 2
16 9 13 0 9 2 16 13 9 13 9 1 0 2 0 9 2
21 13 1 9 2 16 1 9 9 14 13 9 9 2 7 9 9 13 1 15 9 2
9 13 1 9 14 9 0 1 13 2
6 1 9 14 13 9 2
8 1 9 14 9 13 0 9 2
12 9 0 9 14 13 9 2 9 7 0 9 2
6 13 14 12 9 9 2
9 14 9 9 7 0 9 13 9 2
14 0 9 0 7 9 3 13 0 9 0 9 9 9 2
8 0 9 13 3 12 8 3 2
12 1 9 0 9 9 9 7 9 13 0 9 2
16 9 9 13 1 0 9 7 9 1 0 9 2 7 13 9 2
13 2 14 1 9 13 9 0 9 1 9 7 9 2
19 2 9 1 9 9 9 13 2 16 9 9 13 1 9 0 2 1 9 2
6 7 14 13 0 9 2
9 7 13 1 0 9 1 0 9 2
5 7 0 9 13 2
11 9 9 9 13 7 9 1 9 14 13 2
4 9 13 9 2
4 13 0 9 2
12 13 9 1 9 2 3 3 0 1 0 9 2
22 16 14 9 0 14 13 15 13 0 0 9 2 13 0 9 1 9 9 13 0 9 2
6 1 9 14 13 9 2
5 9 13 9 9 2
4 9 13 9 2
15 2 13 9 1 9 13 2 16 9 13 9 9 1 15 2
13 9 13 4 9 0 9 2 0 13 1 9 9 2
6 13 4 12 8 9 2
10 9 13 15 9 1 0 9 1 0 2
6 13 9 2 9 9 2
14 1 9 9 2 1 13 9 9 9 13 9 0 9 2
7 9 0 13 9 9 0 2
9 3 1 0 9 13 15 0 9 2
7 9 13 15 2 13 9 2
4 9 15 13 2
6 9 13 1 0 9 2
27 13 2 16 1 0 9 9 8 2 13 9 9 1 9 0 9 0 1 9 0 1 0 9 9 1 9 2
22 9 0 9 13 13 0 9 1 9 1 9 2 1 9 9 9 1 0 9 1 9 2
5 13 13 1 9 2
9 16 13 2 13 1 15 1 9 2
6 9 13 1 9 0 2
11 2 13 4 15 1 9 9 1 2 2 2
8 2 14 13 13 9 1 9 2
14 2 15 9 13 3 14 0 2 9 13 3 0 9 2
12 2 13 14 0 9 2 7 14 14 13 9 2
9 14 2 3 13 1 9 9 0 2
9 1 13 9 9 13 14 12 8 2
11 9 13 9 2 0 1 9 13 0 9 2
18 1 9 9 1 9 9 0 2 0 7 13 9 13 9 9 9 9 2
13 14 1 9 9 0 2 9 1 15 13 3 13 2
20 0 9 1 9 4 13 1 9 0 9 0 1 9 1 9 1 9 1 9 2
16 3 3 13 4 2 7 0 9 2 0 13 3 2 13 9 2
18 2 13 1 9 9 2 13 9 2 0 1 0 9 13 0 0 9 2
16 0 7 0 9 13 0 9 2 13 1 9 7 0 0 9 2
9 13 9 3 2 13 15 1 9 2
17 13 1 9 2 13 4 0 0 9 7 9 1 0 9 1 9 2
7 13 1 0 9 1 9 2
3 9 13 2
10 14 13 15 9 1 9 13 2 13 2
6 13 1 9 13 9 2
9 3 13 14 4 9 13 1 9 2
10 2 14 13 4 2 16 13 9 9 2
11 9 13 1 9 0 2 13 15 7 13 2
3 3 13 2
4 7 14 13 2
8 13 14 14 9 1 0 9 2
11 9 0 1 9 3 13 9 1 0 9 2
31 16 3 13 1 9 7 13 15 1 9 2 9 1 9 14 14 13 2 3 14 13 15 15 13 13 15 1 15 1 9 2
3 13 9 2
6 14 3 13 1 9 2
2 13 2
5 0 9 13 9 2
7 9 9 9 9 14 13 2
3 13 15 2
7 0 13 3 0 13 9 2
12 1 0 13 9 9 0 4 3 13 1 13 2
5 2 14 13 15 2
5 3 15 13 3 2
15 2 9 13 1 9 2 0 1 9 3 13 1 9 9 2
4 2 13 4 2
6 13 4 9 1 9 2
5 14 15 13 13 2
8 2 7 3 13 9 0 9 2
13 15 13 2 16 13 15 2 16 9 13 0 9 2
6 2 16 13 1 9 2
9 0 9 9 13 13 9 1 9 2
11 3 9 13 9 9 7 13 15 1 9 2
9 1 9 4 15 13 1 9 9 2
8 2 3 13 4 15 1 15 2
8 13 15 2 16 9 13 9 2
3 13 3 2
4 2 9 13 2
15 9 13 9 2 13 1 0 9 2 1 0 13 0 9 2
4 14 13 9 2
4 7 13 9 2
3 2 13 2
5 2 13 2 13 2
7 3 13 4 14 13 9 2
7 2 13 2 16 13 13 2
7 2 13 1 15 9 0 2
7 0 9 2 13 15 13 2
6 16 15 0 9 13 2
3 13 15 2
5 13 9 1 9 2
2 13 2
4 13 15 9 2
13 13 2 16 0 0 2 0 9 13 1 0 9 2
10 13 9 2 3 14 13 3 9 0 2
14 1 0 9 13 2 16 9 9 1 9 13 12 8 2
7 9 9 13 1 0 9 2
10 0 9 2 14 2 13 1 0 9 2
10 9 1 9 13 1 13 1 9 0 2
10 9 13 2 16 13 1 3 0 9 2
15 13 2 16 13 9 3 2 16 13 4 1 15 3 13 2
9 9 0 13 0 9 9 9 0 2
9 0 9 13 9 1 1 9 0 2
10 9 9 2 9 9 2 13 9 9 2
20 13 1 9 2 7 1 0 0 9 2 1 12 9 2 13 14 9 7 9 2
8 7 9 15 14 13 2 2 2
9 0 13 9 9 2 13 9 9 2
18 1 9 9 0 13 0 9 2 7 1 15 0 9 3 13 15 9 2
10 7 9 3 1 9 14 13 2 2 2
8 9 13 4 9 2 2 2 2
14 1 0 9 2 13 1 0 9 0 2 13 0 9 2
7 9 13 0 9 7 9 2
16 4 13 0 9 2 7 1 13 3 0 9 0 13 15 13 2
29 13 13 2 16 9 13 0 9 9 2 16 1 0 9 9 1 0 9 13 14 1 9 9 7 0 9 0 9 2
14 1 9 1 9 7 9 13 9 7 13 15 9 9 2
19 3 9 13 15 9 2 7 9 15 13 2 1 0 9 2 7 13 9 2
15 9 2 1 9 0 2 13 9 9 2 9 0 1 9 2
10 3 2 1 0 9 13 9 9 9 2
6 9 13 0 9 9 2
16 0 9 9 2 13 14 9 0 2 13 0 1 9 9 9 2
4 9 13 13 2
9 14 3 0 13 9 9 1 9 2
8 1 0 14 13 0 9 9 2
11 9 13 9 2 9 7 9 1 12 9 2
11 1 9 13 15 14 13 1 9 9 0 2
10 1 9 0 7 9 0 13 13 9 2
10 1 0 9 1 0 9 13 15 9 2
7 9 13 9 1 9 0 2
19 9 13 9 0 13 3 0 0 9 2 0 13 13 15 1 12 9 9 2
8 9 9 13 13 0 0 9 2
9 9 9 0 13 0 9 1 9 2
6 9 13 9 7 13 2
10 9 7 13 3 14 12 1 9 9 2
19 1 15 9 2 0 1 9 13 7 0 2 13 1 9 0 2 0 9 2
19 9 9 0 1 9 9 13 2 16 1 9 9 3 13 4 9 9 0 2
23 9 9 1 9 14 13 13 1 9 9 7 13 0 9 1 9 3 1 9 9 9 9 2
5 14 13 13 9 2
7 9 14 13 1 0 9 2
14 9 9 13 7 3 14 1 9 9 14 13 9 0 2
17 13 4 15 1 15 1 0 9 2 3 7 14 13 13 1 9 2
10 13 9 7 13 0 9 1 0 9 2
15 0 9 13 9 2 1 16 13 9 13 9 1 9 0 2
6 3 13 15 0 9 2
16 13 9 2 16 15 3 13 7 1 0 9 0 9 13 9 2
4 2 9 13 2
7 13 15 1 9 1 9 2
3 12 13 2
5 13 1 9 9 2
5 2 9 9 13 2
15 13 15 14 13 2 9 0 9 3 13 1 9 7 9 2
11 13 15 0 9 2 14 13 1 9 0 2
10 1 9 13 3 2 7 13 0 9 2
20 0 9 13 4 13 1 9 9 2 0 13 2 16 13 9 1 9 0 9 2
12 9 1 0 9 1 9 13 1 0 9 0 2
5 9 13 9 9 2
7 13 13 0 0 9 9 2
9 14 3 1 9 13 4 0 9 2
8 9 15 3 13 1 9 9 2
6 9 1 0 13 9 2
9 14 0 9 1 15 9 13 0 2
8 9 13 3 1 12 9 9 2
11 9 13 4 3 1 9 1 9 0 9 2
10 9 1 9 9 9 0 14 13 9 2
14 9 13 1 9 1 9 13 14 3 9 0 7 0 2
7 9 0 9 9 13 9 2
18 16 3 14 4 13 3 9 9 0 2 13 13 9 1 9 15 9 2
9 0 9 13 3 13 14 9 13 2
9 16 15 13 1 9 2 13 13 2
12 9 14 3 13 9 2 16 4 13 0 9 2
4 12 13 9 2
8 14 13 4 0 9 1 9 2
3 13 12 2
4 13 12 9 2
3 14 13 2
5 1 12 9 13 2
6 13 1 9 7 13 2
8 9 9 14 13 7 13 9 2
3 14 13 2
13 1 9 0 8 2 9 1 9 13 15 3 0 2
17 3 1 9 0 13 1 9 13 13 15 3 1 0 8 2 9 2
7 0 13 4 1 0 9 2
10 13 3 2 1 9 13 15 1 9 2
5 14 13 1 15 2
4 14 13 9 2
7 2 9 9 14 14 13 2
8 13 9 13 14 1 0 9 2
4 2 7 13 2
6 2 13 9 2 9 2
11 9 13 9 1 12 9 1 9 15 13 2
6 1 9 13 7 13 2
8 9 7 9 13 15 13 9 2
4 9 13 15 2
11 9 9 9 1 9 0 13 13 3 0 2
10 7 9 1 13 9 1 15 14 13 2
8 2 3 13 9 1 9 13 2
5 2 13 15 13 2
5 2 7 9 13 2
9 7 3 13 15 1 9 1 9 2
11 2 9 13 9 1 9 2 0 13 15 2
11 1 0 9 13 15 1 9 7 3 13 2
26 9 9 9 13 3 0 9 13 1 0 9 2 7 1 15 9 13 4 13 2 16 0 9 15 13 2
6 9 3 13 1 9 2
5 9 14 15 13 2
17 9 13 15 1 15 1 9 2 13 1 0 0 9 0 0 9 2
11 9 13 15 1 9 2 13 13 9 9 2
6 13 15 9 13 15 2
8 2 13 2 9 13 0 9 2
6 15 14 4 13 13 2
9 2 14 9 13 2 9 13 2 2
5 2 15 13 9 2
12 16 4 13 9 2 7 13 14 4 1 9 2
4 13 15 13 2
12 16 9 13 2 13 13 0 9 1 0 9 2
18 9 13 14 0 9 2 0 13 1 9 2 1 0 13 15 9 0 2
9 1 9 1 9 4 13 1 9 2
12 7 3 9 9 1 9 13 1 9 0 9 2
10 9 1 15 9 14 3 13 13 0 2
10 13 9 7 1 15 13 15 0 9 2
6 2 13 4 3 0 2
5 2 3 14 13 2
4 9 14 13 2
11 13 4 1 9 7 13 4 1 13 9 2
3 2 13 2
6 13 9 14 3 9 2
23 16 1 9 14 13 9 1 0 0 9 2 9 13 13 9 2 9 0 1 13 9 0 2
7 2 13 9 1 13 9 2
11 13 9 1 9 9 7 0 9 1 13 2
10 0 9 0 13 15 1 9 0 9 2
9 1 0 0 9 9 14 13 15 2
24 13 9 1 0 9 2 13 9 1 9 1 9 2 13 9 1 9 7 13 1 9 9 9 2
12 9 13 9 15 12 9 1 9 9 1 9 2
20 1 9 1 13 9 9 2 9 1 9 0 9 13 1 9 2 0 4 13 2
7 9 0 13 1 0 9 2
15 9 13 0 2 0 9 2 0 9 0 3 13 1 9 2
9 1 0 9 1 9 13 14 9 2
10 2 13 15 13 7 13 1 0 9 2
22 1 9 14 13 14 0 9 2 16 9 12 2 12 7 12 1 9 13 1 9 9 2
4 14 13 15 2
7 0 9 14 13 0 9 2
11 9 9 13 2 16 14 13 9 1 9 2
11 4 4 13 1 9 2 14 13 0 9 2
6 14 13 9 0 9 2
15 9 0 9 13 13 1 0 9 2 16 9 13 9 0 2
5 13 13 12 9 2
18 3 0 9 13 15 3 13 7 13 2 16 3 13 13 9 1 0 2
12 9 9 13 1 9 9 13 1 9 0 9 2
17 1 16 9 13 9 1 0 2 1 9 9 13 13 15 12 9 2
19 13 1 15 12 9 0 2 12 13 1 15 9 7 12 9 7 9 9 2
13 9 9 0 1 9 9 9 9 13 0 9 0 2
7 2 7 13 14 0 9 2
4 2 14 13 2
8 2 7 13 1 9 1 9 2
8 13 4 15 14 9 1 9 2
9 2 7 14 13 1 9 1 9 2
10 1 9 13 9 7 3 14 13 0 2
7 2 16 13 4 1 9 2
6 3 13 1 0 9 2
11 13 15 15 3 2 7 3 13 15 9 2
14 7 3 14 13 2 16 4 13 15 0 7 13 9 2
13 2 13 15 3 2 16 13 1 15 1 0 9 2
10 1 9 13 13 2 9 13 9 9 2
11 14 13 15 2 16 9 9 13 13 9 2
14 0 9 13 2 16 1 9 14 13 9 1 0 9 2
7 3 9 3 3 3 13 2
10 9 13 14 1 9 1 9 1 9 2
6 14 0 9 13 0 2
10 9 9 3 13 0 7 0 9 0 2
5 1 9 15 13 2
16 13 15 2 16 9 13 15 1 9 2 16 15 13 2 2 2
8 9 13 15 1 0 2 2 2
15 1 0 9 2 13 15 15 13 1 15 0 9 1 9 2
16 1 0 9 9 13 0 9 1 9 2 0 3 4 13 3 2
15 9 9 2 9 2 0 9 2 9 9 4 13 7 13 2
16 9 7 9 0 13 9 2 1 0 9 0 1 9 13 9 2
7 1 9 13 15 9 9 2
12 13 15 14 13 9 9 2 0 13 15 13 2
19 9 9 13 9 0 9 2 0 13 13 9 9 9 1 13 9 1 9 2
13 7 0 9 13 9 1 9 13 9 1 9 9 2
5 9 14 13 9 2
6 9 14 13 9 9 2
19 0 13 9 9 1 9 0 2 1 0 9 12 9 4 13 13 0 9 2
4 7 13 3 2
10 1 0 9 9 13 4 0 9 9 2
6 14 9 9 13 9 2
17 9 14 13 2 16 3 4 15 13 9 2 14 13 1 9 9 2
9 3 1 9 13 15 9 1 9 2
8 2 1 9 13 4 12 9 2
5 2 9 13 0 2
15 7 13 3 2 16 0 9 14 13 9 13 1 0 9 2
14 0 9 14 13 2 14 13 2 14 13 13 1 9 2
8 13 9 9 2 13 1 9 2
14 9 0 13 9 9 9 2 0 13 15 13 9 9 2
11 1 9 3 13 15 9 1 9 1 9 2
12 7 14 3 4 13 13 13 0 0 9 9 2
12 7 13 4 2 3 13 1 15 9 1 9 2
7 14 13 0 9 0 9 2
16 3 13 4 9 9 2 0 1 9 0 13 15 1 0 9 2
12 9 14 13 0 9 1 9 7 9 1 9 2
8 13 15 2 16 9 13 13 2
13 7 13 15 1 0 9 2 1 0 15 14 13 2
9 13 9 2 16 1 9 13 9 2
11 9 0 3 13 1 9 13 1 0 9 2
16 9 14 13 15 1 9 9 2 16 13 1 9 0 0 9 2
23 3 3 1 0 9 2 14 1 9 0 13 0 0 9 2 16 9 15 13 13 14 0 2
3 3 13 2
13 3 13 1 9 1 9 7 0 13 1 15 9 2
19 9 0 13 2 16 15 9 0 13 0 1 9 0 2 7 14 9 0 2
21 1 9 2 9 9 13 14 13 1 3 0 9 2 7 9 1 15 4 3 13 2
14 2 14 3 0 3 9 0 14 13 13 1 9 9 2
13 0 13 9 9 13 4 1 13 9 1 9 9 2
4 9 14 13 2
8 13 15 9 1 9 0 9 2
19 1 12 0 0 9 13 3 2 0 13 15 1 9 0 2 13 12 9 2
10 0 9 9 4 14 13 1 0 9 2
11 0 0 9 0 9 13 4 1 0 9 2
21 0 9 9 3 13 0 9 13 2 3 0 9 13 14 3 13 9 9 7 9 2
16 13 1 0 9 1 9 0 2 13 1 13 3 0 9 9 2
10 1 9 0 13 14 7 13 0 9 2
21 15 0 9 0 13 2 16 1 9 9 0 14 13 15 0 9 1 0 9 0 2
17 13 14 0 1 9 0 2 0 13 0 9 13 1 9 0 9 2
19 1 9 13 15 2 16 9 0 14 13 0 9 2 7 13 14 13 9 2
8 13 1 0 9 9 15 9 2
7 1 12 9 9 13 9 2
6 13 0 9 1 9 2
8 1 9 1 9 9 14 13 2
8 13 15 0 9 0 9 9 2
13 9 13 0 9 1 9 13 9 9 13 1 9 2
6 9 14 13 1 9 2
9 13 9 1 9 9 13 1 9 2
9 9 0 13 14 9 9 0 9 2
12 9 9 9 1 9 9 7 9 0 13 0 2
11 13 9 1 9 9 9 14 13 0 9 2
13 16 3 13 2 1 9 9 3 13 14 15 9 2
7 3 9 0 14 13 0 2
21 9 1 9 9 7 9 13 15 3 13 14 0 9 9 2 7 7 9 7 9 2
16 9 9 13 1 9 0 1 0 9 9 0 3 3 13 9 2
11 0 0 9 13 14 1 0 9 0 9 2
27 0 2 0 9 2 0 9 7 9 9 13 2 16 13 1 0 9 1 9 9 3 14 4 13 1 9 2
15 1 9 9 13 14 0 9 1 9 0 2 0 13 0 2
12 13 8 1 9 7 13 9 1 9 2 2 2
14 13 13 9 2 0 3 4 13 2 13 9 0 9 2
16 16 13 1 9 9 7 9 9 0 2 9 13 15 3 0 2
7 9 9 13 1 9 9 2
16 0 9 0 9 7 0 9 0 9 9 0 13 15 14 13 2
11 14 13 14 2 1 12 0 13 13 9 2
12 14 1 0 9 9 9 0 9 9 13 0 2
11 14 3 0 0 9 13 9 0 1 9 2
16 14 0 9 9 9 0 13 9 0 7 13 9 0 9 0 2
8 9 9 13 0 9 1 0 2
11 1 9 1 15 13 0 9 13 9 9 2
6 1 9 9 13 3 2
11 9 9 1 9 0 9 9 13 13 9 2
15 9 1 9 1 0 9 9 13 9 9 13 1 9 9 2
15 9 2 13 1 9 1 9 2 13 15 0 1 9 9 2
9 12 9 0 9 13 9 1 0 2
2 13 2
11 9 0 13 9 1 0 9 7 13 9 2
6 13 9 2 13 13 2
5 13 14 9 9 2
9 3 9 0 2 0 13 15 13 2
7 13 9 13 7 13 9 2
7 9 9 13 15 1 9 2
7 1 0 9 13 13 9 2
12 13 1 0 9 9 14 13 1 9 1 9 2
6 13 1 0 9 9 2
10 14 9 9 9 3 4 13 1 9 2
21 1 9 0 9 1 9 1 0 13 15 1 15 9 9 13 9 9 1 9 9 2
8 13 0 7 13 9 0 13 2
12 13 15 9 2 16 0 9 13 15 9 9 2
5 9 13 1 9 2
6 9 9 13 14 9 2
12 9 9 1 8 2 9 13 1 15 0 9 2
10 0 9 9 9 13 0 9 0 9 2
12 9 13 1 9 1 0 9 12 8 2 8 2
4 2 3 13 2
7 0 9 13 1 15 9 2
10 14 9 13 1 15 9 1 9 0 2
10 14 9 0 13 1 15 1 13 9 2
10 14 12 9 9 7 9 13 1 9 2
8 1 0 9 13 14 12 9 2
8 9 3 13 9 13 15 9 2
15 9 13 0 9 2 16 1 9 13 15 9 9 1 9 2
13 9 13 1 15 0 9 7 1 9 3 15 13 2
16 3 0 9 1 9 2 13 7 13 1 9 2 9 13 9 2
14 13 4 2 16 13 0 9 2 1 9 13 9 9 2
10 14 9 13 1 0 9 1 0 9 2
4 9 13 9 2
8 13 15 15 9 9 1 9 2
17 0 9 13 1 9 9 2 9 2 9 1 9 9 7 0 9 2
9 9 13 3 9 1 3 12 9 2
17 1 9 9 0 9 1 9 1 13 9 13 2 16 4 15 13 2
8 9 1 12 9 13 1 9 2
17 0 9 2 13 3 1 0 9 1 9 1 9 2 13 9 9 2
16 0 9 9 9 13 9 2 16 9 7 9 13 3 13 9 2
7 13 15 15 3 3 3 2
7 1 0 9 13 3 3 2
9 3 13 9 13 1 9 0 9 2
11 16 9 13 1 9 9 2 9 14 13 2
10 13 14 13 2 16 13 9 0 9 2
14 9 1 0 9 13 2 16 13 1 15 9 1 9 2
9 9 7 0 9 13 1 0 9 2
5 2 13 0 9 2
4 4 14 13 2
17 13 15 9 2 9 13 2 9 13 1 9 2 13 9 7 13 2
9 14 13 9 2 13 4 1 9 2
4 14 13 9 2
5 14 9 15 13 2
14 9 14 13 2 7 3 13 15 15 9 1 15 9 2
7 12 9 13 1 9 9 2
2 13 2
2 13 2
3 13 15 2
10 9 13 9 9 3 2 1 0 9 2
8 13 7 9 2 0 3 13 2
9 14 9 14 13 0 9 2 2 2
6 13 15 0 0 9 2
5 3 14 13 9 2
13 3 13 0 0 9 7 3 13 0 9 0 9 2
7 13 15 1 12 0 9 2
7 0 9 13 15 14 0 2
7 9 13 9 1 0 9 2
10 9 1 0 9 13 14 3 0 9 2
3 13 4 2
9 14 15 1 9 13 0 9 9 2
4 7 3 13 2
7 14 15 13 9 7 9 2
9 3 13 4 1 9 9 7 9 2
10 0 9 13 4 1 0 2 13 9 2
16 14 13 4 1 9 13 0 0 9 2 13 1 9 0 9 2
9 14 1 9 13 2 9 9 13 2
7 7 3 13 4 15 9 2
9 13 15 0 9 2 9 13 15 2
7 7 3 13 13 1 15 2
9 13 0 9 7 13 1 9 3 2
3 13 13 2
6 7 7 13 7 13 2
4 13 4 15 2
7 13 9 7 0 9 9 2
4 9 13 9 2
14 9 3 13 15 9 0 9 2 0 3 13 15 9 2
6 1 13 9 13 9 2
5 3 13 9 9 2
15 14 1 12 9 13 15 13 1 13 9 7 0 9 9 2
10 14 13 9 0 9 2 14 13 9 2
6 1 0 9 13 3 2
22 13 0 2 13 9 7 13 9 2 7 9 9 2 9 2 9 7 9 13 9 9 2
4 13 9 9 2
8 9 13 1 9 12 9 9 2
4 14 13 9 2
4 9 15 13 2
7 9 0 13 9 1 9 2
22 9 13 9 2 16 1 9 0 9 9 9 13 1 13 0 9 1 0 0 9 0 2
19 0 13 2 16 9 9 0 4 13 1 9 9 13 9 1 0 9 9 2
22 13 1 9 2 16 9 1 0 9 13 13 9 1 9 0 9 2 9 0 7 0 2
13 1 9 7 9 13 15 0 9 1 3 0 9 2
7 13 15 9 4 14 0 2
6 13 13 0 9 0 2
6 13 0 7 13 9 2
5 13 7 13 3 2
3 13 4 2
11 13 0 9 1 0 7 13 15 1 9 2
5 2 9 14 13 2
6 7 3 15 3 13 2
13 9 14 13 1 0 9 9 1 9 2 13 0 2
11 1 0 9 0 13 15 9 1 0 9 2
8 9 14 13 3 9 1 9 2
15 9 1 9 13 2 16 9 13 14 13 9 14 1 9 2
9 1 9 9 3 13 1 9 9 2
10 4 15 1 15 13 2 1 12 9 2
5 3 1 9 13 2
5 2 13 1 9 2
7 7 3 9 9 3 13 2
7 2 7 13 2 13 9 2
6 13 2 13 2 2 2
4 13 13 9 2
6 13 7 13 1 9 2
13 13 1 9 7 13 2 13 15 1 9 9 9 2
4 13 15 9 2
9 13 14 1 9 1 9 1 9 2
7 13 9 2 13 0 9 2
13 2 13 4 0 9 2 13 2 16 13 2 2 2
3 2 13 2
4 2 3 13 2
4 3 15 13 2
7 2 13 0 9 2 9 2
14 9 0 13 1 12 9 7 13 0 9 1 9 0 2
21 0 9 9 2 13 1 13 0 9 2 13 13 9 1 9 9 1 9 9 0 2
4 9 13 9 2
18 9 9 1 0 9 13 9 7 15 9 2 0 13 1 9 1 9 2
10 13 9 13 7 3 13 1 9 0 2
8 1 9 9 13 9 9 0 2
11 16 1 9 9 14 13 2 9 13 9 2
18 9 2 1 13 2 14 13 3 1 9 2 7 1 9 13 15 9 2
22 15 9 9 0 13 15 1 9 1 8 2 0 2 1 0 3 1 9 13 15 9 2
15 3 9 13 9 9 9 1 9 2 3 13 0 9 9 2
14 13 9 1 9 9 9 9 1 9 1 8 2 0 2
12 9 13 3 9 2 1 0 9 13 0 9 2
11 14 4 13 9 0 2 13 13 14 9 2
15 1 0 9 3 13 4 15 7 3 9 13 15 0 9 2
13 13 4 1 0 9 9 14 12 9 1 0 9 2
19 13 4 9 9 2 16 13 15 9 7 1 0 13 3 13 15 1 9 2
5 13 1 9 9 2
6 13 2 0 9 13 2
9 13 15 1 9 9 1 0 9 2
5 14 13 0 9 2
6 2 13 1 15 9 2
13 2 14 13 15 1 9 0 1 0 9 9 9 2
11 1 9 0 1 9 9 13 15 12 9 2
21 16 0 9 13 9 7 9 2 7 9 13 0 2 13 13 15 1 3 13 9 2
14 13 0 1 0 0 9 2 0 13 3 0 0 9 2
11 1 9 13 9 2 7 9 13 15 9 2
14 13 2 16 3 13 9 0 9 2 7 13 15 15 2
8 13 15 9 2 3 13 9 2
5 3 13 15 9 2
15 2 14 13 0 9 2 14 14 13 4 9 1 15 13 2
11 1 9 13 15 9 2 0 13 13 9 2
9 14 2 3 9 9 14 13 9 2
13 1 9 1 0 12 9 13 9 0 9 7 9 2
6 1 12 9 4 13 2
16 1 9 2 1 9 0 9 0 2 13 15 13 9 0 9 2
19 9 7 9 13 2 16 13 1 9 2 16 13 1 9 13 1 9 9 2
6 1 9 14 13 9 2
7 15 1 9 13 9 0 2
20 0 9 14 13 13 0 9 9 0 1 9 9 2 7 9 0 13 9 9 2
12 3 9 3 13 2 16 13 0 9 1 9 2
11 9 13 15 1 0 9 1 0 9 0 2
13 9 13 15 1 12 9 9 0 9 1 9 0 2
9 9 12 1 12 13 9 13 0 2
13 13 1 13 14 12 9 7 12 9 1 0 9 2
5 12 9 13 9 2
14 13 15 0 9 1 9 9 7 13 15 13 1 9 2
22 3 13 15 13 15 1 9 2 16 1 9 13 1 13 1 9 9 9 13 15 3 2
11 9 14 13 15 1 0 9 13 7 9 2
13 14 12 9 4 13 1 9 1 9 1 9 9 2
6 13 9 1 0 9 2
12 0 9 0 9 13 9 1 9 9 2 9 2
14 1 9 0 9 1 9 0 9 0 13 13 9 13 2
10 9 0 9 13 1 9 0 9 0 2
12 15 13 1 9 9 2 0 13 9 13 9 2
6 2 13 1 9 9 2
8 2 4 9 13 1 9 9 2
10 2 14 4 9 14 3 13 1 9 2
10 1 9 13 9 7 3 13 13 9 2
7 9 13 15 7 13 9 2
11 13 14 13 3 1 9 2 13 1 9 2
12 0 9 13 1 9 7 13 9 1 0 9 2
11 0 9 13 1 9 2 9 7 13 9 2
7 9 13 15 1 9 9 2
13 1 9 13 15 12 9 2 14 13 12 9 0 2
10 1 9 9 7 9 14 13 12 9 2
8 1 9 9 0 13 9 9 2
8 1 0 9 13 15 2 9 2
8 1 9 9 13 15 2 9 2
8 0 9 13 13 1 9 9 2
9 9 13 9 7 9 13 9 0 2
8 2 13 1 9 13 15 3 2
7 2 9 13 9 2 2 2
11 0 9 13 2 16 9 9 13 0 9 2
10 13 15 9 2 13 15 9 0 9 2
8 1 0 9 13 15 2 9 2
10 1 9 0 7 9 13 15 2 9 2
15 16 9 13 15 13 13 9 1 9 2 13 14 0 9 2
6 9 13 1 15 3 2
13 13 13 3 1 9 2 1 9 13 1 9 9 2
5 9 13 0 9 2
8 9 13 15 13 9 1 9 2
18 13 1 9 2 16 0 9 13 15 1 9 2 13 9 1 9 9 2
13 9 2 0 0 9 2 13 9 1 9 9 0 2
10 9 0 13 0 9 0 13 1 9 2
12 9 13 12 9 1 13 9 7 13 9 9 2
21 0 9 9 13 9 1 9 2 0 14 1 9 0 9 13 9 1 0 9 0 2
19 0 9 13 15 1 9 9 0 7 0 7 13 9 1 9 9 1 9 2
15 0 1 13 9 13 15 1 9 9 0 7 0 1 9 2
12 13 15 13 15 1 9 13 1 9 1 9 2
16 1 9 9 13 14 3 12 9 2 13 1 13 1 9 9 2
6 0 15 14 13 4 2
15 13 15 12 2 16 1 9 9 13 4 15 1 13 9 2
16 1 9 9 2 9 9 0 9 0 2 13 4 1 0 9 2
14 1 9 13 4 0 9 9 1 9 0 0 9 0 2
9 13 15 2 16 3 1 15 13 2
18 1 9 9 9 1 9 2 9 2 9 7 9 13 9 1 13 9 2
11 9 1 9 9 0 13 9 9 1 9 2
8 9 13 9 1 9 12 8 2
23 3 1 12 0 9 1 9 13 15 9 0 1 9 9 0 1 9 1 9 1 9 9 2
7 9 9 9 13 9 9 2
7 13 15 1 9 9 9 2
9 1 9 9 13 14 0 9 9 2
12 0 9 9 9 0 13 15 1 9 1 9 2
10 13 2 16 0 9 13 14 9 9 2
9 1 0 9 9 9 13 12 9 2
9 2 13 2 16 9 14 13 9 2
7 13 15 1 9 9 9 2
12 0 9 9 9 0 13 15 1 9 1 9 2
12 13 0 9 13 9 9 9 7 9 1 9 2
7 13 1 15 0 9 0 2
8 1 0 9 14 13 9 9 2
10 12 9 13 9 8 2 9 1 9 2
13 1 12 9 13 4 9 13 1 9 9 1 9 2
12 1 0 0 9 13 12 9 13 1 12 9 2
18 1 9 0 13 9 0 1 0 7 13 9 2 0 13 9 9 9 2
13 1 9 13 9 9 0 2 7 9 13 1 9 2
6 9 9 13 1 9 2
7 9 13 1 15 0 9 2
20 0 9 1 0 9 13 15 14 9 2 0 13 12 1 12 13 1 9 9 2
13 0 9 9 13 15 1 9 0 9 1 0 9 2
9 1 9 1 9 13 0 9 9 2
9 1 9 13 4 3 13 9 9 2
9 1 9 0 13 9 1 9 0 2
10 1 9 13 14 0 9 7 9 9 2
19 1 0 9 9 9 0 1 9 4 13 9 1 9 1 9 1 12 9 2
17 3 9 9 2 1 0 13 4 9 2 13 1 9 1 12 9 2
4 9 13 9 2
16 1 9 7 9 13 9 0 9 2 9 0 1 0 9 0 2
16 1 15 9 13 2 16 3 1 9 0 13 9 1 9 9 2
5 9 13 1 9 2
13 1 9 7 9 13 15 9 7 9 7 9 0 2
17 13 15 2 16 3 0 15 13 14 12 9 9 9 1 9 0 2
3 3 13 2
15 9 13 1 9 1 9 2 13 12 9 9 7 9 9 2
13 9 13 2 3 13 7 13 1 0 9 1 9 2
13 1 0 9 13 9 1 9 7 13 15 3 9 2
20 9 7 9 13 2 13 1 9 7 12 9 9 1 0 9 7 13 1 9 2
13 14 1 0 9 13 9 1 9 1 9 7 9 2
14 12 9 1 9 9 13 9 1 9 1 9 1 9 2
5 14 13 14 9 2
22 13 9 2 9 13 2 16 9 0 3 15 14 13 2 7 1 9 13 12 9 0 2
22 9 13 14 2 16 13 9 9 1 9 9 9 7 0 9 9 7 0 9 1 15 2
6 4 13 1 9 9 2
7 9 1 3 14 13 0 2
4 13 3 0 2
8 0 0 13 15 15 13 0 2
12 1 0 9 0 9 13 15 1 0 9 13 2
13 13 13 2 16 3 13 9 1 9 1 0 9 2
11 3 13 1 0 9 2 13 15 7 13 2
10 3 13 1 9 2 13 9 2 13 2
7 13 15 1 9 9 9 2
6 3 3 13 15 13 2
9 9 3 13 2 13 9 12 9 2
6 2 13 4 0 9 2
4 9 13 9 2
3 9 13 2
6 3 13 4 15 9 2
11 2 14 13 15 9 2 16 14 13 9 2
6 2 14 13 1 15 2
6 2 13 4 1 9 2
5 2 15 15 13 2
5 2 9 15 13 2
6 13 14 4 15 13 2
4 3 15 13 2
3 9 13 2
7 7 1 9 13 1 15 2
13 9 4 13 2 3 3 13 9 2 13 0 9 2
20 9 9 13 1 9 1 0 9 0 9 2 16 13 15 9 1 12 8 8 2
15 9 13 2 16 9 3 13 9 13 1 9 9 9 9 2
8 13 9 9 1 9 1 9 2
5 3 15 9 13 2
11 13 4 1 0 9 7 13 4 15 9 2
11 1 9 2 13 15 1 15 1 9 0 2
16 12 9 1 0 9 13 3 1 9 2 9 2 14 1 9 2
12 14 13 9 2 16 0 9 14 15 14 13 2
20 13 7 1 9 2 16 9 2 1 9 9 2 13 1 9 13 9 1 9 2
21 1 0 9 0 9 13 1 9 9 13 15 3 2 13 15 1 9 1 9 9 2
5 9 14 13 9 2
15 2 9 2 13 15 2 0 13 1 9 9 13 3 9 2
20 13 15 0 9 0 2 13 1 0 9 9 0 7 9 1 9 9 7 9 2
9 9 9 13 13 9 0 1 9 2
16 13 15 2 16 13 9 0 3 4 13 13 1 9 1 9 2
5 3 13 1 9 2
5 13 3 1 15 2
5 13 2 9 13 2
6 13 15 9 1 9 2
11 9 13 15 9 2 13 4 15 1 9 2
5 7 3 13 4 2
3 13 13 2
10 9 3 13 0 9 1 9 1 9 2
4 13 1 9 2
15 13 14 0 9 2 0 9 4 13 1 9 1 15 9 2
22 13 16 9 9 1 9 7 9 2 1 15 13 13 9 9 7 13 9 0 9 9 2
14 9 0 13 12 9 2 16 13 1 15 9 1 9 2
9 13 9 9 0 9 1 0 9 2
15 1 9 0 4 13 1 9 9 9 9 0 9 9 9 2
6 9 1 15 13 0 2
15 13 1 9 13 9 7 13 1 9 2 13 13 9 9 2
9 9 1 15 13 1 9 1 9 2
11 1 0 9 13 1 9 9 9 1 9 2
14 13 14 1 0 9 2 0 13 14 13 1 13 9 2
8 9 13 1 0 9 0 9 2
14 9 13 1 9 9 2 16 1 0 9 13 0 9 2
15 3 13 4 9 1 9 13 2 0 13 15 1 9 9 2
8 9 13 0 9 2 1 9 2
8 1 9 13 1 14 13 9 2
7 1 9 9 14 13 9 2
19 9 9 2 0 13 0 9 8 2 2 14 13 15 1 9 7 13 9 2
10 1 9 13 1 9 1 9 0 9 2
4 9 13 0 2
11 9 1 13 9 7 9 9 13 1 9 2
10 9 3 2 1 9 2 13 1 9 2
11 9 9 9 13 0 9 14 1 0 9 2
14 13 14 0 0 9 1 0 9 1 9 0 9 9 2
8 9 13 1 0 9 9 9 2
11 1 0 9 13 15 15 1 0 9 0 2
10 3 13 15 0 9 1 0 9 0 2
5 13 4 13 9 2
7 9 13 15 1 13 9 2
22 0 13 15 13 1 9 2 1 16 9 13 15 14 1 9 7 13 9 13 3 0 2
7 12 9 13 0 2 2 2
9 9 1 12 0 9 13 1 9 2
14 9 4 3 13 2 7 9 9 13 1 9 9 0 2
10 1 9 13 1 9 1 9 1 9 2
8 9 13 15 9 1 12 9 2
24 1 9 12 9 13 1 9 0 7 9 9 9 0 2 3 1 12 9 9 13 9 9 0 2
9 9 13 0 7 13 12 9 9 2
9 0 9 13 4 1 3 13 9 2
12 13 0 9 9 0 2 1 0 13 0 9 2
8 0 9 13 1 9 0 9 2
5 4 15 3 13 2
23 16 9 9 13 9 2 9 9 13 1 8 2 9 9 13 15 1 9 9 7 9 9 2
11 1 9 9 9 13 15 1 9 0 9 2
8 13 0 2 0 9 1 9 2
8 2 4 13 2 13 0 9 2
11 9 9 13 1 12 0 9 1 0 9 2
19 2 9 13 2 16 13 9 9 1 9 7 3 9 13 3 1 0 9 2
14 13 4 9 1 9 1 9 0 2 3 13 4 9 2
13 9 13 1 9 0 2 16 3 13 0 9 9 2
15 1 0 9 14 13 4 2 16 9 0 1 9 15 13 2
13 13 14 0 9 2 0 1 9 9 7 9 9 2
10 1 0 9 13 0 9 13 0 9 2
10 13 1 9 12 13 1 0 9 9 2
20 9 0 13 1 9 12 9 15 13 2 16 13 1 9 2 14 0 7 0 2
15 9 9 9 13 1 9 13 0 9 1 13 3 0 9 2
25 9 9 9 9 13 2 16 4 13 0 2 13 1 9 9 9 2 0 3 13 9 9 1 9 2
28 9 9 9 9 13 0 9 0 9 2 0 13 15 1 13 9 7 1 0 9 1 9 4 13 13 1 9 2
10 2 9 13 15 1 0 2 0 9 2
13 2 9 13 2 16 1 3 0 9 13 1 9 2
20 1 0 9 13 9 7 9 2 3 3 13 15 7 13 3 9 0 2 0 2
13 14 14 13 1 0 9 14 9 9 9 9 9 2
13 12 14 13 0 9 1 9 13 9 1 9 0 2
8 7 3 13 14 3 2 2 2
9 7 3 15 0 9 13 2 2 2
12 1 9 13 15 13 2 16 9 13 1 9 2
10 2 13 13 2 9 2 9 14 13 2
9 9 13 15 9 7 13 1 0 2
15 13 1 9 2 1 0 13 15 0 9 2 13 1 9 2
9 9 13 15 7 13 1 12 9 2
5 2 14 13 9 2
6 9 15 1 9 13 2
5 13 15 1 9 2
9 3 3 9 13 2 16 13 13 2
14 9 13 2 16 1 9 9 9 13 9 9 0 9 2
17 9 9 0 9 9 9 9 13 1 9 0 9 9 7 9 9 2
8 3 9 13 9 13 1 9 2
24 9 9 9 1 9 13 15 9 13 1 9 0 9 2 16 13 9 9 1 15 9 13 9 2
12 3 14 13 4 2 16 1 0 9 13 9 2
12 15 13 2 16 13 4 9 7 9 15 13 2
8 13 4 1 0 2 0 9 2
6 0 4 13 3 9 2
4 13 15 15 2
7 13 0 0 9 1 9 2
26 13 14 2 16 1 12 9 13 15 9 1 9 2 0 1 9 0 0 9 13 13 9 9 1 9 2
12 12 0 9 13 9 1 9 2 9 2 9 2
13 13 2 16 13 13 9 1 9 1 9 1 9 2
9 13 14 9 1 9 2 13 9 2
23 3 2 1 9 9 9 2 0 13 1 9 9 13 1 0 9 7 13 1 15 0 9 2
8 9 1 0 9 13 0 9 2
11 1 0 9 9 1 13 9 13 12 9 2
6 0 9 13 15 0 2
8 1 9 0 0 9 13 9 2
5 9 1 15 13 2
6 3 9 0 13 13 2
10 13 15 9 9 7 13 9 9 0 2
20 13 1 9 13 15 1 13 9 2 16 13 0 9 7 9 0 1 9 13 2
6 9 14 13 15 9 2
4 13 9 13 2
5 15 14 14 13 2
5 3 13 1 9 2
13 0 9 13 1 9 9 2 16 13 4 1 9 2
8 14 13 1 9 0 9 9 2
16 13 4 1 0 0 0 9 2 1 0 13 15 3 3 13 2
7 3 13 9 9 1 9 2
4 13 7 13 2
14 9 1 9 13 9 9 2 13 4 2 3 13 9 2
6 16 13 9 1 9 2
12 13 15 9 3 1 3 13 2 0 9 0 2
11 13 13 2 16 9 0 13 0 9 9 2
10 1 9 3 13 13 0 9 9 9 2
10 3 9 13 1 9 9 1 0 9 2
7 0 9 14 13 1 9 2
5 13 13 9 0 2
6 9 13 1 9 0 2
16 9 1 9 9 9 13 15 2 16 3 3 14 13 0 9 2
7 9 9 13 13 13 9 2
15 13 15 13 9 0 2 0 13 15 13 9 0 9 9 2
10 9 4 14 13 13 1 9 9 9 2
8 9 0 9 13 9 0 9 2
19 1 9 9 0 9 13 15 13 1 9 1 9 9 9 0 13 1 9 2
17 1 15 9 9 13 1 15 7 13 2 16 13 4 3 0 9 2
4 14 13 15 2
12 13 4 15 1 9 0 7 13 1 0 9 2
7 13 15 2 16 13 3 2
7 13 15 3 13 1 9 2
17 9 9 13 0 9 2 0 13 13 1 9 2 1 0 9 13 2
6 13 14 13 1 9 2
8 1 9 13 13 9 7 9 2
22 13 9 2 0 13 13 9 2 7 1 9 1 9 4 13 1 12 9 13 1 9 2
14 9 2 14 1 9 0 9 2 13 13 3 13 9 2
13 2 0 9 9 0 1 9 13 15 1 12 8 2
9 15 1 12 8 2 4 13 3 2
9 2 3 9 13 1 9 9 9 2
14 3 9 9 0 13 9 9 2 13 15 9 1 9 2
11 2 1 0 9 13 9 13 13 0 9 2
6 2 3 13 3 3 2
4 3 13 3 2
10 2 14 9 3 15 13 1 9 9 2
6 13 3 2 13 9 2
5 3 13 0 9 2
12 9 13 9 1 9 9 7 9 1 9 9 2
17 13 3 13 2 16 1 12 9 0 13 9 9 12 13 9 9 2
6 14 3 15 13 4 2
17 13 9 1 9 2 9 13 15 1 9 2 7 14 13 15 9 2
15 13 4 0 7 0 9 2 13 15 9 13 1 9 9 2
13 7 14 13 9 2 14 14 13 14 3 2 2 2
7 14 13 15 13 2 2 2
14 9 9 13 1 9 2 0 9 0 14 13 9 9 2
16 9 0 9 13 14 15 1 0 9 2 0 9 4 14 13 2
12 1 0 9 0 9 9 9 9 13 0 9 2
13 14 0 9 14 13 14 1 9 0 9 1 9 2
10 9 14 13 15 2 9 13 1 9 2
9 0 9 1 13 9 13 9 9 2
9 13 9 2 16 13 0 13 13 2
24 0 9 9 13 1 9 1 9 13 9 2 7 13 13 2 16 13 4 15 1 9 9 9 2
11 13 9 13 0 9 0 9 1 0 9 2
11 13 15 1 0 9 9 13 1 9 9 2
12 13 9 0 2 16 1 0 9 13 12 9 2
15 0 1 15 13 9 9 2 0 13 1 13 9 0 9 2
15 9 0 13 15 1 13 1 15 9 1 0 9 7 9 2
9 9 0 13 15 1 0 9 9 2
18 9 2 0 15 13 2 3 13 12 9 13 1 0 2 13 14 9 2
11 1 0 9 9 13 13 9 1 0 9 2
20 9 13 1 9 1 0 9 0 9 3 0 2 13 9 0 7 13 0 9 2
10 1 0 9 13 15 14 1 9 9 2
5 3 13 9 9 2
10 9 13 15 1 9 7 13 1 9 2
13 9 13 15 3 3 7 13 14 9 1 0 9 2
7 3 13 9 13 1 9 2
7 13 13 15 13 0 9 2
4 3 13 9 2
10 9 0 13 9 1 9 9 9 0 2
12 9 1 9 0 4 13 1 9 1 9 9 2
9 0 9 13 9 1 9 1 9 2
17 9 13 2 16 15 13 13 1 9 9 2 7 9 14 13 9 2
12 9 9 9 1 9 14 13 9 1 15 9 2
23 0 9 9 13 15 1 0 9 0 9 2 16 9 13 0 9 7 9 13 1 0 9 2
10 9 13 1 0 9 9 1 0 9 2
17 14 13 2 3 13 15 0 9 2 13 2 16 13 14 15 3 2
5 2 13 0 9 2
7 13 3 1 15 2 2 2
9 13 15 1 9 7 13 1 9 2
3 13 9 2
8 2 13 2 14 13 15 13 2
7 14 15 9 14 14 13 2
6 0 9 9 3 13 2
6 2 3 13 13 9 2
17 2 3 14 13 4 2 14 13 2 16 1 0 9 13 14 13 2
13 2 14 13 9 13 1 9 2 14 15 15 13 2
5 14 13 1 9 2
7 9 14 13 15 0 9 2
3 2 13 2
11 9 9 9 1 9 13 1 9 9 0 2
11 1 0 14 9 13 14 12 8 2 9 2
16 1 9 13 1 9 2 9 7 9 13 12 8 2 0 9 2
11 9 9 2 9 9 0 2 13 0 9 2
11 14 14 9 9 13 9 9 2 2 2 2
6 13 14 9 9 9 2
11 9 14 13 0 2 14 13 9 2 2 2
5 2 3 9 13 2
14 9 0 13 13 12 9 2 12 13 9 0 1 9 2
6 1 9 14 3 13 2
18 14 13 4 15 15 13 2 7 15 13 2 16 13 1 9 2 2 2
15 1 0 9 13 15 9 0 2 0 9 9 7 9 9 2
5 9 9 13 9 2
6 1 9 13 9 9 2
22 9 9 2 14 13 13 0 2 0 9 7 0 9 9 2 13 15 7 13 1 9 2
17 1 9 9 9 13 0 9 1 9 2 9 13 1 9 9 9 2
9 9 13 7 9 13 15 15 9 2
18 13 3 2 1 9 2 1 9 13 9 1 0 9 2 13 15 3 2
16 13 15 2 13 14 1 9 9 13 1 9 7 13 1 9 2
14 9 7 9 13 15 2 9 1 9 1 9 4 13 2
7 1 9 1 9 14 13 2
14 13 9 9 9 1 9 2 13 9 7 13 1 9 2
8 13 9 2 13 9 2 13 2
5 9 14 14 13 2
19 1 0 9 13 15 0 2 0 9 9 9 2 13 1 9 13 1 9 2
20 9 9 13 15 1 9 2 13 1 9 2 13 0 9 2 9 13 1 9 2
10 13 15 1 9 1 9 9 9 9 2
7 13 15 13 1 13 9 2
8 3 9 13 9 13 1 9 2
11 9 9 9 9 13 0 9 7 13 9 2
7 14 13 15 15 13 9 2
7 13 9 9 1 9 9 2
10 7 9 13 0 9 8 2 1 9 2
6 8 2 13 13 9 2
7 3 13 13 15 1 9 2
9 13 15 13 2 9 13 4 9 2
9 1 9 13 15 9 0 0 9 2
10 0 9 9 4 13 1 9 0 9 2
13 3 9 13 1 9 2 13 15 1 9 1 9 2
7 9 14 15 1 15 13 2
20 0 9 2 0 7 0 2 3 3 13 15 1 9 2 13 1 9 9 0 2
17 1 9 9 1 9 1 9 9 13 1 9 2 3 13 15 9 2
8 15 0 9 13 9 7 9 2
21 1 0 0 9 1 9 13 4 2 1 9 9 1 9 0 2 9 1 9 9 2
11 1 9 13 4 13 9 0 9 2 2 2
16 13 4 15 1 0 9 7 13 4 15 1 0 9 1 9 2
11 9 13 1 9 9 13 1 0 0 9 2
9 1 0 9 13 4 15 1 9 2
7 3 13 1 15 0 9 2
16 16 9 3 15 13 2 9 14 14 13 0 9 2 0 13 2
12 14 3 13 9 2 13 3 3 0 0 9 2
18 9 13 2 16 1 0 9 14 4 9 2 13 9 9 14 0 9 2
19 9 2 9 13 1 0 9 9 0 7 9 3 13 9 13 1 9 9 2
10 1 9 9 9 13 9 1 9 0 2
5 7 13 13 9 2
6 2 9 3 13 4 2
12 13 4 9 1 9 7 13 4 9 1 15 2
8 7 13 1 9 9 9 0 2
13 16 9 13 2 14 14 0 2 13 4 13 9 2
9 13 7 7 15 2 7 14 9 2
6 14 13 4 9 13 2
5 9 14 9 13 2
13 3 3 2 3 13 1 9 2 13 9 1 9 2
14 14 13 15 13 2 16 13 1 9 9 13 0 9 2
10 3 13 2 16 1 9 13 15 13 2
9 0 9 9 13 9 0 9 0 2
7 3 13 15 14 9 9 2
9 3 13 7 9 13 9 1 9 2
6 3 3 13 9 9 2
10 3 13 15 9 2 9 2 0 9 2
18 2 14 13 15 15 1 0 9 2 7 13 13 2 1 9 15 13 2
10 13 2 16 9 13 14 1 15 0 2
8 13 15 2 16 13 9 9 2
6 1 9 3 13 9 2
7 3 13 13 9 1 9 2
13 9 1 9 2 9 2 13 1 3 0 9 0 2
14 13 14 2 16 9 13 1 9 9 0 9 7 9 2
8 14 9 13 9 1 0 9 2
4 13 15 9 2
10 7 14 0 9 9 13 15 9 0 2
6 0 0 9 13 9 2
7 9 13 9 9 1 9 2
13 13 2 13 0 9 1 9 9 9 9 1 9 2
12 0 9 13 0 9 9 13 9 9 1 9 2
15 1 0 9 9 0 13 15 1 9 7 13 13 9 0 2
12 1 13 15 1 9 13 15 1 9 1 9 2
5 13 9 9 9 2
14 9 9 2 9 0 2 13 9 0 0 9 1 9 2
8 13 1 13 9 9 1 9 2
6 2 13 13 1 9 2
5 13 4 2 2 2
8 13 4 14 0 9 2 13 2
5 9 2 13 9 2
12 13 2 15 13 13 9 0 1 9 1 15 2
3 2 13 2
4 2 14 13 2
5 3 13 15 9 2
5 14 13 9 9 2
10 2 9 13 2 16 0 13 12 9 2
6 13 15 9 9 9 2
7 2 9 2 0 4 13 2
5 2 9 13 15 2
5 2 13 15 9 2
4 9 13 9 2
6 2 13 15 1 9 2
6 13 15 3 1 9 2
3 13 15 2
3 14 13 2
12 9 14 13 15 3 2 9 13 13 1 15 2
5 9 13 15 0 2
3 2 13 2
6 7 3 13 15 3 2
5 9 9 13 9 2
7 9 4 13 1 9 3 2
4 9 14 13 2
19 1 14 12 9 1 9 0 1 13 9 14 13 9 1 13 1 0 9 2
5 13 13 9 9 2
9 15 15 14 13 9 9 7 9 2
6 7 13 15 9 9 2
9 16 9 13 9 2 4 15 13 2
18 3 1 15 2 9 0 9 13 1 9 9 1 9 9 9 9 9 2
13 1 12 13 1 9 13 1 9 12 9 1 9 2
10 1 12 9 13 4 9 1 9 9 2
12 13 4 9 1 9 1 9 9 13 9 0 2
11 3 3 14 13 4 2 16 13 4 9 2
5 2 14 13 15 2
4 2 14 13 2
3 13 9 2
13 13 15 1 9 0 2 9 13 15 9 13 9 2
7 13 9 1 3 0 9 2
5 15 13 0 13 2
18 14 1 12 9 9 9 9 0 13 0 7 0 2 7 9 14 13 2
17 16 16 13 9 2 14 13 9 0 13 15 9 1 9 7 9 2
12 1 9 1 9 8 2 13 1 15 0 9 2
9 2 0 13 1 15 9 1 9 2
14 13 9 1 9 9 2 13 9 9 13 15 9 9 2
14 1 9 1 9 13 12 9 2 1 9 12 1 9 2
13 2 13 4 9 2 13 9 9 1 9 2 2 2
19 13 3 9 9 2 9 9 2 9 9 2 3 1 15 9 13 9 9 2
9 2 14 0 9 0 3 13 9 2
14 2 13 9 2 3 1 12 9 9 13 1 9 9 2
8 2 13 13 1 0 0 9 2
7 4 0 9 13 0 9 2
8 2 13 0 9 1 13 9 2
18 1 0 9 13 15 2 14 1 0 0 9 4 13 15 13 9 0 2
9 14 13 9 2 16 13 1 9 2
12 9 0 9 13 0 9 0 9 9 1 9 2
7 9 13 0 9 9 9 2
9 1 0 9 9 13 0 9 9 2
5 13 2 9 9 2
2 13 2
6 2 13 14 1 9 2
5 2 13 9 9 2
19 2 0 9 3 3 0 9 0 1 9 13 9 9 9 1 0 9 9 2
17 1 12 0 9 0 9 13 7 13 1 9 2 9 15 14 13 2
9 2 13 2 16 1 9 3 4 2
5 13 2 9 9 2
8 2 13 1 9 1 9 0 2
4 2 13 3 2
4 2 13 9 2
6 3 13 2 9 9 2
3 2 13 2
11 13 9 9 9 1 9 13 9 7 9 2
5 2 14 13 9 2
17 2 14 13 2 16 13 2 7 13 4 3 2 9 9 2 2 2
9 14 9 9 9 13 13 0 9 2
6 2 14 13 2 2 2
8 2 3 2 9 9 2 13 2
5 2 13 9 9 2
4 13 1 9 2
4 13 1 9 2
2 13 2
4 13 1 13 2
14 2 3 4 13 9 1 9 9 1 9 9 9 9 2
3 2 13 2
5 13 4 0 9 2
7 2 9 9 2 9 13 2
14 2 14 13 2 9 9 2 13 13 14 1 12 9 2
6 1 9 13 0 9 2
4 2 13 3 2
16 0 9 13 9 13 1 9 9 0 9 13 1 9 9 9 2
5 2 13 9 9 2
8 14 9 9 9 13 13 9 2
8 9 9 13 1 9 4 13 2
3 13 3 2
9 13 14 4 13 1 0 0 9 2
8 2 9 13 1 13 0 9 2
4 9 15 13 2
8 13 1 13 1 9 9 9 2
7 13 2 16 9 9 13 2
4 13 1 9 2
4 13 12 9 2
11 9 13 3 9 1 13 9 9 7 9 2
12 1 0 9 13 4 1 9 1 13 9 9 2
4 13 1 9 2
13 2 13 9 0 9 2 1 9 9 4 1 9 2
3 2 13 2
3 13 3 2
4 9 15 13 2
7 13 2 16 9 9 13 2
4 13 12 9 2
7 9 13 1 13 0 9 2
4 13 1 9 2
14 2 13 2 16 9 1 13 0 9 9 9 9 13 2
7 9 0 2 14 13 4 2
5 9 15 14 13 2
17 2 14 9 1 9 9 7 9 9 13 13 9 1 9 13 9 2
5 13 7 1 9 2
4 9 15 13 2
9 1 13 1 9 9 13 3 3 2
4 2 13 9 2
4 9 15 13 2
4 13 12 9 2
13 13 2 16 9 1 13 0 9 9 9 9 13 2
12 2 13 2 16 9 13 9 9 0 9 9 2
4 13 1 9 2
7 9 13 1 13 0 9 2
12 13 2 16 13 15 9 1 9 13 9 0 2
3 13 9 2
11 1 9 13 4 9 0 0 2 9 9 2
6 2 9 9 4 13 2
11 1 0 13 9 9 13 1 0 9 9 2
5 2 13 9 9 2
4 13 1 9 2
13 13 2 16 9 1 13 0 9 9 9 9 13 2
4 9 15 13 2
4 13 12 9 2
16 9 7 9 9 13 4 9 9 9 9 7 9 9 9 9 2
6 2 13 1 13 9 2
3 13 9 2
16 1 0 9 9 9 4 9 9 9 9 7 9 9 9 9 2
5 13 9 13 9 2
2 13 2
5 2 13 12 9 2
16 1 12 9 13 9 7 9 9 2 7 13 0 9 1 9 2
3 2 13 2
14 2 13 2 16 9 1 13 0 9 9 9 9 13 2
7 9 13 1 13 0 9 2
6 2 13 9 0 9 2
15 2 13 9 2 7 3 15 13 9 1 0 9 2 2 2
9 2 9 9 2 14 13 4 9 2
4 13 1 9 2
4 9 15 13 2
7 9 13 1 13 0 9 2
15 9 0 14 4 13 9 9 2 14 13 14 1 9 9 2
5 13 2 9 9 2
18 2 13 14 1 9 1 9 9 9 0 9 0 2 13 1 9 0 2
10 2 1 13 1 9 9 13 3 3 2
9 2 9 9 13 1 9 4 13 2
6 9 3 15 14 13 2
3 13 9 2
11 0 9 1 0 8 2 13 0 9 9 2
14 3 13 0 2 7 13 1 9 0 7 0 9 0 2
2 13 2
10 13 15 9 7 9 9 1 13 9 2
9 2 9 9 13 1 9 4 13 2
6 1 9 13 9 13 2
3 13 9 2
11 9 13 3 0 2 0 2 0 7 0 2
7 2 14 9 13 0 9 2
7 1 9 14 13 4 9 2
11 1 0 9 1 15 0 9 13 3 0 2
11 1 0 9 9 13 15 1 0 9 9 2
11 3 9 9 13 13 15 1 9 0 9 2
6 13 15 14 0 9 2
4 2 13 9 2
5 13 15 15 3 2
9 14 1 9 0 1 9 13 4 2
5 3 13 15 3 2
10 3 13 1 9 2 13 15 7 13 2
4 9 9 13 2
5 9 13 14 13 2
5 14 9 14 13 2
4 13 0 9 2
16 9 9 4 13 1 0 9 13 9 1 9 1 0 9 0 2
4 14 13 9 2
14 7 14 2 16 4 15 13 2 13 14 4 15 9 2
9 9 13 9 7 13 15 1 9 2
7 3 15 1 9 13 4 2
7 1 9 9 13 15 3 2
23 13 4 1 9 2 7 3 13 4 3 9 9 2 1 0 9 2 0 9 2 0 9 2
5 9 13 9 0 2
11 0 9 9 13 1 9 1 9 9 9 2
21 9 9 2 9 9 9 0 9 9 2 13 3 9 1 9 1 13 9 1 9 2
20 9 1 0 9 0 13 14 9 2 0 13 9 1 12 9 1 9 1 9 2
8 9 13 3 0 1 9 9 2
33 3 13 9 9 1 9 1 9 9 2 13 3 9 13 2 16 9 13 9 13 15 1 9 2 13 9 1 9 9 7 9 0 2
14 9 2 13 1 0 9 2 13 13 15 1 9 9 2
4 9 13 3 2
13 13 15 2 13 12 0 9 7 13 9 1 9 2
10 13 15 1 12 9 7 1 9 13 2
12 1 12 9 9 13 12 3 13 15 1 9 2
10 13 15 3 2 7 3 13 1 9 2
7 14 9 13 15 1 9 2
7 7 3 13 9 0 9 2
6 15 3 13 13 9 2
12 13 4 15 1 15 2 16 13 13 9 9 2
20 3 0 9 14 13 7 1 0 9 14 13 4 2 1 0 9 13 1 9 2
13 1 9 13 13 15 9 9 1 0 1 9 9 2
30 13 4 2 16 14 13 13 15 9 9 9 2 16 15 0 9 13 15 1 9 2 7 1 9 0 13 14 13 4 2
4 9 13 15 2
7 2 3 15 13 0 9 2
7 9 13 2 3 9 13 2
12 9 13 14 3 2 16 0 9 13 13 0 2
8 2 14 3 3 14 14 13 2
4 9 13 3 2
16 13 4 15 0 9 7 13 9 2 0 13 15 1 9 0 2
7 2 15 13 3 1 9 2
12 13 4 1 0 9 7 13 4 9 1 9 2
13 15 14 13 4 3 0 2 7 13 4 1 9 2
6 13 4 3 1 9 2
4 9 13 9 2
8 2 1 9 13 15 3 3 2
14 2 16 15 15 14 13 2 13 13 0 9 2 2 2
7 2 14 13 15 0 9 2
5 2 13 0 9 2
4 9 13 9 2
6 9 13 9 0 9 2
13 9 13 1 12 9 2 1 9 13 15 0 9 2
6 9 3 3 13 9 2
7 1 9 13 15 9 9 2
12 13 15 9 0 1 0 13 1 9 9 0 2
15 9 0 9 13 0 9 9 2 0 9 9 13 1 9 2
7 3 1 9 13 9 9 2
15 9 13 12 9 9 2 9 2 9 2 9 0 2 9 2
8 0 9 13 15 9 13 9 2
12 9 1 9 13 9 0 9 9 0 1 9 2
11 9 7 9 13 3 9 1 13 9 0 2
32 13 15 2 16 9 0 4 13 13 1 9 1 9 1 12 9 7 16 0 0 9 1 9 1 9 1 9 4 13 9 9 2
10 13 15 9 1 9 1 12 0 9 2
8 0 9 13 1 9 1 9 2
4 3 13 0 2
8 3 13 15 9 1 13 9 2
9 2 1 9 13 1 15 0 9 2
10 9 3 13 9 7 13 1 15 9 2
20 13 2 16 13 2 7 14 13 13 0 9 9 7 9 1 9 1 0 9 2
20 7 14 13 2 3 13 1 9 9 13 9 1 13 1 9 9 0 9 0 2
15 13 2 16 13 2 7 14 13 13 0 9 13 1 9 2
6 3 9 13 0 9 2
4 13 0 9 2
7 9 13 1 9 1 9 2
16 13 0 9 1 9 1 9 2 0 9 13 1 9 0 9 2
7 1 9 9 9 13 9 2
10 2 9 1 9 13 15 15 0 9 2
2 13 2
5 2 13 9 0 2
13 9 13 9 9 0 2 0 13 0 9 0 9 2
32 0 1 9 9 9 0 13 13 15 1 0 9 2 7 9 4 13 1 9 0 1 9 1 9 7 14 13 15 0 9 0 2
24 1 9 0 9 1 8 2 0 9 13 9 2 7 9 1 0 0 9 1 15 13 1 9 2
15 14 13 4 1 0 9 7 13 2 16 13 13 0 9 2
7 2 13 15 1 0 9 2
6 14 13 15 1 9 2
10 0 9 13 15 9 2 13 3 13 2
10 2 3 15 13 2 3 15 13 2 2
10 2 14 13 9 7 13 1 0 9 2
10 0 9 8 2 13 14 9 0 9 2
30 13 1 0 9 9 9 8 2 2 13 1 9 9 2 4 13 1 9 9 1 9 2 7 3 13 7 13 1 9 2
9 9 13 15 1 9 0 7 0 2
10 15 9 13 15 1 9 7 9 9 2
6 0 9 13 15 9 2
7 2 13 4 15 1 9 2
11 16 14 15 9 13 0 2 3 13 4 2
9 1 12 9 14 13 1 15 9 2
5 13 4 15 12 2
4 2 13 9 2
8 2 13 1 9 9 9 9 2
10 2 14 13 1 0 9 13 0 9 2
6 2 7 3 9 13 2
3 13 4 2
8 13 4 1 15 3 1 9 2
3 2 13 2
7 7 3 13 2 3 13 2
2 13 2
12 13 4 15 2 13 4 7 13 4 1 9 2
5 13 4 14 9 2
12 13 4 15 9 13 1 9 2 0 1 9 2
11 13 15 1 13 2 16 9 13 15 9 2
11 1 12 13 9 2 16 9 15 15 13 2
8 7 3 13 1 15 0 9 2
8 2 13 2 13 15 7 13 2
7 13 4 15 1 0 9 2
6 9 9 14 15 13 2
7 2 0 9 14 14 13 2
9 9 9 13 0 9 7 13 9 2
6 3 9 13 15 3 2
6 1 0 9 13 9 2
7 9 9 13 3 9 0 2
8 0 13 15 1 0 0 9 2
5 13 13 13 9 2
8 9 9 13 2 16 9 13 2
7 13 3 1 9 9 0 2
4 13 1 9 2
12 0 9 13 15 1 9 0 1 9 1 9 2
13 1 9 1 9 1 9 1 13 9 13 0 9 2
14 2 9 0 13 9 9 0 1 13 0 9 1 9 2
8 7 13 13 1 9 1 9 2
5 2 13 9 0 2
18 15 15 13 2 13 9 2 13 2 3 13 9 2 0 13 15 9 2
8 13 9 2 13 1 15 9 2
19 2 1 9 9 2 0 3 3 3 13 9 7 9 2 14 13 9 9 2
8 2 9 9 13 14 1 9 2
11 0 0 9 13 14 1 0 0 9 9 2
9 9 3 13 1 0 9 0 9 2
12 0 9 13 14 1 9 2 3 2 1 9 2
5 14 13 13 9 2
22 2 0 9 1 9 13 9 13 1 9 1 9 2 1 0 3 13 8 2 9 9 2
11 3 1 9 13 0 9 2 16 13 9 2
18 2 12 1 15 3 13 1 9 1 9 2 7 14 15 9 13 9 2
11 15 14 13 0 9 7 14 13 1 9 2
8 1 9 14 13 15 13 9 2
25 14 13 13 9 2 16 1 9 2 1 9 2 1 9 13 13 9 1 9 2 0 9 14 13 2
15 9 13 9 3 1 9 2 7 13 9 7 9 15 13 2
9 14 13 1 0 9 1 0 9 2
9 2 9 13 0 9 9 9 0 2
11 9 13 15 2 16 9 14 0 14 13 2
7 9 1 9 13 0 9 2
14 13 2 9 4 13 2 13 1 9 2 13 1 9 2
13 16 9 3 13 1 0 9 2 13 4 3 13 2
8 2 13 1 9 13 1 9 2
8 2 1 9 9 0 9 13 2
10 2 14 2 14 4 4 13 1 9 2
6 9 13 15 0 9 2
10 14 3 15 9 13 1 9 12 9 2
11 13 15 14 13 2 9 9 13 2 2 2
13 2 3 13 9 9 2 0 13 1 9 12 9 2
12 3 13 9 4 14 13 9 1 12 9 0 2
24 0 9 9 13 14 2 16 9 0 3 4 13 3 13 2 13 14 9 9 9 7 9 0 2
14 1 0 9 1 0 9 9 13 15 13 0 0 9 2
12 13 9 9 9 0 7 0 2 7 14 9 2
10 0 9 13 3 14 14 13 9 9 2
8 2 14 13 4 9 0 9 2
15 1 9 3 13 9 1 0 9 13 9 9 2 9 13 2
9 0 9 0 13 15 1 15 0 2
10 15 9 13 0 9 1 9 0 9 2
9 9 13 2 16 0 13 1 9 2
11 3 4 13 1 9 1 0 3 0 9 2
7 2 3 1 15 15 13 2
15 7 16 13 9 0 12 9 2 14 13 13 9 9 0 2
14 14 9 9 13 4 1 9 0 2 7 0 7 0 2
17 9 14 13 2 16 9 7 9 1 9 13 15 0 9 7 9 2
13 2 14 0 9 4 13 1 9 1 0 9 0 2
12 2 14 9 9 1 9 14 13 1 13 9 2
9 2 9 13 9 9 3 13 9 2
12 7 0 0 9 13 12 9 2 7 12 9 2
11 3 1 9 13 4 15 1 0 0 9 2
8 3 3 13 7 4 3 13 2
4 9 13 0 2
22 13 1 9 2 3 3 13 15 1 9 9 2 0 3 13 0 9 1 9 13 9 2
13 13 14 0 2 16 0 9 13 9 9 0 9 2
17 3 9 2 0 4 13 1 9 1 9 13 2 13 15 13 9 2
8 2 12 13 14 1 9 9 2
15 1 0 9 9 9 13 9 0 2 0 9 13 1 9 2
9 9 9 1 13 0 9 13 0 2
21 0 9 1 9 7 9 0 13 9 9 7 9 9 2 9 2 9 7 9 9 2
5 13 14 12 9 2
9 1 3 13 9 3 13 2 2 2
29 1 9 0 2 12 9 2 13 15 9 13 0 9 2 13 1 9 1 3 13 9 0 2 9 2 9 7 9 2
9 9 13 1 9 9 13 1 9 2
9 9 13 14 9 1 13 0 9 2
9 2 13 4 3 9 1 9 9 2
11 14 1 0 0 9 3 15 1 15 13 2
18 13 1 9 2 1 0 9 13 3 13 9 0 9 7 9 0 9 2
10 2 14 13 15 0 9 9 9 0 2
8 2 4 13 0 9 1 9 2
11 14 14 13 15 9 9 9 1 9 0 2
11 13 12 9 0 7 13 14 12 9 0 2
26 9 9 13 1 9 14 1 9 0 2 2 3 13 15 1 9 0 2 1 0 13 14 1 9 0 2
5 13 9 0 9 2
8 2 9 1 3 14 4 13 2
7 9 15 13 13 14 9 2
6 7 3 13 14 13 2
13 2 9 9 13 2 16 13 0 9 13 0 9 2
4 3 4 13 2
7 3 9 13 1 12 9 2
6 9 13 1 9 3 2
10 1 14 12 9 13 1 9 9 9 2
12 13 9 0 9 0 2 0 9 4 3 13 2
8 0 9 3 13 1 9 0 2
11 7 16 3 4 13 2 7 4 9 13 2
3 16 13 2
11 2 9 13 15 1 9 13 7 13 9 2
18 13 3 13 9 9 0 2 16 3 13 1 9 7 9 3 13 9 2
6 9 13 2 9 13 2
8 9 13 14 12 9 9 9 2
14 2 9 9 13 12 8 8 2 9 0 9 14 13 2
11 2 9 7 9 0 13 1 9 9 0 2
8 9 13 15 1 12 9 0 2
9 14 9 13 13 9 1 15 9 2
8 3 13 15 9 1 9 0 2
16 0 9 1 12 9 13 2 16 9 0 9 0 3 15 13 2
7 3 0 9 13 15 9 2
11 2 0 13 15 1 9 2 1 9 9 2
10 2 9 1 12 9 13 1 9 9 2
17 13 0 9 9 2 13 9 1 9 1 0 9 2 9 2 9 2
16 2 16 9 7 9 14 13 9 2 7 0 13 13 0 9 2
15 2 1 9 1 13 9 0 9 13 0 9 1 9 0 2
4 9 13 9 2
11 1 9 0 13 15 14 9 0 7 0 2
7 1 9 13 0 9 0 2
14 3 15 13 2 14 13 2 13 2 13 0 3 9 2
10 2 13 4 0 9 2 15 15 13 2
7 9 13 13 9 1 9 2
20 14 3 13 15 1 0 9 0 2 16 13 9 1 9 9 13 1 9 9 2
27 9 13 2 16 1 9 1 13 9 13 15 9 13 15 1 9 1 9 0 9 1 9 13 1 9 9 2
5 13 1 13 9 2
6 3 9 13 15 9 2
6 3 13 3 0 9 2
15 9 9 9 13 0 9 2 13 1 9 13 15 9 9 2
12 13 14 9 1 9 1 0 9 7 9 9 2
9 14 13 9 2 16 13 0 9 2
12 1 0 9 9 13 14 9 13 0 9 0 2
19 13 15 15 2 16 13 14 9 0 13 9 1 9 0 7 13 9 0 2
9 13 2 16 9 14 13 3 0 2
7 13 15 2 16 15 13 2
11 1 0 9 14 13 2 16 9 13 0 2
10 13 9 1 0 9 2 9 13 9 2
7 9 9 13 9 9 0 2
9 1 9 9 1 9 13 9 0 2
4 4 3 13 2
14 4 13 0 9 2 3 1 9 9 13 12 9 9 2
26 14 0 9 9 9 9 13 0 9 7 13 2 16 4 13 15 9 1 9 9 9 7 9 9 9 2
19 9 13 2 16 1 9 14 13 15 0 9 1 9 9 0 13 1 9 2
11 2 14 13 4 15 2 9 13 2 9 2
5 2 13 2 13 2
3 13 15 2
4 3 13 3 2
11 13 4 1 15 9 9 1 9 9 0 2
6 9 4 14 13 3 2
7 13 15 2 3 13 9 2
8 2 1 9 14 13 14 4 2
6 13 1 15 1 9 2
11 2 13 4 15 2 16 3 13 2 9 2
6 2 13 14 4 2 2
15 2 14 13 2 9 2 13 9 1 9 1 9 9 9 2
9 13 2 16 13 0 9 2 2 2
6 13 9 9 2 2 2
11 9 13 1 9 2 13 3 1 0 9 2
5 9 13 3 0 2
6 2 13 9 2 9 2
9 9 1 9 14 13 15 1 9 2
7 14 13 15 15 9 0 2
9 2 14 0 9 13 15 1 9 2
8 2 13 2 16 9 15 13 2
5 9 13 1 9 2
7 2 13 3 2 9 0 2
4 9 13 0 2
7 9 13 9 3 1 15 2
6 9 13 15 1 9 2
8 9 9 13 15 1 9 3 2
7 2 13 4 3 2 2 2
9 13 15 2 16 9 14 13 4 2
6 2 3 15 13 2 2
6 2 15 9 13 3 2
9 2 14 13 2 9 13 2 9 2
9 2 14 13 12 0 1 0 9 2
11 9 13 15 3 2 13 9 9 1 9 2
6 14 13 14 12 0 2
8 13 3 0 9 2 0 9 2
11 13 3 15 9 2 13 15 1 9 9 2
7 9 4 13 1 9 9 2
13 0 9 1 3 14 13 9 1 0 9 0 9 2
7 9 0 9 0 4 13 2
8 13 15 3 1 9 9 0 2
9 0 13 9 1 13 9 1 9 2
7 13 13 13 0 1 9 2
7 3 14 13 1 9 9 2
13 13 9 9 9 2 1 0 3 13 1 12 9 2
10 9 13 1 9 9 1 9 1 9 2
10 9 0 13 9 9 9 0 9 0 2
8 1 0 9 13 15 9 9 2
6 3 13 0 9 0 2
7 1 0 13 0 9 0 2
10 13 15 9 2 9 2 9 7 9 2
12 9 9 0 1 9 0 13 1 15 0 9 2
9 13 0 9 0 13 9 1 9 2
27 15 9 1 9 13 9 1 13 9 2 9 1 9 1 0 9 2 0 1 9 13 1 15 9 0 9 2
9 9 13 15 1 0 9 1 9 2
11 1 0 13 2 16 9 0 14 13 9 2
3 14 13 2
15 14 1 9 9 0 3 14 13 15 15 3 13 1 9 2
10 3 13 15 9 1 9 9 2 2 2
7 12 1 15 13 1 9 2
13 1 9 1 9 12 9 13 13 15 1 9 9 2
12 12 9 2 0 9 13 0 2 13 1 9 2
8 1 9 13 15 14 12 9 2
7 14 2 9 14 13 9 2
21 1 15 9 9 14 14 13 0 9 2 1 0 1 0 9 13 15 9 13 9 2
17 9 9 1 9 9 0 9 13 15 9 1 9 1 8 2 0 2
7 1 9 13 15 1 9 2
7 9 13 1 8 2 9 2
9 9 0 13 1 0 2 0 9 2
12 0 9 13 1 9 2 16 15 1 15 13 2
7 9 13 14 0 2 0 2
5 13 15 14 13 2
7 14 13 14 15 1 9 2
10 9 13 1 15 9 7 13 4 15 2
5 2 13 9 0 2
7 2 13 4 0 0 9 2
8 13 4 2 16 3 15 13 2
5 2 9 13 9 2
7 13 15 1 9 2 13 2
15 1 9 13 9 7 9 13 2 7 9 13 13 9 0 2
16 16 9 13 12 2 1 9 0 13 2 16 12 9 13 0 2
8 9 1 9 13 9 13 9 2
12 1 9 13 15 2 16 13 13 3 1 9 2
20 1 9 13 0 9 1 9 9 9 2 13 1 9 9 2 14 3 13 9 2
18 14 1 9 13 4 15 13 2 12 13 9 1 0 9 1 0 9 2
6 13 15 15 7 13 2
17 9 13 3 14 3 2 13 4 9 0 2 0 7 3 14 13 2
15 0 9 2 0 13 2 13 1 9 2 7 9 14 13 2
3 9 13 2
11 4 13 9 3 0 1 9 14 1 9 2
13 9 0 15 13 9 2 9 2 9 9 7 9 2
10 9 0 13 4 1 0 1 0 9 2
10 13 15 12 9 0 9 1 0 9 2
17 1 9 13 4 3 12 9 1 9 13 3 1 9 0 7 0 2
10 13 4 2 3 0 9 13 1 9 2
9 7 9 1 0 12 9 13 0 2
15 13 9 1 0 9 2 9 7 9 13 15 0 9 0 2
5 13 15 15 3 2
5 2 9 15 13 2
10 2 13 1 9 9 1 9 13 9 2
6 13 4 0 2 9 2
6 2 9 9 13 3 2
5 2 13 1 9 2
10 14 13 4 9 1 9 7 13 4 2
12 16 13 4 13 2 13 15 1 12 9 3 2
9 13 0 2 7 3 14 15 13 2
7 2 9 9 13 1 9 2
6 15 14 3 4 9 2
9 2 15 13 4 3 1 0 9 2
13 1 13 1 9 9 13 1 9 1 9 1 13 2
8 9 13 15 1 9 1 9 2
6 2 14 15 3 13 2
4 3 13 9 2
26 1 0 8 2 13 9 9 0 9 0 2 7 1 0 8 2 13 9 9 9 0 2 0 9 0 2
7 9 13 0 9 1 9 2
4 13 0 9 2
10 7 13 9 1 3 0 9 1 9 2
16 13 15 1 15 13 0 9 9 1 9 2 9 7 9 9 2
3 14 13 2
4 3 13 9 2
16 1 9 14 13 9 0 9 2 13 15 7 3 13 1 9 2
10 2 13 2 9 9 13 2 2 2 2
20 3 9 1 9 0 13 0 9 2 1 9 7 9 13 1 15 14 9 9 2
9 3 13 1 0 9 0 0 9 2
8 13 1 9 0 2 0 9 2
5 3 14 4 13 2
4 3 13 9 2
7 15 0 9 4 3 13 2
7 0 9 13 15 3 0 2
7 9 0 3 13 15 9 2
7 9 13 9 1 9 9 2
24 9 1 9 13 1 9 0 1 12 9 7 9 13 1 0 9 13 9 13 2 13 7 13 2
10 1 15 9 13 15 14 12 0 9 2
10 9 13 15 1 9 0 9 9 9 2
12 9 0 13 2 16 9 13 1 9 9 0 2
23 1 9 2 1 9 0 1 14 12 9 13 15 9 1 9 7 0 9 13 9 9 9 2
5 13 9 0 9 2
11 2 13 2 16 9 3 15 13 0 9 2
6 14 9 13 9 9 2
9 7 9 15 14 1 0 9 13 2
11 9 1 9 13 15 1 9 1 0 9 2
7 7 13 1 9 0 9 2
14 0 9 0 13 3 9 9 7 13 9 9 0 9 2
17 13 15 9 0 2 9 15 1 0 14 13 2 7 0 13 0 2
15 9 3 13 9 1 9 2 16 13 2 3 13 15 9 2
14 3 0 9 13 15 3 2 13 15 9 9 0 9 2
25 9 9 13 15 1 9 2 7 9 7 9 14 13 13 15 1 15 7 9 15 9 13 9 9 2
15 9 13 0 7 0 2 13 1 9 2 16 13 15 9 2
11 16 9 13 1 9 2 9 13 0 9 2
19 13 1 9 9 9 13 9 2 7 9 13 7 13 15 1 9 1 13 2
11 0 9 13 1 9 9 3 13 9 9 2
9 1 0 9 13 9 13 0 9 2
8 0 0 9 4 13 7 13 2
6 1 9 13 0 9 2
8 9 13 0 9 1 0 9 2
15 9 13 15 1 9 9 7 13 13 9 1 0 9 9 2
4 2 13 15 2
10 9 13 9 7 13 1 15 0 9 2
10 2 13 3 2 16 15 1 15 13 2
5 2 9 13 9 2
5 2 13 1 9 2
4 13 15 15 2
6 2 9 13 0 9 2
10 2 13 9 7 13 1 15 1 9 2
9 9 13 1 0 9 1 9 0 2
8 13 2 16 13 0 0 9 2
10 9 13 2 16 9 9 0 13 9 2
8 9 0 13 9 1 9 9 2
15 9 9 13 1 15 9 0 7 9 0 1 9 7 9 2
15 1 9 14 9 13 1 0 9 9 13 9 0 9 9 2
10 9 9 13 12 9 1 0 9 9 2
9 14 1 9 0 9 13 3 0 2
23 9 0 7 0 13 14 0 2 13 0 9 7 9 0 2 7 14 9 0 1 9 0 2
12 1 9 9 13 9 7 9 0 1 9 9 2
4 2 3 13 2
4 9 14 13 2
13 9 13 13 0 2 0 2 1 9 1 9 13 2
9 3 1 9 14 0 9 14 13 2
12 2 7 15 3 9 0 2 0 2 13 13 2
23 9 13 2 16 9 13 3 1 0 0 9 2 3 13 15 2 13 7 13 1 0 9 2
3 3 13 2
6 9 9 13 0 9 2
3 14 13 2
9 2 12 9 2 9 9 2 13 2
9 9 0 14 13 14 3 0 3 2
7 13 9 0 7 9 9 2
16 3 13 15 9 0 2 0 2 0 7 0 0 2 9 0 2
6 2 0 15 15 13 2
7 9 13 15 1 9 9 2
10 7 13 2 16 9 0 13 13 9 2
5 2 13 9 9 2
4 13 9 9 2
5 13 14 9 9 2
5 2 13 2 2 2
7 1 9 9 9 3 13 2
5 14 13 2 2 2
4 13 15 13 2
8 2 9 2 14 13 1 9 2
10 9 0 13 2 16 4 13 2 2 2
6 14 13 15 2 2 2
6 2 14 13 1 9 2
7 13 3 2 13 15 9 2
7 13 9 1 9 2 2 2
7 13 4 15 9 2 2 2
13 7 0 0 9 13 2 16 15 3 13 2 2 2
8 2 13 0 9 9 2 2 2
6 2 13 3 2 2 2
12 3 12 13 14 1 9 9 2 9 13 3 2
4 0 9 13 2
7 9 9 14 13 1 9 2
6 0 9 13 14 9 2
7 3 14 4 13 9 9 2
7 9 3 14 13 1 9 2
18 3 13 1 0 9 9 13 9 13 9 9 1 9 2 9 7 9 2
8 13 15 1 9 9 9 0 2
24 1 9 9 14 13 9 1 9 2 13 14 1 0 9 0 7 0 2 13 15 1 0 9 2
19 9 9 13 9 9 9 0 9 9 9 0 9 1 13 15 1 13 9 2
21 9 9 13 14 2 16 13 13 1 9 0 9 1 9 9 9 1 9 7 9 2
14 2 1 9 9 3 3 13 9 13 9 13 1 9 2
8 9 9 13 13 1 9 9 2
10 3 13 9 2 1 9 0 9 13 2
10 13 2 16 14 3 4 13 13 9 2
13 14 2 3 13 9 2 9 9 0 3 15 13 2
13 13 15 2 13 9 2 13 1 9 7 13 9 2
9 9 13 13 15 1 0 9 9 2
5 13 9 2 13 2
4 2 13 15 2
8 2 13 15 2 13 9 9 2
6 3 13 1 9 9 2
11 9 13 9 1 9 7 13 15 1 9 2
17 16 9 13 15 9 7 13 14 0 9 2 13 1 15 1 9 2
17 1 9 9 9 9 13 3 0 2 16 9 13 9 13 3 0 2
21 9 13 7 9 7 1 9 9 9 13 13 0 9 9 7 13 15 14 0 9 2
8 9 13 9 2 13 9 9 2
5 13 15 1 9 2
8 3 3 13 2 16 3 13 2
7 1 9 13 0 0 9 2
4 13 4 9 2
4 2 14 13 2
5 9 3 14 13 2
6 2 13 15 0 9 2
14 1 9 0 0 9 13 15 2 16 13 15 1 9 2
6 0 0 9 13 9 2
17 9 1 9 13 9 0 1 9 2 0 1 9 13 1 9 9 2
13 3 1 0 9 13 9 9 0 1 0 9 0 2
7 9 13 9 1 12 9 2
8 9 0 13 14 0 9 9 2
6 7 14 15 13 9 2
3 13 9 2
7 0 9 7 14 9 13 2
7 14 13 15 1 0 9 2
2 13 2
4 13 1 9 2
3 9 13 2
2 13 2
11 9 1 9 13 1 0 15 9 0 9 2
8 12 13 15 1 0 9 9 2
8 9 1 9 13 0 9 9 2
14 14 2 1 9 13 3 7 0 9 13 14 4 13 2
12 9 1 9 13 2 16 1 9 0 13 9 2
17 0 9 1 9 13 14 1 9 9 2 0 3 13 9 1 9 2
10 9 15 13 13 9 9 9 9 9 2
18 1 9 3 13 15 13 1 9 0 9 1 0 9 13 1 9 9 2
7 0 9 13 15 0 9 2
6 9 9 3 13 9 2
14 13 15 9 13 3 2 16 0 9 9 14 4 13 2
17 13 1 9 13 1 0 9 9 0 2 3 0 1 9 7 9 2
4 9 15 13 2
11 7 0 13 14 1 9 2 9 1 9 2
12 16 1 0 9 0 9 14 12 14 13 9 2
9 15 9 14 13 2 14 1 9 2
6 2 0 9 14 13 2
7 1 9 9 13 15 9 2
7 3 13 15 3 0 9 2
6 13 4 0 0 9 2
24 1 9 13 9 2 16 13 4 1 0 0 9 2 0 13 15 9 1 9 7 0 9 9 2
8 2 9 13 1 15 0 9 2
6 13 4 15 1 9 2
10 0 9 14 13 14 1 9 9 9 2
9 13 14 15 12 9 2 3 0 2
2 13 2
10 9 13 9 2 7 9 13 15 13 2
8 9 4 13 1 0 0 9 2
9 3 14 15 9 0 13 0 9 2
4 9 3 13 2
5 13 3 0 9 2
5 7 14 13 13 2
7 13 0 9 1 9 9 2
6 14 13 15 1 9 2
13 13 9 9 2 7 9 13 13 9 0 1 15 2
6 3 13 9 7 9 2
6 15 14 13 1 9 2
10 0 9 9 1 9 13 1 0 9 2
9 2 13 4 3 0 7 0 9 2
8 13 14 14 0 9 9 0 2
11 3 14 9 9 13 15 1 9 0 9 2
14 1 15 9 13 15 9 0 2 3 13 4 0 9 2
15 0 9 13 12 9 2 16 13 9 2 9 13 14 9 2
6 0 1 9 13 9 2
20 0 9 2 0 4 15 13 2 1 0 9 1 9 9 13 9 0 1 9 2
9 9 13 15 14 1 9 1 9 2
7 0 9 13 9 7 9 2
8 9 13 1 9 1 0 9 2
15 1 0 9 13 9 0 9 2 7 14 9 7 9 9 2
13 13 1 0 9 8 2 2 9 0 1 0 9 2
7 9 15 13 1 0 9 2
8 13 3 0 9 7 13 9 2
5 9 3 13 9 2
14 9 13 15 9 7 13 13 3 0 9 1 0 9 2
7 3 9 14 13 1 15 2
4 13 13 9 2
6 13 15 13 1 9 2
11 1 9 1 9 0 9 13 1 9 9 2
3 13 9 2
10 16 13 1 9 9 2 13 1 15 2
10 9 2 13 9 2 3 13 1 9 2
8 13 1 9 2 16 13 9 2
10 13 9 0 1 9 9 0 1 9 2
8 1 9 13 3 1 12 9 2
8 2 13 3 0 1 13 9 2
8 13 4 3 12 9 9 0 2
10 9 0 1 9 13 1 9 3 13 2
16 13 2 16 1 9 13 3 2 16 13 4 13 1 9 9 2
4 7 9 13 2
13 2 3 13 4 15 1 9 2 13 4 0 9 2
15 13 14 9 9 2 0 14 13 2 16 13 9 1 9 2
13 9 0 0 9 3 14 13 9 9 1 9 0 2
11 1 9 9 9 1 9 13 15 3 3 2
11 1 9 9 9 3 13 0 9 9 0 2
25 1 15 9 1 0 9 3 13 9 9 0 1 0 9 0 2 13 9 1 9 9 0 2 0 2
7 3 13 9 0 9 9 2
11 1 12 9 13 1 9 0 9 1 9 2
16 9 0 7 0 2 9 2 9 2 9 7 9 13 0 9 2
18 0 9 13 9 1 9 9 1 0 9 9 13 4 14 1 0 9 2
12 0 9 13 1 9 1 9 0 9 1 9 2
5 9 15 13 9 2
10 9 13 0 0 9 2 9 9 9 2
5 13 15 1 9 2
17 1 9 0 9 1 9 9 0 7 0 9 13 1 9 0 9 2
3 13 4 2
5 2 13 1 9 2
8 13 15 2 16 9 13 9 2
13 9 9 13 0 9 9 2 0 0 9 1 9 2
7 9 13 1 9 0 9 2
6 9 13 15 3 0 2
14 1 12 0 9 3 0 9 13 2 7 3 15 13 2
16 1 0 1 9 0 12 0 9 13 1 9 13 1 15 9 2
19 2 9 2 13 15 9 2 7 15 15 13 9 1 9 7 9 1 9 2
5 13 3 12 9 2
7 9 1 15 13 1 15 2
10 13 2 14 13 7 0 9 14 13 2
6 3 14 13 0 9 2
11 0 9 1 0 9 13 9 9 1 9 2
10 0 9 9 13 15 1 9 1 9 2
13 0 9 1 9 13 15 1 9 2 9 7 9 2
13 3 1 9 13 9 9 2 9 9 7 9 9 2
17 7 0 9 1 0 9 13 1 15 7 13 4 13 15 1 3 2
16 9 3 13 2 16 13 15 9 1 0 9 1 9 9 9 2
13 3 3 1 9 8 2 9 13 0 9 1 9 2
25 13 1 15 2 16 4 13 1 3 0 9 2 1 0 13 15 9 1 0 9 1 9 7 9 2
10 9 9 2 9 9 2 13 3 9 2
9 13 12 9 13 9 1 9 0 2
7 9 13 9 9 1 9 2
10 9 1 13 9 1 9 0 3 13 2
5 3 13 9 9 2
8 1 0 9 9 13 0 9 2
19 13 3 1 12 9 2 0 13 1 0 9 2 3 3 13 15 1 9 2
13 13 14 2 16 13 1 9 9 1 3 0 9 2
23 9 1 9 9 9 7 0 9 13 9 1 0 9 0 9 1 9 9 1 9 7 9 2
9 9 9 13 0 9 7 0 9 2
6 9 0 13 3 9 2
4 3 14 13 2
6 3 7 13 7 13 2
13 0 9 13 12 0 9 1 9 13 9 7 9 2
11 1 13 1 0 9 9 13 12 9 9 2
2 13 2
7 3 15 3 13 1 9 2
5 3 15 15 13 2
6 13 15 13 0 9 2
11 13 2 16 9 0 13 15 3 14 3 2
9 9 13 1 12 9 1 0 9 2
10 0 9 9 13 9 1 13 9 0 2
13 1 9 9 1 0 9 13 7 13 15 1 9 2
13 9 1 12 9 9 0 13 3 9 1 9 0 2
14 3 13 2 16 4 13 0 9 1 13 9 9 0 2
8 9 9 13 9 9 0 9 2
20 2 9 13 1 9 2 13 9 2 13 9 2 7 13 12 9 1 0 9 2
13 2 14 0 9 13 0 7 14 13 3 0 9 2
5 3 9 13 9 2
5 13 13 0 9 2
9 3 9 13 15 1 0 9 9 2
10 3 3 15 13 1 13 9 0 9 2
5 3 13 9 9 2
13 1 9 1 9 0 2 0 1 9 13 12 9 2
17 0 9 13 1 9 9 1 9 2 9 9 7 9 13 1 9 2
15 9 8 2 13 14 9 2 13 0 7 13 0 9 9 2
14 9 9 13 9 14 14 0 9 2 0 13 15 9 2
11 9 9 13 15 14 3 0 9 13 9 2
15 13 2 16 15 9 13 9 12 7 16 15 9 13 9 2
4 8 15 13 2
15 14 13 14 14 1 9 0 9 7 13 14 15 9 9 2
4 9 13 9 2
13 15 1 9 9 9 13 14 4 9 13 0 9 2
9 15 3 3 14 4 9 14 13 2
6 7 13 1 15 13 2
14 1 15 9 9 0 4 13 7 13 3 1 9 0 2
10 13 9 9 7 9 2 9 15 9 2
26 16 1 9 9 13 15 0 2 13 1 9 9 2 9 13 1 9 2 7 1 15 13 15 9 9 2
28 9 13 2 16 13 2 13 2 13 15 2 13 2 13 13 13 1 9 9 7 3 13 15 1 15 2 2 2
12 14 13 15 9 9 1 9 0 7 9 0 2
10 1 9 1 9 13 15 0 9 0 2
12 0 13 15 9 0 9 1 9 1 12 8 2
4 13 12 9 2
10 9 9 1 9 3 13 1 0 9 2
7 14 13 13 1 9 9 2
26 3 9 13 9 8 2 0 2 16 9 2 16 13 15 1 9 2 13 13 1 15 0 9 0 9 2
9 1 9 1 9 9 13 15 9 2
8 0 9 13 9 9 1 9 2
9 1 9 9 9 9 13 1 9 2
6 0 13 1 9 9 2
16 0 9 9 3 13 9 0 2 9 0 2 9 2 0 9 2
4 1 9 13 2
9 1 9 9 13 15 13 9 9 2
10 1 15 13 0 9 1 9 1 9 2
28 1 0 9 13 15 1 9 9 2 13 9 2 13 9 0 1 9 0 9 2 13 13 9 0 2 13 9 2
11 13 1 9 9 9 3 13 1 15 9 2
10 0 0 9 3 1 9 13 1 9 2
4 9 3 13 2
9 9 1 0 9 9 13 13 9 2
16 9 13 0 9 9 0 1 0 9 7 9 2 13 1 9 2
9 3 13 1 9 7 3 13 9 2
21 0 3 14 13 13 1 9 9 1 0 9 2 16 3 1 9 13 0 9 9 2
4 13 15 3 2
8 7 9 13 1 9 9 9 2
7 13 14 1 13 15 9 2
4 13 1 0 2
7 9 9 13 1 9 0 2
6 2 9 13 9 9 2
8 1 0 0 9 13 14 9 2
8 2 13 0 0 9 2 9 2
13 7 13 0 9 2 16 3 13 4 2 16 13 2
6 2 13 3 0 9 2
6 2 14 9 13 0 2
25 2 3 13 9 2 16 0 9 1 9 0 13 9 0 2 7 1 9 13 15 1 9 13 2 2
8 3 9 1 13 13 3 0 2
7 1 0 9 13 9 0 2
7 13 14 0 9 1 9 2
4 13 15 12 2
8 14 13 2 3 15 13 4 2
16 13 1 9 1 0 9 1 9 2 1 0 13 15 9 9 2
8 9 0 13 0 9 9 9 2
12 1 9 0 1 9 13 3 3 9 1 9 2
10 13 13 2 3 0 9 13 1 9 2
9 1 0 9 0 9 13 9 9 2
23 9 8 2 13 15 14 2 16 13 1 9 13 0 9 13 9 1 9 0 9 9 9 2
34 1 9 9 2 16 0 9 9 13 15 1 9 2 13 1 15 9 13 1 9 2 1 9 1 9 2 7 13 13 9 1 9 9 2
11 9 9 4 13 1 9 0 0 9 9 2
19 13 4 2 16 14 4 15 13 1 9 2 7 13 15 7 13 4 9 2
4 14 13 9 2
8 7 12 9 14 13 1 9 2
22 7 13 15 15 2 16 9 2 9 7 9 13 3 3 13 1 9 2 9 7 9 2
11 13 0 9 2 16 3 13 13 13 9 2
7 7 14 3 15 14 13 2
12 7 9 1 9 13 0 9 0 2 2 2 2
6 9 13 15 15 3 2
6 9 3 13 1 9 2
5 7 13 1 9 2
13 0 13 3 9 13 7 0 9 13 1 0 9 2
5 9 13 1 9 2
19 1 9 13 9 13 15 9 9 7 13 0 1 9 2 3 1 9 9 2
6 9 14 4 3 13 2
13 7 9 13 1 15 2 13 15 1 9 7 13 2
17 7 9 9 9 1 15 13 2 7 15 15 13 1 12 9 0 2
7 3 3 1 0 9 13 2
40 7 13 9 2 16 3 9 13 2 7 13 0 0 9 2 16 1 15 9 14 3 1 9 9 14 13 2 7 1 0 9 13 9 7 15 1 9 3 13 2
11 7 14 13 2 16 13 15 9 1 0 2
7 13 2 16 14 13 4 2
8 7 14 13 2 16 3 13 2
3 13 13 2
11 9 13 0 9 7 13 1 9 0 9 2
4 13 1 9 2
4 9 14 13 2
7 2 7 9 3 14 13 2
3 14 13 2
6 2 7 3 13 15 2
6 2 16 15 13 4 2
28 9 4 13 1 0 9 7 13 0 9 9 9 7 9 2 1 0 9 0 9 13 9 9 1 9 9 9 2
16 1 9 13 13 9 0 2 0 13 3 1 0 9 13 9 2
24 1 0 9 1 9 13 15 9 2 16 13 2 14 4 13 9 13 15 1 9 13 9 0 2
3 13 9 2
17 3 3 13 15 1 9 1 9 2 0 7 0 1 9 1 9 2
7 13 1 9 12 9 9 2
7 7 14 13 1 9 0 2
10 7 0 13 9 0 9 9 1 9 2
6 0 13 1 15 9 2
7 7 14 13 4 13 3 2
9 13 15 9 9 7 9 0 9 2
2 13 2
8 14 14 4 3 13 9 3 2
10 13 13 2 16 1 9 14 13 9 2
8 7 9 13 14 9 1 9 2
8 3 14 1 9 13 13 9 2
10 3 14 1 0 9 13 15 9 9 2
14 13 15 3 1 9 9 0 2 13 3 0 9 0 2
15 3 13 13 9 9 1 9 2 16 9 14 13 14 0 2
13 3 13 9 7 15 9 2 1 0 13 9 13 2
7 13 1 0 9 12 9 2
8 1 0 9 13 15 13 9 2
16 16 9 3 13 15 1 9 2 13 9 2 16 4 3 13 2
6 9 13 15 13 9 2
7 0 9 1 9 13 3 2
6 2 9 13 3 0 2
7 1 9 13 4 9 9 2
4 13 0 9 2
11 1 9 13 4 3 2 9 13 14 13 2
8 2 13 3 0 9 2 2 2
3 13 9 2
4 9 13 9 2
9 9 0 13 7 13 1 9 9 2
5 3 15 14 13 2
11 2 13 9 9 7 13 2 13 1 15 2
4 2 13 14 2
10 2 14 13 3 2 14 13 1 9 2
4 16 13 0 2
10 12 9 1 13 14 4 1 0 9 2
3 3 13 2
5 3 14 13 4 2
17 1 9 2 1 9 2 13 9 7 9 2 7 1 9 13 9 2
12 3 13 4 0 9 7 13 4 9 1 9 2
6 13 9 7 13 13 2
14 9 3 13 2 7 1 9 9 13 15 9 13 9 2
7 13 9 9 1 0 9 2
4 9 15 13 2
6 2 9 9 14 13 2
5 2 13 14 13 2
7 14 2 14 13 2 9 2
8 2 14 13 9 2 3 13 2
13 16 9 9 3 3 13 1 9 2 13 1 9 2
3 2 13 2
3 13 15 2
6 14 13 9 15 13 2
8 9 4 13 2 9 13 13 2
9 14 13 2 16 13 15 1 9 2
12 2 13 9 1 9 2 3 0 2 0 13 2
3 2 13 2
21 1 9 13 15 9 2 7 15 2 1 9 2 4 13 7 13 3 1 0 9 2
3 2 13 2
8 2 9 13 2 16 13 9 2
9 13 15 1 9 13 2 13 9 2
11 9 13 0 9 13 1 0 8 2 9 2
15 9 1 9 13 9 0 1 12 8 2 7 9 3 13 2
15 9 9 13 2 16 1 12 9 9 14 13 3 0 9 2
11 3 4 0 9 2 1 9 14 12 9 2
14 9 9 2 0 9 9 2 13 3 9 1 9 9 2
3 4 13 2
18 1 9 13 12 9 9 2 1 9 12 13 9 9 0 14 1 9 2
13 1 9 1 8 2 0 2 12 13 15 0 9 2
8 1 0 9 0 9 13 0 2
5 13 15 3 13 2
5 9 13 1 9 2
10 9 13 15 1 9 7 13 1 15 2
12 3 1 9 13 9 2 13 3 1 9 9 2
6 13 9 13 1 9 2
12 3 9 13 9 7 3 1 9 13 1 9 2
10 13 0 9 2 16 13 15 0 9 2
10 1 9 13 15 1 0 9 9 0 2
23 13 9 1 9 2 13 15 9 9 1 9 9 7 14 13 15 3 2 16 13 1 9 2
22 16 9 13 15 14 1 9 1 9 2 9 13 9 1 9 0 9 2 9 7 9 2
10 9 9 13 15 3 9 7 0 9 2
8 9 7 0 9 13 3 3 2
6 0 9 13 0 9 2
7 13 15 1 9 0 9 2
5 9 13 3 3 2
7 9 9 9 9 13 9 2
11 14 13 14 2 3 1 15 1 9 13 2
9 13 13 9 9 1 13 9 9 2
5 13 13 3 3 2
11 1 13 9 7 13 9 9 13 1 9 2
7 9 13 8 2 9 9 2
6 9 13 9 9 9 2
11 9 13 15 1 9 9 1 0 0 9 2
13 12 9 13 1 9 13 0 9 13 1 9 9 2
17 1 0 9 13 4 1 9 9 7 0 9 3 15 1 0 13 2
6 13 0 0 0 9 2
19 0 9 13 4 15 1 9 2 13 4 9 1 9 2 3 13 1 9 2
11 1 9 9 0 13 4 1 9 1 9 2
14 13 15 14 3 2 16 13 4 15 2 9 4 13 2
14 2 1 12 9 1 9 0 13 15 12 0 9 0 2
15 3 9 14 13 1 9 0 13 1 9 0 9 1 9 2
13 1 9 1 0 9 9 9 13 9 9 7 9 2
14 0 9 13 4 9 9 9 1 9 0 1 9 9 2
9 1 0 9 9 13 7 1 9 2
6 9 13 14 12 9 2
9 9 13 9 9 2 13 3 9 2
8 14 9 13 1 9 0 9 2
12 9 13 2 16 13 1 9 1 12 9 9 2
17 1 9 1 9 9 13 15 1 9 0 9 0 1 3 0 9 2
14 13 9 2 16 15 0 9 13 4 9 9 13 9 2
14 1 9 13 9 0 9 0 2 9 9 13 3 0 2
14 9 13 15 1 0 9 2 1 9 9 1 0 9 2
7 13 3 9 9 0 9 2
13 4 15 1 9 0 9 0 0 9 1 9 9 2
4 13 15 0 2
15 1 9 7 9 14 1 9 13 1 9 9 0 12 9 2
18 0 9 0 13 3 0 9 1 13 0 9 9 1 12 1 12 9 2
15 1 0 9 0 0 9 7 9 13 3 13 9 1 9 2
10 9 0 9 14 1 9 13 1 9 2
11 13 14 9 2 1 0 3 14 13 9 2
4 9 13 9 2
18 9 13 14 9 2 16 1 0 9 13 15 0 9 1 9 0 9 2
6 7 3 3 13 4 2
8 2 13 14 4 15 13 9 2
3 13 9 2
13 13 15 1 9 2 13 1 0 9 7 13 4 2
13 13 0 9 1 9 9 9 7 9 9 1 9 2
6 9 0 13 9 9 2
15 3 9 13 2 16 1 0 9 9 9 13 12 9 9 2
14 14 1 0 9 1 9 0 1 9 13 14 12 9 2
9 0 9 13 13 1 0 0 9 2
11 0 9 0 13 13 15 1 9 0 9 2
8 2 13 4 15 15 1 9 2
14 9 13 2 16 14 13 13 0 2 13 9 0 9 2
3 9 13 2
3 13 15 2
4 9 13 0 2
7 15 13 9 1 0 9 2
6 2 3 13 3 13 2
12 1 12 9 1 9 9 13 0 9 1 9 2
15 9 13 2 16 9 2 0 14 13 2 14 13 1 9 2
18 9 9 13 14 0 9 2 13 12 9 9 2 13 1 15 12 9 2
15 3 13 9 2 13 9 2 7 1 9 3 13 1 9 2
13 16 13 15 15 13 1 9 2 13 3 0 9 2
9 1 9 13 1 15 0 9 9 2
9 13 0 9 0 1 13 0 9 2
4 9 13 0 2
12 3 0 13 1 0 9 9 7 13 1 9 2
5 9 13 9 9 2
11 9 8 2 13 9 1 12 9 13 9 2
9 13 13 9 1 9 9 0 9 2
12 7 0 1 9 13 15 1 0 9 7 9 2
10 0 9 0 13 15 14 12 9 1 2
5 9 13 1 9 2
17 13 1 9 2 1 0 13 15 9 0 7 3 13 9 1 9 2
9 13 1 9 9 9 0 9 0 2
10 13 9 1 0 9 2 7 9 13 2
13 14 13 14 1 9 13 9 2 16 13 9 0 2
7 1 9 13 9 1 9 2
8 7 3 9 3 13 0 9 2
18 1 0 8 2 9 13 0 9 1 9 1 0 9 13 1 0 9 2
16 9 9 9 0 2 13 1 9 7 9 2 13 9 12 9 2
8 7 1 9 13 13 9 9 2
12 3 9 9 9 9 13 2 16 13 0 9 2
20 1 9 9 13 9 1 9 2 13 15 13 13 1 9 0 9 2 9 9 2
12 1 9 0 9 13 15 0 9 0 1 9 2
8 9 14 13 15 1 0 9 2
8 13 0 9 0 1 9 9 2
3 13 9 2
13 3 13 15 15 9 0 2 0 9 7 0 9 2
11 1 9 13 1 15 0 0 9 7 9 2
15 0 9 13 9 1 13 9 9 1 9 9 8 2 9 2
7 9 9 3 14 4 13 2
7 9 13 1 9 9 9 2
7 13 13 9 1 0 9 2
14 16 9 13 15 1 13 2 9 9 0 7 12 9 2
14 1 9 0 9 4 13 1 0 9 7 13 1 9 2
13 3 0 9 13 9 2 1 0 9 13 9 9 2
6 1 12 9 13 9 2
9 3 0 9 4 14 1 9 13 2
8 9 9 0 13 4 3 13 2
11 13 14 12 9 2 7 0 9 15 13 2
8 3 9 13 1 9 1 9 2
8 9 1 0 9 13 0 9 2
4 12 15 13 2
13 9 0 0 1 9 9 13 9 9 2 9 9 2
5 9 13 14 4 2
9 1 9 9 4 13 1 9 0 2
5 9 4 3 13 2
4 13 12 9 2
14 1 12 9 9 13 13 1 15 1 9 7 9 0 2
5 9 13 15 3 2
9 9 13 1 0 2 1 0 9 2
6 0 9 13 12 9 2
19 13 15 1 12 9 0 9 0 8 2 9 9 14 13 14 13 15 0 2
17 1 9 9 13 1 9 7 9 1 9 13 15 0 7 0 9 2
6 13 14 13 13 9 2
4 0 13 9 2
15 9 0 9 14 12 9 1 13 13 0 9 1 9 9 2
10 9 9 9 13 15 1 9 9 9 2
5 9 13 9 9 2
11 9 9 13 2 16 1 9 13 14 9 2
8 1 9 9 9 15 14 13 2
9 9 13 13 9 9 7 13 15 2
19 12 9 13 9 9 1 9 2 0 13 15 1 9 1 0 9 1 9 2
5 4 13 7 13 2
4 13 14 14 2
9 3 13 9 13 1 15 14 3 2
4 13 15 3 2
10 13 2 16 13 4 15 1 15 3 2
12 9 13 15 1 9 1 9 3 1 9 9 2
16 3 1 8 2 0 3 9 13 1 9 9 1 9 1 9 2
11 14 8 2 8 2 0 3 13 1 9 2
12 9 9 2 9 2 9 7 9 13 13 0 2
21 13 15 9 1 9 2 9 2 0 9 9 2 9 2 9 1 13 2 9 9 2
4 13 9 0 2
3 13 15 2
14 14 13 9 1 9 2 13 14 13 1 12 8 9 2
5 7 9 15 13 2
5 13 1 0 9 2
11 1 0 9 9 13 9 0 9 9 0 2
16 3 1 9 13 9 13 15 12 0 9 1 9 14 12 8 2
9 13 9 1 9 0 9 0 9 2
17 1 9 2 16 9 3 15 14 13 2 13 15 9 0 9 0 2
19 9 9 13 2 16 9 0 9 1 9 0 13 15 1 0 9 0 9 2
8 13 2 16 15 9 4 13 2
5 3 13 1 9 2
4 9 9 13 2
2 13 2
7 13 4 3 1 0 9 2
7 9 2 9 14 13 0 2
4 0 9 13 2
11 0 9 9 9 13 9 9 1 9 9 2
4 13 12 9 2
10 9 14 4 13 1 0 9 1 9 2
9 9 9 13 3 13 0 9 9 2
12 3 9 9 13 15 1 9 9 7 13 9 2
14 9 13 1 9 13 9 1 0 9 14 1 0 8 2
21 9 9 0 13 1 9 9 0 7 0 2 0 13 9 13 1 9 1 9 0 2
11 1 9 9 13 1 9 9 1 9 9 2
7 1 9 13 4 1 9 2
9 13 2 16 0 9 9 15 13 2
7 9 9 9 13 1 9 2
8 2 13 4 1 0 0 9 2
4 2 14 13 2
4 3 15 13 2
6 2 3 2 13 9 2
3 2 13 2
15 9 0 13 3 1 9 7 9 9 13 15 1 13 9 2
3 13 9 2
10 2 9 1 9 13 0 9 1 9 2
15 2 9 13 1 0 9 9 9 7 13 1 0 9 9 2
3 13 13 2
7 13 15 1 9 7 9 2
11 3 9 1 9 1 9 0 9 13 9 2
8 9 13 9 2 16 15 13 2
9 7 9 15 13 1 0 0 9 2
13 13 9 14 1 9 1 9 1 9 1 9 0 2
3 9 13 2
12 0 9 1 9 9 13 15 0 9 9 0 2
8 16 15 0 0 9 13 9 2
23 13 13 15 9 2 16 9 9 13 2 9 13 2 13 2 7 14 3 9 13 2 2 2
5 13 15 1 9 2
5 13 15 0 9 2
5 4 14 4 13 2
15 0 9 13 9 9 2 0 13 3 1 9 1 9 9 2
12 1 9 9 9 13 15 1 9 14 12 9 2
11 15 9 2 9 0 9 2 13 9 9 2
9 3 1 9 1 9 13 9 9 2
5 9 13 4 3 2
18 0 9 13 4 1 9 9 9 1 9 7 0 9 1 9 0 9 2
21 9 14 13 0 9 1 3 13 9 9 9 2 9 14 3 13 1 13 9 9 2
11 14 9 0 9 13 14 4 1 0 9 2
5 13 15 0 9 2
4 9 14 13 2
9 1 0 9 13 0 2 0 9 2
11 13 9 9 2 0 13 1 9 0 9 2
12 1 0 9 0 9 1 9 1 9 14 13 2
14 1 9 9 9 1 9 1 9 13 9 0 9 0 2
13 9 13 12 9 2 9 13 9 0 7 13 9 2
11 9 13 9 1 9 13 1 15 9 0 2
24 0 9 9 13 15 7 13 12 9 1 9 1 9 1 9 9 2 12 8 1 9 1 9 2
17 1 9 9 2 0 13 1 9 9 2 1 9 13 14 9 9 2
9 13 4 9 9 1 0 9 0 2
8 9 0 13 9 12 8 9 2
7 2 13 15 1 9 13 2
5 2 14 13 2 2
7 2 15 7 3 13 2 2
6 13 4 9 1 15 2
10 2 13 2 13 9 1 0 9 2 2
8 9 9 9 13 1 12 9 2
9 9 0 9 0 13 9 12 9 2
19 1 9 13 15 0 9 9 9 1 9 9 9 0 12 9 0 0 9 2
16 9 9 13 9 9 1 9 13 15 9 9 1 9 0 9 2
6 13 9 0 7 0 2
14 0 9 2 0 2 0 7 0 2 13 9 7 9 2
14 1 0 9 9 0 13 15 9 2 1 0 13 13 2
7 0 9 13 1 9 0 2
13 13 0 9 9 2 9 2 9 2 9 2 9 2
21 9 13 9 2 9 2 9 1 15 2 9 2 9 2 13 15 1 9 1 9 2
10 0 0 9 13 15 1 9 0 9 2
13 1 0 9 9 13 15 0 9 1 9 7 9 2
9 13 15 0 9 7 13 0 9 2
6 9 9 14 13 0 2
12 13 14 12 9 2 1 9 1 9 13 9 2
13 9 15 1 9 9 13 2 7 3 0 9 13 2
11 9 13 15 1 9 9 2 13 9 9 2
8 9 13 14 9 1 9 9 2
11 16 3 13 4 15 3 1 0 0 9 2
7 14 13 4 0 0 9 2
6 13 7 13 2 13 2
14 7 0 9 13 2 16 9 0 13 9 0 7 0 2
5 13 4 15 3 2
4 13 13 9 2
15 13 0 0 0 0 9 2 13 1 0 9 1 13 9 2
25 13 15 2 13 1 0 9 9 0 9 2 4 9 2 4 9 2 4 9 2 4 9 2 2 2
10 13 4 2 16 9 14 0 13 0 2
4 13 9 9 2
9 9 0 14 13 14 0 9 9 2
13 9 13 14 9 7 13 14 0 1 0 9 0 2
12 1 0 9 13 3 13 9 9 1 0 9 2
10 1 9 13 9 14 1 0 9 0 2
19 1 9 0 4 3 13 2 16 13 4 0 9 2 0 13 0 9 9 2
4 9 14 13 2
4 13 13 3 2
4 9 13 9 2
8 1 0 9 14 14 13 9 2
7 14 13 1 15 0 9 2
4 13 15 3 2
8 13 1 15 7 13 1 9 2
18 7 9 9 2 14 14 13 2 13 15 9 7 13 1 15 1 9 2
8 1 0 9 13 12 13 9 2
5 14 13 1 15 2
16 12 0 9 13 15 1 9 7 3 13 15 13 1 15 3 2
9 4 13 16 9 0 7 3 0 2
9 14 9 9 14 13 1 15 9 2
14 13 9 7 13 1 9 14 13 14 0 9 0 9 2
12 9 13 15 3 2 16 13 1 0 9 9 2
9 13 14 2 16 9 3 14 13 2
5 13 14 14 3 2
23 9 9 2 9 9 9 9 1 9 9 2 13 1 9 1 9 2 9 7 9 1 9 2
11 9 3 13 0 9 2 1 13 9 9 2
24 3 0 9 13 9 9 2 13 9 7 13 2 0 9 4 0 2 7 14 14 13 0 9 2
7 3 13 1 9 1 9 2
6 2 13 13 1 9 2
8 13 2 16 0 9 14 13 2
6 15 14 13 1 9 2
13 13 7 9 1 9 4 3 3 13 1 9 9 2
12 9 0 9 13 15 1 9 2 0 13 9 2
12 9 0 9 13 15 1 9 2 0 13 9 2
7 9 13 9 1 0 9 2
18 1 9 9 13 2 13 15 1 9 2 7 1 9 3 13 1 15 2
7 13 15 9 1 0 9 2
5 13 15 1 9 2
7 13 1 15 1 0 9 2
4 14 13 3 2
8 13 13 15 1 9 7 9 2
5 1 0 9 13 2
10 2 13 1 9 1 9 1 0 9 2
3 13 9 2
7 2 9 13 9 1 9 2
18 13 4 1 9 7 13 4 2 16 1 9 0 15 9 13 1 9 2
7 9 9 13 1 9 9 2
9 13 15 1 15 2 13 15 0 2
8 1 9 13 2 13 7 13 2
18 1 9 13 1 9 9 2 13 9 13 1 13 9 9 7 13 9 2
6 13 9 13 15 9 2
3 14 13 2
4 9 14 13 2
6 1 9 13 1 9 2
9 0 9 13 4 15 1 0 9 2
8 9 15 13 2 16 13 9 2
7 13 15 7 13 9 9 2
11 13 3 9 1 9 2 16 13 3 13 2
5 2 9 15 13 2
2 13 2
5 1 9 13 4 2
3 2 13 2
8 2 7 9 2 9 15 13 2
18 9 9 13 1 0 9 2 16 0 9 9 13 15 1 15 9 9 2
16 14 13 15 0 9 1 9 0 9 2 7 13 15 9 9 2
8 9 9 13 1 9 9 9 2
16 9 13 0 9 7 13 15 2 16 3 12 4 9 7 9 2
10 14 4 15 9 13 1 9 1 9 2
10 9 13 1 9 8 2 0 13 9 2
14 9 8 2 13 14 9 9 2 0 13 9 1 9 2
10 9 9 7 9 0 9 13 9 0 2
11 9 13 14 9 0 0 9 9 9 9 2
8 1 15 9 13 15 0 9 2
7 13 2 16 9 13 0 2
5 9 9 13 9 2
10 3 1 0 2 12 9 13 1 9 2
11 9 13 15 14 1 0 9 13 9 9 2
12 9 9 13 3 1 9 1 9 0 9 0 2
6 3 13 9 0 9 2
9 1 13 9 9 0 14 13 9 2
8 14 13 9 0 9 9 9 2
8 1 0 9 9 13 14 9 2
4 14 13 3 2
19 2 13 9 15 9 9 9 2 9 7 9 1 9 9 0 1 12 9 2
12 7 14 9 14 13 15 13 1 0 9 0 2
10 0 9 0 13 1 9 12 0 9 2
11 1 9 13 14 9 13 15 1 0 9 2
7 3 9 9 13 0 9 2
10 1 9 13 15 1 9 1 13 9 2
4 14 13 9 2
15 1 9 13 9 2 9 0 3 14 13 1 9 9 0 2
5 3 15 14 13 2
13 14 12 9 1 12 9 1 0 9 13 1 9 2
9 3 13 15 13 1 8 2 0 2
7 0 9 13 9 7 9 2
10 0 9 13 9 13 1 9 9 0 2
16 9 13 15 13 9 0 1 9 13 2 0 14 13 0 9 2
6 2 9 13 12 9 2
12 14 14 3 13 15 2 16 14 9 14 13 2
5 13 13 0 9 2
11 9 13 0 9 9 14 13 14 1 9 2
7 3 9 13 15 1 9 2
7 13 0 9 1 9 0 2
3 14 13 2
2 13 2
13 9 1 9 0 13 2 16 13 9 1 9 9 2
13 9 9 7 9 1 9 0 9 13 1 12 8 2
5 0 13 14 9 2
3 9 13 2
11 3 3 0 9 13 4 1 9 0 8 2
4 13 0 9 2
10 9 9 13 1 9 1 9 12 9 2
9 1 0 9 9 13 1 13 9 2
20 0 9 1 9 9 13 13 9 1 9 1 9 1 9 0 9 0 1 9 2
15 9 7 9 13 2 16 3 9 9 9 7 9 3 13 2
7 13 14 0 9 1 9 2
13 9 7 9 13 1 9 13 1 0 9 0 9 2
22 1 9 9 1 9 0 2 0 9 13 9 2 9 13 3 0 9 9 0 2 0 2
17 0 9 0 0 9 1 0 9 13 1 9 1 0 9 0 9 2
16 9 3 13 15 1 0 9 2 7 9 9 13 15 1 9 2
7 2 14 9 15 14 13 2
11 1 0 9 9 3 13 7 13 1 9 2
16 13 9 13 0 9 9 0 2 0 9 7 9 9 9 0 2
18 13 3 9 0 9 0 2 13 9 9 1 9 9 0 2 13 9 2
15 2 13 4 14 9 9 1 9 2 0 15 9 14 13 2
21 14 9 0 0 9 0 13 2 16 9 13 9 2 16 13 1 9 9 1 9 2
8 2 9 14 13 13 9 9 2
8 9 13 13 1 9 9 9 2
7 9 9 0 13 12 9 2
8 4 13 7 0 9 0 9 2
5 9 14 14 13 2
8 2 9 14 13 9 1 9 2
9 13 1 9 2 16 3 13 9 2
5 9 9 13 0 2
14 14 13 4 9 1 9 1 9 9 13 1 9 9 2
5 13 9 1 9 2
10 1 9 0 9 13 0 1 9 9 2
8 13 4 3 3 0 9 9 2
9 3 14 14 13 4 0 9 9 2
8 0 9 9 13 14 0 9 2
21 0 9 0 13 12 9 2 7 9 2 9 0 9 1 9 2 13 1 12 9 2
11 2 14 9 9 13 9 0 1 9 0 2
12 15 15 14 13 2 16 13 3 0 1 9 2
9 2 15 14 13 15 1 0 9 2
7 2 13 14 0 1 9 2
7 2 9 13 1 0 9 2
23 14 13 1 9 9 2 9 9 13 13 1 9 9 9 2 9 7 9 13 1 9 9 2
8 1 9 1 15 9 15 13 2
6 0 9 9 13 3 2
7 14 13 15 15 13 9 2
14 1 9 9 9 13 15 13 1 9 1 12 0 9 2
9 3 1 0 9 3 13 15 3 2
15 9 13 9 0 2 0 9 9 2 9 0 0 9 9 2
6 9 9 13 1 9 2
15 13 1 9 9 1 9 1 9 0 8 2 13 3 0 2
10 13 15 14 0 9 9 9 9 9 2
6 1 9 13 9 9 2
11 2 13 13 2 9 13 1 9 9 0 2
11 2 14 14 13 9 0 1 13 0 9 2
8 2 7 9 9 13 1 9 2
5 1 13 13 9 2
7 9 14 13 15 1 9 2
18 0 9 14 13 2 7 0 9 1 0 9 0 9 13 14 9 9 2
17 9 9 9 9 7 9 9 9 9 3 4 13 1 13 0 9 2
8 9 0 9 13 15 3 3 2
10 9 0 9 1 0 9 13 9 0 2
21 14 1 9 13 9 0 0 9 14 13 2 14 9 9 13 0 9 1 15 9 2
14 9 13 0 9 7 3 13 13 15 9 9 0 9 2
8 2 9 13 0 9 1 9 2
15 2 3 9 0 13 1 9 9 1 9 9 1 9 9 2
4 14 9 13 2
6 14 13 14 9 0 2
11 3 14 14 13 2 0 9 13 1 9 2
8 0 9 13 14 9 0 9 2
15 9 1 9 9 0 13 3 2 16 9 0 9 13 0 2
11 3 1 9 9 13 15 1 9 7 9 2
13 1 9 9 13 14 1 9 9 1 0 9 0 2
15 13 16 9 9 0 14 13 13 9 1 9 1 0 9 2
10 9 14 13 0 9 1 0 13 9 2
11 0 9 4 9 13 1 9 0 9 0 2
14 9 13 1 0 9 2 0 13 14 9 9 9 0 2
13 14 13 0 9 9 2 14 13 0 9 9 9 2
10 1 0 8 2 9 1 9 4 13 2
3 9 13 2
17 9 0 9 9 9 13 13 2 16 9 13 9 9 14 13 9 2
7 2 0 9 13 9 9 2
4 13 1 9 2
8 9 0 9 4 13 1 9 2
15 1 9 14 13 2 16 9 13 13 2 16 13 0 9 2
11 13 9 12 0 9 9 9 0 1 9 2
6 12 9 9 13 9 2
6 12 9 13 1 9 2
10 1 9 1 9 0 13 3 12 9 2
6 1 9 13 1 9 2
15 9 9 1 0 12 9 3 13 0 9 1 0 9 9 2
18 9 14 13 13 1 9 2 0 13 2 0 9 2 9 7 0 9 2
17 2 0 9 9 13 1 9 9 0 7 0 9 9 1 9 2 2
11 14 13 14 13 9 9 1 9 0 9 2
17 13 14 9 0 9 2 13 0 9 9 7 13 9 9 7 9 2
8 13 1 13 9 7 0 9 2
6 13 9 0 9 0 2
8 13 15 0 9 9 0 9 2
4 9 13 9 2
11 13 15 13 0 9 2 9 1 0 9 2
17 1 9 1 9 13 15 13 1 9 2 16 9 3 1 15 13 2
6 14 14 13 3 3 2
14 13 15 2 16 9 13 2 7 15 14 13 1 9 2
7 14 13 14 9 1 9 2
15 13 2 16 9 1 9 13 2 7 15 14 13 2 2 2
8 9 13 1 9 2 7 13 2
13 14 13 14 2 3 13 9 7 3 13 0 9 2
6 0 9 13 0 9 2
9 13 15 14 9 9 0 1 9 2
6 13 4 1 9 3 2
9 14 13 9 0 0 9 1 9 2
14 1 9 13 9 0 1 13 9 1 9 13 9 9 2
13 14 13 15 1 9 9 0 2 16 1 15 13 2
18 1 0 9 9 9 13 1 13 0 9 2 0 1 0 9 1 9 2
12 1 9 9 9 13 9 2 16 13 3 13 2
13 1 9 9 9 9 0 13 3 0 2 0 9 2
10 14 3 13 2 14 14 13 1 9 2
6 0 9 14 13 9 2
4 13 3 9 2
12 9 2 3 13 9 1 0 14 13 0 9 2
9 13 9 9 9 9 1 0 9 2
14 9 9 13 15 1 9 2 13 1 9 1 0 9 2
15 0 0 9 9 4 1 9 13 1 9 9 9 9 0 2
13 1 9 0 9 13 9 0 2 7 13 15 9 2
10 3 13 15 15 1 13 9 1 9 2
6 3 1 9 9 13 2
22 1 12 1 12 13 15 1 9 9 9 2 13 9 13 1 9 1 0 9 7 9 2
16 1 0 14 9 0 1 3 12 9 1 15 4 1 9 13 2
6 2 3 14 13 9 2
12 7 9 0 13 3 0 7 0 1 9 0 2
8 14 13 15 1 9 9 0 2
13 2 0 13 9 0 9 2 0 9 13 1 9 2
7 2 12 9 13 9 0 2
6 2 9 9 9 13 2
14 3 1 9 14 13 0 9 7 14 13 0 9 0 2
20 1 9 0 9 2 1 12 9 2 9 4 13 1 9 1 9 1 9 0 2
5 1 9 13 9 2
8 1 9 0 3 9 13 9 2
7 1 12 9 9 13 0 2
11 16 9 15 13 2 13 9 1 13 9 2
10 12 9 1 0 9 0 15 14 13 2
9 3 1 9 9 13 4 9 0 2
6 2 13 1 9 0 2
11 16 9 13 2 4 13 0 9 1 9 2
6 13 9 1 0 9 2
9 1 9 0 13 9 9 9 9 2
19 7 15 2 7 9 9 9 14 13 14 13 15 1 0 9 1 9 9 2
3 9 13 2
6 4 13 1 9 9 2
6 4 14 13 1 9 2
10 1 0 9 13 1 9 0 1 9 2
12 9 9 13 3 1 9 7 13 1 9 9 2
8 13 1 12 8 9 7 9 2
5 3 13 9 0 2
17 9 0 13 9 1 0 9 1 0 0 9 9 2 14 3 13 2
10 1 9 4 13 9 1 9 1 13 2
7 7 9 9 9 4 13 2
7 0 0 9 13 1 9 2
17 1 9 9 1 13 9 13 1 9 2 1 0 0 9 1 9 2
17 9 13 3 1 0 2 12 2 7 0 9 13 9 1 9 9 2
11 0 9 13 9 0 2 9 9 7 9 2
6 9 13 13 1 9 2
5 13 14 1 9 2
5 9 14 13 9 2
17 1 9 9 3 13 9 9 9 2 9 1 9 0 1 9 9 2
12 16 3 9 13 1 15 0 9 1 0 9 2
5 3 3 15 13 2
8 13 2 16 13 15 0 9 2
10 9 9 14 13 2 7 13 1 9 2
17 9 13 1 9 9 2 1 0 9 9 13 15 1 9 13 9 2
8 9 0 14 13 13 12 9 2
10 13 9 1 9 14 13 13 13 9 2
8 9 13 4 13 1 9 0 2
7 13 9 0 9 0 9 2
7 13 9 14 9 0 9 2
3 13 9 2
8 9 13 15 13 1 0 9 2
15 13 14 9 2 16 9 9 3 3 13 14 13 0 9 2
6 13 13 1 0 9 2
8 9 0 13 15 1 0 9 2
7 3 13 2 16 13 0 2
3 14 13 2
4 9 14 13 2
14 9 13 9 2 16 9 14 13 9 2 16 15 13 2
11 13 14 4 13 15 12 9 1 9 9 2
11 13 4 1 9 2 0 9 13 0 9 2
22 16 9 9 13 15 1 9 7 9 2 7 9 0 9 13 14 12 8 2 0 9 2
20 4 13 9 2 7 0 9 3 13 2 1 15 14 2 13 14 9 0 9 2
8 13 1 15 0 9 1 9 2
11 3 13 14 1 9 0 9 1 9 0 2
14 9 1 9 13 1 12 9 1 9 9 13 1 9 2
6 7 3 14 4 13 2
6 9 15 1 9 13 2
3 9 13 2
7 9 9 13 14 1 9 2
10 1 9 0 13 4 14 12 13 9 2
10 9 0 13 13 9 1 12 9 9 2
6 9 3 13 15 9 2
11 14 9 2 1 9 2 13 0 9 0 2
5 13 15 14 9 2
14 0 1 0 9 9 13 15 1 9 1 9 1 9 2
9 7 3 13 15 2 13 0 9 2
25 1 9 13 0 9 2 9 13 9 0 9 7 13 15 9 1 0 9 7 9 2 0 3 13 2
8 0 9 13 0 9 0 9 2
4 1 9 13 2
15 3 9 4 13 7 9 13 1 9 2 7 14 9 9 2
30 7 3 13 4 15 2 16 14 13 14 13 1 9 13 1 9 1 9 9 2 16 1 9 0 9 9 13 15 9 2
9 2 9 13 4 1 9 2 2 2
15 2 7 1 9 9 1 0 9 0 13 15 12 0 9 2
14 9 9 13 2 16 0 9 14 13 3 3 1 9 2
3 2 13 2
9 14 14 13 9 1 9 0 9 2
15 2 3 13 9 2 16 9 13 15 1 9 9 1 9 2
8 13 15 9 2 16 13 9 2
11 9 13 12 9 9 9 7 9 9 9 2
9 1 0 9 9 9 13 9 9 2
13 9 9 13 1 9 9 14 9 1 0 2 9 2
12 16 13 9 2 9 13 9 1 9 7 13 2
24 13 2 16 0 9 0 8 2 9 0 3 9 13 15 1 0 9 1 9 9 2 9 9 2
14 2 13 13 9 2 0 13 13 13 1 0 9 9 2
6 9 0 14 13 0 2
12 7 0 9 1 9 14 13 13 0 9 0 2
3 14 13 2
6 14 13 1 9 9 2
12 7 14 13 13 2 13 2 16 9 14 13 2
7 2 3 1 9 14 13 2
8 2 3 13 4 13 1 9 2
6 14 9 15 14 13 2
8 14 1 9 13 1 9 0 2
21 9 14 12 9 0 2 9 7 9 1 12 0 9 13 13 0 9 13 9 0 2
17 16 13 13 1 9 0 9 0 9 0 2 0 13 0 13 9 2
8 9 13 9 7 13 1 9 2
7 2 13 0 9 1 9 2
3 9 13 2
5 13 15 0 9 2
9 1 9 13 14 1 9 9 0 2
16 9 9 13 1 9 1 0 9 9 0 2 0 13 9 9 2
10 3 9 1 0 12 9 1 9 13 2
6 1 9 13 15 9 2
13 13 15 1 9 9 0 1 9 13 1 9 9 2
9 14 9 13 2 16 9 13 0 2
11 2 3 9 13 0 9 0 9 1 9 2
8 9 13 14 9 13 3 9 2
10 13 9 9 0 0 3 9 1 9 2
7 3 13 0 1 9 9 2
7 7 3 13 9 0 9 2
14 13 15 9 2 16 0 9 0 13 0 9 1 9 2
6 9 13 9 1 9 2
7 0 9 13 4 0 9 2
18 9 9 2 0 1 9 13 9 13 9 0 2 13 0 9 9 9 2
20 16 4 15 13 2 7 1 12 9 4 13 1 9 8 2 12 9 9 0 2
8 0 9 13 14 0 0 9 2
18 9 0 13 13 9 1 9 1 9 2 16 9 0 13 15 1 9 2
14 13 2 14 13 14 3 0 9 2 16 0 13 9 2
8 2 1 0 9 4 0 9 2
9 3 14 13 9 0 1 15 9 2
3 13 9 2
25 14 13 1 9 0 2 13 4 1 0 9 9 2 0 0 9 13 9 13 9 13 1 9 9 2
3 9 13 2
4 13 9 0 2
11 9 13 9 13 0 9 13 1 0 9 2
6 9 13 15 1 9 2
12 3 13 2 16 13 9 0 9 13 1 9 2
17 9 9 13 13 9 3 2 0 9 13 15 7 13 1 0 9 2
6 3 13 15 1 9 2
13 9 13 1 0 9 2 7 15 14 13 9 13 2
9 9 9 13 1 9 9 1 9 2
5 9 9 13 0 2
8 1 9 9 13 15 9 9 2
7 13 13 9 1 0 9 2
18 1 0 9 9 13 2 16 15 0 1 9 9 13 0 7 13 0 2
5 3 13 0 9 2
7 1 12 9 13 9 0 2
5 13 14 9 0 2
6 1 12 9 13 9 2
6 13 1 9 1 9 2
6 13 1 0 9 9 2
6 9 3 13 7 13 2
17 9 13 15 1 9 2 16 13 1 0 9 7 13 15 1 9 2
12 16 9 13 0 9 2 14 14 1 15 13 2
13 2 1 9 0 9 14 13 0 9 1 9 9 2
8 2 1 9 14 13 0 9 2
12 13 1 9 1 9 9 1 9 13 1 9 2
12 9 1 9 9 7 9 13 8 2 9 9 2
14 1 0 9 13 0 9 9 4 12 0 9 0 9 2
17 1 9 7 13 9 13 4 12 8 2 9 7 12 8 2 9 2
11 9 13 4 12 8 2 9 7 9 0 2
11 3 0 13 9 2 9 2 9 7 9 2
11 9 13 1 9 2 9 2 9 7 9 2
16 3 1 9 9 9 0 1 0 1 9 9 13 9 13 9 2
11 9 13 2 16 9 13 0 1 15 9 2
9 12 9 9 13 9 12 9 9 2
13 1 9 1 9 13 9 1 0 9 9 9 9 2
15 13 15 9 1 3 0 9 9 1 9 9 7 0 9 2
18 0 1 9 9 0 0 9 0 13 3 0 0 9 9 13 12 9 2
13 1 9 9 0 9 9 0 13 9 1 0 9 2
7 1 9 13 0 9 9 2
22 9 9 9 9 2 0 9 9 9 7 9 9 9 9 9 13 1 9 9 9 9 2
10 9 13 15 7 13 9 1 0 9 2
8 3 13 9 1 9 9 9 2
12 9 0 13 3 2 16 13 9 9 1 9 2
7 4 15 13 1 0 9 2
12 3 13 1 9 2 13 14 3 0 9 9 2
6 15 13 3 0 9 2
14 9 8 2 14 13 0 0 9 2 0 13 15 9 2
5 9 14 13 15 2
6 9 13 7 9 0 2
7 9 13 14 1 12 9 2
11 9 1 9 14 13 13 1 13 9 9 2
12 9 0 1 9 9 1 0 13 1 0 9 2
8 2 1 9 14 13 4 9 2
12 13 15 9 2 14 0 9 13 15 9 9 2
12 2 13 4 2 16 13 4 15 3 3 13 2
15 14 13 13 0 2 16 1 9 13 4 9 1 0 9 2
9 13 1 0 9 2 0 15 13 2
11 2 13 4 2 16 13 9 14 0 9 2
8 2 9 14 13 1 9 0 2
8 2 13 3 9 0 9 0 2
6 13 15 9 9 9 2
19 13 15 15 2 16 4 13 0 1 0 9 9 2 1 0 9 14 13 2
12 14 13 15 15 2 16 13 4 9 9 9 2
13 14 13 2 14 13 9 13 0 9 1 15 9 2
9 13 15 9 0 13 9 0 9 2
12 9 13 1 3 12 9 1 13 9 1 9 2
21 3 13 15 9 9 0 2 7 3 0 1 15 4 13 13 9 1 9 2 9 2
11 7 9 0 13 2 16 13 1 9 9 2
19 7 3 9 13 14 1 9 2 9 2 9 2 13 14 9 7 9 0 2
8 0 9 13 4 14 12 9 2
12 9 0 1 9 13 9 7 13 3 0 9 2
17 1 0 9 9 13 13 1 9 2 3 13 15 13 1 15 9 2
10 3 13 15 9 9 9 7 0 9 2
27 9 1 9 1 0 9 13 4 14 13 0 9 7 13 0 9 2 7 3 13 4 9 0 9 9 9 2
7 9 14 4 13 12 9 2
19 9 9 13 9 0 9 2 13 9 1 9 2 7 1 9 13 15 9 2
9 1 0 9 1 9 13 3 9 2
15 1 9 9 9 13 1 9 9 2 7 9 13 13 0 2
16 9 13 13 0 9 0 9 7 3 13 1 9 9 1 9 2
8 1 9 9 13 1 0 9 2
4 1 9 13 2
9 16 15 14 13 2 13 3 0 2
16 9 13 2 16 1 9 9 13 1 0 12 9 12 0 9 2
14 9 7 9 2 0 13 2 13 14 2 16 9 13 2
11 14 1 12 9 1 9 13 15 9 9 2
10 2 7 15 9 1 9 4 3 13 2
7 14 14 13 7 14 3 2
7 1 9 9 13 9 9 2
7 1 0 0 14 13 9 2
19 14 2 0 13 9 2 0 13 14 14 0 9 2 9 9 2 0 9 2
6 14 13 3 13 9 2
19 1 9 0 0 8 2 1 0 0 9 0 13 4 3 0 0 9 0 2
5 13 4 9 9 2
7 9 9 1 9 15 13 2
6 13 15 13 1 9 2
6 1 9 9 13 9 2
6 2 13 7 1 9 2
17 14 13 0 9 1 0 9 2 7 14 13 0 9 9 1 9 2
27 1 0 9 13 2 16 1 12 9 2 0 13 1 9 1 9 0 1 9 0 2 9 13 9 0 9 2
19 1 13 3 1 9 9 9 13 12 9 1 12 0 9 9 9 9 9 2
14 0 9 13 0 13 1 9 9 9 1 9 0 9 2
16 9 13 0 9 2 7 1 0 9 12 9 1 9 13 9 2
5 3 3 13 9 2
10 2 0 9 13 0 9 9 1 9 2
9 13 14 9 7 0 9 13 9 2
5 14 9 13 9 2
4 13 1 9 2
5 13 9 0 9 2
15 9 9 9 14 13 1 15 9 1 13 13 15 0 9 2
10 1 9 13 4 1 13 0 9 0 2
19 13 14 15 13 9 0 2 0 13 9 1 13 9 1 9 0 7 0 2
10 3 13 0 9 2 9 13 9 9 2
8 3 13 9 1 9 0 9 2
4 0 14 13 2
15 13 9 2 16 8 2 12 1 12 9 13 13 15 9 2
16 2 9 2 3 13 4 2 16 15 13 0 9 7 0 9 2
6 2 3 15 13 4 2
12 2 7 14 3 13 4 1 9 9 3 3 2
8 0 9 9 9 13 1 9 2
13 9 13 2 16 1 12 9 0 9 13 0 9 2
9 9 13 14 1 9 0 9 9 2
13 0 9 2 0 13 0 9 2 9 13 3 3 2
13 9 1 9 2 0 13 9 0 2 13 14 13 2
15 9 1 9 0 4 13 14 2 3 1 9 13 0 9 2
15 1 0 9 1 9 9 0 13 14 15 12 9 14 9 2
9 0 13 14 9 12 9 1 9 2
10 14 13 13 3 2 16 9 13 0 2
8 2 13 4 0 9 9 0 2
13 9 13 2 16 9 1 9 14 13 0 9 9 2
10 1 9 13 4 15 13 1 9 9 2
6 9 13 15 1 9 2
4 9 14 13 2
19 2 13 15 2 16 13 4 0 9 1 9 2 7 9 14 13 9 9 2
24 3 13 9 13 1 9 0 1 9 7 9 2 9 13 0 9 13 9 1 9 0 9 9 2
6 1 0 9 13 9 2
9 9 0 13 9 0 9 0 9 2
7 13 13 13 15 1 9 2
8 7 14 4 13 9 1 9 2
24 13 15 14 13 2 16 9 13 9 2 0 1 9 13 9 0 9 2 7 13 15 0 9 2
25 1 13 3 9 9 13 2 16 13 13 9 2 16 3 13 15 9 9 2 13 9 9 1 9 2
10 2 0 9 13 9 14 12 9 1 2
14 9 9 13 2 16 13 3 1 9 9 1 9 9 2
14 9 13 9 0 13 9 0 7 13 15 1 0 9 2
4 9 9 13 2
17 0 9 1 9 13 9 0 9 1 13 9 0 2 7 14 9 2
7 9 13 9 1 9 9 2
6 14 4 13 7 13 2
4 14 13 15 2
13 0 1 0 9 9 13 14 0 9 1 9 0 2
11 13 15 9 9 7 3 0 7 0 9 2
8 3 13 4 9 1 9 9 2
11 13 9 9 9 1 0 9 1 9 9 2
13 3 9 1 9 14 3 13 0 13 9 1 9 2
7 9 0 9 14 13 13 2
7 9 13 2 9 13 9 2
5 13 9 9 9 2
7 13 15 0 9 7 9 2
14 2 9 0 13 2 7 8 2 3 13 15 1 9 2
13 9 13 2 16 0 9 4 13 1 13 0 9 2
16 16 9 13 9 2 13 9 2 16 14 13 0 9 1 9 2
4 9 14 13 2
16 14 1 12 9 9 9 13 14 0 2 13 15 15 3 3 2
11 9 1 9 13 9 2 14 13 15 9 2
12 3 13 9 1 9 0 0 9 1 0 9 2
5 9 3 13 9 2
4 13 15 9 2
27 9 9 2 0 7 0 2 3 13 9 7 9 1 0 9 2 13 3 9 0 9 2 9 7 9 9 2
32 2 13 2 16 9 1 9 1 9 0 13 0 9 0 9 7 9 0 2 13 1 9 9 1 9 9 7 0 9 1 9 2
10 9 13 2 16 1 9 13 15 9 2
10 0 9 14 13 9 1 0 9 0 2
9 8 2 9 13 9 0 9 0 2
19 1 9 1 0 9 3 13 15 9 13 3 9 2 9 9 0 7 9 2
16 14 9 13 2 16 1 0 8 2 14 13 4 3 1 9 2
11 14 13 15 1 9 2 14 13 15 9 2
23 3 13 2 13 0 9 1 9 7 13 0 9 1 9 2 3 14 13 15 1 0 9 2
4 9 13 9 2
13 14 3 13 15 2 16 0 9 9 13 1 9 2
14 1 0 1 9 2 9 7 9 9 9 13 15 9 2
5 13 15 1 9 2
3 13 13 2
7 1 9 13 9 1 9 2
4 3 0 13 2
10 1 0 9 13 1 9 0 9 0 2
5 13 1 9 0 2
16 13 15 9 0 2 9 0 7 13 2 16 9 13 0 9 2
8 2 14 13 14 13 0 9 2
8 2 0 2 9 13 1 9 2
21 14 13 15 1 9 1 9 9 9 9 2 7 3 14 0 9 13 1 9 0 2
16 3 14 13 13 15 0 9 2 3 9 1 0 14 4 13 2
5 13 1 0 9 2
5 13 1 15 0 2
9 1 9 13 14 12 0 9 3 2
17 14 9 1 0 9 9 13 0 1 9 2 14 13 14 9 9 2
14 2 3 13 15 1 9 9 1 9 0 1 9 9 2
7 2 14 13 9 0 9 2
15 3 14 4 9 9 9 0 2 9 1 9 1 9 0 2
26 9 14 9 4 15 13 1 9 0 9 0 2 1 0 9 0 13 15 1 9 0 7 9 0 9 2
11 3 4 13 7 9 0 1 9 9 0 2
14 13 4 2 16 4 13 2 13 4 9 1 9 0 2
7 2 3 13 4 1 9 2
13 3 13 2 16 0 9 13 14 13 1 9 9 2
12 0 0 9 13 9 2 7 9 14 13 9 2
13 7 1 15 14 13 9 1 9 2 9 7 9 2
6 2 0 9 13 9 2
16 2 1 13 1 9 9 7 9 9 14 4 15 3 13 3 2
13 1 0 9 0 9 9 4 13 13 0 9 0 2
12 9 13 1 9 9 2 7 9 13 15 13 2
6 9 14 13 13 9 2
15 16 14 13 0 9 2 9 13 13 15 1 9 1 9 2
6 13 9 9 7 9 2
5 13 9 9 9 2
7 0 9 13 0 9 9 2
22 9 13 3 0 2 16 13 15 1 9 9 2 7 14 13 13 1 15 13 2 2 2
15 14 1 8 2 13 9 1 0 9 9 13 13 1 9 2
11 0 0 9 13 9 1 9 9 13 9 2
12 3 0 9 9 13 1 9 13 13 0 9 2
8 12 0 9 13 9 13 9 2
12 2 13 7 1 9 13 2 16 0 9 13 2
5 9 14 13 9 2
15 2 1 0 9 3 15 15 13 2 16 3 12 9 13 2
16 14 0 9 9 1 0 9 4 13 1 9 9 1 0 9 2
9 7 13 0 9 1 13 1 9 2
12 9 13 13 1 9 0 9 14 12 8 8 2
8 1 12 9 13 4 0 9 2
20 1 12 9 1 9 13 15 3 9 0 9 0 1 9 9 0 9 0 8 2
8 1 0 9 9 14 14 13 2
7 13 2 7 13 2 2 2
18 13 9 12 8 2 9 9 7 13 0 1 12 9 9 13 1 9 2
18 1 0 0 9 0 9 9 13 3 9 9 9 7 9 9 7 9 2
15 13 9 2 0 4 1 9 13 1 13 2 3 13 13 2
8 9 9 14 13 15 1 9 2
4 13 15 9 2
18 14 13 9 9 9 1 9 1 9 2 3 13 15 1 13 1 9 2
10 1 9 13 15 3 1 9 9 9 2
8 9 13 2 14 13 13 9 2
8 13 4 14 1 9 1 9 2
5 13 1 9 9 2
10 13 9 1 9 2 13 3 0 9 2
18 0 9 13 1 9 1 9 9 1 9 9 2 3 13 12 0 9 2
14 3 2 16 13 15 13 1 9 2 4 13 1 9 2
8 13 0 9 1 9 9 9 2
11 9 0 1 9 3 13 13 15 9 0 2
9 9 13 12 9 1 13 0 9 2
8 13 13 4 13 1 9 9 2
8 9 13 1 9 9 0 9 2
10 9 1 9 13 1 0 9 9 0 2
10 13 1 9 7 13 1 9 0 9 2
8 1 9 13 9 9 0 9 2
16 9 0 9 13 13 1 9 9 9 7 9 0 9 0 9 2
9 9 0 1 9 13 9 9 9 2
16 9 13 9 9 2 7 13 1 0 8 2 9 7 9 9 2
8 2 14 2 13 14 9 9 2
24 1 9 9 13 15 3 1 9 9 1 9 0 2 13 9 0 7 14 13 15 3 1 9 2
19 13 2 16 13 4 1 0 2 12 1 9 2 13 15 1 9 9 0 2
4 2 13 15 2
11 13 2 16 3 0 9 13 9 9 0 2
11 13 15 0 9 2 9 7 0 9 0 2
10 1 0 9 9 13 1 9 0 9 2
9 16 13 9 9 2 13 13 9 2
4 14 2 13 2
16 13 4 15 9 7 13 15 2 16 13 4 14 14 12 9 2
7 14 9 9 15 14 13 2
16 9 14 13 1 3 2 1 16 13 3 9 13 15 9 0 2
14 14 0 9 13 2 16 9 14 13 9 1 9 9 2
6 1 9 13 0 9 2
8 14 3 13 2 16 9 13 2
15 3 13 9 0 1 9 2 9 2 9 2 9 2 9 2
6 0 9 13 13 9 2
15 16 13 2 13 0 9 2 13 0 9 1 9 13 9 2
9 9 9 7 9 13 1 0 9 2
12 9 0 13 0 9 2 7 14 13 0 9 2
12 0 9 7 9 0 9 9 13 3 0 9 2
7 1 9 13 14 12 9 2
9 3 13 1 15 9 0 9 9 2
10 9 1 9 13 0 9 13 1 9 2
10 13 15 3 0 9 1 13 15 9 2
7 9 13 15 1 9 0 2
5 13 4 14 9 2
15 1 9 13 1 9 2 0 13 9 2 13 1 9 9 2
7 13 15 3 13 14 9 2
15 1 15 1 9 12 8 13 9 13 1 12 9 7 9 2
13 13 4 1 9 7 3 13 4 15 9 1 9 2
7 3 9 13 1 0 9 2
11 9 1 9 13 1 15 9 1 0 9 2
3 13 4 2
4 9 13 3 2
13 13 4 9 1 0 9 7 13 4 0 9 9 2
7 3 13 0 9 7 13 2
4 2 14 13 2
6 2 13 4 1 15 2
5 2 13 1 9 2
5 13 4 1 15 2
4 2 13 15 2
4 2 13 9 2
7 2 1 9 15 3 13 2
11 13 15 13 1 0 9 13 1 0 9 2
9 0 9 13 15 3 0 2 2 2
6 3 13 4 1 9 2
4 13 14 9 2
15 12 9 13 4 1 9 1 9 2 1 0 4 13 13 2
19 7 0 9 13 0 9 2 0 13 1 9 0 2 16 3 13 3 9 2
7 1 9 0 13 9 0 2
10 13 0 2 0 9 13 9 9 0 2
11 13 15 0 9 7 9 15 9 13 0 2
12 9 13 15 0 9 1 0 9 7 0 9 2
6 3 14 13 0 9 2
11 13 1 9 1 12 9 1 9 9 0 2
16 9 0 9 13 9 7 14 13 2 9 13 15 1 0 9 2
12 1 0 9 9 0 9 2 9 13 0 9 2
18 9 8 2 13 15 1 13 15 9 7 1 9 0 3 13 1 9 2
20 12 0 9 13 1 0 2 0 9 9 1 9 1 9 9 9 0 7 0 2
16 0 9 1 0 9 2 0 13 0 9 2 13 15 3 3 2
12 0 9 1 0 9 13 3 1 9 0 9 2
10 1 9 7 0 9 13 14 9 0 2
8 9 0 9 13 15 1 9 2
11 1 9 3 9 0 13 15 1 0 9 2
13 9 13 2 16 9 1 9 9 14 13 12 9 2
17 9 1 9 12 9 9 13 9 1 9 0 9 9 0 1 9 2
9 1 9 9 9 13 12 8 9 2
10 2 1 9 0 3 13 1 9 0 2
9 2 1 0 14 9 3 9 13 2
6 2 14 13 9 9 2
6 2 3 3 9 13 2
12 13 13 9 1 9 1 0 9 7 0 9 2
16 0 9 13 7 9 13 2 9 0 1 9 9 13 2 2 2
8 1 13 9 14 13 0 9 2
6 13 0 9 9 13 2
9 9 13 15 14 3 1 9 9 2
9 4 13 9 14 0 7 3 0 2
10 14 0 9 9 13 15 1 0 9 2
27 13 14 1 13 9 2 3 9 2 13 1 9 1 13 9 7 9 1 9 2 14 13 1 9 1 9 2
3 14 13 2
8 9 3 14 15 13 1 9 2
7 0 9 13 3 1 9 2
18 2 13 9 2 7 15 15 13 2 16 1 0 9 13 15 1 9 2
7 9 13 2 13 9 9 2
6 2 9 3 13 13 2
7 2 13 14 4 13 9 2
6 13 3 7 13 9 2
7 9 1 9 13 15 9 2
11 2 13 2 7 1 9 9 13 9 13 2
5 9 13 3 0 2
5 2 13 1 9 2
4 9 13 9 2
3 2 13 2
6 7 9 14 13 0 2
8 3 13 14 13 15 0 9 2
10 13 7 7 13 9 2 13 0 9 2
13 2 14 13 2 14 13 9 7 14 13 1 9 2
2 13 2
10 2 13 0 7 14 13 15 1 9 2
5 3 9 15 13 2
6 2 9 13 1 9 2
5 2 14 13 4 2
3 2 13 2
8 2 13 1 9 13 2 13 2
6 9 13 15 1 9 2
3 13 9 2
7 2 14 3 13 15 3 2
6 2 7 15 13 9 2
8 14 1 9 13 15 1 9 2
3 13 15 2
3 13 15 2
5 2 4 15 13 2
8 2 13 1 15 2 13 15 2
9 9 1 9 13 9 1 13 9 2
10 13 15 2 16 12 9 13 0 9 2
5 2 14 13 9 2
9 1 13 9 15 15 1 9 13 2
5 13 4 1 9 2
6 13 4 9 1 9 2
5 3 13 0 9 2
5 13 13 1 9 2
4 13 4 9 2
29 9 13 0 1 0 9 0 9 7 13 0 9 2 1 9 2 9 2 0 9 7 9 2 1 9 0 0 9 2
8 1 9 13 14 9 9 0 2
13 13 14 0 9 1 9 0 2 1 9 7 9 2
20 0 9 1 0 9 13 2 13 2 13 9 0 7 13 9 1 12 9 13 2
15 9 13 9 2 13 9 2 13 15 1 9 7 13 9 2
7 14 13 3 9 1 9 2
11 1 12 9 9 14 13 2 13 0 13 2
15 1 9 13 9 1 0 1 9 9 2 0 13 12 9 2
11 13 14 9 1 9 9 13 1 9 9 2
6 2 7 13 4 9 2
4 12 14 13 2
13 13 9 1 9 2 16 9 13 14 1 9 9 2
5 3 13 1 15 2
12 9 13 9 2 16 13 15 15 1 0 13 2
9 2 15 13 2 16 9 13 13 2
11 0 1 9 9 13 2 16 9 13 0 2
6 1 9 13 14 9 2
8 1 0 1 9 14 13 4 2
10 2 14 13 2 3 13 15 0 9 2
8 1 9 9 13 0 9 9 2
11 3 13 15 15 13 2 9 13 0 9 2
14 9 9 0 9 7 9 0 1 9 9 14 13 0 2
11 9 14 1 0 9 13 13 9 9 0 2
8 13 14 1 13 9 1 9 2
6 9 13 0 9 9 2
11 9 14 13 14 9 9 1 0 9 9 2
12 1 9 9 0 1 9 13 9 9 1 9 2
4 3 13 9 2
6 3 13 1 9 0 2
9 2 7 14 14 13 0 9 9 2
11 14 9 14 9 9 1 13 1 9 9 2
14 2 14 3 13 0 9 2 7 9 13 15 1 0 2
10 3 2 0 9 9 1 9 13 0 2
5 13 14 0 9 2
10 0 0 9 13 13 1 12 9 9 2
14 9 14 3 13 1 9 1 0 9 7 13 9 9 2
5 14 13 1 9 2
21 3 7 9 14 13 2 16 1 0 9 2 1 0 9 2 3 15 4 13 9 2
13 2 1 9 13 0 9 2 1 0 13 0 9 2
7 13 1 0 9 2 13 2
4 13 9 13 2
14 0 13 1 9 9 7 3 13 9 9 1 9 0 2
12 0 9 9 1 9 13 9 1 0 9 0 2
16 1 9 9 9 13 9 1 9 9 2 7 9 9 3 13 2
14 9 0 2 0 13 9 1 9 0 2 0 1 9 2
22 9 9 1 9 13 13 13 1 9 9 0 9 7 13 13 1 9 9 9 9 0 2
12 16 3 13 9 9 2 13 3 13 9 0 2
12 9 9 0 13 9 15 9 0 7 9 0 2
11 12 0 9 1 13 9 0 13 1 9 2
7 9 13 9 1 0 9 2
8 9 13 1 9 0 0 9 2
6 1 9 9 13 15 2
21 1 9 9 0 9 13 9 1 9 9 2 0 14 13 9 9 0 7 0 9 2
16 0 13 9 13 15 3 1 9 0 13 1 9 9 9 0 2
14 1 9 0 9 13 1 9 9 13 9 0 12 9 2
5 1 9 13 9 2
12 9 13 0 9 2 0 3 13 1 9 9 2
18 1 3 0 9 0 2 13 1 9 0 2 13 14 9 0 7 0 2
14 2 0 9 0 9 1 9 13 1 0 9 3 12 2
9 13 15 2 16 13 15 0 9 2
20 0 9 13 1 9 3 1 13 9 2 7 13 15 13 0 9 1 0 9 2
11 0 9 9 4 13 13 9 1 0 9 2
7 9 13 15 9 1 9 2
7 13 9 13 9 1 9 2
8 9 4 13 1 9 9 0 2
8 13 15 9 0 9 0 8 2
17 0 9 9 13 9 13 9 9 1 13 9 1 13 9 9 0 2
7 13 1 9 2 1 9 2
6 13 12 9 9 1 2
7 1 9 0 9 3 13 2
6 9 9 13 9 0 2
17 1 0 9 1 12 0 9 13 13 13 15 1 9 2 0 9 2
6 9 13 9 1 9 2
4 4 4 13 2
4 3 13 9 2
5 14 13 15 3 2
8 7 13 2 7 9 14 13 2
4 14 13 9 2
3 13 4 2
8 13 3 0 2 15 7 15 2
6 7 9 3 15 13 2
6 13 0 9 1 9 2
21 9 0 9 9 9 13 2 1 0 9 2 14 0 9 1 0 9 0 9 0 2
14 9 4 13 1 9 9 2 0 1 9 9 9 9 2
4 14 9 13 2
4 14 13 9 2
7 13 1 9 1 9 9 2
5 13 4 1 9 2
7 7 3 15 13 2 2 2
4 3 14 13 2
13 16 13 2 1 0 9 13 15 0 9 2 2 2
12 15 14 14 13 2 3 3 15 1 15 13 2
4 3 13 13 2
5 15 9 14 13 2
8 14 1 9 0 13 4 9 2
10 1 0 9 13 4 3 0 9 9 2
15 13 4 15 1 9 1 9 1 0 9 1 9 1 9 2
6 9 13 1 0 9 2
11 1 9 1 9 9 13 15 12 9 0 2
7 9 0 13 1 9 0 2
20 9 9 13 9 9 2 1 0 13 7 9 2 7 14 9 9 9 9 9 2
9 3 3 13 15 1 9 9 9 2
5 9 3 14 13 2
14 9 1 9 0 1 0 9 13 9 0 7 9 13 2
13 1 9 1 9 7 9 2 0 9 13 13 9 2
15 13 0 1 9 2 1 0 9 13 13 12 1 0 9 2
17 16 0 9 13 3 0 2 13 0 9 1 9 2 9 7 9 2
12 13 0 2 7 0 0 9 0 4 3 13 2
18 9 3 13 0 1 0 9 2 16 1 0 9 13 13 9 1 9 2
5 13 14 13 0 2
15 13 0 2 0 2 0 7 0 2 0 9 2 3 0 2
15 0 9 2 9 2 9 2 0 9 7 9 9 13 9 2
10 4 13 3 9 1 0 9 7 9 2
17 14 13 15 9 2 13 1 0 7 0 9 9 2 0 15 13 2
23 13 0 9 2 9 0 2 13 0 2 13 9 13 7 14 13 13 15 1 9 0 13 2
20 13 14 0 9 1 0 13 0 9 7 9 2 16 15 3 13 1 9 0 2
16 9 13 2 16 9 2 0 13 0 9 2 13 15 1 9 2
17 9 13 15 3 2 9 3 13 9 2 9 0 13 1 9 13 2
4 9 3 13 2
10 9 9 13 1 9 7 13 1 9 2
9 9 13 9 7 13 1 9 9 2
10 9 0 9 13 3 1 0 9 9 2
9 1 9 9 1 9 13 0 9 2
5 0 9 13 15 2
4 15 3 13 2
14 13 9 2 7 14 13 15 0 13 1 9 2 2 2
13 9 9 13 15 1 9 9 2 9 13 1 9 2
11 0 9 0 8 2 13 15 1 0 9 2
13 3 9 13 1 8 2 9 9 13 1 9 9 2
11 0 9 0 9 9 13 15 3 3 0 2
8 1 0 13 1 9 0 9 2
5 3 13 0 9 2
13 13 4 14 2 16 1 0 9 13 15 9 0 2
3 3 13 2
10 1 0 9 13 3 0 1 9 9 2
11 13 15 1 9 7 13 0 9 0 9 2
13 13 2 16 13 2 13 1 9 1 13 1 9 2
13 13 9 0 2 7 14 0 1 0 9 9 0 2
4 13 12 9 2
15 9 1 9 13 15 15 13 2 14 13 2 14 9 13 2
18 1 9 9 1 9 9 9 9 13 9 2 1 0 9 13 13 9 2
9 9 13 1 9 1 0 9 0 2
2 13 2
12 13 9 2 9 0 2 9 2 9 7 9 2
11 9 13 7 13 1 15 13 1 9 9 2
8 13 13 9 1 9 7 9 2
5 13 9 1 9 2
9 9 13 2 9 13 7 3 13 2
7 9 13 2 7 3 13 2
11 9 13 1 9 2 13 7 13 1 9 2
13 14 13 15 7 13 9 2 16 9 15 14 13 2
5 13 3 0 9 2
8 9 13 9 2 0 9 0 2
6 1 9 14 13 9 2
5 13 15 2 9 2
14 0 9 14 15 1 9 13 7 14 1 9 14 13 2
6 14 14 9 9 13 2
8 3 9 13 9 9 7 9 2
9 13 4 15 0 2 16 13 0 2
5 13 1 0 9 2
11 14 13 0 2 13 15 3 7 13 3 2
7 7 13 15 2 16 13 2
11 3 15 9 13 2 16 13 9 1 9 2
21 4 13 9 2 9 2 9 2 9 2 9 7 9 9 2 7 14 13 13 0 2
4 0 15 13 2
7 14 13 13 1 9 9 2
8 1 9 13 0 9 9 9 2
13 3 7 3 1 13 9 13 4 3 1 9 9 2
11 9 3 3 13 2 4 13 1 13 9 2
4 2 3 13 2
3 2 13 2
13 4 13 0 9 9 9 2 0 13 9 0 0 2
9 9 1 0 9 13 0 9 0 2
13 13 15 13 13 1 9 2 13 0 9 1 9 2
7 13 9 7 9 13 3 2
14 9 13 14 9 0 2 16 3 13 15 9 2 9 2
8 9 9 13 3 0 7 0 2
8 13 1 9 9 13 2 13 2
3 13 9 2
4 14 13 15 2
15 14 13 13 9 7 15 2 16 9 13 15 1 0 9 2
5 7 14 13 15 2
15 3 14 13 1 0 9 1 9 7 9 2 13 1 9 2
7 1 9 13 14 0 9 2
4 9 13 9 2
9 13 15 3 1 0 2 0 9 2
4 0 9 13 2
13 9 13 9 2 3 7 13 9 13 1 9 9 2
2 13 2
7 13 0 9 1 9 9 2
5 14 13 0 9 2
7 0 9 0 13 15 9 2
8 7 3 14 3 15 14 13 2
9 9 0 9 1 9 13 1 9 2
10 9 13 1 9 1 12 7 13 9 2
13 9 13 0 9 2 13 15 0 7 0 9 13 2
9 16 13 2 3 14 13 1 9 2
14 3 9 9 13 0 9 7 13 1 0 9 1 9 2
6 13 2 16 13 9 2
6 13 9 1 9 9 2
4 13 0 9 2
6 13 15 1 0 9 2
2 13 2
6 9 13 1 0 9 2
8 1 9 13 9 1 9 0 2
5 13 15 13 3 2
7 9 13 1 15 3 3 2
7 13 15 13 9 1 9 2
7 2 3 15 13 0 9 2
26 13 15 7 13 2 14 13 2 16 9 14 13 1 15 9 7 1 9 13 15 2 16 15 14 13 2
7 14 13 13 2 1 9 2
5 2 3 15 13 2
4 13 15 15 2
12 13 9 2 13 9 1 15 2 13 1 9 2
14 2 13 2 13 2 16 13 9 2 9 13 1 9 2
8 2 13 15 1 13 2 2 2
8 13 15 1 9 9 13 9 2
12 9 13 9 13 1 9 2 13 13 0 9 2
13 1 0 9 15 9 13 9 0 9 7 9 9 2
14 1 9 1 9 13 0 9 1 9 9 1 0 9 2
9 3 3 9 9 13 1 9 0 2
5 13 15 9 13 2
8 13 2 3 13 15 1 9 2
9 13 15 1 0 9 0 13 9 2
5 1 9 13 9 2
11 0 9 13 9 9 1 9 1 9 0 2
7 9 13 9 1 13 9 2
21 9 1 9 9 9 1 9 13 9 2 9 13 9 9 2 7 13 15 1 9 2
13 0 9 13 0 9 1 9 2 13 1 9 9 2
10 9 9 0 13 13 1 15 9 0 2
15 9 13 9 9 13 15 13 9 1 9 7 9 0 9 2
7 14 3 4 15 3 13 2
11 13 12 9 2 13 12 9 7 0 9 2
11 13 9 7 9 0 7 1 9 15 13 2
5 7 13 15 0 2
12 3 13 2 16 14 13 2 3 3 15 13 2
3 9 13 2
7 13 7 3 13 13 9 2
5 14 13 1 9 2
11 9 0 9 13 2 14 14 4 15 13 2
4 13 1 9 2
5 7 13 15 9 2
10 1 9 9 9 13 15 1 9 9 2
9 9 13 15 16 9 1 15 13 2
12 9 2 9 13 0 9 9 1 9 9 0 2
14 1 9 9 2 9 13 3 13 1 0 9 14 9 2
11 13 15 14 0 0 9 13 9 1 9 2
8 13 9 13 9 14 12 9 2
11 0 9 13 2 3 15 13 2 3 0 2
13 0 1 14 12 9 9 13 15 1 9 0 9 2
6 7 9 13 9 13 2
18 13 2 16 14 15 1 9 1 9 13 4 9 2 0 9 13 9 2
14 1 9 13 9 1 9 7 1 9 13 15 13 3 2
18 9 0 2 0 13 1 0 9 9 1 12 8 2 9 1 0 9 2
16 13 4 9 2 9 9 7 9 13 0 9 2 16 4 13 2
20 3 13 4 1 9 1 9 2 0 9 2 7 13 4 1 9 14 1 0 2
6 1 9 3 13 9 2
10 13 9 9 13 13 1 9 0 9 2
6 7 3 3 14 13 2
11 9 9 13 9 1 9 1 9 0 8 2
9 1 9 9 0 0 9 13 9 2
6 9 13 13 9 9 2
7 9 1 15 13 1 9 2
9 0 9 13 0 9 1 0 9 2
9 9 9 7 9 9 13 13 9 2
7 13 15 15 13 9 0 2
6 13 15 1 0 9 2
8 12 9 13 15 3 0 9 2
7 0 9 13 9 9 0 2
20 1 0 9 2 1 0 9 2 13 1 0 0 9 13 1 9 1 0 9 2
7 2 14 13 15 15 9 2
12 13 3 12 0 9 2 7 14 13 13 9 2
19 14 1 13 0 9 1 9 9 13 13 9 1 0 9 1 9 9 9 2
15 9 1 9 13 1 9 2 9 2 9 2 9 7 9 2
7 3 9 13 0 12 9 2
13 1 9 13 9 13 13 1 9 9 9 9 9 2
3 13 9 2
5 9 0 13 9 2
7 9 14 13 9 1 9 2
4 9 13 9 2
5 9 13 1 9 2
10 14 13 2 16 13 4 12 9 13 2
16 1 9 9 9 0 1 9 13 15 1 12 9 1 9 9 2
10 9 13 1 9 2 16 3 3 13 2
7 1 9 9 13 1 9 2
6 13 13 1 0 9 2
8 1 9 1 9 9 13 9 2
6 9 13 1 0 9 2
11 1 0 2 8 0 9 13 9 7 9 2
4 9 13 3 2
8 13 1 9 0 2 13 9 2
5 9 15 14 13 2
8 1 0 9 9 13 13 3 2
19 1 0 2 8 9 13 0 9 0 9 2 13 2 7 9 13 0 9 2
3 9 13 2
5 0 9 13 9 2
10 1 0 2 8 9 0 9 13 9 2
9 1 9 9 13 15 14 9 0 2
5 9 13 15 13 2
9 9 0 9 13 0 9 0 9 2
4 3 13 0 2
10 0 9 9 13 14 9 9 9 9 2
13 3 13 14 13 2 16 9 0 9 3 4 13 2
7 1 12 9 12 14 13 2
6 9 13 14 12 9 2
14 13 14 0 1 0 9 9 2 0 13 9 0 9 2
16 13 0 9 9 9 9 2 1 9 13 0 9 7 13 9 2
7 3 3 13 9 7 9 2
12 9 0 13 13 9 0 1 9 0 9 0 2
13 9 9 9 13 15 2 7 9 7 9 13 9 2
9 1 0 9 14 13 9 1 9 2
14 16 9 13 1 15 13 2 9 13 15 3 2 2 2
10 0 9 13 2 0 9 2 0 9 2
17 3 0 9 0 9 1 9 14 13 2 1 9 1 9 0 13 2
9 14 9 13 2 16 9 13 0 2
5 13 15 9 0 2
12 7 1 9 14 13 2 13 1 9 1 9 2
26 9 1 0 9 13 1 9 2 13 15 0 2 0 9 0 9 2 1 0 13 3 1 9 1 9 2
6 14 9 13 3 9 2
14 1 9 13 14 4 13 15 15 9 14 1 9 9 2
17 9 13 14 2 16 9 1 13 1 9 13 15 14 1 0 8 2
4 15 13 9 2
13 16 14 15 9 13 1 0 9 2 16 3 13 2
18 3 9 13 1 9 12 8 2 9 9 7 14 13 0 0 9 0 2
5 9 13 14 9 2
9 9 13 7 9 1 9 7 9 2
7 7 1 9 13 1 9 2
9 7 15 3 9 13 0 7 0 2
8 14 12 0 9 13 15 9 2
15 1 9 9 8 2 9 3 13 9 9 9 0 1 9 2
10 0 9 1 9 9 13 9 9 9 2
13 9 14 13 14 13 2 16 9 13 1 15 9 2
9 9 0 13 1 0 12 8 8 2
13 1 0 9 9 13 15 1 0 9 13 9 9 2
22 1 0 9 0 9 9 2 13 9 0 2 13 1 0 9 9 13 9 13 9 9 2
29 1 9 9 14 13 1 9 9 9 9 13 9 1 9 2 7 1 9 9 9 14 13 15 9 1 9 9 9 2
14 14 13 14 2 16 9 13 1 9 1 9 13 0 2
12 9 13 9 1 0 9 0 1 9 9 9 2
15 2 3 13 9 2 0 13 15 13 2 16 15 14 13 2
16 3 7 9 2 7 14 9 13 0 9 1 9 9 1 9 2
13 13 14 13 15 1 9 2 13 9 2 13 9 2
25 16 13 9 1 9 13 4 0 9 9 7 13 4 9 1 9 0 2 13 15 12 9 1 9 2
10 14 1 9 9 13 15 9 7 9 2
15 3 9 0 9 9 9 0 13 9 1 9 0 2 13 2
25 1 9 13 15 3 3 2 16 0 9 1 3 13 0 9 13 1 13 1 9 9 13 9 0 2
19 0 9 1 9 1 9 9 13 0 7 0 9 12 9 13 1 9 9 2
19 13 15 15 1 0 9 1 9 1 9 1 0 9 7 13 15 9 0 2
11 13 15 14 1 9 13 9 0 1 9 2
17 9 9 13 1 0 9 9 1 0 9 9 13 9 0 7 0 2
14 9 13 2 16 3 13 4 13 9 9 9 7 9 2
20 1 9 0 2 9 9 1 9 2 13 9 9 2 16 3 0 9 13 15 2
7 3 3 13 1 9 0 2
10 1 0 8 2 13 15 0 13 9 2
11 14 3 13 14 14 13 1 0 9 9 2
11 7 13 14 0 2 0 7 0 2 9 2
3 13 9 2
11 9 13 9 9 13 1 15 0 0 9 2
8 1 9 13 15 7 15 9 2
6 9 13 9 0 9 2
14 9 9 1 0 9 13 14 1 9 9 9 1 9 2
4 9 15 13 2
20 16 15 14 13 1 9 13 2 9 13 1 9 9 2 7 13 13 1 9 2
9 16 14 13 9 15 0 9 9 2
6 1 9 9 14 13 2
21 0 7 0 9 2 3 14 0 2 3 3 13 15 1 0 9 1 9 9 9 2
10 9 13 2 16 14 13 9 3 13 2
11 9 13 2 16 9 13 3 0 3 9 2
10 9 13 2 16 14 13 15 1 9 2
17 9 0 9 13 3 2 16 13 0 9 9 2 13 1 0 9 2
13 0 1 15 1 0 9 14 13 9 9 9 9 2
8 1 9 1 9 13 15 9 2
4 13 1 9 2
7 1 0 9 13 0 9 2
13 1 9 0 9 13 13 1 0 9 1 0 9 2
15 13 15 13 2 13 1 9 7 9 2 16 13 13 9 2
7 1 9 13 15 1 9 2
5 14 9 4 0 2
3 13 9 2
7 1 0 9 9 13 9 2
17 13 3 9 2 13 1 15 9 7 9 2 9 15 13 15 13 2
17 9 2 13 15 1 9 0 1 0 8 2 2 13 1 0 9 2
7 7 3 14 13 13 9 2
10 3 9 13 1 9 13 14 12 9 2
6 14 13 15 13 9 2
14 1 9 9 13 12 9 9 2 7 13 14 12 9 2
11 1 9 1 13 9 9 13 13 9 9 2
13 13 1 9 2 0 13 9 1 9 1 13 9 2
11 1 9 13 15 0 9 2 1 9 9 2
5 13 15 1 9 2
6 13 1 9 0 9 2
6 13 9 9 4 13 2
21 9 13 15 1 9 2 7 9 7 9 14 13 9 2 16 13 15 0 0 9 2
8 1 0 9 3 13 1 15 2
15 14 13 15 9 1 13 2 16 9 0 13 0 1 0 2
17 1 9 13 15 9 9 2 9 9 2 1 9 3 13 1 9 2
15 13 9 7 0 0 9 2 13 15 1 9 0 0 9 2
8 9 13 3 1 0 9 9 2
10 9 13 2 9 13 15 9 7 13 2
5 3 13 12 9 2
9 14 13 15 2 16 13 1 9 2
13 13 1 9 7 13 2 16 13 1 9 0 9 2
13 13 1 9 2 16 13 15 1 9 13 3 3 2
5 9 15 9 13 2
12 13 1 9 2 16 9 13 0 9 2 9 2
7 1 15 9 9 15 13 2
16 13 0 9 1 0 9 7 0 2 0 9 2 0 9 0 2
8 2 13 15 2 16 13 9 2
4 15 15 13 2
16 1 12 9 3 9 4 3 13 1 9 2 16 9 9 13 2
4 13 9 9 2
9 13 3 2 1 9 9 15 13 2
24 13 14 13 1 9 9 2 3 0 2 0 9 7 13 15 2 16 1 15 9 9 9 13 2
14 1 0 9 14 13 4 0 9 7 9 13 1 9 2
12 13 1 15 0 1 9 9 1 3 0 9 2
13 13 14 9 9 2 9 0 2 9 0 7 9 2
8 7 13 3 3 1 9 0 2
3 13 4 2
3 2 13 2
7 2 15 13 13 1 9 2
6 13 9 1 0 9 2
6 2 14 4 13 3 2
2 13 2
6 9 13 15 1 15 2
6 13 15 14 12 9 2
7 2 13 4 15 1 15 2
6 13 1 9 0 9 2
7 13 1 9 9 0 9 2
13 13 3 1 0 9 2 16 13 2 3 15 13 2
5 2 3 15 13 2
9 14 3 13 4 3 13 1 9 2
11 3 13 4 15 9 7 13 4 1 9 2
10 13 4 14 9 1 0 9 1 9 2
8 9 13 3 1 9 13 9 2
9 1 3 13 0 0 2 0 9 2
7 13 9 1 9 9 0 2
14 9 9 13 7 2 16 9 0 13 15 13 1 9 2
6 2 13 13 9 9 2
7 2 14 13 4 9 0 2
6 2 13 2 15 13 2
8 2 13 2 3 2 15 13 2
6 9 3 13 14 3 2
4 3 13 9 2
4 14 13 9 2
14 9 9 14 0 15 13 1 9 9 2 7 14 9 2
10 0 9 9 13 15 9 0 9 0 2
5 15 13 12 9 2
12 9 0 3 13 9 13 13 1 9 1 9 2
23 13 9 9 0 9 1 8 2 12 8 9 2 1 16 1 9 0 9 13 15 3 0 2
7 2 3 9 13 12 9 2
23 1 16 3 14 13 2 3 4 13 0 9 9 2 9 0 9 13 0 9 1 0 9 2
18 0 13 9 15 9 2 3 3 0 2 13 1 0 9 0 9 0 2
8 16 1 9 9 0 4 13 2
12 9 2 9 9 13 1 0 9 0 9 0 2
19 9 2 9 2 0 13 0 9 1 9 2 13 0 9 1 9 7 9 2
15 9 13 2 16 3 13 15 1 9 9 1 9 9 9 2
10 1 0 9 14 4 14 1 9 13 2
6 15 9 13 0 9 2
8 9 13 15 1 9 9 3 2
9 0 9 9 9 13 1 9 9 2
9 1 13 9 2 9 13 0 9 2
6 9 13 14 0 9 2
20 7 13 9 14 0 1 9 2 13 1 0 9 9 1 0 2 3 13 9 2
7 1 9 13 15 15 3 2
7 14 13 9 1 0 9 2
6 13 15 3 1 9 2
8 1 9 13 15 14 9 9 2
10 3 1 13 1 15 13 15 9 9 2
8 7 3 13 2 14 13 3 2
13 4 13 0 9 2 0 1 9 2 1 0 9 2
12 13 0 9 2 7 1 15 13 13 0 9 2
5 13 15 0 9 2
9 9 13 15 9 0 9 7 9 2
11 1 15 9 13 13 12 9 0 7 0 2
16 1 0 1 15 13 4 9 1 9 2 13 9 2 9 9 2
20 3 13 4 0 9 2 1 0 9 2 13 0 9 1 9 0 9 1 9 2
4 13 15 9 2
9 13 9 7 1 9 13 9 9 2
3 13 13 2
11 13 13 15 1 9 2 13 0 9 9 2
11 9 13 15 2 3 13 9 7 9 0 2
11 13 15 14 9 1 9 9 1 0 9 2
17 9 13 14 13 0 9 7 13 1 9 3 1 9 2 13 9 2
4 9 13 9 2
26 9 13 0 7 0 2 7 13 1 0 1 9 9 2 13 1 0 9 2 13 0 0 9 12 9 2
11 7 13 15 0 9 2 3 1 15 13 2
14 13 14 7 9 1 9 2 7 1 9 9 1 9 2
3 13 0 2
4 13 15 3 2
5 3 13 14 9 2
7 13 15 13 14 13 12 2
8 7 14 0 0 9 3 13 2
10 0 9 0 13 15 3 1 9 9 2
17 7 16 14 4 1 0 9 13 0 9 2 13 13 0 9 9 2
13 1 0 9 13 9 0 13 0 9 1 0 9 2
20 9 13 14 2 16 9 4 15 13 1 9 2 16 1 0 9 13 12 9 2
17 1 9 0 9 0 9 13 1 9 13 4 13 14 1 0 9 2
20 13 9 2 13 1 15 3 2 13 1 9 13 9 2 1 15 9 13 9 2
5 1 9 13 9 2
8 9 13 1 9 1 9 0 2
9 0 9 13 0 2 0 13 9 2
4 13 2 13 2
8 2 3 13 1 15 1 9 2
19 2 3 2 3 2 13 2 3 13 4 0 9 13 3 3 1 9 9 2
5 2 13 0 9 2
13 9 1 0 9 13 9 1 9 9 1 9 0 2
16 2 9 13 9 1 9 13 0 13 1 9 7 13 9 0 2
24 9 13 1 9 9 1 13 9 1 9 2 7 9 13 1 0 9 13 9 1 9 9 9 2
11 1 9 9 1 9 13 14 4 0 9 2
5 13 9 9 0 2
4 9 13 3 2
4 9 15 13 2
7 15 9 13 1 9 9 2
10 13 9 2 9 2 13 15 1 9 2
8 7 0 9 13 14 0 9 2
7 3 9 9 9 13 15 2
5 3 4 3 13 2
5 9 13 1 9 2
7 13 9 9 7 3 13 2
10 3 13 15 7 3 13 15 1 9 2
3 13 13 2
5 13 3 9 9 2
2 13 2
4 2 13 9 2
4 9 13 9 2
7 2 9 13 9 1 9 2
11 14 9 9 13 9 9 1 9 0 9 2
16 14 9 13 2 1 9 1 9 2 13 15 9 1 9 9 2
10 14 2 3 9 15 13 1 0 9 2
3 13 9 2
6 3 13 14 4 13 2
9 1 0 9 13 4 0 9 9 2
5 13 3 1 9 2
2 13 2
13 0 9 14 13 13 2 14 13 14 15 0 9 2
10 9 13 1 0 9 1 9 9 0 2
6 9 13 1 9 0 2
6 14 9 9 4 13 2
11 13 1 15 9 2 13 3 7 13 9 2
7 14 9 1 15 13 0 2
5 13 15 1 9 2
11 2 9 3 13 9 1 0 9 2 2 2
11 9 9 13 14 9 7 9 9 9 9 2
5 2 9 13 0 2
5 2 13 14 2 2
11 2 9 2 3 9 13 1 9 2 2 2
5 13 9 0 9 2
8 13 4 0 9 9 1 9 2
3 2 13 2
19 14 13 9 1 9 2 13 4 13 1 9 2 0 4 15 13 1 9 2
8 0 9 9 13 3 1 9 2
11 0 9 9 4 13 14 14 1 12 9 2
14 0 9 9 14 13 15 0 9 1 9 0 2 2 2
17 9 14 13 14 9 1 9 9 13 9 7 13 9 1 9 9 2
8 13 13 1 9 9 0 9 2
11 3 3 13 9 0 2 0 1 9 0 2
7 9 0 13 9 12 9 2
15 1 9 0 9 0 9 2 9 13 0 9 9 13 9 2
12 1 9 0 9 9 13 13 12 8 2 9 2
11 3 13 9 2 3 13 15 1 9 9 2
13 14 1 0 9 13 15 13 7 1 0 9 13 2
5 9 13 0 9 2
8 1 9 0 13 3 9 9 2
10 13 3 9 13 9 13 9 0 9 2
15 1 9 1 13 1 9 9 9 13 9 13 9 1 9 2
6 13 4 14 9 0 2
8 13 4 3 9 9 1 9 2
9 14 1 0 9 13 4 9 9 2
23 14 1 12 9 13 15 2 16 3 0 9 1 13 0 9 13 0 9 9 2 9 9 2
14 1 8 2 9 7 9 13 4 1 0 9 0 9 2
11 9 0 13 15 1 9 0 9 9 9 2
18 12 9 9 9 13 12 9 2 0 1 0 1 0 9 13 0 9 2
13 9 0 3 1 0 9 13 15 1 9 0 9 2
9 9 9 13 0 9 7 0 9 2
20 1 0 9 4 13 13 1 3 13 9 2 9 13 9 2 9 7 0 9 2
13 1 0 9 0 15 13 9 9 1 8 2 0 2
11 9 13 15 13 1 9 2 13 12 9 2
9 9 13 15 1 9 0 2 12 2
10 9 13 9 13 13 0 9 1 9 2
20 9 9 4 13 1 9 0 1 9 1 9 1 8 2 0 1 8 2 0 2
10 13 9 9 1 8 2 9 1 9 2
18 1 9 13 12 9 1 2 1 9 13 14 9 0 0 9 7 9 2
8 9 9 13 4 13 14 3 2
19 1 3 0 0 9 13 13 9 7 9 2 3 13 9 13 15 1 15 2
13 9 13 14 9 0 2 0 13 4 1 0 9 2
18 13 15 0 9 0 2 3 13 9 0 2 7 1 15 0 9 0 2
5 9 13 13 9 2
6 9 13 15 13 3 2
10 9 13 9 1 9 1 0 9 8 2
5 14 13 13 9 2
5 3 15 15 13 2
19 1 9 0 13 9 2 7 15 3 13 15 1 9 9 2 0 13 0 2
6 14 3 13 13 15 2
3 13 9 2
8 0 9 13 9 0 1 9 2
4 9 3 13 2
15 13 1 15 0 2 13 2 16 9 13 14 13 3 0 2
7 3 13 4 0 9 9 2
6 0 9 13 1 9 2
11 13 1 9 0 9 2 0 13 1 9 2
8 0 9 13 15 0 0 9 2
6 13 1 15 14 9 2
5 7 1 9 13 2
8 0 9 9 4 13 1 9 2
8 14 3 13 15 0 0 9 2
8 13 4 9 2 12 0 9 2
7 7 13 0 0 0 9 2
12 7 15 4 13 2 16 1 0 13 9 9 2
27 13 1 0 9 2 9 13 9 2 1 0 13 15 1 0 9 2 7 13 9 2 16 13 13 13 9 2
12 13 3 2 7 13 15 13 2 13 1 9 2
13 13 1 9 1 9 2 3 2 1 9 14 13 2
7 7 9 13 15 13 3 2
2 13 2
5 13 4 0 9 2
13 16 9 0 13 13 15 1 15 2 13 0 9 2
7 9 9 13 1 15 9 2
6 9 13 9 1 9 2
8 13 13 3 0 1 0 9 2
9 0 9 13 1 15 1 13 9 2
11 2 13 4 0 9 2 7 15 15 13 2
10 0 9 1 9 13 15 1 0 9 2
12 1 0 9 13 9 1 13 9 1 0 9 2
6 9 9 9 9 13 2
9 2 9 9 2 14 15 9 13 2
5 2 9 15 13 2
7 2 13 15 1 9 0 2
6 0 9 14 13 9 2
6 2 14 13 4 9 2
12 3 13 2 0 9 14 13 0 9 1 9 2
15 9 13 1 9 2 13 1 9 1 9 9 1 0 9 2
13 9 9 0 3 13 1 0 9 1 9 7 9 2
16 0 9 0 13 9 1 0 9 2 7 9 0 9 13 15 2
19 0 9 0 9 13 7 4 13 2 16 0 0 9 13 15 1 0 9 2
6 3 14 13 9 0 2
6 3 15 13 0 9 2
4 3 9 13 2
5 14 13 9 9 2
7 2 7 9 15 3 13 2
10 2 13 2 16 9 13 9 9 9 2
13 13 1 9 0 9 14 1 9 0 13 13 9 2
12 9 1 0 9 13 4 13 1 9 0 9 2
10 4 13 3 3 2 14 13 9 9 2
14 1 12 9 1 0 9 13 9 1 0 9 9 0 2
8 13 9 7 13 9 7 9 2
8 2 13 15 3 9 0 9 2
10 14 1 0 9 13 3 13 1 9 2
11 9 13 1 12 13 1 9 8 2 9 2
10 0 9 13 14 1 9 1 9 9 2
6 16 9 0 9 13 2
9 2 14 13 14 2 9 13 3 2
8 13 4 7 1 9 1 9 2
5 14 13 0 9 2
4 9 3 13 2
11 3 0 9 13 15 13 0 2 0 9 2
13 9 13 0 1 0 9 1 13 0 1 0 9 2
9 9 13 13 0 9 1 9 9 2
22 0 9 7 9 13 0 9 9 9 2 13 15 1 9 9 7 13 1 0 9 0 2
13 13 1 9 13 9 0 9 7 13 1 15 9 2
6 9 9 13 13 9 2
9 9 13 15 9 9 7 9 9 2
6 14 13 14 9 0 2
13 13 9 1 9 1 9 1 9 7 13 1 9 2
6 2 13 15 1 9 2
14 9 0 7 0 9 13 2 16 9 4 14 3 13 2
7 13 9 7 13 1 9 2
8 13 4 13 9 2 16 13 2
11 13 9 1 9 7 13 0 9 1 9 2
8 9 3 14 13 2 13 9 2
10 13 14 15 13 2 1 9 13 9 2
12 9 13 1 9 1 9 2 7 9 13 9 2
5 13 15 1 9 2
8 2 13 15 7 13 1 9 2
10 9 0 9 9 13 15 7 13 9 2
11 9 13 1 9 9 1 9 1 9 0 2
9 13 1 15 0 7 0 9 9 2
12 13 4 9 9 13 1 9 9 1 12 9 2
16 13 4 9 9 2 0 13 15 9 1 0 9 0 0 9 2
9 16 14 9 13 9 1 9 9 2
6 13 9 7 0 9 2
23 13 1 0 9 7 9 2 16 9 9 13 15 1 0 9 7 13 13 1 9 0 9 2
6 14 13 13 0 9 2
11 13 1 0 9 0 9 2 14 3 0 2
9 2 9 13 1 0 9 9 0 2
11 3 9 4 13 7 3 13 1 9 0 2
26 13 15 13 2 16 14 13 4 2 16 13 13 9 2 16 14 9 9 1 0 9 13 4 1 9 2
9 3 13 15 1 13 9 1 9 2
31 13 7 13 15 9 2 16 1 12 9 13 15 13 1 13 9 2 9 13 15 2 16 13 14 4 13 3 3 1 15 2
13 13 14 1 9 2 7 15 9 1 9 14 13 2
