491 11
54 11 3 13 14 9 15 2 11 7 11 16 13 4 13 1 9 2 13 1 11 7 11 16 13 14 10 10 9 10 0 9 16 13 1 10 9 13 1 9 13 11 13 2 11 7 11 13 1 10 10 9 1 9 2
13 1 10 9 10 2 12 13 9 10 9 12 12 2
16 9 15 14 11 13 1 9 14 9 10 9 1 2 12 12 2
18 7 11 7 11 13 1 9 15 7 13 14 10 9 2 12 12 2 2
16 3 13 13 16 9 10 9 13 7 7 3 1 10 9 11 2
7 15 13 3 13 14 15 2
37 13 1 15 9 11 16 13 14 10 9 1 9 0 2 1 11 11 1 9 9 16 13 14 9 11 3 0 2 16 3 13 1 11 3 16 13 2
18 11 13 15 1 2 12 2 9 12 2 7 2 12 2 9 12 2 2
28 9 15 14 11 1 9 10 9 1 11 2 7 9 15 14 11 1 9 10 9 2 13 14 11 1 10 9 2
35 11 13 1 9 9 2 12 1 9 9 2 16 13 9 1 10 9 1 9 11 1 1 12 9 3 2 12 12 1 10 9 10 2 12 2
23 7 10 9 14 11 2 1 9 9 0 2 12 1 9 9 2 13 14 11 1 9 0 2
28 1 10 9 1 15 13 11 9 2 3 1 10 9 11 3 3 2 12 2 3 13 1 10 9 1 3 13 2
38 9 15 10 0 14 11 7 11 13 1 9 12 0 14 11 9 9 1 9 15 1 10 9 2 12 9 1 10 9 2 7 11 16 13 1 9 12 2
8 3 16 10 9 13 1 9 2
28 10 3 2 16 10 9 10 15 16 2 13 2 7 13 1 9 0 2 13 1 9 9 9 1 9 10 9 2
20 3 16 13 1 15 2 3 1 10 9 10 0 2 13 9 11 12 1 11 2
18 9 15 14 11 11 13 1 10 9 1 10 9 2 1 9 14 9 2
9 1 9 15 13 14 11 9 9 2
7 4 3 13 14 10 9 2
14 1 15 16 13 1 15 9 2 7 16 3 15 13 2
18 12 1 11 13 1 10 9 1 11 7 13 9 0 10 9 9 9 2
24 10 9 12 12 1 10 9 13 9 2 3 1 10 0 16 15 9 0 12 1 15 1 9 2
14 11 4 13 15 3 2 3 1 9 10 9 1 12 2
15 7 10 9 10 0 14 10 9 10 2 12 13 1 11 2
13 12 12 1 10 9 11 9 9 2 1 12 9 2
5 11 13 9 0 2
10 1 11 9 15 13 3 1 10 9 2
15 11 11 13 9 10 9 1 12 9 7 9 9 0 3 2
16 1 9 11 16 13 3 12 9 15 3 9 10 9 10 0 2
9 9 10 9 13 1 9 10 11 2
30 10 9 10 0 13 14 10 9 10 9 11 12 12 7 13 1 15 9 9 0 16 13 14 15 1 10 9 10 0 2
20 9 10 11 13 12 9 1 10 9 10 0 7 13 3 14 11 7 11 11 2
12 12 9 9 0 13 1 9 11 7 1 11 2
23 10 9 9 0 13 14 10 9 1 9 16 13 1 11 7 13 14 11 9 9 12 12 2
14 1 10 9 11 13 3 3 0 1 11 11 12 12 2
4 3 1 9 2
14 11 11 16 13 1 9 1 9 15 13 3 9 9 2
16 10 9 13 1 9 0 12 9 7 13 1 9 1 10 9 2
8 15 13 13 3 1 12 9 2
20 9 13 1 10 9 3 13 14 10 9 11 1 10 9 10 0 1 15 13 2
15 1 11 13 3 16 13 2 7 13 2 9 1 9 0 2
21 10 9 16 13 1 9 10 9 13 2 16 0 1 3 11 11 13 9 10 9 2
21 3 1 15 3 13 2 16 10 9 16 13 1 9 9 10 9 0 1 10 9 2
6 3 13 13 9 0 2
16 10 9 13 1 12 9 2 1 10 9 10 0 7 1 9 2
23 1 10 9 10 12 13 10 9 1 9 12 10 9 10 0 14 10 9 2 11 7 11 2
11 3 13 11 9 7 3 4 13 9 0 2
23 10 9 13 13 1 9 9 15 14 10 9 11 11 11 1 9 15 10 0 14 10 9 2
13 13 13 14 10 9 1 11 11 1 9 10 9 2
19 3 13 10 9 2 16 13 1 9 10 9 1 10 9 16 13 2 13 2
21 10 9 11 11 3 4 13 13 2 10 9 13 1 9 1 16 13 1 9 9 2
45 2 15 13 1 10 9 3 13 13 9 2 2 15 9 1 10 9 16 13 3 10 9 10 0 11 11 2 1 9 1 10 9 10 0 1 10 9 10 0 14 10 9 1 9 2
47 10 9 1 10 9 10 0 7 1 10 9 13 1 9 10 9 1 10 9 1 9 11 14 10 9 10 0 1 11 2 12 1 11 2 16 13 10 11 14 11 1 10 9 10 3 0 2
47 10 9 13 1 12 10 9 1 9 10 9 2 12 12 1 9 10 9 7 2 12 12 1 11 7 1 10 9 10 0 1 9 11 16 13 2 1 15 13 11 12 12 14 11 1 11 2
14 11 13 7 13 2 16 1 10 9 10 0 9 0 2
20 2 10 9 10 0 13 1 10 0 2 7 1 10 9 10 0 13 9 0 2
11 10 9 10 0 13 1 15 1 9 12 2
25 10 9 10 0 13 1 10 9 14 15 7 13 9 2 3 1 10 9 10 0 7 1 10 9 2
17 10 9 1 11 13 1 15 14 10 9 2 7 3 15 10 9 2
15 7 13 9 0 1 11 13 1 15 9 13 1 10 9 2
10 15 13 3 2 7 13 9 1 13 2
8 10 9 13 1 15 9 2 2
15 9 9 9 10 9 11 11 13 3 13 1 9 3 0 2
20 15 13 2 16 3 4 13 9 3 0 1 10 9 10 0 1 1 12 9 2
21 11 11 13 16 10 9 14 15 3 13 1 9 14 9 9 7 3 13 1 9 2
22 9 10 9 11 11 13 13 9 1 10 9 7 13 16 3 11 13 12 12 1 11 2
20 9 10 9 11 11 13 16 11 13 9 0 2 7 13 1 15 9 14 9 2
13 2 13 1 15 12 12 9 1 12 12 1 11 2
29 4 13 1 10 9 14 15 1 9 14 9 1 11 2 11 7 3 1 16 13 9 4 13 1 9 1 0 2 2
17 9 9 10 9 11 11 13 16 10 9 14 15 3 13 1 11 2
15 11 11 11 13 13 9 1 10 9 1 10 9 10 0 2
15 10 9 10 0 13 3 1 9 9 16 13 1 9 11 2
17 3 1 10 9 13 9 9 1 10 9 11 1 10 9 10 0 2
24 10 9 13 2 16 1 10 9 10 0 3 13 9 1 9 7 2 7 9 10 9 1 11 2
14 9 1 12 9 13 3 1 9 10 9 14 9 11 2
22 1 9 15 13 10 9 11 9 9 14 10 9 10 0 10 9 11 10 9 12 12 2
19 1 9 12 10 9 13 9 12 12 7 1 9 10 9 10 0 12 12 2
42 0 13 13 3 14 11 11 2 9 10 9 11 10 9 2 13 1 9 10 9 0 1 10 9 13 3 13 9 15 13 14 10 9 2 3 13 10 9 1 10 9 2
43 1 9 2 9 11 9 9 7 9 8 8 3 13 9 9 1 9 10 9 10 0 2 1 15 3 13 1 10 9 15 9 2 1 3 10 9 1 11 1 10 9 11 2
7 3 15 13 1 12 9 2
17 7 3 16 13 3 1 10 9 1 9 7 9 9 13 9 11 2
16 10 9 13 3 14 11 2 7 9 11 13 10 0 1 9 2
10 11 11 7 11 11 13 9 10 9 2
22 11 13 12 9 2 9 0 2 7 11 13 12 9 7 2 12 9 0 1 10 9 2
23 9 10 9 10 0 13 1 10 10 9 7 3 13 0 1 13 14 9 15 14 11 9 2
10 9 9 9 13 3 9 1 9 15 2
33 7 11 11 7 11 11 2 7 1 9 3 11 11 2 13 10 10 9 0 3 3 9 10 9 11 11 2 11 11 7 11 11 2
19 1 10 9 10 0 13 10 9 0 2 16 9 9 13 13 13 1 11 2
25 10 9 10 0 14 11 1 9 15 13 9 12 2 1 9 10 9 1 10 9 2 12 12 2 2
27 1 10 9 10 12 13 4 16 11 2 16 13 9 0 1 9 10 9 2 3 13 13 3 14 9 15 2
19 7 9 0 14 11 7 11 11 2 9 10 9 2 13 1 10 9 13 2
11 10 9 10 0 13 12 9 1 10 9 2
15 11 11 13 9 2 13 3 1 10 9 7 13 1 9 2
10 15 13 9 12 7 13 9 12 12 2
25 11 13 14 10 9 9 0 7 11 11 2 12 9 1 9 10 9 2 13 13 1 9 12 9 2
10 15 13 3 1 10 9 7 13 9 2
6 10 9 13 9 15 2
17 11 13 12 9 1 9 10 9 7 13 3 12 12 12 1 11 2
5 3 3 12 9 2
21 9 11 13 7 11 11 13 14 10 9 1 1 9 11 7 13 1 2 12 12 2
2 9 2
10 1 12 10 9 10 0 13 3 9 2
32 11 13 1 9 10 9 1 12 9 2 7 3 13 15 11 16 13 12 9 2 12 12 2 16 13 14 10 9 1 9 0 2
37 9 11 2 16 13 3 1 10 10 9 10 0 2 1 15 9 11 2 11 11 2 11 7 11 11 13 14 10 9 10 12 1 9 9 2 3 2
17 9 11 13 14 10 9 10 0 14 9 15 7 14 9 9 15 2
29 12 9 1 10 9 2 9 12 2 13 11 1 9 12 9 1 9 14 11 1 9 1 10 9 2 12 12 2 2
18 11 3 13 13 2 7 3 3 7 13 1 10 9 1 2 12 12 2
10 13 3 10 9 11 11 7 11 11 2
38 9 9 10 9 14 10 11 2 9 11 11 2 13 13 3 9 1 10 9 1 9 10 9 10 0 16 13 1 9 10 9 1 9 9 0 7 0 2
41 9 11 13 14 9 10 9 16 13 1 10 9 9 11 1 10 9 9 11 11 2 7 14 9 9 11 9 11 2 1 9 10 9 1 11 1 9 10 9 11 2
29 9 11 13 3 14 9 9 10 9 3 13 1 9 0 9 1 9 0 1 9 0 2 1 9 10 9 10 0 2
53 9 9 10 9 13 1 10 9 3 14 9 9 10 9 1 9 11 11 2 9 9 10 9 11 11 2 9 9 10 9 2 9 9 9 10 9 11 11 2 9 9 10 9 1 9 9 11 11 7 9 10 9 2
42 1 9 11 3 13 1 11 10 9 1 10 9 10 0 1 10 9 9 11 11 2 1 16 9 9 11 11 13 9 1 9 10 9 10 0 1 11 0 13 14 15 2
15 9 10 9 13 1 10 9 7 13 9 9 1 9 15 2
42 9 15 14 9 9 11 11 13 1 9 9 9 9 11 2 11 11 2 16 13 1 9 2 9 1 9 9 9 11 10 9 11 11 2 16 13 1 10 9 16 13 2
10 1 9 15 13 11 1 9 9 11 2
15 10 9 10 0 14 15 13 9 11 13 1 11 1 11 2
29 10 9 14 9 11 9 11 2 13 1 9 9 16 13 1 9 9 7 13 13 1 9 14 9 10 9 1 9 2
47 9 11 13 1 2 9 10 9 2 2 2 10 9 13 13 7 13 3 2 9 1 9 1 9 2 7 3 13 1 9 16 13 13 1 10 9 16 13 1 9 1 9 1 9 10 9 2
8 10 9 13 4 13 14 15 2
21 4 13 9 9 1 9 9 7 9 16 9 15 13 3 1 10 9 10 15 2 2
22 9 10 11 13 3 9 0 2 14 13 14 10 9 9 10 9 10 9 11 12 12 2
16 1 10 9 10 0 13 11 1 9 0 7 13 1 10 9 2
9 9 15 11 7 11 13 9 0 2
15 9 10 11 2 1 9 0 2 13 14 10 9 1 9 2
9 7 3 2 3 13 1 10 9 2
11 1 10 9 10 2 12 13 9 12 12 2
46 11 10 0 16 13 13 2 16 13 13 14 10 9 1 9 15 10 0 1 3 13 7 13 12 9 1 10 9 10 2 12 2 1 15 13 1 11 7 13 1 10 9 13 1 9 2
21 1 13 16 9 10 11 13 13 2 13 11 7 11 13 14 15 1 9 10 9 2
8 12 12 1 11 1 10 9 2
9 1 9 10 9 13 1 0 3 2
22 11 11 7 11 13 1 10 9 7 1 10 9 10 2 12 13 9 10 11 12 12 2
9 11 13 14 11 1 9 12 12 2
10 3 13 10 9 10 0 14 10 0 2
6 11 13 1 9 13 2
26 9 15 13 13 9 16 13 1 9 15 7 13 1 15 13 9 0 1 10 9 10 13 14 10 0 2
15 11 7 11 2 16 1 10 9 10 0 13 2 3 13 2
20 3 9 15 3 13 1 9 10 11 16 13 9 15 12 12 2 9 12 2 2
8 10 9 13 1 9 7 13 2
9 10 9 1 10 9 13 13 9 2
7 10 9 13 1 9 15 2
7 10 9 13 1 9 0 2
23 1 1 12 9 13 1 11 10 9 11 11 11 2 10 9 1 11 2 7 13 1 11 2
27 15 13 3 9 9 1 9 7 13 14 15 1 9 2 9 11 7 10 9 1 11 2 1 9 1 9 2
29 10 9 13 13 1 15 9 0 2 16 13 9 0 2 9 2 11 2 9 1 10 9 7 9 1 9 9 15 2
38 1 11 12 13 10 9 1 9 10 9 2 11 11 11 11 2 9 11 2 1 9 9 2 16 1 9 15 13 10 9 1 9 15 9 14 12 9 2
17 12 1 10 9 13 10 9 2 7 12 10 13 13 1 10 9 2
15 1 15 13 10 9 13 9 1 10 9 1 9 10 9 2
39 1 10 9 1 9 10 9 13 10 9 13 14 9 10 9 10 0 1 9 9 15 2 1 9 10 9 7 9 15 1 9 15 2 7 16 3 13 9 2
25 1 9 10 9 13 10 9 13 1 10 9 14 10 9 10 0 1 12 9 1 9 9 10 9 2
16 13 2 16 10 9 13 1 9 10 9 3 1 9 10 9 2
13 10 9 3 13 1 10 9 16 13 2 11 12 2
10 3 1 9 12 13 9 1 10 9 2
28 10 9 13 1 10 9 2 16 13 14 10 9 1 9 15 7 13 13 1 15 14 10 9 2 16 16 13 2
38 7 9 15 2 16 13 9 1 10 9 1 9 10 9 10 13 2 13 1 9 9 12 9 9 1 10 9 2 7 1 15 13 9 1 9 10 9 2
21 12 12 9 13 3 2 7 9 15 13 10 9 9 12 2 16 13 1 9 9 2
18 13 2 16 10 10 9 13 1 10 9 1 9 1 9 9 10 9 2
11 1 15 13 2 16 9 10 9 13 3 2
29 1 10 9 16 13 10 9 4 13 14 9 10 9 2 1 9 1 12 12 9 2 13 15 1 9 12 9 15 2
34 16 16 10 9 13 13 14 9 10 9 2 13 1 15 10 9 9 1 9 2 9 13 1 9 2 10 9 10 0 1 9 2 9 2
14 10 9 13 9 9 13 1 10 9 2 1 12 9 2
32 3 2 1 10 9 1 9 10 9 13 2 16 9 9 10 9 13 3 1 9 10 9 1 10 9 2 7 7 10 9 0 2
28 3 2 10 9 13 1 9 10 9 7 1 15 13 9 0 2 16 10 9 4 13 14 15 1 9 10 9 2
30 3 2 10 9 13 13 9 0 1 9 15 2 7 7 15 13 9 13 9 9 1 16 12 10 9 13 1 9 12 2
67 9 9 2 10 9 10 0 11 11 2 11 13 2 16 10 9 13 9 13 3 1 9 10 9 2 7 3 15 3 1 1 12 12 9 2 16 13 1 9 9 16 13 10 9 7 1 9 10 9 1 9 9 2 16 13 1 15 10 9 7 10 9 1 9 10 9 2
63 7 1 10 9 16 13 10 9 13 1 10 9 16 13 1 15 13 10 9 2 16 9 10 9 3 13 1 10 0 7 16 10 9 13 1 9 15 10 0 1 9 10 9 2 1 9 10 10 9 2 1 1 9 9 2 1 9 16 13 1 9 2 2
19 7 7 13 9 15 14 10 9 1 9 2 3 15 4 13 9 1 15 2
37 10 9 13 2 16 1 10 9 10 13 2 13 1 9 1 9 2 9 13 2 16 9 15 10 0 9 16 13 1 10 9 1 9 9 10 9 2
25 10 9 13 2 1 9 11 11 2 1 9 10 9 1 9 2 10 9 10 0 2 9 12 2 2
39 10 9 11 2 16 13 14 9 2 10 9 2 13 2 16 3 10 9 13 14 10 9 1 9 10 9 4 1 10 9 13 14 9 10 9 1 10 9 2
20 7 7 3 2 4 13 16 10 9 4 13 14 9 10 9 14 13 10 9 2
70 3 13 10 9 2 16 7 16 10 9 13 1 15 9 15 1 9 10 9 2 16 13 3 14 10 9 10 0 2 4 13 1 15 9 7 9 16 15 13 1 9 15 1 9 10 9 1 9 10 9 2 16 16 10 9 13 13 1 10 9 1 9 10 9 1 9 9 10 9 2
34 9 10 9 15 13 14 9 15 1 10 9 1 9 15 2 1 10 9 16 16 13 1 15 16 10 9 10 9 1 10 9 13 3 2
85 10 9 11 13 1 9 15 14 10 9 11 2 2 9 10 9 10 0 2 2 16 1 9 10 9 1 10 9 1 9 9 13 2 3 1 15 2 1 10 9 2 13 16 9 0 1 9 15 2 7 7 3 1 9 2 7 9 2 10 9 4 13 9 13 2 16 7 3 13 3 2 13 3 3 1 9 9 2 7 10 9 13 13 2 2
26 7 3 2 1 9 10 9 11 2 13 1 9 10 9 9 9 16 4 3 13 2 16 10 9 0 2
41 15 13 3 1 10 9 2 16 2 9 9 13 9 9 16 9 0 2 7 1 9 15 13 1 10 9 10 9 13 10 1 16 10 9 10 0 13 1 15 2 2
29 7 16 16 13 16 10 9 4 13 2 3 4 13 1 15 9 9 16 1 9 1 3 2 9 9 13 9 9 2
43 1 9 9 2 10 9 13 10 9 11 2 16 9 9 2 10 9 10 0 13 1 12 10 9 13 9 1 9 2 16 9 15 3 13 0 1 12 9 1 10 9 9 2
30 7 7 9 2 9 10 9 13 1 9 2 10 9 2 9 0 16 16 13 9 15 14 15 7 16 16 13 9 15 2
18 3 13 2 16 9 10 9 13 1 12 2 12 7 12 2 2 9 2
34 10 9 3 13 9 2 7 9 15 13 1 12 2 12 7 12 2 2 9 2 7 7 9 10 9 1 9 10 9 13 1 12 9 2
56 15 7 3 2 7 1 9 9 3 13 9 2 9 10 9 7 3 13 9 15 2 16 1 10 16 4 1 10 9 1 9 10 9 13 9 2 9 10 9 3 13 2 7 3 13 1 10 9 9 3 1 9 9 9 2 2
7 1 15 13 12 10 9 2
22 10 9 3 13 1 9 9 10 9 2 7 7 10 9 13 12 9 1 9 10 9 2
32 11 2 1 9 10 9 10 12 14 10 9 2 13 1 15 1 10 9 15 10 0 11 11 1 12 9 9 2 9 7 9 2
10 1 9 0 1 9 15 13 9 15 2
32 1 9 15 13 9 1 9 0 0 16 1 15 10 9 10 0 7 10 0 13 13 1 9 16 13 9 0 7 9 0 9 2
34 9 9 10 2 9 2 2 9 2 1 9 7 1 11 9 14 11 2 13 9 15 10 0 14 11 2 10 9 10 0 16 13 3 2
13 2 2 16 13 14 13 1 15 9 1 9 0 2
24 11 11 13 2 9 2 13 16 9 15 3 0 2 7 0 1 9 0 1 9 7 1 9 2
13 10 9 10 0 13 1 9 3 0 2 7 0 2
11 11 13 9 16 4 13 9 1 9 15 2
50 1 2 9 12 9 16 3 1 9 2 2 9 2 15 13 1 9 0 1 10 13 2 1 10 13 7 1 10 0 1 9 10 9 14 9 7 9 9 0 2 1 9 1 9 9 0 1 2 0 2
30 15 13 3 7 3 1 10 9 10 0 2 7 9 15 3 2 9 2 3 13 1 9 10 9 10 0 7 10 0 2
25 9 12 10 9 1 9 7 1 9 9 13 1 9 1 9 9 15 2 11 2 1 0 7 0 2
21 7 3 2 15 1 9 16 13 1 15 9 2 7 16 13 13 3 1 16 13 2
45 2 10 9 10 9 13 2 2 12 1 9 11 2 1 9 7 9 14 11 11 13 1 15 10 9 10 0 10 13 7 9 10 9 10 0 2 0 2 10 0 3 14 10 9 2
19 3 3 13 9 15 1 10 9 2 10 9 11 7 10 9 11 2 11 2
14 9 13 16 13 12 9 0 2 11 2 11 7 11 2
15 7 1 9 10 9 1 11 1 12 2 0 9 0 12 2
15 15 10 9 10 0 14 10 9 10 0 14 9 2 11 2
20 9 15 13 9 1 13 9 2 11 11 14 10 9 10 0 10 0 10 0 2
28 1 10 9 15 15 9 0 14 9 2 10 9 2 16 3 0 13 13 1 9 2 16 13 1 11 7 11 2
16 10 9 13 13 1 9 1 12 9 2 7 3 15 13 13 2
9 1 12 1 12 13 15 9 0 2
12 9 2 13 9 0 2 3 13 13 1 15 2
38 15 13 9 10 9 10 0 10 0 3 14 10 11 2 16 13 1 11 2 9 15 14 9 2 11 2 7 10 9 16 1 15 13 7 13 11 11 2
10 1 12 13 9 15 14 11 1 11 2
38 1 9 12 13 11 11 7 11 11 1 9 2 16 1 15 13 9 15 1 9 9 15 14 9 9 9 9 11 16 13 9 0 1 9 2 10 9 2
21 11 13 1 9 15 9 13 14 9 10 9 10 0 16 13 1 9 2 10 9 2
14 1 9 11 15 13 9 1 9 0 13 16 13 9 2
25 1 12 13 0 1 10 11 9 0 2 0 16 13 13 1 10 9 10 9 10 0 14 10 11 2
26 1 9 11 10 0 1 11 13 11 1 10 10 9 16 13 1 9 2 10 9 1 9 12 14 11 2
22 15 13 14 10 9 7 13 14 10 9 1 10 9 1 9 2 11 2 3 1 11 2
31 1 12 2 16 10 9 13 14 10 9 10 9 2 0 3 14 11 10 9 10 0 14 9 2 11 13 10 9 10 0 2
11 13 13 16 13 9 15 3 1 9 0 2
11 13 13 3 1 9 2 11 7 1 11 2
19 1 10 9 1 11 7 11 1 12 2 13 11 9 1 9 9 10 9 2
20 10 9 13 1 9 15 1 1 9 9 1 9 15 3 14 9 0 2 0 2
13 10 9 16 13 1 9 15 13 3 13 14 15 2
32 1 9 10 12 13 3 10 9 14 10 9 14 11 2 7 9 15 13 9 9 1 9 9 0 1 15 1 9 2 10 9 2
43 11 11 2 9 9 0 1 11 2 13 1 12 16 9 15 13 9 16 1 10 9 1 11 11 2 16 13 1 12 9 16 13 14 9 15 14 10 9 1 9 10 11 2
14 7 10 9 13 3 1 9 9 1 10 9 10 0 2
20 9 10 11 2 16 3 13 9 1 11 2 13 1 10 9 10 0 1 12 2
20 10 11 3 13 1 10 9 13 9 0 1 10 9 10 9 2 0 14 11 2
28 7 10 9 2 1 13 1 10 9 2 13 4 16 13 9 1 9 15 2 7 15 13 1 9 1 10 9 2
23 3 13 10 9 13 14 10 9 10 0 10 0 1 11 11 2 3 9 2 11 10 0 2
63 9 11 2 9 9 2 11 2 2 9 9 14 9 1 9 2 10 9 2 13 1 9 1 2 11 2 2 16 9 2 9 0 0 0 2 1 9 2 9 11 2 13 3 0 2 7 3 2 3 4 13 3 13 9 16 15 13 9 2 1 0 2 2
44 1 11 10 0 13 10 9 13 9 1 10 9 10 0 1 9 2 10 9 9 0 1 9 15 2 16 9 10 9 2 11 11 2 13 9 1 10 9 1 9 15 10 0 2
21 3 1 12 9 13 16 13 13 1 9 2 11 10 0 7 13 1 9 2 11 2
36 10 9 1 1 3 13 11 1 9 13 9 1 9 0 0 13 1 11 11 2 7 13 13 14 9 10 9 1 11 2 1 2 9 11 11 2
43 9 0 13 1 12 1 11 2 16 11 11 2 9 0 1 11 2 13 1 9 1 2 11 11 2 2 16 9 11 4 13 1 9 0 1 10 9 1 9 2 10 9 2
18 15 3 13 16 4 13 1 9 13 14 10 9 3 1 9 10 11 2
25 3 13 10 9 10 0 1 11 9 0 7 3 13 16 13 16 10 11 13 2 9 0 0 2 2
8 1 9 15 13 3 10 11 2
33 1 16 10 9 10 0 10 12 13 13 3 1 9 0 2 9 1 9 4 13 1 10 9 7 13 11 13 1 9 2 10 9 2
27 7 11 13 0 2 3 13 1 10 9 10 0 10 0 11 2 10 9 0 1 10 9 9 2 10 9 2
13 9 11 13 9 0 1 9 11 2 16 13 9 2
29 1 12 13 11 13 14 10 9 2 16 13 1 9 1 9 15 1 9 14 10 9 14 15 1 9 2 10 9 2
40 15 13 14 10 9 10 0 14 9 2 11 16 13 1 10 9 11 2 16 13 1 1 12 9 0 2 7 13 14 15 1 10 9 10 0 10 0 10 0 2
41 11 2 16 14 15 13 1 10 9 10 12 9 0 1 9 10 11 2 1 10 9 11 11 2 13 9 1 9 2 11 1 12 2 3 1 10 9 12 12 2 2
43 1 12 13 11 10 0 1 11 2 16 13 3 13 1 9 9 10 9 2 1 9 1 9 9 15 14 9 10 9 13 14 11 13 1 11 2 16 1 15 13 1 12 2
20 9 0 14 11 4 2 1 13 1 9 15 10 0 2 13 1 9 1 11 2
26 1 9 12 13 10 9 2 1 9 16 13 1 9 10 9 1 11 2 9 16 13 9 1 10 15 2
17 10 9 3 13 9 16 13 1 9 9 2 11 1 11 1 12 2
27 7 3 13 9 0 0 16 13 3 3 1 0 2 13 10 9 9 1 9 0 14 9 16 13 1 15 2
29 1 12 9 13 10 9 2 16 13 9 10 9 1 9 10 9 7 10 9 14 9 2 10 9 2 14 9 15 2
65 10 9 2 16 1 9 15 13 9 9 2 10 9 10 0 11 11 2 13 1 13 9 0 1 3 16 13 1 9 15 2 9 0 14 9 0 2 1 9 2 10 9 2 7 3 1 9 2 10 9 10 0 7 1 9 2 10 9 10 0 1 9 2 9 2
55 2 7 3 13 3 9 1 9 10 9 2 16 3 4 13 16 9 2 9 15 13 1 10 9 2 7 9 15 3 4 3 13 1 10 9 14 10 9 16 15 0 13 15 2 2 13 9 11 1 9 7 9 14 15 2
22 1 10 9 16 13 3 3 13 9 10 9 2 7 10 9 1 9 2 10 9 13 2
61 1 9 16 13 13 1 9 2 10 9 10 0 1 12 9 0 7 13 2 1 1 12 1 12 2 2 1 9 2 10 9 10 0 1 12 12 2 1 12 12 1 12 2 7 1 9 2 9 10 9 1 12 12 2 1 12 12 1 12 2 2
18 10 9 10 0 1 9 2 10 9 13 2 3 2 1 9 9 0 2
47 16 16 9 10 9 10 0 13 7 13 2 4 9 13 1 9 3 13 2 13 10 9 14 9 9 2 7 13 3 1 10 15 16 13 14 9 10 9 1 13 1 10 9 10 12 13 2
38 1 9 12 13 9 10 9 2 11 9 2 1 10 11 9 1 9 10 9 1 9 1 9 9 2 10 9 2 7 10 9 13 1 10 9 10 0 2
26 10 10 9 13 1 10 9 1 9 2 7 13 1 9 15 10 0 14 10 9 10 0 1 10 9 2
12 10 9 13 1 10 9 9 13 1 9 15 2
57 9 10 9 11 11 13 1 9 0 13 14 10 9 2 9 9 9 2 9 10 9 1 9 10 9 16 15 13 13 1 15 1 12 12 9 2 7 9 9 10 9 13 1 9 0 1 9 2 9 10 9 1 9 1 9 9 2
38 3 13 10 9 14 9 2 9 10 9 7 13 10 9 14 15 2 1 9 13 14 9 15 10 0 14 9 2 10 9 10 0 1 10 9 10 0 2
35 7 9 15 3 13 2 7 13 9 16 13 2 16 10 9 10 0 13 9 10 9 1 9 2 10 9 10 0 1 9 2 9 10 9 2
46 8 2 8 3 9 10 9 3 13 9 2 9 10 9 13 1 9 0 13 1 10 9 10 0 1 10 9 2 7 3 4 13 9 1 16 13 10 9 1 10 9 16 13 1 15 2
53 9 9 11 11 2 16 13 1 9 9 11 2 13 3 1 10 11 9 2 9 1 9 1 9 9 2 10 9 2 16 13 13 14 10 9 1 13 1 9 10 9 10 0 2 16 16 13 4 1 9 10 9 2
18 10 9 16 13 1 10 9 13 9 12 2 7 15 13 1 9 12 2
37 1 9 10 9 2 13 9 9 2 10 9 1 12 9 2 9 2 9 14 10 9 10 0 2 9 2 9 1 9 7 9 2 10 9 10 0 2
22 10 9 10 0 13 1 9 0 14 9 2 9 10 9 7 9 2 10 9 10 0 2
30 1 10 9 10 0 13 10 9 1 10 9 10 0 14 9 0 7 9 9 2 7 9 10 9 13 1 9 9 15 2
48 1 15 2 13 9 10 9 16 13 3 1 12 9 9 2 10 9 2 7 10 9 13 9 9 0 1 9 1 9 7 1 9 1 9 7 9 9 1 9 1 9 1 10 9 7 10 9 2
16 9 10 9 14 12 9 9 2 10 9 13 1 9 10 9 2
37 1 10 9 2 9 14 10 9 10 0 13 9 7 9 9 2 9 9 7 9 2 7 15 13 1 9 1 2 0 2 9 2 0 2 9 9 2
51 1 15 13 1 10 9 2 9 1 10 15 9 9 2 16 13 1 10 9 1 9 14 9 2 10 9 1 9 0 2 14 9 2 10 9 1 9 0 2 14 9 9 7 14 9 10 9 1 10 9 2
16 9 1 9 15 1 9 2 10 9 1 9 13 1 9 3 2
18 9 2 10 9 1 9 13 1 10 10 9 1 9 10 9 10 0 2
27 1 15 13 1 15 9 1 10 9 16 13 3 1 10 9 10 0 7 1 9 9 2 10 9 10 0 2
21 9 2 9 15 13 13 1 9 0 7 1 9 0 2 7 1 9 15 13 9 2
26 9 2 10 9 10 0 13 1 10 9 10 0 2 7 13 9 9 1 9 9 2 10 9 1 9 2
9 10 9 1 15 13 1 9 3 2
23 1 9 15 13 2 16 9 2 10 9 10 0 13 13 9 0 7 13 1 9 0 9 2
28 9 9 13 1 9 2 10 9 10 0 2 1 1 10 9 1 9 9 9 2 16 13 1 10 9 10 0 2
29 1 9 9 15 14 9 11 2 13 9 10 9 1 10 9 10 0 14 10 9 10 9 7 13 9 9 10 9 2
27 3 9 10 9 13 13 9 7 9 9 1 9 2 10 9 2 1 9 1 9 9 2 10 9 10 0 2
20 13 13 9 8 1 10 9 1 9 9 2 1 13 1 9 10 9 10 9 2
31 1 15 13 13 14 10 9 2 16 13 14 9 10 9 13 14 10 9 1 9 9 3 2 14 13 2 16 4 13 9 2
20 1 9 15 13 2 16 16 13 9 9 2 13 10 9 4 13 14 10 9 2
46 1 13 14 9 10 9 1 9 10 9 13 13 9 9 2 16 13 1 9 9 2 10 9 7 9 14 9 2 10 9 1 9 15 2 7 1 9 15 9 2 10 9 1 10 9 2
16 9 9 15 13 1 10 9 2 7 15 13 1 9 10 9 2
19 3 2 13 9 9 9 0 2 16 13 0 1 9 9 9 2 10 9 2
22 9 10 9 13 14 10 9 1 10 9 10 0 1 10 9 10 0 2 1 9 15 2
30 15 3 13 14 9 10 9 1 9 15 7 1 9 2 10 9 1 9 2 14 10 9 13 10 9 1 9 9 2 2
32 9 15 13 1 11 9 13 9 14 9 1 9 2 16 13 1 9 10 9 1 10 9 10 12 7 1 9 10 9 10 12 2
37 10 9 13 1 10 9 10 0 1 11 2 7 13 1 9 9 9 0 2 16 13 1 11 1 1 9 7 13 9 0 3 0 1 9 10 9 2
16 9 10 9 13 9 1 9 10 9 10 0 1 9 10 9 2
35 9 0 13 13 9 13 1 11 7 15 13 1 9 1 11 11 2 16 13 1 10 9 1 11 9 13 1 11 1 9 9 15 14 11 2
31 9 9 10 9 1 10 9 13 1 9 1 9 10 9 1 3 9 15 14 10 9 11 11 2 9 15 14 9 10 0 2
22 1 9 15 13 9 9 10 9 13 9 9 13 1 9 9 15 7 1 9 10 9 2
20 13 9 0 1 9 14 9 9 7 13 3 9 1 9 14 9 9 2 9 2
16 1 10 9 13 10 9 10 0 1 9 0 7 1 9 9 2
15 1 10 9 13 9 1 9 0 2 9 2 9 7 9 2
14 1 10 9 10 12 13 9 1 9 2 9 7 9 2
33 10 9 10 0 13 1 9 10 9 10 12 2 14 13 13 9 1 9 0 7 13 1 15 9 0 7 9 1 9 14 9 0 2
12 14 10 9 13 13 1 10 9 1 9 0 2
30 1 10 9 13 12 9 1 10 9 10 0 2 7 1 9 15 13 9 2 16 13 1 9 15 10 0 1 9 9 2
7 14 10 9 13 1 9 2
15 10 9 13 13 1 9 7 9 15 13 14 9 10 9 2
29 1 10 9 13 12 9 1 10 9 14 10 9 2 16 1 15 13 9 1 9 0 14 11 11 2 11 7 11 2
33 14 10 9 13 1 11 10 9 11 11 11 11 2 11 2 7 15 13 9 9 1 10 9 10 0 3 1 11 2 11 11 11 2
15 9 1 9 9 15 9 2 9 2 9 13 7 9 2 2
14 3 13 1 9 9 9 12 14 9 10 9 1 9 2
9 15 9 9 0 3 2 3 0 2
13 1 9 10 9 13 10 9 2 9 1 9 2 2
36 9 0 1 9 10 9 13 1 9 1 9 12 9 1 10 9 16 9 15 10 0 1 12 10 9 16 13 1 10 9 13 0 1 10 9 2
78 9 9 2 10 9 2 10 9 11 11 11 2 16 13 13 1 10 9 14 9 10 9 1 12 9 2 2 7 11 11 2 13 14 10 9 14 15 1 9 9 10 9 7 9 2 10 9 10 0 2 7 3 12 13 16 3 10 9 13 1 15 7 13 1 15 9 0 1 13 14 15 1 10 9 16 15 13 2
15 3 16 13 9 12 2 13 13 3 1 10 9 10 0 2
23 9 2 13 2 9 9 2 9 0 7 3 13 14 9 9 10 9 1 9 0 7 0 2
35 1 10 9 13 9 0 16 13 14 9 9 15 7 9 15 14 9 0 1 10 10 9 2 11 2 11 2 11 11 11 2 11 7 3 2
25 1 10 9 10 15 2 13 9 0 14 9 7 9 2 7 3 12 9 1 10 9 10 0 2 2
37 1 9 2 10 9 10 0 7 10 0 3 1 9 15 2 10 9 12 13 9 0 0 16 15 9 14 12 9 0 0 2 12 12 12 12 12 2
13 3 3 4 16 0 9 0 0 3 9 15 9 2
18 7 3 15 13 7 13 2 1 2 9 12 9 15 14 9 10 9 2
13 7 10 9 10 0 13 9 2 9 7 9 9 2
21 3 3 13 10 9 16 10 9 1 9 15 16 13 2 7 13 2 13 1 15 2
9 9 2 10 9 13 1 9 15 2
26 9 10 9 14 10 9 2 12 9 1 12 9 16 13 9 1 9 2 2 13 9 10 9 10 0 2
12 10 9 2 10 9 7 10 9 13 1 9 2
24 1 9 0 2 9 11 11 2 10 9 1 9 10 9 7 10 9 2 9 10 9 2 11 2
65 9 9 9 10 9 2 9 2 9 11 11 2 11 2 13 1 9 10 9 2 11 11 2 13 9 9 16 13 2 16 9 10 9 1 10 9 1 9 9 7 9 7 3 9 10 9 7 9 10 9 10 0 3 4 13 1 9 15 1 3 1 12 9 0 2
63 1 9 1 10 9 11 13 9 11 2 11 2 16 9 16 13 1 9 9 9 9 2 10 9 13 1 9 0 9 2 16 13 1 10 9 10 0 10 0 7 13 14 9 15 14 9 1 9 12 1 10 9 1 9 9 7 1 10 9 1 9 9 2
45 2 10 9 7 10 9 10 0 3 13 1 15 16 1 9 15 9 10 9 2 2 13 2 2 7 15 13 1 9 9 15 2 1 13 1 9 9 2 9 0 9 9 9 2 2
60 2 9 7 9 15 3 13 14 9 10 9 16 1 15 13 3 9 9 2 10 9 2 16 9 0 0 9 9 7 9 0 13 9 15 1 9 1 9 15 2 16 9 10 9 16 13 9 1 9 15 10 0 2 2 13 9 11 2 11 2
43 1 9 10 9 7 10 9 16 1 9 9 11 11 2 13 1 9 15 7 1 9 15 1 3 9 0 9 9 0 0 9 2 16 13 3 1 9 10 9 16 1 15 2
26 15 9 10 11 2 9 11 2 14 9 11 2 16 13 14 9 15 14 11 11 2 9 10 9 3 2
17 15 13 1 9 10 12 1 9 15 10 0 14 9 11 2 11 2
63 9 10 9 10 0 16 1 9 15 10 0 14 9 0 15 13 3 1 9 15 14 10 9 10 0 3 2 11 2 9 14 9 9 0 7 13 2 16 1 9 15 9 9 0 16 13 3 1 9 1 9 10 9 2 7 9 0 7 13 13 14 15 2
18 1 15 2 1 9 16 13 2 13 10 9 11 11 9 0 7 0 2
32 15 13 13 1 15 9 0 7 0 7 13 1 9 0 2 16 13 14 9 9 10 9 2 3 1 9 1 9 15 14 11 2
18 1 9 15 15 9 9 9 12 0 2 16 13 1 9 3 2 0 2
15 1 9 15 10 0 13 9 10 9 2 8 9 12 9 2
23 9 15 10 0 4 9 9 0 7 0 2 16 13 9 1 9 10 9 7 9 10 9 2
25 10 9 13 1 9 7 13 1 9 9 1 9 10 9 10 0 2 16 13 14 9 9 10 9 2
29 10 9 10 0 14 10 9 13 1 10 9 1 12 9 0 2 16 13 1 9 0 9 0 1 9 7 1 9 2
17 1 10 9 1 10 9 13 9 0 2 9 1 9 15 10 0 2
27 7 7 10 9 13 13 1 10 9 2 7 0 1 15 2 13 1 9 15 10 0 10 13 14 10 9 2
34 13 9 10 9 16 9 3 9 9 2 16 9 15 0 2 0 7 9 15 0 7 0 2 13 1 10 9 1 9 9 1 10 9 2
44 9 10 9 16 13 1 9 2 9 2 7 10 9 16 1 15 13 9 15 14 9 9 2 1 10 9 16 13 1 15 9 0 2 13 1 10 9 13 0 7 9 9 0 2
28 1 10 0 13 16 9 1 10 15 13 1 9 16 4 13 13 15 2 1 9 9 9 7 1 9 9 0 2
58 7 2 7 1 10 10 9 10 0 2 16 13 1 9 1 9 7 1 9 0 7 0 16 1 15 9 1 9 7 1 9 0 2 13 9 2 9 1 9 0 14 9 9 2 16 1 15 13 1 9 10 9 7 10 0 9 13 2
22 16 13 9 10 11 3 13 10 9 3 2 9 2 7 10 9 10 0 13 13 3 2
19 1 9 15 13 11 2 11 2 16 13 14 10 9 11 1 9 10 12 2
9 15 13 9 9 1 9 9 0 2
83 15 2 7 3 2 9 0 0 2 16 13 14 9 15 1 9 0 14 9 0 7 13 13 1 9 15 1 9 9 0 2 9 10 9 10 0 14 11 11 2 9 10 9 0 10 9 2 9 10 9 2 9 10 9 7 10 9 16 13 1 10 9 14 11 2 10 9 10 0 2 10 9 10 13 2 10 9 9 10 9 7 3 2
12 13 1 15 10 9 14 9 2 9 7 9 2
16 10 9 10 13 10 15 13 1 9 0 9 14 9 0 3 2
12 4 16 1 15 13 10 9 14 9 9 11 2
11 9 10 9 10 0 10 0 0 1 9 2
52 9 11 13 1 9 15 1 9 10 9 10 0 10 13 1 9 15 2 7 9 15 13 1 10 9 10 0 2 16 13 1 10 9 10 0 2 1 9 15 14 9 0 1 1 10 9 10 0 1 9 15 2
15 13 1 15 9 9 10 9 7 10 9 10 0 1 9 2
21 10 9 1 9 11 7 9 15 14 9 0 0 2 13 1 9 10 9 0 13 2
51 10 9 16 9 15 2 3 2 1 9 10 9 16 13 1 2 9 2 16 13 14 9 10 9 1 10 9 10 0 1 10 9 7 10 9 2 13 1 3 1 13 10 0 14 9 10 11 16 13 3 2
58 11 3 13 1 10 9 10 0 10 15 7 15 4 1 9 1 3 10 9 16 13 13 1 10 9 7 1 10 9 7 13 9 0 7 0 0 1 9 15 14 10 9 10 0 2 7 3 16 10 9 13 1 9 1 9 0 0 2
6 9 9 13 9 0 2
23 3 14 13 1 9 1 9 1 9 9 9 16 3 13 9 9 1 3 2 9 14 15 2
26 1 2 15 4 13 9 1 9 0 16 9 15 13 0 1 9 0 16 16 15 13 1 9 9 0 2
37 16 16 9 10 9 1 9 9 13 1 9 10 9 2 13 1 9 10 9 9 2 9 1 9 10 9 2 7 1 9 15 10 9 13 9 9 2
57 10 9 10 0 2 16 13 2 9 9 9 10 9 12 2 2 13 13 13 14 10 9 10 0 1 10 9 1 9 9 10 9 2 7 13 1 15 7 13 9 1 9 1 9 16 13 13 9 1 9 10 9 1 9 9 9 2
24 1 2 9 10 9 2 13 9 10 9 9 2 9 1 10 12 1 10 9 16 13 13 9 2
21 9 10 9 2 16 13 13 1 9 9 16 13 9 9 2 13 9 9 10 9 2
48 7 7 10 9 16 13 1 9 9 0 7 9 1 9 14 9 9 2 13 9 10 9 16 13 1 9 10 9 2 16 1 9 15 13 10 9 2 7 9 10 9 16 13 1 9 15 9 2
8 7 2 10 9 1 9 9 2
25 1 9 10 9 13 9 14 9 9 2 3 1 9 9 9 2 9 2 7 3 1 9 9 0 2
25 1 9 9 10 9 2 13 9 10 9 14 10 9 1 9 10 9 2 1 9 1 9 9 2 2
34 10 9 16 1 10 9 13 7 7 3 1 9 2 9 2 16 3 13 14 9 9 15 1 10 9 2 7 13 1 9 10 9 3 2
32 9 10 9 16 13 1 9 9 16 13 1 9 9 9 13 3 1 3 16 13 2 1 9 10 9 10 0 2 1 9 9 2
15 9 10 9 13 9 1 9 15 16 13 0 1 9 15 2
34 1 9 15 13 9 13 9 1 9 9 10 9 2 1 9 9 2 1 1 9 9 2 2 1 9 0 2 1 9 0 7 1 9 2
42 9 1 10 9 16 13 2 1 2 9 10 9 10 0 2 13 1 10 9 16 13 1 10 9 2 1 13 15 13 14 9 10 9 10 0 7 13 1 9 10 9 2
37 9 10 9 13 13 1 9 1 9 10 9 2 1 10 9 16 16 10 9 16 13 1 10 9 13 13 1 9 1 13 1 9 0 1 10 9 2
18 7 7 13 10 9 13 16 13 1 9 1 12 9 16 13 13 3 2
36 1 9 15 2 3 13 9 1 10 9 10 0 1 9 9 9 1 9 10 9 2 16 13 1 15 9 10 9 16 0 1 10 9 10 0 2
3 0 12 2
22 10 9 16 13 1 9 13 7 13 1 9 9 0 1 9 7 9 14 9 13 0 2
46 10 9 11 2 11 2 9 9 0 1 9 16 13 1 9 0 2 9 11 2 9 7 9 9 13 13 16 16 10 9 13 10 1 10 9 7 10 9 13 2 1 9 2 1 9 2
24 1 1 10 9 15 2 16 9 13 3 2 13 10 9 1 12 1 12 9 13 9 7 9 2
35 1 13 9 0 1 9 15 13 3 1 13 9 12 14 9 7 9 0 14 9 2 9 2 9 7 9 0 2 9 1 9 0 14 9 2
17 12 10 9 2 16 13 1 9 0 1 12 2 13 3 12 9 2
7 15 9 0 1 9 0 2
43 15 13 9 0 1 10 9 10 0 1 10 9 10 0 2 7 13 1 15 9 0 7 0 9 2 13 1 9 0 1 15 16 4 13 1 10 9 0 1 10 9 11 2
27 10 11 7 10 9 9 2 11 2 9 9 1 9 2 14 11 13 9 0 1 10 9 10 0 10 0 2
30 13 10 9 0 7 0 1 10 9 15 2 7 16 16 15 0 2 0 1 9 7 13 1 9 0 2 15 3 13 2
25 10 9 13 3 7 9 10 9 10 0 16 13 1 10 9 13 1 9 11 2 1 10 9 0 2
37 11 11 2 16 13 3 15 2 13 1 9 14 9 9 16 1 15 13 9 0 14 9 2 9 0 7 0 2 9 2 9 2 9 7 9 9 2
17 1 9 0 3 10 9 11 2 11 7 3 10 9 13 9 0 2
26 1 10 9 10 0 13 9 9 1 9 13 1 9 9 7 7 13 14 15 1 9 7 1 9 11 2
22 10 9 10 12 2 9 9 1 11 2 0 1 9 2 9 2 9 7 9 9 0 2
8 10 9 10 9 14 11 0 2
38 10 9 14 15 13 9 0 14 9 11 0 2 9 7 9 7 10 9 11 11 2 16 13 1 9 0 2 9 9 7 9 9 0 1 15 10 9 2
13 9 16 13 1 9 15 13 1 12 9 1 9 2
13 9 9 14 9 10 9 13 12 9 1 10 9 2
32 1 1 10 9 10 0 10 0 7 1 10 9 10 0 10 0 14 10 9 2 15 9 16 4 13 14 15 3 1 9 12 2
26 11 11 2 10 9 14 13 9 0 1 9 7 9 1 10 9 10 9 0 10 0 9 15 10 9 2
27 4 16 3 1 15 1 13 13 10 9 0 1 10 9 10 0 2 7 3 1 15 3 1 13 9 0 2
26 10 9 16 13 1 10 9 1 10 9 11 13 3 9 9 0 1 9 0 2 7 15 3 13 11 2
39 1 11 1 11 7 3 1 11 2 10 11 16 1 15 13 3 3 13 9 15 7 0 14 9 2 9 2 9 0 2 7 1 9 0 9 15 14 9 2
37 10 9 1 15 3 13 1 9 14 11 11 2 16 1 9 10 9 13 1 15 9 9 2 9 7 9 9 16 1 15 13 9 1 9 0 3 2
22 9 14 11 11 11 13 1 9 9 11 0 7 0 1 9 14 9 13 7 9 0 2
24 10 9 13 13 3 7 10 9 13 0 2 7 10 9 13 1 9 9 9 0 7 0 3 2
9 13 3 9 14 11 11 2 11 2
26 1 11 13 11 2 16 13 4 13 13 1 10 9 7 13 10 9 9 1 10 9 1 16 13 0 2
14 7 3 16 13 14 10 9 3 9 3 13 10 9 2
40 9 11 4 13 0 1 9 0 2 7 1 10 9 16 13 3 13 9 14 9 2 3 3 9 1 9 2 7 3 10 9 10 0 3 1 9 7 1 9 2
20 13 16 1 10 9 13 9 0 2 7 1 3 13 1 10 9 1 9 0 2
13 10 9 13 0 2 9 3 1 10 9 10 12 2
24 10 9 3 0 2 4 13 9 9 0 1 9 1 3 1 12 9 2 2 7 10 9 13 2
12 1 3 13 1 11 2 13 1 9 0 3 2
17 10 9 13 1 11 11 2 11 2 9 16 13 1 9 9 0 2
17 10 9 10 13 13 3 2 7 10 9 13 0 9 7 3 13 2
12 9 10 9 10 0 16 13 13 9 11 11 2
28 10 9 2 9 9 9 0 2 13 0 2 7 15 13 1 10 9 10 0 9 0 3 7 1 3 13 0 2
36 3 16 9 10 9 13 0 2 13 1 15 10 9 10 0 7 10 0 14 10 11 2 16 13 1 9 13 1 10 9 10 0 3 1 11 2
5 10 11 13 9 2
31 1 16 10 11 10 0 4 13 3 1 9 14 12 9 2 10 9 16 13 14 9 15 1 9 15 13 13 1 10 9 2
20 13 3 13 10 9 10 0 14 9 9 7 9 10 13 9 15 0 10 3 2
35 7 3 1 13 9 1 9 2 13 10 11 3 3 9 1 10 9 2 7 1 15 13 14 9 10 9 10 0 1 9 16 13 1 9 2
14 10 9 10 0 2 9 1 11 2 13 14 10 9 2
52 10 9 2 16 13 1 9 14 9 7 9 7 1 15 13 1 9 2 11 7 9 9 0 2 13 0 1 9 7 0 1 1 15 16 13 4 13 1 10 9 10 0 3 14 9 9 16 13 1 10 9 2
10 10 9 16 13 1 9 13 0 3 2
23 3 1 9 14 11 11 2 9 1 12 16 13 1 10 9 15 13 1 12 9 13 9 2
10 1 9 15 4 13 1 9 0 3 2
18 13 1 9 16 9 15 13 2 1 10 9 2 9 0 0 7 0 2
33 12 10 9 10 0 16 10 9 13 13 9 11 16 1 15 9 14 9 0 2 10 9 9 2 13 0 0 7 9 0 14 9 2
21 4 3 13 9 1 10 9 15 3 2 7 13 13 1 9 0 16 9 15 9 2
38 10 11 10 0 2 13 1 9 11 16 1 15 13 9 9 2 13 1 9 14 9 7 9 9 2 16 1 16 13 1 15 3 3 9 13 0 3 2
16 3 10 11 2 16 13 1 9 0 7 9 9 2 13 0 2
22 3 13 1 11 2 9 0 9 1 9 13 3 2 9 11 2 9 11 7 9 9 2
25 13 3 11 11 2 15 9 0 0 16 1 15 10 9 13 1 9 14 9 2 9 0 7 9 2
14 12 10 9 13 1 9 1 10 9 10 0 14 15 2
30 1 9 9 13 3 9 13 1 12 9 7 10 9 2 13 9 0 14 9 10 9 0 2 13 1 12 9 1 9 2
42 3 9 15 14 10 9 10 0 1 9 15 2 16 13 1 9 2 9 1 9 9 2 9 11 7 9 9 1 9 9 0 2 2 0 7 13 1 12 1 12 9 2
4 3 0 13 2
31 1 10 9 2 9 9 0 3 7 9 9 0 2 15 1 9 10 9 10 0 7 10 13 16 13 13 13 1 9 11 2
31 11 2 16 13 1 15 9 1 9 10 9 1 11 2 13 13 1 10 9 7 9 13 4 13 16 10 13 13 0 0 2
31 10 9 16 1 15 13 13 0 2 13 1 9 0 7 13 1 9 9 0 1 9 14 9 2 9 2 9 9 7 9 2
8 9 10 11 13 13 3 3 2
13 10 9 10 0 13 3 1 9 13 7 10 13 2
30 9 9 13 9 9 2 14 10 9 14 10 9 13 3 1 1 10 9 10 0 14 9 7 10 9 0 1 9 0 2
25 11 2 11 2 9 9 14 9 16 13 1 9 0 7 1 9 9 2 9 7 9 2 13 0 2
27 10 9 13 1 10 9 16 1 15 13 7 13 14 10 9 14 15 1 12 10 9 10 0 3 1 11 2
22 10 9 2 13 9 10 9 1 9 2 13 13 9 2 7 10 9 13 0 1 9 2
36 16 13 2 1 12 1 10 9 2 3 3 13 10 9 1 10 0 7 10 9 10 0 16 13 1 10 9 3 13 13 1 10 12 1 9 2
29 9 1 12 2 16 13 1 9 0 7 9 9 14 9 10 9 2 13 1 1 12 9 2 3 0 14 10 9 2
22 9 2 16 13 16 15 13 3 7 3 1 10 9 10 0 7 4 13 14 9 15 2
49 9 9 15 14 10 9 10 0 1 9 2 9 4 3 13 14 10 9 3 2 16 16 3 1 3 13 9 11 1 11 7 1 9 11 2 13 10 0 1 12 10 9 10 0 3 1 10 9 2
31 10 9 13 16 1 10 1 10 9 16 13 14 9 10 9 10 15 13 9 0 7 9 0 3 1 10 9 16 15 13 2
17 10 9 16 13 3 4 13 9 1 9 0 1 9 15 10 0 2
28 16 15 3 13 14 9 10 9 10 12 1 9 15 2 13 15 1 9 10 9 10 0 14 10 9 10 0 2
26 3 15 13 1 9 0 2 7 13 1 10 15 10 4 16 15 12 10 9 10 13 9 1 10 9 2
25 11 13 9 0 16 1 15 13 9 0 14 9 9 0 1 9 7 13 14 15 1 9 9 0 2
13 1 9 12 1 11 13 10 9 0 7 0 9 2
23 1 9 0 13 3 10 9 1 9 2 3 16 13 1 10 9 14 9 15 7 9 15 2
27 1 11 0 2 10 11 11 2 13 1 9 13 9 14 9 0 7 0 7 9 0 2 9 1 9 9 2
24 10 9 15 13 0 3 2 7 16 16 10 9 13 9 1 10 9 15 13 0 7 0 9 2
10 10 11 2 1 9 12 2 13 9 2
16 15 13 1 9 0 2 1 9 2 7 13 3 1 9 9 2
15 13 1 12 9 9 2 11 1 9 9 7 0 1 9 2
9 12 10 9 13 0 7 3 13 2
30 10 9 10 0 2 11 2 13 9 0 1 15 16 1 11 3 13 1 9 0 14 9 7 15 13 1 9 1 9 2
10 1 9 12 13 10 9 10 15 0 2
23 1 9 0 14 9 13 9 2 9 7 9 7 7 13 1 9 9 0 14 9 9 11 2
13 10 15 13 1 9 1 9 7 13 0 7 0 2
25 1 9 0 13 10 9 9 1 10 9 7 10 9 16 1 15 13 10 9 13 0 10 3 3 2
32 1 9 13 11 2 9 16 13 1 9 2 9 9 2 9 0 2 9 2 9 0 2 0 7 9 2 16 13 0 7 0 2
16 1 9 10 9 10 9 16 13 1 10 9 13 1 9 9 2
16 1 10 9 14 11 3 15 3 0 13 1 9 1 9 0 2
27 1 1 10 9 15 2 13 9 9 0 11 11 11 1 9 12 2 13 9 9 1 12 1 1 12 9 2
8 10 9 0 3 2 7 0 2
25 15 9 0 1 9 0 1 10 9 10 0 7 10 0 2 1 16 9 15 13 13 1 12 9 2
41 10 9 2 11 11 2 13 9 3 1 11 7 15 13 14 10 9 14 15 2 16 13 1 9 7 1 9 2 2 9 2 2 7 1 15 13 9 9 13 9 2
29 9 13 0 2 13 3 1 9 9 13 7 13 1 9 0 2 13 13 1 9 0 13 10 9 16 1 15 13 2
30 10 9 10 0 1 9 15 13 16 9 10 9 16 13 1 10 9 13 1 9 0 0 0 7 9 15 13 0 3 2
19 9 14 9 9 7 9 1 9 9 7 1 10 9 13 9 0 0 3 2
22 11 1 9 7 9 7 11 1 9 7 9 13 16 10 9 13 3 13 1 10 9 2
19 12 10 9 13 1 9 0 16 13 0 3 7 13 1 9 0 1 9 2
37 1 9 0 10 11 11 2 11 13 0 7 3 0 2 7 7 16 10 9 13 0 1 10 0 2 15 13 2 1 9 0 2 14 9 10 9 2
23 10 11 16 13 1 9 13 9 0 2 3 10 9 10 0 3 16 13 1 9 1 11 2
47 13 9 14 9 9 14 9 10 9 2 11 0 2 7 9 1 9 9 9 16 13 1 10 9 15 10 9 13 1 12 9 2 13 9 9 1 9 12 9 2 9 13 1 1 10 9 2
33 11 11 2 10 9 7 10 9 14 13 1 11 1 12 9 7 15 12 1 9 10 9 10 0 10 0 16 13 9 0 1 11 2
20 13 16 13 10 9 7 9 14 10 9 1 10 9 14 15 2 15 0 3 2
38 9 10 11 16 13 1 9 10 11 10 0 13 3 2 7 10 9 2 16 13 1 9 7 1 15 13 2 13 13 1 9 9 16 13 1 9 15 2
26 9 9 10 9 7 10 9 13 0 9 7 9 0 3 1 9 7 1 9 9 13 13 14 9 15 2
26 10 9 14 9 9 13 13 3 1 9 9 7 1 9 13 1 9 0 2 9 2 9 9 7 9 2
29 7 16 10 9 13 0 2 13 1 15 10 9 14 9 11 7 10 9 14 9 10 13 1 9 9 1 9 15 2
7 1 9 2 9 7 9 2
19 9 15 13 1 10 9 10 0 7 10 9 13 1 11 2 9 0 9 2
9 10 9 13 0 7 3 10 9 2
