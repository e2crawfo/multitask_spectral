489 11
5 13 10 11 11 2
17 11 2 4 13 10 9 1 10 0 9 0 1 10 11 1 9 2
30 1 10 9 0 15 13 1 13 10 9 1 10 9 2 13 16 10 9 4 3 13 1 9 10 9 1 10 9 11 2
6 0 9 1 10 11 2
7 10 0 9 10 0 9 2
34 13 9 1 13 16 10 9 0 1 9 0 2 1 9 7 1 9 0 2 4 13 9 15 13 13 9 15 15 3 4 3 3 13 2
29 15 3 15 4 3 4 13 2 16 10 10 9 13 10 9 0 2 7 10 15 3 2 10 15 13 1 10 9 2
20 10 0 2 0 9 1 10 9 0 1 10 10 2 9 2 13 1 10 9 2
33 3 11 2 13 11 2 2 13 10 9 2 1 10 0 9 2 7 2 10 9 1 11 3 13 1 13 15 1 10 10 9 2 2
5 10 9 1 11 2
57 10 9 1 10 9 2 10 9 13 3 10 9 0 1 10 11 2 13 2 0 9 2 2 7 10 9 4 4 13 1 10 9 7 10 9 0 11 11 4 13 10 9 1 10 9 1 9 1 10 9 1 10 9 1 10 11 2
45 10 0 9 10 9 2 15 13 10 9 1 9 1 11 1 10 11 2 1 11 2 4 13 15 3 1 10 9 2 16 15 13 10 9 2 7 15 3 15 15 4 13 1 13 2
48 11 11 2 0 9 1 10 11 1 11 2 9 1 9 2 12 9 2 12 1 10 15 13 1 10 9 2 2 4 4 13 1 10 10 9 10 12 9 2 1 9 1 10 9 0 11 11 2
18 10 9 1 10 9 4 13 10 9 1 3 2 15 13 3 1 11 2
31 10 9 13 1 10 9 1 10 9 0 7 3 15 1 10 11 3 0 1 10 9 4 4 13 1 10 9 1 9 0 2
30 10 11 15 13 1 9 2 10 9 2 7 2 1 10 9 0 2 1 15 4 13 1 13 15 1 10 9 2 3 2
22 12 9 1 11 2 13 1 9 10 9 2 11 2 7 9 7 12 9 2 11 2 2
7 4 13 3 10 9 3 2
21 11 2 2 9 2 4 13 1 0 9 10 10 9 7 1 15 13 16 13 3 2
14 9 7 9 13 1 10 9 1 10 9 1 10 9 2
7 11 13 1 9 1 9 2
6 7 10 9 4 13 2
24 1 10 9 4 13 10 10 9 1 10 9 0 7 1 3 1 3 13 10 9 1 10 9 2
7 3 4 4 13 10 11 2
7 13 9 1 10 9 2 2
12 10 9 1 3 11 4 13 1 10 9 2 2
6 13 1 10 10 9 2
12 10 9 15 4 13 16 11 3 15 4 13 2
16 3 4 4 13 1 15 1 10 10 0 9 2 11 11 11 2
17 7 16 15 15 4 13 1 10 10 9 2 15 1 11 11 2 2
20 10 9 4 13 2 2 1 10 9 1 9 0 2 10 9 4 13 3 0 2
34 10 9 13 1 9 10 11 13 1 10 9 1 11 2 10 0 9 4 13 1 10 11 0 1 9 7 1 13 9 1 10 0 9 2
13 7 3 15 13 1 9 7 1 9 1 10 9 2
5 15 4 13 2 2
30 9 11 4 13 10 9 1 10 10 9 0 1 13 2 0 2 10 9 1 10 9 7 13 10 9 1 10 10 9 2
14 10 9 15 4 3 13 1 10 2 9 2 1 11 2
9 2 15 15 13 10 9 9 2 2
28 10 9 1 9 3 13 10 0 9 1 10 9 7 10 9 1 10 9 0 2 7 10 9 1 10 9 0 2
14 3 3 12 9 3 13 10 9 13 1 10 9 0 2
17 2 13 1 10 0 9 1 10 9 1 11 2 2 13 10 9 2
8 2 11 2 13 15 11 2 2
26 1 15 15 15 13 2 10 9 3 4 13 10 9 1 10 0 9 0 11 11 1 10 9 1 11 2
55 1 15 2 1 9 2 15 13 12 2 9 2 2 10 9 1 10 9 1 2 11 11 2 7 1 2 11 11 2 2 15 13 10 9 1 10 12 9 2 10 0 13 1 11 2 10 0 2 12 9 3 2 1 11 2
38 4 4 13 2 1 9 1 9 2 3 1 13 9 1 9 3 0 2 12 9 15 4 13 1 10 9 2 1 10 9 0 2 10 9 1 9 0 2
23 7 10 9 3 0 4 13 15 1 11 11 2 9 1 10 11 1 10 9 1 10 11 2
15 10 9 13 1 13 9 0 1 10 9 0 10 10 9 2
16 7 16 1 9 2 13 9 9 2 0 2 0 2 0 2 2
21 10 9 0 15 16 0 13 16 10 12 3 13 9 7 13 10 9 1 10 9 2
22 10 9 1 15 2 13 3 1 10 9 2 15 4 13 3 0 9 1 9 1 9 2
13 10 10 9 7 10 10 9 3 4 4 3 13 2
9 2 4 13 10 0 1 9 3 2
8 11 13 10 9 1 12 9 2
14 3 13 3 9 1 10 9 15 13 9 1 10 9 2
42 7 10 2 0 9 2 3 13 15 2 10 9 3 4 13 1 1 11 11 2 1 15 2 13 2 2 1 9 13 1 13 3 10 9 15 13 1 13 1 15 0 2
27 1 9 2 13 7 13 0 10 9 0 1 11 11 2 15 1 10 9 1 11 15 13 1 10 9 0 2
11 7 3 15 13 1 10 2 3 0 2 2
18 7 2 16 13 10 11 2 15 4 13 10 10 9 2 15 13 2 2
10 10 9 1 10 11 1 11 11 11 2
6 11 2 10 9 0 2
25 9 2 9 1 9 2 13 1 9 1 10 9 13 1 10 9 0 1 10 9 7 1 10 9 2
15 16 3 13 2 10 0 9 13 1 9 1 10 9 0 2
34 15 13 1 13 16 2 3 1 13 15 1 10 0 9 7 1 13 10 9 1 10 10 0 9 2 11 4 13 1 9 1 10 9 2
38 13 13 16 15 13 0 1 10 9 1 9 2 3 10 9 2 15 2 16 10 10 9 13 1 9 7 10 0 9 13 2 2 13 0 7 0 2 2
13 15 13 1 13 1 10 9 10 9 1 3 3 2
11 2 1 15 10 2 11 2 4 13 3 2
23 11 11 13 1 10 9 2 1 10 9 2 1 16 15 4 13 3 15 13 3 1 3 2
18 7 1 10 10 9 13 3 1 11 7 3 3 1 10 11 1 11 2
6 15 13 0 11 11 2
21 7 13 1 15 16 15 13 9 1 10 9 1 9 15 3 13 1 10 9 13 2
36 10 9 1 10 9 3 4 13 15 15 13 10 9 9 2 16 10 9 3 13 2 1 9 2 9 7 9 7 2 16 13 2 4 13 15 2
6 10 11 1 11 11 2
15 13 1 9 10 10 9 2 11 13 1 9 10 9 11 2
11 13 10 9 1 11 1 10 0 9 2 2
10 2 7 10 9 13 3 0 2 2 2
12 13 1 10 9 1 10 9 7 1 10 9 2
10 7 13 15 15 4 13 11 7 11 2
8 7 10 9 13 1 10 11 2
35 3 13 1 10 9 1 10 12 9 2 15 1 10 11 1 11 2 12 9 12 2 13 11 11 13 10 9 1 10 9 1 10 0 11 2
58 9 15 3 13 10 9 7 15 13 3 0 16 10 10 9 2 1 10 9 1 10 0 9 2 13 13 1 10 9 2 1 10 12 9 1 9 0 15 15 13 3 9 1 15 11 3 13 2 3 0 1 10 9 1 15 3 13 2
14 3 4 13 10 9 0 2 15 4 13 1 10 9 2
9 3 10 9 4 13 10 9 0 2
11 10 9 1 11 4 13 10 9 1 9 2
18 13 10 9 0 16 11 1 10 9 3 13 16 15 13 1 10 9 2
20 10 9 1 11 2 1 9 2 4 4 13 3 1 10 0 9 2 1 12 2
8 1 10 12 10 9 1 11 2
54 10 9 3 4 13 10 9 1 9 13 1 10 11 7 1 10 11 1 10 0 9 13 1 10 9 1 10 9 2 1 10 9 1 11 7 11 2 7 13 9 1 10 9 0 13 1 15 13 1 9 11 7 11 2
19 11 11 13 13 1 10 9 1 10 9 7 3 3 1 10 10 9 0 2
15 7 13 15 3 2 16 1 13 3 13 13 1 9 11 2
40 13 3 10 9 1 9 2 1 10 15 4 13 10 9 11 11 2 1 13 1 10 0 9 1 10 9 2 1 13 1 10 9 7 1 10 9 1 10 9 2
38 16 11 13 1 10 9 2 10 9 2 1 10 9 0 3 12 9 2 0 12 7 0 3 1 12 2 4 13 1 13 1 13 1 9 10 9 0 2
20 10 9 2 10 2 11 11 2 2 4 13 1 11 7 4 13 15 1 11 2
19 11 4 13 1 9 2 0 2 1 9 1 10 0 9 2 10 9 3 2
11 9 11 4 13 3 0 1 13 12 9 2
47 9 2 9 9 1 10 11 2 10 9 13 1 10 9 2 7 3 10 0 9 1 9 2 10 9 1 11 13 1 9 1 9 2 1 10 9 1 10 9 2 1 10 9 1 10 9 2
18 13 10 9 1 9 1 9 2 1 9 1 9 3 13 0 13 2 2
24 1 10 9 1 13 2 3 15 13 1 13 16 10 9 3 13 10 9 7 13 1 13 2 2
36 1 15 2 15 1 3 10 9 13 10 0 9 2 1 0 9 13 1 10 9 0 7 10 9 0 13 1 9 2 2 15 13 1 9 0 2
17 10 11 1 10 12 1 12 15 1 10 0 2 0 9 1 9 2
32 10 11 15 13 3 9 1 11 1 10 9 1 10 9 2 16 4 13 1 9 0 10 9 1 11 3 1 10 9 1 11 2
19 15 13 11 2 13 0 7 13 10 2 9 2 1 10 9 1 10 9 2
7 15 13 1 10 0 9 2
12 1 10 12 13 10 0 9 0 1 10 11 2
29 10 3 0 13 15 13 3 1 10 9 1 10 9 1 10 9 2 10 9 15 3 1 10 12 9 13 10 9 2
54 13 1 10 0 9 2 1 10 9 0 2 16 13 10 9 1 10 9 1 10 9 0 1 10 11 2 7 1 10 10 9 13 10 9 13 1 9 2 10 11 0 2 1 10 9 15 13 10 9 2 7 15 13 2
34 13 10 9 2 10 9 2 10 9 2 10 9 0 7 0 2 10 0 9 1 10 9 2 15 13 1 10 0 9 3 1 10 9 2
12 15 13 3 9 1 9 1 0 9 1 15 2
43 10 9 1 11 2 10 0 11 2 9 1 9 0 1 9 7 1 10 9 0 2 10 9 3 1 10 9 2 9 0 7 0 2 0 9 1 10 9 7 1 10 9 2
22 11 11 2 3 2 15 4 13 1 13 10 9 1 10 0 9 1 10 9 3 0 2
25 2 9 2 1 9 0 2 2 9 2 1 9 1 10 9 2 0 7 0 2 9 1 9 0 2
27 0 3 10 9 1 2 11 2 2 10 9 1 9 7 9 1 10 9 15 13 1 10 13 1 10 9 2
17 16 15 13 1 9 1 9 3 15 4 3 13 10 9 1 11 2
12 10 0 1 10 9 2 10 15 1 10 9 2
19 3 1 10 9 0 2 13 9 1 10 9 2 3 1 0 9 1 9 2
35 13 10 0 9 1 10 9 2 13 0 7 0 2 13 3 3 1 10 9 7 3 3 13 9 1 9 1 9 15 13 10 9 0 2 2
33 16 13 10 9 0 13 10 9 1 10 9 0 2 11 1 10 9 2 1 11 11 2 15 13 10 9 7 10 9 1 10 9 2
30 10 9 2 3 2 13 3 15 1 16 13 1 10 9 3 16 15 13 9 1 3 13 3 0 1 2 13 15 2 2
20 15 13 10 9 13 10 9 0 7 10 9 0 13 9 7 9 1 10 9 2
8 13 1 10 9 10 0 9 2
21 13 10 9 3 0 1 3 12 9 7 15 1 3 1 12 13 1 9 1 11 2
18 3 2 3 2 16 3 13 4 15 13 1 13 2 4 13 10 9 2
37 7 13 3 11 11 2 10 9 0 1 10 10 9 2 1 11 2 4 13 10 9 1 11 11 7 10 11 2 7 15 13 9 1 9 10 9 2
45 10 9 1 10 9 0 0 7 9 1 9 2 1 9 9 9 2 13 3 0 1 10 10 0 12 9 1 9 2 7 4 13 1 10 9 1 10 9 1 10 3 0 1 9 2
46 1 9 0 9 7 9 1 9 2 10 9 1 9 4 13 10 9 2 9 1 10 0 9 1 10 9 7 1 10 9 2 2 3 1 15 15 13 1 13 9 7 9 1 0 9 2
5 0 9 3 0 2
36 1 10 13 1 9 1 10 9 0 10 9 1 9 13 3 7 1 10 9 13 1 10 9 10 9 1 10 9 9 13 0 1 10 9 0 2
7 10 9 0 2 10 9 2
22 4 13 1 12 2 12 9 1 10 9 7 4 13 1 10 9 1 13 15 3 12 2
45 2 1 10 9 1 11 4 4 13 10 9 1 9 1 10 10 9 2 13 16 10 9 2 9 1 10 0 9 2 4 13 3 0 2 3 1 10 15 0 3 1 10 9 0 2
18 13 16 4 4 13 10 9 0 1 10 15 4 3 13 10 9 0 2
24 1 15 10 2 13 2 3 13 1 13 10 9 1 9 2 3 13 9 0 1 10 9 0 2
22 10 10 9 4 13 1 15 1 9 2 13 1 9 1 9 2 9 1 9 7 9 2
4 0 13 15 2
19 13 10 9 3 1 12 9 3 7 15 13 3 1 10 9 1 10 9 2
38 10 2 11 1 10 9 2 13 10 9 1 10 9 1 10 11 2 13 1 10 0 9 2 3 1 9 1 10 0 9 0 1 15 4 13 10 9 2
24 1 3 13 3 15 15 13 10 9 15 2 1 10 12 1 9 2 13 3 1 10 10 9 2
18 1 11 2 3 2 15 4 3 13 10 9 7 10 9 1 9 0 2
17 1 10 9 1 9 10 9 15 13 2 1 0 9 2 10 9 2
15 10 9 2 1 3 13 7 13 10 9 1 10 9 0 2
7 9 2 13 12 2 2 2
9 10 9 4 13 1 10 9 0 2
58 10 9 13 10 9 1 9 2 0 3 1 10 0 9 1 10 9 2 7 1 10 0 9 1 10 9 1 9 1 10 9 2 7 1 10 9 15 10 0 9 4 13 1 10 9 0 2 1 10 9 7 1 10 9 1 10 9 2
10 12 2 9 7 9 1 10 9 13 2
22 10 9 1 9 0 1 10 9 1 10 9 13 1 10 9 0 4 13 1 9 0 2
54 16 10 9 4 13 15 2 12 2 1 10 9 13 1 10 9 3 1 13 15 10 9 1 10 10 9 2 3 13 10 9 1 13 15 0 1 9 1 10 9 12 2 7 4 13 10 9 2 12 2 1 10 9 2
15 10 9 4 3 13 9 0 1 9 1 15 1 10 9 2
27 10 9 2 12 2 3 13 10 9 1 10 9 1 10 9 7 9 1 15 4 13 9 1 10 9 0 2
34 10 9 4 2 12 2 13 10 9 0 2 7 13 1 10 9 10 10 9 1 9 7 9 2 12 2 1 10 9 13 2 12 2 2
12 12 2 9 1 9 2 9 2 9 7 9 2
7 12 2 9 1 10 9 2
10 10 9 13 1 12 9 15 13 0 2
67 16 1 9 1 10 9 15 4 13 1 9 1 9 1 10 9 2 1 9 1 9 7 1 9 1 9 2 10 9 0 2 1 9 1 10 9 1 10 0 7 3 1 9 2 4 13 10 9 1 10 9 1 10 9 15 13 9 1 10 9 0 2 12 2 12 2 2
33 10 9 15 1 9 13 1 10 9 10 13 1 0 13 10 10 9 2 3 16 10 9 13 10 9 1 10 9 2 13 12 2 2
45 10 9 4 13 10 9 1 13 7 13 1 10 1 3 1 10 9 10 9 1 9 1 15 2 15 15 13 10 9 2 12 2 12 9 12 2 12 9 12 2 12 9 12 2 2
48 3 2 13 0 10 9 1 9 0 2 0 1 9 2 13 12 2 2 1 15 1 10 9 15 13 10 9 1 10 9 1 9 1 13 15 10 9 1 15 13 1 1 10 9 1 10 9 2
9 12 2 9 1 10 9 1 9 2
23 10 9 1 10 9 15 13 1 9 1 10 3 9 13 1 12 9 2 12 7 0 2 2
27 10 9 13 10 9 1 13 10 9 1 10 9 1 15 13 10 9 2 1 15 4 13 1 10 9 12 2
26 10 9 13 9 1 10 9 1 10 9 15 13 1 10 9 1 10 9 1 10 9 2 9 12 2 2
30 16 10 9 3 4 13 15 1 9 1 10 9 7 13 9 1 15 15 13 10 9 0 1 10 9 2 9 12 2 2
17 10 9 4 13 15 1 15 3 1 10 9 15 13 1 10 9 2
33 10 9 4 13 10 9 15 13 9 1 10 10 9 2 1 10 9 1 10 9 2 1 15 4 13 1 10 9 12 2 12 2 2
48 10 9 1 10 9 7 1 10 9 1 9 2 12 2 4 13 1 13 1 9 2 7 1 9 1 10 9 2 10 9 7 10 9 1 10 9 7 1 10 9 1 15 10 9 0 4 13 2
7 12 2 9 1 10 9 2
26 16 4 13 10 9 7 10 9 13 1 13 15 1 10 9 13 1 9 2 10 9 3 4 13 15 2
23 16 10 9 4 13 7 13 1 0 9 2 10 9 15 13 1 10 9 0 2 12 2 2
5 1 10 9 0 2
28 10 9 0 13 1 10 9 13 1 10 9 1 10 9 1 10 0 9 13 1 10 9 2 12 2 12 2 2
10 12 2 9 1 10 9 1 10 9 2
8 12 2 9 1 10 9 0 2
16 16 10 9 4 13 1 9 2 10 9 13 1 10 9 0 2
5 12 2 9 0 2
15 10 9 13 1 10 9 1 15 15 4 13 1 13 15 2
35 10 9 13 1 10 9 1 10 9 0 13 16 10 9 15 13 1 9 1 10 9 2 1 9 7 1 9 2 12 2 12 2 12 2 2
11 1 10 9 1 9 7 1 9 1 9 2
29 16 15 13 1 9 13 1 13 10 9 1 9 0 2 10 9 4 13 1 9 1 10 9 15 15 4 13 15 2
28 10 9 15 13 9 1 10 9 4 13 0 1 9 0 7 4 13 1 10 9 2 3 3 0 1 10 9 2
18 1 10 13 10 9 10 9 4 13 10 9 1 10 0 9 1 9 2
14 1 10 9 10 9 15 13 16 10 0 9 4 13 2
40 10 9 13 1 9 16 2 1 10 9 0 2 3 13 10 9 13 15 1 10 9 13 1 10 9 0 7 3 13 15 13 0 16 10 9 4 13 10 9 2
43 1 10 9 15 13 1 9 10 9 1 9 2 4 13 1 10 9 1 10 9 10 9 0 2 3 16 3 4 13 3 7 3 16 10 9 3 13 1 4 13 10 9 2
32 10 9 0 1 10 9 0 1 10 9 2 13 1 10 9 1 10 9 2 13 9 1 10 9 3 1 1 10 9 1 9 2
17 3 16 10 0 9 4 13 10 9 2 15 13 13 1 10 9 2
25 10 9 3 15 13 1 9 1 10 15 15 4 13 9 1 9 7 1 9 1 15 1 10 9 2
14 10 9 13 9 0 1 10 9 7 9 1 10 9 2
12 10 9 3 4 13 9 3 1 10 9 0 2
30 10 9 13 1 9 0 7 0 9 10 9 1 10 9 7 10 9 1 10 9 0 2 1 0 9 1 10 9 0 2
16 10 0 7 10 0 13 9 1 10 9 7 1 10 9 0 2
32 10 9 1 9 3 4 4 13 16 3 1 9 0 7 1 9 1 9 0 0 7 1 10 9 1 9 0 13 1 10 9 2
18 1 10 9 1 9 1 10 9 3 15 4 13 0 9 7 0 9 2
26 10 9 15 13 9 0 7 10 15 13 1 10 9 4 13 3 1 10 9 1 10 9 1 10 9 2
34 10 9 1 10 9 2 3 1 13 10 10 9 2 13 9 1 9 1 10 9 7 1 9 1 10 9 3 1 10 9 1 9 0 2
30 10 9 1 10 9 1 10 9 7 10 9 2 3 1 13 10 9 2 13 9 1 10 9 1 10 9 1 10 9 2
23 1 10 9 1 10 9 4 13 10 9 1 9 2 10 9 7 10 9 0 1 10 9 2
43 10 9 1 9 7 10 0 9 1 9 0 13 9 1 10 9 1 10 9 1 10 0 9 1 10 9 0 7 2 1 0 9 13 1 10 9 2 3 1 10 9 0 2
41 10 9 1 10 9 3 4 4 13 1 10 9 1 9 13 1 15 2 1 0 9 2 15 4 3 3 13 1 10 9 1 9 1 10 9 7 1 10 10 9 2
12 10 9 13 13 7 13 10 9 1 10 9 2
29 10 9 1 10 9 4 13 10 9 1 9 0 1 10 9 0 3 1 10 9 0 1 12 9 1 10 10 9 2
33 10 9 0 13 10 9 2 10 9 2 10 9 1 9 1 10 9 1 9 0 2 7 10 9 1 9 1 10 9 1 10 9 2
19 1 9 0 4 13 10 0 9 0 1 10 9 7 10 9 1 10 9 2
47 1 10 9 1 10 11 2 11 11 2 1 15 1 10 9 12 2 15 13 3 10 9 0 1 10 9 0 1 10 9 0 2 0 13 10 9 1 10 9 0 1 9 1 10 9 12 2
33 1 10 9 1 9 1 10 9 15 13 1 13 1 9 10 9 0 0 12 9 12 2 9 12 2 1 10 9 0 1 10 9 2
62 3 1 10 9 1 10 9 1 10 0 9 2 10 9 0 4 4 13 2 16 15 13 9 1 13 1 10 9 13 1 10 10 9 1 10 9 12 2 0 7 0 9 2 7 12 2 9 0 7 0 2 1 10 9 0 12 9 12 2 9 12 2
24 10 9 4 4 3 13 1 9 0 1 10 9 1 10 10 9 7 1 10 9 1 10 9 2
35 2 12 2 1 9 0 2 10 9 0 1 10 9 15 13 9 1 9 7 16 4 13 4 4 13 1 10 9 0 1 10 10 0 9 2
33 2 10 9 4 4 13 1 3 12 9 1 10 0 9 1 9 0 2 12 9 1 11 1 10 9 2 7 10 0 9 7 9 2
30 10 9 1 10 9 4 13 1 10 9 1 9 7 1 9 15 13 3 10 9 3 1 9 13 1 10 0 9 0 2
22 8 2 10 9 0 0 13 1 10 9 1 9 4 13 1 10 9 0 1 10 9 2
32 3 10 9 4 13 10 9 0 1 11 15 1 10 12 10 9 0 1 11 15 13 3 1 10 9 0 1 10 9 1 11 2
15 15 13 10 9 1 10 9 1 10 9 1 10 9 0 2
14 16 4 13 1 10 9 2 15 13 12 9 1 9 2
21 15 13 16 15 13 10 9 0 1 10 9 1 11 7 1 10 9 1 10 9 2
10 7 10 9 1 10 9 3 4 13 2
11 11 11 4 13 10 9 0 1 10 9 2
13 3 1 9 4 13 10 9 1 10 12 1 12 2
20 10 9 4 13 1 10 9 1 10 11 1 10 9 1 10 9 1 10 11 2
30 3 13 10 9 1 15 13 10 9 13 1 10 9 1 12 12 9 7 2 3 2 1 10 12 7 10 12 12 9 2
5 13 10 9 0 2
80 16 11 15 13 13 1 9 1 10 9 13 1 10 2 9 0 2 2 1 15 1 10 12 9 1 10 9 0 1 10 9 0 11 2 9 1 9 1 10 9 1 10 9 1 9 1 10 11 2 11 2 2 13 10 0 9 0 7 15 13 13 10 9 0 11 2 11 2 7 10 9 1 9 1 10 0 0 9 0 2
27 10 9 13 10 12 5 1 10 9 1 10 9 0 15 13 1 10 9 0 1 10 11 7 3 1 15 2
31 11 11 2 9 7 9 2 13 10 9 1 9 1 10 9 0 7 1 11 10 9 1 11 7 3 10 9 0 13 0 2
21 10 9 1 9 2 12 9 2 10 9 1 10 9 13 1 10 9 1 10 9 2
35 1 11 15 13 10 3 0 9 1 9 1 11 1 9 0 15 13 1 10 9 1 11 9 13 12 9 1 10 9 1 10 9 1 11 2
16 15 4 13 3 2 16 13 0 7 0 13 15 16 13 15 2
72 11 2 11 7 10 9 13 1 9 7 10 9 0 1 13 15 4 3 13 2 13 10 9 1 10 9 11 11 2 15 15 13 13 3 1 10 0 9 1 10 9 1 11 11 2 13 1 0 12 9 1 10 9 3 0 7 13 1 10 9 0 2 9 1 10 13 9 1 10 9 0 2
27 1 10 9 7 10 9 1 9 3 1 10 9 2 10 9 1 10 9 1 10 9 4 4 13 7 13 2
7 9 1 13 9 0 0 2
19 10 0 9 2 1 0 9 1 10 9 0 2 4 13 10 9 1 9 2
51 7 1 9 1 10 13 15 1 10 9 1 11 2 15 13 16 10 11 4 13 3 1 13 1 10 3 13 9 11 11 10 9 1 10 9 2 1 9 0 2 1 10 9 3 0 1 10 9 0 0 2
37 10 0 9 4 4 13 1 10 9 1 10 9 1 10 9 2 11 11 11 2 1 13 10 9 0 1 10 9 0 2 15 13 9 3 1 11 2
11 2 10 9 1 10 9 13 10 15 2 2
26 9 0 1 11 1 10 9 15 1 10 9 0 13 10 0 9 0 1 10 9 2 9 13 10 9 2
38 10 9 1 3 12 9 2 13 3 1 10 0 9 3 9 0 4 13 10 9 3 0 2 3 4 4 3 13 1 10 9 2 1 13 1 9 0 2
45 1 10 8 8 11 13 3 13 10 9 1 10 11 2 10 9 0 1 10 0 9 0 15 1 10 9 1 10 9 0 1 11 11 13 1 10 9 12 9 1 12 9 1 9 2
7 10 9 0 13 10 9 2
61 1 12 12 2 10 9 1 12 2 4 13 1 10 9 0 1 10 9 1 9 0 1 10 9 13 1 10 12 5 1 10 12 5 2 1 10 9 1 15 10 9 0 13 1 10 12 5 10 9 7 10 9 0 8 8 3 13 10 12 9 2
39 10 9 2 13 1 10 9 9 9 0 1 11 7 1 10 9 0 1 10 9 1 9 1 11 7 11 11 4 4 13 1 10 9 1 10 9 1 11 2
42 15 4 13 9 1 10 13 10 9 1 10 12 2 12 2 13 15 1 10 9 1 10 9 11 2 3 1 10 9 2 1 10 9 13 16 10 9 4 13 1 9 2
14 15 15 13 10 9 15 13 1 10 9 1 10 9 2
38 4 13 3 10 0 9 16 11 4 13 1 9 1 9 1 10 9 1 9 1 10 9 0 2 3 11 11 13 3 1 10 9 1 10 9 1 9 2
34 1 10 12 15 13 10 9 1 10 9 9 2 10 11 2 7 2 3 1 10 9 0 2 10 0 9 13 1 9 1 10 12 9 2
11 3 10 9 1 10 9 4 13 10 9 2
26 10 9 15 4 13 9 1 10 0 9 2 9 1 10 9 2 1 10 11 0 1 11 1 10 9 2
12 11 7 11 1 9 1 10 9 1 10 0 2
43 7 10 9 1 3 13 10 9 2 15 1 10 9 1 10 9 1 10 9 1 10 10 9 0 2 13 1 12 9 2 0 2 2 1 10 9 1 13 3 10 9 0 2
9 2 3 13 9 0 2 2 13 2
74 7 15 15 13 1 10 9 3 15 13 1 10 9 7 15 13 3 1 13 15 3 16 15 4 13 10 0 9 1 11 2 0 1 10 9 0 2 13 1 10 10 0 9 1 9 0 2 1 9 0 2 1 9 1 9 7 1 0 9 2 9 7 9 2 8 8 2 1 10 9 1 10 9 2
49 1 10 9 15 13 1 9 0 2 1 9 1 10 9 1 10 9 7 1 10 9 0 15 10 0 9 4 13 10 9 1 13 1 10 9 1 9 1 10 9 1 10 9 15 13 10 9 0 2
36 3 1 11 11 10 0 1 10 9 15 13 9 15 15 13 0 2 15 15 3 13 10 9 16 13 2 15 15 16 13 15 13 3 1 9 2
43 13 1 10 10 0 9 2 0 9 11 2 2 13 1 10 9 9 1 11 11 2 3 1 10 9 13 2 10 9 1 10 9 0 7 0 15 3 4 3 13 10 9 2
37 7 13 16 1 9 11 13 9 1 9 3 3 1 11 2 7 1 10 10 0 9 0 1 9 13 3 1 11 2 3 16 10 10 9 13 9 2
7 13 10 0 9 7 9 2
16 9 1 9 1 10 11 1 10 9 1 10 9 0 7 0 2
28 1 10 9 1 10 9 0 15 13 10 9 15 3 15 13 1 11 11 2 1 15 1 11 11 2 7 11 2
7 9 1 10 9 1 9 2
35 1 12 9 1 9 2 3 2 4 4 13 15 15 1 2 11 11 0 2 2 3 1 10 11 11 2 15 4 13 1 12 9 12 9 2
35 3 1 13 15 13 10 9 1 9 0 1 10 9 7 10 0 0 9 1 10 9 11 11 2 15 13 10 9 1 9 1 10 9 0 2
29 16 10 0 9 15 13 10 9 16 1 10 9 4 13 10 9 1 9 7 15 4 13 1 13 15 1 10 9 2
15 10 12 9 10 9 4 13 1 13 1 10 9 1 9 2
63 7 3 11 2 13 1 11 1 10 9 11 11 3 3 1 13 9 7 3 1 13 10 3 0 1 10 9 1 13 10 9 0 0 1 10 9 1 13 10 9 1 10 9 7 13 15 3 1 9 10 0 9 0 1 9 3 0 2 13 10 10 9 2
37 10 12 9 12 4 13 1 9 1 11 11 1 10 9 1 10 9 2 3 13 2 1 10 9 1 10 11 1 10 9 1 10 9 1 11 11 2
20 10 12 9 0 7 10 12 9 15 13 10 9 13 3 9 1 10 0 9 2
81 1 10 12 1 11 13 1 9 1 10 9 0 1 10 9 1 11 11 10 9 2 3 1 10 9 0 13 1 10 9 2 15 13 1 10 9 2 10 9 1 0 9 0 2 15 13 10 0 9 1 10 9 0 1 10 9 0 2 13 10 9 1 10 9 7 1 10 9 0 13 10 9 3 1 11 11 7 11 11 11 2
72 15 4 13 1 10 9 0 1 10 9 0 1 10 9 7 1 10 9 7 1 10 9 0 7 0 1 10 9 2 16 4 13 3 1 10 9 1 10 9 1 10 9 1 10 9 13 2 0 7 0 2 7 1 10 9 1 9 0 7 1 10 9 1 9 0 7 0 13 1 10 9 2
26 1 10 12 10 9 3 4 3 4 13 1 10 0 2 0 9 9 9 2 13 10 9 1 10 9 2
31 1 9 10 9 13 1 9 3 3 0 2 13 10 9 0 7 0 1 9 3 0 2 0 2 1 3 9 1 9 0 2
28 10 9 13 10 0 9 2 7 13 10 9 2 1 15 13 10 0 9 7 15 15 13 1 4 13 10 9 2
22 10 9 1 10 9 13 1 13 13 0 9 0 1 10 9 9 2 13 1 10 9 2
12 10 10 0 9 1 10 9 13 1 13 3 2
51 10 0 9 1 10 9 13 1 10 9 1 2 9 9 2 2 1 9 3 13 9 1 9 1 10 9 1 9 2 7 15 13 1 13 10 9 2 13 10 9 15 13 1 10 9 0 1 10 9 0 2
40 11 13 10 9 1 10 12 2 1 10 0 9 1 10 0 9 1 10 11 1 10 9 2 1 9 1 11 11 11 2 9 1 11 7 9 1 10 9 0 2
23 10 10 0 9 4 3 13 1 10 9 1 10 12 2 13 1 10 9 1 10 9 0 2
50 10 9 0 4 3 13 9 0 7 9 1 11 11 16 3 0 1 10 9 0 7 0 2 16 13 3 1 10 9 1 11 11 2 10 0 9 1 9 0 4 13 3 1 10 12 1 11 11 2 2
23 11 2 8 4 13 3 1 11 2 11 2 2 11 7 11 2 2 13 10 10 9 0 2
55 3 10 9 1 11 1 13 10 9 1 10 11 1 10 9 1 0 9 1 10 9 1 11 15 13 10 9 3 0 1 9 1 10 0 13 15 1 10 9 9 9 7 10 9 1 9 1 10 9 1 9 1 0 9 2
53 10 9 0 1 10 0 9 1 9 1 9 0 13 10 0 9 1 9 7 9 2 11 2 2 10 9 1 9 9 2 9 2 2 10 0 9 0 9 2 11 2 7 10 11 2 11 11 9 9 2 11 2 2
10 10 9 1 10 10 9 4 13 9 2
11 10 9 15 15 13 15 13 9 1 9 2
17 4 13 3 1 9 7 13 10 9 0 2 9 1 10 0 9 2
28 10 9 2 15 13 9 2 9 7 10 0 9 13 2 4 13 1 9 9 0 2 1 11 7 11 1 9 2
23 10 0 9 4 13 1 10 9 7 1 15 13 1 10 9 16 4 13 1 9 10 9 2
25 13 16 10 9 1 9 0 1 10 9 1 9 13 1 10 9 7 1 10 9 7 1 10 9 2
14 3 4 4 13 10 9 11 1 10 9 1 11 11 2
6 3 15 13 10 11 2
5 15 13 11 11 2
6 3 15 13 10 9 2
9 1 10 9 13 10 9 1 9 2
6 3 13 10 9 0 2
11 1 10 15 4 13 10 9 1 9 0 2
13 15 13 10 9 1 10 9 1 2 11 11 2 2
7 1 10 9 13 10 9 2
8 15 13 10 9 1 11 11 2
10 10 15 4 13 10 2 9 11 2 2
11 15 15 4 13 1 10 2 11 11 2 2
9 10 15 4 13 10 11 11 11 2
12 10 9 13 10 9 1 10 9 1 10 11 2
12 15 13 10 9 1 10 11 11 1 10 12 2
11 1 10 9 0 15 13 10 9 1 11 2
11 15 13 10 9 1 10 9 1 9 11 2
11 15 13 10 9 1 10 9 1 11 11 2
16 3 15 13 10 9 1 11 11 2 10 0 9 1 10 11 2
11 13 10 9 1 15 1 10 9 1 11 2
5 15 13 11 11 2
7 10 15 4 13 10 11 2
13 10 9 1 10 9 1 10 11 4 13 1 11 2
13 3 15 4 3 13 12 9 1 10 11 11 11 2
11 15 13 10 9 1 10 9 11 1 11 2
9 3 15 13 10 9 1 11 11 2
10 1 10 9 11 11 4 13 0 9 2
15 10 9 4 4 13 1 10 11 0 1 10 9 1 11 2
6 10 9 13 11 11 2
9 1 10 9 0 13 9 11 11 2
9 15 13 10 9 1 11 1 11 2
9 15 13 10 9 1 10 9 0 2
5 3 13 11 11 2
12 10 0 9 1 10 11 11 13 10 9 0 2
19 10 9 2 1 10 10 11 2 13 9 1 9 1 13 10 0 11 11 2
9 15 13 10 9 1 10 11 11 2
12 15 13 10 9 1 10 11 1 10 11 11 2
7 3 13 10 9 1 11 2
9 15 13 10 11 1 10 11 0 2
8 3 11 11 13 1 10 11 2
11 10 11 11 0 15 13 1 10 9 12 2
11 3 4 13 10 9 11 11 1 10 12 2
17 3 4 4 13 10 9 2 11 1 11 2 2 2 11 2 2 2
7 13 10 9 1 10 11 2
14 10 9 13 1 10 9 0 1 10 12 1 10 11 2
8 3 10 11 11 13 10 11 2
7 15 13 0 10 9 11 2
8 3 15 13 10 9 1 11 2
15 10 9 4 3 0 1 10 9 1 10 9 1 10 9 2
7 3 4 13 10 0 11 2
16 10 9 1 11 13 1 10 12 1 10 9 1 10 11 11 2
11 3 15 13 10 9 3 0 1 10 11 2
8 15 13 10 9 0 1 11 2
6 15 13 0 11 11 2
15 15 13 10 9 1 10 3 0 9 1 9 1 10 9 2
8 1 10 9 4 13 10 11 2
8 15 13 9 1 10 11 11 2
9 15 13 10 9 1 10 9 0 2
9 3 15 13 10 9 13 1 11 2
9 3 15 13 10 9 0 1 11 2
9 15 13 10 9 0 1 10 9 2
19 3 15 13 10 0 9 1 9 13 1 9 15 15 13 10 9 1 11 2
10 3 15 13 16 13 10 9 0 0 2
9 3 13 2 9 0 2 1 9 2
15 10 9 13 1 10 12 10 9 1 11 11 2 11 2 2
9 3 15 13 2 9 2 1 0 2
6 15 13 0 10 9 2
8 3 4 13 10 9 1 9 2
15 1 10 9 4 13 11 11 2 10 9 1 10 11 11 2
8 10 9 4 13 1 10 12 2
8 15 13 10 9 1 10 11 2
8 13 3 15 13 10 9 11 2
5 15 13 11 11 2
8 15 13 10 9 1 10 11 2
8 10 9 4 13 10 9 0 2
13 10 9 13 10 9 1 9 15 13 1 10 9 2
13 3 4 13 10 9 13 1 10 12 1 10 12 2
11 15 13 10 9 1 10 9 1 10 11 2
9 15 13 10 9 1 10 0 9 2
24 13 10 0 15 4 13 10 9 1 11 11 1 9 1 9 1 10 2 11 11 2 1 11 2
11 10 0 13 10 9 0 0 1 15 0 2
12 15 13 10 9 1 10 2 11 11 11 2 2
14 1 10 9 13 10 9 1 9 3 0 2 11 2 2
10 10 9 4 13 10 0 9 11 11 2
15 1 10 9 0 15 13 10 0 9 1 9 1 9 0 2
13 1 10 9 4 13 10 12 9 1 10 9 0 2
7 1 10 9 13 10 11 2
6 10 15 13 10 11 2
10 1 10 9 13 10 9 1 11 11 2
10 3 11 15 13 13 10 11 1 11 2
9 1 10 9 10 11 13 10 9 2
10 1 10 9 15 13 10 2 9 2 2
9 10 9 13 10 9 0 1 9 2
7 1 10 9 13 11 11 2
5 15 13 11 11 2
9 1 10 9 4 13 10 11 11 2
9 1 15 13 10 2 9 2 0 2
7 3 15 13 10 11 11 2
7 10 9 13 10 11 11 2
15 10 9 13 10 9 1 11 1 10 2 11 1 11 2 2
6 15 4 13 10 11 2
8 1 15 13 10 11 1 13 2
7 10 15 4 13 10 9 2
6 15 4 13 10 9 2
7 15 4 13 1 10 11 2
6 10 15 13 10 9 2
5 1 15 4 13 2
8 3 10 11 4 13 10 9 2
76 1 10 9 1 9 7 9 1 9 2 10 9 9 1 11 2 11 11 2 4 13 10 9 1 9 1 10 0 9 0 1 10 11 11 11 11 2 9 1 11 1 3 12 9 2 1 9 1 10 9 1 9 1 10 11 1 10 9 0 1 10 9 1 11 7 11 2 13 1 10 12 9 1 10 11 2
9 1 10 9 11 11 7 11 11 2
71 7 10 9 2 1 10 9 1 11 2 13 9 1 10 9 2 7 13 1 15 16 11 11 2 10 9 1 10 9 0 2 4 4 13 1 10 9 1 10 9 1 10 9 1 11 1 9 0 1 10 9 1 10 9 1 10 0 9 15 10 9 1 11 11 4 13 1 10 0 9 2
15 1 10 0 9 11 10 9 0 13 10 9 1 9 0 2
26 4 3 13 1 11 2 3 10 9 4 13 10 9 1 13 10 9 3 3 1 9 7 10 10 9 2
31 3 16 10 9 13 3 10 9 1 11 2 11 11 2 13 1 10 9 1 10 0 9 2 3 13 1 11 1 11 11 2
16 7 3 13 16 1 11 4 4 13 3 10 9 1 11 11 2
19 10 12 9 2 1 15 11 11 2 9 1 11 2 4 13 1 9 0 2
30 13 9 1 15 10 9 11 1 10 9 1 15 1 10 9 1 11 2 11 11 2 13 1 9 1 9 7 1 9 2
13 2 1 10 9 4 13 10 9 0 1 10 9 2
16 3 4 3 13 1 0 9 0 7 1 10 10 9 1 9 2
30 3 2 2 4 13 11 2 15 4 13 1 9 13 0 9 2 7 15 13 0 2 1 10 9 7 1 10 9 2 2
46 10 9 1 10 9 2 3 2 4 13 10 10 9 7 2 3 1 10 9 0 2 4 4 13 3 10 9 1 10 9 7 15 1 10 9 1 9 15 4 13 10 9 1 10 9 2
11 11 13 0 12 5 1 11 1 12 9 2
14 1 10 0 9 10 9 1 10 9 1 11 11 11 2
13 3 13 9 3 0 1 13 10 12 2 2 13 2
19 0 9 2 3 2 15 4 13 1 10 9 1 9 1 10 9 1 11 2
12 9 2 13 1 10 0 9 12 2 11 2 2
25 10 9 1 10 9 15 3 4 13 1 10 9 1 10 0 9 7 1 10 9 1 9 4 13 2
13 9 1 10 9 1 10 9 1 10 9 1 9 2
117 1 16 4 3 13 3 1 9 1 10 9 2 10 11 13 10 9 1 9 2 3 16 13 2 7 3 13 10 9 7 9 1 10 9 1 9 1 10 9 2 13 15 0 7 0 2 1 9 0 7 1 0 9 2 13 3 13 2 1 10 15 2 10 9 0 1 10 9 2 1 10 9 2 1 10 9 1 10 9 0 7 1 10 3 9 1 9 1 15 7 1 10 9 1 9 0 7 1 0 9 2 1 10 9 7 1 10 9 1 9 2 13 15 0 7 3 2
19 11 11 3 13 9 1 10 0 9 7 3 13 10 9 13 1 10 9 2
19 3 2 9 11 2 13 16 10 9 1 10 9 15 15 13 13 3 0 2
13 13 16 4 13 10 9 2 1 3 3 13 3 2
58 1 15 2 10 0 9 13 13 1 10 10 9 1 9 2 1 1 13 10 9 0 2 10 9 3 0 15 13 1 10 13 1 9 1 10 9 0 10 9 0 1 10 9 10 9 3 2 7 3 10 9 3 2 16 4 4 13 2
26 16 13 0 2 10 9 13 1 10 9 1 9 0 1 10 9 1 10 9 13 1 10 10 9 0 2
46 15 13 16 10 10 9 0 2 1 9 1 10 3 9 2 15 3 3 13 10 9 0 2 2 13 0 7 16 10 0 9 13 1 10 9 1 13 16 13 1 10 9 1 10 9 2
74 1 0 10 9 1 10 9 1 10 9 4 13 3 1 10 9 1 10 9 1 10 8 8 1 10 9 0 1 10 9 1 11 1 11 2 10 0 9 0 1 11 2 10 12 9 0 1 15 4 13 10 9 10 9 1 10 9 7 10 9 0 13 1 10 9 11 1 10 9 1 10 9 0 2
55 10 9 1 10 9 1 10 9 0 2 0 7 1 9 9 0 13 0 7 0 10 9 0 1 10 9 1 9 2 3 10 9 1 9 1 10 9 1 10 9 4 4 13 2 1 2 1 9 2 1 10 0 0 11 2
13 10 0 9 4 3 4 13 7 13 10 9 0 2
26 1 10 9 1 15 10 9 1 9 4 13 9 1 10 0 9 1 10 9 13 13 1 10 0 9 2
37 9 9 2 13 1 15 13 15 1 10 9 9 11 1 10 0 9 7 10 0 9 13 1 10 9 1 13 10 9 7 13 10 9 7 10 9 2
29 9 9 2 16 15 13 13 1 15 13 15 1 16 2 1 10 9 1 10 9 2 4 13 10 9 1 10 9 2
35 13 3 0 16 3 1 10 9 1 15 1 10 9 1 10 11 11 4 13 9 3 0 2 10 9 1 9 3 15 13 1 10 10 9 2
41 4 13 1 10 10 9 15 13 1 10 9 1 10 9 11 2 15 4 13 10 9 1 9 1 9 1 10 9 7 10 9 0 2 7 15 3 3 15 13 3 2
51 10 9 13 13 16 10 9 0 3 13 3 16 13 10 0 9 1 10 9 1 9 1 10 9 0 0 2 0 1 9 1 12 9 7 9 2 7 10 9 1 9 0 0 1 10 9 1 10 9 9 2
77 1 10 10 9 4 13 10 9 1 13 9 1 10 9 0 2 10 9 1 9 7 10 9 0 2 1 9 16 10 10 9 13 2 1 10 9 0 7 3 0 2 1 10 9 0 1 10 9 1 9 7 1 10 9 1 9 1 9 10 15 2 1 0 2 13 10 12 9 0 1 10 9 1 15 4 13 2
19 4 13 10 9 0 1 10 9 7 4 13 10 9 13 1 9 1 9 2
21 10 9 4 3 3 13 16 10 9 3 4 4 13 1 9 1 9 1 10 9 2
47 1 10 9 13 13 3 0 13 15 1 10 9 1 10 9 7 1 10 9 15 4 13 1 13 10 9 0 1 10 9 2 13 16 10 9 15 15 13 13 13 15 1 13 10 9 0 2
35 7 13 1 4 15 13 2 9 9 2 16 10 9 12 2 9 12 1 10 9 1 11 13 10 9 15 13 1 10 9 0 1 10 9 2
32 1 9 13 13 16 13 1 13 1 10 9 1 9 1 10 9 12 2 12 15 3 4 13 10 9 1 9 1 10 0 9 2
41 1 10 9 15 13 10 9 13 1 10 9 15 13 1 13 9 13 1 10 9 1 9 1 13 10 9 1 9 0 7 10 9 1 10 9 1 9 1 9 0 2
47 13 16 1 10 0 9 3 1 3 2 1 9 1 10 9 1 10 9 7 1 15 1 10 9 1 11 2 10 11 13 9 1 9 0 7 0 1 10 9 7 10 9 1 10 10 9 2
21 10 9 13 9 1 13 10 9 2 13 10 15 2 7 1 13 1 10 10 9 2
28 9 7 9 1 9 0 13 10 9 1 13 15 7 1 13 10 9 2 1 10 9 1 9 2 9 7 9 2
19 10 9 13 9 1 13 1 9 1 9 1 10 0 9 1 10 10 9 2
42 10 9 15 13 13 9 1 10 9 0 7 0 15 13 1 15 0 7 1 10 10 9 10 9 0 1 10 9 0 7 13 2 16 0 2 1 0 9 1 9 0 2
19 1 10 9 4 13 10 9 1 9 7 10 9 4 13 10 9 0 0 2
44 1 13 15 1 10 9 0 2 11 4 13 10 9 1 9 9 15 15 13 1 10 9 1 10 9 7 1 10 9 0 2 13 3 9 0 0 1 13 10 9 1 10 9 2
18 3 4 13 10 9 13 1 10 9 15 15 13 3 16 3 13 9 2
15 16 3 13 10 9 2 3 4 13 10 9 1 10 9 2
6 13 3 10 11 11 2
41 2 13 3 0 1 9 0 1 4 4 13 1 10 0 9 1 9 1 10 9 0 1 10 15 1 10 9 1 10 10 9 7 16 10 9 13 1 10 10 9 2
30 10 10 9 1 11 4 13 1 11 11 2 10 10 9 1 10 12 1 10 0 9 1 10 9 1 9 0 1 11 2
19 13 1 13 15 0 10 9 2 13 9 3 1 10 9 3 0 1 11 2
15 1 10 9 2 13 10 9 1 9 7 13 1 10 9 2
7 10 10 9 3 4 13 2
28 10 10 9 1 9 13 13 13 10 9 0 1 10 12 7 1 10 12 1 10 9 7 3 13 1 1 9 2
30 1 11 13 2 3 10 9 7 10 9 2 2 4 3 13 1 13 1 9 1 10 9 15 13 9 1 10 10 9 2
32 10 9 1 15 13 1 10 9 2 7 11 13 1 10 9 16 11 13 2 1 10 9 1 0 9 2 7 2 13 3 2 2
11 10 9 13 10 0 9 0 16 15 13 2
22 11 13 1 13 10 10 9 1 9 0 2 7 3 0 7 3 0 2 7 3 0 2
33 16 13 1 10 9 1 1 15 2 11 13 1 9 10 9 2 13 1 9 0 7 13 9 1 15 15 4 13 1 10 9 0 2
21 2 10 9 1 10 11 11 2 2 15 13 2 2 13 0 2 13 1 10 9 2
16 2 11 13 0 9 1 9 3 15 1 11 11 7 11 11 2
40 3 15 13 1 9 16 11 13 1 13 2 7 9 0 7 10 9 1 10 9 13 16 15 1 10 10 9 4 13 1 9 1 10 9 0 3 1 10 12 2
20 11 4 13 1 10 9 1 10 9 1 10 0 9 12 9 1 10 10 9 2
40 10 9 13 1 10 9 1 9 15 13 10 9 13 10 9 1 15 13 13 10 10 9 2 15 15 4 3 13 1 10 9 1 9 1 10 9 1 10 12 2
23 11 13 1 0 12 9 3 3 13 2 11 0 7 0 12 0 9 2 3 1 11 11 2
23 1 11 2 11 13 3 10 10 9 0 2 1 9 1 10 9 3 0 1 10 0 9 2
25 1 10 0 9 1 11 2 15 4 3 13 1 10 9 3 0 2 15 9 10 9 1 10 9 2
21 1 10 9 1 10 0 7 0 9 2 10 10 9 15 4 13 3 1 10 9 2
42 3 10 0 9 1 9 13 16 15 13 9 1 13 1 9 10 9 0 1 10 9 2 7 10 9 2 1 9 10 9 0 1 10 9 0 2 13 1 10 0 9 2
6 9 0 2 15 0 2
32 10 9 13 3 0 9 3 0 7 0 0 0 15 13 10 9 1 10 9 0 2 13 1 10 0 9 10 9 1 9 0 2
24 10 9 2 1 15 0 2 3 13 10 9 16 3 15 13 15 1 13 15 7 1 13 15 2
5 11 12 2 12 2
12 3 1 10 9 2 10 11 4 13 10 9 2
30 7 2 1 10 9 10 2 10 11 15 4 13 1 10 9 1 13 10 10 9 13 2 13 3 3 0 1 10 9 2
20 1 10 9 2 3 2 10 9 15 4 13 10 9 1 9 15 16 1 9 2
43 13 13 1 10 9 1 9 7 13 15 1 9 7 9 0 2 10 11 13 1 13 1 1 10 9 1 10 9 7 1 10 9 1 9 2 7 1 10 9 1 10 9 2
23 16 10 9 0 13 3 2 10 9 1 10 9 13 3 0 1 15 3 13 10 9 0 2
14 10 10 9 13 9 2 3 1 10 0 7 0 9 2
13 7 3 10 9 13 3 0 1 15 13 10 9 2
50 13 3 0 16 10 0 9 1 10 12 9 1 10 9 2 13 9 1 10 9 0 7 0 1 10 10 9 2 3 13 1 9 1 10 9 1 15 10 9 1 10 9 13 10 9 1 10 10 9 2
18 15 13 10 9 0 1 10 9 0 1 13 9 0 1 10 9 0 2
49 1 11 1 10 9 2 11 7 3 2 13 7 13 10 9 1 10 9 13 9 1 10 9 0 7 1 10 9 1 10 9 2 3 1 10 9 0 2 3 1 10 9 1 10 9 1 10 9 2
21 10 15 13 10 9 1 9 15 4 2 7 3 13 2 4 13 1 10 10 9 2
30 1 10 9 1 10 9 0 2 4 13 1 0 13 9 1 3 13 10 9 1 13 0 9 1 9 0 1 10 9 2
15 15 1 9 4 3 13 2 7 1 3 3 1 9 10 2
26 10 9 0 7 0 0 1 10 9 4 13 3 2 3 15 13 3 3 13 1 10 0 1 10 9 2
8 4 4 13 10 9 1 9 2
30 1 9 2 10 9 4 13 1 13 10 11 3 0 2 3 1 13 10 9 1 10 11 1 10 9 1 13 10 9 2
13 10 0 9 13 16 10 9 3 15 4 3 13 2
50 7 2 16 10 0 13 1 13 10 10 9 1 10 9 0 1 11 11 2 13 10 0 9 2 3 2 9 1 2 9 1 9 2 2 10 0 9 1 10 9 0 13 1 13 10 9 1 10 9 2
29 16 3 15 13 10 9 1 10 9 1 9 0 1 11 2 3 15 13 10 9 1 13 10 9 0 1 10 9 2
21 3 2 16 15 13 1 9 0 2 10 9 13 13 10 9 0 1 1 10 9 2
15 10 11 13 10 9 2 7 3 13 1 9 1 13 15 2
19 3 2 13 10 0 9 0 13 10 0 9 0 7 10 0 9 1 9 2
