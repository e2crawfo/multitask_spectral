2527 17
2 0 9
9 13 3 13 11 0 9 9 9 2
20 3 9 9 9 2 3 9 13 13 9 9 15 2 13 15 4 13 7 13 2
7 3 9 13 3 3 0 2
11 9 13 0 12 0 9 7 12 9 1 2
19 15 13 13 15 13 2 13 9 2 13 0 9 13 9 2 13 9 9 2
25 9 13 3 3 3 0 2 16 0 9 13 0 9 7 9 2 0 9 4 3 13 9 7 9 2
7 0 9 2 16 13 9 2
5 7 16 13 13 2
8 9 11 11 9 13 0 0 2
12 9 13 7 0 9 13 13 13 16 15 13 2
20 16 9 3 13 9 13 9 7 3 13 0 3 0 9 2 4 9 13 9 2
7 9 13 13 2 13 9 2
17 9 4 13 9 2 16 9 13 9 2 15 2 2 9 13 15 2
10 16 9 13 9 2 9 4 13 13 2
4 8 2 8 2
4 7 2 7 2
5 9 13 0 9 2
6 3 9 13 3 9 2
15 11 11 3 13 9 1 7 13 15 3 0 7 0 9 2
10 13 3 0 13 9 7 9 15 9 2
14 9 3 11 11 13 0 9 7 15 4 3 13 3 2
12 15 13 13 9 7 9 9 13 9 9 15 2
8 3 9 13 15 3 3 9 2
19 13 4 16 13 2 13 9 7 3 9 0 9 3 13 9 9 0 9 2
6 15 13 3 4 13 2
2 9 13
12 0 9 4 13 9 9 1 3 0 9 9 2
16 13 9 2 9 2 1 2 7 15 13 3 3 13 3 0 2
12 3 13 7 9 13 9 13 9 0 7 0 2
22 9 4 13 3 0 9 2 15 13 3 3 0 16 3 2 15 15 9 2 5 2 2
12 9 13 15 9 15 9 9 7 13 9 2 5
12 3 4 13 15 9 7 3 3 4 15 13 2
18 13 4 13 2 13 15 9 3 13 9 9 2 7 15 0 7 0 2
14 3 3 13 2 16 9 13 13 9 7 9 1 2 5
12 0 0 13 15 2 16 9 4 13 3 2 5
21 9 13 13 3 2 7 3 0 9 7 0 9 9 7 9 7 0 9 3 9 2
13 9 1 13 2 16 9 4 13 9 9 12 9 2
12 4 13 2 16 9 13 15 9 0 0 9 5
22 13 3 3 15 9 2 16 0 9 9 1 13 0 9 0 16 0 9 7 0 9 2
8 13 3 15 9 3 0 9 2
3 0 2 5
4 9 2 9 2
13 3 13 9 13 2 15 3 2 15 9 3 13 2
13 13 4 3 13 15 9 2 16 13 0 9 2 2
4 13 3 9 2
12 13 15 9 2 3 9 4 13 3 3 9 2
10 15 13 15 9 1 2 9 2 9 2
16 3 13 13 3 15 13 9 2 7 15 9 4 13 0 9 2
38 11 9 9 13 3 0 2 16 16 9 13 9 2 3 9 2 9 9 1 7 9 15 3 15 9 2 2 3 9 3 13 13 9 9 7 13 3 2
14 2 13 15 3 4 13 15 0 9 2 2 15 13 2
11 15 11 13 2 16 2 15 13 13 2 2
23 3 4 13 3 3 2 9 0 9 2 2 16 13 16 11 9 9 9 13 3 13 9 2
11 13 3 15 15 9 2 15 13 13 2 2
19 4 13 2 16 11 13 3 13 9 2 9 2 15 2 15 15 9 13 2
23 13 15 2 15 13 13 15 9 2 16 11 13 9 2 7 11 13 13 7 15 0 9 2
12 15 13 3 13 3 9 2 7 3 3 9 2
6 15 13 15 9 3 2
6 15 15 13 15 9 2
7 7 15 13 3 15 9 2
26 7 16 3 13 15 9 2 3 13 3 2 16 15 13 15 9 7 15 9 2 16 3 15 13 9 2
27 9 13 9 13 9 9 15 7 9 3 9 2 13 3 9 9 2 9 9 7 3 9 7 9 9 9 2
15 15 13 0 9 2 16 15 4 3 15 13 9 13 9 2
10 9 13 15 2 15 13 13 9 3 2
24 15 13 13 3 3 15 13 2 3 13 7 3 3 13 2 7 15 15 13 0 9 7 9 2
12 9 13 3 9 9 9 7 15 9 15 9 2
17 3 15 13 2 16 9 4 13 3 15 9 7 13 15 9 9 2
17 6 2 3 15 13 3 2 16 9 13 3 0 2 16 15 9 2
8 3 15 13 3 13 3 0 5
19 9 13 15 9 3 15 9 7 9 2 0 7 9 2 3 13 13 9 2
18 9 13 3 15 9 2 9 2 9 2 9 2 0 9 9 9 3 2
15 3 13 0 13 15 9 13 2 16 9 13 3 15 15 2
15 9 13 9 9 0 9 13 2 3 15 13 15 9 2 2
19 15 13 0 9 2 9 2 15 13 15 13 2 3 13 7 13 3 9 2
20 15 2 13 9 0 16 9 2 13 3 0 13 2 13 15 15 15 9 13 2
6 15 4 3 13 9 2
22 9 4 13 3 0 9 2 7 9 13 3 0 2 3 0 2 3 2 0 2 9 2
5 3 9 13 9 2
16 15 13 15 9 15 13 13 2 3 9 2 15 13 3 15 2
13 9 9 9 13 3 3 0 2 3 9 9 13 2
21 9 13 13 3 9 7 13 15 9 7 3 9 2 15 13 2 13 2 13 3 2
11 9 9 13 9 2 16 15 13 13 13 2
21 3 15 13 3 0 9 2 16 15 13 13 13 2 16 0 2 9 2 13 9 2
6 15 3 9 15 9 2
10 15 13 15 2 16 13 13 15 9 2
24 16 9 9 15 9 13 0 9 2 15 13 0 13 7 3 13 2 3 13 15 4 9 13 2
10 13 9 3 13 2 16 3 13 9 2
18 7 15 13 15 2 16 0 16 13 15 2 15 13 15 7 13 0 2
18 9 13 9 2 9 7 9 4 13 13 3 0 3 2 16 0 9 2
20 15 13 3 15 9 13 9 2 15 3 15 9 13 3 0 2 16 0 9 2
10 3 9 4 13 3 15 9 3 3 2
10 13 15 9 2 15 15 9 13 15 2
12 15 15 15 13 16 9 7 9 9 9 9 2
20 9 2 9 7 9 13 9 7 9 2 9 13 9 7 0 9 9 3 13 2
13 13 15 9 1 9 9 9 3 9 7 9 1 2
15 13 15 2 16 3 13 3 9 1 2 9 2 3 3 2
16 15 9 13 15 9 2 16 15 13 9 2 16 13 3 9 2
18 3 15 13 15 2 15 9 13 13 9 2 16 9 13 3 2 3 2
23 0 9 13 9 2 15 13 16 13 15 2 2 7 16 9 15 13 2 3 9 13 9 2
8 13 15 15 9 9 15 9 2
12 13 16 15 13 0 2 13 15 13 7 13 2
3 13 15 2
6 16 3 13 15 9 2
8 9 2 9 2 13 15 9 2
14 13 9 0 9 1 9 2 7 0 9 1 9 9 2
11 13 9 9 13 9 7 9 15 13 9 2
19 3 13 3 13 13 9 0 7 0 2 7 15 9 13 15 9 13 9 2
16 16 3 13 15 9 13 2 3 15 13 0 9 9 9 1 2
20 15 13 3 9 7 0 9 2 15 13 9 13 15 9 2 15 15 3 13 2
21 15 13 0 9 2 3 9 2 0 9 2 3 9 2 0 9 9 2 0 9 2
7 9 13 9 3 9 9 2
27 15 15 9 13 9 2 3 16 13 9 15 9 2 9 2 9 2 9 2 9 2 15 15 13 3 9 2
6 3 13 9 13 9 2
36 3 13 15 13 2 16 9 2 9 7 0 9 13 15 0 2 16 15 13 15 13 2 15 1 2 16 15 13 15 13 13 9 9 13 9 2
28 9 4 13 13 9 2 3 16 15 13 15 2 13 15 2 2 16 15 13 13 16 2 13 9 3 3 2 2
9 9 11 2 9 13 3 0 9 2
19 3 9 13 15 15 0 9 2 7 3 13 9 2 15 4 13 0 9 2
20 4 3 13 9 9 9 7 13 15 13 15 2 15 1 4 13 9 3 9 2
8 15 9 1 9 13 0 9 2
12 9 1 11 9 9 9 13 13 13 9 9 2
6 15 13 13 9 9 2
7 9 13 3 13 15 9 2
13 4 13 9 2 7 4 13 9 15 0 9 9 2
21 0 9 2 13 13 12 9 3 9 9 1 2 15 13 13 9 9 9 7 9 2
16 13 3 13 12 9 15 15 9 9 2 15 13 0 9 1 2
17 3 13 2 16 15 13 12 9 9 11 2 15 13 9 0 9 2
41 0 13 2 16 15 13 2 16 9 9 13 13 0 9 9 2 3 3 16 13 11 9 9 2 15 3 13 3 9 9 2 15 13 3 3 9 9 2 3 11 2
36 0 15 9 2 3 3 9 2 9 13 4 13 3 3 2 15 13 3 0 2 7 15 1 13 0 13 2 16 13 9 4 13 9 15 9 2
14 0 13 13 9 11 11 0 9 2 15 15 4 13 2
22 2 2 0 9 2 0 9 9 2 0 9 2 13 15 9 13 9 0 9 9 9 2
22 13 9 13 2 16 0 9 9 4 9 9 3 7 13 13 15 9 9 9 11 9 2
23 12 0 9 9 2 15 4 13 0 9 7 13 9 0 9 2 4 13 3 15 0 9 2
23 11 9 9 13 15 3 0 2 16 9 12 9 13 0 2 0 7 0 9 11 0 9 2
23 9 13 9 4 13 15 9 13 9 2 3 11 9 2 13 3 3 3 0 9 9 9 2
22 9 0 9 13 13 0 2 7 13 2 16 15 2 0 9 9 2 13 3 15 9 2
39 11 0 0 9 0 0 2 0 7 0 9 13 0 9 15 9 2 7 13 13 3 2 15 4 13 0 9 2 15 13 0 15 2 15 13 13 13 15 2
17 3 13 15 0 9 0 9 9 2 15 11 7 11 13 11 9 2
16 13 0 2 16 15 9 13 9 4 13 15 9 15 15 9 2
10 3 13 0 9 9 13 9 13 9 2
7 3 13 9 13 11 9 2
5 15 13 11 9 2
3 15 11 2
18 12 9 13 9 2 11 0 9 0 0 9 2 15 13 15 0 9 2
16 9 4 13 0 9 2 15 13 15 0 9 9 9 12 9 2
11 15 1 13 0 13 15 15 9 0 9 2
17 3 0 9 13 11 9 9 9 0 9 2 15 15 9 4 13 2
14 13 15 0 9 7 9 2 15 13 3 0 9 9 2
75 9 13 0 2 9 15 9 9 9 2 15 13 3 0 9 7 0 0 9 0 9 0 9 2 0 9 9 11 7 11 9 2 9 9 0 9 2 0 7 0 9 9 7 15 9 9 2 0 9 15 9 9 2 0 9 9 9 2 15 13 3 3 9 9 7 9 2 0 9 7 0 9 9 9 2
10 15 9 13 0 9 13 12 9 9 2
16 3 13 9 2 15 13 3 9 9 3 13 0 9 7 9 2
21 0 9 9 13 0 0 9 2 16 4 13 9 9 7 13 3 15 9 13 9 2
12 3 13 9 2 15 13 9 9 9 0 9 2
26 0 9 13 0 9 9 13 0 9 9 7 3 15 2 3 0 9 13 0 9 2 15 9 3 13 2
17 13 0 9 2 16 0 9 9 0 9 13 9 13 0 0 9 2
21 0 9 2 11 9 13 9 13 0 3 2 16 15 13 3 13 11 9 9 1 2
19 16 9 13 13 0 13 2 9 13 15 0 0 2 13 13 3 0 9 2
9 0 7 0 9 1 13 9 9 2
38 15 9 13 0 2 16 7 3 11 4 13 0 9 2 3 3 4 3 13 15 2 16 15 9 9 4 13 9 7 9 9 3 0 9 16 11 9 2
15 3 4 13 13 0 0 9 2 7 0 9 4 13 9 2
11 4 13 2 3 9 1 9 13 9 13 2
15 4 13 2 3 0 7 3 0 9 9 9 9 4 13 2
18 4 13 2 3 9 13 9 9 2 7 3 0 9 9 13 9 13 2
24 11 9 2 8 2 13 9 9 9 2 8 2 1 2 7 11 9 13 9 13 9 0 9 2
19 9 13 3 3 3 2 13 15 13 3 15 9 9 2 16 15 9 13 2
13 9 11 9 13 13 3 0 0 9 15 15 9 2
12 9 13 9 9 2 15 9 13 3 9 9 2
38 15 9 7 15 13 9 2 4 13 3 13 3 15 9 2 15 13 3 9 13 9 9 2 9 9 4 13 9 9 2 15 9 13 13 0 9 11 2
3 11 2 11
9 9 9 13 3 7 13 1 9 2
26 13 13 3 15 4 13 2 13 4 3 13 13 9 13 13 15 15 9 2 15 0 9 11 9 13 2
15 3 13 9 2 9 3 3 2 15 9 7 9 3 3 2
79 9 9 13 9 2 6 3 0 3 13 2 13 13 9 7 9 15 3 13 2 3 9 9 7 0 9 2 0 9 9 2 15 9 15 13 2 13 9 2 9 13 9 2 13 3 13 2 0 9 16 13 2 15 9 13 2 0 16 15 13 9 2 13 13 2 13 13 15 9 16 15 9 13 13 9 2 0 9 2
52 0 13 9 15 9 2 15 13 9 9 2 13 9 16 15 13 8 8 2 13 3 9 15 9 7 13 13 2 9 13 0 7 15 13 9 7 9 3 9 9 1 16 13 3 15 13 2 9 13 3 9 2
18 9 9 13 16 9 2 9 13 9 11 2 0 11 2 15 13 3 2
34 3 3 9 9 13 9 2 9 13 9 2 9 13 13 9 9 9 2 16 13 9 13 13 3 9 13 2 9 13 3 3 0 9 2
10 13 3 3 9 2 16 9 13 3 2
15 13 15 13 9 2 15 13 9 7 13 9 2 13 0 2
24 3 13 2 16 9 9 13 0 9 15 0 9 2 15 13 7 13 9 2 7 13 3 9 2
36 0 9 9 13 9 1 2 13 3 9 2 13 3 9 9 1 2 13 13 9 2 13 3 2 13 9 2 15 9 2 3 2 3 2 3 2
6 0 9 13 9 9 2
17 13 15 9 1 2 15 13 3 9 2 13 16 15 13 15 3 2
1 9
14 9 13 3 3 9 2 16 13 0 9 9 13 9 2
7 4 13 9 13 9 1 2
19 9 13 15 3 3 7 3 3 2 16 3 13 15 1 7 13 13 9 2
9 13 9 3 2 16 9 13 9 2
10 13 9 7 13 0 0 9 1 9 2
12 9 4 13 9 0 9 3 7 13 15 9 2
25 15 13 13 3 3 0 9 2 3 13 15 1 2 7 3 1 2 16 13 13 13 9 15 1 2
15 15 13 15 3 13 2 13 9 9 7 13 15 3 3 2
11 15 3 13 3 3 7 13 15 9 3 2
7 13 7 13 13 9 3 2
11 9 13 0 3 7 15 13 0 0 9 2
6 2 9 2 15 13 2
3 2 9 2
5 0 7 0 9 2
3 3 13 2
3 2 6 2
4 2 13 13 2
10 13 13 2 9 13 7 13 13 9 2
10 2 4 15 9 13 2 13 13 3 2
18 2 13 0 2 9 13 7 13 9 9 13 9 2 15 13 3 9 2
17 13 13 9 7 13 9 2 15 13 13 0 9 9 7 3 9 2
16 15 4 3 13 15 9 13 9 7 0 9 15 9 7 9 2
8 9 13 4 4 3 13 9 2
13 2 3 3 2 9 13 7 13 3 9 13 9 2
4 13 9 9 2
13 9 13 3 0 9 7 9 0 9 13 15 1 2
14 9 13 9 2 13 3 13 15 2 7 13 9 9 2
4 15 13 0 2
20 15 13 3 0 16 15 3 13 2 7 15 13 15 9 3 3 16 13 13 2
5 7 3 15 13 2
13 9 13 3 0 7 13 3 3 2 3 3 13 2
8 3 3 13 9 9 13 0 2
15 4 13 15 9 2 7 13 3 0 7 13 9 3 3 2
12 13 13 15 15 9 2 15 13 13 13 3 2
16 16 9 13 9 2 9 3 13 3 0 7 0 7 13 3 2
12 16 15 3 13 9 9 2 15 13 15 9 2
8 2 3 13 9 7 0 9 2
4 4 13 15 2
18 13 13 3 2 7 0 9 13 3 13 9 9 7 13 15 3 13 2
23 13 13 9 9 2 13 13 15 13 9 2 7 15 13 0 2 0 9 7 13 15 9 2
18 2 9 13 2 15 13 7 13 3 9 3 3 16 15 13 3 9 2
2 11 9
12 11 0 9 11 13 13 15 9 16 0 9 2
20 16 11 13 9 13 2 11 13 13 9 15 2 15 13 11 0 7 0 9 2
16 11 13 15 0 9 9 2 16 9 13 13 11 0 9 1 2
13 11 13 3 13 15 13 9 0 7 3 0 9 2
8 9 11 9 13 3 9 1 2
12 15 9 13 9 9 11 2 15 4 13 11 2
12 15 13 13 9 3 3 0 7 13 15 9 2
15 9 15 2 16 11 13 3 15 13 9 13 11 0 9 2
21 2 15 4 13 3 3 9 2 16 13 13 11 3 0 9 2 11 13 9 11 2
6 2 3 13 15 9 2
8 2 15 13 9 9 1 9 2
3 11 13 2
16 2 16 13 15 9 11 2 13 3 13 13 15 3 0 9 2
11 13 15 0 9 2 15 13 13 15 0 2
13 11 13 11 2 7 13 3 15 13 3 7 13 2
9 11 13 9 7 13 15 3 9 2
17 3 9 13 0 9 11 9 7 9 0 9 13 15 9 11 1 2
9 11 13 7 15 13 9 0 9 2
6 15 9 4 13 9 2
17 11 13 13 9 13 3 9 7 3 9 2 15 15 13 13 0 2
16 11 9 13 15 9 3 0 9 2 3 15 13 3 0 9 2
16 11 7 11 13 13 3 2 3 0 9 2 15 3 13 9 2
10 11 7 11 13 0 7 0 9 1 2
12 9 9 1 13 0 2 13 3 13 0 9 2
10 15 9 1 15 13 9 9 0 9 2
17 15 13 0 9 9 2 3 3 16 3 0 9 13 13 3 9 2
14 11 7 11 13 3 2 15 13 9 13 9 13 3 2
18 15 3 16 11 4 13 9 7 13 9 2 15 13 13 9 9 1 2
5 9 9 13 9 2
18 15 13 4 13 9 9 13 2 16 9 13 0 7 15 9 13 0 2
8 13 3 9 11 13 13 11 2
14 11 13 3 13 11 2 7 13 3 9 9 13 9 2
15 9 13 3 3 2 16 3 9 13 0 0 3 0 9 2
14 9 13 3 3 2 3 15 13 13 9 13 7 13 2
19 16 15 13 9 2 15 1 13 0 9 2 15 15 13 3 13 0 9 2
9 9 13 13 3 9 13 13 3 2
9 11 13 2 13 9 15 13 9 2
11 2 15 13 11 2 11 9 2 9 13 2
10 2 15 13 3 3 16 11 13 0 2
11 16 9 13 2 15 13 13 9 13 9 2
19 2 3 15 4 13 15 11 2 16 15 13 15 16 13 9 2 11 13 2
14 2 3 16 13 2 15 15 13 2 9 13 3 3 2
10 15 13 3 13 9 13 3 15 0 2
10 2 11 13 13 13 9 2 9 13 2
6 2 13 15 13 9 2
12 9 2 9 7 15 9 13 9 13 9 9 2
7 11 13 9 7 9 3 2
12 9 13 9 7 13 9 2 13 9 15 9 2
13 13 13 2 3 11 7 11 13 13 9 15 9 2
10 11 13 0 9 7 9 9 0 9 2
10 2 4 13 0 9 2 11 13 9 2
23 2 9 9 11 4 13 0 9 2 7 3 4 13 15 0 2 15 13 13 11 0 9 2
15 2 9 13 3 3 2 16 3 9 13 0 2 11 13 2
12 2 16 13 13 11 2 13 13 16 13 9 2
8 11 13 2 13 11 13 9 2
12 0 9 15 13 13 9 15 9 16 11 13 2
11 15 13 9 0 9 9 7 11 13 9 2
12 11 13 13 3 9 2 7 11 13 13 9 2
6 3 11 13 15 1 2
20 11 13 1 0 13 0 9 2 7 15 9 13 13 3 16 15 13 9 1 2
6 11 13 9 13 9 2
15 9 4 13 3 7 11 4 13 0 9 13 13 9 1 2
7 13 9 11 13 13 11 2
8 11 4 3 13 13 0 9 2
12 11 13 9 2 15 4 13 0 9 1 9 2
19 11 4 13 12 9 9 9 2 16 15 13 4 13 9 11 9 9 1 2
22 11 13 13 9 11 7 13 2 16 15 13 11 9 16 15 13 11 9 1 11 9 2
12 9 13 0 7 15 9 13 9 9 9 1 2
7 9 13 7 9 9 13 2
15 11 13 9 3 1 11 7 11 13 13 9 13 0 9 2
8 13 9 11 13 15 0 9 2
15 3 13 9 2 3 11 4 13 15 9 15 13 9 9 2
17 15 9 11 13 11 9 7 9 11 13 2 16 9 13 11 9 2
15 3 13 3 11 0 9 2 3 9 13 13 11 0 9 2
2 0 11
8 11 13 9 9 7 13 15 2
7 15 4 3 3 13 3 2
6 9 9 4 13 0 2
7 0 9 9 13 9 13 2
5 15 13 0 15 2
5 15 13 3 9 2
4 13 13 9 2
4 9 13 9 2
7 9 9 11 9 13 13 2
8 9 9 13 9 7 13 3 9
7 3 9 13 3 3 13 2
6 15 15 4 13 3 2
7 15 13 13 16 15 13 15
9 13 9 0 9 2 16 3 13 2
3 9 13 12
3 6 15 15
5 13 9 12 9 2
5 9 13 9 1 2
4 9 13 9 2
7 11 13 0 9 9 3 2
7 11 9 7 9 13 15 2
17 7 16 15 13 13 13 9 3 3 2 15 13 0 0 9 9 2
6 15 13 7 9 13 2
15 9 13 9 9 7 3 13 3 9 2 11 13 0 9 2
7 16 15 4 13 9 9 2
14 15 13 13 0 9 13 2 16 13 3 13 15 9 2
8 2 13 11 7 13 9 2 2
17 15 9 7 15 9 4 13 15 9 2 16 4 13 13 15 3 2
12 11 13 9 2 15 13 13 9 3 13 9 2
8 9 0 9 13 13 3 0 2
24 15 13 13 3 3 16 16 13 15 9 7 6 3 16 3 13 15 2 6 15 3 3 9 2
9 3 13 15 15 0 9 7 9 2
16 9 13 13 15 0 9 2 3 0 9 4 13 3 9 3 2
4 15 11 13 2
11 9 13 13 9 9 7 9 13 0 9 2
2 13 13
12 15 13 9 0 0 11 13 15 9 9 9 2
7 9 13 3 3 9 1 2
10 7 13 9 11 2 15 9 13 3 2
13 15 4 13 15 9 2 15 0 9 13 0 9 2
4 9 13 9 9
12 11 9 13 9 13 13 9 2 7 13 9 2
10 9 13 9 2 16 9 13 15 9 2
12 16 0 13 2 15 4 3 15 1 13 13 2
14 13 3 13 11 9 9 11 9 9 2 16 9 13 2
7 15 13 13 15 13 9 2
3 9 13 2
10 9 9 13 7 13 12 9 9 13 2
7 13 3 2 16 13 15 2
42 9 9 2 13 12 9 9 12 2 9 9 12 7 12 9 9 7 9 7 9 7 9 9 13 9 9 9 13 9 12 7 12 9 2 13 9 12 12 2 2 12 2
91 11 9 9 2 15 13 9 11 9 9 2 13 9 9 13 9 9 12 9 9 12 13 9 9 12 2 12 2 2 0 16 15 13 3 13 9 12 2 12 2 2 7 3 15 12 9 12 7 12 9 2 13 9 9 13 9 9 12 9 9 12 13 9 9 12 2 12 2 2 0 16 15 13 3 13 9 12 2 7 3 15 12 9 12 7 12 9 2 7 13 2
60 16 12 2 9 12 9 12 13 9 9 12 2 12 2 7 12 2 12 2 2 0 16 15 13 13 12 9 9 12 13 9 9 12 2 12 2 2 7 12 9 9 12 13 9 9 12 2 12 2 2 13 9 12 7 12 9 13 0 9 2
25 12 2 9 4 2 15 9 2 13 9 9 7 9 7 9 13 9 13 9 9 0 9 0 9 2
27 12 2 15 9 2 15 9 13 0 16 12 12 9 2 4 13 9 13 3 15 9 7 9 13 9 9 2
14 12 2 11 7 11 4 13 3 13 9 13 9 2 7
17 12 2 15 9 13 9 9 12 2 12 2 13 0 9 9 0 2
5 4 13 15 9 2
2 12 9
5 13 9 12 3 2
16 13 9 0 13 9 9 9 2 9 2 1 9 2 11 2 2
2 12 9
5 13 9 12 3 2
28 9 0 13 9 9 13 9 2 9 2 1 13 9 2 11 2 2 13 9 2 9 2 1 9 2 11 2 2
2 12 9
7 15 9 4 13 15 9 2
7 13 11 12 9 9 12 2
7 9 1 11 11 11 9 9
30 9 9 2 13 12 9 9 12 2 9 12 7 12 9 11 9 9 13 9 9 1 2 11 9 0 9 2 2 12 2
98 11 9 9 2 15 13 9 11 9 9 2 13 9 9 9 13 9 0 9 9 7 0 9 13 9 9 12 9 9 12 13 9 9 12 2 12 2 2 0 16 15 13 3 13 11 2 11 7 11 9 2 7 3 15 12 9 12 9 2 12 9 9 9 7 12 9 2 7 13 2 16 9 9 12 2 12 2 2 0 16 15 13 13 9 12 2 12 2 2 13 0 0 9 9 9 9 1 2
27 13 9 9 11 9 4 13 15 13 9 9 2 15 4 3 13 11 9 2 7 13 9 0 9 13 9 2
18 9 9 11 13 9 9 9 9 9 13 13 3 9 3 13 9 9 2
31 11 4 13 3 12 9 9 0 9 2 9 7 11 11 9 2 7 11 9 13 4 13 3 3 2 13 15 9 1 13 2
37 0 9 13 4 13 11 3 12 9 2 7 9 15 9 1 2 15 13 11 2 11 7 11 0 9 9 9 9 12 1 2 13 4 13 3 9 2
35 11 9 4 13 13 9 7 9 9 2 9 7 9 12 9 13 15 9 12 9 9 13 0 9 9 7 9 9 7 15 9 13 9 9 2
20 11 9 4 13 0 9 9 13 9 13 9 9 2 7 0 9 13 3 13 2
13 3 9 12 12 9 7 12 9 12 9 9 13 2
22 9 9 7 9 13 9 4 13 13 9 0 9 9 2 15 9 15 13 3 13 9 2
23 9 9 12 7 12 2 12 2 4 13 3 2 7 15 9 13 9 13 13 9 9 0 2
5 4 13 15 9 2
2 12 9
70 13 9 12 9 9 2 11 2 12 2 11 9 2 3 2 2 11 11 2 11 2 11 11 11 2 11 2 11 2 11 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 3 13 11 9 2 2 11 2 11 2 11 2 11 2 11 7 11 11 9 2
2 12 9
5 13 9 12 3 2
23 0 13 9 2 11 2 12 2 2 12 2 2 9 9 0 13 9 9 13 0 9 9 2
30 0 13 9 2 11 2 9 9 0 13 9 9 9 7 13 15 3 15 0 9 9 2 15 13 9 9 9 4 13 2
2 12 9
7 15 9 4 13 15 9 2
7 13 11 12 9 9 12 2
6 9 1 11 11 9 9
1 9
2 15 9
3 9 2 2
23 0 9 9 1 13 9 13 3 15 9 1 9 13 9 2 3 3 13 0 13 9 9 2
12 0 9 9 9 13 13 9 3 12 9 9 2
10 15 9 11 13 3 3 15 9 9 2
13 15 15 9 1 3 0 9 13 9 13 9 13 2
11 0 9 9 4 3 13 3 15 9 1 2
13 13 13 3 2 9 2 9 9 7 13 3 9 2
13 9 13 9 13 2 16 4 9 13 13 0 3 2
9 11 4 15 9 13 9 3 3 2
11 0 9 4 3 13 3 7 9 13 0 2
6 4 13 13 9 0 2
6 15 9 4 9 13 2
11 0 9 13 3 2 3 16 3 3 3 2
9 4 13 3 0 13 0 9 13 2
5 13 3 3 13 2
11 4 3 13 13 0 9 7 3 0 9 2
5 11 2 9 0 9
9 9 11 13 9 0 9 0 9 2
12 9 1 9 9 13 13 3 13 0 9 9 2
14 9 9 13 12 12 9 2 15 13 9 12 9 0 2
9 9 13 3 0 0 9 3 9 2
12 9 1 9 13 12 9 7 13 12 12 9 2
10 9 9 9 13 3 12 9 12 9 2
14 9 1 9 9 3 13 13 12 12 9 12 12 9 2
10 0 9 1 9 13 12 9 12 9 2
10 2 9 1 11 0 9 9 13 3 2
14 13 13 0 9 9 3 13 9 7 8 13 0 9 2
16 13 3 3 13 13 9 9 0 9 2 9 11 11 13 9 2
8 11 4 13 0 9 9 3 2
9 9 13 9 1 9 13 0 9 2
13 9 9 9 13 9 9 1 15 9 16 9 9 2
11 11 1 15 9 9 9 9 13 3 0 2
5 11 13 3 3 9
17 12 9 1 13 0 9 3 11 9 9 9 2 13 9 11 11 2
26 13 11 0 9 11 12 9 1 9 9 13 2 16 9 4 13 3 0 0 9 9 2 15 13 9 2
16 11 1 15 13 2 16 9 13 0 3 0 7 0 9 1 2
6 3 0 9 13 11 2
7 15 1 13 11 7 11 2
12 0 13 11 13 0 12 12 9 3 16 13 2
11 3 0 9 13 11 2 3 11 7 11 2
21 9 1 9 13 9 2 15 9 7 9 4 13 9 15 3 2 16 15 13 0 2
15 11 9 9 11 11 9 11 9 13 0 9 1 9 9 2
17 11 13 2 16 11 2 11 7 11 4 13 9 3 12 9 9 2
22 15 9 3 11 2 11 7 11 13 3 0 9 9 2 16 4 13 0 9 13 9 2
17 2 0 9 9 7 0 9 9 13 0 9 9 2 11 13 11 2
18 3 9 13 0 0 9 7 9 3 2 16 13 13 9 9 13 9 2
15 11 1 15 13 2 4 9 13 0 9 13 0 9 9 2
21 9 4 13 12 9 2 13 9 9 7 13 9 2 15 9 13 3 0 9 0 2
7 11 2 9 9 13 13 11
23 11 9 13 9 2 15 1 11 11 2 9 9 12 2 13 13 11 15 9 2 9 13 2
11 11 0 9 1 11 4 13 11 9 9 2
18 9 9 4 3 13 0 2 7 15 9 4 13 9 3 2 11 13 2
6 11 9 13 9 1 2
9 9 0 9 13 12 9 9 9 2
16 11 13 15 15 9 9 0 9 2 16 15 9 13 3 0 2
15 3 9 9 13 9 2 15 13 9 0 0 11 9 3 2
7 9 13 9 9 11 0 2
11 11 7 11 9 4 13 13 15 9 3 2
9 11 11 9 4 15 9 3 13 2
15 11 11 13 0 0 12 12 9 7 11 3 12 12 9 2
10 11 1 11 11 13 9 11 0 9 2
3 11 0 9
11 9 11 7 9 11 13 0 9 0 9 2
12 0 9 1 11 4 13 0 9 3 9 9 2
9 9 13 3 11 7 11 13 9 2
13 11 13 9 13 11 9 13 11 9 7 15 9 2
7 11 9 9 13 11 11 2
13 9 1 11 7 11 13 13 15 2 0 2 9 2
7 9 13 11 11 0 9 2
17 3 9 13 15 2 16 9 13 9 9 13 11 7 11 0 9 2
4 9 9 9 11
17 9 11 11 13 9 9 13 9 7 9 9 9 2 0 9 0 2
9 9 11 11 13 9 9 9 12 2
31 2 13 0 2 16 9 13 3 15 9 7 9 9 2 15 13 15 2 16 9 7 9 13 9 3 7 3 2 11 13 2
26 9 13 2 16 0 9 11 9 9 9 11 11 4 13 13 9 7 9 9 9 2 9 7 9 9 2
13 11 13 3 9 9 9 7 9 1 9 0 9 2
18 11 4 9 1 15 4 13 9 7 13 3 9 2 9 7 0 9 2
18 9 9 9 2 0 9 0 11 13 7 13 15 7 15 9 9 9 2
14 9 13 9 12 9 9 12 9 7 9 9 13 9 2
6 9 13 9 11 11 2
7 9 13 9 12 12 9 2
5 11 9 9 13 9
12 9 13 0 0 9 2 0 9 9 7 9 2
25 11 9 13 9 3 11 9 7 11 11 11 1 9 12 9 2 15 13 9 7 9 7 9 9 2
12 9 13 15 9 2 9 2 9 7 9 2 2
9 11 9 9 11 11 13 9 9 2
8 11 13 9 13 0 11 9 2
24 15 13 9 9 0 9 7 9 13 13 2 13 11 9 9 9 2 15 13 11 0 0 9 2
23 2 3 11 9 4 13 9 7 13 9 2 16 15 13 3 13 9 9 15 9 0 9 2
14 3 11 1 4 13 0 9 2 15 13 13 0 9 2
10 2 0 9 13 13 0 9 0 9 2
16 11 13 2 16 9 13 3 9 2 0 0 9 9 7 9 2
15 9 13 3 13 11 9 0 9 0 9 2 9 7 9 2
15 9 13 9 9 9 2 9 7 9 13 9 3 9 1 2
14 2 9 13 2 16 9 9 7 3 0 9 9 13 2
8 11 13 9 12 9 3 0 2
15 2 0 9 13 3 2 16 9 13 15 7 13 15 1 2
24 9 11 11 11 9 9 13 13 9 2 0 9 11 9 9 3 13 9 9 7 9 13 9 2
22 11 13 13 11 9 11 2 15 9 13 15 2 16 9 4 3 13 13 9 0 9 2
19 11 13 2 16 15 9 9 4 13 15 2 16 13 9 9 7 9 1 2
18 2 9 13 9 2 15 13 0 9 9 7 15 4 13 3 7 3 2
14 11 9 9 4 13 13 9 9 3 2 15 9 13 2
24 3 13 9 9 13 13 9 11 2 15 9 15 4 13 0 9 13 9 2 0 9 7 9 2
18 2 11 13 3 3 9 2 15 9 13 13 9 9 0 2 11 13 2
5 4 0 9 13 2
18 11 0 9 0 9 7 15 9 9 7 9 13 9 13 11 9 12 2
42 11 9 9 9 9 9 7 9 13 9 9 13 13 2 0 9 0 0 9 0 9 13 3 7 9 9 1 2 3 9 9 13 9 9 7 3 9 9 13 9 13 2
20 0 9 9 13 9 2 9 9 7 9 9 13 0 3 0 9 0 9 9 2
16 15 3 13 2 16 9 9 7 9 13 13 3 1 15 9 2
8 9 9 13 13 13 9 9 2
23 3 13 2 16 16 9 13 2 15 13 13 3 9 9 7 9 13 13 9 3 0 9 2
9 9 1 9 13 3 15 3 9 2
16 9 7 9 9 0 9 13 3 0 13 15 0 9 7 9 2
23 9 9 1 9 13 13 0 9 9 2 7 9 9 13 13 3 9 7 2 9 2 9 2
22 9 9 9 13 2 13 0 9 0 9 1 13 3 9 2 16 9 13 9 7 9 2
9 9 13 3 9 9 7 9 9 2
7 9 9 9 13 3 13 2
11 9 13 11 13 12 0 9 0 9 9 2
16 7 9 7 9 9 1 9 9 13 3 3 7 9 13 0 2
14 15 1 9 9 0 13 9 0 7 13 0 9 9 2
10 9 13 9 13 3 0 0 9 9 2
20 9 3 9 13 3 3 15 2 16 0 9 0 9 9 13 3 3 3 3 2
13 9 13 1 9 0 9 2 15 4 13 9 9 2
20 9 13 9 9 13 9 7 9 2 9 9 2 9 7 0 9 7 9 9 2
5 3 13 9 9 2
21 9 13 11 9 9 9 9 9 7 9 9 9 9 7 11 9 9 11 9 1 2
10 9 13 9 11 11 11 9 9 9 2
22 11 11 2 3 12 2 11 2 0 9 12 2 11 2 13 9 7 11 9 9 9 2
15 11 13 3 9 9 11 11 9 7 13 9 9 12 1 2
19 13 9 9 12 15 13 9 11 11 9 12 7 11 9 9 9 9 12 2
14 9 12 11 13 11 9 7 15 13 15 9 9 1 2
36 11 13 9 2 9 7 9 9 2 9 7 9 11 11 9 7 15 13 3 0 9 13 9 9 2 15 13 0 9 13 9 11 9 9 12 2
9 11 13 0 11 13 0 9 9 2
15 15 4 13 9 9 2 3 15 13 13 0 2 0 9 2
5 11 13 0 9 2
15 0 9 13 12 11 11 9 0 9 11 8 11 11 9 2
16 11 9 13 3 3 12 2 16 11 11 13 9 11 0 9 2
17 11 13 3 9 3 7 13 9 9 3 3 13 11 9 9 12 2
10 0 0 11 9 13 11 3 15 9 2
27 0 9 13 9 3 8 8 8 2 0 9 9 2 8 8 2 8 9 9 2 8 2 13 8 0 9 2
13 9 12 2 15 13 12 2 13 3 0 11 9 2
8 9 12 13 9 12 9 9 2
17 0 9 1 5 2 5 7 5 13 15 0 9 0 9 7 9 2
12 5 13 9 12 7 13 0 0 9 13 9 2
9 11 13 3 12 13 9 12 1 2
35 0 9 13 3 13 9 7 15 13 0 0 9 2 3 9 9 2 11 2 8 9 2 11 9 13 9 2 0 8 9 7 0 0 9 2
6 9 13 3 11 9 2
7 0 11 9 9 13 12 2
13 9 12 2 15 13 12 2 13 0 5 9 9 2
17 11 4 13 0 9 12 2 15 13 0 9 7 11 13 0 9 2
22 9 12 13 9 12 9 11 11 2 7 3 13 9 3 9 8 8 8 7 8 9 2
21 0 0 9 5 13 12 2 7 15 13 3 0 9 9 2 8 2 8 8 2 2
12 9 12 13 9 12 7 15 13 9 15 9 2
13 12 0 9 13 3 9 0 9 9 12 0 9 2
20 9 12 13 12 9 9 2 3 9 3 13 9 9 7 9 9 7 9 9 2
9 3 0 9 11 9 9 9 13 2
11 11 11 11 11 13 0 11 11 9 9 2
5 15 13 9 12 2
20 9 13 9 2 15 9 13 9 2 0 9 13 9 7 13 9 13 9 15 2
7 3 9 13 9 13 9 2
15 9 13 0 9 9 2 15 13 3 0 9 0 9 11 2
10 9 9 4 3 13 3 12 12 9 2
18 0 0 9 9 13 0 9 9 12 1 9 9 2 13 11 9 11 2
9 0 9 9 13 3 12 9 3 2
10 9 12 9 13 9 11 13 12 9 2
21 11 9 13 0 9 3 9 9 2 12 9 3 9 13 13 11 12 7 11 12 2
16 11 9 13 3 9 11 9 2 15 9 13 0 11 9 9 2
11 9 12 1 11 13 3 3 3 12 9 2
18 9 9 13 9 7 9 9 9 9 3 9 9 7 15 9 9 13 2
21 3 11 9 13 3 9 12 9 9 7 9 13 9 7 0 0 9 13 9 12 2
24 16 0 9 1 9 4 13 2 0 9 2 7 3 13 2 9 4 3 3 13 9 0 9 2
20 9 13 9 7 9 13 9 15 1 2 16 9 13 3 7 13 3 15 9 2
16 9 7 9 9 9 13 13 0 9 9 7 13 3 9 9 2
9 9 9 4 3 13 3 9 9 2
17 3 0 13 9 7 9 4 13 9 7 15 9 9 13 3 0 2
18 3 3 13 9 9 2 9 7 15 0 9 1 9 9 7 9 1 2
5 9 7 9 13 2
9 9 4 13 3 3 9 9 13 2
12 9 0 9 13 13 9 3 7 13 15 9 2
17 0 9 13 3 3 12 9 2 9 9 13 9 9 4 13 12 2
24 9 7 9 9 13 13 3 9 9 13 9 1 13 9 3 2 9 9 13 3 3 3 0 2
14 9 9 4 13 12 9 9 2 7 13 3 3 0 2
18 9 0 13 3 9 2 15 9 13 9 7 3 9 7 9 1 9 2
18 3 15 13 0 9 9 2 15 9 7 9 13 0 9 7 0 9 2
8 9 13 13 3 9 13 9 2
19 9 9 13 9 9 9 13 9 9 16 15 9 13 13 13 9 0 9 2
12 9 9 13 3 9 2 9 7 0 13 9 2
14 0 9 13 9 3 3 3 9 7 3 3 9 9 2
27 9 9 7 9 2 15 13 13 9 2 13 7 15 9 13 2 16 9 13 13 0 9 9 1 0 9 2
15 9 13 9 1 13 3 13 9 2 7 15 4 13 9 2
27 9 9 4 13 7 13 0 0 9 2 11 11 2 11 11 2 11 11 11 7 11 9 13 0 11 9 2
11 9 1 9 13 9 2 9 7 15 9 2
18 11 9 9 13 11 11 2 12 2 12 2 2 15 13 3 11 11 2
20 11 13 3 15 3 13 0 9 2 15 13 9 12 3 12 9 1 11 1 2
10 0 9 11 13 9 12 13 9 9 2
10 9 13 3 3 9 2 3 9 12 2
9 13 9 13 0 11 9 9 9 2
12 11 9 13 15 12 9 11 9 2 11 9 2
16 9 13 9 13 12 9 2 9 9 5 9 7 9 5 9 2
8 0 9 4 3 13 0 9 2
6 9 12 9 13 9 2
21 11 13 11 9 11 9 2 15 13 3 9 9 7 15 13 0 9 3 9 1 2
18 11 9 13 7 13 3 13 9 2 15 13 9 1 12 9 7 9 2
7 11 11 9 2 3 11 9
14 3 0 9 11 11 4 3 9 1 13 9 11 9 2
10 9 13 11 7 9 9 12 13 9 2
18 11 13 13 9 13 9 9 2 7 13 13 3 0 2 0 9 2 2
11 15 1 15 13 0 13 9 11 11 1 2
5 11 13 3 11 2
19 11 4 13 9 12 2 7 0 11 11 11 13 15 15 9 0 9 9 2
2 9 12
15 11 9 12 9 9 9 12 13 13 9 2 9 7 9 2
4 15 9 13 2
9 9 7 9 7 9 13 12 9 2
8 3 11 7 11 13 12 9 2
14 11 11 13 0 9 2 15 13 9 1 9 3 9 2
8 1 9 9 4 13 9 9 2
10 9 9 13 0 9 11 11 9 9 2
11 11 13 9 3 12 12 9 3 16 9 2
10 9 12 9 12 12 9 13 11 9 2
16 15 9 9 13 0 12 12 9 2 16 9 13 12 3 9 2
16 16 9 13 0 2 9 12 12 9 4 13 15 3 0 9 2
24 9 9 11 11 13 12 12 9 2 11 11 11 12 12 9 2 7 9 11 11 12 12 9 2
12 9 13 3 3 3 12 12 9 9 7 9 2
8 9 13 0 2 12 5 2 2
14 9 0 9 13 0 9 9 7 9 0 9 7 9 2
5 11 9 13 12 12
15 9 0 9 9 12 9 0 9 15 11 3 13 0 9 2
14 0 0 9 9 0 9 7 9 11 11 13 0 11 2
12 11 13 3 3 12 9 2 15 0 13 0 2
7 9 2 15 13 12 9 9
14 11 9 9 4 13 12 9 2 16 13 12 9 9 2
24 11 9 13 9 2 15 13 9 11 9 9 7 11 7 11 9 16 15 13 15 12 9 9 2
9 9 13 9 13 15 9 15 9 2
20 11 9 13 9 2 13 4 13 13 15 2 13 11 9 9 11 11 11 9 2
25 16 3 3 11 13 15 9 9 4 13 11 9 2 15 4 13 11 9 7 4 13 9 9 9 2
6 11 9 13 0 9 9
16 11 9 13 9 2 7 0 0 9 13 3 0 9 13 9 2
7 9 13 9 12 9 1 2
15 9 9 13 3 2 16 3 13 12 9 9 3 9 9 2
8 3 13 0 0 9 0 9 2
8 11 9 13 9 9 13 0 2
9 9 13 9 9 15 9 0 9 2
12 15 9 13 13 9 9 7 9 0 9 9 2
37 11 9 9 9 12 9 13 11 11 13 2 2 3 13 9 2 15 13 3 13 9 7 9 12 7 15 9 2 15 13 9 2 9 7 9 2 2
15 11 1 11 9 13 13 9 1 13 3 3 0 9 9 2
3 11 9 9
21 11 2 11 2 11 9 2 11 9 2 9 9 7 9 13 9 11 0 0 9 2
7 11 13 9 3 9 1 2
10 9 0 9 13 3 9 11 0 9 2
15 11 2 9 7 11 9 4 13 12 9 11 9 9 12 2
13 9 13 0 7 0 0 9 2 9 7 9 9 2
10 9 13 11 13 9 11 0 9 9 2
10 9 0 13 3 12 9 0 0 9 2
12 9 9 13 2 16 15 0 9 13 9 9 2
9 0 9 13 11 3 3 12 5 2
11 9 13 11 13 9 3 11 2 3 11 2
8 9 0 9 13 3 9 9 2
11 9 3 13 0 9 2 16 13 3 13 2
2 13 13
6 9 0 9 13 0 2
11 0 15 13 13 2 7 13 13 15 3 2
6 13 11 11 10 9 2
5 9 13 10 0 2
2 9 15
4 13 0 9 2
27 10 2 9 2 2 15 13 9 2 9 2 9 2 9 2 9 2 9 7 9 2 12 0 9 13 9 2
7 15 13 11 9 1 13 9
15 16 15 13 3 10 9 13 15 1 2 16 15 13 13 2
6 9 13 0 7 0 2
5 13 15 3 0 2
3 10 9 2
12 11 13 9 2 15 13 13 9 3 13 9 2
8 9 13 3 0 9 7 9 2
12 7 13 15 13 10 9 2 16 13 13 0 2
2 0 9
7 10 9 13 0 16 10 9
20 15 3 13 2 16 9 13 3 3 2 10 9 15 13 7 15 3 13 13 2
10 0 0 9 13 13 0 0 7 0 2
10 7 15 13 13 0 0 7 0 9 2
8 16 13 13 2 3 13 13 2
16 3 15 13 3 3 11 11 15 13 11 13 11 12 9 1 2
8 3 0 10 9 9 13 9 2
3 13 10 3
3 11 13 2
4 9 13 9 13
2 9 9
15 0 9 13 13 13 15 13 9 2 16 13 9 13 9 2
13 11 9 11 9 13 9 3 13 3 12 9 1 2
4 9 13 9 2
9 9 13 9 9 9 13 12 12 2
17 11 13 0 9 2 16 11 13 13 13 9 3 13 11 0 9 2
8 3 0 13 9 9 7 9 2
7 10 9 13 3 12 9 2
26 15 13 9 3 2 16 10 0 9 13 3 9 9 7 9 2 2 16 0 9 13 3 0 9 2 2
14 0 9 13 13 9 12 9 9 7 13 3 9 1 2
4 13 3 13 13
9 15 13 15 0 9 3 0 9 2
7 9 13 15 13 3 13 2
6 13 3 3 13 9 2
5 13 15 13 15 2
6 9 1 15 13 3 9
12 11 13 15 9 2 15 13 15 13 0 9 2
3 15 13 13
7 0 9 13 3 9 1 2
11 0 9 9 13 9 2 7 13 9 9 2
5 11 13 3 13 2
12 16 9 13 13 3 2 9 13 13 13 3 2
12 9 11 2 13 3 13 15 2 13 3 9 2
6 0 15 3 13 0 2
14 15 13 3 13 2 16 13 16 3 13 0 9 3 2
8 9 7 9 13 9 3 3 2
2 13 13
11 15 13 3 3 3 16 15 3 15 13 2
6 9 13 3 0 9 2
6 13 13 13 3 9 2
8 9 0 9 13 13 9 0 2
10 9 1 9 13 3 3 13 9 3 2
6 15 13 9 13 9 2
6 13 3 3 13 13 2
9 11 13 11 0 11 9 1 12 2
7 11 13 2 9 16 13 2
14 13 15 3 7 13 11 2 15 15 13 10 3 13 2
7 15 13 15 9 7 3 2
5 11 13 0 9 2
4 15 13 9 2
19 3 12 9 2 9 7 9 9 13 13 9 9 9 2 13 11 9 9 2
9 1 9 15 13 3 9 13 9 2
7 13 2 16 13 0 9 2
12 9 13 0 9 2 15 13 13 13 3 9 2
5 0 13 13 11 2
7 15 13 9 16 3 13 2
12 7 10 9 13 2 7 9 9 13 3 0 2
11 0 13 15 2 16 15 3 13 13 15 2
8 15 1 13 13 13 13 9 2
9 9 13 9 3 0 9 13 0 2
8 9 9 13 0 9 9 1 2
10 0 9 9 13 13 0 7 0 9 2
5 9 13 12 9 2
3 13 9 2
6 9 13 13 13 13 2
10 11 13 9 9 0 2 9 13 9 2
11 15 3 10 10 11 13 16 13 3 9 9
12 9 13 9 7 0 9 7 3 9 13 9 2
20 9 2 15 13 9 2 13 9 0 7 0 2 0 7 0 13 3 10 9 2
3 11 13 9
2 3 0
2 6 13
10 9 13 13 1 9 13 9 13 13 2
3 10 9 11
7 9 1 13 3 13 9 2
10 9 13 9 2 16 9 13 10 9 2
11 13 9 2 15 9 13 13 12 12 9 2
3 3 3 2
16 16 9 3 13 9 3 8 7 9 15 13 12 9 9 1 2
6 13 9 3 9 13 2
13 0 9 9 2 13 11 16 9 9 9 9 13 2
2 9 1
3 13 13 0
4 13 0 9 2
8 15 13 3 13 0 9 1 2
6 11 13 13 9 0 2
5 9 13 13 9 2
6 11 13 13 11 9 2
5 3 15 13 9 2
22 15 13 9 9 2 15 15 13 13 7 13 7 9 2 15 13 15 1 13 3 3 2
22 9 9 3 13 3 3 2 16 10 0 9 13 3 0 9 9 2 3 15 13 13 2
6 9 9 13 13 9 2
16 0 9 9 2 9 7 9 13 13 15 7 13 9 15 15 2
9 13 0 13 9 13 0 9 1 2
11 9 13 3 13 3 7 9 7 0 9 2
9 15 16 13 2 3 9 13 0 2
30 15 13 3 13 3 2 16 9 7 13 9 9 2 0 9 2 1 9 7 3 15 9 13 7 9 13 13 3 0 2
12 15 1 9 13 13 9 9 9 1 9 9 2
5 13 9 9 11 2
8 3 11 9 11 9 13 9 2
9 3 13 13 0 13 9 9 9 2
18 9 13 13 9 9 9 2 11 2 2 16 9 9 13 3 10 9 2
7 7 3 10 9 13 9 2
5 9 9 13 13 2
10 7 13 9 11 2 10 9 13 9 2
11 3 13 0 9 3 2 15 9 13 13 2
14 16 13 9 3 0 9 2 13 12 9 13 9 9 2
2 10 9
11 9 13 15 13 9 7 15 13 15 9 2
5 9 13 0 9 2
9 3 13 0 2 15 15 13 13 2
2 3 11
4 11 13 9 2
2 13 3
5 3 3 13 0 2
8 9 9 12 9 9 13 3 2
4 15 13 3 2
10 3 15 13 2 16 11 13 3 9 2
9 9 9 13 10 9 9 0 9 15
10 9 13 9 9 2 15 13 9 9 2
11 2 13 15 11 13 13 16 10 0 13 2
10 9 13 0 0 16 3 10 10 9 2
4 0 9 9 2
10 13 3 15 1 2 15 3 13 13 2
7 0 7 3 0 9 13 13
5 13 15 9 9 2
6 0 9 15 13 9 2
12 16 15 13 0 2 13 15 3 10 9 3 2
4 15 9 13 2
7 0 9 7 9 13 9 2
4 15 13 9 1
6 15 13 10 3 3 2
3 15 13 9
2 9 1
3 13 0 2
2 11 2
2 13 9
7 11 12 9 13 0 9 2
7 9 9 13 11 3 13 2
5 9 13 3 9 2
3 3 13 9
7 9 13 9 7 9 0 2
7 13 10 9 9 3 13 2
6 11 9 9 13 9 2
14 7 9 13 2 15 1 9 13 13 13 10 0 9 2
7 9 9 13 3 9 3 15
6 9 9 11 11 13 2
6 9 1 9 13 0 2
16 9 12 9 13 13 13 2 10 9 7 9 13 3 0 9 2
2 9 9
25 10 9 13 9 0 2 0 7 0 9 2 7 15 13 2 16 16 15 13 3 2 3 3 13 2
5 9 13 3 13 2
6 15 15 13 13 3 2
3 0 16 15
10 9 13 9 13 13 3 9 9 9 2
8 13 13 13 9 15 3 9 2
5 11 13 9 9 2
5 9 13 7 13 2
11 9 13 0 2 16 13 9 1 13 13 2
6 9 9 13 13 15 2
9 11 13 16 9 9 13 10 9 2
4 13 3 9 2
5 11 7 11 13 9
13 0 16 13 0 9 13 13 9 9 0 9 13 2
9 9 9 9 13 12 9 13 11 2
2 10 9
10 13 3 2 16 15 13 15 3 3 2
6 9 9 13 0 9 2
8 11 13 0 2 16 9 13 3
5 13 10 11 9 2
5 9 13 9 11 2
4 9 13 12 12
6 9 0 15 13 9 2
7 9 13 16 9 13 13 2
6 15 15 13 0 9 2
7 3 10 9 13 9 3 2
14 3 15 9 9 13 2 13 9 1 13 2 0 9 2
8 9 13 3 12 9 11 0 2
9 11 13 0 13 15 3 11 9 2
18 15 13 2 16 9 13 0 2 13 13 15 13 0 3 16 15 13 2
11 3 0 0 9 13 13 3 3 12 9 2
2 0 9
12 10 9 13 3 12 9 9 2 3 0 9 2
4 9 9 13 13
21 9 1 13 0 0 9 2 15 13 11 9 2 7 0 0 9 13 1 13 9 2
14 10 9 15 13 11 11 9 2 15 13 10 9 9 2
9 9 13 13 3 16 13 13 9 2
6 15 13 9 0 9 2
10 0 13 9 2 15 15 13 13 9 2
11 13 15 10 0 0 9 0 9 3 3 2
7 13 13 13 1 9 9 2
5 9 15 3 13 2
7 13 13 13 3 3 9 2
7 0 9 9 13 9 13 2
22 3 13 9 13 2 16 15 3 13 9 9 7 13 3 3 3 16 13 9 13 9 2
3 13 15 1
5 3 16 13 13 2
16 9 2 9 7 9 13 0 13 2 3 9 10 9 13 9 2
3 11 13 13
7 15 13 13 12 12 9 2
8 9 7 9 13 13 0 9 2
8 9 13 15 0 9 0 3 2
3 6 13 13
6 13 13 2 15 13 2
13 10 9 9 13 9 1 13 15 13 2 13 9 2
14 9 12 11 13 9 11 2 9 13 2 9 13 12 2
9 13 0 9 13 2 3 7 3 2
2 3 11
6 9 13 13 10 9 2
5 10 9 13 12 9
14 15 13 13 13 15 2 16 15 13 13 9 9 9 2
8 9 11 7 9 13 12 9 2
8 9 13 0 9 2 3 9 2
4 13 3 13 2
5 15 13 3 9 2
5 11 13 9 9 2
8 11 13 0 9 7 9 13 3
12 7 13 10 9 9 13 13 10 9 2 13 2
2 15 13
7 11 11 9 13 13 9 2
4 12 0 0 9
7 9 13 9 9 16 13 2
4 9 13 9 2
6 3 3 0 3 3 13
16 9 13 13 13 3 9 2 16 9 9 9 13 13 0 13 2
10 11 13 3 1 9 9 13 11 11 2
8 9 9 9 9 13 3 9 9
8 13 2 3 11 13 11 9 2
13 13 9 9 3 13 13 9 13 7 13 0 9 2
8 3 11 1 13 9 1 0 9
13 9 13 13 3 10 10 9 2 15 10 0 13 2
22 10 0 13 3 13 2 16 16 3 9 13 0 9 2 3 3 13 9 13 13 0 2
13 3 11 13 13 13 13 15 2 15 13 13 9 2
10 11 9 9 12 13 9 13 12 9 2
14 10 9 13 3 3 2 0 9 0 9 13 3 13 2
16 9 13 3 3 12 0 9 7 9 2 3 13 3 13 13 2
2 13 13
14 0 0 15 13 13 13 9 13 0 7 13 10 9 2
10 9 9 12 13 0 9 13 9 13 2
6 9 13 3 9 9 2
12 3 13 9 2 16 9 9 9 13 10 9 2
5 10 9 15 13 2
2 13 13
5 15 13 9 9 3
8 11 13 3 3 9 13 1 0
6 11 7 11 13 3 12
3 15 13 3
8 9 13 11 9 7 13 9 2
3 13 9 2
6 9 13 3 13 0 2
5 3 13 13 0 2
5 2 7 13 13 2
4 15 13 9 1
21 9 1 9 13 2 9 13 7 9 9 7 9 13 13 13 9 9 7 9 13 2
12 9 1 9 9 3 13 3 3 13 15 3 2
9 10 12 13 13 11 3 9 9 2
9 13 13 13 9 2 7 9 13 2
11 0 9 15 13 13 9 3 0 9 1 2
9 9 13 13 9 9 9 13 9 2
5 11 9 11 13 9
9 9 13 13 11 1 13 8 7 9
7 9 13 15 13 9 3 2
9 15 13 13 13 3 0 9 1 2
7 11 13 0 9 9 3 2
4 13 16 15 13
5 15 3 13 0 9
8 2 10 9 15 9 9 13 2
3 13 13 9
6 3 3 0 9 13 2
8 13 9 13 3 9 7 9 2
7 11 9 13 13 13 3 2
9 16 13 13 15 2 13 3 3 2
14 9 9 13 2 16 9 13 13 3 9 9 9 9 2
7 15 13 0 9 16 15 2
6 13 9 7 9 15 2
3 13 3 2
5 15 13 3 3 16
7 9 13 3 10 0 9 2
17 7 16 15 13 13 13 9 3 3 2 15 13 0 0 9 9 2
9 11 13 9 13 9 9 9 9 2
9 11 9 13 9 9 7 3 9 2
15 9 12 11 13 0 9 2 15 1 3 0 9 9 13 2
4 13 9 9 2
6 15 13 11 7 11 2
9 9 13 2 16 9 13 13 9 2
5 10 9 13 3 2
10 11 13 3 13 10 9 13 9 9 2
14 16 13 9 9 9 9 1 2 13 9 0 9 9 2
11 9 13 11 2 13 3 0 9 13 9 2
12 11 9 0 9 12 12 9 13 12 12 9 2
6 9 13 13 3 9 2
5 13 9 0 9 11
12 11 13 9 13 3 0 2 16 15 13 11 2
25 3 13 3 0 0 9 2 2 13 9 9 13 9 2 7 13 9 13 9 2 13 9 7 9 2
2 0 9
4 13 13 9 2
7 9 9 13 10 9 9 2
8 10 13 15 13 2 16 13 9
15 0 9 13 3 0 9 9 2 13 3 10 9 9 3 2
11 10 9 12 9 9 13 3 12 0 9 2
4 15 13 0 2
8 0 9 13 10 9 13 3 2
2 13 13
4 3 10 9 2
9 9 13 9 7 9 9 11 9 2
11 11 13 0 9 13 2 7 13 0 9 2
8 12 16 13 3 13 13 0 2
13 15 13 9 2 16 13 3 3 9 9 10 11 2
4 9 13 0 2
9 9 1 9 13 13 3 1 9 2
11 3 9 13 3 13 13 3 9 0 9 2
13 7 3 11 13 11 9 3 0 9 16 11 11 2
8 9 13 0 16 15 13 13 2
19 7 3 15 13 2 16 6 2 15 13 2 15 15 13 2 13 13 0 2
10 9 13 3 0 2 13 9 13 3 0
8 9 13 3 13 11 9 11 2
3 13 13 13
6 13 15 3 3 9 2
12 9 13 0 13 10 9 2 16 9 13 9 2
7 9 10 11 13 9 9 2
8 9 13 13 9 9 12 1 2
7 10 9 13 9 9 11 2
9 13 11 11 9 9 12 9 9 2
6 7 3 15 13 13 2
8 9 13 0 7 9 13 3 2
15 9 1 9 13 0 9 3 9 7 13 9 10 0 9 9
6 10 0 9 13 9 2
5 15 13 13 9 2
11 9 13 3 13 9 9 1 9 9 9 2
13 13 9 13 3 8 7 3 2 3 3 7 3 2
5 15 13 0 9 2
6 11 13 12 13 0 2
10 6 2 3 9 13 15 0 9 9 2
9 3 13 12 11 9 9 13 9 2
12 13 3 9 2 3 9 13 13 13 9 9 2
2 0 9
18 9 13 9 7 0 9 9 2 13 11 2 0 9 13 9 7 9 2
2 9 9
12 7 13 10 9 9 13 13 10 9 2 13 2
3 15 13 2
16 9 13 10 0 0 9 2 7 7 9 7 9 9 13 13 2
7 9 9 13 1 0 9 2
16 13 10 9 2 16 9 13 2 7 15 13 13 3 15 9 2
28 13 3 13 10 10 9 11 1 13 9 0 9 2 15 3 13 13 2 16 9 13 13 9 9 13 12 9 2
6 13 3 3 13 13 2
16 10 9 7 9 2 15 9 15 13 2 13 9 7 9 13 2
14 9 7 9 13 2 9 13 7 0 9 13 9 9 2
2 6 2
13 9 9 1 2 9 13 3 3 9 0 9 9 2
12 15 13 15 2 16 13 3 15 13 0 9 2
4 9 12 9 2
3 13 3 9
9 13 9 0 9 2 16 3 13 2
10 9 9 13 2 9 7 9 13 13 2
4 15 13 3 2
15 11 7 11 9 13 10 9 9 2 15 13 3 3 13 2
14 13 13 3 0 2 16 0 9 13 9 9 0 9 2
5 9 0 9 7 9
2 9 0
13 13 15 0 2 16 9 9 9 13 13 9 3 2
13 15 1 13 13 9 9 9 2 15 13 9 9 2
7 9 11 13 3 3 3 2
3 15 13 15
15 0 9 13 12 9 9 1 2 7 15 1 13 3 9 2
5 9 13 13 13 2
5 9 13 3 0 2
2 13 13
11 11 9 13 3 13 0 2 9 0 9 2
14 15 13 13 0 9 13 2 16 13 3 13 10 9 2
3 13 9 2
13 9 13 7 9 13 9 1 13 3 3 0 9 2
7 10 0 3 13 13 13 2
3 13 3 2
7 12 13 2 15 13 13 2
6 9 2 9 7 9 2
13 9 13 3 9 2 15 9 13 9 13 9 9 2
7 16 15 13 13 9 9 2
14 6 2 15 13 13 2 16 15 13 9 2 11 13 2
12 13 3 9 2 3 9 13 13 13 9 9 2
2 9 9
3 13 0 2
6 15 13 9 9 3 2
9 16 13 0 9 13 10 10 9 2
3 9 0 9
6 11 13 0 9 11 2
8 15 13 16 15 13 12 13 2
11 3 13 0 9 7 13 3 0 9 13 2
14 15 13 9 3 9 2 11 2 9 2 13 15 3 2
6 13 13 2 9 13 2
12 3 9 9 13 3 2 16 15 9 1 13 2
19 15 13 16 9 11 9 7 11 9 0 9 2 16 3 0 9 13 13 2
16 9 13 13 3 3 9 2 16 11 9 13 11 11 9 3 2
4 9 3 13 9
6 13 15 13 10 9 2
6 11 13 3 9 1 2
6 15 13 9 0 9 2
16 15 13 0 9 1 0 16 13 9 7 13 10 9 9 13 2
9 13 9 2 13 15 16 9 13 2
6 13 15 0 9 3 2
19 16 13 2 16 13 13 13 2 15 13 3 3 2 16 13 13 13 9 2
18 3 13 0 13 9 9 1 2 9 13 9 3 16 9 13 13 3 2
13 15 13 13 15 9 2 15 0 9 13 0 9 2
7 13 0 9 7 13 0 2
4 13 0 9 2
5 3 3 9 13 2
5 13 11 3 9 2
10 11 13 15 3 2 3 7 15 13 2
4 9 9 0 9
12 13 15 13 15 13 0 9 3 10 12 9 2
11 15 13 13 15 9 13 9 7 3 13 2
10 15 13 9 13 9 2 15 13 9 2
7 9 9 11 9 13 13 2
9 9 9 13 9 3 1 12 9 2
4 3 13 3 2
8 11 13 9 9 7 13 15 2
4 13 0 9 2
8 7 15 15 13 13 13 13 2
9 15 13 13 9 15 9 13 9 2
12 15 13 7 13 9 9 9 2 11 13 11 2
7 0 9 13 10 9 9 2
2 0 11
9 7 13 9 12 9 2 3 13 2
4 13 3 9 2
7 9 13 3 3 13 9 2
7 13 9 7 9 3 9 2
10 3 10 9 15 13 13 3 0 9 2
6 3 9 13 9 3 2
4 12 9 9 13
9 0 7 0 9 9 13 3 0 2
5 9 13 9 13 2
5 3 13 3 9 2
8 11 9 9 9 13 9 13 2
9 13 9 13 9 2 13 10 9 2
7 13 3 13 13 15 9 2
3 13 15 13
8 2 6 16 13 9 13 13 2
5 12 9 13 9 2
9 3 11 13 3 9 16 3 3 2
7 15 13 3 15 13 3 2
12 13 15 10 9 2 3 15 13 3 9 9 2
4 12 9 9 9
15 13 9 9 2 16 13 15 2 9 13 2 13 13 0 2
3 3 1 9
6 13 15 3 0 9 2
3 13 9 9
12 11 1 13 2 16 9 13 0 9 13 9 2
11 9 9 1 11 13 3 3 9 7 9 2
4 9 13 9 2
12 13 11 0 9 13 3 12 9 11 3 9 2
19 16 7 16 9 13 2 13 9 9 9 3 10 1 9 2 9 7 0 2
2 10 9
13 9 13 11 9 11 2 15 13 0 9 16 11 2
9 9 13 9 13 9 13 2 16 2
15 9 13 3 2 16 9 13 0 13 2 16 15 13 13 2
7 9 13 2 16 13 13 2
6 3 15 13 3 13 2
6 3 15 13 10 9 9
9 9 13 10 9 9 13 0 9 2
3 9 13 2
15 7 3 9 13 9 2 16 13 3 11 2 3 3 11 2
3 13 9 2
11 0 9 0 9 13 9 1 13 15 1 2
14 3 13 15 2 16 9 13 3 0 0 13 0 9 2
14 13 9 13 10 9 3 9 7 13 15 1 10 9 2
9 15 13 12 0 9 13 13 9 2
14 3 0 9 15 13 3 13 3 2 9 10 9 0 2
5 11 13 3 0 9
7 9 1 13 13 12 9 2
11 9 13 10 9 2 15 13 3 9 13 9
4 10 13 9 2
7 15 13 13 15 13 9 2
5 15 13 16 15 13
9 3 3 2 13 15 0 9 3 2
5 3 13 3 9 2
8 0 9 13 0 9 9 9 13
7 13 11 13 3 9 9 2
8 9 13 9 2 13 2 9 2
14 15 13 0 13 15 2 3 9 2 9 7 3 9 2
15 15 13 0 9 9 2 15 13 13 2 7 16 13 13 2
4 15 13 13 2
5 10 15 13 15 2
2 9 9
13 15 13 9 3 13 13 9 2 3 7 9 1 2
16 7 10 10 9 13 10 9 15 13 16 16 15 13 9 0 9
7 13 3 2 16 13 15 2
9 10 9 15 3 13 9 3 9 2
16 11 13 13 2 16 15 13 13 10 9 13 9 0 9 9 2
17 9 13 3 10 9 6 16 13 15 16 9 13 15 13 7 9 2
9 7 9 7 9 13 0 13 9 2
3 15 13 2
4 9 9 11 9
6 3 13 15 3 3 2
3 13 11 2
5 3 15 13 15 2
3 9 11 2
2 12 12
4 13 9 9 2
4 9 13 13 9
10 0 9 2 15 3 13 3 0 13 2
13 13 3 15 0 13 15 13 2 15 13 9 0 2
2 13 9
14 0 9 13 9 7 13 9 15 2 13 9 10 9 2
8 0 9 1 9 13 11 11 2
2 9 9
5 13 0 9 12 2
16 0 9 13 11 15 2 16 9 7 0 9 13 3 0 9 2
11 9 13 9 11 9 2 15 15 13 13 2
9 3 13 13 13 9 2 11 13 2
10 13 13 13 7 13 7 13 0 9 2
8 13 9 7 13 9 9 13 2
7 3 15 13 0 11 13 2
7 9 13 13 9 13 9 2
16 7 3 13 2 16 13 13 13 2 13 10 9 2 13 3 2
7 0 9 9 13 11 0 2
4 13 13 9 2
14 9 13 10 9 2 16 10 9 13 3 0 9 3 2
11 7 15 13 3 10 0 3 13 15 9 2
12 15 13 3 13 15 15 13 15 2 11 13 2
2 9 15
13 3 13 2 15 13 3 2 15 13 7 13 0 2
5 13 15 13 9 2
6 3 10 15 13 13 2
4 2 13 3 2
8 15 1 13 13 15 3 3 2
8 13 13 0 9 13 9 9 2
8 11 7 11 13 3 0 9 2
9 0 9 13 0 2 16 9 13 2
12 10 9 15 13 15 2 3 15 13 10 9 2
6 12 9 9 13 9 2
10 3 13 11 2 3 13 13 15 1 2
15 9 13 9 9 7 3 13 3 9 2 11 13 0 9 2
16 9 13 12 2 7 11 13 13 16 15 13 13 11 9 1 2
20 10 10 9 13 13 0 13 10 9 16 15 13 13 10 9 15 3 9 13 2
8 3 9 13 13 12 9 9 2
15 9 13 13 3 13 13 9 2 13 15 13 15 3 3 2
14 11 11 13 9 1 9 11 11 7 9 11 11 9 2
14 9 1 9 13 3 13 7 13 10 9 0 9 1 2
16 9 1 11 13 0 3 12 2 15 1 11 13 12 0 9 2
1 11
7 10 9 13 13 10 9 2
10 9 3 13 3 7 9 13 9 9 2
3 13 3 2
14 15 13 2 16 13 13 9 2 16 0 13 9 9 2
9 11 13 10 9 16 15 11 13 2
3 9 13 2
10 15 13 9 2 13 3 7 2 9 2
5 13 15 13 15 2
12 15 13 0 9 13 15 13 10 0 9 3 2
5 15 13 3 9 2
17 13 13 2 16 9 0 12 2 12 2 12 9 13 9 11 1 2
7 15 13 2 16 15 13 2
15 9 13 13 0 9 2 15 1 0 9 13 13 0 9 2
3 9 3 2
9 11 13 13 11 7 15 0 9 2
12 9 13 9 2 16 3 8 7 0 9 13 2
10 11 13 9 13 3 9 0 9 9 2
11 16 9 13 13 13 3 2 3 3 13 2
3 0 9 2
5 9 13 13 0 2
9 3 9 13 15 2 13 0 13 9
6 0 9 11 13 9 2
8 15 13 13 3 9 3 3 2
10 16 9 13 2 3 15 13 10 9 2
2 15 1
5 13 3 9 13 9
2 13 9
5 9 13 3 13 2
8 9 13 13 3 3 0 9 2
3 13 9 1
7 11 13 9 9 13 9 2
13 7 9 13 13 10 0 9 2 15 15 13 9 2
11 9 13 15 16 13 13 3 13 0 9 2
2 3 9
2 13 3
5 9 13 9 9 2
12 10 0 0 13 15 13 9 7 9 0 9 2
4 13 15 3 2
13 9 13 9 2 10 9 13 3 3 12 12 9 2
3 0 9 0
9 13 3 9 2 0 13 3 13 2
4 15 13 9 13
12 13 13 0 9 9 2 16 13 9 13 3 2
8 15 3 3 13 10 9 3 9
7 15 13 12 3 15 13 2
3 3 13 9
2 0 9
7 15 13 9 2 15 13 2
4 9 13 9 2
13 13 10 9 3 2 13 13 3 2 7 13 3 2
6 13 15 10 0 9 2
7 8 7 9 13 9 3 2
14 16 9 13 12 9 9 2 15 13 3 13 15 9 2
10 3 10 9 13 3 13 9 9 9 0
2 10 9
6 10 9 15 13 13 2
20 3 12 9 13 0 2 16 11 9 1 9 13 9 2 10 9 10 9 13 2
23 10 9 13 11 9 12 9 2 15 13 0 9 13 9 9 2 16 3 11 13 13 3 2
6 0 13 13 10 9 2
5 11 13 9 9 2
24 11 7 11 2 11 7 11 9 13 9 2 15 13 9 2 7 3 0 13 9 2 0 9 2
16 11 9 9 7 9 13 0 9 13 3 9 7 9 9 1 2
12 7 9 13 15 16 10 9 13 13 3 9 2
7 9 13 13 0 7 0 2
5 15 13 3 9 2
12 9 11 11 13 11 13 15 13 9 9 3 2
7 15 13 3 13 15 13 2
7 13 15 3 13 0 1 2
20 16 11 13 9 2 16 9 13 7 16 0 9 13 13 2 13 13 15 16 2
6 0 3 13 10 9 2
3 0 0 9
11 11 13 0 9 2 9 9 2 9 9 2
9 3 3 13 13 3 16 9 13 2
3 15 1 2
4 9 13 11 2
10 13 13 9 2 9 7 9 3 13 2
3 15 13 9
3 10 9 1
7 9 13 9 12 9 1 2
2 10 9
9 9 11 7 11 13 3 9 0 2
11 13 13 0 9 2 7 15 13 3 13 2
6 9 13 13 9 1 2
15 16 9 13 13 9 9 2 9 13 9 2 7 13 3 2
6 9 13 0 9 9 2
2 13 2
18 9 13 9 0 2 0 7 0 9 7 15 3 11 2 11 7 11 2
8 9 13 13 13 3 12 9 2
12 16 15 9 13 9 2 3 13 15 13 9 2
4 13 11 10 9
5 9 13 10 9 2
30 3 13 9 9 2 15 3 13 13 9 9 9 0 9 7 10 9 10 0 13 13 2 13 1 2 3 9 9 9 2
14 16 13 2 15 13 13 3 13 9 9 7 9 9 2
7 11 11 13 13 0 9 2
8 15 13 13 13 2 13 13 2
9 9 15 13 3 10 7 9 9 2
5 11 13 9 13 2
12 16 0 0 9 13 0 2 13 9 13 9 2
15 13 15 0 2 11 13 11 13 2 13 0 9 9 2 2
2 0 9
20 9 13 13 3 2 16 9 13 13 9 0 9 9 2 15 9 9 13 13 2
9 3 13 9 13 3 3 3 3 2
14 13 9 0 9 9 2 9 7 9 7 9 9 9 2
10 9 13 3 13 2 16 7 16 13 2
8 3 15 0 13 16 13 13 15
16 6 2 13 13 3 3 2 16 10 15 13 10 9 16 15 2
18 16 15 13 9 9 2 9 13 3 11 7 15 13 3 3 15 1 2
5 9 13 9 1 2
22 10 15 13 9 9 15 1 2 16 13 9 3 3 11 9 2 13 3 3 9 1 2
13 9 13 13 13 9 9 2 16 3 13 13 13 2
8 13 13 13 15 16 9 13 9
6 15 13 15 9 3 2
6 9 9 13 0 0 2
10 15 13 13 0 9 2 15 13 15 2
5 9 7 10 0 9
7 9 13 3 0 0 9 2
16 13 3 3 16 11 9 13 0 9 3 0 7 3 13 9 2
14 3 3 3 9 9 13 10 0 9 7 9 7 9 2
5 13 9 10 9 2
4 9 13 3 13
10 7 8 15 9 3 16 15 13 9 2
11 11 9 13 15 9 13 13 13 9 1 2
5 9 13 9 1 2
4 6 15 13 3
8 9 9 3 13 9 11 9 2
9 9 13 9 2 10 9 9 13 2
7 3 13 9 1 0 9 2
4 9 12 1 2
2 13 0
14 11 11 13 2 9 2 11 9 13 15 3 13 9 2
3 13 15 2
5 3 15 13 7 2
2 13 12
3 13 15 2
6 15 13 13 9 9 2
4 7 9 13 2
12 10 9 7 9 13 3 3 0 0 9 3 2
6 0 0 9 13 3 2
31 13 9 7 13 9 13 9 2 10 9 13 13 9 3 16 3 16 13 13 7 13 9 2 0 9 13 2 16 13 15 2
6 0 9 1 9 13 2
12 9 13 3 13 9 9 2 7 13 9 9 2
8 10 15 11 9 13 16 9 2
7 9 13 2 7 13 13 2
3 9 13 12
14 15 13 3 3 15 2 16 13 13 9 0 0 9 2
9 15 13 0 9 10 9 2 3 2
8 15 13 13 11 2 7 3 15
15 3 15 3 9 13 3 3 3 16 3 13 12 9 9 2
15 11 13 9 3 9 13 9 13 2 16 13 15 13 13 2
6 9 13 13 3 3 2
2 3 2
10 9 15 13 13 2 3 12 9 2 2
5 3 13 3 13 2
15 15 13 3 3 3 11 2 3 3 11 2 3 3 9 2
6 13 15 15 13 9 2
10 15 13 3 9 1 2 13 15 13 2
12 9 9 13 13 9 13 9 9 7 9 9 2
6 9 13 16 13 9 2
4 9 13 3 2
6 0 9 13 3 0 2
6 13 16 13 3 9 2
17 3 9 13 13 0 2 3 13 7 13 13 10 9 1 13 15 2
5 0 9 13 13 2
16 9 13 13 10 11 13 9 2 16 3 9 13 3 9 13 2
9 3 11 2 11 13 9 3 11 2
4 10 9 9 2
13 9 9 13 13 0 0 9 2 7 3 13 15 2
14 13 3 3 11 2 16 13 3 15 2 16 13 13 2
5 11 11 13 9 2
5 9 13 9 1 2
5 13 2 13 9 9
13 3 15 13 9 2 13 15 3 13 0 9 15 2
9 15 15 15 13 13 9 1 0 2
13 16 9 13 7 13 2 10 10 9 13 13 3 2
4 9 13 13 0
2 15 13
23 0 3 3 13 15 2 16 9 13 15 16 15 0 11 2 11 7 13 9 11 9 9 2
14 13 3 2 16 9 9 13 2 16 9 13 3 3 2
11 13 3 11 2 15 9 9 13 3 3 2
72 9 10 9 9 7 7 3 15 13 3 3 0 3 16 15 13 3 3 7 3 3 15 3 3 13 0 3 0 13 7 3 15 13 3 15 9 3 0 13 9 7 15 13 13 3 0 9 16 3 13 13 13 15 3 3 3 13 10 9 7 15 13 9 1 10 9 3 3 7 0 7 2
8 13 9 13 9 9 7 9 2
4 9 15 13 9
16 15 13 13 3 3 3 2 11 13 2 16 13 3 0 9 2
2 0 9
4 9 13 0 2
10 9 13 9 9 2 15 9 13 0 2
10 3 13 0 9 11 9 9 11 11 2
17 9 9 11 13 13 10 9 10 9 2 13 15 3 13 12 9 2
11 15 13 13 9 2 0 2 9 7 9 2
5 9 13 9 9 2
3 13 3 2
2 13 9
9 10 0 13 3 3 9 0 9 2
4 16 15 13 13
5 13 15 9 0 2
8 9 0 9 13 13 9 0 2
4 0 16 13 2
2 9 9
10 9 12 9 2 0 7 0 13 15 2
11 6 2 13 3 15 13 3 1 10 9 2
5 6 13 3 3 2
14 15 3 13 15 2 16 8 7 9 9 13 9 13 2
8 3 13 11 13 0 3 9 2
6 9 0 13 12 9 2
10 13 13 9 2 11 2 2 7 9 2
8 13 13 15 13 13 0 9 2
16 13 9 0 9 13 0 13 0 9 7 3 0 13 0 0 2
13 10 9 13 16 9 9 13 9 2 3 3 0 2
8 11 11 13 13 3 13 9 2
12 13 9 1 11 13 13 0 11 9 9 9 2
3 13 9 2
12 15 13 15 11 15 2 16 13 15 15 13 2
10 16 13 13 9 0 2 13 13 15 2
8 10 10 9 13 13 0 9 2
3 15 13 3
10 3 11 13 3 9 13 7 13 9 2
2 13 3
11 0 3 2 10 9 13 3 13 2 11 2
7 11 12 9 13 13 9 2
5 13 13 13 10 9
16 0 9 9 11 13 15 2 16 9 9 9 9 1 13 11 2
10 0 11 9 13 3 9 1 9 9 2
18 11 9 9 3 13 11 13 11 2 11 13 3 13 11 1 3 11 2
9 15 13 9 13 9 7 13 15 2
5 13 3 3 11 2
5 13 9 13 9 2
6 9 1 13 13 3 2
14 3 16 13 9 9 2 3 9 13 9 13 0 13 2
15 11 9 13 10 10 9 9 0 2 0 2 0 7 0 2
3 2 15 2
9 13 2 16 15 9 13 3 0 2
13 15 13 2 10 9 9 2 13 11 11 11 9 2
6 9 13 0 9 0 9
5 15 13 3 9 2
4 9 13 13 2
20 3 15 13 13 12 2 3 3 12 9 2 3 3 7 0 9 3 9 1 2
6 3 2 3 13 11 2
14 9 13 13 15 2 7 13 13 2 13 15 3 15 2
6 15 13 13 15 9 2
8 3 3 9 13 13 9 9 2
2 13 13
5 9 13 9 13 2
13 0 0 9 9 13 1 15 15 2 13 9 9 2
3 9 13 2
10 15 13 11 13 13 3 16 9 1 2
2 13 13
10 9 9 9 13 3 13 2 13 11 2
19 3 15 13 9 9 2 7 16 13 3 15 13 9 2 15 3 13 9 2
6 6 10 9 13 13 2
10 11 13 7 13 0 2 7 0 3 2
6 3 13 10 9 9 2
17 0 9 13 0 9 9 2 13 15 2 13 0 15 7 13 9 2
8 10 12 0 3 13 1 9 2
11 9 13 13 3 16 9 15 13 15 13 2
6 11 11 0 9 13 2
5 3 0 9 0 2
6 0 9 15 3 13 2
5 3 13 9 13 2
7 0 9 9 13 3 11 2
11 0 9 13 3 11 9 2 3 0 9 2
13 9 9 13 11 0 9 2 16 11 9 13 0 2
4 13 15 9 2
5 0 9 7 10 9
22 9 13 0 3 13 2 2 13 13 10 9 2 15 9 7 9 13 13 9 0 2 2
8 15 3 3 13 0 13 3 2
13 2 13 15 13 13 13 10 9 2 15 13 13 2
2 10 0
3 13 11 2
3 9 13 13
13 11 13 3 9 9 0 9 7 10 9 9 12 2
5 9 13 3 9 2
7 9 1 15 3 13 13 2
3 13 3 0
15 16 9 9 9 13 3 0 2 9 13 13 13 0 9 2
26 9 13 2 16 15 13 13 10 9 2 13 2 7 13 0 9 2 16 15 3 13 10 9 3 13 2
14 15 13 3 0 2 16 10 9 13 9 2 16 13 2
21 15 13 13 15 11 1 2 7 10 0 9 2 15 15 9 13 0 9 9 1 2
12 9 13 2 16 9 13 10 9 11 0 9 2
2 9 11
14 9 13 13 3 9 13 3 9 2 16 13 0 9 2
6 9 13 3 3 3 2
4 9 13 9 2
7 13 3 9 9 9 9 2
14 13 3 10 11 2 15 15 1 13 13 3 9 13 2
15 9 13 13 9 1 13 15 2 16 9 13 9 0 9 2
9 15 13 9 13 9 7 13 15 2
6 16 15 3 9 13 2
9 11 13 0 9 13 13 9 9 2
10 6 2 15 16 13 16 15 13 9 2
2 0 9
17 0 13 9 11 11 11 2 15 13 13 0 13 9 9 12 1 2
8 3 9 13 13 9 15 3 2
14 11 11 13 3 15 2 16 10 9 13 13 13 15 2
8 13 15 3 12 12 9 9 2
9 16 9 13 2 15 13 13 3 2
5 9 13 9 15 2
5 16 3 13 0 2
3 13 0 2
7 9 13 3 10 9 1 2
13 0 9 9 13 2 10 15 13 9 7 13 9 2
11 11 3 13 11 7 11 11 13 9 9 2
12 13 15 10 9 3 13 10 0 9 10 10 9
4 9 13 9 9
10 0 9 15 9 13 0 3 10 9 2
7 9 15 13 2 11 13 2
9 15 13 10 9 3 11 9 11 2
6 15 13 15 13 3 2
5 13 3 10 9 2
4 9 13 11 2
30 11 2 13 9 9 9 7 9 9 2 2 13 3 11 2 0 9 15 13 13 0 2 7 13 3 11 11 0 9 2
4 9 13 3 3
10 1 9 9 8 11 13 11 9 9 2
5 13 0 9 7 9
7 0 0 10 10 0 9 2
18 10 9 11 13 0 9 13 10 0 9 2 15 10 9 13 13 9 2
11 10 9 13 13 0 9 2 10 9 13 2
15 15 13 13 13 3 3 2 7 9 7 9 9 13 9 2
13 11 11 1 0 9 13 0 9 13 13 13 11 2
7 2 13 3 15 15 13 2
8 9 13 9 1 13 13 9 2
3 11 9 11
18 9 2 13 2 3 3 16 2 3 2 11 15 13 13 2 13 3 2
6 0 15 13 13 9 2
5 13 13 3 13 2
15 15 13 3 9 3 7 3 3 9 13 7 9 13 1 2
6 9 13 9 7 0 9
8 11 9 13 3 15 16 9 2
13 7 13 13 2 7 13 12 9 2 10 11 9 2
4 13 3 13 2
8 13 13 0 9 9 3 3 2
3 15 13 9
17 10 0 9 13 13 13 2 16 11 15 13 10 9 13 0 9 2
5 9 13 3 3 2
11 13 2 16 15 13 15 2 7 13 3 2
8 9 9 13 13 3 13 9 2
5 16 15 3 13 13
6 9 13 0 9 3 2
2 0 0
14 9 1 2 11 13 11 0 9 7 0 9 9 2 2
11 11 11 16 13 13 0 0 9 13 9 2
4 9 13 9 2
10 11 13 9 2 13 3 13 10 9 2
2 9 9
15 11 13 9 2 16 9 9 13 3 3 9 16 9 9 2
16 13 3 9 9 0 9 13 9 7 9 10 9 10 9 9 2
9 13 11 13 13 9 13 9 9 2
3 11 13 9
10 9 13 11 13 0 9 11 9 9 2
8 6 16 15 13 3 13 3 2
21 9 9 11 13 13 13 2 7 12 9 15 13 3 3 2 9 15 13 13 3 2
5 15 13 13 9 2
7 3 9 13 3 3 13 2
5 9 13 9 9 2
16 9 13 9 13 13 9 2 16 9 13 0 0 7 13 9 2
10 16 13 13 3 2 15 13 13 0 2
12 0 2 0 2 16 13 13 0 9 13 11 2
3 15 13 2
17 16 13 9 9 9 9 2 9 13 0 9 16 13 12 9 0 2
11 9 1 11 13 2 16 15 13 3 9 2
7 15 13 3 0 16 15 2
3 13 3 2
10 12 11 9 9 13 13 0 9 9 2
3 13 15 3
6 9 13 3 13 9 2
3 13 9 9
4 13 13 9 2
2 0 9
9 9 7 9 13 13 13 0 9 2
14 2 13 10 9 3 15 10 9 13 2 2 11 13 2
8 3 0 13 2 15 11 13 2
16 0 9 7 9 13 13 3 3 0 2 16 13 0 16 9 9
4 9 13 3 2
14 9 1 13 0 9 13 9 1 9 3 12 9 9 2
13 9 13 13 13 11 9 3 7 13 0 9 9 2
7 0 9 9 13 13 3 2
11 9 13 0 9 9 2 15 13 9 9 2
2 3 3
2 9 9
10 9 13 9 13 13 0 9 15 1 2
8 9 13 3 13 3 9 9 2
3 9 13 15
4 9 13 9 2
11 9 1 0 9 13 9 7 0 9 1 2
8 9 9 13 0 16 9 9 2
11 3 9 13 12 9 0 9 0 9 11 2
10 13 0 2 16 13 13 9 0 9 2
5 13 3 16 13 2
7 9 13 13 7 13 9 2
14 13 3 16 0 13 2 13 9 9 7 16 3 0 2
13 0 9 1 10 9 1 13 13 9 3 12 9 2
2 13 9
7 3 9 13 12 9 3 2
14 3 9 9 13 13 3 13 9 9 13 3 3 3 2
3 0 9 12
10 16 15 13 9 2 15 13 3 3 2
8 9 11 11 13 3 9 9 2
7 13 2 10 9 3 13 2
5 16 13 10 9 3
12 3 9 13 3 13 2 7 9 13 10 9 2
4 9 13 0 2
11 9 9 9 11 13 9 13 3 9 13 2
2 9 9
8 9 15 13 15 15 3 13 2
11 15 13 3 0 13 2 16 15 13 9 2
12 0 9 9 9 7 9 9 13 3 3 13 2
6 11 9 9 9 9 9
12 0 2 9 7 9 13 13 0 9 0 9 2
19 15 13 3 3 0 7 3 13 15 7 13 9 7 9 7 10 0 7 2
5 15 15 13 0 2
11 9 1 9 13 13 9 0 8 7 9 2
4 9 3 9 2
20 13 0 9 13 10 10 9 9 3 16 11 13 9 13 13 15 13 9 9 2
4 13 9 13 3
3 3 7 3
13 9 15 13 13 0 9 2 16 3 13 13 13 2
3 9 13 13
3 13 0 2
11 9 9 13 2 16 9 13 3 12 9 2
4 9 13 3 13
12 16 0 9 13 9 11 13 0 9 9 9 2
17 16 9 13 2 3 10 9 13 0 9 9 7 15 2 9 13 2
5 9 15 13 0 2
6 10 9 13 3 0 2
16 11 13 3 3 13 2 7 3 13 3 13 13 3 16 3 2
11 13 15 13 0 9 10 9 3 0 9 2
3 13 9 9
8 13 9 3 3 3 16 9 2
5 15 13 0 16 9
5 9 13 3 9 1
6 9 13 1 9 13 2
6 3 0 13 13 9 2
2 13 13
8 3 10 9 11 7 11 13 2
11 3 0 7 0 9 13 0 3 13 9 2
10 16 9 9 13 13 2 9 13 13 0
12 9 13 3 3 13 2 13 9 0 11 9 2
2 13 13
7 13 13 16 9 13 9 2
8 3 9 13 3 3 3 13 2
5 13 15 10 9 2
8 9 13 11 3 3 7 3 2
4 13 9 9 2
13 9 13 3 13 3 12 9 2 16 9 13 3 2
13 16 9 13 0 9 2 13 2 16 13 15 0 2
14 9 9 9 13 13 15 2 16 9 13 0 9 9 2
9 9 13 10 0 0 9 3 3 2
35 3 16 13 11 9 0 9 2 13 2 16 13 13 15 2 13 9 0 9 2 11 2 9 2 11 8 7 9 2 9 11 11 2 12 2
7 15 13 3 0 13 9 2
5 0 9 13 0 2
9 16 13 3 2 15 13 13 0 2
4 10 0 0 9
3 9 13 3
12 9 13 13 3 3 16 13 2 9 13 13 2
4 0 9 7 9
9 3 11 9 13 13 10 0 0 2
2 13 13
12 0 9 2 7 9 15 2 16 3 13 15 2
9 2 7 9 2 15 13 13 9 2
4 15 15 13 2
12 3 3 12 2 7 13 3 12 2 11 13 2
8 9 13 8 7 9 9 9 2
8 16 13 13 2 13 13 9 2
3 15 13 13
7 0 10 9 13 9 9 2
6 9 13 9 13 9 2
7 9 13 3 3 9 1 2
9 9 13 7 10 0 9 13 9 2
12 13 0 13 9 16 9 13 3 12 9 9 2
7 6 6 3 2 11 13 2
3 3 15 13
5 9 13 15 1 2
15 7 13 13 16 3 15 13 13 13 10 10 9 10 9 2
16 2 13 15 13 2 7 3 15 15 13 13 2 2 11 13 2
5 13 2 16 13 2
5 15 13 13 9 2
8 11 7 9 9 13 3 9 2
4 15 13 3 2
17 15 3 13 9 13 0 2 3 9 2 15 15 13 13 9 1 2
3 13 13 13
5 15 13 9 0 9
4 15 15 13 2
12 9 1 9 13 7 3 15 13 13 13 9 2
14 13 0 9 2 16 0 9 13 12 0 9 9 1 2
6 15 13 13 0 9 2
11 9 13 3 9 11 11 0 13 0 9 2
5 11 13 15 9 2
21 9 13 12 9 0 16 0 9 9 7 3 9 0 16 0 11 9 1 13 9 2
7 3 15 13 0 13 9 2
12 0 9 13 13 9 13 9 13 10 12 9 2
13 11 13 3 9 9 2 3 16 15 13 13 0 2
11 15 13 10 12 9 1 13 9 7 9 2
9 9 13 0 7 0 2 3 13 2
6 9 13 3 10 0 9
8 9 13 9 7 9 13 9 2
18 7 3 0 9 2 9 9 2 13 13 9 13 9 13 9 3 3 2
5 15 13 3 3 2
11 9 13 13 0 9 2 15 13 3 9 2
12 7 15 13 3 0 16 3 9 13 3 3 2
7 9 13 3 12 12 9 2
23 2 9 9 13 13 2 16 11 13 13 9 13 2 2 11 0 9 9 11 11 13 9 2
6 15 13 3 0 1 2
15 9 13 3 13 0 13 9 3 3 0 9 2 9 13 2
12 12 0 9 13 13 3 0 9 2 11 13 2
16 9 1 13 9 13 15 2 13 12 9 7 11 9 1 9 2
10 15 13 3 3 0 7 3 0 9 2
8 13 9 7 13 15 3 3 2
2 9 9
5 13 9 9 1 2
5 15 13 13 9 2
7 13 0 2 7 13 13 2
17 15 13 3 15 13 0 3 0 9 9 13 0 0 0 0 0 0
4 3 12 3 2
22 15 13 13 13 0 9 3 2 16 15 13 0 2 7 15 1 2 16 15 13 9 2
21 7 10 10 3 9 13 12 0 0 9 15 16 15 13 10 9 15 15 3 13 2
4 15 11 13 2
3 13 3 2
6 9 0 9 13 9 2
5 13 15 0 9 2
4 0 15 13 2
3 3 15 1
6 13 3 3 0 9 2
7 13 9 2 16 3 13 2
6 9 9 9 13 3 2
7 9 13 13 3 0 9 2
6 10 9 9 15 13 2
14 13 11 13 9 13 2 7 13 13 13 9 3 9 2
11 13 13 15 2 16 9 11 13 13 13 2
7 15 13 12 13 10 0 2
2 9 9
6 13 13 16 13 3 13
15 9 13 3 3 2 13 13 0 13 13 9 1 0 9 2
32 6 16 13 3 3 3 3 10 9 1 3 3 15 13 13 9 3 9 7 7 3 15 13 10 9 3 9 3 6 15 13 13
10 11 1 11 13 13 9 3 0 9 2
12 15 13 13 9 2 15 13 13 9 0 9 2
15 11 13 3 0 9 7 9 2 15 9 13 3 3 13 2
9 3 15 13 10 9 1 0 9 2
6 13 9 11 13 0 9
3 15 3 2
5 13 13 3 12 2
5 13 9 9 13 2
11 0 13 13 3 9 7 9 13 0 9 2
10 15 13 0 9 3 16 13 13 9 2
3 13 13 13
2 0 9
11 9 12 7 9 1 15 13 13 15 12 2
4 13 9 3 2
5 15 13 13 3 2
12 9 13 0 9 13 9 3 3 13 9 1 2
10 11 13 0 9 2 3 0 9 1 2
4 13 13 15 2
14 13 15 13 2 10 9 2 13 0 9 3 10 9 2
12 16 0 13 2 15 13 3 15 1 13 13 2
7 13 2 16 13 13 13 2
10 9 13 3 0 9 9 9 3 9 2
12 9 11 2 13 3 2 13 9 9 9 9 2
6 9 13 9 13 9 2
8 9 13 9 13 3 12 9 2
2 9 1
12 9 9 13 15 3 0 9 13 11 11 1 2
8 9 9 2 0 9 2 0 9
6 13 3 13 3 0 2
9 3 9 9 13 9 3 12 9 2
4 10 9 13 0
2 3 9
11 3 9 13 9 13 3 3 10 3 9 2
14 15 13 11 2 7 15 15 13 9 3 13 0 9 2
12 9 13 0 7 10 0 9 13 0 9 9 2
5 9 13 9 13 9
10 13 9 13 2 3 13 2 13 9 2
4 9 9 13 2
3 15 13 13
5 11 13 3 0 9
6 3 13 13 10 9 2
2 0 9
11 16 11 13 13 9 2 15 13 0 9 2
2 0 9
7 3 0 13 9 1 9 2
9 11 9 13 9 9 13 0 9 9
5 15 13 15 1 2
10 1 11 9 11 13 13 3 3 9 2
3 9 13 2
9 13 3 15 11 2 16 15 13 2
7 15 13 13 2 11 13 2
9 9 13 13 9 7 9 13 0 2
11 13 2 13 15 13 9 7 3 13 15 2
4 13 16 13 13
12 15 13 9 0 0 11 13 15 9 9 9 2
4 15 13 1 15
10 9 7 9 13 13 13 9 10 0 2
10 0 9 13 0 13 3 9 3 9 2
2 0 9
17 15 13 9 13 12 9 0 0 9 2 15 12 9 1 13 0 2
13 15 13 10 9 13 10 0 9 7 13 9 13 9
15 10 0 9 13 3 0 9 7 13 3 13 3 0 9 2
2 13 13
18 15 13 13 9 0 9 2 16 12 9 9 13 13 1 9 9 9 2
8 9 9 13 0 10 9 9 2
8 3 13 11 9 0 11 9 2
6 15 13 15 0 9 2
6 15 13 15 3 9 2
9 7 3 3 15 13 0 9 13 2
10 11 13 11 9 11 11 9 1 11 2
12 10 3 11 7 11 3 15 3 13 10 9 2
6 11 13 9 10 9 2
12 9 0 13 3 9 2 0 13 10 12 9 2
4 13 3 13 2
9 11 13 0 9 2 15 13 13 2
8 13 13 9 9 13 9 1 2
8 9 9 13 9 7 13 3 9
4 3 13 15 9
10 6 16 13 13 2 13 13 3 9 2
4 15 13 9 1
3 9 13 2
16 15 13 2 16 13 0 9 13 2 16 13 3 9 10 9 2
4 15 13 9 2
6 13 13 13 9 9 2
15 3 9 13 10 0 9 2 3 15 13 13 10 9 3 2
7 3 10 9 13 3 13 2
4 15 13 3 2
14 9 13 13 3 3 15 2 16 0 9 13 13 9 2
3 13 15 3
6 9 13 9 13 9 2
15 13 9 3 9 7 12 9 2 10 9 13 13 3 0 2
16 15 3 13 16 3 13 3 3 11 3 3 15 13 10 0 2
2 9 9
7 9 13 9 9 13 9 2
10 3 11 13 13 9 2 7 3 13 3
7 10 0 9 13 13 3 2
25 11 2 11 2 11 7 10 15 13 3 9 13 9 2 9 2 9 7 3 10 0 9 0 9 2
5 3 15 13 3 2
12 13 12 9 9 3 3 7 15 1 13 9 2
13 13 15 2 3 15 2 3 2 3 2 9 1 2
24 15 13 9 1 9 2 3 13 0 9 0 9 2 15 13 9 9 2 13 3 7 13 3 2
19 9 13 13 9 2 16 15 13 9 2 7 15 1 2 0 9 15 13 2
8 13 13 3 13 0 13 0 2
12 9 13 9 2 16 9 13 13 7 9 13 2
5 15 13 9 1 2
9 10 9 13 13 9 12 9 1 2
9 3 13 13 7 13 0 0 9 2
7 10 12 9 9 13 9 2
13 10 9 13 9 2 10 9 13 0 9 11 9 2
14 15 3 3 13 9 16 11 13 13 9 2 11 13 2
4 13 15 13 2
2 13 3
5 15 15 13 15 2
13 16 9 13 15 3 2 11 13 0 3 3 13 2
11 0 9 13 3 9 9 0 9 13 9 2
8 15 3 3 13 10 9 13 2
12 7 15 13 3 0 9 2 7 13 9 3 2
14 11 12 0 3 12 2 12 13 9 7 12 13 3 2
8 9 13 2 16 15 13 0 2
5 15 13 9 3 2
13 0 9 13 13 9 9 3 16 0 9 9 1 13
11 11 15 3 7 11 13 13 9 13 15 3
8 9 1 13 9 13 10 3 2
3 15 13 9
3 15 13 9
5 13 3 15 13 2
5 15 13 0 15 2
6 0 9 1 13 13 2
4 9 13 13 2
4 15 13 0 9
8 10 9 15 3 13 3 13 2
10 11 9 13 9 9 9 9 12 9 2
6 15 15 13 15 3 13
19 16 13 15 13 2 13 9 13 3 3 2 13 0 9 13 0 0 9 2
7 15 13 0 3 11 1 2
7 13 10 3 9 9 11 2
13 9 13 0 9 15 2 15 13 0 9 3 0 2
15 15 13 3 12 9 9 13 15 2 13 3 13 3 13 2
9 13 2 15 10 9 9 3 13 2
6 9 13 11 9 1 2
4 9 13 0 2
7 11 7 11 13 0 9 2
11 11 11 13 13 0 9 13 0 13 9 2
18 11 13 2 16 9 0 9 13 10 12 9 7 9 2 15 13 9 2
33 15 13 16 15 13 15 3 2 7 15 13 3 0 16 15 13 11 9 2 7 13 15 16 15 13 9 2 7 3 15 13 0 9
9 3 13 15 15 0 9 7 9 2
7 13 3 7 9 13 0 2
7 15 13 13 16 15 13 15
20 3 9 10 9 13 0 7 9 15 13 13 3 0 2 16 0 9 13 13 2
16 15 13 15 2 13 11 9 2 7 15 0 13 3 9 3 2
9 11 13 13 13 11 9 11 1 2
7 11 9 13 3 13 3 2
4 15 15 13 2
12 9 9 9 13 0 2 3 3 12 9 13 2
8 10 0 9 11 13 9 9 2
4 15 13 0 2
22 7 0 13 2 15 15 13 0 7 0 3 11 7 13 9 2 7 15 10 0 13 2
2 0 9
19 11 9 1 13 9 13 13 9 1 7 3 13 13 3 0 9 7 9 2
4 9 13 9 2
2 0 11
10 9 13 11 11 13 0 9 9 1 2
9 9 13 9 1 13 9 7 9 2
14 9 9 13 13 0 0 9 2 7 15 13 9 9 2
17 13 13 9 2 13 9 9 3 2 13 0 9 9 7 13 13 2
6 12 9 13 16 13 2
4 9 13 3 2
6 13 10 9 7 13 2
10 11 13 3 9 1 9 9 0 9 2
14 9 13 9 9 7 15 9 2 13 9 7 13 9 2
7 15 16 13 13 3 9 2
6 9 13 13 13 9 2
5 13 15 0 0 2
3 13 15 2
15 7 9 0 0 9 10 0 9 13 3 10 3 0 13 2
7 13 10 3 13 9 13 2
3 9 13 0
7 10 9 13 13 0 9 2
10 6 2 3 15 13 2 6 6 10 11
2 9 9
7 3 3 7 3 15 13 2
19 3 13 13 2 16 15 13 0 9 7 0 9 2 7 0 9 13 13 2
7 9 13 13 3 3 11 2
8 9 13 11 7 11 11 9 2
5 9 13 13 11 2
6 16 13 2 13 9 2
12 0 9 13 13 3 13 3 0 9 16 3 2
8 9 11 13 13 3 0 9 2
27 11 13 9 7 10 9 15 13 2 16 9 13 15 3 10 9 2 16 16 9 13 13 2 3 9 3 2
15 11 13 3 10 9 2 16 12 9 9 13 13 10 0 2
3 15 13 2
13 13 3 9 2 16 0 9 13 13 3 11 9 2
5 13 15 13 16 2
17 13 9 9 13 3 0 3 9 9 2 3 13 0 0 9 9 2
11 11 13 13 3 2 16 15 13 9 9 2
7 9 13 9 8 7 9 9
5 11 13 9 11 2
25 13 13 3 13 9 10 0 9 9 15 13 3 9 7 3 13 3 9 0 9 7 10 0 9 2
8 3 13 2 16 3 13 9 9
4 9 13 9 9
7 9 9 7 9 1 13 2
12 15 13 3 0 15 2 16 13 13 3 9 2
4 3 15 13 9
4 6 10 9 2
2 0 0
4 11 9 12 11
4 13 12 9 2
12 1 9 2 13 9 3 9 2 9 7 9 2
3 11 13 13
10 15 13 13 9 3 9 2 3 9 2
14 3 13 3 10 9 2 13 13 11 9 9 11 11 2
3 13 9 9
6 16 15 13 3 13 2
13 15 13 15 9 3 13 2 16 13 9 0 9 2
2 13 3
8 0 9 1 15 3 13 9 2
9 15 13 13 9 0 9 0 9 2
2 6 2
8 9 13 3 0 9 7 9 2
8 13 0 2 16 13 3 9 2
10 11 13 9 13 7 12 9 13 13 2
5 15 13 9 9 2
6 9 9 3 7 3 2
6 3 13 3 0 9 2
11 9 13 9 7 10 9 0 9 11 1 2
15 0 9 13 11 0 2 10 9 3 13 9 0 12 9 2
12 15 13 9 9 9 2 15 13 13 9 1 2
8 9 13 9 0 15 13 9 2
8 11 9 13 3 9 1 0 2
6 11 11 13 9 12 2
13 3 9 13 13 9 7 10 9 9 9 12 1 2
6 0 9 13 0 9 2
15 11 13 3 9 1 10 9 9 2 15 13 13 13 9 2
7 11 13 3 13 11 9 2
12 11 9 13 9 13 13 10 9 10 0 9 2
5 15 13 2 13 3
7 11 3 13 9 13 9 2
4 13 3 9 2
11 9 9 9 13 13 3 15 3 13 9 2
4 13 3 0 2
3 8 7 9
17 11 9 13 3 15 2 16 11 13 13 13 11 9 1 13 9 2
10 13 10 9 0 9 2 1 0 9 2
8 16 13 9 2 3 9 13 2
12 11 13 9 7 11 15 1 13 9 9 3 2
19 9 9 13 9 3 3 12 9 2 16 3 15 13 11 9 11 12 9 2
10 9 13 3 2 16 13 8 7 9 2
8 9 9 9 13 13 0 9 2
5 12 9 13 13 2
9 9 13 3 0 7 13 9 9 2
22 11 9 9 13 13 11 9 13 12 9 11 2 16 9 13 10 9 13 3 12 9 2
9 10 9 15 3 13 2 11 13 2
13 9 13 9 9 9 13 3 12 9 0 7 0 2
13 9 2 13 3 9 2 3 15 13 15 3 9 2
9 3 13 16 13 3 3 13 13 2
9 15 13 9 16 9 13 9 3 2
5 13 15 15 13 2
8 9 15 13 9 11 9 12 2
7 11 9 9 13 3 0 2
7 3 0 9 13 13 9 2
11 13 15 10 9 13 2 16 15 15 13 2
6 0 9 11 13 0 2
4 13 15 0 2
11 9 13 3 0 13 15 3 13 13 9 2
3 10 9 16
12 3 9 13 13 9 2 3 16 15 13 13 2
8 13 13 2 3 9 11 13 2
10 13 3 3 9 2 3 0 9 13 2
6 0 9 11 11 0 9
19 9 9 13 3 0 9 13 9 7 13 9 9 16 9 0 9 13 9 2
7 9 13 13 11 1 11 2
12 0 9 1 13 13 9 10 13 13 9 1 2
6 11 13 13 15 13 2
2 13 13
3 13 9 2
9 15 13 13 10 9 2 13 13 2
4 9 13 9 2
7 11 9 13 13 11 0 2
20 13 9 13 9 11 3 0 13 9 2 15 1 9 9 13 11 0 9 9 2
9 9 13 3 13 0 13 9 9 2
13 11 1 9 13 9 2 15 13 0 9 16 9 2
9 3 8 7 9 13 9 13 3 2
8 15 13 9 7 13 3 3 2
11 8 13 13 2 16 11 9 13 0 3 2
8 9 13 13 3 16 3 13 13
14 9 13 3 15 2 16 9 3 13 9 13 9 3 2
5 3 3 9 0 9
2 13 9
5 3 15 3 9 2
3 13 9 1
14 15 13 0 9 2 7 3 10 0 9 13 13 9 2
5 3 0 15 13 2
7 9 13 9 1 9 1 2
17 10 9 7 10 9 13 13 10 9 2 16 13 13 13 15 3 2
11 3 16 13 10 9 13 0 2 3 13 2
7 11 9 13 9 1 9 2
3 13 9 1
5 15 15 13 9 2
6 9 13 13 9 1 2
10 9 13 3 3 2 16 13 9 13 2
4 9 13 0 9
10 15 13 15 9 16 9 13 0 9 2
4 15 13 9 2
8 0 9 1 9 13 3 12 9
8 10 9 9 13 9 9 9 2
3 9 9 9
17 3 9 13 3 3 0 7 3 13 7 13 9 2 0 7 9 2
10 16 15 13 2 13 13 13 15 9 2
3 9 15 13
17 11 13 16 15 13 13 9 9 7 12 9 9 16 9 13 3 2
5 9 2 9 7 9
11 13 2 3 3 13 0 9 7 10 9 2
5 13 13 0 9 2
3 9 13 13
15 6 15 16 11 13 2 3 15 13 13 9 3 0 9 2
2 9 13
10 7 15 15 13 13 10 0 0 9 2
5 9 13 3 9 2
8 9 13 3 3 16 13 13 2
11 13 0 16 12 13 7 16 12 13 13 2
5 9 13 10 9 2
5 15 3 9 13 2
11 3 16 11 11 13 10 0 9 9 9 2
4 15 13 9 1
7 9 9 13 9 9 9 2
2 9 9
10 9 13 13 3 12 9 0 12 1 2
5 11 13 13 9 2
6 13 13 9 2 13 13
13 9 13 9 1 12 9 2 3 3 12 9 9 2
8 9 13 13 10 9 7 13 2
11 0 13 9 7 9 13 9 13 9 9 2
9 3 15 13 12 9 1 12 9 2
13 6 2 16 3 3 13 2 3 3 13 15 13 2
6 13 9 15 15 1 2
5 13 9 13 9 2
11 7 10 9 13 9 13 9 1 0 9 2
14 15 9 13 13 13 2 13 11 7 11 13 11 9 2
13 13 15 13 13 13 9 9 3 7 13 15 9 2
10 9 9 13 7 13 12 9 9 13 2
14 16 15 13 9 2 3 9 13 3 0 9 0 9 2
14 13 13 2 16 13 13 9 7 9 0 16 15 13 2
2 9 13
14 3 0 9 2 16 15 13 0 2 11 3 13 0 13
7 9 1 9 13 3 3 2
10 9 2 15 9 13 15 0 7 0 13
13 9 3 9 13 13 3 3 2 7 0 13 13 2
6 15 13 9 7 9 2
15 9 13 9 13 9 9 9 9 2 3 13 10 0 9 2
18 9 13 9 13 3 9 7 13 0 2 16 9 13 0 9 9 1 2
14 9 11 13 3 13 2 7 9 15 13 3 7 3 2
3 13 15 3
3 13 13 2
4 13 13 9 2
6 15 13 9 13 9 2
11 13 3 13 2 16 13 3 13 15 13 2
13 13 3 13 3 2 16 9 13 9 10 9 0 9
17 11 9 9 13 9 13 3 3 3 0 12 9 9 2 12 2 2
13 9 13 9 2 15 9 0 9 7 9 13 9 2
7 9 13 10 3 0 9 2
14 10 2 0 2 9 13 13 3 0 7 13 3 13 2
9 9 13 0 2 7 13 3 0 2
15 15 13 11 9 3 3 13 16 13 10 9 10 0 9 2
5 13 13 10 9 2
9 9 7 9 13 0 9 9 13 2
8 9 1 9 11 13 13 9 2
4 11 13 11 2
5 9 13 3 9 2
10 3 13 9 9 13 3 12 12 9 2
16 11 13 3 0 0 2 2 7 10 9 13 9 7 13 9 2
7 13 0 2 16 9 13 2
10 13 13 2 16 9 7 9 13 15 2
4 11 11 11 9
12 13 11 11 7 9 13 10 9 13 9 9 2
16 13 9 2 16 9 13 10 0 9 9 13 9 9 11 11 2
10 11 13 13 9 15 13 15 3 3 2
30 11 13 13 9 3 2 7 16 13 15 13 13 10 9 15 2 13 15 15 13 2 15 13 13 3 3 3 3 3 2
11 9 9 13 11 9 12 9 13 9 9 2
3 15 13 2
8 2 13 11 7 13 9 2 2
10 13 3 13 9 2 15 13 0 15 2
8 9 13 9 16 13 10 9 2
11 13 9 13 2 16 11 13 3 0 9 2
7 15 13 0 0 0 9 2
8 0 16 3 0 9 13 13 2
8 15 13 13 10 0 11 9 2
13 11 13 13 13 9 1 9 2 3 13 15 9 2
7 15 13 13 15 13 9 2
18 9 13 13 3 9 12 2 3 10 9 9 9 7 9 1 13 0 2
3 13 7 13
6 0 9 13 3 3 2
13 16 10 9 13 3 3 2 15 13 3 3 11 1
12 3 9 16 9 13 9 2 15 13 13 9 12
12 15 15 2 11 13 11 3 9 7 0 9 2
6 13 9 7 13 9 2
2 9 9
5 13 9 13 15 2
9 15 13 13 15 2 7 13 9 2
19 11 11 9 13 0 0 9 9 2 9 7 9 9 7 0 7 0 9 2
2 13 13
2 13 9
16 12 9 2 12 9 7 9 1 15 13 7 13 9 13 9 11
9 9 9 13 9 7 9 1 0 2
11 9 13 15 3 3 3 16 12 9 1 2
6 15 13 3 3 13 2
9 16 13 13 9 3 2 13 13 2
11 0 7 0 13 11 9 3 3 13 15 2
9 3 13 13 0 9 13 13 9 2
4 9 13 0 2
4 11 0 0 9
5 15 13 9 9 2
13 9 9 13 0 2 16 13 9 9 12 3 9 2
34 10 0 7 0 9 15 9 9 2 15 3 13 3 15 2 13 10 10 9 13 3 11 2 11 7 11 2 13 3 3 13 9 3 2
4 13 13 9 2
21 11 13 7 13 9 7 15 9 13 0 9 13 13 0 9 9 9 9 0 9 2
6 11 13 13 9 3 9
11 15 13 9 13 3 2 16 0 9 13 2
15 13 11 2 11 7 11 1 9 15 2 16 11 13 9 2
13 13 13 10 9 2 15 15 13 15 0 7 0 2
2 0 9
5 13 9 7 13 2
7 13 3 3 0 15 13 2
12 11 13 0 9 2 16 9 13 13 13 3 2
14 15 13 3 0 9 2 3 16 15 13 3 0 9 2
10 9 9 13 13 15 13 13 15 3 2
21 13 3 13 9 2 16 9 13 9 3 9 7 9 7 13 9 0 9 7 9 2
8 3 13 13 9 15 1 13 2
6 13 13 2 15 15 13
20 11 13 2 16 13 11 10 9 13 7 13 3 3 0 2 16 15 13 3 2
14 9 9 9 13 13 9 1 3 9 9 2 13 9 2
6 9 9 13 12 9 2
7 9 13 13 3 9 13 2
10 13 3 0 2 16 9 13 0 9 2
9 13 13 3 0 9 1 10 2 9
2 0 9
12 9 13 12 9 7 15 13 13 3 12 9 2
10 3 3 9 13 13 9 9 2 7 2
3 0 9 2
11 15 13 9 2 13 9 7 13 3 15 2
7 13 0 2 16 13 3 2
13 12 9 13 0 11 11 7 12 9 11 11 11 2
10 11 1 9 0 9 9 1 13 0 2
8 3 3 9 3 10 9 9 2
7 15 13 15 7 13 3 2
14 9 13 13 15 2 16 10 9 13 13 3 13 9 2
7 15 13 0 13 13 3 2
6 9 9 9 3 3 3
5 9 13 3 3 2
6 13 3 13 7 13 2
8 11 13 13 9 13 9 9 2
9 3 9 11 9 3 13 3 11 2
5 10 9 13 0 2
2 9 9
7 15 13 0 9 7 13 2
6 13 3 0 9 1 2
6 11 15 15 13 13 2
10 0 9 15 13 13 13 13 2 16 2
12 13 13 9 2 16 11 15 13 13 0 9 2
10 6 16 13 3 12 9 3 11 13 2
3 10 9 1
3 3 0 0
22 9 13 13 9 9 9 2 7 11 13 2 16 10 12 13 0 9 3 9 7 9 2
5 10 9 13 15 2
9 13 9 3 9 7 13 3 3 2
6 15 13 13 3 3 2
19 15 9 13 2 15 13 3 7 3 2 16 3 9 13 9 15 10 9 2
4 15 13 13 2
9 15 13 2 3 13 3 0 9 2
16 15 13 3 3 12 2 13 9 7 9 7 13 9 13 9 2
13 11 9 9 9 13 2 9 13 3 7 9 13 2
10 11 13 11 9 7 13 10 9 3 2
6 13 15 9 7 9 2
10 13 9 2 3 11 9 9 3 13 2
2 0 0
5 13 15 13 9 2
11 12 9 1 13 15 13 15 13 11 9 2
4 13 9 9 2
7 15 13 3 2 0 3 2
14 13 13 9 9 2 3 16 15 9 13 13 9 0 2
17 11 9 11 13 13 0 9 2 16 11 13 16 15 3 3 13 2
8 9 15 13 11 3 13 9 2
8 13 9 9 10 9 1 3 9
12 8 8 9 13 0 7 0 2 15 13 13 2
7 0 16 13 3 13 3 2
5 9 13 3 13 2
11 3 9 13 0 2 16 3 3 15 13 2
12 10 10 0 9 9 9 7 9 13 3 9 2
5 13 3 15 13 2
13 15 15 3 13 2 16 9 13 3 7 13 3 2
21 9 13 3 13 3 13 7 3 13 2 3 13 9 13 7 13 7 13 0 9 2
4 13 13 9 2
11 15 13 3 16 13 0 9 2 9 13 2
11 11 13 9 3 7 13 3 9 9 1 2
7 9 13 11 13 3 9 2
12 13 9 3 13 10 9 10 9 13 7 13 2
7 15 15 13 13 9 13 2
4 9 13 0 13
5 3 10 9 13 2
4 15 13 3 13
8 9 13 13 2 3 13 15 2
18 16 10 9 9 13 12 9 2 15 13 13 3 2 16 15 13 13 9
6 15 3 13 0 9 2
6 10 9 13 0 9 2
6 3 13 13 3 3 2
6 3 15 13 3 3 2
7 9 13 13 15 16 10 15
4 13 0 9 9
5 13 10 12 9 2
6 10 9 13 11 0 2
10 10 9 1 13 13 13 9 9 13 2
20 9 13 13 7 16 13 0 9 2 3 3 15 13 12 9 13 9 3 3 2
12 11 13 0 9 2 13 3 0 3 16 9 2
11 13 13 15 0 9 9 2 9 7 9 2
2 9 9
12 9 11 7 9 11 13 13 9 1 13 9 2
19 11 9 2 9 7 9 9 13 3 0 0 2 3 16 15 13 0 13 2
6 13 13 13 10 9 2
5 11 13 10 0 2
21 16 3 9 7 15 13 13 16 7 10 9 3 16 9 9 3 13 15 10 9 2
11 9 1 11 13 13 13 9 0 9 9 2
2 15 1
3 13 13 2
2 9 9
18 7 16 10 10 9 13 9 3 3 15 13 3 13 16 15 13 13 2
5 9 13 13 9 2
4 15 13 9 2
8 9 13 9 9 1 13 3 2
11 15 13 13 0 9 16 13 0 9 15 13
8 13 10 11 3 13 13 15 3
10 15 13 9 2 15 13 3 3 9 2
4 9 13 12 9
4 13 15 9 2
5 0 13 9 9 2
12 9 13 0 7 0 2 3 13 9 0 9 2
2 13 15
3 9 13 9
5 15 13 3 0 2
2 13 0
14 3 13 9 13 9 2 10 9 13 9 7 9 9 2
13 9 13 3 9 15 2 13 11 9 10 9 9 2
16 16 9 13 9 1 2 9 13 13 13 2 7 9 13 9 2
6 9 13 3 13 0 2
8 9 13 13 9 0 0 9 2
5 15 13 3 3 9
2 7 15
7 13 2 16 15 13 9 2
4 9 13 9 2
8 0 9 9 13 3 2 13 2
5 9 13 13 9 9
8 12 0 9 11 13 9 9 2
5 13 9 12 9 2
6 15 13 2 0 9 2
6 9 13 7 13 3 2
7 0 13 0 9 9 9 2
3 13 13 9
4 15 13 9 2
2 13 3
5 15 9 9 13 2
4 10 0 0 9
4 3 13 9 2
8 13 13 13 15 0 9 3 0
6 13 13 10 9 9 2
9 13 13 2 3 3 15 13 9 2
7 0 9 13 0 9 1 2
10 9 13 0 2 16 15 13 13 15 2
12 10 3 9 7 9 7 9 13 3 9 3 2
5 13 11 13 11 2
19 3 15 3 13 0 9 3 2 15 13 0 9 7 9 16 9 13 9 2
11 13 13 0 2 7 13 0 7 0 9 2
4 13 15 13 2
9 11 11 13 9 13 0 0 9 2
8 9 13 10 9 9 9 11 2
8 9 13 9 2 9 9 13 2
6 13 9 13 3 3 2
9 6 6 2 13 2 16 13 15 2
9 3 9 13 9 7 15 3 9 2
10 9 13 13 12 7 12 16 13 9 2
8 3 13 15 16 13 9 13 2
12 3 15 13 9 7 0 9 3 13 16 15 2
12 0 9 2 11 12 2 13 9 9 13 9 2
12 15 13 9 9 7 9 11 9 0 9 9 2
11 13 9 3 2 7 6 15 10 9 13 2
7 3 13 9 0 7 0 2
20 3 16 3 3 13 3 10 11 9 3 3 3 13 3 15 15 3 13 0 2
6 11 13 9 9 11 2
11 7 8 16 9 13 9 13 0 9 9 2
20 15 13 13 13 3 9 2 13 9 2 9 9 13 13 9 15 13 13 9 2
6 13 3 3 0 9 2
16 9 13 13 10 0 9 2 3 0 9 13 13 3 9 3 2
13 15 15 3 13 2 16 9 13 3 7 13 3 2
9 0 9 13 13 0 9 7 9 2
4 15 9 13 2
10 13 9 2 13 15 13 2 7 13 2
14 16 0 11 13 13 9 0 2 9 13 0 9 9 2
6 13 15 15 2 9 2
8 15 1 9 13 9 9 9 2
7 16 13 9 2 13 3 13
5 13 13 13 13 15
3 2 6 2
18 13 13 15 15 15 13 2 9 0 9 13 3 2 7 15 13 13 2
12 7 9 13 13 9 2 3 9 3 3 13 2
2 10 9
7 9 9 7 9 13 15 2
2 9 15
5 15 13 3 0 2
3 9 13 9
4 13 15 13 2
7 15 13 9 7 13 9 2
4 2 13 15 2
10 9 9 13 9 13 13 15 0 9 2
12 16 11 13 3 9 3 15 13 3 0 9 2
10 9 13 3 15 8 2 3 3 9 2
9 13 3 0 8 2 8 7 9 2
15 9 13 9 13 0 2 3 3 9 7 3 3 16 9 2
17 0 9 9 13 13 9 2 15 13 9 1 7 13 9 9 9 2
10 3 3 7 7 9 13 11 13 9 2
11 13 9 7 9 2 13 9 2 13 9 2
15 13 13 13 9 3 2 7 15 16 13 2 16 13 3 2
10 11 13 13 13 0 0 7 0 9 2
3 6 15 15
5 13 9 0 11 2
5 9 13 11 9 11
6 3 13 9 7 9 2
11 15 13 16 15 13 9 13 16 9 3 2
10 0 9 13 0 11 9 13 0 9 13
9 13 15 3 12 9 10 11 3 2
12 10 0 9 13 0 7 0 16 9 7 9 2
2 13 3
3 3 0 9
12 9 9 13 12 12 9 13 3 12 12 9 2
17 15 13 13 12 1 9 2 13 2 7 13 3 9 13 3 15 2
7 9 13 3 9 9 9 2
8 9 13 9 7 15 0 9 2
6 9 9 9 13 0 2
8 9 13 2 15 15 13 13 2
5 7 0 7 0 9
6 9 13 0 0 9 2
8 3 15 13 15 3 10 9 2
12 1 13 9 3 13 3 9 3 9 7 9 2
4 9 13 3 0
3 13 15 3
3 11 9 11
9 13 10 9 9 1 13 0 9 2
8 3 9 13 9 13 9 9 2
21 7 15 13 3 15 2 16 16 15 13 10 9 9 2 3 15 13 13 10 9 2
26 3 16 15 13 0 3 13 2 13 3 3 2 7 3 13 2 6 7 3 13 3 16 15 13 11 2
8 9 13 9 15 9 13 9 2
7 15 13 9 13 3 9 2
3 13 13 2
12 9 13 0 9 11 11 7 15 13 11 11 2
4 6 0 9 2
10 0 9 9 11 13 13 11 9 9 2
11 16 9 13 9 2 3 3 13 13 3 2
2 12 9
12 13 13 3 0 15 2 16 13 11 9 13 2
5 9 9 7 9 9
10 16 0 13 3 9 2 13 9 15 2
2 0 9
3 13 13 15
9 9 9 13 13 9 7 0 9 2
3 0 0 9
15 9 13 7 0 12 9 2 3 2 3 7 9 9 1 2
14 7 13 2 16 13 3 0 2 16 9 13 10 9 2
4 6 15 15 2
15 3 0 7 0 9 13 13 2 3 3 15 13 13 13 2
12 15 13 16 3 3 13 13 15 13 3 3 2
3 0 9 11
20 15 13 3 9 9 9 12 9 1 7 15 13 3 0 9 11 9 9 9 2
4 13 10 9 2
12 10 9 13 9 9 9 13 3 15 1 13 2
9 7 3 3 0 9 9 12 13 2
13 1 0 11 7 9 9 13 9 13 0 11 11 2
3 9 13 15
2 13 13
4 13 9 0 11
6 15 13 7 9 13 2
10 3 11 9 1 13 9 13 0 9 2
9 11 13 9 9 2 7 0 9 2
8 9 13 9 1 3 12 9 2
2 3 9
7 15 13 13 2 13 9 2
13 13 3 3 3 2 16 15 13 0 9 0 9 2
8 9 11 13 3 0 16 11 2
9 11 0 9 13 9 0 7 0 2
12 16 9 13 2 3 9 13 3 12 12 9 2
4 13 10 9 2
6 13 3 13 0 13 2
7 15 13 11 9 0 9 2
3 9 9 3
5 6 13 0 9 2
2 9 1
18 9 9 13 2 16 13 3 9 1 3 3 0 9 7 9 2 9 2
6 15 13 13 9 13 2
7 3 3 16 3 13 15 2
9 15 13 10 0 9 2 9 13 2
4 9 13 15 2
2 11 9
10 9 13 13 3 9 2 7 3 15 2
2 13 0
14 15 13 13 9 2 15 13 13 9 3 2 13 9 2
6 13 0 9 11 11 2
9 16 9 13 13 0 2 13 15 2
3 16 13 15
6 13 9 7 13 9 2
13 15 13 13 0 0 9 2 16 13 13 9 1 2
8 11 1 13 13 9 0 3 2
9 9 13 9 13 0 9 10 9 2
6 13 9 0 9 1 2
7 15 13 13 0 0 9 2
11 6 3 3 0 16 9 3 13 15 0 2
12 11 13 13 9 9 10 3 10 0 0 9 2
9 3 0 9 3 13 13 3 9 2
7 15 13 13 15 9 1 2
5 15 13 13 13 3
10 13 3 13 9 2 15 13 0 15 2
10 3 9 13 10 9 11 3 0 9 2
13 10 0 13 15 2 16 9 9 9 13 9 9 2
2 0 11
10 13 13 9 2 16 13 9 13 0 2
5 11 13 13 9 2
12 13 10 9 9 7 9 7 13 10 9 9 2
22 11 13 13 15 2 16 10 0 13 11 9 12 12 7 16 9 9 13 13 12 9 2
16 7 13 13 9 9 1 2 3 16 13 3 0 1 3 3 2
11 3 9 11 7 3 11 8 0 9 11 2
7 11 9 13 10 12 9 2
4 9 9 13 3
3 2 15 3
6 13 3 13 3 0 2
9 9 11 13 9 3 9 7 9 2
15 3 13 16 13 3 10 9 16 9 2 7 3 13 3 2
10 13 3 2 16 9 13 3 9 9 2
13 9 3 13 2 7 13 3 3 3 16 10 15 2
13 9 13 13 3 9 2 7 9 15 13 13 13 2
15 9 9 13 3 13 9 2 3 9 13 13 10 9 9 2
3 9 13 9
8 10 0 9 2 9 13 11 2
21 9 13 13 3 2 16 9 13 13 13 9 0 9 1 7 16 15 13 13 9 2
16 3 10 9 7 9 13 0 9 16 15 15 2 3 9 1 2
9 9 13 3 13 0 9 11 9 2
6 9 1 3 13 9 11
15 13 9 9 13 15 13 13 3 13 15 15 15 13 13 2
4 13 15 3 2
19 10 9 15 13 0 7 3 3 3 13 9 2 10 9 13 3 13 13 2
18 3 12 11 13 12 9 9 2 0 9 3 12 2 9 3 12 9 2
9 9 11 9 13 3 1 15 9 2
7 3 12 9 13 3 3 2
7 2 10 9 13 0 2 2
5 9 13 0 0 2
14 13 9 2 16 13 3 9 2 15 13 3 9 2 2
3 3 13 9
20 9 13 13 0 2 16 9 3 13 2 7 3 16 9 9 13 13 15 0 2
13 9 13 3 9 0 9 9 13 15 3 0 9 2
3 10 9 2
12 9 13 3 9 2 10 9 13 11 7 9 2
7 15 13 13 9 3 0 2
6 7 3 15 13 9 2
5 2 15 13 9 2
5 11 9 13 0 9
3 9 0 9
8 0 9 13 13 3 3 3 2
11 15 13 0 16 3 13 13 9 13 9 2
3 15 13 2
10 13 13 13 9 2 7 9 13 9 2
9 9 7 9 9 13 0 9 9 2
14 3 13 13 3 0 13 13 15 9 13 9 13 13 2
2 3 3
16 13 13 3 0 9 2 7 15 13 2 16 9 13 3 15 2
12 13 9 13 3 12 9 2 15 13 3 9 2
6 0 9 9 13 13 2
6 3 0 13 15 13 2
2 3 13
8 3 13 13 13 12 0 9 2
7 13 15 13 10 9 9 2
12 13 3 0 15 1 2 13 9 13 13 9 2
12 16 12 9 1 13 13 9 2 13 9 0 2
8 13 3 3 0 13 10 0 2
2 3 3
8 9 13 13 10 9 7 9 2
7 13 9 9 8 7 9 2
42 3 2 15 13 3 15 1 15 13 0 0 9 7 15 13 3 3 9 3 7 3 10 9 13 15 16 15 13 3 13 2 16 15 13 2 13 13 13 15 2 3 3
8 13 15 3 0 8 3 15 2
13 7 3 3 15 13 13 0 7 0 2 3 0 2
9 3 15 13 13 15 3 9 1 2
10 11 1 12 9 13 13 15 9 9 2
11 16 13 3 0 2 3 13 13 3 13 2
5 13 15 9 1 2
5 15 13 9 3 2
5 2 13 3 9 2
4 15 13 13 13
6 13 11 13 3 9 2
