1929 17
17 10 9 15 13 7 13 9 7 1 10 9 7 1 10 0 9 2
27 3 3 13 0 9 2 10 15 1 15 13 9 1 10 0 9 7 0 9 1 0 9 2 9 7 9 2
37 10 0 9 13 10 9 3 3 2 13 14 13 3 1 10 9 9 7 3 0 9 2 3 13 10 0 9 1 9 10 9 7 10 9 15 13 2
17 13 7 15 10 9 14 13 9 7 1 9 9 9 1 10 9 2
3 2 9 2
15 13 0 9 1 10 9 9 7 10 9 13 10 9 15 2
38 15 1 9 1 10 9 1 10 0 9 15 13 13 14 13 7 13 1 10 0 9 10 9 9 7 10 0 0 9 1 9 10 9 13 10 12 9 2
23 15 13 10 0 0 9 7 13 1 0 9 10 9 14 14 13 3 3 10 9 10 0 2
83 1 9 2 10 9 13 3 10 0 9 0 9 1 0 9 2 7 1 10 9 1 9 10 9 1 9 1 10 0 9 2 3 10 12 10 0 9 13 14 13 1 3 0 9 9 2 9 10 9 2 9 7 9 1 0 9 2 10 15 13 14 13 10 0 9 7 14 13 1 15 9 9 7 9 2 3 10 9 7 10 0 9 2
37 14 13 14 13 13 9 1 10 0 9 15 3 1 10 0 9 2 10 15 2 3 2 3 15 0 9 10 2 2 14 13 14 13 3 0 9 2
25 10 9 9 13 1 10 9 10 9 1 10 15 10 9 13 10 9 1 9 15 2 1 9 9 2
21 10 9 10 15 13 10 9 13 7 14 13 0 7 14 13 10 0 9 10 9 2
46 1 10 9 15 10 9 9 10 9 13 14 13 10 9 1 9 10 9 9 7 9 2 10 15 13 9 2 1 10 0 9 15 9 14 13 10 0 2 10 0 7 7 10 0 9 2
10 10 0 15 9 13 10 9 0 9 2
40 10 0 9 10 9 7 10 0 15 9 14 13 9 1 0 9 2 13 3 9 7 1 15 9 14 13 9 15 14 13 14 13 1 3 9 7 9 0 9 2
35 10 9 13 1 9 10 0 9 9 7 9 2 2 2 1 10 0 9 2 10 9 2 10 9 2 10 9 2 10 3 9 7 10 9 2
70 1 10 9 15 10 0 9 10 9 13 2 13 14 13 2 13 0 9 10 9 3 1 0 0 9 15 13 2 13 3 10 9 1 15 0 9 2 10 9 15 13 10 9 7 2 9 14 3 0 2 10 0 9 9 10 0 9 1 10 9 9 1 15 12 1 10 12 9 9 2
41 13 1 10 9 9 1 0 0 9 2 1 9 10 0 9 1 9 9 2 1 9 1 10 15 13 0 9 9 7 3 7 9 1 0 2 1 10 9 0 9 2
9 13 7 15 13 10 3 0 9 2
11 10 9 14 13 9 9 1 0 10 9 2
13 10 9 10 9 13 1 10 9 7 13 1 9 2
25 10 9 13 1 0 0 9 10 9 1 10 15 10 0 9 13 1 9 10 0 0 1 0 9 2
47 10 9 9 2 9 10 1 9 9 1 10 0 9 2 13 7 2 3 10 9 7 10 0 9 13 9 9 1 9 2 14 13 14 13 0 7 0 9 1 10 9 10 9 1 9 2 2
26 1 9 9 2 1 9 9 1 9 10 9 9 13 10 9 1 14 13 10 9 14 13 10 9 15 2
25 0 9 13 7 2 10 9 13 0 9 2 9 9 2 9 7 9 1 10 0 9 1 15 13 2
20 10 9 9 13 10 9 10 9 9 2 7 10 9 9 13 14 13 10 9 2
16 10 9 15 1 9 9 1 10 0 9 13 1 10 0 9 2
18 7 13 14 13 1 10 3 0 9 2 1 15 10 9 13 12 9 2
19 3 3 13 0 7 14 13 13 10 9 3 3 3 15 13 15 10 9 2
17 10 9 15 9 14 13 0 9 9 1 9 2 13 10 0 9 2
26 15 13 10 9 15 13 1 1 9 9 2 7 13 14 13 15 10 0 10 0 9 15 13 1 15 2
2 12 2
67 3 2 0 9 1 0 9 13 14 13 10 0 9 2 15 13 10 2 9 9 2 1 10 9 10 9 2 1 10 15 13 9 1 10 0 9 2 1 10 9 10 9 10 9 10 15 2 15 1 9 1 10 0 9 2 13 14 13 1 10 0 9 10 9 10 9 2
13 2 2 0 9 13 0 9 1 0 9 10 9 2
37 7 3 1 15 9 2 9 1 10 9 13 9 3 1 10 15 10 9 10 9 13 3 14 13 9 2 7 14 3 14 13 10 9 10 3 0 2
31 1 3 13 3 0 9 9 1 9 10 0 9 7 7 15 9 7 10 9 10 9 13 1 0 9 10 9 7 10 9 2
44 1 9 2 10 0 9 13 9 1 10 9 10 9 2 13 15 2 0 12 9 2 2 7 13 7 2 10 2 13 3 14 13 14 3 9 7 7 9 1 10 0 9 2 2
34 10 0 9 2 2 2 7 0 9 2 3 7 10 0 0 9 9 13 1 0 9 15 0 0 9 7 10 0 0 9 13 0 9 2
17 14 13 3 1 9 15 14 13 3 9 1 0 9 9 10 9 2
23 3 13 0 10 9 15 7 13 14 13 3 0 0 9 9 1 0 9 1 3 12 9 2
27 10 9 13 14 13 10 0 9 15 1 10 9 3 12 9 1 10 9 10 9 1 10 9 15 10 9 2
48 14 13 10 9 7 2 15 7 7 13 10 9 15 13 10 9 1 10 0 7 0 9 2 10 0 9 13 14 15 13 7 13 7 10 9 13 10 0 7 0 0 9 7 9 1 0 9 2
8 12 0 9 13 13 1 9 2
22 1 10 0 9 10 9 13 10 0 9 10 9 1 12 9 10 9 7 1 10 9 2
47 10 9 10 0 9 15 13 3 1 10 9 10 9 2 10 0 9 1 10 12 9 10 12 9 2 3 7 10 9 2 10 15 13 3 1 9 10 9 13 10 9 7 9 10 0 9 2
23 3 2 3 12 9 9 13 13 1 9 10 9 1 9 10 9 2 13 10 12 9 9 2
2 12 2
21 10 2 2 10 2 7 10 2 13 13 10 9 9 1 10 13 9 9 7 9 2
16 0 13 1 9 10 9 10 9 2 7 13 13 7 10 9 2
4 2 2 9 2
35 10 9 13 10 9 15 13 3 1 0 9 10 0 9 13 1 10 0 9 1 10 9 9 7 9 2 10 15 13 2 3 10 9 2 2
50 1 9 10 9 10 12 9 10 9 9 13 1 12 10 9 10 9 2 10 0 9 9 2 9 0 2 7 7 10 3 0 9 2 10 15 1 10 0 9 15 13 2 1 9 2 13 1 10 9 2
18 13 14 14 13 10 9 1 10 0 1 0 1 10 0 7 10 0 2
31 12 1 10 3 0 9 10 9 13 10 9 10 9 10 9 15 13 13 1 10 0 9 15 3 13 1 0 0 10 9 2
27 10 9 13 1 10 9 10 9 2 15 13 10 9 7 13 10 9 10 9 15 15 13 3 10 0 9 2
41 7 2 10 9 13 13 14 13 1 0 9 10 9 7 10 0 13 14 13 1 10 0 0 9 2 0 10 0 9 0 9 2 1 10 9 10 9 9 10 0 2
55 13 0 7 15 9 10 9 14 13 1 9 14 13 7 14 13 10 9 3 1 15 10 0 9 2 10 15 2 1 0 9 2 14 13 10 9 15 7 13 3 2 7 10 0 9 10 15 13 10 0 9 10 9 9 2
52 10 9 13 3 7 10 9 10 0 9 3 1 10 9 13 14 13 1 9 10 9 9 1 10 0 9 7 10 9 10 0 9 7 10 0 9 2 10 0 0 9 7 10 9 10 0 9 10 9 10 9 2
11 10 12 9 13 1 9 12 1 10 9 2
4 15 13 0 2
36 3 1 9 2 3 10 9 13 12 9 2 7 3 13 7 13 12 9 2 1 10 9 12 9 2 10 15 13 10 0 9 10 2 10 9 2
37 10 9 10 9 10 0 9 13 1 10 0 0 9 1 10 9 7 10 9 1 10 9 10 9 9 1 10 2 9 9 2 15 13 1 9 9 2
29 3 2 10 9 9 13 13 1 12 9 9 7 13 1 10 9 2 10 15 13 14 15 13 1 10 9 0 9 2
50 10 9 10 9 13 7 13 3 1 10 9 2 3 3 10 0 14 13 3 0 2 7 10 0 7 0 9 10 9 13 2 1 0 0 9 14 13 1 10 9 7 14 13 1 10 0 9 1 9 2
18 10 9 13 0 9 1 0 9 2 1 9 7 12 9 1 10 9 2
59 13 1 10 9 10 2 9 2 7 13 0 7 0 9 1 9 15 3 1 10 9 2 10 9 7 10 9 2 12 9 2 9 3 10 9 10 9 2 15 14 13 13 1 9 0 7 0 9 10 15 13 7 10 15 7 15 15 13 2
17 10 12 9 2 15 13 10 0 9 2 13 10 15 3 0 9 2
78 1 10 9 15 2 10 9 14 13 14 13 3 3 7 0 9 2 3 7 0 9 2 7 9 15 13 10 9 14 13 0 14 13 1 9 2 3 7 7 10 9 14 13 1 9 14 13 0 9 7 14 14 13 1 10 9 10 9 2 15 13 1 9 15 2 7 3 7 10 9 14 13 14 13 1 0 9 2
7 14 13 14 13 15 15 2
13 7 3 2 12 0 9 2 13 10 9 10 9 2
24 13 7 2 7 10 9 14 13 0 2 14 13 14 13 10 9 1 15 13 3 10 9 15 2
26 3 2 13 14 13 10 9 9 2 10 15 14 13 9 1 9 10 15 13 13 1 10 0 9 9 2
24 15 13 3 1 9 10 9 7 1 9 15 10 9 9 13 1 9 10 9 0 7 0 9 2
1 9
20 10 9 14 13 3 10 9 15 13 7 3 3 10 9 15 13 10 9 15 2
11 10 0 9 14 13 1 9 7 1 9 2
13 13 1 10 9 0 9 9 1 10 0 9 9 2
39 3 1 10 9 12 10 9 10 9 2 14 13 0 9 1 9 10 0 9 7 2 1 9 2 1 9 9 10 0 9 1 9 9 1 9 15 10 9 2
1 9
37 2 14 13 15 9 1 14 13 10 9 10 0 0 7 10 9 13 3 9 10 9 15 2 2 13 10 9 9 9 9 0 9 10 0 9 9 2
1 9
31 10 9 15 13 1 0 9 15 9 9 7 2 3 13 0 10 9 15 2 1 9 15 10 9 10 12 9 9 13 3 2
5 13 3 12 9 2
46 13 3 14 13 7 10 9 14 13 1 9 3 1 10 9 10 12 0 9 1 9 2 3 7 7 15 10 9 10 9 15 14 13 1 9 14 13 10 9 15 13 1 10 0 9 2
20 13 7 13 0 10 9 10 9 15 3 0 9 10 9 9 2 9 7 9 2
19 10 9 12 0 9 2 12 1 10 15 13 1 9 0 9 2 13 1 2
22 3 10 0 9 9 9 13 13 1 12 1 12 9 2 7 13 14 13 10 0 9 2
42 13 7 13 1 9 2 14 13 7 14 13 10 9 15 1 15 7 14 13 0 14 13 10 9 12 1 10 9 3 1 10 0 9 9 7 9 7 10 9 0 9 2
15 10 9 10 9 13 7 13 9 1 9 7 10 0 9 2
16 10 9 15 13 3 15 1 0 15 2 7 13 14 15 13 2
14 0 14 13 7 15 10 9 14 13 3 0 1 9 2
37 10 12 10 9 13 1 12 9 2 7 10 12 1 12 2 15 13 7 10 0 12 9 10 9 13 12 9 1 0 9 3 1 10 9 10 9 2
13 13 10 9 15 1 10 9 10 9 10 2 9 2
16 3 2 10 9 13 10 9 1 9 12 2 7 13 10 12 2
10 14 13 3 14 13 3 0 10 9 2
33 10 9 15 13 14 13 3 7 13 10 9 2 3 2 7 13 1 9 15 1 10 2 9 2 0 15 10 9 14 13 0 9 2
17 10 0 9 13 7 3 7 13 14 13 10 9 10 9 10 9 2
44 10 9 13 1 0 9 12 0 9 3 10 9 7 13 2 3 1 10 9 2 10 0 9 7 10 9 9 2 12 9 2 9 9 2 9 2 9 2 9 2 9 2 9 2
33 1 10 9 15 14 13 14 13 10 0 2 9 10 9 2 2 3 7 14 13 10 9 1 9 9 15 13 1 9 10 0 9 2
54 10 9 13 1 9 2 12 9 3 10 9 2 7 10 9 2 10 15 13 1 9 10 9 2 13 1 9 1 9 2 10 15 1 10 9 15 13 9 2 1 9 12 9 14 13 10 9 15 7 15 12 14 13 2
16 10 9 9 13 12 10 9 7 10 0 12 13 10 9 9 2
56 15 10 9 15 13 10 0 9 9 1 9 2 9 7 9 13 1 10 9 1 12 0 9 2 10 9 10 9 7 10 9 15 13 10 0 9 1 10 9 7 10 0 9 9 15 0 1 10 9 7 10 9 13 1 9 2
21 3 2 10 2 9 13 2 7 10 0 9 14 13 14 13 0 2 3 10 9 2
13 10 9 13 1 9 7 13 1 9 7 10 9 2
36 3 2 13 7 13 0 14 13 10 0 9 15 14 13 1 9 10 9 10 9 10 0 9 7 14 13 10 13 9 10 0 9 15 13 3 2
41 1 10 9 15 2 10 9 9 10 2 2 9 9 2 13 1 0 9 10 9 7 2 1 10 9 7 13 3 0 9 1 10 0 9 2 10 9 13 9 2 2
28 15 1 10 9 15 2 13 10 9 14 13 1 15 0 9 15 13 1 0 15 9 7 14 13 1 10 9 2
19 10 9 13 13 9 7 10 0 0 9 14 13 9 7 10 9 13 2 2
32 10 0 9 3 13 7 13 1 9 15 13 15 10 9 1 9 10 9 2 3 1 10 0 9 0 9 1 9 10 0 9 2
25 9 0 9 13 10 2 7 0 9 9 9 2 0 1 10 15 13 2 13 7 13 10 9 15 2
21 14 13 14 13 7 10 9 15 13 10 0 9 10 0 9 10 9 7 10 9 2
8 3 1 15 13 14 13 9 2
3 2 9 2
40 13 14 13 7 10 9 9 13 3 10 9 9 9 0 9 15 13 10 9 2 13 10 9 7 10 9 10 9 7 13 3 10 9 15 3 0 1 10 9 2
12 13 10 9 1 15 13 10 2 14 13 0 2
19 7 14 13 1 15 2 7 14 13 9 1 15 10 9 1 0 10 9 2
38 1 10 15 13 10 9 9 1 10 9 9 2 7 13 7 1 0 9 9 13 3 0 9 1 10 9 9 9 15 13 1 10 0 3 1 10 9 2
14 15 12 3 13 0 1 9 2 1 15 13 1 9 2
17 10 9 9 14 13 1 10 9 15 10 3 0 9 10 9 12 2
18 15 7 14 13 14 13 1 10 9 3 7 10 2 14 13 0 9 2
8 10 9 0 9 14 13 9 2
38 10 0 9 10 0 12 9 1 9 13 0 1 12 9 7 9 2 12 9 1 9 10 9 2 15 7 15 13 13 9 7 3 12 2 0 2 9 2
30 10 9 10 9 13 10 9 14 13 1 9 15 14 13 14 13 10 9 9 10 2 9 2 1 10 9 15 1 9 2
45 3 13 10 9 2 1 9 2 13 3 14 13 7 1 10 9 10 0 9 9 15 13 10 9 2 15 9 7 9 15 14 13 9 14 13 3 10 9 14 13 9 1 0 9 2
23 10 9 13 3 7 13 0 14 13 10 9 15 13 13 2 1 14 13 14 13 0 9 2
24 13 7 13 0 7 1 9 13 10 9 10 2 1 10 0 9 1 10 0 9 7 10 9 2
9 10 2 13 9 9 10 0 9 2
16 3 2 1 10 9 13 10 9 1 0 0 0 9 10 9 2
26 9 10 9 13 10 9 2 10 0 9 2 1 0 9 10 9 2 15 13 10 9 15 1 9 9 2
3 2 9 2
6 9 13 10 9 10 9
28 3 10 9 2 10 9 13 7 14 13 9 1 12 9 1 9 9 15 1 9 10 9 1 10 9 1 9 2
13 13 3 10 9 10 9 2 10 9 7 10 0 2
24 1 9 2 10 9 15 14 13 10 0 9 15 13 10 9 15 7 14 13 10 9 10 9 2
21 10 9 10 9 13 3 1 10 9 10 9 2 1 9 12 9 1 10 0 9 2
25 10 9 2 13 1 10 0 9 10 9 10 9 15 13 10 9 10 0 0 9 1 10 0 9 2
32 3 9 7 9 13 14 13 0 7 0 9 1 10 9 10 9 1 7 1 15 13 1 9 9 2 10 9 15 13 1 3 2
25 3 1 9 9 9 7 9 15 13 3 9 10 0 9 10 0 9 7 9 13 0 9 0 9 2
13 9 9 13 1 9 0 7 1 0 9 10 9 2
15 1 9 13 7 10 9 15 13 10 9 0 10 9 15 2
3 2 9 2
15 10 9 7 10 9 13 0 10 9 15 14 13 14 13 2
41 10 9 10 9 2 9 9 9 2 13 1 9 15 13 1 0 9 10 2 2 7 10 9 15 14 13 1 10 2 10 9 1 9 10 0 9 9 2 9 9 2
21 3 1 0 9 1 10 0 9 13 9 2 1 10 15 10 9 9 9 9 9 2
19 15 13 1 9 1 9 10 2 10 9 2 1 9 14 13 1 10 9 2
23 13 0 15 15 14 13 10 9 14 13 10 3 0 0 9 1 10 9 10 9 10 2 2
14 10 9 13 10 9 15 1 0 9 10 9 10 9 2
33 13 1 2 9 2 14 13 14 13 7 3 13 10 0 9 10 15 13 13 1 9 2 10 9 13 13 3 10 9 10 0 9 2
23 10 9 9 10 9 2 9 9 2 13 7 2 10 9 13 0 14 13 10 9 0 2 2
26 10 9 9 10 9 13 3 1 10 0 9 2 1 9 9 2 10 0 9 10 9 1 3 0 9 2
23 10 0 13 7 13 10 9 3 1 10 9 7 0 1 15 13 1 7 3 3 1 9 2
19 3 2 3 1 9 2 10 9 12 13 14 13 9 1 0 9 10 9 2
12 3 2 10 0 14 13 14 13 9 1 9 2
60 10 0 9 2 1 10 9 15 2 13 10 9 15 14 13 3 1 10 0 9 2 3 13 1 9 15 1 10 9 10 9 10 9 2 10 9 10 0 9 2 10 12 9 10 9 7 9 9 7 10 9 9 1 9 9 7 9 10 9 2
44 1 9 2 10 0 10 9 9 2 9 9 2 13 7 10 9 13 2 10 0 9 9 2 1 9 7 2 10 9 9 2 9 2 7 0 9 13 3 9 2 1 10 9 2
43 1 15 10 9 2 10 9 0 9 2 10 15 10 9 13 3 2 13 10 9 10 9 9 10 0 9 10 15 13 10 0 9 9 2 1 9 1 10 15 13 1 9 2
15 7 2 15 14 13 14 13 3 9 7 9 1 10 9 2
24 13 10 0 9 2 7 9 3 1 12 9 2 1 10 0 9 10 9 10 9 1 10 9 2
23 10 0 13 10 0 9 9 2 9 9 0 9 2 15 13 14 13 9 1 10 9 9 2
27 7 10 9 13 14 13 1 10 9 2 10 0 9 13 3 1 10 9 2 14 13 10 0 9 10 9 2
15 1 15 10 9 13 3 13 14 13 1 9 10 9 15 2
37 10 0 9 13 2 7 3 14 13 10 9 1 0 9 2 7 13 9 1 9 9 7 9 10 0 0 9 1 10 9 0 9 1 10 9 2 2
34 13 9 3 10 9 15 13 1 15 13 1 0 9 1 10 9 15 2 7 15 13 1 0 15 9 7 14 13 7 9 3 1 15 2
13 9 2 9 0 10 0 9 10 2 13 1 9 9
1 9
17 13 3 13 7 10 9 10 0 9 13 7 1 9 3 10 9 2
17 1 15 13 10 0 9 2 10 9 2 10 9 0 9 7 15 2
53 15 13 7 13 14 13 10 9 10 9 10 0 0 9 3 1 9 0 2 3 1 9 1 10 9 2 7 3 7 1 9 1 10 9 2 1 10 0 9 2 7 13 7 13 14 13 3 10 9 7 10 12 2
23 14 13 10 9 10 0 9 10 9 2 10 15 14 13 7 10 15 13 14 13 1 9 2
11 14 13 1 9 1 9 3 14 15 13 2
27 1 10 9 15 2 10 9 9 10 9 13 7 2 10 0 9 14 13 1 10 9 7 13 3 0 2 2
35 13 10 12 9 3 10 2 9 2 13 3 10 9 15 1 10 0 2 10 9 7 10 9 2 9 15 13 10 9 10 2 0 9 2 2
31 1 9 10 9 10 0 9 13 1 9 2 7 7 14 13 3 3 2 3 1 10 9 10 9 7 10 9 9 1 9 2
60 13 9 9 2 1 10 9 0 9 2 1 9 10 9 2 1 15 13 7 13 0 2 0 9 0 9 2 3 1 10 9 9 9 7 9 9 9 13 10 0 9 7 3 2 1 9 2 13 1 10 9 2 10 15 13 7 15 1 9 2
45 10 9 13 10 9 1 10 9 10 9 10 9 1 9 9 9 2 15 13 10 9 2 7 2 14 14 13 10 9 1 10 9 0 9 9 1 10 9 15 10 9 10 12 2 2
29 10 9 10 9 1 10 0 9 10 9 13 10 0 9 1 9 9 7 9 2 10 15 14 13 1 9 9 9 2
24 1 10 0 9 10 2 13 13 10 9 12 9 9 7 12 9 1 10 15 13 9 10 9 2
13 1 3 10 0 9 13 14 13 10 9 10 9 2
26 1 9 13 10 9 3 7 10 9 14 13 10 0 9 1 13 9 7 1 9 9 9 7 9 15 2
8 14 13 13 3 10 9 9 2
18 13 0 10 9 1 10 9 15 7 15 13 7 13 12 3 0 9 2
14 3 2 1 9 13 9 9 9 7 9 1 0 9 2
10 10 0 9 13 14 13 9 10 9 2
12 13 10 0 9 1 9 3 13 10 0 9 2
21 10 9 10 9 13 1 9 10 9 7 13 3 1 0 1 9 3 1 0 9 2
7 15 13 1 10 9 15 2
23 13 7 13 7 1 0 0 9 14 13 1 0 9 7 1 0 9 0 10 9 1 9 2
9 13 1 10 9 10 9 10 9 2
11 10 12 9 13 1 9 12 1 10 9 2
48 10 2 9 2 13 1 10 9 9 9 3 7 2 13 2 2 10 9 9 13 14 13 3 1 0 0 9 1 0 9 10 9 2 7 14 13 0 9 9 10 9 9 1 9 10 2 2 2
47 7 13 13 1 0 9 2 13 7 10 9 10 9 1 9 14 13 14 13 1 0 10 0 0 9 10 2 2 3 7 14 13 3 10 0 9 1 10 9 7 10 9 1 10 0 9 2
38 10 9 13 3 10 9 15 1 10 9 10 0 9 14 13 10 9 10 9 1 0 10 9 10 0 9 1 10 9 2 15 13 1 10 9 10 9 2
35 7 2 1 10 15 9 2 13 10 0 9 1 10 0 15 9 7 10 9 7 13 3 7 13 9 10 9 14 15 13 1 10 0 9 2
36 10 9 9 13 14 13 0 3 12 9 3 1 10 9 10 9 2 3 7 0 15 14 13 14 13 9 1 10 9 15 7 14 13 15 13 2
33 7 7 10 9 10 9 13 10 9 1 9 10 9 10 9 3 13 15 9 9 14 15 13 10 9 14 13 3 10 9 15 9 2
19 3 13 10 0 9 10 9 2 14 13 14 13 10 0 9 1 9 9 2
7 3 12 9 13 10 9 9
29 10 0 9 2 10 9 2 10 9 7 10 9 10 9 14 13 15 15 13 10 9 7 13 1 0 10 9 15 2
5 14 13 0 9 2
1 9
14 3 2 10 2 13 3 0 1 10 9 1 10 9 2
34 13 10 15 9 10 9 2 10 15 2 3 2 13 10 9 7 10 9 3 1 10 9 0 9 10 0 9 14 13 3 10 0 9 2
38 1 14 13 1 2 9 2 10 9 13 13 14 13 1 0 9 9 10 0 9 10 9 7 10 9 2 1 10 9 7 13 15 9 1 10 0 9 2
8 13 10 0 9 3 10 9 2
10 14 13 14 13 0 9 1 0 9 2
23 10 9 10 9 10 9 13 1 12 2 7 9 1 10 9 13 10 12 9 2 10 9 2
81 3 13 10 9 10 9 2 10 9 15 13 0 0 9 15 13 1 0 9 7 1 9 10 9 10 9 2 3 1 9 2 7 13 3 2 7 15 1 15 10 9 9 2 14 14 13 14 13 3 7 13 14 13 1 0 9 9 10 15 13 10 0 9 10 0 9 9 2 3 7 7 13 9 1 10 9 10 9 15 2 2
42 3 2 10 0 9 10 0 9 13 14 13 1 9 1 10 9 10 9 2 13 7 2 1 14 13 15 0 9 2 10 9 9 9 14 13 3 14 13 10 9 2 2
20 3 2 1 9 13 3 1 10 9 3 1 12 0 9 1 10 9 1 9 2
34 1 9 10 9 2 14 13 10 0 9 2 3 1 15 15 13 10 2 9 10 0 9 2 7 13 10 12 0 0 9 1 9 15 2
17 0 15 13 13 9 2 7 10 9 9 13 10 9 15 3 3 2
34 15 13 7 10 9 14 13 9 1 10 12 9 2 9 7 9 2 1 0 9 10 9 2 2 13 10 9 9 2 9 9 10 9 2
7 10 12 13 1 10 9 2
22 3 7 1 9 9 2 10 9 15 14 13 9 1 9 9 2 0 9 7 3 9 2
7 15 13 3 1 10 9 2
10 10 9 9 13 10 9 2 9 2 2
10 10 0 9 7 9 13 1 10 9 2
8 10 9 1 10 9 13 0 2
20 10 9 13 14 13 10 12 15 9 3 1 12 9 2 3 1 9 10 9 2
22 10 9 10 9 13 10 9 9 1 12 9 2 7 10 0 13 1 10 9 1 12 2
41 10 9 9 10 9 13 3 7 2 10 9 10 9 10 2 1 9 13 9 1 10 9 2 7 10 9 10 9 7 10 9 9 14 13 7 13 9 1 9 2 2
40 10 9 0 1 10 13 9 7 10 0 9 2 10 0 0 1 10 0 9 2 10 9 2 10 15 13 7 13 1 0 9 10 9 13 15 0 9 10 9 2
21 13 3 10 2 9 9 2 10 9 15 2 7 13 1 9 14 13 10 9 15 2
21 13 0 9 9 3 10 0 9 2 3 3 7 3 7 3 0 9 9 1 9 2
18 3 1 15 9 13 10 9 14 13 7 14 13 10 9 1 0 9 2
34 13 1 15 2 7 13 3 0 14 13 10 0 3 1 10 9 15 1 10 0 9 7 14 13 3 10 0 0 1 10 3 9 15 2
29 10 9 10 9 13 3 7 14 13 1 10 9 10 9 1 12 9 7 7 9 15 14 13 10 9 9 2 9 2
49 13 3 1 12 1 10 9 10 9 0 2 0 7 0 0 2 1 15 10 9 15 2 10 15 3 13 2 13 7 13 14 13 10 9 13 10 9 2 7 3 13 14 13 12 10 9 1 2 2
31 15 9 13 10 9 14 13 14 13 3 7 7 10 9 15 13 2 7 10 9 13 14 13 10 9 1 9 2 7 13 2
45 10 9 14 13 14 13 7 13 1 9 9 7 7 1 9 15 13 3 1 9 10 9 13 15 9 3 1 10 3 0 9 10 9 1 3 0 9 2 3 10 9 7 10 9 2
16 3 2 3 13 3 9 1 10 9 15 10 9 10 9 9 2
22 1 9 13 14 13 3 3 1 15 1 10 9 15 13 15 9 1 10 9 10 9 2
6 13 9 1 0 9 2
41 7 13 14 13 15 9 1 9 15 2 15 14 13 10 9 2 3 13 1 15 15 9 2 7 1 10 9 7 13 2 3 2 10 9 9 1 2 9 15 2 2
20 10 9 10 9 13 9 7 9 10 0 9 15 13 1 9 1 10 0 9 2
11 15 13 3 10 9 15 13 15 3 3 2
28 9 9 2 14 13 3 14 13 10 9 1 10 0 9 9 15 13 1 9 15 7 1 10 9 15 15 13 2
36 10 9 10 9 9 1 0 9 13 14 13 1 10 9 9 2 1 10 15 14 13 0 1 10 9 10 2 9 1 14 13 10 9 10 9 2
34 3 2 3 13 10 9 10 0 9 2 10 9 10 0 9 12 13 10 9 10 9 10 9 2 1 10 15 13 13 9 1 10 9 2
32 13 7 7 15 15 15 13 7 1 9 14 13 7 13 14 15 13 3 2 14 13 10 9 10 9 10 0 9 15 1 9 2
45 10 9 15 13 1 9 13 14 13 15 10 9 7 2 7 10 9 3 14 13 7 13 3 7 7 13 9 14 13 0 2 13 10 15 0 9 14 13 15 10 9 1 9 15 2
7 12 0 1 9 1 0 9
18 15 13 10 9 14 13 10 9 10 9 0 9 7 10 9 15 0 2
12 10 9 13 14 13 10 3 3 15 10 9 2
24 10 9 10 9 2 0 9 12 2 2 15 1 10 15 13 13 2 13 1 10 0 9 15 2
37 9 1 10 9 10 9 13 10 9 14 13 1 10 9 10 0 9 1 9 2 0 1 9 2 7 1 0 10 9 13 0 10 9 1 10 9 2
7 13 0 2 0 2 0 2
21 13 7 13 14 13 1 9 1 9 15 9 7 10 0 9 14 14 13 0 9 2
61 7 7 10 9 10 9 13 13 1 9 9 9 9 2 10 15 1 10 9 2 2 2 1 9 13 1 10 9 1 0 2 10 0 9 13 14 13 10 9 7 13 10 0 9 13 3 1 9 9 3 1 10 9 2 7 14 13 1 9 9 2
41 1 9 13 12 9 2 3 3 1 10 9 9 10 0 9 2 10 9 2 10 9 2 10 9 2 3 3 7 10 0 1 9 9 3 1 10 9 7 10 9 2
13 1 9 12 10 9 9 14 13 9 1 10 9 2
19 3 10 9 13 12 3 9 1 10 9 9 1 9 9 2 3 1 9 2
19 3 2 14 13 9 14 13 12 9 3 7 3 1 14 13 9 10 9 2
5 1 9 10 9 2
15 13 14 13 10 9 10 2 9 7 15 13 7 13 3 2
9 10 9 10 9 9 9 13 10 9
21 14 13 3 14 13 10 9 2 9 7 3 10 9 2 9 1 10 0 9 15 2
30 3 13 14 13 15 10 9 2 10 0 9 2 10 0 9 2 10 9 10 9 10 9 1 10 9 7 10 0 9 2
10 3 2 13 3 3 0 1 10 9 2
15 13 1 0 7 3 3 1 0 9 7 3 13 14 13 2
16 10 0 9 10 9 13 1 10 0 9 10 9 7 0 15 2
28 10 9 13 1 0 9 9 2 7 13 10 9 9 1 9 7 9 14 13 1 14 13 7 10 9 0 9 2
19 10 0 13 10 9 10 0 9 1 0 9 2 1 12 2 1 10 9 2
10 10 9 9 13 9 1 14 0 9 2
14 3 2 13 7 13 3 0 9 3 9 10 0 9 2
7 9 9 13 12 9 1 2
9 3 14 13 14 13 7 15 15 2
11 10 9 14 13 3 2 7 10 9 13 2
26 10 9 10 9 13 14 13 15 9 9 10 0 0 9 7 3 15 13 10 9 15 14 13 14 13 2
26 3 2 10 9 13 13 1 9 9 7 13 13 7 13 0 10 9 10 15 13 13 1 10 9 9 2
27 1 9 3 1 10 9 13 0 9 9 2 3 1 12 2 7 7 9 3 9 2 9 2 9 2 9 2
38 10 12 13 10 0 7 10 12 10 0 1 10 0 9 15 13 3 2 9 2 10 0 9 2 3 1 0 9 10 9 9 10 9 9 1 9 9 2
11 10 9 7 10 9 13 3 9 1 9 2
10 13 3 7 13 12 0 9 1 9 2
30 13 7 10 9 9 9 13 1 12 9 12 1 9 7 10 9 15 13 10 0 9 10 9 15 13 9 1 0 9 2
18 10 0 9 15 14 13 14 13 1 9 10 0 9 7 10 0 9 2
25 10 9 10 0 9 13 7 2 10 0 9 1 9 13 10 0 1 9 2 1 10 0 9 2 2
57 10 0 9 10 0 9 13 10 0 9 14 2 13 10 0 9 1 9 15 13 10 0 3 9 1 0 15 9 2 7 15 15 13 0 1 9 1 9 10 9 15 2 1 9 2 1 9 10 9 15 2 7 1 9 9 2 2
32 10 9 1 9 7 9 1 10 9 10 9 13 7 10 9 2 15 12 1 10 9 15 13 1 0 9 2 13 1 0 9 2
27 10 9 2 9 9 10 0 9 13 14 13 9 1 9 1 10 9 14 0 9 2 1 10 9 10 2 2
30 10 9 15 14 13 0 10 0 9 1 10 0 2 10 9 15 13 3 12 0 9 15 13 1 10 9 10 9 9 2
12 1 9 15 3 13 10 9 15 13 14 13 2
28 1 3 2 9 1 10 9 10 9 9 7 1 10 0 0 9 10 0 9 1 10 9 13 1 9 10 9 2
30 3 10 0 9 13 1 0 9 0 9 2 9 2 1 9 10 9 2 7 2 13 10 9 14 13 1 10 9 2 2
57 1 10 9 15 2 10 9 9 13 7 14 13 15 9 1 10 0 9 1 9 15 13 1 9 7 1 15 13 13 9 9 15 10 9 15 13 9 10 9 2 7 1 12 1 10 9 13 7 10 0 10 9 10 9 10 9 2
26 1 9 13 3 12 9 9 2 10 15 10 0 9 13 15 9 1 9 15 1 10 0 9 10 9 2
22 10 9 10 9 13 0 7 13 13 3 1 10 9 15 3 0 0 9 2 10 9 2
25 14 13 14 13 7 1 2 9 7 2 7 13 1 10 9 2 14 13 15 10 9 10 9 15 2
20 1 10 15 9 2 13 14 13 0 9 9 1 9 2 1 9 7 1 9 2
14 10 9 13 0 9 2 7 13 10 0 9 10 9 2
12 13 7 13 0 10 0 9 13 1 10 9 2
34 10 1 9 9 13 3 13 9 9 10 0 9 1 9 1 0 9 1 9 10 9 10 9 15 7 10 9 10 9 15 1 15 9 2
34 13 7 15 0 9 15 13 13 1 10 9 13 14 13 0 9 15 13 1 0 9 9 1 10 9 2 10 3 9 7 10 0 9 2
13 10 9 13 1 10 9 12 0 1 15 10 9 2
20 10 9 13 10 9 9 2 1 9 2 10 15 13 10 9 0 1 10 9 2
21 10 9 2 10 9 13 0 9 2 1 15 14 13 15 1 10 0 9 10 9 2
8 13 3 7 9 15 13 9 2
36 10 0 9 15 2 9 2 9 2 13 1 9 10 0 9 15 2 9 2 3 2 9 10 9 2 15 13 1 10 12 9 15 13 1 9 2
22 3 2 10 9 13 13 0 9 0 9 2 7 0 9 7 9 13 7 10 9 15 2
14 0 1 0 0 9 13 10 9 10 0 9 10 9 2
21 7 14 13 1 9 2 3 10 0 1 15 14 14 13 3 14 13 10 9 15 2
18 13 7 14 13 0 10 9 1 0 9 1 0 7 0 9 15 9 2
11 0 15 13 0 9 7 13 13 1 9 2
12 3 2 10 9 14 13 15 9 1 0 9 2
43 7 2 9 9 2 1 9 9 2 7 13 7 15 14 13 0 15 9 2 13 0 9 1 10 9 9 1 9 3 13 14 13 10 9 2 0 15 14 14 13 15 9 2
29 10 9 15 3 3 13 1 9 10 9 14 13 10 0 9 1 10 12 9 7 14 13 10 0 9 1 10 9 2
27 13 10 0 15 13 10 9 7 13 10 9 3 10 0 9 1 10 9 10 0 9 9 1 0 0 9 2
58 7 13 10 9 2 10 3 3 0 1 10 9 15 13 10 9 2 2 15 13 7 10 9 15 13 10 9 14 14 13 14 13 3 1 10 0 9 7 10 0 7 7 15 9 2 3 10 0 9 7 10 9 9 10 9 15 13 2
8 13 14 15 13 14 15 13 2
31 2 10 12 9 2 7 7 9 2 13 0 7 13 0 1 10 0 2 7 3 13 1 0 9 2 2 13 10 0 9 2
24 3 2 10 9 13 10 9 15 10 9 10 9 7 10 9 10 9 13 7 15 1 10 9 2
20 1 10 12 0 9 10 0 9 13 3 0 1 3 1 10 0 9 10 9 2
29 10 9 10 2 2 9 9 2 13 7 2 10 0 9 9 0 9 14 13 9 1 15 9 7 15 13 0 2 2
17 3 9 13 1 9 7 10 9 10 9 7 10 9 14 13 3 2
10 14 13 14 13 0 9 7 0 9 2
23 10 9 13 10 9 10 9 10 9 9 10 12 2 10 9 9 2 10 15 7 13 3 2
53 3 0 13 10 9 15 13 7 10 2 1 0 9 1 10 9 1 15 13 13 10 0 9 1 10 0 9 0 0 2 9 15 13 3 2 9 1 15 13 0 9 2 2 13 1 9 10 2 9 1 9 2 2
34 10 9 13 10 9 2 13 7 2 10 9 10 9 13 3 1 9 2 7 13 1 10 9 14 14 13 3 9 1 0 9 10 9 2
31 10 0 0 9 9 9 13 10 9 1 10 9 2 3 0 2 3 7 13 14 13 10 9 15 10 9 13 10 9 2 2
30 10 12 9 10 9 9 1 0 15 9 13 9 1 9 15 14 13 10 9 10 0 9 15 1 3 13 10 9 9 2
51 3 1 10 9 10 9 1 10 9 1 9 2 3 10 9 10 9 13 10 0 1 14 13 2 7 14 13 10 9 1 10 9 10 9 2 15 13 10 0 7 10 3 0 1 10 0 9 10 15 13 2
8 13 1 9 15 10 0 9 2
26 3 2 1 9 13 10 9 10 9 9 2 15 13 10 0 9 2 7 7 10 0 9 10 0 9 2
40 10 9 13 7 10 9 14 13 1 9 12 9 9 3 1 0 12 9 1 9 1 9 3 10 9 9 2 10 9 9 9 2 10 0 9 7 10 0 9 2
9 12 1 10 9 13 1 0 9 2
27 13 12 1 10 0 9 10 9 2 7 13 0 0 9 1 10 9 10 9 2 7 13 3 1 10 9 2
40 3 13 0 14 13 7 14 13 3 1 10 9 15 2 7 1 9 10 9 2 7 14 13 14 13 10 0 9 1 10 9 15 14 13 3 1 10 0 9 2
45 10 0 9 13 14 13 2 7 2 7 1 10 9 7 10 9 13 13 2 14 13 14 13 10 9 15 13 10 2 14 13 1 10 9 9 2 10 15 1 9 10 9 13 3 2
40 9 10 0 9 1 9 13 10 9 9 1 9 3 1 9 9 9 10 9 9 2 7 1 12 0 9 15 13 10 9 1 9 15 13 1 3 1 10 9 2
23 10 9 10 9 2 10 9 2 13 3 1 12 9 2 10 15 13 0 9 1 9 15 2
14 10 12 9 14 13 1 2 9 2 2 1 12 9 2
9 13 7 3 13 3 10 9 15 2
7 10 12 9 13 12 9 2
20 13 14 13 3 10 3 3 10 0 9 7 10 9 14 13 3 10 3 3 2
21 13 3 10 9 10 2 9 7 13 10 9 9 1 0 9 14 13 1 12 9 2
10 13 15 9 14 13 9 1 10 9 2
25 10 9 9 9 1 9 15 13 7 13 1 10 9 2 1 10 15 13 3 7 0 9 7 9 2
22 7 2 13 1 9 7 13 0 2 3 7 13 1 10 9 3 7 7 13 10 9 2
10 10 0 9 13 10 9 1 0 9 2
9 10 0 9 13 1 9 10 9 2
15 0 15 13 1 10 0 9 2 1 3 0 7 13 9 2
12 13 12 1 10 0 0 9 10 0 12 9 2
11 10 9 13 10 9 10 9 1 10 9 2
35 2 1 10 9 7 10 9 15 13 10 9 13 3 1 10 3 0 9 2 10 9 10 9 9 13 9 9 2 13 10 9 10 0 9 2
11 9 9 2 13 15 14 13 1 10 9 2
41 13 10 9 15 13 15 7 14 13 10 9 15 3 9 0 9 10 9 1 10 3 2 7 3 13 3 1 10 9 2 1 0 15 13 14 13 3 1 0 9 2
32 13 1 10 0 9 7 13 1 3 3 10 9 15 13 1 9 2 15 13 3 10 9 10 3 9 2 13 14 13 0 9 2
37 10 9 13 3 10 0 9 2 7 14 13 14 13 3 10 0 9 1 10 9 10 9 1 9 1 10 0 9 2 1 9 10 9 15 13 3 2
35 10 9 2 1 10 9 15 1 10 0 9 10 9 1 10 9 15 1 9 10 9 2 10 9 2 13 10 0 0 9 1 12 3 9 2
26 1 10 0 9 10 9 2 10 9 13 1 10 0 9 10 13 9 9 1 10 9 10 1 9 9 2
23 1 10 9 15 13 3 14 13 1 10 9 2 14 13 14 13 12 15 13 3 10 0 2
42 3 2 1 10 9 10 0 9 13 10 9 10 0 9 3 1 10 9 2 15 14 13 1 0 9 7 15 14 15 13 2 9 7 9 2 7 13 10 0 0 9 2
27 14 13 1 9 14 13 9 9 0 1 15 15 13 3 2 3 1 10 15 10 9 9 15 13 3 0 2
11 13 3 7 7 10 0 9 14 15 13 2
31 2 10 9 10 9 9 13 10 9 10 9 9 0 9 1 10 9 3 10 9 15 2 3 7 10 9 15 1 9 2 2
12 14 13 15 13 3 1 15 2 0 9 2 2
27 13 7 10 9 10 9 15 1 10 9 14 13 0 7 14 13 0 9 1 0 9 1 15 13 1 9 2
21 13 3 10 9 9 2 0 3 2 9 10 0 2 2 3 9 1 0 9 9 2
14 10 9 3 1 10 12 9 10 9 13 1 0 15 2
8 13 10 0 9 2 10 9 2
23 3 3 1 10 9 13 10 9 9 2 9 7 9 2 10 15 13 13 1 12 0 9 2
16 3 15 13 2 9 2 13 3 1 10 9 3 0 7 0 2
39 13 3 7 0 9 13 14 13 1 10 9 9 10 0 9 0 9 9 1 9 15 14 13 9 10 9 2 7 13 3 1 15 10 9 10 9 9 9 2
17 13 3 0 14 13 10 9 3 1 10 9 10 12 9 1 15 2
36 1 10 0 9 13 3 14 13 3 1 0 9 9 10 0 9 3 9 2 3 9 2 3 9 1 10 15 14 13 3 1 10 9 10 9 2
16 9 9 9 9 9 2 15 13 14 13 1 9 10 9 15 2
46 0 0 9 13 15 10 9 1 10 9 7 10 9 2 10 9 10 15 13 10 0 9 1 10 9 2 1 10 9 2 12 1 10 12 9 9 2 9 2 10 15 13 7 10 9 2
14 1 0 9 9 10 9 13 0 2 7 1 15 14 2
16 10 9 13 7 0 9 13 14 13 10 9 1 10 9 2 2
34 15 13 10 9 10 9 9 10 9 7 10 9 15 13 7 13 0 15 13 13 10 9 2 1 10 12 3 9 9 2 3 9 15 2
25 3 2 10 9 9 13 1 9 12 1 10 9 9 2 1 9 10 9 10 12 10 9 9 12 2
3 2 9 2
33 10 9 9 9 1 9 15 1 10 9 10 0 9 13 7 10 9 3 13 7 13 3 1 9 7 15 7 14 13 14 13 9 2
26 12 1 10 9 15 13 13 2 3 2 14 13 1 0 10 9 10 0 9 1 9 15 1 10 12 2
43 10 9 7 10 9 9 13 0 14 13 10 13 9 10 9 1 10 9 2 10 15 14 13 3 0 7 0 14 13 1 0 9 1 0 9 1 9 7 1 9 10 9 2
31 1 0 9 15 13 2 10 9 13 14 13 0 9 3 9 7 0 9 2 10 0 9 10 9 7 10 9 10 9 12 2
35 13 1 2 9 2 14 13 14 13 7 10 0 9 10 9 9 13 3 7 10 9 15 13 14 13 3 10 9 7 10 9 7 10 9 2
10 3 2 13 0 3 1 10 0 9 2
12 3 1 10 9 13 10 9 1 10 0 9 2
19 10 0 9 13 13 1 0 9 3 15 13 9 7 9 1 0 9 2 2
48 10 9 13 1 10 12 9 7 10 9 10 9 1 9 1 9 3 2 3 7 1 9 1 9 9 10 2 3 14 13 14 13 3 2 9 10 0 9 10 15 14 13 14 13 10 9 9 2
36 10 0 9 13 7 10 0 9 13 0 9 1 10 9 7 2 9 10 9 13 10 9 10 9 10 0 9 13 7 10 9 10 0 9 2 2
32 10 9 10 2 9 1 9 2 1 2 2 9 9 2 13 1 9 15 1 10 2 7 2 10 9 10 9 13 1 0 9 2
7 1 15 2 1 9 13 2
25 10 9 10 2 9 9 9 13 12 1 15 10 9 2 2 13 10 9 9 10 9 2 9 9 2
39 0 9 15 13 10 9 7 9 9 2 12 2 2 2 9 15 13 0 1 10 9 9 1 0 0 9 9 2 9 2 9 7 1 15 13 7 0 9 2
7 0 1 15 13 10 9 2
20 1 9 2 10 9 9 1 12 9 15 13 10 12 13 10 12 9 10 12 2
29 10 9 9 13 1 10 9 12 9 3 2 1 10 15 10 0 9 15 13 1 9 9 7 10 0 1 9 9 2
29 1 10 9 10 9 2 10 9 13 3 0 3 10 9 10 15 13 14 13 10 9 10 9 9 7 10 0 9 2
9 10 0 9 13 13 10 9 15 2
19 12 9 10 0 9 13 0 1 10 9 15 1 10 9 0 9 1 9 2
37 10 9 3 1 15 10 9 13 14 13 10 9 1 10 0 9 10 9 3 1 10 9 9 2 9 9 2 9 2 9 2 9 2 9 7 9 2
24 3 2 10 9 1 9 13 2 3 7 14 13 10 0 9 7 0 10 0 9 13 1 9 2
24 10 9 13 10 9 1 9 0 1 10 9 15 2 10 15 13 12 1 10 3 0 10 9 2
19 1 15 13 10 9 1 9 2 14 13 0 7 10 9 14 13 0 9 2
22 7 3 13 14 13 7 10 9 15 1 9 9 2 15 3 3 13 2 14 13 3 2
30 3 2 7 14 13 15 0 0 9 2 0 10 9 1 9 14 13 3 14 13 1 10 0 9 0 7 0 9 9 2
20 1 10 15 9 13 7 10 9 9 14 13 3 15 1 9 3 0 9 9 2
11 13 0 7 1 10 9 2 0 9 2 2
21 10 9 9 13 3 15 9 0 9 1 14 13 10 9 10 9 15 13 1 9 2
16 3 1 10 12 10 9 10 0 9 13 10 0 9 1 9 2
12 1 10 9 10 9 13 10 0 0 9 9 2
17 10 9 13 14 13 0 9 9 10 9 7 10 9 1 0 9 2
25 3 13 10 9 15 2 9 2 10 9 13 1 10 9 7 10 0 9 10 0 9 1 10 9 2
17 14 13 14 13 3 9 2 7 0 9 10 0 9 15 13 0 2
26 3 2 10 0 9 10 0 9 7 10 0 0 9 2 3 7 10 9 3 1 10 9 9 2 13 2
17 1 10 12 9 10 9 2 13 3 9 1 10 9 9 10 9 2
1 9
19 10 9 9 7 13 10 0 9 9 7 13 3 3 13 14 13 10 9 2
1 9
23 10 9 10 9 9 13 1 15 3 1 10 9 15 13 14 13 2 13 15 3 1 9 2
6 13 10 9 10 9 2
11 1 9 2 13 10 0 9 1 10 9 2
12 10 12 9 2 10 0 9 13 3 3 0 2
11 9 15 13 10 9 14 13 3 10 0 2
10 7 2 10 9 14 13 10 9 15 2
19 10 9 13 3 0 9 7 9 1 9 3 13 3 0 9 1 10 9 2
38 0 9 13 7 10 0 9 10 9 13 1 12 12 3 1 3 12 9 2 1 10 12 1 10 12 2 9 10 0 9 9 7 10 0 9 1 9 2
8 15 14 13 3 1 10 9 2
4 9 1 9 2
20 1 3 13 14 13 3 1 9 3 7 1 0 9 7 10 0 9 10 9 2
8 10 9 13 0 9 1 9 2
24 3 2 10 9 13 10 9 9 15 13 10 0 9 9 2 1 10 15 7 10 0 9 9 2
13 10 0 13 7 10 9 15 3 1 10 0 9 2
49 10 9 1 10 9 13 3 3 1 0 9 0 9 10 15 13 3 9 10 9 2 1 0 9 7 9 1 10 0 9 2 7 13 3 0 1 10 0 9 1 9 2 1 10 0 9 10 9 2
11 10 0 15 9 13 3 1 15 10 9 2
28 1 9 15 2 10 9 13 13 0 7 0 9 2 9 0 9 7 9 2 15 0 13 10 0 9 10 9 2
20 10 9 13 10 9 15 10 9 3 13 10 9 10 9 3 1 10 9 9 2
29 10 9 9 13 3 7 2 10 9 13 1 0 9 1 14 13 7 10 9 14 13 1 15 15 15 13 9 2 2
33 10 9 13 10 9 15 1 10 12 9 2 7 7 13 7 14 14 13 14 13 1 10 9 15 14 13 0 10 9 15 13 3 2
23 3 1 15 2 13 1 10 9 1 10 9 9 2 10 15 1 0 9 13 0 3 9 2
22 13 15 0 2 3 1 10 9 3 7 1 10 9 2 13 10 2 9 10 9 12 2
23 10 9 13 7 3 1 12 9 10 0 9 10 9 13 1 12 12 1 12 1 12 9 2
21 13 3 10 9 15 13 7 2 10 2 14 13 7 0 9 3 1 0 9 2 2
36 13 3 10 3 0 9 15 13 3 14 14 13 3 10 0 9 9 2 7 3 1 0 9 13 2 1 10 9 15 2 14 13 1 0 9 2
17 3 1 15 13 13 7 10 9 10 9 2 9 2 2 9 9 2
1 9
29 10 9 10 0 9 13 1 9 10 9 14 13 9 1 9 2 1 14 15 13 2 3 13 2 1 10 0 9 2
42 10 9 10 0 7 0 9 3 7 10 0 9 10 0 9 2 10 9 10 0 9 2 3 7 10 9 10 9 1 9 13 10 0 9 15 14 13 14 13 10 9 2
32 10 12 9 15 13 3 1 12 9 13 10 0 10 15 3 13 14 13 15 0 9 1 10 15 13 1 9 15 3 10 9 2
10 10 9 13 14 13 10 9 10 0 9
26 10 9 1 9 2 9 10 9 2 13 7 2 0 1 10 0 1 9 13 13 1 14 13 3 2 2
31 10 9 10 9 14 13 3 10 9 9 9 7 10 0 9 2 7 7 10 0 9 15 13 1 10 9 10 1 9 9 2
36 1 0 9 10 9 2 10 9 9 2 13 14 13 15 10 9 0 9 2 3 13 9 1 10 0 9 10 9 7 10 0 9 10 0 9 2
15 7 2 13 10 9 15 3 1 10 9 15 15 13 0 2
4 2 2 1 2
32 1 0 9 2 14 13 14 13 10 9 10 0 9 1 9 1 9 15 15 13 1 9 7 1 9 15 15 13 3 1 9 2
81 13 3 7 13 0 7 10 9 9 14 14 13 3 14 13 0 9 1 10 9 10 9 7 7 14 13 3 10 9 14 13 10 9 1 10 9 15 13 7 1 10 9 15 14 13 2 3 10 0 3 7 10 0 9 2 3 3 7 14 13 3 9 1 10 3 14 13 14 13 10 9 7 10 0 9 9 13 3 13 0 2
29 1 9 10 9 9 9 9 9 13 10 9 1 0 9 1 10 9 7 10 0 9 10 9 10 9 7 10 9 2
51 1 0 15 2 10 9 10 9 13 14 13 10 9 15 14 13 10 0 9 2 1 9 10 9 7 1 0 0 9 2 1 9 9 7 0 9 2 7 14 13 0 10 9 1 9 10 0 7 0 9 2
10 10 9 13 2 0 2 9 1 9 2
44 3 7 1 10 9 10 12 9 10 0 9 13 14 13 9 9 10 0 9 10 9 13 14 13 10 3 13 9 15 1 9 15 2 3 3 1 9 15 10 9 13 0 9 2
25 3 10 9 7 10 9 15 14 13 10 15 0 9 14 13 3 14 13 3 1 10 9 9 9 2
16 13 7 13 14 15 13 3 13 3 7 3 10 0 15 9 2
16 0 13 7 14 13 10 12 9 9 10 9 3 1 12 9 2
35 3 2 13 7 13 1 9 2 10 9 15 13 3 1 15 13 3 10 9 2 10 15 13 3 15 15 13 10 9 7 14 13 10 9 2
46 3 1 9 10 9 9 13 9 10 9 2 10 0 9 2 10 0 9 9 1 10 9 9 2 10 0 9 2 9 10 9 9 2 9 10 3 9 9 2 7 13 1 0 0 9 2
16 13 1 9 10 0 9 7 10 0 9 7 13 1 9 15 2
47 3 7 13 10 9 10 9 10 0 9 2 10 9 10 9 13 10 9 14 13 3 1 10 9 9 2 13 0 9 9 1 10 9 10 9 2 3 1 9 3 7 1 9 10 0 9 2
42 13 14 13 1 10 9 10 9 7 14 13 7 14 13 10 0 9 7 9 15 14 13 7 15 15 14 13 1 0 9 14 13 1 0 9 1 15 1 15 15 13 2
54 1 14 13 1 2 9 7 1 2 9 2 9 10 9 1 0 9 13 10 9 10 9 1 10 9 10 9 7 14 10 9 10 9 2 0 7 15 2 1 10 15 13 14 13 10 9 0 1 15 9 13 10 9 2
22 3 1 10 9 10 0 9 13 3 1 9 3 9 7 14 13 1 9 10 9 9 2
21 1 9 7 10 1 15 9 15 1 15 14 13 10 9 10 1 9 9 10 9 2
10 9 0 9 1 9 1 9 0 9 2
44 10 9 13 10 0 9 1 2 0 9 9 2 10 0 0 9 1 9 2 1 10 9 2 1 9 9 2 10 9 12 0 9 1 9 9 1 10 9 15 1 9 1 9 2
34 1 0 15 2 10 0 9 10 9 13 10 9 2 7 9 1 10 2 13 7 3 14 14 13 10 0 1 9 2 9 10 0 2 2
18 10 0 9 10 9 9 1 0 9 9 13 13 0 9 7 13 0 2
17 13 10 0 9 7 10 9 1 10 12 2 10 15 13 14 13 2
21 10 0 9 13 3 1 12 9 3 1 15 10 9 1 10 9 10 9 1 9 2
20 3 2 13 14 13 3 0 1 9 10 0 9 7 13 0 1 9 9 15 2
11 13 7 10 9 10 9 13 10 0 9 2
16 13 1 15 9 10 9 14 13 10 9 3 12 9 10 9 2
56 10 9 1 10 15 13 10 9 10 9 2 10 9 10 9 7 10 9 10 9 1 9 15 2 3 1 10 12 9 10 9 15 2 13 10 9 15 14 13 1 10 9 10 9 7 14 13 10 9 2 7 15 13 3 0 2
50 13 14 13 7 10 9 1 10 15 13 14 13 15 10 9 10 9 2 1 14 13 1 9 10 9 15 1 10 9 10 9 14 13 14 15 13 14 13 10 9 15 13 3 15 10 9 1 0 9 2
40 1 12 7 9 2 10 9 0 9 13 1 0 9 10 0 9 10 9 7 13 7 15 13 1 9 7 7 13 10 9 1 10 9 10 9 3 1 10 9 2
32 10 9 15 13 10 9 10 9 9 10 2 7 13 10 9 14 13 10 9 9 9 10 9 15 2 9 15 14 13 10 9 2
30 10 9 9 10 9 13 7 13 0 14 13 9 2 9 9 10 0 9 2 10 15 13 14 13 1 9 10 0 9 2
15 10 9 9 0 9 13 1 9 2 1 9 10 9 9 2
26 10 0 13 2 3 7 3 2 13 14 13 1 10 9 10 0 9 7 9 2 7 0 7 15 9 2
23 3 7 12 9 13 3 1 9 7 14 13 3 14 13 10 9 0 9 1 15 10 9 2
41 3 7 1 10 0 9 3 10 0 15 2 15 13 1 10 9 3 10 9 13 0 9 1 0 9 2 3 10 0 9 10 0 9 13 3 3 1 10 9 9 2
58 1 9 15 2 10 9 10 9 13 7 2 10 9 13 9 1 10 3 7 10 0 9 1 10 9 7 10 9 10 9 2 7 13 7 2 10 9 15 14 13 10 9 1 9 10 9 15 1 0 9 7 14 13 10 9 15 2 2
28 10 9 13 13 1 9 1 2 7 1 2 14 13 10 0 9 15 7 0 9 15 1 10 9 9 1 9 2
37 1 10 9 9 15 2 15 13 1 9 10 9 2 10 9 9 13 3 9 1 2 0 9 2 2 1 10 9 0 0 7 0 9 1 10 0 2
15 3 2 10 9 13 10 0 9 1 10 0 9 10 9 2
16 10 9 1 0 9 7 9 13 3 13 1 10 9 9 2 2
16 13 10 9 10 9 2 10 9 13 14 13 10 0 9 9 2
21 1 10 0 9 2 10 9 9 13 1 9 10 9 2 3 3 13 12 0 9 2
2 12 2
15 15 13 7 13 14 13 10 9 15 7 13 10 0 9 2
27 7 13 3 1 9 1 9 2 10 9 10 9 14 13 0 14 13 1 10 9 7 10 9 9 10 9 2
31 1 12 9 2 10 9 10 9 9 2 9 9 2 13 10 9 9 10 9 2 7 10 9 13 14 13 10 9 1 9 2
27 10 9 2 10 15 13 10 9 10 9 9 7 13 10 9 10 0 2 13 1 9 12 9 7 12 9 2
18 13 3 0 14 13 3 15 10 9 7 14 13 10 9 1 10 9 2
32 10 9 10 9 2 10 15 13 1 0 9 15 13 0 1 0 9 1 10 9 7 10 9 2 13 14 13 10 9 0 9 2
9 2 10 15 13 14 13 3 9 2
24 1 14 13 9 1 0 9 15 10 9 2 13 7 10 0 9 14 13 14 13 3 1 9 2
8 10 0 9 10 9 1 9 2
28 3 1 10 0 9 13 7 10 9 10 9 1 9 1 10 9 15 13 1 10 9 9 1 10 0 0 9 2
26 10 9 10 9 15 13 1 0 9 15 13 7 10 0 9 3 13 0 9 9 1 7 10 0 9 2
30 1 10 9 15 2 13 3 0 10 9 15 13 15 10 9 7 15 13 10 9 0 9 2 10 9 7 10 0 9 2
17 10 9 10 9 1 9 15 13 3 10 0 2 7 10 9 13 2
72 3 0 13 10 9 7 3 1 10 13 9 9 15 13 3 1 15 9 1 10 9 10 9 10 9 14 13 7 10 0 9 0 9 1 10 0 9 3 2 1 15 2 14 13 10 9 1 10 9 2 10 9 1 10 9 10 9 2 10 0 9 2 3 7 10 9 1 10 9 10 9 2
29 10 9 3 1 10 0 9 10 9 1 9 1 9 3 9 7 1 9 1 9 9 14 13 3 0 1 10 9 2
27 7 1 10 12 2 10 9 13 1 10 12 2 14 13 0 0 9 2 10 9 10 9 14 13 14 13 2
21 10 9 13 1 10 0 0 9 2 10 0 9 2 10 0 9 7 10 0 9 2
39 10 9 15 13 0 7 0 10 0 9 7 13 1 9 15 10 9 2 3 7 10 0 9 14 13 0 7 13 7 10 0 9 2 10 9 7 10 9 2
30 10 9 15 14 13 1 10 9 0 9 2 7 10 0 9 15 13 0 2 0 9 1 9 0 9 1 10 13 9 2
28 3 1 10 9 9 0 9 2 13 7 0 9 1 0 9 2 7 10 9 10 9 13 1 0 9 1 9 2
27 10 9 10 9 10 9 2 9 9 2 10 15 13 13 1 10 9 0 9 2 13 0 1 9 0 9 2
11 10 9 10 0 9 13 1 15 10 9 2
34 3 2 10 9 9 13 10 9 9 10 9 2 0 1 10 0 9 3 10 9 9 3 7 10 9 9 2 1 14 13 1 15 9 2
27 13 7 7 2 10 0 9 13 13 9 10 15 13 2 7 14 13 0 2 3 13 2 10 9 14 13 2
21 14 13 14 13 0 14 13 14 13 12 9 7 14 13 1 10 9 1 0 9 2
8 9 13 1 9 1 0 9 2
12 1 2 10 15 14 13 14 13 10 9 15 2
28 1 10 9 15 10 9 13 14 13 1 0 9 7 13 1 0 9 14 13 1 3 13 14 13 9 1 9 2
27 3 13 10 9 2 10 0 9 9 12 2 2 7 13 10 9 1 10 9 1 10 9 1 12 9 3 2
36 10 9 10 9 10 2 7 10 9 10 0 9 1 10 2 7 10 0 9 13 10 9 15 13 10 0 9 2 1 10 9 9 1 10 9 2
31 10 9 15 13 14 13 3 0 9 7 3 1 9 9 1 10 0 9 7 10 0 9 2 10 9 3 13 10 9 9 2
7 1 10 9 13 12 9 2
11 10 9 13 13 3 2 3 1 12 9 2
21 1 13 0 1 10 0 9 2 1 15 13 7 0 0 2 3 0 1 12 2 2
28 7 15 13 10 0 9 1 10 0 9 2 7 10 0 9 2 3 10 0 9 10 9 3 15 13 14 13 2
13 10 9 14 13 10 9 1 10 9 10 0 9 2
20 15 13 3 7 2 1 15 10 9 2 9 1 10 9 15 13 13 1 9 2
3 2 9 2
41 10 9 13 1 0 2 1 3 2 9 15 1 10 9 10 9 2 9 9 9 2 13 7 2 13 13 3 0 9 1 10 14 13 10 9 15 13 10 9 2 2
16 7 2 1 9 10 9 7 10 9 13 13 0 3 0 9 2
31 10 9 10 12 9 10 9 10 9 10 9 1 9 13 15 10 9 2 10 15 13 3 1 9 10 9 0 9 10 9 2
23 1 9 2 10 0 9 2 3 1 9 13 9 10 9 14 13 10 9 15 10 0 9 2
23 1 9 2 1 10 0 9 13 12 1 12 9 1 10 9 10 9 1 10 9 10 9 2
35 10 9 9 9 10 9 2 9 9 2 13 1 9 9 1 15 13 0 9 1 10 9 1 10 0 9 10 0 9 1 10 9 10 9 2
26 10 9 9 13 13 0 1 10 9 1 10 12 0 9 7 13 14 13 3 9 1 9 9 10 9 2
12 15 13 14 13 2 10 9 2 14 10 9 2
48 15 13 10 9 15 1 10 12 9 3 10 9 7 13 3 1 10 0 9 14 15 13 10 0 9 1 3 10 9 2 7 13 14 13 10 9 15 13 10 9 1 9 1 10 9 10 9 2
34 1 10 0 9 15 13 10 9 10 2 9 9 2 2 10 9 9 2 9 2 13 0 1 10 9 1 9 9 15 13 1 10 9 2
20 13 3 14 13 9 15 3 14 13 7 3 1 10 0 9 7 10 9 15 2
7 13 14 13 10 0 9 2
17 14 13 7 1 10 9 15 14 13 10 0 9 3 0 1 9 2
5 9 9 1 0 9
28 1 10 0 9 1 10 9 1 9 13 10 12 0 9 2 10 15 1 10 9 13 1 9 1 9 1 9 2
11 7 2 13 3 3 3 1 10 15 9 2
11 13 3 1 0 0 9 1 9 10 9 2
39 9 15 13 1 10 9 15 13 10 9 10 9 10 9 10 9 1 9 2 13 1 9 10 9 12 1 12 9 1 10 0 9 7 10 9 10 0 9 2
41 10 0 9 0 9 7 0 9 2 3 7 13 10 9 9 1 10 9 10 9 2 15 13 10 9 13 0 1 9 7 10 9 15 13 1 9 13 0 7 0 2
19 15 7 10 9 13 1 10 9 7 13 10 0 9 10 9 15 1 9 2
40 10 9 10 9 13 9 10 0 9 15 13 10 9 7 3 1 10 15 10 9 13 10 9 14 13 3 10 0 9 2 3 1 10 9 10 0 9 7 9 2
13 10 9 13 10 9 10 0 9 7 13 1 9 2
51 10 9 2 13 9 2 1 10 9 9 7 10 9 9 13 10 0 9 1 9 10 9 2 10 0 9 10 9 15 3 13 13 0 2 13 1 0 9 3 1 0 9 7 13 10 0 9 1 10 9 2
32 15 13 3 0 3 3 1 9 9 15 13 10 0 9 9 7 10 0 9 10 0 9 1 10 9 2 10 9 10 0 9 2
5 15 13 10 9 2
32 1 10 2 3 13 13 2 0 9 2 10 9 13 3 0 0 9 2 9 9 2 7 1 9 9 1 10 9 9 10 9 2
9 1 15 2 13 3 10 9 15 2
36 3 2 10 9 9 13 13 7 2 10 9 9 13 3 1 10 9 10 9 15 1 9 2 10 15 13 10 9 0 9 1 10 9 15 2 2
22 12 9 1 10 9 10 0 9 10 9 2 10 9 13 1 12 9 1 9 10 9 2
44 1 10 15 2 10 9 9 13 7 2 10 9 15 14 13 10 9 10 12 13 10 9 10 9 7 10 15 12 0 9 7 10 9 0 10 0 9 1 9 7 1 9 2 2
20 13 7 10 2 9 14 13 14 15 13 1 9 15 7 1 0 9 10 9 2
13 14 13 0 1 10 9 9 10 9 10 9 15 2
32 10 9 14 13 0 7 10 9 13 9 1 9 14 13 0 9 3 1 10 0 9 2 10 15 7 13 1 9 1 0 9 2
32 1 10 9 15 2 14 13 10 0 9 2 10 15 1 3 13 13 10 9 10 9 10 9 9 2 14 13 10 12 1 12 2
29 3 2 3 1 10 9 10 9 1 9 2 1 0 10 0 9 13 0 7 10 9 9 14 13 1 0 9 9 2
32 1 9 2 1 10 9 9 1 9 2 9 10 0 9 10 9 2 7 9 2 12 9 13 10 9 15 2 7 15 12 13 2
11 13 0 7 0 9 2 0 1 10 9 2
27 1 9 10 9 2 10 9 13 10 9 7 10 9 2 13 3 10 9 10 9 2 7 7 0 10 9 2
16 10 0 9 2 10 15 13 1 10 0 10 0 9 13 9 2
40 10 9 13 3 7 13 10 9 1 9 2 1 15 13 10 0 9 10 9 1 9 3 10 2 2 7 13 3 3 10 9 10 9 15 13 13 1 15 9 2
35 1 9 2 10 9 9 13 1 9 9 3 13 9 1 10 9 9 10 2 2 9 9 2 9 15 13 10 0 9 1 10 9 10 9 2
18 10 9 12 2 9 1 10 9 2 13 9 9 9 7 10 9 9 2
20 10 0 9 15 13 13 1 9 1 10 9 1 0 9 13 3 0 9 2 2
26 10 0 9 10 0 9 13 10 9 10 9 9 2 10 15 13 1 2 1 9 9 2 0 9 2 2
9 13 10 9 10 9 10 9 9 2
28 3 2 10 9 13 10 9 0 9 1 9 12 2 1 10 9 10 0 9 1 9 10 12 10 9 9 12 2
39 10 0 9 9 13 13 10 0 9 2 10 0 9 10 15 2 1 10 9 0 0 7 0 9 1 0 15 10 9 2 13 14 15 13 7 14 15 13 2
29 1 0 9 1 9 10 9 13 7 3 7 10 9 0 9 14 13 14 13 3 9 14 13 3 3 10 0 9 2
26 1 10 9 14 13 10 15 14 13 0 10 9 1 10 9 1 10 9 10 9 2 13 10 2 9 2
23 10 9 10 9 15 13 10 13 9 10 0 9 10 9 2 14 13 1 0 10 0 9 2
14 10 0 9 13 14 13 10 9 15 3 1 0 9 2
13 15 13 14 13 1 9 7 14 13 10 9 15 2
11 13 3 0 9 10 9 3 13 10 9 2
29 10 0 9 2 10 0 9 13 9 1 9 1 9 1 0 15 13 3 9 10 9 1 0 0 9 1 10 9 2
12 1 9 15 13 10 9 10 0 0 9 9 2
42 3 2 1 9 10 9 10 9 2 15 13 10 9 10 9 14 13 3 15 9 1 9 10 0 15 9 3 13 3 1 0 9 10 9 15 13 1 10 0 0 9 2
38 1 14 13 10 9 14 13 3 10 9 15 2 7 15 13 1 9 2 10 0 13 14 13 1 10 9 10 9 10 9 10 9 15 13 3 10 9 2
14 10 9 10 9 14 13 13 10 0 9 10 9 9 2
3 2 9 2
43 13 2 10 9 2 10 2 9 2 1 9 10 9 2 3 1 9 10 2 7 10 9 15 13 0 1 3 13 0 9 1 10 9 10 9 9 7 13 10 9 0 9 2
26 10 9 2 0 3 2 9 10 9 2 2 13 10 9 3 2 10 12 0 9 1 10 0 9 2 2
37 1 10 9 15 13 13 7 10 0 9 7 10 0 9 13 1 9 7 13 0 10 0 15 9 2 7 9 10 9 9 2 7 14 15 10 9 2
18 3 2 10 9 9 13 10 9 15 1 10 9 7 14 13 0 9 2
34 10 0 9 15 14 13 14 13 7 0 10 9 14 13 0 1 0 15 7 7 2 7 13 2 14 13 10 9 7 10 9 1 9 2
21 0 7 0 9 1 10 9 13 1 0 9 2 12 1 10 3 0 9 10 9 2
40 7 0 9 9 14 13 10 9 15 13 1 10 9 2 10 2 13 14 13 1 9 14 13 13 9 10 15 14 13 10 9 10 9 2 3 13 3 1 9 2
39 1 10 9 10 9 9 9 13 0 9 1 10 9 15 2 7 1 10 9 10 9 10 9 13 13 7 14 13 0 10 9 15 13 13 10 9 10 9 2
29 1 3 1 9 13 0 9 7 9 9 2 7 10 0 9 2 10 9 10 9 2 14 13 3 7 14 13 3 2
11 10 9 13 9 3 1 9 10 0 9 2
47 15 9 13 7 2 10 9 13 1 9 10 0 2 10 15 13 1 9 9 7 9 12 9 9 2 2 7 15 13 7 2 10 9 13 14 13 3 9 10 9 15 13 1 0 9 2 2
13 10 9 10 9 13 12 1 10 12 0 10 9 2
38 10 9 1 10 9 9 13 14 13 7 0 10 9 7 0 10 9 13 3 2 3 7 1 0 9 13 15 13 9 2 3 15 15 13 1 9 9 2
23 1 9 2 13 0 1 10 9 9 14 13 1 0 9 7 14 13 10 9 10 0 9 2
33 1 9 1 10 0 2 10 9 13 3 10 0 9 7 1 10 9 15 10 9 10 0 9 1 10 0 9 13 3 10 0 9 2
33 1 10 9 15 10 2 13 1 10 9 2 3 1 12 9 15 2 15 1 15 2 3 1 10 3 0 9 9 9 2 13 9 2
1 9
21 13 10 9 10 0 14 13 1 14 13 14 13 3 10 9 9 1 9 10 9 2
2 12 2
10 10 9 15 14 13 13 1 15 15 2
12 13 3 7 10 9 10 9 13 1 0 9 2
27 3 3 1 9 1 10 9 14 13 14 13 7 0 10 9 1 9 14 13 0 9 14 13 9 1 9 2
35 3 1 10 9 10 9 1 0 9 7 9 13 0 1 10 0 9 15 13 1 10 9 10 0 9 10 0 9 1 9 10 9 10 12 2
52 13 1 15 10 15 13 1 10 9 15 10 9 2 7 10 9 15 9 13 1 10 9 10 9 2 10 0 15 2 9 1 10 9 15 13 13 10 12 0 9 7 14 13 3 10 9 14 13 13 0 9 2
34 10 0 9 1 0 9 2 1 9 0 1 10 9 10 2 2 13 7 10 9 13 3 7 0 9 1 9 3 3 13 1 0 9 2
17 1 0 9 10 9 10 0 9 2 13 7 10 9 13 12 9 2
4 2 2 1 2
23 13 0 7 13 10 0 9 9 10 9 7 10 0 9 0 0 9 7 9 10 9 9 2
26 1 15 9 10 9 13 1 0 9 2 15 9 13 10 12 9 2 7 10 9 15 13 10 12 9 2
13 15 13 10 9 15 13 1 9 1 10 9 9 2
28 10 9 13 3 0 7 0 1 12 9 2 1 9 14 13 10 9 1 12 9 10 9 2 3 1 9 9 2
11 1 15 10 9 13 15 10 9 10 9 2
29 1 0 9 2 1 9 10 9 13 7 10 12 13 2 15 15 13 3 10 9 1 9 1 10 0 9 9 9 2
49 3 3 13 10 9 10 9 2 2 1 9 15 2 15 13 10 0 9 10 9 2 14 14 13 14 13 10 9 1 12 9 2 7 15 13 1 15 13 14 15 13 7 1 9 15 15 13 2 2
23 10 0 9 3 13 10 9 3 1 10 12 15 9 1 3 0 9 0 9 7 0 9 2
13 10 9 13 7 1 10 0 9 10 0 9 15 2
6 15 13 10 0 9 2
44 1 9 13 9 1 9 2 9 10 0 9 2 2 3 1 10 9 10 0 9 2 15 13 13 1 9 10 9 2 10 9 13 1 9 10 0 9 15 1 10 9 10 9 2
19 10 0 9 13 14 13 2 7 10 9 7 10 9 13 9 1 0 9 2
13 10 9 13 1 10 9 15 13 0 1 9 9 2
26 10 9 9 13 7 10 9 2 15 14 13 1 1 15 9 2 13 0 9 1 10 9 10 0 9 2
2 12 2
8 13 0 7 13 13 12 9 2
11 10 0 9 3 1 10 9 7 10 9 2
36 1 9 15 2 13 7 10 9 14 13 10 9 7 14 13 10 9 7 10 9 14 13 14 13 15 10 9 9 1 10 9 9 10 0 9 2
17 3 2 13 15 10 9 7 3 1 0 9 2 13 1 0 9 2
18 10 12 9 13 9 10 9 10 0 9 15 13 10 0 9 0 9 2
105 1 0 7 9 10 0 9 13 1 0 9 2 3 3 13 10 9 9 1 10 0 9 1 9 2 9 7 1 10 9 0 9 2 10 9 12 10 15 14 13 14 13 2 3 7 14 13 3 0 14 13 3 10 9 1 9 10 0 9 2 7 1 12 9 2 3 1 9 9 1 10 0 9 1 9 10 9 2 10 9 7 10 9 2 14 13 10 0 9 10 9 12 2 10 15 13 0 1 10 9 12 10 12 9 2
17 10 9 13 1 0 9 10 9 2 13 10 0 7 0 15 9 2
1 9
55 13 14 13 1 9 15 1 10 0 12 7 12 9 7 10 9 9 10 9 14 13 1 10 9 7 10 9 10 0 9 2 7 13 2 7 14 13 1 15 3 2 1 14 13 1 9 14 13 13 10 9 1 10 9 2
44 15 13 1 7 10 9 10 9 13 3 0 7 10 0 0 9 13 7 10 14 13 15 10 9 15 1 15 9 9 13 0 9 7 10 0 9 7 14 13 0 10 15 9 2
6 13 0 9 10 9 2
17 7 2 10 9 13 3 7 13 14 13 1 10 9 1 12 9 2
13 1 10 9 15 2 10 9 13 9 1 9 9 2
35 10 9 2 10 15 3 13 13 0 0 9 13 14 3 1 9 1 0 15 9 7 1 9 1 0 9 15 7 1 9 1 0 9 15 2
30 13 14 13 10 9 15 2 3 1 10 9 10 9 7 1 9 1 10 0 9 2 9 1 9 2 14 13 3 2 2
32 1 10 9 15 13 2 3 1 0 15 0 9 15 13 3 1 9 13 2 10 0 9 1 15 14 13 14 13 1 10 9 2
20 2 13 9 14 13 2 1 9 0 9 7 10 9 9 15 14 13 0 9 2
2 15 2
14 1 15 10 0 13 0 7 10 0 14 13 9 9 2
19 10 0 0 9 13 1 15 10 0 2 0 7 0 9 1 9 10 9 2
17 10 0 0 9 10 9 13 12 9 2 12 1 15 9 10 9 2
46 10 12 9 9 3 1 10 9 9 14 13 3 14 13 1 0 7 0 9 2 3 7 1 0 9 14 13 9 7 9 1 15 9 7 10 9 1 9 14 13 3 10 0 3 13 2
24 7 3 10 0 9 10 9 15 13 14 13 3 7 10 9 3 1 10 9 14 13 3 0 2
8 10 0 9 13 13 10 0 9
71 7 2 0 1 15 1 15 10 9 13 7 10 9 10 0 9 14 14 13 10 3 9 10 9 2 7 1 15 10 9 3 13 0 9 14 13 10 0 9 15 13 2 14 3 1 0 9 1 10 9 10 9 10 9 2 7 3 2 14 13 1 2 9 2 1 9 10 0 9 10 2
31 1 10 9 2 1 10 0 9 13 3 10 9 2 13 9 9 10 0 9 10 9 1 12 0 2 9 9 2 10 9 2
35 13 10 0 9 15 14 13 7 10 0 9 7 9 14 14 13 14 13 3 3 1 10 9 10 0 9 0 9 2 10 15 13 10 9 2
26 10 9 9 13 1 10 9 9 1 9 12 2 1 9 10 0 9 10 9 10 12 10 9 9 12 2
32 3 2 10 9 3 1 10 9 2 3 3 7 10 9 10 9 2 13 13 0 9 2 2 13 10 9 9 2 9 10 9 2
10 13 7 10 9 13 13 10 9 9 2
22 3 2 10 9 2 10 9 7 10 9 13 1 2 7 10 9 13 7 1 10 9 2
38 10 9 15 1 0 10 9 13 14 13 1 9 10 0 9 7 14 13 10 9 14 13 1 9 7 14 13 0 9 9 7 9 1 9 1 0 9 2
23 3 2 10 0 9 10 9 13 2 3 1 15 15 2 10 9 15 13 14 13 1 9 2
30 3 2 10 9 13 10 9 14 13 10 0 9 1 9 10 9 0 9 2 15 13 1 9 1 10 9 1 10 9 2
1 9
21 3 10 0 9 13 15 12 12 9 2 1 9 9 15 13 13 1 10 0 9 2
28 3 14 15 13 3 7 14 15 13 2 7 3 3 13 1 0 9 14 15 13 10 9 15 7 10 9 15 2
5 1 9 10 9 2
12 3 1 10 9 2 13 7 10 9 10 9 2
14 10 12 9 10 0 9 15 13 10 3 0 0 9 2
35 10 9 10 9 2 10 15 13 3 7 9 10 9 15 2 7 3 13 1 12 9 2 13 3 1 9 10 9 2 7 13 14 13 3 2
46 13 3 15 10 9 15 9 1 9 0 9 7 10 0 9 15 13 10 9 9 2 10 15 13 9 1 9 15 7 13 2 3 2 1 10 9 15 2 13 14 13 1 9 10 9 2
9 15 13 10 0 9 10 9 15 2
31 15 14 13 0 10 9 7 1 10 9 15 13 9 14 3 1 9 2 7 3 1 9 9 13 7 13 14 13 10 9 2
26 10 9 13 7 14 13 0 10 0 0 9 1 0 9 7 1 15 13 3 14 13 1 0 9 15 2
20 1 10 9 15 10 9 13 0 9 1 10 9 10 9 1 9 1 9 9 2
31 9 9 2 1 3 1 10 9 15 1 9 9 10 9 2 3 1 10 9 7 10 9 10 9 2 13 14 13 10 9 2
9 14 13 14 13 7 10 0 9 2
71 1 10 9 15 10 9 10 2 2 9 9 2 13 14 13 10 9 2 13 7 10 9 1 10 12 9 14 13 10 0 9 1 9 2 7 10 9 10 12 9 1 9 0 9 2 9 7 9 2 7 10 9 14 13 14 13 3 1 10 9 1 9 2 0 10 0 9 7 10 9 2
10 15 13 3 10 0 9 10 0 9 2
17 10 9 9 10 2 13 1 10 2 7 10 2 1 9 0 9 2
16 10 9 1 10 2 13 7 10 9 15 13 1 9 1 9 2
25 13 7 1 0 9 2 10 2 9 9 13 10 0 9 2 10 0 9 10 0 9 13 3 0 2
18 1 9 13 9 1 10 9 9 2 7 10 9 1 10 9 13 0 2
24 10 9 10 9 9 9 13 2 13 10 3 0 0 9 1 9 15 3 7 3 0 9 2 2
9 2 2 0 9 1 10 0 9 2
18 10 9 10 0 9 10 9 1 9 10 0 0 9 14 13 0 9 2
4 0 9 1 9
8 3 1 10 0 9 9 9 2
35 13 13 1 10 9 15 13 10 9 3 1 10 9 15 13 13 10 0 9 2 3 7 7 13 3 10 9 10 15 13 13 10 0 9 2
20 1 10 9 2 9 13 9 7 0 9 1 0 9 1 0 10 9 10 9 2
23 13 10 0 9 14 13 9 1 10 0 2 0 9 7 14 13 9 10 9 10 9 15 2
22 1 0 9 10 0 9 13 0 3 9 1 9 1 10 0 9 1 9 10 9 9 2
17 13 1 10 9 9 2 9 9 9 9 2 1 10 9 10 9 2
12 10 9 12 13 7 10 9 13 1 0 9 2
17 13 7 10 9 3 1 10 9 10 9 1 10 9 10 0 13 2
48 3 2 1 14 13 10 0 9 14 13 3 10 3 3 1 9 10 9 2 13 14 13 14 13 10 0 0 9 7 0 0 9 15 2 3 7 10 9 15 1 9 15 13 10 9 10 9 2
29 1 10 0 9 13 7 13 1 10 9 15 10 9 3 7 7 13 9 10 9 2 7 13 7 10 9 10 9 2
21 10 9 14 13 14 13 1 9 7 1 12 0 2 3 10 9 7 10 12 9 2
34 3 7 1 2 10 0 9 15 13 13 10 0 9 1 9 12 10 9 13 13 7 10 9 10 2 14 13 9 9 10 0 9 9 2
14 1 9 10 0 9 13 10 0 0 9 1 10 9 2
21 14 13 9 7 13 10 0 0 9 9 7 10 0 2 13 14 13 15 10 9 2
10 10 0 15 9 13 14 13 10 9 2
28 13 0 14 13 10 9 7 7 10 12 9 13 3 10 9 15 7 13 15 15 10 0 13 9 1 9 9 2
19 3 2 3 0 9 2 1 10 9 1 10 9 2 14 13 0 1 9 2
39 10 9 15 13 7 10 0 9 15 13 1 9 2 1 10 9 10 9 15 2 2 9 2 13 1 9 14 13 0 0 9 7 3 13 10 9 1 9 2
6 9 13 10 9 9 2
35 10 9 12 13 10 9 1 9 10 9 2 10 9 12 10 9 9 15 13 10 9 10 0 9 7 13 1 9 1 10 9 9 7 9 2
5 13 3 12 9 2
4 0 9 1 9
17 14 13 14 13 1 0 1 10 9 15 13 1 9 1 10 9 2
9 3 2 13 7 1 10 0 9 2
44 13 10 9 1 10 2 9 2 7 14 1 10 2 9 2 1 0 9 0 9 1 9 9 7 9 10 9 1 10 0 9 2 1 9 10 9 10 9 9 12 10 0 9 2
40 10 9 15 13 10 9 15 1 10 9 10 9 10 9 2 9 10 9 15 1 10 9 2 13 1 0 9 10 9 7 13 1 10 9 3 1 10 9 9 2
34 10 9 9 9 13 1 9 1 10 9 10 9 9 9 2 7 13 1 10 0 0 9 1 9 1 10 9 10 9 10 12 7 12 2
20 10 15 9 2 15 13 1 12 0 9 1 10 9 2 13 7 14 13 0 2
37 14 15 13 3 2 14 15 13 1 9 15 7 1 15 15 15 10 0 13 14 13 2 7 14 13 7 13 14 13 3 7 3 1 15 10 9 2
12 10 9 9 10 9 14 13 7 14 13 0 2
25 10 9 13 9 7 9 1 14 13 1 12 10 9 2 1 10 9 14 13 9 1 9 12 9 2
19 10 9 13 13 1 0 9 2 3 10 12 10 9 13 1 10 0 9 2
15 9 10 9 14 13 10 12 9 0 15 9 7 9 9 2
16 7 13 3 0 14 13 15 3 1 9 3 1 10 0 9 2
17 1 9 15 2 10 9 10 0 7 0 9 9 13 0 7 0 2
10 10 0 9 13 3 14 15 13 3 2
17 2 1 3 13 10 9 1 0 9 7 14 13 3 10 9 15 2
52 7 10 9 13 9 2 13 1 9 10 9 10 9 2 3 10 9 13 3 9 10 9 7 13 10 9 10 9 15 2 10 15 13 1 9 15 0 1 10 9 10 9 2 9 2 7 10 9 2 9 2 2
14 1 7 10 9 15 2 13 1 9 2 13 7 9 2
24 15 13 7 13 7 1 10 0 7 0 9 1 0 2 0 7 0 9 7 9 1 10 9 2
18 13 1 9 10 9 10 9 15 7 1 9 10 0 9 1 10 9 2
22 3 15 10 9 10 0 9 7 9 13 10 9 10 9 15 1 9 9 10 9 9 2
27 1 10 9 13 10 9 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 7 0 7 0 9 2
5 13 3 3 15 2
35 3 15 10 9 13 14 13 10 12 0 7 3 7 10 12 0 2 1 9 10 9 0 9 2 9 10 15 10 9 13 3 7 1 10 2
3 2 9 2
27 3 2 10 9 15 13 14 13 7 10 0 9 3 13 10 9 10 9 2 1 14 15 13 3 0 9 2
27 14 14 13 3 1 0 9 10 9 10 9 9 1 10 0 15 9 7 14 13 0 10 9 10 0 9 2
14 13 0 9 3 1 10 9 9 1 10 9 10 9 2
13 1 10 9 15 2 13 14 13 10 9 1 9 2
26 1 9 10 15 14 13 14 13 13 1 10 9 14 13 9 9 2 7 2 1 15 13 2 9 0 2
14 10 2 9 9 13 10 9 15 13 14 13 7 15 2
34 3 14 13 7 14 15 13 1 9 7 3 7 0 9 13 14 13 7 13 13 3 10 9 10 9 15 13 10 2 1 0 9 3 2
14 1 10 13 9 10 9 2 10 9 9 13 1 9 2
19 0 9 13 7 10 9 1 0 10 9 2 10 15 13 0 1 9 9 2
30 9 9 1 10 0 9 7 0 9 13 7 2 1 10 9 13 12 9 7 10 9 13 1 9 2 9 7 9 2 2
28 10 0 9 2 13 3 0 2 7 13 1 10 9 10 9 1 10 12 9 10 9 9 1 0 9 10 12 2
19 13 7 10 9 15 10 9 14 13 9 10 2 2 14 13 7 14 13 2
18 1 15 10 9 2 10 9 13 3 1 9 14 13 1 10 9 15 2
27 1 9 2 13 13 0 1 12 0 9 1 10 9 2 7 9 13 13 1 12 1 10 12 9 7 9 2
30 2 10 0 9 13 10 0 9 15 2 13 0 9 1 9 7 13 3 1 10 9 10 0 9 2 13 10 9 9 2
21 3 2 1 10 9 15 2 13 14 13 10 9 9 1 9 9 0 10 12 9 2
7 2 1 3 13 0 9 2
6 1 0 9 10 9 2
20 10 9 2 1 10 9 10 9 13 1 0 9 2 10 15 13 3 12 9 2
21 10 9 2 10 9 7 10 0 9 13 14 13 1 9 3 1 10 9 1 9 2
22 3 13 10 0 9 1 9 1 10 9 2 10 15 13 1 0 9 1 9 10 9 2
16 13 7 10 9 15 13 0 7 13 10 9 14 14 15 13 2
39 3 3 1 10 9 10 9 7 10 9 10 9 7 9 10 9 1 10 9 13 0 10 0 9 14 13 7 10 9 13 9 15 15 13 1 9 10 9 2
29 13 9 1 14 13 10 9 15 7 13 14 13 10 9 1 10 9 7 10 9 3 3 7 14 13 9 1 9 2
39 7 7 14 13 14 13 10 9 2 10 9 10 9 1 10 9 7 10 9 13 3 13 7 2 3 3 3 2 13 13 7 13 10 9 14 13 0 9 2
26 10 0 9 10 9 2 10 9 13 9 1 10 0 9 2 10 15 13 0 10 9 15 13 1 9 2
24 3 13 10 0 9 2 13 10 9 7 10 0 9 2 13 1 10 9 3 2 1 0 9 2
28 10 9 13 10 9 1 10 9 9 15 13 10 9 1 9 9 0 0 2 10 15 1 9 13 1 0 9 2
1 9
28 10 0 7 0 9 13 1 10 0 0 9 1 10 9 10 9 7 10 9 15 1 0 9 1 3 0 9 2
21 3 2 13 12 9 2 1 10 15 10 12 13 7 13 1 9 1 10 9 15 2
17 0 10 9 13 3 9 10 9 9 2 7 12 1 15 13 9 2
31 10 9 7 10 9 2 7 14 13 14 13 7 13 1 0 9 2 13 1 10 9 10 0 9 2 10 15 13 3 0 2
6 1 9 10 9 9 2
28 1 10 9 15 2 10 0 9 13 1 10 0 9 14 13 10 0 9 10 0 0 9 2 3 7 3 9 2
9 13 7 13 3 14 15 13 15 2
18 13 9 1 15 13 12 9 1 0 9 2 10 9 7 10 12 9 2
41 10 9 15 13 3 1 10 9 10 2 9 9 7 14 13 14 13 10 0 9 9 9 1 0 0 9 2 7 13 0 14 13 3 0 9 9 9 1 0 9 2
37 1 9 10 9 13 1 10 9 2 13 7 13 1 10 0 9 7 13 14 13 7 7 10 9 13 10 9 15 1 9 2 14 13 1 9 15 2
12 1 0 9 2 13 0 1 10 9 10 9 2
30 1 15 15 13 10 9 14 13 1 10 0 9 1 15 13 10 0 9 1 9 7 10 0 9 1 9 10 0 9 2
36 10 9 14 13 9 1 9 7 1 9 1 10 9 0 0 0 9 15 14 13 1 9 1 9 10 9 10 15 13 14 13 1 9 10 9 2
23 9 13 3 10 9 1 9 10 9 9 2 7 1 9 10 9 10 9 15 13 3 0 2
17 15 13 10 9 9 2 7 15 14 15 13 7 15 15 13 3 2
42 13 3 14 13 10 9 7 0 10 9 9 1 10 9 15 1 15 15 1 12 9 13 10 3 0 9 2 7 7 13 15 1 9 7 1 9 15 2 13 3 0 2
14 10 9 10 9 1 9 13 10 9 15 13 3 0 2
38 10 9 15 10 9 14 13 7 3 14 13 3 3 10 9 10 9 2 1 10 9 1 9 2 2 10 9 0 9 2 10 9 9 7 10 0 9 2
18 15 10 9 1 10 15 10 9 14 13 10 9 13 10 0 9 9 2
18 10 9 13 1 10 9 7 1 9 13 1 0 9 1 9 0 9 2
47 1 0 9 2 13 0 7 15 15 13 3 13 9 3 0 9 7 13 10 13 9 9 2 7 13 14 13 3 9 7 7 1 15 13 0 7 0 9 2 3 14 15 13 3 3 3 2
42 3 2 10 9 10 9 3 1 10 9 0 9 1 0 9 2 10 15 3 14 13 0 1 10 9 15 2 14 13 13 3 1 9 2 12 9 3 1 10 9 15 2
24 3 13 10 0 9 10 9 7 10 9 10 9 15 2 13 13 14 13 7 13 13 0 9 2
19 1 9 13 9 0 0 9 2 3 9 2 9 2 9 7 15 0 9 2
7 3 14 13 14 13 3 2
19 10 15 15 13 2 7 13 7 13 10 9 15 14 13 3 0 7 0 2
51 3 1 10 9 2 10 0 9 13 7 13 1 0 9 7 7 13 15 1 9 2 1 9 14 13 0 2 14 13 7 13 14 13 0 9 3 0 9 2 13 3 1 10 9 14 13 3 1 10 9 2
39 7 13 3 1 9 2 3 13 3 2 13 10 9 1 14 13 10 9 15 7 14 13 3 10 9 15 2 2 13 10 9 9 2 9 9 1 10 9 2
36 3 1 9 2 10 9 13 10 0 9 2 13 10 9 2 1 10 9 7 1 9 1 10 9 7 3 1 10 9 2 3 13 9 10 9 2
44 10 9 13 9 10 9 1 10 9 10 9 2 12 9 2 3 13 10 9 15 9 9 9 2 9 10 0 9 1 10 9 10 9 7 10 9 2 9 2 15 13 10 9 2
36 10 9 9 3 13 7 13 14 13 1 9 2 13 0 0 9 2 3 1 0 0 9 2 3 10 9 10 9 15 7 13 1 0 15 9 2
12 9 1 10 9 10 0 9 13 10 9 9 2
6 14 14 13 14 13 2
90 10 9 15 10 9 9 2 10 15 10 9 13 2 13 10 0 0 9 1 14 13 10 0 9 2 10 15 13 0 9 3 1 10 9 10 9 3 1 10 9 10 9 7 10 0 9 9 2 14 13 3 2 1 10 9 2 7 10 12 0 9 2 10 15 13 14 13 9 9 1 9 9 7 0 9 1 12 7 9 7 10 15 13 3 1 0 9 10 9 2
36 14 13 3 14 13 14 13 0 10 12 9 10 9 1 10 9 1 9 2 1 9 9 7 1 9 2 9 15 14 13 0 9 1 0 9 2
32 10 9 2 3 1 9 2 10 9 7 10 9 2 13 12 1 10 0 9 10 9 2 1 15 13 9 0 9 9 7 9 2
32 13 1 10 0 9 3 1 10 0 9 2 3 7 10 9 3 13 0 10 9 1 10 0 9 2 7 13 1 9 7 13 2
17 7 7 13 2 10 9 13 10 9 1 10 0 9 10 9 9 2
28 10 0 9 2 12 9 10 9 13 13 1 10 9 7 10 0 9 2 7 9 13 13 7 1 0 0 9 2
32 3 1 10 9 2 2 10 9 9 13 14 13 10 9 10 0 9 10 2 2 7 10 9 9 13 14 13 9 1 9 2 2
13 7 13 1 10 9 15 2 13 10 9 1 9 2
91 1 15 10 9 2 1 10 15 10 12 13 9 9 2 2 7 13 3 10 2 9 3 7 10 2 9 2 7 10 12 13 3 1 10 2 9 2 10 0 9 13 10 9 10 0 9 10 1 9 12 9 2 7 14 15 13 0 9 0 9 2 14 15 13 10 9 1 0 9 7 9 1 9 15 7 10 9 1 0 9 2 3 7 14 15 13 3 10 9 9 2
11 10 9 9 13 0 1 9 1 10 12 2
19 1 10 9 15 2 13 1 10 9 14 13 10 9 10 9 10 9 9 2
13 13 0 10 9 1 10 15 13 10 9 1 9 2
23 13 13 9 0 9 1 10 9 15 10 0 9 2 1 15 13 10 0 9 1 10 9 2
57 10 9 7 13 9 1 10 0 9 13 10 9 10 0 9 10 0 9 7 13 14 13 10 9 1 9 7 1 0 9 7 14 13 1 9 14 13 9 2 7 10 9 14 13 3 14 13 7 13 10 9 1 15 10 0 9 2
10 10 9 15 13 0 1 10 9 9 2
21 10 0 9 13 7 2 9 9 13 1 9 10 9 15 2 9 9 7 0 9 2
5 13 10 9 15 2
16 15 14 13 0 9 1 9 10 0 9 10 9 9 1 9 2
8 0 15 13 7 13 14 13 2
37 7 10 9 10 9 2 7 3 1 10 9 10 9 10 9 10 0 9 2 13 14 13 7 10 9 13 15 15 13 10 9 1 10 9 10 9 2
34 10 9 10 0 9 2 9 9 2 7 10 0 10 0 10 9 7 3 9 10 9 2 9 9 2 13 10 9 15 1 9 10 9 2
21 1 10 9 10 0 9 10 9 10 9 10 12 9 13 1 10 9 0 0 9 2
12 0 9 13 3 14 13 3 1 10 9 15 2
8 1 0 9 10 9 1 9 2
10 10 9 13 12 12 10 0 12 9 2
25 13 7 3 1 12 9 13 9 2 7 10 12 10 9 14 13 9 7 7 13 14 13 12 9 2
15 10 9 10 9 10 9 2 10 9 9 9 2 13 0 2
30 1 0 9 10 9 2 3 1 10 9 2 1 10 0 9 1 0 9 7 1 9 12 9 2 13 10 9 0 9 2
15 3 2 10 9 9 13 12 9 1 12 9 10 9 9 2
15 10 9 13 10 0 9 7 10 9 13 10 0 0 9 2
47 3 13 14 13 1 15 15 13 10 9 9 1 9 10 0 15 9 7 14 13 3 1 9 10 0 15 9 10 0 9 7 10 9 1 10 0 9 15 13 10 0 9 1 9 10 9 2
13 9 9 2 13 0 7 15 10 9 13 15 13 2
13 13 1 0 9 10 12 7 13 10 9 10 12 2
18 10 9 13 14 13 9 10 9 1 10 9 15 15 13 10 9 15 2
10 13 10 9 10 9 10 9 1 9 2
23 3 13 2 1 12 9 9 2 10 9 10 9 9 10 9 9 7 10 0 10 9 9 2
33 1 9 2 13 3 9 15 10 9 14 13 1 12 2 14 13 10 9 7 14 13 0 9 1 0 9 1 10 15 13 14 13 2
20 13 3 10 0 9 1 9 10 9 2 3 10 0 9 2 13 10 0 9 2
50 10 9 10 9 2 10 9 10 9 15 13 10 9 2 13 13 1 9 2 1 9 10 0 9 10 9 14 13 0 9 14 13 1 10 9 15 10 0 0 9 2 10 15 13 13 1 0 10 9 2
35 1 15 10 9 2 13 0 10 9 10 0 9 1 12 9 9 15 13 3 1 12 9 9 2 10 15 13 10 0 9 1 0 0 9 2
17 3 1 10 0 9 2 15 9 14 14 13 10 0 9 10 9 2
21 3 1 10 9 13 10 9 0 7 0 9 2 9 2 9 2 0 9 7 9 2
16 13 3 10 9 15 14 13 3 1 9 10 9 7 10 9 2
11 3 10 12 10 9 13 1 10 0 9 2
36 1 9 2 0 9 15 13 1 10 9 9 2 13 12 9 15 13 1 0 9 0 0 1 9 3 9 1 0 9 15 13 10 9 1 9 2
55 3 13 10 0 9 10 9 2 9 9 2 2 10 9 9 9 1 9 13 10 9 9 0 9 2 7 7 2 13 1 9 10 0 9 10 0 9 2 10 2 7 10 9 7 7 3 13 9 1 10 9 10 9 2 2
33 3 1 9 10 9 9 13 3 9 2 9 15 13 9 2 3 9 2 7 3 3 1 9 10 9 10 9 9 13 3 3 0 2
45 3 3 14 13 0 10 9 10 0 9 2 13 0 14 13 3 10 14 9 15 2 3 7 0 9 10 9 10 0 9 7 9 10 9 10 9 10 0 9 3 1 10 0 9 2
8 10 9 13 10 9 10 9 2
15 7 13 14 13 10 9 2 13 14 13 14 13 3 0 2
33 10 0 9 2 14 13 14 13 10 9 14 13 10 0 9 7 14 13 15 0 2 1 14 13 10 0 1 10 0 7 0 9 2
19 10 15 9 10 9 15 13 1 9 10 9 7 10 9 1 9 10 9 2
34 1 10 9 10 9 0 13 2 13 7 14 13 14 13 1 9 15 1 2 10 9 9 7 10 0 9 2 2 3 13 13 10 9 2
55 10 3 9 10 0 9 0 9 2 9 9 2 13 0 9 1 9 2 1 3 13 14 13 1 0 9 7 10 9 13 13 14 13 7 3 14 15 13 14 13 1 9 2 7 13 14 13 9 1 10 0 9 10 2 2
21 1 15 10 9 1 10 9 10 0 13 12 0 2 7 12 13 0 1 0 9 2
66 10 12 9 13 10 9 15 13 1 10 9 10 0 9 7 10 0 9 10 9 2 10 9 15 13 1 10 9 10 9 10 9 14 13 10 9 15 13 10 9 7 1 10 0 9 15 10 9 1 9 15 2 15 13 3 13 1 10 9 2 1 10 9 0 9 2
1 9
27 13 3 7 3 9 0 1 9 10 0 7 10 0 0 0 9 14 13 14 13 10 0 9 1 9 9 2
65 3 1 15 2 1 10 9 10 9 15 3 1 9 13 7 13 10 9 0 9 3 13 10 9 10 13 2 10 9 9 1 9 2 10 9 7 10 9 2 10 9 10 0 9 3 7 10 9 10 9 10 0 9 3 1 10 9 10 0 9 1 10 0 9 2
20 10 9 13 7 10 0 0 9 13 1 9 2 13 0 9 3 7 15 9 2
39 1 15 10 9 2 3 13 2 15 13 0 14 13 10 9 1 10 15 13 1 9 10 9 3 1 10 12 3 3 1 10 9 10 9 9 1 0 9 2
51 3 7 10 9 2 10 9 9 9 1 9 15 2 13 7 10 2 0 9 2 14 13 12 1 10 12 0 9 15 14 13 10 0 9 2 7 10 9 10 9 14 13 3 10 0 0 9 2 10 0 2
9 3 3 10 9 10 9 3 13 2
34 3 1 15 10 9 2 10 0 9 2 9 9 2 7 2 9 9 2 13 0 1 9 10 9 12 15 13 2 7 14 13 9 9 2
22 10 9 2 9 10 9 1 0 15 9 10 0 9 7 10 0 9 13 0 0 9 2
26 10 0 9 13 13 3 1 12 9 9 1 10 12 2 9 1 10 15 10 9 15 13 10 9 15 2
20 10 9 9 2 3 7 10 9 2 13 1 9 7 10 9 15 13 3 9 2
31 10 3 13 1 10 9 10 9 2 10 9 2 7 13 10 9 9 14 13 1 10 9 7 1 9 7 1 10 0 9 2
14 10 14 0 9 15 13 1 9 15 13 9 0 9 2
38 3 1 10 9 10 0 13 10 9 10 2 2 2 10 9 10 15 13 0 9 0 1 10 15 7 0 9 2 3 13 10 9 9 1 9 15 2 2
14 10 9 14 13 14 13 2 7 7 10 0 15 9 2
33 10 0 9 3 1 10 0 9 13 13 9 0 1 10 9 1 14 13 1 0 9 15 7 7 14 13 10 9 15 15 15 13 2
4 9 9 1 9
25 3 1 10 0 9 9 2 13 0 14 13 3 2 1 10 9 10 9 2 7 0 9 1 9 2
29 13 2 3 2 1 9 2 10 9 1 10 9 2 1 9 10 0 9 10 9 7 1 0 9 9 10 0 9 2
17 13 3 10 0 9 1 9 1 0 9 1 10 0 9 10 9 2
7 1 0 9 10 0 9 2
29 3 1 10 0 9 9 13 10 9 15 7 13 10 9 7 14 13 15 10 9 10 9 15 1 9 10 0 9 2
33 1 9 13 3 10 9 10 9 10 0 9 2 13 1 9 10 12 9 1 9 1 10 9 9 3 2 1 10 0 9 7 9 2
34 13 3 3 3 1 9 10 9 7 3 14 13 3 15 10 9 2 7 14 13 10 9 10 9 2 15 13 10 9 15 1 10 9 2
37 10 9 10 9 13 3 1 9 2 1 10 15 10 9 13 10 9 0 9 12 9 7 10 9 15 1 9 2 9 2 2 1 10 15 13 3 2
16 10 9 15 13 1 9 7 3 1 9 7 10 9 13 0 2
11 9 1 9 13 10 0 9 1 0 9 2
14 10 0 9 10 9 13 1 0 9 10 9 10 9 2
12 14 15 13 3 7 15 13 15 3 1 9 2
17 10 9 7 10 9 13 10 9 15 13 3 1 10 0 0 9 2
43 1 9 10 9 10 9 10 9 10 9 10 0 9 13 1 0 9 2 1 2 0 2 9 7 3 1 9 10 0 9 10 0 9 7 10 15 9 9 10 9 10 9 2
8 10 9 13 1 10 0 9 2
24 12 12 9 13 1 0 9 10 9 2 7 10 0 9 13 9 1 10 9 1 10 9 9 2
14 10 0 9 9 13 1 9 7 13 9 1 10 9 2
11 14 13 7 10 9 9 7 9 13 13 2
46 10 0 9 2 7 7 10 0 9 3 1 10 9 7 10 9 2 13 1 10 9 15 0 9 1 14 13 10 9 14 3 14 13 10 9 10 9 7 7 14 13 1 0 0 9 2
63 1 0 15 2 13 10 9 10 9 9 7 10 9 15 1 10 0 9 1 9 15 13 13 1 10 9 2 10 15 13 1 9 10 9 10 9 7 1 9 10 9 10 2 9 1 9 2 7 7 10 0 9 13 1 0 9 9 10 0 9 10 9 2
24 13 1 10 9 15 7 13 7 14 13 14 13 10 0 9 7 14 13 10 9 9 1 15 2
11 10 12 9 13 1 9 12 1 10 9 2
14 3 2 10 0 9 15 14 14 13 3 9 1 9 2
42 3 13 0 2 1 9 10 9 2 0 9 2 3 9 2 9 2 9 2 7 1 0 9 9 2 9 7 9 14 13 14 13 10 9 2 1 9 3 10 0 9 2
7 1 0 9 15 13 15 2
38 1 15 13 1 9 2 7 13 14 13 0 10 9 15 13 3 1 0 9 2 14 13 9 15 14 13 10 9 10 9 2 7 15 13 3 0 9 2
9 14 13 3 1 9 10 0 9 2
24 14 13 14 13 10 9 3 1 15 13 1 9 3 7 3 7 13 7 13 14 13 10 9 2
21 1 9 3 13 10 9 7 10 0 1 10 9 10 9 9 13 1 10 0 9 2
21 10 9 15 13 3 1 9 1 12 9 12 2 7 14 13 7 1 9 10 12 2
4 14 13 3 2
43 1 0 9 3 10 9 14 13 14 13 2 3 2 1 15 15 13 10 9 2 3 2 15 13 15 13 10 9 7 3 1 15 13 14 13 1 15 1 9 1 10 9 2
27 13 3 9 14 13 10 9 10 15 13 7 10 15 13 7 1 9 10 9 14 13 14 13 1 0 9 2
19 1 0 9 15 2 10 9 13 7 13 1 0 9 1 10 9 10 9 2
27 3 13 10 9 10 2 9 2 13 0 10 9 2 7 13 7 15 13 3 10 9 14 13 10 0 9 2
35 3 9 10 9 2 10 9 7 10 9 15 2 13 3 0 10 9 10 9 15 13 13 10 9 0 1 12 9 3 2 10 3 0 9 2
24 3 9 10 9 10 9 9 9 2 1 9 2 13 1 12 9 9 1 10 3 0 9 9 2
39 13 10 9 2 10 15 13 10 9 9 1 0 9 2 10 9 1 10 9 7 10 9 10 9 2 10 9 13 14 13 1 15 10 9 0 9 7 9 2
16 9 13 7 2 0 10 9 10 9 13 0 1 10 0 9 2
26 13 1 9 9 7 14 13 7 10 9 15 13 3 10 0 9 2 2 13 10 9 9 10 0 9 2
20 10 0 9 13 15 9 14 13 1 9 10 0 2 1 9 14 13 12 9 2
20 10 9 2 3 1 10 9 2 13 13 1 9 12 9 10 9 1 10 9 2
19 10 9 10 0 9 14 13 0 2 3 7 13 10 0 9 10 0 9 2
39 13 7 0 9 9 13 13 10 9 10 9 1 9 0 9 2 7 1 10 9 15 1 15 14 13 15 2 10 9 14 13 10 9 0 9 0 10 9 2
35 10 9 10 2 2 9 9 2 13 10 9 15 7 14 13 0 10 0 9 2 13 7 10 0 9 2 1 14 14 13 10 9 0 9 2
33 3 14 13 7 14 13 10 3 2 10 9 14 13 3 10 0 9 2 7 13 3 7 0 9 2 13 9 10 0 9 10 9 2
30 1 9 15 2 10 9 13 1 10 0 9 10 9 1 9 1 10 1 3 0 9 7 14 13 1 9 10 0 9 2
15 3 13 0 2 3 10 9 14 13 0 9 1 10 9 2
44 15 13 10 9 15 1 9 14 13 14 15 13 1 0 9 2 13 1 9 15 1 0 9 10 9 9 10 9 2 9 9 2 13 3 7 14 13 14 13 9 10 9 15 2
13 9 2 13 9 3 1 9 1 14 13 10 9 2
27 10 9 1 0 10 9 9 9 13 10 9 10 9 1 9 3 12 10 9 12 2 12 1 12 0 9 2
19 3 13 14 13 7 10 13 1 9 9 14 13 1 10 9 10 0 9 2
24 10 9 15 13 1 9 15 1 10 0 9 2 9 15 13 10 0 7 0 9 10 9 9 2
7 3 13 14 13 0 9 2
25 3 1 10 9 10 0 9 2 2 10 9 13 7 15 9 13 14 13 9 1 10 9 9 9 2
33 10 9 1 10 9 10 9 3 7 1 10 9 10 9 13 1 0 9 15 13 1 9 1 10 9 9 9 2 2 13 1 9 2
32 10 9 13 1 15 9 10 12 9 10 0 9 3 1 10 0 15 0 9 2 7 3 10 12 9 10 9 0 7 0 9 2
3 3 3 2
17 3 2 10 9 13 10 9 10 9 9 2 12 2 10 0 9 2
19 13 2 3 2 14 13 7 10 9 10 15 13 10 1 9 9 13 0 2
17 1 9 9 13 1 10 9 10 9 2 13 3 10 9 10 9 2
7 1 0 9 13 10 0 9
20 1 2 0 9 0 9 2 1 9 13 9 10 0 9 9 1 9 15 13 2
43 13 14 13 10 0 9 10 9 10 0 9 10 9 1 10 0 9 0 7 0 9 7 13 10 9 15 1 10 0 9 3 1 10 9 10 9 15 13 1 10 9 9 2
16 3 2 10 12 0 10 9 13 1 0 0 9 1 9 9 2
20 10 9 2 1 10 9 15 2 13 7 14 13 10 0 7 0 9 10 9 2
21 0 9 13 7 13 3 1 9 10 9 2 7 15 15 13 3 13 15 10 9 2
16 10 9 2 3 2 13 1 9 9 1 9 7 9 10 9 2
9 2 10 0 9 13 1 0 9 2
4 9 1 9 2
30 3 2 1 9 2 13 9 3 1 10 0 9 2 1 9 10 9 2 9 2 7 10 9 9 14 13 10 9 15 2
44 1 10 9 10 9 10 9 9 13 0 9 2 3 10 9 10 9 2 10 9 9 0 9 7 10 0 9 1 10 9 2 0 10 9 10 9 9 7 10 9 10 9 9 2
18 10 9 10 9 13 1 14 13 10 9 2 10 9 7 10 9 9 2
29 1 9 10 9 1 9 1 10 9 10 9 14 13 10 9 2 3 12 9 13 13 10 9 15 1 10 0 9 2
19 13 3 7 10 0 9 13 0 7 13 10 9 10 9 10 0 0 9 2
11 10 9 2 3 2 13 10 9 1 9 2
44 14 13 14 13 1 2 9 7 13 13 10 9 3 13 14 13 3 3 0 9 7 7 10 9 2 15 13 1 9 14 13 3 10 0 7 0 9 1 9 1 10 0 9 2
6 10 0 9 10 9 2
24 3 2 1 9 2 10 9 13 7 10 9 10 9 3 7 3 3 0 13 1 9 10 9 2
14 3 10 9 13 0 1 10 9 9 10 2 1 9 2
8 15 13 10 9 1 15 13 2
27 10 9 13 12 9 1 15 10 9 9 13 7 14 13 0 2 1 9 10 9 14 15 13 9 0 9 2
3 2 2 2
44 10 2 9 13 1 0 0 9 9 2 13 7 10 9 2 9 2 2 15 13 13 10 9 9 2 13 14 2 13 2 10 0 9 1 0 9 7 10 9 0 9 0 9 2
24 3 2 10 9 9 10 2 13 13 10 1 9 9 2 13 2 0 2 10 0 9 15 13 2
18 1 15 10 9 10 9 13 3 7 12 9 1 0 9 10 0 9 2
1 9
27 10 9 1 9 1 10 2 14 13 14 13 3 7 10 9 10 0 9 13 7 15 14 13 3 0 9 2
28 3 2 13 0 14 13 10 9 3 7 14 14 13 7 10 9 9 9 13 10 0 2 7 3 0 2 9 2
24 3 2 13 0 1 0 10 0 9 7 13 9 15 13 10 0 9 0 9 1 15 1 15 2
22 0 0 9 13 10 9 10 3 13 9 15 14 13 10 0 9 1 9 10 0 9 2
7 15 14 13 12 0 9 2
18 1 0 9 1 10 9 13 10 9 7 10 9 0 9 7 3 9 2
35 3 2 10 0 9 13 3 0 7 0 9 10 0 9 1 9 15 13 0 9 2 3 7 3 1 10 0 9 3 1 10 9 10 9 2
35 10 9 9 10 2 2 9 9 2 13 3 9 1 9 10 0 9 2 1 15 13 10 0 9 1 9 15 13 13 10 9 1 9 15 2
18 3 1 10 12 2 13 14 13 1 9 7 14 13 14 13 0 9 2
22 3 1 10 9 9 10 9 9 9 9 2 10 0 9 13 0 1 0 7 0 9 2
36 10 9 15 10 9 13 1 10 0 9 2 1 15 10 9 10 9 10 0 9 7 10 9 12 10 9 9 10 0 9 13 1 15 15 9 2
23 10 9 10 9 13 7 2 10 9 9 1 10 0 9 14 13 10 9 1 10 2 2 2
7 0 9 1 9 9 1 9
22 10 0 9 13 10 9 2 1 9 10 9 2 1 9 1 9 0 9 7 9 9 2
32 1 10 9 15 13 0 14 13 3 10 0 9 2 14 7 12 9 2 12 1 10 9 10 9 9 7 12 1 9 10 9 2
25 13 7 10 12 12 14 13 14 13 9 12 12 9 2 7 10 12 13 14 13 1 12 9 9 2
27 10 9 13 1 12 10 9 1 10 0 9 10 9 1 10 0 9 7 13 1 0 0 9 12 9 3 2
40 1 10 9 15 3 10 9 10 9 15 13 10 9 2 1 9 3 10 9 10 9 7 3 10 9 10 9 2 7 3 1 9 13 7 3 1 9 10 9 2
34 13 10 9 10 9 7 13 0 9 2 0 9 7 0 9 2 1 10 15 3 9 10 9 2 10 15 13 1 10 0 9 1 9 2
43 1 9 10 0 9 2 7 14 2 13 2 10 0 9 10 9 2 10 9 13 1 0 9 7 0 9 2 7 10 9 10 9 13 3 14 15 13 1 9 10 0 9 2
12 1 3 2 13 13 0 10 9 15 10 9 2
13 15 1 9 15 13 15 2 10 9 10 9 2 2
19 10 0 9 7 10 0 9 1 10 0 0 9 13 0 10 9 10 9 2
26 10 9 15 13 12 9 1 10 9 10 9 9 1 10 9 10 9 10 9 2 1 9 1 0 9 2
35 10 9 13 0 2 7 1 15 13 0 0 9 15 13 2 15 9 2 9 0 9 1 10 9 7 1 10 9 2 9 2 9 7 9 2
17 10 9 13 1 9 9 1 9 7 7 10 0 13 13 14 13 2
1 9
29 14 13 0 3 9 1 10 2 9 7 15 9 3 1 10 9 10 9 7 14 13 10 9 7 10 9 10 9 2
26 10 9 9 13 3 12 9 1 0 9 1 10 0 9 10 9 2 7 13 1 10 9 9 1 9 2
43 14 13 7 14 13 13 1 10 9 10 9 10 15 2 3 13 2 13 10 9 10 9 10 9 9 2 7 10 15 14 13 10 9 10 9 10 9 1 9 3 10 12 2
26 3 2 13 15 10 9 3 0 15 2 7 15 10 9 2 3 15 13 2 13 3 1 10 9 15 2
28 13 1 0 9 7 0 9 2 3 1 10 3 9 2 13 3 14 13 10 9 10 0 9 3 9 10 9 2
11 3 9 10 9 10 9 13 1 12 9 9
20 10 9 15 13 14 13 0 3 3 1 9 9 15 13 10 9 7 10 9 2
47 10 0 9 10 0 9 13 7 2 10 0 10 0 9 10 0 9 2 9 9 2 13 10 9 1 9 9 9 2 10 9 9 1 9 2 10 9 1 10 9 10 9 1 10 9 2 2
29 10 0 9 13 1 10 0 9 9 14 13 1 9 1 10 0 9 9 15 13 9 1 9 1 3 0 0 9 2
5 10 9 1 10 9
28 10 9 13 7 14 13 10 9 10 9 9 9 2 3 9 10 0 9 10 9 1 10 9 10 9 9 9 2
33 1 9 13 9 2 15 14 13 0 10 9 2 10 15 13 7 10 9 14 13 14 13 3 7 1 9 1 10 0 9 1 9 2
82 10 9 13 3 9 10 0 0 9 2 10 0 9 2 10 12 12 0 9 15 13 10 12 9 2 7 9 3 2 13 14 15 13 2 10 9 9 2 10 9 9 12 9 2 10 9 9 2 10 9 9 2 10 9 9 2 10 9 9 2 10 9 9 2 10 9 9 2 10 9 9 7 3 10 9 9 2 3 9 10 9 2
5 12 9 9 1 9
19 3 2 10 9 3 1 9 10 9 2 10 9 13 1 10 9 10 9 2
36 13 0 9 1 15 9 1 9 1 9 7 9 2 9 9 9 2 2 2 7 7 13 1 9 2 10 9 10 9 15 13 14 13 10 9 2
40 15 9 2 15 13 15 9 2 13 1 10 9 10 0 9 9 1 15 9 1 10 15 3 13 2 7 14 13 7 15 13 10 0 0 9 1 10 9 15 2
19 3 2 10 9 9 10 15 13 9 1 10 9 14 13 14 13 1 9 2
1 9
16 3 2 0 9 14 13 10 9 14 13 10 9 1 10 9 2
1 9
7 0 15 14 13 14 13 2
18 0 15 9 13 14 13 10 9 15 7 14 13 1 9 0 0 9 2
12 10 9 15 13 10 0 9 1 10 9 9 2
15 1 10 3 2 10 9 10 2 1 1 0 9 13 3 2
34 1 10 9 1 9 10 9 2 1 9 10 9 2 10 9 15 13 10 12 9 2 12 9 7 12 9 2 7 3 13 15 12 9 2
15 10 12 9 14 13 1 2 9 9 2 2 1 12 9 2
14 10 9 10 9 13 10 9 2 10 9 7 10 9 2
24 7 2 3 1 10 9 10 9 2 14 13 14 13 9 2 7 10 9 13 14 13 9 3 2
24 1 9 10 0 9 13 3 10 9 9 2 9 10 9 9 2 9 2 7 15 0 0 9 2
12 9 10 9 10 0 9 1 10 0 9 10 2
37 1 3 2 10 9 10 9 13 0 2 7 13 7 10 9 2 1 15 13 13 10 9 2 13 0 7 7 15 10 9 1 9 14 13 0 9 2
59 7 2 13 9 3 13 10 9 10 0 9 15 14 13 3 0 2 13 3 9 7 0 7 13 1 15 10 9 14 13 0 1 10 9 1 14 13 13 0 9 7 14 13 13 9 3 1 10 7 10 9 13 0 1 10 9 7 14 2
28 10 0 9 10 2 13 7 2 14 13 10 9 9 10 9 2 1 9 9 1 10 9 3 12 9 9 3 2
31 3 2 10 12 10 9 13 10 9 10 0 9 1 10 9 2 3 7 7 10 0 9 14 13 0 14 13 10 9 15 2
15 3 2 10 3 9 13 1 9 2 9 2 9 7 9 2
31 10 9 13 7 10 9 1 9 10 9 2 3 13 1 10 9 10 0 9 2 13 10 3 0 9 1 10 9 10 9 2
36 1 3 10 0 9 13 1 9 10 0 9 9 10 0 9 2 7 13 0 14 13 3 1 14 13 14 13 10 9 10 9 1 0 0 9 2
1 9
50 10 0 9 2 1 14 13 0 2 13 14 13 1 0 9 1 9 9 2 3 3 13 10 9 10 9 10 9 7 10 0 9 15 13 1 10 0 9 2 10 15 13 14 13 0 2 0 7 0 2
48 3 2 3 1 10 12 9 15 14 13 10 9 2 7 13 15 9 1 10 9 2 10 9 7 10 9 2 14 14 13 3 10 9 15 13 3 1 10 9 10 2 2 10 9 7 10 9 2
18 10 9 9 10 9 13 0 9 3 1 10 9 3 7 1 10 9 2
4 10 9 10 9
32 14 13 14 13 10 9 7 13 14 13 1 0 10 9 15 1 14 13 15 9 14 13 14 13 1 9 15 1 10 9 9 2
12 1 15 14 13 10 9 10 9 7 10 9 2
15 10 12 10 9 14 13 14 13 1 0 9 2 3 13 2
37 2 10 9 13 0 9 2 2 13 10 9 9 10 9 9 1 10 9 10 9 2 2 1 0 10 9 15 13 1 9 2 13 10 0 9 2 2
30 1 10 0 9 15 13 1 9 10 9 9 3 10 9 2 10 12 9 9 13 3 10 9 15 1 10 9 10 9 2
19 10 9 15 13 3 1 9 2 1 15 13 9 10 0 2 15 15 13 2
6 15 13 15 9 9 2
36 1 0 9 0 10 12 2 10 9 9 13 10 12 10 9 2 10 9 9 13 10 12 2 10 9 9 10 12 7 10 9 9 13 10 12 2
20 7 2 13 0 1 12 9 2 7 1 9 10 9 13 13 7 9 1 9 2
13 10 0 9 10 0 9 14 13 1 12 9 2 2
1 9
23 13 3 3 3 7 3 0 9 1 10 12 15 9 9 10 9 2 3 3 7 12 9 2
1 9
14 10 9 10 9 10 9 1 10 9 9 13 14 13 2
12 10 0 9 3 10 0 15 9 13 10 9 2
28 10 9 13 10 0 9 9 1 9 7 12 1 10 0 10 9 2 0 9 12 2 1 10 9 1 10 9 2
24 14 13 15 14 13 7 10 9 13 1 9 10 0 9 3 1 10 3 9 10 0 10 9 2
23 10 9 14 13 3 15 14 13 10 0 2 10 9 7 10 9 7 15 3 9 2 14 2
7 3 2 14 13 1 9 2
22 10 9 13 10 9 10 0 9 2 7 3 1 15 9 1 0 9 13 10 0 9 2
21 14 13 3 14 13 7 1 9 9 14 14 13 3 14 13 9 3 9 1 0 2
31 10 9 9 13 2 3 2 12 2 1 10 9 2 12 2 1 10 9 2 12 2 1 10 9 7 12 2 1 10 9 2
41 1 0 9 2 10 9 13 10 0 7 10 9 10 9 14 13 10 0 9 2 14 13 10 0 9 1 9 10 9 7 10 9 7 14 13 1 10 0 9 9 2
34 1 10 9 10 9 10 9 2 15 9 1 10 9 13 1 9 7 10 9 10 9 15 13 1 9 15 13 3 0 1 10 9 15 2
60 7 10 9 10 9 3 13 10 9 10 9 2 10 9 9 15 13 1 0 2 1 13 9 12 2 9 2 2 7 10 9 0 0 1 0 9 1 2 13 9 7 10 9 0 13 3 10 0 9 9 1 2 2 9 10 15 13 1 3 2
13 13 7 0 14 14 13 7 0 9 10 0 9 2
22 10 9 9 13 10 9 9 1 9 12 2 1 9 10 9 10 12 10 9 9 12 2
26 10 0 2 7 0 9 2 7 3 15 2 9 9 2 3 7 10 2 9 13 1 15 1 0 9 2
30 10 9 9 10 9 13 7 10 9 10 2 13 2 0 9 1 10 0 9 2 14 13 10 0 9 15 1 0 9 2
19 2 3 7 14 13 1 9 15 2 2 13 10 9 2 15 7 14 13 2
52 10 12 9 13 10 9 0 9 1 10 15 13 12 9 2 14 3 1 0 0 9 2 7 1 0 10 9 10 0 9 10 9 2 10 9 15 13 3 3 1 10 0 9 15 13 15 10 9 1 10 9 2
27 10 9 13 1 10 0 9 10 9 1 9 15 13 2 3 2 15 0 9 1 10 12 2 1 10 12 2
20 10 2 13 1 12 9 10 12 2 7 10 3 0 9 13 13 1 12 9 2
45 13 3 2 3 7 15 9 2 7 2 10 9 13 3 14 13 10 0 15 9 7 14 13 10 0 15 9 7 14 14 13 10 9 7 15 13 9 0 9 7 3 10 9 2 2
31 1 15 12 0 14 13 3 13 2 3 1 9 10 9 2 3 13 10 9 9 2 10 15 13 7 10 9 13 3 12 2
42 10 9 14 13 14 13 1 15 0 9 2 1 15 9 2 7 2 14 13 14 13 9 3 1 10 15 9 0 1 10 9 7 14 13 14 13 10 9 10 9 15 2
8 9 2 12 10 0 1 9 2
34 7 10 0 9 13 10 0 9 9 2 3 13 1 9 2 3 1 10 9 10 9 2 13 7 14 13 2 2 13 14 13 3 2 2
57 10 9 9 2 15 13 1 12 9 1 9 9 10 9 9 10 9 2 13 13 9 1 10 9 2 7 13 3 10 9 7 10 2 9 13 13 7 1 14 15 13 9 14 13 14 13 14 13 15 9 1 10 0 9 10 2 2
27 3 2 10 9 13 2 9 2 2 2 9 9 2 2 2 0 9 2 2 7 7 2 9 10 9 2 2
57 3 2 10 9 13 14 13 0 9 2 0 0 9 2 10 0 9 10 9 2 9 1 10 0 9 2 10 9 2 10 9 2 10 9 10 9 9 2 10 9 10 9 2 10 12 9 9 2 2 7 7 9 0 7 0 9 2
24 3 13 13 3 3 10 9 10 0 9 10 9 10 9 2 3 3 10 9 10 9 10 9 2
49 10 9 9 13 7 2 13 7 10 9 10 9 10 9 14 13 1 9 13 9 1 10 9 2 2 7 13 10 9 10 9 7 2 10 9 10 9 14 13 14 13 1 10 0 10 9 15 2 2
1 9
37 9 10 9 13 7 2 10 0 9 13 14 13 10 9 10 0 9 14 13 9 10 9 15 13 1 10 9 9 15 13 7 13 10 0 9 2 2
10 13 15 1 15 13 14 13 0 9 2
27 1 10 9 15 13 7 2 3 1 10 0 15 9 2 10 9 10 9 9 14 13 10 0 15 0 9 2
12 3 13 10 9 2 14 13 14 13 0 9 2
30 1 10 9 10 9 10 9 10 9 10 2 9 2 15 2 1 9 2 13 10 0 9 7 14 13 10 9 10 9 2
29 10 9 13 2 1 10 12 9 9 1 10 9 2 10 0 9 1 10 9 10 9 10 9 7 10 0 9 15 2
33 1 10 9 13 15 14 13 1 12 9 10 9 2 1 15 1 12 9 10 9 2 7 1 0 9 9 3 1 12 9 10 9 2
24 15 13 1 9 15 7 15 13 14 13 1 9 7 9 1 12 9 10 9 15 15 13 3 2
11 3 7 10 9 2 13 2 13 3 9 2
38 10 9 15 2 13 1 0 10 9 10 0 0 9 2 13 10 9 15 14 13 1 3 9 2 3 7 10 9 15 14 13 10 9 3 10 0 9 2
34 13 2 3 2 7 10 9 10 3 0 9 3 10 0 9 9 13 14 13 10 9 10 0 9 14 13 15 10 9 10 0 15 9 2
18 10 9 1 0 9 14 13 3 1 9 0 9 7 1 9 0 9 2
8 2 10 9 15 13 9 9 2
41 10 0 10 9 9 10 9 2 9 9 2 13 7 2 7 15 1 10 0 14 13 14 13 10 12 10 9 2 12 9 10 0 9 14 13 1 12 7 12 9 2
49 10 9 10 9 10 9 10 9 1 10 9 0 9 13 13 10 0 7 13 13 10 9 9 2 10 15 13 3 1 9 7 14 13 10 9 2 14 13 10 9 1 0 9 7 14 13 10 9 2
54 15 10 9 15 13 7 10 0 2 0 9 2 2 10 9 2 10 9 2 10 9 7 10 3 9 2 15 13 7 14 13 10 9 10 9 1 0 9 7 10 9 15 1 10 9 2 15 13 3 10 0 15 9 2
32 10 9 10 0 9 9 9 7 9 9 13 10 0 9 10 9 2 10 15 3 13 2 0 9 2 1 14 13 1 10 3 2
35 3 13 10 0 9 2 0 1 0 9 2 1 9 10 15 13 9 2 9 2 9 2 3 7 9 10 15 13 13 10 0 9 1 9 2
14 10 0 9 13 14 13 10 0 7 10 0 0 9 2
21 13 10 13 9 15 10 0 9 7 14 13 14 15 13 7 15 7 10 2 9 2
26 10 9 10 9 9 7 3 10 0 9 9 10 9 1 10 0 9 2 13 10 9 1 12 3 9 2
47 1 10 9 1 10 0 0 9 9 2 10 15 9 13 10 2 9 9 15 13 3 15 2 10 0 9 13 1 0 9 1 9 0 9 9 1 9 2 3 3 1 0 9 10 9 15 2
26 7 2 13 3 9 10 9 7 10 0 9 13 3 0 7 0 2 7 14 13 3 3 0 10 9 2
20 10 9 1 10 9 7 10 9 2 9 9 2 13 3 0 9 1 10 9 2
31 3 13 14 13 15 10 9 3 13 10 9 10 0 9 2 15 13 10 9 10 9 9 1 14 13 9 1 9 10 9 2
19 7 2 15 15 13 0 9 1 9 0 9 2 15 1 3 14 13 13 2
34 7 13 14 13 0 7 1 0 9 14 13 14 13 9 3 3 14 13 3 10 0 9 1 0 9 7 3 14 13 13 0 15 9 2
20 15 13 7 13 3 13 1 0 9 9 2 10 9 3 13 3 10 3 9 2
3 3 15 2
17 1 10 0 12 9 2 15 10 9 10 9 14 13 0 1 12 2
23 10 9 15 13 3 7 1 12 9 9 1 10 9 2 3 3 7 1 13 9 1 9 2
16 10 9 13 3 10 12 9 7 13 1 0 9 7 0 9 2
25 10 9 13 10 9 10 0 0 7 9 1 10 12 9 13 3 0 9 1 10 15 13 14 13 2
9 13 10 0 9 10 9 10 9 2
7 7 3 13 9 1 15 2
27 10 9 13 1 10 9 10 9 9 9 2 10 15 13 1 9 10 9 2 7 13 10 9 10 0 9 2
44 7 13 1 10 9 15 13 14 13 1 9 10 0 9 2 7 14 13 1 9 1 10 9 15 14 13 3 2 13 3 15 2 7 10 0 9 15 13 14 13 3 14 13 2
21 3 13 10 9 1 9 7 13 7 14 14 13 9 14 13 9 1 15 1 9 2
42 0 10 9 14 13 1 9 10 9 7 1 9 0 9 2 14 13 0 9 1 10 0 0 9 1 10 9 2 1 10 9 7 10 9 10 9 9 10 9 1 9 2
28 1 9 15 13 1 9 10 0 9 13 1 9 10 0 9 14 13 1 9 10 9 10 0 7 0 9 15 2
10 10 9 13 1 0 9 1 9 15 2
26 3 1 0 9 2 3 7 1 9 10 0 9 2 14 13 0 10 9 15 1 0 9 9 1 9 2
30 1 9 15 1 0 9 10 9 2 10 2 9 13 7 10 9 13 0 14 13 3 9 7 14 13 10 9 10 9 2
67 10 0 13 7 10 12 0 2 10 15 13 10 9 10 0 0 9 2 15 10 15 14 13 7 1 10 9 7 10 9 9 10 9 2 10 0 9 13 3 10 0 9 10 0 9 7 3 10 0 9 10 9 13 1 9 2 10 0 9 1 9 7 10 0 1 9 2
25 10 9 14 13 3 3 10 9 9 2 7 3 7 10 0 9 2 1 10 15 13 1 0 9 2
11 15 13 3 14 13 1 0 9 10 9 2
72 10 0 9 7 0 9 10 0 1 9 13 7 2 13 1 9 1 10 9 10 9 2 3 1 12 9 0 9 1 9 14 13 10 0 2 0 9 2 2 3 10 0 9 9 7 10 9 9 15 14 13 1 12 9 7 15 3 1 9 14 13 14 13 10 0 9 7 3 1 9 2 2
32 13 15 10 9 2 13 0 9 1 10 9 10 9 10 9 10 9 1 0 9 2 3 7 1 10 9 10 9 10 0 9 2
40 1 10 12 0 1 9 2 10 12 13 7 2 14 13 10 0 0 9 2 2 7 10 0 9 2 12 2 13 7 2 13 0 3 7 3 1 12 9 2 2
27 10 3 0 2 9 10 9 2 13 0 7 1 9 13 1 0 0 9 2 3 1 0 10 9 10 9 2
28 3 1 15 13 0 10 7 13 7 13 14 13 3 0 9 2 1 10 15 14 13 0 10 9 9 10 2 2
38 13 3 9 0 7 15 9 3 10 2 2 10 0 9 2 10 2 2 10 0 2 2 10 0 9 2 10 2 9 2 10 0 9 7 15 0 9 2
20 3 1 9 2 12 9 13 7 12 9 13 1 10 9 9 0 9 1 9 2
27 3 2 13 1 0 1 10 9 15 2 0 9 2 9 9 9 2 0 9 9 7 0 9 10 0 9 2
24 3 7 10 0 7 0 9 13 1 10 9 7 13 1 9 2 13 3 10 9 1 15 9 2
23 12 9 3 2 1 9 2 13 9 1 9 2 3 1 9 10 2 1 10 0 9 9 2
16 10 9 10 0 9 7 10 9 10 9 1 0 9 13 9 2
13 10 9 13 2 3 2 1 10 9 1 0 9 2
33 15 13 7 10 9 14 13 10 9 15 1 14 13 7 10 0 1 10 9 10 0 9 7 14 14 13 10 9 14 13 10 9 2
23 1 9 10 9 10 9 13 0 9 1 9 2 15 15 13 3 3 10 9 1 0 9 2
48 1 0 9 7 9 9 2 10 9 13 3 0 9 1 9 7 10 9 10 0 7 0 9 2 3 7 10 9 10 0 9 14 13 10 9 9 9 1 9 10 0 9 0 1 1 9 9 2
32 10 0 9 13 9 15 13 10 9 2 1 10 15 10 9 14 13 14 13 1 0 9 12 9 2 7 14 13 10 9 15 2
33 3 13 3 12 9 2 10 9 10 9 2 1 10 0 9 10 9 7 10 0 9 10 0 9 2 10 0 9 7 10 0 9 2
48 14 13 3 0 7 13 15 15 2 7 10 9 14 13 3 0 9 7 14 13 10 9 1 10 9 9 1 10 9 10 9 7 13 3 7 10 0 7 0 9 1 10 9 1 9 10 9 2
25 15 1 10 3 0 9 10 9 13 10 0 9 2 10 0 2 10 9 2 10 9 7 10 9 2
12 3 1 9 2 1 9 2 13 2 3 2 2
16 9 1 2 1 9 13 1 12 12 7 1 9 1 12 12 2
27 10 0 9 10 2 13 7 2 14 13 14 13 10 9 9 10 9 9 9 7 10 9 15 2 9 2 2
23 1 9 10 9 13 14 13 9 1 0 9 10 9 7 14 13 0 9 7 0 9 9 2
39 10 12 15 9 13 10 0 9 2 7 3 13 3 1 10 9 15 13 7 13 14 13 15 0 9 1 10 0 9 7 10 9 15 1 10 9 10 9 2
10 10 9 15 15 13 1 9 10 9 2
22 13 3 3 3 14 13 15 14 13 7 10 9 9 15 13 1 10 9 1 10 9 2
37 7 10 9 13 9 1 9 7 1 9 2 10 9 15 13 1 9 2 13 1 9 2 3 1 9 3 13 13 0 1 12 9 7 13 9 15 2
71 7 2 10 9 15 13 7 2 3 3 10 9 10 9 13 1 15 9 1 15 10 9 2 15 1 15 14 13 1 9 7 13 1 10 0 9 2 14 13 3 14 13 1 15 10 9 2 7 1 9 14 13 14 13 9 1 9 7 1 9 7 14 13 10 9 15 10 9 10 9 2
10 3 10 9 13 14 13 1 0 9 2
29 1 9 10 9 13 7 0 9 3 10 9 13 9 2 13 3 10 9 2 10 15 13 13 1 10 9 10 9 2
32 0 9 13 10 9 10 0 9 1 9 1 0 9 10 9 1 10 9 7 7 1 0 9 14 13 10 0 0 9 1 9 2
19 3 13 10 9 10 9 10 9 2 14 15 13 1 10 9 10 9 9 2
25 7 14 15 13 2 10 9 15 13 1 9 2 0 1 9 7 9 2 10 15 13 0 7 0 2
12 7 15 14 13 15 9 1 10 2 9 9 2
17 15 1 9 14 13 0 7 14 14 13 3 14 13 14 13 9 2
24 10 9 1 10 9 9 7 9 9 2 10 12 13 0 9 7 10 12 9 10 9 10 9 2
13 14 13 14 13 10 0 9 1 9 3 10 9 2
29 15 13 3 0 9 2 7 3 1 9 10 9 10 9 15 13 1 0 1 10 9 10 9 13 10 9 0 9 2
19 1 9 15 9 10 0 9 13 10 0 9 15 10 9 15 13 1 0 9
33 2 3 2 13 2 7 14 13 9 10 13 9 7 10 9 14 13 3 10 9 15 7 3 14 13 1 9 2 13 10 2 9 2
6 13 0 15 10 9 2
30 1 9 15 2 13 15 0 9 14 13 2 1 9 1 15 2 7 10 9 14 13 0 9 9 1 9 9 7 9 2
26 10 9 10 9 1 10 9 13 1 10 0 0 9 2 10 15 13 10 9 10 9 1 10 3 9 2
51 10 9 10 9 2 9 9 2 13 1 1 9 9 1 9 15 1 10 0 0 9 2 2 13 7 2 10 9 9 9 14 13 14 13 13 3 3 7 14 13 13 10 9 15 1 15 0 9 15 2 2
24 3 1 10 9 2 10 9 13 13 0 9 3 10 12 9 7 13 10 9 9 10 9 9 2
22 1 9 13 10 9 10 0 9 10 9 2 10 15 13 1 12 9 9 10 0 9 2
9 13 7 10 9 9 13 10 9 2
14 1 10 9 10 9 14 13 3 10 0 9 10 9 2
24 15 13 0 9 10 9 12 10 9 9 2 10 15 13 1 9 14 13 10 9 1 15 9 2
16 0 13 10 9 7 0 10 9 9 13 1 0 9 12 9 2
36 1 10 9 15 13 3 10 9 9 1 9 10 2 14 13 7 10 0 9 13 13 3 2 3 3 1 10 0 0 9 15 13 10 0 9 2
17 10 9 7 13 10 9 10 9 7 10 9 13 1 0 9 3 2
1 9
10 14 13 3 1 9 14 13 10 9 2
25 3 2 10 1 9 9 13 10 9 2 3 1 9 10 9 7 7 1 9 10 9 7 10 9 2
39 3 1 10 9 2 13 3 7 3 1 10 0 9 10 9 1 10 9 2 10 9 15 13 1 9 14 13 10 0 9 2 13 2 2 13 10 9 2 2
67 1 10 0 10 9 2 10 9 13 1 10 9 3 1 10 9 2 1 2 2 12 2 7 10 9 1 0 9 2 3 10 9 13 10 0 9 1 10 9 15 2 3 1 10 9 12 10 9 2 15 13 1 10 9 10 0 9 2 14 15 13 14 13 1 10 9 2
21 13 7 13 1 10 0 9 2 10 15 3 13 3 7 0 9 3 9 10 2 2
35 3 2 10 9 9 10 9 13 10 9 1 9 9 1 0 9 2 10 15 2 1 12 9 2 13 13 1 9 10 9 15 0 0 9 2
18 10 9 9 13 1 9 9 10 9 7 2 10 9 14 13 0 2 2
2 12 2
20 3 2 13 3 7 10 9 13 10 9 7 10 9 14 13 10 0 15 9 2
15 0 10 9 13 14 13 9 14 13 3 12 9 10 9 2
6 13 7 10 0 9 2
29 3 3 1 10 9 13 10 9 9 2 10 0 9 2 10 15 13 10 0 9 1 10 9 9 1 9 0 9 2
8 12 2 9 1 2 13 9 2
29 10 12 15 9 14 13 14 15 13 1 10 9 7 10 9 10 0 9 15 14 15 13 14 13 1 15 10 9 2
47 7 13 3 13 0 9 1 15 2 13 7 10 0 9 2 10 15 13 10 0 9 2 13 0 3 7 15 9 2 7 10 2 2 10 15 13 10 9 2 14 13 0 3 1 10 9 2
27 14 13 10 9 10 9 3 2 13 10 9 9 2 7 1 12 1 12 9 10 9 10 9 14 13 2 2
4 2 2 9 2
29 13 7 10 0 9 14 13 10 9 14 13 10 15 0 9 14 13 13 10 9 3 10 0 9 13 1 9 15 2
47 10 9 0 9 7 9 15 13 13 1 15 1 10 12 9 13 10 0 9 1 10 9 1 10 0 9 9 2 1 10 0 9 2 10 9 7 10 9 1 10 9 1 10 9 10 9 2
11 10 2 14 13 10 9 9 10 9 9 9
60 13 1 10 9 9 2 1 15 13 12 9 9 2 1 10 9 15 10 0 9 1 9 10 9 10 9 10 9 1 10 0 9 10 0 9 2 1 14 14 13 1 0 9 15 13 1 9 10 9 10 9 7 3 7 10 9 1 10 9 2
32 13 15 14 15 13 7 3 1 10 9 15 13 10 9 10 9 15 1 10 9 9 2 10 15 15 13 14 13 15 10 9 2
5 13 14 15 13 2
39 12 1 10 0 9 10 9 2 15 3 13 3 10 15 10 15 2 13 3 1 10 0 9 1 10 0 0 9 1 10 9 9 1 0 1 10 0 9 2
48 10 9 9 13 2 0 1 9 15 13 1 9 2 7 2 10 0 13 10 9 1 10 9 10 0 9 10 9 9 2 7 7 2 7 10 9 9 13 9 2 13 14 13 10 0 9 2 2
30 10 0 13 9 10 9 9 2 13 10 9 7 13 9 10 9 9 1 14 13 9 2 10 15 14 13 10 0 9 2
19 3 2 10 9 13 14 13 10 9 10 9 15 13 1 10 9 10 9 2
46 7 7 10 0 9 7 10 0 9 13 7 10 9 10 9 13 0 2 10 9 10 9 10 9 9 9 13 1 10 0 9 2 0 9 2 2 13 3 15 15 13 9 9 0 9 2
32 13 0 9 7 1 9 10 9 10 9 10 9 9 9 2 9 9 2 13 14 13 3 9 10 0 9 9 2 9 10 9 2
23 13 7 10 9 1 10 15 13 13 14 13 2 3 2 0 7 14 15 13 1 0 9 2
31 10 9 13 14 13 0 9 7 10 0 9 13 1 9 9 2 1 9 14 13 10 9 10 9 9 2 15 13 1 9 2
7 10 0 9 9 1 9 2
71 10 12 2 0 9 1 10 9 15 2 13 10 9 2 1 10 12 2 10 12 10 0 9 1 0 3 9 2 7 0 9 7 3 7 9 2 13 3 0 9 3 13 10 9 10 0 9 10 12 2 1 10 0 9 14 13 3 10 0 9 10 12 10 9 10 9 15 13 1 9 2
38 7 14 13 10 9 10 0 9 1 10 9 13 9 1 9 7 9 1 7 1 10 9 2 7 3 1 9 2 15 13 13 14 13 10 9 10 9 2
47 10 9 14 13 14 13 10 9 10 9 7 10 9 10 0 1 10 0 9 2 3 10 0 9 15 13 0 1 10 9 10 9 7 10 9 10 0 9 13 14 13 1 9 1 10 9 2
38 10 0 10 9 9 13 10 9 10 9 10 0 9 2 7 10 0 9 13 13 1 10 9 10 9 15 13 1 10 0 9 10 3 9 9 9 9 2
13 9 9 2 10 9 13 0 9 15 10 9 1 9
11 3 2 13 14 13 3 9 1 10 9 2
21 2 10 9 15 1 10 9 13 7 10 0 9 10 9 14 13 1 9 10 9 2
9 1 10 0 9 13 0 0 9 2
9 10 9 1 10 9 13 3 0 2
28 7 2 14 13 14 15 13 10 9 1 0 9 15 14 13 3 3 0 7 0 0 9 1 10 12 9 9 2
18 10 9 13 7 2 10 9 9 13 13 3 1 9 9 7 9 9 2
22 1 15 13 9 1 10 0 9 1 9 9 2 10 0 2 0 7 0 9 10 9 2
18 3 2 13 0 9 9 1 0 9 2 1 10 9 10 9 10 9 2
41 10 0 9 10 0 9 2 9 9 9 2 13 10 9 7 2 13 13 0 9 2 3 1 10 15 10 9 9 13 7 13 9 1 9 1 10 9 10 9 2 2
28 1 9 2 10 0 9 13 15 15 13 13 1 0 9 10 9 10 9 2 7 3 14 13 1 9 10 9 2
16 10 9 9 13 3 1 9 9 2 7 13 9 15 1 9 2
36 1 12 9 1 9 10 2 2 14 13 10 9 9 15 14 13 10 9 10 9 7 10 9 3 1 12 9 2 7 15 14 13 3 7 3 2
8 10 0 15 9 13 14 13 2
41 1 3 2 10 9 10 9 9 10 9 13 1 9 9 0 9 9 10 9 12 9 7 13 1 9 14 13 0 9 10 9 2 9 2 1 9 9 1 10 9 2
26 10 9 13 7 2 10 12 0 9 1 9 1 10 9 10 9 9 14 13 1 12 7 12 9 2 2
36 7 2 0 15 10 9 14 14 13 0 9 2 7 14 13 1 9 10 9 10 0 9 1 0 0 9 2 15 14 13 10 9 7 10 9 2
48 9 1 10 9 2 10 9 9 9 0 9 2 9 2 2 13 7 2 10 12 10 0 13 7 10 0 0 9 13 9 1 9 2 1 10 12 14 13 7 15 13 3 13 9 1 15 9 2
27 13 9 7 13 9 1 15 15 13 14 13 2 14 13 1 3 13 14 13 7 15 13 10 0 9 9 2
28 10 12 9 14 13 1 10 9 12 9 1 10 9 3 13 10 9 2 10 12 1 9 7 10 12 1 9 2
26 1 0 9 13 7 3 10 9 9 10 2 7 13 10 9 10 9 1 10 12 10 9 10 12 9 2
24 3 2 10 9 15 13 3 10 9 10 15 13 1 9 10 2 7 13 0 9 15 10 9 2
7 13 0 12 9 10 0 9
27 10 9 9 13 1 10 9 2 9 2 10 9 10 9 3 1 10 9 15 9 7 10 9 15 2 9 2
30 1 10 9 15 13 3 1 10 0 9 10 9 9 9 1 10 9 9 7 14 13 10 9 15 10 9 3 12 9 2
36 1 0 9 13 12 1 10 3 0 7 0 9 10 9 2 10 15 13 9 7 1 0 9 2 7 3 1 9 13 7 10 0 9 10 9 2
42 1 9 10 9 13 9 7 9 15 13 10 9 15 2 3 10 9 10 0 9 2 10 9 2 10 0 9 2 10 9 2 10 0 10 9 7 10 9 10 0 9 2
11 15 13 10 9 1 10 15 13 14 13 2
5 1 9 10 9 2
12 10 9 2 3 3 2 14 13 10 0 9 2
30 10 9 10 2 2 9 9 2 13 1 9 1 10 0 10 9 3 10 9 10 9 7 13 14 13 9 1 0 9 2
13 13 1 9 10 9 14 13 1 10 0 0 9 2
44 1 3 10 9 10 9 13 10 0 9 2 13 10 9 10 12 9 2 3 10 15 13 15 14 13 10 9 10 0 9 2 0 3 0 9 0 9 2 7 10 0 0 9 2
34 12 1 10 9 15 14 13 3 14 13 10 9 13 7 10 0 9 13 3 1 15 10 0 2 3 15 13 10 0 9 1 10 9 2
31 2 0 13 3 0 0 1 0 9 7 9 15 0 9 10 9 2 15 14 2 13 2 14 13 1 10 0 0 9 2 2
10 9 12 9 0 9 1 0 9 12 2
22 9 9 2 0 9 2 13 3 10 9 1 9 14 15 13 1 10 9 10 9 15 2
32 3 2 1 10 12 2 9 9 2 2 13 10 9 2 9 12 9 2 15 13 1 0 9 9 10 9 9 9 9 1 9 2
36 1 9 12 9 1 10 9 13 10 9 10 0 9 10 9 10 0 13 10 12 9 3 2 3 13 3 9 10 0 0 0 9 2 9 9 2
27 1 9 1 10 12 2 10 9 13 1 12 9 2 3 13 13 1 12 9 1 9 1 10 0 15 9 2
16 7 2 10 0 9 13 1 10 9 10 0 9 10 0 9 2
8 7 2 13 3 10 9 9 2
80 10 0 9 2 1 10 9 10 12 9 9 2 10 15 13 0 1 15 10 9 3 1 10 9 2 7 1 10 0 9 15 13 1 9 2 13 1 9 10 0 9 1 9 10 9 2 7 13 0 9 3 10 7 15 13 1 9 2 3 1 10 12 2 10 9 1 10 15 13 7 10 0 9 13 10 9 15 15 13 2
28 1 10 0 9 2 0 14 13 1 10 9 12 10 9 2 10 9 3 15 15 14 13 3 1 10 9 12 2
10 14 13 14 13 10 0 9 15 3 2
7 0 9 13 7 15 9 2
11 13 7 10 0 9 7 13 1 0 9 2
13 3 1 12 9 9 10 9 13 9 10 0 9 2
18 13 1 10 0 10 9 9 7 3 1 9 12 9 13 1 0 9 2
86 10 9 1 10 0 9 7 9 7 10 0 9 2 10 9 2 10 0 9 13 10 9 15 13 3 3 9 2 10 9 10 9 9 2 9 10 0 0 9 2 10 9 2 10 9 2 13 3 1 9 10 2 0 9 2 15 13 13 10 9 9 12 9 2 10 9 9 10 9 2 10 9 9 7 10 9 13 15 3 1 10 0 9 10 9 2
30 10 0 9 13 0 9 10 0 9 2 7 15 1 10 9 15 13 1 9 10 9 9 2 13 9 1 9 9 9 2
24 10 9 9 13 1 9 15 7 2 10 9 15 13 1 0 9 15 15 13 14 13 10 0 2
31 9 10 9 13 10 9 10 9 7 10 9 9 2 3 3 7 10 9 10 9 2 10 15 13 3 1 14 13 9 9 2
30 15 13 10 9 10 9 1 9 7 10 9 10 9 9 1 9 2 10 0 9 10 15 13 3 1 10 9 10 9 2
25 0 15 13 1 9 10 9 7 10 9 2 1 10 9 7 13 1 9 1 10 9 9 7 9 2
16 7 2 10 0 9 14 13 10 0 9 1 10 9 0 9 2
7 10 9 15 14 13 0 2
20 14 13 0 14 13 3 0 3 13 3 9 2 7 3 9 9 13 10 9 2
24 10 9 10 9 2 7 9 2 2 10 12 0 9 1 9 2 13 10 9 15 1 9 9 2
64 10 9 10 9 13 1 9 2 12 1 10 3 0 9 10 9 2 1 9 12 2 1 10 9 2 13 3 1 9 7 3 1 10 0 9 10 9 10 0 9 10 9 2 12 1 10 3 0 9 10 9 2 15 13 10 9 10 9 1 10 0 0 9 2
14 7 3 7 3 10 12 9 9 13 9 3 1 15 2
23 15 13 10 0 13 9 2 7 10 9 14 13 3 13 10 9 9 10 12 9 10 9 2
23 7 2 13 0 10 9 7 10 13 9 0 9 13 10 9 2 3 3 1 10 9 9 2
24 3 13 10 2 9 2 7 2 10 9 13 14 13 0 10 9 2 3 1 10 9 10 9 2
40 13 7 10 9 14 15 13 0 9 7 7 14 13 14 13 0 9 10 12 9 2 1 0 9 14 14 13 1 9 10 0 9 7 1 9 10 14 13 0 2
16 3 7 1 10 9 10 9 10 9 13 9 9 0 9 9 2
20 15 10 9 13 14 13 9 10 9 10 0 9 1 15 10 9 10 0 9 2
19 10 9 7 10 9 13 0 7 0 9 2 1 9 10 9 10 0 9 2
13 3 13 3 14 13 9 3 1 10 9 10 9 2
5 1 9 10 9 2
1 9
14 1 9 2 13 10 9 7 13 10 9 9 14 13 2
34 10 0 0 9 15 13 1 10 9 14 13 9 10 9 10 9 2 13 10 9 9 1 10 9 9 9 1 10 9 10 9 9 9 2
59 10 9 10 0 9 9 1 10 0 9 9 2 10 9 15 7 10 9 1 9 0 9 2 9 2 9 2 2 10 15 13 1 10 9 10 9 7 13 0 10 9 2 13 10 9 1 10 15 10 9 10 9 13 7 3 13 10 9 2
30 9 9 2 3 14 13 14 13 10 12 9 2 10 2 9 2 10 2 9 9 7 10 2 9 2 1 10 9 15 2
73 13 14 13 14 13 3 2 13 7 14 13 3 13 2 10 9 15 13 3 7 14 13 14 13 7 1 10 9 10 9 10 9 14 13 10 0 9 2 14 13 10 9 7 3 14 13 1 3 1 9 2 9 2 9 7 9 2 9 9 0 2 9 1 10 15 15 15 14 14 13 14 13 2
7 3 15 13 13 1 9 2
20 10 9 15 14 13 14 13 7 14 13 0 3 1 10 9 10 9 1 9 2
12 15 13 3 15 15 14 14 13 14 13 0 2
27 10 9 10 0 9 1 9 13 1 9 9 2 10 0 9 13 3 3 7 10 9 9 0 9 13 9 2
28 10 9 10 9 15 13 14 13 1 9 1 10 9 7 14 13 7 10 12 13 10 9 10 9 0 10 9 2
21 1 0 9 13 3 2 3 13 2 14 13 0 9 9 1 9 0 7 0 9 2
22 3 13 10 9 3 2 7 14 14 13 3 3 0 7 14 13 10 9 0 0 9 2
35 1 10 9 10 9 10 0 9 1 10 9 2 10 9 13 1 9 10 9 3 7 3 13 9 1 9 7 13 9 1 10 9 0 9 2
6 14 13 14 15 13 2
32 1 10 9 15 13 14 13 7 1 0 9 14 14 13 0 10 9 10 9 1 10 9 1 0 9 9 15 13 9 7 9 2
12 3 2 10 9 13 0 9 1 7 10 9 2
24 10 9 9 13 1 0 9 15 13 13 10 9 1 9 9 7 13 9 1 10 9 10 9 2
15 10 9 15 13 14 13 1 9 10 0 9 9 1 2 2
36 1 9 2 10 9 9 7 9 13 1 10 9 9 10 9 15 14 13 10 9 9 1 10 9 10 0 9 1 0 9 3 1 10 9 9 2
24 3 10 12 9 13 10 9 15 2 10 15 7 13 1 0 9 1 10 9 15 2 10 9 2
39 3 2 7 7 13 3 1 10 0 0 9 2 3 13 1 10 9 9 1 10 9 15 13 10 9 15 2 2 9 2 13 3 1 10 9 0 9 9 2
30 13 3 14 13 1 9 10 9 10 9 2 10 9 2 7 14 13 10 9 1 15 10 9 1 9 10 9 10 9 2
11 10 9 15 13 3 1 10 9 10 9 2
30 3 2 3 13 10 0 13 10 9 2 10 15 13 10 9 10 9 2 7 14 13 13 13 9 1 10 9 10 9 2
4 1 9 9 2
27 10 9 13 1 9 9 2 9 2 1 15 10 12 9 13 1 0 9 1 0 9 2 3 1 9 9 2
33 10 12 13 3 0 9 10 9 7 10 9 9 7 9 1 9 9 2 10 12 10 9 9 7 3 10 12 10 0 9 1 9 2
31 13 15 13 1 10 9 7 15 13 14 13 10 9 15 1 10 9 9 10 9 2 7 13 14 13 10 9 1 12 9 2
10 10 2 13 0 9 1 9 10 9 2
30 1 9 13 10 9 14 13 1 0 0 7 14 13 1 0 9 9 0 0 9 1 9 9 2 9 7 1 9 9 2
5 10 9 13 3 2
20 10 9 2 10 15 13 10 9 2 13 3 12 9 1 0 1 12 9 9 2
6 10 0 9 13 13 2
1 9
27 14 13 14 15 13 1 15 7 14 15 13 14 13 14 13 10 9 15 1 0 15 9 15 10 12 9 2
14 10 0 9 13 14 13 3 1 10 9 10 0 9 2
20 1 15 10 9 13 7 10 9 10 3 9 9 9 9 1 9 2 1 9 2
23 3 10 9 9 9 9 13 13 10 0 9 2 13 7 3 1 9 14 13 1 15 9 2
15 10 9 15 13 3 10 9 2 7 7 13 10 0 9 2
18 10 9 13 3 1 9 7 9 15 13 3 1 10 9 15 10 9 2
24 3 3 7 13 1 12 9 9 2 14 13 14 13 10 9 15 13 1 10 9 10 9 15 2
19 1 3 13 3 1 0 9 0 9 9 1 7 1 0 9 10 0 9 2
37 3 2 1 9 2 10 9 9 15 14 13 9 9 1 9 0 9 7 9 0 9 7 0 9 0 9 13 0 7 13 9 1 9 10 0 9 2
25 10 9 1 9 13 10 9 14 13 10 9 15 1 10 9 7 10 9 14 13 9 3 1 15 2
24 10 9 9 1 9 1 10 0 9 2 10 9 7 10 9 15 13 10 9 2 13 10 9 2
26 7 13 14 13 1 9 2 13 0 9 1 15 1 0 9 10 9 2 1 9 1 12 0 0 9 2
20 7 13 14 13 1 9 3 2 13 0 14 13 7 10 9 13 1 10 9 2
37 15 13 3 1 10 9 15 2 15 14 13 7 1 10 9 15 10 0 9 15 13 10 9 15 7 10 0 9 15 13 1 10 9 10 3 9 2
6 13 7 15 13 0 2
35 13 3 7 3 1 10 0 9 9 2 9 7 9 2 10 9 9 13 14 13 14 13 10 9 7 14 13 10 0 9 1 0 15 9 2
32 10 0 15 9 13 1 9 15 7 10 9 15 13 1 9 10 9 9 7 9 13 14 13 1 0 10 9 9 10 2 3 2
24 1 0 9 10 9 13 9 1 10 9 9 9 1 9 2 1 10 9 7 9 15 1 9 2
95 9 9 2 1 10 9 10 0 9 13 0 9 2 10 15 13 3 1 10 9 10 9 2 3 7 10 0 9 2 7 7 1 9 0 9 2 9 7 9 13 10 9 7 0 15 10 9 2 13 3 7 10 9 9 10 15 3 13 3 13 10 0 9 2 10 15 13 2 13 9 3 7 13 10 0 9 1 10 9 9 2 3 1 10 9 10 9 7 3 1 10 9 10 9 2
15 10 9 10 9 13 15 10 9 1 9 15 13 1 9 2
60 7 10 9 13 3 0 7 0 9 1 10 9 10 9 10 9 3 13 7 1 10 9 0 9 2 3 14 14 13 10 0 9 9 2 7 3 14 3 3 10 9 13 10 12 9 10 0 9 2 13 3 7 15 13 3 0 3 7 0 2
23 12 1 10 9 14 13 15 2 7 10 9 10 9 7 10 9 9 13 1 10 13 9 2
21 10 9 13 10 13 9 10 9 14 13 10 9 7 15 13 13 1 10 0 9 2
32 3 2 13 3 7 13 14 13 10 9 10 9 7 10 9 15 7 1 0 9 15 13 14 13 10 0 9 7 14 10 9 2
14 10 9 14 13 1 9 10 9 10 9 15 14 13 2
5 13 10 9 9 2
8 10 9 10 9 13 14 13 2
17 1 9 7 1 9 15 2 13 10 0 9 10 9 7 10 9 2
7 9 1 9 13 10 9 9
33 1 9 2 14 13 15 3 10 9 1 10 9 15 13 10 9 7 13 0 9 1 9 2 1 0 7 0 9 1 10 0 9 2
20 14 15 13 7 13 15 10 9 10 9 2 7 14 13 10 9 2 13 3 2
8 13 10 9 9 0 7 0 2
18 13 14 13 10 9 2 9 9 10 9 2 13 1 10 9 10 9 2
24 10 9 10 0 9 9 9 2 15 13 1 10 0 13 10 9 15 13 10 9 2 9 2 2
21 10 9 14 13 14 13 1 9 15 7 0 9 7 13 10 9 15 13 10 9 2
10 3 2 14 13 14 13 12 3 9 2
16 13 7 14 13 3 15 10 9 7 13 10 9 1 0 9 2
24 7 2 10 0 0 13 7 13 14 13 3 10 9 1 10 9 0 0 9 1 0 10 9 2
22 3 2 10 0 9 1 0 9 14 13 14 13 3 9 2 13 10 9 15 10 9 2
22 3 1 9 2 10 9 14 13 3 14 13 0 10 9 0 10 9 2 13 7 14 2
49 10 9 9 10 9 10 9 0 0 2 9 7 9 14 13 3 14 15 13 2 3 3 13 10 0 9 2 3 13 10 9 10 9 1 9 2 10 9 9 10 9 2 7 10 0 7 10 0 2
22 10 9 10 9 13 1 9 9 2 3 1 9 10 2 7 10 2 7 1 0 9 2
30 12 9 3 2 10 9 13 10 12 9 7 12 9 1 10 9 10 9 10 9 9 13 10 9 10 9 3 1 9 2
19 10 0 9 13 1 0 9 9 9 0 9 2 0 9 7 9 9 9 2
26 3 1 9 2 10 12 10 9 13 7 10 0 9 13 7 10 0 12 13 7 14 13 15 0 9 2
28 10 0 9 13 14 13 0 15 0 9 7 13 15 10 0 14 13 15 9 9 1 14 13 14 13 0 9 2
39 10 9 13 7 1 9 1 10 9 10 9 13 0 9 1 10 0 0 2 0 7 0 9 10 9 9 2 7 14 13 1 9 10 9 9 1 0 9 2
25 10 12 9 10 9 13 1 9 10 9 7 10 0 9 2 3 1 10 9 2 13 1 0 9 2
11 3 2 10 9 13 14 13 10 3 3 2
12 10 9 13 2 3 13 2 14 13 1 15 2
20 10 9 10 9 7 10 9 13 7 10 9 14 14 13 10 9 10 12 9 2
69 14 13 14 13 10 9 0 10 9 1 9 7 2 7 13 15 9 10 15 13 0 9 1 10 9 10 9 10 0 9 2 3 1 10 9 3 10 0 15 2 10 9 10 9 1 15 9 7 1 10 9 12 9 2 3 7 10 9 9 2 13 0 1 10 9 10 9 15 2
10 3 2 0 10 9 13 10 0 9 2
35 3 13 7 10 9 2 9 15 3 13 3 3 9 14 13 1 0 9 10 9 15 14 13 3 1 9 10 9 2 3 7 10 9 9 2
26 1 12 9 2 10 9 13 12 9 1 10 9 9 9 2 12 9 2 7 9 9 2 12 9 2 2
44 10 9 9 13 10 9 7 2 10 9 9 13 1 10 9 10 9 2 9 9 2 7 10 9 9 2 9 9 2 7 15 13 10 0 15 9 1 9 9 9 1 0 9 2
59 15 7 14 13 10 9 9 1 9 2 1 9 10 12 9 13 10 9 15 13 3 1 10 9 9 7 9 1 10 9 9 3 2 7 1 10 9 10 2 2 10 9 7 10 9 1 9 1 10 9 2 10 9 7 10 9 1 9 2
17 13 0 9 10 9 10 9 14 13 3 0 15 9 10 0 9 2
22 15 2 3 9 2 13 10 9 10 0 0 9 2 7 3 7 10 9 15 14 13 2
24 10 9 9 13 10 9 9 7 15 10 9 9 9 2 15 13 1 9 9 9 1 10 9 2
9 13 1 0 9 1 10 0 9 2
26 10 9 15 14 3 14 13 10 9 10 9 1 9 15 7 14 13 3 10 0 9 1 10 9 9 2
11 13 14 13 7 3 10 9 1 10 9 2
34 10 9 10 9 9 2 9 9 9 2 13 10 9 7 2 7 10 9 13 14 13 10 9 1 9 2 14 13 14 13 7 10 9 2
28 13 14 13 0 10 9 14 13 10 9 2 3 13 10 2 9 2 7 14 13 10 12 2 14 13 1 9 2
32 1 10 9 15 13 10 9 14 13 1 0 10 9 14 13 10 0 9 1 9 3 7 14 13 7 14 13 10 0 0 9 2
27 10 9 15 13 1 9 10 9 10 9 14 13 1 9 10 9 0 1 9 9 3 7 1 0 0 9 2
16 12 0 9 2 9 12 9 2 10 9 9 13 3 1 9 2
43 10 9 12 10 9 2 3 13 1 9 10 9 9 1 9 2 15 13 3 1 15 0 9 1 9 1 10 9 9 7 9 1 10 9 10 9 15 3 9 15 10 9 2
48 10 9 9 13 7 2 3 13 0 9 1 9 1 10 9 2 7 13 15 9 2 13 1 9 10 9 7 13 10 9 10 9 2 1 15 13 10 0 9 1 10 9 10 0 15 9 2 2
11 13 2 13 2 14 13 10 9 10 9 2
26 10 0 9 10 9 15 13 10 9 10 9 9 9 2 9 2 13 9 2 9 2 9 7 13 9 2
13 13 14 13 9 15 14 13 10 9 7 10 9 2
26 10 9 10 9 1 9 10 9 13 1 0 9 15 2 10 15 13 3 1 10 12 1 10 12 9 2
28 10 9 13 3 1 0 9 7 3 1 15 13 14 13 10 9 10 9 14 13 10 9 3 3 1 10 9 2
43 1 10 9 10 9 7 10 9 10 2 1 10 9 10 9 13 10 9 1 10 15 9 10 0 9 13 10 9 14 13 1 9 9 1 9 10 2 2 9 0 9 2 2
12 1 9 15 12 7 12 13 0 9 1 9 2
26 3 2 10 0 9 9 10 9 14 13 10 9 7 10 9 13 7 13 14 13 1 9 10 0 9 2
41 7 13 7 3 3 14 13 14 13 15 9 2 7 15 14 13 14 13 3 1 10 0 9 2 14 13 10 0 2 0 9 2 2 3 15 15 14 13 14 13 2
24 10 9 13 3 1 10 0 9 2 13 3 1 10 9 2 1 0 9 7 13 10 0 9 2
14 10 9 13 12 9 1 9 3 0 10 12 2 9 2
20 10 12 9 13 13 1 9 7 9 7 13 0 2 7 14 13 9 1 9 2
24 10 9 9 10 9 14 13 3 1 10 9 2 14 13 7 14 13 10 9 1 0 10 9 2
20 10 0 9 9 10 2 13 3 1 9 15 1 9 2 10 9 7 10 9 2
25 10 9 10 9 7 10 9 14 13 0 9 14 13 10 9 1 10 9 10 9 1 9 10 9 2
28 13 15 2 9 9 2 14 13 10 12 9 10 0 9 15 15 13 1 12 9 2 1 10 9 15 10 9 2
12 10 9 13 10 12 0 9 1 10 0 9 2
17 15 13 3 2 13 10 9 7 10 0 9 2 7 13 3 0 2
22 1 10 9 13 9 2 7 9 13 10 0 9 3 10 0 1 10 3 9 10 9 2
29 3 13 13 3 1 9 10 0 9 1 9 2 10 15 13 3 7 0 9 1 9 15 13 1 9 10 0 9 2
25 10 9 13 10 9 7 13 9 9 2 0 9 9 2 9 0 9 2 9 9 7 9 9 9 2
50 3 2 3 13 10 9 10 9 1 10 3 10 9 14 13 14 13 1 9 2 10 9 1 9 12 13 0 7 13 3 13 7 10 0 9 14 13 10 9 10 0 9 1 9 7 1 9 7 9 2
12 13 1 9 2 10 9 13 9 10 0 9 2
30 10 9 13 7 2 10 9 13 3 9 9 1 9 1 3 12 9 7 13 1 0 7 0 9 1 9 9 15 2 2
32 3 13 2 13 7 13 10 12 9 10 0 9 7 13 10 9 10 9 1 10 9 9 2 9 9 2 9 7 9 10 9 2
22 3 12 9 13 1 10 9 10 9 15 13 3 1 9 10 0 0 9 10 0 9 2
48 15 13 14 14 13 1 9 10 1 9 9 7 2 1 9 1 10 15 15 13 2 15 10 9 9 10 9 13 2 1 10 9 10 9 0 9 2 0 2 9 10 15 13 1 9 14 13 2
17 3 2 9 13 7 1 10 0 9 9 2 9 2 9 7 9 2
1 9
1 9
26 10 0 9 14 13 14 13 10 9 1 10 9 9 14 13 0 9 1 10 9 7 14 13 10 9 2
2 12 2
55 3 1 0 9 13 14 13 10 9 15 1 12 3 9 2 7 13 14 13 10 0 1 10 9 9 1 9 7 9 7 13 1 9 7 9 9 2 9 7 0 9 14 13 3 1 9 15 14 13 10 0 9 1 9 2
47 10 9 13 3 7 10 0 9 15 13 13 1 9 10 0 9 14 13 1 10 0 7 0 9 10 0 9 3 1 9 9 15 15 13 1 12 9 3 1 10 0 9 10 9 10 9 2
32 3 14 13 1 0 9 2 7 1 9 3 10 9 1 10 15 0 9 13 10 0 10 9 3 13 10 9 7 10 9 9 2
9 13 14 13 3 0 3 1 15 2
31 10 2 9 9 13 3 14 13 0 9 7 3 14 13 13 14 13 10 0 9 13 1 10 9 10 9 1 10 9 9 2
64 10 9 9 13 7 2 3 3 10 9 13 13 14 13 15 13 15 13 15 1 10 0 9 14 15 13 2 7 13 7 2 15 14 14 13 3 1 9 10 0 9 2 7 14 13 7 10 0 2 2 7 13 7 2 1 10 12 14 13 9 1 0 2 2
19 0 0 9 2 3 10 9 10 9 9 1 0 9 2 13 1 0 9 2
28 3 13 14 13 12 9 2 9 15 13 1 9 9 12 2 10 0 9 7 13 15 7 10 9 13 14 13 2
34 10 9 10 0 9 1 9 13 3 0 9 2 3 9 13 14 13 10 9 1 0 0 9 10 9 15 10 9 10 0 7 0 9 2
5 1 9 10 9 2
37 1 10 9 10 9 10 9 2 3 13 10 9 10 2 9 2 13 13 1 10 0 9 15 13 7 10 0 13 7 1 10 9 10 2 9 9 2
22 13 7 14 13 14 13 0 1 15 10 9 14 13 3 10 9 10 9 1 0 9 2
19 10 9 1 10 9 9 10 0 9 14 13 1 9 10 9 10 9 15 2
39 10 9 13 0 7 13 1 10 9 1 10 15 3 14 13 0 9 2 7 14 13 10 0 7 0 9 9 10 9 2 7 9 15 13 1 10 0 9 2
27 10 9 15 13 3 10 9 2 3 1 10 9 2 10 9 2 10 9 7 10 0 9 13 9 0 9 2
17 1 9 10 9 2 10 9 13 0 9 1 0 1 15 0 9 2
15 15 10 9 13 1 9 10 9 1 0 9 10 9 9 2
31 13 1 3 1 9 10 9 9 9 9 3 1 10 9 1 10 0 9 7 1 0 9 9 2 1 10 15 13 3 9 2
24 1 12 2 10 9 13 14 13 2 7 10 9 1 10 9 10 9 13 10 12 9 10 9 2
68 9 10 9 9 10 9 10 9 13 1 9 2 1 9 2 1 3 13 10 12 2 12 0 9 2 13 10 9 9 2 13 10 9 1 9 10 9 2 13 3 1 0 9 7 9 7 13 10 9 10 9 2 7 14 13 14 13 1 10 9 15 10 9 14 13 10 9 2
29 10 0 0 1 10 9 10 0 9 2 9 9 2 13 3 9 10 0 9 1 0 0 9 10 9 7 10 9 2
12 9 2 12 9 13 3 1 9 10 0 1 9
15 10 9 10 0 9 9 2 9 7 9 13 0 1 9 2
14 13 15 3 14 13 7 10 9 3 1 10 9 9 2
43 13 3 3 10 9 15 1 9 2 1 15 13 10 9 10 0 9 15 13 3 9 1 10 9 7 13 10 9 10 15 13 1 0 9 10 9 15 13 3 1 0 9 2
24 7 14 13 3 1 10 9 15 7 14 13 14 13 0 10 0 9 2 3 7 10 0 9 2
45 1 14 15 13 3 2 10 0 9 3 1 10 0 9 15 13 9 1 10 9 3 7 10 0 9 1 13 9 3 13 7 10 0 13 14 14 13 9 1 10 15 14 13 9 2
7 13 0 9 3 1 15 2
16 14 13 14 13 7 10 9 15 13 1 0 7 1 0 9 2
28 0 9 2 1 10 15 14 13 7 10 0 9 2 13 14 13 1 9 3 3 13 13 14 13 1 10 9 2
25 10 0 0 9 10 0 9 13 7 2 13 9 1 10 9 9 1 3 0 9 0 1 9 2 2
24 1 10 9 2 10 9 7 10 0 9 2 10 9 13 1 9 7 9 2 10 9 10 9 2
7 13 0 9 1 0 9 2
18 1 9 10 9 2 1 9 2 13 9 2 10 0 9 10 15 13 2
57 10 9 15 2 9 9 2 9 2 3 14 13 0 3 9 9 2 2 13 0 1 10 0 15 9 2 7 7 10 0 9 13 14 13 1 9 7 13 10 9 10 9 10 2 1 10 0 2 3 3 13 1 10 0 0 9 2
54 10 9 7 2 3 10 13 0 9 13 7 0 9 3 1 3 15 3 0 13 0 2 7 1 10 9 10 0 9 1 9 2 2 9 2 2 2 10 0 9 2 9 15 3 9 2 2 10 0 9 13 14 13 2
23 10 9 15 13 10 9 9 13 1 9 14 13 10 9 15 7 13 10 9 10 12 9 2
97 10 3 3 15 13 14 13 13 14 13 10 9 15 1 9 10 9 2 3 1 15 1 10 9 1 9 2 1 0 9 14 2 13 2 2 7 14 15 13 2 10 9 10 9 15 2 7 14 13 0 14 13 12 7 0 1 10 9 10 0 9 15 14 13 14 13 10 9 2 10 9 2 10 9 2 10 9 2 3 7 10 0 9 2 3 10 9 14 13 0 9 14 13 7 3 0 2
39 1 14 13 10 9 1 9 10 9 2 14 13 14 13 10 9 1 9 1 10 9 9 1 10 9 9 2 1 10 13 1 9 9 7 1 9 1 9 2
44 10 9 9 9 13 3 7 2 9 9 1 9 9 1 10 2 7 10 0 9 13 14 13 1 0 9 1 14 13 10 9 9 1 10 9 12 9 9 1 9 1 9 2 2
16 3 2 10 0 0 9 13 0 9 1 10 0 0 9 2 2
26 15 13 1 10 9 2 10 9 2 10 9 9 9 2 10 9 2 10 9 9 1 0 10 0 9 2
48 10 9 15 13 1 10 0 9 2 7 13 7 10 9 15 1 15 2 13 14 13 1 9 10 0 9 2 1 14 13 1 9 15 15 0 9 15 14 13 3 3 3 10 9 10 0 9 2
17 13 7 10 9 15 13 14 14 13 3 9 7 0 9 1 9 2
24 3 2 10 9 15 2 15 13 2 13 10 0 9 10 9 0 10 9 9 1 9 9 9 2
28 3 14 13 14 13 7 1 10 9 15 13 3 0 7 13 7 10 0 9 7 14 13 9 1 10 0 9 2
25 10 9 14 13 10 9 2 3 15 13 10 0 9 7 10 9 1 15 13 13 3 1 0 9 2
38 1 3 2 10 9 13 7 2 14 13 1 9 10 9 9 1 10 9 7 1 15 9 15 14 13 10 9 9 14 13 0 0 9 9 1 9 2 2
15 1 0 1 12 0 9 2 10 9 15 14 13 14 13 2
14 10 0 9 14 13 0 9 7 13 10 0 9 15 2
7 13 14 13 10 9 15 2
4 13 13 9 2
18 13 10 9 1 10 15 0 15 14 13 7 13 14 13 0 0 9 2
15 10 9 13 0 9 1 10 9 7 10 9 10 0 9 2
44 13 7 1 10 0 9 14 13 7 14 13 10 0 9 10 0 9 9 1 9 10 9 7 1 9 10 9 7 7 10 0 9 14 13 9 1 10 0 9 10 9 1 9 2
31 9 1 0 9 13 1 10 9 14 13 9 1 9 9 2 7 10 0 9 14 15 13 10 9 1 9 2 0 9 9 2
11 10 0 9 2 1 9 2 13 0 9 2
30 13 2 9 9 2 9 7 9 9 2 10 0 9 15 13 10 9 14 13 10 9 3 1 10 9 10 9 1 9 2
23 10 9 15 0 9 1 9 15 13 10 9 15 2 13 0 9 7 1 9 7 1 9 2
29 1 12 0 9 9 1 10 9 1 10 9 13 1 0 9 15 13 0 9 2 7 13 10 9 1 3 12 9 2
36 10 9 15 10 0 9 13 7 10 9 10 9 10 9 15 13 0 3 0 2 7 1 9 3 14 13 10 9 14 13 1 9 10 0 9 2
28 13 10 0 9 14 14 13 15 9 3 1 10 9 10 9 2 7 14 13 7 10 9 13 10 9 10 9 2
9 10 3 3 13 15 15 13 3 2
8 3 12 9 13 10 9 15 2
18 10 0 9 10 9 13 10 9 15 7 14 13 10 0 9 1 9 2
9 10 9 15 13 1 9 10 2 2
20 10 9 13 0 7 13 7 13 12 9 1 9 9 2 7 13 3 12 9 2
5 10 9 15 13 2
15 13 7 7 13 3 0 14 13 0 9 1 10 9 15 2
34 1 10 9 15 2 13 10 0 9 1 12 3 0 9 2 1 9 10 0 9 7 1 9 3 10 3 9 13 14 13 0 0 9 2
11 12 0 1 10 0 9 15 13 10 9 2
25 13 1 9 9 12 9 2 3 7 1 9 0 1 9 10 9 2 7 13 9 9 12 2 9 2
17 10 9 13 7 14 13 14 13 9 2 7 10 9 14 13 3 2
46 10 15 9 1 15 13 13 13 10 9 10 9 14 13 0 9 3 1 10 9 1 10 9 2 10 15 13 0 2 14 3 1 10 0 9 10 9 7 7 1 10 9 1 9 9 2
19 10 9 14 13 1 9 7 15 13 13 14 3 10 9 7 7 10 9 2
12 10 0 9 10 9 13 10 9 10 9 9 2
54 10 9 3 13 14 13 10 0 9 10 15 14 13 1 0 9 2 3 13 10 9 10 9 2 7 3 14 13 10 9 10 9 2 10 15 1 10 9 15 13 0 9 2 0 0 9 2 0 0 9 2 0 9 2
11 14 13 2 3 2 10 9 10 0 9 2
23 1 15 10 9 2 10 0 9 10 9 13 14 13 9 1 9 2 13 10 9 10 9 2
12 0 15 10 9 14 13 14 13 10 0 9 2
21 10 9 9 13 0 3 7 9 1 9 14 13 14 13 0 9 7 13 9 15 2
38 10 2 9 13 10 9 15 1 0 1 10 9 15 13 13 1 15 9 7 13 14 15 13 1 0 9 2 0 9 2 9 9 2 0 9 7 15 2
19 1 10 0 9 10 9 10 9 13 7 13 10 9 7 10 9 10 9 2
16 1 9 13 7 10 0 9 10 9 2 10 15 13 10 9 2
39 10 9 1 10 9 14 13 10 9 10 9 2 7 14 13 2 3 9 10 9 15 2 0 9 1 10 9 10 13 9 1 9 2 13 3 10 0 9 2
30 13 10 12 9 3 10 0 9 13 1 0 9 14 13 10 9 9 1 10 9 9 2 3 13 10 0 9 10 9 2
20 1 10 0 12 2 10 12 13 7 13 1 9 0 7 12 1 9 0 9 2
27 14 13 14 13 10 9 2 10 9 15 13 3 1 10 0 9 7 13 10 0 9 10 9 1 10 9 2
4 10 9 9 2
12 14 13 3 14 13 0 14 13 3 0 9 2
27 10 9 13 1 10 9 9 2 10 15 13 9 9 10 9 12 7 0 9 10 9 9 1 10 9 12 2
16 13 10 0 9 10 9 2 15 13 10 0 9 10 0 9 2
12 12 2 9 9 2 10 9 13 9 1 10 9
9 13 9 10 0 9 9 10 2 2
23 10 9 9 10 12 0 9 13 10 9 2 9 15 1 10 9 13 10 9 10 9 15 2
10 13 10 0 9 7 9 10 0 9 2
40 10 9 9 1 10 0 9 15 13 0 9 7 13 7 3 1 0 15 9 1 10 9 10 9 10 9 9 14 13 1 15 10 9 15 10 9 1 10 9 2
65 3 13 14 13 2 1 9 10 9 2 7 1 10 0 15 9 14 13 14 13 3 14 13 10 0 9 9 7 1 10 0 9 2 7 10 9 15 13 9 10 0 9 2 10 15 1 10 9 15 14 13 13 15 9 9 3 1 10 3 14 13 10 9 9 2
8 10 9 10 9 13 0 9 2
21 0 7 0 9 2 9 2 0 9 2 9 2 0 9 2 9 2 9 2 9 2
25 15 9 2 13 3 1 10 0 9 2 3 13 12 7 12 9 9 9 2 0 1 10 0 9 2
4 1 9 9 2
14 13 15 14 13 12 9 10 9 15 1 15 10 9 2
15 1 9 13 10 9 10 0 9 1 0 9 10 0 9 2
16 10 9 13 7 13 10 0 9 1 10 9 9 1 10 9 2
21 14 13 0 9 9 7 3 10 9 14 13 10 0 7 0 9 1 10 0 9 2
31 7 7 10 9 13 15 9 7 9 7 13 14 13 9 0 9 2 10 9 13 14 13 10 0 9 0 2 0 7 0 2
15 10 0 9 13 1 9 1 9 1 10 0 0 9 9 2
55 14 15 13 14 13 1 12 7 12 0 9 2 10 9 2 15 13 10 0 2 10 0 9 10 9 1 3 2 7 3 2 3 13 7 15 2 10 0 9 10 9 2 7 14 13 1 0 9 1 10 9 10 0 9 2
17 3 2 3 1 9 9 2 0 9 2 13 10 0 9 10 9 2
29 0 9 13 7 2 10 9 9 10 2 13 0 9 7 14 15 13 14 13 1 10 9 3 13 10 9 15 2 2
26 3 2 1 15 10 12 9 2 10 9 9 13 3 10 9 10 9 2 13 10 0 1 10 0 9 2
36 10 9 9 13 1 3 3 10 9 0 9 1 14 13 10 9 2 1 7 14 13 14 13 10 9 2 1 9 14 13 13 12 9 7 9 2
13 13 3 7 1 10 9 15 13 3 10 9 15 2
14 10 9 13 9 14 13 10 9 9 9 1 0 9 2
60 13 7 10 0 9 14 13 10 0 9 15 13 10 9 10 9 2 10 0 9 2 10 9 1 0 9 2 10 9 7 10 9 10 9 2 10 9 1 10 9 10 9 2 10 0 9 1 10 9 10 9 7 10 0 9 10 9 0 9 2
44 7 1 0 9 10 9 9 10 9 13 0 9 7 13 3 0 2 7 14 13 3 13 0 14 13 14 13 3 3 10 0 9 1 10 0 9 15 13 1 9 15 9 9 2
22 10 9 15 13 0 10 9 9 1 9 10 9 2 1 10 0 9 7 9 15 13 2
33 3 13 1 0 9 1 10 3 0 9 2 1 10 9 7 10 9 2 14 13 10 9 7 10 9 10 9 9 0 1 10 9 2
12 9 9 13 10 0 9 10 9 1 0 9 2
17 7 14 13 0 0 2 7 14 13 13 1 10 9 3 10 9 2
19 1 10 9 13 9 1 10 9 10 9 2 10 15 13 10 0 0 9 2
11 3 13 3 15 9 9 7 15 9 9 2
30 9 10 9 9 1 9 13 7 2 1 10 9 13 7 12 9 2 7 10 0 13 9 2 9 2 9 7 9 2 2
15 7 15 13 10 9 3 13 2 14 13 3 14 15 13 2
31 10 0 13 7 15 14 13 14 15 13 1 10 13 10 9 15 1 9 2 3 1 10 9 7 0 9 15 13 10 9 2
20 1 10 9 10 9 3 9 2 12 1 12 9 13 7 10 0 9 14 13 2
11 13 10 9 15 1 9 9 7 0 9 2
26 13 13 14 13 9 3 1 2 14 13 1 15 9 10 9 15 13 13 1 9 3 1 10 9 9 2
34 13 0 7 10 0 9 1 10 9 10 0 9 13 14 13 7 14 13 1 10 9 9 7 0 9 10 9 15 13 13 1 10 9 2
18 7 10 9 13 1 15 2 13 14 13 10 9 14 13 9 1 9 2
15 15 13 7 0 9 15 13 0 7 0 1 9 9 9 2
21 13 10 0 9 15 1 15 13 10 2 9 7 13 14 15 13 1 10 9 15 2
13 3 3 2 1 9 13 12 9 9 1 12 9 2
25 14 13 3 1 10 9 10 9 10 9 2 13 2 7 2 0 9 1 10 9 10 9 10 9 2
51 1 9 13 0 7 7 1 0 9 9 9 2 3 7 1 0 9 9 2 14 13 0 7 0 9 2 10 15 13 7 14 13 1 9 7 1 10 0 9 3 7 1 9 9 9 1 10 0 9 9 2
11 3 2 13 3 9 1 0 9 10 9 2
63 10 0 9 10 12 9 1 10 0 9 14 3 13 0 9 9 1 14 13 10 9 10 9 1 9 1 10 9 15 9 0 9 2 7 3 13 10 9 15 13 14 13 10 9 10 9 1 10 15 13 14 13 10 9 9 9 1 15 13 10 9 15 2
26 10 9 13 0 14 13 10 0 2 0 9 2 10 0 9 2 3 15 13 3 10 2 7 10 9 2
22 10 9 2 12 13 3 0 1 0 9 9 15 13 1 9 7 13 1 0 10 9 2
16 15 10 9 13 10 0 7 3 0 9 1 14 13 0 15 2
31 2 1 10 9 1 9 14 13 1 10 9 9 10 9 14 15 13 14 13 10 9 1 12 9 2 2 13 10 9 9 2
16 10 9 15 13 10 12 7 9 1 10 9 10 9 1 9 2
88 14 13 14 13 10 9 15 13 10 0 9 2 7 2 7 13 13 10 9 10 9 10 9 10 9 7 10 9 10 9 15 13 0 1 9 2 14 13 13 10 9 9 1 10 9 7 10 9 2 9 15 13 7 10 12 0 9 7 13 2 3 2 0 0 0 9 2 7 7 10 9 13 3 13 9 14 12 9 10 0 15 9 2 3 1 10 9 2
8 2 10 9 10 9 13 0 2
9 10 9 15 13 10 12 0 9 2
39 13 10 9 9 15 13 10 9 10 9 10 0 2 0 0 9 2 15 13 14 13 7 10 9 10 0 9 9 13 1 10 9 0 0 9 1 0 9 2
38 10 15 9 10 9 13 10 2 2 10 15 13 10 0 9 9 7 0 9 2 15 13 1 10 9 2 1 2 2 12 7 10 0 9 12 7 12 2
19 1 10 12 9 10 9 15 10 12 13 10 9 15 2 3 1 10 9 2
17 1 14 13 15 13 3 13 2 14 13 14 13 1 12 0 9 2
31 0 13 7 10 9 10 9 15 13 13 0 2 7 13 3 1 12 2 7 0 13 15 15 13 10 9 1 9 7 9 2
21 1 10 15 2 0 13 9 7 10 0 9 13 3 1 9 2 7 13 0 9 2
32 3 2 10 9 13 7 1 9 15 14 13 14 13 1 9 14 13 14 13 7 10 9 10 9 9 3 7 10 9 0 9 2
51 10 9 13 13 1 9 7 2 13 14 13 1 0 9 1 14 13 10 9 14 13 2 7 13 13 7 2 13 14 13 1 9 1 10 9 9 9 1 0 9 2 2 7 13 10 9 10 9 1 9 2
8 13 3 7 0 9 1 15 2
16 10 9 13 7 10 9 9 1 9 13 10 2 0 9 2 2
52 3 2 13 0 14 13 7 2 1 9 10 0 9 10 0 9 10 0 9 3 1 10 9 2 10 0 9 13 1 9 1 10 15 13 10 9 10 9 2 7 13 9 1 9 14 13 10 0 0 9 9 2
17 1 15 13 14 13 10 9 9 1 14 13 10 9 1 0 9 2
24 3 10 9 15 14 13 14 13 2 7 13 14 13 3 0 1 14 13 3 9 1 15 9 2
30 10 9 1 10 9 10 9 13 0 2 1 10 9 9 2 9 0 9 1 10 0 9 7 9 10 9 1 0 9 2
30 7 13 1 9 14 13 14 13 1 13 9 10 9 7 14 13 10 9 10 9 3 1 10 9 1 3 13 9 15 2
26 10 0 9 9 10 9 2 9 2 15 13 13 1 0 9 12 9 2 3 1 3 0 1 10 9 2
1 9
25 3 2 10 9 10 0 9 14 14 13 10 0 9 1 10 9 10 9 1 9 9 1 10 9 2
29 7 13 14 13 10 9 1 9 10 9 1 10 9 7 10 0 9 2 13 0 2 0 7 0 0 9 10 9 2
20 9 13 10 0 9 10 2 2 7 10 9 3 0 9 13 9 1 10 9 2
38 10 9 2 10 9 10 9 13 1 9 2 10 15 13 10 9 15 1 10 9 10 9 15 13 3 2 10 9 15 10 9 13 7 13 0 0 9 2
20 13 10 0 2 0 7 0 9 1 10 3 0 9 15 13 10 9 10 9 2
12 1 10 9 10 9 9 13 9 7 0 9 2
48 13 7 14 13 14 13 3 0 9 7 3 14 13 1 10 0 9 10 9 9 7 3 14 13 10 9 3 0 9 2 3 7 14 13 0 7 10 9 10 15 14 13 14 13 10 0 9 2
3 2 9 2
9 13 3 10 9 10 0 1 9 2
7 15 13 12 3 0 9 2
38 15 9 2 1 15 14 13 13 15 9 10 9 1 12 9 13 13 1 9 10 9 9 2 7 3 3 1 9 0 9 13 10 9 10 12 9 9 2
14 7 13 2 3 14 14 13 9 14 13 10 9 15 2
33 15 13 1 10 0 9 9 2 15 13 2 1 9 2 1 10 0 9 14 13 10 9 1 0 9 9 1 10 9 3 13 3 2
36 10 15 0 9 2 10 9 10 9 2 13 12 9 1 10 15 10 9 13 14 13 2 7 3 13 14 13 7 10 9 14 13 15 10 9 2
40 9 2 13 7 2 12 0 9 13 3 1 9 10 9 15 13 0 1 10 9 12 9 2 1 10 15 13 7 12 9 2 0 9 2 1 9 1 9 2 2
11 1 12 9 13 14 13 12 0 9 9 2
51 14 15 13 3 10 0 9 15 10 9 2 3 13 10 9 10 9 10 9 2 3 1 10 15 10 9 9 13 14 13 10 9 10 9 7 10 9 15 14 13 0 9 3 1 10 9 10 1 9 9 2
62 13 2 3 2 10 9 14 13 1 9 0 9 0 9 7 14 13 0 10 9 10 0 9 1 10 9 7 13 10 9 1 10 9 15 13 1 15 10 9 2 3 7 1 10 0 9 9 2 2 2 10 9 10 0 9 2 1 10 9 10 9 2
29 3 2 13 10 9 10 12 9 2 7 12 3 1 10 9 15 13 1 10 9 1 9 10 12 9 13 1 9 2
27 3 2 10 9 13 10 9 10 9 14 13 10 0 15 9 1 0 15 9 2 1 9 0 10 0 9 2
28 10 0 9 1 9 13 9 9 1 10 9 10 0 9 1 9 10 9 2 10 15 9 13 9 12 0 9 2
60 3 2 3 13 10 9 10 9 1 10 9 7 10 0 9 2 10 9 2 3 13 1 10 0 9 2 14 13 7 13 9 1 10 9 3 10 9 10 9 7 15 13 2 3 13 1 9 10 9 10 9 2 0 9 1 10 0 10 9 2
15 10 9 10 9 2 9 9 2 14 13 10 9 15 2 2
48 3 10 9 13 0 0 7 0 2 7 7 0 0 2 7 10 9 15 13 3 1 9 3 7 1 2 2 3 3 10 0 9 12 9 7 15 15 13 7 13 9 10 9 9 13 3 9 2
17 10 9 13 1 10 0 9 9 10 9 2 1 10 0 9 9 2
11 1 0 9 10 9 13 9 7 0 9 2
34 13 1 10 9 10 0 9 10 9 10 9 2 9 2 10 0 9 9 2 10 9 9 7 10 9 13 1 15 10 9 10 9 9 2
32 14 13 2 7 13 1 15 3 1 9 15 2 1 14 13 15 10 9 1 9 7 14 15 13 3 1 10 9 7 10 9 2
27 13 7 10 9 15 2 13 7 10 0 9 15 15 13 2 14 13 1 0 9 2 7 13 1 10 9 2
40 3 3 13 7 10 9 13 13 3 3 0 2 10 9 1 0 9 13 1 10 9 10 9 10 0 9 2 3 7 1 10 9 10 9 7 10 9 10 9 2
37 10 9 10 9 2 9 9 9 2 13 9 1 9 10 9 1 10 9 9 2 10 15 13 1 9 10 9 9 1 10 0 9 0 9 10 2 2
7 10 9 13 10 0 9 9
7 14 13 10 0 15 9 2
15 13 7 0 3 14 13 14 13 10 0 9 15 3 13 2
52 12 1 15 13 10 9 10 0 9 1 9 2 1 10 15 13 3 9 10 0 9 15 13 1 0 9 7 10 15 9 13 10 9 10 0 0 9 7 10 9 1 10 15 13 15 2 2 13 10 2 9 2
15 9 9 2 13 7 14 15 13 10 9 0 15 10 9 2
28 13 14 13 1 9 7 13 14 13 1 9 15 2 1 9 15 7 1 9 15 7 7 14 13 14 15 13 2
10 3 13 14 13 1 0 7 0 9 2
18 14 13 14 13 0 9 7 14 13 14 13 10 9 9 1 0 9 2
26 3 9 10 9 3 10 12 2 3 7 10 12 0 9 10 9 9 2 13 13 1 15 10 0 9 2
21 1 10 9 10 9 2 10 9 2 10 0 9 13 1 2 3 9 10 13 9 2
43 1 10 3 13 3 13 10 0 9 10 0 9 15 13 10 9 10 0 9 1 9 7 13 1 0 9 3 15 13 1 9 2 10 9 10 12 9 7 10 12 9 2 2
15 10 9 10 9 13 14 13 1 9 10 2 9 1 9 2
13 1 9 10 9 13 1 9 9 1 9 13 9 2
28 10 0 9 13 3 3 13 7 2 1 10 9 2 10 0 9 10 9 14 13 3 1 10 9 15 10 9 2
36 9 9 1 9 13 3 10 9 2 7 10 12 9 10 9 13 3 0 1 10 0 9 7 13 3 10 9 10 0 10 9 10 12 2 12 2
11 9 1 9 1 9 10 9 9 10 2 2
20 7 3 10 9 2 9 7 9 2 3 7 10 0 7 0 9 13 1 9 2
12 3 2 13 10 9 10 9 3 3 1 9 2
28 1 9 10 0 9 2 10 2 13 0 10 9 10 9 1 0 9 7 13 9 1 9 10 9 1 10 9 2
19 0 1 12 9 13 2 7 10 9 9 13 1 9 1 9 10 0 9 2
27 14 15 13 15 9 1 9 10 0 9 10 9 7 10 9 7 3 14 13 14 13 3 1 9 10 9 2
25 10 0 9 10 9 13 10 3 0 9 10 9 1 9 2 7 10 9 1 10 9 15 13 0 2
53 15 9 13 3 1 10 9 10 0 9 10 9 14 13 1 9 3 1 10 9 9 15 9 10 0 10 0 9 2 3 0 9 15 13 1 10 9 10 0 9 2 13 1 9 10 9 10 0 9 1 0 9 2
17 1 0 9 0 9 13 10 9 7 1 0 13 10 0 9 2 2
15 10 0 9 7 10 9 9 10 9 13 3 7 3 0 2
18 3 3 10 12 13 7 10 0 9 13 10 9 10 2 1 9 15 2
19 1 10 9 10 0 9 1 0 9 13 7 10 9 1 0 7 0 9 2
25 10 12 9 1 15 13 13 10 9 10 9 7 10 9 1 9 9 10 2 2 1 9 10 9 2
52 13 14 13 3 10 9 2 3 1 10 9 10 9 2 1 10 9 0 9 7 1 10 0 0 9 10 0 9 2 14 13 7 14 13 3 3 9 1 10 0 7 15 9 7 1 15 9 9 0 9 9 2
13 0 13 10 9 10 0 9 1 9 10 0 9 2
7 10 0 15 13 7 9 2
15 1 10 9 2 13 13 1 10 9 10 9 7 10 9 2
17 1 9 13 2 3 2 9 1 9 10 9 10 9 1 0 9 2
57 10 9 10 9 1 10 9 9 13 0 9 1 10 9 1 9 7 13 10 0 0 9 7 10 9 14 13 3 15 1 0 9 10 0 9 10 9 1 9 10 0 9 7 14 13 14 15 13 1 9 1 10 9 15 10 9 2
23 3 10 9 12 9 13 3 1 0 9 2 1 9 10 9 12 9 7 10 9 3 12 2
26 10 12 10 9 13 0 10 9 1 10 9 2 10 15 13 1 10 9 10 0 9 1 10 0 9 2
28 10 9 13 1 12 9 1 9 7 1 9 10 0 13 1 9 2 9 10 9 7 3 10 0 9 10 9 2
31 15 10 9 13 9 2 1 10 9 2 10 9 2 9 2 10 9 2 0 9 2 10 15 14 13 3 1 10 0 9 2
6 10 9 9 3 13 2
42 13 7 10 9 10 0 9 7 9 14 14 13 7 10 0 9 10 9 14 13 1 0 9 7 13 14 13 7 10 0 9 10 9 15 3 3 1 3 13 13 9 2
19 1 0 15 10 9 15 13 13 9 14 13 13 3 0 9 1 10 9 2
26 3 1 10 9 2 13 0 14 13 14 13 0 1 12 10 0 9 2 7 15 13 0 1 13 9 2
25 1 9 15 2 10 9 13 14 13 9 7 9 2 7 10 3 9 13 0 1 0 9 1 9 2
35 3 13 10 9 2 1 15 13 14 13 7 14 13 1 15 15 14 14 13 14 13 2 7 13 14 15 13 7 13 14 15 13 1 9 2
10 9 9 10 9 1 10 9 10 9 2
46 7 10 0 9 13 14 13 1 10 0 9 2 13 9 1 9 10 9 9 7 0 9 2 1 9 10 9 9 1 10 0 9 2 1 9 1 10 9 10 0 9 1 10 0 9 2
8 0 0 9 1 9 7 9 2
1 9
19 9 10 9 13 14 13 2 1 10 12 2 10 3 0 9 1 9 2 2
13 1 14 13 9 2 13 14 13 9 2 3 9 2
12 3 15 13 10 9 15 13 1 9 10 9 2
33 13 3 0 14 13 15 3 2 0 9 7 14 13 10 0 9 1 10 9 15 10 9 10 15 13 3 10 9 3 7 10 9 2
12 14 13 7 0 2 10 9 15 14 13 0 2
27 13 1 9 0 10 9 7 10 0 9 14 13 7 0 10 9 7 0 10 9 14 13 0 7 0 9 2
10 1 10 9 10 9 13 9 10 9 2
24 13 3 7 10 9 14 13 14 13 10 9 9 9 1 9 9 10 15 13 3 10 0 9 2
23 10 9 9 13 1 10 9 9 1 9 12 2 1 9 10 9 10 12 10 9 9 12 2
15 10 9 13 7 2 14 13 1 12 10 9 10 9 2 2
31 1 12 9 10 9 13 3 10 9 10 9 7 12 9 1 10 9 10 0 9 2 10 9 9 13 10 0 9 10 9 2
26 2 13 10 9 9 14 13 10 9 15 1 10 9 10 9 10 9 0 9 2 13 10 9 7 13 2
47 13 3 3 3 1 10 9 15 13 1 10 9 10 9 9 7 0 9 2 3 13 3 2 3 13 10 0 9 2 7 3 14 13 14 13 3 3 10 0 3 7 10 0 7 0 9 2
24 1 10 9 10 9 13 0 9 7 9 1 15 13 3 1 14 13 1 10 9 7 10 9 2
26 10 9 13 7 0 9 13 10 9 9 12 9 9 9 10 9 7 7 13 13 0 9 1 9 15 2
29 2 12 9 2 9 10 9 9 7 10 9 9 2 13 1 12 1 10 9 2 7 13 10 9 7 10 0 9 2
11 3 1 9 10 9 13 10 9 14 13 2
17 10 9 10 9 13 10 0 9 1 12 9 9 2 10 0 9 2
18 3 9 15 10 9 10 9 13 2 3 2 10 0 9 7 10 9 2
37 1 12 10 9 2 1 10 0 9 13 10 9 1 9 10 9 2 14 7 1 10 9 10 9 2 15 13 10 9 15 7 13 10 9 10 9 2
15 3 2 10 9 10 0 9 10 2 13 1 12 9 9 2
24 10 9 13 7 13 1 10 0 9 10 9 9 10 2 1 10 9 2 7 14 15 13 0 2
22 10 9 9 13 7 2 10 9 9 13 1 9 1 10 9 10 9 2 9 9 2 2
22 3 1 9 15 13 13 1 9 9 2 10 9 13 3 14 13 1 10 9 10 9 2
32 10 0 9 2 15 13 10 9 2 13 0 9 1 10 9 10 9 15 7 13 1 0 9 1 10 9 7 13 9 0 9 2
11 13 3 3 1 9 10 9 9 10 12 2
36 10 0 9 1 9 14 13 3 13 1 9 10 0 9 7 10 9 13 13 10 9 10 9 7 15 13 1 10 9 15 13 1 0 0 9 2
17 13 7 10 9 9 14 13 3 1 10 0 9 15 1 10 9 2
36 10 9 10 9 13 0 1 10 9 2 7 7 13 1 0 9 10 9 10 9 2 10 0 9 9 1 10 9 7 9 10 9 10 3 9 2
22 10 9 13 1 10 0 9 9 10 9 7 10 9 10 2 14 13 1 9 10 9 2
9 13 14 13 3 1 9 10 9 2
13 10 9 2 10 0 0 9 10 9 13 1 9 2
21 13 15 3 14 13 15 9 1 9 10 9 9 7 10 9 15 13 1 9 9 2
25 10 0 9 13 9 1 0 9 1 12 9 15 13 3 1 0 0 9 1 9 1 10 0 9 2
58 13 14 13 14 13 7 10 0 9 14 13 14 13 10 9 7 3 13 10 0 9 0 9 9 2 10 9 1 10 9 9 7 9 2 10 0 9 15 14 15 13 2 3 7 15 10 9 1 10 9 9 7 10 9 15 13 3 2
10 10 9 13 10 9 0 9 1 9 12
13 10 9 13 9 3 10 9 10 9 7 12 9 2
4 13 12 9 2
4 2 0 9 2
50 10 9 10 9 10 9 1 9 13 10 12 9 10 0 0 2 10 2 12 9 2 1 10 0 0 2 7 13 1 12 9 2 2 12 9 2 2 2 15 13 10 12 1 10 2 0 2 9 10 2
32 14 13 1 10 15 2 1 15 7 13 15 1 10 0 9 15 10 9 2 14 13 1 9 10 0 15 9 1 15 10 9 2
35 10 9 13 1 9 10 9 1 12 9 12 7 10 9 13 7 2 13 0 7 13 14 13 10 9 10 0 9 3 1 10 9 9 2 2
35 10 9 13 1 10 9 1 9 1 0 9 7 1 9 2 1 0 9 9 13 3 10 2 9 2 7 13 14 13 1 9 1 3 9 2
33 1 0 9 2 10 0 9 10 9 13 9 7 9 2 10 15 13 10 9 15 1 10 9 10 9 15 13 10 9 1 10 9 2
19 1 14 13 0 9 2 13 14 13 1 9 10 9 10 9 15 13 3 2
9 10 9 13 10 9 10 9 9 2
11 14 13 10 9 10 9 15 13 3 3 2
32 1 9 2 10 9 13 9 1 9 10 0 9 2 13 7 10 0 0 9 10 0 9 14 13 10 9 10 9 1 10 9 2
11 10 9 10 9 13 14 13 10 0 9 2
8 10 9 13 1 9 1 9 2
36 9 13 7 2 10 9 13 9 1 12 9 10 9 9 10 9 10 2 0 9 2 7 9 10 9 1 9 15 13 10 12 9 10 9 2 2
21 7 10 12 9 13 10 0 9 7 10 9 10 9 2 10 9 1 9 3 2 2
11 13 0 10 9 7 13 3 7 3 3 2
13 13 12 2 3 10 9 10 9 7 13 9 12 2
35 13 3 7 10 9 10 9 1 10 9 2 10 9 1 10 9 2 10 0 9 2 15 9 10 0 9 2 12 9 7 10 9 10 9 2
20 10 0 15 9 13 1 9 10 0 9 9 7 10 9 9 7 9 10 2 2
14 10 9 13 0 1 15 9 13 3 1 10 0 9 2
15 10 9 1 9 15 13 7 0 9 9 14 13 10 9 2
7 14 13 3 10 9 15 2
21 3 13 10 0 9 7 1 13 14 13 7 10 0 9 13 0 1 10 0 9 2
22 10 2 7 10 0 9 15 13 14 13 10 9 15 1 10 9 1 10 9 10 12 2
25 10 9 13 10 9 10 9 2 1 9 9 7 9 9 10 0 9 13 1 9 1 10 9 15 2
21 13 10 9 9 1 10 9 7 3 10 9 2 12 1 10 15 13 13 1 9 2
18 13 1 10 0 9 2 7 13 3 10 9 1 14 13 10 9 3 2
1 9
17 10 0 0 9 13 13 3 1 0 9 7 1 9 10 0 9 2
14 1 15 7 13 7 3 13 10 0 9 14 13 2 2
15 10 9 2 10 9 13 0 9 7 13 1 10 0 9 2
1 9
18 3 2 15 9 13 7 7 13 1 9 13 15 0 15 13 3 3 2
20 10 0 9 7 10 9 10 2 2 9 9 2 13 13 7 14 13 10 9 2
46 3 13 10 0 9 10 0 9 13 7 2 3 1 10 9 14 13 10 9 1 0 9 7 14 13 0 9 1 0 9 2 10 0 9 2 7 10 9 3 2 13 10 9 10 9 2
32 3 10 2 14 13 14 13 10 9 12 2 10 15 1 9 13 0 9 9 10 9 1 9 9 2 13 10 0 9 10 9 2
23 10 9 13 13 3 9 1 10 9 9 9 10 9 1 9 7 10 9 15 1 0 9 2
22 1 9 10 0 9 14 13 1 9 14 13 3 2 3 14 13 3 10 0 9 15 2
13 13 7 15 10 0 9 14 13 1 9 10 0 2
6 13 10 9 3 9 2
11 10 9 15 13 1 10 14 13 9 9 2
22 1 0 9 9 10 0 9 13 1 10 9 2 7 10 9 13 1 2 12 9 9 2
76 3 13 10 9 10 0 9 2 10 0 9 13 10 9 15 13 1 15 10 9 10 9 1 10 9 2 1 9 2 1 10 0 9 2 10 9 0 9 2 15 13 3 1 10 9 2 1 2 2 12 2 1 14 13 0 9 1 10 0 9 2 10 15 13 13 10 9 15 14 13 3 1 15 10 9 2
21 3 9 10 0 9 13 14 13 10 9 1 10 0 0 9 1 10 9 10 9 2
32 3 13 10 9 9 2 0 10 9 10 0 9 1 10 9 2 2 10 0 9 9 15 13 9 13 10 9 10 0 9 2 2
20 15 9 14 13 14 13 7 1 0 9 7 9 7 1 0 9 1 10 2 2
21 1 9 13 10 9 7 14 10 9 10 9 2 10 15 7 13 1 9 1 9 2
12 0 15 13 10 9 15 3 9 10 0 9 2
29 14 13 14 15 13 10 9 1 14 13 7 10 0 9 14 13 10 9 10 0 9 10 0 2 7 10 9 9 2
11 13 10 0 9 1 10 9 10 0 9 2
53 10 0 9 13 3 7 10 9 15 13 13 1 0 1 12 9 10 2 1 9 9 1 10 9 7 13 1 10 2 14 13 3 1 9 15 13 10 2 9 9 7 9 15 1 2 2 2 3 13 10 2 9 2
15 1 9 10 12 0 9 7 10 0 9 13 10 9 15 2
19 10 9 10 9 13 10 9 15 1 9 10 3 9 10 9 2 9 9 2
21 3 2 3 1 9 13 10 0 9 1 9 2 7 10 9 13 3 1 10 9 2
20 13 10 9 15 13 10 0 0 9 7 13 3 0 13 10 9 10 0 9 2
19 15 13 1 10 9 15 10 9 2 7 14 13 10 9 1 15 10 9 2
10 0 9 1 9 0 1 9 10 9 2
27 1 15 10 9 13 10 0 9 9 2 1 10 0 10 9 7 10 9 14 13 2 13 14 13 0 9 2
41 3 1 0 9 2 10 13 9 2 10 0 9 1 9 9 7 10 12 9 2 10 9 15 14 13 10 0 9 2 10 0 0 10 9 15 13 1 9 10 9 2
33 10 0 9 10 9 10 9 1 2 7 10 0 9 1 10 9 13 9 10 9 15 3 7 3 2 12 9 3 2 13 1 0 2
64 7 13 10 9 0 9 10 9 2 13 3 1 9 3 10 9 1 10 9 7 9 10 9 2 10 9 1 10 0 9 9 2 7 3 10 9 9 1 10 9 0 9 2 1 9 10 0 2 7 1 10 9 15 0 2 9 10 9 1 0 9 15 9 2
7 12 9 13 1 9 10 9
19 10 0 9 13 3 2 13 3 2 10 0 9 2 13 10 0 9 9 2
12 10 0 9 10 9 13 1 9 1 0 9 2
39 3 7 1 10 9 10 0 9 1 9 2 0 0 9 1 0 9 13 1 0 9 7 13 0 9 2 7 3 13 3 1 0 0 9 10 0 9 2 2
27 1 0 9 13 7 10 9 9 2 1 10 15 13 0 9 15 13 0 10 9 1 10 9 3 12 9 2
27 10 9 1 9 7 10 9 10 0 7 0 9 13 10 9 1 9 14 13 15 9 1 10 9 10 9 2
62 14 13 14 13 1 9 10 9 10 9 1 10 9 15 10 9 2 3 3 3 13 2 13 1 9 1 10 9 1 10 9 10 0 9 15 15 13 1 0 15 9 2 1 14 13 3 1 10 9 15 13 3 3 2 3 1 15 15 13 3 3 2
14 3 2 10 9 1 9 9 9 13 1 9 7 9 2
23 7 13 14 13 1 9 10 0 9 15 13 2 3 10 9 13 14 13 10 9 9 9 2
20 13 14 13 14 13 10 0 15 9 2 7 0 9 3 14 13 14 15 13 2
35 10 0 9 2 10 0 9 7 10 9 13 7 10 9 2 9 12 2 14 13 1 10 9 1 9 9 1 9 10 0 9 10 0 9 2
29 3 2 10 9 9 13 9 1 9 7 1 0 9 2 10 15 7 7 14 13 1 0 9 13 9 1 0 9 2
20 10 9 10 9 9 13 10 3 9 10 0 0 9 2 9 12 2 14 13 2
15 3 3 3 14 13 10 0 9 13 14 15 13 9 9 2
43 10 0 9 15 14 13 10 9 0 10 9 7 10 0 9 15 2 1 15 7 15 13 1 9 2 7 3 13 0 10 0 9 15 7 13 0 10 9 9 15 1 9 2
29 1 0 9 13 1 10 0 9 10 9 10 9 1 9 10 9 10 9 9 2 9 9 2 1 10 0 1 9 2
25 10 9 13 10 9 1 9 14 13 10 9 7 14 15 13 1 9 2 2 13 9 10 0 9 2
29 1 0 9 2 9 9 2 3 13 7 10 0 9 10 9 13 1 10 9 10 9 2 1 10 9 9 7 9 2
24 15 10 9 13 10 3 0 1 3 3 10 9 13 9 1 9 1 10 9 10 12 9 12 2
10 7 3 14 13 0 9 10 0 9 2
16 15 9 1 15 13 10 3 0 9 1 10 2 9 7 9 2
16 10 9 10 9 2 10 9 7 10 9 13 1 3 13 9 2
28 1 10 12 0 9 2 10 0 9 13 1 10 0 9 2 1 10 0 9 3 2 0 9 2 3 1 9 2
20 1 10 0 9 13 0 0 9 2 3 10 0 9 1 10 9 15 3 13 2
18 10 9 15 13 0 7 10 9 1 0 9 13 1 9 10 0 9 2
30 14 13 3 1 10 9 2 12 15 13 10 9 10 9 15 10 9 7 14 13 10 0 9 15 13 14 13 3 0 2
1 9
37 10 9 13 3 0 9 1 14 13 10 9 0 9 9 9 9 14 13 10 9 15 1 10 9 7 14 13 14 13 9 10 0 9 1 10 3 2
52 15 13 13 3 0 9 1 0 9 2 7 0 1 15 10 9 13 1 12 0 9 15 2 1 10 15 15 13 2 14 14 13 3 0 1 10 0 0 9 15 13 10 9 2 7 14 13 3 0 0 9 2
13 3 2 10 9 13 10 0 7 0 9 10 9 2
25 3 14 13 1 12 3 9 7 3 1 9 1 10 9 10 9 10 9 1 10 9 10 9 9 2
18 10 9 10 9 13 1 10 13 9 2 10 3 9 14 13 3 9 2
1 9
5 9 9 13 10 9
12 3 1 10 9 13 0 9 1 10 0 9 2
17 10 9 10 9 13 3 10 9 15 13 1 3 7 13 0 9 2
8 13 0 9 2 9 7 9 2
18 15 10 9 13 0 9 1 10 3 9 2 10 9 7 10 0 9 2
18 10 9 10 9 13 2 3 1 3 2 1 9 15 7 1 9 15 2
33 3 1 9 1 0 9 10 9 2 13 7 3 14 13 14 13 0 1 10 12 15 15 13 9 10 9 2 3 0 9 0 9 2
1 9
52 7 7 10 9 13 10 0 9 15 13 1 9 2 13 10 9 15 2 14 13 7 10 9 2 1 14 14 13 1 0 9 10 9 2 14 13 1 0 9 10 9 2 13 10 9 1 0 9 1 0 9 2
8 10 2 13 10 9 1 9 2
40 10 12 0 9 10 9 7 9 9 10 9 9 9 7 10 0 9 9 9 2 10 9 2 13 10 9 1 0 9 7 9 2 15 3 13 10 9 10 9 2
37 10 0 9 9 2 1 10 15 13 3 1 9 7 9 10 15 14 13 14 13 7 3 1 9 2 14 13 7 14 13 1 10 0 9 10 9 2
4 2 2 1 2
27 10 9 13 0 9 2 13 7 1 9 9 7 13 1 9 1 10 9 10 0 9 2 3 13 13 9 2
18 10 9 15 3 13 1 9 10 9 13 10 9 10 9 10 0 9 2
26 10 9 12 13 10 0 0 9 7 13 1 9 15 13 1 10 15 9 3 9 1 0 9 12 9 2
13 3 2 10 9 15 13 1 14 13 3 15 9 2
15 1 15 13 14 13 2 15 13 10 9 7 10 9 15 2
29 15 13 12 1 10 9 1 10 15 13 14 13 0 0 9 2 1 14 13 1 0 9 10 9 1 10 0 9 2
26 3 10 9 10 9 13 3 1 15 14 13 3 1 9 7 7 10 9 15 13 0 14 13 3 3 2
8 10 12 9 13 10 0 9 2
17 10 0 9 3 1 10 3 0 1 9 2 13 9 1 10 9 2
19 10 0 9 1 10 9 7 10 0 0 9 9 13 1 0 9 10 9 2
15 1 0 0 9 13 7 10 9 2 10 9 7 10 9 2
12 13 1 10 9 10 0 9 1 15 10 9 2
15 3 1 12 9 2 10 9 13 10 0 12 1 10 9 2
27 10 9 7 9 13 1 9 10 9 2 1 9 12 9 1 10 9 9 7 13 9 10 9 1 10 9 2
20 10 9 13 10 12 0 9 3 13 1 12 9 10 0 9 1 10 9 9 2
9 10 9 14 13 10 9 1 9 2
23 10 0 9 13 1 9 10 9 1 0 9 2 10 15 10 9 9 13 2 0 9 2 2
64 10 9 15 2 15 3 13 13 2 3 13 14 13 1 0 0 9 7 2 1 15 10 9 2 13 3 10 9 10 2 9 2 10 15 13 7 10 0 9 13 14 13 0 9 1 14 13 14 13 15 10 9 2 7 14 13 10 9 10 9 7 10 9 2
21 3 3 2 7 10 9 13 14 13 3 0 2 14 13 3 14 13 15 10 9 2
46 3 13 10 9 15 10 9 2 7 14 14 13 14 13 3 7 10 9 13 10 9 14 13 1 3 0 9 7 1 0 9 2 7 3 13 14 13 1 9 15 1 10 0 0 9 2
17 9 15 13 14 13 10 9 9 14 13 10 9 3 9 9 15 2
33 10 9 13 3 7 10 0 9 14 13 14 13 13 14 13 1 0 9 10 9 1 10 15 13 14 13 9 1 10 0 0 9 2
9 0 9 1 10 9 12 10 9 2
29 9 9 2 9 9 2 3 13 3 10 9 15 13 2 10 9 1 9 13 3 7 3 0 1 10 9 10 9 2
9 13 0 7 13 1 10 9 9 2
32 7 15 13 2 3 10 9 13 2 3 2 1 9 7 10 9 9 13 2 3 3 2 9 0 9 1 10 9 7 10 9 2
8 13 10 0 9 2 2 9 2
28 3 10 9 9 13 9 1 10 9 10 9 9 7 2 10 9 14 13 14 13 14 13 3 1 15 9 2 2
16 3 2 13 10 9 1 0 9 9 1 0 9 7 0 9 2
37 7 3 15 13 0 2 7 13 7 15 13 9 2 3 7 14 13 14 13 1 0 10 9 2 13 0 9 7 14 14 13 10 9 1 0 9 2
48 1 10 9 15 1 9 10 9 2 10 9 9 13 3 1 10 9 9 2 13 0 1 12 9 2 7 13 10 0 9 2 10 9 2 1 10 9 15 13 3 1 9 1 7 12 9 9 2
36 10 9 10 12 9 10 9 7 9 9 7 10 9 9 10 9 15 10 0 9 1 15 10 9 13 10 9 10 9 14 13 1 10 0 9 2
14 7 2 10 9 9 1 9 13 10 9 1 10 9 2
2 12 2
37 1 10 9 10 9 10 9 13 0 9 2 1 9 3 12 2 10 9 15 1 9 2 10 9 2 10 9 2 10 9 2 10 9 7 10 9 2
31 3 2 14 13 3 13 7 13 14 13 0 9 10 0 9 1 0 0 9 7 13 7 15 15 14 13 10 9 1 9 2
23 10 9 13 7 13 0 14 13 10 9 7 10 9 13 3 9 3 1 10 9 10 9 2
37 10 0 0 9 13 10 2 7 10 0 10 9 2 10 2 15 13 13 1 9 10 2 7 1 0 15 9 13 1 9 15 1 9 14 0 9 2
23 10 9 9 15 13 3 1 9 10 9 13 10 0 9 9 7 9 10 0 9 1 9 2
64 13 10 0 9 9 1 9 7 9 2 1 0 9 9 1 9 9 10 0 9 2 7 3 10 9 10 9 10 9 13 13 10 13 9 1 10 9 10 9 15 2 15 13 14 13 1 10 9 15 1 10 0 9 7 10 0 0 9 15 13 1 0 9 2
20 13 0 10 9 10 9 2 7 13 0 10 9 15 0 1 10 9 0 9 2
56 13 14 15 13 7 10 0 9 14 13 3 14 13 10 9 7 2 3 13 10 0 9 7 10 0 9 2 13 14 13 7 13 0 0 9 7 0 9 1 9 3 13 14 13 10 9 2 10 9 7 10 0 9 10 9 2
46 0 9 7 0 9 0 0 9 13 10 0 9 1 9 9 2 9 1 9 2 9 2 9 7 9 7 3 15 0 9 7 9 2 3 10 2 9 2 7 3 2 9 10 9 2 2
24 10 9 13 14 13 1 10 9 7 10 9 10 9 9 2 14 15 13 3 10 9 15 9 2
34 10 3 13 7 1 10 9 7 13 13 1 10 0 9 2 10 9 13 0 2 13 9 7 2 1 10 9 10 12 9 13 9 2 2
17 1 15 10 9 13 1 3 12 9 10 9 7 10 9 15 13 2
33 9 9 9 9 10 9 2 9 9 2 13 10 9 15 9 7 13 1 10 9 10 9 10 9 10 9 2 9 0 10 9 2 2
5 1 9 10 9 2
38 14 13 7 2 3 13 2 7 10 9 10 0 9 7 10 0 9 1 9 15 13 14 13 10 2 9 9 3 13 10 9 9 13 14 13 1 9 2
19 10 0 9 2 15 13 1 10 9 9 10 9 2 13 0 3 0 9 2
2 12 2
30 13 7 14 13 1 9 2 10 9 7 10 9 15 13 3 15 14 14 13 9 10 0 9 1 9 10 9 10 9 2
6 14 13 1 9 15 2
21 1 15 10 9 2 13 14 13 10 9 1 10 0 2 10 0 7 10 0 9 2
11 10 9 9 13 1 10 9 9 1 9 12
18 13 10 0 1 10 0 9 14 13 9 3 2 1 0 9 7 3 2
10 10 0 9 14 13 3 14 13 9 2
15 10 9 9 10 2 2 9 9 2 13 10 9 0 9 2
37 7 10 0 10 0 9 9 2 9 9 2 13 7 10 9 10 0 9 15 13 1 3 10 9 13 13 1 0 9 9 1 10 9 0 0 9 2
31 10 9 2 10 0 9 10 9 2 3 12 0 9 1 10 9 13 1 10 0 9 15 2 10 0 9 7 10 0 9 2
32 1 10 9 9 9 10 0 9 13 7 2 10 9 9 13 1 9 10 0 0 9 2 10 15 13 10 9 9 1 12 9 2
19 3 13 2 2 10 2 14 13 0 10 0 9 1 14 13 10 9 2 2
15 14 13 0 2 10 0 15 9 0 9 13 1 10 9 2
14 14 13 2 7 2 10 9 9 12 9 10 9 2 2
8 10 9 13 1 12 0 9 2
52 13 7 2 3 1 15 2 13 14 13 10 9 10 9 1 10 9 9 7 2 3 2 14 13 0 9 0 10 9 1 9 0 10 12 9 7 14 14 13 10 9 1 3 0 9 9 3 1 9 0 9 2
19 13 0 10 9 10 0 9 7 13 10 0 9 2 3 13 10 9 9 2
27 1 0 9 13 1 12 9 15 10 9 10 9 2 1 9 2 1 10 9 7 10 9 2 10 0 9 2
47 14 13 14 13 0 1 10 0 9 15 13 13 1 10 9 15 10 9 2 3 1 9 10 9 15 13 3 3 1 10 9 9 1 10 0 9 2 10 15 14 13 0 9 1 10 9 2
21 1 10 9 2 10 9 13 10 9 15 2 15 13 1 15 2 7 13 10 9 2
54 1 10 0 9 2 13 14 13 15 9 3 13 15 10 9 2 3 1 10 9 10 9 9 1 10 9 1 10 9 2 10 9 9 1 10 9 10 0 9 2 10 9 10 0 9 1 12 12 10 0 9 10 2 2
9 9 9 13 1 15 7 10 9 2
15 14 13 2 7 2 10 9 15 1 9 15 2 2 9 2
26 7 3 10 9 1 10 0 9 13 1 0 9 2 13 1 9 10 9 10 9 1 9 0 9 1 2
9 10 0 9 10 2 13 1 9 2
42 7 0 9 13 10 9 10 9 2 10 9 2 15 13 9 1 9 1 10 0 9 15 2 13 1 10 9 15 1 10 9 15 13 14 13 3 1 10 9 10 9 2
18 10 2 13 14 13 10 9 1 10 1 9 9 9 7 9 1 9 2
14 10 0 9 13 1 9 1 10 0 9 1 10 9 2
37 10 0 9 10 0 9 10 15 13 10 9 13 2 13 2 0 2 7 10 9 13 7 14 13 14 13 3 10 9 9 10 9 2 3 9 9 2
20 14 13 2 9 2 1 15 10 9 14 13 15 15 13 1 9 10 9 15 2
8 13 10 9 10 0 9 9 12
15 1 0 9 10 9 13 10 9 10 9 2 9 9 2 2
44 10 0 9 15 14 13 14 13 0 10 0 9 10 0 9 7 10 0 9 2 1 10 9 10 0 9 1 9 0 10 9 1 0 9 2 1 9 0 9 1 9 13 9 2
10 10 9 13 0 10 0 9 10 9 2
16 3 13 14 13 10 9 15 9 9 7 10 9 15 1 9 2
44 13 7 3 1 10 0 9 7 10 3 0 9 1 9 0 9 7 0 9 13 3 9 14 13 3 10 12 9 1 10 9 1 9 2 15 13 7 14 13 0 10 9 15 2
27 3 13 7 13 10 0 9 9 1 10 9 10 0 9 2 13 10 9 2 13 14 13 10 9 10 2 2
10 10 9 10 9 13 10 9 10 9 9
13 3 13 7 13 9 1 14 13 10 9 10 9 2
32 10 9 13 0 2 3 1 15 10 9 3 7 1 15 0 9 2 7 14 13 1 9 3 1 0 9 7 0 9 15 13 2
10 10 9 13 13 10 9 9 10 9 2
9 9 2 0 9 1 9 9 9 2
13 10 0 9 9 7 9 13 10 0 9 10 9 2
21 3 10 9 9 15 13 10 9 14 13 3 10 9 9 1 7 1 10 0 9 2
36 0 9 10 9 10 9 13 1 9 10 9 2 9 1 9 2 2 10 15 10 0 9 13 9 1 10 9 10 9 10 9 1 0 10 9 2
11 10 9 7 9 13 10 9 10 0 9 2
19 3 2 14 13 1 9 9 2 9 7 9 1 10 9 10 9 3 9 2
11 10 9 10 9 13 7 10 9 7 9 2
22 1 0 9 13 3 14 13 10 9 15 1 14 13 10 9 2 3 1 10 0 9 2
40 10 9 10 9 2 1 10 12 9 2 12 1 15 9 10 9 2 7 10 12 9 2 13 1 9 10 0 9 7 13 3 1 9 2 10 9 7 10 9 2
29 15 13 10 3 0 13 9 10 9 9 2 7 10 0 9 13 12 2 7 1 9 12 1 12 9 13 12 9 2
13 15 13 7 10 9 13 10 9 15 1 12 9 2
28 15 13 15 15 2 13 2 14 13 3 7 3 10 9 15 2 7 14 13 3 7 0 9 14 13 0 9 2
11 13 3 1 10 0 9 3 13 10 9 2
6 7 10 9 14 13 2
11 15 13 3 10 0 9 2 15 15 13 2
23 3 2 13 14 13 7 15 12 9 15 10 15 13 3 10 9 1 10 2 0 9 9 2
25 13 3 3 0 14 13 7 2 1 10 9 2 10 9 15 14 13 14 13 1 9 10 0 9 2
26 13 1 9 10 9 10 9 9 9 9 13 7 2 10 9 13 1 9 1 10 9 15 13 3 2 2
8 1 0 9 13 7 14 13 2
23 3 0 10 9 3 1 9 10 9 13 10 9 10 9 10 2 2 10 15 13 1 9 2
28 10 0 1 10 9 15 13 13 1 3 13 3 3 1 9 9 7 1 10 0 7 0 9 15 13 14 13 2
37 10 9 15 1 9 9 1 0 9 13 12 9 2 3 12 9 9 1 10 15 13 0 9 2 7 13 1 0 10 0 9 10 9 10 0 9 2
25 13 7 10 0 9 10 9 13 1 9 2 1 9 10 9 15 10 9 13 2 9 7 9 2 2
10 3 2 13 14 13 1 9 10 9 2
1 9
15 7 13 3 1 10 9 15 10 9 15 2 14 13 9 2
14 13 13 3 3 1 12 9 1 15 13 10 0 9 2
42 13 10 0 9 1 10 9 15 10 9 2 1 10 9 15 13 0 9 2 7 13 14 13 10 9 15 1 9 7 1 9 7 10 9 15 1 10 9 15 10 9 2
31 1 15 10 9 2 9 9 10 9 2 15 13 10 9 1 9 10 0 9 3 1 10 9 0 9 2 15 13 3 0 2
40 3 1 10 9 13 0 7 10 9 1 10 9 1 9 13 1 12 2 7 0 9 13 7 10 9 2 1 10 12 2 13 12 9 2 13 13 12 9 9 2
27 10 9 9 13 9 10 9 10 9 2 7 13 10 9 1 3 15 13 3 1 9 15 9 9 10 9 2
62 13 1 9 7 14 13 10 0 9 7 1 10 9 7 1 10 0 9 2 7 3 10 9 1 10 0 9 9 10 15 2 3 15 2 13 14 13 10 9 7 13 14 15 13 3 2 1 10 9 10 9 2 10 15 13 0 1 12 3 9 3 2
55 14 13 3 10 3 0 9 1 10 9 15 2 7 14 13 14 13 10 9 7 10 9 15 0 9 2 3 13 7 15 2 14 13 10 9 15 13 10 9 1 10 9 7 14 13 14 13 10 9 1 10 0 15 9 2
36 10 0 9 13 12 9 15 13 9 9 3 1 0 9 1 9 2 10 15 13 9 15 13 9 14 13 1 14 13 1 9 1 10 9 9 2
17 10 9 2 9 10 0 9 2 13 13 3 1 9 10 9 9 2
11 1 9 10 9 13 1 0 9 12 9 2
13 3 10 0 9 13 14 13 9 1 10 0 9 2
31 10 9 10 0 9 1 9 13 7 2 3 13 9 10 9 10 12 2 3 13 10 9 15 13 9 1 9 1 3 2 2
20 1 10 2 2 12 9 13 10 9 15 2 10 12 1 9 2 7 12 13 2
22 13 0 7 13 9 2 3 2 10 9 10 9 9 13 1 9 10 0 9 7 9 2
4 0 0 9 2
