29146 17
12 9 9 15 9 13 2 15 15 13 9 0 2
20 13 16 15 7 13 2 15 9 13 2 3 3 0 2 13 13 15 13 9 2
8 1 15 13 1 15 9 9 2
3 13 9 2
5 3 13 3 13 2
7 7 3 13 13 0 9 2
14 15 1 15 13 13 9 9 2 15 13 9 0 13 2
16 9 16 13 0 9 2 0 9 9 13 9 7 13 0 9 2
9 3 13 9 9 9 9 13 9 2
30 16 0 9 13 0 2 2 3 16 0 15 2 7 16 0 3 13 2 2 9 7 13 13 2 9 0 3 9 13 2
17 9 13 0 9 9 0 9 13 1 9 2 15 13 9 9 13 2
20 9 9 13 7 15 13 0 9 2 13 15 3 9 9 9 7 13 0 9 2
20 15 13 9 16 13 3 2 3 12 3 13 1 9 9 7 13 9 0 13 2
12 15 9 13 3 13 9 7 1 9 0 13 2
20 15 16 13 0 9 2 0 13 9 13 1 9 2 0 16 13 15 13 13 2
12 3 13 15 9 2 15 9 0 13 13 12 2
9 3 9 13 0 2 9 13 9 2
12 3 7 13 9 13 1 9 2 13 16 13 2
18 16 13 13 0 9 15 7 3 9 9 13 2 9 15 15 9 13 2
14 13 0 9 9 2 9 9 15 13 13 15 7 13 2
9 3 13 15 15 13 9 0 9 2
9 15 0 9 13 9 13 7 9 2
10 3 13 9 13 13 13 1 0 9 2
7 1 15 13 0 13 9 2
24 13 15 16 13 9 7 15 9 13 13 13 2 7 15 13 13 9 7 15 9 15 13 9 2
7 13 3 0 15 0 13 2
25 9 1 9 9 16 13 13 2 9 1 9 13 9 15 2 0 7 9 1 0 13 13 13 13 2
17 3 13 9 7 15 13 9 13 9 2 7 15 13 13 3 13 2
7 3 13 0 1 0 9 2
6 13 15 9 9 15 2
14 9 7 9 7 13 9 9 0 13 1 9 1 9 2
16 15 16 13 9 0 9 2 3 13 13 2 9 13 2 9 2
9 12 2 16 13 0 2 13 15 2
10 3 2 16 3 13 2 15 13 12 2
7 0 13 16 15 12 13 2
7 3 0 9 0 9 13 2
11 0 9 0 13 9 9 7 3 13 13 2
13 9 3 9 16 13 13 2 9 9 13 1 9 2
7 9 13 13 9 9 9 2
8 15 13 13 2 16 13 9 2
6 9 0 3 9 13 2
16 15 15 13 13 2 15 9 7 9 9 13 2 9 0 13 2
10 15 9 9 1 0 13 2 12 13 2
20 9 13 9 16 13 9 2 0 9 13 13 12 13 9 2 16 15 13 0 2
18 3 13 13 9 13 9 2 9 7 13 9 9 2 0 13 9 9 2
13 15 3 13 7 0 9 13 0 13 0 13 9 2
12 13 1 9 2 9 13 0 2 9 13 9 2
5 15 3 13 9 2
13 16 13 2 15 9 0 13 9 7 0 13 13 2
13 15 3 0 15 13 0 2 0 9 9 13 15 2
14 15 0 9 12 13 2 7 16 0 13 2 13 9 2
6 15 13 0 9 9 2
6 9 13 9 9 9 2
7 3 9 1 15 13 9 2
11 15 9 16 13 15 2 13 13 9 9 2
7 15 3 13 13 15 13 2
14 9 0 2 9 13 9 2 0 13 2 13 13 9 2
24 13 9 9 16 13 9 2 13 15 9 7 13 3 2 16 0 9 13 0 2 13 15 13 2
13 3 9 9 3 0 13 9 0 7 13 9 9 2
12 15 16 13 9 13 13 2 9 13 0 9 2
13 15 16 9 0 13 2 9 13 13 7 9 13 2
7 0 13 9 15 9 15 2
10 13 0 15 13 3 13 15 13 9 2
15 1 9 9 2 16 13 2 13 7 1 9 13 9 15 2
26 3 16 0 13 13 9 9 7 0 9 13 2 13 3 9 13 1 9 13 13 7 9 0 9 13 2
16 9 3 13 0 2 1 15 13 13 9 13 13 9 0 9 2
7 3 13 13 9 15 13 2
18 15 3 3 13 0 15 3 13 15 13 2 7 15 13 0 9 13 2
13 15 15 13 13 9 0 2 3 13 9 0 9 2
22 16 1 9 9 13 9 13 13 2 0 13 9 2 9 15 13 2 3 3 13 13 2
10 6 15 15 2 9 2 9 13 9 2
7 0 9 9 7 9 13 2
9 16 9 13 2 0 0 9 13 2
21 7 15 0 2 16 13 9 13 2 13 9 9 2 15 3 0 9 0 13 9 2
7 3 3 13 9 13 9 2
7 15 9 13 3 9 13 2
5 9 3 13 9 2
22 0 16 9 9 13 9 13 13 13 9 7 13 13 9 9 2 0 13 15 9 9 2
15 3 16 13 9 13 0 9 9 2 15 13 9 9 13 2
16 13 3 13 9 13 15 9 15 9 2 13 13 15 13 9 2
19 9 9 15 3 13 13 3 9 0 9 15 9 2 3 9 9 13 0 2
6 9 13 9 15 13 2
13 15 13 3 1 15 13 2 15 9 9 9 13 2
11 1 9 13 3 9 1 9 9 13 0 2
8 15 13 0 0 15 9 13 2
7 9 1 9 0 13 0 2
13 15 9 9 3 13 13 9 13 2 16 13 13 2
3 0 13 2
11 3 15 13 15 15 13 9 16 13 15 2
16 9 9 16 13 9 0 2 3 9 13 2 7 0 13 13 2
8 9 13 9 9 9 9 9 2
14 13 7 13 3 13 9 2 15 1 9 13 0 9 2
7 3 15 13 16 9 13 2
6 13 0 13 9 9 2
26 9 1 9 16 13 9 2 15 13 9 15 13 2 9 13 9 3 12 3 13 13 2 3 13 12 2
9 9 13 13 9 15 3 13 13 2
10 1 0 9 9 13 1 9 13 9 2
7 15 3 13 15 13 9 2
11 13 9 9 13 9 9 13 0 9 13 2
14 9 13 13 2 9 9 13 2 9 9 3 3 13 2
6 13 9 9 9 0 2
7 15 16 13 9 13 13 2
16 9 13 16 13 0 2 16 9 1 15 9 13 2 3 13 2
16 3 13 9 9 13 2 9 13 0 2 16 0 13 9 13 2
8 15 3 13 13 3 9 13 2
14 0 9 3 3 9 13 2 7 1 9 3 0 13 2
7 9 13 1 9 13 9 2
11 15 16 13 13 13 3 2 9 13 13 2
9 7 13 3 13 3 15 13 13 2
13 15 13 9 0 2 0 7 9 13 1 9 0 2
24 13 9 7 13 9 9 16 13 9 0 13 2 9 0 13 1 15 9 7 13 9 0 9 2
8 0 9 3 13 9 0 9 2
12 9 2 16 13 0 3 13 2 9 9 13 2
6 0 3 13 15 13 2
13 15 2 9 9 2 16 13 3 13 12 13 13 2
3 13 15 2
12 13 16 9 15 2 0 13 7 13 9 9 2
22 3 16 13 16 13 9 2 15 13 13 2 3 7 15 13 2 13 13 0 9 15 2
7 7 3 13 0 9 13 2
20 15 1 15 13 13 15 13 2 15 13 13 9 15 2 7 13 0 13 0 2
12 3 0 0 0 13 2 3 0 0 13 9 2
3 3 13 2
14 7 15 13 15 13 9 13 2 13 16 15 9 9 2
15 1 9 3 9 13 9 7 13 9 0 9 0 13 9 2
10 3 13 15 13 2 16 9 13 0 2
3 15 13 2
14 3 13 9 0 9 7 0 13 9 2 15 0 13 2
4 15 13 9 2
12 3 13 16 13 3 13 15 2 13 13 9 2
14 9 15 13 0 13 9 2 7 13 9 7 13 3 2
15 9 13 13 1 9 9 2 1 9 16 13 2 13 13 2
4 3 13 9 2
3 13 13 2
3 0 13 2
11 16 15 3 13 2 13 0 9 9 13 2
23 9 1 9 13 9 0 13 7 15 1 9 0 13 9 2 15 0 9 13 13 13 9 2
11 15 9 16 13 2 13 9 0 9 13 2
10 15 9 13 13 15 7 13 9 9 2
13 15 16 9 9 3 13 2 0 3 13 9 13 2
8 15 15 9 13 0 9 13 2
14 15 9 0 13 13 13 7 15 0 13 13 0 13 2
25 0 13 9 9 9 13 2 7 13 16 0 9 2 13 13 15 9 9 2 9 16 13 9 13 2
12 7 2 9 16 13 13 9 2 9 13 13 2
7 15 13 9 1 13 13 2
18 6 9 2 3 13 2 15 13 3 0 9 2 9 13 2 13 9 2
12 3 0 13 0 13 2 9 0 16 13 9 2
14 0 9 9 3 13 9 7 13 9 2 9 16 13 2
13 15 13 9 13 13 2 16 0 0 9 13 15 2
8 13 15 2 13 16 15 9 2
18 9 1 9 13 13 9 0 7 9 9 13 2 9 9 9 13 9 2
12 9 16 9 9 13 15 0 13 0 9 13 2
17 3 0 9 16 13 0 2 0 13 0 9 7 15 0 13 9 2
4 13 13 9 2
12 15 13 13 9 7 13 2 3 3 13 13 2
14 0 16 13 15 15 13 2 3 0 13 15 9 15 2
12 9 2 16 13 13 0 9 2 13 9 7 2
11 0 9 13 15 2 7 13 13 0 9 2
6 0 13 3 13 13 2
2 13 2
7 13 9 13 7 13 9 2
17 13 9 9 15 13 2 9 1 13 13 9 7 13 13 0 9 2
8 3 9 1 15 9 15 13 2
14 15 15 13 9 13 0 2 9 16 13 2 9 13 2
23 9 3 16 13 9 7 9 9 13 9 2 9 9 13 1 9 7 9 0 0 13 9 2
21 3 0 3 9 13 2 3 9 15 13 13 9 2 15 15 1 0 13 13 9 2
6 15 13 13 15 9 2
12 15 9 13 13 13 12 7 13 9 0 9 2
3 3 13 2
5 9 13 9 9 2
17 7 0 15 1 9 13 3 13 9 16 0 13 7 15 13 9 2
21 15 13 3 13 9 2 16 13 9 7 13 13 15 2 9 13 2 3 9 9 2
7 3 0 9 9 13 0 2
28 7 16 13 15 13 2 13 9 16 13 9 2 0 1 9 2 9 2 13 13 2 3 16 13 15 9 9 2
20 15 0 16 13 9 2 13 2 3 13 0 13 2 0 7 13 15 3 13 2
6 1 9 13 13 9 2
5 9 13 9 13 2
4 7 0 13 2
15 3 0 9 13 13 1 15 9 0 7 13 13 3 9 2
11 7 2 15 13 9 15 9 2 3 13 2
11 3 13 9 9 13 2 9 16 9 13 2
6 9 0 3 7 0 2
8 3 13 9 0 7 0 9 2
14 1 9 3 13 9 2 13 2 13 2 7 9 13 2
18 9 0 15 9 3 0 13 9 13 9 2 9 7 15 0 0 13 2
14 12 2 13 16 13 15 0 2 9 9 13 13 3 2
12 15 15 13 13 9 9 2 0 3 13 13 2
9 7 3 0 9 2 0 9 13 2
17 13 15 9 0 9 13 9 9 13 0 2 13 13 16 9 9 2
19 13 1 0 15 13 9 2 16 15 0 13 2 16 13 13 0 9 9 2
5 9 0 0 13 2
7 9 1 0 9 9 13 2
7 9 9 13 1 0 13 2
8 9 9 9 9 1 0 13 2
11 3 0 9 9 9 7 0 3 13 9 2
21 7 13 9 16 13 3 9 0 2 9 13 13 2 16 15 1 0 3 9 13 2
11 9 13 7 13 9 13 1 9 0 9 2
16 7 2 3 13 13 1 0 9 2 9 13 13 13 9 15 2
13 15 7 9 16 13 9 2 0 3 13 15 0 2
20 3 13 9 13 9 2 3 9 15 13 7 9 15 2 9 13 13 0 9 2
6 9 13 9 9 13 2
7 9 9 13 3 13 3 2
12 9 13 13 1 15 9 7 9 0 13 9 2
13 0 9 0 3 13 0 2 9 13 0 9 13 2
27 13 9 15 9 9 2 3 13 2 13 1 9 2 3 13 2 0 13 9 13 2 15 0 7 0 0 2
11 15 13 2 16 3 13 2 13 0 9 2
5 9 13 9 13 2
36 1 0 12 9 2 15 9 1 9 9 0 13 13 2 9 13 2 13 0 9 0 2 9 13 0 13 9 13 2 0 9 13 2 7 13 2
11 3 13 9 13 0 1 9 2 13 9 2
7 13 9 9 9 7 13 2
3 13 9 2
9 15 7 13 2 9 0 0 9 2
8 3 0 13 7 9 3 13 2
6 3 0 9 15 13 2
7 1 13 9 13 13 3 2
14 16 3 13 9 0 2 9 7 9 15 13 2 13 2
6 9 1 0 13 9 2
21 15 16 13 0 9 9 7 0 13 13 13 13 2 13 1 9 9 7 3 13 2
6 0 3 9 13 9 2
14 7 16 13 15 13 13 15 2 0 3 15 13 9 2
20 13 9 13 2 16 9 1 0 1 9 0 13 9 2 15 13 3 13 9 2
14 13 9 9 2 13 13 2 3 7 9 3 13 9 2
13 3 13 15 9 13 9 2 0 12 13 0 9 2
6 9 13 9 13 12 2
12 12 13 9 1 9 2 0 13 0 9 9 2
19 15 9 0 0 9 13 0 7 9 13 9 2 9 13 13 7 0 9 2
19 3 9 1 9 13 1 7 9 9 9 13 2 13 9 2 13 0 9 2
8 7 9 13 7 13 13 9 2
7 15 9 13 13 9 9 2
6 0 9 13 9 0 2
22 9 0 13 9 2 16 9 13 13 9 2 0 9 0 9 13 7 0 15 9 13 2
17 15 13 15 2 0 2 3 15 1 9 13 9 7 9 9 13 2
5 9 3 13 13 2
6 9 9 9 13 9 2
8 9 9 13 2 9 3 13 2
10 13 3 7 13 0 0 2 15 13 2
9 13 7 0 2 7 15 15 13 2
15 3 13 0 9 13 13 13 9 2 9 13 16 13 9 2
3 13 12 2
5 0 15 13 3 2
18 15 1 15 9 1 9 13 7 16 13 13 3 9 2 13 1 9 2
8 3 9 9 13 2 9 13 2
7 13 15 0 0 13 9 2
10 16 13 12 2 9 7 0 13 9 2
9 15 13 13 13 9 9 7 13 2
10 15 13 9 9 13 3 1 9 15 2
26 9 9 9 13 0 9 7 13 0 1 9 2 13 9 13 16 0 9 7 9 13 2 7 9 9 2
12 3 13 0 16 12 13 2 16 0 13 13 2
3 15 13 2
12 16 9 13 9 13 2 3 3 13 9 9 2
19 16 15 9 1 9 13 15 7 9 13 9 13 9 2 0 9 13 9 2
32 16 7 13 15 13 9 2 0 15 1 9 9 13 7 15 13 7 0 13 2 0 9 9 13 13 2 16 9 9 13 15 2
21 9 9 13 16 13 2 13 13 2 9 2 1 9 2 16 0 9 13 9 9 2
15 3 3 9 13 9 15 13 15 2 15 13 9 3 13 2
3 3 13 2
12 0 13 9 2 15 15 13 9 1 9 13 2
14 13 15 13 13 7 9 9 2 13 16 9 9 13 2
48 15 2 15 0 9 13 13 9 2 1 15 13 13 9 9 0 12 9 13 9 2 3 1 15 3 13 13 9 9 7 13 3 9 13 7 9 0 9 1 15 13 2 3 3 1 9 13 2
19 15 13 15 13 2 15 0 9 13 13 0 9 2 13 9 0 13 9 2
6 15 16 13 2 13 2
11 16 7 3 2 13 3 15 15 13 0 2
10 3 9 3 13 13 9 2 0 13 2
21 9 0 2 16 15 13 3 13 13 2 9 0 1 9 13 9 7 13 13 9 2
19 15 3 15 9 13 9 2 7 13 0 3 13 2 1 9 13 15 15 2
28 16 16 9 0 9 13 2 16 9 0 2 9 0 3 2 0 13 13 15 0 0 2 7 15 9 13 9 2
19 9 16 15 13 15 7 13 1 15 15 13 0 0 2 3 13 9 9 2
6 15 13 15 13 3 2
16 7 7 13 12 9 13 15 2 3 15 9 7 9 9 13 2
8 9 15 13 13 3 15 0 2
15 15 2 0 15 13 0 9 2 3 9 0 13 9 9 2
16 3 3 13 2 9 2 16 3 13 2 3 15 0 13 9 2
5 13 15 1 13 2
8 0 15 9 13 13 9 13 2
18 9 13 13 13 9 2 3 0 9 1 9 0 9 15 0 3 13 2
12 0 15 13 0 3 13 2 0 16 13 9 2
9 15 3 13 2 13 15 15 13 2
7 13 1 13 0 13 9 2
7 9 0 3 1 9 13 2
3 13 0 2
8 0 9 13 2 0 13 9 2
16 15 3 13 13 3 2 3 9 13 2 13 9 16 13 9 2
9 13 0 9 2 3 13 13 3 2
20 7 15 2 9 16 13 0 2 0 9 9 15 13 7 1 9 13 13 9 2
19 0 9 13 13 2 9 13 2 15 9 13 2 7 0 13 13 13 9 2
17 3 15 13 2 15 0 13 2 9 3 13 2 3 1 9 13 2
10 13 15 15 9 13 2 15 9 13 2
4 15 13 13 2
8 15 13 9 2 15 15 13 2
21 9 0 9 3 13 3 13 13 2 9 7 3 13 2 13 15 3 12 9 15 2
9 13 15 9 13 9 9 0 9 2
8 9 13 1 13 13 13 9 2
11 15 13 1 9 13 9 7 13 9 9 2
17 15 7 13 9 13 9 7 0 13 9 2 7 13 13 0 9 2
10 0 13 9 9 7 9 9 0 13 2
13 13 1 9 15 13 9 2 1 0 9 7 9 2
4 13 15 13 2
8 3 3 15 13 3 3 13 2
14 3 7 0 3 13 0 2 7 0 9 0 13 0 2
6 9 1 9 0 13 2
6 9 15 0 9 13 2
8 9 3 15 13 2 3 13 2
6 13 3 0 7 13 2
9 15 3 13 9 7 0 13 9 2
6 7 9 13 0 9 2
6 13 7 9 13 9 2
8 9 1 9 13 7 9 13 2
4 3 0 13 2
7 13 16 9 9 13 15 2
3 13 15 2
5 9 3 13 15 2
18 7 15 13 9 15 12 13 9 9 13 0 15 7 9 9 13 13 2
5 3 13 0 9 2
10 7 7 3 13 7 3 13 13 13 2
13 15 13 9 3 13 2 15 1 9 0 13 9 2
8 3 0 13 9 2 3 13 2
8 9 13 9 13 9 9 13 2
6 3 13 3 16 13 2
7 7 15 9 13 0 9 2
10 15 2 15 13 3 0 2 13 9 2
12 15 13 9 15 2 13 9 16 0 9 13 2
3 13 15 2
5 15 3 13 13 2
11 3 13 9 9 7 1 9 0 9 13 2
14 3 13 0 15 1 9 13 2 7 0 0 13 9 2
4 13 3 15 2
11 16 13 2 13 9 1 9 9 13 9 2
3 9 13 2
4 13 13 3 2
18 16 13 0 2 13 15 3 2 9 16 13 7 13 2 9 16 13 2
9 9 13 2 3 13 13 2 13 2
4 13 3 9 2
7 1 9 15 13 9 9 2
11 9 13 9 7 2 15 13 15 2 9 2
7 3 1 9 9 13 15 2
7 13 2 15 13 2 9 2
9 13 13 2 0 16 3 13 15 2
6 9 13 3 15 13 2
11 13 15 9 0 15 7 0 0 9 9 2
15 15 2 9 1 9 9 16 13 13 2 3 13 9 13 2
5 15 15 0 13 2
19 3 1 9 13 9 3 0 7 9 13 9 2 9 13 16 9 9 13 2
9 0 9 9 2 7 0 13 9 2
7 0 13 13 7 3 13 2
6 15 9 3 13 9 2
8 9 13 2 16 9 13 13 2
8 9 16 3 13 2 13 9 2
13 3 13 13 9 3 2 3 3 0 3 13 9 2
14 7 0 16 9 13 2 13 15 9 15 13 13 15 2
26 9 15 16 13 9 9 7 0 3 13 9 2 13 1 13 1 0 13 15 2 13 9 13 15 0 2
32 15 16 1 9 0 13 13 7 0 1 9 0 9 2 13 15 2 15 13 3 13 13 2 13 9 9 7 0 13 9 9 2
15 13 15 13 9 9 13 9 1 9 3 7 1 9 13 2
23 3 9 3 9 13 2 3 9 9 13 2 1 15 13 9 0 13 2 9 13 13 3 2
22 16 13 9 2 16 13 9 2 9 13 9 3 13 1 9 13 2 13 1 9 9 2
15 16 13 13 2 9 9 13 2 9 13 2 16 9 13 2
19 9 13 2 3 13 9 13 7 9 13 9 2 13 12 15 9 9 13 2
13 13 1 15 9 9 7 9 13 2 15 9 13 2
9 9 13 9 9 7 13 1 9 2
9 0 0 13 9 2 16 0 13 2
8 13 9 3 9 13 0 9 2
19 1 0 9 3 13 9 2 16 13 9 13 9 2 16 15 9 13 9 2
13 7 0 9 3 7 13 9 13 3 3 13 13 2
9 9 13 9 2 7 3 13 3 2
17 3 7 15 13 2 15 3 13 2 7 15 3 13 2 13 9 2
12 15 13 0 7 13 2 9 0 16 15 13 2
11 9 7 13 0 7 9 13 7 9 15 2
8 13 15 13 15 1 15 13 2
11 15 13 13 3 0 9 0 3 15 13 2
19 9 13 1 15 0 2 15 1 0 13 7 0 9 9 13 13 13 9 2
9 7 15 9 2 0 2 9 13 2
10 15 3 13 9 0 2 15 13 13 2
11 1 9 9 0 16 13 9 2 9 13 2
14 15 16 15 9 0 13 15 2 3 13 1 9 0 2
19 15 16 15 13 2 0 15 3 13 9 2 7 15 13 7 15 15 13 2
9 15 15 13 2 15 15 3 13 2
7 9 1 0 13 9 9 2
7 15 9 0 13 13 15 2
9 9 1 9 13 13 2 9 9 2
13 15 9 15 13 16 3 2 9 12 15 13 9 2
16 3 0 9 7 0 13 9 2 1 0 3 9 16 3 13 2
31 7 16 9 13 0 15 2 9 13 7 9 9 13 2 16 1 9 9 7 9 9 2 1 15 3 13 2 9 15 13 2
3 9 13 2
4 9 9 13 2
6 3 15 0 13 9 2
9 0 13 15 3 13 7 15 13 2
6 3 9 9 13 15 2
12 15 13 9 9 2 16 13 9 3 13 9 2
17 9 1 9 15 13 0 9 9 16 13 2 13 7 3 0 13 2
16 15 13 3 9 3 3 13 9 2 9 13 13 1 0 9 2
3 13 9 2
10 15 15 13 3 7 9 13 9 13 2
3 3 13 2
8 3 13 9 3 16 13 13 2
9 7 16 13 2 16 13 13 0 2
14 3 9 9 13 3 13 2 1 13 0 16 13 15 2
6 3 13 3 9 15 2
6 9 7 13 13 3 2
24 3 15 13 2 15 2 16 13 13 2 13 2 3 13 9 0 0 9 2 3 13 13 9 2
8 3 15 13 0 15 15 13 2
4 3 3 13 2
8 3 15 13 0 7 0 13 2
3 13 3 2
12 13 16 13 9 2 15 13 2 16 13 0 2
13 9 3 0 0 13 2 16 13 9 1 9 12 2
21 15 9 0 1 13 13 2 3 15 13 0 15 13 13 13 0 7 9 13 9 2
7 13 9 9 2 3 9 2
12 15 13 13 9 9 13 9 9 2 9 13 2
11 9 15 15 3 13 2 3 9 13 9 2
18 9 0 9 9 13 2 13 9 1 9 13 0 7 9 13 9 3 2
5 13 13 16 13 2
7 3 13 9 13 3 13 2
18 9 16 13 15 0 13 9 7 9 13 15 2 15 13 13 0 9 2
6 16 3 13 2 13 2
3 3 13 2
15 15 2 15 13 9 2 3 13 9 13 15 2 3 13 2
11 9 13 1 0 13 13 13 7 9 13 2
7 3 0 15 13 13 0 2
12 3 15 13 13 1 9 15 2 0 13 9 2
17 9 9 7 9 9 13 2 9 9 2 9 9 2 9 0 9 2
8 9 13 2 3 0 13 13 2
4 9 13 9 2
8 6 0 2 3 13 13 0 2
10 16 0 13 15 13 2 0 13 9 2
8 9 13 15 3 13 9 13 2
14 9 1 9 13 2 3 13 9 9 16 15 3 13 2
6 3 13 9 13 9 2
7 7 9 13 2 13 9 2
12 9 9 9 13 15 13 7 9 0 9 13 2
7 9 9 9 13 15 13 2
15 13 13 15 15 3 13 13 2 13 16 9 1 9 13 2
13 9 9 0 16 13 9 2 13 9 13 13 3 2
14 9 3 13 12 13 9 2 3 7 13 3 9 13 2
9 3 13 13 15 9 0 13 0 2
7 7 3 1 9 13 13 2
9 9 13 13 2 7 13 13 9 2
21 15 16 0 15 1 9 13 2 13 3 15 9 3 13 0 2 3 15 13 13 2
22 13 15 15 13 2 7 13 13 2 3 16 13 13 15 0 2 13 15 0 9 9 2
10 9 15 9 16 13 13 15 13 13 2
4 13 9 9 2
21 7 9 9 0 13 3 2 7 15 0 13 1 15 9 2 3 3 13 9 9 2
9 16 3 9 13 2 9 13 0 2
7 13 3 2 16 3 13 2
11 13 9 16 13 15 9 2 9 9 13 2
21 3 9 0 3 13 9 13 15 2 16 3 13 13 9 0 7 9 0 13 13 2
12 0 13 15 9 13 2 0 3 16 13 9 2
6 3 13 9 13 9 2
6 3 0 3 13 13 2
4 15 13 9 2
11 13 0 3 2 3 0 9 13 0 9 2
15 13 15 9 2 15 13 9 2 7 3 15 13 9 15 2
6 13 9 15 13 9 2
14 7 3 13 9 2 9 15 0 0 1 0 13 9 2
5 15 13 2 13 2
3 13 9 2
21 15 2 3 13 15 9 9 2 3 13 0 9 13 2 16 9 13 2 3 13 2
9 9 9 9 0 3 13 0 13 2
44 7 7 9 0 9 9 3 3 9 13 7 13 9 9 13 2 15 9 9 0 2 16 9 9 9 0 13 2 13 3 9 9 0 9 13 9 13 7 3 9 13 9 13 2
23 9 7 0 13 2 15 13 2 16 1 0 3 0 9 9 9 13 9 7 1 9 13 2
38 15 9 1 9 9 9 1 0 9 13 1 9 2 3 1 9 9 1 0 13 2 13 9 1 9 15 13 7 3 0 9 1 0 9 1 9 13 2
10 12 1 15 9 9 9 13 9 9 2
29 15 0 9 7 9 13 2 1 15 0 9 9 13 9 13 2 3 9 7 3 1 15 0 0 13 13 9 0 2
20 7 9 15 7 0 2 7 9 7 9 2 1 0 9 13 3 1 9 9 2
15 9 9 12 0 9 9 1 9 9 9 13 9 9 9 2
9 9 0 9 13 13 9 3 13 2
23 15 9 9 0 3 0 9 13 15 13 0 7 0 2 7 1 15 12 9 9 15 13 2
15 9 9 0 15 9 13 2 9 1 9 0 2 9 0 2
9 7 15 3 1 0 9 0 13 2
30 9 9 9 1 9 9 7 9 7 9 0 13 2 16 3 13 15 3 1 0 0 7 7 1 9 9 7 0 13 2
13 0 7 13 9 9 7 13 13 3 7 3 13 2
27 1 9 9 13 0 2 0 9 7 9 9 2 0 9 13 1 9 13 2 9 15 1 9 1 9 13 2
8 9 13 3 0 9 3 9 2
40 7 9 7 0 0 9 13 3 0 13 2 16 9 9 9 13 2 15 9 9 15 9 3 0 9 9 9 13 13 7 13 2 13 1 13 0 0 15 9 2
35 13 9 2 3 3 13 15 0 9 13 2 9 13 0 2 0 9 9 0 2 15 1 9 2 7 9 0 3 9 2 15 1 9 13 2
14 9 9 9 9 7 9 2 9 9 9 2 13 13 2
32 9 2 0 9 0 2 0 1 9 0 9 2 1 9 9 9 0 13 9 13 7 9 9 1 9 9 0 9 0 9 13 2
25 3 15 9 2 13 7 0 9 9 2 9 15 0 9 13 7 3 0 9 3 9 9 13 13 2
19 9 3 0 15 9 3 3 7 9 2 7 7 7 0 9 3 13 9 2
10 2 0 15 9 13 1 0 9 9 2
9 15 13 9 9 13 0 0 2 2
36 13 13 9 9 9 9 9 9 9 9 12 2 9 0 3 1 9 9 2 9 9 1 9 0 2 3 3 9 13 2 3 3 3 13 13 2
61 7 16 9 13 13 2 16 9 9 2 9 0 9 2 1 13 0 9 9 1 9 7 0 15 3 9 13 13 2 13 9 7 3 9 9 2 15 3 0 9 13 13 2 13 7 13 3 0 15 7 0 9 2 13 13 16 15 9 9 13 2
26 9 15 13 3 9 1 0 9 1 9 0 7 9 0 9 2 13 7 9 9 3 7 13 3 13 2
27 3 13 7 3 7 3 9 13 2 13 9 0 2 3 3 13 9 15 7 9 13 2 7 7 3 13 2
36 7 16 9 9 0 7 9 7 13 9 13 15 3 13 2 13 16 1 0 9 9 13 3 13 9 7 0 3 0 1 9 3 1 9 13 2
26 0 9 0 13 13 2 1 9 0 9 2 7 16 9 0 3 15 13 9 9 1 0 9 3 13 2
33 0 13 3 0 9 13 13 0 9 15 0 0 0 7 3 3 13 9 15 9 13 2 15 9 1 15 9 13 1 9 9 13 2
27 7 7 1 9 9 1 9 1 9 3 0 13 7 15 9 0 3 13 15 13 1 9 15 0 9 13 2
4 0 9 13 2
10 12 9 13 9 9 13 1 9 13 2
19 9 3 0 9 13 0 9 9 9 0 13 13 2 16 0 9 1 9 2
37 13 3 9 1 9 1 9 9 9 3 0 1 0 9 1 0 9 9 0 9 9 7 13 13 2 3 13 2 13 3 7 9 9 1 9 9 2
17 9 1 13 9 9 1 9 7 3 1 9 13 13 9 9 13 2
26 16 7 3 13 15 9 7 15 13 2 3 13 16 0 9 13 2 15 3 9 7 0 0 7 13 2
17 3 9 13 9 13 2 13 9 2 9 3 9 9 0 3 13 2
22 13 9 15 3 9 9 3 7 1 9 7 1 9 13 2 3 3 13 13 7 13 2
5 9 0 12 13 2
8 0 9 9 7 9 3 13 2
38 9 13 13 3 9 9 13 13 7 13 2 3 16 9 13 2 9 9 7 7 9 0 7 2 16 13 9 13 2 9 13 9 7 9 13 13 13 2
15 9 7 9 9 3 13 13 15 13 15 9 2 15 13 2
22 7 3 3 0 7 13 2 1 9 9 9 9 13 13 15 13 2 16 0 7 9 2
59 7 13 9 15 9 9 9 2 15 7 0 9 13 2 7 7 0 3 7 0 9 0 1 9 15 1 9 0 9 13 2 1 0 15 13 2 15 15 13 13 2 3 16 9 9 13 9 9 1 9 13 7 1 9 13 13 9 13 2
27 13 7 0 9 15 13 2 7 9 13 9 1 9 13 0 3 1 15 7 9 0 9 0 13 9 13 2
30 13 7 13 9 1 9 13 7 1 9 7 9 2 15 9 13 2 9 9 9 13 2 13 9 12 9 13 12 9 2
45 0 9 13 15 13 7 1 9 9 7 1 0 3 13 2 13 3 13 3 3 9 2 7 7 9 13 9 7 1 0 9 2 9 9 15 3 0 2 9 9 13 3 7 13 2
34 15 9 16 9 1 9 2 9 3 3 1 9 13 2 9 13 12 9 15 13 2 16 9 13 2 9 0 9 13 0 9 9 13 2
18 9 3 3 13 9 13 2 16 9 0 13 13 2 3 9 9 13 2
15 13 15 9 9 0 1 9 9 1 9 9 1 15 13 2
55 7 16 13 9 1 9 1 9 9 13 0 7 9 7 9 13 1 9 2 9 0 1 9 13 2 1 9 13 9 13 13 7 15 13 2 3 0 15 9 2 0 13 13 7 13 2 16 7 15 7 0 0 9 13 2
34 7 3 3 9 0 9 13 2 0 0 9 7 15 13 13 13 0 9 13 2 16 0 9 13 9 9 3 13 13 1 9 15 13 2
30 13 1 9 7 9 9 0 7 9 2 16 0 7 0 2 0 9 13 2 15 0 9 13 3 1 9 9 9 13 2
27 7 9 9 13 13 2 7 9 9 9 13 2 16 9 9 13 2 1 0 15 0 3 1 9 9 13 2
14 7 3 12 3 9 13 13 13 3 15 9 13 9 2
26 3 0 2 1 15 9 9 15 9 0 2 16 13 13 2 9 9 3 13 2 15 0 9 3 13 2
39 13 1 9 9 16 9 9 13 2 15 0 1 9 13 7 0 9 13 13 2 7 0 7 9 9 13 2 0 13 15 2 0 3 1 9 13 13 13 2
38 15 9 9 9 9 9 2 15 13 2 7 0 9 9 0 13 13 9 13 7 1 9 9 13 2 3 3 1 0 15 7 1 9 7 1 9 9 2
36 7 16 9 9 0 9 1 12 9 13 13 1 9 13 2 9 1 9 13 3 15 3 7 13 13 2 3 13 16 13 9 7 9 9 0 2
13 9 13 2 16 15 13 3 13 0 7 1 9 2
16 1 0 7 9 13 3 13 13 1 9 9 2 15 9 13 2
20 9 13 1 0 13 2 13 9 7 13 15 13 12 9 13 2 13 13 2 2
19 13 15 12 1 0 13 0 9 1 9 0 9 13 9 0 9 9 13 2
37 13 15 13 13 15 1 9 13 2 16 13 0 7 15 9 3 3 9 13 2 9 9 9 9 13 2 13 13 7 15 7 13 13 0 9 13 2
32 1 15 16 9 0 9 13 2 9 1 9 7 9 13 2 1 9 9 3 0 3 9 13 2 16 1 13 9 1 9 13 2
7 3 13 9 9 13 13 2
29 0 13 13 7 15 13 2 3 9 9 13 13 7 0 9 9 15 13 2 7 9 0 0 0 9 9 9 13 2
11 7 3 0 7 0 9 0 0 9 13 2
27 13 1 9 9 2 16 9 0 9 13 13 2 13 1 0 1 9 7 9 9 9 12 3 9 3 13 2
23 3 16 1 9 9 9 13 7 13 0 0 9 13 15 13 13 1 9 2 3 13 13 2
29 3 7 1 0 9 13 9 9 9 9 15 2 13 13 3 1 15 9 9 7 3 9 9 13 2 13 13 13 2
38 1 9 9 9 0 9 9 2 15 1 9 1 9 13 2 13 12 9 9 0 7 15 9 9 7 9 13 13 9 0 7 13 9 9 1 0 13 2
46 9 9 9 3 0 7 0 9 7 0 3 13 13 3 2 7 3 3 13 15 1 0 9 13 2 9 2 15 15 9 7 1 9 9 1 9 13 13 2 13 13 7 1 9 13 2
20 13 3 9 13 9 9 7 0 7 1 0 9 9 7 9 9 3 3 9 2
21 0 3 3 2 16 1 9 9 3 13 2 9 13 13 1 0 9 1 9 15 2
19 7 3 3 0 9 1 9 13 1 0 9 13 2 16 1 9 9 13 2
38 7 3 3 12 7 12 9 2 16 2 1 9 9 13 2 9 13 2 9 9 7 9 9 13 13 7 9 2 3 9 1 9 13 2 0 13 13 2
14 7 9 3 0 9 9 13 1 9 13 13 7 0 2
24 9 2 15 13 9 3 13 2 7 9 13 2 15 9 7 9 13 2 16 13 9 9 13 2
13 12 0 9 9 13 7 9 1 15 13 13 13 2
42 1 15 9 9 7 9 0 9 2 16 13 1 0 13 9 2 9 0 13 7 9 13 13 13 13 7 2 3 7 9 13 13 2 9 15 13 13 13 2 3 13 2
28 9 1 9 9 13 16 0 0 7 9 0 13 2 9 0 2 1 15 9 13 2 13 0 9 0 9 13 2
41 3 7 0 9 9 13 7 1 0 13 2 9 9 1 9 13 9 7 3 0 13 7 13 0 9 9 9 9 2 15 13 13 2 13 0 9 9 7 9 13 2
21 9 3 7 9 0 9 9 7 0 2 3 3 13 9 13 2 13 0 0 9 2
11 7 7 0 3 9 9 9 7 9 13 2
31 9 7 9 9 9 7 9 9 1 9 2 15 13 2 13 1 9 2 9 3 13 15 9 9 7 15 7 9 13 13 2
6 9 7 13 9 13 2
28 0 1 9 13 2 16 3 15 0 7 0 7 13 7 3 3 13 2 9 7 9 7 9 3 1 9 13 2
28 13 7 3 9 3 9 15 9 2 9 2 9 2 9 1 9 0 2 3 9 7 9 7 9 2 9 0 2
36 13 7 9 9 12 15 9 1 0 9 13 2 9 7 1 9 9 13 2 1 15 9 7 9 13 15 13 1 9 7 1 0 9 9 13 2
9 0 3 9 3 13 1 9 13 2
60 7 0 9 1 0 7 0 9 9 13 3 7 13 1 9 15 9 9 7 0 9 13 2 16 15 0 9 1 9 9 9 13 13 13 15 1 9 7 9 15 13 2 1 15 3 0 9 9 2 9 2 13 13 2 16 13 0 9 13 2
12 7 3 9 3 0 13 2 3 13 9 13 2
31 7 7 3 7 3 13 0 3 13 13 9 2 3 16 0 1 9 13 2 16 1 0 9 13 16 7 1 12 9 13 2
24 15 9 9 7 9 0 7 7 9 9 3 13 13 1 9 15 9 7 0 3 1 9 13 2
40 9 3 7 9 13 3 13 7 9 0 2 15 9 9 7 9 9 13 2 13 13 9 7 3 13 2 3 0 3 1 9 13 2 3 7 1 15 13 13 2
25 9 9 3 7 3 1 13 9 1 9 15 13 1 3 0 9 9 9 9 7 9 13 3 13 2
14 3 13 13 13 9 2 1 0 7 3 1 0 9 2
15 0 9 12 13 2 0 2 0 2 0 2 3 9 0 2
26 15 13 9 1 9 13 2 16 15 9 13 2 7 9 9 13 9 2 16 1 0 7 13 0 13 2
16 13 7 0 9 9 0 0 2 16 9 0 1 0 9 13 2
8 15 13 0 0 7 9 13 2
19 3 3 13 13 2 16 1 0 9 9 9 7 13 9 3 9 13 13 2
16 1 9 0 7 13 0 7 13 7 7 1 0 9 0 13 2
4 9 3 13 2
16 7 9 3 15 2 7 3 0 7 3 9 2 13 9 13 2
19 9 0 2 16 12 9 13 9 13 9 9 13 2 15 0 7 13 9 2
22 15 3 2 16 13 9 0 13 2 0 15 13 2 16 13 1 9 1 0 13 13 2
20 12 9 3 13 1 9 0 13 2 3 0 3 9 13 1 0 13 9 13 2
11 9 2 16 15 13 9 2 13 9 13 2
43 9 9 13 2 3 16 0 2 0 9 13 2 1 0 9 9 0 9 13 2 16 13 1 0 9 13 1 9 2 3 13 13 7 2 3 1 9 2 7 7 9 13 2
52 7 1 9 0 7 1 9 7 1 9 0 9 9 13 2 7 9 2 7 7 1 9 3 7 9 15 9 0 3 13 13 13 2 0 15 13 2 3 7 9 0 7 9 9 7 15 9 7 15 9 13 2
19 0 9 2 3 9 9 9 7 16 9 1 0 9 13 2 3 13 13 2
30 15 7 2 9 3 9 9 7 0 13 7 1 9 13 2 1 0 9 13 2 7 7 13 1 0 7 15 9 13 2
26 9 0 3 3 9 7 9 2 15 9 9 7 13 2 3 0 7 0 9 2 15 9 13 2 13 2
11 9 9 1 9 1 0 9 0 9 13 2
12 9 7 3 13 9 3 9 9 7 13 13 2
5 3 3 15 13 2
18 9 3 7 9 13 3 13 2 16 16 0 9 9 3 9 9 13 2
22 7 0 0 3 0 13 9 0 13 13 0 9 13 2 15 13 9 0 9 13 13 2
14 9 7 9 7 1 9 7 15 0 9 0 7 13 2
18 9 12 9 9 13 13 3 1 9 9 13 7 15 15 9 9 13 2
58 12 9 1 12 9 2 12 9 13 13 2 13 3 1 12 13 2 0 7 3 2 16 13 2 13 12 0 2 15 13 12 9 2 9 7 3 12 12 9 3 3 13 2 16 9 7 9 9 0 0 9 15 15 9 13 1 9 2
26 12 0 9 1 12 1 12 0 13 2 0 7 12 7 12 7 12 7 12 9 2 12 3 0 9 2
23 7 9 9 0 16 3 1 9 0 9 3 0 9 13 2 9 13 13 0 1 9 15 2
9 9 9 0 13 1 12 9 13 2
34 7 15 1 0 3 9 1 9 7 9 0 0 3 13 16 15 13 2 13 7 7 9 9 9 15 2 15 9 9 15 9 1 9 2
45 9 9 15 3 13 2 16 13 9 9 9 1 9 13 13 7 9 9 1 0 13 2 3 0 9 13 13 2 15 1 13 13 2 3 9 15 13 13 2 16 0 15 13 0 2
22 1 15 3 9 9 3 9 9 9 2 16 9 15 13 13 3 13 2 0 9 13 2
8 1 15 15 9 0 13 9 2
24 15 3 13 9 13 13 15 13 7 1 15 1 9 2 3 9 13 13 9 7 9 9 13 2
7 1 13 9 0 3 13 2
26 7 13 7 15 13 3 1 9 13 7 15 0 9 3 13 2 1 13 13 2 0 9 0 7 9 2
17 15 9 2 16 1 15 3 13 2 15 7 9 15 9 13 13 2
16 13 7 15 15 9 9 13 0 9 2 16 15 0 9 13 2
14 13 3 2 3 13 0 9 13 2 7 1 0 13 2
10 0 9 0 13 2 1 15 7 0 2
18 9 13 9 13 9 7 9 9 2 15 13 3 13 12 7 12 13 2
22 7 3 7 13 9 9 13 13 13 7 2 16 3 1 15 0 9 7 9 9 13 2
10 9 9 9 0 1 9 0 13 13 2
29 13 3 2 16 1 9 9 7 3 13 9 2 9 1 9 13 3 13 2 15 7 9 13 2 3 9 9 13 2
18 9 9 1 15 9 0 9 13 2 15 9 13 13 1 9 9 13 2
21 13 9 1 9 0 0 7 2 15 9 3 0 3 7 9 13 9 7 9 13 2
22 13 9 9 13 13 9 2 16 9 0 1 0 9 9 15 9 13 9 7 13 13 2
32 15 7 9 1 9 0 2 9 3 7 9 9 7 13 2 7 9 9 7 9 7 9 2 3 9 9 7 9 9 7 9 2
23 7 7 0 0 9 3 13 13 2 16 1 9 15 9 7 0 7 13 7 13 9 13 2
25 9 9 1 9 9 7 13 13 7 2 16 15 0 9 3 13 2 15 9 1 9 15 9 13 2
9 1 9 9 0 0 7 13 13 2
44 16 13 9 1 0 9 1 9 2 3 16 3 13 2 0 1 15 9 13 7 9 3 9 0 13 0 9 2 15 0 13 9 9 13 2 1 9 0 13 7 9 1 15 13
25 15 9 7 9 13 9 0 9 1 0 9 0 13 7 13 9 1 0 9 15 13 8 9 9 13
12 15 2 16 3 9 9 13 13 2 1 9 13
24 13 9 9 7 0 9 15 0 9 13 16 15 15 1 15 13 13 7 15 1 15 9 0 13
12 15 3 0 13 9 13 2 9 1 0 9 13
9 3 3 13 3 13 16 1 15 13
13 9 0 13 9 13 7 9 3 12 1 9 9 13
20 9 9 13 7 3 9 13 0 9 1 15 13 7 9 9 9 1 15 13 13
9 15 9 1 15 3 1 9 13 13
26 15 9 9 3 13 13 0 9 9 0 7 0 9 13 9 9 13 2 16 1 0 9 0 9 13 13
7 15 13 9 15 1 15 13
44 16 0 9 9 1 0 9 13 1 15 13 13 7 3 3 3 13 1 15 15 13 9 7 1 9 13 2 9 9 2 7 13 1 0 9 9 2 9 13 13 7 3 9 13
33 15 9 7 9 0 9 9 9 13 7 1 15 15 13 13 1 9 13 7 9 1 9 7 0 9 16 1 9 1 15 13 13 13
5 1 15 9 9 13
16 3 9 13 7 1 0 9 9 8 9 9 9 1 12 9 13
12 9 1 9 9 12 9 7 9 12 9 13 13
24 3 1 0 9 9 15 9 13 15 9 1 9 13 2 9 7 0 9 7 9 0 9 9 13
19 15 9 7 9 1 9 9 9 13 13 7 9 15 1 9 9 13 9 13
15 15 9 2 16 9 7 9 13 2 3 12 9 12 9 13
9 9 13 3 0 1 0 7 9 9
6 15 16 0 13 9 13
17 0 7 2 16 1 15 9 13 13 2 16 13 13 13 1 9 13
7 3 9 0 1 0 9 13
15 3 0 13 9 13 2 0 9 9 0 9 0 1 9 13
17 9 3 1 15 9 1 9 9 13 2 15 13 1 0 9 13 13
51 3 9 13 9 0 9 13 13 13 15 9 16 2 16 13 2 9 2 15 13 8 2 9 9 2 13 7 9 13 2 16 3 13 2 9 9 13 2 15 0 15 9 1 9 13 13 2 7 9 0 13
31 9 9 9 7 9 9 15 15 1 9 13 7 13 13 2 7 16 13 9 0 1 9 9 7 9 9 13 2 12 9 13
16 15 13 7 0 9 1 9 13 2 1 15 9 1 9 9 13
8 15 15 7 0 9 1 9 13
4 15 9 9 13
11 15 1 9 7 9 9 16 13 2 3 13
22 16 1 15 9 9 9 13 2 13 1 9 9 9 1 9 0 3 3 12 9 12 13
14 9 1 9 3 0 1 9 9 2 15 3 13 2 13
29 1 15 9 0 9 9 13 0 15 7 0 2 9 3 12 3 0 2 1 0 9 0 2 16 3 3 3 13 13
8 1 15 9 9 1 9 15 13
9 1 0 9 1 9 0 9 9 13
6 9 13 9 9 3 12
6 9 9 13 13 0 9
13 7 9 7 9 9 3 15 13 16 9 1 9 13
12 7 16 9 13 2 9 0 9 12 9 13 13
6 1 15 0 9 9 13
14 3 0 9 15 3 13 13 0 9 13 7 9 9 13
13 9 0 1 9 7 9 9 13 1 9 9 9 13
48 16 15 15 3 1 9 1 0 13 7 3 1 9 1 0 9 13 2 7 3 0 3 3 15 1 9 13 7 9 13 13 13 13 13 2 3 9 12 15 0 13 2 9 13 2 9 13 13
16 15 7 9 0 9 1 0 9 7 15 15 1 9 13 13 13
20 1 0 9 9 13 7 9 1 9 13 13 2 16 15 9 9 1 9 9 13
70 15 3 13 2 16 13 13 2 9 2 16 9 13 0 9 13 7 3 3 13 13 2 3 1 15 15 13 7 13 9 2 3 9 1 9 13 7 9 13 2 15 3 2 16 9 9 13 2 9 13 2 0 9 2 15 3 0 1 0 9 9 13 2 0 9 3 1 9 9 13
54 3 2 16 3 9 13 2 9 9 13 2 1 0 9 3 13 13 2 7 13 1 9 3 3 13 16 1 9 0 1 0 9 9 0 9 1 15 15 1 9 7 9 9 13 13 13 2 16 1 0 9 0 9 13
10 13 3 9 12 12 0 1 9 13 13
22 3 15 9 13 9 2 16 3 13 9 2 7 13 9 0 2 9 15 9 3 9 13
12 1 15 15 13 9 9 1 15 13 13 12 12
49 15 9 1 8 2 9 2 15 1 9 0 13 1 9 2 9 2 9 2 9 2 9 2 9 2 9 2 15 13 0 9 7 9 13 2 0 13 13 0 15 9 1 9 7 9 9 0 13 13
9 3 3 3 13 2 9 2 9 0
8 3 3 7 9 15 0 15 13
7 15 1 9 15 13 13 9
16 13 0 9 3 13 2 13 3 15 0 9 13 9 0 3 13
6 9 15 13 2 9 13
3 15 3 13
1 13
21 3 3 3 1 9 13 2 13 0 9 9 2 13 7 13 9 1 9 0 15 0
25 1 9 15 2 9 2 13 9 9 3 3 13 2 1 15 13 9 15 15 1 15 0 3 3 13
11 9 9 9 9 7 9 13 13 15 9 13
20 3 15 3 0 13 2 16 8 2 9 9 9 2 9 0 9 13 9 0 13
21 13 2 13 15 3 1 15 9 0 9 16 9 0 0 9 9 0 3 0 9 13
22 13 9 9 1 15 2 9 2 0 7 0 2 3 13 9 0 9 7 3 9 15 9
33 3 3 15 0 9 9 2 3 9 9 2 3 9 9 2 3 9 0 0 2 3 15 0 13 9 9 2 3 15 9 7 9 13
15 13 3 9 16 8 2 9 9 13 16 15 9 0 9 13
3 9 0 13
25 13 13 1 15 9 9 8 2 9 2 0 9 2 9 2 9 2 13 13 1 9 8 2 9 0
15 0 9 9 8 2 9 7 8 2 9 9 13 13 9 0
11 7 3 15 0 3 9 13 13 9 15 9
29 13 7 15 9 9 9 2 3 13 1 9 2 3 1 9 13 2 15 1 9 9 3 15 13 13 2 9 2 13
12 13 2 7 13 3 1 13 2 7 1 13 9
27 13 2 9 13 2 15 13 0 2 13 1 0 9 0 9 3 13 13 2 7 3 15 15 9 7 9 13
18 9 13 1 9 1 9 0 1 9 9 13 2 13 1 9 0 9 9
21 15 7 9 9 7 9 9 1 9 7 3 1 9 13 0 15 3 9 9 0 13
16 3 15 15 15 3 3 13 13 13 0 1 9 7 13 16 13
25 3 3 13 2 16 3 9 3 0 2 3 13 2 3 0 0 13 13 15 15 3 9 13 13 13
31 3 3 15 13 15 15 13 13 2 13 2 7 13 3 16 3 13 2 0 0 7 0 9 13 16 13 15 1 9 0 13
36 7 15 13 2 9 2 15 3 3 13 2 16 7 3 9 9 13 9 0 7 3 13 9 9 13 9 9 0 13 2 16 13 2 16 13 9
2 13 3
13 9 13 0 15 0 9 0 2 15 3 15 13 13
32 13 15 15 1 9 9 15 0 13 1 1 9 12 9 9 2 3 16 0 9 9 9 3 3 0 13 3 0 9 13 9 13
34 3 13 13 15 15 15 9 0 9 2 0 9 13 13 15 1 9 0 3 13 2 16 15 9 9 0 3 15 13 9 13 15 13 13
25 16 15 9 9 15 0 13 0 9 13 13 2 13 15 9 0 9 0 9 2 9 2 9 13 13
20 9 13 2 9 13 2 9 13 15 3 15 3 3 13 7 3 13 7 3 13
6 13 15 3 9 15 0
14 3 13 3 15 13 3 1 9 3 15 1 9 9 0
8 13 3 0 15 9 7 9 9
3 3 13 13
2 15 13
4 13 2 16 13
11 13 7 13 3 1 9 15 15 15 3 13
3 3 9 13
4 15 9 0 13
4 1 15 9 13
21 15 15 13 9 7 1 9 0 9 13 2 7 15 9 13 13 2 15 3 9 13
25 13 13 0 9 0 15 15 15 9 13 7 15 15 15 9 9 1 9 15 1 0 9 13 13 13
9 15 15 9 3 3 9 0 13 13
36 9 0 0 9 13 7 13 2 13 15 15 15 1 15 13 8 13 2 16 15 15 13 15 15 3 0 7 0 9 1 15 15 9 13 13 13
10 15 16 3 13 2 9 2 13 3 13
4 13 3 1 9
2 13 9
1 13
9 3 3 15 9 0 15 0 9 13
11 13 15 3 0 0 2 16 3 2 3 0
2 13 9
12 0 15 9 13 2 3 1 15 7 15 9 13
6 15 13 3 3 3 13
8 3 13 2 3 13 2 3 13
11 3 13 3 1 0 9 0 9 13 9 0
20 7 3 15 9 13 2 9 2 13 13 2 3 0 15 9 2 7 13 9 13
26 16 0 9 0 15 9 1 9 7 9 0 13 13 2 13 9 0 0 9 9 7 9 0 9 3 13
22 3 2 3 15 13 2 1 15 15 13 2 16 13 9 0 1 0 9 9 9 13 13
26 3 3 3 9 0 0 13 2 9 9 0 2 9 9 2 9 0 9 2 9 0 1 9 7 9 13
35 15 9 2 16 15 15 13 0 2 7 15 15 9 7 9 0 0 13 2 13 3 13 2 13 15 15 13 1 9 0 2 1 0 9 0
13 7 16 15 13 13 2 13 1 9 0 0 9 9
22 16 15 2 16 15 3 3 13 2 13 2 13 1 9 0 9 0 7 0 9 9 0
4 15 13 2 9
11 3 13 15 15 13 13 15 3 0 9 13
6 13 1 9 13 9 9
6 13 15 2 3 1 9
10 3 13 2 7 2 16 15 13 2 13
14 15 13 3 2 9 2 15 15 3 1 15 9 13 13
18 1 15 9 13 1 15 9 9 9 15 15 3 13 2 9 15 3 13
9 15 9 0 9 3 13 9 0 13
8 15 13 9 9 3 13 1 9
17 15 15 9 15 9 9 13 3 7 1 9 9 7 1 9 9 13
18 3 16 9 0 9 0 9 9 13 2 3 3 0 0 9 15 9 13
11 13 9 9 0 15 9 0 9 15 13 13
32 1 15 13 15 3 1 13 9 9 0 2 3 1 0 0 9 7 9 2 7 1 0 9 0 7 1 0 15 9 7 9 13
60 3 13 15 15 9 2 9 2 7 15 9 9 13 0 2 16 13 13 15 9 15 13 15 3 9 0 9 7 9 9 13 1 9 1 9 2 9 9 7 9 9 13 9 13 2 9 7 9 0 3 9 15 7 9 0 7 9 9 0 13
21 3 15 0 9 3 13 16 13 13 3 13 0 15 9 7 2 16 13 2 9 13
13 15 13 2 15 13 2 7 3 3 13 7 13 13
17 3 3 15 13 13 15 9 1 9 2 3 13 9 15 7 13 13
21 15 3 15 1 15 13 9 7 13 13 13 2 16 15 0 13 13 1 9 9 13
7 3 3 15 0 13 15 9
5 13 9 3 1 9
14 15 15 1 15 0 9 2 3 1 0 9 7 9 13
18 16 15 1 9 9 13 9 2 9 13 9 2 16 13 0 9 9 13
5 15 15 9 3 13
23 7 16 15 0 9 9 13 3 3 7 13 13 2 13 15 9 9 16 0 9 9 13 13
28 15 2 16 9 9 9 13 9 9 0 7 3 3 15 13 2 13 15 9 7 9 13 2 15 9 7 9 13
23 16 15 9 13 7 13 0 7 3 15 9 0 13 13 2 16 13 2 1 15 9 3 13
25 3 15 9 2 15 0 13 9 0 15 2 13 7 13 7 3 3 9 15 13 16 1 9 0 13
14 15 15 7 3 9 13 7 3 9 13 7 3 9 13
12 15 15 2 9 2 3 13 7 3 3 13 13
14 0 3 15 9 9 13 16 1 15 2 0 9 1 15
15 15 0 9 9 9 2 15 9 7 9 9 0 13 7 0
15 15 3 3 1 13 9 7 9 3 3 1 13 7 13 13
12 0 15 2 16 13 3 13 2 3 16 13 13
33 3 3 15 0 13 1 9 1 0 15 2 15 13 2 9 13 2 0 13 1 15 9 13 13 15 1 0 9 13 2 3 13 13
9 15 1 9 13 7 15 15 9 13
20 15 16 15 2 16 13 2 9 13 2 3 13 13 2 3 16 9 13 3 13
15 15 2 16 15 15 1 9 13 2 16 13 9 9 1 8
5 9 15 13 13 13
18 1 15 3 13 3 1 15 13 13 13 2 7 16 9 8 15 13 13
18 7 3 3 13 1 9 7 1 9 13 13 15 15 15 3 0 9 13
6 13 2 13 2 1 9
20 15 7 13 7 2 16 15 9 13 15 13 15 13 1 9 2 13 15 13 13
20 3 13 2 15 16 13 1 0 9 2 7 3 13 16 13 15 15 1 15 13
20 13 1 9 2 9 2 13 9 0 9 2 1 9 2 16 15 9 13 2 13
2 15 13
7 15 13 2 15 13 15 9
3 13 2 13
9 15 13 9 13 2 15 9 13 13
28 15 15 3 1 15 3 3 9 7 9 13 2 15 3 13 16 15 15 15 13 3 3 13 13 3 1 9 13
3 7 15 13
7 3 15 15 9 9 0 13
32 7 13 2 16 0 9 13 13 1 9 9 13 2 0 9 9 15 2 16 3 1 0 9 0 9 9 0 2 7 1 9 13
17 7 13 0 2 16 3 0 15 13 13 9 7 1 9 0 9 13
20 7 15 16 9 0 13 2 16 9 9 13 2 16 9 9 0 13 3 13 13
22 3 13 9 9 2 16 15 13 2 3 9 15 9 2 16 1 9 9 9 13 2 13
51 16 7 13 0 9 7 9 13 2 13 1 0 13 9 2 13 15 1 9 2 13 13 9 2 13 15 1 0 2 13 9 9 2 13 0 9 2 16 1 15 3 13 1 9 2 7 13 1 0 13 13
57 7 3 15 15 13 2 1 15 3 13 13 13 15 15 1 9 0 13 13 2 15 13 13 7 13 1 9 9 2 1 15 3 9 15 0 15 15 7 0 0 13 0 7 0 13 2 15 9 0 9 0 13 13 2 13 13 13
14 13 3 3 3 15 3 3 0 15 9 13 7 0 13
13 7 3 3 15 15 9 13 9 2 7 15 0 9
12 1 15 15 9 9 13 2 9 13 2 9 13
12 3 15 3 3 9 7 3 9 3 16 0 13
17 13 13 1 13 7 1 0 3 3 9 7 3 9 13 13 0 9
29 3 15 15 9 13 2 15 9 13 2 0 1 9 13 2 16 1 0 9 9 7 3 13 9 0 15 7 3 13
35 1 15 9 9 13 15 13 15 13 9 0 2 13 9 3 3 1 13 9 7 3 1 9 13 2 13 3 3 13 9 9 7 3 9 0
21 13 16 13 0 15 0 9 9 2 9 2 9 9 0 15 15 0 9 13 13 13
34 0 13 2 16 15 1 9 13 2 16 9 3 13 16 9 13 9 0 13 2 7 16 15 15 13 1 15 3 13 9 3 16 9 13
6 8 2 9 2 15 13
16 3 15 1 9 13 2 3 1 9 13 2 3 0 9 13 13
4 15 3 15 13
12 7 3 3 9 1 15 9 0 0 9 9 13
13 7 3 1 15 9 15 1 9 0 13 9 9 13
4 7 9 9 13
20 7 2 16 9 13 9 2 13 9 2 9 13 2 3 15 3 13 9 9 13
16 15 15 0 9 0 9 7 15 9 15 15 15 13 9 9 13
41 7 16 0 9 7 0 9 9 7 9 7 9 7 0 9 9 3 3 15 3 13 7 7 13 2 3 13 15 3 13 16 15 15 9 9 13 9 15 1 9 13
21 7 16 15 15 3 13 2 3 15 9 13 3 16 9 9 13 9 2 3 9 13
19 7 3 0 13 1 15 9 15 7 15 15 13 3 13 7 15 15 13 13
12 15 9 9 0 9 13 7 9 13 3 13 13
21 15 9 9 3 3 0 7 7 0 2 16 1 15 13 2 3 7 3 13 13 13
31 3 13 2 16 15 2 16 13 2 1 0 9 13 2 9 3 0 13 15 3 13 9 13 13 2 9 3 0 15 3 13
17 15 7 0 13 13 15 9 0 9 3 13 2 3 1 9 13 13
32 7 3 3 2 9 13 2 1 15 9 9 7 9 13 2 7 13 16 9 0 9 7 0 9 7 9 9 1 0 9 9 13
35 3 16 1 0 9 15 0 13 2 13 3 1 0 15 9 9 7 9 13 13 2 9 7 13 7 13 13 3 1 9 7 1 9 9 0
44 16 3 9 0 9 0 2 16 9 7 9 13 2 16 9 0 13 2 3 13 13 2 3 3 3 7 3 13 2 3 15 9 15 13 1 9 0 13 15 9 3 0 9 13
26 15 9 13 0 2 13 15 1 0 2 0 1 9 13 2 9 3 2 16 3 3 13 2 13 1 15
23 13 13 9 0 9 2 13 9 9 0 2 13 1 9 9 2 9 7 9 1 13 9 13
12 13 3 13 1 9 0 15 15 1 9 0 13
34 15 9 2 9 2 1 0 9 0 9 2 1 0 9 7 9 1 15 9 15 15 15 0 9 7 9 13 2 13 1 0 9 7 0
71 15 2 9 2 15 15 15 15 9 9 1 9 13 13 2 15 9 15 9 7 9 3 13 2 15 7 15 9 1 0 7 0 9 2 1 9 9 7 9 2 1 9 7 9 9 0 13 7 9 0 0 2 9 9 2 9 9 9 9 1 15 7 0 9 13 0 9 0 7 0 13
40 3 3 2 9 2 8 2 9 2 13 9 2 9 13 2 9 9 3 13 2 15 7 15 9 9 7 9 13 1 9 7 13 7 13 7 15 13 9 13 13
7 13 2 13 2 13 2 13
13 0 3 9 1 9 15 7 9 9 15 1 9 13
11 7 15 3 0 15 9 0 9 1 9 13
28 3 7 3 1 9 0 9 15 13 2 3 1 9 2 3 1 9 2 3 1 9 2 3 3 1 0 9 13
10 9 15 13 13 2 16 13 1 9 13
9 3 3 1 9 0 13 9 0 13
17 1 9 13 9 7 3 13 2 16 15 1 13 9 1 0 9 13
42 16 3 3 0 9 2 16 13 2 13 2 16 0 15 13 13 2 16 15 9 1 9 13 2 16 0 9 2 16 13 9 13 2 0 3 15 9 13 13 7 13 13
29 13 15 3 13 2 9 2 7 15 13 7 13 13 13 7 13 9 3 3 1 15 9 15 1 0 9 13 13 13
13 15 3 15 13 13 2 16 0 9 13 7 3 13
45 7 16 15 13 0 0 13 9 13 2 15 1 15 15 1 15 13 7 13 9 0 15 3 13 2 16 3 0 9 3 13 3 16 13 2 3 13 15 0 9 2 9 2 7 9
28 13 13 8 2 9 7 0 9 13 3 3 13 2 7 15 1 15 7 9 9 7 15 9 9 7 9 0 13
32 7 3 0 13 13 15 15 15 13 3 13 2 3 0 15 1 9 3 13 2 3 0 15 3 13 2 3 0 15 1 9 13
26 7 16 15 13 13 1 15 0 9 13 2 3 3 15 8 2 9 3 3 9 0 7 7 9 9 13
44 7 16 13 2 3 15 3 0 3 3 9 13 16 15 2 16 13 13 2 9 13 2 13 16 15 9 9 13 13 3 13 2 9 3 13 16 3 3 13 13 16 9 3 13
29 15 3 15 9 2 9 2 3 3 3 13 13 13 2 7 3 13 2 16 3 15 3 13 16 1 9 3 13 13
7 3 15 0 15 0 9 13
24 9 15 13 15 13 1 9 13 2 9 7 9 15 9 0 13 1 9 0 9 0 9 13 13
13 13 15 9 2 0 9 0 2 3 13 2 3 0
56 3 15 15 9 1 0 9 7 15 9 15 1 9 0 7 0 8 2 9 13 2 7 15 9 15 1 15 3 13 2 0 9 13 2 13 1 9 13 2 1 0 9 2 1 0 9 2 1 15 15 9 13 16 15 9 13
17 15 15 3 3 16 9 9 0 2 7 3 16 9 9 13 2 13
31 15 15 13 13 1 9 2 15 13 1 9 2 15 3 1 9 13 2 15 13 9 2 15 13 9 2 13 15 0 9 13
18 15 16 3 13 2 13 3 3 9 15 13 15 16 15 15 9 13 13
16 7 15 3 13 13 3 16 15 13 15 13 13 7 3 3 13
26 13 15 13 9 13 2 15 13 9 2 15 9 0 2 15 0 2 15 15 15 0 9 9 7 9 13
9 0 0 9 9 1 15 13 13 13
5 13 1 9 0 9
5 9 15 13 2 13
3 15 15 13
13 6 15 3 13 2 16 15 0 0 9 0 13 13
17 15 13 2 3 13 13 16 15 0 13 13 3 9 1 9 0 13
13 7 3 7 15 13 15 9 0 1 9 13 3 13
5 3 13 3 9 9
4 9 9 15 13
4 0 3 3 13
11 13 2 13 2 6 13 9 15 9 0 13
2 13 9
4 0 9 13 13
7 16 13 13 2 1 9 13
13 15 3 9 7 9 13 7 13 13 15 3 15 13
56 15 0 9 9 2 15 9 2 15 9 2 15 9 2 15 9 2 15 9 9 2 15 9 2 15 9 2 15 9 2 15 9 2 15 9 0 2 15 9 9 2 15 13 2 15 13 13 13 15 15 1 9 3 3 13 13
16 15 9 1 15 9 1 15 13 13 2 15 0 9 3 1 15
13 3 3 15 0 3 1 0 9 9 13 0 1 15
25 15 0 15 13 3 2 9 9 3 13 2 0 9 9 2 0 9 9 3 3 13 7 3 13 13
17 3 3 3 3 3 3 1 9 7 3 1 9 0 9 13 9 13
24 9 3 3 9 7 3 0 3 1 9 0 9 13 9 0 13 15 3 1 15 0 9 9 13
42 7 16 15 13 9 1 0 9 13 13 2 9 13 1 9 0 0 1 9 0 15 15 3 9 9 13 13 2 9 1 9 0 7 0 15 15 3 15 3 9 13 13
32 7 15 3 9 7 9 9 13 9 7 9 7 9 7 9 13 0 1 15 13 2 16 9 9 7 9 9 1 9 7 9 13
13 3 3 3 13 0 9 9 2 3 0 7 13 9
10 15 13 16 9 2 16 9 2 16 9
7 9 0 13 2 9 0 13
9 9 15 3 3 2 9 3 13 13
9 15 3 15 15 13 1 9 9 13
21 7 16 1 9 7 9 9 3 7 9 13 2 13 15 3 13 2 7 3 13 13
32 15 15 13 1 9 2 13 9 0 2 9 0 2 13 9 2 9 13 2 9 13 2 13 9 13 9 0 9 0 7 9 9
25 15 15 13 13 9 15 7 9 3 3 9 2 9 2 9 2 9 13 7 13 3 3 7 3 13
23 15 16 0 9 2 16 13 3 13 2 13 2 3 0 13 15 9 7 0 9 13 9 0
15 0 7 13 9 15 13 2 0 9 15 9 9 0 13 13
9 0 13 0 0 9 9 7 9 13
16 0 9 13 2 3 9 13 2 3 13 9 13 2 3 13 9
11 1 9 15 2 1 9 2 1 9 13 13
8 15 15 15 9 9 13 2 9
4 13 9 9 13
16 15 13 13 15 9 13 2 15 13 13 3 13 1 9 9 13
21 3 7 13 7 13 7 2 16 7 1 9 7 1 15 9 13 2 15 15 13 13
13 7 3 13 15 13 2 9 2 1 15 13 13 9
13 7 15 16 9 13 13 2 15 15 13 15 15 13
12 9 7 3 0 7 3 0 9 9 13 3 13
9 3 7 13 1 9 13 13 2 13
24 7 0 9 2 16 9 9 3 13 13 2 9 1 9 9 9 13 2 9 0 1 9 13 13
26 3 16 9 13 2 15 15 9 13 2 15 13 2 15 3 3 13 16 13 9 7 3 3 16 0 9
16 7 3 9 15 9 9 15 9 1 15 15 13 0 7 0 13
23 3 15 0 15 9 15 9 9 1 9 13 13 1 9 1 0 9 1 9 2 9 13 3
11 16 15 9 0 9 13 3 13 2 13 9
23 15 15 9 13 2 7 13 2 15 1 0 13 2 15 1 9 13 15 9 0 9 13 13
10 1 9 13 15 3 13 13 1 9 13
11 6 9 0 3 3 13 7 3 13 9 0
78 3 16 8 2 9 9 2 9 2 9 0 13 7 13 3 13 2 9 13 2 13 0 2 9 9 13 13 2 7 1 15 9 9 7 9 9 1 9 7 1 9 13 2 3 15 1 15 13 9 9 2 3 13 7 13 0 9 2 3 1 9 7 9 13 2 7 0 0 1 9 13 1 9 9 7 9 13 13
23 7 13 15 15 2 16 15 13 2 3 0 7 0 2 15 3 0 9 7 0 9 13 13
25 13 15 3 2 9 2 15 9 0 7 0 9 13 2 16 3 1 15 15 0 9 7 0 9 13
12 13 3 13 13 1 15 2 16 3 13 1 9
7 7 15 13 2 3 13 13
30 3 15 1 9 0 13 2 9 2 9 0 13 9 16 8 2 9 13 9 9 7 1 9 13 13 2 7 9 3 13
17 7 0 3 15 13 16 15 13 0 3 16 15 13 3 16 16 13
23 7 16 13 9 15 15 2 16 13 13 2 13 13 13 2 15 2 16 13 13 2 15 13
13 7 15 15 9 9 13 13 3 3 15 13 16 13
15 9 13 15 3 0 15 15 3 1 9 16 1 9 13 13
30 3 3 2 16 15 15 3 1 15 9 7 9 13 2 16 7 0 15 9 13 13 2 13 3 16 13 1 9 16 13
14 1 15 15 13 2 15 9 13 2 15 15 13 15 13
39 15 3 15 2 16 0 9 13 13 2 3 3 13 13 16 13 15 15 2 13 9 0 2 7 3 15 15 9 13 3 13 2 16 3 15 13 13 2 13
13 13 3 15 2 9 2 1 15 9 9 15 9 13
13 3 0 9 9 7 9 0 2 16 3 13 2 13
20 0 9 13 15 15 0 1 9 0 0 3 9 13 15 9 13 13 0 9 13
15 15 9 9 13 0 2 13 16 0 2 9 3 7 9 0
9 0 9 13 3 0 7 0 7 0
48 15 3 3 13 2 15 3 13 2 15 3 9 2 3 3 13 9 2 3 3 9 1 0 9 0 13 2 15 9 2 9 2 9 9 13 0 7 1 9 7 1 9 15 1 15 9 13 13
11 15 15 3 3 9 0 16 9 0 13 13
24 15 9 3 3 2 16 13 3 13 2 13 2 7 3 16 3 3 9 7 3 9 3 0 13
10 0 9 13 9 2 9 2 3 9 0
6 15 15 1 9 3 13
23 7 7 3 1 15 13 13 7 13 3 1 9 2 16 13 3 0 16 15 9 13 3 13
29 0 7 9 13 3 3 9 7 3 9 15 7 9 15 0 9 13 2 1 15 9 2 3 3 1 9 15 7 9
23 15 0 9 2 0 2 7 0 7 3 0 13 2 0 7 0 9 2 9 13 2 3 9
11 15 0 9 9 7 13 9 1 0 9 13
14 1 15 9 0 9 2 0 9 2 0 0 7 0 13
24 15 9 3 0 7 0 3 3 13 7 13 7 3 13 7 13 7 7 9 13 7 13 9 13
20 15 16 13 2 16 13 2 3 16 9 13 2 13 15 1 9 0 9 9 13
7 7 3 15 15 15 0 13
8 3 0 15 9 13 1 9 13
12 15 1 9 7 15 13 13 2 15 3 3 9
11 15 7 9 15 9 7 15 9 7 9 13
16 13 3 2 9 2 1 15 3 0 9 9 0 9 7 0 9
12 7 3 9 15 13 7 0 9 7 9 0 13
14 3 1 15 9 13 7 13 9 9 0 9 7 9 13
10 3 7 9 9 7 9 13 9 9 0
18 7 3 15 0 9 2 9 2 9 0 1 15 9 9 7 9 13 13
12 9 0 0 0 15 13 9 2 13 0 3 9
25 3 15 0 13 9 9 7 9 13 13 9 9 2 16 15 13 0 13 9 0 2 7 0 13 9
16 7 15 3 0 9 15 3 13 9 2 16 3 0 13 13 9
11 9 0 13 2 9 2 9 9 0 13 9
10 15 3 0 13 9 9 0 0 9 13
5 3 0 13 13 9
8 3 1 9 9 7 3 9 13
19 1 15 0 9 3 0 13 9 2 7 7 13 0 2 16 3 2 13 9
30 7 15 2 13 15 13 9 9 7 9 1 0 0 13 9 2 6 6 9 9 13 0 2 7 13 15 9 13 9 3
12 3 15 13 15 7 9 7 9 13 0 13 9
15 3 7 9 0 13 7 9 2 13 3 9 15 13 9 13
16 13 1 0 9 7 13 1 9 2 3 3 0 0 9 13 9
16 15 13 2 15 0 9 13 9 2 13 7 1 0 3 9 0
21 1 15 0 9 9 13 0 2 7 0 0 9 13 9 2 15 2 13 2 13 9
11 0 15 13 9 2 7 3 0 13 9 9
43 3 13 13 13 2 9 2 9 7 0 0 9 13 9 2 7 3 0 9 13 9 2 7 15 0 13 9 2 7 9 9 13 13 9 2 7 7 13 1 0 9 13 9
9 13 15 2 3 0 0 13 9 9
6 0 9 9 3 13 9
28 13 15 13 9 0 9 2 3 13 9 9 0 3 2 13 7 1 0 3 9 9 2 7 13 0 13 9 9
12 9 0 13 13 9 2 7 9 0 3 9 13
11 7 7 0 0 13 9 9 13 0 9 9
13 7 9 13 0 0 9 2 0 0 13 9 1 9
9 3 15 3 13 16 13 15 0 15
9 0 16 9 13 2 0 9 3 13
28 16 15 3 9 0 9 13 7 0 0 9 9 2 0 7 7 13 0 9 9 2 0 15 9 2 15 9 13
14 15 15 3 13 0 0 9 2 9 16 0 13 15 9
11 3 7 13 0 0 9 0 3 0 9 9
26 0 13 15 0 13 9 9 3 0 13 9 9 2 0 16 0 13 9 9 2 7 13 0 9 9 9
14 15 15 2 3 3 9 13 0 2 3 13 13 13 9
40 7 3 0 13 9 13 3 9 3 9 2 0 0 9 2 13 3 13 13 9 7 9 13 13 7 9 9 2 3 3 13 13 9 13 9 2 13 13 9 9
14 7 3 13 0 1 9 9 7 13 0 2 9 2 9
6 7 3 13 13 13 9
6 3 0 0 9 13 9
7 3 13 1 0 13 9 9
11 3 15 0 13 9 9 0 13 13 1 0
15 6 3 0 13 2 0 2 9 2 15 0 0 3 13 13
11 3 3 15 13 13 0 0 3 1 9 9
6 15 13 9 0 9 0
12 3 15 3 13 9 15 13 15 3 13 13 9
19 15 13 9 9 9 2 7 15 0 13 9 9 2 7 15 13 0 9 9
6 9 3 15 9 13 13
8 15 7 9 0 9 13 0 9
9 13 0 2 15 2 9 2 13 13
14 15 3 7 0 13 13 9 2 15 3 13 13 0 9
3 3 3 13
11 13 15 0 9 7 15 3 0 9 9 13
12 7 7 15 15 1 15 13 9 7 7 15 13
14 13 0 9 15 0 2 7 15 1 0 0 13 9 13
5 6 0 9 0 13
13 3 0 3 13 9 9 3 15 16 13 13 9 9
14 13 3 3 2 13 2 7 7 15 1 15 15 13 13
5 15 15 13 2 0
21 0 2 13 0 13 9 2 7 0 0 9 13 1 9 2 7 13 1 0 9 9
7 3 13 15 0 0 13 9
6 3 13 3 13 15 15
15 7 16 9 0 3 13 0 9 2 7 15 9 12 0 13
9 3 15 3 9 2 3 15 13 9
6 15 0 9 13 0 9
50 6 2 0 13 3 1 9 13 2 16 15 9 0 9 13 2 7 0 0 13 9 9 2 7 9 0 13 1 9 9 2 7 15 13 13 15 9 13 2 7 7 13 2 15 13 7 3 2 13 0
13 3 0 9 0 13 9 13 7 13 15 13 13 9
15 7 7 3 9 3 13 0 2 7 3 13 0 9 0 15
7 7 7 15 9 13 13 9
5 13 9 0 13 9
15 3 15 3 13 9 13 13 2 16 15 0 0 13 9 9
12 7 3 0 0 13 9 0 1 0 0 13 9
5 3 3 15 13 13
28 3 15 3 9 13 9 13 15 2 9 2 8 7 0 13 9 9 2 7 15 0 13 13 9 7 9 13 0
13 7 15 13 13 9 9 2 7 13 0 3 9 9
13 15 15 0 13 9 9 2 7 13 0 13 13 9
7 15 15 3 9 13 13 9
8 6 13 2 16 15 0 13 13
13 15 9 0 13 13 9 2 7 0 13 9 13 9
14 7 15 3 3 0 9 15 9 13 7 9 0 0 0
14 15 13 2 15 3 13 9 13 2 15 9 0 13 9
14 9 0 13 1 9 3 2 1 15 9 15 3 9 13
9 3 15 13 9 2 3 13 0 9
6 15 15 9 9 13 13
15 7 15 7 0 3 13 9 2 7 3 0 9 13 9 9
14 7 9 9 7 9 13 9 13 2 7 13 9 13 9
16 3 15 16 15 15 13 3 0 9 2 13 15 0 9 0 13
13 7 7 3 9 3 13 9 13 7 9 9 0 13
17 15 15 13 9 9 2 15 0 9 13 2 3 13 9 9 13 0
28 15 13 13 9 13 9 2 9 2 7 0 3 13 9 15 13 3 1 15 13 9 2 7 13 15 13 0 9
14 7 3 13 9 0 13 9 2 9 0 0 9 2 13
7 15 13 0 0 13 9 9
6 3 13 0 9 0 9
20 3 13 13 15 9 9 7 0 9 9 13 9 2 3 3 1 0 13 13 9
6 0 1 0 9 9 13
12 7 16 3 13 13 13 15 2 13 13 9 9
16 3 3 0 13 13 9 2 13 15 1 15 0 2 9 2 9
13 13 15 13 3 13 9 2 7 9 0 13 13 9
15 7 13 0 9 13 0 2 7 7 0 1 9 13 9 0
9 9 15 13 3 15 13 15 13 13
17 7 2 16 15 13 2 0 9 13 2 7 15 1 9 9 0 13
14 13 13 2 16 13 15 2 7 3 13 0 13 13 9
15 7 15 13 0 3 7 9 9 2 15 3 9 3 13 0
13 15 13 0 0 13 9 2 15 3 0 9 9 13
6 15 1 0 13 9 9
14 7 15 13 15 13 9 9 13 1 0 2 9 2 9
37 7 3 3 15 9 13 9 0 0 9 13 9 2 7 13 13 0 9 1 9 0 0 13 9 9 2 16 13 0 0 13 9 3 1 0 9 13
10 13 3 2 16 15 15 0 9 13 0
3 9 9 13
8 7 1 15 9 9 13 0 0
16 7 0 13 7 1 0 9 2 15 13 2 13 2 9 9 13
7 15 3 3 3 0 13 9
16 3 15 9 3 13 13 9 2 15 13 15 2 0 9 2 9
14 3 0 15 0 13 13 9 9 2 3 9 0 13 9
16 7 3 15 13 9 13 9 9 2 7 3 0 3 1 9 13
3 3 0 13
10 3 15 9 15 13 16 0 13 13 9
2 9 13
4 3 15 9 13
7 7 15 13 0 13 9 9
5 3 13 15 15 13
4 13 9 0 9
6 0 1 0 9 13 9
13 3 3 0 0 13 9 13 7 15 0 9 13 0
6 3 3 13 13 9 9
12 7 16 13 13 13 9 2 13 3 13 9 9
11 15 7 3 13 0 7 3 15 13 9 13
7 9 0 13 2 9 9 13
17 15 2 16 3 13 2 0 13 9 2 9 2 16 13 0 9 13
9 7 3 15 0 13 2 0 2 9
8 13 15 3 2 9 2 9 13
28 16 15 13 13 9 9 2 0 7 1 0 13 9 9 2 13 1 15 0 13 9 13 2 7 0 13 13 9
6 15 13 15 13 9 9
5 0 0 13 0 9
14 15 15 0 15 13 9 2 7 7 0 13 3 0 13
9 15 15 3 9 0 2 3 9 13
2 13 15
5 15 13 9 13 13
32 13 15 15 0 13 13 9 7 13 13 2 9 2 3 9 2 7 13 13 9 13 9 2 7 15 3 0 13 2 9 2 9
6 3 15 9 13 13 0
6 0 13 0 1 0 9
26 3 3 0 9 13 9 0 0 13 9 9 2 7 7 3 0 13 9 9 9 13 1 0 9 0 9
6 0 9 0 13 13 9
4 15 0 9 13
18 7 3 0 2 7 13 9 0 7 0 9 7 9 9 0 2 0 12
13 15 13 9 7 0 9 2 15 0 9 13 13 9
9 15 3 16 3 13 13 9 2 13
5 3 0 9 0 13
9 15 15 13 0 2 16 0 13 9
8 7 15 13 2 0 13 15 15
26 15 13 13 0 3 9 0 0 9 13 9 2 7 3 3 0 13 13 9 7 3 3 0 9 13 9
12 7 9 0 13 13 9 9 2 13 0 9 9
7 3 3 15 0 13 13 9
5 13 9 0 13 9
7 3 15 13 13 0 9 9
8 15 13 2 16 15 9 13 13
6 0 15 0 9 13 9
13 15 13 0 9 13 9 2 15 3 0 9 13 9
23 15 7 3 0 13 13 9 7 3 13 0 2 9 2 13 9 2 7 0 0 9 13 9
5 15 13 0 9 0
14 15 15 16 13 13 2 3 0 13 9 7 9 9 13
15 3 15 0 0 9 0 13 2 15 3 13 2 9 2 9
6 13 15 0 13 9 9
7 15 3 1 0 0 9 13
11 7 3 3 0 8 13 9 0 3 13 9
39 0 15 9 0 0 9 13 2 0 0 13 9 2 7 16 3 1 15 13 2 13 15 3 2 0 0 9 7 7 3 9 13 0 9 9 0 13 1 9
12 9 0 1 15 13 9 2 16 3 0 13 9
14 9 0 13 13 1 9 9 2 9 7 0 9 13 9
13 15 0 0 13 13 9 2 15 3 16 13 0 9
14 13 3 13 0 9 9 2 9 2 7 13 13 13 9
14 0 6 3 2 0 13 9 2 16 15 9 15 0 13
21 0 3 0 13 9 9 2 9 7 13 13 3 9 2 16 0 1 0 13 9 9
7 13 15 13 2 3 0 3
15 3 15 3 0 15 13 9 2 1 15 3 15 13 9 13
14 15 15 13 2 16 15 13 13 2 16 15 13 13 9
14 7 1 0 13 15 13 9 2 7 3 13 13 0 9
10 15 0 13 9 9 2 9 9 0 0
27 3 15 2 0 9 0 9 2 13 0 3 13 9 2 7 15 3 13 0 13 9 3 7 13 9 13 9
12 7 7 13 0 9 13 9 2 0 0 13 9
15 2 7 3 3 15 9 13 13 9 2 0 7 9 13 9
11 15 0 3 13 13 9 2 0 13 9 9
14 9 3 9 3 0 15 2 3 15 3 0 13 13 9
12 3 3 13 0 13 9 2 0 0 13 13 9
15 3 0 9 13 0 13 9 2 0 7 1 0 9 9 13
16 15 0 9 2 15 9 0 13 2 7 0 0 15 13 9 9
10 15 0 0 3 13 9 13 13 0 9
12 6 3 13 0 0 9 9 13 9 13 1 9
30 13 16 3 9 13 15 0 2 13 16 7 9 0 7 9 2 3 3 15 0 13 13 9 2 13 7 0 9 1 9
13 3 13 0 0 13 9 2 7 0 0 9 13 9
16 7 15 0 0 15 0 9 9 2 13 0 3 2 9 2 9
25 15 3 0 0 13 9 9 2 15 13 13 13 0 9 16 15 3 0 0 13 9 0 9 13 9
14 7 15 3 0 13 9 9 2 7 9 13 13 13 9
16 1 0 3 13 15 2 0 2 9 2 7 13 13 9 13 9
13 15 15 3 16 15 0 13 9 2 7 0 13 9
12 3 15 3 9 9 7 3 9 9 0 13 9
7 7 13 2 16 13 13 9
5 3 15 0 13 9
14 7 3 15 9 0 13 9 2 7 0 0 9 9 13
9 7 3 13 13 15 2 9 2 9
7 13 2 3 0 13 9 9
6 3 0 13 13 9 9
6 15 0 0 9 9 13
15 7 13 0 0 9 13 9 2 7 9 0 0 0 13 9
14 6 13 2 15 9 7 9 13 0 7 0 9 13 9
28 3 16 15 0 13 9 9 2 0 7 13 13 9 9 2 15 0 0 13 9 9 2 3 7 0 13 9 9
14 15 9 0 13 9 9 2 3 15 3 0 9 9 13
12 16 3 0 13 9 13 9 2 0 9 13 9
14 15 3 13 9 7 0 13 2 7 0 9 13 9 9
13 3 13 13 13 3 9 16 3 0 13 9 13 9
9 3 0 3 13 2 0 9 2 9
8 15 15 13 13 2 9 2 9
13 15 3 0 1 13 9 3 1 9 0 13 13 9
3 3 0 13
5 15 15 15 9 13
6 7 0 9 9 9 0
16 3 15 15 13 2 0 2 16 3 0 0 9 0 13 0 9
32 3 0 15 9 15 0 9 13 2 3 3 0 3 13 9 0 2 16 15 13 3 3 9 2 7 0 13 9 13 0 13 9
16 7 7 0 13 13 9 9 2 7 3 0 0 13 1 9 9
14 6 3 0 13 0 9 1 9 2 13 7 0 9 9
7 7 0 7 13 15 9 9
6 15 3 13 13 13 9
12 0 13 0 13 0 9 7 3 0 9 9 13
13 1 15 0 9 7 0 9 7 13 0 9 0 9
13 7 15 0 13 13 9 2 13 1 13 13 0 9
17 7 3 13 13 15 2 9 2 9 2 7 7 0 0 9 9 13
18 3 15 3 0 13 2 0 9 2 9 2 7 7 13 0 13 9 9
15 7 16 9 0 13 15 9 9 2 15 9 13 15 0 9
14 3 3 3 0 9 13 9 2 16 0 13 9 9 13
23 3 9 0 9 9 3 13 0 0 13 9 2 7 0 0 13 9 9 0 0 13 9 9
8 3 15 13 2 3 0 13 9
6 13 3 9 9 9 9
12 3 0 13 9 9 2 15 13 0 0 9 9
25 15 0 0 13 15 2 9 2 9 0 2 3 2 9 15 3 0 13 2 16 15 0 13 9 9
6 0 3 9 9 13 0
7 15 15 0 0 13 13 9
8 3 15 3 0 9 13 0 9
23 3 13 2 16 15 13 2 9 2 9 13 1 0 9 0 9 2 13 7 0 9 13 13
5 13 0 0 9 9
9 6 2 16 13 2 1 15 13 13
7 3 3 13 0 9 0 9
4 0 9 13 9
14 13 15 3 1 9 2 3 9 0 2 0 0 9 9
17 3 15 13 0 9 7 0 9 2 9 2 7 3 13 3 13 9
11 15 0 0 9 13 1 9 9 0 13 9
14 3 9 9 2 0 16 13 9 2 0 0 9 9 13
11 7 9 0 9 13 3 0 13 13 9 9
11 15 1 0 13 13 9 7 0 9 13 9
5 3 0 13 9 9
5 13 9 2 13 9
21 15 3 13 0 3 9 13 9 13 9 2 7 3 0 13 0 9 9 0 13 9
11 3 13 13 13 9 9 13 0 0 13 9
16 15 16 13 9 9 9 13 13 13 9 2 13 3 0 13 9
6 3 9 13 9 13 9
14 15 3 9 13 9 2 7 15 9 1 0 9 9 13
15 15 2 6 9 2 0 13 13 9 2 0 9 13 13 9
6 9 15 13 0 0 9
15 3 15 13 16 13 13 9 2 7 9 9 0 13 1 9
13 7 15 1 13 13 9 9 0 2 15 13 13 0
6 7 15 13 0 0 9
27 7 15 3 13 0 13 9 2 16 15 13 13 9 9 2 16 15 13 0 13 1 9 0 0 3 13 9
18 7 15 3 0 2 15 13 2 15 13 2 16 1 15 9 3 13 13
15 15 9 0 13 13 9 2 15 13 0 2 9 2 13 9
28 6 3 0 13 9 9 2 7 13 0 0 9 9 2 7 7 15 0 13 9 9 2 7 0 0 13 9 9
16 7 15 9 1 15 2 0 2 13 2 13 9 0 3 0 9
16 7 7 15 13 9 13 13 2 13 2 15 9 13 9 0 13
11 6 15 3 0 2 7 3 15 0 9 13
15 6 15 13 13 0 9 9 0 2 7 1 0 9 13 13
2 3 13
3 3 13 13
2 13 9
1 13
5 0 3 13 15 9
6 0 13 0 13 9 9
6 13 13 0 9 0 9
16 15 0 15 7 1 15 0 9 13 2 7 1 15 0 9 13
15 3 0 13 2 3 0 13 2 3 3 15 0 13 0 9
15 15 15 3 9 2 3 0 13 9 2 7 13 0 9 9
14 13 7 9 2 7 7 9 0 9 2 15 15 0 13
4 9 0 0 13
7 3 15 0 13 13 9 9
9 16 9 7 9 13 2 15 0 13
7 7 7 15 9 0 13 9
5 15 0 13 9 9
15 13 15 13 2 9 2 9 2 7 7 15 3 0 9 13
16 6 13 7 9 13 1 9 9 2 7 15 3 15 13 13 9
14 3 15 0 13 1 9 9 13 2 15 9 15 9 13
7 15 9 7 9 3 13 0
13 3 15 3 0 13 0 13 9 7 0 9 13 9
7 3 1 9 13 9 9 9
7 3 15 0 0 9 13 9
6 15 13 13 0 9 9
25 3 3 0 13 13 9 7 3 0 9 13 9 2 16 9 3 9 13 9 7 9 13 13 13 0
14 0 9 15 0 3 13 9 2 16 3 0 13 15 9
10 7 3 15 13 2 16 13 3 15 13
10 3 2 16 9 13 2 3 3 9 13
7 13 3 13 3 1 9 13
29 0 9 2 15 15 13 13 0 9 2 0 9 13 13 2 16 9 9 13 3 9 2 15 9 0 7 9 13 13
10 7 0 0 9 1 9 7 9 13 13
7 9 9 2 9 9 3 13
17 7 3 0 1 0 9 13 2 9 9 7 9 9 9 0 3 13
7 7 3 9 9 1 9 13
43 3 3 3 1 9 9 2 1 9 9 7 9 13 9 7 9 13 2 9 13 9 0 13 2 0 9 1 0 9 13 2 3 3 9 7 9 13 13 1 9 0 9 13
11 7 9 3 0 9 13 2 15 9 13 13
20 0 16 1 9 9 2 1 9 7 9 9 7 9 13 2 9 3 1 9 13
10 3 9 3 1 0 15 1 3 0 13
9 15 9 13 13 13 2 9 9 13
16 7 0 9 2 13 9 7 9 2 13 7 13 9 3 9 13
10 15 3 1 9 9 9 2 9 9 13
12 15 15 9 7 9 3 13 2 3 1 0 13
23 0 7 9 15 3 15 13 7 13 9 13 2 15 15 9 13 0 9 7 9 0 9 13
10 7 1 0 9 9 0 0 9 9 13
13 0 13 3 13 9 0 2 3 3 13 3 0 13
7 7 9 7 9 0 13 13
11 7 15 13 7 15 9 0 13 2 0 13
22 7 15 3 2 16 8 0 9 13 9 7 9 9 2 3 1 0 0 13 9 13 13
17 15 16 9 13 13 0 9 2 3 1 0 9 0 9 9 13 13
21 7 15 2 16 1 0 0 9 13 2 3 0 9 9 0 3 0 9 7 9 13
9 7 1 9 9 3 3 13 0 13
12 7 15 9 1 9 15 0 13 9 7 9 9
13 1 15 9 9 0 3 13 13 2 3 9 13 13
20 8 2 9 2 0 9 13 2 13 0 9 7 9 7 9 7 9 0 7 0
17 15 1 9 9 0 9 9 9 9 0 13 2 7 3 9 0 13
8 0 9 0 0 3 0 3 13
24 13 3 7 3 1 9 9 0 9 9 0 7 9 9 2 15 0 15 9 13 2 15 3 13
45 9 15 13 13 2 16 1 9 9 9 13 2 3 13 7 9 13 0 9 7 9 2 15 9 9 0 13 7 0 13 2 16 3 13 1 0 7 0 0 7 0 13 13 2 13
24 15 16 1 0 9 13 2 0 9 2 0 9 2 0 0 9 13 2 0 9 13 3 0 13
10 3 3 9 13 7 0 9 9 13 13
25 7 16 9 15 9 9 9 13 3 0 7 3 13 13 2 16 0 9 13 2 9 1 9 13 13
13 3 9 7 9 0 9 13 2 0 1 9 9 13
7 7 0 9 13 1 9 13
24 7 9 9 7 9 13 13 2 13 2 0 0 13 2 9 3 13 2 9 9 7 9 9 13
20 3 16 9 9 13 2 9 7 9 9 13 2 7 3 13 15 13 9 9 13
7 9 0 2 9 9 0 13
15 13 2 15 9 9 0 2 9 9 0 13 2 9 0 13
8 15 3 9 3 9 9 9 13
30 3 16 0 9 15 9 13 9 7 13 9 0 13 2 1 9 7 9 15 13 2 13 9 0 9 7 0 9 15 13
10 15 9 3 13 13 1 9 13 9 0
14 7 15 9 13 15 15 3 13 7 3 9 1 9 13
15 7 9 0 16 0 0 13 2 7 3 15 0 9 0 13
10 7 9 0 9 13 13 9 0 0 13
4 0 9 9 13
33 3 0 9 2 3 7 9 13 13 2 1 9 1 9 9 9 13 2 7 3 1 0 9 7 0 9 15 1 9 7 9 9 13
19 3 0 9 3 9 0 2 3 9 0 0 7 0 13 2 3 9 9 0
3 9 0 13
7 7 9 0 9 1 15 13
16 15 15 9 13 2 9 13 2 13 2 16 0 9 13 2 13
10 15 9 2 15 0 9 7 0 9 13
6 9 0 2 9 0 13
6 9 0 2 9 0 13
30 13 13 2 15 1 9 0 9 9 9 0 0 9 13 2 15 9 9 13 13 13 2 3 15 9 3 15 1 9 13
7 7 3 9 1 0 9 13
12 15 9 0 1 9 3 3 1 9 13 7 13
16 7 16 13 3 9 0 9 2 1 9 9 9 9 1 0 13
15 3 15 15 13 9 0 13 2 3 15 9 13 13 0 9
38 7 9 0 3 15 9 13 2 16 0 15 3 0 13 2 9 9 1 9 13 2 0 15 13 16 13 2 0 1 0 3 13 13 16 15 0 13 13
7 7 9 7 9 0 9 13
6 9 0 2 0 9 13
11 9 7 9 1 15 3 9 3 16 9 13
12 1 9 9 0 2 9 13 2 1 9 0 13
6 15 3 9 0 0 13
13 1 15 9 2 9 2 9 13 2 0 0 13 13
7 15 3 3 13 2 3 13
19 3 16 9 3 9 13 2 9 13 2 9 1 0 7 0 0 7 13 13
16 7 3 3 9 16 9 9 9 13 2 15 3 9 1 9 13
16 7 15 0 9 13 2 15 16 0 9 13 2 9 7 9 13
9 9 9 9 13 2 15 9 0 13
24 15 7 9 0 13 9 7 9 0 13 2 3 0 7 0 13 2 7 3 9 7 3 9 13
26 3 13 16 9 2 9 9 2 15 1 9 13 2 15 15 0 13 2 1 9 9 3 7 3 3 13
13 7 0 9 2 16 9 13 13 2 9 9 13 13
6 3 0 9 9 9 13
24 16 9 9 13 13 7 15 9 9 9 13 2 13 9 2 9 9 13 2 9 1 9 13 13
10 7 1 9 9 9 7 9 1 9 13
19 7 15 9 9 9 2 9 0 9 13 2 7 7 13 15 1 9 9 13
9 3 3 9 13 15 3 13 9 13
23 7 15 15 13 2 15 16 15 15 13 9 0 13 2 1 13 9 13 9 2 9 13 13
6 15 15 13 9 13 9
10 7 15 3 13 13 2 13 1 9 13
9 9 0 13 2 9 9 1 9 13
7 13 9 9 7 9 9 13
6 13 3 3 9 9 13
18 3 9 7 9 2 7 3 9 7 3 9 13 2 7 15 9 9 13
11 15 9 2 3 0 9 13 2 1 9 13
8 9 13 0 9 3 3 9 13
9 7 3 0 9 9 7 9 13 13
5 7 3 9 9 13
10 15 9 0 7 9 13 9 3 3 13
17 3 7 3 9 7 3 9 0 13 2 16 15 0 7 0 15 13
18 13 13 9 2 15 3 13 9 2 15 9 9 13 2 3 3 9 13
14 7 1 0 9 3 16 15 15 15 13 13 15 9 13
24 3 3 9 9 0 0 9 13 2 1 9 0 2 1 9 9 2 0 15 9 1 9 7 9
34 3 13 9 0 9 2 15 1 9 3 3 0 13 2 16 15 13 15 13 13 9 13 9 2 1 0 13 13 9 0 9 0 9 13
11 15 3 9 15 1 9 13 9 13 9 13
5 3 9 9 13 13
7 3 1 9 7 9 9 13
16 7 9 2 15 2 16 3 13 2 13 2 0 9 0 9 13
7 1 15 9 7 9 0 13
11 3 16 15 9 7 9 8 2 0 0 13
15 3 16 1 9 13 9 7 9 2 0 3 0 7 0 13
41 15 9 7 9 13 9 2 3 16 9 0 1 0 9 0 13 7 16 7 0 0 9 2 3 0 13 2 9 7 9 0 0 0 9 13 2 13 9 0 9 13
13 1 9 0 9 2 8 2 9 1 0 9 9 13
11 9 0 2 0 9 0 2 0 9 9 13
19 16 3 13 13 15 13 2 1 0 9 13 2 15 0 9 7 9 9 13
20 13 3 0 9 3 9 15 9 0 2 15 3 9 9 13 16 9 7 0 9
10 15 1 9 7 3 7 3 13 9 13
8 0 1 0 2 9 16 9 13
15 13 3 15 9 15 13 8 2 0 9 3 0 15 9 13
33 16 8 2 9 2 0 15 2 0 9 13 2 15 9 13 1 15 9 13 2 3 13 2 16 9 13 2 3 1 15 9 15 13
13 7 3 3 13 9 1 9 0 2 1 15 9 13
6 1 15 16 3 13 9
16 0 9 8 2 9 7 8 2 9 13 9 9 9 13 9 13
17 3 9 9 9 13 9 13 13 9 13 2 16 1 0 9 13 13
36 1 15 9 7 9 1 9 9 9 13 13 1 9 9 0 8 2 9 7 8 2 9 9 13 2 15 9 13 9 1 9 1 13 0 9 13
10 15 9 13 3 1 9 0 9 9 13
20 7 16 9 13 1 9 9 9 13 2 15 9 1 0 9 9 0 9 13 13
10 16 3 0 9 13 2 15 9 9 13
21 3 9 1 0 9 9 1 9 13 13 13 9 2 16 15 0 9 8 2 9 13
18 7 15 9 1 9 1 9 0 2 15 1 9 13 2 9 13 13 13
12 13 15 3 13 9 15 0 0 0 9 13 13
13 3 9 3 0 9 13 2 7 9 0 0 3 13
6 15 15 9 1 9 13
5 1 0 9 3 13
45 9 16 15 2 15 9 3 13 2 13 13 2 16 2 1 0 0 3 13 2 3 1 9 13 13 0 13 7 13 2 1 0 9 9 13 7 3 0 9 3 13 9 15 9 13
13 3 9 7 9 0 13 15 13 2 3 0 9 13
21 9 0 2 9 1 9 3 13 2 7 3 15 1 9 7 0 9 0 1 0 13
34 7 16 0 7 0 9 15 13 0 7 0 15 2 3 9 13 13 0 7 0 9 13 2 3 16 15 15 15 15 0 7 0 13 13
11 7 15 15 9 13 2 9 3 3 13 13
30 0 9 2 0 0 2 9 7 0 2 0 13 1 9 2 1 9 2 15 0 2 15 2 16 9 0 13 2 0 13
20 3 13 1 9 13 3 9 0 7 0 2 16 0 9 9 13 2 1 9 13
21 7 7 3 2 1 9 7 9 9 2 9 1 9 15 13 2 13 9 2 9 13
7 3 15 9 7 9 0 13
8 3 9 9 13 2 0 9 13
31 7 15 9 2 15 0 9 13 2 13 13 15 9 13 2 15 13 1 13 9 7 9 13 2 15 9 0 7 1 0 13
13 15 0 7 3 9 13 2 15 9 0 3 0 13
26 16 9 9 9 13 2 0 13 2 0 13 2 3 0 9 9 13 13 2 3 0 9 9 0 13 13
16 7 15 13 9 9 2 3 9 0 2 0 9 2 9 0 0
7 3 15 0 13 1 0 9
3 7 7 13
6 9 0 15 9 9 13
13 9 9 9 9 9 9 0 3 16 9 0 15 13
9 7 3 9 7 3 9 1 15 13
24 15 15 2 3 13 2 15 3 9 13 2 16 9 15 9 13 7 15 13 3 16 13 13 13
24 3 9 13 9 0 2 9 0 2 9 2 9 2 9 2 0 9 2 15 9 7 9 9 13
7 1 15 15 9 9 13 13
12 1 15 9 13 0 0 2 0 8 15 13 13
21 13 9 9 2 9 9 9 2 9 9 7 9 2 0 9 0 2 15 15 9 13
27 9 13 7 15 7 9 3 13 1 15 2 15 9 9 15 3 13 13 13 13 9 9 15 2 15 9 13
8 15 15 9 1 9 3 13 13
25 7 1 15 9 13 8 2 0 2 13 3 0 9 2 9 7 9 13 2 15 9 9 9 9 13
8 15 9 3 0 9 13 16 9
35 15 16 3 0 13 2 16 9 3 13 13 2 3 13 9 7 9 13 13 7 13 3 9 2 16 15 0 13 2 3 3 13 16 13 13
26 7 0 9 9 9 13 0 9 9 0 3 13 13 2 7 13 9 1 9 9 15 7 9 13 9 13
22 7 7 3 0 9 9 13 2 7 3 13 9 13 2 16 15 3 0 9 0 13 13
10 7 16 9 13 2 9 7 9 3 13
12 7 9 13 9 13 9 2 9 7 9 2 9
6 15 9 3 9 9 13
26 9 1 9 9 0 13 2 9 9 7 9 9 13 0 9 1 9 15 13 2 15 3 9 13 9 13
20 1 15 15 9 13 13 9 0 13 2 9 13 2 9 15 7 13 15 7 13
13 7 1 15 13 9 2 15 0 3 0 9 9 13
9 9 7 9 3 13 2 3 3 13
10 9 3 13 2 16 3 13 9 3 13
13 7 15 3 3 9 13 2 9 13 2 9 0 13
5 9 7 9 3 13
15 13 9 13 2 9 13 2 9 13 7 0 7 0 7 0
7 3 0 9 7 0 9 13
24 15 9 13 9 9 3 1 0 9 9 13 2 13 2 16 13 13 2 3 15 1 9 9 13
10 7 3 15 3 1 13 9 7 9 13
28 7 7 1 9 2 9 15 9 13 1 9 13 2 16 9 2 9 2 1 15 9 3 13 2 9 9 15 13
8 1 15 9 9 7 9 3 13
36 16 9 9 13 7 9 7 3 9 7 3 9 15 9 1 9 13 3 13 2 13 9 13 7 0 9 13 2 16 15 3 13 9 7 9 13
35 3 9 2 9 9 7 1 15 9 9 2 9 15 0 1 9 0 2 9 2 9 1 9 13 2 3 0 9 2 15 3 0 15 13 13
5 3 9 9 3 13
12 9 9 13 2 13 9 2 0 9 13 9 13
16 15 1 9 13 2 3 0 13 2 13 16 3 13 7 13 13
64 3 2 16 9 13 15 13 2 3 0 9 9 9 13 1 9 2 9 9 2 7 3 9 1 9 15 13 13 15 9 13 1 15 9 2 15 1 13 9 13 2 3 0 1 0 9 0 2 15 9 9 13 2 7 15 1 9 13 13 2 16 3 9 13
5 15 0 9 3 13
40 7 13 7 13 9 8 2 0 9 0 9 0 13 7 1 15 8 2 9 9 13 15 9 9 3 1 13 9 16 13 13 1 9 7 1 0 9 0 0 13
17 9 16 13 2 0 9 9 13 2 3 1 9 9 9 15 13 13
8 3 15 9 13 0 9 3 13
45 15 16 9 13 2 0 9 13 2 16 7 3 9 1 9 13 9 3 13 13 7 3 2 9 0 0 7 15 9 13 2 3 13 13 2 9 1 9 13 2 3 3 9 9 13
22 3 2 16 3 1 0 9 13 2 9 13 2 13 9 9 2 16 15 9 0 9 13
9 15 9 1 9 9 0 9 0 13
21 9 13 2 9 13 2 13 0 9 9 7 9 2 9 7 9 9 7 9 0 13
10 3 1 9 9 9 15 9 9 9 13
35 1 0 9 8 2 9 9 1 9 9 13 2 15 9 13 15 13 2 1 15 13 13 8 2 9 9 13 1 0 9 1 9 12 9 0
9 15 9 13 9 7 0 9 9 13
28 13 2 13 2 7 3 9 7 3 9 15 3 13 2 7 3 9 13 7 3 9 13 2 0 15 9 9 13
21 7 9 0 9 15 15 13 2 16 9 13 7 15 9 0 13 13 1 9 2 9
15 3 13 9 7 15 13 2 16 9 13 13 2 1 9 13
26 3 8 2 9 9 2 7 9 15 13 7 9 13 2 9 13 0 7 0 9 0 2 15 3 13 13
30 7 16 15 13 2 9 2 16 13 13 1 13 9 2 0 9 2 9 0 13 1 9 13 2 16 15 1 15 3 13
17 15 9 13 2 3 15 1 9 9 13 2 16 0 9 1 9 13
14 3 15 0 2 16 3 13 2 13 2 1 9 3 13
4 9 0 9 13
6 3 15 1 9 9 13
33 7 9 7 9 7 9 2 15 13 0 9 2 13 2 15 9 13 2 9 9 13 2 9 9 13 2 9 9 7 0 9 9 13
8 15 3 1 0 9 1 9 13
20 16 15 9 13 2 9 2 9 1 0 9 9 1 0 9 13 1 9 15 9
16 7 3 15 15 13 9 9 9 13 7 3 13 9 0 9 13
6 0 9 9 7 9 13
16 3 15 9 2 7 13 9 13 7 9 9 2 13 1 9 13
31 7 15 3 9 7 3 9 13 2 15 9 9 9 7 9 0 1 9 13 2 7 9 2 15 9 0 16 1 9 3 13
33 15 7 9 13 2 13 0 9 2 9 9 15 9 9 13 13 2 3 15 15 9 13 2 16 13 2 3 9 3 13 9 15 13
18 15 9 7 9 9 9 0 3 13 2 16 9 3 1 15 3 9 13
39 15 0 9 13 2 16 9 9 13 13 2 9 13 2 9 1 9 13 2 3 16 15 0 9 0 13 2 7 16 9 0 0 13 7 1 0 9 9 13
18 1 15 3 13 9 9 2 9 1 9 13 2 15 15 9 9 13 13
5 15 9 3 13 13
18 0 0 9 2 9 13 2 0 15 0 1 0 9 2 9 9 0 13
10 15 1 9 9 1 0 9 3 13 13
13 15 9 3 0 1 0 9 9 0 9 13 13 13
10 9 16 13 13 2 13 13 9 15 13
7 3 9 13 7 0 9 13
9 15 1 9 13 2 1 9 0 13
1 6
31 7 15 9 9 13 1 9 2 9 1 9 0 2 16 9 3 13 9 13 2 1 9 7 9 9 9 1 9 1 9 13
30 15 16 9 13 13 2 9 9 7 9 9 13 2 0 9 9 13 2 1 15 1 9 13 1 9 13 1 9 0 13
19 3 13 2 16 9 9 13 2 9 1 9 9 13 13 2 9 9 9 13
11 15 9 15 9 9 0 3 3 0 13 13
22 7 7 0 9 9 1 0 9 7 3 9 13 9 13 7 3 1 9 9 15 9 13
23 7 3 3 15 0 9 13 2 15 0 9 13 2 7 3 0 9 0 9 9 9 9 13
6 15 3 9 0 13 13
42 7 3 1 9 2 15 9 0 13 2 0 13 2 9 13 2 9 13 2 9 13 2 9 0 9 13 9 13 2 9 7 9 1 9 13 2 16 9 3 13 1 9
38 3 9 0 0 9 2 16 1 0 9 0 9 13 2 0 3 9 2 16 0 9 7 9 9 13 2 15 15 2 16 1 9 13 2 1 9 0 13
21 3 9 2 15 1 9 9 9 9 13 2 0 7 0 9 13 0 9 0 9 13
7 15 7 0 9 9 0 13
18 3 3 13 13 9 13 2 0 9 2 0 9 9 0 3 7 15 13
17 1 15 15 0 7 9 9 13 2 13 9 0 16 3 13 15 13
9 15 3 0 0 1 9 1 9 13
47 7 16 9 2 9 7 9 2 9 9 0 9 13 13 2 9 0 0 9 13 2 15 9 7 9 0 13 2 13 9 13 9 13 2 3 13 7 13 3 13 2 3 15 0 7 0 13
12 1 15 0 9 13 0 9 9 9 1 0 9
9 7 3 15 9 7 3 9 9 13
4 15 9 3 13
20 7 16 9 2 9 1 9 0 7 0 13 13 2 9 9 13 2 9 9 13
8 15 9 2 9 7 0 9 13
20 15 0 2 13 2 1 9 9 13 7 15 9 13 2 16 9 1 9 3 13
18 7 16 3 0 9 13 2 8 2 9 13 13 2 0 9 9 15 13
45 7 16 0 9 9 0 7 0 9 13 2 3 0 9 7 9 9 0 13 2 7 3 15 2 15 9 13 13 2 3 15 13 13 2 16 13 7 0 15 3 13 9 7 9 13
12 13 3 1 9 9 2 15 1 9 3 13 13
46 7 9 2 9 15 9 13 2 16 9 9 13 7 15 2 16 13 2 13 1 9 9 2 13 3 7 3 9 0 13 2 3 16 9 9 0 0 13 2 3 15 1 0 9 13 13
29 3 1 9 2 16 3 9 1 9 13 2 13 9 1 9 9 7 3 13 15 9 13 13 2 15 9 0 9 13
46 7 15 13 13 1 9 9 2 13 9 2 16 1 15 9 9 13 2 9 0 9 9 13 2 2 7 15 2 13 2 15 2 16 3 9 13 13 2 9 13 2 15 0 15 9 13
15 15 16 13 2 9 1 0 9 13 9 13 2 16 15 13
22 9 3 9 7 7 3 0 13 2 15 3 3 13 13 2 16 15 9 9 9 0 13
19 15 15 1 9 9 2 9 13 2 16 9 0 13 7 3 0 9 1 9
6 7 3 9 1 9 13
9 3 9 13 2 16 0 9 9 13
7 3 15 13 9 0 9 13
10 7 9 3 1 9 13 2 15 9 13
15 1 0 9 13 9 0 2 9 9 2 0 9 1 9 9
8 15 15 13 3 13 9 9 0
19 3 9 2 0 9 2 15 9 9 3 13 2 9 0 2 16 13 2 13
29 9 1 9 9 13 9 13 2 16 9 9 3 13 2 15 13 2 3 13 7 13 9 2 16 15 16 3 0 13
19 15 3 9 1 9 0 7 0 2 3 1 9 0 2 9 2 9 9 13
17 7 3 15 2 15 3 9 13 2 3 7 3 1 9 0 3 13
17 0 9 2 9 7 9 9 2 13 2 13 9 0 9 16 9 13
47 7 9 9 1 8 2 15 9 9 13 2 13 16 13 0 9 13 2 16 2 16 9 1 9 8 1 9 13 2 9 2 9 9 9 9 13 13 1 9 9 7 9 0 9 0 9 13
6 7 15 13 15 9 13
28 9 7 9 7 1 0 9 12 3 0 9 9 13 2 16 9 0 9 1 9 7 0 2 15 9 13 2 13
8 9 9 9 13 7 15 9 13
17 0 7 0 2 7 9 9 2 15 1 9 0 9 13 2 9 13
9 3 9 7 9 13 9 1 9 13
11 1 15 13 7 13 9 3 13 1 9 9
8 15 13 7 9 13 0 9 13
23 9 2 3 9 1 0 9 9 13 2 7 15 2 16 9 13 2 13 9 9 1 9 13
14 9 0 2 0 2 9 0 13 2 0 9 1 9 13
9 7 9 1 9 9 1 0 15 13
18 1 9 2 9 2 9 2 3 0 13 9 13 2 15 13 1 9 13
9 3 3 3 15 1 0 9 13 13
18 0 9 13 13 2 0 15 3 0 13 13 7 9 1 9 1 9 13
26 9 1 15 8 2 9 15 0 13 2 16 9 2 0 3 9 13 2 1 9 13 7 13 9 9 13
12 15 9 9 1 9 13 2 15 9 3 13 13
12 15 13 2 1 15 2 15 1 15 13 2 13
13 13 13 2 1 0 9 13 2 7 13 15 9 13
6 13 2 15 0 9 13
8 9 13 1 9 2 7 1 0
5 1 15 9 9 13
11 16 1 9 9 13 13 2 15 9 9 13
6 1 9 13 13 15 13
5 3 13 15 3 13
34 15 9 3 13 2 13 9 15 13 9 1 9 0 13 8 2 9 9 7 8 2 0 9 13 2 16 1 9 0 1 9 9 9 13
7 9 0 13 2 0 9 13
10 9 2 16 9 9 13 2 3 13 13
66 16 1 15 9 9 1 9 13 7 3 3 9 13 13 2 9 3 13 9 1 9 9 15 13 2 9 3 13 15 9 15 1 9 13 2 3 2 16 1 9 13 13 2 9 3 1 9 0 0 13 2 16 15 13 13 2 3 0 7 9 13 16 9 15 9 13
9 15 9 13 0 3 1 9 9 13
8 7 15 0 9 7 9 3 13
16 3 7 0 13 13 2 1 0 9 0 9 13 15 9 9 13
11 9 15 15 9 2 9 13 9 0 13 13
27 7 13 9 13 1 15 13 9 2 9 2 9 2 0 7 3 9 0 2 15 1 9 1 13 9 13 13
4 0 1 9 13
12 9 2 9 3 9 13 2 13 9 1 9 13
22 9 9 2 16 9 13 2 15 9 13 1 9 13 2 0 1 9 1 9 9 13 13
27 3 9 13 7 0 9 15 9 9 1 9 13 2 9 9 9 1 9 2 15 1 9 13 2 3 13 13
24 9 13 1 9 2 1 9 2 3 15 7 15 1 9 9 13 2 3 13 15 2 13 1 9
16 15 9 13 7 9 13 13 1 9 9 2 15 15 13 13 13
8 1 9 0 9 9 12 0 13
14 9 7 9 3 2 15 0 13 2 15 9 13 9 13
19 3 1 9 9 15 13 0 9 2 15 3 1 9 9 13 9 0 0 13
41 3 9 9 2 9 9 2 15 3 9 13 2 9 9 2 0 2 9 9 2 9 2 9 9 2 9 2 9 16 15 9 3 1 9 13 13 9 2 9 9 13
24 3 9 9 13 2 15 3 0 9 0 3 9 13 2 13 9 9 9 8 2 9 1 9 13
33 7 7 0 9 9 9 3 16 9 13 2 9 3 0 2 0 7 15 3 0 13 2 16 15 0 9 1 9 0 7 9 9 13
20 1 15 9 15 9 2 9 1 9 13 13 2 15 1 9 13 1 9 13 13
43 3 15 13 1 9 2 9 2 16 9 13 2 16 15 9 7 9 7 0 1 9 13 13 2 7 3 3 13 1 9 8 2 3 7 9 9 13 7 15 3 1 9 13
32 3 13 9 0 9 13 9 9 0 13 7 15 1 9 13 7 3 3 9 13 2 16 1 15 13 2 15 9 0 9 13 13
24 13 15 9 15 13 9 15 1 9 2 9 13 2 16 3 13 9 1 9 9 0 15 9 13
17 9 9 1 9 9 13 2 16 9 9 0 13 9 9 9 0 13
13 15 9 15 3 13 13 0 15 9 15 1 9 13
36 7 15 9 8 2 9 7 8 2 9 2 7 3 9 2 7 3 9 7 7 0 9 13 13 2 16 1 9 7 0 9 8 2 9 3 13
32 9 13 1 9 9 13 1 15 0 9 0 2 9 1 9 9 9 13 2 16 0 9 2 0 9 13 2 1 9 9 13 13
17 9 7 0 13 2 16 15 3 0 9 2 3 0 9 0 9 13
69 7 16 9 1 0 9 13 13 2 15 3 13 7 13 2 15 15 1 9 7 9 13 13 2 0 15 9 13 2 3 3 16 0 9 0 2 15 9 9 1 9 13 1 9 9 2 7 9 9 7 9 9 13 2 16 9 0 1 9 0 0 13 2 13 1 9 9 9 13
27 9 7 1 9 9 7 9 0 2 0 7 13 2 13 2 1 9 2 2 16 9 13 1 9 1 15 13
30 9 16 15 13 13 2 13 9 2 3 9 7 9 13 2 13 9 13 2 15 1 15 13 13 2 15 1 9 13 13
11 7 15 9 3 0 9 13 1 9 0 13
50 3 8 2 0 9 0 9 13 2 16 15 9 9 13 13 2 1 15 2 15 1 9 13 2 7 3 1 8 2 0 2 8 2 0 2 8 2 9 2 8 2 9 2 16 13 13 2 9 13 13
26 7 15 3 13 9 8 2 9 9 1 9 8 2 9 13 15 13 2 15 1 0 9 9 13 13 13
18 7 9 2 16 1 15 13 13 2 13 9 1 9 15 9 9 13 13
23 0 9 2 9 13 2 15 1 9 0 13 2 1 9 2 9 2 9 7 9 0 13 13
19 3 3 9 9 13 2 16 15 13 2 7 3 15 0 9 3 7 9 13
5 16 13 9 2 13
10 16 9 13 2 15 13 2 9 3 13
19 0 15 9 13 13 2 9 13 2 15 9 7 9 9 7 9 13 3 13
16 7 15 13 13 2 15 9 0 1 9 9 15 3 7 9 13
26 9 0 2 15 1 9 9 13 2 9 9 0 7 0 2 15 9 0 9 13 2 0 7 13 15 13
26 7 16 9 13 1 9 13 13 2 9 0 2 16 15 9 3 3 9 9 9 13 13 2 13 15 13
25 3 9 0 0 2 16 3 0 7 1 9 7 1 9 0 0 9 13 2 3 15 1 9 0 13
15 3 15 15 0 13 2 3 15 1 15 9 13 13 2 13
15 16 9 9 9 9 13 2 15 13 13 2 15 9 13 13
10 15 9 9 13 2 15 13 13 2 13
4 13 9 2 9
5 13 9 1 9 9
6 9 9 13 15 9 8
4 9 7 9 13
4 9 2 9 13
10 3 9 2 9 2 9 7 9 0 13
10 7 2 1 9 0 2 3 15 9 13
14 3 2 15 9 0 7 3 0 3 13 2 15 9 13
8 7 0 0 9 13 2 9 13
21 15 13 1 9 9 13 2 16 15 9 13 2 0 13 2 9 7 9 15 0 13
14 15 0 9 0 1 9 9 13 2 15 9 0 0 13
7 3 1 0 9 0 9 13
11 7 7 13 7 7 13 2 7 3 13 13
13 15 1 0 9 13 2 15 1 9 9 7 9 13
7 3 15 3 13 2 9 13
7 0 9 0 3 9 15 13
22 7 7 0 0 3 13 7 1 9 0 9 15 13 1 9 13 2 16 15 0 0 13
28 8 2 9 2 9 0 7 0 2 3 13 15 13 9 9 0 13 2 7 3 15 1 0 9 9 7 9 13
7 15 9 7 15 9 9 13
17 1 9 0 13 13 2 16 3 9 0 9 9 0 9 13 1 9
5 15 0 0 0 13
9 3 7 7 9 7 7 9 9 13
20 7 2 1 9 0 2 15 1 9 1 9 3 13 2 16 3 9 1 15 13
14 7 0 9 3 13 9 3 9 13 2 7 9 13 13
12 15 7 0 7 3 0 13 1 9 0 9 13
18 16 16 0 13 2 3 13 1 0 9 9 13 2 16 15 1 0 13
11 7 7 15 13 15 1 9 9 0 13 13
5 15 9 13 15 13
12 3 15 2 9 13 2 15 1 0 13 2 13
8 0 0 9 1 9 0 13 13
24 7 3 9 1 0 15 7 3 0 13 2 0 15 9 1 0 7 0 1 0 7 3 0 13
12 0 13 9 12 9 13 2 15 9 0 15 13
10 15 3 13 0 15 7 0 13 0 13
7 15 9 13 7 9 13 13
16 3 16 3 9 13 2 3 0 7 0 3 13 2 0 9 13
9 3 9 9 13 0 9 0 9 13
25 0 9 9 9 16 9 7 0 15 9 2 15 0 9 0 13 2 13 13 2 15 3 9 15 13
14 9 0 7 0 2 15 9 9 0 13 2 9 13 13
7 7 15 9 0 9 9 13
27 3 15 2 15 9 9 9 13 2 0 3 15 13 2 7 3 3 9 13 13 2 3 9 0 0 9 13
23 7 15 15 3 1 8 2 9 7 3 15 9 13 2 7 1 0 9 0 7 0 9 13
19 13 0 9 2 0 9 2 15 3 9 1 9 13 2 9 15 1 9 13
17 3 15 9 1 9 9 9 9 13 2 15 15 9 13 7 15 13
14 0 0 2 9 13 2 7 3 9 7 3 9 3 13
17 7 3 15 9 13 2 3 0 0 9 2 16 3 0 13 2 8
13 9 7 9 0 1 9 2 9 9 1 9 0 13
16 3 2 15 3 1 9 7 9 0 13 2 1 0 9 9 13
5 13 3 13 9 13
17 7 15 15 9 9 9 13 9 13 1 9 2 1 13 0 9 13
26 3 9 7 9 0 15 13 2 15 1 0 9 0 9 13 2 16 1 15 2 15 15 3 13 3 13
8 13 7 15 13 7 13 9 9
3 7 3 13
12 3 15 1 15 3 1 9 13 3 1 9 13
14 15 3 13 2 9 13 15 1 9 0 7 9 0 13
12 16 9 13 9 13 2 0 9 0 0 3 13
11 7 8 2 9 9 13 9 15 9 9 13
23 3 0 15 9 13 2 9 13 2 16 9 7 9 0 13 2 7 16 9 9 15 15 13
19 15 15 13 13 1 9 15 2 15 9 2 9 2 9 7 9 0 9 13
13 9 7 13 13 1 15 3 3 15 1 15 13 13
9 7 0 9 3 13 2 16 13 13
12 15 16 13 16 13 2 16 13 2 3 9 13
6 13 9 9 13 0 13
25 7 2 1 9 0 2 15 15 13 2 15 3 9 2 9 2 9 2 9 0 0 16 9 0 13
9 3 13 1 0 7 7 1 9 9
7 9 7 9 0 1 0 13
29 3 2 9 13 2 0 9 1 15 9 13 2 3 1 9 7 9 0 9 13 13 2 7 0 0 15 9 13 13
18 15 15 7 9 0 0 3 9 9 13 2 3 3 0 9 3 13 13
16 7 15 16 15 0 13 2 3 9 0 0 13 2 9 9 13
7 3 15 15 9 7 9 13
8 3 3 3 15 0 9 9 13
19 16 0 0 13 9 2 0 9 9 9 13 2 3 9 0 1 9 13 13
19 13 3 2 16 3 15 9 13 2 0 1 0 9 2 13 0 1 9 9
16 3 15 9 0 13 7 2 16 0 13 13 2 0 0 13 13
26 3 7 3 8 2 9 0 3 1 15 9 1 9 7 9 13 2 13 0 13 15 2 15 1 9 13
14 13 9 0 1 0 9 0 2 0 2 0 7 0 13
33 3 13 9 15 13 2 15 1 9 1 9 13 2 3 13 2 16 2 16 9 13 2 7 1 9 9 7 1 9 0 1 9 13
28 3 9 0 7 0 3 1 9 7 3 1 0 9 13 2 7 3 3 0 13 9 2 16 1 13 9 0 13
12 3 9 3 15 9 13 2 16 9 1 15 13
17 16 1 0 0 9 0 3 13 2 3 3 13 15 15 7 15 13
11 3 15 3 15 13 2 3 15 9 0 13
11 16 0 9 15 13 13 2 3 0 0 13
11 13 13 9 0 9 9 0 1 0 0 13
9 16 3 13 2 0 0 15 15 13
15 3 9 7 9 2 3 9 7 9 0 9 15 16 15 13
13 7 0 13 2 15 15 0 13 2 15 15 0 13
13 1 15 15 13 9 7 9 2 3 9 2 3 9
5 13 9 2 13 9
12 1 0 7 0 9 0 2 0 9 9 9 13
28 3 15 3 15 15 9 13 2 3 9 9 2 3 9 7 9 13 2 3 13 2 3 9 13 1 0 9 0
4 7 15 15 13
22 13 0 9 9 13 2 9 9 0 9 0 1 9 13 2 9 9 1 9 1 9 13
13 15 13 3 3 7 13 2 15 1 9 13 9 13
11 13 13 13 9 9 1 9 7 3 9 13
15 3 15 15 9 7 9 2 16 15 9 13 2 1 9 13
11 3 9 15 0 13 2 7 15 3 13 15
24 7 9 7 9 9 0 9 13 13 2 3 9 0 13 2 15 15 9 0 3 1 0 9 13
9 3 9 7 3 9 0 9 9 13
9 13 2 13 2 3 13 0 0 13
10 16 9 15 7 9 13 2 3 9 13
4 13 7 0 13
32 1 9 0 8 2 0 9 9 0 9 0 2 16 15 1 9 1 9 13 2 13 13 2 7 15 0 9 0 9 9 9 13
8 15 1 0 9 15 13 2 13
7 3 0 9 15 15 9 13
20 0 13 9 9 2 16 15 9 2 16 9 0 2 16 9 7 9 3 0 13
9 13 9 9 2 16 3 9 9 13
10 7 15 15 1 0 2 9 2 9 13
14 15 16 15 3 9 13 2 3 15 9 1 9 0 13
4 7 3 13 13
5 9 1 9 9 13
9 0 1 9 7 1 9 9 13 9
9 7 3 13 7 7 13 15 13 3
4 15 3 13 13
26 16 9 13 2 9 0 7 3 9 0 9 9 15 13 2 9 9 1 9 13 2 0 0 13 0 13
5 9 0 7 0 13
7 9 9 13 2 16 15 13
32 7 15 0 13 2 0 13 2 15 9 0 9 7 9 2 9 7 9 0 9 13 2 9 13 13 2 15 9 3 0 9 13
9 13 3 0 9 1 0 9 9 13
25 13 0 9 9 13 1 0 9 2 1 15 3 9 9 13 2 9 0 2 9 9 9 1 9 13
23 7 15 0 13 13 9 9 0 9 0 13 2 7 3 9 2 16 9 9 2 9 9 13
35 7 16 9 7 9 9 13 13 2 3 9 0 9 0 9 7 9 9 13 7 2 3 0 9 9 2 0 9 3 3 15 9 9 0 13
10 1 0 0 9 13 2 1 0 0 9
6 15 9 2 15 9 13
8 3 9 1 9 13 13 2 13
12 9 9 13 0 13 2 9 13 15 9 0 13
14 15 0 9 2 9 2 9 0 13 2 16 9 13 13
11 7 9 9 9 2 9 2 7 3 9 13
23 3 9 1 9 7 3 9 1 0 2 7 1 0 9 2 1 0 9 2 1 9 9 13
5 13 16 13 0 13
33 16 2 16 13 2 9 1 9 9 13 2 9 0 9 13 9 15 13 13 2 16 15 15 9 13 2 9 15 1 9 13 13 13
7 15 9 13 9 1 9 13
5 15 13 9 1 9
20 13 1 9 9 2 15 0 13 2 16 3 13 1 9 2 1 12 9 9 13
10 9 13 3 9 7 3 9 0 9 13
19 1 15 9 16 13 13 9 2 9 9 0 2 15 9 13 2 9 9 13
22 3 15 0 1 9 0 0 2 15 0 9 9 13 2 0 9 7 9 0 9 9 13
13 1 9 2 9 2 0 2 9 15 9 9 13 13
27 16 15 9 13 2 9 1 0 9 2 15 7 15 13 7 0 13 2 0 9 13 2 9 1 9 9 13
30 3 2 16 15 0 7 1 9 1 9 13 2 3 13 2 7 0 9 9 9 9 13 2 16 9 3 0 0 12 13
11 7 1 0 9 3 9 0 13 0 9 13
15 0 2 16 15 9 13 2 9 7 9 2 0 13 9 13
12 13 3 0 9 15 13 2 16 9 9 13 13
28 3 9 13 2 15 9 1 15 0 9 13 2 9 9 0 2 3 0 0 9 13 13 9 9 1 9 0 13
22 0 9 1 9 0 0 9 1 9 0 13 15 9 2 16 1 9 3 13 1 9 0
24 7 8 2 9 0 1 12 9 1 9 0 13 2 1 9 9 15 15 13 15 3 13 9 13
25 7 16 9 15 1 9 13 2 9 3 13 7 1 15 9 9 13 2 3 15 9 13 1 9 13
17 7 3 3 9 3 13 2 3 15 0 9 9 0 13 1 9 13
41 7 9 3 13 9 7 9 9 15 13 2 1 9 9 13 2 7 3 9 7 3 9 0 9 2 0 9 13 1 0 9 9 9 13 2 13 1 9 3 3 13
7 3 9 13 15 9 9 13
11 15 7 3 9 7 3 9 13 2 3 13
4 9 9 9 13
16 7 15 15 2 3 0 13 2 13 2 3 16 9 0 9 13
12 3 3 15 9 9 0 13 2 3 15 9 13
12 9 9 0 2 0 1 9 2 0 1 9 13
17 3 1 15 9 13 2 16 3 9 13 2 9 7 0 9 9 13
8 3 13 13 2 9 9 13 13
32 3 15 13 2 16 0 7 13 9 13 7 2 16 9 13 2 13 15 9 2 9 2 9 2 3 9 7 9 1 9 0 13
7 16 13 2 9 15 13 13
7 9 3 2 9 7 9 13
21 16 9 13 2 15 15 13 13 2 7 3 9 7 3 9 15 13 15 9 3 13
11 3 2 9 2 3 15 15 7 15 9 13
10 15 1 9 2 1 9 2 1 9 13
7 15 0 13 13 1 9 0
6 3 3 13 0 0 9
18 13 15 1 0 9 1 9 9 13 2 13 0 9 13 0 0 9 13
11 16 15 0 7 13 9 13 2 15 13 13
8 16 15 13 13 2 9 9 13
6 9 16 9 9 9 13
11 3 1 9 15 0 13 9 2 15 3 13
4 9 1 9 13
17 16 15 13 2 9 2 7 16 9 0 13 2 0 15 9 9 13
15 9 9 9 0 15 13 2 3 9 2 15 3 0 0 13
10 7 9 9 16 13 13 2 13 9 9
29 7 16 9 0 9 13 2 13 0 9 13 2 3 13 3 3 9 13 2 3 9 9 13 0 7 0 9 9 13
16 15 16 13 2 3 13 9 13 13 7 13 9 1 9 0 13
21 3 13 9 9 2 3 9 13 9 9 0 13 2 15 9 9 1 9 7 9 13
26 7 2 16 9 13 1 0 9 7 1 0 9 0 2 12 9 1 9 13 2 0 9 1 9 3 13
20 1 15 9 2 0 0 7 0 2 3 1 0 9 0 15 13 1 0 9 13
19 15 1 9 7 9 1 9 13 2 15 9 0 8 2 9 1 9 13 13
21 7 1 0 9 8 2 9 2 9 0 16 9 13 13 2 8 2 9 9 9 13
19 15 9 0 2 15 9 9 13 2 1 9 2 1 15 0 9 1 9 13
30 15 9 13 0 15 13 13 2 13 2 13 2 16 13 15 1 9 0 1 9 2 1 9 2 1 9 7 9 0 13
5 15 13 9 9 13
14 7 16 0 9 13 9 9 9 13 2 9 3 13 13
4 15 13 9 9
18 16 3 13 13 2 3 1 9 9 13 13 2 0 9 1 0 9 13
6 9 13 2 9 9 13
12 0 0 9 0 3 3 13 2 15 3 0 13
3 0 9 13
27 3 9 1 9 1 0 9 13 2 13 13 2 0 1 0 13 2 9 13 2 0 15 13 2 3 9 13
8 0 9 7 0 9 9 3 13
28 9 3 13 9 2 3 3 13 13 2 0 9 13 2 9 0 1 0 9 13 7 15 13 7 0 3 13 13
6 3 3 1 9 0 13
7 9 7 9 1 0 13 13
25 9 16 13 9 7 15 1 0 13 13 2 0 9 7 0 0 9 1 0 9 13 7 3 13 13
18 7 13 9 2 3 3 13 2 0 9 7 0 9 9 13 1 9 9
14 7 3 15 15 0 13 9 13 2 15 13 9 9 13
18 0 7 2 15 0 9 0 13 2 9 3 2 7 9 3 13 9 13
25 9 7 3 1 0 1 9 9 13 13 2 3 7 13 7 9 9 2 15 13 0 2 1 9 13
17 3 1 0 9 7 3 1 9 7 3 1 9 15 9 0 13 13
8 3 0 0 7 9 9 3 13
12 7 7 3 9 9 0 0 7 0 9 13 13
11 7 0 15 7 13 1 9 7 3 13 13
6 13 3 15 9 0 13
13 3 3 1 0 9 9 2 9 2 9 7 9 13
15 3 13 13 2 7 9 13 9 2 7 3 0 9 13 9
3 13 9 9
12 3 9 0 9 13 9 2 7 9 0 13 9
7 9 9 13 13 9 1 0
7 3 13 9 9 7 0 9
32 9 2 16 9 13 2 13 0 9 2 0 9 13 15 13 9 2 0 1 9 0 13 1 9 2 7 0 0 3 1 13 9
17 13 15 3 9 2 15 2 9 2 13 9 9 2 7 13 0 9
4 13 13 9 9
6 3 13 9 13 0 9
18 0 9 7 3 13 9 9 15 9 9 7 9 13 2 0 13 9 9
14 15 3 0 9 9 1 0 2 13 9 2 9 2 13
7 3 13 13 9 13 1 9
4 3 9 13 9
7 3 15 15 15 9 9 13
14 3 9 1 0 12 13 9 13 2 3 13 1 9 0
16 13 0 9 0 9 1 9 2 15 0 13 9 12 2 9 12
7 13 13 1 9 2 16 9
4 13 9 9 13
17 15 0 13 1 9 3 3 9 2 3 9 0 2 3 13 13 9
1 13
4 7 0 13 13
15 0 9 1 0 13 9 9 2 7 13 9 9 9 1 0
44 9 2 0 9 3 13 9 2 0 15 9 13 9 7 9 9 1 9 2 0 13 9 0 9 13 9 15 2 7 3 13 9 9 7 13 9 9 2 3 3 9 13 13 9
6 3 0 3 13 9 13
21 15 3 0 3 9 13 13 9 2 7 9 7 9 0 15 13 9 7 0 9 9
16 3 9 7 9 0 1 9 9 13 2 7 0 9 1 9 9
7 15 3 0 13 9 0 0
23 3 15 7 7 0 9 7 0 9 2 13 0 9 2 13 2 7 13 13 2 0 2 9
12 9 3 3 9 13 2 16 13 13 0 9 9
3 15 13 13
4 9 13 9 13
9 7 3 3 3 13 13 0 9 9
18 7 2 9 3 13 2 0 1 9 13 9 2 0 16 9 13 13 9
14 3 3 15 13 9 0 2 0 9 13 2 7 13 13
15 9 3 9 13 0 12 9 0 2 7 9 13 9 1 9
4 7 9 0 13
5 1 9 9 9 13
5 13 15 1 9 9
5 7 3 7 13 13
13 3 9 15 2 7 3 9 2 7 3 0 9 13
10 0 9 3 13 9 2 13 7 15 9
15 15 3 13 9 2 7 3 13 13 2 3 0 15 9 13
12 9 0 9 2 15 3 13 2 0 13 1 9
7 7 3 9 13 9 3 13
16 0 1 9 13 0 9 13 13 9 7 9 13 2 0 0 13
11 15 9 13 13 2 7 9 1 9 13 9
12 16 3 13 9 7 0 9 13 2 13 9 9
13 3 0 9 2 6 9 2 0 15 9 7 0 13
7 0 13 7 9 15 3 13
2 0 13
6 13 9 7 0 9 13
17 15 15 1 9 7 12 13 9 13 15 9 2 7 0 1 9 13
15 6 2 16 15 9 13 7 0 9 13 2 15 13 13 13
14 2 13 7 3 0 2 7 3 15 3 9 9 13 0
13 0 13 13 2 7 9 13 2 16 3 13 13 9
7 9 7 9 13 0 9 9
11 13 0 0 9 2 7 9 9 13 13 0
32 7 16 0 9 9 2 16 0 9 13 2 3 0 13 9 2 3 0 13 9 2 7 0 13 13 9 2 13 2 15 13 3
15 13 9 0 0 7 9 7 0 9 9 2 9 0 13 0
10 15 13 0 9 2 7 0 13 9 9
14 7 3 3 13 9 13 13 2 0 3 15 13 9 9
8 15 15 0 0 13 9 9 13
12 0 13 3 13 0 0 2 7 0 13 9 9
10 3 3 13 9 2 7 3 9 13 9
11 7 15 13 7 0 13 2 16 15 9 13
12 3 3 9 0 13 2 7 3 0 13 13 9
8 9 15 13 3 0 7 13 9
3 13 0 9
4 15 0 9 13
9 3 3 9 9 7 9 0 0 13
6 13 2 7 13 13 9
16 9 0 13 9 9 13 2 13 9 2 7 0 13 9 9 15
11 15 0 9 13 9 2 7 0 9 9 13
15 9 15 0 13 9 2 9 1 7 9 9 0 13 7 9
18 16 15 9 9 13 9 2 0 9 15 0 9 13 9 2 3 0 13
34 7 3 2 9 0 16 13 9 9 2 0 2 7 9 13 1 9 9 2 0 13 9 2 16 13 0 13 2 1 9 9 0 13 9
10 3 0 0 3 9 13 2 3 0 9
19 3 9 9 2 3 9 2 13 13 2 7 9 9 13 9 7 9 13 13
21 13 9 2 13 9 9 9 2 7 0 9 9 7 0 9 13 2 13 0 9 9
17 7 15 15 0 0 1 9 13 2 13 9 0 2 7 3 9 13
21 3 15 13 13 2 0 16 9 9 0 1 9 9 9 13 13 2 7 0 13 9
10 3 0 9 0 13 9 2 7 0 13
24 13 9 2 6 2 16 0 9 13 2 7 9 1 9 13 1 9 2 16 0 0 13 9 9
13 3 9 9 13 2 13 15 9 13 2 3 13 13
12 13 15 3 13 13 2 7 9 13 9 13 13
32 3 16 13 1 9 3 13 0 2 13 15 0 2 7 0 1 9 13 9 13 0 1 9 13 2 0 3 9 1 9 9 13
36 3 13 9 0 9 9 9 13 0 2 15 3 0 13 9 2 7 0 9 0 13 9 2 0 13 9 9 13 0 9 2 3 0 13 9 9
14 13 9 3 7 0 13 13 2 7 9 13 1 9 9
15 7 3 3 9 9 1 0 0 13 9 2 7 0 13 9
12 7 15 2 6 2 0 3 13 9 2 0 9
27 9 0 9 7 9 13 0 13 9 2 15 9 0 13 9 2 7 0 3 9 13 2 7 13 3 13 9
15 9 0 9 7 0 13 9 13 2 7 9 13 13 7 13
2 13 9
10 13 13 0 9 2 9 2 13 9 9
20 16 13 9 7 9 13 9 9 7 0 13 9 2 7 9 13 9 13 9 0
23 15 3 9 0 13 9 2 13 9 0 7 9 0 9 2 7 13 9 2 7 13 0 9
35 7 0 9 0 9 9 13 2 7 0 9 9 2 7 9 7 9 2 9 1 0 2 15 3 9 1 15 13 2 7 0 13 1 9 9
15 7 3 3 3 9 1 9 9 13 2 7 9 0 9 13
7 15 13 2 3 13 13 9
27 9 0 13 7 0 0 9 2 0 2 13 9 0 7 9 9 2 15 1 3 0 13 3 13 13 9 9
10 0 15 9 0 9 13 9 1 0 13
6 3 9 9 13 9 9
13 12 3 3 13 9 9 13 2 7 9 13 9 9
9 13 0 9 2 7 0 9 13 9
20 15 0 9 9 9 9 9 7 0 9 9 13 2 7 0 15 2 9 2 9
21 3 0 9 0 13 9 2 7 0 13 9 9 9 2 0 7 3 9 13 13 9
30 3 7 2 0 1 9 9 7 9 2 1 9 13 9 2 7 9 13 13 9 2 7 13 9 13 1 9 2 13 9
14 3 6 3 13 2 0 2 13 9 2 7 0 13 9
8 3 13 2 13 9 15 13 13
7 15 9 3 0 13 9 13
9 7 15 13 9 2 7 9 13 9
10 13 9 0 13 9 0 9 7 9 13
16 13 0 0 1 9 1 9 2 7 1 9 9 0 7 0 9
15 9 1 15 2 7 0 1 9 9 9 7 0 13 9 9
25 1 9 9 7 0 9 13 9 0 2 0 2 15 9 9 3 0 13 13 2 7 9 1 0 13
31 9 1 9 13 2 7 9 0 2 7 0 9 2 7 9 9 13 13 2 7 9 13 9 2 9 7 9 7 9 0 9
37 13 3 13 0 9 9 9 2 7 13 9 13 13 2 7 2 16 13 9 0 1 9 9 13 13 0 1 9 9 2 13 2 7 3 9 13 9
14 0 3 9 7 0 9 9 13 2 7 0 9 13 9
10 13 9 9 2 0 1 9 9 13 9
24 15 9 9 13 2 7 9 13 2 7 0 13 9 9 2 3 0 2 7 0 9 7 0 9
12 13 13 0 13 9 2 7 13 9 9 0 9
15 9 7 0 3 15 3 13 15 2 7 0 3 13 13 9
18 9 2 13 7 7 13 9 2 13 13 6 9 2 15 13 9 1 9
7 15 3 3 13 13 0 9
11 15 0 2 15 13 2 0 7 0 9 13
7 15 2 15 13 9 2 13
8 12 13 9 7 13 15 9 1
6 3 3 13 9 13 13
15 13 9 13 7 9 13 2 0 13 2 7 9 9 13 0
14 7 3 9 13 13 7 0 9 13 3 3 9 9 13
17 7 15 13 9 2 7 15 9 9 15 13 2 15 9 9 0 13
8 1 0 13 9 13 13 9 9
23 9 2 9 2 16 15 13 3 15 2 13 0 7 0 1 9 9 1 0 0 13 9 9
20 1 9 7 9 7 15 13 0 9 0 13 0 9 9 1 9 2 15 13 0
33 15 9 16 0 13 0 9 2 13 7 2 9 3 13 0 2 0 0 13 9 9 2 0 9 7 0 9 13 9 2 7 9 13
4 13 9 0 13
7 13 9 0 2 9 0 0
7 0 9 13 2 9 0 15
11 15 9 13 9 1 0 9 13 7 0 9
9 15 9 0 9 7 0 0 13 9
17 15 9 13 2 15 2 16 9 9 13 2 3 13 0 13 9 9
31 3 16 0 9 13 9 2 0 15 9 7 9 13 0 0 9 13 7 3 7 3 9 2 1 15 9 2 9 7 9 13
6 0 3 9 9 13 13
20 3 15 1 9 9 3 0 15 9 13 2 15 12 15 13 13 0 0 9 9
17 7 16 9 9 13 2 3 15 1 0 9 7 1 0 13 9 9
13 3 15 2 3 0 9 13 9 2 13 13 0 9
10 1 9 13 0 2 1 9 0 13 9
3 0 3 13
11 7 0 9 9 13 13 2 16 9 0 13
15 13 15 9 2 13 0 9 2 9 9 7 9 7 9 9
13 15 16 9 3 13 9 2 15 13 3 9 13 13
29 7 3 2 6 9 2 13 13 13 15 2 16 15 2 15 9 2 15 15 7 13 7 13 2 13 9 9 9 9
8 13 9 7 9 13 13 0 13
24 3 2 16 9 0 13 9 0 0 13 9 2 13 0 13 9 9 0 9 13 7 0 13 9
13 13 16 9 13 9 9 2 9 15 3 9 9 13
9 15 3 9 2 9 15 13 2 13
9 15 3 13 2 15 13 9 2 13
5 13 0 9 9 9
13 15 13 0 9 13 9 7 9 0 13 1 9 9
11 0 9 13 2 0 9 13 3 13 2 13
5 0 13 15 9 9
11 9 13 9 13 9 7 1 9 0 9 9
14 9 3 9 7 0 9 9 13 2 13 16 0 9 9
9 9 13 13 9 2 7 9 13 13
19 13 3 0 9 9 7 3 13 2 13 9 15 2 9 0 2 7 13 0
5 7 3 13 0 9
8 9 0 9 0 13 9 15 13
5 15 15 13 9 9
5 7 3 13 15 13
23 13 1 9 0 9 0 9 9 13 2 7 3 0 3 13 9 13 9 2 3 9 13 9
14 15 3 13 9 2 15 9 9 1 9 0 13 9 9
13 13 15 13 2 7 13 9 9 13 7 3 13 13
18 1 15 13 9 9 2 7 13 9 9 13 1 9 7 3 3 9 13
8 1 9 13 9 2 1 9 9
7 13 9 7 0 13 9 9
16 9 0 13 2 0 9 9 2 3 9 13 2 0 9 9 13
3 13 0 9
7 7 3 9 0 13 0 13
7 3 9 13 2 0 13 9
4 1 9 13 13
12 13 3 9 15 13 13 2 3 13 9 2 9
14 9 9 9 9 13 7 9 13 13 2 9 9 9 13
33 13 3 0 9 9 9 9 2 7 2 15 13 9 0 0 9 0 2 13 2 15 13 13 1 9 9 2 3 9 13 13 13 9
21 0 13 2 15 16 13 9 9 2 9 9 13 13 7 9 0 0 9 13 9 0
7 3 13 1 0 13 9 9
16 7 13 2 16 9 0 3 1 9 9 13 9 7 0 13 9
24 13 3 1 9 13 2 13 9 2 15 9 2 15 9 7 13 9 9 13 7 9 9 13 13
5 9 13 9 13 9
15 3 0 9 13 1 9 7 15 13 13 9 9 7 13 9
10 0 9 13 9 2 0 0 13 9 9
8 9 0 9 2 0 13 9 9
9 9 13 9 2 13 7 9 7 9
10 7 3 9 3 13 9 13 2 13 9
6 3 0 13 1 9 9
14 13 9 7 13 9 9 13 2 7 0 13 9 0 9
16 8 3 9 13 0 13 9 9 2 7 15 0 9 13 0 9
3 13 15 9
17 15 16 9 9 13 0 2 2 3 13 9 0 3 2 13 2 13
3 9 13 0
3 3 9 13
10 13 9 7 9 13 9 0 0 13 9
1 13
12 15 13 7 9 9 13 7 0 13 1 9 9
5 15 9 0 9 13
8 7 15 13 7 9 9 13 9
21 13 13 1 0 9 9 7 9 9 3 7 9 7 9 7 9 1 0 13 0 9
7 3 9 7 9 0 9 13
3 9 9 13
4 13 3 9 9
32 13 15 9 2 9 13 0 0 7 13 9 3 2 16 3 13 2 15 1 9 7 13 9 9 13 2 15 0 9 13 1 9
17 13 1 0 2 16 9 13 2 9 9 2 7 9 13 0 9 9
16 7 2 3 3 0 9 13 9 2 3 3 0 13 0 9 9
22 13 1 9 9 7 9 7 9 9 2 7 9 13 9 7 0 13 9 7 13 9 13
16 7 13 3 9 2 7 13 13 2 1 9 13 9 0 13 9
12 13 9 0 9 9 2 7 13 0 0 9 9
4 0 9 9 13
10 15 9 13 2 15 0 13 0 9 9
15 9 3 9 13 0 9 0 2 9 9 2 7 13 9 9
31 3 16 9 2 16 9 13 9 2 1 9 9 0 9 13 13 2 0 9 7 9 9 13 7 0 9 2 15 3 9 13
15 3 15 0 15 7 3 13 9 9 13 7 15 13 0 9
44 9 16 0 13 9 9 7 13 9 1 12 3 12 0 2 7 13 13 1 12 3 12 0 2 0 12 7 9 9 12 2 9 13 7 9 9 13 7 9 9 13 7 9 9
39 3 9 9 13 2 0 13 9 9 2 9 13 7 9 13 13 2 13 9 2 13 9 13 9 2 7 1 9 0 13 9 9 13 7 9 13 1 9 13
3 13 9 13
17 15 16 13 0 7 13 13 0 9 9 2 9 9 3 9 13 13
3 13 9 9
10 15 3 3 9 3 13 9 0 0 3
5 13 3 3 9 9
16 15 15 2 16 1 15 9 13 13 2 3 9 2 13 2 13
6 15 0 9 13 9 13
3 15 13 13
23 7 7 15 2 13 15 2 16 15 3 9 13 2 15 13 2 9 2 7 15 3 9 13
12 6 3 13 9 13 0 9 7 9 13 13 9
16 3 9 1 15 13 0 0 2 3 13 9 2 7 9 9 13
4 13 2 7 13
10 13 0 13 9 7 9 1 0 13 9
3 0 9 13
14 13 3 0 9 2 3 3 0 2 3 3 9 0 13
26 3 16 13 13 9 9 7 9 2 13 9 13 1 9 9 2 15 9 0 13 9 7 13 1 9 9
53 16 9 13 9 2 13 0 0 9 7 0 13 13 9 9 7 3 2 16 9 2 13 2 9 0 13 13 2 16 13 9 9 2 13 2 9 2 15 9 9 0 0 9 13 2 7 13 13 9 2 0 2 9
6 13 9 13 7 9 13
16 13 9 7 13 9 7 13 13 9 7 9 1 9 0 13 9
30 13 3 2 7 13 9 9 9 0 7 9 9 13 13 2 7 13 15 9 0 13 9 2 7 13 13 13 0 9 9
13 3 13 0 0 9 9 13 9 15 1 7 15 13
25 3 9 0 9 9 13 7 2 7 0 2 13 2 13 9 15 2 7 0 13 7 0 9 9 13
5 13 15 1 9 13
12 9 9 16 9 13 13 2 9 3 1 0 13
5 3 0 12 13 9
4 7 15 13 13
14 13 7 13 9 7 9 13 7 13 9 0 1 9 13
35 3 16 13 7 9 0 15 13 2 3 15 2 3 3 0 2 13 9 13 9 2 7 2 16 1 9 13 2 3 13 3 7 0 0 9
10 15 0 13 7 13 13 2 13 1 9
9 15 3 9 13 2 1 15 9 13
20 1 0 9 9 9 9 13 9 9 9 13 9 2 7 1 0 13 13 9 9
14 3 9 0 13 7 13 9 7 9 13 15 13 9 9
45 3 16 13 0 0 9 9 7 0 0 9 13 9 7 0 0 13 9 9 2 0 9 13 0 9 13 2 7 1 15 15 3 13 1 15 13 9 2 15 0 7 0 0 13 9
14 7 15 1 9 3 0 9 13 2 0 13 9 0 9
17 3 16 9 13 7 9 7 9 2 13 2 7 1 15 13 0 0
18 16 13 9 9 0 2 9 0 0 9 13 2 7 0 9 9 0 13
23 15 3 13 2 7 15 3 2 0 9 2 3 13 2 7 9 0 2 0 9 2 9 13
5 0 9 1 9 13
29 15 9 0 2 7 3 0 9 3 16 1 9 7 9 0 9 2 12 0 9 13 3 9 13 13 1 9 0 9
18 3 9 9 13 13 9 2 13 0 0 9 9 2 9 13 9 9 13
14 3 9 15 9 7 9 7 9 13 2 0 13 9 9
14 3 9 13 2 7 0 13 9 9 13 1 15 9 9
15 15 9 13 15 13 13 9 13 0 2 7 3 9 13 0
14 13 2 7 3 9 13 0 9 3 0 13 0 9 0
19 13 7 13 13 9 9 0 0 9 13 9 8 0 13 0 9 9 13 9
6 13 15 2 13 15 9
9 15 13 2 13 13 7 9 13 0
10 15 13 2 13 13 7 13 1 9 9
19 3 0 13 2 13 0 9 13 9 9 7 0 9 9 13 7 13 0 9
6 9 13 13 1 9 9
27 0 15 13 2 3 13 13 0 7 0 9 9 0 13 2 7 7 15 9 2 15 9 2 15 13 9 13
21 3 9 13 2 9 15 2 9 2 13 2 2 3 9 13 2 13 15 9 2 9
33 15 2 3 9 9 0 0 2 0 0 13 9 9 2 1 9 0 13 9 9 2 13 15 0 2 9 0 2 2 13 2 9 13
5 13 15 9 3 9
12 15 3 13 2 7 15 9 15 15 13 13 13
6 7 9 0 0 9 13
18 9 13 7 13 13 9 9 2 15 13 2 13 2 7 0 15 9 13
40 7 16 0 9 13 13 9 2 16 9 9 13 2 15 9 9 7 3 13 7 3 1 9 13 2 3 9 1 9 13 2 3 9 0 13 7 0 13 13 9
1 13
15 13 9 13 9 0 9 2 13 9 2 15 3 13 13 3
13 13 7 9 7 9 7 9 7 0 0 0 9 9
5 15 13 2 0 13
12 13 0 9 15 0 7 3 1 15 13 9 13
3 3 13 9
3 9 2 13
18 3 9 9 2 3 9 9 2 3 9 9 13 13 9 2 9 15 0
5 9 13 15 9 13
7 0 2 3 13 2 9 13
8 3 2 13 2 13 7 9 13
3 3 13 15
5 15 13 2 13 3
16 3 9 9 2 3 15 13 9 2 3 3 9 7 9 0 13
11 13 2 0 2 13 15 13 2 7 3 13
15 15 0 9 7 9 7 9 7 0 9 13 2 9 13 9
10 1 15 15 7 13 7 13 7 13 13
5 1 15 13 9 9
17 0 3 0 13 2 0 3 0 9 0 2 1 0 15 9 9 13
16 9 9 0 13 2 7 0 1 9 13 2 7 9 13 9 15
16 0 13 0 0 9 13 1 15 9 0 13 2 3 3 13 13
24 13 9 9 2 7 0 13 13 9 9 2 7 0 13 3 13 9 9 2 7 13 9 9 13
20 7 7 3 13 3 13 9 0 9 2 7 16 13 15 9 2 13 13 9 9
11 3 9 7 9 13 15 9 0 2 15 9
21 15 3 13 9 9 9 2 0 13 7 9 13 7 9 0 13 7 9 13 9 13
23 9 13 13 15 7 13 13 9 9 13 0 9 2 13 9 2 13 2 9 16 9 9 13
7 15 3 13 2 13 13 9
7 3 9 13 9 0 13 9
26 0 13 0 9 9 2 1 9 9 2 1 9 9 13 2 9 3 3 0 0 9 13 2 9 9 13
5 13 9 0 1 15
28 15 3 9 13 2 7 13 1 9 9 13 3 13 0 1 9 9 13 0 9 2 3 9 2 9 9 13 9
4 13 3 9 9
18 15 9 2 7 16 9 0 3 13 13 2 9 13 3 2 13 2 0
14 3 13 15 9 2 15 9 2 15 0 2 9 2 9
15 15 9 0 13 2 16 0 9 9 13 7 13 0 9 9
29 9 9 3 0 9 1 9 13 7 0 13 9 2 7 3 0 13 9 13 0 9 2 15 3 0 3 13 9 9
2 13 9
12 13 3 9 9 13 7 16 9 13 13 13 9
9 13 9 9 2 0 15 3 13 9
2 13 9
30 1 15 9 1 0 13 9 0 13 9 2 7 9 0 0 13 9 9 13 7 0 9 9 13 7 9 3 16 0 13
11 15 9 2 15 9 2 15 13 0 0 9
15 1 15 13 9 1 9 9 2 9 9 13 7 9 13 9
10 13 2 7 9 13 2 7 13 1 9
5 7 15 3 13 3
7 13 13 3 7 9 0 13
45 13 1 0 13 9 15 9 7 2 6 9 9 0 7 0 0 13 15 13 9 2 13 2 13 2 9 0 9 2 2 7 9 13 9 2 2 2 16 13 7 0 9 13 0 9
33 16 0 13 9 13 9 2 9 8 9 9 9 13 2 7 7 1 9 9 2 7 15 0 0 9 9 13 2 7 15 0 9 13
3 3 13 15
3 2 13 7
23 3 0 9 7 13 9 9 13 9 2 16 9 13 0 9 9 13 7 13 9 7 13 9
28 3 0 9 13 1 9 7 9 9 9 13 0 1 0 13 9 2 3 9 15 13 2 7 7 13 13 9 13
15 7 0 9 3 13 13 2 16 15 13 3 3 13 9 9
29 15 16 9 3 13 2 2 7 15 13 2 7 15 13 2 13 2 7 13 1 9 0 13 1 9 7 9 13 13
10 9 9 13 7 13 9 9 13 15 9
4 9 3 0 13
25 9 9 9 2 16 0 2 13 2 7 7 3 7 15 7 3 7 15 13 9 2 9 3 0 13
4 13 15 0 9
2 15 13
9 0 0 13 9 2 3 13 0 13
9 9 13 15 13 3 2 3 13 9
4 13 9 13 9
13 3 0 9 13 0 9 2 9 13 7 1 9 13
7 13 15 9 2 13 1 9
8 1 9 9 2 3 13 2 13
3 9 13 13
13 16 9 9 1 0 13 2 13 7 0 13 9 9
21 9 0 7 0 13 9 2 7 1 9 9 3 3 9 13 13 0 7 0 9 13
31 15 3 0 9 16 9 13 13 2 3 13 2 15 9 13 9 2 7 13 13 9 13 9 7 13 0 7 0 13 9 13
13 7 0 16 13 1 9 9 2 13 7 15 13 13
10 9 13 2 13 7 9 15 2 15 13
14 7 15 9 13 7 13 9 7 13 13 7 15 13 13
5 13 0 13 9 9
15 9 1 9 2 15 9 1 9 13 2 9 9 13 9 13
13 13 2 2 3 15 13 13 1 0 9 2 15 9
7 15 3 13 13 9 13 0
11 1 9 3 15 9 2 3 1 9 9 13
13 0 13 0 13 9 7 13 9 13 1 9 9 13
13 15 3 9 0 9 13 2 3 13 9 13 1 0
26 8 3 9 9 9 0 9 3 13 13 7 9 13 2 15 0 9 9 13 13 2 7 9 13 13 9
14 0 9 13 9 9 7 9 0 0 13 9 7 9 9
12 15 16 13 2 0 9 9 1 9 13 1 9
12 3 7 9 13 7 13 9 2 3 9 13 13
19 15 13 2 16 9 2 1 0 9 9 2 16 13 2 13 7 13 13 9
17 13 9 7 13 9 13 13 9 9 7 0 13 13 9 13 9 13
18 15 3 13 0 13 9 7 2 16 9 13 9 9 13 2 9 3 13
15 13 3 2 7 16 13 9 3 13 2 2 15 13 9 13
17 3 9 2 9 0 1 9 2 13 2 1 9 0 0 9 0 13
3 9 9 13
17 3 3 7 9 13 15 13 7 15 9 7 0 9 7 0 9 13
21 9 3 13 9 13 7 13 13 9 2 16 3 0 15 9 2 16 3 13 0 15
3 3 3 13
34 13 9 0 9 13 15 7 9 9 13 0 0 9 13 2 2 13 9 13 7 9 13 13 1 0 9 2 16 0 0 9 1 9 13
28 3 15 9 13 9 2 3 15 13 0 13 9 2 9 2 16 8 15 3 9 13 2 9 1 9 9 13 0
15 7 16 3 13 2 13 1 9 9 13 9 0 7 0 13
16 9 0 7 9 9 9 13 2 15 15 9 15 2 13 2 13
12 7 3 0 9 9 9 1 15 13 9 13 9
11 0 13 13 9 0 13 9 7 13 9 9
11 13 3 9 7 13 9 0 13 13 9 9
23 8 3 9 2 0 13 13 9 15 9 13 0 9 2 7 9 0 13 7 13 0 9 9
20 9 2 13 2 15 1 9 9 9 13 2 13 13 2 7 12 9 9 13 3
13 13 15 7 9 0 9 9 13 7 9 9 13 13
28 3 13 7 3 9 13 9 7 0 9 7 9 13 9 9 0 7 9 1 9 0 13 7 0 1 0 13 9
7 0 0 13 2 9 2 9
39 15 3 7 13 2 13 1 9 9 13 9 7 0 0 9 2 15 13 0 2 13 1 9 9 7 9 7 9 7 0 9 1 9 13 13 7 9 13 9
23 9 15 0 13 9 9 2 13 16 9 3 2 13 2 1 2 7 2 0 13 9 2 13
6 3 15 9 9 15 13
6 7 0 13 15 13 9
14 16 13 9 13 2 9 13 15 0 7 13 15 3 13
29 13 1 9 9 2 9 13 2 13 9 0 9 2 13 9 2 13 7 9 7 9 2 7 9 1 0 13 13 9
9 1 9 9 13 9 16 9 1 15
21 7 9 9 9 13 0 13 7 13 13 2 16 9 9 13 2 7 3 9 0 13
25 3 9 0 13 0 9 2 3 9 0 13 1 9 3 13 13 9 2 7 1 9 13 9 9 13
9 13 15 9 0 7 9 9 13 9
11 13 15 9 15 7 13 13 7 3 13 13
18 7 15 2 16 3 13 0 9 13 2 13 9 0 9 7 15 13 9
21 13 7 13 0 9 9 7 1 0 7 9 9 7 9 9 13 13 0 15 9 9
17 16 9 13 2 13 15 13 15 15 2 7 13 9 9 15 0 0
9 8 7 0 0 9 13 15 13 9
8 3 13 2 9 13 9 0 0
10 16 3 13 9 2 13 7 13 1 15
28 13 3 0 1 0 9 9 0 9 7 13 9 9 2 9 0 7 13 1 9 9 0 13 7 0 13 0 9
21 13 3 0 9 2 15 13 9 0 9 2 7 3 9 0 9 3 13 2 16 9
8 15 13 13 2 3 1 15 13
19 13 3 3 13 0 9 2 7 9 3 0 9 13 3 15 13 1 9 13
5 15 3 13 13 13
25 8 7 3 9 15 2 16 13 9 9 2 1 9 13 2 3 15 9 9 2 15 0 9 0 13
17 7 3 3 15 13 15 9 13 2 7 9 0 13 9 7 13 13
4 13 3 9 0
24 16 15 3 13 9 2 2 13 9 7 15 13 13 1 15 9 13 2 7 3 3 9 9 13
18 7 3 3 13 9 16 2 9 9 13 2 1 15 9 9 9 13 13
16 13 15 9 9 13 1 9 2 7 9 3 13 1 9 9 13
4 0 13 0 13
12 3 13 9 2 7 9 13 9 9 1 9 13
15 3 9 9 13 13 2 3 9 2 7 9 1 9 0 13
21 12 3 9 1 9 15 9 13 2 2 7 16 0 13 13 2 9 15 0 13 13
23 16 3 13 2 1 9 15 0 7 0 9 13 7 3 1 9 15 3 13 2 0 9 13
22 13 15 9 3 0 7 1 9 1 9 13 2 2 1 15 9 9 13 1 15 9 13
11 15 9 1 0 9 3 13 2 13 9 12
18 1 9 7 15 13 9 0 2 0 13 9 2 7 1 9 0 9 13
13 1 9 7 9 13 0 2 1 15 9 0 13 13
11 3 15 16 0 13 2 3 13 9 0 13
26 1 9 7 13 3 3 1 9 9 9 0 7 9 13 2 1 9 13 13 7 3 13 9 13 13 9
18 13 7 0 1 9 13 2 7 15 9 0 9 13 7 9 13 9 13
12 1 13 3 3 9 13 9 1 9 13 9 13
12 3 13 9 9 13 0 7 12 9 0 9 13
10 13 3 1 9 9 9 1 9 15 13
31 3 0 9 1 9 13 2 1 15 9 13 9 0 13 7 9 9 0 7 9 0 3 0 2 1 15 9 15 13 13 13
10 13 3 9 13 2 15 1 9 9 13
9 9 7 9 13 2 7 9 0 9
4 3 13 8 13
14 15 2 3 1 9 13 2 1 15 9 0 9 9 13
28 1 15 9 7 9 0 1 9 13 2 7 0 9 1 0 9 13 2 15 0 2 16 3 13 2 15 13 9
20 12 2 7 3 9 0 9 2 0 3 13 2 0 9 9 7 9 12 9 13
11 7 15 9 0 15 0 13 2 13 9 13
24 15 13 9 16 13 1 9 13 2 13 0 1 9 2 15 1 15 9 13 13 2 2 0 9
12 1 0 3 13 2 16 1 9 15 15 9 13
21 3 16 3 13 0 9 2 9 15 13 13 1 9 7 13 13 2 16 15 9 13
10 7 3 0 13 9 0 2 1 15 13
13 13 7 15 9 9 1 9 2 15 3 13 12 9
17 13 3 0 9 7 9 1 9 9 13 13 13 2 16 9 13 9
15 0 15 13 9 7 3 3 9 15 13 13 16 9 8 9
21 9 0 0 13 2 15 15 9 0 9 15 13 2 0 1 0 2 7 3 3 13
3 15 3 13
3 13 15 15
9 1 9 2 3 13 13 15 13 9
5 9 0 9 9 13
21 3 3 13 9 0 9 1 9 0 13 7 9 13 1 9 7 9 1 0 9 13
13 7 3 1 15 3 3 0 13 9 2 7 3 13
12 15 13 13 2 7 0 9 13 2 3 9 13
16 0 9 3 3 15 0 9 13 2 7 15 15 13 13 16 13
6 13 13 3 9 3 13
14 7 3 0 13 1 15 9 2 15 9 0 9 0 13
15 13 9 0 9 2 1 15 9 9 8 13 13 7 9 9
9 9 7 13 13 9 9 7 9 13
18 13 7 9 1 9 0 13 13 2 7 1 9 0 9 1 9 0 9
19 9 7 0 13 13 9 7 1 13 9 9 0 13 9 9 3 7 3 13
19 7 16 15 3 13 9 2 0 13 9 9 0 13 7 0 9 9 13 13
29 3 3 9 0 9 13 2 9 13 3 15 0 13 1 9 13 2 7 16 3 0 9 15 13 2 0 9 15 13
4 13 3 13 9
14 13 9 1 9 0 7 0 9 2 7 13 9 0 0
11 1 9 7 0 7 0 0 7 0 13 9
35 3 16 15 0 9 9 1 9 13 2 13 3 15 9 13 13 1 9 2 1 15 9 13 0 13 1 9 9 2 0 13 13 15 13 9
17 13 3 0 9 7 9 13 13 9 13 7 13 3 0 9 13 9
14 13 1 15 9 9 9 7 9 13 9 9 9 13 13
7 13 3 2 16 3 0 13
14 13 15 9 3 3 9 13 7 9 1 9 0 13 13
14 15 3 3 13 9 0 2 7 13 15 3 1 9 13
33 3 9 15 0 9 13 13 7 13 9 0 9 2 16 15 15 3 13 9 13 2 16 3 9 9 13 7 9 3 1 9 13 13
23 0 3 9 16 9 9 13 7 9 13 13 2 13 9 7 9 13 9 7 13 3 9 13
11 13 13 9 7 9 1 0 9 9 13 13
23 3 13 0 9 0 7 0 9 2 0 13 13 15 9 1 9 13 2 7 9 13 1 9
4 9 7 9 13
8 0 1 9 9 9 13 9 13
6 3 13 0 15 9 13
10 3 7 0 9 0 15 9 9 0 13
17 3 13 13 9 0 3 13 2 15 1 9 9 13 13 1 15 9
3 6 9 13
3 0 0 13
10 3 3 3 0 13 2 7 3 0 13
23 13 3 15 7 3 9 13 9 0 13 0 3 13 2 16 9 15 9 13 1 0 9 13
18 15 16 1 9 3 7 3 13 2 7 9 0 0 9 13 2 8 13
8 3 13 0 2 16 15 13 9
7 3 13 2 16 13 13 3
9 9 9 13 13 3 3 1 9 0
5 9 3 0 13 9
19 0 7 9 12 13 9 1 9 13 2 1 15 0 7 13 9 9 13 9
9 1 9 7 9 1 9 13 9 13
6 13 9 9 9 0 9
10 7 15 3 0 9 1 0 9 9 13
13 15 16 0 1 3 0 13 9 2 13 13 9 13
4 15 13 9 9
14 15 16 13 2 1 9 12 13 13 7 0 9 9 13
22 15 9 13 3 2 3 1 0 9 2 0 7 9 9 1 9 9 13 2 16 9 13
23 13 7 1 9 9 9 12 2 1 15 9 9 8 0 13 1 9 2 15 3 1 9 13
11 13 9 9 1 9 13 7 9 0 13 13
9 3 3 7 9 3 9 0 9 13
17 13 3 9 7 1 9 13 3 13 9 2 16 13 9 9 13 13
6 13 9 3 9 0 9
3 13 2 13
22 15 13 1 15 9 3 13 9 13 2 3 13 15 2 15 1 15 13 2 15 15 13
15 7 15 2 15 3 3 9 13 2 13 15 13 15 9 13
2 9 13
33 3 13 0 15 13 2 7 13 1 15 2 16 3 0 13 2 3 13 9 13 7 13 2 15 13 9 15 2 15 3 7 3 13
12 9 13 2 9 2 9 13 2 15 9 9 13
6 7 3 2 3 15 13
11 13 15 9 0 2 13 1 9 15 9 13
12 1 9 2 0 9 16 13 15 9 13 2 13
8 15 13 15 13 2 3 0 13
9 7 15 9 13 0 3 16 3 13
11 1 9 2 15 1 15 9 1 9 9 13
8 7 7 13 7 13 15 15 13
3 0 9 13
12 9 2 9 2 9 7 9 0 16 13 2 13
8 1 9 2 3 15 0 9 13
10 9 1 9 13 2 7 15 13 1 9
11 9 0 16 9 13 2 9 1 9 13 13
10 3 7 0 15 13 2 0 1 9 13
13 3 1 15 9 13 2 16 15 1 9 9 9 13
12 7 9 3 0 13 2 15 3 1 9 13 13
3 13 3 9
8 0 3 7 0 7 0 9 13
4 0 13 9 9
6 0 7 9 15 13 13
3 3 0 13
7 13 15 15 1 9 0 13
4 3 0 0 13
3 1 9 13
6 3 13 9 0 9 13
8 15 9 13 2 16 15 9 13
9 13 3 1 9 7 3 13 15 3
6 3 3 9 15 9 13
9 9 2 9 9 1 9 0 9 13
4 15 7 9 13
11 3 15 15 9 9 13 2 3 3 15 13
3 3 13 15
8 9 0 13 3 2 7 3 13
6 15 7 9 0 3 13
9 7 9 13 2 15 9 1 15 13
2 13 7
15 9 9 3 13 2 7 16 3 9 13 13 2 9 1 9
10 7 3 0 9 13 7 7 15 3 13
2 9 13
11 0 9 1 9 13 2 16 15 1 9 13
17 13 3 9 0 2 16 13 16 9 15 13 13 2 15 9 9 13
8 9 2 9 9 9 13 9 0
5 13 3 0 9 9
16 7 3 13 13 9 2 7 0 9 9 7 9 13 9 13 13
12 15 3 13 1 9 15 9 13 15 13 0 13
3 9 13 13
14 13 2 15 13 15 9 13 13 2 15 1 9 9 13
3 15 3 13
6 13 3 3 13 9 13
13 9 0 9 3 13 2 15 15 9 1 9 13 13
13 7 15 9 0 13 13 2 16 15 9 3 13 9
19 9 15 2 1 15 12 9 13 2 1 3 15 9 13 2 7 3 13 9
22 3 15 13 15 9 2 0 9 13 2 0 9 2 9 3 0 2 9 0 7 9 0
7 0 15 9 9 13 7 9
3 13 9 9
2 3 13
5 3 0 9 9 13
5 1 9 15 13 13
13 3 0 9 13 2 7 1 9 7 1 9 9 13
7 7 9 7 3 7 3 13
13 7 3 3 3 9 1 15 13 2 16 9 0 13
6 1 9 9 13 7 0
31 13 13 15 9 2 1 15 13 13 0 9 9 2 7 3 0 2 1 15 9 9 13 0 9 13 2 0 9 0 9 13
17 3 7 0 9 1 9 13 2 3 9 13 2 9 13 13 2 13
5 7 15 3 9 13
39 3 1 13 9 3 15 9 13 2 15 0 13 2 7 0 0 2 9 0 13 7 9 13 0 2 7 13 0 9 9 9 3 13 2 1 15 9 9 13
12 13 9 1 9 13 7 15 1 9 13 9 13
9 3 16 0 15 13 13 9 2 13
10 7 13 2 15 9 15 0 0 13 9
18 3 9 1 9 13 2 15 13 1 9 7 9 7 9 1 9 13 13
18 3 15 2 15 0 13 13 2 1 0 9 13 13 2 3 9 0 13
15 16 3 0 9 13 2 13 13 15 9 0 2 15 15 13
7 3 3 15 9 0 13 13
8 3 7 9 13 7 7 9 0
14 15 9 2 16 3 0 9 15 13 2 1 9 13 13
7 3 3 3 9 1 9 13
15 13 15 9 0 7 9 0 13 2 16 13 3 1 0 13
31 16 15 13 2 9 0 2 9 7 9 13 7 3 9 2 3 9 7 9 13 2 9 9 13 7 9 9 0 0 9 13
9 1 15 9 13 9 9 13 9 13
8 9 13 9 9 7 9 0 13
4 3 9 3 13
7 3 13 15 13 13 0 9
8 13 9 9 7 13 9 3 13
7 1 15 9 9 1 9 13
9 15 9 1 9 13 13 13 9 9
11 9 3 0 16 9 13 2 9 13 9 13
6 16 13 15 2 9 13
4 7 0 9 13
4 3 15 9 13
5 3 0 9 9 13
7 9 13 2 7 3 0 13
5 9 15 1 9 13
10 13 9 9 9 7 15 13 3 3 13
14 9 7 9 13 2 9 9 13 2 7 9 0 3 13
9 7 16 9 9 13 2 9 6 13
5 7 7 3 13 13
5 13 7 3 1 9
5 3 2 3 15 13
5 13 15 1 15 13
3 9 13 13
17 0 16 9 13 2 9 3 15 9 13 2 15 3 0 13 16 9
12 12 9 9 1 9 0 3 13 2 3 9 9
4 3 13 1 0
8 9 15 13 7 3 3 0 9
8 9 7 9 0 13 16 9 9
10 3 3 13 13 2 0 9 7 9 0
10 13 13 3 13 9 16 3 15 13 9
5 9 9 0 13 13
8 3 13 7 7 16 1 9 13
5 7 0 9 9 13
5 0 13 2 9 13
2 9 13
6 15 13 2 15 15 13
5 3 13 7 3 13
4 15 13 15 13
11 1 9 13 7 13 13 9 1 9 3 13
8 3 13 2 15 13 2 16 9
11 1 9 3 15 9 13 2 15 9 0 13
10 0 9 13 2 0 2 9 7 3 9
13 9 15 0 13 2 9 9 2 9 0 7 0 9
13 7 1 9 0 9 13 2 7 13 9 15 0 9
7 13 3 9 2 0 15 13
18 7 16 15 9 13 2 9 13 2 1 15 0 13 2 16 15 13 13
15 7 15 9 2 16 9 0 13 2 0 15 9 9 9 13
6 3 13 2 15 0 13
9 13 7 0 9 2 15 15 3 13
7 15 13 13 2 3 15 13
10 3 9 9 7 1 9 15 9 9 13
8 0 13 7 2 16 9 9 13
7 7 3 13 15 9 15 13
11 7 0 13 2 9 3 13 7 0 16 9
8 13 9 3 3 7 3 0 13
8 3 3 0 13 7 0 9 9
9 7 7 13 2 15 0 7 15 13
6 15 9 13 2 15 9
8 3 15 6 3 9 9 13 13
4 7 3 9 13
4 3 9 9 13
14 9 3 13 2 15 1 9 13 2 13 15 2 13 15
4 3 9 13 13
3 15 13 13
16 9 16 9 0 13 2 9 3 15 13 2 16 15 9 13 13
5 2 7 2 13 9
13 3 13 1 9 0 2 15 9 2 9 2 3 9
6 15 15 13 2 9 13
19 1 0 7 3 0 2 3 2 8 2 13 2 2 7 3 9 13 7 0
12 16 13 3 1 9 2 3 15 9 13 3 9
14 7 3 13 3 7 7 13 2 13 15 13 15 8 13
13 7 3 0 13 2 9 0 13 2 3 0 1 15
18 3 15 9 9 1 9 13 2 9 9 15 13 2 3 13 1 0 13
5 3 9 0 13 0
7 15 9 3 13 3 9 9
15 7 3 15 13 9 12 9 2 15 15 13 9 3 9 0
14 3 3 13 2 0 1 9 9 13 2 3 0 9 13
8 3 13 2 3 13 9 12 9
10 7 16 15 9 13 2 3 3 15 13
8 3 9 13 3 9 2 3 9
19 15 1 15 13 2 3 9 0 13 2 7 16 13 15 9 2 9 0 13
15 15 7 13 13 2 16 7 7 0 7 7 9 15 9 13
12 3 0 13 2 16 15 13 0 15 1 9 13
18 3 0 13 0 9 1 9 2 13 9 2 9 0 2 7 9 9 13
4 3 3 3 13
6 7 0 13 0 3 9
11 3 0 9 0 13 2 16 15 0 3 13
2 9 13
7 13 15 13 9 9 3 13
3 0 9 13
7 15 3 3 13 2 3 13
3 3 9 13
10 3 6 9 0 13 13 2 16 9 13
9 7 13 15 9 2 7 7 15 0
9 3 13 13 13 2 3 0 9 13
10 15 16 3 13 2 13 3 9 13 13
9 7 9 0 0 9 13 7 13 0
8 7 15 7 15 13 2 15 3
15 9 0 13 13 2 1 9 2 9 1 9 2 3 9 13
3 7 13 3
10 13 13 15 9 3 2 13 15 9 3
12 3 0 13 2 3 13 9 15 2 7 3 13
19 3 9 15 13 7 9 0 7 9 9 2 15 13 13 2 16 9 0 13
7 13 9 9 1 9 7 9
5 15 13 15 15 13
8 15 9 13 2 15 13 13 13
8 9 15 9 0 13 16 9 13
10 15 7 9 13 9 9 3 0 9 9
6 15 9 13 13 9 13
4 9 9 3 13
5 9 2 9 13 0
13 3 7 13 2 13 9 2 7 7 15 7 9 13
4 7 15 15 13
15 7 13 2 15 15 9 13 13 9 2 0 9 15 7 0
9 15 16 15 13 2 13 9 0 9
6 13 13 0 9 15 13
8 7 3 2 15 15 15 9 13
11 13 9 8 3 0 2 15 16 13 2 13
4 3 0 9 13
9 13 1 9 9 2 13 15 9 0
12 0 15 9 13 0 2 15 3 15 1 9 13
7 1 9 2 0 3 13 13
12 3 1 0 9 2 13 2 13 2 3 9 0
7 9 3 2 13 2 15 13
4 7 15 15 13
8 13 2 7 15 0 13 3 13
3 9 9 13
6 13 15 2 9 2 13
4 15 15 13 0
10 3 13 0 9 2 7 3 9 9 13
6 13 15 1 9 0 13
3 15 3 13
13 15 9 15 13 2 16 1 9 13 7 13 9 0
11 3 13 2 3 16 9 15 9 9 0 13
5 13 3 3 0 13
7 7 3 15 9 13 9 0
4 3 12 9 13
7 16 13 2 13 1 9 9
12 0 13 7 0 9 2 3 16 1 9 0 13
12 15 15 3 12 9 13 2 7 13 16 9 13
8 13 3 0 9 2 7 3 13
15 13 7 0 3 3 13 2 7 0 2 15 3 13 16 13
13 3 13 9 13 9 13 2 7 15 13 2 0 13
17 13 3 3 9 15 9 0 2 16 13 15 1 9 15 1 9 13
4 13 15 9 9
4 3 15 3 13
10 16 3 13 2 3 9 1 9 3 13
8 9 9 13 2 7 9 3 13
29 3 9 13 2 16 9 13 7 13 9 9 9 13 7 9 0 13 13 15 13 9 2 9 3 9 9 15 3 13
5 7 3 9 15 13
8 13 15 3 9 7 9 1 9
7 13 3 2 0 9 15 13
8 3 1 9 15 13 2 13 9
5 9 15 3 13 13
9 15 0 13 3 0 9 13 3 13
10 13 2 9 2 15 13 15 9 0 13
16 7 3 3 1 9 0 13 13 15 15 13 2 7 9 13 13
10 3 16 15 0 13 2 9 3 13 13
10 0 13 3 13 2 16 13 15 9 13
13 9 13 9 7 9 15 2 7 3 13 0 9 9
14 7 3 3 13 15 1 0 9 2 15 13 2 9 13
13 7 9 9 13 15 13 1 15 13 1 9 3 13
10 9 7 0 2 9 7 8 9 9 13
8 0 9 3 9 9 13 13 13
19 7 3 9 13 13 2 7 3 13 9 0 0 9 13 13 2 7 0 9
4 1 0 9 13
6 13 3 13 16 3 13
25 7 9 3 9 13 1 9 9 13 2 9 7 8 1 15 9 13 7 9 13 16 3 13 2 13
5 15 15 13 0 13
22 9 9 3 13 2 7 3 15 1 9 13 2 1 0 13 15 2 15 15 3 3 13
6 13 0 13 0 7 0
16 3 13 9 9 13 2 16 16 9 13 13 2 1 0 9 13
12 15 3 16 9 3 13 2 1 9 3 9 13
10 13 3 2 16 15 13 2 9 9 0
8 3 13 9 7 13 15 9 13
11 3 9 15 13 16 13 13 2 9 3 13
7 16 13 3 13 2 9 13
31 15 7 0 16 0 13 9 2 13 13 9 15 0 2 3 12 9 9 13 2 7 1 9 9 2 3 15 9 9 9 13
7 13 15 15 9 1 9 13
2 13 15
11 3 13 9 2 16 9 1 9 0 9 13
33 13 15 9 13 7 13 2 3 9 3 0 3 3 13 13 2 0 3 3 2 16 3 0 15 9 13 13 2 16 0 3 9 13
6 13 9 15 3 13 13
3 3 6 13
1 13
9 9 13 13 8 9 7 9 3 13
1 13
12 3 13 9 2 13 9 7 1 0 9 0 13
6 13 3 9 13 7 13
2 13 13
3 13 2 13
22 15 2 0 9 2 3 13 15 13 2 7 13 1 9 9 3 13 15 13 9 13 0
4 15 13 9 13
8 3 6 15 13 2 16 9 13
21 7 3 9 2 15 13 1 9 9 3 13 16 3 0 9 13 2 3 15 15 13
14 13 9 9 9 13 7 9 9 3 7 3 0 9 13
14 7 3 9 2 1 9 9 9 13 9 1 9 13 13
17 7 3 3 9 9 13 13 7 0 9 2 7 9 1 9 13 0
8 15 16 9 3 13 2 13 9
6 9 13 15 0 0 13
11 13 2 16 1 0 9 13 15 9 9 13
3 7 15 3
10 7 3 13 13 2 3 0 0 0 13
9 15 13 7 0 2 16 15 9 13
16 7 16 15 13 0 8 2 3 3 13 2 3 3 0 13 13
5 13 15 2 15 13
8 15 13 15 0 2 3 3 13
4 3 7 0 13
11 13 3 9 15 13 9 0 2 15 3 13
17 13 3 9 13 1 0 9 2 3 13 13 9 7 15 1 9 13
6 7 15 13 9 1 9
10 3 9 1 9 13 7 9 9 3 13
13 15 13 13 15 9 9 13 2 3 3 9 15 13
2 13 3
7 16 13 2 13 15 9 8
5 1 9 3 0 13
6 13 9 0 3 3 12
14 3 9 13 9 0 2 7 9 0 13 3 16 13 13
17 13 9 12 2 15 13 9 0 0 2 3 9 9 1 9 0 13
7 15 16 13 2 9 9 13
13 1 15 13 9 3 13 15 15 13 2 16 0 13
6 7 15 3 15 13 13
9 13 2 1 15 13 2 16 13 0
8 3 3 13 1 15 9 13 9
5 15 13 1 9 13
7 7 9 3 2 9 3 13
17 13 9 13 2 7 1 0 9 2 15 13 2 15 9 13 1 9
18 3 13 9 3 13 7 3 0 0 9 13 15 13 9 0 2 16 13
2 13 15
4 9 9 3 13
10 7 13 1 9 2 16 9 1 9 13
13 2 7 2 13 2 13 3 13 9 15 3 0 9
5 9 7 3 0 13
15 1 9 0 2 15 13 9 2 9 13 9 12 2 9 12
9 13 1 9 1 9 9 12 9 0
3 9 13 0
12 1 9 13 13 2 15 13 3 13 2 9 3
7 13 9 3 15 0 9 13
21 13 9 7 15 13 15 9 13 13 2 16 1 0 9 13 2 1 9 0 13 13
14 3 7 9 9 13 7 9 9 2 15 9 7 9 13
16 3 9 9 7 13 1 9 9 1 9 9 13 7 9 9 13
9 3 9 13 9 7 9 1 9 13
4 9 7 3 13
25 9 0 7 9 13 7 9 13 1 9 7 1 0 9 9 13 2 9 3 13 13 7 9 9 13
9 13 15 0 9 7 13 0 9 13
18 16 3 9 13 13 2 7 13 15 9 13 2 7 9 0 13 3 13
33 13 9 2 8 3 3 9 2 3 1 9 3 0 2 15 3 9 13 3 13 2 7 1 0 9 9 2 16 0 13 9 0 13
12 3 15 13 2 16 15 9 1 0 15 9 13
13 7 7 3 3 13 9 15 2 15 13 13 9 13
6 8 7 3 13 9 0
25 1 9 3 9 13 9 9 2 3 9 13 0 13 2 16 15 13 13 2 0 9 13 1 9 13
16 13 15 9 2 7 3 1 0 9 0 13 2 2 0 9 13
21 3 13 9 3 13 15 9 1 9 13 7 3 9 13 7 3 3 9 13 15 13
7 15 3 13 2 1 0 13
6 7 1 15 9 9 13
7 3 13 15 9 0 2 9
8 15 0 13 0 13 2 0 0
5 9 9 9 13 9
17 0 9 13 9 13 0 13 0 0 2 9 15 0 2 15 0 9
12 3 0 13 9 0 2 16 16 13 9 1 9
13 0 13 13 9 9 0 2 3 13 0 1 9 0
10 7 9 0 2 15 9 13 7 9 13
22 3 3 9 1 9 13 2 16 9 1 9 13 13 2 7 9 1 15 13 9 9 13
9 13 13 9 2 1 15 9 13 13
4 9 0 13 13
9 9 1 9 13 13 7 9 1 9
4 9 7 9 13
4 9 7 9 13
5 9 7 9 13 13
8 9 7 9 13 7 9 9 13
2 3 13
9 9 15 13 2 15 3 13 9 0
8 15 7 0 13 7 13 3 13
10 1 9 2 16 13 15 2 13 3 13
12 3 6 13 3 13 2 7 1 0 9 9 13
1 13
4 15 13 15 13
5 3 9 9 13 9
3 9 0 13
4 7 15 9 9
3 3 3 13
11 7 3 13 15 3 13 2 16 9 9 13
8 9 1 9 13 2 9 0 13
4 9 0 9 13
3 9 13 3
8 9 15 1 9 13 13 15 13
5 9 13 2 9 13
5 12 9 13 7 9
11 9 0 13 2 16 15 1 9 15 9 13
5 12 9 1 9 13
4 9 3 13 13
9 13 2 3 13 2 16 13 3 13
11 15 7 3 0 13 2 16 1 15 3 13
10 1 0 9 13 2 1 15 9 3 13
4 15 0 0 13
2 13 15
3 15 0 13
5 3 13 2 3 13
6 15 9 0 13 16 9
7 1 9 2 15 15 3 13
3 9 12 13
9 9 3 13 2 7 0 13 7 0
7 7 9 0 1 15 9 13
5 3 9 3 13 13
11 7 13 1 9 2 15 15 9 13 3 3
4 9 15 9 13
4 15 13 0 9
7 3 3 13 3 9 1 9
17 1 15 9 9 2 15 1 9 13 2 9 3 3 13 3 3 13
21 15 16 13 9 9 2 13 9 1 9 7 15 7 13 2 7 15 13 2 9 0
8 6 9 2 13 2 9 9 13
3 3 0 13
11 3 0 9 13 2 16 15 15 9 0 13
5 3 3 15 3 13
12 3 15 13 2 7 15 9 2 15 15 3 13
19 3 15 13 2 7 3 13 9 0 2 7 16 13 2 9 0 9 3 13
12 3 2 13 15 1 0 2 9 2 3 9 9
28 7 7 3 7 7 3 3 13 2 16 9 0 1 9 9 3 13 2 7 7 15 13 2 16 6 9 0 13
11 13 2 3 15 13 9 15 0 7 9 0
5 3 2 13 1 9
14 7 15 3 15 13 2 7 3 13 2 16 9 0 13
13 9 15 13 13 2 13 2 7 15 15 0 6 13
25 3 13 9 2 0 7 0 9 2 7 0 9 13 2 9 12 13 1 9 2 1 9 2 1 9
4 13 2 13 9
11 3 13 9 0 9 13 2 16 3 9 13
2 13 15
12 13 15 2 15 1 15 13 7 1 9 3 13
7 15 1 15 13 7 0 13
5 15 13 9 0 2
11 9 13 9 10 2 7 9 10 13 0 2
3 8 12 2
25 9 9 2 15 1 9 13 13 9 13 2 0 13 16 0 13 15 9 0 13 7 15 3 13 2
17 3 1 15 15 9 1 0 13 2 1 9 13 16 0 13 13 2
16 10 7 13 1 9 2 9 7 9 9 1 9 13 0 13 2
13 3 3 15 9 0 13 1 1 10 9 13 13 2
6 9 3 13 9 15 2
18 3 13 1 9 12 15 13 0 7 3 0 2 1 15 13 15 9 2
29 16 0 9 0 13 7 15 13 2 1 15 16 9 2 1 15 0 13 2 9 13 10 9 2 15 9 0 13 2
9 7 0 13 1 9 0 9 0 2
10 7 1 0 9 0 7 10 0 9 2
12 15 3 9 15 13 0 13 2 3 0 9 2
14 3 7 15 9 2 15 9 13 2 9 15 13 0 2
41 16 0 13 9 2 0 15 9 9 13 2 1 9 0 10 3 13 2 13 3 0 15 7 15 9 2 1 15 9 13 12 8 12 2 16 0 9 2 9 13 2
20 9 7 0 0 15 0 13 15 9 1 9 0 13 2 15 3 13 9 9 2
10 3 1 9 2 0 13 9 9 13 2
15 9 7 0 15 9 13 15 13 1 0 9 7 9 15 2
13 0 7 9 7 9 0 13 9 2 16 1 13 2
9 13 3 0 9 0 13 9 9 2
5 15 7 13 9 2
9 13 3 9 13 0 9 15 0 2
8 7 1 15 9 0 9 13 2
20 7 3 1 9 9 0 9 9 13 15 13 1 9 13 2 13 2 8 12 2
18 15 1 15 13 4 2 7 1 15 13 1 9 2 16 9 13 9 2
10 7 7 0 9 9 13 13 9 9 2
21 3 15 2 7 15 9 15 13 9 10 9 2 3 15 13 1 0 9 13 10 2
9 3 7 10 9 13 10 9 9 2
11 3 3 13 9 9 1 9 16 1 9 2
19 15 7 13 12 0 13 7 15 13 16 9 2 15 9 13 2 9 13 2
21 3 16 0 13 9 0 1 0 9 13 7 15 13 2 3 15 13 9 0 13 2
13 13 3 1 9 9 0 0 9 1 9 13 13 2
22 3 9 0 2 15 0 13 9 2 13 13 2 15 13 1 13 2 9 13 9 10 2
45 7 9 1 9 13 2 15 13 1 13 2 7 9 10 13 0 2 1 15 9 1 0 9 13 2 15 9 0 13 2 15 3 9 13 2 3 7 9 0 15 9 15 9 13 2
8 15 13 1 15 9 9 9 2
16 1 10 0 9 9 9 9 13 9 2 0 2 0 7 0 2
31 9 3 2 16 16 9 9 9 13 2 3 0 9 3 15 9 13 3 0 13 2 0 9 15 1 9 13 2 8 12 2
19 0 7 13 16 1 15 9 0 1 0 9 13 2 15 10 1 9 13 2
16 3 2 16 9 9 13 9 2 9 9 0 9 1 9 13 2
23 1 15 8 12 13 16 9 0 9 13 9 2 15 15 13 4 2 13 4 0 9 9 2
12 0 7 13 16 1 15 9 1 9 9 13 2
11 9 3 9 13 1 9 0 2 8 12 2
22 0 7 13 16 3 13 9 9 15 7 9 0 15 2 7 9 7 9 2 8 12 2
34 13 3 1 0 9 9 0 9 13 2 16 0 9 13 2 13 10 9 13 9 15 9 0 13 2 1 10 9 13 2 9 13 0 2
28 16 3 9 9 13 2 15 15 7 0 9 10 9 13 15 9 0 13 2 16 15 10 9 10 7 9 13 2
11 1 0 7 9 0 13 13 2 1 12 2
25 0 2 16 3 3 13 15 13 0 13 13 0 16 1 15 15 13 13 9 13 1 15 9 13 2
32 15 3 9 13 4 0 9 1 9 9 0 15 9 13 13 16 7 15 0 13 2 7 3 1 0 13 7 1 15 9 13 2
38 0 2 16 15 15 2 16 9 7 0 2 3 13 15 1 9 15 9 2 1 15 13 13 2 16 1 0 13 13 1 0 9 2 1 0 1 0 2
5 15 0 15 13 2
13 3 0 13 1 0 9 13 2 15 10 13 13 2
8 15 3 1 9 0 13 13 2
12 3 7 9 15 13 13 15 9 1 15 13 2
10 7 3 0 9 2 9 0 9 13 2
8 15 9 13 0 0 9 13 2
10 16 0 3 10 9 13 9 13 15 2
38 13 7 9 13 3 1 15 9 13 13 2 3 9 9 13 2 16 1 9 2 0 9 9 13 2 0 13 0 13 15 9 13 0 1 9 13 13 2
12 13 7 1 15 15 1 9 13 0 9 9 2
20 15 3 0 13 1 9 15 10 9 0 9 13 2 16 9 13 0 7 12 2
24 15 0 13 1 15 3 9 0 13 13 2 16 13 9 13 2 9 13 12 2 7 15 3 2
13 15 3 9 0 1 9 13 2 13 0 9 9 2
16 16 7 13 15 0 0 15 0 9 3 13 9 2 0 13 2
30 1 3 9 15 9 15 1 15 9 9 13 2 13 9 9 15 2 15 16 2 1 9 9 9 9 13 15 15 13 2
18 13 16 1 9 15 9 9 13 2 13 9 15 15 1 9 15 13 2
24 3 16 9 0 2 15 9 9 13 2 13 9 7 0 2 15 0 15 9 9 0 9 13 2
8 15 3 15 1 9 3 13 2
13 3 1 9 15 13 9 0 0 9 13 3 13 2
14 1 9 10 2 1 9 0 9 2 9 1 9 13 2
23 7 3 15 15 1 9 3 13 2 3 13 0 9 13 2 16 15 1 0 15 9 13 2
18 0 7 1 15 13 9 10 3 13 16 1 15 0 9 13 15 13 2
8 1 13 9 9 9 3 13 2
25 13 3 1 0 9 10 1 0 9 16 13 1 9 16 13 2 7 15 3 15 13 13 0 9 2
11 13 3 15 0 0 15 0 9 13 0 2
9 15 0 15 3 9 0 9 13 2
9 3 1 9 9 15 0 13 13 2
26 12 3 15 12 15 9 15 9 0 13 2 15 15 9 13 13 2 0 13 15 15 3 13 3 13 2
14 16 13 1 0 2 15 15 9 9 0 9 13 13 2
15 9 7 9 0 13 9 0 16 9 0 9 9 0 9 2
14 16 15 9 1 9 0 9 13 2 15 0 9 13 2
10 13 3 9 9 1 0 9 16 9 2
32 3 15 9 9 2 1 15 1 9 9 13 0 9 2 13 0 9 0 7 3 15 9 2 1 15 9 0 1 9 9 13 2
10 0 0 9 0 13 0 16 0 0 2
28 15 3 9 0 10 9 9 10 13 2 7 3 9 1 15 13 15 13 2 7 10 13 15 1 15 0 13 2
31 3 7 0 9 9 1 9 13 15 13 2 16 7 15 9 9 2 1 15 1 9 9 13 2 13 9 9 9 3 13 2
15 3 3 10 15 1 15 9 13 2 9 0 9 13 13 2
15 7 1 10 15 9 10 0 9 13 2 0 9 13 13 2
51 16 3 0 9 13 9 15 15 15 1 9 13 0 13 13 1 15 16 15 13 3 13 2 3 2 7 0 0 2 0 9 13 9 16 15 15 0 9 9 13 0 13 13 1 15 16 9 13 3 13 2
13 3 15 0 13 1 9 15 1 9 13 3 13 2
20 9 3 0 0 9 13 2 15 9 15 9 13 9 9 1 0 13 3 13 2
14 0 3 0 15 13 9 10 0 0 9 13 3 13 2
32 15 3 13 9 9 2 15 1 12 8 13 16 9 10 15 13 1 0 9 2 15 13 0 1 9 2 16 9 9 1 9 2
8 15 3 9 0 9 9 13 2
5 13 3 9 12 2
12 3 9 9 13 2 7 0 1 1 9 13 2
3 7 12 2
9 6 2 9 0 2 13 9 10 2
5 7 12 8 12 2
4 1 9 13 2
27 3 3 10 15 1 9 13 2 16 9 13 3 13 2 3 3 0 13 13 2 16 9 7 0 0 13 2
13 16 9 0 1 15 0 9 13 13 9 13 13 2
30 0 3 9 0 0 13 2 12 1 15 9 9 13 13 2 15 15 10 9 0 9 13 2 15 13 0 9 13 13 2
14 15 7 1 15 0 13 13 15 9 9 0 13 13 2
19 16 9 15 13 2 1 15 9 13 13 2 3 15 0 9 13 13 4 2
12 13 7 12 9 16 3 9 3 9 13 13 2
9 12 13 16 0 9 9 9 13 2
17 1 9 3 0 9 2 15 13 9 9 2 0 13 12 1 9 2
15 15 16 1 9 9 2 1 15 0 0 13 0 1 13 2
20 3 15 9 1 15 13 13 16 0 9 0 9 13 2 15 1 13 9 13 2
7 15 0 13 9 9 0 2
33 13 3 13 1 9 15 15 0 13 13 2 15 15 9 1 9 0 9 3 13 13 16 1 0 9 0 9 13 2 3 9 9 2
5 15 7 13 9 2
15 1 9 3 15 15 1 9 9 13 13 2 0 13 13 2
10 1 3 15 9 9 1 9 9 13 2
16 1 15 0 2 15 1 0 13 2 1 9 9 0 13 13 2
15 3 3 3 16 1 0 9 9 1 13 9 9 13 13 2
19 15 3 9 0 13 13 1 9 9 2 15 3 9 9 0 9 13 9 2
18 0 9 13 16 15 15 1 13 9 9 13 2 3 1 0 9 13 2
22 7 1 15 9 9 2 1 15 13 1 9 9 3 16 1 0 9 9 0 0 13 2
11 7 3 1 0 15 13 2 16 13 4 2
38 7 3 1 15 16 9 9 2 16 0 9 9 9 13 2 3 13 0 1 3 9 9 9 2 7 1 13 13 0 7 13 2 16 13 1 12 8 2
19 13 3 0 9 2 16 0 9 9 1 9 13 13 2 1 0 9 9 2
25 1 9 9 2 15 9 0 9 7 0 13 2 3 16 15 0 2 7 15 3 1 9 9 13 2
22 0 9 13 16 9 9 0 10 9 13 2 1 9 9 10 1 13 2 7 9 9 2
19 7 3 1 0 1 9 13 15 15 4 3 0 13 2 16 9 9 13 2
13 7 0 1 13 1 0 15 0 13 2 0 13 2
29 1 0 3 0 15 13 2 13 3 15 0 2 15 3 13 2 7 15 0 7 0 9 13 2 15 3 9 13 2
17 7 3 13 1 9 9 13 9 7 0 9 1 9 0 9 13 2
17 0 3 0 13 9 16 15 3 15 9 13 13 2 9 13 13 2
16 16 3 10 1 0 13 0 9 0 13 7 1 9 7 9 2
7 15 13 15 8 12 13 2
17 3 3 13 16 7 9 13 1 9 9 10 2 9 13 13 9 2
4 7 9 12 2
8 13 0 9 10 13 1 9 2
13 16 15 15 9 13 3 13 13 9 13 9 13 2
26 13 7 15 3 3 13 9 1 13 13 15 15 9 13 3 13 1 0 9 15 1 9 10 9 13 2
17 7 3 13 13 16 0 13 9 0 13 13 3 15 15 9 13 2
13 15 3 9 7 9 1 15 13 16 13 15 13 2
57 16 3 1 9 9 16 13 1 0 9 13 0 9 2 9 1 0 9 13 2 16 1 13 13 2 13 9 13 1 15 9 16 9 10 1 0 13 13 2 16 3 13 15 13 2 7 9 13 1 15 15 15 9 0 9 13 2
15 7 15 0 0 9 13 2 15 0 9 0 7 0 13 2
10 3 7 1 15 0 0 9 13 13 2
17 9 7 0 2 15 0 13 13 2 0 13 15 0 9 9 13 2
39 1 3 15 9 9 9 13 2 1 15 16 9 1 0 9 1 9 13 2 13 13 15 9 15 0 0 2 15 9 0 0 15 13 0 7 0 9 13 2
15 13 3 0 3 9 1 13 9 13 1 9 9 0 13 2
22 3 3 0 9 0 13 16 15 13 13 1 10 15 15 1 9 13 1 9 0 13 2
14 15 16 0 9 9 0 9 13 2 16 1 13 4 2
27 1 15 3 16 9 1 9 15 13 15 9 13 2 13 1 9 9 16 9 13 15 1 15 15 13 13 2
15 15 3 9 3 13 2 3 9 9 2 15 13 9 9 2
34 13 3 15 3 1 10 9 13 16 15 9 9 15 13 10 9 13 13 2 13 3 15 13 0 15 15 13 7 0 15 15 3 13 2
26 16 3 1 15 9 0 9 13 1 0 9 9 13 2 0 13 9 13 15 0 15 3 9 15 13 2
11 13 3 15 9 1 9 9 1 12 8 2
24 1 3 9 15 9 13 0 9 13 7 0 9 9 13 2 13 13 0 13 9 7 0 0 2
16 1 15 9 13 16 9 13 15 1 0 7 0 13 3 13 2
34 3 1 12 1 8 13 2 16 2 16 9 13 15 1 9 0 13 2 3 15 0 13 3 13 7 13 10 9 15 1 9 9 13 2
28 13 3 1 12 8 7 8 16 1 1 9 0 9 13 13 0 7 0 9 2 13 9 16 0 13 9 15 2
16 1 15 10 13 16 1 9 0 15 0 9 0 9 9 13 2
28 7 3 2 16 15 15 1 9 13 9 0 0 13 3 13 2 3 0 15 9 13 16 3 15 15 13 9 2
6 7 3 13 8 12 2
8 0 1 9 9 13 4 15 2
13 7 12 8 12 15 13 9 15 13 16 9 9 2
8 15 7 13 9 1 9 10 2
14 16 13 15 15 13 9 3 13 9 16 1 9 13 2
29 3 7 9 2 15 9 0 9 3 13 2 9 13 3 0 13 2 3 0 9 13 2 16 12 8 12 2 13 2
19 15 3 0 9 9 15 0 9 2 15 10 0 13 2 13 4 9 13 2
31 15 15 9 7 9 7 9 9 2 13 9 13 2 16 1 13 15 15 0 9 13 2 9 0 13 15 15 9 13 9 2
14 3 1 0 9 9 2 13 9 2 0 9 0 9 2
28 7 2 15 13 0 2 0 9 9 2 16 9 7 0 2 9 9 0 13 2 0 9 7 9 1 9 13 2
60 15 13 2 13 9 9 2 3 9 9 2 3 9 9 2 7 2 15 13 0 2 1 9 9 2 0 9 3 0 0 2 7 0 9 2 1 9 0 13 2 1 15 10 0 9 13 13 2 9 9 13 7 10 15 1 9 13 13 13 2
24 15 9 0 13 7 0 9 13 2 7 0 0 9 9 2 16 2 13 0 2 0 0 13 2
44 15 7 3 3 7 1 9 2 7 1 0 9 13 4 2 0 13 1 15 16 15 15 13 9 0 1 9 13 9 2 15 9 1 15 1 9 13 2 3 10 9 9 13 2
40 15 3 9 9 13 8 12 15 2 3 0 9 2 1 9 13 13 1 9 2 1 15 15 13 1 15 13 4 2 13 9 9 7 9 7 0 9 0 9 2
15 15 7 3 0 9 9 1 9 0 9 0 13 13 9 2
15 16 15 0 13 0 3 13 2 1 1 10 9 13 0 2
35 13 3 10 9 0 16 1 13 3 0 2 7 1 13 3 0 2 7 1 13 3 9 2 9 1 0 9 13 4 1 0 7 0 9 2
18 16 3 13 9 3 10 9 2 1 9 9 2 1 0 10 9 13 2
10 15 0 15 9 9 13 13 9 0 2
19 16 13 1 9 15 0 9 13 2 1 15 9 0 9 13 2 9 13 2
21 13 3 13 13 0 2 9 0 9 13 2 1 15 1 9 13 1 0 9 13 2
18 9 3 9 3 13 16 15 1 0 1 15 0 13 0 9 13 13 2
12 16 0 0 15 13 0 9 7 0 9 13 2
31 9 3 3 13 0 13 2 15 0 0 9 13 9 13 2 16 9 0 15 3 13 13 16 0 2 13 9 9 0 13 2
17 7 13 15 1 9 9 13 2 15 9 3 9 7 9 3 13 2
17 15 3 3 15 0 2 1 9 0 7 0 13 2 1 9 13 2
24 7 9 0 1 9 13 2 10 9 0 3 0 2 1 15 9 15 9 9 1 10 9 13 2
10 15 3 0 9 13 9 15 9 13 2
19 16 0 3 10 0 7 0 9 9 0 9 13 2 16 13 15 9 13 2
20 3 0 9 9 0 7 0 9 10 0 3 13 13 2 16 1 15 9 13 2
11 7 3 13 16 15 9 9 13 0 13 2
9 16 9 9 0 3 13 9 9 2
26 16 7 13 9 9 0 0 9 9 13 2 15 3 15 9 0 13 13 2 15 9 0 13 3 13 2
12 15 3 15 0 9 13 13 2 0 13 13 2
10 1 3 16 7 13 0 13 0 13 2
19 7 15 15 9 13 2 1 3 0 0 13 4 2 9 13 13 13 0 2
31 16 3 0 0 0 0 13 2 16 1 15 9 13 0 13 2 0 13 15 9 15 9 0 13 2 13 9 9 0 13 2
2 3 2
14 15 15 15 13 1 9 9 1 13 2 9 9 13 2
11 16 13 13 2 15 1 9 9 13 13 2
10 9 7 0 13 9 15 0 4 13 2
8 1 15 9 13 10 9 9 2
8 15 3 9 3 0 9 13 2
11 15 3 9 3 0 13 2 0 9 13 2
7 3 3 1 9 13 13 2
17 15 3 15 1 9 0 1 9 13 2 3 13 0 9 13 0 2
2 3 2
13 0 9 9 10 13 2 16 1 0 9 13 13 2
18 16 3 0 9 15 1 9 13 2 1 15 1 9 9 10 9 13 2
7 15 1 9 13 3 13 2
2 0 2
11 15 15 13 0 13 3 13 2 9 13 2
9 0 7 9 3 15 13 3 13 2
14 3 3 1 9 0 15 9 7 9 9 1 9 13 2
8 7 3 9 13 2 8 12 2
11 1 13 9 1 9 10 7 1 9 10 2
8 15 13 9 9 2 15 13 2
11 7 16 13 9 2 1 15 13 3 0 2
5 15 13 3 13 2
16 15 3 9 9 13 2 15 1 12 1 8 1 8 13 3 2
18 15 15 9 13 2 9 0 7 9 0 7 0 15 9 13 13 13 2
25 1 15 0 13 2 15 9 1 9 9 13 2 15 1 9 0 9 13 1 15 13 3 0 13 2
14 3 7 9 9 13 2 7 7 13 9 0 7 0 2
8 7 3 1 15 13 9 13 2
9 15 15 13 0 9 1 9 9 2
37 13 3 13 16 9 3 0 2 1 15 0 9 9 9 13 2 0 9 1 15 0 9 13 2 3 3 0 16 1 13 15 9 9 3 0 13 2
15 13 3 9 10 9 10 9 9 2 1 9 13 15 0 2
10 3 3 9 1 9 9 9 3 13 2
45 0 3 9 1 13 9 9 2 15 0 13 0 9 13 13 13 2 3 15 13 16 1 15 13 15 9 13 2 15 3 3 13 1 15 16 13 9 3 0 7 1 15 13 13 2
23 0 3 13 16 1 3 9 2 15 0 2 15 9 0 13 2 16 13 13 7 13 9 2
20 16 1 9 9 3 0 7 0 9 15 13 13 0 13 2 16 1 13 13 2
20 15 3 9 9 9 13 2 15 3 13 1 9 1 8 2 13 1 3 9 2
8 15 13 13 2 13 2 13 2
9 16 3 13 13 2 13 3 13 2
16 15 3 0 0 13 2 16 3 13 3 2 3 3 13 13 2
21 7 16 15 13 1 15 9 2 7 0 0 9 3 15 13 2 0 9 13 13 2
5 7 13 0 13 2
9 1 9 7 9 13 1 15 9 2
20 1 13 3 0 13 0 9 1 0 9 0 13 13 2 7 1 9 0 13 2
15 1 15 12 9 9 13 13 2 15 0 10 9 13 9 2
19 13 7 0 9 0 2 3 1 9 15 9 2 15 13 12 7 0 9 2
14 7 1 9 9 10 2 15 1 0 13 9 15 13 2
17 1 0 3 9 9 1 9 0 2 15 9 13 13 2 13 13 2
22 7 16 15 9 1 0 9 13 3 13 2 3 13 13 1 15 9 16 9 9 13 2
12 7 16 15 9 2 15 1 9 13 2 13 2
14 1 9 9 9 0 0 13 3 13 2 16 13 4 2
16 0 0 9 13 9 1 3 9 13 1 9 9 0 13 9 2
13 15 3 1 9 0 13 2 3 13 16 9 13 2
24 13 3 1 3 9 13 9 15 0 13 2 1 0 3 9 7 0 2 3 7 1 9 13 2
22 16 15 9 9 15 3 1 10 9 13 2 16 13 15 1 3 0 9 9 9 13 2
41 9 3 13 13 13 2 0 13 1 9 15 9 15 9 13 7 9 13 2 13 9 0 7 0 2 15 15 1 9 9 7 0 13 1 15 9 13 7 9 13 2
37 3 2 16 1 0 1 0 0 13 9 2 1 15 9 9 13 15 9 13 2 13 9 9 7 9 0 7 9 2 3 9 13 2 9 9 13 2
28 13 3 15 1 9 9 13 15 15 1 9 9 0 13 13 2 0 2 13 9 1 15 15 9 1 15 13 2
10 0 2 0 2 1 9 9 1 15 2
13 0 2 7 2 1 9 9 1 15 16 1 9 2
26 1 15 0 15 1 9 1 15 13 13 2 13 13 2 3 15 9 0 9 2 9 15 13 9 13 2
11 15 3 13 2 10 9 1 9 0 13 2
15 1 9 13 16 9 13 13 3 13 1 13 1 15 13 2
42 15 7 9 15 15 13 1 13 9 13 2 0 3 15 13 2 15 13 16 9 13 1 15 13 13 2 3 16 15 0 13 3 13 2 7 3 9 13 13 3 13 2
6 15 3 13 1 15 2
13 15 3 1 15 13 13 13 15 3 13 9 13 2
21 16 2 13 15 13 15 7 15 13 9 2 3 13 16 10 15 13 0 10 9 2
9 3 7 13 15 16 13 9 13 2
11 3 9 9 13 15 15 0 13 3 13 2
14 15 7 1 9 13 1 15 15 13 7 13 9 9 2
10 16 3 3 1 9 3 9 13 13 2
7 7 13 1 9 0 13 2
17 3 15 1 9 7 9 13 2 0 13 15 15 1 0 9 13 2
10 9 7 15 13 0 15 9 9 13 2
17 3 13 16 9 13 1 15 13 13 2 3 1 15 9 9 0 2
2 3 2
13 13 3 13 16 15 13 15 3 13 13 3 13 2
11 15 0 13 0 15 15 13 13 3 13 2
15 3 3 9 15 0 13 13 2 16 15 13 13 3 13 2
6 15 13 1 9 9 2
9 13 16 9 13 1 15 13 13 2
2 3 2
18 9 15 13 13 13 1 15 15 1 15 13 2 16 2 9 13 9 2
14 7 15 9 1 9 9 13 2 16 2 9 13 0 2
36 1 9 7 15 1 15 13 2 16 1 13 2 16 10 9 13 10 9 2 7 16 15 13 15 13 1 9 15 13 2 7 1 9 16 13 2
21 3 3 1 13 2 9 13 2 9 7 13 15 9 2 7 3 1 9 9 13 2
9 7 3 9 13 1 15 13 13 2
2 0 2
9 15 0 13 13 2 1 15 13 2
9 3 3 1 15 13 9 9 13 2
7 7 9 13 0 13 13 2
16 1 1 9 0 9 9 13 16 1 0 9 2 16 1 13 2
8 13 3 1 15 13 9 13 2
2 3 2
11 15 1 15 13 13 13 15 10 15 13 2
5 9 7 3 13 2
19 16 3 9 9 9 13 10 0 9 2 3 0 9 10 0 9 9 13 2
10 1 13 1 15 0 0 9 0 13 2
10 13 3 16 9 13 1 15 13 13 2
21 1 15 3 7 0 15 13 9 13 3 1 15 13 13 16 0 9 13 3 13 2
8 9 13 9 7 9 9 13 2
5 13 7 9 13 2
15 9 3 1 9 15 1 9 13 4 9 9 13 7 13 2
14 9 7 2 7 0 15 13 1 9 2 9 9 13 2
23 1 15 13 16 15 15 1 9 9 13 2 3 0 13 7 16 13 0 7 1 15 13 2
24 9 0 13 1 15 16 3 13 15 13 13 1 15 0 2 7 15 13 1 15 1 15 13 2
10 3 0 3 9 13 1 15 13 13 2
11 1 15 15 16 9 13 2 13 10 9 2
17 7 16 15 15 16 9 13 9 13 3 13 2 13 0 1 15 2
14 16 10 15 10 9 0 13 2 1 15 13 13 0 2
13 15 7 15 9 15 9 3 13 2 13 13 0 2
26 7 3 13 16 1 15 15 13 13 9 2 10 9 15 13 16 9 9 1 9 2 16 12 8 13 2
21 7 13 16 3 2 13 15 9 9 9 2 9 13 13 13 2 16 0 9 13 2
24 0 3 2 16 3 10 13 13 2 3 13 9 13 2 16 9 13 15 15 0 13 3 13 2
9 1 0 0 9 15 13 9 13 2
17 7 3 1 9 15 9 9 2 15 9 13 2 15 3 13 13 2
33 3 16 2 13 16 1 10 1 15 9 9 13 15 15 0 13 3 13 2 3 0 13 15 13 15 0 13 3 13 1 9 9 2
12 15 3 9 0 13 13 9 2 7 9 9 2
20 1 15 7 16 9 13 15 13 15 9 9 2 3 13 9 13 16 1 9 2
14 3 7 13 15 15 0 13 3 13 13 16 1 9 2
17 7 1 15 3 13 16 13 15 1 9 9 15 0 13 3 13 2
10 7 3 15 9 13 13 9 3 13 2
32 3 3 9 13 15 13 7 1 9 7 1 9 15 0 13 13 2 16 15 15 13 13 15 15 0 13 3 13 1 9 9 2
20 7 3 13 2 16 0 9 13 2 9 13 15 0 13 16 13 13 3 13 2
24 3 16 13 13 3 13 2 3 1 9 15 9 13 7 9 2 1 10 9 13 1 15 0 2
28 7 1 9 10 9 2 15 15 13 3 13 1 15 2 7 1 9 15 2 7 3 1 13 15 9 13 13 2
7 1 15 3 0 9 13 2
35 3 16 15 1 15 13 13 16 15 10 9 13 0 2 3 13 15 0 9 1 15 13 13 9 13 2 1 15 16 10 9 13 10 9 2
22 7 16 15 9 13 3 13 2 1 15 9 13 3 1 15 2 7 1 15 9 13 2
6 1 0 3 13 9 2
11 3 3 9 0 9 13 16 0 15 13 2
17 13 7 15 9 0 16 13 0 9 2 15 13 15 9 0 9 2
19 3 3 3 13 16 9 15 1 15 13 13 0 13 9 2 7 9 15 2
16 3 13 16 1 15 9 1 9 13 1 9 15 9 13 13 2
8 1 0 3 1 0 13 9 2
26 3 9 13 3 15 10 13 2 3 3 16 15 3 13 16 15 13 2 16 1 9 1 15 13 13 2
11 7 16 1 15 9 10 13 1 15 9 2
14 1 9 13 16 9 13 13 3 13 7 0 9 13 2
20 13 7 15 15 9 13 9 0 2 1 15 3 0 13 9 13 13 9 13 2
21 13 3 16 9 13 3 13 1 9 13 2 7 1 0 9 9 7 9 4 13 2
18 1 15 7 13 13 4 15 1 9 9 15 15 13 1 13 9 13 2
38 13 3 15 9 9 15 0 15 13 1 15 9 9 2 15 13 1 9 15 13 9 7 9 2 3 15 15 13 1 15 13 2 7 1 9 16 13 2
13 9 7 9 13 3 13 16 13 1 9 15 13 2
10 3 7 9 13 13 13 16 9 13 2
2 3 2
17 16 9 1 13 16 13 2 1 9 9 2 13 13 15 13 9 2
15 9 0 13 1 9 13 9 2 1 9 2 1 12 8 2
15 15 13 9 1 13 9 13 2 13 0 9 7 9 9 2
2 3 2
26 16 9 9 1 9 9 9 13 2 16 1 0 13 2 15 15 10 9 7 0 13 2 13 0 13 2
6 3 7 13 9 13 2
4 13 3 0 2
19 15 7 9 9 15 13 2 7 1 9 9 2 15 1 9 9 13 13 2
6 7 1 15 9 9 2
25 3 2 16 3 13 15 0 9 1 9 0 2 3 13 15 9 1 0 2 16 13 1 12 8 2
12 7 1 9 9 2 15 9 13 13 13 4 2
9 7 3 0 9 13 2 8 12 2
10 0 9 1 15 15 13 4 13 13 2
19 7 15 13 13 2 16 1 9 15 13 9 7 9 2 16 0 9 13 2
22 3 15 13 1 9 15 9 1 15 13 2 15 15 15 13 0 13 2 16 15 9 2
10 3 7 13 1 9 15 13 9 9 2
25 3 3 13 9 1 9 13 2 16 1 9 0 9 10 13 3 9 1 9 13 15 13 9 13 2
23 1 9 7 15 13 9 13 2 3 13 13 1 0 0 9 7 9 2 16 0 9 13 2
14 7 9 9 13 1 0 9 2 16 13 1 9 16 2
10 7 1 3 9 13 9 15 9 9 2
22 3 10 0 9 13 7 1 9 9 0 1 15 2 7 1 15 9 9 1 10 9 2
30 13 3 1 15 16 2 16 9 0 10 7 9 13 2 15 3 9 2 1 15 9 13 1 13 9 13 2 0 13 2
15 7 3 10 9 9 1 9 13 3 1 15 15 9 13 2
6 9 1 13 9 13 2
26 13 3 16 3 13 0 13 1 13 9 13 2 13 1 13 9 15 3 9 7 9 0 9 13 13 2
12 0 7 13 9 15 9 13 1 13 9 13 2
10 15 15 13 13 1 9 9 12 9 2
5 15 0 15 13 2
8 10 15 13 2 1 15 13 2
9 13 7 9 15 13 2 16 9 2
5 3 15 13 13 2
9 7 3 15 13 13 2 7 3 2
16 16 3 13 2 3 13 13 2 16 0 13 13 15 13 0 2
5 7 15 13 9 2
10 16 7 13 2 3 1 15 13 13 2
7 7 3 13 13 1 0 2
8 7 13 13 1 15 13 0 2
7 7 3 13 13 1 0 2
9 3 0 13 13 15 0 13 0 2
9 1 15 7 9 13 12 9 13 2
9 3 2 16 10 13 13 1 15 2
12 7 16 1 13 7 13 3 13 13 1 0 2
7 15 0 13 9 12 9 2
4 0 2 3 2
14 16 15 13 15 2 13 16 1 15 13 9 9 10 2
7 15 2 0 1 15 13 2
7 13 3 16 4 0 13 2
20 3 16 13 9 15 15 2 7 3 9 10 9 2 16 13 9 1 9 9 2
18 3 3 15 3 13 1 15 2 7 10 9 2 7 12 9 1 15 2
10 13 3 15 13 0 2 7 13 9 2
13 1 10 15 13 13 0 2 16 13 1 12 8 2
5 15 13 3 13 2
11 15 15 1 15 13 13 2 4 0 13 2
11 3 1 9 12 9 15 2 13 9 15 2
28 16 3 2 13 12 9 2 15 9 15 13 2 3 15 15 3 4 0 13 2 7 9 15 15 13 15 13 2
11 15 7 15 13 13 15 2 13 1 15 2
16 15 3 9 1 9 13 15 2 13 16 9 1 9 15 13 2
7 7 3 3 13 1 15 2
13 3 15 15 13 1 15 13 2 3 13 1 15 2
11 0 13 3 10 15 13 2 1 15 13 2
21 7 13 15 9 16 9 15 13 13 16 15 15 13 13 15 2 9 3 13 13 2
13 7 3 16 9 3 13 13 7 13 16 1 9 2
4 16 9 13 2
31 16 9 9 1 15 13 2 16 2 16 15 15 13 0 7 1 15 2 3 9 9 2 13 16 10 13 3 13 1 15 2
14 13 7 15 0 2 16 7 15 9 2 13 1 9 2
11 7 3 3 13 15 13 0 7 1 15 2
18 3 13 3 1 9 9 13 16 13 9 13 15 13 16 15 0 0 2
17 7 13 15 0 13 0 2 16 2 16 13 9 2 16 13 15 2
11 15 3 13 13 0 3 16 13 13 0 2
14 16 15 0 13 0 2 16 9 13 9 2 13 0 2
8 0 2 13 1 9 2 3 2
11 10 15 13 1 9 2 3 13 1 15 2
6 13 3 1 9 15 2
7 0 7 15 13 1 9 2
4 16 0 13 2
19 7 15 13 1 9 16 1 15 13 2 16 9 2 15 13 1 9 13 2
11 7 3 15 13 1 9 16 0 7 0 2
9 16 15 13 1 13 7 13 13 2
14 10 7 15 13 2 7 13 1 15 2 7 1 9 2
13 7 16 1 15 2 7 1 9 2 7 1 9 2
22 7 15 2 7 13 1 15 2 16 9 2 7 3 13 1 15 2 16 0 7 0 2
9 3 10 15 13 2 1 15 13 2
5 0 2 13 3 2
10 15 15 13 3 9 7 9 9 15 2
12 7 10 15 13 2 16 3 2 13 1 9 2
11 16 9 13 9 13 1 9 1 16 3 2
11 10 7 15 13 13 1 9 2 16 3 2
10 16 15 13 16 1 16 13 1 9 2
10 3 15 13 9 15 9 13 7 13 2
6 7 3 15 13 15 2
17 13 7 16 9 15 13 10 13 13 2 0 13 9 9 16 9 2
16 9 3 0 13 9 1 16 13 9 13 1 9 1 16 3 2
14 15 3 13 16 0 7 9 2 16 13 1 12 8 2
9 1 9 7 13 15 3 13 9 2
16 13 3 9 1 15 9 2 3 16 13 7 13 13 15 13 2
11 15 3 9 13 9 13 1 12 1 9 2
17 1 15 3 13 0 13 15 13 16 13 15 7 13 7 13 15 2
8 15 1 15 3 13 9 9 2
14 15 3 13 13 1 15 0 15 13 15 2 1 9 2
12 7 13 1 0 15 3 13 0 2 1 9 2
20 15 7 9 2 3 16 1 13 7 13 3 13 13 1 0 2 13 12 9 2
5 15 0 15 13 2
16 16 1 9 7 13 13 1 0 2 13 10 3 0 9 13 2
15 16 10 15 13 13 0 7 9 2 16 13 1 12 8 2
12 10 7 9 15 13 13 2 3 16 13 13 2
11 3 10 15 0 3 13 16 12 15 13 2
12 7 12 15 2 1 13 13 2 13 9 13 2
8 3 10 15 0 13 9 13 2
5 15 7 13 0 2
12 3 0 13 16 1 9 7 13 13 1 0 2
14 16 7 13 0 16 0 13 13 9 13 2 3 13 2
7 13 7 13 13 3 13 2
8 16 13 13 1 0 9 9 2
12 7 9 3 13 3 13 16 1 9 7 9 2
25 1 3 10 13 13 7 13 13 9 2 16 13 4 2 13 16 13 3 12 0 1 9 7 9 2
8 7 3 12 0 13 9 13 2
10 15 13 0 2 16 13 1 12 9 2
8 0 9 1 15 13 15 13 2
36 1 13 7 13 13 2 15 3 12 1 9 1 15 13 2 15 0 13 13 2 16 2 13 0 13 7 13 1 9 2 15 15 13 7 13 2
8 16 0 13 9 13 10 15 2
24 7 16 13 13 7 13 1 9 1 0 2 3 13 15 0 13 2 7 10 13 3 0 13 2
6 3 15 15 13 13 2
7 7 3 15 13 1 9 2
17 0 9 1 15 13 2 16 16 13 9 13 2 13 3 1 0 2
4 7 13 15 2
15 15 15 13 0 2 3 13 13 16 13 15 15 0 13 2
29 7 16 1 0 13 1 13 7 13 2 10 13 3 0 13 2 16 13 16 13 13 2 15 7 13 16 0 13 2
4 3 15 13 2
21 7 3 13 9 15 9 15 13 1 0 9 9 2 15 13 9 13 0 9 0 2
5 0 9 15 13 2
17 16 10 13 13 2 7 15 9 13 0 1 15 2 7 1 9 2
9 16 1 9 2 3 3 13 0 2
11 15 3 13 1 9 0 2 3 13 0 2
7 13 13 3 15 13 13 2
9 7 16 13 3 13 2 3 13 2
4 16 9 13 2
6 3 13 13 15 13 2
9 3 2 16 15 13 2 15 13 2
14 15 7 13 9 1 0 2 16 3 3 15 9 13 2
6 3 0 3 13 13 2
9 16 1 0 13 3 13 0 0 2
17 7 3 15 9 2 10 13 1 15 13 2 3 13 1 9 0 2
12 3 2 16 15 12 13 13 1 9 1 15 2
16 7 12 15 13 1 15 2 0 13 16 15 1 15 13 13 2
30 16 2 16 0 7 0 13 1 9 2 7 1 9 13 0 1 0 2 0 13 16 1 15 15 13 13 0 1 0 2
31 16 3 13 7 13 13 1 15 1 9 2 13 7 13 1 15 1 15 15 13 2 0 13 16 13 13 1 15 15 13 2
14 7 1 15 13 13 9 1 12 15 12 1 15 13 2
11 16 15 3 13 1 15 2 7 1 9 2
15 16 7 13 9 13 0 1 15 2 0 13 0 7 9 2
15 16 7 13 16 13 13 15 9 9 15 13 2 7 15 2
25 16 15 2 3 13 16 13 13 2 7 0 16 13 13 2 7 16 13 13 2 7 1 15 9 2
5 15 7 13 0 2
14 3 13 0 13 13 9 2 13 0 0 13 3 13 2
14 7 3 15 13 1 15 7 3 13 2 15 13 0 2
27 16 7 1 15 9 9 13 2 3 3 16 13 13 1 9 2 7 13 1 9 13 2 7 3 1 15 2
16 1 13 13 9 7 9 9 2 13 16 3 13 13 1 0 2
12 7 3 13 15 0 13 15 3 13 1 15 2
24 16 9 15 13 16 13 9 15 9 16 2 13 10 9 7 9 9 2 3 13 13 1 0 2
17 16 2 16 13 1 9 13 7 13 13 2 3 13 13 1 9 2
8 7 1 15 13 15 15 0 2
20 3 16 15 15 13 1 15 9 9 2 1 15 13 2 16 3 0 7 13 2
14 3 13 16 13 13 15 0 15 3 13 1 15 0 2
35 16 0 2 15 13 16 13 0 13 15 3 13 1 15 0 2 3 13 16 13 3 0 2 3 0 13 9 2 13 16 15 13 13 0 2
11 12 9 2 3 16 15 0 13 3 0 2
6 15 13 2 13 13 2
9 3 2 16 13 15 0 13 0 2
10 15 9 2 16 15 0 13 1 15 2
5 7 15 13 0 2
15 16 15 13 1 15 2 3 13 0 15 15 13 1 15 2
16 3 7 1 13 0 9 0 13 1 15 13 2 3 1 15 2
9 7 2 15 13 2 3 15 13 2
12 3 3 13 13 16 13 15 15 13 1 15 2
20 16 3 13 13 9 2 3 16 15 3 13 7 13 2 7 0 1 15 9 2
25 7 3 16 15 3 13 1 9 7 9 2 3 13 2 16 3 2 13 9 2 13 0 1 9 2
13 13 3 16 12 9 15 13 13 3 7 15 13 2
7 7 3 13 15 15 0 2
7 3 16 15 13 13 0 2
15 3 7 13 13 16 15 9 13 2 3 16 12 1 15 2
10 7 16 12 9 13 15 7 13 15 2
6 7 16 15 13 9 2
6 7 16 9 13 15 2
17 16 13 13 9 2 3 16 15 3 13 7 13 1 15 9 9 2
9 7 16 3 13 1 9 7 9 2
14 7 0 16 15 3 13 0 13 15 2 7 9 9 2
15 13 3 16 13 15 13 12 9 13 0 7 13 15 9 2
31 7 16 1 13 15 15 13 1 15 2 3 1 9 2 9 13 2 3 9 2 16 13 0 1 15 2 13 3 1 9 2
17 0 13 16 0 13 15 9 13 3 13 7 1 15 7 1 9 2
23 13 3 15 15 13 1 15 2 3 9 2 1 13 0 2 9 13 1 15 13 1 9 2
16 0 13 7 13 15 0 13 1 15 0 13 15 15 13 0 2
18 3 0 13 15 9 13 15 13 15 15 7 1 15 7 1 9 13 2
17 16 7 0 13 2 1 10 9 2 15 13 15 13 0 2 13 2
24 16 3 9 13 0 2 16 15 13 2 13 16 9 13 15 15 13 0 7 0 2 13 0 2
12 7 15 9 3 13 13 9 15 15 13 15 2
5 16 3 3 13 2
4 7 3 10 2
5 7 16 0 13 2
6 7 16 3 3 13 2
20 13 3 16 13 13 15 13 15 0 2 15 13 9 9 1 15 9 13 15 2
13 7 3 9 15 3 13 7 1 15 7 1 9 2
29 3 2 1 13 15 13 16 15 13 1 0 13 1 15 9 15 3 13 1 15 9 2 16 9 13 7 9 13 2
11 15 3 9 15 9 13 15 13 1 9 2
19 1 15 13 13 16 15 13 15 13 3 15 9 13 1 15 7 1 9 2
7 7 0 13 15 13 3 2
18 15 3 13 9 13 0 2 1 10 15 9 1 9 0 13 15 13 2
19 13 3 16 0 13 15 13 1 9 15 3 13 7 1 15 7 1 9 2
20 7 13 1 15 9 16 9 9 9 13 9 0 2 7 3 13 13 1 9 2
21 16 13 13 1 9 3 9 15 15 2 7 9 10 0 2 15 13 9 0 9 2
36 7 16 9 3 13 9 15 13 15 2 0 9 2 1 10 0 2 13 1 15 9 15 13 9 13 15 2 15 9 13 3 2 15 13 9 2
24 1 3 10 13 15 13 1 9 2 13 16 9 15 13 9 13 15 2 13 1 9 15 0 2
7 15 13 15 0 1 13 2
7 3 13 13 3 13 13 2
8 0 7 13 13 3 3 13 2
13 13 3 13 0 9 13 3 0 2 15 9 13 2
7 13 7 9 12 13 13 2
11 15 0 13 2 16 13 1 9 9 9 2
7 15 1 0 13 13 0 2
28 7 1 15 13 16 9 0 1 13 9 13 13 1 9 9 9 2 15 13 2 0 13 13 0 16 9 13 2
24 3 16 9 7 9 1 0 13 2 0 13 16 13 13 15 9 15 1 0 13 9 7 9 2
14 16 10 15 1 0 13 2 1 15 9 13 13 9 2
15 1 15 13 15 1 9 1 9 7 1 3 13 1 13 2
20 0 13 2 16 13 1 13 9 0 13 2 3 9 0 2 4 13 1 15 2
7 1 15 13 15 13 13 2
6 15 1 0 3 13 2
24 7 1 15 13 13 16 2 16 0 13 3 13 13 1 15 2 13 16 13 0 1 3 0 2
9 3 3 9 1 9 15 9 13 2
27 16 3 13 7 3 13 1 0 13 0 13 2 7 1 13 15 2 1 15 3 13 1 13 0 0 13 2
28 13 7 9 15 9 1 12 8 2 1 13 3 13 13 1 0 1 9 0 2 7 13 13 1 12 9 0 2
5 7 15 13 9 2
6 7 15 9 15 13 2
16 1 10 9 0 13 0 13 9 0 2 7 0 13 9 0 2
8 7 13 12 2 7 0 0 2
10 13 7 9 2 13 15 15 13 9 2
11 3 2 13 0 2 0 9 13 3 13 2
14 7 16 13 1 9 0 1 0 2 15 9 13 0 2
9 3 10 15 13 2 15 13 0 2
6 15 7 13 0 0 2
8 3 13 13 0 9 0 13 2
4 15 9 13 2
9 13 3 15 9 13 1 9 9 2
17 1 12 3 8 13 16 15 15 13 0 0 2 13 7 0 9 2
31 1 12 7 8 13 13 15 0 0 2 1 15 16 13 12 0 12 15 13 3 0 2 3 13 16 15 13 3 15 0 2
14 15 7 13 1 9 1 15 15 13 0 7 0 0 2
12 1 15 13 13 0 13 15 15 13 0 9 2
5 7 15 13 9 2
13 1 15 3 13 1 9 15 9 13 1 9 9 2
8 15 3 13 9 1 12 9 2
4 7 13 15 2
29 0 13 15 0 7 13 1 12 9 13 3 7 0 16 15 9 2 1 15 10 7 0 13 16 1 0 9 13 2
27 7 1 9 13 9 0 9 1 12 9 13 2 3 16 0 7 1 9 2 7 16 3 7 1 0 9 2
9 13 3 13 15 15 9 9 13 2
5 7 15 13 9 2
9 16 1 9 9 13 13 9 9 2
17 13 3 16 13 15 0 9 2 15 9 13 2 13 15 9 13 2
11 13 7 9 9 13 0 1 9 0 9 2
14 3 0 9 10 9 15 9 10 13 2 10 9 13 2
10 7 3 15 13 3 13 13 15 13 2
10 7 0 15 13 9 13 15 3 13 2
17 3 7 15 9 3 13 2 3 0 1 9 10 1 15 13 13 2
14 3 3 15 9 13 2 3 9 15 1 15 0 13 2
14 13 3 9 15 1 15 9 0 1 10 15 9 13 2
22 3 7 1 9 15 9 13 2 0 15 1 9 13 2 1 15 13 1 0 15 13 2
11 7 3 9 13 2 15 1 9 15 13 2
8 7 3 13 9 9 0 9 2
33 7 16 1 9 9 0 3 13 13 15 2 3 9 2 7 9 15 1 15 9 1 0 9 13 13 2 13 15 13 1 9 0 2
37 16 7 1 0 9 12 15 13 2 7 3 1 0 9 9 13 1 16 1 0 13 13 2 3 12 9 0 1 15 13 2 15 1 0 13 13 2
16 16 2 16 13 9 3 13 9 2 1 15 1 10 9 13 2
15 3 16 13 15 3 13 9 2 13 15 3 1 15 9 2
17 7 3 1 9 1 10 15 15 13 1 15 2 1 9 3 13 2
15 7 3 1 9 15 13 0 9 1 13 16 1 10 13 2
13 3 3 13 9 2 16 3 13 15 1 15 13 2
27 1 13 3 1 9 9 1 9 9 2 13 9 15 15 1 0 3 0 13 2 3 16 9 13 3 0 2
7 15 3 9 0 9 13 2
5 13 3 8 12 2
7 15 9 2 7 3 13 2
3 8 12 2
6 1 15 3 13 9 2
4 7 8 12 2
9 3 13 9 3 9 2 16 13 2
5 16 9 13 0 2
9 1 15 7 13 0 9 13 0 2
15 3 10 15 13 13 7 13 2 1 9 7 9 15 13 2
8 13 7 4 9 13 3 0 2
9 13 3 0 2 13 9 7 9 2
2 3 2
20 15 0 9 13 15 13 2 15 16 9 13 9 9 2 16 13 1 12 9 2
12 9 7 13 3 1 9 2 16 3 13 4 2
5 9 3 3 13 2
10 3 1 15 3 13 0 7 0 13 2
33 3 3 13 9 1 3 9 2 7 3 9 1 9 13 13 2 7 15 9 1 9 15 13 13 2 16 15 1 9 13 3 13 2
13 13 3 13 9 7 9 2 15 9 10 3 13 2
6 1 15 9 9 13 2
2 3 2
18 16 3 3 13 7 3 13 2 1 15 13 4 1 3 13 1 13 2
4 3 1 15 2
9 16 15 3 13 3 13 15 13 2
10 16 7 1 15 2 15 13 0 15 2
8 13 7 4 9 13 0 9 2
5 3 3 13 13 2
15 3 7 13 13 2 16 15 3 13 2 13 9 3 13 2
4 13 3 0 2
2 0 2
17 13 1 9 15 15 13 0 13 7 3 13 2 3 0 7 0 2
10 10 7 15 13 0 13 2 9 13 2
31 16 2 1 1 15 0 15 13 1 12 2 3 13 7 3 13 2 13 2 16 15 13 13 2 16 15 13 1 15 9 2
17 7 1 9 3 13 13 1 0 2 16 1 13 4 1 9 9 2
8 3 13 13 15 15 13 13 2
19 10 7 0 7 13 9 10 9 3 2 7 3 2 7 13 1 15 0 2
15 3 13 7 13 1 0 1 0 15 13 9 10 9 3 2
13 3 13 13 15 0 0 2 15 13 1 15 0 2
14 7 15 9 13 2 1 13 9 0 2 16 13 4 2
13 13 3 9 0 2 1 10 0 1 15 13 0 2
9 13 3 9 1 9 9 9 9 2
8 1 15 3 13 9 9 13 2
7 0 7 9 13 9 13 2
4 13 3 0 2
14 13 7 9 9 7 9 2 3 13 9 1 9 9 2
13 3 2 16 9 13 2 13 16 1 15 13 13 2
8 15 16 13 2 15 13 13 2
15 7 3 7 1 0 13 2 7 13 1 15 15 3 13 2
8 15 7 9 0 9 9 13 2
3 3 9 2
9 15 7 2 9 2 1 0 13 2
3 7 15 2
12 15 7 15 15 13 2 7 9 10 3 13 2
8 16 1 9 3 13 9 0 2
14 16 7 9 0 13 2 0 13 15 3 13 1 9 2
28 10 3 15 1 15 9 13 9 2 1 15 15 13 1 9 13 3 13 2 16 15 13 13 2 13 3 13 2
13 9 7 1 15 3 13 3 13 2 1 13 0 2
9 1 9 3 3 13 9 1 13 2
2 3 2
26 16 15 15 3 13 1 9 3 9 2 0 13 9 1 9 16 1 9 2 3 0 9 13 0 9 2
21 16 9 3 13 15 1 9 2 7 13 16 13 1 9 1 15 15 13 1 9 2
14 10 3 15 13 15 9 1 9 2 13 15 0 15 2
15 9 7 13 0 9 7 0 9 2 16 1 1 13 13 2
9 3 3 13 1 15 15 9 13 2
2 3 2
14 15 15 13 1 15 0 13 2 15 9 13 0 13 2
12 16 15 13 1 15 0 13 2 3 13 9 2
15 10 7 15 13 0 13 2 13 9 2 16 1 13 4 2
8 9 7 13 1 15 0 13 2
7 15 3 9 13 0 13 2
8 15 3 9 1 10 9 13 2
2 3 2
7 15 13 1 16 13 9 2
16 15 3 3 13 15 9 2 3 15 15 13 2 7 15 15 2
12 15 7 3 15 15 13 2 3 13 0 9 2
10 13 3 15 9 2 3 1 9 10 2
18 0 3 9 2 15 9 13 2 15 13 9 13 2 7 13 9 0 2
2 3 2
18 15 2 16 13 4 13 16 13 9 2 3 13 4 13 16 13 9 2
7 3 9 13 9 9 13 2
13 7 9 13 3 0 7 0 2 16 13 1 13 2
9 15 3 13 1 9 2 3 0 2
2 3 2
12 13 15 13 1 9 15 13 1 9 1 9 2
17 3 7 13 15 1 9 1 9 2 16 15 13 9 2 3 13 2
5 3 7 13 13 2
14 3 13 13 15 15 0 2 15 13 1 9 1 9 2
24 7 3 2 16 15 13 13 1 9 1 9 2 13 1 15 15 15 13 2 15 13 1 9 2
8 15 7 1 0 13 3 13 2
15 3 13 13 1 15 15 13 3 9 7 15 9 1 9 2
5 7 15 13 9 2
7 16 1 9 3 13 9 2
9 13 3 1 15 9 3 13 9 2
10 16 9 15 15 13 2 1 9 13 2
2 3 2
6 9 3 13 13 9 2
12 3 13 7 9 1 15 3 13 2 1 9 2
14 9 7 13 13 0 9 0 9 2 16 1 13 4 2
6 15 3 9 3 13 2
2 0 2
16 13 9 0 9 13 15 15 10 1 9 13 16 1 9 0 2
7 1 15 13 1 12 9 2
20 16 3 9 2 15 13 0 9 2 13 9 0 9 2 13 10 1 9 13 2
2 3 2
14 9 3 13 9 15 1 9 16 1 16 13 7 13 2
20 16 3 9 13 0 2 16 13 4 2 15 9 13 13 9 9 1 9 9 2
21 15 7 9 9 0 13 2 15 9 3 1 10 9 2 7 1 15 13 10 13 2
41 1 15 7 9 9 1 9 13 2 15 13 4 13 9 13 15 16 0 9 2 1 15 16 2 16 3 13 15 2 13 13 15 15 9 2 7 3 3 13 0 2
15 3 1 15 15 1 9 1 15 13 2 15 9 9 13 2
14 15 7 13 1 9 15 13 15 1 9 7 9 13 2
20 13 3 2 16 1 12 8 13 2 13 1 15 2 3 10 13 15 13 13 2
13 0 7 15 0 13 2 1 15 16 3 13 15 2
11 9 3 1 15 13 13 15 1 15 13 2
10 13 3 15 1 15 13 1 16 13 2
13 16 12 9 13 1 9 2 3 13 16 9 13 2
19 1 15 7 15 1 15 13 2 3 13 13 15 13 2 7 15 0 13 2
9 3 3 7 13 9 1 3 13 2
9 3 3 13 9 3 9 10 9 2
13 7 3 3 13 13 15 13 2 15 3 0 13 2
23 3 3 9 7 9 0 13 2 15 12 13 9 0 2 15 9 0 2 1 15 9 13 2
7 16 1 9 15 13 9 2
12 1 13 7 13 13 16 1 9 15 13 9 2
10 3 1 10 9 13 13 9 7 9 2
17 3 3 0 13 0 12 13 16 15 13 3 9 2 7 15 9 2
19 15 3 9 13 2 3 13 16 3 13 7 13 2 15 3 13 12 0 2
12 1 15 3 15 9 13 13 16 9 9 13 2
11 13 3 13 1 9 16 13 1 9 0 2
7 1 9 7 15 13 9 2
8 3 13 3 1 15 15 9 2
2 3 2
7 10 9 0 13 10 13 2
13 0 3 9 2 15 9 13 2 1 15 13 13 2
2 3 2
21 10 9 13 9 0 2 3 13 1 9 9 2 16 1 15 13 15 15 9 13 2
12 15 7 13 0 2 13 1 9 1 3 13 2
11 15 9 3 13 2 1 13 1 15 13 2
8 3 13 3 1 15 15 9 2
2 0 2
6 10 9 13 15 13 2
9 16 3 9 13 2 1 0 13 2
17 15 7 1 15 13 0 2 1 12 3 13 16 1 15 13 13 2
9 16 3 13 13 9 2 13 13 2
14 3 3 15 15 13 13 2 16 15 13 9 15 15 2
9 13 3 0 15 2 15 13 0 2
7 13 7 13 9 0 13 2
6 3 9 13 9 0 2
12 7 3 3 13 9 0 2 15 1 13 4 2
2 3 2
23 1 15 9 3 15 13 0 3 0 2 16 1 9 0 9 2 15 3 13 15 0 9 2
15 15 3 13 1 9 9 10 9 2 13 13 1 9 9 2
18 15 7 15 13 1 9 9 10 9 2 13 9 2 1 13 0 9 2
6 9 3 13 0 9 2
7 15 3 9 15 13 13 2
2 3 2
29 1 10 9 9 3 13 15 7 15 9 2 7 15 2 2 7 13 9 1 15 9 15 13 0 15 7 9 15 2
7 3 9 13 0 9 15 2
31 16 9 9 3 13 9 2 9 3 9 0 3 13 9 0 2 7 0 9 9 3 13 1 9 9 15 1 15 9 13 2
22 16 3 9 13 13 2 9 7 9 15 0 13 1 15 2 3 7 1 15 15 9 2
14 7 3 3 13 1 15 0 15 9 15 13 0 15 2
9 3 13 3 15 0 7 0 9 2
2 3 2
7 1 10 9 13 13 9 2
7 1 10 7 9 13 9 2
15 3 13 15 15 13 1 10 2 3 9 2 10 9 13 2
10 16 1 9 15 13 0 7 1 9 2
16 1 15 7 9 13 16 1 9 15 13 13 0 7 1 9 2
17 10 3 15 1 15 15 0 7 1 9 13 2 15 15 13 13 2
14 3 15 13 1 9 9 3 13 13 0 7 1 9 2
9 15 7 0 13 1 15 15 13 2
6 1 15 3 9 13 2
20 1 3 9 13 0 2 16 13 4 2 15 1 15 13 13 0 7 1 9 2
2 0 2
7 9 9 13 9 1 15 2
20 1 9 7 3 13 9 1 15 2 7 13 1 15 0 2 7 9 9 15 2
7 3 15 1 15 13 13 2
2 3 2
17 3 13 15 0 2 3 13 13 15 1 15 15 9 1 15 13 2
9 3 0 13 15 15 13 1 9 2
26 7 1 9 3 13 0 13 15 1 15 15 1 15 15 13 2 1 1 15 13 13 2 16 13 4 2
9 3 13 3 1 15 13 15 0 2
2 3 2
15 10 1 15 13 15 0 7 0 2 13 4 1 15 13 2
12 3 0 13 15 9 13 1 15 13 9 13 2
10 9 7 13 3 0 2 16 13 4 2
11 3 3 13 1 15 13 15 0 7 0 2
6 16 9 3 13 9 2
10 1 13 3 13 16 9 3 13 9 2
14 10 3 9 2 1 13 0 2 13 13 7 9 13 2
10 9 7 3 13 13 2 16 13 4 2
5 3 9 3 13 2
2 3 2
8 10 15 13 15 9 1 9 2
8 3 0 13 9 0 1 0 2
7 9 7 1 0 13 0 2
6 10 7 9 13 15 2
7 3 10 9 13 1 9 2
15 9 7 3 13 1 9 2 7 9 0 2 16 13 4 2
6 3 9 3 13 9 2
2 3 2
12 16 9 13 9 2 13 16 13 15 9 0 2
19 3 9 0 3 13 1 15 13 2 16 9 13 2 15 16 9 9 13 2
14 3 7 13 9 0 2 1 13 0 2 16 13 4 2
7 10 7 9 0 0 13 2
6 9 3 3 13 9 2
2 0 2
5 10 9 13 13 2
15 15 3 1 9 0 8 1 13 13 1 12 9 7 9 2
10 15 7 9 13 9 7 9 13 13 2
16 16 3 9 13 9 2 9 7 9 10 15 0 9 13 13 2
9 7 3 9 3 13 0 9 10 2
4 15 13 9 2
5 3 13 3 9 2
2 3 2
7 9 0 0 13 16 0 2
9 13 7 15 13 9 1 9 9 2
4 3 7 9 2
12 7 1 9 9 13 9 9 2 16 7 9 2
12 3 1 10 0 13 15 0 1 9 9 13 2
9 10 7 9 1 9 13 13 0 2
9 3 1 10 9 13 15 13 0 2
13 16 3 9 13 9 2 3 13 0 7 0 9 2
2 3 2
9 15 9 3 13 9 13 13 0 2
18 15 7 9 13 10 9 13 0 2 1 1 15 13 1 15 9 9 2
11 15 3 15 15 13 0 2 9 3 13 2
5 15 7 13 9 2
5 3 3 13 9 2
2 3 2
15 13 9 9 1 15 13 13 1 9 9 2 1 15 9 2
23 1 10 9 0 13 16 0 13 3 13 7 1 15 7 1 9 2 16 1 1 13 13 2
8 9 7 9 13 0 9 0 2
13 3 0 9 15 3 13 7 1 15 7 1 9 2
17 15 7 9 13 0 16 13 2 15 16 13 13 7 13 13 3 2
16 7 3 9 13 13 13 2 1 15 16 13 3 1 9 13 2
22 15 3 9 1 9 13 16 1 9 13 2 16 2 13 9 2 13 1 9 9 9 2
12 3 0 9 9 3 13 9 7 9 1 9 2
17 15 7 1 15 0 13 9 9 16 1 0 13 0 2 13 9 2
6 9 3 3 13 9 2
2 3 2
8 15 9 0 13 9 1 9 2
7 9 0 9 13 9 0 2
7 3 3 13 1 15 9 2
18 7 3 9 2 15 13 0 9 2 7 13 9 7 13 9 1 9 2
4 0 3 13 2
16 16 9 9 15 13 0 2 7 3 13 9 13 2 7 0 2
17 9 0 15 13 2 16 13 1 12 8 7 1 12 9 7 9 2
10 9 7 13 3 13 0 13 9 0 2
10 7 3 1 15 9 13 13 9 0 2
14 16 7 1 9 13 3 13 13 9 0 2 3 13 2
17 0 9 15 13 9 0 1 9 0 2 13 9 0 1 9 0 2
21 15 13 15 9 2 7 13 1 9 2 7 1 9 0 2 7 1 15 15 9 2
9 7 9 0 13 0 10 9 13 2
16 3 13 16 1 0 13 9 2 0 13 2 16 9 15 13 2
10 7 13 13 16 1 0 16 13 9 2
9 13 3 16 15 13 1 0 9 2
11 7 3 13 7 13 7 9 13 1 9 2
8 15 0 13 4 1 12 9 2
16 16 7 3 13 9 0 9 13 13 1 9 2 3 3 13 2
7 13 9 0 15 13 8 2
7 13 9 15 15 13 8 2
8 9 3 15 13 1 9 0 2
21 13 3 13 15 9 15 9 1 9 1 15 13 15 9 2 1 15 9 13 13 2
13 13 3 15 12 9 1 8 9 15 1 3 13 2
13 3 3 3 1 15 9 13 15 7 15 9 13 2
26 16 7 13 1 9 13 13 2 13 13 1 9 1 9 9 1 9 2 1 0 9 1 0 9 13 2
27 16 3 13 8 2 15 9 13 1 9 15 13 0 9 9 1 15 13 0 9 13 0 9 2 3 8 2
21 7 3 15 9 15 13 8 15 2 13 9 13 2 1 13 9 13 1 9 13 2
12 13 3 16 1 0 9 13 9 13 7 0 2
4 15 13 0 2
12 3 3 9 0 9 13 13 13 1 9 15 2
11 16 7 9 0 9 13 0 2 3 13 2
8 15 9 13 13 13 9 0 2
15 7 9 0 9 13 1 9 0 2 16 9 0 13 0 2
7 3 9 0 9 13 0 2
4 0 3 13 2
38 16 15 9 13 15 9 13 9 0 2 9 15 9 2 13 9 9 2 13 1 9 0 2 16 3 15 13 0 9 2 3 1 0 9 9 13 13 2
17 7 3 9 13 13 9 13 2 0 7 9 1 0 9 13 13 2
18 7 3 3 2 1 16 13 1 9 9 2 13 1 9 1 15 9 2
13 7 9 3 13 13 1 9 15 2 7 3 13 2
15 3 7 9 1 9 9 13 1 9 9 1 15 13 15 2
11 9 7 1 15 15 13 2 13 13 0 2
7 3 9 13 13 9 0 2
4 15 13 0 2
8 7 1 15 9 0 13 9 2
25 15 12 13 2 16 13 13 16 15 9 15 13 0 9 2 3 13 0 2 16 13 1 9 0 2
8 13 7 9 13 1 9 15 2
14 7 1 15 13 16 0 13 13 0 15 13 13 0 2
13 7 16 15 13 15 13 9 15 0 2 13 0 2
19 16 2 16 15 13 9 15 0 2 16 9 13 2 13 9 2 13 0 2
10 7 1 9 15 13 13 9 9 13 2
19 16 15 0 13 0 2 16 9 0 13 2 9 15 13 0 9 16 15 2
17 15 7 0 9 13 16 13 0 13 13 9 2 1 0 15 13 2
6 3 13 15 13 0 2
12 7 0 13 13 16 13 9 1 9 9 13 2
18 16 3 13 13 1 9 9 9 1 10 9 15 13 9 1 9 15 2
11 13 3 0 0 2 15 1 13 9 13 2
29 0 9 13 16 2 16 9 13 2 15 9 13 13 15 9 15 3 13 13 9 2 16 9 0 3 13 13 9 2
40 7 1 15 13 13 16 1 9 13 3 13 16 3 13 9 13 9 16 9 0 9 0 2 7 16 3 13 9 1 9 16 9 0 2 15 13 1 9 9 2
15 3 3 13 1 9 0 16 3 13 9 7 9 1 9 2
15 16 7 9 2 3 13 13 9 16 9 2 15 9 13 2
38 0 9 13 16 2 16 15 9 13 9 13 2 16 1 13 9 13 2 1 9 7 13 3 13 15 13 9 0 2 13 16 15 9 13 13 9 0 2
8 7 3 9 0 1 9 13 2
26 1 15 7 1 15 13 16 9 0 1 9 10 13 13 2 7 9 9 13 1 15 15 13 9 0 2
18 7 15 9 13 13 9 2 15 1 9 0 9 13 13 1 15 9 2
18 9 10 13 0 2 9 7 10 0 2 16 9 10 0 13 9 10 2
10 15 7 9 13 9 2 1 12 8 2
23 3 0 13 2 1 15 2 16 15 15 13 1 15 0 3 13 2 13 9 13 1 15 2
8 13 3 16 0 13 1 9 2
6 15 13 0 1 15 2
8 7 3 15 1 15 9 13 2
12 16 1 9 0 10 9 15 13 2 13 13 2
8 3 3 13 16 13 10 9 2
22 13 3 1 9 0 2 1 9 2 1 12 8 2 9 1 3 2 7 3 1 13 2
12 7 3 3 13 16 13 15 9 1 3 13 2
10 13 3 16 15 9 9 3 13 0 2
53 16 2 16 13 16 1 9 0 3 13 9 3 0 1 13 2 15 13 9 9 2 13 3 1 15 9 3 0 2 15 13 9 13 2 1 13 9 13 2 1 12 9 7 9 2 16 9 13 9 16 13 3 2
21 7 3 0 13 13 16 2 1 9 13 1 9 2 13 13 1 9 1 9 9 2
10 9 7 1 15 9 9 13 7 9 2
11 3 9 15 0 13 16 9 13 13 0 2
8 9 7 3 13 15 9 9 2
11 0 1 9 15 9 13 0 2 16 9 2
46 7 3 3 13 16 9 13 13 0 1 9 13 2 16 1 0 13 2 16 3 13 16 1 15 9 15 13 1 12 9 7 9 0 2 1 9 15 0 3 13 1 9 16 1 9 2
29 0 9 13 1 15 16 3 13 13 0 16 15 15 13 9 0 2 13 9 0 2 1 15 13 15 13 3 13 2
22 16 15 9 15 13 1 9 15 2 3 3 0 9 13 13 16 15 9 13 16 1 2
28 16 9 9 13 13 2 7 2 16 1 13 15 9 0 3 13 2 0 9 13 13 1 15 9 2 1 9 2
16 7 1 15 13 13 16 9 3 13 16 13 2 16 13 4 2
15 7 3 2 16 13 9 15 3 13 2 13 15 3 13 2
16 1 10 7 15 13 13 9 1 13 2 16 9 9 13 13 2
17 7 3 2 3 13 1 15 2 10 9 15 13 0 13 3 13 2
16 7 15 0 13 3 13 2 3 13 1 15 16 0 9 13 2
9 7 3 3 16 1 0 9 13 2
19 13 3 13 9 1 9 13 9 13 2 15 3 13 1 15 13 9 0 2
24 7 9 15 1 15 0 13 13 7 3 13 2 13 7 3 13 2 13 13 9 9 1 15 2
5 15 13 13 0 2
8 7 3 13 0 13 13 0 2
23 7 3 15 13 1 9 9 13 2 15 13 1 15 9 1 13 2 13 3 9 1 13 2
24 3 7 15 0 9 0 2 1 9 2 13 0 9 9 9 0 13 2 1 16 9 13 9 2
32 7 13 9 1 9 16 15 15 1 15 13 1 9 13 7 3 13 2 13 1 15 9 9 2 16 13 13 0 1 9 13 2
10 3 9 13 15 9 1 13 1 0 2
17 7 3 13 15 0 13 1 15 9 9 2 15 3 13 1 15 2
10 9 7 13 15 13 7 13 1 9 2
28 7 3 15 1 15 13 1 9 1 3 13 2 3 13 2 16 15 13 2 1 9 9 13 1 15 9 13 2
22 0 9 13 16 1 13 9 3 13 0 9 3 3 13 9 0 1 9 16 1 9 2
9 3 3 13 16 13 3 1 9 2
28 7 1 15 13 16 13 7 0 1 9 7 9 7 9 13 1 12 9 2 16 13 1 12 7 1 12 8 2
12 7 3 0 1 12 15 13 9 13 1 15 2
15 1 15 7 15 13 9 2 3 13 13 7 0 16 0 2
11 3 13 9 13 1 15 9 9 3 13 2
51 15 7 13 7 0 2 16 9 13 12 9 2 12 0 2 15 13 13 9 2 7 1 15 13 16 9 15 13 13 9 2 7 15 13 2 15 13 0 9 2 1 15 13 16 9 15 13 13 0 9 2
20 7 3 13 16 9 0 15 3 13 1 9 2 13 13 9 3 0 1 9 2
18 7 9 15 13 1 9 13 16 13 0 2 1 15 9 13 16 13 2
12 3 2 16 13 2 13 16 13 1 3 9 2
19 13 3 0 13 16 9 15 3 13 1 9 13 9 2 7 13 1 9 2
13 3 13 1 9 0 2 7 3 1 9 10 9 2
24 9 7 15 13 1 9 3 13 13 16 1 9 9 2 16 13 4 16 9 3 13 9 0 2
10 7 3 13 1 9 1 9 10 9 2
11 3 13 2 16 13 2 16 13 1 9 2
12 1 15 3 2 13 13 9 2 13 9 9 2
2 0 2
25 15 9 15 13 1 13 0 13 13 0 7 0 2 15 16 13 0 1 9 0 13 13 7 13 2
29 15 7 15 13 7 13 3 1 15 9 15 13 1 13 1 9 9 1 1 9 2 1 3 13 0 2 3 13 2
11 7 3 15 9 13 13 9 0 7 0 2
14 9 7 0 13 0 7 0 2 16 13 1 12 8 2
8 3 13 0 9 3 13 9 2
2 3 2
28 15 9 15 13 1 9 15 13 1 9 1 9 2 13 13 0 2 16 2 1 13 4 1 9 2 9 13 2
21 16 3 9 0 13 0 2 13 16 13 1 9 15 13 3 7 10 9 1 9 2
23 15 7 3 13 15 9 7 15 9 1 9 2 1 10 3 13 0 1 15 7 1 9 2
12 3 9 0 9 3 13 9 7 9 1 9 2
13 9 7 0 9 13 0 13 2 15 13 16 13 2
5 15 7 13 9 2
10 9 3 7 13 9 7 9 1 9 2
48 16 7 0 13 2 1 9 10 2 16 9 9 13 0 2 16 1 13 2 3 0 13 16 9 15 3 13 7 1 9 9 2 7 1 9 9 0 2 1 3 13 9 9 1 9 9 13 2
8 3 9 13 10 9 3 13 2
8 15 7 9 13 13 0 9 2
5 13 3 8 12 2
17 9 13 9 2 7 15 15 15 13 2 1 9 7 9 13 13 2
6 13 3 12 8 12 2
9 9 9 0 2 0 2 0 9 2
4 7 8 12 2
10 0 9 1 15 15 13 4 13 13 2
11 15 3 3 9 7 9 13 2 0 13 2
24 1 15 7 13 9 0 9 0 2 15 3 13 16 9 0 2 16 9 7 9 7 15 3 2
13 7 3 0 9 9 9 13 2 7 15 13 9 2
12 1 15 3 15 13 13 9 13 9 7 9 2
7 15 3 1 13 9 13 2
21 3 2 1 9 7 9 13 1 9 1 15 2 13 0 9 13 13 9 1 9 2
12 15 3 13 9 13 13 1 12 9 7 9 2
11 1 15 13 13 16 13 9 13 9 0 2
14 1 0 7 0 9 1 9 13 2 13 9 13 10 2
35 15 3 9 13 0 13 15 9 9 7 9 1 15 13 9 13 2 16 9 2 9 2 9 2 9 7 3 2 9 13 1 13 9 9 2
36 13 3 9 13 9 0 0 2 9 2 9 7 9 0 15 9 0 9 13 2 3 7 9 2 15 15 0 9 9 1 0 9 13 9 13 2
22 15 10 9 13 9 16 1 0 13 1 9 13 2 1 15 3 13 13 16 9 9 2
9 7 3 15 1 0 13 13 13 2
6 16 9 13 10 9 2
15 1 13 7 13 13 16 9 13 10 9 2 9 7 9 2
17 1 10 3 15 15 3 13 10 9 7 9 2 13 15 13 9 2
32 1 3 1 15 13 10 9 2 16 15 1 15 13 1 15 9 2 15 15 9 13 13 15 9 2 7 3 15 13 10 9 2
17 16 3 15 3 13 10 9 2 13 15 1 15 13 1 15 9 2
8 7 3 13 1 15 13 9 2
15 3 3 9 1 9 13 1 9 9 2 16 9 1 9 2
9 13 4 7 1 9 15 13 9 2
6 9 3 13 10 9 2
2 3 2
15 0 15 13 13 1 9 7 9 9 15 3 13 9 15 2
7 9 3 13 15 13 9 2
11 0 7 9 9 13 15 1 9 3 13 2
11 0 3 9 13 1 9 15 1 9 15 2
11 1 9 7 3 13 15 9 2 16 13 2
9 15 3 13 1 15 1 9 15 2
6 13 3 15 10 9 2
2 0 2
28 9 15 1 9 0 3 13 2 7 1 0 7 1 0 13 2 13 9 15 3 1 15 0 13 1 15 13 2
27 3 3 13 16 9 7 9 7 0 13 9 2 16 9 3 13 1 15 0 0 2 7 13 1 9 0 2
16 0 3 9 0 3 13 1 15 0 2 7 13 1 0 9 2
14 3 3 13 16 15 9 2 7 9 2 13 10 9 2
30 15 3 9 7 9 9 7 9 13 1 9 13 15 7 15 9 2 16 3 9 9 7 9 9 13 7 9 1 0 2
12 3 3 13 16 9 2 7 9 2 13 9 2
24 7 0 9 13 1 15 0 13 7 1 15 13 2 1 3 13 1 15 9 2 16 13 4 2
10 0 3 9 13 1 9 2 16 13 2
5 9 13 10 9 2
2 3 2
24 9 9 7 13 9 15 7 15 13 1 15 15 9 16 9 2 1 9 1 10 9 9 13 2
18 7 15 9 13 13 15 9 9 2 1 13 0 9 2 16 13 4 2
6 9 3 13 10 9 2
2 3 2
18 15 3 13 10 9 2 15 13 1 15 15 1 15 16 9 1 9 2
13 3 7 1 9 9 13 9 2 16 13 2 9 2
12 7 1 9 15 13 9 2 16 1 13 4 2
8 13 3 16 15 13 10 9 2
9 16 1 9 15 13 9 7 9 2
24 1 15 7 15 1 13 4 2 0 13 13 16 1 9 3 13 15 9 7 9 16 10 9 2
17 13 4 3 1 15 13 15 1 15 0 13 13 2 15 9 13 2
45 15 3 9 15 0 13 2 16 13 15 9 15 3 13 15 15 13 2 7 13 0 15 9 7 13 2 16 1 15 13 9 9 2 7 15 0 7 0 2 16 9 13 1 15 2
22 16 0 9 2 15 9 3 13 13 15 13 1 15 0 2 16 7 9 1 15 13 2
25 16 7 0 9 2 13 16 7 9 3 13 1 9 2 7 15 1 15 9 2 7 9 1 9 2
25 0 12 13 1 9 15 15 13 1 15 13 2 16 2 16 1 15 13 2 3 3 13 0 9 2
30 1 0 0 13 16 15 9 0 13 1 9 15 1 15 0 13 13 2 16 10 15 13 1 9 9 2 13 15 0 2
7 7 3 3 13 15 9 2
11 9 3 3 13 9 15 3 13 10 9 2
32 7 1 15 13 13 16 15 9 3 0 13 1 9 15 2 16 3 3 13 16 15 13 2 7 13 3 1 9 15 15 13 2
18 7 3 15 9 1 15 0 13 2 7 15 13 3 1 15 0 13 2
8 15 7 9 13 9 3 13 2
21 16 16 15 9 13 13 1 15 9 2 13 16 15 9 0 15 13 1 15 9 2
11 7 15 15 13 1 15 13 13 15 9 2
15 3 15 9 15 13 0 1 15 15 13 1 15 0 13 2
6 3 3 13 9 15 2
12 15 7 15 13 1 1 15 13 2 13 9 2
13 3 3 15 13 9 9 2 7 15 9 9 0 2
27 16 7 3 13 13 15 9 1 15 9 2 3 15 9 0 13 1 15 1 15 13 9 10 1 9 15 2
7 7 3 13 15 16 0 2
2 3 2
6 15 13 1 10 9 2
13 15 3 3 13 10 9 2 3 13 1 15 13 2
7 9 7 13 1 15 13 2
6 3 9 13 10 9 2
2 0 2
35 16 9 9 3 13 10 9 2 3 7 9 15 13 13 2 1 9 0 13 0 2 16 13 4 2 13 16 3 9 13 15 1 9 15 2
18 10 7 15 13 15 15 3 13 1 9 15 2 13 15 1 15 9 2
18 15 3 15 1 15 3 13 12 2 16 13 2 13 1 15 9 13 2
9 9 3 13 15 9 1 15 9 2
21 7 3 1 15 15 13 1 9 15 9 2 7 1 9 15 2 7 1 15 15 2
20 16 0 9 2 9 7 13 1 15 9 2 13 16 15 13 15 15 9 13 2
15 15 7 13 0 2 16 0 1 9 13 9 13 16 9 2
19 16 3 15 15 15 13 9 13 2 13 13 16 13 9 2 15 13 0 2
19 2 16 13 16 15 13 15 9 13 1 9 0 2 15 9 13 1 15 2
6 15 3 3 13 0 2
19 13 3 15 9 0 13 1 9 15 9 2 1 15 9 13 9 0 9 2
12 3 7 3 13 1 9 0 2 7 1 0 2
9 16 7 15 13 1 15 15 9 2
18 10 7 15 13 9 1 15 9 2 4 13 2 7 3 13 9 0 2
14 9 7 13 0 9 3 13 9 2 16 1 13 4 2
13 3 15 9 15 13 9 3 2 3 13 9 9 2
10 0 13 3 16 9 9 9 10 13 2
2 0 2
5 9 9 15 13 2
20 3 3 13 13 15 1 15 16 13 1 9 2 7 1 15 16 13 1 9 2
20 10 7 15 13 9 15 0 1 15 13 2 15 13 1 15 16 9 1 9 2
9 9 3 7 9 1 15 3 13 2
22 16 3 0 9 13 15 16 10 9 2 13 16 9 7 9 15 13 16 9 7 9 2
16 13 4 7 1 9 15 13 1 9 2 7 15 13 0 9 2
10 3 3 9 9 13 15 16 10 9 2
2 3 2
13 10 15 15 3 13 13 16 13 0 2 13 13 2
23 7 15 9 1 15 13 15 9 7 15 9 2 13 13 16 13 0 2 3 9 7 9 2
15 3 10 9 1 15 13 15 9 7 15 9 2 13 13 2
10 9 7 3 13 13 2 16 13 4 2
8 15 3 9 9 13 10 9 2
2 0 2
9 10 9 13 1 15 16 13 9 2
23 15 3 9 15 9 3 13 10 9 2 13 1 9 10 2 7 9 15 2 3 15 9 2
27 15 7 13 1 9 15 2 3 13 13 0 9 2 16 15 15 15 13 1 15 16 13 2 13 15 0 2
11 9 7 13 0 9 2 15 15 13 0 2
7 9 3 9 13 10 9 2
20 15 7 0 9 9 1 9 4 13 2 15 1 13 1 9 2 8 12 13 2
11 16 13 1 15 9 9 2 15 9 15 2
4 15 13 15 2
3 9 13 2
5 15 13 15 13 2
5 3 13 9 9 2
15 15 13 13 15 1 15 2 13 10 0 9 13 15 13 2
13 15 7 9 4 13 1 13 9 7 9 15 9 2
12 3 13 16 15 0 9 13 10 9 7 9 2
8 15 3 9 0 9 13 4 2
9 13 3 9 2 1 9 1 8 2
19 9 3 13 9 9 2 7 0 9 2 7 13 9 2 7 0 9 9 2
21 9 3 13 2 1 9 1 8 2 16 0 9 13 15 9 7 1 15 13 9 2
7 16 1 9 3 13 9 2
22 1 15 3 9 1 9 13 16 9 1 15 9 15 13 13 2 7 15 15 0 13 2
23 15 3 9 3 13 13 15 15 3 13 1 9 10 2 16 15 15 13 13 15 15 13 2
9 15 3 13 0 7 0 16 9 2
8 7 3 15 9 15 13 13 2
7 0 7 9 13 15 9 2
10 3 15 13 15 3 13 1 10 9 2
7 15 3 9 15 13 13 2
2 0 2
19 10 15 13 15 0 2 13 9 3 13 2 1 13 1 9 15 15 13 2
16 16 3 15 0 13 1 9 2 13 16 15 13 1 15 9 2
13 7 3 9 9 13 15 0 9 2 7 15 15 2
12 16 15 15 2 13 16 15 13 1 0 9 2
39 15 3 13 15 9 2 7 0 7 0 2 1 15 13 2 16 15 9 13 1 15 2 15 16 13 15 15 13 16 13 15 9 2 15 3 13 1 9 2
9 3 9 13 7 13 1 15 9 2
5 15 13 1 13 2
12 16 7 15 0 9 13 9 9 15 15 13 2
23 0 13 7 16 13 9 15 1 16 13 13 15 2 16 3 15 1 15 13 15 1 9 2
34 3 13 2 16 1 9 13 15 9 2 16 1 15 7 15 13 7 13 9 15 2 16 0 13 0 9 1 9 9 7 13 1 9 2
6 3 3 9 13 13 2
6 15 0 0 13 4 2
2 3 2
24 10 9 9 13 1 15 16 9 1 9 2 15 16 9 15 9 13 13 9 9 1 9 0 2
12 7 1 9 15 13 9 2 16 1 13 4 2
8 1 15 3 15 9 13 13 2
2 3 2
13 15 13 15 0 2 13 15 9 1 10 9 0 2
11 9 3 1 15 13 4 13 7 3 13 2
15 16 3 9 13 15 0 15 13 2 13 16 15 13 0 2
6 15 0 1 13 4 2
2 0 2
20 15 13 15 9 2 3 13 15 13 1 15 2 16 9 3 13 1 9 9 2
8 7 9 13 15 1 15 13 2
7 1 9 3 15 13 9 2
4 0 3 13 2
9 15 0 13 1 9 16 1 9 2
6 9 7 13 10 9 2
12 3 15 13 1 15 2 0 9 1 15 13 2
9 9 7 13 15 15 15 13 15 2
15 15 3 9 13 12 16 1 15 15 0 13 16 9 9 2
11 15 3 13 9 13 16 1 15 0 13 2
8 13 3 16 9 13 15 13 2
2 3 2
12 9 3 13 1 9 2 16 9 13 1 9 2
13 15 7 3 13 1 15 2 13 3 13 1 15 2
8 3 13 15 9 13 1 9 2
13 15 7 0 13 0 9 13 2 15 13 9 0 2
8 0 3 9 3 9 3 13 2
9 1 15 7 9 3 0 9 13 2
16 3 9 2 1 9 1 8 2 13 16 1 9 15 13 9 2
22 1 15 7 9 13 2 9 15 1 9 9 13 13 2 15 13 15 9 0 9 13 2
12 16 0 9 3 13 13 1 9 15 9 0 2
26 13 3 1 13 13 16 1 15 0 9 3 13 15 13 15 13 15 9 0 2 16 13 9 1 9 2
15 0 13 3 15 13 1 9 16 10 13 15 9 0 13 2
14 3 3 13 13 9 1 9 16 13 9 0 7 0 2
42 3 3 0 2 13 9 2 3 13 9 1 15 13 9 2 15 13 1 9 9 1 9 0 2 7 13 9 1 15 13 0 9 2 15 1 15 9 3 13 0 9 2
23 16 3 0 9 1 15 15 13 13 9 0 2 15 9 3 13 1 9 16 15 13 13 2
12 7 15 9 0 13 10 9 2 16 13 4 2
12 3 9 0 3 13 13 1 9 16 15 13 2
11 1 15 13 13 16 3 13 1 15 13 2
6 15 0 1 13 4 2
2 3 2
18 10 15 15 13 15 13 1 15 16 13 13 2 13 1 9 9 15 2
15 7 0 9 3 13 15 9 1 9 2 16 1 13 4 2
7 7 10 9 13 10 9 2
14 3 9 10 3 13 13 15 9 0 1 15 15 13 2
2 0 2
24 10 15 1 15 9 13 9 1 9 7 13 0 9 2 7 13 15 9 9 2 7 9 9 2
17 15 7 13 15 9 0 2 13 9 13 9 7 13 0 9 13 2
8 15 1 15 13 3 13 0 2
13 3 13 16 13 7 15 9 9 2 7 9 9 2
30 7 16 15 13 1 9 0 2 15 3 13 13 15 9 9 2 16 3 13 4 16 9 9 3 13 15 1 9 15 2
8 13 3 16 13 9 9 0 2
9 7 3 9 13 13 1 9 0 2
6 15 0 1 13 4 2
2 3 2
20 15 13 15 1 9 15 9 0 2 3 13 15 9 2 7 0 9 1 9 2
19 0 3 13 9 13 9 9 1 9 2 3 7 13 9 9 16 13 9 2
7 3 9 3 13 9 9 2
26 7 16 1 9 13 15 1 15 13 9 0 2 13 16 15 13 15 15 13 9 0 15 9 7 9 2
11 3 15 3 13 2 13 9 9 1 9 2
18 15 7 2 3 9 1 9 2 13 15 0 9 2 16 1 13 4 2
20 13 3 16 1 0 9 15 13 13 15 13 15 9 0 2 16 9 13 9 2
8 16 9 3 13 1 15 9 2
14 1 15 7 1 9 13 16 9 3 13 1 15 9 2
20 3 10 15 13 1 15 9 2 13 15 1 15 1 15 9 9 13 1 9 2
13 15 3 13 1 9 15 3 13 1 15 15 9 2
11 15 7 1 9 13 0 2 16 13 4 2
9 0 13 3 9 13 1 15 9 2
2 0 2
17 16 9 13 1 9 2 7 13 1 9 9 2 7 1 9 9 2
6 1 9 9 3 13 2
11 9 3 3 13 13 0 9 7 0 9 2
19 1 9 3 9 13 3 13 2 16 9 15 13 9 2 3 13 15 9 2
25 15 10 9 13 9 10 2 7 3 3 4 13 1 15 2 15 13 3 13 2 16 13 1 13 2
6 9 7 13 15 9 2
7 3 3 13 1 15 9 2
2 3 2
15 15 13 1 9 1 9 13 1 15 15 1 15 9 13 2
7 15 9 1 0 3 13 2
23 13 7 10 15 13 1 15 9 2 1 9 9 13 16 1 10 9 1 15 15 13 13 2
11 9 3 15 1 9 13 13 1 9 9 2
7 15 7 1 9 0 13 2
7 9 3 1 9 3 13 2
2 0 2
9 15 13 1 9 1 9 10 9 2
7 9 3 13 1 15 13 2
8 7 9 9 13 15 10 9 2
19 1 15 3 13 15 1 9 2 16 3 9 13 9 2 15 13 15 9 2
9 13 3 16 9 3 13 1 9 2
15 16 7 9 3 13 13 9 2 13 1 9 1 15 9 2
15 16 9 13 9 2 13 9 15 13 1 15 13 1 9 2
36 15 7 9 13 9 2 3 3 16 9 13 1 9 9 2 16 3 9 13 3 1 9 9 2 7 13 9 13 1 15 15 13 1 9 9 2
23 15 7 13 13 15 13 1 15 15 13 1 9 2 16 9 13 1 9 15 1 15 13 2
8 7 3 1 15 9 13 13 2
8 13 3 16 9 3 13 9 2
13 3 1 15 1 9 13 16 9 3 13 1 9 2
19 1 15 3 13 16 9 13 3 13 2 16 10 9 13 1 9 7 9 2
25 13 3 16 3 13 9 1 15 13 2 16 1 9 2 16 9 9 13 9 15 1 15 13 9 2
36 13 7 15 13 16 2 16 9 9 9 0 13 3 13 2 16 9 3 13 9 2 9 3 13 1 9 15 13 2 7 3 13 1 9 9 2
21 3 9 13 9 1 15 2 15 9 13 13 2 1 15 13 4 15 3 13 9 2
17 7 1 15 13 13 1 13 16 1 9 9 3 13 9 1 15 2
22 1 15 3 15 13 9 3 13 13 9 2 16 3 13 4 16 9 3 13 9 9 2
9 0 7 1 15 16 13 1 15 2
9 16 15 3 13 13 16 9 3 2
13 13 3 9 1 15 1 15 16 3 13 1 15 2
5 15 13 9 0 2
21 15 7 13 9 9 13 2 16 3 9 3 13 15 13 9 2 7 15 3 13 2
20 13 3 16 9 9 13 15 9 2 16 9 13 9 15 13 13 3 1 9 2
29 9 7 9 1 9 13 2 16 9 9 1 9 2 7 3 1 9 9 13 16 13 9 15 13 13 3 1 15 2
6 15 7 9 3 13 2
8 3 3 13 9 16 10 9 2
10 3 13 16 15 9 13 1 9 9 2
17 7 3 7 1 15 9 2 1 13 4 15 3 13 1 9 9 2
8 16 9 3 13 9 0 10 2
18 1 15 7 13 15 9 15 13 9 15 15 13 16 9 0 15 9 2
11 3 9 15 13 1 9 9 7 9 9 2
15 0 7 9 7 13 9 9 7 9 9 2 16 13 4 2
13 0 13 3 9 9 15 13 15 0 15 9 13 2
2 3 2
16 9 1 3 3 13 1 16 13 9 2 16 1 15 10 13 2
43 16 3 9 13 1 3 2 13 16 7 15 9 13 1 15 9 13 2 3 16 9 0 13 0 9 1 9 2 7 16 9 13 1 15 16 15 9 0 9 1 9 13 2
24 7 0 15 13 0 2 16 9 3 13 13 15 9 1 9 15 9 13 9 2 16 13 4 2
17 13 3 16 9 1 15 13 16 13 0 9 2 15 13 9 9 2
17 9 7 0 3 13 15 9 2 7 13 15 9 2 16 13 4 2
15 16 16 9 0 13 0 9 10 2 13 10 0 13 12 2
2 0 2
9 9 0 0 13 15 15 13 9 2
10 9 7 1 15 9 13 15 3 9 2
17 9 3 13 13 9 13 2 7 0 9 2 15 13 15 13 9 2
30 16 3 9 0 13 9 15 9 2 13 16 9 2 15 13 10 9 2 13 15 9 2 7 3 3 13 13 1 15 2
6 15 0 1 13 4 2
2 3 2
40 15 13 0 0 2 3 13 15 1 0 16 0 9 2 16 9 3 13 15 1 9 7 9 7 15 9 16 9 2 15 13 9 9 13 1 10 13 7 13 2
8 9 3 13 15 0 13 9 2
24 15 13 16 1 9 7 9 13 0 9 2 3 15 9 0 2 7 9 0 2 7 15 9 2
18 0 16 0 7 15 9 0 13 15 1 10 9 13 16 1 9 0 2
19 16 3 9 13 9 0 2 9 3 13 15 9 16 15 13 1 9 3 2
17 13 7 4 1 9 13 15 3 0 1 9 2 7 1 9 9 2
9 3 13 3 9 15 9 0 10 2
2 3 2
16 9 1 15 13 13 9 1 9 2 7 9 9 1 3 9 2
20 3 3 9 9 13 9 7 9 9 2 16 16 9 13 9 7 9 3 9 2
17 13 3 16 15 9 3 13 9 2 3 13 13 15 15 9 13 2
15 16 3 9 13 10 9 9 0 2 13 16 13 9 9 2
14 15 13 0 2 1 15 13 0 2 16 1 13 4 2
2 3 2
9 13 16 9 15 9 13 1 0 2
8 3 3 13 13 9 7 9 2
14 16 3 13 2 13 16 9 13 15 9 1 0 13 2
12 7 3 15 0 13 2 7 15 9 0 13 2
39 16 0 9 2 1 12 13 9 10 13 1 9 13 2 13 16 9 15 13 13 2 3 13 0 9 2 7 0 9 13 2 15 3 13 9 2 7 9 2
19 16 7 15 9 0 13 2 13 16 13 1 15 2 15 13 1 9 9 2
9 3 15 9 3 9 7 9 13 2
7 7 3 13 15 13 0 2
30 15 3 9 0 9 13 2 16 13 9 13 7 13 2 16 13 9 12 2 7 15 1 10 13 2 16 8 12 13 2
15 16 3 9 10 2 3 13 15 10 2 3 7 1 10 2
27 15 3 13 15 9 13 15 7 9 2 15 0 9 2 3 9 2 9 7 9 13 2 16 13 8 12 2
20 16 3 9 13 9 10 2 3 3 13 0 9 13 9 2 16 9 13 9 2
10 15 7 9 12 13 15 13 13 9 2
7 0 13 15 9 9 13 2
17 13 3 1 9 9 2 12 8 8 8 2 9 10 13 0 9 2
23 1 15 13 13 15 9 0 10 9 9 13 2 3 13 15 9 15 9 0 13 3 13 2
21 3 16 9 13 10 9 0 2 3 13 1 10 2 7 1 10 2 3 15 10 2
19 1 3 9 1 10 13 2 13 1 10 9 1 10 13 7 1 10 13 2
23 1 15 0 16 13 16 9 13 9 10 2 13 16 1 9 1 10 15 0 9 9 13 2
41 15 3 15 13 9 3 13 13 2 13 1 12 8 1 8 8 2 16 15 9 7 9 7 15 9 13 1 9 15 2 16 13 13 1 9 7 9 9 1 9 2
12 0 15 15 1 15 9 13 2 13 9 9 2
52 16 3 15 15 0 13 1 9 13 7 13 2 13 0 9 2 15 15 13 9 2 3 13 15 9 0 2 7 9 0 10 2 3 13 16 15 15 0 13 7 0 1 9 13 3 13 2 7 1 9 13 2
15 3 3 9 13 13 1 0 9 2 16 1 15 9 13 2
13 16 3 13 0 1 9 2 3 3 1 9 9 2
20 3 16 9 15 9 13 13 2 9 3 13 2 7 0 13 1 10 15 9 2
28 0 7 9 13 1 9 3 0 1 9 2 7 3 1 9 9 2 7 0 1 9 2 7 3 1 9 9 2
26 3 1 15 15 16 9 2 3 13 7 13 13 2 3 13 13 16 9 3 13 9 0 2 7 0 2
16 3 1 15 15 10 9 1 10 15 13 16 15 15 13 13 2
22 3 9 1 9 1 9 13 16 9 0 1 15 9 10 9 1 15 13 7 3 13 2
13 0 15 15 1 15 9 13 2 13 0 9 9 2
27 16 3 9 1 9 9 13 2 13 15 15 1 0 9 13 15 15 13 1 15 2 9 13 2 3 0 2
14 3 3 13 1 0 13 1 9 15 15 13 1 15 2
27 1 15 3 15 13 9 2 16 3 13 15 15 1 15 0 13 2 3 3 9 0 2 16 9 15 13 2
10 9 7 9 13 16 9 15 9 0 2
43 0 3 15 15 1 15 13 13 2 13 9 13 15 13 9 1 10 9 13 2 3 13 16 3 3 13 1 9 3 15 9 2 7 16 9 9 15 15 9 10 9 13 2
14 3 3 0 13 13 9 1 9 2 7 9 1 9 2
8 16 9 3 13 9 15 9 2
20 13 3 16 9 3 13 9 10 2 0 13 13 16 9 3 13 15 9 9 2
18 3 0 9 3 13 13 15 9 15 3 13 15 9 2 16 13 4 2
13 15 7 13 15 9 0 2 3 13 15 16 9 2
9 0 13 3 9 13 15 15 9 2
2 0 2
11 9 9 3 13 15 9 2 7 13 9 2
6 9 7 13 15 9 2
7 3 3 13 9 9 9 2
2 3 2
17 1 13 9 7 9 13 15 13 2 15 13 15 9 9 7 9 2
8 9 7 13 1 9 9 15 2
7 1 9 7 15 13 9 2
10 0 13 3 9 13 9 13 15 9 2
2 3 2
15 15 1 15 13 9 2 0 13 15 15 13 9 1 15 2
10 10 7 9 15 9 13 9 1 15 2
18 1 3 9 13 9 0 2 3 0 13 9 2 3 13 13 15 9 2
2 3 2
10 15 15 13 13 1 9 9 2 3 2
18 16 9 13 9 15 0 2 1 15 13 0 13 2 9 13 13 15 2
9 7 13 15 13 13 7 3 13 2
6 15 3 1 15 13 2
12 15 7 13 3 2 3 13 9 9 1 15 2
16 13 3 1 13 15 13 15 0 13 2 15 13 15 9 9 2
16 7 3 9 2 15 13 0 13 2 3 13 9 9 13 15 2
9 13 7 15 9 0 13 9 9 2
13 15 3 13 2 15 9 13 13 1 9 9 9 2
16 16 3 13 15 13 13 7 13 2 3 13 0 7 0 13 2
25 9 3 9 9 9 13 1 15 9 0 3 0 2 15 3 13 9 9 13 15 3 15 9 15 2
7 15 7 9 9 13 9 2
5 13 3 1 9 2
9 13 4 9 10 1 9 2 9 2
4 7 9 12 2
7 13 9 13 7 15 13 2
9 0 9 9 15 13 7 0 9 2
50 3 3 0 9 13 2 15 13 9 13 9 9 7 3 9 15 9 2 7 1 15 9 2 9 13 2 13 15 9 13 9 2 3 9 9 2 7 9 9 2 16 9 13 0 3 9 9 7 9 2
16 15 13 2 13 13 16 9 7 9 15 3 0 0 9 13 2
27 9 3 13 2 1 12 8 2 16 15 9 13 9 13 9 9 2 3 9 16 3 13 9 13 9 9 2
4 1 9 0 2
31 16 7 15 15 13 7 13 2 9 13 16 15 15 3 13 2 9 3 15 3 13 15 16 10 9 2 13 0 9 9 2
12 7 13 0 9 2 15 3 13 15 9 9 2
11 10 3 9 15 9 13 15 1 10 9 2
19 15 3 9 13 9 1 10 9 16 1 15 0 13 2 7 3 1 15 2
15 3 3 1 9 15 9 13 9 2 13 10 9 1 9 2
25 3 9 1 16 10 9 13 1 15 0 9 9 0 7 0 2 13 13 1 15 0 7 0 0 2
20 3 16 15 13 15 13 15 9 13 2 15 15 9 13 13 15 15 9 13 2
30 7 9 15 13 10 9 2 13 13 1 15 13 9 2 16 2 16 13 15 9 13 2 15 15 1 9 9 13 13 2
28 3 15 0 15 1 9 9 13 1 9 13 9 2 15 15 1 9 10 13 2 7 3 3 1 15 13 9 2
21 9 3 2 15 13 10 9 2 16 1 13 4 2 13 9 1 15 9 15 9 2
11 3 13 3 13 15 9 15 15 9 13 2
23 16 7 10 9 7 9 13 9 1 16 13 2 3 10 9 13 15 1 16 0 3 13 2
30 9 7 2 16 13 9 0 2 3 1 15 0 13 3 9 2 16 1 9 1 15 13 15 9 2 13 1 3 9 2
7 1 9 3 10 9 13 2
5 13 3 0 9 2
15 15 0 15 3 13 2 3 13 0 1 9 15 9 0 2
20 3 3 15 13 9 1 10 15 13 2 7 13 9 1 15 0 9 7 0 2
2 3 2
10 10 0 1 15 9 0 13 16 13 2
9 9 3 13 1 9 7 1 9 2
7 3 0 9 13 13 9 2
8 13 4 7 9 13 0 9 2
4 13 3 9 2
2 0 2
17 15 9 13 16 13 9 2 0 7 1 16 13 9 1 9 9 2
16 15 3 15 15 9 13 9 7 13 9 0 2 13 9 13 2
5 15 7 9 13 2
4 13 3 9 2
2 0 2
9 15 13 16 1 16 13 1 9 2
8 9 3 13 9 9 1 9 2
18 0 13 3 9 15 1 9 13 2 13 1 0 9 16 13 9 9 2
25 0 13 3 9 9 0 13 16 13 9 9 13 2 15 16 9 13 13 1 9 15 1 15 13 2
30 1 9 7 9 0 13 9 1 12 0 15 9 13 2 16 1 13 13 2 1 15 13 10 9 2 16 1 13 13 2
26 13 3 15 9 13 1 15 9 15 2 13 1 9 0 13 16 13 1 9 15 2 3 7 1 0 2
5 13 3 9 9 2
2 3 2
40 1 15 9 13 15 9 1 9 15 2 1 15 10 15 13 15 9 13 2 16 1 15 15 13 3 7 0 9 13 2 15 1 9 10 9 3 7 0 13 2
15 16 0 13 13 9 1 10 9 2 7 0 1 10 9 2
19 15 7 15 13 9 10 9 3 13 13 15 16 9 2 15 13 10 9 2
10 15 3 15 13 9 15 15 9 13 2
7 15 3 13 10 0 9 2
41 15 13 16 2 1 13 9 0 13 9 7 9 2 13 4 15 1 9 2 15 13 15 10 9 2 16 13 8 12 2 1 15 13 13 1 15 10 9 9 13 2
11 9 3 2 1 12 8 1 8 8 13 2
19 9 3 15 9 13 13 2 7 0 7 0 15 9 1 15 13 7 13 2
19 13 3 13 16 9 9 13 13 3 13 16 9 9 3 1 15 9 13 2
12 15 3 13 3 4 2 7 9 13 13 13 2
52 7 16 10 15 13 2 1 9 1 9 13 4 7 1 3 9 1 9 16 13 4 2 3 0 9 13 13 2 3 0 13 2 16 9 0 13 1 9 13 2 16 15 1 3 9 13 2 7 13 9 0 2
28 1 15 3 9 9 9 13 3 0 15 13 13 1 9 0 2 7 15 3 15 13 1 9 0 1 10 9 2
12 7 3 9 9 13 13 2 1 15 8 12 2
10 13 9 16 7 9 10 0 9 13 2
4 1 9 9 2
18 1 15 7 3 1 9 13 9 1 9 13 7 3 13 2 13 13 2
24 9 3 1 10 9 13 3 13 1 15 1 9 7 9 2 0 13 3 15 1 15 9 13 2
18 1 9 3 9 13 16 9 15 0 13 1 15 13 1 16 9 13 2
24 3 9 9 1 9 13 13 3 0 2 7 1 15 9 7 15 9 2 9 15 9 0 13 2
13 9 3 1 9 9 9 13 13 1 16 9 13 2
34 3 13 16 9 1 9 13 0 9 13 1 9 0 9 2 1 15 9 1 15 9 13 2 9 15 9 0 13 2 16 3 12 9 2
15 7 3 9 10 15 0 0 13 1 15 10 9 0 13 2
23 1 15 3 3 10 0 13 2 16 3 9 3 15 9 13 9 7 3 15 1 9 13 2
20 3 3 7 9 10 9 9 13 2 7 1 15 1 10 9 13 7 9 3 2
20 7 3 13 16 0 9 3 9 1 15 7 9 13 2 16 1 13 8 12 2
8 13 9 1 9 7 9 10 2
9 3 9 13 2 1 15 9 12 2
12 15 3 0 13 9 2 7 15 9 13 15 2
4 7 1 9 2
7 9 2 15 0 13 15 2
15 15 7 9 9 13 2 15 1 12 8 1 8 8 13 2
7 15 0 13 9 7 0 2
18 0 3 2 1 9 15 15 3 13 9 0 2 15 1 15 13 13 2
11 0 7 2 1 16 13 13 0 10 9 2
13 1 3 15 9 13 13 9 9 0 16 1 0 2
11 0 3 15 13 15 15 13 9 7 9 2
33 16 3 15 15 1 9 9 13 2 1 9 15 1 15 13 9 13 2 15 1 15 9 13 2 9 3 0 13 2 3 7 9 2
8 7 3 9 13 15 9 13 2
7 3 7 9 0 0 13 2
11 3 7 3 13 13 9 13 15 9 13 2
9 3 7 13 13 9 9 0 13 2
17 16 7 9 13 10 9 13 0 2 15 3 10 9 0 0 13 2
10 0 3 0 0 13 16 9 9 13 2
18 3 9 9 1 9 13 7 3 13 7 15 1 15 13 3 0 13 2
15 9 7 13 1 9 3 15 13 0 2 3 7 1 0 2
11 3 3 9 9 13 2 7 3 1 0 2
7 15 9 1 9 13 13 2
28 1 15 3 13 13 15 1 9 13 7 3 13 13 2 15 7 1 15 3 13 2 15 3 3 7 15 9 2
43 16 3 10 9 9 13 1 9 13 7 1 15 9 13 2 15 9 0 9 1 9 13 2 1 9 13 7 1 15 9 2 16 13 9 2 9 2 9 2 7 15 3 2
41 15 0 9 3 9 13 1 9 0 9 2 1 9 13 3 13 16 1 9 7 9 2 1 15 15 13 12 9 15 13 13 2 16 15 9 13 9 1 9 9 2
17 3 7 13 10 9 13 1 13 9 9 13 2 16 9 7 9 2
10 3 15 9 13 0 9 9 7 9 2
14 0 3 15 9 9 9 13 15 1 0 9 9 13 2
9 3 1 9 13 3 13 16 0 2
28 15 0 3 9 13 1 9 9 15 9 13 2 1 0 9 13 2 16 0 9 2 0 9 2 7 15 3 2
20 13 7 15 13 9 9 1 9 13 2 3 1 15 1 15 13 9 4 13 2
12 3 3 1 9 13 2 10 9 1 9 13 2
10 3 9 9 13 15 9 15 9 13 2
35 9 7 10 2 1 9 13 9 13 2 15 9 3 13 15 1 9 0 13 2 1 15 15 13 9 7 13 9 2 1 9 7 9 9 2
31 9 0 1 15 9 13 3 0 2 7 0 2 3 3 0 2 13 7 9 13 3 0 2 7 3 0 2 3 9 13 2
13 3 9 10 2 15 13 16 0 2 13 1 9 2
16 15 0 16 0 2 13 3 16 15 13 2 7 16 15 13 2
39 7 3 1 10 9 1 15 13 2 3 1 9 13 2 9 13 2 15 9 3 13 2 16 9 13 15 13 9 9 13 2 16 13 1 9 9 7 9 2
12 3 9 13 16 3 0 2 9 7 16 9 2
21 7 3 1 15 15 9 9 13 13 2 7 0 3 1 15 1 15 13 9 13 2
16 13 3 2 16 9 13 2 3 9 7 13 1 9 7 13 2
7 13 3 2 1 9 9 2
7 13 0 2 1 13 9 2
49 9 7 9 15 1 9 13 9 13 2 1 9 1 15 13 13 3 13 16 7 1 9 2 16 1 13 9 0 7 0 2 7 3 1 9 15 1 15 2 16 1 13 0 9 2 7 0 9 2
28 3 3 1 9 13 13 15 13 2 7 15 3 13 2 7 15 15 15 13 1 15 2 16 1 1 13 13 2
12 16 0 9 7 9 9 0 0 9 3 13 2
19 1 13 3 13 13 16 0 9 7 0 9 13 1 9 15 9 3 13 2
19 3 3 10 9 1 9 15 13 9 13 13 16 9 1 10 9 0 13 2
14 15 3 9 1 10 9 13 9 2 16 9 1 9 2
19 9 7 3 16 0 13 1 9 9 2 9 1 15 13 3 15 0 13 2
27 1 15 3 9 9 0 13 2 3 0 16 9 13 2 7 16 9 1 15 15 13 2 13 15 0 9 2
22 1 15 7 9 1 15 9 13 9 2 13 7 0 15 9 1 9 9 2 16 9 2
19 7 3 9 7 9 2 15 1 9 13 9 0 2 9 13 1 12 9 2
22 3 7 10 9 2 15 9 15 1 0 9 13 2 9 1 12 15 9 13 13 0 2
20 15 3 9 3 13 15 1 10 9 2 1 15 15 13 13 2 16 13 4 2
32 3 3 0 9 13 3 0 1 15 16 9 13 2 7 16 2 1 16 0 13 2 9 15 2 15 0 15 13 2 15 13 2
25 3 7 13 9 2 16 9 13 2 16 1 9 9 13 9 13 13 2 1 15 9 1 9 13 2
21 13 7 9 9 16 9 1 9 2 1 9 2 7 15 3 2 16 7 15 9 2
14 15 7 0 13 13 1 9 0 7 1 9 0 0 2
18 9 3 0 9 13 10 15 9 0 0 9 13 2 7 3 15 0 2
25 9 3 2 3 13 9 2 3 15 12 0 13 13 2 1 15 13 9 9 3 13 16 1 0 2
16 9 3 0 1 10 15 13 1 15 0 1 15 9 9 13 2
26 3 3 7 9 1 12 0 10 9 0 9 13 2 15 9 15 2 3 0 0 2 1 15 0 13 2
9 1 15 13 9 0 9 9 13 2
33 16 3 15 3 13 13 0 16 1 9 13 1 15 2 13 16 9 15 9 15 13 2 0 13 2 16 7 9 1 9 13 0 2
20 16 7 15 9 16 13 13 13 7 15 9 0 13 2 12 9 3 15 13 2
12 15 13 15 15 15 1 9 13 2 8 8 2
11 1 9 15 13 9 12 7 9 15 12 2
10 16 15 1 9 7 9 15 0 13 2
15 1 15 7 13 16 15 1 9 7 9 15 13 0 13 2
27 3 9 15 3 13 9 1 9 0 15 1 15 9 13 2 9 1 15 9 13 1 0 9 13 3 13 2
13 3 3 0 13 0 9 1 9 13 2 7 9 2
27 9 15 9 13 9 2 9 1 9 0 9 3 13 2 1 13 7 0 13 15 1 9 0 7 0 13 2
13 13 3 16 1 9 7 9 15 15 0 13 13 2
2 0 2
23 16 15 9 1 9 9 13 2 9 9 0 3 13 16 1 15 13 9 15 9 9 13 2
24 3 3 0 13 9 15 13 1 9 2 7 1 9 2 1 15 16 9 9 13 9 0 3 2
19 9 7 15 2 3 16 3 0 9 13 2 3 3 13 1 15 9 13 2
24 3 15 13 1 9 15 3 13 15 13 0 2 16 1 13 13 2 15 1 15 9 3 13 2
12 0 13 3 15 0 1 9 7 9 15 13 2
2 3 2
22 10 15 1 0 0 13 2 7 13 9 2 7 9 2 7 9 2 7 9 7 0 2
34 1 9 7 15 13 16 9 7 16 9 2 16 1 13 4 2 7 3 7 16 9 2 7 3 16 9 2 15 1 9 7 9 13 2
24 7 15 15 13 13 2 16 1 13 4 2 7 3 15 1 15 13 7 16 9 7 16 0 2
7 3 0 1 9 9 13 2
11 13 3 15 1 9 7 9 15 0 13 2
2 3 2
15 15 0 1 0 13 2 15 15 1 0 1 9 0 13 2
13 9 7 7 1 9 7 1 9 13 13 15 0 2
10 15 3 0 1 9 7 9 15 13 2
2 0 2
16 10 15 1 0 13 0 2 1 9 15 15 13 1 15 13 2
10 3 9 13 13 9 2 7 9 9 2
8 1 9 7 15 13 1 9 2
20 3 10 15 13 13 1 9 13 2 7 3 0 13 7 3 1 10 9 9 2
11 13 3 15 1 9 7 9 15 0 13 2
2 3 2
15 15 13 1 15 1 0 7 0 2 0 13 0 3 13 2
17 3 0 1 9 0 13 2 16 9 1 9 9 1 16 13 9 2
24 16 3 13 0 9 1 9 7 9 2 13 16 9 3 13 1 9 9 1 16 1 9 13 2
5 15 13 13 0 2
37 15 7 1 9 7 9 15 13 15 9 2 7 1 0 7 0 2 1 1 9 10 13 0 2 13 3 9 3 15 9 2 7 0 3 15 9 2
22 1 15 7 9 13 1 9 2 16 9 13 9 3 16 13 15 9 2 7 9 13 2
12 0 13 3 15 1 9 7 9 15 0 13 2
12 16 3 10 9 13 1 9 7 9 0 0 2
27 1 13 3 13 16 3 15 1 9 7 9 15 13 2 1 0 9 13 2 16 15 15 13 1 9 0 2
30 3 1 15 15 13 1 9 0 2 15 9 7 9 13 12 1 15 2 7 3 1 9 13 16 12 9 0 9 13 2
12 3 3 9 13 12 13 15 13 9 1 15 2
13 3 7 3 13 1 9 15 1 9 13 7 9 2
16 13 3 1 3 9 9 9 9 7 13 2 16 1 13 13 2
13 3 3 1 0 9 15 1 9 7 9 15 13 2
2 0 2
16 16 13 0 9 2 15 9 1 9 13 2 7 0 9 9 2
15 9 7 1 9 13 15 9 9 2 16 1 1 13 13 2
11 13 3 16 3 13 1 9 1 0 9 2
2 3 2
19 16 12 1 0 1 0 9 13 2 1 12 15 3 13 13 1 9 15 2
13 3 9 9 3 13 1 9 2 7 1 9 9 2
18 1 15 7 15 1 9 15 13 1 0 9 13 2 16 1 13 13 2
13 3 3 1 0 9 13 3 1 9 7 15 9 2
2 3 2
6 9 9 9 9 13 2
22 16 3 15 13 1 9 7 9 16 0 0 2 15 9 13 13 13 1 9 1 9 2
9 15 0 13 1 10 13 1 0 2
2 0 2
15 3 15 9 1 15 13 16 1 15 9 15 1 15 13 2
33 7 16 9 13 1 9 7 9 3 0 2 15 1 15 9 1 9 13 2 1 9 15 9 13 13 15 0 1 16 1 9 13 2
21 3 3 13 7 13 1 9 16 9 13 9 2 0 2 7 16 15 15 3 13 2
48 16 7 13 16 1 3 9 0 1 9 13 15 3 13 2 16 3 15 9 13 13 16 3 13 1 9 9 0 7 3 1 15 2 1 0 13 16 0 1 9 7 9 13 13 1 9 0 2
7 7 3 3 13 0 0 2
11 16 15 15 13 1 9 7 9 13 0 2
35 3 3 1 13 13 16 15 15 1 9 7 9 15 13 2 13 7 0 7 0 2 7 0 2 15 13 2 1 9 7 9 1 15 12 2
5 15 3 0 13 2
38 12 9 2 1 16 0 13 9 1 15 12 2 16 1 9 1 12 9 9 13 0 16 15 13 2 9 16 15 0 2 9 16 0 2 9 16 9 2
46 15 9 2 1 16 12 13 9 7 9 2 3 1 15 15 2 7 1 12 15 2 16 9 1 9 7 9 13 1 16 9 1 9 9 13 2 3 16 9 7 9 1 15 0 13 2
26 3 3 9 1 9 7 9 15 3 13 0 1 0 9 2 13 3 15 9 13 0 2 7 9 0 2
20 1 3 7 0 9 9 13 15 1 9 7 1 9 3 2 3 0 3 15 2
13 3 9 9 13 9 9 2 16 13 9 0 9 2
50 16 3 15 15 13 0 1 9 2 13 3 9 0 2 15 13 0 7 1 9 9 7 1 9 9 2 16 9 13 0 9 7 9 2 16 9 13 9 9 2 7 9 2 16 9 1 9 9 13 2
19 7 3 9 13 0 1 9 16 1 9 7 1 9 9 7 1 9 9 2
63 16 0 15 15 13 0 1 9 2 13 0 1 9 2 3 1 0 3 13 15 9 1 9 7 1 9 9 2 16 9 13 15 13 1 0 2 0 13 0 9 15 13 1 9 2 16 9 9 2 7 16 15 9 1 9 13 2 3 3 1 9 13 2
20 7 3 13 16 0 13 0 9 9 2 7 9 13 1 0 0 1 9 9 2
35 3 3 2 16 1 9 15 1 9 9 13 2 9 9 1 9 7 9 15 13 1 0 13 1 9 1 10 9 2 7 9 9 1 0 2
8 3 7 13 13 1 10 13 2
10 16 0 9 13 1 9 3 13 0 2
26 13 3 1 13 16 2 16 9 1 9 13 15 9 13 2 3 3 13 0 2 16 3 13 9 15 2
35 3 16 0 9 12 0 9 15 9 13 13 1 9 0 2 3 9 10 1 0 9 15 0 13 2 16 1 0 9 9 1 15 13 13 2
36 7 3 1 12 2 9 10 0 13 3 13 0 7 0 2 16 15 0 9 0 3 13 16 15 1 9 0 15 13 13 2 16 1 13 4 2
12 1 7 0 9 0 9 9 13 15 9 13 2
22 7 3 2 1 3 1 15 9 13 2 13 15 3 13 0 2 16 9 3 12 13 2
18 3 3 13 15 9 9 2 1 9 1 0 9 9 16 9 13 13 2
8 15 9 10 1 9 9 13 2
26 1 15 3 0 13 16 9 10 1 9 0 3 1 0 9 13 13 7 13 2 16 9 3 13 0 2
27 16 3 9 10 1 9 9 1 0 9 13 2 16 13 4 2 13 3 15 15 10 15 13 3 12 13 2
20 3 3 9 9 15 13 9 13 13 2 16 7 9 9 2 16 15 0 13 2
42 7 3 9 9 13 1 9 0 2 15 13 9 9 2 1 13 2 9 13 0 7 9 2 3 16 16 15 9 1 9 13 2 1 9 13 2 9 0 1 9 13 2
49 7 1 15 9 3 9 10 9 1 9 13 1 15 9 9 2 9 13 2 16 1 13 2 9 13 1 9 2 16 7 3 13 15 9 2 15 13 9 2 7 15 9 2 15 13 1 9 13 2
5 16 9 13 0 2
13 1 9 7 0 2 15 13 2 9 15 13 13 2
12 15 3 15 15 0 13 2 13 0 9 15 2
14 3 9 13 15 15 0 13 13 7 9 15 0 13 2
6 9 7 13 9 15 2
16 3 3 15 9 13 16 13 0 9 2 16 13 1 12 9 2
10 1 15 3 15 0 13 15 9 13 2
12 7 3 13 16 15 10 9 13 16 0 9 2
7 13 4 7 9 13 9 2
4 13 3 0 2
2 3 2
13 13 4 1 13 15 0 13 0 2 15 9 13 2
7 13 7 16 13 3 0 2
5 16 13 16 13 2
13 9 3 2 1 13 0 13 0 2 13 0 13 2
15 13 7 0 15 2 7 16 13 0 2 7 16 13 0 2
7 15 0 13 16 13 0 2
16 3 13 9 3 13 1 15 2 7 1 16 13 15 9 9 2
6 9 0 13 1 15 2
12 0 3 13 2 15 9 13 2 13 0 0 2
2 3 2
15 9 13 15 10 13 2 16 9 0 9 13 2 12 9 2
9 10 7 13 13 9 1 10 9 2
12 15 13 1 15 16 15 1 9 10 13 9 2
31 13 3 9 9 9 13 2 3 7 1 9 9 1 9 13 9 2 15 13 9 13 2 3 1 9 13 2 1 12 0 2
14 9 7 13 9 9 3 1 9 2 16 1 13 4 2
5 13 3 0 0 2
2 0 2
8 9 9 7 9 1 9 13 2
14 15 3 13 7 1 15 9 9 2 7 1 15 9 2
10 0 3 9 15 13 9 7 9 15 2
9 15 7 1 15 13 16 9 13 2
9 13 7 9 7 9 1 15 13 2
19 3 7 9 9 13 15 16 0 13 13 2 16 13 1 9 1 12 9 2
10 9 0 9 13 1 15 16 13 0 2
4 15 13 9 2
7 15 3 13 13 1 13 2
10 1 15 13 9 13 0 15 7 9 2
6 15 7 9 9 13 2
16 13 3 4 1 16 15 13 9 13 2 16 1 15 9 0 2
5 13 3 0 0 2
7 15 13 15 1 9 13 2
10 16 0 9 9 15 15 13 13 9 2
5 7 8 12 13 2
11 0 13 9 13 1 15 2 9 13 15 2
6 16 9 13 15 9 2
11 1 15 7 13 13 16 9 13 10 9 2
9 13 3 9 1 15 13 9 15 2
19 7 9 3 0 13 9 9 2 7 13 15 10 9 2 16 1 13 4 2
9 13 3 15 9 2 3 3 0 2
2 3 2
10 9 15 13 9 15 2 16 13 4 2
25 9 7 0 9 3 13 1 15 13 1 15 2 7 16 15 1 15 9 13 2 16 1 13 4 2
17 9 3 9 3 13 15 13 10 9 2 7 10 9 13 10 9 2
2 3 2
12 15 9 15 3 13 10 9 2 0 13 0 2
17 15 7 1 9 13 2 15 1 15 13 2 1 15 9 13 9 2
23 15 7 1 0 3 13 0 13 2 16 1 9 0 3 13 1 0 2 0 3 13 9 2
6 9 7 9 9 13 2
26 13 3 13 1 15 9 0 2 15 3 0 13 0 1 9 1 15 15 2 7 13 1 9 10 0 2
5 15 7 9 13 2
6 13 3 9 10 9 2
2 3 2
12 15 15 13 13 15 13 2 15 7 9 15 2
11 15 3 13 9 13 2 9 7 9 13 2
10 7 9 13 15 9 2 16 13 4 2
9 3 13 3 0 0 2 7 0 2
2 0 2
11 10 0 10 9 7 15 15 13 12 13 2
12 3 2 16 13 15 7 15 2 3 9 13 2
10 9 7 13 3 0 2 16 13 4 2
10 3 15 13 0 3 13 15 16 15 2
5 13 3 10 9 2
12 1 15 3 13 16 15 15 9 13 10 9 2
6 1 15 13 8 12 2
6 15 0 16 0 9 2
8 16 1 9 3 13 13 9 2
13 1 15 7 0 13 16 1 9 3 13 13 9 2
32 9 3 7 9 2 7 10 15 1 9 13 2 15 1 15 13 13 2 16 15 15 13 7 9 13 15 1 9 7 9 13 2
39 15 3 13 15 13 12 9 13 2 3 15 13 2 16 15 13 9 13 13 0 7 0 2 15 7 9 10 9 9 13 2 16 15 0 1 15 13 13 2
13 9 7 13 9 2 3 0 0 2 16 13 4 2
10 3 13 3 1 15 13 15 3 9 2
10 7 3 9 1 15 3 13 3 13 2
2 0 2
29 15 15 13 13 9 15 9 2 15 3 13 3 13 16 13 2 16 9 3 13 13 9 7 9 16 9 13 13 2
11 7 0 9 13 15 9 2 16 13 4 2
18 3 9 2 15 13 9 13 2 1 15 9 13 3 13 16 13 13 2
13 15 13 0 2 1 13 0 2 16 1 13 4 2
2 3 2
20 1 9 13 10 9 2 15 0 1 15 13 13 2 16 13 1 9 1 13 2
14 16 3 9 1 15 13 2 3 13 0 2 7 0 2
12 3 7 9 1 15 13 13 16 13 9 15 2
13 15 3 9 13 2 15 9 13 2 16 13 4 2
15 1 9 7 3 13 13 15 0 13 2 16 3 1 9 2
8 9 3 1 9 13 3 13 2
2 3 2
5 9 9 13 13 2
7 9 7 9 1 9 13 2
6 3 9 9 1 9 2
21 9 7 7 9 1 9 2 15 13 0 9 2 13 3 13 2 16 1 13 4 2
8 1 9 3 9 13 3 13 2
2 3 2
8 9 13 15 1 16 13 9 2
10 3 0 13 1 16 13 13 1 9 2
10 3 9 7 9 13 2 7 9 13 2
6 9 7 9 13 9 2
8 15 7 1 9 13 3 13 2
4 3 7 9 2
2 3 2
16 16 9 13 15 1 10 13 2 3 9 15 9 13 16 3 2
15 15 7 13 15 1 9 0 9 2 13 0 7 1 9 2
27 9 3 1 15 13 0 7 1 9 1 16 13 15 9 2 16 13 15 13 0 1 15 15 1 9 13 2
21 9 7 13 3 13 2 7 15 13 13 1 15 0 7 1 9 2 16 13 4 2
8 9 3 1 9 13 3 13 2
6 15 3 0 9 13 2
6 13 3 0 0 9 2
12 9 9 13 2 7 9 1 15 3 13 15 2
5 7 1 9 12 2
10 13 1 9 9 2 7 1 0 9 2
7 16 9 13 10 9 9 2
11 13 3 1 13 16 9 13 10 9 9 2
11 9 3 15 13 9 15 2 16 13 4 2
19 9 7 2 1 13 0 9 2 10 9 10 9 9 13 2 16 13 4 2
7 10 3 9 10 9 13 2
7 7 3 13 10 9 9 2
2 3 2
30 15 1 9 13 0 2 3 13 15 16 16 13 15 9 15 15 1 9 13 2 16 9 13 13 16 15 9 9 13 2
17 7 9 13 0 1 9 2 10 0 15 1 9 2 16 13 4 2
12 3 15 13 0 16 16 13 15 9 0 9 2
7 13 3 15 9 10 9 2
2 3 2
33 1 15 0 13 1 9 2 9 7 9 13 1 15 16 13 0 2 13 16 15 13 0 7 16 13 9 2 7 16 13 1 9 2
11 9 3 0 13 1 15 10 9 9 13 2
9 15 7 9 13 2 16 1 13 2
7 13 3 9 10 9 9 2
15 15 13 16 9 2 10 9 9 13 2 13 2 9 12 2
6 15 13 15 10 9 2
9 7 8 12 2 13 1 0 9 2
8 13 15 10 9 0 1 15 2
6 16 9 13 0 9 2
10 1 15 7 13 16 9 13 0 9 2
17 3 9 0 13 15 9 0 2 16 9 9 13 0 16 9 12 2
11 9 3 15 7 9 13 9 7 9 9 2
23 7 0 9 13 1 10 15 16 0 9 1 0 2 1 13 10 9 9 2 16 13 4 2
6 13 3 15 0 9 2
2 3 2
16 15 15 1 9 13 2 0 13 16 15 15 4 1 9 13 2
17 7 9 13 0 1 10 9 2 15 0 1 9 2 16 13 4 2
6 13 3 15 0 9 2
2 3 2
15 15 13 0 1 15 9 13 9 15 15 13 1 15 9 2
6 9 3 0 13 9 2
12 1 9 7 10 13 9 9 2 16 13 4 2
6 13 3 15 0 9 2
2 0 2
16 16 0 13 15 13 0 9 2 3 0 13 15 13 9 9 2
30 7 9 13 0 9 9 2 16 1 15 7 9 7 9 9 13 13 2 7 15 15 1 10 9 13 2 16 13 4 2
6 13 3 15 0 9 2
8 15 13 15 13 12 8 12 2
7 3 13 0 16 13 9 2
5 16 9 13 12 2
12 15 7 13 2 0 13 9 3 13 16 12 2
9 3 3 0 13 13 12 0 9 2
11 15 3 1 9 13 2 1 12 3 13 2
10 9 7 13 0 9 2 16 13 4 2
5 9 3 13 12 2
2 3 2
12 13 4 9 13 3 9 2 15 15 9 13 2
12 16 3 13 0 9 2 13 13 0 3 9 2
5 15 7 13 0 2
31 3 16 15 15 13 15 9 2 7 15 9 13 2 15 13 1 15 16 15 13 0 9 2 3 13 1 15 1 3 13 2
7 0 13 3 0 9 13 2
2 3 2
15 15 0 13 12 13 2 0 13 1 12 13 16 1 0 2
9 7 9 9 13 16 0 13 13 2
14 3 3 9 9 0 13 9 15 13 1 9 1 9 2
10 0 7 10 13 13 1 12 0 9 2
7 3 13 3 13 0 9 2
2 0 2
12 0 13 12 9 0 7 0 1 0 9 13 2
21 3 2 16 3 13 2 15 15 13 9 9 2 7 10 15 13 9 12 9 9 2
13 15 3 13 1 0 9 2 9 3 13 0 0 2
15 16 7 3 3 13 2 15 15 13 3 13 3 3 3 2
11 1 15 13 16 9 3 13 0 7 0 2
10 9 3 0 7 12 13 1 12 9 2
35 9 3 15 3 3 13 2 0 13 13 2 16 13 1 9 9 2 1 15 9 0 1 9 13 7 1 9 13 2 9 7 0 1 0 2
14 7 0 9 13 12 7 0 2 16 1 9 13 4 2
8 3 13 15 9 0 13 12 2
2 3 2
10 9 0 13 1 0 16 1 10 9 2
23 3 13 1 15 9 0 2 15 0 9 13 13 2 1 10 15 13 13 0 3 0 13 2
24 7 10 9 0 9 13 13 1 12 0 2 1 15 3 13 15 0 15 15 9 13 1 15 2
19 3 1 9 0 15 13 9 0 9 2 3 13 15 15 3 13 1 15 2
6 15 7 9 9 13 2
7 3 13 3 16 12 9 2
2 0 2
32 10 0 13 1 3 2 9 15 1 3 13 1 9 15 1 15 12 2 16 9 9 9 1 3 13 1 9 15 9 1 9 2
26 3 16 15 0 1 9 15 13 2 3 13 13 1 0 9 1 16 13 0 2 16 1 15 3 13 2
22 7 13 13 1 0 13 2 16 3 13 13 16 12 9 13 1 15 1 16 13 0 2
29 7 3 7 9 0 1 3 13 1 9 2 7 13 13 1 15 12 0 13 2 15 1 9 15 13 10 15 13 2
35 10 7 9 15 9 13 13 1 3 2 1 16 15 1 15 13 16 9 9 13 1 0 2 7 15 1 9 0 2 16 1 1 13 13 2
14 7 15 13 1 9 2 1 13 3 7 1 0 9 2
12 3 15 15 9 3 13 16 12 9 7 9 2
8 7 1 15 9 3 13 15 2
13 3 13 3 16 12 10 9 9 2 15 9 13 2
2 3 2
16 16 13 12 15 15 13 13 2 13 16 13 1 9 9 13 2
14 13 3 16 13 1 15 15 13 12 3 2 7 15 2
10 7 3 13 7 15 7 15 13 13 2
14 15 7 9 13 13 2 1 15 2 16 1 13 4 2
10 0 13 3 13 0 15 15 13 13 2
6 7 3 7 0 9 2
2 0 2
25 15 1 15 13 2 1 15 13 13 1 9 13 2 7 13 1 9 9 13 15 9 2 7 3 2
23 16 3 13 2 3 13 15 0 2 16 10 15 13 9 15 13 1 9 15 2 13 9 2
6 3 15 9 13 9 2
12 7 3 9 15 15 13 13 2 7 15 15 2
25 16 9 15 2 1 15 9 13 13 9 15 2 16 1 1 13 13 2 9 13 13 9 15 9 2
7 7 9 13 13 1 15 2
6 3 15 13 15 9 2
7 7 3 3 13 1 15 2
20 16 7 9 15 9 13 15 15 2 16 3 15 15 13 2 15 9 3 13 2
11 7 16 15 9 13 2 9 13 3 13 2
19 3 2 16 13 15 15 2 15 12 15 13 13 2 3 13 12 7 12 2
9 3 9 0 15 13 13 1 15 2
8 7 3 15 13 13 1 15 2
47 16 7 15 1 15 13 13 0 1 9 13 13 2 7 15 13 16 15 13 1 9 9 13 2 16 13 13 1 9 9 2 7 15 13 16 9 13 13 1 15 2 16 9 13 1 0 2
28 16 0 9 2 13 16 2 3 13 9 13 2 13 15 15 1 15 9 13 2 16 15 13 9 2 13 13 2
16 7 3 2 1 9 13 13 9 13 2 1 15 13 3 13 2
11 16 7 0 9 2 15 3 13 3 13 2
18 3 9 13 9 3 13 9 9 2 7 1 15 13 9 9 1 9 2
21 9 3 9 0 13 1 9 0 2 7 3 13 13 9 9 16 13 0 7 0 2
19 3 3 15 13 9 13 3 1 9 1 9 7 3 3 1 9 9 13 2
7 15 13 0 2 1 12 2
19 0 2 16 15 15 13 13 2 10 9 13 10 9 2 16 1 13 4 2
11 0 2 16 3 13 13 9 1 15 15 2
4 15 13 0 2
13 3 13 3 0 13 0 15 15 13 13 1 15 2
2 3 2
17 16 13 12 9 2 7 15 9 9 1 15 13 0 2 7 0 2
9 16 0 2 15 13 1 9 0 2
15 3 15 13 9 15 15 9 0 13 2 16 9 13 13 2
14 16 7 13 0 2 13 16 1 15 13 1 12 9 2
12 7 3 13 16 1 15 13 12 9 1 9 2
17 7 3 15 9 13 1 15 1 12 9 2 7 1 15 7 15 2
12 16 1 12 2 3 3 13 12 7 12 3 2
10 12 3 3 13 12 9 16 0 13 2
18 16 7 13 15 7 15 9 1 15 2 3 15 13 10 9 10 9 2
11 7 15 13 1 9 13 2 16 13 4 2
11 3 15 15 12 13 15 15 13 9 9 2
8 3 3 0 13 13 12 9 2
2 0 2
27 15 15 15 13 15 13 16 13 15 13 2 0 13 15 13 2 16 9 15 9 3 13 15 1 15 0 2
14 7 15 15 13 13 10 9 13 13 16 13 15 13 2
8 3 0 13 16 15 15 13 2
12 7 3 0 13 16 13 0 15 15 13 13 2
9 7 1 13 0 13 13 0 9 2
3 9 0 2
30 16 3 15 15 13 13 3 13 15 13 16 13 13 2 13 16 9 10 9 3 13 0 1 15 2 7 1 15 13 2
12 15 7 1 16 13 9 13 13 1 10 15 2
6 15 13 9 15 13 2
16 3 15 13 13 13 1 15 3 1 15 16 13 9 1 9 2
9 15 13 1 9 15 15 13 13 2
16 13 3 16 15 15 13 13 13 13 1 15 16 13 15 13 2
2 3 2
19 9 13 15 9 9 7 4 1 15 13 1 15 9 2 7 1 15 15 2
9 16 1 15 13 16 13 3 9 2
11 16 1 15 2 3 0 13 16 15 13 2
13 15 3 15 13 9 9 2 3 13 13 0 0 2
7 0 3 13 13 0 9 2
2 0 2
16 16 13 0 9 2 13 16 9 9 3 13 12 9 1 15 2
13 13 3 13 15 13 9 0 1 15 7 1 15 2
22 7 15 13 0 2 16 9 0 3 13 9 7 9 0 7 13 2 16 1 13 4 2
16 7 3 9 0 13 9 15 9 2 16 13 13 1 9 9 2
7 0 13 3 13 0 9 2
2 3 2
8 9 0 15 9 13 3 12 2
12 7 15 9 13 9 10 2 16 1 13 4 2
8 0 13 3 13 16 12 9 2
2 3 2
26 1 15 9 9 13 9 15 13 9 2 3 15 10 9 1 13 13 2 16 1 15 1 3 9 13 2
8 7 0 9 13 0 13 9 2
7 13 3 1 15 0 9 2
7 15 3 9 1 0 13 2
2 0 2
29 1 15 9 13 9 1 15 9 13 2 7 3 1 15 9 13 12 0 2 15 13 9 10 15 1 15 9 13 2
16 15 3 13 1 15 12 9 2 13 16 1 15 12 9 13 2
6 7 10 1 9 13 2
11 13 3 13 12 3 15 13 9 10 9 2
4 15 9 13 2
2 3 2
19 1 15 9 15 15 13 9 13 2 3 1 9 13 0 9 2 7 9 2
21 0 3 9 12 13 9 2 7 1 15 0 9 13 15 15 13 9 2 9 13 2
14 3 7 9 2 15 13 10 9 2 13 12 0 13 2
12 15 7 9 0 9 3 1 0 9 13 13 2
5 3 8 12 13 2
11 13 2 9 2 9 9 10 9 12 13 2
4 7 8 12 2
8 3 13 15 9 15 1 15 2
4 7 8 12 2
8 12 9 2 12 9 2 8 2
9 15 7 9 13 0 9 9 13 2
37 16 0 15 12 9 0 13 13 2 1 15 10 15 15 9 13 13 4 13 2 10 9 0 9 9 13 2 7 0 9 9 7 9 7 9 9 2
23 15 3 9 13 3 1 0 9 13 2 16 0 9 2 7 3 9 7 9 2 9 13 2
4 16 15 9 2
9 3 13 0 15 1 9 2 9 2
9 7 3 2 15 13 2 9 13 2
9 7 0 3 1 0 9 9 13 2
20 3 3 15 9 13 0 9 2 12 0 13 9 2 15 15 15 9 3 13 2
31 15 3 9 9 10 9 13 2 16 13 9 7 9 3 12 2 7 0 9 13 2 1 3 9 0 9 9 9 13 13 2
5 16 9 13 0 2
37 1 7 0 9 13 2 16 9 13 2 3 13 9 9 13 9 9 2 1 13 4 0 12 9 13 2 15 7 1 15 9 7 9 7 9 13 2
16 1 3 9 0 0 13 3 13 2 1 13 4 15 0 13 2
12 13 3 13 16 1 0 9 9 0 15 13 2
23 15 3 0 9 3 1 12 13 2 3 3 1 9 2 7 3 1 0 9 9 7 9 2
16 13 3 15 3 7 0 0 1 9 15 1 15 10 9 13 2
10 13 3 9 9 1 9 9 7 13 2
7 15 7 9 12 15 13 2
12 3 1 15 15 15 15 9 13 2 0 13 2
15 1 3 9 15 1 9 10 13 2 13 9 9 10 9 2
12 7 3 13 9 0 0 13 1 9 10 9 2
20 3 7 9 13 16 1 15 15 3 9 0 13 2 15 13 13 0 16 0 2
11 13 13 3 1 15 9 9 9 0 13 2
15 3 7 3 16 0 0 13 2 16 1 9 0 7 0 2
8 3 3 9 13 4 9 13 2
12 3 1 9 15 15 4 13 13 2 0 13 2
9 7 1 15 1 15 0 9 13 2
22 7 1 9 0 0 3 13 2 16 15 13 9 10 9 7 9 2 7 13 0 9 2
7 7 3 9 0 13 13 2
15 10 3 15 1 10 9 13 13 2 1 9 15 9 13 2
21 9 7 3 13 1 15 9 2 7 15 9 10 9 9 13 2 16 1 13 4 2
4 13 3 0 2
2 0 2
25 10 9 15 13 9 13 1 15 1 15 13 2 16 15 13 1 15 2 13 1 15 1 9 13 2
8 9 3 1 15 13 15 13 2
25 13 2 16 9 13 1 15 13 2 9 9 1 15 3 13 2 16 13 15 1 9 9 13 13 2
41 9 7 13 9 15 9 1 15 13 2 16 7 13 9 1 9 2 16 13 4 2 7 9 10 13 15 9 7 9 2 1 15 13 10 9 2 16 1 13 4 2
6 13 3 15 13 0 2
2 3 2
38 1 9 13 15 15 13 9 3 2 16 9 0 2 15 15 13 9 3 2 16 9 2 16 1 13 4 2 15 15 13 9 7 9 2 16 9 10 2
22 7 9 2 1 13 1 9 2 3 13 9 13 2 16 7 1 15 2 3 7 0 2
25 1 3 9 0 13 0 1 10 9 2 13 16 9 2 15 13 9 0 2 13 0 1 10 9 2
2 3 2
12 3 9 15 9 13 2 3 0 13 9 13 2
24 3 10 9 15 13 9 2 13 9 10 9 2 15 7 3 13 15 9 2 13 1 9 9 2
14 9 7 13 9 0 1 10 9 2 16 1 13 4 2
4 13 3 0 2
2 0 2
7 15 9 0 13 0 13 2
10 3 1 0 7 0 9 13 0 13 2
22 16 3 15 9 13 13 2 13 16 13 9 15 1 15 15 15 13 0 9 15 9 2
16 7 9 0 3 13 13 15 9 2 16 15 13 0 1 15 2
10 3 9 10 13 0 2 7 15 0 2
2 3 2
15 10 15 13 15 9 2 3 13 9 3 15 9 0 13 2
32 7 3 13 13 15 9 2 7 3 13 2 15 0 13 15 9 16 1 15 15 1 10 9 13 9 7 15 9 13 10 9 2
5 15 7 9 13 2
11 15 3 9 13 13 15 0 7 9 9 2
6 13 3 0 1 9 2
2 0 2
8 9 10 1 0 1 13 13 2
16 15 9 13 16 2 15 9 13 13 2 9 10 0 13 13 2
15 3 7 13 15 9 9 1 0 16 13 15 9 0 0 2
14 13 3 13 15 9 0 0 2 15 13 13 0 9 2
5 7 15 13 9 2
5 9 3 13 0 2
2 3 2
8 9 3 13 13 1 10 9 2
16 9 7 10 3 13 13 16 1 9 2 15 13 0 10 9 2
10 3 3 13 15 13 9 10 0 9 2
15 16 3 10 13 13 15 0 13 2 13 9 13 3 13 2
2 0 2
25 9 0 3 13 13 1 9 13 2 16 15 13 1 10 9 2 15 7 13 9 15 7 9 9 2
6 9 7 9 9 13 2
8 7 9 3 13 9 0 13 2
20 13 3 1 9 0 2 15 3 13 13 16 1 9 0 2 16 1 13 4 2
7 13 3 9 9 13 0 2
9 15 7 9 13 1 13 9 9 2
13 15 3 13 2 3 3 13 9 1 9 0 9 2
29 3 15 13 3 13 0 1 13 3 9 3 13 1 9 1 9 13 2 16 0 9 9 13 1 13 9 16 9 2
19 7 15 15 3 3 13 2 0 13 1 9 2 7 13 15 9 1 9 2
18 3 2 16 9 13 4 16 3 0 3 13 2 13 9 9 13 0 2
19 15 7 9 2 3 1 15 15 13 9 9 2 13 1 13 9 0 9 2
37 13 3 9 13 9 0 9 2 16 15 0 13 2 13 15 9 9 0 0 9 9 13 16 9 1 0 13 9 9 16 1 0 4 13 1 9 2
15 15 7 9 13 2 1 9 13 3 13 9 9 13 0 2
33 3 7 1 9 2 1 15 2 7 1 0 2 1 15 2 13 2 15 13 13 1 9 15 15 3 13 2 1 13 0 13 9 2
11 7 3 2 15 13 9 7 9 2 13 2
11 13 7 9 9 0 13 1 9 9 0 2
18 3 2 3 9 0 0 13 7 13 2 3 0 9 0 1 9 13 2
34 13 3 2 1 9 13 13 15 9 13 9 9 2 16 9 9 2 15 15 9 13 2 3 13 13 2 7 0 2 7 3 9 0 2
2 0 2
12 15 9 3 13 0 3 15 9 9 13 0 2
16 15 3 15 9 13 0 2 13 16 13 9 1 9 9 0 2
6 7 9 9 13 0 2
8 13 4 3 1 15 13 0 2
17 1 3 3 13 2 15 9 10 9 1 15 2 13 15 13 0 2
9 15 7 9 0 9 9 9 13 2
4 13 3 9 2
13 0 9 7 0 3 2 7 9 15 3 13 9 2
22 15 3 9 13 0 9 9 2 15 10 0 13 0 9 9 2 3 1 15 9 13 2
61 0 3 9 13 2 13 2 9 0 9 1 9 9 13 2 1 9 2 15 13 0 0 9 9 2 7 1 9 2 15 13 0 9 0 9 9 2 7 1 9 9 0 2 1 15 15 13 15 9 2 7 13 15 0 9 2 13 0 10 9 2
42 7 1 13 4 1 13 9 9 16 3 13 15 9 0 2 7 15 13 16 13 13 0 9 15 9 0 2 13 16 7 13 9 7 9 1 9 0 15 13 0 9 2
5 16 9 13 13 2
10 1 13 7 13 13 16 9 13 13 2
32 13 3 4 1 16 1 13 7 13 3 13 0 1 0 13 2 7 13 0 10 13 2 16 0 13 2 1 12 0 13 15 2
10 13 7 15 15 13 1 9 7 9 2
16 0 3 3 13 15 13 2 16 1 15 13 13 7 3 13 2
15 9 3 13 1 0 13 15 13 7 16 13 13 7 13 2
26 1 9 7 15 13 1 9 7 9 2 13 7 13 13 13 13 2 0 7 7 13 13 13 3 13 2
34 1 3 15 15 13 10 0 13 2 15 9 13 2 13 13 3 3 13 2 13 16 13 1 9 15 13 9 13 15 16 0 1 13 2
7 3 7 16 0 0 9 2
22 3 9 0 3 13 9 0 2 7 15 13 9 2 1 7 9 9 3 13 16 0 2
22 15 7 15 13 0 7 0 0 2 13 0 15 15 13 0 7 0 16 3 7 3 2
9 13 3 0 13 13 0 16 13 2
11 7 3 13 13 15 13 15 2 13 13 2
24 0 3 3 7 15 0 0 13 13 2 16 13 15 13 13 9 1 15 16 15 16 0 13 2
17 13 3 9 13 13 13 9 16 0 13 13 15 2 16 9 13 2
2 3 2
21 15 0 13 13 16 13 9 0 3 1 15 0 13 15 2 7 1 13 3 0 2
8 3 0 13 13 0 9 9 2
30 13 3 2 1 10 13 13 1 15 9 15 13 1 13 2 16 9 1 15 13 0 13 2 13 0 9 7 0 9 2
11 9 7 1 9 0 3 13 16 1 9 2
12 13 3 0 13 2 15 9 13 2 13 13 2
2 0 2
22 1 15 9 13 13 16 13 1 9 13 9 15 15 13 1 9 2 7 3 1 0 2
23 10 7 13 15 13 1 9 2 13 1 0 13 2 15 9 13 2 16 9 1 9 0 2
19 1 3 1 9 13 0 13 1 9 2 0 13 16 0 13 13 1 9 2
7 0 13 3 9 13 13 2
2 3 2
11 1 15 15 9 13 13 16 13 1 9 2
14 15 9 13 16 9 13 13 1 9 1 9 1 9 2
15 3 7 9 13 0 7 3 0 2 16 9 13 9 9 2
12 9 7 13 1 9 13 12 1 9 9 13 2
27 3 2 16 1 15 4 9 13 1 9 16 13 1 9 2 13 9 15 1 15 13 13 16 13 1 9 2
9 13 4 7 1 9 13 3 0 2
4 13 3 13 2
2 3 2
31 9 15 9 13 15 1 15 9 9 13 2 16 1 13 4 2 7 1 15 15 9 1 15 13 2 16 3 1 0 13 2
11 1 9 7 9 0 13 16 15 13 0 2
14 3 1 15 15 13 3 10 2 13 1 15 10 9 2
5 9 3 13 13 2
2 3 2
21 10 15 13 13 1 15 9 2 7 15 13 15 9 2 7 13 15 9 1 15 2
11 15 3 3 1 15 16 1 15 9 13 2
7 0 7 13 1 9 13 2
8 3 3 1 9 0 9 13 2
12 3 3 3 13 3 7 1 0 2 7 0 2
5 15 3 13 9 2
27 1 3 15 3 13 15 9 2 16 9 9 3 13 2 13 16 15 13 9 1 15 2 15 13 9 9 2
24 15 7 13 15 13 10 9 2 7 13 1 15 13 2 15 9 13 2 16 1 1 13 13 2
9 3 7 13 9 9 13 16 13 2
5 9 3 13 13 2
2 0 2
10 10 15 13 0 2 13 1 15 9 2
11 3 9 0 13 0 0 2 16 9 9 2
19 7 9 1 9 0 13 13 0 2 16 0 2 7 3 1 9 10 9 2
12 13 3 16 13 1 15 9 9 7 3 13 2
21 15 7 9 13 3 13 16 13 2 1 3 13 15 9 1 10 9 16 1 9 2
19 7 1 13 13 15 13 13 2 16 13 0 2 3 3 0 13 13 13 2
19 9 3 2 15 13 9 0 0 2 1 15 10 15 13 2 13 13 13 2
8 15 7 9 3 9 0 13 2
7 13 3 9 12 1 9 2
7 0 9 13 7 0 9 2
3 7 12 2
7 1 15 13 9 7 9 2
3 1 9 2
8 0 13 4 9 10 1 15 2
4 7 8 12 2
8 3 9 9 9 7 9 9 2
16 15 7 9 9 1 3 1 9 13 16 1 13 9 9 13 2
19 3 9 2 15 1 9 9 13 2 13 1 8 2 15 13 13 7 13 2
7 16 13 9 13 10 9 2
16 1 15 7 16 9 13 13 2 13 16 10 13 13 10 9 2
21 13 3 13 9 13 1 15 13 2 3 1 15 0 13 2 16 9 13 1 13 2
14 3 3 15 13 0 1 15 16 13 2 7 13 13 2
10 15 7 13 1 9 2 13 0 9 2
15 13 3 9 13 0 9 2 7 0 9 2 7 15 9 2
9 3 9 13 10 9 7 10 9 2
2 3 2
9 13 13 1 9 16 9 1 9 2
12 7 9 0 13 15 9 2 16 1 13 4 2
7 3 7 13 0 15 9 2
12 9 7 0 13 9 9 2 15 13 9 9 2
9 13 3 16 13 0 13 15 9 2
2 0 2
13 9 0 13 9 16 9 0 2 16 9 16 9 2
34 9 7 7 9 9 13 15 15 9 2 16 13 13 2 16 13 4 2 1 15 9 13 15 0 2 7 1 9 2 16 1 0 13 2
17 16 3 10 9 3 13 10 9 2 15 13 10 9 0 7 9 2
10 7 3 3 13 1 9 9 7 9 2
5 3 3 13 0 2
2 3 2
5 13 13 9 13 2
19 16 3 9 13 3 13 10 13 2 13 16 13 1 15 16 9 1 9 2
9 7 3 1 9 13 9 7 9 2
9 15 13 0 2 16 1 13 4 2
2 3 2
7 10 9 13 1 10 9 2
18 16 3 9 9 13 15 16 0 9 2 13 9 15 15 15 1 15 2
15 7 3 9 3 13 10 9 2 1 9 15 13 9 15 2
34 16 7 0 13 13 15 9 2 0 13 16 13 15 13 0 2 0 7 0 2 7 9 3 13 2 7 10 15 1 0 9 13 4 2
24 3 13 3 9 1 9 13 2 7 1 0 15 13 13 2 7 15 9 7 9 1 13 13 2
11 16 9 1 15 15 13 16 1 10 9 2
22 1 15 7 15 1 13 4 2 0 13 16 9 0 15 15 9 0 13 16 10 9 2
18 9 3 0 9 0 13 0 9 2 16 9 15 9 9 13 0 9 2
12 0 7 9 0 13 15 9 2 16 13 4 2
20 13 3 15 15 0 9 9 7 9 16 15 0 9 16 10 9 9 0 13 2
5 15 1 13 13 2
2 3 2
16 1 9 0 13 9 13 9 2 16 1 9 0 9 9 13 2
11 13 3 9 0 1 9 16 9 1 9 2
18 16 3 9 0 15 15 9 0 13 16 15 2 13 1 9 9 15 2
10 15 13 3 13 2 16 1 13 4 2
2 0 2
12 9 0 1 9 1 9 15 13 9 0 13 2
8 9 15 9 10 1 9 13 2
14 1 9 7 3 13 15 13 9 2 16 1 13 4 2
13 3 3 13 1 9 15 15 9 1 15 0 9 2
2 3 2
7 9 0 9 13 15 13 2
18 16 3 1 9 0 13 15 0 9 1 9 15 2 9 15 13 13 2
9 7 3 0 9 2 7 15 9 2
25 15 3 0 9 3 13 13 2 16 3 0 9 3 13 0 1 15 2 7 15 9 13 15 0 2
18 7 3 13 13 1 9 0 9 15 1 9 15 15 13 15 9 9 2
8 15 3 9 13 15 1 15 2
35 3 7 1 15 2 16 3 15 13 9 7 0 2 13 7 15 9 15 3 10 7 15 9 13 0 2 7 3 3 10 9 15 0 13 2
4 7 1 15 2
7 13 3 15 9 0 15 2
14 3 0 13 16 1 15 13 15 9 0 1 15 9 2
2 3 2
10 13 9 13 15 9 2 16 13 4 2
20 16 3 13 1 15 9 15 3 13 10 9 2 13 1 15 15 1 10 9 2
4 15 13 0 2
12 3 3 13 1 15 9 15 3 13 10 9 2
6 16 9 13 9 15 2
11 1 15 7 0 13 16 15 15 9 13 2
18 1 3 1 9 0 9 1 9 13 13 2 1 12 9 0 9 13 2
10 12 13 16 9 0 9 9 13 13 2
7 15 13 16 9 9 13 2
13 15 3 3 13 0 3 9 1 13 0 9 13 2
25 15 7 0 9 15 13 9 0 15 9 0 13 2 13 15 9 3 15 2 13 7 9 15 3 2
6 15 3 9 9 13 2
2 3 2
14 9 0 0 13 1 15 16 1 9 7 0 9 13 2
21 15 3 13 1 10 9 1 10 9 7 0 9 13 2 15 13 0 1 10 9 2
12 7 10 0 13 1 16 13 12 9 1 13 2
10 15 7 9 13 13 2 16 13 4 2
18 3 2 1 13 0 3 2 7 15 15 0 13 12 2 0 15 13 2
2 3 2
16 1 15 15 9 13 16 9 1 9 7 13 1 9 12 13 2
9 0 7 9 13 3 9 1 9 2
10 15 3 13 1 9 7 0 1 9 2
14 9 7 9 1 15 9 0 13 2 16 1 13 13 2
21 1 3 9 0 7 9 0 13 12 2 1 13 2 0 13 16 9 9 15 13 2
10 9 3 13 7 10 9 7 10 9 2
2 3 2
13 10 15 13 1 15 1 9 0 2 13 1 15 2
10 9 7 0 13 1 9 1 9 0 2
19 3 9 0 9 7 9 0 12 7 15 13 2 1 9 10 13 10 13 2
6 9 3 13 9 10 2
9 3 15 2 1 15 13 10 9 2
2 0 2
13 9 9 2 16 7 15 9 9 2 1 9 13 2
11 3 3 13 9 9 9 3 13 9 0 2
15 7 9 0 13 9 0 2 1 13 9 9 7 0 9 2
18 9 7 9 0 13 3 0 2 1 13 15 9 0 2 16 13 4 2
5 9 3 15 13 2
2 3 2
8 9 10 9 1 9 0 13 2
24 1 15 7 9 1 9 13 13 0 13 13 9 2 1 9 0 15 13 2 15 9 13 13 2
6 0 7 0 9 13 2
6 9 3 0 15 13 2
6 15 7 9 0 13 2
16 13 3 9 2 12 8 12 2 16 9 9 13 3 0 9 2
10 16 9 0 7 1 15 0 15 13 2
14 1 13 7 13 16 9 0 7 1 15 0 15 13 2
16 15 3 0 9 4 0 7 1 15 1 9 13 15 9 13 2
9 9 3 9 15 13 9 9 13 2
16 7 15 15 9 13 15 13 15 16 10 9 2 16 13 4 2
14 3 13 1 15 0 7 1 15 15 13 15 16 15 2
2 3 2
10 0 13 3 0 0 7 1 15 13 2
9 12 3 9 3 13 3 0 13 2
10 9 7 15 3 13 2 16 13 4 2
24 16 3 13 15 15 3 0 7 1 15 13 2 13 16 9 15 13 1 9 15 1 9 15 2
6 15 7 13 15 0 2
8 3 3 9 0 13 1 0 2
4 15 13 0 2
2 0 2
6 9 9 13 1 9 2
18 16 3 9 13 15 7 15 1 15 3 0 9 2 13 0 9 0 2
20 3 7 10 9 13 1 0 13 2 7 15 9 0 13 15 3 13 10 9 2
7 15 15 0 13 13 4 2
18 13 3 15 1 9 4 13 3 0 7 1 15 13 2 16 10 9 2
2 3 2
16 9 2 1 16 13 13 1 10 13 2 13 1 9 9 15 2
23 16 3 15 15 4 13 1 9 0 7 1 15 2 13 16 15 13 1 9 9 15 15 2
9 15 13 0 2 16 1 13 13 2
2 3 2
5 13 13 9 13 2
10 1 3 15 9 9 13 16 9 13 2
13 15 3 13 1 15 16 13 12 1 15 15 13 2
22 16 3 15 15 1 9 4 0 13 1 15 2 13 15 15 9 15 2 7 15 0 2
4 15 13 0 2
2 0 2
7 1 0 13 13 9 13 2
23 16 3 13 0 13 1 9 3 0 13 7 1 15 2 13 16 9 9 13 1 0 13 2
14 7 3 7 13 0 9 13 2 7 9 13 9 9 2
9 15 15 0 13 1 13 0 13 2
21 13 3 16 15 15 4 0 7 1 15 13 1 9 2 15 13 15 16 10 9 2
2 3 2
22 9 0 9 7 9 13 1 15 15 4 1 15 7 0 13 2 1 15 13 15 9 2
29 16 3 9 15 1 15 13 3 1 15 7 0 13 2 15 9 0 9 7 9 13 1 15 15 13 15 1 15 2
16 15 7 13 0 2 1 10 9 13 15 9 2 16 13 4 2
17 3 3 0 13 16 13 1 9 0 7 1 15 13 15 1 15 2
7 16 9 13 15 1 15 2
21 1 15 7 16 15 13 0 7 1 15 2 16 15 1 15 1 15 13 13 13 2
10 9 3 9 0 13 1 9 10 9 2
9 3 7 13 13 15 1 9 13 2
11 15 7 9 13 1 10 9 9 13 15 2
14 1 3 10 9 0 13 2 13 13 16 3 15 13 2
2 3 2
16 10 9 1 10 9 0 13 9 2 1 10 9 13 15 0 2
17 10 7 15 13 1 15 2 13 1 15 1 9 15 1 15 13 2
24 16 3 9 15 9 13 9 2 1 15 13 1 10 9 0 2 9 13 10 1 15 13 0 2
13 15 7 13 1 15 1 9 0 2 1 15 13 2
10 9 3 9 15 1 15 1 15 13 2
2 0 2
23 15 13 9 9 15 2 13 10 15 1 9 15 0 13 13 7 15 15 13 1 10 9 2
11 9 7 1 10 9 13 16 13 15 9 2
11 1 3 9 15 13 2 13 15 13 9 2
9 15 13 3 13 16 13 0 13 2
6 15 13 15 1 15 2
7 15 3 15 15 9 13 2
7 3 9 13 15 1 15 2
25 13 3 15 12 9 2 13 9 13 15 3 0 7 1 15 13 2 15 0 16 1 9 10 13 2
16 15 3 9 13 9 13 2 1 12 8 1 8 8 2 13 2
15 3 1 9 0 15 13 2 7 1 12 9 9 13 10 2
3 7 1 2
7 0 9 15 13 13 15 2
9 15 3 9 13 13 9 0 9 2
7 3 1 9 1 9 13 2
13 13 1 13 0 10 2 3 1 15 13 15 13 2
9 16 9 13 0 9 1 10 9 2
50 16 0 15 13 16 9 1 15 9 3 13 9 16 0 2 3 13 15 16 13 9 2 1 15 16 9 13 13 1 9 15 15 2 13 13 16 9 13 10 15 9 16 1 3 13 13 7 1 9 2
9 15 13 13 9 1 0 9 15 2
12 1 15 7 9 2 9 13 9 10 9 13 2
13 15 7 1 1 13 15 13 2 7 1 0 13 2
19 3 3 15 1 15 9 13 13 15 3 4 1 15 13 7 13 7 0 2
8 13 7 9 2 13 15 9 2
21 15 3 13 1 15 9 13 13 13 9 7 10 9 0 15 13 1 9 7 9 2
16 7 9 15 13 7 10 9 0 15 13 1 15 7 9 15 2
10 16 3 15 9 13 2 3 13 4 2
11 15 7 13 2 13 16 1 15 0 13 2
22 15 13 2 13 3 16 1 15 0 13 2 7 3 1 10 9 0 1 1 0 9 2
8 3 9 13 15 13 1 9 2
23 15 7 13 13 0 7 0 9 1 9 2 13 3 10 15 1 9 13 2 0 7 0 2
15 9 3 0 1 9 9 13 2 1 16 13 1 3 13 2
2 3 2
24 10 15 13 1 9 2 13 9 1 9 15 13 1 0 13 9 2 16 9 13 13 9 13 2
22 9 7 9 13 9 1 9 2 1 10 9 13 10 13 2 15 7 13 16 13 9 2
13 13 3 13 10 0 2 1 16 13 13 1 15 2
2 0 2
8 9 9 3 13 13 1 9 2
5 13 3 9 0 2
11 13 3 1 15 9 9 9 1 9 13 2
34 3 7 1 9 15 9 1 9 9 13 2 16 9 13 1 12 2 7 3 15 9 1 9 9 13 9 13 13 1 0 16 13 13 2
13 13 3 16 9 1 9 13 1 9 15 9 13 2
9 13 7 9 0 13 9 9 13 2
8 3 7 9 9 9 9 13 2
23 0 7 9 9 3 13 13 1 9 15 9 0 2 16 10 3 9 13 1 9 13 13 2
19 13 3 15 0 9 2 15 1 15 1 10 15 13 2 13 9 10 9 2
7 9 3 13 9 16 13 2
2 3 2
7 15 9 13 2 9 13 2
16 13 3 1 15 10 9 16 1 0 9 2 16 1 13 4 2
11 15 7 13 1 0 3 2 3 9 13 2
19 13 3 15 15 13 0 15 9 2 3 0 9 2 15 13 0 9 15 2
12 3 15 9 3 13 9 1 9 16 1 9 2
20 16 3 9 13 9 10 13 10 1 0 2 13 16 3 0 13 9 1 9 2
2 3 2
12 15 13 9 15 2 13 1 15 9 15 9 2
21 1 15 7 9 9 2 16 13 9 2 13 12 7 0 2 16 13 1 12 8 2
18 9 3 2 16 13 9 10 13 1 0 9 9 2 13 16 13 9 2
8 9 7 1 9 13 3 13 2
9 13 3 9 16 13 1 3 13 2
2 0 2
27 15 13 9 15 9 0 2 13 9 15 9 15 13 13 2 16 15 13 9 2 13 16 13 3 7 0 2
10 7 1 0 9 13 13 0 9 9 2
34 16 3 9 13 15 13 9 0 9 2 3 7 0 2 16 1 15 10 9 0 13 2 16 1 13 4 2 13 16 13 10 9 9 2
11 7 3 1 9 15 1 15 13 0 9 2
2 3 2
12 15 13 9 15 2 13 10 15 13 1 15 2
6 7 9 13 15 9 2
11 3 13 10 15 13 1 15 1 9 0 2
19 7 10 1 0 9 13 1 15 1 9 0 2 1 15 13 10 9 9 2
9 15 3 13 9 0 1 10 9 2
2 3 2
12 15 13 9 15 2 13 16 15 9 13 0 2
13 3 3 9 9 13 9 15 13 15 0 0 13 2
8 0 7 9 0 13 1 9 2
12 13 3 9 15 9 15 9 15 0 13 13 2
13 7 1 15 13 9 9 16 0 9 9 9 13 2
8 3 9 9 0 0 15 13 2
10 9 3 1 9 13 9 1 0 9 2
2 3 2
18 1 9 7 15 13 13 9 1 9 16 1 10 9 13 1 3 13 2
29 16 3 9 9 1 10 9 3 13 2 13 15 0 13 2 16 7 15 15 13 9 3 13 9 2 15 10 13 2
15 15 1 9 13 9 2 1 12 1 9 7 1 12 0 2
7 15 3 9 9 0 13 2
5 13 3 8 12 2
11 13 9 10 15 13 2 7 13 3 0 2
4 7 8 12 2
9 3 13 15 9 0 1 9 15 2
8 10 0 7 13 13 9 15 2
11 9 1 13 15 9 13 13 1 9 0 2
19 7 16 9 13 1 9 0 9 13 2 13 13 9 15 15 13 13 0 2
16 3 7 15 9 3 13 13 16 0 13 13 9 13 1 9 2
25 15 3 13 7 13 15 16 9 0 2 7 3 1 9 9 13 15 9 2 15 1 0 4 13 2
20 7 13 13 9 0 2 7 3 13 1 9 15 9 2 15 1 0 13 13 2
11 7 3 13 13 3 9 0 1 15 13 2
13 15 9 2 13 9 13 2 13 13 2 13 9 2
16 3 9 9 0 1 9 13 3 13 2 1 7 1 9 13 2
14 15 3 16 13 2 7 15 13 1 13 9 13 9 2
49 3 1 9 13 13 1 9 9 2 16 1 15 9 9 9 13 3 13 2 15 1 9 10 9 13 2 13 16 10 9 1 13 1 15 13 2 7 1 13 1 13 2 1 10 9 13 10 13 2
6 15 0 1 13 4 2
2 3 2
31 1 10 15 13 1 9 10 4 13 1 15 2 16 1 13 2 0 13 2 16 9 13 1 9 13 2 1 15 13 4 2
12 15 7 13 9 9 1 9 2 16 1 13 2
15 3 9 13 3 0 13 9 9 1 15 16 3 0 13 2
16 3 3 1 15 9 13 9 16 0 0 1 15 13 1 15 2
2 3 2
18 0 1 9 13 9 1 9 2 16 7 0 1 9 13 9 1 9 2
19 1 0 16 0 1 9 13 2 13 15 1 9 2 16 7 1 9 13 2
28 3 7 9 13 13 9 2 7 0 13 9 2 16 1 9 13 0 9 2 16 3 1 9 7 0 12 13 2
22 16 3 0 9 13 1 9 15 2 13 16 9 10 13 1 9 2 7 0 0 15 2
8 7 3 13 15 13 1 9 2
4 15 13 0 2
6 3 15 13 15 0 2
2 3 2
6 13 13 13 1 13 2
29 3 3 13 13 9 9 1 15 13 1 9 0 1 15 16 9 9 9 13 2 7 13 16 13 1 15 9 0 2
28 1 15 3 9 13 16 3 13 13 16 9 0 13 13 1 15 15 9 1 0 2 7 9 7 9 7 9 2
17 3 3 9 0 2 3 1 15 10 9 2 13 1 15 0 9 2
5 15 3 13 0 2
16 16 3 9 1 15 13 1 9 13 2 3 7 15 9 13 2
20 3 7 1 9 13 0 1 15 0 13 13 13 0 2 1 15 9 13 9 2
16 13 3 9 0 13 1 9 2 1 10 0 3 13 15 13 2
12 16 3 15 13 0 9 2 3 7 0 9 2
39 3 3 13 13 16 1 15 16 15 9 1 13 13 2 15 9 0 13 2 7 15 9 1 15 9 13 2 16 15 13 1 9 10 2 3 1 9 15 2
21 1 15 3 16 0 0 13 1 15 0 9 2 3 13 13 16 9 0 9 13 2
4 9 13 9 2
17 13 7 9 0 13 13 2 16 13 13 15 9 13 1 9 13 2
50 7 16 1 9 10 1 0 9 9 2 16 13 0 2 13 2 13 13 16 9 0 13 1 15 1 9 10 3 13 1 0 9 2 7 13 16 9 15 13 1 9 10 2 1 15 13 9 1 9 2
16 13 7 1 9 1 3 9 16 1 0 9 2 13 9 15 2
23 3 7 3 16 15 13 13 9 13 1 13 2 16 9 13 1 13 2 7 13 1 13 2
26 7 13 9 1 9 15 13 2 1 15 16 9 13 2 15 13 9 0 9 16 9 2 13 9 15 2
30 0 7 13 13 16 9 2 1 9 9 13 2 13 13 1 15 15 9 9 13 2 15 13 9 15 2 15 13 9 2
6 7 15 3 0 13 2
17 15 16 9 13 0 9 13 7 13 2 1 15 1 9 9 13 2
36 7 9 15 0 13 2 16 3 13 9 16 13 1 9 0 2 1 15 1 9 9 3 13 2 7 15 3 13 13 16 9 15 9 13 13 2
38 15 7 9 13 2 1 13 3 9 0 9 2 13 15 1 9 0 15 13 9 1 9 2 15 13 13 16 0 9 9 2 16 15 13 9 13 9 2
36 1 15 3 16 9 0 15 13 9 9 7 13 9 2 13 9 9 0 2 13 16 9 9 13 15 9 0 2 16 15 13 15 2 15 13 2
23 7 1 15 16 9 13 13 0 15 9 2 13 16 9 2 13 3 9 2 9 15 13 2
16 9 7 0 15 15 9 13 16 9 10 2 16 1 13 4 2
9 7 3 9 10 13 9 10 9 2
35 1 15 3 13 16 9 9 0 2 16 15 13 2 15 13 9 15 2 3 0 13 9 15 9 13 2 7 3 10 15 13 0 9 9 2
29 3 3 1 12 9 0 2 15 13 0 9 2 7 1 12 9 13 2 15 13 9 0 2 0 13 1 9 13 2
12 15 0 9 12 7 0 13 0 9 10 0 2
25 7 3 0 7 0 15 13 13 16 12 7 15 0 2 16 0 9 2 13 0 9 7 9 0 2
26 3 2 1 0 9 13 9 9 0 9 2 16 15 1 0 9 0 13 2 15 0 13 16 0 13 2
23 1 0 16 0 15 0 13 2 15 13 15 9 12 13 2 16 9 7 9 16 13 9 2
15 1 15 13 16 9 1 9 0 9 3 13 2 7 0 2
21 3 1 9 15 9 13 13 1 13 2 13 9 9 2 16 7 9 1 9 9 2
11 9 3 13 1 13 13 16 9 15 13 2
18 13 3 2 16 9 1 0 0 9 13 2 16 15 13 0 9 0 2
6 15 15 13 13 4 2
22 16 3 9 13 2 1 12 8 2 9 7 9 9 2 15 15 13 2 13 0 9 2
21 3 1 9 2 12 9 13 7 13 2 9 9 13 2 16 13 1 0 7 0 2
7 0 7 13 7 1 9 2
9 3 12 9 13 7 13 13 9 2
13 9 3 0 1 0 2 7 0 13 2 9 13 2
17 1 15 7 15 1 15 0 13 2 3 3 15 13 9 16 9 2
16 3 15 15 1 9 15 9 13 15 9 9 13 13 3 13 2
11 3 3 13 9 9 16 1 9 9 13 2
23 9 0 15 15 13 1 9 13 2 3 13 13 13 2 16 12 15 1 15 9 3 13 2
20 7 1 15 1 0 13 13 0 3 2 7 1 9 0 15 15 13 0 3 2
19 3 9 15 15 0 13 13 13 16 0 9 0 2 13 15 15 1 15 2
23 13 3 13 9 16 0 9 0 2 12 9 13 2 7 0 16 0 9 0 9 1 13 2
24 0 3 1 9 13 13 0 0 9 0 16 3 2 7 9 9 15 2 16 15 9 13 0 2
19 1 15 15 9 2 0 9 2 13 16 0 1 9 2 13 0 0 0 2
26 0 7 9 1 15 9 10 9 13 2 3 3 1 9 9 2 7 1 9 9 2 16 1 13 4 2
19 9 7 10 2 3 0 7 0 2 1 15 16 15 13 2 13 9 15 2
12 3 7 9 13 16 1 16 13 1 0 9 2
30 9 3 0 15 15 13 0 15 1 9 10 13 13 2 13 1 15 15 9 13 2 7 1 15 1 15 9 13 15 2
19 3 2 13 9 10 16 0 1 9 9 7 3 9 2 13 0 9 9 2
20 16 0 16 0 1 9 9 7 3 9 2 0 9 0 2 7 3 1 15 2
19 3 3 13 16 9 0 2 16 13 0 9 2 13 13 16 0 9 0 2
11 3 1 15 9 0 9 1 10 13 13 2
42 16 0 0 9 12 13 1 0 9 15 2 9 7 13 9 9 2 13 1 9 0 9 15 7 9 9 13 13 2 1 16 15 15 13 1 9 0 13 0 9 0 2
45 3 2 1 15 13 1 16 9 13 0 9 9 15 13 15 9 1 15 2 13 16 9 9 1 9 0 3 13 0 7 13 16 1 16 9 13 9 0 7 0 9 13 0 15 2
25 7 1 15 9 13 16 9 15 9 13 9 7 15 9 2 7 9 9 0 1 9 0 13 13 2
20 1 15 3 0 13 9 9 13 9 2 1 15 13 10 15 1 9 0 13 2
6 16 9 10 3 13 2
11 1 15 7 0 13 16 9 10 3 13 2
41 9 3 10 3 0 9 13 3 13 2 16 2 1 9 1 9 13 13 1 9 2 16 0 3 9 13 2 13 16 9 3 13 0 1 12 9 2 15 13 0 2
25 13 7 1 12 9 2 16 15 13 15 9 13 0 9 0 9 2 16 15 9 13 13 7 13 2
21 9 7 0 2 15 9 13 1 15 16 4 15 13 1 9 2 10 13 12 9 2
21 13 3 12 9 13 1 9 0 2 16 9 15 13 9 1 12 13 3 13 9 2
12 3 7 0 13 1 9 9 15 13 1 9 2
16 7 3 13 16 2 16 15 0 13 15 9 13 2 3 13 2
33 3 3 13 15 0 2 3 9 1 9 2 7 0 3 13 9 2 3 0 9 7 3 9 2 16 1 12 15 9 10 9 13 2
16 1 15 3 13 13 16 15 0 12 9 13 2 3 13 13 2
15 10 7 15 9 13 2 12 9 13 2 15 13 10 9 2
6 10 3 3 13 13 2
2 3 2
10 9 0 3 13 15 9 16 13 9 2
18 3 7 9 1 9 13 3 3 9 13 2 16 9 3 13 1 15 2
12 9 3 15 9 1 9 13 1 13 1 9 2
13 0 3 1 15 3 9 3 13 2 3 3 13 2
13 15 7 13 1 12 9 13 2 13 3 4 13 2
15 15 3 9 12 13 2 9 1 15 13 7 3 13 15 2
14 10 7 15 13 1 0 9 1 12 9 0 13 13 2
8 13 3 9 10 9 9 13 2
14 15 13 13 15 1 15 9 10 2 1 15 10 13 2
11 9 3 2 13 9 10 2 3 10 13 2
2 0 2
32 9 0 0 13 0 13 13 12 3 9 2 1 3 9 1 9 13 2 13 0 13 9 9 15 13 0 2 7 15 13 0 2
17 9 7 0 13 12 9 2 15 13 10 9 2 16 13 4 1 2
11 3 3 0 2 7 3 10 10 13 13 2
2 3 2
22 9 1 9 13 3 13 2 7 9 1 9 2 1 9 13 9 9 1 0 7 0 2
16 1 9 7 0 13 13 9 15 2 16 1 1 13 13 13 2
8 15 3 13 1 9 0 9 2
8 7 3 10 15 13 3 13 2
2 3 2
13 13 9 13 15 10 9 2 16 1 1 13 13 2
20 1 9 7 0 3 13 0 7 0 2 7 13 15 3 2 16 1 13 4 2
14 3 7 9 9 13 0 7 0 2 7 10 3 13 2
2 3 2
26 10 9 13 12 1 15 13 3 9 13 7 3 9 2 16 3 13 0 1 9 2 13 0 1 9 2
12 9 7 0 3 13 1 9 7 3 9 13 2
11 3 3 13 9 0 2 7 10 3 13 2
8 15 7 9 9 0 9 13 2
15 13 3 8 12 2 16 1 9 3 13 9 7 9 9 2
7 16 9 9 3 13 0 2
12 1 15 7 13 16 1 9 3 13 0 9 2
22 1 15 3 13 0 9 2 3 10 3 13 2 7 16 15 13 9 2 15 13 9 2
11 9 7 10 3 9 13 2 16 13 4 2
8 3 13 3 1 15 0 9 2
2 3 2
16 13 9 7 3 13 13 3 1 9 2 15 3 16 1 13 2
12 13 4 7 16 9 0 15 9 13 1 9 2
9 15 3 9 13 1 15 0 9 2
2 3 2
19 10 9 0 15 13 13 15 15 9 16 10 9 0 2 15 13 15 9 2
16 9 3 0 13 13 10 9 2 3 7 15 9 13 15 13 2
14 1 9 7 10 9 13 10 9 2 16 1 13 4 2
9 3 13 3 1 15 9 0 9 2
2 3 2
11 9 0 3 13 3 13 1 10 0 9 2
16 3 7 9 2 15 13 0 2 13 1 9 2 7 1 9 2
19 16 3 9 13 0 13 1 10 9 2 1 10 9 13 3 13 0 9 2
6 15 0 13 4 1 2
2 0 2
19 13 4 16 15 13 13 1 9 10 2 3 7 1 15 9 0 9 13 2
10 10 7 9 1 9 1 15 9 13 2
38 3 9 7 13 9 15 9 1 13 9 0 15 9 13 13 2 7 13 13 9 15 9 13 1 9 3 1 0 9 2 7 0 9 1 9 7 9 2
8 3 13 3 1 15 0 9 2
2 3 2
5 9 15 9 13 2
16 9 7 3 13 7 9 7 15 9 13 2 16 1 13 4 2
7 3 3 9 13 0 9 2
31 16 0 9 15 15 13 9 3 13 7 13 7 13 13 9 13 2 15 13 15 9 2 16 0 9 1 9 13 2 13 2
10 6 2 3 13 7 13 15 13 9 2
8 15 3 13 15 8 12 13 2
8 9 9 0 13 0 1 9 2
8 3 9 3 13 1 9 13 2
7 16 9 9 3 13 0 2
14 1 15 7 0 13 16 0 9 3 13 0 7 0 2
21 3 3 0 13 10 9 16 1 12 13 1 15 13 2 16 13 1 9 1 9 2
20 3 3 1 15 15 13 7 13 16 13 15 9 1 13 13 2 3 15 13 2
21 15 3 13 3 13 2 7 9 13 2 16 7 9 0 13 1 15 16 0 13 2
17 13 4 7 16 9 3 13 12 1 15 3 0 2 16 3 10 2
16 3 3 15 9 13 0 7 0 2 16 10 9 7 9 13 2
2 3 2
9 10 13 15 9 13 9 7 9 2
22 3 3 13 2 13 9 2 1 9 13 2 16 1 15 15 16 9 13 9 3 13 2
17 9 7 13 10 9 12 2 15 13 10 9 2 16 1 13 4 2
7 3 13 3 10 9 0 2
2 3 2
12 10 0 9 13 15 1 9 7 15 1 9 2
8 3 9 1 9 13 1 9 2
14 1 0 7 9 9 9 3 13 2 16 1 13 4 2
7 3 13 3 15 9 0 2
2 0 2
9 1 10 9 0 13 15 13 13 2
8 3 9 13 3 9 13 9 2
8 3 7 9 13 9 13 13 2
19 1 0 7 9 15 13 13 13 2 1 13 15 9 2 16 1 0 13 2
8 9 3 9 3 13 13 0 2
2 3 2
17 15 15 0 13 2 1 9 15 13 13 2 16 13 1 0 9 2
14 7 1 9 3 13 13 9 16 0 2 3 16 0 2
12 10 3 9 13 10 9 2 16 1 13 4 2
7 9 3 9 3 13 0 2
2 3 2
16 10 9 0 13 13 1 0 13 15 13 13 3 7 3 13 2
16 15 3 1 15 13 0 9 9 2 13 3 13 13 3 13 2
11 15 7 13 9 0 2 16 1 13 4 2
10 13 3 9 0 3 13 13 3 13 2
12 9 7 13 15 9 9 13 1 12 1 15 2
7 3 13 3 0 9 0 2
2 3 2
13 15 13 0 1 15 13 9 15 15 1 9 13 2
10 3 9 3 13 0 16 1 15 0 2
18 0 7 1 10 9 13 2 3 9 2 7 9 2 15 13 9 9 2
11 9 3 9 3 13 0 2 7 0 3 2
2 0 2
19 1 9 10 9 13 13 2 15 16 15 13 0 9 2 16 1 13 4 2
9 7 1 9 0 9 13 0 9 2
32 3 15 1 15 13 0 13 13 15 15 1 15 13 2 7 1 15 15 1 15 13 13 9 13 13 1 15 1 15 13 13 2
10 1 9 7 0 13 15 13 1 15 2
20 15 7 0 13 1 15 13 13 2 7 1 15 13 9 13 13 1 0 0 2
10 3 0 13 16 0 15 9 13 9 2
7 0 3 9 3 13 0 2
2 3 2
11 1 9 9 13 15 15 9 13 1 13 2
13 3 3 9 13 1 9 13 15 9 1 9 13 2
12 0 7 9 13 10 9 2 16 1 13 4 2
10 3 3 13 1 15 13 1 9 9 2
12 13 3 9 15 15 9 1 0 9 13 13 2
10 7 1 15 16 1 9 10 15 13 2
28 15 3 13 4 3 13 0 2 1 15 9 15 13 1 15 3 16 9 1 9 2 7 16 9 1 9 13 2
14 7 1 15 16 9 9 15 13 16 9 13 3 13 2
13 13 3 13 9 16 13 2 7 3 16 13 13 2
13 15 7 9 2 9 13 2 3 0 9 9 13 2
5 13 3 8 12 2
8 10 0 7 13 13 9 15 2
19 15 3 13 13 3 13 1 15 15 0 7 13 2 7 9 13 7 13 2
8 16 9 3 13 13 7 13 2
17 1 15 3 13 13 16 9 0 3 13 1 9 9 13 7 13 2
7 13 3 10 13 9 10 2
9 9 7 10 3 13 13 7 13 2
6 13 3 15 16 13 2
7 1 15 7 15 13 9 2
10 3 3 13 1 9 9 13 7 13 2
2 3 2
13 15 15 9 13 7 13 13 4 3 1 15 13 2
26 9 3 7 9 9 3 13 16 1 15 15 16 1 15 13 15 13 2 13 15 15 13 7 3 13 2
23 16 3 9 13 1 9 9 13 7 13 2 13 16 3 12 9 10 13 2 7 3 15 2
6 15 0 1 4 13 2
2 0 2
9 1 9 3 13 13 0 7 0 2
17 9 7 7 9 0 13 9 15 15 15 13 2 15 13 15 9 2
12 1 9 3 0 9 9 7 9 13 3 13 2
2 3 2
8 0 9 9 13 15 15 13 2
32 3 1 15 3 13 9 16 1 9 2 1 9 7 7 9 13 2 16 7 9 15 13 0 3 13 0 2 1 15 7 13 2
17 1 9 7 0 3 13 15 1 9 2 7 0 15 1 15 13 2
15 1 0 3 9 3 13 9 7 9 7 0 0 9 9 2
2 0 2
21 9 1 9 13 7 13 13 9 1 15 9 13 2 3 1 9 15 13 1 9 2
19 16 3 9 0 1 9 13 1 9 9 13 7 13 2 13 9 15 13 2
10 15 13 0 2 16 1 1 13 13 2
2 3 2
9 9 13 7 13 0 9 0 13 2
8 9 3 9 9 9 3 13 2
15 3 9 15 9 13 9 13 9 2 3 13 0 13 9 2
9 9 7 7 9 9 15 9 13 2
20 16 3 9 9 13 13 7 13 2 13 16 10 13 3 13 12 3 7 0 2
10 7 3 3 10 9 3 13 12 3 2
13 1 10 9 0 13 10 9 2 16 1 13 4 2
11 3 7 1 15 13 15 13 16 0 13 2
17 3 9 10 2 1 13 12 7 0 2 0 13 10 0 7 9 2
15 7 3 1 15 9 10 9 7 9 3 9 7 9 13 2
7 15 7 0 9 9 13 2
11 13 3 9 12 3 3 9 10 9 10 2
6 7 3 1 9 13 2
14 9 13 9 9 2 15 13 1 9 7 9 9 13 2
10 9 3 13 2 12 8 1 8 8 2
20 3 0 9 2 15 13 2 13 10 2 7 0 0 7 0 0 7 0 0 2
8 16 1 9 3 13 9 0 2
40 1 15 7 13 16 2 16 0 9 9 3 15 13 1 9 9 13 7 13 2 3 3 13 1 15 9 2 15 2 1 9 2 0 1 9 7 9 9 13 2
41 1 3 9 9 13 9 9 7 9 2 1 16 9 13 13 15 13 7 3 13 15 3 13 2 1 15 1 9 9 13 15 9 13 2 3 1 9 15 15 13 2
46 3 3 1 9 9 13 16 15 13 9 13 2 1 9 3 13 0 2 13 0 0 2 7 15 15 9 13 13 7 13 2 13 13 9 13 2 16 3 3 13 1 9 16 9 13 2
28 9 7 10 0 9 2 1 15 3 13 9 7 9 2 13 3 0 9 9 2 7 3 9 2 16 13 4 2
13 7 3 15 15 9 0 13 13 13 9 7 9 2
11 3 3 13 9 1 9 0 9 10 9 2
2 0 2
33 1 15 0 7 13 7 13 2 15 3 0 2 3 13 1 15 2 3 13 9 13 7 9 0 2 1 9 7 9 1 9 13 2
17 0 7 2 3 13 1 15 2 3 13 15 9 7 9 1 9 2
27 3 1 15 7 0 7 0 13 13 2 7 3 13 2 1 15 13 9 0 1 9 1 9 9 7 9 2
26 9 3 0 2 13 15 15 13 2 13 9 9 1 15 9 1 9 2 16 13 15 16 15 9 9 2
65 3 2 16 15 0 2 7 3 9 2 3 13 1 15 0 7 0 2 3 9 13 15 15 13 13 3 1 15 3 13 0 2 16 13 1 12 1 9 2 16 1 9 13 13 0 2 16 7 9 13 15 9 2 7 9 9 1 3 2 7 15 9 1 13 2
50 3 9 13 2 1 16 13 16 15 7 15 9 9 2 1 16 1 9 13 2 7 0 0 2 16 9 9 3 13 3 2 16 16 13 9 0 2 7 0 1 15 9 2 16 9 9 13 16 0 2
23 13 3 2 1 0 2 16 9 0 0 0 13 2 3 13 0 2 13 10 9 16 10 2
2 3 2
30 0 9 9 3 13 2 16 1 10 9 0 13 15 9 1 15 9 1 15 9 9 7 9 13 2 16 1 13 4 2
40 9 7 10 2 13 0 2 3 13 1 0 10 9 2 16 3 13 1 9 9 9 7 9 2 16 7 1 0 0 13 1 9 9 13 2 7 9 9 15 2
23 9 3 1 10 0 9 15 9 9 13 15 9 10 13 1 15 9 2 7 13 7 0 2
17 7 9 13 9 10 1 15 9 9 2 16 3 1 1 9 13 2
10 3 7 1 15 0 9 9 13 9 2
2 3 2
26 1 9 10 9 9 13 2 3 10 9 1 15 13 2 16 1 13 4 2 9 9 15 13 3 13 2
15 7 0 13 9 9 2 16 13 1 9 2 1 12 9 2
6 3 9 1 9 13 2
8 7 15 13 15 13 1 9 2
5 13 7 9 0 2
5 16 9 13 9 2
10 1 13 7 13 16 15 9 13 9 2
15 9 3 15 9 13 9 2 7 0 9 2 16 13 4 2
7 13 7 9 13 10 9 2
35 15 3 13 2 1 13 0 9 2 16 13 4 2 3 13 15 9 9 13 2 7 13 1 15 9 2 16 7 1 0 9 1 13 4 2
9 13 3 16 0 9 13 15 9 2
2 3 2
9 9 13 15 9 9 2 1 9 2
11 9 7 13 10 9 2 16 1 13 4 2
6 3 13 3 10 9 2
2 3 2
16 1 9 15 0 13 13 2 1 13 10 9 2 15 15 13 2
11 7 9 13 1 9 2 16 1 13 4 2
11 16 3 3 13 0 2 13 16 13 0 2
6 9 3 13 10 9 2
2 0 2
28 16 0 0 3 13 1 9 7 1 9 2 1 9 2 9 3 3 0 13 2 1 16 0 9 0 9 13 2
45 3 9 13 2 1 10 0 2 16 9 9 13 9 9 15 9 15 13 4 15 2 16 15 9 13 4 1 15 13 0 9 2 7 3 0 15 9 15 13 1 9 0 2 13 2
6 7 9 13 10 9 2
17 3 2 7 1 9 9 13 7 1 9 9 2 9 13 10 9 2
12 15 7 13 9 9 1 15 13 2 8 12 2
8 15 13 9 2 9 7 9 2
6 16 9 13 0 9 2
21 15 7 13 2 0 13 16 1 9 13 0 9 2 15 15 9 7 9 13 13 2
11 9 3 9 3 13 2 16 7 9 9 2
12 9 7 3 0 13 0 2 7 13 15 9 2
8 3 1 15 9 13 3 13 2
2 0 2
16 9 3 13 1 13 15 15 13 2 16 7 9 1 0 0 2
19 10 7 9 0 9 15 13 1 9 9 13 15 15 13 2 16 13 4 2
13 0 13 3 1 0 9 9 7 9 7 9 13 2
2 3 2
20 9 1 0 9 3 13 2 7 1 9 3 2 1 15 1 9 0 13 13 2
14 9 7 0 3 13 0 7 0 2 16 1 13 4 2
10 3 3 13 13 1 15 9 7 9 2
2 3 2
19 3 15 9 0 13 9 2 3 15 0 9 13 0 2 0 1 15 13 2
19 3 15 15 9 13 1 9 2 9 0 7 9 13 16 1 0 9 13 2
11 7 9 0 9 13 1 9 9 1 13 2
17 3 10 0 13 1 15 16 0 0 7 1 15 7 3 1 9 2
8 1 15 7 9 0 3 13 2
10 1 15 3 0 0 13 0 9 13 2
2 0 2
9 9 0 13 15 9 9 1 13 2
14 1 7 9 0 3 13 9 0 13 2 7 3 0 2
15 0 3 13 13 0 9 9 2 9 7 13 9 0 13 2
15 7 0 9 9 13 1 10 9 16 9 0 1 9 9 2
6 13 3 1 9 9 2
11 13 3 16 1 9 0 3 13 13 9 2
2 3 2
8 9 9 0 1 9 3 13 2
9 3 13 16 0 13 9 9 0 2
20 1 15 3 0 13 15 9 13 2 16 9 3 15 13 2 7 3 1 0 2
10 9 7 0 1 10 9 13 9 9 2
22 3 13 16 9 15 13 9 9 2 16 9 13 9 9 15 1 3 9 13 16 13 2
14 15 3 13 9 9 0 1 9 15 9 1 9 0 2
18 9 7 13 1 9 9 0 7 9 3 13 1 9 2 7 1 9 2
21 16 3 3 13 0 9 9 0 1 9 2 9 13 1 9 2 3 1 9 0 2
19 7 3 1 9 13 9 2 16 15 15 13 1 9 2 15 13 1 9 2
19 15 3 9 13 1 9 0 7 9 2 7 15 9 1 9 0 13 13 2
2 3 2
12 16 0 13 9 9 2 3 0 13 9 15 2
10 0 3 13 0 13 7 13 0 13 2
12 9 7 1 9 13 3 13 2 16 13 4 2
8 3 13 3 1 15 13 9 2
7 15 13 15 13 8 12 2
5 13 7 9 0 2
4 7 8 12 2
9 3 13 9 16 9 2 16 13 2
5 7 12 8 12 2
11 9 9 13 7 9 1 15 3 13 15 2
9 16 0 9 13 0 7 0 9 2
17 1 15 7 15 13 4 0 13 16 0 9 13 0 7 0 9 2
22 16 3 13 9 9 1 9 2 3 7 1 9 2 16 13 1 9 2 1 12 8 2
11 7 15 3 16 0 7 9 15 3 13 2
15 13 3 0 1 13 9 15 13 7 3 9 15 3 13 2
8 7 0 9 13 0 7 9 2
9 3 7 10 9 13 0 7 0 2
2 3 2
10 15 1 9 15 13 2 9 15 13 2
10 7 9 9 13 0 2 16 13 4 2
9 10 3 9 13 0 7 0 9 2
2 3 2
12 9 1 10 9 1 15 13 16 13 9 13 2
12 9 7 9 13 9 2 16 13 1 12 0 2
21 1 3 1 9 0 13 3 15 9 7 15 13 2 10 9 13 0 7 0 9 2
2 0 2
13 15 15 13 9 1 15 9 2 13 9 15 9 2
6 3 10 9 13 0 2
8 7 0 9 13 9 10 9 2
23 9 3 10 9 13 1 9 15 13 1 9 2 1 15 3 9 10 0 13 16 13 9 2
24 9 7 9 13 1 9 0 2 15 13 9 9 2 16 1 13 2 16 9 9 1 9 9 2
9 3 3 0 13 9 16 13 9 2
34 1 3 9 13 0 9 7 0 0 2 13 16 9 9 15 15 9 13 2 16 15 13 0 10 9 2 16 9 13 2 1 12 0 2
11 0 3 9 13 0 2 0 7 9 9 2
7 9 13 13 9 9 0 2
12 13 7 15 15 9 0 9 0 9 13 13 2
8 1 15 3 13 12 9 13 2
7 0 13 1 15 9 9 2
26 1 3 9 9 13 9 13 2 3 13 1 15 9 0 0 13 13 2 16 10 9 1 15 9 13 2
21 3 7 1 15 15 0 9 0 13 15 0 9 13 2 16 9 7 9 7 3 2
12 9 7 10 2 16 0 13 2 0 3 13 2
15 0 3 0 9 0 0 13 0 2 15 0 1 9 13 2
11 7 3 15 9 13 16 9 0 13 13 2
8 0 13 16 0 3 3 13 2
15 7 3 3 13 1 9 2 7 3 13 7 3 3 13 2
21 0 13 3 13 2 16 1 15 15 3 13 3 13 13 9 2 15 0 0 13 2
11 15 7 15 3 13 2 0 13 3 13 2
18 0 3 13 3 13 2 16 0 9 9 13 3 0 2 16 13 4 2
16 0 2 1 15 16 3 10 0 1 9 13 2 7 15 13 2
12 3 1 15 0 9 13 3 13 16 16 13 2
9 0 3 9 13 15 13 3 13 2
15 9 7 10 15 13 1 13 2 1 0 13 2 13 13 2
9 13 3 13 13 15 15 9 13 2
11 16 3 3 13 13 13 2 3 0 13 2
17 3 7 1 13 0 3 13 13 1 15 9 2 7 0 9 15 2
16 13 7 13 10 9 9 13 0 7 0 2 16 1 13 4 2
19 0 13 3 16 9 15 1 0 13 13 2 1 15 9 2 16 13 4 2
11 1 15 3 13 13 16 0 13 3 13 2
11 0 13 1 15 16 15 0 9 13 9 2
14 9 7 2 16 13 2 3 13 16 1 10 9 13 2
11 3 3 0 13 13 16 1 15 13 13 2
18 9 7 9 1 15 13 1 9 13 16 1 13 2 1 15 9 13 2
18 0 3 13 16 9 1 3 0 15 9 1 9 13 2 9 0 13 2
6 0 13 1 0 9 2
9 0 3 2 16 3 2 13 0 2
21 3 10 15 13 1 13 9 3 13 2 1 9 15 15 13 16 15 9 9 13 2
6 3 10 9 0 13 2
10 0 7 13 0 2 1 0 1 9 2
8 0 3 13 16 9 0 13 2
7 0 13 1 15 9 0 2
19 1 3 9 9 1 9 0 3 13 2 9 3 0 1 9 9 13 13 2
6 0 7 9 0 13 2
13 3 3 15 9 13 16 9 15 0 1 0 13 2
10 0 13 1 9 15 1 15 0 13 2
41 1 3 13 13 15 9 1 13 2 9 7 1 9 13 3 13 2 16 1 13 4 2 13 13 16 9 9 7 9 3 3 13 2 7 0 9 15 13 1 9 2
9 9 3 3 16 1 9 13 13 2
19 7 1 15 13 16 3 13 9 1 0 9 2 1 15 9 7 9 13 2
6 9 13 1 0 9 2
29 1 15 7 9 9 2 16 3 0 9 9 13 2 13 13 9 13 1 0 13 2 16 15 15 13 9 0 13 2
11 0 2 3 2 13 16 0 9 0 13 2
11 0 2 16 13 15 15 3 13 1 9 2
9 0 2 16 13 13 0 0 9 2
7 0 2 16 13 9 9 2
6 0 2 16 13 0 2
11 0 2 16 13 15 0 7 0 1 9 2
11 0 2 16 13 9 7 9 15 7 9 2
5 16 9 0 13 2
11 0 3 13 16 0 9 9 3 13 13 2
13 13 3 4 1 16 9 13 15 16 13 9 15 2
7 9 7 9 13 9 0 2
14 15 3 9 9 13 9 2 16 13 15 13 1 9 2
20 0 7 3 13 9 0 2 7 13 9 0 1 0 2 16 13 1 12 0 2
17 9 3 13 9 15 1 15 3 0 1 0 2 7 3 1 0 2
2 3 2
26 13 9 1 15 13 9 9 2 0 13 9 15 13 2 16 2 13 9 0 7 9 15 2 13 9 2
36 0 7 9 13 1 9 13 7 9 13 2 16 9 9 1 15 9 7 15 9 2 16 9 9 0 1 9 7 9 2 16 13 1 12 0 2
20 3 2 16 15 13 1 9 9 0 2 3 15 13 1 9 9 16 13 13 2
26 15 3 13 9 9 2 7 15 1 15 9 13 2 7 9 1 9 13 2 15 3 13 13 9 0 2
13 7 9 9 1 1 9 7 9 13 7 9 13 2
20 1 3 10 13 13 10 9 2 13 16 13 10 15 13 15 9 1 15 9 2
26 1 15 3 9 13 2 16 1 0 9 2 10 15 9 15 9 13 2 1 13 0 7 0 13 9 2
22 1 15 9 7 9 3 13 0 2 1 9 13 9 1 9 7 9 13 9 1 15 2
7 9 3 9 0 3 13 2
2 0 2
15 9 9 9 3 13 13 16 15 9 0 7 9 0 13 2
12 3 3 9 13 9 9 16 0 7 0 13 2
13 7 0 7 0 13 9 2 7 1 15 9 9 2
22 16 3 9 2 13 9 10 2 9 13 9 0 9 2 13 16 9 13 0 7 0 2
38 16 7 3 9 13 0 16 13 9 9 7 3 13 9 0 2 16 9 7 9 2 3 3 9 13 0 16 13 9 9 7 3 13 15 7 15 0 2
8 13 3 16 9 9 0 13 2
2 3 2
16 16 9 13 15 10 9 2 3 13 10 13 2 16 13 4 2
26 7 1 15 16 13 10 9 13 16 1 15 13 10 9 13 16 1 0 13 9 2 16 1 13 4 2
16 3 13 16 1 15 9 13 10 9 9 16 1 0 9 9 2
18 15 7 3 13 16 15 0 9 13 2 1 1 15 15 13 9 13 2
9 0 13 3 15 0 9 3 13 2
2 3 2
40 1 10 9 13 15 0 13 16 9 0 1 0 15 13 7 3 13 0 2 9 0 9 15 13 1 0 2 7 13 3 9 15 2 16 13 1 9 7 9 2
17 3 12 9 9 15 13 1 10 15 12 9 9 13 7 1 0 2
11 7 9 0 1 9 13 0 16 1 9 2
22 15 3 9 0 9 13 2 9 3 2 9 7 9 2 15 9 12 10 0 9 13 2
12 13 3 0 0 2 15 15 9 7 9 13 2
2 0 2
24 0 9 1 9 9 3 13 2 16 10 2 7 3 1 10 9 13 9 9 2 16 1 13 2
16 7 3 15 9 15 1 9 15 13 2 13 1 9 0 9 2
11 0 7 9 3 13 9 16 1 0 13 2
12 3 0 9 9 13 9 2 15 1 0 13 2
15 0 3 9 15 1 15 9 13 2 15 1 1 0 13 2
2 3 2
16 0 0 13 1 9 13 1 9 7 9 2 16 1 13 4 2
19 3 7 13 9 15 1 9 13 9 16 13 0 16 13 4 13 1 9 2
16 15 7 13 16 13 3 7 3 2 7 1 13 16 13 0 2
15 9 3 15 13 9 0 0 2 13 0 0 16 13 0 2
19 15 3 9 7 13 9 2 7 3 13 13 2 7 15 15 13 1 9 2
22 15 9 16 13 13 0 10 9 2 15 10 9 3 13 2 0 3 15 13 9 9 2
2 3 2
11 9 0 13 0 7 13 2 16 9 9 2
16 9 3 15 13 9 9 3 13 13 13 10 9 1 9 9 2
33 7 9 0 13 13 13 10 9 1 9 9 2 16 1 9 0 9 13 9 0 1 15 9 2 9 7 0 3 13 13 9 0 2
10 9 7 10 13 1 9 13 7 13 2
36 1 15 3 13 2 16 9 1 9 0 13 1 9 9 0 1 9 0 0 2 1 9 7 9 13 1 0 1 9 9 9 0 1 9 13 2
35 9 3 9 0 2 1 4 1 10 9 13 2 10 9 9 13 3 13 1 15 16 13 3 0 2 7 0 1 1 9 15 9 0 13 2
16 1 9 7 13 1 9 9 13 2 16 3 1 9 9 13 2
14 7 3 9 9 9 0 3 13 13 1 1 9 0 2
28 9 7 9 9 0 2 1 13 1 1 9 0 2 1 15 13 10 9 2 13 1 1 9 9 0 7 0 2
11 9 3 0 13 13 0 2 3 7 0 2
2 3 2
23 13 9 15 9 1 9 13 2 3 9 13 0 2 16 0 3 13 2 15 3 9 13 2
10 15 7 13 9 3 9 0 9 13 2
5 13 3 8 12 2
9 3 13 15 9 0 1 9 15 2
7 9 3 0 13 8 12 2
3 3 13 2
11 1 9 13 2 7 1 0 15 15 13 2
13 13 3 1 13 15 9 1 0 13 3 0 13 2
25 3 15 15 9 0 13 2 16 0 13 2 13 3 7 9 7 9 9 2 16 0 9 0 15 2
8 16 9 13 15 15 3 13 2
14 3 13 13 16 9 3 13 9 15 3 15 3 13 2
21 16 3 1 1 13 13 2 15 13 9 9 0 1 9 13 15 0 1 9 10 2
34 13 7 15 9 0 1 10 9 2 16 0 13 13 1 15 16 15 9 1 15 13 2 16 13 9 9 2 1 9 2 1 9 9 2
5 3 7 1 0 2
16 15 3 13 9 0 9 1 9 15 16 3 3 13 13 13 2
2 3 2
21 9 0 9 13 1 9 15 16 9 9 1 9 2 1 1 10 9 13 9 9 2
13 9 7 10 9 9 3 15 15 3 4 13 13 2
14 9 3 9 1 15 9 13 1 0 9 1 9 9 2
13 3 15 13 1 9 9 13 9 15 3 0 13 2
12 3 3 15 13 9 15 15 3 13 9 13 2
2 3 2
22 9 13 15 1 15 1 10 9 16 13 9 15 15 1 15 13 2 16 1 13 13 2
35 7 2 1 9 9 13 0 9 2 16 1 13 4 2 15 7 15 9 13 9 7 9 13 2 0 13 16 9 9 15 13 9 0 9 2
15 13 3 15 9 10 9 1 0 0 16 1 15 15 13 2
30 16 3 9 0 9 7 9 9 10 13 2 13 15 15 9 3 0 1 15 15 13 2 7 3 1 15 15 3 13 2
2 0 2
22 9 10 2 1 15 9 15 13 15 15 13 2 9 13 13 3 15 15 3 13 9 2
12 13 3 9 7 9 9 13 10 3 9 13 2
24 9 7 0 13 1 9 13 15 15 13 3 0 9 2 7 3 0 2 16 1 1 13 13 2
10 13 3 3 15 15 3 13 9 13 2
2 3 2
22 9 15 1 10 9 13 13 3 16 13 2 16 13 9 9 0 1 9 9 0 9 2
10 7 9 9 13 1 9 10 1 9 2
20 15 3 13 2 15 13 10 9 2 15 3 10 9 13 2 16 1 13 4 2
10 15 3 13 16 3 15 3 13 13 2
2 0 2
11 13 9 9 3 13 2 16 7 15 9 2
7 13 3 15 3 3 13 2
6 15 1 9 9 13 2
9 9 7 9 9 0 7 0 13 2
14 9 3 9 1 15 9 9 13 16 9 0 1 0 2
45 3 3 15 0 15 9 0 13 2 15 3 13 15 9 0 2 2 15 3 9 13 9 9 2 7 15 0 15 1 0 13 2 15 3 9 0 2 7 9 1 0 13 2 13 2
20 3 2 1 9 9 3 13 2 9 2 15 3 1 9 13 2 15 9 13 2
17 3 2 1 0 9 3 13 2 15 9 7 9 9 0 13 9 2
8 15 9 3 1 9 13 13 2
27 9 3 1 9 13 2 16 0 13 2 3 3 15 9 15 1 9 13 3 2 9 3 9 9 9 13 2
18 9 0 2 15 13 1 9 2 1 15 9 1 9 13 0 9 13 2
24 15 3 1 15 9 9 13 2 13 0 3 0 15 2 16 9 15 9 9 13 13 7 0 2
16 0 7 3 13 15 0 13 16 15 2 16 9 9 3 13 2
18 15 3 1 15 9 9 13 2 0 9 1 15 10 9 13 3 0 2
12 7 3 15 15 9 9 13 2 3 13 13 2
15 13 3 16 15 15 1 9 9 3 13 2 9 9 13 2
12 1 15 3 9 13 16 9 3 13 9 13 2
12 3 3 10 3 13 15 13 9 1 15 9 2
18 15 3 15 3 13 7 13 7 13 2 1 9 13 3 15 9 0 2
18 3 3 13 15 16 13 0 1 15 2 7 16 13 0 1 9 0 2
13 15 3 1 15 13 1 9 13 1 9 0 9 2
29 15 0 15 13 0 2 13 7 0 15 2 13 9 1 16 13 1 10 9 2 7 1 0 9 2 7 1 15 2
7 7 15 9 13 9 9 2
37 3 3 9 9 15 1 15 3 13 2 13 0 9 15 13 1 10 9 2 7 3 15 15 13 1 15 2 16 15 9 13 0 10 9 10 9 2
11 7 3 9 15 9 9 13 1 9 10 2
15 3 10 9 13 0 1 0 15 3 13 7 13 7 13 2
15 15 3 13 9 9 15 9 2 1 15 13 9 1 9 2
15 9 3 15 9 15 13 1 15 2 4 1 15 0 13 2
26 3 3 3 13 13 9 16 15 9 13 9 2 7 1 9 9 2 7 1 9 10 2 7 1 15 2
6 15 9 9 3 13 2
12 15 7 15 13 4 3 9 0 9 9 13 2
5 13 3 8 12 2
11 9 9 10 2 16 13 2 13 4 10 2
7 3 7 1 9 13 10 2
4 7 8 12 2
8 16 15 13 1 9 13 15 2
57 13 7 1 13 16 3 13 13 2 16 15 13 2 9 0 0 13 2 16 13 15 1 9 0 3 2 16 15 13 9 15 2 3 16 15 2 7 16 13 1 9 2 1 13 4 16 0 9 15 13 1 0 16 13 1 15 2
7 16 9 13 0 13 0 2
23 1 15 7 3 0 13 13 16 13 0 1 0 9 0 9 13 2 7 3 13 13 13 2
19 13 3 9 9 3 13 16 1 16 0 13 2 3 7 1 16 0 13 2
21 13 3 2 1 0 13 2 13 3 13 2 7 3 9 13 15 0 13 13 13 2
10 13 3 16 3 13 15 0 13 13 2
14 1 15 7 0 13 2 1 15 9 3 13 3 13 2
23 13 7 1 0 3 13 2 7 15 3 3 13 1 13 16 0 13 2 7 16 0 13 2
17 3 15 9 9 13 1 15 13 13 9 2 16 15 9 13 13 2
15 10 3 9 15 1 13 13 16 0 13 2 0 13 13 2
23 0 7 9 9 1 0 13 1 15 15 15 9 9 13 16 0 13 2 16 1 13 4 2
14 13 3 16 1 13 15 13 9 1 0 9 0 13 2
2 3 2
12 13 1 0 13 1 16 15 1 10 9 13 2
16 13 3 3 1 10 9 13 16 3 13 1 15 13 7 13 2
10 0 0 3 13 1 10 9 16 13 2
51 1 15 0 16 15 15 1 15 13 2 3 13 3 1 9 2 1 15 13 0 2 16 1 13 2 1 15 16 1 15 13 2 3 13 9 7 3 9 2 7 0 9 2 16 1 0 13 13 3 13 2
26 0 7 9 1 0 13 9 3 0 1 9 15 13 1 9 10 2 7 3 1 9 15 13 1 15 2
12 15 3 13 15 13 0 9 1 13 7 0 2
2 0 2
17 16 1 9 0 0 13 9 2 3 1 9 13 0 16 3 13 2
26 7 2 1 9 13 10 2 16 1 1 13 13 2 13 3 0 9 13 2 7 3 15 15 13 13 2
11 13 3 1 9 16 13 13 7 3 13 2
2 3 2
14 9 13 10 9 9 3 13 2 3 3 1 15 13 2
23 3 2 1 1 15 1 9 9 13 2 13 3 16 0 3 1 9 9 13 2 7 9 2
17 16 7 1 15 9 13 9 9 2 3 0 9 13 9 9 13 2
15 15 3 13 15 1 15 13 13 1 15 9 0 9 13 2
2 3 2
10 9 3 13 13 0 15 9 13 13 2
7 13 3 9 13 13 9 2
10 9 7 0 9 13 7 0 7 13 2
36 16 3 0 13 13 2 15 9 13 13 13 2 3 16 9 13 0 13 2 16 9 3 0 13 2 16 9 9 13 0 2 1 9 0 13 2
17 9 7 9 2 16 13 9 9 13 1 15 2 13 3 9 13 2
15 15 3 9 13 9 3 13 2 1 13 9 0 13 13 2
2 3 2
19 9 9 0 3 13 7 9 16 3 15 9 9 13 16 9 15 13 13 2
30 9 7 2 1 13 9 15 9 2 15 13 9 2 13 15 9 3 0 1 15 2 7 3 1 9 1 15 10 9 2
14 9 7 13 1 10 9 0 13 16 13 1 15 13 2
9 13 3 9 15 13 7 13 13 2
12 3 3 0 9 9 7 9 9 9 3 13 2
14 13 3 1 13 3 9 9 13 1 9 13 13 13 2
19 3 3 0 9 0 9 13 2 1 13 1 9 0 0 9 0 13 13 2
21 9 7 1 9 13 3 13 0 15 9 2 16 1 15 13 2 7 13 15 0 2
23 3 3 13 2 16 15 15 13 1 9 13 13 13 2 16 15 9 13 13 7 15 13 2
24 1 13 3 13 16 2 16 10 9 9 0 0 13 2 1 15 1 10 9 15 0 13 13 2
42 3 2 1 13 2 9 13 2 7 13 2 15 0 2 0 15 13 1 0 9 7 9 13 2 3 9 1 15 13 9 2 9 15 15 15 1 9 13 13 13 0 2
21 3 7 13 0 9 0 9 2 15 2 1 9 9 13 2 1 10 0 15 13 2
44 9 15 2 16 9 9 1 0 13 2 3 13 13 15 13 13 3 3 13 2 16 9 13 9 15 13 16 13 3 13 2 7 3 13 13 1 9 16 3 1 10 9 13 2
25 15 13 2 3 13 13 9 9 2 16 15 3 13 2 3 13 2 3 1 15 9 2 3 13 2
28 9 3 13 1 15 16 9 1 15 13 2 13 9 2 7 3 9 13 2 15 13 1 13 2 9 13 2 2
17 3 9 9 13 7 0 1 0 9 13 2 15 3 15 3 13 2
8 7 1 15 13 1 9 13 2
30 3 2 16 15 1 9 13 16 0 13 2 3 0 13 13 15 9 13 2 16 0 13 9 13 1 15 16 13 13 2
25 15 7 3 0 13 0 2 7 2 16 1 15 13 2 9 13 2 7 1 9 2 7 9 9 2
12 15 3 0 13 0 2 16 13 13 2 13 2
43 3 7 2 16 0 1 0 13 2 16 13 2 15 13 13 2 0 13 13 2 13 15 1 9 13 2 7 13 2 13 0 2 1 9 0 13 2 7 13 2 13 0 2
23 7 3 1 15 2 7 1 10 0 15 9 9 1 13 13 13 2 1 9 7 9 13 2
13 16 7 9 0 13 13 2 3 9 9 0 13 2
9 13 3 8 12 2 1 0 9 2
13 9 7 9 13 16 13 2 7 9 9 7 9 2
11 7 8 12 3 13 15 13 1 9 15 2
7 1 9 1 1 9 13 2
4 7 9 12 2
5 13 15 1 3 2
6 16 13 2 13 15 2
6 16 9 13 9 9 2
12 3 13 13 16 9 9 9 7 9 9 13 2
20 10 3 15 15 9 13 13 1 9 2 16 10 9 13 2 16 1 13 4 2
13 9 7 15 13 1 9 2 15 1 9 1 9 2
14 13 3 9 10 3 9 9 2 7 15 1 15 13 2
12 9 7 1 9 13 15 13 1 9 7 9 2
13 13 3 16 9 15 15 13 1 9 7 9 13 2
2 0 2
15 3 9 13 10 9 15 13 2 16 1 9 9 13 9 2
15 10 3 9 13 2 10 9 13 2 1 15 10 9 13 2
8 13 7 1 9 9 7 9 2
45 3 2 1 9 15 13 1 10 9 2 1 15 13 15 9 9 2 13 0 9 15 9 2 1 15 13 3 10 9 2 10 9 9 13 2 1 9 9 0 1 9 0 0 13 2
9 13 3 9 7 9 7 9 9 2
2 3 2
27 16 9 10 13 0 7 1 15 10 9 9 2 3 10 13 13 0 2 7 1 15 10 0 9 0 9 2
23 16 3 9 13 10 9 13 9 15 9 2 3 13 10 13 7 13 13 10 9 7 9 2
2 3 2
26 9 3 0 13 9 1 16 1 15 13 2 7 3 1 16 13 1 9 10 2 16 1 1 13 13 2
8 13 3 9 9 1 10 9 2
22 7 0 13 1 9 1 9 7 9 9 2 16 9 0 13 1 10 9 1 9 9 2
27 16 3 9 0 13 15 10 9 1 10 9 0 2 3 9 1 9 13 9 9 2 1 15 13 10 9 2
11 7 0 9 13 1 10 15 1 13 13 2
8 13 3 9 7 9 7 9 2
2 3 2
28 9 3 0 13 9 0 16 15 2 7 15 2 9 0 2 1 9 0 13 3 0 2 13 3 1 9 13 2
14 9 7 7 9 9 0 13 7 1 9 7 1 15 2
38 1 3 9 9 13 1 9 15 15 2 9 7 13 15 9 15 1 15 2 3 7 15 9 9 0 9 0 13 2 13 16 9 9 7 9 9 13 2
7 15 7 9 9 0 13 2
5 13 3 1 9 2
6 13 9 7 9 9 2
3 8 12 2
6 9 7 9 1 9 2
6 3 3 9 9 9 2
3 8 12 2
7 15 13 15 13 1 9 2
32 9 7 15 13 9 1 10 9 2 1 15 1 15 13 9 13 7 3 13 2 13 9 9 1 12 2 7 9 9 0 13 2
15 3 7 13 9 0 9 2 1 15 13 15 9 7 13 2
27 7 3 13 9 1 9 0 2 15 9 13 2 9 9 9 2 16 3 9 2 15 13 2 3 13 13 2
5 16 9 13 0 2
9 1 15 13 13 16 9 0 13 2
16 13 3 15 13 9 9 15 1 15 13 2 16 1 0 13 2
11 15 7 13 9 0 2 16 0 13 9 2
8 13 3 10 15 15 13 9 2
5 13 3 0 0 2
2 3 2
12 9 10 9 9 13 2 16 1 1 13 13 2
21 9 7 3 13 13 9 16 13 10 1 15 13 2 1 1 15 9 9 3 13 2
18 10 7 9 2 1 13 0 2 16 13 4 1 2 1 0 15 13 2
6 13 3 9 0 9 2
2 0 2
29 16 9 9 1 10 15 13 15 15 9 13 2 16 13 4 2 13 16 3 0 13 9 9 2 7 3 9 9 2
20 7 1 9 0 13 0 1 9 2 16 3 9 2 16 9 13 1 12 9 2
26 13 3 9 0 2 16 9 2 15 13 9 9 2 0 9 9 13 16 13 15 13 1 15 1 9 2
7 13 3 9 9 10 9 2
2 3 2
10 9 9 10 16 15 0 0 15 13 2
35 7 1 13 9 0 2 16 1 13 4 2 1 15 0 13 0 13 9 13 2 16 7 15 12 15 2 7 0 0 13 9 0 13 13 2
13 7 3 3 13 0 9 15 15 13 15 13 13 2
10 15 3 13 15 1 9 10 0 13 2
2 3 2
6 9 9 13 10 13 2
17 16 3 10 9 13 0 2 16 13 4 2 3 10 13 13 0 2
13 16 7 15 13 13 1 13 2 3 0 1 0 2
23 16 3 1 13 10 2 15 13 13 2 13 13 13 2 7 9 1 10 13 0 13 13 2
2 0 2
22 9 13 0 0 3 0 13 0 2 7 3 2 16 13 1 9 2 1 12 1 9 2
19 15 1 15 13 16 9 3 13 1 13 0 2 16 9 2 7 3 13 2
42 7 16 13 0 9 2 7 13 15 9 2 16 0 9 2 7 0 9 2 3 16 15 7 10 13 0 1 9 2 16 15 13 0 2 0 15 13 0 9 16 9 2
24 3 15 15 7 10 3 13 9 13 7 13 1 15 9 7 9 2 7 3 1 15 13 13 2
16 3 13 1 9 9 2 15 13 0 0 2 16 1 13 4 2
16 1 3 9 9 15 13 2 15 13 15 3 15 0 0 13 2
2 3 2
31 3 15 9 13 0 7 0 1 13 2 3 1 12 13 0 13 2 16 7 10 9 2 3 13 0 2 3 13 3 13 2
15 9 7 0 1 9 7 9 13 0 2 16 1 0 13 2
13 13 3 1 12 2 15 13 10 9 2 0 13 2
2 3 2
11 9 0 13 9 0 2 16 7 15 9 2
7 15 3 9 0 15 13 2
14 7 15 1 15 13 1 9 9 10 13 15 9 0 2
9 13 7 1 9 1 10 9 0 2
6 9 7 3 13 0 2
9 3 7 9 9 0 13 7 9 2
9 13 3 16 9 10 3 0 13 2
2 3 2
17 1 9 10 13 0 0 1 9 2 13 3 1 0 9 9 13 2
34 16 9 0 3 13 0 3 9 2 13 16 7 0 13 0 9 0 16 0 2 7 16 9 0 3 13 10 9 15 13 0 1 9 2
11 15 15 13 0 2 16 1 1 13 13 2
2 3 2
7 0 9 13 16 13 9 2
13 3 9 0 13 1 15 0 13 2 3 9 13 2
23 13 7 15 1 9 10 9 13 9 0 13 9 1 9 2 3 7 9 3 0 9 13 2
17 1 3 9 1 9 13 10 3 2 3 3 13 13 0 16 13 2
2 0 2
16 10 9 1 15 9 9 13 2 7 1 15 9 13 0 9 2
17 16 3 9 15 9 13 2 3 7 15 15 9 13 15 9 13 2
29 1 9 7 9 0 15 9 13 16 12 2 1 3 1 0 9 2 7 1 12 9 2 15 13 9 9 2 13 2
8 3 7 3 0 13 1 9 2
10 7 3 1 9 9 15 9 9 13 2
8 3 7 0 2 15 9 13 2
11 15 3 13 1 9 0 0 7 13 9 2
14 7 3 2 1 13 13 2 15 13 15 13 3 0 2
8 15 7 13 15 1 9 13 2
7 7 9 15 3 13 9 2
15 13 7 1 13 3 9 10 0 3 13 2 16 9 0 2
16 13 3 9 10 1 9 0 3 1 9 2 15 15 9 13 2
10 0 13 2 16 9 10 0 13 13 2
4 0 7 0 2
12 0 13 2 16 9 10 0 1 0 9 13 2
13 3 3 13 1 0 1 12 9 2 16 9 0 2
23 0 13 1 15 13 2 16 9 10 2 16 1 0 9 0 13 2 3 13 3 0 13 2
11 7 3 0 13 3 13 16 0 15 13 2
18 15 3 13 1 9 0 2 15 3 0 13 2 3 1 12 9 13 2
19 0 13 2 16 9 0 13 15 15 13 7 15 3 13 2 16 13 4 2
23 13 3 3 9 9 2 15 13 16 0 2 1 16 0 2 13 0 2 0 9 3 13 2
24 16 2 1 0 9 9 13 2 16 15 13 2 0 16 0 13 16 1 9 10 9 13 13 2
7 15 13 3 0 9 9 2
6 3 7 9 3 13 2
31 3 2 16 3 13 2 3 13 0 1 16 13 0 2 7 1 16 1 10 9 15 13 7 16 13 13 2 16 13 4 2
38 13 3 16 9 0 3 13 9 9 2 16 9 15 13 2 16 0 7 13 9 2 7 13 7 13 2 1 9 1 15 9 13 0 2 1 9 0 2
7 13 3 0 9 0 9 2
19 13 3 9 0 15 7 13 7 13 7 13 2 15 3 13 1 9 9 2
17 7 13 3 0 15 13 1 10 9 15 7 13 7 13 7 13 2
16 3 2 3 1 9 1 9 0 13 2 13 13 1 9 0 2
6 3 3 0 13 0 2
10 16 3 13 2 15 0 9 15 13 2
5 16 9 0 13 2
20 15 7 13 2 13 13 16 9 13 0 2 7 16 15 9 15 9 3 13 2
22 16 3 15 9 0 13 0 2 3 1 13 10 9 13 2 16 3 1 0 9 13 2
11 9 7 0 9 1 13 9 13 9 0 2
17 9 3 0 3 13 1 9 13 2 7 3 1 15 16 15 13 2
22 1 3 13 0 9 1 13 2 16 1 13 13 2 13 16 15 9 1 1 13 13 2
22 7 9 9 7 9 1 10 9 13 1 9 7 9 1 9 2 15 13 1 9 9 2
15 3 15 0 1 9 9 2 1 0 9 10 9 2 13 2
2 3 2
28 10 15 13 2 1 15 15 13 7 15 15 13 2 9 13 2 7 9 0 9 13 2 7 1 15 9 13 2
14 15 3 9 13 2 1 9 1 9 2 9 13 0 2
5 3 3 13 13 2
18 13 3 16 15 2 1 15 13 2 0 13 2 7 0 13 9 0 2
17 1 9 7 13 0 15 9 3 0 16 0 9 13 13 1 0 2
13 16 3 15 9 13 0 9 2 0 3 13 15 2
11 7 3 13 16 15 9 13 15 1 15 2
5 15 1 13 4 2
20 16 3 15 15 1 15 13 2 15 0 2 0 9 13 15 2 15 13 0 2
2 0 2
33 9 9 0 0 13 15 9 0 2 1 9 0 13 1 9 9 15 13 1 15 16 1 9 2 16 1 9 13 2 1 12 0 2
14 16 3 9 13 15 15 9 0 2 0 13 9 0 2
21 15 7 13 3 13 16 13 7 0 7 0 2 1 15 9 7 9 9 0 13 2
16 13 3 16 9 13 3 0 0 2 7 3 15 15 0 13 2
2 3 2
9 9 13 1 13 3 13 1 15 2
16 15 13 3 1 9 9 2 16 13 13 9 13 1 9 10 2
35 1 9 7 13 13 1 13 9 13 2 7 15 16 2 16 0 13 2 1 0 13 13 2 7 15 16 1 9 0 1 15 0 9 13 2
13 15 3 1 9 13 3 13 2 16 1 13 13 2
28 3 3 13 0 9 0 9 9 2 7 3 13 1 0 9 2 1 16 10 1 15 13 2 16 1 13 4 2
2 3 2
16 9 15 3 13 0 15 1 0 13 2 7 15 1 0 13 2
12 3 9 15 1 0 13 2 3 13 1 0 2
28 9 3 15 3 13 1 0 7 0 2 3 13 13 0 2 7 15 15 1 0 3 13 2 16 1 15 13 2
14 3 15 9 13 0 7 0 2 7 15 9 13 15 2
9 3 2 9 0 2 9 0 13 2
7 1 9 7 3 13 3 2
11 3 15 9 7 9 15 7 10 15 13 2
14 3 3 15 9 15 9 13 1 15 16 15 0 13 2
25 15 7 13 15 13 8 12 1 0 9 2 16 13 3 1 10 9 2 7 15 13 13 1 15 2
16 13 7 1 13 16 9 15 1 13 13 2 13 9 3 13 2
21 9 3 9 13 1 15 1 15 0 9 13 2 7 3 1 10 15 1 9 13 2
19 1 0 3 9 2 1 15 2 13 3 0 0 1 9 2 7 3 9 2
21 3 9 0 9 10 13 1 0 9 1 1 9 1 9 2 15 13 0 1 9 2
15 3 7 1 0 9 13 9 9 3 1 0 13 3 13 2
19 0 3 9 13 0 1 9 13 2 1 15 10 13 2 16 1 13 4 2
13 13 3 16 15 9 3 13 9 9 1 12 0 2
21 3 3 13 13 16 0 9 3 13 15 1 15 15 13 10 9 9 3 0 13 2
28 7 1 15 9 13 16 0 0 13 16 13 2 16 3 13 15 9 0 7 0 2 7 0 9 9 0 13 2
5 16 9 13 9 2
9 3 13 13 16 9 13 3 9 2
8 9 3 13 2 9 13 13 2
11 7 9 13 10 0 9 2 15 9 13 2
5 13 3 9 9 2
2 3 2
8 0 9 1 9 3 13 0 2
11 15 3 3 13 1 9 2 7 3 13 2
17 9 3 15 13 0 2 3 13 9 2 7 3 1 9 9 13 2
30 16 3 1 9 2 1 10 0 9 2 13 10 9 9 2 16 1 13 4 2 13 16 1 15 13 9 15 9 13 2
7 7 3 13 3 9 0 2
2 3 2
5 0 13 9 9 2
11 1 15 3 15 9 13 0 16 0 13 2
15 0 7 3 0 13 9 13 0 2 7 3 9 13 0 2
17 16 3 0 13 13 15 13 2 3 0 13 3 13 15 3 13 2
9 9 3 9 3 1 9 9 13 2
18 7 2 1 0 9 13 9 1 9 2 3 13 15 13 15 0 9 2
6 13 3 15 9 9 2
2 0 2
10 9 13 9 9 2 16 1 13 4 2
7 7 1 9 9 13 9 2
9 13 3 13 15 12 3 13 15 2
13 3 7 0 2 15 15 13 2 0 15 9 13 2
16 9 15 0 9 1 15 13 0 2 16 2 15 9 13 9 2
5 13 3 9 9 2
15 9 7 9 15 13 1 9 13 2 16 1 12 8 13 2
4 13 3 9 2
14 7 1 13 9 2 15 15 13 15 16 9 13 9 2
2 3 2
26 16 9 13 10 9 9 2 16 1 13 4 2 7 3 1 15 9 13 7 13 2 13 16 13 0 2
21 3 16 15 9 9 13 0 2 7 16 9 9 13 0 2 16 13 1 12 0 2
13 7 1 0 13 9 9 7 9 2 16 3 13 2
7 3 13 16 9 13 9 2
5 7 1 13 9 2
2 3 2
15 9 13 3 0 9 2 7 3 9 2 16 1 13 4 2
30 9 7 2 1 13 9 1 9 2 13 9 3 13 16 13 1 15 15 9 15 13 2 16 7 1 10 15 9 13 2
11 13 7 15 9 9 7 1 9 7 9 2
10 15 3 13 13 2 13 3 3 13 2
5 3 9 13 9 2
7 7 3 13 1 13 9 2
2 3 2
14 16 9 13 15 15 1 15 2 0 13 15 13 0 2
16 15 7 13 9 0 2 1 15 16 1 9 10 0 9 13 2
28 1 9 7 0 13 15 15 13 1 13 9 15 13 1 15 15 13 2 16 13 1 15 15 13 9 1 9 2
6 3 3 9 9 13 2
4 13 3 9 2
2 3 2
37 1 15 9 9 3 13 1 15 15 1 15 9 13 2 3 1 9 15 13 1 9 2 7 1 9 2 1 16 1 9 9 3 15 1 9 13 2
16 15 7 3 13 1 9 2 16 0 13 2 16 1 13 4 2
8 15 3 13 16 9 9 13 2
15 15 7 13 15 13 8 12 2 16 9 9 3 13 9 2
4 8 12 13 2
6 9 7 9 1 9 2
4 7 1 9 2
8 13 10 1 15 3 4 13 2
5 7 9 12 13 2
12 15 13 9 9 2 7 13 9 2 3 13 2
19 13 7 16 1 9 9 7 9 15 15 13 9 0 2 7 15 9 10 2
31 3 1 9 10 0 9 1 0 9 0 13 7 0 2 15 15 13 1 9 13 1 9 0 2 1 15 13 9 1 9 2
30 3 7 9 13 13 2 16 1 9 1 15 9 3 15 13 2 16 16 9 13 1 9 2 3 3 9 1 9 13 2
37 7 16 9 13 1 9 9 2 3 9 13 9 2 15 9 13 9 1 9 2 13 16 9 10 13 15 9 13 9 2 16 4 13 13 1 9 2
15 16 3 13 13 16 1 15 9 9 13 9 9 7 9 2
20 9 7 0 2 15 15 9 13 1 9 2 3 13 9 13 9 7 15 15 2
27 3 16 13 15 1 9 15 3 13 15 2 13 1 9 16 9 15 1 15 9 13 16 9 9 1 9 2
13 3 13 16 15 13 0 1 9 15 13 10 9 2
11 7 1 13 16 13 15 3 16 0 13 2
12 13 3 15 2 13 15 2 16 1 13 4 2
10 3 0 7 9 2 7 9 7 9 2
23 7 15 13 9 9 15 9 13 1 12 1 9 2 13 2 7 3 9 13 2 7 0 2
5 0 3 3 13 2
11 13 7 9 13 13 2 7 13 1 15 2
22 16 0 15 3 13 0 2 3 1 9 2 2 15 13 2 7 9 13 2 7 0 2
25 7 13 13 9 9 2 15 13 16 1 15 13 16 9 15 13 3 1 9 2 15 9 13 9 2
29 7 9 13 16 3 13 9 1 15 16 13 1 9 1 15 15 2 7 1 15 16 13 15 7 13 3 1 9 2
32 3 13 16 2 16 9 15 9 15 13 16 2 13 15 2 3 13 15 9 2 15 13 0 9 2 15 9 13 9 7 9 2
33 16 9 15 13 15 3 13 15 9 13 2 1 9 7 10 13 4 13 13 1 15 2 7 3 15 15 13 9 0 15 9 13 2
6 7 1 13 7 0 2
18 3 2 13 16 9 15 0 13 2 13 9 15 13 15 3 13 9 2
28 7 16 2 13 15 2 13 9 1 15 13 4 13 9 2 0 13 16 13 9 13 2 7 9 13 0 9 2
34 13 3 16 2 16 9 1 9 9 13 15 13 15 2 16 1 13 4 2 3 3 3 13 16 15 9 13 0 16 1 9 13 9 2
8 3 9 13 3 9 9 9 2
17 3 13 9 1 9 16 9 1 10 9 2 3 16 9 1 9 2
14 7 3 1 9 9 0 13 16 9 1 9 9 13 2
11 16 9 3 13 13 16 16 13 9 9 2
8 3 1 15 0 9 13 0 2
13 3 15 2 15 13 1 9 2 15 13 1 9 2
5 16 9 13 13 2
16 13 15 15 1 0 9 9 13 2 3 13 13 1 9 9 2
13 1 15 3 16 9 13 13 2 13 16 13 13 2
20 1 3 9 13 13 9 0 9 2 13 16 9 13 2 16 3 2 13 13 2
6 13 7 13 1 13 2
13 0 13 3 16 13 9 2 16 3 2 13 13 2
5 9 7 13 9 2
19 1 3 13 9 13 2 16 1 1 13 13 2 13 9 3 1 9 9 2
4 13 3 13 2
2 3 2
31 15 13 15 9 2 13 1 15 9 9 1 15 15 13 1 9 9 2 16 9 0 1 10 9 13 15 0 7 15 0 2
20 1 13 7 7 13 13 9 9 13 7 0 2 1 10 9 13 1 15 9 2
21 13 3 13 9 13 7 13 1 15 15 13 13 7 0 1 16 13 1 9 9 2
11 3 7 15 13 1 15 16 13 7 13 2
30 3 1 15 3 13 9 9 1 13 7 13 2 16 13 7 13 13 1 16 9 13 1 9 7 9 2 1 9 15 2
17 13 7 9 13 7 13 1 9 15 13 1 9 1 9 7 9 2
9 3 10 13 7 9 13 7 13 2
7 9 3 0 1 9 13 2
11 1 3 9 13 13 2 13 16 13 13 2
2 0 2
12 15 15 13 10 9 2 13 9 16 13 9 2
16 15 7 13 3 2 13 16 1 15 0 13 15 13 0 9 2
12 15 7 9 13 13 10 9 7 9 10 9 2
23 15 3 1 10 9 2 0 3 1 9 2 0 1 0 9 2 13 0 9 1 9 0 2
10 15 3 15 13 2 7 15 3 13 2
18 3 15 15 3 13 2 0 9 10 9 9 13 1 13 15 15 13 2
8 15 7 13 2 13 1 15 2
13 15 3 0 9 2 15 9 13 2 13 3 13 2
19 1 3 15 13 13 2 13 15 9 2 15 13 15 10 9 7 10 9 2
2 3 2
11 13 2 3 9 13 2 3 0 13 13 2
15 7 9 13 2 7 10 13 13 9 2 16 1 13 4 2
6 3 13 13 15 0 2
15 9 7 0 13 1 9 2 16 9 0 13 1 9 9 2
6 13 3 1 9 9 2
2 3 2
27 9 1 9 13 3 13 7 15 13 16 13 9 2 15 9 13 9 7 9 2 1 15 13 15 1 13 2
12 3 9 0 3 13 2 7 9 0 1 9 2
12 7 9 9 0 13 9 9 7 9 1 15 2
10 13 3 9 1 9 2 16 1 13 2
7 13 3 16 15 13 13 2
2 3 2
12 1 9 9 2 1 13 9 2 0 13 9 2
9 3 9 10 9 13 1 10 9 2
15 13 3 16 13 2 7 13 16 13 2 7 3 1 15 2
39 7 15 13 16 9 15 13 9 2 2 16 9 2 3 1 9 9 0 7 13 2 7 1 9 9 0 2 13 9 2 13 15 10 9 2 15 13 9 2
8 0 3 13 13 0 13 9 2
2 3 2
7 0 13 15 15 9 13 2
11 7 3 0 13 9 15 15 13 1 15 2
8 9 7 0 13 9 1 13 2
12 16 3 0 13 15 2 13 0 13 15 9 2
16 0 3 9 0 13 1 9 13 2 15 0 13 1 15 13 2
2 0 2
36 9 7 9 1 9 3 12 9 13 1 9 2 3 7 9 0 2 15 13 13 9 2 13 1 15 9 1 9 2 3 1 0 7 1 0 2
41 3 9 9 1 15 9 13 2 13 9 9 15 13 1 9 2 15 13 9 9 2 7 9 9 13 15 13 2 13 15 9 1 9 9 13 2 15 13 9 9 2
10 9 7 15 13 3 15 9 16 15 2
11 15 13 0 0 2 15 0 1 13 4 2
11 15 13 3 0 9 1 9 15 13 15 2
30 15 3 3 0 13 9 0 2 7 13 2 16 3 13 2 15 9 2 7 9 0 2 1 13 13 2 15 13 9 2
6 13 3 1 9 9 2
9 15 7 9 9 9 0 9 13 2
5 13 3 1 9 2
7 10 15 13 2 9 13 2
4 7 8 12 2
5 9 15 15 13 2
7 16 9 9 13 15 9 2
14 1 15 7 13 16 10 9 3 13 15 16 10 9 2
13 9 3 13 13 13 16 13 13 2 16 13 4 2
12 13 7 13 1 9 10 2 16 1 13 4 2
4 3 7 13 2
8 13 3 9 9 15 15 9 2
2 3 2
11 16 13 13 9 13 2 3 7 13 13 2
18 15 3 13 9 1 9 13 2 3 7 13 1 15 13 2 16 9 2
24 7 13 9 13 15 9 2 16 1 13 4 2 15 16 15 13 9 13 2 16 1 13 4 2
8 13 3 7 0 13 9 15 2
8 3 7 9 9 13 15 9 2
2 0 2
22 1 10 9 13 16 9 13 2 13 16 9 2 15 13 9 0 2 1 10 9 13 2
7 13 7 13 15 9 9 2
10 13 3 16 9 1 9 10 13 13 2
7 10 3 9 13 10 9 2
2 3 2
45 16 9 13 15 13 0 9 2 1 0 9 13 15 13 1 9 2 13 16 9 13 15 16 9 9 2 13 16 0 9 13 1 15 16 9 1 9 2 7 16 13 9 1 9 2
6 15 10 1 13 4 2
13 3 13 3 0 16 0 9 13 15 13 0 9 2
8 16 0 13 9 13 0 9 2
14 1 15 7 0 13 16 0 0 9 13 13 15 9 2
11 9 3 13 13 9 9 2 16 13 4 2
16 15 7 15 1 9 0 13 13 0 9 2 16 1 13 4 2
12 0 3 9 13 15 1 15 0 13 0 9 2
2 3 2
14 0 13 1 9 16 13 1 13 2 16 1 13 4 2
16 7 0 15 13 13 1 9 2 1 9 13 1 9 0 9 2
26 16 3 9 0 13 15 0 13 16 15 9 9 2 13 16 15 15 13 0 0 9 2 15 15 13 2
6 15 0 1 13 13 2
2 3 2
52 0 13 13 15 13 9 13 2 1 3 13 2 13 13 16 13 2 9 15 13 13 2 7 16 13 2 3 13 13 2 13 1 9 9 16 13 1 9 0 2 15 13 0 13 2 15 13 9 13 1 15 2
19 16 3 9 15 15 0 13 16 15 2 13 16 15 15 13 15 9 13 2
11 7 10 13 13 10 9 2 16 13 4 2
8 3 15 15 13 15 9 13 2
7 15 13 1 9 0 9 2
2 3 2
9 15 13 0 13 13 10 0 9 2
14 3 9 4 1 15 13 2 7 1 15 15 13 13 2
17 0 7 9 13 15 9 2 16 15 13 0 9 2 16 13 4 2
8 15 3 13 0 13 10 9 2
2 0 2
10 15 9 1 10 9 0 1 9 13 2
18 3 9 9 1 9 13 2 16 13 1 9 2 1 12 9 7 9 2
17 9 3 1 0 13 10 0 9 2 7 0 9 2 7 3 9 2
11 0 7 9 15 1 0 13 16 15 9 2
9 3 0 9 0 9 13 9 0 2
40 1 7 9 0 13 9 13 7 10 15 15 1 15 13 13 2 0 13 0 16 15 9 0 13 15 13 2 15 13 2 15 13 12 2 7 15 15 13 3 2
10 16 9 2 13 15 2 13 3 15 2
13 15 7 13 13 16 2 13 15 2 13 3 15 2
18 15 3 13 13 9 0 2 15 13 13 15 15 13 1 9 9 9 2
14 13 7 15 9 0 9 9 2 16 1 13 15 13 2
20 1 15 3 16 13 15 13 2 3 15 13 2 15 1 15 16 1 9 13 2
2 3 2
15 15 15 15 4 1 15 1 15 13 7 13 2 9 13 2
20 15 3 1 15 13 2 13 13 0 2 7 3 13 7 13 2 3 0 13 2
11 15 7 9 9 10 1 15 13 7 13 2
29 3 7 1 15 0 7 0 13 2 16 1 1 13 13 0 2 7 0 0 13 1 10 9 2 15 1 0 13 2
16 13 3 9 9 9 1 15 16 10 9 7 9 13 7 13 2
2 0 2
31 15 13 15 1 15 7 1 15 2 13 1 13 10 1 15 15 13 2 16 15 13 9 1 15 2 13 16 10 0 13 2
18 7 9 10 9 1 15 7 1 15 13 7 13 2 16 1 13 4 2
18 10 7 15 9 13 15 10 9 1 9 9 2 16 1 13 15 13 2
19 13 3 16 9 2 1 15 15 16 13 7 13 15 2 13 7 13 15 2
2 3 2
12 9 2 13 15 2 13 10 15 1 15 13 2
15 10 7 3 13 1 15 1 0 9 2 16 1 13 4 2
10 9 3 2 13 15 2 3 15 13 2
2 3 2
23 3 15 13 9 9 2 3 10 9 1 0 15 13 7 1 3 13 2 16 1 13 4 2
12 9 7 9 1 15 13 16 1 15 15 13 2
20 3 3 9 13 9 7 3 13 2 3 9 13 9 1 0 13 9 9 15 2
11 0 7 9 13 9 1 9 9 7 9 2
29 3 13 10 9 0 1 0 2 16 1 15 0 4 13 2 7 0 1 9 2 15 15 1 15 10 9 9 13 2
2 3 2
4 9 13 9 2
13 7 9 9 10 13 15 0 7 1 15 13 15 2
15 3 0 0 13 15 2 7 2 13 15 2 13 10 15 2
7 15 7 9 0 9 13 2
5 13 3 8 12 2
13 13 3 10 15 13 2 7 15 15 13 15 13 2
10 16 9 12 9 9 15 7 15 13 2
15 15 7 13 2 13 16 9 12 9 9 15 7 15 13 2
34 10 3 9 12 9 2 7 12 9 2 13 1 9 7 1 9 0 9 2 16 15 9 13 9 7 9 2 15 13 0 9 1 9 2
36 1 7 15 13 1 9 3 2 15 15 1 9 13 13 9 13 1 9 2 7 3 9 13 1 15 16 9 0 1 9 2 16 9 1 9 2
24 1 3 9 10 15 13 1 15 16 1 9 2 16 13 4 2 12 9 9 13 15 7 15 2
2 0 2
14 15 9 13 7 13 2 1 15 10 9 13 7 13 2
22 9 7 9 13 3 0 1 16 1 15 13 2 7 3 1 16 15 13 0 1 15 2
11 15 3 9 13 9 2 15 9 15 13 2
24 7 3 13 13 15 9 9 13 15 13 15 7 3 13 15 9 2 1 1 15 15 13 0 2
16 15 3 9 15 9 13 15 2 13 15 0 7 15 1 15 2
15 15 0 1 15 3 13 16 16 13 15 2 16 13 4 2
19 13 3 16 15 7 15 3 15 7 15 9 9 13 2 7 12 7 15 2
2 3 2
25 16 1 1 13 13 2 1 9 0 9 9 13 1 16 13 13 9 2 7 1 15 1 9 13 2
23 16 3 1 15 9 13 9 15 9 13 2 3 13 9 2 16 3 16 15 13 1 9 2
23 16 7 9 15 13 1 9 1 0 2 3 9 1 15 15 13 1 9 1 0 7 0 2
20 3 16 9 13 1 9 2 3 1 9 13 9 7 9 15 15 13 1 9 2
20 16 3 15 13 13 9 7 15 15 13 1 9 2 13 15 9 1 15 9 2
14 15 7 1 9 13 13 0 2 1 13 1 10 9 2
16 13 3 16 3 2 7 15 9 9 2 9 13 15 7 15 2
2 3 2
25 1 9 3 13 15 2 16 15 9 13 15 7 15 15 2 13 16 3 13 1 15 12 9 9 2
4 15 13 0 2
10 3 12 0 9 3 13 3 12 9 2
2 3 2
13 1 10 9 9 13 13 1 13 16 13 1 13 2
29 16 3 13 15 9 9 0 15 13 15 1 15 2 0 1 9 15 13 15 2 1 15 13 15 15 13 0 9 2
4 15 13 0 2
2 0 2
10 13 9 13 10 9 2 16 13 4 2
9 7 1 9 3 13 16 12 9 2
8 3 3 13 3 16 12 13 2
2 3 2
8 13 13 9 1 16 13 13 2
32 16 3 12 9 13 15 7 15 2 16 9 10 13 0 10 2 3 12 9 13 15 7 15 2 16 10 9 13 9 10 9 2
8 16 13 9 0 9 3 13 2
15 1 15 7 13 16 13 9 3 13 9 7 9 0 9 2
6 3 9 1 9 13 2
24 16 3 13 0 15 9 13 13 1 15 15 9 2 13 16 3 13 1 15 12 3 9 9 2
5 15 13 1 13 2
2 3 2
11 13 4 16 9 15 13 16 13 9 10 2
13 15 3 9 13 15 1 9 15 13 1 9 15 2
8 7 10 1 9 15 12 13 2
22 13 3 15 1 15 1 9 15 2 3 0 0 7 0 13 2 16 1 1 13 13 2
10 13 3 16 9 13 3 13 0 9 2
2 3 2
18 0 9 7 9 13 0 9 2 16 15 13 0 9 2 16 13 4 2
16 9 7 13 3 13 9 1 9 0 2 7 9 1 9 15 2
17 3 7 9 13 13 7 9 1 9 0 2 7 9 1 15 9 2
2 0 2
42 15 1 9 7 9 13 2 16 9 13 1 16 13 13 15 9 1 13 2 9 7 3 2 7 1 0 1 16 9 13 1 9 0 2 15 13 13 7 1 15 13 2
15 7 1 15 9 7 9 2 15 13 9 2 13 1 9 2
21 0 7 7 0 2 15 13 9 2 13 1 9 2 16 9 13 2 1 12 0 2
21 15 7 15 1 0 15 13 2 3 13 9 15 2 1 7 9 13 0 9 9 2
10 9 3 13 1 9 3 13 15 9 2
9 16 0 9 1 0 9 15 13 2
42 1 15 3 13 16 3 13 15 13 2 1 13 9 0 2 16 13 15 9 1 15 9 2 16 13 15 13 9 9 15 13 1 15 13 2 3 7 13 15 1 0 2
10 3 13 13 1 9 13 1 9 13 2
13 3 7 13 0 9 16 13 13 1 0 3 0 2
10 13 3 9 0 7 0 3 9 0 2
16 3 10 9 3 13 16 3 1 0 7 0 15 1 15 13 2
2 3 2
20 9 9 1 15 13 16 9 13 1 9 1 9 0 2 15 13 9 13 9 2
20 7 3 0 9 9 2 7 7 0 15 1 9 0 9 13 2 16 7 9 2
9 9 3 9 1 0 9 15 13 2
2 0 2
14 1 9 2 1 12 8 2 0 9 9 13 1 0 2
20 12 3 1 16 15 0 13 1 15 15 13 1 0 2 16 9 13 1 9 2
14 15 1 16 9 0 13 1 3 2 16 7 9 9 2
7 0 7 9 13 1 0 2
26 9 7 2 1 15 16 13 15 16 9 13 2 13 15 15 13 1 15 16 1 9 2 16 13 4 2
19 13 3 9 9 15 0 1 15 2 7 9 9 0 1 9 10 1 3 2
8 9 7 9 13 1 0 9 2
6 13 3 3 0 9 2
2 3 2
20 16 9 3 13 0 9 1 15 13 0 2 13 16 1 0 13 9 9 9 2
37 3 13 3 0 16 15 9 0 10 0 9 13 1 9 0 2 7 0 0 9 15 0 2 15 9 13 2 15 1 10 9 13 2 16 1 13 2
20 16 7 9 0 13 0 2 13 0 2 16 13 16 0 3 15 0 13 9 2
9 13 3 16 9 3 0 9 13 2
2 3 2
9 9 13 2 16 3 2 13 13 2
12 7 9 13 3 0 9 2 16 1 13 4 2
6 13 3 3 0 9 2
21 15 7 9 9 13 2 15 2 9 12 2 1 0 9 9 0 9 13 2 13 2
19 13 9 9 16 13 0 2 7 0 1 15 9 2 7 3 1 10 3 2
11 13 9 10 15 13 2 7 13 3 0 2
9 16 9 13 3 15 15 3 13 2
23 16 7 13 13 1 9 13 1 13 2 9 15 13 13 16 9 3 13 16 15 15 13 2
18 3 0 13 3 13 2 7 2 12 13 2 13 15 2 16 9 13 2
18 16 3 13 13 1 9 13 1 13 2 15 13 13 16 15 15 13 2
2 3 2
11 9 13 1 13 2 16 7 9 7 9 2
19 3 7 13 13 3 9 9 2 7 9 2 7 9 2 16 15 15 13 2
10 3 7 13 13 13 16 15 15 13 2
35 1 15 7 13 0 13 2 16 0 13 13 0 2 16 7 10 9 2 7 3 13 16 15 15 9 13 2 16 15 13 15 3 3 13 2
21 13 7 1 15 15 16 15 15 3 13 1 15 2 13 1 9 7 1 15 9 2
19 3 15 13 3 15 15 3 13 1 15 2 9 13 1 16 1 15 13 2
7 15 7 3 13 0 13 2
16 3 1 15 13 15 13 15 13 2 16 9 10 13 1 13 2
41 16 3 0 9 3 13 1 13 15 3 13 16 1 16 13 1 15 7 1 15 9 2 13 16 9 3 13 15 15 16 16 13 15 13 1 15 7 1 15 9 2
18 15 7 3 13 13 7 16 9 3 15 3 13 13 13 3 1 15 2
54 3 2 16 9 13 1 9 13 1 10 9 2 15 13 9 13 2 9 7 3 0 13 9 13 1 15 2 7 3 1 0 9 2 7 9 13 1 13 3 0 1 16 13 1 13 2 7 3 1 16 13 1 15 2
31 13 3 16 2 1 9 13 13 9 2 13 16 15 13 13 9 9 2 16 7 9 15 0 13 9 13 15 13 9 9 2
11 9 7 13 1 13 13 13 1 9 15 2
11 1 15 3 13 13 1 13 16 13 15 2
48 3 7 0 13 13 9 1 16 13 1 15 2 7 1 16 13 1 0 9 2 16 3 0 13 9 13 1 15 2 16 13 15 13 1 9 2 7 15 13 7 13 7 13 4 1 0 9 2
35 16 3 3 9 15 3 13 16 1 13 2 9 3 13 9 13 1 15 3 16 13 1 13 2 7 16 13 1 0 9 2 15 13 13 2
29 9 3 0 9 13 1 9 3 13 1 16 13 1 0 9 1 15 9 2 7 3 0 1 16 13 1 9 13 2
24 13 3 9 9 15 3 13 3 2 13 1 15 9 2 7 3 0 13 1 16 15 15 13 2
25 7 13 0 1 9 13 1 13 2 7 13 1 13 2 7 13 1 13 2 7 9 1 13 9 2
8 3 13 13 9 1 13 13 2
8 3 3 13 13 15 1 13 2
22 7 13 7 13 7 13 13 9 13 1 0 9 2 1 15 9 3 9 3 13 13 2
11 16 9 1 9 13 10 9 7 10 9 2
25 1 15 7 15 1 13 4 2 13 16 9 1 9 13 10 9 7 10 9 2 7 13 0 13 2
23 13 4 3 1 16 9 13 10 9 7 10 9 16 0 9 2 15 13 15 9 13 15 2
19 1 10 3 13 13 10 9 7 10 9 2 16 9 1 10 9 13 9 2
9 0 13 7 9 3 13 15 9 2
7 13 3 13 1 9 3 2
11 15 13 0 2 1 10 13 13 10 9 2
11 0 13 3 16 13 10 9 7 10 9 2
2 3 2
22 15 13 1 9 13 10 0 9 2 16 9 1 9 13 10 9 2 7 13 13 9 2
14 7 9 13 15 13 16 0 9 2 16 1 13 13 2
13 0 3 13 15 13 2 7 13 13 15 3 13 2
2 0 2
16 1 0 7 1 0 9 15 9 15 13 16 9 0 1 0 2
23 16 3 1 9 13 1 0 9 2 3 1 0 7 0 9 10 13 7 13 1 9 13 2
18 7 1 0 9 1 9 13 0 9 0 2 15 0 15 9 13 13 2
13 3 9 0 13 9 0 2 16 3 13 0 13 2
19 7 3 2 16 0 9 3 13 15 9 16 15 2 1 9 13 15 13 2
2 3 2
15 10 2 16 13 2 13 9 2 15 13 0 7 0 9 2
13 10 7 2 16 13 2 10 9 0 13 10 9 2
9 0 3 3 9 10 9 13 0 2
13 9 7 15 13 1 15 13 2 16 1 13 4 2
8 9 3 1 9 13 15 13 2
2 3 2
18 10 9 7 9 15 1 9 13 2 9 13 0 2 16 1 13 4 2
16 13 7 9 13 0 9 0 9 2 1 1 15 3 9 13 2
6 3 1 9 0 13 2
6 3 1 9 13 15 2
6 7 3 13 15 13 2
10 16 9 3 1 9 13 15 1 15 2
36 16 7 0 9 13 0 9 7 0 9 1 9 2 13 15 13 16 3 15 1 9 13 2 1 10 15 13 13 10 9 2 16 1 13 4 2
12 7 3 0 13 13 16 3 13 15 1 9 2
10 13 3 15 16 13 1 9 10 9 2
20 9 7 3 1 9 13 1 15 15 13 1 9 2 16 9 1 15 13 13 2
25 3 3 13 0 9 2 1 9 9 15 13 1 13 2 15 9 13 0 1 15 3 13 0 13 2
31 1 3 0 9 1 15 13 13 2 3 7 1 15 15 15 13 2 15 13 15 9 16 15 13 1 15 16 13 10 9 2
2 3 2
20 1 9 13 13 0 9 9 2 15 1 9 13 13 13 9 16 13 9 9 2
38 3 2 16 9 15 2 16 3 2 9 13 2 3 9 7 9 2 15 3 3 9 15 13 13 1 9 9 15 9 13 15 13 2 16 3 1 9 2
11 13 3 9 15 13 2 3 15 3 13 2
24 0 3 15 0 9 2 1 15 9 2 3 13 13 3 13 2 15 3 13 13 0 9 9 2
7 15 7 15 13 1 9 2
16 13 3 9 2 1 15 9 2 13 3 13 15 9 1 9 2
10 7 1 9 13 9 1 15 10 9 2
8 10 3 1 15 13 0 9 2
12 13 3 9 13 3 13 15 9 15 1 15 2
10 3 3 1 9 13 13 15 1 15 2
2 0 2
16 9 2 13 9 10 2 13 13 15 1 15 16 9 15 13 2
24 1 7 0 9 13 0 2 13 0 9 0 2 7 15 9 16 1 15 9 15 3 13 13 2
31 16 3 2 1 15 16 13 9 10 2 13 1 9 15 15 15 13 2 13 16 13 13 0 9 2 0 9 13 10 9 2
24 15 13 13 0 2 16 2 16 13 2 13 2 1 10 9 13 9 13 9 2 16 1 13 2
11 3 3 1 9 13 3 15 15 3 13 2
2 3 2
20 0 9 2 1 15 16 13 1 9 2 13 1 9 15 1 9 1 9 13 2
15 0 3 13 13 9 13 1 9 2 7 3 13 9 9 2
21 7 9 15 3 1 9 13 1 9 2 3 13 0 15 13 1 15 16 13 9 2
13 1 9 7 13 15 3 1 9 2 16 1 13 2
14 3 3 0 13 16 9 15 13 1 15 16 13 15 2
2 0 2
13 9 13 1 9 16 9 1 9 2 16 1 13 2
17 7 9 2 16 13 15 13 9 2 3 3 1 9 13 9 13 2
11 3 7 9 1 9 13 15 1 15 13 2
34 13 3 13 3 9 15 1 15 1 9 13 2 3 7 1 9 13 2 1 3 2 1 15 16 13 7 13 15 2 13 7 13 15 2
5 15 7 9 13 2
29 16 3 13 13 15 2 13 1 15 16 13 15 13 15 9 2 16 1 15 15 9 13 16 13 15 9 1 13 2
16 7 16 13 15 13 2 1 15 13 16 13 15 9 15 13 2
14 13 3 15 7 16 9 13 2 7 16 1 9 13 2
18 13 7 10 1 9 2 16 1 15 13 13 2 1 9 13 0 9 2
18 3 7 0 9 1 9 13 15 13 2 15 1 15 13 16 1 9 2
13 7 1 15 0 13 9 15 13 2 3 7 13 2
28 3 7 10 13 15 1 9 15 9 13 13 2 10 7 13 15 1 9 15 2 1 15 13 2 15 9 13 2
13 9 13 1 9 16 9 15 1 15 3 0 13 2
14 13 3 13 9 16 9 15 15 13 3 1 9 13 2
19 16 3 9 9 9 15 13 3 13 3 1 15 2 13 15 1 15 13 2
12 10 7 9 15 13 1 15 13 3 1 9 2
8 3 1 15 9 13 0 13 2
7 13 3 9 9 1 9 2
17 3 3 13 9 9 2 1 15 15 13 9 2 16 1 13 4 2
2 3 2
27 16 9 1 9 2 16 3 2 13 4 13 2 16 15 13 13 13 3 13 2 13 0 0 9 13 0 2
2 3 2
13 16 0 13 9 15 1 13 10 13 2 0 13 2
8 0 7 15 1 15 13 13 2
17 3 3 1 15 13 13 15 1 9 7 0 2 16 1 13 4 2
2 3 2
49 16 15 13 1 15 0 15 13 3 3 1 12 16 1 15 13 16 1 15 13 2 13 16 9 7 15 15 13 1 15 1 15 15 13 2 15 0 1 13 4 2 7 16 1 15 13 1 12 2
13 7 3 13 15 15 0 2 15 15 13 1 12 2
7 15 7 15 0 13 13 2
10 1 15 3 13 15 9 13 13 0 2
17 12 9 2 1 9 15 2 15 9 2 1 9 15 1 15 13 2
18 1 9 3 15 2 16 3 13 4 10 9 2 1 15 1 12 13 2
31 3 15 1 9 9 13 2 7 13 13 9 1 15 2 16 13 1 9 13 2 15 3 13 4 9 1 15 1 15 13 2
42 1 9 7 15 1 15 13 2 13 15 9 1 15 9 16 9 9 9 1 15 13 2 7 3 15 13 13 2 16 9 2 15 0 9 13 13 1 15 9 0 13 2
31 15 7 1 9 9 3 13 2 7 3 1 15 9 2 16 15 13 13 2 7 1 15 13 1 15 2 15 1 15 13 2
11 3 7 13 1 0 9 9 15 1 15 2
17 3 9 15 1 15 15 13 2 1 3 15 9 10 9 4 13 2
10 3 3 13 9 15 1 0 9 13 2
5 0 7 7 9 2
91 16 3 1 0 9 15 13 9 2 3 3 1 9 15 13 13 1 10 13 16 13 1 9 1 15 2 16 0 13 13 9 15 7 3 13 9 2 7 3 13 13 9 15 13 2 3 0 1 15 7 3 1 13 2 7 16 13 3 13 0 9 1 0 9 2 15 13 0 9 0 9 2 1 9 15 3 0 2 7 0 0 13 16 3 13 0 9 9 1 9 2
73 3 1 13 2 9 13 15 13 2 0 13 13 0 3 0 2 7 0 2 15 9 15 3 13 15 0 1 15 9 2 7 16 3 0 13 13 7 0 13 13 2 16 9 13 1 12 8 2 16 0 13 12 9 0 13 0 0 2 3 3 1 15 9 2 1 1 0 3 13 9 7 9 2
10 9 3 9 13 9 0 9 3 13 2
9 15 9 0 13 2 12 8 12 2
7 9 1 9 9 3 13 2
28 16 7 0 9 1 10 13 3 13 2 3 3 13 13 16 15 15 13 2 16 16 1 13 1 15 0 13 2
48 1 3 9 13 9 16 0 9 13 2 9 7 0 3 13 0 1 15 9 2 1 15 13 10 9 2 16 9 9 1 15 13 1 10 9 9 13 2 3 13 9 9 0 1 15 0 13 2
24 9 3 0 13 3 0 0 9 2 15 13 9 15 2 7 3 15 9 2 16 1 13 4 2
16 15 3 13 16 9 15 0 9 7 9 2 3 16 15 9 2
19 7 3 9 0 1 15 13 16 10 9 13 2 3 16 1 10 9 0 2
9 2 3 7 7 1 10 9 13 2
34 16 2 1 1 15 13 3 0 0 1 9 2 15 9 13 1 15 2 1 7 13 1 15 0 1 9 15 2 3 0 1 15 13 2
10 3 7 0 9 13 1 10 13 0 2
11 3 3 13 1 13 0 15 1 9 13 2
22 9 3 10 12 7 15 9 13 15 7 15 2 7 9 15 1 15 13 0 7 0 2
24 9 7 15 1 15 13 1 9 15 2 3 3 0 7 0 2 7 0 7 0 2 7 0 2
13 15 3 0 13 2 7 0 7 0 0 13 13 2
10 16 9 13 15 15 1 15 9 9 2
23 1 15 7 13 13 16 2 16 9 1 13 15 0 13 0 2 13 3 15 0 1 9 2
8 13 3 4 0 9 0 13 2
16 1 15 7 0 2 16 3 13 15 2 3 13 3 3 13 2
12 15 3 13 13 15 15 15 13 3 7 0 2
20 16 3 0 9 13 0 2 13 16 15 13 2 0 13 1 9 15 15 13 2
2 3 2
5 10 0 13 0 2
9 9 7 13 15 13 4 13 0 2
11 16 3 9 10 2 3 7 13 9 13 2
4 13 3 0 2
16 7 3 0 13 2 16 9 9 3 13 0 9 1 15 13 2
6 3 13 0 1 9 2
2 3 2
6 15 9 13 2 13 2
11 9 3 15 3 13 2 16 7 15 9 2
17 7 3 13 3 3 13 15 13 13 2 16 3 13 13 10 9 2
8 3 3 13 3 13 15 13 2
24 13 3 0 1 9 15 13 15 13 2 16 7 13 2 15 7 0 0 2 7 0 9 13 2
2 0 2
40 15 13 15 2 0 13 15 15 0 13 1 15 2 16 13 1 9 15 9 2 7 1 9 2 7 16 1 0 9 15 15 13 1 9 13 13 1 15 9 2
7 15 1 9 13 3 13 2
43 16 3 9 2 13 15 2 13 15 15 1 15 2 0 13 15 13 10 15 15 1 13 1 15 1 9 13 2 16 0 13 9 13 9 0 13 2 13 16 13 9 13 2
9 16 9 9 3 13 0 1 15 2
16 1 15 13 16 9 9 3 13 13 15 15 13 1 15 0 2
21 3 3 13 15 1 15 9 13 2 16 9 13 9 2 1 15 13 0 13 0 2
20 15 7 13 15 2 13 15 15 15 1 15 13 2 16 13 9 13 9 9 2
22 16 3 0 13 15 15 13 1 15 16 13 13 2 0 13 15 13 15 15 15 13 2
12 7 3 0 13 15 13 15 15 13 0 0 2
2 3 2
24 16 1 13 4 2 9 2 13 10 9 2 15 13 10 9 2 13 10 15 16 13 15 9 2
28 1 15 7 16 15 13 9 9 16 3 2 3 13 1 15 13 9 0 9 2 3 0 2 15 13 9 13 2
13 3 13 3 9 13 15 15 13 9 9 16 3 2
26 16 7 9 9 16 13 9 13 13 0 2 3 9 9 16 3 13 16 15 13 3 9 7 3 9 2
13 3 13 3 9 13 16 9 7 9 13 3 0 2
18 15 7 13 1 10 1 15 0 2 15 1 15 9 13 16 9 13 2
10 9 3 9 3 13 13 1 15 0 2
2 0 2
8 9 3 13 16 15 9 13 2
14 15 3 15 3 13 1 9 2 3 13 13 1 9 2
33 7 15 15 13 1 15 0 3 13 1 9 2 1 15 15 13 2 16 9 1 9 3 13 9 9 2 15 1 9 13 3 13 2
13 1 0 3 9 3 13 13 15 1 15 13 0 2
2 3 2
14 1 16 15 15 13 1 9 2 3 15 13 1 9 2
8 7 0 13 15 3 13 13 2
6 3 3 13 13 0 2
18 3 7 13 1 9 2 15 3 13 16 15 15 13 7 13 13 0 2
15 16 0 9 3 13 9 1 9 2 7 15 9 0 13 2
18 1 13 7 13 13 16 0 9 9 3 13 2 7 9 0 9 13 2
15 13 3 9 10 15 13 1 9 15 13 2 16 13 4 2
15 7 15 9 1 9 10 9 13 16 13 13 2 3 0 2
7 3 13 15 9 13 13 2
26 9 7 0 9 13 16 3 0 13 15 9 13 13 2 7 3 16 15 9 13 16 9 13 15 13 2
35 3 7 1 9 0 2 1 9 13 13 0 2 13 15 10 9 3 0 3 1 9 2 7 3 3 1 9 2 15 13 15 9 15 9 2
8 3 9 0 9 9 3 13 2
2 0 2
21 9 0 13 9 9 10 9 16 15 9 0 2 3 1 15 0 13 10 9 9 2
9 9 7 0 13 16 13 15 13 2
9 15 3 10 9 9 1 0 13 2
7 13 3 9 15 13 13 2
2 3 2
13 9 0 1 15 9 13 2 16 13 1 12 0 2
22 13 7 9 0 15 9 13 0 2 1 9 13 1 9 0 2 15 3 13 16 13 2
8 1 9 7 0 9 13 13 2
11 3 3 13 13 9 0 9 16 10 9 2
52 3 13 2 16 9 13 13 0 2 16 3 9 0 13 13 2 9 13 13 2 16 13 1 15 15 1 9 9 13 2 15 3 13 13 1 0 9 9 2 16 9 13 2 15 13 9 0 2 13 1 9 2
7 13 3 9 15 13 13 2
2 3 2
13 9 1 9 1 9 3 13 13 9 0 1 9 2
23 9 7 13 15 1 9 3 9 0 2 7 0 9 15 13 1 9 2 16 1 13 4 2
13 1 9 3 0 3 13 13 1 9 13 9 0 2
6 15 7 0 13 9 2
20 3 3 13 1 15 13 1 9 0 2 16 9 13 2 16 13 2 13 0 2
10 0 3 9 3 13 1 9 13 9 2
32 3 3 13 2 16 9 13 15 2 16 15 1 9 13 2 7 16 15 0 13 0 7 0 2 16 9 15 13 2 15 13 2
7 13 3 3 13 13 0 2
7 16 0 9 13 9 13 2
12 13 7 1 13 13 16 0 9 9 13 13 2
11 9 3 13 9 13 15 15 13 1 9 2
19 9 7 13 9 10 16 9 2 10 7 15 13 16 15 15 13 1 9 2
14 10 3 9 13 9 3 13 15 15 13 0 1 15 2
2 3 2
15 9 0 13 1 9 15 16 1 9 2 16 0 1 9 2
15 3 7 13 15 1 0 9 1 16 15 13 1 9 9 2
16 13 3 16 9 0 13 9 3 9 13 15 0 9 1 0 2
2 3 2
22 16 1 13 4 2 13 16 9 15 13 2 13 1 9 16 13 15 15 1 15 13 2
12 15 7 15 9 13 2 13 9 3 15 13 2
19 9 3 3 9 13 15 15 13 1 15 2 13 16 13 15 1 15 13 2
10 3 3 13 13 1 13 0 9 9 2
32 9 13 9 13 9 1 15 16 9 13 2 13 7 9 13 1 15 16 9 0 13 2 13 7 9 0 13 16 13 9 15 2
10 3 3 13 0 9 1 15 9 13 2
16 3 9 0 7 13 1 9 0 2 7 1 15 15 15 13 2
52 9 7 0 2 16 1 15 0 9 1 9 13 2 15 13 0 9 0 2 1 15 3 3 13 1 9 2 7 3 1 15 15 9 7 9 13 0 2 16 1 15 15 13 0 1 9 7 9 15 9 0 2
26 0 7 9 13 1 9 1 15 15 1 15 0 13 2 16 7 15 3 13 15 15 13 1 0 15 2
29 3 3 9 0 9 13 0 9 2 3 9 2 3 7 9 15 13 1 9 2 9 0 0 2 0 1 13 15 2
8 16 0 9 15 13 13 9 2
19 16 7 15 9 0 9 13 13 2 3 3 13 16 9 15 13 15 9 2
7 9 3 9 13 13 9 2
8 9 7 0 9 13 10 9 2
14 15 3 13 9 9 13 2 15 13 3 15 10 13 2
11 15 7 1 9 13 15 13 9 9 13 2
13 7 12 15 13 15 9 16 9 13 1 0 9 2
10 7 3 13 9 1 12 15 15 13 2
12 13 3 16 3 13 9 15 13 1 9 9 2
17 3 16 13 12 9 2 3 13 9 2 16 1 1 9 13 4 2
19 9 7 12 9 13 7 10 9 7 10 15 2 1 10 9 13 10 9 2
26 1 13 7 13 9 15 13 10 13 1 9 1 0 9 2 16 1 15 13 9 13 16 16 9 13 2
16 15 3 9 0 13 2 15 9 13 1 9 9 10 10 13 2
4 1 15 9 2
5 10 1 9 13 2
14 7 8 12 13 16 9 13 9 10 1 10 9 10 2
7 16 1 9 13 0 9 2
12 1 13 7 13 13 16 1 9 0 9 13 2
16 3 0 9 13 9 15 15 3 9 15 13 2 7 0 9 2
14 3 1 15 13 0 9 9 15 16 13 13 7 13 2
15 9 7 15 1 15 3 1 9 13 2 16 1 13 4 2
7 9 3 0 9 13 13 2
2 3 2
23 9 0 1 15 1 15 1 10 9 3 13 2 13 3 1 10 9 2 16 1 13 4 2
24 7 1 15 9 13 1 10 9 0 9 13 16 1 13 9 9 13 2 3 9 9 16 0 2
7 3 1 9 13 0 9 2
2 3 2
19 1 9 2 1 12 8 2 9 13 9 2 9 7 15 15 1 9 13 2
29 1 3 9 15 16 9 13 2 15 0 16 15 1 9 13 2 13 16 9 15 13 9 3 2 9 7 15 9 2
8 9 7 3 1 0 9 13 2
6 9 3 0 9 13 2
2 3 2
13 9 1 15 16 13 0 9 2 13 10 9 9 2
14 15 7 0 13 0 9 2 15 9 1 15 3 13 2
7 15 3 9 0 9 13 2
9 15 3 1 15 9 9 13 13 2
15 3 0 13 15 15 9 13 2 1 9 2 1 9 0 2
13 15 7 15 3 13 16 0 9 2 15 9 13 2
8 16 1 9 3 13 9 9 2
13 1 13 7 13 13 16 9 9 1 9 3 13 2
20 1 3 0 9 3 13 15 9 2 7 0 1 0 2 16 13 1 12 9 2
22 15 7 15 9 1 9 13 13 2 1 13 15 0 9 2 16 1 1 13 4 0 2
10 13 3 16 1 9 3 13 0 9 2
2 3 2
21 10 0 9 1 15 9 0 13 2 13 1 9 7 9 9 2 7 1 15 3 2
23 15 15 1 9 0 13 13 2 15 16 3 13 9 7 9 1 9 2 16 1 13 4 2
8 3 13 3 1 15 0 9 2
2 3 2
30 1 10 0 9 13 0 13 1 10 0 2 0 7 0 9 2 15 9 13 16 3 9 2 16 13 2 9 13 9 2
22 7 3 13 0 9 1 10 0 9 0 13 2 1 13 3 0 2 16 1 13 4 2
11 13 3 16 1 9 3 9 13 3 13 2
2 0 2
18 10 9 15 13 1 9 2 13 1 12 13 2 1 9 7 9 9 2
22 9 3 9 13 1 15 12 2 16 7 9 2 7 1 15 9 13 15 13 7 13 2
26 0 7 9 3 13 1 15 1 12 1 15 15 13 4 2 16 1 9 10 9 2 16 1 13 4 2
10 3 13 3 1 15 9 1 9 15 2
2 3 2
7 10 9 13 15 9 13 2
13 9 7 13 3 0 1 9 2 1 13 0 9 2
15 13 3 9 3 2 7 15 9 15 9 1 15 9 13 2
10 3 3 10 9 9 9 1 9 13 2
17 15 7 9 13 1 9 3 0 9 10 9 2 7 3 9 9 2
8 10 3 9 1 9 9 13 2
19 15 3 9 3 13 9 0 2 15 9 1 9 13 3 1 9 0 9 2
7 15 7 13 9 7 9 2
17 3 15 9 13 9 3 13 2 16 9 9 13 9 0 7 13 2
14 9 3 7 9 1 15 15 9 1 9 13 3 13 2
2 3 2
25 9 9 15 9 3 0 13 1 9 7 9 2 7 3 1 15 16 0 15 15 13 1 15 15 2
7 3 3 9 7 9 13 2
31 16 3 9 15 15 13 1 9 15 1 9 9 13 2 9 3 13 2 7 15 9 9 13 13 2 3 1 9 0 9 2
17 9 7 2 16 13 9 9 2 3 3 9 3 13 2 7 13 2
21 15 3 9 3 13 13 2 9 10 9 2 15 15 13 16 15 9 13 3 13 2
13 9 3 1 9 13 3 13 2 3 9 10 9 2
8 7 0 7 9 15 3 13 2
2 0 2
24 16 0 9 13 9 9 15 9 13 1 9 2 3 3 2 7 0 0 2 13 9 1 9 2
13 9 7 13 9 15 13 13 2 16 9 9 13 2
28 0 3 9 10 9 9 1 9 13 2 7 16 3 13 16 13 1 9 2 7 16 13 9 9 15 13 13 2
2 3 2
5 9 9 9 13 2
21 3 7 9 9 9 13 2 3 0 16 9 9 13 2 7 3 16 9 9 13 2
2 3 2
16 1 9 0 9 13 3 13 16 15 15 13 0 13 16 0 2
22 7 13 16 1 0 9 16 15 9 13 9 13 15 2 1 15 9 12 13 9 15 2
15 0 7 9 1 15 0 9 15 13 2 7 1 15 13 2
13 9 7 13 0 9 2 15 9 13 10 13 0 2
8 15 3 9 15 13 13 9 2
31 7 13 13 16 15 15 13 0 0 7 3 13 15 0 2 13 16 9 2 16 10 9 13 1 9 2 16 1 13 4 2
39 9 3 1 9 0 13 13 2 3 1 10 9 9 2 3 0 16 9 9 9 13 2 7 3 16 13 1 9 15 2 7 3 13 9 15 16 9 15 2
2 3 2
10 15 9 13 13 1 9 7 13 9 2
10 3 0 13 1 15 16 9 13 9 2
10 0 0 13 1 15 16 9 13 9 2
9 9 7 13 9 9 15 1 9 2
31 9 3 1 9 0 13 1 9 10 9 2 3 0 16 9 9 13 2 7 3 3 13 9 9 1 9 1 0 13 13 2
19 3 2 15 15 9 15 9 13 7 1 15 13 2 0 9 1 9 13 2
13 16 1 9 13 9 7 9 3 3 13 0 9 2
25 13 7 15 9 15 2 16 9 3 13 1 16 9 2 15 3 1 9 10 9 13 13 0 9 2
7 15 7 13 9 7 9 2
6 13 3 9 0 9 2
31 7 3 9 9 2 15 13 9 2 7 9 9 15 13 1 9 2 15 4 9 13 2 9 1 10 9 9 0 9 13 2
14 1 15 7 0 13 16 9 7 9 0 1 9 13 2
16 16 3 9 7 9 13 13 9 9 0 2 3 7 9 0 2
54 15 3 13 13 9 7 13 9 2 7 1 9 7 1 9 2 16 16 9 0 9 13 0 16 0 2 16 0 9 13 9 7 9 0 2 9 7 0 9 7 9 1 9 2 16 3 7 9 9 13 0 16 9 2
8 7 9 9 9 1 9 13 2
43 13 3 1 9 0 2 15 13 9 2 0 9 1 9 9 9 9 0 2 1 15 13 16 1 9 0 13 9 2 1 9 15 1 9 0 2 1 0 7 13 9 0 2
25 16 3 1 9 9 2 15 13 1 9 0 2 13 15 9 0 2 3 1 9 0 9 15 13 2
31 1 3 9 7 9 9 3 13 1 10 9 2 7 0 16 9 13 2 1 9 7 13 1 10 9 2 3 7 16 9 2
8 13 16 3 0 9 3 13 2
2 3 2
11 9 7 9 13 15 9 9 1 10 13 2
21 9 7 1 15 2 15 13 10 0 13 2 0 13 2 3 1 15 10 9 13 2
12 15 3 1 10 9 1 15 0 13 7 13 2
2 3 2
14 9 13 15 9 9 2 16 13 1 9 2 12 8 2
7 13 3 9 16 9 9 2
13 7 9 9 9 13 1 13 2 16 1 13 13 2
18 16 3 10 13 2 1 10 9 2 13 0 2 0 13 13 15 0 2
2 0 2
35 15 0 1 10 0 13 2 3 1 13 2 16 1 9 2 16 13 0 0 9 2 16 9 1 3 13 2 1 15 16 12 13 9 15 2
22 10 7 9 13 0 9 9 2 16 1 1 13 13 2 7 1 15 9 15 15 13 2
9 13 3 16 9 1 10 9 13 2
9 13 3 1 15 0 9 7 9 2
7 13 7 9 7 9 9 2
25 3 9 13 1 9 0 13 2 9 7 15 3 13 2 7 0 9 9 1 13 13 1 9 9 2
17 3 9 13 0 1 13 9 2 16 0 13 2 9 7 1 0 2
19 1 15 13 16 9 0 1 15 13 2 13 7 7 1 15 7 1 15 2
6 16 1 9 13 9 2
13 0 7 13 7 9 1 9 13 1 9 9 15 2
14 15 3 13 0 1 9 9 2 16 13 9 13 13 2
13 9 7 13 9 10 7 15 2 16 1 13 13 2
10 1 15 3 9 7 15 7 15 13 2
2 3 2
12 1 9 9 13 16 9 15 13 16 13 15 2
46 15 3 9 15 13 0 16 1 15 9 13 2 1 9 13 2 16 15 13 9 13 16 15 13 2 7 9 16 15 13 0 7 0 2 1 9 13 9 7 9 2 1 15 7 15 2
10 7 9 13 9 15 1 16 13 15 2
19 13 3 15 13 1 16 1 15 0 13 2 16 3 12 13 1 9 15 2
9 9 3 0 13 7 15 7 15 2
2 0 2
43 1 15 0 13 7 13 10 9 0 9 2 16 15 13 9 9 16 13 13 7 13 9 13 2 13 13 16 13 1 13 15 13 16 1 15 15 13 1 15 15 9 12 2
23 1 15 13 0 9 9 13 1 15 16 9 12 13 1 15 16 1 12 1 15 15 9 2
11 1 15 13 1 9 16 9 13 0 9 2
17 3 3 15 3 13 13 12 1 13 13 0 2 3 13 9 13 2
27 3 3 13 15 15 13 9 9 2 7 9 9 2 7 15 3 2 16 15 15 0 15 13 0 9 9 2
19 7 3 2 3 15 1 15 13 13 13 3 0 13 2 3 9 13 0 2
26 3 3 9 15 13 1 15 9 2 13 13 9 15 13 1 0 9 7 1 15 9 2 7 0 13 2
27 15 7 3 10 9 13 2 3 15 9 2 15 10 13 2 13 0 7 0 9 2 1 15 13 10 9 2
15 13 3 1 9 9 3 0 0 2 7 3 9 7 0 2
2 3 2
14 9 1 9 9 3 13 15 13 9 2 1 13 9 2
8 7 1 9 15 13 1 9 2
22 3 9 13 15 9 3 0 1 13 2 7 3 2 16 9 15 13 15 0 1 13 2
38 3 7 9 1 9 1 9 0 1 9 9 13 2 3 7 0 1 9 13 2 16 16 1 13 13 15 15 13 9 2 3 3 0 13 16 13 2 2
11 3 3 9 13 0 9 1 9 10 9 2
5 13 3 1 9 2
2 3 2
10 9 13 1 13 13 2 16 9 13 2
38 1 3 2 1 9 7 9 13 7 13 2 9 13 13 3 13 13 2 13 9 1 9 13 2 16 3 13 15 3 13 4 1 9 2 13 1 9 2
13 3 7 9 0 13 0 9 7 0 7 9 13 2
8 9 7 13 10 15 1 13 2
18 16 3 13 15 9 7 15 9 2 13 15 15 1 9 15 0 13 2
8 9 3 7 15 7 15 13 2
2 3 2
6 10 9 9 13 9 2
31 9 3 7 9 3 13 16 13 9 2 9 7 9 3 13 16 1 9 15 13 9 13 2 1 15 7 10 15 9 13 2
13 7 1 9 13 9 7 9 2 16 1 13 4 2
6 3 1 9 13 9 2
13 13 7 15 13 16 9 3 3 15 16 15 13 2
22 16 3 9 7 9 9 0 0 13 2 9 13 3 13 2 1 15 10 9 3 13 2
2 3 2
18 15 15 15 1 9 1 9 9 13 2 1 3 7 0 1 15 13 2
16 7 3 3 15 15 13 2 7 3 1 15 16 1 15 13 2
22 13 3 16 2 1 15 9 9 13 1 12 0 9 2 0 9 1 12 9 13 13 2
16 1 15 3 16 13 7 13 2 1 15 9 0 15 13 13 2
19 9 0 15 15 13 2 15 3 13 13 15 15 9 13 2 1 9 13 2
37 3 7 15 15 13 2 0 3 7 0 13 13 2 3 7 13 2 7 0 15 15 2 15 15 13 2 7 1 15 15 1 9 7 0 13 13 2
13 15 3 9 1 0 9 9 1 3 7 0 13 2
7 15 1 9 13 3 13 2
19 3 9 9 1 9 15 13 13 2 10 7 0 9 12 7 15 9 13 2
10 9 7 1 3 7 0 0 13 13 2
21 12 3 9 2 1 9 15 15 13 2 1 16 15 3 13 13 15 13 0 9 2
19 15 9 1 9 9 2 1 16 13 15 13 15 2 0 9 2 0 13 2
22 0 3 3 9 2 15 13 13 16 9 15 15 3 13 2 1 16 15 0 13 9 2
15 0 7 9 13 3 13 2 15 9 15 1 15 13 4 2
37 13 3 1 13 16 1 10 9 15 13 15 1 9 0 13 13 16 9 7 9 2 2 16 15 3 1 15 3 1 9 2 16 1 15 2 13 2
13 15 7 1 9 13 9 7 9 2 9 9 13 2
5 13 3 1 9 2
8 9 1 0 10 1 1 9 2
22 8 12 2 13 0 9 13 1 15 2 13 0 9 2 15 9 13 2 16 13 4 2
13 8 12 2 9 13 1 9 1 12 9 9 13 2
17 9 3 13 2 1 12 8 2 16 9 3 13 12 7 0 9 2
9 9 3 9 9 13 2 8 12 2
3 13 9 2
7 8 12 2 9 0 13 2
9 8 12 2 15 3 9 13 15 2
9 9 3 15 13 9 9 9 9 2
22 15 13 9 9 2 12 8 1 8 8 2 13 16 0 9 3 13 15 1 9 13 2
42 13 3 3 15 9 2 15 1 9 10 0 9 13 2 1 0 9 1 9 13 2 3 3 0 2 16 13 4 2 7 0 2 1 9 7 9 2 7 15 9 13 2
22 13 7 9 2 16 3 9 1 9 9 1 15 9 13 1 15 15 1 9 0 13 2
12 9 3 1 9 13 2 16 7 13 1 9 2
15 13 3 3 9 13 2 16 1 9 10 9 15 13 13 2
4 1 15 9 2
7 1 13 1 0 9 15 2
20 0 0 13 16 1 10 9 9 9 13 2 16 7 15 1 9 9 13 15 2
4 3 1 9 2
10 9 7 0 9 2 13 7 0 0 2
31 13 3 3 13 2 16 1 0 7 0 9 10 9 13 15 0 13 2 7 13 15 0 13 2 16 7 9 13 13 13 2
9 3 8 12 2 13 15 13 9 2
17 16 7 15 0 13 3 13 2 13 1 15 16 13 12 8 12 2
10 9 1 9 3 13 2 7 9 13 2
7 13 7 1 9 9 13 2
16 3 9 7 9 2 15 1 9 0 13 2 9 13 10 9 2
7 9 3 1 9 9 13 2
6 9 0 1 9 9 2
10 3 3 13 13 13 2 3 9 13 2
29 13 3 9 13 2 16 13 15 0 15 15 15 13 7 13 2 16 7 1 15 13 9 1 15 15 15 13 13 2
20 7 15 13 9 12 13 9 2 7 9 13 1 9 15 2 16 3 13 9 2
17 7 13 16 3 13 9 2 7 13 4 2 16 3 13 15 13 2
34 1 13 7 13 9 15 0 13 9 9 2 9 2 9 2 7 10 3 9 2 1 9 2 3 13 15 1 9 0 0 7 0 13 2
7 3 1 9 13 13 9 2
12 13 13 7 13 13 3 9 1 9 13 13 2
29 13 3 2 16 9 15 13 0 9 2 10 9 9 1 15 3 13 2 3 7 9 15 10 9 1 15 3 13 2
7 9 7 13 9 15 0 2
11 3 1 15 13 0 2 7 9 15 0 2
10 13 3 9 0 10 9 10 9 13 2
13 3 15 15 1 9 1 9 13 2 16 1 15 2
22 9 3 3 13 0 13 1 15 15 15 13 2 7 1 9 10 2 1 13 3 0 2
20 7 3 1 15 10 9 13 13 2 1 10 9 13 10 9 2 16 13 4 2
12 3 13 3 9 15 15 9 2 7 10 9 2
2 3 2
12 9 0 9 13 2 3 0 1 9 7 9 2
7 3 7 13 9 13 13 2
7 1 9 7 13 9 9 2
23 9 3 1 15 3 13 16 9 2 16 9 2 7 16 13 2 15 13 9 0 7 9 2
2 3 2
6 9 9 15 0 13 2
13 1 9 7 15 13 1 9 2 7 0 1 9 2
8 1 15 3 9 13 3 13 2
2 3 2
6 9 1 9 9 13 2
12 15 1 9 3 3 13 2 16 1 13 4 2
15 3 7 9 15 1 9 1 9 13 2 7 0 1 9 2
38 1 7 9 0 13 15 0 9 13 2 0 7 9 13 0 2 0 7 0 2 15 3 1 0 9 9 13 2 16 15 9 13 2 9 13 3 13 2
10 9 3 0 9 1 9 0 9 13 2
12 3 7 9 9 0 13 15 15 9 0 13 2
7 3 7 9 13 3 13 2
9 3 7 3 9 16 15 9 13 2
2 3 2
9 3 9 9 9 1 0 9 13 2
13 3 15 15 0 9 3 13 2 13 3 0 13 2
18 0 3 0 9 13 13 2 15 9 7 9 0 13 1 9 0 9 2
15 15 3 9 15 1 0 9 13 2 15 1 9 15 13 2
7 15 1 9 13 3 13 2
17 9 3 15 1 9 13 2 1 15 9 9 13 16 1 0 9 2
19 3 7 9 1 9 13 16 15 1 9 13 2 15 0 1 9 7 9 2
11 1 9 7 9 3 13 2 16 13 4 2
9 3 7 3 9 1 9 13 13 2
2 3 2
27 3 9 3 1 9 0 9 13 2 7 1 9 0 2 1 15 0 9 13 13 2 16 13 1 12 9 2
12 1 9 7 3 13 0 9 2 7 0 9 2
16 13 3 16 1 9 3 9 13 3 13 2 3 1 0 9 2
30 9 7 1 15 9 13 2 15 13 1 9 9 1 15 0 9 15 13 0 1 9 2 16 13 9 7 9 7 0 2
14 1 15 9 13 9 2 9 2 7 0 9 7 9 2
45 3 2 16 0 9 3 1 9 13 13 2 9 13 7 0 9 13 2 1 1 9 13 2 7 3 0 1 9 13 1 9 2 16 7 13 13 9 15 1 9 1 9 15 9 2
26 15 0 9 13 1 9 9 1 15 0 9 2 16 13 9 2 9 2 9 2 9 2 7 15 3 2
20 1 15 9 2 9 7 3 9 13 9 2 9 2 9 2 7 15 3 9 2
15 15 3 1 9 0 13 3 13 2 15 16 1 9 13 2
12 13 3 1 9 0 1 9 2 1 9 9 2
7 16 13 15 12 8 12 2
7 3 13 0 16 9 10 2
4 7 8 12 2
6 13 0 2 13 0 2
11 16 1 9 13 9 0 15 13 1 9 2
31 13 7 9 15 9 0 9 13 15 3 1 9 2 7 1 9 13 2 16 9 2 9 2 9 2 9 2 9 7 9 2
42 1 7 9 1 9 7 9 9 13 2 9 7 15 13 15 9 9 7 9 2 0 9 3 13 2 7 3 9 2 1 0 9 2 13 15 1 15 1 0 9 13 2
2 3 2
16 3 9 9 15 9 7 9 13 2 15 13 9 9 1 9 2
11 1 9 7 13 9 7 9 15 13 9 2
7 3 15 9 13 3 13 2
2 0 2
21 15 10 15 1 9 1 9 13 2 9 0 1 0 9 13 2 16 1 13 4 2
10 9 7 9 13 1 9 13 9 13 2
15 3 9 13 2 1 12 8 2 16 9 13 0 9 0 2
7 13 3 0 9 1 9 2
6 7 3 13 8 12 2
6 10 9 13 15 9 2
2 3 2
23 0 9 2 1 15 15 13 15 1 15 2 13 1 12 1 9 10 2 16 1 13 4 2
23 9 7 13 9 1 13 9 13 2 16 1 9 2 1 12 8 2 9 13 0 9 0 2
6 13 3 1 9 9 2
8 7 15 13 15 13 9 12 2
7 1 15 13 9 7 9 2
2 3 2
18 13 4 1 16 1 15 16 9 13 15 2 13 15 15 13 1 15 2
11 15 7 1 9 15 13 2 13 13 15 2
14 13 3 1 9 9 2 15 13 15 15 10 13 13 2
5 3 1 9 13 2
6 0 9 7 9 13 2
2 0 2
33 16 1 13 4 2 9 0 1 15 9 13 10 2 15 9 13 1 15 15 13 1 9 2 7 3 1 9 7 3 1 9 15 2
26 3 3 13 15 10 9 13 1 15 16 15 3 15 13 2 7 16 15 13 13 15 13 16 9 9 2
31 13 7 3 1 15 0 1 9 13 2 7 1 15 9 7 9 9 2 13 9 9 2 16 13 1 9 2 1 12 9 2
18 9 3 13 0 0 2 7 2 16 9 13 2 15 0 0 13 13 2
18 3 10 15 9 1 15 1 10 9 15 9 13 2 15 13 9 13 2
11 15 7 15 9 9 13 2 13 1 9 2
9 13 15 9 10 2 10 13 9 2
4 7 8 12 2
8 15 13 10 13 7 3 13 2
2 3 2
33 10 15 1 9 9 13 2 0 13 16 15 9 13 16 13 2 7 0 13 2 7 0 9 1 0 9 13 2 16 1 13 4 2
28 15 7 1 9 9 13 2 16 1 9 1 12 8 13 2 16 1 10 13 7 13 15 15 15 13 15 13 2
7 13 3 1 9 9 9 2
4 3 8 12 2
5 13 7 9 0 2
4 7 1 9 2
5 10 9 10 9 2
34 16 15 7 9 13 15 1 15 9 13 15 13 9 1 0 2 15 9 13 3 13 2 16 9 2 9 2 7 15 3 15 0 13 2
20 16 3 15 1 13 9 13 15 9 0 2 1 15 9 13 13 9 3 13 2
11 16 9 3 1 9 3 13 9 3 13 2
32 1 3 9 13 15 9 2 16 13 1 12 8 2 0 7 9 3 13 0 2 16 1 13 4 2 3 13 15 13 13 13 2
4 3 9 12 2
4 15 13 9 2
7 3 15 15 3 13 9 2
4 7 9 12 2
9 1 15 13 9 2 7 13 15 2
20 1 7 9 15 15 13 1 13 13 7 13 13 2 15 13 9 1 9 13 2
7 13 3 3 9 1 9 2
5 7 1 9 9 2
5 3 9 13 13 2
22 3 15 13 1 0 9 13 2 1 9 9 13 2 16 13 9 12 2 1 15 9 2
6 9 10 0 0 13 2
5 7 16 13 13 2
9 13 3 3 1 9 13 13 13 2
19 0 3 9 3 1 9 9 9 13 3 13 2 1 15 1 15 15 13 2
4 3 8 12 2
9 15 0 13 15 2 7 13 15 2
4 7 9 12 2
9 15 1 15 13 2 16 13 15 2
14 1 9 3 15 9 13 13 2 3 10 13 9 13 2
11 3 3 15 13 9 9 2 7 0 0 2
19 3 9 13 2 12 8 1 8 8 16 9 13 9 16 10 1 9 13 2
5 1 15 8 12 2
6 13 15 1 0 9 2
20 13 7 13 16 9 1 15 13 13 9 2 1 10 9 1 9 0 3 13 2
20 3 3 1 13 13 2 15 13 7 13 2 0 9 13 2 7 15 9 13 2
22 1 3 16 1 9 0 13 2 1 15 3 9 13 2 16 0 1 9 13 9 0 2
26 9 3 13 2 1 16 13 0 9 0 2 1 15 9 13 16 1 9 0 13 2 1 15 9 13 2
8 1 15 9 9 13 3 13 2
16 1 0 16 9 13 1 10 9 13 2 13 3 9 0 13 2
21 16 3 9 9 0 2 16 9 7 9 2 9 13 2 3 7 9 10 9 0 2
12 13 3 13 9 1 9 0 9 16 1 9 2
20 3 16 9 9 15 13 1 9 7 9 2 3 9 9 15 13 1 15 0 2
8 3 7 0 9 10 0 13 2
22 3 15 13 13 7 13 2 9 15 0 9 13 2 16 9 9 15 13 1 9 9 2
37 15 0 9 2 15 9 0 3 13 2 3 13 0 1 0 9 2 7 0 1 0 9 2 15 10 9 0 9 13 2 16 13 1 15 0 9 2
6 16 1 9 13 9 0
13 1 0 7 9 0 13 3 13 16 9 0 13 2
49 16 3 9 1 9 9 9 13 2 1 9 2 1 9 0 2 15 7 9 0 15 13 2 7 15 13 16 13 15 2 16 13 4 2 15 13 10 0 9 2 0 13 16 15 0 9 13 13 2
4 3 9 12 2
4 0 9 13 2
4 7 8 12 2
13 10 9 1 9 9 13 2 7 1 15 13 3 2
16 9 3 13 2 1 9 0 2 16 13 0 9 2 3 0 2
2 3 2
39 16 9 13 9 9 1 0 9 2 7 10 9 7 9 9 13 2 7 1 15 0 0 9 13 2 16 1 13 4 2 0 13 16 1 15 0 9 13 2
16 2 3 3 15 4 1 9 13 2 16 9 10 1 9 13 2
5 3 12 8 12 2
5 9 9 9 13 2
2 3 2
29 16 0 9 15 9 1 9 9 13 2 9 7 3 9 1 10 13 2 16 1 13 4 2 13 3 1 15 9 2
4 3 9 12 2
6 15 13 9 7 9 2
13 15 3 9 1 9 13 0 10 2 16 9 0 2
7 16 9 3 13 13 9 2
16 1 15 7 15 13 4 2 13 13 16 9 3 13 13 9 2
10 9 3 9 13 1 15 15 3 13 2
20 10 7 9 9 13 9 9 2 1 10 9 13 10 9 2 16 1 13 4 2
6 3 13 3 9 13 2
2 3 2
18 9 3 1 9 13 16 15 9 1 9 13 2 1 0 1 0 0 2
30 1 3 9 9 13 9 13 2 3 13 9 13 1 9 16 15 9 13 15 16 9 2 7 15 1 9 13 3 13 2
14 1 0 7 9 3 13 13 9 2 16 1 13 4 2
9 3 3 9 15 13 1 9 13 2
2 0 2
10 9 13 0 9 2 16 1 13 4 2
16 0 7 9 3 13 15 9 9 2 16 7 0 0 9 0 2
9 0 3 9 3 13 13 1 9 2
2 3 2
18 1 9 13 9 9 2 9 3 13 13 1 9 16 1 9 1 9 2
21 9 7 0 1 9 13 3 13 2 1 15 13 13 16 13 15 2 16 13 4 2
6 3 13 3 13 9 2
14 7 3 13 16 0 9 1 15 0 13 4 1 9 2
8 15 7 13 15 13 8 12 2
6 9 0 7 1 9 2
4 7 8 12 2
14 0 13 9 10 2 9 2 7 13 1 9 3 13 2
30 1 15 7 13 9 0 2 15 1 9 13 9 3 13 7 1 9 13 2 7 0 2 15 13 9 1 0 9 13 2
13 16 9 15 13 2 7 9 15 9 15 13 13 2
13 1 15 7 13 16 9 15 9 9 13 3 13 2
15 16 3 9 15 13 1 9 2 3 9 15 13 1 9 2
8 3 15 15 13 2 9 13 2
7 15 0 15 13 2 0 2
23 16 3 9 9 1 9 13 3 13 2 16 13 4 2 0 13 16 15 9 15 9 13 2
2 3 2
36 9 9 1 15 1 15 13 2 16 1 13 4 2 16 2 13 7 13 10 9 7 10 9 13 15 13 2 1 16 0 13 2 1 9 9 2
20 15 3 13 15 9 1 9 15 1 15 13 2 16 1 15 13 10 9 9 2
12 15 7 13 9 15 9 2 16 9 0 13 2
12 3 15 9 15 3 13 16 15 9 0 9 2
7 3 9 15 9 13 9 2
4 15 3 13 2
2 3 2
9 1 0 9 10 15 9 13 13 2
20 16 3 15 15 15 13 9 13 2 13 15 3 13 2 16 15 13 15 9 2
16 13 3 9 10 3 13 15 15 1 9 13 7 13 7 0 2
20 13 4 3 1 16 2 16 9 15 13 2 13 16 15 13 15 1 15 13 2
5 15 7 13 0 2
23 15 3 13 2 16 9 1 9 15 1 9 13 2 16 3 13 9 15 9 13 13 0 2
25 0 16 0 13 9 9 2 16 2 16 13 15 10 9 2 3 13 15 10 15 15 10 9 13 2
6 15 3 9 9 13 2
2 3 2
17 15 15 13 1 10 9 0 0 2 0 1 0 9 0 13 13 2
24 10 7 9 10 9 10 9 13 2 1 16 3 2 16 9 9 2 9 9 2 9 10 9 2
14 0 3 3 9 15 9 13 2 1 15 13 10 9 2
8 15 7 13 15 13 8 12 2
12 13 10 15 13 2 7 15 13 15 15 13 2
7 13 7 0 9 15 13 2
4 7 15 0 2
22 0 9 2 1 15 16 9 2 13 9 2 13 15 9 13 2 13 0 9 3 13 2
16 3 9 9 13 13 2 3 15 3 13 13 2 13 9 13 2
5 1 15 8 12 2
17 15 9 1 9 10 16 13 1 9 10 2 7 9 0 3 13 2
10 10 3 15 13 15 13 2 13 9 2
16 15 7 3 13 9 16 9 0 2 15 0 13 9 7 9 2
21 15 7 9 13 1 15 16 9 13 15 0 9 15 13 3 13 1 9 0 9 2
11 7 3 13 13 2 1 3 15 13 13 2
30 3 3 2 16 13 9 9 7 9 0 2 15 13 3 13 1 9 7 9 15 2 13 15 13 15 9 13 7 9 2
5 1 15 8 12 2
4 9 9 13 2
4 7 15 9 2
12 13 10 15 13 9 2 13 10 15 13 9 2
7 9 0 7 0 13 9 2
5 16 9 13 13 2
16 1 15 7 15 3 13 4 2 1 9 13 16 9 13 13 2
9 13 4 3 9 13 13 7 13 2
9 13 7 7 13 3 16 13 13 2
5 13 3 9 13 2
2 3 2
17 13 1 15 15 13 4 16 13 4 1 15 2 3 1 15 13 2
44 7 1 15 15 15 13 1 15 13 2 15 9 9 3 13 2 1 9 13 13 2 16 9 0 9 13 2 3 7 9 7 9 13 2 7 9 0 2 15 9 15 13 13 2
20 0 3 15 0 1 15 13 15 13 15 2 13 1 9 7 13 2 16 13 2
7 3 15 0 0 13 13 2
18 15 0 10 1 15 0 13 2 7 13 2 7 13 13 2 7 13 2
27 7 16 9 0 1 9 13 2 0 10 15 15 13 15 1 0 9 2 16 3 13 1 9 2 13 13 2
10 3 13 2 13 7 13 9 9 13 2
18 7 9 0 3 1 15 2 7 1 15 13 2 1 13 0 9 13 2
6 0 3 15 13 13 2
2 3 2
12 0 9 10 9 13 13 2 16 1 13 4 2
7 13 7 13 15 9 9 2
9 3 13 1 9 9 3 13 13 2
6 0 3 9 13 13 2
5 15 3 13 13 2
7 15 3 9 0 9 13 2
9 13 3 8 12 2 1 9 9 2
7 13 2 13 15 1 0 2
4 7 1 9 2
10 9 10 7 9 10 13 1 9 0 2
6 16 9 13 10 9 2
11 1 15 7 0 13 16 9 13 10 9 2
21 9 3 13 13 15 13 1 15 9 13 2 16 9 3 13 1 9 15 16 13 2
18 13 7 13 13 15 9 15 2 16 13 1 9 2 1 12 1 9 2
35 1 3 1 15 9 13 13 16 9 13 2 1 15 13 9 2 16 1 0 9 2 13 16 13 15 13 15 16 15 9 1 15 9 13 2
11 9 7 13 10 9 2 16 1 13 4 2
8 13 3 10 13 7 10 9 2
2 3 2
16 15 13 13 15 13 2 16 13 1 9 2 1 12 1 9 2
6 3 13 13 9 13 2
11 9 7 13 10 13 2 16 1 13 4 2
8 13 3 10 13 7 10 9 2
2 0 2
23 16 9 3 13 10 9 2 1 13 13 2 16 13 4 2 13 16 13 13 1 9 9 2
15 10 7 15 13 1 9 2 13 1 15 15 13 1 15 2
11 9 3 13 1 15 0 2 1 15 13 2
9 15 13 0 2 16 1 13 13 2
2 3 2
15 16 13 13 9 2 16 13 4 2 13 1 15 13 9 2
17 16 3 3 13 15 10 9 2 13 15 1 15 15 3 13 15 2
5 7 3 13 13 2
5 15 1 13 4 2
6 13 3 9 10 9 2
8 7 15 13 15 13 8 12 2
4 15 13 9 2
6 16 9 9 13 0 2
10 1 15 7 13 16 9 15 13 0 2
9 15 3 13 13 16 1 9 9 2
7 15 7 1 15 13 13 2
10 10 3 9 13 1 9 15 1 15 2
18 0 13 3 16 9 13 13 2 1 15 13 10 9 2 16 13 4 2
2 3 2
15 10 15 15 3 13 7 3 3 13 2 13 1 15 9 2
18 15 3 15 1 3 13 1 13 13 2 16 15 3 13 2 3 13 2
13 0 7 9 3 13 15 9 2 16 7 0 9 2
14 3 3 3 13 13 7 3 3 13 2 7 3 13 2
6 13 3 9 15 0 2
2 3 2
13 1 15 9 13 13 2 16 3 9 13 1 9 2
17 3 7 1 9 0 13 15 9 1 15 9 2 16 3 1 9 2
20 16 3 9 13 15 9 2 13 16 15 3 1 9 13 2 7 15 3 13 2
13 13 7 7 13 9 15 13 9 2 16 13 4 2
12 3 15 9 3 13 9 2 7 13 15 3 2
4 13 3 0 2
2 0 2
10 9 3 0 13 2 16 1 13 4 2
16 15 7 13 7 13 13 2 7 1 13 9 13 2 0 13 2
19 3 9 15 13 1 9 2 13 7 1 9 2 9 7 1 9 15 13 2
16 9 3 7 13 13 2 7 13 13 2 7 1 13 9 13 2
6 13 3 15 9 0 2
11 15 13 15 13 8 12 2 1 9 9 2
5 13 15 1 0 2
4 12 8 8 2
8 15 13 0 9 7 9 0 2
5 16 9 13 0 2
9 13 7 1 13 13 9 13 0 2
9 15 3 0 9 0 9 13 9 2
12 1 3 9 13 13 2 10 0 9 13 9 2
32 3 7 13 1 0 9 16 15 1 9 3 13 13 2 15 3 13 9 0 7 1 9 13 2 7 16 15 3 13 0 9 2
13 3 9 3 0 13 2 16 15 2 7 15 13 2
4 13 3 0 2
2 0 2
21 15 13 0 13 7 13 1 0 9 15 13 9 1 15 2 7 15 13 15 9 2
9 9 7 1 15 13 9 9 15 2
8 3 9 7 9 1 9 13 2
9 3 7 9 13 9 13 9 9 2
7 9 7 9 13 1 12 2
14 0 2 1 10 9 2 16 3 13 13 1 15 13 2
20 13 7 9 1 15 13 1 15 3 13 15 1 15 9 2 16 13 7 13 2
24 3 3 13 9 15 15 13 9 2 7 13 13 0 2 16 3 13 1 15 13 15 13 9 2
27 9 0 7 9 1 15 13 15 13 1 15 2 13 9 13 2 3 13 2 7 13 1 15 16 1 9 2
12 7 3 15 9 0 9 3 13 9 7 9 2
11 0 2 1 9 9 2 16 13 9 9 2
19 3 1 9 9 3 13 1 15 9 2 7 1 9 9 7 1 9 9 2
6 0 2 1 9 9 2
13 7 1 15 1 15 0 9 13 1 13 9 0 2
17 0 2 1 9 9 2 16 3 9 2 0 2 0 7 0 13 2
33 15 7 13 9 9 2 1 13 13 2 7 10 9 9 9 13 2 7 13 9 13 2 16 1 15 9 13 2 16 1 13 4 2
19 15 7 15 13 2 15 13 0 0 2 9 2 1 10 9 2 7 0 2
4 13 3 0 2
2 3 2
21 1 9 9 10 13 2 16 2 15 13 2 3 13 15 13 2 1 13 0 9 2
15 13 3 15 13 0 15 9 13 3 1 10 15 13 13 2
12 3 9 13 16 9 13 9 10 9 9 13 2
18 7 15 13 0 9 16 10 9 1 15 9 13 2 16 1 13 4 2
6 15 3 13 0 0 2
2 3 2
18 16 15 13 15 15 13 2 3 0 13 2 16 15 9 3 4 13 2
13 15 3 15 13 13 2 15 13 2 15 0 13 2
39 13 4 7 1 16 9 3 13 15 2 1 1 15 0 10 9 13 2 7 15 13 1 15 16 1 9 16 15 13 2 7 0 16 15 13 13 10 9 2
5 13 3 15 0 2
2 3 2
11 13 4 1 16 9 3 13 13 15 0 2
22 0 13 7 15 15 13 15 3 13 2 1 15 15 9 13 1 9 2 16 13 4 2
10 3 15 13 13 15 13 15 3 13 2
6 15 3 13 2 13 2
10 7 15 0 13 2 16 1 13 4 2
19 13 3 0 2 1 16 1 15 0 13 13 15 15 13 7 15 0 13 2
11 15 3 9 0 9 13 2 12 8 8 2
8 15 13 10 9 0 7 13 2
6 16 9 13 10 9 2
10 1 15 7 13 16 9 13 10 9 2
12 9 3 15 13 0 9 15 2 16 13 4 2
11 1 7 13 16 15 9 13 13 10 9 2
6 15 3 13 10 9 2
2 3 2
20 9 2 1 13 0 9 2 13 15 15 15 13 13 2 7 13 2 0 13 2
11 13 4 7 1 16 9 0 13 10 9 2
7 10 3 9 13 15 9 2
2 3 2
8 15 1 9 10 13 15 13 2
24 15 3 13 15 1 15 3 13 2 7 1 15 13 9 9 12 1 15 13 2 16 13 0 2
32 1 3 9 10 15 13 1 10 9 2 15 13 10 9 2 13 16 15 2 16 13 10 9 7 10 9 2 3 13 10 9 2
2 3 2
7 12 0 9 13 13 0 2
15 16 3 15 12 13 15 15 13 2 15 0 7 9 13 2
9 9 7 13 4 1 0 9 13 2
13 9 3 0 9 13 13 1 15 16 13 0 9 2
7 3 9 7 9 13 15 2
6 13 3 9 10 9 2
12 16 9 0 9 7 0 13 13 10 15 9 2
10 0 7 1 13 13 13 9 0 9 2
12 3 3 15 0 13 9 2 3 9 0 13 2
25 3 2 16 15 1 9 9 13 0 13 2 15 9 10 9 13 15 9 15 15 3 9 13 4 2
9 0 7 13 9 15 13 15 9 2
6 15 1 9 13 4 2
7 15 3 13 0 9 0 2
2 3 2
22 1 9 1 9 13 2 16 13 4 2 16 13 0 9 2 7 0 9 1 9 13 2
27 7 15 2 10 0 2 0 15 13 16 15 2 15 9 13 16 2 16 15 13 15 0 2 3 0 13 2
24 0 3 13 9 1 10 9 2 15 13 15 2 16 15 0 1 9 15 3 13 15 15 13 2
10 3 3 9 13 2 7 9 13 9 2
2 3 2
25 15 1 9 13 2 0 13 15 15 1 9 13 16 9 9 9 13 1 15 9 16 1 9 13 2
8 9 7 1 9 10 0 13 2
6 15 15 15 13 13 2
16 15 3 15 1 15 13 13 0 9 2 16 1 13 13 13 2
15 7 3 13 16 15 15 1 15 0 13 2 9 0 13 2
8 0 3 9 10 15 9 13 2
2 0 2
11 9 1 9 9 9 13 2 16 13 4 2
10 15 7 15 0 9 15 9 13 13 2
38 15 13 3 0 1 15 16 13 9 0 2 7 16 12 9 9 15 3 9 13 16 13 2 7 10 15 2 15 13 7 15 3 13 2 0 7 0 2
14 1 15 7 13 13 15 3 13 0 2 7 9 13 2
37 7 15 9 2 15 13 0 0 2 15 3 9 13 13 16 9 13 2 1 15 9 9 13 16 9 0 2 7 15 9 13 13 9 16 10 9 2
21 7 13 15 15 9 15 10 3 15 9 13 13 2 13 2 16 3 0 9 13 2
15 15 3 15 9 15 13 2 3 10 12 7 15 9 13 2
8 0 3 9 1 10 0 13 2
2 3 2
14 3 15 3 13 13 2 3 15 9 7 9 9 13 2
9 9 7 0 1 0 9 9 13 2
29 15 3 9 15 9 13 13 9 9 15 13 1 9 15 3 2 7 0 16 3 1 9 13 2 7 1 0 13 2
26 0 7 13 13 1 9 15 3 0 13 2 10 7 13 9 13 2 16 13 15 1 9 0 7 9 2
16 0 3 9 1 0 13 0 2 16 9 9 13 3 9 13 2
2 3 2
54 9 2 7 9 0 15 0 13 9 10 1 15 9 13 2 1 15 13 0 0 9 2 16 15 13 0 9 2 9 2 9 2 7 9 0 15 13 0 9 2 13 3 0 13 0 9 2 0 15 9 2 0 9 2
2 0 2
15 9 0 9 13 13 1 15 16 10 9 13 1 9 9 2
13 1 0 3 9 2 13 9 15 7 15 0 9 2
21 1 0 0 2 3 9 12 9 2 7 9 7 9 7 9 2 7 15 0 9 2
14 0 3 9 7 0 3 13 16 15 9 15 9 9 2
20 13 3 1 12 2 1 9 2 3 1 9 2 9 2 9 2 9 7 9 2
19 13 7 9 13 9 1 15 2 7 0 9 1 10 9 2 1 0 9 2
16 1 9 0 13 0 9 1 15 10 9 2 16 1 13 4 2
6 1 9 13 0 9 2
9 1 9 13 10 9 9 7 9 2
10 1 9 13 9 10 9 15 3 13 2
15 15 3 15 0 0 13 2 9 13 7 9 1 9 9 2
2 6 2
5 9 13 1 13 2
14 13 4 1 10 9 10 2 7 1 13 9 10 13 2
3 8 12 2
12 9 15 9 9 13 3 13 16 15 9 13 2
18 1 9 3 9 7 9 9 7 9 9 13 2 9 0 9 9 13 2
13 1 15 3 15 13 4 13 16 9 15 9 13 2
14 13 7 0 9 9 2 16 9 13 2 1 12 0 2
20 12 3 15 1 15 13 13 7 13 15 13 9 2 16 13 2 13 7 13 2
24 15 0 15 1 0 9 13 2 15 13 9 13 15 1 15 13 2 16 13 2 13 7 13 2
7 15 7 13 9 13 9 2
13 0 3 1 15 16 13 2 13 2 13 7 13 2
16 15 0 1 15 16 9 1 9 13 2 7 15 13 7 13 2
40 16 0 0 9 9 13 13 2 0 0 9 13 2 9 7 0 0 13 13 7 9 15 2 13 16 0 13 9 13 9 0 7 15 13 0 2 16 9 9 2
8 15 3 1 9 0 0 13 2
11 9 3 7 9 9 9 13 7 9 9 2
19 0 3 13 9 2 16 0 13 9 2 9 13 15 9 2 7 3 9 2
13 0 0 2 15 16 13 9 13 2 9 9 13 2
13 3 0 13 15 1 9 3 1 9 1 9 13 2
20 1 0 3 9 9 1 13 9 3 13 2 16 4 13 1 9 7 9 0 2
25 3 2 1 0 0 9 9 2 13 3 1 0 9 13 2 1 15 3 9 13 7 13 1 9 2
9 15 3 9 1 13 9 13 13 2
25 13 3 0 9 9 2 1 13 2 13 4 1 10 9 10 2 16 9 1 0 13 7 13 13 2
40 13 0 1 9 9 2 1 13 2 7 1 13 9 10 13 2 16 1 13 9 15 13 9 7 9 2 7 10 15 13 1 9 1 9 16 1 9 0 13 2
9 16 9 9 0 13 1 9 9 2
14 3 3 0 13 9 1 9 0 13 1 9 0 13 2
15 0 3 2 16 1 13 9 0 9 3 13 13 7 13 2
17 15 3 15 9 13 2 15 9 13 0 2 3 1 9 9 13 2
9 9 7 10 9 9 1 9 13 2
6 1 15 1 9 13 2
5 10 1 9 13 2
20 3 1 13 9 0 9 13 13 2 16 1 9 13 1 15 9 10 9 13 2
5 13 3 8 12 2
11 13 15 2 3 9 2 1 10 9 10 2
31 3 2 1 9 13 2 0 13 4 9 10 1 15 2 13 4 2 7 3 13 1 15 2 7 13 0 9 9 1 13 2
5 9 9 10 8 2
14 1 9 0 9 15 13 1 0 9 13 13 2 13 2
10 0 9 10 2 7 9 10 13 3 2
21 0 2 15 9 1 9 9 9 9 13 2 7 1 13 1 9 9 9 9 13 2
10 13 3 16 9 13 13 9 13 13 2
6 7 3 13 8 12 2
30 16 9 7 9 15 2 3 9 7 9 7 9 9 2 13 4 2 3 9 2 13 16 15 13 15 2 0 13 15 2
5 7 8 12 13 2
17 0 9 1 15 15 13 4 13 13 2 0 3 9 15 7 9 2
10 1 15 7 9 9 9 13 7 9 2
11 3 13 8 12 0 13 9 10 1 9 2
9 15 3 13 15 2 3 9 9 2
12 0 2 15 9 9 9 1 9 0 9 13 2
32 15 3 9 7 9 1 0 9 0 13 4 2 15 1 15 0 4 13 2 16 1 9 15 9 2 16 1 0 9 13 4 2
35 16 3 9 9 2 9 7 9 3 9 9 13 2 15 9 0 9 2 9 9 1 0 9 13 13 13 2 9 9 13 0 1 15 13 2
5 3 1 9 13 2
16 13 15 2 9 2 1 9 10 2 7 1 9 9 10 13 2
7 7 3 1 9 9 13 2
25 13 1 9 9 10 2 3 15 9 2 7 16 13 9 10 13 15 2 16 1 15 13 9 9 2
8 7 8 12 2 13 1 15 2
37 1 15 15 13 9 2 3 9 2 15 13 9 1 15 9 2 3 13 13 15 15 13 2 3 0 0 2 3 15 9 2 16 1 0 13 4 2
12 0 2 15 9 9 1 15 9 0 9 13 2
18 13 4 3 1 0 9 16 9 2 13 15 2 1 15 10 15 13 2
28 1 3 0 9 9 1 9 0 13 2 7 1 9 0 9 15 9 9 13 2 13 1 9 15 0 9 9 2
8 15 13 15 13 12 8 12 2
15 15 0 10 2 13 9 9 9 13 2 1 15 9 13 2
12 3 3 13 16 9 9 13 1 9 9 0 2
6 7 3 13 8 12 2
10 9 13 9 9 2 7 15 13 13 2
6 1 9 9 9 15 2
13 16 13 9 9 13 1 13 9 15 13 1 9 2
17 13 3 0 9 9 3 0 1 9 9 2 7 3 1 9 13 2
20 9 3 15 1 9 13 2 3 1 9 9 13 2 1 16 0 9 9 13 2
5 15 7 0 13 2
51 0 3 2 1 15 16 9 9 13 1 15 13 3 16 15 15 3 13 16 1 15 13 2 0 9 7 9 13 2 15 1 9 15 13 13 2 16 13 15 15 9 15 9 13 2 1 15 13 8 12 2
27 15 7 9 2 7 9 2 7 13 9 2 7 9 9 2 7 0 9 2 7 9 7 9 2 9 13 2
14 0 2 1 15 16 15 15 9 0 13 9 15 13 2
8 15 3 1 9 1 9 13 2
25 15 3 9 9 15 3 13 2 15 3 13 16 16 15 9 13 2 16 16 9 13 13 12 9 2
21 15 7 0 9 13 9 9 3 13 2 16 15 0 9 13 3 13 15 9 9 2
12 1 15 3 16 9 9 13 2 13 9 13 2
8 7 1 15 9 13 8 12 2
7 0 9 9 7 9 13 2
22 1 15 9 13 15 9 9 2 7 0 9 2 7 9 9 2 15 9 16 9 13 2
20 0 0 2 1 15 16 0 9 1 9 13 15 13 1 15 16 9 9 13 2
51 16 13 1 15 15 12 9 9 13 2 7 15 9 3 1 0 9 2 7 1 9 9 1 9 13 13 2 7 15 3 15 9 2 7 10 7 15 2 0 9 13 2 7 15 13 1 13 9 13 13 2
7 15 3 10 0 13 9 2
6 1 15 13 9 12 2
9 16 15 13 13 0 2 13 15 2
4 7 8 12 2
12 9 13 15 2 15 3 13 13 1 9 13 2
2 0 2
39 9 2 15 1 9 1 9 13 16 1 0 9 2 1 15 16 13 9 9 2 7 1 13 9 15 9 1 0 2 15 9 15 13 13 13 15 0 13 2
49 16 13 1 15 15 9 9 9 13 2 1 15 13 8 12 2 1 9 9 13 13 2 15 9 13 2 7 1 15 15 9 9 9 13 2 7 9 9 13 0 2 7 16 15 0 9 13 9 2
35 3 3 13 0 13 15 9 15 13 15 13 1 9 9 15 1 9 15 13 2 16 1 9 0 13 2 16 9 13 1 9 1 9 9 2
31 3 9 1 9 13 1 0 1 9 9 2 7 9 9 1 9 13 2 1 15 9 13 13 2 16 15 15 15 9 13 2
17 7 3 15 15 1 9 13 9 16 0 9 13 2 13 1 9 2
18 16 3 13 9 9 7 1 9 9 15 2 13 15 7 3 13 15 2
18 7 8 12 15 13 7 13 2 7 13 2 12 3 13 9 9 0 2
9 16 15 13 1 9 9 7 9 2
31 0 13 7 1 13 16 9 1 9 13 9 9 0 16 1 15 13 15 9 9 2 7 16 9 1 15 13 1 0 9 2
12 7 3 15 9 13 13 9 2 7 9 0 2
10 3 9 0 15 13 1 16 3 13 2
11 3 7 1 0 9 9 0 9 9 13 2
30 9 7 0 15 13 2 3 16 3 2 16 9 16 9 13 2 7 16 0 9 13 2 7 1 15 9 15 9 13 2
6 16 3 8 12 13 2
7 9 9 0 13 9 15 2
9 3 9 13 13 0 10 0 10 2
13 7 1 15 3 15 1 9 7 9 7 0 13 2
16 9 3 13 15 15 15 1 9 0 13 2 16 9 13 3 2
33 0 7 15 0 13 1 9 15 15 13 1 16 13 1 9 13 2 16 2 16 13 1 9 13 2 16 13 9 13 2 7 3 2
22 3 3 13 1 9 9 9 13 16 0 9 9 13 2 16 9 9 2 7 9 9 2
24 3 3 7 0 1 9 15 9 13 15 9 2 7 0 15 15 13 15 16 13 9 9 0 2
19 16 15 0 1 9 0 1 9 7 0 13 2 1 15 7 15 9 13 2
39 3 9 9 13 1 0 9 9 2 0 7 1 9 0 2 16 13 2 16 3 0 4 13 2 7 16 15 1 9 9 13 2 7 16 9 9 13 0 2
14 3 7 15 0 9 13 13 2 3 1 9 9 13 2
5 1 15 8 12 2
9 15 13 9 10 7 9 1 9 2
12 7 1 15 15 2 3 0 2 9 0 13 2
12 7 3 3 1 9 9 0 2 9 0 13 2
15 3 7 1 9 0 9 13 10 9 9 1 10 13 13 2
11 3 3 13 16 3 15 9 15 9 13 2
29 3 1 9 9 2 15 9 1 15 13 7 1 15 2 1 9 9 13 2 0 13 9 1 9 7 0 1 9 2
23 1 9 0 9 2 15 9 3 16 1 9 1 9 13 2 0 13 9 9 7 3 9 2
16 7 3 13 9 2 16 9 9 0 2 15 15 13 15 13 2
28 3 2 1 15 9 2 1 15 15 1 9 1 15 1 0 9 4 13 2 1 15 15 1 15 13 13 13 2
3 9 13 2
37 13 7 15 9 9 2 16 0 13 1 9 9 1 9 2 0 2 1 15 9 2 0 0 1 15 9 13 7 13 9 2 3 1 9 13 9 2
9 16 9 13 16 13 15 9 13 2
21 13 3 15 1 0 13 4 2 13 3 16 13 9 16 13 15 13 9 7 9 2
19 13 4 3 1 2 1 9 9 2 13 15 0 9 0 2 15 9 13 2
9 0 7 9 10 9 1 9 13 2
7 9 3 15 13 9 13 2
2 3 2
20 13 4 1 0 9 2 1 9 15 2 13 15 0 13 0 2 15 9 13 2
16 0 7 13 1 15 9 9 13 9 10 9 15 13 15 9 2
29 1 3 0 1 9 9 13 1 9 2 1 15 9 9 13 0 13 13 4 2 13 16 9 13 0 9 9 13 2
2 0 2
21 15 1 15 15 13 2 0 15 13 0 13 2 16 9 0 2 7 9 3 13 2
11 13 7 15 9 1 15 13 9 1 9 2
11 3 15 9 1 15 13 16 1 9 13 2
11 10 3 9 9 13 4 13 15 9 13 2
13 7 9 13 9 9 2 16 1 0 9 13 4 2
13 3 15 13 13 15 9 9 2 15 13 9 13 2
2 3 2
21 9 9 1 9 9 13 16 13 15 0 13 2 16 13 1 9 2 1 12 9 2
13 9 7 13 0 9 2 16 1 0 9 13 4 2
17 15 3 13 13 15 15 0 9 1 9 2 16 3 13 9 13 2
2 3 2
16 13 4 1 0 9 16 9 13 10 9 15 13 1 9 9 2
19 1 9 7 9 13 16 13 9 7 9 9 2 16 13 1 12 1 9 2
19 1 3 0 9 13 9 2 3 13 15 9 13 9 10 15 1 9 9 2
7 7 3 13 15 9 13 2
2 3 2
18 3 15 9 9 13 9 2 3 9 10 13 1 0 13 7 3 13 2
19 9 3 2 16 13 0 2 0 0 13 2 16 7 13 0 2 3 13 2
20 9 7 0 2 15 9 13 2 9 13 16 9 9 13 2 16 1 15 13 2
6 9 7 9 9 13 2
60 1 3 1 9 15 1 15 13 13 3 0 1 9 1 15 13 2 16 13 13 7 13 2 7 3 1 9 15 1 0 13 2 1 15 15 13 13 2 0 3 9 13 2 1 15 16 9 13 2 3 0 13 7 13 2 7 3 13 9 2
8 7 3 13 15 13 9 13 2
7 15 13 15 13 9 12 2
10 15 13 0 7 0 7 0 1 9 2
7 16 1 9 13 9 0 2
17 1 15 7 13 16 9 13 13 2 7 16 15 13 9 0 13 2
13 9 3 0 13 9 13 1 15 1 16 13 15 2
8 9 7 13 13 15 9 13 2
6 3 13 15 13 13 2
2 0 2
16 16 9 0 13 9 1 9 2 3 9 0 13 9 1 9 2
17 15 3 1 15 13 16 13 9 2 13 0 1 15 16 13 9 2
6 7 9 13 13 9 2
6 3 13 15 9 0 2
2 3 2
15 0 9 10 9 1 15 13 2 16 1 0 9 13 4 2
8 9 7 0 1 9 9 13 2
10 15 3 3 0 9 13 3 9 13 2
8 9 3 0 9 3 13 13 2
2 3 2
7 10 15 13 13 13 13 2
21 3 15 3 13 13 2 0 13 13 2 7 15 0 13 13 2 0 13 3 13 2
12 9 7 13 13 7 13 2 16 1 13 4 2
16 3 13 13 13 2 7 9 15 13 13 0 2 7 3 0 2
7 15 13 15 1 9 13 2
5 13 13 2 9 2
3 7 3 2
14 9 10 9 2 7 9 10 1 1 9 15 13 9 2
7 16 9 9 13 15 9 2
14 1 15 7 0 13 13 16 0 9 13 15 9 9 2
10 9 3 0 13 15 1 16 13 9 2
35 9 7 13 9 15 2 3 7 13 9 9 1 15 9 15 3 13 15 13 15 2 1 1 15 15 13 9 2 16 1 0 9 13 4 2
6 13 3 15 10 9 2
2 3 2
14 10 13 15 3 13 10 9 2 13 13 9 9 15 2
21 1 9 7 15 13 13 0 2 1 13 15 10 9 2 16 1 0 9 13 4 2
6 13 3 15 10 9 2
2 0 2
12 9 0 1 9 9 13 2 16 1 13 13 2
17 10 7 0 9 1 15 10 9 13 2 16 1 0 9 13 4 2
11 0 3 9 3 13 15 1 15 9 15 2
13 9 7 13 10 9 2 16 1 0 9 13 4 2
5 13 3 10 9 2
2 3 2
14 1 9 15 9 3 13 15 9 2 15 9 13 9 2
9 3 9 0 1 0 9 9 13 2
15 1 9 7 3 13 13 15 9 2 16 1 0 13 4 2
6 9 3 13 10 9 2
2 3 2
17 10 15 13 1 15 2 13 1 15 15 13 1 15 16 1 0 2
11 15 0 9 13 1 9 16 1 0 13 2
6 13 3 13 1 15 2
11 15 7 1 15 13 2 1 10 9 13 2
11 15 7 15 15 13 2 13 15 0 9 2
9 15 3 9 9 13 15 0 9 2
7 16 9 9 13 15 9 2
15 1 15 7 13 13 16 9 9 3 13 15 16 10 9 2
13 15 3 12 7 15 13 15 2 15 3 13 15 2
11 0 7 9 13 15 9 2 16 13 4 2
17 15 3 9 13 15 9 2 16 1 0 9 13 4 1 0 9 2
7 15 3 9 1 15 13 2
11 3 1 9 3 13 15 9 7 15 9 2
2 3 2
9 9 15 9 13 9 15 9 15 2
10 13 3 1 9 16 9 0 1 0 2
15 0 7 9 3 13 15 16 15 2 1 13 15 9 9 2
11 1 9 3 3 13 15 9 7 15 9 2
2 0 2
14 16 9 0 13 15 13 2 3 9 15 13 15 13 2
11 7 0 9 13 15 9 2 16 13 4 2
7 3 10 13 13 10 9 2
7 7 15 9 13 10 9 2
5 7 3 16 0 2
2 3 2
13 9 15 3 13 9 9 2 13 15 16 9 9 2
10 3 7 9 12 1 12 9 9 13 2
11 1 9 7 3 13 13 15 1 9 9 2
15 1 9 3 10 9 3 13 15 1 10 9 7 10 9 2
6 15 9 1 9 13 2
37 16 0 15 13 15 15 9 2 1 0 9 3 13 15 16 15 9 2 0 13 1 13 16 9 3 13 1 9 16 9 9 2 7 16 9 13 2
69 7 16 9 9 1 15 13 1 9 9 2 13 3 9 0 9 13 1 15 2 16 13 1 9 1 12 8 2 0 13 16 9 13 1 9 1 9 1 13 2 1 9 9 2 3 1 9 1 9 16 1 9 13 2 16 9 10 0 9 15 13 2 0 3 9 7 15 9 2
35 3 2 16 15 9 9 13 15 3 1 15 13 13 7 13 1 13 2 9 15 3 13 1 9 9 16 1 9 13 2 3 1 9 9 2
8 3 7 9 13 13 7 13 2
16 9 3 9 2 0 13 2 3 13 3 9 2 7 0 9 2
16 9 3 7 9 1 9 3 13 16 9 2 7 0 16 9 2
44 13 3 1 13 16 9 9 15 9 13 2 16 13 2 13 2 13 9 2 7 0 2 3 13 0 9 2 1 15 15 9 1 9 13 15 15 9 2 15 13 12 7 15 2
23 3 7 9 9 12 9 9 3 13 2 1 15 15 1 0 9 13 4 2 0 13 13 2
9 16 1 9 13 15 0 1 9 2
40 1 7 9 9 13 9 10 9 2 9 7 9 9 13 2 16 13 4 2 9 7 0 1 13 13 2 0 13 16 15 0 13 13 1 9 1 9 10 9 2
2 3 2
17 3 13 13 15 0 13 1 15 16 1 0 15 0 13 1 15 2
26 7 9 15 0 13 1 9 2 3 1 10 9 2 15 1 9 13 2 16 13 4 2 1 15 13 2
9 9 3 1 13 0 1 9 13 2
2 3 2
5 9 13 9 15 2
12 9 7 2 16 7 10 9 2 15 0 13 2
7 13 3 15 0 1 15 2
2 0 2
6 9 1 13 0 13 2
13 9 7 3 0 15 15 2 7 3 15 9 13 2
9 3 15 0 13 1 9 1 15 2
2 3 2
11 13 13 0 1 13 2 7 13 1 13 2
13 9 7 13 13 7 13 3 13 2 16 13 4 2
6 13 3 1 15 9 2
2 3 2
7 0 9 15 13 0 0 2
13 13 4 7 1 0 15 13 0 9 7 0 9 2
9 13 3 16 0 1 9 0 13 2
13 16 9 13 1 9 1 9 3 13 0 1 9 2
16 3 7 9 15 13 1 10 9 2 0 1 9 13 3 13 2
24 3 3 1 15 13 13 16 9 1 9 2 1 1 15 15 13 9 16 1 0 9 13 4 2
8 7 3 13 13 15 9 9 2
32 1 3 0 13 15 1 10 9 1 15 3 15 13 2 16 9 13 1 9 2 13 16 9 9 15 15 15 13 1 15 13 2
23 15 7 15 15 13 1 15 13 2 3 1 15 13 2 1 7 13 7 13 1 15 13 2
11 13 3 16 9 9 1 15 0 13 13 2
15 7 3 3 13 1 15 13 2 16 1 0 9 13 4 2
10 3 13 3 3 9 1 9 1 9 2
2 3 2
12 13 4 1 0 16 9 10 9 13 0 9 2
17 13 3 9 1 15 9 16 0 1 9 10 2 15 15 9 13 2
23 3 1 15 16 9 13 7 3 13 2 9 7 9 0 7 0 13 2 1 9 1 9 2
22 0 7 16 1 9 0 13 2 3 9 1 9 1 0 3 13 2 7 1 9 3 2
24 3 1 9 2 1 12 8 2 0 13 0 2 3 16 15 13 2 7 16 15 13 1 15 2
9 13 3 9 1 9 3 13 0 2
2 3 2
38 9 13 13 1 9 3 0 9 15 15 13 9 2 7 9 15 15 13 1 9 2 16 7 15 9 13 2 7 9 15 13 7 0 9 7 0 9 2
19 7 15 15 13 9 1 15 15 3 13 9 7 9 2 3 13 9 0 2
25 15 13 16 13 0 9 9 1 15 2 1 9 0 1 9 13 0 0 2 15 10 15 13 0 2
26 9 7 3 15 13 1 15 15 13 9 16 1 15 15 13 9 2 16 3 13 1 15 16 15 13 2
12 3 3 13 1 15 1 9 0 1 15 13 2
2 0 2
18 15 15 1 0 13 2 0 13 15 13 2 7 1 15 7 1 9 2
23 9 7 15 1 0 13 1 9 2 16 16 13 9 7 9 15 9 15 1 0 13 13 2
29 16 3 13 15 9 0 1 9 13 2 13 16 15 9 1 0 13 2 7 3 16 13 7 1 15 7 1 9 2
8 15 0 1 0 9 13 4 2
7 3 13 9 1 9 13 2
16 3 7 13 13 16 9 13 13 13 0 16 9 15 1 9 2
26 1 3 9 13 0 9 7 0 9 2 13 1 15 3 9 2 15 13 15 9 2 9 9 15 13 2
14 7 16 15 3 13 9 15 2 13 3 0 9 13 2
5 7 3 1 0 2
17 3 3 9 15 9 1 9 15 13 2 13 9 15 1 9 13 2
2 3 2
8 0 13 9 15 15 0 13 2
23 13 3 15 1 15 15 1 15 13 2 16 1 9 13 15 13 3 2 7 1 9 3 2
13 15 0 13 1 15 15 13 2 16 1 9 0 2
14 1 9 0 3 13 15 13 3 0 13 2 7 13 2
12 3 3 13 15 9 16 1 9 15 15 13 2
18 3 3 13 13 16 9 15 9 1 9 13 2 13 9 15 1 15 2
34 1 3 13 4 16 3 13 1 15 0 2 7 3 13 1 15 2 13 16 7 13 0 1 9 9 2 1 15 16 15 13 1 15 2
23 9 3 10 2 13 15 13 1 15 2 13 9 15 1 15 2 16 1 9 3 3 13 2
20 7 3 3 13 16 15 9 13 1 9 13 9 2 7 15 15 1 9 13 2
13 3 10 15 2 16 9 2 9 2 15 9 13 2
11 9 0 13 0 2 7 1 9 13 3 2
6 7 3 9 13 0 2
22 1 15 3 15 16 9 10 13 9 0 9 13 1 15 9 2 15 13 0 1 15 2
15 16 7 0 0 13 7 13 1 15 16 9 13 1 15 2
27 13 3 1 15 16 0 9 3 13 16 0 9 1 15 13 2 16 15 9 3 13 2 16 13 13 9 2
28 15 3 13 9 10 13 0 2 7 0 13 1 15 15 13 1 15 0 2 16 3 15 0 1 0 9 13 2
35 7 3 15 13 3 0 2 3 13 0 9 7 0 9 2 7 1 15 0 13 13 2 16 9 0 13 9 16 9 2 7 9 16 9 2
15 15 3 15 16 0 0 1 9 13 2 15 0 9 13 2
7 16 9 13 10 9 13 2
23 16 0 13 4 16 9 13 15 13 9 2 13 0 13 16 15 1 15 13 16 1 15 2
21 10 3 15 15 13 3 1 16 15 13 2 1 15 9 13 15 2 16 0 9 2
23 3 15 9 3 13 2 0 7 0 13 2 3 0 13 16 13 1 15 7 1 16 15 2
13 0 13 7 15 12 12 13 7 15 1 16 15 2
24 15 3 1 15 1 16 15 13 2 15 3 13 2 16 13 12 9 12 13 0 3 13 0 2
14 16 3 15 12 13 2 3 13 15 1 16 15 13 2
55 0 13 3 15 12 1 12 13 3 16 1 15 1 9 13 2 7 13 7 12 13 15 9 2 16 9 13 9 9 9 13 2 1 3 15 0 13 2 7 13 16 15 0 13 9 15 2 16 12 9 9 13 9 13 2
9 9 7 13 1 10 15 15 13 2
27 0 13 3 13 15 12 15 15 13 9 13 2 7 13 15 13 13 1 9 2 7 15 15 13 9 13 2
19 13 3 16 1 15 15 15 13 9 13 2 13 10 15 15 15 9 13 2
13 9 7 1 13 3 9 13 15 15 13 9 13 2
10 1 15 3 13 10 15 15 9 13 2
16 16 7 13 16 9 3 13 9 0 2 15 0 13 9 13 2
19 3 3 1 0 0 13 2 7 1 9 2 7 3 13 13 9 1 12 2
2 0 2
21 15 15 13 1 10 9 2 3 1 15 9 2 13 1 15 7 13 13 3 13 2
29 16 3 9 15 0 13 7 13 2 3 15 9 13 2 16 7 1 9 13 2 1 15 9 13 7 13 9 13 2
35 16 7 2 9 7 9 9 0 13 2 15 13 13 2 3 13 16 15 3 0 13 1 15 9 2 7 1 15 15 2 1 15 9 13 2
21 15 3 15 0 13 16 15 2 3 13 15 1 10 9 3 2 7 1 15 9 2
15 15 3 13 9 10 1 15 9 15 0 13 15 9 9 2
22 3 7 15 0 0 13 13 13 9 9 1 10 0 2 7 15 0 0 9 10 0 2
13 9 7 13 0 9 2 16 1 0 9 13 4 2
10 15 3 13 9 10 1 15 9 13 2
2 3 2
16 1 9 9 13 13 9 9 2 15 16 9 9 10 13 13 2
58 3 13 16 2 16 9 0 13 1 9 0 2 3 15 15 0 13 1 9 0 2 13 1 15 9 0 2 16 1 0 9 9 15 7 15 13 9 0 9 9 2 7 9 13 0 9 9 1 9 2 1 13 9 7 3 9 0 2
6 10 7 0 13 9 2
14 13 3 16 1 10 9 13 15 9 15 13 13 9 2
11 0 7 9 9 13 2 16 1 13 4 2
9 13 3 10 15 13 1 9 13 2
2 3 2
22 15 1 9 13 2 13 9 10 15 1 9 13 2 16 9 13 9 10 13 16 3 2
13 9 7 13 9 1 9 10 2 16 13 15 9 2
26 10 7 15 9 13 9 1 9 2 16 9 15 13 10 9 3 13 13 16 12 16 1 0 13 4 2
8 9 3 13 9 13 10 15 2
2 3 2
34 10 15 13 0 13 7 3 13 2 13 9 15 2 16 1 15 13 1 15 15 13 2 7 3 13 13 15 15 15 15 1 12 13 2
24 3 2 1 1 0 13 3 13 2 13 16 13 15 0 15 13 9 10 0 9 7 3 9 2
30 0 7 15 13 13 9 10 9 2 1 15 3 1 0 13 3 13 2 7 3 13 13 1 15 15 13 1 15 13 2
15 15 7 3 13 13 16 12 2 16 1 0 9 13 4 2
5 7 15 13 9 2
14 13 3 10 15 1 15 13 1 15 16 1 9 13 2
2 0 2
15 9 1 15 0 13 9 16 9 13 2 16 1 13 4 2
23 15 7 10 9 7 9 10 9 9 13 2 16 1 0 13 4 2 7 3 13 0 10 2
6 13 3 15 10 0 2
14 15 7 3 13 16 15 15 4 13 13 3 1 15 2
34 15 3 13 4 13 1 15 7 3 1 15 2 16 2 16 13 4 3 1 15 9 2 13 1 15 13 2 16 3 13 1 15 13 2
8 15 3 13 13 16 1 9 2
2 3 2
11 0 1 9 13 9 2 16 9 1 9 2
15 9 7 13 9 9 7 0 9 2 16 1 0 13 4 2
19 15 3 13 10 9 13 2 0 1 13 4 16 15 3 13 13 16 12 2
6 15 7 0 13 9 2
5 13 3 1 9 2
15 15 13 9 7 9 2 9 2 7 10 15 1 15 13 2
4 7 8 12 2
13 10 1 15 13 4 2 7 1 15 13 4 15 2
4 7 8 12 2
18 1 15 10 2 1 15 10 2 7 1 15 10 2 15 9 1 9 2
17 1 15 7 13 0 0 9 2 15 13 9 15 3 13 9 13 2
16 7 3 15 15 13 9 3 13 9 9 9 2 7 0 9 2
9 16 9 1 15 13 9 1 9 2
17 1 15 7 13 16 9 9 1 9 13 1 15 13 16 1 9 2
15 16 3 13 15 9 9 2 7 13 15 15 2 7 3 2
16 16 3 2 13 13 2 3 16 9 15 9 13 1 15 13 2
38 16 7 15 15 13 2 7 13 13 1 0 2 15 3 13 0 1 9 0 2 16 9 13 1 12 0 2 7 13 13 1 15 0 15 15 3 13 2
9 15 3 3 13 13 16 15 9 2
31 13 4 3 1 0 9 16 15 3 13 9 15 9 2 7 13 13 15 1 9 15 9 3 13 9 13 2 16 13 4 2
16 13 3 16 9 1 9 15 9 3 13 9 13 1 15 13 2
2 3 2
10 15 9 1 9 13 13 1 15 9 2
17 13 3 1 9 13 13 9 15 9 2 13 13 1 15 13 9 2
7 15 7 9 13 9 0 2
6 9 3 13 0 13 2
16 9 3 15 13 1 9 9 13 1 15 13 2 13 9 0 2
14 9 7 13 9 16 9 0 13 2 16 1 13 4 2
10 3 15 1 10 9 9 13 3 13 2
2 3 2
25 3 15 9 13 0 2 3 13 0 9 9 2 16 3 9 13 9 2 3 1 0 9 15 13 2
7 13 7 13 0 16 13 2
16 13 3 15 9 0 2 16 3 9 13 2 16 9 7 3 2
22 13 3 16 1 9 15 3 13 16 13 7 13 2 13 15 9 15 13 0 13 9 2
6 15 7 13 13 9 2
9 9 3 3 13 3 13 7 13 2
20 10 7 15 3 13 13 9 1 9 16 1 9 13 2 13 0 13 7 13 2
12 13 3 15 1 9 13 1 9 7 9 15 2
12 3 3 0 13 13 9 1 9 1 9 13 2
2 3 2
16 15 13 3 1 9 7 9 3 13 0 9 15 15 13 9 2
21 3 3 1 9 7 9 13 9 1 3 9 0 2 7 9 15 1 3 9 15 2
11 9 7 13 0 13 9 2 16 13 4 2
12 3 3 15 13 13 3 1 9 7 1 9 2
11 7 3 15 13 13 13 9 1 15 13 2
2 0 2
9 15 9 15 0 13 2 15 9 2
9 13 7 15 9 1 16 9 13 2
27 15 3 9 13 13 9 13 15 9 9 9 13 15 13 9 1 9 15 13 2 7 3 1 15 9 10 2
33 3 9 2 1 12 8 2 13 16 9 0 2 13 9 1 9 2 13 1 0 9 13 9 1 9 2 3 1 9 1 15 13 2
22 9 7 3 13 9 9 1 15 15 13 2 7 1 15 10 9 2 16 1 13 4 2
22 3 0 9 10 9 13 16 13 9 0 15 2 3 0 9 13 2 3 9 1 9 2
14 1 15 7 9 13 10 9 15 9 1 13 3 13 2
10 9 3 9 13 3 13 1 10 9 2
2 3 2
12 9 13 1 9 16 13 9 15 1 15 13 2
15 9 3 15 13 9 16 1 15 2 13 0 16 1 15 2
11 3 13 9 1 15 9 16 13 9 15 2
21 15 3 9 9 1 0 13 13 9 0 7 9 2 7 15 9 9 2 1 15 2
26 9 7 3 13 9 15 15 0 13 1 15 0 13 2 16 10 9 13 10 9 2 16 1 13 4 2
9 3 3 1 13 9 13 9 13 2
2 3 2
28 10 9 15 1 13 13 9 13 2 13 9 13 10 9 2 16 15 13 1 9 9 2 15 13 1 9 9 2
21 15 3 13 1 9 13 15 13 1 10 9 0 2 7 3 3 13 9 1 15 2
9 9 7 3 13 15 9 1 9 2
33 3 3 1 9 13 9 1 9 15 2 16 13 1 9 2 1 12 9 2 1 3 0 9 13 0 0 2 16 1 0 13 4 2
12 9 3 3 13 9 13 1 15 1 9 13 2
2 3 2
6 0 9 0 13 9 2
15 3 3 13 15 9 0 7 0 2 7 9 0 7 0 2
20 15 3 1 15 13 16 13 2 15 13 9 9 2 3 15 9 13 1 13 2
19 3 9 15 13 1 0 13 0 2 16 9 13 9 0 3 1 9 0 2
16 9 0 0 13 9 9 2 3 7 9 13 2 16 9 9 2
13 3 13 3 12 9 15 13 1 9 1 9 0 2
9 15 7 9 13 15 9 0 0 2
7 15 3 15 9 0 13 2
7 3 3 9 1 9 13 2
2 0 2
24 15 1 9 9 13 15 9 7 15 9 2 13 12 15 13 1 15 2 7 9 1 15 12 2
10 13 3 9 1 12 13 13 1 15 2
26 15 9 7 9 13 1 9 2 15 1 0 9 9 13 13 0 2 16 13 3 10 15 13 1 9 2
22 16 3 13 15 9 0 9 13 2 13 7 16 15 13 1 15 2 7 15 1 0 2
18 7 1 9 13 0 9 7 0 9 2 7 13 13 1 15 0 9 2
17 13 3 2 16 13 15 9 13 0 9 2 16 15 15 13 9 2
2 3 2
13 15 13 1 9 0 2 13 13 9 15 15 13 2
17 16 3 3 4 13 2 3 4 1 15 13 2 16 3 13 4 2
61 1 9 7 7 9 15 13 9 16 2 16 1 12 7 15 15 3 13 9 3 9 2 9 13 0 9 16 9 2 16 9 13 0 9 2 3 0 13 2 13 9 9 0 13 2 15 13 1 15 2 16 9 3 13 1 9 16 1 9 9 2
7 7 9 13 9 1 9 2
21 3 13 16 9 2 15 13 9 0 2 13 0 15 0 2 7 1 13 9 15 2
9 3 3 10 9 13 9 1 9 2
2 3 2
12 9 0 15 9 13 2 16 13 9 1 9 2
13 9 7 13 9 10 15 13 2 16 1 13 4 2
7 9 3 13 9 9 0 2
4 15 15 13 2
8 0 3 9 9 13 3 13 2
12 15 7 9 0 9 13 2 13 2 8 12 2
8 1 9 13 9 9 7 9 2
14 15 3 13 15 13 16 1 9 13 15 1 9 13 2
26 1 15 7 13 9 0 9 15 13 9 3 15 9 13 2 15 16 9 0 9 3 13 15 9 13 2
14 1 15 9 13 2 10 0 2 16 1 15 15 13 2
8 15 3 1 0 9 0 13 2
24 1 0 7 9 2 15 13 15 9 0 2 9 3 13 2 15 15 1 10 9 13 0 13 2
8 16 9 3 13 9 7 9 2
28 15 7 13 2 0 13 16 9 9 2 15 13 1 9 13 7 9 13 2 3 13 9 7 9 2 0 13 2
14 9 3 10 7 9 13 9 13 1 9 1 16 3 2
18 1 15 7 9 3 13 15 1 9 15 13 9 2 16 3 13 4 2
7 3 3 13 9 7 9 2
2 3 2
48 0 9 7 9 13 1 15 9 2 7 16 13 1 12 9 2 16 0 2 16 13 1 9 9 7 9 7 1 9 9 2 7 16 13 1 12 9 9 2 16 9 7 9 1 9 7 9 2
7 15 7 13 13 1 9 2
18 9 3 3 3 13 2 7 15 15 9 15 13 9 2 16 13 4 2
9 3 3 13 3 7 9 7 9 2
2 3 2
15 1 10 9 7 9 13 13 15 15 15 13 3 7 0 2
7 15 3 15 9 9 13 2
30 16 7 15 9 9 1 9 13 2 3 13 13 15 15 15 7 15 15 13 2 16 15 13 3 13 2 7 9 13 2
6 3 13 3 9 9 2
2 3 2
25 13 16 9 7 9 9 13 15 15 13 1 9 7 9 2 16 13 4 13 9 9 7 9 9 2
14 3 13 10 9 13 9 7 9 9 2 15 13 0 2
21 7 1 15 2 15 13 3 13 2 16 2 16 13 9 2 15 13 7 3 13 2
20 1 15 7 9 9 2 1 15 13 9 2 3 3 13 15 2 7 13 4 2
25 1 9 7 3 13 15 13 2 16 2 16 15 9 13 16 9 7 9 2 13 15 13 15 9 2
6 15 13 1 9 9 2
8 9 3 3 13 9 7 9 2
8 3 13 15 15 1 9 13 2
47 1 15 7 13 9 13 9 1 9 13 1 9 9 7 9 2 16 16 13 9 2 16 10 9 7 9 2 13 1 15 9 2 7 16 13 3 9 13 1 9 2 16 9 13 1 9 2
17 3 3 13 9 9 2 7 15 9 9 13 1 9 1 15 13 2
7 7 3 13 1 9 9 2
11 3 15 13 15 1 13 13 16 1 9 2
29 13 3 9 13 9 15 1 9 13 3 2 16 3 9 10 13 12 7 15 9 16 3 13 0 2 7 3 13 2
24 13 7 2 16 9 9 15 13 2 16 9 15 13 2 7 7 0 13 2 7 15 9 13 2
16 1 3 9 13 0 13 1 13 2 13 3 9 13 9 15 2
9 10 7 9 1 9 1 9 13 2
8 4 3 1 9 1 9 13 2
16 3 3 15 9 13 2 16 15 9 0 15 1 15 13 13 2
35 16 9 7 9 2 16 1 15 3 13 2 3 7 1 15 13 2 1 9 13 9 9 2 7 2 16 1 15 13 2 3 15 13 13 2
2 3 2
24 9 3 13 1 15 9 2 16 3 13 13 1 0 2 7 1 15 13 2 16 0 9 13 2
18 3 3 15 9 9 13 2 15 15 9 13 2 7 3 1 0 13 2
7 16 1 9 3 13 9 2
11 13 3 1 13 16 10 9 1 9 13 2
6 3 9 0 13 9 2
13 9 7 3 13 9 2 7 9 9 2 16 9 2
7 3 15 13 1 15 9 2
2 3 2
24 1 10 9 0 13 15 0 1 15 0 2 16 0 13 1 15 0 13 0 13 16 1 0 2
19 1 9 7 7 3 9 2 15 13 3 0 9 2 3 13 13 15 0 2
7 3 3 13 3 15 9 2
2 3 2
20 1 10 9 1 15 13 9 2 13 13 1 13 4 2 16 13 1 12 9 2
8 15 7 1 9 3 13 13 2
12 16 13 15 13 13 4 9 2 13 15 9 2
34 15 3 13 13 15 9 1 15 9 13 2 16 15 3 13 1 13 4 2 7 3 1 9 2 3 3 13 13 9 13 2 7 13 2
12 13 3 16 13 13 1 9 15 9 13 13 2
6 15 13 1 9 9 2
8 0 13 3 1 9 9 13 2
2 0 2
8 10 9 0 1 9 13 13 2
9 0 3 7 0 1 9 13 9 2
15 3 7 13 9 2 7 9 2 7 15 1 15 13 9 2
8 15 3 1 9 0 0 13 2
10 3 1 9 9 0 13 13 0 9 2
27 9 7 1 9 13 9 9 13 1 9 7 9 2 16 2 16 15 1 3 9 3 13 2 1 0 0 2
45 1 15 3 13 13 9 1 9 2 7 15 9 2 16 15 1 15 13 9 2 13 0 2 7 1 9 2 16 1 9 0 7 1 9 2 7 1 9 7 9 2 16 1 9 2
6 15 7 0 13 0 2
26 12 9 2 16 15 9 15 13 9 9 2 13 0 1 9 7 9 2 16 13 1 15 13 1 9 2
26 15 9 2 16 15 9 13 1 9 1 15 9 2 16 13 9 0 13 1 9 13 1 9 1 9 2
19 15 7 9 0 9 3 13 0 9 13 2 16 9 3 13 3 7 0 2
10 7 1 9 13 9 2 9 3 13 2
7 3 9 1 9 9 13 2
11 13 3 16 1 9 3 13 13 15 9 2
2 3 2
20 9 1 9 9 1 9 9 13 2 15 3 13 13 1 9 1 9 9 13 2
16 3 2 16 9 3 9 13 13 1 9 2 15 13 1 9 2
44 7 3 13 16 2 16 0 3 13 1 0 9 1 9 2 3 1 9 0 1 9 13 2 7 15 9 13 1 9 0 2 7 0 9 0 1 9 13 2 1 15 13 13 2
34 1 9 7 15 13 1 9 9 2 7 15 13 9 1 13 15 3 1 9 15 13 2 1 13 0 2 16 1 0 15 9 13 4 2
8 13 3 16 9 13 1 9 2
17 3 3 15 2 16 13 2 13 4 2 16 3 13 7 13 4 2
15 7 3 13 16 9 0 9 9 1 0 13 13 2 13 2
8 1 9 13 9 9 7 9 2
8 15 3 9 9 9 9 13 2
11 15 13 13 0 2 16 1 12 9 13 2
6 16 15 9 13 13 2
15 1 15 7 0 13 16 15 9 13 15 1 9 9 13 2
21 15 3 9 13 16 13 2 15 16 13 9 7 13 13 3 2 7 13 7 13 2
15 3 7 13 15 1 15 9 13 2 16 13 1 12 8 2
9 9 7 3 13 9 16 1 9 2
8 15 7 9 13 16 1 9 2
10 15 3 13 1 9 9 2 13 0 2
10 9 7 2 16 13 4 3 13 9 2
11 15 3 13 1 9 15 1 9 9 13 2
2 3 2
15 10 9 15 13 16 13 2 1 9 13 15 1 15 13 2
55 13 3 7 13 13 9 13 7 9 2 15 16 10 9 13 15 0 2 3 2 16 9 2 3 1 15 9 15 13 2 13 16 1 9 13 2 13 16 3 1 13 7 13 15 9 9 13 2 15 1 9 13 3 13 2
12 10 7 9 3 13 16 13 2 16 13 4 2
13 15 3 13 1 9 9 16 1 9 7 9 13 2
12 9 7 3 13 9 7 9 2 16 13 4 2
8 3 15 9 13 15 13 13 2
2 3 2
58 1 9 7 13 13 15 13 0 2 3 13 13 0 15 9 13 15 3 15 10 9 13 2 16 1 0 13 9 2 1 12 8 2 16 9 1 9 2 15 15 15 13 2 3 13 13 9 0 9 2 1 15 0 9 1 9 13 2
38 15 7 9 15 10 9 13 2 16 15 13 2 16 2 1 10 9 13 1 9 15 9 13 2 15 0 1 15 10 9 13 13 15 13 15 9 9 2
20 15 1 15 9 13 13 2 1 10 9 13 9 2 15 16 10 9 13 0 2
11 3 15 9 13 15 13 1 15 15 9 2
6 15 13 1 9 9 2
2 0 2
7 13 3 13 16 9 0 2
32 3 3 13 0 9 9 15 2 3 9 3 1 9 13 1 9 13 13 2 16 15 13 1 9 9 13 2 16 15 1 9 2
41 3 2 16 3 9 13 13 2 13 10 13 9 9 2 7 3 0 13 9 9 15 15 13 15 9 13 2 13 10 9 15 13 13 1 9 9 15 1 9 13 2
15 15 7 9 9 13 0 2 16 13 1 9 1 12 9 2
14 15 3 9 13 15 13 2 15 13 1 15 15 13 2
2 3 2
18 13 7 13 2 13 7 13 2 13 3 13 2 16 13 1 12 9 2
18 9 7 13 3 13 13 10 9 16 1 9 2 15 13 0 13 3 2
9 3 0 13 15 9 13 16 13 2
7 9 7 15 1 15 13 2
21 7 3 2 16 3 13 15 13 1 9 2 16 1 9 13 2 9 13 3 13 2
7 15 3 9 13 13 13 2
36 13 3 9 9 15 13 9 0 9 9 9 9 13 2 1 9 9 13 3 13 16 15 15 13 13 2 15 16 15 13 0 9 7 9 9 2
6 16 0 9 13 13 2
20 1 13 3 13 13 0 16 9 13 0 9 9 2 7 16 15 0 13 13 2
26 1 3 1 9 9 13 9 9 2 15 16 0 9 0 13 9 2 13 16 0 9 13 0 9 0 2
18 9 7 13 0 9 2 15 16 15 15 13 2 10 7 15 13 15 2
13 13 3 9 0 9 0 9 2 15 13 9 0 2
2 3 2
20 1 15 13 4 16 9 13 9 2 16 15 13 13 1 15 1 15 3 13 2
15 15 7 15 15 13 13 2 1 15 15 13 0 9 13 2
11 0 3 9 13 9 2 16 0 15 9 2
2 3 2
44 9 10 9 0 13 2 16 3 9 1 9 9 0 13 2 7 9 1 9 9 15 13 1 9 2 7 0 9 0 9 0 2 0 0 0 2 16 13 9 2 1 12 9 2
6 9 7 13 13 0 2
7 15 1 9 10 9 13 2
14 9 3 0 13 13 9 0 7 0 2 15 9 13 2
19 15 0 9 3 13 9 13 0 2 7 9 13 15 2 16 9 7 0 2
22 9 7 0 1 9 13 2 15 15 13 2 16 3 13 15 13 15 13 1 9 0 2
9 1 15 9 13 15 9 7 15 2
10 3 1 9 13 13 15 9 7 15 2
7 3 9 13 0 9 9 2
2 0 2
20 15 4 13 1 15 9 2 3 13 13 0 9 15 9 2 7 0 7 0 2
41 9 3 2 16 13 10 9 9 2 3 13 13 0 9 9 2 16 2 1 9 10 4 1 15 13 2 13 16 13 15 15 9 2 1 13 15 15 13 1 9 2
19 7 3 13 16 13 0 13 3 9 0 9 15 15 13 9 0 15 9 2
18 7 3 13 16 13 10 9 9 13 13 1 9 0 16 0 1 0 2
17 10 7 15 9 1 9 13 9 13 1 15 2 16 1 13 4 2
16 0 13 3 16 13 9 13 16 16 0 7 13 1 9 15 2
12 9 7 3 13 16 1 13 15 1 9 9 2
9 13 3 9 9 16 13 13 13 2
10 9 7 3 13 9 2 16 13 4 2
9 15 3 9 1 9 13 15 13 2
2 3 2
30 9 13 1 9 15 1 13 2 16 13 0 1 9 0 7 13 7 13 15 2 7 3 9 0 13 1 13 1 9 2
15 3 13 16 13 15 13 0 9 1 15 15 1 9 13 2
6 15 13 1 9 9 2
4 3 15 13 2
18 13 3 16 15 15 1 9 13 13 2 7 16 0 9 7 16 9 2
2 3 2
32 10 9 0 13 9 0 9 1 15 9 0 7 0 15 2 16 9 0 13 9 13 7 13 2 7 9 13 1 9 9 13 2
27 16 3 15 9 13 15 13 1 9 16 9 0 13 2 13 16 15 13 1 15 9 13 7 0 10 9 2
27 9 7 13 9 0 9 13 0 1 9 9 16 9 13 0 9 2 1 15 13 16 0 9 9 0 13 2
16 0 3 13 9 9 16 9 9 2 7 9 9 16 9 9 2
27 13 3 15 4 13 1 0 9 0 13 15 13 0 1 9 9 16 9 2 15 13 9 13 9 0 13 2
5 15 7 13 0 2
33 3 3 15 13 0 2 3 13 0 1 9 9 2 16 0 13 9 16 9 1 9 9 2 16 9 13 2 1 9 1 9 9 2
15 0 13 3 16 15 9 13 2 7 16 0 9 7 0 2
2 3 2
21 15 4 1 15 9 13 2 3 13 13 0 15 9 9 2 13 3 15 15 9 2
31 13 7 13 9 15 9 1 15 2 16 9 13 9 0 9 1 9 2 3 7 0 2 15 16 15 4 13 1 0 9 2
19 15 7 13 9 15 1 15 2 13 13 9 0 15 1 15 13 7 13 2
16 15 3 13 13 1 9 2 15 15 13 15 15 13 1 9 2
12 0 13 3 15 9 13 13 9 15 1 9 2
2 0 2
19 1 10 9 13 1 16 9 13 2 13 9 9 13 1 9 9 15 9 2
12 3 0 15 3 13 1 9 9 2 3 13 2
31 15 3 9 13 1 9 7 9 7 9 2 15 9 13 13 13 1 9 0 9 16 3 2 15 16 10 9 13 15 0 2
22 15 7 15 13 9 13 2 13 13 0 15 15 9 7 9 16 1 9 9 7 9 2
13 3 1 16 13 15 15 2 15 13 1 15 13 2
35 15 3 15 9 13 13 2 13 1 10 9 13 9 15 16 3 1 15 16 13 9 7 9 2 3 7 3 1 15 16 13 1 15 13 2
15 10 3 9 13 13 1 10 9 15 3 13 10 0 13 2
26 3 3 13 2 7 0 15 13 9 15 9 13 0 2 15 13 10 9 13 9 2 16 1 13 4 2
2 3 2
76 1 10 15 13 1 15 13 16 13 2 13 2 16 15 13 13 15 0 13 2 16 15 3 13 1 15 2 7 1 9 2 1 15 0 15 15 0 3 13 2 16 2 16 1 0 13 0 2 13 3 7 0 7 13 2 7 0 1 15 2 16 13 1 3 0 2 13 7 1 9 2 3 0 13 13 2
50 3 3 2 1 13 15 9 2 16 9 7 9 2 9 3 13 1 15 2 16 1 3 9 2 9 7 1 9 2 16 3 1 3 9 0 2 7 1 3 9 15 2 16 9 13 2 1 12 9 2
14 1 3 15 13 3 1 3 9 2 9 1 15 13 2
12 13 3 16 1 15 15 13 1 15 9 13 2
7 3 9 0 13 1 9 2
14 15 7 13 0 9 0 2 15 13 9 9 16 3 2
14 15 0 13 9 13 1 9 2 7 15 9 1 15 2
18 1 3 13 9 3 1 9 13 13 13 2 13 16 0 9 13 13 2
17 15 7 9 0 9 9 13 2 15 9 10 13 13 2 8 12 2
8 1 9 13 9 9 7 9 2
10 9 3 2 1 0 10 9 2 13 2
16 15 0 13 9 9 13 15 9 2 15 10 13 9 15 9 2
7 9 3 13 3 13 9 2
30 1 15 7 13 15 9 9 15 13 9 13 0 9 13 2 7 1 15 4 13 0 2 7 3 15 9 1 1 0 2
5 16 9 10 13 2
14 1 15 7 13 16 0 9 3 13 1 15 12 9 2
25 16 3 0 9 13 13 2 1 15 0 13 4 13 15 1 10 9 13 3 13 16 1 9 9 2
27 3 7 13 10 9 13 2 15 3 13 13 1 9 7 9 2 15 13 3 13 2 7 0 10 9 0 2
13 15 3 2 3 0 13 2 13 9 0 9 13 2
17 15 7 9 13 0 0 9 3 1 9 2 13 13 1 12 9 2
19 13 7 0 2 16 2 16 1 0 13 2 13 13 9 1 9 0 9 2
30 13 3 3 1 9 2 16 15 9 7 15 9 13 0 9 1 9 9 2 16 9 9 2 15 13 9 7 13 9 2
10 9 3 9 3 13 13 1 12 9 2
2 3 2
37 10 9 9 1 15 10 15 13 1 15 10 1 15 7 0 9 15 13 13 2 16 0 1 10 15 13 2 16 9 13 2 15 13 9 13 9 2
21 9 7 0 13 1 15 9 13 2 7 9 13 15 0 9 2 16 1 13 13 2
12 3 1 10 15 15 13 15 9 9 3 13 2
23 16 3 1 15 3 9 9 15 13 2 3 13 1 15 9 9 16 3 2 7 15 9 2
12 9 7 9 13 13 9 2 15 13 3 9 2
13 10 3 9 13 15 1 15 9 3 9 3 13 2
7 15 7 13 15 9 13 2
11 13 3 16 15 9 3 13 2 9 13 2
2 3 2
7 10 9 13 16 9 13 2
13 1 3 9 9 15 9 13 9 10 9 1 13 2
9 9 3 13 9 2 7 9 9 2
17 9 7 13 9 9 2 1 15 10 9 13 2 16 1 13 4 2
22 13 3 10 9 0 9 2 1 10 15 13 15 3 13 9 15 15 13 9 1 9 2
8 15 7 13 0 15 9 13 2
7 10 3 1 15 9 13 2
2 0 2
7 10 9 0 13 9 0 2
11 9 3 1 9 13 2 16 9 1 9 2
18 3 13 7 9 1 9 13 16 13 9 16 1 9 15 13 1 9 2
25 0 3 13 9 16 13 9 0 9 15 15 1 9 13 13 2 1 3 15 13 0 1 9 9 2
36 7 1 15 9 13 16 10 15 13 1 9 9 0 7 0 2 13 13 1 9 1 9 0 15 13 1 9 0 2 15 13 0 0 1 9 2
21 16 7 9 0 13 0 9 9 9 9 2 3 9 13 0 9 9 15 9 13 2
18 15 3 13 1 9 9 13 2 15 15 9 1 10 9 0 13 13 2
26 1 9 7 9 13 13 10 15 9 13 3 13 2 16 1 9 9 0 13 10 15 9 0 3 13 2
5 10 3 9 13 2
2 3 2
14 16 9 15 3 13 9 15 9 2 13 1 12 13 2
14 12 9 2 1 15 16 3 13 1 9 9 7 9 2
9 9 3 10 13 15 0 15 9 2
24 3 9 15 13 1 9 9 2 3 13 13 0 7 9 2 9 7 13 2 15 3 13 13 2
23 15 9 2 1 9 9 2 15 13 9 9 0 2 16 9 0 0 3 13 13 9 13 2
37 0 9 2 1 9 13 1 9 2 1 15 9 13 3 13 2 16 0 3 13 13 9 2 16 10 9 3 13 13 1 9 2 1 15 13 9 2
11 15 7 15 9 13 15 9 13 0 9 2
28 7 3 1 9 9 15 15 0 13 13 2 1 10 9 2 16 13 9 2 13 15 0 2 16 1 13 4 2
20 3 3 1 9 9 2 1 13 4 16 9 13 1 10 9 1 9 7 9 2
21 3 3 1 9 9 2 1 15 13 9 9 2 15 3 0 13 13 16 1 9 2
18 15 3 1 13 3 13 9 2 1 2 15 13 2 9 1 9 13 2
14 7 3 1 9 9 15 9 13 3 13 1 9 9 2
22 13 3 16 0 9 3 13 1 15 9 2 7 0 10 13 2 15 13 15 13 0 2
11 15 13 16 3 0 9 9 13 15 13 2
9 13 3 8 12 2 1 9 9 2
4 15 9 0 2
7 13 1 15 7 13 9 2
4 7 9 12 2
5 13 16 10 13 2
8 7 9 12 2 1 9 9 2
8 3 13 0 1 9 10 9 2
42 1 15 7 13 15 9 9 15 13 1 9 0 13 12 9 3 2 16 9 15 1 15 9 13 13 2 7 16 9 3 13 15 13 16 1 16 9 9 0 15 13 2
6 1 15 13 9 12 2
8 16 15 13 0 2 13 15 2
8 16 9 3 13 1 9 9 2
19 1 15 7 13 16 9 13 1 9 3 1 9 9 2 7 1 9 9 2
12 10 3 9 1 9 9 9 13 1 12 9 2
19 7 3 13 16 10 0 3 13 15 9 2 16 13 9 2 3 7 0 2
15 0 7 9 3 13 1 12 9 3 2 16 1 13 4 2
12 9 3 3 13 1 9 9 2 7 1 9 2
2 3 2
13 15 3 13 9 2 13 0 9 2 16 13 4 2
44 0 7 3 13 1 9 13 15 3 2 16 13 2 9 3 13 2 16 13 0 1 9 2 9 7 9 9 7 15 9 2 1 15 16 15 15 13 9 9 2 9 3 13 2
12 0 3 13 0 9 15 1 9 9 3 13 2
24 15 7 15 15 13 13 15 13 7 15 3 13 2 13 1 9 9 2 7 3 1 9 9 2
12 9 3 3 13 1 9 9 2 7 1 9 2
2 3 2
13 15 9 15 9 13 1 16 9 13 13 1 15 2
7 10 3 9 13 15 0 2
17 10 7 15 13 1 15 2 13 1 15 1 9 15 1 15 13 2
26 1 3 9 13 1 9 10 13 2 16 1 13 4 2 13 16 9 9 15 13 1 15 1 9 0 2
5 3 1 9 13 2
22 9 7 3 13 15 9 16 13 9 2 15 9 13 9 13 2 15 13 9 16 9 2
11 9 3 1 9 13 2 3 1 9 9 2
2 0 2
11 1 9 2 1 12 8 2 0 13 9 2
13 12 15 13 1 9 7 13 9 15 2 16 13 2
15 15 15 13 1 0 7 13 9 13 2 16 13 1 9 2
28 0 7 9 3 13 13 1 9 15 9 15 3 13 1 9 2 1 10 9 13 10 9 2 16 1 13 4 2
18 13 3 16 13 1 9 15 9 15 13 1 9 7 13 3 9 15 2
17 3 7 3 13 16 9 13 7 13 2 9 3 13 7 13 13 2
11 3 3 1 9 9 2 7 1 9 9 2
2 3 2
31 9 13 1 9 1 15 0 13 13 16 0 3 13 1 9 2 7 1 15 9 13 2 16 1 9 13 2 1 12 0 2
13 0 7 9 1 9 13 13 9 1 9 7 9 2
16 15 3 15 9 13 2 13 1 9 16 1 9 1 15 13 2
6 15 3 1 0 13 2
11 3 9 9 13 1 13 9 1 9 13 2
8 0 7 13 13 7 1 0 2
29 1 15 3 16 15 0 1 9 13 13 2 13 9 15 9 2 7 15 15 13 1 9 2 7 13 9 1 15 2
5 15 0 13 13 2
18 1 3 9 13 0 9 2 3 13 1 9 9 2 7 9 7 9 2
2 3 2
13 15 1 15 13 2 0 13 15 15 1 15 13 2
21 10 3 15 13 1 15 2 13 13 1 15 15 1 15 13 2 16 1 0 13 2
13 15 7 10 9 3 13 9 2 3 1 15 13 2
12 13 3 3 1 15 9 2 3 3 15 13 2
13 13 3 0 9 15 9 13 16 15 9 9 13 2
11 3 13 7 15 15 9 9 16 1 9 2
18 13 3 9 2 15 13 0 9 2 1 9 13 2 3 1 9 9 2
2 3 2
13 0 9 13 0 9 2 16 7 0 0 0 9 2
10 7 0 9 9 13 0 16 9 9 2
17 15 3 0 0 13 16 13 9 2 16 1 12 15 13 9 0 2
8 9 7 9 1 9 13 9 2
21 15 1 15 13 16 9 13 15 1 15 15 1 9 13 2 16 15 1 9 9 2
15 3 9 2 15 13 0 9 2 13 9 15 13 1 9 2
2 0 2
29 1 15 15 13 16 2 16 13 15 9 2 0 13 9 15 13 1 9 15 15 13 1 9 7 13 15 3 9 2
22 3 1 9 0 13 9 2 15 13 1 9 2 16 9 0 2 15 13 1 9 9 2
9 0 7 9 13 0 1 10 9 2
14 3 15 13 1 9 10 1 9 2 3 1 9 9 2
2 3 2
27 9 13 1 9 9 1 9 9 2 9 7 3 13 1 0 9 9 2 7 1 15 9 15 13 10 9 2
34 1 3 10 9 13 1 16 1 9 13 2 16 9 13 9 2 13 16 9 1 9 1 9 1 9 9 13 16 9 0 1 9 0 2
17 9 7 0 15 13 1 9 0 16 15 0 2 7 16 15 9 2
15 3 13 16 0 9 13 0 2 7 3 1 9 9 13 2
8 15 3 9 0 9 15 13 2
5 13 3 1 9 2
6 10 15 13 9 13 2
4 7 8 12 2
8 15 13 10 1 13 9 10 2
8 7 9 2 1 9 1 9 2
7 10 9 9 9 9 13 2
3 7 1 2
12 15 3 10 13 13 2 15 9 15 13 13 2
15 1 15 7 13 9 15 9 15 13 9 13 1 9 9 2
7 16 9 13 1 10 9 2
13 1 15 7 13 16 9 9 10 13 1 10 9 2
9 9 3 1 13 1 15 9 13 2
7 9 3 13 13 9 9 2
11 9 7 13 9 1 9 2 16 13 4 2
32 1 3 1 9 3 13 16 0 9 2 15 7 13 16 13 15 2 15 13 13 0 13 2 13 16 10 9 1 10 9 13 2
2 3 2
6 10 9 13 15 0 2
23 3 13 16 1 15 13 15 9 1 16 13 9 15 9 2 16 9 13 1 9 15 9 2
18 7 1 15 9 1 9 2 16 3 2 13 9 15 9 1 9 9 2
25 16 3 1 9 9 0 13 9 9 9 0 2 3 13 16 12 2 16 9 0 12 13 12 3 2
11 10 3 9 0 13 9 1 9 15 9 2
10 9 7 13 1 9 2 16 13 4 2
10 3 1 9 15 9 9 1 9 13 2
2 0 2
11 1 9 2 1 12 8 2 13 0 13 2
27 9 3 15 13 3 13 16 1 9 9 7 9 13 1 3 2 7 1 15 9 15 2 15 13 9 15 2
12 9 3 15 1 3 13 1 9 15 1 9 2
23 13 7 9 7 9 15 1 3 13 0 13 9 2 13 7 1 15 1 9 9 9 13 2
12 7 3 13 16 10 9 1 9 15 13 13 2
11 3 7 1 0 9 9 0 15 9 13 2
22 9 7 15 4 1 9 13 2 9 1 3 13 3 0 2 1 13 3 7 1 0 2
12 7 3 13 16 9 9 1 9 13 15 13 2
10 9 3 1 10 9 9 1 9 13 2
2 3 2
29 15 15 13 1 9 2 7 13 0 2 16 9 9 2 15 13 9 13 2 7 13 1 0 9 2 15 0 13 2
12 7 3 13 16 9 13 4 1 9 16 13 2
10 0 7 9 13 9 2 16 9 13 2
12 13 3 10 9 13 1 9 16 9 1 9 2
13 7 9 1 9 10 9 7 9 9 1 9 13 2
11 3 7 9 10 9 1 9 15 9 13 2
6 15 7 0 9 13 2
5 3 13 1 9 2
5 10 1 9 13 2
4 7 8 12 2
5 9 9 13 9 2
19 1 15 7 13 15 9 15 13 10 1 0 0 9 13 2 1 15 9 2
7 15 0 13 15 3 13 2
18 1 13 7 13 13 16 2 16 9 13 0 2 15 3 13 3 13 2
10 13 3 4 1 1 9 13 9 0 2
14 9 0 0 1 15 3 13 3 1 1 0 4 13 2
7 1 7 15 9 13 13 2
11 15 3 9 3 13 15 13 9 0 13 2
8 15 7 3 13 2 13 4 2
15 0 3 3 9 0 1 13 13 2 9 7 0 1 13 2
14 3 1 15 0 13 9 1 13 15 9 13 9 9 2
19 1 3 1 9 0 9 3 13 2 15 1 10 9 13 2 9 3 13 2
11 3 13 3 9 13 9 2 7 15 3 2
2 3 2
7 15 9 0 9 9 13 2
13 9 3 2 15 9 0 3 13 2 13 3 13 2
29 13 7 0 13 16 3 13 13 1 0 9 9 2 16 16 3 13 13 7 13 2 7 13 2 7 13 7 13 2
2 0 2
13 1 13 15 13 13 2 13 16 1 15 13 13 2
2 3 2
7 9 10 1 9 15 13 2
7 9 7 9 9 9 13 2
6 15 3 9 13 13 2
2 3 2
21 1 9 13 1 9 9 2 9 7 1 9 9 2 13 16 7 13 7 13 13 2
2 0 2
6 7 13 7 9 13 2
11 15 3 3 13 16 15 15 13 4 13 2
20 0 7 7 13 13 2 7 13 7 13 2 1 15 10 1 9 7 9 13 2
2 3 2
52 16 9 0 9 7 9 13 9 13 2 15 7 9 9 13 16 13 9 15 9 2 16 9 3 13 13 0 1 9 2 13 16 9 13 3 13 15 13 1 9 9 16 13 9 2 7 13 9 16 4 13 2
8 15 7 13 3 2 13 13 2
12 0 3 3 1 9 9 13 15 9 9 13 2
18 13 7 9 9 1 10 13 2 16 9 9 1 13 15 7 9 15 2
7 13 7 9 13 3 9 2
23 15 3 9 3 13 2 16 13 3 12 7 15 13 7 3 13 2 15 13 0 13 3 2
2 3 2
7 9 0 7 0 13 13 2
30 13 3 2 16 13 0 7 0 2 16 13 0 7 3 0 2 7 16 13 13 7 0 2 16 13 13 7 3 13 2
17 3 15 9 3 13 16 9 3 13 13 13 3 13 15 1 15 2
2 0 2
10 1 9 15 9 0 13 9 15 9 2
34 16 3 9 3 13 13 9 3 13 7 3 13 2 7 3 13 13 16 9 13 15 10 9 0 15 13 2 16 16 9 3 13 9 2
2 3 2
68 1 9 15 9 2 16 0 2 9 7 9 2 13 1 0 9 0 9 2 1 15 9 9 13 2 13 16 0 15 9 9 13 3 13 2 16 16 9 3 13 0 1 9 2 7 16 9 13 1 9 1 9 3 13 0 2 7 16 0 0 3 13 12 9 0 12 13 2
13 15 3 13 16 9 3 13 13 16 13 3 13 2
6 3 15 3 9 13 2
15 15 3 9 13 15 13 16 13 2 7 15 13 16 13 2
11 13 3 15 15 13 9 9 13 16 3 2
7 15 3 9 13 3 13 2
10 3 10 15 13 9 2 13 4 13 2
11 1 15 7 13 16 9 3 13 13 9 2
14 3 1 9 9 13 13 16 9 10 1 15 9 13 2
14 15 13 1 9 15 15 13 9 2 16 1 0 13 2
12 15 3 9 2 3 13 9 13 15 0 15 2
30 3 15 15 9 1 15 3 13 2 0 13 1 13 7 1 10 9 15 15 1 15 13 2 15 1 9 9 13 13 2
14 0 3 9 13 3 13 16 15 13 1 9 1 15 2
9 3 9 9 15 13 1 9 10 2
10 3 13 16 2 13 9 2 13 9 2
19 16 3 9 15 13 13 15 1 9 3 13 1 13 2 3 13 9 15 2
2 3 2
16 16 15 13 1 9 9 2 15 3 13 13 15 3 13 13 2
18 15 7 13 3 13 2 13 13 16 13 15 1 0 9 9 13 13 2
22 3 15 0 13 13 2 0 13 3 13 2 7 15 0 13 13 2 0 13 3 13 2
38 13 7 1 15 16 3 13 9 13 15 3 13 2 7 3 13 0 7 0 2 16 1 9 13 15 13 2 0 13 7 0 2 16 1 0 13 4 2
12 3 13 4 1 16 9 3 13 13 15 9 2
8 3 13 16 9 13 3 13 2
12 0 13 4 1 16 9 9 3 13 13 0 2
15 3 3 3 13 13 15 15 4 1 15 13 2 3 13 2
12 13 3 16 15 15 9 13 3 13 1 13 2
10 3 13 0 9 7 13 7 13 13 2
27 3 7 13 3 9 7 13 7 13 2 16 15 9 7 9 0 13 2 3 7 16 13 13 9 1 13 2
18 3 9 0 9 9 9 3 13 16 1 9 2 16 1 0 13 4 2
24 7 3 10 15 9 2 9 3 13 13 0 15 15 13 13 2 7 15 0 13 2 13 13 2
9 3 3 13 9 0 9 1 13 2
16 16 7 13 13 2 13 0 2 16 13 9 7 9 9 0 2
17 16 7 9 13 1 9 2 3 7 1 9 7 9 16 13 4 2
33 0 3 9 3 13 13 15 15 13 3 13 2 7 13 15 15 13 13 2 15 3 13 13 15 13 3 13 2 7 13 15 13 2
26 7 15 9 13 7 13 15 2 16 3 13 3 13 13 2 3 3 0 2 7 1 9 7 1 9 2
9 16 0 9 3 13 1 13 9 2
70 16 7 13 4 16 0 9 1 13 9 3 13 2 7 1 15 16 1 9 9 3 13 2 7 1 9 7 9 2 16 15 9 13 16 15 9 7 9 1 13 9 3 13 13 2 7 3 13 1 9 9 2 16 3 1 9 9 2 13 13 16 15 9 7 9 15 9 9 13 2
36 13 4 3 1 16 9 10 15 15 1 15 13 13 13 10 9 13 2 1 15 10 3 13 0 13 1 0 9 2 16 9 9 13 1 9 2
25 16 3 9 0 1 9 13 3 13 2 16 1 13 4 2 0 13 7 1 15 9 0 9 13 2
2 3 2
6 0 9 9 1 13 2
23 0 7 2 15 9 13 13 2 13 3 13 16 0 13 15 13 2 16 3 9 0 13 2
24 15 7 15 1 9 13 13 1 9 0 2 1 10 15 1 9 9 1 13 9 7 9 13 2
17 0 3 7 15 0 9 13 2 3 1 0 9 13 16 15 13 2
7 7 3 0 9 13 13 2
20 0 3 9 2 15 9 0 9 13 2 16 1 13 4 2 10 9 9 13 2
11 3 3 1 9 1 15 7 15 9 13 2
2 3 2
10 1 13 4 16 0 9 0 13 9 2
11 9 7 1 15 9 9 9 13 1 9 2
10 9 3 0 9 1 13 9 3 13 2
2 0 2
26 16 0 9 9 1 9 15 2 3 1 9 13 2 13 2 15 13 9 15 15 1 15 13 1 9 2
22 15 7 13 3 13 2 1 1 13 4 16 9 13 3 15 3 13 7 13 7 13 2
11 3 3 9 13 1 9 15 9 7 9 2
2 3 2
15 0 9 13 1 9 1 15 13 16 9 9 1 9 13 2
23 15 7 9 15 13 1 10 15 13 13 1 9 13 15 9 2 16 9 0 1 10 9 2
22 9 7 13 0 9 13 9 2 1 15 1 10 9 13 0 9 9 2 16 13 4 2
15 3 9 0 1 10 15 9 9 3 13 2 10 9 13 2
15 3 3 10 2 3 13 1 15 2 13 4 1 9 13 2
10 3 3 0 9 1 15 13 9 13 2
7 15 13 15 1 9 13 2
15 0 9 2 7 0 9 15 2 7 9 15 3 13 9 2
40 1 15 7 13 15 9 9 13 16 1 15 16 9 15 13 2 13 1 15 1 9 15 9 9 2 16 3 10 9 13 0 7 0 13 2 16 9 0 13 2
26 13 3 16 2 16 0 9 1 0 9 3 13 2 15 3 15 13 13 9 15 1 10 9 0 13 2
5 16 9 12 13 2
11 10 1 9 2 9 7 9 13 2 9 2
9 16 0 9 1 13 9 3 13 2
20 1 15 3 13 13 16 7 15 9 2 1 15 13 2 1 13 9 9 13 2
8 9 3 10 9 13 13 13 2
13 9 7 9 13 9 13 2 16 13 1 1 13 2
17 9 3 1 15 15 13 4 13 15 15 9 1 9 9 13 13 2
25 16 3 9 0 1 0 9 3 13 2 16 13 4 2 13 16 7 0 9 13 9 1 9 13 2
2 3 2
9 15 13 1 9 13 15 3 13 2
16 13 4 7 1 16 9 1 15 1 15 15 13 1 9 0 2
16 3 3 1 9 0 9 15 9 13 2 7 1 15 0 9 2
7 15 1 9 9 9 13 2
24 13 3 1 13 13 16 9 3 1 9 13 4 1 9 9 16 1 9 9 9 1 9 13 2
18 9 3 2 1 9 2 1 12 8 2 1 15 13 2 15 9 13 2
10 0 7 9 9 15 13 15 15 13 2
12 15 3 0 9 9 1 9 9 13 3 13 2
2 3 2
26 1 9 9 13 13 15 15 10 13 2 9 9 13 9 15 15 15 10 13 2 16 1 9 0 13 2
14 15 3 13 13 10 13 15 9 1 9 9 15 13 2
16 15 3 9 15 0 15 10 15 13 2 3 13 13 9 9 2
11 7 1 9 9 13 0 13 15 10 13 2
8 3 3 9 1 9 9 13 2
2 3 2
27 15 13 15 15 16 1 15 16 0 13 1 15 2 7 15 13 1 15 7 1 15 2 9 15 15 13 2
36 3 3 9 13 9 9 2 16 13 9 1 15 2 9 9 2 16 1 15 13 9 15 13 2 10 9 0 1 9 2 1 15 9 10 13 2
21 7 9 1 15 13 2 7 13 15 15 1 15 13 2 16 1 1 13 0 13 2
12 9 3 3 13 9 1 9 1 15 9 9 2
2 0 2
15 1 15 9 15 13 1 15 13 0 15 15 13 1 15 2
16 15 3 15 13 0 0 1 10 9 2 13 9 1 15 3 2
13 15 7 13 1 9 9 2 3 13 1 15 3 2
7 13 3 1 15 15 13 2
20 9 3 2 1 13 0 9 7 0 9 2 9 1 9 3 13 1 9 9 2
7 15 13 15 8 12 13 2
9 15 0 13 15 2 7 13 15 2
12 16 1 15 7 1 15 7 1 15 13 10 2
4 7 9 12 2
9 15 1 13 15 2 16 13 15 2
9 10 15 1 9 13 2 10 13 2
25 1 15 7 13 9 15 13 13 16 9 3 13 13 16 15 13 2 16 3 13 13 16 15 13 2
12 3 3 1 9 9 9 13 2 16 13 4 2
24 16 7 0 9 9 15 13 13 15 15 13 13 13 2 13 3 15 0 2 15 13 9 9 2
6 15 3 0 13 13 2
26 15 3 0 9 13 16 9 7 0 9 1 13 2 1 9 2 15 13 2 16 9 0 13 2 13 2
14 9 7 15 7 9 13 16 15 15 9 1 9 13 2
15 16 3 15 0 9 0 13 2 15 9 1 9 9 13 2
44 13 3 12 9 15 15 13 1 9 15 1 15 2 16 3 1 15 13 13 15 1 15 13 2 16 13 13 9 16 15 1 9 9 13 2 16 15 15 13 9 15 15 13 2
29 15 3 9 9 1 9 9 9 3 13 2 1 3 13 15 13 15 13 13 15 9 13 2 7 15 15 9 13 2
9 15 9 13 15 15 13 1 15 2
13 15 3 13 1 9 15 13 15 1 15 9 13 2
17 16 9 13 13 13 9 7 9 2 16 1 15 9 13 3 13 2
10 0 7 9 15 0 13 1 15 9 2
11 3 13 3 1 9 9 15 13 9 9 2
2 3 2
13 9 10 9 9 1 9 13 2 16 1 13 4 2
19 3 13 7 0 2 16 9 10 9 13 13 2 16 13 15 1 15 13 2
11 15 3 0 13 13 0 2 3 7 13 2
22 13 4 3 1 0 9 16 9 1 9 13 10 9 13 2 3 7 1 9 13 15 2
10 3 3 1 9 13 0 9 9 9 2
2 0 2
24 13 4 16 9 13 9 1 9 3 1 9 9 2 7 1 9 9 2 7 9 2 7 9 2
14 15 3 9 9 0 9 13 13 16 9 1 9 13 2
11 13 3 13 13 15 13 1 9 15 9 2
8 9 7 0 13 9 9 13 2
13 15 3 1 9 15 13 2 1 9 9 15 13 2
34 16 3 9 9 3 13 13 13 1 9 9 15 9 9 13 9 2 3 3 1 15 9 9 15 10 9 13 9 2 16 9 0 13 2
17 0 3 9 13 2 13 13 1 9 9 9 2 16 0 13 9 2
26 16 0 0 9 13 15 9 13 10 9 7 9 9 1 9 13 2 3 9 9 1 9 0 9 13 2
16 3 3 13 13 16 9 15 15 13 13 15 3 15 3 13 2
9 15 15 9 7 13 0 7 0 2
9 15 3 9 1 9 13 16 13 2
25 7 3 15 9 3 13 1 9 9 0 13 1 9 9 2 1 15 13 3 13 16 9 9 13 2
19 15 7 1 15 3 13 9 0 13 2 16 13 1 9 2 1 12 9 2
26 3 3 0 13 13 16 9 1 9 9 9 1 9 13 2 15 9 16 1 9 7 9 15 13 13 2
19 16 7 15 9 9 13 2 13 3 9 9 13 1 9 0 9 1 0 2
10 13 7 0 3 0 9 2 7 9 2
11 3 3 1 0 0 9 13 13 3 13 2
11 1 0 0 9 13 9 2 9 3 0 2
20 3 16 15 15 13 0 0 2 13 3 0 1 9 2 0 1 0 9 13 2
15 13 3 13 16 2 13 9 2 13 9 1 15 13 9 2
32 16 0 15 13 0 0 2 13 0 1 9 2 3 1 0 0 9 13 1 0 2 16 9 13 13 13 1 15 16 9 13 2
25 3 7 15 0 13 2 16 9 7 9 13 1 15 15 13 0 9 2 1 15 15 13 9 0 2
34 9 7 15 13 1 0 1 9 16 13 0 9 2 3 13 0 9 2 7 0 2 16 2 16 15 13 13 2 0 13 15 0 13 2
11 1 3 15 9 1 9 9 9 13 0 2
20 0 2 16 13 13 9 1 15 9 9 1 15 15 9 15 1 9 13 0 2
25 16 3 15 0 13 9 13 2 13 13 16 9 7 9 13 2 7 3 1 15 0 13 3 13 2
33 0 2 16 13 9 9 1 12 9 1 15 2 16 2 16 9 7 9 9 13 13 2 13 13 16 0 9 13 2 1 15 13 2
33 7 16 9 13 13 2 13 13 9 7 9 2 7 15 3 15 9 13 1 9 9 2 16 7 15 7 15 1 0 9 13 9 2
69 0 2 16 1 15 9 13 0 9 1 10 9 7 9 7 9 2 1 15 13 9 3 1 9 7 3 1 15 15 9 2 16 2 13 16 9 9 13 13 2 13 1 15 9 13 16 9 7 9 1 15 13 2 7 9 2 7 15 3 9 2 3 0 16 0 2 15 13 2
19 1 15 10 2 16 0 13 2 9 9 9 3 13 2 7 10 9 13 2
16 13 7 7 15 9 9 1 9 9 1 16 15 13 0 0 2
22 15 3 9 13 1 9 0 1 9 2 16 1 9 0 2 7 1 9 13 7 13 2
17 7 15 9 9 1 0 9 9 9 13 3 13 3 1 9 13 2
18 3 3 0 9 9 13 13 2 15 13 0 13 2 16 1 13 4 2
16 15 7 3 9 9 2 7 9 13 13 2 16 1 13 4 2
30 15 0 15 9 13 2 9 13 3 13 16 1 0 9 9 2 1 15 13 13 9 16 15 13 1 15 13 1 9 2
19 7 3 1 9 0 7 0 2 15 13 3 1 0 9 9 9 0 13 2
19 1 15 3 16 15 9 1 9 4 13 2 0 13 15 0 7 0 13 2
21 7 1 15 16 15 9 13 13 0 9 2 0 13 16 12 9 0 12 13 13 2
14 15 7 9 13 1 9 9 1 9 13 0 7 0 2
17 16 1 15 9 9 13 3 13 2 7 3 1 9 9 9 13 2
29 1 9 7 9 2 16 3 9 13 13 2 13 13 9 0 1 9 13 13 2 16 1 9 9 9 9 0 13 2
23 3 3 1 13 9 9 9 0 1 9 13 7 3 1 9 9 2 7 3 1 15 9 2
12 7 3 9 13 0 7 0 10 13 7 13 2
8 3 3 1 13 13 0 9 2
43 15 3 15 2 0 9 13 2 13 9 3 13 13 16 15 13 2 16 3 13 13 2 7 15 15 13 16 10 13 0 9 2 1 15 15 9 7 13 1 9 7 13 2
9 15 1 9 13 13 13 9 0 2
43 16 7 10 1 9 9 13 16 1 0 9 2 15 1 13 9 3 13 16 1 15 13 9 2 3 3 1 15 0 9 1 9 13 2 16 13 0 15 13 10 13 13 2
34 2 15 13 15 13 2 1 15 16 1 9 10 3 1 9 13 13 2 1 13 1 9 13 13 9 15 1 9 10 3 1 9 13 2
14 13 3 15 1 9 13 15 0 7 0 0 13 13 2
18 15 3 9 0 7 0 0 13 13 1 15 3 13 9 1 3 13 2
20 15 7 9 3 4 1 9 1 9 13 16 1 15 9 13 9 1 3 13 2
16 15 3 13 1 15 16 9 1 15 13 1 9 1 15 9 2
29 15 3 9 1 15 7 3 13 9 2 7 2 16 13 2 3 13 0 1 15 9 2 3 13 9 1 3 13 2
9 15 3 0 7 0 0 13 13 2
35 16 7 13 16 15 15 13 1 15 2 3 13 1 15 1 15 13 2 7 3 10 9 13 9 1 3 13 2 2 0 13 15 3 13 2
14 13 3 9 13 15 9 1 15 13 15 13 1 15 2
9 15 3 3 13 16 1 9 9 2
44 3 3 7 9 13 3 13 9 1 3 13 2 7 9 13 9 16 15 13 9 7 15 13 9 13 2 1 3 1 9 9 13 1 9 9 2 7 1 9 2 16 13 4 2
2 3 2
21 1 15 9 13 1 0 9 1 9 13 2 13 15 15 13 15 9 15 13 13 2
43 1 15 7 16 13 9 13 9 1 13 1 9 2 3 1 9 2 3 13 16 13 15 9 13 15 1 9 13 7 15 15 13 13 2 1 15 16 13 1 9 9 13 2
11 15 3 13 9 15 0 9 13 0 13 2
2 3 2
23 1 0 9 13 16 9 13 10 9 13 2 16 3 1 15 15 13 15 15 13 9 13 2
11 9 3 9 13 13 15 0 3 0 13 2
11 13 7 0 0 3 13 1 9 9 13 2
17 15 3 13 15 13 0 15 3 10 9 9 13 2 16 9 9 2
18 15 3 13 15 9 3 4 13 1 9 16 3 15 13 13 0 0 2
6 3 15 0 9 13 2
2 0 2
23 3 15 3 13 1 15 15 1 15 13 9 2 3 9 2 3 3 0 13 1 3 9 2
14 3 3 15 13 0 9 2 3 3 13 1 3 9 2
19 15 7 9 13 2 0 13 1 3 9 1 15 16 13 9 1 3 9 2
37 15 3 15 13 9 0 2 7 1 15 1 3 9 13 2 15 13 13 2 1 15 16 13 9 9 0 2 16 1 15 3 13 9 1 3 9 2
6 15 7 13 0 0 2
9 3 3 15 13 1 9 13 9 2
34 13 13 3 16 2 16 9 13 9 13 16 13 1 0 9 2 13 13 1 9 2 3 1 9 9 2 16 9 9 2 16 13 4 2
12 16 0 13 1 9 0 2 13 9 13 0 2
46 15 3 13 15 9 3 1 9 13 2 15 3 13 2 1 9 13 15 9 2 16 9 9 15 0 9 13 1 15 16 3 1 0 13 13 2 16 15 1 0 13 3 13 0 0 2
13 0 7 16 15 9 9 1 9 13 2 0 13 2
16 16 7 2 15 3 13 2 15 13 7 13 2 0 9 13 2
11 9 7 1 0 9 9 13 1 9 13 2
34 3 16 1 10 0 9 2 15 13 9 7 9 2 9 13 3 13 2 15 1 9 9 0 9 13 2 0 9 1 10 13 0 13 2
18 1 15 7 9 2 1 16 13 13 9 2 0 13 9 0 1 9 2
12 12 3 9 2 1 9 1 9 15 15 13 2
51 7 16 9 2 1 15 15 13 2 9 1 9 13 2 15 7 13 13 2 13 3 7 3 13 2 1 9 9 0 9 15 0 13 2 16 9 16 1 0 13 13 2 7 9 16 15 9 13 0 0 2
18 9 7 2 1 15 15 13 2 9 13 2 7 1 15 9 9 13 2
10 3 1 15 13 9 1 13 1 15 2
12 15 13 7 16 9 15 13 9 3 1 9 2
26 7 3 3 13 15 9 1 3 13 2 7 1 10 9 3 13 1 9 13 2 16 13 1 9 13 2
33 7 16 9 15 10 9 13 15 9 9 2 16 3 3 13 9 1 15 9 2 7 1 13 1 3 13 2 16 13 1 9 0 2
19 1 15 0 9 3 13 15 9 9 2 13 3 1 9 9 1 15 9 2
27 7 3 3 13 1 15 9 13 2 7 9 13 13 1 15 9 9 1 9 2 16 13 1 9 7 0 2
11 9 3 9 3 13 9 1 15 15 13 2
16 3 3 13 0 9 9 12 16 1 15 16 13 15 9 9 2
13 9 0 13 13 9 1 16 13 1 13 9 9 2
16 15 7 9 13 13 0 7 0 10 2 15 13 1 9 0 2
17 3 0 13 16 10 15 7 0 13 7 1 0 13 2 0 13 2
29 15 7 3 3 13 2 0 13 2 16 1 9 13 2 16 9 15 3 13 7 9 15 13 1 15 16 13 9 2
29 15 0 9 1 9 0 13 1 9 0 9 1 9 1 9 9 7 9 2 16 13 3 9 1 15 3 0 13 2
28 16 3 9 0 9 13 9 13 7 13 7 13 2 0 13 0 9 15 9 7 9 7 9 0 1 15 13 2
26 0 2 16 9 13 9 0 0 2 7 15 13 9 7 9 9 2 0 13 15 7 9 7 0 13 2
37 0 9 13 1 9 9 0 1 9 9 0 1 9 13 9 7 9 2 16 0 13 9 2 16 1 9 13 2 0 13 2 7 9 9 0 13 2
16 9 0 9 13 7 3 1 15 13 2 7 3 1 9 13 2
14 0 7 9 9 0 13 9 9 15 13 1 9 0 2
22 16 3 15 9 1 9 9 0 13 2 3 7 9 1 9 9 1 15 9 13 9 2
7 3 3 13 16 9 13 2
28 13 3 15 13 1 9 15 1 15 9 13 2 16 13 7 13 2 7 1 9 15 1 15 13 2 16 13 2
31 3 1 0 9 9 2 13 1 9 1 15 9 13 9 2 9 9 15 2 16 1 15 9 15 0 13 1 15 9 13 2
27 1 3 9 4 13 1 9 1 9 0 2 0 13 15 13 2 7 0 1 9 13 1 9 1 9 0 2
16 1 0 7 9 9 2 13 1 9 9 9 3 1 9 13 2
27 16 3 9 13 0 2 0 13 15 13 9 13 2 3 3 0 13 15 13 2 15 16 1 0 13 13 2
32 7 1 13 13 3 9 13 12 3 1 9 0 1 10 9 7 13 0 9 1 12 9 13 13 2 16 0 9 1 13 9 2
17 3 10 13 16 12 9 2 15 13 9 1 9 15 1 9 12 2
86 9 7 15 13 1 9 13 7 13 1 9 7 13 2 3 3 13 1 9 13 2 7 3 1 9 15 9 7 13 9 9 2 15 7 15 9 13 9 1 13 15 9 9 2 16 9 16 1 15 13 9 2 7 13 9 13 1 0 9 2 7 1 0 9 13 0 7 9 2 0 9 16 13 9 9 1 13 2 16 9 3 13 1 0 0 2
33 13 3 2 1 15 16 13 9 2 16 1 13 13 9 1 13 2 7 1 9 13 9 1 13 2 16 13 15 13 1 0 9 2
28 7 16 3 9 13 1 13 1 9 9 1 15 13 0 0 9 0 2 13 9 9 2 16 1 9 13 3 2
50 16 0 3 13 0 0 9 15 9 2 3 13 9 9 2 7 9 0 2 16 13 1 9 9 2 15 13 1 9 13 0 2 3 3 13 1 0 9 0 2 7 3 3 13 9 0 2 7 0 2
10 0 13 1 9 9 9 1 9 0 2
13 3 0 9 13 1 9 9 1 13 9 9 0 2
7 3 3 13 1 9 9 2
22 3 9 13 1 9 3 13 0 0 9 2 15 13 9 9 2 16 13 0 9 13 2
11 3 3 9 1 9 0 13 13 9 9 2
29 1 13 3 13 16 9 15 13 1 9 13 2 1 15 13 1 9 9 3 2 1 15 0 1 9 9 7 0 2
38 16 3 15 9 1 15 1 9 13 9 2 13 0 0 7 1 9 7 1 0 2 13 9 0 1 9 13 2 16 1 15 15 13 1 9 7 3 2
45 16 7 3 13 0 0 7 0 13 2 3 13 9 1 9 13 16 1 9 9 15 13 1 13 2 16 1 15 15 13 3 1 10 9 7 1 9 9 2 7 1 9 15 0 2
13 3 3 13 3 7 1 9 2 7 16 1 0 2
10 1 9 7 0 13 1 9 9 0 2
11 12 3 9 2 16 13 0 1 9 9 2
15 7 3 1 15 2 15 9 13 9 1 9 7 1 9 2
17 9 3 1 3 13 1 3 9 13 2 3 1 0 7 1 0 2
20 1 9 3 0 2 9 9 13 9 1 10 9 2 1 15 9 13 15 13 2
21 3 13 16 1 9 9 13 9 0 1 9 2 16 0 1 9 9 13 1 0 2
49 1 9 7 0 2 3 9 13 1 13 1 9 3 13 9 2 16 3 3 3 13 1 13 15 7 15 15 13 1 9 3 13 9 2 16 9 3 0 1 15 7 15 13 13 2 7 0 9 2
14 15 0 9 13 1 9 9 1 16 13 0 1 9 2
24 7 15 13 9 3 0 2 7 13 2 16 13 0 13 16 9 13 0 16 13 13 9 9 2
8 16 3 13 0 9 3 13 2
15 1 13 7 13 13 16 3 13 0 9 13 1 0 13 2
26 16 3 9 9 2 7 15 12 9 2 0 13 13 2 13 16 9 15 13 1 15 2 7 1 15 2
8 1 15 3 15 13 3 13 2
13 13 4 3 1 16 10 9 13 13 1 0 9 2
28 15 7 3 13 9 1 15 2 0 13 16 9 13 1 15 13 2 16 15 0 13 13 2 0 13 3 13 2
36 7 3 15 1 15 13 16 13 13 2 1 15 13 16 3 13 13 3 9 2 7 1 13 2 16 3 13 3 9 2 7 3 16 13 9 2
30 16 7 15 9 9 13 1 15 2 13 16 13 1 15 9 15 13 0 2 16 15 13 0 9 2 13 9 1 15 2
10 9 7 0 13 7 0 2 7 9 2
18 1 0 0 13 16 9 0 13 13 2 1 15 16 9 0 13 13 2
10 1 9 3 9 9 1 9 0 13 2
18 16 3 9 3 0 13 13 1 9 9 2 7 9 0 13 13 0 2
16 9 7 3 13 1 15 9 1 9 9 2 16 1 13 4 2
13 3 13 3 0 0 9 13 9 13 1 9 0 2
8 0 7 9 13 1 9 0 2
40 15 3 15 13 1 9 2 9 1 9 3 13 16 1 16 9 1 15 7 3 13 13 2 16 9 9 1 9 2 7 3 3 3 13 2 16 9 1 9 2
26 9 7 0 9 2 1 15 9 1 9 13 2 3 13 15 13 16 10 9 2 16 1 0 13 4 2
31 15 3 1 9 3 13 2 7 3 1 13 2 1 13 1 15 13 2 7 3 1 3 13 2 1 13 1 15 9 0 2
6 15 10 1 13 4 2
8 3 13 3 9 13 0 0 2
9 7 3 0 13 13 9 3 13 2
2 3 2
19 15 13 1 9 2 3 13 0 0 2 16 9 16 9 15 13 13 0 2
32 9 7 3 1 9 9 2 7 1 9 13 9 1 9 2 16 13 4 2 7 1 9 13 9 13 2 16 1 0 13 4 2
8 3 3 13 0 0 9 13 2
8 7 3 0 13 15 3 13 2
2 0 2
40 13 4 1 16 9 3 13 15 9 15 13 1 15 2 3 1 15 13 7 1 9 13 2 16 9 13 1 9 7 13 1 9 2 7 15 13 13 15 13 2
13 7 15 9 13 9 2 1 16 9 13 15 13 2
29 7 3 13 0 16 9 13 9 3 13 2 1 3 3 13 0 9 13 16 9 13 3 2 16 1 0 13 4 2
9 3 3 13 0 16 9 3 13 2
2 3 2
15 1 9 1 9 3 13 15 1 9 16 1 9 15 9 2
20 1 15 7 9 9 9 13 2 16 0 0 9 9 13 2 16 1 13 4 2
8 3 3 1 9 9 9 13 2
16 7 3 0 13 2 16 9 0 13 2 16 9 1 0 13 2
2 3 2
40 13 4 1 16 0 9 1 9 13 3 13 1 9 1 0 9 15 1 15 0 13 13 2 3 9 2 7 1 9 1 15 9 2 15 3 13 1 15 13 2
19 9 7 9 1 15 15 3 13 1 15 0 13 2 3 13 15 3 13 2
10 13 3 2 16 15 13 2 16 13 2
18 3 3 0 13 16 3 13 4 2 16 15 13 3 13 1 15 0 2
7 15 3 13 9 3 13 2
10 9 13 13 9 9 1 9 9 13 2
34 7 16 0 9 13 16 9 3 7 1 9 13 2 7 15 13 13 4 2 13 9 15 13 2 16 13 16 3 1 9 13 9 9 2
12 0 2 7 2 13 9 15 13 1 9 9 2
8 0 2 15 13 1 9 9 2
17 0 2 15 13 1 9 9 9 2 1 15 13 1 0 13 13 2
13 1 9 7 9 2 1 9 9 13 13 9 3 2
14 10 9 15 3 3 13 2 13 1 15 7 1 9 2
30 1 15 3 2 16 9 15 3 3 13 2 13 13 7 16 1 0 13 2 7 16 1 0 13 2 16 13 0 0 2
52 1 9 7 2 16 9 9 13 1 0 13 9 15 0 9 13 1 15 2 7 1 0 2 16 2 1 9 13 9 13 2 13 13 2 7 1 0 2 16 1 1 0 13 9 13 1 15 9 1 0 13 2
17 9 7 3 13 7 1 15 7 1 9 2 16 1 0 13 4 2
7 9 3 3 15 9 13 2
10 1 10 7 9 9 13 1 9 13 2
5 3 3 9 13 2
2 3 2
9 9 13 1 9 13 1 9 15 2
6 7 9 9 13 0 2
23 15 13 1 9 9 9 9 2 7 13 16 13 1 9 1 15 0 9 2 15 13 0 2
9 3 9 1 9 13 1 0 13 2
2 0 2
9 13 9 13 2 0 13 9 13 2
26 16 3 3 2 13 9 2 3 0 13 9 13 2 0 3 13 2 9 13 2 9 13 7 3 13 2
9 9 3 9 1 9 13 0 3 2
12 15 7 13 0 2 13 15 15 13 1 9 2
13 13 3 13 15 9 15 13 16 9 13 1 9 2
8 7 3 0 9 3 13 0 2
8 7 9 13 9 0 9 9 2
14 15 3 13 9 2 7 3 1 9 15 1 9 13 2
6 15 3 13 13 9 2
5 15 13 13 0 2
18 13 3 0 16 2 1 9 1 0 13 2 16 9 3 13 1 0 2
2 3 2
21 9 1 9 3 13 10 13 13 1 15 13 16 1 15 1 0 13 15 3 13 2
50 7 15 3 13 1 15 9 2 16 1 13 9 9 1 13 2 7 9 15 13 9 2 3 0 13 1 9 2 16 1 13 9 15 1 15 9 13 2 7 3 1 13 9 15 9 0 15 3 13 2
33 16 3 9 13 0 2 3 9 13 2 16 13 9 1 15 2 16 1 9 9 3 13 9 9 2 16 13 9 9 9 13 9 2
39 7 1 15 13 16 2 1 15 13 15 13 7 3 3 13 2 13 16 7 15 13 1 9 9 2 15 13 13 2 7 16 9 3 13 0 1 15 13 2
14 13 7 9 9 13 2 16 13 15 0 13 10 9 2
28 9 7 0 13 2 16 15 3 13 13 15 0 2 7 13 15 9 15 3 13 2 7 16 13 9 15 13 2
16 13 7 16 15 9 3 13 16 13 2 1 0 13 16 13 2
9 3 3 0 9 9 15 13 13 2
34 7 15 9 7 9 9 15 13 13 2 7 15 15 13 13 1 0 9 9 2 1 15 15 13 0 16 15 0 2 16 1 13 4 2
11 0 3 13 16 1 0 9 1 9 13 2
2 3 2
14 9 1 9 3 13 12 15 16 1 9 12 1 15 2
12 7 16 15 13 9 2 3 13 2 13 9 2
13 16 3 15 13 9 2 3 13 9 12 1 15 2
19 7 1 15 1 9 1 15 15 13 0 15 13 9 2 16 7 1 9 2
7 15 3 9 13 9 9 2
11 3 9 7 1 3 9 15 13 13 9 2
9 12 3 3 9 3 13 15 0 2
11 7 1 15 9 9 15 13 16 9 9 2
21 1 15 7 3 13 13 15 9 9 2 16 1 12 3 13 15 13 16 1 15 2
18 0 7 1 9 2 15 15 13 0 7 0 2 16 1 0 13 4 2
15 13 3 16 9 9 0 15 13 1 13 9 1 15 9 2
19 7 3 9 10 13 1 15 16 3 9 1 9 15 13 2 7 8 3 2
26 13 7 16 3 13 9 15 1 15 16 3 9 1 9 15 0 13 2 1 13 9 9 15 4 13 2
13 13 3 1 9 2 16 13 2 16 9 3 13 2
2 3 2
19 15 15 13 1 9 2 9 13 1 9 2 7 0 1 15 15 9 13 2
30 13 3 16 2 9 15 9 15 13 2 15 15 13 1 9 15 9 15 13 7 13 2 16 13 0 9 15 1 9 2
19 9 7 9 1 0 9 13 13 0 9 2 15 0 13 13 0 9 9 2
34 1 3 9 0 1 15 9 15 9 15 13 1 15 7 1 9 1 0 9 13 16 15 9 9 1 9 13 1 0 9 1 15 9 2
28 3 3 13 13 16 15 0 9 15 13 1 9 2 16 3 13 3 13 1 15 13 9 2 1 15 13 13 2
2 3 2
43 1 9 0 9 13 2 3 15 9 13 16 10 1 9 13 1 9 15 2 16 15 15 1 9 13 2 7 16 9 13 16 15 13 16 0 13 2 1 15 15 9 13 2
20 1 7 10 9 9 13 16 13 9 2 1 16 0 13 2 3 9 9 13 2
9 3 7 9 0 9 13 0 9 2
6 9 7 0 0 13 2
15 15 3 13 16 15 1 0 13 2 3 15 13 9 3 2
15 15 3 13 1 0 9 13 2 16 9 15 1 0 13 2
15 15 3 13 1 9 9 13 1 15 13 16 9 3 13 2
10 9 13 13 9 9 13 1 9 9 2
15 13 7 7 15 2 1 9 9 13 2 15 15 13 13 2
15 15 3 3 13 9 1 3 13 2 0 13 15 3 13 2
14 15 7 13 1 9 1 15 3 13 9 1 3 13 2
17 3 3 13 13 9 1 3 13 16 1 15 15 13 9 9 9 2
19 9 3 1 13 7 3 13 13 9 1 9 7 9 2 15 9 13 9 2
16 9 0 3 13 9 0 2 1 0 13 9 13 1 10 9 2
46 7 15 9 13 1 15 3 13 9 9 9 2 7 16 3 3 13 9 2 16 9 0 2 16 1 13 2 7 3 13 0 2 16 9 0 2 15 15 9 13 2 15 0 3 13 2
8 15 3 9 0 13 3 13 2
7 3 15 0 13 3 13 2
2 3 2
23 15 9 3 13 1 9 15 13 10 9 13 2 16 1 9 2 16 1 15 15 0 13 2
26 7 15 9 13 15 13 9 13 3 1 15 13 9 2 7 1 3 13 2 16 9 0 7 0 9 2
9 0 3 13 2 1 0 3 13 2
8 13 3 16 15 13 3 13 2
9 15 7 13 13 2 3 3 13 2
8 15 3 3 13 16 13 13 2
2 3 2
32 16 15 1 0 13 13 2 13 16 13 2 7 13 2 7 15 2 15 15 13 3 16 13 9 2 16 0 16 3 13 9 2
15 13 3 9 7 9 15 13 1 13 1 16 13 13 9 2
13 9 7 0 3 13 1 9 15 7 15 3 0 2
11 15 7 15 15 13 3 7 0 2 13 2
19 3 13 2 1 9 15 1 0 13 2 15 9 13 1 0 7 1 13 2
16 13 3 16 15 9 7 13 0 2 7 13 15 9 1 15 2
5 9 3 3 13 2
4 3 7 0 2
6 7 3 9 3 13 2
12 9 3 3 0 13 2 16 1 0 13 4 2
2 3 2
23 10 9 2 15 13 15 0 2 13 13 9 0 1 9 2 15 3 13 0 13 1 9 2
8 0 13 7 9 9 0 13 2
9 13 3 16 9 0 9 13 0 2
2 3 2
15 16 9 13 0 2 13 9 13 0 2 1 13 9 9 2
13 7 1 13 0 13 0 2 1 9 13 9 0 2
6 7 9 13 13 0 2
18 3 3 13 13 13 9 16 13 3 2 16 7 9 13 13 1 9 2
10 3 7 3 13 9 13 7 9 0 2
7 15 3 13 9 15 3 2
13 7 3 15 3 13 13 1 15 9 0 7 0 2
9 7 3 15 13 13 0 7 0 2
14 13 3 16 0 2 15 13 9 13 2 13 1 0 2
2 3 2
6 13 7 13 7 13 2
14 16 3 1 9 15 13 15 9 2 13 15 13 3 2
5 9 7 13 3 2
37 3 2 16 9 3 3 13 2 13 13 0 3 9 15 16 9 2 7 0 2 16 3 13 3 0 2 13 16 3 9 15 13 0 1 9 15 2
13 0 7 7 0 3 13 13 1 9 16 9 13 2
8 3 9 0 7 0 9 13 2
14 7 3 13 9 13 16 13 2 7 0 13 16 13 2
6 13 3 9 13 0 2
12 9 7 13 9 2 15 1 9 13 3 13 2
23 9 7 15 3 13 9 2 15 13 1 9 2 1 13 3 0 2 16 1 0 13 4 2
8 13 3 15 9 13 0 13 2
2 0 2
15 0 9 3 15 13 16 15 15 13 2 13 16 15 13 2
10 16 15 13 9 13 2 13 9 13 2
9 13 3 10 0 13 0 15 13 2
15 7 0 13 1 15 15 13 15 9 2 9 3 13 3 2
23 13 3 15 13 9 15 13 13 0 2 13 7 9 0 2 7 3 3 1 15 15 13 2
33 16 3 15 1 15 9 13 10 9 2 13 13 3 2 16 13 4 2 13 16 13 9 2 7 10 15 1 15 13 2 13 0 2
7 15 7 9 3 13 9 2
8 3 13 15 1 9 13 0 2
15 15 3 7 3 9 13 13 1 9 9 16 9 13 3 2
9 9 1 13 9 9 1 9 9 2
15 13 3 13 15 9 2 1 9 15 9 2 1 15 13 2
13 15 3 1 10 0 13 2 0 13 0 13 0 2
20 0 3 9 9 15 9 13 2 16 7 0 9 1 0 0 1 9 9 13 2
11 9 7 1 9 13 2 16 1 9 9 2
29 15 7 13 1 9 2 3 13 13 3 7 1 10 2 16 9 15 1 9 1 10 9 13 2 3 13 13 0 2
14 3 9 15 1 10 1 9 13 2 3 13 13 0 2
11 0 7 9 13 10 9 1 15 15 13 2
6 13 3 15 13 0 2
12 16 3 15 4 13 2 13 1 15 4 13 2
14 15 16 3 13 4 2 13 3 7 15 1 15 13 2
21 3 13 7 15 1 0 13 2 16 3 15 9 13 2 1 3 13 0 0 13 2
11 13 3 13 1 15 0 15 3 4 13 2
12 10 7 9 15 3 3 13 2 13 4 13 2
12 3 13 15 1 15 0 10 13 2 13 0 2
21 15 7 3 13 9 2 16 15 3 13 13 9 15 9 2 16 1 0 13 4 2
13 13 3 16 15 1 9 13 0 2 3 0 9 2
2 0 2
17 16 15 3 15 13 15 9 3 7 0 2 13 15 13 0 13 2
14 15 3 13 13 2 3 15 9 15 3 7 0 13 2
17 10 7 15 1 0 13 13 2 3 15 9 15 13 3 7 0 2
10 13 3 15 1 15 9 13 7 9 2
10 10 7 9 7 9 1 15 9 13 2
5 13 3 9 0 2
26 1 7 9 13 0 15 15 13 1 9 2 1 1 15 13 9 2 13 1 15 13 13 15 9 0 2
24 7 1 15 3 13 0 1 0 13 2 13 13 1 15 0 9 3 1 0 13 7 3 13 2
2 3 2
15 10 15 1 0 13 13 2 16 13 2 0 13 15 13 2
14 16 3 3 2 0 13 15 13 2 7 0 3 13 2
11 7 3 3 13 3 9 7 3 13 13 2
11 7 15 13 0 13 2 13 9 9 13 2
12 13 3 1 15 1 0 13 13 9 9 13 2
21 7 1 15 1 0 13 3 13 2 13 13 15 0 9 15 3 13 13 1 0 2
2 3 2
7 15 9 13 13 16 13 2
7 1 15 3 13 16 13 2
8 3 3 13 2 16 3 13 2
12 7 16 13 2 13 15 13 15 13 9 9 2
13 3 3 9 2 1 13 9 2 1 9 13 13 2
10 10 3 15 13 2 13 15 9 13 2
19 7 1 15 1 0 13 3 13 2 13 0 9 3 13 13 2 7 0 2
20 1 15 0 13 15 1 9 13 0 2 1 15 9 9 7 9 13 3 13 2
17 15 3 9 13 15 15 16 9 13 2 13 0 9 13 3 13 2
23 1 15 9 0 13 2 15 13 15 1 9 3 13 2 7 10 13 13 1 12 9 0 2
13 9 9 1 13 7 0 15 15 13 1 9 9 2
10 13 3 13 13 9 3 1 9 13 2
10 7 0 2 15 15 1 9 9 13 2
24 3 3 13 16 1 15 7 1 9 9 13 16 9 15 1 0 13 13 2 16 0 9 13 2
12 9 3 9 13 13 9 9 16 13 9 9 2
21 3 3 13 13 16 1 9 13 0 9 16 15 9 13 2 3 1 9 1 9 2
23 9 7 0 9 3 13 9 9 1 9 2 1 9 10 13 10 9 2 16 1 13 4 2
10 3 7 9 9 9 9 13 13 13 2
23 7 3 13 16 2 16 0 9 9 13 0 2 16 15 9 13 0 2 16 0 9 13 2
12 13 4 3 1 16 9 13 9 1 9 9 2
42 3 7 3 16 13 15 15 15 9 0 2 16 1 15 9 9 9 13 0 1 9 9 7 9 2 16 1 13 13 4 2 7 13 16 10 13 7 13 13 10 13 2
14 9 7 1 9 7 9 13 1 9 9 7 9 9 2
17 16 7 1 9 13 9 13 15 15 9 2 3 7 13 15 9 2
22 3 3 0 9 13 16 15 15 13 2 7 16 3 13 2 16 9 16 3 9 13 2
27 3 2 16 15 13 1 15 13 0 1 9 13 2 13 1 0 9 1 0 9 2 15 9 1 0 13 2
23 15 3 13 13 9 9 1 0 13 2 9 7 3 1 0 2 7 3 1 1 0 13 2
34 1 15 3 13 16 2 16 9 13 0 9 9 9 1 9 2 3 3 13 16 15 9 0 13 2 15 13 0 2 16 0 9 13 2
16 13 3 9 0 2 13 15 9 2 3 7 9 0 1 9 2
13 15 3 13 1 9 9 2 7 16 0 3 13 2
12 0 7 9 9 13 16 13 15 15 9 13 2
20 16 7 15 15 13 16 9 13 2 3 13 9 0 9 2 7 0 1 15 2
19 9 7 2 16 13 4 2 16 13 15 13 15 2 3 13 15 13 3 2
26 3 3 13 2 1 15 16 9 13 0 9 2 16 9 13 16 9 13 2 7 16 9 9 13 13 2
22 1 15 7 15 1 9 0 13 13 2 1 13 2 16 9 9 13 1 16 15 13 2
8 3 1 13 9 13 13 9 2
16 9 7 13 2 3 1 9 10 9 2 7 1 9 10 13 2
24 7 3 2 16 9 0 9 13 9 9 2 16 13 0 2 3 9 9 1 9 13 9 13 2
24 1 15 3 13 16 0 9 3 13 9 2 16 3 3 13 2 9 13 2 16 0 9 13 2
17 3 1 9 0 13 3 0 16 15 9 13 2 7 16 3 13 2
23 15 3 13 15 13 3 9 13 2 3 13 2 16 3 13 9 13 16 9 1 0 13 2
20 3 13 7 1 15 9 9 9 15 9 15 9 13 2 16 1 0 9 13 2
8 3 15 9 3 13 7 9 2
34 9 7 9 2 15 13 9 2 3 13 9 2 7 13 0 3 2 3 13 0 7 0 2 1 9 13 0 2 16 1 0 13 4 2
52 3 13 3 13 9 15 9 1 15 0 13 1 15 13 9 2 1 15 9 9 0 7 0 15 13 13 2 16 13 9 13 1 13 3 1 15 13 15 9 9 1 9 13 2 7 3 1 15 13 7 13 2
34 15 3 9 13 16 15 9 1 9 0 13 1 15 9 13 2 16 13 1 0 9 2 1 15 13 9 1 9 2 3 7 15 9 2
11 9 7 3 1 9 13 7 9 7 9 2
19 3 13 3 9 3 3 7 3 0 1 15 13 2 7 0 3 3 3 2
7 16 1 0 1 9 13 2
46 0 3 9 2 16 1 9 13 2 3 7 1 9 13 13 2 7 16 13 1 15 9 7 9 2 1 15 13 2 13 13 9 3 3 1 15 9 7 1 15 9 13 16 1 15 2
31 1 15 7 9 2 1 15 3 13 9 2 7 1 15 0 9 10 13 2 3 13 9 13 3 3 7 3 3 13 4 2
17 15 9 16 15 13 13 2 13 1 9 2 16 13 0 1 9 2
56 7 0 1 9 15 9 2 1 15 3 13 9 2 7 1 15 3 9 13 2 3 13 13 9 3 3 7 3 0 2 16 1 15 13 1 13 9 9 2 7 0 3 3 3 2 7 3 1 3 9 2 7 1 15 9 2
23 1 15 7 13 2 0 9 13 1 9 9 2 15 0 13 13 9 1 15 15 9 13 2
11 9 7 0 9 3 13 13 16 15 9 2
32 3 7 13 1 15 9 13 1 9 2 16 9 13 1 9 9 2 1 9 15 13 0 7 0 2 3 16 15 15 13 13 2
11 7 3 13 13 16 1 15 9 9 13 2
16 7 3 13 1 15 9 13 15 2 16 9 13 16 13 9 2
6 15 3 13 10 9 2
13 13 3 16 13 1 9 16 9 13 1 9 9 2
44 1 13 3 9 3 1 9 2 0 9 9 1 9 3 13 13 16 9 9 0 2 7 3 13 13 9 9 1 9 15 13 1 9 2 16 15 13 9 15 13 13 1 9 2
19 3 1 15 16 9 0 15 13 1 9 2 3 13 13 16 9 13 0 2
36 7 13 0 9 0 3 13 2 1 15 16 3 13 13 1 9 2 16 0 9 13 13 2 7 13 13 1 9 1 15 16 13 3 3 13 2
17 10 3 9 13 9 1 9 10 9 2 13 1 15 13 10 9 2
20 3 3 0 9 13 13 1 10 9 9 9 13 2 16 10 9 0 9 13 2
36 3 7 13 13 15 9 1 9 9 2 16 9 0 10 9 13 2 16 3 13 1 0 9 0 9 13 2 7 16 13 13 1 15 15 13 2
16 9 7 0 9 1 9 1 15 0 13 16 9 3 3 13 2
43 1 15 3 13 13 16 10 15 1 15 15 13 10 9 9 2 7 16 9 15 3 13 1 3 9 13 2 16 9 1 9 0 2 7 1 13 16 13 9 13 7 13 2
9 15 0 15 13 2 9 9 13 2
14 3 3 1 9 9 15 13 15 9 9 15 13 13 2
9 9 9 15 13 1 9 9 13 2
18 0 3 7 1 9 9 13 15 15 15 1 15 9 13 1 9 13 2
26 9 3 13 15 1 9 13 2 1 15 0 9 1 15 13 2 13 9 9 2 16 1 13 4 13 2
19 9 7 9 3 13 15 15 15 13 9 2 3 13 2 16 1 13 4 2
26 16 3 9 9 2 1 15 16 13 9 1 3 9 2 13 9 1 9 2 15 3 9 13 15 9 2
16 3 2 9 15 3 1 9 13 2 15 9 9 3 13 13 2
18 3 7 13 13 0 9 3 13 2 1 9 15 13 1 9 9 15 2
16 0 3 9 13 3 2 1 15 13 0 9 2 13 9 9 2
18 3 2 1 1 9 9 9 13 2 15 9 9 9 0 13 3 13 2
11 9 3 9 3 13 15 13 9 13 13 2
16 3 3 13 16 1 9 9 13 13 13 16 0 13 3 0 2
16 16 7 0 13 15 1 15 13 1 0 2 13 16 7 13 2
13 3 9 9 9 9 0 13 1 9 3 3 13 2
21 0 3 9 0 9 1 9 9 2 1 15 0 9 13 2 13 0 9 3 13 2
23 3 9 3 13 15 9 16 1 9 0 3 1 9 13 2 3 7 1 1 9 9 13 2
13 3 7 0 13 13 9 0 13 2 1 13 13 2
15 9 3 0 2 1 9 13 2 9 9 3 13 16 13 2
43 1 3 0 7 0 7 9 9 13 0 7 0 7 9 9 2 1 9 9 2 13 16 15 9 13 9 0 7 9 13 16 15 13 1 9 13 9 7 9 0 9 9 2
29 3 13 3 10 9 3 13 2 16 10 9 1 9 13 13 0 1 0 7 0 1 9 2 15 13 13 9 0 2
20 13 7 9 3 13 0 2 13 13 0 9 9 13 9 0 7 15 13 9 2
63 7 13 9 9 16 13 1 15 15 3 9 7 3 9 1 15 16 9 2 1 15 13 13 15 9 7 3 9 2 13 13 2 7 3 13 2 16 3 1 9 15 0 2 15 3 3 13 13 7 13 2 13 15 13 16 9 9 3 7 3 16 9 2
11 15 3 10 9 13 0 2 15 13 0 2
32 16 7 0 13 3 9 9 16 15 9 16 9 13 2 3 13 15 13 16 13 9 13 16 13 3 13 2 16 0 9 13 2
21 3 0 15 13 16 9 13 2 3 13 15 9 9 1 9 2 7 0 1 9 2
23 1 3 13 16 9 13 9 1 3 9 2 13 16 3 13 15 9 9 1 15 3 13 2
33 16 2 1 13 16 1 9 15 13 2 3 13 16 15 9 13 1 9 15 13 13 1 9 9 2 7 16 3 13 9 15 0 2
10 3 7 9 13 9 15 9 13 13 2
22 9 15 2 16 3 13 13 9 9 0 2 16 13 1 12 8 2 3 7 9 0 2
25 9 7 9 15 13 13 3 9 13 2 1 15 0 9 13 2 13 9 9 15 13 9 1 9 2
26 3 3 13 15 9 13 3 2 16 9 9 0 2 1 15 13 9 10 9 2 16 1 0 13 4 2
14 13 3 16 9 1 9 13 3 13 1 9 9 13 2
9 9 9 15 13 1 9 9 9 2
17 13 7 13 16 7 1 9 9 9 15 9 13 13 13 1 15 2
25 0 3 9 9 13 1 15 15 13 2 1 15 0 9 13 2 9 13 1 15 13 15 15 13 2
22 16 3 10 10 9 1 9 13 2 15 0 13 2 1 0 9 1 0 9 0 13 2
20 3 9 9 13 0 9 9 3 13 2 13 15 7 15 9 7 15 9 13 2
49 7 3 0 2 3 0 16 13 13 9 13 2 13 9 13 0 1 15 0 9 2 16 0 2 0 2 7 3 2 13 1 13 13 15 13 16 13 2 1 15 16 1 9 1 9 15 13 13 2
39 0 0 2 3 0 2 9 9 13 2 1 13 9 1 9 13 2 13 16 3 13 15 13 1 9 1 9 16 1 9 2 7 1 15 1 9 1 9 2
16 15 7 13 2 15 13 9 1 15 9 2 13 9 9 0 2
19 15 3 13 16 13 15 9 2 16 9 7 9 2 3 7 16 13 0 2
11 9 3 0 13 2 15 1 15 9 13 2
28 0 7 1 9 9 13 2 13 1 0 15 9 13 1 12 0 9 9 2 16 1 9 15 13 1 13 13 2
18 1 15 7 9 15 9 1 9 3 13 0 13 15 1 15 15 13 2
8 3 3 13 15 9 13 9 2
18 7 15 3 9 3 13 0 0 2 15 13 0 9 1 15 15 13 2
46 7 2 16 15 15 13 2 3 0 9 9 15 13 13 2 1 9 9 9 7 9 13 2 1 15 7 15 9 9 1 12 0 9 13 3 13 9 12 9 1 15 2 16 13 4 2
29 1 15 7 1 0 9 13 3 9 9 13 2 7 1 9 0 2 15 13 9 0 7 15 15 13 13 1 9 2
26 15 3 1 15 9 3 1 15 9 9 9 13 2 16 13 15 13 15 9 7 9 1 15 9 13 2
17 1 15 13 16 7 0 9 1 9 13 2 15 1 9 9 13 2
19 3 9 9 13 3 13 16 1 9 2 16 13 13 13 9 1 3 9 2
30 9 15 15 1 15 13 13 3 15 15 3 9 3 13 2 1 15 0 16 12 15 13 1 15 2 16 9 1 9 2
10 7 9 9 13 1 15 15 13 13 2
29 3 15 15 9 13 2 3 15 13 15 9 2 16 13 13 16 2 16 13 13 2 15 9 15 13 3 7 0 2
21 1 15 3 13 16 3 13 15 9 0 13 9 15 9 13 2 16 0 9 13 2
22 15 3 13 0 1 15 15 1 9 13 9 13 2 15 16 9 13 9 13 1 9 2
20 0 7 13 9 13 4 2 16 13 2 1 9 9 2 1 15 7 13 13 2
11 7 1 9 9 2 1 15 15 9 13 2
17 15 3 0 1 15 9 13 2 16 13 1 9 2 1 12 8 2
22 15 3 9 15 13 9 2 3 13 15 9 15 13 9 7 9 2 16 0 13 9 2
24 7 3 13 16 3 13 0 13 2 7 1 13 16 13 0 13 16 13 2 3 15 9 13 2
29 1 15 7 15 1 9 13 2 13 0 13 0 1 15 0 9 2 1 15 9 2 1 12 8 2 15 13 9 2
12 13 3 1 15 16 7 0 9 1 13 13 2
21 3 13 3 3 13 1 9 9 1 15 15 1 9 13 2 1 15 13 9 13 2
16 1 15 7 15 3 13 1 9 2 3 13 0 13 16 9 2
13 3 3 0 13 16 15 13 13 9 3 3 13 2
5 15 9 0 13 2
3 8 12 2
8 1 9 13 9 9 7 9 2
7 7 8 12 1 9 13 2
7 16 15 13 1 9 8 2
10 9 15 15 13 13 9 3 13 0 2
18 13 7 15 9 1 15 13 1 13 9 3 3 13 2 13 1 15 2
9 9 3 13 10 9 9 4 13 2
12 9 7 13 9 13 15 15 1 9 9 13 2
2 3 2
26 1 15 9 1 9 4 13 2 3 13 13 13 4 1 15 9 2 7 3 13 16 4 13 1 15 2
10 7 1 13 16 13 9 1 3 9 2
2 3 2
6 16 0 3 13 13 2
19 16 7 9 3 13 2 4 3 0 13 2 16 15 13 4 2 13 4 2
14 13 7 0 9 7 9 9 13 2 16 9 3 13 2
2 3 2
17 13 16 0 13 9 2 1 1 9 7 9 13 3 1 0 13 2
2 0 2
22 13 16 1 9 13 13 13 1 0 2 16 9 13 3 2 15 13 13 9 3 13 2
15 3 9 9 13 9 2 7 15 15 2 7 3 1 0 2
2 3 2
12 13 16 13 0 2 3 0 9 13 9 0 2
35 15 7 9 16 3 3 1 9 13 2 16 9 13 2 13 13 0 2 16 13 9 0 1 0 9 13 2 7 3 0 1 0 9 9 2
15 7 3 13 13 13 15 13 15 1 15 15 9 9 13 2
35 15 3 0 13 2 9 1 9 13 9 15 1 10 9 13 2 0 13 1 15 15 13 15 1 9 2 16 9 3 13 16 1 9 9 2
10 9 7 0 13 13 3 1 9 13 2
26 1 15 7 15 1 9 13 2 15 3 13 0 2 16 3 16 9 13 1 9 13 2 13 10 0 2
9 15 3 0 13 2 3 13 0 2
37 15 3 15 13 1 15 15 13 2 0 15 13 13 1 15 3 13 2 13 3 1 15 13 2 3 7 15 16 13 1 15 2 16 1 9 0 2
11 1 15 13 3 13 16 13 1 3 13 2
9 15 3 0 13 2 3 13 13 2
24 3 0 2 16 3 13 3 1 9 2 13 3 13 1 9 2 16 3 15 0 13 13 13 2
11 15 3 9 13 13 13 2 16 13 13 2
15 1 10 7 3 2 16 9 3 13 2 3 13 13 0 2
11 7 3 7 9 2 15 3 13 12 0 2
8 15 3 0 13 2 0 13 2
13 3 15 13 0 1 15 9 9 13 15 13 13 2
22 1 15 7 16 13 9 0 2 13 16 13 0 1 9 1 2 7 13 1 9 1 2
6 3 0 13 9 13 2
8 15 3 0 13 2 3 13 2
27 16 9 13 1 0 13 13 0 2 1 9 2 1 9 3 13 2 16 13 9 13 1 9 0 3 13 2
15 7 3 13 9 1 15 0 2 16 15 9 1 13 13 2
19 1 9 7 3 3 13 2 15 3 13 0 2 1 15 15 13 9 0 2
6 15 7 9 13 9 2
12 13 3 9 9 16 13 15 9 7 3 9 2
15 3 7 13 9 2 16 13 9 2 16 4 13 1 9 2
6 13 3 16 4 13 2
8 15 7 1 9 13 0 13 2
12 7 3 9 3 13 0 0 2 16 0 13 2
14 15 3 9 9 13 13 3 0 9 3 13 1 9 2
25 15 0 16 1 10 9 3 13 16 9 13 2 7 13 2 1 15 2 7 3 0 2 1 15 2
18 15 7 13 9 1 9 2 13 16 15 9 1 15 9 1 9 13 2
18 15 0 1 9 3 13 16 13 15 0 9 1 15 15 9 3 13 2
17 13 7 0 13 1 15 13 1 9 0 9 2 16 1 13 4 2
15 9 3 0 9 1 9 9 13 15 9 16 1 13 13 2
18 0 7 13 0 9 7 9 1 15 16 9 15 1 15 3 3 13 2
20 1 15 3 13 0 16 9 15 1 15 1 15 9 13 2 16 3 3 13 2
18 13 3 16 3 13 1 9 9 2 7 16 9 10 13 0 1 13 2
14 15 3 13 13 0 9 2 16 9 13 9 9 13 2
14 1 15 7 15 13 4 2 13 13 0 9 0 9 2
6 15 15 13 9 0 2
29 15 9 9 0 2 1 15 1 15 9 9 13 13 2 7 1 9 2 7 1 15 9 2 7 3 9 7 9 2
10 1 10 3 15 13 15 1 9 0 2
5 15 9 0 13 2
8 8 9 9 3 13 1 9 2
19 13 7 15 15 1 9 9 13 2 13 13 15 15 13 13 1 9 9 2
13 1 15 0 13 13 16 9 9 3 13 1 9 2
11 9 3 3 13 16 1 0 15 15 13 2
14 15 3 13 1 9 7 3 2 3 13 13 1 9 2
27 13 4 7 1 15 9 13 4 1 15 9 3 13 9 1 3 13 2 16 13 9 0 2 7 1 9 2
9 9 3 15 0 13 13 1 9 2
9 13 7 1 10 9 1 3 13 2
8 15 3 9 3 13 1 9 2
2 0 2
29 1 9 13 3 1 0 15 15 13 2 9 7 3 9 13 9 2 3 7 9 2 15 3 13 9 9 1 12 2
20 15 15 9 13 1 9 2 3 13 9 2 7 9 15 15 9 13 1 9 2
7 9 7 9 13 1 9 2
7 0 7 15 9 1 9 2
20 9 3 9 1 9 3 13 13 1 9 2 7 9 15 9 9 13 13 0 2
2 3 2
24 1 9 13 9 7 9 9 0 2 16 13 4 2 1 15 9 13 13 9 15 1 9 13 2
15 13 4 7 1 16 0 9 9 1 9 3 13 1 9 2
9 1 15 3 9 9 13 3 13 2
34 13 7 16 0 9 9 1 9 13 2 1 0 13 1 9 13 15 7 1 3 13 2 7 1 15 12 0 2 16 3 13 1 9 2
11 3 13 3 0 16 9 9 13 1 9 2
2 3 2
11 9 1 15 0 13 15 15 13 1 9 2
21 16 3 0 13 1 9 1 15 13 2 9 13 13 0 13 1 9 1 9 0 2
10 9 7 9 13 0 9 7 9 9 2
11 13 3 9 7 9 13 9 13 7 13 2
27 9 7 7 9 9 13 1 9 1 15 7 13 2 1 13 7 3 7 1 0 1 10 9 15 9 13 2
23 3 7 9 9 13 1 9 1 15 7 13 2 3 1 9 2 15 13 9 1 9 0 2
2 0 2
16 15 9 13 1 13 1 9 7 9 2 9 13 1 13 13 2
21 15 7 9 9 9 13 9 2 15 13 9 1 9 7 9 2 16 1 13 13 2
27 7 1 9 10 9 15 13 13 2 16 3 13 1 10 9 2 1 10 9 13 0 2 16 1 13 4 2
12 13 3 16 9 0 13 1 9 13 7 13 2
6 3 13 3 1 9 2
10 9 3 13 13 15 1 9 9 13 2
11 9 7 0 13 1 9 7 9 9 15 2
8 3 13 3 9 9 1 9 2
2 3 2
14 15 15 13 0 7 0 1 9 2 13 9 9 15 2
20 7 9 7 9 0 13 1 9 9 15 1 3 2 15 1 9 13 3 13 2
15 1 15 3 9 0 1 10 9 13 2 15 13 0 15 2
13 15 3 9 9 0 7 9 15 13 9 9 0 2
8 3 13 3 9 9 1 9 2
39 15 7 9 0 9 13 2 16 13 8 12 2 16 2 1 0 13 2 1 9 13 9 9 7 9 2 13 2 13 9 9 1 9 2 7 3 1 15 2
26 16 3 0 9 9 2 7 3 9 9 1 9 13 13 2 3 1 9 2 7 3 9 7 9 0 2
3 3 13 2
11 13 9 10 15 13 2 7 13 3 0 2
22 1 15 7 13 9 0 0 13 9 0 0 7 12 2 1 15 10 13 9 7 9 2
25 15 3 0 13 13 9 9 15 1 0 13 2 3 1 15 13 9 13 2 7 1 9 0 9 2
58 0 3 13 9 9 7 9 13 0 9 0 2 3 0 9 15 9 7 13 9 2 9 7 9 2 1 15 9 2 15 13 13 0 2 1 9 13 13 2 13 13 9 1 9 2 1 12 13 0 9 2 3 9 2 9 7 9 2
7 3 13 9 9 13 0 2
7 15 1 13 13 13 0 2
9 16 9 3 13 0 9 9 9 2
18 1 15 7 0 13 16 9 9 3 13 1 9 9 16 1 0 9 2
18 1 9 3 15 13 13 13 16 0 2 15 16 9 1 0 0 13 2
16 1 15 16 12 3 13 2 15 16 1 0 13 0 13 13 2
13 3 7 13 15 0 13 2 7 0 13 9 9 2
11 13 4 7 16 9 9 3 13 1 9 2
13 13 3 16 3 13 1 9 9 16 1 0 9 2
2 3 2
16 15 15 13 1 9 9 2 3 13 1 9 16 1 0 9 2
24 9 3 13 0 13 1 13 16 9 2 16 9 3 13 9 9 16 1 16 4 13 1 9 2
21 3 2 16 15 9 13 9 9 7 9 9 2 3 13 1 9 16 1 9 0 2
27 7 1 15 13 16 15 15 13 1 9 16 1 9 0 2 13 1 9 9 2 16 9 7 15 9 9 2
7 9 7 13 1 9 9 2
5 15 1 15 13 2
21 9 3 13 15 0 1 9 2 7 16 3 15 13 2 15 13 1 9 1 9 2
22 9 3 3 13 9 9 16 0 9 2 7 3 1 0 9 3 13 16 13 15 9 2
9 9 7 9 1 9 13 1 9 2
13 9 3 9 3 13 1 9 9 16 1 0 9 2
2 0 2
16 9 9 3 13 13 1 9 16 1 15 15 1 9 13 13 2
32 0 7 13 1 3 13 1 9 15 3 13 1 13 9 13 2 16 13 1 9 0 2 15 3 13 0 2 16 15 9 13 2
11 3 3 13 13 0 9 9 9 9 9 2
2 3 2
12 15 13 10 9 9 13 2 13 9 10 9 2
18 15 3 1 15 13 9 1 15 13 12 1 15 0 7 1 15 13 2
18 7 16 9 15 9 13 9 9 9 2 13 13 9 1 15 13 13 2
25 13 7 16 9 15 13 9 1 15 2 1 15 16 1 13 4 10 15 15 13 2 1 9 13 2
8 3 15 13 9 9 1 9 2
11 3 3 0 9 9 9 13 13 9 9 2
2 3 2
23 1 10 9 13 1 9 2 3 13 0 1 0 2 7 1 0 2 7 0 13 1 9 2
16 10 7 9 13 1 9 1 9 13 2 16 1 1 13 13 2
13 13 3 1 9 0 1 0 2 7 3 1 0 2
13 9 7 0 13 9 2 1 13 9 7 9 15 2
20 3 3 13 15 9 9 1 15 9 2 7 3 15 9 13 16 13 15 9 2
27 3 3 9 9 1 9 2 15 13 1 9 2 13 1 9 2 7 3 9 4 13 0 16 0 9 13 2
27 1 15 7 13 9 9 13 0 9 0 2 1 9 3 13 1 12 13 2 15 3 9 13 9 9 13 2
12 7 15 15 13 0 9 0 1 9 9 13 2
9 16 9 9 3 13 1 9 9 2
18 1 13 3 13 13 16 9 9 9 3 13 9 2 7 3 9 9 2
24 16 3 0 9 1 15 13 9 9 2 13 13 1 3 2 13 16 15 9 13 15 12 9 2
9 3 0 3 13 16 1 15 12 2
12 7 3 15 13 13 0 9 7 12 9 9 2
20 16 0 0 9 3 13 1 3 13 2 9 15 1 9 9 13 13 1 9 2
6 9 3 9 13 0 2
6 15 0 1 13 4 2
2 3 2
15 1 0 9 3 13 3 13 9 13 2 16 9 1 9 2
10 0 3 2 16 3 2 3 13 12 2
20 9 7 13 13 13 9 1 3 3 0 2 1 16 1 0 12 1 15 13 2
15 0 13 3 16 9 9 3 13 13 1 9 9 3 13 2
2 0 2
14 15 13 9 10 9 2 3 13 13 0 9 9 9 2
16 7 16 0 9 1 0 13 2 0 13 16 13 9 10 9 2
19 13 3 9 13 2 1 10 9 13 1 12 0 9 2 16 1 13 4 2
16 15 7 13 9 13 15 7 9 15 1 15 2 16 13 4 2
11 3 13 3 13 0 9 9 9 9 9 2
2 3 2
40 16 9 9 13 1 9 7 9 0 9 2 0 15 13 2 15 7 0 13 2 1 9 9 7 9 2 3 16 10 9 13 1 0 9 2 9 7 1 0 2
9 9 3 7 9 13 1 10 9 2
10 3 13 7 13 12 0 9 10 9 2
25 1 3 15 15 13 1 15 2 13 1 15 15 13 1 15 2 13 0 0 9 13 1 15 9 2
12 1 15 7 13 15 15 1 9 10 15 13 2
7 15 3 9 3 13 0 2
5 15 7 13 0 2
14 10 3 15 13 2 16 13 9 2 0 13 13 0 2
9 9 3 10 15 13 7 13 13 2
11 9 7 13 2 16 1 13 15 10 9 2
7 9 7 13 15 10 13 2
19 3 13 3 9 1 9 13 1 12 0 9 15 12 13 0 7 15 0 2
2 3 2
7 10 9 13 16 13 9 2
9 16 0 13 9 2 15 9 13 2
10 9 0 10 2 16 3 2 0 13 2
10 10 3 9 2 16 3 2 0 13 2
13 16 15 3 1 15 0 13 2 3 13 13 9 2
17 16 7 13 9 9 0 2 13 13 1 15 0 2 16 13 4 2
15 0 13 3 9 1 9 13 1 12 9 2 0 7 0 2
2 0 2
21 16 10 9 2 16 3 2 0 13 2 9 3 2 16 13 0 2 13 3 9 2
22 3 9 7 2 16 3 2 3 13 13 9 13 2 1 10 9 13 16 13 9 9 2
6 13 7 15 15 0 2
15 9 3 2 16 13 3 2 3 13 13 9 1 15 13 2
18 3 13 3 13 9 9 1 12 0 9 15 1 15 13 9 10 9 2
2 3 2
26 15 13 1 9 9 2 3 13 9 1 15 2 7 13 1 9 2 16 1 15 13 9 13 1 13 2
20 7 9 1 9 15 3 13 13 16 1 9 9 2 1 10 9 1 9 13 2
7 9 3 13 15 10 13 2
16 9 3 3 13 9 1 15 2 7 1 9 13 1 9 9 2
10 3 3 13 13 12 0 9 10 9 2
2 3 2
6 0 9 13 0 9 2
14 15 3 15 1 12 9 13 2 3 13 13 9 0 2
8 9 7 7 9 15 9 13 2
9 15 3 9 9 13 7 9 13 2
17 3 13 3 2 1 9 9 7 9 1 9 13 2 13 9 0 2
2 0 2
11 15 3 3 13 2 7 0 7 0 13 2
14 15 7 13 2 16 13 2 0 13 2 16 13 4 2
10 13 3 0 13 15 16 13 3 9 2
6 15 7 13 9 13 2
17 9 3 2 16 3 2 13 9 13 2 7 15 9 13 15 9 2
17 9 7 3 13 9 1 15 13 2 16 10 9 13 16 13 9 2
21 7 3 13 1 15 9 9 13 13 9 2 1 9 13 15 0 2 16 1 9 2
22 13 3 16 9 3 13 9 1 15 13 2 7 13 1 9 1 9 9 1 15 13 2
28 3 13 3 12 12 7 1 15 9 9 2 7 0 10 9 13 12 0 9 2 1 15 9 13 9 1 9 2
7 15 13 15 9 12 13 2
21 15 9 2 7 3 13 15 9 2 13 9 7 13 9 2 13 9 7 13 9 2
6 15 9 13 10 15 2
4 7 8 12 2
16 9 7 9 2 9 7 9 2 9 7 9 2 1 9 13 2
4 7 15 12 2
5 1 9 9 13 2
7 3 7 1 9 0 9 2
15 7 3 13 1 10 9 9 12 1 12 2 12 1 12 2
51 13 7 9 13 0 2 7 13 2 16 13 15 15 1 15 0 13 2 7 3 15 13 0 2 16 9 2 16 1 10 9 15 9 9 13 2 3 9 13 0 2 7 0 9 9 2 16 13 15 0 2
13 7 1 0 9 13 9 9 1 9 15 9 13 2
5 3 13 9 12 2
10 16 13 9 1 9 15 9 3 13 2
7 7 15 13 15 9 13 2
13 3 9 2 15 15 10 9 13 2 13 1 9 2
17 7 13 9 13 1 9 1 15 0 13 15 0 13 1 9 13 2
10 1 15 7 13 9 13 0 9 0 2
7 15 9 0 13 1 9 2
22 13 3 12 0 9 13 2 9 7 9 2 15 9 13 13 9 9 2 9 0 9 2
24 1 15 13 2 16 9 13 2 1 12 8 2 15 12 2 9 7 9 2 0 9 0 13 2
24 13 7 7 9 12 0 2 9 7 9 2 7 3 1 9 9 13 2 7 1 9 0 9 2
21 13 3 15 12 13 9 1 15 10 15 13 2 16 13 1 9 2 1 12 0 2
24 15 7 0 9 9 2 15 3 1 0 9 4 0 13 2 15 13 9 9 9 0 13 13 2
43 15 0 13 9 2 1 15 0 4 13 2 15 1 9 0 9 13 2 13 12 15 13 9 2 15 13 4 9 2 7 3 9 2 7 0 9 2 15 15 9 0 13 2
11 16 9 0 9 9 3 13 0 9 9 2
39 1 15 3 13 13 16 9 9 3 13 1 9 0 9 2 16 15 13 13 16 9 2 1 13 12 7 0 2 13 3 12 9 2 15 13 9 0 13 2
35 15 2 16 9 0 9 13 3 13 2 1 3 13 9 0 7 13 15 1 9 13 2 13 15 9 2 16 1 15 3 9 15 13 13 2
22 7 3 3 9 1 9 9 13 2 16 13 9 2 9 9 13 2 1 15 0 13 2
17 15 3 9 15 9 9 3 12 9 13 2 7 0 9 13 9 2
11 15 7 9 9 1 9 10 9 13 13 2
20 15 7 1 9 13 13 15 1 9 0 9 13 7 3 1 15 12 9 13 2
10 9 3 9 7 9 0 13 1 9 2
2 0 2
21 15 15 13 0 1 9 13 2 13 16 1 0 9 1 15 15 13 0 1 9 2
7 13 3 9 0 13 9 2
29 0 7 1 10 9 13 13 9 0 2 1 15 9 0 13 2 16 7 1 9 0 9 9 13 0 16 9 12 2
19 13 3 9 0 16 1 9 0 13 1 9 2 15 1 13 13 0 9 2
23 3 3 9 9 2 1 15 9 13 0 2 13 1 9 0 2 7 3 1 9 9 0 2
2 3 2
16 0 13 15 15 13 0 1 9 13 16 1 9 1 9 9 2
15 0 7 1 9 13 13 9 7 9 15 2 16 13 4 2
19 9 3 13 13 16 15 9 1 15 13 16 0 9 13 1 9 9 0 2
2 3 2
34 1 10 9 13 13 2 16 13 1 9 2 13 16 9 9 0 13 1 9 9 0 2 16 9 0 7 0 7 9 13 1 9 0 2
22 9 7 9 1 0 9 13 1 9 13 1 9 2 1 13 1 9 2 16 13 4 2
7 9 7 10 1 9 13 2
30 16 3 1 9 9 13 15 9 0 2 13 16 9 15 7 9 13 1 9 9 0 2 15 13 0 9 1 9 13 2
15 15 7 13 9 7 9 9 0 2 15 13 3 0 9 2
27 3 3 13 9 1 9 7 9 1 9 0 9 2 7 3 9 0 9 13 1 9 7 9 1 9 13 2
2 3 2
32 16 9 9 0 7 9 15 13 0 9 9 0 2 3 0 9 7 0 1 0 2 13 9 9 7 9 13 1 9 9 0 2
38 1 9 3 15 1 9 13 2 9 15 1 9 13 13 2 13 1 9 0 15 13 1 9 2 16 9 15 13 1 9 2 1 9 15 13 1 9 2
19 9 7 9 7 9 3 13 13 1 9 13 16 13 3 9 13 7 13 2
23 13 3 1 9 0 9 0 9 13 7 13 2 7 15 9 15 13 2 16 1 13 4 2
43 16 3 1 9 15 13 1 9 13 9 1 9 2 1 15 15 1 9 13 2 13 1 0 9 0 13 0 7 0 2 3 13 0 9 2 1 15 15 1 13 9 13 2
2 3 2
21 9 13 1 9 13 1 9 15 13 2 3 1 15 2 16 1 9 7 1 9 2
26 9 7 13 13 1 9 2 16 13 4 2 7 13 15 9 13 0 2 1 3 13 1 10 9 13 2
15 13 3 16 13 9 10 1 15 16 15 9 13 7 13 2
17 7 1 15 9 13 12 9 2 13 7 0 9 15 1 15 13 2
8 13 3 3 0 13 1 0 2
2 0 2
38 16 1 13 4 2 9 0 3 13 1 12 9 2 7 15 15 9 13 2 16 3 15 9 13 3 13 2 3 13 3 0 2 1 0 15 13 13 2
19 16 7 1 12 3 13 16 12 2 3 13 16 16 9 1 12 9 13 2
28 3 13 3 13 16 2 16 9 13 12 7 3 0 2 1 15 9 13 3 13 16 13 15 1 15 9 13 2
2 3 2
9 13 4 1 16 0 9 13 13 2
27 0 7 13 9 15 3 13 13 1 9 16 1 9 2 16 10 15 3 13 13 1 9 7 9 9 13 2
16 3 3 9 13 13 2 1 10 9 13 1 0 7 1 9 2
18 15 7 13 10 0 9 2 7 10 9 0 2 7 3 15 9 0 2
13 13 3 13 10 3 0 1 9 13 15 9 9 2
7 15 13 15 13 8 12 2
8 1 9 13 9 9 7 9 2
3 9 12 2
13 15 3 13 4 9 2 15 0 3 9 13 13 2
12 7 3 3 13 9 9 13 13 1 9 0 2
28 13 7 1 13 9 9 2 15 13 16 9 2 13 15 2 13 12 9 0 2 1 15 3 13 9 7 9 2
39 15 2 16 13 9 2 13 9 0 2 16 0 13 15 1 16 13 1 9 2 13 9 9 2 16 0 13 15 1 16 13 1 9 2 13 9 9 0 2
17 13 3 9 15 0 0 2 15 13 9 3 13 9 2 7 9 2
9 15 9 13 0 9 9 13 9 2
16 16 9 9 3 13 1 15 1 0 9 13 1 9 0 9 2
22 13 7 15 0 0 15 13 9 10 0 13 9 2 7 1 15 9 0 9 4 13 2
6 15 9 9 0 13 2
18 3 3 0 9 2 1 15 15 9 13 2 1 15 9 13 13 13 2
13 10 3 15 13 1 9 13 2 13 1 0 13 2
17 0 13 3 16 1 15 9 0 1 9 13 9 15 0 9 13 2
2 0 2
20 0 9 7 1 15 9 13 1 9 9 2 7 3 13 1 15 9 16 0 2
12 3 3 9 13 1 9 13 2 7 9 0 2
11 15 15 9 13 2 1 9 10 9 0 2
20 9 7 0 3 13 13 1 15 1 10 9 13 2 1 3 13 16 9 3 2
10 10 3 9 1 9 13 1 15 9 2
17 0 13 3 16 1 9 0 1 9 13 15 9 10 0 9 13 2
2 3 2
10 10 15 13 2 1 15 13 16 13 2
7 13 3 13 9 1 9 2
11 3 3 15 13 13 13 16 15 13 9 2
13 9 7 3 13 9 3 7 9 3 2 7 9 2
8 9 3 3 13 16 1 9 2
11 9 0 13 15 15 13 2 13 3 9 2
7 3 13 16 9 0 13 2
11 15 3 0 13 13 2 3 9 1 9 2
14 3 13 3 15 9 13 9 0 2 7 15 13 9 2
2 3 2
15 0 9 9 1 9 3 13 13 1 15 13 1 9 3 2
30 10 3 9 1 9 13 1 9 13 1 9 13 2 16 9 3 13 13 1 10 9 2 7 3 13 15 9 1 9 2
14 7 10 9 1 9 0 0 13 16 13 9 1 9 2
39 1 3 9 0 3 13 1 15 0 2 7 15 9 13 13 9 2 3 13 13 1 9 16 7 1 9 15 9 2 7 1 9 9 1 15 7 15 9 2
25 0 13 3 16 0 9 9 1 9 13 1 15 13 9 3 2 7 1 15 15 13 9 15 9 2
2 3 2
20 9 1 9 13 0 0 9 1 9 2 1 13 9 3 0 2 16 13 9 2
10 0 7 1 9 0 9 13 1 0 2
10 9 3 1 9 13 1 9 1 9 2
9 0 7 9 1 9 13 9 0 2
10 10 3 9 1 9 13 13 9 0 2
24 15 3 15 3 13 13 13 9 0 2 3 13 13 1 15 9 15 3 13 13 16 1 9 2
18 15 13 13 9 15 3 13 13 16 13 9 1 9 2 16 13 4 2
25 1 9 7 0 3 13 13 0 9 0 16 13 13 9 13 2 16 9 15 3 13 16 1 9 2
27 0 3 9 15 9 2 1 15 9 3 13 9 0 1 9 0 9 1 9 2 13 16 13 1 0 13 2
2 3 2
25 16 15 13 9 0 9 7 15 2 16 15 9 7 12 9 2 3 9 9 13 15 15 7 9 2
40 9 7 15 0 7 0 13 13 9 1 9 1 9 15 13 1 9 2 3 7 1 9 1 9 13 2 1 13 13 13 0 13 2 16 13 9 1 12 0 2
20 7 3 0 9 9 1 9 13 13 1 9 1 15 9 13 2 3 13 9 2
19 7 7 13 16 15 13 13 9 0 2 7 1 13 2 15 13 1 9 2
2 3 2
15 16 9 13 0 1 9 2 3 13 0 9 16 0 9 2
11 9 7 13 1 9 2 7 3 1 9 2
10 0 3 9 9 0 13 0 9 13 2
2 0 2
32 1 10 9 13 15 0 2 1 15 13 9 9 15 1 9 13 13 2 16 9 1 9 1 9 2 15 13 9 9 1 9 2
29 7 10 13 9 15 13 9 0 2 16 13 9 2 1 15 13 1 9 2 7 16 9 13 2 0 9 13 13 2
16 0 13 3 13 16 9 9 1 15 13 16 1 9 10 9 2
34 7 3 13 16 2 1 13 15 9 2 8 12 2 9 2 16 13 9 1 9 9 7 9 13 2 13 3 10 1 0 9 13 13 2
29 7 9 13 2 8 12 2 16 1 0 13 4 0 2 7 15 1 9 13 7 15 1 9 2 7 0 7 0 2
11 16 9 9 3 13 1 9 7 9 9 2
24 3 13 13 16 9 9 3 13 1 0 9 0 9 0 9 2 16 13 9 2 1 9 8 2
81 13 3 13 0 0 9 7 9 2 15 13 13 0 9 9 7 9 13 1 9 1 0 9 2 1 0 9 13 3 1 9 0 7 1 9 0 2 15 15 9 13 13 2 3 16 15 9 13 0 2 15 0 2 15 9 1 9 2 15 1 0 13 2 13 4 13 10 9 1 9 13 1 9 9 2 1 9 9 2 13 2
20 13 3 16 9 1 0 10 9 0 10 9 0 13 2 7 10 0 7 0 2
24 15 1 0 9 9 4 13 2 15 13 9 0 7 0 2 15 1 15 13 7 3 7 0 2
37 7 1 15 0 9 1 9 0 1 0 9 4 13 2 16 15 13 9 1 0 9 2 15 9 0 3 1 0 9 2 15 3 9 1 9 0 2
32 7 1 9 0 9 13 9 0 9 9 13 2 16 0 9 0 0 9 13 2 16 9 0 9 0 9 9 15 9 15 13 2
8 15 7 9 0 13 0 13 2
15 3 3 15 13 0 1 9 2 3 13 0 1 9 9 2
16 0 7 1 9 13 13 9 0 2 15 13 1 9 13 9 2
10 1 10 3 9 15 13 9 0 9 2
15 3 9 9 1 0 9 0 9 13 2 3 1 9 9 2
2 3 2
23 16 10 9 0 1 9 4 0 13 2 13 13 16 12 15 1 10 9 1 15 3 13 2
17 15 7 13 1 9 0 9 15 12 1 15 3 13 2 13 0 2
14 3 2 1 13 9 2 15 9 7 9 9 13 0 2
9 15 13 0 2 16 1 13 4 2
2 0 2
12 15 13 15 0 2 3 13 1 15 1 9 2
18 9 3 9 2 7 0 9 2 13 9 13 2 1 15 15 0 13 2
24 16 3 1 9 0 9 13 4 0 9 0 9 2 15 9 0 13 10 9 0 2 7 0 2
5 15 7 13 0 2
38 1 3 9 0 13 15 0 2 13 16 10 9 0 13 13 12 9 2 3 9 2 9 2 7 9 0 2 7 9 0 9 2 15 9 13 13 2 2
9 7 15 13 0 9 9 0 13 2
52 3 3 13 15 9 15 0 13 9 0 2 15 9 7 9 13 2 7 9 0 7 9 9 2 16 9 13 9 7 0 9 13 9 7 9 7 15 3 9 2 1 15 16 13 9 9 13 2 15 13 0 2
18 13 3 16 9 9 0 3 13 9 9 2 15 13 1 9 0 9 2
2 3 2
42 16 15 15 13 0 3 13 1 9 0 9 2 9 7 0 15 9 13 13 15 1 13 9 7 9 1 9 0 9 2 13 16 9 15 9 1 15 9 3 13 0 2
6 3 7 9 13 0 2
21 9 7 2 7 9 2 1 9 2 7 9 2 13 13 1 9 0 7 9 15 2
14 3 10 3 2 15 13 0 1 0 9 2 13 0 2
2 3 2
34 16 15 9 0 3 13 16 13 15 9 15 9 13 2 7 3 16 4 3 13 2 15 9 13 3 13 15 1 15 2 7 1 9 2
21 1 15 7 15 1 9 13 3 13 15 9 2 16 3 13 1 15 12 1 15 2
11 3 3 13 15 9 9 0 7 9 13 2
19 13 3 16 9 3 13 15 9 2 7 9 2 7 9 2 7 15 3 2
2 0 2
14 15 15 1 9 13 2 13 1 0 7 1 0 13 2
27 9 3 7 9 13 13 7 13 2 7 0 1 9 2 15 13 0 9 15 9 3 13 1 15 9 0 2
41 16 3 9 0 15 9 13 4 1 13 9 7 9 2 13 16 13 3 13 15 9 2 7 3 0 16 9 0 13 15 9 0 2 7 3 16 13 3 9 0 2
12 15 13 1 0 9 2 15 9 15 9 13 2
38 15 7 7 1 9 13 13 0 2 1 15 13 9 7 9 13 13 9 7 13 0 2 7 1 9 0 2 15 9 1 9 15 9 13 13 15 13 2
2 3 2
25 1 9 1 9 13 3 13 2 16 13 1 9 9 0 1 15 9 13 2 13 15 15 9 13 2
10 15 3 13 12 15 15 3 13 15 2
22 7 3 15 1 9 9 3 13 2 0 9 7 13 0 16 9 9 1 9 9 13 2
2 3 2
32 10 9 13 7 1 9 9 2 15 1 0 9 13 2 3 1 9 0 13 2 1 9 2 13 3 13 2 7 1 9 0 2
17 15 1 9 9 13 3 13 2 1 15 9 13 1 9 7 9 2
13 7 3 13 16 15 9 13 13 0 7 15 0 2
18 3 2 1 9 2 9 9 13 16 9 2 15 12 15 13 7 13 2
20 3 3 2 16 13 1 9 0 9 0 13 2 13 16 13 1 15 9 9 2
2 3 2
35 16 9 0 1 9 13 13 2 3 13 0 1 0 9 0 9 9 1 9 0 13 2 16 7 1 9 9 13 0 9 1 9 0 13 2
23 16 7 9 0 1 9 13 3 13 2 3 1 9 3 1 9 0 4 3 9 0 13 2
14 0 13 7 9 0 9 1 0 16 0 9 1 3 2
32 16 3 1 9 9 3 0 9 1 10 9 13 1 15 9 13 2 3 13 9 0 13 1 15 16 1 0 9 9 0 13 2
2 3 2
20 16 9 9 0 13 9 9 0 2 0 9 7 9 0 9 13 9 9 0 2
17 4 3 9 0 13 3 16 0 9 0 9 3 13 2 7 0 2
18 4 3 13 9 0 2 15 13 10 9 0 2 7 1 12 3 9 2
9 13 7 1 15 0 9 1 9 2
12 13 3 0 2 0 12 15 9 13 1 9 2
7 15 3 13 13 0 9 2
2 3 2
42 16 9 0 9 13 0 9 0 9 0 9 2 13 13 16 9 3 13 3 12 9 1 9 2 13 16 12 3 0 9 3 13 4 1 0 9 16 15 9 13 13 2
12 15 7 13 1 9 2 16 12 3 3 13 2
18 13 3 1 9 16 13 12 9 1 9 2 7 3 1 9 0 9 2
2 3 2
39 1 9 0 3 13 13 16 1 9 2 13 7 1 10 9 2 1 15 0 13 2 1 15 16 0 9 13 2 13 13 16 0 9 13 15 13 1 9 2
13 15 13 0 9 9 13 15 0 1 0 9 13 2
9 15 3 9 9 0 9 0 13 2
20 16 1 0 9 0 9 15 9 13 13 9 2 13 9 16 13 0 2 8 2
7 7 3 1 10 3 13 2
11 13 9 10 15 13 2 7 13 3 0 2
35 1 15 0 13 13 16 9 0 7 0 3 4 13 16 0 13 15 13 2 15 13 0 0 9 2 7 3 1 15 9 0 9 7 9 2
35 13 7 9 3 13 16 2 1 15 3 1 9 2 7 0 13 2 3 13 1 9 16 0 13 2 15 9 9 13 2 1 9 13 13 2
21 9 7 2 16 1 13 4 2 1 15 9 2 7 1 0 9 9 1 9 13 2
8 3 9 9 9 9 3 13 2
25 3 2 1 9 15 13 0 16 9 9 0 2 3 13 0 9 13 9 15 16 15 9 13 9 2
16 3 3 9 9 13 15 9 15 13 13 2 16 9 13 0 2
34 9 3 10 2 9 2 3 13 15 0 1 10 9 0 2 16 13 10 9 0 2 16 0 9 9 1 0 13 2 7 3 13 0 2
9 15 13 0 9 9 9 1 9 2
13 13 7 1 13 13 15 13 0 0 9 9 9 2
25 1 3 10 9 13 10 9 1 9 13 1 16 9 13 13 2 3 15 13 9 3 9 9 13 2
27 13 3 16 3 15 13 0 2 3 13 3 0 2 7 3 13 15 0 9 2 9 9 9 13 1 9 2
6 9 7 13 9 9 2
17 10 3 9 1 9 13 1 9 13 13 9 2 3 9 13 13 2
44 7 9 9 9 3 13 13 9 13 1 12 0 9 9 2 16 2 1 9 13 9 2 15 13 1 9 0 7 13 2 1 9 13 13 7 0 2 16 9 13 1 9 9 2
15 15 1 13 13 3 13 2 3 3 9 13 13 9 0 2
23 13 3 13 9 7 9 1 9 13 2 1 15 16 13 1 15 9 9 9 1 9 10 2
2 0 2
23 16 15 13 1 9 13 1 9 9 0 2 3 15 13 1 9 13 13 1 9 0 9 2
23 3 7 9 0 9 9 13 1 9 16 1 9 13 12 3 15 1 15 9 13 1 9 2
30 3 2 16 15 9 15 9 13 1 0 9 2 13 12 15 3 2 9 15 3 3 13 13 1 9 16 1 13 0 2
15 1 15 7 16 9 0 13 1 9 2 9 13 9 9 2
16 3 3 13 9 9 9 1 0 16 13 12 3 9 10 9 2
20 1 15 3 13 9 1 9 13 2 16 9 9 9 13 1 0 16 1 12 2
2 3 2
15 3 15 1 0 13 9 0 2 3 9 1 15 9 13 2
12 1 9 7 13 9 2 7 9 9 1 15 2
42 9 3 13 9 13 1 9 9 16 3 0 0 13 7 3 1 9 15 13 13 2 16 1 0 1 15 0 13 2 16 0 13 9 15 13 7 13 16 15 13 3 2
29 3 7 13 9 1 9 15 9 13 16 13 1 9 13 9 7 9 2 16 9 13 15 1 0 2 7 0 15 2
20 13 3 2 1 15 16 1 9 13 9 9 9 2 16 0 9 1 9 13 2
2 3 2
8 0 9 12 9 13 13 0 2
7 13 3 15 7 3 0 2
7 10 7 9 9 13 13 2
8 13 3 13 1 0 9 9 2
17 9 13 3 0 9 16 13 0 2 16 16 13 12 3 9 9 2
9 0 7 9 13 13 15 0 13 2
10 3 13 15 13 16 0 13 9 9 2
2 3 2
13 9 9 13 9 9 2 16 0 15 15 13 0 2
15 3 3 13 1 9 0 9 9 1 9 9 1 12 9 2
29 13 3 1 9 0 13 3 0 16 0 13 9 2 7 16 13 3 0 9 9 2 7 1 13 0 9 1 9 2
2 3 2
14 10 15 13 1 9 2 13 9 10 9 1 9 13 2
9 3 3 9 1 9 15 13 0 2
20 9 7 13 9 16 13 1 9 2 7 3 1 9 9 2 16 1 13 4 2
11 9 3 9 0 13 1 9 1 15 13 2
11 9 7 0 13 3 0 13 1 12 3 2
28 1 3 9 0 0 13 2 16 1 0 13 4 2 9 15 13 16 0 0 9 9 13 16 16 12 3 13 2
2 0 2
12 9 1 0 0 9 13 3 13 13 0 9 2
13 7 9 9 0 13 0 15 15 13 1 15 13 2
12 13 3 0 9 0 2 16 9 15 9 9 2
9 3 13 3 9 9 9 9 13 2
15 15 7 9 13 3 13 2 16 9 7 9 9 3 13 2
41 13 3 9 7 9 1 9 13 3 1 9 2 3 1 9 9 2 3 1 9 15 9 2 7 9 2 7 1 0 9 9 9 9 13 13 15 0 13 15 13 2
7 15 13 15 13 8 12 2
19 13 9 10 15 13 2 7 13 3 0 2 1 1 0 13 16 13 0 2
28 16 0 3 13 1 10 9 0 2 3 7 10 3 0 2 1 9 0 2 15 13 0 7 0 9 1 9 2
10 16 13 1 9 0 15 9 0 13 2
28 15 3 13 9 9 1 9 2 13 3 1 9 13 13 2 3 1 9 9 13 2 15 13 0 1 15 13 2
31 7 13 0 2 16 1 0 9 9 9 13 1 10 9 0 13 2 13 13 16 15 9 0 13 2 1 0 9 9 13 2
12 3 3 9 0 9 13 16 1 10 13 9 2
25 3 7 9 1 10 9 2 7 9 0 1 10 9 2 13 0 9 2 16 1 15 1 9 13 2
17 1 15 3 16 0 9 0 9 13 2 13 9 1 10 13 9 2
55 13 7 1 10 9 0 7 10 9 16 10 9 9 13 1 10 9 7 10 9 2 1 15 15 9 13 2 16 7 10 9 3 0 9 13 16 0 13 9 13 2 16 9 16 0 13 9 2 7 9 16 0 13 13 2
25 1 3 9 9 9 9 9 13 2 16 1 13 4 2 0 13 1 9 9 16 15 9 13 13 2
2 0 2
8 9 0 1 9 13 1 0 2
17 16 7 9 7 9 9 13 1 0 9 2 3 9 1 9 0 2
26 13 3 2 1 13 0 9 2 13 15 9 15 1 9 13 3 0 1 9 9 2 7 3 1 9 2
22 15 3 3 13 13 16 1 9 9 7 9 2 16 7 15 9 15 1 15 9 13 2
13 13 3 2 1 9 0 0 2 13 15 9 0 2
2 3 2
33 1 15 16 9 0 9 9 1 9 13 2 13 2 16 1 13 4 2 3 0 16 9 0 13 2 7 3 16 1 15 9 13 2
21 13 7 9 15 15 1 13 16 3 0 13 15 9 9 2 7 3 15 9 13 2
20 13 3 2 1 0 9 9 2 16 13 15 9 15 13 15 9 15 9 13 2
12 13 4 7 1 16 9 13 1 9 7 9 2
9 13 3 15 9 13 13 7 13 2
2 0 2
14 9 9 1 9 13 13 1 9 9 15 13 1 9 2
11 9 3 13 15 0 1 9 1 15 13 2
30 9 7 9 13 3 1 9 3 1 15 9 13 15 13 1 9 2 16 9 9 13 15 13 13 9 1 9 9 13 2
26 3 0 1 15 9 13 2 16 9 9 15 13 0 1 9 9 2 13 0 1 9 15 13 1 9 2
9 13 7 9 13 0 9 16 0 2
21 9 7 9 9 13 1 9 1 9 2 16 3 9 15 9 1 9 1 9 13 2
20 13 3 0 0 9 3 0 0 9 9 1 9 2 7 0 2 3 0 13 2
14 9 7 1 15 9 13 9 2 13 9 0 1 15 2
11 13 3 9 1 9 2 16 1 13 4 2
19 13 3 1 0 9 0 13 15 9 1 15 1 9 0 9 0 9 13 2
10 7 15 13 13 9 1 10 9 0 2
2 3 2
27 1 9 9 15 15 13 9 16 10 9 2 15 9 15 13 13 1 9 9 1 15 2 16 1 13 13 2
42 9 7 12 13 1 15 0 2 12 9 2 3 1 9 9 2 16 9 9 0 13 1 9 13 1 9 2 15 9 2 1 9 2 16 9 9 13 1 9 7 9 2
29 1 15 3 16 9 9 9 13 1 9 9 0 2 13 16 0 9 9 1 9 13 3 0 1 13 2 7 13 2
8 13 7 0 9 0 9 13 2
6 13 3 13 9 0 2
2 3 2
21 1 10 13 13 9 0 1 0 13 9 0 1 10 0 7 0 2 16 3 13 2
11 13 4 7 16 9 1 15 10 9 13 2
12 7 15 13 1 0 9 2 16 1 15 9 2
29 3 3 13 0 9 13 7 13 9 2 3 1 9 9 2 1 9 10 9 0 9 2 7 3 9 9 2 13 2
32 16 3 7 1 15 9 13 9 9 9 13 2 13 4 9 0 2 15 9 0 13 2 3 9 9 2 7 0 1 9 0 2
13 3 15 13 13 1 13 2 7 15 0 9 13 2
6 16 9 0 13 13 2
9 15 7 9 0 0 13 13 13 2
17 13 3 10 9 9 2 1 9 13 15 10 13 2 16 9 13 2
22 3 7 9 1 15 3 15 9 13 2 13 0 9 2 16 13 16 9 13 13 3 2
19 1 15 7 15 9 0 13 2 13 9 0 2 15 13 1 0 7 0 2
16 1 15 0 15 13 2 13 9 0 7 0 2 15 13 9 2
7 9 3 0 13 13 9 2
2 3 2
16 15 13 1 15 2 13 1 15 15 13 1 15 16 1 0 2
19 3 7 2 1 9 2 1 12 8 2 13 1 15 13 1 0 13 15 2
22 1 9 3 9 2 15 13 13 1 15 2 13 1 0 9 2 15 13 13 1 15 2
26 13 7 1 9 13 15 15 3 13 15 1 13 2 7 13 9 9 2 16 0 2 9 7 9 0 2
10 3 3 13 1 15 13 7 3 13 2
14 13 3 16 13 9 1 15 0 15 15 13 1 13 2
14 0 7 1 9 13 13 9 0 2 16 1 13 4 2
8 15 3 9 15 13 1 13 2
24 15 7 13 0 9 2 1 15 9 15 13 9 10 9 2 16 1 15 13 13 7 3 13 2
7 9 3 0 13 13 9 2
2 0 2
19 9 15 9 13 9 1 15 15 13 9 2 1 10 9 13 16 13 9 2
12 13 3 16 1 9 9 13 9 9 13 9 2
19 9 3 15 3 13 1 15 13 1 9 2 13 9 15 9 3 13 9 2
21 16 15 0 13 9 15 13 1 15 15 1 15 13 2 9 3 13 13 9 13 2
26 9 7 0 2 1 15 13 9 7 9 0 2 3 13 1 15 15 13 9 2 7 1 0 9 0 2
19 1 1 9 0 15 13 13 1 10 9 2 15 7 13 13 15 9 13 2
10 7 3 15 13 0 2 3 13 15 2
15 3 3 0 13 15 3 2 7 13 2 15 13 15 9 2
37 1 9 3 0 9 0 7 13 13 3 4 13 1 15 9 0 2 7 4 13 1 15 1 0 0 2 15 13 1 9 2 7 13 1 0 0 2
38 3 2 16 3 13 13 15 2 16 15 12 9 13 13 7 15 13 13 2 3 15 13 3 13 15 1 15 2 7 9 1 0 0 7 9 1 9 2
17 16 3 9 13 9 2 13 15 13 2 15 13 1 0 7 9 2
26 16 0 15 13 1 9 13 1 15 1 9 13 1 9 7 9 0 9 2 3 15 13 9 16 13 2
7 3 3 13 9 10 9 2
39 9 7 13 2 1 15 9 0 13 2 13 1 15 9 2 16 1 15 13 7 3 13 2 16 13 1 9 9 2 15 9 13 7 13 7 1 15 13 2
14 9 3 0 15 13 1 13 2 16 13 10 9 9 2
4 13 3 9 2
2 3 2
10 0 13 13 13 0 2 7 9 0 2
15 7 1 13 9 9 0 15 13 1 0 16 9 1 0 2
15 3 13 1 9 7 9 7 9 2 13 9 0 7 0 2
12 9 7 0 3 13 1 15 2 7 13 10 2
20 3 7 1 9 0 9 13 2 1 12 1 9 2 16 13 15 13 10 13 2
10 9 3 0 9 13 1 10 15 13 2
12 15 7 13 0 9 2 16 1 10 15 13 2
13 3 1 12 9 9 13 16 13 7 0 7 0 2
6 9 3 0 13 9 2
9 16 9 0 13 0 9 1 13 2
13 1 15 7 13 16 13 9 13 0 9 1 13 2
18 16 3 9 13 2 0 13 2 15 16 1 9 0 9 13 1 13 2
17 9 7 0 13 15 13 2 16 13 9 10 9 2 16 13 4 2
9 13 3 13 9 0 9 1 13 2
2 3 2
7 0 13 15 15 9 13 2
14 15 3 3 13 15 9 13 2 3 13 0 1 13 2
18 15 7 3 13 7 13 16 1 15 13 2 3 13 15 15 9 13 2
10 0 3 13 15 15 9 1 13 13 2
6 7 15 0 9 13 2
9 3 13 15 13 1 13 7 13 2
16 13 7 13 9 1 9 7 9 7 9 13 2 15 13 13 2
12 15 3 15 0 0 13 15 1 13 15 13 2
14 15 7 9 13 15 1 13 13 16 1 9 10 13 2
14 13 3 2 16 15 1 13 13 2 16 10 9 13 2
6 15 3 0 9 13 2
16 13 3 9 0 3 0 3 9 7 9 2 3 7 0 9 2
16 0 7 2 15 0 1 15 13 2 7 3 0 9 7 9 2
17 0 0 3 0 9 2 7 3 0 9 2 15 13 0 9 13 2
2 3 2
14 9 13 13 9 13 1 16 13 1 9 0 7 13 2
20 9 3 0 1 13 15 13 1 9 15 13 15 13 0 7 13 1 9 13 2
20 16 3 13 1 13 15 13 2 13 16 1 15 9 9 13 15 13 1 13 2
22 15 3 13 3 13 16 15 9 9 7 13 2 1 15 1 15 13 9 7 13 13 2
15 15 3 0 15 1 13 13 15 0 9 7 13 9 13 2
6 15 7 13 0 0 2
15 0 3 0 15 3 0 1 13 2 7 3 1 13 13 2
14 0 16 15 13 0 1 13 2 15 13 0 9 13 2
2 0 2
22 1 9 0 3 13 9 7 9 16 13 0 9 2 15 16 9 7 9 1 0 13 2
7 9 7 13 0 0 0 2
22 1 15 3 16 1 9 9 13 9 7 15 9 2 13 16 0 9 9 13 1 0 2
8 7 0 13 1 9 0 0 2
11 13 3 9 9 0 13 1 0 7 0 2
12 9 3 9 1 0 3 13 13 1 12 3 2
7 13 3 10 0 0 9 2
2 3 2
36 9 9 13 15 7 1 15 16 15 13 9 2 16 15 9 13 2 16 9 7 9 2 7 16 13 9 1 9 13 1 12 2 16 0 9 2
16 0 3 9 13 9 9 15 0 2 7 1 15 9 13 15 2
5 0 7 1 15 2
19 15 3 13 9 1 13 3 13 1 9 1 12 2 0 13 0 9 13 2
6 3 7 13 10 0 2
15 9 3 13 3 0 15 7 15 9 2 7 15 9 0 2
33 3 2 1 9 1 9 13 13 9 2 1 10 7 13 7 13 13 13 13 2 9 9 0 3 4 13 1 9 16 1 9 0 2
21 15 3 13 15 1 9 9 2 13 9 13 1 15 2 15 9 0 1 0 13 2
11 10 3 0 0 9 13 1 9 9 13 2
14 15 13 0 9 13 2 15 13 13 0 1 9 9 2
7 16 9 0 3 13 9 2
11 1 13 7 13 16 15 9 0 13 9 2
11 15 3 9 13 15 13 16 1 9 9 2
23 3 7 2 16 15 15 15 15 13 2 7 9 9 13 2 0 3 0 2 0 7 0 2
28 9 7 3 13 9 15 13 1 15 9 9 2 1 15 15 13 7 13 15 7 9 2 0 1 9 7 0 2
7 15 3 9 13 13 9 2
2 0 2
15 15 9 13 15 9 9 0 13 16 1 9 10 9 13 2
16 9 7 3 13 2 7 3 13 1 15 16 13 9 10 9 2
5 13 3 1 13 2
10 13 7 1 16 13 1 15 9 13 2
7 15 3 9 0 13 9 2
2 3 2
11 9 9 9 15 9 13 9 9 1 9 2
35 9 3 15 9 1 9 15 9 3 13 16 1 15 16 13 1 0 9 1 15 9 13 2 7 15 16 9 9 2 1 15 9 13 0 2
13 15 7 13 1 9 2 13 1 15 1 9 9 2
10 3 9 3 13 1 9 16 16 13 2
17 16 3 9 13 9 2 9 9 0 3 13 1 15 16 16 13 2
12 13 7 9 9 1 9 15 15 1 15 13 2
10 3 3 9 13 0 2 7 0 0 2
5 15 13 13 0 2
6 15 3 9 13 9 2
2 3 2
16 15 13 16 1 10 9 2 15 16 9 13 9 13 1 15 2
13 16 3 9 13 9 2 9 15 9 9 3 13 2
6 3 3 13 16 9 2
6 15 7 13 13 0 2
8 13 3 0 15 3 13 9 2
6 9 3 3 13 9 2
2 3 2
13 16 9 13 13 9 2 7 13 13 2 7 0 2
13 9 7 13 0 9 13 0 2 16 1 9 13 2
10 13 3 13 9 2 16 9 13 13 2
5 15 7 13 0 2
15 1 15 3 9 13 13 13 9 0 2 16 1 13 4 2
9 9 7 9 13 3 0 1 13 2
15 1 0 3 13 9 9 13 2 7 0 9 9 7 9 2
20 13 3 0 2 15 13 9 0 1 10 9 2 13 3 9 15 13 9 0 2
6 9 3 3 13 9 2
2 0 2
8 0 13 12 9 15 3 13 2
5 1 13 13 13 2
14 12 7 9 15 3 13 7 13 2 16 12 15 13 2
6 3 13 3 9 9 2
2 3 2
7 15 9 9 13 1 9 2
27 13 4 3 1 9 16 15 9 1 15 13 16 1 9 2 3 3 16 12 9 15 13 13 7 15 13 2
7 9 7 1 15 13 13 2
12 13 3 15 3 0 1 9 2 7 1 15 2
5 3 13 3 9 2
2 3 2
18 9 9 1 9 3 13 2 7 9 1 9 2 16 1 9 4 13 2
8 9 7 9 13 1 9 13 2
17 9 3 2 16 13 9 2 3 13 15 13 2 7 3 1 0 2
7 9 3 13 3 13 9 2
27 15 13 16 0 9 9 0 9 13 2 1 15 9 13 9 0 13 2 1 15 8 12 2 9 9 13 2
22 13 7 8 12 13 7 1 15 2 3 0 9 2 9 9 2 15 13 10 9 0 2
16 1 15 7 13 9 0 0 2 15 15 9 16 0 13 13 2
18 3 7 9 13 13 9 2 7 9 7 9 7 9 2 7 15 3 2
22 15 3 9 1 9 0 15 13 4 13 2 13 9 13 9 13 2 16 9 0 13 2
6 16 9 0 13 0 2
10 1 15 7 13 16 9 0 13 0 2
10 15 3 1 9 7 9 9 13 9 2
12 0 3 9 9 3 16 1 0 9 13 13 2
24 15 3 9 9 13 1 9 3 13 16 1 16 1 9 1 9 13 12 0 9 1 0 13 2
8 13 3 9 2 9 0 13 2
10 13 4 7 16 15 9 13 13 9 2
11 13 3 16 3 13 1 9 7 9 13 2
2 0 2
16 16 9 3 13 1 15 9 2 3 9 3 13 1 15 9 2
20 15 3 1 9 13 0 1 9 7 9 13 2 13 13 1 9 7 9 0 2
12 9 7 3 13 13 13 1 9 7 9 0 2
15 9 3 9 13 13 0 9 1 15 16 1 9 0 13 2
12 1 7 16 13 0 9 2 13 12 1 9 2
9 3 7 9 13 13 1 9 0 2
11 3 13 3 9 13 1 9 7 9 13 2
2 3 2
19 9 15 1 9 7 9 9 3 13 3 9 2 7 3 9 2 7 9 2
8 15 3 13 13 15 13 9 2
7 13 7 13 9 1 9 2
7 3 7 9 1 9 13 2
16 16 3 9 13 13 13 1 9 7 9 2 13 13 15 9 2
8 9 7 13 1 15 0 9 2
11 3 7 9 13 3 13 9 2 7 9 2
18 16 3 13 13 9 9 2 3 13 7 9 7 9 2 7 3 9 2
6 15 7 13 13 0 2
11 3 13 3 9 13 13 1 9 7 9 2
2 3 2
13 9 9 0 9 9 13 1 9 16 1 9 0 2
9 13 3 0 7 1 0 15 13 2
12 1 12 3 9 9 0 2 10 9 9 13 2
18 9 7 9 1 9 13 13 13 9 15 2 3 7 9 2 7 13 2
30 16 7 3 13 15 13 15 2 13 0 1 15 2 16 9 9 1 9 16 1 13 2 7 16 9 0 9 1 9 2
24 16 3 9 13 1 9 7 9 13 2 9 9 13 13 9 13 9 15 9 15 13 15 13 2
23 7 3 13 9 9 2 15 13 16 9 9 13 9 2 7 9 9 2 7 3 1 15 2
5 15 13 13 9 2
11 3 13 3 13 9 13 1 9 7 9 2
2 3 2
12 10 15 13 1 15 13 1 15 1 9 13 2
22 16 3 9 13 13 1 9 7 9 2 9 9 13 1 9 0 2 16 13 1 9 2
15 16 3 1 9 3 13 0 9 2 3 3 13 1 9 2
2 3 2
13 9 0 2 1 9 15 13 1 9 2 13 0 2
6 3 7 15 3 13 2
25 1 7 16 13 1 9 2 3 13 0 2 7 12 0 13 9 0 15 2 16 12 1 15 13 2
8 3 3 13 9 0 1 9 2
10 3 9 3 13 13 1 9 7 9 2
2 3 2
13 9 3 13 15 9 1 0 16 1 9 7 9 2
24 9 7 3 13 1 15 16 13 9 2 7 3 13 7 13 13 2 13 7 1 13 1 9 2
14 3 3 13 9 1 9 16 1 9 7 1 9 0 2
12 3 13 16 9 13 0 13 2 16 7 0 2
12 15 13 15 9 13 2 12 8 1 8 8 2
16 1 0 9 9 13 0 10 9 2 15 16 0 7 0 13 2
8 16 9 0 3 13 9 0 2
23 1 15 7 13 16 9 0 13 9 13 2 3 7 13 1 9 16 9 15 1 9 13 2
18 9 3 1 13 1 9 13 3 15 0 13 9 2 7 9 1 15 2
24 16 3 9 0 13 3 9 2 13 16 13 9 0 2 16 7 16 13 1 9 7 9 13 2
2 3 2
19 9 15 1 15 3 13 2 3 13 1 15 13 2 13 7 9 1 15 2
21 16 3 9 0 3 9 13 2 13 16 15 3 13 2 7 9 1 15 7 9 2
10 7 3 13 13 9 1 9 7 9 2
8 15 13 0 2 16 13 4 2
2 0 2
23 16 9 13 9 1 9 7 3 1 15 0 2 13 16 15 15 13 1 9 13 1 9 2
18 3 3 9 15 13 9 9 13 2 3 13 15 15 1 9 3 13 2
21 1 3 9 9 1 9 3 13 9 9 1 9 2 0 13 16 9 13 9 0 2
2 3 2
33 13 16 9 13 9 3 0 7 9 13 2 15 13 1 9 7 16 13 16 9 13 13 1 9 7 9 2 13 7 0 1 9 2
19 3 0 9 2 13 9 15 9 9 2 0 0 9 2 13 9 15 9 2
22 16 3 0 13 9 13 13 1 9 7 9 2 0 13 16 13 9 3 0 7 0 2
11 16 1 9 0 13 13 9 7 15 13 2
35 3 13 7 13 16 2 16 9 0 3 13 0 2 7 1 9 7 9 13 2 7 1 9 13 16 9 0 2 16 1 15 0 9 13 2
19 13 3 1 15 15 9 1 15 16 3 13 15 1 15 9 7 15 13 2
13 16 3 9 13 0 2 15 1 15 9 15 13 2
83 16 3 1 15 15 9 3 13 0 2 16 13 13 1 9 15 2 13 3 13 13 2 3 7 13 12 1 9 15 2 16 1 9 2 16 13 12 9 13 9 7 15 15 13 1 9 2 16 13 16 9 2 1 10 9 0 2 13 0 2 15 3 0 13 1 15 9 0 2 3 3 15 13 13 9 7 13 0 2 16 1 9 2
23 16 3 3 13 9 1 15 9 2 3 13 15 9 15 13 15 13 15 15 13 1 9 2
12 9 7 2 16 13 9 2 3 13 13 0 2
19 13 7 13 1 15 15 13 1 9 2 16 9 9 13 15 1 9 9 2
14 15 3 15 13 9 0 2 3 13 13 16 12 3 2
10 13 4 7 16 9 13 10 9 0 2
10 15 3 15 1 15 13 13 10 9 2
18 13 3 1 10 9 15 13 1 15 2 13 15 15 9 7 9 15 2
2 0 2
21 9 0 2 16 13 13 2 3 13 13 16 12 2 16 13 9 15 0 13 13 2
20 16 3 9 9 1 15 13 13 2 3 13 15 15 13 9 7 15 13 9 2
12 3 3 3 13 9 3 2 7 9 7 9 2
22 13 7 9 0 9 2 13 9 9 0 2 16 15 9 15 13 0 9 13 0 9 2
25 3 3 2 16 15 15 15 13 9 13 0 16 9 2 9 13 1 15 0 3 13 13 16 12 2
36 16 0 3 13 9 2 16 9 2 7 1 15 16 13 15 7 15 9 2 16 9 13 2 3 13 0 16 3 13 13 1 15 13 16 12 2
18 13 3 16 2 1 9 13 9 0 2 15 15 1 15 13 10 9 2
2 3 2
9 0 13 16 13 0 9 3 0 2
29 9 3 15 3 13 0 2 10 9 13 13 2 7 3 2 16 12 15 13 9 2 3 13 15 12 1 15 13 2
13 9 7 0 13 13 0 2 16 3 13 15 13 2
10 0 13 3 13 15 9 0 1 0 2
2 3 2
19 16 13 15 9 1 15 0 2 15 13 15 16 16 13 9 16 13 9 2
19 15 3 13 1 15 3 16 3 2 3 13 15 16 1 9 2 9 9 2
13 3 2 16 13 1 9 13 2 15 9 15 13 2
12 9 7 1 15 13 3 13 9 16 13 9 2
26 15 10 9 13 1 15 13 2 7 3 13 13 1 0 1 9 2 15 13 0 2 16 1 13 4 2
13 15 3 9 15 13 0 2 13 16 13 3 13 2
8 15 3 9 13 13 10 9 2
2 0 2
11 9 15 13 15 1 15 7 3 1 15 2
16 3 13 0 9 3 13 1 9 9 2 16 13 15 1 15 2
11 7 15 9 13 10 9 13 15 1 15 2
5 15 3 13 13 2
10 15 3 9 13 10 9 13 10 9 2
2 3 2
22 1 10 9 13 16 13 9 2 0 9 2 15 13 9 2 13 13 1 9 9 9 2
16 3 7 15 13 9 1 9 3 15 9 13 1 9 9 0 2
17 9 3 13 9 9 0 1 12 7 15 15 1 9 1 9 13 2
15 9 3 13 1 9 15 13 15 9 16 15 13 13 9 2
7 15 3 1 15 9 13 2
16 15 3 3 13 2 13 1 1 13 16 9 0 13 0 9 2
17 15 3 0 13 13 1 9 9 9 2 16 3 13 15 9 9 2
13 15 7 13 13 2 1 15 9 7 10 9 13 2
12 10 3 9 7 9 13 1 9 16 9 13 2
17 0 3 9 13 16 13 15 9 2 16 0 13 16 13 0 9 2
2 0 2
9 15 9 13 0 9 1 0 9 2
11 9 3 9 13 15 9 16 1 13 4 2
24 15 7 13 15 1 0 9 10 2 3 13 15 16 1 9 9 2 16 9 15 9 1 9 2
13 15 3 9 13 10 15 1 0 9 1 9 15 2
12 15 7 13 15 1 9 2 3 13 9 15 2
14 0 13 3 16 9 15 9 1 9 0 13 15 9 2
28 15 13 16 9 12 0 9 9 13 13 15 13 2 16 15 0 0 13 16 10 9 3 13 15 16 10 9 2
10 16 1 9 0 13 13 9 7 9 2
16 1 15 7 0 13 16 1 9 0 13 13 9 9 7 9 2
24 1 15 3 13 15 12 15 12 13 9 15 2 9 12 15 1 15 13 16 9 9 1 9 2
8 15 3 13 16 1 0 9 2
26 1 9 7 0 13 13 12 2 3 9 15 2 7 9 15 2 15 3 13 15 9 2 16 13 4 2
8 15 7 9 13 9 9 13 2
10 15 3 9 13 1 15 16 9 13 2
13 13 3 16 1 15 13 9 13 9 9 7 9 2
2 0 2
10 15 13 15 1 9 2 13 13 9 2
7 9 3 13 13 15 9 2
27 13 4 7 1 16 10 15 9 13 9 1 0 9 2 7 1 15 15 9 13 13 16 9 1 15 13 2
11 15 3 9 13 9 13 16 15 9 15 2
9 15 7 15 9 13 2 9 13 2
10 3 9 2 16 3 2 1 9 13 2
10 1 15 3 9 13 13 9 7 9 2
2 3 2
13 10 13 15 13 1 15 15 13 16 9 1 9 2
10 1 15 3 15 13 13 13 9 15 2
18 13 7 4 1 16 0 9 13 0 9 2 10 7 15 13 15 9 2
13 13 3 9 10 13 1 10 9 16 9 1 9 2
2 3 2
9 9 15 1 9 13 13 1 9 2
9 9 3 13 15 0 16 13 9 2
17 9 7 15 9 13 1 9 13 1 15 9 2 16 1 13 4 2
12 15 3 9 13 1 10 9 13 16 9 15 2
14 1 15 13 16 1 15 9 13 13 9 9 7 9 2
15 16 3 13 15 13 1 9 7 9 2 7 9 7 9 2
25 3 13 7 15 9 9 1 9 7 9 2 7 1 9 7 9 2 16 15 13 1 9 7 9 2
29 0 3 2 16 9 3 13 15 9 9 2 3 13 10 9 13 9 2 16 0 0 13 2 7 9 13 9 9 2
15 0 7 16 15 9 3 13 0 9 9 2 7 9 15 2
12 15 3 9 13 9 1 15 13 13 16 13 2
11 9 7 3 13 1 9 2 7 1 15 2
16 3 9 3 13 13 15 13 2 7 15 9 13 15 15 13 2
15 0 2 16 7 9 13 15 9 2 7 15 13 1 9 2
17 13 3 9 1 15 9 16 9 1 13 2 7 9 1 0 13 2
12 3 16 1 15 3 9 13 15 9 16 9 2
39 1 15 3 1 9 1 9 7 9 13 9 13 9 13 2 16 13 9 9 2 15 9 13 15 9 2 16 0 13 9 9 13 3 13 15 0 9 9 2
22 3 1 9 1 9 7 9 7 9 7 9 13 13 15 15 13 2 7 3 15 9 2
13 9 3 13 13 15 13 2 1 16 13 13 9 2
18 15 7 15 9 13 15 15 13 2 7 15 9 13 15 9 13 9 2
41 1 9 7 0 2 15 3 13 1 9 7 9 13 2 16 13 4 2 7 1 15 15 9 13 9 0 2 9 13 15 13 2 15 7 9 13 9 7 15 13 2
39 7 1 15 1 15 13 0 3 9 9 7 9 2 15 3 13 1 9 7 9 2 15 1 15 13 1 15 13 7 9 2 7 1 15 13 7 15 13 2
15 1 9 7 13 1 9 7 9 13 0 9 9 7 9 2
12 0 3 15 9 2 15 13 1 9 7 9 2
28 0 0 1 15 9 3 13 7 9 2 15 3 13 13 1 15 13 7 9 2 7 1 15 13 7 15 13 2
17 3 3 13 16 9 9 7 9 13 1 0 16 9 9 7 9 2
8 3 9 7 9 13 9 0 2
8 9 7 7 9 13 9 0 2
29 7 1 15 15 3 13 9 7 9 16 3 2 13 0 9 0 7 0 13 2 16 13 7 13 2 13 7 13 2
32 15 0 13 0 9 7 9 16 3 2 16 13 7 13 7 15 3 2 15 13 0 9 0 2 7 15 9 13 9 0 13 2
6 16 9 0 13 0 2
12 1 15 7 13 13 16 10 9 0 13 0 2
10 10 3 9 13 1 9 9 1 9 2
8 0 3 9 1 9 9 0 2
9 9 7 1 15 1 9 9 0 2
8 9 3 13 2 13 9 13 2
12 1 9 3 9 13 0 0 15 15 13 9 2
16 3 7 3 13 9 9 7 9 2 3 3 13 13 9 15 2
4 3 7 9 2
14 13 4 7 16 15 9 0 13 13 1 9 7 9 2
7 15 3 9 0 13 0 2
2 0 2
28 15 1 15 15 13 2 1 9 7 3 7 0 15 13 2 16 0 1 15 3 13 9 2 1 9 7 9 2
17 3 9 3 13 3 0 13 0 2 9 7 3 13 0 13 0 2
8 9 7 1 15 13 1 9 2
8 1 15 3 13 1 16 15 2
9 15 7 13 9 1 16 13 9 2
27 9 3 15 3 13 15 9 2 13 13 9 2 1 16 13 9 2 16 9 13 9 1 16 13 13 0 2
26 9 0 15 13 15 9 2 3 13 13 9 2 16 2 16 15 9 13 9 2 3 13 13 3 0 2
12 13 4 7 1 16 9 0 13 15 9 0 2
7 0 13 3 16 13 13 2
4 13 3 0 2
2 3 2
10 1 10 9 2 13 9 2 13 9 2
18 3 3 13 15 1 3 3 9 2 16 7 13 15 1 3 3 9 2
21 1 9 7 0 2 16 13 4 2 9 13 15 9 2 15 7 9 13 16 9 2
11 16 3 9 0 13 2 13 1 10 9 2
5 15 13 3 0 2
7 10 3 9 0 13 0 2
2 3 2
13 1 10 15 13 2 13 16 13 9 1 3 9 2
19 16 15 3 13 1 15 3 13 9 1 3 9 2 15 3 13 13 0 2
11 1 9 7 0 3 13 9 1 3 9 2
14 0 13 3 1 13 16 9 0 13 0 0 15 9 2
40 0 7 0 15 9 3 13 16 9 1 9 15 16 15 9 13 1 9 1 13 2 16 9 3 13 1 9 16 9 1 9 16 15 9 13 1 9 1 9 2
19 3 7 1 15 9 0 13 9 1 3 9 1 15 9 0 16 9 9 2
15 1 9 7 0 3 13 9 2 7 15 13 9 0 0 2
10 3 1 15 3 13 9 1 3 9 2
4 13 3 0 2
2 3 2
22 1 15 13 9 9 7 9 2 15 15 13 9 0 9 2 7 0 9 2 13 0 2
10 3 3 1 9 0 9 0 13 0 2
19 7 1 9 0 15 15 13 9 0 9 7 9 2 13 15 15 9 0 2
6 3 9 15 13 0 2
12 15 7 13 0 16 1 15 16 10 9 13 2
7 3 10 0 9 13 0 2
2 0 2
13 10 15 13 7 13 1 15 2 7 13 1 9 2
9 9 7 0 3 13 1 15 13 2
7 10 3 9 13 1 0 2
19 9 3 2 1 13 1 16 13 9 9 2 3 13 13 1 15 13 9 2
23 3 2 16 1 3 13 9 15 13 13 13 9 2 13 16 15 13 1 9 15 1 3 2
8 3 0 13 15 0 15 13 2
20 7 1 15 13 10 15 13 1 15 2 7 13 0 2 7 13 1 0 13 2
7 15 7 15 9 0 13 2
20 15 9 13 2 16 1 9 15 3 15 1 10 9 13 0 2 13 13 0 2
10 0 3 7 0 1 9 3 13 0 2
18 3 3 15 13 2 3 3 15 13 2 1 9 3 12 15 13 15 2
9 9 3 0 3 13 0 1 15 2
6 0 7 7 1 9 2
9 3 3 13 9 7 9 3 0 2
10 13 7 4 1 16 9 0 13 0 2
5 13 3 3 0 2
2 3 2
5 9 13 9 15 2
12 15 13 13 9 9 2 16 1 9 4 13 2
8 3 13 16 10 15 13 13 2
12 13 4 7 1 0 16 10 15 13 13 9 2
28 13 3 10 15 13 13 9 2 16 1 15 13 2 7 15 9 7 9 9 1 9 13 2 16 13 1 9 2
15 9 7 0 3 13 9 2 7 9 7 9 1 9 13 2
9 3 7 1 15 7 1 9 13 2
5 13 3 3 0 2
2 3 2
11 10 15 13 2 13 1 15 16 15 13 2
8 3 7 15 13 13 15 13 2
13 15 7 9 0 13 13 15 9 15 13 1 9 2
6 3 13 13 15 13 2
19 15 7 13 1 9 0 2 13 16 13 1 15 1 9 15 2 3 0 2
18 15 0 3 1 9 0 13 2 13 13 9 0 2 7 3 13 15 2
6 0 3 13 9 13 2
6 9 3 13 13 0 2
2 3 2
12 16 0 13 9 9 2 3 0 13 9 9 2
29 9 7 0 9 3 13 16 1 9 10 9 2 16 9 1 3 0 2 7 9 1 0 0 2 7 3 1 15 2
15 13 7 0 9 2 16 9 13 3 1 9 1 9 9 2
25 15 3 9 9 3 13 13 9 2 1 3 13 9 9 15 3 1 9 13 2 16 1 13 4 2
25 13 7 16 7 13 1 9 10 9 2 16 15 13 3 0 2 3 0 13 0 0 2 7 3 2
7 9 3 15 9 13 0 2
2 0 2
6 0 13 0 9 9 2
11 3 9 1 9 7 0 1 9 13 12 2
22 15 3 13 0 16 13 0 2 13 13 9 16 3 2 16 9 7 0 13 12 9 2
12 0 7 2 16 13 0 2 13 0 7 0 2
7 0 3 9 13 9 0 2
10 13 0 2 16 3 2 3 16 13 2
10 13 3 1 15 3 9 2 7 9 2
16 3 7 0 9 9 13 1 16 13 0 2 16 3 13 0 2
6 13 3 9 13 0 2
2 3 2
7 15 13 1 9 10 9 2
12 1 9 3 9 15 9 13 13 9 9 15 2
16 9 7 3 13 1 9 2 7 1 15 16 13 1 9 13 2
26 13 3 1 0 9 9 7 9 2 13 9 7 0 7 9 9 2 16 13 1 9 2 1 12 9 2
18 9 3 9 13 13 16 9 10 13 1 9 2 7 1 13 1 9 2
10 9 7 15 9 0 13 9 7 9 2
8 0 13 3 9 13 13 0 2
2 3 2
7 0 13 0 9 13 0 2
6 9 3 15 13 3 2
20 7 15 13 0 13 9 0 2 3 0 16 13 13 1 9 2 7 3 9 2
4 15 3 13 2
25 0 3 9 15 3 13 1 9 2 16 9 0 13 9 9 1 15 13 2 7 9 0 13 9 2
24 15 0 1 9 2 1 0 9 0 9 2 15 0 9 1 15 13 2 16 0 13 13 3 2
9 15 7 9 13 9 0 9 13 2
31 15 9 13 16 7 15 15 9 13 2 13 13 1 9 10 9 0 2 7 15 15 9 13 2 13 15 1 9 10 9 2
29 15 3 9 9 15 9 13 9 1 13 9 0 3 16 13 3 15 1 9 2 0 13 9 0 3 1 15 9 2
25 15 7 9 3 13 1 15 9 2 7 0 1 13 9 0 1 15 9 2 3 3 0 13 9 2
41 15 3 9 13 7 1 15 13 15 9 13 1 9 13 2 16 3 15 15 3 13 9 16 16 3 2 13 9 16 3 2 3 7 3 2 16 9 0 3 13 2
27 13 3 13 0 9 2 3 1 9 2 16 9 0 2 15 1 15 13 2 0 13 2 7 3 13 9 2
15 15 3 15 15 9 0 13 7 13 2 13 15 0 9 2
7 15 7 13 10 9 13 2
10 10 3 9 13 0 9 13 13 3 2
7 3 0 13 16 13 13 2
2 3 2
12 15 13 13 7 13 2 1 15 9 13 15 2
11 15 3 13 9 1 9 7 1 3 9 2
13 7 9 13 3 13 13 13 16 1 9 0 9 2
14 3 3 13 1 9 2 15 13 13 2 16 13 4 2
22 3 7 13 15 9 1 3 9 15 16 1 0 9 2 1 16 13 3 13 15 9 2
10 7 1 15 0 9 15 13 13 0 2
25 3 16 9 13 0 7 13 1 9 15 13 1 15 2 7 3 1 9 9 2 16 1 13 4 2
20 3 3 16 9 2 15 13 9 9 2 3 13 9 15 15 13 0 9 15 2
12 13 4 7 16 0 9 0 13 16 13 0 2
8 3 15 15 1 9 3 13 2
9 13 3 9 0 1 10 9 0 2
19 15 13 15 1 9 2 13 9 1 9 2 13 9 7 0 9 2 13 2
15 13 15 1 0 7 1 9 9 2 1 15 13 9 13 2
52 9 3 2 1 12 8 1 8 8 2 13 16 1 0 9 9 13 0 7 0 9 2 7 13 7 13 2 7 13 9 0 7 0 2 1 0 9 7 9 7 9 9 13 2 7 13 1 0 7 13 9 2
9 1 15 9 9 0 13 9 13 2
27 1 7 1 13 4 9 0 3 13 9 7 9 15 1 9 13 2 13 13 3 15 9 0 9 13 13 2
15 13 7 0 0 16 9 0 3 13 9 13 1 9 9 2
10 15 3 13 2 13 1 3 13 13 2
20 15 3 13 16 1 15 15 13 9 15 2 15 13 13 0 7 0 1 3 2
10 9 7 0 3 13 1 9 1 0 2
9 13 3 0 2 16 1 13 4 2
6 3 13 3 9 0 2
2 3 2
15 15 13 2 9 3 13 2 3 13 9 2 7 9 3 2
13 3 16 9 13 2 3 13 9 2 7 9 3 2
9 3 9 13 1 9 15 15 13 2
8 15 7 0 13 13 9 0 2
9 13 3 0 2 16 1 13 4 2
11 3 3 13 9 0 13 9 1 9 9 2
16 0 7 13 16 9 0 3 13 13 9 1 9 9 0 13 2
7 9 3 3 16 9 13 2
20 13 3 13 15 13 0 3 2 16 9 7 9 7 9 2 15 13 9 0 2
11 3 3 1 9 9 9 0 9 13 13 2
22 1 15 7 13 16 7 9 2 7 9 7 9 2 1 9 0 7 9 12 13 13 2
9 10 3 15 1 9 13 3 13 2
12 13 3 15 9 9 15 9 0 9 13 13 2
34 9 3 0 13 15 13 2 7 3 1 3 13 3 0 1 0 9 2 7 3 1 9 9 7 9 2 16 13 9 10 13 1 13 2
35 7 16 2 16 13 0 0 9 2 13 1 10 0 13 9 2 3 2 16 13 1 9 7 9 2 13 15 13 13 3 7 15 13 3 2
14 9 3 0 13 3 15 9 0 9 2 16 15 13 2
12 3 7 13 1 15 2 16 1 15 3 13 2
18 16 3 13 15 9 15 9 0 3 13 2 13 3 13 2 16 13 2
9 1 15 9 13 16 13 15 13 2
13 15 3 9 13 0 13 13 9 0 9 1 9 2
19 13 3 9 0 1 9 7 13 15 2 1 13 0 7 3 1 9 13 2
10 15 7 9 3 13 9 2 7 9 2
10 3 13 15 9 1 9 0 1 12 2
14 0 3 2 16 15 9 15 15 13 0 13 13 0 2
8 15 1 9 0 3 13 13 2
9 3 9 3 13 13 16 0 15 2
18 9 7 0 2 16 13 0 2 13 13 9 0 2 16 13 1 15 2
11 15 3 9 13 0 9 2 7 9 0 2
20 9 3 16 9 9 2 7 3 13 9 13 1 0 2 1 15 13 3 13 2
11 9 7 0 13 0 3 1 9 9 13 2
10 3 3 13 15 0 15 9 1 13 2
10 0 2 16 9 9 13 0 1 0 2
9 9 7 9 13 1 15 15 13 2
9 3 3 13 1 16 13 7 13 2
9 15 7 13 1 16 13 1 9 2
11 9 0 13 1 15 2 3 1 0 15 2
4 3 15 13 2
6 1 15 13 0 9 2
30 16 1 9 9 2 15 13 1 0 2 13 13 13 0 15 15 13 2 7 3 13 13 1 15 2 7 13 1 15 2
30 9 7 9 2 15 13 9 0 2 1 13 1 0 2 13 9 13 13 1 15 15 13 2 7 13 1 15 1 9 2
11 3 3 9 0 13 9 13 1 9 9 2
12 15 7 13 1 15 9 2 3 13 12 0 2
8 13 3 12 1 13 7 13 2
7 15 3 13 13 12 0 2
8 3 3 13 12 3 7 9 2
8 13 7 9 3 13 13 0 2
11 3 7 13 12 1 13 13 13 12 0 2
21 12 7 0 0 13 2 7 16 0 2 7 16 0 2 7 16 15 13 9 12 2
14 1 9 7 0 7 9 3 13 13 12 15 13 0 2
8 13 3 15 13 13 1 12 2
12 7 3 16 13 0 2 16 9 0 15 13 2
19 13 3 13 3 1 9 0 7 9 13 3 13 12 16 15 13 9 12 2
17 1 12 7 13 3 13 15 9 12 16 16 1 9 0 7 9 2
10 1 9 3 7 9 3 13 9 12 2
9 3 3 13 15 9 9 7 0 2
15 15 3 13 13 2 3 9 0 9 15 9 0 13 13 2
8 13 7 0 13 15 13 0 2
12 1 12 3 9 9 13 3 13 13 15 12 2
10 9 3 15 13 15 15 1 15 13 2
13 9 7 0 13 9 9 13 2 16 1 13 13 2
5 0 7 7 9 2
16 3 3 13 15 12 13 2 16 13 2 1 9 0 7 9 2
2 3 2
8 9 7 9 1 15 9 13 2
9 10 3 9 1 9 7 9 13 2
9 9 7 0 7 9 13 0 9 2
9 3 3 13 0 12 13 9 15 2
2 0 2
12 10 15 15 9 13 1 9 2 13 13 0 2
17 7 16 9 0 13 9 9 2 13 16 9 15 13 1 9 0 2
9 3 3 9 9 13 1 9 9 2
14 13 3 16 9 0 3 13 0 2 16 1 13 4 2
2 3 2
14 0 13 15 15 9 13 1 9 2 13 1 9 13 2
20 9 7 13 1 9 13 13 1 9 2 7 16 7 13 9 7 9 1 9 2
8 3 13 3 0 9 9 9 2
8 3 3 9 15 13 1 9 2
2 3 2
13 15 9 13 0 9 2 13 7 9 9 0 13 2
25 15 3 13 1 16 13 9 2 7 9 0 9 13 13 0 16 15 9 2 1 9 9 9 13 2
18 16 7 9 0 13 9 9 2 13 16 9 15 13 15 7 9 0 2
16 1 9 3 7 9 13 15 12 0 2 15 13 1 9 12 2
16 13 3 7 9 9 0 0 9 2 7 9 15 9 1 9 2
7 15 1 13 13 13 0 2
9 9 9 1 13 9 0 1 9 2
19 1 15 7 7 0 9 15 13 2 13 16 15 9 0 13 13 9 9 2
29 7 16 15 9 15 9 9 13 13 2 15 1 9 0 7 9 13 13 13 2 13 15 9 1 15 9 9 13 2
34 9 3 13 2 7 15 0 2 16 9 0 3 13 9 16 9 9 2 7 0 16 9 0 2 13 9 13 1 9 16 9 1 9 2
19 7 3 13 9 7 9 3 13 16 1 9 9 2 1 15 1 13 4 2
5 15 7 13 9 2
14 1 13 3 9 3 13 15 12 0 2 16 13 4 2
9 1 13 7 9 7 9 13 9 2
21 13 3 16 9 3 13 12 0 2 7 1 13 7 9 0 2 7 9 1 9 2
43 1 15 7 13 2 9 13 16 9 3 13 15 13 1 9 7 9 2 7 16 15 9 13 9 13 9 2 16 9 3 13 15 13 1 9 7 9 2 7 9 13 9 2
6 15 7 13 0 13 2
10 9 3 7 9 13 15 0 7 0 2
28 15 7 3 13 16 9 7 15 9 3 13 1 9 9 7 9 2 7 15 9 15 13 9 2 1 9 13 2
9 9 3 3 13 15 0 7 0 2
20 0 13 3 9 7 9 13 9 13 9 2 3 7 15 1 9 7 9 13 2
2 3 2
14 0 13 16 15 15 13 0 1 9 2 13 9 12 2
21 13 7 9 12 2 3 1 9 15 1 15 13 9 2 7 1 16 13 1 9 2
52 0 3 13 9 12 9 13 1 9 13 2 15 13 12 2 7 3 1 9 13 13 0 9 2 16 13 0 9 1 13 2 1 3 9 13 9 7 9 2 13 15 13 0 9 7 9 2 13 7 9 0 2
35 16 7 9 13 15 9 0 2 1 15 3 13 9 2 16 13 2 13 3 15 9 0 15 7 9 2 16 13 7 13 7 13 7 3 2
22 15 3 13 1 15 9 15 13 9 9 2 1 15 13 16 3 13 9 7 9 9 2
17 13 3 1 9 7 9 12 13 2 7 16 3 13 1 9 0 2
8 15 7 9 1 9 9 13 2
17 15 3 9 13 13 7 13 2 16 1 9 0 2 13 15 9 2
18 3 9 13 15 9 13 16 1 15 13 2 13 7 16 1 15 13 2
22 3 3 9 13 13 9 13 9 9 7 0 16 3 13 9 16 13 7 9 16 13 2
6 7 15 13 3 13 2
19 16 2 16 13 9 1 12 1 9 2 13 13 1 15 13 1 0 0 2
17 3 3 13 9 13 1 0 0 2 16 3 13 15 13 1 13 2
14 9 3 9 13 7 13 1 13 2 7 1 0 0 2
23 15 7 15 13 13 9 2 15 1 15 13 2 16 13 9 3 13 1 0 15 9 9 2
8 9 3 13 9 0 15 9 2
20 9 3 0 3 15 13 1 13 16 13 7 9 2 7 16 15 15 0 13 2
10 15 0 13 13 0 1 9 1 0 2
12 3 13 3 9 0 1 9 0 1 9 13 2
2 3 2
19 16 9 13 0 9 13 7 13 2 3 15 9 13 13 9 7 13 9 2
9 3 7 12 9 13 13 7 13 2
23 16 3 1 13 9 0 15 13 16 9 7 9 16 0 2 15 13 9 9 7 15 9 2
8 9 3 0 13 15 9 0 2
6 13 3 7 9 0 2
9 3 3 2 13 9 2 13 13 2
11 9 3 0 2 3 0 9 2 13 0 2
5 15 3 0 13 2
15 3 1 9 9 3 13 2 7 1 15 1 13 9 13 2
2 0 2
8 0 3 13 9 1 10 9 2
21 16 3 9 3 13 9 16 16 9 0 2 9 7 9 15 3 13 9 1 9 2
12 13 3 9 2 13 9 7 9 15 15 9 2
6 15 7 13 0 0 2
29 3 9 7 9 7 9 7 3 9 1 9 9 3 13 16 0 2 1 15 15 9 0 9 13 2 15 9 13 2
15 3 3 13 9 9 0 16 9 0 2 7 16 9 9 2
2 3 2
12 0 3 13 9 1 10 9 2 7 3 9 2
22 16 3 9 13 9 3 16 9 2 9 13 3 1 9 2 7 3 13 9 1 15 2
7 13 7 13 15 9 13 2
7 3 3 9 13 1 9 2
2 3 2
29 0 7 13 1 9 9 1 15 2 7 1 15 9 13 2 1 3 13 0 1 9 1 9 2 7 1 13 3 2
26 16 3 9 13 9 0 16 9 2 13 16 1 13 9 7 9 3 13 15 9 2 7 1 9 9 2
17 7 3 9 2 15 13 1 9 9 7 9 2 3 13 9 0 2
5 15 13 0 0 2
2 3 2
21 10 13 15 3 15 13 16 1 15 13 13 7 3 13 2 7 13 7 3 13 2
13 7 9 2 1 9 9 2 13 9 16 13 15 2
11 13 3 1 9 9 13 9 7 3 13 2
27 16 3 3 13 15 16 16 9 0 2 13 1 9 9 13 1 9 1 13 2 7 3 13 15 1 13 2
5 15 13 13 0 2
12 16 7 16 9 0 9 9 13 2 3 13 2
16 15 15 15 13 1 9 9 9 9 2 13 9 7 9 15 2
11 9 7 1 9 13 9 9 1 9 13 2
6 13 3 13 9 13 2
17 9 7 1 9 13 13 0 1 9 2 1 9 7 13 13 9 2
7 13 3 9 9 9 13 2
2 0 2
34 16 3 13 7 3 13 3 13 0 9 7 0 9 2 7 13 2 13 7 13 12 13 2 15 12 15 13 1 15 16 9 1 9 2
30 13 3 16 9 13 0 9 7 9 2 7 16 13 13 9 7 9 2 15 9 13 9 9 13 2 7 9 9 0 2
9 13 7 7 13 13 9 7 9 2
10 13 3 7 13 7 13 9 7 9 2
9 7 9 3 16 9 9 7 9 2
6 13 3 9 9 9 2
2 3 2
14 0 15 13 15 9 0 1 15 9 16 9 1 9 2
14 9 7 3 15 13 1 9 16 13 9 7 9 15 2
8 9 3 13 9 7 9 9 2
8 3 9 13 9 7 9 9 2
13 16 0 2 0 7 0 3 13 1 9 12 9 2
14 13 7 13 9 1 9 9 13 3 1 13 9 13 2
15 13 3 9 3 13 15 9 1 15 0 2 0 7 0 2
23 3 2 16 9 0 13 9 9 2 3 13 1 15 13 16 15 0 9 9 9 13 13 2
10 16 7 15 13 0 2 3 13 13 2
14 15 13 15 15 1 0 9 2 13 1 3 1 9 2
15 0 3 13 13 0 1 9 2 16 9 13 9 7 0 2
30 16 3 9 0 2 0 7 0 13 0 9 7 9 1 15 2 15 15 1 15 9 15 13 2 1 3 13 1 9 2
15 7 1 9 0 13 9 2 1 0 9 2 1 0 13 2
17 13 3 15 9 1 9 2 9 13 9 2 7 2 9 13 0 2
5 13 7 1 15 2
20 3 9 1 16 13 9 2 9 13 2 7 9 1 16 13 9 2 0 13 2
12 13 3 15 1 15 9 9 2 0 7 0 2
32 16 7 13 16 2 3 13 9 0 13 2 3 13 13 9 13 1 9 2 15 16 9 15 1 3 9 13 2 15 3 13 2
18 3 9 0 1 0 2 7 0 1 0 2 13 16 9 9 1 9 2
12 3 0 0 2 7 0 0 0 1 9 13 2
9 0 3 1 9 13 9 16 9 2
40 16 3 15 9 13 9 13 13 1 15 2 15 3 13 1 15 9 13 1 15 15 13 1 9 2 7 1 15 15 13 1 9 7 9 2 16 13 9 13 2
5 15 7 13 0 2
32 16 1 15 9 13 1 15 2 15 15 13 0 13 1 15 1 9 2 16 1 13 2 9 13 0 2 7 2 9 13 0 2
20 7 3 1 15 9 13 1 15 9 13 1 9 9 2 16 9 1 9 0 2
6 3 7 1 0 13 2
26 3 3 9 1 15 13 1 9 2 7 1 0 2 7 3 3 13 9 1 9 9 2 7 1 0 2
11 3 3 13 9 13 1 15 9 13 9 2
2 3 2
8 1 15 15 13 9 7 9 2
6 12 3 13 1 9 2
15 1 3 1 9 15 9 13 9 2 1 9 3 13 9 2
20 16 3 13 1 9 0 9 16 0 9 2 9 3 13 12 9 2 7 0 2
8 7 1 9 9 9 9 13 2
18 16 13 12 1 9 3 13 13 12 0 2 1 9 9 13 0 9 2
2 3 2
22 3 13 13 9 2 16 3 1 9 0 7 9 3 13 12 0 2 7 1 9 3 2
19 10 3 15 13 15 1 13 0 2 13 15 0 2 1 13 1 9 15 2
11 15 7 9 0 13 9 0 1 9 9 2
8 13 3 9 9 7 15 15 2
12 15 3 1 0 9 0 13 9 2 0 13 2
29 1 3 9 0 13 9 0 2 0 3 0 1 9 13 7 1 9 2 13 16 9 0 13 0 2 7 0 0 2
19 7 3 7 9 7 9 13 12 0 2 7 15 9 7 9 1 9 9 2
2 0 2
44 16 9 2 1 9 9 2 3 13 15 1 9 7 9 13 2 7 13 9 13 9 2 7 15 13 0 1 9 0 2 7 1 12 9 2 16 12 13 2 7 1 12 15 2
20 16 7 1 12 7 12 2 13 16 9 3 13 12 2 7 13 12 7 12 2
9 13 3 12 9 2 7 3 12 2
64 16 7 15 13 1 9 0 3 2 3 3 16 13 9 0 13 9 9 2 7 9 0 13 9 13 7 13 13 9 2 13 3 9 2 3 16 9 3 13 9 2 7 13 9 2 3 1 9 0 15 13 9 2 7 16 9 3 13 2 7 13 9 13 2
21 15 1 13 9 2 0 13 12 9 9 13 13 1 15 2 0 2 0 7 0 2
2 3 2
26 1 12 7 0 3 13 13 12 16 3 13 15 13 2 16 12 15 15 13 1 15 16 9 1 9 2
15 3 3 1 9 7 9 13 12 2 15 9 0 15 13 2
28 16 7 1 9 13 0 9 2 3 15 13 1 3 16 9 7 9 2 7 10 13 16 9 15 7 9 9 2
20 13 3 2 16 13 1 13 15 12 2 13 9 7 9 2 16 13 15 13 2
24 15 7 3 13 13 9 2 1 3 9 13 1 9 2 15 9 13 16 13 9 2 9 13 2
14 13 3 16 13 15 0 13 15 13 1 15 0 12 2
13 7 15 3 13 9 16 15 0 15 1 15 13 2
22 16 3 15 3 13 13 9 0 2 7 3 13 12 1 15 2 13 3 13 15 13 2
18 1 3 3 13 13 1 0 2 13 13 1 15 15 13 1 15 12 2
6 7 15 0 13 9 2
12 13 3 1 12 9 7 9 12 3 9 13 2
2 3 2
33 16 15 15 13 1 9 9 1 9 2 13 1 0 13 2 13 16 16 15 13 15 13 1 15 9 2 3 0 1 0 9 9 2
8 15 3 1 9 9 3 13 2
15 13 3 9 0 1 9 2 0 1 9 2 0 1 9 2
8 15 7 13 13 0 2 0 2
31 0 3 16 15 9 9 13 15 3 13 13 15 9 9 2 3 9 2 1 15 1 13 4 16 3 13 9 15 9 9 2
48 0 2 16 0 13 16 1 15 9 9 13 0 9 9 9 2 16 13 1 9 15 13 13 2 16 15 9 13 9 7 9 7 9 15 13 2 7 0 15 9 9 13 13 2 13 7 13 2
15 1 15 13 16 0 9 9 1 12 7 15 9 9 13 2
13 3 3 13 0 9 1 15 2 0 9 9 13 2
2 0 2
23 0 9 15 3 13 1 12 9 2 3 13 15 3 1 13 2 16 9 15 9 13 0 2
6 15 1 13 3 13 2
9 13 7 16 0 9 9 13 15 2
9 1 3 12 13 13 2 15 13 2
19 13 3 16 15 9 2 7 9 15 13 15 0 9 2 13 1 12 9 2
46 15 7 9 3 13 13 9 2 3 16 15 9 13 1 15 3 13 9 2 3 13 2 7 16 2 16 9 15 9 7 9 13 9 16 3 2 13 1 10 9 2 15 13 13 0 2
19 7 3 13 16 13 9 15 9 15 12 2 1 15 15 9 13 15 9 2
4 15 13 9 2
16 13 3 16 10 9 9 15 13 1 15 2 1 9 12 13 2
9 7 3 3 13 1 15 0 9 2
11 15 7 13 15 13 1 9 1 8 9 2
58 7 12 9 13 13 1 12 9 2 16 9 7 15 9 13 2 12 0 2 15 13 9 2 7 13 4 9 2 7 15 0 2 15 9 13 2 7 13 12 15 7 13 9 1 9 15 7 9 10 9 13 2 7 15 10 9 13 2
9 16 9 0 9 3 13 9 13 2
19 13 7 7 15 15 9 13 1 13 16 9 0 3 13 13 9 16 9 2
21 13 3 16 9 2 3 15 9 0 13 2 13 15 9 13 3 13 15 16 9 2
32 7 15 13 13 2 0 2 1 9 9 15 13 2 1 15 9 13 2 16 13 13 2 7 0 9 2 7 0 2 7 0 2
11 15 3 13 13 1 15 16 13 9 9 2
29 3 2 1 9 15 15 13 16 2 16 9 0 13 10 9 9 0 16 1 9 1 15 13 2 13 16 10 13 2
13 16 9 2 15 13 10 9 9 2 13 10 9 2
15 16 3 13 1 15 15 9 2 15 9 13 13 15 9 2
8 3 15 13 16 1 15 9 2
19 7 0 13 1 9 0 2 16 13 1 15 15 9 7 9 1 9 0 2
11 15 7 13 13 2 16 13 13 15 9 2
30 7 0 16 13 9 15 9 2 16 2 1 1 9 7 9 13 12 2 13 16 9 13 15 1 9 15 15 13 9 2
17 0 13 3 9 0 13 13 9 2 7 13 9 7 9 15 9 2
2 3 2
19 16 13 9 15 9 0 2 13 15 9 9 15 9 2 7 9 9 0 2
15 15 3 15 13 15 9 9 2 3 13 15 1 10 9 2
7 9 7 0 13 9 0 2
9 3 1 15 13 16 13 1 9 2
9 9 3 0 13 9 16 13 0 2
6 7 3 3 13 0 2
5 15 13 13 0 2
2 3 2
9 9 0 3 13 0 9 15 13 2
18 16 3 15 13 9 9 0 7 9 0 2 7 9 0 13 9 13 2
4 15 13 0 2
2 0 2
16 0 13 1 9 13 9 0 2 16 13 1 9 1 12 8 2
8 9 7 0 13 3 9 0 2
23 13 3 1 15 9 0 1 9 2 16 1 15 13 0 2 1 15 13 0 0 1 9 2
9 3 13 3 9 0 9 1 9 2
36 1 15 7 13 4 9 7 15 0 2 16 15 13 2 1 13 9 0 2 15 13 9 2 13 13 1 9 1 9 2 7 3 13 9 9 2
47 7 16 15 9 15 1 15 13 2 7 1 15 13 2 16 15 15 9 13 2 13 3 9 15 13 15 2 13 16 9 13 1 9 13 9 9 0 2 16 0 1 9 13 9 9 0 2
12 3 1 9 0 7 9 13 1 9 13 12 2
11 15 3 13 9 13 13 2 13 9 0 2
14 13 7 15 13 9 2 15 13 9 15 15 9 13 2
10 1 15 3 9 3 9 0 15 13 2
11 16 7 15 0 13 7 0 0 13 13 2
6 13 3 9 13 13 2
9 13 7 15 15 9 0 9 13 2
30 1 15 3 16 9 0 9 13 4 1 9 1 15 9 2 3 13 9 16 13 13 2 7 0 16 13 1 9 13 2
2 3 2
24 3 9 13 1 9 13 9 9 0 2 16 9 0 1 9 13 9 9 0 2 7 15 9 2
28 9 7 13 13 1 9 16 9 0 1 9 1 13 15 13 1 9 2 7 15 9 15 13 2 7 3 9 2
26 0 3 9 13 9 0 1 9 0 1 9 15 1 15 13 2 7 9 0 1 9 15 13 1 9 2
12 15 7 9 3 13 9 13 2 7 0 13 2
16 3 7 13 9 9 0 15 3 13 15 13 2 7 13 0 2
12 0 7 13 16 0 7 0 13 16 9 13 2
12 3 3 9 9 13 16 1 15 16 15 13 2
8 3 3 0 13 13 9 9 2
2 3 2
23 10 13 1 9 0 13 9 2 7 3 1 0 2 16 7 13 10 1 9 0 13 13 2
11 9 7 13 13 1 9 16 1 9 0 2
14 3 3 13 1 9 0 9 2 7 3 1 9 0 2
2 0 2
10 15 15 15 13 2 13 13 9 15 2
9 15 3 13 16 1 16 13 9 2
13 9 7 3 13 15 16 1 15 15 13 9 15 2
18 3 7 9 13 9 13 9 2 1 15 16 9 1 9 13 7 13 2
10 9 7 13 2 7 3 16 1 9 2
16 3 7 9 2 13 1 9 15 13 2 13 15 9 9 0 2
15 13 3 9 0 0 13 15 2 7 3 0 1 10 9 2
2 3 2
19 9 1 9 7 0 1 9 13 12 2 16 9 1 9 7 0 1 9 2
20 3 7 9 1 9 7 0 1 9 2 16 7 9 1 9 7 0 1 9 2
15 9 3 9 2 1 16 13 1 9 2 3 13 0 9 2
39 3 3 3 13 12 1 9 1 9 7 1 16 13 1 9 13 2 16 7 9 9 13 0 1 9 1 16 13 1 9 2 7 0 1 16 13 1 9 2
17 3 7 0 13 15 9 0 1 16 13 1 9 2 1 9 13 2
15 3 3 13 15 1 16 13 12 1 9 0 16 9 15 2
27 3 3 13 13 0 15 13 9 0 15 2 16 1 16 13 1 9 0 2 3 13 15 2 7 1 0 2
12 13 7 15 15 15 9 13 2 9 13 4 2
32 9 3 1 9 13 2 13 9 2 13 0 9 16 13 13 9 2 3 7 16 9 0 2 1 16 13 12 1 9 1 9 2
35 7 0 9 1 9 9 13 13 9 0 2 16 13 13 9 0 2 3 7 16 4 13 9 2 1 16 13 12 1 9 0 13 1 9 2
2 3 2
16 16 13 9 9 13 2 3 13 9 9 9 2 13 15 9 2
10 1 9 16 13 0 9 1 9 13 2
14 1 9 7 13 9 9 2 3 13 7 13 1 9 2
8 3 7 9 13 9 9 9 2
17 7 3 1 9 13 9 9 1 9 13 16 1 9 2 3 13 2
7 3 9 13 9 9 9 2
6 7 9 13 1 9 2
14 13 3 9 9 9 2 15 13 2 16 13 9 0 2
7 15 7 13 9 16 9 2
6 13 3 9 9 9 2
6 7 1 13 9 15 2
2 3 2
18 15 13 1 9 15 9 2 3 13 15 9 2 16 9 13 9 0 2
12 9 7 1 15 15 13 9 2 13 9 0 2
15 13 7 9 0 1 9 2 1 9 13 2 13 9 9 2
18 13 3 13 9 2 15 2 1 9 2 13 9 13 1 9 1 9 2
9 1 15 3 13 3 13 9 9 2
15 3 3 13 9 9 1 0 9 1 15 16 13 9 13 2
2 0 2
25 16 9 9 13 1 15 16 13 0 7 9 13 2 15 13 1 9 0 2 13 0 7 9 13 2
14 7 9 2 3 16 1 9 13 2 13 1 9 0 2
12 1 15 3 3 13 9 2 15 13 0 9 2
20 3 3 13 9 9 13 1 15 16 9 13 9 13 9 0 15 9 13 9 2
14 16 9 3 13 9 1 9 0 2 7 1 9 0 2
8 15 7 9 13 1 13 9 2
37 13 3 13 9 16 9 13 9 1 0 1 9 15 9 13 0 2 15 13 15 9 0 2 15 13 0 9 2 9 15 15 0 13 15 0 0 2
30 15 7 0 9 13 13 9 0 2 7 13 15 1 3 2 16 9 15 13 13 7 0 2 13 7 13 1 9 0 2
56 7 16 1 15 9 2 3 1 0 7 0 2 13 9 16 13 9 9 13 2 1 15 13 0 9 2 16 13 15 9 13 9 9 0 2 3 13 9 13 9 9 7 9 2 1 15 9 13 16 13 9 1 0 9 9 2
20 7 1 9 15 9 13 9 12 1 15 1 9 7 1 15 15 13 1 13 2
11 7 1 9 15 7 9 13 9 9 9 2
12 3 9 9 13 1 15 9 0 16 1 9 2
19 7 15 9 0 1 9 13 9 2 1 15 13 9 0 2 16 9 13 2
13 16 7 15 13 0 2 7 0 13 2 0 13 2
22 9 3 9 13 1 9 16 9 0 1 0 2 16 13 1 9 2 1 12 1 9 2
16 9 7 0 1 15 13 9 9 0 2 16 9 13 1 13 2
26 1 15 3 13 15 9 9 2 13 1 15 13 15 9 9 15 13 1 15 9 16 9 0 1 0 2
30 7 9 13 0 9 1 15 9 2 3 13 7 13 2 15 13 9 9 16 13 9 2 16 9 13 2 1 12 9 2
24 3 13 1 9 13 15 9 15 0 13 9 9 2 15 15 13 1 13 16 9 0 1 0 2
32 15 7 3 13 13 9 0 13 2 16 9 13 9 13 13 0 7 3 13 9 2 16 9 13 2 15 0 13 1 9 0 2
25 3 3 13 0 16 1 9 0 2 15 13 9 0 2 9 9 13 2 1 15 1 15 9 13 2
2 3 2
36 15 13 9 9 0 2 3 13 13 1 9 9 9 16 13 9 0 2 16 15 13 9 9 0 2 3 13 1 9 9 9 16 13 9 0 2
31 13 7 16 9 2 7 3 9 15 1 15 13 2 16 0 7 0 2 13 9 9 0 2 16 9 13 1 9 1 9 2
23 3 3 1 13 9 2 7 15 15 2 15 9 13 13 1 9 9 9 16 13 9 0 2
8 9 7 13 1 9 9 9 2
31 15 13 1 9 2 1 12 1 9 2 15 2 13 9 9 2 13 0 2 15 9 13 2 0 2 15 13 0 10 9 2
13 3 3 9 13 13 9 15 0 1 9 0 13 2
2 0 2
19 10 13 15 2 1 16 13 9 2 1 12 8 2 13 1 13 7 13 2
12 9 7 2 16 7 15 9 2 13 13 15 2
8 3 13 7 13 13 9 15 2
8 0 7 13 1 9 13 9 2
7 3 9 10 0 13 9 2
17 7 13 13 16 0 9 0 13 13 2 16 9 0 13 0 0 2
36 1 13 7 13 7 0 9 2 15 13 9 0 2 7 0 2 15 13 13 9 0 2 16 13 1 9 2 1 12 1 9 7 1 12 8 2
8 3 9 0 13 15 9 9 2
8 7 13 0 7 0 1 15 2
12 3 1 15 9 13 2 7 3 1 9 0 2
2 3 2
19 9 0 13 3 13 9 9 15 1 15 16 13 0 10 9 0 1 0 2
20 15 3 9 15 9 15 13 13 1 0 10 9 0 2 13 13 9 15 9 2
5 9 7 13 3 2
13 10 3 15 15 13 13 13 9 2 3 15 13 2
7 13 3 9 9 1 0 2
20 13 3 2 16 13 9 1 10 0 2 1 0 9 9 2 13 7 0 3 2
19 9 3 3 13 13 9 15 9 9 2 7 13 15 9 15 13 9 9 2
14 10 7 9 9 13 9 15 9 1 0 9 0 13 2
7 3 9 1 0 9 13 2
24 3 7 9 13 2 1 12 1 9 2 16 9 1 9 13 2 0 7 7 0 1 9 0 2
20 1 16 7 9 0 7 0 1 9 13 2 3 7 9 9 2 7 1 9 2
22 9 7 9 3 13 0 1 9 2 3 1 15 9 13 13 2 7 13 1 15 9 2
49 15 3 3 13 9 10 9 2 16 13 9 15 9 13 2 7 1 15 13 3 9 0 1 9 13 2 3 0 7 0 2 15 13 1 9 0 2 16 7 1 10 9 2 15 3 13 16 13 2
14 15 7 13 0 2 7 0 15 0 9 7 0 9 2
21 13 3 9 0 1 15 13 2 1 15 1 0 13 2 7 3 0 1 9 0 2
2 3 2
27 16 15 13 13 13 16 1 9 0 1 15 13 2 3 15 13 13 13 16 1 9 0 15 1 15 13 2
24 0 3 13 13 13 3 0 16 13 15 13 13 15 2 7 3 16 13 1 15 9 16 13 2
12 13 7 15 13 13 16 13 1 12 1 9 2
24 1 3 9 13 9 13 2 16 3 9 13 2 13 16 13 1 15 15 9 15 13 13 13 2
7 15 7 9 13 9 0 2
13 13 3 16 9 3 13 13 9 0 16 9 13 2
26 3 13 3 9 9 0 1 9 1 9 13 1 9 2 7 15 9 0 13 9 1 9 16 15 15 2
7 15 7 9 13 9 13 2
10 13 3 16 9 13 9 13 0 9 2
15 12 9 2 16 9 15 13 1 15 2 13 0 1 9 2
21 15 9 2 16 9 0 13 13 13 1 15 2 7 3 16 9 13 3 13 15 2
9 13 13 7 16 15 9 13 0 2
22 15 3 13 9 15 9 13 13 2 7 15 9 15 0 13 13 2 7 1 13 13 2
17 1 15 3 16 13 15 16 13 13 2 3 13 15 16 13 13 2
16 13 7 13 13 13 13 2 1 13 15 13 13 2 1 9 2
25 3 3 13 9 13 13 1 15 16 9 1 15 13 4 13 1 9 2 1 15 13 1 13 13 2
6 9 3 13 9 0 2
2 3 2
14 9 13 9 15 3 13 15 1 15 15 9 3 13 2
7 13 7 13 13 9 0 2
8 13 3 13 9 9 16 3 2
13 9 7 3 13 9 0 2 7 3 13 9 9 2
10 3 3 9 9 13 13 9 9 13 2
16 0 7 7 13 13 9 13 13 16 9 0 13 13 1 15 2
20 3 3 15 13 13 13 7 13 1 9 0 7 0 2 16 13 0 1 9 2
11 3 7 13 15 0 16 9 4 15 13 2
16 3 7 13 15 13 13 7 13 16 9 0 7 0 15 13 2
23 3 3 1 9 13 13 16 13 13 13 16 9 0 2 15 13 9 13 2 4 15 13 2
2 3 2
48 15 13 15 13 13 16 13 9 15 13 2 7 15 16 3 13 9 7 13 1 9 1 13 2 16 15 13 9 13 13 3 16 13 0 2 7 15 16 3 4 13 0 7 13 1 10 9 2
20 9 7 13 1 9 13 3 3 3 13 9 13 2 7 13 9 16 3 13 2
17 13 3 1 13 1 0 9 1 15 13 2 16 13 1 12 9 2
31 3 3 1 15 13 13 13 16 9 0 2 15 13 13 9 2 13 13 15 2 7 16 3 4 13 7 13 1 9 0 2
8 3 2 9 13 2 3 13 2
2 3 2
8 9 13 15 15 13 1 13 2
13 13 3 15 13 9 2 7 9 15 13 1 9 2
25 7 13 13 2 15 13 9 15 9 15 13 9 2 3 13 13 9 0 2 7 13 15 9 0 2
16 1 15 3 16 15 9 13 2 13 16 3 13 9 9 15 2
14 3 7 9 9 3 13 1 9 0 7 1 9 0 2
11 9 7 1 15 13 2 1 15 13 13 2
16 3 7 9 0 13 1 15 2 7 3 1 9 1 15 13 2
2 3 2
8 9 9 13 13 1 9 13 2
16 9 7 13 2 16 13 13 2 3 13 13 16 1 9 0 2
6 9 3 1 3 13 2
22 9 7 0 3 13 13 1 9 0 2 1 13 9 13 9 2 7 0 1 9 0 2
14 9 3 3 13 1 9 0 2 7 0 1 9 0 2
2 0 2
13 9 1 9 2 16 9 13 2 13 9 9 13 2
33 9 7 13 9 13 0 9 2 15 0 13 13 9 0 2 1 15 13 9 16 9 1 9 2 16 9 13 2 1 12 1 9 2
19 13 3 9 1 9 2 15 13 9 9 2 13 1 9 0 2 16 0 2
2 3 2
10 0 13 16 9 0 9 13 1 9 2
9 9 7 9 0 13 1 9 9 2
10 13 3 1 9 2 15 13 9 0 2
10 3 13 3 9 0 15 9 0 9 2
12 3 13 16 13 15 9 16 9 7 9 15 2
2 3 2
11 15 13 13 1 9 2 13 3 13 9 2
13 3 9 13 1 10 9 2 16 9 0 1 0 2
25 3 9 13 2 1 12 1 9 2 16 2 16 15 9 9 13 1 9 2 16 0 13 9 13 2
7 9 7 9 0 13 9 2
36 13 3 9 2 1 12 1 9 2 16 9 13 13 1 15 2 3 13 2 16 4 13 1 9 1 9 1 9 13 2 15 3 13 1 9 2
10 3 9 0 3 13 3 1 9 13 2
2 0 2
50 15 13 15 9 1 9 2 4 15 1 9 13 15 1 15 15 9 13 3 13 2 16 9 13 2 1 12 9 1 9 2 16 2 16 9 13 9 0 1 9 9 2 16 9 13 15 9 9 0 2
16 7 9 9 0 13 1 9 0 2 1 15 0 13 13 9 2
8 9 3 9 0 0 13 9 2
9 3 13 3 1 9 1 9 13 2
2 3 2
30 16 13 1 9 1 9 13 2 3 13 9 15 13 1 9 13 16 9 0 2 3 13 3 0 2 7 3 15 0 2
17 3 13 7 13 9 3 1 9 13 2 16 15 3 13 15 9 2
17 15 7 9 3 1 9 13 2 16 9 13 2 1 12 1 9 2
14 13 3 15 9 16 0 9 2 1 15 9 3 13 2
10 3 13 3 9 1 9 13 1 9 2
2 3 2
14 1 10 9 3 15 13 9 0 3 9 0 15 9 2
16 3 3 13 15 9 0 1 9 15 3 13 15 9 0 0 2
9 7 9 13 3 13 0 16 9 2
15 3 7 9 0 13 1 15 0 16 1 9 1 9 13 2
8 7 3 9 13 13 3 13 2
2 0 2
16 1 9 13 13 9 9 0 0 2 1 15 1 0 9 13 2
14 16 3 9 0 13 9 13 2 1 15 13 0 9 2
13 3 3 13 15 1 9 2 16 9 3 13 0 2
20 16 7 13 16 9 13 3 13 9 0 2 3 13 13 16 15 13 9 9 2
12 15 13 3 13 9 0 2 16 13 9 13 2
5 13 3 0 9 2
11 12 1 9 9 13 2 15 1 9 13 2
4 15 15 13 2
2 3 2
14 9 0 13 15 13 9 2 16 13 1 12 1 9 2
13 16 3 9 0 13 9 13 2 7 15 13 15 2
5 15 13 13 0 2
15 13 3 15 1 15 16 9 9 1 9 2 16 9 13 2
8 15 7 13 2 1 9 13 2
26 9 3 0 2 1 16 13 1 15 0 2 13 9 13 2 7 13 1 9 1 15 16 0 1 9 2
17 1 7 16 13 15 2 1 9 13 1 9 1 9 1 9 13 2
11 3 15 1 9 3 13 1 15 9 13 2
6 7 15 13 3 13 2
22 9 3 0 1 15 13 2 1 15 2 13 15 2 16 13 1 9 0 1 9 13 2
16 0 3 13 13 9 16 1 9 1 3 9 16 16 13 15 2
15 3 3 1 15 16 13 15 2 13 1 9 1 3 9 2
2 3 2
20 1 15 2 13 1 9 1 13 9 3 13 15 1 15 13 2 7 1 15 2
15 1 15 7 15 3 13 15 1 15 2 3 13 15 13 2
24 3 3 9 9 0 13 1 15 16 0 13 1 13 9 2 16 13 15 9 1 12 1 9 2
2 3 2
13 0 13 9 0 3 0 13 16 12 1 15 13 2
12 3 3 12 9 0 9 3 13 16 1 9 2
27 16 3 9 0 13 9 13 7 9 1 9 13 2 13 16 7 13 1 9 3 9 13 2 7 1 0 2
11 15 7 13 2 13 16 15 13 9 13 2
29 16 16 15 13 9 0 16 13 15 9 0 2 9 7 0 13 15 1 15 16 13 9 13 2 7 0 15 13 2
7 7 0 16 13 1 0 2
6 15 7 13 0 0 2
8 3 3 9 0 13 9 13 2
6 3 13 3 9 13 2
8 16 13 9 13 1 9 9 2
27 7 16 15 9 9 13 9 9 13 1 15 16 13 9 3 13 2 13 0 16 13 9 13 1 9 9 2
57 0 3 2 16 9 1 12 1 9 2 13 9 13 16 13 9 0 9 9 0 9 9 13 2 7 3 13 16 15 13 9 0 13 1 10 9 2 3 16 13 9 13 2 1 9 15 13 2 16 13 1 9 9 7 9 9 2
14 3 7 2 1 15 9 2 13 13 15 9 9 0 2
6 15 3 13 16 0 2
9 13 3 16 15 9 13 9 9 2
8 7 13 1 15 15 3 13 2
18 1 9 7 7 0 9 15 13 3 0 2 7 13 9 15 9 13 2
39 3 3 1 15 13 9 13 1 0 9 9 2 7 1 0 9 15 9 2 16 15 13 16 15 9 9 13 0 1 0 2 3 13 1 0 0 9 9 2
21 3 2 16 13 1 15 13 15 2 13 2 7 15 0 13 13 16 0 1 0 2
26 7 13 9 9 16 9 13 13 2 13 16 3 13 0 1 9 3 9 13 9 2 16 1 15 9 2
21 3 3 9 0 13 2 15 4 13 7 2 15 4 13 2 7 2 15 13 0 2
17 15 13 13 3 1 15 15 13 0 15 2 3 3 1 0 9 2
27 16 7 2 16 15 13 2 9 0 13 1 9 7 15 2 0 13 9 2 3 13 2 16 13 9 10 2
5 15 13 1 0 2
7 15 3 13 1 9 0 2
2 3 2
10 1 12 1 9 9 13 1 9 9 2
9 7 1 9 3 13 13 0 9 2
14 3 13 3 9 1 9 0 2 7 13 15 9 15 2
2 3 2
18 1 12 1 9 2 13 13 1 9 0 2 13 15 9 9 2 13 2
10 1 9 7 9 15 13 9 7 13 2
11 1 15 0 13 16 9 0 13 15 9 2
16 3 7 0 1 15 15 3 13 2 13 9 9 0 2 13 2
9 13 7 9 15 13 7 13 9 2
15 1 15 0 13 9 13 15 9 0 2 15 9 0 13 2
12 13 3 13 9 1 9 9 2 7 1 9 2
6 3 16 0 13 13 2
7 1 9 9 1 9 0 2
34 15 3 9 9 13 2 9 13 9 0 13 15 9 1 15 2 16 3 9 0 1 9 13 1 9 1 12 1 9 2 13 15 13 2
31 16 0 13 3 13 15 9 0 13 9 9 2 13 13 9 3 13 13 1 15 0 9 2 7 13 9 9 1 9 0 2
39 13 3 9 0 9 9 13 9 13 1 9 1 13 9 9 13 2 15 3 13 1 9 2 7 1 15 13 15 9 13 2 1 15 9 9 13 13 9 2
14 15 7 1 9 1 15 13 9 13 2 13 9 0 2
14 7 3 13 13 16 1 9 13 1 15 13 9 0 2
14 13 7 1 0 9 15 9 9 7 9 9 13 0 2
19 13 3 9 1 12 1 9 2 16 13 4 2 16 9 0 13 0 9 2
12 15 7 13 0 13 1 15 9 13 9 9 2
23 15 3 3 13 2 13 16 1 15 9 9 13 2 16 13 1 9 7 9 7 15 3 2
16 3 3 9 13 9 13 13 1 9 7 9 9 2 16 13 2
20 1 15 7 9 13 16 9 0 13 15 9 1 9 0 1 13 9 9 13 2
15 9 7 15 3 13 15 9 0 13 2 7 13 13 9 2
11 13 3 9 15 2 7 9 12 1 15 2
8 7 15 0 13 1 9 9 2
32 13 3 9 1 15 9 0 3 13 13 15 9 0 2 7 1 13 3 13 13 9 2 16 13 0 10 9 0 7 0 15 2
17 15 1 9 3 13 13 2 16 15 3 13 13 2 7 3 13 2
14 3 3 9 9 13 1 9 2 7 1 15 13 13 2
2 0 2
28 16 15 15 13 9 1 9 0 2 13 15 16 13 9 2 7 3 1 9 9 13 2 13 16 10 9 13 2
12 1 9 7 13 9 15 1 0 1 9 13 2
11 3 7 15 13 13 1 9 7 9 0 2
26 15 0 0 13 9 2 13 9 1 9 9 7 9 1 15 16 9 13 1 9 9 2 3 7 9 2
2 3 2
18 9 13 0 9 13 1 0 2 13 9 0 2 13 1 9 1 15 2
10 13 3 15 9 1 15 15 13 13 2
14 15 3 10 3 13 13 1 9 2 7 1 9 13 2
12 13 3 1 9 9 16 9 0 13 9 15 2
2 3 2
12 9 13 0 0 7 13 13 2 16 9 9 2
10 3 7 15 13 0 2 3 13 0 2
9 3 13 3 9 13 0 10 9 2
11 10 7 9 0 2 16 3 2 13 0 2
29 3 7 1 9 2 15 13 9 1 9 9 0 2 13 9 2 1 12 1 9 2 16 13 0 0 9 1 9 2
11 0 13 3 1 9 9 13 15 9 0 2
10 9 7 0 13 0 9 0 1 15 2
19 13 3 9 2 1 12 1 9 2 16 9 0 13 15 13 7 13 9 2
9 9 3 0 3 13 1 9 9 2
2 0 2
24 16 9 15 9 1 15 9 13 2 13 9 15 3 13 9 15 2 1 9 0 13 9 0 2
10 9 7 9 0 3 13 9 9 0 2
36 13 3 9 2 1 12 1 9 2 16 9 3 13 9 9 2 7 9 15 9 2 0 7 9 13 9 2 1 15 13 9 16 9 1 9 2
10 3 3 13 9 0 13 1 9 9 2
8 0 3 0 9 7 9 0 2
2 3 2
13 13 13 15 9 1 15 0 13 13 15 9 0 2
10 15 7 9 13 9 2 7 3 9 2
12 13 3 16 9 13 2 7 2 9 1 9 2
19 13 3 15 9 1 9 13 2 1 9 3 13 2 15 13 9 15 9 2
10 9 7 13 9 9 1 9 13 0 2
7 3 13 3 9 15 9 2
5 13 7 9 0 2
19 13 3 9 2 1 12 1 9 2 16 9 0 13 15 9 13 7 13 2
7 3 13 3 9 0 9 2
24 16 7 13 16 9 13 9 1 15 13 9 0 13 1 9 1 9 13 2 15 13 3 13 2
44 16 2 1 9 1 9 13 13 9 13 2 13 16 3 0 13 1 9 0 2 1 15 13 9 13 2 7 1 15 9 0 2 15 13 13 9 9 2 16 7 1 9 13 2
9 15 7 9 1 9 13 9 0 2
9 9 3 0 13 3 13 1 9 2
2 3 2
14 9 3 13 0 9 16 1 16 4 13 1 9 0 2
27 15 7 3 13 13 16 13 1 15 9 0 2 15 3 4 13 1 9 0 2 7 15 13 9 0 9 2
10 13 3 13 15 9 0 1 15 0 2
5 15 13 9 0 2
2 3 2
8 9 0 1 9 13 9 9 2
9 9 7 3 13 9 2 7 9 2
8 9 3 13 9 9 1 9 2
20 13 3 1 9 15 9 1 0 9 2 16 1 9 9 13 9 1 9 9 2
12 9 3 0 3 13 15 9 2 7 9 15 2
2 0 2
18 9 13 9 7 9 0 1 9 9 15 0 2 15 3 13 9 0 2
19 15 7 13 9 7 9 1 16 13 1 9 2 7 1 16 13 1 9 2
28 1 3 9 15 13 15 16 9 9 1 9 2 0 13 16 9 0 15 13 15 16 9 15 1 9 0 13 2
10 16 9 3 13 9 2 16 13 9 2
15 13 7 9 9 1 9 0 2 0 13 9 9 1 9 2
6 13 3 9 13 9 2
22 1 15 7 13 13 4 1 15 16 13 1 0 9 13 1 15 0 9 15 13 9 2
18 15 3 9 13 2 16 0 2 1 0 13 2 0 0 1 0 13 2
21 3 7 1 15 9 15 9 13 13 1 15 13 4 9 9 2 7 1 15 0 2
26 13 4 3 1 16 9 9 0 2 7 9 0 2 13 9 9 0 7 0 2 7 0 3 9 9 2
9 9 7 13 1 9 0 7 0 2
9 3 13 3 9 13 9 9 9 2
9 3 0 13 16 15 9 13 9 2
2 3 2
21 9 2 1 13 15 13 1 0 9 3 0 1 15 2 0 13 16 13 9 0 2
12 3 9 15 13 0 2 7 13 3 7 0 2
10 9 7 13 9 0 2 7 3 0 2
10 15 1 9 3 13 15 9 7 9 2
6 9 3 3 13 9 2
2 3 2
8 9 3 13 9 9 9 0 2
11 13 3 9 13 2 7 3 3 3 13 2
8 9 7 13 9 1 10 9 2
6 3 13 3 9 9 2
2 0 2
11 9 13 9 7 13 9 2 15 9 13 2
29 1 9 3 15 13 3 15 1 9 7 9 0 2 15 3 3 1 15 13 2 1 15 13 2 16 13 1 13 2
6 15 7 3 13 9 2
6 3 13 3 9 9 2
18 13 7 4 13 1 15 16 3 13 15 9 13 9 2 7 15 9 2
43 9 3 13 16 13 2 7 3 1 15 15 13 0 1 9 2 16 9 9 7 3 2 9 7 16 0 9 2 1 9 15 15 13 1 9 0 2 16 1 9 9 9 2
6 16 9 3 13 9 2
11 0 7 13 9 13 9 13 9 13 9 2
18 3 3 13 9 13 9 0 2 7 0 2 1 15 13 13 9 13 2
11 15 3 9 1 9 1 9 13 13 9 2
7 9 7 9 13 15 9 2
12 3 7 13 16 7 13 2 7 3 0 9 2
9 10 3 9 13 9 13 7 9 2
17 7 9 13 13 9 7 13 15 2 7 13 9 2 16 7 9 2
9 13 3 7 13 2 16 7 9 2
14 1 15 10 13 16 9 3 13 9 2 16 7 9 2
2 3 2
9 9 9 3 13 9 9 16 9 2
19 3 9 13 9 15 9 2 9 2 9 7 9 2 9 2 9 7 9 2
18 3 7 13 13 15 9 13 9 7 9 2 7 10 15 1 9 13 2
6 3 13 3 9 9 2
2 0 2
4 9 13 0 2
12 12 9 2 15 9 2 15 9 2 9 9 2
23 9 7 3 13 9 2 16 13 16 15 9 9 13 9 15 9 9 2 15 3 13 13 2
27 0 3 13 9 9 2 16 2 1 1 0 9 9 13 0 9 7 9 9 2 0 9 9 13 0 9 2
17 15 3 9 13 9 7 9 7 9 2 1 13 1 0 9 13 2
5 15 13 13 0 2
6 3 13 3 9 9 2
6 16 9 3 13 9 2
12 13 7 7 15 3 13 2 13 9 13 9 2
14 15 9 16 13 0 7 0 2 13 15 3 0 13 2
16 13 3 2 1 13 15 9 0 2 13 13 1 9 7 9 2
12 13 7 1 9 7 9 2 15 13 13 9 2
11 3 13 15 15 13 9 2 7 15 9 2
19 9 7 3 13 13 9 2 16 9 3 13 1 15 16 1 9 7 9 2
5 9 3 13 9 2
11 3 3 13 9 2 1 15 9 13 9 2
2 3 2
7 0 13 12 9 13 3 2
10 9 7 3 13 3 1 9 16 13 2
6 3 13 3 9 9 2
2 0 2
5 10 9 0 13 2
11 10 7 0 13 15 13 7 13 9 15 2
16 16 3 9 13 9 2 13 15 15 13 7 15 3 13 9 2
9 13 3 2 9 13 2 9 13 2
30 7 16 15 3 13 0 2 13 7 13 1 15 0 7 0 2 15 13 9 2 7 13 13 1 0 2 15 13 0 2
6 3 13 3 9 9 2
2 3 2
31 16 1 13 4 2 7 1 12 9 13 2 10 13 15 13 1 12 2 15 15 13 13 7 3 13 2 7 15 13 13 2
6 7 9 13 13 15 2
12 13 7 1 15 13 9 2 13 7 13 9 2
7 9 3 13 13 3 13 2
12 15 7 9 13 16 13 2 16 1 13 4 2
6 9 3 3 13 9 2
2 3 2
12 1 13 4 16 13 3 13 13 9 15 9 2
5 13 7 9 9 2
11 9 3 2 1 0 0 2 3 13 9 2
15 15 7 15 15 13 4 13 9 13 9 2 0 13 13 2
27 13 3 9 13 9 2 1 15 16 9 13 9 3 1 9 9 2 1 3 9 13 1 9 1 9 0 2
6 7 16 9 13 9 2
6 7 16 13 1 9 2
7 13 7 13 9 15 13 2
18 7 1 15 3 13 4 16 9 9 13 0 9 9 9 1 9 13 2
22 9 3 3 13 9 16 1 9 2 16 2 1 13 9 9 2 13 1 9 13 9 2
18 13 3 9 1 9 2 3 16 13 1 13 2 7 16 9 1 9 2
14 16 7 15 9 13 0 1 9 2 16 1 13 4 2
27 13 3 1 15 9 0 16 13 15 3 13 9 2 3 13 2 9 13 3 13 2 15 0 1 9 13 2
16 3 15 9 2 8 12 2 1 9 0 13 2 13 1 9 2
15 9 7 9 13 1 9 10 2 7 9 9 1 13 9 2
8 1 13 9 7 9 13 15 2
15 15 7 0 13 16 15 0 9 9 1 9 13 3 13 2
5 15 3 0 13 2
7 9 3 1 10 9 13 2
9 15 7 9 1 9 9 3 13 2
39 15 1 15 13 2 16 3 13 0 7 13 2 3 9 13 2 7 2 16 1 9 13 2 13 15 9 2 7 0 1 15 9 2 16 10 9 0 13 2
8 3 13 3 15 9 7 9 2
2 3 2
7 9 3 13 0 16 0 2
17 13 3 10 0 9 1 9 0 2 1 13 9 9 1 9 0 2
11 9 7 13 0 0 2 16 1 9 13 2
6 13 3 9 1 9 2
2 0 2
9 9 9 3 15 13 16 1 0 2
28 15 1 15 13 2 16 9 0 2 15 13 0 9 9 2 3 13 16 1 0 2 1 15 7 9 15 13 2
14 9 7 13 0 2 16 9 2 9 2 7 9 9 2
8 3 13 3 15 9 7 9 2
2 3 2
9 15 9 15 13 2 7 10 9 2
24 9 3 3 13 15 2 7 13 15 13 2 7 15 0 9 13 2 16 13 1 9 1 9 2
10 9 7 13 15 2 7 13 15 13 2
8 3 13 3 15 9 7 9 2
2 3 2
6 9 13 1 13 0 2
19 9 7 3 13 1 9 0 2 3 15 13 0 2 13 0 3 0 13 2
8 13 3 15 9 0 7 0 2
7 1 13 9 0 13 9 2
16 15 7 9 0 13 16 15 13 9 0 3 13 15 16 9 2
6 15 3 13 13 0 2
8 9 3 13 3 1 15 9 2
13 15 9 13 16 2 13 0 2 13 7 13 15 2
11 15 3 13 16 1 15 0 9 0 13 2
15 9 7 1 15 3 13 2 1 15 9 9 1 15 13 2
8 3 13 3 15 9 7 9 2
2 3 2
25 9 3 13 16 0 7 0 2 1 9 13 9 13 1 9 1 9 2 16 13 1 9 1 9 2
7 9 7 0 7 0 13 2
7 3 13 3 9 0 9 2
2 0 2
8 0 13 15 13 13 7 13 2
18 7 9 13 9 0 16 0 9 2 16 9 13 2 1 12 1 9 2
11 0 13 3 16 13 15 9 0 7 9 2
2 3 2
15 13 4 1 12 1 9 16 9 3 13 9 15 9 9 2
7 9 7 13 9 0 13 2
9 3 13 3 15 9 7 9 0 2
7 15 13 15 13 9 12 2
14 15 13 15 1 9 9 2 7 1 0 9 13 15 2
21 1 15 13 13 16 9 13 15 9 0 1 9 7 9 2 15 13 1 15 9 2
8 15 9 0 13 13 9 9 2
15 1 13 3 9 13 13 16 0 9 13 13 9 16 9 2
30 16 3 9 0 3 13 9 0 16 9 2 16 9 13 2 7 13 15 0 1 9 2 16 13 9 2 7 16 9 2
42 7 3 9 15 9 13 2 13 9 1 0 9 2 16 13 9 2 7 9 2 16 9 2 7 9 2 16 9 2 7 9 2 7 9 2 7 9 2 16 0 13 2
12 13 16 9 0 13 0 9 9 13 16 9 2
7 15 3 3 13 13 0 2
13 1 15 3 16 15 13 9 0 15 2 12 13 2
15 15 12 13 2 16 9 13 9 13 0 15 15 13 9 2
17 9 7 13 2 3 0 2 7 0 2 15 15 13 7 13 9 2
14 3 13 15 2 3 16 9 7 9 13 1 12 9 2
12 15 3 13 1 9 0 1 15 15 13 9 2
22 7 15 9 13 1 15 13 9 13 2 15 13 12 1 9 2 1 9 7 9 13 2
28 3 7 13 9 0 2 1 15 16 13 0 2 16 13 4 2 13 0 9 13 9 2 3 9 10 13 9 2
29 3 13 3 9 16 15 13 9 1 15 13 9 7 9 15 2 1 9 3 13 16 1 9 2 7 3 15 13 2
24 13 7 13 16 9 0 9 10 9 0 13 3 13 2 16 13 12 9 9 0 7 9 0 2
14 0 3 9 13 0 9 13 2 7 0 9 0 9 2
16 15 7 13 13 16 15 9 15 9 9 13 16 13 9 0 2
5 3 13 7 3 2
25 13 3 9 0 16 13 7 9 1 15 9 13 2 9 7 0 16 9 2 7 1 0 9 9 2
15 15 3 13 9 0 13 9 9 0 2 15 13 9 0 2
9 15 7 9 0 9 9 13 13 2
40 3 3 13 9 0 9 13 0 9 9 2 16 15 9 1 9 9 9 13 9 9 2 16 9 2 15 13 0 7 0 9 13 2 7 9 1 9 9 13 2
22 3 7 0 9 13 2 1 12 8 1 8 8 2 16 0 9 13 9 0 9 9 2
43 13 3 13 15 0 1 9 9 2 3 9 0 0 13 2 15 13 1 9 0 9 2 3 1 9 0 2 15 13 0 9 1 9 0 9 2 16 1 9 13 13 13 2
26 7 3 13 16 9 0 13 13 3 15 9 7 0 0 7 0 2 16 13 9 0 2 9 3 9 2
39 3 7 0 13 15 12 1 9 0 7 9 0 16 1 9 9 7 15 9 2 7 9 3 2 16 3 9 3 13 9 2 1 15 7 9 13 3 12 2
19 16 7 13 12 9 9 7 9 2 3 3 13 16 9 3 13 9 9 2
14 3 2 3 9 13 0 2 3 1 10 9 13 9 2
13 15 13 13 9 9 2 1 15 9 15 9 13 2
7 15 3 13 1 16 13 2
17 3 9 15 9 13 9 9 2 7 15 1 9 10 9 13 9 2
47 13 3 15 9 9 2 15 1 15 9 13 16 1 15 15 13 9 15 13 9 9 2 16 0 2 0 2 0 7 0 2 0 2 0 2 0 7 0 2 7 15 0 2 16 9 9 2
12 3 15 13 9 3 0 2 7 0 13 9 2
47 1 15 13 9 13 9 2 15 16 3 15 13 1 15 13 15 3 13 13 1 9 13 2 3 3 13 15 9 9 9 2 16 13 1 9 0 2 15 13 15 9 2 16 9 13 9 2
64 1 15 3 13 15 9 15 9 13 1 15 13 15 13 9 9 13 2 16 9 13 0 1 15 9 13 2 16 13 9 9 2 15 3 13 3 0 9 9 0 1 13 9 0 7 0 2 7 15 9 9 0 2 16 13 9 9 9 13 2 15 13 15 2
20 1 15 9 13 15 9 0 0 9 3 0 1 13 2 7 3 0 1 13 2
30 7 3 13 13 1 9 1 15 7 0 9 13 13 2 3 9 3 3 13 16 13 9 0 2 16 13 9 0 9 2
19 13 3 7 13 3 13 13 7 13 2 16 15 13 0 1 13 9 9 2
33 1 10 7 15 9 13 9 0 0 9 3 3 1 9 9 2 15 13 13 2 7 3 13 13 1 9 15 13 1 9 0 3 2
6 7 15 13 9 0 2
9 3 13 3 13 1 15 9 0 2
35 3 13 16 15 9 15 9 13 2 15 13 9 0 2 7 13 9 9 0 2 3 13 0 13 1 9 7 15 13 2 16 15 9 0 2
13 15 15 9 0 13 2 1 15 3 13 9 0 2
33 16 3 15 13 9 0 13 9 15 1 15 9 0 13 2 3 9 7 9 2 1 15 15 13 16 0 13 9 1 13 9 0 2
15 9 9 15 1 13 16 9 0 3 13 13 9 16 9 2
16 15 7 13 2 3 13 0 13 15 1 13 13 1 13 4 2
7 1 0 3 9 0 13 2
21 3 3 9 7 9 13 12 9 9 13 2 7 1 15 12 13 12 9 9 13 2
20 9 3 9 3 13 15 9 13 9 2 7 13 2 7 9 13 15 9 13 2
31 15 7 0 13 2 9 7 9 1 15 9 13 2 3 3 0 13 16 15 13 9 12 9 2 7 16 13 9 15 9 2
24 3 3 9 0 7 9 2 15 3 13 13 0 9 9 2 16 13 2 13 12 9 16 9 2
21 3 7 13 9 0 13 9 0 2 16 9 15 13 1 9 2 16 0 9 13 2
23 3 3 13 1 9 16 9 13 2 7 1 9 0 13 2 7 15 9 2 16 13 4 2
24 7 3 1 15 16 9 0 13 9 16 9 2 13 15 1 9 13 2 9 13 1 9 13 2
13 13 3 1 9 13 7 15 9 2 7 9 15 2
9 1 9 3 10 13 9 15 9 2
7 1 9 0 9 0 13 2
36 16 3 9 9 1 9 0 13 2 13 16 9 9 15 13 15 9 9 2 13 9 15 9 9 1 15 9 15 13 2 16 9 13 9 9 2
18 16 7 9 15 3 13 1 9 0 2 9 15 3 13 9 15 9 2
31 7 1 15 13 9 13 13 2 3 16 9 9 15 13 9 9 2 7 9 0 2 13 9 9 16 9 13 15 9 9 2
38 3 13 7 0 2 16 9 1 10 9 13 9 9 2 16 10 15 9 13 1 9 2 7 1 15 10 15 9 13 15 9 9 2 16 0 9 13 2
28 3 3 13 4 16 9 0 3 13 15 9 15 13 0 13 9 2 7 13 1 10 15 9 0 1 9 13 2
27 3 7 9 13 13 1 9 2 3 2 3 3 13 1 9 1 13 2 16 7 3 1 13 13 1 9 2
23 15 3 9 13 16 15 15 9 10 9 13 13 2 3 13 9 0 9 3 13 16 9 2
32 9 3 9 15 13 1 9 0 2 16 13 0 7 0 7 13 2 3 13 13 16 9 0 3 13 13 9 16 9 13 9 2
27 13 3 3 16 13 16 0 9 2 15 9 13 9 0 2 3 13 15 9 9 3 1 15 10 13 9 2
7 7 15 3 10 9 13 2
15 1 9 3 0 15 10 13 2 13 15 0 13 7 13 2
9 9 7 13 1 9 16 1 9 2
18 3 13 16 7 9 9 15 13 2 16 9 0 3 13 9 16 9 2
58 16 3 13 9 9 1 9 9 3 13 2 9 7 15 9 9 13 2 3 13 16 9 13 15 9 2 1 9 13 0 2 1 3 13 9 2 7 9 15 9 2 16 1 9 13 9 2 1 12 1 9 2 16 13 15 9 9 2
9 3 3 13 9 9 0 1 9 2
53 16 7 1 15 16 9 13 9 13 0 7 13 2 3 13 13 15 13 9 7 9 9 15 13 9 15 9 2 13 1 15 15 13 1 9 0 1 9 2 1 15 15 13 9 1 0 9 9 0 15 9 13 2
15 16 15 9 10 9 13 2 13 7 9 15 15 9 13 2
5 15 7 13 0 2
12 15 3 9 7 3 9 13 2 0 13 13 2
23 13 3 16 2 1 15 9 15 9 9 9 13 2 16 3 13 9 15 13 9 9 0 2
12 1 15 15 9 7 9 13 3 1 9 0 2
24 7 3 0 9 9 13 2 1 3 13 9 1 9 2 7 1 9 0 13 2 16 13 4 2
12 16 1 9 9 13 13 9 13 9 16 9 2
35 7 16 9 0 13 10 9 13 1 9 7 9 9 2 13 13 16 0 13 13 2 1 9 9 2 9 1 10 9 15 9 13 16 9 2
19 13 3 9 2 1 9 9 2 16 1 9 7 13 0 13 13 1 0 2
22 3 13 16 0 13 13 1 15 0 13 2 15 7 13 1 0 9 2 7 13 15 2
32 7 1 15 12 13 0 2 3 16 0 0 13 15 2 15 9 2 16 15 13 1 15 2 3 13 0 15 15 13 1 15 2
21 3 13 16 13 15 1 9 13 1 12 9 2 15 12 13 13 7 15 13 13 2
18 13 3 0 15 13 13 1 12 9 2 15 12 13 13 7 15 13 2
6 10 7 3 13 13 2
14 0 3 0 2 3 9 2 13 13 2 1 9 9 2
32 3 7 1 12 1 9 13 13 16 9 13 13 2 7 1 15 13 1 15 13 9 9 3 0 1 15 2 7 3 1 15 2
13 13 3 2 1 9 9 2 15 9 13 9 13 2
24 13 7 1 12 0 2 16 1 9 9 13 13 15 15 13 3 0 2 7 15 15 13 13 2
19 15 7 15 13 3 0 2 13 16 0 2 7 0 16 1 15 15 13 2
20 13 7 16 3 16 0 9 9 2 15 13 9 9 2 7 16 0 0 9 2
12 3 13 16 0 13 3 13 13 0 7 0 2
23 3 15 15 1 15 13 2 3 9 2 13 13 7 13 0 9 16 15 2 16 13 13 2
15 13 3 9 13 2 1 9 9 2 1 9 0 7 9 2
33 7 15 13 1 12 1 9 2 16 13 16 15 13 0 7 9 2 16 9 2 7 16 15 3 13 15 2 7 0 2 3 9 2
13 13 7 16 9 3 13 9 0 2 1 9 9 2
11 13 3 0 9 2 15 3 13 9 9 2
39 7 1 15 13 2 13 9 16 15 1 9 0 13 9 2 13 10 15 9 2 16 13 13 16 15 0 13 9 15 3 13 15 9 9 2 3 9 0 2
26 3 13 3 13 16 9 13 9 0 1 9 2 7 13 13 16 9 1 10 9 13 9 0 16 9 2
42 3 3 7 9 0 2 15 13 1 10 9 9 0 2 7 9 10 9 9 2 1 10 9 13 2 0 2 1 9 9 9 0 13 3 1 15 9 7 16 9 15 2
27 15 7 15 13 4 1 9 9 2 3 13 3 13 1 9 9 2 1 15 15 13 7 3 7 15 13 2
9 3 9 2 1 9 9 2 13 2
36 7 15 3 0 13 2 3 1 15 9 2 3 9 2 13 9 7 9 7 10 9 2 16 15 0 13 9 2 3 1 9 7 9 2 13 2
6 16 9 0 13 9 2
45 1 13 7 13 13 8 9 0 9 13 2 7 13 13 15 0 3 9 9 13 2 7 9 2 16 13 9 2 7 9 15 2 16 15 13 2 7 3 9 0 2 16 15 13 2
11 13 4 3 16 9 13 9 16 9 15 2
8 9 7 13 9 1 10 0 2
17 1 15 3 13 9 16 13 9 15 9 2 7 3 1 15 15 2
27 3 7 13 15 12 13 1 9 7 9 16 9 2 15 9 13 1 9 2 16 13 9 2 1 12 0 2
11 3 9 7 9 13 15 16 9 7 9 2
24 13 3 13 15 13 0 1 9 7 9 2 16 3 1 13 2 3 1 13 7 1 9 9 2
19 1 13 3 2 16 1 9 15 9 13 9 2 13 15 9 0 7 9 2
10 9 3 10 9 10 13 1 10 9 2
20 3 13 9 13 9 2 7 3 9 13 9 2 7 0 12 9 13 15 9 2
18 1 9 7 9 9 1 9 13 9 1 9 2 16 13 0 1 13 2
21 3 7 9 9 15 13 0 0 15 9 2 15 9 13 13 0 1 9 7 9 2
12 16 9 13 15 1 15 7 15 1 15 9 2
18 1 15 7 13 13 9 15 1 15 9 13 2 7 15 1 0 9 2
9 13 3 0 9 1 0 0 13 2
12 9 7 13 9 9 0 2 3 12 9 3 2
23 13 3 1 15 9 2 7 3 1 12 9 3 2 1 10 9 2 1 15 13 9 9 2
14 3 7 9 13 9 15 9 16 3 13 9 0 9 2
33 16 3 13 9 15 7 3 9 2 3 13 9 0 15 9 2 16 9 9 2 15 13 9 15 7 3 0 9 2 13 9 0 2
22 16 7 13 9 0 15 7 9 2 13 1 15 16 1 15 13 9 7 15 7 9 2
13 3 2 15 13 2 7 15 7 9 13 15 9 2
11 3 9 13 7 9 15 3 13 16 0 2
28 16 3 9 13 9 0 9 2 9 7 13 1 15 15 13 9 2 13 16 13 1 10 9 1 15 9 9 2
7 16 7 15 2 0 13 2
18 1 3 15 13 1 9 1 9 2 13 15 9 13 16 9 13 9 2
5 13 7 9 0 2
16 12 3 9 2 16 13 15 1 9 2 16 0 13 9 0 2
18 15 9 2 16 13 15 1 9 9 2 16 9 7 9 13 9 9 2
12 13 3 15 7 1 9 2 7 1 9 9 2
22 15 7 7 9 1 9 13 9 3 13 16 1 9 2 3 16 13 9 9 9 13 2
13 15 7 7 9 1 9 9 13 1 9 1 15 2
28 1 15 3 9 13 2 15 1 15 9 13 2 1 15 9 13 16 13 15 1 15 7 15 1 15 9 15 2
20 3 9 2 16 1 15 9 9 13 1 15 9 2 3 7 1 15 9 15 2
11 1 7 13 1 9 15 1 9 13 9 2
13 3 3 3 13 13 16 15 9 13 1 15 9 2
42 16 3 13 15 9 15 3 13 9 9 2 16 13 9 9 9 2 3 13 9 9 2 1 15 3 13 16 12 9 2 7 0 13 13 15 15 13 1 15 9 9 2
32 7 13 15 0 13 15 15 13 9 3 3 13 0 16 9 2 7 3 0 0 13 16 9 1 3 13 2 16 1 13 4 2
18 3 13 7 9 9 2 1 13 15 9 0 2 13 9 9 3 0 2
9 16 15 9 13 9 1 10 9 2
14 3 7 15 9 13 0 7 0 2 3 13 0 9 2
23 3 9 2 15 13 0 1 9 9 2 16 0 1 9 2 13 0 1 9 7 0 9 2
30 3 13 0 9 1 10 9 13 2 15 0 9 9 0 9 13 13 2 16 9 9 2 9 9 2 7 3 1 15 2
14 1 15 9 9 13 0 9 1 9 2 9 0 0 2
41 15 3 9 1 15 9 13 4 9 13 1 15 9 9 2 16 1 15 9 2 1 9 1 9 9 9 2 13 13 1 9 2 16 15 9 15 15 9 9 13 2
30 9 3 9 2 1 15 9 1 9 15 13 2 13 0 1 9 2 1 15 9 1 15 9 9 7 15 3 9 13 2
10 16 9 0 3 13 12 1 10 9 2
31 1 13 7 0 13 3 13 12 9 0 10 9 15 13 7 15 13 7 15 13 2 16 9 2 1 12 1 9 2 13 2
12 13 4 3 16 9 9 13 9 0 16 9 2
18 0 13 7 12 9 13 16 12 9 2 16 0 9 1 0 9 13 2
6 13 3 1 3 13 2
8 3 13 3 9 12 10 9 2
2 3 2
6 15 9 13 0 9 2
9 15 3 13 9 9 2 15 9 2
17 9 7 13 1 9 16 9 15 2 16 9 13 1 12 1 9 2
21 16 3 0 13 16 9 13 9 9 2 3 0 13 16 9 12 9 13 9 15 2
2 3 2
37 9 2 1 12 1 9 2 13 0 1 15 16 2 13 1 9 2 15 1 0 0 13 2 16 13 13 2 1 0 9 2 15 9 15 9 13 2
19 3 13 3 0 16 9 9 13 9 9 2 7 9 9 15 9 16 9 2
21 7 15 13 9 9 9 1 9 9 2 15 13 9 9 15 9 1 9 15 9 2
14 3 13 3 0 9 15 9 13 15 9 16 15 9 2
11 7 9 15 9 13 1 15 15 9 13 2
13 9 3 1 9 13 1 9 9 1 12 1 9 2
10 3 13 3 12 9 15 7 15 9 2
2 0 2
8 1 15 15 13 9 7 9 2
7 12 3 7 9 15 13 2
8 7 15 13 9 1 10 9 2
8 3 7 9 9 13 9 9 2
9 0 13 3 0 9 13 9 12 2
8 9 7 15 9 13 9 0 2
9 0 13 3 10 9 13 12 9 2
33 16 7 13 16 9 0 15 9 13 15 1 9 0 15 2 7 1 3 3 13 12 9 2 16 13 12 9 2 15 13 3 13 2
11 0 3 9 15 9 13 7 13 9 15 2
23 16 7 9 0 9 13 13 2 3 9 0 9 13 13 2 16 9 13 2 1 12 9 2
28 3 13 16 2 16 15 9 13 9 1 9 2 1 9 2 1 12 1 9 2 3 13 9 1 15 15 13 2
22 15 7 15 13 9 2 7 9 1 9 2 13 9 0 2 16 13 1 12 1 9 2
9 13 3 15 9 9 1 9 0 2
34 16 3 15 9 13 15 9 0 1 15 9 2 3 7 15 9 0 2 7 12 7 15 2 13 16 13 12 9 2 7 3 12 9 2
5 15 13 0 13 2
9 3 13 3 12 9 0 10 9 2
42 15 7 9 13 9 13 2 1 12 1 9 2 13 16 9 0 13 15 1 9 10 2 3 1 9 0 2 15 12 9 13 9 1 15 13 2 15 13 1 0 0 2
18 7 3 9 0 13 1 0 2 3 9 10 9 2 7 9 10 9 2
15 16 7 15 9 15 13 2 13 1 15 15 1 13 4 2
18 13 4 3 1 16 3 13 0 9 13 16 3 0 9 0 13 15 2
22 13 7 16 13 9 13 1 15 16 9 13 13 2 3 9 13 9 1 13 3 13 2
18 1 3 13 9 2 15 1 9 13 13 13 1 9 9 16 0 9 2
31 7 15 15 9 3 4 13 1 16 4 13 1 9 2 16 3 13 1 9 0 2 7 4 13 1 0 9 1 9 13 2
16 9 7 2 1 16 4 13 1 9 2 3 13 9 9 0 2
14 3 3 3 13 15 15 9 1 15 16 1 9 0 2
14 7 13 13 9 2 16 3 13 0 9 15 7 15 2
2 3 2
17 15 13 9 1 15 15 13 1 9 2 7 1 15 15 13 9 2
16 9 7 2 1 16 4 13 2 13 3 1 9 1 9 0 2
21 3 1 9 2 1 16 13 2 3 13 15 9 9 9 0 2 15 13 9 9 2
15 7 3 13 15 15 9 0 13 2 3 4 13 1 0 2
2 3 2
27 15 1 15 9 13 15 13 2 13 9 0 2 7 3 9 0 2 16 13 1 9 2 1 12 1 9 2
11 9 7 3 13 9 0 2 7 9 0 2
17 13 3 9 9 13 1 9 1 9 2 16 13 1 9 1 9 2
14 3 13 3 15 9 15 13 2 1 15 9 9 13 2
2 0 2
10 9 15 4 13 1 9 2 0 13 2
11 15 7 15 15 9 13 2 13 13 12 2
6 3 9 12 13 12 2
21 3 3 1 9 2 16 13 13 1 0 2 16 4 13 1 9 2 9 9 13 2
2 3 2
33 15 15 9 13 9 2 13 3 13 13 1 15 9 16 13 2 15 9 3 3 13 12 7 15 9 2 7 3 15 2 3 15 2
21 9 7 3 3 15 13 1 12 9 2 7 15 1 0 13 2 7 15 13 13 2
22 9 3 9 7 1 9 13 9 2 7 1 15 13 9 10 9 2 15 13 9 0 2
49 16 7 13 16 15 9 3 13 9 1 15 9 2 7 1 9 1 15 13 9 2 3 0 2 0 7 0 2 15 13 0 9 2 15 9 1 12 1 9 2 0 9 13 2 3 13 15 9 2
31 16 2 1 9 0 13 9 0 1 0 2 15 9 13 7 13 2 7 13 9 0 1 15 13 2 3 13 9 9 0 2
16 9 7 1 9 0 3 13 16 13 9 2 7 16 13 9 2
16 3 3 13 16 13 1 15 0 15 15 13 9 16 13 9 2
2 3 2
22 9 0 2 1 13 1 9 2 3 13 15 15 13 2 1 13 3 13 9 15 9 2
22 15 7 15 13 2 13 15 15 9 13 9 2 1 13 13 0 9 9 13 15 9 2
28 3 13 3 15 9 9 1 9 0 2 7 15 9 13 15 1 15 9 0 13 1 0 2 16 9 13 13 2
2 3 2
32 9 0 3 13 9 1 9 0 2 15 13 9 2 16 1 10 9 15 13 9 16 1 9 13 13 0 9 7 13 9 0 2
10 9 7 15 3 3 15 13 1 15 2
19 0 13 3 16 9 1 15 7 13 9 9 0 2 7 1 15 13 9 2
10 3 3 13 16 13 9 3 13 13 2
2 3 2
28 15 15 15 13 7 13 2 13 9 1 15 13 9 3 0 3 1 9 15 2 7 3 3 1 9 7 9 2
34 1 15 3 9 3 13 16 12 13 2 7 12 9 0 2 16 13 13 0 13 2 7 0 9 0 2 1 9 13 3 1 12 9 2
16 9 7 0 13 15 13 9 2 16 13 9 1 12 1 9 2
24 16 3 9 0 15 7 15 9 13 12 7 15 9 2 0 13 3 13 15 13 12 7 15 2
5 15 13 13 0 2
9 3 0 9 0 13 13 9 12 2
11 0 13 3 9 0 13 12 15 7 15 2
16 16 7 13 16 15 13 13 1 9 9 2 15 13 3 13 2
20 16 3 13 4 2 12 9 12 9 13 0 1 0 9 1 15 13 15 9 2
34 13 7 7 13 2 7 3 2 3 13 9 13 1 0 9 2 7 13 1 15 9 3 9 15 9 2 16 13 1 9 1 12 0 2
12 3 13 3 12 13 9 0 13 1 9 9 2
2 3 2
28 9 15 13 1 9 0 16 0 3 1 0 2 1 16 9 13 2 1 12 1 9 2 16 13 15 13 13 2
19 13 7 15 0 13 1 0 9 0 7 9 2 3 1 9 15 1 9 2
42 1 12 3 0 13 3 1 12 0 2 3 13 7 13 2 13 7 13 2 3 7 1 12 13 13 1 12 0 0 13 2 7 12 3 2 16 9 13 0 9 9 2
38 1 3 9 0 12 9 3 13 13 1 12 9 2 9 7 13 1 9 1 15 2 16 13 12 9 7 15 9 2 3 13 13 0 13 1 12 9 2
21 7 15 13 2 16 13 15 9 9 2 16 13 1 9 9 9 2 9 7 9 2
30 1 9 3 9 9 0 3 13 16 1 0 9 9 2 16 13 16 15 13 15 13 16 13 9 2 7 16 13 9 2
9 7 15 12 13 3 13 10 9 2
13 3 3 13 16 15 13 9 13 15 9 7 15 2
2 3 2
22 9 0 13 9 2 3 1 16 13 15 9 2 7 16 13 9 0 2 1 9 9 2
29 15 7 9 12 13 2 15 9 9 13 2 7 1 12 9 7 1 0 2 1 0 9 9 2 15 0 13 9 2
17 9 3 9 3 13 13 9 16 13 15 13 9 0 9 12 9 2
10 7 3 3 13 12 9 9 0 9 2
2 3 2
16 0 9 9 9 13 9 0 2 16 15 9 13 13 1 9 2
13 9 7 2 16 13 12 2 3 13 16 1 9 2
29 16 3 9 0 13 12 10 9 2 0 13 16 9 9 15 1 9 2 13 9 9 2 13 15 9 1 10 9 2
4 15 13 0 2
9 3 13 3 9 0 12 1 10 2
20 7 1 15 13 16 9 9 9 3 13 9 0 2 7 9 0 7 9 0 2
6 15 3 13 3 13 2
23 3 2 16 13 9 2 1 12 9 2 1 0 9 13 0 9 2 7 0 3 9 13 2
21 1 9 7 9 0 13 9 9 1 15 2 7 1 15 9 13 13 1 9 9 2
11 9 3 9 13 1 9 0 2 3 0 2
2 3 2
6 9 13 1 9 9 2
14 3 9 13 9 13 13 2 16 9 13 1 12 0 2
10 9 7 9 13 0 2 16 7 9 2
10 13 3 1 15 9 15 13 0 0 2
12 9 7 0 3 13 0 0 2 7 0 9 2
7 3 13 3 9 9 9 2
2 3 2
17 1 15 13 0 9 13 1 2 1 1 13 9 0 1 9 13 2
33 13 7 1 15 13 9 1 13 9 9 1 9 0 13 2 16 9 13 13 7 0 13 1 9 9 1 0 9 9 0 7 0 2
43 7 15 9 13 1 15 9 16 1 9 13 2 16 3 13 1 9 9 7 9 9 2 1 16 13 9 2 1 12 1 9 2 9 0 9 7 0 9 13 3 0 9 2
13 1 9 7 9 13 9 13 16 1 0 9 9 2
25 13 3 16 9 9 13 9 15 13 2 16 13 1 13 0 2 16 7 15 9 9 1 15 13 2
2 3 2
28 9 13 9 13 1 9 9 2 3 9 2 15 1 9 15 9 13 1 15 16 0 13 0 9 1 9 13 2
19 9 7 15 13 1 9 9 2 3 13 9 2 7 15 13 1 9 9 2
26 3 3 9 15 0 13 13 2 13 9 9 2 7 9 15 9 9 2 3 0 2 13 1 0 13 2
23 3 0 13 16 9 9 3 13 1 9 0 2 16 9 13 13 2 7 3 1 9 0 2
2 3 2
39 16 12 13 9 0 10 9 2 13 13 9 0 3 13 2 16 9 3 13 2 16 13 2 7 0 3 9 13 2 16 9 13 0 0 2 16 9 13 2
15 7 16 9 13 0 2 7 13 0 2 13 13 13 0 2
10 3 9 0 1 0 13 1 9 0 2
9 3 3 1 0 13 15 9 0 2
18 1 15 7 9 7 9 13 0 1 13 16 16 1 15 13 9 0 2
11 9 3 3 13 0 1 13 2 7 9 2
21 7 13 9 9 2 16 9 3 13 1 9 2 7 1 15 13 1 13 0 13 2
51 7 1 15 13 9 13 2 16 9 0 13 0 9 2 1 12 15 13 9 2 3 1 9 0 2 1 15 7 13 9 2 3 1 9 2 16 3 9 0 9 13 0 2 3 9 1 9 7 9 0 2
7 15 7 9 13 3 13 2
13 0 3 13 16 9 7 9 0 13 1 15 0 2
14 9 7 0 13 2 1 0 3 1 15 13 1 9 2
30 0 13 3 8 9 0 2 15 9 0 13 9 7 13 2 13 1 9 2 16 9 0 13 1 9 15 13 1 9 2
2 0 2
17 15 13 15 3 13 2 16 13 13 4 13 1 13 2 1 9 2
13 7 9 0 1 10 13 7 10 13 1 9 0 2
19 3 3 15 13 1 15 13 2 16 9 0 4 13 1 9 1 9 0 2
37 7 13 13 8 9 15 0 13 1 9 0 2 13 13 2 16 9 0 3 0 13 2 7 13 15 13 2 3 1 12 1 9 13 13 9 9 2
11 3 1 9 10 3 13 9 1 9 0 2
11 3 3 1 9 13 13 0 9 10 9 2
2 3 2
8 13 13 1 13 1 9 13 2
8 7 9 1 15 13 1 9 2
11 3 15 13 1 15 2 13 13 7 0 2
2 3 2
35 1 9 13 0 9 16 9 2 13 16 13 3 13 2 7 1 15 13 16 12 9 13 9 1 0 9 0 2 15 1 0 9 0 13 2
16 3 13 13 16 9 13 1 0 9 0 2 1 12 9 13 2
19 9 7 0 15 13 3 2 16 9 2 15 7 13 2 16 9 7 9 2
5 3 7 9 13 2
12 13 3 16 9 0 7 13 2 7 13 13 2
2 0 2
31 1 9 0 0 13 13 16 15 1 15 13 1 9 2 3 13 2 7 3 13 13 2 1 16 13 9 13 10 3 13 2
7 13 3 9 1 9 13 2
13 0 3 0 13 13 16 13 1 9 0 3 13 2
2 3 2
37 16 1 9 15 13 1 15 9 0 3 13 15 9 0 2 16 3 13 1 9 15 15 13 1 15 2 0 9 2 1 15 9 13 15 15 13 2
14 7 15 15 15 13 2 16 9 13 0 2 16 13 2
10 3 3 9 0 13 15 9 1 9 2
15 3 3 13 9 13 1 9 2 16 13 9 13 0 9 2
2 3 2
13 1 15 13 13 16 9 0 3 13 9 1 13 2
7 15 7 1 9 0 13 2
10 7 3 15 9 7 9 13 1 13 2
9 15 13 0 0 7 1 9 9 2
52 16 7 13 16 2 0 9 2 3 13 9 1 13 15 15 9 0 13 1 9 13 2 3 16 9 0 13 0 1 0 2 15 13 1 9 2 15 13 16 3 1 9 13 9 2 13 16 3 13 13 9 2
15 9 3 0 2 16 7 15 9 2 13 1 9 10 9 2
8 1 7 10 9 13 9 9 2
12 3 13 3 0 2 7 13 15 1 15 0 2
18 15 9 13 2 16 1 9 0 9 0 13 2 1 15 15 13 13 2
24 15 3 9 15 13 9 0 1 9 15 13 2 1 9 0 2 7 15 9 16 13 9 0 2
12 1 3 2 13 15 16 1 15 13 9 0 2
10 3 15 13 1 9 0 16 9 13 2
16 7 1 9 1 15 13 2 13 15 3 9 7 9 10 9 2
9 3 15 13 1 9 16 9 13 2
26 1 3 9 9 13 1 9 9 13 15 9 0 2 1 15 13 9 0 16 0 1 13 7 1 9 2
18 16 3 9 0 3 13 9 2 3 13 1 9 16 13 1 9 9 2
2 3 2
12 9 0 13 15 9 7 9 13 2 1 9 2
30 16 7 9 0 13 12 10 7 0 2 13 16 1 15 3 4 13 10 9 0 15 15 1 15 9 4 13 7 4 2
29 15 3 10 2 15 1 9 0 13 2 3 15 13 13 15 13 9 0 2 13 10 15 4 7 4 1 15 13 2
5 15 13 13 0 2
24 1 15 7 9 13 13 2 13 16 15 3 13 1 9 0 16 1 16 13 15 1 10 9 2
21 7 16 3 13 15 9 1 10 7 15 9 13 2 7 15 13 12 2 13 15 2
7 7 13 15 9 13 13 2
25 3 3 16 9 0 3 13 12 2 3 13 15 15 9 13 1 9 0 16 13 9 1 15 13 2
13 7 16 13 9 3 13 0 9 13 2 3 13 2
25 1 9 0 13 4 9 1 9 0 13 2 13 13 1 15 2 16 13 9 2 1 12 1 9 2
18 3 13 16 15 15 9 3 13 2 13 1 9 10 3 13 1 13 2
44 7 13 1 9 2 16 1 9 10 13 13 9 0 9 15 13 2 16 9 13 9 1 9 9 15 13 2 16 13 1 0 7 0 2 15 3 13 13 0 9 9 7 0 2
48 7 1 15 9 13 2 1 12 8 2 16 15 15 3 13 9 9 2 16 13 9 13 2 3 13 9 15 13 15 1 9 1 9 2 16 13 13 2 7 13 15 13 1 9 9 16 13 2
46 16 7 1 9 0 13 9 0 10 9 2 15 13 13 16 13 12 7 0 2 9 9 1 9 0 13 16 13 15 15 3 13 9 1 13 1 9 15 2 15 3 1 9 3 13 2
30 1 3 15 9 13 1 9 0 1 16 4 13 1 9 1 9 0 2 15 9 13 13 2 1 13 2 13 10 9 2
5 15 13 0 0 2
9 3 3 15 13 9 1 13 9 2
9 3 13 3 12 7 0 9 0 2
14 1 9 9 2 15 13 9 0 3 13 1 9 0 2
9 13 0 9 13 13 15 9 13 2
22 13 3 2 1 10 9 1 9 2 16 1 9 0 3 13 9 0 16 16 9 13 2
20 15 3 1 15 13 13 2 16 2 16 9 13 13 1 9 0 2 9 13 2
26 1 15 3 13 9 1 9 2 16 13 15 1 0 1 9 2 7 0 9 1 9 13 13 1 9 2
32 3 13 16 2 16 9 7 9 4 13 12 1 0 7 13 2 1 16 13 9 15 2 13 9 1 9 1 9 7 1 9 2
54 9 7 15 13 9 3 13 1 9 2 13 3 13 9 0 2 7 9 9 0 2 16 9 2 15 13 9 9 13 1 9 2 7 9 2 15 13 2 1 15 2 9 9 13 1 9 2 16 1 9 13 9 9 2
26 15 7 13 3 9 16 13 9 3 13 9 2 16 13 15 9 0 2 1 15 13 9 9 0 9 2
17 7 1 15 2 9 0 2 13 15 1 3 9 2 13 1 9 2
16 13 7 16 9 0 13 9 0 2 7 16 3 13 9 0 2
18 3 13 16 0 13 16 9 0 13 1 9 0 2 16 16 13 9 2
66 13 3 16 7 15 9 0 13 1 15 9 0 2 7 1 15 9 13 9 0 2 7 13 16 9 0 13 1 15 13 2 1 15 13 9 0 10 16 9 1 9 15 13 1 9 2 7 13 16 9 0 13 1 9 0 1 0 1 15 9 13 2 16 9 13 2
22 0 7 15 12 13 0 2 16 9 13 1 9 13 9 0 2 13 0 1 9 3 2
13 0 7 13 9 9 2 15 13 9 2 1 0 2
27 3 13 0 2 16 16 13 9 2 13 9 0 1 9 0 10 1 9 13 2 15 13 15 15 9 13 2
49 16 0 15 13 1 15 16 3 3 13 9 1 9 1 0 13 2 7 1 3 13 13 1 9 15 0 13 2 13 16 13 15 15 13 16 13 9 9 13 15 9 9 1 13 1 15 9 0 2
13 7 3 1 13 13 0 9 1 9 1 15 9 2
7 13 0 13 16 9 13 2
27 13 3 15 9 13 16 9 2 1 9 1 9 2 13 9 3 13 1 9 0 2 7 1 9 9 0 2
13 1 15 13 16 9 9 0 3 13 1 9 0 2
20 7 16 13 13 2 15 9 2 3 1 9 2 9 7 15 13 1 9 9 2
18 13 3 9 9 0 13 15 9 13 2 1 15 9 13 1 9 10 2
21 15 7 13 1 12 9 13 2 15 13 9 13 1 15 2 9 1 9 10 13 2
21 3 7 13 2 3 1 9 13 9 2 3 1 12 7 0 9 13 9 10 13 2
11 3 3 13 16 9 10 3 13 1 0 2
20 15 0 13 1 15 16 15 13 15 9 2 13 9 0 15 13 1 9 15 2
48 13 7 16 1 15 16 9 0 13 0 15 13 1 9 2 13 9 9 13 1 13 0 2 7 16 9 9 9 2 3 9 7 0 7 0 2 13 13 9 1 13 9 9 13 2 13 0 2
22 13 3 16 9 10 3 3 13 1 13 1 9 13 2 3 3 1 0 7 0 13 2
16 1 9 3 1 15 15 1 13 2 13 1 15 15 1 13 2
22 3 3 13 0 16 1 15 16 9 13 1 9 0 2 16 13 1 13 9 9 13 2
9 9 7 9 10 9 0 4 13 2
28 13 3 16 0 3 13 13 9 1 13 9 9 13 2 7 0 13 9 1 13 15 15 9 13 1 0 13 2
16 13 3 16 1 9 1 9 13 13 9 1 9 10 10 0 2
7 3 13 13 13 15 13 2
8 7 15 0 13 1 15 9 2
29 3 2 1 9 13 13 0 7 3 15 9 15 13 2 3 1 15 13 9 9 1 9 10 2 15 13 15 0 2
2 0 2
12 15 13 1 15 2 13 1 15 1 9 13 2
12 9 7 9 0 13 3 0 16 9 9 0 2
25 1 3 9 13 1 9 0 1 9 13 2 1 15 2 13 1 15 2 0 3 13 1 9 0 2
2 3 2
6 9 0 13 9 0 2
18 16 3 1 0 9 13 15 13 13 2 0 0 15 13 1 9 0 2
2 3 2
29 13 16 0 15 1 9 9 9 13 1 0 9 2 1 0 9 13 1 12 2 16 9 0 13 0 10 9 0 2
27 13 3 7 13 2 15 1 9 9 0 13 1 0 9 2 13 16 1 0 9 2 3 1 9 2 13 2
2 3 2
10 9 13 2 1 15 2 13 10 9 2
25 16 3 13 15 13 15 16 13 16 13 9 13 2 15 13 12 9 2 3 3 13 15 16 15 2
5 15 13 13 0 2
25 13 3 16 15 9 13 1 9 9 2 15 13 2 1 12 1 9 2 16 9 0 13 9 9 2
17 15 15 15 13 13 16 15 13 9 0 9 2 16 9 9 13 2
2 3 2
20 3 13 16 16 9 0 13 9 2 13 13 13 1 15 2 16 3 9 13 2
8 3 3 13 9 15 0 9 2
40 13 3 2 1 12 9 2 16 1 13 13 9 1 9 0 1 9 2 7 3 13 9 1 15 13 1 9 2 3 7 2 16 3 13 2 13 1 15 9 2
7 3 3 13 9 9 13 2
20 13 3 2 1 12 1 9 2 16 9 15 13 1 9 0 16 0 1 9 2
17 3 13 16 9 0 13 1 9 0 1 9 2 3 1 9 13 2
13 9 7 15 13 1 0 13 2 3 13 0 13 2
14 9 3 0 13 1 9 9 1 9 0 1 13 9 2
25 1 0 3 13 9 2 3 13 1 9 9 1 15 9 2 7 15 13 0 9 1 9 7 9 2
30 7 15 13 16 9 13 2 1 12 1 9 2 16 2 1 15 9 2 3 9 0 2 15 13 2 13 13 1 9 2
9 15 7 13 1 13 13 1 15 2
17 13 3 7 3 9 0 3 2 3 3 0 7 1 13 7 13 2
16 9 0 1 9 0 13 2 16 13 15 16 13 1 13 9 2
6 3 13 3 16 13 2
20 7 3 2 1 3 13 1 0 9 2 3 13 1 9 0 2 15 13 0 2
19 7 1 15 3 13 16 9 0 13 0 0 2 15 13 1 10 9 0 2
9 9 9 15 13 13 9 9 0 2
17 1 13 7 9 9 0 15 9 13 2 15 13 13 0 3 13 2
19 13 3 16 10 9 15 13 12 1 9 7 13 1 9 2 13 1 9 2
18 15 3 13 12 9 7 0 1 9 2 13 1 9 7 13 1 9 2
30 16 3 9 0 1 0 9 4 13 1 9 2 1 13 12 1 9 2 13 16 4 13 1 15 7 1 15 1 9 2
25 3 7 1 9 15 13 9 15 2 16 3 13 9 15 1 9 9 9 0 2 7 13 9 0 2
6 15 13 1 9 9 2
14 13 3 16 13 1 9 15 13 9 9 15 13 9 2
14 10 7 9 13 1 9 15 13 9 2 13 9 0 2
15 13 3 16 9 15 9 13 1 15 1 15 13 9 15 2
18 16 3 9 0 13 1 9 9 2 3 9 13 13 1 9 15 9 2
9 13 3 16 9 0 13 9 0 2
13 7 1 13 16 3 13 15 7 13 1 9 0 2
8 15 3 13 1 9 9 0 2
14 3 9 0 3 13 1 0 9 2 7 13 12 10 2
2 3 2
30 16 9 0 13 15 1 15 7 1 15 9 2 13 16 9 13 13 15 9 1 15 7 1 15 2 12 0 1 9 2
27 1 3 9 13 1 9 0 9 13 9 0 2 13 16 2 13 9 0 2 13 9 0 1 9 1 0 2
18 9 7 7 9 15 13 15 1 9 7 0 1 9 2 13 9 0 2
15 15 3 13 13 9 0 2 16 0 13 0 2 3 0 2
12 0 13 3 9 0 4 13 1 0 9 9 2
9 0 13 3 16 13 12 1 10 2
2 3 2
8 9 9 15 13 13 1 9 2
13 7 3 15 9 2 7 15 9 0 2 3 9 2
25 0 13 0 13 2 16 3 9 13 9 10 1 9 16 13 9 10 1 15 13 15 0 1 9 2
7 15 13 13 1 9 0 2
10 13 3 16 15 9 9 13 1 9 2
11 15 13 3 13 16 13 12 9 0 15 2
10 0 3 13 9 0 13 12 10 9 2
22 16 7 13 9 9 3 13 2 16 13 4 2 3 9 13 1 15 13 0 0 13 2
43 13 3 9 0 13 12 9 1 0 9 2 0 7 1 9 2 16 3 3 13 1 15 9 2 16 9 9 3 13 1 9 7 9 1 15 2 7 0 16 13 9 15 2
13 7 3 13 16 13 9 0 1 13 13 1 9 2
33 16 3 9 0 1 10 9 13 16 15 9 1 9 13 2 3 15 9 13 1 15 9 0 1 15 16 1 15 9 9 9 13 2
27 7 3 13 9 0 2 7 1 13 9 0 2 15 13 9 9 2 1 9 2 3 3 9 1 9 13 2
21 0 0 9 15 13 2 1 15 16 3 13 1 15 15 13 2 7 15 15 13 2
13 9 3 13 1 9 0 3 13 15 16 15 13 2
24 1 3 1 15 15 13 13 10 9 7 9 2 13 16 10 9 13 1 9 13 1 9 0 2
5 15 13 13 0 2
12 15 3 9 1 15 15 13 16 0 7 0 2
11 7 3 1 15 15 13 1 10 9 13 2
39 13 15 3 9 0 13 1 9 0 1 13 16 15 15 13 2 3 16 15 15 13 2 16 7 9 9 1 9 3 13 15 15 13 2 7 15 15 13 2
23 15 0 15 13 2 13 15 9 9 13 1 9 2 16 7 9 1 9 13 9 0 13 2
16 1 15 3 13 4 9 7 9 16 9 1 10 9 13 13 2
24 7 3 13 16 2 16 9 13 1 0 2 16 0 13 1 9 1 15 13 2 16 9 13 2
23 16 16 1 9 9 0 13 16 9 9 13 2 3 3 13 16 15 13 9 9 7 9 2
11 15 3 13 13 1 9 2 3 13 13 2
10 3 3 12 9 13 7 0 7 0 2
11 9 3 13 0 9 2 7 9 0 9 2
23 3 3 7 9 13 9 1 9 0 13 2 1 9 0 2 16 7 1 9 0 13 13 2
12 15 7 9 13 1 9 9 0 1 9 13 2
13 15 3 13 9 9 3 2 3 0 9 0 15 2
33 0 7 2 16 9 9 7 9 3 13 16 1 15 9 2 13 3 9 9 9 7 9 3 13 9 13 2 7 15 13 13 0 2
28 7 3 15 12 3 13 2 16 0 3 13 1 9 2 7 16 9 2 13 0 2 13 9 15 13 1 9 2
42 16 7 13 9 9 9 7 9 13 1 9 13 2 13 1 9 9 0 1 15 13 2 15 4 0 13 1 9 13 2 3 13 1 9 7 9 9 2 15 15 13 2
23 7 3 9 0 3 13 13 0 2 16 3 13 13 9 0 2 1 13 3 1 9 0 2
13 3 3 13 13 9 12 9 0 15 13 7 15 2
21 1 15 3 13 13 12 13 9 15 7 15 2 1 9 13 9 15 13 9 9 2
17 7 13 2 1 15 16 13 12 13 2 16 13 12 7 15 9 2
11 7 15 13 0 16 9 0 13 9 0 2
21 15 3 13 12 9 13 0 9 13 2 7 1 15 13 16 12 9 1 0 13 2
14 3 3 13 9 0 9 16 13 0 9 0 1 0 2
30 7 1 15 13 16 2 16 9 0 13 0 9 7 15 9 2 16 3 13 0 9 2 7 9 3 2 16 15 9 2
16 3 3 15 15 13 13 9 2 13 15 15 13 13 0 9 2
30 13 3 13 15 9 0 7 13 2 16 13 15 9 13 9 3 13 1 15 0 2 15 9 13 2 7 3 0 13 2
8 7 15 15 13 9 13 9 2
21 15 9 13 16 2 1 15 16 13 9 9 0 0 9 2 13 16 1 9 13 2
19 7 3 1 15 1 15 9 13 1 15 9 13 2 13 3 13 0 9 2
18 16 7 9 13 3 1 9 2 15 13 15 15 13 9 13 9 0 2
19 9 7 0 13 1 10 9 2 15 13 9 0 2 16 7 10 15 9 2
21 3 2 1 9 0 3 13 0 2 3 13 1 9 13 1 15 16 13 0 9 2
2 3 2
39 1 9 0 2 16 3 13 0 9 9 15 13 0 1 12 9 2 16 9 7 9 2 3 7 9 15 13 0 1 10 9 2 16 15 9 7 15 9 2
25 15 7 9 13 9 1 9 0 7 13 0 9 0 7 12 2 7 3 15 9 13 1 15 9 2
28 15 3 13 2 3 1 15 16 9 13 1 9 0 13 0 9 2 3 9 0 13 12 1 10 2 7 0 2
2 3 2
21 9 0 2 1 9 13 2 13 0 1 9 0 9 2 15 3 1 15 13 0 2
15 7 13 13 16 15 0 9 13 9 15 15 9 0 13 2
19 1 9 3 9 2 16 15 3 13 2 13 9 15 15 13 1 9 9 2
18 3 3 13 2 16 9 0 13 12 2 16 9 0 13 1 0 9 2
40 16 7 13 16 9 0 1 9 0 13 2 3 13 15 13 2 7 15 13 2 3 3 13 16 1 9 15 9 15 13 2 7 10 13 2 7 9 15 13 2
6 10 7 13 13 0 2
11 12 9 1 0 2 13 3 15 3 13 2
13 15 9 1 0 2 1 16 13 1 15 9 9 2
40 3 7 9 7 9 0 13 15 9 0 2 7 13 15 13 7 13 9 0 2 15 13 13 1 0 2 7 13 10 7 9 0 9 2 15 13 13 1 0 2
11 7 1 15 1 9 7 0 13 1 9 2
12 1 15 7 15 13 4 3 0 9 13 9 2
21 16 3 13 9 1 9 7 9 13 9 12 2 9 3 0 13 2 9 7 3 2
26 13 3 9 12 3 1 15 15 13 2 3 3 3 1 9 0 15 13 2 7 3 1 15 9 9 2
16 3 3 13 16 15 9 9 13 9 1 9 16 9 13 9 2
17 3 3 15 13 9 15 15 1 9 13 2 7 15 15 1 9 2
16 9 3 3 13 9 0 2 13 9 1 9 1 9 10 9 2
10 9 0 13 9 1 9 1 9 9 2
13 1 15 3 13 9 0 2 15 9 1 0 13 2
7 9 3 13 9 13 13 2
33 13 3 16 2 1 15 9 1 12 0 13 2 9 15 13 1 15 9 3 13 15 9 13 1 9 9 13 2 16 13 1 0 2
20 3 3 13 1 9 7 9 15 9 0 13 1 9 9 2 7 9 0 3 2
22 15 0 13 9 1 15 9 13 15 0 9 13 1 13 9 9 2 16 13 1 0 2
11 3 1 9 0 13 15 0 9 1 9 2
23 7 3 9 9 0 9 3 13 9 2 7 3 13 1 9 2 16 9 10 13 1 9 2
16 9 7 9 0 9 13 7 1 9 2 7 1 9 1 9 2
12 0 3 1 9 9 2 1 9 0 2 13 2
15 1 15 7 15 13 13 7 9 7 9 2 9 13 9 2
13 16 15 3 1 0 9 13 2 9 15 13 13 2
12 3 7 9 2 16 15 13 13 2 13 13 2
8 15 7 9 0 13 9 13 2
25 1 15 3 15 13 2 13 9 0 1 9 2 3 9 2 7 15 15 0 13 2 3 0 9 2
17 7 3 9 13 0 2 7 1 9 2 1 9 2 7 1 9 2
51 13 3 15 9 13 13 16 13 13 13 2 13 3 9 9 9 1 15 13 2 16 10 9 1 13 13 9 2 7 15 9 1 9 13 2 7 13 9 0 2 1 15 1 9 9 13 9 0 1 13 2
42 7 16 0 9 13 15 13 16 13 9 0 9 2 15 13 15 0 2 3 1 9 13 16 9 13 9 13 2 9 7 0 13 2 16 7 9 13 9 9 1 13 2
21 3 3 13 9 1 9 1 9 2 3 9 0 9 2 7 0 2 16 13 4 2
33 3 2 1 9 13 13 9 9 13 1 9 0 16 1 9 2 9 9 0 15 13 1 15 16 13 12 9 9 1 9 7 9 2
15 9 3 0 13 3 13 15 1 0 2 1 13 9 0 2
12 3 15 9 3 13 1 13 2 1 15 9 2
12 16 9 13 3 13 9 13 2 7 15 9 2
31 1 15 3 13 13 16 7 9 13 13 12 1 10 2 16 9 3 13 2 7 9 2 15 3 13 9 0 13 12 10 2
16 1 3 9 7 13 13 13 2 13 16 15 0 13 0 0 2
13 9 7 0 13 1 13 16 0 0 7 0 15 2
18 13 3 15 1 15 13 16 9 1 9 2 16 13 1 12 1 9 2
31 16 3 9 0 13 15 9 0 2 13 1 9 9 2 16 13 4 2 7 9 13 13 3 3 2 7 3 13 12 10 2
2 3 2
32 9 13 3 13 9 0 9 16 15 1 15 13 2 0 16 9 13 2 1 3 13 1 9 2 7 16 1 15 13 9 0 2
13 3 3 13 15 16 15 15 13 9 0 1 13 2
8 15 7 13 15 15 13 15 2
7 3 10 9 13 15 0 2
8 13 3 9 13 13 9 0 2
17 7 3 2 1 9 0 13 9 9 2 9 13 3 13 9 13 2
2 0 2
23 16 9 0 13 1 9 0 2 15 13 1 9 2 3 9 0 13 1 9 13 1 9 2
52 7 9 0 13 1 9 0 2 3 1 9 15 9 13 3 2 7 1 9 9 15 9 2 3 15 13 1 9 2 16 15 9 13 1 9 15 13 1 15 9 7 1 15 9 2 16 13 9 1 12 0 2
41 16 3 9 0 13 9 9 7 3 13 9 13 2 16 13 4 2 9 13 2 1 15 9 13 9 0 1 15 2 3 13 15 9 13 2 7 15 9 0 9 2
2 3 2
16 9 13 9 1 15 13 1 9 2 15 13 13 15 9 13 2
9 15 3 9 9 13 1 12 0 2
14 13 7 16 9 10 13 1 9 13 16 1 0 9 2
23 16 3 9 13 13 15 9 13 2 15 13 7 0 9 1 9 15 7 0 1 9 13 2
2 3 2
31 16 9 13 13 15 9 13 2 13 16 15 9 13 0 7 3 13 2 7 3 13 13 16 3 13 7 13 1 10 9 2
9 9 7 15 13 13 9 0 9 2
10 7 3 15 3 13 2 7 3 3 2
12 16 3 3 2 3 3 15 13 1 9 10 2
10 7 3 13 9 16 9 13 0 9 2
17 3 13 16 7 3 13 2 7 16 3 13 1 9 10 9 13 2
2 3 2
24 9 9 13 1 10 9 15 13 1 15 9 2 13 12 2 16 9 9 13 12 1 10 9 2
18 9 7 0 0 13 13 7 0 2 7 1 13 15 9 13 1 15 2
8 0 3 13 0 1 9 13 2
5 15 3 0 13 2
29 13 7 13 16 9 13 3 13 3 1 15 13 2 7 3 3 9 13 0 9 2 7 0 16 13 1 15 13 2
16 13 7 1 15 1 9 0 9 2 15 9 13 1 10 9 2
9 7 3 13 9 13 1 10 9 2
32 7 1 15 3 13 16 3 10 9 13 15 15 13 9 2 16 3 10 13 9 9 0 13 2 7 0 15 13 13 7 13 2
10 13 7 16 15 9 3 13 3 13 2
45 15 3 9 15 13 1 0 1 13 2 13 16 13 7 9 9 0 1 13 9 0 1 9 13 13 2 16 9 13 2 7 16 13 9 16 13 0 9 2 16 9 7 9 13 2
8 0 7 15 3 13 13 13 2
14 16 9 0 1 10 9 13 1 9 1 9 0 9 2
13 3 13 1 15 16 0 1 9 7 1 9 9 2
39 3 7 13 15 1 15 9 13 13 9 15 2 13 0 1 9 15 2 16 9 13 1 15 0 9 2 16 9 9 13 1 9 9 1 9 9 7 9 2
15 15 7 0 13 1 9 0 15 13 13 15 9 0 9 2
25 3 9 0 3 0 1 9 3 13 0 2 16 13 9 1 12 0 2 1 12 13 9 13 15 2
32 9 7 15 13 1 9 9 13 7 13 2 13 2 3 1 15 16 1 9 0 13 15 13 2 7 1 15 16 15 15 13 2
22 3 3 2 3 1 15 13 2 9 0 13 15 9 16 13 9 0 1 9 13 13 2
2 3 2
20 9 13 0 9 1 9 1 0 13 10 9 1 0 2 7 1 13 1 9 2
39 16 3 15 9 13 1 9 13 3 13 10 9 1 9 0 2 7 0 13 15 1 13 2 3 13 9 9 1 9 0 16 9 1 9 2 16 9 13 2
2 3 2
31 1 15 9 3 13 1 15 0 1 13 2 7 1 13 7 9 2 7 0 1 13 2 3 13 7 13 9 0 1 13 2
49 15 13 9 0 2 7 1 9 9 9 7 9 15 13 9 2 1 12 8 7 8 8 2 13 16 1 9 13 9 2 1 0 9 12 9 2 1 0 9 0 9 2 15 13 9 9 7 9 2
14 13 7 15 9 9 0 15 15 1 9 9 0 13 2
24 13 3 16 10 9 9 0 1 10 9 13 9 1 13 9 15 13 1 9 1 9 13 13 2
21 3 7 2 15 9 2 13 16 9 13 9 0 2 9 7 0 13 1 9 13 2
28 0 7 16 1 0 13 9 1 15 16 13 0 9 7 13 9 0 2 13 3 13 16 9 13 13 9 13 2
25 15 3 13 13 0 9 13 16 9 9 13 0 13 1 0 9 2 0 7 9 13 1 9 13 2
9 15 13 1 9 9 1 12 0 2
18 3 3 13 0 15 13 9 0 1 13 2 16 9 9 1 0 9 2
2 0 2
18 9 0 1 15 9 13 3 0 1 9 0 2 7 13 9 10 9 2
7 9 3 13 9 7 9 2
31 7 0 13 1 15 9 9 16 15 0 9 1 9 3 9 13 2 1 9 0 10 9 2 16 13 1 9 13 1 9 2
11 13 7 13 0 9 15 13 1 15 9 2
15 3 3 13 13 1 15 9 13 2 16 3 13 9 0 2
8 15 3 9 1 9 3 13 2
10 3 15 13 10 9 13 13 1 9 2
2 3 2
5 9 9 13 9 2
36 3 9 13 1 9 3 13 1 9 9 9 2 7 0 3 2 16 13 1 9 0 3 2 1 16 9 2 1 12 8 2 13 15 13 9 2
15 9 7 15 13 1 9 2 13 1 9 9 0 7 9 2
23 15 7 9 15 13 13 9 0 1 9 2 13 1 9 10 2 3 0 1 9 9 13 2
11 3 13 1 15 13 15 0 9 15 9 2
6 15 7 13 9 13 2
12 3 13 3 9 13 2 7 15 9 9 10 2
2 3 2
12 1 9 15 13 13 9 0 1 9 0 15 2
23 7 16 3 9 15 13 1 9 2 13 15 9 0 2 16 13 1 9 9 0 1 9 2
21 16 0 9 15 13 1 9 2 13 15 9 0 2 16 13 1 9 0 1 9 2
9 9 7 13 9 1 10 9 13 2
38 15 7 0 7 0 9 13 13 2 15 3 13 1 9 15 2 16 9 13 1 0 2 7 3 1 9 2 16 9 13 0 1 9 13 0 1 9 2
25 13 3 1 9 9 13 15 0 9 3 9 13 7 0 2 7 15 1 9 1 9 9 13 13 2
2 3 2
16 16 9 13 13 15 9 13 2 0 13 16 13 1 9 9 2
30 9 7 15 9 13 0 9 15 0 9 2 13 9 0 2 16 9 13 7 13 2 7 15 3 15 0 9 9 13 2
28 1 3 9 3 13 13 16 9 9 13 2 16 9 13 13 15 9 13 2 13 16 13 3 13 9 0 9 2
14 7 3 9 3 13 13 1 15 16 13 0 7 0 2
2 3 2
12 15 13 16 1 15 9 15 0 1 15 13 2
20 3 9 2 1 12 1 9 2 13 16 15 13 7 13 2 13 9 7 9 2
14 7 15 9 2 3 9 0 7 9 13 2 13 9 2
13 9 3 13 1 9 2 7 13 9 0 1 9 2
14 3 3 15 1 9 15 9 13 16 15 1 15 13 2
23 13 3 16 9 15 13 15 9 2 3 9 0 7 13 2 13 9 15 1 15 0 13 2
47 16 7 13 16 15 9 13 9 3 13 9 13 15 2 16 9 13 2 3 1 13 4 16 9 9 0 15 2 16 13 15 9 13 2 15 15 13 2 3 13 1 15 16 1 15 13 2
7 0 3 13 1 9 13 2
34 13 3 9 13 1 9 0 13 1 9 0 2 16 9 1 9 0 15 1 9 13 1 9 2 16 13 1 9 9 1 12 1 9 2
13 9 7 9 3 13 9 9 2 7 0 9 0 2
13 3 7 9 15 9 13 1 3 9 9 9 13 2
24 3 7 9 2 1 15 16 13 1 15 9 0 9 13 1 9 13 2 13 13 9 9 13 2
2 3 2
25 15 15 3 13 13 1 0 9 16 1 15 16 13 1 0 9 2 3 13 1 13 16 15 13 2
21 3 9 0 3 13 1 13 16 15 13 2 16 10 9 15 13 1 9 0 13 2
24 9 3 2 13 1 0 0 2 13 1 9 2 7 3 1 9 13 1 10 9 1 1 9 2
34 9 7 0 9 13 13 2 15 0 9 13 9 13 2 15 13 9 0 2 1 15 13 3 9 0 2 15 13 1 9 2 13 9 2
18 16 3 9 13 13 15 9 1 9 2 15 9 9 13 1 9 0 2
12 3 3 13 9 13 15 2 7 9 1 15 2
14 7 3 3 13 9 10 9 2 7 13 9 7 9 2
13 7 13 15 9 0 7 9 0 2 15 13 9 2
10 3 13 3 9 13 9 13 1 9 2
14 16 3 13 0 9 0 7 13 1 12 9 9 13 2
56 13 7 3 15 15 13 0 2 16 12 7 15 9 2 3 10 9 2 13 1 9 1 10 0 2 15 13 1 9 0 2 7 13 15 9 2 15 13 9 13 2 1 15 13 1 16 13 1 9 2 7 1 16 13 9 2
15 3 3 13 16 13 7 0 9 13 1 12 9 9 13 2
12 16 15 7 0 13 2 15 9 7 0 13 2
23 15 3 13 15 9 15 13 1 15 1 9 7 1 15 1 9 2 16 1 9 0 13 2
14 9 3 13 9 0 7 9 0 2 9 7 1 0 2
11 15 7 9 13 13 1 9 0 7 9 2
26 13 3 9 0 15 1 9 1 15 9 13 1 9 2 7 1 15 13 1 9 15 1 9 9 13 2
27 13 3 9 9 0 9 2 7 2 16 1 13 13 2 1 15 13 9 0 2 16 10 9 0 13 3 2
27 1 15 7 3 13 16 13 15 7 15 9 13 2 15 13 1 15 16 9 10 15 7 15 9 13 13 2
10 10 3 9 13 1 9 13 1 13 2
21 13 3 15 9 0 1 9 1 13 9 9 0 1 15 2 15 13 9 9 0 2
11 7 15 3 13 9 9 0 13 15 9 2
30 15 3 3 13 1 9 0 2 1 13 9 9 0 3 1 9 0 2 15 13 9 0 2 7 13 3 1 9 0 2
6 3 3 13 0 9 2
27 7 3 2 16 1 15 9 15 9 13 9 2 13 13 9 0 13 1 10 9 13 2 13 0 1 9 2
14 3 3 13 9 1 9 2 9 7 9 9 1 9 2
8 1 0 7 13 1 9 0 2
23 13 3 1 9 0 9 0 1 9 2 13 15 0 9 2 7 15 9 9 13 9 13 2
22 13 3 1 15 9 15 13 1 9 1 13 9 9 0 2 7 15 13 9 9 0 2
16 13 3 15 15 13 1 9 2 1 15 15 13 1 9 0 2
17 16 3 12 13 1 9 1 15 1 15 9 15 1 15 9 13 2
16 3 9 9 13 1 9 1 9 9 15 9 15 13 1 9 2
18 7 3 9 0 2 15 13 1 9 2 15 9 13 7 13 1 3 2
46 9 7 0 3 13 1 9 1 9 9 15 13 1 9 1 9 15 15 13 3 2 7 1 16 15 9 13 1 15 9 2 16 3 4 13 1 9 13 0 2 1 15 13 0 9 2
12 7 3 9 9 13 1 9 13 9 9 0 2
12 7 3 9 9 3 13 9 2 7 9 13 2
14 1 15 9 13 16 15 13 1 0 16 9 1 9 2
42 15 7 9 3 0 13 16 9 2 3 1 15 16 13 0 7 0 9 2 13 3 1 9 16 13 9 13 0 9 2 16 15 9 13 10 9 9 0 15 13 9 2
12 1 15 1 9 13 3 2 1 9 0 0 2
15 13 3 0 9 2 3 0 9 13 2 1 0 7 13 2
22 15 3 0 13 1 9 10 16 1 15 15 13 0 2 15 13 16 9 9 1 9 2
14 3 0 9 0 15 13 15 0 2 13 1 10 13 2
23 16 7 9 0 10 9 0 13 1 13 9 9 13 2 13 16 15 13 9 13 9 13 2
13 13 3 9 1 9 1 0 2 16 9 1 0 2
11 16 3 3 3 13 2 3 3 3 13 2
19 15 7 0 15 9 0 0 13 2 9 13 13 0 1 15 2 3 9 2
11 3 3 13 15 0 13 9 13 1 0 2
22 16 7 15 13 0 2 13 16 2 3 15 13 1 15 3 0 2 3 13 1 15 2
5 15 13 13 0 2
17 3 3 13 15 0 15 13 9 0 2 15 1 15 13 0 0 2
27 3 9 4 13 1 13 16 15 15 13 15 0 2 3 13 15 13 0 1 15 2 7 16 13 1 0 2
9 3 13 16 13 9 15 15 13 2
6 7 15 13 9 13 2
13 1 15 3 13 9 13 2 16 13 0 15 13 2
10 15 7 3 13 9 9 0 15 0 2
21 3 15 13 15 9 10 9 13 9 9 13 2 7 0 1 9 9 13 13 9 2
20 16 3 13 9 9 1 9 13 16 13 9 13 2 7 3 16 13 15 9 2
31 16 0 0 9 1 13 13 13 15 13 9 9 13 13 1 9 15 16 15 15 3 13 1 9 13 2 16 13 9 13 2
62 13 3 2 0 2 16 2 16 1 10 9 13 15 16 9 1 15 9 2 7 15 13 1 9 1 10 15 13 15 9 2 7 15 9 13 3 0 2 15 13 10 15 13 15 9 2 16 15 13 9 1 9 2 0 13 7 1 9 13 15 9 2
23 7 3 3 2 3 15 1 9 13 16 9 2 13 9 2 0 2 1 15 13 10 0 2
39 15 0 2 15 1 9 13 16 13 9 2 13 9 1 15 13 10 13 2 3 0 1 9 2 2 3 9 13 2 15 13 16 9 2 7 3 16 9 2
14 15 7 13 9 13 9 2 13 13 16 13 16 9 2
18 15 3 9 9 13 9 9 13 9 9 2 16 3 13 15 0 9 2
8 15 7 1 0 13 9 13 2
17 1 15 0 13 16 9 13 3 13 9 13 2 7 3 15 9 2
18 13 3 13 16 9 0 7 13 13 9 9 2 7 16 13 1 9 2
7 15 3 15 13 9 13 2
2 3 2
6 9 15 15 15 13 2
46 16 1 10 9 1 15 13 9 7 9 2 13 15 3 9 2 15 13 1 9 1 15 15 13 15 9 2 7 15 3 9 2 15 13 9 1 9 2 16 1 0 13 9 7 9 2
23 7 9 0 13 15 9 1 15 13 9 7 9 2 1 3 13 9 13 7 3 1 9 2
40 13 3 1 9 9 0 15 3 9 2 15 13 1 9 1 10 0 2 15 13 9 0 2 7 15 3 9 0 2 15 13 10 1 9 2 7 13 9 13 2
26 15 3 9 2 1 9 9 2 13 1 9 9 2 7 3 15 13 1 9 1 9 15 9 13 9 2
2 0 2
12 9 13 16 9 13 13 16 9 15 13 9 2
14 9 7 3 13 16 15 1 15 13 2 7 15 13 2
18 3 13 3 9 13 15 9 13 1 15 13 2 7 13 15 9 0 2
17 3 7 13 9 9 16 9 13 13 9 9 13 2 16 13 9 2
11 13 13 9 13 10 2 15 13 16 9 2
37 15 3 13 9 9 2 16 9 9 3 13 2 16 13 9 13 1 15 15 13 15 0 1 15 7 16 13 2 1 15 16 13 1 15 15 0 2
15 13 3 13 9 3 15 13 2 7 9 15 13 10 13 2
29 7 3 13 13 16 9 13 13 9 1 9 15 9 13 1 0 9 9 2 1 16 15 13 9 13 13 9 9 2
40 16 9 15 9 4 13 1 0 2 16 13 9 1 12 0 2 7 3 13 16 13 9 9 13 2 15 13 9 2 15 4 13 1 9 2 13 13 1 9 2
20 7 13 9 1 16 13 1 9 7 9 2 16 10 9 7 9 13 13 9 2
17 7 15 13 2 16 13 15 9 9 13 13 9 16 9 9 13 2
21 3 13 2 16 15 9 2 3 13 2 13 13 7 0 7 0 7 9 9 13 2
25 15 7 12 15 13 9 13 2 12 1 13 1 9 0 13 2 3 16 13 0 7 16 13 13 2
11 0 2 3 16 13 0 2 1 9 13 2
30 13 3 0 16 3 13 0 16 9 2 7 3 13 16 2 0 13 13 2 0 13 2 16 3 13 1 9 1 0 2
24 0 0 3 13 1 9 0 2 13 16 13 1 9 1 0 2 7 15 15 13 9 1 13 2
11 3 3 1 12 0 9 0 13 1 13 2
8 1 0 9 13 7 9 13 2
9 1 0 7 3 13 13 1 0 2
11 15 12 9 13 13 1 12 9 2 13 2
15 3 3 0 13 9 0 2 7 9 2 3 0 2 9 2
16 1 3 13 16 9 13 13 16 9 0 2 7 0 16 9 2
10 1 15 7 0 13 12 0 2 3 2
7 9 13 0 0 7 9 2
20 7 0 2 15 13 16 0 7 9 2 13 13 7 0 2 16 1 13 4 2
5 3 0 3 9 2
8 15 0 1 15 0 3 13 2
25 9 1 15 13 0 0 7 9 2 16 13 1 15 16 9 7 9 9 1 0 7 9 1 9 2
10 9 7 0 13 0 3 7 9 9 2
12 9 3 13 13 9 3 13 2 7 9 9 2
36 13 7 16 7 1 15 9 9 13 13 16 9 13 13 15 9 13 2 7 16 13 13 15 9 15 1 13 1 0 2 3 16 3 13 9 2
24 16 7 13 16 13 9 9 13 2 3 13 15 16 9 9 13 1 9 2 16 1 13 4 2
3 3 13 2
8 15 7 13 1 9 9 9 2
11 1 15 9 13 16 13 9 13 1 0 2
15 3 1 9 13 15 13 13 7 13 2 3 7 1 0 2
8 15 7 0 13 1 9 9 2
21 3 1 15 9 13 1 9 0 2 16 13 1 9 0 16 15 0 13 16 0 2
15 1 15 3 15 1 9 13 2 15 13 9 7 15 13 2
12 9 3 0 2 7 15 13 4 2 15 13 2
30 0 3 1 15 16 9 0 2 16 13 9 13 2 15 13 1 15 15 13 2 13 13 16 9 0 13 16 15 0 2
19 7 9 1 13 16 9 0 13 9 3 0 2 7 15 9 13 16 13 2
15 3 13 13 13 16 1 15 16 13 9 2 13 15 0 2
22 7 13 0 16 15 13 1 9 0 2 16 15 3 1 13 1 9 7 0 1 9 2
33 9 3 13 9 1 9 0 1 9 2 7 0 9 0 13 9 1 9 0 9 2 7 15 9 9 1 9 13 15 0 1 9 2
34 13 3 13 16 2 16 9 13 1 9 0 7 13 2 15 13 13 1 9 1 9 2 13 16 9 1 9 13 15 9 13 1 9 2
3 3 13 2
18 15 0 1 9 2 9 0 1 12 13 2 3 7 2 7 1 9 2
40 15 3 9 1 9 7 9 1 0 9 13 2 3 16 9 1 9 13 0 9 2 9 0 2 1 12 7 15 15 13 1 9 1 9 2 13 0 9 9 2
22 0 0 13 2 3 13 9 3 9 0 9 2 16 9 3 13 1 9 16 1 9 2
33 13 3 16 9 15 13 1 9 2 7 0 2 16 13 1 9 2 0 13 9 16 9 1 9 2 7 15 13 1 12 7 15 2
33 3 3 3 2 3 0 2 16 9 0 13 1 9 1 9 13 2 15 13 9 2 16 13 2 7 3 1 15 9 0 13 9 2
19 3 13 1 12 8 2 16 1 13 13 15 13 16 13 1 9 1 9 2
20 3 3 1 9 15 13 9 9 0 2 16 13 1 9 2 1 9 1 9 2
3 3 13 2
11 7 3 3 3 13 2 7 3 3 13 2
11 1 15 13 9 9 1 9 7 9 0 2
32 1 3 13 1 9 0 16 3 3 13 2 7 3 3 13 2 16 13 1 9 1 0 2 3 13 2 16 3 13 9 15 2
15 9 7 1 15 13 9 16 13 15 0 2 16 3 13 2
11 3 3 13 15 3 13 7 3 3 13 2
3 3 13 2
8 13 7 15 0 15 0 13 2
7 15 3 13 13 1 13 2
15 3 3 15 0 13 13 2 16 3 15 13 1 9 0 2
13 7 13 13 1 0 2 16 3 15 13 1 13 2
54 13 3 16 13 1 15 15 13 15 2 3 1 9 1 9 2 1 15 13 2 16 15 0 1 9 10 13 13 2 3 13 9 2 15 13 1 9 1 9 2 3 2 15 9 9 15 13 9 2 13 0 7 13 2
22 7 3 13 16 15 0 9 13 0 7 0 2 3 1 9 3 13 2 1 13 13 2
10 16 9 0 2 13 9 2 3 13 2
14 1 13 3 0 13 13 9 0 3 13 2 13 9 2
10 13 4 3 1 10 9 0 13 0 2
12 9 7 9 13 15 9 0 2 16 13 4 2
7 13 3 9 0 0 13 2
2 3 2
11 15 9 13 1 15 1 15 13 10 9 2
12 15 3 9 13 0 2 3 1 9 7 9 2
11 9 7 9 0 13 1 9 15 1 9 2
7 13 3 9 9 7 9 2
11 1 9 7 3 3 13 3 3 0 13 2
21 9 7 9 13 1 15 16 9 9 9 3 13 2 7 15 1 9 13 7 13 2
12 3 3 9 9 13 1 15 16 1 9 13 2
26 16 7 13 16 9 9 13 1 9 15 1 9 1 9 2 9 7 1 9 1 9 2 3 13 13 2
26 9 3 9 13 9 7 9 15 2 16 15 13 1 16 13 9 2 7 0 9 9 13 0 15 9 2
14 3 13 3 13 9 15 9 16 1 16 13 15 9 2
26 16 3 9 1 9 10 13 1 13 9 2 0 9 10 1 9 10 3 13 1 15 16 1 9 13 2
2 3 2
9 0 0 9 1 9 13 15 0 2
11 0 3 9 9 2 16 3 2 13 13 2
11 1 15 3 13 1 0 7 9 7 0 2
9 13 7 0 13 7 0 16 3 2
7 9 7 13 13 0 13 2
6 3 9 0 13 0 2
2 0 2
7 0 13 9 0 13 3 2
7 7 9 0 13 0 13 2
12 15 13 1 15 16 9 13 15 1 10 13 2
18 9 7 1 9 13 13 3 0 16 3 2 16 0 9 2 7 0 2
16 13 3 9 9 1 9 2 15 13 0 7 1 10 9 13 2
2 3 2
16 15 15 13 1 15 2 13 1 15 1 9 15 1 15 13 2
12 9 7 9 13 1 9 0 16 13 0 9 2
15 13 7 0 9 16 13 0 2 0 2 7 1 13 0 2
6 3 9 0 13 0 2
14 7 2 16 1 4 13 2 9 0 13 15 9 0 2
6 13 3 9 0 0 2
2 3 2
8 9 0 13 13 16 9 0 2
23 7 15 15 15 13 1 9 0 1 9 0 13 2 13 0 1 10 9 2 3 9 0 2
12 0 3 0 9 0 2 15 13 0 9 0 2
14 3 7 9 0 2 15 9 0 13 9 2 13 0 2
2 0 2
10 13 13 0 13 2 16 3 9 13 2
12 7 9 13 13 9 0 2 16 1 13 13 2
18 1 3 0 9 2 16 3 2 13 0 2 0 0 9 13 13 0 2
16 3 7 9 0 2 15 9 13 9 13 2 16 1 13 13 2
2 3 2
21 15 9 13 16 7 1 9 0 2 7 1 9 10 9 2 7 1 9 10 9 2
12 1 9 3 0 2 16 9 13 1 9 0 2
14 1 9 7 10 9 2 16 2 13 9 13 9 0 2
18 1 9 7 9 2 16 9 9 13 13 9 9 2 15 13 15 9 2
10 7 9 0 3 13 13 1 9 0 2
19 3 13 3 15 15 0 2 1 1 9 0 15 13 0 7 0 10 0 2
8 0 7 7 1 9 10 9 2
17 13 4 3 1 16 9 0 13 9 3 13 1 9 1 10 9 2
21 0 7 7 1 9 10 9 2 16 3 13 13 15 9 16 0 2 16 1 13 2
8 15 3 9 9 0 13 13 2
2 3 2
16 16 9 13 1 9 9 2 13 16 15 9 13 1 9 9 2
34 16 7 15 9 9 13 13 9 2 15 3 13 16 1 9 2 16 3 9 9 13 9 0 2 16 9 13 13 9 2 1 9 3 2
5 15 1 15 13 2
15 16 3 15 9 1 15 13 15 9 2 3 13 9 13 2
19 13 7 16 2 15 9 0 13 13 2 16 9 13 2 16 9 0 13 2
22 3 13 9 2 1 12 1 9 2 16 2 16 0 13 9 0 2 13 3 16 0 2
36 1 3 9 13 9 9 15 3 13 9 2 16 1 13 13 2 15 3 13 2 7 1 15 7 1 9 2 1 9 7 1 15 15 9 9 2
37 16 7 1 9 9 13 9 7 9 1 9 9 2 15 3 13 1 9 15 9 2 7 1 9 9 15 9 13 2 3 9 2 0 7 0 9 2
7 13 3 16 9 13 0 2
11 3 7 9 0 2 15 13 0 15 9 2
7 15 3 13 1 9 9 2
19 13 3 2 1 12 1 9 2 16 9 13 9 15 13 2 7 3 13 2
22 16 7 15 3 13 13 1 15 9 13 15 13 9 0 7 13 2 1 13 13 13 2
10 3 13 1 15 9 9 1 12 0 2
23 3 13 2 1 9 13 2 16 9 13 13 2 9 0 0 13 3 1 15 15 13 9 2
13 16 3 13 9 2 3 9 13 2 7 3 0 2
10 1 15 15 9 13 9 9 13 9 2
17 7 15 13 2 3 13 2 16 7 7 0 15 13 2 13 13 2
18 3 1 15 15 13 2 16 16 13 9 15 2 3 10 2 7 9 2
26 1 15 13 2 1 13 1 9 2 16 13 9 2 15 13 9 9 2 1 9 13 2 3 1 9 2
31 13 7 1 13 9 9 16 2 16 13 9 13 9 2 3 3 13 15 3 13 7 1 13 0 2 16 9 9 15 13 2
20 3 1 9 15 9 9 0 13 2 13 15 1 9 13 2 7 9 15 13 2
7 13 7 9 0 9 13 2
8 13 3 1 9 1 8 9 2
21 0 9 13 13 9 0 2 15 7 13 9 13 2 7 9 10 7 9 0 13 2
21 7 1 9 13 2 16 9 13 2 7 1 0 9 2 16 9 2 16 0 13 2
16 1 15 7 13 9 0 2 1 15 9 9 13 2 8 12 2
13 1 15 13 4 2 7 1 15 13 16 3 13 2
10 7 1 15 9 9 13 2 8 12 2
12 12 13 9 9 7 9 2 7 0 15 9 2
9 16 13 9 2 3 7 15 13 2
11 0 13 10 2 7 15 13 9 9 0 2
21 16 3 3 1 9 10 7 0 13 2 13 1 15 16 1 9 9 3 13 13 2
18 16 13 9 1 9 10 3 13 2 7 9 13 1 15 15 13 15 2
11 0 3 13 9 0 9 15 9 9 13 2
12 9 13 9 13 13 9 2 7 9 15 2 2
14 13 7 15 9 13 13 9 0 3 13 13 1 9 2
26 16 3 9 0 13 1 9 9 2 16 1 13 4 2 13 3 9 2 3 13 9 1 10 9 13 2
20 3 13 15 12 13 2 7 16 0 9 0 13 13 2 7 16 13 12 3 2
19 15 13 13 1 9 15 15 13 13 0 0 15 15 13 12 1 10 9 2
21 7 15 13 9 13 3 2 16 9 13 2 7 1 13 3 0 2 16 13 9 2
2 0 2
8 9 0 13 9 9 1 9 2
15 7 2 16 13 0 9 1 9 9 2 13 15 13 0 2
19 16 3 15 13 15 13 12 1 9 2 3 0 13 15 13 0 1 9 2
13 3 13 7 13 1 9 13 1 9 9 16 0 2
18 3 3 13 13 1 9 7 9 2 16 1 13 4 1 10 9 0 2
8 13 3 16 13 0 1 9 2
22 3 7 1 9 9 13 9 1 15 9 2 16 10 15 13 1 9 1 9 2 13 2
15 13 3 16 3 16 13 1 9 13 2 13 1 9 0 2
7 9 7 13 9 1 9 2
9 3 7 9 9 13 1 9 0 2
4 15 13 9 2
11 3 0 13 16 9 0 0 13 1 9 2
2 3 2
22 13 3 13 0 2 1 13 9 9 2 13 16 9 0 1 10 9 13 1 9 9 2
12 16 3 9 13 1 0 2 9 13 1 0 2
6 3 7 9 13 0 2
13 7 16 9 13 0 2 0 9 13 4 1 15 2
23 16 3 9 13 13 1 9 1 10 9 2 13 13 9 0 13 3 1 9 9 0 13 2
5 15 7 13 0 2
9 3 0 9 3 13 13 1 9 2
16 13 3 2 16 9 13 0 2 16 9 3 13 0 1 9 2
2 3 2
15 15 13 15 7 13 1 15 1 10 9 2 13 15 0 2
6 15 3 13 9 9 2
15 16 3 9 3 13 9 13 2 13 16 9 0 9 13 2
15 3 9 13 9 1 9 2 15 13 13 1 9 7 9 2
10 7 13 0 16 3 13 15 9 0 2
13 3 3 1 15 15 13 1 9 2 13 9 12 2
8 3 9 0 3 13 15 9 2
2 0 2
11 0 13 15 9 13 15 3 13 15 9 2
8 7 10 9 9 13 1 9 2
6 15 3 13 1 9 2
36 3 9 9 0 13 1 9 0 2 7 1 9 0 2 7 1 15 9 15 13 1 9 2 15 13 7 13 2 7 1 15 13 9 1 9 2
37 9 3 10 9 15 13 1 9 0 2 13 1 9 0 2 7 15 15 13 1 15 9 0 2 16 15 13 9 9 2 16 9 2 9 7 3 2
29 13 7 16 3 13 9 1 15 9 0 13 2 3 9 15 13 9 2 15 3 15 13 1 15 16 9 1 9 2
19 3 2 16 9 3 13 13 1 9 2 3 9 0 3 13 13 1 9 2
21 13 3 9 1 13 9 13 9 1 15 16 13 0 9 2 3 9 0 7 0 2
22 1 15 13 16 2 1 13 9 15 9 9 1 15 13 2 16 3 13 13 1 9 2
28 3 7 9 13 16 3 1 9 13 9 2 7 16 15 13 1 9 0 2 15 13 9 0 2 15 13 0 2
24 7 1 15 13 2 1 12 1 9 2 16 13 9 13 15 0 13 2 3 9 7 0 9 2
20 7 1 12 1 9 2 13 16 3 13 2 1 9 2 15 15 13 1 9 2
12 3 3 13 16 15 9 9 13 13 1 9 2
14 7 3 9 15 13 2 1 15 9 13 13 1 9 2
18 15 7 9 2 16 0 13 2 16 1 13 4 13 2 13 13 13 2
24 7 0 13 13 16 15 13 13 3 13 7 13 2 3 13 9 7 9 2 15 1 10 9 2
24 16 3 9 12 13 1 15 2 9 7 9 15 3 1 15 13 2 3 2 1 15 9 0 2
23 9 3 7 9 3 13 13 1 3 13 7 3 0 13 2 16 0 9 1 0 9 13 2
15 3 3 13 16 9 7 9 13 15 3 1 9 7 9 2
18 16 3 9 9 13 1 9 2 9 15 1 9 13 2 7 0 9 2
22 16 7 3 2 13 3 0 13 9 1 9 9 2 3 3 1 9 2 7 9 15 2
13 3 7 3 16 13 9 7 9 15 9 1 9 2
16 13 4 7 16 9 0 13 9 1 10 9 1 9 3 13 2
20 3 13 16 13 3 9 1 16 13 9 2 3 3 9 9 13 9 9 9 2
18 7 3 3 13 16 2 13 9 2 13 9 9 2 16 0 9 13 2
11 1 15 3 1 0 13 9 1 0 9 2
25 3 3 15 9 9 13 9 1 9 2 7 0 15 15 13 1 9 0 2 7 1 0 9 9 2
23 13 3 16 15 13 9 9 15 9 7 15 2 7 3 13 15 9 7 15 9 1 9 2
22 9 3 9 1 9 13 13 3 9 9 1 9 2 16 15 13 9 15 9 7 15 2
28 3 3 15 9 13 1 9 9 0 15 9 2 7 13 1 0 9 9 2 7 13 1 0 9 9 1 9 2
20 15 3 9 13 13 15 9 7 3 15 2 15 7 15 2 7 3 1 10 2
25 3 7 9 13 1 9 3 13 9 2 16 7 15 15 9 13 2 3 1 9 1 9 3 13 2
9 13 3 9 1 9 10 9 9 2
22 15 0 9 13 2 7 3 1 9 7 9 3 13 12 1 15 2 7 12 1 9 2
11 16 7 9 13 2 13 15 13 9 13 2
16 3 13 16 15 0 9 13 1 9 13 2 7 1 13 9 2
16 9 7 0 9 13 2 15 9 9 13 1 0 9 0 13 2
14 15 3 9 0 13 2 13 9 0 1 9 3 13 2
32 15 0 13 16 1 10 9 13 15 12 13 15 13 10 0 2 3 9 13 2 1 15 2 7 1 15 9 0 2 1 15 2
29 15 7 13 9 1 10 9 1 9 13 2 7 2 16 13 9 13 9 2 13 15 9 0 9 13 1 13 9 2
11 7 15 13 0 9 2 1 15 1 13 2
17 15 0 2 10 13 13 2 13 3 13 9 9 13 9 13 0 2
19 9 3 0 9 1 15 15 3 13 1 3 9 2 13 9 0 1 9 2
6 15 13 3 13 9 2
7 7 13 9 9 7 9 2
19 15 7 15 9 13 2 1 15 13 3 13 2 1 3 13 9 9 13 2
11 0 3 13 9 9 1 15 13 3 13 2
26 3 1 12 8 7 1 12 9 7 9 2 13 3 13 0 9 1 9 0 2 3 7 1 9 0 2
18 0 3 13 1 15 15 9 13 0 9 9 2 15 9 9 3 13 2
23 3 13 3 0 2 16 16 9 13 9 13 2 16 4 15 0 13 2 16 0 9 13 2
4 9 3 13 2
14 15 13 13 7 13 1 9 9 13 1 9 7 9 2
12 16 7 13 1 9 9 13 2 0 3 13 2
16 13 3 9 0 0 7 0 13 2 16 13 9 1 12 9 2
10 3 2 13 9 2 13 1 10 9 2
10 3 3 9 0 15 13 2 7 0 2
7 13 3 15 1 9 12 2
14 0 7 9 13 9 1 9 12 2 16 1 13 4 2
14 3 2 16 13 1 9 2 0 15 13 2 3 0 2
40 16 7 9 0 3 13 9 1 9 16 1 9 15 9 2 9 7 0 13 1 9 15 2 1 15 13 16 9 0 13 9 7 9 2 9 7 0 9 9 2
21 15 7 0 9 13 2 15 9 13 13 1 9 16 1 9 13 2 13 13 0 2
10 13 3 9 15 15 1 9 3 13 2
7 3 7 13 13 7 13 2
18 15 7 1 9 0 13 2 16 13 9 9 0 7 0 2 3 13 2
21 13 3 13 16 15 9 13 9 13 1 9 7 9 13 2 16 7 15 9 13 2
9 15 3 1 15 13 1 15 13 2
28 9 3 9 0 16 13 9 13 2 16 13 0 1 9 3 13 2 3 9 15 15 7 9 15 13 13 9 2
31 3 7 13 9 0 15 2 15 13 13 2 16 3 13 1 9 3 1 9 0 13 2 13 3 9 1 9 2 3 9 2
34 3 2 16 13 9 1 9 2 3 13 13 1 9 2 7 3 13 16 1 9 0 7 0 2 1 15 9 13 2 16 1 13 13 2
18 7 1 15 13 2 3 1 15 9 2 7 0 13 2 13 9 13 2
10 9 0 13 9 13 15 0 1 9 2
46 3 7 15 9 2 15 13 13 2 13 1 9 1 15 9 1 0 9 13 2 15 13 9 2 7 13 1 15 2 1 9 9 15 13 0 1 9 1 9 13 2 1 15 1 13 2
15 1 15 3 16 1 0 2 0 9 13 13 1 9 13 2
7 15 9 3 1 0 13 2
18 3 9 2 16 13 1 9 1 9 0 2 13 0 1 13 15 9 2
19 3 7 9 9 2 15 1 0 9 13 9 2 0 13 9 1 13 0 2
34 9 3 13 2 16 0 9 3 13 2 7 13 15 9 9 7 9 13 2 13 1 13 2 1 0 9 2 15 15 9 9 0 13 2
19 7 15 0 3 13 1 13 7 9 13 2 3 3 13 9 1 0 9 2
5 7 0 15 13 2
34 16 2 1 9 0 2 16 1 13 4 2 1 0 9 7 0 9 2 3 1 9 13 9 7 9 2 13 1 9 2 13 1 0 2
25 3 7 2 16 0 13 1 9 13 2 9 13 9 13 3 1 9 13 2 7 0 9 15 13 2
22 3 3 2 16 13 10 1 9 0 9 2 13 9 13 2 13 3 15 9 13 9 2
41 13 7 2 1 13 9 1 0 9 13 2 16 1 9 1 9 7 8 9 13 2 3 13 1 9 1 9 13 2 16 13 0 13 1 9 15 15 15 0 13 2
26 15 13 9 13 13 3 15 15 13 1 9 2 1 9 0 1 9 0 0 13 2 16 1 13 4 2
20 1 15 0 9 9 2 16 13 13 2 13 2 7 15 3 2 13 9 13 2
8 3 3 13 16 13 9 9 2
16 7 3 13 9 0 9 1 0 7 0 2 1 15 9 0 2
18 7 3 1 9 13 3 13 1 9 2 16 9 13 1 9 1 9 2
13 13 7 3 1 0 9 9 2 15 13 1 9 2
30 3 9 13 2 1 12 8 2 16 9 12 0 9 13 2 7 1 12 2 16 1 9 9 13 9 0 2 7 13 2
28 1 0 9 13 9 3 13 9 2 16 7 9 2 3 13 3 2 1 16 13 9 9 2 1 9 13 13 2
13 3 3 1 13 9 13 3 13 9 9 13 0 2
8 16 9 0 9 3 13 0 2
15 1 15 7 15 13 4 2 0 13 0 9 3 13 0 2
14 3 3 13 4 16 15 9 0 9 13 1 9 13 2
14 1 9 7 0 3 13 13 15 9 0 9 0 9 2
6 3 3 13 7 13 2
23 15 1 15 13 2 16 10 9 15 9 0 13 2 3 1 9 13 7 3 1 9 13 2
13 10 3 9 0 13 9 2 7 10 9 0 9 2
12 15 3 13 9 9 0 15 13 13 1 9 2
16 1 3 10 9 15 9 13 2 3 13 9 0 1 9 13 2
7 3 2 13 9 2 13 2
2 3 2
10 10 9 13 1 9 4 13 1 9 2
19 3 3 9 13 13 9 0 9 2 16 13 15 2 16 1 1 13 13 2
15 7 2 16 9 0 13 13 9 2 13 9 1 9 13 2
7 3 13 9 13 1 9 2
20 7 1 13 1 9 15 13 13 7 13 2 16 9 13 2 1 12 1 9 2
12 3 9 0 2 16 1 9 13 2 13 0 2
4 15 13 0 2
2 3 2
16 1 15 9 15 13 13 1 15 9 2 13 0 9 15 9 2
14 0 3 13 15 10 13 2 3 3 16 15 0 0 2
40 1 0 7 3 13 15 9 1 9 0 2 16 16 13 1 9 2 16 1 15 13 9 9 2 1 15 9 13 2 15 3 13 7 1 9 7 1 9 0 2
17 3 7 3 1 0 9 9 16 13 9 2 15 13 9 9 13 2
19 3 2 1 9 0 3 13 16 15 7 3 2 0 13 16 13 9 0 2
6 7 3 13 9 0 2
9 3 13 3 9 0 0 0 9 2
2 0 2
28 1 9 9 13 2 16 13 1 9 1 12 8 2 1 15 13 9 15 9 16 1 9 1 15 10 9 13 2
10 9 7 0 9 10 13 1 13 9 2
26 3 3 13 1 0 2 9 7 9 2 16 1 16 13 0 9 7 0 2 1 15 13 10 15 9 2
13 15 3 9 15 13 1 9 9 0 16 1 9 2
9 3 3 13 15 15 9 1 9 2
8 15 7 9 9 0 9 13 2
15 13 3 8 12 2 1 9 0 2 9 15 1 9 13 2
3 3 13 2
7 1 9 9 9 15 13 2
7 7 1 9 1 8 9 2
18 0 9 13 9 0 13 2 3 1 15 0 2 0 9 1 9 13 2
21 9 3 2 1 12 1 9 2 13 16 0 9 9 13 1 15 16 0 1 0 2
14 1 15 7 13 9 9 2 15 13 3 0 9 0 2
9 13 3 13 13 0 9 13 0 2
16 15 3 13 15 9 1 15 13 2 7 15 13 1 15 0 2
19 7 9 0 1 0 13 15 9 1 15 1 15 3 13 9 2 3 13 2
15 3 13 13 1 12 2 15 12 13 13 7 15 13 13 2
14 3 2 1 9 13 13 2 13 16 9 0 13 13 2
6 3 13 1 15 0 2
10 3 3 13 1 9 13 2 9 13 2
13 15 3 0 1 9 13 15 1 15 3 13 9 2
18 1 15 7 3 13 13 2 1 7 0 13 2 7 13 1 0 13 2
7 13 3 16 13 3 0 2
29 1 15 3 13 13 9 9 15 13 10 9 13 0 2 16 3 9 13 13 15 2 10 7 13 15 13 13 0 2
11 9 3 3 13 16 13 15 1 15 13 2
8 15 7 1 15 3 13 13 2
13 3 13 2 1 15 2 16 13 15 3 13 13 2
13 7 3 13 16 9 10 9 13 0 2 3 0 2
42 3 7 15 9 1 15 13 13 1 13 2 16 1 2 1 9 9 2 15 13 16 13 2 15 15 13 15 13 2 13 1 15 9 2 7 3 13 15 9 1 15 2
18 3 0 7 1 13 2 7 3 1 13 13 9 9 0 0 9 13 2
22 13 3 16 13 13 9 15 15 9 13 2 7 15 2 3 13 2 13 9 1 13 2
13 3 2 13 9 2 13 16 13 9 9 1 9 2
10 15 7 15 13 4 2 13 13 0 2
10 3 3 13 13 13 2 7 3 13 2
16 3 1 9 13 13 9 9 13 1 0 2 1 15 9 13 2
30 3 7 13 13 0 9 13 1 0 16 13 9 1 0 2 16 3 13 13 13 9 9 1 0 9 2 16 13 13 2
21 3 9 13 9 1 9 1 9 7 0 9 2 15 13 9 9 2 3 7 9 2
12 15 3 13 16 9 13 0 2 9 0 0 2
23 3 13 16 9 13 1 9 1 16 13 1 9 2 3 7 9 2 7 1 16 13 0 2
13 9 3 9 13 1 9 0 2 3 7 9 9 2
2 3 2
14 0 9 13 0 0 0 2 16 9 9 2 9 0 2
10 15 7 9 0 1 9 0 9 13 2
17 3 9 9 13 13 1 9 1 10 9 2 9 9 1 10 0 2
16 16 7 15 9 13 1 9 0 2 15 9 13 10 0 0 2
17 3 9 0 15 13 0 2 3 1 15 13 2 1 10 3 9 2
13 3 9 2 15 3 13 9 0 2 10 0 13 2
8 13 3 3 13 1 9 0 2
2 3 2
25 9 13 1 9 0 2 3 7 9 2 16 15 13 9 0 2 3 0 13 15 13 2 7 3 2
14 15 3 9 13 9 9 1 0 2 7 9 1 0 2
8 9 3 9 13 1 9 0 2
14 9 0 9 1 9 0 2 15 9 13 1 0 9 2
20 15 7 9 13 2 9 13 13 15 2 0 13 13 1 15 15 1 9 13 2
9 15 3 9 13 13 16 4 13 2
7 3 9 13 10 13 13 2
22 7 3 3 13 1 0 16 15 13 1 15 13 2 13 0 13 1 15 9 13 15 2
19 7 1 15 13 9 2 15 13 0 13 1 9 9 2 13 15 13 15 2
8 15 7 13 13 0 2 0 2
16 0 3 2 16 13 4 16 10 15 13 1 15 2 13 9 2
16 3 2 1 9 3 13 9 2 0 13 15 13 16 1 9 2
28 0 16 2 1 13 16 3 13 9 2 13 7 16 3 13 1 9 2 15 7 13 13 1 15 9 7 9 2
32 0 13 16 15 1 15 13 13 7 13 2 7 13 2 16 15 13 13 15 2 16 12 9 15 13 13 7 15 9 13 13 2
18 7 15 9 13 9 13 15 2 16 9 13 13 2 7 9 13 13 2
36 7 16 9 9 3 13 13 9 2 16 13 9 9 2 15 0 9 13 2 3 3 1 15 9 0 13 13 2 7 13 9 0 1 15 9 2
18 16 3 9 13 2 1 12 1 9 2 16 13 7 13 13 9 15 2
14 3 7 9 3 13 9 13 1 9 2 7 9 9 2
34 3 2 1 13 9 13 15 2 13 1 15 13 16 15 13 1 9 9 2 1 0 15 15 13 1 15 9 2 15 3 13 1 9 2
9 3 3 9 13 13 2 7 0 2
10 1 15 13 13 10 9 9 13 0 2
20 3 15 1 15 13 9 2 7 1 15 13 9 2 7 1 15 9 13 13 2
19 7 3 13 4 16 9 9 0 2 15 13 13 2 3 13 13 1 9 2
12 0 7 3 15 13 1 9 15 15 13 13 2
16 3 10 15 1 9 0 9 13 2 0 1 9 15 9 13 2
6 3 7 9 9 13 2
14 1 15 13 16 7 15 13 13 9 9 0 1 9 2
11 3 3 13 9 0 16 1 9 7 9 2
14 3 9 15 13 13 9 2 13 9 13 9 9 9 2
13 3 3 13 9 13 9 1 13 2 16 9 13 2
13 3 3 13 16 15 9 9 0 13 13 1 9 2
13 1 15 1 9 13 13 16 9 0 1 9 13 2
7 16 9 0 13 1 9 2
37 7 16 15 9 13 7 13 13 7 9 13 13 2 13 15 13 16 2 1 15 9 0 9 13 3 13 2 16 7 9 13 13 2 7 13 3 2
8 15 3 13 15 9 13 13 2
13 3 15 15 3 13 13 2 13 9 16 13 3 2
29 15 7 13 9 16 13 3 3 1 15 0 13 13 3 13 2 16 3 15 13 9 13 2 3 9 13 1 9 2
13 10 7 15 13 13 2 13 3 0 13 3 13 2
11 15 3 3 13 13 2 7 13 3 13 2
2 3 2
17 9 0 2 16 13 0 2 3 2 3 13 1 15 2 13 0 2
4 13 3 0 2
17 10 7 0 13 0 2 16 15 0 13 13 2 0 13 3 13 2
11 1 9 7 9 0 13 9 1 9 0 2
12 0 3 9 2 1 15 9 13 13 9 9 2
2 0 2
11 15 3 13 9 15 0 10 0 9 13 2
19 13 7 0 9 0 13 0 9 2 1 15 9 13 4 1 13 9 0 2
27 16 3 3 1 0 15 9 0 13 13 15 9 13 2 13 3 0 0 0 9 13 2 7 0 15 13 2
6 13 3 0 13 0 2
4 15 13 0 2
9 3 3 15 13 1 9 0 9 2
23 13 3 8 12 2 16 9 9 0 13 9 10 15 13 2 7 13 1 10 9 15 13 2
10 15 7 3 13 16 3 0 9 13 2
15 3 3 1 0 9 0 13 13 2 7 1 9 9 13 2
26 1 15 3 7 0 9 15 2 9 9 13 2 13 9 0 2 16 13 0 2 3 7 1 0 13 2
40 3 15 13 9 0 1 15 9 13 0 2 3 0 2 13 15 1 0 13 2 7 3 3 9 13 2 3 7 1 9 13 2 15 9 1 13 9 9 13 2
49 15 0 13 9 0 13 0 1 15 12 15 1 10 9 13 1 9 2 13 15 15 12 1 0 13 2 7 15 13 9 13 3 2 16 13 9 7 2 1 15 2 3 9 0 2 16 13 9 2
8 15 3 13 13 7 9 9 2
17 3 2 1 9 13 2 13 15 3 0 0 2 7 3 0 13 2
14 15 0 0 9 13 2 0 9 13 2 9 0 13 2
42 16 3 2 1 9 0 2 15 13 0 1 9 2 0 3 9 0 3 13 2 7 15 1 9 2 7 0 1 9 0 2 13 4 2 7 3 15 1 0 9 13 2
19 15 3 9 0 1 0 9 9 9 13 13 2 7 1 15 0 15 13 2
26 15 3 9 1 3 1 0 13 2 15 9 15 3 0 13 2 1 9 2 7 1 9 1 9 13 2
12 7 1 0 13 13 13 9 3 13 9 13 2
16 16 3 3 13 12 10 9 0 16 13 2 3 1 13 4 2
29 3 13 1 15 9 13 15 13 0 9 13 9 2 7 3 13 15 1 9 13 2 7 1 0 7 1 9 9 2
7 15 3 13 9 15 9 2
13 13 4 3 1 9 13 9 16 9 7 9 15 2
20 9 7 2 16 13 0 0 9 2 3 2 1 12 7 15 2 9 13 0 2
8 13 3 15 1 9 1 9 2
19 0 3 13 9 2 15 13 9 0 2 16 13 9 2 15 13 9 9 2
2 3 2
8 15 9 0 13 0 9 13 2
11 3 13 1 9 7 9 13 15 1 9 2
17 0 7 13 15 15 13 15 1 9 2 16 15 13 15 1 9 2
21 15 3 13 15 1 9 13 15 1 9 2 15 7 13 1 9 13 15 1 15 2
15 15 7 1 9 13 2 3 0 13 15 15 13 1 15 2
13 9 3 0 13 4 13 9 16 4 1 9 13 2
9 3 3 13 4 1 9 15 13 2
2 0 2
9 10 9 1 10 15 13 13 0 2
16 9 7 2 1 13 9 2 16 13 4 2 13 9 9 0 2
11 3 2 13 1 15 1 9 2 13 0 2
10 13 7 13 0 0 1 9 0 9 2
18 3 3 13 9 9 16 9 4 0 13 1 9 13 2 16 9 13 2
2 0 2
14 16 9 4 13 1 9 2 13 13 3 4 9 13 2
10 7 3 15 13 0 2 7 1 9 2
20 16 7 0 2 10 7 0 13 1 9 2 13 3 9 1 9 13 1 9 2
12 9 3 2 15 1 15 13 2 13 15 0 2
5 15 13 13 0 2
11 3 2 9 0 9 9 13 16 9 0 2
10 1 9 7 0 15 13 0 7 0 2
7 0 3 0 1 9 0 2
18 16 7 0 9 4 9 13 2 0 3 9 1 15 9 13 9 13 2
20 9 7 0 3 13 1 9 16 13 15 13 2 16 13 1 9 0 7 0 2
7 9 3 3 12 9 13 2
14 3 3 1 9 10 9 13 9 13 16 13 15 13 2
11 7 10 13 9 0 9 2 13 9 13 2
13 1 9 3 13 16 9 13 15 9 1 9 13 2
4 15 13 9 2
15 7 16 1 15 9 3 13 13 15 0 2 16 13 4 2
30 7 16 0 2 7 15 13 1 9 2 1 13 1 9 2 3 13 13 0 15 15 13 1 9 2 7 15 9 13 2
2 3 2
17 1 15 0 13 10 9 2 9 13 13 9 2 7 3 1 0 2
15 9 7 13 1 9 16 9 1 9 2 16 1 13 4 2
17 3 3 13 9 1 9 13 1 9 9 2 7 3 1 9 9 2
28 16 7 13 16 15 13 9 0 2 3 13 9 7 13 1 9 13 2 1 0 9 2 2 15 13 13 0 2
16 16 15 15 0 13 1 0 2 13 9 2 16 9 7 0 2
19 16 3 13 9 7 13 1 9 0 1 9 13 2 13 9 9 9 13 2
17 7 3 1 15 13 9 13 3 13 9 1 15 2 7 1 9 2
2 3 2
21 10 15 15 13 9 15 1 9 9 2 13 13 0 9 2 15 13 15 9 9 2
17 9 7 0 7 0 2 1 15 13 9 13 2 13 15 9 9 2
8 3 3 13 13 13 0 9 2
25 0 13 3 16 2 1 0 9 2 0 13 3 7 13 3 2 7 0 3 15 2 3 15 13 2
23 16 7 13 16 7 1 9 7 1 9 9 13 2 7 0 9 2 2 15 13 3 13 2
10 15 3 13 1 9 0 13 16 13 2
10 9 7 13 13 9 9 16 9 13 2
24 7 0 1 0 15 13 16 1 13 9 13 9 15 15 0 13 2 7 13 1 9 0 9 2
8 3 3 13 9 13 16 13 2
19 9 7 15 1 15 9 13 13 2 1 13 2 1 15 2 9 10 13 2
30 7 13 13 16 9 1 0 9 13 1 0 0 13 1 9 2 16 13 1 0 2 16 9 3 3 13 1 0 9 2
8 3 3 13 13 1 9 13 2
16 13 3 16 9 2 16 13 1 9 2 3 13 9 0 9 2
2 3 2
34 10 9 13 1 9 12 9 1 3 3 13 2 13 9 0 2 16 13 1 15 2 13 13 2 13 1 9 9 15 3 1 13 13 2
21 9 7 0 13 2 1 15 13 9 9 2 3 13 9 1 9 9 13 13 13 2
18 1 3 1 15 9 13 9 7 9 13 3 13 2 13 16 13 0 2
13 7 3 9 9 3 13 1 9 2 7 1 9 2
11 15 13 13 0 2 1 13 16 1 0 2
36 16 7 3 13 16 3 1 9 2 7 1 0 9 9 9 13 2 7 1 0 9 2 2 15 3 3 13 13 2 16 9 1 9 4 13 2
10 15 3 9 13 1 13 9 10 9 2
32 3 7 8 12 2 1 0 13 13 2 13 9 16 13 0 2 7 3 1 10 2 13 9 10 15 13 2 7 13 3 0 2
19 16 3 9 13 1 9 13 2 13 13 16 15 9 13 13 13 9 15 2
20 3 13 7 1 9 0 9 13 9 1 9 9 13 2 7 3 1 0 13 2
12 3 3 1 0 9 13 4 16 9 9 13 2
2 3 2
15 3 13 1 9 0 9 1 0 9 15 15 13 9 13 2
11 9 7 1 9 9 13 9 0 7 0 2
32 3 3 13 13 9 0 9 2 1 13 0 9 2 9 13 15 13 2 1 15 1 9 15 13 3 13 2 16 1 13 13 2
28 15 7 9 13 2 1 13 9 0 1 9 4 13 2 13 16 9 0 9 9 13 13 2 7 1 15 9 2
25 3 1 9 15 13 13 2 7 1 9 9 9 0 7 0 0 15 13 2 3 15 9 2 13 2
7 7 15 9 13 3 13 2
12 9 3 9 9 13 2 7 1 15 13 0 2
15 16 3 13 9 7 9 13 15 0 2 3 13 9 9 2
4 15 13 0 2
6 13 3 13 1 9 2
7 3 1 15 0 9 13 2
33 7 3 13 8 13 9 3 13 9 1 9 2 1 3 8 12 13 2 1 9 9 2 13 9 10 15 13 2 7 13 3 0 2
2 3 2
9 1 0 3 13 9 16 1 9 2
25 16 3 1 9 9 13 15 13 4 2 16 9 9 13 2 1 15 13 15 9 2 1 9 13 2
7 0 3 13 16 9 13 2
22 15 13 0 9 2 1 15 13 2 8 12 2 16 10 1 9 2 9 7 9 13 2
9 3 7 7 15 13 0 0 9 2
30 13 3 8 12 1 9 7 9 2 16 2 1 3 13 4 7 15 0 7 0 13 2 13 4 2 16 0 13 0 2
27 3 3 2 16 15 9 13 2 15 15 9 13 2 1 3 15 1 15 9 13 4 2 16 13 8 12 2
22 13 7 1 2 1 1 9 9 13 2 0 1 9 9 13 2 15 3 3 13 13 2
11 7 3 2 15 13 2 1 15 13 13 2
2 3 2
13 0 13 13 16 9 0 7 13 9 2 7 3 2
41 13 7 0 1 15 15 13 2 16 13 9 2 16 15 13 9 15 2 3 13 9 1 0 15 13 1 9 15 2 16 0 13 15 9 13 7 15 13 1 9 2
24 7 3 2 16 3 13 0 0 9 9 1 13 2 3 13 1 9 15 9 0 7 0 9 2
4 15 0 13 2
26 3 1 9 13 1 15 9 2 1 15 9 1 9 13 2 1 15 1 13 0 9 7 9 9 13 2
45 16 3 9 0 1 13 9 13 2 9 7 15 13 1 0 1 0 9 13 2 16 9 13 9 0 7 9 2 13 13 9 9 7 9 2 3 4 9 0 1 0 9 9 13 2
13 9 7 3 13 1 9 0 2 16 1 13 13 2
9 3 3 4 13 9 1 9 0 2
34 16 7 9 0 3 13 9 1 13 2 7 1 15 13 1 9 4 13 2 13 13 16 2 16 9 13 2 10 9 9 13 1 15 2
22 15 7 0 13 2 13 9 2 15 13 9 9 0 13 1 9 9 2 9 9 13 2
15 3 9 13 2 1 15 9 13 2 0 10 9 9 13 2
18 13 3 13 16 2 16 9 13 2 1 13 13 2 9 13 9 13 2
53 15 3 0 13 2 15 9 9 13 13 16 15 2 15 13 2 13 13 1 15 15 1 9 13 2 9 13 2 16 2 1 15 3 13 15 15 0 13 2 9 13 15 15 0 4 13 2 1 15 9 15 13 2
12 1 15 3 13 16 13 3 13 15 16 13 2
16 3 3 1 15 9 1 9 13 16 13 9 9 13 9 9 2
20 15 7 9 9 13 15 1 16 10 9 13 2 7 3 15 1 15 13 13 2
9 3 3 13 13 9 7 9 0 2
13 7 3 9 3 13 9 0 2 7 15 9 0 2
5 15 13 13 0 2
2 3 2
15 0 9 9 15 13 15 1 15 9 13 13 1 10 9 2
15 7 1 10 0 9 13 7 13 9 13 13 1 9 9 2
13 3 9 9 0 13 15 9 7 9 1 9 0 2
9 9 3 9 13 13 1 9 9 2
8 1 15 3 9 13 13 9 2
5 15 13 13 9 2
20 3 3 1 15 16 13 9 2 9 13 13 2 7 3 15 13 16 9 13 2
2 3 2
34 16 15 9 0 1 15 15 1 9 13 13 2 3 13 9 16 1 0 9 2 15 15 13 2 7 13 1 10 15 9 7 0 13 2
35 3 7 13 13 2 13 9 1 15 15 13 0 9 2 13 9 1 9 2 7 3 3 3 9 0 9 1 15 1 15 13 2 13 13 2
20 1 15 3 0 13 16 1 9 0 2 1 15 15 13 2 13 9 1 0 2
7 3 3 0 13 9 13 2
2 3 2
31 16 3 13 9 0 9 9 16 9 2 15 13 9 1 10 1 9 16 1 9 2 16 15 13 0 2 13 15 1 10 2
15 3 13 7 1 10 15 9 1 9 2 7 0 1 9 2
13 13 3 16 9 9 13 15 0 2 3 7 9 2
24 15 7 3 13 0 15 2 13 1 15 15 13 0 2 16 3 1 0 1 9 13 10 0 2
12 3 3 9 9 13 1 15 16 1 9 13 2
2 3 2
23 1 9 3 13 1 12 2 12 9 13 13 0 12 9 2 16 9 9 2 7 9 0 2
21 9 3 1 13 12 9 2 13 15 12 0 9 2 15 1 15 7 0 9 13 2
26 15 7 13 13 15 1 15 13 10 1 9 13 2 16 1 9 13 10 9 2 15 13 1 15 0 2
7 15 3 13 15 16 9 2
17 0 3 9 10 13 9 2 7 15 15 13 1 15 9 16 3 2
20 1 15 9 13 0 9 9 2 16 3 13 3 13 7 13 2 7 15 3 2
26 15 3 0 9 9 10 0 13 2 9 7 1 15 2 16 1 9 13 9 3 0 16 0 1 9 2
2 3 2
14 15 15 1 9 1 15 13 2 3 13 9 1 9 2
10 7 15 9 9 1 15 1 0 13 2
25 16 3 15 15 9 13 2 3 13 13 16 15 13 0 9 2 16 7 0 13 15 13 1 9 2
10 3 7 15 9 9 13 9 1 9 2
5 0 3 0 15 2
13 3 3 0 13 9 9 16 9 13 16 9 13 2
2 3 2
20 16 10 9 13 9 15 13 2 13 13 16 15 9 1 9 9 0 9 13 2
8 15 3 13 13 13 9 9 2
19 16 3 9 9 13 0 2 13 0 9 0 13 7 13 1 15 9 9 2
35 7 3 13 13 9 13 9 0 2 16 0 9 0 9 13 2 7 13 13 2 16 9 13 13 2 16 15 13 3 15 2 3 15 9 2
17 15 7 13 13 16 13 9 13 9 2 7 3 9 3 13 0 2
21 16 3 13 0 9 3 3 13 2 3 15 0 13 16 1 9 1 0 13 13 2
25 3 3 4 15 0 13 2 16 1 9 13 2 16 2 16 4 1 15 13 2 3 13 15 13 2
18 15 7 13 0 2 16 2 9 13 13 2 12 0 9 13 3 13 2
16 3 7 0 13 9 1 9 2 13 9 9 1 9 1 9 2
5 15 7 13 0 2
7 3 3 9 1 9 13 2
13 16 7 13 0 12 9 0 9 13 2 3 13 2
13 9 3 0 3 13 9 1 3 2 7 9 0 2
6 3 7 9 9 13 2
9 9 7 1 9 13 1 9 0 2
9 13 3 9 9 1 15 0 13 2
10 3 7 3 16 15 9 13 9 9 2
17 13 4 3 1 16 13 9 0 2 7 16 15 15 9 9 13 2
25 13 3 16 1 9 1 0 9 15 9 13 2 9 7 9 9 13 2 15 9 15 1 13 4 2
15 16 3 13 0 9 2 0 13 16 13 0 9 15 13 2
6 3 3 12 0 13 2
2 3 2
9 13 4 1 9 13 9 16 9 2
18 9 7 13 13 0 9 13 2 1 15 13 1 3 16 9 7 9 2
7 0 3 9 0 9 13 2
8 3 3 12 9 0 9 13 2
2 0 2
8 9 9 13 13 10 0 13 2
8 3 3 15 9 13 15 0 2
19 9 7 2 16 3 13 9 9 2 3 3 13 13 16 3 13 9 15 2
9 13 3 1 0 13 9 7 9 2
9 13 3 1 9 9 13 9 9 2
2 3 2
15 1 15 15 13 7 13 2 0 13 1 9 13 15 9 2
30 1 3 9 7 9 13 9 1 9 2 1 15 15 13 7 13 3 13 9 15 2 16 13 1 15 15 1 9 13 2
17 7 16 12 9 0 9 13 13 0 2 13 15 9 9 1 9 2
14 15 9 1 9 13 2 15 13 9 13 9 9 13 2
30 13 3 7 15 15 2 16 2 1 9 9 13 9 2 16 7 9 2 13 16 15 13 12 9 15 13 9 9 12 2
10 3 3 13 0 12 9 0 9 13 2
11 1 15 3 13 16 7 9 13 1 9 2
8 15 7 9 0 9 9 13 2
5 13 3 1 9 2
6 15 13 0 9 15 2
20 16 3 15 3 9 9 13 2 3 7 3 10 13 2 7 12 0 9 13 2
9 15 3 1 9 1 8 9 13 2
20 9 9 13 3 13 1 9 1 10 0 9 2 7 3 13 2 16 9 13 2
4 9 9 13 2
18 9 7 15 13 9 1 0 13 2 7 3 9 13 2 0 13 13 2
38 15 3 0 13 2 9 13 9 16 13 3 2 13 13 2 7 13 16 9 7 9 9 3 15 13 1 15 15 13 2 7 1 15 15 13 7 13 2
9 3 7 1 13 9 9 3 13 2
23 3 3 1 15 16 9 13 9 16 13 3 2 13 13 16 3 13 2 7 16 3 13 2
2 3 2
14 1 9 3 13 15 1 15 13 9 2 16 13 9 2
24 16 3 9 13 9 16 13 3 2 3 3 13 13 16 9 13 3 2 16 16 15 9 13 2
23 16 7 13 16 15 9 1 0 13 2 4 13 15 15 13 13 2 3 15 13 1 0 2
23 15 0 0 13 2 1 9 9 2 15 13 9 2 13 13 16 13 9 9 13 13 0 2
9 12 9 2 3 1 15 15 13 2
9 15 9 2 3 1 15 15 13 2
23 7 16 3 9 13 13 0 3 1 15 15 13 2 13 9 9 15 13 2 3 7 13 2
18 16 7 9 13 13 0 3 1 15 15 13 2 13 13 9 13 0 2
12 3 7 9 13 3 13 0 2 7 0 9 2
22 1 13 3 13 9 0 15 9 10 13 9 2 1 0 15 13 1 9 1 9 13 2
18 3 3 13 13 16 9 13 0 2 7 16 9 13 13 1 15 0 2
14 13 3 1 0 9 2 16 1 9 0 0 10 9 2
20 1 15 7 0 13 9 2 3 16 9 1 9 2 7 16 9 1 0 9 2
9 3 0 13 9 9 7 9 15 2
21 1 9 7 9 13 13 1 9 9 2 16 7 1 9 9 13 13 1 9 13 2
14 15 3 13 13 1 9 0 2 13 13 0 0 9 2
15 3 13 13 1 9 9 0 9 9 2 3 7 15 9 2
23 16 0 3 3 13 13 1 9 9 2 13 1 15 15 1 13 4 1 1 9 9 13 2
13 15 3 0 13 2 1 9 0 2 9 3 13 2
23 0 3 9 13 3 1 9 2 3 7 3 1 9 2 1 0 0 0 9 13 13 9 2
17 9 7 0 3 13 0 1 9 2 7 0 9 2 16 13 4 2
11 3 3 13 9 0 16 9 1 0 13 2
11 1 15 3 13 9 1 15 15 0 13 2
22 3 3 13 2 8 12 2 16 9 13 9 10 2 7 16 13 1 10 9 15 13 2
38 16 3 9 7 9 9 1 9 13 7 3 1 9 2 3 9 9 13 13 1 9 1 0 9 13 2 3 7 1 0 9 2 15 0 1 9 13 2
26 7 3 2 1 10 9 0 13 12 9 16 7 10 9 2 3 13 13 9 16 9 3 0 9 13 2
15 13 7 13 16 1 9 3 13 13 16 9 0 13 0 2
13 15 3 13 13 1 15 15 1 10 9 3 13 2
6 13 7 15 13 0 2
16 15 3 13 13 1 15 15 3 13 2 3 16 3 3 13 2
53 3 7 1 12 8 2 1 9 0 1 9 15 9 13 2 3 13 16 15 9 13 1 9 2 15 3 9 1 9 13 2 7 3 13 13 9 1 15 13 16 15 15 1 9 13 2 7 13 16 13 1 9 2
8 16 9 3 13 1 9 9 2
11 1 15 3 13 9 3 13 1 9 9 2
16 13 4 3 1 0 9 13 0 2 7 15 15 1 0 13 2
12 9 7 0 3 13 1 9 2 16 13 4 2
9 3 3 9 13 13 1 9 0 2
2 0 2
11 13 4 1 16 9 15 9 9 13 13 2
11 9 7 0 13 9 9 2 16 13 4 2
7 3 3 13 1 9 0 2
2 3 2
17 10 15 1 15 13 15 2 13 1 9 1 15 15 13 1 15 2
20 9 7 9 3 13 1 9 1 15 2 1 13 0 9 2 16 1 13 4 2
14 0 13 3 16 1 9 9 13 9 2 7 15 15 2
2 3 2
10 15 1 15 13 15 2 15 9 13 2
11 9 7 13 3 0 2 16 1 13 4 2
10 0 13 3 16 1 15 15 13 13 2
2 0 2
13 1 9 0 13 9 1 9 7 9 7 15 13 2
13 9 7 13 3 0 2 7 1 15 7 1 9 2
9 3 3 9 13 13 1 9 0 2
2 3 2
15 1 13 4 16 9 13 9 0 2 1 15 15 9 13 2
10 1 9 7 0 13 7 9 7 9 2
24 13 3 1 15 9 0 2 15 13 9 1 10 0 2 7 9 13 2 16 1 1 13 13 2
9 3 13 3 9 0 1 9 0 2
2 3 2
20 1 9 0 13 3 0 2 3 13 15 9 15 13 9 16 13 15 9 15 2
14 9 7 0 0 13 13 16 12 2 16 1 13 4 2
13 13 3 16 10 9 13 3 9 12 3 1 9 2
6 7 15 1 13 4 2
8 3 13 3 9 1 9 0 2
9 13 7 15 9 1 0 9 13 2
8 15 3 13 15 9 0 13 2
30 3 0 9 9 13 13 2 7 15 13 9 2 7 9 2 7 15 15 9 13 2 7 1 9 15 9 9 13 13 2
19 3 10 15 15 13 9 2 9 13 2 16 13 1 9 1 12 1 9 2
9 7 3 13 9 13 1 9 0 2
28 7 1 15 9 13 9 9 2 15 13 9 13 15 9 0 1 0 9 13 2 15 15 9 0 9 13 13 2
36 15 7 9 1 13 4 2 7 1 15 16 13 4 9 3 13 9 2 7 1 15 16 13 4 9 3 0 9 3 13 2 7 15 0 9 2
24 15 0 13 9 10 9 13 12 2 7 13 3 2 7 13 7 0 3 2 16 1 13 4 2
23 7 16 15 9 13 0 9 13 13 2 13 9 10 2 3 9 15 13 2 13 0 9 2
24 3 7 1 15 10 9 0 9 9 2 13 9 13 13 2 13 4 13 16 9 13 13 9 2
11 15 7 9 1 9 9 10 1 13 4 2
14 13 7 7 1 15 9 9 10 1 9 15 9 13 2
22 13 3 2 15 0 13 0 9 2 15 9 1 9 9 13 13 16 9 2 1 9 2
9 3 13 13 9 1 9 0 13 2
15 7 3 1 9 1 15 9 13 13 16 9 9 13 0 2
23 1 15 3 13 13 15 8 12 2 16 13 4 2 13 9 1 9 7 9 10 2 13 2
15 13 9 9 1 9 9 2 7 13 1 9 15 9 9 2
12 1 15 15 13 13 16 9 13 1 9 0 2
18 15 3 1 9 15 13 2 15 9 15 1 15 13 2 1 15 13 2
18 7 3 13 9 13 16 15 0 1 9 1 9 1 15 13 13 4 2
25 7 9 13 3 13 9 13 15 9 0 2 1 1 13 9 0 13 2 15 1 9 13 3 13 2
13 3 15 9 3 13 0 15 0 9 16 15 9 2
12 15 3 9 13 1 13 1 9 9 9 13 2
20 3 7 9 13 9 9 1 9 1 9 1 15 9 13 2 3 1 9 9 2
30 1 15 7 1 9 9 9 13 13 2 16 2 1 1 15 9 9 13 0 9 9 13 2 1 15 9 0 9 13 2
23 3 3 9 13 1 9 9 9 13 2 16 9 9 9 13 2 3 15 1 10 9 13 2
31 3 7 15 0 13 1 9 15 2 3 13 13 4 9 2 9 1 9 15 13 2 3 7 15 10 9 9 1 15 13 2
8 16 9 0 3 13 1 9 2
18 1 13 7 13 13 16 9 0 3 13 1 9 2 3 1 9 13 2
18 15 3 9 9 3 13 13 1 9 2 7 15 9 1 9 13 13 2
16 3 3 9 13 9 16 7 13 2 1 15 13 16 13 9 2
19 1 0 0 2 15 9 9 13 1 9 2 15 9 3 13 1 9 9 2
17 9 7 9 0 7 0 3 13 13 1 9 2 16 1 13 13 2
15 9 7 9 0 3 13 1 9 0 2 16 1 13 4 2
15 3 9 0 7 0 1 9 9 13 2 3 7 9 0 2
8 7 9 9 1 9 9 13 2
15 3 9 0 7 0 13 13 1 9 9 2 3 7 0 2
2 3 2
16 16 9 0 1 9 9 13 13 2 15 3 13 13 16 0 2
46 12 9 2 16 13 13 1 9 9 2 3 1 9 13 1 9 13 2 16 9 13 1 9 2 16 13 1 9 0 2 15 13 13 2 1 15 13 9 12 1 9 7 0 1 9 2
15 13 7 9 9 13 2 1 15 9 13 13 9 13 9 2
27 15 9 2 16 13 1 9 13 9 0 9 0 2 16 3 9 0 13 13 1 9 9 2 7 3 9 2
9 0 7 15 13 0 2 0 9 2
32 0 16 2 1 9 0 13 9 9 7 0 9 2 15 0 0 13 9 13 0 9 1 9 2 1 15 13 0 15 9 13 2
27 3 3 13 13 16 13 9 1 9 13 2 16 7 3 9 0 9 1 9 13 2 16 13 1 9 0 2
31 0 16 2 1 9 2 15 13 0 7 0 9 9 0 2 3 13 15 9 9 9 2 3 13 13 1 9 1 9 9 2
5 3 7 9 0 2
5 0 3 13 0 2
15 9 3 0 15 13 1 9 2 13 1 9 9 13 9 2
11 3 3 15 13 13 9 15 13 1 9 2
16 7 10 9 15 13 9 1 9 9 2 13 9 1 9 13 2
24 9 3 9 13 15 1 9 1 9 2 7 3 13 1 9 9 9 2 15 13 1 13 9 2
32 3 2 16 1 15 3 13 9 9 0 2 9 9 3 13 16 1 15 15 13 13 9 2 7 3 13 1 9 1 9 13 2
30 16 3 9 0 13 1 9 1 9 0 15 13 1 9 2 13 16 9 10 13 13 1 9 2 16 9 15 9 0 2
6 15 0 1 13 4 2
12 15 3 9 9 0 13 1 9 1 9 9 2
2 0 2
17 10 9 15 13 1 9 1 9 9 2 13 9 13 1 9 9 2
12 15 3 13 9 13 2 1 9 1 9 13 2
10 9 7 0 3 13 13 1 9 9 2
26 3 3 1 13 4 16 15 9 0 13 15 13 9 2 1 13 15 9 1 9 2 16 1 13 4 2
11 3 3 9 0 13 1 9 1 9 9 2
12 7 3 2 7 1 9 9 15 13 1 9 2
2 3 2
8 15 9 0 13 1 10 9 2
20 7 9 0 13 15 9 9 2 1 13 9 1 10 9 13 2 15 13 13 2
9 15 3 9 0 13 13 9 0 2
15 7 10 9 9 15 13 1 9 2 13 1 15 9 0 2
16 13 3 9 0 13 0 9 2 9 2 9 2 7 9 9 2
15 3 3 13 13 1 13 9 0 1 9 15 13 1 9 2
2 3 2
20 0 13 13 15 0 9 7 1 9 9 13 2 7 3 1 15 9 0 13 2
13 7 9 0 13 15 0 9 2 16 1 13 4 2
23 3 3 13 13 16 13 1 9 9 2 7 16 13 1 9 1 9 0 15 13 1 9 2
12 7 3 15 9 1 9 9 9 0 13 13 2
2 3 2
18 16 9 15 13 9 16 15 13 2 9 15 13 9 16 15 13 13 2
21 9 7 9 3 13 9 16 9 0 13 13 2 1 13 0 2 16 1 13 4 2
11 7 3 9 9 13 9 16 9 13 13 2
9 7 9 9 13 0 9 9 9 2
11 3 13 3 9 9 9 9 9 1 9 2
22 1 15 7 13 9 0 7 0 15 2 15 13 9 1 9 13 2 16 1 9 9 2
11 16 9 0 13 1 9 1 9 1 9 2
18 1 15 7 15 13 4 2 13 13 16 0 9 9 0 13 1 9 2
17 10 3 15 1 9 13 7 13 1 15 7 1 9 2 7 13 2
22 9 7 0 3 13 1 15 2 1 3 13 13 1 9 7 9 2 16 1 13 4 2
5 7 13 1 9 2
22 1 3 13 9 9 2 13 1 9 9 2 15 13 1 9 0 9 2 15 13 4 2
31 1 3 9 0 1 0 13 13 2 3 3 13 0 2 7 13 9 2 16 1 13 4 2 13 16 13 1 9 1 9 2
10 13 4 7 1 16 0 9 13 13 2
9 0 3 15 9 0 1 9 13 2
2 0 2
19 10 15 15 9 3 13 10 9 2 13 10 9 9 2 16 1 13 4 2
8 9 7 0 3 13 10 9 2
11 15 3 0 9 13 2 16 1 13 4 2
7 13 3 9 0 10 9 2
12 7 15 1 15 13 9 2 1 15 3 13 2
29 15 0 3 13 9 1 15 2 7 0 1 15 2 3 1 15 13 2 7 15 13 2 16 9 9 13 9 13 2
27 9 7 0 15 13 0 1 15 9 2 16 13 1 10 9 0 2 7 9 15 13 15 0 2 9 13 2
20 9 3 1 15 13 10 13 2 1 9 15 9 2 15 13 1 9 9 13 2
20 7 2 1 9 0 3 13 9 9 10 2 3 13 13 1 15 16 1 9 2
7 13 3 16 1 15 13 2
5 7 3 2 13 2
21 1 3 9 13 9 0 9 2 16 1 13 4 2 13 16 1 0 9 0 13 2
2 3 2
18 15 15 13 12 9 2 13 15 9 13 1 9 2 16 1 13 4 2
21 9 7 13 1 9 9 0 2 15 3 13 15 13 13 1 9 16 1 9 9 2
11 9 3 0 13 1 9 1 9 1 9 2
2 3 2
26 15 13 1 9 1 15 9 2 13 1 15 7 15 15 13 9 13 1 15 9 2 7 15 9 0 2
37 9 7 3 13 3 13 1 9 16 13 15 15 15 13 9 13 2 16 13 1 9 13 1 9 7 9 2 15 13 1 15 16 13 9 1 9 2
23 3 3 13 9 15 1 15 15 13 15 9 13 2 1 13 9 0 2 16 1 13 4 2
20 13 3 16 3 13 1 9 1 15 9 16 1 15 16 13 1 15 9 0 2
11 15 7 9 13 0 9 0 7 0 9 2
20 0 3 9 13 1 15 16 13 9 10 9 1 9 13 2 15 13 9 13 2
18 9 3 3 13 13 1 9 16 1 0 7 0 9 2 15 13 9 2
2 3 2
6 9 9 13 9 15 2
18 3 3 9 9 13 1 1 0 9 13 2 7 1 9 7 15 9 2
28 9 7 9 0 7 0 9 15 13 16 1 9 7 9 13 15 9 9 7 13 1 0 9 2 15 9 13 2
9 3 1 15 13 0 10 9 9 2
10 15 3 13 13 0 9 2 8 12 2
58 1 3 2 1 9 15 9 13 2 15 9 15 9 13 2 16 1 13 2 13 9 0 9 13 2 7 0 1 15 2 1 9 13 2 9 15 1 9 13 13 2 13 2 13 9 9 1 9 9 2 7 13 1 9 15 9 9 2
12 1 15 7 13 9 13 9 1 9 4 13 2
10 9 1 13 16 9 0 13 1 9 2
9 13 7 15 15 13 13 13 13 2
33 1 3 9 13 9 16 13 9 0 2 9 7 9 0 9 7 15 9 13 2 13 16 9 0 9 13 15 9 1 9 15 9 2
13 15 7 13 12 9 2 15 9 13 13 1 9 2
20 9 3 0 9 2 16 7 15 9 2 1 9 15 13 1 9 1 9 13 2
17 13 7 15 1 9 9 0 7 0 1 9 2 16 1 13 4 2
11 13 3 16 3 9 0 1 9 9 13 2
2 3 2
17 16 13 9 1 9 1 9 9 2 0 9 13 9 9 16 9 2
16 7 2 1 13 9 7 3 9 2 13 9 0 7 3 0 2
19 15 3 0 3 13 0 1 9 0 9 13 2 16 7 1 10 9 13 2
41 15 7 8 9 0 13 1 9 16 13 0 2 16 7 15 9 13 1 9 16 13 9 0 2 16 9 13 16 9 0 13 13 15 1 9 2 15 1 13 4 2
14 13 3 16 9 9 0 13 1 9 15 13 1 9 2
2 3 2
13 9 2 1 13 9 9 2 13 9 1 10 9 2
16 7 1 15 15 13 12 1 9 2 13 12 9 7 12 9 2
20 16 3 13 0 9 2 7 1 13 0 9 2 13 16 13 13 0 1 9 2
13 13 3 12 9 12 9 13 1 9 9 7 9 2
13 13 7 16 9 13 1 9 9 15 13 1 9 2
18 3 7 1 15 13 9 2 15 13 15 9 2 7 3 1 9 13 2
2 0 2
14 9 13 15 0 1 9 1 9 15 13 1 9 13 2
22 10 7 9 0 13 15 0 1 9 1 15 16 13 9 13 2 1 15 13 15 9 2
18 9 3 0 2 1 15 13 9 9 2 13 1 9 15 13 1 9 2
2 3 2
4 0 3 13 2
8 15 13 9 9 2 13 9 2
19 7 2 16 9 13 1 9 2 15 13 9 9 9 15 3 1 9 13 2
5 3 9 9 13 2
5 15 15 9 13 2
16 13 7 1 9 15 9 9 13 2 15 9 1 15 15 13 2
4 13 7 3 2
12 1 9 7 9 13 12 2 15 13 9 12 2
25 16 3 9 13 0 16 9 2 7 9 0 16 9 2 15 13 0 7 0 15 2 15 13 0 2
7 3 3 13 9 7 9 2
8 7 9 13 13 1 9 9 2
10 3 7 1 9 9 9 1 9 13 2
2 3 2
19 0 13 13 9 9 15 3 15 9 1 9 13 2 7 0 15 15 9 2
35 16 3 9 9 1 9 13 2 9 0 9 9 13 2 15 12 13 9 12 2 3 9 2 15 9 2 3 9 7 0 9 2 0 13 2
5 15 13 13 9 2
12 1 12 3 7 15 9 13 9 7 9 9 2
8 13 7 9 9 13 9 9 2
4 3 7 9 2
2 3 2
68 1 10 15 13 1 9 2 10 9 9 13 3 13 9 1 9 2 16 9 3 13 2 16 13 1 9 2 7 1 15 15 9 2 16 9 7 9 7 9 7 9 7 9 9 13 1 0 9 2 7 3 13 9 7 13 2 15 9 0 2 1 9 2 3 13 15 0 2
7 13 7 9 13 9 9 2
18 1 9 3 9 9 13 9 0 2 3 7 1 15 0 9 9 13 2
2 0 2
14 15 15 13 15 9 7 9 2 13 13 15 9 9 2
15 7 1 9 9 15 9 9 7 9 2 7 15 9 13 2
17 1 3 16 9 7 9 9 13 2 7 9 9 3 7 3 13 2
23 3 0 13 9 9 0 2 7 3 9 9 0 2 7 3 2 9 13 2 9 9 0 2
8 3 15 13 9 9 7 9 2
9 7 9 9 9 13 1 9 9 2
6 3 7 9 9 9 2
2 3 2
24 15 13 15 2 13 1 9 15 15 13 2 16 9 15 13 9 2 13 15 9 1 9 9 2
14 13 7 9 9 2 7 15 9 2 13 0 9 13 2
14 15 13 3 9 9 15 13 1 9 9 1 15 13 2
7 9 3 13 1 9 9 2
17 3 7 9 13 2 1 12 1 9 2 16 9 13 0 9 9 2
10 15 7 3 13 16 9 13 1 9 2
10 3 9 1 9 15 13 1 9 13 2
8 13 3 9 0 1 9 9 2
8 7 3 1 9 9 9 13 2
2 3 2
6 15 13 16 1 9 2
5 9 7 13 0 2
5 15 13 1 12 2
8 0 3 2 16 1 13 13 2
18 0 2 16 1 9 13 9 0 7 9 9 2 15 13 9 13 9 2
27 0 2 16 9 9 9 13 2 16 1 15 9 13 2 1 9 2 15 13 0 2 3 13 13 1 13 2
6 13 3 9 1 9 2
8 7 3 1 9 9 9 13 2
2 0 2
33 16 9 3 13 1 9 2 16 13 4 2 7 13 13 1 9 9 2 13 16 0 13 9 2 7 3 15 13 9 1 0 13 2
14 7 16 15 13 0 2 13 0 16 9 13 1 9 2
16 15 3 13 1 15 2 13 15 0 2 16 9 13 1 9 2
5 15 7 13 0 2
7 3 3 9 13 1 9 2
6 9 3 3 0 13 2
11 13 3 13 16 9 3 1 9 9 13 2
4 9 9 13 2
22 1 0 0 13 9 9 2 13 13 15 1 13 9 7 9 9 0 2 7 0 9 2
39 0 3 13 13 0 13 9 15 13 16 9 9 15 13 1 9 1 0 9 2 3 13 1 15 9 2 7 9 9 2 1 15 13 2 7 1 9 9 2
21 16 3 15 13 0 2 3 9 3 13 9 2 1 10 9 1 9 7 9 13 2
31 9 3 9 3 13 1 9 0 0 2 7 1 0 9 2 1 15 0 1 3 13 13 13 13 2 15 13 0 13 15 2
8 15 3 13 2 13 15 9 2
15 3 13 1 13 13 9 9 0 2 1 9 15 0 13 2
9 7 0 13 15 0 1 9 9 2
17 3 13 7 13 13 15 1 9 15 1 15 13 2 3 1 15 2
21 3 2 1 9 13 13 1 0 9 2 7 3 13 2 3 13 15 13 9 9 2
26 7 3 13 13 16 1 9 1 15 9 13 9 1 10 9 13 2 15 3 9 3 13 1 9 9 2
18 3 2 1 9 13 9 16 9 2 3 13 16 9 15 13 0 9 2
7 13 7 9 9 9 0 2
17 3 13 3 1 9 9 1 9 9 9 2 7 0 9 7 9 2
45 3 7 9 13 2 1 12 1 9 2 16 9 7 9 3 13 9 9 13 16 13 9 2 3 9 13 2 1 3 15 15 9 13 9 2 13 9 9 13 2 3 3 13 9 2
31 13 3 2 16 1 9 9 13 1 9 2 16 9 9 13 0 1 9 2 16 13 1 9 0 2 16 1 12 13 12 2
16 9 3 2 16 3 1 4 13 9 13 2 3 13 9 0 2
12 10 7 9 0 13 9 0 2 3 15 13 2
20 16 15 0 9 9 0 13 2 3 13 1 9 13 2 7 1 3 9 15 2
10 3 3 9 9 13 1 15 9 9 2
9 10 7 9 13 13 1 9 0 2
12 7 3 3 13 0 16 15 1 9 0 13 2
19 7 16 0 13 16 13 1 9 9 2 1 15 16 1 13 9 13 13 2
18 7 16 13 16 1 10 9 1 15 9 3 13 2 3 0 9 13 2
9 7 3 13 13 2 15 15 13 2
43 16 1 9 9 1 9 3 13 9 9 2 7 9 2 1 9 9 2 3 15 9 9 2 15 13 9 0 2 16 3 13 2 13 0 9 9 1 9 2 7 3 9 2
26 7 16 9 9 0 13 9 16 9 0 2 0 9 13 1 9 9 13 2 15 13 9 13 9 0 2
15 3 2 9 3 13 7 13 2 15 13 16 13 9 0 2
41 0 7 2 9 9 13 2 15 9 13 0 2 3 3 1 9 9 9 2 7 1 9 0 9 2 1 15 13 9 13 9 1 0 13 2 1 9 1 9 9 2
22 1 3 15 9 2 13 16 15 9 15 9 3 13 9 0 3 2 7 3 9 0 2
11 7 3 15 9 0 0 3 7 3 13 2
17 7 0 13 16 3 3 2 7 0 13 9 0 1 9 1 9 2
12 7 0 16 9 13 9 0 2 16 7 9 2
7 15 10 13 0 1 9 2
13 13 3 3 0 9 2 3 16 9 0 13 0 2
14 15 3 0 15 9 0 13 13 15 13 0 1 9 2
21 15 0 13 1 0 2 15 13 0 2 1 13 1 9 2 16 13 1 12 0 2
26 9 7 9 0 2 1 13 4 1 9 13 1 9 13 1 9 13 2 1 9 13 0 1 9 9 2
35 16 3 15 13 0 15 9 0 13 2 15 0 15 13 1 15 2 13 3 0 9 0 2 1 9 13 16 9 0 2 9 13 2 13 2
14 15 13 0 2 16 1 13 4 2 7 9 0 13 2
70 3 3 15 9 15 1 9 13 7 13 0 2 13 9 2 7 1 9 9 13 9 2 7 2 1 15 13 16 1 0 9 1 9 15 13 9 0 2 16 15 0 2 13 9 9 16 13 1 9 9 9 2 15 13 9 16 0 13 2 3 1 9 9 13 2 3 16 9 13 2
11 3 3 13 13 15 2 7 13 1 9 2
9 7 15 13 13 1 0 9 9 2
10 3 3 13 13 9 9 9 9 0 2
41 3 16 9 0 3 13 10 9 16 13 9 0 7 0 2 15 15 13 2 1 13 13 3 9 2 7 16 9 0 3 13 1 9 15 9 2 7 1 9 9 2
19 7 3 13 13 9 0 2 15 9 13 13 9 13 2 15 3 3 13 2
21 3 3 9 1 9 9 13 1 9 13 2 7 13 1 13 9 7 0 9 9 2
4 0 7 0 2
13 1 15 3 13 9 1 9 2 7 0 1 9 2
17 1 0 7 7 0 9 2 13 16 3 13 15 9 9 15 13 2
46 13 3 16 9 9 2 0 3 1 0 7 0 9 2 3 13 1 9 13 2 7 1 9 0 13 1 9 15 2 7 13 1 9 9 0 9 2 15 9 13 13 0 13 1 9 2
16 15 3 9 0 15 13 1 9 13 1 9 9 1 1 9 2
7 9 3 13 3 13 15 2
18 3 0 13 9 9 2 3 9 2 7 3 3 16 13 1 0 9 2
48 16 3 9 0 9 3 13 1 9 2 15 16 15 15 13 9 0 9 0 2 1 9 3 9 15 2 13 13 9 9 2 1 0 9 0 2 1 0 9 9 7 0 9 1 15 9 13 2
10 7 3 13 0 9 7 9 15 13 2
27 7 13 9 16 15 0 13 7 3 3 13 2 16 0 3 13 9 13 2 7 13 16 1 9 1 9 2
16 7 3 3 13 16 13 2 7 16 1 15 1 0 13 13 2
26 7 13 0 16 15 9 9 3 13 0 2 7 13 0 9 0 2 16 15 3 13 1 9 7 9 2
25 3 3 13 15 9 0 2 7 15 9 2 7 0 9 0 13 0 0 2 16 13 1 12 9 2
34 3 3 15 9 13 0 7 3 13 1 9 9 2 3 13 13 0 9 0 2 15 9 1 9 0 13 2 7 1 13 0 9 0 2
32 7 3 1 9 9 7 9 1 15 13 9 9 2 13 0 9 7 9 0 2 7 1 13 9 2 16 9 12 13 9 15 2
35 9 3 0 2 15 0 13 2 1 9 13 9 9 2 13 2 7 13 9 9 2 15 13 0 7 0 3 2 7 3 9 13 9 9 2
17 15 7 13 2 13 9 0 1 0 13 2 16 13 13 9 9 2
10 15 3 13 2 0 13 13 1 9 2
34 15 3 0 13 2 13 9 0 15 9 9 1 9 7 1 0 13 2 1 15 16 9 1 15 0 13 2 2 13 15 0 3 13 2
24 16 3 9 0 1 9 7 0 13 1 9 9 2 13 3 9 2 16 7 15 15 13 9 2
35 16 3 9 15 13 9 2 1 15 9 9 13 1 15 16 13 0 2 3 9 0 9 1 9 0 0 9 13 1 15 16 13 3 0 2
23 9 3 1 0 13 15 15 13 0 3 2 7 1 13 7 9 7 15 9 1 9 13 2
14 3 13 16 3 1 9 9 13 2 7 1 9 13 2
42 9 7 0 1 9 2 1 13 1 0 9 9 0 2 1 15 13 16 15 9 9 4 1 9 7 9 1 9 13 2 7 1 9 9 13 2 7 1 15 9 13 2
30 0 3 9 9 1 9 13 3 13 1 9 0 2 1 15 13 9 9 2 7 1 9 0 2 1 15 13 9 9 2
12 3 3 13 13 9 9 2 7 0 9 9 2
20 15 0 0 13 2 13 0 13 9 16 9 2 3 13 0 9 1 9 13 2
35 3 9 0 1 15 9 13 2 3 13 2 7 15 13 9 15 13 3 0 7 0 2 1 15 13 9 7 9 3 2 16 1 13 13 2
22 15 0 0 13 2 0 9 9 3 13 1 12 13 2 13 13 1 0 9 3 13 2
13 16 3 13 4 1 3 2 13 15 13 12 9 2
17 3 9 13 0 13 1 9 9 0 13 0 16 3 15 9 0 2
20 3 13 16 9 15 1 9 13 1 0 9 2 3 0 13 0 9 16 9 2
49 13 7 3 16 9 0 9 13 1 15 1 13 1 15 3 13 9 9 2 16 9 0 1 9 9 13 2 1 15 3 13 13 9 9 2 15 13 15 9 2 16 13 13 1 15 13 7 13 2
44 1 3 10 9 9 0 13 1 9 16 9 1 0 7 0 9 2 15 13 1 12 7 15 13 15 13 9 2 9 9 1 15 9 13 2 7 3 1 15 15 13 9 9 2
22 9 3 9 13 3 7 9 9 3 0 9 7 0 2 7 3 9 9 3 9 0 2
19 7 9 9 13 9 0 2 15 9 9 13 3 13 2 7 13 1 15 2
6 3 13 9 1 0 2
25 3 3 9 15 0 1 9 13 2 16 9 9 15 0 13 1 0 9 2 1 15 9 9 13 2
12 9 0 9 13 1 9 9 2 15 13 9 2
10 3 3 9 9 0 13 2 7 9 2
14 9 7 15 13 1 9 9 15 13 0 2 3 0 2
13 3 3 13 9 16 9 15 9 13 0 9 13 2
12 15 0 0 13 2 13 16 3 1 9 13 2
25 16 3 13 16 9 9 13 0 16 9 13 2 7 1 13 2 3 13 16 15 9 13 0 15 2
11 3 3 9 13 10 9 2 7 10 9 2
10 13 7 16 15 9 15 13 15 0 2
5 15 3 13 9 2
7 3 9 9 13 0 9 2
26 9 13 1 16 13 1 9 1 9 2 3 1 16 9 13 1 9 9 2 3 3 13 3 1 9 2
24 9 3 0 2 1 15 13 1 9 1 9 2 3 1 3 13 9 2 13 0 9 16 9 2
11 3 7 3 13 0 9 2 7 9 3 2
24 1 0 13 0 9 2 3 1 9 0 9 2 3 13 0 7 0 9 2 7 3 1 15 2
29 7 3 13 2 16 9 1 9 9 3 13 7 0 9 2 16 13 0 9 3 9 7 9 2 16 0 9 13 2
11 9 3 9 15 13 2 7 9 7 9 2
16 16 9 9 13 1 15 13 9 9 0 2 9 7 0 13 2
17 7 3 13 16 9 9 9 13 0 2 1 13 15 1 15 13 2
25 13 13 3 1 9 9 13 10 15 15 9 0 3 13 2 16 9 2 9 2 9 2 7 0 2
24 1 15 13 3 13 16 15 9 15 15 9 0 13 2 1 9 9 13 2 16 0 9 13 2
42 16 7 9 9 13 13 1 9 9 0 16 13 9 9 2 3 13 9 0 7 9 15 9 13 2 16 0 9 13 2 7 13 16 9 9 9 13 0 1 9 9 2
27 15 7 0 13 2 9 9 13 2 7 1 15 9 15 9 0 13 2 9 3 13 0 2 9 7 0 2
20 16 3 13 1 9 13 2 13 0 15 13 2 0 7 16 13 1 9 13 2
24 3 3 9 9 13 13 9 3 1 0 7 0 9 2 7 9 9 13 2 16 1 13 4 2
9 0 3 7 10 9 10 9 13 2
15 3 3 15 9 13 1 9 13 2 7 1 9 9 13 2
23 15 7 0 13 1 9 9 1 9 9 2 2 13 3 1 13 3 13 0 16 1 9 2
10 3 7 9 9 3 13 2 7 9 2
24 1 9 7 9 13 9 0 7 0 1 9 9 2 15 3 13 2 7 13 2 9 0 13 2
22 7 3 2 16 9 9 9 13 0 2 13 16 9 13 1 9 2 16 0 9 13 2
7 13 3 15 1 15 0 2
17 12 9 1 15 9 2 7 9 7 15 3 13 15 13 1 9 2
20 7 3 13 0 15 1 15 13 2 16 9 13 1 9 2 7 9 1 9 2
13 15 9 13 15 1 15 2 3 2 1 9 15 2
14 7 3 15 13 1 15 2 13 0 9 7 9 0 2
15 15 7 9 9 13 1 9 2 16 7 10 9 1 9 2
24 1 7 13 16 1 9 7 9 3 13 12 1 9 2 16 13 15 13 9 3 13 9 9 2
12 16 15 15 9 16 0 13 9 0 16 9 2
29 16 0 13 4 9 15 0 9 13 16 9 2 3 9 0 2 13 13 3 15 15 9 15 9 0 16 9 13 2
30 7 3 1 9 0 2 16 4 13 9 0 2 0 2 4 13 15 1 15 9 13 2 7 16 9 15 1 0 13 2
9 3 0 9 1 9 0 13 13 2
16 16 7 15 9 0 9 0 13 16 9 16 0 2 0 13 2
14 16 3 15 9 13 2 7 13 9 13 2 7 0 2
7 3 7 13 13 9 13 2
18 16 13 15 9 0 13 0 9 2 1 10 9 2 1 10 9 13 2
15 1 13 3 9 13 0 9 13 3 3 1 9 9 13 2
21 7 3 2 16 13 9 0 2 3 9 0 2 16 13 9 13 2 13 13 13 2
20 3 3 13 16 9 9 7 9 9 2 15 9 9 13 2 13 9 0 9 2
9 9 7 0 0 13 9 9 0 2
20 13 3 2 16 9 0 13 15 9 13 2 16 15 13 15 9 1 9 0 2
15 9 3 15 13 15 9 1 9 0 2 16 13 9 0 2
12 3 3 13 9 1 9 1 15 9 7 9 2
22 0 7 7 9 0 2 13 9 7 9 7 9 7 9 2 13 13 9 0 16 9 2
11 15 3 15 9 13 0 1 15 7 9 2
22 15 3 9 7 9 13 9 9 7 15 9 2 16 15 9 13 2 7 0 1 15 2
7 0 7 9 0 9 13 2
28 16 3 15 9 15 13 9 4 13 9 0 2 13 9 2 15 9 7 10 9 15 2 15 9 2 4 13 2
6 15 7 0 13 0 2
13 3 15 9 9 13 1 9 9 7 15 0 9 2
16 3 3 15 9 9 2 7 0 9 2 9 0 13 16 9 2
2 3 2
35 16 15 0 9 13 15 9 0 16 9 2 7 13 9 3 2 7 13 15 9 2 3 15 13 1 9 0 7 0 2 16 13 1 9 2
10 16 7 13 9 3 2 3 13 9 2
11 10 3 9 9 13 15 0 9 1 9 2
16 9 7 3 13 15 9 1 9 13 2 16 1 16 13 9 2
19 13 3 15 3 13 9 15 1 9 9 13 2 7 15 9 2 7 13 2
17 9 3 9 13 1 13 0 2 3 1 13 2 7 3 13 15 2
12 3 3 13 16 2 1 15 9 2 4 13 2
33 16 7 13 9 0 15 13 13 9 7 9 15 2 15 9 9 2 1 9 15 13 9 15 9 2 13 1 9 9 13 9 9 2
5 15 13 9 15 2
14 3 3 9 0 13 13 16 9 15 9 7 9 15 2
2 0 2
24 3 15 9 13 0 9 0 2 3 13 0 2 3 3 1 9 13 2 7 0 1 9 0 2
20 9 7 15 13 0 9 0 16 9 13 2 1 7 15 13 13 9 9 0 2
11 13 3 9 9 0 1 10 9 9 13 2
24 1 3 0 9 13 0 9 2 0 13 16 0 9 2 15 13 9 0 2 4 13 9 9 2
2 3 2
34 16 9 9 2 7 15 9 15 2 4 13 0 9 2 15 13 9 0 2 13 16 2 3 15 9 13 0 9 2 13 0 1 9 2
9 15 7 3 13 2 7 3 0 2
28 3 9 0 13 1 9 16 9 2 1 3 13 0 9 2 7 0 2 15 13 3 0 2 15 13 1 9 2
15 3 3 9 0 13 15 9 2 7 9 15 2 16 9 2
2 3 2
9 10 13 0 9 1 9 9 13 2
15 3 9 7 9 13 1 13 0 7 0 2 0 7 0 2
10 1 9 7 9 0 13 9 15 9 2
10 3 3 13 0 16 1 15 13 9 2
11 0 3 13 16 9 0 13 15 16 9 2
2 0 2
17 9 16 1 15 13 0 2 3 0 9 13 0 2 3 9 13 2
20 16 3 15 9 9 13 15 13 9 13 2 0 13 16 13 15 9 0 13 2
31 15 3 13 9 9 2 15 13 0 0 7 0 7 0 9 2 1 16 7 2 3 0 1 9 1 9 2 10 9 13 2
21 15 7 9 0 13 13 9 0 2 1 13 9 9 3 13 9 9 2 7 9 2
8 15 13 0 1 13 7 13 2
12 3 3 13 0 15 9 9 4 13 9 0 2
2 3 2
10 10 9 13 15 9 1 9 0 13 2
12 3 9 0 2 16 3 4 13 2 13 0 2
5 9 9 9 0 2
7 9 7 9 9 7 9 2
14 9 7 9 9 7 9 2 15 13 15 9 1 9 2
17 7 1 9 3 13 15 9 15 13 1 9 2 7 0 9 0 2
6 3 13 3 9 13 2
24 16 7 13 16 9 0 2 16 3 13 9 9 7 9 15 16 9 2 13 3 15 16 9 2
10 0 3 2 1 9 15 13 0 13 2
27 1 3 9 9 3 13 1 15 0 2 3 13 15 9 15 13 9 0 13 2 1 15 15 9 0 13 2
2 3 2
26 16 15 9 0 13 15 9 0 16 9 0 0 2 13 9 9 15 9 13 1 9 0 15 0 13 2
12 3 15 9 0 9 3 13 1 13 0 0 2
24 0 7 13 13 16 9 15 9 0 3 13 1 13 15 13 9 15 9 2 7 15 9 13 2
23 3 13 3 13 16 15 9 0 13 15 9 0 0 16 9 2 16 15 3 13 16 9 2
2 3 2
13 9 9 0 13 1 15 9 13 16 1 9 0 2
13 0 3 13 1 3 9 0 9 0 9 0 13 2
43 1 15 7 13 9 9 2 7 15 0 2 15 13 0 13 9 9 0 2 9 0 2 9 0 2 9 0 2 7 15 0 13 9 13 13 2 3 7 15 9 0 13 2
20 13 3 9 13 9 7 9 13 9 0 15 13 2 1 9 0 7 9 9 2
9 16 13 15 9 0 9 3 13 2
14 1 13 7 13 13 13 15 9 0 9 3 3 13 2
16 13 4 3 1 2 9 13 2 9 9 2 3 0 2 13 2
28 7 16 3 9 9 15 13 2 13 12 10 2 16 15 13 2 1 9 13 15 13 1 10 9 1 9 13 2
13 7 3 13 13 2 16 9 0 15 1 9 13 2
31 16 7 0 9 0 13 2 9 13 2 13 15 9 0 1 9 13 2 3 1 13 4 16 9 3 13 1 9 1 9 2
16 13 7 9 13 1 9 13 1 9 2 1 0 13 9 9 2
16 15 7 15 13 1 9 2 13 0 13 15 15 13 1 15 2
19 13 3 15 9 0 2 9 1 9 0 2 15 1 15 13 1 9 13 2
2 0 2
13 10 15 13 1 9 9 2 13 1 9 9 13 2
28 13 7 15 15 13 1 9 9 2 3 7 1 9 9 2 16 0 13 1 9 9 2 3 7 1 9 9 2
21 15 7 13 1 9 9 2 3 7 1 9 9 2 3 13 0 10 9 9 13 2
7 0 3 9 13 0 9 2
24 9 7 0 1 10 9 13 16 13 1 15 13 2 1 13 1 15 9 2 16 0 4 13 2
13 1 9 7 9 1 15 13 3 13 16 15 13 2
28 3 13 3 1 9 9 0 1 10 9 16 13 9 13 2 16 13 15 1 9 15 0 9 2 15 13 9 2
9 13 3 15 9 0 9 3 13 2
2 3 2
12 9 0 1 10 9 13 9 9 1 15 0 2
7 9 7 0 13 0 0 2
13 13 7 15 1 15 9 10 2 15 13 9 0 2
31 13 3 16 2 16 9 9 1 9 0 13 0 1 9 9 2 3 9 0 2 15 13 9 2 13 9 1 9 9 0 2
15 13 3 15 9 0 3 13 9 2 0 1 9 9 9 2
2 3 2
22 16 13 15 0 1 15 9 2 13 1 15 2 1 9 9 2 15 1 9 15 9 2
7 9 3 9 0 13 0 2
17 9 7 15 13 1 9 2 13 9 0 2 16 3 13 9 0 2
17 13 3 15 9 15 13 9 0 1 15 0 2 7 9 0 13 2
13 10 7 9 1 15 0 1 9 2 13 9 0 2
12 9 3 9 13 9 0 2 16 1 13 13 2
9 13 3 15 9 0 9 3 13 2
6 10 3 9 9 13 2
2 0 2
14 9 13 13 1 9 2 16 9 1 9 13 3 13 2
12 9 3 15 9 0 13 9 2 9 7 9 2
8 7 15 9 0 13 1 9 2
11 13 3 13 15 1 9 9 3 1 9 2
9 10 7 9 0 1 9 9 13 2
6 15 3 13 0 0 2
9 1 0 3 3 13 13 7 13 2
36 13 3 15 9 1 9 13 2 1 0 9 2 15 9 13 2 15 3 13 1 9 2 16 1 13 4 2 7 1 9 2 15 13 9 13 2
2 3 2
35 16 1 15 12 13 15 9 2 7 15 15 13 1 15 15 13 0 9 2 7 15 2 15 13 3 9 7 0 10 13 2 1 15 13 2
16 13 7 15 9 13 1 9 0 7 9 2 16 1 13 13 2
13 9 7 13 1 15 2 16 13 1 10 9 0 2
10 0 3 0 13 9 0 9 3 13 2
2 3 2
17 9 9 13 13 13 10 9 2 16 9 13 9 7 9 9 13 2
8 7 13 13 0 9 9 0 2
11 13 3 9 0 15 13 15 13 13 9 2
22 13 7 2 1 13 9 1 9 0 3 13 2 3 13 9 16 16 0 13 1 0 2
7 15 7 13 0 9 13 2
15 9 3 9 13 13 16 13 15 15 13 1 9 10 0 2
24 16 7 3 13 16 15 15 3 13 1 15 0 2 7 13 0 1 9 2 13 0 9 13 2
54 16 3 1 10 0 13 13 9 15 1 9 15 2 13 16 1 9 0 2 15 13 13 1 9 2 13 15 0 9 13 15 15 13 1 15 0 2 3 13 9 1 0 2 7 1 15 3 1 9 1 10 9 13 2
2 3 2
7 9 13 3 1 12 0 2
32 9 0 2 0 7 2 3 1 15 13 2 0 2 13 13 1 9 15 3 13 7 1 15 7 1 9 2 16 1 13 4 2
9 0 3 9 13 1 0 9 13 2
36 9 7 9 13 0 2 0 2 7 2 3 1 15 13 2 0 13 2 7 1 0 9 2 13 0 15 9 1 9 2 16 1 9 9 13 2
15 13 3 13 0 9 15 3 13 7 1 15 7 1 9 2
12 15 7 9 13 16 13 2 16 1 13 4 2
18 9 7 0 13 9 2 13 1 9 1 9 9 2 16 13 1 9 2
14 13 3 13 0 9 15 7 13 9 7 13 9 13 2
13 9 7 0 13 1 15 9 2 16 1 13 4 2
9 13 3 0 9 0 9 3 13 2
24 15 7 13 9 9 2 12 8 1 8 8 2 13 1 9 16 2 16 0 2 7 0 13 2
13 1 15 7 13 9 9 2 15 13 9 3 13 2
12 7 9 0 0 2 15 13 10 9 0 13 2
18 9 3 9 15 13 16 15 9 2 1 9 0 2 1 9 13 13 2
17 7 10 15 13 10 9 2 0 7 0 2 13 9 0 15 13 2
5 1 9 9 13 2
31 13 13 7 16 9 13 13 3 0 13 15 9 0 1 9 2 7 16 13 15 9 15 13 9 13 1 9 2 7 0 2
36 13 3 16 3 13 15 9 1 9 15 1 15 13 3 13 2 1 15 16 10 9 15 13 1 9 2 13 1 9 15 9 2 15 0 13 2
13 9 3 13 9 2 9 7 13 13 1 9 13 2
55 3 13 16 3 13 15 9 13 1 15 3 13 15 9 1 9 2 16 2 1 9 0 13 1 9 13 16 1 9 2 16 13 15 9 13 16 15 15 13 2 13 15 9 1 15 13 16 1 9 2 15 13 9 0 2
42 3 1 15 13 16 3 13 0 9 13 16 9 13 2 7 15 13 13 2 1 9 2 3 1 3 13 0 9 0 15 9 2 16 3 3 13 13 0 9 15 0 2
7 15 7 9 3 13 9 2
25 1 15 3 15 13 1 9 2 13 9 1 9 2 16 15 13 1 12 9 2 3 7 1 0 2
28 3 2 16 9 0 13 1 9 13 16 1 9 2 16 15 13 2 3 13 13 0 9 9 13 1 9 9 2
49 13 3 13 16 13 15 9 13 9 9 16 15 15 13 0 9 9 0 2 16 2 16 9 0 13 1 9 15 1 15 13 2 15 13 13 15 9 15 1 9 3 3 13 0 2 7 13 13 2
15 7 3 15 9 15 9 3 13 3 0 2 7 16 0 2
3 13 3 2
10 3 9 7 9 0 0 13 15 13 2
6 0 3 13 0 13 2
17 13 3 13 16 13 0 0 9 0 1 9 13 16 13 9 0 2
11 9 3 0 1 10 9 13 10 9 0 2
14 13 3 13 9 1 13 9 1 9 15 1 0 9 2
27 13 7 15 0 9 13 1 0 9 1 10 9 9 3 2 15 3 9 13 16 9 2 16 1 13 13 2
41 7 16 9 9 0 1 10 9 15 1 9 9 13 2 16 1 13 4 2 13 9 9 13 9 2 15 16 3 13 9 16 9 2 13 3 0 9 15 9 13 2
23 0 7 9 9 0 3 13 1 13 2 1 13 13 13 1 0 15 9 2 15 13 13 2
21 13 3 7 15 9 9 9 0 2 15 3 13 0 9 15 9 2 7 0 9 2
2 0 2
28 16 9 1 9 13 1 10 9 0 2 3 9 1 9 13 1 9 9 2 16 13 1 15 15 13 1 9 2
42 16 3 9 1 9 13 13 0 9 10 9 0 2 3 9 1 9 13 13 0 7 13 1 9 9 2 16 3 3 13 9 0 16 13 13 1 9 9 1 9 13 2
35 13 3 0 9 9 2 15 1 9 13 2 16 1 15 9 9 13 13 2 15 9 13 15 13 0 1 9 9 2 7 0 1 9 0 2
10 7 1 3 9 0 13 13 15 0 2
13 9 3 0 13 9 9 16 13 9 15 1 9 2
23 3 13 16 0 13 9 9 0 16 0 2 7 1 9 0 0 13 9 9 13 16 13 2
15 13 7 9 0 9 13 1 9 0 9 15 13 15 0 2
16 13 3 15 9 0 1 15 15 13 0 7 0 9 13 9 2
2 3 2
18 9 0 13 13 16 15 15 13 1 9 0 2 13 9 7 9 0 2
7 0 3 13 13 1 0 2
15 3 13 16 0 2 3 1 15 13 2 13 3 0 13 2
30 7 3 13 16 9 0 2 3 0 2 1 3 13 0 2 3 0 2 16 3 15 3 13 0 9 1 9 1 15 2
26 16 7 0 9 0 13 0 2 16 0 0 2 3 9 0 10 9 2 16 0 7 0 0 7 0 2
12 13 3 1 9 0 9 13 10 9 0 9 2
7 3 3 13 9 0 9 2
2 3 2
12 9 9 0 3 13 1 9 2 7 1 9 2
19 9 7 15 13 1 9 2 13 9 13 7 0 16 9 15 13 1 9 2
9 3 9 1 9 13 1 9 9 2
23 3 13 3 13 0 9 9 15 13 1 9 2 15 13 9 13 2 16 13 9 0 9 2
17 3 7 1 15 13 16 9 13 13 9 15 0 2 16 0 13 2
62 1 3 3 13 1 13 9 9 13 16 1 0 2 13 15 9 13 15 9 1 15 2 7 3 9 15 2 16 2 16 15 3 13 9 7 9 7 15 9 2 7 13 13 15 9 0 2 13 15 9 15 9 0 2 13 15 13 15 9 1 15 2
5 15 3 13 0 2
36 0 3 0 13 9 0 13 15 9 1 0 2 7 9 15 2 1 9 13 1 9 9 15 0 2 16 3 15 9 2 15 13 0 9 9 2
25 16 1 9 9 9 13 9 7 9 2 3 7 15 9 7 15 9 2 15 13 9 9 7 9 2
24 3 3 3 13 9 13 13 9 15 0 2 7 13 15 9 0 15 2 3 0 13 0 13 2
12 7 3 15 9 13 0 13 15 9 9 0 2
2 3 2
14 3 13 15 0 1 10 9 0 16 1 10 9 0 2
11 0 3 9 13 15 1 9 13 3 13 2
17 1 15 13 16 15 13 9 13 13 0 13 9 2 3 7 0 2
26 9 3 9 2 9 9 2 7 9 9 2 1 0 13 13 1 9 2 16 13 0 1 9 3 13 2
11 9 7 13 13 1 9 0 1 10 9 2
20 0 3 9 1 15 13 0 16 1 9 0 2 1 9 7 9 13 9 15 2
9 1 0 7 3 13 13 7 13 2
9 13 3 9 9 13 9 0 9 2
6 15 7 13 0 9 2
5 13 3 8 12 2
13 12 12 13 15 2 7 3 12 12 12 13 15 2
18 7 9 2 12 8 8 8 2 13 16 9 15 9 13 10 0 9 2
20 1 15 7 13 9 13 9 13 1 9 9 0 2 7 1 9 9 0 13 2
39 7 9 9 9 2 15 13 9 9 15 1 9 13 2 3 13 9 9 13 2 7 9 1 15 9 2 16 16 9 0 13 9 9 2 7 3 1 15 2
10 16 1 9 13 3 13 0 12 9 2
21 1 15 7 15 1 15 9 13 4 2 13 13 16 3 13 0 9 13 12 9 2
12 13 4 3 1 16 9 13 13 15 9 0 2
14 9 7 9 13 15 13 9 2 15 13 9 9 9 2
7 3 9 0 13 9 0 2
12 0 3 9 13 13 3 13 16 13 0 9 2
2 3 2
11 15 13 15 9 13 7 9 2 13 9 2
11 9 3 15 1 9 13 2 13 9 9 2
10 15 7 1 9 2 13 9 1 9 2
20 9 7 13 3 13 3 9 2 7 15 13 9 15 2 7 15 13 16 9 2
9 0 13 3 16 13 0 12 9 2
2 0 2
29 1 15 13 0 9 1 12 9 1 9 0 2 16 9 9 2 15 3 13 0 13 1 12 9 2 13 1 0 2
14 3 3 1 9 0 3 13 16 12 9 1 12 9 2
20 9 7 13 9 13 13 1 12 9 2 15 16 13 0 2 16 1 13 4 2
12 3 3 13 13 0 9 1 15 9 15 9 2
2 3 2
20 15 15 13 9 1 15 2 0 13 15 15 13 9 9 2 1 9 9 13 2
14 9 3 9 0 13 9 0 16 9 9 1 12 9 2
9 9 7 0 0 13 1 9 13 2
23 3 3 13 1 9 0 16 13 0 1 9 0 2 16 16 13 0 1 9 1 15 9 2
2 3 2
8 9 13 13 9 16 9 0 2
17 7 1 9 0 2 1 15 9 2 3 13 16 12 9 12 9 2
39 3 16 15 15 13 1 15 9 10 9 2 7 16 1 12 9 13 9 9 9 1 13 15 1 0 1 15 15 9 13 2 16 0 13 1 9 7 9 2
15 0 3 3 1 9 13 3 13 16 12 9 1 12 9 2
10 16 9 13 7 9 3 13 12 9 2
15 1 15 7 0 13 16 9 3 13 15 9 1 9 13 2
16 0 3 13 9 9 0 1 9 13 16 12 9 13 1 15 2
13 7 9 13 10 1 3 9 13 2 16 13 4 2
8 0 3 3 9 13 1 9 2
2 0 2
10 15 9 13 0 9 1 9 10 9 2
12 15 3 13 0 9 13 2 15 13 0 9 2
12 9 7 9 0 7 9 13 3 13 12 9 2
27 3 1 9 9 13 3 13 13 9 2 16 13 13 1 9 9 0 2 15 1 9 13 9 16 9 9 2
9 9 3 0 13 9 1 9 13 2
2 3 2
25 15 13 1 15 9 2 3 13 13 15 9 1 15 15 3 13 1 15 9 2 7 13 9 9 2
8 9 7 13 13 1 15 9 2
10 9 7 3 2 7 13 9 9 0 2
26 0 13 3 16 9 13 15 9 1 9 13 2 16 9 9 13 15 9 1 15 2 15 13 13 0 2
2 3 2
8 1 0 9 9 13 9 15 2
9 9 3 13 9 2 15 13 9 2
11 0 7 9 9 13 7 9 0 13 13 2
11 13 7 3 15 9 13 9 13 7 9 2
24 3 9 13 1 9 13 2 3 7 9 13 2 1 3 13 9 0 2 1 15 13 13 9 2
11 3 13 3 9 0 7 9 13 12 9 2
9 3 13 9 7 9 1 9 13 2
11 13 7 13 1 15 13 9 1 9 13 2
25 1 9 3 0 15 13 0 9 12 9 13 2 9 9 1 9 0 13 2 9 9 1 9 0 2
28 9 3 0 2 1 15 13 9 9 2 13 0 1 9 9 9 0 2 1 15 13 9 0 9 2 3 0 2
31 16 3 9 13 3 13 1 9 7 9 13 2 16 1 13 2 13 2 3 13 1 15 1 15 9 7 9 0 13 13 2
12 13 3 13 16 0 9 9 9 9 9 13 2
32 3 3 1 0 9 9 13 15 3 9 2 3 9 1 15 7 9 9 2 15 0 0 2 3 9 1 15 7 9 1 9 2
28 7 15 9 13 1 0 13 12 9 1 15 15 9 9 13 2 16 9 1 9 2 7 9 0 1 9 0 2
15 1 9 3 12 9 15 9 13 2 1 16 13 9 0 2
26 1 15 9 2 1 12 8 2 13 16 9 9 13 16 9 2 1 15 9 13 7 13 9 9 13 2
17 1 15 9 1 9 2 16 12 9 13 7 13 2 0 9 13 2
16 9 3 13 9 13 1 15 16 9 0 1 13 9 9 13 2
39 7 16 1 9 1 9 7 9 13 9 13 3 9 2 15 7 15 13 1 15 13 9 7 0 2 13 16 9 9 13 1 0 2 9 0 0 1 0 2
14 7 3 1 9 7 9 13 12 16 1 9 7 9 2
49 7 16 12 7 15 13 9 15 1 9 7 9 13 2 3 9 3 13 15 0 9 1 9 2 7 13 15 9 15 9 9 2 16 2 16 9 13 9 9 13 2 9 15 13 9 12 9 13 2
12 15 3 9 15 0 1 9 13 2 0 13 2
41 3 13 16 13 9 7 9 16 9 15 9 13 2 1 15 9 13 16 9 9 2 1 15 16 9 15 13 9 2 13 13 1 9 7 9 16 1 13 7 13 2
29 16 3 13 15 9 0 2 15 3 1 15 13 13 2 7 13 16 13 12 9 2 15 12 13 13 7 15 13 2
9 1 15 3 9 9 13 9 9 2
17 1 9 7 15 1 16 13 1 15 9 9 2 13 15 9 0 2
36 1 15 3 13 16 2 16 15 9 13 3 13 2 7 0 1 15 2 16 1 13 4 1 9 0 2 3 13 1 15 13 7 9 7 9 2
11 15 13 0 15 15 1 2 1 9 13 2
46 13 3 1 13 16 2 1 0 9 1 9 13 13 1 16 0 9 13 2 1 12 7 9 3 13 0 9 2 16 3 13 1 9 13 12 0 1 9 2 7 12 0 13 15 0 2
6 3 7 9 12 13 2
5 15 13 9 9 2
45 7 9 13 2 12 8 0 9 2 16 16 1 15 9 9 13 9 0 2 0 7 9 2 3 1 15 9 13 9 0 2 0 7 9 2 7 1 15 9 0 2 0 7 9 2
24 1 15 7 13 9 9 2 15 13 1 9 10 9 0 0 13 4 2 1 15 3 9 13 2
31 9 7 15 1 3 9 13 2 16 15 13 13 9 2 15 3 13 2 7 15 9 2 15 0 9 2 13 1 9 13 2
9 13 4 3 15 9 9 0 13 2
11 7 16 9 3 13 15 9 1 9 13 2
14 7 15 9 13 1 3 2 7 3 1 9 9 0 2
9 16 9 13 3 13 9 1 0 2
16 1 13 13 13 16 9 13 3 13 0 9 1 9 1 0 2
16 0 3 1 10 9 13 4 13 1 9 2 16 0 1 9 2
31 10 3 9 0 1 0 9 13 2 13 9 0 2 7 1 13 13 9 0 13 2 1 9 0 1 9 0 13 3 13 2
15 9 7 13 3 13 9 0 15 13 2 16 0 4 13 2
9 3 3 0 9 1 9 0 13 2
2 0 2
7 9 9 13 13 9 9 2
28 9 7 0 9 13 13 9 16 9 0 9 0 2 1 9 9 0 13 9 1 9 9 2 16 1 13 13 2
13 9 7 9 0 9 13 9 2 16 1 13 4 2
20 15 13 0 1 9 9 16 9 0 1 9 13 2 16 1 9 9 0 13 2
22 9 3 9 13 3 13 13 9 13 1 9 2 16 1 15 0 13 9 2 7 9 2
12 13 3 16 9 9 9 13 13 15 9 9 2
16 15 7 13 9 9 1 9 9 0 16 15 15 13 0 9 2
20 9 3 13 3 13 9 0 1 0 2 7 13 15 15 13 1 15 3 0 2
2 3 2
7 1 9 9 13 9 0 2
25 7 15 15 13 1 15 0 2 13 0 1 9 0 15 15 3 13 0 16 16 15 13 15 0 2
10 3 7 13 13 10 0 1 0 13 2
8 3 0 3 13 1 15 0 2
9 3 7 0 13 15 13 9 10 2
26 9 3 9 13 2 1 13 0 9 10 2 3 13 0 1 0 13 2 7 15 13 1 15 0 9 2
2 0 2
13 9 9 0 15 9 0 13 9 9 7 9 15 2
14 9 7 13 13 9 1 15 13 2 3 1 9 15 2
14 9 3 0 15 13 0 15 3 13 13 1 15 9 2
25 10 7 0 1 0 13 13 1 15 9 0 13 2 16 0 10 1 9 2 15 13 1 9 0 2
9 9 3 13 3 13 9 1 0 2
2 3 2
44 16 9 0 13 9 1 9 9 0 2 7 1 15 13 1 9 3 1 10 9 0 2 3 9 0 2 9 1 9 0 13 2 13 1 9 1 10 0 2 16 1 13 13 2
24 7 15 15 13 1 9 0 1 9 0 2 13 1 9 10 9 2 1 15 13 1 9 0 2
20 9 3 13 2 15 13 1 9 0 1 9 0 0 2 13 9 1 9 0 2
18 9 3 13 9 1 0 2 3 13 9 1 9 0 2 7 1 9 2
9 9 3 13 3 13 9 1 0 2
2 3 2
9 9 9 0 3 13 1 9 9 2
13 9 7 9 13 2 1 13 0 2 13 1 13 2
16 15 3 13 3 13 1 9 0 2 3 16 1 15 9 13 2
19 13 7 1 15 16 1 9 13 3 13 9 13 7 0 2 16 9 0 2
18 9 3 0 7 13 1 9 0 13 1 15 16 13 9 0 1 0 2
14 3 9 13 13 15 13 9 1 0 13 13 0 9 2
14 9 7 0 13 15 13 1 9 1 10 9 0 13 2
19 1 3 9 13 3 13 9 1 0 2 3 13 1 15 9 13 7 0 2
22 3 7 9 2 1 12 1 9 2 9 0 7 13 13 2 13 15 1 9 13 13 2
15 3 0 13 1 15 16 0 9 9 9 13 13 3 13 2
23 0 3 9 1 15 13 1 9 2 3 7 1 9 2 16 1 9 2 16 1 9 13 2
8 3 0 1 13 9 13 9 2
21 0 7 9 2 1 16 13 9 2 3 13 1 9 2 1 13 1 9 0 13 2
19 1 3 9 13 3 13 0 9 1 0 2 1 15 9 9 0 15 13 2
11 3 13 3 16 0 9 15 3 13 9 2
14 16 3 0 9 13 1 9 2 3 3 13 1 9 2
6 3 9 13 9 0 2
11 3 3 13 16 15 15 0 13 1 9 2
9 7 3 13 9 13 13 1 9 2
20 9 7 0 10 13 9 2 1 15 16 1 9 9 13 2 15 13 13 9 2
25 7 3 13 16 1 9 7 9 3 10 9 13 9 13 7 0 2 3 7 1 13 15 15 13 2
11 13 3 15 15 13 13 0 1 0 9 2
17 3 1 15 9 2 7 1 9 7 1 15 9 0 9 0 13 2
20 13 7 7 13 13 0 0 13 1 9 2 7 1 15 9 0 13 13 9 2
8 16 9 9 13 3 13 9 2
13 1 15 7 13 16 9 9 13 13 3 13 9 2
14 15 3 13 3 1 9 2 3 1 9 2 13 9 2
12 9 7 9 13 13 1 9 2 16 13 4 2
10 3 13 3 3 13 9 7 3 3 2
2 0 2
35 10 9 13 13 15 9 9 1 9 1 10 9 15 13 15 3 2 16 15 3 13 15 1 9 2 16 9 3 13 2 16 3 3 13 2
20 9 7 13 13 9 13 2 16 1 13 13 2 7 13 15 9 9 16 13 2
12 13 3 16 1 10 9 13 16 13 9 3 2
2 3 2
12 9 13 13 1 9 9 0 2 1 9 9 2
8 9 7 9 0 13 3 0 2
9 13 3 9 13 13 0 7 3 2
17 15 7 15 13 16 3 13 13 9 0 2 1 13 9 9 0 2
27 3 2 16 0 9 9 0 2 15 13 9 15 2 13 0 2 0 3 0 9 9 13 2 15 13 13 2
2 0 2
16 10 15 3 13 7 3 3 13 2 13 1 15 7 1 9 2
26 3 7 15 15 15 3 13 2 3 3 2 13 1 9 15 13 1 9 0 2 16 13 1 12 9 2
24 7 9 13 3 13 1 15 2 16 3 13 9 2 7 13 1 9 2 16 3 13 13 9 2
16 3 9 0 2 15 13 13 2 13 1 15 0 2 3 13 2
7 3 12 9 13 13 15 2
53 16 7 9 13 13 15 15 13 1 15 0 2 16 13 4 2 1 15 7 0 13 9 13 2 9 3 1 9 13 15 13 1 15 0 2 16 1 0 13 2 13 16 9 13 13 2 16 0 9 2 9 13 2
8 15 3 7 15 7 15 13 2
11 15 3 15 15 15 13 16 9 0 15 2
11 9 3 0 13 16 9 13 1 9 0 2
19 13 7 9 1 9 0 2 16 9 0 13 9 1 9 0 1 9 0 2
15 15 7 13 1 16 13 9 3 2 7 1 16 13 9 2
13 3 7 9 13 9 9 9 15 1 15 13 9 2
11 0 7 9 0 13 9 13 1 9 15 2
19 9 3 0 10 3 13 15 16 1 9 0 2 15 13 9 1 9 0 2
30 7 1 15 13 9 2 1 12 1 9 2 16 13 0 16 7 15 2 3 1 9 1 9 13 2 16 1 9 0 2
14 9 7 13 13 1 10 9 16 9 13 1 9 0 2
16 3 15 15 15 1 9 10 13 2 3 1 15 9 15 9 2
59 1 7 10 9 13 1 16 1 13 13 9 13 2 12 7 9 13 13 0 15 1 0 9 9 2 13 7 1 3 1 9 2 16 1 13 13 2 13 13 16 12 15 15 3 13 3 1 0 9 9 2 7 0 3 1 0 9 9 2
12 13 3 15 16 12 9 13 13 9 0 15 2
30 1 15 7 9 0 13 13 9 10 9 2 7 0 1 15 9 13 13 9 10 9 2 15 16 15 9 13 15 0 2
16 3 3 1 0 9 13 13 9 9 16 1 9 13 9 9 2
14 1 9 7 9 0 13 16 1 9 13 9 10 9 2
19 1 9 7 3 0 9 9 13 1 9 13 2 9 7 1 9 9 9 2
20 15 7 9 13 13 9 13 0 9 2 1 3 13 12 9 1 0 9 13 2
27 13 3 9 13 9 0 1 9 9 13 2 3 1 9 9 13 2 7 9 9 2 0 7 9 13 9 2
34 7 15 13 15 1 9 1 9 13 2 16 9 13 15 13 1 15 7 15 13 1 15 2 1 9 10 9 2 16 15 13 9 15 2
25 7 1 0 4 13 16 9 13 0 3 13 13 1 9 7 9 2 3 13 13 16 1 9 9 2
11 13 7 0 9 13 2 16 1 13 4 2
10 3 13 3 12 9 13 13 15 9 2
2 3 2
13 13 4 16 0 9 0 10 13 1 9 0 13 2
8 3 13 3 12 15 1 15 2
32 15 7 9 13 13 1 0 9 0 2 0 0 16 9 7 9 2 1 15 15 13 0 9 2 7 0 16 15 9 0 9 2
14 3 3 12 15 13 1 15 2 7 10 0 1 9 2
28 3 3 2 1 13 2 15 9 13 13 9 2 0 9 2 1 9 10 9 2 1 15 0 13 9 16 9 2
15 9 7 13 15 16 0 9 2 15 10 1 15 9 13 2
18 3 7 15 9 12 9 13 13 13 15 2 1 12 3 13 9 15 2
44 13 13 3 16 2 1 15 3 9 1 10 9 13 0 9 9 10 15 9 2 15 15 2 1 0 9 2 13 13 15 0 9 2 1 15 15 15 15 1 0 9 13 13 2
7 15 7 3 0 13 13 2
18 13 3 0 9 9 9 0 2 15 3 13 10 9 7 9 9 0 2
8 15 3 13 13 2 13 13 2
28 1 7 10 9 13 1 9 9 2 3 13 0 10 9 9 13 16 13 1 15 9 15 9 7 10 9 15 2
32 15 7 9 15 9 13 3 13 16 9 0 2 15 3 13 1 15 9 7 9 9 2 7 13 0 9 7 9 0 15 9 2
12 15 13 0 9 0 2 16 1 0 13 4 2
23 10 7 15 9 2 1 13 13 1 15 9 7 9 9 2 3 13 13 0 9 15 9 2
11 13 3 16 0 9 1 10 9 10 13 2
31 15 7 9 13 1 10 9 13 2 9 9 2 10 9 3 2 9 7 0 3 2 7 1 0 9 2 16 1 13 4 2
14 1 15 7 16 9 15 13 0 2 0 13 15 9 2
43 3 2 1 9 13 1 10 9 3 13 9 13 15 9 2 15 2 1 10 9 13 2 13 3 9 1 9 0 15 15 9 13 2 7 15 9 13 9 15 16 13 0 2
26 3 7 13 0 16 15 9 13 0 2 16 3 13 4 16 15 9 0 9 9 13 3 13 16 0 2
31 16 7 9 9 13 3 13 0 7 13 2 3 9 0 1 15 13 3 13 13 0 2 7 13 1 15 9 7 9 9 2
10 3 1 9 15 9 13 0 3 9 2
16 3 7 15 9 13 13 0 2 3 15 9 13 0 9 0 2
27 7 3 13 0 13 2 3 0 13 1 9 0 9 7 0 2 7 1 15 2 0 9 7 9 9 13 2
15 7 3 9 0 1 9 0 13 13 0 13 7 3 0 2
21 7 15 13 15 9 2 12 8 0 9 2 13 2 16 9 0 13 9 3 0 2
14 7 1 9 1 9 13 16 9 0 13 9 3 0 2
20 0 7 15 9 13 1 9 2 15 1 12 2 3 1 9 10 2 10 13 2
18 9 7 1 9 0 2 15 1 15 0 13 9 0 0 7 15 13 2
16 3 13 3 1 9 0 1 9 0 0 9 2 16 1 15 2
27 1 9 16 9 2 1 15 13 15 1 9 3 2 0 9 13 16 1 9 9 2 1 15 13 9 13 2
26 13 3 15 1 9 3 2 13 13 0 7 3 1 9 2 13 7 1 9 13 13 9 7 1 9 2
27 9 7 10 2 16 9 9 13 1 9 0 2 3 13 9 13 16 15 0 0 13 13 0 9 1 15 2
18 3 1 9 9 3 13 0 2 7 1 13 7 9 2 16 1 15 2
18 9 7 0 15 13 1 9 13 2 13 0 9 2 1 0 13 0 2
10 7 3 3 13 0 9 2 7 9 2
27 13 3 0 9 2 1 9 9 13 1 9 0 2 15 3 13 0 2 3 1 0 15 13 7 0 13 2
23 1 9 3 12 13 7 9 7 9 0 2 7 3 0 9 7 13 2 1 9 9 13 2
20 9 3 15 16 13 4 2 1 12 0 13 13 2 3 1 9 0 7 0 2
13 9 3 1 12 2 15 13 10 9 2 13 10 2
9 9 7 1 0 13 0 9 13 2
15 15 3 2 3 9 13 9 2 3 1 0 0 13 13 2
17 3 15 15 13 0 9 2 13 9 0 13 1 9 1 9 13 2
31 1 7 9 13 2 1 10 9 13 2 13 1 9 1 9 15 15 9 13 2 3 13 13 16 13 13 1 10 3 9 2
16 15 13 3 9 9 0 16 13 2 16 13 1 12 1 9 2
55 7 13 3 13 16 15 15 13 1 9 2 7 15 1 9 3 2 16 9 0 1 9 9 13 12 9 1 9 7 15 1 9 2 7 16 9 0 10 1 3 13 13 2 13 9 1 15 0 2 1 15 0 1 9 2
31 1 3 15 9 13 3 13 7 1 15 7 1 9 2 16 13 4 2 10 15 13 1 15 1 9 2 13 13 1 9 2
16 15 13 1 9 1 9 2 7 3 13 1 15 7 1 9 2
21 13 3 1 15 9 7 9 3 1 9 0 2 16 1 9 0 3 1 9 0 2
18 9 3 9 0 3 13 1 10 9 16 3 13 1 9 1 15 9 2
16 7 0 9 9 13 0 13 1 9 0 2 3 1 9 0 2
15 9 7 0 10 0 15 13 9 0 2 15 13 16 9 2
15 3 3 13 9 13 15 9 0 16 13 1 9 1 15 2
27 7 1 15 13 1 9 1 9 2 16 9 13 0 9 2 16 3 15 9 9 15 13 0 1 9 0 2
13 7 3 1 3 0 9 12 9 13 15 13 13 2
35 9 7 15 13 13 16 2 1 9 13 1 9 13 0 2 3 13 13 16 1 15 9 0 12 1 15 13 2 7 1 9 15 9 13 2
25 15 3 16 9 15 1 9 0 13 2 13 13 9 0 1 15 16 3 13 1 10 9 0 9 2
8 3 13 16 1 9 13 13 2
28 15 3 13 13 9 9 13 2 1 12 8 2 16 1 9 13 1 9 3 13 9 2 13 2 7 15 13 2
10 15 7 16 13 2 13 9 3 0 2
16 0 3 2 16 9 1 9 13 13 1 9 2 1 9 9 2
15 0 13 7 13 3 12 9 13 13 12 15 16 13 15 2
2 3 2
17 10 9 7 13 13 1 10 9 2 15 9 13 2 16 9 9 2
9 3 7 15 13 15 9 9 13 2
21 3 13 7 13 0 16 12 9 13 13 9 15 2 1 13 15 9 13 1 15 2
12 0 3 13 16 12 13 1 15 1 9 10 2
2 0 2
5 13 13 9 13 2
9 3 13 7 9 9 13 9 0 2
21 13 3 16 0 9 3 13 2 16 1 9 10 15 13 2 7 3 1 9 15 2
2 3 2
10 0 13 1 9 3 1 15 15 13 2
20 15 7 9 13 9 16 0 9 2 15 13 1 10 1 9 2 9 7 9 2
21 0 3 13 16 9 13 1 9 10 13 1 15 2 7 3 1 9 15 1 15 2
28 7 15 3 13 0 13 1 9 9 2 15 13 16 13 13 1 15 16 13 1 9 13 12 1 9 1 9 2
23 3 9 13 2 16 13 1 15 0 9 2 3 3 1 15 13 16 1 9 15 13 12 2
10 3 7 9 13 15 13 1 9 10 2
13 7 1 15 13 15 9 2 7 13 2 7 13 2
14 1 7 9 9 2 13 13 1 9 9 1 9 0 2
17 3 3 12 9 13 13 15 1 15 9 13 2 16 15 0 13 2
12 0 3 9 2 3 15 10 9 13 7 13 2
11 9 0 0 2 3 15 13 16 10 9 2
20 3 7 9 13 2 12 8 1 8 8 2 16 0 9 0 13 3 9 9 2
6 16 9 13 13 0 2
20 1 13 3 9 0 9 13 3 0 13 15 9 13 2 7 3 9 9 0 2
27 1 3 9 15 13 9 0 9 2 3 15 1 9 13 2 13 16 10 9 2 3 9 0 2 0 13 2
10 1 9 7 0 13 3 9 9 0 2
6 15 3 9 13 13 2
2 3 2
31 1 9 9 13 16 9 9 2 16 1 13 4 2 13 16 1 9 0 13 0 15 13 1 9 2 16 0 9 13 0 2
29 1 3 9 13 13 1 9 0 2 13 16 15 15 13 1 9 0 1 9 0 2 13 1 9 13 1 9 0 2
16 15 3 13 1 15 2 13 1 15 1 9 15 1 15 13 2
2 3 2
36 16 9 13 13 9 0 2 16 9 13 2 15 13 1 9 9 0 13 15 9 16 9 2 15 16 13 13 2 9 7 13 13 16 0 9 2
7 13 7 7 13 1 9 2
17 13 3 13 15 15 13 1 9 9 0 16 9 13 1 10 9 2
14 9 3 15 15 13 7 13 2 13 0 1 9 13 2
25 3 7 9 2 1 9 1 9 2 13 16 1 9 15 13 1 9 2 13 9 15 13 1 9 2
15 13 3 9 13 3 0 9 13 2 7 3 9 9 0 2
24 3 2 16 13 9 0 7 0 9 2 16 0 9 2 0 3 9 9 0 2 3 0 9 2
43 16 0 9 9 13 13 1 9 2 13 10 9 1 15 13 1 9 2 13 7 9 13 10 9 7 9 9 2 0 13 16 9 13 15 13 10 9 0 7 15 9 15 2
22 1 7 9 1 9 9 13 13 1 9 2 13 15 13 16 9 13 3 13 9 0 2
11 9 3 13 16 9 0 13 9 9 13 2
18 7 16 0 13 2 9 13 13 9 13 1 10 9 15 13 1 9 2
14 3 3 9 15 13 1 9 2 13 9 9 0 10 2
22 9 7 9 0 1 9 9 13 13 0 2 1 9 9 13 2 3 1 9 9 0 2
19 3 3 13 9 16 15 9 13 13 9 9 9 13 2 16 0 9 15 2
6 16 9 13 13 0 2
51 16 0 9 9 1 9 9 13 13 0 16 1 9 10 2 7 0 1 15 16 1 15 15 13 2 1 9 9 0 9 13 3 0 13 9 0 1 9 9 7 9 2 16 9 10 2 7 3 1 9 2
49 1 3 9 9 1 9 13 13 13 0 2 3 13 2 1 16 13 1 9 10 2 13 9 13 0 2 15 1 9 13 2 15 16 9 9 10 1 3 13 13 9 16 12 13 0 1 9 12 2
47 3 2 16 9 9 9 3 13 13 1 9 9 7 9 2 16 1 15 9 13 2 3 9 9 9 3 13 13 1 9 9 13 2 15 13 9 0 2 16 1 15 9 1 10 9 13 2
50 9 0 9 9 13 2 1 13 0 9 2 3 15 12 7 0 13 2 13 13 1 9 9 9 7 13 2 3 16 1 15 9 13 3 0 9 9 7 9 2 7 3 9 2 13 13 1 10 9 2
20 7 13 16 9 1 15 13 2 13 0 2 7 16 13 0 2 1 9 9 2
2 3 2
12 15 13 9 9 2 13 7 0 2 7 13 2
14 3 9 9 13 1 0 2 9 0 13 1 12 3 2
13 9 3 2 3 13 0 2 3 3 13 7 13 2
9 1 0 0 9 9 13 7 13 2
19 3 13 16 0 9 0 2 15 12 9 0 13 2 12 9 9 0 13 2
11 9 7 0 13 9 9 9 16 9 13 2
17 15 7 0 13 0 7 0 1 12 9 2 3 1 9 7 9 2
20 9 3 13 2 15 13 9 2 13 15 9 9 1 12 9 2 3 1 9 2
2 3 2
16 9 9 0 0 9 13 1 9 10 2 7 1 9 9 13 2
17 1 9 3 10 13 1 9 9 2 1 9 1 9 0 7 13 2
10 3 1 15 0 13 3 13 1 15 2
13 1 9 7 9 13 13 9 0 3 1 9 9 2
26 13 3 9 0 1 9 10 1 0 0 9 9 0 2 15 16 3 13 1 9 13 2 7 9 0 2
15 13 7 0 3 0 9 2 7 9 2 15 13 9 9 2
20 9 3 9 9 13 15 9 13 2 7 3 0 9 9 2 7 3 9 13 2
17 3 13 3 0 9 13 9 13 2 16 9 10 0 13 3 13 2
2 3 2
28 16 9 0 13 1 9 13 2 1 9 9 2 1 9 13 13 7 13 1 9 2 13 16 13 0 15 13 2
5 15 13 15 0 2
5 3 0 0 13 2
22 9 3 2 15 13 1 9 2 13 15 0 2 15 3 13 13 1 9 13 1 9 2
12 13 3 13 16 9 13 0 13 15 0 9 2
9 3 9 13 0 9 13 10 3 2
46 16 0 9 1 9 13 13 1 9 2 16 9 1 9 13 0 1 9 2 15 7 3 13 3 13 0 1 9 2 0 13 16 9 9 13 13 9 0 0 2 16 3 1 13 4 2
19 7 13 13 16 3 10 15 13 13 1 9 15 9 0 9 13 1 9 2
44 1 3 9 13 13 3 13 2 7 1 15 13 9 10 9 2 1 9 15 13 2 16 13 9 0 2 16 15 13 1 13 9 2 7 2 16 13 0 2 16 13 12 15 2
12 3 7 15 15 9 13 2 3 10 9 13 2
28 9 3 0 2 1 0 9 13 2 13 12 2 15 13 2 7 1 15 3 9 13 10 15 1 12 9 13 2
28 10 3 13 16 12 0 16 4 1 12 13 2 16 7 9 10 3 13 0 1 3 13 7 13 16 12 15 2
12 15 0 15 1 0 9 13 2 3 13 3 2
15 7 3 2 16 13 9 12 2 3 13 13 1 9 12 2
10 13 3 1 9 9 13 15 9 9 2
17 3 3 9 2 0 13 2 1 3 13 9 9 2 7 9 9 2
27 9 7 0 2 16 1 12 2 15 13 10 9 2 10 13 2 7 10 9 13 10 9 2 10 3 13 2
23 3 1 9 15 3 13 15 9 2 7 10 13 13 15 3 9 2 13 1 10 9 9 2
2 6 2
10 9 0 9 7 9 0 1 10 9 2
7 16 3 13 9 9 10 2
15 16 1 9 15 13 10 9 9 2 7 9 9 15 13 2
15 16 15 13 9 7 15 13 15 2 7 0 9 15 13 2
3 8 12 2
43 12 13 0 9 2 15 9 9 0 13 2 15 9 13 2 1 0 4 13 2 15 1 10 9 9 10 13 9 13 2 16 3 0 0 9 2 7 7 9 10 13 13 2
20 9 7 15 13 3 9 9 2 7 1 10 9 9 2 16 1 0 13 0 2
9 3 13 13 16 13 10 13 9 2
10 3 1 15 15 10 9 13 2 13 2
33 15 7 9 1 9 1 15 13 9 13 2 16 15 1 15 13 7 0 9 9 13 2 7 9 9 2 1 13 15 9 0 9 2
16 15 7 15 1 9 13 9 2 15 1 9 1 9 15 13 2
23 9 3 7 9 13 9 0 9 2 3 0 13 16 15 1 9 13 2 1 9 15 13 2
25 9 7 0 15 9 1 10 13 9 2 15 13 1 9 13 1 15 15 9 9 13 1 15 13 2
31 0 13 3 16 9 2 15 13 1 15 0 9 7 10 9 1 10 9 9 13 2 10 9 9 13 2 1 15 3 13 2
20 7 13 15 15 1 15 9 13 2 16 7 13 15 15 1 15 9 3 13 2
17 13 3 2 16 9 1 13 7 13 2 3 3 7 1 13 9 2
13 15 0 9 9 1 0 13 9 2 1 9 9 2
19 15 3 3 1 9 13 4 16 2 9 13 2 15 9 13 7 9 13 2
19 3 7 15 3 0 13 13 2 7 7 15 13 1 0 9 1 13 9 2
18 15 16 1 10 9 0 13 9 2 1 0 9 13 1 0 9 13 2
9 13 7 16 1 1 10 9 13 2
18 15 0 2 9 9 2 15 1 10 9 3 13 2 7 1 15 13 2
46 15 15 2 0 13 2 16 1 9 0 13 3 13 9 2 3 1 0 9 1 9 1 9 15 13 3 13 2 7 0 9 0 13 13 2 16 13 9 0 2 15 9 3 0 13 2
19 15 0 2 0 13 2 0 9 13 13 9 2 15 3 1 15 9 13 2
8 3 2 12 13 2 15 13 2
20 7 0 1 9 0 1 0 9 13 2 15 3 9 1 15 9 3 13 13 2
19 1 15 13 16 7 15 15 1 9 0 9 13 13 2 9 0 13 13 2
19 3 7 15 0 9 2 16 1 15 9 13 4 2 3 9 15 9 13 2
23 15 3 2 0 13 9 2 9 13 2 16 15 0 9 13 2 0 13 15 0 13 9 2
52 9 3 2 1 15 16 13 9 2 9 2 1 15 16 13 0 9 2 3 15 13 1 10 9 9 13 2 9 2 1 15 16 13 9 0 1 10 9 2 16 2 16 13 0 13 2 10 3 15 9 13 2
7 0 7 15 13 9 9 2
33 7 3 3 1 0 2 15 2 15 9 13 2 1 15 13 0 9 2 15 13 15 2 7 3 13 2 16 3 13 9 9 10 2
34 3 0 1 0 2 15 2 3 16 13 3 1 0 9 2 1 9 3 0 13 3 13 2 13 2 16 1 9 15 13 10 9 9 2
32 3 0 1 0 9 2 15 10 9 9 13 2 3 0 9 2 7 3 0 9 0 9 13 2 13 2 7 9 9 15 13 2
24 0 0 15 0 9 9 13 2 16 0 13 16 15 15 1 9 4 13 2 1 15 3 13 2
12 7 15 13 15 13 2 16 15 13 9 8 2
51 16 3 1 0 9 1 9 0 9 13 4 2 1 0 7 1 9 9 15 2 1 16 13 9 10 9 7 9 2 13 1 15 0 9 13 1 9 9 7 9 15 2 1 16 13 9 10 9 7 9 2
18 13 3 15 9 13 2 16 0 13 1 15 1 16 13 9 10 9 2
13 0 2 1 9 0 15 2 1 16 10 9 13 2
12 0 2 1 0 9 2 16 13 9 9 13 2
7 16 10 9 13 1 9 2
14 13 13 3 0 2 16 10 9 1 13 13 15 9 2
19 1 15 3 15 0 1 9 13 2 15 13 13 9 1 15 13 9 9 2
32 15 3 13 13 13 9 2 13 7 1 15 13 13 1 9 13 2 16 13 1 9 13 1 9 2 7 9 13 1 0 9 2
18 7 13 2 3 1 15 2 3 15 13 1 9 13 13 2 7 3 2
13 16 3 9 13 9 13 2 3 13 9 9 9 2
9 10 7 9 9 1 15 0 13 2
20 3 3 1 15 9 15 9 13 2 7 1 9 3 9 2 1 9 7 9 2
9 3 7 9 1 9 0 9 13 2
27 9 0 3 3 13 1 15 13 2 16 9 1 9 2 9 1 9 2 3 7 3 2 16 13 7 13 2
18 7 16 3 9 13 1 15 13 2 9 9 13 1 9 1 15 13 2
15 16 7 3 13 1 15 13 2 9 9 13 1 15 9 2
21 13 3 16 10 9 1 13 13 9 2 3 3 9 15 2 3 15 1 9 13 2
2 3 2
19 1 10 9 1 9 2 15 13 0 9 13 2 1 15 9 3 13 15 2
18 16 9 9 13 1 1 9 2 15 0 13 2 3 13 1 15 0 2
15 7 1 9 15 9 13 13 15 1 15 9 3 13 15 2
7 15 3 9 1 0 13 2
18 15 3 13 0 2 16 2 1 0 3 13 13 2 9 13 3 13 2
11 15 3 13 1 15 1 15 0 13 13 2
7 10 3 9 13 1 9 2
2 0 2
20 16 9 9 13 1 0 2 13 16 7 1 15 9 13 15 13 2 7 3 2
14 16 3 13 15 13 2 9 15 13 13 1 0 9 2
15 15 7 13 0 2 0 13 13 2 1 3 13 0 13 2
20 15 7 0 13 13 2 0 13 13 2 7 15 0 13 13 2 0 13 13 2
15 0 13 3 16 9 13 13 15 13 1 15 13 9 0 2
63 16 7 1 15 9 3 13 15 13 2 13 9 3 9 13 7 1 9 9 0 2 16 16 9 13 16 13 2 13 7 16 13 2 13 7 16 13 2 7 1 9 9 2 16 13 9 16 13 9 2 15 13 16 13 9 13 2 15 13 16 13 9 2
30 3 7 13 0 13 1 0 7 1 9 0 2 16 7 1 9 9 2 16 13 1 12 8 2 9 3 13 13 9 2
20 7 1 9 2 16 7 1 9 2 1 13 12 0 9 2 16 1 13 4 2
10 3 13 3 0 16 9 1 0 13 2
10 13 3 13 15 15 13 9 9 13 2
7 10 3 9 13 1 9 2
2 3 2
25 1 15 15 13 1 9 2 10 0 1 0 9 7 0 9 13 9 9 0 7 9 0 9 13 2
28 16 3 9 9 3 13 1 15 13 2 7 9 2 16 13 4 2 13 1 0 2 13 9 0 1 0 13 2
9 15 13 0 2 16 1 13 4 2
11 0 13 3 16 9 9 13 1 15 13 2
2 3 2
11 10 9 7 13 1 9 2 7 1 9 2
13 1 9 7 1 9 3 13 0 16 13 1 9 2
17 13 3 13 1 9 15 15 1 9 13 2 7 1 15 9 13 2
7 15 3 13 13 1 9 2
33 16 7 1 9 13 13 15 9 9 1 15 1 9 13 13 2 3 1 9 0 13 9 0 9 2 1 15 9 1 15 9 13 2
9 3 9 13 9 2 7 9 9 2
18 16 3 9 1 9 13 1 9 13 1 10 9 2 3 9 1 9 2
7 10 3 9 13 1 9 2
2 0 2
26 9 3 13 16 1 15 15 13 1 9 2 7 3 13 15 1 9 16 13 1 15 1 15 3 13 2
16 9 3 13 1 9 16 13 1 13 2 3 7 9 7 9 2
31 7 9 13 1 15 15 13 1 9 2 16 1 9 3 0 13 2 7 1 15 15 13 1 9 2 16 13 1 9 0 2
18 3 3 9 1 9 2 16 9 1 9 7 1 13 2 13 1 9 2
2 3 2
15 16 9 3 13 1 15 9 13 2 10 9 13 15 0 2
16 16 7 0 15 13 1 0 2 3 3 12 15 13 16 15 2
16 3 1 13 1 15 3 13 15 9 16 1 15 13 1 12 2
6 0 3 13 16 13 2
14 10 3 9 13 1 15 13 9 2 15 13 9 15 2
30 13 7 15 9 15 3 13 13 1 9 2 16 9 0 7 0 2 7 9 15 1 9 13 2 16 9 9 7 3 2
13 1 15 15 13 13 16 13 15 9 3 1 9 2
16 7 13 16 9 0 3 13 1 15 9 2 7 15 13 9 2
18 9 7 0 3 13 9 2 1 15 0 13 1 9 15 1 9 13 2
14 3 7 13 1 9 2 16 1 13 16 3 0 13 2
37 9 7 15 13 1 9 2 3 13 1 9 2 7 1 15 13 9 7 0 9 2 16 9 9 9 13 13 9 9 9 2 15 13 1 9 9 2
12 7 15 1 15 9 13 2 16 1 9 9 2
23 1 15 7 13 0 0 9 2 15 13 10 13 1 9 9 2 9 0 1 9 3 13 2
7 16 10 9 13 1 9 2
13 1 15 7 0 13 13 16 10 9 13 1 9 2
18 3 3 0 13 10 9 13 1 9 2 16 15 9 13 1 15 13 2
13 15 7 1 15 9 13 13 2 13 13 13 15 2
12 3 3 13 1 15 16 1 15 9 1 15 2
10 15 7 13 13 15 2 13 15 0 2
7 3 10 9 13 1 9 2
2 3 2
15 9 13 1 15 13 9 9 7 13 2 7 15 15 13 2
11 15 7 13 1 9 9 2 16 13 9 2
7 3 9 13 15 10 13 2
9 10 3 9 7 9 13 1 9 2
2 3 2
25 10 9 7 9 1 9 15 9 13 13 2 7 16 13 1 9 7 9 2 7 16 1 0 13 2
10 15 7 15 15 13 9 2 9 13 2
6 7 3 10 13 13 2
9 10 3 9 7 9 13 1 9 2
2 0 2
9 10 9 7 9 13 1 15 9 2
15 16 3 15 9 13 9 2 0 13 16 13 9 0 9 2
31 16 7 9 13 9 0 9 2 0 13 16 13 13 15 9 13 1 9 13 2 1 15 3 13 0 2 16 13 9 0 2
10 15 7 13 13 9 15 13 9 9 2
9 10 3 9 7 9 13 1 9 2
2 3 2
8 10 9 13 1 16 13 9 2
7 13 7 13 1 15 0 2
6 3 13 1 9 15 2
7 9 7 10 13 9 9 2
11 3 9 3 13 16 1 9 13 1 9 2
7 10 3 9 13 1 9 2
2 3 2
11 9 1 9 13 1 9 16 13 15 9 2
35 9 7 1 9 2 16 13 1 9 2 16 13 4 2 3 3 13 15 9 2 1 3 13 9 9 2 7 13 1 9 13 15 1 15 2
13 9 7 1 9 3 13 15 9 16 1 9 9 2
14 0 3 3 13 16 1 9 9 2 15 13 9 9 2
28 3 7 9 1 9 3 13 7 13 1 15 9 16 1 16 13 9 2 1 9 1 9 13 9 1 15 9 2
7 10 3 9 1 9 13 2
2 3 2
20 15 9 13 13 9 7 13 9 2 16 15 9 13 13 1 3 7 13 3 2
6 10 7 13 9 13 2
15 3 9 1 9 15 9 15 13 2 16 13 15 16 9 2
19 10 7 9 0 2 3 13 1 9 2 3 13 9 2 15 13 9 15 2
6 10 3 13 1 9 2
2 3 2
17 15 13 1 15 9 9 1 9 15 2 13 1 9 7 9 13 2
35 13 7 1 9 9 13 7 3 7 0 15 0 13 2 16 1 9 9 3 13 13 16 13 9 2 7 9 9 3 13 16 9 13 13 2
16 16 3 15 13 1 9 0 9 2 15 13 1 9 7 9 2
5 7 15 13 0 2
20 3 15 15 13 3 7 0 2 3 13 0 7 0 2 7 15 13 1 0 2
10 0 3 9 13 1 15 15 0 13 2
8 7 0 0 15 13 1 9 2
8 10 3 9 13 9 1 13 2
2 3 2
12 10 15 13 13 1 9 9 1 13 7 9 2
9 13 3 13 7 13 1 15 13 2
20 15 7 13 2 1 13 1 9 2 13 1 9 2 7 3 1 9 7 9 2
9 1 9 3 13 1 9 1 9 2
13 3 7 13 7 9 3 1 13 7 13 13 9 2
8 15 13 15 9 13 9 13 2
6 9 13 15 10 13 2
18 7 9 2 12 8 2 1 0 9 2 13 16 10 9 7 9 13 2
8 16 9 13 1 9 1 9 2
13 1 15 7 13 16 9 1 9 13 1 9 9 2
20 15 3 1 9 13 0 1 15 15 13 13 1 9 2 0 13 1 9 13 2
12 9 7 0 13 1 9 2 15 13 10 9 2
7 13 3 9 1 9 13 2
2 3 2
28 9 1 9 7 9 13 15 9 1 9 9 2 16 1 15 9 9 13 9 0 2 7 1 9 9 13 9 2
18 9 7 13 1 16 13 1 9 0 2 3 1 15 15 9 9 13 2
9 1 7 16 13 2 3 13 9 2
6 13 3 9 13 9 2
12 15 3 13 13 9 9 2 13 1 9 9 2
5 15 7 13 9 2
6 13 3 9 1 9 2
2 3 2
9 1 15 13 9 0 7 9 13 2
17 0 7 13 1 15 1 9 2 1 9 7 1 9 7 1 9 2
9 15 3 0 1 9 7 9 13 2
40 9 3 2 1 13 1 12 9 2 13 1 9 1 9 15 7 9 9 3 13 2 16 2 1 13 1 9 9 2 13 1 9 1 9 9 7 9 9 9 2
8 7 1 15 9 9 13 3 2
19 1 9 3 9 1 16 13 9 2 1 9 7 9 9 1 16 13 9 2
14 3 7 9 7 9 9 13 1 9 2 7 1 9 2
6 3 3 13 1 0 2
17 13 7 0 9 3 1 9 13 2 13 0 15 1 9 13 0 2
9 3 15 13 1 9 13 1 9 2
19 13 7 1 15 16 13 1 9 15 13 2 15 9 15 9 1 9 13 2
19 9 3 9 1 9 7 9 1 15 13 1 9 2 9 0 13 1 9 2
8 7 0 13 13 1 10 9 2
28 7 3 1 15 9 13 9 7 9 1 15 2 16 2 1 15 13 1 0 1 0 2 13 0 7 13 0 2
17 9 7 13 1 16 9 13 9 1 9 2 7 9 1 9 0 2
9 9 7 1 16 4 13 9 13 2
19 10 3 15 13 13 1 10 9 13 1 9 2 13 7 1 9 1 9 2
17 3 2 1 10 9 7 13 13 1 9 2 9 13 1 9 9 2
2 0 2
12 1 9 1 9 7 9 15 2 9 13 9 2
10 1 15 3 13 9 15 13 16 9 2
36 16 3 13 1 15 15 3 13 9 13 2 13 1 9 2 16 2 16 15 13 13 9 2 7 13 9 13 15 13 9 2 15 13 1 9 2
21 7 10 9 1 9 13 1 15 1 15 13 15 1 9 9 2 16 1 0 13 2
15 16 3 15 3 13 0 2 7 0 2 15 13 1 9 2
11 9 3 1 9 3 13 9 16 1 9 2
25 1 3 13 1 0 13 0 9 1 9 7 1 9 2 9 3 13 1 9 15 9 16 1 9 2
20 15 13 16 9 13 2 12 8 1 8 8 2 16 9 13 1 9 7 9 2
16 9 15 13 13 16 9 3 13 1 9 2 7 9 15 2 2
9 13 7 15 15 15 9 9 13 2
17 15 3 13 1 9 9 2 13 13 0 7 0 7 1 0 9 2
21 9 7 13 3 13 0 7 0 2 7 16 1 0 9 2 7 3 7 1 0 2
8 1 0 3 3 9 9 13 2
31 1 9 3 1 9 1 0 13 13 2 1 0 13 1 9 13 2 16 13 9 1 9 2 16 13 9 2 1 12 9 2
9 3 3 13 9 13 13 1 9 2
2 3 2
12 9 1 12 8 2 13 13 16 9 13 0 2
42 7 15 13 1 15 16 15 0 13 0 2 0 7 13 13 0 0 3 13 0 13 2 7 0 13 3 13 0 13 2 7 1 15 16 9 13 0 3 0 13 9 2
10 3 13 3 9 1 9 7 9 13 2
2 3 2
9 10 9 0 13 9 13 1 9 2
10 9 7 13 9 0 2 16 7 9 2
27 9 3 15 2 15 13 9 13 9 9 2 13 13 1 9 2 16 3 9 7 9 2 15 13 9 9 2
24 16 7 13 9 9 0 13 2 13 13 16 9 13 13 7 1 9 15 2 7 1 9 15 2
19 9 3 1 9 15 13 1 15 16 13 15 15 15 13 4 7 13 13 2
19 16 3 9 3 13 9 2 3 13 15 9 2 16 3 4 13 15 13 2
25 16 3 9 9 0 3 13 2 3 13 9 2 16 16 13 4 13 2 3 3 13 13 16 13 2
26 13 3 9 16 3 13 9 2 15 13 4 7 13 13 2 16 13 9 2 15 3 3 13 9 9 2
21 10 7 9 2 16 0 7 13 13 2 13 15 15 15 13 4 13 7 13 13 2
10 1 9 3 3 13 3 13 9 9 2
33 9 7 2 1 13 9 1 10 9 2 10 3 13 4 13 2 15 3 13 15 13 2 1 1 15 12 15 13 13 9 1 9 2
12 15 3 15 13 13 15 15 15 1 9 13 2
19 3 3 13 13 9 16 13 9 9 2 7 13 13 9 16 13 9 9 2
34 9 3 9 3 2 13 1 9 2 3 13 9 9 2 7 13 1 15 15 13 9 2 13 9 15 2 16 9 9 9 13 9 9 2
35 7 16 3 9 7 9 7 9 3 13 13 16 1 16 13 1 9 2 16 3 9 13 9 1 9 1 9 1 15 13 2 13 9 0 2
11 3 7 2 13 9 15 2 7 3 0 2
9 9 3 13 9 2 13 9 0 2
16 9 7 13 9 9 2 3 13 9 0 2 7 13 9 9 2
13 9 7 9 7 9 13 1 9 2 13 9 9 2
23 7 16 15 9 13 13 15 9 7 15 9 2 0 13 16 15 9 1 9 0 9 13 2
25 15 3 13 2 13 13 16 3 10 15 13 1 9 2 13 13 0 7 0 2 16 0 9 13 2
47 16 3 15 13 1 9 2 13 13 1 15 15 13 13 7 3 7 0 2 3 13 0 7 0 2 16 1 15 15 13 9 9 13 2 16 1 9 9 13 9 2 3 13 0 7 0 2
9 13 7 0 16 13 16 1 0 2
15 9 3 9 0 2 16 13 1 9 13 2 13 3 3 2
9 3 3 9 12 4 13 9 15 2
25 3 9 3 13 0 7 16 1 0 2 16 9 3 3 13 9 0 2 7 15 2 16 13 4 2
25 16 7 13 15 9 15 13 15 15 13 13 13 2 13 0 7 0 9 2 16 1 13 9 0 2
23 15 3 3 13 1 9 1 15 15 13 13 2 7 13 15 13 2 1 9 13 9 13 2
12 9 7 9 13 1 0 9 1 9 9 0 2
40 3 16 9 13 9 0 2 15 9 13 1 9 2 7 3 13 0 2 16 1 9 13 13 1 15 13 2 16 3 15 9 7 3 7 0 13 15 9 9 2
11 13 7 0 16 15 9 0 15 13 9 2
16 1 9 7 0 9 13 1 9 15 0 2 16 13 13 9 2
13 3 0 3 13 2 7 0 2 1 15 13 9 2
48 16 3 15 9 15 13 2 13 13 9 9 1 9 7 3 7 0 2 13 9 0 3 0 2 7 7 3 7 0 2 16 13 1 15 15 13 13 9 1 9 2 15 9 13 4 9 9 2
7 3 9 9 3 13 0 2
28 13 7 0 9 16 1 15 15 13 2 13 15 13 16 1 0 2 16 1 15 2 13 1 9 2 13 9 2
44 16 7 3 0 15 13 16 1 0 15 9 9 1 9 13 2 1 15 13 16 0 13 1 9 2 15 16 0 13 15 0 2 7 3 0 13 1 0 2 1 15 13 9 2
11 1 0 7 15 9 13 9 9 1 9 2
29 1 15 13 16 2 16 9 1 9 13 2 13 3 0 2 16 0 9 13 2 16 3 1 15 2 7 1 9 2
12 9 3 13 0 9 2 15 15 1 15 13 2
44 9 7 13 15 3 15 15 13 1 15 2 3 16 0 3 13 2 16 15 13 9 1 9 9 9 2 3 13 9 9 2 7 9 2 9 7 13 3 0 2 7 9 9 2
25 0 1 15 9 0 13 15 13 13 0 9 2 3 13 9 2 7 13 15 0 2 7 1 15 2
17 7 3 15 9 9 7 13 13 13 0 2 16 9 9 1 9 2
9 15 7 9 13 9 1 0 9 2
19 3 3 13 9 9 1 9 9 2 7 1 13 7 9 9 1 9 9 2
15 9 3 3 13 9 9 3 1 9 9 2 7 3 15 2
23 3 3 13 1 9 9 0 16 3 13 9 2 7 16 13 9 2 15 13 3 13 9 2
12 15 3 16 13 13 9 2 13 9 1 15 2
19 16 0 13 3 13 9 2 3 13 16 16 13 13 15 16 13 13 9 2
20 3 3 9 1 9 3 4 1 15 13 2 7 1 9 2 9 0 1 15 2
23 13 3 1 13 16 15 15 13 0 9 2 3 13 1 9 1 9 9 2 16 9 0 2
22 15 0 3 13 0 2 7 15 9 2 3 13 13 1 9 1 15 2 7 1 9 2
7 16 9 3 13 15 9 2
12 1 15 7 13 16 15 9 13 1 15 0 2
21 9 3 2 16 13 4 2 15 13 15 16 9 15 15 15 13 4 7 13 13 2
10 3 3 1 10 13 9 15 9 0 2
13 9 7 3 13 15 9 2 7 13 9 1 9 2
9 9 3 3 13 15 9 1 9 2
2 3 2
7 15 1 10 9 13 9 2
9 16 7 13 9 2 13 15 9 2
20 3 2 16 9 13 15 10 13 2 13 15 9 9 13 2 1 10 13 13 2
10 1 15 3 15 9 13 15 9 13 2
6 9 7 7 9 13 2
9 15 3 13 0 1 16 9 13 2
6 15 3 9 0 13 2
2 0 2
10 10 9 7 13 9 2 7 4 13 2
19 9 7 3 13 13 9 2 16 15 13 2 13 16 13 9 13 7 9 2
7 7 0 3 13 4 13 2
9 3 15 9 9 13 9 7 9 2
9 15 3 9 1 10 9 13 0 2
2 3 2
6 15 13 1 10 0 2
10 15 3 13 15 13 15 0 7 13 2
11 10 7 9 13 13 9 2 16 13 4 2
10 15 3 9 2 16 3 2 13 0 2
2 3 2
7 10 9 13 15 9 0 2
12 16 3 13 1 9 9 2 13 15 9 9 2
41 16 0 13 1 9 9 2 13 16 1 9 15 9 13 2 7 3 15 9 13 0 2 16 9 15 9 3 13 0 2 16 9 13 0 9 2 16 13 0 9 2
13 15 7 13 1 15 0 2 3 13 13 15 0 2
16 1 9 3 9 13 9 15 15 13 15 13 13 7 13 15 2
17 9 3 2 1 13 15 15 13 0 9 2 3 13 13 15 0 2
17 3 7 15 0 13 15 2 13 15 9 2 7 9 16 15 13 2
8 15 3 9 13 1 15 0 2
2 0 2
15 15 13 9 15 2 7 15 13 9 2 7 13 9 15 2
10 1 9 3 13 15 1 9 7 9 2
31 9 7 2 16 3 2 13 9 9 2 1 13 9 9 2 7 9 15 13 10 13 2 7 9 15 15 13 9 9 13 2
12 15 3 13 9 15 2 16 3 2 13 9 2
7 9 3 3 13 9 15 2
2 3 2
7 9 1 9 7 9 13 2
21 9 7 2 16 3 2 9 13 2 16 1 16 15 13 9 2 1 15 13 9 2
6 9 3 0 15 13 2
12 13 3 9 1 9 2 16 1 15 9 13 2
10 7 13 3 9 13 2 3 15 0 2
8 7 13 1 15 9 1 9 2
9 7 9 3 13 15 16 1 9 2
16 10 3 15 13 2 15 9 13 2 16 13 9 2 9 13 2
7 9 3 3 13 15 9 2
2 0 2
18 13 4 1 0 15 2 16 10 9 2 15 9 13 2 13 1 9 2
10 9 7 13 9 9 2 1 0 13 2
21 1 3 9 9 9 13 3 13 2 0 13 15 9 2 16 13 9 2 13 9 2
7 15 13 15 8 12 13 2
11 13 9 10 15 13 2 7 13 3 0 2
4 7 8 12 2
7 10 13 0 1 9 10 2
5 7 12 8 12 2
5 10 9 9 0 2
33 7 9 2 8 12 1 8 8 2 13 16 9 3 13 13 2 3 1 15 2 7 15 1 13 2 3 9 2 16 9 7 9 2
16 1 15 7 13 9 9 2 13 15 9 1 10 9 13 0 2
17 9 15 13 13 16 9 13 9 7 9 15 2 7 9 15 2 2
9 13 7 15 9 13 9 13 13 2
9 1 0 3 9 0 15 9 13 2
16 9 7 13 9 0 1 15 9 2 3 1 9 7 9 0 2
20 16 3 9 1 10 9 13 0 9 2 3 0 9 13 0 9 1 10 9 2
8 7 0 1 9 9 7 9 2
8 9 3 13 13 9 15 9 2
10 13 3 15 9 2 7 15 9 0 2
2 3 2
6 15 0 13 9 15 2
13 16 3 15 13 2 15 0 13 9 7 9 0 2
8 7 9 7 9 13 13 0 2
6 9 3 13 9 15 2
2 3 2
13 9 7 9 13 13 9 0 1 9 2 1 9 2
9 15 7 9 13 9 7 9 15 2
20 3 3 9 3 13 9 7 9 2 7 3 15 3 13 2 3 13 13 9 2
8 9 3 13 15 9 7 9 2
2 3 2
8 10 15 13 2 13 9 15 2
6 9 7 13 16 9 2
7 13 3 9 7 13 15 2
10 9 3 2 16 9 2 13 9 15 2
2 0 2
15 1 15 13 3 7 0 2 13 16 13 9 15 13 9 2
10 9 3 7 9 3 13 3 7 0 2
8 13 7 1 0 12 15 0 2
12 13 3 2 16 13 2 16 9 13 9 15 2
2 3 2
5 9 7 9 13 2
6 13 7 9 1 9 2
7 3 13 9 15 7 9 2
8 15 7 9 3 0 13 13 2
21 9 3 7 9 1 0 0 9 13 2 16 0 9 13 2 16 0 1 9 13 2
13 1 15 3 15 1 9 9 13 2 15 13 0 2
8 9 7 9 13 9 7 9 2
21 3 1 9 9 0 13 2 16 7 0 9 1 9 9 0 2 16 9 1 9 2
27 16 3 9 7 9 13 1 0 9 1 9 2 7 9 9 2 13 16 1 0 0 9 13 9 7 9 2
9 12 7 9 13 13 12 9 0 2
6 0 7 9 13 9 2
14 13 3 16 1 9 9 13 15 1 0 0 7 0 2
19 15 3 1 0 13 9 1 9 15 13 1 9 2 13 1 9 10 0 2
16 15 0 13 9 1 9 0 9 9 2 13 1 9 10 0 2
23 9 7 15 2 16 13 9 9 2 13 3 15 9 2 16 0 1 9 2 7 15 3 2
17 3 7 1 15 9 13 9 2 7 9 3 1 13 1 9 13 2
11 7 13 15 13 9 12 2 13 9 15 2
45 7 3 7 9 2 1 16 13 9 0 1 9 0 2 13 15 15 13 1 9 10 9 2 7 15 15 1 15 13 0 2 9 7 9 2 16 13 9 9 2 15 13 9 9 2
17 1 15 3 13 16 9 7 9 13 0 1 16 1 9 0 13 2
20 3 7 0 13 2 16 0 9 13 2 7 9 9 13 9 2 16 13 9 2
26 15 3 9 13 13 9 16 9 7 9 2 16 13 1 0 2 13 9 0 2 1 15 0 9 13 2
26 10 3 0 0 7 15 13 9 2 16 9 7 9 2 7 12 9 7 15 9 2 16 9 7 9 2
38 13 3 9 0 7 9 7 9 2 3 1 16 13 9 9 9 2 1 15 13 9 2 7 1 9 9 7 9 13 1 15 9 15 13 13 9 9 2
37 16 9 0 13 9 9 3 16 13 0 2 7 16 13 15 9 2 7 0 13 9 9 3 1 9 9 2 7 9 15 9 1 15 13 9 9 2
61 13 3 13 16 9 13 9 7 9 13 9 2 3 1 0 9 2 1 1 0 12 9 2 1 15 15 13 15 9 2 15 3 13 2 7 1 9 9 2 15 13 9 7 9 13 0 9 7 0 9 2 7 1 15 15 13 13 12 0 0 2
25 1 9 3 13 2 0 2 12 2 0 2 0 2 13 2 13 2 9 2 13 2 7 0 9 2
28 1 9 7 2 0 2 0 2 0 2 0 2 0 2 13 2 0 2 9 2 15 9 0 2 7 0 9 2
22 3 7 7 1 0 9 0 9 13 9 2 1 9 15 9 2 3 0 1 15 9 2
8 13 3 7 15 9 15 9 2
12 3 0 13 15 0 13 2 1 15 13 0 2
17 10 3 0 12 13 9 2 7 15 13 2 3 9 15 13 13 2
19 16 0 7 0 13 9 2 0 0 7 0 13 0 2 3 1 9 13 2
35 16 3 10 9 7 9 1 9 9 13 2 10 7 9 7 9 1 9 9 2 3 1 0 15 1 9 13 13 2 15 1 9 9 13 2
12 7 1 15 9 7 9 9 0 10 13 13 2
15 1 15 3 13 15 9 13 9 2 1 15 0 9 13 2
42 1 3 16 9 7 9 2 15 13 9 9 2 7 13 13 0 9 2 4 13 9 0 9 7 9 0 2 9 15 13 1 15 9 7 15 9 2 13 9 7 9 2
17 1 9 3 2 3 9 2 1 16 3 2 3 13 15 9 9 2
36 1 15 3 1 12 8 1 8 8 2 13 9 2 16 9 3 13 1 9 16 9 9 2 1 15 0 13 0 7 0 2 3 15 9 9 2
31 9 3 13 13 9 3 0 13 9 9 2 16 13 4 2 7 0 1 15 2 16 13 9 13 9 16 13 15 9 9 2
13 1 15 9 13 9 9 13 16 13 15 9 9 2
14 13 7 15 15 3 7 0 9 2 1 9 1 9 2
15 3 3 15 9 13 2 13 7 13 2 16 0 7 0 2
18 13 3 0 15 13 1 9 3 13 2 7 0 0 3 1 9 13 2
17 3 7 3 9 13 15 13 3 13 9 2 3 3 1 0 13 2
25 9 7 13 3 3 15 9 13 2 16 9 7 9 2 16 0 9 13 2 7 1 9 9 13 2
19 16 9 0 13 3 0 13 13 9 9 2 3 3 0 1 9 9 13 2
49 13 3 9 13 1 9 2 3 3 9 15 13 2 7 9 15 13 2 16 0 9 13 2 7 15 9 15 13 16 9 15 0 13 15 0 2 16 9 7 15 9 13 13 16 9 9 13 0 2
11 9 3 0 13 2 16 9 1 0 13 2
15 12 9 2 1 16 13 9 9 2 7 13 1 12 9 2
8 7 3 15 9 13 13 9 2
9 15 9 2 1 16 13 9 9 2
15 7 3 9 7 9 13 9 2 16 9 13 15 13 13 2
6 16 9 9 13 9 2
13 1 13 7 13 13 16 9 3 13 16 1 0 2
28 16 3 15 9 13 9 9 2 9 7 3 13 16 9 9 2 16 13 4 2 13 15 9 13 9 0 9 2
2 3 2
8 15 3 13 2 15 13 9 2
8 10 3 9 13 13 9 15 2
11 9 7 3 13 9 15 2 16 13 4 2
8 9 3 3 13 13 15 9 2
13 13 3 16 1 15 13 9 2 16 15 13 9 2
2 3 2
14 15 13 0 7 1 15 15 9 2 13 1 0 9 2
17 16 3 9 13 1 15 15 9 2 13 1 0 9 2 3 9 2
5 15 7 13 0 2
9 3 13 4 16 10 9 13 9 2
14 9 3 1 15 3 13 9 15 2 7 0 1 9 2
11 10 7 9 1 9 13 1 9 1 15 2
18 0 7 9 13 13 1 15 9 2 7 9 3 13 13 1 15 9 2
7 9 3 13 4 1 9 2
2 3 2
15 10 9 7 13 9 2 7 9 2 7 9 2 7 9 2
10 9 7 3 13 13 7 9 7 9 2
17 13 4 3 1 16 3 9 9 2 7 9 1 9 2 13 9 2
17 0 3 13 13 9 2 1 15 13 1 16 13 9 7 9 13 2
15 7 3 13 13 9 2 1 13 1 9 2 16 13 4 2
8 9 3 3 13 13 15 9 2
14 16 3 15 13 9 9 2 13 16 4 1 9 13 2
43 1 7 9 7 9 13 13 2 12 7 13 3 13 13 9 15 16 1 9 2 16 0 13 2 16 13 1 12 9 2 13 16 9 3 13 13 9 0 9 16 1 9 2
17 15 7 9 1 0 13 13 7 1 9 9 2 7 1 9 9 2
45 1 9 3 9 2 16 1 9 13 9 9 2 1 15 13 16 9 13 0 7 9 13 2 16 2 1 9 9 13 13 0 2 13 0 9 7 9 0 2 15 13 15 9 9 2
13 13 7 9 2 16 13 9 2 16 9 9 13 2
17 3 3 13 1 16 13 15 9 2 7 1 16 13 15 1 9 2
10 16 3 3 9 13 2 3 3 13 2
16 3 3 9 13 1 9 1 9 9 2 16 9 13 13 9 2
33 1 15 13 16 9 3 13 9 13 2 7 13 2 16 9 3 13 1 9 13 16 16 13 13 9 2 7 1 15 3 13 13 2
33 1 15 7 13 16 9 9 7 9 13 1 9 9 2 7 15 15 15 13 1 9 9 2 16 1 9 9 13 9 1 9 9 2
10 15 3 9 13 2 7 9 7 9 2
24 1 9 0 9 2 9 1 9 13 1 9 2 3 1 9 9 9 2 7 1 9 9 15 2
26 16 3 9 13 0 1 13 9 9 2 0 13 9 13 1 9 2 16 1 0 9 13 1 9 9 2
17 7 15 13 1 15 9 9 2 16 9 0 3 13 1 9 9 2
38 15 3 9 0 13 9 13 1 9 10 9 2 15 16 3 13 2 3 1 15 13 13 1 9 2 7 3 0 16 13 1 9 9 15 13 1 9 2
34 1 9 7 9 9 2 1 9 9 13 16 9 15 1 9 13 9 15 9 2 3 3 1 9 12 9 2 0 13 15 9 13 9 2
20 7 15 9 3 13 9 9 13 1 9 2 16 1 13 13 2 7 15 9 2
14 3 3 1 0 13 16 9 1 9 3 13 1 9 2
8 15 7 9 7 1 0 13 2
15 9 3 1 10 9 13 9 2 7 0 9 1 15 13 2
8 1 0 7 13 15 15 13 2
23 3 3 1 9 9 13 13 0 9 2 1 9 9 0 9 7 0 13 2 7 3 13 2
16 9 3 3 13 9 2 15 9 13 2 7 3 9 7 9 2
10 0 3 13 13 9 9 2 3 0 2
17 16 3 13 13 2 13 3 1 15 0 2 3 0 1 15 0 2
21 0 3 3 1 15 2 16 9 0 1 0 9 13 2 3 7 1 15 9 13 2
10 3 9 0 3 13 0 2 7 0 2
5 9 7 0 13 2
14 7 3 13 4 16 1 15 0 9 13 16 1 9 2
17 9 3 0 3 13 1 9 7 9 9 2 7 0 13 1 9 2
11 1 9 7 0 13 1 9 12 0 9 2
18 15 12 13 9 0 2 3 9 9 2 15 13 9 1 13 9 9 2
12 3 15 9 1 9 13 2 15 13 15 9 2
30 9 0 13 1 9 9 0 2 15 13 15 13 9 7 9 2 15 13 9 9 2 12 1 13 13 2 15 1 13 2
9 15 7 9 0 13 1 9 13 2
11 0 3 0 9 1 9 0 13 9 13 2
4 0 9 0 2
3 0 9 2
9 0 9 9 2 15 13 9 9 2
11 9 7 9 13 3 13 9 7 9 0 2
14 3 3 1 9 3 9 0 13 16 1 16 13 0 2
22 3 2 16 9 13 9 0 2 7 9 0 0 13 2 0 7 2 16 15 13 0 2
17 15 7 1 9 0 13 16 9 0 13 13 9 1 9 3 13 2
10 9 3 3 13 9 9 2 7 9 2
14 3 3 9 13 9 9 9 7 0 13 2 7 13 2
14 9 0 15 9 13 0 9 2 0 13 1 9 9 2
14 13 3 1 9 0 0 9 2 7 15 9 9 0 2
30 15 3 9 0 9 2 1 15 13 2 0 9 13 2 1 15 9 9 0 7 13 7 13 2 16 7 9 13 9 2
10 0 3 9 7 9 13 13 7 13 2
27 13 3 16 0 9 1 0 9 9 0 7 0 13 2 7 0 3 1 15 9 0 13 2 16 0 13 2
12 1 9 3 9 13 13 9 7 9 9 0 2
7 13 7 15 9 13 9 2
19 1 3 9 13 13 1 9 0 9 2 13 13 9 1 9 1 9 0 2
11 15 3 9 16 13 0 2 3 13 9 2
8 3 3 9 1 13 0 13 2
7 15 9 9 0 13 13 2
24 16 7 9 13 0 2 3 13 9 0 2 15 9 3 13 13 2 7 3 9 1 0 13 2
20 13 3 13 16 9 1 9 13 3 13 0 2 16 13 9 1 15 9 13 2
22 7 3 0 7 0 2 3 3 13 1 15 0 13 2 0 3 13 0 7 1 9 2
4 13 3 0 2
11 3 3 9 0 2 16 13 1 0 13 2
9 15 3 15 13 13 2 13 13 2
11 15 3 0 9 9 9 1 0 0 13 2
9 9 3 0 13 1 9 0 9 2
36 1 3 0 9 13 1 9 0 9 2 0 13 2 13 7 1 13 16 13 15 1 9 0 9 13 2 16 13 1 9 1 13 1 9 9 2
25 13 4 7 16 1 9 9 0 12 9 9 13 2 3 9 0 2 7 9 13 2 15 13 9 2
26 1 7 15 0 13 0 9 2 3 15 9 0 13 13 9 15 9 2 7 15 15 2 7 15 15 2
19 16 3 9 0 0 9 13 9 0 0 2 3 9 0 9 13 9 15 2
35 3 2 1 9 0 9 7 0 9 13 13 2 15 7 13 0 9 2 7 9 13 9 7 0 9 2 3 9 15 2 7 9 15 13 2
19 1 3 9 13 1 9 13 1 9 9 13 15 0 9 2 13 13 9 2
30 1 7 9 1 9 13 1 9 0 0 2 7 15 9 15 15 9 13 1 0 9 0 2 13 1 9 9 9 0 2
16 13 3 1 9 9 9 9 9 1 9 2 7 1 0 9 2
20 1 9 3 2 16 1 2 1 13 9 9 2 9 1 9 0 1 9 13 2
36 1 9 0 13 2 16 1 9 1 15 9 13 13 15 3 13 2 7 3 7 15 9 2 0 2 7 3 9 1 15 13 3 1 0 9 2
7 15 7 9 9 0 13 2
11 3 1 9 15 9 13 13 7 3 13 2
22 3 13 1 9 15 16 9 9 13 2 7 1 9 13 2 7 16 15 7 15 13 2
8 7 3 15 9 13 9 0 2
22 16 3 9 15 13 2 7 13 9 15 2 3 13 9 2 16 9 1 9 0 13 2
6 15 3 13 9 9 2
19 3 3 3 1 0 7 1 0 13 16 9 1 9 3 13 16 1 9 2
6 16 9 13 1 9 2
14 1 13 3 13 13 16 10 9 13 1 15 9 13 2
20 9 3 3 13 13 1 15 13 2 1 3 13 9 13 2 16 1 13 4 2
9 13 3 16 9 13 1 15 9 2
18 10 7 9 2 1 13 9 15 2 9 15 13 2 16 1 13 13 2
8 10 3 9 1 9 15 13 2
2 3 2
10 9 9 15 13 2 16 1 13 13 2
10 9 7 7 9 13 1 15 9 13 2
14 9 7 9 13 9 1 9 1 9 2 15 9 13 2
9 3 1 15 9 13 9 7 9 2
15 9 3 2 15 9 13 2 13 1 9 15 16 1 9 2
2 0 2
9 1 15 13 15 9 2 16 13 2
7 3 7 16 16 13 9 2
12 13 3 9 0 13 2 1 9 9 13 0 2
14 3 7 13 2 0 13 2 9 2 16 13 1 9 2
10 3 3 9 9 13 16 1 15 13 2
8 13 3 16 9 13 1 9 2
2 3 2
12 9 3 13 16 1 9 2 7 1 9 3 2
15 10 7 15 13 1 9 2 13 1 15 15 13 1 15 2
30 13 3 3 1 9 13 2 15 13 9 9 1 13 2 13 9 15 15 13 9 9 1 15 2 3 16 13 9 15 2
14 3 15 13 1 9 2 13 1 15 15 13 1 15 2
34 7 1 9 7 9 13 13 2 12 7 13 3 13 13 15 9 2 7 13 15 2 13 15 0 9 13 9 16 9 9 9 13 13 2
9 3 13 7 9 2 16 9 13 2
22 3 9 0 13 16 7 9 2 1 10 9 2 16 3 2 13 9 2 16 13 4 2
14 3 13 7 9 16 3 9 13 1 9 16 1 9 2
19 9 3 15 13 3 9 2 7 3 9 15 13 9 2 15 13 9 15 2
13 3 3 3 9 13 1 9 15 13 16 1 9 2
18 9 3 3 13 3 9 0 2 7 3 9 15 2 15 3 13 9 2
13 3 13 3 1 9 16 1 9 2 7 1 9 2
19 0 7 9 3 13 16 1 9 1 9 15 13 2 7 15 1 9 13 2
14 7 1 15 15 9 2 16 9 9 13 1 9 9 2
21 9 7 9 2 15 13 9 9 2 13 1 9 2 15 13 9 16 9 1 9 2
7 16 9 3 0 13 9 2
16 13 7 1 13 16 2 15 13 9 2 3 13 15 9 13 2
12 3 3 13 16 13 9 9 2 16 9 13 2
6 9 7 9 13 9 2
5 13 3 3 9 2
24 7 1 13 9 1 0 13 2 3 7 1 9 9 13 9 2 13 1 0 1 9 13 9 2
12 9 7 15 1 9 13 13 2 13 13 13 2
15 3 0 9 3 13 0 9 2 16 1 0 9 13 4 2
10 13 3 16 3 15 13 9 1 9 2
15 3 16 1 13 15 0 13 2 13 15 3 1 9 13 2
36 3 7 13 13 2 16 13 15 2 16 13 9 2 1 15 9 13 15 7 0 2 1 0 13 2 9 3 13 13 2 16 1 0 9 13 2
25 3 16 1 0 9 0 13 2 3 1 0 0 2 7 3 1 0 13 2 3 15 3 13 13 2
15 7 3 1 15 9 9 3 0 13 13 13 0 1 9 2
22 0 3 15 2 15 0 13 2 0 13 1 9 0 16 0 0 2 16 15 9 13 2
14 15 7 1 9 15 9 1 9 13 2 3 13 13 2
12 3 3 9 3 1 9 4 13 2 13 0 2
9 7 3 1 0 9 3 13 13 2
11 3 9 13 13 13 0 2 7 0 0 2
17 3 3 3 0 13 1 9 1 9 0 9 9 2 9 13 15 2
5 13 3 15 13 2
18 1 13 3 0 13 16 9 0 9 15 13 13 13 2 16 9 9 2
10 13 7 16 13 9 15 13 9 9 2
23 15 3 2 16 9 13 2 13 9 9 2 1 16 13 9 1 9 9 15 13 1 9 2
15 3 3 0 13 1 9 1 15 9 2 3 0 13 9 2
57 9 7 13 0 9 1 9 2 3 3 1 0 9 15 9 9 2 7 1 15 16 15 9 9 13 2 7 1 15 16 9 13 1 0 9 16 1 9 9 13 13 2 16 9 3 13 0 9 0 2 3 1 15 3 9 13 2
14 13 3 9 1 9 3 13 0 16 1 9 15 13 2
10 15 3 13 15 15 4 13 1 9 2
27 13 3 16 9 13 1 9 9 2 15 3 13 15 9 2 1 15 13 9 15 9 2 15 13 15 13 2
24 3 3 15 9 13 1 15 1 9 9 13 9 2 3 13 2 3 9 1 9 0 13 3 2
9 7 3 3 1 9 13 13 9 2
14 15 7 9 9 1 9 3 13 1 0 1 0 13 2
20 3 9 0 7 9 10 13 4 2 7 13 1 15 9 1 15 13 3 13 2
27 3 13 3 7 9 15 0 2 7 9 0 9 1 0 13 2 16 1 15 13 1 0 9 9 1 9 2
10 1 0 7 13 15 9 1 0 13 2
11 3 9 7 9 1 10 9 9 3 13 2
8 13 3 9 13 1 0 13 2
9 3 0 9 9 7 9 0 13 2
9 7 0 9 1 13 1 0 13 2
17 15 3 13 9 13 2 13 3 13 15 13 2 7 3 1 0 2
18 3 7 9 3 1 9 0 13 2 3 0 13 1 0 7 13 9 2
15 15 13 1 15 1 15 1 13 9 3 4 9 9 13 2
12 1 0 3 1 9 9 9 0 9 13 13 2
11 3 3 0 13 2 7 3 9 13 13 2
7 16 9 13 15 9 9 2
24 1 13 7 13 13 16 2 16 9 3 13 9 1 15 2 15 3 9 13 13 9 1 9 2
15 15 3 13 1 15 16 1 9 2 13 16 13 15 9 2
13 13 3 7 1 9 9 2 7 1 15 0 9 2
13 9 7 13 1 9 16 1 9 2 16 13 4 2
7 13 3 16 9 13 9 2
2 3 2
19 15 13 1 9 1 15 13 2 3 13 1 9 15 15 16 1 15 9 2
9 15 3 9 13 15 13 1 9 2
13 9 7 13 9 15 15 15 13 4 7 13 13 2
8 1 15 3 15 13 9 13 2
16 13 3 9 1 9 15 13 1 9 1 15 7 1 10 13 2
8 13 3 16 9 13 15 9 2
2 3 2
14 15 13 15 1 10 9 2 13 15 1 15 15 9 2
14 10 3 1 15 15 13 15 0 13 16 15 15 13 2
18 3 9 3 13 3 16 1 15 13 2 7 9 13 16 1 15 13 2
22 9 7 3 13 1 9 15 15 13 2 1 13 9 15 15 13 4 15 7 13 13 2
16 3 13 16 9 3 13 15 9 2 7 1 15 7 1 9 2
2 0 2
14 10 0 13 1 15 0 2 16 9 13 1 15 9 2
25 7 10 9 13 15 9 2 1 0 9 2 1 15 3 13 15 9 2 16 1 0 9 13 4 2
13 10 3 9 13 15 9 2 1 15 13 1 9 2
7 16 9 13 9 1 9 2
20 1 15 3 13 16 9 2 16 3 13 9 1 15 2 13 3 9 1 9 2
32 16 3 15 13 9 15 1 15 2 15 15 13 15 2 13 9 15 1 9 2 16 0 15 13 9 2 13 9 9 1 9 2
8 10 7 9 13 1 15 9 2
9 9 7 10 13 15 15 9 9 2
20 9 3 13 3 9 9 2 7 3 1 0 2 7 0 13 1 9 7 9 2
27 3 3 13 9 1 0 1 9 2 16 15 13 15 9 2 1 9 13 1 9 7 13 1 9 0 9 2
7 9 3 13 1 9 9 2
2 3 2
10 9 13 9 15 2 16 1 13 13 2
17 9 7 13 9 1 9 1 9 0 2 16 9 7 9 1 15 2
8 9 3 13 15 9 1 9 2
2 3 2
8 1 9 9 13 9 1 9 2
8 9 7 1 9 13 15 9 2
26 3 3 13 13 9 1 15 2 16 9 3 13 9 1 15 16 13 13 2 7 1 15 16 13 9 2
9 16 3 15 13 2 15 13 9 2
13 9 3 13 15 9 3 1 15 2 7 1 9 2
2 3 2
13 1 10 9 9 13 2 13 9 13 1 9 9 2
18 1 9 3 9 0 16 1 9 13 13 9 13 9 1 9 7 9 2
15 1 9 0 9 0 2 16 1 9 9 13 1 9 9 2
15 1 9 0 9 0 2 16 12 9 3 13 15 9 9 2
19 1 9 0 9 0 2 16 0 9 13 9 2 16 1 15 9 13 13 2
17 13 3 16 9 13 9 1 9 2 7 3 13 13 9 1 15 2
6 16 3 13 0 9 2
18 1 15 7 13 16 3 13 13 15 0 9 2 15 13 10 9 9 2
22 0 3 9 13 13 1 9 10 9 2 16 7 0 9 13 15 13 3 13 1 9 2
20 3 13 7 13 15 9 3 13 1 9 2 1 13 4 16 9 13 1 9 2
6 3 15 13 0 0 2
2 3 2
26 16 15 13 0 0 2 13 16 1 9 10 13 0 2 16 7 0 0 13 15 1 10 9 0 13 2
17 15 7 13 0 2 1 9 3 13 15 9 2 16 1 13 4 2
12 0 13 3 13 0 9 2 15 13 0 9 2
2 3 2
12 15 15 13 0 9 2 3 4 1 15 13 2
11 10 7 9 13 1 0 2 16 13 4 2
7 3 13 3 9 0 9 2
2 0 2
12 9 3 13 16 9 9 2 16 1 13 13 2
7 0 7 9 13 9 0 2
8 9 3 3 13 13 0 9 2
2 3 2
26 1 15 15 13 1 9 2 13 0 15 15 13 1 15 2 0 13 16 13 0 15 15 13 1 9 2
15 9 7 3 13 16 1 9 7 1 9 2 16 13 4 2
9 0 13 3 16 9 13 0 9 2
2 3 2
11 10 9 13 9 1 9 2 16 13 4 2
13 0 7 9 3 13 9 7 1 15 7 1 9 2
11 9 3 3 13 13 0 9 1 15 9 2
2 3 2
10 9 1 15 0 13 15 15 1 9 2
13 7 9 3 13 9 16 1 9 2 16 13 4 2
8 9 3 3 13 13 0 9 2
19 1 15 7 13 9 9 2 13 15 0 9 2 15 13 9 0 10 0 2
7 16 9 15 9 13 9 2
22 16 7 10 9 13 1 0 2 16 1 13 4 2 13 0 16 15 9 9 13 9 2
10 10 3 9 13 1 9 1 10 9 2
17 13 3 16 7 15 9 13 9 2 7 9 9 13 3 9 9 2
5 15 13 15 9 2
2 0 2
10 9 9 15 13 1 15 13 9 15 2
8 9 7 15 9 13 1 9 2
10 3 3 9 13 9 2 15 10 13 2
8 15 3 9 9 13 15 9 2
2 3 2
22 15 1 15 15 13 1 1 15 13 2 7 1 15 13 1 15 13 2 13 9 15 2
17 15 7 2 16 9 0 13 2 1 15 13 2 3 1 15 13 2
9 16 0 15 13 2 1 15 13 2
8 9 3 15 9 13 15 9 2
7 9 7 15 13 9 15 2
9 15 3 13 1 9 16 1 9 2
2 3 2
28 15 9 13 1 9 15 15 13 9 2 7 15 15 9 3 13 2 16 15 13 9 2 1 15 13 1 9 2
20 15 7 3 13 2 13 1 9 3 1 15 13 2 16 13 1 13 7 9 2
14 7 15 15 13 9 2 3 13 1 9 16 1 9 2
23 3 9 2 15 13 9 9 13 2 3 13 1 15 16 1 9 9 2 15 13 15 9 2
15 3 7 15 15 9 3 13 2 13 1 9 16 1 9 2
6 9 3 10 13 9 2
11 16 10 13 1 12 9 2 15 13 9 2
15 1 15 7 13 16 10 13 1 12 9 16 1 0 9 2
24 16 3 15 13 1 15 16 1 9 16 16 15 13 9 2 3 13 16 9 16 9 13 9 2
11 15 3 13 0 9 2 13 0 10 9 2
18 7 0 9 13 12 3 2 15 13 9 2 16 1 0 9 13 4 2
13 10 3 13 16 1 9 1 12 9 15 13 9 2
2 3 2
30 15 13 0 1 15 9 2 13 9 10 15 15 13 15 9 2 16 9 2 15 13 0 2 13 9 9 1 15 9 2
15 0 3 9 2 15 13 9 2 13 9 9 1 10 9 2
21 3 7 13 9 15 9 15 13 9 2 1 15 13 9 2 13 3 16 13 9 2
10 1 15 7 13 15 2 7 15 3 2
8 9 3 0 13 10 9 9 2
2 3 2
13 1 15 9 9 9 0 13 3 9 16 9 0 2
11 3 9 0 3 13 9 16 1 9 0 2
23 15 3 15 13 9 0 1 9 9 0 2 13 16 13 3 9 0 15 16 9 0 0 2
17 7 9 13 0 9 1 9 9 0 2 1 13 0 1 9 9 2
11 13 3 3 9 15 9 16 15 9 0 2
2 0 2
51 1 10 9 13 13 16 0 9 13 9 10 13 9 2 16 2 16 9 13 16 13 9 2 13 7 16 13 2 13 7 16 13 2 13 7 16 13 2 13 16 9 13 9 7 9 7 9 7 15 13 2
19 7 10 13 1 0 9 9 13 1 12 0 9 2 15 13 9 10 9 2
21 7 1 15 2 1 9 13 9 9 2 10 13 1 9 16 9 13 1 9 0 2
8 13 3 16 10 9 13 9 2
2 3 2
10 9 0 13 1 9 0 16 1 9 2
8 9 3 9 13 1 9 15 2
11 3 7 9 9 13 0 16 9 12 9 2
19 9 7 0 2 15 13 9 2 13 9 0 2 1 1 15 0 9 13 2
19 9 7 15 15 9 0 13 2 13 9 0 15 7 15 15 1 15 13 2
15 10 3 9 13 16 1 9 1 12 9 2 15 13 9 2
2 3 2
8 1 9 9 13 9 1 9 2
22 3 16 0 9 13 10 0 9 2 3 1 9 0 9 13 16 13 10 9 0 9 2
11 15 3 13 0 9 2 13 1 9 10 2
21 13 7 0 9 10 9 9 2 13 10 1 10 9 2 7 1 13 1 10 9 2
16 3 13 16 10 9 0 9 13 1 0 9 1 9 10 0 2
14 9 7 0 9 10 13 9 2 16 1 0 13 4 2
21 9 7 15 15 15 9 13 16 10 9 2 15 13 15 2 16 1 0 13 4 2
22 10 3 15 4 13 7 1 15 0 2 7 13 9 0 2 1 9 13 16 1 9 2
6 10 7 9 13 3 2
17 3 2 16 1 0 13 2 15 13 13 15 1 15 3 13 9 2
9 10 3 13 1 9 16 1 9 2
2 3 2
12 9 0 15 13 2 16 13 13 2 13 15 2
29 13 3 13 1 15 1 15 2 7 16 15 3 1 15 9 13 2 15 13 1 9 10 7 0 7 0 7 0 2
24 9 7 13 9 0 9 10 2 15 3 0 2 15 7 13 15 9 2 16 1 13 13 0 2
7 13 3 15 9 9 10 2
2 3 2
20 9 1 15 9 9 13 2 7 1 15 10 15 9 13 16 13 9 1 9 2
12 9 3 3 13 16 1 9 2 16 13 4 2
9 1 9 7 9 1 9 9 13 2
25 3 9 13 9 15 9 9 2 7 0 9 15 9 9 2 1 9 9 2 7 1 13 1 9 2
12 9 3 0 13 9 16 13 9 13 16 9 2
12 3 3 13 15 1 9 0 16 1 9 0 2
8 13 3 9 0 0 10 9 2
20 13 7 0 10 9 0 13 0 9 13 2 15 9 13 2 16 1 13 4 2
7 9 3 13 0 10 9 2
7 15 13 15 13 8 12 2
7 0 1 15 13 4 9 2
4 7 8 8 2
10 15 13 9 7 8 2 0 7 0 2
6 3 9 13 9 9 2
9 13 3 13 3 9 13 10 9 2
7 15 3 1 13 13 0 2
15 3 3 13 0 9 10 9 16 3 13 0 10 1 13 2
24 9 7 15 13 15 2 3 16 9 13 1 13 1 16 13 1 9 2 13 3 1 13 0 2
28 15 3 13 1 15 9 15 9 10 9 13 2 16 9 13 9 1 10 9 1 0 2 15 3 13 9 15 2
45 15 7 9 13 15 2 16 13 13 1 13 2 3 3 1 13 13 2 16 13 9 15 15 15 10 9 7 9 13 13 2 16 9 3 9 1 10 9 2 7 9 9 1 9 2
15 9 3 3 13 9 9 16 15 1 15 9 10 9 13 2
2 3 2
15 9 13 3 0 9 9 2 7 0 9 2 16 13 4 2
19 9 7 1 9 9 13 2 3 13 13 0 9 2 7 13 3 9 9 2
19 3 13 3 9 3 13 9 9 3 15 13 2 7 0 3 15 13 13 2
2 0 2
45 16 15 13 1 9 15 3 13 2 7 1 15 9 15 13 2 13 16 9 1 15 13 15 13 1 9 9 2 16 16 9 13 1 9 2 15 13 9 2 15 9 10 9 13 2
11 9 7 3 13 15 13 1 9 15 9 2
14 13 3 10 9 3 9 2 16 1 0 9 13 4 2
36 13 3 16 9 13 9 9 2 3 16 15 13 7 13 1 9 2 7 3 16 15 15 1 9 13 2 7 15 0 9 2 16 15 9 13 2
2 3 2
14 13 16 15 9 9 13 1 9 15 9 1 9 13 2
46 9 7 15 13 0 9 10 9 2 3 3 13 3 10 9 15 13 2 7 3 10 9 15 13 2 16 3 13 1 9 16 15 13 13 2 7 0 1 9 9 2 1 15 13 13 2
27 9 3 3 13 1 9 16 1 9 15 15 13 2 7 16 1 15 15 10 9 13 2 1 15 13 9 2
6 16 10 13 13 9 2
14 1 15 7 16 13 0 9 2 9 13 0 9 13 2
25 16 3 9 10 1 9 16 1 0 9 13 16 15 9 13 2 13 16 0 9 9 13 9 13 2
2 0 2
12 9 13 13 9 9 16 9 13 1 9 9 2
7 3 9 13 13 9 9 2
13 7 9 3 13 9 9 16 13 3 0 9 15 2
11 10 3 13 2 16 0 9 2 9 13 2
2 3 2
9 1 9 0 13 16 9 13 0 2
24 3 7 16 15 13 13 2 0 13 13 2 7 13 15 16 13 2 16 9 3 7 9 3 2
24 1 15 7 9 13 10 16 9 13 2 15 13 15 9 0 2 1 10 13 0 3 9 13 2
9 10 3 13 3 0 9 9 13 2
2 3 2
12 9 10 13 13 15 9 0 9 2 3 9 2
6 9 3 13 15 0 2
13 9 7 9 13 16 13 10 0 1 9 1 15 2
6 1 15 3 9 13 2
13 13 3 9 10 1 0 9 13 16 1 0 9 2
2 3 2
20 10 9 1 10 9 7 9 13 1 15 9 16 1 9 2 16 1 13 4 2
18 1 3 7 15 1 9 13 2 1 3 13 0 9 2 15 9 13 2
16 10 3 1 9 10 7 9 13 1 0 9 16 1 9 0 2
6 3 9 13 0 9 2
16 13 3 1 15 15 13 4 16 13 1 9 13 0 10 9 2
11 15 7 15 0 13 9 9 2 13 9 2
13 13 3 9 1 15 16 13 9 0 16 13 0 2
22 9 7 9 3 13 15 9 16 1 9 13 2 16 0 9 15 9 13 1 10 9 2
12 0 3 9 0 13 2 3 15 1 12 13 2
16 15 3 0 9 10 9 9 13 2 16 1 0 9 13 4 2
21 3 2 1 15 1 3 13 0 1 3 13 9 2 15 0 9 13 15 9 9 2
33 15 3 13 9 13 2 13 2 0 13 2 0 13 2 7 15 15 1 9 7 9 13 13 2 16 15 0 9 13 15 0 9 2
10 3 15 0 9 13 15 9 13 9 2
9 1 15 7 9 15 13 3 13 2
14 13 4 3 1 0 16 15 9 13 13 15 10 9 2
20 3 2 16 1 16 9 15 13 2 0 13 2 3 13 7 15 15 10 9 2
22 15 15 13 10 9 2 7 15 15 9 9 0 13 2 16 7 15 9 9 13 9 2
2 3 2
9 3 10 9 1 12 9 9 13 2
22 3 15 9 9 7 9 13 2 3 15 1 15 15 13 2 13 13 9 7 9 13 2
27 15 0 9 1 9 7 9 13 13 2 15 13 9 13 7 9 13 2 7 1 15 15 2 3 1 9 2
7 0 3 9 10 9 13 2
17 9 0 0 9 13 1 15 15 13 2 9 7 13 1 15 15 2
14 1 15 7 0 9 9 3 9 13 3 1 15 9 2
37 3 15 1 9 7 9 13 15 9 9 9 13 2 3 16 3 13 1 9 9 1 15 9 2 7 1 13 7 1 15 15 9 9 1 15 9 2
13 7 3 13 9 0 2 15 1 15 9 10 13 2
9 15 0 9 3 13 15 9 9 2
28 3 3 1 9 13 9 1 15 9 2 7 1 15 9 9 13 9 1 15 9 2 16 13 1 9 7 0 2
63 16 0 9 13 9 1 9 15 15 9 13 13 2 0 13 16 1 15 9 15 3 13 15 9 9 2 13 9 9 2 15 3 13 3 13 9 15 9 13 15 9 9 2 7 15 15 13 9 1 10 9 2 7 0 0 15 15 9 13 15 10 9 2
51 1 7 0 13 16 9 3 13 13 16 3 13 9 1 15 2 16 9 13 9 13 1 9 2 3 0 13 16 9 13 15 9 9 2 0 13 16 1 15 0 9 9 13 9 0 7 9 9 13 13 2
9 15 1 0 9 9 13 3 13 2
20 13 3 15 9 0 9 13 2 16 0 9 1 9 2 3 0 9 1 9 2
15 1 9 3 15 9 1 9 7 9 13 2 9 9 13 2
51 1 3 9 13 9 1 9 1 15 13 2 9 0 13 9 15 2 9 0 13 13 9 13 1 9 2 9 3 13 1 15 0 2 9 0 13 16 9 13 9 2 9 0 1 16 13 1 9 1 9 2
28 7 16 15 13 0 16 13 9 2 3 3 13 16 9 2 15 13 9 0 1 9 2 13 0 0 1 9 2
12 9 3 0 13 2 9 7 3 1 9 13 2
37 3 3 0 15 0 13 16 13 9 2 7 16 13 13 9 2 7 2 3 16 3 1 9 13 2 16 4 13 1 9 2 1 15 15 13 0 2
21 9 3 3 13 0 13 9 1 15 16 13 9 9 2 1 15 13 9 1 13 2
12 13 7 1 15 0 13 0 2 1 9 15 2
33 1 15 13 16 9 3 0 13 9 16 9 2 1 16 9 13 2 12 8 1 8 8 2 16 9 15 13 1 13 7 3 13 2
20 3 7 15 3 13 2 3 9 1 16 13 9 13 2 13 9 2 3 9 2
8 1 15 13 16 3 13 0 2
7 15 3 13 9 16 9 2
11 13 7 15 9 9 9 1 9 0 13 2
16 3 2 16 13 4 2 9 1 15 10 9 0 9 13 9 2
14 9 7 13 10 9 3 13 1 12 2 7 1 0 2
12 15 3 13 1 0 13 2 0 1 9 13 2
17 3 9 1 15 13 13 0 2 0 7 13 2 9 0 1 0 2
18 3 7 9 9 15 9 0 9 13 2 3 3 1 0 9 13 13 2
13 16 0 9 9 3 13 13 2 0 13 1 0 2
60 7 3 13 16 2 16 0 7 0 9 13 3 0 2 9 7 15 1 9 0 2 13 0 7 3 1 9 0 2 9 3 9 13 0 15 0 15 2 16 9 9 7 9 2 16 3 13 13 1 9 9 7 9 2 15 13 9 7 9 2
37 0 13 3 1 13 16 2 16 9 1 10 0 9 9 7 15 10 9 13 2 9 3 1 9 10 9 3 13 1 0 10 9 2 7 1 0 2
25 3 2 16 15 15 13 0 16 13 2 3 3 13 0 0 13 16 15 13 15 1 15 9 13 2
35 16 9 15 2 9 13 2 9 13 0 2 13 3 0 1 15 2 3 16 13 9 7 16 13 9 2 3 3 0 0 2 7 3 0 2
20 3 3 15 9 15 13 13 7 0 13 0 2 16 15 15 0 13 16 13 2
10 9 0 0 15 13 13 7 13 0 2
51 16 7 9 15 13 1 0 9 9 16 1 9 2 0 7 9 13 15 3 1 10 15 1 0 13 9 2 9 7 9 3 0 1 9 10 13 2 7 1 10 15 15 1 10 9 13 2 16 13 4 2
40 0 13 16 9 13 1 9 16 1 9 3 0 1 9 0 2 7 3 1 15 15 15 13 13 1 9 2 7 3 1 0 9 2 15 3 13 1 9 9 2
12 16 9 13 0 13 9 1 15 16 13 9 2
17 1 15 7 13 16 9 13 0 9 3 1 15 16 13 9 15 2
11 13 3 1 0 9 9 13 1 10 9 2
10 1 10 7 9 12 9 13 9 15 2
14 3 1 15 3 9 13 0 9 2 16 13 15 9 2
2 3 2
14 9 13 1 0 9 16 13 0 2 16 1 13 4 2
10 1 9 7 9 13 16 15 9 13 2
8 15 3 13 16 13 9 9 2
14 13 3 0 9 1 15 9 13 2 16 13 15 9 2
2 0 2
13 9 1 9 9 9 13 2 16 1 13 13 0 2
13 15 7 1 15 16 13 9 15 2 13 1 9 2
17 9 3 0 13 1 15 2 9 7 1 9 3 2 16 13 4 2
7 13 3 15 9 13 9 2
23 1 7 15 9 1 15 15 13 2 13 0 9 2 1 15 9 13 13 1 9 0 9 2
12 13 3 9 0 9 1 15 16 13 15 9 2
2 3 2
17 15 9 13 16 9 13 1 9 9 2 7 16 9 13 15 9 2
11 13 3 9 1 9 1 15 13 1 9 2
19 9 7 13 15 13 0 3 0 3 1 9 15 2 7 3 3 1 9 2
20 16 3 1 9 13 9 0 9 1 15 13 2 3 9 1 15 15 13 9 2
18 1 3 9 2 16 13 2 13 1 13 9 0 2 3 3 9 0 2
23 9 3 13 1 9 9 3 0 3 1 9 15 2 7 3 3 1 15 16 13 15 9 2
17 3 7 13 9 1 9 9 16 9 1 9 9 2 16 13 4 2
13 13 3 9 0 13 9 1 15 16 13 9 15 2
2 3 2
12 3 0 9 13 15 16 13 15 15 0 13 2
9 15 3 9 13 15 15 13 13 2
12 15 7 13 1 10 9 2 13 1 0 9 2
15 1 15 3 15 13 1 0 9 2 16 13 15 9 13 2
31 16 0 9 2 16 3 2 0 13 13 2 0 13 16 13 1 0 9 1 15 9 16 13 15 9 2 13 0 1 9 2
2 3 2
16 0 13 15 1 15 9 16 13 15 13 2 16 3 13 4 2
12 15 3 9 0 13 9 2 16 15 9 13 2
27 1 3 1 0 13 9 13 1 0 9 2 15 0 15 13 2 16 0 9 13 1 15 8 13 15 9 2
17 3 9 13 2 12 8 0 9 2 16 10 0 13 9 9 13 2
9 1 16 9 13 2 12 8 12 2
4 9 13 13 2
8 3 9 9 13 1 10 9 2
20 1 13 7 0 13 13 16 0 1 15 9 15 13 1 9 2 13 15 9 2
7 9 3 2 1 9 9 2
14 3 15 9 13 9 16 15 13 2 16 13 7 13 2
15 15 0 13 9 9 16 1 15 13 2 16 13 7 13 2
14 15 0 9 13 9 13 9 13 1 15 13 3 13 2
8 15 0 13 1 9 7 9 2
9 0 0 2 1 9 0 0 9 2
11 3 7 9 13 16 13 2 13 7 13 2
31 3 0 13 16 15 15 13 7 13 3 2 1 15 16 13 16 13 2 13 1 0 9 3 1 15 16 13 1 15 9 2
20 15 0 13 7 13 2 16 3 2 13 1 0 9 1 15 16 13 15 9 2
15 15 0 1 15 16 13 13 2 13 0 9 3 1 15 2
24 9 7 9 2 1 16 13 9 0 2 13 16 13 3 2 3 7 16 13 2 16 1 9 2
11 13 3 9 16 2 13 2 15 13 13 2
9 7 0 13 1 9 7 15 9 2
26 3 9 9 15 13 16 13 0 9 3 1 15 16 13 1 15 9 2 3 13 0 9 7 0 3 2
6 9 0 0 13 13 2
12 3 9 9 15 13 13 0 9 3 1 15 2
22 3 3 1 0 9 2 16 9 0 13 1 15 3 1 9 1 15 0 13 1 9 2
21 7 1 15 0 10 9 13 2 16 1 3 1 15 0 13 9 2 13 1 9 2
32 0 3 7 9 0 1 10 9 13 1 15 16 13 1 9 9 15 0 13 1 9 2 16 7 15 13 13 15 0 9 13 2
28 3 3 0 9 10 9 13 1 15 13 1 9 2 16 15 15 9 13 1 9 0 2 15 3 13 3 13 2
38 3 2 1 9 0 13 1 9 1 3 16 9 0 1 9 2 9 10 13 1 15 16 15 9 15 1 3 13 1 9 0 2 15 3 3 13 13 2
19 16 0 13 13 2 13 9 9 15 13 0 9 1 15 16 13 9 15 2
18 13 7 15 9 1 15 16 13 9 7 9 7 15 9 1 15 9 2
19 9 3 9 0 2 16 13 2 13 1 9 7 9 15 13 1 15 9 2
34 3 13 7 9 16 9 0 13 1 9 15 9 2 16 15 9 9 13 0 9 0 2 1 3 9 13 13 0 15 15 13 1 9 2
25 13 3 13 1 9 13 2 1 3 13 3 13 0 13 2 7 1 9 0 13 15 9 1 15 2
44 13 3 13 9 13 2 15 13 9 9 2 3 3 0 9 2 7 9 9 0 1 9 9 2 7 1 9 9 10 2 1 15 16 15 9 9 10 13 2 7 15 13 9 2
50 0 7 9 0 2 16 13 0 9 9 2 3 13 9 15 2 7 9 13 1 9 13 1 10 9 2 3 3 0 9 2 7 1 15 1 0 9 13 3 1 0 9 2 1 15 16 9 15 13 2
33 13 7 16 15 2 16 13 9 0 9 2 15 13 9 9 15 2 3 13 1 9 0 9 2 1 15 9 13 1 9 7 13 2
10 0 7 0 9 9 13 0 7 0 2
7 9 0 0 7 3 13 2
29 3 7 1 9 0 7 9 3 13 9 1 9 2 16 1 15 15 13 12 9 2 7 16 0 9 1 0 9 2
36 16 3 9 0 1 15 9 9 13 1 9 15 9 7 15 2 3 9 9 0 13 1 0 0 9 0 2 15 1 9 13 7 13 7 13 2
47 1 0 2 16 13 4 2 15 9 13 2 16 13 2 13 1 0 9 16 13 1 15 9 2 9 7 13 15 16 13 9 2 13 16 9 15 1 9 13 13 16 1 9 13 1 9 2
18 3 3 15 9 13 0 7 3 9 2 3 0 1 15 9 9 13 2
26 3 13 16 1 0 7 9 9 15 9 13 13 2 13 9 9 15 13 9 2 16 1 0 9 9 2
8 1 9 7 9 9 15 13 2
11 3 9 0 13 1 9 0 1 9 9 2
19 1 9 0 9 13 13 1 9 1 9 13 2 1 16 9 13 9 13 2
13 1 9 7 13 13 2 13 1 9 1 9 0 2
7 3 15 9 9 9 13 2
8 16 9 0 13 9 1 0 2
5 0 0 1 0 2
5 15 9 9 13 2
20 0 3 1 9 13 9 13 9 9 2 3 0 9 0 2 3 0 9 9 2
15 1 15 7 9 3 13 1 0 7 0 0 9 7 0 2
19 0 3 9 9 15 13 9 0 2 7 1 15 13 9 16 1 0 9 2
7 13 3 9 1 9 13 2
5 15 0 1 13 2
7 1 15 9 13 1 9 2
5 9 0 1 9 2
7 9 3 13 9 15 9 2
24 16 0 1 15 9 13 7 13 1 9 2 1 9 13 1 9 9 13 3 9 1 9 15 2
11 3 13 16 9 13 13 1 9 0 9 2
7 9 0 1 13 9 13 2
6 9 1 9 9 13 2
12 7 15 3 9 7 0 1 15 0 7 0 2
10 9 0 13 10 9 9 1 15 9 2
10 15 3 1 9 2 15 0 1 9 2
35 3 7 1 9 0 4 13 2 3 13 1 15 15 9 13 2 16 3 15 15 0 9 9 13 16 9 2 16 1 0 9 15 9 13 2
5 15 0 1 9 2
25 3 1 9 9 2 7 1 9 1 13 9 2 0 9 0 13 2 3 15 9 1 9 15 13 2
11 7 1 15 10 0 13 1 0 9 9 2
13 3 7 1 9 1 9 13 2 1 9 13 9 2
6 10 13 1 9 15 2
17 7 9 13 2 1 12 0 2 16 9 13 0 9 1 10 9 2
41 16 3 9 15 9 13 1 9 2 9 7 15 13 1 9 16 1 0 9 15 9 2 0 13 16 9 9 9 13 1 9 16 1 0 9 1 9 0 7 0 2
17 15 13 16 8 12 2 13 16 9 9 0 13 1 9 10 9 2
8 16 9 9 13 1 9 0 2
13 1 13 3 13 13 0 9 9 9 13 15 0 2
12 15 3 1 0 9 13 13 9 9 10 9 2
7 13 3 10 9 15 0 2
33 9 7 0 2 1 16 13 1 9 10 2 13 0 9 2 15 13 9 0 2 15 3 13 9 10 0 9 2 16 1 13 13 2
35 9 3 9 3 13 1 9 1 0 9 2 16 9 0 2 7 1 9 15 0 9 0 2 1 15 15 13 9 0 16 9 1 9 0 2
9 13 7 9 1 9 1 16 13 2
9 13 3 9 0 1 15 0 9 2
2 3 2
15 10 15 13 2 0 13 1 15 13 2 16 0 13 4 2
7 9 3 9 1 15 13 2
36 7 3 15 15 13 3 13 1 15 2 7 13 15 13 2 3 16 9 1 9 7 13 13 13 15 2 16 12 9 15 13 13 7 15 13 2
20 16 7 3 13 2 10 7 13 15 13 0 7 13 2 13 16 9 13 13 2
7 3 7 15 9 16 0 2
22 3 3 0 2 1 1 15 3 13 9 7 9 2 7 0 2 1 3 13 9 9 2
8 13 3 16 13 1 9 0 2
15 16 7 13 1 9 0 2 7 15 13 0 2 7 0 2
10 7 16 3 0 2 3 13 16 13 2
12 15 3 9 13 16 13 2 16 1 0 13 2
8 13 3 7 15 1 15 13 2
17 1 7 3 13 13 1 0 1 9 2 13 13 1 0 13 0 2
17 15 7 13 3 1 9 13 2 13 13 0 2 16 1 0 13 2
14 9 3 9 2 15 13 0 0 2 13 1 0 9 2
2 3 2
17 9 0 7 0 13 1 13 7 13 13 2 16 13 1 12 9 2
20 3 3 13 13 16 9 1 15 13 13 7 9 13 2 15 3 13 16 9 2
25 16 7 9 9 13 0 2 7 3 13 1 15 9 16 9 7 9 2 3 7 9 0 13 0 2
23 16 3 13 16 0 7 0 2 13 16 13 1 13 1 15 2 7 1 13 13 1 9 2
5 15 7 13 0 2
18 3 15 9 9 13 2 3 3 13 9 2 7 9 15 13 3 13 2
11 13 3 16 13 15 9 1 13 1 9 2
8 3 7 0 2 16 13 4 2
3 3 0 2
2 0 2
27 16 9 9 9 13 0 9 2 1 9 15 2 13 16 9 9 9 13 9 0 9 2 16 7 1 9 2
27 16 3 9 0 3 13 13 2 13 3 9 9 2 1 15 3 13 9 0 2 16 7 10 15 0 9 2
15 3 7 13 13 16 9 0 13 9 0 9 16 9 0 2
50 3 3 9 13 9 9 0 2 16 15 9 2 1 10 9 2 13 15 9 2 1 15 13 1 9 10 9 13 1 9 15 2 15 16 13 13 2 13 13 9 2 16 9 1 10 9 13 13 3 2
16 9 7 0 2 1 10 9 2 3 3 13 12 3 16 15 2
9 3 3 9 0 9 13 0 9 2
12 13 3 16 9 9 15 13 15 1 9 13 2
2 3 2
6 9 3 1 12 13 2
14 3 15 13 1 9 2 3 13 15 9 2 16 13 2
5 15 13 1 0 2
18 15 3 1 15 9 13 9 2 0 13 16 13 9 1 15 13 9 2
8 9 7 1 9 10 13 3 2
15 15 3 13 2 16 3 2 0 15 13 7 3 7 0 2
10 0 13 3 16 9 13 9 1 15 2
16 13 3 9 1 9 2 15 15 13 1 9 16 12 1 0 2
10 13 3 15 0 15 13 3 7 0 2
15 16 3 9 9 13 1 9 3 2 13 13 1 15 9 2
8 15 0 13 2 1 13 0 2
18 3 13 3 9 9 1 9 16 1 9 0 2 7 3 1 9 13 2
2 3 2
31 10 9 15 13 1 9 16 1 9 0 2 13 16 2 16 9 1 15 13 0 2 16 9 1 15 13 0 7 1 9 2
12 16 0 13 3 0 2 13 7 3 1 9 2
22 16 3 9 9 13 0 2 1 13 1 13 0 2 1 9 1 13 13 1 13 13 2
5 15 7 13 0 2
11 1 9 3 0 15 13 0 7 1 9 2
11 0 13 3 16 9 0 9 0 13 9 2
18 13 3 9 0 15 15 9 0 2 7 1 9 2 16 1 13 13 2
8 13 3 9 0 1 9 0 2
9 3 3 13 13 9 0 13 0 2
25 13 3 13 9 15 0 2 3 0 1 0 9 2 7 3 1 0 2 16 13 1 9 0 9 2
10 15 3 3 13 13 0 9 9 0 2
24 13 3 15 0 1 9 0 15 9 0 13 1 2 9 3 13 9 9 1 15 1 15 13 2
10 9 7 0 1 9 0 9 13 1 2
26 3 13 3 0 9 9 0 2 7 0 9 9 0 2 15 13 9 2 15 13 0 9 1 9 0 2
21 3 3 9 0 9 2 3 1 0 9 2 3 13 0 2 7 3 0 7 0 2
18 3 0 1 9 0 13 0 2 3 9 0 13 0 9 1 15 9 2
13 15 7 0 13 16 9 13 0 9 1 10 3 2
20 13 3 7 13 15 1 16 13 1 9 2 13 0 7 13 1 16 13 9 2
31 9 7 0 2 1 10 9 13 2 13 16 1 9 0 15 13 1 15 3 2 16 9 0 1 15 9 2 16 13 4 2
32 15 7 13 1 9 0 7 0 2 15 2 1 10 9 13 2 3 13 0 1 10 9 2 7 1 9 10 9 13 15 9 2
12 9 3 9 0 7 0 13 9 0 9 15 2
10 9 0 9 0 13 9 15 0 9 2
22 3 3 13 15 13 16 0 13 2 16 9 0 7 0 2 15 1 15 13 1 9 2
52 9 3 0 7 0 13 0 9 1 0 9 15 15 13 1 15 2 7 3 1 15 13 1 9 2 16 9 9 9 2 15 13 1 9 2 3 13 15 0 16 13 13 2 16 13 15 0 16 13 0 15 2
19 9 7 0 3 13 9 1 9 0 2 7 1 15 15 13 1 9 13 2
18 3 3 13 0 2 3 1 9 0 2 7 0 2 3 1 9 0 2
34 16 7 9 9 13 0 1 0 9 2 3 13 9 7 9 0 9 2 1 15 16 9 1 0 15 13 2 7 3 13 13 1 12 2
27 16 16 9 13 1 12 1 10 9 2 3 9 13 1 12 1 10 9 2 15 9 13 0 1 12 9 2
23 13 3 1 13 16 1 9 0 3 13 1 9 7 9 1 15 3 2 7 9 1 15 2
11 15 3 13 1 9 0 7 0 1 12 2
31 0 3 2 16 9 9 13 13 1 0 7 0 1 12 9 2 3 2 16 0 13 1 15 2 3 1 9 13 1 15 2
18 0 2 16 12 9 15 12 13 1 9 2 7 15 13 2 13 0 2
35 16 7 13 1 9 0 7 0 3 0 9 2 7 0 2 16 1 15 13 0 2 3 1 15 0 13 2 16 15 13 1 12 9 9 2
11 7 3 13 9 0 2 7 12 7 0 2
23 3 7 13 1 9 0 9 2 16 9 9 3 13 1 15 3 13 2 16 3 13 4 2
26 9 3 15 13 9 0 13 1 15 9 2 3 13 0 9 15 15 13 2 7 13 12 9 7 0 2
18 3 15 3 1 9 9 13 16 0 2 7 3 16 0 1 9 13 2
47 3 13 7 2 3 1 0 9 2 3 9 0 13 1 9 0 13 2 15 13 9 15 2 7 1 9 13 2 7 3 15 9 0 13 1 9 0 2 7 15 2 7 13 9 0 13 2
23 7 0 3 0 1 9 2 15 0 13 9 13 2 16 13 16 9 0 13 1 9 0 2
8 3 13 9 3 15 9 13 2
37 16 7 9 0 1 9 0 13 2 16 13 4 2 9 7 9 0 13 1 9 1 9 2 0 13 16 9 7 9 15 9 13 1 9 9 13 2
11 1 15 3 13 9 0 9 2 7 9 2
16 9 7 13 9 9 9 1 10 9 2 15 13 1 9 0 2
9 13 3 16 13 16 9 0 9 2
26 4 3 9 7 9 9 9 1 9 0 13 7 13 16 1 0 9 2 1 9 0 0 16 1 9 2
33 13 7 16 9 15 15 13 7 13 1 0 9 2 13 1 9 15 2 16 9 9 13 1 9 9 2 7 1 15 13 1 9 2
27 10 3 9 15 13 1 15 9 2 7 10 9 2 13 1 9 0 15 13 1 9 15 9 2 7 15 2
26 7 1 15 13 9 2 1 9 1 8 2 16 9 15 13 1 9 2 13 1 9 15 13 1 9 2
33 7 3 1 15 13 9 9 2 16 9 13 13 9 9 15 13 1 9 2 16 9 13 15 1 15 0 2 7 13 0 9 0 2
16 15 0 13 15 1 9 13 2 7 13 9 9 1 9 9 2
67 16 0 10 15 13 1 15 1 15 2 3 1 9 2 13 1 15 1 9 10 9 2 9 7 0 13 1 9 0 2 9 7 0 13 1 10 9 10 9 1 15 9 2 0 13 16 9 0 13 1 9 10 9 1 9 0 2 7 1 13 10 9 9 1 0 9 2
17 3 3 3 13 0 13 15 0 9 9 9 13 7 13 1 9 2
23 13 3 1 9 16 13 1 9 1 9 13 2 1 9 15 9 13 1 9 13 1 13 2
34 16 3 9 13 9 1 9 13 1 9 13 2 3 9 0 13 9 1 9 0 1 13 0 2 1 15 13 10 9 7 9 7 9 2
12 3 3 13 16 15 9 9 13 9 9 13 2
16 3 9 0 13 0 13 13 1 9 2 16 9 1 15 13 2
15 7 1 15 9 9 13 13 13 1 9 2 16 9 0 2
30 0 3 13 16 15 3 15 9 13 2 13 13 1 9 2 7 13 9 0 9 2 7 13 0 9 2 7 0 9 2
10 3 13 7 9 7 15 7 15 13 2
24 3 1 15 16 13 1 10 9 2 13 1 9 2 1 15 1 3 0 13 1 3 13 9 2
15 1 0 16 13 1 15 16 13 0 2 13 1 0 9 2
8 9 3 13 15 16 0 13 2
16 9 7 15 7 15 0 13 16 13 0 16 13 9 0 9 2
19 1 15 3 13 1 0 9 2 16 13 1 0 9 2 7 3 1 13 2
11 3 13 16 10 13 0 9 3 0 9 2
9 9 7 10 15 9 13 13 0 2
12 12 3 9 2 1 16 13 15 0 9 9 2
15 7 3 13 9 10 0 1 13 9 2 15 1 13 13 2
10 15 9 2 1 16 13 15 9 9 2
26 7 3 13 0 9 9 16 13 9 9 7 15 9 2 7 15 15 13 1 9 7 9 9 10 9 2
7 0 0 9 2 9 9 2
13 7 3 13 0 9 1 13 9 0 2 16 9 2
12 0 7 9 2 9 9 9 13 1 10 9 2
17 7 3 9 2 15 13 1 9 2 1 10 9 10 9 13 9 2
33 1 15 13 16 3 15 13 9 9 2 7 13 1 9 9 2 3 9 9 0 13 2 7 3 1 13 1 15 9 13 7 13 2
9 3 0 1 0 9 0 9 13 2
6 9 0 1 9 9 2
6 9 0 1 9 9 2
14 9 7 2 15 13 9 1 9 2 1 9 15 9 2
28 3 3 0 13 1 15 16 9 2 16 3 2 13 0 2 16 3 15 13 0 2 3 1 13 9 10 13 2
42 7 16 1 15 9 15 13 9 13 0 7 9 10 15 13 15 9 2 13 16 9 2 15 13 1 9 9 7 10 9 0 13 2 1 10 9 13 0 10 9 13 2
12 16 7 15 9 13 1 15 2 13 15 9 2
25 15 3 13 16 15 13 1 15 16 13 15 9 2 13 1 0 9 2 7 3 13 1 10 9 2
30 3 13 3 9 16 9 9 0 2 7 9 9 15 2 13 13 0 1 15 9 15 13 7 13 2 15 13 15 0 2
27 3 3 13 1 15 16 1 0 9 2 7 2 13 15 9 2 13 10 9 2 7 0 9 16 0 9 2
9 16 13 9 13 9 10 0 9 2
30 1 7 10 9 2 3 9 13 2 13 1 9 16 1 9 0 2 1 15 7 9 13 10 16 1 9 15 15 13 2
16 0 9 15 0 9 1 15 13 2 3 1 0 9 13 15 2
13 3 13 16 15 13 9 0 9 2 3 13 9 2
12 0 3 9 15 9 13 9 2 16 13 4 2
14 13 3 15 16 0 9 9 13 3 3 15 0 13 2
33 0 7 13 15 9 1 15 16 1 15 9 15 15 9 13 2 15 13 16 15 15 13 1 0 9 2 16 16 13 15 15 9 2
12 9 3 0 13 1 0 9 16 1 0 9 2
2 3 2
8 0 9 15 9 13 9 15 2
6 13 3 0 9 15 2
14 3 15 1 0 9 3 15 13 2 13 0 7 0 2
8 13 7 13 0 9 9 0 2
6 15 3 13 9 15 2
13 15 3 13 9 1 15 9 2 15 13 0 9 2
17 7 0 1 9 15 3 13 1 15 13 2 16 13 13 7 13 2
29 1 7 3 9 1 9 9 13 2 1 15 3 13 2 13 16 3 13 9 15 15 9 2 3 15 9 13 9 2
20 7 3 13 9 0 2 15 9 13 2 13 9 1 9 15 9 15 13 13 2
11 13 3 9 13 13 0 9 15 0 9 2
15 13 7 15 13 0 3 9 0 9 13 1 13 0 0 2
33 3 3 15 15 13 0 0 15 7 15 0 9 2 13 0 0 0 2 7 3 15 0 9 13 9 2 3 10 0 0 13 9 2
25 7 3 9 0 0 9 13 13 1 0 0 15 15 13 0 0 2 3 15 9 13 1 13 9 2
22 15 0 9 9 0 9 13 13 15 9 0 2 15 13 3 9 15 15 1 15 13 2
17 7 0 9 0 13 16 3 13 13 0 0 0 2 1 15 9 2
16 13 3 15 1 13 15 15 13 0 0 16 9 9 1 9 2
16 7 0 13 16 9 15 9 0 2 3 9 2 13 13 9 2
16 13 4 3 1 16 10 9 0 9 1 15 13 2 13 9 2
19 9 7 0 2 16 13 9 1 9 0 9 2 13 3 0 10 9 13 2
17 1 3 0 9 3 13 0 9 2 13 3 9 0 9 15 9 2
17 15 7 13 13 10 9 0 1 15 16 15 13 2 16 13 4 2
11 13 3 13 9 0 1 9 16 1 9 2
2 3 2
26 16 9 9 13 13 1 9 16 1 9 1 9 9 2 3 9 0 1 9 9 2 16 1 13 13 2
41 9 7 9 13 2 16 13 1 9 0 9 2 3 3 3 13 9 9 2 7 13 1 9 9 1 0 9 2 16 1 13 13 2 16 0 1 15 9 13 13 2
24 9 3 15 0 13 1 0 9 13 2 15 13 15 1 0 9 2 3 16 9 9 9 0 2
2 0 2
7 15 0 13 10 9 0 2
33 9 7 0 3 13 2 7 13 2 7 13 1 9 0 2 16 0 3 1 15 13 13 2 16 1 9 9 15 13 1 9 9 2
10 13 3 0 9 9 13 15 9 9 2
2 3 2
10 15 13 1 0 9 16 1 0 9 2
14 15 3 1 15 15 0 9 13 2 13 0 9 15 2
12 9 7 13 0 9 0 1 15 16 0 13 2
14 15 3 9 13 1 10 9 2 7 15 13 10 15 2
35 1 9 7 15 9 3 13 9 1 16 13 9 2 16 1 16 13 1 9 7 9 2 16 9 3 9 13 13 2 16 1 0 13 4 2
16 7 1 15 16 13 9 2 0 13 9 1 16 13 15 9 2
15 3 15 9 13 15 13 10 15 2 16 1 0 13 4 2
10 13 3 9 13 0 9 10 0 9 2
2 3 2
17 15 13 3 1 15 0 2 13 1 15 15 13 3 1 15 0 2
22 3 3 13 13 1 0 1 9 9 2 16 9 9 13 2 1 3 13 0 13 0 2
14 10 7 9 7 9 7 9 0 13 3 1 15 0 2
11 3 1 15 9 3 13 13 2 7 13 2
8 9 7 0 13 1 15 0 2
7 3 9 15 13 15 13 2
18 7 13 15 9 1 9 0 15 3 13 1 15 9 2 16 9 0 2
33 3 3 15 9 0 2 15 13 1 9 13 2 13 15 9 13 2 3 16 1 15 3 9 13 2 3 13 3 13 1 0 9 2
15 15 13 3 13 2 16 9 1 15 13 2 15 13 9 2
20 13 3 9 0 1 0 2 7 0 10 0 9 1 9 9 2 16 1 9 2
42 1 10 7 9 7 9 13 1 15 13 13 0 9 15 13 0 7 0 15 2 16 9 0 2 1 15 13 9 9 2 15 13 9 15 2 13 0 7 0 9 0 2
32 15 7 9 15 13 9 0 1 15 9 0 2 3 1 15 10 15 13 2 3 1 15 13 10 9 2 7 9 1 13 9 2
20 15 7 0 9 15 13 1 9 9 16 1 0 9 2 3 7 9 0 13 2
12 13 3 9 0 9 0 10 0 9 7 9 2
2 3 2
29 1 10 9 7 13 13 13 16 9 0 9 7 9 13 0 9 10 2 16 9 9 9 13 9 10 1 15 13 2
11 1 10 7 9 9 2 9 13 0 9 2
10 3 9 13 9 2 13 15 10 9 2
28 9 7 0 2 15 13 9 2 13 9 0 2 15 13 0 7 0 2 3 7 9 3 13 16 9 9 13 2
12 9 7 0 2 13 9 9 2 13 3 9 2
9 9 3 9 13 9 10 9 0 2
16 9 7 7 9 9 13 0 2 7 1 13 0 9 0 0 2
22 13 3 0 9 15 9 2 7 10 9 7 9 15 2 13 0 0 2 15 13 9 2
2 0 2
11 0 13 10 9 9 13 9 15 15 13 2
21 3 1 9 15 15 13 2 15 9 13 2 9 0 13 13 2 13 7 9 13 2
9 7 13 9 16 13 1 0 9 2
11 7 3 9 15 13 13 16 0 9 13 2
11 13 3 9 0 13 0 9 3 0 9 2
7 0 7 10 9 9 13 2
8 13 3 0 9 9 13 9 2
2 3 2
9 15 9 13 0 9 13 9 13 2
7 9 7 0 13 9 0 2
18 13 3 0 13 9 15 2 15 0 9 13 2 16 1 0 13 4 2
12 3 4 7 15 13 9 0 16 0 9 13 2
29 3 13 3 1 9 0 2 15 13 0 9 2 15 0 9 2 16 0 9 13 2 15 13 0 9 16 0 9 2
9 13 3 0 9 9 15 9 9 2
2 0 2
21 9 2 15 0 9 13 1 10 3 2 3 0 7 0 13 2 3 3 13 9 2
26 3 13 9 1 12 1 9 2 16 9 0 13 3 13 13 1 0 2 16 3 3 13 3 16 0 2
21 15 3 0 1 15 13 1 16 0 2 3 13 1 0 2 7 1 15 13 13 2
7 15 7 13 1 9 13 2
12 3 3 15 0 13 2 3 0 9 13 13 2
12 13 3 9 0 9 1 13 1 15 13 9 2
14 15 7 3 13 13 15 16 0 0 2 15 9 13 2
8 13 3 9 0 9 0 9 2
15 0 7 9 9 2 7 15 0 9 2 9 7 9 13 2
17 15 3 13 15 10 9 0 13 16 0 9 2 7 1 15 3 2
12 13 3 9 7 9 0 15 9 0 13 9 2
7 15 13 15 13 8 12 2
9 0 9 9 2 16 15 9 13 2
4 7 8 12 2
12 15 13 9 0 2 16 13 15 2 9 0 2
24 15 3 9 9 1 0 9 2 13 2 16 0 9 9 13 13 0 2 3 1 9 0 0 2
7 3 9 13 1 9 9 2
62 16 0 0 9 10 9 13 1 9 3 0 13 2 7 3 1 9 9 2 13 7 13 15 7 1 15 9 13 2 13 15 13 16 0 9 2 7 0 9 9 2 3 13 1 13 9 2 7 3 1 13 2 7 15 15 9 9 15 13 1 15 2
31 0 1 9 9 13 9 2 15 13 9 9 2 0 7 2 15 13 9 9 2 3 13 9 9 16 16 7 15 13 9 2
17 3 3 13 9 13 0 9 1 9 9 2 7 3 1 9 9 2
2 3 2
20 0 9 9 13 9 2 15 13 9 16 9 9 2 16 1 12 8 9 13 2
20 16 3 9 9 13 0 9 2 13 16 0 9 3 13 1 9 9 16 9 2
2 3 2
11 9 13 3 1 15 13 16 3 1 15 2
10 0 3 13 13 1 15 3 13 13 2
13 15 7 13 9 0 9 2 16 3 1 15 13 2
14 13 3 0 9 3 1 9 9 16 9 2 16 13 2
2 3 2
12 1 9 0 9 0 10 13 2 1 13 0 2
7 0 7 13 9 16 9 2
9 3 3 13 13 9 9 16 9 2
2 0 2
8 9 13 13 9 9 16 9 2
8 3 9 13 9 1 10 9 2
12 9 3 9 13 15 9 13 2 1 15 13 2
9 9 3 9 13 0 16 9 9 2
19 3 3 13 0 9 2 15 13 9 2 13 1 9 9 16 1 9 9 2
7 15 7 13 0 0 13 2
21 1 3 9 13 0 9 0 9 2 13 16 1 15 0 9 13 15 13 15 0 2
19 9 7 3 13 0 0 9 2 7 10 9 13 2 16 13 9 1 0 2
14 15 3 9 13 1 15 16 9 9 15 13 1 9 2
11 15 3 3 9 13 2 13 9 0 3 2
18 15 0 13 9 0 2 7 9 0 13 2 1 15 0 7 0 13 2
15 15 0 13 9 0 2 7 9 9 0 13 2 3 9 2
22 9 3 2 1 16 13 9 2 3 13 0 0 9 2 7 0 1 16 1 9 13 2
9 9 7 1 15 0 13 0 9 2
18 9 3 7 9 1 9 9 13 0 7 0 2 3 16 1 9 9 2
2 3 2
27 1 10 9 15 13 1 10 9 2 9 13 0 0 9 15 9 2 16 9 0 0 13 16 13 15 0 2
6 15 7 9 13 9 2
5 0 3 13 9 2
10 9 3 9 13 0 0 16 9 15 2
9 0 3 15 9 13 10 9 15 2
9 3 13 3 9 9 0 13 13 2
10 15 7 13 0 9 2 15 13 9 2
12 0 13 3 16 9 7 9 13 15 9 9 2
2 3 2
28 1 10 9 15 13 13 1 10 9 2 0 13 16 9 15 9 13 1 9 15 2 7 3 13 1 10 9 2
22 16 3 9 13 15 13 2 0 13 13 16 13 9 15 2 7 13 16 13 15 13 2
11 3 15 13 15 9 13 2 15 9 13 2
28 3 13 16 7 13 1 0 2 7 2 16 13 13 1 0 13 2 15 3 13 15 13 2 7 15 9 0 2
15 0 13 16 0 13 3 13 15 13 2 7 15 15 0 2
11 0 7 13 0 9 13 15 9 7 9 2
7 3 1 15 13 15 13 2
10 0 13 3 9 0 1 9 9 13 2
2 0 2
13 15 1 15 15 13 9 15 2 13 9 10 9 2
13 13 3 0 9 1 13 1 15 15 9 9 13 2
11 0 7 9 3 13 1 0 1 9 9 2
28 3 15 9 15 13 9 1 13 7 13 7 13 2 15 13 15 15 15 13 16 0 9 2 7 0 7 0 2
19 3 7 0 13 0 9 15 16 15 13 7 0 2 15 13 1 9 9 2
16 9 3 2 7 9 2 1 9 0 3 16 1 9 9 13 2
2 3 2
20 16 15 9 9 13 15 9 2 15 9 13 7 13 2 7 13 2 7 13 2
9 0 13 7 16 13 13 0 9 2
13 13 3 9 1 16 9 13 1 15 15 3 13 2
7 15 7 13 9 0 9 2
8 13 3 3 13 13 0 9 2
24 13 3 9 3 0 16 13 2 7 3 16 3 13 2 1 9 16 13 16 3 13 9 13 2
17 7 16 9 3 13 9 13 2 15 13 1 15 16 9 13 13 2
23 15 3 13 13 9 15 13 9 2 16 13 2 15 1 13 13 0 2 1 13 0 9 2
8 0 7 7 9 13 0 9 2
28 15 3 13 9 9 13 9 2 7 16 9 3 13 13 2 7 16 0 13 13 2 7 16 1 13 13 13 2
7 3 13 3 9 0 9 2
10 15 3 9 9 13 13 0 15 9 2
2 3 2
12 16 9 13 0 9 2 15 1 15 13 13 2
5 15 7 13 0 2
12 13 3 15 9 13 1 15 1 15 13 9 2
22 3 9 15 13 0 7 13 9 2 0 13 7 13 2 15 7 0 2 0 7 13 2
10 13 3 16 13 0 7 13 1 15 2
11 3 13 3 15 0 9 2 15 13 9 2
2 3 2
8 13 9 9 13 1 9 9 2
10 3 9 0 13 1 10 9 1 9 2
13 1 0 7 13 9 1 9 2 7 3 1 13 2
39 13 3 16 9 15 9 9 9 13 15 13 0 1 9 0 13 2 16 1 9 9 2 15 13 1 9 9 2 7 1 9 0 2 15 13 1 9 9 2
12 16 3 13 9 2 9 1 13 9 0 13 2
9 0 3 13 16 9 13 0 9 2
2 3 2
23 9 15 15 13 13 16 9 9 1 15 9 13 2 16 9 13 9 9 1 15 9 13 2
30 16 7 9 1 9 13 1 9 7 13 1 15 2 3 9 0 13 9 0 1 9 0 2 15 3 13 9 3 13 2
24 0 7 13 13 16 9 9 9 0 3 13 13 1 9 0 2 7 9 9 15 1 15 13 2
14 16 3 15 0 9 13 16 9 13 2 3 13 15 2
11 13 7 15 16 1 15 13 1 9 0 2
10 15 13 2 3 9 2 13 9 9 2
12 7 3 9 15 3 13 9 2 7 13 9 2
11 7 3 9 13 9 0 2 7 13 15 2
10 0 3 3 7 15 9 9 13 9 2
2 3 2
43 16 15 9 13 15 9 0 9 2 15 15 9 13 3 9 0 1 15 0 13 9 15 2 16 15 15 9 13 9 2 13 3 13 9 9 2 3 7 13 2 7 13 2
8 9 7 0 9 0 13 9 2
18 15 3 9 9 13 0 15 9 7 9 2 1 15 0 13 1 9 2
5 15 7 13 13 2
8 3 13 3 13 15 3 13 2
17 13 3 0 9 9 1 13 9 1 9 0 2 3 1 9 9 2
14 3 3 1 15 15 13 4 2 13 9 1 0 13 2
33 3 3 2 16 9 1 15 16 13 9 0 9 2 13 9 9 2 1 15 0 13 16 13 0 15 9 9 2 16 0 9 13 2
21 3 1 15 15 16 13 0 9 2 13 16 3 13 9 15 2 16 1 13 13 2
22 7 3 13 16 10 15 15 9 15 9 13 2 13 9 15 9 2 16 0 9 13 2
7 13 3 15 9 15 0 2
8 0 9 2 16 13 3 9 2
8 15 9 2 16 1 9 13 2
20 16 9 9 1 16 3 13 9 2 13 15 1 15 9 9 13 2 3 9 2
8 3 3 9 13 16 1 15 2
15 3 7 1 9 9 13 15 13 2 16 13 9 13 9 2
54 9 0 1 9 9 2 13 3 15 15 13 1 9 13 2 16 9 0 15 2 16 15 15 13 1 9 9 2 16 9 2 15 13 1 9 9 2 7 3 15 15 13 1 15 16 9 9 13 13 2 16 9 9 2
22 15 3 15 13 9 9 1 16 3 13 9 2 13 9 15 2 16 9 13 9 9 2
17 7 0 0 9 15 9 2 15 13 3 9 15 2 13 9 15 2
13 15 7 13 9 9 1 9 2 3 13 9 9 2
6 3 9 13 9 15 2
8 9 3 7 9 13 1 9 2
17 16 3 9 13 9 9 2 3 3 13 9 3 13 7 9 13 2
10 3 1 15 13 9 16 9 13 0 2
28 0 13 9 1 10 9 2 16 9 7 9 0 2 16 13 9 2 3 3 13 9 9 2 7 3 1 13 2
54 15 3 15 13 9 1 0 9 9 13 2 7 1 13 9 13 13 2 3 13 9 9 2 7 3 1 13 2 16 9 9 2 7 9 9 2 7 15 3 2 1 15 13 9 2 1 12 9 2 16 0 13 9 2
43 9 7 13 9 9 2 3 3 16 1 15 13 9 1 10 9 2 7 13 1 15 9 2 16 9 13 1 10 9 1 9 9 2 7 13 0 9 15 13 1 9 9 2
12 3 1 9 13 7 13 9 13 1 15 13 2
28 3 1 12 9 9 13 16 9 13 9 16 9 9 2 15 3 13 1 15 15 13 9 2 7 3 1 13 2
27 7 7 16 9 3 1 15 13 9 7 1 15 2 13 0 9 16 9 13 0 9 2 16 0 9 13 2
22 3 9 2 16 3 13 0 9 2 13 3 0 9 13 2 1 1 9 9 9 13 2
13 3 7 0 13 9 15 13 1 13 2 16 9 2
20 15 3 0 9 9 13 2 16 13 9 9 0 2 1 15 9 10 13 4 2
12 1 2 9 13 16 0 9 9 13 3 13 2
21 15 7 13 1 0 2 16 9 0 3 13 13 9 2 13 2 16 0 13 9 2
32 7 15 15 13 1 9 2 15 13 13 9 7 13 15 2 7 15 13 15 3 13 9 9 2 16 9 9 13 1 9 0 2
21 3 3 13 1 9 9 2 16 1 9 13 9 2 15 13 2 13 9 10 9 2
11 7 3 9 15 13 0 2 13 0 9 2
15 0 3 13 1 12 9 0 2 1 1 10 9 13 9 2
26 7 16 9 13 9 3 2 3 13 12 9 2 3 1 12 9 15 13 2 7 1 9 10 9 13 2
26 7 1 15 9 9 0 7 0 13 12 2 3 0 16 9 13 1 9 9 2 7 3 0 1 9 2
26 7 3 13 16 15 3 13 9 9 3 0 2 1 1 9 10 13 9 0 2 3 0 2 7 0 2
37 3 15 13 0 9 9 2 3 3 3 1 15 15 13 1 9 10 2 3 1 9 0 2 7 3 3 1 15 15 13 1 9 10 2 3 9 2
52 9 3 10 3 13 12 9 0 9 9 13 2 3 16 1 9 9 13 2 1 15 13 0 9 9 1 0 9 2 7 16 15 15 1 9 13 12 7 0 2 13 1 9 10 2 3 16 0 1 9 13 2
13 7 9 13 3 12 9 0 2 3 9 7 9 2
29 9 7 9 3 3 13 1 10 9 2 15 0 13 2 16 13 1 9 7 9 2 15 15 13 1 15 9 9 2
22 13 3 9 9 1 9 9 2 7 13 9 15 9 7 13 9 7 9 7 0 3 2
44 3 13 15 13 2 16 1 9 13 15 9 9 7 9 7 15 15 13 1 9 2 7 1 0 13 15 9 9 2 7 1 0 13 15 9 15 9 1 15 15 13 1 9 2
18 13 3 9 1 15 10 9 2 13 1 9 2 13 1 9 1 15 2
33 7 3 0 13 15 2 9 2 9 7 9 2 3 16 9 13 1 9 13 1 9 9 2 9 1 9 2 9 1 9 1 15 2
40 7 3 0 13 15 2 12 2 0 7 9 2 16 9 9 13 1 10 9 16 1 9 13 4 2 7 9 1 16 13 9 2 7 9 1 16 13 1 9 2
26 3 3 13 13 1 9 15 9 1 16 13 3 9 1 9 2 7 1 0 9 2 7 1 9 9 2
15 7 15 13 15 16 13 9 0 7 0 0 2 3 9 2
12 7 9 13 9 13 2 1 13 9 0 9 2
9 3 2 9 0 0 13 16 0 2
11 7 9 0 13 9 10 1 15 9 0 2
14 7 16 1 9 13 9 0 2 3 1 9 9 0 2
9 3 3 9 0 13 10 9 0 2
20 3 7 3 1 9 2 16 9 2 1 13 9 0 2 13 12 9 15 9 2
37 7 3 13 16 0 9 9 13 9 2 16 13 1 9 16 9 0 9 15 9 13 2 16 13 9 0 7 0 2 15 13 3 9 7 9 15 2
26 1 0 13 2 16 9 0 13 9 15 2 1 15 13 9 2 15 13 9 13 15 2 16 9 0 2
18 9 7 0 3 13 15 9 13 9 2 16 13 4 2 1 8 8 2
31 1 0 13 2 16 16 1 9 0 13 9 7 9 9 1 9 2 3 9 3 13 10 9 2 16 9 9 3 13 9 2
30 16 13 2 16 9 13 1 9 9 9 2 7 3 9 9 2 1 15 13 2 16 9 13 9 9 2 7 9 15 2
12 3 10 9 2 3 13 1 15 2 0 13 2
42 3 1 13 2 9 13 9 15 3 13 9 9 2 1 9 2 15 13 0 2 1 9 13 9 9 2 15 1 9 13 2 3 3 3 1 9 2 7 3 1 9 2
39 13 13 2 16 9 1 9 13 15 9 2 15 16 15 2 1 13 9 2 13 9 10 1 9 15 13 2 1 13 9 2 7 3 13 9 1 9 9 2
31 16 7 13 9 0 2 13 9 9 2 1 9 9 15 9 2 1 9 2 0 0 2 13 9 7 9 1 9 10 9 2
21 1 0 13 2 16 16 12 9 13 1 9 2 9 13 13 3 9 15 15 13 2
18 13 9 15 3 13 9 9 2 9 3 13 9 9 7 9 1 9 2
6 9 3 13 9 9 2
9 7 9 13 9 9 2 7 9 2
31 7 0 13 16 3 1 9 13 0 13 1 9 9 1 15 13 9 2 16 1 15 13 9 2 1 9 15 13 9 9 2
20 7 9 13 1 9 9 2 1 15 9 13 2 13 9 0 2 7 9 0 2
19 7 3 9 13 1 15 9 12 2 13 1 9 9 2 7 3 1 9 2
16 7 15 9 9 13 1 0 9 2 15 13 9 13 1 9 2
31 1 0 13 2 16 1 13 9 13 9 2 13 0 9 1 15 16 9 9 13 13 3 0 2 16 13 9 10 1 9 2
16 16 9 2 3 0 13 2 16 3 9 13 9 10 1 9 2
14 3 9 13 13 2 16 3 3 1 15 13 9 9 2
58 3 3 13 1 9 1 9 2 16 1 9 13 15 15 13 9 7 13 15 0 1 9 9 2 16 13 13 1 9 7 1 15 9 13 2 7 0 9 13 2 15 13 1 9 9 1 10 9 7 3 1 10 9 2 16 13 9 2
31 3 2 10 15 13 9 9 2 4 13 1 15 7 1 9 2 1 15 2 16 15 9 13 2 1 9 2 16 9 15 2
21 13 3 9 9 1 15 13 9 2 7 15 9 9 7 9 9 13 9 9 13 2
11 7 15 9 9 13 13 9 1 9 13 2
65 13 3 13 9 2 16 2 1 1 10 9 0 13 15 13 9 9 7 15 1 9 13 2 16 1 9 9 9 9 13 9 2 7 15 13 1 9 13 2 16 3 1 9 15 2 2 3 13 16 2 1 9 0 13 9 9 0 2 1 9 13 13 9 0 2
56 0 7 0 13 15 13 0 1 15 15 1 9 10 13 2 7 15 13 10 9 2 16 1 0 2 7 2 16 1 9 2 15 9 13 9 2 16 13 2 9 13 13 0 2 7 9 2 16 13 2 9 13 0 13 0 2
19 3 2 10 9 0 15 9 13 1 9 0 15 2 16 13 1 9 9 2
8 3 9 15 13 0 9 9 2
14 3 15 9 13 7 9 0 2 7 0 9 15 9 2
20 0 7 7 9 13 9 15 2 7 9 9 1 9 2 0 9 1 9 0 2
23 13 3 0 9 13 2 1 15 16 13 9 9 15 13 2 7 3 13 0 9 1 15 2
16 9 3 0 9 13 3 1 15 15 13 9 9 10 9 0 2
32 7 9 9 13 3 1 15 15 3 13 9 2 16 3 0 13 7 13 1 9 3 13 9 9 2 16 13 1 9 1 15 2
36 9 3 13 1 15 1 9 15 2 7 3 13 2 16 7 15 15 9 2 15 1 15 0 13 2 7 1 16 13 1 15 2 13 1 15 2
11 7 9 0 3 13 13 9 16 13 8 2
25 13 3 15 9 7 9 9 1 9 10 9 2 3 9 2 13 9 2 7 15 15 13 9 9 2
25 1 0 3 13 2 16 9 13 3 15 9 15 13 1 9 9 0 7 0 15 9 3 13 0 2
17 9 7 3 13 9 9 2 1 3 13 1 15 2 7 1 15 2
11 7 3 9 2 15 13 9 2 0 13 2
18 7 3 9 3 13 1 15 2 7 3 1 9 2 16 13 1 9 2
25 3 3 13 3 9 1 16 13 9 15 9 2 7 16 13 9 13 15 2 16 9 13 9 9 2
12 9 3 13 9 13 2 0 7 0 9 13 2
5 7 9 13 9 2
27 13 3 15 9 15 3 13 9 1 15 2 7 3 1 15 2 16 9 0 2 16 9 15 2 16 0 2
39 7 9 15 13 1 12 2 7 16 13 0 1 9 7 1 9 2 16 9 0 2 7 9 2 7 0 2 7 16 13 0 15 2 15 0 9 3 13 2
10 16 3 13 9 2 9 13 9 9 2
12 7 3 13 2 16 9 7 13 9 7 9 2
6 3 3 13 9 0 2
11 3 9 9 3 13 9 16 13 12 8 2
6 3 3 13 9 0 2
19 3 2 15 9 0 13 1 15 3 13 2 1 10 9 13 1 15 0 2
14 16 3 9 13 9 0 2 3 13 1 15 3 13 2
29 15 3 13 2 16 9 13 13 1 9 7 9 2 15 3 13 15 13 2 15 13 9 9 7 15 0 7 0 2
25 7 15 3 13 13 0 2 16 15 9 13 0 2 16 1 15 16 13 1 9 7 1 9 9 2
22 15 7 3 13 16 13 9 0 9 9 2 1 15 9 9 13 0 1 9 1 9 2
35 7 3 9 0 2 16 13 0 1 10 9 2 3 13 15 9 2 7 13 0 1 15 9 1 9 9 0 2 1 9 0 3 13 0 2
10 3 13 16 0 9 0 13 15 9 2
20 7 0 9 15 13 1 9 2 13 9 2 1 15 3 13 2 16 13 8 2
17 3 9 9 13 1 15 9 2 7 3 9 3 13 16 1 9 2
39 16 3 13 2 16 9 9 13 0 9 13 1 9 2 3 13 1 15 2 16 1 9 9 9 3 13 9 2 7 1 9 2 15 13 9 9 1 9 2
18 7 3 1 9 9 2 1 16 13 0 9 2 13 1 15 0 9 2
13 9 7 3 13 9 2 7 9 1 9 7 9 2
23 3 1 10 15 1 15 13 9 1 9 7 9 2 13 3 9 1 15 13 7 15 13 2
13 1 9 7 1 9 7 9 15 13 13 13 0 2
14 13 3 13 15 13 15 9 9 2 15 13 9 9 2
42 13 3 13 15 13 15 9 15 13 1 9 9 1 9 2 16 9 2 0 1 13 16 9 2 15 13 15 2 15 13 9 2 3 13 9 9 2 1 15 13 9 2
33 1 7 1 9 9 2 7 9 2 3 13 16 13 13 7 9 2 13 13 13 7 13 15 9 0 2 3 13 9 9 7 9 2
24 16 7 13 15 9 15 3 13 13 1 9 7 9 2 15 9 7 13 9 10 2 7 3 2
21 3 9 7 9 13 13 9 7 9 7 9 0 2 16 15 9 3 13 1 0 2
24 1 0 3 13 2 16 9 3 13 13 1 15 15 13 9 9 15 2 16 7 15 15 9 2
35 7 16 9 13 9 0 2 3 13 1 9 2 15 13 15 1 9 7 9 1 9 2 15 13 9 1 15 2 15 3 13 15 9 0 2
33 3 1 9 13 9 9 7 15 13 2 7 3 1 15 9 2 16 15 9 3 13 9 0 0 2 16 15 15 13 2 7 9 2
10 9 3 13 3 13 16 9 15 9 2
24 7 0 13 16 15 9 0 2 1 15 9 2 3 13 1 15 9 2 7 13 3 9 13 2
33 1 0 13 2 16 16 9 13 1 9 9 15 9 2 9 13 0 1 9 15 13 3 0 16 3 13 10 9 2 16 13 9 2
17 3 13 0 9 10 3 1 9 0 2 15 9 3 13 1 9 2
37 7 15 9 13 9 0 13 2 15 3 3 13 10 9 9 9 15 13 1 9 15 2 16 13 4 2 1 8 8 2 7 15 9 13 9 9 2
18 1 0 13 2 16 10 9 13 15 9 0 9 2 15 13 9 0 2
15 3 3 9 3 13 1 9 15 2 0 13 1 9 15 2
13 1 9 7 9 3 13 1 9 9 2 9 0 2
24 13 3 2 16 9 3 13 13 2 7 13 9 0 2 16 13 9 2 7 16 13 9 9 2
13 3 13 1 9 0 2 15 3 13 9 1 15 2
13 1 3 9 13 9 0 2 9 15 13 1 9 2
9 1 2 9 0 13 15 9 9 2
8 7 9 13 9 0 9 13 2
30 12 13 2 16 13 4 9 13 1 9 16 1 9 2 7 16 3 13 9 2 7 3 9 2 16 13 9 1 9 2
24 9 7 13 1 9 16 15 9 1 15 15 9 7 15 9 15 13 9 2 16 1 9 0 2
17 3 16 13 9 16 13 9 7 9 2 13 1 15 9 9 15 2
22 9 7 16 13 9 0 2 13 3 0 1 9 2 1 16 1 15 9 13 0 9 2
16 7 15 9 9 0 13 13 15 9 9 2 16 13 15 9 2
35 1 0 13 2 16 9 3 13 1 9 7 1 9 9 2 16 1 9 2 7 16 9 1 9 2 7 3 3 13 16 13 1 0 9 2
38 1 9 15 9 13 13 2 16 16 15 0 13 1 9 2 9 13 15 9 2 7 3 15 9 2 16 9 3 13 9 2 7 9 2 7 15 9 2
13 9 7 2 15 13 1 9 9 2 13 9 0 2
12 3 3 9 13 13 2 16 9 13 16 9 2
10 7 9 15 13 9 2 13 16 0 2
11 3 3 13 0 13 16 1 9 10 9 2
9 3 1 9 0 9 2 7 9 2
5 7 9 13 0 2
11 15 3 13 7 13 1 15 15 13 9 2
19 7 3 1 9 9 15 13 1 9 0 9 2 7 3 13 0 9 0 2
13 7 9 9 13 15 9 1 15 2 0 7 0 2
39 15 7 3 13 2 16 1 9 7 9 2 13 13 7 13 2 7 3 1 0 2 16 9 13 9 1 9 9 2 16 13 7 13 2 7 9 1 9 2
21 7 1 15 13 3 9 9 0 7 9 0 15 9 2 15 13 9 9 7 9 2
33 7 3 3 13 9 16 1 9 9 9 13 15 9 2 7 13 9 1 15 2 1 7 16 13 9 0 15 9 2 13 9 9 2
35 15 9 13 0 13 2 0 2 16 1 10 9 9 13 9 9 2 0 13 16 15 9 15 9 13 1 9 2 15 3 13 1 9 9 2
67 0 9 13 3 13 1 9 15 9 2 1 15 13 1 15 9 0 2 15 13 1 0 9 2 16 9 13 2 7 1 15 16 1 10 9 13 1 9 9 7 9 2 0 9 13 0 9 2 16 9 0 3 13 1 9 9 2 15 13 3 9 2 7 1 9 0 2
35 0 2 16 13 13 1 0 9 2 3 3 9 10 3 13 16 13 9 2 16 9 0 9 2 16 1 9 13 1 15 9 13 9 13 2
10 1 2 9 3 13 15 15 13 9 2
7 7 9 13 9 0 9 2
10 7 9 3 13 9 1 15 9 0 2
9 3 2 10 9 13 1 9 15 2
12 3 13 16 9 13 15 9 13 13 1 9 2
24 13 3 16 10 9 1 9 15 0 13 2 16 9 0 1 9 2 7 9 0 1 9 0 2
41 7 13 13 9 9 9 1 9 0 2 16 13 9 9 0 1 9 1 15 9 2 15 13 9 9 15 9 0 13 2 16 9 1 15 3 13 2 16 13 4 2
56 7 15 9 13 13 0 3 1 9 7 9 15 9 13 2 7 1 9 9 13 2 7 9 2 16 3 1 0 9 2 15 13 9 9 2 9 13 0 1 9 9 0 2 16 15 9 13 13 1 9 2 16 1 15 9 2
26 1 0 13 2 16 9 13 1 9 3 3 16 9 13 2 1 16 13 9 9 2 7 3 16 9 2
15 9 7 3 13 9 15 9 7 9 2 15 0 13 13 2
22 7 3 15 13 1 9 9 16 9 0 2 7 13 16 1 9 9 9 15 0 13 2
11 7 3 13 9 15 2 15 0 13 0 2
33 9 7 13 9 13 9 1 9 9 15 13 1 15 9 13 1 15 2 7 3 1 9 15 13 0 13 1 9 9 1 15 13 2
57 16 3 9 1 9 13 9 9 9 2 7 15 9 13 0 1 9 13 1 15 9 13 2 15 13 3 9 9 15 9 2 7 3 9 15 13 9 9 0 2 15 9 1 9 13 2 3 3 7 1 9 9 13 9 9 9 2
31 1 0 13 2 16 15 13 13 0 2 7 1 9 0 2 16 9 13 9 0 2 7 1 9 9 2 16 9 13 0 2
21 13 3 1 9 0 7 9 13 2 13 15 9 16 0 2 7 15 9 16 9 2
15 7 16 13 1 9 0 16 9 0 2 1 9 13 9 2
30 7 16 1 9 0 9 13 15 9 16 9 13 15 1 9 9 2 16 13 4 2 8 8 2 3 13 16 13 9 2
69 7 3 13 1 9 10 16 1 9 9 2 7 9 1 9 0 7 0 2 16 1 0 13 1 9 0 2 13 9 9 10 1 15 2 16 13 16 9 9 0 13 15 9 2 7 13 9 0 2 0 3 16 13 9 0 2 7 13 1 15 9 0 2 15 9 1 15 13 2
19 1 0 13 2 16 9 3 13 13 1 9 1 9 0 2 7 0 0 2
17 3 2 16 15 13 9 0 1 9 9 2 3 9 1 13 9 2
12 7 9 0 13 1 9 9 2 16 13 9 2
49 16 7 13 1 9 0 2 16 1 9 0 2 16 9 7 9 7 3 2 9 13 3 7 0 13 1 13 9 2 3 3 1 9 9 1 15 9 9 9 13 0 7 0 0 1 13 9 10 2
10 7 3 3 13 1 9 0 9 9 2
37 16 3 9 13 9 0 9 1 15 9 2 15 16 13 9 0 0 2 3 9 13 7 13 10 9 2 16 13 9 0 9 2 15 13 9 0 2
41 7 3 13 16 15 9 15 9 9 10 13 2 13 15 15 9 15 0 1 9 13 2 16 3 9 13 1 9 0 2 7 3 15 9 13 15 9 1 10 9 2
21 15 3 9 13 13 3 13 1 9 2 16 1 15 16 13 0 9 1 9 10 2
24 15 3 3 13 13 2 16 15 9 13 2 16 7 1 0 9 2 7 1 9 1 9 9 2
24 7 1 9 10 13 7 9 0 1 9 9 2 7 9 0 2 15 3 3 13 0 7 0 2
15 13 7 9 9 2 16 13 1 9 15 15 13 15 9 2
7 15 3 9 13 9 13 2
54 7 16 9 3 13 16 1 15 16 13 1 15 9 9 2 3 15 9 3 13 1 15 9 9 2 7 7 9 16 13 9 0 2 16 16 1 9 13 9 2 7 9 2 16 13 9 0 2 16 1 9 9 13 2
21 7 15 13 1 15 1 9 0 7 9 7 9 0 2 3 7 1 9 9 0 2
15 15 7 15 13 1 9 9 0 2 3 13 13 9 9 2
26 7 15 13 9 10 0 2 15 1 0 13 2 15 10 13 1 9 9 2 16 9 2 9 7 3 2
21 7 1 9 9 2 3 16 13 2 7 16 9 9 1 9 9 2 13 9 9 2
56 7 3 13 16 15 1 9 7 16 1 0 2 7 16 9 1 9 7 16 1 0 2 7 16 1 9 2 7 16 9 1 9 2 7 16 1 13 2 16 9 13 1 9 2 7 16 1 9 0 2 16 1 0 13 13 2
24 3 13 9 2 16 9 15 13 1 9 9 2 7 9 1 9 9 2 7 9 1 9 9 2
29 1 9 16 1 15 9 2 15 9 2 3 13 1 15 2 0 13 13 1 0 2 1 10 9 13 1 15 0 2
39 1 0 13 2 16 16 9 13 1 9 0 2 3 9 13 2 7 9 9 2 9 3 13 2 16 7 15 9 0 2 16 1 9 2 7 3 9 0 2
12 15 9 9 13 1 9 2 16 13 9 9 2
33 7 3 1 15 15 13 1 9 10 2 7 3 1 9 13 9 9 0 10 15 1 15 13 2 16 9 9 1 9 9 10 9 2
6 9 3 0 9 13 2
32 16 7 13 9 9 15 13 2 3 9 13 0 2 13 15 9 7 9 12 1 15 2 9 9 13 2 3 16 13 9 15 2
21 0 9 13 2 16 13 9 15 1 9 9 13 9 2 15 13 2 7 15 13 2
15 16 7 13 9 1 9 9 2 0 13 2 7 13 9 2
11 16 7 13 1 9 9 2 3 0 13 2
17 7 9 3 13 9 2 16 9 2 3 13 1 15 2 0 13 2
13 7 13 10 0 1 9 9 9 2 16 13 9 2
26 7 1 15 3 1 9 9 13 3 13 2 16 9 13 0 2 7 1 9 0 13 9 2 3 13 2
23 3 9 15 9 13 13 9 2 1 16 15 13 1 9 9 9 2 15 13 9 0 13 2
41 1 0 13 2 16 15 9 9 3 13 9 0 0 1 9 9 2 16 15 9 0 2 16 13 9 0 16 15 13 2 7 16 9 0 2 16 13 16 15 13 2
31 16 7 9 0 13 0 2 3 13 9 15 9 2 1 16 15 9 9 3 3 13 9 9 16 9 2 7 16 15 0 2
30 13 3 2 16 1 13 2 9 13 0 9 2 9 13 0 2 16 9 0 13 13 10 15 1 9 1 9 9 9 2
15 3 2 10 9 13 9 15 9 13 1 9 2 1 9 2
19 7 2 16 13 9 2 9 2 15 10 9 13 2 9 0 13 3 13 2
33 1 0 13 2 16 16 9 13 1 9 0 2 3 0 13 16 9 3 13 9 0 2 7 13 16 10 15 13 2 9 0 13 2
50 16 7 13 1 9 0 2 3 13 10 9 13 2 3 16 15 1 15 3 13 0 9 2 1 15 13 0 9 7 0 7 0 9 2 1 9 2 7 16 15 9 9 13 2 9 13 15 15 9 2
37 7 16 1 15 9 13 13 15 1 15 13 9 2 15 13 3 9 13 2 3 3 1 15 13 9 9 2 1 16 9 7 9 13 9 13 9 2
12 3 2 1 9 2 12 9 9 0 9 13 2
16 7 0 13 1 10 15 9 0 2 16 9 2 9 7 3 2
19 10 3 13 1 13 9 0 1 9 13 13 9 7 13 7 15 0 9 2
29 0 13 2 16 1 9 13 9 9 7 9 2 16 9 13 9 9 2 3 3 13 15 9 1 9 7 1 15 2
19 7 3 9 3 13 9 3 2 7 1 9 1 9 7 9 2 13 15 2
15 7 3 13 9 1 9 16 9 13 9 1 9 7 9 2
29 7 15 9 3 13 2 16 13 9 1 9 7 9 2 3 3 1 15 9 13 13 9 13 2 1 15 13 9 2
43 1 7 13 13 9 13 2 7 15 9 13 13 9 2 15 9 13 2 13 16 15 13 0 1 0 9 2 15 13 1 9 9 2 16 0 1 9 2 7 13 1 9 2
19 7 3 1 9 13 9 16 9 7 9 13 9 13 9 2 1 15 13 2
25 16 16 13 15 16 15 13 2 3 9 13 9 2 16 13 9 15 2 9 9 9 2 9 9 2
51 1 0 3 13 2 16 0 13 9 1 9 7 9 13 2 7 0 1 9 13 13 3 9 1 9 7 9 2 3 3 13 2 16 9 1 9 7 9 7 9 2 3 3 1 15 9 7 1 15 9 2
18 1 0 13 2 16 9 0 3 13 9 16 1 9 9 1 15 13 2
24 7 16 9 1 15 13 15 9 9 2 3 13 2 3 7 15 9 2 15 1 15 9 13 2
15 7 9 9 13 1 9 9 2 15 13 9 13 9 15 2
7 3 9 13 9 9 13 2
18 9 0 2 16 1 9 1 9 7 9 2 7 1 9 7 15 13 2
18 9 7 0 13 7 1 9 2 7 9 2 7 1 9 2 7 9 2
22 1 3 12 13 9 9 13 2 1 15 16 9 13 9 2 13 12 16 13 1 9 2
25 7 1 0 9 9 2 15 13 13 1 15 2 13 16 13 9 9 2 7 16 13 1 9 9 2
20 13 3 15 9 1 9 7 9 2 1 16 12 9 1 9 10 13 1 15 2
13 0 13 9 1 9 9 2 16 13 16 9 15 2
32 16 0 9 9 13 9 13 15 9 1 15 9 15 13 2 16 13 1 15 13 12 9 2 3 9 13 9 2 7 13 15 2
16 16 15 9 13 0 2 3 13 1 15 1 15 9 9 13 2
19 7 3 0 2 15 16 3 13 2 3 1 15 7 15 9 13 9 13 2
13 7 1 13 13 2 13 9 1 15 15 9 13 2
17 7 9 1 9 2 16 9 3 13 9 2 7 9 13 9 15 2
38 7 3 1 12 7 15 13 9 12 9 2 16 9 13 0 2 3 13 0 13 1 12 9 2 16 9 1 15 13 2 3 9 2 3 13 1 15 2
38 16 7 13 0 7 0 2 3 0 13 13 2 16 3 13 9 1 9 2 7 3 1 9 13 2 16 13 4 2 8 12 2 8 12 2 8 12 2
16 7 9 7 9 2 1 15 13 9 9 1 0 2 13 0 2
18 7 16 9 0 2 16 9 7 9 7 3 2 15 3 13 1 0 2
18 3 7 9 9 2 15 1 15 9 13 2 0 3 13 2 7 0 2
29 13 3 1 0 15 9 0 2 16 9 2 15 1 9 3 0 1 9 13 2 7 3 1 2 13 15 1 9 2
22 3 1 16 1 15 9 13 9 9 2 9 0 13 2 16 13 3 0 15 9 0 2
19 7 3 3 13 0 1 9 10 2 7 1 9 2 16 13 9 7 9 2
17 7 9 9 13 1 9 7 9 2 15 13 13 7 0 7 9 2
22 7 13 3 3 1 9 13 2 16 9 13 16 9 2 7 15 9 0 13 16 0 2
28 16 16 3 13 9 1 9 1 9 9 2 3 2 16 13 15 13 1 9 0 2 13 1 0 9 16 0 2
38 7 15 9 7 9 0 7 0 2 1 9 13 13 1 0 7 0 1 9 2 15 16 9 9 13 1 9 2 7 9 9 1 9 2 16 13 4 2
22 7 1 9 0 3 13 15 13 1 9 15 13 0 2 3 0 2 7 9 13 13 2
17 0 2 16 1 0 15 13 16 9 2 7 16 9 0 15 13 2
11 3 15 13 1 9 9 2 15 13 0 2
19 16 10 15 9 0 1 15 10 9 13 16 15 1 15 15 13 2 13 2
20 15 9 13 2 16 10 9 7 9 13 7 1 9 7 1 9 2 1 9 2
23 16 3 0 2 13 16 13 0 9 2 16 3 15 13 9 2 7 15 9 0 3 0 2
57 16 3 13 1 15 15 13 1 9 2 16 9 9 13 13 2 16 9 7 9 2 7 15 9 0 13 9 13 9 2 3 13 1 15 15 13 1 9 2 16 9 15 13 1 9 9 2 13 13 2 7 15 9 13 9 9 2
25 3 0 3 13 9 1 9 2 7 0 4 13 1 15 2 16 9 9 2 7 9 9 7 3 2
13 3 2 9 9 0 15 13 16 13 9 0 15 2
26 1 3 15 9 9 9 13 0 16 9 2 13 16 9 13 9 9 1 9 2 7 3 13 1 9 2
34 1 0 13 2 16 3 13 0 9 1 9 7 9 2 16 9 0 13 15 9 13 9 9 0 7 0 2 7 13 2 7 3 9 2
9 7 9 13 0 13 9 9 0 2
19 3 2 9 3 13 1 9 16 1 16 13 1 9 9 15 1 15 13 2
15 7 1 9 2 16 9 9 2 16 9 7 9 1 9 2
23 3 2 15 15 13 9 0 9 2 13 13 9 0 2 16 0 9 13 1 0 9 13 2
27 1 0 13 2 16 9 3 13 9 9 1 9 3 9 13 15 9 2 7 0 3 13 15 9 1 9 2
23 7 9 0 3 13 9 2 13 9 9 2 15 13 9 2 16 9 13 9 9 1 0 2
18 15 7 9 15 13 9 2 13 15 9 2 7 9 1 9 9 13 2
19 7 9 9 9 13 16 15 9 9 7 9 13 1 13 1 15 15 13 2
25 0 2 16 10 9 7 13 1 9 9 2 16 0 7 9 2 7 9 9 2 16 9 7 9 2
15 15 9 13 2 16 9 9 1 9 15 3 13 16 0 2
11 16 9 9 0 13 1 9 0 9 0 2
21 7 15 13 13 13 2 16 1 0 9 9 7 9 13 1 9 7 9 9 13 2
26 9 7 15 13 15 9 9 2 1 16 0 13 2 13 15 9 7 9 2 16 15 9 9 13 9 2
42 16 3 9 13 1 9 2 15 3 13 16 13 2 7 1 15 3 13 1 13 0 9 9 13 2 7 9 2 16 1 13 4 2 12 8 2 8 12 2 8 12 2
18 3 3 13 15 15 13 1 9 1 16 13 2 16 16 13 9 9 2
28 15 7 9 0 1 15 13 9 9 2 13 3 1 13 7 3 1 0 2 16 3 13 9 9 1 9 0 2
15 3 2 1 9 1 9 7 1 9 3 13 9 16 9 2
14 7 9 16 4 13 1 9 2 13 9 7 9 9 2
28 1 3 1 0 3 13 9 16 9 2 15 13 1 15 9 2 13 16 15 13 1 9 0 2 13 1 9 2
19 1 13 16 10 13 12 1 9 2 7 13 9 3 0 2 7 3 9 2
8 16 3 9 2 3 0 13 2
50 1 0 3 13 2 16 1 13 16 10 13 12 1 9 2 9 1 3 3 13 9 9 1 9 0 2 7 3 1 9 9 2 16 9 9 13 9 9 2 3 0 9 2 15 1 0 10 12 13 2
13 7 3 15 13 2 16 0 15 13 1 9 9 2
17 7 15 3 1 15 3 13 0 2 16 9 3 13 15 16 13 2
30 7 3 1 9 0 3 15 13 1 9 16 0 2 7 16 1 15 0 2 3 13 13 16 13 16 9 13 9 9 2
29 7 3 9 13 9 9 9 15 15 13 9 2 15 9 13 2 7 3 1 9 0 2 7 0 2 7 9 13 2
57 7 3 15 13 2 15 13 13 9 9 1 8 9 3 1 2 16 13 1 9 3 9 0 2 16 13 9 0 9 10 15 15 1 9 13 2 16 0 1 0 3 13 0 7 9 2 7 0 13 2 15 13 9 9 1 13 2
21 7 1 15 3 13 9 16 1 9 0 2 15 13 1 15 9 7 0 7 0 2
18 7 16 15 9 9 13 15 9 0 2 3 15 13 13 13 12 9 2
16 7 9 2 15 13 9 9 1 9 2 7 1 15 9 9 2
37 16 7 13 0 2 3 2 16 9 13 9 15 13 9 15 9 2 13 9 13 9 15 9 15 13 9 9 9 0 2 16 9 13 9 9 9 2
25 7 3 3 13 1 9 15 9 2 7 1 9 9 16 9 13 9 2 7 0 16 9 13 13 2
12 7 9 13 1 9 9 13 1 15 15 13 2
21 15 7 13 13 1 15 1 9 9 7 0 7 0 2 13 16 9 15 1 15 2
8 16 9 0 13 9 0 9 2
8 9 7 3 13 1 9 9 2
16 1 3 9 13 1 9 2 13 16 3 13 13 0 9 13 2
16 16 9 15 15 13 0 2 13 13 1 0 1 9 9 0 2
30 15 0 9 9 13 13 1 0 1 9 3 7 3 0 2 3 9 9 2 16 1 13 16 9 13 9 1 9 10 2
21 16 15 13 9 15 9 2 13 13 13 1 9 15 2 16 9 13 13 1 9 2
5 7 1 13 9 2
34 16 7 13 13 15 9 15 13 15 9 9 2 15 3 9 13 13 2 3 1 9 13 7 1 15 0 13 2 7 9 13 7 15 2
13 3 1 15 15 9 1 13 9 1 0 3 9 2
18 16 1 9 9 13 2 3 9 7 9 2 13 12 9 7 12 9 2
16 3 2 10 9 13 9 15 15 13 9 3 1 15 10 9 2
37 0 1 9 0 12 13 2 3 9 2 7 9 2 16 15 13 1 0 2 13 1 9 9 2 15 3 13 13 7 13 1 15 2 7 1 15 2
15 1 0 13 2 16 9 13 1 9 9 7 9 1 0 2
17 9 7 9 7 9 3 13 0 9 1 9 15 2 7 9 9 2
16 1 0 13 2 16 9 13 1 9 9 2 7 9 13 13 2
15 3 2 15 13 1 15 9 2 13 16 13 15 1 15 2
28 7 9 15 15 9 3 0 13 1 9 2 13 15 0 15 9 15 9 13 1 9 2 3 9 0 1 9 2
27 3 15 3 0 13 13 16 9 2 15 13 9 0 9 2 3 7 9 7 9 2 15 13 1 9 9 2
23 16 9 13 16 9 15 2 16 13 0 2 7 9 16 9 15 2 16 13 0 7 0 2
34 7 13 15 9 1 9 10 2 15 13 1 0 15 13 15 12 1 9 2 15 12 15 13 2 16 9 1 15 13 13 9 0 0 2
23 7 9 13 15 0 1 9 2 15 13 9 2 7 15 0 2 15 15 13 9 1 0 2
19 16 15 13 16 9 2 16 9 2 7 15 16 0 1 9 2 16 9 2
25 1 0 3 13 2 16 16 9 7 9 13 15 9 2 3 13 9 2 16 12 16 9 15 13 2
26 1 0 13 2 16 3 13 3 3 9 1 9 2 7 1 9 9 2 16 13 4 2 1 8 8 2
21 7 16 9 3 13 16 9 12 9 2 3 3 13 13 16 12 9 13 12 9 2
22 7 3 13 9 9 0 7 0 2 3 7 9 7 9 2 15 13 0 16 9 9 2
28 1 0 13 2 16 15 9 15 13 1 9 9 2 13 12 0 2 15 12 13 15 9 2 7 15 9 9 2
8 15 3 13 1 9 15 9 2
31 1 1 9 10 9 7 9 13 2 15 16 15 13 9 0 7 0 2 13 9 15 13 13 1 9 2 7 13 9 3 2
12 16 7 9 9 13 9 2 3 9 13 9 2
6 3 9 9 9 13 2
16 3 13 16 10 9 1 15 13 13 1 9 2 13 0 9 2
40 16 7 3 13 1 15 0 2 7 3 9 15 0 2 3 13 9 7 9 13 2 3 10 9 3 1 15 0 3 13 7 13 9 9 2 16 9 1 9 2
45 15 7 13 0 2 16 15 13 13 9 15 7 9 15 2 7 1 15 13 2 16 9 3 13 13 9 16 13 9 9 7 15 15 13 13 2 16 9 13 13 2 7 9 13 2
19 13 3 1 9 13 9 15 0 2 16 9 1 9 13 9 0 10 9 2
24 7 3 16 9 13 1 9 13 15 9 2 3 13 0 13 2 1 16 3 9 3 0 13 2
71 7 3 1 10 15 13 1 9 9 7 9 13 15 9 2 16 10 9 13 10 9 2 1 15 13 1 15 9 2 16 13 9 3 1 9 2 7 13 3 1 9 2 7 3 1 15 2 16 13 9 3 13 15 1 9 2 7 3 1 15 2 3 15 1 9 7 9 0 13 13 2
30 1 0 3 13 2 16 1 9 1 9 3 13 9 0 16 16 13 13 13 1 13 15 9 9 2 7 1 15 9 2
35 7 3 15 9 13 13 1 13 9 1 9 1 9 15 1 15 13 2 16 7 9 9 13 13 9 0 1 9 2 16 1 9 10 13 2
18 0 2 16 15 15 3 13 9 4 13 2 7 9 13 3 13 9 2
32 16 9 16 1 9 9 13 13 13 15 9 2 3 1 9 7 9 2 1 9 9 15 13 1 15 2 13 9 15 7 15 2
19 7 16 1 9 10 3 13 16 9 2 3 9 10 13 0 9 9 9 2
40 1 0 3 13 2 16 2 16 1 13 13 2 9 1 15 9 0 13 7 13 0 2 16 9 3 13 2 7 0 2 16 1 9 7 1 9 15 0 13 2
22 7 3 13 9 7 9 9 15 15 1 9 13 2 7 9 7 9 2 16 13 4 2
37 7 3 15 15 13 2 16 0 13 16 13 2 0 16 13 2 13 13 1 9 10 2 15 1 9 13 1 9 0 2 7 1 9 1 9 0 2
9 7 9 13 1 9 9 7 9 2
24 7 15 13 13 2 16 9 9 15 1 9 13 2 13 9 16 13 16 9 15 7 9 9 2
14 7 9 2 1 15 16 1 9 13 9 2 9 13 2
26 3 2 9 13 1 12 8 16 16 10 9 13 1 9 1 0 9 2 3 13 1 9 1 0 9 2
13 7 15 15 13 9 2 16 9 9 1 9 13 2
55 13 13 2 16 2 16 9 0 13 0 9 2 12 1 9 1 16 13 1 9 2 15 1 9 1 16 13 1 9 9 2 3 3 1 9 0 2 7 0 2 3 3 9 0 13 0 9 2 16 13 9 1 12 8 2
16 7 3 9 9 1 9 13 9 13 2 15 13 16 9 0 2
10 9 3 13 1 8 2 15 13 9 2
12 9 3 9 1 9 13 2 15 9 9 13 2
38 16 3 1 9 13 9 13 1 9 15 13 9 0 9 2 1 16 9 0 9 9 13 2 3 3 9 0 9 13 2 1 16 9 13 9 9 13 2
22 3 15 13 9 3 13 2 7 1 9 15 9 13 9 0 1 15 13 1 9 13 2
27 3 2 16 13 4 2 9 15 13 1 9 15 13 2 16 9 9 2 15 13 1 9 9 2 1 9 2
18 7 9 9 13 1 9 9 15 13 1 9 9 2 7 3 1 0 2
24 9 3 2 16 1 13 13 2 8 8 2 13 9 16 13 2 7 3 16 13 1 9 13 2
24 3 3 15 9 13 1 9 9 9 7 9 2 16 9 9 3 13 1 9 16 16 9 13 2
16 16 13 9 2 15 13 15 3 1 9 13 2 16 9 15 2
6 3 2 9 13 9 2
9 13 3 1 8 2 15 13 9 2
21 7 9 0 3 13 15 9 2 16 7 0 9 2 15 13 9 2 13 15 9 2
19 7 0 16 3 2 3 13 13 9 2 1 10 0 12 9 1 9 13 2
24 7 3 9 2 1 9 10 9 2 13 9 9 1 9 2 9 0 0 2 7 9 15 9 2
15 7 3 9 9 7 9 13 1 9 2 15 9 13 9 2
18 1 9 3 15 0 9 0 13 15 9 15 13 2 16 9 7 9 2
19 15 7 9 7 13 1 9 7 9 2 7 1 9 2 7 1 9 15 2
9 1 9 2 16 9 13 1 9 2
17 7 15 13 0 2 16 9 7 13 9 9 2 7 13 9 9 2
20 3 9 0 13 13 9 0 9 10 16 13 9 9 2 16 3 9 15 13 2
10 7 1 16 13 9 9 7 3 9 2
27 7 3 15 9 0 13 13 1 9 2 3 16 1 9 2 7 16 13 1 13 2 7 16 9 1 9 2
19 1 0 13 2 16 9 13 1 9 16 9 13 9 2 7 13 9 0 2
49 3 3 9 9 13 13 9 9 2 7 1 0 9 0 2 16 13 1 9 0 9 7 1 9 9 7 9 2 7 1 0 9 0 15 9 13 1 9 7 9 15 9 2 16 1 9 9 0 2
45 3 0 9 1 15 2 3 13 13 9 1 15 2 16 13 1 15 9 1 15 13 9 1 9 1 9 2 7 1 0 2 16 1 9 7 9 2 7 9 2 7 1 10 3 2
30 7 1 15 3 9 13 13 13 9 2 1 13 9 3 3 13 1 9 7 9 2 7 9 13 3 1 9 7 9 2
35 7 1 3 9 15 13 13 3 2 7 1 9 2 16 1 0 9 9 2 15 13 9 13 2 13 15 9 7 9 2 15 15 0 13 2
16 3 3 13 0 7 0 1 9 9 2 16 3 13 9 0 2
29 3 2 1 9 13 15 9 1 9 2 13 16 1 10 9 7 12 0 13 9 15 2 7 15 1 12 9 13 2
18 0 9 13 9 1 15 13 9 2 1 15 9 9 9 13 9 13 2
27 7 3 13 16 15 13 1 9 1 9 1 9 9 2 7 1 9 2 3 13 1 9 9 16 1 9 2
20 3 13 16 9 2 15 13 9 1 9 7 1 9 2 3 13 1 9 9 2
16 7 3 9 13 9 9 2 1 16 13 9 0 9 7 9 2
15 3 9 16 13 1 9 9 9 2 3 13 1 9 9 2
37 15 7 13 9 9 2 13 9 2 16 3 9 9 1 9 7 9 13 2 1 15 9 13 2 13 1 15 9 9 1 9 2 7 9 1 9 2
45 1 0 3 13 2 16 15 13 1 9 13 1 9 9 7 1 9 9 15 13 1 9 0 2 16 9 15 13 1 9 9 2 3 13 9 15 15 13 1 9 2 7 3 9 2
20 7 3 13 15 9 2 7 10 15 13 9 1 9 9 2 13 16 0 13 2
33 3 1 9 3 3 13 9 9 2 7 3 15 9 13 1 15 9 2 7 10 9 15 13 9 7 1 9 9 7 1 9 9 2
24 1 2 15 9 13 3 1 9 0 2 1 15 9 13 13 2 3 7 1 9 0 1 9 2
34 7 3 13 15 9 1 15 13 15 3 13 2 16 1 9 13 9 9 1 9 13 2 3 13 13 16 15 9 13 9 1 9 15 2
17 3 16 13 15 15 9 2 3 13 9 15 9 2 7 9 3 2
35 7 13 0 2 16 16 15 13 13 13 9 9 2 3 7 9 2 1 16 1 15 13 9 0 9 2 16 9 9 1 9 9 15 13 2
21 15 9 10 3 13 13 2 16 3 13 0 0 13 16 1 0 9 1 15 13 2
22 7 3 9 10 13 3 13 0 2 16 13 9 0 2 15 13 1 9 1 0 0 2
60 16 3 9 9 13 15 1 9 2 1 16 13 1 9 9 16 9 9 13 2 7 1 16 13 1 9 7 9 16 9 13 2 3 3 9 9 9 15 9 13 1 9 0 2 16 9 13 2 7 15 1 9 0 2 15 9 9 0 13 2
32 7 15 13 9 9 2 7 9 13 1 15 16 1 9 3 0 13 9 0 2 1 15 13 9 10 9 9 2 16 13 9 2
16 3 2 10 9 13 1 15 9 13 2 16 1 9 13 15 2
10 15 9 2 1 16 13 1 13 9 2
33 7 15 16 13 1 0 2 16 9 13 9 1 15 13 2 3 13 1 9 2 1 16 13 9 9 2 7 13 15 13 1 9 2
39 7 3 2 16 9 13 3 13 9 9 7 9 2 16 15 1 15 9 13 9 2 15 9 3 13 9 2 3 3 13 0 9 9 9 2 7 13 3 2
13 7 1 15 10 9 9 13 2 3 15 9 13 2
20 1 15 2 16 13 9 1 15 9 15 9 13 13 2 16 9 9 9 0 2
10 13 12 9 1 9 2 7 13 15 2
22 7 9 0 2 15 1 15 13 0 1 10 9 2 3 7 0 13 2 13 1 9 2
24 7 0 9 2 15 2 3 1 15 13 2 13 13 0 9 9 2 13 1 9 1 15 13 2
13 10 3 9 1 0 9 16 0 13 2 9 13 2
30 15 7 4 1 10 9 13 1 12 2 16 13 2 15 1 15 9 13 2 7 13 9 9 2 15 1 15 9 13 2
8 16 15 13 7 9 7 9 2
11 3 3 12 8 13 2 16 9 13 9 2
12 7 9 15 13 13 9 9 2 9 9 13 2
18 7 1 9 9 9 15 9 13 13 2 16 15 3 9 7 9 13 2
24 16 3 15 13 0 9 1 9 15 13 13 2 3 13 1 15 9 2 16 9 15 9 13 2
18 16 3 9 9 3 13 2 3 13 9 13 2 7 9 1 9 13 2
17 16 13 9 9 2 1 15 13 9 2 7 9 13 0 9 9 2
18 12 15 13 9 9 13 1 9 1 15 16 15 13 13 1 9 9 2
27 7 16 9 9 13 1 9 1 15 15 13 1 9 2 13 16 3 9 9 13 1 15 16 13 1 9 2
10 3 2 9 13 9 12 1 9 12 2
28 13 13 2 16 9 13 9 1 9 12 2 7 3 15 13 16 9 15 13 9 9 2 16 1 12 8 13 2
13 7 1 15 16 13 12 9 2 16 12 0 9 2
16 7 1 15 16 12 15 0 13 9 2 13 15 15 0 13 2
8 9 3 13 1 9 1 9 2
16 7 9 7 9 9 13 15 13 2 16 7 13 13 9 13 2
12 16 9 0 3 13 1 9 2 7 1 9 2
14 1 9 3 13 9 9 2 7 1 15 13 9 9 2
16 9 7 15 9 0 13 1 9 2 15 13 9 9 13 9 2
23 1 0 13 2 16 16 9 0 13 1 9 1 9 2 3 9 9 13 1 13 1 9 2
38 7 16 9 0 1 9 13 13 9 3 13 9 2 16 9 3 13 9 1 9 0 2 3 3 13 0 1 9 2 15 13 0 9 2 3 9 13 2
15 3 13 16 1 15 9 15 13 1 9 9 2 3 13 2
13 7 3 13 3 1 15 9 15 13 1 9 9 2
9 7 3 9 7 9 1 15 9 2
46 0 9 3 2 1 16 9 1 9 13 9 15 15 13 1 9 9 2 16 10 9 13 1 9 2 7 13 9 15 13 9 2 7 15 9 13 13 2 7 13 1 9 13 15 13 2
15 9 3 3 13 1 9 13 9 9 2 7 13 9 0 2
9 7 13 9 0 2 13 9 9 2
9 13 3 9 13 9 7 9 15 2
17 0 7 9 2 15 9 13 9 2 13 9 9 0 13 1 15 2
12 3 10 9 13 1 0 9 16 1 9 0 2
27 7 15 13 1 15 15 1 9 2 7 1 15 1 9 2 13 9 1 15 15 2 3 13 9 1 9 2
25 3 1 15 1 15 9 13 2 16 9 13 9 15 3 13 2 7 1 9 13 1 9 9 13 2
28 3 9 13 7 0 3 3 15 13 1 10 15 15 1 9 13 2 7 1 9 2 15 1 9 1 9 13 2
11 7 0 3 9 0 3 13 7 13 4 2
25 1 0 13 2 16 9 0 2 16 13 2 3 13 1 15 9 13 2 16 13 1 9 9 9 2
10 7 9 7 13 3 13 9 9 15 2
15 10 9 0 15 9 13 15 9 2 7 0 2 7 0 2
20 15 13 1 15 16 3 13 0 15 13 9 0 1 12 2 7 0 1 15 2
15 3 9 2 15 13 9 9 2 3 13 13 9 0 9 2
9 3 15 9 9 13 15 9 0 2
13 16 10 15 13 2 13 13 13 1 9 7 9 2
23 1 7 1 15 9 2 15 3 16 13 0 2 3 3 13 9 0 2 1 3 13 0 2
26 3 9 1 9 3 13 15 2 7 9 13 15 9 2 15 1 15 13 13 2 3 1 15 9 13 2
10 9 0 13 3 13 13 16 1 9 2
18 7 3 3 13 0 9 2 15 13 1 15 16 0 9 0 13 9 2
22 15 9 15 0 13 9 15 13 2 9 13 2 15 13 9 2 13 13 9 1 9 2
30 7 3 1 15 9 13 9 9 2 15 13 16 10 9 13 1 9 2 7 9 0 3 13 16 13 9 1 9 9 2
11 7 3 16 13 13 1 15 13 1 9 2
11 7 15 13 3 9 2 3 9 7 9 2
9 3 9 2 3 16 1 9 13 2
27 0 13 9 2 0 1 15 2 3 16 10 9 13 1 9 1 9 0 2 3 7 9 16 13 9 13 2
17 7 9 0 13 3 9 2 7 9 2 13 9 1 9 1 9 2
24 7 15 9 0 1 10 9 13 3 9 15 9 13 2 15 3 9 13 2 7 9 9 13 2
28 3 3 13 2 15 9 13 2 16 13 13 9 2 7 16 13 15 1 15 2 16 3 13 9 2 7 9 2
9 3 9 0 13 1 9 9 0 2
21 7 3 1 15 9 3 3 13 9 1 9 9 0 2 7 3 1 9 9 0 2
7 7 9 3 13 1 9 2
13 3 9 1 0 13 9 9 10 2 15 9 13 2
30 16 7 9 0 13 1 9 0 2 16 3 13 9 16 1 9 1 9 15 2 3 9 0 13 1 9 1 13 9 2
16 3 3 9 13 16 1 9 9 2 15 13 3 7 3 13 2
12 7 1 15 13 10 13 3 3 1 9 0 2
10 3 16 9 13 9 2 3 9 9 2
26 16 13 1 9 2 15 9 13 1 13 15 2 16 15 9 2 1 15 13 9 9 2 13 9 9 2
12 16 15 3 13 16 9 15 9 2 7 9 2
16 13 13 2 16 9 7 9 13 1 3 2 16 9 7 9 2
36 3 9 15 9 7 9 1 9 13 2 16 1 10 9 0 2 16 9 13 9 2 7 9 15 13 1 9 9 2 13 9 15 13 1 9 2
15 7 3 3 13 1 9 1 15 2 3 16 13 9 15 2
31 7 3 10 9 9 7 9 13 1 9 0 9 2 7 1 15 13 2 16 13 0 13 16 9 0 2 15 13 9 9 2
59 7 16 0 13 15 1 15 16 0 13 0 15 2 3 10 9 0 13 1 9 9 0 3 13 2 15 9 9 0 9 13 2 7 1 15 3 9 0 2 3 9 0 2 13 13 9 0 13 1 9 9 2 16 1 12 1 9 13 2
23 3 1 9 9 1 9 13 1 0 13 2 13 16 9 3 13 9 0 2 16 9 9 2
29 7 9 13 9 13 1 9 15 9 1 15 9 13 13 2 16 15 9 3 13 13 1 15 9 2 16 13 9 2
38 1 0 13 2 16 1 15 9 9 13 2 16 9 9 13 2 16 9 13 1 9 16 9 1 0 2 16 9 1 9 2 7 3 16 9 1 9 2
25 7 3 13 16 9 9 0 0 13 9 16 9 9 2 7 9 9 2 16 1 12 1 9 13 2
14 7 15 9 13 1 15 16 15 13 15 0 16 9 2
10 15 7 9 9 7 15 9 9 13 2
20 1 9 7 9 3 13 1 0 9 2 7 9 13 9 2 7 9 13 9 2
12 1 0 13 2 16 1 9 13 15 9 9 2
12 7 3 15 9 13 0 2 3 0 9 13 2
12 3 9 9 13 3 0 16 9 9 7 9 2
14 1 7 10 9 9 0 0 13 2 3 0 13 9 2
23 16 3 9 9 9 13 16 9 2 3 3 16 9 0 3 13 9 0 1 15 13 13 2
12 1 3 9 13 9 2 0 9 13 0 9 2
14 3 13 16 9 0 13 13 9 2 15 13 0 9 2
11 3 2 0 9 3 13 9 0 16 9 2
6 7 9 13 0 9 2
16 3 2 3 9 13 0 2 3 3 13 1 9 9 7 13 2
17 13 13 2 16 13 15 9 2 3 9 0 2 9 3 13 13 2
29 13 2 16 1 15 9 13 2 16 13 9 0 1 15 0 1 9 0 2 7 7 15 7 9 1 9 9 13 2
17 16 15 13 12 9 2 1 12 8 2 9 2 9 2 7 9 2
20 3 2 1 15 2 9 7 9 7 9 13 1 15 2 16 1 12 8 13 2
24 9 7 15 13 9 9 3 13 1 15 1 15 9 13 1 9 2 7 1 15 9 7 9 2
19 7 12 15 13 9 9 2 3 9 7 9 2 15 1 15 0 9 13 2
26 9 3 13 9 1 9 9 13 2 7 3 1 9 10 15 9 13 2 16 13 9 2 1 12 8 2
9 3 2 1 0 9 13 0 9 2
10 7 1 9 9 0 13 9 9 0 2
21 1 0 13 2 16 0 9 15 3 13 13 1 9 1 9 2 13 1 9 9 2
23 3 15 9 0 13 1 15 9 13 1 9 9 7 13 2 7 9 0 2 0 2 0 2
16 12 3 9 13 3 0 2 16 3 13 13 1 9 7 9 2
9 3 9 13 13 1 9 7 9 2
10 13 16 9 13 13 1 9 7 9 2
18 7 9 9 2 1 16 13 9 2 13 16 13 13 1 9 7 9 2
30 9 3 13 1 8 9 16 9 2 13 0 2 3 9 7 9 2 13 1 0 2 3 1 9 2 1 1 9 13 2
16 1 3 9 13 1 9 9 2 13 16 1 9 7 9 13 2
9 7 9 9 9 13 9 7 9 2
36 1 3 9 15 13 1 9 9 2 13 15 9 2 3 16 1 15 13 2 13 16 3 9 2 15 13 1 15 9 2 1 9 7 9 13 2
9 7 15 13 13 1 9 7 9 2
16 3 13 9 1 8 1 8 2 16 9 0 9 13 3 13 2
13 3 3 13 3 9 2 7 3 13 9 9 15 2
17 16 9 0 13 9 2 3 16 13 9 0 2 7 16 13 15 2
21 3 9 13 1 9 3 4 13 16 1 9 2 16 13 9 9 2 16 13 9 2
19 7 3 16 9 15 13 13 9 2 9 13 1 15 3 4 13 1 9 2
8 7 3 1 9 15 3 13 2
19 15 3 9 13 2 16 9 0 3 13 0 2 16 16 1 9 9 13 2
21 7 15 3 13 9 1 9 15 9 2 1 10 9 1 9 1 9 9 0 13 2
18 7 13 15 1 15 2 7 0 2 7 13 1 9 0 2 7 0 2
36 1 3 12 0 13 12 9 2 7 1 9 0 3 13 15 9 2 13 16 10 9 16 13 1 15 13 15 9 2 7 13 2 13 15 15 2
10 3 13 16 15 9 13 13 9 9 2
32 1 9 1 9 7 9 13 2 9 9 2 15 9 7 9 13 2 1 9 9 1 9 13 2 16 9 1 9 9 7 9 2
14 7 13 1 15 9 2 7 9 2 15 13 9 10 2
14 7 16 15 9 13 9 2 13 13 1 9 7 9 2
28 7 3 9 7 9 2 15 13 9 9 2 1 3 13 2 3 13 1 9 9 16 9 2 7 0 16 9 2
29 3 9 13 13 2 16 1 12 15 2 3 9 2 9 2 7 9 2 1 15 0 9 13 1 9 9 16 9 2
18 3 7 13 16 10 15 13 1 9 9 2 13 13 1 9 7 9 2
21 9 3 0 13 9 3 16 13 9 0 2 7 16 13 15 2 3 1 9 13 2
21 7 9 13 9 16 13 9 0 2 3 13 15 2 16 9 1 9 13 9 0 2
30 1 0 13 2 16 9 3 0 2 15 13 10 9 2 16 9 0 2 1 15 9 3 13 2 15 9 13 13 9 2
19 7 9 0 0 15 3 13 10 9 2 9 9 15 13 2 13 9 13 2
15 3 2 10 9 2 3 13 1 15 2 0 13 7 0 2
6 7 9 13 9 0 2
18 7 9 0 2 15 13 9 9 2 3 13 9 0 2 7 3 0 2
19 7 1 9 1 15 13 13 1 15 16 1 15 16 9 0 13 3 13 2
20 1 0 3 13 2 16 9 0 3 13 16 1 9 2 1 15 13 9 13 2
30 7 9 15 3 13 0 2 3 13 9 13 2 7 1 10 9 13 1 9 15 15 3 1 9 13 13 16 9 0 2
13 16 9 9 9 13 1 15 16 1 0 13 0 2
16 1 0 13 2 16 9 15 4 13 1 9 2 13 0 13 2
34 16 3 0 13 2 1 15 9 7 9 13 9 16 1 9 9 2 13 16 9 0 7 0 2 3 13 1 15 9 2 13 12 3 2
28 3 15 13 1 15 2 13 15 9 2 15 16 13 1 15 1 9 2 3 1 0 9 2 15 3 15 13 2
41 15 9 1 9 13 13 2 13 2 16 15 9 13 15 9 1 15 2 16 9 0 7 0 13 12 2 16 0 9 1 15 0 9 13 2 13 1 0 9 9 2
15 3 3 12 9 9 2 0 9 13 7 13 3 13 13 2
14 7 15 9 13 1 9 1 9 13 2 16 9 0 2
20 7 10 9 7 9 15 13 1 0 9 9 2 13 1 0 7 0 1 9 2
27 1 0 3 13 2 16 16 9 13 9 0 2 16 7 9 2 3 9 3 13 9 1 9 16 1 9 2
14 7 9 9 7 9 13 9 9 7 9 2 16 13 2
30 3 13 2 1 9 3 13 13 1 9 7 9 2 7 12 13 1 9 1 15 9 2 16 3 13 3 1 9 13 2
16 16 1 9 9 13 1 9 9 2 7 9 13 1 9 9 2
14 7 3 1 9 9 13 9 2 7 1 9 9 9 2
21 3 7 3 16 9 13 9 2 7 9 9 2 1 15 13 9 2 7 15 13 2
11 7 16 9 13 9 15 2 3 0 9 2
9 7 9 9 15 2 3 0 9 2
12 3 15 13 13 1 9 7 9 7 1 15 2
11 7 3 13 16 9 13 9 16 9 9 2
26 0 9 0 13 1 15 15 0 1 9 13 2 1 15 13 1 9 7 9 13 0 16 9 1 9 2
20 7 9 16 13 9 15 9 2 3 13 1 9 9 16 9 2 7 16 9 2
26 1 3 9 3 13 9 16 1 16 13 9 2 13 16 13 0 3 13 13 13 1 9 9 1 9 2
10 3 2 15 9 7 9 13 15 0 2
33 7 9 7 9 13 15 9 2 16 0 10 9 1 9 13 9 13 2 15 9 0 13 9 2 16 9 1 8 12 1 8 13 2
22 15 3 13 2 16 9 3 13 1 9 9 16 9 2 7 16 9 2 1 13 9 2
21 7 1 15 9 0 7 9 0 3 13 1 9 9 16 9 2 7 0 16 9 2
22 7 3 13 16 13 1 9 9 16 9 2 7 3 16 9 2 16 13 9 15 9 2
19 7 3 13 15 9 2 16 9 15 13 9 0 2 15 3 13 9 9 2
11 15 0 13 9 7 9 2 16 9 0 2
24 15 15 9 13 13 2 16 1 9 7 9 9 9 7 9 13 2 16 1 1 9 13 4 2
45 1 15 3 16 9 9 9 7 9 13 2 13 1 9 15 15 9 9 13 2 16 9 2 7 3 2 1 15 9 0 13 2 1 15 16 0 13 13 9 13 1 12 1 15 2
27 1 0 3 13 2 16 9 3 13 0 9 2 16 9 12 13 0 15 2 7 16 9 12 0 13 15 2
18 16 9 15 9 13 2 15 13 1 9 9 3 13 2 16 13 9 2
14 16 15 15 13 9 16 13 9 2 13 9 9 0 2
15 3 2 1 8 1 9 13 2 16 10 9 13 0 9 2
8 3 13 16 9 1 9 13 2
19 1 9 0 0 9 9 13 13 15 1 9 9 2 7 13 16 9 15 2
28 7 3 13 9 9 1 9 9 2 7 9 1 9 9 2 16 9 13 9 13 2 15 9 13 9 9 0 2
31 7 15 9 9 0 7 0 13 9 1 9 13 2 16 9 0 2 16 9 0 13 1 9 9 2 1 15 9 15 13 2
13 7 3 16 15 13 1 12 9 0 9 15 13 2
26 7 3 9 0 9 13 13 2 16 9 15 1 9 13 4 9 1 13 2 4 3 9 13 1 13 2
25 3 7 3 13 1 9 9 2 1 3 13 9 7 9 15 15 1 9 13 2 3 9 7 9 2
42 3 2 15 15 13 1 15 15 1 9 1 9 13 2 16 1 10 9 13 0 9 2 1 15 13 9 3 0 2 3 1 0 2 7 1 15 0 2 3 1 9 2
18 13 13 2 16 2 1 9 7 9 13 13 9 0 9 13 3 0 2
13 7 3 13 3 2 16 13 1 15 0 9 0 2
12 7 3 13 16 15 9 13 0 9 3 13 2
18 7 3 1 0 9 13 2 3 9 15 13 0 2 7 0 0 9 2
9 7 15 9 9 9 3 13 0 2
20 13 3 15 0 1 9 2 15 13 0 9 15 2 16 9 9 1 9 9 2
32 7 1 15 9 13 0 9 9 1 9 0 13 2 3 3 16 13 0 2 7 16 13 0 0 2 16 15 0 9 0 13 2
53 0 3 13 0 3 1 9 2 3 1 9 2 15 13 9 9 1 9 9 2 1 15 13 16 9 9 15 9 0 13 0 2 15 9 13 0 1 13 2 16 3 1 15 2 15 13 15 9 1 0 0 9 2
24 7 15 9 13 2 16 9 0 0 1 9 0 13 9 2 16 9 1 9 10 9 13 10 2
23 1 0 13 2 16 9 13 2 16 9 0 0 3 13 0 1 9 0 2 15 13 13 2
18 16 10 15 13 9 1 9 0 2 13 0 1 0 2 7 3 0 2
10 13 16 9 1 9 0 0 3 13 2
14 15 3 13 2 16 9 1 9 13 0 9 0 13 2
18 3 1 1 9 13 9 9 9 0 2 1 3 9 10 0 13 13 2
27 7 3 1 15 9 15 13 2 16 1 9 15 9 0 1 15 0 7 15 13 9 9 16 15 0 13 2
33 15 0 13 2 16 1 9 0 15 13 2 13 9 0 2 1 16 1 0 9 13 13 15 9 9 2 15 3 13 13 1 15 2
9 16 9 9 3 13 16 1 9 2
18 3 15 9 13 2 3 13 9 15 0 0 2 16 13 1 9 13 2
12 3 13 3 9 13 2 3 13 9 7 9 2
14 7 1 15 9 1 9 13 9 9 15 13 1 9 2
23 7 9 13 9 9 2 3 0 3 1 9 2 7 3 3 1 9 2 15 13 9 9 2
17 3 9 1 9 0 13 9 9 3 1 15 2 3 9 7 9 2
24 9 7 15 13 1 9 9 2 13 0 9 0 1 9 0 13 2 16 13 0 0 1 15 2
41 7 3 1 15 0 3 13 2 15 13 1 9 2 16 1 9 15 9 1 9 7 9 2 16 3 9 9 0 2 15 1 0 13 2 13 9 0 1 9 13 2
21 7 3 3 9 0 15 13 1 9 9 2 13 9 9 2 3 3 1 9 0 2
16 16 15 15 9 13 1 15 9 0 13 2 15 9 0 13 2
32 3 2 1 0 9 13 16 9 13 10 15 13 0 9 2 16 1 15 15 13 13 2 0 0 16 15 9 13 9 0 13 2
16 16 16 15 13 9 0 1 9 0 2 3 9 0 1 9 2
29 1 0 3 13 2 16 1 9 9 3 13 15 9 9 15 9 15 13 7 13 13 2 16 13 1 0 7 0 2
16 1 15 3 9 15 0 13 9 13 1 9 2 9 0 13 2
25 1 3 9 13 9 9 2 13 1 15 9 9 13 1 9 15 13 13 2 7 9 1 9 0 2
18 3 9 9 7 0 15 9 13 1 9 0 2 9 13 9 9 0 2
28 1 0 3 13 2 16 16 9 0 9 1 15 13 1 9 9 2 3 3 1 9 15 2 1 15 0 13 2
42 1 0 13 2 16 9 9 7 9 2 1 16 13 1 0 9 2 13 9 9 1 15 7 9 15 2 3 9 7 9 2 1 9 9 7 9 2 16 9 13 9 2
34 3 3 1 9 9 13 15 9 9 13 2 16 13 1 9 2 15 15 0 13 2 1 15 15 9 9 13 2 16 15 3 9 13 2
18 13 7 1 0 15 9 0 3 0 7 1 10 9 7 1 10 9 2
34 7 3 9 0 13 2 16 13 1 9 0 2 15 9 3 13 0 15 15 9 7 9 2 3 13 13 1 9 7 1 13 1 9 2
20 7 9 9 3 15 13 1 9 9 15 9 16 13 1 10 9 0 1 15 2
16 3 3 1 9 9 13 9 9 9 2 7 3 15 0 13 2
38 0 13 1 9 9 0 2 1 15 3 15 13 9 9 7 9 2 7 9 2 16 9 7 9 1 0 7 9 0 1 0 2 7 9 0 1 0 2
15 3 13 16 15 9 1 9 9 13 13 1 9 1 9 2
8 7 9 3 13 13 9 0 2
8 3 7 9 9 0 13 13 2
15 16 9 0 13 3 13 1 9 15 13 1 9 9 13 2
45 16 9 0 3 13 1 9 9 2 7 1 9 9 2 15 15 1 9 9 13 2 7 13 1 9 13 1 9 15 9 9 2 1 16 1 9 13 1 9 9 1 13 9 0 2
20 7 3 13 2 16 9 9 0 15 9 1 9 13 13 2 7 0 7 0 2
12 3 3 16 15 9 13 2 7 16 0 13 2
21 1 0 13 2 16 9 9 10 3 13 9 0 13 2 15 3 13 9 0 9 2
13 16 13 1 15 16 1 9 13 9 9 1 9 2
29 7 15 9 0 13 15 15 9 9 13 13 2 16 0 0 7 0 13 3 13 2 7 1 15 13 15 0 13 2
26 16 9 0 9 3 13 1 9 9 15 13 9 2 7 1 9 9 1 9 13 2 16 13 9 0 2
20 1 0 13 1 9 9 1 0 9 2 3 13 1 9 13 2 7 0 13 2
11 7 13 13 2 9 1 0 9 13 9 2
9 0 13 2 9 13 1 0 9 2
9 0 13 2 9 1 0 9 13 2
8 12 3 9 1 9 0 13 2
18 15 3 13 3 13 2 16 13 9 15 9 7 3 9 13 15 9 2
17 7 3 13 9 9 13 2 9 13 9 9 7 13 1 15 9 2
27 7 3 1 10 9 13 9 1 9 1 9 2 0 13 9 15 15 9 3 13 16 15 15 9 9 13 2
19 7 15 13 9 1 9 0 3 2 7 3 16 9 13 2 15 0 13 2
23 3 2 1 9 3 13 13 9 9 2 16 13 4 2 3 13 9 13 16 16 9 0 2
7 3 7 3 1 9 9 2
35 16 0 9 9 1 9 2 1 16 1 15 13 13 9 15 1 9 2 13 1 9 9 2 7 9 15 1 9 13 1 9 9 0 13 2
20 7 3 1 9 0 2 1 15 15 9 13 1 9 13 2 13 9 9 0 2
7 3 7 16 9 1 9 2
20 1 0 13 2 16 9 13 2 3 9 2 13 9 1 12 9 16 9 15 2
16 7 9 13 13 1 9 13 9 3 16 9 2 7 16 9 2
12 16 3 13 16 9 13 9 2 7 3 13 2
10 15 3 9 15 13 13 16 13 3 2
10 16 12 9 0 3 13 13 1 15 2
20 1 0 13 2 16 9 3 13 1 9 16 1 9 2 7 16 9 1 9 2
18 1 0 13 2 16 9 15 13 1 15 9 2 3 13 16 1 9 2
11 3 13 16 1 3 9 0 9 3 13 2
27 13 13 2 16 9 1 9 10 0 9 3 13 13 7 3 9 16 1 0 2 7 1 0 9 9 13 2
15 7 15 13 2 16 13 1 9 0 15 13 0 9 9 2
17 3 3 15 13 3 0 2 3 13 0 2 16 0 13 1 9 2
54 1 0 13 2 16 16 9 1 9 15 9 13 0 1 10 9 2 16 9 2 16 13 9 9 2 15 7 13 1 12 9 13 15 2 16 9 2 3 3 9 1 10 9 0 9 0 13 9 9 2 9 7 9 2
27 1 0 13 2 16 15 9 7 13 2 13 15 13 13 0 2 7 1 9 3 2 7 1 9 7 9 2
11 7 15 13 9 1 9 1 9 7 9 2
8 16 13 3 1 9 15 9 2
21 7 3 9 15 9 13 13 9 9 1 9 0 9 2 1 15 13 9 0 0 2
40 7 1 15 9 15 9 3 13 1 9 1 9 2 7 9 13 1 9 13 1 9 2 16 9 1 15 13 2 13 0 1 0 9 9 2 1 15 9 13 2
20 7 16 15 9 13 0 2 13 1 9 3 13 7 13 1 15 7 1 15 2
22 7 15 13 9 0 9 2 1 15 13 9 0 7 13 16 1 15 13 1 9 10 2
32 7 16 10 9 13 1 9 2 15 13 9 7 13 9 9 2 3 9 13 1 15 15 13 1 15 9 9 2 16 1 0 2
26 1 3 9 9 13 0 2 7 1 0 2 13 16 15 9 13 1 9 3 13 7 0 16 1 0 2
11 15 7 13 9 15 13 1 9 9 9 2
16 15 0 13 2 15 9 13 2 1 15 13 9 0 7 0 2
14 15 0 15 13 13 9 2 7 15 13 1 13 9 2
12 9 3 15 13 9 2 1 15 9 13 0 2
64 1 0 13 2 16 16 1 9 0 2 1 15 9 3 13 1 9 2 16 9 13 9 2 7 9 13 2 7 9 9 13 1 9 1 9 9 15 13 2 3 3 9 2 15 13 0 9 2 13 0 9 13 9 2 7 1 15 13 2 3 9 7 9 2
34 3 2 15 13 9 2 0 13 9 13 1 9 2 16 9 9 9 13 2 16 16 13 12 9 9 2 9 13 1 15 9 3 13 2
17 3 3 13 13 9 9 13 1 9 0 16 9 0 1 9 0 2
17 1 13 7 1 9 0 2 15 1 9 9 13 9 1 15 13 2
6 7 0 3 1 9 2
26 15 3 13 9 12 9 2 15 13 12 9 0 2 15 16 0 9 1 0 9 13 2 16 13 9 2
10 7 9 9 13 12 9 1 10 9 2
26 3 2 1 9 13 2 16 1 9 0 0 13 10 9 2 1 9 13 13 4 1 9 9 7 9 2
15 15 1 15 13 0 9 10 2 13 0 9 1 15 9 2
12 16 16 13 15 9 1 9 2 13 0 13 2
14 7 1 9 15 13 1 10 9 2 3 13 15 9 2
9 16 9 9 9 13 1 9 9 2
11 16 16 9 13 9 2 3 9 13 9 2
14 7 9 0 15 13 1 9 2 3 13 1 9 9 2
13 16 16 13 1 9 12 2 13 15 9 9 15 2
55 15 7 9 9 13 13 1 8 9 7 9 7 1 0 15 9 2 1 15 16 1 9 2 3 1 15 13 2 13 1 9 1 10 9 2 7 13 13 1 0 3 2 13 16 1 16 13 1 12 13 1 9 1 15 2
59 3 1 3 13 15 9 0 0 15 9 9 1 9 15 9 13 2 16 3 13 0 2 16 9 13 2 16 9 0 15 2 3 0 2 3 13 15 0 2 16 13 1 12 9 7 9 2 13 16 1 15 15 13 1 9 0 9 9 2
27 7 13 13 2 16 9 16 13 1 9 9 2 15 9 13 2 3 16 15 13 1 15 9 1 15 9 2
15 3 3 13 9 16 1 9 9 2 1 15 13 1 9 2
28 3 2 1 9 0 1 15 13 13 1 9 1 10 9 0 2 3 13 15 15 9 13 16 1 9 10 9 2
24 3 3 12 9 13 1 9 2 3 16 13 0 7 3 9 2 13 9 1 9 15 0 0 2
15 9 3 1 9 9 13 2 3 13 1 9 1 9 9 2
30 3 16 9 9 13 0 2 3 3 2 13 1 9 0 2 3 13 15 9 15 2 16 3 1 15 13 10 15 9 2
41 7 3 16 13 16 9 9 1 10 9 2 15 9 9 13 2 3 13 16 9 13 1 9 0 2 13 1 9 1 9 9 2 7 13 1 9 1 9 9 0 2
12 0 3 9 15 13 1 9 13 1 9 0 2
24 1 0 3 13 13 2 16 1 9 2 13 10 3 13 1 9 9 2 7 3 1 9 9 2
27 7 16 9 3 13 9 2 3 16 9 9 9 9 13 2 0 13 4 9 0 2 7 3 1 9 13 2
7 3 0 9 3 9 13 2
19 3 2 16 15 9 9 15 13 2 7 13 9 9 13 2 7 9 0 2
8 3 13 16 13 9 9 0 2
13 16 13 2 16 3 13 15 15 9 2 7 15 2
14 7 1 15 0 9 13 1 9 0 2 13 4 9 2
18 3 13 9 15 13 1 9 15 12 9 2 16 13 1 9 15 0 2
9 7 1 2 10 9 13 1 9 2
15 16 3 9 0 13 1 9 9 2 13 16 9 15 13 2
20 3 2 16 15 13 9 0 1 0 9 2 3 15 13 9 0 1 9 0 2
9 3 0 13 13 9 1 10 9 2
25 1 16 13 9 9 2 9 0 13 15 1 15 0 13 9 9 0 2 15 13 13 1 10 9 2
15 16 10 9 15 13 9 2 13 0 1 9 7 9 9 2
47 7 3 2 16 10 9 13 1 9 2 15 9 0 13 0 2 16 13 9 1 12 8 2 1 9 3 2 16 13 15 13 9 0 15 3 15 13 1 10 9 16 15 13 9 1 9 2
29 7 16 9 0 3 13 2 3 13 15 9 9 9 10 2 3 3 13 1 10 9 2 16 13 9 1 10 8 2
17 3 16 13 12 9 2 13 15 2 1 16 9 12 13 9 15 2
12 7 3 13 0 9 2 13 15 13 15 9 2
23 15 3 13 15 13 15 1 12 9 2 13 12 9 10 0 9 13 2 7 15 1 15 2
29 15 0 13 15 1 0 9 2 3 3 13 1 3 2 7 15 9 13 2 15 9 9 1 9 7 9 13 4 2
12 15 3 13 9 15 0 15 1 12 9 13 2
32 7 16 1 0 9 13 13 2 13 15 9 3 13 12 12 9 2 7 15 15 15 13 1 9 1 15 2 16 0 1 9 2
9 16 9 9 15 13 1 9 0 2
17 16 2 1 9 2 0 9 15 13 1 9 2 13 1 9 9 2
24 3 3 13 15 9 0 1 9 0 7 9 9 2 16 13 0 0 1 9 0 7 9 9 2
24 7 3 2 1 3 0 9 13 4 2 13 3 3 1 0 9 9 13 15 9 1 9 9 2
31 16 9 13 1 9 9 9 9 2 13 12 0 9 2 7 3 1 9 0 13 4 9 0 0 2 7 3 9 0 13 2
17 7 15 9 9 13 2 16 10 9 0 13 9 0 1 9 9 2
9 3 13 10 15 9 0 13 9 2
18 3 15 13 16 1 15 9 1 9 2 9 13 9 7 9 7 9 2
43 7 3 13 9 15 0 2 15 13 9 1 9 12 9 2 13 15 13 2 16 0 9 4 13 1 0 9 0 2 7 16 10 9 0 9 0 9 1 9 9 13 4 2
40 7 15 13 0 13 2 16 13 13 9 9 2 15 13 9 1 13 13 1 9 0 3 1 0 9 2 13 7 3 1 0 2 3 3 1 9 0 7 0 2
20 3 0 13 9 13 1 9 0 1 15 16 13 9 0 7 0 1 15 9 2
26 3 15 9 15 9 13 2 0 13 2 3 12 1 9 9 2 7 1 9 9 2 3 1 9 0 2
13 1 0 13 2 16 3 13 9 12 2 7 0 2
21 3 3 9 9 13 2 16 15 13 9 0 7 0 9 9 2 1 15 0 13 2
25 1 0 13 2 16 9 0 13 13 9 9 0 1 9 2 15 16 9 13 9 2 16 9 13 2
35 7 3 13 9 9 7 9 1 9 3 2 16 13 9 1 9 9 2 9 3 1 10 9 0 13 1 9 2 1 13 3 9 0 2 2
14 9 0 1 9 9 2 16 0 13 3 0 7 0 2
17 7 0 9 0 9 13 2 16 13 9 2 1 15 9 0 13 2
18 7 1 15 13 13 13 2 16 1 9 13 1 9 0 9 7 9 2
35 16 13 1 9 9 0 2 3 13 13 9 9 3 13 0 9 9 2 16 1 12 9 13 13 15 0 9 2 16 1 12 9 0 9 2
11 16 9 13 0 7 0 2 1 9 9 2
8 7 0 16 9 13 9 9 2
12 0 2 16 9 13 9 1 15 13 9 9 2
43 16 3 9 13 9 1 9 0 13 2 16 1 12 8 13 2 3 13 9 2 7 9 15 1 9 9 15 13 2 2 3 1 9 13 9 1 9 9 2 13 0 13 2
17 7 1 15 9 9 1 0 1 9 13 2 16 9 13 9 0 2
23 1 0 13 2 16 1 9 9 9 9 13 4 3 1 9 0 2 15 13 1 9 0 2
32 7 1 9 9 13 9 0 1 9 2 16 13 1 9 2 16 13 2 16 9 0 9 0 9 13 2 7 1 9 15 13 2
21 1 3 9 0 13 1 9 9 1 9 7 9 2 13 16 9 9 13 3 13 2
23 7 1 9 0 9 13 9 2 7 15 9 0 1 15 2 7 9 0 15 2 1 15 2
19 16 3 9 13 16 9 3 13 9 0 9 2 16 1 9 13 13 9 2
14 3 13 16 9 15 1 15 13 2 3 13 9 0 2
13 7 16 9 0 9 13 9 2 3 13 16 0 2
53 7 3 13 15 2 15 13 13 15 2 16 9 13 9 0 2 13 9 13 7 0 1 9 2 7 16 2 16 9 2 13 9 0 15 9 2 7 1 15 13 1 16 3 1 9 13 2 15 15 9 13 9 2
15 1 0 13 2 16 9 0 2 13 1 9 1 9 9 2
29 7 3 13 16 9 15 1 9 1 9 13 2 9 9 13 2 7 1 9 0 13 2 16 13 1 9 15 9 2
21 16 3 9 9 13 1 9 0 9 2 1 16 13 1 9 9 0 1 15 13 2
31 7 1 9 3 13 0 2 16 7 9 0 2 0 1 9 13 3 9 13 2 16 9 3 13 1 9 13 13 9 0 2
17 1 0 13 2 16 9 9 0 1 9 9 1 10 9 0 13 2
23 3 2 1 9 2 9 13 15 13 1 9 13 16 15 1 9 2 7 16 9 1 9 2
24 3 0 9 1 15 13 13 2 13 1 16 9 13 1 9 9 2 16 13 9 1 12 8 2
11 7 9 0 13 15 9 13 9 9 0 2
19 3 13 16 9 9 13 1 9 0 15 2 7 3 1 15 13 1 9 2
18 1 9 7 9 0 2 16 9 0 13 9 9 2 3 3 13 9 2
21 7 0 9 13 13 15 13 9 2 7 0 13 13 13 2 16 13 1 12 8 2
34 15 9 9 13 2 16 9 1 15 13 9 0 2 15 3 13 16 0 13 1 9 0 9 9 2 7 1 15 15 1 9 9 13 2
21 7 3 13 13 9 1 15 13 9 0 13 1 9 2 7 15 13 13 9 9 2
22 7 1 3 13 13 9 0 9 15 7 9 2 16 13 15 9 2 16 9 15 13 2
18 7 3 9 2 15 13 9 0 2 13 9 13 2 3 9 7 9 2
24 1 15 7 13 13 2 16 13 2 0 9 2 15 13 9 3 0 2 13 9 13 7 13 2
19 9 7 9 2 15 13 9 3 0 2 16 0 13 4 2 13 9 0 2
62 1 0 3 13 2 16 2 16 9 13 1 12 9 7 9 2 9 9 13 0 2 3 16 9 15 0 13 15 9 0 2 7 16 15 9 0 13 15 9 16 15 9 13 4 13 1 15 9 2 3 13 9 13 15 9 0 2 16 13 1 15 2
13 9 3 3 3 13 1 9 2 7 3 1 9 2
9 7 3 3 13 15 9 13 15 2
12 3 2 15 9 13 9 0 1 9 10 9 2
23 7 9 3 1 0 9 9 0 13 2 15 13 1 9 2 15 15 9 1 9 9 13 2
21 1 0 13 2 16 16 9 7 9 3 13 9 0 9 2 3 7 9 7 9 2
20 7 3 16 9 9 0 1 9 9 13 2 3 3 1 15 1 0 9 13 2
14 3 13 16 3 13 13 9 9 7 9 1 15 9 2
32 1 9 7 9 2 15 13 9 0 2 15 13 15 2 13 9 13 1 9 0 2 1 15 13 9 0 2 15 0 9 13 2
41 7 1 15 9 10 9 0 13 1 9 15 13 1 9 2 16 9 13 2 12 1 8 2 8 12 2 1 8 2 7 9 1 12 8 2 16 9 9 1 9 2
13 1 0 13 2 16 0 13 15 1 15 9 13 2
10 7 13 16 15 9 3 0 13 15 2
23 13 9 9 2 15 13 0 0 15 16 13 0 1 9 7 0 1 9 2 1 9 13 2
24 1 0 13 2 16 15 9 15 10 9 13 2 3 13 15 0 2 7 0 9 2 7 9 2
25 3 13 9 16 9 15 13 1 9 2 13 13 9 2 15 16 1 15 9 13 15 1 9 13 2
9 9 3 13 1 9 2 3 0 2
26 9 7 0 0 13 2 3 1 15 9 1 15 13 2 7 1 9 1 9 2 16 13 1 12 8 2
8 3 13 1 9 7 9 13 2
19 7 10 15 1 15 13 9 9 7 13 9 2 13 1 9 7 9 13 2
12 7 3 3 13 13 9 0 2 7 9 13 2
8 16 9 13 9 15 9 13 2
9 7 1 9 0 9 9 13 0 2
11 3 1 15 9 13 0 2 0 0 9 2
14 3 2 9 0 3 13 9 0 2 16 7 9 9 2
14 7 10 15 13 9 2 13 3 0 9 13 9 9 2
15 1 3 9 13 9 0 2 13 16 1 9 13 3 13 2
8 7 15 13 0 9 7 9 2
24 1 3 9 13 9 9 2 13 16 7 1 15 9 10 13 9 9 2 7 1 9 9 10 2
17 16 15 15 1 15 13 9 0 2 3 13 13 9 7 9 15 2
26 10 7 9 1 9 9 13 9 0 2 16 13 0 9 0 9 7 9 2 16 1 12 1 9 13 2
29 16 7 1 9 9 10 13 9 9 2 1 15 13 1 9 2 7 3 1 15 15 13 9 15 2 13 12 9 2
25 12 13 16 12 9 9 13 9 0 9 2 3 9 0 2 7 9 0 2 1 15 9 9 13 2
64 7 3 13 9 0 15 9 9 13 2 3 1 9 7 15 13 2 16 1 2 8 12 1 9 2 7 1 12 2 8 12 2 1 15 9 13 4 2 15 3 9 9 1 15 9 3 13 2 16 3 13 13 0 16 1 9 10 2 7 13 1 9 9 2
13 7 1 15 13 16 13 3 13 9 16 1 9 2
43 7 16 15 15 13 0 2 3 13 15 9 15 13 9 9 15 2 7 15 10 9 2 3 15 15 13 0 2 3 13 15 9 15 13 9 9 15 2 7 15 10 13 2
13 1 9 3 13 13 9 2 15 13 9 9 15 2
38 3 7 13 9 13 15 15 3 13 15 7 9 9 10 2 16 9 0 13 9 15 13 9 9 15 2 16 13 15 9 3 9 2 16 9 13 9 2
14 15 3 9 13 1 13 1 9 9 2 16 9 0 2
22 7 9 2 16 1 12 1 9 13 2 3 13 9 0 2 1 3 13 9 9 15 2
13 15 1 15 10 9 13 2 16 13 10 9 0 2
25 16 3 9 13 1 9 9 2 16 13 15 0 2 13 16 9 0 1 15 13 2 3 4 13 2
30 15 13 16 13 15 9 13 9 1 9 0 7 1 9 0 2 16 3 13 16 13 15 2 7 3 16 13 9 0 2
22 7 3 2 16 9 0 3 13 0 1 9 15 13 2 3 7 9 0 2 16 13 2
31 16 16 13 9 10 0 0 2 3 13 13 0 1 15 15 13 1 9 15 2 1 15 13 2 16 9 0 1 9 13 2
14 1 9 7 15 3 13 9 9 2 15 9 9 13 2
23 7 3 13 13 16 9 0 9 13 1 9 2 16 7 15 9 9 13 1 9 10 9 2
14 7 1 13 2 16 0 13 0 9 13 12 9 9 2
8 7 9 0 13 9 15 9 2
9 3 2 9 13 9 9 7 9 2
24 7 13 9 0 15 13 1 9 1 13 10 9 13 2 16 9 13 1 9 1 13 10 9 2
16 7 3 15 15 13 9 0 2 13 9 2 7 9 1 9 2
30 7 3 15 13 2 16 9 0 15 15 13 16 9 0 2 1 16 4 13 16 13 1 15 9 15 4 13 1 9 2
51 13 3 2 16 9 1 9 2 15 13 0 2 13 12 1 10 2 7 0 2 7 13 3 13 1 9 13 7 0 2 3 16 9 13 13 16 9 15 2 7 1 9 9 0 13 3 1 15 9 13 2
23 1 3 13 9 1 9 13 1 9 10 2 13 16 9 13 13 9 1 9 16 9 15 2
32 16 13 16 9 9 0 15 13 2 13 1 0 1 9 2 7 1 9 2 1 15 9 15 3 13 1 9 0 16 9 15 2
10 16 9 9 0 13 1 15 9 13 2
20 7 13 16 9 13 3 15 13 1 0 16 9 15 2 7 16 9 1 9 2
21 7 9 13 13 1 9 2 13 16 9 9 0 2 1 15 12 13 9 1 9 2
31 0 2 16 13 16 3 13 0 16 16 9 13 13 0 7 13 0 2 3 9 0 2 16 9 13 0 2 3 9 0 2
65 13 3 2 16 1 9 13 15 13 1 9 0 3 16 9 1 9 2 15 9 16 1 15 3 13 12 0 2 9 15 1 15 13 1 15 15 13 0 1 13 9 2 3 1 9 13 2 15 12 9 13 13 9 2 15 13 1 15 2 7 1 15 9 0 2
25 0 2 16 2 16 13 4 2 9 15 13 9 9 0 2 3 13 15 9 1 9 7 1 9 2
46 7 3 2 13 10 13 9 2 13 1 9 2 9 0 13 3 13 1 9 2 7 1 9 3 13 2 7 1 0 0 13 2 7 13 1 9 9 1 0 9 2 16 15 9 0 2
33 3 3 13 16 12 9 13 13 13 1 9 9 10 9 0 2 15 13 9 0 2 7 13 9 9 10 15 2 15 13 9 13 2
18 15 3 13 13 10 9 0 2 1 15 13 16 1 16 13 1 9 2
24 1 0 3 13 2 16 9 3 13 13 9 0 16 13 9 9 16 9 0 3 1 9 0 2
30 1 3 1 9 9 1 9 9 13 13 2 3 9 13 0 2 7 3 13 9 2 3 3 13 13 9 1 9 9 2
11 7 9 1 9 0 2 15 13 0 9 2
16 1 7 13 1 15 9 0 15 3 13 3 9 15 13 9 2
15 7 9 13 9 9 0 2 16 15 15 0 9 9 13 2
41 3 16 1 9 13 4 2 13 15 7 13 0 1 9 2 7 3 10 9 9 13 1 9 9 2 7 16 13 12 3 9 2 7 3 13 9 13 1 13 9 2
30 1 3 9 9 13 3 13 13 16 1 16 13 9 16 9 15 2 16 13 4 2 13 16 3 13 13 16 1 9 2
38 1 15 3 13 16 1 9 0 13 0 7 9 0 2 13 15 9 9 2 1 15 9 15 9 9 13 13 2 7 1 15 7 9 13 9 9 13 2
16 7 3 13 9 9 2 7 9 10 13 1 13 15 1 9 2
7 15 3 9 13 15 0 2
17 7 9 9 0 13 1 9 0 1 9 13 2 15 9 9 13 2
14 7 15 13 13 1 15 9 0 2 13 0 7 0 2
6 9 0 0 9 13 2
30 16 15 13 9 0 16 1 9 0 2 15 16 9 9 13 0 0 2 15 9 10 9 13 2 7 1 9 0 13 2
17 16 15 9 3 13 9 0 9 0 2 7 15 9 13 9 15 2
32 1 0 3 13 2 16 9 15 13 9 0 2 3 13 15 9 1 9 15 13 9 0 2 16 13 0 15 1 10 9 0 2
18 16 3 1 9 9 9 0 13 2 3 3 1 9 9 9 0 13 2
37 16 0 9 9 9 13 2 1 15 15 13 13 16 15 13 15 0 3 13 2 13 16 15 9 13 1 9 9 9 15 0 1 9 9 3 13 2
34 15 7 15 13 3 13 16 7 1 9 15 9 1 9 9 2 15 9 1 9 15 13 2 7 1 15 16 15 9 4 1 0 13 2
29 7 3 13 16 1 9 15 9 2 7 1 0 13 2 7 1 9 15 9 13 2 1 9 9 9 9 13 4 2
17 16 9 0 3 13 9 15 13 2 7 1 15 1 9 0 13 2
14 7 9 3 13 9 1 9 9 2 7 1 9 9 2
26 3 16 1 9 9 13 9 0 1 9 2 3 3 1 9 1 9 0 13 13 10 9 7 9 0 2
29 7 16 2 16 9 13 2 15 15 13 13 13 13 9 2 9 13 1 9 3 13 9 7 9 0 1 15 13 2
30 16 1 9 9 3 13 2 7 1 9 13 13 2 9 9 3 13 1 13 9 15 9 13 2 7 13 1 9 13 2
30 9 7 2 15 15 9 9 13 2 3 0 9 7 9 0 9 13 2 7 3 9 13 15 15 15 1 9 13 13 2
5 0 1 9 9 2
11 16 9 15 13 9 2 3 13 15 0 2
8 9 7 0 15 0 13 13 2
24 9 7 9 1 16 1 9 0 13 2 0 13 13 2 15 16 15 13 0 9 0 9 13 2
16 15 3 13 2 16 9 9 3 13 1 9 16 13 9 9 2
19 3 16 13 15 9 9 1 15 9 13 9 2 7 1 15 9 13 9 2
9 15 3 9 0 0 9 0 13 2
13 16 1 15 9 13 9 15 9 1 13 9 0 2
14 16 10 9 15 13 1 15 9 0 2 13 9 0 2
14 15 13 1 9 9 0 2 16 13 1 12 1 9 2
40 7 3 2 1 10 9 13 15 9 2 7 0 13 12 9 13 0 9 0 2 13 2 16 0 9 0 13 9 13 15 9 0 2 16 0 13 13 9 0 2
20 7 3 3 13 15 9 15 9 13 9 2 7 15 13 9 2 16 9 13 2
20 7 16 9 13 1 12 8 9 3 13 9 7 9 0 1 9 7 0 9 2
13 15 3 13 1 13 9 9 1 9 7 1 9 2
24 7 3 13 16 9 13 1 9 13 9 9 13 1 9 13 2 7 3 1 9 13 3 13 2
11 16 1 9 9 0 3 0 13 9 0 2
30 3 15 13 2 16 1 10 9 2 1 9 2 1 9 9 13 2 13 15 9 13 1 9 0 2 1 15 3 9 2
27 7 3 3 13 1 15 13 1 9 2 16 13 9 0 15 13 9 0 1 13 2 16 3 13 9 0 2
20 16 16 9 13 1 9 9 2 15 3 9 9 3 13 0 2 7 0 3 2
11 15 3 9 9 9 13 2 7 9 9 2
9 3 7 9 13 1 9 7 9 2
30 7 16 9 0 13 9 0 0 1 9 1 0 0 2 16 9 7 9 2 7 9 9 2 7 9 9 2 7 3 2
51 1 0 13 2 16 9 0 13 9 13 2 3 16 13 13 13 1 9 1 9 9 0 2 3 13 1 9 9 2 7 1 9 15 2 1 16 13 9 2 7 1 9 15 3 9 0 1 9 13 13 2
26 7 16 1 9 9 13 9 1 9 9 2 7 1 9 13 9 0 2 1 15 15 9 1 9 13 2
28 3 2 16 13 9 1 12 8 2 0 13 16 13 0 9 15 12 9 13 1 9 9 2 7 15 1 9 2
14 16 1 9 9 9 9 3 13 16 1 16 13 9 2
27 13 3 2 16 15 13 2 16 9 7 9 13 12 13 2 1 15 3 13 12 2 16 13 9 0 9 2
12 7 9 0 13 9 15 9 15 13 9 0 2
30 1 3 9 0 13 9 10 9 0 2 13 16 1 9 15 9 13 0 9 1 9 2 0 0 9 0 15 13 13 2
10 7 1 9 2 16 9 0 9 13 2
17 3 1 9 0 13 9 0 2 3 13 15 9 1 9 0 13 2
15 16 15 3 13 16 1 15 16 9 13 9 1 15 9 2
17 9 7 0 3 13 15 1 9 2 1 0 13 2 7 9 13 2
21 7 13 9 0 2 15 13 13 1 9 9 2 16 15 9 0 2 16 13 4 2
15 7 16 9 1 15 9 13 1 9 1 9 1 9 13 2
14 7 16 1 9 13 9 2 16 13 9 1 9 9 2
11 7 0 9 13 3 1 10 1 9 0 2
24 0 7 13 3 2 1 9 2 1 10 9 0 2 16 15 13 10 9 0 13 1 9 13 2
20 7 1 9 7 9 2 9 0 0 13 1 0 9 2 7 9 0 1 0 2
9 16 3 0 9 13 2 7 9 2
25 3 13 3 9 0 2 13 1 12 9 2 7 15 13 1 0 9 9 2 7 15 13 1 9 2
23 1 0 13 2 16 9 0 7 1 9 13 13 2 7 13 9 0 2 3 1 9 13 2
29 7 3 3 13 13 1 15 9 15 0 9 13 1 15 1 9 9 15 13 1 9 2 16 13 1 15 9 0 2
22 0 1 15 15 13 1 8 1 9 2 16 9 0 13 9 13 13 2 16 13 9 2
18 7 1 15 13 9 2 13 9 0 7 10 15 9 0 1 15 9 2
10 16 1 0 9 9 13 1 9 9 2
10 3 1 9 9 13 13 9 1 9 2
41 15 3 9 9 13 9 0 3 1 9 9 13 2 15 13 10 13 2 16 1 9 9 0 15 13 10 13 2 7 15 13 9 0 13 1 15 13 9 0 0 2
13 16 10 9 0 13 13 2 16 1 12 8 13 2
15 15 15 13 3 9 7 3 15 15 2 3 13 13 9 2
17 3 1 12 8 9 13 16 9 9 3 13 9 1 9 15 0 2
32 7 0 1 15 16 1 0 15 13 13 16 9 0 2 16 9 7 9 15 9 3 13 9 13 2 1 15 13 1 10 9 2
20 7 3 13 13 2 16 15 9 1 9 0 7 15 9 0 13 3 1 9 2
12 16 13 9 10 9 0 13 1 9 13 13 2
10 3 9 0 2 16 9 9 7 9 2
46 15 0 2 16 9 7 9 15 2 15 13 9 15 0 1 9 9 13 9 9 0 2 13 3 9 0 7 0 1 9 13 2 15 16 9 9 0 3 13 15 0 2 7 15 9 2
24 3 13 16 13 7 13 1 9 13 13 1 9 7 9 2 7 3 9 3 2 7 9 13 2
41 7 1 15 13 9 1 12 8 2 7 1 15 9 13 1 12 1 9 2 9 0 7 0 3 1 0 13 2 13 15 13 9 0 1 15 16 9 13 13 9 2
16 15 0 9 13 1 15 9 2 7 16 15 1 15 13 13 2
11 7 3 13 10 9 13 1 9 0 13 2
31 1 0 16 13 1 9 9 0 13 1 10 10 9 2 13 1 15 9 15 0 16 9 15 3 13 1 9 16 1 9 2
12 16 7 13 2 13 9 13 15 9 7 9 2
44 15 7 9 3 13 0 1 9 9 16 13 9 7 9 13 1 9 9 2 3 3 13 9 1 0 9 2 2 7 13 9 0 2 16 13 9 9 1 9 9 13 9 9 2
23 15 7 9 13 9 0 2 3 1 9 9 16 1 9 9 2 16 9 15 15 9 13 2
14 7 3 7 9 0 7 15 9 0 1 9 15 13 2
14 16 13 16 9 0 1 9 9 13 2 16 9 13 2
34 7 0 13 2 16 1 9 9 0 13 9 0 7 15 9 0 1 16 1 15 16 9 13 9 9 2 7 15 0 9 7 15 9 2
16 7 1 10 9 13 9 1 15 16 9 15 1 3 9 13 2
18 7 9 7 9 13 12 9 2 1 9 13 9 2 15 1 15 13 2
10 3 3 13 13 9 9 1 9 9 2
13 7 9 13 9 9 2 16 1 12 1 9 13 2
25 16 13 2 16 9 3 13 9 7 9 2 7 1 9 3 13 16 13 9 2 7 16 13 9 2
14 7 9 13 9 1 9 10 2 7 1 15 9 10 2
28 16 0 9 2 3 1 12 9 3 13 0 9 2 16 9 1 9 3 13 16 13 9 2 9 10 3 13 2
44 16 7 0 9 2 1 1 9 7 9 3 13 12 15 13 9 16 16 9 13 9 9 2 13 16 9 13 9 1 9 2 7 3 13 15 1 9 9 2 15 13 3 0 2
20 7 3 1 9 2 1 3 13 9 1 15 13 2 7 9 15 1 15 0 2
11 7 1 9 13 3 13 9 13 1 9 2
16 3 13 15 9 15 13 15 9 2 1 10 9 0 0 13 2
20 7 15 9 13 9 1 12 1 9 2 13 16 9 13 9 9 7 9 15 2
24 13 7 16 13 9 13 9 13 2 7 13 9 13 9 2 16 15 9 1 9 13 0 9 2
13 3 15 9 3 13 13 9 7 9 16 15 9 2
22 7 16 9 13 9 1 9 9 1 9 2 3 9 9 1 15 9 13 1 15 9 2
21 7 16 9 1 15 13 2 7 3 2 15 9 13 1 9 0 15 9 7 15 2
44 16 3 13 9 15 15 9 13 0 7 3 13 2 1 15 9 9 9 13 1 15 16 13 15 9 2 13 16 1 9 9 9 3 9 13 2 1 15 16 0 1 15 13 2
18 7 3 15 9 13 1 10 9 2 7 3 9 13 9 2 9 13 2
36 16 0 9 3 13 9 0 1 15 13 2 7 13 1 9 9 2 3 1 15 9 13 9 2 13 16 9 3 9 13 2 7 1 9 13 2
25 1 0 13 2 16 2 16 13 9 1 12 1 9 2 9 3 15 9 13 9 1 15 9 0 2
29 7 3 13 9 3 13 1 9 9 16 15 9 2 15 3 13 16 1 9 9 2 7 15 9 13 16 13 9 2
23 1 0 13 2 16 9 0 1 15 9 13 13 9 7 15 15 2 1 16 13 9 0 2
54 7 15 13 2 16 9 13 0 13 2 3 1 16 13 9 2 7 1 16 13 9 2 3 13 13 3 1 0 15 1 15 13 2 16 15 13 9 10 7 15 15 13 9 2 16 3 13 9 13 15 16 9 9 2
13 3 3 1 15 16 13 9 13 16 1 9 13 2
30 1 9 7 0 9 0 13 3 13 2 1 1 0 13 2 15 13 9 9 1 9 2 1 9 9 13 1 15 9 2
29 1 0 3 13 2 16 9 15 13 2 16 9 9 13 1 9 9 2 7 3 1 9 9 2 15 9 0 13 2
34 0 2 1 9 0 15 13 3 0 1 9 13 2 3 13 13 13 12 9 0 16 9 13 1 12 15 9 16 12 13 0 7 13 2
23 13 13 2 16 1 15 9 13 12 13 2 3 9 15 13 9 2 7 0 15 13 9 2
37 1 10 3 13 9 1 15 13 9 9 2 9 15 13 16 0 7 9 13 2 7 9 15 13 16 9 7 9 13 2 16 1 12 1 9 13 2
24 7 1 9 0 0 13 1 9 9 13 2 7 1 15 9 13 16 13 9 1 9 9 0 2
6 0 9 9 2 3 2
12 3 9 1 9 2 7 1 9 9 13 9 2
18 16 3 0 9 13 9 13 2 9 0 9 2 3 9 2 13 13 2
24 3 1 9 0 9 9 15 13 15 13 2 16 3 1 9 9 13 2 7 16 0 9 13 2
35 16 7 1 9 9 13 2 3 9 13 2 7 1 9 0 2 15 15 15 9 2 1 15 3 13 13 2 13 13 2 16 1 9 13 2
32 7 3 13 16 3 3 1 9 9 0 13 9 9 2 1 13 9 1 9 9 13 2 16 9 1 9 2 7 9 1 9 2
14 7 15 3 13 15 1 15 13 2 16 9 9 9 2
20 3 2 1 9 0 3 13 9 13 9 0 2 7 9 15 13 1 9 0 2
18 9 9 2 9 9 13 9 16 15 9 2 7 9 0 16 15 9 2
12 16 9 0 15 13 2 3 13 9 0 9 2
20 0 3 9 15 13 9 1 9 9 2 16 13 1 9 13 3 13 15 9 2
17 7 9 0 15 13 1 9 9 2 13 9 0 7 13 1 15 2
30 3 16 13 2 9 0 9 13 1 15 1 9 0 13 2 3 3 13 2 9 9 13 2 1 15 1 9 9 13 2
26 3 3 13 13 16 15 13 9 16 15 1 9 10 13 2 7 9 15 13 2 7 0 2 7 0 2
22 3 0 9 13 2 1 1 9 7 9 3 13 15 0 2 16 1 12 8 9 13 2
10 9 7 3 13 9 9 2 16 0 2
13 3 13 16 13 15 9 2 1 9 0 15 13 2
24 1 3 13 9 13 13 9 9 0 2 15 3 13 13 16 7 1 9 9 7 1 9 0 2
13 16 7 13 0 2 3 13 16 9 13 9 9 2
13 3 3 13 15 9 1 9 9 15 15 0 13 2
20 16 7 9 0 13 9 9 1 9 0 2 3 9 13 9 9 1 9 0 2
11 3 2 9 13 13 9 10 9 7 9 2
37 7 3 15 13 2 16 9 7 9 0 13 2 3 3 16 13 0 1 9 2 7 16 1 9 7 9 13 12 16 1 9 7 15 15 13 9 2
14 1 0 13 2 16 9 15 9 13 9 9 16 9 2
27 9 3 13 9 9 1 9 9 2 16 3 10 9 9 1 10 9 13 2 15 16 15 9 13 9 0 2
32 3 3 13 1 10 9 7 9 13 2 16 15 15 9 9 13 2 13 9 9 15 1 15 13 2 15 9 1 10 9 13 2
14 16 13 16 9 13 9 9 2 15 13 13 9 9 2
24 15 7 15 1 15 13 2 9 7 9 1 15 13 2 7 1 10 9 13 2 16 9 13 2
37 1 0 13 2 16 9 13 1 12 9 13 13 1 9 2 3 0 2 7 0 2 1 16 15 9 13 13 15 1 9 2 16 9 13 13 0 2
30 3 13 13 3 16 3 13 0 9 1 13 2 7 16 0 9 13 9 9 2 7 1 9 13 9 1 15 0 13 2
17 3 2 10 9 13 1 9 15 15 13 2 1 0 0 13 9 2
6 7 9 13 9 9 2
50 16 7 9 1 15 16 13 9 9 2 13 1 15 9 1 15 13 9 2 0 13 16 13 1 15 9 1 15 13 9 2 7 1 0 7 1 0 2 1 16 15 9 1 0 1 9 13 16 15 2
14 12 3 9 13 15 13 9 2 7 15 13 9 9 2
19 1 0 13 2 16 9 15 13 1 9 15 13 0 9 7 3 0 15 2
18 3 7 9 3 13 13 9 9 2 7 3 9 1 15 9 0 13 2
19 3 15 3 0 13 2 9 13 0 9 9 2 7 9 2 15 9 13 2
9 3 0 2 16 9 13 9 9 2
45 16 15 9 15 3 13 1 15 0 2 13 9 1 9 9 2 7 13 9 15 13 7 9 1 0 9 2 7 0 1 9 2 1 15 9 9 13 3 13 2 16 1 15 13 2
22 1 0 3 13 2 16 15 13 1 9 15 15 13 9 0 2 7 15 13 9 0 2
15 9 3 0 15 13 9 15 2 3 13 15 9 15 9 2
42 7 3 13 16 9 15 13 9 9 1 16 13 15 2 13 13 0 1 16 13 9 15 15 2 16 9 1 9 2 7 9 9 2 1 15 9 13 2 7 9 13 2
9 7 16 9 2 15 13 9 9 2
29 1 9 7 9 1 9 3 13 9 9 2 1 15 15 1 9 10 13 2 16 9 2 1 9 1 15 15 13 2
16 7 9 13 2 16 9 3 13 1 9 2 16 1 9 9 2
13 1 0 13 2 16 9 9 13 13 1 9 9 2
10 16 1 0 9 13 13 1 9 10 2
26 7 15 3 9 3 13 13 9 9 2 15 13 9 3 9 13 4 7 13 2 1 9 7 1 9 2
29 7 16 0 9 13 9 9 16 15 9 15 2 3 1 0 0 9 13 13 1 15 9 9 16 13 1 9 15 2
32 1 0 13 2 16 1 15 15 13 1 9 9 2 13 16 9 1 9 13 1 9 9 15 1 15 13 2 16 1 0 13 2
24 9 7 3 13 1 9 16 13 2 16 13 1 9 0 7 0 2 15 13 9 1 9 9 2
14 3 3 13 9 9 16 16 13 9 1 9 9 15 2
54 1 0 13 2 16 16 9 9 0 0 13 9 9 13 7 9 13 2 16 13 0 9 9 2 15 3 13 15 9 0 13 1 15 2 16 3 15 13 1 9 15 9 0 13 1 9 2 16 9 2 7 15 3 2
20 3 7 9 15 15 9 13 2 9 9 13 1 15 15 16 3 9 9 13 2
24 16 9 13 1 9 1 9 15 9 2 1 10 15 13 1 15 2 13 1 15 1 9 13 2
19 7 15 13 1 15 16 3 1 9 9 9 1 9 1 9 13 9 9 2
9 7 15 13 0 15 15 9 13 2
23 1 3 9 9 1 9 13 2 13 16 15 15 13 2 1 9 1 9 9 15 13 13 2
27 13 3 16 13 9 0 9 1 15 16 13 9 15 13 9 15 9 2 15 9 1 9 0 1 9 13 2
17 16 13 3 1 15 9 7 9 2 16 9 13 9 10 1 9 2
17 13 3 16 9 0 2 3 1 15 13 2 13 10 9 7 9 2
15 3 0 15 13 1 13 10 9 2 16 1 13 10 9 2
55 1 3 9 13 7 10 15 9 1 9 9 9 13 2 15 16 13 9 1 9 13 9 15 15 13 2 16 1 12 8 13 2 13 16 9 0 1 15 9 13 1 9 2 16 15 13 9 0 2 15 1 9 13 13 2
26 9 0 0 3 13 1 9 1 15 9 16 1 15 15 13 1 9 9 2 7 1 9 0 13 13 2
19 3 3 16 9 9 3 1 15 9 9 13 3 15 0 1 9 9 13 2
21 7 13 16 15 3 12 9 13 2 15 13 0 2 16 13 1 9 9 7 9 2
12 7 1 9 9 7 9 2 7 3 13 13 2
24 13 3 16 16 9 13 2 7 0 9 13 2 1 16 15 13 2 9 9 3 13 1 9 2
28 7 1 15 2 3 15 15 13 1 9 7 9 9 3 13 2 16 15 15 13 15 9 2 0 13 7 13 2
11 3 3 16 15 15 13 9 2 3 13 2
17 7 15 1 9 9 13 1 9 2 16 13 9 7 9 13 9 2
31 13 3 2 16 15 9 13 13 15 13 1 9 7 1 9 1 9 7 9 2 16 7 1 15 15 15 13 9 1 9 2
22 15 16 3 1 15 15 13 2 7 1 9 3 2 3 13 3 9 2 7 3 9 2
13 16 13 16 9 13 13 1 13 2 1 0 0 2
34 7 15 9 9 1 9 13 0 13 4 2 3 16 3 0 1 9 7 9 13 9 2 7 3 1 15 16 9 13 1 9 1 9 2
43 1 0 13 2 16 16 9 9 13 0 1 10 9 2 3 13 16 13 13 1 9 13 0 2 7 0 3 2 3 3 1 12 9 1 9 2 7 1 12 9 1 9 2
20 3 9 13 1 9 9 10 16 9 2 1 1 9 9 13 7 1 9 9 2
19 9 1 12 8 2 13 2 16 13 9 7 9 3 13 1 15 9 0 2
6 9 7 9 9 13 2
41 7 16 0 13 1 9 1 9 15 1 15 9 2 16 9 13 2 3 3 1 15 13 15 9 13 2 2 13 16 1 9 9 13 0 7 0 16 1 9 0 2
26 1 0 3 13 2 16 9 0 13 13 1 9 16 9 2 1 16 13 9 15 9 2 7 16 9 2
12 16 0 13 16 13 9 2 3 0 9 13 2
14 16 9 15 13 9 9 13 2 13 1 9 7 9 2
21 0 7 3 13 1 9 1 16 13 9 16 9 2 7 1 16 13 15 16 9 2
15 9 7 0 13 1 15 1 9 2 16 9 13 9 9 2
10 9 3 13 4 3 16 9 15 9 2
6 7 9 13 9 9 2
9 7 9 9 0 13 1 9 10 2
18 9 15 1 9 9 13 2 1 9 9 13 2 16 1 9 0 13 2
21 3 7 0 13 16 9 1 0 9 9 13 2 16 0 9 7 9 9 9 13 2
15 3 1 9 15 3 13 16 12 9 0 9 16 15 13 2
18 7 1 2 1 12 1 9 9 13 2 16 9 9 1 9 9 13 2
23 15 3 13 9 7 9 1 9 7 9 9 2 7 1 15 12 2 15 13 9 9 15 2
15 15 15 13 9 1 15 2 1 15 15 1 9 9 13 2
9 7 15 9 9 2 9 9 13 2
28 13 7 15 9 9 3 1 15 2 7 1 9 2 1 9 9 13 2 1 16 1 9 0 13 0 9 13 2
16 7 15 13 3 13 16 15 1 9 13 2 1 9 13 9 2
8 7 15 9 13 1 9 9 2
16 16 1 15 16 9 13 15 2 13 16 9 13 15 3 13 2
13 7 15 13 1 9 1 9 2 7 3 1 0 2
29 3 9 13 1 9 0 2 3 1 9 9 9 2 15 9 9 13 2 7 1 9 9 9 2 1 15 9 13 2
12 9 3 9 13 9 2 16 13 9 1 9 2
23 9 7 12 7 9 15 2 16 9 9 7 9 9 2 13 3 15 9 2 7 13 9 2
17 7 1 15 16 9 10 13 2 13 2 7 3 16 9 2 13 2
14 1 15 7 16 9 10 0 13 9 15 9 2 13 2
16 16 13 1 9 13 2 15 9 10 13 2 9 9 13 13 2
8 7 3 15 9 9 15 13 2
14 15 7 13 1 9 16 1 16 9 7 9 15 13 2
9 9 3 13 9 10 1 9 13 2
18 7 16 9 9 3 13 9 9 2 3 13 1 9 9 9 9 9 2
26 16 3 1 0 3 13 13 12 9 0 0 9 13 15 9 9 2 3 3 13 13 12 0 9 9 2
53 3 16 9 0 1 15 16 13 12 9 2 13 9 15 9 2 3 3 9 1 15 16 15 16 0 9 13 2 15 13 15 9 3 13 2 13 1 9 0 15 13 2 1 15 13 9 0 9 2 1 9 9 2
31 9 0 2 15 13 9 13 1 12 9 2 16 13 9 9 15 2 3 13 9 9 9 15 2 16 13 1 9 7 9 2
30 9 7 1 13 9 13 0 1 10 9 9 0 2 3 13 9 9 9 2 16 1 10 9 2 16 13 1 12 8 2
58 13 7 15 9 0 16 9 0 2 9 15 13 1 9 3 2 3 9 0 15 16 13 9 0 7 1 9 2 3 15 3 13 9 0 9 2 16 13 9 2 16 9 3 13 9 1 15 2 7 1 9 2 3 9 9 15 13 2
34 16 3 9 7 9 3 13 1 9 2 16 1 12 13 4 2 8 12 2 7 1 9 2 3 3 3 13 1 9 2 7 1 9 2
35 7 1 9 15 13 16 9 2 3 13 2 16 15 9 13 1 9 7 9 2 15 3 13 1 15 0 15 0 9 13 2 16 13 4 2
7 9 0 13 15 0 9 2
25 16 3 13 15 9 7 9 15 9 0 2 13 13 0 9 16 7 13 9 9 2 13 13 9 2
19 16 13 1 9 2 15 13 9 10 1 9 13 2 1 15 13 9 9 2
19 3 7 9 9 2 1 15 9 13 2 13 3 9 15 15 9 13 13 2
28 7 16 0 9 15 15 13 2 13 9 1 9 9 2 3 3 9 1 9 9 9 13 2 13 0 1 9 2
20 1 15 3 13 15 9 15 13 1 9 2 7 15 9 2 7 1 9 9 2
7 7 13 9 1 9 9 2
19 7 15 13 7 9 2 7 9 2 7 9 2 15 1 15 1 9 13 2
23 7 16 9 9 13 1 9 9 2 7 9 13 7 9 13 2 7 1 9 13 9 13 2
36 1 0 3 13 2 16 16 9 15 9 9 13 2 13 9 1 15 9 1 9 9 9 13 2 3 3 13 9 15 1 15 1 9 9 13 2
15 7 3 1 15 9 9 13 13 2 16 9 13 9 15 2
16 3 3 15 9 13 16 9 15 2 1 16 1 9 9 13 2
15 7 9 9 1 9 3 4 13 1 9 2 16 9 13 2
10 7 3 9 9 1 9 9 15 13 2
13 1 0 13 2 16 9 9 1 9 13 0 13 2
13 7 3 3 1 9 13 2 1 15 10 9 13 2
27 7 3 9 13 13 2 3 1 15 16 1 9 13 13 2 7 16 9 13 9 1 9 2 16 9 15 2
30 3 16 1 9 9 1 9 7 1 9 2 13 15 9 0 7 0 2 3 3 9 9 9 1 9 1 15 9 13 2
38 7 3 13 16 9 9 9 3 13 2 16 15 3 0 9 1 15 13 13 16 3 1 9 13 13 2 7 3 1 16 1 0 1 9 15 9 13 2
16 3 2 9 0 15 13 9 2 13 1 9 0 15 13 9 2
17 3 2 16 9 0 13 9 1 9 2 3 0 13 9 1 9 2
8 7 9 0 3 13 12 9 2
9 3 2 9 13 9 1 9 9 2
14 3 1 0 9 13 9 1 9 2 16 13 7 13 2
16 7 9 9 13 9 2 15 13 0 2 16 0 13 9 9 2
33 16 3 3 15 9 13 13 1 15 9 2 7 15 9 1 15 9 2 7 15 0 1 15 9 2 3 7 15 9 1 15 9 2
31 13 13 2 16 15 13 13 0 15 9 15 13 15 1 9 10 9 2 1 15 1 15 9 13 2 16 9 0 13 3 2
14 9 7 1 15 9 13 9 2 13 15 9 7 9 2
10 7 9 0 1 9 13 1 9 9 2
23 13 13 2 16 9 13 9 1 9 9 2 15 13 9 9 2 16 3 9 9 3 13 2
15 9 7 9 13 9 7 9 2 15 13 15 9 7 13 2
7 9 3 0 0 9 13 2
44 3 9 7 9 3 13 9 1 16 1 9 0 13 2 7 3 1 9 15 13 9 2 16 9 15 13 1 9 0 2 7 3 1 9 0 2 16 1 12 1 9 9 13 2
21 1 0 13 9 1 15 15 13 4 2 16 9 13 9 9 1 15 9 0 13 2
25 7 3 9 7 9 9 0 7 0 1 9 0 9 13 2 16 7 15 9 13 1 0 9 9 2
44 7 1 15 9 13 13 9 2 7 13 13 9 2 16 15 9 0 13 1 10 9 2 2 16 1 15 9 3 13 13 0 9 7 1 15 2 7 13 1 9 0 7 13 2
46 13 2 16 1 12 7 9 13 2 13 16 1 15 1 15 9 13 9 2 9 1 15 9 7 9 13 2 16 13 1 0 2 16 9 15 13 9 1 9 2 13 3 9 1 9 2
9 3 13 16 0 9 13 0 9 2
37 7 16 3 9 9 9 13 9 9 2 16 1 15 15 9 3 13 2 3 3 3 13 13 9 9 2 16 13 0 9 0 2 7 3 1 15 2
25 7 16 9 3 13 9 1 9 2 7 1 9 2 3 3 0 13 9 1 15 9 15 9 13 2
11 3 1 9 9 3 13 9 1 15 13 2
12 9 7 2 7 9 2 9 1 10 0 13 2
10 7 3 15 9 9 1 9 4 13 2
15 0 3 3 13 9 16 9 3 1 10 9 13 1 9 2
28 7 16 9 1 10 9 3 1 9 13 2 15 9 9 13 2 2 3 15 13 2 3 0 2 13 13 13 2
15 13 3 0 13 1 9 7 9 2 7 1 9 7 9 2
36 15 0 13 1 3 2 7 1 15 12 1 15 9 13 2 13 16 9 7 9 2 16 9 13 9 16 9 15 2 7 9 13 1 9 0 2
49 15 9 13 9 9 9 2 16 13 13 9 1 9 7 9 2 16 15 13 1 9 2 16 13 9 1 9 2 7 15 1 9 15 2 16 16 9 13 13 9 2 3 7 9 13 13 15 9 2
50 7 13 16 13 9 0 13 1 9 0 9 7 1 9 2 16 12 9 1 9 10 13 1 9 13 0 9 2 16 9 9 2 7 9 9 2 7 9 3 13 13 16 12 15 2 7 3 1 9 2
15 12 9 16 13 9 9 2 7 3 13 9 16 13 9 2
35 15 9 13 13 9 1 9 2 16 13 9 13 9 9 2 3 3 13 13 9 2 16 13 9 1 10 9 2 1 15 13 15 10 9 2
24 15 9 13 13 9 1 9 16 13 9 9 2 16 3 13 13 9 2 7 1 9 15 13 2
26 7 13 2 16 13 9 1 9 13 7 13 9 9 2 7 3 1 15 13 15 9 15 9 1 9 2
83 1 3 15 9 13 0 2 7 1 15 13 0 9 13 1 9 7 9 9 2 7 3 15 9 9 9 0 13 2 13 16 3 13 2 9 3 13 2 13 9 9 2 16 1 9 9 9 9 13 2 7 1 9 9 9 2 7 1 9 0 9 1 9 0 9 13 2 7 0 9 15 9 0 13 2 3 9 0 15 1 15 13 2
39 16 3 2 13 2 9 1 9 7 9 9 13 2 1 10 9 13 2 9 9 9 3 13 2 7 0 9 13 2 7 0 9 9 9 9 9 9 13 2
77 3 1 9 13 9 0 2 7 1 9 2 16 13 9 15 2 7 1 9 2 16 13 9 15 2 7 13 1 15 2 0 13 16 9 15 13 9 2 7 3 1 9 9 2 16 13 9 1 9 0 2 7 1 9 0 9 2 16 13 9 13 2 13 3 9 3 1 9 9 2 3 3 1 9 9 15 2
39 1 0 13 2 16 1 9 0 13 7 13 0 1 9 7 9 9 13 2 13 12 12 9 2 16 12 0 9 13 2 16 1 12 9 0 13 12 9 2
17 7 3 1 13 2 9 9 13 12 9 2 13 9 9 7 9 2
11 13 16 3 13 9 15 1 9 9 13 2
14 9 3 15 13 15 1 15 16 1 9 0 0 13 2
8 3 1 15 9 15 3 13 2
18 3 1 9 15 13 9 1 9 2 13 16 1 0 9 15 3 13 2
17 7 13 16 7 9 7 9 13 9 15 2 1 0 1 9 0 2
8 3 1 0 9 15 3 13 2
17 7 1 2 9 15 1 9 13 13 1 13 7 9 9 1 9 2
7 3 1 0 13 9 15 2
13 3 2 9 13 9 1 3 1 9 1 9 15 2
7 3 1 0 13 9 15 2
34 13 16 10 0 9 1 0 13 2 7 9 7 9 0 2 0 7 0 2 7 0 9 15 13 1 9 9 7 9 2 15 9 13 2
16 7 15 3 9 9 9 13 2 16 15 9 0 13 9 13 2
29 7 3 9 0 3 1 15 9 15 13 2 9 13 2 7 16 13 9 15 9 2 0 3 2 7 13 9 13 2
18 15 13 3 13 2 1 0 9 13 0 9 2 7 15 9 13 9 2
10 1 0 13 2 16 9 13 1 9 2
14 9 7 0 9 13 9 0 2 1 15 9 9 13 2
35 3 3 9 0 13 9 15 13 1 9 15 13 15 9 2 16 1 15 9 2 1 15 13 1 15 9 9 3 2 16 13 1 9 0 2
19 3 3 13 13 16 9 1 15 9 13 2 16 1 15 15 13 9 15 2
37 3 1 9 15 9 9 9 13 13 2 16 13 15 13 9 2 7 3 0 2 2 13 16 9 0 2 16 3 13 9 2 13 16 9 3 0 2
31 15 7 13 15 13 1 15 16 13 9 9 3 13 16 9 2 7 3 16 9 2 16 9 13 2 1 15 9 9 13 2
29 1 0 13 2 16 1 15 16 9 13 2 13 16 15 13 9 9 1 9 9 2 16 1 15 13 12 9 0 2
8 9 7 9 9 13 3 13 2
18 7 3 1 15 16 9 0 12 13 13 2 13 9 15 13 15 9 2
23 1 0 13 2 16 2 16 1 12 1 9 13 2 15 15 15 13 0 2 13 9 15 2
27 3 1 9 0 3 13 13 9 1 9 0 2 13 16 15 15 9 13 7 13 2 13 9 0 7 0 2
31 3 3 0 0 9 13 13 2 7 9 15 0 0 2 16 9 9 13 4 16 9 15 2 3 16 1 15 12 15 13 2
24 3 7 13 2 16 1 9 9 1 9 3 13 9 15 2 1 15 1 9 1 15 9 13 2
15 7 3 9 3 13 9 16 9 2 16 9 13 9 15 2
25 1 0 13 2 16 16 9 0 3 13 13 1 9 2 3 9 3 13 9 9 2 7 1 0 2
21 16 3 1 9 7 9 15 13 0 1 9 15 1 0 13 1 9 16 9 0 2
47 7 16 9 9 1 9 13 9 13 13 0 7 0 2 15 9 13 0 1 9 9 2 3 3 1 0 9 13 15 13 2 15 13 13 16 13 1 0 9 2 16 9 7 9 7 3 2
22 0 3 1 15 16 9 9 13 1 9 2 13 15 9 1 15 9 1 9 13 13 2
19 3 2 9 2 1 13 9 2 13 0 9 2 3 9 0 1 15 13 2
40 16 9 13 1 9 2 3 16 1 15 9 1 15 9 13 2 9 0 13 2 3 3 1 15 9 1 15 9 13 2 16 9 0 13 4 2 3 13 13 2
20 1 0 13 2 16 9 13 9 0 7 13 2 3 9 9 2 7 9 9 2
20 16 1 15 9 1 15 9 13 9 2 3 1 0 9 9 2 13 9 0 2
16 1 0 13 2 16 9 16 13 0 9 2 13 3 9 9 2
13 9 7 3 13 16 9 9 13 2 7 9 3 2
9 9 7 3 13 0 9 16 9 2
32 1 15 9 2 15 1 15 9 13 2 13 13 9 13 9 9 2 3 9 7 9 2 1 15 16 1 9 0 10 9 13 2
23 9 3 15 15 13 2 13 9 9 2 15 13 9 0 1 9 13 13 1 9 1 9 2
26 3 3 1 15 2 16 9 1 12 8 13 2 9 9 13 1 9 7 9 2 7 1 15 9 15 2
31 9 7 3 13 1 9 7 1 9 1 15 2 1 3 13 0 2 7 16 9 1 15 2 1 3 13 9 16 9 15 2
18 7 13 9 7 9 15 2 16 9 13 3 2 7 13 9 1 9 2
53 1 0 0 9 9 13 4 2 15 3 9 0 9 13 16 1 0 13 3 13 2 3 3 13 9 0 9 2 7 9 2 16 9 9 1 15 16 13 9 15 10 9 1 15 13 2 3 13 1 9 1 9 2
10 9 13 9 2 9 2 7 9 9 2
40 1 9 7 0 3 13 9 0 3 2 15 9 13 0 2 7 3 0 2 2 7 13 13 9 15 9 15 1 9 13 13 2 1 9 2 7 1 9 0 2
23 3 3 13 13 16 9 15 13 1 15 9 2 13 1 15 2 7 13 9 2 7 0 2
26 9 3 15 1 15 3 13 2 3 13 2 7 0 13 2 7 9 13 9 9 2 7 13 9 9 2
15 7 3 3 13 0 16 15 9 0 1 13 13 9 0 2
21 3 13 16 9 0 13 1 9 2 0 13 1 9 1 9 0 16 13 15 13 2
16 3 3 13 1 13 13 1 9 1 15 9 1 9 9 13 2
19 7 13 13 16 13 4 1 9 9 3 2 15 3 1 9 1 9 13 2
11 13 3 9 13 0 16 13 9 1 9 2
20 7 3 9 0 1 15 13 9 2 13 9 2 15 13 9 15 7 10 9 2
27 16 7 13 9 2 9 15 13 9 2 13 7 13 15 15 13 9 2 16 9 13 9 15 15 13 9 2
21 3 7 9 9 2 15 9 9 1 15 15 13 13 2 3 13 1 9 7 9 2
24 12 9 16 7 9 13 0 7 9 0 13 1 15 9 2 16 13 1 9 9 1 9 9 2
36 1 3 10 9 13 9 13 2 16 9 0 13 1 9 15 9 1 15 9 1 15 13 9 15 9 2 3 13 9 15 9 1 9 15 9 2
11 3 3 1 15 0 9 13 13 15 9 2
35 3 2 1 10 9 0 9 0 13 9 10 1 9 15 0 15 9 13 3 13 2 16 9 1 9 9 2 15 0 9 9 13 3 13 2
16 1 0 13 2 16 9 7 9 2 3 13 1 9 16 9 2
31 16 16 9 13 1 9 9 2 9 13 3 13 1 9 13 2 1 15 13 1 9 2 16 1 9 1 15 0 13 4 2
18 15 3 15 9 13 2 13 9 15 9 2 16 9 0 9 13 13 2
42 7 16 1 9 13 9 0 13 13 9 9 9 2 3 3 13 1 9 0 9 1 15 9 13 16 1 9 2 1 16 13 1 9 9 2 16 13 1 0 9 9 2
16 7 3 15 9 3 13 1 12 9 0 13 2 15 13 0 2
28 1 0 7 9 9 15 9 13 2 3 9 7 9 0 9 13 2 7 9 2 7 1 9 0 9 13 4 2
14 3 9 9 7 9 9 0 0 13 15 1 15 9 2
13 16 2 16 13 9 2 15 9 9 0 9 13 2
25 7 1 2 10 9 0 13 1 15 1 9 15 9 2 16 7 9 9 13 1 15 1 10 9 2
12 9 7 13 15 9 1 9 2 7 1 9 2
20 7 3 9 13 2 16 1 9 9 13 9 2 7 9 9 1 15 13 9 2
41 7 16 3 0 9 13 1 9 2 7 1 9 13 2 3 13 4 1 13 15 9 2 1 15 13 9 1 12 8 2 7 1 13 3 15 9 2 16 13 9 2
21 9 7 2 1 9 15 9 7 9 13 9 2 13 12 9 2 1 9 12 8 2
15 7 15 13 9 9 2 15 16 9 2 15 7 16 9 2
14 3 2 3 13 0 9 9 1 9 16 9 1 9 2
16 7 1 9 9 13 9 9 2 16 0 9 13 1 0 9 2
11 1 0 13 2 16 9 13 9 13 15 2
12 7 3 13 16 1 0 9 0 13 9 13 2
19 3 2 9 2 16 13 9 2 13 15 9 9 2 16 9 13 9 9 2
14 7 3 13 1 9 9 16 9 2 15 13 9 9 2
25 16 3 9 0 1 15 9 3 13 13 9 15 9 2 0 0 9 0 13 13 9 15 15 9 2
37 1 9 7 15 3 3 13 16 15 0 13 2 16 13 1 13 9 7 9 2 15 15 3 13 9 0 2 7 1 9 2 16 15 13 9 13 2
59 1 3 0 9 7 0 15 13 2 3 15 13 0 1 9 2 7 0 9 9 13 0 1 15 13 1 9 2 7 1 15 0 13 2 1 15 13 1 15 15 13 2 13 2 16 13 13 9 2 16 0 9 13 1 0 9 9 0 2
21 1 0 13 2 16 9 0 3 13 0 9 16 1 15 13 2 16 9 1 9 2
7 9 9 13 2 3 9 2
29 1 0 3 13 2 16 16 9 13 15 9 15 9 13 1 9 13 2 3 3 9 2 7 10 15 13 0 9 2
8 7 1 2 15 9 13 9 2
5 7 9 13 9 2
17 15 13 9 9 15 10 0 13 2 16 9 13 9 16 9 9 2
29 1 2 13 2 1 0 13 2 16 1 9 9 13 2 13 13 0 7 13 2 1 15 9 9 0 9 13 13 2
30 13 2 16 9 0 13 9 2 3 16 13 9 15 9 2 7 16 3 13 9 15 9 2 7 15 9 1 15 13 2
31 9 0 0 13 9 2 3 16 13 9 3 0 2 13 3 7 9 7 9 2 2 7 1 9 15 9 9 13 9 15 2
18 0 3 13 3 3 9 2 7 3 9 9 2 3 13 13 9 15 2
12 16 7 9 9 2 13 1 9 2 7 9 2
6 9 7 3 13 9 2
27 7 16 15 13 9 2 13 2 16 15 9 1 9 7 9 2 15 13 9 9 2 3 13 15 0 0 2
17 7 9 2 0 13 2 13 13 9 7 9 2 1 15 13 9 2
26 3 3 13 13 2 16 13 1 12 9 3 13 9 15 9 13 2 7 9 1 15 13 2 3 9 2
14 9 15 7 2 7 9 12 3 13 15 9 7 9 2
7 10 3 9 0 13 9 2
6 7 9 13 9 0 2
23 9 3 0 2 13 15 13 9 16 15 15 13 2 16 13 9 7 9 16 15 15 13 2
23 1 0 3 13 2 16 9 13 9 2 3 3 16 15 9 13 9 7 9 2 7 0 2
22 16 3 9 1 9 7 9 13 1 15 0 2 13 1 9 15 9 9 0 1 15 2
64 16 7 3 13 1 15 0 2 3 13 1 9 9 15 9 2 7 0 15 15 13 2 13 9 1 9 1 15 15 15 13 2 16 16 13 9 13 1 9 2 7 9 1 15 13 13 2 7 3 15 0 13 2 13 16 9 9 13 9 9 1 15 0 2
21 7 16 13 9 2 3 13 1 9 9 15 9 9 2 16 9 3 13 9 0 2
14 3 2 9 3 13 13 2 16 9 13 15 3 9 2
16 16 3 9 3 4 13 9 0 3 9 2 13 9 15 0 2
12 16 9 13 1 9 13 2 7 3 13 13 2
13 7 9 13 3 1 9 13 2 3 3 1 9 2
15 3 2 9 13 13 1 9 13 2 16 9 13 13 0 2
18 7 9 13 1 15 9 9 7 1 15 9 9 2 13 0 0 9 2
34 9 3 13 9 0 2 15 3 3 13 1 9 13 1 15 9 9 2 7 13 1 15 9 0 9 2 15 13 15 1 9 0 9 2
40 16 1 15 2 9 13 9 2 9 13 13 9 9 9 2 7 9 9 13 1 9 2 7 1 15 2 9 13 9 2 9 3 13 9 9 9 13 1 9 2
22 16 9 3 13 9 9 13 1 9 2 7 9 9 2 16 13 1 1 8 1 0 2
29 1 0 13 2 16 1 13 2 9 13 9 2 9 9 3 1 9 13 13 0 2 7 3 1 9 13 9 13 2
32 3 3 13 16 13 13 1 10 15 13 9 13 1 15 9 9 2 16 3 13 1 15 1 9 9 13 2 7 1 9 9 2
34 7 3 15 3 13 1 9 2 9 13 9 2 7 13 15 0 1 15 15 13 1 9 2 16 9 3 13 9 9 9 13 1 9 2
16 7 9 9 9 1 0 13 8 12 2 12 2 9 9 13 2
49 1 0 13 2 16 9 3 13 0 2 7 9 9 2 13 9 2 7 16 9 9 13 2 16 0 9 0 16 13 2 16 13 9 2 0 9 2 1 9 9 2 7 9 13 2 7 13 13 2
9 9 7 7 9 13 13 1 13 2
17 13 3 9 9 2 1 15 13 15 1 9 2 16 9 7 9 2
43 7 3 2 1 3 13 7 1 9 7 1 9 2 3 13 1 15 13 2 16 9 9 13 0 2 16 13 9 2 15 13 13 1 9 2 1 9 15 13 9 1 9 2
20 7 15 13 9 2 15 1 9 0 13 2 13 9 0 2 13 15 13 0 2
19 7 9 2 15 13 9 9 2 13 0 15 15 9 1 15 13 15 9 2
63 1 0 13 2 16 16 9 13 1 12 1 8 2 10 15 9 7 9 1 9 9 13 13 2 7 13 13 1 9 13 1 15 0 13 9 2 1 9 9 13 0 9 2 16 13 1 8 12 2 7 13 13 1 9 9 2 1 16 9 13 9 9 2
16 7 1 9 9 9 13 0 9 9 2 16 9 9 1 15 2
34 15 0 13 13 2 16 9 1 15 13 2 7 0 2 16 9 7 9 2 7 3 9 15 13 13 2 7 0 2 16 9 13 13 2
7 3 3 13 9 16 9 2
41 7 3 15 15 13 1 9 9 2 15 9 13 1 9 7 1 0 7 1 9 2 7 1 0 7 1 0 2 16 9 3 13 0 12 2 7 9 13 9 15 2
19 7 1 15 16 9 13 1 15 2 13 16 13 15 9 9 13 1 9 2
7 7 9 9 9 9 13 2
17 7 13 16 13 15 9 9 13 7 13 2 16 13 9 1 15 2
32 1 0 13 2 16 15 9 1 0 13 1 9 9 2 16 7 9 9 13 1 9 9 15 9 9 13 2 16 13 1 9 2
13 3 13 15 9 13 1 15 13 2 15 0 13 2
34 1 0 13 2 16 16 10 9 13 1 15 13 1 13 2 16 7 13 0 2 13 15 1 9 2 2 3 3 13 1 9 9 9 2
27 16 7 13 15 9 0 0 15 3 13 10 9 2 13 3 9 3 1 9 2 15 13 13 1 9 15 2
22 7 15 9 3 13 13 2 16 3 4 1 15 13 2 16 16 13 9 1 15 13 2
10 7 1 15 3 9 0 13 13 9 2
47 7 16 9 15 4 13 1 15 2 1 9 13 13 3 1 9 13 15 9 2 3 0 3 1 9 0 2 16 3 0 3 13 9 13 0 2 7 15 9 2 15 9 15 13 0 13 2
35 7 0 13 16 3 13 13 3 1 9 15 9 2 16 3 13 15 9 1 10 9 9 15 2 16 15 15 13 1 13 1 9 15 9 2
9 13 7 9 15 9 15 13 0 2
83 1 0 3 13 2 16 16 1 9 0 9 13 1 10 9 2 13 9 1 9 2 7 13 1 9 12 1 9 2 7 1 15 13 9 12 0 9 2 3 3 10 9 9 0 13 1 0 9 9 0 2 15 13 12 9 1 10 2 7 15 9 13 1 15 1 9 0 2 16 13 1 0 1 9 2 13 3 1 12 9 1 9 2
37 3 2 1 9 7 9 3 13 15 9 0 2 16 7 1 9 7 9 2 16 1 9 0 7 9 13 9 0 2 15 3 13 0 15 9 0 2
54 15 9 13 15 1 9 2 16 13 9 1 9 9 2 3 16 13 1 9 1 9 9 13 2 3 9 13 2 16 9 13 1 9 9 2 3 16 0 13 1 9 7 9 2 7 9 13 1 9 9 1 9 9 2
47 1 0 13 2 16 15 13 15 13 0 15 1 15 2 15 13 0 0 2 16 3 9 9 0 1 15 13 0 15 9 2 16 15 13 1 15 16 9 1 9 2 1 13 9 0 15 2
35 1 0 9 13 2 16 15 9 0 13 1 9 13 16 13 1 9 0 2 1 15 13 1 9 2 16 15 13 16 1 16 13 1 9 2
18 15 9 1 9 9 7 9 2 16 9 0 3 13 4 0 15 0 2
30 1 9 7 13 1 15 9 16 9 10 0 13 1 15 3 0 1 9 9 2 7 3 1 9 9 7 9 0 9 2
6 7 15 9 9 13 2
37 16 3 9 0 9 13 1 13 2 13 16 1 0 9 13 15 13 2 16 3 9 0 3 0 13 1 15 1 9 9 2 7 3 1 9 9 2
14 3 13 1 9 1 9 2 16 10 9 13 0 9 2
32 1 15 7 16 15 13 15 0 2 13 16 13 1 9 15 0 9 1 15 13 13 9 2 16 1 9 2 9 0 15 13 2
27 7 1 15 16 15 13 0 0 2 13 16 9 10 15 0 9 13 2 16 16 1 9 13 0 9 9 2
29 7 3 13 16 15 15 13 1 9 12 7 0 2 9 0 9 7 9 13 2 15 15 13 1 9 9 0 9 2
18 9 7 13 13 9 9 16 4 13 2 16 1 15 13 9 1 9 2
20 3 16 1 9 7 9 13 12 9 2 3 9 13 7 9 13 13 12 13 2
49 1 0 13 2 16 9 13 9 15 13 1 9 2 3 1 15 9 15 9 13 1 9 2 7 1 15 16 9 15 13 16 9 9 13 2 16 13 1 15 2 7 15 9 13 9 10 15 9 2
20 10 7 15 13 1 9 1 9 15 2 13 0 2 16 15 9 13 1 15 2
25 3 1 9 0 3 13 0 2 13 16 9 9 1 15 9 0 13 1 9 2 4 13 1 15 2
19 7 1 15 16 13 9 13 16 15 9 9 13 9 16 9 15 13 13 2
49 1 0 13 2 16 12 9 3 13 1 15 1 15 15 13 13 1 9 2 7 1 15 15 3 13 2 15 0 13 7 1 9 2 7 1 9 15 9 3 15 13 2 1 15 13 9 3 0 2
18 7 9 0 2 1 13 9 0 9 0 2 13 3 0 9 16 0 2
68 1 0 3 13 2 16 1 15 9 3 13 16 16 13 10 15 1 9 0 13 13 2 16 16 9 0 13 1 0 9 3 1 15 9 15 1 9 0 13 13 2 16 9 15 1 9 15 13 13 2 3 3 9 0 13 1 9 0 15 3 15 1 9 9 13 13 13 2
23 16 3 15 13 9 15 16 9 13 16 9 2 3 15 9 9 13 2 13 3 9 9 2
18 3 9 13 1 9 9 3 1 15 3 16 9 2 16 13 9 9 2
21 9 7 9 1 0 9 13 13 1 15 1 15 16 9 0 1 15 13 0 0 2
11 16 3 9 13 13 2 3 9 13 13 2
25 13 7 9 7 1 9 10 2 1 16 13 9 0 2 7 1 9 10 9 2 16 13 9 15 2
20 1 7 16 13 9 16 9 2 3 3 13 16 15 0 2 7 16 13 15 2
19 3 3 3 13 1 15 2 7 1 9 2 16 15 9 13 13 9 13 2
40 7 16 3 9 3 13 0 2 7 9 9 0 2 3 3 13 13 1 15 2 7 9 1 15 2 7 1 9 2 16 9 13 2 16 13 1 12 1 9 2
56 7 16 9 3 13 1 0 1 9 13 2 1 9 0 3 13 1 9 1 9 0 16 13 1 0 2 7 1 9 0 2 15 13 0 9 2 3 3 13 9 1 9 2 7 13 9 15 2 16 1 16 13 9 9 2 2
29 1 0 13 2 16 16 1 9 9 2 9 3 13 0 3 1 9 2 13 3 9 2 1 15 9 13 9 9 2
23 13 7 9 0 2 3 1 9 2 16 13 9 7 1 9 2 3 3 10 2 7 15 2
47 13 3 1 9 0 13 2 3 3 1 9 2 15 13 0 1 15 2 15 13 1 0 1 10 9 9 2 1 16 1 9 9 13 2 1 15 3 9 9 13 2 1 16 13 15 9 2
65 7 3 2 1 9 1 10 9 13 9 9 2 7 9 7 10 15 9 13 9 9 2 7 1 9 1 9 9 13 0 2 3 1 9 9 1 9 2 7 1 9 9 1 15 9 15 13 1 9 0 2 1 15 9 13 9 1 9 9 2 16 1 0 13 2
10 3 3 0 9 10 9 13 1 9 2
10 3 2 9 13 13 1 9 13 9 2
12 7 9 9 0 2 9 3 0 2 13 0 2
65 7 3 1 9 9 9 15 1 9 3 13 9 13 2 16 15 1 9 15 9 2 1 9 10 9 0 9 13 2 16 15 0 13 2 7 3 1 9 9 0 2 16 15 13 9 13 2 7 9 15 3 13 2 7 15 9 1 9 13 13 15 9 9 13 2
28 1 0 13 2 16 9 13 13 13 9 2 3 16 13 9 9 2 7 16 13 13 1 13 9 1 9 10 2
32 1 0 13 2 16 3 13 13 16 9 13 1 9 1 9 9 2 16 9 0 3 13 0 1 15 9 2 16 13 9 9 2
29 15 7 3 13 1 0 9 2 15 13 9 0 2 7 1 9 2 15 13 9 13 7 0 15 9 0 3 13 2
28 1 0 13 2 16 9 13 3 1 15 15 9 13 2 16 13 9 0 1 9 2 1 15 9 13 4 13 2
21 9 7 9 13 9 2 16 13 1 12 8 2 16 15 13 9 15 9 15 13 2
32 7 3 16 13 0 9 2 13 3 0 9 2 16 9 13 7 13 1 9 7 9 2 7 9 13 7 13 1 9 7 9 2
30 1 0 13 2 16 16 13 13 9 2 3 9 7 9 13 9 7 9 13 1 9 2 16 7 15 9 1 9 13 2
28 3 16 15 9 13 9 0 9 1 0 15 9 13 15 9 2 3 15 9 13 0 9 1 0 9 7 9 2
17 7 1 0 9 1 9 13 2 3 1 9 9 2 7 1 9 2
42 7 15 7 1 9 1 9 9 2 16 1 2 8 12 2 8 12 2 8 12 2 13 4 2 16 9 9 1 9 13 3 2 16 13 9 15 2 7 1 9 0 2
59 16 7 9 1 10 9 13 9 9 2 9 7 13 16 13 9 13 2 3 1 15 9 9 3 1 9 13 2 13 16 4 13 13 1 9 9 2 16 3 13 9 1 9 3 1 15 9 15 0 15 13 13 7 1 9 7 1 9 2
18 1 0 13 2 16 9 9 13 1 9 9 2 16 9 7 9 9 2
11 1 15 9 13 4 2 1 15 13 4 2
18 13 3 9 0 2 12 9 13 9 2 7 15 13 0 9 13 9 2
10 15 9 13 0 13 9 1 13 9 2
12 0 3 13 13 9 2 16 13 9 1 9 2
22 7 0 13 9 0 1 9 0 9 2 16 13 15 2 9 9 13 2 16 9 9 2
26 3 2 16 15 9 3 13 13 1 0 1 0 9 2 3 12 9 1 0 3 13 13 0 7 0 2
12 3 3 13 13 2 16 9 9 13 9 9 2
12 1 0 13 2 16 9 3 13 13 9 9 2
61 1 0 13 2 16 16 15 15 13 1 9 0 1 9 9 3 13 13 1 9 9 2 16 15 13 13 0 0 7 15 9 2 3 3 15 15 13 1 9 0 16 13 9 9 2 3 13 13 1 9 9 2 16 16 13 9 2 7 15 3 2
33 3 2 9 3 13 1 9 16 1 9 13 9 9 2 15 13 16 9 1 9 13 2 16 1 15 9 9 13 0 1 15 9 2
35 1 0 13 2 16 16 15 9 9 2 15 13 9 1 9 9 2 4 13 1 9 2 3 3 3 13 4 9 7 9 9 2 9 13 2
10 3 2 10 9 13 1 9 15 13 2
8 7 9 9 0 13 9 0 2
11 16 3 13 15 2 1 9 0 15 13 2
30 7 3 13 2 16 1 9 9 0 13 16 13 7 3 13 2 7 3 16 13 2 16 13 1 9 9 2 7 3 2
46 1 3 13 1 15 9 0 9 2 7 9 9 2 13 1 12 3 13 9 2 7 1 15 2 7 13 9 1 9 9 1 9 9 2 16 3 13 2 7 13 2 16 1 0 13 2
25 1 0 13 2 16 9 0 9 0 10 9 13 2 15 13 3 9 13 2 7 3 9 9 9 2
17 13 3 1 9 9 16 13 2 16 13 1 9 0 16 13 13 2
9 7 9 7 9 13 1 9 15 2
8 9 7 15 13 1 9 9 2
13 7 3 9 3 13 9 9 2 7 13 9 0 2
33 13 3 0 13 1 0 9 16 15 13 9 9 13 2 8 12 2 7 16 1 0 9 13 1 9 2 1 15 3 1 3 13 2
26 16 13 15 1 9 1 15 13 0 9 2 3 3 1 0 13 15 0 9 2 16 13 9 1 9 2
22 9 7 13 0 2 3 1 9 15 13 9 0 9 2 7 1 9 15 13 9 0 2
21 13 3 16 15 9 13 2 3 1 9 9 13 2 16 9 9 13 9 9 13 2
18 3 3 0 7 0 15 0 13 2 13 16 15 15 13 13 10 9 2
16 7 15 3 9 2 7 9 2 16 3 13 0 2 9 13 2
32 9 7 2 16 13 1 12 1 9 2 16 15 2 13 15 2 16 3 1 9 3 3 15 2 7 9 2 15 13 9 15 2
22 16 3 9 1 0 9 9 13 2 15 9 0 13 0 15 9 13 0 1 9 9 2
51 13 13 2 16 13 9 9 13 0 7 0 9 9 3 1 15 15 13 1 9 2 7 3 3 1 9 9 2 15 9 2 7 3 9 2 13 2 16 3 7 9 9 13 13 15 1 15 9 13 13 2
14 7 3 13 1 9 0 2 16 9 13 1 9 9 2
13 13 3 15 1 9 0 2 3 16 13 9 0 2
17 1 0 3 13 2 16 9 3 13 3 1 9 2 7 1 9 2
16 9 7 9 3 13 9 2 16 1 13 2 15 1 9 13 2
10 9 3 13 13 2 1 13 9 9 2
10 3 2 10 9 13 9 1 0 9 2
7 3 9 3 13 9 9 2
9 3 2 12 9 3 13 0 9 2
8 3 2 9 9 13 9 15 2
9 3 2 9 9 13 1 9 10 2
6 7 9 9 13 9 2
12 3 2 15 9 1 9 13 15 9 1 9 2
20 0 9 15 15 1 16 10 13 7 13 13 10 9 1 13 7 13 1 15 2
33 15 7 9 7 13 1 9 15 9 2 1 16 10 9 13 1 9 9 1 15 13 2 7 13 1 9 13 9 2 15 13 9 2
17 7 3 10 9 15 13 1 9 13 1 9 9 2 13 9 9 2
14 15 3 9 15 1 9 9 13 13 2 13 10 0 2
28 3 1 15 9 2 15 13 9 15 2 13 0 9 2 1 16 13 9 15 13 2 1 9 1 9 7 9 2
17 3 1 9 2 15 13 9 9 2 13 9 0 15 7 15 9 2
17 3 1 15 13 9 0 1 9 0 9 2 7 9 1 15 13 2
11 7 3 1 15 3 9 13 1 9 9 2
21 1 0 13 2 16 1 9 15 13 9 1 9 9 7 9 0 2 13 9 9 2
14 7 9 9 13 1 9 15 13 1 9 13 7 13 2
25 3 1 12 9 12 9 3 13 3 13 1 15 9 2 13 16 13 9 7 9 2 9 0 13 2
9 3 7 9 0 13 1 9 9 2
21 12 7 9 12 9 3 13 3 13 2 16 9 13 1 9 1 9 9 7 9 2
15 3 2 9 0 3 13 9 13 2 16 13 1 9 13 2
21 3 9 0 2 15 13 9 0 2 3 13 2 16 13 1 9 1 12 1 9 2
15 7 9 0 13 3 1 9 7 9 13 16 15 9 0 2
40 7 16 15 13 1 16 13 1 9 7 1 10 9 2 9 7 13 0 1 9 0 2 3 9 9 2 1 15 13 9 0 2 13 15 15 13 0 1 9 2
24 1 0 13 2 16 9 0 3 13 1 16 1 10 9 13 2 7 1 16 13 1 15 0 2
13 7 13 2 16 9 0 3 13 0 1 9 9 2
23 3 13 9 9 1 9 2 0 13 2 13 16 1 9 0 15 9 0 13 1 9 10 2
43 7 1 15 13 16 9 3 13 13 1 13 2 16 9 15 0 15 0 13 9 9 2 3 9 2 9 9 10 13 2 7 3 13 15 0 1 9 9 2 16 13 9 2
22 3 0 1 15 9 9 9 13 15 9 15 15 13 2 7 9 1 15 15 3 13 2
18 16 3 9 13 9 13 1 9 2 15 13 1 9 0 9 1 15 2
12 3 2 0 13 1 13 1 9 1 0 9 2
12 10 7 0 13 1 16 13 1 9 10 0 2
13 16 9 2 16 13 1 9 0 2 13 7 13 2
27 0 16 9 7 9 3 13 9 9 15 13 15 9 2 13 15 1 15 2 7 13 15 16 13 1 15 2
28 7 16 10 15 13 9 15 2 13 12 1 15 2 3 1 9 13 13 12 1 13 2 15 4 13 9 13 2
16 15 7 13 1 9 10 9 2 15 13 9 13 7 9 9 2
13 7 15 9 13 0 15 0 2 3 9 10 13 2
28 7 16 9 3 13 13 1 9 15 13 15 1 9 10 9 2 16 1 9 2 3 7 13 16 13 1 9 2
16 1 0 13 2 16 9 13 13 13 2 16 13 13 10 9 2
44 16 3 13 1 15 16 9 13 2 15 3 9 13 2 16 0 3 13 4 9 13 2 2 3 15 15 13 2 3 3 13 2 16 13 1 9 2 15 9 0 13 0 9 2
40 1 15 3 16 9 13 13 1 13 2 13 13 13 1 0 13 2 7 1 1 2 16 15 13 13 13 3 13 2 16 9 13 1 0 13 2 7 1 0 2
39 7 16 15 13 1 15 13 16 1 1 1 10 9 3 13 2 16 12 12 13 9 2 3 15 9 9 13 15 9 2 15 13 1 15 13 1 13 13 2
46 16 0 15 1 15 13 16 13 15 15 1 15 13 2 16 9 0 3 13 9 16 13 9 15 9 1 9 13 2 3 13 16 1 13 9 15 2 15 1 9 10 3 13 2 13 2
17 15 13 13 15 13 12 0 2 16 13 0 2 7 9 7 9 2
14 7 15 13 13 9 2 16 9 13 13 13 9 13 2
27 1 0 13 2 16 15 9 0 1 13 9 2 15 13 15 1 0 9 2 9 15 13 2 16 1 13 2
26 7 15 9 1 9 0 13 7 13 13 2 16 7 9 12 13 13 2 1 15 1 12 3 9 13 2
9 13 16 9 3 13 9 15 9 2
9 10 3 9 7 13 0 7 0 2
31 7 9 3 13 9 0 9 2 16 3 1 15 9 13 15 9 2 7 3 13 9 0 2 16 13 9 7 9 15 9 2
8 3 9 15 9 13 9 9 2
13 7 9 13 13 9 10 9 2 16 13 9 0 2
6 3 9 3 13 9 2
25 7 3 9 13 3 9 9 16 9 2 7 3 9 2 15 3 13 1 9 3 9 10 15 9 2
18 3 2 9 0 7 9 3 13 1 15 9 2 16 13 1 12 8 2
6 3 15 3 13 9 2
22 7 15 9 13 10 9 7 9 1 9 10 2 1 15 0 0 13 2 7 0 0 2
35 3 2 15 15 13 0 2 3 1 0 2 13 0 9 15 2 16 9 13 3 9 9 2 9 9 2 7 9 9 2 16 13 12 8 2
7 3 15 13 9 15 9 2
8 3 2 9 3 13 13 0 2
8 7 9 13 9 10 15 9 2
22 1 0 9 13 2 16 9 1 10 15 9 13 7 16 9 7 16 9 7 16 9 2
13 0 3 13 16 13 9 13 15 9 1 9 9 2
14 7 1 15 9 13 9 7 9 1 10 15 9 0 2
13 7 3 9 13 9 9 15 10 2 16 9 0 2
12 7 15 13 12 9 15 9 13 9 15 9 2
12 1 0 3 13 2 16 9 13 9 0 9 2
6 7 9 0 13 0 2
18 7 1 15 3 13 16 9 3 2 16 13 9 0 13 9 0 9 2
33 15 9 13 9 0 1 15 9 15 13 2 7 1 15 9 9 13 2 16 0 9 13 9 0 10 9 2 7 0 9 10 9 2
22 7 15 9 0 3 13 16 13 12 9 1 13 2 16 13 3 3 13 1 9 13 2
26 7 15 9 9 13 9 15 9 0 2 16 9 15 9 1 9 9 13 9 15 3 13 2 9 9 2
18 3 1 9 9 1 15 9 15 9 13 2 15 0 13 9 15 9 2
18 7 3 9 2 15 13 9 9 2 13 9 9 2 15 13 9 0 2
9 7 3 9 13 9 9 7 9 2
25 7 3 9 2 15 13 9 9 9 2 13 15 1 9 0 2 13 9 7 9 7 9 7 9 2
26 1 0 13 2 16 9 0 13 1 15 9 1 13 7 9 2 16 13 1 9 2 3 7 9 0 2
24 7 3 15 9 15 13 1 9 9 2 13 3 9 2 15 13 9 2 1 9 9 0 9 2
18 7 9 15 13 15 9 2 13 1 9 0 9 1 9 1 0 9 2
23 7 15 9 7 9 13 15 9 1 10 9 2 7 3 15 9 7 9 15 13 1 0 2
15 0 9 13 13 1 15 16 15 9 13 10 9 7 9 2
25 7 0 1 15 15 13 9 2 13 1 9 16 1 9 2 16 9 13 9 2 7 9 13 9 2
32 7 16 15 13 0 9 1 15 9 13 13 2 3 15 13 0 1 15 9 3 13 13 2 16 13 1 0 1 12 9 0 2
19 7 1 2 9 16 13 2 16 1 15 0 13 2 3 0 1 15 13 2
12 7 9 7 9 1 13 9 2 9 15 13 2
31 13 7 0 9 2 3 9 15 13 9 0 16 3 2 16 9 2 7 9 15 13 9 9 16 3 2 16 9 13 9 2
58 16 7 9 9 15 13 0 0 2 3 13 1 9 7 9 2 3 15 13 3 13 15 9 15 9 2 7 15 9 2 16 13 16 16 1 0 13 0 2 7 1 0 2 13 15 15 9 13 2 3 15 9 9 2 7 15 9 2
20 3 15 13 9 15 0 1 10 0 2 16 15 13 9 0 1 10 9 0 2
9 15 9 1 15 16 13 9 9 2
17 7 9 0 13 9 10 1 9 2 16 13 1 9 13 1 0 2
13 3 2 0 9 12 9 3 13 13 1 15 9 2
31 9 7 9 2 15 13 1 9 16 1 0 9 2 13 16 1 9 0 13 2 16 3 9 9 13 1 9 1 0 9 2
13 9 7 13 1 9 15 13 1 9 9 7 9 2
29 7 3 15 9 9 9 9 7 9 13 2 16 3 13 1 0 2 16 0 9 3 13 13 1 13 9 12 9 2
13 3 2 12 9 15 9 3 13 13 1 12 9 2
46 13 13 1 0 9 2 16 16 1 0 13 15 9 10 13 1 9 2 7 16 9 0 13 15 1 0 1 0 2 16 13 15 15 13 9 15 13 2 3 3 13 15 1 9 9 2
37 0 3 13 2 16 13 15 9 13 1 9 2 16 9 13 1 9 9 2 7 9 9 1 9 0 2 16 15 1 0 13 2 0 1 0 13 2
21 13 7 13 13 9 2 16 9 9 2 1 16 13 1 9 2 13 1 9 0 2
33 1 0 9 13 13 2 16 15 9 2 15 13 9 2 13 10 9 13 1 9 2 7 16 9 0 3 13 16 9 1 9 15 2
18 7 1 9 15 13 9 2 13 0 15 15 13 9 16 15 13 9 2
12 3 2 15 13 9 9 1 15 13 9 15 2
7 7 9 13 9 13 0 2
13 9 3 0 2 16 13 9 2 9 13 3 13 2
7 7 9 9 13 9 0 2
23 1 0 3 13 2 16 9 15 7 13 9 1 15 7 1 15 2 15 9 13 13 9 2
33 9 7 15 13 9 1 15 2 16 3 13 9 1 15 2 13 13 9 3 16 0 13 9 2 7 16 15 15 13 9 9 13 2
44 7 16 9 13 0 0 2 15 1 9 3 13 2 7 3 3 0 9 13 2 3 9 13 0 3 0 0 2 15 13 0 1 0 13 1 13 2 7 3 0 15 3 13 2
44 15 0 15 1 15 13 9 2 3 0 2 7 0 2 13 1 15 2 16 16 9 9 0 2 1 15 0 13 2 13 1 15 16 1 9 9 2 7 3 13 3 9 9 2
19 3 1 15 9 13 3 15 9 9 2 1 16 0 9 13 16 0 9 2
31 3 13 9 7 9 2 16 13 9 9 1 15 1 15 9 9 15 13 2 7 9 2 15 2 13 9 9 9 15 13 2
57 7 1 15 13 9 15 13 1 9 0 1 15 16 13 9 9 1 15 1 15 9 9 15 3 13 2 7 0 0 2 7 0 0 2 1 15 13 9 2 7 3 3 2 7 3 0 2 7 9 2 15 13 9 0 9 0 2
22 3 7 9 3 9 13 2 3 9 13 2 16 9 3 3 13 9 2 3 9 13 2
57 7 3 3 1 9 9 13 9 9 3 0 1 9 9 2 15 9 9 9 3 13 2 7 13 1 9 0 9 2 2 7 3 1 9 2 7 9 2 7 0 9 1 15 10 13 13 9 1 8 1 0 9 13 1 0 9 2
80 1 0 9 13 2 16 1 10 9 0 13 16 9 1 10 9 9 13 15 1 15 13 2 15 3 13 1 15 9 2 16 9 1 9 13 2 16 13 1 9 7 9 9 2 16 16 9 0 13 1 9 9 2 9 9 13 2 7 9 3 1 9 9 13 2 16 0 13 9 2 3 13 9 9 2 16 1 15 9 2
16 0 15 13 15 9 2 13 16 9 13 2 15 13 9 9 2
16 0 1 9 2 15 13 9 9 2 1 15 10 9 3 13 2
25 7 13 2 16 15 3 13 9 2 16 16 1 0 9 7 9 13 1 15 2 3 7 1 0 2
13 7 13 3 3 13 9 9 3 4 13 1 9 2
31 15 15 3 7 3 13 0 2 16 15 1 15 13 9 9 7 9 1 0 2 16 0 13 2 9 13 2 7 15 3 2
21 12 9 3 1 9 15 13 13 1 9 2 7 3 13 1 15 2 3 9 9 2
13 7 3 13 9 0 2 15 1 15 9 9 13 2
6 0 13 1 9 9 2
6 0 13 9 13 9 2
14 0 13 2 3 13 13 9 15 13 0 9 2 3 2
11 0 13 9 9 15 13 1 9 2 3 2
5 0 13 9 9 2
7 0 13 9 9 1 0 2
7 7 15 13 0 9 13 2
31 3 2 0 15 13 1 9 16 15 12 2 16 13 9 13 2 13 9 13 2 16 3 9 1 9 13 2 7 0 3 2
29 1 0 13 2 16 1 9 2 15 13 9 13 2 13 13 9 7 9 7 9 7 10 15 1 9 13 13 13 2
20 7 9 13 3 9 3 2 7 3 1 0 9 13 2 16 15 13 1 9 2
44 3 16 13 9 4 2 16 9 3 13 1 9 2 3 7 16 15 9 13 0 13 9 13 2 3 3 9 2 15 9 9 13 2 13 9 15 13 1 9 15 9 13 13 2
34 1 0 13 2 16 15 15 13 1 9 2 13 3 3 1 9 9 2 7 3 3 1 9 0 2 7 9 15 15 13 1 9 0 2
20 15 3 13 2 16 1 0 9 2 16 0 9 13 2 15 9 1 13 13 2
26 7 3 9 0 15 9 13 3 9 13 2 7 3 9 13 2 16 1 9 9 15 2 9 9 13 2
25 9 3 0 13 2 15 3 9 13 9 9 2 7 0 9 9 2 16 15 9 13 7 9 13 2
15 9 13 0 9 0 9 2 16 9 13 2 7 9 13 2
9 3 13 13 2 0 7 0 9 2
9 3 2 10 9 13 0 7 0 2
31 7 9 3 13 9 0 0 9 2 16 1 15 13 2 7 3 9 0 2 1 9 0 3 13 9 0 2 7 1 0 2
9 3 9 15 9 13 9 0 9 2
7 7 15 15 13 9 0 2
10 9 7 0 13 1 15 9 15 13 2
10 3 3 13 15 9 7 9 9 15 2
7 7 9 13 9 0 9 2
51 13 3 9 9 1 15 16 13 2 16 9 13 2 7 9 13 9 3 1 9 2 1 15 16 13 2 0 9 0 9 2 7 9 9 9 0 2 3 1 9 0 2 1 15 16 13 2 16 9 13 2
34 1 0 13 2 16 9 13 3 0 1 9 2 1 16 13 1 0 9 9 2 7 3 1 9 0 2 16 1 9 9 9 15 13 2
17 7 16 13 1 9 0 2 15 13 16 9 13 3 9 0 9 2
25 1 0 13 2 16 1 0 2 16 9 15 13 9 2 3 13 9 1 9 2 1 9 9 13 2
21 15 3 13 9 0 9 0 9 13 2 7 1 9 13 2 16 0 9 0 9 2
69 1 0 3 13 2 16 16 9 0 13 0 2 3 1 0 15 9 13 9 2 7 1 15 13 2 16 13 2 9 13 9 2 3 3 1 1 9 9 3 13 9 0 2 7 0 1 9 9 7 9 2 3 13 9 16 9 9 1 15 13 2 7 1 15 9 16 9 13 2
21 7 1 12 15 3 13 13 2 3 13 15 12 13 2 7 12 13 13 9 15 2
29 1 3 9 7 9 13 3 13 2 13 16 1 15 3 13 13 9 2 16 13 1 9 9 2 7 9 1 9 2
32 7 16 9 13 13 1 9 1 9 13 2 16 13 4 2 3 9 13 0 2 7 9 0 2 1 9 15 10 0 9 13 2
57 1 0 13 2 16 9 1 16 13 1 9 2 7 9 1 16 13 9 2 3 13 15 9 9 2 7 1 16 15 13 9 1 9 9 9 13 2 15 13 15 9 2 16 1 9 13 9 13 9 2 7 3 9 1 9 13 2
16 15 3 13 13 16 9 0 2 15 3 13 9 9 15 9 2
43 7 3 9 3 13 13 1 15 12 9 2 16 3 13 9 0 2 16 1 15 13 2 7 1 15 15 9 1 9 2 7 3 1 9 2 16 13 13 1 12 9 9 2
19 3 1 13 2 15 13 9 1 9 0 2 7 13 2 15 13 0 9 2
29 3 3 13 1 15 1 15 15 13 15 1 10 9 2 7 15 13 0 9 2 7 9 2 15 3 13 16 9 2
27 3 9 0 7 0 9 13 0 1 9 0 13 1 9 2 3 7 1 9 9 0 2 15 13 1 0 2
58 7 16 10 9 13 9 0 2 15 13 15 16 13 9 15 2 13 1 9 15 13 15 16 13 9 2 16 9 13 10 9 13 0 1 9 9 2 3 3 0 9 13 9 0 2 1 15 13 9 0 9 2 13 1 0 9 0 2
9 9 3 0 13 1 9 10 9 2
17 7 3 9 0 1 15 13 15 9 7 9 13 0 9 1 9 2
25 1 15 13 16 15 15 13 1 9 16 9 13 9 2 13 1 9 2 16 3 2 16 9 0 2
18 7 3 16 15 13 9 1 9 0 2 3 15 13 1 13 9 9 2
46 7 16 9 0 3 13 9 13 1 15 9 0 2 7 1 9 9 2 16 13 4 2 7 9 13 13 1 15 1 9 9 2 16 13 9 9 1 9 2 1 15 9 3 13 13 2
26 0 2 16 1 9 3 13 9 9 1 0 9 9 2 16 13 1 9 3 0 2 7 1 9 0 2
53 0 2 16 13 1 15 1 9 9 2 7 3 1 0 9 1 9 2 16 9 9 13 1 9 0 3 0 1 9 9 1 9 2 16 3 1 0 9 15 9 7 9 15 13 1 9 2 16 9 13 1 9 2
29 15 12 13 1 9 1 9 2 16 3 1 0 13 9 2 15 13 9 9 2 16 13 16 13 1 9 1 9 2
22 1 0 13 2 16 9 9 15 13 1 9 0 7 0 2 3 13 15 9 1 9 2
23 9 3 0 3 13 1 15 9 1 9 13 2 7 1 15 9 2 16 13 1 12 8 2
27 16 3 13 1 13 10 9 2 15 13 9 7 9 13 2 7 13 15 1 9 1 9 9 1 9 13 2
37 7 15 3 13 13 2 16 16 1 9 13 0 13 9 0 16 9 9 2 3 1 9 9 13 13 0 9 9 2 16 3 13 0 16 13 9 2
5 12 9 1 9 2
43 9 7 13 0 3 9 9 2 7 1 15 13 9 2 15 9 1 15 13 13 2 16 1 0 3 0 13 2 7 9 9 2 7 1 15 13 9 2 15 15 9 13 2
28 7 3 13 15 9 2 16 0 15 13 1 15 9 9 2 16 3 1 0 0 9 3 13 16 13 10 9 2
95 16 3 13 9 0 13 9 2 7 0 9 13 1 9 2 7 13 1 9 13 15 9 1 9 9 15 13 2 3 3 13 10 0 2 2 7 3 1 9 1 9 9 1 9 13 1 9 9 9 1 9 1 9 2 3 1 9 15 1 9 1 9 13 2 0 13 9 2 15 13 1 9 0 9 9 2 0 9 2 15 13 1 9 1 9 2 0 9 15 13 1 9 9 13 2
15 1 9 7 9 1 9 9 7 9 13 3 0 16 9 2
15 13 16 3 13 1 15 9 2 15 13 15 1 9 13 2
9 3 3 13 9 15 1 9 15 2
14 3 15 13 9 9 1 9 13 2 7 1 9 0 2
29 3 13 2 16 9 9 9 13 3 0 1 9 0 7 0 9 2 16 9 1 9 0 13 3 1 9 7 9 2
27 13 3 3 1 9 0 9 1 15 16 13 9 3 2 1 9 7 9 0 1 9 2 7 3 1 9 2
14 1 0 13 2 16 9 13 1 9 9 1 15 13 2
13 1 0 9 13 2 16 9 9 1 9 10 13 2
15 7 3 9 9 13 15 1 15 9 7 9 7 9 13 2
24 7 16 9 9 9 15 13 13 1 0 2 3 15 13 10 9 13 2 16 1 9 13 13 2
53 7 16 3 15 9 15 13 1 9 15 15 3 13 7 15 15 13 0 2 16 1 15 15 13 0 2 9 13 16 13 2 1 15 7 15 3 13 2 0 15 13 2 3 0 9 1 9 7 0 13 9 9 2
15 3 1 3 13 9 13 1 9 9 2 13 16 13 9 2
13 1 0 13 2 16 1 9 13 9 1 13 9 2
8 1 0 3 13 1 9 9 2
7 1 0 13 1 9 9 2
5 0 13 9 9 2
14 0 13 15 9 1 9 9 2 7 13 15 2 3 2
7 1 0 13 9 0 9 2
11 1 0 15 9 0 1 9 13 2 3 2
5 12 1 9 15 2
12 9 13 9 9 0 2 13 1 9 13 9 2
10 3 2 9 7 9 13 1 9 9 2
11 7 15 15 9 13 1 9 7 9 9 2
33 16 7 10 0 3 0 13 9 15 15 13 2 3 9 0 3 13 15 0 13 9 2 7 15 15 13 15 15 13 0 9 15 2
41 7 16 1 9 13 15 9 16 9 13 1 9 2 7 9 1 0 2 7 0 1 9 2 3 9 3 0 13 2 15 13 3 9 9 2 0 7 15 13 9 2
8 3 7 0 13 9 7 9 2
15 3 7 9 0 13 9 7 9 7 0 2 0 7 9 2
32 7 16 9 2 1 13 9 2 15 9 13 2 3 9 0 15 13 15 13 9 7 9 15 7 0 2 7 0 15 13 9 2
13 7 13 9 1 15 15 13 2 1 9 9 13 2
8 7 9 9 13 9 0 9 2
17 7 1 15 9 13 1 9 9 2 1 15 13 9 7 9 0 2
43 16 7 0 3 13 1 9 1 9 0 2 7 1 9 2 3 3 13 16 9 13 1 9 9 16 16 0 13 2 7 13 13 1 9 9 2 2 3 3 13 1 9 2
42 1 0 9 13 2 16 9 15 9 13 7 9 9 1 15 16 13 2 9 2 7 9 1 15 16 13 2 13 9 2 7 9 1 15 16 13 2 1 9 9 13 2
24 1 0 13 2 16 3 3 13 9 2 16 15 15 13 1 9 9 2 15 13 1 9 9 2
40 15 7 9 7 13 15 9 2 16 9 2 7 15 15 9 2 7 3 1 9 13 13 1 9 9 2 7 3 1 15 13 9 2 7 13 9 1 9 13 2
16 0 1 9 1 13 2 1 16 1 9 13 13 13 0 13 2
12 0 3 1 9 15 13 2 15 1 9 13 2
11 0 3 1 9 15 2 15 9 13 9 2
15 3 15 9 2 15 15 13 8 2 13 1 9 9 0 2
23 13 16 9 9 0 3 13 1 15 9 2 15 15 13 1 9 9 7 9 7 9 0 2
46 7 1 9 15 9 13 8 8 12 2 16 13 2 13 10 9 2 3 13 13 16 15 15 13 13 1 9 9 2 16 15 9 13 2 13 3 1 13 9 9 2 3 3 9 9 2
9 3 13 16 3 13 1 9 9 2
14 7 15 9 13 1 9 1 9 2 15 13 9 9 2
16 3 0 13 1 9 9 13 9 1 9 9 16 1 9 9 2
15 13 16 13 15 15 1 15 9 13 2 13 1 9 9 2
7 9 3 15 9 13 13 2
18 3 2 15 15 13 2 15 13 15 2 13 1 9 1 13 9 9 2
13 3 13 13 9 9 2 16 13 2 15 13 15 2
18 7 0 9 13 9 9 2 16 13 1 9 0 2 16 1 8 13 2
8 3 7 3 9 9 13 13 2
13 3 2 12 9 1 9 9 13 1 13 9 9 2
6 3 13 13 9 9 2
19 3 3 13 0 9 1 9 15 13 1 9 9 2 16 1 9 0 9 2
7 3 7 9 9 1 9 2
15 3 2 1 9 0 3 13 16 9 13 7 13 13 9 2
16 3 7 16 1 9 9 15 13 7 13 2 13 9 15 9 2
11 3 2 9 3 13 9 15 16 1 9 2
9 3 3 13 13 7 13 1 9 2
7 3 13 15 1 9 13 2
11 3 2 9 13 13 1 9 1 13 9 2
4 3 13 9 2
34 13 13 1 0 9 2 16 9 0 9 0 13 3 1 9 15 13 2 7 9 0 1 15 13 2 16 9 0 13 9 1 9 13 2
31 7 16 0 13 15 9 15 0 2 3 9 9 13 7 0 0 2 3 9 9 13 2 7 9 9 0 15 13 9 9 2
18 1 0 13 2 16 9 9 3 13 16 9 0 3 2 7 16 0 2
31 7 16 15 13 16 1 16 9 13 2 3 1 9 9 0 13 16 13 15 15 1 9 13 2 16 12 1 15 13 13 2
39 1 0 13 2 16 1 9 15 9 0 3 13 13 9 9 2 16 0 15 13 2 16 13 3 1 9 2 7 13 15 13 9 13 1 9 0 15 13 2
17 7 3 1 9 15 13 0 13 9 13 2 16 3 13 3 13 2
23 7 13 2 16 15 9 13 9 1 15 10 9 3 2 7 9 13 13 9 1 9 9 2
17 7 16 15 9 13 0 2 3 13 16 9 9 13 9 9 13 2
64 1 0 9 13 2 16 16 9 9 13 1 9 0 2 7 0 13 1 9 9 16 3 9 2 3 16 15 13 13 9 2 7 15 0 13 2 3 15 13 13 9 9 3 1 15 15 13 1 9 9 1 0 9 9 0 2 15 9 10 15 9 3 13 2
22 16 7 15 13 1 9 1 9 9 2 16 15 13 2 3 13 9 2 7 9 13 2
23 1 9 7 0 0 13 15 13 9 13 2 1 15 13 15 9 2 16 15 13 9 13 2
21 7 3 3 1 10 9 9 13 1 9 9 2 7 15 3 1 15 9 13 13 2
23 15 0 13 2 16 9 13 3 13 1 9 9 2 7 16 1 15 9 9 9 9 13 2
26 1 0 3 13 2 16 1 9 9 2 1 9 9 13 9 9 3 1 13 2 7 3 3 1 13 2
19 9 7 13 1 9 3 13 1 9 9 2 16 1 15 9 9 3 13 2
14 7 9 13 13 1 9 9 2 16 9 1 13 13 2
11 7 3 13 1 9 1 15 3 1 12 2
10 0 2 16 9 9 1 9 3 13 2
51 3 7 15 13 15 15 13 1 9 9 2 16 3 13 13 2 16 15 13 15 2 3 3 13 13 2 7 0 1 15 2 15 13 16 13 9 9 13 1 9 9 2 7 16 9 9 13 1 9 9 2
57 15 7 0 16 9 15 15 13 2 0 13 2 3 16 9 13 2 16 13 1 13 2 3 16 3 13 9 9 15 9 13 13 2 7 1 9 9 2 15 15 9 13 2 15 3 1 0 9 13 13 2 15 9 1 9 13 2
13 7 3 3 13 2 0 0 2 1 9 9 13 2
18 7 13 15 9 9 2 3 1 9 2 16 0 3 13 16 0 13 2
18 7 3 1 15 3 13 9 9 3 1 9 2 7 0 3 1 9 2
38 1 0 13 2 16 9 15 9 13 2 3 4 1 9 13 3 1 9 2 16 1 0 9 15 9 13 2 16 1 9 13 2 7 0 3 1 9 2
17 7 15 13 15 15 13 2 16 4 13 9 0 2 7 3 0 2
18 7 1 15 9 9 15 13 1 9 15 0 4 13 1 13 9 15 2
41 16 7 9 9 15 9 13 2 3 16 13 9 3 1 0 0 2 3 3 13 3 1 9 2 16 16 9 13 13 15 13 1 9 9 2 13 3 1 9 9 2
34 1 0 9 13 2 16 1 9 15 0 13 2 16 16 13 15 15 13 1 9 9 2 3 13 9 2 7 15 15 13 2 0 13 2
17 7 16 1 10 9 9 13 1 9 9 3 15 15 9 13 13 2
13 7 15 13 2 16 9 9 3 13 1 9 9 2
19 13 3 16 1 9 9 9 13 1 9 13 13 2 15 13 1 9 9 2
19 0 3 9 9 13 13 1 9 9 2 16 1 15 13 9 1 15 9 2
28 7 9 9 13 13 16 3 13 1 9 3 1 9 9 2 7 1 9 9 2 16 9 3 13 1 9 15 2
36 16 16 13 2 13 15 13 1 9 2 3 13 1 15 0 9 13 2 13 16 3 13 13 9 15 13 9 2 7 3 7 13 15 9 13 2
11 16 16 13 0 9 2 3 3 13 9 2
18 16 16 13 2 1 9 9 0 7 9 0 2 13 9 15 9 13 2
23 3 1 15 15 13 9 3 13 2 16 3 13 0 9 2 7 13 3 13 13 9 9 2
12 7 0 1 13 9 7 9 13 9 13 9 2
28 3 16 13 15 1 9 9 13 2 7 13 15 3 1 9 9 2 7 16 13 1 9 9 2 3 13 9 2
14 1 0 13 2 16 9 15 13 9 9 15 13 9 2
5 7 3 13 9 2
33 1 0 13 2 16 1 15 13 3 1 9 9 2 16 15 13 1 9 0 2 16 13 1 9 0 2 16 1 12 9 10 13 2
11 3 13 1 9 9 2 15 13 15 13 2
36 1 0 9 13 2 16 1 9 9 13 1 12 2 3 9 2 9 9 2 7 9 2 15 13 2 16 15 15 13 7 13 2 3 13 9 2
46 7 16 9 9 13 15 9 9 2 9 7 3 13 9 9 16 9 10 9 2 3 15 13 2 16 16 13 9 7 13 7 13 2 3 16 3 13 9 9 7 9 2 15 13 9 2
34 7 16 9 3 1 9 7 9 13 13 15 9 2 3 15 13 0 9 2 16 13 7 9 0 2 7 9 0 15 13 1 9 9 2
23 7 1 15 1 0 13 2 16 16 13 15 9 16 13 9 13 2 3 3 13 12 9 2
45 16 7 3 13 0 9 2 7 9 3 13 9 2 16 16 13 2 1 9 9 0 2 7 9 2 7 9 2 7 15 3 2 16 9 3 13 2 3 13 1 9 9 9 9 2
18 13 3 16 9 9 1 9 9 13 3 13 2 1 9 13 9 13 2
8 7 9 9 0 13 1 9 2
32 7 3 1 9 1 9 9 13 13 13 9 9 7 1 9 9 1 15 16 0 13 2 1 9 2 7 1 9 1 9 9 2
30 1 0 13 2 16 9 0 13 13 15 3 13 9 1 9 2 1 13 0 15 3 13 9 1 9 15 9 15 13 2
9 3 2 9 3 13 1 9 10 2
10 7 9 4 13 1 9 2 8 8 2
29 7 15 9 4 9 13 1 9 12 9 1 9 0 2 16 9 13 1 9 2 9 1 9 2 9 0 1 9 2
27 3 13 2 16 8 8 2 3 4 9 13 1 1 9 1 15 9 13 16 1 9 13 2 7 4 13 2
14 1 7 16 13 1 9 9 2 13 3 9 3 13 2
23 7 3 13 9 2 7 1 15 13 9 2 16 9 13 9 9 2 9 7 3 13 9 2
22 15 7 13 3 13 2 16 9 1 9 15 9 7 9 13 2 13 15 1 9 13 2
11 0 3 15 13 1 15 16 1 15 9 2
15 3 13 16 15 15 9 15 13 9 2 13 15 9 13 2
29 7 1 3 13 9 0 2 16 9 0 1 9 3 13 2 13 16 9 13 13 9 15 2 15 9 9 9 13 2
7 7 9 15 9 9 13 2
36 1 0 13 2 16 16 1 12 9 13 0 9 2 1 15 9 13 0 12 9 3 13 7 13 15 1 9 15 2 7 15 13 3 9 15 2
33 13 13 1 0 9 2 16 1 9 15 1 9 9 10 0 9 13 2 7 3 9 1 9 0 2 16 3 13 1 9 13 9 2
14 7 15 3 13 9 9 2 3 13 9 2 7 13 2
18 7 15 15 13 9 3 13 9 2 16 3 13 13 9 7 13 9 2
48 13 13 1 0 9 2 16 0 13 2 12 13 3 9 2 15 1 9 13 1 13 9 9 2 1 15 9 13 8 8 2 12 2 13 10 9 2 13 15 1 9 9 7 9 7 9 0 2
13 3 2 1 9 0 13 9 0 16 15 9 0 2
17 3 2 10 9 15 9 13 13 9 15 2 16 9 13 1 0 2
14 7 3 3 13 16 9 0 13 2 15 3 13 9 2
11 1 0 13 2 16 13 0 9 9 15 2
12 0 3 9 3 13 13 9 2 7 0 0 2
8 3 2 9 13 0 16 9 2
10 7 15 9 13 4 16 13 13 9 2
27 1 0 13 2 16 15 9 13 13 9 2 16 9 3 13 16 13 1 12 8 2 7 13 1 9 9 2
10 7 3 3 13 0 1 9 7 9 2
32 7 15 13 0 2 3 16 15 9 2 1 9 2 15 13 16 13 2 9 7 9 15 13 2 7 16 3 13 13 9 9 2
16 3 3 13 13 13 2 16 13 9 9 2 7 13 9 13 2
13 16 3 1 9 13 9 7 9 2 3 7 9 2
12 7 16 13 9 0 7 9 2 3 13 9 2
31 9 7 0 2 1 13 15 0 2 13 16 13 9 2 15 13 1 10 9 1 9 0 2 7 15 0 1 9 3 0 2
47 7 9 0 3 13 16 13 9 15 13 16 13 15 2 7 0 1 9 9 2 16 1 9 9 1 9 13 2 16 1 12 8 2 8 12 2 8 12 2 8 12 7 12 2 13 4 2
34 15 3 13 13 9 2 16 1 15 3 13 9 1 9 2 1 13 12 9 7 12 9 2 7 13 3 1 9 2 16 7 3 13 2
7 7 0 3 1 9 9 2
24 7 15 9 13 2 16 1 0 9 13 1 15 9 2 16 3 13 13 2 15 15 13 8 2
17 1 9 7 9 13 0 13 2 3 9 2 9 9 2 7 9 2
37 15 7 3 13 13 1 3 16 13 12 9 2 16 1 9 13 2 15 3 9 1 9 13 2 10 0 9 1 15 2 7 15 15 1 9 9 2
28 7 0 3 1 10 15 9 13 9 9 1 13 9 7 9 2 3 0 1 9 9 13 2 7 1 9 9 2
32 15 13 2 16 1 9 7 1 15 9 15 13 1 9 9 13 2 3 13 0 9 2 7 13 9 9 1 9 1 9 13 2
18 7 3 16 9 13 2 7 15 0 13 15 9 0 13 2 13 13 2
67 1 0 13 2 16 16 9 9 13 13 1 13 9 10 3 13 2 16 0 1 9 0 9 9 13 0 2 16 3 9 13 3 0 2 3 16 3 3 13 0 9 16 9 13 2 16 0 13 2 7 0 9 3 13 2 9 3 13 2 16 13 3 1 9 0 9 2
55 1 0 9 13 2 16 16 0 7 15 0 13 9 13 2 7 9 13 13 2 0 9 13 2 16 9 3 13 9 1 9 13 2 7 1 9 0 2 15 13 1 13 1 9 0 1 13 2 7 1 9 9 1 9 2
24 3 16 13 9 2 1 15 9 0 3 13 2 16 13 1 9 9 2 13 9 7 9 9 2
38 3 16 13 1 0 15 9 13 1 9 15 15 13 1 9 9 2 13 0 3 13 1 15 9 2 13 15 2 16 3 13 13 2 1 9 9 8 2
36 16 7 13 2 15 13 15 2 3 13 9 2 16 3 13 13 9 2 16 1 2 8 12 2 8 12 2 8 12 2 8 12 2 13 4 2
36 0 3 13 9 2 16 12 13 0 7 15 0 2 12 13 9 2 7 15 13 2 16 15 9 9 13 16 1 15 13 13 9 7 9 9 2
20 16 16 9 13 13 2 13 13 9 9 2 15 15 3 13 13 15 9 13 2
12 1 9 7 9 1 2 8 12 2 13 4 2
17 1 0 13 1 9 9 15 15 1 15 13 1 9 15 9 13 2
15 1 0 13 15 15 13 1 9 9 2 3 9 7 9 2
4 12 1 9 2
41 7 13 16 1 9 7 1 9 9 3 13 9 1 9 7 9 15 9 2 16 9 0 7 15 15 1 9 13 13 13 1 0 9 1 9 0 2 16 9 13 2
13 3 3 1 9 8 8 13 15 1 9 9 0 2
41 1 0 13 2 16 16 9 9 2 3 9 2 13 9 9 1 0 9 2 3 15 9 3 13 3 1 9 2 7 1 9 9 2 7 9 2 16 7 9 9 2
9 3 2 9 9 15 0 9 13 2
20 7 1 9 9 13 9 2 16 13 1 9 2 15 9 13 9 9 9 13 2
13 15 9 1 2 8 12 2 13 9 13 9 9 2
14 3 3 13 1 9 9 0 15 9 1 9 9 13 2
20 7 3 13 2 16 9 9 3 13 15 9 2 7 9 9 1 9 13 9 2
23 15 7 9 0 9 3 13 9 9 2 7 3 13 15 9 0 2 16 9 9 7 9 2
35 1 0 13 2 16 16 9 9 0 13 0 2 3 16 13 9 9 2 7 16 13 1 0 9 1 9 2 3 3 9 9 0 9 13 2
13 15 13 16 13 1 9 2 15 13 1 9 9 2
6 3 9 9 13 9 2
8 13 16 9 9 3 13 9 2
11 7 0 3 13 15 9 13 2 9 13 2
17 3 1 15 9 9 9 13 2 13 16 9 9 3 13 15 9 2
27 3 1 3 13 15 1 15 9 9 9 13 2 16 13 1 9 0 13 2 13 16 15 9 3 13 9 2
14 3 2 9 15 13 9 2 1 15 9 1 10 13 2
8 3 15 9 3 13 15 9 2
6 9 7 1 9 13 2
9 13 16 15 9 9 3 13 13 2
14 7 1 13 9 1 9 9 13 9 13 15 9 15 2
11 3 7 1 9 9 15 9 15 13 13 2
20 1 3 1 9 15 13 9 1 9 1 9 2 7 3 13 13 1 15 9 2
12 7 1 9 9 3 13 9 15 1 0 9 2
11 3 7 1 9 15 13 13 9 1 9 2
12 3 2 16 9 13 9 13 2 3 7 9 2
11 7 1 9 9 3 13 9 1 9 15 2
18 3 2 9 13 1 9 9 2 16 0 13 9 15 3 13 9 9 2
16 3 3 13 9 9 13 1 9 2 16 3 13 2 9 9 2
12 13 16 9 15 3 13 1 15 9 15 9 2
11 7 9 15 9 13 13 3 1 9 9 2
8 3 9 9 15 9 13 9 2
31 7 3 15 9 9 13 1 9 13 2 16 13 1 9 9 15 13 2 1 15 9 13 2 1 13 2 9 9 10 8 2
14 7 1 13 2 16 9 13 0 1 9 16 1 9 2
10 16 3 9 15 13 2 0 0 9 2
18 7 3 1 16 1 15 9 13 9 2 3 13 9 15 9 9 13 2
29 16 3 9 13 1 9 7 9 2 3 13 9 2 16 15 13 9 9 1 9 2 15 13 9 9 1 0 13 2
24 1 0 13 2 16 15 13 16 9 1 9 7 9 15 13 1 9 7 9 1 0 9 9 2
15 7 3 13 2 16 9 15 9 13 2 16 3 4 13 2
27 0 2 16 9 1 9 13 9 9 0 2 16 15 3 1 15 8 13 2 16 13 9 9 16 9 13 2
30 1 0 13 2 16 9 9 1 15 15 3 13 1 9 9 2 13 13 1 0 9 9 2 16 9 9 1 10 13 2
13 7 3 1 15 3 13 16 15 9 13 13 9 2
30 1 0 9 13 2 16 16 9 13 13 15 9 9 2 16 13 9 2 3 1 9 9 13 13 15 15 1 9 13 2
9 7 3 12 13 1 9 15 9 2
13 7 3 3 13 15 9 9 1 9 1 9 13 2
33 1 0 13 2 16 9 15 13 1 9 2 3 13 1 9 9 2 7 1 9 9 2 15 13 1 9 9 9 1 9 9 9 2
14 7 3 0 1 0 13 9 9 2 7 1 9 13 2
13 1 0 9 13 2 16 9 9 13 1 13 9 2
44 7 3 1 15 9 15 15 13 1 15 9 0 13 2 7 3 1 9 15 9 2 9 9 13 15 15 9 13 2 3 7 15 9 15 1 9 9 13 2 16 13 1 9 2
40 1 15 7 9 15 13 1 9 9 2 16 9 1 15 9 7 9 2 9 9 13 15 13 1 9 9 2 3 15 13 1 9 9 2 16 15 0 15 13 2
37 7 3 1 9 9 2 16 13 4 2 13 1 9 9 2 13 16 15 9 15 13 9 13 2 13 9 9 2 7 13 9 16 7 15 9 9 2
12 7 3 9 9 15 13 9 13 1 9 9 2
13 16 1 15 9 7 9 3 13 13 16 12 9 2
24 1 0 3 13 2 16 1 12 9 7 9 2 15 15 9 13 2 3 13 13 16 12 9 2
16 7 15 15 13 9 7 9 1 9 13 15 9 1 13 13 2
16 7 15 2 3 3 13 2 13 9 13 15 13 9 15 9 2
18 3 2 15 13 13 1 9 15 13 2 16 15 13 1 15 13 9 2
29 7 13 9 15 16 13 9 9 2 16 1 0 1 15 16 9 15 1 15 9 13 1 15 9 2 13 9 0 2
64 1 0 9 13 2 16 1 10 9 7 9 13 2 7 9 2 3 13 16 0 9 13 13 1 0 9 1 9 15 2 16 9 15 13 1 9 9 2 13 9 9 9 0 2 15 9 13 2 7 15 13 0 9 2 3 9 9 2 9 0 2 3 0 2
24 7 3 9 13 13 2 16 1 9 15 13 2 7 3 13 16 9 13 9 10 13 1 15 2
21 7 15 15 13 9 7 9 2 13 15 9 13 1 13 9 2 16 13 1 9 2
17 1 0 13 13 2 15 15 9 13 2 3 9 7 9 2 3 2
6 1 0 9 2 3 2
8 9 0 13 15 15 3 13 2
5 0 1 9 15 2
9 3 2 9 9 13 1 9 10 2
17 7 1 9 13 12 9 2 12 1 9 9 2 15 1 9 9 2
17 9 3 13 9 9 2 3 15 13 2 16 13 9 1 12 8 2
26 3 9 15 13 9 0 1 15 13 2 13 3 13 9 0 2 7 9 1 9 2 7 9 9 0 2
11 7 0 9 13 15 13 9 13 10 9 2
32 1 0 13 2 16 9 15 13 1 9 15 9 2 3 13 9 9 0 2 7 1 9 1 15 2 16 1 12 8 13 4 2
26 7 16 1 9 9 0 13 2 16 9 7 9 2 7 3 2 3 1 15 9 9 13 9 12 13 2
16 1 0 13 2 16 9 15 13 2 16 15 9 13 15 9 2
20 7 15 0 13 2 16 12 9 13 12 2 7 15 15 15 15 1 9 13 2
18 7 9 4 13 1 0 9 2 16 9 9 9 13 13 2 8 8 2
46 1 0 13 2 16 9 15 13 1 9 15 15 15 1 9 13 13 2 15 9 13 1 9 2 3 7 1 15 15 13 1 9 1 9 9 2 15 13 1 9 2 16 1 13 4 2
16 7 9 13 15 15 9 13 1 9 9 2 16 9 7 9 2
20 1 0 3 13 2 16 9 7 9 4 13 1 9 13 15 9 3 0 9 2
7 3 13 1 9 15 9 2
8 12 1 9 15 9 0 13 2
8 12 1 9 15 13 15 9 2
12 3 15 13 9 9 2 3 15 13 9 10 2
14 13 16 15 3 13 9 9 9 2 15 13 9 10 2
10 3 1 13 9 3 13 9 9 9 2
14 3 2 9 9 13 1 9 15 13 1 15 9 9 2
10 3 1 15 9 3 13 9 15 9 2
15 13 16 3 3 1 15 9 13 9 2 15 13 9 10 2
10 3 15 3 13 9 2 13 7 13 2
26 3 2 15 15 3 13 1 9 9 2 3 13 13 1 0 9 2 1 15 9 2 16 3 1 15 2
13 3 15 3 13 1 9 2 7 3 3 9 13 2
8 13 16 9 15 3 13 13 2
36 1 9 3 9 13 13 15 15 1 9 13 1 9 13 9 2 16 1 9 9 13 2 15 15 13 2 7 1 9 9 2 13 15 9 9 2
6 3 3 13 13 9 2
11 7 1 9 15 9 13 15 13 1 9 2
15 3 1 1 15 9 3 13 9 9 2 13 16 13 0 2
18 7 9 9 3 13 16 1 15 16 9 9 13 1 9 1 9 13 2
16 7 1 9 9 9 13 2 13 9 1 9 2 7 13 9 2
12 13 16 9 15 1 9 13 2 3 13 13 2
33 13 13 1 0 9 2 16 1 9 15 9 13 16 13 15 1 15 9 9 13 2 16 1 9 9 9 13 2 15 9 13 9 2
9 7 3 15 9 13 9 15 9 2
32 15 3 13 2 16 0 2 15 13 9 9 1 9 2 1 10 9 9 0 13 2 7 3 9 13 2 1 15 15 3 13 2
27 7 15 9 13 9 2 13 2 0 13 13 2 16 0 9 0 13 2 7 3 9 13 1 15 0 13 2
24 7 3 15 13 2 16 13 3 1 15 9 9 2 3 7 1 15 2 7 1 15 9 0 2
12 0 13 2 1 13 2 16 9 13 15 13 2
26 7 3 15 13 2 7 0 2 16 0 15 3 3 13 2 7 15 3 13 13 2 7 9 13 13 2
16 7 3 9 3 1 15 9 13 1 9 15 13 1 9 9 2
15 1 15 7 9 9 13 1 9 15 13 1 9 9 13 2
29 3 15 9 15 1 9 13 2 3 13 1 9 2 7 3 15 15 1 9 9 13 2 3 2 15 13 9 10 2
23 7 3 3 13 13 1 9 3 0 15 15 13 1 9 2 7 3 15 15 13 1 9 2
19 7 3 16 9 15 13 1 9 2 3 13 1 9 2 3 7 13 9 2
14 9 3 9 15 9 13 1 9 1 9 0 3 0 2
9 15 7 9 9 1 9 9 13 2
18 7 3 3 13 13 15 15 3 13 1 9 9 9 2 1 0 13 2
52 3 1 15 9 1 15 15 9 9 13 2 13 16 9 13 13 9 13 2 7 9 0 13 0 9 2 16 1 9 13 2 16 9 0 2 15 9 9 13 2 13 0 9 2 15 0 9 13 1 9 13 2
14 3 13 16 9 9 13 15 15 9 0 1 9 13 2
22 7 3 15 13 13 9 1 9 2 15 13 9 10 2 15 15 15 13 4 2 13 2
31 16 7 1 9 9 7 9 13 1 13 7 13 9 1 9 0 7 0 2 3 1 9 0 13 9 7 9 1 9 9 2
25 3 15 3 13 13 9 15 9 2 15 13 9 10 2 16 1 15 3 13 15 13 7 3 13 2
16 3 1 15 9 0 13 13 9 9 15 2 16 1 9 0 2
16 7 3 9 9 1 9 15 13 1 9 9 2 13 3 13 2
28 1 0 9 13 2 16 2 16 13 4 2 9 9 9 1 10 9 13 13 2 3 1 16 13 16 1 13 2
22 7 3 1 9 9 13 12 9 9 2 7 15 9 16 13 1 10 9 1 9 13 2
39 1 9 7 9 1 15 2 13 9 13 9 9 2 7 9 3 0 15 9 16 13 1 9 2 7 16 13 0 1 0 9 0 2 16 3 9 9 13 2
16 3 13 16 0 1 15 9 12 9 13 2 15 13 9 10 2
47 7 15 3 13 3 13 2 16 1 1 9 3 13 16 15 13 9 13 9 2 3 13 9 0 1 9 1 9 2 7 1 9 3 2 15 13 0 2 7 9 13 3 13 9 15 9 2
22 7 16 13 15 9 15 2 3 13 4 9 2 16 3 15 9 3 13 1 9 9 2
38 16 7 1 0 9 0 15 9 13 9 7 9 2 13 7 9 1 9 0 7 0 2 3 1 9 0 13 9 0 2 15 13 2 9 7 13 9 2
13 7 1 9 9 13 13 7 9 9 7 9 15 2
26 1 0 13 2 16 2 16 13 4 2 15 9 2 13 7 13 1 15 10 2 3 13 1 9 9 2
16 3 9 9 9 13 1 15 3 9 2 15 13 9 9 10 2
45 13 16 9 9 9 13 1 15 3 9 2 15 13 9 9 10 2 7 15 15 13 2 0 7 0 9 2 9 9 2 15 1 15 7 1 0 13 1 9 9 3 13 1 9 2
25 9 3 13 13 1 15 15 13 1 9 9 15 9 2 16 9 9 15 9 0 13 1 9 0 2
8 3 3 13 1 9 15 9 2
9 3 9 15 13 3 13 1 9 2
22 3 1 15 9 15 13 13 15 9 9 1 15 13 9 2 13 16 3 13 1 9 2
15 7 1 13 16 8 12 2 12 2 13 13 9 9 9 2
32 3 15 13 1 9 9 2 16 9 3 13 9 1 1 9 15 2 15 3 13 2 15 3 13 1 9 2 16 13 9 9 2
21 3 2 1 9 13 1 9 9 13 13 9 1 15 13 9 2 16 1 13 13 2
8 3 3 13 13 1 9 13 2
16 3 2 1 9 9 3 13 13 15 15 3 13 1 9 9 2
8 3 3 13 13 1 9 9 2
16 3 2 15 15 13 13 9 9 2 3 13 13 1 9 9 2
6 3 9 13 1 9 2
20 1 3 15 3 13 1 9 9 13 2 7 1 9 9 1 9 13 9 13 2
11 7 1 9 9 3 13 9 1 9 9 2
11 15 3 13 2 16 15 13 3 1 9 2
13 15 13 9 9 10 2 16 9 15 9 13 0 2
30 3 15 0 13 2 16 15 15 13 2 13 1 9 2 1 15 15 15 13 3 13 9 1 15 2 7 13 9 9 2
17 9 3 3 13 9 7 9 9 13 2 7 13 7 13 9 13 2
9 7 3 13 16 13 1 9 9 2
29 3 7 15 9 9 0 13 9 15 2 16 9 1 15 9 3 13 15 0 2 3 3 15 15 9 13 1 9 2
11 7 15 9 13 3 13 13 1 15 9 2
14 9 7 3 13 9 3 1 9 2 7 3 1 9 2
23 7 16 9 0 13 1 9 2 3 2 9 13 2 1 0 1 9 9 13 9 9 13 2
35 1 9 7 2 9 7 9 2 15 13 3 15 1 13 4 1 9 9 2 8 12 2 8 12 2 8 12 2 8 12 2 12 7 12 2
13 3 3 13 1 9 13 9 9 13 3 9 13 2
31 7 1 9 13 13 1 9 2 7 9 9 0 13 2 16 13 9 2 9 15 3 13 3 13 2 16 1 15 0 15 2
20 3 1 9 9 3 13 13 2 9 13 2 16 15 9 13 13 4 1 9 2
28 7 1 13 15 9 13 1 9 8 8 2 1 15 2 3 0 9 2 3 9 9 2 13 9 0 1 9 2
8 7 9 13 13 9 0 9 2
16 9 7 0 13 9 13 1 0 13 2 7 1 15 9 13 2
23 7 3 13 13 2 16 1 9 13 2 16 7 1 15 9 9 2 13 15 9 1 9 2
53 7 15 9 3 13 9 13 9 0 1 9 2 15 13 9 15 0 9 1 9 10 2 7 13 9 0 2 16 9 15 13 1 9 1 9 0 9 2 7 16 9 9 1 9 2 16 1 2 8 12 13 4 2
7 3 9 13 15 1 13 2
8 13 16 9 13 15 1 13 2
15 16 3 15 13 9 1 9 2 3 15 13 9 1 9 2
9 3 7 9 9 13 1 9 9 2
11 3 0 12 9 15 13 1 9 12 9 2
15 7 1 12 9 9 15 13 3 1 13 2 16 13 4 2
8 3 7 9 9 13 9 9 2
9 3 9 0 3 13 0 1 13 2
23 7 1 0 9 9 2 3 13 0 9 9 1 9 2 1 9 9 13 9 1 9 13 2
8 3 1 9 9 9 4 13 2
26 3 1 9 13 2 15 9 9 13 1 9 0 2 3 2 15 3 16 13 8 2 3 13 13 9 2
15 7 9 9 1 13 0 13 15 15 1 9 15 13 13 2
22 13 13 1 0 9 2 16 15 13 2 16 0 9 3 13 9 10 16 13 9 0 2
12 7 15 3 13 13 2 16 9 9 13 13 2
15 3 16 9 13 13 7 1 3 13 2 3 9 13 13 2
16 7 3 13 1 15 2 16 9 13 3 13 15 0 1 13 2
28 1 0 13 2 16 12 9 1 15 9 3 13 1 12 9 16 12 9 13 2 16 1 0 9 13 12 9 2
14 7 0 9 13 1 0 2 15 13 9 7 9 3 2
42 1 0 9 13 2 16 15 13 16 9 15 2 1 15 9 13 2 16 13 4 2 16 1 15 13 1 15 2 3 13 9 2 1 0 1 15 15 13 1 9 9 2
33 1 0 13 2 16 1 15 9 13 13 9 9 1 9 0 13 2 3 9 15 3 13 2 16 9 9 13 1 9 0 13 13 2
19 7 3 15 3 13 1 9 2 16 13 4 1 2 8 12 2 8 12 2
11 7 1 2 1 9 15 9 13 9 9 2
59 7 16 1 15 3 13 16 9 0 2 15 1 15 9 0 15 13 2 16 9 1 0 9 12 9 2 3 16 9 3 13 2 15 9 13 3 13 9 0 2 16 7 1 9 0 9 13 13 13 1 9 2 16 9 1 9 15 13 2
29 7 15 13 2 16 9 1 15 9 3 13 9 9 2 7 9 1 9 9 2 3 9 2 7 9 2 3 9 2
18 3 9 15 15 13 9 2 1 15 3 13 2 16 1 12 8 13 2
34 9 7 0 13 1 9 1 0 3 13 2 16 9 13 4 1 15 2 3 16 15 15 9 13 9 1 15 9 2 16 3 13 9 2
14 3 3 13 9 1 15 16 9 2 7 1 15 0 2
8 3 2 9 9 13 13 9 2
14 7 1 9 3 13 9 1 9 2 7 0 1 9 2
14 7 12 13 9 9 0 7 9 2 16 9 7 9 2
10 0 1 9 9 2 15 9 13 9 2
60 1 15 3 13 16 1 9 0 3 13 9 1 9 9 2 7 1 9 9 1 9 13 9 2 7 9 13 1 9 9 2 15 13 13 7 13 2 1 9 3 13 9 9 7 9 2 7 1 9 7 9 0 2 15 1 9 13 3 13 2
24 9 7 3 13 13 2 16 9 9 3 13 3 16 9 0 13 1 9 2 7 13 1 9 2
29 16 7 13 9 0 13 1 9 2 7 13 13 9 2 16 9 15 13 1 9 2 7 13 9 2 16 9 0 2
57 16 7 13 13 9 2 13 1 7 1 2 7 15 1 15 2 7 15 1 9 2 16 15 9 0 9 13 1 15 9 15 2 16 9 9 0 3 13 9 9 2 16 13 1 9 9 0 2 15 13 1 9 2 7 13 15 2
31 7 1 15 9 15 13 15 1 15 15 2 7 15 1 9 15 2 3 13 1 9 0 13 3 0 9 2 7 0 9 2
15 12 9 16 1 9 13 1 9 2 16 9 13 1 9 2
25 1 0 13 2 16 9 1 15 9 3 13 2 16 9 3 13 13 1 9 2 7 1 9 0 2
16 7 3 1 9 0 13 3 0 2 1 9 9 3 13 9 2
13 13 13 1 15 2 3 1 16 13 1 9 10 2
15 9 7 13 13 15 9 0 2 1 16 1 0 9 13 2
21 9 7 0 1 9 15 9 13 9 0 2 1 15 1 2 8 12 2 13 4 2
12 3 7 13 13 1 9 13 2 3 9 9 2
9 13 16 3 9 0 9 13 13 2
10 9 3 0 3 13 13 1 9 0 2
20 7 13 13 9 9 0 2 16 13 16 15 9 2 16 13 1 12 1 9 2
24 3 1 9 15 1 9 13 2 3 0 13 2 16 1 15 13 2 13 16 9 0 9 13 2
40 7 9 0 9 3 13 1 15 9 0 2 16 16 13 2 13 16 13 1 9 2 15 13 9 0 9 0 2 1 15 3 13 15 2 16 1 13 8 13 2
8 3 9 0 9 13 16 9 2
12 7 9 0 13 9 2 16 13 1 12 8 2
16 1 3 9 13 2 13 16 9 9 1 15 13 9 2 13 2
49 3 2 1 9 1 8 1 9 9 2 7 1 12 8 2 13 1 9 13 9 1 9 0 15 9 1 0 7 0 2 15 3 13 13 0 9 1 0 9 9 2 1 9 3 13 16 1 9 2
6 3 7 9 0 13 2
15 7 1 2 13 9 7 9 0 2 15 13 16 9 0 2
12 3 3 13 13 15 9 13 16 9 0 13 2
24 7 16 13 3 9 0 9 2 13 1 15 3 16 1 9 0 2 16 13 15 0 1 9 2
9 3 13 16 3 13 9 0 9 2
14 1 0 9 13 2 16 9 9 0 3 13 1 9 2
21 15 7 1 15 13 9 2 3 13 9 3 7 9 3 2 7 9 13 1 9 2
7 7 3 9 9 3 13 2
15 7 9 0 3 13 15 0 2 7 13 13 1 9 0 2
13 3 1 9 9 3 13 2 3 9 0 3 13 2
18 0 2 16 9 3 0 13 1 9 0 2 7 1 9 0 9 13 2
16 1 0 3 13 2 16 15 9 13 15 1 13 9 0 13 2
16 7 13 16 9 15 3 13 13 16 9 9 13 16 16 9 2
34 15 7 0 9 13 1 15 2 3 13 3 1 9 2 7 3 1 9 2 3 9 0 9 2 16 13 2 13 3 13 3 16 9 2
21 1 0 13 2 16 9 3 13 9 15 13 0 10 0 1 15 7 1 10 9 2
55 3 16 1 9 0 1 16 13 9 15 2 3 13 15 2 3 13 9 9 15 2 7 3 1 9 7 3 1 9 1 15 9 0 15 2 1 16 13 13 13 9 1 0 9 2 16 3 13 0 2 7 0 9 9 2
45 1 0 13 2 16 16 9 3 13 13 9 0 1 15 2 13 3 13 9 9 15 13 1 10 9 16 9 2 16 13 1 15 16 9 1 9 13 2 7 9 1 9 9 13 2
21 7 0 1 13 9 2 13 9 2 15 9 0 13 2 16 9 12 13 9 15 2
25 3 3 1 9 9 7 9 7 9 9 13 13 9 15 0 15 13 9 0 1 15 9 13 9 2
26 16 7 3 13 9 0 15 4 1 9 13 1 15 9 13 9 2 13 9 0 0 2 3 9 9 2
25 1 0 13 2 16 9 15 13 1 9 0 1 9 2 3 13 9 0 2 16 3 13 9 13 2
7 9 3 9 13 1 9 2
28 7 16 1 9 13 9 2 9 9 2 15 13 9 1 15 2 3 13 16 1 9 9 0 2 15 13 9 2
31 3 1 3 13 13 15 13 1 15 9 9 2 16 3 13 1 9 16 9 2 7 1 9 16 9 2 13 16 3 13 2
15 3 2 16 15 13 9 0 1 9 2 3 0 1 9 2
15 7 1 9 0 13 9 2 16 13 1 1 9 13 9 2
26 12 9 16 13 1 9 1 9 10 2 15 3 7 1 9 13 13 2 16 15 9 13 1 15 9 2
16 9 3 1 9 10 13 9 1 9 2 7 9 13 9 15 2
17 16 3 13 9 1 9 13 9 2 13 9 9 13 7 3 13 2
25 1 0 3 13 2 16 1 9 0 9 1 15 13 9 15 2 15 3 3 13 1 9 1 15 2
16 15 0 9 13 15 13 1 1 9 0 2 16 9 7 9 2
13 9 3 3 13 2 16 13 15 2 7 15 13 2
39 7 3 7 15 13 1 15 2 16 9 13 9 0 2 7 9 3 13 2 16 9 9 13 9 9 0 2 7 9 0 0 13 15 9 15 13 9 0 2
29 3 13 16 9 9 0 13 15 15 13 9 3 9 9 2 3 9 2 1 15 13 9 2 7 3 15 3 9 2
18 3 3 13 9 16 1 0 9 1 15 9 3 13 16 1 1 9 2
52 7 3 16 15 13 13 9 13 2 9 3 13 1 9 2 13 9 2 16 13 1 9 0 2 1 1 15 3 13 15 0 7 13 9 2 7 0 1 9 3 13 16 9 13 13 2 0 9 1 15 13 2
47 16 7 9 13 9 1 13 1 15 9 9 3 13 15 13 2 3 15 9 13 13 0 9 2 16 3 13 10 15 9 13 2 16 15 13 1 9 2 13 0 2 7 3 0 9 0 2
74 1 7 9 1 15 13 2 1 15 9 9 13 2 16 13 4 2 1 15 13 1 9 9 7 9 2 12 9 3 3 13 1 12 16 1 15 2 3 13 13 0 7 0 9 1 9 2 16 15 0 13 2 3 1 15 15 13 1 9 0 2 3 13 1 15 0 10 9 3 1 0 15 9 2
12 1 0 3 13 2 16 9 9 13 0 9 2
20 7 3 2 1 9 15 9 3 13 9 16 1 0 9 2 3 13 9 10 2
39 3 1 10 9 2 1 15 13 9 7 9 3 2 7 9 7 9 3 2 1 15 13 2 3 13 13 9 1 9 7 9 1 9 1 9 1 0 9 2
40 7 16 9 7 15 9 13 1 1 9 9 2 16 1 13 13 2 13 15 9 13 0 9 0 15 15 2 1 15 13 7 9 0 7 0 2 7 9 0 2
28 16 3 1 9 0 13 9 9 1 13 15 9 2 3 1 15 0 9 13 9 9 16 15 9 13 1 15 2
36 3 3 13 16 13 13 15 9 15 13 1 9 3 2 7 15 13 1 9 2 16 15 9 9 0 13 2 13 16 9 13 13 13 1 9 2
14 1 15 7 9 13 2 1 2 8 12 2 13 4 2
12 3 2 9 9 3 13 3 0 9 16 9 2
10 7 9 1 9 9 13 9 1 9 2
12 15 7 13 2 16 9 4 13 1 15 9 2
54 1 0 9 13 2 16 9 3 13 13 16 9 0 1 9 13 13 1 9 2 13 1 9 16 13 9 1 9 2 16 15 13 9 1 1 2 7 3 16 13 15 13 1 9 16 9 2 16 15 13 1 9 0 2
27 7 16 9 0 0 13 2 0 13 13 9 15 7 9 3 1 9 9 2 7 1 15 9 9 0 13 2
8 3 2 9 13 13 9 13 2
15 7 1 9 9 9 3 13 16 13 9 9 1 9 9 2
16 3 2 9 3 13 16 1 9 2 16 7 9 16 1 9 2
17 3 2 10 9 13 1 9 13 9 1 9 2 16 1 9 13 2
14 7 16 9 13 3 1 9 2 13 15 9 1 9 2
18 15 9 13 16 13 3 9 0 2 7 1 15 13 10 9 15 13 2
16 7 3 0 0 13 0 9 0 1 9 13 16 9 1 9 2
10 7 3 9 3 13 9 16 9 9 2
6 3 9 0 9 13 2
24 7 3 2 1 15 9 13 9 13 1 9 2 3 13 9 13 1 9 2 9 0 9 13 2
15 9 3 13 1 8 1 8 16 9 0 9 13 3 13 2
24 7 15 12 13 12 9 0 9 2 3 9 7 9 2 3 0 7 0 9 13 9 9 2 2
6 7 9 1 9 9 2
44 7 16 9 13 9 0 15 3 13 1 15 2 9 7 13 1 15 2 3 9 2 3 3 13 1 15 15 13 3 13 1 15 2 9 16 9 2 7 1 13 16 15 9 2
21 7 3 0 9 9 13 9 2 15 13 13 1 9 15 15 9 7 0 7 0 2
18 3 1 13 9 0 13 15 13 9 16 1 9 2 15 13 9 9 2
28 7 1 15 1 9 13 15 9 15 9 2 16 1 13 9 7 9 0 1 15 2 13 13 1 9 7 9 2
19 7 16 9 0 13 2 15 3 13 3 13 9 3 2 7 9 1 9 2
11 3 3 13 13 1 9 15 13 9 3 2
10 7 10 13 13 9 1 9 7 9 2
16 1 3 9 15 13 9 3 2 3 13 13 13 15 1 15 2
20 7 15 9 13 9 1 12 8 1 9 2 15 13 9 13 13 9 9 0 2
7 16 15 9 13 9 3 2
14 7 9 13 0 9 13 2 16 13 1 8 12 9 2
9 7 3 9 13 9 1 9 0 2
16 3 2 16 15 9 1 0 9 9 13 2 3 7 9 13 2
16 7 3 9 15 13 1 9 0 1 9 9 2 15 0 13 2
30 7 3 7 9 13 7 9 2 7 9 2 15 3 3 13 9 9 2 7 9 9 2 15 13 9 2 7 9 9 2
30 7 16 9 15 13 1 9 9 2 7 9 1 9 9 2 3 9 3 13 16 13 9 2 15 13 1 15 9 9 2
29 1 0 9 13 2 16 1 9 0 9 0 3 13 0 9 9 2 7 13 13 9 0 7 0 2 16 0 9 2
17 7 3 9 3 0 13 1 9 0 2 7 3 1 9 9 0 2
16 3 9 15 3 0 13 1 9 0 2 7 3 1 9 0 2
15 7 3 2 16 1 13 13 1 9 0 2 3 7 3 2
32 1 0 3 13 2 16 15 3 13 3 3 9 13 2 16 9 13 9 0 2 1 13 1 9 15 15 13 0 9 15 0 2
16 9 7 9 13 3 13 0 13 2 7 0 9 9 7 0 2
21 7 9 15 2 15 13 9 2 13 13 1 9 10 2 16 9 13 1 9 9 2
17 1 0 3 13 2 16 9 13 13 0 2 16 3 13 9 9 2
22 7 3 15 13 1 9 1 15 13 16 9 1 9 0 2 7 15 13 16 9 9 2
24 13 3 15 9 9 1 9 15 2 16 9 13 9 9 2 7 9 9 9 2 16 13 4 2
30 16 9 13 13 3 1 9 3 2 16 15 15 9 15 0 13 1 9 9 2 3 13 1 9 9 2 7 15 3 2
29 16 3 9 13 1 12 8 2 7 1 8 1 9 9 2 1 9 0 7 0 13 13 9 0 1 9 9 0 2
17 15 3 13 13 9 9 2 16 1 0 9 9 0 9 0 13 2
13 3 7 9 1 9 9 0 13 9 13 7 0 2
23 15 7 13 1 9 1 9 9 0 2 15 13 15 9 1 13 7 1 15 1 15 13 2
20 7 15 13 9 9 9 13 15 15 1 9 13 2 9 3 13 1 9 0 2
64 3 16 9 15 4 13 16 13 7 13 7 15 9 15 13 0 9 0 9 2 7 9 9 2 7 10 15 9 2 3 3 13 15 16 13 13 15 9 0 2 7 15 9 2 16 1 9 10 3 13 16 13 3 9 2 7 3 9 0 2 16 13 4 2
68 7 3 7 1 13 13 3 9 1 9 0 9 1 9 2 16 1 9 0 9 0 1 9 2 13 9 1 9 2 7 15 3 13 1 0 13 2 16 3 9 1 0 13 2 7 15 9 9 0 13 9 9 1 9 1 15 2 16 3 15 13 13 9 1 9 7 9 2
53 1 0 13 2 16 16 16 9 13 1 9 2 3 13 16 9 9 13 12 2 3 9 9 7 9 9 2 7 12 3 2 16 13 9 2 3 3 9 15 3 13 13 12 2 7 12 3 2 3 9 3 0 2
19 7 16 9 3 13 13 15 9 2 15 9 13 1 9 2 15 13 0 2
27 7 3 15 13 2 16 13 9 0 9 2 7 15 13 15 9 15 13 9 2 7 3 13 16 9 13 2
16 7 15 3 13 13 2 16 9 9 3 13 13 2 7 13 2
7 15 3 13 13 1 9 2
16 3 2 16 9 0 13 15 1 15 9 9 2 3 9 0 2
11 7 9 0 0 13 1 9 1 9 9 2
29 1 0 13 2 16 9 0 0 15 9 13 9 1 9 2 1 9 0 13 1 9 1 9 0 2 16 13 4 2
12 7 3 3 13 0 1 9 0 7 15 9 2
18 16 7 9 0 15 13 1 9 9 2 3 9 15 13 1 9 9 2
16 15 13 13 15 3 13 9 7 9 7 9 13 1 9 13 2
23 1 15 7 9 9 16 9 13 2 3 9 13 2 3 16 13 9 2 7 9 13 13 2
52 7 16 9 13 9 0 13 2 16 13 4 2 3 0 7 9 7 13 13 2 16 1 10 9 2 16 13 13 9 7 9 7 9 2 15 3 1 0 13 13 2 16 1 2 8 12 1 9 2 13 4 2
26 1 0 3 13 2 16 9 9 13 13 3 1 15 15 13 9 3 13 2 7 3 1 9 15 13 2
30 7 0 15 9 13 2 16 1 9 3 13 9 0 9 2 13 13 3 1 9 2 7 1 9 2 3 1 9 9 2
26 7 13 0 15 15 13 2 16 9 1 9 9 9 1 9 13 2 16 9 3 13 1 13 9 9 2
56 3 1 3 9 3 1 9 9 7 9 7 9 2 3 13 1 9 9 2 7 1 9 2 16 13 2 3 13 4 9 2 16 13 15 15 13 1 9 9 2 3 9 7 9 1 9 13 2 7 9 7 9 1 9 13 2
29 1 0 3 13 2 16 9 0 15 13 1 0 9 9 2 16 13 2 15 13 2 16 16 15 9 13 7 9 2
36 1 0 13 2 16 1 15 9 13 15 9 2 3 15 0 9 2 7 15 9 2 3 9 13 2 15 13 9 15 9 2 15 13 9 9 2
14 7 15 12 13 9 13 2 16 3 1 9 9 13 2
11 3 9 1 9 13 15 13 2 12 13 2
36 9 3 13 9 7 0 2 15 9 1 9 9 13 2 0 13 2 16 13 7 9 7 9 7 9 2 7 15 15 15 1 9 9 13 13 2
31 7 15 3 13 13 2 16 12 9 3 13 13 16 12 9 2 16 12 9 16 12 9 2 7 12 9 3 16 12 9 2
17 16 1 9 0 3 0 13 9 0 2 7 3 9 1 9 15 2
13 7 9 15 1 9 13 2 13 13 16 9 0 2
29 15 9 13 15 9 13 9 9 0 2 16 1 10 9 9 7 9 9 13 13 2 16 0 13 2 13 9 9 2
8 7 3 15 9 9 9 13 2
9 7 1 2 9 0 9 13 13 2
25 15 9 13 9 9 10 13 2 1 13 2 8 12 2 12 2 3 16 15 13 2 7 16 15 2
21 1 0 13 2 16 0 1 15 13 9 2 13 9 9 2 16 9 13 9 9 2
14 15 0 13 9 9 2 16 9 7 9 2 3 9 2
11 7 9 0 1 9 0 1 15 9 13 2
20 1 0 9 13 2 16 9 15 13 1 9 1 15 16 9 13 2 12 13 2
25 3 16 13 1 13 9 1 9 7 1 9 15 13 9 13 2 16 15 15 13 1 9 1 9 2
22 7 13 9 9 1 9 13 0 2 3 1 9 0 9 1 9 2 7 1 9 9 2
33 13 7 1 9 15 13 1 9 0 13 2 15 1 9 10 9 13 15 15 13 1 10 9 2 0 13 16 15 9 13 9 13 2
61 3 3 15 9 13 1 10 9 2 16 9 15 13 0 9 1 9 13 2 0 1 9 13 13 9 13 1 9 1 9 2 15 9 10 9 13 2 7 9 0 1 9 1 9 0 2 15 9 9 13 1 9 0 15 13 2 15 13 3 13 2
36 9 7 15 0 1 9 13 2 3 13 9 0 1 9 9 2 7 15 1 9 13 2 16 1 9 15 13 1 9 9 2 16 13 9 0 2
36 9 7 15 3 13 9 2 16 9 7 9 2 0 1 9 13 2 15 13 1 9 0 2 7 0 1 9 1 9 0 9 2 16 13 4 2
45 1 0 3 13 2 16 9 1 9 9 3 15 13 16 9 0 2 7 16 9 0 2 15 9 13 2 16 9 9 13 2 9 1 9 13 2 3 16 9 2 7 16 9 0 2
25 7 1 9 3 13 9 0 2 15 9 13 9 0 13 2 7 3 15 15 13 2 15 13 15 2
22 1 15 7 15 4 13 13 3 2 16 9 0 2 13 1 9 13 0 9 1 9 2
56 1 0 9 13 2 16 16 1 9 0 2 1 15 12 9 13 7 15 13 2 1 15 16 9 12 13 9 15 2 13 13 13 1 15 2 3 1 9 2 15 9 13 7 9 13 2 13 13 9 9 1 0 9 1 15 2
15 7 9 9 7 9 9 13 1 9 0 2 15 13 9 2
11 7 0 1 9 15 13 1 9 7 9 2
28 16 1 9 9 0 9 13 9 9 3 13 15 2 7 9 13 9 9 3 13 15 13 9 1 9 9 0 2
26 1 9 7 9 0 15 13 1 15 9 10 15 1 15 9 13 0 15 9 2 16 9 7 9 9 2
31 7 3 1 9 0 16 9 12 13 9 15 1 15 16 9 12 13 7 15 13 2 9 9 13 15 13 1 9 9 0 2
12 7 3 1 9 9 0 13 0 9 15 9 2
25 7 16 9 7 9 7 9 13 1 15 9 7 9 2 3 3 1 9 9 0 9 9 0 13 2
15 16 9 0 13 2 13 9 9 9 2 1 15 9 13 2
22 16 9 0 13 9 9 2 7 1 15 13 9 10 15 1 15 3 13 13 9 9 2
35 3 1 9 9 7 9 9 2 16 1 13 13 2 15 13 16 9 12 9 7 9 15 2 13 16 1 9 9 0 9 9 13 9 9 2
17 1 15 3 9 13 9 1 9 15 13 9 2 7 9 1 9 2
13 16 9 15 13 9 2 13 9 1 9 9 0 2
9 7 9 13 0 1 9 9 0 2
22 7 1 15 9 15 9 13 13 3 0 9 9 0 2 1 16 9 0 13 9 0 2
50 16 9 15 13 3 1 9 0 2 3 13 1 9 0 2 7 16 9 13 1 15 9 7 9 9 3 13 13 2 7 0 2 3 3 13 1 9 0 9 2 16 3 13 1 9 13 1 9 9 2
22 3 2 9 9 7 9 9 15 13 1 9 16 9 12 9 7 9 15 1 9 0 2
15 3 2 9 15 13 3 7 0 2 3 13 3 1 9 2
11 15 9 9 13 1 15 0 1 9 9 2
24 0 7 13 16 10 0 1 9 13 0 2 3 0 2 16 3 13 9 3 13 0 15 9 2
18 1 0 9 13 2 16 9 9 13 9 9 15 15 13 1 9 13 2
12 7 9 9 13 0 9 9 15 15 13 9 2
7 16 9 13 2 9 13 2
27 7 16 13 13 9 16 0 13 2 13 7 2 16 0 3 13 2 3 13 13 9 1 9 15 7 15 2
12 7 3 3 13 3 9 12 9 7 9 15 2
11 1 0 9 13 2 16 0 13 9 9 2
24 15 3 9 13 15 13 3 7 0 1 9 1 0 2 7 1 9 1 9 0 2 16 9 2
10 7 3 15 9 3 0 1 9 13 2
27 15 7 9 13 15 3 13 3 7 0 2 7 3 7 3 2 16 9 15 13 1 0 2 16 9 0 2
17 7 15 9 7 13 0 1 9 2 7 13 7 13 16 13 4 2
52 15 7 9 0 9 15 13 2 16 3 13 3 7 0 1 9 1 0 2 15 16 15 9 10 0 0 13 7 1 15 13 1 9 0 2 7 3 13 3 7 0 1 9 1 10 9 2 16 13 1 9 2
15 7 3 15 9 3 13 0 1 9 2 16 7 9 0 2
16 7 3 16 13 2 13 13 7 13 2 16 9 0 0 13 2
30 7 15 9 13 9 2 16 15 9 13 1 10 13 2 15 16 10 13 3 13 9 9 16 15 9 2 16 7 9 2
68 7 3 16 1 9 13 9 9 0 1 9 2 7 1 15 9 9 15 9 2 7 1 15 9 0 9 2 15 13 9 1 9 2 7 1 15 9 9 2 3 9 9 13 1 9 2 7 1 15 9 13 9 9 2 7 9 0 9 2 15 13 3 9 0 1 13 9 2
17 7 9 15 13 1 9 2 16 9 1 9 2 16 9 13 9 2
16 1 0 13 2 16 9 13 1 9 0 3 1 9 15 13 2
21 7 13 2 16 9 9 3 13 9 1 9 2 16 9 13 9 1 9 15 13 2
16 3 3 13 9 9 13 15 9 1 0 2 15 0 3 13 2
12 0 13 9 9 2 16 13 9 9 9 13 2
25 7 0 9 0 2 16 9 9 13 9 1 15 13 2 15 13 9 0 9 13 2 15 9 13 2
24 1 9 7 9 9 1 9 13 1 15 9 0 13 2 15 9 9 13 1 9 9 1 15 2
11 7 1 0 3 13 9 2 7 0 9 2
31 7 9 9 13 1 15 9 2 16 13 1 9 9 2 16 1 2 8 12 2 8 12 2 8 12 2 8 12 2 13 2
20 7 3 1 15 15 13 0 9 2 16 13 15 9 2 15 1 15 13 13 2
35 1 0 3 13 2 16 16 1 9 7 9 3 13 9 1 9 1 9 2 7 1 9 9 1 9 2 3 3 7 1 9 7 0 9 2
28 1 0 9 13 2 16 16 9 9 15 13 13 1 9 2 3 13 9 2 3 7 9 15 9 13 9 9 2
21 7 3 15 15 13 15 9 2 13 15 9 2 7 15 15 9 1 15 9 13 2
12 7 0 9 3 13 15 9 9 1 9 15 2
24 7 0 3 16 13 15 9 13 15 9 10 9 13 2 16 1 9 13 2 7 1 9 13 2
23 1 0 13 2 16 0 9 1 15 9 13 9 9 1 15 9 2 16 9 13 7 13 2
11 7 3 3 13 16 13 1 15 9 9 2
23 3 16 1 9 7 9 1 15 9 13 12 9 2 3 3 1 9 13 2 7 9 9 2
28 1 0 9 13 2 16 1 9 1 15 13 9 7 9 2 9 13 1 9 9 0 2 7 9 1 9 9 2
39 7 3 1 9 13 1 15 9 13 16 9 2 7 9 9 16 9 2 0 15 9 3 1 9 13 13 1 9 13 2 7 3 1 9 2 1 9 9 2
24 1 0 13 2 16 1 9 9 3 13 1 9 9 2 7 1 9 0 1 9 2 3 9 2
22 7 16 9 9 3 13 1 12 9 2 3 9 9 3 13 9 1 12 15 9 9 2
4 12 1 9 2
21 16 9 9 13 1 10 9 7 1 10 9 2 1 1 15 9 9 13 7 9 2
10 7 9 15 9 0 13 3 15 9 2
44 1 0 3 13 2 16 9 15 9 3 13 1 9 9 7 9 2 15 13 1 9 15 2 16 13 16 3 15 9 13 9 7 9 2 1 15 13 12 9 2 7 15 9 2
13 7 1 15 9 9 9 7 9 9 9 3 13 2
34 1 0 13 2 16 9 15 13 9 15 9 2 16 13 2 7 3 15 9 1 10 9 13 9 2 3 13 1 15 2 1 9 0 2
12 16 15 9 13 12 9 1 9 1 9 9 2
7 3 15 9 13 15 9 2
9 13 16 15 9 3 13 15 9 2
23 1 3 9 9 13 1 9 2 7 3 1 9 2 13 16 9 13 1 15 15 9 13 2
14 7 9 15 9 3 13 13 7 1 0 7 1 9 2
7 3 9 3 13 15 9 2
13 7 15 13 3 1 9 9 13 9 16 15 9 2
28 3 1 3 13 15 9 0 13 1 10 1 15 9 2 16 0 9 13 2 13 16 15 9 3 13 15 9 2
26 3 2 1 9 3 13 9 16 1 9 9 2 16 13 9 9 9 13 9 13 2 16 1 13 4 2
7 3 3 13 15 9 9 2
6 9 7 13 9 9 2
13 3 1 15 13 9 0 9 2 13 16 13 9 2
16 13 16 9 15 9 13 13 1 9 0 2 7 3 1 0 2
28 7 9 9 3 13 1 9 9 16 1 9 0 2 16 1 13 2 15 13 9 10 2 7 2 15 13 15 2
9 3 13 13 9 15 9 9 0 2
15 3 2 1 9 9 13 13 9 9 2 15 13 1 9 2
31 3 2 1 15 9 13 3 9 1 9 15 9 2 13 15 9 9 13 1 9 9 8 2 7 15 13 0 15 9 9 2
10 3 13 16 1 15 13 9 15 9 2
15 7 1 2 15 15 13 9 9 2 1 10 13 16 13 2
8 3 9 15 9 13 9 0 2
17 3 1 9 9 13 1 9 2 13 16 9 15 9 13 13 9 2
11 13 16 13 9 3 13 13 9 15 9 2
23 16 1 9 15 9 13 9 1 9 2 16 13 1 9 2 2 15 3 13 1 9 13 2
6 3 3 13 13 9 2
20 7 1 9 15 9 3 13 9 1 9 0 2 7 3 1 9 7 1 9 2
6 3 9 13 13 0 2
18 13 13 1 0 9 2 16 15 13 16 15 9 13 1 9 15 9 2
21 9 7 9 3 13 1 9 13 2 1 1 0 15 13 13 2 16 1 9 9 2
21 7 3 9 15 9 15 9 13 13 1 9 2 15 13 9 15 9 2 16 13 2
19 7 1 15 13 2 16 0 13 2 16 13 9 13 2 16 7 15 9 2
17 7 3 9 9 2 16 1 10 13 13 2 13 1 0 9 13 2
17 7 0 9 9 2 15 13 9 15 9 2 15 13 1 9 9 2
10 7 9 15 9 3 13 1 9 13 2
21 1 0 13 2 16 15 9 15 13 1 9 9 2 3 9 0 2 1 10 13 2
9 7 1 9 9 13 9 9 13 2
35 1 0 9 13 2 16 9 15 9 13 9 0 2 16 13 1 9 9 2 7 1 9 9 9 2 15 0 9 0 13 1 9 15 9 2
16 7 3 1 15 9 3 13 13 9 0 9 16 1 13 9 2
24 1 0 13 2 16 1 15 9 15 13 1 9 2 3 2 1 15 0 9 2 3 13 9 2
41 1 0 13 2 16 9 15 0 9 2 15 1 9 15 13 9 2 3 13 9 15 9 2 7 13 15 9 1 9 2 16 9 9 13 1 9 15 1 15 9 2
14 1 0 9 13 2 16 13 9 13 13 9 15 9 2
25 1 0 3 13 2 16 9 15 9 13 13 1 9 9 2 3 7 9 9 1 9 1 9 13 2
26 1 0 13 2 16 1 9 13 13 9 0 2 7 15 3 13 1 9 2 16 13 9 1 9 13 2
14 9 15 9 15 9 13 9 2 15 13 9 15 9 2
14 7 1 13 16 15 13 13 9 15 3 13 9 9 2
21 7 9 15 9 3 13 9 2 15 3 13 1 9 7 9 2 16 1 9 13 2
13 15 13 1 15 16 1 9 9 9 15 9 13 2
19 3 0 1 0 9 13 2 16 1 15 9 13 2 15 3 13 1 9 2
10 13 16 9 15 9 9 1 9 13 2
7 16 9 9 13 1 9 2
20 3 1 9 15 9 13 13 9 1 9 0 1 9 9 2 16 1 15 9 2
18 3 2 1 9 9 3 13 13 9 16 1 15 15 13 1 9 9 2
12 3 3 13 1 15 13 9 1 9 15 9 2
11 7 1 9 15 9 3 13 9 1 9 2
34 3 7 1 9 15 9 13 1 15 13 9 2 16 13 1 13 2 13 9 2 16 0 9 10 13 2 1 15 15 9 9 3 13 2
21 7 3 1 9 9 13 9 9 1 9 15 13 2 7 13 9 9 1 0 9 2
22 3 15 9 9 13 13 16 9 9 13 1 9 9 2 16 13 2 13 15 7 15 2
22 1 0 13 2 16 9 0 13 1 9 1 15 1 16 1 15 13 13 1 9 10 2
15 7 3 1 15 15 16 9 0 13 2 1 9 9 13 2
24 7 15 13 1 9 2 16 3 1 0 1 15 9 13 9 1 0 9 1 9 7 13 9 2
23 13 13 2 16 2 16 13 4 2 15 13 9 15 13 2 7 9 1 0 13 1 9 2
25 7 16 0 9 9 13 13 9 7 9 0 2 3 1 15 9 9 1 9 9 13 9 0 13 2
20 1 0 13 2 16 3 0 13 13 0 9 2 7 3 0 9 1 9 9 2
45 7 3 15 13 2 16 3 13 1 9 13 9 7 15 9 13 2 16 9 13 7 9 13 2 7 3 1 0 9 2 15 13 9 9 2 7 3 1 0 2 15 13 9 9 2
33 1 0 13 2 16 1 9 9 13 9 0 2 16 16 1 15 3 13 1 15 2 13 3 1 15 3 1 9 9 2 15 13 2
14 10 3 9 0 9 13 15 9 15 13 1 9 9 2
26 1 0 3 13 2 16 9 15 9 0 13 2 13 9 15 9 2 3 7 9 9 15 13 15 0 2
15 3 2 10 9 13 9 2 13 15 1 9 7 9 10 2
38 1 0 13 2 16 16 9 9 7 9 9 3 13 1 9 0 2 7 1 9 2 3 9 0 7 9 13 9 0 13 9 15 2 15 13 9 9 2
14 3 2 3 13 13 9 7 13 9 2 3 13 9 2
27 7 1 0 9 13 13 9 2 16 13 9 0 1 13 2 7 13 9 2 16 13 9 1 0 9 13 2
25 3 2 0 13 1 9 9 9 2 15 13 9 2 16 9 2 16 9 16 9 1 9 9 0 2
36 16 7 1 9 13 1 9 9 13 9 9 15 9 2 1 15 9 0 13 13 9 2 3 1 15 15 9 13 2 9 13 13 9 7 9 2
27 1 0 13 2 16 16 9 0 9 1 9 13 2 3 9 9 9 1 15 13 2 16 13 1 12 8 2
12 3 2 9 9 3 13 1 9 16 1 9 2
17 7 1 9 9 13 9 2 9 9 2 16 13 1 12 1 8 2
26 7 1 15 15 13 1 9 2 15 13 9 9 2 13 9 2 16 1 9 7 9 7 9 7 15 2
25 7 1 0 9 3 13 13 9 16 9 2 16 9 13 1 9 9 0 2 7 9 0 1 9 2
20 1 0 13 2 16 9 13 9 9 9 15 13 1 15 9 2 16 7 9 2
30 9 9 13 9 3 13 2 7 3 13 13 2 16 13 15 0 15 9 9 3 13 2 7 3 1 9 9 4 13 2
27 1 0 13 2 16 9 3 13 1 9 2 1 15 15 13 9 2 16 1 9 2 1 15 13 1 9 2
23 9 7 13 1 9 15 15 13 2 16 15 9 9 13 9 2 7 16 9 10 13 9 2
44 16 3 0 9 13 9 1 15 2 3 9 15 13 9 9 2 7 9 1 15 2 3 9 0 2 3 9 0 13 9 1 15 2 9 7 9 2 9 1 15 2 9 0 2
42 3 1 1 0 9 13 10 15 13 1 9 9 2 16 13 9 15 13 9 9 2 7 13 9 2 3 9 9 0 1 9 2 13 3 16 0 9 13 9 16 0 2
19 7 15 9 0 9 1 12 1 9 13 2 13 9 9 16 9 9 13 2
25 1 0 13 2 16 9 3 13 1 9 0 16 13 1 9 15 13 2 7 3 16 9 1 9 2
52 7 13 2 3 1 15 2 7 13 0 9 0 9 1 9 9 0 9 2 3 9 2 7 9 9 15 13 9 1 9 0 2 16 13 1 9 9 1 9 9 2 7 3 1 10 15 1 9 9 7 9 2
43 3 16 10 9 9 9 13 15 9 1 15 3 13 16 9 9 0 13 9 2 7 13 9 13 2 3 1 0 9 2 1 15 15 9 9 13 2 3 13 13 9 9 2
11 9 7 0 13 13 9 1 9 10 9 2
28 3 3 15 9 2 1 15 13 9 9 1 9 2 13 0 9 9 15 13 15 9 2 16 9 1 9 13 2
27 3 7 15 9 15 9 13 2 3 13 9 0 7 1 15 15 9 1 15 13 9 2 7 9 15 9 2
54 1 0 13 2 16 16 9 9 13 9 13 2 16 1 13 4 2 3 1 15 16 13 2 7 1 15 16 13 2 3 15 9 2 15 13 2 13 9 0 1 13 2 3 1 15 16 13 2 7 1 15 16 13 2
17 3 7 13 15 9 15 2 7 15 1 13 4 13 1 9 9 2
26 1 0 13 2 16 15 13 13 1 0 15 7 1 9 9 2 3 16 1 0 9 9 9 10 13 2
16 3 2 15 9 13 9 1 10 9 2 7 0 15 9 9 2
15 7 9 13 1 9 16 9 1 9 2 7 9 1 9 2
20 7 9 13 2 15 13 9 0 9 0 2 16 9 15 2 3 13 15 13 2
25 7 9 9 3 13 1 3 13 1 9 2 1 13 9 0 2 7 0 9 0 1 15 13 9 2
8 3 9 9 3 13 15 9 2
22 0 2 16 9 15 13 9 15 2 3 13 9 7 9 16 9 2 7 13 9 3 2
9 3 7 9 3 13 1 3 9 2
46 3 2 9 9 0 13 1 9 16 9 9 1 9 2 16 0 15 13 1 9 9 1 9 2 7 0 1 9 2 16 13 1 9 1 12 8 2 7 9 15 13 1 12 1 9 2
26 7 16 9 13 0 2 7 15 13 0 2 16 9 13 1 15 16 9 1 9 2 16 13 12 8 2
26 15 0 13 2 16 9 3 13 9 0 16 9 9 2 7 0 0 2 16 9 0 2 7 9 9 2
19 1 0 13 2 16 15 15 13 1 9 1 9 2 13 1 9 1 9 2
45 13 7 2 16 9 13 1 12 8 2 7 1 8 1 9 9 2 1 9 0 7 0 1 9 0 13 9 3 13 2 1 15 13 9 9 2 16 0 9 1 0 9 13 13 2
14 3 7 1 9 9 0 1 9 3 9 15 13 15 2
33 7 3 9 1 15 9 13 2 15 9 13 2 13 0 9 1 15 15 1 15 13 4 2 16 15 9 15 9 1 15 9 13 2
66 1 0 13 2 16 16 9 0 3 13 9 0 9 2 7 9 0 15 2 7 9 1 15 9 13 0 15 9 2 3 9 9 2 15 13 9 13 1 9 0 1 0 13 2 3 13 0 9 9 13 2 7 13 9 0 2 7 9 1 15 9 13 0 1 9 2
39 9 7 0 1 15 9 9 3 13 15 9 0 16 9 0 2 16 16 13 15 9 0 0 15 2 13 15 9 0 2 7 3 1 15 13 1 9 9 2
26 7 3 9 9 1 9 13 16 9 9 0 1 10 9 3 1 15 16 13 1 9 9 1 10 9 2
17 3 1 9 0 13 2 15 9 9 0 0 13 3 1 3 13 2
10 9 7 0 9 3 13 9 1 9 2
64 7 13 2 16 15 0 7 0 9 3 13 1 15 0 2 16 1 9 9 13 13 2 16 13 1 9 0 2 15 9 2 15 15 1 9 13 2 3 1 9 13 2 7 1 9 15 9 9 1 9 13 2 1 3 13 15 9 9 7 15 9 1 9 2
44 7 3 15 9 13 4 1 9 0 9 2 16 3 13 15 9 13 1 9 13 2 16 13 1 15 9 13 2 15 9 3 13 2 9 3 13 2 9 7 1 15 9 13 2
16 1 0 13 2 16 1 9 7 1 15 9 15 13 0 9 2
15 15 3 13 2 16 15 1 9 13 9 15 7 9 9 2
19 9 9 1 16 13 9 2 9 7 15 1 16 1 15 15 9 9 13 2
41 15 9 13 9 2 15 0 13 2 16 9 15 3 13 9 9 3 2 7 9 15 15 1 9 9 2 7 13 15 13 1 9 9 7 9 2 13 1 15 15 2
10 7 15 9 15 2 9 7 9 13 2
21 0 7 9 13 9 9 0 2 13 7 16 9 13 15 15 9 13 9 7 9 2
51 0 3 7 13 9 9 2 16 13 9 1 15 9 2 16 9 15 3 13 1 9 9 2 7 13 15 2 15 16 9 3 13 1 15 9 15 13 9 7 9 2 16 13 12 8 2 16 13 9 9 2
13 3 13 15 9 9 2 3 13 15 9 9 9 2
37 16 7 13 16 15 9 1 9 1 9 13 0 7 0 2 15 1 15 9 13 2 16 9 13 1 9 2 15 13 9 0 2 16 1 9 0 2
35 1 9 7 2 15 13 9 0 2 13 15 9 2 16 1 9 0 2 15 0 9 13 1 13 15 15 13 2 16 1 12 1 9 13 2
21 7 1 9 0 13 1 16 13 9 2 15 9 15 13 2 7 13 2 9 13 2
12 7 9 9 2 3 9 2 13 1 9 9 2
30 7 3 3 13 1 9 15 13 1 9 2 16 9 3 13 15 9 1 9 2 7 1 9 2 1 15 13 9 15 2
12 3 7 9 13 0 2 16 3 1 9 0 2
35 13 13 1 0 9 2 16 2 16 13 1 12 1 9 2 9 13 15 1 9 3 0 1 9 9 7 9 2 7 3 1 9 9 0 2
29 1 0 3 13 2 16 9 0 13 13 1 9 1 9 2 7 1 9 9 1 9 2 7 1 9 9 1 9 2
48 16 15 13 15 13 15 9 13 2 1 15 13 1 9 9 2 16 9 2 7 15 12 9 2 15 9 13 1 9 2 15 1 15 13 2 7 3 13 15 9 13 2 16 7 15 9 9 2
20 15 0 9 13 1 9 13 1 9 1 9 2 3 1 9 9 1 9 9 2
24 7 15 9 3 13 2 16 1 9 9 9 0 1 10 9 13 2 16 12 1 15 3 13 2
17 7 3 3 13 15 9 15 13 1 15 9 13 1 9 1 9 2
56 7 1 15 16 9 1 9 0 13 9 13 2 9 15 13 1 9 0 2 16 9 13 2 3 7 9 13 1 9 9 0 2 16 7 15 9 2 16 3 13 1 15 9 16 15 9 2 7 9 13 3 13 9 16 13 2
26 7 15 13 15 13 9 0 9 2 16 0 9 13 15 13 0 9 9 2 1 15 13 0 9 9 2
24 13 3 3 1 15 16 13 15 15 13 1 9 9 7 9 2 15 9 1 9 0 9 13 2
23 1 0 3 13 2 16 9 0 3 13 15 15 13 2 1 10 9 2 7 1 10 9 2
29 3 16 15 9 15 3 13 9 9 0 13 1 9 1 9 9 0 2 3 13 16 13 9 9 2 7 9 9 2
50 3 3 15 9 13 9 1 12 1 9 2 1 13 0 9 2 7 1 13 16 15 9 13 13 7 1 9 3 1 15 15 13 9 7 9 1 15 2 7 1 9 3 1 15 15 13 9 7 9 2
19 13 7 16 9 9 3 13 9 1 9 0 2 16 16 13 1 15 9 2
19 1 0 13 2 16 1 9 0 7 0 9 0 13 13 1 9 9 0 2
11 7 9 0 7 13 13 9 1 9 0 2
21 7 15 9 3 13 16 1 9 9 2 15 13 13 9 2 16 7 10 15 9 2
23 3 1 10 9 13 15 9 0 2 1 10 13 13 1 9 15 9 9 2 16 13 9 2
24 1 0 13 2 16 9 3 9 3 0 13 9 9 2 7 3 9 9 2 16 1 13 13 2
32 3 2 10 15 13 1 9 1 9 15 2 13 0 1 15 2 16 1 15 15 13 0 1 15 2 16 13 1 12 1 8 2
12 7 9 0 1 9 13 1 9 1 15 9 2
14 15 13 1 9 2 12 15 13 1 9 1 9 15 2
16 9 3 1 16 13 1 12 9 2 3 13 9 1 15 9 2
8 3 13 1 9 1 15 9 2
29 7 3 2 1 9 15 13 0 9 9 2 1 9 7 9 15 13 2 13 3 0 16 2 9 13 2 9 13 2
31 0 13 7 16 15 13 1 0 16 16 13 9 9 0 1 9 0 2 13 1 9 15 13 1 9 2 1 15 3 13 2
17 9 3 13 9 9 2 13 15 1 12 2 1 16 13 1 15 2
28 7 16 1 9 0 3 9 13 9 1 9 2 3 9 13 13 15 2 16 13 3 1 15 9 9 0 9 2
20 7 3 1 9 15 13 15 9 1 9 15 15 3 13 2 3 1 9 9 2
14 16 3 9 3 13 9 2 3 9 0 3 13 0 2
19 13 3 1 15 16 9 1 9 13 2 16 13 15 9 1 15 9 0 2
30 7 16 1 9 0 9 13 9 3 2 3 13 4 9 9 1 15 9 15 0 13 9 2 7 13 1 15 0 9 2
42 7 3 15 13 2 16 13 9 2 1 15 9 0 0 13 2 13 1 9 9 13 2 15 13 9 9 2 1 15 2 9 15 9 0 0 13 2 3 3 9 13 2
35 0 7 9 15 9 9 13 2 13 1 13 9 0 2 16 13 15 16 9 9 2 7 3 13 15 1 15 9 9 2 16 9 13 9 2
24 0 2 16 9 15 9 9 13 2 13 1 9 13 2 13 15 9 9 3 9 13 10 9 2
21 15 3 15 1 9 9 13 1 9 2 13 3 1 9 9 2 16 1 9 9 2
21 13 7 15 9 13 0 1 9 7 9 7 0 9 2 15 10 1 9 9 13 2
17 7 3 13 9 7 9 2 7 0 9 1 0 7 0 7 3 2
12 0 3 7 9 9 13 16 1 9 9 13 2
13 9 7 13 9 3 0 16 9 2 7 16 9 2
44 3 16 1 9 9 13 15 0 2 16 13 9 9 2 13 9 0 2 3 1 9 9 13 15 16 13 9 2 16 3 13 13 7 0 1 13 9 1 10 9 7 9 9 2
34 3 7 0 13 9 13 1 15 3 2 7 3 1 15 2 16 13 1 9 0 0 7 0 2 16 1 15 9 15 13 1 9 15 2
15 13 3 9 9 13 2 15 13 9 1 15 0 7 0 2
34 1 9 7 9 3 13 15 9 7 9 13 1 0 9 2 7 0 9 2 16 9 3 13 9 16 1 16 1 9 13 13 9 0 2
21 13 3 15 9 13 1 15 15 1 9 0 0 2 16 9 13 1 9 1 9 2
57 15 9 1 9 0 1 9 15 13 1 9 2 16 13 1 10 9 0 2 1 15 3 13 16 1 9 13 9 0 2 15 1 0 0 13 2 16 9 15 13 1 9 13 1 9 13 0 1 15 2 7 1 9 9 13 0 2
11 7 9 9 1 9 0 13 13 9 15 2
23 9 16 1 9 13 2 13 1 9 16 1 15 7 9 13 12 2 16 1 9 7 9 2
9 7 9 3 13 9 15 9 0 2
13 3 2 0 13 13 9 1 9 16 9 1 0 2
14 7 9 9 0 7 0 3 13 16 9 13 9 9 2
23 3 13 16 15 9 13 13 16 9 2 9 7 16 9 13 2 16 9 13 9 9 9 2
22 16 7 9 15 1 15 15 16 1 9 10 9 13 2 13 9 9 15 9 0 13 2
45 1 0 13 2 16 9 9 0 3 13 13 9 9 16 9 0 15 2 16 9 9 15 13 2 7 13 9 15 16 13 15 1 0 9 2 16 9 13 9 9 13 15 1 13 2
28 3 13 0 9 13 16 13 15 0 2 16 9 13 9 1 9 13 9 2 7 9 13 9 13 1 9 9 2
13 12 9 16 9 9 2 16 1 15 13 12 0 2
72 16 7 9 1 9 3 13 15 9 2 15 13 9 7 13 9 2 13 3 15 15 0 9 1 9 15 1 9 9 15 2 1 15 13 3 1 9 2 15 9 15 0 1 9 13 13 2 1 16 3 13 1 0 9 2 15 9 0 1 9 13 2 3 9 2 15 9 9 9 13 13 2
51 0 7 7 0 13 15 1 15 15 13 15 15 13 9 9 2 15 2 16 8 12 2 8 12 2 8 12 2 8 12 2 1 12 2 13 4 2 3 13 13 2 3 7 3 13 2 1 0 9 9 2
52 16 3 13 15 9 9 2 15 13 15 7 15 2 13 15 1 9 2 15 15 15 13 2 3 13 9 9 1 15 13 2 16 15 3 13 13 1 15 9 9 2 1 15 13 0 9 2 1 15 9 13 2
42 16 7 9 1 15 9 13 2 15 13 15 7 15 2 15 7 9 15 2 7 15 15 13 1 9 13 15 1 9 13 2 15 9 3 0 0 2 7 3 13 13 2
24 1 0 9 13 2 16 15 15 13 0 1 15 2 13 13 1 15 2 16 1 9 9 13 2
10 13 3 13 2 1 15 9 0 13 2
22 3 2 16 1 13 8 13 2 0 1 9 9 13 2 1 15 0 1 10 13 13 2
26 7 15 1 9 7 9 9 13 16 15 0 9 13 15 13 2 16 9 9 13 13 0 16 9 0 2
14 1 0 13 2 16 9 13 7 9 9 13 0 13 2
40 7 16 9 13 1 9 9 2 9 9 0 3 13 9 9 16 9 9 13 2 16 3 9 13 1 15 13 15 9 9 2 16 9 0 2 15 9 13 0 2
19 1 0 13 2 16 1 9 9 4 9 0 9 13 2 15 1 3 13 2
14 3 2 9 9 13 0 9 1 15 13 13 0 9 2
13 7 12 15 13 0 9 0 2 3 9 7 9 2
21 1 12 0 2 3 9 7 9 2 3 13 9 0 15 2 7 13 1 9 9 2
31 7 3 12 9 2 3 9 2 9 7 9 2 9 13 2 16 9 13 15 9 0 15 3 13 2 16 3 3 9 13 2
52 13 3 7 9 2 1 15 13 3 13 16 9 9 13 1 9 1 9 9 2 1 7 9 13 0 2 7 9 1 3 2 7 3 9 2 16 1 15 9 3 13 9 0 1 9 10 9 2 12 9 13 2
53 7 3 15 13 2 16 10 9 13 1 9 2 7 9 0 7 0 1 15 13 2 16 3 13 16 1 9 13 9 13 1 9 10 0 1 15 16 0 9 13 2 1 13 1 0 13 2 7 0 15 0 13 2
55 7 15 3 13 0 2 1 9 0 9 13 9 9 0 2 16 9 0 13 9 13 13 13 2 16 1 9 0 1 9 2 16 1 9 13 13 16 1 9 10 9 9 13 2 15 1 9 9 13 2 16 9 9 13 2
31 13 3 2 16 9 16 13 0 16 13 9 9 2 0 9 7 9 2 0 3 13 0 2 16 15 9 9 9 9 13 2
14 1 0 3 9 13 1 15 9 0 1 9 13 13 2
10 1 0 13 16 0 13 1 9 9 2
21 7 16 13 0 1 9 9 13 1 9 13 2 3 3 13 13 9 13 1 9 2
10 1 0 13 16 0 1 9 9 13 2
10 1 0 16 1 9 9 0 2 3 2
12 7 1 1 9 0 13 15 13 2 13 8 2
9 12 3 0 1 9 9 4 13 2
8 3 0 1 9 9 4 13 2
10 13 16 0 1 9 9 3 4 13 2
6 3 1 9 9 13 2
6 3 1 9 9 13 2
7 3 3 13 1 9 0 2
10 3 0 1 9 13 1 9 9 0 2
12 13 16 0 1 9 3 13 1 9 9 0 2
7 7 13 4 1 9 0 2
11 3 1 9 9 13 2 3 1 9 0 2
9 3 13 16 3 13 1 9 0 2
15 3 2 1 15 9 9 1 9 13 15 1 10 13 13 2
30 7 0 1 9 9 0 3 13 13 1 10 2 0 7 0 2 16 9 3 13 3 13 13 13 1 13 9 9 0 2
7 3 3 13 1 9 0 2
10 3 1 9 3 13 10 1 9 0 2
12 3 2 1 15 9 0 13 1 15 13 4 2
16 1 15 9 0 13 4 2 0 13 2 16 13 1 0 13 2
7 7 13 4 1 9 9 2
6 3 1 9 0 13 2
9 3 0 0 9 1 9 0 13 2
19 7 1 0 9 2 1 15 0 13 1 15 16 13 2 1 9 9 13 2
17 3 1 0 9 1 15 13 1 15 16 13 2 13 1 9 0 2
21 16 3 1 0 9 1 15 13 16 1 15 13 1 9 2 1 9 10 9 13 2
7 7 3 1 9 0 13 2
11 7 3 1 9 0 0 1 9 13 13 2
21 1 0 13 2 16 9 3 13 1 9 0 2 1 15 13 4 2 7 3 13 2
28 13 13 1 0 9 2 16 2 16 1 13 4 2 0 1 13 13 2 1 9 0 13 1 9 15 9 13 2
42 1 0 13 2 16 16 0 1 15 16 0 13 4 2 0 9 13 2 3 3 13 1 9 9 2 1 15 0 13 4 2 7 1 9 0 2 1 15 1 9 13 2
36 1 0 3 13 2 16 9 13 3 13 9 9 2 7 13 3 1 15 2 13 1 9 9 2 7 1 9 9 2 15 1 9 0 3 13 2
12 3 2 9 7 9 13 0 9 16 15 9 2
19 15 13 3 13 2 16 1 9 15 1 15 13 2 3 13 15 9 13 2
22 7 15 1 9 9 2 3 1 9 9 2 3 9 0 2 15 1 9 9 13 0 2
36 9 0 0 7 9 7 0 7 10 9 13 13 7 1 15 7 1 9 2 7 1 9 9 15 9 13 2 7 1 9 9 15 9 3 13 2
48 1 7 9 0 13 1 15 9 9 0 9 2 9 7 0 9 2 16 13 9 2 13 0 9 2 13 16 7 1 15 9 0 9 9 13 2 7 1 15 1 15 9 1 9 0 9 13 2
34 1 0 13 2 16 16 9 1 9 7 9 13 2 3 9 0 13 1 9 2 3 1 9 2 16 9 15 9 13 9 9 15 0 2
34 16 3 9 13 1 9 16 1 9 2 7 9 1 9 2 16 13 1 12 1 9 2 3 7 9 9 13 1 9 9 16 1 9 2
14 1 0 13 2 16 9 13 1 9 3 9 0 9 2
21 7 15 3 13 10 9 15 13 9 2 15 13 9 0 9 2 13 9 1 9 2
62 15 0 15 13 9 2 15 13 9 0 9 2 3 13 9 1 9 2 7 1 15 13 9 15 9 15 13 13 2 7 12 0 10 2 13 9 2 15 13 9 9 2 13 0 2 7 13 1 9 9 2 7 0 1 15 9 9 2 15 13 4 2
25 1 0 13 2 16 1 9 12 13 13 2 3 9 9 2 7 9 15 2 1 15 9 13 9 2
9 7 1 9 10 9 13 15 9 2
22 7 3 15 9 3 13 15 9 2 7 15 9 9 2 7 9 2 16 1 13 4 2
22 7 15 9 13 15 15 13 9 1 9 2 7 13 9 2 7 9 2 7 15 3 2
12 3 7 15 15 13 1 9 16 9 1 9 2
18 15 7 3 13 13 15 0 9 2 16 9 7 13 13 13 12 9 2
21 13 3 16 9 15 13 9 10 13 9 2 13 15 9 13 1 9 1 9 10 2
40 15 0 13 2 16 16 9 9 3 13 1 0 9 2 16 1 16 13 9 13 2 3 9 13 9 3 13 1 15 7 15 2 16 1 16 13 0 9 0 2
24 7 3 16 9 13 9 13 1 9 9 2 13 9 13 2 15 13 12 7 15 1 0 13 2
22 12 3 9 13 13 9 2 16 13 9 1 15 9 9 2 7 3 1 15 9 9 2
42 1 15 7 16 9 13 9 2 13 16 13 1 15 9 9 1 9 10 9 2 16 3 1 15 9 13 2 16 13 15 9 9 9 1 9 2 7 1 9 1 9 2
13 16 3 13 1 9 9 0 2 3 13 13 9 2
29 3 3 9 13 1 9 7 9 2 13 9 9 1 9 13 15 13 3 2 7 1 9 1 15 13 1 9 0 2
79 1 3 1 15 9 13 0 15 9 2 15 9 13 7 13 2 9 15 15 9 13 1 13 9 13 2 3 13 9 15 9 13 1 9 13 2 16 13 0 9 2 7 15 9 13 1 9 13 1 9 10 2 16 13 0 2 7 13 15 9 13 2 15 13 9 10 16 9 2 16 15 13 15 13 2 7 15 13 2
37 7 15 13 1 15 9 13 2 3 15 9 13 15 13 1 9 9 1 9 2 16 15 15 9 13 9 10 2 3 13 1 15 13 1 9 0 2
49 15 3 3 13 13 16 0 9 13 0 9 9 10 2 7 16 1 15 7 9 10 13 12 0 2 16 1 0 1 9 7 9 0 2 7 16 9 9 0 1 9 10 13 16 9 9 1 9 2
55 16 3 15 12 2 15 12 13 9 15 2 13 1 15 0 2 9 12 12 1 15 2 3 3 9 1 0 9 2 13 16 9 9 1 9 2 16 9 7 9 13 1 0 2 15 9 15 13 1 9 16 9 1 9 2
32 7 3 1 1 9 13 9 0 2 7 15 9 0 13 2 16 3 1 15 9 2 9 0 15 13 1 9 16 9 1 9 2
34 16 3 1 9 0 15 15 13 9 2 7 9 2 13 12 9 0 2 3 1 9 15 9 13 2 7 15 9 2 13 12 1 13 2
33 1 9 7 0 9 1 15 13 3 13 13 9 15 9 2 16 15 9 13 9 9 15 2 16 3 13 13 16 9 13 9 15 2
31 7 16 15 9 1 15 13 13 9 3 2 15 13 15 13 9 15 9 2 7 13 15 13 15 9 2 16 13 1 9 2
18 1 9 7 13 13 15 9 1 9 3 9 2 7 9 0 3 9 2
32 3 16 13 15 9 1 15 13 15 3 13 15 1 15 1 15 15 13 0 1 15 2 15 9 1 15 13 13 9 15 13 2
17 15 9 13 2 16 13 9 0 13 1 9 2 7 10 9 9 2
17 7 3 2 1 9 0 13 9 0 2 13 13 9 15 9 13 2
19 1 13 7 2 15 15 13 13 9 15 13 2 16 1 9 9 13 9 2
28 1 0 13 2 16 9 3 13 1 9 15 9 1 9 13 1 15 9 13 2 15 9 10 13 1 15 13 2
29 7 2 16 13 9 2 9 10 9 9 10 13 2 16 15 9 9 10 13 2 15 9 3 13 1 9 0 9 2
20 7 1 0 15 15 1 9 15 13 9 10 2 13 2 7 13 15 3 13 2
32 1 0 13 2 16 9 9 16 13 10 9 15 3 9 13 2 3 3 13 15 9 0 2 15 13 3 9 9 10 1 0 2
14 7 1 15 9 13 2 16 9 13 13 13 1 9 2
23 1 0 13 2 16 1 9 15 9 1 9 13 2 15 0 9 13 3 9 9 15 13 2
28 7 3 15 9 13 16 9 10 13 9 2 13 15 9 0 2 7 16 15 9 13 1 15 3 9 7 9 2
18 7 0 0 13 13 1 9 9 13 2 16 9 3 3 13 1 9 2
21 7 15 13 9 0 15 13 15 9 1 0 9 2 16 1 9 9 1 13 9 2
15 7 3 3 9 0 3 13 1 9 2 3 13 9 9 2
14 7 3 13 16 9 1 9 13 15 9 13 9 9 2
14 3 2 9 9 13 1 9 9 2 15 13 9 9 2
14 7 9 2 15 13 9 9 2 13 15 15 13 13 2
19 1 0 13 2 16 9 3 13 9 3 2 15 13 9 9 2 7 9 2
21 7 3 9 13 13 3 0 1 9 2 15 13 9 9 2 7 3 1 9 9 2
28 7 9 15 3 13 1 15 0 2 3 13 15 9 1 9 9 2 16 3 13 9 16 16 13 9 15 9 2
8 7 3 9 9 13 9 9 2
28 7 9 15 13 1 15 0 2 13 15 9 16 13 9 15 0 2 7 15 9 2 1 16 13 9 15 9 2
14 7 15 9 13 1 9 15 0 13 16 13 15 9 2
20 13 13 2 16 1 9 9 13 9 15 13 2 13 1 9 15 13 9 9 2
15 15 7 1 9 0 16 1 15 9 2 16 0 13 4 2
26 1 15 3 9 13 9 9 1 9 1 9 15 15 13 4 1 9 1 9 2 16 1 9 1 0 2
14 1 9 7 0 2 1 16 9 13 9 3 7 0 2
15 9 7 0 13 9 15 13 2 1 15 16 13 9 13 2
17 3 1 9 13 9 13 9 15 13 9 10 9 0 16 9 0 2
21 7 1 13 9 9 1 9 2 15 15 9 13 9 2 3 1 9 9 1 9 2
44 1 0 13 2 16 16 1 9 12 0 3 13 13 9 9 15 15 13 2 16 1 15 2 16 15 1 9 10 9 13 2 3 9 12 9 13 9 15 13 2 16 9 15 2
22 3 1 1 15 0 9 9 0 13 3 9 9 10 2 13 16 0 13 9 10 13 2
21 3 2 9 13 1 12 1 9 2 16 16 9 13 13 9 9 0 2 13 10 2
34 3 13 2 16 1 9 0 3 9 7 9 13 1 0 9 2 16 9 15 13 1 9 13 2 9 0 1 9 0 13 1 9 15 2
22 7 1 9 0 13 15 1 9 15 9 2 16 9 13 1 9 9 2 7 1 0 2
23 1 0 13 2 16 9 13 13 9 13 9 0 2 16 3 9 9 13 13 9 9 0 2
24 7 3 16 9 13 13 9 9 0 2 13 16 9 0 13 10 1 15 15 13 9 9 13 2
12 0 7 9 3 13 9 15 9 9 10 13 2
25 13 13 2 16 1 15 16 9 9 1 9 13 2 13 16 9 0 13 9 10 3 16 9 0 2
16 9 7 3 13 0 16 16 0 13 9 15 13 0 15 9 2
36 0 3 9 1 9 1 15 9 13 1 0 7 9 15 2 3 16 16 12 13 0 2 7 15 2 16 0 1 0 9 1 9 13 15 9 2
14 9 7 15 13 0 9 2 10 9 7 9 0 13 2
15 7 3 9 7 9 9 3 15 13 16 1 10 9 9 2
19 1 7 0 9 13 9 13 13 1 9 9 1 9 13 15 13 7 13 2
39 9 3 9 10 13 1 9 0 15 1 9 13 13 13 1 9 2 15 16 9 15 9 15 13 1 9 10 16 0 1 9 2 16 13 1 12 1 9 2
23 7 3 13 16 1 10 15 15 9 10 13 2 0 13 1 9 0 2 16 3 9 13 2
26 7 16 9 13 2 15 13 1 15 0 0 2 13 9 9 0 2 3 9 10 13 0 1 9 15 2
25 9 7 0 9 0 2 16 3 13 13 1 9 0 2 13 3 13 1 9 13 15 13 10 9 2
20 16 3 0 9 13 15 9 0 2 3 3 13 0 15 9 2 16 9 0 2
21 15 3 0 13 16 1 9 13 9 0 1 15 16 13 0 0 9 16 9 0 2
14 0 1 9 9 0 9 1 9 15 9 13 0 13 2
11 13 7 1 9 0 0 13 9 9 0 2
17 7 3 9 15 1 15 9 13 9 0 0 2 13 13 9 13 2
43 9 3 9 1 9 9 1 10 9 0 2 7 3 0 2 3 13 1 15 0 16 16 13 10 15 13 1 9 13 2 1 15 0 9 9 15 13 2 16 1 13 13 2
27 9 7 1 9 10 13 3 13 7 1 15 9 1 9 13 2 7 1 15 9 13 2 16 1 13 13 2
49 1 13 3 13 16 15 9 1 9 9 9 9 2 7 3 9 2 13 13 2 16 13 10 9 0 2 1 15 9 10 1 9 9 13 2 7 15 9 10 2 1 15 9 15 1 9 0 13 2
65 1 0 3 13 2 16 1 9 2 1 15 16 1 9 13 2 16 15 0 13 9 2 16 9 2 7 15 15 2 3 13 13 16 9 9 2 15 13 10 9 13 2 13 2 7 16 13 4 15 15 9 2 7 0 2 7 0 2 1 15 13 1 9 9 2
21 7 15 13 9 9 2 15 9 13 9 9 1 13 1 0 0 9 1 13 9 2
16 3 16 9 13 13 2 7 9 13 1 15 9 13 4 15 2
35 1 0 13 2 16 9 0 13 1 15 15 13 1 9 1 10 9 2 3 15 9 2 7 1 15 15 13 1 15 16 9 0 1 9 2
28 7 13 9 2 16 9 9 1 9 13 9 1 13 2 7 9 0 15 9 2 16 13 16 9 13 1 9 2
20 15 3 13 16 15 9 13 13 9 10 1 9 13 2 16 9 7 9 9 2
17 7 3 1 15 3 13 13 1 9 15 9 15 10 9 0 13 2
31 13 13 2 16 16 9 13 9 9 2 3 1 15 15 13 0 9 7 9 2 15 15 1 9 9 15 13 2 13 0 2
17 13 3 16 1 9 13 15 9 2 7 1 9 13 15 1 9 2
13 3 10 9 0 13 1 9 3 16 9 1 9 2
10 1 15 9 13 9 0 2 16 9 2
42 15 7 13 1 9 0 7 0 2 16 1 0 9 13 0 16 1 9 2 16 9 1 9 2 7 1 0 0 9 13 1 0 2 16 3 0 1 15 9 9 13 2
24 1 15 7 9 13 0 9 2 1 15 9 0 13 15 13 2 16 1 15 9 13 0 9 2
14 1 0 9 13 2 16 9 13 9 9 2 7 9 2
27 3 1 9 9 1 15 13 16 9 9 9 13 2 15 13 16 13 15 9 7 16 9 2 7 16 9 2
25 1 9 7 1 9 12 13 2 3 9 0 2 9 2 7 9 0 2 3 0 2 7 9 9 2
22 16 0 9 13 15 16 9 1 0 9 15 13 1 9 1 9 2 3 13 9 9 2
11 3 9 1 15 9 3 13 15 9 13 2
27 16 3 13 15 2 13 16 13 1 9 1 9 13 2 1 10 9 13 1 15 9 15 13 9 9 13 2
15 7 9 9 13 1 9 0 3 13 15 9 1 9 13 2
16 3 3 9 9 3 13 13 15 2 1 3 13 15 0 9 2
26 10 7 3 9 13 0 13 2 16 9 2 16 13 13 9 9 7 9 2 13 9 9 1 9 0 2
24 7 3 15 13 2 16 16 9 13 1 15 9 13 9 9 0 2 3 7 9 1 15 9 2
19 7 16 13 1 9 2 1 9 13 2 16 15 9 13 3 13 1 13 2
26 7 13 9 15 1 9 13 2 7 3 15 9 13 2 1 15 15 13 16 13 3 13 15 16 13 2
12 7 16 1 9 4 13 2 13 15 9 13 2
24 7 13 0 16 2 1 9 0 9 13 2 0 13 1 9 1 9 2 16 9 13 13 13 2
16 7 3 15 13 13 2 16 9 1 15 9 15 13 9 13 2
21 7 1 15 16 1 9 1 9 13 2 13 15 9 1 9 13 7 3 7 0 2
23 3 9 13 2 16 3 13 0 15 1 15 9 15 13 0 9 2 16 1 9 0 9 2
24 1 0 13 2 16 9 13 9 9 1 9 16 13 2 16 13 9 2 3 7 16 13 9 2
29 1 0 13 2 16 9 9 16 3 13 9 13 7 13 2 13 3 15 9 0 1 9 0 9 2 13 9 9 2
13 3 2 0 13 12 9 15 9 13 1 15 9 2
18 7 9 13 13 15 9 0 1 9 9 0 2 1 15 13 9 13 2
14 3 1 15 3 13 13 0 9 15 9 1 9 13 2
15 3 2 1 15 9 10 9 13 16 9 0 1 15 13 2
13 3 16 13 9 13 2 9 0 1 15 3 13 2
21 7 3 13 16 3 13 1 9 13 15 9 0 1 9 13 2 1 15 13 13 2
14 3 7 13 2 16 1 15 13 9 0 1 9 13 2
37 12 13 1 9 9 2 15 13 2 16 9 10 0 3 13 15 9 16 9 13 13 2 16 9 0 3 13 13 1 9 0 16 16 1 9 13 2
35 7 9 0 1 13 15 1 9 13 2 15 13 13 2 13 9 0 1 9 15 2 15 13 9 1 9 13 2 7 13 15 1 9 0 2
33 7 1 13 15 13 1 9 13 2 9 15 13 13 1 15 2 16 9 0 13 13 1 9 2 1 9 13 15 13 1 9 13 2
40 0 2 16 1 15 9 1 9 0 13 2 3 13 0 15 13 2 16 15 9 13 15 13 2 1 0 0 13 9 0 1 9 0 16 9 0 1 9 0 2
23 1 0 13 2 16 9 0 13 3 13 3 12 9 1 15 9 15 0 1 9 0 13 2
29 3 15 13 15 9 1 9 13 13 2 7 9 15 3 13 1 9 0 9 13 0 7 0 9 9 13 1 9 2
18 1 0 13 2 16 1 9 10 13 9 0 2 3 16 9 13 13 2
44 13 7 3 9 0 1 9 0 2 1 9 3 13 2 3 16 1 9 0 2 7 1 9 0 1 9 0 7 9 9 2 16 3 9 15 13 1 13 2 15 9 15 13 2
22 7 1 9 0 9 2 9 15 1 9 13 16 9 13 13 2 3 13 1 9 0 2
22 13 13 2 16 1 10 9 13 1 9 2 15 13 9 13 13 2 0 13 13 9 2
7 12 1 9 1 9 13 2
14 15 1 9 15 13 9 9 2 7 1 9 9 13 2
21 1 15 3 9 15 13 1 9 1 9 13 2 15 9 1 10 9 13 9 9 2
88 1 3 10 9 13 1 9 2 9 7 3 13 1 15 13 0 2 1 15 9 3 13 13 1 9 9 0 2 16 1 15 9 3 13 9 2 15 13 9 9 2 16 1 0 2 16 3 13 9 1 9 0 2 16 15 13 0 2 13 9 16 13 9 0 2 16 16 9 0 13 1 13 16 13 1 9 1 9 2 16 13 1 9 0 1 9 0 2
40 7 1 15 9 15 13 1 9 15 13 9 9 2 7 15 9 2 13 1 1 0 2 16 3 9 13 3 0 2 15 16 9 9 0 13 15 9 9 13 2
8 9 7 0 9 7 9 13 2
14 3 3 9 13 0 1 9 15 2 3 9 7 9 2
17 9 3 2 1 13 9 13 2 3 13 16 1 9 1 9 13 2
27 7 3 1 9 15 0 1 15 9 1 9 3 0 13 2 0 0 3 13 2 7 3 1 9 9 13 2
30 1 0 3 13 2 16 9 1 9 9 3 13 0 0 2 16 1 9 0 2 16 3 13 16 1 9 1 9 13 2
9 9 3 0 13 1 9 3 0 2
13 3 1 15 9 3 13 15 13 15 9 1 0 2
17 7 9 0 13 1 9 0 2 15 13 13 9 13 0 7 0 2
22 1 0 13 2 16 15 9 13 9 1 9 9 13 7 1 9 9 13 2 3 0 2
15 7 3 9 15 13 1 9 13 2 13 15 9 7 9 2
29 7 16 13 16 9 13 13 1 9 15 7 13 7 13 1 0 9 2 3 13 13 16 15 9 1 9 9 13 2
33 3 3 1 3 9 13 1 16 9 15 13 1 9 2 7 9 1 9 2 16 3 0 0 2 1 15 9 13 2 9 13 13 2
19 7 9 13 13 1 15 0 16 9 1 9 13 13 9 15 13 1 9 2
27 3 3 9 0 15 13 9 1 9 1 9 13 2 16 3 13 3 16 13 2 0 13 9 13 7 0 2
30 16 3 9 9 13 3 13 1 9 9 1 9 0 2 16 1 13 4 2 15 9 13 13 16 15 9 0 9 13 2
92 1 0 13 2 16 13 13 1 0 9 1 0 9 2 1 15 16 1 15 13 15 9 2 16 9 1 0 3 13 1 9 9 1 10 0 0 9 2 16 0 9 1 9 7 9 13 9 13 2 16 13 3 2 7 13 1 9 0 2 1 16 0 13 1 9 2 16 13 13 9 15 1 9 0 1 9 2 7 3 1 9 0 2 16 1 2 8 12 2 13 4 2
24 3 1 10 9 13 0 1 9 0 9 13 2 15 15 2 1 15 9 2 3 13 3 13 2
22 9 7 9 7 9 15 0 2 15 9 0 1 9 13 2 13 1 15 9 7 9 2
34 3 13 15 9 9 15 1 9 3 13 13 1 15 9 2 1 15 15 13 1 9 1 15 9 2 16 15 1 9 13 1 15 9 2
30 16 3 13 16 9 13 9 13 2 1 15 9 13 9 0 2 15 9 9 9 13 1 0 3 13 1 13 9 15 2
30 13 16 13 1 9 1 9 9 13 2 16 9 13 2 15 1 15 13 9 13 2 13 9 9 1 9 7 15 15 2
63 7 1 15 2 1 15 9 15 13 1 9 2 13 1 9 9 13 2 3 16 7 15 9 7 13 1 15 13 0 15 1 13 9 13 2 16 13 1 9 0 2 16 13 9 0 2 7 16 9 0 13 15 9 1 15 1 15 9 15 13 9 13 2
30 3 2 16 9 1 9 13 9 1 3 9 0 1 15 13 1 9 13 2 13 15 9 13 15 9 2 16 13 4 2
16 3 1 15 16 15 13 16 9 2 13 15 7 15 9 13 2
13 0 7 3 13 13 9 0 7 0 2 1 15 2
30 1 15 3 13 9 0 2 15 13 15 16 9 2 13 0 7 0 2 9 0 13 2 15 13 0 2 13 9 13 2
26 1 3 9 13 2 1 9 2 13 13 15 9 13 0 2 0 13 16 9 13 13 9 9 1 9 2
16 9 9 2 16 13 9 2 13 0 2 16 9 9 13 0 2
20 16 3 3 13 9 13 13 0 1 9 1 9 2 0 13 16 13 9 15 2
20 7 3 0 9 2 16 13 1 9 0 13 9 0 15 15 9 0 13 9 2
28 16 9 13 3 13 9 15 9 2 3 16 1 15 13 13 2 15 9 13 13 9 15 9 1 15 0 13 2
15 13 3 16 12 9 3 1 9 13 13 16 1 9 10 2
31 13 3 0 2 16 0 13 13 16 9 13 15 13 1 9 0 13 1 15 7 16 9 1 9 2 7 16 9 1 9 2
23 12 7 9 3 13 12 16 12 15 13 1 15 16 9 1 9 2 7 16 9 1 9 2
24 13 3 16 9 13 13 1 0 9 9 1 9 7 16 9 1 9 2 7 16 9 1 9 2
42 15 7 13 1 12 9 2 15 15 13 16 9 15 2 16 2 1 9 7 9 13 1 0 16 1 9 2 13 16 15 2 3 9 2 13 3 9 15 2 3 9 2
32 13 3 16 2 1 13 0 4 15 13 1 9 2 15 13 15 9 15 2 16 3 9 13 13 15 2 16 13 9 13 0 2
37 16 3 10 13 1 9 4 1 15 13 1 9 2 3 9 13 9 13 15 16 9 2 7 13 1 15 9 2 16 3 9 13 1 9 1 9 2
50 16 9 13 13 9 13 2 3 13 15 16 1 9 13 13 1 9 2 1 15 9 2 16 7 9 0 2 16 9 0 15 13 1 15 9 16 9 1 9 2 9 7 13 1 13 16 9 1 9 2
42 1 9 13 2 9 13 3 13 13 15 16 9 16 1 15 16 13 9 0 13 2 15 3 13 9 1 15 16 15 9 13 9 13 7 15 13 2 3 13 13 9 2
16 3 3 13 13 9 15 16 1 16 13 1 9 15 13 0 2
28 16 1 9 13 13 9 13 2 15 3 13 16 9 13 13 9 15 7 15 9 0 2 7 16 13 9 15 2
15 13 7 9 15 3 1 0 13 0 2 1 15 15 13 2
42 16 7 13 16 3 13 15 9 9 1 15 13 0 9 13 2 16 1 15 13 13 9 13 2 15 3 13 16 16 15 13 0 3 13 9 9 13 1 13 9 13 2
26 3 3 1 15 16 10 0 0 13 2 13 16 3 9 9 13 13 15 9 16 1 15 13 9 13 2
29 1 15 16 9 13 13 15 16 9 3 16 1 15 13 9 13 2 13 16 9 9 1 9 13 0 2 1 9 2
55 13 3 1 12 9 1 8 2 16 1 0 9 2 1 15 10 0 13 4 2 9 1 15 13 2 7 1 15 7 1 15 7 1 9 0 7 0 9 15 13 2 9 9 13 2 7 3 13 9 0 9 1 15 13 2
12 9 7 10 13 1 9 1 10 9 9 13 2
18 0 9 2 3 16 15 9 9 1 9 13 9 15 13 9 10 9 2
23 16 16 9 13 9 2 7 1 9 10 13 9 1 15 15 9 2 7 15 9 2 13 2
46 9 0 1 15 13 15 1 10 9 2 13 16 13 15 9 2 7 3 9 15 2 16 9 9 15 13 1 9 9 2 13 15 9 1 9 9 15 13 1 9 2 7 0 9 15 2
64 1 7 9 9 15 13 3 13 16 13 9 1 15 9 13 15 15 13 9 9 13 2 0 13 13 15 16 1 9 0 9 13 13 13 15 9 9 3 1 15 9 0 2 1 0 9 13 15 1 15 0 2 7 1 0 13 4 16 9 15 13 13 9 2
28 1 15 3 9 9 2 13 13 16 9 15 13 1 15 0 2 13 7 9 3 2 7 9 1 9 7 9 2
35 15 3 15 1 9 7 9 13 13 2 3 13 15 13 9 2 16 9 1 15 13 3 13 1 15 9 2 16 15 9 9 13 3 13 2
37 15 7 15 3 13 0 16 3 0 13 9 2 13 15 13 9 2 16 9 10 13 15 16 1 15 15 13 13 2 16 1 0 13 1 9 0 2
16 16 0 9 10 1 15 13 3 13 2 15 9 9 13 13 2
21 1 3 9 9 13 0 2 15 0 13 16 9 3 1 9 0 15 13 9 15 2
21 15 3 0 0 13 3 16 0 9 1 9 0 2 7 16 9 1 9 15 13 2
11 7 3 13 13 9 15 9 1 9 0 2
10 13 3 1 0 9 13 0 15 13 2
10 9 15 0 3 13 15 16 15 13 2
11 9 3 13 15 0 16 9 10 15 13 2
20 13 7 9 9 0 13 16 15 0 9 13 9 9 15 13 2 16 13 4 2
11 9 3 13 9 13 2 9 0 9 13 2
25 1 15 7 16 9 13 13 9 9 2 13 16 15 0 9 13 9 16 9 0 2 16 13 4 2
29 0 13 3 16 15 15 13 9 15 9 0 2 13 15 9 9 2 16 9 15 13 15 9 15 15 13 0 9 2
14 9 7 0 13 0 9 0 9 0 2 7 15 13 2
24 0 13 3 16 15 9 13 0 9 15 9 13 2 16 1 15 16 15 0 9 9 13 13 2
14 15 13 0 9 0 16 1 15 9 1 15 9 13 2
10 9 7 0 13 9 9 10 9 13 2
8 15 9 2 1 0 9 9 2
25 16 0 9 13 1 15 16 13 13 2 1 15 16 13 0 9 1 9 9 13 1 15 1 0 2
19 3 3 0 0 13 0 2 16 13 3 9 13 9 2 15 13 9 9 2
16 7 13 0 0 2 16 9 1 15 0 3 13 1 9 13 2
38 9 7 9 13 13 3 1 9 13 2 3 1 9 15 9 13 2 7 1 16 9 13 15 9 12 1 15 2 16 9 1 9 2 7 9 1 9 2
16 10 9 1 3 9 13 1 3 9 13 9 15 13 9 9 2
13 9 7 0 15 0 9 13 2 13 15 0 9 2
19 15 16 13 9 0 9 13 2 3 3 9 13 13 15 1 15 13 15 2
14 1 15 7 3 3 1 0 9 9 1 9 9 13 2
43 16 0 9 9 13 9 15 13 9 9 2 9 7 15 9 13 0 9 13 2 9 15 13 9 13 2 16 1 13 13 2 0 13 16 1 9 15 9 13 9 0 9 2
37 3 13 16 0 9 7 9 9 13 7 15 9 2 7 9 9 7 9 2 9 0 1 15 9 13 2 13 9 0 2 16 13 1 12 1 9 2
19 15 3 9 3 13 9 9 16 16 13 9 16 9 0 13 1 15 9 2
22 9 3 13 2 7 9 15 2 1 1 9 13 1 15 1 9 2 16 13 15 0 2
47 1 15 7 13 15 13 1 9 9 9 2 15 2 1 15 16 13 13 9 9 9 13 2 13 10 9 13 9 2 7 16 15 9 13 1 12 9 2 16 3 3 9 9 13 1 13 2
52 1 10 9 13 13 15 15 13 0 1 9 7 0 1 9 2 13 0 9 0 9 2 16 9 9 2 15 13 0 9 9 2 0 13 16 9 9 7 9 7 9 2 15 13 1 9 9 2 15 13 9 2
12 15 3 9 7 9 13 1 15 16 13 9 2
47 10 9 15 13 15 9 2 13 16 9 15 9 15 13 15 9 2 16 9 0 7 0 0 13 9 15 2 1 15 13 0 7 0 2 7 3 9 9 15 13 13 13 2 15 13 9 2
13 13 4 3 1 0 16 7 9 7 9 13 15 2
25 15 7 9 9 13 13 4 2 13 15 9 2 7 0 7 0 2 16 1 9 9 13 1 9 2
10 3 3 13 9 7 9 13 1 9 2
28 7 16 9 0 9 9 13 2 16 1 0 13 4 2 13 13 16 0 9 3 9 0 7 0 1 9 13 2
57 16 3 10 15 1 15 3 13 2 1 15 15 13 1 15 13 13 2 13 16 9 9 15 3 13 1 15 13 7 1 9 2 13 1 9 15 1 15 1 9 13 2 16 9 1 9 13 13 15 9 15 9 15 1 9 13 2
25 7 1 15 9 13 9 9 0 13 15 9 13 2 15 13 9 13 15 0 2 1 16 15 13 2
12 9 2 0 13 10 9 0 1 9 13 13 2
17 0 7 9 13 13 9 9 2 15 1 9 9 9 9 13 13 2
37 15 7 9 13 13 16 15 9 0 13 13 1 15 9 16 0 9 2 16 9 0 7 0 2 15 3 13 13 1 15 13 16 9 0 13 13 2
10 3 13 16 15 9 1 9 9 13 2
12 7 0 9 15 9 2 15 15 13 0 0 2
8 3 10 9 9 13 13 9 2
19 15 7 15 13 1 9 9 3 13 9 3 2 7 9 1 9 7 9 2
18 3 10 9 1 15 13 2 3 1 9 2 7 1 15 2 3 9 2
16 13 3 16 13 3 13 9 3 2 7 9 1 9 7 9 2
25 7 9 13 2 16 13 9 2 13 9 9 15 13 1 9 2 7 3 15 9 1 9 7 9 2
9 13 7 9 13 9 0 16 0 2
22 16 3 9 0 15 13 1 9 0 13 0 9 2 0 3 9 0 13 15 0 9 2
21 3 13 7 15 0 9 13 9 2 16 15 13 1 9 2 1 15 13 9 0 2
14 16 9 0 13 13 9 9 16 9 0 13 1 13 2
50 1 3 1 15 15 13 16 13 2 16 9 3 13 13 16 15 13 13 2 7 16 1 15 13 13 2 3 7 9 0 13 2 7 13 13 1 15 16 13 4 13 1 9 1 9 2 15 13 9 2
22 7 3 13 16 10 15 13 15 9 3 13 2 13 15 0 1 15 15 13 0 9 2
29 7 0 3 1 15 15 13 0 9 2 0 9 3 13 2 15 3 13 1 9 15 9 13 2 16 15 13 15 2
27 16 15 9 0 2 16 13 1 9 0 2 15 3 1 9 13 9 10 0 9 2 3 13 9 9 0 2
33 15 7 13 1 9 15 2 13 9 0 3 15 3 2 7 3 15 1 15 9 13 2 16 1 9 9 13 1 9 9 9 9 2
20 1 15 13 16 1 9 9 0 13 9 0 2 16 13 0 1 9 0 9 2
40 1 9 7 15 1 9 13 2 13 9 0 1 9 0 2 3 9 0 2 15 13 0 0 2 3 13 16 10 13 1 9 1 15 9 2 13 1 9 15 2
17 7 1 15 2 1 13 15 9 0 13 9 0 2 1 9 0 2
20 1 13 7 9 9 2 16 13 9 9 9 2 13 3 1 9 0 9 0 2
14 3 13 7 0 16 9 13 9 9 2 16 1 9 2
19 9 7 1 9 13 2 1 13 0 9 2 13 1 13 0 9 1 13 2
19 3 9 15 13 0 1 9 7 0 1 9 2 3 9 2 13 3 0 2
19 13 7 9 9 15 9 1 9 13 13 13 2 9 13 3 16 13 9 2
31 0 13 3 16 9 3 13 13 15 15 2 1 13 13 1 9 2 15 13 9 1 9 2 7 1 9 2 15 13 9 2
35 7 1 15 10 9 13 1 10 9 2 1 15 13 15 9 2 3 13 2 1 10 9 16 9 2 16 9 15 13 1 9 1 9 13 2
22 16 7 1 0 1 9 9 13 13 1 9 9 9 13 2 13 9 7 0 1 3 2
18 3 3 9 13 13 1 9 3 9 15 9 2 7 9 1 15 13 2
30 9 0 2 1 13 13 1 9 7 9 2 13 1 0 9 16 13 9 2 15 9 2 1 12 8 2 13 0 15 2
11 7 1 15 2 1 16 13 9 2 13 2
12 9 3 0 3 13 13 0 9 1 15 9 2
60 9 7 9 9 13 1 9 0 9 2 16 0 9 13 9 15 9 9 1 15 13 2 7 13 15 2 7 3 13 15 1 13 2 16 9 13 9 1 0 9 2 15 3 3 13 9 1 15 13 9 2 7 13 2 7 13 15 0 9 2
14 9 7 13 15 9 13 9 15 2 15 13 9 9 2
12 9 7 1 15 13 0 9 2 3 13 13 2
18 13 3 9 1 9 13 1 9 2 3 9 13 13 9 16 15 9 2
19 9 7 3 13 12 9 9 13 2 7 1 9 10 13 16 9 9 13 2
8 1 9 0 9 13 1 9 2
38 9 15 1 9 1 9 13 13 2 1 9 15 13 15 9 1 10 9 13 2 16 7 9 9 15 13 1 9 2 1 15 13 15 13 1 9 9 2
19 3 9 0 13 9 0 2 10 7 9 0 3 13 1 15 9 0 13 2
12 7 15 15 9 13 2 13 15 15 9 13 2
15 0 7 1 0 9 13 9 3 0 2 16 1 13 4 2
13 1 15 7 9 9 15 9 9 1 9 9 13 2
14 16 7 9 10 9 9 9 13 2 13 1 15 9 2
5 0 2 9 9 2
7 0 7 2 16 1 9 2
25 15 0 15 13 9 2 9 15 15 13 0 9 9 15 13 1 9 2 16 9 0 9 9 9 2
12 0 7 9 9 9 1 15 9 0 9 13 2
7 9 3 1 9 0 13 2
29 3 15 9 13 0 9 2 3 13 13 0 7 1 15 3 0 13 9 9 2 3 9 13 13 2 16 7 9 2
20 15 7 13 13 9 7 9 15 9 13 2 16 10 9 0 13 0 7 13 2
10 3 15 9 1 9 10 0 13 13 2
36 7 15 9 3 0 13 2 16 9 3 13 2 16 9 13 7 13 2 7 13 0 1 9 7 13 0 7 0 9 2 15 1 9 3 13 2
23 15 9 0 15 13 1 15 15 13 1 9 7 9 9 2 16 10 9 13 1 10 9 2
31 15 7 9 13 0 7 3 3 15 9 15 13 2 1 9 2 15 13 1 9 1 0 9 2 7 1 9 9 7 9 2
17 1 15 9 15 13 4 13 7 13 1 15 9 13 13 1 9 2
8 3 10 9 13 1 9 10 2
32 9 7 0 3 0 0 13 2 16 13 1 0 0 9 9 2 16 13 2 15 13 9 9 9 0 13 2 13 15 0 3 2
29 15 1 9 13 2 1 15 9 13 9 2 3 15 1 15 9 0 9 3 13 2 7 0 1 15 13 1 9 2
17 9 7 1 15 0 13 2 16 9 13 0 2 1 15 9 13 2
11 3 3 1 9 13 9 9 9 1 9 2
9 1 9 7 9 13 9 9 9 2
44 1 3 9 13 1 15 9 13 9 2 9 7 15 1 16 13 9 2 13 1 9 9 2 15 13 15 10 9 0 2 0 13 16 9 15 13 15 16 0 9 13 1 9 2
20 3 13 9 2 1 12 8 2 1 9 13 2 13 16 13 0 15 7 0 2
16 3 1 9 9 13 3 13 16 1 16 12 13 13 16 15 2
44 1 15 9 2 1 12 8 2 9 2 1 15 9 9 7 9 13 2 13 9 2 1 15 9 13 1 9 7 9 9 2 16 1 15 13 13 16 9 9 0 9 9 13 2
16 1 9 7 9 2 1 15 9 9 13 2 13 7 9 9 2
8 13 7 15 9 9 1 9 2
8 13 16 9 9 13 9 15 2
13 13 3 2 16 13 0 9 2 16 13 0 9 2
11 13 3 1 9 9 0 9 9 1 9 2
33 1 3 9 0 13 1 16 15 13 15 13 2 13 1 15 15 1 3 9 16 13 1 15 0 7 9 2 1 15 13 9 9 2
42 15 0 1 15 9 13 3 13 2 7 9 1 9 13 2 16 3 15 15 13 3 13 9 3 2 7 9 3 2 15 1 15 3 13 9 9 2 7 9 1 15 2
18 3 7 13 9 7 9 1 15 12 13 13 16 13 15 9 1 15 2
16 16 7 13 13 15 13 2 0 13 16 0 9 0 9 13 2
14 3 13 16 15 9 13 9 0 2 15 0 9 13 2
20 7 1 0 9 2 0 9 9 13 13 2 13 1 9 9 7 1 9 15 2
39 1 3 13 15 9 9 2 13 0 7 13 9 9 2 13 16 15 15 9 13 13 7 0 0 2 13 1 15 15 13 3 0 2 7 15 9 13 0 2
14 1 9 7 9 7 9 7 9 13 9 9 7 9 2
23 1 15 13 0 13 9 0 1 9 7 9 2 7 9 7 0 2 7 9 7 9 13 2
11 9 7 1 0 13 9 7 15 15 13 2
15 1 0 0 9 2 15 3 3 13 9 2 3 15 15 2
12 1 15 9 13 16 13 9 15 7 9 15 2
7 15 7 13 0 9 15 2
17 15 9 2 1 9 2 15 13 9 13 2 7 15 1 9 13 2
14 13 3 2 15 13 9 2 13 10 9 7 9 13 2
16 3 9 13 9 13 16 9 15 2 9 7 10 9 9 13 2
40 15 7 13 1 9 1 9 0 1 9 15 9 2 16 15 13 1 15 1 15 9 2 3 13 1 9 0 2 16 13 3 0 0 9 15 13 1 3 9 2
17 3 15 9 9 7 9 13 13 16 13 13 9 15 13 0 9 2
40 1 9 3 0 15 13 2 16 9 15 13 1 9 9 1 9 0 2 3 13 0 7 1 9 2 16 3 13 13 9 0 15 9 9 13 1 9 10 9 2
22 3 13 7 1 9 9 16 9 15 15 13 1 10 9 2 3 16 15 0 9 13 2
14 13 3 16 10 9 0 13 1 15 9 1 9 13 2
36 15 3 3 13 0 1 9 9 2 15 13 1 12 8 2 16 9 15 13 1 9 2 3 13 1 9 13 2 7 1 9 15 13 1 9 2
34 9 3 0 13 0 9 15 9 13 13 1 9 0 2 3 9 1 15 15 13 16 13 1 9 15 9 2 16 1 9 0 15 9 2
17 3 3 15 13 9 13 3 9 0 2 16 13 9 1 0 9 2
20 3 2 1 15 9 13 3 13 15 13 0 9 1 9 0 7 13 10 9 2
13 3 9 0 13 15 1 9 13 1 9 0 9 2
10 9 3 9 1 10 13 13 9 0 2
18 0 13 7 16 15 13 15 9 0 1 0 16 13 9 15 0 13 2
22 1 9 7 15 9 3 13 15 9 0 2 7 13 9 0 1 9 2 15 13 9 2
9 13 3 9 9 2 7 15 3 2
34 1 9 7 3 13 9 16 13 1 9 1 15 9 2 16 9 13 2 1 10 9 2 1 10 9 7 9 0 2 1 13 15 0 2
14 1 9 3 13 0 9 0 1 9 2 16 13 4 2
51 16 0 9 1 0 13 3 9 0 2 13 15 13 16 15 13 16 9 9 2 15 13 9 9 2 13 15 9 1 9 0 2 3 1 16 9 13 2 7 1 16 13 9 9 2 15 13 9 1 9 2
35 1 9 3 9 9 13 3 13 2 16 0 9 9 13 2 7 10 9 9 13 13 1 15 16 13 9 9 13 9 2 16 1 15 13 2
17 9 7 0 13 9 9 1 0 10 9 9 2 3 13 13 9 2
32 1 0 9 9 9 13 1 9 2 7 9 9 9 1 9 2 16 7 1 15 9 9 13 1 9 2 7 9 1 0 9 2
45 13 3 12 8 2 12 3 3 9 13 1 15 2 7 1 9 7 9 2 9 7 9 13 2 16 15 15 13 2 3 16 3 13 9 2 7 16 15 9 13 15 1 13 15 2
26 3 3 7 9 9 2 1 1 0 9 0 9 13 2 15 13 15 9 7 3 9 2 7 0 13 2
22 16 1 9 0 15 13 1 9 2 3 1 9 0 7 0 15 13 1 9 7 9 2
18 7 15 13 9 15 0 9 13 1 9 2 16 3 13 13 9 13 2
12 9 3 13 9 1 9 16 4 1 9 13 2
11 9 7 7 9 13 9 9 16 9 9 2
19 15 9 1 9 0 9 13 13 1 0 9 2 7 0 1 9 0 9 2
22 1 9 3 1 9 0 9 13 9 9 2 7 9 9 13 1 9 2 15 13 9 2
41 9 0 3 13 1 9 13 1 0 9 16 1 16 13 1 9 0 9 2 16 9 9 3 3 13 9 1 9 9 16 1 15 9 2 16 16 13 1 9 9 2
17 13 7 15 9 15 1 9 13 13 2 16 15 9 7 9 15 2
28 15 7 3 13 16 13 9 13 9 1 15 9 7 9 2 7 3 1 15 9 13 2 7 3 13 1 15 2
18 13 3 9 0 13 15 9 7 9 1 9 13 2 3 16 3 13 2
11 15 13 1 9 15 13 1 9 10 9 2
19 3 13 16 9 13 15 0 9 7 9 2 1 15 13 13 1 9 13 2
7 15 7 13 1 0 9 2
32 13 3 2 1 15 16 9 13 1 0 9 1 0 9 2 16 13 15 15 9 2 1 15 15 9 9 15 13 13 0 9 2
23 3 9 9 2 15 9 1 9 13 1 13 1 0 9 2 15 9 7 9 9 13 13 2
31 9 1 15 9 13 1 15 9 2 13 3 9 15 9 2 16 9 1 9 9 13 9 7 9 1 9 1 15 0 13 2
23 13 4 7 16 9 0 13 13 9 15 1 9 1 15 13 1 0 9 2 15 9 13 2
21 7 1 15 9 2 15 1 13 3 13 9 13 2 13 1 9 9 9 0 13 2
40 13 3 2 1 8 12 1 1 9 9 13 2 3 9 13 4 13 15 0 9 2 7 15 13 2 9 9 13 2 1 9 9 13 2 7 9 13 16 9 2
43 7 13 1 0 9 13 2 15 13 0 9 2 9 7 9 10 9 2 1 15 0 13 13 15 9 2 1 15 13 10 9 9 2 0 10 15 9 2 15 0 9 13 2
21 9 13 2 8 12 2 16 9 2 16 13 15 9 9 13 2 1 9 9 13 2
22 1 9 7 9 3 15 13 16 9 0 2 16 1 9 9 3 13 15 16 0 9 2
22 13 7 9 15 4 13 1 9 9 0 2 3 3 16 9 9 0 13 1 9 0 2
29 13 3 2 1 8 12 1 1 9 9 13 2 3 9 13 4 13 15 0 9 2 7 15 13 2 9 9 13 2
15 3 3 9 9 13 9 1 9 2 16 1 9 13 13 2
20 1 9 0 15 9 9 13 2 16 15 15 1 15 13 2 13 1 15 9 2
9 0 3 0 9 10 0 9 13 2
9 15 7 9 3 13 9 9 13 2
16 9 7 9 1 9 9 3 13 9 0 2 7 0 0 9 2
34 9 7 3 0 3 13 0 16 13 2 13 3 9 9 7 0 13 2 7 13 15 16 15 13 2 13 3 9 9 9 15 9 13 2
15 15 3 1 0 9 13 0 13 16 9 13 13 9 13 2
20 3 0 9 15 9 13 1 0 13 9 2 9 13 1 12 7 0 15 9 2
20 9 3 15 1 15 9 13 2 7 1 15 13 0 2 7 1 15 13 0 2
56 16 3 10 9 13 9 15 9 13 2 7 1 9 9 13 2 13 16 15 9 13 13 1 9 9 2 7 1 15 13 2 7 3 15 15 9 13 0 7 0 2 3 9 0 2 1 0 9 2 13 0 9 7 3 9 2
16 3 3 9 0 0 13 2 7 3 13 15 1 10 9 9 2
24 9 3 13 1 9 1 9 0 16 13 13 2 16 9 0 13 9 1 9 0 1 0 9 2
25 9 7 0 1 9 15 13 1 10 9 2 13 9 1 0 9 7 0 9 2 15 1 9 13 2
18 3 3 13 16 1 9 0 13 1 13 9 1 0 9 7 0 9 2
19 3 3 15 13 10 9 9 2 16 1 9 0 15 13 16 13 7 13 2
12 9 0 13 4 1 9 13 1 9 10 9 2
9 16 3 13 15 13 1 9 0 2
12 3 9 2 16 9 13 2 13 9 1 9 2
39 15 3 9 0 9 3 13 2 1 15 13 12 9 2 16 12 9 2 1 15 9 2 8 12 2 1 9 13 2 15 1 1 9 9 13 2 3 9 2
27 3 9 2 1 1 12 9 13 12 9 2 3 13 13 16 1 9 7 9 2 16 13 3 1 15 9 2
27 7 1 15 2 3 13 0 9 1 9 16 9 9 1 9 2 3 1 9 9 2 3 3 1 9 9 2
33 1 1 9 9 13 2 3 9 13 4 15 13 0 9 2 7 15 13 9 9 13 2 1 9 9 13 2 7 9 13 16 9 2
39 0 3 3 13 9 9 9 7 9 2 7 3 9 9 7 9 2 7 3 3 0 13 15 9 13 2 15 1 1 9 9 13 2 13 15 9 9 13 2
22 0 9 9 13 1 15 16 13 1 9 9 13 2 1 15 16 13 2 9 9 13 2
31 0 13 3 9 1 9 13 2 7 3 1 9 2 1 15 16 13 2 15 1 1 9 9 13 2 16 1 9 13 9 2
28 15 3 9 13 13 0 9 2 9 13 7 9 2 1 15 13 9 9 1 15 15 13 1 9 7 9 13 2
33 13 3 9 9 13 1 15 16 0 9 15 13 2 16 7 9 15 13 13 2 16 9 9 13 2 3 3 16 9 9 3 13 2
12 13 4 3 1 16 9 9 9 13 3 13 2
28 1 3 9 9 13 9 2 16 13 4 2 0 13 16 9 9 13 9 9 2 16 3 9 1 9 13 13 2
25 16 3 0 9 3 13 13 9 9 2 7 7 3 15 0 9 2 1 15 0 9 9 9 13 2
15 0 13 7 9 0 1 9 9 13 2 1 13 15 9 2
12 15 3 1 9 13 2 15 9 13 3 13 2
16 9 13 1 9 16 9 1 9 2 7 16 9 1 0 9 2
12 13 7 9 13 13 9 2 7 9 0 9 2
28 9 13 2 8 12 1 0 9 2 16 1 1 9 9 13 2 13 15 2 9 9 13 2 1 9 9 13 2
23 15 3 9 2 16 0 9 13 2 3 0 13 1 9 9 2 16 3 1 9 9 13 2
32 13 3 16 13 1 9 9 2 15 0 13 1 0 1 9 9 2 3 1 9 9 2 7 3 13 15 2 1 9 9 13 2
20 13 7 2 12 15 1 1 9 9 13 2 3 9 13 4 13 15 0 9 2
20 0 13 3 13 16 9 15 13 1 9 2 3 1 9 9 2 7 0 9 2
15 13 7 9 0 1 15 16 13 9 2 16 7 9 0 2
20 3 3 13 9 16 13 9 9 2 7 0 3 13 9 16 13 9 9 10 2
8 9 3 9 0 13 15 9 2
14 13 7 13 16 1 0 13 12 9 2 3 1 13 2
23 13 3 9 2 8 12 2 1 0 9 2 16 2 1 1 9 9 13 2 9 9 13 2
14 3 7 13 13 16 13 15 9 9 2 7 9 9 2
23 7 3 2 16 15 13 9 9 7 9 9 2 1 3 9 9 13 2 3 13 9 9 2
14 7 3 13 13 16 9 9 1 0 1 13 4 13 2
19 7 3 13 13 16 9 9 4 13 1 13 2 16 3 3 13 9 9 2
12 7 7 13 13 16 9 9 13 13 9 9 2
12 3 3 13 16 13 9 9 2 7 15 15 2
21 7 3 13 13 2 1 9 9 2 16 1 0 2 3 1 13 2 13 12 9 2
23 7 16 3 9 13 9 7 9 2 0 9 13 9 7 9 9 0 13 1 15 9 9 2
23 7 16 9 7 9 13 9 9 0 2 13 4 9 9 1 13 9 15 9 1 9 13 2
23 15 3 15 9 13 9 7 9 2 3 13 9 0 2 16 3 15 9 13 13 9 9 2
17 7 16 1 9 7 9 13 15 12 2 16 1 9 7 9 9 2
18 13 4 3 1 0 9 16 9 7 9 13 2 7 15 9 13 13 2
6 9 7 13 0 9 2
17 10 3 9 9 13 15 9 7 15 9 2 16 3 13 1 9 2
14 16 3 9 9 13 0 9 16 9 2 13 15 9 2
24 1 9 7 9 3 13 12 9 2 15 13 0 1 0 9 7 9 2 3 13 1 9 9 2
26 16 3 0 9 0 9 3 9 13 2 13 16 1 9 15 15 0 9 13 2 15 13 1 0 0 2
14 3 9 13 9 9 2 1 15 15 9 13 0 9 2
17 3 13 16 2 16 0 9 13 0 9 2 3 13 7 0 9 2
7 9 3 9 13 9 13 2
18 1 15 0 15 13 1 9 7 9 13 2 13 13 0 7 9 15 2
18 9 7 2 1 13 0 9 2 3 13 9 9 2 7 3 9 15 2
71 9 3 16 0 9 13 2 3 7 9 13 2 7 9 9 7 9 2 7 9 7 9 9 13 2 3 7 3 9 13 15 15 13 9 2 13 15 15 1 9 13 9 2 3 3 13 9 0 0 13 10 9 2 7 0 1 10 2 2 15 3 13 1 9 1 15 13 9 9 15 2
19 3 3 1 9 7 9 13 12 9 2 1 9 7 9 0 9 13 9 2
20 7 13 1 9 0 9 16 15 13 0 0 9 15 15 3 3 13 9 15 2
38 15 3 13 15 9 13 13 0 9 1 9 16 0 9 13 3 9 9 3 13 7 13 2 7 3 0 9 1 9 9 13 2 7 9 13 15 9 2
26 9 3 13 16 9 2 15 13 9 7 9 10 9 7 9 2 15 9 0 7 3 9 9 13 13 2
14 0 7 9 13 0 9 2 16 7 15 15 9 0 2
30 9 0 7 9 2 7 3 9 2 3 13 13 16 1 15 2 1 7 9 3 13 1 15 0 2 7 13 1 15 2
23 13 4 3 9 9 3 3 13 13 16 9 13 1 9 13 2 7 13 9 13 16 9 2
40 15 3 0 9 13 1 10 0 13 2 16 1 1 15 13 2 16 9 0 0 9 13 1 9 16 1 15 9 2 1 15 13 9 0 2 3 3 1 9 2
25 15 0 0 13 4 2 1 15 13 16 9 13 1 0 9 13 1 9 2 3 7 1 9 9 2
23 15 3 9 9 2 7 1 0 7 1 15 9 13 2 3 15 9 13 2 3 9 0 2
26 13 3 13 4 9 9 16 0 2 16 1 9 15 13 9 7 9 2 1 13 1 9 7 9 13 2
11 7 15 13 0 9 13 7 9 15 13 2
21 3 2 1 1 9 9 9 13 2 3 13 7 9 13 9 2 7 9 15 13 2
14 9 3 2 1 13 9 2 13 3 13 16 1 9 2
8 3 13 9 2 13 9 0 2
20 7 3 1 9 0 9 9 13 0 13 2 1 9 0 1 9 13 3 13 2
34 3 1 15 9 0 13 9 2 1 15 13 15 0 9 2 7 0 2 16 1 0 1 0 13 2 7 0 2 16 1 9 1 9 2
68 16 3 9 0 9 2 15 9 15 13 3 1 9 9 2 7 9 9 13 2 15 15 1 15 15 13 1 9 9 7 9 2 16 15 9 1 15 9 13 2 3 9 0 2 15 9 3 13 2 7 15 13 2 7 15 9 13 1 15 2 7 1 13 15 9 1 15 2
12 9 3 9 9 13 2 16 9 13 9 9 2
32 3 7 13 0 9 9 7 13 9 2 16 9 9 2 9 2 7 9 9 7 9 2 7 15 3 15 1 9 0 13 9 2
36 15 7 9 13 13 15 9 13 2 7 1 9 15 9 13 2 16 9 9 13 7 16 9 10 13 1 15 2 7 16 9 13 1 9 9 2
13 9 3 15 9 0 13 2 13 9 15 13 9 2
14 7 15 15 9 13 2 13 9 1 15 13 9 9 2
8 13 3 1 10 9 9 9 2
10 7 0 3 15 9 2 7 9 9 2
20 0 7 1 15 13 13 15 9 2 15 13 13 9 15 2 9 1 9 13 2
18 15 3 3 0 1 9 7 9 0 13 2 7 3 1 9 7 9 2
59 1 15 3 9 2 13 13 16 9 2 16 1 13 4 2 1 9 0 9 2 15 9 0 13 1 15 15 15 1 0 9 13 2 3 9 15 2 1 15 13 10 9 13 2 16 16 9 9 0 13 2 3 9 1 9 13 0 13 2
36 7 15 3 9 2 16 3 13 0 3 1 0 9 2 13 3 3 0 1 9 1 9 2 16 3 9 13 10 0 9 2 15 13 9 9 2
18 3 16 9 15 13 3 13 2 3 13 16 9 3 1 9 15 13 2
8 15 7 13 9 2 3 13 2
14 1 0 13 13 2 9 13 2 15 13 13 9 9 2
18 3 9 0 2 15 13 9 9 2 13 1 9 2 16 0 4 13 2
21 9 3 13 2 15 15 9 4 13 2 1 9 15 1 15 13 16 13 0 9 2
16 12 9 2 1 16 13 9 0 9 2 16 1 9 9 13 2
31 7 3 9 15 9 15 13 15 16 9 0 15 2 1 15 1 9 7 9 13 2 1 15 13 9 0 16 13 12 9 2
22 3 3 13 0 9 0 1 12 7 15 2 1 15 12 13 1 9 0 2 13 9 2
24 16 16 0 9 13 13 9 2 13 9 3 13 15 15 13 15 15 1 9 7 0 1 9 2
21 7 3 0 9 3 13 15 15 2 7 13 1 9 15 13 15 15 16 9 0 2
32 13 3 2 16 9 2 16 13 9 0 1 9 2 3 13 15 16 9 0 2 15 1 10 9 15 13 2 16 13 12 9 2
19 15 9 13 9 16 13 9 0 2 1 15 13 9 15 13 1 9 9 2
8 0 3 9 13 0 13 13 2
12 12 9 16 1 9 13 13 9 0 9 13 2
37 7 3 2 1 1 9 3 13 15 9 0 16 9 0 2 16 13 4 2 3 13 13 16 9 13 2 16 13 9 0 2 9 13 13 1 15 2
35 15 9 13 9 13 9 15 13 7 13 1 9 0 9 2 15 3 15 13 1 9 0 9 13 16 15 13 9 0 1 9 0 9 0 2
16 3 16 9 9 3 13 1 15 13 2 3 13 9 9 13 2
53 1 9 0 2 3 13 13 16 13 15 9 13 1 9 9 1 9 2 16 0 13 15 1 15 2 16 2 1 1 9 9 13 15 15 9 2 16 13 12 1 9 2 15 0 9 13 3 13 0 2 7 0 2
12 13 7 15 16 9 9 15 13 7 9 15 2
12 7 13 9 9 1 16 13 9 13 1 9 2
10 9 0 15 13 1 16 13 9 9 2
14 9 7 9 0 3 13 3 9 2 7 9 7 9 2
16 0 13 16 9 15 13 13 1 9 7 9 2 16 7 9 2
11 0 13 3 16 9 7 9 12 13 9 2
11 3 3 9 13 9 1 9 16 1 9 2
11 13 3 3 1 15 9 0 1 15 9 2
12 3 9 15 9 3 13 16 1 9 1 9 2
13 3 9 7 9 0 9 15 0 13 1 15 9 2
15 7 0 15 13 13 15 9 13 1 9 7 9 9 13 2
7 9 13 9 16 9 9 2
7 10 7 9 13 13 9 2
19 13 7 1 9 9 16 9 0 13 9 9 2 15 13 7 1 9 13 2
23 13 3 9 0 10 1 9 9 2 16 3 9 0 9 0 9 13 2 0 9 3 13 2
15 3 3 15 9 13 1 9 2 3 15 9 9 13 9 2
27 3 15 9 13 1 9 0 9 2 16 13 0 2 0 2 1 9 7 9 0 2 7 9 10 9 9 2
12 7 15 15 13 13 9 9 1 9 1 9 2
56 9 7 0 1 9 3 13 0 1 9 1 9 2 7 1 0 7 1 0 2 16 1 15 0 13 1 9 3 1 9 9 2 3 16 3 3 13 0 15 9 1 15 9 13 2 7 15 13 2 0 9 9 9 0 13 2
30 3 7 9 15 13 1 0 9 1 10 9 2 1 9 0 13 3 13 1 9 9 2 16 13 1 9 15 9 13 2
20 3 3 15 9 9 1 9 13 13 2 1 9 3 1 15 9 0 13 13 2
10 7 3 9 0 0 13 2 16 0 2
42 13 3 13 9 9 7 1 9 9 16 9 9 0 13 2 16 13 15 9 2 7 3 1 15 16 13 15 9 2 16 0 2 9 9 2 9 13 9 7 3 9 2
18 3 3 0 1 9 9 13 2 15 10 13 13 2 3 0 7 0 2
56 7 13 13 16 9 0 9 13 2 16 9 0 13 1 3 1 9 1 9 2 16 15 9 3 13 15 1 9 13 2 16 16 9 0 13 9 1 12 3 2 13 1 9 1 15 2 16 13 7 1 9 9 0 9 9 2
29 1 15 3 0 0 9 13 1 13 2 16 9 9 2 3 9 0 2 0 13 1 9 2 16 1 0 4 13 2
39 16 1 9 9 2 9 15 13 9 9 2 13 0 7 9 2 9 9 9 2 15 13 9 7 13 9 2 3 13 12 8 12 2 16 0 9 9 13 2
11 0 2 3 13 1 15 9 9 7 9 2
10 13 16 1 9 13 9 9 7 9 2
19 10 3 15 13 9 2 13 13 1 9 7 9 2 16 9 13 9 9 2
9 3 9 13 13 1 9 7 9 2
9 3 9 1 9 7 9 13 13 2
8 3 13 13 1 9 7 9 2
21 7 1 2 10 9 1 9 7 9 13 9 2 9 3 0 13 15 0 13 9 2
10 3 9 3 13 13 1 9 7 9 2
12 3 0 13 16 9 13 13 1 9 7 9 2
31 0 2 16 10 9 1 9 7 9 13 9 7 0 1 10 9 2 3 13 16 13 0 1 9 2 1 16 9 13 9 2
12 3 0 13 16 9 13 13 1 9 7 9 2
29 0 2 16 15 9 13 1 10 9 2 3 1 16 15 15 13 1 10 9 2 3 15 13 1 15 16 13 9 2
18 15 3 0 13 7 1 15 9 2 13 16 13 0 7 1 15 9 2
15 13 3 1 9 10 9 2 7 3 13 1 9 7 9 2
45 1 0 13 16 9 15 13 0 1 9 13 1 9 2 15 3 13 13 1 15 2 1 13 0 9 13 2 9 0 2 3 13 1 15 2 16 15 15 13 2 13 13 1 0 2
34 7 15 9 15 3 13 0 1 9 2 7 13 1 15 0 2 1 15 15 13 2 16 3 13 13 1 15 2 7 3 9 13 9 2
25 1 15 9 13 13 2 16 1 9 13 1 9 7 9 2 0 13 16 13 9 7 9 7 9 2
41 1 15 3 15 3 13 13 1 9 7 9 2 1 15 9 3 13 1 9 0 2 3 1 15 9 2 7 15 9 1 15 13 2 13 16 15 9 13 9 0 2
35 7 3 2 1 9 3 13 13 1 9 7 9 2 16 13 4 2 13 16 9 13 10 9 2 10 9 2 7 15 15 3 1 9 13 2
26 0 2 16 9 13 9 10 9 7 9 2 3 3 9 7 9 13 1 9 2 16 16 13 15 13 2
30 15 3 1 12 13 9 2 3 13 1 15 13 9 2 16 13 16 9 3 13 9 0 9 2 16 1 15 13 9 2
23 9 7 3 13 13 9 2 16 9 0 3 13 13 9 2 16 13 9 1 8 1 8 2
66 1 3 1 9 3 13 9 2 7 0 9 2 16 9 3 13 2 7 9 9 7 9 2 7 1 15 13 15 9 7 9 2 7 15 9 7 9 2 7 1 15 13 9 9 7 9 2 7 9 7 9 2 0 13 16 9 15 9 13 13 2 7 13 3 0 2
39 15 7 16 13 13 1 13 9 2 16 3 13 15 15 3 13 15 2 13 1 0 13 15 15 3 13 1 9 0 2 2 3 1 15 9 15 13 0 2
19 3 2 1 9 13 15 9 2 7 0 15 9 2 15 9 13 13 13 2
30 3 2 9 13 9 2 13 3 9 2 1 9 1 9 9 2 16 9 9 2 15 13 9 2 13 9 15 3 13 2
6 7 9 13 9 9 2
24 9 7 0 1 9 9 13 3 13 1 15 9 2 7 0 1 15 9 2 9 3 13 9 2
12 7 3 9 7 9 2 15 13 0 9 9 2
27 9 7 15 13 9 9 2 13 9 13 2 16 7 13 13 0 15 15 13 1 9 2 3 7 15 13 2
17 1 0 13 16 9 13 9 0 2 3 7 9 15 13 9 9 2
22 15 3 13 9 2 16 16 13 2 3 15 9 13 9 10 9 2 7 3 15 9 2
20 7 15 13 1 9 1 9 2 15 3 9 9 13 15 9 2 16 0 9 2
25 13 13 16 2 1 9 13 1 9 7 9 1 9 2 0 13 9 2 1 0 9 13 1 9 2
32 15 3 13 0 2 15 13 1 15 9 1 15 9 2 7 1 15 9 2 7 15 3 0 13 0 2 7 0 1 10 9 2
25 15 9 13 0 2 15 13 1 9 1 15 9 2 7 3 1 15 9 2 7 1 3 7 0 2
18 0 9 13 15 0 2 15 13 1 15 9 2 7 3 1 15 9 2
28 1 3 10 9 13 15 0 16 13 9 2 13 7 15 1 10 9 2 0 13 16 1 9 13 9 9 9 2
26 16 3 9 13 13 1 15 9 1 10 9 2 13 9 1 13 7 13 1 9 2 1 15 9 9 2
50 16 7 9 3 13 13 1 15 9 2 13 9 2 7 3 1 15 9 9 2 16 15 15 13 1 9 9 2 13 3 1 15 9 9 2 3 3 16 13 9 9 1 9 9 2 7 1 9 9 2
50 16 3 13 15 9 2 15 3 1 9 13 2 9 15 3 3 13 13 1 9 9 9 2 3 3 3 16 13 9 9 9 1 15 9 9 7 9 2 7 1 0 9 2 16 15 9 13 0 10 2
27 1 0 13 16 3 13 13 9 9 1 9 1 9 1 9 1 15 9 9 7 9 2 7 1 9 3 2
42 9 7 2 1 13 9 0 2 13 9 9 0 2 15 9 0 13 2 16 9 3 13 16 1 9 2 7 1 9 9 13 1 9 2 3 13 16 9 13 9 9 2
33 7 3 2 1 13 2 9 13 0 16 9 2 16 9 16 9 2 7 15 9 2 1 9 13 9 0 2 0 13 9 16 9 2
33 13 3 16 15 15 13 0 1 13 2 0 13 1 13 2 9 3 0 13 16 9 9 13 2 1 3 9 1 9 13 9 0 2
9 0 2 9 13 2 13 1 9 2
4 0 13 9 2
19 3 1 0 13 13 1 13 2 16 0 13 15 9 2 1 15 13 9 2
33 1 0 3 13 16 0 7 9 1 9 3 13 15 2 16 1 15 9 13 2 3 1 9 2 7 1 15 2 9 13 16 0 2
20 7 16 9 13 1 9 2 9 7 13 9 2 0 0 13 1 9 9 0 2
54 1 7 15 13 15 15 13 2 1 10 9 2 9 7 13 15 2 7 15 1 15 1 9 13 2 1 15 16 15 13 9 7 0 2 0 13 16 9 13 2 7 15 15 13 1 15 2 7 15 15 13 1 15 2
29 13 7 1 9 9 7 9 9 2 7 0 2 7 13 15 2 7 15 13 1 9 2 3 13 16 9 9 13 2
15 15 7 9 13 1 9 2 16 1 9 15 1 9 13 2
37 1 9 7 13 9 1 9 2 7 1 9 2 7 1 15 3 2 16 15 2 16 13 9 2 13 2 7 13 1 15 15 15 13 1 10 9 2
38 1 0 13 16 15 9 13 1 9 15 2 3 1 15 9 9 2 13 15 9 2 9 7 9 2 16 9 13 9 2 9 7 9 2 16 13 9 2
30 15 7 15 13 0 9 9 2 13 13 0 2 7 15 9 1 15 13 2 16 9 7 9 2 7 9 1 9 15 2
17 9 7 7 9 9 13 15 9 9 2 1 10 9 13 15 0 2
42 3 0 9 9 13 1 9 2 15 13 1 10 9 0 2 0 0 15 9 13 1 9 2 9 7 9 2 7 3 2 0 0 9 15 13 1 16 1 9 10 13 2
13 13 7 3 7 9 1 9 2 7 9 1 9 2
28 9 3 1 9 2 16 9 2 16 13 9 2 13 1 9 1 0 9 2 7 1 13 12 2 13 1 15 2
32 9 0 13 1 9 2 16 9 2 1 15 13 2 0 13 1 0 2 7 1 15 16 13 1 9 2 13 9 13 15 9 2
21 9 7 13 1 9 1 15 13 2 7 3 0 1 16 13 9 2 13 9 0 2
8 13 3 3 9 3 13 9 2
33 9 7 3 13 1 9 2 7 3 1 15 15 9 13 2 3 0 1 16 15 13 1 9 9 3 13 1 9 2 13 9 9 2
30 1 0 13 16 9 9 13 16 9 15 2 15 9 13 2 16 9 2 15 13 1 9 9 2 13 15 9 1 9 2
31 16 3 13 1 0 1 16 13 9 2 0 13 16 10 13 1 9 2 13 15 9 2 7 3 9 15 13 13 1 9 2
54 7 16 9 2 1 16 13 1 12 9 0 2 13 1 9 1 0 9 0 2 15 13 13 0 2 13 13 0 1 15 2 16 9 13 13 1 10 9 2 7 3 13 0 1 15 2 16 13 1 9 1 9 0 2
30 16 7 13 1 0 1 16 13 9 2 3 0 13 16 15 15 9 13 1 9 2 13 0 13 2 7 15 9 0 2
68 16 7 13 15 9 13 3 13 1 9 2 7 1 15 0 2 16 15 1 9 13 2 13 3 0 1 15 2 16 3 9 3 13 7 13 1 15 9 2 7 16 9 13 3 0 13 9 2 7 3 13 10 9 2 0 13 16 15 15 9 4 13 7 13 1 13 9 2
26 1 0 13 16 15 15 16 9 9 13 15 3 1 0 2 13 1 15 16 9 13 9 3 1 9 2
29 3 3 9 0 2 3 1 9 2 3 13 0 0 2 7 1 15 2 16 15 9 3 15 13 16 1 9 0 2
40 13 3 16 13 15 9 0 1 9 2 16 9 7 9 2 3 3 13 0 1 9 2 16 9 10 13 13 1 15 9 1 9 2 7 1 15 9 1 9 2
37 13 13 3 16 9 2 15 13 9 0 2 0 13 2 3 0 2 1 16 13 1 15 0 9 2 7 0 2 1 16 13 1 15 9 7 9 2
28 3 10 9 0 15 9 0 13 13 2 1 3 1 9 0 13 9 2 0 13 16 1 13 9 13 13 9 2
25 16 16 13 9 0 13 9 2 13 16 13 15 1 15 9 2 16 15 13 9 16 1 10 9 2
18 3 2 1 9 15 2 16 3 2 13 9 2 13 16 13 15 9 2
30 1 9 7 15 13 1 9 2 3 9 15 13 1 9 9 2 1 9 7 13 1 15 2 15 15 13 1 9 9 2
36 13 7 0 9 2 3 9 9 2 16 9 7 9 13 9 9 2 7 9 7 9 9 9 2 7 3 9 9 2 1 15 3 13 15 9 2
60 16 13 3 1 9 0 2 15 1 9 9 13 2 9 3 13 15 1 15 9 9 2 16 13 9 9 2 16 1 9 9 10 9 13 1 15 9 9 2 16 7 13 9 1 9 2 15 13 1 9 2 3 3 13 15 1 15 9 9 2
21 7 9 13 0 2 13 3 1 9 12 9 2 16 9 13 0 7 0 9 13 2
35 3 1 9 9 13 9 7 1 9 0 2 16 9 15 13 13 1 9 9 0 15 2 7 3 1 9 0 2 16 9 13 15 9 9 2
28 1 9 0 0 2 9 3 13 15 9 9 2 16 9 13 15 9 9 2 7 3 3 13 0 1 9 0 2
44 9 0 0 2 16 13 15 9 0 2 15 3 15 13 1 9 15 16 9 1 9 2 3 13 15 9 15 9 2 16 9 13 9 2 7 15 13 16 1 15 16 13 9 2
22 3 1 15 9 3 13 9 1 3 9 2 7 3 3 9 13 0 7 0 1 9 2
25 1 0 13 16 9 13 0 2 16 3 13 13 9 9 2 13 3 9 2 16 9 1 15 13 2
34 7 3 1 9 2 9 10 9 2 13 16 9 9 13 1 9 2 15 3 13 1 9 9 0 2 16 9 7 9 2 7 15 3 2
30 1 15 7 15 0 2 15 13 1 9 13 9 15 2 16 15 9 9 13 9 2 7 15 13 9 0 1 10 9 2
26 1 15 7 15 0 2 15 9 13 9 15 2 15 3 9 9 13 9 2 7 15 9 9 13 9 2
66 16 3 9 15 3 13 9 9 2 13 9 1 9 2 16 9 1 3 9 2 3 16 9 13 9 1 15 15 13 1 9 9 2 16 13 9 2 7 1 15 15 13 1 9 2 16 7 9 9 13 9 1 15 16 13 15 9 2 3 1 15 16 13 3 9 2
28 1 0 13 16 0 15 15 13 1 9 9 3 9 1 9 2 0 13 1 15 2 16 10 9 13 1 9 2
19 7 0 15 15 13 1 9 9 3 13 1 9 2 13 1 15 0 13 2
36 16 7 13 12 7 15 9 2 15 13 9 0 9 2 7 15 13 9 13 2 13 13 1 15 9 7 9 0 13 2 7 9 1 15 13 2
22 0 2 16 9 9 13 15 9 15 2 16 1 13 4 2 15 15 9 13 13 13 2
13 3 13 3 15 9 13 13 9 13 13 9 9 2
34 7 15 15 9 1 15 9 13 13 13 2 16 10 9 13 4 13 1 15 9 7 9 2 7 9 2 7 15 9 2 7 15 3 2
45 3 2 16 15 9 0 15 3 13 10 9 2 13 9 1 15 9 15 13 15 9 7 13 15 1 9 2 3 0 9 13 9 13 16 13 1 9 2 1 15 13 9 1 9 2
37 1 0 13 16 1 9 0 3 13 9 9 2 7 15 9 1 9 13 2 13 9 1 15 9 9 2 16 1 9 0 0 1 9 0 0 13 2
30 15 3 15 3 13 9 16 1 9 0 2 13 13 15 0 2 15 16 9 10 2 1 15 13 2 13 9 15 9 2
22 16 3 13 9 13 9 1 9 2 3 13 9 1 15 2 7 13 15 9 1 15 2
40 7 3 2 1 9 13 1 10 9 13 4 13 9 9 7 9 9 1 9 2 1 9 9 15 2 13 1 9 13 16 13 9 13 0 2 7 9 13 0 2
42 13 13 16 10 15 13 1 15 15 13 10 9 2 13 16 13 15 9 15 13 1 10 9 2 16 2 16 9 13 13 9 9 2 13 16 13 15 9 1 15 9 2
18 1 7 15 9 13 13 9 1 9 2 15 9 9 13 9 0 9 2
17 1 0 13 16 9 1 9 9 3 13 13 0 16 13 9 9 2
35 9 7 10 2 16 1 15 9 13 2 13 9 1 9 0 2 3 0 3 13 15 16 15 13 9 1 9 2 7 15 1 3 13 13 2
16 13 3 9 2 1 9 1 8 2 16 9 3 13 0 9 2
12 9 7 0 13 0 9 2 16 1 13 4 2
31 1 0 3 13 16 9 1 9 0 13 3 13 2 16 13 1 15 15 13 2 13 3 1 15 13 2 16 13 16 13 2
38 9 7 1 15 3 13 15 0 0 2 7 3 15 15 13 2 3 13 16 10 9 1 15 13 1 13 15 0 0 2 13 1 9 2 16 13 9 2
29 15 7 13 1 13 9 0 2 13 15 3 16 0 2 7 16 15 15 13 2 16 9 13 16 15 15 13 0 2
21 1 0 13 16 13 9 1 9 2 13 13 9 1 9 7 9 13 1 15 13 2
56 3 15 9 3 15 13 2 7 13 15 0 2 16 9 15 13 2 3 3 3 16 13 15 16 15 15 9 7 9 2 7 16 13 9 2 1 15 9 9 13 2 15 3 0 9 9 13 2 16 9 9 9 13 9 0 2
53 16 10 9 3 13 9 9 13 2 13 9 9 3 1 15 9 2 7 13 2 3 16 15 13 7 0 13 1 9 2 1 9 13 0 7 15 9 2 16 9 1 12 9 2 0 7 0 9 1 15 9 13 2
61 1 13 7 15 9 0 13 0 2 13 13 16 10 9 1 9 0 13 2 1 15 13 2 0 13 0 2 7 1 9 7 1 9 3 2 16 9 0 0 13 0 1 9 7 9 2 9 7 9 3 13 0 0 1 9 2 7 1 9 3 2
36 9 0 15 3 13 1 15 9 2 7 1 15 2 16 3 13 9 0 2 2 16 13 1 16 13 1 15 2 3 13 13 7 9 7 9 2
42 7 16 9 0 1 15 0 3 13 13 1 16 13 2 7 13 15 1 9 9 13 13 9 1 9 2 3 2 16 13 4 2 13 15 9 9 13 9 1 15 9 2
10 3 3 13 9 15 2 7 15 9 2
40 3 2 1 9 9 13 15 15 9 2 7 15 15 15 13 2 16 1 13 4 2 0 13 16 1 15 9 15 0 0 13 9 2 15 3 13 1 10 9 2
18 3 2 9 13 2 1 9 1 8 2 16 9 0 9 13 3 13 2
12 7 9 0 13 9 0 2 16 1 13 4 2
57 7 7 1 9 1 15 15 13 1 15 2 15 15 9 13 2 16 9 15 15 13 1 9 9 2 13 1 9 9 2 15 0 13 1 9 9 2 13 1 9 9 1 9 13 2 1 16 13 16 9 13 0 2 7 9 0 2
39 1 0 13 16 9 10 3 13 9 0 0 1 16 1 15 13 2 13 2 7 13 15 1 9 9 2 1 15 13 15 15 13 2 7 13 15 15 13 2
14 7 3 13 9 0 1 9 9 2 7 13 15 15 2
42 1 15 9 2 13 13 16 13 1 3 13 1 15 13 2 16 3 13 15 13 16 9 10 3 2 7 13 13 4 13 9 3 9 15 2 3 9 13 13 1 13 2
7 9 7 9 13 1 9 2
21 3 7 1 13 16 9 2 1 16 13 3 0 2 1 15 3 13 1 15 9 2
26 9 3 2 16 13 9 13 15 9 2 3 1 15 13 2 16 0 1 15 13 9 2 1 15 13 2
26 1 0 13 16 9 0 3 13 9 0 2 15 13 1 9 2 16 1 16 4 13 1 9 1 9 2
43 16 3 1 13 4 2 13 3 13 9 13 1 15 0 2 7 13 1 13 16 9 7 9 15 2 16 9 13 9 13 2 16 3 9 13 9 2 3 13 13 9 0 2
18 1 9 7 3 13 9 15 13 15 16 10 9 2 16 1 13 4 2
49 1 0 13 16 13 13 9 13 3 3 1 10 9 2 7 1 10 9 2 1 15 13 1 9 2 16 9 7 9 15 2 9 3 3 13 1 9 2 7 9 15 2 16 13 1 12 1 9 2
33 3 3 15 13 13 1 9 10 2 16 9 0 13 9 0 9 2 3 10 9 13 1 9 15 13 9 9 2 16 9 1 9 2
15 3 1 15 9 0 13 0 9 2 15 13 9 1 9 2
17 7 10 9 2 1 15 15 9 1 0 9 13 2 9 15 13 2
30 9 7 9 13 9 9 2 15 16 9 13 1 10 9 2 3 13 16 9 9 13 9 9 2 16 9 13 9 9 2
22 7 13 13 16 9 0 2 16 13 9 13 1 15 15 13 9 2 3 13 9 9 2
27 7 0 9 0 3 13 9 9 1 16 13 3 1 13 2 16 13 15 9 1 9 2 15 13 1 9 2
34 1 3 9 0 1 13 15 13 2 1 13 15 9 13 2 2 3 13 13 9 2 16 13 1 12 1 9 2 16 13 1 12 8 2
35 15 13 1 15 2 16 9 0 7 0 3 13 9 1 9 10 2 7 1 9 3 2 3 16 13 9 1 9 10 2 3 1 9 13 2
25 16 0 1 9 0 13 15 9 7 9 2 15 2 15 1 3 13 2 3 13 16 1 9 0 2
45 3 2 1 9 0 9 15 13 3 0 1 9 2 1 15 13 9 0 2 7 3 1 1 9 2 16 1 13 2 0 13 16 9 9 1 1 0 15 13 2 15 1 9 13 2
18 7 13 0 1 9 9 2 16 13 0 15 9 2 7 3 9 3 2
19 15 7 3 13 2 16 9 15 13 15 13 1 9 9 15 13 9 9 2
16 7 13 15 2 13 16 15 9 13 9 1 9 0 1 9 2
13 1 9 7 0 1 9 2 3 13 9 13 9 2
34 15 16 13 0 9 0 13 2 7 3 1 16 0 13 2 0 3 13 15 1 9 9 1 9 2 3 1 9 9 1 9 0 0 2
21 9 3 9 2 0 9 13 2 3 1 9 13 9 15 9 2 1 15 9 13 2
38 9 7 15 9 1 15 13 2 1 12 13 13 2 7 16 13 9 15 15 13 9 2 7 16 13 9 9 15 2 1 16 9 0 13 13 1 13 2
17 1 10 3 15 3 1 9 13 2 0 13 9 13 9 9 15 2
15 9 7 3 13 1 9 2 16 16 9 9 13 1 15 2
20 1 15 3 9 13 9 9 13 1 9 0 2 16 1 15 15 13 1 9 2
17 7 15 13 13 9 9 2 16 9 13 9 13 9 15 9 13 2
37 16 3 9 3 4 9 13 2 7 4 13 1 9 1 9 13 2 16 1 13 2 0 13 16 1 9 0 13 9 2 1 9 15 9 4 13 2
47 7 1 13 15 13 9 2 1 9 12 12 8 2 9 13 0 15 9 7 9 9 0 7 0 2 16 15 13 3 13 2 7 1 15 0 7 3 15 9 15 13 2 15 0 9 13 2
40 15 7 3 0 9 3 13 2 0 13 13 2 16 15 13 9 13 13 1 9 13 16 15 13 2 3 7 16 9 15 13 2 15 13 9 13 9 1 9 2
20 9 3 9 1 9 9 13 15 1 15 13 2 1 15 9 9 1 9 13 2
38 16 9 2 16 13 9 9 1 9 2 13 13 9 2 16 7 13 9 9 16 1 15 13 2 1 15 16 13 15 13 15 2 13 9 7 9 9 2
18 3 2 9 13 9 0 2 15 3 13 13 9 2 1 15 13 9 2
28 7 16 15 13 9 13 1 9 2 3 3 1 9 2 13 3 9 9 1 9 2 3 3 15 1 9 9 2
34 9 3 1 9 9 13 10 9 15 1 9 13 9 2 7 15 15 13 9 3 13 2 16 9 7 15 15 2 13 1 15 15 9 2
29 7 3 13 16 9 0 13 0 1 9 1 9 10 2 13 3 9 0 2 15 13 9 9 15 13 1 9 9 2
39 1 7 10 9 13 0 1 16 13 0 9 9 10 2 0 13 16 9 2 16 13 13 2 13 0 16 13 9 9 13 2 15 13 9 15 16 13 13 2
22 7 16 13 9 3 15 13 16 13 9 15 1 9 13 2 3 0 13 7 13 0 2
30 7 15 13 13 7 13 2 3 1 10 9 15 9 13 1 13 2 7 13 15 9 13 1 9 2 7 13 1 15 2
25 7 3 2 16 0 13 9 7 9 9 2 3 12 13 9 0 9 2 1 15 10 9 13 0 2
45 15 9 2 16 3 13 1 15 15 13 1 15 9 7 9 2 16 9 0 13 13 12 2 3 16 13 12 9 2 16 9 13 12 1 9 12 9 2 7 1 9 10 9 13 2
7 3 3 9 0 13 13 2
30 13 3 9 0 0 0 7 1 15 2 16 13 1 9 9 2 3 13 15 9 9 0 13 2 16 13 1 9 9 2
48 7 1 0 0 9 3 13 0 9 2 16 1 9 2 7 16 1 0 2 1 15 3 16 2 1 9 9 2 3 13 13 9 0 2 16 7 15 0 2 1 10 9 2 13 13 9 9 2
22 13 13 16 2 16 9 13 9 1 0 9 2 3 9 0 13 13 1 9 9 13 2
58 3 2 16 9 0 3 13 1 9 15 15 13 1 10 9 2 13 7 13 1 15 0 7 13 2 16 9 1 15 15 13 13 12 9 2 3 7 1 15 15 13 13 9 2 3 9 0 3 13 1 13 9 15 9 15 9 13 2
39 7 3 2 9 0 7 0 13 1 9 0 2 7 13 2 15 13 9 2 7 13 13 2 16 13 1 12 8 2 7 3 3 13 15 2 16 9 13 2
10 9 0 0 13 15 1 10 9 13 2
22 7 15 3 13 1 15 9 2 15 3 13 1 9 10 9 2 7 1 9 0 9 2
46 13 3 15 2 15 13 15 2 3 13 9 1 9 7 9 2 15 13 15 1 9 2 7 0 3 1 9 9 2 7 9 1 15 13 2 7 9 1 15 13 2 13 15 1 9 2
20 7 3 13 9 2 15 1 9 13 15 1 9 2 13 15 1 9 7 9 2
29 15 0 0 13 15 2 3 0 13 9 1 9 9 2 7 3 3 1 9 15 13 9 9 2 15 1 15 13 2
20 7 3 13 9 2 15 9 9 13 9 3 1 9 13 2 7 1 9 13 2
46 7 16 3 9 9 15 13 9 9 2 1 9 13 2 3 3 1 15 13 15 9 10 9 2 7 10 9 2 7 4 15 13 1 9 2 15 9 1 15 13 13 1 9 9 13 2
38 16 3 1 9 2 13 16 9 1 15 13 9 9 2 3 9 0 2 13 15 15 13 9 9 2 7 15 13 15 15 13 9 3 2 1 13 9 2
18 1 0 13 16 13 13 13 9 1 9 9 2 3 7 1 9 13 2
39 3 15 9 9 13 3 9 1 9 7 1 13 2 16 9 9 1 9 9 13 9 0 7 0 2 1 9 7 15 13 1 9 2 13 9 0 7 0 2
36 1 0 13 16 2 16 1 9 9 0 3 13 9 2 7 3 9 2 10 9 0 9 13 9 0 1 9 0 1 10 9 2 16 1 15 2
21 16 3 9 0 13 9 1 9 1 10 9 2 3 9 13 9 1 10 9 0 2
21 15 7 9 1 10 9 0 15 13 9 2 16 16 3 13 15 2 13 1 15 2
26 3 7 9 0 1 9 13 1 9 0 2 0 9 13 2 16 3 2 1 13 15 2 13 1 15 2
54 1 0 13 16 12 7 15 9 2 3 1 15 2 13 9 9 16 13 2 15 13 9 9 2 7 9 16 13 2 16 9 2 16 13 1 9 3 2 3 13 1 15 16 13 7 3 13 1 9 2 16 1 9 2
29 1 15 9 2 13 4 16 2 1 9 13 9 1 10 9 2 15 9 13 1 9 13 2 15 13 1 9 0 2
45 1 9 7 3 13 16 2 16 15 13 13 1 15 9 0 2 3 1 9 0 15 13 13 2 13 3 13 15 15 3 13 9 7 0 2 3 7 13 13 15 15 3 13 9 2
27 3 3 9 0 13 9 7 9 2 7 9 2 15 13 9 15 9 2 7 9 12 2 15 13 9 15 2
48 16 3 1 9 0 13 13 9 2 1 0 9 15 13 1 15 0 2 3 12 9 15 4 1 9 9 2 7 15 1 9 9 2 1 9 1 9 13 2 16 3 13 9 9 1 9 0 2
21 7 3 15 9 9 13 1 15 9 2 7 15 1 15 2 13 1 0 0 9 2
29 3 2 1 9 2 1 12 8 2 15 9 0 13 15 9 2 3 9 13 0 16 9 2 7 9 16 9 0 2
25 1 10 3 9 15 13 2 16 3 15 9 9 13 9 15 13 2 3 13 0 15 9 1 13 2
19 1 0 3 13 16 9 13 1 0 15 13 1 9 9 3 13 1 9 2
53 1 0 13 16 2 16 0 9 3 13 15 13 2 7 3 13 3 13 2 13 3 13 9 0 9 0 2 13 16 15 13 2 9 13 9 0 2 0 7 0 2 9 3 0 13 9 9 0 2 7 13 15 2
17 7 16 3 9 13 0 7 0 2 0 3 9 7 9 13 9 2
22 7 16 1 9 13 9 15 9 2 0 9 15 9 2 15 13 15 9 2 13 9 2
29 3 9 1 15 9 13 16 9 13 15 13 0 9 2 0 3 9 13 15 13 9 2 7 13 1 0 9 9 2
25 3 2 9 13 2 1 9 9 2 16 9 2 15 13 15 16 9 2 13 9 1 9 7 9 2
21 15 7 15 13 13 1 9 7 9 2 13 9 9 2 15 7 9 7 9 13 2
23 3 2 9 13 2 1 9 9 2 16 9 13 9 2 9 7 2 3 9 2 13 9 2
9 7 7 9 7 9 13 13 9 2
32 3 1 9 13 1 9 7 9 2 9 13 3 0 9 2 7 0 9 2 7 9 1 9 7 9 0 2 16 13 9 9 2
42 7 9 1 15 9 7 1 15 9 2 13 9 9 7 9 2 9 3 7 9 7 9 13 1 9 9 2 7 15 9 7 15 9 7 15 9 13 1 9 15 9 2
23 7 13 15 1 9 1 9 1 9 7 9 2 16 1 13 4 2 1 1 9 0 13 2
20 1 0 13 16 9 13 1 9 7 9 2 13 16 13 9 2 1 9 9 2
17 3 7 9 13 2 1 9 1 8 2 9 0 9 13 3 13 2
30 7 16 1 15 13 2 13 1 9 10 9 2 15 3 13 9 0 2 7 13 9 0 9 2 16 3 9 13 13 2
27 1 15 3 9 13 9 2 7 9 2 7 9 2 9 2 16 9 13 9 13 2 7 9 13 9 13 2
39 15 13 9 0 2 15 13 1 13 7 0 9 2 7 15 9 13 9 15 3 13 1 15 9 2 7 13 1 13 2 1 16 9 13 1 12 7 0 2
9 1 0 13 16 9 13 9 9 2
24 13 7 3 12 9 1 0 2 16 13 1 15 15 13 8 12 2 15 1 1 9 9 13 2
34 13 3 9 9 9 1 0 9 2 1 16 9 0 13 1 9 9 2 3 13 16 3 13 1 3 9 1 9 2 7 1 13 9 2
33 16 16 13 1 9 9 2 3 13 0 2 16 13 9 2 0 9 13 9 2 3 2 15 1 15 15 15 13 9 2 13 9 2
22 1 15 2 1 13 0 9 2 9 0 13 2 1 13 0 9 0 2 13 9 9 2
15 0 13 3 16 9 13 9 1 9 2 15 13 9 13 2
37 7 3 15 13 0 9 13 2 3 0 7 9 13 9 2 16 9 0 13 9 16 3 0 2 3 1 9 13 13 2 16 13 15 0 1 9 2
46 3 15 15 16 1 9 0 13 15 9 9 13 7 13 2 1 9 7 13 3 13 15 9 2 7 9 3 2 13 16 9 2 7 1 13 9 2 1 0 13 1 9 16 1 9 2
55 9 3 9 9 9 0 3 13 2 13 3 9 2 12 1 8 2 3 13 15 9 9 2 16 9 3 13 2 16 15 13 3 0 13 1 9 2 15 3 13 9 16 9 13 2 15 7 13 13 2 7 0 3 13 2
17 1 8 9 3 1 9 9 13 2 3 13 2 7 9 9 13 2
36 3 13 13 0 9 13 1 9 13 2 1 15 15 9 9 13 2 7 0 9 15 1 9 10 2 16 9 10 13 1 9 1 9 9 13 2
11 7 9 2 7 9 2 1 0 13 0 2
22 1 0 13 16 9 2 16 13 1 9 1 9 9 2 13 9 13 1 15 1 15 2
25 15 3 9 9 13 13 9 15 2 16 15 15 13 15 2 13 9 15 2 16 13 9 15 0 2
12 3 9 13 1 9 13 2 16 7 15 0 2
34 16 3 9 7 9 13 12 9 2 1 9 9 13 1 15 9 9 2 3 13 12 9 9 0 2 1 9 9 13 1 15 9 9 2
28 1 0 13 16 2 1 13 2 9 7 9 13 12 9 9 0 2 13 12 9 2 15 13 9 13 1 9 2
17 3 0 9 13 9 1 9 2 0 0 1 15 2 1 9 13 2
41 3 1 15 9 2 13 13 16 2 1 9 0 13 1 10 9 2 16 0 1 9 2 7 9 1 9 2 10 15 1 15 15 13 2 3 1 15 13 9 9 2
22 16 16 13 2 15 13 13 9 2 15 0 13 1 9 9 0 2 16 3 13 9 2
47 13 3 16 9 13 13 9 2 16 9 3 13 9 2 15 13 9 9 2 7 9 1 9 13 2 7 13 16 9 13 13 9 2 16 9 3 13 9 9 2 7 15 9 1 15 13 2
32 7 3 9 15 13 16 9 2 9 7 16 9 9 2 1 15 3 1 0 2 3 1 9 13 2 9 13 16 9 12 9 2
13 13 7 1 9 13 9 15 13 15 15 13 9 2
36 9 7 13 9 3 13 13 9 2 16 1 9 15 9 2 15 13 15 9 2 16 1 13 2 15 9 13 0 9 2 15 9 13 9 9 2
36 7 0 2 16 1 0 2 13 9 2 3 13 9 2 13 12 9 13 12 9 2 7 12 9 12 9 2 16 13 15 0 13 1 9 9 2
21 1 0 13 16 9 2 0 13 2 13 13 16 15 15 13 9 2 16 9 9 2
22 1 0 7 2 9 13 9 15 3 13 13 16 15 2 16 1 13 13 7 13 9 2
49 7 3 13 12 0 2 15 12 13 9 2 7 15 9 9 2 16 16 13 2 9 13 0 9 2 7 3 13 12 0 13 9 12 0 2 16 1 13 2 9 9 13 15 2 3 9 0 9 2
15 16 3 9 0 13 16 9 9 9 2 13 9 9 13 2
13 15 3 13 10 9 2 16 13 1 10 9 0 2
36 7 3 1 15 16 13 12 9 12 9 2 13 9 1 9 9 2 3 13 15 13 9 16 9 2 15 13 2 16 13 12 9 1 15 9 2
31 9 7 2 16 1 15 13 9 2 3 1 15 13 9 7 9 2 3 7 9 7 9 9 0 13 1 9 13 1 9 2
19 1 9 7 3 13 12 9 1 0 9 16 9 9 2 16 9 9 13 2
22 3 9 13 15 9 2 16 13 0 2 13 1 0 1 0 2 3 7 16 13 9 2
26 1 0 7 9 0 13 1 9 9 2 16 13 4 15 3 0 13 7 0 12 2 16 1 13 4 2
20 1 0 13 16 9 13 1 15 9 9 2 3 13 9 7 9 2 7 9 2
29 3 3 15 9 9 13 1 9 2 16 1 13 2 9 13 2 16 15 9 13 9 9 9 13 2 15 13 9 2
39 1 0 3 13 16 15 9 9 2 16 13 1 9 0 1 15 2 16 9 13 3 13 2 13 3 1 9 0 1 15 2 16 9 13 13 1 0 9 2
24 16 3 9 13 1 15 9 9 2 3 9 2 0 13 1 0 9 2 1 15 13 1 9 2
19 7 9 13 1 15 9 9 2 3 9 0 2 13 12 7 0 1 9 2
22 7 15 9 9 3 13 1 9 10 9 16 13 1 9 2 16 13 9 16 9 0 2
21 1 0 13 16 9 2 16 13 12 1 0 9 2 13 15 9 1 9 9 0 2
14 3 2 0 9 2 1 0 13 2 13 1 9 9 2
23 7 12 9 3 15 13 1 15 16 9 2 1 9 1 15 15 13 9 2 13 3 13 2
29 1 0 13 16 2 16 3 13 0 9 9 2 16 13 15 0 2 13 16 12 9 15 13 1 15 1 9 9 2
10 3 0 13 9 9 1 15 9 13 2
11 15 3 13 1 0 2 16 15 9 9 2
29 3 2 1 1 9 9 13 2 16 13 1 15 15 13 9 2 13 13 9 13 1 9 2 7 15 3 13 9 2
25 16 3 0 9 13 9 9 7 9 2 13 16 1 0 15 13 0 7 9 2 16 9 7 9 2
26 1 9 7 13 13 1 9 9 2 3 3 1 9 3 2 7 3 1 9 13 2 16 9 1 9 2
12 9 7 3 13 16 9 2 7 16 9 9 2
20 3 2 15 9 13 16 1 10 9 2 3 3 0 1 0 13 16 1 9 2
9 9 0 1 9 9 2 16 9 2
34 0 3 2 16 1 15 16 15 12 13 13 2 0 13 15 9 13 1 15 0 15 2 16 1 9 13 7 1 9 2 7 1 9 2
21 15 0 2 1 16 9 13 1 9 2 16 9 9 13 1 9 1 10 9 0 2
34 1 9 0 15 13 1 9 7 9 2 15 13 1 9 2 13 3 9 9 1 9 2 13 3 1 9 10 7 9 9 7 9 9 2
31 16 7 1 0 3 13 0 7 0 2 7 9 7 9 2 1 9 2 3 2 1 9 13 2 13 15 9 15 1 0 2
40 16 0 13 1 9 9 9 1 9 2 13 9 3 0 2 13 9 9 7 9 2 16 2 13 1 9 1 9 16 13 0 7 13 2 13 9 7 9 9 2
47 3 3 9 0 3 13 13 9 0 2 16 9 9 13 2 7 13 15 10 9 2 16 13 15 9 0 2 16 9 13 15 9 2 9 3 13 15 13 1 0 2 1 9 13 9 9 2
13 15 9 13 2 16 9 13 9 9 1 15 13 2
27 0 13 7 16 12 9 3 13 16 12 9 0 2 1 15 9 13 9 2 3 15 15 13 2 15 13 2
44 7 9 1 15 9 13 2 3 13 12 3 2 7 13 0 2 1 16 13 0 9 13 2 3 15 9 13 2 3 13 15 15 13 9 2 7 15 13 7 13 15 9 13 2
18 15 3 13 1 9 2 13 1 9 15 1 15 13 2 1 15 9 2
12 0 7 9 3 13 0 2 7 15 9 0 2
62 13 7 13 16 15 13 1 15 2 15 9 15 13 16 9 0 2 7 15 13 9 0 2 16 9 13 13 1 9 2 7 13 9 0 2 16 9 13 13 1 9 2 7 13 9 0 2 1 15 3 1 15 15 9 13 0 2 7 3 13 15 2
33 10 7 13 15 1 10 9 2 13 15 0 3 1 9 15 13 16 9 13 13 0 13 1 9 0 2 15 9 9 13 13 9 2
27 16 3 9 16 9 9 13 2 13 3 9 0 2 13 15 1 9 9 2 16 9 0 1 15 9 13 2
24 9 7 0 2 1 9 13 2 13 9 13 2 3 7 13 15 13 13 2 3 9 13 9 2
27 15 3 13 3 13 16 1 0 9 9 2 9 3 12 9 3 13 16 1 9 2 15 1 0 3 13 2
7 9 7 13 1 9 9 2
11 9 7 1 9 3 13 9 2 7 9 2
37 7 15 13 9 9 2 15 13 1 9 15 9 7 9 2 15 3 9 13 1 16 13 15 3 7 0 0 2 16 13 9 7 0 9 1 9 2
34 3 7 9 0 13 0 3 1 9 2 3 1 15 9 9 7 9 2 7 3 13 9 0 2 16 13 0 9 1 10 9 7 9 2
9 0 7 13 9 0 1 9 9 2
16 0 7 9 9 13 9 2 3 10 9 13 9 1 10 9 2
14 0 7 9 13 9 2 3 10 9 13 1 10 9 2
41 15 3 13 1 12 9 2 13 13 0 2 16 0 15 9 13 2 16 16 13 9 13 0 9 1 9 2 7 3 13 13 0 2 16 12 15 9 9 15 13 2
28 13 3 13 0 9 2 16 13 9 9 2 7 3 1 0 2 16 9 0 13 1 9 2 7 0 1 13 2
39 1 9 3 0 2 1 9 9 2 16 3 1 9 0 9 13 13 9 15 9 13 2 16 1 13 4 2 3 1 15 9 13 13 9 1 15 9 13 2
28 1 0 13 16 9 13 1 9 0 9 0 2 16 9 9 13 1 9 9 2 1 15 9 1 9 1 0 2
39 16 2 16 9 13 2 12 1 8 2 9 0 3 4 13 0 9 1 9 0 2 7 1 9 1 0 9 9 2 9 0 15 7 9 9 13 15 13 2
27 0 0 13 2 13 1 9 1 9 0 7 9 2 15 13 0 2 7 13 9 13 1 9 1 9 0 2
12 7 13 13 16 9 1 9 13 1 13 9 2
47 15 3 15 13 9 9 16 13 9 2 13 13 9 9 2 3 0 1 16 13 15 1 9 0 2 7 1 16 13 15 1 9 0 2 7 3 1 10 15 15 13 1 9 15 15 9 2
38 1 0 3 13 16 9 1 12 8 13 1 13 0 2 15 13 1 9 1 9 2 7 0 7 0 3 7 13 1 9 1 9 15 1 0 9 13 2
22 1 0 13 16 9 15 3 13 16 9 3 4 13 2 7 16 3 4 13 1 9 2
21 7 9 2 1 15 9 9 12 12 8 13 2 13 9 0 2 15 0 9 13 2
52 1 15 9 2 13 13 16 1 9 15 9 3 0 13 9 2 16 9 13 9 13 2 9 3 13 13 9 1 9 2 1 9 1 15 13 2 7 15 13 9 1 15 1 13 2 7 13 9 0 9 13 2
13 0 13 7 16 15 15 0 13 2 13 9 13 2
28 15 7 9 9 13 16 13 2 16 1 0 9 2 1 0 9 2 15 9 0 13 2 15 1 9 9 13 2
27 7 3 13 13 16 1 0 9 13 9 10 9 2 15 1 13 9 2 15 13 9 0 1 9 0 13 2
28 3 2 9 9 7 9 13 7 9 3 13 1 15 9 2 16 13 1 12 8 2 16 9 9 13 9 13 2
23 1 0 13 16 9 13 3 13 9 9 16 16 13 9 9 13 2 15 10 9 13 13 2
17 3 9 13 13 0 13 2 1 9 13 0 15 15 13 1 9 2
47 16 9 0 13 0 7 0 16 9 2 1 15 16 9 0 13 0 16 9 0 2 3 9 0 9 2 15 13 9 1 15 1 9 2 13 0 16 0 2 15 13 9 1 15 1 9 2
15 7 7 15 9 13 9 0 3 1 9 2 7 13 9 2
18 7 1 2 0 13 13 15 1 15 9 2 16 1 9 0 7 0 2
21 7 9 0 7 1 15 2 15 13 15 1 9 0 7 0 2 13 15 1 13 2
22 9 7 7 9 2 7 15 3 2 3 13 9 16 15 13 2 7 16 15 15 13 2
27 16 3 9 7 9 2 7 3 2 15 3 13 2 3 13 13 16 13 2 3 3 13 13 13 16 13 2
27 3 3 13 16 9 2 13 9 2 15 13 1 9 10 9 2 13 9 9 2 15 13 9 0 0 9 2
30 1 9 7 0 3 13 13 15 1 15 13 15 2 16 13 15 1 10 9 2 1 15 13 9 2 1 13 9 0 2
44 0 3 13 9 2 16 13 9 1 9 1 15 13 13 9 2 16 9 13 13 9 9 1 9 15 0 2 7 13 1 9 7 9 0 2 15 3 13 9 16 13 1 9 2
26 3 15 9 13 0 9 9 2 3 7 9 15 2 16 9 13 9 2 7 15 9 13 13 9 9 2
28 15 7 9 13 9 3 1 9 9 15 2 16 9 13 9 13 2 7 9 9 9 2 7 15 13 9 9 2
24 15 3 9 13 1 10 9 2 7 13 9 1 15 13 1 9 2 7 13 9 1 15 15 2
21 1 7 16 13 15 9 7 9 2 13 9 2 1 16 9 9 13 1 9 9 2
33 7 15 15 13 1 9 12 12 8 15 13 2 15 13 2 15 13 2 13 3 15 1 10 9 2 13 1 9 2 13 1 9 2
11 1 15 3 9 9 7 9 13 15 9 2
19 7 1 9 0 3 13 15 9 16 9 0 2 15 13 9 0 7 0 2
9 3 3 1 9 9 13 9 0 2
12 3 15 9 3 13 1 9 2 7 1 9 2
9 13 13 16 15 9 13 1 9 2
19 15 15 13 3 13 1 9 9 2 7 0 1 9 13 2 13 9 9 2
30 7 15 13 15 1 9 9 2 16 13 13 1 9 7 9 2 16 3 9 13 1 9 1 9 2 13 15 0 13 2
15 15 0 13 9 13 7 13 1 9 13 2 1 9 9 2
8 7 15 13 15 1 9 9 2
46 3 3 13 16 9 0 9 3 13 0 2 7 15 15 13 2 7 3 2 1 13 7 13 3 13 0 16 9 0 2 16 1 13 4 2 9 3 13 13 7 13 2 7 13 13 2
26 1 0 3 13 16 9 13 13 1 9 2 9 13 2 3 16 15 13 1 15 2 7 1 9 3 2
14 1 0 13 16 9 0 1 9 13 1 9 9 0 2
39 1 0 13 16 1 9 9 0 13 9 0 2 15 13 9 0 2 15 13 3 1 9 2 7 1 9 15 2 7 13 13 16 15 9 13 1 9 13 2
31 7 15 0 13 13 2 13 9 2 15 13 1 9 1 9 2 15 13 1 9 2 7 1 3 9 2 15 13 1 9 2
17 7 3 13 13 9 1 9 2 9 7 9 1 9 2 13 9 2
21 16 9 0 13 9 2 7 13 9 2 3 13 16 9 13 1 9 1 13 9 2
22 3 0 1 15 13 16 13 9 1 15 9 7 3 1 15 2 1 9 9 1 9 2
30 7 15 3 0 13 1 9 2 15 3 13 9 7 9 2 7 13 0 1 15 2 16 15 13 9 0 9 7 9 2
36 1 0 13 16 2 16 9 13 1 9 13 0 1 9 10 9 2 3 13 1 9 1 9 1 9 1 15 13 7 13 2 16 1 0 13 2
18 1 0 13 16 2 13 9 2 13 9 1 9 9 15 13 9 9 2
20 1 13 7 1 9 2 15 13 4 7 13 2 13 16 9 15 13 9 9 2
13 0 2 16 9 13 1 9 2 7 3 1 0 2
8 9 7 9 13 1 9 0 2
25 3 3 9 13 1 9 1 9 2 7 0 1 0 1 9 13 4 9 2 16 13 0 9 13 2
28 1 0 3 13 16 9 1 9 13 1 9 1 15 13 2 15 12 3 13 12 2 7 3 3 13 16 12 2
18 9 7 0 2 15 13 9 2 16 1 13 4 2 13 1 9 13 2
13 1 7 9 13 1 9 2 9 0 13 1 0 2
31 9 7 0 3 13 9 2 16 2 16 13 1 12 8 2 9 9 13 16 9 2 1 15 9 13 1 9 7 9 9 2
26 3 2 10 15 13 9 1 9 2 13 13 1 9 2 13 15 9 2 16 9 1 9 13 1 9 2
27 7 9 13 9 1 9 2 16 3 1 13 9 2 13 9 2 1 7 13 15 9 2 13 9 1 9 2
20 3 2 1 13 9 2 13 9 2 1 7 13 15 9 2 13 9 1 9 2
16 3 3 13 13 16 9 13 15 9 2 7 15 9 7 9 2
34 7 1 3 9 7 9 13 9 2 3 0 2 7 0 2 16 16 10 9 13 9 9 2 3 10 9 2 16 3 2 13 9 9 2
31 7 3 9 13 9 13 9 1 0 2 16 1 16 13 9 0 2 16 7 1 0 13 9 9 0 2 16 13 15 9 2
44 15 7 12 9 9 3 13 15 1 15 2 3 1 16 13 9 15 2 7 1 16 15 9 13 2 3 10 9 13 1 15 9 2 7 10 15 13 16 9 2 13 9 15 2
58 9 7 9 7 9 13 12 7 15 2 3 9 1 9 2 7 13 9 1 9 0 2 16 9 0 2 15 13 9 9 0 7 9 13 2 7 13 9 1 9 1 15 7 1 9 0 2 16 9 0 2 15 13 9 9 7 9 2
30 0 13 7 16 9 1 15 15 13 9 2 9 15 13 2 7 9 15 2 7 3 10 9 1 9 2 9 15 13 2
28 9 7 15 9 3 13 13 1 9 2 16 13 9 1 9 2 7 1 9 2 16 13 9 1 9 7 9 2
28 13 3 3 9 1 9 15 9 13 1 9 2 15 3 3 13 1 9 2 3 0 13 1 13 9 7 9 2
31 16 13 1 9 0 7 0 9 2 9 3 7 9 2 1 15 13 7 13 9 9 1 9 9 2 3 13 13 1 0 2
15 9 3 0 13 9 7 9 9 2 9 7 0 13 9 2
17 12 9 2 1 9 9 2 7 15 9 2 15 13 1 9 9 2
15 9 3 15 13 1 9 9 7 9 9 2 13 9 9 2
36 7 16 13 0 9 9 2 9 7 9 7 9 9 15 13 2 15 13 1 9 9 2 7 7 9 2 16 13 9 1 9 2 13 9 9 2
13 9 7 0 9 3 13 2 7 13 3 9 9 2
31 1 9 3 7 9 9 2 16 1 9 13 1 9 13 1 9 15 9 9 2 16 1 9 9 13 9 9 9 7 9 2
36 16 3 2 3 9 13 9 1 9 2 3 9 13 9 10 2 3 3 3 9 13 0 2 3 9 7 9 9 7 9 2 13 1 9 9 2
19 7 15 13 1 9 2 16 9 3 13 13 9 9 2 7 13 9 0 2
28 13 4 3 16 15 9 2 16 10 9 13 15 9 1 15 13 9 7 9 2 13 10 9 15 9 7 9 2
18 0 13 7 16 9 15 0 9 13 1 9 13 2 13 9 9 0 2
13 16 7 9 13 9 15 2 3 9 13 15 9 2
23 3 10 9 7 9 7 9 1 9 1 9 9 13 2 9 7 7 9 1 9 1 9 2
18 0 2 13 16 9 13 15 2 13 3 9 13 13 1 9 7 9 2
10 13 16 9 13 13 1 9 7 9 2
17 7 9 13 1 9 2 9 0 1 9 2 16 13 1 12 8 2
14 3 10 15 13 1 9 2 13 13 1 9 7 9 2
8 3 13 13 1 9 7 9 2
17 3 13 9 2 1 9 1 8 2 16 9 0 9 13 3 13 2
9 3 9 13 13 1 9 7 9 2
6 3 2 9 13 9 2
10 15 3 13 9 3 2 13 9 0 2
12 3 3 13 9 3 2 7 13 9 1 9 2
10 3 2 9 0 13 7 13 1 9 2
12 9 3 15 3 13 1 9 2 13 9 0 2
13 7 9 9 3 13 0 2 16 10 9 13 13 2
7 3 9 9 13 1 9 2
13 13 13 16 15 13 9 13 13 1 9 7 9 2
34 3 1 15 13 13 16 15 1 15 13 9 0 1 0 2 13 15 3 9 2 7 15 15 13 15 9 13 3 0 2 13 9 15 2
35 7 1 15 13 16 15 13 9 0 0 7 0 2 16 13 16 9 0 9 3 13 13 1 9 0 2 16 9 9 13 13 1 9 0 2
27 3 3 13 0 16 9 0 7 0 13 1 12 9 9 2 16 3 12 7 15 9 9 13 0 7 0 2
19 3 13 16 15 9 9 13 15 13 9 0 2 7 15 15 13 9 0 2
41 15 1 15 9 13 2 1 15 9 15 13 9 7 9 2 3 3 15 13 2 16 1 9 13 2 16 9 1 9 13 0 9 2 15 9 3 13 1 16 3 2
34 1 9 7 0 15 13 15 13 1 0 9 2 3 9 2 7 15 15 13 2 3 9 2 3 1 15 13 9 2 7 1 15 9 2
24 9 3 13 9 2 16 1 15 13 1 9 15 9 2 7 9 2 7 9 2 7 15 15 2
23 3 7 9 3 13 9 2 3 13 9 9 2 15 13 16 9 9 13 2 7 9 9 2
17 7 9 0 13 1 9 1 15 9 9 2 3 3 13 1 9 2
23 1 0 13 16 2 16 1 9 3 13 9 9 7 9 2 13 3 1 15 9 7 9 2
12 0 3 9 7 9 2 1 15 13 9 15 2
26 13 3 9 2 7 13 16 15 9 13 3 1 9 2 3 13 9 9 1 15 9 16 9 1 9 2
38 7 15 13 15 1 15 13 2 16 9 13 13 1 15 13 7 15 13 2 7 1 9 7 15 13 2 16 9 13 2 3 15 13 13 15 9 0 2
23 9 7 0 13 9 1 9 9 2 7 9 1 9 9 2 15 13 1 9 1 15 13 2
22 9 7 0 13 13 13 1 10 9 2 7 0 1 16 15 9 3 4 13 1 15 2
37 1 0 3 13 16 1 9 3 13 9 15 13 9 13 2 13 1 9 0 2 7 13 1 9 9 2 16 9 13 1 13 2 16 1 13 4 2
17 15 3 15 13 9 7 13 9 2 13 1 9 2 7 13 0 2
26 16 3 9 3 13 13 1 9 7 9 2 16 13 4 1 2 13 16 0 13 13 12 9 12 9 2
23 3 13 16 10 9 0 13 12 9 2 7 16 13 1 15 15 15 9 9 16 9 0 2
22 1 0 13 16 3 7 0 2 1 16 13 1 9 7 9 12 9 2 3 13 9 2
22 7 1 16 13 1 9 0 9 2 3 13 9 2 16 16 13 16 9 13 13 9 2
40 15 9 13 2 16 15 13 16 1 15 2 16 9 15 1 9 13 2 3 2 1 9 13 15 9 0 2 16 1 13 13 2 0 13 16 15 9 13 0 2
17 9 7 1 15 13 9 2 15 3 13 9 9 1 16 13 9 2
8 9 0 13 9 9 1 9 2
18 9 3 1 9 7 9 13 13 9 1 15 2 16 9 13 1 9 2
23 7 16 15 9 13 1 10 9 2 16 13 1 9 2 16 13 4 2 3 13 13 9 2
12 7 9 3 13 9 16 9 2 16 13 4 2
19 1 0 13 16 9 13 13 9 2 3 3 16 9 2 7 0 16 9 2
16 3 7 3 13 9 13 1 15 2 16 9 3 13 15 9 2
28 15 13 1 10 9 9 2 12 3 13 9 0 12 9 2 7 12 13 0 13 2 16 13 13 0 9 13 2
26 1 0 13 16 7 3 9 7 9 13 1 9 1 15 9 9 2 1 9 13 9 2 3 7 9 2
55 16 1 9 2 7 1 9 0 9 2 3 13 13 0 9 1 15 9 13 0 2 7 1 15 9 13 1 9 9 9 2 7 13 13 0 9 2 3 16 1 0 15 9 13 7 9 1 9 2 7 9 9 1 9 2
48 7 1 9 9 13 16 15 15 13 2 15 15 13 3 7 0 2 7 3 1 15 3 9 13 9 2 0 15 13 1 15 7 15 9 2 3 13 16 1 0 3 13 9 15 0 3 13 2
18 7 9 1 15 9 13 2 13 15 1 9 1 15 13 1 0 15 2
21 7 3 13 16 2 16 13 15 9 2 3 3 1 15 9 13 9 13 7 13 2
17 7 9 0 9 13 3 13 2 16 9 13 2 1 9 1 8 2
12 3 9 3 13 9 0 2 15 13 1 13 2
27 1 0 13 16 9 0 15 13 9 0 2 15 9 13 13 9 2 16 9 13 1 9 16 9 1 9 2
8 7 1 15 9 13 3 9 2
57 9 7 0 15 3 13 10 9 2 7 13 1 15 16 9 1 9 2 13 13 9 9 2 7 0 15 15 13 9 2 3 3 9 13 1 9 2 9 0 15 13 9 2 3 13 15 9 2 13 9 2 15 13 9 9 2 2
7 7 15 9 0 13 9 2
23 13 13 3 15 15 9 13 2 13 1 9 13 16 9 15 2 16 9 13 15 9 13 2
24 13 7 2 1 15 16 9 9 13 1 9 2 16 10 13 1 9 2 1 15 9 15 13 2
29 7 3 13 16 1 9 0 9 3 9 13 9 9 2 16 9 9 1 0 15 13 16 13 9 9 15 7 15 2
30 3 7 9 1 9 13 13 13 1 9 2 3 16 9 9 13 15 9 1 15 13 2 7 16 15 9 13 9 15 2
38 0 7 9 13 9 1 15 9 0 9 1 9 2 1 9 7 9 9 9 3 0 13 1 9 2 7 13 3 12 2 3 15 9 2 1 15 9 2
43 9 3 0 9 2 3 9 2 13 9 0 9 2 16 13 9 9 2 7 3 1 15 9 13 13 15 16 1 9 2 7 1 9 10 9 0 13 2 3 3 9 13 2
44 9 7 9 1 9 2 15 13 3 1 9 2 3 3 1 0 9 2 0 13 1 9 9 15 13 1 9 2 7 9 9 15 13 1 9 1 9 1 9 7 1 9 0 2
25 3 15 13 13 9 0 2 3 13 9 0 13 1 9 0 2 16 0 13 15 1 9 9 13 2
23 16 3 9 0 13 1 9 3 0 16 9 2 13 16 9 0 13 9 3 0 16 9 2
32 7 16 9 0 13 1 12 9 0 0 2 15 9 9 13 1 0 9 0 2 13 16 9 0 13 12 9 0 1 13 0 2
14 7 1 9 1 9 13 16 9 0 13 9 3 0 2
17 7 3 13 16 15 9 13 0 2 3 1 0 15 13 15 15 2
42 7 3 15 13 9 13 9 1 3 9 2 16 9 15 13 9 9 1 15 9 2 16 3 9 13 9 0 9 1 9 2 3 9 9 13 13 9 0 9 1 9 2
41 15 7 13 2 1 15 16 9 13 9 9 2 16 15 9 13 15 13 2 7 16 13 1 15 0 2 3 3 0 9 13 16 13 1 15 0 2 16 13 0 2
18 3 3 7 16 15 1 9 0 15 13 16 9 0 0 2 13 15 2
18 9 7 2 1 13 0 2 13 15 9 0 2 7 1 15 0 9 2
15 3 13 16 1 10 9 2 15 13 10 9 2 15 13 2
28 3 15 9 13 9 13 1 9 0 2 3 7 9 15 15 13 1 9 15 9 2 7 13 3 9 0 3 2
20 16 3 7 9 9 1 9 13 9 0 2 1 0 7 13 13 9 0 3 2
42 0 13 7 16 1 9 13 1 9 3 0 15 15 1 9 0 13 2 7 3 15 15 13 9 9 2 13 3 9 15 9 9 2 7 3 1 9 7 3 1 9 2
32 7 1 15 3 9 1 9 13 9 10 2 7 3 1 9 7 3 1 9 2 16 1 15 13 16 1 9 15 1 9 13 2
31 7 15 9 9 9 9 2 15 13 15 13 9 1 0 9 2 13 9 9 3 0 3 1 9 2 7 3 3 1 9 2
28 1 0 13 16 9 13 0 1 9 0 2 15 3 13 9 9 7 3 1 9 0 2 7 3 1 9 9 2
29 16 0 9 0 13 1 16 9 13 9 9 15 13 1 0 9 2 1 9 13 2 3 15 13 9 0 7 0 2
16 7 9 0 1 10 9 13 1 10 9 2 15 13 15 9 2
19 9 7 9 13 7 9 15 1 15 13 2 7 9 15 13 1 9 15 2
44 3 13 1 9 0 2 16 9 15 13 1 9 9 2 3 13 1 15 13 9 2 7 1 9 2 15 13 9 16 15 13 2 7 1 9 2 15 13 9 1 9 16 13 2
27 1 0 3 13 16 9 0 1 9 0 13 1 9 10 2 7 1 0 13 1 15 13 2 16 13 4 2
26 7 15 3 13 1 15 15 9 13 2 3 9 0 9 13 16 13 15 10 9 2 15 13 9 15 2
37 3 2 9 13 2 1 12 8 2 16 16 15 9 13 9 1 9 2 3 1 15 13 9 7 12 2 7 3 13 9 15 13 15 9 7 12 2
11 7 9 13 9 0 2 16 1 13 4 2
19 3 2 10 15 13 1 15 9 2 1 15 16 13 2 13 9 1 15 2
21 11 13 15 13 1 9 12 15 12 13 9 15 9 0 15 15 9 9 15 9 13
8 15 15 9 9 9 1 15 13
11 9 1 9 11 9 1 9 11 7 11 13
42 0 15 0 13 9 3 16 1 9 7 9 9 3 13 3 7 1 15 9 3 13 7 15 15 1 13 9 13 13 0 7 13 9 15 1 11 13 15 1 3 9 13
29 15 1 9 9 3 0 9 9 13 16 3 0 9 1 9 13 16 7 15 9 15 13 7 15 1 15 9 9 13
8 1 9 3 0 13 7 0 11
23 15 11 11 11 11 9 9 9 13 9 9 13 7 9 13 16 1 9 15 1 15 9 13
10 0 13 16 9 15 13 0 11 9 13
9 15 1 9 9 13 0 0 9 13
25 1 9 3 9 7 1 9 9 7 9 0 15 9 13 13 15 1 9 12 9 12 1 9 12 13
38 0 9 13 7 9 11 13 13 15 15 1 13 13 13 9 7 9 3 0 9 13 9 3 0 13 16 1 9 9 9 13 1 0 9 9 7 9 13
9 1 0 9 13 9 15 3 13 13
6 1 0 9 9 9 13
6 1 0 9 13 11 13
6 15 15 9 1 9 13
29 3 7 11 9 9 11 15 0 9 9 1 9 13 7 3 9 0 13 16 0 13 13 15 7 9 15 1 9 13
10 15 15 9 15 7 9 0 9 13 13
25 0 9 13 1 15 9 7 9 13 13 7 9 13 1 12 0 7 0 9 0 11 15 13 13 13
7 0 9 13 9 1 9 13
8 9 15 11 1 9 9 13 13
7 13 9 13 13 16 9 13
28 9 13 9 9 11 1 9 15 15 9 3 9 12 12 3 13 7 15 9 9 7 15 15 0 9 13 3 13
21 16 9 1 0 9 13 9 9 15 13 13 9 7 9 1 9 9 13 11 13 13
12 3 7 13 9 3 9 13 16 15 15 9 13
23 3 3 15 1 0 9 0 13 13 13 9 15 15 9 3 12 9 3 12 0 0 9 13
20 9 15 1 15 15 1 13 13 13 16 9 9 9 13 0 1 15 9 13 13
9 12 9 0 9 15 15 9 13 13
40 13 9 7 9 7 9 0 16 0 13 9 9 15 9 7 13 3 1 15 13 9 7 15 1 11 13 7 1 9 0 13 11 7 13 13 1 15 9 15 13
9 13 3 9 12 15 9 9 13 13
9 9 3 0 13 16 3 0 13 13
28 0 1 9 15 3 0 7 0 3 16 1 9 9 7 9 15 3 13 13 11 13 15 7 3 15 9 9 13
9 0 9 9 13 0 7 9 9 11
23 9 15 7 13 16 3 0 9 1 9 0 13 13 7 9 13 16 1 15 9 15 13 13
14 15 9 1 9 13 9 13 15 9 1 9 11 15 13
13 0 9 13 1 9 12 9 0 11 11 11 11 9
29 11 16 15 13 13 15 1 9 15 9 13 13 13 1 9 13 7 3 0 13 9 1 11 0 13 7 1 11 13
49 3 1 15 9 9 0 13 13 9 1 15 13 0 9 15 9 11 7 11 0 9 13 15 13 15 13 1 9 1 15 9 9 1 9 13 3 16 15 9 13 15 13 16 15 9 15 15 13 13
21 11 16 9 13 11 11 9 13 9 7 15 1 9 13 7 1 9 13 13 3 13
17 3 7 9 0 9 13 9 1 9 9 13 13 1 9 7 9 13
17 3 16 9 13 13 16 9 15 13 13 9 13 9 15 1 13 13
41 3 0 9 15 15 1 13 9 7 15 1 9 13 1 9 11 15 1 9 11 13 1 9 11 15 9 9 1 9 13 12 9 12 9 1 9 9 12 9 7 13
5 0 9 13 9 13
11 9 13 16 3 16 15 0 13 13 13 13
38 9 0 9 13 9 13 9 7 0 13 15 9 11 3 0 9 9 13 3 3 3 3 3 16 13 13 13 9 9 7 9 9 7 9 13 0 9 13
13 13 12 1 9 9 15 9 0 1 9 13 3 13
18 0 16 15 9 13 3 13 9 1 11 9 13 16 15 9 1 9 13
37 11 9 7 9 1 9 0 13 7 9 13 9 16 1 0 9 11 9 1 9 13 7 9 9 13 0 9 13 7 3 0 9 15 9 13 13 13
33 3 9 13 7 1 9 13 16 1 9 15 9 13 13 9 7 16 1 15 13 13 9 16 9 9 13 9 16 1 9 7 9 13
22 15 16 13 13 0 1 9 9 13 16 9 0 9 0 9 9 0 3 7 0 0 13
11 1 0 9 0 9 15 13 11 11 9 13
13 3 9 7 9 7 9 9 0 13 9 9 13 13
20 0 0 9 13 1 11 15 13 9 0 9 0 1 9 9 0 9 9 0 13
4 3 1 9 9
6 1 9 1 11 9 13
7 15 13 1 9 1 11 0
19 9 3 1 9 7 9 9 15 9 13 7 1 9 9 13 15 7 9 13
25 3 15 15 9 1 9 0 13 13 16 3 1 9 9 15 9 13 9 1 9 13 9 13 3 13
23 3 9 15 1 11 9 9 7 13 9 15 1 11 13 7 13 15 1 9 9 15 13 0
17 15 9 13 11 3 13 15 13 16 15 9 9 13 1 9 9 13
24 9 13 11 15 1 9 9 7 9 1 11 13 0 9 3 16 9 1 15 9 13 13 3 13
7 15 9 9 7 9 13 13
40 3 1 9 11 0 13 13 12 3 9 9 9 0 9 13 0 3 9 1 9 11 0 13 1 0 9 1 9 12 1 9 13 1 0 9 13 15 3 9 13
9 15 13 7 0 13 0 9 15 13
9 0 15 9 13 7 1 0 9 13
19 0 9 12 16 9 13 9 15 9 11 11 9 13 7 15 9 1 9 13
20 3 7 9 7 9 9 0 15 9 9 11 0 9 9 0 13 15 0 9 13
28 15 1 9 11 3 3 0 7 3 0 9 13 13 16 15 9 11 11 9 11 11 9 11 0 9 15 11 13
18 0 9 13 0 9 9 16 13 13 9 1 11 13 13 7 3 9 13
25 9 0 15 9 13 16 15 15 15 9 12 3 13 16 9 13 0 12 9 13 13 9 1 15 13
11 15 9 11 9 13 15 9 0 9 9 13
5 15 3 1 11 13
22 16 9 9 0 1 9 13 1 0 9 13 7 3 13 9 3 15 11 13 7 13 13
28 16 0 12 9 13 13 16 15 15 9 13 15 9 13 3 13 16 1 0 9 7 15 3 9 13 7 15 13
17 15 3 1 9 0 7 15 13 16 3 9 13 3 9 7 9 13
20 3 3 13 16 0 9 3 13 1 9 9 0 7 9 9 9 13 7 9 13
4 0 11 3 13
24 3 15 3 9 13 16 0 9 15 9 0 13 9 13 7 3 3 13 3 3 9 9 0 13
11 15 16 15 9 15 0 13 3 13 3 13
18 7 3 13 16 3 7 13 1 15 13 3 13 3 7 1 9 13 13
29 3 16 0 9 13 13 3 3 0 9 16 15 0 9 1 9 1 9 13 16 9 16 9 16 9 13 9 13 13
39 16 15 3 13 3 16 9 1 15 15 13 16 15 15 13 13 13 7 16 9 1 9 15 15 9 7 15 13 3 16 9 3 13 15 1 15 9 13 13
15 11 13 3 9 1 0 15 13 13 16 9 13 3 13 13
6 15 9 9 0 13 9
4 0 9 13 13
7 0 9 9 1 0 9 13
30 0 13 11 9 7 15 1 9 12 12 15 1 15 9 7 9 7 15 9 13 13 13 15 13 15 1 9 9 9 13
17 15 3 0 9 13 0 9 1 9 9 9 13 7 0 1 15 13
16 11 15 1 9 13 7 3 13 1 9 9 9 9 9 7 13
10 3 3 11 9 9 15 13 3 13 13
19 3 1 9 3 3 9 1 9 0 3 13 7 3 9 3 3 0 9 13
22 0 3 9 15 9 11 9 13 3 13 3 13 16 9 1 11 9 13 1 15 13 13
5 9 1 9 13 9
4 13 13 13 13
81 3 15 3 13 13 7 9 13 15 9 9 9 13 13 13 15 9 15 0 9 1 9 13 1 0 11 7 11 15 0 9 13 15 9 13 9 15 13 0 7 9 9 7 1 15 13 9 3 15 13 16 16 3 7 13 3 7 1 9 13 13 3 0 9 3 0 9 1 15 3 13 3 16 0 1 9 15 9 13 9 13
15 13 0 15 9 1 9 3 13 15 3 0 13 3 0 9
12 0 0 7 0 9 9 13 16 9 13 15 13
11 1 0 15 9 15 7 1 9 13 9 13
6 0 1 15 13 3 13
23 3 3 16 0 9 13 11 13 13 15 15 15 1 9 13 7 1 0 9 3 3 13 13
22 11 0 9 11 11 11 9 13 13 7 16 0 0 0 9 13 13 3 9 13 11 13
8 13 1 0 15 15 1 9 13
5 0 3 1 15 13
3 13 13 0
14 15 13 11 9 9 0 1 9 1 9 9 0 9 0
13 0 9 7 15 9 0 13 7 9 1 13 0 13
35 0 9 9 15 9 3 13 7 1 15 13 3 7 3 3 7 3 1 0 9 3 13 7 0 9 9 9 1 9 9 3 0 7 0 13
16 15 1 9 9 13 9 1 9 7 0 15 13 1 15 9 13
31 13 7 13 9 1 0 9 13 3 15 9 11 7 9 16 15 9 9 15 13 7 11 9 1 0 9 9 7 9 13 13
15 9 9 9 3 3 1 9 7 3 1 0 15 13 9 13
38 13 3 1 13 11 16 9 0 0 0 3 9 13 13 9 15 9 13 1 11 7 15 9 3 9 15 9 11 9 13 11 13 15 9 0 13 9 13
55 15 9 13 16 1 0 9 0 9 13 16 1 9 9 9 13 16 9 1 15 13 13 16 15 15 3 3 9 15 7 9 7 3 0 15 13 16 1 9 9 13 3 13 9 13 3 1 15 7 0 13 7 9 13 13
22 0 15 9 12 13 16 11 9 0 1 9 0 9 0 1 15 9 0 9 9 9 13
31 3 16 15 13 11 1 15 13 13 7 0 9 13 1 11 11 11 9 11 9 0 15 15 0 15 9 9 13 1 15 13
21 3 13 15 15 0 1 9 1 11 13 13 7 13 15 3 15 1 15 1 15 13
19 13 7 13 16 1 15 9 9 7 0 1 15 9 13 13 7 9 13 13
34 13 15 0 13 0 3 7 15 1 15 0 3 15 9 13 3 16 16 15 9 0 3 7 1 0 11 0 0 1 9 13 1 15 13
15 15 9 7 9 3 3 1 13 9 7 3 1 9 15 13
9 15 3 7 9 0 7 9 9 13
22 3 16 15 15 1 11 0 13 16 15 0 9 9 1 0 13 15 13 3 15 9 13
11 15 1 9 13 16 0 11 9 1 15 13
5 13 13 9 13 13
20 0 15 1 15 9 13 13 16 7 9 0 9 7 15 9 15 9 7 9 13
2 9 13
5 15 1 15 13 13
7 15 0 13 15 9 13 13
8 13 16 1 0 9 15 9 13
6 0 15 11 9 13 13
11 11 9 13 16 15 13 15 1 13 13 13
4 13 13 0 13
5 15 15 9 13 13
18 0 1 0 9 0 9 15 9 13 1 15 13 9 7 15 1 15 13
21 11 11 15 9 0 0 13 7 1 9 11 11 7 3 1 11 11 13 1 9 13
39 0 9 16 0 9 1 11 13 0 1 9 9 3 3 12 7 12 9 13 3 7 3 3 1 9 13 7 15 9 7 11 13 13 11 9 13 1 15 13
18 13 9 15 1 11 13 13 1 9 13 15 15 1 0 9 7 9 13
7 11 15 9 1 0 9 13
2 9 13
16 0 9 15 13 9 9 13 7 12 9 12 1 15 9 9 13
32 3 0 9 16 3 9 13 3 9 9 13 13 7 16 1 11 9 9 3 0 7 0 3 3 12 9 12 13 9 0 13 13
9 3 9 1 9 13 7 11 13 13
11 0 9 1 9 11 11 9 9 9 9 13
41 9 7 16 9 13 9 13 1 15 13 3 3 16 3 0 9 13 9 3 13 7 3 16 9 0 13 13 13 13 9 7 9 13 15 1 0 9 13 7 13 13
18 16 15 9 13 9 15 11 1 9 9 13 9 7 15 13 9 9 13
11 0 3 1 9 0 0 9 13 9 12 0
23 1 0 9 12 9 15 1 11 0 3 13 7 15 9 13 3 16 1 15 0 9 9 13
11 9 1 15 15 9 13 9 1 12 9 13
13 15 0 9 13 15 9 9 13 1 0 15 9 13
20 11 3 15 3 15 1 9 13 9 16 13 15 9 9 9 13 13 15 9 13
9 9 9 0 9 13 3 9 9 13
8 15 13 9 13 1 15 9 13
44 9 0 1 9 13 9 16 0 15 9 12 9 9 13 7 13 16 9 15 13 3 7 13 3 7 9 13 3 3 13 13 0 16 3 13 9 13 9 9 13 7 0 9 13
18 3 9 13 7 9 13 7 16 9 13 3 12 9 9 3 15 13 13
43 13 9 7 13 15 9 7 9 15 9 12 3 12 9 9 13 7 0 9 13 1 9 15 1 9 13 13 13 7 15 13 9 15 1 9 15 13 3 13 7 9 13 13
14 3 16 13 15 9 3 13 0 15 3 13 1 9 13
8 0 1 9 7 9 15 15 13
17 3 0 0 9 16 1 9 0 1 9 13 13 13 9 13 15 13
36 1 0 9 3 1 9 13 13 3 16 1 9 9 13 7 1 9 0 1 15 13 9 13 7 0 1 9 9 7 9 7 9 13 15 7 13
10 3 16 13 13 9 9 7 15 13 13
9 3 11 9 7 12 1 9 13 13
14 1 0 9 3 9 12 12 13 15 7 0 9 3 13
15 11 1 9 9 9 7 13 16 15 9 16 7 15 9 13
9 15 9 13 1 15 9 15 13 13
11 9 15 9 9 13 9 1 9 1 15 13
30 15 16 15 1 9 13 15 7 1 9 13 3 7 13 13 9 13 7 15 1 0 9 15 3 13 15 9 13 13 13
12 3 16 11 13 9 9 9 15 1 15 13 13
54 16 0 13 7 13 9 13 3 9 12 12 0 9 15 9 13 7 9 13 16 9 13 9 13 7 9 9 13 16 1 0 9 9 15 9 7 13 7 3 13 13 13 0 9 1 9 9 13 1 11 9 7 9 13
19 15 3 11 13 15 1 9 13 0 16 13 7 13 16 15 13 13 13 13
9 0 15 9 9 9 13 1 9 13
29 9 9 9 1 9 15 3 13 13 13 13 7 16 15 9 13 3 15 13 15 9 13 9 13 16 0 9 9 13
36 15 0 3 9 13 16 13 0 9 3 9 13 13 16 1 9 9 9 15 1 11 13 1 15 9 1 9 9 13 7 0 11 9 9 7 13
14 9 13 9 16 0 9 13 13 16 1 9 15 13 13
17 15 0 9 13 15 7 3 1 0 9 9 7 9 3 15 13 13
37 1 9 9 9 13 13 9 0 13 7 1 11 13 15 1 9 3 9 13 13 15 9 9 13 15 15 9 13 13 7 3 3 3 9 9 9 7
15 9 13 9 9 12 12 9 12 12 9 12 9 12 9 12
6 9 15 13 3 12 12
16 15 15 9 13 9 13 3 11 13 13 13 9 12 12 7 12
13 9 9 13 0 3 11 9 9 9 1 11 13 13
16 13 16 15 9 0 11 1 9 0 13 15 7 11 13 9 13
12 15 13 15 9 15 1 0 9 1 15 13 13
21 0 9 13 9 9 13 7 9 13 16 15 13 3 15 0 9 13 13 1 15 13
28 0 9 13 0 9 9 15 1 13 1 11 13 13 7 16 15 3 1 0 1 15 15 7 9 1 15 13 13
29 3 3 15 0 13 7 13 16 15 15 13 13 3 16 15 15 13 13 3 16 16 13 13 0 1 9 15 13 13
6 13 13 1 0 11 9
5 11 0 9 13 12
7 0 0 9 13 9 0 9
7 0 3 3 12 12 11 13
14 16 9 7 9 7 9 9 9 0 7 0 13 13 0
10 3 13 1 11 1 12 7 12 12 9
11 0 9 13 13 15 9 15 9 15 9 13
55 15 9 9 7 13 15 7 15 9 7 9 0 9 7 9 0 3 1 11 13 13 13 9 9 13 0 9 7 9 13 9 13 15 3 7 9 13 3 7 9 1 9 0 13 3 7 13 16 0 1 0 9 7 9 13
18 12 15 13 1 15 9 9 15 13 3 13 16 13 7 9 15 9 13
24 1 15 9 15 1 9 13 7 11 1 9 13 9 13 16 0 3 7 9 13 3 7 9 13
54 7 3 0 9 3 9 13 13 3 16 11 9 9 1 0 9 13 0 7 9 9 0 15 13 0 0 11 13 7 3 1 0 9 0 9 13 13 3 16 0 9 3 9 12 9 12 1 15 13 15 9 7 9 13
17 3 7 3 13 13 0 1 9 9 3 7 0 9 9 1 0 13
43 11 3 16 3 9 9 9 13 15 9 13 13 1 11 3 7 3 13 9 0 15 9 13 7 1 15 15 9 9 7 13 16 15 9 3 1 9 7 1 9 15 13 13
6 3 13 15 9 3 13
33 16 15 1 11 9 7 0 13 9 15 9 0 13 13 15 9 13 16 9 13 15 9 15 9 13 1 9 13 9 7 15 13 13
18 0 16 13 11 13 3 13 16 1 15 9 15 1 15 13 0 9 13
29 11 7 9 15 7 9 7 0 9 7 9 9 0 13 13 16 0 9 9 11 13 11 7 15 1 11 9 13 13
15 0 9 1 11 13 15 15 13 0 9 9 1 11 13 13
19 13 11 0 1 15 9 15 0 9 13 15 0 13 7 0 9 13 9 13
9 15 9 13 7 1 0 9 0 13
16 0 9 13 11 9 9 9 13 13 7 13 15 0 9 9 13
14 0 15 13 9 7 9 15 7 9 13 11 9 9 13
5 0 9 13 9 13
56 7 1 15 0 9 15 13 3 15 0 9 13 7 13 13 1 0 16 9 9 9 7 3 9 1 9 13 1 9 7 9 13 9 13 0 7 9 13 1 11 7 9 13 15 1 0 9 9 0 0 15 7 9 0 13 13
45 3 3 9 13 11 13 7 1 11 0 0 9 13 9 0 0 13 3 7 15 9 0 7 0 13 13 16 1 15 11 13 3 3 9 9 7 13 1 9 13 7 3 1 11 13
6 15 9 3 3 13 13
13 0 3 11 0 15 9 0 9 13 16 13 3 13
16 0 9 11 13 16 15 0 1 11 9 13 15 1 15 13 13
10 16 15 0 15 13 0 1 15 13 13
28 3 15 3 7 1 9 1 0 9 11 13 13 15 11 13 3 7 9 1 0 9 7 9 1 12 9 13 13
19 15 3 0 13 15 1 15 11 15 9 13 7 11 7 3 9 0 9 13
14 0 9 1 11 13 3 1 15 11 9 1 0 9 13
48 16 0 15 9 7 0 9 13 16 1 9 15 9 7 9 1 9 13 13 0 15 9 7 0 9 13 16 1 9 13 13 13 3 7 1 0 9 13 15 7 13 13 0 13 15 1 15 13
11 3 16 15 9 9 3 1 11 1 11 13
19 3 9 15 13 1 9 13 9 7 13 16 15 0 13 9 15 13 0 13
14 16 3 13 15 9 7 0 0 9 7 9 1 15 13
35 16 3 13 15 16 11 11 11 11 9 9 13 16 15 11 9 13 15 9 9 0 13 13 9 0 7 9 9 0 13 15 9 9 3 13
16 1 0 11 13 9 13 9 16 15 13 15 15 13 3 13 13
14 3 9 0 13 3 1 0 9 7 1 15 9 13 13
20 16 15 9 0 3 13 3 15 9 13 3 13 15 1 9 0 1 15 9 13
15 9 15 16 9 9 13 7 9 13 7 13 13 0 13 13
11 0 11 9 13 15 15 9 9 15 0 13
26 9 15 9 13 3 13 3 7 0 3 7 15 9 9 9 13 16 1 15 13 15 13 9 7 3 13
3 16 13 13
16 13 15 0 9 0 1 9 15 1 9 12 9 3 13 9 13
14 0 0 9 11 9 13 7 9 1 9 7 1 9 13
13 9 13 16 9 15 3 1 11 13 13 9 15 13
9 15 3 9 3 13 9 11 13 13
13 9 3 9 12 9 1 9 11 13 15 11 13 13
6 0 13 11 7 11 9
12 3 9 0 3 3 13 13 0 9 1 11 13
8 15 16 13 3 15 13 11 13
38 3 15 9 15 1 9 9 13 0 13 1 0 9 9 15 7 9 9 3 13 16 0 1 13 9 13 9 3 16 9 11 3 9 13 3 0 9 13
26 0 9 15 13 3 3 9 12 3 9 13 9 13 0 9 3 16 9 0 9 1 15 9 9 9 13
9 0 9 13 9 13 7 1 9 13
14 3 11 0 0 0 7 9 13 13 7 9 3 9 13
61 16 0 9 1 11 9 0 9 7 9 13 1 9 15 9 7 9 7 9 15 0 9 9 9 0 9 7 9 1 9 13 13 3 9 15 1 0 13 3 9 3 7 9 9 13 13 13 0 3 9 15 9 13 16 3 3 15 9 9 7 13
18 15 15 15 9 13 15 15 1 13 0 13 13 13 16 15 9 13 13
8 0 9 13 16 9 9 13 13
14 13 1 9 7 15 9 13 7 1 9 15 0 9 13
5 3 0 9 9 13
21 0 9 7 9 3 3 15 15 0 1 9 9 13 9 9 7 15 7 9 13 13
34 15 15 1 0 3 0 13 13 3 15 9 13 7 9 9 7 9 9 15 13 1 15 7 11 7 9 0 16 3 3 13 13 13 13
22 0 3 11 13 16 9 13 7 9 13 13 3 13 9 13 9 3 7 1 9 9 13
8 11 15 9 3 9 0 9 13
9 3 0 3 3 15 1 9 13 13
20 15 3 13 13 15 9 7 9 9 13 15 3 7 15 3 7 9 0 9 13
10 7 3 1 15 9 7 1 0 9 13
14 13 0 9 9 9 15 9 9 7 9 1 11 11 13
18 13 3 3 1 11 0 9 15 3 15 9 7 9 15 1 15 13 13
24 1 15 13 13 3 13 1 15 0 9 3 16 15 3 0 1 9 13 0 3 0 7 9 13
46 16 15 0 9 7 9 9 13 0 16 13 13 13 9 9 13 9 11 16 0 9 9 15 7 9 13 3 7 15 9 13 13 3 1 9 7 13 3 13 3 9 7 9 3 9 13
18 15 9 1 9 0 7 0 9 13 0 3 15 3 13 15 9 13 13
22 15 15 9 1 9 0 9 9 7 9 13 13 3 16 7 1 9 9 13 7 13 13
4 0 15 13 9
6 1 9 15 0 9 13
15 16 3 13 9 13 3 7 9 13 13 15 15 0 9 13
21 13 3 15 9 9 13 3 13 7 3 9 13 9 13 7 15 9 13 9 13 13
32 3 15 15 1 0 9 13 13 13 7 0 9 1 0 9 9 13 16 3 3 13 13 3 1 15 9 7 9 7 9 0 13
22 3 16 3 15 13 3 15 1 0 0 9 13 1 15 3 13 15 7 15 0 9 13
11 0 9 11 7 13 3 7 1 9 13 3
43 0 9 13 0 1 9 13 13 15 9 0 7 9 7 9 9 13 13 13 0 7 0 11 1 9 9 15 9 13 16 1 15 0 9 13 15 7 13 1 9 13 0 13
14 3 0 9 1 9 9 7 0 9 9 13 16 11 13
31 15 9 13 7 9 13 1 11 16 1 9 15 0 9 13 16 12 3 12 9 9 0 9 13 1 0 9 3 13 13 13
21 0 9 16 9 3 13 1 9 0 13 13 11 9 1 15 12 9 12 7 12 13
21 15 3 1 9 13 15 1 15 13 13 16 3 13 15 7 0 1 9 13 13 13
40 3 13 9 11 3 7 15 1 9 13 13 16 15 15 3 13 13 3 13 0 7 1 9 13 1 15 0 9 7 0 1 15 9 13 15 9 13 16 9 13
8 9 9 13 13 1 0 9 0
19 3 3 16 9 3 3 7 1 15 13 11 13 16 15 9 1 9 11 13
8 13 15 16 1 9 1 15 13
4 15 1 9 13
45 11 16 3 7 9 13 9 13 13 3 7 9 15 9 9 13 13 0 13 13 15 9 0 9 13 3 0 9 9 0 15 3 3 13 13 16 9 3 0 16 15 9 13 13 13
12 13 15 1 9 0 9 0 9 13 1 9 13
10 9 13 0 7 1 15 9 0 3 0
11 0 9 0 3 9 1 9 11 7 11 13
7 3 3 13 13 1 9 13
11 9 11 15 9 13 9 12 1 0 9 13
6 3 9 11 0 9 13
13 11 1 9 16 13 7 1 15 0 1 9 13 13
20 0 16 3 7 9 3 7 9 13 0 13 9 7 9 15 7 9 0 9 13
38 13 3 3 0 3 7 0 9 9 15 1 9 13 15 9 9 3 3 7 0 1 15 13 13 3 15 9 0 11 9 9 13 3 3 16 15 9 13
21 9 0 0 13 9 16 9 7 9 3 3 15 15 13 7 9 9 9 0 13 13
13 15 3 1 9 9 0 13 15 15 13 15 13 13
32 13 3 0 15 9 1 9 13 3 7 9 7 15 9 9 13 9 13 16 15 9 9 9 13 13 3 3 15 3 11 13 13
6 11 1 9 11 0 13
5 1 15 9 0 13
12 13 11 15 3 15 9 7 13 7 13 1 9
11 9 13 1 11 1 15 13 9 15 9 13
9 9 13 9 9 15 9 13 13 13
8 3 15 9 7 9 15 9 13
12 15 11 9 1 15 13 13 7 1 15 9 13
11 0 15 9 1 15 12 9 13 7 13 13
9 16 3 13 13 15 3 0 13 13
16 16 9 13 13 0 13 1 9 13 15 15 9 1 0 9 13
16 9 9 0 15 9 7 9 3 9 13 13 7 15 0 9 13
16 0 9 9 13 16 3 13 3 13 7 16 9 3 13 7 13
8 15 3 1 11 13 3 9 0
11 3 1 0 9 9 9 0 11 9 9 13
3 15 15 13
5 3 1 15 9 13
8 9 15 0 13 11 3 0 15
22 3 0 13 3 13 16 1 15 9 9 13 3 3 15 13 0 16 1 15 9 15 13
15 13 15 13 13 11 9 16 9 1 11 13 15 13 9 13
32 3 16 15 13 0 15 9 9 7 9 0 0 13 13 15 15 1 15 1 15 9 13 13 15 15 9 7 9 15 9 13 13
26 3 16 13 7 0 9 11 15 13 0 15 0 9 13 7 15 9 13 13 1 15 15 9 7 9 13
13 0 1 11 1 0 9 13 13 3 9 13 3 13
25 3 7 15 3 7 9 0 9 13 16 3 13 9 13 3 7 15 13 11 3 13 11 3 9 0
23 9 13 13 9 7 9 1 11 11 11 15 9 0 13 3 7 1 9 13 3 7 9 13
14 3 16 0 15 9 13 13 9 0 0 13 1 11 9
23 16 0 1 9 13 11 13 13 9 11 3 9 13 7 1 15 13 9 9 7 1 15 13
19 11 13 9 13 15 7 1 15 13 15 7 13 16 15 3 9 1 9 13
39 16 1 9 9 13 13 15 9 1 9 11 13 15 11 9 13 9 7 1 15 15 9 13 0 7 9 9 3 13 0 0 9 9 7 13 0 9 13 13
7 9 3 11 1 11 9 13
17 13 15 1 0 9 15 1 15 13 13 3 7 13 13 13 1 15
18 16 7 3 9 9 13 7 16 15 3 13 1 15 9 15 1 15 13
22 13 11 9 13 3 13 3 3 3 16 3 0 9 9 13 3 13 16 9 1 15 13
59 0 13 13 11 11 11 11 11 11 9 0 9 7 9 9 15 9 1 11 11 9 9 13 13 7 1 9 7 1 9 0 9 15 0 3 11 0 9 13 7 16 1 15 13 9 9 3 13 1 15 13 7 3 11 11 15 9 11 13
10 0 13 15 13 11 13 7 1 15 13
16 15 16 1 15 1 9 11 13 9 15 0 13 15 1 15 13
7 13 13 13 7 1 9 13
14 0 9 9 13 7 12 9 12 1 11 9 1 9 13
31 3 0 9 1 9 11 15 9 13 7 12 9 12 1 15 9 13 0 9 16 9 9 7 15 1 9 7 9 13 11 13
26 1 0 9 9 0 12 11 1 9 15 9 13 7 9 13 13 16 16 13 11 9 13 15 9 3 13
4 0 9 3 13
8 9 0 13 9 15 15 9 13
4 9 12 13 12
16 3 9 9 0 7 0 15 1 15 9 0 0 15 9 9 13
5 1 15 15 9 13
6 0 16 15 13 0 13
8 16 15 0 9 13 9 13 13
36 3 15 9 15 13 11 13 16 3 9 13 1 0 9 15 1 9 9 13 3 9 12 1 0 9 0 9 13 9 7 0 13 1 15 9 13
11 0 7 0 9 1 9 13 0 9 13 13
18 3 3 9 12 12 0 1 15 9 11 13 15 9 15 13 7 9 13
14 9 3 11 3 3 13 12 9 9 13 0 9 13 13
9 13 9 12 3 9 13 7 9 9
24 0 9 9 15 11 1 9 15 9 15 13 3 7 1 0 9 13 9 13 9 7 13 9 13
13 3 3 3 3 15 13 13 3 9 9 1 9 13
7 3 3 3 1 9 13 13
14 9 9 15 9 11 0 7 13 7 13 9 1 9 13
36 16 1 9 13 11 3 11 9 3 13 0 13 9 16 1 9 0 9 13 16 9 9 15 9 7 9 13 3 9 13 1 9 13 3 7 3
14 15 3 13 3 13 9 9 13 16 1 0 9 9 13
13 3 0 9 11 9 15 9 15 3 13 13 13 13
23 9 15 1 9 9 1 9 0 13 16 3 9 9 0 1 9 9 13 16 1 9 9 13
34 3 3 3 9 15 9 9 13 3 7 13 0 9 9 9 9 9 9 9 9 15 7 9 15 9 7 9 13 16 15 9 1 9 13
15 11 0 9 0 9 7 9 13 16 15 9 15 15 9 13
14 15 1 0 9 16 0 9 3 0 9 13 13 9 13
24 3 15 3 1 9 9 13 9 13 3 7 9 3 3 7 13 16 9 9 1 9 13 3 13
6 13 9 3 9 13 13
11 3 9 3 1 9 15 9 13 9 9 13
15 13 13 0 15 15 1 0 13 7 9 9 13 7 3 13
21 16 9 9 1 0 9 13 7 1 9 13 13 1 0 9 3 9 15 15 9 13
13 3 0 7 9 13 13 13 7 9 13 15 9 13
12 1 0 13 11 15 9 13 1 9 13 15 13
6 0 15 13 9 15 13
24 12 13 11 9 12 0 9 15 9 15 1 13 0 0 9 11 9 15 1 11 13 1 9 13
5 15 1 0 9 13
8 12 9 0 0 13 0 13 13
19 11 11 11 16 1 9 1 9 0 9 13 13 1 0 11 9 9 13 13
39 15 3 9 11 3 0 3 0 9 9 13 16 9 0 9 11 15 0 7 9 13 1 9 9 15 13 13 3 7 15 9 1 0 9 7 9 15 9 13
5 9 9 15 13 0
9 3 11 11 13 7 1 15 13 13
14 0 9 1 11 13 9 15 1 9 11 13 9 13 13
14 15 3 15 0 11 13 13 13 13 0 1 15 9 13
19 11 12 9 12 0 9 13 3 3 3 9 9 13 1 9 1 9 9 13
3 9 11 13
9 15 1 0 11 1 9 13 13 13
38 16 13 11 1 0 11 3 16 3 13 0 1 15 9 13 9 7 3 11 0 13 15 9 15 0 13 11 9 13 1 9 0 13 9 7 1 15 13
35 3 16 1 0 9 13 3 15 3 9 3 1 11 13 13 3 9 0 9 13 7 13 1 11 3 13 3 15 9 7 9 9 0 9 13
19 1 0 3 16 1 11 1 0 7 15 15 1 13 9 9 13 3 9 13
9 15 3 3 0 9 9 15 13 13
25 0 9 9 7 13 11 12 9 1 0 11 0 13 7 13 9 1 0 11 15 13 11 11 9 13
10 15 16 3 9 9 13 13 1 9 13
24 13 9 9 0 7 9 15 0 9 13 16 15 15 1 15 13 13 15 7 1 0 9 0 13
11 15 3 15 13 9 13 9 1 12 9 13
13 9 0 13 9 13 9 7 3 12 1 9 9 13
51 0 15 9 1 9 13 9 7 15 1 11 13 15 1 0 13 0 7 13 15 15 9 16 3 9 3 9 9 7 15 15 0 9 7 0 9 13 12 9 12 7 9 1 15 13 13 13 16 1 15 13
18 16 1 15 13 15 9 15 7 1 9 13 7 15 1 9 13 3 13
40 0 9 13 13 1 9 11 7 3 13 1 9 9 3 13 9 7 15 0 9 13 13 0 7 13 15 9 15 9 15 11 13 9 9 7 1 15 9 13 13
18 15 1 9 13 16 0 9 9 0 15 9 0 7 9 1 9 0 13
28 1 9 15 15 15 13 13 9 13 3 16 9 9 7 13 15 15 9 1 0 9 9 1 0 9 13 13 13
12 0 1 15 9 7 9 7 9 7 9 9 13
4 9 15 13 0
6 9 0 0 7 9 13
16 3 13 9 11 1 0 1 9 9 7 9 0 9 15 9 13
8 9 13 9 12 13 12 0 12
11 3 9 15 3 0 1 15 13 3 7 13
22 12 12 9 9 12 12 9 12 12 9 12 12 9 12 12 9 7 9 3 9 12 12
13 9 9 9 9 15 12 9 9 13 13 3 12 12
9 15 15 1 0 3 1 9 13 13
24 15 11 9 3 13 13 3 9 0 0 7 9 13 9 9 13 16 1 0 9 12 9 13 13
16 15 13 13 16 15 9 9 1 9 9 13 7 15 9 13 13
41 16 15 9 9 1 12 9 13 1 15 13 13 3 7 3 3 13 1 0 15 13 9 7 1 9 13 9 11 15 13 1 0 9 9 9 13 13 7 3 9 13
33 15 9 7 9 12 9 9 9 13 7 1 15 15 13 0 1 9 13 7 9 1 9 0 7 9 16 1 9 1 15 13 13 13
5 1 0 9 9 13
16 3 9 13 7 1 0 9 9 11 11 11 9 1 12 9 13
11 1 0 9 9 9 9 11 13 12 9 12
8 15 1 9 0 9 9 13 13
5 3 0 9 13 13
7 9 0 3 9 9 13 0
4 15 3 3 13
14 3 16 0 9 9 7 9 13 1 9 13 9 13 15
31 16 9 13 9 13 11 9 0 9 7 9 1 15 15 3 9 13 12 1 15 15 9 1 9 1 11 13 9 1 15 13
23 3 1 0 9 11 0 9 13 15 9 1 11 13 9 7 9 9 7 9 0 9 9 13
19 15 9 7 9 1 9 9 9 13 13 7 9 0 1 9 9 13 9 13
31 3 3 1 9 13 9 7 9 13 15 9 9 7 3 13 13 13 1 9 11 15 9 13 7 1 12 9 3 12 9 13
13 15 9 3 9 7 9 13 3 12 9 12 9 13
14 11 3 7 1 9 9 7 1 0 9 9 9 13 13
90 3 15 3 13 0 13 9 1 9 1 9 13 9 0 7 0 3 0 9 3 9 13 13 3 1 9 13 3 1 1 9 13 3 9 9 13 13 13 7 1 15 9 9 9 13 7 1 9 3 13 3 1 9 13 1 15 9 0 9 0 9 13 3 9 12 7 1 0 9 9 13 3 7 9 13 16 16 9 13 9 16 3 9 13 1 9 13 15 13 13
26 0 13 12 9 15 3 13 1 9 13 16 16 15 9 13 9 13 13 0 12 9 1 9 1 9 13
9 9 13 3 0 1 15 7 9 9
6 0 16 15 13 9 13
15 15 3 16 1 0 9 13 13 16 13 13 0 1 9 13
7 3 9 0 1 12 9 13
14 3 15 13 9 13 0 9 9 15 11 15 1 9 13
16 9 3 1 0 9 1 9 11 13 15 13 1 15 9 13 13
20 11 0 13 1 11 15 9 7 0 9 9 9 9 7 9 13 7 1 15 13
10 9 13 15 1 9 13 0 15 9 13
17 1 15 9 0 0 13 13 9 9 13 0 7 15 13 9 13 13
39 9 3 7 1 13 9 7 1 9 13 9 15 13 13 3 7 15 1 9 0 13 13 9 13 7 15 9 0 13 13 9 13 13 0 13 9 15 15 13
28 7 15 1 9 3 9 9 13 1 15 13 3 13 16 3 1 15 3 1 9 9 13 7 0 9 9 0 13
19 1 0 9 1 0 9 0 3 9 15 13 16 11 7 9 9 9 13 13
12 0 13 16 3 13 3 7 15 9 13 3 13
35 0 9 13 0 9 0 1 9 7 9 9 13 15 0 9 3 7 9 16 15 15 0 9 9 13 7 9 13 13 13 16 0 9 9 13
9 0 11 11 7 11 11 11 9 13
8 11 11 9 1 9 12 13 13
28 15 0 13 7 0 12 9 13 0 9 15 13 13 16 1 0 9 1 15 13 13 13 3 7 9 15 9 13
24 0 16 13 1 9 13 3 7 15 9 3 7 9 13 13 9 13 9 15 1 9 15 9 13
13 3 1 15 9 0 15 9 15 13 15 13 9 9
13 1 9 9 13 13 15 7 1 9 3 13 13 13
28 3 0 9 11 16 15 9 1 9 7 9 13 1 9 9 15 0 9 13 9 13 7 0 9 1 9 11 13
22 15 1 9 13 13 16 0 1 9 13 13 1 9 9 9 7 9 0 13 13 3 13
11 3 15 1 9 9 9 1 9 0 9 13
37 3 9 1 9 13 9 13 9 7 13 9 9 15 3 7 13 3 9 3 7 13 7 9 9 13 9 1 11 1 9 13 7 13 9 16 13 13
26 11 9 13 0 9 7 15 11 9 12 9 9 7 15 1 9 13 1 9 9 13 9 7 1 9 13
50 15 16 15 15 7 15 1 9 11 13 7 1 0 9 11 1 9 3 12 9 12 13 15 0 3 1 9 13 9 1 11 13 7 9 13 13 15 1 15 9 7 9 13 3 7 1 9 0 9 13
22 3 16 1 9 13 9 7 3 13 9 9 7 1 9 13 9 15 9 9 1 9 13
15 1 0 11 3 1 9 9 13 9 9 1 15 13 13 9
10 9 15 9 1 9 7 9 9 0 13
26 13 1 15 9 15 13 9 1 11 1 9 13 15 9 9 7 13 7 1 9 13 7 9 0 9 13
19 15 16 13 9 9 1 15 9 13 15 9 7 9 16 3 9 13 13 13
29 11 9 11 7 9 9 15 15 1 9 13 7 13 13 7 16 13 9 0 1 9 9 7 9 9 13 12 9 13
15 0 13 15 7 9 1 9 13 1 0 9 1 9 9 13
8 15 15 15 7 15 1 9 13
4 15 9 9 13
10 15 1 9 9 7 11 16 13 3 13
6 15 13 9 1 15 9
6 13 9 0 0 7 9
12 13 15 3 7 9 13 3 7 15 9 9 13
21 16 1 15 9 9 9 13 13 1 9 11 9 1 9 15 3 3 12 9 12 13
18 1 0 9 15 9 13 9 7 3 9 13 3 1 9 7 9 0 15
9 3 0 15 13 16 0 9 9 13
10 13 3 1 15 9 9 7 13 1 9
20 9 15 7 1 9 1 9 0 13 1 0 9 13 15 1 9 9 9 3 13
64 16 1 0 9 0 7 9 0 11 13 3 9 13 15 1 0 3 3 1 9 13 13 0 9 9 9 15 9 13 9 1 9 13 7 0 13 1 0 9 9 0 9 13 3 7 13 15 9 16 0 9 1 9 13 0 7 9 0 9 13 0 1 9 13
12 15 13 9 7 13 13 16 0 3 13 3 13
13 0 9 16 9 9 15 13 3 13 15 9 9 13
9 9 9 13 0 15 9 15 9 13
12 9 1 0 3 0 1 9 11 15 3 13 13
26 1 0 9 0 9 9 13 0 0 7 0 9 3 12 0 0 1 0 9 0 16 3 3 3 13 13
8 1 0 9 9 1 0 15 13
6 9 13 9 9 3 12
6 11 9 13 13 15 9
13 7 9 9 7 9 3 15 13 3 9 1 9 13
6 1 15 0 9 9 13
14 3 12 9 15 3 13 13 0 9 13 9 7 9 13
13 9 15 1 9 9 7 9 13 1 9 9 9 13
43 16 15 0 3 1 9 1 15 13 7 3 1 9 1 15 9 13 3 7 15 3 3 15 1 9 0 9 0 13 13 13 13 3 9 12 15 0 13 9 13 9 13 13
22 0 3 13 7 13 0 9 1 9 13 16 3 12 9 7 1 9 7 1 9 9 13
16 0 3 9 0 9 1 15 9 7 15 15 1 9 13 13 13
6 11 15 12 9 13 13
10 9 13 15 13 9 16 1 9 13 13
4 1 9 13 9
8 15 0 3 9 13 9 13 13
2 9 13
2 9 13
10 15 9 0 9 9 9 7 9 9 13
43 0 9 12 9 13 9 9 7 9 9 16 0 9 13 15 13 13 3 3 3 0 15 13 3 1 15 13 13 7 16 1 9 0 7 9 0 9 11 13 3 13 9 13
17 15 1 9 7 9 9 15 3 11 9 13 7 1 15 15 13 13
17 11 0 9 13 1 13 9 15 9 9 13 13 7 1 9 0 13
9 7 1 0 3 13 9 13 13 13
28 9 0 13 0 9 7 3 0 1 13 9 16 3 3 1 9 13 7 3 1 9 13 9 7 9 13 9 13
57 13 9 3 3 9 9 7 9 9 3 3 9 0 9 7 9 13 16 0 9 15 15 1 9 9 13 9 7 0 3 3 13 13 9 13 3 7 0 9 13 3 7 15 1 15 9 9 13 13 3 7 1 12 15 9 13 13
10 3 1 0 9 9 9 3 9 0 13
43 9 0 7 0 9 3 1 0 9 9 13 9 13 9 7 9 13 9 7 13 9 3 0 0 9 13 3 1 9 0 1 9 13 7 13 13 13 9 0 9 15 13 13
18 15 13 9 3 13 7 1 9 0 13 3 13 9 13 9 1 9 13
24 3 15 1 9 0 12 9 0 7 0 13 9 15 1 13 13 1 9 0 1 0 9 9 13
39 3 0 3 9 1 9 7 1 0 9 13 16 1 0 9 11 0 7 3 0 1 15 9 0 13 15 9 0 9 9 11 15 9 9 13 1 0 9 13
34 0 9 9 15 0 7 9 9 15 1 15 3 13 15 0 9 9 13 13 16 15 1 9 13 13 9 13 7 3 15 1 9 9 13
17 3 15 15 1 9 13 9 9 7 13 15 7 15 1 9 13 13
50 15 15 9 13 9 9 15 1 9 9 9 13 0 15 9 9 1 9 13 1 11 13 16 9 9 9 13 9 13 7 3 13 13 9 9 9 9 13 13 7 1 15 9 13 13 13 15 9 9 13
12 9 13 13 7 9 9 7 15 9 13 9 13
144 11 1 0 9 9 1 0 9 13 3 15 13 9 7 1 12 9 13 0 9 13 9 15 0 1 9 13 9 13 0 9 15 9 13 9 7 13 9 13 0 9 15 3 9 7 13 7 13 1 0 9 11 11 11 0 9 0 0 7 9 13 16 3 15 13 3 13 0 13 0 7 3 15 1 0 13 9 9 13 7 9 13 9 3 7 1 9 1 0 9 13 13 7 1 15 9 13 7 9 13 1 0 13 3 7 15 13 9 15 13 13 9 1 0 9 13 16 15 3 1 9 13 1 0 9 13 9 7 3 13 0 13 9 9 13 7 9 13 13 16 3 9 13 13
28 15 9 9 13 9 7 13 9 16 1 15 15 1 9 9 3 1 0 15 9 9 13 13 3 9 9 13 13
26 11 16 0 9 15 3 13 3 13 1 9 13 9 9 13 16 3 15 9 13 7 13 9 1 9 13
21 15 13 16 15 15 9 13 3 7 13 16 13 1 9 13 3 13 7 3 13 13
41 0 9 0 9 9 13 13 16 15 3 15 9 13 13 9 13 9 13 9 13 9 13 3 0 0 13 9 3 16 9 9 9 13 15 1 9 9 15 0 9 13
60 3 9 3 1 0 9 9 0 9 13 16 16 0 15 13 0 13 13 7 1 15 9 13 0 13 7 13 9 15 13 3 1 9 9 1 15 13 7 9 13 13 16 3 3 0 9 9 13 13 13 13 13 0 9 13 0 9 13 0 9
7 15 0 1 0 9 9 13
49 0 9 13 7 3 1 9 9 7 9 9 13 0 9 15 3 1 9 9 7 1 9 7 9 13 13 0 9 13 16 9 15 13 13 15 0 13 15 15 13 9 9 1 11 13 15 7 15 13
25 7 1 13 9 9 1 12 1 12 9 1 9 12 12 3 1 12 15 9 13 13 15 13 13 13
31 15 11 16 1 0 7 0 13 9 13 3 13 15 7 9 7 9 13 13 7 0 13 16 1 9 7 9 15 15 7 13
18 9 1 15 3 13 16 15 9 9 9 13 0 9 13 1 9 9 13
14 0 9 9 7 13 15 15 1 12 9 3 9 13 13
6 15 9 0 0 9 13
10 3 0 9 9 7 0 9 1 9 13
40 15 13 1 9 9 7 13 15 16 9 1 9 15 7 11 13 0 9 15 15 1 13 7 13 3 13 1 9 11 13 9 1 15 7 9 12 12 9 3 13
26 0 1 15 9 0 9 1 0 13 16 3 9 13 3 13 13 9 15 15 9 13 0 15 9 9 13
16 7 0 9 9 15 0 1 9 9 13 0 7 9 1 15 13
15 3 9 9 12 1 9 12 12 0 7 9 13 9 15 13
23 3 9 13 9 13 9 3 13 13 3 13 1 9 7 13 9 16 0 9 1 0 9 13
31 15 3 9 7 15 9 3 9 0 9 3 3 15 9 1 9 9 15 9 15 9 13 0 9 9 1 9 15 13 13 13
18 15 15 3 0 13 0 7 15 9 13 1 15 15 13 13 9 3 13
23 15 13 16 1 0 9 13 15 9 1 9 0 13 3 1 0 1 9 13 1 15 13 13
20 1 0 11 13 15 3 9 15 3 3 15 9 13 16 16 9 9 13 15 13
8 7 9 15 13 9 3 9 13
17 15 15 15 1 9 13 13 0 7 13 16 15 9 9 0 9 13
10 9 13 1 15 0 15 15 13 13 13
44 9 0 9 1 9 1 9 15 13 1 9 13 3 16 3 9 9 9 7 9 9 9 13 7 3 3 9 0 3 3 13 13 13 7 1 9 13 9 13 0 9 9 13 13
59 0 3 13 3 13 13 9 16 9 13 15 9 13 7 3 3 13 13 3 1 0 15 13 7 13 9 3 9 1 9 13 7 9 13 15 3 3 9 9 13 9 13 0 9 3 3 0 1 15 9 9 13 15 9 3 1 9 9 13
10 13 3 9 12 12 0 1 9 13 13
19 3 0 9 13 9 16 3 13 15 7 13 9 15 9 0 9 0 11 13
12 1 15 15 13 9 9 1 15 13 13 12 12
39 0 9 1 11 11 15 1 9 12 13 1 9 9 9 9 9 9 9 15 13 0 9 11 7 13 0 13 13 15 0 9 1 9 9 7 9 0 13 13
33 0 9 13 15 11 13 0 0 9 1 0 9 13 13 16 1 0 9 15 1 11 13 9 1 11 13 15 15 9 13 13 13 13
16 15 9 11 16 1 11 11 7 13 13 0 9 1 15 13 13
18 1 0 7 9 1 9 11 9 12 9 13 13 15 1 0 9 13 15
33 16 1 11 13 11 11 11 1 9 0 7 9 9 1 9 9 9 7 13 15 1 9 9 7 9 11 7 9 11 1 0 11 13
14 0 13 16 9 13 13 16 1 0 9 9 13 9 13
41 11 0 15 9 13 9 7 0 15 13 13 1 15 3 9 9 7 13 7 9 13 13 9 12 1 9 13 7 0 1 0 0 9 9 1 9 9 15 13 11 13
13 15 9 13 1 9 3 0 13 9 0 9 3 13
20 16 0 1 12 9 9 13 0 9 0 13 9 13 0 0 1 0 13 9 13
6 0 9 9 9 7 13
61 15 15 1 9 13 16 3 9 9 13 9 7 13 9 13 3 16 9 3 0 0 13 9 12 7 0 3 15 9 13 9 13 13 13 1 9 13 3 3 16 1 9 9 16 15 1 9 1 9 13 7 9 13 3 0 3 9 15 13 13 13
33 13 16 15 1 15 9 13 9 9 13 7 9 3 3 9 9 7 3 0 9 9 11 13 13 7 0 9 0 9 13 15 13 13
41 0 9 13 11 16 3 7 9 9 9 7 3 13 13 3 7 1 9 0 7 9 3 13 13 16 9 13 9 7 13 15 1 9 13 13 9 3 13 9 13 13
17 0 3 9 13 0 13 1 0 9 9 3 9 9 13 7 9 13
21 0 9 13 3 16 0 9 15 13 13 7 13 9 13 9 1 15 9 9 13 13
6 9 9 7 1 9 13
42 15 3 0 9 3 13 3 7 15 3 9 1 9 0 13 7 15 9 9 13 9 13 13 3 13 7 9 13 7 0 13 16 9 9 9 13 9 13 15 0 9 13
77 16 3 3 9 12 3 13 7 3 3 9 7 3 9 15 13 7 9 3 13 0 7 15 9 13 7 9 13 13 9 7 13 3 1 0 13 9 11 11 11 0 9 9 15 0 9 0 13 9 13 7 3 11 11 9 9 9 7 9 0 7 9 1 11 13 7 12 13 9 9 13 16 9 13 0 9 13
34 3 13 9 3 9 0 13 3 13 9 7 3 3 9 13 13 15 7 1 9 13 3 13 9 1 9 13 7 15 9 9 1 9 13
22 15 13 13 13 7 3 15 9 9 13 3 7 13 15 13 3 7 15 13 9 9 13
43 3 13 9 15 15 1 9 13 9 13 3 13 13 7 1 9 12 3 12 15 9 9 1 9 13 13 3 0 9 13 0 13 1 9 13 7 3 1 9 3 0 13 13
54 15 9 13 16 3 9 13 11 13 7 15 15 1 9 9 13 13 15 13 9 13 3 9 9 13 0 9 15 0 9 9 13 1 9 13 13 7 15 9 13 7 9 13 0 9 1 9 3 1 9 13 3 7 13
34 0 9 13 16 15 1 9 11 13 11 13 7 3 13 9 1 11 13 13 16 15 3 9 13 7 9 13 13 0 9 1 11 13 13
5 15 9 0 13 9
19 15 16 1 0 9 9 9 13 9 9 7 9 0 1 0 9 9 9 13
21 15 1 9 13 11 11 13 1 9 11 11 9 1 11 11 11 1 11 11 1 9
52 0 13 9 3 0 9 15 9 0 9 0 16 7 9 13 9 0 15 1 11 13 13 7 9 7 9 9 0 0 13 7 1 0 9 9 7 9 0 9 13 15 13 15 15 3 15 0 9 13 13 13 0
19 1 0 13 9 13 11 7 11 16 1 15 15 15 9 15 11 13 13 13
58 0 9 0 13 3 13 9 0 7 0 9 0 1 9 11 11 7 13 7 3 13 9 1 15 9 1 15 13 15 3 0 9 13 0 7 15 9 9 13 13 0 7 9 13 16 1 0 9 15 1 0 13 13 3 9 9 13 13
32 15 1 9 11 1 11 0 13 16 0 13 3 9 3 0 13 1 9 11 15 13 1 11 9 1 9 13 9 9 7 13 13
14 0 9 3 13 0 16 3 1 9 9 13 1 9 13
27 0 13 9 13 9 9 13 1 9 9 9 7 9 13 3 7 15 9 1 9 9 3 1 15 13 13 13
46 7 3 16 15 1 9 13 3 15 0 9 13 9 3 7 15 9 13 9 3 7 0 9 3 9 13 13 9 9 9 13 7 3 0 13 9 1 13 9 3 1 0 7 0 11 13
24 0 13 9 9 13 9 1 9 1 9 13 9 1 11 3 11 3 9 13 13 3 0 13 13
13 9 15 1 0 9 9 9 9 9 9 9 9 13
10 9 1 11 15 1 0 9 13 13 13
42 13 0 9 9 13 15 3 13 7 3 0 11 1 0 9 13 9 13 9 9 9 13 1 9 9 13 9 3 9 9 1 0 16 0 9 13 0 9 15 0 13 13
14 3 11 11 9 1 9 15 0 9 11 13 1 9 13
26 11 11 1 9 0 12 7 0 9 9 1 11 13 13 16 1 0 9 9 1 11 13 7 0 9 13
18 11 11 11 9 1 9 12 1 9 9 9 7 13 15 0 9 13 13
27 11 11 9 9 0 7 9 15 1 9 7 9 0 7 13 9 13 13 13 7 16 3 13 1 9 13 13
5 15 3 0 9 13
41 13 0 9 3 9 9 16 13 1 0 9 9 7 3 7 9 9 13 16 1 9 15 9 13 15 13 3 9 12 9 3 7 9 16 3 13 9 9 1 9 13
6 3 15 9 9 9 13
39 7 16 3 9 9 3 13 13 9 9 7 9 7 0 9 9 13 15 9 13 13 0 9 9 13 15 9 0 9 13 15 15 13 15 7 1 0 9 13
10 3 15 9 1 0 9 13 13 7 13
14 9 3 0 3 15 9 16 3 9 7 9 9 13 13
12 9 3 13 7 3 9 1 9 9 9 7 13
11 9 0 13 1 9 1 15 9 7 9 13
12 9 1 0 1 9 9 13 9 0 9 9 9
6 9 1 9 0 9 13
42 9 1 9 9 7 3 13 7 1 9 9 7 0 9 9 7 3 15 13 3 0 0 16 0 9 11 0 7 9 9 13 7 0 9 9 13 9 3 3 3 13 13
28 1 0 9 15 9 0 9 9 13 16 12 9 7 9 9 13 0 1 9 9 1 9 9 0 13 0 7 0
24 13 16 16 15 9 13 7 9 13 3 7 1 9 13 3 7 1 9 13 15 9 7 9 13
8 15 9 15 15 9 9 13 13
25 0 13 9 11 3 13 3 0 9 13 3 7 9 9 13 9 13 3 7 15 13 13 13 13 9
25 15 3 13 7 3 1 9 13 13 3 12 9 15 0 7 15 9 9 0 13 1 9 15 0 13
25 3 7 3 11 15 9 13 7 9 9 9 7 15 0 9 13 13 13 15 13 7 15 9 9 13
6 9 3 13 3 13 13
28 9 3 13 3 0 9 9 1 0 9 13 16 3 7 1 0 9 3 3 9 13 13 7 13 1 9 3 13
19 12 13 0 9 9 13 1 15 9 0 13 13 7 9 3 0 9 0 9
30 0 13 9 13 1 9 15 15 9 3 13 7 3 3 16 1 9 11 7 15 9 9 13 16 15 3 3 9 13 13
15 15 3 9 7 9 0 3 13 0 9 1 9 1 9 13
19 13 3 13 9 16 0 0 7 0 9 13 9 0 9 13 1 9 9 13
18 15 16 9 13 13 13 0 9 16 0 9 15 13 9 9 9 13 13
23 7 3 13 1 0 9 9 3 9 13 0 3 9 7 9 13 16 15 1 9 13 3 13
9 15 3 9 1 9 13 0 13 9
25 3 0 15 13 13 16 0 1 15 9 9 9 1 9 13 16 1 9 3 12 3 1 9 9 13
26 3 16 15 9 15 3 0 9 1 15 15 9 7 9 13 3 13 3 9 15 3 13 1 12 9 13
7 3 15 15 7 15 11 13
17 1 15 3 3 11 13 13 16 3 1 0 9 1 9 9 9 13
8 3 15 9 13 0 1 9 13
19 16 0 1 9 13 11 11 11 1 0 9 15 1 11 13 1 9 9 13
16 0 13 11 7 9 9 13 0 15 9 15 13 1 15 9 13
23 7 0 0 9 9 9 9 7 9 15 13 16 9 9 13 13 9 13 15 7 1 11 13
40 11 0 15 9 9 9 15 13 16 11 1 15 12 12 9 13 3 7 13 9 13 9 13 16 3 3 3 9 1 9 11 13 7 3 15 9 9 3 15 13
13 0 7 9 9 13 16 3 1 9 9 9 13 13
19 0 13 9 9 0 15 9 7 0 13 9 1 0 15 9 9 15 1 13
15 0 0 9 9 7 13 16 1 9 13 7 15 13 13 13
10 15 3 1 9 1 15 13 9 9 13
28 15 9 0 11 1 9 13 13 3 7 3 13 16 0 9 11 3 1 9 9 13 7 1 11 9 13 9 13
17 15 3 13 13 13 15 9 9 3 13 13 3 13 1 9 13 13
24 0 9 13 3 3 11 0 7 9 1 9 13 16 1 15 13 13 9 16 13 7 1 9 13
18 15 9 13 0 3 13 9 9 9 7 13 15 9 9 13 1 9 13
12 9 13 9 13 7 3 1 0 0 3 9 12
6 11 15 13 13 9 13
13 13 9 1 15 15 13 9 3 12 9 9 13 13
25 13 13 9 9 9 9 7 9 9 9 7 0 9 9 16 3 12 3 15 9 13 7 3 9 13
11 15 13 0 9 9 15 13 0 9 15 13
23 3 12 9 7 1 0 9 11 7 1 11 9 11 13 0 13 9 7 15 15 3 11 13
22 3 3 1 9 13 9 0 7 0 13 9 3 0 7 3 13 1 9 13 9 15 13
52 0 3 9 11 11 16 1 11 13 15 3 3 13 13 0 9 11 13 16 13 1 0 9 15 9 13 3 0 3 9 11 11 11 9 9 13 13 13 7 3 11 11 9 9 13 13 3 0 15 9 13 13
33 3 9 0 13 9 9 7 13 0 3 9 0 11 7 11 7 11 15 13 9 11 9 0 1 0 9 3 13 1 9 9 9 13
17 3 9 15 13 7 13 15 3 0 9 15 1 9 1 9 13 13
6 0 15 13 13 9 13
33 13 13 3 7 3 16 9 0 9 0 1 15 9 0 11 9 13 13 15 3 15 1 9 7 1 0 9 9 9 13 13 13 13
11 15 0 9 13 11 1 9 9 9 13 13
7 15 3 13 9 9 7 13
47 0 3 9 13 3 9 1 9 9 7 13 15 9 13 3 0 9 3 16 0 9 1 15 9 9 7 13 3 9 15 15 0 9 13 13 13 9 1 11 13 15 7 1 9 16 13 13
7 15 9 13 9 13 13 13
24 7 1 0 9 15 15 13 9 15 1 9 9 11 15 9 9 13 1 12 0 15 0 9 13
17 3 7 3 9 9 13 13 15 15 15 13 15 15 9 13 9 13
34 1 0 11 9 13 13 9 1 0 9 9 13 16 1 9 9 13 3 7 3 13 13 13 1 9 3 16 0 9 9 13 1 11 13
32 3 3 9 13 16 9 7 9 9 7 9 13 0 9 15 3 13 13 13 13 9 3 3 13 13 9 1 15 13 9 13 13
12 13 3 1 0 9 9 15 13 0 11 0 11
5 3 9 9 7 13
12 15 9 0 1 9 7 0 9 9 9 13 13
19 9 3 15 13 15 3 1 11 11 15 9 13 0 7 9 9 0 13 13
12 0 9 9 0 9 13 9 13 9 15 13 13
14 0 9 1 9 13 3 15 0 13 13 0 9 9 13
47 0 16 1 9 7 0 9 9 9 7 15 15 3 13 13 3 0 13 13 13 9 9 13 1 9 9 13 7 16 1 9 9 0 0 15 13 13 13 1 9 7 1 9 0 9 13 13
11 0 9 13 1 9 13 9 9 15 9 13
37 0 9 13 11 16 15 9 7 9 9 9 15 9 0 1 13 13 7 15 9 13 13 3 3 13 16 1 9 13 13 15 15 13 1 9 9 13
74 3 16 15 9 13 15 0 9 13 9 9 9 7 13 9 7 15 1 9 3 3 11 13 9 9 7 13 7 1 9 9 13 9 7 9 13 13 16 3 1 9 3 7 3 3 13 9 7 1 9 0 13 3 3 13 9 13 9 9 11 13 3 0 13 9 1 0 9 9 13 0 7 9 13
15 11 9 9 13 16 0 9 9 7 15 13 15 13 13 13
58 0 3 13 13 13 0 9 15 9 9 13 0 1 9 13 7 0 9 13 16 1 9 9 13 13 15 9 9 7 1 9 13 3 1 0 15 13 9 13 7 0 13 3 1 9 9 13 16 3 1 0 13 7 15 9 13 13 13
20 3 3 9 1 0 9 13 15 13 9 15 3 1 9 9 13 13 3 13 13
13 0 13 9 0 9 11 15 11 13 9 7 3 13
15 15 1 9 13 9 9 9 9 9 9 9 9 9 9 9
12 0 0 9 9 9 13 16 9 13 0 13 13
41 0 3 9 11 16 3 13 3 9 13 3 16 15 11 13 9 9 7 13 15 1 9 13 3 7 1 15 3 9 1 9 13 13 0 9 3 13 13 3 9 13
10 15 3 0 9 3 0 9 9 13 13
24 3 16 13 0 9 15 9 13 13 13 7 13 0 7 9 7 9 13 3 15 15 7 15 13
32 1 15 9 9 16 11 13 9 7 13 13 3 7 9 3 13 13 13 1 9 15 3 1 15 9 9 13 7 1 15 9 13
20 15 3 9 13 15 7 1 9 13 7 0 13 3 0 9 13 0 1 15 13
39 0 9 0 9 0 9 13 16 3 9 7 0 9 1 15 13 15 0 9 13 0 9 13 9 13 16 9 3 13 7 9 9 3 1 9 9 13 3 13
27 3 13 15 15 9 9 9 7 13 11 9 13 7 1 9 9 7 0 3 9 15 3 9 13 1 9 13
31 0 15 13 13 9 15 13 9 11 11 11 11 9 9 9 7 3 9 0 9 9 9 11 13 3 3 1 9 3 11 13
15 9 13 13 16 1 9 0 9 13 9 13 7 9 9 13
9 9 9 13 3 0 7 0 9 15
16 0 12 9 13 13 1 15 3 0 12 9 13 9 1 9 13
8 0 15 3 13 15 7 0 13
8 0 3 3 9 3 1 9 13
20 7 0 7 0 9 1 15 15 13 3 7 3 9 13 12 1 9 13 9 13
16 3 7 3 9 7 0 9 9 7 9 13 3 7 13 1 9
33 15 9 7 9 9 7 0 9 7 9 9 16 1 9 15 9 7 9 13 15 3 1 9 13 7 9 13 7 0 9 9 9 13
27 7 1 0 15 9 13 16 9 0 3 9 1 9 13 15 15 1 9 0 13 9 9 0 7 13 1 9
20 9 13 9 3 3 16 15 9 13 15 13 13 3 16 15 9 1 15 13 13
33 3 3 9 15 3 9 13 15 7 0 13 9 9 13 3 13 7 15 13 1 15 13 0 7 0 0 0 9 0 16 13 9 13
23 0 9 3 1 9 13 7 9 13 9 7 0 13 9 13 1 15 15 3 16 9 13 13
10 3 1 15 9 0 9 3 0 13 13
23 3 0 13 13 9 3 3 1 15 9 13 9 0 9 13 0 9 9 15 9 13 3 13
13 3 12 1 9 1 9 3 12 9 12 9 13 13
15 1 0 9 13 9 15 13 9 0 7 0 3 13 9 9
27 15 3 16 13 0 9 13 0 0 3 16 11 13 3 7 1 15 9 13 7 0 1 9 0 13 9 13
26 0 16 9 0 3 9 13 1 9 9 7 9 9 13 3 13 3 0 15 13 7 3 0 0 7 13
10 1 0 9 13 9 7 9 15 3 13
18 1 9 3 9 13 7 0 9 11 9 13 1 11 13 15 9 9 13
10 0 1 15 9 9 9 9 9 7 13
62 0 15 13 16 3 7 9 13 1 9 9 3 7 3 13 1 9 9 13 13 15 1 15 9 9 7 13 7 9 9 13 3 13 7 15 0 9 12 9 9 13 0 0 7 9 13 15 1 9 9 1 9 0 13 1 9 1 11 1 15 9 13
31 0 13 9 7 15 13 3 16 0 9 9 15 1 11 13 0 13 9 13 7 15 15 9 13 0 9 9 15 15 9 13
25 0 1 9 11 0 13 7 9 9 13 16 13 1 9 13 0 7 0 3 9 13 15 0 13 13
41 13 3 0 0 9 16 7 9 3 0 13 13 7 15 15 15 1 15 9 13 7 13 13 7 9 1 9 9 13 15 7 1 9 13 15 7 3 9 13 13 13
29 0 9 7 9 13 1 0 3 9 9 13 15 15 1 9 13 3 13 16 0 9 13 7 0 1 9 15 13 13
25 3 16 13 0 15 13 13 13 13 13 13 9 1 3 15 9 1 9 13 7 15 16 1 11 13
7 15 15 13 1 15 13 0
18 15 9 13 9 3 3 13 7 1 9 9 7 9 15 13 9 9 13
18 9 0 13 9 7 13 9 1 0 9 13 13 15 1 9 13 9 13
15 1 15 16 0 9 9 13 9 1 15 13 15 0 13 9
31 9 3 7 0 9 0 9 13 3 7 3 13 16 13 16 9 13 16 9 9 13 1 9 13 15 9 13 13 3 7 13
7 0 3 13 13 0 13 9
11 7 15 9 13 7 13 0 13 15 9 13
12 15 12 9 13 15 3 9 3 0 0 13 13
10 0 3 1 9 13 15 15 3 13 13
7 1 0 11 15 13 13 13
11 15 15 1 15 9 13 13 16 1 11 13
12 3 7 0 13 15 15 9 13 3 13 0 13
15 3 7 15 1 11 13 9 15 13 0 3 9 1 9 13
4 0 15 9 13
16 9 0 15 1 15 13 13 7 9 13 1 9 0 1 11 13
7 3 16 3 15 9 13 13
9 3 0 3 11 1 15 13 13 13
19 13 3 0 9 9 1 15 15 9 1 13 13 7 9 1 9 1 9 13
17 11 16 1 9 3 3 9 12 12 13 3 13 13 1 15 9 13
9 15 1 9 13 3 16 3 13 13
19 15 16 9 7 9 15 9 13 9 13 0 9 15 1 11 13 15 13 13
8 1 0 9 13 15 9 9 13
16 0 15 11 0 0 13 13 16 9 9 13 9 15 15 13 13
13 3 15 3 3 12 9 12 9 9 13 0 9 13
11 3 0 9 3 0 13 16 1 15 9 13
26 3 1 9 15 1 15 9 13 13 15 13 16 9 9 13 7 16 0 13 13 3 15 1 9 3 13
34 3 0 13 9 15 1 9 13 13 7 9 0 7 15 13 0 1 9 13 7 3 13 13 16 3 3 9 13 16 1 9 9 15 13
21 1 0 9 0 11 0 0 9 13 15 9 1 9 15 9 13 9 1 9 15 13
12 0 16 9 13 1 9 9 13 0 1 9 13
8 0 9 13 13 3 13 3 13
23 16 13 0 9 13 13 7 0 9 15 3 9 13 3 13 13 9 15 9 13 7 13 13
27 0 13 9 11 3 7 3 15 9 13 3 7 9 13 13 1 15 15 1 9 7 9 13 9 3 9 13
28 13 3 16 9 9 13 9 7 13 0 12 13 13 7 13 9 9 3 3 1 15 9 12 9 9 13 13 13
8 15 1 9 13 15 9 13 13
16 0 15 9 9 13 9 7 16 0 9 13 13 13 9 13 13
20 9 0 13 7 3 12 12 9 13 3 1 9 9 13 16 15 13 9 13 13
36 15 15 9 3 13 7 9 9 15 7 9 15 3 7 9 13 3 7 9 13 9 13 13 9 3 1 9 13 7 9 13 7 9 9 13 13
16 15 9 16 9 7 9 13 9 15 0 9 9 13 1 9 13
17 15 9 15 3 9 13 13 3 15 13 7 1 9 9 7 9 13
18 3 0 9 9 9 7 3 1 15 15 9 13 11 7 13 3 13 13
6 1 15 13 11 9 13
46 9 1 9 9 13 16 15 13 13 9 13 9 7 0 13 15 1 9 13 7 16 1 9 11 7 11 13 0 9 13 0 9 13 0 15 1 9 13 7 3 9 9 9 9 13 13
9 11 15 15 1 9 13 13 9 13
15 0 9 9 7 9 13 15 9 13 13 15 1 15 13 13
4 0 11 9 13
12 0 9 13 0 1 9 11 13 15 11 13 13
32 15 0 13 0 16 16 13 9 3 3 13 16 1 11 13 15 3 9 15 13 13 16 13 7 13 7 13 9 0 9 11 13
37 13 3 16 0 9 9 9 7 9 15 3 13 13 13 7 9 11 13 3 7 9 13 1 9 15 15 1 11 1 9 9 13 15 7 1 0 13
23 1 15 16 11 9 13 15 13 15 15 15 11 7 9 13 15 13 13 9 0 9 11 13
20 16 15 0 9 1 11 13 3 9 13 3 15 15 13 9 7 9 1 11 13
10 0 15 1 9 9 7 0 9 3 13
28 0 13 9 7 9 0 9 11 13 7 0 0 9 13 3 1 0 9 9 16 9 7 9 9 0 0 13 13
7 9 0 9 1 13 9 13
9 11 0 1 9 15 13 11 13 13
19 7 9 13 3 7 3 0 13 13 3 7 15 3 7 9 0 9 13 13
23 3 16 0 9 13 9 13 1 9 9 9 7 9 3 0 15 13 7 3 3 13 9 13
4 9 9 0 13
46 0 16 9 13 1 9 13 9 7 13 3 9 9 3 1 9 7 3 7 3 16 1 9 9 13 0 3 0 12 1 0 9 13 9 9 0 1 0 9 1 9 7 9 9 13 13
26 15 13 7 1 0 9 13 0 13 9 9 7 0 9 9 16 15 0 9 9 15 13 0 3 13 13
10 0 13 9 13 13 7 9 9 7 13
53 7 9 3 9 7 1 0 9 9 3 13 15 1 9 13 7 1 15 9 13 9 9 13 7 15 3 1 9 0 9 16 16 9 9 16 7 9 13 9 9 13 1 9 13 0 9 0 9 9 13 7 9 13
12 9 12 15 9 13 13 13 15 9 13 9 13
12 11 1 15 9 9 0 9 13 1 9 9 13
8 3 1 0 9 1 15 9 13
36 3 9 1 0 9 15 9 13 13 13 9 13 13 15 15 1 9 7 9 1 15 13 9 15 13 15 7 15 13 15 7 1 9 7 9 13
33 11 0 9 1 15 9 13 15 9 9 7 13 9 7 13 15 1 9 9 13 7 0 9 15 13 16 1 9 13 0 1 15 13
10 0 13 13 9 3 9 0 15 0 13
8 3 9 9 13 7 3 13 13
47 15 3 11 13 15 0 9 13 15 9 9 9 13 13 16 9 9 13 16 9 13 16 9 9 13 9 3 12 1 11 13 3 7 1 9 7 1 9 13 13 15 1 11 13 9 7 13
59 0 9 9 0 11 16 1 0 9 16 15 11 1 9 13 0 13 9 3 1 11 13 13 16 15 3 0 9 9 15 3 13 9 13 7 16 9 9 1 9 13 13 3 0 15 9 13 13 16 3 9 13 9 9 13 9 9 9 13
6 15 15 3 9 13 0
41 3 13 1 15 3 9 3 7 15 13 9 9 3 7 15 7 15 9 13 3 7 15 9 9 13 7 15 9 13 3 7 15 13 1 0 9 9 0 9 13 13
16 1 0 13 3 16 9 13 0 13 13 11 11 1 9 0 13
11 0 13 16 13 15 9 1 15 3 3 13
17 3 9 3 1 0 9 7 15 0 9 1 0 9 13 9 13 13
27 3 9 15 13 7 1 9 13 1 9 1 0 9 9 1 15 9 13 15 13 9 13 7 9 9 0 13
47 15 13 3 13 13 7 16 1 0 9 13 15 9 13 7 1 15 3 11 15 0 9 13 9 3 13 15 7 9 7 9 13 7 15 15 0 13 13 15 7 9 1 0 9 0 13 13
19 0 13 15 13 13 9 13 7 16 9 0 9 13 15 7 3 3 13 13
42 16 1 0 9 11 9 13 9 13 1 0 9 9 1 15 9 13 15 15 1 0 9 9 13 16 9 0 7 15 9 0 9 9 0 13 15 7 0 15 13 13 13
38 0 15 11 3 3 13 13 16 3 7 1 9 9 13 13 3 7 9 13 1 9 9 9 13 3 7 0 0 9 9 11 13 13 0 15 9 9 13
6 15 13 15 1 9 13
25 9 3 12 0 13 13 7 3 3 13 1 12 13 9 13 15 3 9 0 13 9 9 9 7 13
3 0 9 13
26 0 9 11 11 11 7 11 11 11 9 1 9 7 1 0 9 9 1 15 1 15 9 3 13 13 13
14 11 11 11 9 1 0 9 15 3 13 13 9 13 13
27 1 15 16 3 3 13 13 0 9 9 3 0 1 0 9 11 13 7 3 1 15 9 13 9 9 0 13
20 15 9 0 13 9 7 3 9 0 9 13 16 1 9 0 1 9 9 13 13
18 0 1 13 3 0 9 13 16 0 9 3 13 1 9 0 1 9 13
45 3 9 9 7 9 13 7 15 1 11 13 7 15 13 13 13 13 7 3 9 0 9 3 7 3 0 9 13 16 16 0 7 0 9 13 1 9 7 1 9 15 9 1 15 13
29 0 13 7 9 7 9 12 9 13 0 13 9 7 13 9 3 12 9 12 1 0 9 13 0 7 0 9 9 13
64 13 1 0 9 0 9 16 9 1 9 3 1 0 13 3 13 9 3 0 9 13 9 0 7 0 9 9 13 3 7 1 9 13 7 1 9 13 7 1 9 13 13 16 0 7 1 9 7 3 1 9 13 15 9 0 0 9 3 9 13 7 9 13 13
22 15 9 15 13 7 0 3 9 9 0 3 0 9 7 9 15 1 0 13 9 13 13
6 15 9 0 9 15 13
19 3 7 9 9 7 9 9 7 0 9 9 13 9 13 7 3 3 9 13
29 7 15 9 13 3 1 9 9 15 0 9 9 13 13 9 16 0 9 9 3 13 13 13 9 16 13 9 9 13
9 15 3 15 9 0 7 9 9 13
15 0 16 9 0 13 15 1 9 13 7 1 9 9 13 13
13 3 15 13 1 15 16 0 9 13 0 1 9 13
5 13 13 1 15 3
18 9 3 13 15 9 3 1 9 15 0 1 9 13 13 13 9 13 13
3 0 0 13
8 15 1 9 0 1 0 9 13
20 15 16 13 11 9 0 9 3 0 9 9 13 13 7 15 13 13 0 9 13
17 15 16 1 9 13 15 15 13 1 9 9 13 7 15 1 9 13
14 3 7 3 13 13 16 9 9 13 7 9 13 3 13
7 0 12 1 0 9 11 13
15 3 1 0 9 11 11 13 15 3 13 1 11 1 11 13
18 0 0 1 9 13 16 1 15 9 9 11 9 13 13 7 1 9 13
20 3 9 13 13 7 1 13 9 0 9 9 1 9 13 7 1 9 16 13 13
24 11 13 16 16 3 1 9 9 13 9 1 15 13 9 1 9 13 13 15 9 13 9 7 13
5 15 0 9 3 13
10 9 1 0 9 13 0 9 15 13 13
18 3 15 1 9 13 13 9 7 3 13 7 15 9 7 15 11 13 13
28 0 9 9 13 1 9 0 16 13 1 11 13 9 12 1 15 3 13 13 15 9 13 1 0 9 0 9 13
15 15 3 9 13 16 9 13 3 0 9 1 9 13 9 13
21 0 9 13 16 13 9 0 15 9 0 9 0 1 11 13 13 15 7 0 13 0
32 3 12 9 7 0 9 15 11 1 9 13 9 13 7 0 15 1 9 13 13 9 13 3 7 15 15 9 7 13 7 13 13
26 0 9 13 0 16 13 9 9 0 7 9 13 1 13 0 0 0 15 3 13 13 0 9 9 13 13
35 3 7 3 9 13 15 15 13 13 7 15 13 15 1 13 9 13 9 7 16 15 13 13 1 11 13 9 1 0 9 1 9 13 3 13
73 15 9 13 9 11 15 1 9 1 11 13 1 15 13 16 7 9 7 9 7 9 9 13 13 7 9 9 1 9 9 13 15 0 13 3 0 16 1 9 11 9 13 0 13 13 13 9 13 9 9 7 15 13 7 9 1 9 13 16 0 13 7 9 13 15 3 9 13 9 1 11 13 13
15 3 3 9 13 3 1 9 13 7 15 3 1 9 13 13
25 3 11 16 3 15 9 13 3 7 1 9 9 15 7 1 15 16 9 13 13 13 0 15 13 13
17 3 16 0 9 1 9 13 12 9 13 0 16 13 3 3 13 13
57 16 0 13 9 1 9 12 13 13 15 13 12 3 7 15 1 0 9 9 9 13 16 9 9 1 9 13 9 3 1 9 13 15 15 1 9 9 1 9 13 11 13 9 0 16 9 13 1 0 9 13 15 1 9 11 9 13
35 11 0 15 13 13 15 0 1 9 13 9 9 15 1 9 13 15 1 1 0 9 13 1 0 12 1 9 13 0 13 7 3 15 13 13
22 16 3 3 1 9 13 15 1 9 13 7 3 13 7 13 9 1 15 9 9 13 13
22 3 16 15 1 0 9 13 9 9 12 13 0 13 9 3 15 13 13 3 1 9 13
20 3 13 13 9 1 13 13 3 13 0 13 0 0 9 13 7 9 7 9 13
6 9 0 13 1 9 9
22 9 3 3 1 9 13 7 3 9 13 16 16 0 1 9 9 13 0 1 15 9 13
9 15 9 13 15 9 0 11 9 13
5 3 15 9 9 13
5 15 15 1 9 13
24 15 13 1 13 9 7 13 9 0 13 9 13 15 15 9 13 7 0 9 13 1 9 9 13
12 16 0 13 15 15 13 15 13 1 9 0 13
17 13 13 0 0 9 9 15 7 15 1 9 13 7 9 1 9 13
12 0 9 3 0 9 9 9 7 13 1 9 13
39 11 16 0 15 0 9 13 13 13 16 16 13 9 13 9 9 13 3 13 9 3 12 15 11 11 1 15 3 13 13 15 1 13 9 1 9 1 9 13
14 15 0 9 13 15 9 7 9 13 13 0 1 15 13
11 3 15 3 3 7 9 13 15 1 9 13
11 0 9 9 1 9 13 1 11 1 9 13
25 0 11 9 9 15 3 13 13 15 7 1 9 13 13 16 0 9 9 0 9 9 9 13 3 13
16 15 0 9 13 3 1 0 9 9 13 15 15 0 1 9 13
39 15 1 9 16 13 13 9 3 12 7 1 9 13 9 15 11 1 11 13 13 13 9 9 13 3 3 3 0 15 9 13 7 16 15 13 13 9 13 13
14 16 0 9 13 15 13 3 1 9 9 3 12 12 13
11 15 9 13 11 15 1 9 9 15 9 13
18 16 3 9 15 1 9 13 9 13 9 9 13 0 7 15 9 13 13
19 11 0 9 11 11 9 1 0 9 15 1 11 13 1 9 15 9 13 13
22 15 16 1 9 9 3 15 13 3 13 15 9 0 9 13 13 15 3 1 9 11 13
33 3 11 11 7 11 11 9 15 1 9 9 9 13 15 15 9 13 9 13 9 13 16 9 15 15 1 0 9 13 15 1 11 13
8 3 12 3 9 1 11 9 13
2 0 13
13 0 9 13 1 9 11 9 12 9 1 9 13 13
31 11 11 11 11 9 13 1 9 11 1 11 3 3 13 13 9 13 15 9 13 16 3 0 13 9 9 13 0 7 13 13
30 1 9 13 9 7 3 13 0 3 15 1 15 9 13 13 7 0 3 3 16 1 0 9 9 3 0 3 9 13 13
14 1 9 1 9 9 13 3 0 3 15 1 0 13 9
11 0 15 0 13 13 15 1 9 3 9 13
17 15 9 11 0 13 1 11 13 16 1 9 0 9 9 9 13 13
12 3 16 13 9 9 13 0 7 1 9 13 13
26 15 9 13 9 9 1 15 13 15 13 15 0 9 0 13 9 15 7 0 13 13 15 9 1 9 13
13 13 9 15 11 9 13 15 7 1 0 9 13 13
8 16 3 13 15 9 9 13 13
15 0 13 9 9 7 13 1 0 11 13 7 3 1 9 13
38 3 16 13 13 15 9 0 9 9 1 0 15 9 9 3 12 0 9 15 3 13 9 7 0 12 13 13 3 7 3 13 1 0 16 0 9 13 13
9 0 9 15 3 13 13 13 9 13
28 15 1 9 0 12 7 9 12 1 9 9 13 16 0 3 7 1 9 13 3 7 9 13 9 7 0 13 13
19 0 9 3 3 0 11 9 13 0 7 13 9 9 11 7 3 3 13 13
12 1 0 9 12 1 9 1 15 13 11 7 11
15 1 15 0 16 3 1 11 9 7 9 13 13 1 15 13
21 15 15 7 15 1 9 13 3 7 1 9 9 0 13 13 15 7 1 9 13 13
44 7 16 3 15 9 1 0 9 7 9 11 13 7 9 15 9 13 1 11 13 7 1 15 3 9 1 15 13 13 16 9 13 3 13 13 16 1 15 13 11 9 1 11 13
23 3 13 9 1 15 9 15 7 16 11 13 1 15 1 9 13 15 9 7 9 15 9 13
37 11 16 13 15 1 9 15 13 15 7 15 9 1 13 9 13 3 16 9 1 9 13 13 15 1 0 9 9 13 11 1 15 1 12 9 13 13
21 0 13 1 15 9 0 7 15 15 15 3 13 13 11 13 7 13 16 1 9 13
38 9 3 3 9 9 1 15 13 0 3 11 13 16 3 9 15 1 15 13 13 3 0 13 13 15 9 1 15 3 3 13 15 3 0 1 15 9 13
24 15 13 9 3 11 15 9 1 15 13 7 15 3 1 0 1 15 9 13 0 3 0 9 13
10 0 9 13 11 1 9 11 1 9 13
21 3 13 12 9 15 1 9 13 13 9 13 9 13 3 13 7 3 3 13 13 13
25 1 15 0 15 1 15 9 13 13 1 11 0 9 9 15 1 13 13 16 16 0 13 9 11 13
13 13 3 1 0 11 0 1 15 3 1 15 13 13
21 0 15 1 13 1 0 13 16 15 0 9 0 0 9 0 9 0 1 9 9 13
14 13 3 16 1 9 9 11 13 15 1 11 9 9 13
16 15 9 9 3 13 3 7 13 7 13 9 9 1 11 13 13
7 15 9 1 15 9 11 13
22 0 15 3 9 13 13 16 1 11 13 3 16 0 13 9 13 3 16 9 13 15 13
22 16 15 3 15 13 13 15 9 13 13 9 11 13 13 0 13 7 13 16 1 9 13
17 15 13 9 11 16 15 1 9 11 13 13 0 15 1 11 13 13
3 9 0 13
13 9 13 13 16 15 13 1 9 11 13 0 9 13
6 0 1 0 1 11 13
33 15 9 13 11 16 0 9 0 9 13 13 7 13 15 9 13 11 13 16 3 15 9 13 13 13 16 15 15 7 9 0 13 13
37 3 9 3 12 1 15 9 13 16 9 9 9 13 15 0 9 0 9 1 0 9 13 13 13 9 16 1 9 11 13 9 3 3 15 15 9 13
11 3 0 13 9 9 9 7 13 1 9 13
15 3 15 13 9 11 1 9 9 1 9 0 11 9 13 13
21 0 3 13 13 7 15 9 13 15 7 9 13 13 3 13 0 15 0 7 13 9
8 0 3 13 13 13 9 7 13
7 3 9 9 1 11 15 13
6 0 13 0 3 12 12
20 0 1 9 11 0 11 9 13 1 11 11 11 11 11 11 11 9 9 13 13
65 3 1 11 11 9 13 16 0 1 9 1 9 9 0 9 13 15 1 0 11 9 9 13 1 9 13 7 1 15 13 13 0 13 3 1 0 9 1 9 11 13 0 13 11 9 16 16 15 13 1 9 9 13 3 3 15 0 9 13 7 3 0 13 9 13
45 15 16 11 7 9 0 7 9 13 3 13 1 15 9 12 1 13 9 7 13 7 13 9 13 7 15 9 9 15 1 11 11 13 7 9 7 9 13 15 9 0 9 7 9 13
9 0 0 9 13 7 9 13 3 13
13 13 0 9 9 13 1 15 13 9 7 1 9 13
6 11 15 9 7 9 13
44 15 9 13 11 16 3 9 13 13 9 9 9 13 0 15 9 13 1 9 9 1 9 3 13 7 1 9 0 7 9 9 13 1 9 9 0 9 13 3 15 1 9 13 13
44 3 3 9 13 0 12 13 9 1 0 1 9 9 13 7 16 0 7 13 7 13 13 0 9 7 9 9 13 7 15 9 9 13 13 7 9 1 9 13 7 9 15 13 13
9 0 3 13 9 3 1 9 9 13
30 9 11 0 9 3 13 13 16 0 1 9 9 9 7 13 9 9 7 9 0 13 13 16 15 13 13 9 11 9 13
17 0 9 1 9 13 0 9 1 9 1 9 13 0 7 9 3 13
14 13 15 9 11 15 0 0 9 13 13 1 9 9 13
10 3 9 13 9 7 13 9 1 11 13
9 13 1 9 15 3 13 1 9 9
18 3 11 13 9 13 9 9 7 13 16 0 9 13 9 3 9 13 13
7 9 13 12 0 9 13 13
13 3 9 9 9 7 13 13 9 9 15 13 1 9
7 13 9 11 9 7 13 9
15 0 9 11 13 0 7 9 7 9 1 9 9 7 11 13
23 11 1 9 9 15 1 13 13 16 15 7 1 0 9 7 1 0 15 13 9 9 13 13
21 13 9 0 9 9 0 9 9 7 13 15 0 1 11 1 9 1 11 9 3 13
6 1 0 13 9 11 13
8 3 1 9 13 9 1 9 13
23 0 3 0 13 9 13 16 15 9 13 16 13 9 7 15 1 9 13 7 1 0 13 13
8 15 1 9 0 12 1 9 13
16 0 15 13 9 9 9 0 1 9 9 7 13 15 7 3 13
17 11 13 9 1 11 11 9 7 11 11 9 3 7 13 9 13 3
4 9 9 7 13
11 15 9 13 9 9 1 15 9 13 9 13
17 0 9 13 9 15 9 13 13 16 7 11 7 15 9 9 15 13
12 0 13 9 11 9 1 9 9 9 1 9 13
39 16 0 1 11 13 9 0 13 9 9 7 9 11 1 12 9 15 1 15 9 13 13 13 3 7 1 15 3 3 9 9 13 16 12 13 9 9 11 13
10 13 9 1 12 9 12 9 9 13 13
32 11 9 13 9 13 9 15 13 15 13 9 9 12 9 9 13 1 12 9 0 7 9 1 9 13 7 12 9 13 9 9 13
11 13 1 11 7 9 0 9 9 9 7 0
13 0 3 7 0 13 1 9 13 3 7 9 13 13
23 13 3 3 16 9 13 13 15 15 9 7 9 1 0 3 13 7 0 9 0 9 9 13
17 3 0 1 9 13 16 1 0 0 9 9 0 0 9 13 9 13
6 0 9 9 0 9 13
13 0 3 1 9 1 9 1 0 9 9 1 9 13
51 3 9 0 1 9 13 16 9 13 1 15 16 0 9 1 9 13 0 13 13 9 9 9 13 3 7 15 13 9 16 0 9 3 0 9 3 13 7 13 13 3 13 9 13 7 0 9 13 9 3 13
15 15 13 13 11 16 15 1 9 13 0 13 9 9 3 13
15 3 13 3 9 7 1 9 15 13 13 13 9 15 13 9
6 9 13 7 0 9 13
21 3 9 1 9 13 9 7 13 13 7 0 9 9 1 9 13 0 9 1 9 13
27 0 3 1 9 15 13 13 0 9 1 15 13 13 9 3 13 3 13 7 0 9 1 9 13 0 9 13
14 15 11 9 13 0 9 13 0 13 0 3 9 9 13
11 3 9 15 9 13 13 9 9 15 9 13
13 1 0 9 11 15 9 9 13 13 15 1 9 13
13 11 15 1 9 13 1 9 13 9 7 9 13 13
13 11 16 1 9 1 9 13 12 1 9 11 13 13
9 15 12 13 16 9 1 15 9 13
11 13 7 13 9 0 9 9 0 9 9 13
19 0 1 9 1 9 9 13 16 15 1 0 3 9 13 0 9 9 7 13
33 9 15 3 9 13 7 1 9 13 13 15 9 1 15 9 13 15 13 3 7 1 15 9 9 1 9 13 3 7 1 15 9 13
15 13 7 13 16 15 13 16 0 9 9 0 1 0 9 13
6 16 0 9 13 13 13
9 13 11 9 13 1 9 9 13 13
3 9 9 13
6 9 9 7 1 9 13
6 0 13 9 9 0 13
4 9 0 9 13
26 9 13 16 9 13 15 7 15 1 9 1 9 13 13 0 7 0 9 9 9 1 0 13 9 13 13
13 13 16 0 9 1 9 13 15 7 1 15 13 13
31 0 13 13 7 0 9 13 13 9 15 16 0 9 1 9 9 13 1 15 15 9 7 9 15 13 3 1 0 9 15 13
8 9 3 13 0 9 15 13 11
13 0 3 3 13 7 1 0 9 13 9 1 9 13
9 1 0 9 9 9 9 9 13 13
16 15 7 0 9 9 3 13 13 16 15 1 9 1 0 9 13
18 15 3 15 13 7 13 3 13 3 7 3 16 13 15 1 15 13 9
8 0 0 9 13 1 9 0 11
8 3 15 9 13 13 1 12 9
12 16 11 1 11 13 0 9 0 13 9 0 9
32 15 16 1 15 3 13 16 0 9 3 13 1 9 0 7 15 13 9 9 7 11 15 13 15 7 1 15 0 9 9 7 13
52 9 3 0 13 0 7 15 9 9 13 3 9 13 16 0 9 9 1 9 1 15 13 9 7 1 0 9 9 13 7 3 13 13 15 15 1 9 9 13 7 9 0 9 1 9 13 13 11 7 0 9 13
41 9 11 13 9 9 9 9 13 0 9 13 0 1 11 13 16 15 15 15 1 15 9 13 0 9 7 0 9 15 13 13 0 9 15 9 9 7 13 9 9 13
23 15 16 13 1 11 9 13 15 15 1 0 9 15 9 1 9 13 13 15 9 1 9 13
4 0 0 3 13
7 3 0 7 3 13 9 13
15 0 3 9 9 13 16 3 0 9 13 0 9 9 9 13
14 1 15 11 0 9 15 15 13 9 7 9 9 13 12
14 3 9 3 9 13 9 15 15 13 1 15 15 13 9
10 1 0 0 15 13 9 15 9 1 9
10 7 1 0 12 9 0 13 9 0 9
15 1 0 0 9 9 9 9 13 0 7 0 13 1 15 9
27 3 3 1 15 9 0 0 7 13 7 16 15 13 9 13 16 9 13 16 1 9 1 9 9 13 0 13
4 9 9 7 13
12 16 15 7 0 7 9 15 9 3 13 9 13
6 0 9 1 15 13 0
3 0 15 13
11 9 15 9 7 13 16 15 1 9 9 13
11 3 7 15 13 9 13 3 7 9 15 13
17 0 13 7 16 15 1 0 13 9 13 7 16 13 0 0 9 9
6 3 3 9 1 9 13
17 15 0 9 9 1 9 9 15 9 0 11 0 13 13 1 9 0
13 3 15 3 15 9 13 13 15 7 9 9 7 13
12 9 1 9 13 13 3 7 9 3 1 0 13
16 0 13 9 7 15 9 0 1 9 13 7 1 9 9 7 13
6 0 3 9 9 13 13
7 3 9 0 0 1 9 13
25 15 15 12 1 9 13 13 16 3 7 1 9 9 13 13 3 7 15 15 13 9 13 3 9 13
13 3 3 0 13 16 9 9 9 1 13 7 9 13
26 1 0 0 13 13 3 13 9 7 1 15 1 9 13 1 15 7 0 3 1 9 13 13 9 9 13
4 0 9 13 9
45 15 16 13 9 7 15 9 13 15 3 1 11 9 3 13 13 16 7 0 9 13 7 13 13 15 1 9 13 7 15 16 15 13 9 9 7 0 3 0 1 15 9 9 7 13
6 0 12 9 9 7 13
61 0 13 15 9 3 0 0 7 1 0 9 15 13 13 0 0 15 7 1 9 9 7 13 7 1 9 9 13 7 15 13 13 9 7 1 0 0 9 13 16 1 9 9 16 9 9 13 3 13 9 0 9 13 13 3 7 0 9 13 13 9
12 15 0 9 9 13 15 13 9 9 0 9 13
17 9 15 15 1 9 7 9 7 15 9 13 13 0 9 0 13 13
11 7 16 0 9 9 13 3 1 0 9 13
4 0 13 0 9
5 0 15 9 9 13
5 0 9 7 9 9
10 0 1 9 9 9 7 13 9 0 13
9 1 0 11 7 11 7 11 7 9
9 1 0 0 3 15 0 9 13 9
11 0 16 9 13 13 15 15 9 13 3 13
11 0 1 9 0 9 13 9 9 0 13 13
26 3 7 3 13 16 13 15 9 7 13 1 15 13 7 13 13 13 0 7 0 9 9 1 9 13 13
14 9 15 15 1 11 9 0 13 15 7 1 9 13 13
12 1 0 9 9 15 9 3 9 9 7 9 13
13 9 0 7 9 7 9 9 3 13 16 9 9 13
38 1 0 9 9 0 3 1 0 13 16 15 9 3 1 13 16 9 9 13 13 1 1 15 13 3 13 9 7 0 9 1 0 1 9 9 13 0 13
17 9 15 9 1 9 9 9 13 0 1 15 0 9 13 1 9 13
11 9 1 9 3 1 9 9 9 7 13 9
35 7 16 9 0 9 13 13 15 9 13 7 1 9 16 9 1 9 13 1 9 1 0 9 9 13 7 16 13 13 9 7 15 9 13 13
8 9 13 1 9 9 0 7 0
31 15 7 15 0 9 13 13 1 9 13 3 9 7 3 1 0 9 9 7 9 15 1 15 13 13 13 0 9 13 3 13
54 15 9 3 15 9 9 13 13 13 9 13 16 15 15 1 9 0 1 0 9 7 9 13 16 1 9 13 3 7 1 15 15 13 16 3 9 0 7 0 0 9 13 7 1 9 13 7 1 0 9 9 13 13 13
5 9 15 13 13 13
7 15 13 1 9 13 9 13
9 1 9 0 3 1 9 13 3 13
13 3 3 7 9 13 15 9 0 13 3 7 9 13
17 9 9 15 0 13 15 13 7 15 3 9 13 11 7 11 7 11
5 0 3 9 3 13
10 9 15 1 9 7 1 9 9 0 13
6 1 9 9 7 9 13
9 15 3 0 13 0 1 15 13 9
9 0 9 13 0 9 9 7 13 13
11 1 9 3 0 9 9 13 1 0 13 9
10 3 7 15 9 9 0 7 9 13 0
28 7 9 7 9 1 9 0 9 9 7 9 15 3 13 15 7 15 9 13 13 9 13 7 9 3 15 13 13
57 0 9 0 13 9 16 0 9 13 9 9 13 9 13 16 0 9 13 13 0 7 0 9 13 16 3 1 9 7 9 13 13 16 15 13 9 9 15 1 9 9 9 7 13 16 9 9 9 13 16 15 15 9 1 0 13 13
12 9 0 9 13 3 3 1 15 13 9 9 13
14 0 0 9 13 13 9 0 13 3 7 15 3 13 13
10 3 0 15 13 0 13 0 9 9 13
20 16 9 9 7 13 13 7 13 9 15 0 9 13 7 9 9 7 13 9 13
20 9 15 13 9 15 1 9 15 9 13 7 15 9 13 7 9 13 9 13 13
19 15 1 0 13 3 13 1 9 7 9 9 13 15 7 0 9 3 9 13
5 9 13 9 3 13
10 15 15 1 9 1 15 13 1 9 13
2 0 13
8 0 7 15 9 13 9 7 13
22 7 13 3 9 16 9 9 9 13 3 9 13 1 9 9 9 7 9 1 11 9 13
17 15 9 1 0 9 0 9 15 13 0 7 13 9 7 0 9 9
17 3 16 1 0 9 9 9 15 3 9 13 0 9 7 9 9 13
15 3 13 13 0 7 13 9 3 15 3 0 1 0 9 13
13 0 11 9 15 3 13 13 9 12 9 9 0 13
10 3 3 3 13 13 3 7 9 9 13
19 13 1 9 7 9 7 9 9 0 7 9 11 9 13 1 9 9 7 9
15 3 15 13 3 0 1 9 9 0 7 9 9 1 9 13
15 0 7 1 15 9 9 13 13 15 0 1 9 13 3 13
13 1 15 15 3 13 1 0 7 9 13 13 0 13
23 13 9 9 9 15 1 0 9 1 9 12 9 13 0 3 7 0 0 15 15 0 13 9
6 0 13 9 9 7 9
5 0 9 9 7 9
5 13 3 15 13 9
40 0 13 0 9 9 7 9 9 7 9 3 13 0 7 13 9 7 9 1 9 9 7 13 3 7 9 9 13 3 7 16 15 13 9 13 13 15 7 13 13
11 1 15 15 13 7 3 3 3 13 9 13
29 15 1 9 16 13 13 1 9 3 15 13 13 15 0 9 7 1 9 13 7 13 9 3 16 9 9 15 13 13
13 3 16 15 9 13 0 9 9 13 7 3 0 13
7 0 13 9 15 15 9 13
6 9 7 9 7 9 9
16 0 9 15 13 7 0 9 3 7 9 3 7 9 15 13 13
5 0 3 9 13 13
11 7 13 1 9 7 13 3 0 3 13 13
12 9 9 7 9 7 9 3 1 15 9 9 13
14 0 3 13 1 9 9 13 7 1 0 9 1 9 13
27 11 16 1 9 9 13 9 15 1 9 13 9 9 13 16 3 1 13 3 15 9 9 13 13 3 13 3
49 7 16 3 9 9 15 9 13 7 16 15 9 13 13 9 9 0 9 15 9 9 13 1 9 9 12 13 7 1 0 9 9 9 12 13 9 7 9 12 9 13 9 13 0 7 0 9 9 13
28 15 16 13 9 13 1 9 11 13 1 11 9 11 11 11 1 15 9 13 16 15 9 9 7 9 9 13 13
14 13 16 9 1 9 13 13 16 15 15 9 3 9 13
5 11 3 13 13 13
12 3 1 7 15 9 13 9 0 1 9 0 13
14 15 9 1 0 11 13 15 1 9 1 0 9 13 13
11 3 3 1 15 9 3 1 9 0 13 9
44 3 3 0 13 9 16 1 15 0 3 7 0 13 3 7 15 9 1 15 13 16 9 7 9 13 3 0 13 9 15 0 9 15 1 15 13 13 9 9 7 13 15 13 9
35 7 0 13 13 16 9 13 9 3 13 3 9 9 15 13 9 9 3 9 7 9 13 9 9 9 7 15 0 1 9 3 9 15 9 13
3 13 9 13
27 11 9 15 9 3 3 13 16 9 13 3 13 7 9 13 7 0 9 9 13 16 0 9 13 13 0 13
10 7 3 13 1 9 9 15 15 13 13
10 15 9 1 11 9 9 1 0 9 13
12 15 0 11 13 0 9 15 13 15 9 13 13
11 0 1 15 9 13 15 15 7 15 0 13
42 11 9 0 9 9 15 3 1 11 9 13 9 3 13 16 9 9 7 9 13 3 13 15 9 13 11 15 0 9 9 13 9 15 0 1 11 11 7 9 13 15 13
37 9 9 7 1 9 7 9 9 15 13 1 9 9 7 9 1 11 13 13 16 15 1 9 9 13 16 7 15 9 15 13 1 11 12 13 9 13
8 16 3 13 9 15 15 13 13
11 3 9 1 12 9 13 9 15 9 11 13
4 15 9 9 13
14 0 3 13 1 0 9 9 3 11 7 11 13 9 13
17 0 3 0 9 9 13 3 16 0 9 9 0 13 16 9 9 13
14 9 9 9 0 13 12 1 15 15 3 13 1 11 13
12 0 9 9 7 11 11 11 13 12 7 9 13
18 13 9 11 11 1 9 12 1 11 3 1 15 9 15 9 13 13 13
24 15 1 0 12 1 9 11 15 13 1 11 0 7 11 9 13 13 3 1 0 9 13 11 13
19 13 1 9 0 15 13 13 15 1 9 0 9 15 1 9 13 9 13 13
27 11 11 7 13 16 9 0 9 13 13 1 0 9 13 16 3 13 9 13 7 9 9 15 9 9 13 13
21 13 3 3 13 9 0 15 3 9 3 9 15 15 9 13 7 1 15 9 13 9
18 3 15 7 9 0 7 9 0 7 9 0 9 9 7 9 15 13 13
30 0 9 9 13 0 0 7 9 9 13 3 1 9 9 13 15 3 13 0 1 13 7 13 9 13 7 1 0 9 13
9 15 3 1 9 9 1 9 9 13
16 3 7 9 9 0 3 13 7 9 0 0 7 9 0 13 13
28 3 1 0 9 9 3 9 13 13 13 16 3 1 13 15 13 16 15 9 1 13 13 3 1 15 9 9 13
6 13 1 0 9 9 11
30 15 13 9 9 1 13 9 16 3 1 9 9 9 3 0 9 13 3 16 0 9 13 1 0 9 9 7 9 9 13
5 0 3 9 3 13
20 0 1 15 9 9 13 9 7 13 0 15 1 9 11 1 9 9 7 13 13
12 3 3 1 9 9 13 7 15 13 9 13 13
15 13 7 13 9 3 13 9 13 15 15 0 3 9 9 13
19 13 9 12 12 9 15 13 0 11 1 15 13 1 9 9 7 9 3 13
4 0 9 9 13
5 0 1 9 13 13
8 0 9 9 15 13 0 9 13
4 13 9 3 13
11 3 0 9 1 9 9 7 13 3 9 13
8 15 1 9 13 11 1 9 13
18 7 12 1 9 15 15 13 0 0 7 0 13 9 15 13 3 13 0
5 12 9 11 13 13
16 9 0 13 16 3 9 3 13 13 3 7 15 13 1 9 13
10 13 9 9 15 13 13 9 1 0 13
10 15 11 13 13 0 9 15 0 9 13
100 11 15 15 0 9 9 11 1 0 9 9 1 9 13 7 3 9 3 15 1 9 13 9 13 0 9 13 1 9 9 11 9 13 16 3 9 13 3 7 15 1 9 15 9 13 3 15 13 9 15 0 9 3 9 13 16 3 1 9 13 3 13 15 15 9 9 13 15 12 13 9 0 7 9 13 7 3 13 9 1 12 9 12 13 13 12 9 13 1 0 9 13 15 1 7 9 12 3 9 13
8 0 13 1 9 1 9 0 13
46 0 0 9 9 9 9 13 3 7 0 0 15 13 9 1 0 9 1 9 13 13 3 3 13 13 13 1 15 9 9 16 9 13 3 3 16 15 1 9 13 9 13 15 9 3 13
13 0 15 9 0 13 7 3 0 9 9 1 9 13
10 13 9 1 0 9 16 15 9 13 13
9 0 9 9 0 1 15 9 7 13
10 0 13 9 7 15 1 15 9 9 13
13 3 7 3 9 13 3 7 15 1 9 15 13 13
5 15 9 3 13 13
20 0 0 15 1 9 9 13 11 7 7 11 9 15 1 0 9 13 1 9 13
15 0 9 15 13 13 9 9 3 1 9 13 15 13 3 9
12 13 13 15 7 0 13 16 0 9 1 9 13
25 13 0 1 9 13 11 11 11 15 0 9 1 11 13 15 9 0 9 13 7 9 3 0 9 13
9 13 13 9 7 1 0 9 13 9
8 13 9 1 0 7 1 9 13
9 13 0 9 0 9 15 1 9 13
6 13 9 11 0 13 9
5 3 1 9 13 13
16 0 9 13 0 15 13 3 16 1 9 13 13 9 7 9 13
7 3 13 9 9 15 9 13
2 13 9
8 3 3 15 9 13 15 13 13
13 3 13 7 9 0 0 1 9 9 9 7 9 13
8 15 13 3 0 16 9 9 13
6 9 9 3 13 9 13
10 13 3 9 13 15 3 13 1 9 13
8 3 13 9 1 15 9 9 13
5 9 1 9 9 13
9 3 3 13 15 1 9 9 7 13
7 15 9 13 16 3 13 13
10 15 16 1 9 13 7 0 15 13 9
11 0 0 3 13 9 15 1 9 3 13 13
25 3 1 15 13 9 11 11 9 0 15 15 13 13 1 0 9 13 0 7 1 12 15 1 9 13
10 0 13 9 9 7 0 9 9 9 13
43 3 15 15 1 9 13 15 3 3 9 9 0 13 3 7 1 0 15 13 9 13 3 7 0 15 13 15 9 9 7 13 13 13 7 15 1 9 13 13 0 1 9 13
27 9 15 0 1 0 9 0 9 9 9 1 0 13 9 0 9 13 16 3 13 9 0 9 13 3 13 13
12 9 9 0 9 13 9 1 9 0 1 9 13
28 7 0 13 3 1 9 9 9 16 0 9 16 11 11 13 1 9 1 9 13 9 3 13 13 1 0 11 9
27 3 15 9 9 13 16 3 13 9 13 15 9 9 15 1 9 13 13 3 7 0 9 9 9 13 13 13
5 15 9 11 9 13
41 13 0 9 9 3 13 12 16 9 9 13 13 13 3 0 3 9 9 13 13 3 9 1 0 9 9 13 13 3 3 3 16 3 1 0 9 9 7 9 0 13
25 15 15 9 3 13 13 16 9 15 0 9 11 13 16 11 9 13 1 9 9 13 0 11 9 13
17 11 3 1 13 9 13 9 0 13 9 1 0 9 1 15 9 13
9 15 9 7 15 9 15 15 13 13
5 9 1 15 9 13
85 7 3 1 0 9 13 13 0 1 15 9 13 9 16 3 13 1 15 11 1 9 13 9 3 3 3 13 1 9 13 16 9 13 13 7 0 9 13 15 15 0 1 11 9 13 13 3 9 9 13 3 7 3 1 0 9 13 13 7 0 9 7 9 15 13 7 3 13 15 9 9 7 13 3 0 9 9 3 12 15 0 9 15 13 13
42 0 9 13 9 9 11 12 9 9 11 9 13 9 7 1 0 9 11 13 1 9 9 7 9 9 13 13 7 1 11 15 0 0 9 13 0 9 13 9 0 9 13
4 0 9 13 13
36 15 16 9 7 9 13 12 9 1 9 9 12 1 9 12 0 1 9 9 11 1 9 13 9 7 9 13 3 13 1 11 1 9 13 13 13
7 3 1 15 11 9 9 13
16 9 1 9 9 15 11 1 9 13 9 9 9 7 9 9 13
15 16 0 9 13 3 13 15 9 13 0 13 9 13 15 9
17 9 15 15 15 0 9 13 13 0 9 9 13 15 3 9 13 13
13 3 9 13 9 3 0 9 15 13 0 0 0 9
10 3 0 3 13 3 16 15 15 13 13
12 3 15 13 15 13 16 0 13 0 15 9 13
23 15 3 9 13 13 13 0 0 9 15 15 9 1 0 9 13 11 13 1 9 9 0 3
11 9 15 0 13 13 11 7 11 7 11 11
8 13 15 1 0 7 13 7 13
8 16 9 13 13 15 3 11 13
10 11 16 13 13 9 3 13 0 13 9
8 1 15 15 3 13 11 0 13
22 11 1 11 13 13 15 3 0 7 1 9 7 9 13 16 15 13 3 13 8 11 13
6 7 0 1 15 15 13
9 15 9 3 13 13 11 13 1 11
24 15 13 3 1 15 15 3 13 15 16 1 15 9 13 0 9 13 13 3 16 9 13 9 0
6 9 0 13 3 13 9
7 16 13 9 9 13 1 15
8 0 13 0 13 0 3 0 9
11 13 15 15 0 13 16 1 15 9 3 13
5 7 0 0 9 13
8 7 13 15 1 15 15 13 13
30 11 9 15 1 11 11 16 0 9 13 13 13 1 15 9 11 11 11 1 0 9 15 15 9 0 9 13 1 11 13
23 3 13 0 9 1 15 13 11 11 7 11 11 7 15 15 13 9 13 16 9 13 11 11
3 3 13 9
7 13 15 11 16 13 1 11
10 9 3 15 13 16 0 11 9 15 13
3 15 13 0
11 13 7 15 7 11 9 0 9 1 15 9
16 3 13 13 3 0 11 9 3 11 1 15 0 3 9 15 13
3 13 0 11
29 3 1 9 0 9 9 3 0 15 1 15 15 11 15 9 13 3 9 0 13 0 13 15 7 9 15 13 7 9
24 3 13 0 15 13 13 3 13 7 3 9 0 13 7 3 3 1 13 15 0 9 9 3 13
32 1 15 13 16 15 0 13 7 15 13 9 13 13 16 3 9 0 9 0 15 9 13 16 15 15 15 9 7 9 1 15 13
11 3 16 13 1 15 13 0 9 13 15 13
17 13 3 1 15 9 13 7 3 15 9 3 3 13 3 3 13 13
5 13 15 15 9 13
3 13 3 3
3 3 15 13
13 11 11 11 11 11 11 9 9 15 13 13 0 11
6 1 15 3 3 15 9
9 15 1 15 1 15 9 13 3 3
7 0 9 11 9 15 13 13
11 13 16 13 13 0 0 15 13 1 9 9
5 16 3 13 3 13
14 3 3 0 9 13 9 15 9 0 9 0 9 15 13
11 1 15 9 15 13 0 15 15 9 13 13
9 3 0 9 3 13 13 16 11 13
25 9 15 13 9 15 13 13 7 3 16 13 13 16 0 1 9 3 13 7 1 9 0 9 3 13
10 0 9 9 1 15 11 11 13 13 13
17 15 3 15 1 9 0 13 1 15 9 7 1 9 15 1 15 13
9 9 15 15 13 15 13 1 11 13
8 3 7 3 13 11 9 15 13
5 13 15 1 9 13
12 15 3 13 16 15 1 15 3 0 7 13 13
21 15 1 15 3 13 1 15 9 13 13 7 13 13 15 7 0 1 9 13 9 0
13 15 1 9 16 13 15 13 3 1 15 16 13 13
9 11 0 13 1 15 0 9 3 13
11 0 1 15 13 16 15 15 13 1 15 13
5 0 9 15 15 13
15 3 3 16 3 15 13 13 3 1 15 1 9 0 13 13
14 3 3 13 15 9 15 13 13 13 1 0 9 15 13
4 13 11 9 9
4 15 0 9 13
3 0 9 13
9 0 15 3 11 16 1 15 13 13
9 13 3 0 13 15 3 3 9 13
11 15 3 0 7 0 9 9 1 11 11 13
22 15 16 0 13 3 3 0 9 1 9 9 0 13 13 3 1 15 16 13 13 9 13
10 15 1 15 1 11 13 3 15 0 13
17 13 9 11 0 15 16 7 11 0 15 7 11 0 13 9 0 9
12 3 13 3 13 0 3 9 3 0 0 9 13
8 15 15 3 9 13 15 3 13
8 1 0 13 3 15 3 13 13
5 0 15 1 0 13
12 15 16 13 13 11 9 7 15 9 7 9 13
24 15 9 13 7 15 9 13 13 7 0 7 0 11 9 15 9 1 0 1 15 9 15 13 13
16 3 15 15 15 0 1 9 0 7 9 9 13 13 1 0 13
34 3 3 13 16 15 3 15 0 13 16 7 15 9 13 7 0 15 9 9 7 0 15 7 7 15 9 7 15 9 0 9 9 7 13
26 16 1 15 13 1 9 15 9 13 15 0 15 15 9 13 16 11 9 9 1 15 13 15 15 13 13
23 15 16 13 0 13 0 9 1 15 13 15 7 13 3 9 7 13 3 0 7 13 3 13
21 3 1 15 15 3 3 1 15 1 15 13 13 13 3 13 15 16 7 13 7 13
13 3 3 1 11 15 0 13 13 13 15 13 9 13
15 1 0 3 9 15 15 13 16 3 1 15 9 11 13 13
27 7 13 16 7 9 15 9 13 7 16 15 15 1 15 3 9 13 13 13 11 15 9 1 9 3 15 13
33 3 16 0 9 9 15 11 13 15 9 9 15 0 13 13 3 15 0 13 13 1 15 1 0 9 16 0 13 15 13 0 0 13
24 7 1 15 0 15 15 13 12 15 13 9 13 13 16 7 9 1 13 3 7 9 13 0 13
27 15 13 3 16 15 9 1 15 13 0 1 15 13 13 13 15 13 3 7 15 13 7 13 0 15 9 13
9 15 3 15 13 13 1 15 3 13
22 15 16 1 15 13 13 15 3 7 0 13 13 3 15 13 3 7 0 13 3 15 13
21 1 0 9 15 1 11 13 13 15 3 13 15 13 3 15 13 16 9 9 13 13
5 0 9 13 15 13
20 15 15 13 7 15 15 13 13 15 0 13 3 13 13 15 1 9 15 13 13
12 3 15 1 15 9 7 9 12 0 1 9 13
4 11 9 3 13
5 11 0 9 9 13
14 13 16 13 7 15 13 7 15 13 15 1 15 3 13
10 3 13 3 16 15 13 1 9 9 13
12 15 3 13 1 0 9 16 0 1 0 15 13
13 15 15 13 13 16 15 3 0 9 1 9 15 13
27 11 9 3 15 13 15 13 9 13 1 11 7 1 15 3 1 0 9 13 7 15 1 13 9 8 11 11
4 9 15 13 3
7 0 13 3 15 15 13 13
14 15 0 3 13 16 15 3 0 3 3 16 3 13 13
14 15 13 15 1 9 7 15 13 13 13 15 3 3 0
9 1 9 3 13 15 7 15 9 13
7 11 11 3 13 15 13 3
16 15 9 9 15 15 16 1 9 13 13 13 1 15 9 13 13
5 1 15 13 3 13
10 9 15 7 9 1 15 11 7 9 13
24 15 15 13 1 15 9 15 13 13 7 13 0 9 13 16 0 13 3 13 3 1 15 3 13
18 15 15 1 0 9 13 13 15 15 11 7 0 13 13 7 0 9 0
13 0 15 9 9 6 0 7 15 0 3 15 13 13
13 0 16 15 15 13 13 3 15 15 13 13 13 13
12 11 11 3 1 9 0 3 15 1 15 13 13
35 3 13 7 15 7 9 7 0 15 15 0 9 7 15 9 7 15 9 13 13 3 0 3 3 7 13 7 3 15 15 9 9 7 13 13
16 3 1 0 9 3 9 13 16 1 15 13 1 15 3 13 13
11 11 9 15 15 9 13 7 15 3 9 13
7 15 3 13 3 13 3 13
31 3 3 15 1 15 9 13 16 7 3 15 3 13 15 11 13 3 15 15 11 7 0 15 13 15 13 11 3 15 15 11
25 3 1 0 9 15 0 0 0 9 13 16 16 0 13 3 13 13 0 15 0 9 1 0 9 13
11 9 0 7 9 1 15 1 15 13 3 13
16 15 0 9 13 0 11 15 15 13 16 13 13 7 9 15 13
6 15 8 3 13 15 13
7 13 1 15 16 0 3 13
9 11 15 13 7 15 15 9 8 8
44 16 13 1 0 13 0 15 1 0 15 16 13 1 11 3 3 16 3 13 11 9 1 9 15 13 9 15 1 15 13 13 13 7 0 0 9 1 9 13 15 15 1 15 13
14 3 13 13 16 9 15 13 15 9 9 3 0 13 13
11 3 15 1 15 9 13 7 3 3 13 13
28 15 15 16 15 9 3 13 3 3 3 7 13 3 7 13 1 0 3 16 0 1 9 9 0 9 15 13 13
8 0 15 13 13 3 0 13 13
12 3 3 13 0 1 15 13 16 15 9 0 13
14 3 9 15 13 15 1 9 9 13 13 7 9 0 12
9 9 15 13 15 13 16 0 9 13
12 3 15 15 15 9 3 13 16 0 9 9 13
10 1 9 13 3 13 16 3 13 7 13
5 0 9 13 0 9
6 3 0 16 9 0 13
45 1 9 15 7 15 15 13 13 7 15 3 0 0 9 15 15 13 13 15 3 3 3 13 1 15 7 13 16 13 3 3 13 15 15 13 15 13 13 0 9 3 15 15 13 9
24 15 3 15 7 13 1 15 7 13 16 15 16 15 13 13 3 3 15 0 7 1 15 13 13
4 11 15 9 13
3 9 15 13
19 7 15 9 13 3 7 3 12 9 15 3 1 0 9 13 0 9 13 13
16 3 13 9 0 11 16 13 3 3 1 11 1 15 0 9 13
23 7 16 15 13 3 3 0 9 15 15 13 1 15 13 3 13 3 3 9 3 13 13 9
70 16 13 0 3 0 15 9 7 15 15 3 3 3 13 13 15 9 13 3 13 15 3 15 3 1 9 15 13 15 3 7 9 15 3 7 15 9 3 13 3 13 3 15 0 3 3 9 7 15 9 0 0 13 16 3 0 13 0 15 16 15 13 7 16 9 15 13 13 3 13
36 7 16 0 13 3 16 15 3 13 15 1 9 15 13 0 1 15 9 13 3 0 13 13 0 13 3 15 13 0 9 0 7 1 0 9 0
5 3 0 13 1 11
9 15 13 15 11 15 13 3 3 13
11 3 3 0 9 3 3 9 7 3 9 13
6 9 3 15 13 15 13
5 15 15 3 13 13
10 0 15 15 9 13 3 9 3 0 9
13 15 15 0 13 3 0 9 3 0 13 13 3 13
7 13 1 11 11 11 13 13
13 7 16 1 0 0 13 15 15 0 0 0 0 13
2 9 13
2 11 13
3 8 7 8
5 7 13 3 8 8
18 3 15 0 9 13 3 11 13 11 13 13 0 7 9 13 9 1 9
12 3 13 0 16 0 15 9 13 13 15 16 13
12 9 15 13 3 0 9 11 13 9 7 9 15
13 3 13 3 13 3 7 3 13 7 3 15 9 13
2 0 13
1 13
12 13 7 9 0 16 15 9 13 1 0 9 13
7 0 9 11 9 11 11 13
5 11 15 0 13 13
4 9 11 3 13
26 11 11 11 9 13 15 13 1 9 0 13 9 11 11 16 1 9 13 15 7 1 9 9 13 7 13
6 15 15 3 13 3 13
13 15 3 1 15 13 3 13 7 6 13 1 13 0
16 3 9 0 9 15 11 13 15 7 3 3 9 9 13 13 13
6 15 13 3 1 15 13
6 3 11 11 11 11 9
5 13 15 12 3 9
10 12 1 11 11 15 11 3 13 15 13
7 0 15 15 0 15 9 13
15 15 13 15 3 9 9 13 3 9 13 9 3 0 9 9
18 15 9 13 3 1 15 13 1 13 7 3 13 0 16 3 13 0 9
14 15 3 15 13 15 9 3 0 13 13 16 15 9 13
32 15 3 15 13 13 1 11 15 9 3 13 1 11 13 13 3 7 3 15 0 0 13 3 1 11 13 7 15 1 11 9 13
13 3 3 7 0 9 3 7 0 3 0 9 13 13
25 13 3 1 9 1 15 15 9 0 9 15 7 3 13 0 9 9 16 7 13 7 13 7 13 13
25 3 3 13 3 15 3 13 13 9 13 7 13 15 9 9 15 7 13 9 3 7 15 0 13 13
36 13 3 7 1 13 9 0 0 7 1 9 1 9 0 13 3 0 9 13 7 0 0 1 13 9 13 9 3 9 7 9 3 3 13 9 9
6 0 16 3 0 13 11
17 9 3 0 0 9 3 0 3 9 9 0 0 15 3 1 9 13
5 15 13 1 9 0
3 13 1 9
16 1 15 15 13 0 9 0 16 3 13 15 13 0 16 3 13
13 15 3 9 7 1 15 0 7 9 0 7 9 0
6 15 3 3 1 15 13
9 7 13 16 0 15 13 13 13 3
9 15 13 9 16 15 3 15 15 13
7 3 1 9 9 9 9 13
4 9 11 9 13
25 1 0 9 11 9 11 11 13 9 13 16 0 9 15 0 13 7 13 1 9 9 7 1 9 13
5 11 3 3 13 3
7 0 9 9 11 13 1 9
2 9 13
10 15 3 0 15 0 1 9 13 3 13
15 13 16 0 13 1 0 13 1 0 0 9 0 9 9 13
25 15 3 0 9 13 3 15 13 1 15 15 1 15 13 16 3 13 13 13 13 15 3 13 3 13
1 13
1 13
2 3 13
7 3 7 3 16 0 13 13
2 15 0
2 15 0
2 15 0
2 15 0
2 15 0
7 7 0 1 15 13 3 3
20 3 3 7 3 15 3 13 13 7 0 9 9 15 13 9 0 1 9 3 13
5 9 9 3 13 13
6 9 3 13 9 3 13
9 8 15 13 11 7 9 13 9 15
11 3 3 16 1 15 13 13 3 15 8 13
6 1 0 9 0 13 15
9 9 15 13 16 15 9 15 8 13
4 0 15 15 13
1 15
1 3
6 9 9 0 9 13 3
1 13
10 11 0 0 9 13 7 3 13 1 9
3 15 0 13
5 1 15 0 9 13
6 3 11 11 11 11 9
27 13 16 0 13 13 1 15 3 13 13 7 3 3 13 16 0 3 0 9 9 13 7 0 13 1 0 9
9 0 9 11 15 13 13 1 15 3
2 0 0
3 0 3 0
2 3 13
12 3 11 9 9 0 9 9 11 1 9 13 11
15 9 13 1 9 0 7 13 1 0 0 9 0 9 9 8
15 13 1 15 13 3 15 9 1 9 13 15 9 0 9 13
9 15 3 13 1 0 9 1 9 13
16 3 11 9 1 9 1 11 13 15 1 9 7 1 13 9 13
28 13 3 13 1 9 16 15 0 9 9 8 13 15 7 16 13 13 15 13 3 1 15 3 1 0 9 13 13
52 11 16 13 0 13 9 1 15 16 0 13 9 15 9 15 13 13 3 7 1 15 9 13 13 3 3 13 15 16 13 9 16 9 16 0 16 13 15 9 13 3 9 3 9 3 9 13 3 15 9 15 13
24 0 0 9 15 15 3 15 9 15 15 11 13 13 13 1 9 1 9 13 0 8 3 3 13
3 0 11 13
40 13 9 13 3 11 13 15 9 15 15 13 7 13 0 9 15 15 3 0 9 13 1 15 3 15 15 9 0 3 3 13 16 15 15 9 1 11 9 13 13
17 0 9 15 3 11 13 7 3 1 0 3 3 15 13 13 3 13
2 15 0
1 9
21 3 0 13 8 1 9 9 1 0 9 1 9 11 1 13 9 9 1 9 1 9
7 13 3 1 0 9 9 15
6 0 3 15 9 3 13
3 9 8 8
2 15 0
2 15 0
24 3 16 9 13 9 1 9 9 13 13 0 9 0 0 9 11 9 9 11 7 9 16 13 13
8 11 3 9 9 9 0 13 9
4 9 0 9 13
8 9 13 3 16 15 13 16 13
17 9 11 9 0 13 16 15 13 9 9 0 9 0 9 0 3 9
8 13 3 3 15 11 0 3 0
5 0 9 9 9 13
2 9 13
29 16 13 0 9 3 13 11 1 9 15 3 13 11 16 9 9 13 1 9 13 9 1 12 11 15 9 9 13 13
6 1 0 9 3 12 13
3 13 9 13
4 11 9 3 13
5 15 3 13 15 13
3 13 9 0
8 7 3 3 0 15 3 13 13
11 11 9 13 0 0 0 0 15 9 9 9
33 0 0 12 9 3 0 16 0 16 9 0 16 0 16 8 7 9 3 8 16 11 1 0 9 1 15 1 15 9 13 13 13 13
9 3 0 1 9 15 1 15 0 13
14 3 7 15 3 9 11 13 13 3 9 0 9 7 9
9 7 13 15 0 1 9 1 11 15
8 3 16 1 0 13 8 9 13
5 15 9 13 15 13
17 11 9 15 0 9 0 9 13 3 0 13 16 16 13 13 0 9
5 1 11 1 9 13
4 13 9 3 13
2 13 9
15 15 15 13 3 13 15 9 0 9 13 13 15 3 3 0
1 3
13 3 3 13 16 3 15 0 9 3 15 15 9 13
38 3 16 7 9 0 3 13 7 1 0 8 7 13 7 13 7 0 9 7 9 9 0 9 13 8 8 8 13 7 7 13 16 1 15 7 13 7 13
14 0 1 9 0 1 15 1 0 9 13 15 0 11 13
16 15 15 13 0 13 15 1 15 9 13 7 3 15 1 15 9
12 3 3 11 13 13 15 15 1 15 13 13 9
5 3 13 13 15 13
1 3
25 13 1 15 15 13 1 9 15 3 1 9 15 13 13 7 3 13 13 3 15 3 3 13 13 13
17 3 16 15 3 13 13 1 9 0 0 3 15 1 0 9 13 13
23 16 3 0 1 9 13 1 15 7 15 9 1 9 13 9 0 15 15 9 7 15 9 13
11 15 9 1 11 1 11 1 0 0 9 13
7 3 13 13 9 9 9 9
5 3 3 15 9 13
12 15 3 0 9 9 15 3 3 9 9 0 13
67 3 3 3 11 13 16 9 1 9 11 9 9 13 1 15 15 15 1 0 9 13 3 9 9 1 15 3 13 15 13 7 16 3 13 16 7 15 7 9 13 15 0 9 13 13 13 9 13 9 9 3 7 13 15 1 9 3 15 13 3 0 7 0 16 3 13 13
53 15 3 16 13 13 13 11 9 15 16 13 13 16 11 0 9 13 15 1 9 9 13 3 13 0 3 13 0 1 9 13 7 9 3 0 9 13 7 13 9 13 9 13 1 9 16 0 0 9 13 13 3 13
30 3 16 9 13 13 9 0 16 9 3 9 0 9 0 13 9 3 0 9 0 15 13 16 3 9 13 3 13 0 13
9 3 3 3 0 1 9 0 9 13
12 0 9 0 9 9 3 3 0 3 3 13 9
23 0 3 0 13 15 9 13 0 3 13 15 0 1 15 0 7 13 13 7 9 9 3 13
15 3 16 15 9 1 9 0 9 13 0 13 9 15 9 9
3 15 13 9
7 13 15 13 11 15 13 3
10 15 13 15 0 9 7 3 3 13 13
33 15 15 9 3 0 13 13 3 7 0 16 13 15 9 11 9 13 13 7 16 9 11 11 16 15 3 9 13 13 15 9 13 13
6 3 0 13 15 9 0
19 3 9 9 16 15 3 1 15 3 9 9 13 13 9 7 3 9 15 13
14 1 15 3 0 9 3 13 15 1 13 9 13 9 13
10 13 0 9 15 3 13 13 3 9 13
6 12 0 9 9 3 13
4 13 9 1 9
4 3 3 7 13
3 13 9 9
4 13 9 15 13
9 8 8 8 8 8 8 8 8 8
17 13 11 1 0 0 0 9 15 1 15 9 1 15 0 1 15 13
3 13 1 15
1 13
1 13
1 13
23 3 0 9 0 0 9 9 12 9 3 0 3 13 16 0 13 9 3 13 13 3 13 15
8 12 13 15 9 3 3 9 13
12 15 11 16 13 15 15 15 13 9 1 15 13
9 13 3 3 13 9 9 7 9 9
10 13 3 15 3 13 9 9 7 15 15
81 9 0 9 0 15 15 15 9 15 0 13 13 15 0 15 9 7 9 9 15 13 7 13 13 16 15 15 9 13 13 13 13 1 9 12 0 9 16 9 13 12 9 9 0 0 7 0 9 13 9 7 9 15 13 7 15 15 3 3 9 0 3 9 13 13 13 15 11 7 11 7 11 7 0 0 9 9 13 3 13 13
23 7 3 16 15 1 9 0 13 3 3 16 13 0 0 13 9 0 9 0 13 9 1 9
36 3 3 3 13 16 9 16 9 16 9 9 16 9 9 13 13 16 3 9 9 7 9 9 1 0 15 13 15 9 15 0 15 13 9 9 15
15 13 3 13 7 0 9 15 15 0 7 9 0 9 8 13
9 11 9 15 1 9 13 3 13 13
9 9 1 0 15 9 13 7 13 13
14 11 0 13 1 9 3 9 0 0 9 3 9 0 9
5 1 15 13 0 13
20 3 0 3 13 13 0 3 7 9 3 7 9 13 0 9 9 15 8 15 13
32 3 3 3 1 9 13 13 15 9 0 13 1 0 9 0 7 0 9 13 1 15 13 3 16 12 9 13 9 0 13 16 13
21 9 13 0 9 15 15 3 7 13 3 7 13 13 16 7 13 0 7 13 0 13
2 13 11
5 3 9 0 13 9
3 13 15 9
7 13 0 1 9 0 0 9
4 9 13 0 9
4 9 3 13 13
10 15 13 9 13 0 7 15 13 13 13
9 1 12 9 0 9 0 0 13 13
3 13 1 9
3 13 0 9
6 13 15 15 1 11 13
5 13 7 3 15 0
8 0 13 13 3 1 9 13 13
7 15 13 9 0 1 9 0
8 13 13 9 15 15 11 9 13
3 13 3 0
9 9 13 13 16 11 15 9 15 13
6 0 3 11 9 9 13
3 9 13 13
5 13 13 13 9 13
5 13 13 15 3 13
6 15 3 13 12 9 13
8 12 16 9 3 13 15 15 13
6 0 9 13 13 7 13
11 1 9 9 7 9 3 0 13 3 3 13
11 3 3 0 15 3 13 13 15 9 3 13
24 13 13 9 9 1 9 7 3 0 3 16 15 0 9 0 9 9 0 0 13 13 1 9 13
43 13 0 16 0 0 9 9 0 7 0 9 15 1 0 11 3 13 13 7 6 0 7 0 9 13 1 15 13 3 3 16 15 0 9 9 0 9 0 1 9 11 11 13
12 3 7 9 7 9 0 8 1 15 0 9 13
4 3 13 9 9
35 1 15 15 0 13 15 11 11 9 7 1 15 3 7 9 3 7 9 13 7 15 11 15 9 13 13 13 1 15 3 9 0 9 13 13
4 15 15 3 13
6 3 9 1 3 13 13
25 0 13 1 9 0 16 15 9 1 9 13 16 3 13 3 13 16 13 16 3 13 0 9 3 13
8 13 0 9 11 11 3 3 13
7 13 3 13 13 7 3 13
3 7 6 15
17 13 3 9 0 15 15 11 3 13 13 16 0 13 13 9 9 13
24 15 1 15 13 15 1 11 13 3 13 3 13 16 13 7 13 16 15 1 0 9 3 3 13
16 7 3 3 13 13 9 15 3 16 15 3 1 9 3 13 13
13 7 13 16 11 16 0 9 13 3 1 0 9 13
10 11 15 9 9 13 0 7 9 11 13
18 1 15 3 3 3 13 16 3 13 0 15 13 3 7 3 13 15 13
3 3 15 13
9 11 16 15 1 15 15 9 13 13
6 1 15 15 15 3 13
12 15 16 12 1 9 13 13 0 1 15 9 13
5 7 0 3 0 13
5 13 15 13 1 11
7 15 15 15 1 15 9 13
3 15 13 13
25 0 15 9 9 7 9 9 7 9 11 9 15 13 13 1 9 15 1 15 1 15 9 0 9 13
30 15 15 13 16 13 3 3 7 3 3 1 9 9 3 7 3 13 15 13 9 3 9 15 13 3 7 3 13 3 13
21 7 3 0 15 0 13 16 3 13 16 15 0 7 11 7 1 0 9 3 13 13
24 15 16 13 13 7 15 13 13 16 15 13 1 15 3 3 9 7 9 7 9 0 9 7 15
29 3 15 13 1 11 9 15 9 15 9 3 0 9 7 1 13 7 1 13 9 15 13 15 1 15 15 15 13 13
11 7 0 9 9 3 13 3 13 13 3 13
9 13 3 16 16 13 15 3 13 15
18 3 3 13 16 15 1 0 9 13 13 0 3 15 13 15 3 13 13
41 1 0 9 15 1 15 11 13 7 1 9 15 1 0 7 11 1 9 15 7 1 9 13 13 3 0 9 13 13 7 15 1 15 13 13 9 15 9 0 13 9
48 3 16 3 13 7 0 9 13 0 3 9 7 0 0 7 13 0 9 16 3 13 9 7 9 3 9 7 0 15 9 13 15 1 15 15 7 9 7 9 7 9 13 13 3 0 3 13 13
6 15 15 16 13 15 13
22 3 1 15 15 15 3 13 3 13 15 13 15 15 7 15 3 13 7 1 15 3 13
25 0 9 9 15 3 13 0 1 15 13 15 9 7 0 7 0 9 7 15 9 7 15 0 9 13
32 3 7 15 1 15 7 15 15 13 3 13 1 9 13 9 16 15 9 15 1 9 9 15 3 15 3 13 9 1 0 9 13
14 0 3 9 9 9 9 3 7 15 15 3 7 15 13
15 13 3 13 3 7 13 1 15 0 9 7 9 7 9 15
13 13 15 3 7 9 15 9 15 0 7 9 9 0
24 3 15 3 15 0 3 3 9 15 15 13 7 3 9 9 15 15 0 15 1 13 13 3 13
2 15 13
47 1 0 3 9 15 1 9 15 0 13 3 13 7 1 0 9 15 3 1 9 13 3 16 9 13 9 13 7 1 0 0 9 1 15 15 3 3 3 3 1 9 9 15 9 7 15 13
29 3 3 9 15 3 9 3 9 3 9 3 0 9 3 0 3 0 3 0 13 3 15 0 7 0 9 7 9 13
22 3 3 0 13 0 1 0 9 9 15 1 15 15 7 9 15 15 13 7 13 13 13
16 3 7 0 15 13 13 7 0 15 15 13 3 13 15 9 13
10 15 3 1 9 0 0 0 0 7 13
11 13 3 15 13 15 9 3 1 9 13 13
19 15 3 0 3 3 13 13 1 9 9 13 16 1 15 15 1 13 13 13
39 15 1 9 13 16 15 9 3 13 13 7 0 0 9 13 3 3 7 3 13 13 9 3 15 13 13 0 1 9 7 1 9 3 0 3 0 7 0 13
6 6 15 9 9 3 13
8 15 15 3 3 13 7 3 13
7 15 0 1 9 7 3 0
9 3 16 0 13 0 13 11 15 13
7 0 9 0 9 7 9 9
11 0 13 9 16 16 15 13 3 13 1 9
30 0 3 9 13 13 3 1 15 13 7 16 0 9 7 0 13 0 7 1 15 1 9 9 7 9 13 13 3 7 3
10 3 7 3 9 13 13 7 9 9 13
22 12 3 3 13 11 9 13 7 13 13 1 15 1 9 9 13 3 13 9 0 15 11
15 3 15 13 9 9 7 15 13 3 13 0 1 15 13 0
7 15 15 9 3 13 3 13
4 9 0 13 3
3 13 11 3
3 13 15 13
16 13 15 13 13 7 13 3 1 15 1 15 9 13 9 0 0
8 11 13 9 13 1 9 3 13
5 12 3 0 13 13
18 11 1 15 13 1 11 13 7 11 1 0 15 13 1 11 11 13 13
2 15 13
5 15 15 13 1 15
1 15
6 0 13 7 1 15 9
5 13 13 13 16 13
11 3 0 3 13 15 3 13 16 3 3 13
1 3
6 13 3 9 8 7 0
37 15 3 15 3 9 7 9 9 15 9 7 9 13 15 15 15 7 1 0 9 9 7 1 0 15 0 7 15 15 9 7 9 9 13 13 3 13
18 3 13 1 15 13 16 3 9 13 3 1 9 7 9 7 0 11 13
12 3 0 0 15 0 7 9 13 1 15 9 0
4 9 0 3 13
30 3 16 3 13 9 13 9 0 16 1 9 13 9 9 13 13 1 0 9 15 13 15 1 7 13 3 7 13 3 13
3 3 15 13
4 15 3 3 13
8 0 13 3 15 15 13 13 7
18 7 0 3 9 9 15 7 9 13 3 7 15 0 9 7 0 9 13
21 7 0 13 3 15 13 3 13 0 7 3 13 7 13 7 15 0 9 7 9 13
9 1 9 0 3 16 9 13 0 3
21 3 16 15 3 15 1 15 9 13 13 13 3 13 3 13 9 0 3 13 3 13
46 3 1 9 15 0 3 13 9 13 1 9 9 0 1 15 15 13 3 15 13 9 13 9 7 13 9 0 13 7 15 13 9 9 7 9 15 3 9 13 15 7 9 13 7 13 9
5 13 15 13 3 13
14 9 13 13 0 15 15 15 1 15 9 13 1 9 13
3 15 0 9
2 13 9
3 13 9 0
12 3 0 9 12 9 9 0 1 15 12 13 13
9 3 7 9 9 13 7 9 9 13
11 15 9 0 9 13 16 0 9 11 3 13
8 3 11 11 9 11 15 9 13
6 11 3 15 13 9 13
17 16 0 9 0 9 3 13 0 15 11 3 11 3 11 0 3 13
3 3 13 13
12 9 3 15 13 7 11 9 15 9 15 13 13
20 15 1 9 11 11 13 0 7 13 16 0 9 1 9 0 9 1 9 11 13
20 11 13 9 0 7 15 13 7 13 9 15 16 13 9 9 13 0 0 1 11
12 11 3 9 6 9 0 3 0 7 1 9 9
12 3 0 15 11 3 13 9 1 3 13 3 13
13 0 3 13 13 1 11 3 0 0 3 15 13 0
9 7 3 8 8 8 8 15 13 13
5 11 9 15 1 9
3 0 3 13
16 12 13 15 13 9 3 7 9 3 3 15 13 9 7 9 11
19 15 0 9 15 13 0 15 0 3 9 13 3 7 15 1 9 9 13 13
12 3 15 13 0 1 9 15 13 16 9 13 13
6 3 3 9 13 13 13
44 3 13 15 9 13 7 16 1 0 15 13 0 3 1 15 3 13 13 13 15 3 7 16 13 0 13 3 15 13 3 13 16 9 15 0 13 16 3 3 1 0 9 13 13
10 3 16 0 13 13 13 7 13 9 15
7 3 13 16 15 3 3 13
6 3 11 11 11 11 9
32 3 3 16 15 0 13 9 15 13 15 3 3 16 3 0 9 13 13 3 15 13 3 15 13 7 1 13 3 13 0 3 15
21 7 1 0 7 0 9 15 13 16 15 1 15 13 9 1 15 1 9 7 9 13
15 7 3 15 3 0 13 9 13 9 15 13 1 9 0 13
18 3 16 15 9 15 0 13 13 3 1 15 15 15 13 15 3 13 13
11 7 1 9 0 3 3 3 0 9 13 9
20 3 9 9 15 9 3 0 13 7 9 1 9 13 1 9 9 7 1 9 13
24 7 0 9 0 3 13 13 16 16 1 0 15 0 9 13 12 9 9 0 13 15 1 9 13
15 0 0 1 15 11 13 16 15 12 3 9 9 0 13 13
12 15 3 15 15 1 15 8 13 16 0 3 13
6 0 3 9 3 15 13
10 0 9 1 11 9 9 3 13 9 11
6 15 15 0 13 1 9
15 1 0 15 9 0 9 9 15 0 13 15 1 9 9 13
11 13 9 0 15 11 11 11 11 9 0 13
14 9 7 9 15 9 11 13 3 7 13 1 15 9 13
17 12 9 3 13 16 9 0 0 9 13 15 1 0 9 1 9 13
12 0 0 9 0 9 13 13 11 0 15 9 13
7 11 3 1 9 13 9 13
10 15 3 0 1 9 9 13 15 9 9
10 9 3 7 11 3 15 3 13 13 9
13 15 13 3 7 9 9 13 7 9 9 13 13 13
7 7 0 0 9 13 9 13
34 0 13 1 9 0 16 3 0 1 9 0 13 13 0 15 9 9 9 15 3 9 0 7 13 3 3 1 11 11 1 9 13 13 13
3 0 3 13
7 0 13 3 13 1 9 0
82 15 3 3 3 9 0 0 13 9 7 0 9 0 15 7 0 9 13 13 3 13 0 9 9 1 9 0 13 7 0 13 7 13 9 13 7 16 3 11 9 9 9 7 9 13 3 13 15 0 3 1 9 13 16 1 15 0 3 13 3 3 0 9 0 0 13 9 15 3 3 15 13 13 15 0 15 9 7 0 9 13 13
33 3 3 15 15 3 3 1 9 15 13 11 13 1 0 9 16 1 9 3 3 7 3 0 7 9 0 15 9 9 7 9 9 13
41 15 3 3 13 15 3 7 3 0 9 7 3 13 0 16 9 7 3 0 16 9 13 3 9 0 16 13 15 0 15 9 13 15 15 1 11 1 9 0 9 13
23 1 0 15 15 0 9 13 16 15 15 1 15 9 0 7 1 9 0 0 0 9 13 13
12 7 15 3 9 7 9 3 15 9 3 13 13
5 15 13 3 3 13
12 13 3 0 9 0 0 0 9 15 15 9 13
25 3 15 15 13 1 13 13 1 15 9 9 13 13 15 9 3 13 0 3 1 9 0 1 9 13
19 7 3 13 13 1 11 11 9 15 1 0 9 13 7 13 0 9 3 13
9 3 9 15 9 13 3 3 13 13
14 15 16 15 9 3 1 9 9 15 13 13 15 13 0
39 1 15 16 15 13 15 9 0 3 0 0 7 13 3 13 15 15 16 13 11 11 1 15 12 13 15 15 3 0 13 0 9 13 3 9 15 7 8 13
12 1 15 16 15 13 0 9 15 0 13 7 0
12 0 9 13 16 15 9 1 15 0 9 15 13
4 3 15 13 13
3 8 3 8
10 16 13 3 1 9 15 15 3 13 13
9 3 3 8 13 0 7 8 15 13
10 3 0 15 1 0 9 7 9 13 13
5 15 3 15 13 3
26 11 0 15 13 9 3 15 0 9 7 3 0 7 0 15 13 13 7 0 15 13 15 15 15 9 13
19 16 1 0 15 11 13 3 11 15 0 15 1 15 9 13 15 15 3 13
6 0 3 9 9 0 13
10 7 3 15 13 13 9 1 15 15 13
32 3 15 1 0 9 15 15 3 1 15 7 15 7 3 13 13 0 13 3 13 15 7 3 7 9 0 7 9 0 7 9 13
12 3 13 13 3 16 15 9 13 3 1 15 13
22 15 1 15 1 9 0 13 13 15 3 7 3 7 3 7 1 15 9 9 15 3 13
34 3 3 7 1 9 15 15 9 13 13 3 7 1 15 9 1 0 9 13 7 15 1 15 13 15 13 0 15 0 15 3 13 7 0
45 3 3 13 9 15 3 1 9 15 9 3 0 7 6 9 0 3 3 0 3 15 9 0 9 1 15 13 16 9 0 9 9 9 13 9 13 7 1 9 9 1 15 9 9 13
21 7 3 1 15 3 13 13 15 3 16 15 0 13 0 7 16 0 15 13 0 13
17 0 3 1 15 13 7 13 16 3 13 16 15 15 13 3 13 13
30 15 0 9 0 15 13 7 0 15 15 13 13 3 3 3 3 13 7 3 16 15 1 0 13 3 1 15 0 9 13
11 3 3 13 11 3 13 8 8 8 8 8
4 8 8 8 8
16 15 3 3 13 9 15 7 13 1 15 3 7 1 9 15 13
27 1 9 3 15 15 9 13 7 16 3 0 13 7 16 9 15 3 0 7 16 1 9 15 13 3 15 13
13 1 9 3 1 15 13 3 3 0 9 13 1 9
6 3 16 15 13 0 13
6 15 9 16 15 13 13
20 13 9 9 9 3 13 16 3 7 13 15 13 7 0 3 9 3 9 9 13
5 11 15 13 0 9
11 12 13 16 9 13 1 11 3 0 9 13
3 13 13 13
3 0 13 3
2 0 0
10 1 15 9 13 1 15 3 13 9 15
10 13 15 0 15 13 0 3 0 0 13
6 15 16 13 13 1 15
3 7 15 13
22 3 16 1 9 15 13 11 11 11 9 0 9 7 15 15 9 0 15 11 11 13 13
17 16 15 1 9 0 13 13 11 9 15 13 3 13 15 13 16 13
25 3 16 15 13 16 15 1 15 13 13 13 1 9 9 9 9 3 7 9 15 16 9 3 15 13
17 3 7 0 0 9 15 13 7 0 15 13 0 13 15 3 9 13
12 15 15 9 1 15 7 9 9 15 3 13 13
20 1 15 13 13 15 3 3 1 0 9 3 3 13 9 11 11 1 15 13 13
12 3 16 15 15 3 13 13 15 1 15 13 13
31 3 15 0 13 3 3 0 15 7 0 13 13 7 3 13 13 0 0 16 9 13 7 3 9 3 3 13 16 15 13 13
18 15 3 9 0 11 9 7 15 15 9 9 7 3 15 3 0 9 13
10 15 15 11 3 15 15 9 13 3 13
7 3 3 3 13 1 11 13
13 15 15 15 3 13 13 13 16 15 3 7 3 13
2 15 13
3 13 0 9
14 3 3 15 13 16 13 15 15 13 3 13 15 9 13
15 15 16 15 13 9 13 16 7 11 13 7 1 0 9 11
8 13 3 13 15 15 9 9 13
21 9 3 7 15 13 7 0 3 13 16 3 15 15 15 13 9 9 13 15 3 13
41 13 3 15 0 16 1 0 9 15 0 13 13 9 0 15 11 7 16 15 1 0 0 0 13 9 13 16 8 8 7 8 13 13 16 15 3 13 9 15 0 13
6 15 12 13 1 9 3
3 0 1 11
4 0 1 13 9
6 0 16 9 1 9 13
4 0 16 11 13
9 0 15 13 1 9 3 3 11 13
7 0 1 9 15 9 9 13
4 0 1 9 3
25 0 0 8 13 16 13 7 16 15 3 9 3 9 15 13 0 1 9 13 7 15 13 7 15 13
6 15 3 15 15 3 13
32 3 13 15 13 3 15 13 7 3 13 15 9 13 13 3 7 13 16 3 3 16 9 13 7 3 16 13 13 15 3 13 3
9 3 3 13 15 9 9 3 13 13
9 3 13 3 3 16 13 1 0 9
8 3 15 15 13 7 15 15 13
18 7 3 3 9 13 7 16 3 3 9 11 13 13 3 15 15 3 13
2 15 13
9 13 9 8 7 3 3 13 9 0
51 15 1 9 16 1 9 13 13 9 7 9 15 13 15 11 9 9 13 16 1 11 9 15 13 13 3 7 0 9 13 13 15 13 16 9 3 15 13 13 0 9 0 13 3 0 15 15 9 9 13 13
33 3 16 15 0 0 9 13 1 9 3 7 15 1 15 13 13 7 3 15 13 13 1 15 7 15 1 9 13 15 15 0 13 13
5 1 11 0 9 11
5 3 12 9 11 11
2 3 13
4 3 13 13 3
7 3 3 3 16 13 3 13
2 15 13
8 3 3 3 1 15 13 7 13
14 3 3 16 9 13 13 1 15 3 13 9 9 9 13
1 13
18 3 15 13 0 9 13 7 9 15 0 13 0 9 12 15 0 9 13
4 13 3 0 13
4 3 0 13 9
1 13
6 7 15 0 13 3 0
18 15 1 9 9 13 3 7 3 1 11 7 3 1 11 16 15 3 13
9 16 1 0 9 13 3 3 13 13
42 16 15 15 9 0 9 1 11 9 13 13 3 13 15 15 9 9 1 0 13 13 7 3 9 13 13 16 16 1 15 13 15 3 9 0 1 9 0 9 13 13 3
16 15 1 15 9 1 15 15 0 13 3 13 3 3 1 15 13
10 15 3 3 13 15 13 9 0 13 9
7 0 13 0 15 3 13 13
4 9 0 3 13
1 15
27 3 3 16 15 15 13 16 15 3 13 0 13 3 3 3 13 13 9 15 13 0 9 9 0 3 15 13
50 3 3 16 9 0 15 15 1 9 0 15 9 7 9 13 9 13 15 3 9 9 15 9 13 13 16 9 0 1 9 13 15 1 9 13 15 3 13 3 15 3 13 13 16 13 16 13 13 15 13
13 7 3 0 0 9 13 7 0 9 13 3 9 0
12 13 3 3 1 11 8 3 3 1 11 9 9
12 15 0 3 1 9 13 15 1 9 13 9 13
3 13 0 11
2 13 9
5 9 9 9 3 15
4 15 0 9 13
4 13 7 13 11
28 3 3 9 1 9 13 3 3 9 13 13 15 15 15 15 9 3 7 0 9 15 1 15 13 9 0 13 13
2 15 3
5 0 13 9 13 13
6 15 13 16 3 3 13
6 3 9 7 3 9 13
6 7 3 15 13 8 8
6 13 11 3 7 3 3
11 13 3 16 11 13 9 3 3 11 9 13
5 15 16 13 3 13
7 3 3 13 3 9 0 9
12 11 15 13 13 1 15 16 11 13 15 13 9
10 16 9 15 13 11 7 0 9 13 11
1 15
8 0 9 3 1 0 0 9 13
5 3 1 9 0 13
7 11 15 15 13 7 13 15
21 0 7 0 3 15 13 3 16 15 0 0 9 9 0 9 3 0 7 0 0 13
5 1 11 13 13 9
17 11 15 1 9 1 9 13 7 3 15 13 1 9 15 13 1 15
10 3 15 11 13 13 15 9 0 11 13
12 15 1 15 9 15 1 15 1 9 15 13 13
14 11 3 3 1 15 13 15 9 15 9 15 13 15 13
6 0 15 15 13 13 0
10 7 3 0 3 3 3 0 16 13 13
5 15 13 0 9 13
4 1 11 13 9
5 1 15 15 13 13
15 3 7 3 0 15 9 0 13 13 3 7 15 1 9 13
5 7 13 3 13 3
4 15 15 8 13
11 6 0 9 7 3 3 0 13 3 1 11
7 8 7 8 13 15 11 13
4 15 0 9 13
11 8 16 9 13 15 3 13 3 12 9 13
4 15 15 9 13
6 1 15 3 13 3 13
5 1 9 0 3 13
3 1 9 13
2 9 13
15 3 3 1 15 13 11 13 1 9 15 9 15 3 13 13
23 13 3 16 15 13 1 11 9 15 13 13 1 15 7 16 3 3 13 13 1 15 3 3
3 13 3 13
3 13 16 13
5 11 13 13 11 13
13 15 9 11 9 13 13 7 11 13 3 13 0 13
9 3 15 9 15 7 9 0 3 13
9 9 9 16 13 13 15 8 8 13
16 3 16 15 0 3 13 11 13 9 8 0 9 3 3 13 0
16 3 8 8 8 8 8 8 8 8 8 8 8 8 8 8 8
3 13 3 0
17 0 16 13 3 13 0 3 16 15 13 0 9 16 1 9 13 13
5 13 9 3 0 9
40 3 7 3 13 13 9 0 1 15 13 15 9 7 0 9 7 13 15 13 3 0 3 13 1 11 7 11 7 3 13 15 1 15 13 11 3 13 16 3 13
10 3 13 1 15 11 0 13 11 11 9
23 3 13 0 9 15 0 1 11 16 13 3 1 11 9 1 9 1 9 9 1 9 9 9
11 7 15 8 15 0 13 15 13 1 9 0
23 3 9 15 0 1 9 9 15 7 3 9 9 9 7 13 0 13 7 13 9 9 7 0
4 15 3 11 13
3 9 13 13
4 7 11 11 13
2 9 13
22 13 15 0 16 11 9 1 15 13 1 15 3 15 15 1 15 13 13 0 9 3 13
16 3 16 9 9 13 13 13 15 13 16 1 11 15 9 13 13
21 16 1 15 15 13 3 13 15 3 13 15 15 3 13 13 13 16 9 11 13 13
11 3 0 13 16 13 3 3 13 3 7 13
6 11 3 3 13 1 11
2 13 9
3 7 3 13
29 0 3 15 13 1 0 9 9 0 3 7 11 15 3 3 13 1 9 13 7 0 9 0 9 15 9 13 13 13
32 3 3 1 11 15 13 9 0 3 3 3 13 7 0 3 7 15 3 13 1 9 11 13 3 7 13 16 1 15 0 3 13
4 7 15 0 13
15 15 15 13 1 9 0 7 3 15 9 13 13 13 16 13
4 3 3 13 0
8 13 3 15 3 1 9 0 13
3 11 9 13
2 15 13
10 1 9 0 15 13 16 11 0 13 13
10 15 1 3 7 1 0 13 7 1 0
12 1 9 13 11 16 13 16 0 13 15 15 13
5 15 13 3 13 11
29 0 9 3 0 9 0 15 0 13 12 9 9 9 0 7 3 3 16 15 0 13 3 11 7 9 13 1 9 9
23 13 3 7 3 13 11 0 7 11 13 7 3 1 0 9 9 15 13 7 1 15 9 13
11 7 0 9 7 0 13 8 8 8 8 8
9 15 3 15 9 16 15 0 13 13
8 3 15 15 9 1 9 13 13
9 15 3 9 1 15 1 9 12 13
5 7 13 13 7 13
10 16 3 13 13 15 15 9 7 3 13
8 3 6 13 1 3 13 0 9
11 3 16 15 8 15 1 3 13 3 3 13
50 1 0 9 13 15 9 15 11 13 15 9 15 13 13 7 15 9 13 3 3 9 9 11 7 11 7 3 15 13 1 11 11 11 7 3 15 0 9 7 3 15 0 3 7 16 11 13 15 9 13
8 15 3 12 15 1 0 13 13
3 13 9 15
14 7 15 15 0 15 13 13 7 0 9 7 15 9 8
18 3 3 16 15 13 13 0 13 13 3 13 0 1 15 9 9 13 13
60 15 3 1 11 1 15 13 3 7 3 15 1 15 9 13 7 15 1 11 11 13 7 15 3 13 8 8 13 7 15 9 11 15 13 13 13 1 15 13 16 0 15 13 15 1 9 13 13 9 7 3 13 1 0 9 1 15 1 15 13
5 3 3 13 15 9
16 16 15 0 9 13 13 16 9 13 0 9 15 3 0 9 13
11 3 3 13 13 9 16 1 15 13 3 13
13 3 7 9 15 13 15 13 11 0 9 7 9 13
8 3 1 9 13 9 3 13 0
7 3 8 15 13 0 9 13
5 15 13 16 11 13
47 7 6 13 9 0 1 13 7 8 3 7 3 13 8 3 13 7 15 9 13 15 15 3 0 9 13 13 15 3 13 3 3 11 13 7 0 9 15 13 3 3 15 13 9 3 11 13
6 15 3 0 11 9 13
10 7 15 13 0 13 0 9 0 9 9
32 13 9 3 1 11 3 0 13 15 11 3 13 3 15 13 1 15 15 15 1 12 9 0 7 0 13 3 15 13 15 13 15
4 3 3 3 8
13 3 8 15 15 12 13 0 9 7 3 0 3 13
20 3 15 3 15 8 3 13 0 7 0 0 15 1 9 7 3 1 15 13 9
11 13 15 13 15 9 13 9 7 9 0 13
7 3 1 9 13 15 13 13
2 15 15
1 3
8 3 15 13 3 13 13 16 13
6 9 3 1 15 12 13
6 15 0 3 13 15 13
7 0 16 13 15 15 3 13
8 3 15 13 16 15 3 13 13
37 1 11 15 1 15 13 3 15 0 13 15 7 3 13 15 9 13 1 15 13 16 13 7 3 13 16 15 13 7 13 7 3 1 9 15 13 13
2 15 3
7 1 9 13 16 11 13 13
6 9 0 9 13 3 13
2 15 13
7 13 15 1 13 0 15 9
19 15 16 0 13 7 16 3 13 9 15 13 7 9 7 9 9 0 9 0
3 15 13 13
13 0 0 1 13 9 11 3 13 0 7 9 11 13
12 0 0 9 9 13 15 15 9 1 0 9 13
8 0 9 13 9 0 1 0 9
7 15 15 15 9 13 1 11
7 3 3 11 9 15 13 13
7 11 7 0 0 9 0 13
2 13 3
11 13 15 0 1 0 9 9 1 15 3 13
17 7 0 15 13 13 13 15 13 3 3 3 1 0 12 9 13 15
9 16 13 3 15 0 13 0 3 13
8 3 3 13 15 13 3 16 13
18 3 3 16 13 13 1 9 3 13 7 13 9 13 0 9 1 9 13
14 13 3 13 15 9 11 8 8 8 8 8 8 8 8
6 1 9 15 9 13 13
4 11 15 9 13
7 1 8 16 15 13 3 13
16 9 16 1 15 3 13 1 9 3 13 6 15 9 9 13 11
1 13
3 13 15 9
1 13
2 15 13
1 13
4 15 3 1 11
2 3 13
15 15 3 1 15 1 0 9 9 0 15 9 0 7 0 13
17 3 16 15 1 0 9 15 3 13 13 9 0 13 3 3 16 13
7 16 15 1 9 13 15 0
8 7 13 11 9 13 1 15 13
9 3 15 9 1 11 1 15 9 13
8 15 3 0 1 9 9 13 0
10 3 13 13 13 9 3 7 13 0 13
3 13 15 13
10 15 15 13 9 16 13 15 11 13 13
4 15 15 13 0
10 7 13 9 15 16 13 3 15 13 13
5 1 0 13 13 9
19 3 16 13 13 15 13 0 9 9 0 0 3 1 0 13 16 9 13 3
4 15 11 13 13
4 3 13 1 11
12 15 7 1 0 7 11 7 1 0 13 16 13
8 9 0 13 15 7 13 15 0
38 3 16 15 13 11 9 9 15 11 13 0 13 3 16 15 13 0 1 11 9 3 15 1 15 13 3 0 15 13 7 13 0 13 15 1 15 13 13
26 0 3 15 3 13 13 15 0 8 16 1 11 13 1 15 13 13 3 13 13 15 0 13 15 13 0
28 16 3 15 1 15 13 13 15 3 13 1 9 13 16 13 0 15 0 9 1 9 3 0 15 0 9 9 13
4 15 13 0 8
28 3 3 9 13 16 13 9 0 1 0 9 1 9 3 3 1 0 9 7 3 1 0 3 9 11 13 15 13
10 16 3 1 15 13 13 0 1 15 13
19 3 15 13 7 0 9 3 13 9 0 1 9 0 13 13 3 3 3 13
37 0 9 11 7 3 9 0 15 9 15 0 9 15 0 7 0 15 0 7 0 13 15 15 9 9 0 13 15 9 15 9 9 15 0 9 0 13
9 13 3 3 9 13 7 3 13 13
19 15 15 13 3 7 9 3 7 1 11 13 16 0 9 13 15 0 9 13
22 3 16 13 0 9 9 16 15 3 1 9 7 1 12 9 0 13 13 15 3 13 13
9 3 0 13 13 15 13 9 9 9
17 13 0 9 0 3 3 15 15 15 13 7 3 0 0 15 13 11
3 9 0 13
4 7 0 3 3
4 3 13 15 13
7 11 15 1 11 13 13 3
6 11 13 3 13 1 0
15 7 16 1 0 13 3 13 3 1 3 13 13 3 15 0
4 13 13 15 9
5 9 11 13 3 13
18 13 3 8 16 13 13 15 9 9 3 8 3 3 3 7 3 3 13
9 3 13 16 13 15 9 15 13 13
5 1 11 9 9 0
7 13 15 3 3 1 12 9
2 13 15
20 9 3 15 13 11 16 13 15 9 3 3 13 11 15 13 3 15 15 13 11
24 3 9 15 3 3 15 11 7 3 15 1 9 0 3 7 3 15 13 0 3 15 13 13 13
12 3 3 16 15 1 13 9 13 13 13 15 13
37 3 16 3 15 0 13 3 0 9 15 1 15 3 13 13 13 0 15 9 0 15 3 3 9 7 3 9 15 7 9 15 11 13 13 13 16 13
11 3 16 1 0 9 3 13 11 15 3 13
6 3 11 15 15 15 13
2 0 3
6 13 0 11 0 13 13
9 0 3 9 13 7 13 15 9 13
6 13 1 15 11 15 13
12 13 9 15 9 11 11 15 13 15 1 9 13
9 6 0 9 15 12 9 15 13 12
4 13 3 3 13
3 7 13 8
7 3 3 9 1 15 1 9
7 0 1 15 15 3 13 0
2 15 13
5 11 13 9 9 13
2 15 13
10 7 0 3 11 7 16 15 13 0 13
1 13
7 3 15 11 11 11 13 9
6 13 9 13 13 1 9
6 3 13 15 13 8 8
34 3 3 13 1 15 9 3 1 0 9 15 13 1 9 0 1 9 11 1 9 8 1 9 11 1 9 13 1 11 1 11 9 7 9
8 15 3 15 9 13 9 0 8
15 13 1 9 8 7 3 3 13 15 0 1 15 8 3 13
3 0 13 13
14 15 16 3 1 15 13 3 13 0 13 3 7 3 0
3 11 3 13
12 0 9 13 7 9 3 3 0 3 0 15 8
22 9 13 9 0 9 3 3 15 13 7 15 13 13 3 13 3 15 15 15 0 3 13
5 11 13 13 15 9
12 13 15 0 9 8 8 8 8 8 8 8 8
23 3 13 0 9 3 0 13 9 0 0 9 13 13 15 15 13 7 1 15 1 0 13 13
15 3 15 15 9 13 13 1 15 13 3 15 3 0 0 13
6 3 6 1 9 3 13
8 3 3 0 9 9 15 13 13
12 16 3 1 0 8 13 8 11 13 15 9 9
3 3 13 9
6 15 1 9 15 9 11
8 15 9 3 1 11 0 9 13
3 13 15 13
11 15 3 13 15 0 3 3 3 15 13 13
13 15 16 9 1 0 13 13 1 0 3 15 3 13
8 3 3 13 13 3 1 13 9
28 3 15 13 3 15 3 13 15 13 3 16 0 15 11 16 15 15 9 13 13 7 16 0 9 8 13 13 13
19 15 3 3 3 13 13 16 0 9 15 3 13 13 8 3 1 0 9 13
9 1 13 16 15 3 13 13 15 13
6 9 13 3 9 9 0
3 7 13 9
5 11 11 0 13 9
3 3 15 13
8 13 3 15 9 9 13 13 15
17 6 9 0 16 15 3 16 15 1 15 13 13 1 15 9 0 13
4 7 3 0 13
8 0 15 13 7 0 9 7 9
10 7 3 3 13 1 15 3 7 13 9
10 3 3 0 1 9 0 3 1 9 15
10 7 3 0 0 15 9 9 9 7 13
13 0 3 13 3 13 15 13 13 15 13 1 9 0
18 11 3 0 9 9 1 9 9 15 13 3 15 9 1 15 9 9 0
5 3 1 11 9 13
1 13
13 13 9 9 16 15 15 16 3 3 15 1 11 13
14 7 0 3 3 0 13 16 16 15 13 0 9 13 13
23 3 3 0 3 13 3 16 7 13 16 7 13 9 0 0 9 15 13 3 15 9 13 13
7 16 0 3 13 6 15 11
1 13
2 13 11
4 0 13 11 13
8 15 15 9 13 16 1 0 13
27 3 16 0 3 13 1 0 3 3 1 0 0 3 3 16 16 15 0 15 13 1 0 15 13 3 1 3
10 11 0 13 9 15 7 9 1 9 0
11 13 3 15 0 9 13 15 15 9 0 13
6 7 3 15 15 9 13
9 15 15 3 7 8 8 8 9 13
16 13 15 7 3 13 3 9 13 0 13 1 15 1 9 0 13
2 15 13
5 13 3 0 3 13
21 3 1 15 15 0 9 13 1 9 15 0 13 13 13 15 15 15 13 0 15 13
6 0 15 0 9 3 13
13 15 9 16 0 0 13 3 3 9 12 12 13 13
8 0 15 9 1 0 13 3 13
10 15 15 13 12 9 9 9 15 13 13
8 11 3 15 3 3 15 13 13
6 15 3 3 3 13 13
12 3 3 0 8 15 9 11 13 9 15 13 13
12 0 9 15 13 13 13 3 3 15 1 15 13
7 1 9 0 13 15 3 13
11 11 1 9 3 13 3 3 15 13 3 13
6 1 9 13 0 9 13
5 3 3 11 15 13
1 15
3 0 3 13
6 13 15 13 13 9 11
31 3 6 15 15 3 3 0 9 3 0 9 0 9 15 13 0 15 15 3 3 9 7 3 9 3 3 9 15 7 9 13
13 3 16 1 0 15 9 13 3 3 15 13 13 9
36 3 3 0 13 16 16 0 9 13 11 9 15 1 11 9 15 16 0 15 8 8 8 3 15 13 0 3 8 8 15 1 15 9 13 13 13
6 13 3 15 11 3 13
14 16 1 11 9 9 13 1 15 3 13 8 8 8 8
3 15 13 13
11 3 3 13 0 9 9 15 16 15 13 13
12 3 3 13 16 15 13 16 9 15 13 7 13
9 0 3 15 13 13 13 1 9 9
9 13 15 1 9 9 9 1 9 13
15 3 3 15 9 13 15 1 15 9 13 7 13 13 3 13
25 13 16 15 0 3 11 1 11 1 0 9 13 13 7 16 15 13 15 13 15 15 1 0 9 13
15 8 8 8 3 15 1 13 1 0 9 13 0 11 7 9
5 3 15 3 3 13
7 0 15 13 3 15 9 13
4 7 15 15 13
8 9 3 13 3 3 1 9 13
17 3 16 15 15 13 16 13 15 13 15 3 0 3 13 15 0 13
12 15 1 11 13 7 9 0 13 16 0 0 13
5 3 3 13 3 13
3 8 8 8
13 15 3 0 0 9 9 15 9 0 15 9 9 13
19 15 16 13 0 3 13 3 0 7 0 9 9 13 16 0 0 13 3 13
2 15 3
7 15 0 0 1 15 13 13
11 3 3 13 16 1 15 9 0 9 15 13
18 3 3 13 0 1 11 3 3 3 13 16 7 9 7 9 9 15 13
23 9 0 3 3 15 8 13 3 3 3 8 15 15 1 9 3 13 3 1 0 0 7 0
16 13 3 15 13 16 11 9 1 9 1 9 12 0 13 3 15
7 0 3 9 3 3 0 13
8 13 3 0 3 16 0 13 13
3 7 0 3
9 15 3 13 15 11 13 1 15 9
9 15 3 3 13 16 15 9 13 13
16 13 3 8 8 8 7 1 15 1 15 3 8 13 3 15 13
9 15 1 15 9 13 8 8 8 13
19 13 3 3 7 3 16 13 13 7 9 7 9 3 0 13 15 3 13 0
15 7 0 9 15 3 13 12 9 15 13 3 7 9 15 13
11 8 13 3 13 0 15 13 15 15 9 13
7 0 13 7 3 13 9 11
13 0 9 0 9 0 0 9 3 9 9 1 0 13
16 0 1 9 3 9 7 9 13 0 16 13 9 9 13 9 13
27 7 16 3 13 8 8 1 0 9 0 9 3 13 13 9 16 15 13 3 3 3 9 3 3 9 0 13
15 0 3 1 9 9 1 9 3 7 1 9 13 0 3 13
20 13 3 0 9 9 1 9 9 16 9 13 3 3 9 13 3 3 1 9 0
4 3 13 13 0
11 11 13 3 13 16 9 9 13 13 16 13
8 7 1 9 0 3 13 0 13
13 15 13 3 13 15 3 3 3 0 9 13 3 3
19 1 11 3 3 13 1 9 0 15 16 13 9 7 3 0 9 9 9 13
16 7 0 7 9 1 9 11 3 13 3 7 1 9 9 15 13
11 0 7 0 13 7 3 13 16 13 16 13
4 3 3 13 15
3 3 13 13
2 13 13
3 7 15 13
3 15 0 13
13 1 11 13 7 0 15 9 13 3 7 3 3 13
6 15 13 15 7 13 13
8 3 7 15 9 3 7 9 13
20 0 15 13 7 1 9 0 0 9 7 1 0 9 15 15 0 13 7 12 13
8 7 15 15 13 0 3 11 13
14 3 7 15 13 13 3 7 3 13 1 9 15 13 9
10 15 3 3 13 13 3 15 15 3 13
5 3 13 7 3 3
4 0 1 0 9
10 9 11 9 7 15 15 13 3 15 13
15 3 7 13 15 13 15 0 1 9 7 13 15 1 9 13
4 9 8 3 8
2 15 0
3 3 3 13
4 15 3 15 13
8 15 3 8 7 3 8 8 8
29 13 15 3 13 3 0 3 0 3 3 15 9 9 9 13 3 0 9 15 3 13 3 6 3 13 3 3 3 13
8 0 0 3 3 0 9 13 13
18 11 1 9 13 3 7 3 13 7 3 13 16 0 9 15 13 13 9
7 16 9 3 13 15 13 13
20 15 3 3 7 13 1 0 9 1 0 9 3 7 13 16 15 13 15 3 13
2 13 9
8 9 9 3 9 7 9 13 13
8 3 9 3 9 3 9 9 13
10 9 0 11 9 1 15 11 3 13 13
5 15 9 15 13 0
4 3 13 13 13
7 0 9 9 13 3 7 0
16 3 7 0 9 13 0 9 16 1 9 1 9 11 13 13 13
8 16 3 7 9 3 7 9 13
9 7 0 0 1 9 7 9 13 13
9 11 16 13 13 9 11 9 13 13
11 0 3 13 13 16 0 9 0 11 13 13
3 13 11 3
6 9 11 1 11 13 13
5 0 9 3 0 13
4 3 9 13 13
14 3 13 15 13 13 1 0 9 13 7 13 16 3 13
19 3 13 9 15 13 13 3 13 7 13 3 12 9 15 3 9 13 3 9
5 15 3 11 15 13
2 9 13
7 13 9 1 15 15 3 13
7 11 13 9 1 15 3 0
9 1 15 3 15 0 13 7 15 13
7 11 13 13 1 15 9 13
6 15 13 13 1 9 13
15 15 15 0 1 9 13 3 7 3 1 0 0 8 15 0
6 13 3 0 1 0 0
6 15 1 0 15 13 9
6 11 15 15 13 13 9
9 0 9 0 9 7 15 0 3 13
2 13 13
3 15 3 0
2 3 13
2 3 13
6 7 3 16 13 0 13
1 15
2 0 13
4 0 13 13 15
7 7 0 13 13 7 6 3
19 3 1 15 7 16 0 13 15 13 13 3 15 7 16 3 13 15 3 13
8 1 0 9 15 11 15 11 13
4 0 13 8 8
6 9 11 13 1 15 13
7 15 13 9 7 9 15 11
8 11 3 15 13 13 15 9 13
10 11 1 9 15 3 13 3 1 9 13
3 11 13 15
6 11 13 15 0 7 13
1 13
1 13
3 3 15 13
26 7 16 3 0 9 15 9 9 9 3 13 13 7 13 13 0 13 16 13 0 16 3 13 13 3 13
5 11 3 15 13 9
5 11 13 3 13 9
12 13 3 15 3 13 13 1 15 3 15 13 13
2 13 9
7 16 13 13 13 1 9 9
8 16 9 13 1 11 15 3 13
7 1 9 0 3 1 15 13
8 3 3 9 0 16 15 13 13
11 3 3 16 13 15 0 1 15 13 8 13
33 3 3 0 15 9 9 13 16 16 15 15 15 13 13 13 13 13 9 15 1 9 13 3 7 13 7 3 3 13 3 9 15 13
8 11 9 9 7 9 1 9 13
7 0 15 9 1 0 9 13
8 0 3 15 3 13 3 9 0
5 0 3 13 13 13
9 7 16 13 15 13 13 1 15 3
16 15 16 15 13 3 3 3 13 13 13 16 13 16 13 16 13
8 7 13 9 7 13 16 13 3
10 16 13 11 13 15 3 13 15 9 13
5 13 15 3 3 3
8 9 11 1 0 9 1 3 13
4 1 11 9 13
10 9 0 7 3 13 15 7 13 3 0
3 13 7 13
7 1 9 0 15 15 15 3
28 0 13 7 0 13 0 3 13 16 3 13 0 9 9 9 13 15 0 13 9 0 3 3 0 16 3 1 9
12 3 3 0 1 9 13 15 16 3 13 13 13
12 7 3 0 13 13 9 16 13 13 1 9 13
11 3 3 9 9 9 0 9 11 13 16 13
24 3 13 3 3 3 13 15 1 13 3 9 9 0 13 13 16 3 9 13 3 13 9 13 13
9 7 13 3 16 9 9 9 13 13
16 7 16 3 3 13 3 3 13 1 9 3 13 15 7 13 13
20 3 0 15 9 0 9 3 1 9 13 13 9 13 9 13 9 3 15 13 13
5 9 0 0 9 13
7 0 9 13 0 0 3 9
20 15 3 13 13 13 15 3 0 1 9 0 1 9 9 0 13 3 0 3 0
3 3 13 13
10 3 15 3 15 3 15 3 15 13 13
8 6 9 12 11 0 0 3 3
46 3 16 13 1 9 13 3 3 13 13 7 3 11 16 11 7 11 16 11 0 15 9 13 13 0 13 13 9 3 15 0 15 1 15 13 7 13 9 9 3 13 3 1 0 9 13
20 16 15 13 1 0 9 15 0 9 13 13 3 0 13 9 16 13 15 13 9
22 3 0 1 0 9 11 9 3 13 0 16 0 9 3 13 1 9 15 15 13 13 13
33 15 6 0 16 7 15 15 3 13 3 13 7 13 3 0 9 3 7 0 1 9 7 3 0 9 16 15 9 9 9 7 9 13
8 3 3 9 15 13 0 9 13
25 15 16 9 1 9 9 13 16 13 0 9 9 9 13 13 11 9 15 13 13 9 16 13 1 11
8 0 16 3 13 9 13 3 13
2 15 13
7 13 15 15 15 9 9 13
6 3 3 9 15 13 13
8 11 13 15 15 13 13 1 15
4 15 0 13 13
7 9 13 15 0 13 15 9
11 15 3 15 13 3 3 9 1 9 0 13
12 0 9 9 9 3 15 16 15 1 9 13 13
3 11 15 13
3 11 13 3
13 15 15 13 3 15 13 15 1 9 13 16 13 13
4 3 13 11 13
6 13 3 16 0 13 13
5 3 15 9 3 13
1 13
1 13
3 15 13 0
6 15 9 13 0 13 13
17 16 13 15 13 1 9 9 0 9 1 15 15 0 13 9 13 13
12 16 3 3 9 15 7 9 13 13 15 1 0
8 15 3 0 3 9 3 9 13
9 9 13 15 7 15 7 11 1 15
16 0 16 0 3 13 3 13 16 15 13 15 15 0 9 15 13
29 0 7 1 0 9 16 0 13 13 0 3 3 3 0 3 1 9 3 9 13 7 13 15 15 1 15 9 13 13
13 15 16 3 13 3 15 15 13 7 15 3 13 13
17 3 3 15 13 16 1 9 0 7 9 1 15 9 7 9 15 13
6 9 0 15 1 9 13
11 1 9 7 1 0 9 15 0 0 9 13
15 15 3 3 3 15 15 13 9 7 3 1 9 0 13 13
1 13
3 13 9 9
14 1 0 9 13 16 15 0 9 15 13 3 3 13 13
11 3 15 7 9 9 13 15 7 9 7 9
2 3 13
7 13 15 13 15 16 15 13
26 0 1 11 15 13 13 15 15 13 13 0 0 1 0 11 13 0 13 15 15 0 13 3 13 0 3
11 7 0 13 0 13 16 15 13 15 1 15
10 7 0 13 1 15 16 16 0 13 9
6 9 15 7 9 3 13
10 15 15 9 15 9 15 9 9 13 13
18 1 9 0 15 13 1 15 13 3 0 9 15 9 1 15 15 13 15
4 9 3 9 15
10 7 15 3 13 13 0 11 3 7 13
13 3 13 3 15 9 13 13 7 3 13 0 15 13
14 9 11 0 9 7 3 0 9 7 3 3 0 15 13
7 1 15 13 13 15 9 13
18 3 16 0 9 15 13 7 16 13 9 9 3 13 15 13 0 13 13
37 3 3 0 15 13 13 11 15 9 3 15 9 13 13 7 1 0 9 13 1 15 13 9 7 15 13 15 7 9 3 3 13 15 15 13 13 15
22 15 3 3 15 15 13 13 3 13 0 9 15 13 0 7 15 1 0 9 9 7 13
16 1 15 15 3 13 13 1 0 9 0 9 15 13 9 7 13
13 7 8 15 9 3 0 9 13 7 13 7 11 13
6 0 1 15 13 7 13
13 15 1 9 16 15 13 3 3 3 13 16 13 13
3 16 13 13
3 16 13 13
20 0 3 13 15 15 1 9 7 9 15 15 7 0 13 15 1 9 7 9 13
6 9 9 0 9 3 13
7 9 3 15 9 9 0 13
13 0 15 13 15 16 9 3 13 3 13 0 13 11
3 13 16 13
16 15 11 9 13 3 15 15 13 16 15 0 3 7 0 13 13
13 13 3 15 7 3 13 3 13 9 15 0 7 0
11 7 9 13 3 13 3 3 9 0 3 9
20 11 0 0 15 9 11 16 13 13 13 15 13 16 1 15 9 9 11 9 13
33 3 13 1 9 9 7 1 15 3 9 13 3 13 9 1 0 9 13 16 13 15 0 13 1 15 9 1 11 9 13 15 7 13
8 0 11 1 9 13 0 1 11
5 9 13 1 9 13
14 13 11 3 13 15 3 1 11 13 3 7 0 3 3
2 13 13
10 3 11 11 9 11 9 15 1 11 13
26 15 0 13 13 11 9 13 16 15 9 13 3 7 3 15 13 13 16 3 11 11 13 0 16 13 9
6 1 15 15 11 9 13
42 13 11 9 13 1 15 15 11 13 3 7 1 15 3 3 11 13 13 16 13 9 9 16 1 9 1 9 11 11 13 1 15 9 11 13 15 13 0 9 1 11 13
15 13 9 9 16 11 16 13 13 15 1 9 13 1 9 13
8 15 13 15 1 9 0 13 13
12 15 7 3 13 13 16 11 9 3 1 11 13
7 3 9 9 1 9 13 13
16 3 0 15 15 13 1 9 0 13 3 15 3 13 13 7 13
18 3 11 1 9 15 13 15 1 9 3 13 16 13 9 7 0 9 13
37 3 15 1 9 3 0 3 9 13 15 13 11 11 1 15 13 13 1 15 13 11 11 0 15 1 11 11 13 11 11 15 9 13 13 3 9 13
19 15 3 13 7 13 9 13 9 9 15 13 11 11 15 7 11 9 13 13
16 3 9 13 1 11 11 11 1 9 7 16 13 13 13 9 13
12 15 15 3 15 15 13 13 3 13 7 3 13
7 9 3 0 1 15 9 13
4 7 3 9 13
3 3 9 13
3 3 13 13
2 15 13
3 15 15 0
19 15 3 1 0 9 13 9 7 3 13 13 3 7 3 9 15 0 9 13
16 11 1 11 13 15 13 1 9 7 9 1 15 9 15 9 13
11 15 13 9 9 9 9 15 1 9 13 13
4 13 16 15 13
22 3 3 15 13 13 1 15 1 9 1 15 9 15 1 15 13 0 9 0 15 9 13
15 7 15 13 1 0 13 15 0 13 3 3 13 7 16 13
6 3 3 0 13 3 13
8 7 15 13 9 0 8 8 8
28 3 6 0 15 9 11 3 0 9 3 3 3 3 15 9 1 9 13 16 1 11 9 7 1 0 9 9 13
13 3 13 3 7 3 3 7 3 3 7 3 13 13
11 15 15 0 13 1 15 15 13 13 3 13
4 7 15 15 13
7 3 3 13 15 1 0 9
3 3 15 13
11 0 1 9 15 13 1 15 3 0 15 3
4 9 0 15 0
6 0 15 9 15 0 9
14 15 3 9 7 9 7 9 15 13 0 9 9 13 13
2 3 13
8 7 13 15 15 9 7 13 9
3 13 16 13
11 15 1 9 15 13 13 9 16 15 3 13
11 15 3 3 13 16 1 9 11 13 9 13
13 0 9 15 1 13 16 1 15 1 15 9 0 13
23 9 15 9 13 16 3 13 9 3 1 15 9 3 13 13 3 1 9 11 3 3 9 13
24 7 3 13 1 0 9 16 15 13 13 15 11 13 1 15 3 3 13 15 0 9 13 1 11
14 3 3 1 15 3 13 16 1 15 13 9 0 9 13
10 9 13 0 13 7 0 9 15 9 13
3 13 16 13
3 13 3 11
12 3 0 9 13 3 15 13 9 16 15 13 13
5 3 3 3 15 13
17 7 15 13 16 1 15 11 3 13 3 15 0 1 9 13 9 15
13 7 3 16 13 1 0 9 7 9 15 9 13 13
10 16 15 3 13 13 7 13 15 13 13
15 9 15 3 13 3 9 13 16 1 11 3 15 13 3 13
21 3 9 11 1 13 1 9 9 16 3 11 1 15 13 13 7 16 11 13 3 13
9 3 15 13 16 15 13 16 3 13
7 3 13 3 7 15 13 13
6 15 15 11 3 13 13
8 15 1 9 1 15 15 0 13
3 7 0 3
4 13 3 16 13
8 11 15 7 3 7 0 13 9
5 1 15 15 13 13
9 16 3 13 11 3 15 13 3 13
13 16 13 1 9 16 13 15 13 1 13 15 13 13
13 3 15 13 16 16 15 0 3 13 16 0 9 13
4 15 3 0 13
8 9 15 15 15 3 15 0 13
3 13 16 13
30 3 13 15 0 16 15 11 7 11 13 13 15 7 1 0 13 1 15 7 16 1 11 13 7 1 0 9 15 9 13
7 15 9 13 1 11 3 11
3 15 15 13
5 15 3 3 7 13
4 13 3 1 0
3 11 13 3
20 0 9 9 15 15 1 15 9 13 7 15 9 1 9 0 0 9 15 9 13
11 13 9 15 3 13 16 13 3 15 9 13
3 13 3 9
4 9 13 3 13
11 13 15 0 9 3 3 0 1 9 3 0
8 7 9 9 16 13 3 13 0
6 3 1 11 7 0 9
3 3 1 15
4 13 3 13 0
5 3 16 13 11 13
5 3 3 13 16 13
12 16 15 1 9 13 12 13 16 1 15 9 13
11 0 3 13 16 15 3 15 9 9 7 13
16 15 3 13 15 15 13 3 16 9 0 3 13 15 15 13 13
31 3 13 16 13 9 15 1 15 13 1 0 9 7 9 3 3 9 15 3 0 16 7 15 9 13 7 15 1 0 9 13
6 15 13 9 0 13 13
11 0 9 13 3 3 1 9 3 1 9 9
16 1 9 0 13 15 13 15 15 13 15 9 15 13 13 13 9
8 15 16 0 13 3 16 13 13
10 3 7 13 1 11 7 3 1 11 13
17 9 3 1 11 3 9 15 13 7 16 1 9 3 15 13 13 13
14 15 3 15 3 7 15 9 13 3 7 3 13 13 13
22 15 3 3 1 15 7 0 13 16 15 9 15 3 15 9 9 3 3 0 9 9 13
3 13 15 13
3 13 16 13
3 13 3 11
28 11 13 13 1 15 15 1 9 1 11 3 13 13 16 7 11 3 13 0 0 9 7 9 0 13 16 3 13
9 3 0 3 13 11 16 3 11 13
21 0 13 7 11 3 13 3 7 1 0 9 15 0 13 3 15 1 11 3 3 13
15 16 15 0 9 13 3 13 13 16 3 13 0 3 13 0
10 7 0 13 3 13 3 0 16 13 3
19 3 3 15 15 9 0 13 7 13 3 3 0 13 9 3 15 9 0 13
15 7 7 9 0 13 7 0 0 3 15 13 3 15 9 13
6 3 11 9 15 3 13
10 9 13 1 11 1 11 11 15 3 13
19 3 3 0 1 0 15 9 7 9 0 9 13 13 11 13 3 7 13 15
4 11 11 3 13
8 9 15 7 11 13 1 15 9
18 9 1 9 0 3 3 15 13 13 3 15 7 13 7 1 15 13 13
6 11 3 13 13 13 15
5 11 15 13 13 9
1 13
2 3 9
30 1 9 15 9 13 15 9 15 9 13 15 16 0 7 0 9 13 13 3 3 3 13 1 9 3 1 9 15 9 13
10 15 3 9 13 7 13 13 3 3 13
15 7 3 3 3 13 3 7 0 9 15 9 15 1 3 13
25 3 16 15 13 7 13 9 13 13 15 9 15 9 13 3 3 9 16 15 13 15 13 0 3 13
12 15 7 15 9 9 7 9 1 9 1 13 13
6 15 0 15 13 7 13
5 11 15 0 9 13
8 9 9 15 1 11 13 13 15
31 11 9 16 1 11 13 1 3 7 11 13 3 3 13 15 13 16 15 0 13 9 16 15 3 13 15 0 15 9 3 13
53 3 15 13 13 11 3 1 15 13 7 3 13 3 15 0 13 1 15 9 9 15 13 13 9 13 3 13 16 7 0 0 15 0 9 0 1 9 13 7 15 9 9 13 7 13 9 0 13 7 1 0 13 13
13 7 3 0 13 15 3 13 16 1 15 13 3 13
17 13 15 9 0 1 9 3 0 7 9 13 7 9 13 1 9 15
9 0 9 9 0 9 3 13 9 13
8 1 0 15 9 15 13 9 13
5 3 15 9 13 9
13 3 15 15 9 13 1 15 3 15 0 13 3 13
12 13 15 11 3 13 15 9 15 9 15 9 13
7 7 15 1 0 15 3 13
12 3 13 15 13 15 13 15 3 9 7 0 13
13 3 16 3 13 15 13 13 15 7 9 15 13 13
15 16 3 15 13 0 13 15 0 9 13 3 13 3 0 13
5 11 15 3 13 9
11 15 3 12 1 9 1 9 13 9 0 9
13 15 3 3 0 9 7 9 9 3 15 13 11 13
12 15 16 3 13 3 11 13 13 1 9 15 13
7 9 15 1 11 13 15 13
3 13 3 11
10 13 15 13 3 1 3 13 1 15 9
6 0 13 3 15 13 11
7 15 13 3 13 13 3 13
9 16 3 15 13 0 13 15 15 13
8 3 3 15 15 13 3 9 0
15 3 15 15 15 13 13 7 3 3 15 15 13 13 15 13
25 3 16 15 3 3 7 3 3 13 7 9 0 13 13 13 15 0 0 13 15 1 15 9 3 13
20 15 3 3 1 0 9 3 1 0 9 0 9 9 9 9 0 9 0 15 13
19 13 13 15 13 3 13 15 13 15 13 9 15 9 15 9 15 9 15 9
37 15 15 16 0 9 9 13 16 0 13 3 15 0 3 7 13 13 16 13 16 7 0 9 9 7 13 7 15 15 0 0 13 0 0 13 7 13
3 3 9 13
32 3 3 3 13 13 16 13 7 16 13 16 0 3 7 13 15 3 13 16 1 9 15 1 15 9 9 13 7 3 0 3 13
37 0 3 13 16 3 13 15 15 13 3 16 9 7 9 0 13 3 7 1 15 3 0 13 16 7 9 13 7 16 13 3 3 13 3 15 0 13
17 15 3 3 13 3 0 1 9 1 15 13 13 16 3 3 15 13
3 13 3 11
24 15 7 15 9 7 15 0 9 3 0 3 9 7 9 15 9 7 16 15 3 13 3 11 13
16 16 13 9 15 13 16 9 13 15 15 9 13 1 15 15 13
8 15 15 3 13 9 9 9 13
3 13 3 13
3 13 3 13
10 15 16 13 3 15 15 9 7 9 13
6 11 9 0 0 7 13
8 1 15 13 15 16 15 0 13
2 13 3
2 3 13
18 3 15 15 13 16 15 13 16 3 13 13 16 15 3 15 15 3 13
4 9 13 1 9
10 15 0 13 0 9 9 7 9 9 13
7 13 3 15 3 1 9 13
16 13 3 3 15 13 16 0 0 13 7 3 13 16 3 13 13
3 3 13 13
8 15 16 13 15 13 13 13 13
5 16 3 13 3 13
13 15 3 3 0 1 9 13 1 9 15 1 9 15
9 3 15 3 13 13 16 1 15 13
11 13 15 3 13 3 3 9 3 13 15 13
9 3 13 0 13 3 7 13 15 13
3 13 3 11
4 15 15 11 13
31 15 1 9 16 9 13 13 15 7 15 1 15 13 3 13 3 16 13 15 13 3 7 15 9 3 0 9 13 13 3 13
17 15 3 9 15 13 13 15 15 0 13 13 15 13 15 13 15 13
7 1 9 9 13 0 9 13
13 15 16 13 3 13 16 13 15 9 15 9 15 13
27 16 15 3 13 3 0 15 9 3 3 13 13 13 16 3 15 13 13 16 15 3 3 7 13 3 7 13
17 3 16 13 15 13 15 3 9 9 1 9 13 15 3 9 0 13
23 3 16 13 11 15 13 15 3 1 15 9 13 0 13 3 15 15 13 15 13 9 13 13
5 11 9 15 13 13
11 15 15 0 16 0 13 3 15 0 13 13
2 13 3
14 1 15 9 0 13 9 1 11 15 1 15 13 7 13
5 9 3 13 13 13
8 15 13 13 0 13 13 1 15
23 16 15 0 13 13 15 13 13 15 9 16 13 15 15 0 9 3 7 15 9 13 13 13
9 13 15 15 0 9 1 0 9 13
16 15 16 15 9 15 1 9 13 3 3 13 15 13 7 3 13
14 15 1 9 9 7 0 9 9 0 3 13 15 3 11
22 7 3 13 3 1 11 3 15 3 13 3 1 0 9 3 13 1 13 1 0 9 9
23 1 11 3 3 13 3 13 16 3 15 0 9 13 7 9 3 15 13 3 3 3 11 13
10 3 16 15 1 9 13 15 1 11 13
7 3 3 13 3 3 7 13
3 13 3 11
17 3 16 15 15 12 3 1 9 13 15 15 13 15 7 15 7 15
13 7 16 15 0 15 13 3 1 15 0 9 13 13
18 13 13 15 9 13 13 3 3 16 3 13 7 3 16 13 0 9 15
15 0 13 3 7 0 9 13 13 15 3 7 1 0 9 13
11 9 3 3 3 3 13 9 0 7 3 13
5 3 0 9 13 9
14 0 3 13 3 7 9 0 9 7 9 0 9 3 13
3 15 3 13
34 3 16 13 15 15 15 15 13 13 7 1 15 11 15 3 3 0 13 1 0 9 13 16 3 13 3 1 15 9 15 3 0 9 13
10 0 16 13 13 15 13 13 15 16 13
4 7 0 3 13
6 11 9 15 13 3 13
6 1 9 9 3 13 13
3 7 15 11
5 15 3 13 13 13
12 7 11 0 9 13 1 15 9 3 3 13 11
7 15 16 15 13 3 3 13
5 11 9 13 9 11
7 7 3 0 11 13 1 9
9 15 3 3 15 9 3 15 13 13
44 15 16 15 3 15 7 9 0 9 13 3 13 16 3 13 12 1 15 9 15 7 9 7 9 15 3 3 13 13 13 3 3 13 16 15 3 15 3 9 7 9 15 13 13
6 1 15 3 0 13 3
50 3 7 0 3 13 16 15 3 15 9 0 9 13 13 13 7 3 16 3 15 13 7 13 3 13 13 7 13 3 13 13 15 15 15 13 13 9 3 7 13 13 15 13 0 15 13 9 1 9 13
13 7 15 3 9 13 9 15 15 13 9 3 0 15
32 3 16 3 3 15 7 15 13 15 15 11 3 0 9 13 1 0 9 13 15 0 15 13 3 13 7 13 3 7 9 3 13
3 3 15 13
6 15 3 0 3 3 13
11 3 15 3 15 0 7 16 15 9 9 13
15 16 15 1 11 13 1 9 13 13 15 7 3 13 3 13
7 16 3 15 13 3 13 0
10 16 13 15 13 3 13 0 9 9 13
8 3 7 15 15 9 13 3 13
17 15 16 3 13 13 13 13 7 3 13 13 13 13 3 15 3 13
9 3 15 3 15 9 13 7 3 13
21 0 0 13 13 1 9 13 1 9 13 15 16 3 15 1 13 13 13 13 0 13
9 3 13 0 15 13 15 13 7 3
4 3 3 13 15
12 1 15 0 0 13 15 9 13 16 3 9 13
7 15 3 13 13 13 7 3
3 1 9 3
6 3 3 11 15 13 13
16 3 3 15 15 15 13 7 1 9 13 7 16 13 13 11 13
3 15 1 9
3 15 1 9
3 13 3 13
8 7 16 3 13 15 3 3 13
9 0 16 13 13 15 1 9 15 13
9 16 3 9 15 13 15 13 15 9
80 3 11 16 15 13 15 9 1 9 15 16 7 1 15 0 3 13 9 13 7 15 15 3 15 13 3 16 3 13 16 7 15 13 13 13 1 9 15 15 9 13 0 11 3 13 1 15 13 13 7 13 15 15 15 13 9 13 7 13 15 15 16 3 3 9 13 3 15 3 13 3 16 13 13 13 7 1 15 15 13
11 15 16 15 9 13 3 15 3 15 9 13
13 15 9 13 16 15 1 15 3 13 3 15 13 13
24 3 16 13 9 0 9 0 13 15 3 1 9 13 13 0 9 15 3 1 9 15 13 3 13
42 3 13 16 15 1 15 13 7 13 13 15 7 3 13 13 13 15 16 15 13 7 15 13 13 3 13 3 13 7 16 0 9 3 15 7 15 0 1 15 13 13 13
16 16 15 13 15 13 9 13 15 9 9 13 13 13 13 7 13
2 13 3
10 0 9 15 0 13 9 9 15 3 13
15 3 15 13 3 16 1 15 15 13 3 13 15 13 3 13
2 13 3
15 1 11 9 9 15 0 3 7 0 13 1 3 3 1 3
13 15 3 9 11 11 11 9 1 15 1 11 13 13
22 15 3 9 15 13 13 13 7 13 3 9 1 11 11 9 15 7 15 1 9 9 13
19 7 3 11 9 13 15 1 15 9 13 3 3 13 1 9 3 9 11 13
14 3 13 1 15 0 9 0 7 3 3 16 11 9 13
16 0 15 1 15 0 9 13 1 15 9 13 13 0 3 15 13
10 13 1 15 9 15 15 1 15 12 13
12 15 15 7 13 15 13 7 13 9 15 3 13
11 3 13 9 13 15 9 16 0 9 15 13
5 15 9 3 3 13
14 1 15 13 13 16 7 9 15 15 0 7 9 0 13
2 13 3
30 9 15 3 0 13 16 13 11 15 1 9 13 9 15 11 3 13 7 16 1 11 15 9 15 13 13 13 9 3 13
14 3 15 15 13 7 13 13 11 9 7 13 15 1 9
19 16 13 15 1 9 13 7 16 13 13 9 15 15 13 1 0 9 15 0
19 3 11 9 9 0 15 15 3 3 13 15 13 9 0 13 13 9 9 15
5 15 3 9 13 0
10 3 7 3 15 13 13 3 7 3 13
11 13 13 15 16 15 15 13 1 15 13 13
20 3 0 9 15 9 1 15 13 16 15 1 15 13 13 9 7 9 11 13 13
28 16 15 9 0 9 13 15 13 1 11 13 13 16 7 9 15 9 13 7 16 13 15 1 0 9 13 3 13
27 7 7 1 9 3 1 15 9 13 7 16 15 13 13 3 3 0 0 9 7 13 7 15 3 13 3 13
2 9 13
10 15 15 9 3 1 0 9 13 15 15
11 7 3 15 9 3 0 3 13 3 15 9
48 7 3 16 13 13 13 15 9 13 13 7 15 1 9 3 13 3 7 0 7 0 9 0 7 0 9 3 7 11 0 7 9 3 7 9 0 9 9 3 7 0 9 11 9 7 0 9 15
11 15 11 7 9 1 9 13 7 15 13 3
90 15 13 7 13 11 11 16 15 15 0 0 0 7 9 9 9 13 16 15 1 15 9 13 7 13 13 16 13 15 13 16 0 15 7 15 13 16 15 15 9 13 7 11 9 15 13 13 0 13 11 9 7 15 13 15 16 13 15 3 13 13 16 3 13 16 13 15 7 1 9 15 3 13 3 15 9 13 13 7 9 1 15 1 9 3 3 7 3 3 13
12 15 3 3 13 7 9 15 13 13 9 3 13
10 13 15 3 13 16 15 0 9 13 13
17 3 15 13 1 9 16 15 9 16 9 16 9 15 15 13 3 13
6 15 13 13 16 13 9
15 7 15 13 1 9 3 13 15 9 13 15 15 9 15 9
25 1 15 13 1 9 13 3 13 9 7 0 9 15 13 16 1 15 9 0 13 15 1 7 1 15
30 15 0 9 7 9 15 15 13 3 3 13 13 1 15 1 11 7 3 1 15 13 16 13 13 3 15 0 1 9 13
10 1 0 9 16 15 3 15 13 13 15
6 1 15 15 13 3 9
5 7 15 15 13 3
39 16 9 15 1 15 9 13 16 15 9 1 15 1 0 13 15 15 13 9 13 13 7 15 0 9 15 9 7 13 7 13 13 3 7 16 3 13 13 13
26 16 15 13 15 13 13 1 9 15 15 3 1 15 1 15 13 7 13 13 13 15 9 7 13 0 9
16 15 3 3 3 13 15 15 1 15 9 13 0 3 1 15 15
17 13 15 13 15 13 15 13 1 15 13 15 7 15 1 15 9 13
14 3 7 3 13 13 7 1 9 3 13 7 15 13 13
3 13 3 11
14 12 9 13 0 16 0 13 9 1 15 15 1 15 13
20 15 3 13 1 9 3 3 3 1 15 13 13 1 11 7 3 15 9 3 13
2 13 3
30 16 3 1 15 11 9 7 11 15 13 13 13 3 13 15 15 9 3 13 16 3 13 1 15 15 13 7 15 13 13
12 15 3 11 9 15 13 3 3 13 13 1 11
7 15 9 15 0 9 13 13
13 7 3 16 13 9 13 13 15 13 16 1 15 13
11 15 16 13 1 15 3 13 16 13 3 13
19 11 15 1 15 9 15 7 9 7 9 7 9 13 9 15 0 13 11 9
12 3 3 15 1 15 13 15 0 13 1 0 9
17 15 11 13 16 15 1 7 1 15 15 13 13 7 13 1 15 15
14 13 9 9 3 15 9 3 15 15 15 15 0 3 13
26 15 16 1 11 16 13 1 11 3 15 13 13 7 16 15 0 13 9 1 15 13 16 0 0 11 13
21 3 16 1 15 15 13 13 16 13 15 7 1 15 13 15 3 3 15 9 13 13
9 15 3 7 9 7 3 9 3 13
3 13 3 11
37 3 0 9 1 15 13 12 13 3 1 15 15 13 16 0 9 9 0 13 15 7 15 1 9 13 13 1 11 9 1 11 9 1 0 11 9 13
13 1 0 9 1 9 15 9 3 13 7 3 13 9
40 1 15 16 3 15 9 1 0 9 13 13 13 1 15 1 15 9 0 0 15 9 0 3 3 0 13 16 13 15 9 13 9 16 0 9 3 1 15 9 13
14 15 3 13 1 9 7 9 15 15 1 15 9 3 13
9 7 15 13 13 7 3 15 3 13
16 0 9 13 0 1 9 16 15 1 15 9 0 9 3 13 13
12 0 9 15 11 15 9 7 1 15 13 13 13
22 13 3 11 13 16 3 7 16 3 3 13 3 7 1 9 3 7 1 9 13 15 9
10 7 13 3 13 13 9 0 9 15 13
8 3 16 15 13 15 3 13 13
22 0 16 7 9 0 3 13 7 16 3 3 13 13 7 13 12 15 9 9 9 13 0
50 16 15 1 0 9 13 13 15 1 9 9 7 9 0 13 15 1 9 0 13 13 13 13 1 9 15 3 13 3 13 15 7 15 15 13 13 13 13 1 0 9 9 9 7 13 0 0 9 15 13
8 7 0 1 0 9 9 3 13
6 9 3 9 15 3 13
32 15 0 13 9 9 15 16 15 15 1 15 15 13 13 3 1 15 13 16 0 9 9 16 13 0 3 3 15 0 9 13 13
7 3 7 15 1 11 13 13
14 13 3 1 9 3 0 9 0 9 9 13 13 15 13
11 3 1 9 15 13 0 9 9 15 3 13
51 3 11 7 0 13 13 13 7 15 13 7 3 12 9 9 1 9 1 15 13 3 13 7 7 16 13 0 9 3 13 0 1 13 3 13 13 16 15 13 13 16 13 15 3 15 3 15 9 13 13 13
8 0 9 3 13 0 9 9 13
4 7 13 3 15
9 12 9 15 13 16 9 13 13 0
6 3 3 13 3 0 13
16 13 3 16 9 3 13 13 16 0 15 9 0 15 15 13 13
13 7 16 13 15 1 9 13 9 15 11 11 13 11
3 0 15 13
62 16 3 15 13 3 15 9 3 3 15 9 15 13 13 13 7 15 16 11 9 13 15 15 0 3 13 16 7 15 15 13 0 13 1 15 3 13 9 15 9 15 11 15 15 0 13 1 9 7 9 9 15 13 3 13 9 12 0 0 13 15 9
9 15 1 11 13 16 0 9 9 13
11 15 1 15 13 0 9 3 15 9 13 13
2 13 3
24 3 16 1 15 13 15 9 9 9 13 13 16 13 3 15 13 13 3 13 15 15 3 13 0
24 16 15 7 13 13 7 13 3 9 15 13 13 3 13 16 0 0 9 0 15 13 13 13 13
10 3 16 9 9 15 13 15 13 9 13
12 3 16 9 1 15 0 13 13 13 15 3 13
21 3 16 13 16 3 15 13 0 0 0 1 9 13 13 0 9 9 13 15 9 13
17 3 13 16 7 9 9 13 7 16 9 13 9 0 13 9 13 13
66 13 15 3 0 9 16 0 0 9 3 3 1 15 13 9 15 13 16 1 15 13 13 13 13 3 1 15 9 15 3 3 0 3 13 7 3 0 7 0 3 7 3 3 13 13 13 9 13 16 16 1 0 0 9 15 13 15 9 13 13 13 15 3 13 3 13
10 0 1 15 13 13 9 13 3 0 13
13 13 3 0 13 15 1 0 9 12 9 3 9 13
15 13 3 0 3 13 7 0 9 11 7 11 15 9 3 13
18 0 9 3 13 7 0 9 15 9 13 13 1 15 13 7 3 3 13
11 3 0 9 16 0 3 13 15 3 0 13
19 1 15 1 15 9 9 15 11 13 13 1 15 13 15 1 0 9 13 13
23 3 7 3 7 0 1 9 13 16 15 9 9 15 13 15 1 15 9 1 15 0 9 13
14 7 16 0 7 16 15 13 15 1 3 13 13 0 13
17 0 1 15 13 13 9 15 15 15 13 16 15 1 3 3 13 13
15 9 15 1 11 9 1 9 9 15 1 15 13 13 13 13
6 15 13 13 1 15 13
11 1 15 9 7 1 9 0 15 3 13 13
13 15 13 16 15 1 9 15 15 13 15 0 16 13
66 13 3 16 3 13 15 1 9 15 13 3 7 0 3 7 0 3 15 0 3 7 3 1 0 15 1 15 9 3 1 9 9 15 0 0 7 15 15 0 9 9 15 7 3 9 9 7 13 9 9 13 3 9 15 13 0 7 9 9 9 9 1 13 9 15 13
22 3 0 15 3 13 1 0 9 3 13 9 12 1 13 9 9 7 3 9 15 15 13
27 15 3 13 16 3 13 7 16 3 13 9 15 9 13 9 15 13 3 0 9 9 15 0 3 3 0 13
29 15 3 1 15 9 15 3 13 13 13 13 9 15 0 0 7 1 9 9 7 1 9 0 9 3 3 13 13 13
28 3 16 15 7 13 13 1 15 13 7 3 9 7 9 13 3 15 13 3 15 15 13 3 1 15 9 13 13
13 3 11 13 13 0 0 9 15 9 13 13 1 15
3 11 13 3
22 3 15 11 15 13 3 0 15 0 9 15 9 0 9 13 7 0 9 7 15 0 11
21 3 13 16 11 13 9 11 0 9 15 9 7 9 0 9 11 9 9 0 13 13
16 3 1 9 3 13 9 3 13 16 3 1 15 1 9 9 13
32 1 9 3 13 16 15 15 9 9 9 13 13 15 15 3 3 13 1 0 9 15 15 0 15 9 13 3 13 7 13 7 13
29 1 15 9 0 16 13 15 9 13 0 7 9 7 9 15 3 1 11 13 1 9 7 7 1 0 11 0 9 13
10 3 1 9 15 13 9 3 9 9 13
63 0 9 16 13 9 0 9 7 9 1 9 3 3 1 9 13 9 11 15 9 9 9 13 13 16 1 0 9 9 1 9 13 7 1 15 9 9 3 3 9 3 3 0 11 13 15 7 0 13 9 7 1 15 3 16 15 13 13 13 7 3 9 13
32 16 13 9 16 3 15 13 13 9 13 1 11 7 11 13 13 9 9 1 15 9 16 1 11 13 16 0 9 13 9 7 13
18 15 9 9 13 16 9 9 0 0 7 0 9 15 9 13 13 13 9
10 3 9 0 7 15 9 15 11 13 13
16 0 9 12 16 13 15 9 13 7 1 15 15 0 15 13 13
11 0 15 9 0 3 0 13 0 11 3 13
7 11 0 13 15 13 9 0
4 9 9 11 13
13 15 13 3 3 3 16 1 9 15 15 3 9 13
7 15 16 13 9 9 0 13
6 9 9 1 9 9 13
3 9 0 13
8 1 9 0 3 13 3 13 13
8 3 13 15 0 15 9 3 13
12 3 3 9 0 9 9 9 0 3 13 3 13
18 15 13 7 13 16 13 13 0 7 9 13 16 15 15 9 13 3 13
5 0 9 15 9 13
12 3 15 15 15 0 13 13 0 3 13 3 13
3 3 15 13
13 3 3 13 11 3 3 13 0 13 13 15 13 9
4 3 0 0 13
25 0 15 13 9 15 15 13 7 15 13 9 7 15 9 15 3 13 16 1 0 0 16 1 0 0
10 1 0 13 9 13 13 0 9 1 9
4 13 1 9 3
28 13 9 13 3 1 15 7 16 3 1 13 13 15 7 3 16 3 3 13 3 3 9 9 9 15 15 13 13
7 3 9 9 15 13 3 13
8 15 15 16 3 13 3 13 3
8 15 3 13 16 9 15 13 13
10 3 3 0 1 9 13 15 11 15 13
14 13 3 9 9 1 15 13 15 3 9 13 1 9 13
11 13 16 15 7 11 13 7 15 9 9 13
4 3 13 9 0
6 13 15 9 15 13 9
16 1 15 11 15 13 0 15 9 0 13 13 15 13 1 13 13
29 3 11 11 1 15 9 9 13 9 9 9 13 9 13 9 15 7 9 15 1 9 13 1 9 1 9 13 1 9
13 16 13 9 9 1 9 11 15 1 12 13 11 13
7 1 9 3 0 9 13 13
42 16 9 0 13 9 13 15 9 13 9 11 13 9 9 1 15 9 13 16 15 9 13 13 9 13 15 9 13 13 15 9 9 13 11 13 7 11 1 15 0 9 13
7 13 9 15 1 9 9 13
4 0 9 15 13
2 3 13
3 13 3 3
10 3 9 9 13 13 0 15 1 15 13
8 0 9 9 3 13 13 0 15
22 15 9 9 9 1 9 9 13 9 3 0 3 3 0 9 12 12 0 3 12 12 12
13 15 9 3 3 3 1 0 15 7 3 1 9 13
1 13
4 15 3 9 13
13 13 0 3 9 15 16 3 7 13 3 7 3 13
5 3 0 3 3 13
20 3 0 15 11 11 0 13 0 15 3 15 3 13 15 15 9 13 13 0 13
5 15 3 1 15 13
10 15 13 16 3 9 11 15 15 7 13
10 16 13 15 13 13 1 0 15 9 13
12 15 15 1 11 13 3 13 13 16 15 9 13
22 15 16 13 15 13 0 16 16 9 9 0 9 13 13 13 0 9 13 3 15 9 9
25 7 13 15 9 13 7 13 7 13 9 13 7 3 15 13 1 9 9 1 15 3 13 3 0 13
8 7 0 3 9 0 15 9 13
4 0 3 3 13
11 13 0 15 15 3 7 13 13 3 7 13
2 0 13
3 0 3 13
18 9 9 13 13 1 0 9 15 15 13 1 9 15 13 15 0 15 0
6 15 1 9 3 3 13
6 0 15 15 13 8 13
6 13 1 9 7 1 9
2 15 13
9 0 9 3 13 13 9 1 9 15
15 13 9 11 15 1 9 9 9 9 13 7 1 9 3 13
10 11 9 9 3 13 9 9 1 9 15
9 1 0 3 9 15 3 9 9 13
2 3 13
5 9 3 9 9 13
15 3 3 16 9 13 13 0 3 0 0 7 9 7 3 9
2 13 13
6 13 3 15 9 13 13
15 1 0 9 9 9 13 1 15 3 3 11 9 3 11 13
17 13 16 15 15 13 3 13 9 15 9 0 3 3 13 1 9 13
11 3 3 16 0 9 13 13 13 15 1 15
4 9 9 9 9
3 0 0 15
5 13 1 9 11 11
8 15 13 15 1 3 9 9 13
2 9 13
29 3 11 9 0 15 13 1 11 3 13 7 13 3 13 13 16 3 9 0 1 9 9 13 9 15 1 13 9 13
11 0 9 11 11 1 9 15 1 0 9 13
10 3 1 0 11 9 11 11 13 9 0
7 13 9 1 15 9 0 0
9 0 13 7 0 15 1 0 9 11
3 3 9 3
2 3 11
18 11 9 13 9 13 13 11 3 6 9 15 1 15 9 9 15 0 9
2 11 13
9 0 3 16 9 15 3 13 9 13
34 11 13 11 9 15 0 1 9 3 13 16 0 15 9 9 9 9 15 9 13 15 7 15 9 13 13 15 1 15 9 0 1 9 13
3 9 0 11
2 0 11
2 0 11
10 0 3 0 16 11 1 9 13 9 13
12 11 16 13 9 13 9 1 9 13 3 13 13
10 11 13 1 9 0 9 9 0 1 9
4 9 9 12 0
2 13 9
2 13 9
10 11 3 13 16 15 0 9 1 9 13
7 15 13 16 1 9 9 13
6 15 9 0 1 9 13
5 13 1 9 9 11
1 13
9 0 15 13 0 7 0 11 11 9
2 3 9
3 9 9 15
7 3 0 15 13 9 9 0
4 11 9 3 13
6 11 9 0 3 15 13
2 0 9
16 15 9 15 0 13 13 0 15 1 0 9 13 9 15 3 9
3 13 9 13
8 0 15 0 13 7 0 0 13
4 9 13 3 13
10 9 11 16 3 13 13 13 1 11 13
3 3 13 13
3 1 15 13
14 3 3 15 0 7 0 9 13 13 3 7 0 9 13
9 15 9 3 13 3 3 3 16 13
4 9 0 13 13
16 11 9 3 9 1 9 15 16 3 13 13 0 13 9 9 13
10 15 9 1 15 15 9 13 15 0 13
7 0 15 11 13 3 1 9
13 13 3 15 15 13 1 11 15 7 1 15 9 13
28 15 1 15 9 13 13 3 16 13 15 15 3 3 3 0 13 7 16 0 0 13 15 15 9 0 0 7 13
3 0 3 13
3 0 13 13
9 15 9 13 3 1 15 1 15 13
6 3 13 16 1 15 13
33 7 13 15 13 1 15 9 12 15 15 11 13 9 1 0 9 15 7 13 16 13 9 1 15 9 13 15 15 0 3 13 8 13
6 7 0 16 15 13 0
14 0 3 3 13 13 16 13 1 0 9 13 7 11 13
8 3 3 7 0 13 7 13 11
4 9 13 13 3
8 16 13 13 12 0 9 0 13
3 7 0 3
3 13 3 15
12 15 13 1 15 13 15 13 13 7 3 1 15
5 3 3 15 13 3
10 13 1 15 1 15 13 7 3 13 9
1 15
6 7 13 0 0 0 9
19 3 13 0 15 13 9 1 0 9 3 13 13 7 3 13 16 15 13 9
6 13 13 13 13 1 15
11 3 0 13 9 16 1 15 1 9 0 13
4 0 13 15 13
5 3 3 15 9 13
11 13 15 15 13 13 15 13 3 3 16 13
26 15 6 15 9 13 13 0 0 9 16 15 15 13 13 1 0 15 3 3 3 13 15 13 3 13 13
19 13 0 16 7 0 3 13 7 15 13 15 9 15 3 13 13 15 11 13
6 15 9 13 13 15 13
3 13 13 13
20 7 15 1 0 16 15 9 13 15 3 0 13 13 13 3 15 1 11 9 13
2 9 13
16 16 15 15 13 15 15 13 13 13 9 16 1 15 15 13 13
1 13
3 13 3 3
9 9 15 16 3 13 13 15 3 0
3 9 11 13
6 15 1 9 0 1 9
4 13 3 1 15
2 3 3
3 15 3 15
2 7 13
7 9 15 15 13 9 7 9
7 1 11 3 3 13 3 13
49 9 0 7 0 9 7 1 0 9 9 0 9 13 13 15 7 0 0 7 0 3 13 16 15 9 3 13 3 16 11 7 15 7 6 16 3 13 9 16 15 15 9 9 13 1 15 9 13 13
7 3 15 0 15 9 3 15
12 3 15 3 16 13 9 3 3 15 13 0 9
3 0 13 9
3 15 13 3
12 0 3 0 16 3 13 3 13 16 3 0 13
9 15 16 13 13 7 1 9 9 13
7 3 13 3 15 3 13 13
3 3 13 13
10 15 3 0 15 3 3 13 3 13 13
3 0 3 13
2 8 8
2 8 8
11 3 6 13 7 11 13 15 13 1 9 13
13 1 15 9 3 1 15 13 13 7 15 12 9 13
11 9 3 0 3 13 15 3 11 13 13 13
3 6 0 9
6 7 0 3 13 3 0
3 15 3 0
15 16 15 13 16 13 0 0 1 15 13 3 0 0 9 15
42 7 6 1 13 13 16 15 13 3 0 9 9 3 13 3 3 9 0 13 0 16 15 13 7 3 16 8 15 15 1 13 13 1 13 13 0 7 15 9 9 13 13
7 15 3 3 3 1 15 15
41 9 11 3 15 13 15 15 9 16 13 13 13 16 1 15 13 3 9 13 15 7 16 13 13 7 16 15 15 3 13 13 13 9 9 15 3 13 13 11 15 13
14 15 8 9 15 15 15 0 1 11 15 9 0 3 13
5 13 9 12 3 11
3 0 9 13
20 1 11 16 13 15 0 9 13 9 0 15 13 7 0 13 15 13 15 9 0
4 3 11 15 9
5 15 9 15 9 13
3 15 3 13
13 15 9 13 16 11 13 9 13 3 3 16 13 15
4 1 15 13 0
5 15 9 1 9 13
2 9 13
2 11 13
2 15 13
2 3 13
5 8 8 8 8 8
10 15 13 3 9 11 13 7 13 3 13
11 3 1 9 16 13 8 8 8 8 8 8
6 13 15 1 9 15 13
16 1 9 13 15 1 15 13 0 13 3 0 7 0 3 15 9
2 15 0
2 15 0
2 15 0
5 8 8 8 8 8
12 3 3 16 11 15 9 13 9 13 13 15 9
11 15 0 3 0 15 9 16 15 9 9 13
1 13
6 3 13 3 16 15 13
5 11 3 13 16 9
2 15 13
7 13 3 13 16 9 3 13
4 13 13 15 3
5 3 3 15 13 13
15 9 3 16 9 13 13 3 3 3 3 0 9 1 11 13
30 1 11 8 8 8 8 8 8 8 8 8 8 3 13 0 8 15 7 16 1 0 7 16 1 9 7 16 9 0 3
5 12 0 16 0 3
8 3 1 0 9 13 16 0 0
30 15 3 0 3 3 15 15 3 9 3 13 13 9 13 13 9 3 13 3 16 7 0 7 3 3 3 3 1 0 13
35 16 3 0 13 15 13 16 13 16 3 3 0 3 1 9 0 13 9 9 13 3 13 15 0 0 3 9 0 1 15 3 13 3 0 15
7 1 11 1 15 3 13 9
2 13 9
1 13
16 1 11 11 15 13 13 9 0 3 15 13 3 7 15 3 9
8 3 3 0 7 0 7 0 0
6 15 16 3 13 13 13
11 13 1 11 10 0 11 13 9 7 13 0
2 13 9
1 13
3 0 3 9
11 15 13 16 15 1 15 13 16 3 13 13
17 1 15 15 15 13 16 7 8 15 13 7 8 8 8 13 3 13
11 7 9 13 0 9 15 1 15 3 13 13
25 15 13 1 11 16 15 13 9 13 7 0 9 15 13 7 1 15 1 0 9 7 1 15 3 13
8 3 15 13 15 13 15 0 13
3 13 16 13
21 3 13 13 3 9 13 9 9 13 13 3 0 9 0 7 1 9 15 13 15 13
5 15 3 1 11 13
8 15 3 9 13 16 9 13 13
7 1 15 3 3 6 13 13
8 13 3 1 15 1 0 1 15
10 15 3 13 15 13 13 3 11 9 13
8 1 15 0 16 15 13 13 13
14 16 11 13 15 15 9 13 7 9 15 16 3 13 0
16 11 9 1 15 13 15 16 11 0 15 1 13 1 15 3 13
5 0 9 11 1 11
8 11 0 13 9 11 13 1 9
6 16 15 13 0 13 13
5 15 3 13 9 11
8 3 15 13 0 9 0 7 0
4 3 0 3 13
48 7 6 16 1 0 9 13 7 9 1 9 0 3 9 13 7 13 13 7 1 0 15 9 15 13 1 9 11 13 3 1 0 9 0 15 1 7 1 15 13 3 1 15 15 1 13 13 13
26 15 9 7 0 15 7 15 0 13 13 15 13 13 7 13 11 16 13 16 13 15 15 1 0 9 13
5 11 1 0 9 13
8 1 15 3 3 13 16 0 13
10 13 15 9 15 15 13 12 9 12 3
2 13 0
4 13 13 0 15
7 3 0 15 9 13 13 13
10 13 15 11 11 1 15 1 0 13 3
14 15 16 13 11 15 7 15 3 13 16 9 1 9 13
3 13 9 3
17 15 15 9 13 7 3 16 13 7 16 15 11 13 1 15 13 13
17 15 3 13 9 1 9 0 3 6 13 11 15 15 15 7 15 13
5 8 8 8 8 8
21 3 16 9 0 3 13 1 15 15 0 9 15 0 15 9 15 11 15 0 9 0
12 3 3 16 3 13 3 9 0 3 15 9 13
15 15 15 1 1 11 13 15 3 7 13 3 16 15 9 13
4 1 15 9 13
5 15 11 15 9 13
3 11 11 13
10 7 15 1 15 1 9 11 3 11 13
6 3 15 13 1 11 13
6 11 3 13 3 13 13
8 9 3 9 11 13 7 9 3
9 0 15 16 11 0 13 13 15 13
10 7 16 15 13 3 13 1 15 1 11
3 3 15 13
4 13 9 9 9
8 3 9 13 16 13 3 3 11
5 9 15 15 0 13
8 15 1 0 13 3 13 15 13
5 3 11 15 3 13
4 11 3 13 13
2 15 13
1 13
2 11 9
16 15 16 13 13 13 15 1 9 15 1 9 13 13 13 3 3
11 3 7 13 15 3 13 7 13 15 3 13
22 7 6 13 9 0 7 0 9 9 0 7 15 9 9 13 0 8 13 1 15 15 0
10 3 13 8 7 16 13 15 15 13 13
17 11 3 15 0 9 13 13 0 3 3 0 15 11 11 3 3 9
3 6 9 0
8 1 9 0 13 13 1 15 3
14 0 3 7 3 15 13 8 8 8 8 16 3 9 13
19 11 15 15 1 9 13 0 15 11 3 13 13 13 3 3 13 16 3 13
6 16 3 3 13 3 13
20 13 9 1 15 13 16 15 15 9 13 3 3 3 16 0 13 3 0 3 11
21 13 3 15 13 15 9 1 0 9 1 15 15 1 9 13 15 3 13 15 3 13
33 15 13 16 15 3 0 13 3 1 11 9 3 1 11 11 7 16 15 3 1 9 1 9 0 13 3 15 0 3 13 13 1 15
6 16 15 13 3 13 15
11 3 3 15 15 9 7 0 7 0 13 13
3 11 13 13
3 13 16 13
22 1 11 0 15 0 9 0 9 11 13 11 3 13 1 15 7 1 15 13 11 11 11
28 3 6 15 0 13 11 15 1 15 9 13 7 15 0 1 15 9 8 3 7 3 15 0 3 7 3 0 13
7 9 0 15 13 15 13 13
20 3 3 15 1 0 9 3 3 1 3 15 7 9 7 9 0 7 0 13 13
10 7 9 15 9 7 1 15 9 9 13
21 7 13 16 9 15 13 3 9 11 7 9 0 3 13 7 3 3 13 0 9 11
8 13 15 13 13 15 1 15 9
24 13 7 0 3 1 9 8 13 15 7 3 13 16 15 3 13 1 11 3 13 13 15 3 13
24 9 3 15 1 15 3 9 0 9 3 13 16 3 13 15 13 3 1 15 13 13 15 15 13
4 3 0 9 13
5 3 11 7 11 13
2 11 13
16 1 15 13 13 8 9 9 9 9 0 3 9 0 9 3 13
3 3 13 12
9 11 3 13 9 13 15 9 9 13
8 11 1 0 9 13 15 9 13
3 15 9 15
11 13 13 3 9 15 3 13 16 9 11 13
10 1 15 13 0 13 7 0 3 3 11
9 13 1 11 15 3 15 1 11 13
8 13 1 9 3 0 7 0 9
4 7 0 3 13
3 3 11 9
6 15 13 3 13 16 13
5 16 3 13 9 13
10 7 15 3 0 15 3 1 9 15 3
6 3 0 15 15 1 13
5 1 0 0 13 15
4 13 3 1 11
2 3 13
5 9 1 15 9 13
5 13 3 15 1 9
2 13 9
4 8 8 8 8
1 13
5 0 3 3 3 13
2 6 9
2 6 9
11 1 15 11 9 13 15 9 9 13 3 13
2 11 13
1 13
6 7 3 9 7 9 13
4 9 15 9 13
15 11 13 3 16 7 9 13 7 9 7 9 9 7 11 13
6 0 9 13 13 16 13
7 0 9 13 15 9 11 13
8 0 15 3 13 3 9 13 13
15 7 1 15 3 16 13 13 7 9 3 13 13 0 9 13
7 11 13 1 15 1 9 13
5 3 15 11 13 11
4 11 13 16 13
5 9 13 0 0 0
2 13 3
3 13 3 3
4 13 9 9 0
11 1 15 16 11 3 13 1 0 9 3 13
10 1 11 9 9 13 3 15 13 1 11
5 13 9 13 15 13
18 0 3 13 13 16 0 7 0 9 13 13 15 11 7 0 7 0 13
22 11 13 13 13 7 15 13 7 13 16 3 3 13 16 13 11 15 7 3 15 0 13
11 9 15 3 0 9 13 16 9 0 9 13
23 1 9 9 15 15 13 7 0 3 3 15 13 3 13 7 3 13 3 13 16 13 1 15
11 7 0 9 9 3 3 9 15 3 9 13
13 0 13 0 7 0 9 15 15 11 11 9 15 13
8 1 15 13 3 7 0 3 3
12 11 9 7 9 7 9 13 15 15 9 9 13
10 3 1 9 13 15 16 3 0 3 13
4 3 13 1 0
14 11 1 15 1 15 13 13 1 15 9 16 3 13 9
5 7 13 9 9 15
12 13 9 11 11 11 11 12 11 9 11 7 11
28 3 13 16 1 0 9 13 9 3 11 1 15 15 8 13 15 13 16 3 1 9 0 13 15 15 13 15 13
5 3 3 9 13 13
18 9 3 15 15 3 13 0 13 13 7 0 3 0 9 15 15 3 13
23 16 1 0 9 15 13 9 13 11 3 15 3 13 7 13 0 15 1 8 9 0 15 11
20 16 1 11 11 13 1 11 0 7 0 9 3 0 0 9 13 13 1 13 9
18 3 16 0 3 3 13 13 1 9 0 13 15 13 13 3 7 3 13
17 13 11 3 13 3 0 13 16 9 15 9 1 3 0 9 3 13
6 0 9 8 13 3 13
9 0 9 0 0 3 13 13 3 13
8 1 9 11 16 13 13 15 9
8 3 13 0 9 11 3 13 9
8 7 1 15 15 3 11 15 13
3 11 3 13
11 0 3 15 0 13 13 7 16 0 13 13
6 16 13 12 0 15 0
6 9 0 7 0 13 13
13 0 15 15 13 13 13 3 9 15 3 13 3 9
11 15 3 7 15 1 7 1 11 1 9 13
6 11 9 13 13 1 11
6 9 13 9 13 13 3
8 1 11 9 3 0 7 9 13
15 9 9 15 0 9 1 9 13 15 3 3 15 13 13 13
7 1 11 16 13 15 13 13
3 11 9 13
4 11 11 9 13
24 16 13 15 13 0 9 13 8 7 3 13 9 15 9 3 0 7 13 9 1 9 1 9 9
21 0 12 0 3 13 16 11 13 9 13 3 3 0 9 11 11 13 9 11 11 13
16 15 16 3 13 13 13 15 15 9 1 9 11 13 11 3 13
6 3 15 13 13 16 9
19 13 3 1 0 9 15 11 11 15 13 11 13 1 11 15 13 13 15 13
25 15 6 15 13 13 1 15 9 13 3 1 9 13 7 1 15 0 16 1 15 3 7 3 3 13
4 3 3 15 13
4 3 13 13 9
6 3 13 1 9 9 15
17 15 1 15 3 3 3 13 16 0 3 13 3 13 7 3 13 13
22 15 16 13 15 1 11 13 13 1 15 9 15 13 13 15 0 13 7 1 11 15 13
16 13 15 13 15 3 13 9 7 9 15 3 1 15 13 3 13
29 7 16 9 7 9 15 15 13 0 13 3 7 1 11 3 7 11 3 7 1 11 15 3 1 15 0 13 13 9
18 3 7 3 0 13 9 15 15 16 13 3 13 15 0 9 15 13 13
64 9 13 9 16 11 11 9 9 1 9 13 15 15 7 15 9 11 1 9 13 16 0 3 9 13 16 13 15 9 13 16 12 9 13 15 15 13 13 16 9 0 13 15 13 3 13 7 12 0 15 15 13 1 13 9 0 13 13 16 3 3 9 3 13
22 0 9 3 9 7 9 7 9 0 9 16 13 13 13 13 1 11 13 9 13 9 11
4 3 11 13 0
6 13 0 7 3 13 13
23 11 3 13 9 0 11 3 13 7 3 3 3 0 13 16 3 13 9 0 11 3 11 13
11 11 15 7 15 11 9 0 1 9 3 13
2 15 0
3 0 13 9
3 0 9 9
15 7 15 9 1 0 11 11 11 9 9 13 16 9 9 13
11 9 13 1 9 9 16 9 1 0 9 13
3 13 9 9
2 11 13
10 9 15 0 0 9 13 9 1 9 13
5 3 11 3 13 15
1 13
1 13
5 3 3 15 3 0
10 9 13 16 3 9 13 3 9 13 13
6 16 15 13 9 0 13
3 13 13 3
3 13 3 0
3 9 1 9
14 1 0 9 3 13 9 0 15 9 13 13 1 9 0
7 13 9 13 15 16 0 13
10 3 3 9 13 15 0 9 9 9 13
8 7 9 3 13 13 15 13 3
3 3 3 13
8 3 13 1 11 7 11 3 15
3 3 11 13
8 1 15 15 13 7 3 13 15
3 15 13 15
5 11 11 3 13 13
5 12 9 13 9 13
3 11 1 11
5 11 1 11 11 11
7 11 1 11 7 1 11 11
6 15 13 13 1 15 13
4 3 13 16 13
10 1 0 3 12 9 15 15 13 15 13
4 0 9 9 13
8 13 3 9 9 13 13 0 9
22 3 0 3 13 13 3 7 9 9 13 15 1 0 9 3 7 15 9 9 3 1 9
10 1 15 15 13 15 9 7 9 13 13
11 11 1 0 9 9 3 3 13 0 0 9
6 0 3 15 13 13 0
2 15 13
2 15 0
7 1 9 3 13 13 0 9
3 13 9 0
21 3 1 9 0 9 0 9 0 13 7 13 13 15 7 13 0 9 16 12 9 13
7 3 13 0 9 9 3 0
1 13
5 15 15 0 9 13
7 3 16 9 13 9 13 13
5 13 15 15 3 13
1 15
4 0 13 3 13
12 3 15 7 9 3 15 13 13 13 15 9 13
3 3 3 13
2 3 8
4 3 11 0 9
2 9 9
4 7 3 12 13
3 9 0 13
4 3 13 3 13
1 13
5 15 3 0 3 13
16 13 15 11 15 3 3 9 7 9 7 3 9 7 9 0 9
9 15 13 9 0 15 13 1 15 13
6 15 3 3 13 3 13
2 15 0
7 15 9 15 13 12 15 13
7 13 15 15 15 15 13 13
28 0 15 13 9 3 7 3 15 1 15 9 13 15 7 9 3 13 1 9 1 15 15 13 1 9 7 9 15
6 9 15 7 9 15 13
7 3 13 3 13 7 3 13
12 9 15 1 7 15 16 13 1 15 0 9 13
3 15 8 13
9 9 0 9 15 9 3 13 3 13
3 0 9 13
8 15 0 6 9 13 1 15 9
3 7 13 15
12 9 13 1 9 7 13 0 9 9 9 3 0
7 15 3 11 1 0 9 13
5 9 0 15 9 9
18 13 3 11 15 11 11 3 13 16 3 13 13 3 13 7 15 13 11
12 7 15 13 3 7 3 15 13 3 15 9 13
3 3 9 13
6 0 15 9 3 13 3
3 15 15 0
1 3
20 13 11 13 15 9 9 3 11 11 13 15 1 11 9 9 13 11 9 0 13
3 3 13 3
4 11 13 3 13
12 0 3 11 7 11 9 1 9 7 11 11 9
8 11 3 13 15 0 0 3 13
9 0 15 13 3 0 0 1 9 13
8 11 1 9 15 9 1 11 13
16 1 11 9 7 1 11 13 3 12 9 13 1 9 11 0 3
13 13 11 9 13 15 9 13 3 9 9 1 11 13
7 11 11 13 3 1 11 13
28 15 16 7 9 1 15 13 15 7 15 7 15 9 7 3 16 13 7 13 15 9 13 13 7 3 13 3 13
6 3 6 0 9 15 13
13 15 3 1 15 16 9 13 7 15 7 11 15 13
8 1 15 0 9 13 11 3 13
5 6 13 15 15 9
3 6 0 9
6 6 9 9 7 9 0
3 6 9 13
10 15 6 15 3 13 13 0 15 9 8
8 7 16 13 3 15 3 13 13
12 3 11 13 13 9 7 0 0 8 1 9 13
7 3 3 3 16 15 13 9
11 9 9 13 9 13 3 3 1 15 11 13
4 0 15 3 13
3 15 3 0
3 7 6 15
14 13 3 15 15 13 13 11 7 1 9 3 13 1 3
3 7 15 0
13 11 0 9 15 3 15 3 3 13 7 3 13 9
2 15 13
14 1 0 9 15 15 1 15 9 13 0 0 9 9 13
14 15 9 1 15 13 15 16 15 13 1 15 1 15 13
13 15 3 7 15 1 9 13 9 7 15 13 0 9
17 15 3 13 15 13 16 15 0 13 16 0 15 9 16 0 13 9
11 1 13 3 15 13 3 13 11 15 16 13
11 7 13 15 9 1 9 3 0 9 7 0
15 15 3 15 3 3 9 13 13 13 16 0 9 15 9 13
15 3 13 1 0 0 0 9 0 9 1 15 15 13 1 9
5 15 9 15 3 13
19 16 13 1 0 16 1 15 9 13 1 0 15 9 15 7 0 1 15 13
18 1 15 15 13 1 15 15 13 15 7 15 1 15 1 9 1 0 13
3 0 3 9
5 3 1 0 13 13
7 16 1 11 11 13 9 13
3 13 0 9
10 3 16 13 3 11 11 13 15 13 9
3 15 9 13
17 15 13 15 3 3 13 13 0 0 7 3 9 3 3 9 7 9
13 15 3 1 15 3 13 16 13 11 16 9 15 13
9 3 11 6 13 15 0 15 13 3
1 13
4 15 13 3 13
4 3 15 0 13
8 3 3 7 3 9 9 7 13
2 13 13
6 15 3 11 1 9 13
2 0 13
2 15 0
11 15 15 9 0 15 0 15 9 15 13 13
12 7 0 13 15 3 15 0 9 3 0 11 13
31 11 1 11 13 7 11 1 15 3 3 13 15 7 13 3 7 15 1 0 13 13 7 16 13 13 13 0 9 15 15 13
2 15 13
18 0 1 15 13 3 0 3 3 13 16 13 15 3 13 9 13 7 13
33 0 13 16 16 13 9 15 13 13 1 15 15 11 13 16 13 13 13 16 13 3 13 15 6 15 15 3 7 0 13 3 7 0
7 11 11 3 13 11 0 9
10 15 15 1 15 13 15 1 9 13 13
16 3 16 0 13 9 1 0 13 16 0 9 13 1 0 1 11
8 3 13 1 15 9 0 9 13
18 15 13 15 9 0 3 13 0 3 16 13 15 13 1 15 13 15 9
14 13 1 0 9 3 11 15 15 1 9 9 9 13 13
6 13 1 11 3 0 11
5 3 1 15 3 13
2 3 3
17 16 11 13 7 0 7 3 3 7 11 16 0 3 9 0 3 13
2 3 13
4 3 13 3 9
7 1 15 0 13 15 13 13
13 3 3 13 13 16 15 13 1 15 9 3 13 13
16 0 9 3 0 15 13 7 3 1 15 15 13 16 13 3 13
4 7 13 1 0
16 13 13 15 15 9 13 0 0 9 3 16 13 3 0 0 13
10 0 15 3 13 0 3 13 1 9 15
16 15 15 13 15 9 13 3 3 3 15 13 13 16 1 11 13
12 1 9 0 13 1 15 13 16 15 13 15 13
7 15 16 3 13 0 9 13
5 7 15 1 11 13
6 3 13 1 0 1 11
11 3 15 15 9 0 13 13 0 1 15 9
10 3 3 13 1 0 11 13 1 15 9
7 3 3 3 13 3 15 13
6 15 1 9 0 9 13
1 13
7 1 15 9 15 13 13 13
13 0 3 3 13 1 15 15 0 3 1 0 13 13
6 15 0 9 11 11 13
4 13 3 3 13
5 0 13 1 15 0
14 3 13 16 15 13 8 1 15 15 3 13 15 13 13
6 1 11 13 15 1 9
6 11 15 9 15 13 0
3 11 13 3
5 1 11 1 0 3
11 3 13 0 9 15 15 0 9 13 15 13
11 1 15 15 0 0 9 13 1 0 1 11
16 7 0 3 15 11 13 15 0 11 3 3 15 13 0 9 11
12 0 13 15 15 9 1 0 15 0 7 0 9
6 7 9 13 15 0 13
20 1 0 0 15 13 15 13 13 3 0 13 13 16 15 13 7 15 13 8 13
3 13 15 9
12 3 13 15 16 15 15 13 13 11 11 13 0
10 3 16 3 9 13 13 3 9 3 13
9 3 13 1 0 9 15 13 1 11
4 1 11 13 3
5 16 3 9 3 13
6 15 3 13 13 3 11
14 7 3 13 16 9 9 0 13 1 15 3 13 9 9
6 1 11 7 11 16 13
11 1 0 15 11 16 3 3 8 13 6 9
6 3 3 0 15 13 13
9 3 1 0 7 3 3 16 1 11
18 15 1 11 13 0 15 13 3 16 0 9 1 15 13 3 1 15 13
2 7 13
3 9 3 13
19 1 15 9 15 13 1 12 9 15 11 13 13 16 1 15 13 13 16 13
4 0 15 9 13
3 13 1 15
6 3 3 13 9 15 13
4 15 3 13 12
9 3 15 1 15 9 0 9 9 13
13 3 9 7 9 7 3 16 15 0 13 1 11 13
10 9 7 15 7 11 1 15 9 3 13
4 3 13 15 13
4 3 15 0 13
10 3 3 13 3 15 11 3 13 0 13
14 13 3 15 15 9 15 3 3 9 15 7 3 9 13
3 15 13 11
12 3 3 11 1 0 9 15 15 13 13 9 13
13 15 11 15 1 11 8 1 9 0 13 1 15 13
31 3 15 0 13 13 15 1 9 3 1 15 13 13 15 13 3 3 11 13 13 16 7 3 13 3 9 13 7 16 13 3
8 7 16 13 3 13 13 0 3
3 11 13 3
3 15 13 3
9 0 3 15 0 1 9 0 9 13
8 13 3 9 0 1 0 15 9
16 7 1 15 0 3 1 13 13 13 13 11 3 13 7 3 13
19 15 3 3 13 13 15 3 3 13 16 15 16 13 13 1 15 9 3 13
10 3 3 3 13 15 7 13 15 7 13
2 13 15
15 0 3 3 13 16 13 15 13 1 11 9 13 16 13 13
11 3 13 15 9 7 3 16 13 9 9 15
11 3 7 3 1 9 0 0 9 1 15 13
9 3 3 3 13 15 1 11 3 13
20 7 3 16 9 13 15 13 15 1 3 13 15 11 0 9 13 0 9 0 9
12 15 16 9 1 11 7 1 11 13 13 11 3
11 9 0 0 13 7 1 0 15 13 13 0
28 15 7 0 9 1 15 3 13 3 16 1 9 13 7 11 9 1 15 3 3 9 3 13 13 0 3 9 11
14 15 16 3 13 11 3 3 13 16 13 0 3 13 13
17 11 13 9 11 15 13 1 9 9 15 16 11 9 13 1 9 15
21 0 15 3 13 13 1 11 11 9 15 7 0 11 13 3 0 9 15 15 13 13
36 15 3 9 15 7 0 13 3 16 1 9 15 13 9 16 0 0 9 0 9 15 0 15 1 13 13 3 16 11 15 13 0 13 13 13 13
13 13 3 0 16 0 15 16 15 13 13 3 3 13
5 3 9 0 13 13
5 15 3 13 3 0
27 16 0 13 16 13 1 9 16 0 11 13 11 3 15 15 3 13 15 7 0 13 3 13 0 11 1 9
3 13 1 11
17 13 3 1 11 1 11 1 11 3 7 3 16 3 13 11 15 13
3 9 13 0
9 13 3 1 9 9 9 7 15 13
28 11 13 3 16 3 7 11 7 11 9 15 15 7 11 7 15 9 11 3 7 8 15 13 13 13 0 1 9
13 11 13 9 13 9 15 3 13 7 11 13 0 13
12 9 3 0 11 13 1 9 3 3 13 13 0
7 9 13 13 7 9 15 13
22 15 13 15 13 3 15 9 13 13 15 9 15 11 13 3 1 3 7 3 13 16 13
11 15 0 3 9 13 15 1 15 3 13 13
38 0 3 16 3 13 16 0 3 13 13 3 1 9 3 15 13 13 13 1 15 7 1 15 15 1 0 1 11 16 9 15 13 15 9 16 15 0 13
14 0 15 3 13 16 13 3 3 15 13 16 13 16 13
7 7 3 13 15 15 9 13
4 9 3 3 13
23 11 3 3 3 13 13 7 3 0 13 7 6 1 0 16 15 13 3 7 15 9 13 13
18 16 11 3 13 13 3 3 0 9 11 3 7 1 15 9 0 15 13
8 3 6 15 15 9 3 1 15
9 7 15 1 15 0 15 13 3 13
2 0 13
15 3 9 3 7 1 15 7 3 7 3 3 7 1 15 9
7 15 13 9 0 15 1 9
2 3 3
8 0 13 9 9 7 0 9 13
11 15 13 13 1 0 1 15 3 15 13 13
17 0 13 0 9 16 15 9 3 13 16 3 15 9 1 0 9 13
6 6 9 3 0 15 9
5 6 0 0 8 8
1 13
5 3 3 1 9 13
6 3 13 7 13 0 13
15 3 0 0 13 3 9 3 13 7 9 3 7 13 0 9
18 3 0 7 3 7 3 7 1 15 9 3 3 3 7 13 7 13 3
7 3 13 15 8 16 0 13
6 0 15 8 0 9 13
4 3 0 3 3
18 3 6 3 3 3 0 9 15 13 15 1 11 15 1 11 9 13 13
17 7 3 3 15 9 7 3 11 3 15 16 13 1 9 0 15 13
24 3 16 15 13 15 13 1 0 9 15 13 13 15 13 3 15 0 13 16 15 13 1 15 13
3 15 13 3
4 15 3 3 0
16 3 11 15 7 15 3 11 13 7 3 1 9 0 9 3 13
22 15 13 16 3 13 15 9 1 15 13 16 13 15 13 3 15 9 3 3 11 13 13
15 3 3 3 3 3 13 3 16 3 13 13 13 16 3 13
12 16 9 15 13 1 9 16 13 15 13 13 13
13 3 13 13 3 13 9 9 3 3 0 9 9 13
4 11 3 1 0
8 16 0 9 3 13 13 3 0
10 3 15 13 3 0 9 15 3 11 13
12 11 15 3 13 15 13 11 13 1 11 3 13
12 15 3 11 3 13 15 13 0 3 0 3 13
3 3 0 13
7 13 3 9 15 1 0 3
12 15 0 3 13 11 13 16 3 12 0 13 9
5 13 0 3 11 11
2 13 9
4 15 0 11 13
4 15 13 9 13
18 15 3 9 1 11 0 1 9 13 3 7 6 13 15 3 15 13 15
9 13 15 13 15 9 7 9 9 15
4 3 13 9 15
11 15 13 16 0 0 13 8 8 8 3 13
12 15 3 1 15 13 3 13 16 15 13 13 9
9 16 15 3 13 13 15 1 15 0
10 3 3 9 0 13 7 3 13 13 0
9 3 13 16 16 15 13 13 0 13
6 3 13 1 15 15 13
8 3 13 3 8 3 1 11 13
5 11 3 13 3 15
5 15 0 13 3 13
15 1 11 7 0 9 15 1 0 9 13 7 6 9 15 13
20 3 15 11 13 15 13 1 15 15 1 0 9 9 0 9 13 15 15 0 13
49 7 16 11 15 1 13 16 13 1 15 11 8 13 15 11 9 13 0 13 13 7 11 7 3 0 11 15 1 11 13 15 3 3 15 11 13 11 13 13 16 15 1 15 13 13 15 15 9 13
5 3 13 1 15 3
6 15 9 13 1 15 9
6 15 13 11 15 9 13
3 13 3 15
4 15 0 15 13
7 13 9 1 15 13 9 11
1 13
1 13
17 11 15 15 9 13 13 1 15 3 3 13 3 15 15 3 3 13
8 13 16 15 13 7 3 16 13
8 9 0 13 13 7 0 9 0
5 0 9 11 11 13
12 3 1 11 1 11 9 0 15 15 3 11 13
4 3 1 11 3
2 3 11
2 3 11
4 3 13 9 0
6 15 15 0 9 13 13
17 3 13 1 9 15 13 3 7 15 11 13 16 15 8 8 0 13
23 1 11 1 15 3 3 13 1 11 13 9 7 15 15 9 15 3 1 11 15 3 3 8
50 7 15 1 0 9 9 7 6 0 1 9 0 9 9 13 8 3 13 16 15 1 11 15 13 9 0 9 13 9 1 15 15 3 15 13 3 0 3 11 9 0 13 13 9 15 7 15 13 13 13
10 15 13 13 1 11 1 11 1 0 9
9 15 3 9 16 11 13 13 15 13
22 15 9 13 15 13 1 9 9 3 13 1 9 16 15 13 13 0 13 9 15 13 13
4 3 15 15 13
13 3 16 15 11 13 15 1 15 9 13 0 13 13
6 0 13 1 15 16 13
6 3 13 3 1 0 9
12 13 1 9 7 1 9 7 3 1 9 0 9
28 1 9 9 9 7 1 0 9 15 15 3 11 7 0 1 9 11 3 13 7 13 15 13 7 15 1 15 13
15 1 15 15 13 3 13 0 9 9 15 3 1 9 13 13
23 7 3 13 13 0 9 15 1 15 13 0 7 13 7 3 3 16 1 15 9 13 13 9
22 15 9 11 9 15 13 11 7 16 1 9 15 3 13 13 15 0 3 11 7 11 13
3 0 11 13
5 3 15 15 13 13
4 3 0 3 3
3 13 1 0
17 1 9 16 11 13 3 0 13 7 13 13 16 13 0 16 13 3
16 3 13 15 9 3 7 16 15 13 1 0 0 9 15 3 13
13 3 1 11 15 1 9 15 9 13 3 7 15 13
16 16 15 9 13 3 7 0 1 15 3 7 3 15 9 9 13
6 16 3 13 9 15 13
3 13 11 3
3 0 13 11
7 1 9 15 13 15 13 3
9 1 0 9 16 15 13 8 8 13
27 3 3 0 15 15 13 13 3 9 0 3 13 9 9 3 9 9 13 1 11 9 7 15 3 1 3 13
4 15 11 13 3
6 13 15 15 13 9 15
7 15 3 15 1 11 15 13
17 13 15 1 9 0 13 1 9 0 9 0 9 0 13 0 9 9
21 15 13 16 15 3 13 0 1 9 0 3 15 13 1 15 15 15 13 15 13 13
26 15 15 0 13 13 16 3 15 13 15 0 16 15 15 13 13 3 7 0 8 15 15 13 15 13 0
6 13 9 0 9 7 9
3 0 0 13
3 11 13 3
2 15 0
24 7 13 0 3 15 9 13 3 13 3 0 9 0 15 3 0 9 9 7 9 15 0 9 13
23 3 9 11 15 13 16 11 11 11 13 7 16 9 15 9 13 0 15 9 13 12 9 0
4 3 0 3 13
6 9 9 9 9 15 13
7 7 13 3 13 13 16 9
4 16 13 13 13
8 3 3 13 13 15 16 11 13
6 3 13 16 0 9 13
4 3 13 0 9
17 0 9 1 9 15 16 13 16 0 15 15 1 13 9 15 13 13
10 11 9 3 13 7 13 3 7 13 13
12 9 11 13 3 16 0 9 13 1 9 1 11
15 3 1 11 13 16 1 11 9 13 16 13 1 9 15 13
4 9 9 13 13
5 3 3 13 15 9
16 3 3 1 15 3 13 3 0 3 9 0 13 16 15 13 13
14 15 3 3 13 9 9 13 1 9 9 7 9 15 9
24 16 1 0 9 7 9 13 9 9 7 13 1 9 3 13 15 13 9 16 15 0 9 15 13
14 3 13 1 0 9 16 0 15 0 13 9 3 15 13
22 0 9 1 0 7 3 0 1 0 9 15 13 13 3 13 9 11 9 11 3 9 11
24 13 15 15 3 13 8 13 3 13 8 15 13 9 9 9 9 15 3 9 7 9 13 15 0
2 15 13
22 13 3 0 9 16 15 13 9 1 15 3 7 1 9 3 7 1 9 3 7 1 15
13 3 0 1 9 9 13 1 9 1 9 1 9 15
5 6 3 9 15 13
9 9 9 9 15 11 3 9 15 13
12 11 16 13 15 13 1 0 9 15 13 11 3
3 3 9 13
15 1 9 9 13 7 3 13 9 15 1 9 13 15 15 13
11 15 3 13 1 0 9 13 16 3 13 13
7 15 1 9 13 15 13 9
14 1 15 16 3 13 7 11 13 11 13 13 9 3 15
14 3 9 13 13 1 9 16 1 9 13 1 15 13 9
8 0 9 13 0 9 15 13 9
4 3 3 15 13
24 15 3 16 0 15 1 15 13 13 3 1 9 15 13 15 1 9 13 16 15 9 13 1 15
6 3 15 3 8 9 15
4 11 15 0 13
3 7 3 13
14 11 15 11 9 15 9 1 9 13 13 15 1 1 9
11 16 1 9 15 13 0 9 9 13 0 13
20 11 1 15 13 15 15 1 13 1 15 0 7 0 9 13 7 15 15 13 13
16 13 15 13 1 0 9 7 1 15 13 15 7 13 7 15 13
10 15 1 11 3 15 16 0 13 13 13
7 16 15 15 13 0 9 13
8 13 3 13 3 0 1 15 13
23 7 3 0 9 9 7 9 13 0 13 16 3 13 15 15 11 13 15 0 12 9 11 13
8 3 9 13 16 15 13 1 9
5 15 15 9 3 13
11 3 3 13 9 1 13 9 15 13 13 9
17 7 0 11 15 13 13 0 13 3 3 15 9 15 3 3 13 13
8 3 13 11 13 16 3 3 13
21 15 3 0 13 3 13 15 15 9 3 13 1 15 13 13 15 1 11 13 1 3
22 7 16 7 11 13 16 7 1 11 9 11 13 9 11 11 9 9 9 1 0 3 9
6 11 3 13 13 1 11
6 0 1 9 13 1 9
28 15 9 16 11 13 13 13 3 13 7 0 3 15 15 8 16 15 1 13 7 13 3 13 9 15 13 7 9
22 15 16 13 3 7 0 3 1 15 9 13 12 13 16 9 1 0 9 9 11 13 13
14 3 16 15 1 9 13 3 13 15 16 9 3 15 13
5 0 3 16 13 11
11 16 13 7 3 16 13 0 9 3 15 13
12 13 9 7 16 9 3 13 0 13 13 3 9
22 3 13 0 1 9 11 3 13 0 1 13 9 0 9 7 3 13 1 9 1 15 13
16 9 3 0 13 3 15 13 13 15 0 13 15 7 9 7 9
7 9 1 9 1 9 0 13
4 3 0 9 13
12 13 3 15 7 16 3 13 3 13 8 9 15
22 7 15 13 16 15 9 13 13 16 0 1 9 15 9 1 3 13 16 11 13 9 0
7 3 15 13 9 16 15 13
7 0 9 13 15 9 9 11
7 3 15 13 9 9 9 9
11 11 15 13 1 11 7 16 9 13 13 11
7 15 16 13 11 3 13 3
28 16 1 11 13 3 1 15 1 15 15 9 16 7 15 15 15 13 7 15 15 15 13 15 7 13 13 13 13
11 15 15 11 9 3 13 16 15 0 3 13
7 7 3 13 9 3 7 13
7 13 3 9 7 0 7 0
10 13 3 3 15 3 15 0 13 3 0
4 7 3 13 15
33 1 15 3 13 16 15 11 13 16 11 13 7 3 1 11 13 13 3 7 13 3 13 16 1 11 0 13 3 3 3 15 3 13
9 1 0 9 13 1 11 16 13 11
13 9 15 9 1 15 13 13 3 7 13 16 0 13
21 9 15 15 3 11 0 13 13 15 7 15 3 13 3 7 13 7 0 13 3 13
4 3 7 3 13
16 1 11 7 15 9 15 1 9 1 11 13 0 15 0 13 13
17 16 13 0 15 9 13 15 15 1 9 15 9 9 13 0 9 9
6 3 15 3 13 16 13
1 13
2 3 13
9 7 3 13 16 8 8 13 8 8
12 9 3 15 15 9 13 0 9 16 13 15 13
4 0 9 15 13
1 13
3 9 13 3
7 3 13 11 11 7 11 13
4 15 13 8 8
6 3 3 13 15 0 9
18 11 16 13 13 15 3 15 13 13 0 9 9 15 15 15 3 13 3
11 3 1 9 0 15 13 3 13 11 3 13
12 3 13 9 0 13 0 7 9 15 9 13 0
17 15 0 11 3 11 12 9 13 7 11 9 11 12 9 11 12 13
2 15 0
2 15 0
5 3 9 13 1 11
31 1 0 9 16 0 1 9 9 13 13 1 11 1 11 9 0 15 11 13 0 9 16 0 11 7 0 9 11 15 13 13
21 16 9 12 1 11 11 9 13 0 13 13 9 1 0 9 11 3 13 11 3 13
9 3 3 9 1 11 13 1 11 9
3 11 13 3
6 15 9 13 9 0 0
6 3 3 0 9 9 13
8 9 0 0 11 9 15 0 13
3 9 13 13
22 9 0 9 13 0 0 15 1 11 13 1 11 11 9 3 3 0 3 7 15 7 15
10 3 9 12 13 13 7 13 11 3 13
27 3 13 3 13 15 8 13 3 8 8 8 8 9 9 15 7 11 15 11 13 9 13 7 9 9 13 13
16 15 1 9 0 9 11 9 9 9 13 15 7 13 0 3 9
7 13 1 11 15 9 1 9
3 13 3 11
8 13 13 9 0 0 15 13 0
32 3 0 9 0 0 13 9 7 0 9 0 15 9 11 11 7 0 9 0 7 11 11 11 11 11 0 7 0 9 9 9 9
8 3 9 0 13 3 9 3 9
12 15 1 11 15 9 0 9 15 9 1 9 13
20 9 0 9 9 0 0 9 9 0 9 0 9 9 0 0 15 0 9 9 13
11 0 3 11 9 3 15 9 13 0 9 13
3 9 13 3
9 16 0 13 1 9 9 13 1 3
11 3 9 1 9 9 3 13 13 11 9 13
2 0 3
4 7 1 0 13
12 3 7 3 15 0 9 13 15 9 9 13 13
26 15 1 9 15 15 3 9 0 13 13 15 13 0 9 3 7 15 3 9 15 0 13 3 9 0 13
2 15 13
2 13 0
14 15 15 3 13 3 7 3 13 15 1 0 9 13 13
2 3 8
3 3 0 8
19 8 8 9 7 9 7 16 9 15 8 15 3 3 8 13 9 9 7 13
6 3 1 11 3 9 3
5 11 13 3 13 13
6 15 3 3 13 3 15
4 3 13 3 15
13 7 3 13 0 9 9 15 9 9 1 9 15 13
2 13 15
5 3 15 11 3 13
9 7 13 0 1 15 15 3 13 13
12 13 3 16 16 1 9 13 16 11 13 15 13
6 0 15 16 13 15 13
14 13 1 0 15 15 3 13 1 15 0 9 3 3 13
13 15 3 11 9 15 13 0 7 3 3 0 9 13
8 3 15 11 9 13 13 3 13
11 0 1 11 7 15 9 13 7 15 15 13
9 9 0 16 11 13 13 3 3 13
14 11 1 11 11 3 3 0 13 7 15 13 13 13 13
12 15 16 11 13 11 9 15 9 9 0 13 13
3 15 13 3
15 11 15 9 0 13 13 1 15 3 13 1 11 11 13 13
15 15 3 0 13 9 16 13 9 3 3 9 0 3 9 15
9 11 1 9 13 7 1 15 3 13
23 15 3 13 11 1 9 0 13 16 7 3 13 7 0 1 15 0 1 15 7 1 15 13
3 7 0 3
9 13 16 13 7 16 13 3 13 11
4 3 7 3 13
19 15 15 7 11 7 0 11 3 13 7 3 1 9 0 7 13 13 0 15
25 15 13 15 3 1 15 13 1 9 11 13 9 16 15 15 15 7 9 9 13 13 16 15 9 13
4 15 15 0 13
4 3 15 13 0
8 3 13 11 15 9 0 3 13
8 13 15 3 3 13 7 3 13
33 11 11 9 11 11 9 15 0 0 9 13 1 15 15 1 15 13 15 15 13 3 0 15 3 13 15 1 15 13 13 13 0 9
12 13 0 3 1 11 1 11 9 7 15 15 8
9 3 3 13 1 11 0 7 9 13
34 3 7 11 9 9 9 1 9 15 13 3 7 13 11 15 9 13 13 11 9 1 15 13 13 16 1 15 9 0 0 9 11 13 13
16 15 3 9 0 9 0 1 9 13 13 13 3 0 15 9 13
3 0 13 13
4 11 3 13 13
44 1 0 9 0 13 16 16 11 1 9 9 0 3 13 11 15 9 1 9 13 16 0 9 13 3 13 9 15 16 13 13 13 13 3 7 1 0 9 9 0 9 0 9 13
25 3 16 15 15 13 15 3 9 3 13 13 13 7 3 3 16 15 13 15 9 9 9 0 9 13
7 7 13 15 0 15 9 13
8 13 16 13 3 13 7 15 13
24 16 0 8 13 0 15 9 15 13 13 11 15 3 13 7 13 15 1 13 13 9 13 3 13
12 13 3 3 3 11 1 9 9 1 11 9 13
4 1 0 8 0
5 13 9 15 15 13
4 13 15 9 15
6 3 3 13 15 13 9
11 3 15 11 9 9 0 13 15 13 3 13
8 11 9 15 13 3 1 15 13
11 11 15 9 7 3 9 7 0 9 9 13
11 0 9 0 0 13 12 0 0 1 0 9
10 3 15 13 16 13 11 11 15 3 13
10 7 3 15 15 0 3 13 1 0 13
33 13 13 15 9 3 3 13 13 3 15 9 15 13 9 9 13 13 3 7 1 9 0 3 7 1 15 15 1 3 1 11 11 9
32 15 3 13 7 0 9 13 3 3 1 9 3 3 15 13 15 9 1 15 3 15 13 13 16 15 13 13 16 9 13 9 13
4 1 15 13 15
9 15 9 13 11 9 9 7 11 13
30 11 11 15 11 9 0 9 7 3 3 13 13 1 11 16 3 0 9 13 16 9 0 0 15 3 13 9 15 13 13
7 3 13 1 9 0 3 13
18 0 1 11 13 13 11 3 3 6 13 13 15 9 11 9 3 7 0
23 3 3 3 11 13 13 0 9 11 15 9 15 12 9 9 15 15 15 13 9 3 9 13
10 9 0 16 1 9 9 13 0 9 13
4 0 9 0 12
13 1 0 9 15 0 13 15 9 15 3 9 13 13
13 9 9 8 13 3 7 13 1 15 9 0 0 9
8 7 3 15 15 0 13 1 15
4 13 16 15 13
6 15 3 15 0 13 13
27 9 3 3 1 11 13 16 3 9 15 15 0 13 15 3 13 1 0 15 11 9 3 15 13 15 13 13
13 3 15 9 0 9 13 9 13 13 11 0 7 0
8 1 3 1 11 16 3 0 13
4 13 3 1 9
12 0 16 13 3 13 1 9 13 1 9 13 13
10 13 3 1 9 11 11 7 11 9 3
5 3 15 13 13 3
9 3 13 1 11 9 16 15 13 13
7 15 3 0 7 15 0 13
3 13 9 15
4 3 13 1 11
14 9 13 11 15 15 9 9 1 11 11 11 7 11 11
6 15 15 0 1 9 13
3 11 3 13
6 11 1 15 1 9 13
11 13 13 13 15 11 9 16 15 9 9 13
2 13 9
5 13 15 15 13 13
4 15 0 15 13
6 11 11 13 13 9 15
9 15 13 11 1 11 11 15 0 15
10 16 9 13 13 9 9 15 13 16 13
2 9 13
1 13
16 11 15 9 15 9 13 0 11 1 15 9 13 7 0 13 9
3 3 13 11
2 15 0
19 16 15 9 15 13 16 1 15 9 11 13 7 1 15 11 13 16 9 13
6 0 1 9 1 11 9
3 13 15 13
2 13 13
10 13 3 1 15 1 9 9 16 9 13
13 9 3 3 3 13 7 3 0 13 15 1 15 13
2 13 9
6 3 13 11 7 13 9
18 3 16 15 1 9 0 0 15 13 13 1 9 0 0 1 9 13 0
2 15 13
1 13
18 3 0 13 9 9 11 11 7 9 16 15 11 13 9 1 0 9 13
4 3 13 9 9
9 13 12 9 9 0 9 1 0 9
15 3 15 11 9 0 9 11 13 13 0 16 15 9 9 13
16 13 9 11 9 9 16 3 7 9 3 7 15 15 13 9 13
2 9 13
20 3 3 13 1 9 9 15 15 13 0 9 9 16 1 9 9 13 9 0 13
22 3 13 9 9 16 1 0 9 9 13 3 16 15 9 15 9 13 3 0 7 16 0
21 13 15 15 3 13 7 0 13 9 12 15 13 0 15 13 13 13 3 0 3 0
6 13 16 15 1 12 13
1 3
6 13 0 1 15 13 11
1 15
4 15 15 13 13
3 13 12 12
2 9 13
1 15
5 9 13 13 9 13
1 13
3 1 9 13
4 0 15 13 13
3 13 16 13
5 13 16 9 3 13
5 13 9 9 3 13
9 0 13 16 1 9 13 13 3 13
4 13 15 15 13
11 15 15 0 11 15 0 1 9 0 3 13
7 15 3 0 3 3 0 13
14 3 7 0 9 0 0 3 13 7 3 0 0 0 13
9 15 16 11 3 13 13 3 0 13
25 7 9 15 3 13 3 16 9 9 3 13 13 13 16 15 13 13 1 9 9 16 0 0 9 13
10 0 15 13 16 15 9 13 3 13 13
27 1 15 3 8 8 11 11 11 9 13 1 15 1 9 0 13 9 16 9 9 0 9 9 1 9 0 13
10 13 15 3 9 11 11 13 16 9 13
4 3 9 0 3
22 13 1 11 9 15 16 0 9 13 1 15 15 3 13 13 3 16 0 9 7 9 13
11 1 8 13 0 15 15 11 9 16 11 13
3 7 13 13
7 1 11 9 0 9 15 13
10 3 11 1 9 1 9 0 13 3 13
6 11 3 13 0 9 13
13 11 11 13 13 15 11 9 15 7 13 1 15 13
12 9 15 3 3 13 3 16 11 13 7 3 13
18 15 3 13 3 8 8 3 3 13 3 7 8 15 13 7 9 13 15
17 0 1 11 15 15 9 13 13 3 13 7 13 13 15 15 15 13
15 15 3 15 13 1 0 15 13 11 9 7 11 7 11 13
17 3 3 8 0 9 15 13 7 3 13 16 3 0 13 16 15 13
6 3 15 9 13 13 3
13 16 15 8 1 11 15 9 3 1 11 13 3 13
4 7 13 3 3
18 11 3 1 15 1 9 3 3 7 8 9 13 16 15 1 15 13 13
7 3 3 9 15 9 13 9
28 15 3 13 13 3 0 3 0 13 13 13 9 7 9 9 15 15 13 9 15 13 13 3 7 3 3 7 3
8 15 13 1 0 9 9 9 3
6 1 9 1 9 1 9
19 3 3 9 6 15 0 9 7 0 9 13 7 3 0 13 3 15 0 9
27 0 0 9 11 3 13 15 15 3 13 3 13 13 16 0 3 13 7 3 13 3 15 9 7 0 9 9
34 16 11 3 11 9 15 1 15 13 13 9 15 13 3 3 13 7 3 0 0 9 15 0 1 9 13 13 15 0 3 13 7 13 13
23 3 13 1 11 15 15 15 9 15 9 13 13 15 3 13 13 7 3 15 13 16 15 13
4 15 13 3 13
12 3 1 11 3 13 16 9 15 15 13 0 13
9 3 15 1 9 13 0 9 9 13
8 3 1 11 9 12 13 13 13
20 11 3 3 1 0 9 3 13 12 3 0 15 3 16 13 1 9 0 13 13
5 15 3 3 3 13
10 0 15 9 9 0 12 7 0 1 9
2 9 13
6 15 3 9 15 9 13
4 11 9 9 13
9 15 3 1 9 11 15 3 13 13
17 9 9 12 12 7 0 13 7 15 15 3 3 13 3 15 7 15
10 3 3 13 3 1 9 13 13 13 9
12 11 3 15 13 15 1 15 9 13 1 9 11
12 7 6 15 3 13 15 0 9 0 15 9 0
15 3 7 9 13 15 13 7 3 1 11 11 9 7 9 13
7 3 7 3 1 9 15 13
14 15 3 13 15 3 13 16 3 13 9 13 16 3 9
5 3 12 15 3 13
7 7 15 15 13 1 9 13
12 3 13 1 9 15 13 15 3 0 13 3 15
18 3 3 9 15 13 1 15 13 9 9 13 11 11 7 11 11 9 15
3 15 15 13
12 13 3 7 3 9 13 13 15 1 0 0 9
4 3 11 0 13
9 13 16 13 16 15 0 15 3 13
21 3 1 9 15 13 7 9 1 11 7 1 0 11 9 13 15 7 9 13 3 13
29 7 0 9 0 13 15 9 11 11 9 0 15 9 13 15 3 7 15 3 11 13 3 7 15 3 16 9 11 13
6 3 16 15 0 3 3
21 13 3 9 11 7 3 13 9 9 15 13 1 9 9 11 13 16 9 9 12 13
21 3 15 15 9 13 9 16 15 0 9 11 3 13 9 13 16 9 1 9 3 13
12 0 1 9 13 11 0 1 15 15 1 11 13
16 0 3 13 11 15 9 13 15 15 9 1 9 15 13 9 13
9 13 3 0 15 13 15 0 16 13
8 13 9 13 15 13 1 9 15
5 13 1 9 16 13
13 9 0 3 15 13 7 15 15 13 16 3 11 13
5 7 0 0 11 13
8 15 1 15 1 15 0 9 13
12 1 15 3 3 16 13 15 3 3 8 13 13
4 13 3 15 0
38 3 0 0 9 3 1 15 13 7 3 15 13 13 15 3 13 0 15 15 1 15 15 9 13 16 15 15 1 0 9 3 0 9 13 15 0 3 13
7 3 15 9 13 9 11 13
6 3 15 0 13 15 13
5 3 1 11 3 13
13 7 13 15 13 8 0 15 13 15 15 1 9 13
5 13 15 15 9 13
10 15 9 15 13 1 15 3 15 9 13
1 13
10 1 15 12 8 13 1 11 11 11 9
19 0 3 1 9 3 13 3 15 9 0 13 15 9 0 9 3 9 13 13
6 15 3 13 16 13 9
12 13 13 15 9 0 9 16 9 13 13 1 0
24 3 3 0 13 9 11 11 9 9 13 9 7 13 16 15 0 7 3 11 15 3 13 13 13
7 8 8 8 0 1 9 9
3 15 3 13
13 15 1 9 1 9 13 1 0 9 13 11 3 9
14 1 11 15 15 13 13 7 1 15 7 1 11 15 13
7 15 3 1 15 3 3 13
8 7 13 15 1 15 0 9 13
7 13 3 9 0 15 9 13
10 3 3 13 0 1 11 3 0 1 11
24 3 13 11 15 9 3 0 15 3 13 3 3 16 13 3 9 11 9 1 15 1 0 9 13
10 15 13 15 15 13 3 3 3 1 11
5 11 9 15 3 13
12 3 3 15 15 15 9 13 3 15 0 0 13
10 7 13 1 15 1 0 0 16 11 13
9 1 11 15 9 15 9 13 3 13
8 3 9 13 13 7 13 0 13
8 7 3 8 16 0 13 15 13
4 15 3 13 8
5 11 9 13 1 15
6 11 9 0 9 13 13
3 13 3 9
7 15 3 13 16 13 3 13
6 11 15 3 1 9 13
6 9 3 13 15 3 13
16 7 9 3 7 0 3 7 0 13 13 3 7 15 15 7 0
5 11 11 3 13 13
7 13 11 11 11 15 16 13
4 13 3 13 9
4 0 13 8 11
7 11 16 9 15 13 3 0
7 1 11 9 15 13 13 11
4 11 15 9 13
3 11 3 13
10 0 3 13 3 3 11 15 1 13 13
3 0 9 13
10 1 0 9 7 0 9 9 15 13 13
7 15 15 1 9 0 13 13
4 8 11 13 13
6 13 16 15 0 0 13
3 0 9 13
4 3 11 13 13
8 15 13 13 13 16 3 13 9
6 3 13 1 0 9 9
1 13
5 12 3 9 13 11
8 15 0 13 15 13 3 16 9
8 15 15 3 16 3 3 3 13
15 15 3 1 11 13 16 0 1 15 9 13 1 15 9 15
9 13 3 9 0 15 9 12 9 12
6 13 1 13 3 11 13
11 15 9 15 1 15 13 13 15 9 0 13
3 13 0 11
2 15 13
3 0 13 9
6 3 0 9 1 9 15
50 15 3 13 8 7 0 1 11 11 11 9 9 0 1 15 16 3 9 13 13 16 3 13 3 13 1 9 0 0 7 13 13 11 1 15 0 1 15 15 9 13 9 13 16 9 1 15 13 15 9
13 0 3 9 13 1 0 15 8 16 12 9 13 13
17 15 12 13 0 1 15 13 1 9 9 1 9 0 1 9 1 9
5 1 0 0 1 9
7 0 1 0 9 13 8 13
11 13 15 1 0 9 15 9 1 9 0 13
7 9 3 13 16 0 9 13
2 9 3
1 13
2 15 13
5 3 15 8 13 13
10 15 3 13 0 13 11 0 7 11 9
3 13 1 9
2 9 13
1 13
5 13 16 15 0 13
10 8 8 9 15 15 9 13 13 3 11
2 15 3
12 9 13 3 0 15 1 16 13 13 15 9 13
5 16 3 13 1 9
10 13 15 3 15 0 16 15 15 3 13
4 7 3 8 8
2 13 0
17 1 9 11 8 8 8 7 15 15 0 13 1 15 9 13 3 15
9 11 0 11 9 15 13 9 3 13
11 1 0 3 15 13 1 8 11 13 13 9
9 15 13 0 9 9 9 9 0 13
23 3 6 15 16 1 9 0 0 15 0 11 1 11 13 13 1 11 9 11 9 9 0 13
3 6 8 0
27 3 0 1 11 7 9 16 3 13 0 9 13 7 15 3 8 7 15 0 3 9 13 13 3 0 1 9
14 15 3 3 13 8 1 11 13 1 11 13 13 1 9
2 13 11
9 13 3 15 0 1 0 9 9 13
13 3 3 11 0 9 1 9 0 16 1 0 13 13
7 15 11 9 9 13 3 13
12 3 3 13 11 16 15 1 11 15 9 13 13
6 3 15 1 15 15 3
6 0 15 11 13 15 13
7 15 15 13 13 7 13 13
7 3 0 3 7 3 3 0
10 0 15 15 0 1 0 3 9 9 13
3 13 3 3
2 8 8
5 3 15 1 15 13
4 8 8 8 8
8 3 7 3 15 13 3 7 13
12 7 0 9 15 3 0 13 15 15 13 13 13
11 1 11 11 3 3 15 13 15 0 3 13
3 3 13 3
16 3 11 9 1 15 13 7 9 3 13 7 1 9 7 1 9
12 0 3 0 0 13 9 15 9 9 15 3 13
5 11 15 9 9 13
13 9 15 0 15 13 16 15 3 13 16 15 9 13
13 0 3 11 7 0 3 16 15 15 3 3 3 13
6 3 15 3 9 15 13
15 9 13 9 3 0 13 9 0 9 13 15 15 3 13 13
6 11 3 0 0 9 13
9 3 3 13 8 8 7 0 0 13
9 6 3 15 0 9 15 3 13 8
7 7 13 13 15 13 15 9
4 13 0 13 13
3 13 3 11
4 13 16 13 11
10 1 15 15 13 8 8 8 8 8 8
12 1 11 11 9 3 7 15 3 7 0 9 13
9 11 15 15 13 3 11 13 3 0
3 13 3 0
40 15 13 16 13 11 15 13 1 3 3 3 15 1 1 9 13 7 16 11 13 3 3 13 1 9 0 1 9 15 15 1 9 0 13 13 3 1 15 9 13
12 13 3 15 9 15 13 11 1 11 13 0 13
12 0 15 1 11 11 0 9 7 11 3 9 13
27 0 11 15 3 13 1 12 9 7 9 9 13 7 9 7 9 0 1 15 16 11 9 13 3 13 3 13
4 3 13 9 0
3 7 9 13
6 13 13 11 1 11 11
8 3 15 13 16 1 15 13 13
3 13 3 11
5 11 11 9 11 13
7 16 15 13 1 0 9 13
4 0 15 13 8
5 13 3 0 3 0
4 12 3 13 13
5 13 11 8 11 13
8 3 0 13 16 15 3 11 13
1 13
6 3 15 0 13 1 15
4 13 13 15 9
5 13 0 9 9 0
17 7 3 15 13 13 7 15 1 15 9 0 13 9 0 7 3 13
3 13 16 13
5 1 0 9 9 0
14 7 15 13 3 13 7 13 16 3 1 15 15 9 13
7 1 11 15 13 15 9 13
4 11 3 13 11
7 11 3 13 11 7 9 15
8 11 3 13 11 7 11 1 11
4 11 3 13 11
4 11 3 13 11
4 11 3 13 11
4 11 3 13 11
4 11 3 13 11
6 11 3 13 11 1 11
4 11 3 13 11
5 11 3 13 11 9
10 11 3 9 13 11 1 15 15 13 11
4 11 3 13 11
4 11 3 13 11
4 11 3 13 11
4 11 3 13 11
4 11 3 13 11
4 11 3 13 11
4 11 3 13 11
4 11 3 13 11
4 11 3 13 11
4 11 3 13 11
10 11 3 13 11 7 9 15 1 9 11
4 11 3 13 11
4 11 3 13 11
4 11 3 13 11
4 11 3 13 11
4 11 3 13 11
4 11 3 13 11
4 11 3 13 11
4 11 3 13 11
14 11 3 13 11 9 11 1 15 13 13 11 15 13 11
9 7 1 11 3 1 9 11 9 12
9 7 1 9 11 3 1 11 9 12
5 11 3 9 3 13
17 16 13 13 9 15 11 11 16 13 13 13 1 9 13 1 9 0
15 11 3 9 15 16 13 0 7 13 15 13 13 3 13 15
9 11 9 11 13 13 13 11 9 15
10 15 3 1 15 13 13 1 9 0 13
3 13 3 9
9 15 3 0 13 9 15 1 9 15
16 0 3 0 13 13 16 13 15 15 13 13 1 9 1 9 13
8 6 9 1 9 13 7 13 9
11 7 13 9 15 11 15 13 13 15 1 9
9 7 3 13 15 16 13 9 15 0
5 7 13 9 15 11
19 16 3 13 13 11 1 11 11 1 9 11 9 6 9 1 9 13 11 13
7 3 13 15 13 13 9 9
11 13 3 11 9 13 13 7 15 11 1 0
14 7 13 15 9 9 7 9 9 13 1 15 3 11 13
4 3 0 13 15
6 3 3 13 13 1 9
11 7 15 11 9 11 3 0 13 1 9 11
10 1 15 3 13 9 15 13 9 15 11
14 3 11 3 13 9 3 13 1 15 9 9 15 13 15
6 7 13 0 1 11 13
11 7 16 13 13 15 16 7 15 13 13 15
22 15 16 13 9 13 7 6 9 15 13 1 9 13 15 3 16 13 13 3 3 13 9
13 7 13 9 13 9 1 11 9 15 7 13 13 15
11 7 13 9 15 13 15 9 9 9 7 9
17 7 9 13 1 9 16 13 1 11 1 15 9 13 13 1 9 15
11 15 16 13 6 9 9 13 1 9 11 13
18 13 7 13 9 7 9 15 7 13 1 11 7 13 3 3 16 13 15
10 13 13 3 16 11 13 9 1 13 15
7 7 13 3 3 1 9 11
5 1 11 13 9 15
35 3 11 13 16 13 13 1 9 13 13 3 7 13 13 15 9 15 13 1 11 7 1 15 9 15 1 9 7 3 1 9 15 13 1 9
10 3 13 13 15 13 13 1 11 9 13
9 9 1 11 13 13 9 7 9 0
10 11 13 9 15 7 13 13 16 3 13
13 13 3 11 6 13 9 9 1 9 11 1 11 13
12 13 7 13 9 7 9 15 7 13 1 9 11
14 13 3 16 11 13 1 11 1 11 9 15 13 3 13
8 7 13 1 9 13 1 9 11
18 7 13 13 1 9 15 13 11 16 13 15 13 13 1 9 16 9 13
13 1 9 3 0 13 11 9 13 1 9 11 7 13
2 9 13
4 13 3 9 9
10 0 13 3 15 13 13 1 11 9 13
4 9 13 1 9
4 0 13 9 15
14 0 3 11 13 9 1 9 9 7 9 0 1 9 15
8 9 3 15 13 9 7 9 0
22 3 13 1 15 11 7 15 11 7 15 9 1 11 7 13 1 11 1 15 13 9 15
12 13 3 0 9 7 9 13 1 9 15 13 15
9 9 9 15 13 15 13 1 0 9
5 13 3 9 0 9
6 7 3 13 13 1 15
8 3 3 9 1 9 9 13 13
13 15 3 9 15 3 13 9 0 13 7 1 9 13
8 15 3 15 13 1 9 1 9
15 15 3 1 15 13 13 0 15 13 15 3 13 0 9 13
8 15 15 13 1 9 0 7 9
5 15 9 1 9 15
4 7 13 9 15
5 9 3 13 9 0
5 11 3 13 15 13
10 15 1 15 13 13 7 15 13 1 15
5 13 3 11 13 15
2 13 3
7 3 3 13 15 13 15 9
3 3 13 15
10 7 13 9 9 13 3 9 13 1 15
6 7 6 9 1 9 13
12 3 11 13 13 1 9 1 9 16 13 1 9
10 7 16 13 12 9 7 12 9 3 13
5 7 13 9 13 15
10 16 9 9 13 13 16 9 0 9 13
3 15 13 13
15 3 1 9 0 13 9 7 1 15 9 15 13 1 9 9
16 3 13 15 9 1 0 9 7 13 15 1 9 9 7 13 15
7 16 9 9 13 13 15 3
3 13 0 11
3 3 13 13
5 3 13 9 9 15
8 3 13 15 9 1 9 0 3
8 0 15 15 13 16 13 13 15
4 3 13 15 11
2 13 11
2 13 13
4 3 13 15 9
7 7 6 9 13 7 13 15
10 16 3 13 16 11 13 13 13 1 11
8 3 13 15 13 13 1 11 9
30 9 11 7 9 11 9 9 1 11 11 9 9 15 13 1 9 9 13 0 7 13 1 9 7 9 9 9 13 13 15
7 3 13 11 13 7 13 9
1 13
4 13 3 9 9
9 13 1 15 7 13 15 13 9 9
8 3 0 3 13 9 13 13 15
3 7 13 15
10 0 3 3 13 9 7 9 13 13 15
22 7 13 11 0 11 13 1 9 15 7 13 9 9 7 13 15 9 7 15 9 1 9
29 7 13 9 15 1 0 11 7 13 15 15 3 13 0 9 7 9 13 7 15 9 13 7 0 7 9 7 13 15
18 7 13 13 15 9 0 1 11 7 11 7 11 7 11 7 1 1 11
21 13 3 9 13 1 9 7 16 13 13 1 15 9 15 7 13 9 15 13 15 13
6 0 0 16 15 13 9
9 0 15 13 7 13 9 16 15 13
6 0 0 16 15 9 13
7 0 0 9 16 15 9 13
6 0 0 16 9 9 13
11 0 15 9 13 1 9 16 15 13 9 9
18 0 13 16 13 15 7 13 15 13 7 13 15 0 1 15 13 1 15
10 13 7 13 16 9 15 0 13 1 9
19 15 16 9 13 1 15 13 1 9 13 3 3 16 13 3 7 13 1 9
4 15 13 9 9
26 3 13 9 13 1 9 13 3 7 13 9 7 13 15 1 9 7 1 9 16 13 15 15 1 9 13
19 3 13 9 15 1 9 16 13 15 0 9 7 13 9 15 15 1 9 13
8 13 13 16 13 13 9 7 9
5 3 13 13 7 13
4 6 3 13 15
17 16 13 9 7 9 9 12 7 12 9 3 13 1 9 16 15 13
11 15 3 13 7 13 0 0 13 1 9 9
18 13 3 15 16 16 13 9 15 3 3 9 7 9 3 13 1 9 9
5 13 16 13 13 0
2 3 13
6 15 3 13 9 13 9
5 15 3 13 15 16
8 15 15 13 9 15 9 13 9
9 15 3 13 9 15 8 9 13 9
6 7 3 13 13 9 15
26 13 13 0 15 3 16 13 1 9 1 15 16 3 13 15 0 9 7 9 13 15 9 7 1 9 13
3 6 13 15
7 3 13 3 16 13 0 9
5 13 16 13 13 0
2 3 13
5 15 3 13 15 16
13 15 16 9 15 0 13 15 13 15 7 13 1 15
13 7 16 0 9 15 13 15 13 15 7 13 1 15
14 13 15 16 13 12 9 15 3 0 9 15 13 1 9
3 13 13 3
8 15 13 9 15 13 0 9 9
5 15 3 13 15 16
11 15 15 13 9 15 13 9 9 13 15 13
6 3 13 16 13 13 0
2 3 13
48 15 3 13 15 3 13 3 3 7 1 9 16 9 9 13 3 7 1 9 16 9 13 9 15 3 7 1 11 16 9 13 0 9 3 7 1 9 15 13 16 3 13 12 9 0 13 7 0
8 13 3 9 15 13 13 3 3
8 15 3 0 0 13 1 0 13
4 13 16 13 13
7 9 1 9 7 9 1 9
13 7 16 15 15 13 1 0 9 15 13 0 3 0
16 7 15 15 13 15 1 9 13 7 9 15 13 13 15 3 9
11 7 15 15 13 12 9 13 1 0 15 12
7 7 13 13 1 15 3 13
4 13 16 13 13
8 13 9 15 7 9 13 9 15
4 15 3 13 15
9 15 9 15 13 13 1 0 7 0
6 7 13 1 0 7 0
10 16 3 13 15 15 15 13 15 9 13
5 3 3 9 0 13
5 3 3 0 0 13
11 13 3 15 0 3 3 9 15 0 0 13
11 13 16 9 15 13 1 9 16 13 1 15
21 16 3 13 9 13 9 13 1 15 3 9 13 1 9 7 1 9 16 13 1 9
3 6 13 15
3 13 9 15
26 15 3 13 9 13 9 15 15 13 9 15 16 13 9 15 1 0 7 9 15 15 13 1 0 13 15
21 7 16 13 3 13 3 9 15 13 1 9 7 1 9 9 13 13 16 13 1 9
3 13 9 15
17 15 3 16 13 1 1 9 15 7 13 9 15 13 9 15 1 0
7 13 3 13 3 13 3 0
7 13 3 16 1 9 15 13
4 13 3 13 15
11 13 3 9 15 15 9 13 15 16 13 15
4 3 3 15 13
9 9 15 15 1 9 13 13 9 15
9 13 9 15 3 1 9 3 1 9
11 7 3 13 15 1 9 7 13 15 1 0
14 16 3 13 9 9 15 13 3 15 9 15 0 9 15
11 16 3 3 13 9 3 9 15 13 9 15
8 16 3 13 13 13 3 9 0
8 13 3 9 15 16 13 9 13
7 6 13 15 16 13 9 15
22 15 3 16 13 13 9 15 7 9 15 13 16 13 9 13 7 9 15 15 13 1 0
22 13 3 15 9 1 9 3 3 7 9 3 7 9 13 7 3 9 3 13 3 7 13
10 3 3 13 9 15 3 13 3 9 15
4 9 9 13 9
10 16 13 9 15 0 0 9 15 0 13
11 16 3 9 15 0 13 0 9 15 0 13
12 16 3 9 15 1 15 13 9 13 9 15 13
5 15 13 12 9 13
14 7 3 12 9 13 7 0 13 7 12 13 7 0 13
16 3 13 15 3 0 13 9 15 15 13 3 7 9 15 15 13
12 3 9 0 13 3 9 7 9 0 13 3 9
14 13 9 9 16 3 13 3 7 13 3 7 13 1 9
6 7 9 15 0 13 0
6 3 15 3 0 13 0
11 15 3 15 13 13 13 1 9 15 9 12
6 7 1 9 15 0 13
5 13 9 9 3 13
20 16 3 9 9 15 3 13 7 3 1 9 13 9 3 13 3 3 15 0 9
5 13 3 0 13 13
8 15 13 7 15 13 7 15 13
5 0 3 15 9 13
8 13 3 9 15 16 0 15 13
7 13 3 3 9 7 9 15
5 7 15 0 13 15
7 0 3 9 0 13 15 0
5 13 13 16 3 13
6 1 15 3 9 13 13
8 7 1 15 9 13 13 13 15
15 15 3 13 9 1 9 9 15 7 9 1 9 15 3 13
5 7 3 13 9 15
6 13 13 9 1 9 15
16 9 13 3 9 1 9 15 7 3 13 13 9 1 9 9 15
4 13 13 0 9
4 13 7 13 15
3 13 7 13
4 13 7 13 15
5 15 3 15 13 13
4 7 15 13 13
16 7 15 13 1 15 9 15 16 13 9 15 9 3 9 13 15
8 7 16 9 13 3 9 13 15
23 16 3 15 16 13 0 13 0 13 9 15 3 3 9 15 15 1 9 13 13 0 13 15
6 0 13 3 9 7 9
21 13 1 0 9 16 0 9 7 0 9 15 13 1 9 7 0 13 15 13 1 15
10 3 0 9 7 0 9 15 13 1 9
6 7 0 13 15 13 15
5 3 3 13 9 0
5 1 9 15 13 15
9 3 13 1 9 9 7 1 9 9
7 3 15 9 0 9 0 13
14 3 13 9 0 9 0 13 3 7 9 0 9 0 13
12 15 9 15 3 13 9 0 13 7 1 9 13
6 3 1 9 15 13 15
15 7 15 13 9 9 15 15 1 9 13 15 13 1 9 9
6 0 13 15 1 0 9
20 9 9 3 1 9 15 13 7 1 15 9 9 13 7 1 15 9 9 0 13
5 7 3 13 0 16
3 3 13 15
19 15 3 15 13 9 15 0 7 13 15 13 9 0 15 13 9 15 1 9
17 7 13 9 7 13 9 7 13 9 7 13 1 9 0 7 3 13
21 7 15 15 13 9 15 0 7 3 13 15 0 13 9 0 15 13 9 15 1 9
21 7 13 9 7 13 9 7 13 9 7 13 1 9 0 7 13 7 13 9 15 0
3 7 13 13
10 16 13 11 9 0 13 9 1 9 15
13 13 3 13 15 3 9 13 3 3 9 15 7 9
10 16 3 13 1 9 13 13 15 9 0
6 9 16 13 13 15 13
2 13 13
6 7 3 13 13 9 15
4 7 13 0 11
3 13 15 13
14 7 13 13 15 9 7 13 9 15 13 11 1 9 0
12 16 3 13 11 13 1 15 9 13 15 7 13
10 9 9 15 13 1 9 9 7 3 13
4 7 13 9 13
9 9 3 13 0 16 13 1 9 15
8 7 3 13 9 7 13 9 15
11 3 3 15 9 13 1 9 13 1 15 9
6 7 13 0 13 7 13
5 7 15 13 7 13
7 7 9 15 13 0 7 13
9 13 3 11 13 13 7 13 15 13
6 3 13 0 9 1 11
21 13 3 15 16 0 1 9 7 9 13 7 13 1 11 7 11 7 11 1 9 9
7 9 3 9 13 1 9 0
6 3 13 9 7 9 9
4 7 13 11 9
6 13 7 3 13 13 15
7 7 13 13 9 1 9 0
13 7 16 13 11 1 9 11 13 9 15 13 7 13
18 7 13 9 9 7 15 3 13 13 16 13 15 13 13 1 11 9 13
7 15 9 15 13 7 9 13
11 13 3 11 9 0 1 15 13 13 1 9
6 7 13 12 9 13 0
5 9 13 15 3 13
4 7 13 15 11
7 9 9 13 7 9 9 9
7 15 3 1 9 15 13 0
4 11 3 13 0
8 13 15 7 13 0 13 0 15
10 7 13 15 1 9 13 13 15 9 15
13 7 6 9 0 13 13 1 9 3 16 9 13 9
3 15 3 13
6 7 13 7 13 15 13
1 13
3 7 13 15
11 3 13 13 9 7 9 7 13 13 9 0
5 3 9 13 13 13
10 15 13 0 16 7 9 7 9 13 15
26 7 16 13 1 9 1 9 9 13 15 12 13 9 1 9 13 0 3 3 16 15 13 13 1 9 0
4 7 6 13 13
6 13 3 1 9 13 15
10 13 3 3 3 1 0 9 9 0 13
5 9 3 13 15 13
3 7 13 0
1 13
6 3 0 13 13 1 9
15 7 6 9 13 0 9 1 9 1 9 7 13 13 1 9
12 7 13 1 9 13 15 3 1 0 15 9 13
7 7 6 0 9 13 1 11
9 7 13 15 13 16 13 1 9 15
10 7 13 1 9 13 7 13 1 9 15
7 7 13 11 9 0 13 9
2 13 9
4 13 15 9 15
2 0 13
7 7 16 13 11 9 15 13
7 3 15 13 0 1 9 15
9 15 13 0 13 13 15 9 7 13
3 13 7 13
3 3 13 9
1 13
7 7 13 7 13 1 9 15
12 13 3 9 13 7 13 9 15 13 9 0 9
12 7 16 13 3 11 13 9 13 1 9 11 9
3 7 13 0
2 13 15
5 7 13 13 13 15
6 7 13 9 13 9 15
4 3 11 13 13
8 3 13 9 13 9 7 3 13
5 13 3 13 15 13
5 9 13 7 3 9
7 3 3 13 13 0 7 9
7 3 13 1 15 9 11 13
11 3 15 7 9 13 3 9 3 15 3 13
8 13 3 9 16 13 1 15 9
3 7 3 13
9 15 3 13 9 9 0 1 9 0
10 13 3 9 15 1 9 7 0 9 13
8 3 7 13 9 0 1 9 0
9 3 13 9 7 9 13 7 9 13
10 7 9 0 1 9 0 13 7 0 13
13 0 0 13 1 15 6 9 12 13 7 13 15 13
8 7 13 13 9 1 15 7 13
8 7 13 11 13 15 7 9 15
16 7 6 9 15 9 9 13 12 9 13 3 7 13 9 9 15
4 13 3 1 15
7 16 13 3 9 15 0 13
7 3 11 13 7 13 15 13
1 13
6 9 9 15 15 0 13
1 13
7 3 13 3 13 9 7 13
3 7 13 15
13 7 16 13 13 9 13 7 13 9 15 7 13 9
8 7 13 9 0 1 0 9 0
12 7 13 3 11 13 13 15 12 0 13 7 13
4 13 15 9 11
4 7 13 15 11
2 13 15
2 3 9
5 3 13 9 15 13
5 1 9 15 13 15
5 7 13 13 9 0
6 7 13 13 0 11 13
9 0 3 13 13 15 1 0 9 0
10 13 3 0 6 13 15 9 0 9 13
5 3 13 3 1 11
3 9 3 13
5 1 9 9 13 9
22 7 13 11 9 15 7 9 13 1 9 15 7 13 9 9 7 13 15 9 7 15 9
16 13 3 9 13 13 15 16 13 13 7 13 3 9 3 13 9
3 9 3 0
3 9 3 0
10 13 3 9 9 16 13 9 1 9 15
6 12 3 9 9 13 0
36 0 11 15 13 11 7 11 9 15 11 11 7 11 9 15 11 7 11 11 7 11 9 7 11 11 7 11 11 0 7 11 11 15 3 13 15
8 0 12 13 11 13 15 7 13
11 1 9 9 3 13 7 1 9 9 3 13
5 13 3 13 13 16
3 13 9 9
2 0 13
2 0 13
2 9 13
2 3 13
2 3 13
6 0 3 13 9 9 15
12 1 15 9 7 9 13 13 15 1 15 0 13
5 7 3 13 16 13
6 13 3 1 9 13 15
10 7 16 13 9 0 13 9 15 1 15
22 7 15 3 13 15 3 7 13 9 15 13 3 1 9 7 1 9 13 9 1 9 15
3 6 13 15
9 6 15 13 15 3 9 1 0 9
9 13 3 0 3 9 7 0 3 9
4 13 3 1 9
11 13 3 15 1 9 7 1 9 15 13 15
14 7 1 9 7 1 9 13 1 15 1 9 0 7 9
10 16 3 13 15 13 13 3 7 15 13
14 3 3 15 13 15 13 7 9 9 15 15 13 1 15
9 7 13 9 1 9 7 9 15 13
7 7 13 9 15 1 9 15
8 15 3 13 1 9 0 0 13
10 16 3 13 15 1 9 0 13 1 15
4 6 3 13 15
8 3 13 9 11 16 13 9 9
11 3 13 9 1 9 3 7 9 1 9 15
4 3 3 13 15
11 15 3 0 15 3 13 7 0 15 3 13
8 15 13 15 1 9 13 1 9
8 7 15 1 9 13 13 1 9
12 7 13 13 15 15 13 9 9 3 3 13 13
13 7 3 15 13 15 13 7 9 7 9 13 1 9
5 3 12 9 9 13
11 7 12 1 0 3 13 1 9 1 9 15
3 13 3 13
5 0 9 0 13 15
18 15 3 15 13 15 1 9 13 3 15 15 1 9 15 15 13 1 9
17 15 3 13 15 1 9 13 3 15 15 1 9 15 15 13 1 9
8 13 13 16 13 13 9 1 9
6 3 13 9 13 7 9
17 13 3 13 9 1 9 15 7 9 1 9 15 7 9 1 9 15
5 7 9 9 9 15
13 7 15 3 13 9 15 7 13 15 3 13 15 0
6 15 13 9 15 13 0
9 7 15 13 9 15 1 15 13 15
5 15 13 15 15 13
9 7 15 15 13 13 15 15 15 13
9 15 13 9 1 9 9 9 9 13
10 7 15 13 0 1 9 0 9 0 13
10 7 13 13 16 13 11 13 12 9 15
15 11 3 16 13 1 9 9 11 13 12 1 9 15 13 0
8 15 13 15 13 13 7 15 13
5 7 13 11 13 0
7 13 13 11 15 13 7 13
2 0 13
2 0 13
2 0 13
2 0 13
9 7 0 13 15 3 13 13 1 15
10 0 3 13 13 11 13 1 9 1 11
5 15 13 1 9 13
3 9 9 13
4 7 15 13 13
8 6 15 0 13 1 9 9 13
4 7 15 13 13
1 9
7 0 3 13 1 15 13 13
14 6 15 13 9 15 1 9 15 15 13 9 15 1 15
3 6 13 15
8 3 13 1 13 9 0 11 9
15 1 9 3 11 9 3 3 9 9 9 13 7 0 13 0
9 15 3 9 7 9 3 1 11 13
10 7 16 13 13 15 13 11 15 13 13
5 15 13 9 13 13
6 0 13 9 13 1 9
4 15 13 0 13
5 13 15 7 3 13
11 13 3 11 3 7 13 3 7 13 7 13
2 9 13
8 13 9 9 13 7 13 7 13
10 6 9 0 7 9 9 9 7 9 9
7 7 13 13 9 1 9 15
6 6 15 11 6 15 11
21 3 16 1 11 7 11 13 13 9 15 13 13 1 15 3 1 9 7 9 9 13
10 11 7 11 3 13 1 9 9 3 15
8 7 15 11 3 3 1 9 13
22 3 1 9 13 16 16 1 11 13 13 9 15 13 13 1 15 3 13 3 1 0 9
13 3 13 15 16 9 11 3 13 1 9 9 3 15
6 1 0 9 13 11 13
18 13 15 9 9 9 7 9 16 13 0 1 0 7 0 7 13 15 0
7 15 15 13 13 1 9 15
12 3 7 9 15 13 3 9 7 15 13 9 13
13 13 1 15 15 15 13 7 13 13 7 15 13 15
15 13 9 15 1 15 7 13 1 15 16 0 13 7 0 9
5 7 13 9 9 15
10 9 3 15 0 13 7 9 15 0 13
8 1 0 9 13 11 9 1 9
9 9 3 15 13 13 13 9 7 13
4 3 0 13 15
12 3 13 15 13 11 3 13 7 15 1 15 13
24 3 13 1 9 9 7 9 9 13 15 3 13 15 13 3 7 0 15 1 15 13 3 0 9
16 7 3 13 1 9 16 9 9 1 9 9 13 7 1 9 13
8 13 3 15 16 9 0 13 0
13 16 3 13 15 13 9 13 7 3 9 3 13 0
7 9 13 3 9 9 3 9
8 7 16 3 13 13 1 9 15
11 7 13 15 13 16 13 9 13 16 13 15
4 15 3 13 0
21 15 13 1 15 9 15 13 9 12 7 16 13 0 9 1 9 3 13 7 13 15
6 3 3 0 13 9 9
4 3 13 9 13
3 3 13 9
3 13 9 15
8 7 13 7 13 13 9 3 0
9 7 13 13 15 0 7 13 15 15
7 7 13 15 16 0 15 13
9 3 13 15 13 13 1 11 9 13
13 6 9 15 15 13 0 15 1 15 3 13 9 15
9 13 9 15 1 15 7 9 9 13
13 3 13 3 7 13 3 7 13 15 1 9 9 15
14 9 13 3 13 7 9 13 3 13 16 13 1 9 9
17 3 13 13 15 9 13 0 7 0 7 13 15 3 16 13 7 13
5 3 0 13 9 11
4 9 3 13 13
9 0 3 13 9 3 1 11 9 9
7 11 3 13 9 15 13 15
6 15 9 13 1 15 13
10 7 15 9 7 9 13 1 15 3 13
5 3 3 13 9 15
12 7 16 15 1 11 13 9 9 15 1 15 13
14 16 3 15 1 9 9 13 9 3 13 1 15 9 9
16 7 3 13 15 13 1 9 0 7 9 15 13 16 3 13 0
5 7 3 9 0 13
15 15 3 13 15 1 1 15 13 7 15 3 13 15 1 13
3 3 13 15
5 9 3 9 3 13
9 7 15 13 9 1 9 9 13 15
18 15 3 13 1 9 0 3 13 15 3 7 1 0 9 3 7 1 0
9 9 9 3 13 0 13 16 13 0
6 1 9 3 9 9 13
7 0 9 1 0 9 13 0
8 7 0 9 1 0 9 13 0
10 1 9 3 15 13 7 1 9 15 13
9 3 13 15 15 1 9 7 9 13
6 9 13 1 15 9 13
4 15 13 13 0
9 7 9 3 13 15 3 9 11 9
24 3 3 13 11 1 9 9 12 9 7 12 9 3 13 9 9 1 9 9 12 9 7 12 9
17 9 9 13 1 9 1 9 0 7 13 15 16 9 13 1 9 11
19 9 9 13 1 9 1 9 0 7 13 15 16 13 1 9 9 13 9 11
6 7 6 0 3 11 3
16 16 3 0 9 13 1 9 13 1 9 9 13 9 7 3 13
2 3 13
6 13 1 9 15 3 13
15 3 13 7 13 12 15 9 15 1 0 15 7 13 13 3
7 7 13 0 9 0 0 0
15 3 15 13 1 9 6 9 15 7 9 13 3 13 13 15
4 13 3 15 15
10 6 9 15 7 9 15 3 13 13 15
6 3 15 13 13 15 13
9 15 13 9 15 7 15 13 9 15
7 7 13 9 1 9 15 13
19 15 3 13 9 9 15 15 1 9 13 15 15 7 9 7 9 7 9 13
13 7 13 13 1 15 9 0 3 16 1 9 13 13
6 7 15 9 13 1 9
8 7 13 13 15 0 1 9 13
5 6 13 15 13 13
13 7 16 13 15 13 1 9 7 13 9 7 13 15
10 15 3 13 1 9 3 3 13 9 0
9 7 3 13 13 16 3 13 9 9
6 7 13 9 7 13 15
15 15 3 13 1 9 0 7 13 9 15 0 15 0 15 0
5 15 13 9 13 13
5 7 13 9 13 15
5 3 1 9 13 15
4 15 13 13 0
8 3 15 13 13 13 9 9 9
5 0 3 3 13 13
10 15 3 3 13 3 15 13 13 1 15
16 3 1 9 13 15 16 13 3 13 7 13 3 13 3 7 13
6 7 13 15 9 11 13
5 9 13 7 3 13
6 7 13 13 7 3 13
28 13 13 3 9 9 0 7 9 3 13 7 9 15 13 16 9 13 7 9 13 7 9 13 7 13 7 13 15
11 15 3 0 9 16 13 7 9 15 16 13
23 6 3 13 15 16 0 9 7 0 13 13 15 13 7 3 13 7 13 15 13 7 3 13
7 0 13 15 1 9 13 13
17 15 3 1 9 13 13 0 13 15 9 13 7 3 1 9 13 0
9 3 13 3 1 15 9 7 13 0
9 13 3 9 7 9 1 9 3 13
24 15 3 13 13 1 9 0 13 15 9 13 7 9 9 0 7 9 9 13 9 7 1 9 13
28 15 3 1 9 0 13 13 0 13 15 13 9 7 13 7 9 13 7 13 15 3 12 15 3 12 3 15 12
5 15 9 13 0 13
15 16 3 13 9 13 9 15 7 13 9 1 0 9 7 13
7 13 3 9 9 9 13 15
8 9 3 0 9 13 1 9 15
4 3 3 13 9
3 7 13 0
4 0 9 0 13
4 9 3 13 15
2 7 13
11 3 16 3 13 9 13 3 1 15 3 9
9 13 3 9 7 13 15 9 1 13
6 9 3 13 1 9 15
5 15 9 13 15 13
13 0 13 9 9 9 9 15 13 9 13 1 9 15
6 15 0 3 13 15 9
5 15 9 13 13 15
17 0 13 9 9 9 15 13 9 13 1 9 9 12 16 13 13 0
23 0 15 13 13 11 1 9 1 9 7 1 9 3 13 15 16 13 15 13 13 1 9 13
5 13 0 1 9 9
6 3 13 9 13 1 9
7 7 13 1 15 9 15 13
5 13 15 9 9 9
7 15 13 0 9 13 9 9
4 9 3 13 9
7 0 3 9 0 13 9 9
5 9 3 9 13 0
5 9 3 9 9 13
4 9 3 9 13
12 3 3 13 9 7 9 13 3 13 1 9 9
6 7 13 15 1 9 9
6 3 13 9 7 9 9
9 3 0 13 3 9 1 9 9 15
4 15 13 9 13
13 0 13 9 9 9 0 1 9 15 15 13 9 13
10 3 0 13 9 9 9 9 13 0 9
14 13 3 12 0 9 13 7 13 15 15 13 7 13 15
13 15 16 13 13 13 7 1 9 13 13 0 1 9
4 0 3 3 13
5 3 13 1 9 9
14 13 9 7 13 0 1 0 0 7 13 15 1 9 9
6 3 13 9 7 9 9
3 13 0 15
1 3
20 3 15 9 13 1 9 9 0 13 9 9 9 15 13 1 9 15 0 7 0
10 7 13 13 16 13 11 9 0 13 3
15 7 13 1 9 15 13 15 1 9 15 3 16 13 7 13
6 3 0 9 0 7 9
5 3 0 13 9 9
15 3 9 15 13 11 7 9 15 11 7 11 7 11 7 11
8 7 9 15 3 15 1 15 13
4 11 3 13 15
13 3 13 9 1 9 16 1 9 15 7 1 9 15
9 7 3 13 3 9 0 1 9 0
8 1 0 9 13 11 9 9 11
4 7 13 9 15
4 0 13 11 9
10 15 13 1 0 7 3 9 13 1 15
7 11 3 13 11 7 13 15
4 13 3 0 11
5 3 13 15 13 15
11 7 13 0 13 13 9 16 3 9 15 13
12 9 3 9 11 13 9 11 1 0 7 13 11
11 3 1 9 13 13 15 13 15 13 1 15
15 3 0 13 1 9 15 13 15 13 3 1 9 9 11 9
4 7 13 13 9
10 1 9 3 7 15 15 3 13 13 13
9 7 13 9 15 13 9 7 13 0
4 7 13 13 11
12 15 16 13 11 13 3 1 9 1 9 9 3
10 7 16 13 9 13 13 15 0 1 9
13 7 13 13 9 0 7 13 13 15 7 13 0 15
9 9 3 13 13 1 15 9 15 13
7 0 13 9 7 9 3 13
4 11 3 13 15
4 13 0 15 13
2 13 15
9 3 13 3 3 12 9 7 12 9
3 15 13 15
4 13 0 15 3
26 7 16 13 9 13 1 9 13 12 9 7 12 9 13 1 9 13 7 13 7 13 9 9 9 3 9
7 7 13 9 12 9 9 0
11 13 3 13 9 12 12 9 13 9 7 0
8 7 13 9 13 1 9 0 13
6 9 3 13 0 13 3
7 9 3 1 0 9 13 9
4 13 3 0 9
10 0 3 9 9 13 1 15 13 1 9
2 9 13
4 7 1 9 13
7 3 7 11 13 13 15 13
2 15 13
2 13 13
4 13 3 11 13
11 9 16 15 13 13 15 13 1 15 1 9
1 13
12 7 13 11 1 9 13 1 9 16 13 1 11
5 13 3 9 0 13
6 7 16 13 13 13 13
7 7 3 11 13 9 13 15
3 7 13 0
4 0 9 3 13
10 15 3 1 9 13 13 7 13 15 13
4 3 9 9 13
7 7 16 13 13 1 9 11
18 7 16 13 15 9 9 0 13 1 0 9 0 7 13 15 15 3 13
9 7 13 15 16 7 9 9 15 13
10 3 13 1 15 1 11 9 7 9 13
6 3 9 15 13 9 0
5 15 3 13 13 0
9 3 3 15 13 13 9 1 9 15
3 3 9 13
4 13 9 7 9
8 7 15 13 9 7 9 9 13
3 15 3 13
7 9 15 13 1 15 15 13
8 7 0 13 9 9 1 9 15
7 9 3 13 1 15 11 13
5 9 0 9 15 13
7 9 3 15 3 13 1 15
9 1 9 3 13 15 13 9 9 9
7 7 13 1 15 9 13 15
3 13 7 13
6 3 13 9 15 13 15
7 13 16 9 13 9 13 13
4 3 0 13 13
9 15 9 15 3 13 9 15 0 13
2 13 0
4 0 13 9 0
10 0 3 16 0 9 13 0 1 9 13
5 13 3 11 13 15
3 3 0 13
6 3 3 15 1 9 13
15 3 13 16 15 15 1 9 13 1 9 13 7 1 9 13
12 15 3 13 1 9 1 9 13 7 15 13 9
13 1 9 3 13 9 0 9 9 9 9 0 9 9
5 0 13 15 13 9
8 3 13 3 9 13 3 13 9
10 7 13 3 11 13 1 9 11 7 11
6 9 15 3 1 9 13
5 15 3 13 15 9
7 7 13 9 15 13 15 13
6 13 15 16 13 1 15
4 15 3 13 13
10 3 13 13 3 1 9 15 13 9 11
7 3 0 13 7 13 15 13
3 15 13 13
3 3 0 13
2 3 9
12 3 3 9 13 1 9 15 13 1 9 9 15
5 3 13 11 13 0
6 6 9 0 13 9 15
4 13 15 3 13
9 7 16 13 3 11 13 1 9 11
6 7 13 1 9 13 3
6 7 13 15 1 9 15
14 7 13 15 3 16 9 13 13 0 13 0 13 0 13
4 7 13 9 11
6 11 3 13 9 15 13
13 13 9 16 9 3 13 15 1 7 3 13 15 13
4 7 13 15 9
11 3 3 15 1 9 9 0 16 13 9 0
4 7 13 0 11
3 3 0 13
4 12 7 0 9
7 7 13 9 16 13 1 9
18 7 13 12 9 7 9 7 9 13 13 7 13 9 15 7 9 13 9
9 7 15 13 1 9 13 12 9 0
11 13 3 15 13 12 12 9 1 0 7 9
6 7 13 9 13 1 9
5 7 13 1 9 11
9 7 13 15 16 9 1 9 13 15
5 3 0 13 13 15
3 13 9 13
4 0 13 3 9
2 7 3
2 3 9
4 13 3 0 9
5 9 3 9 13 13
6 9 0 7 0 9 13
8 7 9 3 13 15 3 9 11
11 7 16 13 9 15 1 9 13 13 9 13
3 15 13 0
8 13 7 13 1 9 9 7 9
7 3 0 13 1 15 13 16
3 9 3 13
4 13 3 11 13
14 3 13 3 7 13 12 9 12 12 9 7 3 9 13
9 3 3 13 16 3 1 9 13 15
6 13 1 9 9 7 9
15 3 13 16 3 13 13 1 9 9 7 1 9 9 7 9
7 13 3 11 1 9 11 11
5 7 13 9 15 13
6 15 13 9 13 9 9
3 3 0 13
6 15 3 15 15 13 13
4 13 11 11 13
6 15 13 11 9 9 0
5 13 3 11 13 15
4 0 13 11 11
14 3 9 7 9 3 13 15 7 9 15 15 1 9 13
22 7 15 13 15 16 15 13 11 7 1 0 9 13 9 15 7 9 9 3 13 1 15
6 7 15 13 9 9 9
9 7 15 13 1 9 13 13 1 9
12 3 13 9 15 16 15 13 16 15 13 11 11
27 3 13 11 13 9 15 16 13 15 13 11 7 0 13 1 0 7 9 7 9 9 7 13 7 0 9 13
8 7 13 15 11 13 13 0 13
4 13 1 15 9
4 3 13 15 0
4 15 13 13 11
3 13 1 15
5 3 11 13 9 15
17 16 15 13 1 15 13 13 15 3 0 7 13 9 15 7 13 15
9 15 3 13 9 15 0 13 13 15
9 15 3 13 9 15 1 15 13 15
13 15 3 13 9 16 9 0 13 9 3 15 9 13
8 7 15 13 9 9 1 9 15
12 9 3 9 13 13 1 9 9 15 1 9 15
3 6 13 15
20 7 1 9 12 13 11 11 7 11 7 11 9 15 7 13 0 1 9 0 3
5 7 13 13 1 15
6 7 13 9 15 3 9
8 9 3 15 13 13 0 3 9
10 7 6 13 0 11 7 11 1 15 13
6 13 3 11 13 1 11
14 16 13 13 3 12 9 15 12 7 11 12 7 11 12
8 3 15 13 6 9 0 13 15
10 0 13 9 15 0 1 15 15 3 13
2 15 13
10 7 13 9 13 1 9 15 7 13 3
6 7 13 11 7 13 15
3 13 7 15
9 13 3 9 15 15 13 3 0 11
8 7 13 0 1 9 13 11 13
9 15 13 9 16 9 9 1 0 13
9 15 3 9 13 16 11 13 0 13
5 3 0 13 13 15
7 11 3 13 13 7 13 15
17 13 3 15 16 11 3 13 7 3 13 15 7 13 1 15 15 13
9 3 13 9 16 1 11 9 13 15
14 7 16 13 1 9 13 1 15 9 9 13 1 15 13
10 7 13 15 9 15 7 3 13 13 15
3 13 11 13
3 3 13 15
5 13 3 0 1 15
16 7 13 15 11 7 13 1 15 9 7 13 13 9 1 0 9
6 3 15 3 13 13 0
2 13 0
3 1 9 15
13 6 3 13 15 16 13 9 3 9 9 13 9 0
9 13 3 7 13 7 15 0 13 15
8 13 3 15 1 11 13 0 11
7 9 9 13 13 1 9 9
4 7 13 13 3
12 7 16 13 11 13 15 9 13 1 11 7 13
5 9 15 3 13 9
1 13
1 3
8 7 16 13 9 13 15 11 13
8 9 9 1 15 13 9 7 9
3 7 0 13
2 1 9
3 13 0 11
4 3 0 13 9
11 16 3 3 13 15 13 1 9 7 13 9
7 7 0 9 15 0 13 13
6 7 13 9 15 13 9
7 15 13 0 13 1 9 9
11 7 13 11 0 13 15 1 0 15 7 13
3 6 13 15
12 16 13 13 7 13 3 0 3 13 1 9 9
13 15 3 13 15 3 0 0 3 13 0 1 9 9
11 7 15 13 12 0 0 1 9 15 15 13
25 15 3 13 12 1 0 0 15 1 15 13 13 15 16 13 9 0 1 9 15 7 13 1 9 9
4 6 9 1 9
7 3 6 9 1 15 9 13
15 16 3 9 15 7 9 15 13 15 13 15 7 13 1 15
20 0 15 13 1 9 13 0 7 0 3 12 9 7 12 9 13 13 1 9 0
12 7 16 9 15 13 15 13 15 7 13 1 15
15 0 15 13 0 1 9 13 3 12 9 13 13 1 9 9
7 13 16 13 12 1 0 0
17 13 3 15 16 9 15 1 9 3 13 9 9 15 15 1 9 13
7 13 3 9 9 13 15 13
20 7 16 13 16 13 15 6 13 15 16 13 1 15 3 3 1 12 15 3 13
17 3 3 13 9 1 9 15 15 1 9 13 16 13 12 1 0 0
16 16 3 13 1 15 9 15 13 7 13 15 1 15 7 15 0
7 16 15 13 13 13 9 15
22 16 3 3 15 13 13 15 1 3 12 7 12 16 1 9 12 9 7 12 13 15 9
7 3 16 3 13 15 13 9
12 16 3 3 9 3 13 13 15 3 0 7 9
9 15 13 1 9 13 13 3 1 9
25 3 13 15 16 16 12 1 15 13 1 9 1 15 9 15 13 13 0 1 9 15 15 1 9 13
15 3 3 13 12 7 12 13 1 9 15 3 13 1 0 15
6 3 13 11 1 15 13
10 9 3 13 1 15 9 15 7 13 15
2 3 3
3 13 0 11
14 3 13 13 9 9 9 9 15 13 9 13 1 9 15
14 7 16 13 9 13 13 13 15 12 15 13 12 12 9
7 13 3 9 0 13 15 13
8 9 13 1 15 7 15 13 15
11 13 3 9 9 0 13 15 7 13 13 15
14 13 3 9 0 13 12 1 9 15 15 13 15 12 9
5 7 13 13 15 13
7 7 13 9 15 13 15 13
8 9 13 1 15 7 15 13 15
3 0 3 13
9 13 3 9 15 15 13 13 13 3
10 7 13 7 13 9 15 15 15 13 13
5 3 13 0 9 15
3 7 13 0
14 3 3 13 3 15 13 9 15 3 3 15 15 13 13
11 7 13 9 15 13 15 9 16 13 0 13
16 3 3 9 15 0 13 15 16 3 13 15 9 15 1 9 15
28 7 13 13 16 13 11 9 0 13 1 11 7 13 1 9 11 1 11 7 13 13 15 9 0 7 13 15 3
4 15 13 13 15
12 3 13 16 15 13 1 9 0 7 9 13 15
2 7 13
8 3 3 3 13 12 7 12 9
7 15 3 9 13 9 3 13
2 13 0
9 15 3 11 13 13 9 9 7 13
3 13 0 16
6 1 9 3 3 3 13
15 13 3 15 16 15 13 9 15 3 1 9 7 15 13 13
4 13 15 9 15
10 16 3 13 9 9 1 9 3 13 13
2 15 13
9 3 15 13 9 0 7 15 13 13
10 13 3 9 15 1 9 9 3 13 13
8 7 13 9 15 13 13 1 9
4 15 13 13 13
4 9 3 13 15
4 11 3 13 15
9 13 0 7 13 15 13 1 15 13
5 0 13 3 9 9
7 7 16 13 15 9 13 3
6 7 6 12 13 13 0
9 9 0 15 0 13 16 13 9 0
4 12 13 0 9
8 16 3 13 1 9 13 13 9
2 13 0
1 15
3 11 3 13
23 3 9 13 3 13 3 13 9 3 0 9 13 13 9 7 9 7 13 9 15 3 15 0
3 13 0 9
3 15 0 13
3 13 0 11
16 16 13 0 13 13 13 15 13 7 13 0 7 13 9 1 9
4 7 13 13 15
7 16 13 3 9 9 13 0
5 13 3 13 0 9
5 11 3 13 9 15
10 6 13 15 16 0 0 13 1 9 9
4 7 3 13 15
5 15 3 13 0 13
5 13 3 11 13 0
5 1 9 0 0 13
6 1 9 3 15 0 13
5 3 13 11 13 15
8 6 15 13 15 7 13 13 15
4 15 3 13 15
29 6 13 15 16 15 15 13 13 15 1 9 16 13 9 9 1 9 9 15 13 3 15 1 9 12 13 12 9 11
8 0 3 13 0 0 7 0 0
17 0 13 3 9 9 9 9 9 15 13 3 3 13 9 1 9 15
13 9 3 13 1 9 1 9 0 13 15 1 9 15
14 7 13 1 9 0 13 15 13 1 9 0 7 0 13
11 13 3 15 1 9 7 15 0 13 13 15
3 0 3 13
3 7 13 3
11 1 0 3 13 7 13 15 13 7 13 0
3 13 15 16
3 15 15 13
2 13 0
5 13 3 15 1 9
10 16 3 3 13 13 13 9 9 9 15
11 16 13 3 15 1 0 9 13 13 0 9
10 13 3 3 0 13 13 16 0 13 13
6 13 3 3 15 0 9
16 0 0 12 9 13 7 0 0 15 13 15 13 9 9 7 9
6 3 0 13 12 15 13
5 9 3 13 15 9
6 3 1 9 13 15 1
9 13 3 3 0 0 13 3 3 15
7 7 3 13 15 15 13 13
9 3 9 15 0 13 16 15 0 13
7 3 13 0 0 7 0 0
11 7 13 11 11 13 12 9 3 7 13 0
29 6 13 11 7 9 9 13 9 9 7 9 7 13 15 9 7 13 15 9 1 13 7 13 7 13 7 0 9 13
16 3 13 1 15 9 9 11 1 9 15 13 7 13 15 1 15
2 15 13
2 13 0
18 13 16 13 0 12 9 15 12 1 9 15 7 12 1 9 1 9 15
4 13 3 11 13
3 13 15 13
2 13 15
1 13
4 9 3 15 13
19 13 3 1 9 15 7 9 3 13 15 13 15 7 15 13 13 1 9 15
8 7 13 12 13 13 1 12 9
8 11 3 13 15 1 15 7 13
6 13 16 9 9 13 15
8 7 15 0 13 9 13 1 15
10 7 15 13 1 15 0 13 13 15 9
15 3 9 9 3 13 13 7 13 7 13 9 15 9 1 0
21 7 13 15 1 11 13 13 15 9 0 7 6 12 0 13 1 9 13 16 11 13
3 7 13 13
5 9 13 15 9 11
6 9 3 13 15 16 13
5 3 0 3 13 13
5 9 13 15 9 11
2 13 0
5 9 16 13 9 15
7 13 3 15 11 13 9 15
7 7 3 13 7 13 13 15
17 7 16 13 11 7 13 11 1 9 9 3 11 13 12 9 13 15
16 13 1 9 15 1 15 13 7 3 13 9 13 7 9 1 15
4 13 7 13 15
12 7 16 15 15 15 13 13 16 9 0 9 13
12 0 3 13 13 16 13 15 13 13 1 9 13
3 13 9 11
14 6 9 15 13 15 0 7 13 1 9 7 9 9 9
8 13 3 9 13 3 13 0 11
5 7 13 9 7 9
11 7 13 1 15 9 15 7 15 3 13 13
8 0 3 9 13 9 15 1 9
10 15 3 13 9 1 9 7 13 1 9
7 0 15 13 13 1 9 9
3 6 1 0
9 7 16 13 11 13 13 0 9 13
3 15 13 0
3 9 3 13
7 0 13 11 9 1 11 11
22 7 13 11 1 9 9 7 13 15 13 7 13 1 9 7 9 0 7 9 13 9 13
2 13 13
6 15 3 13 15 9 9
9 7 13 1 15 0 7 0 1 9
3 7 13 15
24 13 3 9 9 7 9 0 15 13 7 9 13 1 9 7 13 6 9 11 13 13 7 13 15
4 13 15 0 13
4 11 3 13 15
3 3 13 16
7 1 9 9 7 13 13 9
3 3 7 13
6 3 3 13 1 9 13
10 7 13 9 9 12 1 9 13 1 15
11 7 15 13 1 15 3 9 3 7 13 0
7 3 1 15 9 13 1 0
6 7 13 9 13 13 13
3 3 3 13
5 13 3 11 13 15
24 16 13 9 7 3 13 3 3 1 9 13 7 3 16 9 0 13 13 7 13 15 1 9 13
8 7 15 15 13 1 9 13 13
15 7 16 13 1 9 13 1 15 13 9 9 7 0 9 13
5 1 15 9 0 13
4 13 11 13 0
6 13 15 3 15 12 9
13 15 16 13 15 3 15 15 13 1 15 9 0 13
9 9 11 3 13 1 9 7 1 9
6 16 13 1 9 13 15
5 3 3 3 13 0
7 16 3 13 1 9 13 9
4 7 13 11 13
1 13
4 13 0 7 15
9 3 15 13 15 1 15 9 0 13
4 15 3 15 13
7 9 13 3 13 1 9 15
4 0 3 13 13
5 3 3 9 13 13
6 13 3 1 0 13 3
4 3 0 13 13
2 13 9
3 7 3 13
6 15 1 12 13 9 9
1 0
12 6 13 15 16 9 7 9 13 15 1 9 9
12 13 3 1 15 11 1 9 9 7 3 13 15
6 9 3 7 9 13 15
10 15 3 13 3 9 13 3 16 13 15
3 15 9 13
27 9 13 9 9 15 13 9 7 9 13 15 7 13 1 15 9 7 13 9 7 13 15 9 7 3 13 13
14 16 3 9 9 13 13 9 15 1 9 16 13 9 15
8 3 3 13 1 15 9 15 13
3 13 9 15
7 9 3 13 9 13 1 15
3 0 13 9
1 13
6 13 15 7 13 9 15
8 7 13 15 13 1 9 7 13
9 16 3 13 9 9 15 13 9 0
3 0 3 13
11 7 9 13 15 9 15 13 15 9 9 15
3 13 0 11
4 3 13 1 9
10 9 15 13 13 0 13 13 1 9 9
11 1 9 13 13 0 7 13 0 1 9 15
15 3 13 15 16 13 1 15 9 9 7 13 9 13 9 15
7 7 15 13 1 9 0 13
11 7 13 15 13 13 9 16 3 9 15 13
9 7 13 11 13 3 1 9 15 13
12 0 13 13 9 9 9 9 15 13 9 9 15
11 7 13 9 15 13 13 1 9 7 13 13
5 3 13 15 9 13
2 13 13
12 6 9 15 13 9 15 7 0 13 7 15 13
14 0 3 13 7 13 15 1 9 15 15 3 1 9 15
6 9 3 16 13 13 13
11 7 13 9 15 13 9 0 7 9 0 13
4 3 13 9 15
11 9 3 13 13 7 15 13 13 3 13 0
11 13 3 1 9 9 7 15 13 13 1 9
13 7 13 9 15 1 9 13 15 15 13 0 7 0
14 13 3 9 16 13 13 7 13 3 9 3 13 9 0
3 7 13 0
3 3 0 13
4 3 13 9 9
10 13 9 15 7 9 13 15 1 9 0
6 3 13 9 7 9 9
7 0 3 13 13 0 3 13
8 7 13 15 9 15 1 9 13
18 9 13 16 0 13 7 9 9 1 9 13 7 3 13 15 9 1 15
5 3 3 13 9 9
6 13 9 13 11 7 3
6 13 3 11 9 15 13
4 15 15 13 9
4 13 15 9 9
4 7 13 0 11
6 15 13 9 0 7 9
2 13 15
1 11
6 13 3 15 13 11 11
5 7 15 13 9 9
8 7 13 13 13 7 13 15 13
4 7 13 15 13
3 9 11 13
18 16 15 13 13 3 13 9 16 13 9 15 9 0 7 13 9 9 15
6 13 3 1 15 12 9
6 7 0 9 13 13 13
7 3 0 7 0 3 1 0
7 3 3 15 3 9 13 13
4 15 3 13 15
5 13 3 11 13 0
7 13 13 9 3 7 9 9
9 1 9 3 3 7 13 3 7 13
7 7 13 3 9 9 1 9
13 1 9 3 0 3 13 15 13 13 1 9 13 15
6 3 13 9 0 7 13
10 9 3 13 16 9 13 9 13 1 12
10 7 13 15 12 1 15 9 9 13 15
7 9 15 13 9 0 1 9
3 13 0 11
18 13 9 9 15 1 0 9 15 7 1 0 9 15 7 1 0 9 15
6 0 13 0 7 0 9
5 0 3 0 13 0
7 13 3 9 13 15 11 13
5 15 15 13 1 11
3 15 9 13
2 13 15
1 11
2 13 0
9 3 3 11 1 9 13 15 9 13
4 13 9 9 15
10 16 3 11 13 15 9 3 9 15 13
6 7 15 13 13 15 9
11 3 7 13 13 15 1 0 9 15 3 13
10 3 11 13 13 1 9 7 9 15 13
7 1 9 11 13 9 7 9
8 15 3 15 13 15 13 7 13
6 1 9 3 15 13 13
5 13 3 7 3 13
9 15 3 9 15 13 16 13 1 9
7 13 3 9 15 7 13 9
20 13 3 0 9 1 9 7 0 9 1 9 7 9 1 9 7 13 1 9 9
5 15 3 13 13 9
5 12 3 13 9 15
5 15 3 15 9 13
7 7 9 13 13 15 1 9
4 3 7 13 9
7 15 0 13 15 13 9 15
5 15 3 15 13 13
5 7 15 15 13 13
13 6 3 15 9 7 9 9 16 13 9 9 1 9
9 15 3 3 13 3 7 13 13 13
26 6 15 9 7 9 9 16 13 9 7 0 16 13 12 9 7 16 13 13 13 15 9 9 0 3 15
6 15 13 1 9 15 13
7 15 3 13 1 9 9 13
7 7 15 13 1 9 15 13
10 15 3 13 1 9 15 13 1 0 13
11 0 15 3 0 13 9 7 9 15 13 9
15 15 3 13 1 9 13 1 15 7 1 15 15 1 0 13
15 7 15 13 1 9 13 1 0 7 1 15 15 13 1 0
24 6 15 9 7 9 9 16 13 9 7 9 7 9 7 13 15 0 13 9 9 7 9 7 9
7 0 13 13 7 0 3 13
7 9 0 13 9 9 3 13
19 9 0 13 3 15 3 13 9 7 9 16 13 3 15 15 1 3 13 0
26 6 15 9 7 9 9 16 0 13 9 13 15 1 3 13 9 0 3 3 0 13 9 0 7 15 9
9 3 3 15 1 3 3 13 9 0
7 3 3 0 13 9 7 9
13 16 13 1 9 9 15 3 13 9 15 1 9 9
13 3 9 13 15 3 0 16 9 13 15 15 9 13
6 7 15 13 9 9 15
8 9 9 9 3 13 1 9 9
18 1 0 13 7 13 7 1 15 13 1 9 15 7 13 1 9 1 9
28 16 13 1 15 15 9 0 15 13 13 1 9 1 9 11 0 3 1 9 11 9 11 15 13 1 9 7 9
3 6 13 15
27 11 11 15 13 9 7 13 15 15 1 15 13 13 3 13 13 9 15 3 9 13 9 15 1 9 7 13
6 6 13 15 9 15 13
3 13 3 15
6 3 15 13 3 16 13
6 0 15 13 1 9 9
9 7 13 9 15 16 13 15 9 9
5 15 3 13 13 15
12 6 13 15 3 13 0 9 1 9 15 3 13
12 13 3 15 1 9 9 13 1 15 9 3 13
13 13 15 3 0 13 7 15 9 9 15 7 9 9
5 7 13 11 13 15
5 13 16 15 15 13
7 0 3 13 1 9 15 13
3 7 0 13
3 13 16 13
8 13 3 0 13 7 3 13 9
18 13 3 9 1 9 7 9 1 9 7 13 9 7 9 7 9 1 9
6 0 3 15 9 13 9
8 3 13 15 1 9 7 13 15
8 7 13 9 15 9 1 9 15
11 7 3 13 0 7 3 13 7 9 13 3
9 15 3 13 3 1 9 0 0 13
12 7 13 0 9 9 1 0 9 1 9 15 9
4 7 3 13 9
26 16 3 13 9 9 15 13 13 1 11 9 13 1 9 0 15 13 13 3 15 1 11 13 13 1 9
11 7 15 1 9 3 13 13 15 1 9 15
9 7 15 1 9 3 13 13 9 15
18 6 3 0 7 13 1 0 9 13 3 16 3 13 9 15 9 7 9
16 13 3 3 9 0 15 3 13 1 9 9 3 3 3 7 13
6 7 1 13 13 9 0
12 3 16 15 15 13 6 3 11 7 3 13 13
5 13 3 9 7 9
16 7 13 9 0 7 9 3 16 1 9 13 16 13 13 3 13
3 6 13 15
10 16 3 13 15 6 1 9 13 13 13
3 6 1 0
2 13 13
23 3 3 1 9 9 0 9 13 7 9 3 13 9 15 7 9 13 1 9 7 9 9 13
8 7 3 13 9 9 9 1 9
6 7 3 13 15 9 9
13 7 13 9 9 13 1 9 9 1 9 0 7 9
9 7 13 9 15 1 9 7 9 0
14 7 13 13 15 1 12 9 1 0 9 3 1 9 15
6 1 9 3 9 13 9
13 3 3 15 16 13 0 15 13 16 3 13 1 9
4 9 7 9 13
5 9 3 15 3 13
15 1 9 3 0 7 9 15 13 3 7 9 9 3 9 0
11 3 3 1 9 11 3 13 3 9 9 9
38 3 3 13 1 9 1 9 13 7 13 13 7 9 13 3 1 0 9 15 13 1 9 11 7 3 13 16 13 9 7 13 15 3 13 3 9 9 9
5 3 12 13 1 9
4 12 13 1 9
5 12 13 7 12 13
21 0 3 13 16 16 13 9 9 15 9 9 13 13 13 3 7 3 13 13 9 15
14 3 7 3 15 13 13 16 15 13 9 9 9 13 13
20 15 13 13 0 9 7 0 15 13 9 15 1 9 15 16 13 0 9 1 9
11 0 0 9 15 16 13 9 15 13 3 13
10 6 13 15 16 1 15 0 15 13 15
6 3 13 9 7 9 9
7 3 0 13 9 9 12 9
9 15 13 9 15 13 1 9 7 9
10 7 12 0 13 9 3 13 9 15 1
9 0 3 13 9 1 9 15 1 9
8 9 3 13 9 13 15 7 13
6 0 3 9 9 13 13
3 13 1 15
9 3 13 15 9 0 7 13 9 15
4 0 3 13 13
9 13 15 1 9 15 16 9 15 13
14 3 3 3 13 15 7 15 13 3 1 13 7 13 15
6 16 3 13 13 13 9
13 7 15 13 13 13 1 15 1 9 7 13 13 9
4 9 9 13 15
4 3 0 13 13
3 6 13 15
2 13 15
8 13 3 16 13 9 3 7 9
16 13 3 15 12 9 13 7 13 13 1 15 7 13 13 15 12
8 3 15 12 13 13 13 15 12
13 1 0 3 9 13 9 9 0 7 13 9 1 15
11 7 13 15 12 9 13 13 15 12 9 13
5 9 12 9 15 13
5 6 15 12 13 13
4 13 0 9 15
5 6 0 9 7 0
5 13 1 9 9 15
5 9 12 9 13 15
5 6 15 12 13 13
4 13 0 9 15
5 6 9 0 7 0
9 16 1 0 13 0 1 0 15 13
5 13 1 9 9 15
8 13 3 3 15 12 9 13 13
9 7 13 13 7 13 9 15 1 9
5 6 13 15 15 13
6 13 3 9 15 13 15
15 9 0 7 0 13 16 13 3 3 13 7 13 3 3 13
17 13 3 15 13 9 15 0 7 13 15 13 3 15 15 13 1 9
12 13 3 1 15 9 7 13 15 15 13 12 9
6 15 3 13 13 7 13
12 15 3 15 3 13 3 15 13 13 13 1 15
6 3 13 9 7 9 9
19 16 3 13 9 9 1 9 15 7 15 9 1 15 3 13 1 9 9 15
17 7 13 1 15 15 9 7 13 15 1 3 3 9 13 9 1 9
11 7 13 9 3 1 0 15 9 3 1 0
9 3 13 9 0 15 1 0 15 13
4 13 0 9 15
7 13 13 15 9 1 9 9
6 13 3 7 13 15 13
4 0 7 13 15
4 0 7 13 15
7 1 9 13 7 13 1 15
5 3 13 15 0 13
12 9 3 15 13 13 7 13 13 7 13 15 9
8 3 3 15 13 9 7 13 15
4 7 0 7 13
5 7 13 9 13 0
10 3 13 12 1 0 9 15 0 15 13
8 3 13 7 0 15 1 0 13
14 13 1 15 13 1 9 0 15 13 13 9 7 9 15
7 13 3 7 3 13 15 13
6 13 7 3 13 15 9
6 9 13 7 3 13 15
8 0 7 1 9 7 3 13 15
5 3 13 3 15 13
4 3 13 0 13
3 6 13 15
10 3 3 13 12 1 0 0 3 15 13
6 7 13 0 1 9 0
5 0 3 1 9 0
12 13 16 1 9 9 13 7 9 9 13 16 13
15 3 13 13 9 9 7 0 9 1 9 9 9 15 13 11
9 7 9 13 16 11 9 13 7 13
10 3 1 9 9 16 3 9 13 1 9
24 16 3 13 11 1 11 1 9 11 0 13 1 15 9 13 9 9 0 7 13 1 9 15 13
6 13 3 9 13 13 13
4 3 15 9 0
5 13 3 11 13 0
4 15 0 13 9
6 9 0 13 13 1 15
6 3 3 0 13 15 1
12 13 3 0 9 0 1 9 15 1 13 15 13
3 6 13 15
16 3 13 13 0 9 1 0 9 13 3 15 0 13 1 9 15
3 7 13 0
9 15 13 15 13 7 15 15 15 13
6 3 0 13 15 12 0
7 7 3 13 9 16 15 13
8 0 3 9 13 9 1 11 13
3 3 11 13
8 13 1 9 1 15 7 13 15
4 9 15 3 13
7 1 15 13 9 1 9 15
10 7 13 9 3 13 0 11 7 13 9
7 9 3 13 13 1 12 9
4 7 13 0 13
9 6 13 15 16 12 15 15 13 13
4 3 15 13 9
10 15 13 15 1 9 1 9 0 15 13
9 9 3 9 13 3 13 13 1 0
18 6 3 9 10 1 15 9 9 13 0 13 15 16 13 3 13 9 0
7 13 3 11 15 13 15 13
4 3 15 13 9
2 13 0
2 15 13
4 0 13 9 15
5 7 13 9 9 13
4 7 13 0 13
4 13 1 0 15
14 0 13 3 9 15 0 9 15 1 0 13 1 9 9
3 13 3 15
21 3 13 3 1 0 9 9 3 1 9 0 3 0 13 15 1 0 1 9 9 15
7 7 9 13 13 1 9 9
9 15 15 9 13 1 15 1 0 9
3 13 13 3
6 13 9 7 13 9 9
7 16 3 13 13 15 1 11
5 13 3 11 13 0
10 3 16 15 13 13 1 15 15 3 13
3 13 0 11
13 6 13 15 16 1 0 9 16 9 13 3 15 13
5 3 7 15 9 13
14 3 13 11 1 0 1 9 15 13 11 7 13 9 15
7 13 3 16 13 3 7 13
12 7 13 11 7 12 9 11 13 13 7 0 13
3 3 13 0
7 0 13 9 15 3 1 9
6 13 3 7 13 15 1
10 15 9 16 0 13 13 1 15 9 0
11 7 13 1 9 7 13 15 13 7 13 11
8 3 3 13 12 9 13 15 1
8 13 7 13 16 3 13 1 9
7 9 3 0 13 9 3 0
6 3 3 13 7 13 13
14 9 15 16 3 13 0 9 13 16 13 0 13 9 15
5 13 3 9 15 13
11 7 13 0 3 13 7 13 3 0 9 13
4 13 3 7 13
10 6 13 9 7 9 9 13 1 9 13
1 13
1 13
5 6 13 15 15 13
8 15 3 13 15 13 0 9 13
5 15 13 13 15 13
2 13 15
2 6 9
4 7 13 13 15
4 13 7 0 11
4 9 1 15 13
22 7 6 12 1 0 15 13 1 11 13 9 13 9 15 7 13 9 9 9 13 9 15
4 3 13 0 11
6 13 9 15 1 9 15
7 15 3 15 13 9 9 13
8 3 3 13 9 16 3 13 13
6 1 0 9 13 11 9
10 3 1 9 13 1 9 7 9 13 15
9 0 3 0 13 13 16 13 9 9
6 3 9 15 13 15 13
14 3 0 13 11 13 1 11 9 9 3 9 7 0 13
11 11 3 13 15 1 3 3 1 9 9 9
9 7 13 3 13 1 9 16 13 9
8 7 3 13 16 0 0 9 13
8 3 3 13 12 0 9 7 13
9 13 13 9 9 7 1 9 13 0
6 7 13 9 9 13 0
9 15 13 1 15 15 0 1 15 13
3 11 3 13
5 7 9 9 13 0
14 13 15 1 9 0 16 13 15 16 15 13 11 9 9
2 15 13
13 3 13 9 9 13 1 0 9 7 13 1 9 9
7 3 9 9 13 9 15 13
1 13
4 15 3 13 9
4 6 3 13 9
3 15 15 13
4 3 0 13 13
8 15 3 9 1 9 15 13 13
3 13 15 11
5 15 13 15 15 13
6 11 3 13 3 1 9
7 7 13 1 15 12 9 13
6 3 15 1 11 9 13
6 3 0 13 1 15 13
3 13 15 13
6 3 0 13 1 11 9
6 7 3 13 1 9 16
3 3 13 9
9 7 1 0 13 15 13 7 13 11
6 3 7 15 1 0 13
7 3 7 9 15 0 15 13
9 3 13 13 7 13 16 3 13 9
4 7 3 9 13
5 7 13 3 13 3
17 3 3 13 9 13 15 9 9 7 0 9 1 11 16 15 9 13
9 7 13 13 15 7 13 11 11 9
19 3 13 11 15 15 13 16 13 13 9 13 13 12 0 9 9 7 0 13
4 13 13 9 0
3 3 0 13
3 15 1 15
6 7 13 0 1 9 13
6 9 3 9 13 0 13
10 3 13 13 15 1 9 16 9 9 13
11 9 3 13 13 1 0 9 9 1 9 9
13 1 0 13 13 9 10 11 9 9 3 1 0 9
10 3 13 13 15 13 13 1 11 9 13
11 7 13 12 0 9 13 15 13 1 9 11
10 11 3 13 1 9 7 13 15 9 13
4 15 13 9 9
2 15 13
10 7 16 13 1 9 9 7 0 15 13
4 3 13 0 11
7 3 13 15 1 15 13 9
12 7 3 13 15 1 15 9 3 16 13 9 3
8 13 3 3 13 0 15 13 11
5 13 3 0 13 11
10 15 13 13 15 11 7 11 15 13 11
11 13 3 0 1 9 13 1 0 9 15 13
5 15 15 7 0 0
9 0 3 13 13 3 1 9 1 15
13 9 3 9 7 0 13 9 16 13 11 11 3 13
6 15 13 15 1 12 13
3 3 0 13
1 11
3 13 0 11
2 13 15
1 13
3 13 0 9
5 3 0 3 13 13
1 13
17 13 3 11 16 15 13 7 3 9 13 13 9 13 9 1 9 13
7 0 15 13 1 9 0 0
2 15 13
8 9 15 1 15 7 1 9 15
4 3 13 0 11
12 3 9 9 13 11 1 9 13 1 15 0 9
21 7 13 15 9 0 13 15 7 13 9 1 9 13 1 9 15 7 9 1 9 15
7 7 9 13 1 15 13 13
3 6 9 9
10 7 13 1 15 13 9 7 13 9 15
17 7 16 13 15 13 15 9 7 13 15 9 15 7 13 15 16 13
6 0 13 16 13 9 15
8 7 13 15 9 13 1 9 13
5 7 16 13 13 13
13 16 3 13 15 13 9 15 9 13 7 13 13 15
8 7 13 1 9 15 9 15 13
5 0 13 11 9 9
14 3 13 13 1 15 12 9 12 1 0 7 12 1 0
9 13 3 13 15 13 9 15 7 13
10 3 3 9 9 13 1 9 7 0 13
3 15 0 13
6 15 0 3 13 0 13
11 16 9 11 13 13 3 1 9 7 13 15
3 13 1 9
5 13 3 15 16 13
3 13 3 16
3 9 9 13
14 1 0 3 9 9 13 13 1 0 9 3 1 9 0
9 7 1 9 0 13 11 9 0 13
4 8 8 8 8
2 0 13
8 9 15 9 15 3 15 13 15
7 15 3 3 13 7 13 13
3 11 13 0
17 7 3 13 12 1 15 13 9 13 9 7 13 9 7 13 15 13
6 13 16 13 11 13 15
8 11 3 3 13 9 0 13 9
13 7 6 9 9 13 13 1 12 9 1 0 3 3
12 7 9 13 13 7 9 13 13 7 9 13 13
7 7 0 9 0 15 13 13
14 7 13 1 9 1 9 15 13 1 0 9 7 13 0
18 9 3 7 15 1 15 13 13 11 13 9 7 0 15 13 13 3 13
15 13 3 3 9 0 1 3 15 13 13 11 1 11 13 15
19 16 3 3 13 13 13 15 9 0 1 11 9 11 15 3 0 9 13 11
8 0 13 1 11 7 13 9 11
5 3 11 13 13 9
19 7 13 9 11 13 0 9 0 7 13 0 1 9 15 0 15 13 1 9
9 7 13 9 0 1 9 9 7 13
11 13 3 3 11 11 7 0 11 13 1 9
9 9 13 13 16 9 10 13 3 13
4 1 12 9 13
3 13 1 0
6 7 13 0 9 0 0
3 13 0 11
2 13 9
1 13
9 0 3 13 13 9 13 9 1 9
16 9 3 9 15 13 1 0 9 13 11 11 7 0 11 13 9
6 7 6 9 13 13 0
8 7 13 13 9 7 13 1 15
6 13 3 9 15 3 9
5 7 9 15 3 9
12 1 9 3 15 13 13 9 7 13 13 3 0
3 13 13 15
8 13 3 16 11 15 13 13 13
3 3 13 3
4 13 3 3 13
6 13 9 3 13 13 9
8 7 3 13 13 9 15 16 13
6 7 6 13 15 1 11
3 6 13 15
14 7 13 3 1 9 1 9 7 0 9 13 13 9 15
6 7 6 11 13 0 13
1 13
10 0 3 13 7 13 9 15 7 13 15
2 13 13
1 13
3 3 15 13
18 15 16 13 6 15 1 9 13 1 9 7 13 9 9 15 15 13 13
11 7 13 1 0 9 13 9 0 13 9 13
12 13 16 9 15 9 13 7 13 13 15 15 13
14 7 16 0 13 13 1 9 15 13 15 7 0 15 13
8 3 0 13 9 13 3 13 13
12 12 3 9 13 1 11 1 9 3 13 0 11
3 15 3 13
7 7 13 11 13 13 15 13
10 13 13 15 15 9 1 9 7 1 9
22 13 3 13 15 9 13 15 1 9 9 7 9 7 9 0 13 15 13 15 15 13 15
12 7 6 15 15 1 13 15 9 3 1 9 9
6 9 9 11 11 9 9
6 3 13 13 1 11 9
3 13 9 9
4 0 13 9 15
32 13 11 1 9 13 7 13 9 9 1 9 9 7 13 1 0 15 11 9 7 9 0 7 13 1 0 1 11 9 13 9 15
18 7 13 11 13 9 9 7 9 0 1 9 15 7 9 7 9 0 13
3 7 13 13
14 13 0 15 1 15 15 3 13 0 13 13 9 9 15
4 15 13 15 9
6 0 3 13 15 9 0
12 13 11 1 11 11 7 13 13 1 11 1 11
17 7 3 13 1 9 13 13 9 7 9 3 9 13 7 13 1 15
6 7 9 13 13 1 9
5 15 13 9 15 0
3 1 15 13
16 7 3 9 13 15 1 9 7 13 1 9 12 9 7 12 9
4 7 13 1 11
8 13 7 1 9 7 9 13 0
4 13 7 13 9
22 7 13 1 9 11 13 11 7 11 9 15 13 9 1 9 13 3 9 7 13 15 11
9 13 1 15 7 13 15 13 9 9
7 7 3 13 9 13 13 15
17 7 13 3 3 13 11 11 7 11 9 15 7 15 1 9 13 9
4 7 3 13 0
12 7 13 9 15 11 1 9 1 9 13 13 15
7 7 3 9 13 9 13 15
11 13 3 13 15 3 9 13 7 3 3 9
9 7 13 1 9 15 9 1 9 0
3 7 13 13
6 15 15 7 15 11 9
3 13 13 15
3 13 15 13
6 7 13 13 15 11 13
5 13 7 13 1 9
10 7 13 13 15 3 16 13 1 15 13
3 15 13 0
14 15 9 0 0 16 1 9 3 9 0 13 7 13 15
9 7 13 9 15 3 1 15 9 11
15 7 3 13 1 9 13 1 9 11 7 11 1 11 7 11
6 7 3 13 15 1 0
7 7 13 13 15 13 9 15
8 7 3 13 15 9 7 13 15
7 7 13 15 9 13 1 9
19 7 13 0 15 13 0 9 7 9 0 13 7 3 13 13 15 16 13 15
12 7 9 3 13 13 13 1 0 9 3 7 13
10 7 13 13 15 11 7 15 1 0 13
3 15 13 15
3 7 13 0
10 13 1 0 9 7 9 16 3 3 13
4 1 0 3 13
7 7 13 1 15 0 13 15
4 7 9 13 13
5 16 13 13 15 13
5 7 13 15 13 0
1 13
1 13
11 7 16 13 3 13 1 15 9 7 13 13
9 7 13 15 3 13 0 7 13 15
2 7 13
15 13 15 9 9 7 13 1 9 15 15 13 11 1 9 0
27 7 3 13 11 1 9 7 13 13 16 1 9 13 7 13 0 3 16 3 13 3 1 9 7 13 15 9
10 7 13 13 1 15 9 15 1 12 13
13 7 16 3 13 13 15 0 1 9 13 9 3 13
8 7 13 13 9 1 15 9 13
8 16 13 3 11 9 0 13 9
4 9 13 15 9
4 15 0 3 13
7 15 13 13 9 3 0 9
13 15 3 13 11 9 15 16 3 13 1 15 13 0
6 15 0 13 1 9 15
17 15 13 0 13 9 13 15 9 7 13 13 7 13 9 15 7 13
14 16 3 13 16 9 13 9 9 1 9 13 9 13 9
2 15 13
1 13
15 7 13 9 13 1 15 3 16 13 15 7 13 9 13 16
3 3 3 13
15 7 13 13 3 1 9 15 7 9 13 1 15 7 13 15
12 7 16 13 13 11 11 13 1 9 7 13 0
2 13 15
5 7 13 13 13 15
19 7 13 13 16 13 1 9 0 0 9 7 9 3 13 1 11 7 9 15
7 13 3 0 15 7 13 15
10 3 1 9 7 9 13 7 13 9 15
5 0 13 11 13 0
9 3 3 13 0 9 7 15 3 13
7 3 3 13 13 0 7 9
7 7 13 9 11 7 9 13
5 7 13 7 13 0
6 3 9 11 7 9 13
5 15 3 9 3 13
9 15 9 13 15 1 9 3 13 13
8 13 3 9 3 13 1 15 9
6 7 3 13 1 0 9
7 15 9 9 0 13 9 0
10 3 13 9 0 1 0 7 0 9 13
8 7 15 13 9 0 1 9 0
10 3 13 9 9 7 9 13 7 9 13
17 7 13 13 3 16 9 13 1 9 7 9 15 13 13 7 13 9
7 6 15 13 9 15 3 13
3 7 13 0
16 3 13 15 13 11 3 9 13 7 13 15 7 15 1 15 13
26 3 13 1 9 9 1 11 9 9 7 9 9 13 15 3 13 13 3 9 7 13 15 15 1 15 13
3 7 13 15
10 9 1 9 13 13 7 3 9 1 9
4 7 13 3 9
7 7 13 3 9 13 9 0
6 7 13 9 13 9 0
3 13 1 0
3 7 13 15
6 13 9 3 13 7 3
5 9 0 13 7 13
12 7 13 15 1 9 13 1 9 9 15 13 9
3 13 9 15
7 7 13 7 13 13 9 0
8 7 11 1 9 15 13 1 9
19 7 0 9 1 11 7 11 13 13 15 7 1 11 7 1 11 7 1 11
14 7 15 1 11 7 11 9 0 13 15 13 13 1 15
13 7 13 9 15 16 9 15 13 1 9 16 13 15
8 7 9 0 16 0 13 13 15
3 7 13 13
4 15 13 9 9
7 7 3 13 15 16 13 0
4 7 13 1 15
12 7 13 16 13 12 1 0 7 16 13 15 13
9 7 13 0 9 13 9 7 13 9
41 7 11 11 7 11 9 11 7 13 15 9 11 15 13 9 9 7 11 7 11 7 11 7 11 7 11 7 11 11 7 11 7 11 0 7 11 11 15 7 13 0
4 7 13 1 9
11 7 13 3 9 3 16 3 13 3 9 13
7 7 16 13 15 13 13 15
7 13 3 16 1 9 13 13
7 7 13 15 1 9 13 0
5 3 13 11 11 13
13 7 16 9 1 15 3 0 13 3 13 9 0 13
17 7 16 11 13 1 15 3 0 13 13 7 3 13 13 7 9 13
17 15 13 9 0 13 1 9 13 16 3 0 13 7 3 9 15 13
13 6 13 15 16 15 13 9 9 9 7 9 15 13
16 15 3 13 1 9 0 3 13 9 1 0 7 9 13 0 9
2 3 13
6 7 13 9 15 7 9
3 7 13 15
9 6 9 15 7 9 15 3 13 15
4 7 13 15 13
7 15 13 9 15 7 9 15
9 7 13 15 15 1 9 15 13 13
6 6 9 15 7 9 15
14 15 3 13 9 9 0 9 15 7 9 15 7 9 13
12 7 13 15 1 9 0 7 13 0 1 9 15
1 13
5 6 13 13 1 13
13 7 16 13 15 13 1 9 7 13 9 7 13 0
10 15 3 13 1 9 3 3 13 9 0
9 7 3 13 13 16 3 13 9 9
6 7 3 13 13 9 13
7 7 3 16 3 13 9 13
10 7 13 9 7 13 0 7 9 3 13
6 7 15 13 1 9 0
16 7 13 9 13 7 13 7 13 12 12 7 12 12 7 12 12
2 7 13
5 15 13 9 13 13
14 7 16 13 0 13 15 0 15 1 15 13 1 12 9
3 7 13 15
6 15 13 13 9 9 9
8 13 9 0 7 3 15 9 13
4 15 13 9 13
24 0 3 13 15 1 9 3 13 9 7 16 13 3 13 11 7 13 9 15 13 13 1 9 15
8 7 0 13 3 15 1 9 13
9 15 16 13 9 3 1 9 13 0
9 7 3 13 9 1 15 7 0 13
9 3 13 9 7 9 1 9 3 13
22 0 13 15 9 13 7 9 9 7 9 9 7 1 0 9 13 13 9 7 1 9 13
3 7 13 0
10 3 13 9 16 1 9 13 7 1 9
5 3 16 1 9 13
8 3 3 13 15 0 15 3 13
10 3 7 13 13 0 7 16 1 3 13
6 16 15 13 9 13 13
3 13 15 13
10 1 15 9 13 13 13 15 7 13 15
10 7 15 3 13 3 15 13 13 1 0
2 7 13
26 3 13 9 9 3 16 9 13 9 1 9 7 13 7 13 9 7 9 7 9 13 7 13 16 13 0
13 3 3 9 13 3 9 3 9 3 0 9 1 9
11 7 16 15 13 9 3 13 9 16 13 9
4 15 13 9 9
5 7 15 9 13 0
17 3 9 9 15 16 13 13 1 9 0 13 15 9 15 13 1 9
10 7 0 0 9 13 15 9 3 13 13
6 1 9 3 3 13 15
6 3 3 9 15 13 15
9 7 13 0 0 9 16 3 13 13
10 7 13 9 13 15 3 3 13 1 9
6 7 15 9 13 1 0
15 7 13 13 9 0 9 7 9 13 1 9 3 16 13 9
8 7 13 15 1 9 1 9 13
7 9 3 1 15 13 16 13
8 7 13 13 13 9 7 13 9
1 13
3 7 13 9
5 7 13 13 9 0
3 7 13 0
3 15 0 13
3 3 13 9
11 15 13 13 0 16 7 9 7 9 13 15
8 7 13 1 9 9 1 9 9
16 16 3 9 7 9 13 13 9 7 9 13 7 15 13 15 13
16 7 3 9 7 9 1 9 7 1 9 13 13 7 13 15 9
9 13 3 11 1 3 13 7 13 15
5 7 13 9 0 13
8 15 15 7 15 11 9 9 0
4 13 15 1 9
3 13 3 0
3 7 13 15
4 15 15 9 13
3 7 13 15
7 11 9 15 13 16 0 13
9 7 13 15 3 16 15 13 1 9
9 13 3 3 1 9 9 9 0 13
5 7 13 15 9 13
7 7 13 9 0 13 1 9
16 7 0 9 9 13 13 1 9 1 12 12 7 13 13 1 9
12 15 3 13 15 13 7 13 1 9 7 1 9
7 7 13 13 13 15 13 13
4 7 13 1 11
14 7 13 0 15 1 9 13 13 13 7 0 9 7 13
15 7 13 0 15 13 3 13 13 15 15 9 13 7 1 9
9 7 13 15 13 16 13 1 9 15
17 13 1 9 15 1 15 7 13 0 15 15 9 13 7 13 13 15
11 7 13 7 13 13 1 11 15 15 13 11
3 7 15 13
18 7 16 13 11 1 9 3 1 9 13 9 0 1 0 7 13 1 9
20 7 13 15 1 9 9 11 7 13 15 13 1 9 15 7 13 15 3 13 16
5 9 15 1 9 13
1 13
9 13 9 1 15 16 0 13 7 13
10 13 3 16 16 7 9 15 13 0 13
7 7 3 13 13 9 9 15
8 7 13 9 16 13 13 1 9
17 7 3 11 13 1 15 3 0 9 15 13 1 15 13 1 9 13
4 15 13 9 15
5 7 13 15 9 15
6 13 9 13 15 7 13
7 7 13 13 15 15 0 13
4 0 3 13 15
6 9 9 15 15 0 13
9 13 1 9 7 13 0 1 9 15
12 3 15 13 13 1 9 13 16 9 15 13 13
4 15 3 13 9
8 11 3 9 15 13 13 13 9
3 3 3 13
14 7 3 13 15 13 15 3 11 7 11 7 11 9 11
4 7 13 13 15
4 15 13 7 13
6 9 3 13 13 7 13
3 7 13 15
20 15 3 13 15 13 9 7 9 9 7 15 15 1 13 7 13 3 13 9 13
5 8 8 15 13 13
3 9 15 13
1 13
4 13 3 9 12
4 7 13 9 0
8 7 13 0 3 16 15 15 13
5 7 13 13 0 13
5 7 13 0 9 15
7 7 13 9 13 1 9 13
8 7 0 13 13 1 9 15 13
4 3 0 0 15
14 3 0 13 9 9 11 9 11 7 11 7 11 7 11
8 3 3 9 15 3 15 1 13
4 7 13 1 0
17 3 13 9 1 9 3 1 9 15 7 1 9 15 7 1 9 15
13 7 3 13 3 9 15 13 16 0 0 13 9 13
11 7 13 1 9 15 7 13 9 1 9 13
3 7 13 12
11 7 13 15 13 0 7 13 0 9 9 0
3 7 13 15
9 3 13 1 9 3 13 16 13 3
6 7 13 13 16 9 13
11 7 9 0 13 7 13 9 0 0 7 13
13 7 13 11 9 0 3 13 13 9 15 7 13 16
5 11 9 13 1 0
6 7 3 13 9 1 0
4 15 3 13 16
3 15 3 13
4 15 13 11 13
8 15 15 13 11 0 1 0 13
21 0 3 11 13 7 13 11 7 13 15 1 9 1 11 9 11 9 15 16 13 15
4 13 3 11 11
7 3 13 15 13 9 9 15
4 11 3 13 0
7 7 13 13 15 3 7 13
16 7 16 9 0 13 11 9 15 9 13 9 7 9 7 0 11
17 16 7 13 9 15 11 7 13 7 13 11 3 7 13 9 13 9
8 13 1 15 15 13 7 13 15
4 7 13 0 16
8 15 13 13 15 3 9 9 15
6 15 16 13 13 9 15
2 15 13
3 7 0 13
10 16 7 13 3 1 9 1 9 13 13
10 13 16 3 13 15 1 9 9 11 9
13 7 13 9 1 9 13 7 1 3 13 13 15 13
9 7 13 9 13 13 9 15 1 9
11 7 13 15 1 9 7 13 9 15 1 9
9 7 13 0 9 7 9 13 9 15
9 15 13 9 15 13 7 13 9 15
5 7 13 0 1 9
8 13 3 1 0 9 7 13 3
7 13 3 15 13 7 13 0
5 7 3 13 9 13
9 7 13 1 9 13 1 0 9 3
7 7 13 15 13 7 13 0
11 7 0 3 1 15 9 13 3 7 13 15
6 7 13 13 0 9 11
10 7 16 3 9 0 13 13 9 15 13
14 13 0 16 13 1 0 9 7 9 13 15 9 15 13
4 7 13 13 0
3 13 0 13
3 7 13 15
9 13 13 9 12 9 7 13 15 13
3 7 13 15
3 13 7 13
4 7 16 13 13
12 7 13 0 16 13 13 15 1 9 1 0 9
9 7 13 1 9 1 0 7 1 0
22 7 13 12 9 7 12 9 13 1 9 13 7 13 9 7 13 9 15 16 13 1 15
5 7 12 9 13 15
6 7 13 15 7 13 13
7 13 3 15 13 12 12 9
18 7 3 13 9 15 13 9 16 13 15 1 9 1 11 16 15 13 9
8 7 16 13 15 13 1 9 13
22 7 13 15 13 1 13 13 3 9 0 15 7 1 0 9 9 13 1 15 13 1 9
4 7 13 13 15
13 3 0 3 13 15 13 1 9 13 9 13 7 13
7 15 3 15 13 7 13 13
1 13
2 15 13
2 13 13
9 7 13 1 0 1 9 7 13 9
5 3 3 13 1 9
5 13 3 9 0 13
9 7 16 13 13 1 9 11 7 13
18 7 13 0 9 0 13 1 9 15 15 15 3 13 13 3 13 15 13
29 7 3 13 1 9 7 1 9 7 9 1 9 13 0 7 13 15 16 7 9 9 15 13 7 3 13 15 0 13
12 7 13 1 15 9 7 15 1 9 13 1 11
16 7 16 13 15 1 9 15 0 9 15 13 3 13 13 9 13
14 9 3 7 15 9 16 3 13 9 3 13 13 9 0
17 7 15 0 13 15 13 13 0 13 9 9 7 9 7 9 7 9
6 7 13 15 9 7 9
5 3 0 13 13 15
9 3 13 11 1 15 9 3 13 13
5 9 0 9 15 13
7 9 3 15 3 13 1 15
9 1 0 3 15 13 13 9 9 9
11 13 3 9 9 13 9 9 9 9 7 9
3 7 13 0
3 11 3 13
6 13 9 15 7 9 15
8 7 15 13 9 7 9 9 13
3 15 3 13
34 16 13 9 9 7 9 8 15 13 9 15 1 15 15 13 7 3 3 13 15 15 13 9 15 7 9 13 9 9 1 9 15 15 13
6 7 0 0 9 0 13
6 7 13 3 9 13 0
6 16 15 13 9 13 13
12 7 16 13 1 9 1 9 13 15 9 15 9
3 7 13 0
5 3 7 15 0 13
12 3 13 16 15 3 13 1 9 3 13 15 13
16 3 3 13 1 9 15 7 1 9 7 1 9 13 13 15 9
10 13 3 16 15 1 9 13 0 13 9
22 1 3 3 1 9 9 9 0 13 9 9 9 9 9 9 9 9 9 0 9 9 9
9 7 3 13 13 1 9 11 7 11
10 7 13 9 15 13 13 7 3 13 13
18 9 3 3 3 13 1 15 15 13 9 9 0 13 7 13 1 9 15
6 13 3 9 9 11 9
9 7 13 15 16 9 13 1 9 15
3 15 13 0
4 13 3 13 9
10 3 13 3 0 13 9 9 7 13 9
3 7 13 0
4 1 0 9 13
5 13 9 1 9 15
13 7 16 13 9 15 13 9 13 1 9 7 9 13
16 7 3 13 1 9 11 13 1 11 1 9 11 1 0 9 11
13 7 13 15 0 7 0 7 13 15 16 13 0 9
11 7 13 15 1 9 3 13 9 15 1 9
8 7 13 1 9 13 7 13 0
15 7 3 13 13 9 15 7 13 13 9 9 15 7 13 3
6 7 13 0 16 15 13
8 3 3 15 13 0 3 0 13
5 7 3 3 13 13
3 3 15 13
7 7 0 13 13 7 0 13
3 13 1 9
11 3 6 3 9 13 15 3 7 13 15 13
7 15 3 1 15 1 3 13
5 7 13 15 9 15
9 3 0 13 15 3 13 9 1 9
9 7 13 15 3 9 13 15 13 12
6 7 13 9 13 1 9
4 7 13 9 0
6 7 15 13 7 13 13
13 7 13 7 13 13 7 13 15 13 1 9 12 9
3 7 13 15
11 7 3 13 9 1 9 15 13 1 9 11
16 7 13 9 7 13 13 1 15 13 1 0 9 1 9 13 15
4 7 13 9 13
8 6 13 15 16 13 9 0 9
8 7 13 15 13 3 13 1 9
5 7 13 13 13 9
10 7 3 12 9 3 13 15 1 1 9
1 13
7 13 1 9 9 7 9 11
6 7 13 1 15 13 16
5 15 13 11 13 0
6 15 13 16 9 3 13
5 3 13 3 7 13
5 3 13 13 9 15
4 9 13 3 13
16 3 7 13 3 12 9 13 1 12 12 3 3 9 9 0 13
2 13 15
11 3 3 12 9 1 12 12 3 9 9 13
3 7 13 15
1 12
3 7 13 15
3 3 3 13
13 7 13 11 7 13 15 0 7 13 15 16 0 13
13 7 13 1 9 15 13 9 15 13 15 16 15 13
5 13 9 3 9 13
7 3 3 13 9 1 9 15
3 7 13 13
8 7 13 13 3 16 13 3 15
7 7 13 0 1 9 15 13
4 13 1 9 15
7 7 16 1 9 13 15 13
5 15 15 13 13 9
6 15 13 0 13 11 9
2 15 11
6 15 3 3 12 1 9
3 3 13 0
6 15 3 15 15 13 13
4 13 11 13 15
3 15 13 11
27 7 13 13 0 16 13 9 9 0 13 7 13 1 0 7 1 0 9 7 9 7 13 7 1 12 9 13
4 7 3 9 13
7 7 13 15 11 13 13 15
10 15 13 7 13 9 15 13 13 11 13
14 13 1 15 11 16 3 13 15 9 13 7 15 13 9
8 7 13 9 1 9 15 13 15
16 16 15 13 1 15 13 13 15 0 7 13 9 15 7 13 15
9 15 3 13 9 15 0 13 13 15
8 7 15 13 9 9 1 9 15
28 15 3 15 13 13 7 15 9 1 9 0 0 7 9 7 9 9 13 15 16 13 1 9 9 15 1 9 0
3 7 13 0
20 6 13 15 16 13 15 1 3 13 15 3 13 9 16 13 9 9 13 1 9
24 7 1 9 12 13 11 11 7 11 7 11 7 13 0 1 9 0 3 0 7 13 13 1 15
18 7 9 15 13 13 13 0 3 3 9 15 9 1 9 3 13 0 13
6 7 13 0 11 1 11
5 7 13 11 13 11
12 7 13 12 9 15 12 7 11 12 7 11 12
5 3 3 13 15 13
4 13 3 9 13
6 7 13 13 9 13 15
6 7 13 9 1 9 13
5 0 13 9 15 0
11 7 3 13 15 3 13 3 11 3 15 1
19 7 13 0 1 9 13 0 16 15 15 13 13 3 16 9 9 1 0 13
4 7 13 15 13
11 15 3 13 9 7 9 16 11 13 13 3
4 15 13 13 0
6 11 16 13 3 13 15
12 7 3 13 13 1 9 9 16 0 13 7 13
15 7 13 1 9 15 13 9 0 1 15 7 9 13 1 0
12 7 3 15 9 13 15 13 13 7 13 13 15
3 7 13 15
6 7 13 12 1 9 13
9 9 13 9 15 1 15 13 9 0
13 15 3 15 13 13 15 7 13 7 13 9 7 13
10 7 13 9 15 16 13 0 7 3 13
7 6 9 0 3 1 15 13
3 3 15 13
4 13 0 1 15
3 7 13 15
6 7 13 1 9 13 13
12 7 13 9 15 15 9 13 1 15 0 15 13
3 3 0 13
13 7 3 15 7 1 9 7 1 9 13 16 15 13
8 7 16 15 13 13 15 13 15
4 11 3 13 0
6 16 13 13 15 0 13
8 7 3 13 9 9 1 9 13
3 13 9 15
12 7 16 13 11 13 9 13 13 9 0 13 0
3 13 1 15
6 7 3 3 13 1 15
21 7 13 7 3 13 15 13 1 15 7 13 13 3 0 3 16 0 13 16 13 13
9 11 3 13 9 15 13 0 7 13
10 7 16 13 1 9 9 15 3 13 15
6 3 15 3 13 13 15
11 0 9 1 15 13 13 3 1 9 7 9
5 3 7 13 15 13
8 13 3 9 15 7 13 0 16
14 9 9 13 1 9 9 7 13 15 7 13 0 9 13
4 3 0 13 9
4 7 13 15 13
3 7 13 11
6 15 16 3 13 13 15
7 7 13 13 12 7 13 0
11 16 15 13 0 13 13 15 0 7 15 9
8 7 13 9 13 15 1 0 15
6 15 16 13 13 13 0
12 15 12 1 0 9 9 13 1 9 15 15 13
12 7 15 15 13 3 15 13 7 15 15 15 13
4 13 0 11 13
15 9 13 15 1 9 15 13 9 15 3 13 15 7 13 15
3 13 13 15
16 15 13 3 15 13 9 1 9 15 7 13 3 3 13 1 15
9 15 3 3 13 1 15 1 15 13
20 15 3 9 13 15 9 9 1 9 15 16 11 13 6 13 15 3 13 9 15
24 7 15 13 12 1 0 0 13 1 15 0 13 15 3 16 13 9 0 9 15 7 1 9 13
8 7 16 13 15 9 15 13 0
26 0 13 15 0 13 1 9 3 12 9 13 13 1 9 1 9 0 3 9 15 3 13 7 9 3 13
8 7 16 9 15 15 13 13 0
25 0 13 15 0 13 1 9 9 3 12 9 13 13 1 9 9 3 9 15 3 13 7 9 3 13
8 15 3 9 13 7 15 9 13
3 0 13 9
9 3 16 9 0 13 1 15 0 13
9 13 1 15 9 7 9 13 1 15
9 7 3 13 13 1 9 11 1 11
6 7 13 3 9 1 15
12 7 13 9 13 15 16 13 9 9 13 13 15
4 15 15 13 11
2 15 13
7 11 13 9 9 13 7 13
4 15 13 11 13
8 1 9 9 15 13 15 9 0
10 1 9 3 9 0 7 9 13 15 9
6 7 13 12 1 9 12
8 3 3 3 13 12 7 12 9
10 7 1 9 3 9 15 1 0 13 15
3 7 13 0
11 15 13 9 15 7 15 13 9 13 1 15
10 7 16 9 13 9 15 7 15 13 13
7 7 13 0 0 16 13 0
9 15 16 13 11 3 13 7 13 0
9 13 0 13 1 15 7 3 13 15
5 0 13 3 9 9
11 15 3 13 9 9 3 0 3 13 1 0
10 7 13 15 7 13 9 1 0 13 15
14 7 16 13 13 1 9 13 15 9 13 1 15 13 15
8 9 0 15 13 16 9 0 13
4 15 15 13 0
5 15 0 3 12 9
20 9 13 3 13 3 13 3 13 3 0 9 13 3 9 13 13 9 15 7 9
5 7 0 13 13 0
9 11 3 13 15 13 15 7 13 0
3 12 15 13
1 13
2 7 13
2 13 15
6 15 13 1 9 13 13
5 13 3 13 9 0
6 7 13 11 13 9 15
6 9 3 13 1 9 15
6 3 11 3 13 13 0
13 3 13 9 1 9 9 13 3 0 13 1 9 9
8 15 3 13 13 1 15 3 0
5 7 15 13 0 13
5 7 13 0 11 13
8 1 9 0 13 7 3 1 9
6 15 3 0 13 1 9
8 6 15 13 15 7 13 13 15
3 6 13 15
50 15 13 15 13 9 7 9 7 9 7 9 7 9 7 9 7 9 1 15 7 1 9 15 3 13 3 3 3 1 9 0 9 7 9 7 9 7 9 7 9 7 9 1 9 7 1 9 0 9 0
8 0 3 13 0 0 7 0 0
7 13 3 1 9 13 1 11
6 7 13 0 11 7 13
3 7 13 13
11 7 13 3 12 13 0 13 15 13 15 13
4 7 0 9 13
10 7 13 1 0 11 7 11 9 11 13
7 9 13 16 15 13 13 15
4 3 0 13 15
5 15 13 16 13 15
2 7 13
16 13 15 16 12 1 9 15 7 15 1 9 15 13 1 9 15
4 11 3 13 15
12 13 13 9 15 15 13 7 9 15 15 13 13
4 3 0 13 15
1 13
4 11 3 13 15
12 9 3 15 15 13 13 7 9 15 15 13 13
16 13 3 1 9 15 7 1 9 3 13 15 13 7 15 13 13
9 7 13 12 13 13 1 11 7 11
6 11 3 13 15 13 0
14 3 3 13 3 1 15 7 15 13 13 0 13 15 9
10 7 15 13 1 15 0 13 13 15 9
19 3 3 9 9 3 13 16 13 15 7 16 13 7 13 9 15 9 1 0
3 7 13 11
19 7 13 15 1 11 7 9 15 7 0 9 9 11 11 0 13 1 9 13
11 15 16 13 16 11 9 13 13 13 7 13
5 9 11 11 13 15
5 3 0 3 3 13
6 7 13 11 13 0 13
5 7 13 0 13 15
2 0 13
1 13
2 13 15
8 15 13 9 15 13 13 1 15
4 15 13 15 13
4 0 3 13 15
4 11 3 13 0
1 13
5 9 15 15 0 13
8 7 3 13 7 13 15 1 9
17 7 16 13 11 7 11 1 9 9 13 12 1 9 15 7 13 0
4 13 0 7 13
17 7 16 15 15 13 15 13 13 16 9 0 13 7 3 0 13 3
10 7 13 13 9 13 1 9 3 1 9
7 7 15 1 3 13 13 0
4 15 13 13 9
10 15 13 15 3 13 0 11 7 13 15
5 7 13 9 1 11
7 0 3 9 15 13 1 9
10 15 3 9 13 1 9 7 13 1 9
8 7 15 13 7 15 13 13 13
1 6
7 0 15 13 9 9 15 11
3 6 1 9
5 7 13 11 1 9
8 7 15 9 16 13 1 11 13
15 16 7 13 1 3 9 13 9 13 16 15 3 13 1 15
9 7 16 13 1 15 15 13 1 9
5 3 3 13 9 9
4 7 13 13 15
4 7 13 9 15
3 7 13 11
8 7 9 0 7 9 13 9 13
9 7 3 13 16 15 9 13 1 9
4 7 13 13 15
11 3 13 13 16 9 15 9 9 13 15 9
6 15 3 13 15 9 9
10 15 13 9 9 7 9 13 3 15 13
8 7 16 9 13 13 13 1 9
5 7 13 11 13 15
6 9 6 9 15 13 13
5 7 13 11 13 0
3 13 9 9
3 6 13 15
23 15 13 0 9 13 7 13 1 9 7 3 13 1 9 15 7 13 16 15 13 13 13 15
3 3 13 15
16 15 16 15 3 13 3 9 15 15 1 9 13 13 15 9 15
4 7 13 3 11
14 7 16 13 1 9 13 1 15 0 9 7 9 7 0
3 7 13 0
5 1 15 9 0 13
9 7 15 15 13 0 9 16 0 13
5 11 3 13 13 0
6 13 15 3 15 12 9
8 9 11 1 9 13 7 1 9
2 13 15
6 3 0 13 15 1 13
10 16 13 1 9 13 3 3 3 13 15
4 7 13 1 9
2 13 9
8 15 3 13 11 16 3 9 13
4 7 13 13 11
9 3 15 13 15 1 15 9 0 13
6 7 13 0 1 9 13
20 9 13 9 7 13 9 7 13 9 7 13 9 7 13 15 9 7 3 13 13
14 7 13 1 9 1 9 9 16 1 9 13 1 9 9
7 15 13 15 13 7 13 0
7 7 3 13 1 0 15 9
7 7 0 9 13 7 9 13
14 3 3 12 13 9 0 3 0 13 1 15 0 13 16
5 9 3 13 1 3
3 0 13 9
1 13
2 13 15
4 7 15 13 9
8 7 13 15 13 7 13 1 9
8 13 7 13 9 7 13 9 15
5 3 7 9 0 13
11 1 9 13 13 0 7 13 0 1 9 15
4 7 13 15 13
3 7 13 9
8 13 3 16 1 15 9 0 13
4 7 13 15 13
4 15 13 13 15
9 9 13 16 0 13 7 3 13 15
13 3 7 3 13 1 9 9 7 1 9 9 9 13
6 15 13 9 15 13 0
3 15 15 13
5 13 15 9 16 13
3 3 0 13
6 15 13 9 0 7 9
2 13 0
1 11
5 13 3 11 13 0
4 7 13 1 15
10 7 13 1 15 9 15 13 9 3 13
4 7 13 15 13
4 12 3 9 13
10 7 0 13 9 7 13 13 3 13 9
7 7 0 13 15 7 13 13
5 7 3 0 13 9
3 7 0 3
4 7 3 13 9
6 0 15 13 13 3 9
5 12 3 13 15 9
5 7 13 11 13 0
10 3 3 13 3 13 9 3 7 9 9
17 16 3 1 13 13 3 7 13 3 7 13 7 13 3 9 1 9
17 1 13 3 16 13 3 13 1 9 11 1 9 3 13 0 9 13
10 15 13 9 11 7 9 11 7 9 11
4 15 3 3 13
5 11 3 13 15 16
4 0 15 9 13
2 13 11
6 9 9 15 9 12 13
24 7 13 9 9 15 1 0 9 15 7 1 0 9 15 7 1 0 9 15 7 1 0 9 15
4 0 13 0 9
4 0 3 0 0
4 7 13 0 9
14 3 9 1 9 13 16 12 13 7 3 13 15 1 15
30 7 16 13 1 0 9 7 1 0 9 7 1 0 9 7 1 0 9 7 13 9 3 15 0 0 13 15 9 7 9
8 11 3 13 16 3 13 13 0
6 3 13 3 1 9 9
6 7 15 3 13 15 13
7 7 13 11 13 13 1 9
7 3 13 9 11 9 13 11
4 13 9 9 15
11 13 1 0 15 16 13 9 15 9 9 15
11 0 3 11 13 15 9 7 3 13 9 15
6 7 0 9 15 3 13
6 7 13 15 1 9 15
24 13 1 9 15 13 1 9 13 7 13 1 9 7 1 0 9 13 1 9 7 0 9 1 9
12 15 13 9 9 1 9 0 9 0 13 0 9
17 7 13 11 1 9 13 3 9 13 9 1 9 7 0 0 13 0
14 6 13 15 16 9 0 0 0 15 13 15 13 1 9
8 15 3 1 15 15 13 0 13
12 0 3 1 9 15 15 15 13 13 0 9 15
11 7 16 13 1 9 13 0 12 1 9 15
7 9 13 15 9 7 15 9
5 7 13 11 13 0
5 13 0 15 0 9
18 7 16 13 1 9 9 1 9 13 15 3 11 7 11 7 11 7 11
9 7 15 9 13 3 0 15 13 13
6 7 13 11 13 13 0
5 13 16 15 15 13
10 0 3 13 1 9 15 13 16 15 13
3 7 0 13
9 16 13 3 9 7 9 9 3 13
3 7 3 9
16 13 3 9 1 9 7 9 1 9 7 13 9 1 9 7 9
5 13 3 15 3 0
19 13 3 15 9 7 1 9 13 7 1 9 7 9 13 1 15 1 9 0
8 7 1 15 9 0 13 13 9
9 7 16 13 15 13 13 13 15 13
10 7 15 13 15 13 1 0 9 15 13
9 13 3 9 9 1 9 7 9 9
9 7 13 9 1 9 7 9 13 15
7 7 13 9 15 1 9 15
20 16 3 13 9 9 13 3 3 13 15 13 13 3 15 1 11 13 13 1 9
17 7 15 1 9 3 13 1 9 3 7 13 16 13 15 1 9 15
11 7 15 1 9 13 3 13 3 13 9 15
8 6 3 0 7 13 1 0 9
20 13 3 9 0 9 0 15 3 13 1 9 9 15 13 9 3 3 3 7 13
10 7 16 13 9 9 3 13 0 15 9
7 7 1 13 15 13 13 9
14 7 3 16 15 15 13 6 3 13 11 6 3 3 13
3 15 3 13
4 6 13 15 15
15 7 1 0 9 1 9 0 9 13 7 9 3 13 9 15
13 7 3 13 9 9 13 1 9 1 9 0 7 9
19 7 3 13 9 15 7 13 13 15 1 12 9 1 0 9 3 1 0 9
5 1 9 3 13 9
16 16 3 9 15 0 13 7 13 13 9 13 16 1 0 13 9
14 3 3 15 16 13 0 13 13 16 1 0 13 1 9
4 9 7 9 13
5 9 3 15 3 13
1 13
3 13 7 13
5 13 3 3 9 13
22 3 9 15 3 13 13 9 15 7 13 9 15 9 15 9 7 9 13 16 13 13 3
6 13 3 3 9 9 13
16 3 7 0 9 7 9 9 7 3 3 16 13 3 13 15 13
1 13
12 7 13 0 9 7 9 3 15 9 13 7 13
2 13 3
9 3 1 9 0 16 3 9 13 9
18 7 16 13 11 1 9 11 0 7 13 13 9 13 9 9 9 0 0
7 7 13 9 13 1 9 15
12 13 3 15 3 13 1 15 3 0 7 13 16
6 15 9 0 9 13 13
3 11 3 13
2 13 15
4 15 0 0 13
6 0 9 13 13 1 15
6 3 3 0 13 15 1
6 7 16 13 13 0 13
5 15 3 3 3 13
4 15 13 0 13
3 6 13 15
16 3 13 13 9 0 1 0 9 3 15 13 0 13 1 9 15
14 7 11 11 12 1 12 13 1 0 9 16 13 15 0
4 15 13 13 13
6 7 13 15 9 15 13
6 7 13 3 0 3 13
10 7 0 9 9 3 9 13 13 15 9
9 3 13 13 7 13 15 16 13 9
11 13 15 7 3 13 13 9 9 16 9 13
10 3 13 9 15 3 9 1 9 15 13
7 7 15 15 13 9 0 13
4 7 3 13 15
8 7 13 9 15 7 13 1 9
8 7 13 3 13 0 7 13 9
6 9 3 13 13 1 12
13 6 13 15 16 12 1 15 15 13 15 13 15 1
2 3 15
3 15 13 0
9 12 1 12 15 13 15 1 1 9
10 7 9 3 9 13 3 13 13 1 15
17 6 3 9 0 1 15 9 9 13 0 0 16 3 13 13 9 0
6 7 13 0 13 11 9
1 13
4 0 13 9 15
5 7 13 1 0 15
3 7 13 0
10 0 13 9 15 0 9 15 1 0 13
21 6 13 15 16 3 3 13 1 9 9 3 1 9 0 3 0 13 0 1 9 9
7 7 9 13 13 1 9 9
5 15 13 1 9 0
3 3 13 13
5 13 9 7 13 9
4 11 3 13 15
8 3 16 15 13 13 7 3 15
4 7 13 0 11
18 6 13 15 16 15 3 1 9 0 16 3 9 9 13 3 15 13 13
10 3 16 13 15 3 13 15 3 15 13
5 3 3 7 15 13
7 7 13 1 9 15 9 11
4 7 13 9 15
9 7 13 11 7 11 7 11 15 1
5 7 13 13 7 13
3 7 13 0
4 13 3 7 13
17 7 16 13 3 13 1 9 7 13 16 16 13 13 13 1 15 9
2 7 13
6 11 9 15 0 15 13
5 13 9 0 1 15
6 7 13 7 13 15 13
3 7 13 11
5 3 13 12 9 13
8 13 7 13 16 3 13 1 9
3 9 3 0
3 9 3 0
7 7 3 13 13 0 9 13
6 7 13 3 13 15 13
6 7 13 3 7 13 0
1 13
2 13 9
7 6 13 9 9 1 9 9
1 13
1 13
6 6 15 15 13 3 13
27 7 3 15 13 13 11 11 12 1 12 7 1 0 9 1 9 7 9 1 0 9 7 1 9 7 1 0
4 13 15 7 13
8 7 16 13 3 13 1 15 13
1 9
4 7 13 13 15
9 3 0 9 13 1 15 7 13 15
15 12 3 15 1 13 13 9 13 9 0 9 7 13 0 9
5 7 13 11 13 0
10 3 1 9 13 1 9 7 9 13 15
4 7 16 13 9
7 3 9 15 13 15 15 13
9 9 3 15 13 0 13 9 1 0
3 7 13 15
8 3 0 13 9 0 13 1 15
6 7 13 11 1 0 9
8 7 13 15 9 7 9 7 0
13 11 3 1 3 13 13 15 3 3 1 9 0 9
3 3 7 13
7 0 3 9 0 13 1 15
5 7 13 9 3 13
10 7 15 13 0 9 13 1 15 13 16
4 15 13 15 13
12 15 13 9 0 0 7 1 9 15 3 0 13
6 7 3 13 13 9 0
10 3 13 15 1 15 15 15 13 1 0
8 3 0 9 13 15 7 13 15
5 15 13 11 9 13
4 11 3 13 0
2 15 13
13 7 13 9 9 1 0 13 9 7 13 1 9 9
7 0 3 9 13 9 15 13
2 13 9
3 15 15 13
16 7 13 15 13 15 7 13 9 15 7 9 15 13 7 13 15
1 13
5 7 9 9 15 13
13 7 16 13 11 1 9 3 13 12 1 9 0 9
9 7 16 13 11 13 15 13 0 13
4 3 0 13 13
8 3 7 13 3 7 13 15 13
8 7 13 3 1 9 7 9 13
4 3 0 3 13
8 7 1 0 3 15 13 13 11
4 3 1 0 13
4 3 7 9 13
5 13 9 0 15 13
5 7 3 3 9 13
9 7 13 13 11 9 15 13 15 11
7 16 9 13 3 3 15 13
20 7 3 3 9 13 0 9 1 0 7 9 7 0 9 13 11 13 7 13 11
4 7 13 15 11
4 15 13 9 9
2 15 13
7 7 13 15 0 9 1 0
6 11 3 3 13 15 13
3 3 13 15
5 13 1 15 15 13
12 1 9 3 0 13 13 0 12 1 13 15 13
15 13 3 15 13 11 15 1 0 13 13 15 1 9 13 9
6 11 3 13 15 7 13
5 13 13 15 9 9
9 13 3 16 1 9 13 15 0 9
9 9 3 13 9 16 3 11 13 15
6 11 3 3 13 13 0
6 15 3 13 13 9 9
2 13 15
4 15 3 0 13
4 3 0 3 13
2 13 15
15 11 3 13 9 13 13 0 11 7 13 11 9 13 16 13
22 9 3 13 15 3 1 9 9 7 13 0 9 7 13 15 9 7 13 15 13 0 9
4 7 13 13 15
3 6 9 9
12 7 16 13 15 13 0 9 7 13 15 9 15
6 7 13 0 16 13 15
17 7 13 13 15 11 0 13 1 9 9 11 7 11 16 13 9 15
11 7 13 0 1 11 9 15 13 13 11 9
6 7 13 15 13 0 9
3 7 3 13
13 7 13 15 13 9 15 13 9 1 15 15 15 13
4 13 3 9 0
6 7 13 9 9 15 13
2 9 9
14 7 1 15 13 12 9 12 1 0 7 15 1 0 15
6 7 13 13 9 15 13
5 7 1 0 13 13
9 7 13 13 15 13 9 15 7 13
17 6 15 13 9 7 1 12 9 13 0 13 15 3 0 13 1 9
10 3 3 0 9 13 1 15 1 9 13
11 11 9 11 13 3 1 9 16 13 7 13
8 7 15 1 15 13 13 13 15
14 7 13 9 0 9 13 13 1 0 9 3 1 9 0
8 7 9 0 13 11 9 0 13
4 8 8 8 8
3 15 13 13
8 9 15 9 15 3 15 13 15
3 6 11 13
1 13
7 13 16 13 11 1 13 15
6 11 3 13 9 0 13
11 7 9 9 13 13 1 12 1 3 3 3
12 13 3 9 15 1 0 13 16 3 13 13 13
6 3 9 0 9 9 13
14 1 15 7 11 11 7 11 11 0 7 11 9 7 11
19 7 16 13 1 11 13 15 7 13 15 3 15 0 15 3 1 15 13 11
6 11 3 13 16 3 13
9 7 13 9 13 15 16 3 0 13
8 7 16 13 1 9 13 9 11
25 11 3 13 9 7 13 15 13 9 7 13 15 1 9 15 13 13 1 9 7 13 9 1 9 9
9 11 3 11 7 11 11 13 3 13
11 7 3 3 12 9 13 1 9 13 3 9
4 7 13 1 3
7 15 13 15 9 1 9 9
4 13 3 0 3
14 7 13 1 9 13 0 13 1 0 13 9 0 7 13
3 15 13 0
2 13 13
1 13
3 3 13 3
5 6 9 3 13 15
13 7 13 7 13 9 15 7 11 16 13 15 1 11
6 3 0 13 13 1 9
6 13 3 15 9 7 9
4 7 15 15 13
14 13 3 3 0 9 13 3 11 11 1 15 13 12 9
11 0 13 13 0 15 1 15 13 13 7 13
12 7 0 13 16 13 7 13 13 1 15 3 13
15 1 0 3 12 1 15 13 13 13 1 15 9 13 1 9
5 7 0 13 13 0
5 3 13 0 12 13
15 7 13 9 0 7 9 9 16 0 15 13 15 13 3 13
8 13 1 9 0 13 9 15 9
7 15 13 7 13 13 0 13
5 15 3 3 13 13
7 9 3 15 15 13 0 13
5 1 9 15 9 13
3 9 13 0
8 7 16 0 15 13 3 15 13
16 7 9 3 16 13 13 15 13 13 1 9 7 13 1 0 9
12 0 3 13 13 3 9 13 7 9 13 13 9
49 16 3 0 13 13 13 9 15 1 15 13 13 9 3 13 15 15 1 9 0 13 7 9 13 9 13 13 3 15 13 1 9 15 3 1 9 15 13 0 11 16 13 15 9 1 15 13 13 9
13 13 1 9 11 9 11 9 15 9 11 1 9 11
10 7 9 0 1 9 11 7 9 15 11
15 13 3 0 0 1 9 13 1 15 9 7 9 9 1 9
16 7 3 13 0 9 3 16 13 11 0 7 0 13 1 9 15
10 13 3 0 9 9 13 1 0 9 9
10 7 11 13 13 13 7 9 13 1 15
5 13 3 1 0 9
8 3 13 11 16 13 13 9 15
12 7 9 15 11 13 15 9 7 13 9 15 11
12 7 13 9 15 7 9 7 0 1 9 15 13
5 13 3 0 1 9
15 7 9 7 9 3 13 7 9 0 13 3 1 9 9 15
25 7 15 13 1 0 1 9 7 9 11 16 13 9 9 1 9 7 0 1 9 0 13 9 9 0
5 7 13 11 1 9
3 3 0 13
11 15 3 13 9 7 9 15 13 1 9 15
5 7 13 9 13 15
7 15 13 11 15 13 1 9
10 7 13 13 13 1 15 7 0 15 13
26 7 6 13 13 7 3 13 13 3 1 9 15 0 13 1 15 16 3 13 9 15 15 13 1 9 15
14 13 3 3 13 13 1 0 7 13 16 9 13 1 9
8 7 15 13 13 0 7 13 0
13 7 13 13 16 13 13 9 9 15 13 1 9 15
15 1 0 3 9 13 11 9 15 7 13 15 9 12 13 16
13 3 15 13 9 1 9 15 13 13 9 15 1 9
27 1 9 3 0 13 13 9 11 1 9 1 9 11 15 9 11 1 9 13 9 15 9 13 11 1 9 11
4 7 9 9 11
3 6 9 0
4 0 15 1 9
14 15 16 13 13 13 1 9 15 7 13 15 13 0 9
4 7 13 9 15
3 3 13 11
5 13 3 9 1 9
12 6 13 1 9 7 13 9 7 13 9 15 11
13 7 13 1 9 11 1 0 7 9 15 3 13 9
5 13 3 11 1 9
5 7 13 9 13 15
10 9 0 13 1 15 7 9 0 13 15
9 3 7 3 15 13 0 13 9 9
12 7 6 11 0 15 3 15 13 9 1 9 15
17 7 0 9 13 0 0 15 13 0 16 3 13 0 1 9 15 9
3 6 9 9
5 13 15 1 9 15
5 7 13 1 0 9
8 7 13 1 9 11 7 13 11
13 7 13 13 3 13 9 11 11 13 9 1 9 15
6 7 13 13 9 0 11
6 7 13 9 0 7 13
11 7 3 0 15 16 13 9 9 15 1 15
18 6 3 3 13 13 9 9 15 1 9 15 13 1 9 9 1 9 15
13 7 0 15 13 16 13 15 15 13 13 15 1 9
3 7 13 11
13 7 13 9 15 1 9 0 15 16 13 9 9 15
16 6 3 1 0 0 15 13 15 9 16 13 15 0 15 13 13
13 7 0 9 15 7 9 15 1 9 7 9 13 15
5 13 0 9 9 15
7 13 13 1 9 7 13 0
3 13 13 0
4 7 0 13 0
18 13 11 9 15 13 9 3 13 13 1 9 15 11 7 9 15 1 9
6 7 13 13 1 9 15
9 11 3 13 13 9 13 7 13 9
9 7 13 13 1 9 0 13 13 9
7 7 13 15 9 9 15 11
5 7 13 9 15 13
4 3 7 13 11
5 7 13 1 0 16
9 15 13 1 9 15 15 13 0 9
5 7 13 9 13 13
4 7 13 13 0
13 13 13 3 3 9 15 7 9 15 7 13 13 9
8 7 13 13 9 1 15 9 15
9 7 1 15 0 11 13 15 9 0
9 7 13 15 15 13 1 9 15 13
5 15 13 9 0 13
6 3 9 9 13 1 0
10 0 9 11 16 13 7 13 9 9 15
33 7 13 9 9 15 1 9 11 9 15 3 13 13 1 9 0 15 1 9 13 9 15 9 1 9 15 7 1 9 15 15 13 15
41 1 13 9 1 9 15 7 13 9 15 0 9 13 15 13 1 11 9 15 13 15 15 16 1 9 1 9 9 15 13 13 0 1 9 7 9 1 15 15 9 15
6 7 15 9 9 0 13
47 13 3 1 9 9 13 9 15 1 13 9 9 9 15 1 9 9 15 1 9 9 9 15 1 15 13 15 13 1 0 13 0 15 1 9 7 1 9 9 13 1 13 9 15 1 9 9
6 9 3 13 7 13 9
11 7 13 1 9 3 1 9 9 15 1 11
15 13 13 3 1 9 0 13 9 1 11 11 16 13 0 9
9 7 13 15 16 13 0 1 15 9
32 13 3 3 11 1 11 1 9 11 1 11 9 11 15 13 11 3 16 13 1 9 7 9 11 16 13 1 11 13 15 9 0
11 13 13 3 1 13 3 13 13 9 16 13
21 7 13 9 15 0 7 9 15 13 7 13 15 1 9 16 3 13 15 9 1 9
14 7 9 13 1 9 0 13 7 13 9 9 1 9 15
16 7 6 9 9 13 1 0 7 9 9 13 0 7 13 9 0
4 7 13 0 9
2 13 13
8 13 9 9 13 7 13 1 9
13 7 3 13 13 1 9 9 9 0 13 9 7 13
12 9 1 0 9 7 1 9 9 1 9 0 9
10 7 13 13 3 13 1 15 9 1 9
4 9 13 1 3
16 13 3 11 7 13 0 9 15 13 13 15 13 9 7 13 15
3 7 13 13
12 13 3 13 1 9 15 13 13 0 1 9 0
10 11 3 13 15 9 0 13 1 9 15
19 7 13 13 9 13 7 13 9 1 15 15 13 7 13 3 13 13 1 0
22 7 16 13 13 9 12 16 13 13 13 9 15 11 15 13 13 1 9 16 1 9 13
49 7 16 13 13 9 9 15 1 9 11 13 0 1 11 16 13 15 9 3 13 13 1 9 9 16 15 0 13 9 0 9 13 7 16 13 9 1 15 13 13 1 9 9 9 9 7 12 9 9
18 7 6 9 13 1 11 15 9 11 7 9 0 0 7 0 13 9 11
6 7 9 0 13 1 15
6 7 13 1 9 1 9
21 7 16 13 9 11 9 15 16 13 1 9 9 1 15 3 15 13 15 1 9 15
31 3 13 9 15 9 1 9 15 1 9 16 13 9 15 9 15 15 13 1 9 15 9 9 1 9 9 7 9 9 15 11
13 7 13 9 15 7 9 13 1 0 15 13 1 0
10 7 13 0 11 7 13 1 11 9 15
16 6 13 13 0 1 9 7 9 0 1 11 7 1 9 15 13
12 7 15 0 9 13 9 16 13 1 0 9 9
15 0 13 1 9 0 7 13 1 9 15 9 12 1 9 15
19 7 0 9 3 1 9 12 15 3 13 1 9 9 7 9 13 9 7 9
7 7 0 0 9 13 13 9
15 7 3 13 15 1 9 9 13 13 1 11 1 9 15 11
7 9 3 13 7 13 0 9
6 7 9 9 13 1 0
13 7 13 9 15 1 15 9 1 11 1 9 0 9
16 13 3 0 13 1 9 13 9 9 7 13 15 1 0 7 0
9 7 3 13 13 13 1 11 13 15
17 7 13 13 1 9 13 0 1 9 13 1 0 13 13 0 7 13
11 13 3 15 15 15 13 1 9 7 9 15
6 7 13 9 15 1 0
5 9 15 13 15 3
8 6 9 15 7 15 13 13 15
5 15 13 16 15 13
11 13 16 1 0 15 9 15 13 13 15 13
10 7 15 3 13 9 15 13 13 1 0
7 7 13 1 15 7 13 11
4 7 13 0 0
11 7 11 13 9 9 7 9 1 9 7 9
43 9 3 0 9 11 11 13 11 11 11 9 3 11 11 11 3 9 15 9 11 7 11 9 7 11 11 9 1 9 9 11 7 11 13 13 9 9 1 11 11 9 1 9
4 9 13 1 9
3 13 9 9
4 0 13 9 15
9 15 9 13 7 15 9 7 9 13
10 7 13 0 1 0 7 0 1 9 0
6 7 13 15 9 9 9
9 9 9 15 13 15 13 1 13 9
3 9 13 11
12 13 3 15 16 13 9 1 9 0 13 9 11
8 3 3 9 1 9 9 13 13
11 15 3 9 3 13 9 13 7 1 9 13
5 7 13 15 9 13
3 15 3 13
4 13 3 13 0
10 13 3 3 9 16 13 7 13 1 0
3 9 15 13
5 3 0 13 1 15
8 15 0 3 15 13 13 15 13
6 13 3 15 3 9 13
4 15 13 3 15
3 7 13 0
6 15 13 3 7 9 13
20 13 3 9 7 13 15 1 9 15 1 11 16 3 15 13 11 13 11 13 15
5 15 3 9 13 15
12 13 3 0 15 15 3 13 0 13 9 9 15
8 15 15 13 1 9 0 7 9
15 15 9 1 9 15 7 13 9 15 7 13 9 1 9 15
5 9 3 13 9 0
7 0 3 7 15 13 13 9
29 11 3 9 16 13 1 0 1 11 9 9 15 7 1 15 0 15 13 11 13 3 0 1 15 7 13 11 1 9
6 7 9 1 9 13 13
5 15 13 9 15 13
4 1 15 13 15
237 7 0 11 13 13 3 9 12 3 13 9 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 11 15 13 9
9 11 3 0 9 0 13 13 1 11
12 7 13 1 9 1 9 9 12 7 13 1 9
6 7 15 13 1 9 0
4 13 3 0 9
5 7 13 1 0 11
3 13 13 16
11 3 1 9 0 13 9 7 1 15 9 9
17 7 13 0 9 7 13 0 15 9 9 9 1 9 9 7 13 15
17 15 13 9 0 0 7 9 0 16 15 13 13 7 15 13 13 0
9 15 3 16 13 1 15 13 15 15
2 13 13
8 9 9 15 13 7 0 0 13
8 16 9 9 13 13 15 3 3
25 13 13 3 16 9 15 13 1 15 16 13 15 7 16 1 9 13 15 16 3 13 1 9 9 15
5 7 13 11 13 0
2 13 13
5 3 13 9 9 15
17 7 13 13 11 1 9 9 1 11 7 9 13 1 0 9 1 0
10 7 15 13 1 9 15 7 13 1 15
18 7 13 11 3 13 13 7 13 1 9 15 9 9 1 9 7 13 13
9 7 3 13 9 13 9 3 13 13
10 9 9 1 15 1 16 13 15 13 0
19 13 15 13 9 9 7 0 9 13 13 1 9 13 9 9 13 7 9 9
8 7 16 13 9 13 9 7 13
6 13 3 13 1 0 16
8 3 13 13 0 9 1 9 15
5 7 15 9 0 13
12 7 13 1 9 9 15 13 1 9 15 7 13
3 7 13 0
5 3 13 15 0 9
4 9 13 15 0
2 13 3
11 6 13 15 16 15 9 0 13 1 9 15
4 1 9 13 15
25 0 9 13 1 9 11 1 11 3 13 13 9 9 12 7 9 12 16 13 13 9 0 1 15 9
14 7 1 15 0 13 13 11 3 1 11 11 1 9 9
8 7 15 15 13 13 3 11 0
9 7 13 13 15 1 9 9 0 13
16 7 13 0 3 1 9 9 1 15 9 0 13 13 16 13 15
7 15 3 13 1 0 0 13
11 7 13 1 11 9 11 3 7 13 0 9
11 7 13 1 9 15 16 1 9 13 9 15
13 7 1 9 13 9 13 9 0 7 13 9 0 13
1 13
3 13 13 15
2 0 9
5 7 13 0 11 13
5 13 7 13 1 0
14 7 16 13 0 9 1 0 13 1 0 15 7 0 13
11 7 13 13 9 1 15 7 13 1 3 13
14 15 13 0 9 16 1 9 7 9 13 0 9 7 13
9 7 13 9 1 0 1 15 9 9
5 7 13 0 1 15
6 7 13 1 0 13 9
3 7 13 0
5 7 3 13 13 0
14 16 9 3 13 15 15 13 0 0 9 13 0 1 15
7 3 0 0 9 13 13 15
10 13 3 3 9 1 0 13 7 13 16
4 15 13 9 9
17 13 3 9 13 13 1 0 9 7 9 13 15 7 13 3 1 15
7 7 13 0 16 13 1 15
4 15 0 13 16
12 3 15 9 13 15 13 9 9 16 3 13 13
6 7 13 13 1 9 11
18 13 13 3 16 9 13 1 15 16 13 9 9 7 15 13 1 9 11
7 7 13 12 9 13 1 9
6 9 3 13 7 13 9
7 3 13 3 13 13 1 11
9 13 1 0 7 13 9 15 1 9
5 7 13 11 13 0
7 9 1 0 9 13 15 13
6 1 9 3 15 13 9
8 7 16 0 13 13 9 9 0
4 13 3 9 15
9 7 13 7 13 0 9 3 16 13
8 13 1 15 16 9 9 13 9
26 9 3 13 15 7 15 15 1 0 13 1 9 9 15 13 3 3 11 7 11 9 11 15 13 9 11
5 7 13 1 11 11
2 13 13
6 1 0 3 9 13 13
10 7 13 1 9 9 13 15 13 13 0
6 9 16 13 13 15 13
6 7 13 9 13 0 13
1 13
6 7 3 9 13 1 0
7 7 15 13 0 16 15 13
16 7 13 13 15 9 7 13 1 9 15 3 13 11 1 9 0
6 13 3 3 9 1 0
7 15 3 13 1 9 7 13
6 7 13 13 1 12 9
4 7 15 13 13
7 7 9 13 9 1 13 15
10 7 6 9 13 1 9 9 15 13 9
8 7 13 15 13 7 13 1 15
12 7 3 13 15 9 0 13 1 9 13 1 9
5 15 9 3 13 13
5 9 13 15 9 15
7 7 13 13 9 7 9 13
6 15 13 0 15 13 9
10 3 13 3 11 9 15 13 13 1 0
5 15 13 1 9 15
12 15 13 0 13 13 15 9 7 13 13 7 13
2 13 9
2 15 13
1 13
8 13 9 15 7 13 1 9 15
9 7 3 13 1 0 13 1 15 13
7 7 9 13 15 7 13 9
6 7 13 13 9 13 16
15 7 1 0 13 7 13 9 9 11 13 1 9 7 13 0
2 13 15
7 7 13 15 13 13 13 15
9 7 13 15 9 0 11 1 9 15
12 7 13 9 0 9 7 15 15 1 0 13 13
10 7 13 9 7 9 15 13 1 9 15
6 7 13 11 13 1 0
8 3 13 13 0 7 9 1 9
5 3 0 13 1 15
16 3 9 11 13 3 7 9 13 3 3 9 15 3 13 7 13
3 15 15 13
11 3 13 9 9 16 1 0 13 9 13 13
10 13 3 9 7 16 13 13 1 0 9
5 3 13 1 0 9
11 3 3 0 13 7 0 3 13 9 1 0
8 7 15 13 9 0 1 9 0
11 3 13 9 0 9 7 15 13 7 9 13
11 7 9 0 1 9 0 13 13 7 15 13
7 7 15 13 0 3 13 0
2 13 3
3 0 0 13
18 13 13 3 1 9 0 16 13 1 9 13 9 15 9 7 13 13 9
7 15 13 15 3 13 1 9
6 7 13 11 1 15 13
14 3 0 13 15 13 11 16 13 15 7 15 1 15 13
25 3 13 1 9 9 7 9 9 13 7 13 7 13 0 15 1 15 13 15 3 13 13 3 3 9
4 7 13 0 16
6 9 13 9 9 3 9
13 13 13 3 3 1 15 9 16 13 1 9 7 13
10 7 13 3 9 7 9 15 0 13 0
7 7 13 9 15 13 9 0
5 13 7 13 1 0
3 7 13 13
5 13 3 1 0 11
14 13 15 16 13 9 3 13 7 3 9 0 13 7 13
5 7 13 15 13 9
3 13 9 15
5 7 13 13 9 15
16 13 13 3 1 0 9 13 1 9 13 7 13 13 1 9 9
8 7 16 9 13 13 13 9 15
41 7 13 12 1 15 15 3 9 13 11 15 13 11 7 11 9 15 11 7 11 11 7 11 11 7 11 11 11 7 11 15 13 11 11 11 7 11 11 15 13 9
8 7 13 1 0 13 1 9 0
28 7 9 9 15 7 9 0 9 1 15 11 7 11 7 0 11 7 11 15 13 16 13 15 7 13 1 9 15
7 7 15 13 1 9 0 13
8 7 15 13 9 1 9 15 13
7 0 0 16 15 13 9 9
6 0 15 3 13 16 13
21 0 13 16 15 13 9 7 16 13 15 7 13 7 13 9 15 3 0 1 9 9
6 13 1 0 9 7 13
7 6 3 9 15 0 1 9
7 1 0 3 13 9 9 15
7 6 15 15 13 13 16 13
9 6 15 15 13 3 16 13 7 13
7 6 16 3 15 13 15 9
5 7 15 13 15 13
3 13 9 15
5 13 0 15 15 13
3 13 13 15
9 15 15 15 13 1 9 13 3 0
11 7 1 15 15 13 15 9 3 9 13 13
13 15 3 13 15 13 7 15 13 15 15 13 3 13
12 7 3 13 16 13 15 9 3 15 13 0 3
6 3 3 9 13 15 13
16 7 16 13 0 15 15 13 15 15 13 9 16 3 9 0 13
13 7 16 0 13 0 1 15 13 13 15 9 13 15
11 3 13 9 15 7 13 7 0 13 15 13
17 7 13 9 15 0 7 13 9 0 16 15 0 13 1 0 7 0
9 13 3 0 3 3 9 15 0 13
5 13 13 7 3 13
5 13 13 7 3 13
4 13 7 13 15
11 9 0 0 7 13 7 13 13 1 9 15
5 13 3 0 3 9
5 3 13 0 0 13
5 3 0 1 9 13
5 3 13 9 1 9
7 0 3 15 13 3 9 15
8 15 3 13 9 1 9 9 15
20 7 3 13 13 9 15 9 13 13 9 1 9 15 0 1 9 15 9 3 13
16 3 13 3 9 0 15 13 9 0 3 7 9 0 13 9 0
7 15 3 9 1 9 15 13
7 3 7 3 1 9 13 9
6 3 7 1 9 13 9
9 0 9 1 0 9 9 15 13 0
7 7 0 9 1 0 13 0
6 1 9 3 9 9 13
14 0 13 9 13 9 15 13 1 0 7 13 9 1 9
13 9 3 13 13 13 9 9 0 7 3 13 15 13
5 13 3 13 1 9
16 15 3 13 7 3 13 0 13 9 13 9 15 1 9 1 9
8 1 15 13 13 9 7 3 13
7 7 13 13 9 9 0 0
11 16 3 13 15 9 15 1 9 9 13 11
8 9 3 15 9 3 13 13 13
18 7 16 13 1 11 13 1 15 0 9 13 15 16 13 7 13 9 15
12 3 0 16 13 1 11 13 15 3 13 15 16
6 0 13 16 0 0 13
9 13 3 9 15 7 9 15 13 15
5 11 3 13 1 0
14 7 16 3 3 3 13 1 9 13 1 15 9 9 13
3 9 13 13
9 3 3 0 13 16 1 9 15 13
12 3 3 15 9 13 1 9 13 13 1 15 9
6 7 13 0 13 7 13
5 7 15 13 7 13
7 7 9 15 13 0 7 13
11 15 13 11 13 13 7 13 13 15 9 13
3 6 13 15
6 3 1 11 0 9 13
4 7 13 13 3
9 7 13 1 0 9 15 7 9 0
13 16 3 13 9 9 7 6 13 13 9 0 9 15
4 7 0 9 13
6 7 9 9 0 1 0
10 15 16 13 9 9 13 1 15 13 0
2 13 13
5 0 3 15 13 13
2 7 13
1 13
8 7 13 15 13 13 7 13 13
5 7 13 0 9 15
20 13 3 15 9 7 13 9 13 16 9 0 13 1 15 7 16 9 13 9 15
13 7 13 0 9 1 0 11 1 15 7 15 3 9
12 7 13 12 1 9 15 11 7 13 1 9 13
8 15 13 15 13 13 7 15 13
7 16 3 13 1 15 9 13
8 15 13 15 13 13 7 15 13
18 1 0 3 9 13 0 1 9 7 9 7 9 0 7 0 0 13 9
4 7 13 13 0
20 13 13 11 15 13 7 13 16 0 13 0 13 0 13 0 13 0 13 0 13
11 7 16 13 9 11 13 13 1 11 1 9
5 15 13 1 9 13
3 9 9 13
4 7 15 13 13
12 6 15 1 9 0 13 7 9 1 9 9 13
4 7 15 13 13
1 9
4 3 0 3 9
6 0 13 1 15 13 13
13 6 13 9 15 1 9 15 15 13 9 15 1 15
3 13 3 15
9 0 1 13 9 9 11 9 15 13
11 7 15 9 13 3 9 13 9 13 9 11
16 9 3 7 9 0 9 9 13 1 15 3 0 3 13 1 15
12 0 13 9 13 1 9 7 13 1 3 7 13
6 13 15 9 7 3 13
4 13 7 3 13
14 13 3 11 9 3 7 13 9 3 7 13 9 7 13
2 9 13
8 13 9 9 13 7 13 7 13
8 7 13 13 9 1 15 9 15
5 7 13 9 9 13
18 7 6 9 15 13 1 9 9 3 13 16 13 1 9 9 13 9 9
23 7 13 3 1 9 15 9 13 13 9 15 7 9 9 15 13 7 13 9 15 7 9 13
10 13 3 9 15 13 15 13 1 15 13
16 0 16 13 9 13 3 15 7 15 9 15 13 15 16 9 13
6 7 13 11 13 1 0
5 11 13 15 15 13
5 12 9 13 15 9
6 12 13 9 12 15 12
7 3 13 0 3 13 13 15
5 15 3 15 3 13
3 13 11 13
6 13 16 15 15 0 13
4 3 0 13 15
2 3 13
3 13 0 9
4 13 1 9 15
5 9 9 15 3 13
10 0 3 9 13 9 15 7 9 15 13
4 9 15 3 13
10 0 3 16 15 13 3 13 13 9 15
5 9 9 15 3 13
6 0 3 9 13 9 15
6 15 3 0 13 3 13
4 13 3 1 0
3 13 15 9
8 7 13 15 3 13 13 1 15
7 15 13 0 15 3 9 13
4 13 3 1 9
5 9 15 15 0 13
4 7 13 13 3
14 16 3 9 0 13 7 1 9 13 1 15 13 1 9
6 13 15 13 13 9 15
15 7 16 13 15 13 1 9 7 13 13 7 9 9 13 0
5 7 15 13 1 9
7 7 13 13 16 3 13 9
11 7 15 13 1 9 7 3 13 9 13 0
5 7 13 13 9 0
3 0 13 13
9 13 3 15 9 15 15 13 0 9
3 15 15 13
7 15 13 13 13 9 9 9
12 0 3 1 9 16 13 3 13 7 13 3 13
4 13 3 0 9
7 15 3 1 9 13 15 13
13 3 13 9 7 13 9 1 9 15 16 13 0 13
11 3 15 1 9 15 16 13 1 9 13 9
9 15 1 9 13 7 1 9 9 13
23 15 3 1 9 13 0 13 15 13 7 1 9 7 9 7 9 9 13 13 7 3 13 9
21 15 3 1 0 9 0 13 15 1 9 0 7 0 13 9 13 7 9 13 1 9
19 15 3 9 13 13 15 9 7 1 9 13 7 1 9 13 16 13 13 9
4 13 3 3 13
17 15 3 13 13 0 7 15 3 13 3 15 13 15 13 13 1 0
16 13 3 1 0 9 7 9 15 7 3 13 13 1 15 1 9
4 7 13 13 0
5 15 13 13 1 15
13 9 15 7 9 15 0 13 15 9 9 13 7 13
6 13 13 3 1 12 9
3 13 1 9
2 7 13
14 13 3 0 13 7 13 9 9 1 9 7 13 7 13
5 13 3 13 15 13
2 9 13
4 7 13 13 9
3 13 3 0
7 15 13 13 13 13 1 3
13 15 13 0 13 16 7 9 13 7 9 7 13 15
9 13 3 1 9 9 15 13 1 11
28 7 16 13 13 1 9 13 0 9 15 15 13 9 3 9 0 7 9 3 13 3 7 1 9 13 7 1 9
7 15 3 13 11 13 1 0
5 7 13 9 0 13
2 13 15
8 13 3 9 0 16 13 1 9
11 0 3 9 13 0 7 13 9 7 9 13
8 7 13 9 13 1 9 1 9
5 13 3 0 11 13
4 15 15 9 13
10 3 0 13 11 16 13 9 0 1 15
10 7 13 0 16 13 0 16 1 9 13
3 7 13 0
9 13 3 9 1 9 7 13 1 9
11 7 9 13 9 1 9 1 9 7 13 13
14 15 3 13 13 15 13 13 7 13 1 9 7 1 9
27 13 3 13 15 13 13 7 13 1 11 7 13 9 13 1 15 9 13 13 7 0 9 1 9 15 7 13
12 13 3 0 3 15 13 3 0 13 13 1 11
15 7 13 0 15 9 9 9 16 13 1 15 16 9 0 13
6 15 3 13 9 13 13
5 13 3 15 11 13
9 13 9 15 7 13 15 15 13 9
10 7 13 1 0 9 13 15 0 13 11
9 13 13 3 16 13 11 13 0 9
5 13 3 15 13 15
12 7 6 13 9 15 9 11 7 15 9 9 13
23 7 13 1 9 11 13 15 16 13 1 9 15 16 9 0 13 0 3 9 12 7 0 13
7 7 13 16 13 1 9 13
6 7 3 13 9 9 15
3 7 13 11
5 15 13 15 15 13
10 13 3 15 13 11 7 15 1 0 13
8 9 9 15 13 7 13 7 13
3 15 15 13
3 7 13 11
7 3 15 13 9 1 15 13
4 3 15 13 0
6 9 9 15 15 0 13
3 13 1 9
10 3 0 13 13 1 9 9 13 15 16
4 13 13 9 15
3 13 13 0
2 13 13
5 13 3 7 0 13
6 13 3 15 7 13 0
3 3 0 13
2 13 13
5 3 13 13 7 13
7 7 13 15 13 16 13 13
2 9 13
8 7 13 13 9 15 7 13 3
5 7 13 0 13 13
16 13 3 12 9 13 0 9 7 9 1 15 9 3 16 9 13
9 7 13 0 13 9 9 7 13 0
4 7 13 1 0
4 15 13 1 9
11 7 1 15 9 13 3 13 7 3 3 13
18 7 15 3 13 15 13 1 9 0 3 9 9 15 13 1 9 1 0
9 13 3 13 1 9 13 7 13 3
36 13 3 11 9 15 15 13 1 15 7 13 3 16 13 1 15 16 11 13 1 0 1 15 3 16 11 13 1 15 3 16 9 12 1 0 13
3 11 15 13
9 15 3 13 0 1 15 13 15 0
4 7 13 13 15
11 7 13 0 13 3 1 9 0 15 13 11
7 15 16 13 9 13 13 0
15 7 13 0 7 13 0 1 9 9 7 15 15 9 13 13
9 9 3 13 13 7 13 12 13 0
21 13 9 16 13 1 9 9 7 15 3 13 13 7 13 9 16 3 1 9 0 13
4 15 13 0 13
3 3 0 13
6 13 3 3 9 12 12
5 13 3 1 9 15
6 13 0 13 1 9 0
3 7 3 13
4 7 13 13 15
13 13 3 12 9 7 12 9 13 1 9 7 13 0
6 7 13 15 7 13 13
12 7 13 13 16 0 13 13 13 1 0 3 9
4 7 13 0 13
5 15 15 13 13 9
5 3 0 13 7 13
12 11 9 15 3 11 15 16 9 12 1 0 13
3 13 3 0
6 15 3 15 15 13 13
11 3 0 13 0 13 16 15 13 0 13 16
20 13 9 9 0 13 7 13 1 0 7 9 9 7 9 7 13 7 0 9 13
4 13 3 1 15
17 16 15 13 1 15 13 13 15 15 7 13 9 15 3 7 13 15
9 15 3 13 9 15 0 13 13 0
10 3 15 13 9 15 1 15 0 13 0
16 15 3 13 9 16 13 0 9 15 3 0 13 7 9 15 13
21 3 15 15 13 7 15 9 0 9 9 13 16 13 1 9 15 7 9 7 0 9
12 13 15 3 13 15 3 13 9 16 13 9 9
22 13 13 3 1 0 9 3 9 12 7 13 11 7 11 7 11 7 13 1 9 16 13
14 7 13 13 16 13 9 9 15 0 7 9 15 0 13
7 7 6 12 9 13 1 0
17 13 3 11 7 11 13 1 9 7 13 9 15 15 13 13 1 11
9 11 3 7 15 1 0 13 13 9
12 7 13 13 9 15 7 12 9 15 13 1 0
32 7 13 13 16 13 1 0 13 11 1 11 9 0 13 15 3 13 7 13 12 9 12 15 7 12 11 7 12 11 13 15 13
7 7 9 13 13 1 9 13
5 0 13 9 15 13
2 15 13
8 7 16 13 9 13 13 11 0
14 7 15 13 7 15 13 1 0 9 15 1 0 15 13
14 13 13 3 1 13 9 13 0 1 9 13 0 9 0
7 7 6 9 1 9 13 13
8 13 1 9 15 16 0 13 15
10 7 13 9 15 16 13 0 7 3 13
4 13 3 11 13
12 6 9 0 7 0 3 13 1 15 7 13 15
4 13 3 9 15
8 7 16 13 13 0 9 7 13
13 7 13 11 9 0 7 13 9 7 13 0 9 15
11 15 7 13 1 15 15 13 13 1 9 15
7 13 15 1 9 15 9 0
14 3 0 13 9 0 7 13 13 1 15 16 3 13 0
7 7 13 13 15 1 0 9
9 13 3 9 1 15 15 15 0 13
15 3 11 13 9 9 0 13 9 13 15 1 15 7 13 0
9 15 13 9 0 1 9 15 15 13
10 3 15 0 13 1 15 15 0 0 13
4 13 3 11 13
16 9 13 15 1 9 15 13 9 7 13 15 16 3 13 15 1
2 13 13
9 15 3 3 13 1 15 1 15 13
16 13 13 3 16 13 9 9 15 7 15 9 15 13 16 13 11
6 7 13 9 1 9 15
10 7 3 13 15 16 9 15 13 13 11
9 16 13 3 9 15 11 7 11 13
11 9 13 13 16 9 13 1 9 7 13 0
4 7 13 13 0
11 13 13 3 13 0 1 9 13 15 1 0
4 13 15 3 13
4 7 13 0 11
8 9 3 9 3 13 3 9 13
4 13 3 1 0
2 13 15
3 0 3 13
8 9 13 15 3 13 13 9 15
6 13 16 0 13 0 15
3 15 3 13
3 7 13 0
12 13 15 9 7 3 13 15 13 0 15 3 13
4 13 1 0 11
13 15 13 9 15 1 9 7 13 3 0 13 9 9
8 1 0 3 13 9 3 15 12
16 7 13 0 0 1 9 15 1 15 9 7 9 3 13 0 13
3 9 3 0
9 13 3 9 9 16 13 9 1 9
1 13
8 6 15 13 15 3 9 1 9
14 13 13 9 3 7 9 3 7 9 7 15 1 9 13
6 1 15 9 13 3 13
3 9 0 9
11 7 16 3 13 9 9 13 1 0 9 15
6 0 3 13 9 9 15
6 13 13 1 9 1 9
12 7 1 15 9 13 7 13 15 13 15 13 15
10 7 13 0 15 1 0 13 7 13 0
5 13 1 15 9 9
13 1 15 9 13 7 3 13 15 13 1 9 15 13
11 3 9 15 13 15 1 9 15 13 1 15
7 3 0 13 16 13 9 9
6 6 15 11 6 15 11
21 3 16 1 11 7 11 13 13 9 15 1 15 13 13 3 1 9 7 9 13 13
10 3 11 7 11 3 13 1 9 3 15
11 7 15 11 3 1 9 13 3 1 9 13
5 15 15 13 15 13
6 7 15 15 13 15 13
9 15 3 15 13 13 15 15 15 13
7 13 13 3 12 1 9 13
7 13 11 3 9 1 9 13
14 6 13 15 9 13 1 9 7 9 7 1 15 9 9
4 7 15 15 13
9 3 1 0 13 13 16 9 15 13
9 13 3 16 9 15 13 13 1 9
8 1 0 9 13 9 0 7 13
18 13 15 9 9 9 7 9 16 13 0 1 0 7 0 7 13 15 0
7 15 15 13 13 1 9 15
6 7 13 1 9 15 13
6 0 9 15 13 15 13
23 13 3 15 16 0 9 7 9 13 13 15 15 13 7 3 13 7 13 15 13 7 3 13
10 7 6 15 9 0 13 13 0 7 13
6 9 15 13 9 0 13
5 3 0 13 1 15
2 3 13
3 0 13 13
3 13 7 0
2 3 13
4 0 13 7 13
9 0 3 13 13 15 0 13 1 11
5 7 15 13 15 0
15 9 15 13 1 11 1 11 7 13 1 9 15 3 13 15
6 7 9 13 13 0 13
8 13 3 16 9 15 13 0 9
11 3 3 9 16 13 1 9 7 13 15 13
8 9 3 15 9 13 13 1 15
6 7 13 15 9 13 13
9 7 13 13 9 15 13 9 7 9
11 7 0 9 13 12 9 7 13 9 7 13
3 9 0 13
8 7 15 13 15 16 13 13 15
12 15 0 12 13 15 0 13 0 15 13 1 9
5 15 13 9 1 0
4 7 13 0 11
5 13 7 15 13 3
25 7 9 15 11 9 13 0 1 9 15 7 0 13 9 9 11 15 3 13 1 9 9 13 9 0
6 11 3 13 1 0 9
4 15 13 7 13
12 9 3 13 15 9 16 9 15 13 15 0 13
6 13 3 0 16 15 13
8 11 11 0 13 7 13 1 0
4 3 12 13 0
18 7 13 13 16 13 1 9 15 13 3 13 13 12 1 9 15 1 15
10 9 13 15 13 3 3 11 13 9 15
3 7 13 0
3 16 13 13
4 9 13 9 15
3 13 9 15
12 7 13 15 9 15 16 3 0 13 15 13 15
4 7 13 1 0
13 15 15 13 9 7 13 1 0 0 9 7 13 0
20 9 13 15 12 9 16 9 15 13 1 9 1 15 7 3 13 15 13 1 0
6 7 0 1 3 13 13
4 13 15 0 13
12 3 9 13 13 7 9 15 15 1 13 1 9
6 3 13 13 7 13 15
4 7 15 15 13
4 13 7 13 15
3 13 7 13
4 13 7 13 15
5 15 3 15 13 13
4 7 15 13 13
3 7 13 13
11 15 3 1 15 9 13 9 3 9 13 0
8 7 16 13 9 3 13 0 9
23 16 3 15 16 13 0 13 0 9 13 9 15 3 3 9 15 1 9 13 9 0 13 15
8 7 13 13 9 7 0 13 0
11 7 16 13 9 13 13 0 7 13 13 9
5 15 3 1 15 13
6 1 11 9 9 13 9
9 7 15 13 9 1 9 13 1 15
8 15 3 16 13 9 15 13 15
7 3 13 1 11 13 15 9
12 16 3 15 1 11 13 9 9 15 1 15 13
5 3 15 9 15 13
13 3 16 1 9 9 13 9 3 13 1 15 9 9
12 16 0 13 13 9 15 1 9 13 15 15 13
18 16 3 0 0 13 13 15 0 9 15 13 1 15 13 7 9 15 13
8 15 3 13 15 1 1 15 13
12 16 0 9 13 1 9 13 1 9 0 13 9
6 13 1 9 15 3 13
6 7 16 13 13 9 13
14 7 3 13 7 13 12 15 9 0 15 7 13 13 3
7 7 13 0 9 0 0 0
14 13 13 3 16 0 13 13 9 15 9 1 9 13 0
9 0 9 15 15 13 7 9 15 13
8 3 0 15 13 9 9 7 13
5 9 3 13 13 13
10 9 13 7 9 3 13 0 3 9 11
13 3 3 11 13 9 9 3 13 3 9 9 9 0
12 9 9 13 1 9 1 9 9 0 7 13 0
13 3 13 1 9 9 13 9 11 7 6 0 11 3
11 9 9 13 1 9 1 9 0 7 13 0
19 15 9 13 7 1 0 13 3 7 1 9 7 1 9 16 15 13 9 13
6 9 9 15 13 9 15
10 16 9 15 13 0 0 9 15 0 13
10 13 3 16 9 15 1 15 13 9 13
21 16 3 9 15 0 0 13 3 13 15 9 9 13 0 0 7 3 9 9 13 15
11 7 16 13 13 0 15 9 16 13 1 15
3 7 13 13
5 7 13 9 1 0
11 3 15 9 15 1 3 13 9 7 9 13
10 15 3 3 13 15 0 13 9 7 9
15 0 3 15 13 15 1 3 13 3 15 15 1 3 13 13
6 7 6 15 0 13 15
18 7 6 15 9 16 13 9 7 9 7 15 9 7 13 9 7 9 9
8 0 3 13 13 7 0 3 13
14 6 15 16 13 3 9 15 3 13 7 9 13 3 13
8 13 3 15 1 9 0 13 0
7 9 0 13 3 15 9 13
3 3 0 13
21 3 15 9 0 6 16 13 9 9 15 13 3 13 7 0 12 9 15 3 13 9
5 9 3 15 13 0
17 3 13 16 13 9 9 15 16 3 15 15 13 15 3 13 15 9
39 13 1 0 9 7 9 7 1 0 13 7 13 16 13 9 15 9 15 13 13 1 9 9 1 9 0 1 9 11 3 1 9 11 15 13 1 9 7 9
3 3 13 15
4 13 1 0 9
8 6 15 9 0 16 13 9 9
8 0 3 13 7 15 15 13 13
29 16 0 1 0 13 13 9 7 9 0 3 13 7 9 15 13 1 0 13 7 13 13 15 1 9 15 16 13 15
7 13 1 9 9 15 13 9
19 3 15 1 9 13 1 9 13 7 15 1 9 13 13 1 9 13 1 9
5 13 3 15 9 15
15 3 13 1 0 15 13 9 7 1 0 3 13 0 15 13
5 13 3 15 15 13
10 13 15 15 16 13 13 9 13 1 9
3 3 13 15
2 0 13
3 13 3 13
4 0 9 0 13
3 13 3 15
17 15 15 13 13 1 15 1 9 3 9 9 13 1 0 1 9 9
10 15 3 13 15 1 9 13 1 9 9
10 7 15 15 13 9 1 9 9 13 0
9 15 3 15 1 9 0 13 3 13
21 16 3 13 15 1 9 7 1 9 7 9 13 0 13 3 7 15 13 7 15 13
6 13 3 15 15 1 9
9 9 13 9 15 16 13 15 1 9
4 3 0 13 15
9 9 15 15 13 9 7 9 1 15
4 13 7 1 0
18 13 7 13 1 15 9 16 3 1 9 15 9 15 13 1 0 15 13
6 13 3 9 1 0 13
7 9 15 0 0 9 9 13
2 7 13
2 0 13
6 13 9 15 7 0 13
15 7 3 13 15 15 13 13 15 7 0 15 7 13 9 15
8 9 13 0 0 13 1 9 0
1 13
1 13
1 13
8 0 0 9 9 15 13 1 15
5 15 3 13 15 13
11 3 13 15 15 13 7 3 13 1 9 0
5 13 7 1 9 15
3 3 13 15
11 13 0 13 9 15 13 3 7 9 15 13
19 13 9 16 3 13 3 7 13 15 3 13 9 3 7 9 7 9 13 0
6 3 3 15 0 13 0
12 16 3 3 15 0 13 13 15 1 0 0 13
4 13 9 3 13
2 3 13
2 3 13
3 13 3 15
21 16 3 9 15 3 1 9 13 7 3 1 9 13 9 3 13 3 3 15 0 9
9 7 15 13 13 15 13 7 15 13
5 7 13 1 3 13
7 9 3 15 13 16 0 13
9 3 13 9 9 7 0 15 13 15
4 13 13 0 9
7 3 13 9 15 13 15 9
19 13 15 9 15 3 13 9 3 13 1 9 3 9 3 13 3 7 9 13
10 3 3 9 15 13 3 3 9 15 13
26 13 9 15 13 7 9 13 7 15 0 9 13 9 15 3 13 1 9 16 16 13 7 13 3 13 15
9 0 9 0 15 16 13 9 13 13
19 7 16 13 1 0 9 7 16 1 0 9 13 7 3 13 0 13 9 0
20 0 3 13 16 16 13 9 9 15 9 9 13 13 3 7 3 13 13 9 15
12 3 15 13 13 16 15 9 3 13 9 9 13
10 9 1 15 13 0 9 7 3 1 15
3 13 3 9
20 15 13 13 0 9 7 0 15 13 9 1 9 15 16 13 0 1 9 9 9
10 0 0 9 15 16 13 9 13 3 13
10 3 13 15 16 1 15 15 13 13 0
19 0 3 9 15 13 9 9 15 7 3 13 7 3 13 1 9 15 13 0
10 15 3 3 13 7 13 0 9 13 0
8 7 15 13 0 0 13 1 15
10 9 13 13 1 9 7 15 13 16 13
10 9 3 13 13 7 3 13 3 16 13
7 13 16 9 13 13 1 9
3 3 13 15
2 7 9
25 13 9 1 9 7 9 1 9 15 9 1 9 7 9 1 9 9 1 9 15 7 9 1 9 15
8 16 13 9 13 1 9 3 13
2 9 13
3 7 3 13
10 7 16 9 13 13 16 9 13 7 13
7 9 9 9 7 9 13 13
6 0 3 9 3 3 13
11 15 3 3 1 15 15 3 13 15 0 13
8 3 13 3 16 3 0 9 13
17 13 3 15 0 1 9 13 0 1 9 15 9 11 13 1 9 15
4 7 13 13 0
13 13 16 0 9 1 15 9 9 13 16 0 13 13
3 3 13 15
7 7 16 9 13 15 3 13
26 3 0 12 7 12 1 15 13 9 1 11 7 13 15 13 16 7 15 9 13 1 15 9 13 1 11
3 3 13 15
4 13 3 0 9
17 9 9 13 15 13 1 9 15 7 13 13 9 1 0 7 3 13
5 13 3 1 9 9
15 6 9 12 13 16 15 13 13 9 1 9 0 7 3 13
3 13 3 0
5 3 15 3 9 13
5 3 0 13 13 0
14 9 13 0 3 0 9 3 16 13 1 0 7 13 9
7 13 3 13 1 9 15 9
11 7 6 9 15 13 9 9 9 12 7 12
9 7 13 13 3 7 3 13 3 13
10 15 16 13 11 13 1 15 7 13 0
6 9 13 13 1 9 15
11 7 13 0 9 7 3 13 13 7 13 9
10 13 3 9 13 16 9 13 11 13 9
11 1 0 3 13 7 13 7 3 1 9 9
15 9 15 15 9 3 13 9 15 7 9 1 9 7 13 13
20 0 3 9 11 15 13 11 6 12 7 12 9 3 13 13 1 9 0 9 9
8 7 16 0 13 13 15 0 15
11 7 15 9 13 1 0 15 3 13 1 15
2 13 3
11 15 0 13 9 9 7 15 0 13 13 0
15 7 13 7 13 13 1 9 0 7 9 9 13 1 9 15
3 7 3 13
14 0 13 9 15 13 9 13 1 9 9 12 16 13 0
12 7 13 1 9 7 9 13 7 9 13 1 11
4 13 3 0 15
6 9 3 0 13 15 13
5 15 3 13 1 0
16 16 3 13 9 9 7 13 9 7 13 3 13 7 13 9 13
3 9 13 15
4 7 13 13 15
3 3 13 13
10 13 1 15 7 13 7 1 9 15 13
3 7 13 15
4 13 15 3 13
23 3 13 9 7 9 9 16 13 11 7 11 7 11 7 15 9 1 9 9 15 3 13 3
15 7 13 1 9 7 9 7 9 7 9 7 13 1 9 9
13 7 6 13 0 15 13 0 7 13 0 15 13 0
8 1 0 9 13 15 9 13 0
3 7 13 0
1 13
3 13 9 0
16 3 13 15 3 7 3 7 0 13 16 3 13 9 13 1 11
25 11 11 15 13 9 7 13 15 15 13 1 15 3 13 13 9 15 3 9 9 15 1 9 7 13
5 6 13 15 9 15
11 13 3 15 16 3 13 15 16 13 16 13
6 0 15 13 1 9 9
8 7 6 9 15 0 13 1 0
11 7 13 11 13 1 9 0 7 9 13 16
3 3 0 13
7 15 3 13 13 15 7 13
5 7 13 1 0 13
15 15 15 9 7 9 1 9 13 7 3 3 13 0 9 9
7 7 3 13 1 0 13 0
14 13 3 3 1 13 9 13 3 0 9 13 13 1 0
10 7 13 15 15 15 7 0 13 13 15
8 7 3 13 1 9 0 9 13
17 7 16 13 13 13 13 1 0 9 16 16 13 15 15 13 13 15
3 9 13 0
7 3 13 15 9 1 3 13
6 3 15 15 15 13 13
5 7 15 15 13 13
7 13 3 3 15 15 15 13
9 0 16 13 15 1 3 13 13 0
7 0 15 13 9 1 9 9
4 3 15 13 15
8 9 15 13 9 0 7 13 0
15 7 13 9 15 9 9 13 13 16 13 16 3 13 13 15
5 7 13 3 15 13
3 0 13 15
9 9 13 7 3 13 13 7 13 0
3 13 15 13
3 7 0 13
8 9 9 13 12 7 13 13 0
2 13 15
3 13 15 13
3 7 15 13
7 9 13 7 3 3 13 13
7 7 13 9 13 0 9 15
10 7 0 7 0 7 0 7 0 13 3
3 7 13 9
9 9 13 13 3 13 7 3 9 13
4 7 13 9 9
5 13 1 9 7 9
7 7 13 13 16 13 9 15
13 13 3 15 16 15 9 0 15 13 13 13 9 15
5 7 13 13 1 0
15 7 15 3 13 9 15 7 13 1 15 3 13 13 15 9
35 15 3 1 15 13 9 13 3 3 13 13 9 15 0 13 16 13 1 13 16 16 13 9 7 3 13 13 15 15 13 13 13 15 13 16
8 0 9 13 13 7 3 13 13
27 7 15 9 13 13 9 1 15 9 3 13 3 13 16 13 1 12 12 13 15 15 1 12 12 13 1 15
12 3 3 0 3 13 9 13 13 15 15 9 13
16 3 3 15 1 15 15 3 13 15 15 13 3 13 15 13 9
8 16 3 9 3 13 1 15 13
13 3 7 1 9 3 7 1 9 0 13 7 3 13
10 13 3 13 15 9 7 9 16 13 0
7 7 13 9 7 9 13 16
7 0 9 13 7 13 1 0
7 7 13 1 0 9 0 13
29 15 1 15 9 15 13 12 9 7 16 13 12 1 0 3 13 12 12 1 9 7 13 1 0 15 13 16 13 0
9 7 13 9 13 9 7 9 13 0
8 13 15 16 13 9 15 15 13
22 13 15 16 3 9 13 1 9 1 12 9 9 13 3 1 12 12 0 15 3 13 9
8 7 16 13 13 9 7 9 13
7 13 15 16 13 9 15 13
13 3 13 15 9 13 1 9 9 1 12 9 9 13
2 13 3
6 7 13 0 1 0 9
8 9 13 15 9 9 15 15 13
4 7 13 0 9
22 7 3 1 0 9 13 15 0 9 3 13 13 1 9 0 7 3 13 9 15 13 3
8 7 13 7 13 12 9 9 0
9 7 13 0 1 9 15 16 13 9
10 7 13 13 9 15 1 9 15 9 13
5 1 15 3 13 13
6 15 9 9 15 13 9
5 15 3 3 9 13
9 13 7 13 1 9 15 7 13 0
15 9 13 1 9 7 1 15 7 3 3 13 0 13 9 15
6 7 13 13 1 9 15
23 16 3 3 3 13 13 0 9 15 7 9 13 13 7 13 13 1 9 15 7 13 13 0
7 9 13 1 9 7 1 15
7 3 3 13 0 13 9 15
6 13 3 9 1 9 15
17 3 13 9 0 7 13 0 7 13 9 1 9 15 7 9 1 9
22 7 13 9 13 7 13 7 13 7 13 16 0 9 15 13 13 7 13 13 7 13 13
3 7 13 13
10 7 16 13 7 13 9 13 9 7 9
4 15 7 13 0
13 9 15 13 7 13 9 15 9 13 16 0 0 13
6 13 13 3 7 13 13
7 9 3 0 13 13 13 0
6 3 0 13 13 9 15
10 6 3 9 13 15 7 3 9 15 13
10 7 3 13 15 9 16 1 9 15 13
11 9 15 3 15 1 13 7 15 15 15 13
17 13 3 7 13 13 16 9 15 0 13 13 7 13 13 7 13 13
6 13 3 7 1 9 15
7 9 15 13 0 15 13 9
10 7 0 13 13 1 0 16 13 0 15
6 7 13 0 7 13 0
5 15 0 13 1 15
4 13 9 9 15
5 13 3 9 1 15
9 15 13 16 9 15 13 1 15 9
3 13 3 13
2 13 13
14 13 15 13 16 16 13 13 1 9 13 15 1 9 15
8 13 3 0 9 9 15 13 0
4 3 13 9 15
3 3 0 13
3 13 9 15
3 7 13 3
2 13 12
3 3 15 13
4 15 3 3 13
2 15 13
3 12 9 9
6 13 9 15 7 13 12
11 3 9 0 9 0 9 9 1 9 15 13
4 7 15 15 13
14 13 15 9 1 9 9 16 16 13 13 15 1 0 9
10 15 0 13 1 0 3 1 0 0 13
11 7 15 1 0 0 13 3 1 0 0 13
14 16 3 1 0 9 0 3 13 15 0 13 15 13 15
6 15 9 13 12 9 13
13 7 3 12 13 7 0 13 7 12 13 7 0 13
8 13 3 15 0 9 15 13 0
3 7 13 0
3 7 13 0
7 15 13 15 13 15 1 9
5 9 3 13 9 15
6 9 7 9 3 1 11
11 1 15 9 9 13 7 15 1 0 9 13
13 3 13 3 9 7 9 13 3 1 9 12 9 13
7 7 15 13 1 9 13 13
13 9 15 13 0 7 13 9 7 9 7 13 3 3
22 7 13 15 0 9 11 15 13 1 9 15 9 0 13 13 1 9 15 13 1 9 0
8 7 3 9 13 7 13 9 15
10 13 13 3 3 0 7 13 13 1 9
16 13 9 15 16 13 1 9 13 11 1 3 7 11 1 9 15
4 7 15 13 13
23 9 11 13 15 7 13 11 16 13 9 9 15 1 9 16 13 9 15 16 13 1 0 9
12 9 13 16 13 0 1 9 15 7 11 3 0
4 3 3 0 13
3 15 3 13
2 7 13
26 13 3 15 9 16 13 15 1 9 9 15 13 3 12 9 16 13 0 16 3 0 13 1 9 0 9
4 7 13 0 11
4 13 11 7 9
2 13 0
3 3 9 11
10 7 16 15 1 0 13 1 15 9 13
13 16 11 7 9 3 13 3 16 15 1 0 13 13
5 7 1 9 15 13
6 0 13 16 3 13 9
6 6 3 0 1 15 13
21 0 13 0 16 9 0 13 1 9 15 7 13 1 9 3 16 13 12 1 0 0
2 13 15
6 7 16 9 13 13 0
4 7 13 9 9
3 13 15 9
3 13 3 9
18 16 13 9 3 9 9 13 0 9 9 13 7 13 1 9 7 13 15
14 15 3 15 13 9 13 7 13 15 13 1 9 13 0
2 3 13
1 13
10 3 9 13 9 0 16 13 15 15 13
2 3 13
11 3 3 15 16 13 15 15 13 13 15 13
3 9 0 13
4 15 13 13 13
13 7 13 13 16 13 1 11 13 1 0 11 7 11
14 7 16 13 15 9 13 15 12 9 0 15 13 1 3
4 7 13 9 13
4 15 3 13 13
1 13
3 13 15 9
7 7 13 13 16 13 13 13
25 12 3 1 0 3 13 16 13 13 13 13 1 0 9 13 9 7 13 1 9 1 9 15 9 13
4 7 0 13 9
4 13 3 11 13
4 3 12 13 13
3 7 13 0
1 13
1 13
6 3 9 15 15 0 13
12 13 3 1 9 3 13 9 9 13 15 7 13
6 3 13 9 9 1 9
8 3 7 13 6 3 7 6 3
4 7 13 1 9
3 7 13 15
2 6 3
2 6 3
5 13 13 3 7 13
21 3 3 9 13 1 1 9 1 15 15 1 9 13 13 3 13 9 9 1 9 15
11 3 3 13 0 0 13 7 13 1 9 0
3 13 7 13
14 9 13 7 13 1 9 3 1 9 15 13 11 1 9
7 3 3 13 13 1 9 11
3 13 7 13
3 13 7 13
1 13
1 13
8 1 0 13 15 9 9 9 13
16 1 0 9 15 13 1 9 7 9 15 1 9 3 13 13 0
8 7 15 1 9 3 3 13 3
7 15 13 9 15 13 13 0
6 7 15 13 0 13 15
2 13 15
7 0 9 13 12 1 9 12
5 12 13 13 1 12
5 12 13 7 0 13
3 12 1 9
5 12 13 7 0 13
2 3 9
3 15 13 15
6 3 13 9 3 13 9
14 9 15 13 1 15 9 15 9 3 13 7 9 3 13
12 9 3 15 13 1 9 0 7 13 1 15 13
5 13 15 1 0 15
5 7 13 1 0 9
6 1 0 3 13 1 15
3 13 3 9
5 13 15 9 9 13
7 13 15 16 3 13 9 0
9 3 9 9 13 13 13 9 1 9
16 13 3 3 1 15 15 1 15 13 3 0 7 13 0 9 0
7 12 9 13 1 9 16 13
5 12 9 7 0 9
6 9 13 0 1 15 13
4 13 3 1 9
11 7 9 1 3 13 13 3 9 1 9 13
5 7 13 9 15 13
5 9 0 13 15 9
2 13 15
8 13 0 13 1 9 15 1 0
11 3 15 15 15 13 13 7 15 15 13 13
9 13 3 1 0 3 9 16 15 13
9 13 9 13 1 15 7 13 15 13
5 0 13 3 9 9
3 6 13 15
11 15 3 13 9 9 3 9 3 13 1 0
6 7 13 15 15 9 13
7 9 0 15 13 9 0 13
4 13 3 15 11
4 15 15 13 0
2 9 13
2 3 13
2 3 13
3 3 9 13
4 3 0 9 13
5 13 9 15 7 9
2 15 13
6 0 15 13 1 9 15
12 15 15 13 13 7 13 0 7 13 9 1 9
2 7 13
2 13 15
9 0 0 13 13 13 16 0 13 3
7 13 3 0 11 0 13 13
9 3 0 15 9 13 1 9 9 13
14 3 13 3 9 1 9 9 13 3 0 13 1 9 9
5 7 15 13 0 13
9 15 0 13 1 9 0 13 1 9
3 13 3 11
8 6 15 13 15 7 13 13 15
3 15 13 15
3 6 13 15
30 15 13 15 13 9 7 9 7 9 7 9 7 9 1 9 9 7 3 13 0 0 1 0 9 7 1 9 13 9 0
14 6 13 11 7 13 15 15 13 13 1 9 1 9 9
9 13 3 9 7 13 7 13 7 13
17 7 15 15 0 13 7 13 9 0 0 1 15 7 3 13 15 13
12 13 13 3 16 13 11 0 15 13 1 9 13
9 7 16 13 9 13 13 15 0 13
7 13 3 15 16 11 9 13
3 7 13 13
7 7 15 13 13 15 16 13
5 15 3 3 3 13
4 9 11 13 15
6 7 16 13 13 0 13
4 15 15 13 13
3 3 0 13
3 9 16 13
1 13
5 9 15 15 0 13
8 7 3 13 7 13 0 13 9
8 7 15 9 3 13 13 9 9
5 7 6 9 9 11
8 7 0 13 9 9 7 15 0
6 7 13 13 11 15 13
13 7 13 13 1 9 9 16 13 0 16 3 13 13
13 7 16 13 1 9 13 11 13 0 7 13 1 15
11 11 13 13 16 3 1 9 15 13 15 13
7 7 13 13 7 13 0 13
11 7 16 13 15 13 13 16 1 9 9 13
7 6 9 0 15 9 13 0
7 7 16 15 15 13 13 0
13 3 9 9 0 13 13 15 16 3 0 9 13 11
10 13 3 9 9 13 7 0 13 15 13
19 0 0 13 13 13 9 15 16 13 3 11 7 16 13 16 3 9 9 13
2 13 3
12 9 15 0 13 1 9 0 13 15 9 7 13
13 13 3 12 9 15 13 0 12 9 7 13 1 0
5 9 3 15 13 0
5 13 0 13 1 15
7 7 13 13 16 13 13 9
13 7 13 13 9 15 13 9 16 13 3 15 13 13
4 13 3 0 13
6 9 9 15 12 9 13
3 7 13 0
14 6 0 9 16 1 0 0 13 13 9 13 1 12 9
3 7 0 13
6 3 15 13 1 12 9
4 7 0 13 13
9 9 6 9 15 15 13 13 1 9
7 13 3 15 16 9 0 13
9 13 15 3 13 7 13 15 3 13
2 13 15
7 1 9 15 15 13 9 0
8 7 3 3 13 9 15 1 9
8 7 15 13 1 9 3 13 0
3 7 13 13
11 13 1 0 9 7 13 0 15 12 9 13
3 7 13 15
4 9 13 12 9
7 13 3 15 16 15 13 13
12 1 15 3 15 3 13 3 15 13 13 1 15
7 7 0 13 13 13 1 11
19 7 13 13 16 13 1 11 7 11 1 9 15 13 9 13 12 9 15 13
6 13 1 9 15 3 13
12 1 15 13 13 9 9 13 15 15 3 9 13
4 13 0 7 13
10 7 16 15 15 13 3 13 3 13 15
5 16 9 9 15 13
7 7 13 3 13 0 13 9
3 15 13 9
3 3 0 13
5 3 9 15 0 13
5 7 13 0 1 11
8 7 13 9 15 1 9 13 11
8 13 3 0 13 9 15 1 9
7 0 15 13 9 1 9 9
7 9 1 9 7 9 1 9
4 9 13 9 15
3 15 15 13
8 13 15 16 16 0 13 9 13
10 7 3 13 13 9 13 1 0 13 16
14 16 13 3 15 3 3 1 0 9 15 15 1 9 15
5 16 13 9 1 15
13 7 13 15 9 15 9 7 13 15 7 13 15 3
25 1 9 13 15 7 9 15 1 15 13 7 3 13 1 15 9 1 9 15 16 3 13 9 9 15
3 13 13 16
5 9 15 9 9 13
6 15 3 13 0 9 9
6 7 13 13 3 1 9
6 7 3 13 15 13 0
7 15 3 9 13 13 13 0
25 7 13 13 1 12 9 13 0 9 1 9 7 13 13 9 9 7 9 1 0 7 13 13 1 0
7 13 15 1 15 9 0 13
5 13 3 13 1 0
5 13 15 3 15 9
2 13 15
7 3 0 13 1 15 13 16
5 16 13 1 9 13
5 3 3 3 13 0
9 16 3 13 1 9 9 0 13 15
6 0 13 3 11 9 13
4 7 11 13 0
10 3 7 15 13 15 1 15 9 0 13
7 9 13 9 7 13 15 9
6 7 15 3 13 0 9
13 7 1 9 13 1 9 9 16 1 9 9 13 0
5 15 13 13 15 0
5 7 13 0 9 13
10 0 3 0 3 13 7 13 9 13 0
5 15 7 0 13 13
2 15 13
4 13 9 15 0
5 3 16 0 13 13
8 15 16 13 9 13 1 15 13
9 0 13 9 13 0 16 15 13 9
6 7 13 0 1 9 13
6 15 3 13 0 9 9
1 13
5 0 3 13 15 13
7 15 13 3 0 15 13 13
10 9 15 13 13 0 13 13 1 9 9
7 15 15 13 1 0 9 13
6 1 15 3 13 13 0
15 7 13 9 9 7 9 13 1 0 9 0 9 7 13 9
8 13 3 16 1 15 13 9 0
4 7 13 0 13
7 9 13 16 3 13 7 13
10 7 3 13 9 7 1 9 9 9 13
7 13 15 13 9 11 7 3
7 13 3 9 0 13 1 15
3 15 15 13
3 13 15 9
5 15 13 9 7 9
3 7 13 0
11 13 3 15 11 13 11 7 15 9 13 9
8 7 3 13 9 15 13 1 9
6 7 13 1 9 15 13
12 13 3 15 9 15 13 13 9 7 13 15 13
27 9 11 13 15 16 9 15 13 13 13 9 7 0 1 9 13 16 13 15 9 15 9 7 13 9 9 15
4 12 3 9 13
10 7 13 13 0 7 0 13 13 1 9
11 3 3 15 12 7 3 13 9 7 13 13
6 0 15 13 13 3 9
7 1 9 3 15 15 13 9
5 3 12 13 15 9
4 7 13 0 11
8 9 9 0 13 7 13 1 9
6 3 7 3 3 13 13
12 0 3 9 13 7 9 13 9 16 13 9 9
7 9 3 3 13 0 7 0
4 15 3 13 15
5 13 3 15 9 13
3 9 3 13
7 7 3 3 13 15 15 13
6 3 13 11 9 11 13
7 7 0 11 13 1 9 9
4 13 9 9 15
5 11 3 9 0 13
5 7 3 9 15 13
7 13 3 15 9 13 9 15
30 13 1 9 15 13 13 1 9 7 13 9 1 9 7 0 9 1 9 7 0 9 1 9 15 13 9 9 13 0 9
11 13 3 13 15 15 13 9 15 1 9 0
10 13 3 7 15 9 0 13 9 13 12
2 7 13
11 3 13 15 16 9 0 0 0 3 15 13
13 0 3 1 15 15 13 0 15 9 15 15 13 13
13 7 15 13 1 9 15 9 0 7 9 13 13 13
15 0 15 13 13 9 1 15 3 13 9 1 9 15 3 13
10 9 3 0 13 7 15 9 1 13 13
2 15 13
3 13 16 13
8 0 3 13 1 9 15 13 16
2 15 13
5 13 3 13 1 0
8 16 3 13 9 7 9 13 13
3 3 13 0
8 13 9 1 9 7 9 1 9
17 9 0 13 1 9 7 9 7 9 9 7 1 9 7 9 0 13
23 7 1 0 15 13 15 9 15 7 13 13 1 9 7 9 13 1 9 7 9 1 9 15
5 13 3 15 1 9
9 13 3 1 9 15 3 13 3 13
15 13 3 1 9 7 9 7 0 7 9 7 9 13 1 15
7 7 9 1 9 15 3 13
6 1 9 15 13 9 15
13 16 3 13 13 1 9 11 3 13 16 13 9 15
14 3 15 1 11 13 13 1 9 7 15 1 0 15 13
19 7 15 1 9 3 13 1 15 16 9 9 0 13 16 13 15 15 13 13
8 6 3 0 7 13 1 0 9
10 13 3 9 0 1 9 7 9 9 0
4 3 9 9 13
13 7 3 13 9 9 13 1 9 1 9 0 7 9
13 0 3 13 13 13 7 13 9 15 16 13 9 15
4 7 13 0 9
5 13 9 7 15 9
11 16 13 3 1 15 9 13 16 3 13 9
13 3 3 15 16 13 0 13 13 16 3 13 9 9
11 6 13 15 16 3 13 9 0 16 15 13
5 9 3 15 3 13
23 13 3 15 16 3 13 9 15 1 9 7 9 7 9 0 9 7 13 1 15 0 9 0
12 3 9 3 13 1 15 15 13 1 9 15 9
19 13 3 15 9 13 16 0 13 13 0 15 15 13 13 7 13 1 9 9
6 13 3 9 13 1 9
9 9 3 13 13 1 9 15 13 9
10 7 15 9 13 1 15 1 9 13 15
8 13 3 9 0 9 15 13 9
11 13 3 11 1 11 15 13 11 12 1 12
14 7 13 7 13 13 1 9 9 7 9 3 0 13 15
9 7 13 13 7 13 13 9 0 13
10 7 13 7 13 9 16 13 0 1 9
10 13 3 9 9 1 15 3 13 13 9
6 7 13 11 7 11 13
6 13 13 15 9 16 13
3 3 13 13
11 6 13 15 1 9 13 15 9 9 9 13
12 13 15 1 9 1 15 13 7 13 9 9 9
3 13 15 9
9 3 13 9 3 9 1 9 15 13
10 7 15 15 13 9 0 9 7 3 13
9 13 3 13 3 13 0 7 13 9
3 7 13 0
9 9 13 0 9 13 15 1 16 13
7 7 13 9 9 13 7 13
5 13 7 13 1 15
13 13 3 15 16 3 13 1 9 9 16 9 9 13
11 7 13 9 9 13 7 13 7 13 15 13
8 0 13 9 15 15 1 15 13
6 3 3 9 16 13 13
12 0 13 9 0 9 1 9 15 15 1 15 13
10 3 6 9 13 15 15 1 13 1 9
7 3 6 10 9 1 15 13
14 7 15 13 13 1 15 15 13 1 15 15 0 13 13
12 13 13 3 3 9 1 15 15 15 13 13 0
3 13 3 15
8 7 15 9 13 1 15 0 13
4 15 3 3 3
9 7 15 0 13 1 15 13 3 0
6 7 15 9 13 3 9
3 3 15 13
9 15 3 1 0 15 13 3 15 13
10 15 3 13 15 13 15 1 1 9 15
3 13 3 9
10 11 11 6 11 13 15 16 13 3 9
10 15 3 13 1 15 16 3 13 9 15
7 7 15 3 13 13 9 15
3 15 13 15
3 7 0 13
3 13 15 11
3 7 13 15
13 3 13 15 1 9 7 9 7 9 3 15 13 15
3 3 0 13
1 15
3 13 3 15
9 7 3 15 13 9 13 3 7 9
13 13 3 15 16 3 0 15 13 13 13 13 1 15
8 3 15 15 13 1 15 9 13
3 3 0 13
5 9 6 9 12 3
4 3 0 13 15
2 3 13
8 7 13 13 1 9 1 9 9
6 13 13 3 0 3 9
10 7 15 13 13 1 15 3 9 13 9
5 7 13 9 13 13
8 9 16 13 13 9 0 1 15
7 3 3 15 9 7 15 13
8 13 3 0 9 1 9 13 15
6 7 13 1 9 3 13
11 7 13 13 9 15 3 9 9 13 1 9
15 7 16 13 1 9 7 13 1 9 15 13 15 13 1 9
2 15 13
1 13
5 13 16 13 1 9
5 3 15 13 6 9
15 7 15 13 11 12 1 12 13 15 7 13 11 16 13 15
5 11 3 13 15 11
4 9 9 9 13
12 13 3 0 15 1 15 13 15 13 13 13 15
4 13 3 11 13
3 13 3 3
7 7 16 13 9 15 13 15
16 13 3 11 1 15 15 13 1 15 9 9 7 9 9 7 0
8 3 1 9 13 1 9 7 9
12 16 3 15 1 13 1 9 3 13 9 1 15
8 7 0 13 9 15 7 9 9
5 11 3 13 1 3
13 15 16 13 9 15 13 1 9 7 15 13 13 13
5 3 0 1 0 13
5 3 0 13 15 13
4 9 3 13 0
7 7 1 0 15 13 15 13
5 3 15 1 0 13
4 6 9 3 13
10 7 9 13 3 9 12 15 15 13 13
4 3 7 9 13
3 7 13 11
4 9 13 15 13
7 7 3 3 0 13 13 9
14 7 13 9 13 11 7 13 13 11 9 9 3 13 16
6 7 13 3 11 13 3
8 7 9 15 13 0 13 15 13
7 7 13 15 7 13 9 15
6 13 15 13 15 15 13
7 7 15 0 13 13 1 15
20 7 3 13 13 9 13 0 9 7 9 9 7 9 7 13 0 1 9 15 13
6 16 15 13 11 13 15
6 16 15 13 3 13 15
10 16 3 7 13 3 13 15 3 7 13
11 1 0 3 13 9 9 13 1 0 9 9
3 13 3 15
2 15 13
5 15 13 16 15 13
3 3 0 13
6 0 3 13 1 9 15
9 7 13 15 9 15 13 0 1 11
5 13 3 13 0 13
16 0 13 13 9 15 7 13 9 13 11 7 13 15 11 9 13
5 11 3 13 15 13
4 3 0 13 13
2 15 13
6 15 13 9 1 0 9
4 3 0 13 13
12 13 9 13 1 0 11 7 13 1 11 3 3
9 11 3 13 11 13 16 9 9 13
19 7 3 13 16 1 11 9 13 13 15 1 11 15 3 0 11 13 0 9
7 11 3 13 11 13 13 3
5 13 3 0 0 9
9 13 3 9 9 7 9 3 13 15
7 13 3 0 11 1 9 15
9 7 13 13 9 0 7 13 1 11
10 7 13 13 9 11 7 11 1 0 9
6 3 3 9 13 1 3
12 11 3 13 9 9 7 9 7 9 13 1 0
25 13 15 0 9 3 13 9 7 6 15 1 15 13 15 9 13 1 9 0 1 0 1 15 15 13
4 13 3 0 13
9 3 3 13 13 15 1 9 0 12
6 13 3 3 0 9 13
6 13 0 7 13 15 11
13 15 13 1 9 15 13 1 9 7 9 13 1 9
10 3 3 11 13 13 1 0 13 13 11
4 3 0 13 13
1 13
6 0 3 3 13 1 0
5 15 3 0 13 0
6 15 9 9 13 1 15
5 13 3 0 7 13
8 3 0 13 9 0 13 16 13
4 7 13 9 15
6 7 11 13 13 9 15
15 13 3 0 15 15 1 9 7 9 13 13 1 9 15 13
7 7 13 0 9 13 1 11
13 13 3 0 0 9 9 7 9 15 13 7 13 15
6 13 3 1 0 11 13
22 9 11 13 13 1 15 7 1 15 0 13 7 1 9 15 16 6 13 9 1 15 13
12 0 0 7 9 15 3 13 7 9 15 3 13
4 3 13 13 9
3 13 1 15
2 13 15
10 13 3 3 15 12 0 1 15 16 13
20 7 16 13 1 9 15 13 11 3 13 15 7 9 12 1 0 7 0 1 0
3 11 3 13
3 9 13 0
5 3 3 13 15 13
6 13 3 9 15 13 9
3 15 0 13
9 15 0 13 16 0 13 11 9 13
8 16 15 13 9 9 0 15 13
13 13 3 7 9 13 1 0 9 0 7 0 7 0
4 0 13 9 9
10 12 3 1 0 15 13 9 13 15 13
11 16 15 13 11 0 13 15 3 0 7 15
10 3 7 15 13 9 16 1 0 9 13
4 7 15 3 3
4 3 0 9 13
4 7 13 1 11
8 9 13 15 16 13 1 9 15
4 7 13 0 11
3 6 13 15
16 13 3 3 9 0 7 9 13 13 1 0 9 3 1 0 9
10 7 13 13 9 7 9 9 13 13 0
6 7 13 9 0 11 13
7 9 1 9 15 13 9 15
9 13 3 9 15 13 13 13 9 13
5 3 0 9 0 13
18 7 15 9 15 15 3 13 1 9 0 7 13 15 13 13 9 15 13
12 7 6 9 9 11 15 13 9 9 0 7 0
17 0 3 13 9 7 9 15 1 11 9 11 15 13 3 0 9 9
8 0 13 1 11 7 13 9 11
16 7 13 13 9 7 13 15 1 9 13 1 15 3 15 13 13
7 7 9 13 9 7 9 13
6 7 13 13 9 7 9
6 7 9 3 13 1 9
6 7 13 9 13 1 9
7 7 13 3 13 9 9 11
18 7 13 13 16 9 13 13 1 0 6 12 9 13 1 0 1 9 13
11 16 13 3 7 13 9 1 9 13 1 0
5 15 13 13 1 0
5 3 13 3 7 13
5 7 13 13 9 15
20 13 3 11 11 7 11 7 11 11 7 0 15 1 15 13 15 13 1 9 0
13 7 13 13 1 0 3 9 9 0 7 3 13 0
6 11 3 13 13 1 9
14 7 13 13 9 0 13 7 13 15 1 13 15 13 13
20 7 6 12 1 0 13 0 9 1 9 15 13 1 9 9 12 1 11 9 11
10 7 15 13 1 3 1 0 15 15 13
9 7 13 13 16 13 7 15 1 13
4 7 13 1 0
12 15 13 0 9 15 13 1 3 13 7 13 0
8 7 13 12 15 9 11 13 15
16 15 0 9 13 1 11 7 3 13 15 13 13 1 0 0 9
3 15 0 13
1 15
2 7 13
17 1 11 9 15 13 9 9 0 1 9 7 9 1 9 7 15 9
8 15 3 13 16 15 13 13 11
12 7 3 1 0 15 0 9 3 16 0 13 13
30 7 7 9 15 1 15 13 15 15 1 9 13 1 9 7 3 13 9 15 13 13 15 3 9 9 13 15 13 15 13
7 7 13 15 1 15 1 9
6 7 3 13 3 9 13
4 15 3 3 13
5 7 15 13 1 15
24 6 0 7 0 9 1 13 1 15 15 13 13 9 3 0 13 13 11 7 3 13 1 9 15
6 7 15 15 13 3 13
4 7 13 0 13
10 13 15 1 16 13 7 13 13 3 9
4 7 13 1 0
16 7 13 13 16 13 1 0 13 9 7 13 7 13 7 13 0
8 7 13 13 9 15 7 13 15
6 7 15 13 1 9 15
15 3 9 15 13 13 1 15 16 13 1 9 7 13 15 9
12 7 13 13 12 7 15 15 1 15 13 13 16
6 13 9 3 7 13 11
15 7 15 13 15 13 13 1 9 7 3 13 15 1 9 9
12 16 0 3 13 11 13 1 0 15 7 13 15
2 9 15
2 15 13
8 13 3 7 13 13 15 9 13
3 7 13 15
9 13 9 15 7 9 16 0 15 13
14 13 7 13 16 9 9 7 9 3 13 3 15 13 13
9 7 16 0 13 13 15 9 7 9
10 3 3 0 3 13 7 13 1 9 13
5 13 3 15 15 13
9 7 16 13 1 15 13 9 13 15
4 7 13 1 15
30 0 13 9 15 13 13 1 15 16 3 13 15 1 16 3 13 13 15 15 13 13 1 9 11 7 9 7 9 1 15
5 15 3 13 9 0
8 7 15 13 9 9 15 1 15
10 15 3 13 1 9 16 13 9 1 0
12 13 3 15 3 1 11 7 13 9 15 13 15
10 7 15 13 13 13 1 11 1 9 0
9 7 13 3 1 9 13 7 13 9
1 6
13 1 9 13 9 7 9 13 1 9 7 9 13 9
5 15 1 15 13 13
9 7 1 15 13 13 15 15 13 13
9 1 15 9 13 7 9 13 9 9
9 13 9 13 1 9 15 9 13 11
14 0 13 1 9 16 9 13 1 9 16 15 13 1 0
10 3 13 0 9 7 16 9 13 1 9
10 13 9 0 15 13 15 9 13 1 9
14 1 9 13 7 9 1 15 13 13 7 9 15 3 13
16 3 3 13 15 13 15 9 9 9 13 0 15 13 1 9 15
19 15 3 1 9 3 7 1 9 9 3 7 1 9 9 7 1 9 13 13
13 7 13 9 15 9 3 0 1 9 0 9 7 9
8 11 9 13 1 15 7 13 13
5 0 13 15 13 15
13 15 1 15 13 13 1 15 13 13 16 0 15 13
11 7 1 9 15 15 15 13 7 9 1 9
6 3 9 1 11 13 13
4 9 15 13 3
18 7 0 13 9 11 3 13 9 1 11 9 7 9 1 15 16 13 15
3 15 15 13
10 7 13 13 7 3 13 7 13 13 16
4 3 13 15 11
3 7 13 15
2 15 3
3 11 13 15
3 9 13 15
2 7 13
1 3
3 13 3 15
2 15 13
7 16 9 13 0 15 13 15
5 15 13 1 15 0
1 13
7 13 9 9 3 13 11 9
7 7 15 13 13 13 1 9
6 7 13 15 7 13 15
14 15 3 13 16 15 3 13 11 3 7 11 3 7 9
4 13 15 11 13
4 15 13 1 9
8 0 3 15 13 15 15 3 13
22 15 13 15 1 15 13 13 15 1 15 13 13 15 15 3 13 0 16 13 15 9 9
7 6 9 9 15 13 9 9
5 0 13 1 15 13
13 1 15 13 9 15 1 15 13 13 16 0 15 13
14 7 15 13 15 7 16 13 11 3 13 15 1 9 13
6 7 9 13 11 13 16
11 13 9 13 3 9 1 9 7 13 1 15
4 7 15 13 15
16 1 15 13 9 13 7 13 1 15 0 13 15 13 1 9 0
8 7 9 13 16 0 13 9 9
10 0 9 3 13 11 7 1 9 15 12
5 7 13 11 13 13
3 6 9 9
10 7 13 15 12 9 13 7 13 13 11
9 13 3 11 7 13 15 13 13 15
3 15 13 15
7 9 15 13 13 9 3 13
3 13 7 13
11 13 7 13 3 13 7 1 15 13 9 0
5 9 3 13 3 0
17 13 3 11 9 11 11 12 1 12 15 13 1 11 7 13 13 15
9 13 0 3 9 15 11 7 13 15
5 7 13 15 1 11
5 13 3 15 11 13
5 15 13 11 9 11
9 1 0 13 13 1 11 7 13 11
4 7 13 15 11
2 13 15
9 13 3 11 1 11 9 11 7 11
13 15 13 11 1 9 7 9 13 11 9 11 1 11
4 7 13 15 11
6 1 11 13 15 0 13
3 13 15 11
10 13 11 11 13 1 15 7 13 1 15
8 6 3 9 1 15 9 3 13
3 13 15 11
5 13 11 7 13 15
10 16 15 11 13 16 13 1 9 13 15
5 13 15 11 7 13
5 9 15 13 9 9
4 15 13 9 11
8 16 13 15 13 15 1 9 13
3 0 0 13
4 6 6 13 15
12 13 9 13 7 9 9 13 7 13 1 9 9
14 7 9 0 9 13 13 1 11 11 7 13 9 11 3
11 13 13 3 3 7 11 7 9 15 1 9
8 7 13 9 13 9 11 1 15
3 9 3 13
6 15 15 7 15 13 9
4 13 9 15 9
4 15 13 15 13
16 13 3 3 0 9 12 13 1 9 9 13 0 9 0 7 0
3 13 15 11
3 13 9 9
6 7 13 15 3 1 0
4 7 13 15 11
24 16 3 13 9 9 9 13 7 3 13 3 13 9 3 13 15 13 9 13 9 9 7 13 15
15 15 9 3 0 9 13 7 1 13 13 3 15 15 0 13
6 15 13 0 9 3 3
18 0 13 9 9 11 1 11 11 7 13 9 15 7 13 1 15 9 15
14 1 0 13 11 15 7 9 15 7 9 15 7 9 15
6 7 3 13 3 0 9
9 7 3 13 9 9 7 13 11 11
13 7 13 1 9 13 9 7 9 7 9 7 0 13
6 7 0 15 9 13 13
3 13 0 3
7 13 13 9 9 15 9 9
8 13 3 13 9 15 16 13 13
5 9 9 15 13 15
6 13 3 9 7 13 15
7 15 9 13 15 16 0 13
5 13 11 7 13 15
14 12 7 12 9 13 13 9 0 7 15 12 9 13 0
7 0 3 13 1 9 9 15
20 16 3 13 1 0 13 13 9 15 16 0 13 7 13 9 7 9 15 13 11
19 16 3 13 11 1 9 1 9 9 0 13 1 9 15 13 9 15 15 13
26 0 3 11 3 13 15 3 0 15 3 16 15 13 15 7 16 9 15 3 13 16 15 9 13 1 9
7 15 3 13 15 13 1 9
9 13 3 9 1 9 11 9 9 9
7 9 13 16 1 9 13 9
5 13 11 7 13 15
4 6 6 13 15
10 16 15 13 13 3 3 13 13 9 9
4 13 1 15 11
7 3 13 9 13 16 9 13
10 3 13 1 9 9 15 3 13 7 13
4 6 6 13 15
14 16 15 13 13 1 9 7 9 3 13 13 1 9 9
8 7 15 13 13 1 9 9 13
5 3 13 16 13 15
4 13 15 13 3
16 9 3 13 13 7 9 15 13 7 3 13 3 13 7 3 13
8 3 13 15 15 13 13 1 9
4 3 13 0 13
5 13 11 7 13 15
7 15 13 9 11 7 0 13
13 16 0 13 15 7 3 13 3 16 13 15 0 13
16 7 15 13 1 9 3 15 13 1 9 9 9 15 13 1 9
24 7 3 11 13 9 1 9 3 13 13 9 9 16 15 15 13 1 0 3 13 7 13 9 0
22 3 3 13 9 9 16 9 15 0 13 16 15 15 13 1 15 3 13 7 13 9 0
6 15 13 1 15 3 13
15 15 3 3 13 3 13 13 16 3 13 1 9 0 9 9
16 0 13 3 9 16 9 13 1 9 7 13 9 3 9 3 9
5 13 3 15 0 9
16 15 3 13 9 13 1 9 16 13 15 9 16 1 9 13 13
10 1 0 13 11 7 9 15 1 11 9
7 7 3 13 1 15 7 13
7 3 3 13 13 1 9 11
11 13 13 3 9 1 9 11 1 9 1 9
7 7 13 1 11 7 13 15
19 9 15 13 15 1 1 11 15 15 9 13 6 0 13 7 15 13 1 15
4 13 11 7 13
8 0 15 15 9 13 16 13 15
9 3 13 11 7 16 13 13 1 0
13 9 3 9 15 13 7 13 15 9 13 1 9 9
6 0 3 9 15 13 13
6 0 13 13 15 3 13
6 15 3 13 1 15 13
11 15 13 1 9 1 9 13 7 1 9 13
7 15 1 9 13 1 15 13
5 7 9 15 15 13
7 15 3 13 9 9 9 13
7 3 3 1 9 13 9 9
9 9 13 9 7 15 13 1 9 15
7 15 13 1 9 13 9 0
14 15 3 0 13 9 3 13 9 7 9 9 13 1 15
30 3 3 13 11 16 13 9 16 11 0 9 13 7 13 3 11 16 11 3 13 7 9 15 13 11 7 13 3 1 11
6 13 3 15 13 1 11
9 11 3 13 1 9 13 3 1 9
4 9 13 3 0
6 13 9 1 11 13 9
3 13 15 11
3 13 15 13
9 9 3 15 13 1 9 16 9 13
6 13 3 15 9 0 0
13 3 15 9 16 13 13 1 15 13 15 13 9 0
5 13 11 7 13 15
23 16 13 9 9 7 15 13 15 13 15 13 15 13 15 3 13 1 15 7 13 15 9 0
3 13 15 9
10 9 3 1 15 13 13 7 9 0 13
5 3 3 13 9 0
22 3 15 0 13 9 15 11 15 13 15 9 7 15 1 15 13 7 9 15 7 9 15
5 13 11 7 13 15
8 15 15 13 1 9 0 13 3
4 13 1 15 9
13 9 13 15 0 9 16 3 13 3 7 13 3 13
3 13 15 11
7 13 13 9 15 7 13 3
4 13 9 7 13
3 3 13 9
3 13 15 11
3 3 13 9
3 0 3 13
3 13 15 9
6 9 13 16 9 13 15
16 9 15 1 9 0 13 7 15 13 16 11 13 9 3 13 13
3 13 15 11
18 9 13 15 16 13 9 3 3 7 1 9 0 3 7 1 11 13 9
9 15 13 15 13 16 9 1 9 13
15 7 13 9 7 3 13 3 0 9 13 9 1 9 7 9
3 9 13 9
11 7 15 15 13 15 1 9 7 9 13 13
3 13 15 9
7 13 16 11 13 15 13 11
7 16 3 13 0 15 13 15
6 15 13 15 13 15 1
11 7 3 13 9 15 7 13 16 1 9 13
6 15 3 13 15 13 7
13 13 3 9 15 9 7 13 1 9 7 13 0 9
1 13
8 13 9 15 13 15 15 15 13
4 3 15 13 11
5 3 13 15 9 13
2 9 13
4 0 3 13 15
7 15 9 13 13 15 15 13
5 3 15 13 15 13
3 13 15 11
14 15 9 13 16 13 9 15 15 13 15 16 13 9 15
3 6 13 15
12 13 9 15 7 13 9 16 0 13 3 1 9
20 7 15 13 9 13 7 13 9 1 9 0 16 3 15 13 3 13 7 15 13
16 1 0 3 13 9 0 16 15 13 15 13 7 15 13 15 13
8 15 13 15 13 15 15 3 13
15 1 9 3 0 0 13 1 15 9 1 9 9 9 13 16
5 13 15 15 15 13
5 7 13 3 12 9
7 7 3 0 13 1 9 15
4 7 9 13 16
6 3 3 1 15 9 13
11 0 3 13 7 13 16 0 13 3 9 9
10 1 12 3 9 13 3 7 13 1 11
17 16 3 13 1 11 13 15 9 16 15 13 15 13 11 1 9 0
10 13 3 3 1 11 11 3 13 9 9
8 7 13 15 9 15 9 13 11
22 0 16 13 16 11 13 1 11 1 11 13 1 15 7 13 15 16 13 7 13 9 15
3 13 3 13
5 13 3 11 1 15
7 16 9 7 9 13 3 13
4 13 1 15 9
1 13
3 9 15 13
9 13 9 9 15 13 15 11 7 13
14 3 3 15 13 9 13 15 7 13 13 16 9 15 13
9 13 3 9 1 15 1 15 3 13
10 7 13 15 16 3 9 0 13 15 9
12 13 3 9 16 0 9 13 1 15 13 15 11
3 9 15 13
12 0 3 0 9 13 11 16 13 1 11 1 11
10 1 0 13 9 0 9 7 13 11 11
13 13 3 11 1 0 9 15 13 3 11 12 9 13
12 1 0 13 9 0 13 0 0 0 13 9 9
13 13 3 15 9 3 12 7 12 9 13 1 9 15
14 0 1 13 11 13 7 13 16 0 3 9 13 13 15
3 13 0 13
3 13 15 0
3 13 15 11
6 13 13 9 15 7 13
6 7 3 0 13 13 9
6 7 13 9 15 7 13
6 13 3 9 1 0 9
6 13 9 0 15 13 13
2 9 13
2 13 15
5 13 9 15 7 13
3 13 3 15
7 15 13 0 9 15 13 15
5 13 9 15 7 13
9 15 3 15 0 13 13 13 15 13
7 11 3 13 9 13 1 9
4 6 0 13 13
8 3 13 13 16 3 15 15 13
9 3 13 9 11 16 0 13 1 9
4 11 3 13 15
8 9 15 3 3 13 7 15 13
22 3 3 3 13 15 9 13 16 3 3 13 9 7 3 9 15 13 9 0 15 13 9
6 13 3 11 7 13 15
12 3 13 9 1 15 13 15 3 15 13 9 13
9 15 3 0 13 0 3 9 3 13
11 9 3 13 9 7 15 13 15 15 15 13
13 3 3 9 13 0 7 13 3 3 9 15 13 13
6 3 7 3 9 13 15
12 7 9 15 13 9 16 15 13 9 3 13 9
10 15 3 13 9 3 13 9 15 13 0
16 6 6 13 15 16 13 9 7 3 13 3 0 13 9 9 9
4 7 15 13 13
19 3 3 9 13 9 1 15 3 0 3 13 3 9 9 13 1 15 3 0
11 7 9 13 15 7 9 13 16 9 9 13
15 7 13 15 0 13 1 9 9 15 3 0 13 1 9 9
8 3 13 15 1 15 0 13 15
19 3 13 13 7 9 15 0 13 16 3 13 9 15 7 9 15 15 13 15
7 15 13 15 9 13 1 15
10 7 13 16 0 13 9 15 13 1 15
8 15 13 1 11 7 9 13 9
7 15 3 3 1 9 9 13
7 7 0 13 16 15 0 13
9 15 3 13 13 1 9 1 9 15
6 15 3 13 9 0 11
10 7 15 13 15 9 15 9 13 1 15
11 3 7 9 15 3 13 3 7 9 15 13
16 7 9 15 3 13 1 15 13 16 15 13 0 0 15 3 13
10 13 9 16 15 13 1 15 9 0 13
8 7 0 13 15 9 13 1 15
9 7 3 13 13 1 15 16 9 13
10 7 13 15 16 9 9 3 13 1 15
8 16 15 13 1 9 15 0 13
18 3 13 15 13 15 9 1 3 13 7 9 15 1 0 13 9 3 13
9 13 13 16 15 13 13 15 1 9
9 13 15 13 15 11 1 15 15 13
8 16 3 13 11 13 3 3 15
5 1 15 3 0 13
10 16 3 0 9 3 13 3 15 9 13
11 13 3 1 9 11 7 3 13 1 9 15
7 13 3 9 9 9 0 9
16 16 13 3 9 11 7 13 16 9 0 13 1 15 13 1 11
6 3 13 9 16 13 0
5 0 3 13 13 15
6 15 3 13 15 13 13
3 13 15 11
11 12 9 9 3 13 15 16 15 0 15 13
12 13 9 12 0 15 13 12 9 0 7 12 9
6 7 0 15 13 1 0
3 13 3 11
3 13 9 13
6 13 3 9 0 1 9
7 13 3 9 9 3 12 12
4 13 3 9 11
12 7 16 9 13 13 13 3 7 1 9 3 13
16 13 3 7 13 12 9 9 1 12 9 0 15 13 0 15 13
10 0 3 9 16 13 15 13 9 13 16
9 0 13 3 9 15 13 13 1 9
20 11 3 16 13 16 13 13 16 13 15 7 13 15 9 13 3 1 9 0 0
10 3 3 3 13 13 13 9 15 1 9
9 7 1 13 9 13 1 9 1 11
11 7 9 3 13 13 7 3 13 1 15 11
19 16 13 3 3 9 12 7 12 13 11 13 1 9 7 0 9 13 7 13
2 15 13
2 13 13
14 13 3 13 15 1 9 7 3 13 9 1 9 15 13
31 0 9 9 15 13 1 9 13 16 9 15 3 13 3 3 12 7 16 3 13 1 9 15 11 1 9 7 0 9 15 13
14 15 3 13 9 1 11 1 9 3 13 9 9 13 9
20 16 3 13 9 16 11 3 13 3 3 7 9 15 13 9 7 13 11 13 11
4 9 3 3 13
5 13 15 11 7 13
14 13 15 3 16 13 9 7 16 13 1 9 7 13 13
16 13 3 9 15 13 7 15 13 1 9 0 15 9 9 15 13
5 0 3 9 13 9
4 13 3 1 15
6 15 13 16 13 9 9
11 0 13 9 9 16 13 1 15 15 13 0
3 13 3 15
10 15 3 15 13 9 16 13 7 13 15
9 9 15 9 13 1 9 3 13 13
6 9 1 9 13 15 13
4 13 3 15 11
4 6 6 13 15
12 9 3 9 13 15 13 1 9 7 13 9 9
4 13 3 1 15
6 9 3 13 15 9 0
4 13 3 15 11
14 15 13 1 15 3 13 7 15 13 1 15 3 13 3
10 7 13 15 16 7 13 15 7 3 13
8 15 15 13 15 9 1 15 13
15 3 13 1 9 3 16 13 9 15 7 9 15 15 13 15
23 0 13 3 9 15 15 13 15 9 16 15 15 13 15 3 13 1 15 7 13 0 0 9
28 0 13 3 9 9 15 15 13 15 16 15 15 13 9 7 13 1 15 13 9 0 7 13 15 15 1 0 9
7 13 3 9 1 0 16 13
7 15 13 9 15 1 9 13
12 3 0 13 11 9 11 15 15 13 9 7 9
5 3 3 13 0 16
6 13 3 11 7 13 15
4 13 13 1 3
18 15 13 13 1 15 16 9 15 13 15 13 15 7 15 13 15 0 9
4 13 13 1 9
5 7 13 15 0 9
10 15 15 13 1 9 7 13 13 1 15
3 0 13 9
7 15 13 1 15 13 9 0
4 15 13 9 9
9 9 15 13 1 9 9 7 13 13
14 0 13 9 1 9 13 16 16 15 1 15 13 3 13
8 15 13 9 0 15 1 9 13
9 16 15 13 1 0 9 13 1 0
11 7 9 15 15 13 9 15 13 1 9 9
4 13 3 15 11
4 6 6 13 15
14 16 13 9 9 9 7 13 15 9 3 13 9 1 15
11 15 13 15 9 7 13 15 9 13 9 0
7 7 15 13 15 1 0 9
6 9 3 15 3 13 9
6 7 9 15 3 13 9
15 15 13 15 9 7 13 15 9 1 15 13 7 15 1 0
16 0 13 9 15 1 9 13 3 3 13 9 15 9 7 0 13
7 15 13 0 9 13 1 0
7 0 13 1 9 13 1 11
7 0 3 13 1 9 15 13
4 0 13 0 9
4 15 13 15 13
15 13 3 11 1 15 3 0 16 13 1 0 9 15 13 15
3 0 15 13
4 9 3 13 15
10 9 15 15 13 13 15 9 7 9 13
8 7 13 15 1 15 15 3 13
13 13 3 1 9 11 15 13 13 7 15 13 13 15
2 7 13
16 3 13 15 16 15 13 13 1 15 16 13 15 13 1 9 15
7 1 0 0 9 15 13 3
5 13 3 11 1 12
5 13 3 15 11 11
4 9 1 15 13
4 9 9 0 13
11 7 15 13 7 13 16 15 13 11 9 9
3 13 15 11
5 3 15 15 12 13
5 13 3 11 11 11
10 0 3 13 13 15 16 13 12 1 12
11 3 3 13 1 11 13 16 13 15 9 13
8 13 3 1 0 9 0 9 9
6 13 3 1 15 9 15
15 13 3 7 13 1 11 16 3 9 15 13 9 15 15 13
12 15 3 1 0 15 13 7 13 0 1 3 13
7 3 3 9 15 13 1 15
4 13 3 15 11
4 9 15 3 13
5 3 13 9 13 15
14 15 3 13 16 15 9 13 1 0 16 9 15 0 13
6 15 13 1 9 0 0
13 15 3 13 1 9 0 0 16 15 9 3 13 13
18 3 3 13 9 15 3 3 15 13 1 9 0 3 3 7 3 1 0
9 9 3 13 15 1 9 0 7 13
3 3 13 0
8 7 9 0 1 15 13 1 9
2 0 13
3 15 3 13
4 3 7 13 9
11 3 3 9 0 13 13 11 1 9 7 13
4 7 13 9 13
7 3 0 9 13 16 3 13
5 13 15 11 7 13
10 15 9 3 13 15 7 15 15 13 15
9 15 1 15 3 0 13 9 0 13
17 15 3 13 9 15 15 13 0 0 0 13 7 9 1 0 3 13
6 7 15 1 15 13 9
4 15 15 13 13
4 13 9 7 13
2 9 13
4 15 15 13 13
5 13 11 7 13 15
18 3 11 13 15 9 3 16 1 11 13 7 1 9 7 1 9 13 9
8 13 13 1 9 7 0 9 13
5 13 3 15 1 11
6 3 0 13 15 13 13
8 7 6 3 13 7 15 15 13
8 3 3 13 9 16 0 13 11
5 7 0 13 3 13
8 11 3 16 13 15 13 3 13
16 7 1 15 0 3 13 7 13 0 15 13 15 15 15 3 13
11 15 13 15 16 1 15 13 7 15 15 13
4 13 3 15 13
11 7 15 13 1 0 9 16 3 13 9 15
9 1 9 3 0 13 1 15 7 13
11 11 16 13 3 0 9 13 3 15 0 13
7 13 9 9 13 1 0 0
9 7 13 9 7 9 9 16 13 15
6 3 0 9 15 1 13
7 7 13 1 15 15 13 15
5 13 15 7 3 13
8 7 3 13 15 15 3 13 13
6 13 3 9 1 15 0
8 3 0 13 13 16 3 13 15
9 3 1 9 9 13 13 7 13 9
6 15 13 0 9 15 13
11 1 0 3 9 0 9 13 11 7 13 13
8 16 15 13 13 1 15 7 13
14 15 13 1 15 3 13 9 9 1 9 15 13 9 0
11 0 3 13 1 9 15 13 13 13 1 15
9 3 3 13 9 16 11 3 13 13
10 1 0 3 9 16 13 0 9 15 13
4 0 13 3 9
3 0 13 11
5 3 1 11 11 13
4 3 9 13 16
11 1 9 11 7 11 9 3 13 11 13 11
8 9 3 13 13 1 9 1 15
7 15 3 1 15 13 13 15
6 7 15 13 1 0 9
4 7 13 15 0
4 3 3 13 15
8 3 3 13 13 9 3 0 9
4 13 3 15 9
5 3 3 15 13 13
10 3 15 1 9 13 1 15 7 1 9
9 7 9 0 15 3 13 9 13 13
14 3 9 15 13 9 16 13 1 15 3 7 13 15 13
4 13 7 13 15
5 3 3 15 9 13
7 7 13 13 15 1 9 15
6 11 3 13 1 9 9
16 7 9 3 13 1 9 7 15 9 13 1 15 7 13 13 15
9 13 3 9 7 9 9 1 9 13
8 9 0 9 3 13 13 1 9
9 1 9 3 11 13 15 0 9 13
4 15 3 15 13
9 0 3 13 13 15 16 13 13 15
10 16 3 13 13 15 13 15 7 13 15
10 15 1 9 13 15 0 1 0 9 13
7 7 3 15 13 13 1 9
8 7 13 0 7 9 1 0 13
6 13 3 15 11 13 15
3 9 3 13
3 15 15 13
2 15 13
3 13 3 11
4 3 15 15 13
7 3 3 13 13 15 11 13
4 15 13 9 9
11 15 13 15 3 13 1 9 7 13 9 9
4 13 3 15 9
6 15 1 15 0 9 13
5 9 15 3 13 0
12 7 16 15 9 13 1 15 0 0 13 9 15
8 15 3 13 3 13 7 3 13
4 15 1 9 13
4 15 3 13 15
19 7 16 13 15 9 15 0 13 16 0 3 13 7 15 7 15 15 13 9
12 7 1 9 15 13 13 16 12 9 9 0 13
17 15 13 15 9 13 1 15 0 7 9 13 1 15 15 13 15 9
3 13 3 15
8 3 7 15 13 3 7 9 15
8 16 15 13 3 3 9 15 13
9 0 9 13 13 1 9 13 1 9
9 7 15 13 15 16 3 13 9 15
5 13 3 3 15 11
10 15 13 7 13 15 7 1 9 15 13
7 3 15 13 15 3 13 13
3 13 3 9
7 3 15 13 15 3 13 13
3 7 13 15
4 15 1 3 13
4 15 1 0 13
5 15 1 9 0 13
6 15 3 13 1 0 9
8 13 3 15 16 13 1 9 15
11 16 3 3 13 16 15 13 13 1 9 15
3 13 15 11
5 9 16 7 13 15
23 0 13 1 15 13 7 13 7 15 13 15 0 13 7 15 15 13 1 15 0 13 1 9
7 7 3 13 16 9 15 13
4 13 3 15 11
22 16 13 9 9 3 13 16 15 13 7 1 15 0 13 15 7 3 13 15 9 0 13
7 7 15 15 13 15 1 13
8 3 15 15 13 13 15 13 3
9 13 3 11 1 0 15 13 15 9
17 16 15 13 1 9 15 3 9 15 13 7 13 9 7 9 13 15
2 13 15
7 9 11 13 7 15 13 3
3 3 15 13
2 0 13
5 6 6 13 15 16
7 15 15 13 9 9 13 9
4 9 13 1 0
8 16 3 9 15 13 3 0 13
5 13 16 9 11 13
11 7 13 15 13 16 9 15 3 13 1 15
6 15 15 13 1 9 13
4 13 7 13 15
4 9 15 11 13
3 13 15 11
15 3 3 13 15 13 9 15 9 15 13 13 15 13 1 9
4 0 11 3 13
5 15 13 9 9 15
3 13 3 15
4 12 9 13 9
4 13 3 15 11
8 16 9 9 15 13 13 3 15
7 15 3 1 9 13 7 13
5 3 9 15 3 13
6 16 3 13 13 9 15
5 15 1 9 9 13
16 0 9 13 1 9 7 1 9 3 13 16 3 13 9 1 15
12 16 13 9 1 0 13 16 9 13 7 9 15
8 15 3 16 9 13 3 13 15
7 15 1 15 13 15 1 9
8 16 9 13 3 15 3 13 15
9 3 15 3 13 16 1 9 3 13
6 13 3 9 7 13 15
2 13 11
4 15 9 3 13
8 7 13 9 15 7 15 13 15
6 15 3 3 13 9 15
5 13 15 13 7 13
4 6 6 13 15
3 13 3 9
8 11 13 13 7 9 7 15 13
10 16 15 9 15 13 3 13 9 1 0
10 3 15 0 13 9 15 11 15 13 13
4 3 9 13 13
4 15 15 0 13
2 13 11
9 16 15 13 15 0 9 15 15 13
4 15 3 13 15
11 7 16 13 16 3 13 15 13 0 15 9
7 7 13 15 7 9 15 13
8 11 9 15 13 16 13 9 15
5 7 13 7 13 13
5 13 3 9 1 15
7 12 9 3 13 7 11 13
3 13 15 11
5 16 11 13 15 13
7 13 3 9 16 13 1 15
8 11 3 13 15 7 13 1 9
7 7 13 13 9 0 1 9
5 7 13 15 9 15
10 9 15 13 0 7 9 15 16 0 13
2 13 11
15 3 7 0 13 3 7 9 15 7 16 13 9 9 1 0
7 3 1 9 13 9 13 9
20 0 16 13 13 1 9 7 13 9 1 9 7 13 9 1 9 15 7 13 15
1 13
7 13 1 9 11 15 13 13
7 13 3 7 13 7 13 13
11 3 9 7 15 13 15 3 16 0 13 13
7 3 0 13 15 13 7 13
2 0 13
5 3 7 0 13 15
3 0 13 16
2 15 13
3 13 3 15
5 3 13 13 9 15
1 13
7 7 13 9 15 7 13 15
6 13 1 9 11 7 13
2 13 15
3 3 13 0
1 13
1 13
7 13 15 1 9 15 0 13
7 3 3 13 15 9 3 13
4 0 3 13 15
9 9 13 15 1 9 7 13 7 13
10 3 13 0 9 1 9 16 9 3 13
2 15 13
7 3 13 9 9 0 9 13
5 7 9 13 1 15
9 15 15 13 1 15 15 13 9 15
4 0 3 13 16
2 9 13
17 3 13 3 9 1 0 16 0 13 7 13 16 13 9 15 15 13
11 0 13 9 15 15 15 13 16 0 13 13
4 3 3 3 13
6 13 15 9 15 7 13
5 3 3 3 13 13
7 7 15 15 13 9 15 13
2 15 13
2 9 13
4 15 1 15 13
13 3 3 13 9 16 16 15 15 13 11 1 9 13
5 3 9 15 13 16
2 15 13
10 13 3 3 9 15 13 0 7 13 15
3 13 9 9
7 15 13 16 0 9 9 13
3 13 3 0
4 16 9 13 13
3 13 3 0
4 3 13 15 9
2 13 15
5 13 15 3 7 13
4 15 3 13 13
7 3 3 15 13 9 15 13
4 13 15 7 13
4 15 9 0 13
5 0 3 13 3 13
6 13 0 9 7 13 15
14 1 0 3 0 13 16 15 13 3 13 7 13 15 9
7 13 3 16 9 9 3 13
12 7 16 15 9 9 13 7 9 15 13 0 13
11 1 9 3 13 13 16 13 15 9 0 13
9 16 13 0 1 9 3 13 13 15
4 13 7 13 15
4 7 13 15 3
6 13 11 16 13 15 3
6 7 16 13 15 13 15
5 15 13 1 9 9
4 13 0 7 13
7 15 13 9 16 13 1 15
4 7 13 15 11
10 7 13 15 7 15 13 15 1 15 13
4 7 13 13 15
3 13 15 11
17 1 9 15 1 0 9 13 16 15 3 13 13 7 15 13 0 13
11 7 13 1 9 15 1 15 13 7 13 15
5 3 3 15 0 13
3 13 15 11
6 16 0 13 3 13 9
1 13
4 6 6 13 15
16 15 3 13 1 9 1 9 9 7 13 3 0 9 13 7 9
8 15 3 13 1 9 9 13 9
16 0 9 13 7 9 9 15 13 7 0 9 13 3 7 13 15
8 7 16 0 9 13 1 15 13
8 7 9 0 13 16 13 9 15
5 0 9 13 15 11
7 0 3 3 13 15 13 15
5 6 6 13 15 16
4 15 13 9 9
12 15 3 13 9 13 7 9 7 3 13 15 9
3 15 13 9
6 1 15 16 15 13 13
10 9 3 13 3 16 13 7 13 7 13
8 15 13 16 9 13 7 3 13
4 15 13 9 0
19 9 7 15 3 13 9 15 3 13 9 0 13 9 13 7 13 9 7 13
6 7 9 13 7 13 9
13 9 3 13 16 9 13 7 3 13 1 15 1 9
4 15 13 9 0
8 3 13 15 9 3 15 13 9
6 7 9 15 13 1 9
10 7 15 9 13 15 3 13 1 0 9
15 7 0 13 15 13 7 9 15 13 7 13 12 9 12 9
5 15 13 15 1 15
4 7 15 13 15
13 1 15 0 9 13 13 15 7 9 13 3 13 15
9 9 3 13 13 1 9 1 9 0
5 13 3 0 1 15
4 9 13 7 13
3 15 15 13
2 15 13
6 3 9 13 0 9 13
9 13 13 3 9 1 11 7 9 13
7 13 3 15 9 7 13 15
4 3 9 15 13
7 16 15 13 11 13 15 3
3 13 15 11
5 13 15 7 3 13
13 9 15 15 13 1 9 9 15 0 9 13 1 15
12 9 15 9 15 13 7 15 13 15 7 13 15
8 9 15 15 13 15 0 15 13
8 7 15 13 13 1 9 9 15
5 15 7 9 12 13
6 13 9 9 16 13 15
3 13 15 11
8 0 9 0 13 15 1 9 15
6 1 15 15 9 15 13
3 13 15 11
9 3 13 13 1 9 15 16 15 13
2 9 13
31 16 0 13 9 1 15 9 9 13 13 7 3 13 13 9 15 9 13 7 13 1 9 15 13 16 13 16 13 9 9 13
9 16 3 13 9 9 15 13 13 15
24 16 3 13 3 16 15 3 13 13 9 13 16 13 7 13 16 1 15 13 9 7 15 1 9
4 13 3 15 13
5 7 13 1 9 15
5 11 3 9 13 15
9 15 3 15 13 11 1 0 0 13
5 7 0 13 1 15
14 13 3 15 13 11 1 11 1 9 11 7 11 9 15
17 11 3 13 15 13 9 9 7 13 9 15 9 15 15 9 11 13
6 13 3 9 1 15 13
5 9 6 15 13 13
5 13 3 11 13 15
13 3 3 13 16 13 3 3 13 1 0 9 12 9
6 3 1 0 13 9 15
4 13 1 11 3
3 13 15 9
10 9 3 13 15 9 13 7 3 13 3
2 13 11
5 3 12 9 13 9
11 16 3 13 9 13 16 9 3 13 1 15
4 11 9 15 13
7 7 13 16 1 9 13 15
4 13 3 9 15
5 9 16 13 0 13
6 13 3 11 1 9 15
8 0 3 13 16 1 9 9 13
3 11 13 13
14 7 13 1 15 16 13 16 3 13 3 7 13 1 15
7 13 3 15 16 13 1 15
3 13 3 11
9 7 13 15 12 9 3 1 9 13
8 13 3 11 1 11 3 9 12
15 0 3 1 9 13 1 11 7 11 16 13 15 1 9 15
4 11 3 3 13
5 13 3 11 1 11
9 9 16 13 3 9 15 3 13 13
3 13 0 11
3 13 9 15
3 13 15 11
8 13 16 13 1 9 1 0 9
5 15 13 9 7 9
9 15 13 1 15 3 16 0 13 13
12 7 15 15 13 7 13 1 15 3 13 1 0
2 13 0
14 3 9 15 13 16 15 13 11 9 9 15 1 9 13
12 7 16 0 13 13 7 13 11 9 15 9 13
5 9 13 7 13 15
6 3 3 13 11 1 9
10 7 13 3 1 0 9 3 13 15 11
24 9 3 15 13 1 15 1 9 7 13 15 16 13 11 16 3 13 7 13 13 13 15 13 16
6 13 1 9 16 13 3
16 11 3 16 13 3 13 11 13 15 13 1 9 15 7 13 15
21 11 3 3 13 15 13 7 9 15 13 1 15 13 13 9 7 13 15 0 7 13
3 3 13 15
4 9 13 7 13
4 7 13 13 11
3 13 3 9
4 6 3 13 15
5 15 3 13 1 15
13 3 13 0 15 13 9 0 13 16 3 0 3 13
8 13 3 9 7 9 13 13 15
2 13 9
8 13 15 11 9 15 15 13 13
3 9 3 13
3 0 3 13
3 13 15 11
9 3 13 15 16 16 13 13 9 9
3 13 3 9
19 15 3 13 16 3 15 13 7 1 9 15 13 13 16 13 16 15 15 13
6 0 16 13 9 0 13
3 11 13 3
17 7 3 13 15 13 13 13 9 7 9 9 7 9 0 9 13 13
3 13 11 15
5 13 15 7 13 13
15 0 3 1 9 15 13 1 11 7 13 15 13 13 1 15
13 15 3 1 15 13 1 9 7 13 15 15 13 11
8 15 13 16 0 9 0 9 13
18 16 13 15 3 15 13 1 15 7 13 0 7 13 15 7 9 7 9
12 12 3 1 15 11 16 13 9 9 0 13 15
20 15 13 15 3 7 13 16 13 15 16 12 13 9 1 9 7 3 0 9 13
8 0 3 1 15 3 0 3 13
29 7 16 13 9 9 0 13 16 11 13 13 1 9 7 3 3 1 9 7 3 16 9 9 15 13 13 13 1 12
8 1 0 3 9 13 16 13 15
25 11 3 3 3 1 3 13 1 9 7 13 1 9 1 9 1 9 15 13 11 7 3 13 1 9
8 15 13 16 3 13 1 9 0
16 13 3 9 7 9 9 16 16 15 13 3 13 13 16 13 15
15 11 3 1 12 9 9 13 11 3 13 11 13 15 13 11
16 13 3 15 9 3 7 11 13 11 3 12 13 1 13 1 15
17 11 3 13 9 9 9 0 0 13 9 11 7 13 9 15 9 15
7 7 9 13 13 1 9 9
12 13 3 12 1 9 15 11 11 15 13 15 13
3 13 3 11
6 0 3 3 13 15 1
5 15 3 3 3 13
23 13 3 9 0 1 9 16 3 13 7 13 3 1 11 3 7 16 11 13 15 13 1 0
19 13 3 9 9 16 3 11 13 16 0 1 0 13 1 9 7 13 1 11
25 1 0 3 9 0 15 13 1 9 0 1 13 16 13 11 11 13 9 9 7 13 1 15 7 13
9 6 0 15 13 1 9 9 9 11
4 13 13 9 11
8 6 9 15 13 13 1 9 9
18 7 3 13 13 11 3 13 13 16 0 13 13 1 15 7 0 13 15
18 9 3 13 9 15 13 1 15 3 11 13 1 9 7 13 15 1 0
12 3 7 1 13 15 9 16 13 15 13 0 9
7 9 3 13 1 15 3 0
4 13 16 15 13
13 13 3 9 15 1 0 15 13 16 13 1 9 0
14 0 3 13 1 11 15 13 1 11 11 7 13 15 13
4 9 13 11 13
6 11 3 7 11 13 11
5 11 3 13 15 13
6 13 9 16 13 9 9
4 6 6 13 15
7 16 3 13 13 0 9 13
19 15 13 9 15 13 15 7 15 13 9 15 1 0 9 1 9 0 13 15
15 16 15 15 13 15 13 7 3 13 15 3 7 9 15 13
8 16 15 15 13 13 15 9 15
3 7 15 13
6 9 13 15 1 9 0
6 7 3 13 1 9 0
5 13 3 9 1 9
5 7 13 7 3 13
10 9 3 15 13 7 13 13 9 13 13
2 15 13
4 9 15 13 13
9 3 1 15 9 0 13 7 1 15
4 3 9 13 9
12 7 15 16 13 13 1 9 15 13 1 15 0
8 0 3 13 13 15 9 13 13
3 13 15 9
9 15 13 1 9 16 11 13 1 0
4 7 3 15 13
4 13 13 9 9
4 13 3 15 11
17 13 16 9 13 16 3 9 15 13 7 15 13 1 9 13 3 13
10 16 9 13 13 1 9 16 9 9 13
11 0 13 13 11 7 13 7 13 15 1 15
18 16 3 0 9 13 1 15 3 13 1 15 16 9 11 9 13 15 13
5 9 15 13 9 15
6 7 9 9 15 13 13
8 3 3 13 13 16 3 13 11
8 3 7 1 9 0 13 1 15
10 7 1 9 3 13 16 1 9 3 13
8 13 3 9 9 3 3 9 9
5 11 3 13 7 13
14 15 13 1 15 3 13 1 15 7 1 15 15 13 15
9 7 15 13 15 13 15 15 13 15
15 15 9 1 9 13 16 15 15 13 1 15 1 9 3 13
13 7 16 15 13 9 15 7 3 13 15 3 13 15
12 15 13 15 7 3 13 9 15 13 15 13 15
32 9 15 13 13 0 13 15 1 0 9 16 15 1 15 0 3 13 13 7 15 13 15 9 15 15 9 13 15 13 7 15 13
8 7 13 16 9 15 9 0 13
10 15 3 15 13 3 13 15 9 3 13
18 1 9 3 0 9 13 11 16 13 15 9 16 13 1 0 9 1 9
11 16 13 15 15 13 1 0 1 9 13 15
45 7 9 13 16 9 3 13 1 9 16 13 15 11 11 11 13 16 15 13 15 9 1 9 7 16 1 9 13 7 1 9 13 13 1 9 7 13 9 15 7 16 13 9 13 15
16 3 13 9 1 9 7 13 13 9 9 7 13 9 15 13 13
5 9 15 15 13 9
5 13 11 7 13 15
6 15 15 13 15 13 3
3 13 3 3
3 13 15 11
6 3 13 15 9 1 0
3 13 11 15
4 13 15 11 11
3 13 15 11
11 15 13 13 3 13 16 13 7 13 0 0
7 7 15 0 13 7 3 15
7 13 3 15 13 15 13 15
2 3 13
4 3 13 0 15
4 13 15 13 15
3 15 13 15
3 7 3 13
2 13 3
16 16 3 15 13 15 9 9 7 9 3 15 13 0 0 13 9
13 9 3 13 15 16 3 15 13 15 3 3 15 13
4 6 6 13 15
8 3 7 9 0 15 15 13 0
8 16 0 13 0 13 16 13 15
5 3 1 15 15 13
4 7 16 13 9
10 15 13 15 1 9 13 1 15 9 15
13 3 13 15 16 13 16 13 16 13 13 16 15 13
4 6 6 13 15
9 15 3 15 13 13 15 15 15 13
7 1 0 13 11 13 13 9
5 7 13 13 7 13
10 6 6 13 15 16 12 1 15 13 15
13 13 3 13 12 1 9 15 1 9 11 15 13 11
8 13 3 0 11 11 7 13 15
5 15 13 1 15 13
3 9 15 13
2 13 11
7 0 13 15 15 13 9 13
8 7 1 13 9 13 11 11 11
8 7 1 9 3 13 1 0 11
4 15 13 13 3
9 0 3 15 13 13 1 15 13 15
7 16 3 13 0 9 13 3
3 13 3 9
5 16 3 13 13 11
11 3 13 13 9 9 7 9 13 13 1 15
14 16 9 13 13 1 15 7 9 13 15 1 15 3 0
4 7 3 13 15
17 13 15 7 3 13 9 3 15 13 15 3 13 13 3 15 13 3
8 3 13 15 16 3 15 13 3
13 1 0 13 15 16 15 9 13 16 9 13 1 3
4 13 15 11 11
3 9 3 13
2 13 11
8 3 15 13 3 13 15 3 13
3 13 3 3
5 9 15 1 15 13
2 13 11
5 9 15 1 15 13
4 6 6 13 15
7 3 13 9 16 15 3 13
4 3 13 9 15
7 13 1 9 7 1 15 13
7 1 9 9 15 9 0 13
22 7 16 13 7 13 15 9 3 13 7 13 15 1 15 0 16 3 13 15 3 15 13
8 7 3 15 13 13 7 9 13
3 13 15 11
4 9 13 3 13
5 7 3 13 9 13
3 13 15 11
7 15 13 9 7 9 7 9
7 15 13 1 9 3 1 15
3 13 15 11
7 9 13 15 9 7 13 15
3 13 15 11
10 0 9 15 1 13 7 3 13 15 11
6 15 13 15 13 3 9
3 3 15 13
3 13 15 9
10 9 15 15 13 15 1 15 0 3 13
11 3 13 16 15 1 9 7 9 1 15 13
5 3 1 9 0 13
4 6 6 13 15
20 15 13 1 15 9 15 15 13 3 15 13 7 0 0 13 16 15 1 9 13
13 7 15 13 1 9 15 0 13 16 13 9 1 9
9 16 15 13 15 1 9 15 0 13
30 7 15 13 9 7 15 9 13 15 16 13 15 1 1 0 9 9 15 9 3 13 13 16 3 13 15 3 7 13 15
12 15 3 13 15 16 1 15 13 7 1 15 13
3 13 1 15
8 3 0 7 9 15 3 3 13
10 15 3 13 15 16 15 13 7 15 13
19 1 0 9 15 13 16 15 13 1 9 15 7 15 1 15 7 15 1 15
12 15 13 9 15 7 13 15 0 13 15 13 15
9 7 15 13 15 7 13 15 15 0
6 13 15 11 3 0 11
13 9 15 13 13 16 15 13 13 15 0 7 3 9
21 16 15 13 15 9 15 13 7 9 15 13 15 7 1 15 13 7 9 1 15 13
8 15 3 13 15 9 15 3 13
13 7 9 15 13 3 13 15 7 15 15 13 15 9
7 0 13 13 15 1 15 13
3 9 13 15
4 9 15 13 15
7 3 3 9 13 15 13 15
7 3 13 9 15 3 7 13
5 13 7 13 1 15
14 16 13 15 13 3 16 13 1 9 16 9 0 15 13
11 7 3 13 15 16 13 16 16 13 13 13
11 13 3 9 9 0 7 1 15 3 13 15
15 7 3 13 9 16 13 9 7 3 9 13 15 9 3 13
1 13
2 13 3
4 15 13 9 0
20 15 9 1 15 3 13 9 13 15 7 15 15 13 9 13 15 16 9 3 13
10 3 15 0 13 1 9 15 13 13 15
21 3 9 3 13 13 9 1 15 3 0 16 13 1 9 3 3 15 16 1 15 13
5 15 13 9 15 9
18 15 13 1 15 7 15 1 15 0 13 9 0 16 1 15 15 13 13
21 16 15 1 15 3 13 13 3 3 9 7 13 7 13 15 7 1 9 13 7 13
16 16 13 1 15 7 9 15 1 15 13 15 13 13 7 13 15
14 1 0 13 13 9 15 16 9 0 13 7 13 15 9
4 13 1 9 15
14 0 13 13 15 16 9 15 1 15 13 7 9 15 13
10 0 13 9 15 16 13 3 3 13 15
13 0 0 9 15 13 16 9 15 15 13 1 9 15
10 15 9 15 13 16 13 15 15 13 15
12 3 3 13 15 9 16 9 13 15 13 9 15
14 15 3 13 9 16 15 15 13 1 9 15 0 13 15
29 3 15 15 13 7 15 13 15 7 13 15 16 13 7 9 13 7 9 15 13 16 15 13 9 1 9 15 13 15
9 16 1 9 13 9 15 15 13 13
16 16 3 1 9 3 13 7 15 13 15 1 9 3 13 15 9
7 13 9 15 15 15 13 15
6 3 13 9 0 9 15
7 16 15 13 13 3 15 13
7 16 9 15 13 3 15 13
14 7 0 15 13 15 1 9 15 16 13 15 15 13 15
10 16 3 13 7 13 13 15 9 3 13
7 15 15 13 3 9 15 13
13 16 9 3 13 1 15 15 15 15 13 9 3 13
11 3 3 7 13 7 13 7 15 7 9 15
11 7 16 13 9 15 1 9 15 13 13 16
4 9 15 13 3
31 16 3 13 9 15 15 13 15 1 9 9 9 15 1 9 13 0 9 13 1 15 7 15 9 13 16 1 9 15 1 13
7 0 13 13 15 16 3 13
4 1 9 13 15
15 7 0 13 13 15 16 16 13 9 15 13 16 15 13 15
11 0 3 15 1 9 3 13 16 15 1 13
14 3 3 13 1 15 15 15 13 7 15 1 15 13 15
2 3 13
10 7 16 0 13 13 15 9 13 9 15
5 7 15 9 13 15
5 13 15 16 15 13
7 16 3 13 13 15 1 15
8 1 9 3 16 3 13 1 15
12 1 9 3 16 1 9 13 7 3 3 13 15
9 1 9 3 16 9 9 0 13 13
10 3 0 13 15 13 7 3 13 13 3
11 16 3 13 0 9 9 13 15 1 15 9
17 3 3 13 1 15 3 0 7 15 13 13 7 15 13 13 13 15
6 15 15 13 9 15 13
3 3 13 16
16 0 7 3 3 13 15 7 3 0 7 13 15 16 13 1 9
7 13 3 1 9 15 1 3
22 15 13 0 15 13 15 0 7 3 13 15 7 3 0 7 13 15 7 16 13 1 9
2 13 3
5 15 13 0 15 13
3 13 15 13
10 13 3 11 16 13 15 13 7 13 15
7 1 0 13 1 15 16 13
9 6 6 13 15 16 13 7 13 15
3 9 3 13
9 15 3 13 7 9 15 13 1 9
9 9 16 13 9 13 16 13 9 15
7 7 15 3 3 3 9 13
8 3 3 13 15 7 13 9 15
7 7 9 15 15 13 1 15
8 7 1 0 9 15 3 13 15
9 16 15 13 9 1 9 15 13 15
8 3 3 3 13 15 1 9 15
8 13 7 13 16 9 15 13 0
15 13 9 3 3 3 1 9 13 15 7 3 1 9 13 15
6 0 9 1 9 15 13
10 7 3 13 15 16 15 13 9 1 15
16 0 3 9 13 15 16 15 15 13 7 13 16 15 1 9 13
7 13 1 9 7 13 1 9
4 13 15 9 15
4 6 3 3 13
14 3 13 16 13 15 7 3 9 13 15 16 15 15 13
7 1 0 13 16 1 9 13
3 13 15 11
2 3 13
15 6 13 9 7 3 13 16 13 15 1 0 7 15 0 13
9 7 3 13 0 16 9 15 1 13
4 1 9 9 13
3 15 13 9
4 0 13 13 11
6 7 13 9 1 9 13
3 9 13 9
23 13 9 15 16 9 15 13 15 3 13 15 9 15 9 16 15 15 13 15 13 15 9 0
16 0 13 3 9 0 16 13 15 0 0 9 7 15 13 11 11
5 15 15 13 1 9
9 13 9 15 9 15 13 15 1 9
6 15 13 7 15 15 13
4 7 9 15 13
10 3 13 16 15 15 13 15 1 15 13
7 3 9 15 13 15 13 15
16 7 15 13 7 13 3 16 1 15 13 7 13 16 15 15 13
4 15 1 15 13
13 3 1 9 13 7 1 0 15 13 15 16 15 13
5 7 13 13 1 15
16 7 3 3 13 1 9 7 0 1 9 13 7 15 1 15 13
16 9 0 13 15 1 9 15 15 13 15 16 13 12 3 3 15
10 16 13 1 15 15 13 15 1 9 15
4 15 13 15 13
11 7 15 1 0 13 3 9 9 16 9 13
5 3 3 1 15 13
14 7 0 13 1 9 16 13 9 15 13 1 15 3 0
11 1 9 3 13 3 3 15 3 13 1 9
4 13 15 1 9
4 9 15 9 13
11 3 15 13 1 9 3 15 13 15 1 9
14 7 1 15 15 13 15 0 16 13 3 0 13 1 9
45 3 1 0 3 13 3 7 3 1 15 15 13 13 1 9 15 1 15 16 15 12 13 3 15 9 1 15 7 15 1 15 16 3 0 1 15 12 13 16 9 13 16 15 15 13
15 7 15 9 15 13 15 13 15 16 13 12 3 15 12 13
27 9 15 13 15 13 16 3 15 13 3 0 13 15 1 16 13 9 15 15 13 15 16 13 15 1 9 9
4 15 3 15 13
7 7 0 13 16 15 15 13
21 7 0 13 15 9 15 7 0 13 16 9 15 13 15 1 0 13 7 15 1 0
22 0 16 13 11 13 13 1 9 15 1 9 11 3 13 9 1 15 13 15 7 9 15
17 13 3 3 11 15 13 15 0 9 16 3 11 13 3 1 9 15
19 11 3 16 13 9 7 1 9 7 9 9 13 3 1 9 7 9 7 9
2 15 13
2 13 15
3 13 15 11
2 15 13
9 13 3 3 11 15 13 15 1 15
12 3 3 13 15 15 13 13 3 7 13 1 9
4 3 3 15 13
3 0 3 13
2 11 9
2 13 11
7 16 3 15 13 13 0 13
6 3 13 9 15 13 16
8 15 13 15 3 13 1 0 15
7 11 3 11 13 9 13 15
5 13 3 9 9 11
4 13 3 11 11
4 13 9 1 9
8 9 15 13 15 9 3 13 0
6 7 13 15 1 11 3
9 13 3 9 11 15 13 9 9 0
14 13 3 11 15 9 13 9 16 13 12 9 13 1 9
13 9 3 0 13 0 9 7 13 1 11 1 9 9
6 11 3 13 1 9 3
11 13 3 9 15 15 13 0 9 7 13 9
3 7 13 11
5 13 3 11 9 0
2 13 0
2 3 13
10 13 3 1 15 3 11 13 7 13 15
11 9 3 13 11 1 9 15 7 1 9 15
3 13 15 11
5 15 3 13 13 9
18 15 3 13 1 9 7 1 9 3 15 9 13 7 1 0 13 13 15
3 15 15 13
6 6 0 13 15 13 15
3 3 13 9
3 13 15 11
8 16 3 13 13 9 13 1 0
6 16 3 3 15 15 13
8 7 13 15 11 13 1 11 9
8 13 3 11 11 13 7 13 15
3 13 3 15
2 3 13
11 13 12 1 9 9 0 15 15 13 11 9
8 3 15 15 13 1 9 1 0
4 3 3 13 11
4 7 3 9 13
7 13 3 11 1 11 1 9
3 13 3 3
12 7 15 3 13 1 9 16 3 13 7 13 9
6 15 9 13 1 9 0
4 13 7 13 15
9 16 3 13 0 9 3 15 13 15
4 13 3 15 11
9 13 15 15 7 1 9 15 13 15
4 13 3 15 9
5 15 3 13 13 15
11 3 9 11 13 15 13 13 15 13 9 13
4 15 13 9 9
3 7 13 11
12 1 15 3 0 0 13 7 15 15 13 1 15
2 13 11
4 3 15 9 13
7 9 15 7 9 13 15 15
2 15 13
7 9 15 3 13 1 9 0
7 3 3 15 9 3 13 3
4 13 3 15 11
4 3 9 13 15
2 13 11
6 15 13 16 9 13 15
15 15 1 0 13 13 7 1 0 13 1 9 16 9 13 9
3 13 15 11
3 15 13 9
6 15 15 13 1 15 9
10 13 3 9 15 16 12 13 15 1 9
6 13 3 13 15 9 9
4 13 3 15 13
4 3 0 7 11
7 3 3 13 11 11 7 13
9 7 9 13 9 1 9 13 9 15
5 7 9 0 13 15
3 6 9 9
4 7 13 15 9
7 13 3 11 3 7 13 15
13 6 13 15 15 3 16 13 16 1 15 15 9 13
3 7 13 15
2 6 9
9 16 3 13 15 9 7 9 13 13
1 13
3 13 15 11
5 13 15 15 7 13
7 15 3 3 13 1 15 9
13 15 9 13 7 1 9 13 13 16 9 9 15 13
8 16 3 13 11 0 9 3 13
5 7 13 13 9 3
4 7 13 1 11
3 3 13 15
4 13 3 15 11
3 15 3 13
2 13 11
11 3 13 9 1 15 15 16 15 13 13 3
8 3 15 13 15 15 0 9 13
5 3 13 11 13 15
4 9 3 13 13
7 16 0 13 3 13 9 11
9 11 3 16 13 0 9 13 3 11
4 13 3 9 9
3 9 3 0
3 7 13 9
3 6 9 15
3 0 3 13
1 13
1 13
3 9 15 13
2 13 9
5 3 13 9 3 11
7 3 3 13 15 0 16 13
5 13 3 11 7 13
27 7 13 15 9 13 1 15 15 13 11 9 3 11 3 15 13 7 1 15 15 12 3 7 3 0 3 11
9 13 3 7 9 11 7 13 1 9
3 13 3 13
22 0 3 9 0 13 9 16 3 9 13 9 3 13 13 11 7 13 13 3 3 7 3
5 13 3 11 9 9
8 13 13 9 9 7 16 15 13
3 9 13 9
2 13 11
3 15 13 13
17 9 3 16 13 15 13 9 15 7 13 12 9 15 9 9 7 9
8 13 3 9 0 3 13 1 0
4 3 9 13 13
5 13 13 9 15 15
6 7 1 9 15 13 9
5 7 9 3 0 13
16 13 3 1 9 11 9 15 7 9 9 15 11 11 7 11 11
13 16 13 3 11 9 7 9 13 15 13 13 9 15
4 9 6 9 15
3 6 9 15
12 3 13 11 16 3 15 13 13 16 13 9 13
1 13
6 9 3 13 13 9 0
10 0 3 9 0 9 9 13 13 9 15
6 16 3 13 11 9 13
2 13 13
26 9 3 16 9 13 16 3 13 1 9 9 9 13 3 0 9 0 9 13 11 16 13 15 9 7 13
3 13 3 9
27 1 11 3 16 13 3 13 15 3 0 3 13 15 9 7 12 9 9 9 15 13 7 3 13 9 7 9
5 7 15 13 9 13
5 7 0 13 15 9
10 7 0 13 16 0 13 16 3 15 13
7 13 13 3 0 16 9 13
5 7 3 15 9 13
4 13 1 15 13
22 1 0 3 13 11 11 1 11 3 16 13 9 11 0 3 1 9 9 16 13 9 11
6 13 3 7 13 9 11
18 13 3 3 11 15 13 1 11 9 3 13 9 9 7 9 3 9 12
15 13 3 9 11 7 13 15 9 1 9 3 9 9 13 13
8 13 3 1 9 3 13 13 9
11 3 3 1 9 9 16 1 13 9 13 11
13 12 3 9 11 11 13 3 16 3 9 13 1 9
6 7 13 9 13 1 9
17 13 3 7 13 1 11 11 7 1 15 9 15 13 11 7 13 15
11 13 3 11 7 0 15 9 7 13 1 9
16 13 3 12 3 7 0 15 9 13 3 11 7 13 0 1 9
7 7 16 15 13 13 13 9
31 13 3 11 11 13 15 7 13 1 9 7 13 9 13 7 9 15 13 1 9 15 3 1 9 13 7 3 13 1 12 9
11 3 3 13 3 0 9 15 13 0 1 9
4 7 13 7 13
10 3 3 13 9 16 13 15 1 0 13
8 13 3 3 1 15 3 0 9
9 16 3 13 13 15 7 13 1 9
19 7 13 12 9 1 0 13 12 1 9 7 12 1 9 3 13 13 9 11
3 9 15 13
3 13 15 16
3 13 9 15
5 7 13 3 13 15
10 0 16 13 13 13 3 7 13 11 13
6 7 3 13 16 11 13
3 9 15 13
7 0 13 16 9 13 13 15
14 9 16 15 13 15 13 15 3 13 15 7 15 15 13
3 13 15 11
1 11
4 13 0 13 15
1 9
3 15 13 9
6 3 3 13 1 9 15
8 13 3 1 9 15 7 13 15
13 13 1 9 15 7 9 15 7 9 15 7 9 15
6 13 11 11 13 9 16
6 13 9 7 0 13 15
20 16 13 3 3 9 0 12 9 7 9 13 13 3 13 9 1 9 9 13 11
7 7 13 1 0 7 13 15
2 9 15
6 13 13 3 9 13 9
4 13 3 15 3
2 9 15
8 3 13 15 9 3 15 13 15
7 0 16 13 13 7 13 15
3 13 9 0
5 15 13 9 13 15
4 15 13 13 13
2 13 9
4 0 3 13 15
23 16 13 1 9 15 9 9 7 13 9 15 1 9 9 7 13 9 15 1 9 15 3 13
13 7 1 9 12 3 13 9 15 3 7 11 1 15
10 13 11 9 13 7 13 1 0 7 13
2 9 15
3 3 13 11
6 7 13 13 0 7 0
5 9 15 7 9 15
3 13 15 11
4 16 13 15 13
6 0 15 3 13 7 13
18 0 3 7 15 9 13 11 1 9 9 15 15 3 13 13 1 9 0
20 0 3 13 13 16 13 16 11 13 11 9 9 7 16 13 9 13 1 9 15
3 13 3 3
25 13 3 11 11 7 11 15 13 11 7 11 15 13 1 11 11 7 9 11 7 15 1 9 15 12
2 13 13
2 13 15
5 13 3 15 15 1
6 7 13 7 13 1 9
5 7 0 9 15 13
7 3 3 13 9 16 11 13
4 13 3 15 11
4 9 3 9 13
1 3
2 13 15
7 13 1 9 9 9 7 13
2 13 3
8 13 3 9 0 15 13 11 11
2 9 13
18 11 11 16 13 16 9 13 9 13 15 13 3 0 7 13 15 1 9
5 15 3 9 9 13
13 3 3 13 1 9 13 9 13 7 9 13 7 9
3 13 15 11
6 13 1 9 15 13 3
8 3 16 0 13 3 13 13 9
3 13 15 11
1 13
1 13
13 7 15 13 13 13 15 15 15 13 13 16 9 13
11 0 3 3 13 13 11 9 16 13 1 0
7 16 3 13 13 11 11 11
2 13 15
7 3 9 15 13 16 13 15
2 13 15
3 13 9 15
3 13 15 3
4 11 11 13 15
7 3 9 15 13 16 13 15
3 13 9 15
3 13 15 3
4 11 11 13 15
7 13 13 11 16 13 15 3
2 13 15
3 7 13 15
4 9 15 15 13
3 13 9 15
4 6 6 13 15
9 16 13 0 13 15 7 13 3 13
15 16 3 13 13 9 15 7 15 15 13 7 13 3 3 13
9 0 3 13 13 15 9 13 13 9
6 7 0 16 13 13 15
2 13 15
19 13 11 13 0 9 15 13 11 13 15 7 13 1 9 1 9 15 7 13
7 0 3 16 13 11 13 11
4 9 0 3 15
3 13 15 11
10 16 3 15 13 13 16 13 15 1 15
3 15 15 13
11 13 3 9 0 1 9 16 9 0 3 13
8 7 3 13 15 11 3 13 7
10 16 3 15 13 13 16 13 15 1 15
8 13 3 3 15 0 15 13 11
15 15 16 13 1 0 3 0 13 9 13 15 15 13 13 9
1 6
27 0 3 9 13 1 15 6 11 15 13 11 13 7 13 3 1 9 15 13 9 1 9 0 15 13 13 13
22 15 7 13 15 0 0 1 9 15 1 0 9 1 9 12 13 15 7 13 1 9 9
17 7 13 13 15 1 11 3 13 7 13 9 9 15 13 1 9 15
5 3 11 3 13 9
6 3 15 13 13 15 13
3 13 3 15
13 3 13 15 13 9 7 9 15 9 13 1 15 9
25 7 13 9 13 9 0 1 15 7 13 15 9 1 11 7 1 15 11 7 11 7 3 1 0 9
8 7 16 0 13 13 0 13 13
7 7 9 13 15 1 9 15
18 16 13 1 9 13 0 6 12 9 13 1 0 1 9 0 15 3 13
17 0 11 15 13 13 1 15 1 9 3 13 3 13 15 13 1 9
16 3 13 13 11 1 9 15 13 11 15 13 1 11 9 13 9
16 0 15 13 13 3 1 9 1 9 7 11 9 11 7 9 15
10 7 1 9 0 13 11 1 0 9 13
7 13 3 9 9 3 3 12
21 9 9 13 13 9 15 13 9 0 1 9 11 1 11 15 13 9 15 15 13 11
11 3 13 13 1 15 7 13 13 9 9 0
6 7 13 13 15 9 15
15 7 0 13 13 15 13 11 3 16 13 9 0 9 15 11
4 0 13 9 9
11 13 9 15 13 7 3 13 15 13 1 15
5 7 9 15 13 15
42 13 3 1 0 9 15 15 1 13 13 1 15 9 15 13 7 13 1 15 9 11 13 1 9 11 3 1 9 15 13 13 1 15 9 9 15 15 1 13 12 1 0
13 7 13 12 11 15 13 11 15 13 13 11 7 11
29 15 9 15 9 13 15 13 15 13 1 0 12 12 13 9 9 0 7 9 1 15 13 13 11 16 13 1 9 15
9 7 13 9 15 7 13 9 1 11
6 7 13 13 1 12 9
11 7 16 13 9 9 13 15 3 1 0 9
12 7 13 0 13 9 3 9 13 7 1 0 15
17 7 13 13 15 9 0 7 13 13 15 9 3 9 0 13 13 0
15 13 3 1 11 13 0 9 0 1 15 9 15 1 9 13
6 13 3 15 7 13 13
8 3 15 6 0 15 13 9 13
11 7 3 15 13 15 9 15 1 15 13 13
44 9 7 9 7 9 7 15 13 11 7 11 7 11 11 7 11 11 7 11 11 7 9 11 15 13 1 11 7 9 0 9 3 7 9 9 7 9 13 13 15 15 9 9 9
8 13 3 15 7 13 1 3 13
5 15 3 13 13 16
4 9 0 13 0
16 9 0 7 15 13 11 0 0 15 0 13 7 9 13 9 15
13 3 3 3 15 13 0 0 13 16 13 9 9 0
9 7 0 13 15 13 13 1 9 11
5 7 13 1 0 9
2 13 9
24 13 1 9 15 1 15 9 7 13 9 15 7 9 15 7 0 15 9 13 7 0 15 9 13
17 7 13 9 1 9 3 7 9 1 9 3 9 7 9 7 9 9
2 7 13
7 15 15 13 9 9 0 13
5 9 9 13 9 0
36 11 9 9 13 1 9 1 15 9 7 9 7 9 15 13 1 0 9 1 0 15 3 15 13 0 0 9 7 9 9 13 1 9 0 13 13
14 15 9 13 13 9 9 3 16 0 13 13 0 1 15
5 11 3 13 1 15
12 13 9 1 15 3 16 1 0 15 13 16 13
5 0 13 15 9 9
6 13 15 9 1 9 15
27 9 9 13 3 13 1 15 1 9 11 16 7 13 13 7 13 13 7 9 15 13 1 15 3 1 0 9
39 9 3 16 13 7 13 16 9 13 13 0 9 1 9 9 15 13 1 9 15 13 13 13 1 9 11 16 3 7 13 13 1 9 3 7 9 15 13 9
9 0 11 13 9 15 15 15 9 13
18 9 3 9 13 7 9 9 0 13 1 9 13 0 15 15 13 7 13
6 3 3 11 13 1 9
3 13 3 15
11 13 1 0 15 16 13 9 15 9 9 15
19 3 3 13 15 9 11 16 7 9 15 7 11 9 13 0 11 15 15 13
13 0 13 13 13 9 7 13 1 11 7 1 0 9
4 15 13 9 9
7 11 3 1 0 9 13 13
12 7 13 15 15 1 9 11 11 1 9 9 15
5 7 13 9 0 9
17 15 3 13 9 7 9 15 7 15 15 3 13 15 13 9 9 15
7 15 3 13 9 15 13 13
10 7 13 13 1 0 9 9 3 12 12
12 13 3 13 1 9 9 7 9 9 9 7 9
5 13 3 15 9 9
16 0 3 9 7 9 1 9 13 1 11 7 9 13 0 1 0
10 15 3 15 13 13 3 7 13 15 0
12 9 7 9 13 7 13 0 15 3 15 9 13
10 9 3 13 15 0 13 3 1 15 0
11 7 15 9 15 13 0 1 9 9 15 13
16 15 13 3 1 9 9 15 13 0 16 13 9 1 13 1 9
14 15 16 13 11 7 11 13 13 1 9 13 16 9 13
8 13 3 1 15 11 1 11 13
3 13 1 15
11 3 0 13 1 15 13 15 15 13 1 15
6 9 7 9 3 13 15
6 15 3 13 0 15 13
15 7 13 15 9 0 13 15 7 3 13 13 9 15 7 9
5 7 13 13 7 13
12 7 13 1 0 1 9 13 7 13 7 13 9
9 7 13 15 9 15 13 7 13 9
14 13 3 0 16 15 13 15 1 9 13 1 0 9 9
17 16 13 3 11 7 11 13 15 9 1 15 1 9 15 13 11 13
6 13 3 11 13 1 9
18 9 9 15 13 1 0 7 15 15 13 16 15 9 7 9 13 0 13
12 15 3 0 7 0 13 7 13 9 9 13 15
13 9 3 9 13 15 9 13 1 0 15 15 9 13
13 7 1 9 9 15 0 15 13 7 13 13 9 15
14 7 9 15 1 15 13 13 0 9 0 1 9 15 15
13 9 3 15 13 1 9 15 9 13 11 15 13 3
46 13 3 7 13 16 13 15 9 16 16 13 9 9 1 9 9 7 13 15 15 13 13 15 11 11 15 13 9 3 13 3 1 9 9 15 15 13 13 9 1 9 0 15 1 9 9
4 11 3 13 16
11 9 15 13 9 9 15 1 9 15 3 15
2 13 3
10 15 9 15 3 13 9 0 13 1 9
14 7 15 9 1 11 7 3 15 13 13 7 13 9 0
8 7 1 9 15 13 15 9 9
17 15 3 9 13 9 15 13 15 13 15 16 13 15 15 1 9 15
23 13 3 0 1 9 13 9 7 9 9 7 9 13 16 13 9 7 13 1 11 9 1 0
12 7 13 1 15 9 7 13 15 1 9 1 0
4 13 3 3 9
7 7 13 13 9 9 12 12
31 13 13 3 1 0 16 13 9 15 7 0 7 9 1 11 7 11 9 9 7 11 7 11 7 11 7 3 13 1 9 0
10 1 15 9 7 1 15 9 13 0 15
8 3 11 13 9 0 13 1 15
47 9 9 7 0 16 15 3 13 1 9 9 0 1 15 0 0 13 13 0 13 15 15 7 15 9 11 16 1 9 11 11 9 15 15 13 15 9 13 1 0 1 0 0 13 1 15 0
15 0 13 9 15 13 13 1 15 13 15 13 13 1 9 9
7 7 3 13 1 15 15 9
16 3 7 3 9 15 13 1 9 13 9 1 15 13 15 0 13
12 9 3 13 13 1 15 15 13 13 15 13 13
5 7 13 1 3 13
4 15 13 9 0
17 3 3 0 9 13 13 1 15 15 13 1 11 0 7 3 13 13
16 7 16 3 13 1 9 13 15 16 3 13 1 9 0 15 9
13 7 13 15 13 16 3 13 3 7 13 1 9 11
8 11 3 7 11 13 13 1 15
12 16 0 13 1 9 9 15 3 13 3 9 13
13 9 3 13 3 12 9 1 15 13 13 9 0 9
16 13 3 13 1 15 7 13 15 15 1 15 9 9 7 0 13
10 15 16 13 3 13 9 1 9 7 13
26 9 15 15 13 9 7 9 7 9 7 15 15 1 15 13 15 9 0 1 9 9 15 11 9 15 13
8 3 13 9 7 9 13 13 0
14 13 9 9 7 9 13 1 12 1 9 7 1 11 15
30 13 3 3 1 9 0 1 0 9 15 11 15 13 11 7 11 11 1 9 7 9 11 13 15 9 15 7 9 13 13
35 7 3 9 13 1 9 15 7 13 9 15 1 15 9 13 9 15 1 15 16 9 15 13 9 7 9 7 9 13 1 9 0 9 15 11
12 7 13 13 15 9 0 7 13 9 9 1 9
8 9 3 13 13 9 7 9 12
15 3 7 15 15 15 13 15 15 13 13 7 13 0 15 0
10 7 9 0 13 9 9 9 11 11 9
7 7 9 0 13 1 15 0
8 3 7 3 15 13 13 1 0
18 3 3 9 9 7 9 13 13 13 9 15 15 13 7 13 1 9 9
7 13 3 0 3 15 9 13
8 7 13 9 15 1 9 9 13
3 13 3 11
15 11 3 13 11 9 15 13 15 9 0 7 13 1 9 9
10 3 13 15 13 7 13 1 15 13 9
7 3 13 1 9 15 0 9
6 3 13 13 9 7 9
8 13 3 11 0 9 13 7 13
8 13 3 0 13 15 7 13 13
4 13 3 15 11
6 13 15 16 0 9 13
3 3 0 13
2 3 0
4 11 3 1 15
7 15 3 13 15 13 9 9
7 3 13 1 9 15 7 13
6 13 3 0 13 0 0
14 7 13 13 9 0 1 0 9 7 1 15 15 13 0
11 1 9 3 9 13 9 7 9 0 1 9
7 7 13 3 15 1 9 11
7 0 3 15 13 13 15 0
4 7 13 15 9
14 13 3 3 9 0 9 11 13 0 7 13 1 9 0
3 15 13 15
17 13 3 9 9 7 15 15 1 0 13 15 13 9 9 13 13 9
12 9 3 9 1 9 13 9 9 7 13 15 13
11 13 7 13 13 1 9 9 15 9 9 0
9 15 16 13 13 9 1 9 7 13
16 13 3 9 9 7 15 1 15 13 13 9 7 15 0 9 11
13 16 13 3 9 7 13 9 3 13 0 13 13 13
12 9 3 13 13 1 15 9 7 9 13 1 9
5 13 3 15 3 13
15 3 13 3 0 9 9 9 7 9 9 13 1 0 15 13
13 6 9 15 13 1 9 13 1 9 13 7 13 9
10 3 13 9 1 9 7 13 0 1 9
5 13 3 9 16 13
6 7 13 15 9 9 13
14 13 13 15 16 13 1 9 0 7 6 13 11 9 15
8 7 13 13 1 15 9 9 0
6 13 3 11 7 9 13
6 13 13 9 3 3 9
15 0 9 9 7 9 13 9 15 1 13 9 11 7 9 9
15 7 15 13 9 0 9 7 9 0 15 13 9 15 13 15
23 13 3 15 1 9 9 9 11 9 9 0 0 9 13 3 1 0 9 13 13 7 1 0
10 9 9 13 15 1 9 0 15 13 13
16 1 0 3 9 13 11 13 13 15 15 15 13 9 9 3 12
15 15 13 13 7 15 15 13 15 13 13 7 13 13 1 9
13 1 0 13 11 9 1 9 9 7 13 9 1 15
10 3 15 13 7 15 3 13 15 13 13
7 13 1 9 0 7 13 0
15 16 3 1 9 13 3 13 13 15 16 3 3 9 13 13
3 13 3 0
13 7 13 9 13 13 16 13 1 9 11 7 13 15
17 7 0 3 13 13 1 9 9 16 0 13 13 1 9 11 9 13
15 15 3 9 1 9 7 1 9 3 13 13 7 13 11 11
21 1 9 3 0 13 9 9 13 13 9 9 1 9 3 16 13 1 9 0 9 15
6 13 3 12 9 9 13
8 15 3 9 7 9 9 13 13
6 7 13 9 1 15 9
23 7 13 11 9 0 9 7 9 0 7 11 7 11 7 11 7 11 7 11 7 11 9 0
5 0 13 1 9 9
5 7 13 13 15 9
11 7 9 9 13 7 13 9 9 1 11 3
6 0 3 9 9 13 9
13 11 3 0 9 7 9 13 9 7 9 0 1 9
9 7 3 13 13 9 7 9 15 13
15 3 13 9 15 13 15 13 15 13 9 9 1 11 7 9
7 13 3 9 7 0 7 9
13 7 13 13 15 7 13 1 9 7 13 9 0 13
11 9 0 3 13 13 9 1 9 0 7 9
18 13 3 15 13 16 11 9 0 13 9 0 7 13 9 15 13 15 11
14 7 13 15 15 15 13 1 9 13 9 15 3 9 9
9 13 3 9 9 16 0 3 15 13
18 9 9 13 9 15 11 16 13 1 11 16 13 1 11 7 13 1 0
15 13 1 9 15 7 1 9 15 7 13 1 9 15 15 13
9 3 13 1 9 9 7 13 1 11
17 7 3 16 13 13 9 15 13 0 1 9 0 1 15 3 15 13
10 7 3 13 0 9 1 15 3 9 9
16 7 13 13 0 15 1 9 7 9 15 1 15 16 3 13 9
5 13 13 3 9 16
18 7 9 15 13 13 15 13 9 7 1 0 13 7 13 15 1 9 0
9 7 3 13 11 7 13 15 9 0
3 7 11 11
4 7 11 12 9
7 7 9 13 11 13 1 11
23 7 13 9 1 15 7 13 15 1 15 9 15 7 13 15 9 7 9 1 9 11 13 11
11 7 13 15 9 1 11 7 1 15 9 15
12 16 13 3 11 13 9 1 11 13 9 15 3
15 7 1 0 13 13 11 1 9 15 7 13 13 11 9 15
5 7 13 11 1 11
7 7 13 13 15 7 9 15
20 7 13 13 1 11 7 13 13 1 9 15 13 11 9 9 1 9 11 9 11
27 16 13 3 9 9 15 13 13 9 11 13 9 7 13 13 1 11 16 13 9 15 1 11 15 3 13 11
12 0 13 9 15 13 9 16 13 9 15 16 13
9 15 13 13 12 9 1 9 9 15
13 13 3 0 13 15 9 11 7 13 15 15 1 9
16 7 13 13 11 15 9 9 7 13 0 1 9 7 1 9 15
17 7 16 13 15 9 13 13 0 7 13 9 15 15 9 13 13 9
12 13 3 13 9 16 9 1 9 15 13 9 0
4 3 0 3 13
6 0 3 9 13 0 13
3 9 9 13
4 3 15 13 15
8 15 3 9 13 0 13 15 13
8 15 15 13 9 7 9 1 15
6 13 3 11 1 9 0
11 7 13 13 9 1 9 11 3 13 9 12
15 7 13 9 12 13 0 1 9 9 11 9 1 9 9 9
9 7 13 0 16 13 13 13 9 9
12 15 9 9 15 9 11 7 9 11 7 9 11
6 13 3 11 3 13 13
4 13 3 0 9
4 13 9 9 15
17 13 13 9 9 15 15 13 1 11 7 9 15 13 7 13 13 15
8 7 3 13 7 13 15 1 11
19 0 13 0 13 9 7 9 1 9 11 7 1 0 9 7 1 9 9 12
7 0 13 11 15 13 9 11
9 9 15 13 9 1 9 15 3 15
20 0 13 15 13 1 9 1 9 1 9 15 13 15 1 9 11 7 1 9 15
6 15 13 9 9 13 15
17 15 13 13 9 15 7 13 7 13 13 9 15 1 11 13 1 11
14 11 3 0 15 13 15 1 9 11 13 15 13 13 15
9 13 3 9 7 13 15 13 9 9
6 3 13 13 1 9 9
12 3 9 7 9 13 15 9 12 1 9 9 11
14 7 13 9 11 7 9 9 15 11 9 15 13 13 15
5 7 13 15 1 11
19 9 9 13 9 15 1 9 3 13 13 1 11 16 13 0 1 9 15 13
34 15 3 13 13 9 15 1 11 1 9 9 15 13 9 1 9 9 15 3 1 9 11 15 13 9 1 9 7 13 16 13 9 9 11
3 3 9 13
4 9 15 9 13
5 9 3 9 9 15
12 15 9 13 15 13 9 7 15 9 9 15 13
6 3 9 15 13 0 15
12 0 9 7 0 9 7 9 15 3 9 0 13
5 3 9 15 3 15
7 15 9 3 13 13 9 15
9 15 13 9 1 9 9 7 3 13
11 13 3 0 13 9 15 7 13 9 1 15
18 16 3 13 0 9 0 13 1 9 13 9 9 7 11 13 1 0 9
2 7 13
11 6 13 9 13 7 9 9 1 0 13 9
13 13 3 9 0 13 9 15 7 9 13 3 1 15
6 7 13 15 1 9 13
11 7 9 13 9 15 1 9 9 15 13 11
6 13 3 9 13 9 0
6 9 3 13 0 0 9
5 7 16 0 13 13
6 11 3 13 13 9 15
24 13 13 3 1 0 9 9 0 1 9 15 13 11 7 15 13 13 1 9 11 7 11 1 9
11 13 3 11 9 0 7 13 9 0 1 0
15 11 3 13 9 1 9 13 7 13 9 7 9 13 1 9
9 11 3 13 1 9 11 13 0 11
11 0 3 15 15 13 9 0 13 9 0 13
7 0 3 9 7 0 13 13
8 13 13 3 0 9 1 0 9
19 9 3 15 9 11 15 3 13 1 9 9 13 9 11 13 13 15 15 0
9 15 13 15 1 0 3 1 0 13
7 0 13 9 9 15 13 0
16 16 3 13 11 13 1 9 9 7 9 11 11 13 9 7 9
5 3 11 3 0 13
9 13 3 9 7 9 0 13 13 13
18 16 3 13 9 15 13 11 16 13 11 9 9 13 1 0 11 7 11
10 15 16 13 13 1 15 16 13 9 0
14 3 3 1 15 0 13 7 13 3 13 1 9 9 11
9 3 13 9 1 0 7 13 9 0
12 13 3 15 0 9 16 15 13 9 13 9 0
5 11 3 13 1 15
13 9 15 15 1 13 1 9 16 9 9 13 9 13
8 9 3 15 3 13 0 1 9
7 9 3 13 1 0 9 15
11 7 13 9 16 3 13 15 0 9 9 15
10 1 9 3 9 7 9 9 13 15 13
14 13 15 1 15 1 9 16 15 13 1 15 0 15 13
15 7 0 3 13 7 13 9 9 13 11 7 0 9 9 13
8 9 3 9 13 13 1 11 13
13 13 7 13 1 0 1 9 15 13 1 11 1 11
3 7 13 13
19 7 6 9 0 9 0 11 9 11 15 13 1 15 9 15 13 13 1 11
10 7 13 13 1 9 15 13 7 9 11
7 13 7 13 15 1 9 0
10 13 3 11 13 0 13 11 9 7 13
5 13 3 13 15 13
2 15 13
8 7 3 13 16 3 15 13 15
7 9 3 9 15 13 13 0
6 3 9 1 9 13 13
6 1 9 9 15 13 13
4 9 0 15 13
6 3 13 1 9 9 15
5 13 3 9 11 13
2 13 15
11 1 15 9 13 0 1 15 7 1 15 15
9 7 16 13 1 9 13 1 15 9
2 6 9
4 15 13 15 13
4 7 13 13 9
11 7 13 15 1 9 11 7 9 7 13 15
15 16 3 13 1 9 9 9 13 11 7 3 3 13 15 9
6 13 3 1 9 15 13
14 11 3 13 13 1 11 7 13 13 9 0 16 13 11
7 7 3 13 15 9 1 9
8 7 13 1 9 13 9 13 15
5 11 11 15 15 13
2 15 13
3 15 13 9
2 7 0
6 15 13 11 15 15 13
12 7 13 7 13 9 7 13 15 15 15 13 13
10 13 3 11 1 9 13 7 9 15 13
7 1 9 3 0 13 13 11
12 7 13 12 9 3 13 7 3 13 3 7 13
7 13 3 15 9 11 9 11
7 7 13 1 0 1 9 9
1 11
3 3 0 13
3 6 15 9
8 7 13 1 9 11 11 9 0
3 6 3 13
13 7 13 9 11 9 13 7 13 15 9 16 9 13
3 13 3 11
14 9 13 1 0 1 9 0 15 0 0 15 13 1 11
13 7 3 13 9 1 9 9 13 15 15 13 9 15
5 13 3 1 15 9
11 15 3 13 0 15 13 15 1 9 15 13
5 7 13 15 9 13
19 11 9 9 13 15 11 15 13 15 1 9 15 13 16 13 7 13 9 0
11 7 3 13 1 9 15 3 9 7 9 13
4 7 13 13 13
6 7 16 13 9 13 13
10 13 3 1 9 15 13 11 1 9 15
7 13 3 15 15 13 7 13
12 3 0 13 15 13 1 11 15 15 13 9 0
15 11 3 3 13 7 13 9 15 13 11 13 16 0 13 11
11 16 13 3 9 0 9 13 9 16 15 13
7 0 3 13 13 11 9 15
10 13 3 3 9 9 7 9 16 15 13
12 13 3 9 15 9 1 9 13 15 13 1 9
7 11 3 13 0 13 1 9
22 7 13 0 3 1 9 13 9 7 16 13 13 15 7 3 1 11 3 13 1 9 11
15 7 13 1 0 13 7 13 1 11 7 3 13 1 9 9
5 0 3 13 13 15
10 15 1 13 9 13 15 11 7 13 11
22 9 3 1 0 11 7 11 7 11 13 9 7 13 13 1 9 9 7 9 0 9 13
14 13 13 3 11 16 13 0 13 3 1 0 15 13 11
4 7 13 0 11
5 11 13 15 11 11
4 13 7 13 15
3 7 3 13
5 15 13 13 1 9
12 1 11 3 13 15 9 9 11 15 13 13 11
9 0 13 0 9 0 7 9 15 13
7 15 16 13 13 15 1 9
20 16 3 3 13 11 1 11 9 13 16 11 13 1 15 13 12 9 1 15 13
6 3 13 13 3 1 15
6 13 3 11 13 1 0
7 7 16 13 13 0 1 9
8 13 3 15 3 11 13 9 13
5 7 13 1 9 13
5 3 0 13 9 15
4 7 13 11 13
6 13 3 0 9 13 15
9 7 16 13 0 7 9 13 15 0
7 0 3 13 13 1 0 11
5 7 13 0 1 9
29 9 3 15 13 1 11 9 11 9 9 15 13 11 0 7 13 9 1 15 9 15 13 9 0 9 7 13 9 3
1 11
7 3 0 13 15 9 13 13
3 15 13 9
3 13 3 0
11 9 15 7 9 15 13 1 9 1 9 9
13 7 3 13 9 1 11 7 13 11 15 15 13 11
11 0 13 1 11 15 9 15 13 9 1 9
18 0 3 9 9 0 13 7 13 9 13 11 1 0 16 13 1 9 0
5 7 16 13 13 13
8 13 3 15 13 1 15 9 9
29 7 13 9 13 7 13 9 15 3 9 0 12 9 13 1 9 1 9 1 15 13 15 9 7 13 9 7 9 9
6 7 13 13 9 1 15
2 13 11
4 7 13 7 13
3 13 3 11
6 7 9 3 3 1 15
7 15 9 13 16 15 0 13
6 0 3 13 13 1 3
7 7 3 13 13 9 1 9
24 7 16 1 15 13 11 15 13 9 15 13 6 9 15 13 13 1 11 13 9 11 13 1 9
12 7 16 13 13 16 11 15 13 11 3 13 9
8 11 3 13 1 9 13 9 15
5 6 9 12 13 15
5 6 15 13 15 13
6 15 9 13 1 15 13
2 15 13
29 11 9 9 0 7 13 9 7 9 13 1 0 9 9 9 13 1 9 0 13 15 1 9 15 7 13 9 1 15
5 13 3 15 13 9
17 0 3 9 13 13 13 1 15 7 15 1 9 1 11 13 13 15
5 0 3 9 13 11
3 7 13 13
5 11 3 13 15 13
1 13
5 3 15 0 9 13
10 7 13 1 0 13 7 13 0 15 13
4 13 7 1 0
12 15 13 3 13 13 9 0 13 7 13 1 9
6 1 15 1 9 13 13
2 13 3
3 7 11 13
26 1 3 0 9 3 1 0 9 13 13 9 0 1 9 15 7 6 9 13 1 15 1 9 0 7 13
13 11 13 13 9 15 7 9 15 13 13 1 9 9
10 13 3 1 11 7 13 11 15 13 11
8 0 13 1 9 11 9 1 9
5 7 15 3 13 13
16 3 3 15 15 1 9 15 13 13 15 15 15 13 13 1 9
5 13 3 11 9 13
9 9 13 9 11 13 9 1 11 11
4 0 13 15 9
18 15 13 15 13 13 9 1 0 11 13 3 1 11 1 9 15 13 11
25 11 1 11 3 13 15 9 9 0 7 9 15 13 13 7 13 15 13 1 9 16 9 13 1 0
6 15 3 13 13 1 9
29 0 9 13 0 9 7 13 15 0 13 3 15 9 7 9 13 1 9 15 15 13 7 13 1 0 16 13 1 0
19 7 13 15 13 9 7 13 16 15 13 15 13 13 1 9 9 0 7 0
16 0 15 9 9 13 9 9 13 1 9 15 15 15 13 1 15
18 7 13 1 9 0 15 13 1 11 16 3 1 9 9 9 0 13 13
8 13 3 0 13 9 7 13 9
3 3 13 11
8 7 13 15 1 9 11 11 13
7 3 13 15 16 13 15 9
15 13 3 9 7 9 15 13 1 11 16 3 9 13 9 9
14 16 13 3 11 1 11 13 1 0 15 13 1 9 13
10 3 13 1 9 9 13 7 13 1 0
28 15 13 1 9 11 13 7 13 1 9 9 9 13 9 15 3 9 0 12 9 13 1 9 7 13 3 1 15
15 1 15 13 13 7 13 0 9 7 9 7 9 7 9 9
5 13 11 13 7 13
2 13 3
11 3 9 16 0 7 0 3 13 1 9 15
6 13 3 9 3 1 9
7 15 9 13 15 3 0 13
6 0 3 13 13 1 3
16 7 6 3 12 9 13 1 9 1 15 13 13 1 11 1 15
14 13 3 15 1 3 12 9 0 7 13 13 1 9 9
13 13 3 15 3 13 9 1 9 15 13 7 13 15
22 13 1 11 7 13 11 15 13 11 15 13 15 9 1 15 0 13 15 7 0 9 15
15 16 3 13 13 13 9 0 1 15 3 3 1 15 1 9
7 13 13 3 9 9 3 13
4 11 3 13 9
5 15 3 13 9 0
4 7 13 9 13
8 3 3 9 9 9 1 9 13
26 7 0 3 15 13 13 1 9 15 13 13 1 11 13 3 11 7 11 7 11 15 13 9 3 0 9
20 13 3 15 1 15 9 0 7 0 15 16 13 11 13 3 1 9 13 9 11
6 7 13 9 9 1 15
8 0 7 9 13 13 13 1 9
11 13 3 9 1 9 9 15 13 11 1 0
5 7 13 11 3 11
18 7 13 15 9 9 13 1 9 16 13 9 0 7 0 9 0 7 9
6 7 13 13 9 0 9
7 13 13 3 11 16 13 11
5 15 16 13 13 11
7 7 9 0 13 13 1 9
11 7 13 9 0 3 16 13 3 11 9 0
9 1 0 3 9 13 1 11 9 11
22 7 13 12 1 15 9 11 13 1 9 9 0 13 1 0 9 9 15 13 13 1 11
12 0 3 9 13 11 9 9 16 13 15 1 9
6 13 3 11 9 11 9
9 13 3 16 13 9 13 13 7 11
4 13 3 9 9
18 15 16 13 13 1 9 13 12 9 9 13 15 13 1 9 13 15 9
6 7 11 3 13 1 9
11 9 3 13 1 9 1 9 1 9 1 15
6 7 9 1 9 13 9
7 13 7 9 11 13 15 13
2 13 3
6 7 13 9 1 9 15
5 13 3 9 1 15
6 13 7 13 15 9 15
3 7 13 3
7 13 15 9 15 7 13 15
12 7 13 13 7 13 16 0 13 15 13 1 9
14 13 3 0 7 0 9 13 1 9 0 15 13 1 9
5 15 3 13 13 15
5 7 13 13 9 12
6 7 3 13 9 1 15
6 7 11 1 15 13 13
18 13 7 13 1 9 11 9 11 15 13 13 11 3 13 0 13 7 13
11 13 3 15 9 9 13 9 1 13 9 11
18 7 16 13 9 11 1 9 3 13 9 7 3 13 13 13 11 1 9
1 13
6 0 3 13 3 15 13
3 0 3 13
3 9 15 13
7 16 3 13 13 15 7 13
15 13 3 15 9 16 13 13 3 9 13 15 1 9 13 7
5 13 11 7 9 0
6 7 13 13 1 15 9
15 11 3 16 13 15 7 3 13 9 13 1 9 13 15 13
9 13 7 1 11 1 11 3 13 13
6 13 3 13 9 7 9
14 13 3 9 11 13 9 0 13 1 9 7 13 1 15
3 9 3 13
5 9 9 7 3 9
12 3 3 13 15 9 9 3 16 3 13 9 9
5 7 13 1 9 13
16 11 3 7 11 13 13 1 11 13 9 13 11 15 13 13 11
30 13 3 1 9 15 13 11 9 7 9 1 15 11 7 11 15 13 11 7 11 0 7 11 15 13 11 9 0 7 11
10 13 15 11 7 11 1 9 15 13 15
10 3 13 7 13 13 7 15 9 13 0
9 7 15 3 13 1 9 0 13 11
4 7 3 13 11
10 7 16 13 11 13 9 9 1 9 9
6 13 3 3 11 1 9
9 3 13 11 7 11 13 13 9 9
12 11 3 15 3 11 13 9 0 13 1 15 13
18 6 0 15 9 7 15 9 9 9 9 15 9 3 13 13 9 9 0
16 7 3 6 9 9 1 15 7 13 0 3 13 9 3 1 9
8 7 3 13 1 15 9 7 9
7 7 13 13 15 15 9 13
10 3 9 16 13 13 13 13 1 9 9
13 7 16 1 11 13 11 7 15 1 15 13 11 11
6 7 13 9 9 9 13
12 1 9 3 9 7 9 13 9 9 1 15 13
12 9 9 16 15 13 1 15 9 9 1 9 13
8 13 3 11 7 9 9 13 13
7 9 9 7 15 13 9 13
33 9 9 11 13 9 15 7 9 13 16 13 9 1 9 11 7 1 9 13 13 15 1 15 7 1 12 9 9 9 15 13 1 9
18 7 13 9 12 1 9 11 9 13 15 9 15 3 1 12 7 12 9
9 7 1 0 13 9 3 1 11 9
13 7 13 0 9 11 9 11 9 1 9 11 9 12
7 7 13 0 13 0 11 9
5 15 3 9 13 13
13 13 11 9 11 9 1 9 15 15 13 15 9 15
21 0 9 1 9 1 9 13 11 9 11 13 11 1 9 9 15 9 9 15 9 11
7 16 13 3 11 9 15 13
7 15 15 13 13 3 13 15
12 7 6 13 1 15 15 3 13 0 9 9 13
15 16 13 15 15 1 15 13 13 13 15 1 9 13 1 9
6 9 3 13 15 1 0
16 15 13 13 1 9 0 0 15 3 13 1 15 1 11 1 11
8 15 3 3 13 9 15 1 9
20 7 15 15 13 0 15 1 9 15 9 13 13 16 0 9 13 9 15 13 11
7 3 3 1 9 0 13 13
4 9 15 13 15
15 16 3 13 15 1 0 3 3 3 13 1 9 3 13 16
5 3 7 3 3 13
6 3 13 0 15 13 9
9 11 3 15 9 16 13 9 9 13
9 7 13 13 1 9 15 7 13 9
7 15 3 9 13 3 13 9
13 0 3 13 15 9 9 16 1 0 15 9 9 13
9 13 3 16 13 15 13 13 1 9
21 13 9 7 13 7 13 16 9 13 15 1 9 15 9 15 3 13 16 15 13 15
14 16 13 13 9 13 13 0 9 7 13 9 11 7 11
9 15 13 13 15 16 13 1 9 9
10 0 3 9 3 0 9 13 13 9 9
15 13 3 9 9 13 13 9 7 13 0 15 1 11 13 13
6 3 3 11 7 11 13
14 7 16 13 0 7 0 15 13 0 9 6 13 1 9
5 3 3 13 15 9
13 13 15 1 9 9 16 13 1 9 3 1 9 9
8 7 13 3 13 13 1 9 0
7 13 3 9 9 1 0 9
17 9 3 13 0 9 7 0 7 0 9 7 13 9 1 11 7 11
6 7 13 15 1 9 15
7 9 3 13 9 7 9 0
19 13 13 3 11 16 3 13 9 9 7 13 3 16 13 9 7 9 0 9
14 15 3 0 13 9 13 7 1 9 13 9 9 1 9
22 0 3 9 13 13 3 13 1 9 9 13 9 9 15 13 9 7 9 13 1 9 15
6 7 15 3 13 1 9
4 15 3 1 9
34 16 3 13 13 9 9 7 9 1 9 15 16 9 13 7 13 15 13 13 1 9 11 11 7 11 7 0 1 9 9 7 3 13 13
4 0 13 11 13
14 15 13 15 7 13 16 13 9 16 0 13 13 0 9
5 13 1 9 15 0
4 7 13 7 13
12 9 3 16 13 15 13 11 13 9 15 3 13
4 7 13 11 11
3 11 3 11
17 9 3 11 15 13 1 9 9 7 9 1 9 13 1 9 13 13
16 15 3 13 9 11 7 11 13 9 15 13 1 9 13 7 13
4 9 15 0 13
29 3 15 0 13 0 15 9 13 15 1 0 0 13 1 9 0 15 13 9 7 9 7 9 7 15 15 1 15 13
11 15 1 0 9 13 15 9 13 1 9 15
23 7 3 3 1 9 15 3 0 13 13 1 9 13 9 7 9 0 13 9 7 9 9 15
8 13 3 15 1 11 7 11 9
16 13 3 15 9 13 13 9 7 0 9 13 13 1 11 1 11
24 16 13 9 0 7 13 0 13 13 11 7 11 7 11 13 9 9 13 16 13 1 9 7 16
9 1 0 9 13 15 13 1 9 9
18 7 16 13 0 1 0 9 9 7 13 1 9 13 15 9 1 15 13
14 13 7 11 13 11 7 13 1 11 9 9 13 1 11
13 7 3 13 11 3 13 13 9 9 1 9 15 13
17 16 3 13 7 13 9 13 15 13 9 1 0 16 13 9 9 9
9 16 13 1 9 11 3 13 0 13
30 13 3 9 3 0 11 7 11 1 0 13 16 13 11 7 11 7 15 15 1 0 1 9 7 9 1 11 1 0 9
12 0 3 13 1 9 13 11 7 11 13 9 9
6 7 13 9 0 15 9
19 16 3 13 11 13 13 1 9 7 1 9 7 0 13 15 9 13 1 0
10 13 3 15 1 9 9 15 13 13 16
8 13 13 15 13 3 13 9 11
9 13 7 9 7 0 13 1 9 0
21 9 9 15 13 16 1 0 9 1 15 13 9 1 9 15 13 9 9 9 7 13
25 7 15 13 9 9 9 13 13 0 9 0 3 3 15 7 15 13 1 15 7 0 9 13 9 15
20 3 3 15 13 9 13 9 1 9 9 15 3 7 9 15 3 7 15 13 13
10 7 1 9 9 11 13 13 3 3 0
4 13 3 15 9
16 7 13 11 7 11 13 15 13 9 9 7 9 1 9 1 15
6 7 16 13 13 11 13
4 9 9 13 15
3 3 13 13
30 1 0 13 7 13 9 11 15 13 7 13 15 13 7 13 0 16 13 0 9 9 7 15 9 1 15 13 13 9 15
4 13 9 13 0
7 0 1 9 13 9 9 15
29 1 15 15 13 3 13 15 15 1 9 13 1 9 7 13 1 15 16 13 15 1 9 9 7 9 7 13 7 9
19 11 3 1 9 0 13 1 0 9 15 15 13 1 9 3 1 15 9 13
29 3 13 9 7 0 1 15 9 13 9 1 15 7 13 11 1 11 7 11 11 15 13 11 7 11 9 0 1 9
16 9 7 0 9 0 15 13 11 7 11 7 11 9 1 9 9
12 13 3 11 7 11 15 3 0 15 9 13 0
26 13 13 3 9 0 7 15 15 3 13 15 9 3 0 3 16 13 15 1 13 9 7 9 13 7 9
6 1 15 13 15 3 13
1 13
5 0 3 13 13 11
5 7 13 9 13 9
16 11 3 7 11 3 0 16 13 9 9 0 13 13 9 7 13
15 13 3 3 9 13 13 1 9 1 9 1 15 15 13 0
8 1 15 3 9 13 1 11 11
14 13 13 9 1 0 9 1 15 13 9 9 3 15 13
11 11 3 13 15 1 13 3 11 15 13 11
21 11 3 13 15 15 13 1 15 1 9 7 3 13 1 15 1 9 3 13 13 15
15 13 13 3 9 3 16 13 1 3 7 11 13 11 13 11
7 13 3 11 7 11 13 9
6 13 3 1 11 7 11
14 7 6 9 15 13 3 9 11 9 9 11 0 9 0
6 0 13 11 15 1 13
11 7 13 13 15 1 9 15 13 1 0 9
8 13 3 15 16 9 15 9 13
18 16 3 13 9 13 15 13 9 15 13 13 1 9 7 0 15 13 11
15 13 3 11 7 11 9 13 13 1 0 9 13 9 1 11
8 16 13 3 1 11 13 13 11
6 7 3 13 15 9 11
6 16 3 13 11 13 11
10 9 9 15 13 13 7 13 15 7 13
5 13 1 11 13 15
17 3 3 9 13 3 13 13 1 11 0 13 16 13 15 9 13 15
10 7 3 11 15 13 0 9 11 9 9
8 13 3 1 0 9 9 15 13
13 9 3 9 13 13 1 9 1 9 3 13 9 13
6 7 13 13 9 15 13
11 7 15 9 9 11 9 9 9 13 9 13
10 16 3 13 13 7 9 15 13 13 13
12 16 13 15 0 9 13 13 1 9 15 7 13
21 13 13 3 13 15 1 9 9 15 13 9 9 13 15 15 9 0 13 9 15 13
7 0 13 11 7 15 13 13
11 0 9 9 9 0 13 15 13 15 9 9
5 0 3 13 0 9
7 13 3 11 7 13 9 13
9 13 15 1 9 11 11 13 1 15
18 13 3 9 15 16 13 9 9 15 13 11 7 11 13 1 9 1 9
8 0 9 13 9 15 16 13 9
14 7 13 9 15 3 13 15 13 3 7 13 16 13 9
5 7 13 9 1 15
8 7 9 13 9 15 13 9 13
16 7 16 0 9 15 13 13 15 1 9 13 9 16 3 13 15
16 15 16 0 9 13 13 15 1 0 9 7 9 15 13 1 9
9 0 3 9 11 7 11 13 13 9
6 7 13 13 3 9 15
5 7 0 9 13 13
17 13 3 9 9 7 13 13 9 9 13 9 13 15 13 13 13 13
6 13 3 11 0 9 13
4 15 13 15 0
4 0 3 3 13
5 13 7 9 13 13
6 7 13 13 11 7 11
8 9 15 15 13 13 16 0 13
3 3 0 13
11 13 1 9 11 7 0 13 15 7 9 15
13 7 13 13 15 9 9 1 15 15 13 1 9 15
10 7 13 15 1 0 9 9 13 9 15
8 7 13 13 15 7 15 15 3
18 16 13 15 1 9 15 13 15 9 7 13 13 1 15 9 15 13 9
9 7 16 9 13 13 13 9 9 13
4 13 9 16 13
6 3 3 13 13 1 9
4 11 3 13 15
9 13 15 3 0 9 0 13 1 9
5 7 3 3 15 13
2 3 3
6 7 13 7 0 15 13
6 13 7 13 16 9 13
7 13 3 1 9 13 1 11
9 7 13 9 13 13 15 7 13 13
12 16 3 13 11 7 11 13 11 3 13 9 9
28 1 9 3 11 13 1 15 7 1 9 12 13 15 1 9 13 7 13 16 11 13 13 7 13 1 0 7 16
8 0 13 11 11 15 15 13 15
23 7 15 1 15 13 7 13 13 11 7 11 7 1 13 9 7 9 0 7 9 0 3 0
9 7 13 9 11 13 15 13 1 9
15 7 16 3 13 15 13 11 7 15 9 1 9 9 13 16
12 7 0 15 1 9 11 13 9 15 13 13 11
8 13 3 9 7 9 9 13 0
10 7 13 3 1 11 7 1 0 13 15
11 9 3 3 1 9 13 11 7 11 1 11
7 15 16 13 1 9 9 13
14 7 0 3 13 1 15 7 0 9 0 7 9 3 0
22 16 3 13 1 11 9 16 3 11 13 13 1 11 9 9 13 7 3 13 7 13 9
11 3 7 3 11 13 9 16 13 3 1 9
24 15 3 13 11 13 3 11 7 13 9 1 15 1 11 7 11 16 3 3 13 1 0 13 13
15 11 3 16 11 15 13 13 9 15 1 15 13 9 13 9
18 13 3 1 9 1 9 7 13 7 1 9 1 15 9 1 15 15 13
12 15 3 0 7 0 9 13 1 15 7 15 13
2 15 3
5 0 9 13 9 13
6 16 11 7 9 13 15
7 7 13 15 1 11 13 13
6 0 3 15 13 9 15
7 13 3 13 15 13 0 13
17 0 3 15 7 9 9 1 15 15 13 3 7 13 7 13 15 0
8 9 0 1 15 3 0 15 13
13 13 3 7 13 9 15 13 3 9 1 15 13 13
2 0 9
8 15 3 13 13 0 15 13 15
38 9 15 13 9 7 15 15 1 15 13 0 9 7 9 16 13 9 3 1 0 9 13 3 7 9 0 13 13 15 16 15 13 15 9 7 9 7 15
8 1 15 3 13 7 13 7 13
6 3 3 15 15 9 13
21 9 3 16 13 9 3 13 13 9 7 9 7 9 9 9 7 9 9 9 13 0
38 7 9 3 0 9 13 9 3 13 9 16 15 3 9 13 3 16 13 9 1 15 13 13 9 1 9 1 9 1 15 13 9 13 15 13 15 1 0
8 16 13 3 9 0 15 3 13
3 15 3 13
5 13 15 1 0 3
6 3 11 13 1 0 15
13 1 15 7 11 11 7 9 9 11 7 15 1 15
29 7 13 15 9 9 11 0 9 15 3 13 1 11 7 11 9 15 3 16 13 11 13 15 9 1 11 13 1 15
10 7 16 0 13 9 13 1 15 7 13
4 13 3 0 9
16 16 13 3 1 11 11 7 11 13 9 11 13 9 13 11 11
10 13 3 15 7 13 13 9 13 1 15
5 9 15 1 9 15
2 0 15
9 11 3 9 13 9 1 15 9 15
7 7 0 9 13 13 7 13
7 13 3 9 9 1 9 11
28 13 13 7 13 7 3 13 1 16 15 13 15 1 7 15 13 15 16 13 15 16 9 13 15 0 1 0 9
11 13 3 9 7 12 9 13 1 15 9 9
17 11 3 9 11 13 12 9 9 1 11 7 13 15 1 9 13 16
7 1 9 0 13 9 13 9
9 13 3 11 13 9 13 11 1 9
14 16 3 9 13 1 9 7 9 7 9 15 15 0 13
5 9 15 0 13 13
5 7 13 15 1 9
9 13 3 15 11 9 9 13 1 9
6 7 15 15 11 9 13
23 11 3 16 3 13 9 0 9 13 13 11 7 1 15 11 7 11 15 15 13 1 11 9
3 13 3 9
7 13 7 11 7 0 3 13
10 7 13 11 13 7 13 9 7 13 11
17 7 13 3 0 9 13 13 13 1 9 0 9 7 11 13 15 9
14 9 3 15 11 9 0 9 9 0 13 11 0 1 9
5 0 13 13 9 9
15 7 13 9 13 7 13 3 15 15 13 11 13 3 9 11
7 0 3 13 3 13 1 9
14 15 16 13 11 7 11 13 15 7 3 13 15 9 9
8 15 16 13 13 0 0 15 13
18 13 13 3 16 11 13 11 16 11 13 0 9 13 11 7 13 15 9
4 13 7 1 15
5 3 9 0 13 13
4 3 0 1 15
7 7 3 16 9 0 13 13
3 0 3 13
2 15 13
3 1 11 9
19 11 13 9 9 9 13 1 15 15 13 13 1 15 16 13 0 13 1 11
8 0 13 13 13 1 9 9 11
16 7 16 13 0 9 11 13 9 0 1 15 7 13 9 7 13
6 13 3 15 9 3 12
15 13 3 9 1 9 13 1 12 9 13 7 13 1 9 9
19 0 3 13 13 1 9 3 16 15 15 13 1 11 13 9 9 9 7 9
30 9 7 3 15 9 13 1 9 11 3 16 3 1 0 13 1 9 15 9 7 9 7 13 1 15 9 7 9 0 13
19 13 3 15 3 1 13 0 9 13 1 15 15 13 9 0 9 9 11 13
12 13 3 15 11 0 9 9 12 9 15 0 13
6 13 3 9 0 13 15
5 11 13 7 11 13
4 15 3 15 13
12 0 3 0 13 13 15 9 7 9 15 13 11
11 7 13 9 1 15 0 7 13 9 9 11
9 0 7 13 13 13 7 13 9 15
14 0 3 1 0 15 13 0 13 13 9 7 13 1 15
7 3 3 9 9 13 7 13
15 0 3 13 13 11 1 9 13 11 7 11 13 11 13 16
8 16 13 3 13 15 3 11 13
11 13 13 3 1 0 9 9 3 0 1 9
14 11 3 15 9 9 13 9 0 11 13 9 3 0 9
10 15 13 7 15 15 0 9 13 9 13
9 9 13 16 1 0 9 9 13 15
26 7 13 7 13 16 3 3 11 7 3 0 11 11 0 13 13 0 9 13 16 3 13 9 15 9 13
8 0 13 13 13 9 7 13 13
3 0 11 0
9 11 3 13 13 1 9 3 13 9
19 15 3 3 1 11 9 15 13 9 15 13 1 15 13 16 15 13 1 9
4 15 3 15 13
4 13 3 9 13
7 7 0 13 15 1 9 13
8 1 9 3 13 11 13 15 9
15 15 3 13 9 13 9 13 13 12 15 3 1 9 12 13
6 7 16 13 9 9 13
17 9 0 15 3 13 9 15 13 0 9 9 13 0 11 11 7 9
14 16 3 0 13 3 13 13 15 13 13 7 15 3 13
12 13 3 9 0 3 7 0 3 7 13 9 15
20 3 16 11 7 15 1 15 13 9 13 1 15 9 9 0 13 7 1 9 13
2 13 3
11 16 15 3 0 9 13 1 0 9 13 13
18 16 3 13 9 13 11 9 7 13 15 13 7 13 13 16 13 1 11
14 16 3 13 9 0 7 13 15 13 0 9 13 1 11
14 3 16 13 9 12 13 13 0 9 1 9 13 1 11
7 13 7 9 16 13 1 11
22 13 13 3 15 11 11 0 9 3 11 7 11 7 11 0 7 11 9 3 11 7 11
6 0 16 13 13 15 11
21 15 3 13 1 9 9 1 11 7 13 1 15 11 1 9 12 3 13 13 9 12
22 1 12 3 9 16 13 1 13 9 11 13 15 13 1 0 13 7 9 3 1 0 9
26 13 3 15 9 9 11 1 9 16 13 9 0 13 3 11 13 9 13 1 0 9 3 7 13 13 0
8 1 15 16 13 11 13 1 15
3 7 13 13
2 13 13
6 9 3 15 1 15 13
16 13 3 13 7 9 7 13 3 7 13 3 1 9 3 13 13
9 13 3 9 13 7 13 13 3 3
10 15 3 13 9 13 1 11 3 13 11
16 7 3 13 0 9 13 1 11 7 15 13 11 7 0 13 11
12 13 3 11 13 11 16 15 9 0 13 1 11
11 13 3 16 0 15 13 16 9 9 13 11
9 1 11 3 13 11 13 0 3 9
10 15 16 13 1 15 7 3 13 13 15
32 15 13 1 0 9 15 13 13 1 11 3 15 1 1 15 9 13 13 9 1 15 9 7 9 7 9 15 15 13 1 9 9
28 3 15 13 0 16 13 15 7 13 15 3 7 1 9 13 9 7 9 1 9 9 7 9 1 9 15 11 11
4 7 15 0 13
19 7 3 6 15 13 16 3 3 13 9 15 15 15 1 15 13 13 9 9
11 3 13 15 0 9 16 0 13 1 9 15
9 3 3 13 16 13 15 9 9 15
19 13 15 7 0 9 1 15 15 9 0 13 9 13 9 9 15 13 9 15
14 15 13 16 13 1 9 15 9 0 1 15 3 13 9
13 7 1 15 0 13 9 13 0 16 13 9 1 15
19 7 3 13 15 9 7 9 9 15 15 0 13 13 7 13 9 1 13 15
7 9 7 9 7 9 15 13
17 15 13 15 16 3 13 13 13 0 7 13 9 9 11 16 15 13
6 0 13 3 13 3 13
11 7 16 0 13 13 9 15 1 15 0 13
6 0 3 9 13 13 15
20 7 13 1 9 11 13 15 13 3 1 9 15 13 16 3 9 15 3 13 13
20 16 3 13 13 16 13 13 1 15 0 9 13 11 7 0 9 11 7 3 11
9 7 16 13 9 13 1 11 13 13
15 16 13 3 11 7 13 15 1 9 13 1 11 7 13 11
7 13 3 9 13 3 9 12
8 15 11 13 1 9 16 13 11
15 7 13 9 13 13 13 15 15 1 9 7 9 3 1 9
6 7 13 9 1 9 13
5 0 3 13 1 15
8 15 3 9 13 1 11 13 11
8 7 13 9 13 9 12 1 0
6 15 3 9 13 13 11
7 0 3 13 9 12 9 13
13 7 16 13 1 9 15 13 15 1 11 9 9 11
8 15 16 13 1 15 13 9 11
4 0 13 9 0
15 9 15 13 9 0 3 13 1 11 9 7 13 1 9 9
13 15 16 13 13 15 7 15 9 0 13 16 13 11
5 3 13 11 7 13
7 15 13 13 7 13 9 15
8 7 16 15 13 3 13 13 13
3 9 9 13
18 13 3 3 1 9 1 11 15 1 13 1 15 13 11 15 0 0 9
8 7 16 13 11 3 13 15 9
14 0 3 9 13 11 15 1 1 11 15 7 13 13 0
14 15 16 13 13 1 0 15 13 9 1 9 1 9 15
9 3 0 16 13 13 9 13 7 15
9 13 9 3 12 13 1 9 15 13
27 13 3 1 15 16 9 13 1 11 15 15 1 9 13 9 13 3 13 13 15 9 15 3 7 1 9 13
4 3 13 13 9
4 13 3 15 13
6 0 3 13 15 15 13
8 13 15 9 12 9 13 1 15
13 0 13 13 15 16 0 7 13 1 0 16 13 9
16 7 13 15 16 15 1 15 13 13 13 7 13 3 15 13 9
22 3 11 13 9 0 9 13 1 0 13 1 9 13 9 9 9 16 13 1 15 15 9
15 13 3 11 0 1 9 1 15 15 13 16 1 9 13 11
10 13 7 13 9 0 7 13 13 9 9
7 7 13 11 13 15 1 9
5 7 3 13 13 9
12 13 3 15 13 13 13 9 9 16 0 13 11
9 15 3 13 9 7 9 13 1 0
9 15 16 13 9 7 9 13 13 11
10 3 13 9 13 15 7 13 13 9 12
6 15 3 15 13 1 9
13 7 16 3 13 0 13 1 9 13 13 15 1 9
13 7 16 13 1 9 13 16 13 1 9 1 9 9
5 13 3 9 9 13
2 13 15
9 7 16 13 13 1 9 11 13 9
7 3 13 15 13 15 1 15
2 15 13
12 15 9 13 3 0 1 11 11 3 0 9 9
3 13 3 15
5 13 15 13 1 9
21 7 16 0 13 11 13 1 9 13 9 1 9 7 0 9 13 13 13 0 9 13
11 9 9 7 9 13 15 1 15 3 13 9
12 16 13 3 16 0 9 13 1 0 3 13 9
2 7 13
26 15 0 9 13 13 3 1 9 13 7 13 1 9 9 7 9 3 9 9 9 15 13 7 15 0 3
17 13 13 3 13 15 7 13 11 0 9 3 1 9 13 15 9 0
8 7 13 1 9 13 9 13 15
5 11 11 15 15 13
3 15 3 13
3 15 13 9
4 13 7 1 15
8 7 15 15 1 13 9 3 13
9 9 3 3 13 15 15 13 15 1
3 15 13 9
5 9 3 13 1 15
3 13 13 11
10 7 3 15 13 1 15 15 15 13 13
15 7 16 3 13 1 9 9 0 1 9 13 1 9 13 11
3 11 9 13
7 7 15 0 9 13 1 15
3 3 0 13
4 7 3 15 13
1 13
8 13 7 13 9 15 13 9 15
21 13 13 3 13 15 1 11 7 13 1 9 13 15 1 9 9 7 13 0 13 15
18 9 15 13 16 15 13 13 1 9 7 13 1 9 15 15 13 1 15
16 7 16 13 9 11 9 15 15 13 7 13 7 13 9 13 0
4 7 13 1 15
8 13 16 15 1 9 3 13 15
5 13 1 9 0 9
6 3 3 9 13 15 13
32 13 3 15 7 13 9 15 7 9 13 1 9 13 9 13 15 1 9 7 9 13 7 13 15 16 13 1 15 9 3 13 15
8 3 9 0 7 0 13 15 13
9 15 13 9 13 1 9 7 13 13
3 15 13 13
6 0 3 9 9 0 13
5 13 3 9 13 0
3 15 9 13
3 3 0 13
3 7 13 9
7 15 0 9 9 0 13 13
3 7 11 13
5 15 3 3 13 13
9 3 3 13 1 0 15 15 13 13
13 9 3 13 16 13 16 9 0 13 7 16 13 15
6 7 13 11 13 1 0
14 9 9 15 15 9 0 13 13 1 9 3 1 0 9
10 9 3 9 11 13 13 15 13 9 15
5 3 11 1 15 13
5 13 15 9 9 0
13 7 15 13 13 15 1 9 7 1 9 13 15 13
4 7 15 13 13
4 0 9 9 13
3 13 13 3
5 9 9 15 3 13
14 13 3 11 16 12 9 13 9 7 0 9 13 1 9
5 9 9 15 9 13
2 9 9
7 1 9 7 9 0 15 13
15 7 16 0 13 13 13 9 1 9 7 9 7 13 13 9
12 9 3 13 3 13 9 3 7 9 3 7 9
5 13 13 3 9 0
6 7 13 15 9 13 13
6 15 0 13 1 9 0
4 15 3 3 13
7 9 3 13 3 15 3 13
17 13 3 15 1 0 9 9 13 16 13 13 11 7 3 13 1 0
16 7 3 1 9 15 1 9 15 9 13 13 1 9 13 9 0
32 1 15 16 13 11 1 9 7 9 9 9 9 0 1 9 13 9 1 9 1 9 9 13 15 9 7 15 15 15 1 3 13
7 7 3 3 13 13 9 12
24 9 3 15 13 9 15 13 1 9 15 1 9 9 15 16 1 9 9 15 13 3 1 9 15
13 7 13 7 13 9 3 3 9 15 13 0 1 9
21 16 3 9 15 9 3 13 3 15 9 13 13 0 9 9 3 13 0 15 13 9
5 15 3 3 13 9
4 15 3 9 9
4 15 9 0 13
2 13 15
7 15 9 9 7 9 0 13
4 3 9 9 3
10 0 15 13 13 9 7 15 13 13 9
6 3 3 1 0 15 13
8 3 1 0 3 15 3 13 13
3 0 15 9
7 9 3 15 13 3 13 9
6 3 15 13 15 15 13
3 15 3 13
5 9 3 15 15 13
8 6 9 15 15 13 15 13 9
7 3 3 13 9 9 7 9
4 3 3 15 13
5 15 3 13 9 9
5 7 15 9 15 13
7 7 16 13 9 15 13 0
5 16 7 13 9 13
9 16 7 3 13 16 7 13 9 13
5 3 3 13 0 15
8 3 15 3 13 0 7 15 0
21 13 3 15 9 16 13 15 15 9 7 9 1 9 15 15 13 13 7 13 1 0
11 0 9 3 11 9 15 3 13 7 15 9
37 11 13 9 11 11 1 9 9 7 11 9 9 9 15 13 11 13 1 11 11 13 0 1 15 15 13 9 9 15 11 11 1 15 9 15 7 15
7 13 9 0 7 9 0 13
23 7 13 9 9 1 9 15 0 13 15 13 9 1 9 1 9 15 15 15 9 0 9 13
8 16 15 9 13 15 13 9 13
5 13 0 1 9 15
11 15 3 15 0 13 7 3 1 0 13 13
9 15 7 13 0 9 7 13 9 9
4 15 3 15 13
6 15 3 13 15 3 13
12 3 16 12 12 9 13 1 11 7 3 0 9
46 15 3 0 9 0 3 9 3 13 3 0 15 15 3 13 13 1 9 9 15 11 11 13 15 7 15 9 1 9 9 11 13 0 9 11 1 9 9 16 9 0 13 1 9 9 11
31 3 3 13 15 3 13 16 15 15 9 13 13 9 7 0 7 9 13 7 0 7 0 7 0 1 0 9 3 7 9 13
6 13 3 3 13 7 9
15 16 15 9 9 13 0 7 0 13 13 1 0 3 13 0
11 3 13 3 9 13 9 7 9 1 0 9
4 3 13 15 9
6 9 3 9 13 0 9
26 3 15 13 1 9 15 0 3 13 9 9 3 13 15 9 7 0 13 1 9 15 13 9 15 3 13
32 3 3 16 13 15 13 9 7 1 9 7 1 9 16 13 9 0 7 9 0 15 3 12 9 9 1 15 15 7 15 1 0
7 0 3 15 1 9 13 0
7 3 15 13 9 9 13 9
16 16 7 3 13 16 7 13 7 15 15 13 15 1 9 9 13
7 9 15 13 3 3 15 11
10 3 3 9 1 9 3 3 9 1 9
4 15 3 1 9
12 0 3 15 13 12 7 0 9 13 0 3 13
22 7 15 3 13 9 1 9 3 9 3 9 3 9 3 9 3 9 9 9 9 9 9
4 16 7 9 13
4 16 7 9 13
4 16 7 9 13
8 3 13 13 9 13 15 13 0
22 3 15 1 9 13 9 13 7 9 7 9 16 9 9 13 3 13 15 13 7 15 13
5 0 9 15 0 13
6 7 9 9 9 0 13
9 3 16 0 3 13 3 7 11 13
5 0 11 1 9 13
5 15 0 0 3 0
6 7 15 0 0 3 0
12 16 3 15 13 13 0 9 7 15 13 7 13
6 13 3 15 0 9 13
12 9 15 7 9 1 9 9 15 7 9 11 11
25 16 7 3 13 1 15 9 7 9 16 7 13 1 15 9 15 13 1 9 15 9 15 3 15 13
27 3 3 13 13 15 9 1 9 15 15 13 13 1 11 16 1 9 13 13 1 9 3 16 13 15 3 13
20 7 0 1 15 0 9 9 13 16 3 13 13 1 15 7 1 9 15 13 0
8 15 1 0 9 13 15 7 13
14 1 15 13 16 3 3 13 13 3 15 1 9 1 15
16 16 1 0 9 15 15 1 15 13 9 1 0 9 13 1 15
5 3 9 15 0 13
10 3 3 15 13 15 3 15 13 7 13
31 7 0 9 13 3 13 1 15 16 0 9 13 7 1 15 13 1 11 7 3 1 11 13 1 15 7 1 15 13 1 11
13 7 15 13 1 9 13 16 13 1 15 13 7 3
17 0 3 9 16 9 15 15 13 1 15 3 13 1 0 13 7 3
28 9 3 9 11 11 15 1 15 1 15 13 13 1 15 7 11 7 11 3 13 13 7 3 7 13 1 0 13
8 3 3 9 9 13 1 0 13
9 3 7 1 15 6 9 1 9 15
13 15 3 13 15 15 1 1 11 7 15 13 15 9
15 15 3 9 9 13 1 9 15 16 13 15 3 13 1 11
10 3 16 13 9 15 7 9 13 9 15
17 3 16 1 3 3 13 7 13 16 3 0 9 13 15 0 9 13
11 3 3 13 3 0 13 9 9 7 1 9
9 7 3 1 9 1 9 1 11 13
9 7 3 13 7 0 7 0 13 0
19 15 3 15 13 13 1 9 11 16 13 15 0 9 3 13 7 0 7 0
5 16 7 0 13 15
10 9 0 13 15 7 1 9 9 13 15
10 15 3 13 9 9 0 3 13 9 16
7 1 15 1 15 13 1 9
18 0 13 15 0 9 13 16 15 13 9 1 9 0 0 3 0 1 9
11 3 0 9 9 9 0 13 15 1 9 11
24 13 9 1 11 1 9 12 7 1 9 13 7 1 9 13 9 13 13 0 9 3 1 0 9
4 1 0 9 13
8 6 0 0 0 13 13 1 15
10 13 3 3 15 0 13 15 3 0 13
21 3 0 0 13 16 3 0 3 13 1 9 15 9 13 15 1 9 7 3 1 9
9 3 3 13 9 3 3 13 1 9
2 13 3
3 15 15 13
6 15 15 13 9 3 13
6 1 0 9 3 13 9
19 9 7 16 13 13 9 1 15 9 15 15 0 13 0 9 13 1 9 9
5 13 3 13 9 15
43 9 13 9 3 3 11 13 9 7 15 0 13 1 15 16 0 13 13 9 9 1 9 16 13 15 15 0 9 3 13 9 7 9 7 15 0 9 7 16 13 0 7 0
18 11 7 11 9 11 11 15 0 1 11 11 15 13 11 1 9 7 9
12 9 15 7 9 1 9 9 15 7 9 11 11
19 7 1 15 9 3 3 3 3 13 11 1 9 15 7 1 9 7 1 9
35 13 3 0 1 15 9 1 9 7 0 9 1 9 13 16 1 9 11 3 1 9 13 13 9 15 16 13 15 15 1 15 13 1 15 9
2 13 9
3 13 0 9
2 13 9
2 9 3
4 15 13 9 0
8 0 3 13 16 1 0 13 13
9 13 3 15 9 13 15 1 9 11
12 7 3 15 0 13 13 7 1 3 7 1 15
74 9 13 13 9 3 1 15 9 3 3 0 13 16 13 9 15 7 13 9 15 15 15 1 3 3 16 3 15 0 1 15 13 1 9 9 1 9 15 7 9 1 15 9 15 7 9 15 13 1 9 0 9 9 16 0 13 9 9 1 15 3 13 16 3 0 13 1 9 13 9 0 15 15 13
12 7 13 9 15 13 7 1 9 7 1 9 15
20 0 3 15 0 9 13 13 7 13 1 9 11 11 16 1 9 13 15 9 13
18 3 16 15 3 13 9 15 1 9 0 13 7 3 13 1 0 16 13
14 9 3 1 15 0 13 9 13 9 15 3 13 7 0
7 3 0 16 3 13 15 13
9 13 3 9 7 15 13 0 0 13
7 7 15 11 13 3 15 13
22 7 0 9 9 13 13 9 0 13 9 15 13 15 7 13 1 9 15 15 13 9 9
10 0 3 13 16 1 0 9 13 9 0
7 9 3 9 0 9 9 0
21 0 9 1 12 7 0 9 13 13 16 13 13 15 0 9 13 7 13 0 9 13
11 3 13 15 9 9 15 9 9 1 9 15
10 3 3 9 13 9 9 0 1 15 13
7 3 3 3 13 15 0 15
8 3 3 15 13 13 3 3 0
17 7 1 15 13 3 3 1 9 3 3 1 15 3 0 13 1 9
10 15 3 15 9 13 9 0 13 9 9
13 13 3 15 13 0 15 3 0 13 1 9 11 9
10 3 3 1 9 9 13 3 13 15 11
9 9 3 1 0 13 11 11 7 11
5 15 0 3 13 9
6 9 0 7 9 13 13
13 15 3 0 9 13 13 3 1 12 13 13 15 9
14 15 13 9 15 16 9 15 13 15 13 9 3 3 13
7 6 15 9 3 0 9 13
6 3 9 9 13 9 9
6 3 3 13 1 0 15
4 15 3 3 9
4 3 3 9 9
5 3 9 0 15 9
11 1 15 7 0 15 1 9 13 9 13 13
5 3 9 0 13 0
17 13 3 3 9 1 9 3 3 1 15 13 9 0 15 13 9 9
15 16 13 16 3 13 9 13 15 7 9 15 3 13 1 15
12 15 13 15 13 15 7 9 15 3 13 9 13
6 13 15 9 16 13 0
6 13 15 9 16 13 9
9 13 15 9 16 13 15 15 1 9
15 13 15 9 16 0 13 7 9 9 1 15 13 7 13 0
12 15 13 9 3 15 15 13 16 11 3 13 11
10 7 0 9 3 13 9 16 9 9 13
8 15 3 13 3 13 0 1 9
6 3 1 0 13 16 13
5 3 7 6 15 13
9 15 3 13 0 6 13 9 0 0
10 15 3 13 13 0 9 16 9 13 9
4 0 13 13 15
4 13 9 1 9
15 9 11 11 15 13 0 9 3 13 9 15 15 13 13 3
20 7 13 13 1 9 15 9 15 11 15 9 13 9 9 7 9 11 11 15 13
16 0 15 13 7 15 13 9 9 7 13 15 15 1 15 13 13
7 11 12 9 15 13 1 11
15 9 15 7 9 1 15 15 13 7 15 13 7 15 13 13
10 7 1 12 9 15 1 9 9 15 13
13 6 13 1 9 7 13 15 15 9 7 15 15 13
8 7 13 15 1 15 15 9 9
1 3
1 6
8 15 13 9 7 9 9 7 9
15 13 1 9 1 0 9 7 13 1 15 9 0 3 9 13
5 15 13 13 1 9
10 7 13 13 16 13 9 15 13 15 1
6 7 13 13 12 9 0
16 7 1 0 12 9 0 9 9 13 9 7 13 1 9 9 9
18 9 3 15 7 9 13 0 3 9 0 3 9 7 9 15 3 9 9
7 7 13 1 9 15 9 12
9 7 1 9 15 9 15 9 0 13
10 7 16 13 15 13 1 9 15 3 0
2 13 13
17 15 13 0 7 0 7 0 7 13 0 7 6 13 13 1 9 9
6 7 13 9 9 7 9
13 13 3 15 13 7 15 13 7 15 13 13 1 0
6 12 9 9 13 12 9
6 7 9 12 12 9 13
4 9 11 9 13
10 7 13 15 15 15 13 9 7 3 13
4 7 13 15 9
11 7 9 13 7 13 1 9 15 7 3 13
9 7 13 1 15 16 9 15 0 13
5 0 13 3 3 13
7 7 13 9 7 0 9 13
11 7 0 13 16 13 9 9 15 7 15 13
8 15 13 9 13 15 9 13 9
5 7 9 11 9 13
10 0 13 0 7 0 15 13 0 7 13
9 13 9 15 7 9 15 7 0 13
16 7 13 1 0 15 15 13 9 13 7 3 13 7 13 9 11
6 15 0 13 15 13 13
10 6 13 13 9 1 15 1 9 16 13
5 7 13 9 9 12
10 13 0 3 1 9 7 13 15 9 9
5 7 9 11 9 13
8 0 13 15 13 9 15 9 0
7 13 3 13 3 9 13 11
9 7 13 9 15 7 3 13 9 15
6 7 13 1 15 0 16
16 13 3 13 9 11 15 13 11 13 9 1 9 11 13 7 13
7 3 13 7 15 13 9 9
13 16 3 13 15 3 7 13 1 0 1 9 9 15
10 13 13 15 9 0 7 13 0 9 0
12 7 1 9 9 0 13 15 15 13 3 15 13
5 7 9 11 9 13
10 0 13 9 9 15 13 9 3 9 9
5 7 9 15 0 9
18 13 9 15 7 9 7 9 7 9 7 9 15 7 9 15 0 0 0
17 13 9 11 15 15 13 9 13 7 13 9 15 13 7 13 1 9
7 7 13 0 9 16 9 13
5 6 13 15 1 9
14 7 15 13 1 15 1 9 0 16 9 13 1 9 15
17 7 9 15 13 1 9 7 13 15 9 16 15 13 13 9 7 9
7 7 13 15 15 1 9 15
7 15 3 13 0 15 11 13
7 3 15 15 13 13 16 13
22 7 15 13 7 15 13 3 1 9 9 15 13 0 9 1 9 7 13 0 1 9 0
4 3 9 9 13
5 7 13 0 9 0
8 15 13 9 13 15 9 13 9
5 7 9 9 11 13
10 0 13 15 13 12 9 9 7 12 9
8 13 13 7 13 0 15 13 13
9 3 3 13 9 15 0 1 9 15
13 1 9 3 13 3 13 7 13 7 13 7 9 13
14 16 3 3 13 13 3 9 7 13 15 9 13 1 15
9 7 13 15 1 1 0 16 0 13
25 15 13 3 13 9 0 7 3 13 9 15 1 9 9 7 13 9 15 1 9 15 7 1 9 15
8 15 13 9 13 15 9 13 9
9 0 13 0 7 0 15 13 9 11
5 15 13 7 15 13
5 7 13 7 15 13
3 13 9 15
15 6 13 1 9 11 15 13 15 9 13 7 3 13 7 13
28 7 13 16 15 13 15 16 13 9 9 15 7 15 15 13 1 9 9 15 13 13 1 9 0 13 13 1 9
2 13 3
14 15 13 13 0 9 1 9 9 15 7 3 3 13 3
25 7 13 1 15 9 9 15 7 9 9 9 15 0 11 15 13 1 9 1 9 15 7 9 15 0
8 15 13 9 13 15 9 13 9
5 7 9 11 9 13
2 0 13
4 13 9 15 16
5 3 0 13 7 0
7 0 13 7 13 7 15 13
14 7 13 16 15 13 0 7 0 7 0 7 0 7 0
28 13 15 13 1 15 9 13 13 16 0 13 7 9 0 13 7 3 13 9 9 15 7 9 13 9 15 16 13
6 15 15 13 13 7 13
5 13 3 7 9 13
6 6 13 1 9 7 13
19 16 15 13 9 15 7 13 9 13 1 0 7 13 1 0 7 15 15 1
8 15 13 9 13 15 9 13 9
3 1 0 13
17 7 6 9 13 1 9 7 9 0 15 13 3 9 13 15 1 13
10 13 3 7 13 15 15 13 13 1 0
4 3 13 1 9
11 7 6 9 13 13 1 9 7 1 9 13
10 7 15 13 0 13 9 9 9 7 0
9 7 9 13 1 9 9 0 9 0
15 7 1 0 9 7 1 9 9 12 0 0 9 3 7 3
23 7 9 0 0 9 7 0 9 0 9 7 0 9 13 9 3 9 7 0 9 0 9 13
8 7 12 9 0 15 13 9 0
8 7 1 9 7 3 0 13 9
8 7 9 3 13 9 7 9 13
15 0 0 0 9 9 0 15 13 7 15 13 7 15 13 13
37 7 16 13 10 0 9 7 9 7 9 13 1 9 13 1 9 9 13 12 0 1 13 1 9 7 13 13 1 9 9 7 13 9 15 1 9 13
15 7 13 1 9 13 1 9 9 13 3 7 3 13 9 12
19 7 15 13 1 9 3 7 1 9 3 7 1 9 13 9 3 7 13 0
15 7 15 13 0 16 15 0 13 13 13 9 3 7 13 15
6 7 12 1 0 13 15
2 3 13
14 6 13 9 1 9 11 9 11 13 9 7 12 9 15
24 7 16 13 9 12 0 7 12 0 13 1 9 13 0 9 7 9 0 0 9 15 13 9 0
5 7 13 0 9 13
4 7 13 1 9
20 0 13 9 15 13 13 13 9 7 9 7 9 7 9 7 9 7 9 7 9
15 13 1 9 7 9 9 7 9 7 9 7 9 1 9 9
4 7 12 9 13
1 6
3 7 0 13
2 7 13
1 13
2 7 13
9 7 16 13 9 0 13 0 9 13
1 13
5 7 13 15 9 0
24 7 15 13 1 0 13 13 15 16 13 9 1 9 7 16 3 15 13 7 13 13 0 9 0
9 7 16 13 9 0 13 0 9 13
10 7 15 13 1 15 13 9 1 9 15
9 7 13 3 9 1 0 12 0 13
14 0 9 9 7 12 0 9 9 7 9 7 9 3 13
3 13 7 13
4 7 6 9 0
28 7 15 13 3 9 0 9 7 9 13 15 7 13 13 0 9 1 12 9 9 13 9 9 7 9 7 9 9
18 7 16 13 0 9 13 1 9 9 13 1 9 9 7 1 9 15 13
17 3 9 0 7 0 3 13 7 13 9 15 1 0 15 13 1 9
7 7 13 13 0 0 9 0
22 7 13 13 0 16 13 9 3 0 16 13 9 15 7 9 15 15 13 13 3 7 0
6 7 13 16 13 9 0
7 7 9 0 13 13 3 9
15 7 9 9 13 1 9 3 9 13 9 15 16 9 0 13
6 7 9 13 3 9 13
23 7 9 9 7 9 7 9 7 0 7 0 7 15 9 7 9 13 15 1 9 7 9 9
5 7 13 9 7 9
4 7 15 13 13
28 1 0 13 12 9 13 1 12 9 9 13 12 9 9 16 13 9 1 9 3 7 1 9 3 7 1 15 9
12 7 13 0 9 13 1 9 9 13 9 9 0
17 13 13 9 3 7 9 3 7 9 16 13 9 9 15 1 9 15
12 7 13 9 13 12 12 13 1 15 9 9 11
5 1 9 11 12 12
5 1 9 11 12 12
5 1 9 11 12 12
5 1 9 11 12 12
5 1 9 11 12 12
5 1 9 11 12 12
5 1 9 11 12 12
5 1 9 11 12 12
6 1 9 11 12 12 13
5 7 13 9 0 13
9 9 9 15 15 13 1 9 7 9
12 7 15 9 13 1 9 9 7 0 7 12 0
12 7 13 1 9 9 1 9 15 7 13 9 13
1 6
7 7 13 12 1 0 13 15
8 0 15 13 13 9 0 15 13
3 7 3 13
3 7 13 0
4 9 15 15 13
3 7 13 15
17 0 13 15 13 1 9 0 7 13 9 15 7 13 15 1 9 9
14 3 13 1 9 9 7 13 15 9 7 9 1 9 15
13 7 16 13 9 0 13 13 9 1 9 3 0 9
8 7 13 12 9 13 1 9 9
6 7 13 13 0 12 9
11 7 15 9 13 7 13 1 9 13 9 0
18 7 13 13 0 9 0 16 13 9 9 15 1 9 0 15 13 1 9
12 7 13 9 9 1 9 9 1 9 9 1 9
14 7 13 9 9 7 13 0 1 9 9 7 13 1 9
10 7 13 13 9 7 9 7 9 7 9
5 7 0 9 9 13
31 7 3 9 0 9 13 13 13 1 9 7 13 13 0 9 9 9 7 13 13 0 9 9 15 13 9 7 0 9 9 13
5 7 0 9 9 13
19 7 13 1 9 9 0 13 3 9 7 13 1 0 9 9 7 1 9 9
24 7 9 9 13 11 7 13 13 0 9 9 1 9 7 0 9 13 13 1 9 16 0 13 13
5 7 0 9 9 13
28 7 13 13 0 9 9 7 0 9 9 7 0 9 9 16 13 0 9 15 7 9 3 13 9 0 7 9 3
16 6 6 6 13 1 9 1 0 9 9 12 9 15 13 9 13
15 7 13 9 1 9 13 1 9 7 13 13 0 9 9 9
4 7 13 9 9
8 7 13 9 9 3 9 9 0
9 7 13 13 9 7 9 1 9 9
17 7 1 9 13 9 1 9 7 13 13 0 9 3 13 9 9 9
11 7 1 9 0 13 9 9 7 3 13 15
8 7 9 9 0 9 13 1 9
6 7 9 15 3 9 9
18 7 13 9 3 9 0 7 9 9 15 3 9 9 9 0 13 1 9
10 7 13 9 0 9 7 9 1 9 15
6 9 15 13 9 9 12
3 6 12 13
7 6 13 3 12 6 1 0
19 7 13 9 12 1 9 9 0 15 13 1 9 9 13 0 9 15 13 9
10 13 12 9 15 13 13 1 9 0 11
21 7 13 13 12 9 15 13 13 1 9 7 9 7 9 7 9 16 13 0 9 9
3 13 9 15
6 7 3 13 9 1 9
19 7 15 13 1 15 13 9 0 7 0 7 0 7 9 9 13 3 9 9
10 7 1 9 15 13 9 7 9 7 9
11 9 3 9 1 9 15 13 7 1 9 15
7 3 9 0 0 9 13 9
4 7 1 0 13
66 7 0 9 15 3 13 13 1 0 9 3 7 9 13 1 9 9 15 16 3 13 9 7 9 0 7 0 7 0 7 0 7 0 15 3 7 13 13 3 7 13 3 7 13 7 3 13 9 1 9 15 3 7 1 9 15 3 7 1 9 15 3 7 1 9 15
7 7 13 1 9 15 9 13
11 7 13 9 15 0 1 9 0 3 1 9
8 7 13 9 0 3 16 9 13
8 7 16 13 13 12 9 13 13
6 7 13 9 1 9 13
6 13 15 13 13 12 9
4 7 13 15 13
15 7 9 15 13 13 1 9 7 1 9 13 9 15 1 9
20 7 1 9 9 0 9 16 13 9 13 7 13 9 9 3 13 1 9 15 9
12 7 9 15 13 1 9 3 13 15 1 7 13
12 13 9 0 1 9 9 13 1 9 7 1 9
10 7 13 1 9 13 15 16 13 15 9
3 7 13 15
4 13 7 13 0
13 7 13 13 9 15 7 1 9 15 13 0 3 9
9 7 13 9 1 9 9 7 13 15
3 7 13 15
8 7 13 13 15 9 0 9 13
11 13 7 13 9 9 7 9 7 13 1 15
12 9 3 15 13 3 9 13 3 7 3 13 15
11 7 13 12 9 15 7 13 9 12 13 9
12 0 13 12 9 7 12 9 1 9 9 9 13
15 7 16 15 15 13 13 9 13 1 9 0 7 13 9 15
10 7 16 15 13 15 13 3 13 15 13
20 7 16 13 9 15 9 15 13 1 9 13 1 0 9 7 13 15 7 13 0
19 7 9 15 1 9 9 0 15 13 3 11 7 11 3 7 9 15 13 13
17 7 13 1 9 7 9 7 9 7 9 9 15 1 12 9 7 9
8 7 9 15 3 13 13 1 9
8 7 13 9 13 1 0 7 13
14 7 9 13 3 16 0 12 9 13 15 15 13 1 9
13 7 1 9 12 7 9 9 9 1 9 13 1 15
14 7 13 1 9 15 7 9 0 13 1 15 15 13 15
2 13 3
6 7 13 1 9 1 9
5 7 13 0 9 15
13 7 1 0 9 13 13 9 0 7 0 9 9 13
9 7 13 13 1 9 9 9 12 12
11 7 0 1 9 13 13 7 13 9 9 9
3 6 0 13
5 6 6 0 13 3
15 13 13 9 0 9 9 15 7 11 15 7 13 1 9 9
19 7 12 0 15 1 9 9 13 1 9 15 13 1 9 15 7 13 9 13
33 7 13 13 9 7 13 9 15 7 9 0 13 7 13 9 9 15 9 7 0 7 13 9 15 0 7 0 7 13 15 15 13 9
7 7 13 13 9 9 1 9
20 7 13 13 9 9 15 1 9 15 7 13 13 9 7 9 7 9 7 9 0
6 7 9 0 13 1 9
15 9 13 9 7 9 1 9 15 7 1 9 15 9 9 12
7 7 13 13 15 9 1 9
19 7 1 9 15 12 9 7 9 15 13 0 9 9 9 7 13 15 1 9
14 7 9 13 1 9 15 13 13 16 16 13 9 15 13
12 7 13 9 0 15 13 13 15 9 1 9 0
28 7 13 13 9 15 1 9 7 1 9 15 7 9 13 1 9 3 13 9 13 1 9 16 3 13 0 9 12
6 7 13 13 9 1 9
13 11 7 9 15 13 1 9 7 9 13 7 9 15
17 7 13 13 9 0 0 9 0 15 13 9 7 11 15 13 0 9
11 13 13 1 9 7 9 15 1 0 13 13
20 7 15 13 0 1 9 9 7 1 9 9 15 7 3 13 9 15 3 1 9
8 3 13 9 7 15 13 1 15
17 6 9 7 9 16 13 9 1 15 13 9 0 13 16 0 9 13
15 7 16 13 9 16 13 13 1 9 13 13 9 15 13 0
27 7 13 13 9 12 9 9 0 16 13 1 9 1 9 15 3 13 1 9 7 9 7 9 9 1 9 9
18 7 13 9 9 7 13 9 9 15 7 13 9 15 13 9 1 9 15
6 7 13 13 9 1 9
17 7 13 13 9 1 0 1 9 15 15 13 9 9 7 13 9 11
24 7 13 1 9 9 13 13 9 12 7 9 12 7 1 9 15 12 9 7 1 9 15 9 9
18 7 9 15 13 0 13 9 7 9 15 3 9 7 9 15 3 9 9
9 7 13 0 9 9 15 7 9 0
9 7 12 1 9 15 3 13 1 9
7 7 13 13 0 9 1 9
7 7 13 9 16 13 9 9
4 7 13 9 13
3 15 0 9
9 7 13 13 15 9 13 0 7 9
8 7 13 13 0 9 13 9 12
20 7 13 9 15 1 9 1 9 13 9 15 7 9 15 7 15 15 1 9 13
21 7 13 13 15 9 1 15 9 7 9 7 9 7 9 7 13 15 15 15 13 9
5 16 15 13 9 13
6 15 1 9 1 9 13
8 15 1 9 13 13 15 9 13
6 0 13 9 7 9 0
9 7 9 0 9 15 13 1 9 15
15 7 13 9 7 13 1 15 13 9 0 15 13 13 9 9
28 7 13 13 9 1 9 15 13 13 0 13 1 9 9 13 13 1 9 16 13 9 9 15 13 9 9 7 13
14 7 13 13 0 16 13 9 9 9 16 7 13 9 9
8 7 13 15 3 13 9 9 13
23 7 13 15 0 7 0 7 0 7 0 7 0 7 9 13 9 1 0 9 7 1 9 15
3 0 9 13
6 15 13 9 13 9 9
5 7 9 15 13 12
23 7 6 9 13 1 9 11 7 1 0 12 12 13 9 15 7 9 9 15 13 1 9 15
14 7 13 9 1 9 3 9 9 0 7 3 9 9 0
10 7 9 15 13 3 9 13 1 9 15
13 7 13 3 9 0 1 9 7 1 12 9 7 0
14 7 15 13 13 9 3 0 12 12 15 13 13 1 9
8 0 13 15 1 9 3 13 13
3 9 3 13
8 7 1 9 15 3 13 13 9
3 1 9 13
26 7 13 0 9 13 1 0 9 13 9 0 16 13 13 1 9 7 1 15 9 7 9 7 9 7 9
11 13 9 7 13 0 9 16 13 9 9 15
13 7 13 15 15 13 9 7 9 7 9 7 9 9
6 7 15 9 13 13 13
1 13
4 13 11 0 0
10 7 15 9 0 13 13 0 13 9 0
8 7 9 9 15 1 9 9 13
11 0 9 0 13 15 13 9 9 7 9 11
6 7 13 9 1 9 13
1 13
6 0 0 15 1 9 13
9 3 3 13 9 16 13 1 9 15
5 9 3 0 13 0
14 7 13 15 13 1 9 9 15 1 9 7 13 13 9
15 7 15 9 13 1 9 15 13 1 9 13 7 15 9 0
10 7 15 9 1 9 15 13 9 1 9
9 7 13 9 0 15 13 9 0 13
18 7 13 9 9 15 1 9 7 13 9 9 7 13 1 9 9 9 0
18 7 13 13 9 1 9 7 13 9 1 9 3 1 9 9 1 9 12
26 7 13 3 9 0 13 9 7 15 15 13 9 7 9 0 7 9 9 15 13 1 9 0 13 9 9
8 0 7 0 9 15 9 9 0
4 7 1 0 13
28 7 6 13 13 9 9 9 1 9 7 13 12 9 13 12 9 1 9 13 9 9 0 7 13 1 9 9 0
18 7 12 1 12 9 13 12 9 12 9 0 0 9 9 13 1 9 9
12 7 13 13 9 9 1 9 9 7 1 9 15
12 7 15 13 13 1 9 16 13 12 9 12 9
9 7 13 9 0 1 9 13 12 9
28 7 13 0 7 13 9 15 1 9 7 13 13 9 0 7 0 1 9 15 13 9 9 7 15 15 13 9 15
13 7 0 13 9 15 1 9 7 13 13 9 3 0
15 7 0 13 9 15 1 9 7 1 9 9 7 13 13 9
5 7 13 9 9 13
2 0 13
4 7 13 9 13
9 3 9 9 0 0 7 0 9 15
22 7 13 9 9 0 7 13 9 9 13 9 1 0 9 3 7 13 9 16 13 0 9
8 7 0 13 9 15 1 9 9
12 7 13 13 9 15 0 7 13 9 15 1 9
10 7 0 13 9 15 1 9 0 0 11
11 7 13 9 15 16 13 9 9 1 9 9
19 7 13 1 9 9 7 1 9 9 7 1 9 9 9 12 0 1 9 9
21 13 3 9 9 13 9 7 13 1 9 0 9 13 0 1 9 1 9 0 9 0
14 0 15 13 7 13 9 15 16 0 13 7 13 9 15
9 7 13 0 1 9 15 13 3 11
16 7 0 13 9 15 1 9 7 13 9 0 1 9 1 9 13
2 13 13
4 7 9 9 13
15 7 11 0 13 1 9 1 9 13 15 9 9 9 9 15
9 7 15 9 13 7 9 3 13 13
16 7 13 12 1 12 9 15 13 12 9 7 13 13 15 1 13
16 13 15 9 9 0 15 13 1 9 0 1 15 13 13 9 9
10 7 13 13 15 13 9 1 9 9 15
7 7 13 15 1 9 1 9
16 7 13 9 13 1 9 0 0 9 9 13 9 12 7 9 12
6 7 1 9 15 9 13
7 11 0 9 9 7 9 9
8 7 13 13 16 13 0 9 0
4 7 13 15 9
2 3 13
17 15 15 13 9 9 7 9 15 13 15 15 13 9 12 7 12 9
16 9 15 13 13 7 3 13 7 13 13 1 9 7 1 9 13
22 7 13 13 9 15 3 13 13 9 1 9 9 1 9 9 13 9 16 13 7 3 13
13 12 9 12 9 13 1 15 9 13 7 9 12 13
2 12 13
3 15 3 13
8 7 16 13 13 0 0 9 13
8 7 1 12 13 7 1 9 13
8 7 12 9 15 13 12 9 13
13 15 9 3 13 7 9 3 9 12 9 13 1 9
12 7 1 0 13 15 9 13 1 9 13 9 0
23 7 13 7 13 15 1 0 9 9 15 1 0 13 13 7 1 9 13 16 13 9 9 15
22 7 9 15 9 9 13 1 15 7 15 0 7 0 13 1 15 7 3 0 3 3 13
19 9 0 15 0 13 13 1 15 3 13 1 9 9 15 13 7 13 7 13
15 7 9 9 7 0 7 9 13 7 9 3 13 1 15 3
10 7 15 9 15 9 3 13 1 15 3
8 7 9 9 3 13 1 15 3
11 1 0 13 3 9 0 9 0 1 9 13
7 7 9 15 13 1 9 9
5 9 3 9 13 0
11 0 15 1 9 9 9 13 13 7 13 15
12 7 1 9 15 13 9 0 16 1 15 13 9
23 7 13 9 7 9 9 7 9 15 13 1 13 9 1 0 15 13 1 9 7 1 9 15
15 7 13 9 13 1 9 13 9 9 7 9 0 1 9 15
14 7 13 13 0 1 0 15 13 13 1 9 1 9 15
14 7 15 3 13 13 1 9 9 13 13 13 1 9 9
7 7 13 9 0 1 9 13
26 0 3 7 0 7 0 7 9 7 9 7 0 7 9 7 15 9 9 0 13 1 9 13 9 7 9
24 7 13 15 1 9 1 9 0 7 0 7 13 15 9 0 11 13 1 9 1 9 13 9 9
14 7 9 1 9 13 13 7 9 15 0 13 15 3 9
12 7 9 3 13 9 3 7 9 16 13 1 15
6 7 13 9 1 9 15
10 7 9 9 13 9 15 7 9 1 0
8 7 13 9 7 9 9 1 0
13 7 9 9 7 9 1 0 13 7 9 15 13 0
14 16 15 13 1 0 13 9 1 0 9 13 1 9 0
29 7 16 15 13 1 9 9 9 0 13 9 9 15 1 9 9 7 1 9 0 7 1 0 15 13 13 1 9 0
3 13 1 9
32 3 13 13 1 15 9 3 15 3 9 10 1 15 13 13 7 13 9 0 0 0 7 3 0 7 1 9 13 9 0 9 11
16 0 3 9 3 15 9 13 13 13 1 0 9 3 13 9 9
17 1 0 3 9 16 13 3 3 13 9 0 10 15 15 1 13 13
4 3 3 15 13
18 13 3 1 0 9 1 9 9 3 12 12 3 1 9 10 15 13 0
10 10 3 9 15 13 13 16 13 9 13
30 0 13 3 9 0 7 0 1 15 9 11 13 13 0 9 16 0 11 13 1 9 9 7 13 3 12 9 7 12 9
15 0 13 3 9 1 15 13 13 9 15 9 3 1 3 13
9 3 9 0 3 13 13 1 10 9
28 0 3 9 10 13 1 15 9 10 9 13 3 0 11 16 13 9 9 15 3 13 13 15 9 1 9 1 9
4 3 3 13 13
29 15 3 13 1 0 9 3 13 1 11 13 9 9 3 13 16 1 0 13 9 10 9 7 3 13 15 1 9 9
9 9 3 10 1 9 3 12 13 13
5 7 0 9 9 13
21 0 3 10 1 15 9 13 0 9 3 13 9 9 3 13 13 1 0 10 15 13
51 7 16 0 15 15 1 9 13 3 13 13 3 3 15 13 13 3 0 10 0 1 15 13 9 9 0 0 13 15 10 16 16 13 1 0 3 0 10 9 15 13 13 3 1 15 13 7 16 9 0 13
45 0 3 3 0 13 7 1 9 9 13 0 3 13 16 16 15 0 13 10 0 15 0 11 13 15 13 1 15 13 9 9 3 13 3 13 16 1 0 9 0 13 16 3 15 13
19 0 3 16 13 1 9 9 3 13 9 13 7 16 3 13 3 13 3 13
25 15 3 9 3 13 13 9 7 13 1 9 15 13 15 3 3 3 9 15 3 13 13 15 15 9
7 3 3 9 3 13 1 9
23 3 3 13 1 0 9 7 3 3 9 0 1 10 9 7 9 15 3 13 13 13 9 0
36 7 3 3 13 11 9 15 13 9 0 15 13 7 3 1 0 9 16 9 15 13 3 13 16 3 3 7 1 9 13 13 3 0 9 3 13
15 1 0 9 3 3 13 9 16 9 15 13 13 9 13 13
30 9 3 0 13 1 9 10 9 9 0 11 3 13 13 9 1 15 15 13 9 3 13 9 9 1 0 9 15 9 13
8 15 3 9 13 1 15 9 0
48 16 3 13 9 13 1 0 9 7 13 1 9 0 9 6 3 13 9 13 1 9 15 15 0 9 13 9 0 7 9 1 0 9 7 3 3 13 9 7 15 0 15 0 13 13 1 0 9
29 13 3 3 15 9 3 7 3 3 3 15 9 15 3 13 1 9 0 15 13 15 3 7 9 7 9 3 13 13
10 3 3 1 10 9 9 10 0 15 13
14 15 3 13 3 15 3 0 9 7 9 3 13 0 11
38 3 16 10 9 0 11 0 0 13 3 16 3 9 13 3 3 1 9 9 10 15 13 7 1 0 15 0 13 7 1 0 15 1 9 13 0 9 13
31 3 0 9 1 9 15 9 13 7 9 13 7 9 3 1 15 9 16 1 10 9 9 15 9 13 15 3 9 15 13 13
8 3 3 10 0 13 13 0 13
39 3 13 15 9 10 3 13 0 11 16 3 13 1 9 9 16 13 3 9 16 0 10 13 13 9 7 0 9 15 13 7 15 15 3 13 13 13 13 15
68 0 3 15 13 13 9 0 9 16 1 0 9 3 13 15 13 1 9 9 9 15 13 1 9 9 10 0 3 1 15 13 13 10 9 15 3 3 13 1 10 0 1 15 13 7 16 13 0 9 16 3 3 0 13 16 3 15 13 3 0 13 3 16 0 0 15 3 13
30 11 3 7 11 7 9 0 7 9 0 0 15 13 11 3 7 3 3 9 9 0 3 1 15 3 13 16 13 3 13
7 15 3 0 15 0 0 13
31 13 3 15 9 15 13 13 13 3 3 13 1 0 9 9 9 1 15 13 1 15 9 15 15 13 13 15 9 13 1 11
32 3 0 13 9 11 3 13 0 11 9 3 13 1 9 11 9 3 15 13 13 9 13 15 15 3 11 3 13 13 1 9 9
21 13 3 3 9 0 15 13 0 0 11 1 13 9 3 3 0 0 0 15 13 13
16 13 3 3 3 9 7 9 0 7 13 13 0 9 1 9 9
17 15 3 15 7 3 15 13 3 16 3 13 3 0 9 1 9 13
39 13 3 3 3 9 13 3 1 15 9 3 3 3 13 9 7 9 15 13 1 0 9 3 13 0 11 1 12 0 16 0 11 13 1 9 9 1 9 11
25 1 0 3 9 16 3 9 3 13 3 9 0 13 1 9 13 9 1 15 1 15 13 13 0 0
11 3 3 1 0 3 3 9 1 9 13 13
16 13 13 3 3 3 0 9 1 9 11 7 13 12 9 0 9
44 7 3 0 9 13 13 15 13 3 0 13 16 3 15 13 3 9 15 0 13 7 9 15 13 3 13 7 3 1 9 10 15 3 13 9 13 15 13 10 9 15 13 9 9
34 3 3 1 9 0 9 13 15 3 13 16 3 13 9 0 0 9 7 9 1 0 9 3 13 9 15 9 3 1 3 13 7 13 9
12 7 3 3 13 9 9 13 1 9 9 3 0
30 0 13 3 9 15 0 13 1 15 13 13 9 11 1 9 15 13 1 0 9 3 9 13 0 7 9 1 9 9 0
17 1 0 3 9 9 13 0 13 9 0 0 1 15 9 0 9 13
19 9 3 13 3 3 3 13 0 11 3 15 13 9 13 9 9 15 7 0
21 7 1 0 3 9 16 13 9 0 13 3 7 3 16 3 3 13 9 13 3 13
15 7 13 13 9 1 9 3 7 3 3 3 1 9 1 9
15 7 3 16 3 13 13 15 9 1 9 1 9 1 0 10
6 7 3 3 13 3 9
16 7 15 9 3 13 13 9 16 3 3 13 9 3 3 13 13
50 7 16 15 9 3 13 16 1 9 10 0 15 13 1 0 13 15 13 0 9 15 0 13 3 13 9 11 16 11 13 1 9 9 7 13 3 3 0 3 13 1 0 0 9 3 15 0 10 9 13
37 3 1 0 9 0 9 3 13 7 13 9 10 1 15 13 13 9 0 11 1 9 13 3 3 0 9 1 15 13 1 9 0 11 3 15 13 9
4 13 9 9 15
8 9 3 1 15 13 9 0 13
14 7 3 3 0 9 3 13 13 1 9 3 15 13 13
11 3 1 0 9 13 13 3 1 3 9 0
30 15 3 3 13 1 3 13 9 9 15 13 1 0 9 0 1 15 9 0 11 13 9 11 13 9 0 9 3 13 9
23 13 3 9 0 1 0 9 3 13 0 11 1 11 9 11 1 15 9 13 13 9 15 13
23 13 3 3 1 0 9 15 15 9 13 1 15 9 3 1 3 3 9 13 3 13 9 13
17 13 3 9 3 9 11 13 13 0 11 1 9 1 9 13 1 9
16 3 13 15 9 3 13 13 9 10 13 0 11 15 13 15 11
16 3 13 9 10 1 15 13 0 11 9 11 3 13 13 1 11
9 3 13 9 3 9 11 13 9 9
11 13 3 3 10 9 3 15 13 9 7 9
33 7 3 3 0 15 13 13 1 9 0 11 13 13 1 0 9 15 13 1 0 9 15 13 13 9 9 15 13 0 11 13 13 15
27 15 3 15 3 13 3 13 16 3 13 13 0 7 16 13 9 15 9 0 11 15 3 13 15 3 13 13
41 0 13 3 9 3 13 13 9 13 9 9 9 11 1 9 11 16 1 0 9 9 11 13 13 3 15 13 16 0 11 13 1 9 9 7 13 3 7 3 7 3
15 3 3 13 13 16 13 9 7 0 15 13 13 1 9 9
27 3 13 13 15 7 10 9 1 15 13 1 11 13 3 9 7 13 13 0 15 13 9 1 9 11 16 13
26 3 3 0 9 13 3 1 0 9 3 0 15 3 1 9 7 9 13 1 9 9 1 9 13 3 13
12 15 3 15 13 13 1 9 15 13 3 3 13
68 7 16 3 9 1 15 9 13 13 3 13 1 0 0 7 0 15 1 15 13 13 13 0 7 3 13 16 13 15 9 15 15 9 3 13 3 3 3 10 15 0 3 13 9 13 15 15 9 13 1 15 9 0 9 13 7 3 1 15 9 13 15 15 3 1 9 0 13
21 0 3 1 10 0 15 1 9 9 7 1 0 9 13 13 13 15 3 1 11 13
5 15 3 0 9 13
23 7 3 3 16 13 11 15 13 1 9 9 12 12 7 12 3 15 13 3 1 13 9 13
22 7 0 9 3 13 13 3 1 9 15 13 1 9 11 3 3 13 13 3 3 0 13
11 9 3 3 3 3 13 7 0 9 13 0
25 0 3 15 3 13 13 1 9 15 9 15 9 7 9 13 1 15 9 15 13 7 3 13 1 9
5 9 3 9 9 13
24 3 7 3 3 1 0 9 1 9 0 13 9 3 15 9 13 13 1 0 9 3 9 0 13
25 1 0 3 9 1 1 9 13 13 1 15 9 3 13 1 9 13 7 3 3 3 13 15 1 9
46 9 3 11 13 1 9 9 11 3 1 0 9 13 13 1 9 15 13 15 13 3 1 0 9 3 1 1 9 13 7 13 15 3 1 9 0 7 3 15 3 9 15 15 13 13 13
16 9 3 11 1 0 9 3 13 13 1 9 0 11 13 9 15
19 1 11 3 16 13 3 15 13 3 3 3 3 13 16 9 9 0 3 13
90 3 16 9 11 3 13 15 13 15 3 1 11 13 3 16 13 15 9 15 9 11 13 1 11 13 13 16 13 3 1 9 0 15 9 3 1 9 15 3 13 13 11 9 3 13 16 1 11 1 9 11 13 15 13 1 9 15 13 11 15 9 1 9 11 13 3 3 0 9 3 13 15 13 9 11 9 11 15 3 9 11 9 13 7 0 3 3 15 11 13
38 13 3 1 11 15 13 1 9 0 3 1 11 9 9 12 1 9 3 3 1 9 16 1 9 9 13 1 9 7 9 15 15 13 3 1 9 1 9
24 1 0 3 9 0 15 15 1 13 0 13 9 7 9 13 15 0 9 15 3 15 1 9 13
30 3 15 13 13 9 15 3 3 13 13 9 11 3 13 16 3 13 0 3 13 0 3 3 1 3 13 3 3 3 13
10 7 3 13 0 9 16 13 1 9 0
6 3 3 11 13 13 15
16 3 9 13 3 3 13 9 1 9 15 3 3 13 1 9 0
17 3 3 15 1 9 13 3 3 1 15 9 7 9 11 13 13 15
5 3 1 0 9 13
23 3 15 13 9 1 9 0 1 9 9 15 0 13 3 9 11 16 13 9 1 15 13 13
19 11 3 13 13 15 15 13 1 0 9 3 13 13 3 7 3 3 3 11
9 3 0 13 9 3 13 13 9 9
26 11 3 9 15 13 9 11 13 13 15 1 0 9 1 0 3 9 3 3 9 11 13 13 3 9 9
31 11 3 9 15 13 10 9 15 13 3 13 11 9 15 11 13 3 13 13 1 9 11 3 13 9 7 0 15 15 13 9
25 3 0 9 9 13 7 9 7 9 0 0 9 1 15 0 13 3 15 13 3 13 1 9 15 13
16 3 10 9 3 13 11 15 3 11 1 9 11 9 3 0 13
5 3 1 9 11 13
6 9 3 0 3 0 13
8 3 3 9 15 9 11 3 13
15 1 0 9 11 13 9 15 7 9 1 9 11 1 9 11
11 15 3 16 13 1 9 11 1 0 11 13
12 15 11 9 3 9 13 3 16 3 12 9 13
12 13 0 16 3 0 13 1 9 7 0 9 13
10 9 3 0 3 13 13 1 3 0 13
29 3 3 3 15 15 13 3 3 12 9 0 0 1 15 13 12 9 13 0 15 13 13 0 9 15 13 11 7 11
11 3 13 3 16 9 11 1 9 15 15 13
12 7 13 3 3 9 9 15 13 1 9 13 13
8 0 3 13 0 9 1 11 13
18 3 15 15 13 9 0 9 3 13 15 3 15 13 15 15 13 9 9
9 15 3 0 9 15 11 13 13 13
16 3 13 3 0 9 3 3 0 1 9 7 0 13 9 3 3
8 3 3 1 9 9 3 13 13
28 15 3 16 15 13 13 13 7 3 15 13 0 3 13 7 13 1 0 9 15 13 3 3 3 1 10 9 9
46 3 3 0 15 0 0 9 13 3 16 11 3 13 16 9 11 13 15 3 0 16 1 0 13 13 1 15 9 15 1 11 7 13 15 15 16 0 13 3 7 3 1 9 11 13 13
20 15 3 3 0 0 13 16 0 9 15 13 1 9 11 3 1 0 9 9 13
27 7 3 3 15 9 3 13 15 0 9 0 7 3 9 9 0 15 3 3 1 0 9 1 15 1 11 13
7 0 3 0 9 1 9 13
26 3 1 0 1 9 13 13 7 3 7 3 13 1 9 13 7 3 13 1 15 9 15 3 3 0 13
18 15 3 3 3 13 9 15 15 1 9 0 9 13 3 1 9 0 13
29 3 3 16 9 0 13 1 11 15 13 1 11 9 15 13 15 13 1 11 1 11 7 3 3 3 13 3 13 9
45 13 3 3 3 1 9 11 9 13 3 1 9 15 13 9 7 9 15 13 9 7 1 9 7 9 0 7 9 0 9 13 3 1 9 9 11 1 9 0 15 13 3 9 9 11
3 7 15 0
10 0 9 13 15 3 13 3 13 9 11
50 7 16 0 9 3 0 13 3 13 15 13 3 11 7 1 11 13 3 16 1 0 13 13 9 15 13 9 11 13 1 11 3 1 9 9 0 11 7 3 3 13 3 3 1 9 11 13 7 3 11
11 13 3 1 11 13 1 9 3 0 13 11
18 7 3 13 3 13 9 1 0 9 11 1 15 9 13 13 1 9 11
21 7 3 1 9 11 9 15 13 3 9 15 1 11 13 13 1 11 15 13 1 11
31 3 13 0 9 7 13 9 13 3 9 13 3 1 11 15 13 1 9 11 1 0 9 1 15 13 9 13 11 13 1 15
33 13 1 9 11 9 11 15 13 1 9 11 1 9 11 7 13 9 11 15 15 13 9 11 1 9 7 13 1 9 0 1 15 13
21 3 3 9 15 11 15 13 1 15 3 13 3 7 1 0 9 15 9 13 13 13
28 3 3 9 0 13 13 15 3 3 0 3 9 11 7 11 7 0 9 11 13 9 1 0 9 9 15 13 11
19 3 3 9 1 9 9 11 7 9 15 3 13 13 1 0 9 1 3 13
10 9 3 0 13 0 1 9 11 1 11
8 3 0 13 9 1 15 13 13
14 7 13 9 11 11 1 11 11 7 11 1 11 12 9
16 0 3 9 13 3 1 9 11 3 11 9 11 13 13 9 9
10 13 3 11 9 15 1 15 3 13 13
25 0 3 13 9 3 13 13 11 1 9 0 9 11 9 9 3 1 9 0 15 13 13 1 9 11
18 0 13 10 9 3 13 0 11 9 9 9 11 3 1 9 1 9 15
23 13 3 9 15 11 1 0 9 3 7 3 3 3 9 15 7 3 9 15 13 1 9 11
13 7 3 1 9 13 13 9 7 9 9 13 13 3
35 15 3 15 3 9 13 16 3 1 9 13 13 13 3 3 13 9 3 13 9 0 1 9 13 3 9 12 13 1 9 7 3 13 3 9
13 0 3 9 13 9 3 13 3 1 9 13 13 13
14 7 3 3 16 13 9 13 13 13 16 13 1 9 11
5 13 3 15 0 9
31 16 13 13 9 15 13 1 9 15 13 15 13 11 9 11 13 13 13 16 3 13 9 15 13 16 1 9 13 3 9 0
20 15 16 13 15 3 0 13 13 13 7 3 13 1 9 13 13 9 15 15 13
8 7 3 7 15 3 13 1 11
12 9 3 0 13 3 3 0 7 15 3 9 13
10 0 3 0 9 13 13 15 13 3 3
8 3 3 1 9 15 13 15 13
19 3 3 1 9 7 9 1 0 13 1 9 9 0 0 3 7 0 9 0
19 3 13 15 3 3 10 0 9 15 3 13 15 13 0 9 0 7 0 9
3 3 0 13
12 0 13 9 15 13 0 11 9 11 1 0 9
26 0 3 7 1 0 9 0 15 3 13 1 9 0 15 3 13 13 15 9 13 13 15 1 13 9 11
26 3 3 13 1 0 9 13 1 9 9 11 15 13 3 13 3 3 16 9 15 0 13 1 9 13 13
15 3 3 13 0 16 9 3 13 13 1 9 3 3 13 13
21 1 15 9 1 0 9 3 9 13 13 9 3 3 0 3 9 13 3 9 13 13
8 3 3 13 0 0 15 13 0
2 15 13
24 3 13 13 0 11 1 9 16 3 13 13 9 0 15 9 13 16 0 13 15 1 9 13 13
10 3 9 0 3 13 13 1 3 3 13
13 15 3 0 3 0 3 15 13 1 0 15 13 13
22 3 3 3 13 13 9 7 15 15 1 0 9 0 1 9 13 13 3 3 3 13 13
14 3 3 15 13 9 9 15 13 9 7 9 0 13 15
38 16 13 13 9 15 13 13 1 9 11 13 1 9 9 7 1 9 0 1 9 3 3 13 3 13 13 7 13 7 13 15 0 15 13 9 0 15 13
8 3 15 13 3 3 13 13 3
20 3 1 9 10 9 13 9 3 13 11 1 9 0 15 9 1 15 3 13 13
17 13 3 1 3 3 3 11 15 1 11 13 7 3 11 15 1 11
11 3 13 13 9 3 13 15 13 1 9 9
23 1 0 3 9 13 9 11 15 3 7 3 3 11 15 3 11 0 1 0 12 1 3 13
16 1 0 3 10 9 15 15 13 3 9 9 3 1 9 13 13
16 9 3 3 13 9 9 11 13 13 15 15 9 3 1 9 13
11 7 15 13 9 0 16 9 0 3 3 13
5 9 3 10 3 13
8 9 3 0 13 9 0 13 13
16 3 9 16 13 9 15 13 7 3 13 15 1 0 9 3 13
21 3 9 9 0 15 13 1 11 13 15 16 3 15 9 13 1 15 3 13 9 0
15 3 1 0 9 13 13 15 1 3 11 15 13 9 9 11
10 0 3 9 15 15 13 1 9 13 13
8 3 3 3 3 0 9 15 13
22 3 13 13 15 16 1 0 9 3 0 11 7 9 11 1 0 9 13 9 3 13 13
6 3 7 9 3 13 9
25 3 1 10 9 9 15 13 9 15 13 1 9 13 13 13 15 9 13 3 15 13 13 1 9 9
23 0 13 9 1 15 13 11 9 11 11 0 1 13 9 11 7 13 9 3 13 3 13 13
22 7 3 3 13 15 15 13 1 9 9 13 1 11 7 9 15 15 13 13 13 1 11
45 0 3 0 9 13 3 13 1 11 1 13 9 0 9 9 15 0 13 1 0 9 13 3 9 13 15 9 16 3 3 1 0 9 13 16 3 9 13 13 3 9 9 15 13 13
33 3 3 13 13 1 11 1 0 15 3 13 13 9 15 9 13 3 15 3 9 9 13 3 9 1 11 3 1 11 13 1 9 12
19 11 3 13 3 9 11 15 1 13 13 11 1 9 11 1 9 11 7 11
26 1 15 9 13 13 1 9 11 9 9 0 3 7 0 13 9 7 9 16 9 0 3 13 7 0 3
11 3 1 0 9 9 13 0 15 13 3 11
26 1 0 3 9 15 13 1 0 9 13 1 0 9 13 9 3 3 0 7 13 3 13 13 9 7 0
16 3 3 1 0 9 13 7 3 1 9 0 9 13 9 0 0
8 3 3 1 10 9 9 0 13
18 0 13 9 9 11 15 13 13 3 11 3 3 13 9 11 13 0 9
25 3 1 0 9 15 13 0 9 13 1 9 15 9 15 13 9 13 15 9 3 13 0 9 8 11
20 3 0 13 9 3 13 11 9 9 0 15 13 9 7 9 3 13 13 15 13
27 3 3 3 0 13 13 1 9 7 6 13 13 13 0 9 0 9 7 9 15 15 3 13 13 3 1 9
32 3 16 13 3 1 9 3 13 13 9 3 13 13 0 9 1 9 0 11 13 13 3 9 12 0 9 0 7 3 13 9 13
36 16 3 13 13 15 0 0 9 3 0 7 1 9 3 13 15 13 15 0 9 13 1 9 15 9 7 9 0 3 3 13 9 0 9 0 13
5 3 0 1 15 13
14 16 3 13 3 0 13 1 9 3 13 15 0 0 9
26 3 3 3 3 16 15 3 3 15 13 13 9 7 9 3 13 3 7 1 9 7 9 0 9 3 13
36 3 6 0 9 15 13 13 1 9 11 7 9 0 0 13 15 9 13 13 0 11 1 9 11 9 9 13 1 11 3 15 13 0 11 9 11
21 3 3 16 13 13 13 13 0 11 1 11 1 11 13 1 15 3 3 13 0 9
5 3 13 0 0 9
6 6 3 13 1 12 9
9 3 16 13 6 3 9 13 15 3
17 3 3 9 15 13 13 7 13 16 13 15 1 9 3 3 13 13
36 3 3 13 13 1 15 9 3 1 9 0 16 13 3 1 9 0 3 0 3 13 15 1 0 9 9 0 3 7 0 15 1 3 0 9 13
6 3 13 15 0 0 9
23 1 3 0 9 3 3 13 0 9 3 8 8 8 8 15 13 15 15 13 3 9 0 11
17 3 7 0 9 0 9 1 0 9 13 13 15 16 13 1 0 9
39 3 3 3 1 0 9 3 3 1 0 9 13 13 9 7 13 13 0 9 13 3 9 0 7 0 15 9 15 13 13 3 1 9 0 13 3 3 3 13
62 0 3 9 0 13 15 3 16 3 1 0 9 3 1 9 15 13 13 1 0 9 15 13 1 9 15 13 8 11 15 1 0 9 13 3 13 3 1 9 1 9 7 9 13 9 7 9 7 3 1 9 3 1 9 0 11 13 3 15 15 13 13
34 7 3 3 13 3 1 9 11 1 9 9 0 16 3 15 9 13 3 1 3 13 9 0 9 11 15 13 11 3 0 13 9 11 11
24 3 13 3 3 1 3 9 1 15 13 0 0 7 3 13 9 0 11 15 9 1 9 9 13
13 7 3 3 7 3 9 9 13 1 9 13 9 15
13 7 3 1 0 9 13 9 15 9 3 15 13 9
19 3 15 3 13 3 0 13 13 15 13 0 9 3 0 9 3 9 15 13
7 3 3 13 0 1 9 13
13 3 13 15 0 15 15 1 9 13 15 13 9 9
14 3 0 9 15 13 1 0 9 13 1 11 0 13 11
25 7 3 3 3 9 9 13 15 15 3 13 0 15 13 13 13 3 3 13 13 9 15 3 0 9
29 7 3 3 13 9 0 9 1 3 1 9 0 3 1 1 9 11 13 13 15 9 0 7 0 3 15 13 1 0
46 15 0 9 9 9 3 13 1 3 9 15 13 1 9 13 15 7 13 1 9 11 16 13 9 7 9 9 0 1 15 15 13 13 16 13 1 0 9 15 15 13 13 3 3 13 13
10 15 9 16 13 13 13 1 9 15 11
38 15 11 1 3 1 0 9 13 13 0 9 15 13 3 3 16 9 1 9 3 13 1 15 9 7 3 3 13 13 9 13 13 3 16 9 1 9 13
14 0 3 9 15 9 13 15 13 3 13 0 3 1 3
22 13 3 3 3 9 13 9 3 13 13 1 11 9 13 1 0 9 1 15 13 12 9
85 3 1 9 9 13 0 9 16 3 12 9 0 13 1 15 1 11 13 13 3 15 9 0 1 15 9 9 15 13 7 3 3 13 1 9 9 13 13 13 9 16 3 1 11 11 13 1 13 0 9 15 3 0 7 3 0 9 13 13 16 3 13 13 3 7 3 3 3 9 9 1 9 0 11 9 3 9 0 0 13 13 15 13 1 11
23 15 15 3 13 16 1 9 13 9 15 11 13 13 1 9 15 1 11 9 1 11 9 13
13 3 9 1 0 9 1 11 9 3 13 0 9 13
38 3 15 13 13 9 15 16 15 0 13 15 3 15 13 3 9 9 15 3 3 1 9 0 15 13 1 11 13 7 0 9 1 11 0 7 0 9 13
26 7 16 0 9 3 0 7 0 13 7 0 15 3 15 13 3 13 9 16 3 3 3 3 13 9 11
31 3 3 13 1 11 1 0 9 1 9 9 13 1 9 11 1 15 3 3 13 13 13 9 0 11 7 0 7 3 0 13
35 3 3 16 3 13 15 9 13 7 9 3 3 0 7 3 13 13 3 3 3 0 9 7 3 1 9 9 13 9 11 13 13 9 11 11
26 7 3 3 13 9 1 9 15 13 1 9 15 9 1 9 13 13 15 13 11 15 9 3 1 3 13
15 3 3 9 1 9 3 0 7 9 7 9 13 7 9 0
7 0 3 9 0 9 9 13
8 3 7 9 3 13 1 9 15
10 3 3 13 13 1 9 11 9 15 11
26 3 3 1 9 13 9 7 0 15 9 13 13 1 9 0 3 7 3 3 3 0 0 0 11 3 13
28 7 3 3 13 1 0 9 9 0 3 7 3 3 0 9 13 15 1 9 15 3 1 9 1 0 9 13 9
69 7 16 0 9 10 9 9 3 0 7 9 7 9 13 15 3 13 15 16 13 15 9 9 9 3 0 9 15 13 16 1 9 3 9 13 1 0 9 3 3 16 3 13 15 9 13 3 0 1 13 0 13 15 3 3 9 13 9 3 7 3 15 13 3 16 13 13 15 13
28 3 3 13 15 3 1 9 11 9 7 3 13 15 9 15 3 0 3 15 13 0 0 9 7 16 1 9 13
15 1 15 11 9 13 1 3 3 13 0 9 3 0 7 0
5 3 13 15 0 9
14 6 9 11 15 16 13 9 13 15 16 13 3 9 9
24 3 13 3 3 9 3 1 0 9 13 15 13 9 15 13 11 3 3 15 13 15 9 1 9
11 7 3 13 15 1 10 9 3 0 9 13
21 15 9 16 13 11 9 1 9 3 9 13 11 1 11 9 3 13 13 1 0 9
10 13 3 0 9 13 9 7 13 9 0
14 7 3 11 9 9 13 1 9 1 15 9 15 3 13
3 7 3 13
17 9 11 15 13 15 16 15 9 13 9 0 7 6 3 9 13 15
35 15 16 13 13 9 13 9 10 13 9 1 3 0 9 13 13 1 9 3 1 9 9 16 3 3 13 9 3 16 3 0 9 1 9 13
17 7 3 3 9 13 13 16 3 9 13 7 13 1 9 0 0 9
19 3 3 16 13 15 15 9 13 13 1 9 13 9 15 13 15 1 9 13
17 3 9 0 15 13 9 1 9 0 1 0 9 15 0 9 9 13
21 3 13 0 9 13 10 9 1 9 7 13 15 9 1 10 9 3 15 9 13 13
25 1 0 3 9 7 1 0 9 15 13 9 9 3 0 9 15 13 1 0 9 9 9 1 3 13
12 1 0 9 0 9 3 1 3 13 3 9 9
31 0 3 9 15 9 13 3 13 13 1 0 9 16 3 15 13 7 12 9 15 13 15 13 9 3 3 3 3 1 3 13
11 3 3 3 3 15 9 3 13 3 1 3
19 7 3 13 9 15 0 13 13 3 13 15 3 13 1 15 15 13 1 11
15 15 9 11 3 1 0 9 13 13 3 3 3 13 3 13
16 3 9 0 13 1 0 9 16 9 3 13 3 1 0 9 13
37 7 16 0 9 1 0 9 13 3 0 11 9 15 11 15 13 0 15 9 13 1 9 13 0 9 13 1 0 9 3 3 16 0 9 1 9 13
10 16 3 0 15 13 0 9 13 1 15
15 13 3 1 9 1 15 13 13 11 9 1 0 9 15 13
24 16 3 13 1 9 10 13 9 13 9 7 13 15 3 10 9 7 3 13 15 13 13 3 9
47 0 3 13 15 0 10 13 3 16 1 0 9 15 11 9 1 10 9 13 13 1 9 9 3 1 0 9 13 16 15 0 16 15 0 1 10 9 13 7 3 9 15 0 13 1 10 9
21 13 3 15 3 1 10 9 0 15 13 3 9 11 7 16 15 3 9 13 13 15
28 7 16 1 9 9 15 13 3 0 15 13 13 16 3 3 15 1 15 13 16 15 3 0 1 15 1 9 13
7 3 3 0 13 15 3 13
15 3 16 9 15 11 13 7 13 1 9 13 15 9 9 15
20 7 3 3 13 3 0 3 15 13 3 1 3 13 3 1 11 16 3 3 13
21 3 1 9 0 13 13 11 3 13 13 0 11 3 13 13 1 11 13 9 1 11
13 13 1 9 15 7 1 9 9 15 7 13 1 11
18 3 3 16 13 15 13 1 11 3 3 13 1 9 15 13 1 9 10
28 13 3 3 9 9 10 3 0 7 9 9 7 0 7 9 7 9 15 3 15 15 9 3 13 13 13 15 13
30 16 3 13 1 10 9 13 13 9 7 13 10 9 1 11 13 3 12 9 7 13 9 7 3 13 15 9 13 13 3
13 3 13 13 15 13 1 9 0 3 13 9 0 11
5 7 13 15 0 9
19 6 9 3 13 0 11 9 9 0 11 15 13 11 7 0 3 15 13 13
27 3 9 15 13 1 9 9 9 0 3 13 3 9 11 3 3 9 3 13 13 15 13 0 15 9 9 11
88 3 3 0 15 1 9 3 3 13 16 0 7 3 9 9 9 0 3 13 3 3 15 15 9 7 9 3 13 15 3 3 13 15 3 13 13 3 16 0 13 9 3 3 0 13 15 15 15 13 13 7 16 13 15 3 16 1 9 9 7 1 9 0 3 15 13 1 9 15 16 0 13 16 3 9 13 0 7 16 13 15 9 13 9 0 9 15 13
13 3 9 13 3 13 16 1 9 15 3 13 3 13
30 13 3 3 3 9 1 9 9 7 1 9 0 0 15 13 13 1 13 0 3 9 15 13 7 13 1 15 15 3 13
24 1 0 3 9 1 0 9 7 0 9 16 15 3 1 9 13 3 15 0 13 7 3 9 13
39 3 3 15 1 0 9 13 9 10 3 3 9 0 11 13 1 9 0 3 3 0 9 3 1 12 9 1 9 1 0 9 13 9 3 13 9 11 7 11
14 7 16 9 0 9 3 13 13 1 9 13 1 15 13
9 13 15 9 16 13 15 15 13 13
9 13 9 15 13 7 13 15 16 13
3 3 15 13
19 0 11 1 9 11 7 11 9 7 11 9 9 13 1 9 1 0 9 13
37 11 3 7 11 3 13 3 1 0 9 13 3 16 0 3 13 16 3 9 11 16 13 11 9 11 9 11 9 9 15 11 15 13 11 1 11 13
14 3 9 13 13 3 13 1 11 0 11 3 13 1 15
13 11 3 1 15 7 11 3 13 9 9 15 9 13
7 7 3 3 3 13 3 15
26 3 3 9 0 13 16 1 13 0 11 3 13 9 0 11 7 3 0 11 3 13 3 13 9 11 0
22 3 15 13 3 13 9 10 3 0 11 13 9 15 13 11 9 11 0 7 13 15 9
25 1 0 9 13 3 9 10 1 9 15 13 3 9 11 0 7 16 13 13 13 15 1 7 13 15
15 3 3 0 9 3 13 3 0 7 9 7 0 9 13 3
17 0 3 13 1 0 9 3 13 9 10 9 3 13 3 11 1 15
12 9 10 9 15 13 0 9 13 3 3 1 11
28 3 3 3 1 11 9 13 12 7 3 3 1 11 15 13 9 9 15 9 13 12 7 3 3 9 9 3 13
15 0 3 9 3 0 13 15 13 1 9 9 7 9 7 9
16 7 0 0 13 13 13 3 3 0 0 9 7 0 9 13 13
34 15 3 1 9 9 7 0 9 13 15 13 9 7 15 3 13 15 0 13 7 3 15 3 1 9 13 15 3 13 0 3 15 13 9
19 3 13 13 9 15 9 3 15 9 13 3 7 1 9 9 7 9 9 0
25 16 9 3 3 13 13 15 9 1 9 10 3 13 0 11 9 0 11 15 9 0 9 13 1 11
14 1 15 9 9 13 13 3 3 0 9 0 3 7 0
20 13 3 9 1 9 13 9 10 0 3 15 13 0 11 1 9 15 3 3 13
46 7 3 3 13 9 1 9 13 1 9 1 0 9 1 9 15 7 9 9 13 7 15 15 13 13 15 1 9 15 3 13 13 0 9 13 7 13 0 9 15 0 13 1 9 0 13
27 3 3 9 13 13 13 15 7 15 15 15 1 13 3 13 9 9 13 0 3 15 0 9 13 1 9 15
30 7 16 10 9 1 9 0 13 1 1 13 13 15 1 0 9 9 0 3 3 1 12 9 1 9 1 15 9 9 13
15 0 3 9 3 9 13 13 3 9 11 0 15 9 13 11
12 3 13 13 15 1 10 9 9 11 0 9 11
12 13 13 3 15 9 3 13 13 11 9 9 15
34 7 3 3 1 9 9 13 15 13 13 0 9 7 0 9 15 15 3 1 0 9 13 13 13 13 13 1 9 7 9 15 13 1 11
27 7 16 1 11 0 9 15 13 1 11 13 9 0 11 0 13 3 16 3 3 13 3 16 3 1 0 13
15 3 13 1 11 13 1 15 9 1 9 3 11 15 13 11
12 7 3 3 13 9 11 13 1 9 15 13 11
10 7 0 9 13 1 9 15 13 11 11
10 3 16 13 13 1 9 3 0 1 9
9 13 3 3 9 3 0 1 0 9
33 7 16 3 1 0 11 15 9 13 1 9 1 9 7 0 13 1 9 3 12 12 9 13 3 13 3 16 9 15 13 13 3 13
15 3 3 1 0 9 15 15 13 3 9 1 9 9 7 9
7 0 3 9 9 7 9 13
15 15 15 16 13 15 9 0 7 15 13 13 3 7 13 13
30 7 16 13 1 9 9 3 0 13 3 1 10 9 7 1 0 9 0 15 13 9 1 15 13 9 15 9 3 0 13
28 3 3 9 13 13 1 13 9 1 0 16 3 0 13 7 3 13 16 3 13 15 13 1 9 15 3 13 13
39 3 3 16 13 1 9 9 13 9 1 9 3 7 3 3 7 13 15 9 0 11 9 11 9 15 13 0 15 15 13 13 0 7 3 13 1 15 9 13
42 7 3 3 13 3 9 13 3 0 9 7 9 3 9 3 9 15 3 13 7 13 9 7 9 13 13 11 1 9 15 3 13 9 0 1 9 9 13 13 3 9 15
17 7 3 13 0 9 1 9 15 13 11 15 13 1 9 11 3 13
42 7 3 15 9 13 9 11 7 13 9 3 0 1 0 9 15 13 13 15 13 11 11 7 11 13 11 3 1 0 9 0 11 1 3 15 0 3 15 3 13 13 9
35 1 15 9 9 9 15 16 0 1 15 9 13 3 9 13 1 9 11 9 15 1 11 13 15 13 11 1 9 0 7 0 9 11 9 9
33 16 3 3 1 0 1 9 13 16 15 3 9 13 13 7 0 13 16 9 13 13 13 15 9 13 7 3 16 15 9 13 9 13
18 15 3 9 9 15 0 15 13 13 16 7 1 9 7 3 1 9 13
24 16 3 13 9 15 15 9 0 9 3 1 9 0 13 0 15 13 13 13 16 3 13 0 13
35 3 0 9 1 9 9 13 15 9 11 7 13 15 9 7 9 3 3 13 7 3 3 0 7 3 0 1 9 7 9 15 3 13 3 13
15 7 1 0 9 3 1 9 13 9 7 9 13 3 3 9
6 7 1 0 9 13 9
10 3 3 3 13 13 3 13 0 9 13
6 13 3 15 9 15 13
3 3 13 9
6 3 13 9 7 13 0
28 7 1 0 13 9 1 1 9 15 1 9 15 13 7 0 15 12 7 12 13 13 3 7 3 13 9 3 9
17 3 9 0 3 13 15 3 1 11 7 13 9 7 9 16 13 9
39 3 13 7 3 13 7 3 13 1 9 1 11 15 13 1 9 3 3 3 7 3 3 3 13 9 3 13 0 7 3 13 1 1 9 3 15 1 9 13
18 9 3 0 15 13 3 9 3 15 13 9 3 15 15 9 13 1 11
9 13 15 9 7 9 7 13 9 0
8 13 3 9 0 7 3 9 3
18 6 7 13 9 7 13 7 13 3 3 7 3 3 3 9 13 9 15
4 13 9 7 9
29 7 1 3 13 13 1 9 13 15 9 7 13 1 9 15 13 1 9 7 12 1 9 13 9 0 3 13 13 9
11 7 9 13 0 9 3 0 0 13 13 3
3 15 13 15
2 13 9
4 15 9 0 13
19 3 13 9 9 16 15 3 13 9 13 9 7 3 13 9 13 9 1 9
17 3 13 9 7 3 13 9 9 7 13 16 15 13 0 13 9 15
9 3 13 0 9 7 3 13 9 11
7 7 13 9 1 9 13 0
5 3 3 15 9 13
7 3 16 13 13 3 13 9
3 3 13 9
4 3 13 15 9
22 7 1 0 3 3 9 3 15 9 13 3 1 9 7 3 3 3 13 3 3 1 9
17 7 3 1 9 9 13 3 1 11 3 3 1 9 3 3 1 9
22 9 3 0 0 3 0 13 7 9 0 13 3 1 11 3 3 1 9 7 3 1 9
13 0 9 3 1 9 12 3 13 1 9 7 1 11
39 0 3 9 15 13 0 9 1 9 9 13 15 15 9 15 13 13 1 0 9 7 3 1 9 1 9 15 13 9 1 11 3 3 3 9 1 0 0 13
14 16 3 13 16 1 9 9 3 13 3 13 7 3 13
16 7 13 9 3 7 3 3 9 7 13 9 1 0 9 7 9
18 3 7 9 7 9 3 13 13 1 0 9 1 9 1 9 15 15 13
14 16 3 0 9 13 3 13 9 7 13 1 9 1 11
27 13 9 15 7 13 15 9 1 11 3 3 9 0 13 7 3 13 13 9 13 9 15 1 9 7 13 15
6 3 13 9 15 1 9
17 3 13 9 13 7 0 9 1 15 9 13 7 3 9 7 9 15
22 13 3 0 12 9 7 13 9 12 6 3 9 13 1 9 11 16 0 9 11 13 9
19 7 3 3 13 9 1 9 13 9 7 13 1 9 7 13 9 9 9 0
26 15 16 13 13 0 9 7 9 13 15 9 7 0 9 16 3 0 13 13 1 9 9 1 15 0 13
16 13 3 9 13 9 7 13 1 9 1 9 7 15 9 1 0
6 3 13 0 7 13 9
34 3 3 13 15 9 1 9 15 7 3 1 0 9 13 15 9 1 11 7 9 13 7 9 3 1 9 7 1 0 9 7 9 13 9
11 9 3 3 9 7 9 13 1 11 1 9
14 1 0 3 9 7 9 16 15 13 3 1 9 9 13
11 16 15 13 13 1 9 15 7 13 15 13
33 1 9 3 16 0 9 13 7 13 1 9 0 15 13 11 15 9 1 11 13 1 9 7 13 15 1 9 15 3 3 13 9 0
21 3 3 3 9 3 13 16 1 15 9 15 13 15 13 13 7 1 0 15 9 13
17 15 9 3 3 0 9 13 16 3 13 9 1 9 7 1 9 9
13 16 3 13 9 13 1 9 13 15 9 1 9 11
8 13 15 9 0 3 3 9 3
14 7 3 3 13 9 13 9 7 3 13 1 9 9 9
10 3 13 9 9 7 3 13 9 1 15
23 3 13 9 9 16 13 9 15 15 3 13 7 3 13 15 9 13 1 9 0 7 3 13
7 13 3 9 15 1 9 13
13 7 3 13 16 3 3 1 0 7 0 9 13 9
9 3 3 1 9 3 13 1 9 0
49 0 3 1 15 3 0 13 15 13 16 9 7 9 0 3 13 3 15 9 13 3 15 3 3 3 3 15 1 9 7 0 7 0 7 1 9 3 3 0 7 3 0 16 1 10 9 13 15 13
40 7 16 0 9 3 0 9 1 9 0 13 15 13 15 1 11 13 15 13 1 9 15 13 11 12 3 9 0 15 13 0 1 9 1 11 13 3 3 13 13
17 3 3 1 11 16 16 13 9 0 3 13 13 3 9 1 9 0
6 0 15 13 1 9 9
4 7 0 15 13
32 7 16 1 9 15 9 13 3 13 3 13 7 3 13 1 11 0 9 15 13 9 9 13 13 15 13 3 9 16 3 9 13
20 3 16 13 13 3 3 1 11 13 9 7 15 1 15 3 9 3 1 9 13
5 13 3 3 12 9
2 3 0
13 13 15 9 7 13 15 15 1 9 15 16 15 13
10 9 3 3 1 9 3 13 7 9 13
19 3 3 3 13 15 9 9 13 0 13 15 15 1 9 0 15 13 1 11
17 15 3 9 13 0 9 9 7 11 7 9 7 1 11 0 13 13
10 3 1 9 7 9 7 9 15 15 13
8 3 7 16 9 13 0 0 13
9 9 3 15 9 0 0 13 0 9
39 3 15 13 1 9 9 0 15 11 1 0 9 15 1 15 9 9 15 13 13 9 9 7 9 0 3 9 0 3 11 7 1 9 7 0 9 0 1 11
17 7 16 13 1 9 13 3 0 9 9 1 9 0 15 13 1 11
38 7 16 16 13 7 13 0 9 7 13 9 15 3 0 10 9 7 3 3 16 9 9 13 13 13 1 9 1 11 1 9 7 3 13 9 3 0 9
11 0 3 9 3 3 1 9 1 9 0 13
10 15 3 9 3 1 10 9 13 1 11
5 0 0 3 0 9
36 0 9 1 11 15 13 1 9 15 13 1 9 9 0 3 3 15 3 13 7 3 13 3 0 9 1 11 15 13 1 11 3 1 12 12 9
4 0 9 1 11
4 0 9 1 9
20 7 3 3 1 12 9 0 15 9 7 0 9 13 1 15 9 0 15 3 13
32 1 11 3 1 0 12 9 3 0 9 13 7 10 9 13 1 9 7 1 15 9 0 9 7 1 9 15 1 0 9 13 13
40 3 1 10 9 15 15 9 1 11 13 1 9 3 9 0 9 15 13 3 1 9 1 9 1 11 13 9 7 9 13 16 9 3 13 0 9 3 1 11 3
23 1 9 3 7 9 0 9 0 9 15 3 13 1 11 3 3 9 7 3 0 9 7 9
22 3 0 9 9 13 1 11 7 15 13 7 9 15 13 15 1 0 9 7 3 1 9
47 13 3 15 9 7 3 9 3 1 0 9 13 9 3 0 9 13 9 1 9 11 7 11 7 13 15 11 7 11 9 9 11 7 1 9 15 15 13 13 9 7 1 9 10 15 13 9
15 7 3 13 15 1 9 15 9 13 13 9 7 3 13 9
15 3 3 1 15 0 1 9 13 3 3 12 9 13 1 9
24 3 3 12 9 13 16 0 9 7 9 3 13 13 12 9 9 15 9 0 13 7 3 13 13
11 1 0 3 9 3 3 3 0 9 9 13
36 7 3 3 1 12 9 13 12 9 0 7 12 9 16 3 13 12 9 13 3 3 13 13 9 12 7 12 15 13 15 3 13 9 15 13 0
28 3 3 3 3 3 0 9 13 7 13 15 0 9 9 13 13 1 9 0 15 13 9 15 13 1 11 1 9
16 7 3 9 1 9 13 1 11 13 1 9 3 3 0 9 13
8 0 3 16 13 13 15 9 0
19 9 0 0 9 15 13 3 3 1 11 7 1 9 3 3 0 9 0 13
21 3 0 9 3 1 9 0 1 11 13 3 3 0 9 7 13 3 1 3 15 3
27 3 1 0 13 1 11 7 13 15 0 9 1 0 13 13 16 1 9 0 3 0 13 16 3 1 0 13
21 3 1 0 7 0 7 9 3 13 3 9 13 1 0 9 13 3 1 10 9 0
17 0 9 3 3 13 1 3 1 11 7 13 15 15 3 3 1 3
7 3 3 1 0 7 1 0
40 1 0 3 16 9 13 3 15 13 0 9 0 9 7 0 9 1 0 1 11 13 16 1 0 9 13 16 9 9 13 3 0 7 0 9 3 3 1 9 13
7 7 3 1 0 1 11 13
19 3 16 3 1 0 9 9 13 0 9 7 0 9 7 1 0 1 11 13
12 3 16 3 9 13 9 7 9 7 9 13 3
14 16 3 13 13 9 3 1 9 9 13 9 3 1 11
16 3 13 9 7 9 13 9 7 13 9 0 1 11 7 1 9
16 9 3 9 1 0 9 15 13 0 3 13 3 3 1 0 9
12 0 9 3 3 15 13 3 0 9 7 0 9
26 0 9 3 3 15 13 3 0 9 7 3 1 0 1 11 13 7 3 3 1 9 3 1 11 13 9
35 7 0 9 9 1 11 13 1 0 9 15 1 11 13 13 1 9 3 1 3 15 13 1 9 9 3 13 13 1 15 9 3 15 13 9
12 13 3 9 1 11 3 3 16 13 9 1 9
2 9 9
6 15 15 3 1 3 13
26 9 3 15 13 9 1 11 1 9 13 0 13 9 16 0 9 15 13 9 13 3 9 1 11 13 13
6 3 3 0 9 13 0
11 15 3 13 3 13 9 9 15 13 1 9
10 3 13 16 3 13 0 15 13 3 0
27 3 0 9 13 3 9 1 0 16 0 15 13 0 15 13 15 13 9 0 9 16 9 0 13 9 16 13
15 7 3 13 0 9 3 3 13 3 9 3 16 13 1 11
38 9 3 9 3 0 13 1 0 16 15 3 13 0 9 1 9 15 13 9 0 7 0 3 3 13 1 0 9 3 9 13 1 9 11 0 15 13 9
35 9 3 16 13 3 3 3 3 13 7 1 15 9 15 13 0 13 1 9 9 9 0 7 3 7 3 3 3 13 3 9 13 3 3 13
30 9 3 3 0 13 16 15 15 13 3 3 13 9 9 7 9 3 3 9 0 7 3 0 9 3 13 3 1 9 13
25 16 15 3 13 1 10 9 15 3 13 13 0 9 9 3 3 13 1 0 0 1 0 0 9 13
10 15 3 3 0 13 0 13 1 0 0
9 15 3 3 0 1 0 1 0 13
13 15 3 13 15 13 13 7 12 15 3 13 15 13
13 3 7 0 13 15 3 13 3 7 0 13 15 0
34 9 3 15 0 9 0 13 16 3 7 9 15 13 3 13 3 7 9 13 3 7 15 15 1 9 13 7 3 9 7 9 0 1 9
7 0 3 9 3 13 3 13
31 7 13 0 9 9 0 9 9 1 11 13 1 9 9 0 9 3 1 11 13 1 9 3 1 3 9 3 9 13 1 11
17 3 0 9 7 0 7 0 7 0 7 0 3 13 3 0 1 0
41 0 3 9 16 13 15 13 3 3 12 13 1 0 16 9 13 0 9 15 3 3 13 3 3 0 9 15 13 3 3 16 9 15 1 10 12 9 1 11 13 13
22 0 3 9 15 13 0 9 1 11 13 9 1 9 0 15 1 11 13 13 1 12 9
13 13 3 0 9 0 9 3 7 9 3 9 3 9
16 3 3 3 13 15 3 13 9 13 13 9 7 13 9 3 9
13 7 3 3 16 13 15 9 0 13 15 1 11 13
11 11 3 15 13 11 13 3 0 9 1 9
27 13 3 1 11 1 11 3 1 12 9 1 0 9 9 13 1 9 1 0 9 1 15 13 9 11 9 11
30 3 3 16 13 9 13 0 15 9 7 9 3 13 13 12 9 7 12 9 7 13 10 9 1 9 3 13 9 11 9
15 7 3 13 9 7 13 15 3 3 3 1 11 1 9 13
25 1 11 3 16 13 13 3 15 15 9 13 16 3 3 0 9 7 3 9 15 1 9 0 13 9
10 13 9 3 7 9 0 10 9 7 9
34 3 3 16 13 9 13 9 15 13 13 9 1 0 9 7 13 10 9 15 13 13 1 9 16 13 11 1 11 1 12 9 9 7 0
21 3 3 0 9 0 13 16 3 1 9 13 13 1 12 9 9 13 0 13 1 11
16 1 9 3 3 1 0 9 15 1 9 3 13 9 12 9 13
13 13 3 15 1 9 3 1 11 7 13 9 1 9
46 15 3 9 15 13 0 15 13 1 9 0 15 3 13 9 0 13 1 9 9 0 15 9 13 1 11 7 1 9 3 1 3 13 9 3 0 3 13 1 9 1 9 0 15 13 9
19 3 3 9 13 16 1 11 13 15 13 1 9 3 9 13 13 7 3 9
20 16 3 13 13 15 1 9 1 9 0 7 16 13 9 13 9 9 7 13 3
6 3 13 9 0 7 13
8 3 15 9 0 1 11 13 13
18 9 3 0 15 9 13 1 9 9 15 13 1 11 1 9 7 3 9
9 13 9 7 9 0 9 10 7 9
3 9 3 3
26 7 16 13 15 13 9 0 13 1 9 1 11 15 13 1 0 9 1 15 13 9 1 9 7 3 13
14 3 15 9 3 0 9 13 13 3 16 9 0 13 3
6 3 3 9 13 7 9
21 7 3 16 13 13 9 0 13 10 9 1 9 3 9 1 9 7 9 13 9 13
6 0 15 13 1 9 9
9 3 3 1 0 9 9 3 9 13
11 3 0 9 1 0 1 9 7 9 13 3
6 0 15 13 1 9 9
30 7 3 13 9 1 0 9 3 3 15 9 13 3 13 16 0 13 1 9 0 9 15 13 15 9 13 15 9 15 9
45 7 1 0 9 3 1 9 7 3 1 11 1 0 9 3 9 15 7 3 16 15 9 13 7 16 15 9 3 13 9 13 7 3 3 7 3 16 13 9 3 3 3 13 1 11
18 3 16 13 13 16 3 13 3 13 9 13 3 9 1 9 7 13 9
20 3 15 9 15 13 0 9 13 15 9 13 1 9 0 13 3 1 3 1 11
12 3 3 1 0 7 1 0 13 15 15 0 0
7 9 3 0 9 7 9 13
3 13 3 9
8 9 3 13 3 16 13 9 13
12 3 16 13 13 9 3 1 9 1 11 13 9
19 1 15 3 13 13 1 11 13 12 9 13 9 13 9 3 0 7 13 9
9 3 0 9 3 15 13 3 0 9
38 0 0 13 0 9 16 9 3 16 9 13 13 1 9 7 13 13 1 11 7 3 1 11 9 13 13 15 0 9 3 13 1 9 15 13 1 9 11
40 1 15 9 16 13 13 13 9 1 9 1 15 9 13 9 13 9 7 13 9 9 7 13 10 9 13 9 9 15 13 13 1 9 1 1 11 15 13 3 13
6 7 15 0 9 13 9
26 3 3 3 0 13 13 9 13 9 3 3 0 13 9 7 13 1 9 15 1 9 15 3 3 3 9
25 9 3 1 9 13 7 13 9 7 13 10 9 3 11 11 13 1 9 13 15 15 13 16 13 9
25 15 9 3 3 13 13 0 9 7 9 13 0 9 16 15 13 15 13 3 13 1 9 1 0 9
10 3 13 9 13 9 3 0 7 13 9
16 3 0 9 13 15 1 9 0 15 9 13 3 1 3 1 11
6 3 1 0 7 1 0
11 12 3 9 1 9 1 11 13 15 15 9
9 3 3 13 15 9 13 15 13 13
10 3 3 16 13 9 13 9 9 7 13
19 9 0 9 15 1 9 15 13 1 11 13 16 0 9 15 13 3 9 0
22 13 3 9 9 13 1 9 13 3 12 9 3 13 9 7 13 9 3 9 7 13 15
16 13 3 0 9 12 1 0 9 3 13 1 9 3 0 9 3
20 13 3 3 3 9 13 1 11 13 9 13 1 9 9 7 3 0 7 13 9
33 7 3 15 13 13 1 9 15 16 13 16 3 16 13 15 13 1 11 1 9 0 1 15 13 9 1 15 0 9 9 1 9 13
17 7 3 3 1 9 9 3 0 3 7 9 7 9 0 9 7 9
23 9 3 0 1 9 13 1 15 9 13 13 9 0 9 13 1 0 9 15 1 0 9 13
21 7 3 3 9 9 3 0 13 3 1 11 1 9 1 0 9 3 13 9 1 9
12 7 3 3 3 9 7 9 7 9 0 9 13
15 9 3 10 15 13 15 13 9 3 3 9 7 9 0 13
34 7 3 3 16 13 13 9 9 13 1 11 1 9 7 13 0 9 3 13 9 3 13 13 1 9 7 13 3 9 9 7 13 7 0
7 1 0 3 9 9 13 0
28 13 3 9 7 15 9 13 3 9 0 9 7 9 13 3 12 9 0 7 13 10 9 1 9 3 13 9 15
5 13 16 13 1 9
44 7 3 3 1 9 3 1 0 9 1 11 9 1 9 13 3 1 3 0 9 9 7 13 1 9 7 9 0 0 16 3 0 9 3 13 13 3 7 3 1 9 13 1 11
11 9 3 0 3 12 13 13 1 9 15 9
10 16 3 13 13 1 11 13 3 9 0
3 3 13 9
10 3 13 10 9 1 9 3 13 13 9
25 15 9 1 16 13 13 0 9 7 9 0 9 13 1 9 16 3 3 1 9 9 9 15 13 13
11 7 3 1 0 9 13 1 9 9 1 9
11 13 1 9 0 9 15 13 3 9 9 13
16 3 13 9 1 11 3 1 9 7 3 1 0 9 3 1 9
13 1 9 3 3 3 13 13 3 9 3 0 13 13
26 3 3 13 10 9 1 9 3 13 9 1 11 7 15 15 13 13 11 1 9 13 7 1 9 3 13
35 3 3 13 9 9 13 15 16 7 0 9 13 7 3 13 13 0 9 16 3 13 7 13 9 1 9 15 15 1 0 9 0 9 13 13
10 7 3 13 15 3 13 15 13 13 15
40 13 3 3 15 1 9 15 13 15 7 3 7 1 9 3 0 9 15 13 13 3 16 1 0 9 3 1 0 0 9 9 13 13 1 9 15 15 15 13 13
26 1 9 3 0 3 3 13 3 15 13 1 0 9 15 13 1 9 16 9 7 9 3 1 9 9 13
12 3 13 13 3 1 9 15 7 3 0 13 13
16 16 3 13 13 1 9 9 13 1 9 15 9 1 9 0 13
7 9 3 15 1 9 13 13
28 0 3 3 3 13 16 9 13 16 12 7 12 15 9 13 3 0 3 9 13 15 1 9 13 0 9 7 13
30 7 16 13 3 13 15 13 9 7 13 1 0 9 3 3 1 9 15 1 9 13 3 13 16 15 13 13 3 3 13
27 7 3 3 15 9 13 12 7 12 0 13 15 3 1 9 3 1 9 13 9 7 9 7 3 13 9 13
6 9 3 15 13 1 13
10 13 9 11 7 9 10 1 15 9 13
3 13 3 9
2 3 0
30 3 1 9 0 15 9 13 1 12 9 13 1 0 13 16 0 1 0 9 13 1 15 3 15 13 0 9 9 13 13
37 3 3 3 0 9 15 13 3 13 1 9 16 7 9 7 9 13 16 10 9 9 13 15 13 3 9 3 0 7 0 3 15 13 1 9 7 11
11 3 3 15 9 15 13 3 16 3 13 13
19 9 3 9 13 1 9 7 1 0 3 1 0 15 15 13 16 13 9 3
16 13 3 1 9 7 1 9 9 7 1 9 3 1 9 9 13
10 3 7 3 3 1 9 13 9 3 13
8 3 13 1 9 3 13 9 13
39 7 3 1 9 0 3 1 9 0 3 3 13 9 7 13 9 16 13 15 9 16 15 13 9 13 1 9 9 13 3 1 9 3 3 1 9 9 13 13
26 7 3 1 0 12 9 13 9 15 15 13 13 15 3 3 13 13 7 15 13 13 15 3 3 13 13
11 3 3 13 9 15 9 3 0 0 9 13
16 1 0 3 9 7 9 0 9 7 9 0 9 13 16 0 13
20 1 0 16 13 15 3 9 0 13 13 3 10 9 1 9 1 11 3 13 9
7 15 13 3 13 9 7 9
39 3 3 3 9 13 13 1 1 9 3 15 1 9 0 1 9 13 7 13 15 15 1 0 9 1 9 0 15 1 9 13 13 13 3 1 3 1 0 9
8 9 3 13 1 9 13 1 11
5 0 3 13 13 9
2 13 9
3 3 13 9
10 7 3 15 13 1 9 3 15 13 13
10 15 3 3 13 3 13 3 3 1 3
23 9 3 13 3 15 13 15 7 0 13 7 0 7 0 9 13 3 9 7 9 3 1 3
14 0 3 9 13 15 1 3 15 1 0 9 15 3 13
9 9 3 15 9 1 9 13 1 0
18 1 0 3 3 3 13 9 7 13 9 0 1 9 0 15 13 1 9
8 9 3 0 3 13 3 1 15
29 13 9 1 9 11 13 12 9 7 3 13 9 9 1 15 7 3 13 1 9 0 1 15 3 1 9 15 9 13
14 13 3 15 9 13 3 3 1 15 7 13 9 13 9
44 7 1 13 9 9 1 9 0 3 1 9 13 1 11 7 3 3 13 10 9 9 9 13 9 7 3 3 13 9 7 0 1 9 13 1 9 16 3 13 7 3 3 13 9
13 0 3 9 13 9 9 0 9 15 9 3 1 15
29 3 3 10 9 0 3 13 3 3 1 15 7 9 15 13 9 1 12 9 0 3 3 3 13 1 9 3 1 0
46 3 3 0 9 13 7 0 9 3 1 12 9 9 15 3 1 9 3 1 9 0 3 1 11 7 1 9 7 1 11 7 3 1 11 3 7 3 3 1 11 7 3 16 9 0 13
6 0 9 3 1 11 13
4 0 9 1 11
3 9 1 9
14 0 3 9 15 13 0 3 1 9 0 15 13 1 9
40 10 3 12 9 0 3 1 9 9 1 15 9 7 15 9 15 13 15 13 13 7 15 15 9 13 9 7 9 3 7 3 3 3 1 9 15 13 1 11 13
2 13 9
33 13 9 3 1 9 15 1 11 13 1 15 13 9 1 15 13 11 9 3 3 1 11 15 13 1 0 9 1 15 9 13 1 9
18 7 16 13 13 9 7 9 13 13 3 3 1 11 1 9 13 9 9
37 3 16 13 13 13 9 0 9 7 9 13 9 7 13 10 9 1 9 3 0 9 9 1 0 9 3 10 9 3 1 11 13 13 9 13 13 9
26 15 13 3 3 12 1 9 3 3 13 15 13 11 3 13 13 7 13 15 15 9 16 9 13 0 13
4 3 13 16 13
20 0 13 13 3 9 13 9 3 0 7 13 15 1 9 15 3 9 3 9 0
17 3 0 9 15 13 9 0 3 1 0 15 9 1 9 1 11 13
8 3 1 9 15 3 13 3 13
2 13 9
6 13 9 0 9 7 9
8 3 3 1 9 13 1 11 3
8 3 3 3 15 13 15 3 3
18 7 16 13 9 13 3 15 9 7 15 9 13 9 1 9 3 1 11
10 0 3 9 13 1 11 15 9 13 13
23 13 3 9 3 1 11 3 1 9 7 3 15 9 3 1 12 1 9 13 9 3 1 11
11 3 16 13 13 3 13 9 0 9 7 9
22 13 3 3 10 9 1 9 3 0 9 13 13 9 3 13 9 7 13 11 3 0 13
6 7 3 15 0 9 13
18 1 9 3 3 1 0 15 13 9 3 3 15 13 3 15 9 15 13
18 3 3 0 9 3 0 9 3 1 11 1 9 0 3 1 3 0 13
7 3 3 1 0 7 1 9
21 0 3 9 3 1 9 15 13 1 9 0 13 1 9 7 3 13 1 11 1 9
17 0 9 3 7 0 9 16 0 9 3 15 13 1 11 13 7 3
4 13 9 9 15
70 9 3 0 1 9 15 13 0 9 3 15 1 0 15 13 0 9 1 11 13 1 9 13 13 3 9 1 9 1 11 1 15 9 9 13 3 13 13 9 15 9 3 15 13 0 9 0 13 9 9 15 3 16 3 9 7 9 13 13 3 9 7 9 7 3 3 13 15 1 11
31 13 1 11 16 13 9 9 10 9 15 3 0 9 13 15 13 9 9 7 3 3 15 13 1 11 15 0 13 3 0 9
7 13 3 15 15 0 13 13
2 13 9
2 3 9
24 13 15 0 15 13 13 1 9 3 0 9 13 13 7 0 13 9 1 9 16 1 9 0 13
26 3 3 9 13 13 1 9 15 9 3 1 12 1 9 13 9 1 11 7 16 9 0 0 1 11 13
19 3 16 13 13 13 10 9 1 9 9 3 13 9 16 15 9 13 15 13
40 3 9 1 0 0 15 13 13 16 15 13 9 1 11 15 3 9 13 3 3 1 9 9 13 13 9 1 9 3 0 13 13 3 3 13 13 3 1 9 9
18 3 13 9 15 9 13 3 3 7 3 16 13 9 13 9 9 7 13
35 13 3 15 9 15 1 9 15 13 15 7 3 1 9 13 9 9 15 13 1 11 15 3 13 3 16 15 0 13 1 9 15 3 15 13
62 3 3 13 13 1 9 9 15 13 1 11 3 13 1 11 15 13 1 0 9 3 13 9 1 9 7 3 13 9 7 9 13 15 9 13 3 9 13 13 9 13 3 9 0 9 10 7 9 9 3 15 13 3 0 9 13 16 7 9 7 9 13
12 13 3 3 10 9 1 9 3 13 1 9 9
15 13 3 3 1 9 9 3 13 1 9 9 1 9 1 9
37 16 3 0 13 13 13 9 3 0 7 9 3 0 13 3 7 1 9 13 1 10 9 15 3 0 1 11 13 15 13 1 15 9 13 13 9 9
3 13 3 9
2 13 9
5 13 9 7 3 0
8 3 13 3 7 3 3 1 9
17 16 3 13 1 9 9 3 9 13 7 13 9 0 7 12 1 9
31 1 9 3 16 3 13 3 1 9 0 0 13 1 9 3 9 9 3 0 13 16 3 7 3 13 3 1 9 16 13 9
18 7 13 9 0 15 13 1 0 9 15 9 13 1 9 1 9 7 9
10 3 1 11 16 13 13 13 9 7 9
2 13 9
2 13 9
2 3 0
16 7 3 3 15 9 0 3 1 12 1 9 13 9 3 1 11
21 3 16 13 13 13 9 0 13 9 7 9 13 9 13 9 7 3 0 7 13 9
19 9 3 13 13 15 1 9 9 7 3 13 15 1 9 15 9 9 3 0
27 3 3 1 15 9 0 15 13 1 9 3 0 9 15 3 13 13 9 9 7 0 15 3 13 1 0 9
20 3 3 0 9 3 0 13 3 0 9 15 13 16 3 1 9 0 1 11 13
35 3 16 0 9 13 3 13 1 9 0 9 9 1 9 1 11 9 9 9 15 3 0 9 13 7 3 9 7 9 3 1 9 13 1 11
21 16 3 0 9 3 13 3 16 9 7 9 3 1 9 0 3 1 9 13 1 11
3 9 15 13
8 9 3 3 9 13 1 9 0
28 9 3 13 13 3 16 9 13 0 1 15 9 13 0 9 16 3 13 0 1 9 0 13 16 9 13 1 11
4 3 3 1 0
11 3 3 1 9 1 9 3 13 0 9 13
12 0 3 7 0 9 3 0 1 11 13 1 9
12 7 0 3 13 13 3 13 0 15 13 1 9
14 3 15 13 9 15 1 9 0 13 7 15 9 13 9
11 0 13 1 10 12 9 15 13 3 13 0
7 7 3 13 12 7 12 9
6 16 3 9 1 9 15
10 7 3 3 13 9 9 15 15 13 13
5 3 0 9 13 0
3 3 9 13
6 3 0 3 13 7 0
10 3 0 9 15 13 3 0 1 9 13
19 7 16 13 1 9 13 1 0 15 15 13 13 9 13 15 9 15 9 0
8 3 1 9 3 1 9 13 13
17 16 15 3 9 13 16 9 13 15 15 13 3 3 3 13 1 9
11 0 3 9 9 16 13 1 9 13 13 13
28 9 13 3 3 0 16 15 13 1 9 1 10 9 12 15 13 3 3 1 9 13 16 9 13 13 1 11 0
45 7 3 13 9 9 1 9 1 9 0 7 13 15 1 9 1 9 15 13 13 3 9 3 9 13 3 9 9 7 9 3 7 3 3 15 13 13 1 9 15 13 7 13 7 0
14 9 3 3 3 13 3 3 9 13 0 9 15 13 3
18 13 1 11 1 0 9 12 13 15 9 3 13 3 7 3 0 13 3
7 3 7 3 3 3 1 9
4 0 3 9 13
13 7 3 3 13 13 9 12 1 15 13 3 13 9
17 15 9 9 3 3 15 9 9 13 15 0 9 3 3 7 3 3
4 3 3 9 13
37 7 3 13 16 1 0 9 15 0 13 9 3 13 1 9 16 15 13 1 0 9 12 15 13 1 9 0 3 1 9 0 16 1 12 9 13 9
36 9 3 13 9 9 16 0 9 13 0 15 1 13 13 1 9 1 15 15 13 7 13 1 9 3 3 13 7 13 1 9 1 0 15 3 13
30 9 3 13 9 9 3 0 3 3 1 9 13 9 1 11 7 13 9 1 0 7 3 12 9 13 1 9 1 9 12
22 9 3 9 0 15 13 15 13 9 0 3 3 13 15 13 16 13 15 15 3 13 13
27 3 1 9 1 9 13 9 9 7 3 12 7 12 13 9 1 9 15 7 9 1 9 15 7 13 9 9
9 13 3 9 9 13 15 9 7 13
16 1 0 12 9 9 15 13 13 9 3 7 3 3 1 9 13
17 13 3 3 1 9 9 7 3 9 15 9 3 13 3 3 9 13
17 9 3 15 13 9 0 15 13 0 9 16 3 9 13 13 3 13
25 7 16 13 15 1 9 13 16 1 9 9 13 13 1 12 9 0 1 9 13 1 9 1 11 13
11 16 3 9 13 9 9 0 13 15 3 13
8 0 3 9 9 15 13 1 11
8 13 3 9 16 15 9 15 13
17 13 3 9 0 7 13 0 9 13 13 16 3 1 9 13 9 15
17 3 3 3 9 15 13 16 15 3 13 13 1 15 15 13 3 13
52 7 16 1 0 9 9 9 7 3 7 3 13 9 3 15 1 15 3 15 3 9 3 3 3 16 9 16 3 13 3 3 3 13 7 3 3 3 3 13 3 9 15 9 3 13 3 13 16 15 13 15 13
21 9 3 15 1 9 13 16 3 13 3 13 3 13 15 3 13 1 9 16 3 13
32 3 15 3 0 13 15 13 15 3 7 3 3 7 3 13 16 13 7 0 13 15 16 13 15 9 7 9 0 15 3 13 15
42 3 9 9 13 3 0 9 15 1 11 13 15 9 13 13 13 9 7 3 0 9 15 13 1 11 15 13 1 0 9 3 9 13 1 9 0 9 3 0 13 13 9
16 0 3 9 0 9 1 0 9 13 16 9 9 13 13 0 9
32 7 0 1 9 0 13 16 0 9 13 9 15 3 0 11 13 9 9 15 13 13 1 9 9 7 13 3 13 13 1 9 11
9 0 3 9 9 16 13 12 9 13
41 3 1 0 9 13 15 3 13 9 3 3 9 7 9 1 0 9 15 13 3 1 11 7 11 7 1 11 7 11 3 0 9 13 7 3 1 0 15 9 7 9
18 15 13 3 15 3 15 0 9 1 11 13 1 0 9 7 3 0 9
20 0 3 3 9 3 9 0 9 1 9 0 3 15 1 15 9 0 9 11 13
3 7 15 0
25 13 15 0 9 13 15 1 0 9 0 9 13 3 16 3 15 9 0 13 15 9 1 0 9 13
30 0 3 9 9 0 9 15 9 13 15 3 1 9 7 1 9 7 3 1 0 9 0 9 0 13 3 1 9 7 9
36 3 0 9 1 11 15 13 1 9 15 13 1 10 9 1 15 13 9 1 9 1 9 1 15 9 13 9 10 1 15 13 9 9 1 9 9
3 0 3 9
