1219 11
15 10 0 9 4 1 12 9 2 9 7 9 2 11 2 2
8 9 13 15 0 1 0 9 2
10 9 13 1 9 1 9 2 9 2 2
12 3 9 15 15 13 1 12 7 12 9 13 2
11 9 1 9 1 9 12 13 3 1 11 2
23 16 9 1 10 9 13 10 3 9 1 10 9 9 1 3 12 9 4 9 0 1 11 2
9 1 12 9 9 4 9 12 9 2
21 9 4 10 9 2 15 13 1 12 9 1 9 1 9 1 10 9 1 0 9 2
10 3 1 3 9 13 2 13 3 9 2
8 9 1 10 0 9 13 9 2
5 3 13 9 0 2
8 1 9 12 4 9 12 9 2
11 15 13 10 9 1 14 13 1 1 11 2
12 9 2 15 13 9 2 13 1 9 1 9 2
4 15 13 9 2
14 9 4 15 13 15 4 0 9 7 0 3 1 9 2
39 16 10 0 9 3 4 0 3 2 4 15 3 13 9 2 16 15 4 0 3 10 9 15 13 12 7 10 12 9 3 3 2 3 1 9 12 9 2 2
24 1 9 1 0 9 4 1 11 0 9 1 10 9 13 9 2 16 15 13 3 0 0 9 2
5 15 4 13 11 2
15 11 4 15 13 2 15 4 13 0 9 1 3 12 9 2
14 10 0 9 2 1 15 0 9 13 2 4 9 12 2
11 9 1 0 9 7 9 4 13 1 11 2
14 1 0 9 13 3 9 7 3 4 9 3 13 9 2
8 9 4 3 13 9 1 9 2
16 9 13 1 9 0 9 1 9 2 9 7 1 9 1 9 2
1 9
10 7 9 7 11 13 9 1 0 9 2
1 9
3 9 7 9
3 9 7 9
6 1 9 4 3 13 2
1 9
1 9
3 9 7 9
4 9 2 0 2
5 0 9 2 0 2
22 16 10 9 4 0 13 2 16 15 13 7 3 3 13 16 10 0 9 13 0 9 2
5 3 9 13 9 2
8 2 13 3 9 12 3 2 2
1 9
31 9 1 9 4 1 9 12 12 9 1 9 1 10 0 9 7 9 10 9 3 13 9 7 12 9 1 12 0 9 3 2
7 3 13 1 0 9 9 2
9 1 9 13 10 0 9 1 9 2
11 0 9 4 1 9 12 12 9 1 9 2
19 0 9 1 11 13 15 2 1 9 2 16 15 13 0 9 1 12 9 2
31 9 1 9 13 3 1 9 1 10 9 1 10 0 9 1 10 12 0 9 2 13 9 12 2 11 10 0 9 2 2 2
9 0 9 13 12 9 1 0 9 2
30 13 15 0 9 1 3 7 12 9 13 9 1 9 1 10 9 9 2 15 13 2 0 9 9 13 0 9 3 2 2
17 1 9 1 10 0 9 13 9 2 15 13 1 10 9 1 9 2
8 1 9 13 10 0 9 0 2
27 4 15 13 3 9 4 15 13 15 1 14 13 10 0 9 1 10 0 9 1 9 1 9 1 10 9 2
68 2 10 9 4 4 0 2 12 2 12 9 2 12 2 12 9 2 12 2 12 9 2 12 2 12 9 2 12 2 12 9 2 12 2 12 9 2 12 2 12 9 2 12 2 12 9 2 12 2 12 9 2 12 2 12 9 2 12 2 12 9 7 12 2 12 9 2 2
27 16 10 0 9 1 9 12 13 12 9 2 0 10 9 1 3 12 9 2 13 9 12 2 12 2 12 2
6 0 0 9 4 12 2
13 16 9 4 12 9 2 13 0 11 1 0 9 2
11 14 13 13 16 10 0 9 13 1 9 2
22 1 0 9 15 4 0 12 13 0 9 2 13 2 11 10 0 9 2 2 9 12 2
1 9
15 9 1 9 13 15 1 7 1 10 9 15 13 12 9 2
8 9 4 15 1 9 7 11 2
17 9 13 14 13 3 9 7 1 7 1 9 2 3 0 1 9 2
15 7 1 0 9 7 0 9 13 15 3 0 9 1 9 2
17 13 15 9 1 7 9 7 11 4 10 0 9 13 0 9 3 2
5 0 9 13 0 9
8 9 13 3 0 1 0 9 2
7 7 15 13 0 9 3 2
17 9 13 12 9 1 10 9 3 15 1 9 4 0 7 12 9 2
12 15 15 4 13 0 9 1 9 4 13 15 2
15 1 9 13 10 0 9 15 13 9 1 0 9 1 9 2
11 7 3 15 13 3 1 14 13 0 9 2
12 13 16 0 9 1 9 3 4 15 7 9 2
14 2 1 9 4 15 13 1 10 0 9 1 9 2 2
5 0 9 13 0 9
15 15 15 13 1 14 13 3 9 1 1 9 13 0 9 2
18 9 13 1 12 9 1 10 9 15 13 1 9 2 3 3 1 9 2
14 15 13 16 9 1 0 9 4 13 1 3 12 9 2
4 11 10 0 9
4 11 13 12 2
11 9 15 15 13 3 13 3 9 1 11 2
9 1 10 9 4 3 3 9 13 2
19 1 14 13 0 9 1 11 13 1 9 16 15 13 12 9 1 0 9 2
14 1 0 9 15 4 0 15 1 9 12 13 0 9 2
41 3 13 15 15 4 0 12 3 0 9 1 12 9 1 14 13 0 11 2 15 15 4 0 12 13 3 12 9 2 3 2 15 15 4 0 12 13 3 12 9 2
16 15 15 4 0 12 7 3 13 3 13 0 9 1 12 9 2
8 15 4 3 3 13 0 11 2
25 9 12 4 3 13 3 12 1 0 9 2 9 12 4 13 3 12 7 9 12 4 13 3 12 2
2 0 9
18 0 9 4 10 9 1 3 9 7 13 1 9 15 10 9 0 13 2
7 9 9 13 1 0 9 2
5 0 9 4 0 2
32 15 13 16 9 13 16 9 1 9 13 1 3 7 10 0 9 2 3 12 9 1 10 0 9 7 12 9 1 12 9 3 2
14 3 9 2 3 1 9 2 1 0 9 4 13 9 2
15 9 13 16 9 1 9 13 12 9 7 3 13 0 9 2
17 15 13 3 16 9 4 0 1 12 9 1 16 9 4 4 13 2
23 1 9 4 3 9 13 3 16 9 3 13 12 9 7 9 4 0 0 9 7 12 9 2
20 9 4 3 13 1 3 0 9 16 9 3 13 3 0 9 7 12 0 9 2
16 9 2 15 4 0 1 10 9 7 0 9 2 13 1 9 2
24 9 13 1 9 2 15 13 0 7 9 9 3 12 9 1 9 7 15 13 9 1 0 9 2
22 9 13 1 10 9 1 3 12 9 1 9 2 1 9 12 12 9 1 9 0 2 2
11 16 9 4 10 0 9 13 3 3 9 2
25 9 13 1 0 9 9 2 16 9 3 4 13 15 0 7 1 0 9 3 13 9 1 0 9 2
10 9 4 4 13 16 9 13 12 9 2
16 15 15 4 0 13 3 9 1 9 16 9 13 1 12 9 2
19 9 13 12 9 1 9 2 1 9 12 4 15 12 9 1 9 0 2 2
21 1 9 7 9 7 9 7 9 4 15 13 1 0 9 15 13 14 13 1 9 2
6 15 13 1 10 9 2
14 2 9 2 13 1 2 0 9 2 7 2 9 2 2
10 3 13 15 1 2 10 0 9 2 2
25 7 15 4 0 14 13 16 10 0 9 4 0 3 1 10 9 16 0 9 1 9 13 1 9 2
22 1 3 10 9 13 15 1 9 0 9 7 9 2 9 2 9 2 9 2 9 3 2
27 7 7 13 15 3 3 13 10 9 15 13 2 7 3 13 15 1 10 9 15 3 13 9 1 9 3 2
21 10 0 9 1 10 9 4 16 9 2 9 2 1 9 7 9 13 10 0 9 2
27 3 13 12 9 7 9 2 9 1 10 9 4 3 4 9 2 1 11 4 9 2 9 3 12 9 2 2
20 0 9 0 1 9 4 9 2 9 2 3 9 1 13 7 9 2 0 9 2
29 15 4 3 13 10 9 9 1 0 9 7 9 9 2 9 2 9 2 9 2 9 2 9 2 9 3 1 9 2
14 10 9 1 14 13 13 10 9 9 7 9 4 0 2
20 1 9 2 3 2 13 3 0 9 7 3 3 0 10 9 15 13 1 9 2
16 9 13 3 15 1 9 1 9 2 1 9 1 10 0 9 2
9 9 13 0 0 9 1 10 9 2
19 7 10 0 9 4 3 0 3 15 4 13 15 10 9 1 0 9 9 2
29 10 9 2 3 1 11 13 9 10 9 1 10 9 2 15 4 3 3 0 7 10 0 9 1 0 11 7 11 2
3 9 4 0
10 1 10 9 4 9 3 13 15 0 2
13 9 3 1 0 2 9 2 13 1 10 0 9 2
19 7 10 9 2 3 12 9 1 9 9 13 2 13 15 3 3 1 15 2
12 11 13 3 10 9 2 9 7 9 7 11 2
9 11 13 1 3 0 9 7 11 2
10 10 9 9 4 0 2 0 3 0 2
10 0 7 0 9 13 1 9 1 9 2
16 15 13 3 12 9 2 15 13 15 1 10 0 7 0 9 2
9 9 1 10 9 4 4 3 0 2
14 1 9 3 0 0 9 2 11 2 13 0 0 9 2
11 1 9 7 11 13 10 9 1 0 9 2
29 9 1 11 9 11 4 13 3 0 14 13 15 3 1 0 9 1 10 0 9 7 10 9 14 13 15 1 9 2
9 1 11 13 12 0 9 7 9 2
21 15 1 10 9 2 15 1 9 13 0 2 13 10 9 3 0 7 3 10 0 2
25 1 12 9 3 13 15 9 1 11 2 1 11 7 1 11 2 12 9 16 9 13 13 1 11 2
11 10 0 9 4 13 3 1 12 1 11 2
15 1 11 2 11 7 11 13 1 9 9 3 3 0 9 2
6 10 0 9 4 4 0
38 3 9 9 13 1 9 4 11 7 11 9 1 9 0 1 10 0 9 2 1 14 13 10 0 9 2 15 13 11 2 11 2 11 2 11 7 11 2
23 15 15 3 13 2 10 9 9 0 9 2 4 13 7 15 1 10 3 0 9 1 9 2
15 14 13 10 9 13 14 13 15 7 13 15 1 0 9 2
33 12 7 9 9 1 11 2 11 2 11 2 11 3 13 10 0 9 1 9 1 9 2 9 2 9 2 9 2 9 2 9 2 2
6 9 13 1 10 9 2
17 15 4 3 13 7 9 2 9 3 13 3 1 7 9 1 9 2
19 1 0 9 4 15 13 1 16 9 1 10 0 9 13 9 1 9 9 2
18 10 0 9 4 3 10 0 9 1 16 15 13 9 13 3 1 9 2
13 3 13 10 0 9 9 1 10 9 3 1 11 2
41 1 3 9 13 10 9 1 0 9 2 15 1 0 9 3 13 2 9 2 2 9 2 2 13 0 9 2 15 15 4 13 9 1 2 9 4 4 13 10 9 2
17 9 2 7 9 7 9 2 13 3 3 1 0 9 3 1 9 2
15 9 9 2 1 9 12 9 2 1 12 9 3 3 0 2
31 1 15 15 4 13 4 11 10 3 0 2 7 3 15 13 9 7 9 10 3 0 2 9 1 1 9 12 9 1 9 2
9 3 13 11 1 12 9 1 9 2
21 9 0 9 13 3 1 12 9 9 1 9 2 7 9 4 0 3 9 4 0 2
20 3 4 15 3 12 9 2 1 9 9 12 9 16 10 0 9 1 9 13 2
5 9 4 3 0 2
9 10 0 9 4 3 13 1 9 2
8 7 9 4 0 1 9 9 2
30 15 4 9 1 16 0 9 3 13 1 0 9 2 16 9 9 1 9 4 13 7 16 9 1 9 7 9 4 13 2
29 9 4 13 3 3 2 15 13 3 3 16 10 9 13 0 9 7 3 2 7 15 15 13 13 1 3 0 9 2
20 1 9 13 9 10 0 9 2 3 3 3 3 10 0 9 13 10 0 9 2
20 1 0 9 4 9 3 0 2 16 9 3 12 9 13 1 9 1 0 9 2
18 14 13 9 2 13 9 7 13 9 1 10 9 4 1 0 9 0 2
24 10 3 0 9 9 1 0 9 13 9 7 9 1 10 9 2 3 15 3 13 9 7 9 2
9 10 0 1 9 13 15 1 9 2
33 3 15 3 3 3 4 13 9 13 10 9 2 15 1 10 9 2 9 2 9 2 9 7 9 4 10 0 7 0 9 1 9 2
4 9 9 13 2
6 7 15 13 3 9 2
16 3 1 10 0 9 1 9 13 15 3 0 1 15 7 15 2
6 3 4 9 13 3 2
10 3 4 15 13 10 0 9 1 9 2
13 15 4 3 13 16 9 4 0 3 9 4 0 2
15 0 9 13 15 15 3 3 15 13 10 9 1 10 9 2
3 9 7 9
16 0 0 9 7 9 2 9 7 9 13 3 3 1 0 9 2
16 3 13 3 12 9 9 4 0 1 9 2 12 9 1 9 2
8 3 12 9 13 1 9 9 2
18 0 9 1 9 13 0 9 1 11 2 11 7 11 7 13 3 9 2
29 9 13 2 1 10 9 15 13 2 1 11 4 12 9 3 0 7 1 11 2 1 11 7 11 12 9 3 0 2
27 1 16 9 0 9 13 3 4 9 1 9 1 9 3 0 7 3 2 3 7 1 10 9 3 3 0 2
20 1 10 9 13 9 1 9 7 3 1 9 7 1 10 0 9 2 9 2 2
24 1 11 7 0 9 2 3 10 0 13 1 0 9 2 13 15 3 7 15 15 13 1 15 2
22 4 9 13 7 10 0 9 13 2 4 9 1 0 9 1 9 13 3 1 9 12 2
26 10 9 9 13 1 16 9 1 9 1 9 4 13 9 1 9 2 15 1 0 9 13 9 7 9 2
17 9 1 9 4 0 13 3 1 10 3 9 1 10 0 9 11 2
21 15 4 13 9 1 9 2 9 2 1 9 1 10 9 2 11 2 11 9 2 2
28 3 13 15 3 0 9 2 9 7 9 2 4 13 2 7 13 3 3 0 15 4 16 9 13 3 0 9 2
11 3 3 4 15 13 1 10 9 1 9 2
21 1 9 13 3 9 1 3 9 7 9 2 9 2 9 2 9 7 0 0 9 2
1 9
14 3 15 4 13 15 4 15 13 1 9 3 15 13 2
19 1 9 4 15 13 2 16 9 13 1 9 2 9 2 16 15 3 13 2
14 3 13 15 3 9 1 3 0 7 0 9 13 1 2
15 15 15 4 3 12 9 4 13 9 9 1 14 13 15 2
14 4 15 7 15 3 12 9 13 3 0 9 1 9 2
19 3 15 4 13 15 13 15 16 0 9 13 0 0 7 0 9 1 15 2
8 9 13 3 9 14 13 15 2
4 3 13 9 2
19 15 13 3 16 10 9 1 9 9 13 9 1 9 1 10 0 9 9 2
20 15 4 3 13 1 16 0 9 15 3 4 4 13 1 9 4 4 0 9 2
6 10 0 9 13 9 2
10 9 4 13 1 9 1 14 13 0 2
7 9 13 9 1 10 9 2
9 15 13 3 9 7 9 1 9 2
18 15 13 9 3 1 0 9 7 15 4 0 14 13 9 9 7 9 2
13 13 9 9 12 2 9 9 12 7 9 9 12 2
6 15 13 15 1 9 2
1 9
1 9
16 16 10 9 13 4 1 9 9 3 4 13 1 16 9 13 2
5 10 9 13 9 2
10 15 4 13 1 9 1 0 9 3 2
19 3 4 3 0 9 13 7 16 15 4 3 1 14 3 13 14 13 3 2
18 16 3 10 0 9 4 13 9 4 15 7 15 13 10 0 1 9 2
22 16 15 13 9 4 15 0 14 13 9 1 9 7 1 9 2 15 4 0 1 9 2
10 9 13 1 1 14 13 9 10 9 2
24 16 15 4 13 9 1 3 1 9 2 15 15 4 13 2 13 9 7 1 9 1 0 9 2
1 9
26 16 9 4 13 15 1 15 2 0 2 1 3 12 9 2 4 15 7 15 13 16 9 13 1 9 2
6 15 13 16 9 13 2
15 3 1 9 1 9 4 9 13 1 0 9 1 0 9 2
18 7 1 9 7 9 4 9 13 15 1 9 15 4 13 9 1 9 2
15 16 15 1 9 13 4 0 14 13 9 4 0 9 13 2
18 9 13 3 16 15 4 13 9 2 3 9 4 13 7 1 0 9 2
10 13 3 9 9 12 7 9 9 12 2
16 15 13 15 1 9 2 9 2 9 7 9 2 9 7 9 2
19 14 13 10 9 4 10 0 9 7 9 7 13 10 0 9 1 10 9 2
14 10 0 9 13 15 3 3 3 0 16 15 4 13 2
19 7 14 4 0 7 0 1 9 4 0 7 0 7 13 1 16 9 13 2
25 10 0 9 1 9 13 13 3 3 3 15 4 13 1 10 9 10 9 7 13 15 0 7 0 2
19 16 9 4 0 7 0 10 9 1 9 2 13 10 0 9 3 1 15 2
22 4 15 0 4 10 0 9 7 10 0 9 3 4 15 7 3 3 9 1 0 9 2
18 3 4 3 9 15 15 4 3 1 9 14 13 7 9 7 9 1 2
16 9 13 3 13 10 0 9 1 14 13 1 1 14 13 15 2
12 16 0 9 1 9 13 9 3 13 9 9 2
3 9 7 9
21 10 9 13 1 3 15 4 13 1 10 9 1 9 7 10 9 15 13 1 15 2
9 10 9 4 13 9 1 0 9 2
20 9 13 3 3 1 3 9 13 3 2 7 3 1 15 7 3 9 7 9 2
29 3 9 4 14 13 7 9 2 10 9 15 4 14 13 7 3 9 13 13 3 1 0 9 1 10 9 15 13 2
20 1 15 9 13 9 10 0 9 1 9 7 9 2 7 3 1 9 7 9 2
32 15 4 0 14 13 2 16 9 15 13 15 0 1 10 0 13 3 0 7 0 1 15 7 15 15 3 13 9 7 0 9 2
32 3 13 15 10 9 1 9 15 9 13 3 1 2 3 10 0 9 15 3 7 3 13 15 15 1 14 4 3 13 10 9 2
11 9 13 0 9 7 0 9 1 14 13 2
31 15 4 0 16 10 0 9 1 9 7 9 4 13 3 1 15 15 13 15 2 3 16 15 1 9 13 15 0 7 0 2
23 10 9 15 13 9 13 15 3 0 7 13 16 15 3 4 13 10 9 15 15 4 13 2
27 7 2 3 16 9 15 4 4 3 1 9 4 0 2 4 15 13 15 15 15 13 1 0 7 0 9 2
20 3 4 10 0 9 1 9 13 2 7 9 3 1 10 0 4 3 3 0 2
28 9 4 3 13 2 16 9 13 15 0 1 9 2 7 15 13 1 9 2 1 10 9 7 15 13 15 3 2
23 15 4 0 16 9 4 13 10 9 2 3 4 13 9 1 10 0 9 7 13 1 9 2
9 13 3 9 0 3 10 0 9 2
24 15 4 3 3 0 7 4 3 13 15 0 16 15 3 4 13 13 7 13 13 15 1 9 2
14 9 4 3 0 7 4 3 13 1 9 1 10 0 2
27 4 9 13 1 9 2 9 7 1 0 9 13 3 2 4 15 0 2 16 9 13 15 3 3 7 0 2
1 9
16 9 9 13 1 10 0 9 2 1 3 0 3 1 10 9 2
18 10 9 9 4 0 7 15 0 2 9 13 13 3 15 1 0 9 2
28 15 4 13 2 16 10 9 4 0 1 10 9 2 3 3 15 13 14 13 2 7 0 1 14 13 7 3 2
11 15 13 3 9 1 14 13 1 10 9 2
8 10 9 13 1 10 0 9 2
16 1 10 0 9 13 15 0 9 10 9 2 3 13 15 3 2
12 0 9 13 1 3 0 2 0 4 9 9 2
23 1 10 0 9 13 9 3 1 9 2 9 13 9 7 15 4 3 13 3 10 0 9 2
19 15 4 3 13 9 7 16 9 13 1 9 3 4 15 14 13 15 1 2
12 3 1 12 9 9 13 15 15 14 13 3 2
27 3 3 4 9 13 3 9 7 9 3 15 13 1 9 7 15 13 1 14 13 3 7 13 1 10 9 2
11 15 13 9 7 13 15 13 1 1 9 2
18 15 4 13 15 3 1 9 2 3 16 15 3 13 3 7 13 15 2
15 9 13 3 3 1 9 1 9 0 1 10 9 1 9 2
22 15 13 13 1 9 7 3 13 9 3 1 10 0 9 2 3 10 9 7 10 9 2
20 1 9 13 9 4 13 1 9 2 7 13 0 13 15 3 1 1 12 9 2
16 15 13 1 10 9 15 13 1 10 9 7 13 15 1 9 2
6 15 13 3 0 9 2
12 0 9 7 0 0 9 4 4 0 7 0 2
13 1 0 9 13 10 0 9 13 15 3 7 13 2
9 10 9 13 7 13 3 1 9 2
25 15 13 15 15 13 3 7 3 13 10 9 3 15 4 13 3 15 15 4 13 3 7 13 15 2
22 7 0 9 13 3 3 4 15 13 1 14 3 1 9 13 15 1 10 9 7 9 2
22 1 9 13 10 9 9 13 10 0 9 2 7 10 0 13 3 13 3 10 9 3 2
12 10 0 0 9 13 13 15 1 12 9 9 2
11 1 10 9 13 9 3 1 9 7 9 2
16 3 1 9 1 9 4 15 0 16 15 13 7 13 1 9 2
22 9 13 1 10 0 9 2 3 13 0 9 2 9 2 3 9 3 13 1 0 9 2
14 1 9 13 10 0 0 9 13 2 15 3 13 9 2
21 14 13 1 3 9 13 2 13 3 15 13 7 13 15 0 9 4 10 0 9 2
31 15 13 3 15 15 13 1 9 0 9 2 3 15 13 1 10 3 0 9 1 10 0 9 0 14 13 10 9 1 9 2
1 9
18 9 4 10 0 2 7 7 9 3 10 0 2 7 1 9 7 9 2
7 9 13 15 15 9 13 2
15 9 13 3 9 7 9 10 3 0 9 1 9 7 9 2
25 7 2 16 9 13 0 1 9 7 3 3 15 3 2 4 15 13 9 10 0 9 1 10 9 2
24 9 13 15 3 1 10 0 0 9 7 15 13 3 0 9 2 15 13 10 0 9 1 9 2
7 9 13 3 9 1 9 2
12 15 4 0 16 9 13 3 0 9 7 0 2
22 15 4 3 0 16 9 13 1 9 9 1 9 2 3 16 15 4 13 10 0 9 2
58 15 4 3 3 0 14 13 9 1 15 16 15 13 0 9 1 9 2 15 3 3 13 15 0 1 10 0 15 4 13 9 3 1 15 0 2 7 16 9 4 13 7 10 0 9 1 9 7 9 4 15 0 1 7 9 7 9 2
7 13 9 3 1 9 9 2
18 10 0 9 4 14 3 13 10 9 13 7 13 1 9 10 0 9 2
19 15 4 3 3 13 15 1 9 2 7 4 13 16 15 13 1 15 0 2
14 10 0 9 13 3 15 1 3 0 9 1 10 9 2
16 9 4 3 10 9 13 10 0 9 7 4 3 3 13 15 2
28 15 13 0 9 7 0 9 1 14 13 15 15 1 9 7 15 13 3 13 3 16 15 13 1 1 15 0 2
1 9
21 10 0 9 13 3 14 13 7 15 4 3 13 15 1 14 13 15 0 7 0 2
21 1 15 13 15 1 9 7 9 2 15 13 3 10 9 7 13 3 3 10 9 2
26 13 9 9 4 15 13 1 2 16 15 4 0 7 1 10 0 9 2 15 3 4 13 3 1 9 2
18 2 9 2 13 0 9 3 3 1 14 4 13 1 7 13 1 9 2
1 9
23 15 4 0 16 9 13 3 2 7 16 15 3 13 1 9 4 15 15 14 13 15 1 2
19 13 15 3 13 3 10 9 2 16 15 0 9 4 4 0 14 13 1 2
8 9 4 3 4 0 7 0 2
9 15 4 4 3 0 7 3 0 2
9 9 4 13 3 7 9 4 0 2
17 15 3 13 0 2 13 0 1 9 7 13 1 0 9 7 9 2
22 10 3 0 9 4 16 9 13 15 0 7 13 9 1 14 13 3 1 9 10 9 2
14 14 13 9 3 15 4 0 13 3 14 13 3 15 2
14 0 0 9 13 15 3 0 1 9 1 10 0 9 2
8 7 3 13 9 10 0 9 2
21 13 13 0 9 1 9 2 13 7 13 1 9 7 13 1 14 4 3 1 15 2
11 9 7 9 4 9 3 13 3 3 1 2
6 9 9 13 1 9 2
14 15 4 3 13 3 7 12 9 16 15 13 3 3 2
13 15 13 3 1 9 2 16 15 4 10 0 9 2
13 9 1 10 9 13 3 3 9 3 15 13 15 2
7 9 13 3 3 7 3 2
11 1 9 13 15 3 10 9 9 1 9 2
8 3 3 12 13 10 0 9 2
5 3 13 9 13 2
12 12 2 3 12 9 3 2 4 15 12 9 2
12 12 2 3 12 9 3 2 4 15 12 9 2
12 12 2 3 12 9 3 2 4 15 12 9 2
10 9 12 7 3 3 4 15 12 9 2
17 7 15 13 1 9 16 9 3 4 13 10 0 9 3 1 9 2
9 3 1 12 9 4 9 3 0 2
11 10 9 1 1 9 4 14 13 7 0 2
12 12 9 9 1 9 4 13 0 9 1 9 2
12 4 13 9 9 3 3 16 3 10 9 13 2
6 15 13 3 3 9 2
25 9 9 4 0 1 9 15 13 0 9 7 1 10 9 15 13 9 10 9 15 9 7 9 13 2
9 15 13 0 10 9 15 13 9 2
3 13 9 2
9 13 15 15 15 13 15 1 9 2
23 15 4 3 13 10 9 2 7 15 0 13 16 10 9 3 4 0 12 9 16 9 13 2
9 7 3 9 11 11 4 13 15 2
14 2 4 15 13 9 1 10 9 16 15 13 15 2 2
32 10 0 9 11 11 11 4 1 2 9 2 2 11 2 9 12 2 13 10 10 0 9 9 1 10 0 9 1 9 7 9 2
18 15 13 15 0 1 9 2 7 3 14 13 13 10 10 9 4 0 2
5 15 4 9 3 2
14 15 13 16 15 4 0 1 12 9 2 16 3 3 2
56 3 3 16 9 13 3 3 2 7 15 13 16 1 10 9 4 9 9 3 0 1 9 1 9 1 0 9 2 0 9 7 9 1 0 9 16 15 13 1 10 0 9 15 13 10 0 9 1 9 9 1 3 3 12 9 2
39 16 9 1 0 9 9 13 9 9 13 13 9 2 13 9 3 9 16 15 4 13 7 13 3 10 9 2 3 13 3 10 9 15 3 4 0 14 13 2
56 15 4 13 9 1 9 1 9 2 13 1 9 7 9 1 9 2 10 9 3 15 3 4 13 10 9 1 10 9 1 9 1 9 2 10 9 1 9 7 9 2 1 0 9 7 0 9 2 10 9 3 9 13 7 9 2
1 0
71 3 10 0 9 13 13 1 10 9 3 15 4 13 3 3 7 3 1 0 9 2 13 3 1 9 9 13 9 2 4 13 1 9 2 13 10 10 9 1 9 2 13 10 9 2 0 1 9 7 13 1 0 9 1 9 2 3 13 15 3 7 9 2 7 15 4 3 3 3 0 2
29 10 0 15 4 13 1 9 13 16 9 4 13 1 10 0 9 7 16 9 1 0 7 0 3 13 0 7 0 2
11 15 4 0 16 11 13 3 1 10 9 2
25 7 9 1 0 11 2 15 13 12 9 1 9 9 2 13 3 3 9 1 9 1 9 10 9 2
24 16 10 9 9 4 13 3 7 3 1 11 0 9 2 4 15 3 13 1 10 0 9 9 2
3 13 3 3
20 3 13 9 1 11 1 14 12 7 13 10 0 9 7 3 13 15 1 9 2
6 15 13 3 3 3 2
5 15 4 0 9 2
20 9 1 9 7 9 4 3 14 13 0 7 0 10 9 15 13 3 1 9 2
6 9 13 0 7 0 2
15 9 13 1 10 9 1 10 9 3 9 3 3 4 13 2
6 11 13 11 7 9 2
20 15 13 1 9 16 9 9 4 0 1 12 9 1 9 7 12 9 1 9 2
6 1 9 13 15 3 2
12 9 1 9 13 3 2 0 3 1 9 9 2
15 9 13 0 7 13 15 1 9 1 14 13 9 1 9 2
1 3
15 11 13 3 10 9 1 12 9 7 10 9 1 12 9 2
14 11 9 13 1 10 9 1 9 7 13 10 0 9 2
21 9 12 13 9 13 10 9 1 12 9 1 12 9 1 9 7 12 9 1 9 2
13 9 4 3 13 1 12 1 12 9 1 12 9 2
25 3 4 15 13 9 1 9 2 9 7 0 0 9 1 10 9 15 3 13 15 1 9 1 9 2
28 3 1 14 13 10 9 1 10 0 9 13 15 12 0 9 1 9 2 0 16 15 3 3 13 3 1 9 2
2 0 9
13 10 0 9 4 11 2 13 13 10 0 1 15 2
10 9 9 13 1 9 1 12 1 9 2
14 15 13 16 9 1 9 13 1 12 7 12 9 9 2
14 9 13 3 3 1 16 15 13 9 2 0 1 9 2
7 12 9 13 1 10 9 2
22 9 13 1 0 9 1 9 2 7 3 15 13 9 13 9 7 9 3 3 7 3 2
11 9 13 7 9 7 15 0 1 0 9 2
35 9 7 11 4 3 13 15 7 9 2 3 9 3 4 13 2 9 13 0 9 7 9 13 7 13 1 9 1 16 15 13 15 1 15 2
31 9 1 10 2 0 2 9 4 1 3 10 9 1 11 2 11 7 11 2 7 15 13 14 13 3 15 1 10 0 9 2
20 11 11 1 11 13 12 9 12 2 13 12 9 3 7 3 12 9 9 12 2
26 7 15 4 9 15 3 13 1 9 2 7 1 9 2 1 0 9 7 1 9 2 0 1 12 9 2
1 9
29 15 4 1 9 13 3 1 9 0 9 1 9 2 3 16 15 3 15 13 3 4 9 1 9 0 9 3 3 2
25 10 10 0 2 9 1 9 1 9 7 9 7 9 2 9 7 10 0 9 2 4 9 1 9 2
29 11 13 1 0 9 3 9 13 3 10 3 0 9 2 3 13 3 9 1 9 3 16 9 13 13 15 1 9 2
36 15 13 3 7 0 7 0 9 1 3 0 9 4 13 10 2 0 9 2 1 0 9 7 3 15 3 1 0 0 9 13 15 0 9 3 2
1 9
36 16 15 4 13 15 16 10 0 9 4 0 1 9 2 3 4 11 0 1 16 9 2 10 0 9 2 4 0 14 13 15 1 3 1 9 2
5 15 4 13 9 2
14 16 15 3 4 13 15 3 12 9 1 9 1 9 2
17 7 15 13 10 0 9 15 13 13 3 9 9 13 1 3 3 2
29 2 15 13 10 0 9 1 10 0 9 14 13 10 0 9 1 9 3 3 3 16 10 0 9 4 3 0 2 2
9 9 4 13 15 1 14 13 9 2
19 15 13 3 12 9 11 1 9 2 15 4 3 7 0 0 9 1 11 2
10 9 13 3 3 1 12 9 1 9 2
11 9 13 9 3 1 12 9 11 1 9 2
4 9 9 1 9
17 1 9 13 12 1 12 1 9 9 12 1 11 2 0 2 9 2
9 7 3 0 13 9 3 1 9 2
6 9 9 1 3 12 9
20 1 12 9 13 15 3 12 9 2 3 9 15 13 3 7 12 9 9 0 2
5 15 1 11 9 2
7 2 15 13 9 1 9 2
7 10 0 9 4 4 0 2
9 9 7 0 9 4 4 3 0 2
15 10 0 9 4 13 0 1 15 1 9 1 10 9 2 2
11 2 9 1 10 0 9 2 9 12 2 2
22 11 4 13 10 9 1 2 0 9 2 2 10 9 14 13 1 0 9 1 9 9 2
8 1 9 13 15 1 11 9 2
17 9 13 10 9 15 4 13 3 9 13 1 9 1 9 1 9 2
27 9 13 3 1 11 9 2 11 12 2 9 12 2 12 2 7 0 9 7 9 9 2 9 7 9 2 2
17 1 10 9 15 15 13 14 13 10 3 9 13 12 9 1 9 2
7 1 10 9 13 12 9 2
8 9 9 4 13 1 12 9 2
14 3 3 15 13 3 4 15 13 13 1 3 12 9 2
29 10 12 15 13 10 9 4 13 16 15 4 13 10 9 1 9 2 7 16 9 0 7 0 9 4 4 13 15 2
6 3 4 9 3 0 2
19 10 9 15 13 3 9 1 10 0 2 0 9 2 12 13 3 10 9 2
11 9 4 13 10 9 1 14 13 1 3 2
9 9 13 14 13 0 9 7 9 2
4 3 13 9 2
5 1 9 10 9 2
17 3 0 13 3 1 9 2 7 10 0 9 1 9 4 13 9 2
13 15 4 9 7 11 2 11 2 11 7 11 13 2
1 13
20 9 1 9 4 3 0 16 9 9 15 7 4 13 7 13 2 9 2 13 2
11 3 4 15 3 3 13 1 9 1 9 2
11 1 9 13 15 12 9 0 9 1 9 2
16 3 13 15 15 1 9 15 13 9 1 10 9 9 0 9 2
9 3 13 15 3 15 15 13 15 2
7 10 9 13 3 1 9 2
16 3 3 15 13 16 10 0 9 4 9 3 4 15 10 9 2
11 9 4 9 1 10 0 0 1 9 9 2
11 9 13 3 7 3 13 1 9 1 9 2
1 0
48 3 10 2 0 2 2 9 13 4 15 13 2 9 13 3 1 2 15 13 3 0 9 7 9 2 3 13 9 0 7 15 13 1 9 7 13 3 2 16 15 3 13 9 14 13 1 9 2
10 10 0 9 4 16 9 13 0 9 2
17 15 13 1 16 9 13 1 10 0 9 7 3 13 9 1 9 2
8 9 4 3 0 1 9 9 2
7 15 4 3 0 7 0 2
15 15 13 3 3 10 0 9 15 13 1 14 13 9 3 2
14 9 13 9 9 16 9 7 0 9 3 4 3 0 2
5 15 13 1 9 2
6 15 13 7 13 9 2
9 10 9 4 3 3 0 14 13 2
28 15 13 14 13 9 3 3 0 2 3 0 1 9 9 2 3 16 15 4 9 1 0 9 7 9 1 9 2
9 0 9 4 11 7 11 3 13 2
15 7 10 0 9 2 9 7 9 1 9 2 4 3 0 2
14 0 9 2 6 2 7 15 4 3 15 14 13 1 2
11 10 9 9 4 3 14 13 9 1 9 2
14 10 0 9 13 9 16 10 9 4 4 13 1 9 2
17 7 1 0 9 13 15 1 9 16 10 0 9 13 10 0 9 2
1 15
15 11 13 3 10 0 9 14 3 13 10 9 13 1 9 2
17 3 13 15 15 13 1 9 0 9 2 10 9 15 4 0 15 2
16 0 9 15 13 0 7 3 0 9 4 11 2 11 7 11 2
12 0 9 1 11 4 3 13 9 1 0 9 2
16 1 11 2 11 7 11 4 10 0 9 3 13 13 10 9 2
14 14 13 9 1 9 2 10 0 9 2 3 10 9 2
4 10 9 0 9
25 12 9 1 9 2 15 4 15 15 3 13 1 9 1 10 9 15 4 13 15 14 13 7 13 2
15 3 3 1 9 13 15 12 9 1 14 13 10 0 13 2
24 9 13 3 12 9 3 1 9 7 1 9 2 12 9 9 1 9 1 9 2 12 1 9 2
30 9 2 11 2 11 2 11 3 2 13 10 3 0 9 1 10 9 1 9 2 12 9 2 7 9 2 12 9 2 2
15 9 13 12 9 1 9 7 9 1 9 2 9 12 9 2
16 9 13 12 9 1 9 9 2 7 3 12 9 1 9 9 2
14 9 9 4 3 3 0 7 10 9 1 9 1 9 2
13 3 10 0 9 4 9 2 4 7 13 7 13 2
6 9 9 13 10 9 2
6 9 13 3 7 9 2
14 1 9 1 9 12 9 1 11 13 12 1 9 12 2
5 15 4 12 9 2
11 12 13 12 1 9 1 10 9 1 9 2
7 15 4 3 3 12 9 2
11 3 9 1 15 1 9 4 3 12 9 2
8 0 9 1 9 4 12 9 2
16 15 13 16 9 2 15 13 3 9 2 4 13 3 1 9 2
16 1 0 9 1 11 7 11 13 3 7 10 9 1 12 9 2
6 9 4 0 1 9 2
24 1 10 9 15 13 3 9 1 9 13 15 3 10 0 9 15 3 13 3 12 7 0 9 2
9 15 13 1 0 9 2 0 9 2
16 9 9 1 9 13 3 7 9 9 2 12 9 1 12 9 2
35 15 4 13 3 16 16 9 4 13 10 9 14 13 3 0 12 2 3 13 12 9 9 7 9 2 12 9 0 7 15 15 13 1 9 2
15 3 12 9 1 9 1 11 7 11 4 9 2 12 2 2
17 9 3 13 3 3 9 13 1 9 9 9 1 9 1 0 9 2
15 0 9 13 3 12 9 9 2 16 9 3 13 12 9 2
11 9 1 11 4 13 1 3 9 1 9 2
25 1 9 13 9 7 9 16 9 1 9 13 0 9 2 9 2 9 7 9 4 3 0 14 13 2
7 15 4 10 9 1 9 2
8 3 13 1 9 9 7 9 2
21 7 9 1 10 0 9 4 10 9 15 13 3 0 9 1 9 7 9 1 9 2
15 3 4 9 0 0 2 7 10 9 1 9 4 15 3 2
34 2 9 1 9 1 1 15 9 4 13 1 3 9 1 9 1 0 9 1 11 2 13 9 11 11 11 2 9 1 9 9 1 11 2
29 2 3 13 15 16 9 1 11 4 0 7 3 3 3 13 15 9 1 16 7 9 2 9 7 9 4 3 0 2
20 9 1 9 1 10 3 9 13 1 10 0 9 15 13 1 10 9 1 11 2
2 0 9
17 1 9 4 15 13 0 9 1 10 9 9 1 7 11 7 11 2
17 9 1 10 9 13 16 0 11 13 1 0 0 9 9 7 9 2
23 2 9 4 13 0 7 3 3 3 4 15 10 9 2 13 7 9 9 1 9 7 9 2
19 7 10 9 7 9 1 15 4 3 13 1 9 1 9 3 0 0 9 2
20 9 1 9 13 1 3 1 9 1 10 9 1 14 13 9 1 9 1 9 2
10 2 3 13 15 3 12 9 3 9 2
7 7 10 9 4 3 0 2
18 10 0 3 9 13 15 3 0 2 13 9 11 11 1 0 9 9 2
2 0 9
24 2 3 4 15 0 16 0 9 3 13 9 1 16 9 3 4 0 7 9 2 13 11 11 2
13 2 15 4 3 0 1 16 11 13 0 9 9 2
7 7 15 4 10 0 9 2
14 2 7 9 0 9 13 3 1 9 1 10 3 9 2
13 15 13 16 9 1 9 13 3 1 10 3 9 2
17 2 10 0 9 4 15 3 13 1 9 11 11 2 13 11 11 2
15 12 9 1 12 13 0 7 3 12 1 12 4 3 0 2
11 10 0 0 9 13 0 0 9 1 9 2
16 3 0 4 15 1 0 0 9 1 9 1 9 12 0 9 2
27 15 4 15 1 10 10 9 15 0 9 11 11 1 0 9 1 11 13 3 1 10 9 1 12 0 9 2
8 1 9 13 11 11 1 9 2
25 10 12 9 4 13 1 12 9 2 1 0 9 1 9 2 3 1 9 7 12 9 1 9 9 2
12 1 10 0 7 0 9 13 3 9 11 11 2
6 0 9 4 2 0 2
14 0 0 0 9 13 0 1 10 9 2 13 11 11 2
15 10 0 9 2 0 9 7 0 9 13 1 10 0 9 2
27 3 13 15 1 9 10 0 9 9 2 3 12 9 2 15 1 9 13 0 9 15 1 0 9 13 9 2
14 1 10 9 13 12 9 9 15 13 1 0 0 9 2
22 2 3 13 3 16 15 13 1 9 1 9 15 13 10 0 0 9 2 13 11 11 2
15 7 1 10 9 4 0 9 3 0 1 9 7 1 9 2
22 0 9 1 9 7 1 0 9 1 9 4 13 9 1 7 1 10 9 2 13 9 2
16 10 0 9 7 0 9 4 1 10 9 9 13 1 0 9 2
21 10 0 9 1 9 1 9 13 3 1 10 9 15 4 13 0 9 1 10 9 2
5 0 9 13 0 9
19 9 9 1 10 0 9 13 3 1 0 9 1 16 9 4 0 7 3 2
18 0 7 10 9 13 1 1 9 1 15 1 10 9 15 13 0 9 2
13 12 9 1 9 1 9 11 9 4 0 1 9 2
9 10 9 4 10 9 2 13 15 2
8 15 13 1 0 9 0 3 2
9 15 4 2 13 14 13 15 2 2
8 10 9 1 9 13 3 0 2
10 10 0 9 1 9 13 3 1 9 2
34 9 15 3 4 13 9 1 0 9 2 15 3 4 13 15 1 10 0 9 7 13 10 3 0 9 1 9 13 3 9 1 10 9 2
23 10 9 9 15 13 16 15 13 9 2 15 13 9 1 9 2 4 3 13 9 1 9 2
17 9 1 9 4 4 10 9 1 10 9 1 9 2 13 11 11 2
17 10 3 0 9 1 9 4 13 10 0 9 3 3 9 4 0 2
2 0 9
21 15 13 3 1 14 13 9 1 9 3 7 10 9 4 13 3 1 10 0 9 2
19 15 4 13 16 15 3 4 13 0 9 7 10 0 9 2 13 11 11 2
18 3 13 9 7 16 9 4 0 7 3 10 0 9 1 9 1 9 2
19 3 0 9 2 15 13 15 7 0 1 0 9 2 13 3 10 0 9 2
15 16 9 13 1 7 3 13 3 13 10 0 9 1 9 2
18 2 15 4 0 3 3 0 14 13 0 9 1 9 2 13 11 11 2
29 7 15 13 16 9 13 16 0 9 2 3 1 9 1 9 1 9 2 4 4 13 10 9 1 10 9 15 13 2
21 7 0 9 1 9 13 1 9 1 9 7 9 7 0 9 13 1 3 0 9 2
27 9 4 13 10 9 15 1 9 7 0 13 1 14 13 10 9 1 9 9 15 1 0 9 13 15 15 2
25 1 15 4 10 0 9 4 0 7 0 0 7 13 3 14 13 7 10 9 1 10 0 9 9 2
26 1 15 3 4 9 4 3 0 7 13 15 0 9 7 4 3 13 1 0 9 15 13 7 0 9 2
25 15 13 9 1 10 9 15 13 10 0 9 1 10 9 15 1 9 13 1 9 2 9 7 9 2
24 1 0 9 4 15 3 13 15 0 7 0 9 2 1 0 9 13 15 3 3 1 10 9 2
37 15 13 10 9 1 16 9 1 9 9 1 9 1 9 4 9 1 10 0 9 7 15 4 13 3 1 15 16 1 10 9 4 10 9 3 13 2
18 15 13 3 3 3 16 15 13 9 3 10 0 9 4 1 0 9 2
24 15 13 1 10 0 15 1 9 0 4 13 13 3 1 10 9 1 9 15 4 13 1 9 2
27 9 1 10 3 0 9 4 16 15 1 0 9 13 16 15 1 10 9 4 13 0 9 1 10 0 9 2
32 15 13 15 3 1 9 3 9 1 9 9 3 3 4 9 7 1 9 13 1 10 0 9 1 9 1 10 9 15 13 9 2
24 10 0 9 4 13 1 10 0 9 7 3 1 16 9 1 9 7 9 1 10 9 4 0 2
2 13 9
21 1 0 9 4 9 13 10 0 9 1 9 7 13 3 10 0 9 1 9 9 2
22 9 13 3 3 1 9 1 9 3 3 1 15 1 9 7 4 13 1 9 0 9 2
16 15 4 1 0 10 9 3 13 1 9 15 13 1 3 9 2
23 10 0 9 4 13 1 2 9 2 1 10 0 9 7 4 3 13 0 9 1 9 9 2
18 15 13 1 15 1 11 3 15 13 10 9 1 0 9 1 0 9 2
15 3 15 13 1 0 9 1 15 13 10 0 15 3 0 2
11 2 13 3 1 15 1 3 0 9 2 2
8 2 13 10 9 1 15 2 2
32 10 9 15 13 4 1 15 13 10 0 9 2 3 1 9 1 11 2 10 9 3 7 9 2 9 2 9 7 9 4 0 2
19 11 4 13 1 15 1 9 1 10 0 9 2 9 9 11 11 1 11 2
1 9
20 15 4 13 15 14 13 7 13 16 9 3 3 13 1 9 3 10 9 13 2
27 15 4 3 1 0 9 1 9 0 14 13 3 0 9 1 9 3 1 16 15 4 0 2 13 9 11 2
25 15 4 1 10 0 9 13 10 0 9 1 14 13 16 15 4 13 1 16 9 9 4 13 0 2
20 1 0 11 9 1 11 13 3 7 9 1 10 9 15 3 13 2 9 9 2
35 16 3 3 10 9 7 3 3 4 13 10 9 1 10 9 15 13 3 2 3 4 15 10 0 9 2 7 1 10 0 7 10 0 9 2
31 10 0 9 4 3 3 14 13 3 10 9 3 9 13 1 10 0 9 2 3 10 9 3 10 9 1 9 4 13 13 2
25 1 10 9 15 13 1 0 9 1 9 1 11 2 10 3 9 2 13 3 9 14 13 10 9 2
11 15 4 3 3 9 1 10 9 1 9 2
1 9
34 1 9 1 10 0 9 15 13 16 9 13 1 9 7 13 10 9 1 9 3 13 2 3 9 13 2 10 0 9 3 3 1 9 2
28 10 9 2 15 3 0 13 9 4 1 10 9 13 1 10 9 3 15 13 10 9 15 1 0 9 4 13 2
45 3 15 13 10 0 9 3 15 13 13 9 9 13 10 0 9 3 1 9 7 15 4 1 9 1 9 13 9 9 2 16 15 4 0 7 13 1 9 15 13 1 10 0 9 2
18 9 13 3 3 10 0 9 15 13 1 9 1 10 0 9 1 9 2
27 10 0 9 4 1 9 1 14 7 1 10 3 0 9 13 3 1 9 2 1 9 13 3 1 9 9 2
2 1 9
40 1 9 15 13 10 9 1 9 2 9 7 9 1 9 9 2 13 3 10 9 1 10 0 9 1 9 2 1 9 7 1 10 9 15 13 1 9 1 9 2
37 15 13 3 16 15 0 10 2 0 2 9 13 10 0 9 1 9 1 10 0 9 7 16 10 9 1 0 7 0 9 4 13 1 9 1 9 2
37 10 9 15 13 9 4 13 1 9 9 7 3 13 15 1 9 1 9 1 10 0 2 9 2 12 0 9 2 15 4 13 1 9 1 12 9 2
30 15 4 3 10 0 9 7 3 13 0 9 1 0 9 1 9 0 10 9 1 9 2 1 10 9 7 3 9 13 2
19 3 3 9 4 0 4 9 1 9 13 15 1 10 9 1 10 0 9 2
2 12 9
34 9 13 3 3 0 9 1 9 7 10 3 9 7 10 3 9 2 7 0 10 9 4 0 1 9 7 13 3 16 9 13 1 9 2
28 16 9 1 9 4 3 0 14 13 7 3 13 1 9 1 9 2 13 3 9 15 9 14 13 3 0 9 2
11 15 13 1 15 9 15 13 3 1 15 2
25 15 4 1 10 9 16 9 9 1 9 7 10 0 9 1 10 0 9 13 7 0 7 0 9 2
26 9 11 11 1 0 9 4 13 10 0 9 1 10 9 15 4 13 1 14 13 9 3 1 10 9 2
22 0 9 13 16 10 9 1 12 9 2 3 12 9 4 4 13 3 1 9 0 9 2
13 9 13 3 0 9 1 10 12 15 13 3 3 2
17 15 4 3 13 3 1 14 13 9 1 3 9 2 9 7 9 2
50 15 4 13 0 14 13 0 9 1 9 1 9 1 10 9 15 13 2 7 1 10 9 15 1 9 4 13 1 10 0 9 4 9 0 2 7 1 10 9 3 0 7 15 9 13 1 10 0 9 2
32 1 10 9 9 2 3 0 13 15 3 2 1 0 9 4 9 13 16 15 13 1 3 0 9 15 9 9 3 4 13 15 2
34 1 10 9 3 9 3 3 4 10 0 0 9 2 13 9 14 13 9 1 10 0 9 1 10 9 1 10 9 15 13 1 9 3 1
16 9 13 10 0 9 1 9 7 13 3 10 9 1 9 9 2
18 15 13 3 1 9 1 9 2 3 1 15 1 9 7 13 1 9 2
15 1 10 9 13 9 7 10 9 15 13 9 0 1 0 9
11 9 11 11 13 10 2 9 2 1 9 2
10 15 4 4 13 0 9 1 10 0 9
18 1 3 9 13 9 10 0 3 9 1 9 9 1 10 3 0 9 2
17 9 4 0 1 9 15 4 0 1 9 2 7 13 3 0 9 2
10 10 0 9 1 9 4 10 0 9 2
19 9 1 9 1 11 13 3 0 9 7 3 12 9 7 13 3 3 1 9
6 9 4 9 1 0 9
20 1 10 0 4 0 9 13 9 1 9 7 9 1 9 1 9 7 3 9 2
13 16 15 4 13 9 0 7 9 7 3 4 0 2
21 7 10 0 9 13 3 16 9 4 1 9 14 13 10 0 9 7 3 13 15 2
12 9 1 15 13 3 1 9 10 0 0 9 2
10 7 3 9 1 15 4 13 0 9 2
23 3 4 9 9 1 10 9 7 9 0 1 0 9 9 2 7 0 9 4 3 3 0 2
9 10 9 15 13 1 15 13 9 2
3 9 7 9
11 10 9 13 10 9 3 1 0 0 9 2
11 15 13 15 0 2 9 13 2 13 15 2
27 15 13 3 3 16 10 0 9 13 9 7 4 10 0 9 1 10 0 9 1 9 1 0 7 0 9 2
32 16 10 0 9 13 0 2 4 9 13 10 9 1 3 9 2 10 9 9 2 15 13 1 16 0 9 1 9 13 1 9 2
13 0 9 13 3 7 3 7 13 9 1 0 9 2
21 15 13 0 9 3 7 4 13 1 2 9 2 7 9 2 9 7 2 9 2 2
13 11 4 1 10 9 1 9 13 0 9 1 9 2
12 15 13 15 1 16 9 13 3 3 9 13 2
44 16 15 13 3 1 9 2 7 16 9 13 3 3 0 9 2 7 16 9 13 3 16 9 13 0 2 4 15 13 0 7 0 7 1 3 3 0 16 15 3 3 4 13 2
1 9
21 0 9 7 10 0 4 13 0 7 13 1 10 3 7 3 0 9 2 10 9 2
27 15 4 3 0 14 13 10 9 1 0 9 1 9 7 10 9 15 3 13 9 7 15 3 13 13 9 2
13 10 0 9 2 7 9 7 9 2 13 3 9 2
14 15 13 0 0 9 7 4 13 1 0 7 0 9 2
21 15 4 0 14 13 1 0 7 0 9 16 0 9 4 13 0 9 7 9 9 2
13 0 9 9 1 9 0 7 0 9 4 3 0 2
11 3 3 13 4 0 9 13 1 0 9 2
9 0 9 13 3 0 14 13 15 2
13 15 13 10 0 7 0 9 2 15 10 3 0 2
16 1 0 9 4 0 9 13 1 16 15 4 13 10 0 9 2
11 15 13 15 0 2 2 1 0 9 2 2
13 15 4 13 15 7 9 2 9 2 9 7 9 2
9 3 13 15 1 9 1 9 9 2
10 1 0 9 13 0 9 10 0 9 2
16 15 13 10 12 0 1 10 3 0 9 2 10 0 7 9 2
3 10 0 9
13 0 9 13 1 3 0 9 1 0 9 3 9 2
11 9 4 13 3 0 16 10 9 13 0 2
19 1 0 9 4 15 13 9 3 2 7 15 4 3 13 0 9 1 9 2
10 15 4 13 1 10 9 7 13 0 2
6 3 9 9 4 13 2
9 1 9 4 9 1 9 3 0 2
11 10 9 4 3 0 1 9 7 1 9 2
12 3 12 9 1 9 4 13 7 13 10 9 2
5 9 2 10 0 9
10 3 3 0 7 10 0 9 4 9 2
17 16 15 13 10 3 0 9 1 10 0 9 2 4 15 3 0 2
19 3 9 1 15 15 13 4 3 13 1 0 9 7 1 9 1 10 9 2
10 1 11 13 12 9 1 9 1 9 2
7 9 9 13 3 0 9 2
19 3 4 15 3 9 1 12 0 9 7 10 0 9 1 9 1 0 9 2
9 15 13 1 9 1 9 7 9 2
6 9 1 9 4 13 2
10 9 2 0 9 7 9 4 0 9 2
16 10 0 4 3 13 0 7 0 2 13 1 9 7 13 9 2
15 1 0 9 13 9 0 7 0 14 13 1 9 7 9 2
32 1 0 9 4 15 13 3 10 9 1 10 0 3 3 0 7 9 3 0 2 16 10 9 13 3 0 7 3 3 3 0 2
28 16 15 1 3 0 9 1 0 9 4 13 0 9 1 0 9 2 13 15 15 16 9 4 4 13 1 9 2
10 10 0 9 13 1 14 13 10 9 2
5 0 9 1 0 9
22 16 0 1 9 0 9 13 0 7 0 4 9 13 1 0 9 7 3 13 15 1 2
12 0 9 4 3 9 2 9 2 9 7 9 2
6 9 1 9 7 9 2
9 10 0 9 4 3 13 10 9 2
18 3 4 15 1 9 7 1 0 9 13 3 9 1 0 7 0 9 2
17 15 4 13 9 7 9 7 9 2 0 9 7 9 7 9 3 2
21 10 9 4 13 7 13 3 0 9 1 14 13 9 2 7 15 13 3 0 9 2
21 7 13 9 1 9 3 0 1 15 7 7 13 15 10 0 9 1 9 7 9 2
27 1 10 0 12 9 4 10 0 0 9 1 9 13 7 13 2 15 13 3 0 7 3 0 9 1 9 2
13 15 13 9 7 4 13 0 9 1 9 1 0 2
4 0 9 1 9
23 3 1 10 9 4 13 10 9 1 9 2 15 13 9 1 10 9 1 10 0 1 9 2
18 1 15 13 0 9 2 15 13 10 0 9 1 9 1 9 1 9 2
27 15 4 13 15 16 10 9 1 9 13 1 16 9 1 0 9 1 9 13 3 1 9 7 9 7 9 2
10 1 9 13 9 7 9 4 13 9 2
17 15 13 3 10 0 7 10 0 9 2 13 9 12 7 12 2 2
7 9 4 13 1 12 9 2
10 10 0 13 1 10 0 2 0 9 2
15 3 10 9 1 15 13 0 9 7 13 15 1 14 13 2
24 1 11 13 10 9 2 11 2 15 9 1 9 9 4 13 1 14 13 9 1 9 7 9 2
15 1 12 4 15 13 10 9 0 9 1 9 1 10 9 2
22 15 1 15 4 9 2 15 13 10 3 0 9 7 15 1 9 13 1 0 0 9 2
11 1 0 9 4 15 3 13 1 0 9 2
13 9 4 3 13 10 9 9 2 15 13 10 9 2
8 9 2 1 10 9 9 13 2
18 10 9 1 3 3 0 9 2 9 2 4 13 0 9 7 0 9 2
24 15 1 15 2 9 2 13 1 9 11 7 13 7 10 0 9 1 9 7 3 1 0 9 2
19 10 0 4 11 2 15 13 1 9 7 9 7 3 7 0 9 7 9 2
15 3 0 9 13 10 0 9 1 9 2 1 15 13 9 2
26 15 4 10 0 9 1 10 3 0 2 9 2 2 15 1 10 9 9 3 4 10 3 0 0 9 2
20 15 13 15 4 0 7 13 1 0 9 2 3 15 3 3 13 15 3 3 2
17 10 0 9 1 9 4 10 0 2 0 9 2 15 13 1 9 2
12 1 15 13 9 2 3 10 3 0 4 11 2
23 15 13 3 7 3 1 0 9 7 9 7 4 3 0 2 15 13 16 15 13 7 9 2
16 3 4 15 0 7 4 3 1 11 4 14 13 1 0 9 2
14 15 13 3 0 9 1 0 7 3 0 7 0 9 2
39 15 13 1 9 0 9 7 4 13 1 9 2 7 15 4 1 0 9 4 13 9 2 15 4 10 3 0 9 1 0 9 7 15 0 9 13 9 1 2
24 10 0 9 2 15 4 13 15 4 13 9 1 0 9 2 4 9 9 2 3 0 1 9 2
7 15 13 3 1 0 9 2
1 9
29 1 0 9 4 15 13 7 13 3 1 10 9 9 2 15 13 0 0 9 1 3 9 7 15 3 3 13 9 2
11 1 0 9 4 15 4 0 1 9 9 2
18 1 11 13 15 3 1 11 9 1 9 2 3 1 9 1 0 9 2
6 9 13 1 0 9 2
22 1 10 9 13 9 7 1 9 2 10 9 15 13 1 9 2 13 15 9 1 9 2
19 10 9 4 3 13 9 2 16 15 13 0 9 1 9 1 14 13 15 2
24 7 15 4 13 9 9 2 3 3 16 15 4 13 15 13 9 1 10 9 7 9 1 9 2
10 1 10 0 9 13 9 1 0 9 2
5 9 13 1 9 2
4 9 1 9 2
18 15 4 3 13 9 1 9 0 7 0 9 14 13 10 9 1 9 2
10 15 13 16 15 4 13 3 0 9 2
17 1 11 4 0 9 1 0 9 7 9 13 10 0 9 1 9 2
20 15 13 15 1 10 9 4 2 13 0 9 2 7 13 10 2 0 9 2 2
21 9 13 16 15 3 13 10 0 9 1 9 7 4 4 0 2 3 7 3 0 2
3 9 7 9
22 3 3 13 4 9 7 9 2 3 0 7 0 9 2 4 0 1 10 9 7 3 2
19 15 4 13 15 1 9 1 10 9 1 9 1 14 13 1 10 0 9 2
27 16 15 1 9 4 0 7 1 0 9 13 0 9 4 15 3 13 2 7 15 4 3 13 15 1 9 2
28 1 10 9 13 15 10 0 9 1 10 0 9 3 2 7 1 3 10 9 13 15 0 9 1 9 7 9 2
13 0 1 9 7 9 4 16 15 13 10 0 9 2
12 1 0 9 13 15 10 9 1 9 7 9 2
31 1 9 1 9 7 0 9 13 15 1 16 0 9 2 15 13 10 0 9 1 9 2 4 13 7 3 7 3 13 1 2
6 15 13 7 10 9 2
18 0 9 13 3 0 9 1 0 9 2 3 16 10 0 9 13 1 2
24 16 9 7 0 0 9 7 9 13 0 9 2 4 9 3 13 1 10 0 9 1 10 9 2
5 9 13 3 1 9
16 0 9 1 9 7 9 13 3 1 16 9 13 15 1 15 2
10 15 13 3 0 9 1 14 13 9 2
11 1 0 7 0 9 4 3 10 9 13 2
24 15 13 10 9 7 9 1 9 1 9 7 3 7 3 0 0 7 0 9 16 3 9 13 2
9 9 13 9 7 9 7 4 0 2
5 3 0 4 9 2
14 3 1 10 9 9 3 1 9 4 9 7 9 13 2
30 9 4 13 12 9 2 7 16 9 13 13 0 9 1 9 1 9 7 9 7 0 1 9 1 9 2 9 7 9 2
12 0 9 1 9 4 10 0 15 3 13 9 2
11 15 13 3 0 9 16 15 13 3 3 2
21 10 3 0 0 9 13 10 9 2 7 15 13 3 0 9 7 13 3 0 9 2
14 15 13 9 2 15 4 13 1 9 16 0 9 13 2
37 10 9 2 15 3 13 0 9 2 3 9 7 9 2 13 3 10 0 9 2 7 15 4 13 1 10 0 0 9 7 1 0 9 1 0 9 2
26 9 1 9 7 9 1 0 9 4 13 10 0 9 2 3 1 9 2 16 9 13 1 7 9 13 2
16 10 0 9 13 3 1 16 10 9 3 13 1 9 7 9 2
3 9 7 9
21 3 9 4 13 1 9 7 9 2 4 15 3 13 9 1 10 0 9 1 9 2
9 1 9 13 3 9 1 9 9 2
26 15 1 9 13 3 1 9 7 9 2 15 13 1 16 9 7 9 3 13 10 0 9 1 0 9 2
35 10 0 9 2 15 3 4 0 16 10 9 4 4 13 1 9 7 9 2 4 3 1 0 9 13 9 1 14 13 9 1 9 7 9 2
21 3 13 10 2 9 2 1 16 10 0 3 13 1 3 0 9 1 9 1 9 2
22 1 10 9 13 10 3 0 7 0 9 2 3 15 4 13 13 9 14 13 1 9 2
17 1 10 9 3 4 9 13 3 0 16 15 13 10 0 9 9 2
28 9 7 9 4 1 9 2 9 2 9 7 0 9 13 13 9 7 9 1 9 1 10 9 15 13 13 9 2
24 9 1 9 13 16 15 7 15 4 13 9 14 13 10 3 0 2 3 0 7 3 0 9 2
7 9 1 9 7 3 3 9
16 1 9 13 9 3 1 9 1 9 7 1 9 1 0 9 2
9 15 13 0 14 13 7 13 9 2
12 15 4 1 9 13 16 10 0 9 13 9 2
6 9 13 1 0 9 2
24 9 1 12 9 7 9 13 15 0 1 9 2 7 10 9 4 10 0 1 10 9 1 9 2
12 10 9 15 4 3 0 1 0 9 13 3 2
14 9 4 0 1 14 13 1 14 13 10 9 1 9 2
14 15 13 3 10 0 9 1 9 15 13 1 0 9 2
8 1 9 13 3 9 1 9 2
12 9 13 13 3 9 1 10 0 9 1 9 2
13 15 13 9 7 9 1 14 13 0 9 1 9 2
18 10 9 1 0 9 4 3 10 9 15 13 1 9 15 13 3 9 2
21 15 4 3 1 9 13 10 9 1 0 9 2 3 16 10 9 13 9 1 9 2
10 3 0 9 13 3 13 9 1 9 2
14 16 12 9 13 12 2 4 0 9 9 12 3 12 2
22 9 13 2 15 13 9 1 9 7 9 2 3 0 9 1 9 13 0 9 1 9 2
27 15 13 16 10 0 9 1 9 3 3 4 13 1 9 7 2 7 10 9 1 10 0 9 2 0 9 2
9 10 0 9 4 3 1 15 0 2
16 9 13 14 13 7 10 0 0 9 1 9 1 9 4 13 2
19 15 4 0 16 9 13 0 9 1 10 0 9 1 9 15 15 13 1 2
7 10 9 4 13 0 9 2
17 9 1 0 13 3 0 7 0 9 4 13 9 9 1 9 9 2
20 9 4 3 13 1 9 1 9 2 15 15 3 4 13 1 9 10 0 9 2
16 1 14 13 1 0 9 7 1 14 13 9 3 13 3 9 2
7 15 13 0 9 1 9 2
15 15 13 0 9 1 16 9 7 9 4 4 13 1 9 2
18 15 13 9 2 3 16 0 9 3 4 13 1 1 9 1 0 9 2
7 15 13 3 10 0 9 2
17 9 1 9 15 13 1 12 13 3 1 10 9 15 13 10 9 2
25 1 9 0 3 13 15 3 10 0 9 2 15 13 15 1 9 2 9 7 9 1 9 1 9 2
24 1 10 9 13 15 13 9 1 9 1 9 2 7 3 1 9 13 15 10 0 9 1 9 2
5 10 0 9 13 9
9 1 9 13 10 3 0 9 9 2
11 9 1 15 4 13 0 1 9 1 9 2
19 15 4 13 1 14 13 3 9 2 13 9 7 3 13 9 1 0 9 2
25 1 16 10 9 4 13 13 9 4 15 4 3 0 16 15 1 9 13 3 12 9 1 12 9 2
14 15 4 3 4 0 1 9 2 9 2 9 7 9 2
17 0 9 1 10 0 9 4 4 13 3 12 9 1 10 9 9 2
8 3 3 4 0 9 14 13 2
14 1 9 13 2 9 2 3 0 9 7 9 7 9 2
9 9 13 3 0 3 9 4 13 2
6 9 4 3 3 13 2
20 1 14 13 3 1 10 9 4 15 3 3 0 14 13 1 9 7 13 9 2
9 15 4 3 3 13 7 13 9 2
14 0 9 1 9 7 9 4 3 0 4 13 9 9 2
16 1 10 0 9 4 15 15 13 0 9 4 13 15 7 3 2
6 9 13 9 1 9 2
11 9 13 3 2 3 7 3 9 4 13 2
11 9 1 15 4 10 9 7 9 9 13 2
21 7 9 1 9 13 9 1 0 9 1 9 7 9 1 9 2 3 9 1 9 2
18 9 13 3 2 1 0 9 2 1 10 0 9 1 10 9 15 13 2
17 0 9 7 0 9 13 3 3 9 14 13 9 1 14 13 9 2
12 9 3 1 9 12 13 9 9 1 0 9 2
5 9 9 1 0 9
28 1 14 13 9 2 9 7 9 1 0 9 15 13 3 0 2 13 9 1 9 1 1 9 9 3 0 9 2
4 0 9 1 9
17 1 10 0 9 15 13 3 12 4 9 13 0 0 9 1 9 2
7 15 4 13 14 13 9 2
17 9 4 4 3 0 16 15 4 13 1 14 13 9 1 0 9 2
24 9 4 13 1 10 0 9 2 7 9 4 13 15 10 9 1 16 9 3 4 13 0 9 2
9 9 4 3 13 9 7 0 9 2
16 0 10 9 7 9 4 13 16 10 0 9 13 10 0 9 2
9 3 12 4 10 0 9 3 13 2
6 10 0 9 4 13 2
12 1 9 4 10 0 9 1 10 9 13 15 2
39 1 9 14 13 10 0 9 1 15 4 13 3 9 2 10 9 13 16 10 9 1 10 9 1 10 9 15 4 13 3 15 4 0 2 13 3 1 9 2
28 1 10 9 1 9 1 9 13 3 10 9 1 10 9 2 13 3 2 15 4 13 1 9 1 9 1 9 2
4 3 13 9 2
26 15 4 1 9 9 13 15 1 16 10 9 15 13 0 9 7 9 1 0 9 13 15 3 0 9 2
12 15 13 3 3 1 9 10 9 12 0 9 2
11 3 13 15 10 0 9 7 9 1 9 2
8 9 13 1 9 14 13 9 2
14 1 3 9 4 15 13 16 10 0 9 13 9 3 2
2 9 9
8 1 9 13 15 9 1 9 2
9 15 13 3 3 13 10 0 9 2
20 9 13 16 15 4 13 3 15 4 13 16 9 3 3 13 1 10 0 9 2
8 1 9 13 9 3 12 9 2
12 1 9 1 9 13 15 3 1 3 12 9 2
22 15 4 3 3 13 3 1 16 9 1 9 3 3 4 13 3 1 9 3 9 13 2
8 9 1 10 0 9 4 0 2
24 1 9 13 9 1 0 9 1 12 9 9 2 7 2 1 3 0 9 2 1 10 0 9 2
22 1 9 9 4 15 4 0 14 13 9 9 1 3 0 9 1 9 7 9 1 9 2
10 9 4 3 13 3 2 3 1 9 2
17 9 4 13 9 1 0 9 15 13 1 9 1 9 1 9 9 2
21 16 9 4 0 2 4 0 9 13 0 7 15 15 13 9 2 15 4 13 0 2
23 3 10 9 1 9 9 4 16 15 4 0 14 13 9 1 10 0 9 3 15 13 9 2
5 15 4 13 9 2
29 7 10 9 1 16 9 13 1 9 4 9 1 3 10 9 7 9 4 13 3 0 9 3 16 15 13 0 9 2
6 1 9 13 9 3 2
19 3 4 0 3 0 2 0 9 4 3 0 7 0 9 3 1 9 9 2
27 10 9 2 15 3 13 0 9 2 4 13 7 3 0 2 3 3 15 13 1 9 1 0 9 1 9 2
7 12 2 0 9 7 0 9
9 9 12 13 10 0 9 1 9 2
9 3 13 12 9 9 1 0 9 2
14 10 0 9 13 16 9 13 1 9 1 9 7 9 2
10 15 13 3 9 0 9 1 10 9 2
16 10 9 14 13 3 9 1 0 9 7 14 13 9 4 13 2
18 10 0 9 13 3 1 16 9 3 1 12 13 3 1 10 0 9 2
27 9 1 10 3 10 0 9 9 1 10 9 12 0 9 4 3 4 13 15 7 1 9 1 9 7 9 2
14 10 9 15 4 13 1 9 12 13 3 1 10 9 2
21 1 14 13 9 9 1 9 1 0 9 7 9 4 3 12 13 0 7 0 9 2
41 10 9 2 15 13 3 7 3 4 0 1 10 9 1 16 9 3 13 1 9 2 13 1 9 1 0 12 9 2 9 2 9 7 9 9 7 1 0 9 9 2
9 3 12 9 4 0 1 0 9 2
7 4 15 13 3 1 9 2
8 9 1 11 4 4 3 0 2
12 9 9 14 2 13 3 2 9 4 3 13 2
22 1 0 0 9 4 15 13 9 1 12 9 1 9 12 1 3 12 1 9 1 9 2
28 1 9 1 9 1 9 1 9 2 0 9 7 0 9 1 9 4 9 1 0 9 3 3 13 9 1 9 2
10 15 13 15 4 10 0 9 1 9 2
4 9 13 9 2
11 1 0 9 13 15 3 14 13 3 9 2
4 9 13 9 2
8 1 9 4 9 13 1 11 2
6 9 13 9 1 11 2
7 9 13 10 9 2 9 2
15 9 4 2 13 15 2 13 3 16 9 4 13 1 9 2
13 16 9 1 10 9 13 1 9 4 10 9 13 2
13 3 9 13 1 9 2 4 9 13 1 0 9 2
12 1 11 13 9 2 15 13 9 1 0 9 2
12 9 2 3 1 9 2 13 0 9 1 0 2
15 10 9 4 3 1 0 9 3 0 9 1 10 0 9 2
19 16 0 9 13 16 9 13 1 9 2 4 15 14 4 13 1 0 9 2
19 13 3 9 13 1 9 2 13 3 10 9 3 9 13 9 7 9 13 2
14 15 3 13 16 10 9 3 13 9 2 3 13 15 2
11 0 9 14 13 9 13 14 13 3 3 2
9 9 4 3 15 15 13 1 9 2
27 13 15 3 9 1 16 10 9 4 13 3 14 13 2 4 15 0 16 10 0 9 4 13 9 1 9 2
15 13 15 3 0 9 1 9 9 7 9 4 15 13 3 2
33 3 2 7 1 3 0 0 9 2 4 15 13 9 1 10 9 3 9 4 13 1 7 0 9 7 1 10 9 10 9 13 1 2
9 3 3 13 11 1 10 0 9 2
24 9 13 12 9 9 2 12 9 9 15 13 1 10 9 7 12 3 15 1 15 15 4 9 2
10 2 9 2 9 9 12 9 12 2 2
3 9 7 9
4 9 7 9 2
16 3 13 15 2 3 0 4 15 1 0 9 7 1 0 9 2
7 0 9 2 15 4 15 2
6 4 15 10 0 9 2
4 9 7 9 2
10 9 1 9 2 9 1 9 7 9 2
11 9 2 4 15 13 1 15 7 0 9 2
6 15 13 3 10 9 2
12 9 9 13 1 3 7 12 9 9 1 9 2
9 1 12 9 13 9 9 4 0 2
13 10 0 9 4 16 9 3 13 1 9 1 9 2
6 3 3 4 9 0 2
18 12 9 1 9 10 9 4 3 13 15 0 7 9 13 1 0 9 2
14 15 13 13 1 9 2 9 2 7 9 2 9 2 2
9 9 4 3 0 7 13 0 9 2
20 10 0 1 15 13 1 11 2 1 11 7 11 7 1 11 7 1 0 11 2
18 9 4 1 9 9 1 0 9 7 3 1 10 0 9 1 0 9 2
14 15 13 3 3 14 13 10 0 9 1 9 7 9 2
37 9 9 13 3 1 16 15 1 10 9 13 1 9 1 7 1 9 4 13 3 1 10 9 1 3 0 9 7 0 9 1 14 4 13 0 9 2
9 1 9 1 9 13 9 0 9 2
16 15 4 4 13 1 15 3 15 3 13 10 9 1 0 9 2
35 15 1 9 3 0 9 4 1 9 4 14 13 13 10 9 3 16 9 9 4 13 9 3 2 3 3 9 13 1 0 9 1 10 9 2
8 9 1 9 4 13 3 0 2
8 9 4 3 13 1 0 9 2
9 15 4 4 9 7 9 1 9 2
24 15 4 4 9 15 13 3 1 14 13 7 13 9 2 9 7 9 2 9 2 9 7 9 2
19 15 4 4 9 1 9 1 9 1 9 1 0 2 0 7 0 9 3 2
11 9 4 13 1 0 9 7 3 3 11 2
10 7 9 4 1 15 13 1 0 9 2
25 3 13 0 9 1 9 12 3 12 9 0 9 2 3 10 0 9 13 1 11 2 11 7 11 2
17 1 10 9 13 11 12 9 0 1 0 9 1 11 7 0 9 2
15 11 2 11 7 11 13 1 10 9 1 3 12 9 15 2
6 9 4 13 3 9 2
13 3 4 15 3 0 16 0 9 13 3 1 9 2
12 11 4 13 9 1 14 13 10 9 1 9 2
20 9 12 13 15 10 0 9 1 12 9 9 2 12 4 15 13 1 12 9 2
21 9 13 12 16 9 1 9 4 13 2 3 16 15 3 12 13 12 9 1 9 2
12 9 4 3 14 13 3 7 12 9 9 3 2
15 3 12 9 1 9 13 1 11 7 10 9 1 0 9 2
29 10 0 9 2 10 0 0 9 1 9 2 13 1 11 2 0 0 9 9 2 2 15 4 10 0 9 1 9 2
7 11 9 4 14 13 9 2
12 3 13 10 9 1 10 0 9 1 10 9 2
9 11 4 11 9 1 9 7 9 2
13 3 10 9 1 11 2 3 9 13 10 9 0 2
17 9 1 9 13 9 7 13 1 10 9 1 10 0 9 1 9 2
9 9 1 10 9 13 1 11 9 2
7 3 13 9 1 10 9 2
15 15 13 3 3 0 9 15 13 9 1 0 9 1 9 2
5 9 11 12 9 12
16 15 13 3 10 1 15 0 9 1 15 15 13 1 10 9 2
14 10 9 1 15 9 3 13 4 1 9 13 10 9 2
16 1 9 1 10 0 9 13 15 3 9 14 13 15 7 9 2
19 1 9 10 0 9 2 13 3 3 12 9 9 2 12 9 1 9 9 2
32 15 13 1 3 12 9 1 2 9 2 2 13 3 12 9 1 9 7 13 1 9 10 9 1 9 1 3 12 9 1 9 2
21 1 11 13 9 10 9 1 10 9 15 4 0 1 10 0 9 1 11 7 11 2
8 11 13 10 0 1 10 0 2
16 9 4 3 3 3 0 7 11 2 11 13 3 12 9 9 2
16 1 10 9 9 1 9 9 13 11 1 0 12 9 1 9 2
11 9 13 10 9 1 3 12 9 1 9 2
18 1 12 9 1 9 4 9 3 2 3 3 3 2 12 9 1 9 2
11 12 13 12 9 1 10 0 9 1 9 2
14 1 9 13 3 12 9 9 2 12 9 1 9 9 2
11 10 9 1 2 9 2 4 3 12 9 2
10 15 13 1 0 12 9 1 9 9 2
12 15 13 3 10 9 1 9 1 3 12 9 2
9 12 9 1 0 9 9 4 9 2
14 12 9 13 9 2 12 9 9 2 12 9 9 9 2
9 9 13 3 12 9 1 10 0 2
22 9 1 9 7 9 4 3 12 9 2 3 12 1 9 2 1 10 9 1 12 9 2
31 1 11 13 15 3 12 9 1 10 9 2 1 11 3 12 2 1 11 3 12 2 1 11 3 12 2 1 11 3 12 2
7 15 13 3 0 1 9 2
6 10 9 13 1 15 2
10 15 13 0 14 13 10 9 1 15 2
7 15 13 3 3 1 15 2
14 10 0 9 13 15 16 15 13 9 1 10 0 9 2
24 3 4 15 13 0 9 2 15 4 13 9 0 1 0 9 7 3 4 13 10 9 1 15 2
12 15 13 15 1 10 9 3 15 13 1 9 2
14 16 15 13 9 13 15 13 3 1 10 9 15 13 2
10 6 2 10 9 1 11 1 11 11 2
12 15 13 15 1 9 9 15 15 13 3 1 2
12 15 13 3 1 9 7 13 10 9 1 9 2
15 15 13 15 9 2 3 16 15 4 13 3 11 11 9 2
28 10 9 13 1 16 15 4 13 10 9 9 7 16 12 1 15 1 10 9 4 13 9 11 0 1 0 9 2
5 3 13 10 9 2
13 2 9 9 4 14 4 0 7 14 13 9 2 2
9 15 4 13 1 9 1 9 9 2
15 9 4 13 7 9 0 9 1 9 7 3 3 10 0 2
20 15 4 3 13 1 15 15 3 4 4 13 10 0 9 15 10 0 9 13 2
23 9 4 13 10 0 9 1 15 2 13 10 9 2 13 10 9 7 3 13 10 0 9 2
28 1 15 4 15 13 16 15 4 0 1 10 9 2 7 16 15 3 13 15 13 10 9 3 3 14 13 1 2
14 10 3 9 1 9 13 1 9 7 9 9 1 9 2
18 15 13 9 7 9 2 1 15 9 2 15 13 9 3 2 13 15 2
28 15 13 3 1 16 15 13 9 15 13 10 9 7 10 9 1 14 13 15 0 7 10 3 0 9 1 9 2
12 9 7 9 4 3 1 0 9 10 0 9 2
22 3 13 10 9 9 7 10 9 1 16 15 4 15 0 2 7 4 13 15 3 3 2
5 15 13 1 9 2
11 9 4 13 10 9 1 10 0 0 9 2
8 9 7 10 9 4 3 13 2
22 3 3 4 15 0 1 12 3 0 9 14 13 10 0 9 1 0 9 7 0 9 2
15 1 16 15 13 9 13 15 0 14 13 9 3 1 9 2
19 3 4 15 7 15 14 13 10 9 9 2 7 15 13 1 1 14 13 2
26 15 4 3 3 9 1 16 9 4 13 10 0 9 3 3 3 7 16 9 13 10 0 9 1 9 2
14 9 13 15 3 7 3 16 15 13 15 14 13 3 2
14 9 13 10 0 9 7 0 1 14 13 3 10 9 2
16 9 1 9 4 3 4 0 2 7 15 4 4 1 0 9 2
17 3 4 10 9 13 15 1 14 13 7 13 10 0 9 1 9 2
6 3 13 15 3 9 2
10 3 13 9 10 0 9 1 9 9 2
14 13 10 9 15 13 9 1 10 9 1 10 3 0 2
14 15 4 3 0 16 10 9 4 13 0 9 1 9 2
35 4 15 3 13 15 16 9 15 13 1 10 9 1 9 2 9 2 9 2 4 3 0 7 2 3 2 1 9 14 13 9 1 10 9 2
5 3 13 15 3 2
15 3 9 3 7 1 10 9 13 15 10 9 9 7 9 2
32 15 4 3 13 1 10 3 9 3 3 3 2 1 10 9 4 15 3 13 16 15 4 4 13 1 15 15 15 3 4 13 2
18 15 2 7 15 1 15 2 4 13 16 3 9 13 3 4 15 0 2
14 7 3 13 15 1 9 3 15 13 14 13 3 9 2
22 1 9 4 15 3 0 14 13 2 7 15 13 15 2 16 10 9 13 9 1 9 2
10 7 13 15 9 1 1 9 9 3 2
12 9 4 0 7 4 3 13 1 3 0 9 2
9 9 13 1 15 2 15 13 3 2
5 9 9 4 0 2
15 9 13 10 9 16 15 3 1 9 7 9 13 3 3 2
6 7 13 15 3 3 2
12 16 15 3 13 3 4 3 10 0 9 13 2
24 9 4 13 3 10 0 9 1 2 3 0 7 0 9 13 15 1 0 3 9 1 9 2 2
17 3 12 9 1 9 13 1 10 0 9 1 3 12 9 1 9 2
22 9 13 3 0 10 9 14 13 10 0 9 1 9 2 3 3 10 9 1 1 9 2
6 3 4 15 13 15 2
10 3 4 3 9 0 1 10 0 9 2
10 3 13 10 9 3 1 9 7 9 2
25 7 15 4 13 0 9 2 3 15 15 4 13 1 9 7 9 7 9 15 13 15 14 13 9 2
24 7 9 4 15 3 13 1 9 7 9 2 15 4 13 3 0 14 13 2 13 3 0 9 2
16 11 11 4 13 0 9 1 10 0 9 7 10 0 0 9 2
8 15 4 13 1 15 9 13 2
35 9 2 9 2 9 2 15 4 10 0 9 15 13 15 3 1 2 7 15 13 0 14 13 15 15 3 7 3 3 15 13 15 1 9 2
29 7 10 0 9 4 16 9 1 10 0 0 9 7 9 4 13 2 9 4 3 3 10 0 9 1 14 13 9 2
48 15 4 3 10 3 0 9 2 0 1 10 9 9 1 9 7 9 2 1 10 9 1 9 7 9 1 9 1 9 2 1 9 7 9 2 6 3 2 0 9 2 7 0 2 0 2 9 2
25 7 3 13 15 3 3 10 9 1 9 2 15 7 15 1 10 9 2 1 10 9 1 0 9 2
39 10 0 9 4 0 7 10 9 1 10 0 9 15 15 13 1 9 2 9 7 1 9 1 9 1 9 9 4 15 3 13 1 15 1 10 0 0 9 2
20 10 0 9 4 3 9 3 13 9 2 16 9 4 13 2 3 1 0 9 2
59 0 9 9 7 0 9 9 13 3 9 1 0 9 7 9 1 12 9 2 7 9 13 3 3 3 15 15 13 2 3 16 9 1 0 9 13 10 9 1 9 2 7 1 10 3 0 9 2 1 9 2 16 9 1 0 9 13 9 2
14 9 14 13 0 9 4 0 1 9 14 13 1 9 2
86 16 15 13 1 9 7 9 13 13 15 15 3 1 10 0 9 2 9 10 0 7 0 9 1 0 7 0 9 15 13 1 9 1 0 9 2 9 2 10 3 3 0 9 1 9 9 2 10 0 9 3 12 9 13 15 3 1 10 0 9 2 7 3 9 3 3 13 3 1 10 0 9 1 10 0 9 2 3 10 9 1 10 0 9 9 2
17 7 3 9 2 10 3 0 9 2 1 0 2 0 2 0 9 2
31 1 9 0 9 2 1 15 0 2 13 10 0 9 16 9 4 0 2 3 3 0 7 3 0 7 9 15 13 1 9 2
17 10 3 9 13 15 3 1 14 13 9 1 9 2 3 1 9 2
44 3 9 13 7 10 9 1 9 15 4 13 15 1 15 10 0 4 13 1 9 1 9 7 9 2 3 7 10 9 15 13 4 2 3 10 9 13 10 0 9 1 14 13 2
20 15 13 3 10 12 9 1 9 0 9 1 10 0 9 1 10 0 1 9 2
21 10 9 4 3 0 1 9 0 2 7 13 3 10 9 14 2 13 2 10 9 2
20 3 16 15 13 1 9 7 9 4 15 13 9 1 0 9 2 3 1 9 2
33 7 1 9 1 15 2 3 1 10 0 9 2 4 15 13 9 1 16 15 13 1 0 0 9 1 14 13 3 0 9 7 0 2
10 0 9 7 3 0 9 4 0 9 2
15 14 13 10 0 9 3 13 3 7 14 13 9 1 9 2
42 3 4 9 1 3 0 9 0 2 3 11 11 1 9 3 9 13 10 0 9 1 9 2 7 3 10 9 4 13 9 1 10 0 16 9 7 9 3 13 1 9 2
19 9 13 9 1 9 7 13 3 1 10 1 15 0 9 1 9 7 9 2
16 15 1 10 0 4 15 13 3 9 3 13 1 10 0 9 2
31 9 13 1 9 1 9 7 4 1 9 1 9 3 3 0 1 15 2 15 15 3 4 13 10 0 9 7 10 0 9 2
7 9 4 13 0 1 3 2
48 15 13 1 10 9 3 16 10 9 15 13 3 13 3 7 13 1 9 7 9 1 10 0 2 10 0 7 0 9 15 1 9 4 13 0 1 9 7 3 3 0 7 9 1 10 0 0 2
28 3 10 0 13 3 13 13 2 1 9 13 15 3 15 7 10 9 1 0 9 2 3 1 10 0 9 3 2
37 9 1 10 9 13 0 9 1 9 2 9 2 9 2 10 0 9 2 15 3 13 0 9 1 10 0 4 1 9 4 0 14 13 1 9 9 2
23 7 3 13 15 3 15 14 13 1 2 15 4 4 0 7 0 3 14 13 15 10 0 2
25 15 4 0 14 13 9 1 10 0 9 1 12 0 9 2 15 10 9 3 4 13 9 0 0 2
41 7 15 13 3 1 9 3 9 13 2 13 3 7 13 13 1 10 0 0 15 3 13 13 15 15 2 10 0 2 0 2 3 15 0 9 1 9 1 9 3 2
69 13 15 13 1 15 9 13 2 9 7 9 2 9 7 9 2 0 0 14 13 1 7 13 1 2 9 1 0 9 2 9 2 9 2 10 0 9 7 10 9 14 13 1 2 15 15 13 9 7 15 15 13 1 2 15 13 3 14 13 3 2 7 15 4 15 13 3 1 2
7 9 14 13 1 10 9 2
10 3 3 9 7 0 1 9 0 9 2
40 15 4 13 3 3 2 7 1 10 9 13 15 16 15 3 13 1 16 9 4 0 7 0 7 0 2 9 15 1 7 1 15 4 13 10 0 9 3 0 2
31 15 4 3 13 1 16 15 1 9 13 0 7 3 1 10 0 9 14 13 10 9 3 0 1 9 3 9 0 9 13 2
38 15 4 13 1 16 9 13 3 3 3 1 9 2 16 10 3 3 0 9 13 3 0 9 2 16 10 0 9 1 12 7 12 9 13 10 0 9 2
31 15 4 3 3 14 13 15 16 10 0 13 9 1 10 9 1 12 7 12 9 2 3 3 16 15 4 0 1 15 0 2
19 15 13 3 3 16 15 3 13 1 14 4 13 9 1 14 4 13 9 2
18 15 4 3 13 10 9 16 15 13 13 3 3 0 1 10 0 9 2
29 3 13 15 3 13 16 10 10 9 4 13 3 3 15 13 2 9 1 0 0 9 0 1 9 2 9 7 9 2
20 15 1 15 4 3 13 14 13 1 0 0 9 7 13 0 0 9 1 9 2
26 15 4 13 15 3 3 1 9 0 9 2 15 4 3 3 13 3 1 10 3 0 9 2 1 9 2
26 7 9 2 7 4 15 10 9 2 2 13 1 3 3 0 9 2 7 4 10 9 4 13 10 9 2
31 0 1 10 9 3 0 9 1 9 7 1 9 3 3 13 3 15 2 3 9 13 1 3 0 9 1 10 3 0 9 2
39 7 3 3 9 4 3 0 1 14 13 3 1 9 9 13 15 10 9 3 16 15 4 13 10 9 9 16 3 4 15 13 14 13 10 13 13 0 9 2
36 13 15 13 9 11 7 13 9 1 10 0 9 2 0 7 0 9 1 9 2 4 15 3 13 13 0 9 3 3 2 3 3 2 3 3 2
30 1 9 1 14 13 9 1 10 0 0 9 4 15 13 15 1 10 0 9 2 15 13 9 1 9 2 9 2 9 2
40 3 4 1 9 7 9 13 9 1 9 2 9 1 9 2 9 2 9 1 9 2 3 10 9 2 9 2 9 1 9 7 9 2 9 2 3 10 0 9 2
28 1 0 9 3 9 2 7 15 15 4 13 15 2 1 0 9 2 1 10 9 0 9 9 2 9 2 9 2
47 9 9 13 15 15 3 1 9 0 9 1 0 7 0 9 2 0 9 7 9 2 3 15 4 13 15 3 1 9 7 1 10 9 2 7 7 0 7 0 9 3 15 13 10 0 9 2
10 7 10 0 9 4 3 9 7 9 2
22 15 15 4 13 9 4 15 1 9 0 9 7 15 4 13 2 13 7 13 15 3 2
41 10 0 9 4 13 10 2 0 9 2 7 10 9 7 0 9 2 1 15 4 13 7 9 7 9 2 15 1 0 0 9 2 7 15 1 9 1 9 7 9 2
17 0 7 9 4 4 9 1 0 9 2 7 9 14 13 1 9 2
36 9 15 13 1 14 13 3 0 10 9 2 3 4 9 3 13 1 9 2 4 4 13 3 1 10 0 9 7 4 13 1 10 3 3 9 2
43 9 4 1 10 0 9 13 0 9 1 9 7 0 9 2 9 4 13 9 14 13 1 9 2 9 4 13 7 13 2 3 4 10 0 0 9 7 9 13 0 9 3 2
37 2 1 9 4 15 3 3 15 14 13 10 0 9 3 1 9 2 3 9 4 13 2 0 9 4 4 13 9 2 0 9 2 3 1 9 2 2
49 1 9 1 10 0 9 3 9 7 9 4 10 0 2 1 9 2 9 2 9 7 9 2 2 10 0 9 15 3 13 10 0 0 9 2 13 9 7 9 10 0 9 2 1 0 9 1 9 2
24 9 13 1 2 10 2 9 2 7 13 9 3 15 13 2 7 9 9 13 9 1 0 9 2
47 9 7 9 4 1 9 0 9 13 0 9 14 13 0 3 2 7 15 4 0 1 10 0 9 3 7 9 3 4 13 15 0 1 10 3 0 9 2 16 9 4 3 0 1 0 9 2
19 9 13 10 0 0 7 10 0 0 9 0 15 15 3 13 10 0 9 2
10 0 9 4 3 10 0 9 7 3 2
35 9 13 10 9 16 15 13 3 0 2 7 2 16 9 3 3 4 0 1 10 9 2 4 15 3 1 0 9 13 3 0 9 14 13 2
21 10 9 15 4 10 9 1 10 9 9 15 3 13 1 9 4 0 1 0 9 2
21 3 3 4 10 3 0 9 14 13 10 0 9 2 7 15 4 3 13 10 0 2
18 15 4 13 10 0 2 0 9 2 3 0 14 13 3 10 0 9 2
15 15 13 3 0 16 15 1 9 13 16 9 13 0 9 2
36 14 1 10 9 3 13 16 10 9 4 0 2 1 9 2 4 1 10 0 0 9 4 3 0 2 1 15 13 15 3 3 3 15 15 13 2
23 15 13 3 16 9 4 0 1 0 9 2 7 9 4 13 10 0 9 1 9 1 11 2
8 15 4 3 3 13 15 9 2
30 3 4 3 15 9 13 3 0 1 0 9 1 9 7 3 13 15 1 15 3 0 16 15 13 9 1 14 13 9 2
13 7 4 15 0 1 9 7 3 4 10 9 13 2
3 3 15 2
36 16 9 13 4 3 3 0 2 7 16 15 13 15 3 13 15 13 10 9 1 9 1 16 12 9 13 1 15 15 4 13 1 12 9 3 2
14 15 4 3 3 3 9 1 10 0 9 1 0 9 2
15 10 2 0 2 9 4 13 15 15 7 3 3 13 15 2
35 3 0 4 16 9 1 9 7 9 13 1 10 9 15 13 9 1 9 7 9 1 10 9 15 1 10 0 9 7 1 9 4 3 0 2
20 0 9 11 13 3 1 10 9 10 9 2 0 2 1 3 0 9 1 9 2
33 1 9 4 9 13 7 10 9 14 13 9 7 3 13 9 1 10 9 3 10 0 4 13 9 1 15 0 1 3 9 1 0 2
13 9 4 10 9 1 2 0 9 1 0 9 2 2
19 3 13 9 1 0 9 2 15 7 15 4 3 3 13 15 0 1 9 2
19 10 0 9 4 13 7 13 15 1 0 9 1 16 10 9 4 3 13 2
24 1 9 13 15 3 1 9 9 2 1 9 7 1 16 15 1 9 13 3 9 13 1 9 2
30 9 9 16 9 1 9 9 4 13 1 0 9 7 16 15 7 15 1 10 9 4 13 1 9 4 1 10 0 0 2
19 10 0 9 2 15 4 13 1 10 9 2 4 14 1 9 13 10 9 2
20 1 10 9 9 15 15 13 1 4 15 13 1 14 3 13 15 15 4 0 2
30 1 10 3 0 4 13 9 9 14 13 9 1 15 2 14 13 14 13 1 2 9 2 1 9 1 1 2 9 2 2
13 9 2 9 7 9 0 9 1 15 13 3 9 2
10 1 10 9 4 3 10 9 3 0 2
20 1 10 0 4 3 9 1 14 13 1 0 9 1 10 0 13 10 0 9 2
17 1 9 4 15 3 0 14 13 16 9 13 3 2 1 0 2 2
3 9 7 9
29 0 9 11 11 13 1 10 9 10 9 2 2 1 9 1 9 2 3 15 13 10 0 9 9 1 9 1 11 2
36 1 9 13 3 2 16 10 9 4 13 7 0 1 10 0 9 9 7 16 10 9 1 0 9 3 3 13 1 10 9 15 13 3 1 9 2
11 10 9 13 15 3 15 13 9 1 0 2
14 15 4 1 9 9 13 9 1 9 1 9 7 9 2
16 16 10 0 9 13 10 9 1 9 3 4 9 7 9 13 2
13 9 4 3 0 1 10 9 3 9 3 4 0 2
22 9 0 9 4 3 10 0 9 4 13 2 7 9 1 10 9 4 3 13 1 9 2
21 9 4 3 1 10 9 0 2 3 16 9 1 9 1 10 0 13 9 7 9 2
17 9 1 9 1 10 9 13 9 1 9 1 0 9 7 0 9 2
20 9 13 3 10 0 2 9 13 1 0 9 2 9 15 10 0 9 3 13 2
20 9 0 9 2 10 0 9 1 9 9 2 13 16 10 9 1 10 9 13 2
18 15 13 3 1 16 9 13 1 10 3 0 9 1 9 1 9 9 2
22 10 0 9 1 14 13 3 9 1 9 13 3 3 3 16 15 4 13 9 1 9 2
22 3 13 1 10 9 3 9 16 15 1 10 0 9 1 9 4 13 3 10 0 9 2
27 9 4 10 0 0 9 14 13 3 9 1 9 7 3 13 16 9 13 10 0 9 15 13 1 10 9 2
14 10 0 9 16 9 4 9 9 13 1 10 0 9 2
10 9 4 10 9 2 7 10 0 9 2
13 15 13 9 1 9 9 7 1 15 7 1 9 2
13 9 1 9 13 9 7 9 13 3 1 0 9 2
27 2 9 4 1 11 0 2 13 15 1 9 2 7 1 10 0 9 13 9 9 10 0 7 3 0 9 2
13 15 4 13 15 10 0 9 1 9 7 10 9 2
6 4 15 0 1 9 2
21 9 4 16 15 1 10 0 9 3 3 4 13 3 9 1 14 13 10 0 9 2
8 15 13 3 16 15 13 15 2
30 10 0 0 9 15 13 9 13 1 16 15 3 0 13 3 9 7 0 9 7 13 3 3 9 1 9 1 9 9 2
20 3 13 16 10 0 9 4 4 0 1 0 9 2 7 0 9 4 3 13 2
27 16 15 3 4 3 0 1 16 10 1 10 9 0 9 4 9 2 3 13 15 3 16 15 13 0 9 2
16 15 13 1 9 16 15 4 13 9 1 15 15 4 13 9 2
7 3 13 3 9 0 9 2
25 15 13 10 9 0 1 15 9 4 1 16 9 2 1 7 1 9 2 13 1 16 9 13 15 2
5 15 4 13 9 2
9 15 0 9 4 1 0 9 12 2
14 15 4 3 0 14 13 15 2 15 13 3 3 1 2
15 15 4 3 2 13 15 2 2 2 3 3 12 9 2 2
15 9 4 0 3 14 13 15 1 0 9 2 13 15 2 2
17 15 13 10 0 9 13 9 1 0 16 9 3 3 4 13 9 2
19 1 9 4 15 13 16 3 10 9 4 4 13 10 0 9 1 9 9 2
14 3 4 3 15 7 15 1 0 9 13 9 1 9 2
17 15 15 13 13 3 4 10 0 9 1 10 9 15 9 9 13 2
32 16 15 2 13 15 2 10 9 2 3 1 9 3 9 1 9 9 13 2 4 9 3 4 0 16 9 13 2 3 0 9 2
26 1 9 15 13 9 4 15 4 10 9 16 1 9 4 13 2 2 13 15 15 7 9 7 9 2 2
25 10 0 9 4 1 0 9 13 9 7 13 1 16 9 1 9 9 13 1 9 1 10 0 9 2
40 3 4 15 4 0 16 15 13 9 9 1 10 3 0 9 1 9 2 3 15 4 13 7 1 9 1 9 7 1 0 9 1 15 15 13 10 3 3 9 2
17 3 13 15 1 0 9 16 2 15 4 4 0 14 13 15 2 2
8 15 13 3 3 15 4 0 2
22 16 15 4 13 1 0 9 14 13 9 13 15 15 1 14 3 1 9 13 1 9 2
14 0 9 4 3 4 10 0 9 2 3 9 1 15 2
23 10 0 9 1 16 15 3 13 15 2 15 4 3 13 15 2 4 15 3 13 1 9 2
20 15 4 13 7 10 9 1 10 0 9 14 13 9 7 7 10 9 1 9 2
16 1 10 9 9 13 1 9 4 15 3 0 13 9 9 1 2
32 3 4 15 13 3 2 16 4 10 9 13 10 0 0 9 7 9 13 9 3 4 10 9 13 1 9 7 16 9 13 9 2
27 1 10 9 4 10 0 9 13 1 14 13 3 10 3 0 9 15 13 3 9 13 1 9 7 1 9 2
34 1 10 9 4 15 13 10 0 9 9 2 15 13 1 14 13 9 9 1 7 15 3 13 10 9 1 15 15 13 1 10 0 9 2
15 16 9 4 13 15 1 0 9 4 1 10 0 9 0 2
24 15 15 15 13 3 13 4 7 16 9 3 3 4 0 7 16 15 1 10 9 3 4 0 2
16 3 7 3 4 3 10 0 9 13 0 2 7 3 13 9 2
6 9 7 9 13 3 2
29 3 4 9 7 9 13 1 10 0 9 2 7 10 0 13 1 3 9 10 9 1 10 9 15 1 9 4 0 2
25 4 9 13 7 13 9 13 9 3 3 10 9 1 10 9 15 15 13 7 13 1 3 1 9 2
10 3 3 9 1 15 13 0 1 9 2
27 15 4 13 16 10 15 15 3 13 1 15 16 10 9 4 13 10 9 13 9 1 16 9 7 9 13 2
7 15 13 0 9 1 9 2
14 15 4 0 3 3 0 9 13 1 9 1 0 9 2
16 1 10 0 0 9 4 15 3 1 10 9 13 9 3 0 2
8 3 13 15 1 0 0 9 2
1 9
8 9 4 3 3 0 1 9 2
15 1 9 9 13 3 1 0 0 9 0 1 9 1 0 2
13 3 16 15 3 13 1 9 9 4 15 10 9 2
25 10 0 9 13 3 0 14 13 3 10 9 1 9 2 3 16 15 1 9 13 1 9 9 2 2
12 10 0 9 13 1 9 9 2 3 1 0 2
11 1 0 2 9 2 4 15 13 0 9 2
29 9 4 13 1 10 2 0 2 1 3 0 9 7 16 9 9 13 3 2 15 13 0 7 0 9 1 0 9 2
6 3 4 10 9 13 2
26 15 4 3 13 16 9 13 1 9 2 7 15 4 13 0 9 16 0 9 3 13 0 9 7 15 2
12 15 13 1 9 10 9 7 9 1 0 0 2
14 1 14 13 9 13 15 10 9 7 15 13 15 0 2
23 15 4 1 9 13 13 10 9 0 1 9 9 1 2 7 10 9 13 10 9 1 9 2
18 15 13 3 2 16 15 4 13 1 10 9 15 13 15 13 9 9 2
18 10 0 9 13 3 1 15 15 13 1 0 9 0 9 1 0 9 2
19 9 9 13 3 0 9 1 10 0 9 2 7 10 9 4 13 1 9 2
21 15 4 3 9 9 14 1 0 13 9 1 9 2 15 4 10 9 1 0 9 2
29 10 0 9 1 9 7 9 4 13 9 1 9 2 9 4 13 10 0 9 7 9 4 13 0 9 1 10 0 2
12 3 4 15 13 9 1 9 2 16 9 13 2
