4477 11
18 11 13 10 9 15 13 1 9 11 2 9 11 2 11 11 2 11 2
21 10 9 9 3 13 1 9 7 1 13 10 9 7 13 10 9 16 15 13 9 2
30 9 10 13 1 9 11 15 13 9 11 11 7 11 2 7 1 9 12 1 11 11 1 9 9 15 3 13 1 9 2
49 1 9 0 2 12 9 9 2 11 7 11 2 11 13 10 9 9 1 9 1 9 11 2 16 13 9 1 1 9 2 9 3 3 13 12 7 12 9 9 1 9 9 9 11 1 3 13 9 2
16 11 9 9 13 12 2 12 9 2 1 1 9 9 11 11 2
22 11 11 15 3 13 9 15 3 15 13 10 13 1 11 11 1 13 13 1 11 11 2
11 11 3 15 0 9 13 9 9 1 9 2
27 11 10 3 13 1 9 0 1 9 11 2 11 11 2 2 11 11 11 2 7 9 2 11 11 11 2 2
10 16 13 10 9 15 13 13 9 9 2
35 9 9 11 11 10 13 1 10 9 0 1 1 1 9 11 11 2 11 15 9 9 13 13 1 11 11 11 1 9 9 2 12 2 12 2
17 15 3 1 10 0 9 9 15 13 16 9 1 11 11 3 0 2
23 9 10 13 9 15 13 2 11 11 2 9 13 0 12 9 1 11 15 13 1 9 10 2
19 11 11 13 10 9 1 11 11 11 2 11 2 11 2 13 1 11 11 2
48 9 10 13 1 9 13 13 0 2 1 13 9 16 9 9 13 1 11 1 3 3 0 1 9 1 13 9 0 9 10 13 1 9 9 9 11 11 11 12 1 12 9 9 9 1 9 0 2
10 11 10 13 1 11 11 12 1 11 2
19 14 13 9 9 11 2 13 1 9 2 9 0 2 7 9 9 13 9 2
17 11 11 11 13 2 2 9 15 1 0 14 13 9 11 2 11 2
18 11 11 7 9 9 0 13 1 9 9 12 2 12 7 12 2 12 2
7 9 10 9 1 9 9 2
10 9 15 15 13 2 7 9 15 13 2
19 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 7 11 11 2
8 9 9 0 0 7 0 0 2
8 10 9 9 5 9 9 11 2
13 3 3 15 14 13 9 15 0 3 10 9 10 2
29 11 2 11 13 11 11 5 11 11 11 11 11 2 15 13 1 9 12 9 9 9 11 11 1 9 12 2 12 2
55 11 7 11 13 9 9 11 11 15 13 12 9 0 2 2 11 7 11 2 2 2 11 11 2 2 7 2 11 11 11 2 2 7 9 13 9 2 9 15 13 1 9 2 9 9 11 0 7 9 2 9 11 5 11 2
44 9 10 3 13 1 9 9 15 13 9 1 9 0 15 3 13 1 10 9 9 0 2 7 9 9 9 15 13 9 1 9 2 7 13 9 15 3 13 13 9 1 9 9 2
16 11 13 11 1 9 11 11 2 11 11 11 2 11 2 11 2
17 11 1 9 13 9 1 11 2 11 11 12 13 11 0 7 0 2
15 11 11 11 2 2 13 10 9 7 9 9 9 9 11 2
26 9 2 9 2 1 11 11 11 11 13 3 1 2 11 11 2 16 1 11 13 1 9 2 11 2 2
16 11 13 10 9 1 9 11 11 2 11 11 2 11 11 11 2
23 9 9 11 2 11 11 2 3 13 1 10 9 1 11 7 3 0 1 9 9 9 9 2
11 11 11 2 2 13 10 10 9 9 11 2
24 13 11 11 2 9 12 11 13 1 9 12 11 2 16 9 9 11 2 7 11 13 9 11 2
9 9 11 2 9 11 13 11 3 2
18 10 9 1 11 7 9 2 9 13 1 9 2 15 3 13 9 9 2
33 11 11 11 2 13 10 10 9 11 11 11 15 13 1 11 11 11 2 15 13 1 11 2 11 2 11 11 11 9 11 2 11 2
6 3 11 3 13 13 2
73 1 9 11 2 11 11 11 11 9 2 9 10 3 13 10 9 9 11 1 9 2 11 11 11 11 2 2 9 1 2 11 11 2 11 11 2 11 2 2 9 9 13 1 2 11 11 11 2 2 11 1 2 11 11 11 2 2 9 1 2 11 11 11 11 11 2 11 2 7 3 9 3 2
38 9 0 3 3 13 1 10 9 1 9 9 1 9 9 0 2 9 11 2 2 7 1 9 1 12 9 9 2 9 9 9 2 11 2 11 11 2 2
21 11 11 13 1 9 9 9 9 7 13 9 9 12 5 2 7 13 9 9 9 2
24 11 0 11 12 13 9 1 11 15 13 9 7 9 9 11 2 1 9 1 9 9 9 12 2
10 10 12 5 11 13 1 1 9 9 2
15 7 2 9 10 3 13 11 11 15 3 13 9 13 13 2
13 13 13 1 12 1 12 12 9 9 11 1 9 2
9 15 13 10 9 7 12 10 9 2
13 11 13 3 13 12 9 11 7 11 13 10 9 2
15 10 9 13 11 11 2 16 13 3 3 9 11 1 9 2
13 9 15 3 13 0 1 11 2 3 13 13 15 2
30 1 9 7 9 0 2 11 0 1 9 9 11 2 9 2 9 9 2 9 11 2 7 9 9 9 2 9 0 11 2
37 16 7 7 2 11 13 11 11 13 1 9 11 2 7 10 9 2 11 3 13 13 1 9 11 15 3 2 3 0 10 16 3 10 13 9 11 2
18 11 13 9 7 13 2 2 1 9 13 9 1 9 15 14 13 9 2
15 3 9 10 13 1 9 0 2 3 1 9 11 1 11 2
4 9 9 9 2
10 10 11 13 1 12 1 11 11 11 2
43 1 9 2 11 11 11 11 2 2 12 2 2 1 9 9 2 10 9 0 15 9 10 13 0 2 0 12 9 1 9 2 3 13 9 9 9 15 13 12 9 1 9 2
27 9 10 13 1 11 11 2 7 13 11 11 2 11 2 11 2 11 11 2 11 2 11 11 2 7 11 2
19 10 3 9 9 2 9 9 2 7 9 2 9 0 15 13 11 2 11 2
23 9 15 13 1 11 11 1 2 11 11 1 9 11 1 2 11 2 11 11 7 11 11 2
19 2 11 11 2 3 15 13 9 15 11 13 9 2 15 13 9 9 9 2
22 9 9 11 15 3 13 10 9 13 9 9 9 15 0 13 9 7 9 0 1 9 2
37 16 2 9 0 11 11 15 13 9 11 11 2 11 11 9 11 11 2 13 13 9 1 13 11 11 7 11 11 16 3 13 9 0 1 11 11 2
5 15 9 9 10 2
16 11 13 9 15 13 1 9 11 2 11 11 2 11 2 11 2
38 11 11 2 9 11 2 11 11 11 2 11 2 2 13 1 9 11 12 1 13 11 11 11 15 3 13 1 9 0 1 9 11 11 1 15 11 11 2
14 9 13 9 1 9 9 15 0 7 9 0 15 13 2
12 9 10 13 11 2 11 2 11 11 11 2 2
7 15 13 9 0 11 11 2
33 9 9 11 13 9 15 13 9 2 9 15 13 9 1 10 9 9 1 9 3 13 2 12 1 1 3 13 0 13 9 9 3 2
28 13 10 9 3 14 0 2 16 15 13 16 11 1 9 15 0 3 13 9 10 9 9 1 13 9 1 9 2
28 10 10 9 13 9 9 16 9 9 3 13 13 1 9 12 2 9 11 11 3 13 9 16 9 0 3 13 2
16 9 11 2 11 7 11 13 1 9 11 11 11 1 9 12 2
24 16 9 11 3 13 2 15 3 13 1 9 9 1 13 9 9 9 9 11 1 11 11 11 2
25 1 9 15 3 0 2 11 3 13 9 2 11 2 13 9 0 2 0 1 15 1 9 9 9 2
16 9 0 13 9 1 9 11 1 13 9 7 13 9 9 9 2
8 9 10 13 1 9 11 11 2
23 11 13 10 10 9 15 13 1 11 11 11 2 9 11 11 2 11 11 11 11 2 11 2
19 16 13 1 11 11 2 11 13 9 15 1 11 11 9 9 1 9 12 2
18 11 13 9 9 15 13 9 0 7 3 13 9 7 3 13 1 0 2
23 1 9 11 1 15 3 13 3 0 16 15 13 2 16 13 3 2 3 3 3 13 9 2
12 3 9 9 10 9 15 3 1 9 9 10 2
10 3 14 13 0 10 3 13 13 11 2
17 9 9 9 11 13 1 11 2 11 2 11 2 11 11 2 11 2
18 9 10 13 9 1 13 2 13 2 7 13 9 2 9 9 9 0 2
33 9 12 2 11 7 9 11 2 12 2 13 1 9 13 2 16 3 15 13 9 13 9 15 0 2 15 9 1 9 15 0 13 2
29 1 11 11 12 2 1 9 9 12 2 12 9 9 1 11 11 2 10 9 1 9 9 13 11 11 1 13 11 2
25 1 9 12 2 11 13 9 1 12 9 9 1 11 11 2 9 11 2 9 9 11 2 11 2 2
39 1 9 12 2 3 11 11 12 15 13 11 11 11 11 11 11 11 11 11 11 2 9 9 12 2 2 15 13 1 9 9 9 15 13 1 11 11 3 2
11 3 0 9 13 9 1 9 11 7 11 2
18 1 12 1 12 2 15 13 1 9 2 9 9 11 2 11 1 11 2
26 12 2 1 9 0 15 13 9 11 2 9 9 2 15 13 9 2 13 1 9 2 15 13 9 0 2
16 11 11 11 11 13 9 9 9 15 0 1 11 1 9 12 2
23 9 10 13 1 9 9 15 3 13 10 10 9 9 15 13 7 13 9 1 9 9 9 2
17 11 2 2 13 11 11 11 1 9 12 1 12 7 12 1 12 2
5 16 2 15 9 2
36 11 9 9 1 13 1 9 10 13 1 9 1 13 9 9 2 3 16 9 0 10 13 1 9 0 15 3 2 3 3 13 9 2 9 2 2
8 3 15 3 13 2 11 2 2
35 11 11 12 11 13 1 9 9 9 12 11 2 3 13 1 11 11 12 11 2 2 16 9 14 13 16 9 13 1 9 1 11 11 11 2
19 16 11 13 9 11 1 9 12 7 13 3 1 9 12 2 12 7 12 2
10 9 13 11 13 1 11 10 9 11 2
16 11 10 3 13 12 9 7 9 9 2 7 12 9 9 9 2
10 11 1 9 9 10 13 9 9 9 2
9 3 15 3 13 9 7 9 9 2
36 13 11 2 7 3 13 9 1 10 9 11 11 2 14 13 16 11 3 3 13 9 2 11 3 9 1 11 11 2 9 15 12 10 3 0 2
20 11 13 9 1 9 11 2 11 11 11 2 11 1 11 2 11 2 11 11 2
24 1 13 9 15 3 0 1 9 11 12 11 2 16 3 13 10 9 9 7 9 15 3 13 2
35 1 9 11 2 9 11 13 1 12 2 12 2 3 1 9 15 0 2 1 13 9 2 9 7 9 2 9 15 13 11 11 7 9 9 2
19 1 9 11 3 13 1 9 2 7 3 13 9 9 9 0 1 9 9 2
17 15 13 9 1 10 9 13 11 7 1 10 9 10 0 7 0 2
18 9 0 3 13 9 9 9 2 9 2 7 13 9 3 9 9 9 2
14 9 15 3 13 1 9 9 10 13 1 9 15 13 2
27 11 13 1 9 1 9 0 2 11 11 2 11 11 2 2 7 10 9 0 13 11 11 2 11 11 2 2
8 1 9 9 13 13 9 9 2
14 13 16 9 1 9 9 13 9 9 2 14 9 9 2
14 1 11 3 13 9 11 15 13 1 9 1 9 12 2
19 2 9 15 3 13 9 1 11 2 11 3 13 9 1 9 1 10 9 2
4 11 3 13 2
17 1 9 9 3 13 1 11 1 9 11 11 16 11 11 13 9 2
22 15 13 9 0 1 9 9 12 11 2 11 12 2 7 16 15 13 0 1 11 11 2
14 1 9 11 3 13 1 9 9 16 15 7 9 13 2
17 3 2 3 13 9 9 7 9 1 9 1 13 11 1 1 9 2
66 2 5 2 2 11 12 2 13 9 0 15 13 3 12 9 2 2 11 2 11 2 11 12 2 13 9 12 15 3 13 12 1 9 2 7 11 2 11 12 2 13 9 12 15 3 13 12 1 11 2 11 3 13 9 1 12 9 9 7 13 10 10 9 11 0 2
48 3 9 11 11 2 15 13 11 2 1 9 11 2 12 2 7 9 9 11 11 2 1 9 12 2 15 13 1 9 11 2 1 9 15 13 3 2 3 11 11 2 11 11 2 7 11 11 2
13 9 13 9 9 15 13 3 13 0 9 9 0 2
14 10 9 15 13 3 1 12 9 3 13 1 10 9 2
14 11 15 13 9 9 9 13 3 1 9 2 0 9 2
39 1 11 11 13 1 11 9 12 11 12 9 12 2 12 11 12 11 11 2 2 9 9 9 13 1 3 1 13 9 9 0 13 9 11 15 13 9 12 2
19 10 9 0 1 9 11 11 2 11 11 2 11 2 11 11 7 11 11 2
22 9 10 13 1 11 7 13 1 9 12 1 9 12 1 10 9 1 11 12 9 9 2
28 1 9 1 9 2 11 13 16 3 9 11 15 13 1 9 9 9 7 9 10 3 13 1 9 13 9 11 2
24 16 9 11 13 13 1 9 0 2 11 13 1 9 1 9 11 9 11 2 11 2 1 11 2
7 2 0 15 3 9 11 2
23 1 9 9 2 11 13 16 9 12 15 13 2 0 2 13 9 15 13 2 9 9 2 2
19 11 13 9 1 13 9 9 9 7 11 9 13 2 13 11 13 1 11 2
46 11 10 13 9 0 1 9 10 7 9 5 9 9 0 10 2 16 1 9 0 3 13 10 9 15 0 3 13 9 9 15 13 13 9 1 13 9 1 9 1 9 9 3 13 9 2
14 9 11 2 11 13 1 2 11 2 11 11 11 11 2
17 9 11 1 9 0 12 11 12 1 9 0 13 9 11 15 0 2
13 3 13 1 9 15 13 9 9 0 1 9 9 2
62 11 13 1 9 11 1 9 9 11 1 11 1 9 2 7 13 2 9 9 11 1 11 2 11 2 11 2 1 9 11 1 11 11 1 11 11 12 1 9 12 11 12 2 9 11 11 11 13 2 11 11 11 11 2 2 11 11 11 2 11 2 2
8 15 15 0 13 9 9 10 2
17 1 9 9 9 9 2 11 3 13 16 9 13 1 9 0 10 2
15 9 9 10 13 1 9 11 11 2 15 13 2 0 2 2
24 11 0 9 7 11 11 13 9 15 13 13 9 9 0 16 13 2 13 7 13 1 1 9 2
79 1 9 11 15 13 11 11 11 13 16 9 11 2 11 2 11 9 12 13 9 0 1 11 15 9 10 1 9 9 11 11 11 2 9 0 10 13 9 1 9 11 2 11 9 11 2 11 2 11 2 7 9 1 11 9 15 13 9 9 11 2 11 2 11 2 7 13 3 12 9 9 2 9 2 7 12 9 9 2
22 9 10 13 16 9 9 1 10 9 13 2 10 9 3 13 13 10 9 9 15 0 2
13 9 3 0 0 1 9 0 13 7 9 0 0 2
39 11 11 13 1 12 9 0 2 11 11 7 11 11 2 7 11 13 0 1 9 11 2 15 13 9 15 1 2 11 2 11 2 13 2 0 7 0 2 2
27 11 13 9 9 2 2 9 9 2 2 1 9 7 13 9 9 11 1 11 11 11 1 9 12 1 12 2
33 16 13 10 9 15 13 9 2 13 15 1 15 2 2 3 15 13 9 15 3 2 16 13 1 10 9 10 1 9 15 0 10 2
23 9 10 3 13 9 9 1 9 0 10 2 1 11 2 11 11 11 2 2 11 7 11 2
11 9 10 13 9 9 9 0 13 9 11 2
13 11 13 9 0 1 9 11 11 11 2 11 2 2
37 11 13 11 1 11 11 11 1 9 12 9 12 1 10 9 0 0 2 15 0 1 11 1 9 12 7 12 0 1 9 9 1 10 9 1 12 2
29 1 9 12 2 9 9 12 1 11 2 11 2 11 7 11 1 11 13 9 13 1 9 11 11 11 1 9 12 2
22 9 12 2 9 3 13 9 7 9 1 9 9 13 9 1 9 9 1 9 15 0 2
17 10 9 9 9 13 3 13 9 0 1 13 0 9 15 3 13 2
9 2 1 9 15 13 1 9 9 2
32 1 11 11 13 13 11 11 1 9 12 11 12 2 9 10 13 1 10 9 0 1 11 13 11 11 11 11 1 12 11 12 2
17 11 11 3 13 1 9 9 0 13 1 9 15 13 0 7 0 2
10 9 9 13 7 9 9 13 1 9 2
23 11 11 2 11 13 10 10 9 1 9 11 11 2 11 11 11 2 11 11 11 2 11 2
10 16 11 0 2 9 15 3 13 15 2
19 11 11 11 10 15 13 11 7 9 11 11 13 3 0 1 9 12 10 2
15 1 10 1 9 9 13 10 9 13 9 1 0 2 0 2
15 9 10 13 9 9 15 0 2 3 13 1 9 11 11 2
15 1 9 12 2 1 11 11 2 9 9 9 13 1 11 2
9 10 9 1 12 11 12 1 11 2
14 15 3 13 10 9 15 1 10 13 13 3 11 11 2
17 9 15 13 1 9 0 2 13 3 9 7 9 2 13 1 9 2
15 11 3 13 1 9 15 0 2 16 3 13 9 15 0 2
41 1 0 2 9 9 13 9 2 10 3 10 9 7 9 1 9 9 13 1 13 7 14 13 2 3 10 10 9 7 9 3 13 13 10 9 15 13 1 9 9 2
37 16 9 14 2 11 14 13 1 1 9 9 2 3 1 9 2 9 0 13 1 9 14 2 11 2 9 13 9 11 15 3 13 1 13 9 10 2
19 9 10 13 9 9 10 3 13 9 9 11 11 7 13 9 13 9 0 2
6 9 13 2 11 2 2
14 1 9 0 3 13 11 11 13 10 10 9 0 9 2
48 9 11 13 9 1 12 9 15 0 2 1 9 9 9 0 13 9 0 2 15 10 1 1 13 9 1 9 12 9 1 9 9 9 2 9 9 2 9 1 9 0 0 2 0 7 0 2 2
25 1 12 9 12 9 2 9 9 9 9 2 2 11 2 13 1 9 9 0 11 7 10 9 9 2
23 15 13 1 1 12 9 1 9 12 2 12 2 7 13 1 11 11 11 11 1 9 12 2
19 11 13 10 9 15 13 1 9 11 11 2 11 11 2 11 11 2 11 2
54 9 2 9 15 13 1 9 11 13 2 9 2 9 11 15 13 1 11 13 2 9 2 9 11 15 13 1 11 1 9 12 2 9 10 13 1 12 9 3 9 11 15 13 1 11 7 9 11 15 14 13 1 11 2
11 11 2 9 15 13 9 9 11 13 9 2
6 9 15 14 13 3 2
52 9 15 3 0 15 13 1 10 9 9 9 9 10 13 11 11 15 1 9 12 13 1 13 1 3 13 16 9 9 13 9 2 13 1 9 2 2 10 9 15 13 1 11 11 15 9 0 13 3 10 9 2
43 11 13 13 12 9 12 1 9 9 2 12 11 7 12 11 11 2 10 9 1 9 12 15 13 1 9 11 11 13 1 9 10 9 1 9 9 2 16 14 13 1 9 2
19 11 11 13 10 9 15 13 1 9 11 11 2 11 11 2 11 2 11 2
45 9 10 3 13 1 10 9 3 2 7 16 9 9 11 11 11 3 13 1 9 11 7 9 11 11 11 2 11 11 11 11 11 11 13 13 11 7 3 3 13 9 1 13 11 2
49 9 9 2 12 1 12 9 2 13 12 9 0 11 11 2 3 13 16 15 14 3 13 11 2 11 9 1 11 5 11 1 9 11 13 1 9 1 12 9 7 12 9 13 12 9 7 12 9 2
23 1 9 11 11 2 11 11 11 13 9 9 11 11 11 2 11 10 3 13 9 9 9 2
21 7 9 2 11 11 2 1 11 2 1 11 2 14 9 7 9 11 3 13 0 2
18 9 10 0 7 3 0 16 15 3 0 13 9 9 9 2 2 9 2
20 3 14 15 1 13 3 9 15 3 15 13 10 13 11 2 1 9 0 0 2
12 16 1 15 11 3 13 9 2 11 7 11 2
11 9 10 13 1 9 11 11 1 10 11 2
12 1 9 11 12 2 13 10 9 1 9 10 2
13 11 3 13 9 1 9 11 11 1 12 11 12 2
11 3 11 2 11 11 7 11 3 13 11 2
28 11 13 9 9 15 13 1 9 9 11 9 9 2 9 2 2 16 1 11 9 10 3 13 9 2 9 2 2
18 11 11 11 13 9 9 9 11 2 11 11 2 15 13 1 9 12 2
33 1 11 2 9 15 13 9 2 9 10 13 11 11 11 7 11 1 9 9 9 9 7 9 11 11 11 11 1 9 9 7 9 2
30 11 13 1 10 9 16 3 13 9 9 15 13 0 15 9 15 13 9 13 7 3 13 1 9 15 13 9 2 9 2
41 3 13 12 9 0 1 9 10 2 16 2 11 7 11 2 2 2 15 15 11 2 2 7 2 11 11 2 2 16 12 9 13 9 2 9 15 15 3 13 9 2
7 9 10 13 1 9 12 2
11 11 2 11 2 11 13 9 9 1 11 2
6 3 11 13 1 9 2
23 16 15 13 13 9 1 9 13 1 1 9 1 13 9 11 2 11 13 13 10 1 9 2
12 9 0 9 10 13 2 9 11 7 11 11 2
29 11 11 11 11 13 9 9 9 11 15 13 1 11 11 7 13 1 11 11 2 11 11 2 11 11 7 11 11 2
6 13 9 1 11 11 2
27 9 11 11 11 11 11 3 13 10 9 7 9 2 9 9 11 11 11 11 15 9 3 13 9 2 12 2
31 1 9 0 13 9 9 1 9 13 9 9 0 1 9 12 7 12 2 9 10 13 16 11 13 1 9 1 13 9 10 2
45 11 2 11 13 0 1 9 9 11 2 1 0 9 11 2 11 13 1 9 11 2 11 11 2 7 11 2 13 10 9 1 9 2 9 15 10 0 9 13 11 1 11 7 11 2
14 11 13 16 9 11 15 3 13 3 3 3 13 9 2
21 13 11 11 2 11 13 9 9 2 9 12 9 9 2 11 2 7 2 11 2 2
16 10 10 15 0 13 9 11 15 13 1 9 11 7 11 13 2
20 11 9 10 13 1 9 12 2 12 2 7 1 13 1 11 2 7 11 2 2
26 15 0 13 9 9 2 2 10 9 13 1 9 10 1 9 9 2 9 2 2 1 9 15 13 9 2
21 9 15 3 0 1 11 1 10 9 9 11 11 2 11 3 13 11 1 13 9 2
32 3 11 11 13 1 9 1 10 3 13 0 7 10 1 9 3 13 2 9 10 13 9 9 11 1 9 7 9 2 9 0 2
33 1 15 9 13 1 3 13 9 10 9 2 11 3 13 9 9 0 1 10 9 1 9 2 15 10 10 9 13 9 9 9 11 2
10 11 2 11 2 13 9 9 1 11 2
12 11 11 3 8 13 9 7 9 13 9 9 2
17 11 13 9 15 13 1 11 11 7 11 11 2 15 13 1 12 2
37 1 9 12 2 12 11 1 11 1 12 11 2 11 13 12 9 2 13 11 13 12 9 0 3 2 3 7 9 12 9 1 11 11 1 9 12 2
24 1 12 2 11 11 11 11 13 12 13 0 7 12 13 0 2 13 9 9 9 1 12 9 2
22 1 7 10 2 16 9 15 3 13 1 13 9 7 9 2 14 0 3 13 1 9 2
19 9 10 13 1 9 12 7 13 1 11 2 11 11 11 7 11 11 11 2
19 11 11 13 10 9 0 0 11 15 13 13 1 13 9 1 10 9 0 2
18 11 11 13 9 9 15 3 13 9 9 9 11 11 11 1 9 12 2
16 11 2 11 11 11 11 2 2 13 11 11 1 11 11 11 2
14 11 11 13 9 0 2 1 13 9 12 11 5 9 2
21 11 10 3 13 1 0 7 9 15 0 13 11 11 2 15 3 13 9 9 11 2
11 3 2 0 9 10 0 7 14 13 9 2
27 9 9 10 1 11 11 2 3 11 2 16 10 9 13 10 13 13 11 2 9 12 13 9 9 1 11 2
15 10 2 10 9 9 15 13 13 9 9 7 9 15 0 2
13 11 14 13 9 0 10 9 0 15 13 9 0 2
14 11 13 9 1 9 11 2 11 2 11 11 2 11 2
15 9 9 16 0 0 0 2 7 1 9 0 0 1 9 2
24 11 11 16 13 9 0 1 11 2 15 13 1 9 9 11 11 13 1 9 15 9 2 11 2
15 9 10 13 12 1 12 9 7 9 15 13 1 11 11 2
47 5 11 11 7 11 11 5 11 11 11 5 11 11 11 5 11 11 7 11 11 5 11 11 5 11 11 5 11 11 5 11 11 5 11 11 7 11 11 11 5 11 11 7 11 11 11 11
11 11 2 9 10 14 3 13 9 9 11 2
15 7 11 11 11 1 9 9 11 11 7 13 9 1 11 2
22 11 14 13 9 9 1 11 7 3 13 2 13 1 10 10 9 11 15 13 1 11 2
12 3 11 2 11 7 11 13 9 9 0 10 2
24 11 11 2 11 11 2 13 9 1 9 11 15 13 1 13 9 3 9 15 3 13 9 0 2
11 9 9 13 9 1 9 9 0 1 9 2
22 1 9 0 1 10 9 9 9 11 2 11 11 11 11 13 13 10 10 9 9 0 2
16 11 3 13 9 9 1 11 2 9 1 13 1 9 9 3 2
20 11 11 13 1 9 1 9 11 11 11 11 11 11 7 13 1 12 9 9 2
12 9 10 3 13 1 9 2 9 2 7 9 2
27 9 9 10 3 13 1 9 2 7 3 13 9 10 3 1 9 2 9 0 2 13 1 11 11 2 11 2
29 11 2 11 2 11 11 2 3 13 9 9 9 9 10 7 13 9 9 13 7 9 9 11 11 2 11 11 2 2
14 1 9 2 11 2 11 2 1 0 13 9 7 9 2
30 1 9 12 2 11 11 11 7 11 11 11 13 13 12 7 13 11 11 11 7 11 11 11 13 9 13 11 11 11 2
11 16 9 13 2 9 1 13 0 3 0 2
34 9 9 2 9 9 9 1 11 11 11 11 7 9 0 1 11 11 1 11 15 13 1 11 2 11 2 13 1 13 9 1 9 10 2
11 0 15 13 1 9 11 13 11 2 11 2
33 1 0 9 9 2 1 9 12 2 3 13 13 12 9 11 7 13 9 9 9 9 9 9 0 11 2 11 11 11 2 11 2 2
9 9 9 3 13 16 13 11 11 2
35 9 1 9 15 13 11 11 11 3 13 1 9 13 2 7 9 13 16 9 10 3 13 1 9 9 15 9 13 1 9 0 15 13 0 2
20 9 10 13 9 0 1 9 11 7 11 16 3 13 9 9 9 7 9 11 2
6 11 13 1 9 0 2
10 3 15 13 1 9 11 1 12 2 2
10 15 3 0 7 0 2 0 1 11 2
28 9 9 11 11 11 9 10 13 9 9 12 9 15 13 9 11 2 11 2 7 11 11 2 11 1 11 2 2
22 11 2 11 13 1 11 11 1 9 2 9 11 7 11 1 9 2 7 11 11 11 11
21 3 13 3 9 15 14 13 9 7 7 13 1 15 1 9 15 7 9 15 13 2
14 11 13 9 1 9 11 2 11 2 11 11 2 11 2
19 11 10 13 1 9 2 9 2 9 2 9 9 2 9 2 9 7 9 2
5 13 1 11 11 2
36 1 9 9 12 2 12 2 11 12 3 13 9 9 13 12 15 13 1 11 11 11 11 11 2 12 11 11 13 1 11 7 9 11 11 11 2
23 16 9 0 15 13 1 9 1 9 9 7 9 9 2 16 9 10 9 3 3 13 0 2
24 9 0 15 2 11 11 11 11 11 13 1 9 12 14 0 16 13 9 1 9 11 11 11 2
28 9 10 13 1 11 11 2 10 9 9 11 2 1 9 12 2 1 10 9 1 11 2 9 12 7 12 2 2
10 3 14 9 0 10 3 13 13 9 2
35 1 12 1 11 2 11 11 11 13 7 13 9 1 10 9 7 9 15 3 13 9 2 9 0 2 11 11 2 11 2 12 2 12 2 2
18 11 11 2 2 13 10 11 1 9 9 11 1 11 2 11 2 11 2
13 3 1 9 12 2 9 11 13 1 9 11 11 2
25 11 9 10 13 9 9 11 15 0 7 0 1 9 11 2 11 1 9 2 9 7 9 2 9 2
18 1 10 2 9 1 9 13 1 9 15 3 13 1 9 9 9 13 2
25 1 1 11 2 11 3 13 9 0 16 13 1 9 11 11 1 11 11 7 11 11 1 9 11 2
7 9 15 3 13 9 10 2
77 3 1 9 11 2 16 9 11 1 11 11 13 9 2 16 11 11 11 10 13 1 11 11 15 13 9 9 1 11 11 1 9 10 13 9 9 13 11 2 11 11 2 2 9 9 2 11 5 11 11 2 7 11 2 11 2 2 11 11 2 11 11 2 15 13 1 9 9 9 11 11 11 11 2 11 2 2
14 1 9 9 2 9 9 13 9 1 9 9 15 0 2
21 1 9 9 9 13 11 13 9 13 9 13 12 1 9 11 11 1 1 2 1 2
18 16 9 13 1 11 7 11 7 3 2 3 13 0 1 9 11 11 2
21 9 9 3 13 9 9 15 13 9 2 11 7 13 9 2 9 0 0 1 9 2
12 11 11 13 9 9 1 11 15 13 9 9 2
10 11 9 9 9 3 3 13 13 9 2
17 11 11 2 11 11 2 7 11 11 13 9 0 1 9 11 11 2
11 9 0 9 1 9 9 0 11 1 11 2
14 11 11 13 9 1 9 10 2 16 13 1 9 10 2
6 15 13 9 13 11 2
15 15 3 13 1 9 2 11 2 16 15 13 10 9 0 2
5 11 0 13 9 2
15 1 10 9 11 13 2 2 3 15 14 13 9 9 10 2
12 13 9 11 2 11 13 10 9 11 11 11 2
16 11 11 13 9 11 15 13 1 9 12 1 13 1 11 11 2
9 14 3 13 9 2 14 0 13 2
24 16 13 12 9 12 1 9 2 1 9 12 2 11 11 13 9 2 11 11 11 2 1 11 2
11 1 9 12 2 11 13 9 1 12 9 2
13 11 13 1 9 11 2 9 2 9 2 9 2 2
10 9 9 13 1 9 11 2 12 2 2
6 11 10 13 9 12 2
22 9 0 13 9 2 9 15 9 13 1 11 11 11 2 7 15 13 9 1 11 11 2
43 11 11 11 13 10 10 9 15 13 1 11 15 3 0 10 13 13 13 11 11 12 11 2 3 13 9 7 9 15 13 3 13 9 9 13 13 2 15 13 1 9 11 2
55 11 3 13 11 2 11 2 11 1 9 2 9 11 11 0 1 11 2 1 11 11 11 11 12 2 11 11 11 11 11 7 11 11 11 11 1 11 2 14 13 3 3 9 9 0 1 11 2 3 11 11 11 11 11 2
22 9 11 13 1 9 0 16 9 12 11 12 2 1 9 11 11 9 12 13 1 1 2
15 15 13 10 9 2 11 11 2 7 10 11 2 11 11 2
71 9 2 12 2 15 0 16 2 16 11 3 0 2 12 2 13 9 0 10 3 1 9 2 2 12 2 13 1 15 0 2 2 9 15 3 15 13 1 9 15 2 2 12 2 15 3 15 13 1 9 15 7 1 9 15 2 12 2 15 3 15 13 2 9 15 15 13 1 15 2 2
14 11 2 11 11 2 2 13 9 9 9 9 13 11 2
18 11 13 9 9 0 1 9 11 7 10 10 1 9 9 0 1 11 2
8 9 10 15 13 1 9 9 2
13 9 10 3 13 1 9 9 2 9 1 9 11 2
7 9 11 11 2 2 11 2
17 11 11 13 9 1 11 11 2 11 11 2 11 11 11 2 11 2
6 15 9 13 3 0 2
31 16 1 9 9 12 2 12 2 9 9 1 11 9 9 14 13 9 9 9 11 2 11 9 13 1 11 1 0 9 12 2
16 9 9 10 13 1 12 9 12 7 13 9 1 12 11 12 2
32 12 2 3 13 1 13 9 0 10 1 12 9 9 15 3 13 2 1 9 7 9 9 2 9 2 9 2 7 0 9 2 2
20 12 12 9 3 2 12 9 11 13 13 3 11 2 11 2 7 11 2 11 2
13 11 9 12 9 1 9 13 9 1 9 9 9 2
19 11 11 11 11 13 1 12 5 9 9 11 2 11 11 11 1 9 9 2
15 9 9 0 1 9 10 13 9 2 9 7 9 2 9 2
20 11 13 11 7 13 13 9 9 1 3 2 3 2 13 9 15 0 1 3 2
12 11 13 9 15 13 1 11 11 11 2 11 2
12 10 9 9 1 9 15 13 2 11 11 2 2
66 9 0 13 16 14 13 7 14 13 9 2 2 9 9 2 7 2 15 13 2 2 16 9 10 2 11 3 3 13 2 2 2 16 1 9 1 9 11 9 11 7 15 13 10 13 7 13 9 1 11 2 14 3 2 0 1 11 11 2 16 15 13 3 1 11 2
29 1 1 2 13 11 15 13 13 11 11 11 2 15 1 9 12 13 11 11 11 2 2 16 9 3 13 1 11 2
14 11 13 9 1 9 11 2 11 2 11 11 2 11 2
22 9 10 1 9 13 1 10 9 0 16 9 9 13 1 9 9 2 9 10 13 3 2
19 9 1 0 11 11 2 11 11 2 11 11 2 11 11 2 7 11 11 2
19 1 9 12 9 11 12 1 12 9 1 12 9 13 15 0 1 9 12 2
36 11 11 15 13 9 9 9 10 13 9 11 16 9 9 2 1 0 11 11 2 9 1 9 11 11 2 2 9 11 11 11 7 0 2 0 2
34 1 9 0 2 12 11 12 2 11 1 12 3 13 1 9 1 9 9 11 5 11 11 1 11 11 11 2 7 13 2 11 11 2 2
32 11 9 9 3 3 13 1 9 9 9 3 2 9 10 13 16 14 3 9 1 9 13 9 15 13 3 1 9 9 9 9 2
13 11 11 11 3 13 9 0 1 9 11 11 11 2
27 9 15 3 13 13 11 15 13 12 9 2 13 11 11 7 11 2 12 2 2 7 11 11 2 12 2 2
7 11 2 11 11 2 11 11
17 16 3 11 13 9 15 1 10 3 13 9 9 13 9 9 0 2
21 0 9 7 9 13 11 9 11 9 1 10 9 2 7 3 13 10 9 1 9 2
6 11 13 9 9 9 2
14 2 9 0 15 3 3 13 12 9 10 2 2 13 2
23 15 13 13 9 9 15 0 7 9 15 0 2 9 3 13 1 0 11 1 11 11 11 2
24 11 11 11 11 2 11 11 2 11 11 11 2 3 13 11 2 13 9 9 11 9 1 11 2
15 7 16 2 11 2 10 9 11 2 13 9 2 9 10 2
8 0 10 14 9 1 11 11 2
23 11 11 13 11 11 2 11 2 11 2 7 11 2 2 9 11 15 13 9 1 11 11 2
10 13 14 13 2 15 11 13 9 3 2
41 11 9 13 9 9 3 2 11 2 13 9 9 2 2 13 9 9 2 9 9 2 9 9 2 2 11 2 0 2 2 9 2 9 9 2 2 7 13 9 9 2
15 15 13 1 11 1 9 12 11 12 2 13 9 11 12 2
26 11 13 9 10 1 9 15 0 2 1 10 9 13 1 13 9 0 2 15 13 3 13 9 10 9 2
23 9 9 13 1 1 9 9 1 12 9 9 11 1 9 11 12 16 9 15 0 9 11 2
15 1 9 13 2 11 11 3 13 11 11 9 2 11 2 2
4 9 1 11 2
4 13 1 9 2
26 15 14 9 1 9 2 9 7 9 9 11 15 12 9 2 16 15 13 9 2 9 1 9 9 10 2
12 1 11 2 9 1 9 13 1 1 9 0 2
22 9 11 3 13 11 11 13 3 0 1 9 1 9 0 1 9 11 7 9 9 9 2
19 11 12 3 13 9 11 13 9 9 0 15 14 13 9 1 13 9 1 2
29 11 1 9 11 11 13 1 12 9 1 11 7 11 1 12 11 12 1 12 2 12 7 13 9 1 9 9 9 2
3 11 12 2
21 15 13 9 1 9 7 9 1 9 2 9 1 13 10 9 1 1 9 9 13 2
41 9 2 9 9 12 2 8 2 11 11 3 13 1 11 11 1 11 1 11 11 12 9 2 11 11 2 8 2 9 9 12 1 9 9 1 9 2 12 9 12 2
22 11 11 11 7 3 13 1 9 11 11 2 12 11 12 2 13 10 9 9 13 11 2
20 12 2 1 9 10 9 9 1 11 11 11 2 16 11 11 1 9 13 0 2
13 11 13 10 9 1 11 11 2 11 11 2 11 2
18 11 1 11 3 13 1 9 15 7 13 11 1 9 1 9 12 9 2
11 13 9 1 9 0 1 11 7 9 0 2
24 11 13 16 11 13 1 9 11 2 1 9 11 13 9 0 13 9 7 13 1 11 7 9 2
48 11 13 9 11 15 11 7 13 10 9 1 13 9 15 1 13 9 3 0 1 9 1 11 10 2 11 3 13 9 12 9 3 1 9 9 11 1 11 7 11 2 13 2 7 3 13 11 2
15 11 2 11 2 2 13 9 9 9 11 15 13 1 11 2
5 9 3 9 10 2
41 11 13 9 7 9 9 16 15 13 1 0 7 0 3 13 10 9 9 9 2 15 13 3 13 13 9 9 0 15 3 13 16 15 3 13 9 9 7 9 9 2
27 16 11 7 9 2 9 13 16 11 13 1 9 10 2 15 3 13 16 11 3 13 9 10 1 15 0 2
13 3 15 3 3 13 9 1 11 2 7 13 9 2
24 3 12 9 3 2 1 12 11 2 11 13 12 9 1 9 12 2 12 1 0 9 13 11 2
34 16 3 13 1 11 2 11 11 11 3 13 9 0 9 7 9 13 11 11 1 11 2 11 2 9 9 1 11 11 15 3 9 11 2
33 11 3 13 7 13 9 9 15 9 1 10 9 13 15 13 1 11 7 0 13 1 9 2 11 2 11 12 2 12 2 12 2 2
11 9 10 3 13 1 11 11 11 11 11 2
73 1 9 12 2 11 13 12 9 11 11 2 11 9 1 11 11 2 15 13 9 0 2 11 13 9 0 2 9 9 12 2 9 2 0 7 9 0 2 2 9 9 13 0 2 0 2 9 2 7 0 2 11 2 9 10 3 3 13 1 9 2 11 9 7 9 9 9 13 9 0 1 1 2
23 3 9 9 11 1 9 3 13 1 9 15 0 7 3 3 9 1 11 1 11 11 11 2
34 3 1 13 12 9 9 9 2 15 3 13 1 12 9 9 9 15 0 15 14 3 13 11 2 7 7 9 2 9 1 9 13 11 2
29 11 10 9 10 13 1 11 11 2 11 2 2 15 13 9 15 0 1 15 13 12 9 0 2 11 7 11 2 2
15 9 12 11 9 13 9 9 0 7 13 1 1 9 9 2
21 11 11 13 9 12 1 9 11 11 11 11 11 1 11 7 11 11 2 10 11 2
27 1 9 12 15 13 10 9 0 1 9 9 1 9 9 9 2 7 3 3 15 13 13 9 9 14 13 2
17 11 11 1 11 2 11 2 2 13 12 11 2 2 13 1 11 2
17 11 11 3 13 9 9 11 15 9 9 9 11 13 9 9 11 2
9 3 9 11 1 11 3 13 0 2
30 11 11 11 11 1 9 13 3 15 13 11 11 11 5 11 11 2 3 11 11 11 2 11 2 1 11 1 9 12 2
15 16 15 13 13 9 16 9 9 10 0 1 9 1 9 2
19 16 13 1 9 9 2 11 3 13 1 9 15 3 13 13 1 9 0 2
23 1 9 12 11 12 2 9 9 1 9 15 15 13 2 11 2 13 1 9 11 11 11 2
54 11 11 13 1 11 2 10 9 9 15 13 11 2 2 1 13 9 9 9 2 15 9 9 11 3 13 2 13 14 1 9 2 14 0 7 9 15 3 13 2 9 0 7 9 11 1 12 2 12 5 1 9 2 2
16 1 9 0 2 11 13 9 1 9 10 9 16 15 13 9 2
57 11 2 9 9 7 0 3 13 1 13 9 9 2 12 9 7 12 9 2 1 10 9 1 11 11 2 1 9 15 13 9 9 2 13 9 2 9 10 15 3 13 9 9 2 7 13 9 2 9 0 15 13 1 9 1 11 2
12 9 9 0 1 0 9 0 2 13 13 0 2
12 11 11 11 13 9 9 0 1 11 2 11 2
19 11 13 9 0 2 12 2 2 7 9 9 15 13 9 13 1 9 12 2
16 9 10 15 13 9 0 1 9 9 9 15 13 9 10 9 2
20 1 9 9 11 11 2 11 3 3 13 9 9 7 14 9 9 15 3 13 2
26 10 2 10 9 15 13 13 11 11 2 11 2 11 11 2 15 3 13 9 9 7 3 13 9 11 2
6 3 9 15 1 11 2
25 3 3 1 9 9 2 13 1 9 9 15 0 15 13 1 10 0 2 3 11 15 13 1 0 2
7 9 13 3 3 12 9 2
38 1 9 11 2 9 2 11 2 11 2 11 2 11 2 7 11 2 9 2 3 13 1 9 2 9 0 15 0 2 15 13 1 9 9 1 9 9 2
16 9 9 1 9 10 13 2 15 15 13 15 13 9 10 2 2
19 11 11 11 13 2 11 2 15 13 2 11 11 2 15 13 1 9 11 2
14 15 14 9 9 3 3 13 9 9 9 2 9 11 2
21 1 9 10 2 9 1 9 9 3 14 3 0 7 9 3 13 1 9 9 0 2
20 16 3 2 15 3 13 1 10 9 9 1 11 11 15 13 9 11 1 11 2
41 11 13 9 9 1 11 11 11 11 1 9 1 11 2 10 9 15 1 10 13 1 10 9 9 2 16 15 13 1 13 1 9 13 1 0 7 14 13 1 9 2
15 1 10 2 0 13 11 11 1 11 11 9 12 2 12 2
14 9 10 13 1 9 11 7 3 13 1 10 9 11 2
19 1 9 9 12 2 12 2 11 3 3 13 9 11 1 9 9 2 9 2
8 9 1 9 9 12 5 12 2
12 9 10 13 1 11 11 1 9 9 11 11 2
10 9 3 13 14 3 0 1 11 11 2
29 11 3 13 3 1 15 13 7 3 9 11 3 13 9 9 11 2 15 14 3 13 3 1 9 9 11 3 0 2
32 13 0 9 2 11 8 13 13 15 10 9 2 10 9 9 0 2 15 3 0 9 9 11 13 1 10 9 2 11 11 2 2
7 9 9 0 12 9 0 2
16 10 10 10 9 15 3 13 9 9 15 1 0 13 1 9 2
12 15 3 13 9 11 11 11 1 11 11 11 2
23 1 15 15 13 3 9 9 0 2 10 9 3 13 1 1 9 9 9 9 7 9 0 2
85 13 9 9 1 11 15 13 1 11 11 11 11 11 15 13 1 13 9 7 9 1 9 9 11 11 11 11 2 13 10 10 9 9 16 11 2 11 11 15 13 16 9 9 9 9 9 13 1 9 9 7 9 9 10 9 9 2 9 9 2 7 11 11 11 15 13 9 9 15 0 7 13 1 13 11 11 11 11 2 9 2 1 9 10 2
19 11 7 11 11 2 11 11 2 13 9 0 1 9 9 2 9 7 11 2
12 11 13 13 9 1 1 1 7 1 9 9 2
34 13 9 9 16 11 11 13 9 2 9 9 11 12 2 11 11 1 12 2 7 11 2 9 11 11 12 2 11 11 11 1 12 2 2
25 1 9 10 2 3 9 15 13 13 9 1 11 15 13 2 7 1 9 3 13 3 1 13 9 2
17 9 10 13 9 9 12 8 2 9 7 9 12 9 2 12 2 2
22 11 13 9 15 3 13 9 9 0 2 3 13 9 2 9 2 9 7 9 9 0 2
10 9 13 9 0 1 9 7 9 9 2
36 10 2 10 9 11 1 12 9 10 13 1 9 9 2 15 13 9 9 0 2 7 9 9 2 15 13 9 9 13 11 12 2 2 12 2 2
19 11 15 13 1 9 2 9 11 13 9 9 11 7 9 9 1 9 11 2
29 16 3 2 11 13 1 9 1 13 10 9 9 2 1 9 1 9 13 9 9 0 15 13 1 9 2 9 0 2
61 9 9 1 9 11 11 13 1 9 9 11 11 11 13 9 9 12 5 7 9 12 5 15 13 1 9 11 11 12 5 12 1 9 9 12 7 12 5 12 1 9 11 12 2 1 13 9 9 9 2 13 9 9 0 1 9 0 12 9 12 2
26 15 3 13 9 11 11 7 9 10 13 9 9 11 11 11 7 9 9 9 11 11 2 11 2 11 2
25 16 3 13 2 11 13 10 9 15 13 9 9 1 9 1 11 11 2 11 10 13 9 9 9 2
26 15 13 9 10 7 9 1 11 11 1 9 12 1 9 12 16 15 13 13 1 10 9 0 1 9 2
22 11 11 13 10 9 1 9 0 11 11 15 3 13 1 11 7 11 2 11 5 11 2
14 16 9 2 9 13 2 11 13 9 15 13 1 9 2
17 3 1 9 10 15 3 3 13 9 1 9 9 1 1 9 0 2
64 11 11 11 13 13 9 15 13 1 11 1 11 1 12 9 12 2 11 11 11 13 9 2 9 15 1 0 13 1 9 2 1 9 1 9 7 9 11 11 11 2 1 10 13 9 9 9 7 9 11 11 11 2 11 11 2 12 1 11 11 12 11 12 2
15 11 9 10 13 1 12 9 15 13 11 11 1 11 11 2
11 3 3 1 11 7 11 1 15 3 13 2
9 11 9 13 9 7 9 1 0 2
10 11 13 3 14 11 11 15 13 0 2
12 11 11 13 10 9 15 13 1 11 11 11 2
13 11 13 9 15 13 1 11 11 2 11 9 9 2
20 10 0 9 13 10 13 9 15 13 1 11 2 16 15 13 9 0 3 13 2
24 9 9 11 3 13 3 1 9 9 0 2 7 9 9 11 13 3 1 9 9 0 2 0 2
18 11 2 9 11 2 11 1 11 2 13 10 9 1 9 11 1 11 2
23 16 11 1 11 2 11 13 1 11 11 2 10 9 0 15 3 13 1 9 9 1 11 2
21 1 9 9 2 9 9 13 2 11 13 12 9 15 13 11 1 11 11 11 11 2
7 3 11 3 13 1 11 2
5 2 9 11 11 2
9 3 16 9 10 3 13 12 9 2
13 3 2 2 3 16 11 13 9 15 13 1 11 2
24 1 9 10 2 15 13 1 9 9 11 11 2 7 9 10 13 9 0 1 9 12 2 12 2
17 3 0 2 3 13 12 9 1 12 9 9 1 0 7 3 0 2
114 11 11 13 10 9 9 1 9 11 1 11 15 13 2 5 11 11 11 11 5 11 11 11 11 5 11 11 11 5 11 11 11 5 11 11 11 5 11 11 11 11 5 11 11 11 11 5 11 11 11 11 5 11 11 11 11 5 11 11 11 11 5 11 11 2 11 11 11 5 11 11 11 11 11 5 11 11 11 11 5 11 11 11 11 5 11 11 11 11 11 5 11 11 11 11 5 11 11 2 2 11 11 11 11 5 11 11 11 11 11 5 11 11 11
25 9 2 11 11 2 13 9 9 9 9 11 11 7 1 9 11 12 3 13 13 9 11 11 11 2
21 9 0 10 13 9 0 7 13 9 9 1 11 2 11 11 1 11 11 11 11 2
21 1 9 15 3 0 2 9 10 3 13 1 10 9 9 9 9 7 9 9 9 2
7 3 13 10 9 1 11 2
15 1 9 9 2 9 10 13 1 9 9 13 1 9 9 2
26 11 11 13 10 9 1 11 11 11 15 13 9 9 12 9 2 7 9 12 2 12 9 2 12 2 2
16 11 7 11 13 9 0 15 3 13 1 9 9 1 10 9 2
33 11 2 2 13 10 9 1 11 11 2 11 2 13 1 9 9 11 11 2 9 9 2 12 2 9 12 2 2 12 2 12 2 2
17 9 9 11 13 9 9 15 13 1 11 11 16 1 9 11 11 2
10 16 16 14 3 2 11 14 13 9 2
62 15 13 10 9 0 1 9 9 9 9 1 9 12 5 12 13 1 9 11 2 9 9 0 14 13 1 9 9 2 7 3 13 9 9 9 15 3 1 0 9 13 9 0 3 0 3 13 9 0 12 1 9 0 7 13 1 9 9 15 14 0 2
9 3 9 13 2 9 9 11 9 2
15 11 11 13 9 1 11 11 2 16 9 9 13 11 11 2
36 11 13 3 3 9 1 9 12 2 12 15 13 1 9 9 9 15 3 3 9 1 1 9 11 2 15 13 9 11 1 11 11 3 12 3 2
28 11 11 1 11 11 13 3 2 2 7 14 13 9 2 16 15 10 15 3 0 1 11 2 3 13 1 9 2
22 11 13 10 10 9 15 13 1 11 11 11 2 11 11 2 11 11 11 11 2 11 2
7 9 1 11 11 11 11 2
16 9 9 1 9 0 3 0 7 13 9 15 0 1 9 0 2
16 1 9 12 2 9 10 13 9 1 12 9 7 12 9 9 2
11 9 9 9 2 2 3 9 15 15 13 2
21 11 10 13 1 10 9 0 7 0 1 11 11 2 1 11 11 1 9 11 11 2
13 11 3 13 9 1 11 11 11 2 7 11 11 2
11 9 11 13 1 9 9 2 11 11 2 2
23 11 11 2 2 13 10 9 9 9 13 11 15 13 1 9 11 12 3 13 1 9 9 2
5 11 13 9 11 2
17 15 14 0 13 3 9 1 9 9 1 11 11 10 13 1 9 2
21 15 13 13 9 2 9 10 13 9 15 13 9 9 7 13 9 1 9 2 9 2
21 11 11 11 2 2 13 9 9 9 9 11 7 9 10 13 1 9 9 11 11 2
7 11 13 1 9 13 0 2
30 0 9 12 2 11 3 13 9 1 9 9 1 9 2 13 9 2 9 10 13 1 9 11 15 3 13 9 9 0 2
28 11 10 3 3 3 13 1 9 3 7 3 1 9 9 9 2 9 9 2 9 9 2 0 2 7 9 13 2
26 1 9 2 12 9 10 13 9 2 9 2 7 9 2 9 0 13 9 0 2 9 2 7 9 2 2
13 11 13 12 5 9 9 11 11 2 9 11 11 2
32 11 10 13 1 11 11 1 1 9 2 1 11 1 1 9 2 1 11 11 11 1 1 9 7 1 11 11 11 1 1 9 2
9 1 9 12 2 11 13 11 11 2
19 1 10 2 9 9 9 0 1 11 1 0 13 7 9 9 7 9 9 2
27 11 11 13 9 15 1 9 16 11 7 11 11 11 2 1 10 1 13 1 9 9 2 9 2 7 9 2
17 9 10 13 12 2 12 10 13 9 10 2 12 1 9 11 11 2
14 11 13 1 9 11 11 11 11 1 12 9 2 12 2
17 9 9 10 13 1 9 2 11 11 11 2 2 11 11 11 2 2
36 1 9 12 2 15 3 13 11 2 2 2 11 11 7 9 2 11 2 15 0 1 0 7 1 12 9 10 2 11 13 10 9 1 11 11 2
30 11 11 3 13 9 1 9 9 11 2 11 11 2 15 3 13 1 11 1 2 9 11 2 2 7 9 9 11 11 2
22 1 13 11 3 13 9 1 10 9 2 13 10 9 11 7 11 15 13 9 9 0 2
14 1 9 11 12 2 9 11 13 7 11 13 1 11 2
18 3 3 1 10 9 3 13 9 9 1 1 13 9 10 14 13 13 2
18 1 10 11 11 11 11 3 13 1 9 1 13 13 1 13 9 10 2
40 9 10 1 13 1 11 11 1 11 11 2 9 1 10 11 7 9 11 11 11 2 11 11 3 13 1 11 11 11 11 2 10 11 15 13 1 11 11 11 2
28 1 9 12 2 11 13 9 11 2 7 13 9 9 9 15 13 0 0 12 1 9 2 7 13 9 1 11 2
18 11 11 13 9 9 9 1 11 11 11 2 11 2 11 11 2 11 2
20 1 9 10 15 13 1 11 11 11 1 11 11 11 13 1 11 11 2 11 2
7 11 11 13 9 11 11 2
21 13 9 7 9 2 9 2 9 11 11 13 3 9 0 15 0 1 9 7 9 2
36 1 10 2 11 11 11 3 13 9 9 11 1 9 11 1 11 11 2 1 13 13 9 15 13 1 2 9 15 3 13 9 1 11 11 2 2
19 11 9 1 13 7 9 9 15 9 1 9 15 3 13 1 9 9 0 2
12 9 7 9 13 9 9 15 13 1 9 11 2
15 1 11 11 7 11 13 9 0 2 16 9 11 11 11 2
17 11 3 13 2 2 3 14 15 13 13 15 3 0 7 0 9 2
30 9 0 2 1 9 9 7 9 0 9 9 0 13 0 2 9 9 0 3 13 1 9 9 7 3 13 1 9 0 2
15 1 12 9 12 2 9 10 9 9 0 1 9 2 12 2
9 9 9 10 13 9 1 9 11 2
9 9 10 13 1 9 9 11 11 2
11 11 11 11 13 10 9 11 1 11 11 2
32 16 9 11 11 2 11 14 0 16 15 3 13 1 11 11 2 15 1 0 9 7 9 2 9 2 9 10 13 1 9 11 2
6 15 13 2 3 9 2
40 11 11 11 13 9 9 9 0 15 13 11 2 11 11 11 2 11 2 1 11 11 1 9 12 2 12 1 9 11 2 11 2 2 11 2 11 2 7 3 2
18 1 10 9 15 13 1 11 11 2 12 2 12 5 13 1 9 9 2
15 16 9 12 9 9 10 3 0 2 15 3 13 9 0 2
31 1 9 15 13 9 1 9 2 9 2 2 9 13 2 16 1 9 9 9 1 9 2 9 9 3 0 13 1 9 13 2
27 11 3 3 13 9 9 2 11 2 15 13 9 0 11 11 2 16 1 12 3 13 9 1 9 9 11 2
34 11 2 9 10 9 1 9 15 13 1 12 2 11 11 11 11 2 11 11 11 11 2 11 15 11 11 2 7 11 15 11 11 2 2
14 9 10 3 13 1 9 0 2 11 2 16 14 9 2
50 10 9 9 9 9 0 13 1 9 9 9 13 9 9 2 1 1 9 11 2 11 3 13 1 9 0 12 11 11 11 13 1 11 2 12 9 2 7 11 2 12 9 2 1 9 11 7 11 11 2
18 16 10 2 9 3 13 13 9 2 9 9 2 1 2 9 9 2 2
10 3 11 13 7 13 11 1 12 9 2
21 11 11 13 10 10 9 15 13 1 9 11 2 11 11 11 2 11 11 2 11 2
15 11 9 1 9 10 13 11 11 13 13 9 9 9 11 2
9 9 13 1 9 0 15 13 9 2
15 1 11 12 2 11 13 10 9 9 11 1 9 1 13 2
30 0 9 1 9 11 11 11 2 11 11 1 13 9 1 11 11 11 13 9 1 12 2 12 9 13 9 11 11 11 2
30 11 11 15 3 3 13 12 9 9 11 11 2 3 13 11 11 1 11 11 11 2 7 2 9 15 13 1 9 2 2
33 11 11 2 2 13 9 9 9 0 11 11 0 15 13 1 11 2 7 3 13 1 9 0 7 9 0 1 9 11 11 11 11 2
11 9 10 13 9 1 9 10 9 9 0 2
14 11 13 9 1 11 11 2 11 2 11 11 2 11 2
20 9 11 13 9 9 1 9 11 11 11 2 11 11 2 11 11 11 2 11 2
11 11 11 13 12 2 11 11 7 11 11 2
19 11 1 3 13 9 1 9 9 2 1 9 9 2 7 13 1 9 9 2
12 10 1 9 10 3 13 1 9 13 1 9 2
18 11 13 16 9 15 11 13 3 9 9 15 0 7 0 2 9 2 2
72 13 10 9 9 1 3 13 7 13 9 9 10 15 9 10 3 13 1 11 11 12 2 12 1 13 11 11 2 12 9 12 1 9 7 9 11 11 11 13 9 15 13 1 9 9 9 9 11 13 9 1 12 5 2 13 9 9 15 13 9 9 0 2 9 9 10 1 11 1 11 11 2
32 1 9 13 11 7 13 11 2 9 9 10 9 7 9 2 2 15 3 13 13 11 2 13 10 9 2 7 13 9 9 11 2
11 11 1 9 12 2 13 9 1 12 9 2
18 11 11 13 10 10 9 1 11 11 2 11 11 2 11 11 2 11 2
8 11 13 9 0 1 9 11 2
58 1 9 9 15 0 1 9 9 9 2 13 1 12 9 16 9 9 15 13 9 9 13 1 12 2 12 9 1 9 12 2 12 5 7 9 9 9 9 13 9 9 1 12 2 12 9 2 9 9 15 3 3 13 1 9 9 9 2
12 11 11 13 3 1 11 11 7 3 11 11 2
23 9 0 1 11 3 13 9 15 16 9 0 13 1 9 11 11 2 9 0 9 3 13 2
8 16 9 13 11 12 3 13 2
19 15 3 3 13 1 11 11 11 11 11 12 1 11 11 2 11 11 11 2
20 9 9 13 1 9 12 2 12 9 0 2 11 5 12 2 1 12 11 12 2
32 11 2 11 2 2 13 11 11 2 11 11 2 11 11 1 13 0 7 11 11 7 11 11 1 9 0 1 9 9 9 10 2
9 11 3 13 1 9 9 7 9 2
44 9 9 13 1 11 11 11 2 13 9 9 1 9 9 2 9 2 9 9 0 9 1 9 0 2 7 9 0 9 2 9 2 9 9 7 9 2 1 9 9 7 9 0 2
20 1 9 9 9 2 11 13 10 9 2 11 11 11 2 13 12 11 12 2 2
20 9 0 2 11 11 2 13 9 1 9 2 9 15 13 9 7 13 9 9 2
20 9 9 10 13 11 11 2 11 11 2 11 11 2 11 11 2 7 11 11 2
14 11 13 9 1 9 11 2 11 2 11 11 2 11 2
20 11 13 11 2 1 13 1 11 2 2 13 11 2 3 15 3 13 3 11 2
11 9 10 3 13 10 9 9 0 9 9 2
61 1 12 1 12 2 11 13 9 2 9 7 9 1 11 2 11 7 11 1 9 9 7 1 13 0 1 0 1 11 11 7 11 11 2 11 9 13 11 11 2 11 0 1 10 9 0 13 9 9 1 9 9 2 7 9 9 1 9 2 9 2
29 1 9 12 2 11 11 13 9 15 0 15 13 1 9 11 2 11 11 2 16 11 11 13 9 9 1 12 9 2
7 9 15 13 13 9 11 2
25 11 13 11 1 13 9 1 11 2 11 2 7 11 13 1 13 13 9 2 14 13 16 13 9 2
14 15 3 13 1 9 0 1 9 12 1 9 12 9 2
11 11 13 1 9 12 1 13 13 11 11 2
21 15 13 1 9 12 9 1 11 11 9 12 2 1 3 13 9 9 1 9 12 2
14 11 13 9 1 11 11 2 11 2 11 11 2 11 2
69 9 9 11 11 11 2 9 3 13 1 9 2 11 11 11 2 11 13 1 12 9 15 13 2 16 9 9 7 9 11 1 9 0 2 9 9 13 12 2 12 9 5 9 7 9 13 12 2 12 11 2 16 13 9 1 12 5 2 12 5 7 9 9 13 12 2 12 9 2
45 11 11 13 9 9 11 11 1 9 2 11 3 13 13 12 9 3 2 11 2 9 2 2 11 11 2 11 2 2 11 11 2 11 2 2 11 11 2 11 2 2 7 11 11 2
17 11 13 9 15 13 1 11 11 2 11 11 2 11 11 2 11 2
22 11 11 11 2 13 11 11 2 13 9 1 13 9 15 0 2 7 3 13 9 9 2
22 11 11 13 10 10 9 15 13 1 11 11 11 2 11 11 11 2 11 11 2 11 2
14 1 9 2 11 13 9 11 11 1 9 15 13 11 2
22 2 7 2 3 15 13 1 0 1 10 9 2 7 14 1 15 2 7 14 3 0 2
7 3 9 13 9 9 9 2
19 9 10 3 13 1 9 1 0 3 10 9 3 13 16 3 0 1 9 2
22 15 3 13 7 13 12 9 9 11 11 11 11 13 12 2 11 2 11 2 7 11 2
15 1 9 9 13 2 9 9 13 9 10 9 1 13 9 2
86 9 9 13 10 9 9 15 13 9 1 13 1 9 15 3 3 1 9 1 9 9 2 15 13 9 9 0 12 5 2 2 9 9 10 13 11 11 2 9 1 9 11 15 13 9 11 2 11 11 2 1 9 2 7 11 11 2 9 11 15 13 13 9 1 9 9 2 11 11 2 7 10 9 9 2 9 9 2 15 3 13 1 9 9 2 2
48 3 13 13 1 12 12 9 2 3 9 11 11 13 3 3 3 3 0 1 11 11 2 16 3 1 1 10 1 9 9 3 15 3 13 11 11 15 9 13 12 2 12 9 0 11 11 11 2
19 11 15 3 13 1 10 9 11 11 7 9 2 9 2 9 2 7 9 2
11 1 12 2 11 11 13 9 11 12 11 2
11 9 10 13 9 13 1 3 0 9 12 2
11 1 9 10 15 13 13 10 9 9 0 2
30 15 3 13 9 9 9 7 9 9 0 1 11 2 11 2 9 2 7 13 10 13 9 1 13 13 9 1 9 0 2
21 1 9 2 9 0 2 9 13 1 11 11 15 13 1 9 11 13 12 9 11 2
18 11 13 9 12 9 1 11 11 2 11 11 11 2 11 11 2 11 2
9 0 9 11 1 11 7 11 3 2
15 11 11 2 12 9 13 9 9 11 2 11 9 11 12 2
34 11 9 11 13 1 1 12 9 2 3 11 11 2 13 1 11 11 7 11 11 2 7 11 11 2 13 1 11 11 7 11 11 2 2
20 11 11 10 13 1 9 1 13 9 0 16 13 1 0 9 7 1 9 10 2
50 16 1 9 9 2 9 9 11 5 11 15 0 2 1 11 11 11 11 1 11 2 11 11 11 2 11 11 11 7 11 11 1 11 3 13 9 9 9 3 3 3 13 9 9 7 9 9 9 11 2
18 11 11 10 1 9 11 13 1 9 11 11 11 11 7 11 11 11 2
47 11 11 11 3 13 9 11 1 11 1 11 11 2 16 9 10 14 9 12 9 11 11 13 1 11 7 11 2 16 10 10 9 9 9 9 10 13 0 1 9 3 13 9 11 7 11 2
11 0 1 9 10 13 1 12 1 12 9 2
15 14 2 9 2 0 15 1 15 2 14 3 0 1 9 2
30 1 9 10 2 11 13 1 9 11 12 1 11 11 2 3 13 11 11 1 9 11 2 11 11 11 11 11 2 12 2
15 9 9 11 11 13 1 9 9 9 11 10 15 13 11 2
97 1 9 11 2 9 11 11 9 12 13 9 1 9 9 11 15 13 11 11 7 1 9 0 2 1 9 2 9 11 3 13 9 2 9 2 7 1 9 13 9 11 12 2 12 9 11 13 13 9 1 9 9 9 9 0 2 15 3 1 9 9 16 9 2 9 11 11 2 3 13 7 11 2 11 11 2 3 13 9 9 11 1 0 3 13 13 1 10 9 9 13 1 11 1 12 9 2
9 11 10 9 1 9 9 9 11 2
17 9 10 3 13 3 1 11 7 9 2 9 13 9 9 11 11 2
33 16 2 13 3 15 13 16 3 13 12 9 9 2 15 9 13 0 7 3 13 2 16 15 10 3 13 3 0 7 3 0 13 2
10 3 2 11 13 1 9 7 13 9 2
17 15 3 13 1 9 0 11 15 13 1 9 11 11 2 11 11 2
15 11 13 9 1 11 11 2 11 11 2 11 11 2 11 2
23 1 9 12 2 1 9 1 9 11 7 9 2 15 13 11 13 9 0 0 2 11 12 2
16 10 2 10 9 9 13 1 3 12 9 9 2 13 7 9 2
21 11 11 3 13 10 9 2 13 1 11 11 2 11 11 2 11 11 2 11 11 2
11 11 1 9 12 2 13 9 1 12 9 2
30 9 11 12 2 11 13 13 9 9 0 1 9 12 2 11 2 2 7 1 9 11 2 11 13 9 9 12 2 11 2
14 1 9 9 3 13 9 1 13 9 0 7 9 9 2
14 11 1 9 13 9 2 15 2 3 2 14 3 0 2
16 11 13 10 10 1 3 9 9 15 9 13 1 9 9 11 2
82 11 3 13 1 10 9 9 11 2 15 3 13 1 14 0 2 8 2 11 7 7 9 2 16 2 11 11 3 13 1 9 12 2 12 2 3 13 1 0 9 11 1 11 11 2 7 13 1 9 2 9 1 12 2 12 1 9 1 11 11 2 15 3 13 1 2 9 2 0 12 1 11 11 2 11 10 3 0 1 11 11 2
18 11 13 9 15 13 1 11 11 11 2 11 11 11 2 11 2 11 2
28 1 10 9 1 11 11 11 2 1 9 2 9 0 11 13 1 9 2 9 1 9 0 7 9 15 1 11 2
25 11 13 9 15 0 2 3 15 3 13 9 0 1 13 13 9 2 7 15 3 13 9 1 9 2
15 15 3 13 9 0 1 2 11 11 2 1 12 11 12 2
13 2 11 9 1 9 15 3 0 3 3 13 3 2
14 11 2 2 11 13 10 2 10 9 11 15 13 0 2
13 10 9 13 9 0 1 9 1 9 12 11 12 2
15 9 16 9 13 2 15 13 12 9 1 11 7 13 0 2
12 9 10 3 13 3 1 11 12 7 11 12 2
21 15 13 9 9 11 11 2 9 9 1 11 13 12 9 2 12 2 12 9 2 2
34 11 11 2 11 2 7 9 9 13 9 7 9 9 2 9 9 2 7 0 1 9 9 7 9 1 11 11 7 1 3 12 9 0 2
18 11 13 10 9 15 13 1 11 11 2 11 11 11 2 11 2 11 2
7 9 15 13 0 2 0 2
17 11 13 1 9 9 9 9 2 9 2 9 2 7 9 0 9 2
7 7 3 3 9 9 10 2
22 1 13 11 2 11 2 9 10 9 9 2 7 13 10 9 7 9 2 9 1 9 2
21 11 13 1 9 9 2 7 9 13 9 9 11 11 2 11 11 1 13 9 0 2
32 9 9 9 11 3 0 1 11 7 11 11 2 1 9 9 1 1 11 11 7 11 11 2 7 1 9 9 2 16 9 11 2
21 11 11 2 2 2 11 2 11 11 2 13 10 9 11 15 13 1 9 9 9 2
10 1 10 9 3 13 1 13 9 0 2
18 15 13 9 11 11 11 11 11 12 2 1 9 11 9 12 11 12 2
10 3 11 3 13 9 9 11 7 11 2
34 15 13 9 9 12 1 9 1 12 9 1 9 12 2 12 1 11 11 2 10 9 9 13 9 12 9 9 1 11 11 7 11 11 2
9 11 11 13 9 11 1 11 11 2
26 9 10 13 13 1 9 11 2 11 11 2 2 7 9 2 0 2 11 2 10 9 0 11 9 9 2
18 11 13 10 9 15 13 1 9 11 2 11 11 2 11 11 2 11 2
17 9 15 13 1 11 11 10 13 1 0 1 11 11 7 11 11 2
38 11 9 0 13 1 10 9 5 9 2 7 10 1 3 3 13 9 2 11 9 9 13 9 7 9 1 11 2 11 13 10 10 9 0 15 3 0 2
14 9 10 13 9 3 0 1 1 9 2 9 9 0 2
24 16 15 3 11 13 9 2 11 2 1 9 2 7 2 7 15 3 16 2 10 9 13 9 2
27 9 10 13 9 0 15 13 16 0 3 13 7 13 1 9 2 9 0 1 1 9 7 1 9 2 9 2
49 1 9 11 2 11 1 9 13 9 9 2 9 2 7 9 2 2 2 1 9 7 9 9 9 11 13 10 9 2 3 7 2 1 9 9 11 1 1 9 9 13 9 9 13 10 9 2 2 2
11 2 9 2 1 11 15 1 11 7 11 2
20 3 9 2 9 2 13 1 11 11 2 9 2 7 2 9 11 13 13 9 2
12 12 9 2 2 15 13 9 9 9 1 11 2
6 3 3 15 13 9 2
16 11 11 13 3 1 9 11 11 11 1 9 9 11 11 11 2
8 3 0 9 2 3 0 13 2
21 1 9 9 2 15 13 0 2 7 13 1 9 16 9 3 3 2 3 13 1 2
28 9 0 13 2 11 11 2 15 13 1 10 12 12 11 11 15 13 1 9 12 2 12 1 9 1 12 12 2
23 16 1 13 9 7 3 13 1 11 11 11 11 12 2 11 2 11 2 2 9 11 0 2
16 3 2 10 9 0 3 13 9 1 9 11 2 11 1 12 2
29 9 9 9 10 13 13 2 0 1 11 11 11 11 2 16 9 2 9 15 3 13 0 13 9 9 15 0 3 2
12 9 13 9 11 11 1 13 9 9 15 13 2
17 1 9 12 11 12 2 11 11 12 9 11 11 1 9 9 10 2
18 11 11 11 13 1 11 2 7 11 13 9 9 1 10 9 1 11 2
25 11 13 10 9 1 11 2 11 11 2 11 15 13 12 5 1 0 11 7 12 5 1 0 11 2
17 7 1 9 15 13 13 15 13 1 11 3 1 9 1 9 0 2
23 9 11 9 15 3 0 13 13 11 11 11 7 11 11 2 9 10 3 13 12 9 10 2
49 16 10 11 11 3 3 13 1 11 11 11 11 7 13 12 9 9 1 11 11 7 11 11 2 9 13 1 9 0 1 11 11 1 9 12 7 13 9 12 2 12 15 13 13 1 11 11 11 2
10 16 3 10 9 9 0 3 13 9 2
22 13 1 11 11 5 11 9 11 11 2 15 13 11 11 11 11 1 9 0 9 12 2
14 11 11 2 11 2 2 3 13 0 1 9 9 11 2
17 11 3 14 13 9 9 16 9 3 13 1 9 1 9 10 3 2
48 1 9 11 1 11 15 13 3 1 9 9 2 9 11 13 9 0 1 9 11 2 1 9 11 2 9 11 13 13 9 2 9 2 9 2 9 9 2 2 9 0 2 7 9 9 1 9 2
76 13 9 9 9 2 15 13 11 11 11 11 11 11 11 11 2 16 13 11 11 2 13 11 11 11 11 2 7 1 11 11 13 11 11 11 2 9 11 10 13 1 9 10 2 9 2 15 13 2 11 11 2 2 16 15 3 9 9 9 12 1 9 11 2 1 9 12 15 13 11 11 11 1 9 9 2
16 9 10 3 13 1 9 11 11 11 11 2 12 2 12 2 2
24 11 11 13 3 1 11 11 7 11 11 1 11 12 1 13 7 13 9 1 9 9 9 0 2
24 9 3 3 14 13 1 9 7 10 9 9 3 13 1 9 10 2 7 10 9 13 9 9 2
37 9 9 11 11 13 1 9 0 7 9 9 2 1 9 9 13 1 12 5 11 2 12 5 11 7 9 9 13 1 12 9 2 12 9 10 9 2
13 2 3 2 9 2 13 13 9 2 16 14 13 2
30 1 10 9 7 9 2 11 11 13 3 2 3 10 11 7 10 11 1 9 1 13 9 9 9 7 9 1 1 9 2
12 9 10 3 13 10 9 1 13 1 9 11 2
27 9 11 15 3 13 1 9 11 11 7 11 11 13 0 9 2 12 0 2 9 9 1 9 9 11 11 2
8 11 9 13 9 7 9 0 2
18 11 11 11 2 13 9 2 13 10 9 9 15 13 1 9 1 9 2
15 9 9 9 15 13 10 9 3 9 10 13 3 12 12 2
38 1 1 9 10 13 9 9 11 7 9 15 2 9 9 15 13 1 15 13 2 7 13 9 11 0 2 0 1 9 11 0 1 9 7 9 9 11 2
14 11 13 9 1 11 11 2 11 2 11 11 2 11 2
10 15 3 9 9 13 9 1 9 10 2
15 11 13 9 0 12 1 11 7 9 7 9 0 1 11 2
17 9 12 11 0 3 13 1 9 12 11 12 3 1 9 11 11 2
48 11 11 15 13 13 10 9 1 9 0 11 11 0 2 7 3 3 14 3 13 11 11 2 3 15 13 9 0 1 13 11 11 7 13 3 13 2 10 13 11 11 11 15 3 13 1 9 2
29 16 9 10 3 13 9 2 16 9 15 0 1 9 9 3 13 9 7 9 15 13 1 9 2 9 15 3 0 2
8 16 9 10 13 1 9 9 2
19 11 9 13 10 9 9 15 13 3 13 7 3 13 16 14 13 9 9 2
20 11 11 15 3 13 13 13 9 9 2 16 10 3 1 9 9 7 9 3 2
23 11 13 10 9 1 11 11 2 11 11 11 2 11 2 7 13 9 9 7 9 11 11 2
36 1 9 12 2 11 13 1 11 11 2 10 9 11 11 2 7 13 12 9 9 2 9 11 11 11 11 7 11 11 11 15 0 13 11 11 2
23 9 11 13 1 9 2 9 10 2 1 9 11 12 2 9 9 11 13 12 2 12 9 2
7 9 15 13 9 10 1 2
6 2 9 9 3 0 2
3 3 13 2
45 1 9 11 2 11 7 9 9 0 1 11 11 3 2 0 1 11 1 9 9 2 10 9 0 13 9 7 9 1 13 1 9 2 9 2 9 2 7 9 15 13 9 9 2 2
15 9 2 9 1 11 10 13 1 9 9 7 9 0 11 2
5 9 9 2 11 2
26 10 0 11 2 11 12 2 11 2 2 11 2 11 12 2 11 2 2 7 11 3 13 1 9 10 2
36 11 9 13 1 12 9 1 9 11 11 1 12 11 12 2 16 9 9 1 9 9 2 15 1 9 3 13 9 2 13 1 9 12 2 12 2
13 11 11 13 1 9 11 11 11 11 11 9 12 2
14 15 0 1 13 13 10 9 9 15 13 1 9 10 2
13 10 9 13 13 10 9 15 0 1 9 1 9 2
8 11 3 13 16 11 3 13 2
9 11 1 13 9 9 1 11 11 2
20 11 3 13 1 9 9 1 13 9 9 2 9 2 7 9 1 9 7 9 2
19 10 13 9 0 0 15 13 9 11 2 11 11 11 1 10 0 9 9 2
19 9 15 0 13 9 13 9 0 1 10 9 2 13 1 9 9 1 9 2
12 11 11 11 12 13 1 11 2 11 1 12 2
10 3 15 10 3 13 7 9 13 15 2
13 9 9 0 3 13 1 9 0 7 0 2 0 2
6 9 10 13 9 11 2
45 9 10 13 9 1 12 9 1 9 2 9 0 1 11 2 11 2 11 11 7 11 1 11 11 11 1 11 9 11 12 7 13 10 10 9 9 0 1 9 2 13 9 9 2 2
24 9 9 11 1 13 9 11 2 9 11 11 11 2 7 11 11 3 13 10 9 9 1 9 2
20 1 12 9 2 13 12 9 9 15 13 1 11 7 13 11 1 12 11 12 2
18 11 11 15 13 1 9 12 2 12 13 9 1 9 9 12 1 9 2
42 9 10 13 11 11 2 11 2 16 7 1 9 11 11 1 9 12 2 13 9 2 9 9 7 9 0 15 13 9 9 15 3 0 7 14 13 9 1 9 9 0 2
21 11 11 1 9 11 2 11 2 3 13 1 9 11 2 11 1 9 9 11 11 2
13 9 9 13 9 9 15 13 9 9 1 9 9 2
19 1 9 2 9 11 13 9 7 11 13 16 9 9 11 13 1 9 0 2
35 1 11 2 11 2 11 11 2 11 2 11 11 2 13 9 9 9 2 12 2 1 11 11 2 11 11 2 7 11 11 2 11 11 2 2
20 1 9 0 2 11 13 11 11 15 12 1 9 2 11 2 1 9 11 11 2
26 9 10 3 3 13 1 10 9 13 2 10 9 13 16 11 11 3 13 0 9 10 2 14 3 13 2
19 11 11 2 2 9 13 11 11 11 11 2 13 10 9 7 9 13 11 2
29 15 3 13 1 9 0 1 11 2 11 2 11 2 11 2 11 11 2 11 2 11 11 2 11 11 2 7 11 2
18 1 10 9 2 9 11 1 11 3 13 9 2 16 13 3 11 0 2
19 9 2 9 9 0 0 3 13 10 9 2 1 9 14 13 9 9 9 2
16 11 11 3 0 13 13 9 11 7 11 11 11 2 11 2 2
39 3 13 9 11 2 11 13 13 1 9 2 11 11 2 11 11 2 2 15 13 1 9 2 9 9 9 9 9 1 11 2 3 13 16 11 3 13 9 2
23 16 1 9 10 2 15 3 13 2 13 3 13 9 0 2 1 13 9 1 9 15 13 2
37 13 9 3 12 2 12 9 2 11 3 13 9 9 9 15 13 11 2 1 3 13 9 3 1 12 9 15 13 1 9 9 15 13 1 12 9 2
15 9 14 0 1 9 13 9 1 11 11 1 9 9 11 2
16 3 9 1 9 13 3 2 7 13 1 9 0 1 1 1 2
25 11 13 9 1 15 13 7 15 13 9 9 9 9 7 9 11 11 15 0 1 11 1 9 10 2
15 1 9 9 11 2 11 13 9 9 1 9 11 11 11 2
13 1 9 10 15 13 1 9 1 9 11 11 11 2
17 11 0 10 13 9 11 11 11 1 9 9 9 9 1 1 11 2
25 3 11 13 1 13 1 11 1 15 3 13 9 1 9 10 7 13 9 1 11 1 9 12 9 2
14 11 13 10 9 9 2 9 2 11 2 12 9 2 2
11 11 10 13 9 9 10 0 13 9 11 2
20 11 3 13 9 9 2 1 11 2 7 3 9 9 9 2 1 9 9 2 2
10 11 9 13 10 10 9 15 13 9 2
24 1 13 9 9 11 2 11 11 13 1 9 11 11 11 2 1 0 1 11 2 11 7 11 2
16 11 13 9 11 0 1 11 11 2 9 13 12 2 12 9 2
14 1 13 9 11 2 10 9 13 1 11 11 2 11 2
19 9 9 12 2 12 5 2 13 0 7 0 0 7 13 9 9 1 9 2
17 1 9 9 2 15 13 13 9 9 7 13 13 9 9 9 11 2
15 1 9 15 0 2 13 2 13 9 13 1 9 15 0 2
11 1 13 9 2 9 9 9 14 3 13 2
23 11 2 3 13 9 9 0 9 9 2 15 13 1 9 7 13 1 9 2 9 7 9 2
15 11 11 13 9 9 10 9 15 13 1 11 11 1 12 2
24 11 15 13 2 16 16 10 3 11 3 13 9 9 1 11 2 9 9 7 3 13 9 9 2
23 9 9 9 9 9 0 13 11 2 11 2 7 11 9 9 13 2 13 2 1 9 11 2
23 1 13 9 9 2 10 9 1 11 3 13 1 9 9 2 1 1 11 2 11 7 11 2
17 11 13 9 15 13 1 11 11 2 11 11 2 11 11 2 11 2
74 9 0 9 13 13 9 9 16 9 10 9 3 3 0 0 1 9 9 2 1 9 10 10 9 13 3 13 7 13 9 10 2 10 1 10 9 2 3 1 9 10 10 9 3 13 10 9 1 9 7 3 13 9 1 9 15 13 9 7 13 9 1 9 7 3 1 9 15 9 0 13 10 9 2
16 11 13 9 2 9 2 15 13 1 11 11 2 11 2 11 2
28 9 10 13 1 13 9 2 9 2 2 13 9 0 7 13 9 9 0 15 13 9 7 9 1 9 7 9 2
20 10 9 15 13 10 13 1 9 2 9 0 1 9 7 9 9 1 9 11 2
14 7 3 3 9 13 9 1 15 15 3 13 13 9 2
23 16 1 11 2 16 1 9 9 15 13 16 13 11 15 13 9 2 11 7 9 7 9 2
12 3 11 3 13 10 9 9 1 9 1 9 2
17 16 15 13 2 15 13 9 11 7 13 1 9 11 11 11 11 2
5 9 9 13 12 2
13 10 9 15 13 13 1 9 11 3 13 9 10 2
13 11 11 13 1 3 1 12 9 1 12 2 12 2
21 11 11 0 9 13 0 9 3 1 12 9 7 9 9 3 1 12 2 12 9 2
18 11 13 10 10 9 1 11 11 2 11 11 2 11 11 11 2 11 2
11 11 9 9 12 3 13 9 1 13 9 2
25 11 11 11 11 2 2 7 13 3 1 11 11 11 11 2 13 9 9 11 11 15 13 1 11 2
9 11 10 13 9 0 11 2 11 2
27 9 10 13 1 11 11 2 11 15 13 9 7 9 9 15 13 7 12 9 1 9 15 13 9 1 15 2
41 11 11 11 13 1 9 9 11 15 13 1 9 9 7 9 9 2 16 1 10 9 13 1 1 9 9 2 9 7 9 13 9 9 9 1 0 9 11 1 11 2
13 9 9 7 11 11 3 13 7 13 9 15 13 2
13 11 11 13 9 15 13 1 9 9 11 5 11 2
38 9 10 13 9 15 0 1 10 10 9 0 9 11 2 2 11 11 11 2 2 15 13 1 9 0 11 11 11 2 9 9 11 11 2 7 11 11 2
69 11 11 11 11 12 11 13 10 11 11 11 15 13 1 9 9 11 0 15 13 1 11 11 11 11 11 2 12 2 11 11 15 9 10 13 1 11 11 11 15 13 1 11 2 11 2 11 11 2 11 2 11 2 11 12 11 13 9 15 13 3 13 1 0 7 0 2 0 2
12 11 13 10 9 1 11 11 2 11 2 11 2
25 11 2 11 11 2 11 11 2 11 2 7 11 2 11 3 0 13 1 9 1 9 9 1 13 2
13 3 15 3 13 9 2 9 2 9 2 7 9 2
14 9 0 9 11 11 3 13 0 7 9 9 15 0 2
18 1 9 12 2 15 13 1 11 7 13 11 11 11 7 11 11 11 2
28 1 11 11 2 15 13 1 9 12 7 9 12 13 0 9 0 16 9 9 7 9 11 13 9 15 3 0 2
33 9 15 13 13 9 15 13 1 10 9 2 9 2 15 13 1 1 9 2 9 2 7 9 2 9 2 15 13 1 9 9 9 2
12 1 10 9 10 3 11 3 13 1 9 0 2
17 11 13 9 15 13 1 11 11 2 11 11 2 11 11 2 11 2
39 9 9 10 13 13 1 9 12 15 13 1 9 9 0 1 11 1 11 11 2 16 13 13 9 13 1 11 11 11 2 11 7 11 11 11 11 2 11 2
19 11 10 13 1 12 9 2 11 11 11 11 7 11 9 2 7 11 11 2
19 11 11 3 13 9 1 9 2 1 9 7 9 9 2 7 3 1 9 2
27 1 9 9 12 2 9 2 9 9 13 9 9 9 7 16 3 13 10 9 9 2 9 9 14 3 13 2
16 11 11 11 13 0 3 13 9 1 13 11 11 1 9 9 2
17 1 9 10 2 11 11 11 13 9 13 1 9 11 1 12 9 2
12 11 11 11 13 9 9 15 13 11 1 11 2
10 15 13 9 13 9 7 13 9 9 2
20 11 2 9 13 0 7 0 7 13 10 9 0 2 11 2 1 9 1 9 2
39 1 9 12 11 12 16 11 11 13 11 11 1 9 9 11 2 15 13 9 12 15 13 1 9 9 1 13 9 11 16 9 13 7 13 14 0 13 9 2
9 3 2 15 15 13 11 11 10 2
10 11 2 11 13 9 9 9 2 9 2
36 13 1 11 2 11 1 11 11 2 9 1 9 9 10 9 9 13 11 7 10 9 9 9 13 11 2 11 13 9 9 7 9 9 1 0 2
9 9 0 0 13 10 9 0 0 2
14 13 9 10 2 10 9 13 1 9 1 11 11 13 2
4 0 9 0 2
47 9 11 1 0 13 1 10 9 2 3 1 9 9 2 9 11 11 13 9 2 9 15 13 0 2 16 13 15 1 13 12 12 2 3 13 1 10 9 9 10 13 11 16 11 11 11 2
25 7 3 9 11 11 1 9 9 9 10 3 13 1 9 7 9 11 11 10 1 0 7 14 0 2
18 11 13 10 9 1 11 15 13 1 12 7 12 2 13 1 11 11 2
61 16 9 2 9 0 15 13 1 10 9 9 9 3 9 11 2 1 9 2 2 11 11 2 1 9 9 2 2 13 2 12 9 2 2 9 2 1 9 2 2 7 1 9 13 9 9 7 9 1 9 2 9 7 1 0 13 9 9 7 9 2
24 11 1 10 9 11 9 11 2 11 2 11 2 11 2 9 11 11 11 2 13 9 9 11 2
23 1 9 10 9 9 1 9 11 13 1 10 9 0 2 7 13 0 1 13 9 0 0 2
6 9 0 2 3 14 2
12 11 13 1 9 10 7 15 13 10 9 9 2
25 9 10 1 9 13 2 1 0 2 11 11 15 13 13 9 7 11 11 11 15 13 13 11 11 2
14 11 11 11 13 9 1 12 9 1 13 13 12 9 2
7 15 13 1 9 11 11 2
19 11 13 1 13 9 1 9 9 11 2 7 11 13 9 7 9 1 9 2
13 9 9 15 15 3 13 1 9 0 15 14 13 2
12 11 11 13 10 9 9 0 1 9 11 11 2
15 11 10 13 1 11 2 15 13 1 9 0 1 9 10 2
36 3 3 11 13 1 9 11 2 11 2 11 2 7 11 13 9 11 2 11 2 11 1 9 11 2 11 2 11 13 1 11 2 11 12 2 2
34 11 10 13 10 9 11 11 7 3 1 9 9 11 11 2 16 9 0 13 9 2 9 10 3 13 10 9 9 7 9 9 9 11 2
11 9 13 16 11 11 0 11 13 11 11 2
21 9 0 3 9 9 0 3 13 9 13 9 9 2 11 2 7 13 0 7 0 2
6 9 9 0 11 11 2
24 9 9 0 1 9 3 13 9 1 11 11 11 2 3 13 1 11 11 2 1 11 11 11 2
23 9 9 10 13 1 9 12 7 13 9 9 9 1 0 9 12 2 12 7 12 2 12 2
21 9 10 13 10 9 9 0 16 13 9 1 13 9 9 1 9 2 9 15 13 2
40 11 11 11 2 2 13 9 12 9 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 11 7 11 11 2 15 13 11 11 1 11 1 9 12 2
30 13 1 11 11 2 9 13 1 12 9 2 13 13 12 1 9 2 2 7 13 3 3 1 13 13 11 11 9 11 2
16 9 0 12 11 2 11 11 13 1 11 13 11 1 9 12 2
18 16 9 11 2 11 1 12 2 9 0 13 1 0 2 11 1 9 2
12 9 9 9 11 10 13 10 9 0 7 0 2
50 11 3 13 1 10 9 1 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 11 2 7 11 10 9 11 0 13 16 11 11 11 3 13 7 3 13 1 9 9 11 1 9 9 2
13 11 3 13 1 10 7 3 10 9 0 15 13 2
13 9 0 13 11 11 15 13 1 9 9 11 11 2
15 11 13 10 9 1 11 11 2 11 11 2 11 11 11 2
18 11 13 2 2 11 2 3 11 3 13 2 11 11 2 1 9 3 2
22 11 2 11 2 9 9 5 9 11 11 2 11 2 2 7 9 13 1 9 9 10 2
14 3 9 11 7 11 13 10 9 15 13 9 9 15 2
20 11 11 11 7 11 11 11 2 11 11 2 13 15 0 1 12 9 11 11 2
10 9 1 9 1 9 15 14 3 13 2
28 9 2 7 3 13 1 9 2 13 10 9 15 3 13 1 9 2 13 15 13 1 10 9 2 3 1 9 2
17 11 11 13 10 11 11 11 2 11 11 2 11 11 2 11 11 2
24 11 11 11 2 2 2 13 9 9 9 15 13 1 11 1 11 2 11 10 13 1 9 12 2
11 11 1 1 13 0 2 9 13 9 9 2
11 9 11 11 11 3 0 1 9 9 9 2
20 13 10 9 15 13 1 9 16 9 12 15 0 14 13 1 9 10 2 12 2
6 2 15 15 13 13 2
5 3 11 13 9 2
25 9 10 13 10 9 11 0 2 7 3 3 13 11 1 11 2 16 2 9 11 3 13 9 11 2
47 11 13 9 9 7 3 9 7 9 9 15 3 3 0 0 0 2 14 0 9 9 0 15 13 3 9 0 11 9 2 2 9 0 15 13 11 11 9 15 13 2 13 9 11 2 11 2
33 16 1 9 9 3 3 13 12 9 13 1 10 9 2 9 9 9 2 3 1 9 9 9 13 9 0 15 3 13 1 9 0 2
24 9 9 11 11 13 1 9 11 7 3 13 1 11 11 2 11 11 7 13 9 1 11 11 2
28 9 9 11 11 13 9 2 0 2 9 9 2 1 1 9 9 1 11 1 0 13 7 13 1 9 9 9 2
11 3 9 10 13 9 1 9 11 11 11 2
46 1 9 7 9 15 2 11 13 1 12 9 2 9 7 9 2 15 13 1 9 2 9 7 9 2 9 7 10 9 9 7 9 13 9 2 9 7 9 2 9 9 15 13 9 9 2
4 9 7 9 2
52 9 11 13 10 12 9 0 13 9 0 7 0 1 11 2 13 9 15 0 2 13 9 9 15 0 1 9 9 1 13 7 13 9 15 1 3 13 1 9 9 9 15 3 13 2 13 2 7 13 9 9 2
17 11 11 13 9 15 13 1 11 11 2 11 11 2 11 2 11 2
14 14 15 10 13 1 9 0 2 16 15 3 13 15 2
12 11 11 13 1 12 9 2 1 11 7 11 2
55 9 9 9 15 13 1 11 11 13 9 1 9 9 7 9 1 9 1 9 2 1 9 9 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 7 11 2 11 2 1 9 9 2 9 9 1 11 11 3 0 2
20 11 13 9 9 9 2 7 13 1 13 7 9 9 11 2 1 10 9 9 2
27 1 11 2 9 9 2 9 11 1 11 2 11 2 11 11 2 11 11 11 2 13 1 9 11 1 11 2
9 9 0 1 11 13 11 2 11 2
8 11 13 3 0 11 3 13 2
21 15 13 9 3 1 9 9 9 9 2 9 3 2 16 15 14 3 13 3 3 2
13 9 9 0 1 11 3 13 1 9 1 9 0 2
45 1 0 2 9 10 13 13 9 2 9 9 2 11 11 11 2 11 11 11 7 11 11 11 2 11 11 11 2 11 11 2 11 11 2 11 2 11 2 7 11 11 7 11 11 2
17 10 9 10 13 12 9 3 2 11 11 2 11 11 7 11 11 2
24 11 13 9 1 11 2 16 11 11 2 9 12 2 12 2 13 11 7 11 1 9 13 9 2
31 13 9 10 9 9 15 13 10 9 9 7 13 9 2 9 7 9 9 16 3 1 9 2 9 7 9 2 9 9 0 2
8 16 13 11 9 9 3 13 2
7 12 9 10 3 3 13 2
30 2 10 9 2 9 10 2 1 9 1 9 12 2 1 9 11 1 9 2 2 13 1 3 9 1 11 0 7 11 2
26 11 11 7 9 9 2 11 11 2 13 9 9 9 0 2 9 1 11 11 1 0 9 12 2 12 2
28 11 11 2 15 13 2 13 1 9 9 11 2 13 9 9 1 9 10 15 13 9 1 11 9 9 15 0 2
17 9 9 1 9 12 15 13 1 11 11 1 9 9 9 11 11 2
6 7 9 1 11 0 2
15 9 13 1 12 2 12 9 15 13 2 7 9 13 0 2
15 9 0 15 13 9 0 2 13 2 13 1 9 9 9 2
16 11 9 1 11 13 2 9 10 13 9 11 7 1 9 9 2
25 1 9 12 2 12 2 7 12 2 9 9 0 1 9 11 2 3 9 9 13 9 15 3 13 2
13 0 3 16 9 2 9 9 2 1 13 9 9 2
45 11 11 11 13 1 11 11 1 9 2 9 2 7 9 2 16 9 9 15 13 1 9 9 3 13 1 9 9 10 1 9 15 0 2 3 12 2 12 1 1 12 2 12 2 2
19 3 2 3 9 10 3 13 1 13 9 9 1 11 2 7 14 11 0 2
23 9 10 13 9 1 9 7 9 1 9 1 13 1 9 15 3 0 16 13 2 7 3 2
34 16 9 9 15 3 3 13 1 9 9 13 9 9 2 9 9 7 9 9 15 13 1 9 9 1 1 9 7 9 9 15 0 9 2
41 11 11 2 15 13 9 0 13 9 1 12 2 12 2 1 1 9 11 11 2 13 13 9 0 1 11 11 1 11 2 15 13 9 0 1 13 9 1 9 12 2
31 3 9 9 2 11 2 9 2 11 2 15 9 0 1 9 11 11 3 13 9 9 13 1 11 11 11 11 1 9 12 2
17 3 2 9 3 13 9 1 9 15 13 7 9 9 9 1 9 2
31 1 13 9 12 10 2 10 9 1 9 9 1 11 13 11 11 9 1 13 9 1 13 1 9 11 11 11 1 11 11 2
21 1 9 15 13 2 11 3 0 1 11 11 15 13 9 9 1 9 1 9 12 2
23 7 9 10 13 10 9 9 15 9 13 1 9 0 1 9 11 15 13 1 11 13 11 2
27 16 13 3 0 1 9 15 13 1 9 2 9 9 9 13 10 9 0 1 9 1 9 0 7 9 0 2
10 1 9 9 11 11 7 13 11 11 2
22 9 3 0 16 11 11 2 11 2 10 9 2 1 11 11 13 9 1 9 1 12 2
19 13 11 11 1 12 1 9 9 11 7 9 9 9 9 9 9 9 11 2
4 9 13 11 2
47 1 9 9 3 13 9 9 15 13 1 9 12 1 11 11 1 12 9 2 9 9 1 12 9 2 11 11 1 12 9 2 9 9 1 12 9 2 7 9 5 9 9 9 1 12 9 2
10 11 11 13 9 13 12 2 0 9 2
22 1 10 10 9 9 13 9 0 2 9 15 13 1 9 2 16 15 13 10 9 10 2
9 3 15 13 15 13 9 1 9 2
36 11 11 1 11 3 0 1 9 9 11 11 11 15 13 1 9 12 9 2 11 11 11 13 1 11 11 11 15 3 3 0 13 9 13 11 2
39 9 2 9 0 1 9 11 11 12 7 11 11 12 2 15 13 9 9 11 11 2 11 11 2 11 11 2 2 13 9 9 2 9 9 12 2 1 11 2
11 1 9 12 9 10 13 9 1 12 9 2
30 9 0 15 14 3 13 0 1 9 16 0 13 1 9 7 9 1 9 9 11 1 11 15 13 1 9 1 9 12 2
20 11 11 13 10 10 9 1 11 11 11 2 11 11 11 2 11 11 2 11 2
14 9 13 9 1 9 11 2 11 11 2 11 2 11 2
19 9 1 9 10 13 9 10 9 9 2 9 7 9 2 1 9 15 13 2
15 11 15 14 3 13 9 3 3 0 2 13 9 9 0 2
22 11 11 11 2 11 2 15 13 1 9 12 11 12 2 13 9 12 9 9 11 12 2
11 11 1 9 12 2 13 9 1 12 9 2
29 9 13 9 13 9 9 0 1 11 2 11 2 7 11 2 9 3 13 9 9 9 0 7 13 9 0 1 9 2
4 9 9 11 2
10 3 15 13 13 2 9 9 9 2 2
28 11 11 11 13 9 9 11 15 13 1 10 9 0 2 7 1 9 2 9 2 7 9 9 0 2 9 2 2
31 9 13 1 9 9 11 9 12 2 16 9 11 11 11 3 13 7 11 11 7 11 11 13 9 0 9 9 1 9 11 2
16 16 11 11 13 1 12 11 12 2 15 13 1 10 10 9 2
25 7 3 16 13 9 9 1 9 11 11 2 11 13 1 13 9 7 13 9 0 15 13 11 11 2
8 1 11 10 13 9 11 11 2
8 11 13 1 11 11 7 11 2
10 9 10 13 3 2 13 2 9 0 2
17 11 11 3 13 1 9 9 15 13 2 13 2 2 2 13 2 2
11 11 11 11 11 11 11 13 9 9 12 2
34 11 11 13 9 0 15 13 1 10 9 11 11 1 11 10 1 11 7 11 3 10 9 13 7 13 9 3 13 9 2 9 15 0 2
30 1 9 9 15 13 9 12 2 11 13 9 1 13 10 9 2 11 13 9 15 0 1 10 9 0 7 10 9 0 2
23 1 9 12 2 12 10 2 15 13 9 7 9 13 9 1 11 11 7 3 13 1 11 2
10 9 3 13 1 10 9 9 7 9 2
15 15 3 13 1 11 11 11 1 9 11 11 2 11 9 2
2 11 11
32 3 0 3 2 9 11 3 13 1 9 1 9 2 1 9 1 9 1 9 11 1 11 7 9 11 11 11 1 11 2 11 2
12 11 11 1 11 11 13 10 9 1 11 11 2
13 11 13 9 9 9 9 9 0 1 9 9 11 2
15 11 11 11 11 11 13 9 1 12 12 1 9 12 12 2
9 15 13 16 15 13 1 3 13 2
10 11 13 9 9 1 9 11 11 11 2
22 11 11 10 13 1 10 9 2 11 2 11 2 11 2 3 11 5 11 2 7 11 2
39 11 3 13 2 2 12 9 10 13 1 13 12 12 9 2 9 12 2 11 11 13 1 9 0 2 11 11 1 10 9 1 11 2 9 11 2 11 2 2
21 9 3 13 1 12 9 2 9 9 7 13 9 7 9 1 9 2 9 9 0 2
12 11 11 12 13 9 12 1 11 11 1 12 2
15 11 11 13 9 9 15 13 1 9 9 1 12 9 9 2
36 1 9 9 9 2 1 9 9 15 3 14 0 2 15 13 13 10 9 1 9 9 10 9 2 16 1 9 2 15 13 13 1 9 9 10 2
13 11 11 13 10 9 1 11 11 2 11 2 11 2
8 3 9 10 14 13 1 11 2
23 9 10 13 9 9 0 1 9 1 9 9 0 2 7 12 2 0 9 1 9 2 9 2
20 9 9 7 9 9 1 9 10 13 9 9 15 0 1 9 7 9 15 13 2
51 16 9 10 13 1 9 0 1 13 9 11 2 11 11 3 13 16 1 10 9 13 9 5 11 5 15 13 1 9 9 9 2 9 2 5 11 5 2 5 11 5 2 5 11 5 2 2 7 3 3 2
34 1 9 9 2 9 15 13 1 2 9 9 9 2 10 3 13 9 9 15 13 7 13 9 1 9 15 13 1 11 1 11 7 11 2
7 9 10 13 9 9 12 2
36 1 9 9 11 11 11 11 11 11 0 13 9 0 11 11 11 2 1 9 2 1 9 10 2 9 3 13 3 1 12 12 9 2 12 2 2
5 3 9 9 11 2
17 13 9 10 2 11 12 13 1 13 9 7 15 13 13 9 9 2
20 11 11 11 0 13 10 9 1 9 0 7 3 13 1 9 9 10 9 9 2
55 13 12 9 11 11 3 12 1 13 9 0 1 0 7 0 15 13 2 13 7 9 0 9 0 9 2 7 13 7 13 9 2 9 9 9 7 9 0 9 2 7 12 1 13 7 13 9 9 9 9 7 9 9 9 2
59 3 11 11 13 9 1 11 11 2 16 1 9 11 11 9 11 11 2 11 11 14 3 13 9 1 11 2 9 11 1 11 2 13 3 1 11 1 9 12 1 13 11 1 9 11 2 11 2 7 11 2 16 13 16 13 9 15 0 2
25 1 9 9 2 9 15 13 9 13 9 0 2 9 9 15 13 1 9 9 7 3 9 9 0 2
24 1 9 9 1 11 2 11 13 7 13 13 13 1 11 2 7 3 9 1 9 7 9 13 2
8 15 13 9 1 13 9 15 2
14 11 11 13 10 9 1 11 11 11 2 11 2 11 2
20 15 13 9 9 1 9 12 1 11 11 11 7 13 9 9 1 11 11 11 2
9 9 10 13 9 0 11 2 11 2
36 16 3 14 13 1 9 2 10 9 3 13 1 12 9 9 9 9 7 9 15 13 9 9 1 9 2 7 3 3 3 13 9 1 15 9 2
8 3 2 11 13 11 1 11 2
14 9 10 13 9 15 0 9 10 13 11 11 9 10 2
20 11 11 11 13 1 11 11 13 11 11 2 11 11 11 2 12 11 2 12 2
13 5 9 5 11 13 1 11 2 11 2 11 11 2
8 1 9 13 9 2 9 0 2
33 11 0 16 13 1 9 10 9 13 9 9 16 13 11 2 3 11 3 2 3 13 2 16 9 9 13 3 1 9 2 1 9 2
22 1 1 9 12 7 12 2 11 3 3 13 1 9 9 1 10 9 9 12 9 9 2
9 11 13 10 9 1 9 9 9 2
20 2 11 2 13 13 9 12 1 11 2 9 9 7 9 1 9 9 11 11 2
17 10 10 9 9 9 9 2 9 10 13 1 13 1 9 1 9 2
12 11 11 11 13 9 9 15 3 13 1 11 2
12 15 9 13 9 2 9 0 1 13 10 9 2
11 9 13 11 11 2 11 11 11 11 11 2
22 11 11 13 10 10 9 15 13 1 9 11 11 2 11 11 11 2 11 11 2 11 2
38 11 11 11 11 11 2 2 12 11 12 11 11 2 12 11 12 11 2 11 2 11 2 11 2 13 9 11 15 13 9 1 10 9 2 1 9 9 2
11 3 11 2 3 13 9 1 13 9 0 2
11 11 1 9 12 2 13 9 1 12 9 2
33 9 9 0 1 9 10 9 13 9 11 11 11 15 13 1 11 16 13 13 1 9 0 1 13 9 9 9 1 11 7 11 11 2
43 9 3 13 9 2 16 13 0 9 0 2 9 9 2 9 2 7 9 1 9 0 2 9 1 9 0 2 11 2 7 9 1 9 0 7 9 15 13 9 15 0 3 2
18 1 13 2 11 13 1 9 9 11 15 13 13 7 13 11 12 9 2
22 9 12 10 13 2 11 11 2 0 15 13 2 13 1 11 11 1 9 12 11 12 2
14 11 13 10 9 1 11 11 2 11 11 11 2 11 2
6 3 13 2 3 13 2
22 16 9 11 13 13 2 11 11 13 9 1 9 2 0 1 9 9 7 9 1 11 2
14 1 10 2 11 1 9 9 11 13 11 2 13 9 2
23 11 2 11 2 11 7 11 13 13 7 13 7 16 3 13 12 11 15 3 13 1 11 2
24 11 11 2 11 2 13 9 9 9 9 12 15 13 1 11 11 11 2 11 11 2 11 11 2
10 11 15 13 1 9 13 1 9 9 2
15 1 10 2 15 13 10 9 9 15 0 7 10 9 0 2
29 9 10 13 1 1 10 9 11 2 10 9 9 7 10 9 9 12 7 7 9 15 13 1 1 10 9 9 9 2
39 10 13 9 1 9 0 2 15 1 9 3 13 9 11 11 11 7 9 9 12 9 2 11 11 2 7 13 13 9 11 12 15 13 9 10 1 11 11 2
7 11 13 9 1 12 12 2
10 15 13 7 13 9 9 1 9 10 2
30 11 11 2 11 13 1 9 2 9 1 10 9 2 13 11 2 11 11 7 11 11 11 2 1 9 9 1 9 9 2
6 15 11 10 15 3 2
23 9 10 2 11 11 13 1 9 12 2 12 1 12 9 1 9 9 9 9 1 11 11 2
10 7 3 15 0 1 12 9 12 12 2
20 9 9 11 11 13 9 15 0 15 13 1 11 11 15 0 2 11 11 11 2
15 10 9 3 13 1 3 1 12 9 2 13 1 9 9 2
14 1 1 11 13 9 9 2 9 11 2 11 7 11 2
30 9 9 3 1 2 3 12 9 1 9 9 1 9 9 2 7 9 3 3 13 2 0 13 1 9 9 7 9 9 2
26 11 11 13 9 1 9 0 3 13 9 0 9 15 13 1 9 9 2 16 11 14 3 13 1 9 2
2 13 2
23 11 1 13 10 10 9 1 9 11 11 11 2 11 11 11 11 2 11 11 11 2 11 2
22 11 11 11 13 1 11 11 7 13 11 2 13 1 11 2 2 1 13 13 11 2 2
31 16 10 13 12 9 9 2 7 10 1 9 0 2 9 15 3 13 15 12 12 12 9 1 9 7 13 13 15 0 10 2
18 11 10 13 7 13 9 7 9 15 0 7 13 9 9 7 10 9 2
16 9 10 13 12 1 12 9 7 9 15 13 1 11 11 11 2
12 9 9 9 7 9 13 0 9 9 15 0 2
8 11 10 13 1 9 9 9 2
17 16 16 10 9 3 13 9 1 11 3 16 11 14 3 13 1 2
8 3 2 9 11 3 3 13 2
14 11 13 9 1 11 11 2 11 2 11 11 2 11 2
18 11 13 1 9 1 11 2 11 11 2 7 9 1 11 2 11 11 2
7 9 13 16 11 13 9 2
23 1 12 2 15 13 13 11 11 11 11 2 11 2 15 9 13 9 2 9 11 7 11 2
18 11 13 10 10 9 1 11 11 11 2 11 11 2 11 11 2 11 2
38 11 11 13 1 12 5 1 9 11 2 3 13 1 12 9 9 1 13 9 0 11 11 11 2 9 9 0 10 13 3 13 1 11 11 1 12 9 2
16 0 9 11 16 13 16 11 13 9 1 9 15 3 13 9 2
31 7 16 14 13 1 9 0 7 3 3 2 9 9 7 9 9 9 2 13 9 10 3 13 2 9 9 2 1 10 9 2
19 1 13 9 13 9 0 3 3 1 12 9 7 9 1 9 1 12 9 2
56 11 11 13 9 2 9 9 0 11 2 1 2 11 15 13 1 10 10 9 7 13 1 9 9 10 3 15 13 1 9 2 7 1 9 9 10 13 9 15 3 13 9 1 11 13 11 13 9 0 9 7 9 15 13 0 2
13 10 9 2 3 10 11 7 11 13 1 9 9 2
10 11 10 3 1 13 10 9 11 11 2
14 11 13 9 1 9 11 2 11 2 11 11 2 11 2
23 16 15 3 11 13 1 9 9 1 9 11 1 11 1 13 9 11 7 13 3 9 15 2
33 1 1 12 9 13 9 10 13 2 9 9 2 2 3 13 9 2 9 9 2 2 16 9 10 2 13 1 1 11 1 12 5 2
17 11 3 13 1 9 1 9 2 3 3 9 0 15 15 13 1 2
12 10 12 11 9 13 1 11 1 12 2 8 2
16 1 9 10 2 11 7 11 14 3 13 3 16 13 3 0 2
11 9 9 11 1 11 2 11 13 1 9 2
18 15 13 1 11 11 1 9 12 9 7 13 1 9 12 1 9 9 2
26 1 10 9 11 11 13 9 9 12 9 7 9 9 9 12 9 2 13 1 12 9 0 7 9 11 2
24 16 2 13 9 12 11 12 2 11 13 13 1 11 5 11 7 13 1 9 0 15 3 0 2
8 14 13 9 1 9 15 13 2
13 3 13 1 9 2 9 0 2 9 2 7 9 2
9 10 9 13 9 10 1 9 0 2
24 16 13 1 9 7 9 0 2 9 10 9 10 13 0 1 9 0 2 16 3 13 1 9 2
8 9 13 1 9 12 11 12 2
61 15 13 12 9 9 15 3 13 9 1 9 1 9 1 9 9 1 9 2 9 9 7 9 0 11 2 16 9 0 13 1 0 2 9 10 14 13 9 9 2 16 13 16 9 2 9 1 9 9 9 15 0 7 9 9 3 13 10 9 0 2
13 11 3 13 9 10 1 9 11 11 11 1 11 2
20 16 2 13 3 9 9 15 13 16 9 11 7 9 11 13 12 9 15 0 2
40 1 9 12 11 12 11 13 13 9 9 11 2 11 13 1 12 9 2 9 2 2 10 2 10 13 1 9 0 2 10 9 13 3 13 10 9 2 9 2 2
16 1 10 2 15 13 13 11 11 11 10 15 1 13 9 0 2
27 1 9 11 11 15 13 1 9 11 7 11 2 7 1 9 15 13 3 0 7 12 9 13 0 2 0 2
10 11 2 2 13 10 10 9 0 11 2
16 3 11 3 15 3 13 1 11 7 11 15 3 13 9 9 2
11 11 3 13 9 2 11 0 0 1 11 2
22 11 13 13 9 9 12 9 1 9 11 2 11 11 11 11 15 13 13 12 11 12 2
27 16 0 9 11 16 9 9 10 2 16 15 13 1 1 9 2 16 3 15 3 13 1 11 16 9 10 2
10 16 9 9 1 9 7 9 1 9 2
51 9 9 11 14 3 13 1 9 9 2 7 3 13 1 12 9 1 9 0 2 1 9 11 11 11 9 11 11 13 9 2 9 9 11 1 2 9 2 9 15 13 13 2 7 2 9 2 9 0 2 2
11 15 13 13 2 13 2 9 9 9 10 2
30 16 14 9 0 1 13 11 11 11 16 15 3 13 12 9 1 13 9 9 10 2 14 0 3 9 11 11 11 13 2
33 11 3 13 1 9 9 0 1 9 9 9 2 9 2 2 16 3 13 1 9 2 9 10 2 3 9 2 1 9 9 1 9 2
14 16 2 9 0 3 13 7 3 13 1 9 9 11 2
7 3 9 7 9 15 13 2
14 11 1 9 9 2 1 9 9 2 9 7 1 9 2
34 13 9 11 11 11 11 2 11 2 1 11 11 11 2 11 2 2 11 9 11 11 13 9 9 9 2 12 9 2 10 12 9 12 2
18 11 13 12 9 10 13 9 12 2 12 1 9 12 9 0 1 11 2
14 7 3 13 13 9 11 15 13 1 11 11 1 9 2
15 10 9 2 9 9 15 0 2 11 11 2 13 9 11 2
11 3 13 11 13 9 1 9 9 9 9 2
32 9 1 9 11 2 15 13 1 13 9 2 3 13 9 0 9 1 9 2 15 13 9 9 3 13 2 16 3 13 9 0 2
14 11 13 9 1 11 11 2 11 2 11 11 2 11 2
20 16 15 13 9 15 13 1 9 9 10 2 16 14 13 9 13 11 11 11 2
8 11 10 13 1 9 9 11 2
13 15 0 13 9 1 9 11 15 13 1 9 9 2
48 11 10 13 1 11 2 11 11 2 11 11 1 9 9 2 11 11 2 11 2 11 11 1 9 9 2 11 11 2 11 2 11 11 1 9 9 7 11 11 2 11 2 11 11 1 9 9 2
9 11 13 9 15 13 3 16 9 2
18 11 13 10 9 15 13 1 11 11 2 11 11 2 11 11 2 11 2
7 1 9 1 9 11 11 2
26 9 1 11 11 11 1 11 11 7 9 2 9 13 9 11 7 9 3 1 11 13 13 9 1 11 2
8 9 10 1 13 1 9 11 2
27 9 2 9 13 9 0 13 9 0 7 0 15 13 9 2 9 9 1 9 9 2 9 2 7 9 0 2
15 11 13 10 9 9 13 0 15 13 1 9 11 11 11 2
6 9 15 13 11 11 2
13 15 3 13 1 11 11 11 1 9 12 1 12 2
47 9 9 3 13 9 11 11 12 1 13 16 11 11 12 14 9 2 13 9 11 2 11 2 16 10 3 13 9 11 16 11 11 12 13 9 15 13 16 14 3 13 2 16 1 13 9 2
40 9 2 9 11 2 11 13 9 9 9 15 13 1 9 9 7 9 1 13 9 9 16 9 13 1 10 9 9 7 9 1 9 15 0 1 13 9 9 9 2
12 11 3 13 13 11 7 13 13 13 9 9 2
15 13 1 9 11 1 1 9 7 3 13 9 9 11 11 2
14 1 9 12 11 12 2 9 10 13 9 1 12 9 2
17 9 2 11 9 2 7 9 2 11 9 2 10 13 9 1 11 2
14 3 11 7 11 3 13 1 9 3 3 9 1 15 2
8 14 3 0 13 0 1 9 2
11 9 10 13 9 9 12 9 5 12 2 2
5 9 1 9 12 2
2 15 2
15 11 9 3 15 13 1 11 2 1 9 9 0 7 9 2
24 11 11 11 2 2 13 9 0 12 1 11 11 7 13 11 2 1 9 9 11 11 2 11 2
22 1 9 11 7 9 0 11 2 11 13 9 0 1 9 2 9 9 0 7 9 0 2
41 9 2 3 0 9 13 9 1 13 9 2 14 0 16 13 9 9 7 9 9 1 11 7 1 9 9 11 1 11 7 11 3 13 1 9 9 9 7 1 0 2
29 11 11 11 2 11 11 2 11 11 2 13 9 11 2 11 11 2 2 16 15 13 1 14 13 9 9 3 13 2
13 1 9 12 13 3 13 11 11 11 2 11 2 2
20 11 11 13 10 10 11 15 13 1 11 11 2 11 2 11 2 11 2 11 2
30 11 3 1 10 13 9 9 11 2 15 7 13 13 1 11 1 9 2 9 0 16 11 13 11 3 13 9 9 15 2
16 11 11 2 11 2 13 9 9 1 11 1 9 9 7 9 2
29 1 9 12 2 11 2 11 11 11 13 1 9 1 9 0 15 13 1 9 9 7 9 11 11 2 1 9 11 2
26 1 9 1 11 11 11 10 2 11 13 1 10 10 9 11 2 11 11 2 13 9 15 13 13 9 2
24 12 16 15 14 13 9 2 16 13 15 1 9 2 16 3 10 11 13 1 1 9 1 9 2
23 11 11 1 11 13 1 9 9 9 11 9 11 12 2 12 2 3 1 9 12 11 12 2
19 1 12 9 13 9 1 9 2 10 11 7 11 3 13 9 9 1 9 2
8 11 13 9 15 13 9 9 2
20 11 13 10 9 1 11 11 15 13 9 1 11 11 2 11 11 11 2 11 2
27 1 9 10 9 1 9 11 11 2 15 13 1 9 11 11 1 11 11 2 3 3 13 1 9 9 10 2
34 1 9 10 2 9 11 11 11 9 11 11 13 9 11 15 3 0 7 13 9 11 13 0 7 13 9 13 9 13 10 2 9 9 2
17 9 9 10 13 1 11 11 11 2 13 9 9 11 0 1 11 2
12 5 11 11 5 11 2 11 2 11 2 11 2
61 11 11 11 11 11 2 2 13 10 9 13 11 15 13 0 16 13 1 9 0 1 11 11 11 2 12 2 2 11 11 2 12 2 2 11 11 2 12 2 2 11 11 11 11 11 2 12 2 2 11 11 2 12 2 7 11 11 2 12 2 2
18 16 0 11 13 12 9 2 9 2 13 10 9 9 9 7 13 9 2
13 9 10 14 3 13 16 3 13 13 1 0 0 2
30 9 15 0 9 9 7 11 2 13 1 9 1 9 15 0 2 3 0 13 2 7 3 9 1 9 0 7 9 0 2
11 9 10 13 1 0 1 11 11 7 11 2
18 9 13 9 13 11 11 11 11 2 11 11 11 2 1 12 11 12 2
26 2 16 13 9 0 2 9 1 12 9 13 1 9 1 9 9 2 2 13 9 11 11 11 2 11 2
37 9 2 9 0 13 9 2 9 13 1 9 12 2 12 9 2 13 1 9 9 2 13 0 1 12 9 2 0 2 13 0 7 13 9 1 9 2
27 10 9 11 11 3 3 13 1 10 9 1 9 1 9 9 1 9 9 9 11 7 9 9 11 1 9 2
59 9 12 2 11 11 2 11 9 12 2 11 11 11 2 11 9 12 2 11 11 11 2 11 2 11 11 11 5 5 9 12 5 5 9 10 2 15 3 13 1 9 12 11 12 2 13 9 12 9 7 12 11 2 11 9 1 9 12 2
21 9 0 1 9 9 0 13 9 2 9 2 9 14 0 9 7 9 9 15 0 2
42 1 11 11 11 11 13 1 9 11 2 9 9 9 3 13 1 9 9 11 11 11 15 13 11 2 11 3 13 13 9 11 13 11 11 11 16 11 13 9 1 11 2
20 1 9 15 0 10 2 9 13 2 16 3 1 9 0 9 13 1 9 9 2
29 11 11 11 11 13 13 9 9 11 11 2 15 3 13 9 11 1 9 9 11 11 7 11 11 1 9 14 13 2
40 11 11 15 9 12 2 5 13 12 9 9 10 1 9 9 1 9 9 7 13 12 9 9 1 11 2 1 9 9 11 11 11 11 11 11 7 11 11 11 2
33 16 9 13 1 9 2 9 1 3 0 2 7 3 0 1 15 11 12 2 2 16 9 11 11 11 7 9 1 9 2 9 0 2
36 1 9 9 2 10 9 1 9 11 11 13 7 13 3 11 11 2 16 9 10 10 9 10 15 1 9 1 9 15 0 13 1 0 9 9 2
9 15 3 13 1 9 11 1 9 2
14 11 13 9 1 11 11 2 11 2 11 11 2 11 2
10 11 2 11 11 2 11 2 11 12 2
20 1 9 11 3 13 9 9 9 11 11 2 1 1 12 2 12 9 10 9 2
26 1 9 11 2 11 9 13 9 9 12 2 12 9 13 9 1 9 9 9 12 1 9 12 2 9 2
15 9 13 1 12 9 15 13 10 9 9 9 12 2 12 2
21 11 11 13 10 10 9 15 13 1 11 11 2 11 11 11 2 11 11 2 11 2
21 15 9 12 1 12 9 9 2 9 15 13 9 11 10 2 9 13 11 7 11 2
10 16 10 9 0 11 11 13 11 11 2
37 1 9 12 11 12 2 1 12 9 1 11 13 2 2 1 10 9 9 1 11 11 11 9 11 9 2 11 2 9 9 11 11 11 13 9 13 2
11 15 3 13 1 9 0 1 11 7 11 2
24 1 9 2 9 0 9 9 11 2 10 9 9 13 13 9 15 3 13 1 9 9 7 9 2
21 1 12 1 12 9 9 0 11 13 1 9 10 13 9 1 11 11 7 11 11 2
52 15 13 2 2 3 15 13 10 9 9 0 1 9 2 2 11 11 10 13 11 13 10 9 3 2 0 15 13 9 11 2 2 11 2 2 11 2 5 2 11 2 12 9 2 2 11 11 2 12 2 2 2
14 9 9 15 13 1 9 9 7 9 9 14 3 13 2
11 1 9 10 2 13 9 1 13 9 10 2
22 9 9 10 1 9 13 1 11 2 16 16 9 9 13 9 9 0 3 13 1 11 2
19 9 0 1 9 1 11 1 9 9 9 2 1 9 9 13 1 11 11 2
14 13 1 11 11 2 7 13 1 11 11 7 11 11 2
57 1 9 0 9 11 3 13 9 9 1 9 9 11 2 9 9 0 1 9 9 2 7 9 9 15 13 1 1 9 11 2 11 9 11 3 0 1 9 9 9 2 15 9 13 1 9 2 9 9 1 9 9 11 7 9 0 2
4 0 9 0 2
9 1 0 15 13 7 14 3 13 2
17 11 13 10 9 1 9 11 2 9 9 11 2 11 2 9 11 2
16 16 9 9 13 0 2 16 9 9 9 9 10 3 13 9 2
45 1 9 12 2 15 13 9 2 11 11 2 15 1 9 9 3 13 11 11 2 2 11 3 13 9 1 9 2 9 11 0 2 1 0 2 11 2 11 2 11 2 11 7 11 2
39 11 11 14 3 2 16 9 9 0 9 11 15 13 9 0 13 9 9 9 0 1 13 16 13 9 7 9 15 3 0 3 1 13 9 2 3 1 9 2
18 16 11 15 13 13 2 13 7 13 9 2 9 15 13 1 11 10 2
49 16 10 9 11 2 11 11 2 13 13 9 11 1 11 1 9 12 11 5 12 9 2 1 9 11 11 9 9 11 11 10 3 0 2 13 1 11 2 10 9 1 9 9 11 2 1 1 11 2
8 11 11 11 7 9 1 9 2
21 9 10 2 11 11 9 1 11 2 11 11 12 11 2 12 11 2 11 2 11 2
24 9 9 3 13 1 13 9 1 9 2 7 3 13 9 2 7 1 13 9 1 9 0 9 2
14 11 13 1 12 9 10 13 11 2 13 1 11 11 2
20 16 9 0 1 15 11 12 2 9 11 13 1 10 9 9 1 9 11 11 2
12 9 10 13 9 1 11 11 11 12 1 9 2
35 9 12 9 1 11 2 2 11 2 11 11 2 15 13 1 9 12 2 13 1 10 10 9 0 11 11 1 12 9 2 12 2 12 2 2
27 11 11 2 7 11 11 11 2 13 10 9 9 13 9 9 0 15 13 1 9 9 7 9 0 1 9 2
33 16 3 2 10 9 9 9 7 9 0 1 9 1 9 2 9 11 13 1 13 1 0 2 9 3 1 9 2 9 1 11 13 2
33 11 13 1 9 9 7 9 2 9 1 9 11 12 1 9 12 2 16 15 13 9 1 9 16 13 9 0 2 16 11 13 2 2
21 9 14 13 3 13 9 1 9 9 2 9 9 14 13 3 13 13 1 9 13 2
13 11 11 13 3 13 9 9 10 16 13 9 9 2
64 9 9 11 7 11 3 13 1 9 9 1 9 1 9 11 7 9 11 2 12 5 11 11 2 12 5 9 2 11 7 11 2 5 9 2 11 2 11 2 2 11 2 5 9 2 11 2 2 7 9 5 9 2 11 2 2 7 9 1 9 11 13 9 2
20 9 9 1 12 9 2 15 0 1 12 2 12 9 2 9 0 2 9 2 2
61 7 12 9 13 1 9 12 9 9 0 2 9 9 9 9 0 13 9 0 9 0 9 10 2 9 0 2 0 7 3 12 9 13 1 9 0 2 9 10 13 9 1 9 12 2 3 2 7 12 9 13 9 2 9 10 14 13 1 9 0 2
24 15 13 1 9 0 1 9 12 2 13 1 12 9 9 7 13 9 1 9 11 2 11 11 2
5 10 9 13 9 2
18 1 9 10 9 3 13 7 3 0 1 13 9 16 3 13 1 9 2
23 11 11 2 11 11 2 11 2 13 9 9 1 11 11 7 11 11 15 13 1 11 11 2
23 9 0 9 1 12 2 12 13 9 9 9 11 2 1 9 11 12 1 11 11 15 13 2
13 1 9 11 3 11 13 1 9 7 9 2 2 2
19 1 10 9 3 13 16 1 9 10 14 13 9 1 13 1 1 9 0 2
8 7 9 13 11 3 13 0 2
15 3 13 10 9 9 12 9 11 9 2 9 1 9 12 2
19 9 10 11 11 9 11 11 13 1 12 11 15 13 1 9 1 11 11 2
15 11 13 9 1 11 11 11 2 11 2 11 11 2 11 2
20 15 15 3 13 16 11 3 13 13 1 13 9 9 12 9 1 11 11 12 2
66 11 11 13 9 9 9 11 9 9 11 11 11 9 9 9 11 11 11 11 2 13 9 11 11 2 11 13 10 10 9 15 3 13 7 9 15 3 13 2 0 1 9 2 0 1 9 2 0 1 9 14 3 13 2 13 9 11 2 15 3 12 14 13 15 12 2
12 7 1 0 13 9 9 0 2 3 11 11 2
20 3 11 11 13 13 12 9 15 13 1 9 11 1 9 12 2 12 1 11 2
23 11 2 9 15 13 1 11 11 13 11 2 11 2 11 2 11 2 11 2 11 7 11 2
15 11 13 9 15 13 1 11 11 2 11 2 11 2 11 2
20 8 2 11 11 13 1 10 9 9 15 13 1 7 9 9 1 9 11 11 2
7 11 10 3 13 9 11 2
14 9 1 9 0 13 9 0 15 3 3 13 9 9 2
24 1 10 3 2 9 11 3 13 9 2 7 3 11 13 1 10 10 9 0 1 11 11 11 2
29 11 2 2 9 2 9 7 9 2 13 9 15 13 13 9 1 9 2 13 13 2 3 9 2 9 2 7 9 2
27 9 11 15 13 3 14 3 13 9 9 16 0 2 0 3 13 1 9 2 9 9 0 1 10 9 9 2
14 11 13 9 1 11 11 2 11 2 11 11 2 11 2
11 1 9 11 3 13 9 0 10 1 9 2
19 3 3 13 9 13 1 9 9 11 1 11 11 1 9 11 11 12 10 2
20 1 12 9 12 3 13 9 9 16 11 11 3 13 9 11 7 13 1 9 2
84 9 2 15 13 1 2 11 2 7 11 2 11 3 13 12 9 1 9 1 11 2 11 2 9 9 2 11 2 11 7 11 13 1 9 11 2 11 2 11 2 11 13 11 14 13 11 2 11 9 2 16 9 13 15 13 9 13 9 2 16 16 11 13 2 11 2 11 13 16 13 9 2 9 13 3 2 3 1 9 2 9 15 0 2
14 12 9 9 13 2 1 9 9 2 9 7 9 11 2
8 10 9 2 3 13 9 11 2
30 1 1 11 11 7 11 11 2 9 11 13 1 12 9 1 12 9 16 1 1 9 11 13 1 12 3 1 12 9 2
9 1 2 1 9 9 1 9 10 2
14 16 13 11 1 11 2 2 9 15 13 1 15 10 2
10 9 2 9 9 9 11 13 1 13 2
23 9 9 1 9 9 2 9 13 1 9 12 9 2 7 9 10 13 1 9 1 13 9 2
16 1 9 9 11 11 11 11 9 0 1 9 2 9 7 11 2
8 11 9 10 14 13 9 9 2
12 9 9 10 13 9 11 11 2 10 9 11 2
28 1 9 9 9 9 12 2 11 13 16 11 3 13 12 5 1 9 11 11 1 10 9 2 13 9 9 11 2
20 11 11 13 9 0 0 11 2 11 11 1 9 0 9 15 13 1 9 9 2
21 11 2 12 13 9 9 15 3 0 1 9 11 3 13 9 9 9 1 9 11 2
27 9 13 9 1 11 11 7 11 11 2 11 2 11 11 2 13 1 9 9 12 2 7 13 1 10 9 2
5 9 15 13 0 2
12 11 11 0 9 13 1 11 1 11 11 12 2
20 13 1 9 9 11 9 7 11 13 10 11 11 13 0 1 9 9 1 0 2
9 1 10 2 13 3 9 9 11 2
15 11 13 9 9 1 9 11 3 13 9 9 1 9 10 2
15 11 11 13 9 9 13 12 2 12 9 11 1 9 12 2
8 3 11 11 13 1 11 11 2
30 11 9 10 3 13 1 9 11 12 2 16 0 9 9 1 9 1 11 11 11 2 16 13 3 1 9 12 1 12 2
23 9 2 11 11 13 9 11 7 13 9 2 9 1 11 16 9 3 13 16 15 13 0 2
33 11 11 10 1 0 13 1 10 9 0 1 9 11 11 2 11 2 10 9 9 12 15 13 1 11 11 11 1 9 10 11 11 2
21 15 3 9 9 9 11 11 2 11 11 11 2 7 11 11 1 11 9 11 11 2
16 1 10 9 2 15 3 14 13 3 1 12 9 1 12 9 2
17 11 11 7 11 11 13 9 0 9 9 1 9 15 13 1 11 2
47 16 16 9 15 13 7 0 9 3 9 0 11 15 14 13 9 10 13 9 0 1 9 10 2 16 3 15 3 13 13 9 11 15 13 9 10 16 13 9 2 9 9 9 11 11 10 2
58 9 9 0 1 11 1 0 13 11 11 2 11 11 2 11 11 11 2 11 11 11 2 7 9 11 15 13 1 9 11 2 11 11 2 11 11 11 2 7 11 11 11 15 13 1 9 11 2 11 11 7 11 11 1 9 11 11 2
9 15 3 13 13 9 9 11 3 2
16 9 10 13 12 1 12 12 12 9 15 13 1 11 11 11 2
12 11 11 2 16 9 13 2 13 1 9 9 2
21 9 10 13 1 9 9 11 11 2 7 9 13 9 1 9 2 9 2 7 9 2
42 11 0 9 13 1 11 12 1 11 13 2 1 9 15 3 13 1 9 11 11 12 7 11 11 12 16 15 12 9 13 16 9 9 0 1 9 11 12 7 3 13 2
18 16 11 2 11 2 11 13 2 3 15 13 9 11 2 7 9 11 2
42 9 11 15 12 9 1 11 11 3 13 1 9 2 9 2 11 11 2 12 2 12 2 11 11 2 12 2 12 2 2 15 1 9 3 2 3 13 2 9 10 9 2
18 9 9 12 13 9 9 2 13 1 11 11 2 11 2 9 9 9 2
12 1 12 9 13 9 1 9 11 13 9 11 2
34 0 9 9 13 1 11 11 2 15 13 1 9 1 2 12 1 9 0 11 11 15 13 1 9 1 2 12 2 16 11 13 9 10 2
13 16 9 15 8 13 1 9 10 3 0 7 0 2
8 11 11 13 9 1 12 9 2
25 1 9 12 2 15 13 1 11 1 13 0 1 11 11 7 13 9 11 2 11 11 7 11 11 2
13 9 9 3 13 13 9 7 9 1 9 7 9 2
17 1 9 12 2 9 10 13 9 9 1 12 9 7 12 9 9 2
12 11 3 0 1 9 7 13 9 1 9 10 2
35 16 9 2 9 11 11 0 1 0 13 9 2 9 1 9 0 2 15 3 0 1 9 9 2 9 9 2 9 9 9 2 7 9 9 2
54 9 9 10 13 1 9 13 10 9 9 0 2 13 1 1 11 2 11 2 11 2 7 11 2 11 9 1 9 12 13 9 12 9 2 3 12 9 9 9 9 12 11 2 2 9 15 14 0 1 10 9 9 11 2
9 1 9 11 13 16 11 3 13 2
29 1 9 9 9 0 11 11 11 2 11 11 11 13 11 11 7 11 11 1 12 2 7 13 9 9 12 9 3 2
14 11 13 9 1 9 11 2 11 2 11 11 2 11 2
12 11 10 13 1 9 11 11 15 13 11 11 2
25 9 1 9 9 0 11 2 1 9 9 15 13 9 13 9 1 9 9 1 13 9 9 9 9 2
58 9 10 13 1 0 1 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 7 11 11 1 15 13 1 9 11 2 12 11 12 1 9 9 11 1 9 9 13 11 11 11 11 11 11 11 15 13 9 1 11 2
17 11 9 9 11 11 13 1 13 1 12 9 15 13 13 12 9 2
32 11 13 9 0 11 7 13 9 0 7 9 0 1 12 9 1 10 9 2 3 9 0 1 12 9 7 9 9 7 9 0 2
9 11 13 1 11 11 7 11 11 2
14 9 7 9 1 11 13 9 1 13 9 1 9 13 2
9 14 15 15 13 15 11 13 11 2
16 10 9 3 13 9 2 9 0 7 3 13 1 13 1 9 2
8 11 12 3 13 1 11 11 2
58 1 13 9 1 9 9 11 1 9 2 9 11 2 16 1 9 12 11 13 10 9 0 1 9 9 9 15 13 1 9 2 2 11 11 11 11 2 1 9 12 2 9 10 13 16 9 9 0 2 7 3 3 13 9 2 9 9 2
54 1 9 12 2 1 11 11 13 1 9 9 1 9 9 15 0 11 11 2 11 11 13 9 0 2 11 2 11 11 2 9 11 2 11 2 11 2 2 16 11 11 11 11 11 2 11 2 13 9 10 1 11 11 2
21 1 9 2 9 0 2 11 13 9 15 3 0 1 9 9 1 13 9 1 13 2
29 13 9 11 11 13 11 11 11 11 11 1 9 12 11 2 12 2 11 3 0 1 11 7 13 13 9 1 11 2
13 1 13 2 15 13 11 11 11 16 9 10 13 2
31 11 7 11 13 10 9 9 9 2 9 15 13 1 12 9 12 1 11 7 13 1 9 2 9 10 13 1 11 2 11 2
17 11 9 0 9 13 11 11 11 11 11 15 13 1 9 9 9 2
40 11 9 10 3 13 1 9 9 2 1 1 9 7 0 2 15 3 13 9 0 1 9 7 9 7 9 2 1 13 9 2 9 13 2 9 9 9 5 9 2
27 11 11 2 13 1 9 0 11 11 2 13 9 9 9 2 0 1 9 7 9 2 15 13 1 11 11 2
12 1 9 10 2 15 13 9 11 11 11 11 2
23 13 11 11 11 2 11 1 9 9 9 1 9 0 2 2 15 3 9 13 13 1 9 2
16 1 9 12 2 9 10 13 9 1 12 9 7 12 9 9 2
12 11 13 9 15 13 12 5 1 9 9 11 2
26 11 9 9 7 9 11 3 13 10 9 15 0 2 16 1 0 9 2 16 9 1 9 13 14 0 2
14 11 12 13 9 12 1 9 9 9 11 11 2 11 2
15 3 13 1 9 2 13 9 2 2 11 2 13 9 0 2
22 11 3 13 10 9 2 1 7 1 9 2 7 10 9 1 15 13 9 15 14 0 2
9 11 10 13 9 12 9 1 9 2
12 9 10 13 1 9 2 9 11 15 0 13 2
24 1 9 2 3 1 12 5 9 2 9 13 3 0 1 9 2 3 10 9 9 3 13 3 2
21 7 9 10 3 13 0 1 9 9 11 1 9 1 12 16 3 13 1 9 0 2
33 9 9 2 3 13 1 9 11 13 1 9 12 9 7 13 1 11 11 11 11 11 2 11 2 11 2 2 9 9 1 11 11 2
24 11 9 9 9 13 1 13 9 10 1 2 9 0 2 13 1 9 15 13 9 15 3 13 2
10 9 10 13 1 11 2 11 2 11 2
11 11 11 11 2 11 3 13 1 9 9 2
34 1 9 12 2 9 10 13 9 9 1 12 9 7 13 9 9 12 12 2 2 9 10 13 9 9 9 12 2 12 9 5 12 2 2
16 11 11 13 9 1 11 11 11 2 11 2 11 11 2 11 2
29 11 13 16 9 0 1 9 9 9 13 1 13 9 2 7 9 1 13 2 12 9 3 0 2 1 0 2 9 2
32 2 12 2 11 13 1 9 11 11 2 12 1 11 11 11 11 12 5 11 11 1 13 10 11 11 1 9 11 11 9 11 2
20 11 2 2 13 9 15 13 1 1 9 9 2 9 13 12 9 2 12 2 2
15 9 10 1 1 2 11 11 11 13 10 9 0 2 1 2
22 11 13 9 9 9 0 2 0 9 9 16 9 7 9 2 7 9 2 7 9 2 2
11 16 15 3 13 2 3 3 13 11 13 2
15 13 1 11 1 9 12 5 7 13 1 12 2 12 2 2
10 13 1 0 9 2 9 15 15 13 2
29 1 9 2 10 9 13 1 9 2 9 2 9 2 9 9 2 7 9 2 9 9 0 3 1 9 2 9 0 2
19 9 10 1 12 11 12 13 9 0 15 13 9 2 9 0 1 9 11 2
9 11 10 3 13 1 9 0 0 2
28 11 2 9 10 2 9 1 9 7 9 9 9 3 13 9 10 9 13 0 1 9 2 9 1 9 9 0 2
15 9 9 3 12 9 1 12 9 2 7 3 13 12 9 2
22 11 11 7 11 3 13 11 1 9 2 7 1 9 12 2 15 13 9 0 11 11 2
19 15 13 1 11 7 1 11 2 13 9 12 1 9 12 9 1 9 9 2
7 9 15 3 15 13 9 2
24 3 2 7 13 1 9 11 7 11 2 1 9 11 13 1 11 2 7 1 9 11 1 11 2
18 1 9 9 11 0 13 13 9 2 9 9 7 9 2 9 9 0 2
25 12 9 10 13 1 0 2 11 9 13 9 2 13 9 2 7 13 9 1 10 11 1 9 10 2
15 1 9 9 15 13 2 13 14 7 13 9 9 13 9 2
6 11 9 13 13 9 2
9 9 10 13 9 12 1 9 12 2
16 11 13 16 9 10 3 3 3 9 1 9 9 9 7 9 2
24 11 13 10 10 9 0 1 9 10 2 16 9 15 3 13 0 7 9 9 1 9 11 11 2
19 11 13 10 10 9 15 13 1 9 11 2 11 11 2 11 11 11 2 11
21 11 11 11 11 13 10 9 0 15 13 1 9 11 11 2 11 11 2 11 11 2
24 1 9 12 12 12 2 12 2 12 2 9 11 2 11 11 2 11 11 11 13 9 1 11 2
32 11 11 13 9 9 1 9 9 2 11 11 11 2 11 3 13 9 0 1 9 11 11 11 12 7 13 12 9 0 1 9 2
21 1 9 9 11 2 9 10 9 1 13 13 9 0 9 3 3 13 1 9 0 2
32 15 13 1 11 11 1 9 2 11 11 2 15 3 10 9 7 9 11 11 2 11 11 2 11 2 2 1 13 9 1 9 2
39 11 9 10 13 11 11 2 9 11 2 11 11 2 15 9 13 7 13 13 9 11 1 9 11 11 11 12 2 11 14 13 16 9 12 9 13 3 9 2
11 3 11 3 14 3 3 13 9 1 11 2
31 1 9 9 9 1 11 11 12 11 12 13 16 15 1 11 11 13 1 9 9 11 11 15 1 0 13 1 12 11 12 2
14 12 9 9 10 13 9 15 3 0 1 1 9 9 2
10 3 16 15 14 3 13 1 9 10 2
14 9 13 9 1 9 11 2 9 2 9 0 2 9 2
13 14 13 9 0 1 13 0 13 13 9 9 0 2
11 11 1 9 12 2 13 9 1 12 9 2
20 1 11 11 11 9 12 13 9 9 1 12 9 2 3 11 11 7 11 11 2
21 9 2 0 2 1 15 13 1 9 9 2 9 10 2 14 9 15 0 7 14 2
49 9 12 12 5 12 1 11 11 15 13 1 9 9 1 13 12 9 2 12 9 1 11 11 11 7 12 9 1 11 11 2 7 15 13 1 11 2 11 1 9 0 1 9 12 5 12 1 11 2
12 11 11 13 9 11 11 0 1 11 2 11 2
23 1 9 12 11 12 2 15 13 9 11 3 9 13 9 3 9 13 1 13 2 11 11 2
13 3 3 7 9 9 13 0 1 7 13 9 10 2
28 1 9 9 13 15 0 1 11 11 11 7 9 10 9 1 9 12 1 9 2 10 9 11 3 13 9 10 2
13 13 9 12 2 15 13 9 9 9 9 2 9 2
34 1 9 12 2 9 12 13 11 11 7 13 1 3 2 3 1 11 11 2 11 11 2 11 11 2 7 11 11 15 13 9 3 9 2
8 9 10 13 10 9 9 9 2
18 11 11 5 11 11 11 13 10 9 13 9 5 9 5 9 1 11 2
8 11 10 13 9 1 9 9 2
17 9 11 2 11 2 7 11 11 1 11 11 13 9 10 2 10 2
43 9 9 9 2 13 9 9 9 2 1 12 9 10 13 14 3 1 12 9 15 3 13 1 9 2 9 9 9 7 9 2 7 10 9 0 9 15 3 13 7 13 9 2
8 9 1 9 11 7 11 11 2
41 9 9 10 3 13 1 10 9 9 9 2 11 11 11 13 9 11 2 11 11 2 15 13 1 11 11 11 11 1 11 2 11 7 13 1 9 11 1 11 11 2
35 13 3 9 9 2 15 13 1 11 11 1 12 11 12 1 9 9 9 11 11 2 10 11 11 2 1 9 13 9 9 15 13 11 11 2
9 1 9 12 11 3 13 9 0 2
37 2 11 11 11 2 13 9 11 1 9 0 9 7 9 9 11 11 2 11 11 11 11 2 10 9 12 9 13 0 1 9 9 9 12 11 12 2
8 11 10 13 9 1 12 5 2
21 10 9 13 1 9 11 2 1 12 9 9 11 11 7 9 9 11 11 7 11 2
36 9 10 13 12 9 15 14 13 1 9 12 15 2 11 11 2 11 11 11 11 11 2 9 10 13 1 5 12 1 11 12 16 9 0 9 2
26 11 11 3 13 1 9 12 2 12 16 11 11 11 3 13 1 11 11 16 3 9 9 13 1 1 2
8 9 9 0 12 1 11 11 2
21 11 2 11 2 9 0 9 13 1 11 2 11 11 2 9 9 11 11 2 11 2
14 15 13 9 16 13 9 11 2 11 1 13 9 15 2
24 11 11 13 10 10 9 15 13 1 9 11 2 11 2 11 11 11 2 9 11 11 2 11 2
15 15 13 1 0 13 9 1 9 11 1 10 9 15 0 2
71 11 12 3 13 9 13 10 9 11 11 15 13 2 1 9 9 12 11 11 15 14 13 1 11 11 9 12 11 11 9 12 2 1 9 9 9 12 1 12 9 15 13 2 7 9 11 11 2 16 13 12 2 12 2 12 2 12 7 12 9 9 2 1 11 11 11 1 9 9 12 2
43 13 3 9 1 9 9 7 9 14 13 2 7 16 15 0 2 15 3 14 13 9 9 2 9 1 9 15 13 2 7 9 9 0 13 0 2 13 11 13 10 9 9 2
15 14 2 9 2 0 15 1 15 2 14 3 0 1 9 2
36 9 9 2 11 13 16 11 16 13 0 1 9 9 9 12 2 16 15 0 1 0 13 9 7 3 13 10 9 15 3 13 1 9 9 12 2
24 1 9 2 9 7 9 9 9 15 13 9 2 0 1 9 2 3 3 3 13 1 9 9 2
21 15 13 1 11 11 16 9 13 11 11 2 1 9 12 2 1 9 12 9 15 2
21 1 7 10 1 9 11 11 2 9 11 3 13 2 9 0 2 7 2 9 2 2
30 9 13 11 13 2 2 13 9 9 9 1 9 0 2 1 9 1 9 2 7 1 15 3 13 9 1 9 9 2 2
46 11 10 10 2 10 15 3 13 9 1 9 9 9 2 9 10 13 12 12 2 9 2 1 9 12 9 9 0 2 0 2 9 0 12 12 2 7 3 13 1 12 9 14 2 9 2
15 1 9 9 2 3 1 12 9 13 9 9 10 10 9 2
15 11 11 2 11 11 10 9 0 1 9 0 1 9 12 2
40 9 11 13 10 10 9 9 1 9 2 9 2 9 2 9 2 7 9 9 13 9 2 13 1 9 9 9 2 9 9 7 9 1 9 15 1 1 9 9 2
76 9 13 10 9 0 15 13 2 11 11 2 2 10 9 15 13 1 11 11 11 1 9 12 2 8 10 13 9 0 7 9 0 1 13 9 9 1 11 2 13 12 1 9 9 13 2 9 9 13 9 2 9 0 15 3 3 13 7 13 1 1 9 9 15 3 13 9 1 9 1 13 9 1 13 9 2
7 9 0 15 0 14 13 2
12 16 13 9 9 2 9 3 13 1 9 11 2
36 1 9 2 9 11 2 11 1 9 10 13 10 9 1 11 1 9 2 11 11 11 2 2 15 13 1 0 9 11 11 2 11 11 0 2 2
15 1 9 10 11 11 13 9 1 11 2 11 11 7 11 2
20 11 11 3 1 0 13 1 16 15 13 9 2 9 2 1 9 2 9 2 2
12 11 13 13 1 9 7 3 0 13 9 0 2
16 9 0 1 9 9 13 1 9 7 9 2 15 13 1 13 2
24 11 7 11 3 3 13 1 0 2 16 11 3 13 9 2 16 9 13 0 1 9 7 9 2
26 11 7 9 15 13 1 10 9 2 9 2 11 2 9 2 1 9 0 7 13 1 13 1 9 0 2
63 1 9 1 9 1 9 0 2 9 0 1 9 3 13 1 11 11 11 11 2 11 2 11 12 13 9 9 1 13 9 9 2 15 13 10 9 15 13 1 9 7 10 9 9 0 9 15 13 1 12 9 9 9 9 9 12 9 7 9 9 9 11 2
86 9 9 2 9 15 0 13 9 0 12 11 2 13 9 12 11 7 9 0 0 12 11 2 1 9 12 9 9 9 15 0 13 9 9 1 0 12 2 12 9 2 3 9 12 2 12 9 2 9 9 12 2 12 9 2 9 9 12 2 12 9 2 9 5 9 12 9 2 9 12 2 12 9 16 15 0 9 13 9 9 15 3 13 12 9 2
14 11 13 10 9 1 11 11 2 11 11 11 2 11 2
22 1 9 12 2 10 9 13 1 10 9 9 7 9 2 7 11 13 7 13 9 10 2
11 9 13 1 9 2 9 2 7 9 0 2
10 11 11 13 1 11 11 7 11 11 2
15 9 2 9 10 13 1 9 9 9 10 13 9 15 13 2
22 11 3 13 1 12 9 3 13 16 16 15 13 9 15 2 3 15 13 1 9 0 2
9 3 15 3 13 11 1 11 13 2
4 3 15 13 2
10 10 9 13 10 9 9 0 1 11 2
13 15 13 9 1 11 16 3 13 1 11 13 9 2
24 3 11 13 1 9 9 1 9 11 11 1 9 12 11 12 2 1 9 0 12 2 12 12 2
57 16 7 2 11 11 1 9 15 3 0 1 11 2 15 13 7 13 1 9 11 1 12 3 1 9 12 1 11 11 2 13 2 2 11 11 2 11 2 10 3 15 13 1 9 2 9 9 2 1 9 11 0 1 9 9 11 2
9 9 13 11 11 2 11 0 11 2
18 9 10 13 9 12 15 13 1 9 11 1 2 0 2 12 11 12 2
13 1 9 10 11 13 9 0 3 2 11 11 2 2
12 9 10 9 0 0 13 12 12 9 1 9 2
12 16 11 13 9 11 2 15 3 13 1 11 2
20 1 9 10 1 9 9 2 11 1 9 13 10 10 9 0 15 13 1 11 2
34 11 10 13 1 9 9 2 13 12 2 12 9 8 12 9 1 9 9 12 2 12 9 13 1 9 12 9 7 9 12 2 12 9 2
42 11 5 11 13 9 1 9 12 16 11 11 2 7 11 11 13 1 11 11 7 9 10 13 9 13 11 11 11 2 9 10 13 1 9 12 2 16 13 13 1 11 2
7 9 9 1 12 9 12 2
18 9 9 15 13 1 9 10 13 9 2 9 2 9 0 2 9 9 2
13 11 10 13 9 9 9 12 2 12 9 5 9 2
19 11 13 9 9 9 11 2 7 13 16 9 9 11 3 13 1 9 11 2
30 9 2 11 11 2 3 13 1 9 11 2 16 9 11 3 13 9 2 9 10 0 2 0 7 3 3 13 11 11 2
12 3 15 13 15 1 11 2 13 15 1 11 2
31 16 11 13 1 9 1 11 2 1 0 0 3 13 1 9 9 11 2 11 11 1 11 9 10 3 13 9 0 1 9 2
9 9 10 13 1 9 12 1 11 2
14 16 13 9 15 0 1 9 10 2 9 13 9 9 2
22 2 16 16 15 13 9 7 9 15 13 1 9 7 1 3 2 3 15 3 13 9 2
28 13 3 9 9 9 2 1 0 9 11 2 11 11 2 11 2 11 11 2 11 11 11 2 7 11 11 11 2
9 15 15 13 1 9 10 13 9 2
18 9 13 11 3 13 1 9 0 7 13 1 11 11 11 2 11 2 2
7 11 1 11 11 13 13 2
37 3 11 11 3 13 9 9 1 9 11 11 11 1 9 9 9 13 1 11 11 2 7 13 11 11 11 1 11 11 11 16 3 13 11 11 11 2
34 9 9 11 11 13 9 15 3 0 1 9 9 9 9 1 9 10 1 9 12 2 1 12 9 1 9 12 13 12 9 1 9 12 2
30 9 9 9 10 13 1 9 12 11 12 1 10 9 1 9 11 11 1 11 11 15 13 1 12 9 2 9 11 11 2
3 1 9 2
19 11 11 11 13 9 0 1 9 9 12 2 12 12 2 13 13 12 9 2
28 9 10 9 11 11 13 1 11 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 7 1 11 2
18 11 13 10 9 1 9 9 11 2 11 11 2 11 11 11 2 11 2
15 13 9 0 1 9 9 11 11 15 13 1 12 11 12 2
15 11 13 10 9 9 9 13 9 13 2 1 9 9 11 2
27 11 9 13 9 15 13 9 9 2 9 0 2 1 9 2 9 2 9 7 9 1 10 9 7 9 0 2
13 11 11 11 13 9 9 15 13 9 11 1 11 2
16 9 10 13 12 10 9 2 11 11 13 1 9 12 11 12 2
29 1 9 12 2 9 13 1 11 2 11 11 2 2 12 5 11 2 11 5 11 2 12 5 11 5 12 5 12 2
17 9 10 13 1 11 11 2 11 11 2 7 2 11 11 11 2 2
14 11 13 9 1 11 11 2 11 2 11 11 2 11 2
23 13 1 9 9 1 9 9 2 9 3 13 1 9 0 1 13 0 15 13 9 9 0 2
25 11 2 9 11 14 3 13 15 13 1 9 10 2 1 11 11 2 11 11 2 7 10 9 0 2
18 1 10 2 1 12 9 13 13 11 11 2 11 7 11 1 11 11 2
24 15 13 9 1 10 9 2 16 14 0 3 15 13 1 9 7 13 1 9 11 3 11 11 2
24 1 9 11 2 11 13 9 11 11 15 3 13 9 15 13 9 9 15 7 3 13 9 0 2
19 13 9 10 2 9 3 13 9 9 10 1 13 9 15 13 1 9 0 2
15 13 12 9 9 15 3 13 1 9 2 9 9 1 11 2
19 1 9 10 2 12 9 10 15 13 1 10 9 13 9 9 0 7 9 2
23 11 11 13 11 13 11 13 9 1 9 9 2 7 13 1 13 9 2 9 11 1 9 2
27 11 11 11 2 2 2 13 10 9 9 11 7 11 11 11 12 2 12 1 12 11 12 1 12 11 12 2
23 11 11 13 10 10 9 15 13 1 9 11 2 9 11 11 11 2 9 11 11 2 11 2
8 12 2 8 10 9 2 13 2
14 1 9 11 2 9 1 11 15 13 12 9 2 13 2
6 11 3 13 1 9 2
7 9 15 13 16 11 13 2
30 9 10 9 0 1 10 9 15 13 11 11 1 0 13 2 13 9 7 13 9 9 2 15 15 14 13 9 1 10 2
17 1 1 9 9 2 9 9 13 0 0 3 13 13 1 11 11 2
15 11 13 9 9 15 13 9 2 16 9 1 0 0 9 2
7 9 9 9 10 13 12 2
22 9 9 13 10 9 15 13 1 9 9 7 9 9 7 1 13 9 1 9 7 9 2
40 11 11 2 11 2 11 2 11 11 2 13 9 11 11 11 2 11 11 2 11 13 9 11 2 11 2 9 13 10 11 7 9 13 10 11 15 13 1 11 2
42 1 9 11 12 2 11 14 13 9 13 11 2 7 1 9 0 7 9 9 15 13 1 11 2 0 1 9 15 15 3 0 2 11 13 9 9 15 0 7 13 0 2
21 11 11 2 11 11 7 11 11 3 13 1 11 11 11 2 11 11 7 11 11 2
10 11 13 11 11 7 9 13 11 11 2
9 11 9 10 0 13 1 9 0 2
14 1 13 14 13 9 9 0 2 11 11 1 13 9 2
13 1 9 10 2 13 10 9 15 13 9 0 11 2
7 9 9 9 9 3 13 2
10 1 9 10 2 15 13 9 9 11 2
28 1 9 11 12 2 15 13 11 11 11 1 11 1 9 13 9 11 11 1 13 9 11 11 1 1 9 11 2
26 11 13 9 9 0 0 7 13 1 10 9 1 9 11 2 11 11 2 12 2 12 2 1 9 12 2
25 9 9 3 13 9 9 9 3 13 1 0 7 13 1 9 2 7 16 10 9 9 3 13 0 2
17 11 13 9 9 15 13 10 9 11 1 9 9 13 1 9 11 2
15 11 2 9 9 15 7 13 13 9 13 2 0 7 0 2
14 11 11 13 9 1 9 11 2 11 2 11 2 11 2
23 1 13 9 10 2 11 14 13 9 1 9 2 7 16 3 13 9 2 15 13 1 11 2
15 16 10 2 9 15 3 13 11 2 14 3 13 9 2 2
59 1 9 2 9 11 1 9 9 9 13 2 11 13 10 9 9 3 0 1 9 2 13 11 11 11 11 11 2 11 11 11 11 2 15 14 13 7 15 3 0 2 16 13 9 3 0 1 9 2 9 0 2 11 11 0 2 7 11 2
13 3 2 9 9 1 9 10 13 1 9 9 0 2
12 11 11 7 11 13 2 2 9 15 13 13 2
22 1 9 10 2 9 3 13 1 9 9 0 2 9 9 1 9 9 9 1 9 2 2
10 3 9 9 11 15 13 1 1 9 2
19 11 11 3 13 9 9 15 13 9 11 1 9 9 9 9 1 9 11 2
30 1 9 11 13 11 2 11 11 7 11 2 9 11 2 9 9 2 1 9 11 2 9 2 9 2 11 2 11 2 2
5 0 9 9 15 2
12 11 11 13 9 9 9 15 13 1 9 11 2
18 11 10 13 1 12 11 12 1 11 2 11 11 1 9 11 11 11 2
17 3 2 3 13 10 9 2 3 2 11 11 11 11 11 11 2 2
19 9 9 1 9 7 1 9 2 9 3 13 1 9 11 2 7 11 0 2
20 10 9 10 13 13 2 3 13 1 13 9 3 7 3 13 1 13 9 0 2
6 1 10 2 9 13 2
21 11 13 1 10 9 1 9 11 2 15 13 9 9 15 0 1 1 9 15 13 2
54 9 10 3 13 13 1 9 11 1 9 12 2 16 14 13 9 15 0 1 1 9 12 2 16 11 2 11 11 11 2 15 3 3 13 11 2 13 1 11 11 2 12 9 3 11 11 12 1 0 13 9 11 11 2
11 15 13 13 11 2 7 3 13 13 11 2
16 11 13 10 9 1 11 11 2 11 11 2 11 11 2 11 2
33 9 10 3 13 1 9 11 2 1 9 9 1 9 9 2 9 7 9 0 2 0 15 13 9 0 2 1 9 13 12 9 9 2
23 11 11 13 10 10 9 15 13 1 9 11 11 2 9 11 11 2 11 11 11 2 11 2
24 11 3 13 1 9 11 11 2 11 2 11 2 2 11 2 11 11 7 11 1 13 1 11 2
5 16 9 15 13 2
22 9 2 9 10 1 9 9 11 13 9 2 9 2 11 2 11 2 11 2 7 11 2
9 3 1 11 13 9 15 13 11 2
17 10 9 13 10 11 7 11 1 13 9 9 7 13 1 9 9 2
24 13 11 11 11 2 10 9 9 15 13 2 7 9 11 2 1 9 12 3 13 13 9 10 2
37 9 9 15 13 9 3 3 13 1 9 12 2 12 1 12 2 12 2 1 13 12 9 9 0 3 11 11 7 11 11 15 3 13 1 9 9 2
26 9 0 13 1 9 9 9 11 11 1 11 11 2 11 2 7 11 2 7 9 0 13 1 9 9 2
23 11 11 2 11 2 11 11 11 2 13 9 15 13 1 11 11 2 11 2 13 11 11 2
16 15 13 1 10 9 1 9 7 9 0 7 3 13 1 13 2
7 11 13 9 9 15 0 2
66 9 9 13 1 10 9 0 2 1 11 16 11 13 12 2 12 11 2 7 11 13 12 2 12 11 2 9 9 1 9 13 1 13 9 13 9 12 1 5 1 12 11 2 11 11 7 9 1 11 0 10 3 13 7 13 1 0 13 1 13 9 9 9 7 9 2
48 15 13 9 9 11 11 7 3 3 13 3 9 11 11 7 1 9 3 13 9 15 13 1 9 9 10 9 1 13 9 9 9 9 13 14 13 1 0 9 13 1 2 9 9 2 11 11 2
15 9 10 13 1 9 9 0 9 9 11 11 2 11 11 2
19 12 1 9 11 13 1 11 2 7 9 9 11 15 13 9 10 3 13 2
16 16 9 13 9 13 9 2 13 9 9 10 13 1 9 10 2
14 16 9 10 13 2 2 1 9 11 3 13 9 10 2
35 11 10 13 1 9 9 1 9 11 13 9 11 11 9 12 2 12 11 2 3 13 11 11 11 2 11 11 11 11 2 7 10 9 11 2
20 3 9 13 9 13 1 9 2 9 9 13 9 2 7 9 9 13 9 9 2
34 11 3 13 11 13 1 1 13 11 11 2 11 13 1 11 2 11 13 2 13 1 9 9 9 9 9 1 9 15 13 1 9 0 2
31 9 9 9 2 13 9 0 1 9 11 0 2 2 1 9 10 11 2 10 9 2 9 11 2 13 1 9 1 9 11 2
29 11 9 9 2 9 9 7 9 9 0 2 13 9 9 7 9 9 13 10 9 9 15 3 13 1 9 9 0 2
15 1 10 2 9 11 3 13 1 11 1 9 15 3 0 2
60 16 12 7 3 9 15 13 1 9 9 1 9 9 9 9 9 2 9 15 13 3 13 1 9 9 2 7 2 7 15 3 13 12 0 0 2 13 9 2 16 9 13 1 13 9 0 15 13 9 16 9 2 15 13 3 13 1 9 12 2
31 11 2 12 2 11 11 13 9 9 11 11 15 13 1 11 11 11 2 1 9 1 9 9 9 11 1 9 0 11 11 2
18 16 14 13 9 0 1 9 9 1 9 2 15 3 13 1 9 0 2
22 9 11 5 11 11 13 13 11 11 1 9 11 11 7 13 13 9 9 12 7 12 2
25 16 13 9 1 11 2 9 11 11 13 9 9 11 1 13 1 11 1 13 7 12 9 9 13 2
13 11 13 9 15 13 1 9 11 1 11 2 11 2
12 9 3 13 7 9 3 2 9 13 1 9 2
15 9 15 3 13 3 1 9 11 2 11 2 11 7 11 2
21 16 13 9 11 7 11 15 10 3 13 2 11 11 2 13 1 13 9 11 11 2
9 11 2 11 11 3 14 13 11 2
33 16 14 13 1 9 1 11 2 9 11 11 2 11 11 11 13 2 16 14 3 3 2 1 1 11 7 9 2 9 1 9 0 2
27 11 11 13 9 11 11 2 10 9 11 2 15 13 1 11 11 2 11 11 11 1 11 2 11 11 2 2
25 14 13 9 0 15 13 2 3 11 11 1 10 9 15 13 9 1 13 9 2 9 11 1 9 2
39 3 13 10 9 1 9 9 9 16 13 11 11 11 11 2 10 9 1 11 11 11 15 13 1 9 11 7 11 13 9 12 7 12 15 14 13 1 9 2
21 1 11 13 1 12 9 2 11 13 1 9 2 2 13 1 9 15 3 13 9 2
36 9 13 1 9 1 11 11 2 11 11 1 11 11 11 7 9 9 9 1 9 11 2 11 11 2 1 11 11 11 7 9 1 11 11 11 2
2 11 2
18 10 9 13 1 12 9 16 9 2 9 2 9 2 9 2 7 9 2
14 14 2 0 15 1 9 2 2 3 15 13 1 9 2
33 3 9 0 11 11 2 11 11 13 13 9 1 13 9 0 12 2 12 13 3 1 11 11 15 13 13 1 9 1 12 2 12 2
14 11 13 9 1 11 11 2 11 2 11 11 2 11 2
24 9 0 13 9 9 0 15 13 1 12 2 12 7 12 2 12 2 9 2 9 9 9 0 2
59 13 15 13 1 9 9 11 1 9 13 9 0 9 13 1 11 15 13 10 9 9 15 0 1 9 9 1 9 2 13 3 15 13 9 9 11 7 9 3 13 16 9 9 13 1 9 16 1 9 0 2 9 13 9 1 13 9 9 2
19 9 15 0 10 3 13 9 13 13 2 13 1 0 2 0 1 11 11 2
45 11 11 15 13 1 9 9 12 2 12 3 13 9 2 13 9 9 11 1 9 7 3 13 9 15 0 1 9 11 11 2 11 11 2 15 1 9 13 3 0 1 10 9 9 2
32 13 12 3 13 1 9 9 9 9 15 3 13 1 11 1 9 1 15 15 13 1 9 11 1 11 11 15 13 1 9 0 2
26 11 11 11 12 13 9 0 1 11 11 11 2 11 11 13 1 11 11 1 12 11 1 12 11 12 2
17 1 11 2 1 9 10 11 13 13 1 9 7 13 13 9 0 2
33 1 10 9 2 9 13 1 10 9 9 15 0 2 7 13 2 13 1 0 9 0 2 3 15 13 9 2 13 0 0 9 2 2
14 1 9 12 11 12 13 9 11 11 11 11 7 11 2
21 11 9 13 10 10 9 15 13 1 11 11 2 11 11 2 11 11 11 2 11 2
40 3 3 1 9 12 2 11 11 13 2 1 12 9 2 13 9 9 9 10 10 11 11 1 11 15 13 12 9 10 16 3 3 13 12 10 9 1 9 11 2
17 11 11 7 11 11 13 9 0 1 9 7 9 1 3 2 3 2
6 3 15 15 13 11 2
6 11 3 13 1 11 2
91 11 11 9 13 10 9 9 0 15 3 13 1 9 11 7 11 11 1 11 11 2 16 10 9 0 15 13 1 9 9 11 2 11 11 11 11 10 13 9 9 1 12 9 10 3 13 1 9 12 1 12 11 7 13 1 9 0 3 12 11 2 1 0 9 13 1 9 12 11 15 3 13 1 9 11 9 2 9 9 9 9 1 9 9 0 15 13 1 11 11 2
22 1 9 3 13 9 2 9 1 9 11 1 2 10 9 0 2 15 13 2 9 13 2
25 13 2 11 13 9 1 9 11 1 11 15 3 13 1 9 11 11 1 9 12 11 12 1 11 2
19 11 3 3 13 1 9 11 11 11 1 11 11 7 9 9 9 11 11 2
14 11 13 9 1 9 11 2 11 2 11 11 2 11 2
14 11 13 10 9 1 11 11 2 11 11 11 2 11 2
14 15 0 13 10 9 1 11 2 9 11 2 11 11 2
15 11 13 9 1 11 11 2 11 11 2 11 11 2 11 2
10 3 15 10 13 7 13 13 9 10 2
7 0 14 2 2 0 14 2
14 11 11 11 2 12 9 12 9 2 2 9 11 11 2
14 11 13 15 12 15 13 9 1 9 0 11 1 11 2
18 1 9 12 2 12 2 9 0 1 9 9 13 1 11 11 2 11 2
47 11 10 13 10 9 2 1 1 11 11 12 7 11 12 2 9 9 9 9 10 13 1 12 5 12 2 11 7 12 5 12 2 11 2 11 11 11 12 12 9 7 11 12 12 9 9 2
13 11 13 1 11 2 11 11 7 13 1 11 11 2
12 11 13 11 2 15 13 9 1 9 13 11 2
26 11 10 3 13 1 9 10 9 1 13 1 9 0 11 11 11 11 11 11 11 11 11 11 11 11 2
30 9 9 10 3 13 1 9 1 9 2 9 9 15 0 2 9 9 15 0 2 7 9 9 16 9 10 13 9 0 2
14 11 13 9 1 11 11 2 11 2 11 11 2 11 2
18 2 11 11 2 16 7 2 15 15 13 9 1 11 2 11 7 11 2
20 9 9 15 13 1 11 11 1 9 10 13 11 11 11 2 11 11 11 2 2
8 9 15 1 9 9 3 13 2
56 3 2 3 15 13 2 9 0 7 13 9 0 2 16 10 10 9 13 1 13 9 11 2 1 9 15 9 10 2 11 7 10 9 0 13 11 11 13 9 2 7 11 13 10 2 10 12 9 7 13 15 13 13 9 13 2
18 1 9 13 1 9 9 2 9 11 13 0 7 3 13 1 9 9 2
16 1 9 12 2 9 13 12 9 2 7 1 9 12 12 9 2
43 15 13 1 9 12 11 12 1 9 12 1 12 13 9 1 11 11 2 11 11 11 2 11 2 11 11 11 9 11 11 11 11 7 11 11 2 11 11 11 2 11 2 2
25 12 2 12 9 10 3 13 9 1 11 7 1 9 12 2 3 12 5 9 11 3 13 9 11 2
8 11 13 9 0 1 9 10 2
22 11 13 9 12 9 15 13 1 9 11 2 9 11 11 2 11 11 11 11 2 11 2
31 1 9 2 9 0 13 9 15 2 10 10 9 13 13 11 11 2 13 15 1 13 9 7 9 0 1 9 0 11 10 2
39 11 13 9 10 9 2 9 2 9 2 7 9 0 15 13 9 9 7 9 15 13 10 9 15 13 0 2 1 9 9 2 9 2 9 9 2 7 9 2
37 11 11 13 1 12 9 12 1 11 11 11 1 11 11 2 13 1 11 1 12 9 2 7 3 13 1 9 0 9 2 11 2 1 9 12 11 2
21 16 16 10 10 1 9 9 13 13 3 2 15 3 13 9 15 13 7 15 0 2
28 1 10 9 2 15 3 13 9 2 9 0 15 3 13 1 9 2 15 13 9 0 1 13 9 9 9 9 2
13 11 13 9 9 11 2 11 2 11 11 2 11 2
13 1 12 9 4 2 3 13 9 15 3 12 9 2
15 11 13 10 9 1 11 11 2 11 11 11 11 2 11 2
10 7 3 11 13 1 9 1 10 9 2
11 3 11 3 13 9 7 11 1 9 9 2
7 9 9 9 10 13 12 2
17 1 9 9 10 2 11 11 13 9 1 13 7 9 13 1 0 2
21 11 11 13 9 9 9 11 11 15 0 1 9 1 12 9 2 12 1 11 11 2
9 9 15 11 13 2 11 7 11 2
10 11 1 13 9 9 1 9 9 9 2
8 11 13 9 9 12 9 11 2
34 9 0 1 12 9 9 2 9 3 13 9 0 1 9 9 2 9 9 7 9 2 7 13 9 10 9 9 1 10 9 1 10 9 2
26 1 10 9 15 13 2 13 9 2 9 11 9 13 1 11 11 11 2 15 13 3 9 1 9 9 2
16 15 3 13 9 9 2 7 1 9 12 15 13 1 11 11 2
29 1 9 9 9 9 2 10 9 9 9 3 3 13 9 1 10 2 10 9 1 1 9 2 1 13 9 1 9 2
27 11 1 11 2 11 2 11 11 11 2 12 11 12 2 12 11 12 2 13 10 11 11 2 11 2 11 2
16 1 1 9 2 11 11 3 13 1 9 9 0 1 9 10 2
30 11 9 1 9 11 11 15 13 1 11 2 9 9 9 15 13 0 2 0 1 11 11 7 11 2 3 13 1 11 2
35 1 9 11 2 9 11 11 2 11 2 9 2 3 3 12 9 1 9 2 9 0 2 11 11 2 11 2 11 2 11 11 2 11 2 2
28 9 10 2 11 7 11 13 9 1 9 15 13 1 12 9 9 9 9 11 2 7 15 13 0 9 15 13 2
25 11 13 9 9 15 3 0 13 1 9 2 9 9 14 3 0 2 14 0 7 14 13 1 9 2
16 11 11 9 11 11 13 11 11 11 11 11 11 11 15 12 2
14 1 9 9 10 2 11 7 11 13 1 13 9 10 2
34 16 10 2 11 13 9 7 13 1 11 2 15 14 13 9 1 13 9 7 13 10 3 9 1 9 10 2 16 9 3 13 15 2 2
33 16 2 9 12 2 9 11 13 9 9 2 9 9 2 0 13 9 2 9 0 2 0 2 1 9 9 2 9 9 10 2 10 2
9 11 13 7 13 9 0 1 0 2
3 9 10 2
10 14 2 11 14 3 13 1 11 14 2
57 1 9 1 9 9 2 9 13 11 11 2 15 13 1 11 2 11 2 13 1 9 7 13 9 2 9 1 9 2 2 11 9 11 2 15 13 15 3 0 7 3 0 1 9 9 11 2 11 15 13 15 0 1 1 10 9 2
11 9 9 10 13 1 13 1 9 7 9 2
6 9 14 13 1 0 2
20 11 10 14 3 13 1 9 16 9 9 1 9 12 3 13 1 11 11 11 2
18 11 10 13 9 15 0 1 9 11 11 2 1 9 9 9 11 11 2
3 11 12 2
16 1 9 13 9 2 11 13 9 1 9 13 1 13 9 9 2
10 9 10 3 3 13 9 1 10 9 2
14 9 9 13 10 9 9 9 10 13 1 9 9 9 2
36 11 2 9 0 11 3 13 11 11 7 9 2 9 1 11 11 15 13 1 11 11 11 2 11 11 2 7 9 9 1 11 11 1 1 9 2
7 10 9 9 10 3 13 2
23 2 11 11 1 11 2 13 9 9 9 11 15 0 7 3 13 1 11 3 1 9 9 2
22 11 3 13 9 1 11 12 9 1 12 9 1 12 9 0 1 3 13 1 11 11 2
44 1 1 9 9 2 9 9 1 11 10 3 13 9 11 2 11 9 0 1 9 11 10 2 3 13 1 0 13 12 9 15 3 13 9 9 16 9 3 13 1 9 11 10 2
17 11 11 11 11 13 0 9 9 9 0 13 0 7 0 1 13 2
16 14 13 9 15 13 9 1 13 1 9 2 1 9 9 9 2
7 3 15 10 3 13 9 2
15 16 9 10 11 11 3 13 3 1 9 9 9 9 11 2
30 11 3 13 1 11 11 11 11 11 15 13 1 11 2 11 2 7 13 9 13 9 0 15 13 1 9 12 11 12 2
23 15 13 10 9 15 13 1 11 2 11 11 2 7 13 9 0 15 7 13 1 9 0 2
24 11 11 2 13 9 2 1 0 9 9 15 3 0 13 11 2 16 9 15 3 0 14 13 2
13 11 11 11 2 2 13 10 9 7 9 9 11 2
14 11 11 13 1 9 12 9 9 1 11 7 13 12 2
34 3 3 13 9 10 10 9 3 13 9 1 10 2 10 9 1 3 13 11 11 11 11 2 12 9 2 3 13 9 9 9 1 9 2
30 11 15 0 1 9 11 7 13 1 9 0 10 2 13 9 1 9 9 3 13 9 9 13 7 13 9 7 9 9 2
15 3 3 9 7 9 13 2 16 9 14 13 9 7 9 2
21 9 1 9 13 9 1 13 11 2 11 9 2 11 1 11 12 1 9 11 12 2
30 15 3 13 9 0 10 9 2 1 10 9 10 10 9 0 12 2 12 1 10 9 13 2 13 1 9 2 9 9 2
19 11 11 0 7 13 0 2 13 1 9 2 9 9 7 13 2 3 9 2
7 11 3 13 1 9 0 2
19 9 12 2 13 9 9 1 9 0 15 13 9 11 11 7 9 2 9 2
24 11 11 11 2 15 3 13 1 11 2 13 9 9 9 1 11 15 13 1 10 9 1 11 2
19 16 11 11 3 13 9 15 0 2 16 13 9 9 11 11 1 9 9 2
39 1 12 3 2 11 3 13 10 9 13 11 11 11 15 13 10 9 1 9 11 2 3 11 1 9 1 11 11 11 11 2 15 13 1 9 9 15 0 2
7 11 11 13 1 9 9 2
19 9 9 1 9 10 13 10 9 7 9 0 2 3 1 9 11 7 11 2
29 11 11 11 11 13 10 10 11 11 15 13 1 11 2 15 13 1 11 2 11 2 11 11 12 11 2 11 11 2
25 9 2 9 11 15 13 13 9 1 9 9 15 1 9 15 3 0 1 3 3 13 9 15 0 2
20 11 10 9 2 9 13 1 10 9 9 1 10 9 0 0 2 2 11 2 2
7 16 9 3 3 14 0 2
21 0 13 1 9 0 1 9 9 7 9 9 1 9 9 11 11 11 11 11 11 2
9 11 9 10 13 1 11 2 11 2
44 11 9 13 10 10 9 9 2 9 9 2 1 9 9 9 11 2 15 13 9 5 11 5 7 5 11 5 2 16 13 13 9 11 2 16 9 10 13 2 11 2 7 11 2
26 1 12 11 12 2 12 9 1 13 2 11 13 1 9 9 7 13 9 1 11 11 11 2 11 11 2
15 16 10 2 10 9 3 13 1 11 11 11 1 9 9 2
51 1 9 16 11 3 13 9 9 0 9 2 11 13 0 1 2 11 11 11 2 7 13 12 9 0 2 2 11 2 7 2 11 2 2 15 9 13 9 9 9 1 9 12 9 2 2 11 11 11 2 2
21 3 9 12 2 12 2 15 13 1 11 11 1 11 11 3 13 1 9 0 9 2
12 16 7 10 2 15 13 1 9 7 10 9 2
28 15 13 13 9 9 9 2 9 9 9 2 9 7 9 9 12 2 13 1 13 1 11 1 9 15 13 11 2
13 1 9 12 2 15 13 9 9 11 11 11 11 2
11 13 3 9 2 9 9 13 9 13 11 2
14 9 9 10 13 9 9 9 0 11 1 9 15 0 2
11 1 10 9 7 9 11 3 13 9 9 2
22 9 12 2 12 9 12 11 12 2 2 9 12 9 12 9 12 2 2 9 9 13 2
15 11 11 13 2 2 9 15 13 3 3 13 1 15 13 2
13 12 9 1 1 10 9 13 12 0 0 1 9 2
33 1 9 11 9 10 2 9 3 13 1 9 9 7 9 1 13 15 13 3 0 7 0 16 3 15 3 13 9 9 3 1 9 2
18 1 9 12 10 10 11 7 11 11 13 11 11 2 13 9 11 11 2
18 9 12 9 10 2 11 2 13 1 9 1 9 11 1 11 2 11 2
32 11 3 3 13 9 1 10 10 9 15 13 1 11 3 11 11 2 9 10 15 0 13 9 11 11 2 11 11 2 1 11 11
21 15 3 9 13 1 10 10 9 9 9 15 0 15 14 13 1 9 9 11 12 2
24 11 7 11 7 11 2 13 9 7 9 15 13 11 1 9 9 2 9 3 13 9 0 9 2
21 1 9 2 13 3 9 2 1 1 9 2 15 13 9 9 0 7 9 9 0 2
19 11 13 10 10 9 15 13 1 11 11 2 11 11 2 11 11 11 2 11
7 11 13 3 9 15 0 2
10 14 13 15 13 2 9 0 14 13 2
13 15 13 10 9 11 11 11 2 11 11 11 2 2
37 11 11 1 1 11 11 11 11 3 2 3 13 12 5 2 12 5 11 1 9 9 3 2 3 12 9 5 9 1 9 9 12 2 12 9 11 2
17 11 11 13 9 9 9 2 11 2 9 2 1 11 11 1 11 2
31 1 9 9 11 11 2 9 11 11 14 3 13 1 9 11 2 7 11 2 16 3 13 1 9 11 11 15 13 9 11 2
11 1 9 10 0 2 3 11 13 9 9 2
28 11 13 2 2 3 15 13 0 2 11 11 2 1 9 2 10 9 2 10 9 15 14 3 13 2 10 9 2
21 11 2 9 10 3 13 16 9 2 9 11 3 13 1 3 0 7 1 3 13 2
17 11 11 13 9 15 13 1 11 11 2 11 11 2 11 2 11 2
29 11 11 7 9 11 2 1 9 11 2 11 11 2 13 10 9 11 11 15 3 13 1 10 0 9 11 11 11 2
11 11 11 13 9 9 11 1 12 2 12 2
26 13 12 9 0 15 13 1 9 2 9 9 2 9 0 2 9 9 2 2 9 15 13 2 7 9 2
28 11 3 13 11 2 11 2 7 11 1 9 2 9 7 9 2 9 1 10 1 9 2 9 7 9 2 9 2
45 3 1 9 13 11 2 11 2 11 11 11 11 11 2 9 11 2 11 2 11 2 11 11 2 16 13 7 15 13 1 11 2 2 16 13 9 13 9 11 2 11 11 2 11 2
12 9 11 13 9 1 9 9 15 13 1 13 2
11 9 13 9 12 1 12 5 2 13 0 2
24 11 2 9 9 15 3 13 2 1 9 9 2 9 2 9 2 7 9 2 13 9 15 0 2
4 3 2 3 2
76 11 11 11 2 12 11 13 10 9 9 9 9 9 15 13 1 9 0 9 11 11 11 11 2 11 2 7 3 2 3 9 9 2 9 1 10 11 2 11 3 13 1 9 2 12 9 2 16 2 11 13 11 16 15 13 9 13 10 11 2 12 9 13 1 9 9 9 7 3 1 13 9 9 1 9 2
13 9 7 9 15 3 13 3 13 1 13 9 0 2
23 11 10 3 13 13 2 9 2 7 13 9 11 2 11 7 0 2 0 1 9 11 11 2
25 1 9 9 12 2 15 13 9 9 9 11 11 2 7 1 9 11 12 15 13 1 12 9 0 2
6 10 0 9 13 9 2
15 11 10 13 1 11 11 11 7 9 5 12 2 12 9 2
12 11 11 13 9 9 7 9 9 1 11 11 2
16 9 9 9 3 13 1 9 15 2 16 13 3 9 9 9 2
8 9 9 11 13 1 11 11 2
30 1 9 11 2 9 13 10 9 1 13 11 0 2 15 13 9 9 0 7 13 1 9 9 1 13 9 9 0 0 2
8 11 13 13 9 15 13 13 2
64 11 11 13 9 11 2 9 9 2 9 9 9 15 1 9 9 13 1 0 1 9 13 1 9 2 13 9 0 5 11 2 16 9 9 2 9 2 9 13 2 9 9 9 15 3 13 13 0 7 0 0 13 1 9 3 3 13 13 2 13 1 9 2 2
10 11 11 11 11 11 13 9 11 12 2
18 1 9 10 2 9 15 13 1 10 9 9 15 0 13 9 2 9 2
29 11 13 1 9 0 16 13 9 12 9 0 1 11 7 9 2 9 9 10 9 1 9 11 11 11 2 11 2 2
9 0 9 9 11 2 11 7 11 2
30 0 1 11 1 9 1 11 9 9 9 1 11 11 12 11 13 1 9 12 9 9 2 13 1 11 11 1 11 12 2
25 9 13 12 9 2 12 11 12 2 7 9 13 12 2 12 12 16 9 9 13 12 9 5 12 2
23 11 7 11 11 13 9 1 9 11 0 1 9 9 1 11 7 9 11 1 11 1 9 2
9 2 3 15 14 3 13 11 11 2
18 11 11 13 9 9 9 1 9 11 2 11 11 2 11 11 2 11 2
15 9 0 0 7 0 10 13 1 11 11 7 11 9 9 2
39 15 10 3 13 1 9 13 9 11 11 10 2 15 3 15 13 1 13 9 2 9 1 9 10 2 15 13 9 1 9 10 2 1 3 11 7 11 13 2
12 15 13 9 12 11 11 2 12 2 12 2 2
10 11 11 11 3 13 1 12 11 12 2
12 11 5 9 9 3 3 13 9 1 9 9 2
16 15 13 1 11 11 12 1 11 11 2 11 1 12 11 12 2
39 16 9 13 1 9 12 9 1 11 1 9 12 2 15 13 9 15 13 12 9 13 9 9 1 10 9 2 7 15 3 13 1 10 9 9 11 15 0 2
21 11 11 11 15 13 1 9 12 1 11 2 13 13 7 13 1 10 9 9 0 2
40 9 15 13 12 7 3 2 9 7 9 9 7 9 15 13 9 15 0 7 0 0 2 15 13 1 9 9 2 9 2 7 9 9 7 9 9 9 15 13 2
17 9 1 9 11 13 9 11 11 1 13 9 15 13 1 11 11 2
35 1 13 9 11 11 11 2 11 13 9 11 11 2 15 13 11 11 7 11 11 1 11 2 1 9 0 1 15 7 13 15 1 13 9 2
18 9 10 13 9 12 9 2 12 5 2 7 13 9 9 1 12 9 2
11 7 0 0 9 11 16 11 9 9 0 2
24 11 11 2 1 9 9 9 11 2 13 10 9 15 13 3 0 1 9 9 9 9 1 11 2
45 11 11 11 13 11 11 12 2 12 2 13 1 12 11 12 1 11 11 2 11 11 2 11 2 13 1 9 12 2 12 9 9 11 2 11 11 13 11 11 1 9 12 2 12 2
60 11 9 9 0 1 9 9 13 11 11 11 11 11 2 11 2 15 13 9 12 1 11 11 11 2 11 2 7 13 1 9 2 9 1 10 9 1 11 11 2 11 9 10 2 11 15 0 13 11 11 11 11 2 11 2 12 1 11 11 2
11 3 13 12 9 1 9 2 9 9 0 2
24 7 15 13 16 9 15 13 9 7 2 15 13 2 9 10 2 15 13 9 9 11 15 13 2
33 9 10 3 13 9 9 0 9 2 9 0 1 11 2 1 9 9 2 9 0 1 9 11 1 1 9 14 13 9 2 7 9 2
19 16 2 12 9 9 15 13 1 9 9 9 15 3 13 1 12 9 9 2
17 16 9 0 9 13 2 10 9 2 9 2 1 9 14 3 13 2
17 9 0 13 1 11 11 2 11 10 13 16 9 9 2 9 0 2
10 15 13 1 9 2 9 9 15 0 2
17 1 10 9 3 3 13 10 11 2 10 1 13 1 9 11 15 2
32 1 12 1 12 11 12 2 11 7 11 13 10 9 9 2 9 15 0 1 9 7 9 2 9 9 1 11 11 2 11 11 2
7 11 11 13 9 9 9 2
46 9 9 9 15 13 13 1 9 11 0 3 13 9 9 9 9 9 2 9 2 9 9 9 2 2 9 2 15 13 9 9 9 9 1 9 15 0 2 3 3 13 7 13 1 9 2
19 11 11 3 14 0 13 7 3 1 9 9 11 11 11 9 10 3 13 2
13 9 13 9 2 16 1 9 9 13 9 3 2 2
16 11 13 10 9 1 11 11 2 11 11 2 11 11 2 11 2
16 9 13 2 7 15 3 13 10 9 1 9 2 11 11 11 2
8 3 10 9 14 13 9 10 2
2 13 2
22 1 9 12 2 10 2 9 9 11 3 3 13 1 10 9 11 1 9 2 1 11 2
59 1 13 2 1 9 0 9 9 13 13 9 16 2 9 7 9 1 9 2 9 9 7 9 9 0 2 9 9 9 0 13 2 9 2 9 2 9 7 9 13 9 2 9 2 9 7 9 2 9 5 9 2 9 9 2 9 7 9 2
50 9 15 13 1 9 9 9 2 9 9 9 2 9 10 13 12 9 11 1 11 11 11 12 1 11 2 13 2 11 11 2 2 2 11 11 2 2 7 2 11 11 2 2 1 1 11 2 11 2 2
28 10 13 9 1 9 15 13 1 13 1 9 9 2 2 11 13 16 15 13 13 9 7 9 0 9 2 9 2
24 1 9 12 9 9 1 9 12 11 12 2 11 11 7 11 11 13 1 11 1 9 1 11 2
13 7 13 11 13 9 1 9 11 11 1 13 9 2
32 1 9 2 9 9 9 13 9 1 9 0 11 2 1 9 10 2 12 9 10 13 9 0 0 1 9 0 1 13 10 9 2
21 11 10 13 1 9 11 11 11 2 7 13 12 1 12 9 15 13 1 11 11 2
25 13 13 16 3 1 0 2 15 13 11 1 13 1 11 11 7 14 3 13 1 3 13 1 11 2
24 16 9 9 10 9 3 13 12 9 1 9 0 1 10 9 2 16 9 10 13 1 9 0 2
29 1 12 2 12 2 12 2 7 12 2 11 13 11 11 16 13 1 12 9 0 1 11 7 9 12 1 11 11 2
11 9 12 2 12 13 9 0 1 9 10 2
22 11 12 9 0 1 11 13 9 12 1 9 9 11 15 13 0 1 9 9 1 11 2
21 9 11 11 13 1 13 9 15 13 16 11 13 9 0 2 15 13 1 9 11 2
28 11 11 13 12 9 9 2 13 1 0 1 9 13 2 1 10 2 11 11 13 2 9 9 2 1 10 2 2
23 11 9 2 11 2 11 2 2 11 11 11 2 11 2 13 2 12 11 12 12 2 11 2
7 11 9 10 13 1 11 2
10 11 9 13 1 9 9 7 9 9 2
10 11 11 3 13 9 9 9 9 9 2
10 2 3 9 15 3 13 14 3 13 2
14 11 10 13 9 11 7 11 15 13 1 11 11 11 2
20 16 2 1 11 3 9 13 1 9 11 15 13 9 2 3 9 11 9 12 2
27 15 3 13 9 2 9 1 9 9 7 13 1 9 0 2 9 10 3 13 1 9 2 9 1 9 9 2
13 1 12 1 11 15 13 11 11 1 9 9 11 2
31 1 9 15 0 2 9 9 13 1 9 7 9 9 2 9 2 9 9 9 9 2 9 9 2 9 2 7 0 2 0 2
21 11 13 9 9 1 11 7 3 9 11 2 11 2 11 1 11 11 11 11 11 2
25 11 11 13 9 9 9 15 13 1 11 11 7 13 1 0 1 11 1 9 9 9 11 11 11 2
26 9 9 2 9 2 11 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11
31 9 2 9 10 13 1 0 1 9 14 9 11 2 3 9 11 2 11 2 11 2 11 2 11 2 11 2 11 7 11 2
29 2 2 9 12 9 2 9 9 9 2 13 9 0 1 9 11 0 2 2 9 9 11 1 11 11 2 11 11 2
15 1 13 3 9 9 9 2 9 13 1 9 2 9 11 2
32 12 9 1 10 9 11 10 3 11 11 2 11 2 11 7 11 13 11 1 12 7 12 9 11 11 11 15 13 13 9 11 2
50 1 9 15 0 2 13 1 12 11 12 2 13 9 12 9 1 11 2 15 13 1 12 9 11 2 3 2 11 2 11 7 11 2 11 16 1 12 9 11 2 3 2 11 2 11 7 11 2 11 2
16 9 13 15 13 9 0 0 2 3 9 0 2 9 0 2 2
16 11 11 2 2 2 2 13 9 0 15 13 1 11 9 9 2
27 1 9 9 9 3 13 9 0 1 9 1 13 1 9 0 2 13 9 9 2 11 7 9 2 1 13 2
21 11 13 10 10 9 15 13 1 11 11 2 11 11 11 2 11 11 11 2 11 2
8 2 16 3 15 3 13 13 2
19 16 7 10 9 9 15 13 2 7 9 9 9 1 9 10 14 3 13 2
18 1 9 12 9 2 9 9 11 2 11 13 1 13 9 9 1 9 2
40 9 9 10 13 2 11 13 11 11 2 9 9 2 2 1 9 11 2 11 13 11 2 11 2 11 2 11 2 9 2 9 2 0 5 0 2 3 0 2 2
20 10 9 11 2 11 11 2 9 9 7 9 9 15 1 13 13 9 7 9 2
12 11 11 13 9 0 1 11 1 9 11 11 2
16 16 3 13 12 9 2 11 13 1 9 9 1 13 9 0 2
18 14 11 11 13 11 11 11 15 13 9 12 2 15 13 14 10 11 2
40 11 11 10 13 12 9 9 11 2 11 11 11 11 2 15 13 1 2 9 9 9 10 13 1 2 9 10 11 13 9 11 11 7 9 11 11 11 11 11 2
19 11 11 10 13 9 11 1 11 7 3 13 10 9 11 16 15 13 0 2
15 16 12 3 13 7 14 9 15 13 1 9 9 15 0 2
23 9 10 13 9 9 1 9 11 11 11 2 11 11 11 2 7 11 11 11 11 1 11 2
13 10 9 0 2 9 2 13 1 9 9 1 11 2
7 9 10 13 1 9 12 2
11 11 11 10 11 13 10 9 1 9 11 2
16 15 3 13 2 14 1 9 7 9 2 7 14 3 1 9 2
8 3 11 11 3 13 11 11 2
63 14 1 9 11 0 2 15 13 9 2 9 1 13 9 9 9 2 1 11 7 11 1 9 12 2 2 1 0 13 9 9 1 9 2 11 1 11 11 13 1 12 13 12 1 9 10 9 2 11 13 1 9 2 7 0 1 1 9 9 12 2 12 2
20 1 9 9 2 12 9 9 13 13 2 11 11 2 9 9 11 1 0 0 2
27 1 9 11 2 1 9 9 9 13 0 2 1 9 9 9 15 13 7 9 16 9 9 9 13 9 9 2
13 11 3 13 16 14 13 9 0 2 3 9 13 2
25 1 9 13 2 9 0 11 11 11 2 11 2 0 1 11 11 11 2 13 11 11 13 11 11 2
20 9 9 7 9 9 3 13 3 0 2 3 1 9 2 9 0 3 13 9 2
71 1 13 11 11 16 9 11 11 13 9 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 9 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 12 2 7 11 2
26 3 16 10 11 11 13 7 11 11 13 1 13 9 9 11 7 11 1 13 13 11 11 1 9 12 2
9 1 10 13 11 11 1 11 11 2
24 11 2 10 9 9 11 7 11 2 13 9 9 11 11 2 1 1 9 9 9 9 2 11 2
16 11 11 11 11 13 10 9 9 15 13 1 11 11 2 11 2
15 1 9 12 2 11 13 7 10 9 0 16 11 1 11 2
16 16 11 13 1 9 9 11 11 11 2 9 13 1 11 11 2
6 3 2 11 13 11 2
12 11 3 13 1 9 10 9 9 1 9 0 2
21 9 10 13 1 9 12 1 9 2 1 9 11 11 11 3 13 9 9 11 7 11
11 3 9 13 9 1 9 2 9 9 10 2
16 11 2 11 9 15 13 3 13 1 13 7 13 1 9 10 2
32 7 10 2 11 11 7 11 1 11 7 9 2 9 9 9 2 1 11 2 11 2 11 2 11 2 7 11 2 3 13 9 2
14 11 13 9 11 11 2 9 0 13 1 13 9 11 2
30 16 14 13 9 1 9 9 2 10 9 3 13 16 9 9 13 9 2 9 2 9 2 9 2 9 1 9 7 9 2
21 11 13 10 10 9 15 13 1 11 11 11 2 11 11 11 2 11 11 2 11 2
32 11 13 1 11 11 2 2 9 11 11 2 2 1 11 11 11 11 2 15 13 10 10 9 9 11 11 11 2 11 11 2 2
13 11 1 0 13 0 2 1 13 12 9 1 3 2
42 9 0 0 9 13 9 0 15 13 9 9 0 7 11 2 9 9 9 2 1 9 9 13 9 0 15 13 9 2 9 7 9 9 11 11 15 13 9 1 10 9 2
9 1 9 15 13 11 11 1 12 2
20 1 9 12 2 12 9 9 12 11 12 2 10 9 13 1 11 2 9 9 2
21 9 10 3 3 1 13 9 2 3 16 3 0 16 9 9 0 13 9 7 9 2
23 3 2 1 9 10 1 12 9 11 13 9 9 9 11 11 15 13 1 11 2 11 11 2
18 9 13 1 9 2 11 11 2 15 3 13 1 9 9 1 11 11 2
36 16 11 14 3 3 13 9 9 0 2 15 3 3 13 9 1 11 11 11 2 11 13 1 9 16 2 14 13 15 13 1 9 9 9 2 2
25 11 0 0 12 2 8 13 12 12 1 13 12 7 12 9 1 9 7 13 1 12 12 9 9 2
17 10 9 9 0 3 13 1 9 1 9 2 9 7 9 15 13 2
44 9 10 13 9 9 0 15 13 13 9 1 11 1 12 9 3 2 3 2 9 15 9 13 1 11 11 11 7 13 1 11 11 2 1 9 9 12 1 9 12 7 3 13 2
38 9 10 13 9 11 11 7 11 2 9 1 1 9 11 11 13 9 13 9 9 2 9 9 2 9 9 7 9 2 7 9 9 1 9 9 9 9 2
8 9 9 1 9 9 9 11 2
17 14 3 13 16 13 9 10 3 13 9 9 9 9 9 11 10 2
12 1 9 12 11 11 3 13 1 1 9 9 2
40 11 2 0 1 11 2 13 10 10 9 1 1 9 9 11 7 11 11 2 9 11 11 2 15 3 13 9 9 9 9 15 13 1 1 11 11 7 11 11 2
14 11 7 11 2 13 9 9 11 1 9 9 11 11 2
18 9 9 10 2 1 13 10 11 1 10 9 2 3 2 3 13 0 2
17 1 9 9 12 2 11 11 3 0 1 9 12 1 9 11 11 2
15 0 13 14 13 2 16 13 2 15 9 3 13 13 10 2
9 11 13 1 11 11 11 1 12 2
6 9 3 0 13 3 2
29 11 13 9 1 9 0 1 11 2 9 1 1 11 11 11 11 1 9 12 3 13 13 13 7 13 9 7 9 2
20 11 11 2 11 2 12 11 12 2 12 11 12 2 13 10 9 7 9 11 2
18 9 0 11 11 13 9 2 9 0 2 11 7 9 11 1 9 0 2
28 9 10 13 1 9 12 9 9 1 9 2 11 11 13 9 0 11 2 13 1 9 11 2 13 2 9 2 2
16 1 9 12 2 9 9 11 11 11 13 9 10 2 9 13 2
29 1 9 12 15 13 11 7 13 11 2 11 2 11 7 11 2 16 3 1 9 10 11 13 1 11 11 7 13 2
18 16 11 11 13 1 12 5 12 9 2 3 1 11 15 13 9 0 2
22 11 11 11 13 10 10 9 15 13 1 11 11 2 11 11 11 2 11 11 2 11 2
13 15 13 11 11 11 11 1 9 12 1 9 12 2
8 15 13 15 0 13 10 9 2
15 11 9 13 1 9 15 13 9 9 2 9 7 9 15 2
28 9 10 3 13 9 0 15 1 13 9 9 16 3 13 2 7 15 3 3 13 12 9 3 1 9 15 0 2
6 16 2 9 10 13 2
25 11 3 13 2 2 16 9 15 13 1 11 2 3 15 13 16 9 15 0 15 13 11 3 13 2
26 9 9 9 15 13 7 9 15 14 13 7 9 9 1 1 9 10 13 9 9 11 11 1 12 9 2
16 11 14 13 9 9 1 13 9 9 2 16 13 9 9 0 2
19 11 10 3 13 10 9 3 1 9 11 2 7 3 13 9 2 9 0 2
11 11 1 9 12 2 13 9 0 12 9 2
19 9 9 0 7 3 0 1 9 2 9 2 9 2 9 9 7 9 9 2
21 12 2 11 11 11 11 2 11 11 2 2 13 9 9 0 1 9 9 15 0 2
12 1 10 11 2 1 11 3 13 1 9 9 2
13 9 3 13 9 10 7 13 9 9 1 9 9 2
28 3 14 3 13 10 2 11 11 2 11 2 9 9 11 11 11 2 11 2 10 13 11 2 13 2 1 9 2
49 11 15 3 9 11 11 11 9 9 10 1 10 1 12 9 0 2 3 3 13 9 9 2 9 7 9 9 1 11 2 7 9 10 15 13 1 13 1 9 9 1 13 1 1 10 9 9 0 2
36 1 12 11 12 9 9 1 9 12 2 12 1 9 11 2 16 11 11 11 11 13 9 9 12 2 12 1 9 11 2 13 9 11 7 9 2
17 16 11 11 13 9 2 9 13 9 9 7 13 9 9 9 9 2
5 0 16 15 13 2
18 11 7 12 9 13 1 11 2 7 9 0 11 13 13 15 9 3 2
14 9 10 13 9 0 7 0 1 9 9 7 9 9 2
150 11 9 15 3 13 1 11 13 9 9 9 9 11 11 11 15 13 12 5 1 9 11 2 9 9 9 9 11 11 15 13 12 5 1 9 13 1 9 11 2 9 9 9 0 15 13 12 5 1 9 15 13 1 9 11 11 2 11 11 11 11 11 11 11 12 2 8 2 9 1 9 11 1 11 1 9 11 11 9 2 11 11 11 11 11 11 11 11 11 11 13 9 11 11 11 9 2 9 11 11 2 11 11 11 2 11 12 2 8 2 11 11 2 9 2 9 11 1 9 11 9 2 11 11 11 11 11 11 11 2 11 11 12 2 8 2 11 11 2 2 9 1 0 2 1 11 1 9 11 11
21 11 11 11 2 3 13 1 11 2 2 13 0 1 11 11 1 9 12 2 12 2
10 11 13 1 9 11 1 11 1 11 2
23 7 7 9 13 1 14 13 1 9 1 9 12 2 7 3 13 9 11 1 9 9 9 2
25 16 3 2 13 3 15 13 16 9 10 13 9 9 0 9 11 2 9 1 11 2 11 11 13 2
55 11 2 9 0 13 1 13 9 9 1 2 9 0 1 9 2 9 2 2 2 13 9 0 2 13 9 1 13 9 2 9 9 1 9 1 9 13 9 2 9 2 7 13 1 13 9 1 3 2 3 13 9 9 9 2
17 9 10 11 11 3 13 9 11 2 16 16 13 9 16 13 9 2
22 16 3 13 9 7 10 9 1 1 9 7 9 13 2 3 3 10 9 15 1 9 2
36 11 13 10 9 15 13 1 9 9 2 3 9 10 13 1 13 1 9 15 13 2 13 2 13 2 7 13 2 7 13 9 15 13 1 9 2
7 11 11 3 13 9 11 2
18 3 10 9 13 2 14 9 9 13 9 0 2 2 11 11 12 2 2
11 11 11 3 13 13 11 1 9 9 9 2
5 3 9 9 10 2
16 15 13 3 2 2 3 15 13 9 1 1 11 11 16 13 2
17 9 11 1 11 11 11 11 11 11 11 13 1 9 13 9 11 2
16 9 0 11 13 9 7 9 13 0 11 1 9 9 13 0 2
18 1 10 2 15 3 13 9 1 9 9 9 15 7 9 2 9 13 2
12 3 15 14 9 11 15 9 0 13 1 11 2
20 1 9 9 9 2 9 3 13 3 0 2 13 1 9 9 7 13 15 0 2
19 3 1 9 12 2 10 9 11 13 11 2 11 13 1 11 1 11 11 2
8 15 0 9 0 1 9 0 2
7 11 10 13 1 9 12 2
22 11 9 13 9 0 1 11 2 7 10 9 9 12 13 9 9 1 9 7 9 0 2
9 15 13 1 9 9 1 9 12 2
40 1 9 0 1 11 7 11 11 2 9 1 9 13 9 1 11 11 2 11 7 11 11 7 11 2 13 11 11 2 9 2 2 7 3 13 11 1 9 9 2
39 11 11 13 9 1 9 9 7 9 2 9 9 9 1 11 1 9 12 1 11 7 11 2 10 9 1 9 15 13 1 9 9 11 2 11 2 11 11 2
13 9 2 1 13 2 13 11 3 13 1 9 9 2
46 16 2 11 13 9 2 11 2 7 13 10 9 7 9 15 15 13 1 9 9 11 11 11 11 2 16 3 1 9 11 1 9 2 9 9 11 15 13 9 10 7 0 0 13 15 2
26 16 2 10 9 3 13 1 9 9 1 10 9 1 13 9 9 1 9 9 2 9 7 13 9 9 2
17 3 13 1 9 3 3 9 2 9 2 7 9 15 3 15 13 2
24 9 10 13 9 9 15 13 9 9 0 15 13 9 9 9 15 3 13 1 9 7 9 9 2
32 1 10 9 11 11 13 1 12 9 7 12 9 2 16 13 9 10 1 9 11 11 15 13 1 12 9 2 2 16 2 11 11
17 1 13 3 2 9 9 13 13 2 13 1 9 9 7 9 9 2
27 11 13 13 9 11 2 11 13 12 9 0 2 11 11 7 11 11 2 7 11 11 1 9 12 2 12 2
17 9 10 13 1 9 10 9 1 9 9 9 11 1 13 9 9 2
29 16 9 2 13 9 9 2 7 3 9 10 15 13 2 16 3 15 3 13 9 0 2 3 15 13 1 15 0 2
14 11 13 9 1 9 11 2 11 2 11 11 2 11 2
32 9 2 9 10 2 10 9 9 3 13 9 1 1 9 2 9 9 15 2 9 7 9 2 2 13 16 9 3 13 1 9 2
12 10 9 3 13 9 10 1 7 1 9 9 2
17 9 13 1 12 9 1 9 11 1 9 12 1 11 11 2 11 2
11 11 11 11 11 13 10 9 15 13 11 2
16 9 10 13 1 9 12 1 9 1 10 9 0 1 9 11 2
30 11 2 1 9 11 2 13 9 9 7 9 0 2 1 9 1 1 9 9 10 13 12 9 9 15 13 12 9 11 2
5 11 10 9 9 2
26 10 13 1 9 9 1 1 11 11 7 11 2 2 11 13 9 11 11 2 2 7 9 1 9 10 2
8 9 1 10 9 11 13 11 2
7 9 15 3 13 1 11 2
42 1 12 2 9 11 13 13 12 2 7 11 13 9 11 11 2 1 12 2 10 9 13 9 2 16 13 13 13 10 9 3 1 9 12 2 11 11 11 1 9 10 2
24 1 13 9 2 9 3 13 9 0 2 9 9 2 7 13 9 1 9 0 1 12 9 9 2
15 9 13 3 9 1 9 0 16 13 9 0 1 11 11 2
14 7 12 2 13 12 9 15 3 13 13 1 11 11 2
15 1 13 9 2 11 1 11 7 11 1 9 13 1 13 2
9 9 13 1 9 9 7 9 0 2
20 9 10 13 1 9 11 2 11 2 15 13 1 9 0 14 9 1 10 9 2
19 1 9 2 1 9 12 9 10 13 1 12 5 11 2 9 1 9 0 2
10 9 9 13 11 11 11 1 9 0 2
14 11 10 13 1 9 11 11 2 16 11 13 9 9 2
11 11 13 3 1 11 2 11 2 7 11 2
16 9 2 9 9 13 1 11 11 2 9 2 13 0 9 9 2
52 11 11 15 13 12 2 12 2 9 9 7 13 12 2 12 2 9 2 16 2 11 2 11 2 11 2 7 11 2 13 7 11 15 13 1 11 2 11 2 11 2 11 2 10 13 10 9 1 11 1 11 2
15 11 13 10 9 0 13 1 11 11 2 1 9 9 11 2
12 11 11 13 9 0 11 2 11 2 7 11 2
23 9 10 13 9 9 1 9 11 12 1 9 1 11 7 11 2 1 9 11 11 2 11 2
13 11 11 13 9 1 11 11 2 7 13 11 11 2
37 15 13 10 9 0 15 13 1 9 9 15 0 0 2 9 7 9 0 2 15 3 13 9 0 1 9 0 9 7 9 11 1 13 1 9 10 2
33 1 13 2 11 13 9 9 11 1 11 11 2 1 12 1 9 12 13 12 1 9 12 2 16 3 1 12 9 11 13 10 9 2
18 11 13 9 13 9 9 9 2 9 2 9 7 9 3 9 7 9 2
33 9 10 13 9 2 9 9 1 14 13 10 9 9 9 10 2 3 1 9 16 9 9 9 9 12 2 12 13 3 0 13 9 2
24 16 16 13 1 10 1 9 13 0 15 3 13 11 11 15 9 3 10 9 0 11 11 11 2
10 3 11 13 13 11 1 3 13 9 2
16 9 10 13 1 1 13 9 2 9 7 9 9 1 9 11 2
21 1 9 9 2 9 3 0 13 1 9 2 13 2 13 9 1 9 1 9 0 2
18 9 0 9 11 13 16 9 2 9 9 10 13 1 13 13 1 9 2
26 9 0 15 3 13 13 11 11 3 13 13 11 11 1 13 9 9 2 3 1 13 9 1 11 11 2
16 16 9 15 3 13 16 9 9 13 1 9 9 14 9 13 2
25 1 11 11 11 11 11 2 1 9 12 14 13 9 1 11 15 13 1 12 9 0 1 10 9 2
30 9 15 12 13 11 11 2 15 13 9 15 15 13 9 11 11 2 16 9 13 9 2 9 11 11 2 15 13 11 2
27 11 9 11 11 12 13 9 9 15 13 1 9 12 11 12 1 9 12 2 12 9 1 11 11 2 11 2
22 15 3 13 9 9 7 9 2 9 11 15 13 9 9 9 0 2 11 11 11 2 2
35 9 9 11 11 13 1 9 9 1 9 0 2 11 2 2 9 13 11 2 11 2 7 11 2 9 7 9 11 7 11 2 7 9 11 2
7 11 7 9 13 0 9 2
35 1 12 12 9 15 9 11 11 13 1 9 9 2 13 9 9 2 15 13 1 9 0 15 3 13 1 11 7 9 10 3 13 1 11 2
39 11 11 13 1 1 9 12 7 12 2 11 2 11 2 11 3 13 9 2 0 2 0 1 11 2 11 2 11 2 7 11 2 11 2 11 2 12 2 2
24 1 9 2 11 13 9 15 13 9 11 9 2 11 2 1 9 11 1 9 1 13 9 9 2
28 1 9 10 2 9 11 2 9 13 16 11 2 12 1 0 13 1 11 11 11 2 11 2 1 9 11 12 2
10 11 11 13 9 7 9 9 11 13 2
25 1 11 2 11 11 13 11 11 11 11 2 11 11 2 11 11 11 11 2 7 11 11 11 11 2
8 9 10 13 10 9 9 3 2
19 11 11 13 1 11 11 11 1 13 1 11 11 11 2 11 11 1 11 2
42 9 15 13 1 13 9 9 1 11 11 7 9 9 1 11 11 7 9 11 11 2 14 1 2 15 11 12 13 12 9 1 11 11 2 10 9 9 11 7 9 9 2
31 11 15 13 1 9 2 11 11 11 11 2 10 9 13 9 9 12 2 3 13 1 9 11 12 2 12 1 0 11 12 2
13 9 0 2 1 9 9 11 13 10 10 9 9 2
16 9 9 11 2 11 2 11 2 7 11 1 9 12 9 0 2
18 11 13 9 12 7 1 9 10 15 13 9 11 11 1 9 2 9 2
9 9 10 2 9 3 13 1 9 2
21 1 0 2 9 12 3 1 0 13 1 9 9 0 1 10 9 13 10 10 10 2
13 11 11 13 1 9 1 9 11 1 9 11 11 2
19 10 10 9 11 16 11 11 13 1 13 13 9 13 9 9 1 9 10 2
21 9 0 2 3 13 1 9 0 7 9 0 2 3 3 13 9 9 1 9 3 2
13 9 15 13 1 11 7 11 16 13 9 15 0 2
14 16 9 0 1 11 7 11 13 3 1 9 9 12 2
13 3 9 11 7 11 3 13 1 13 10 9 10 2
29 11 3 13 16 13 13 0 2 7 1 3 13 2 2 16 9 2 9 11 13 1 11 11 1 9 9 9 9 2
50 13 15 2 2 11 2 10 9 15 0 9 7 13 3 11 2 7 15 0 0 1 1 10 9 11 2 3 13 9 9 1 9 10 9 0 2 16 15 13 15 1 9 7 13 9 15 3 13 2 2
16 9 13 11 2 9 9 9 2 11 2 7 9 9 1 11 2
17 11 2 15 3 13 11 2 13 16 15 3 13 9 11 15 0 2
20 10 9 9 0 1 11 13 1 9 12 9 13 9 9 11 13 1 9 0 2
59 9 9 0 7 3 0 1 9 9 15 3 3 0 1 9 9 1 9 9 11 11 1 9 9 10 13 1 2 1 12 12 9 9 13 1 9 2 12 12 9 9 2 12 12 12 9 9 13 9 2 7 12 12 9 1 9 15 0 2
16 11 13 11 2 2 13 0 2 7 13 2 9 15 0 2 2
3 0 9 2
5 9 1 11 11 2
21 11 13 1 2 11 2 11 2 11 2 11 2 11 2 11 2 11 11 2 11 2
22 11 11 12 13 9 1 13 11 1 13 9 11 12 16 13 9 9 9 1 9 12 2
20 15 13 11 11 1 12 2 12 7 3 13 11 11 11 11 1 12 2 12 2
13 11 13 10 9 1 11 11 2 11 11 2 11 2
24 1 9 11 11 13 12 11 11 2 16 11 12 15 13 1 9 7 11 12 15 13 1 11 2
25 11 11 11 2 2 13 9 9 9 9 11 15 13 1 11 11 1 11 11 2 15 13 1 9 2
26 15 13 1 11 11 2 2 9 9 15 15 13 10 7 9 3 15 15 13 1 15 1 9 0 10 2
15 15 3 13 13 9 0 1 9 1 11 2 1 9 12 2
18 11 11 13 9 12 1 13 1 11 11 15 1 9 1 9 13 9 2
23 11 11 3 13 10 9 1 11 11 11 11 2 11 11 7 13 1 9 1 13 9 10 2
8 11 3 13 11 1 9 0 2
27 11 9 9 11 11 13 9 13 12 5 2 11 11 2 1 9 12 9 1 9 3 2 3 12 5 12 2
33 11 3 13 11 7 10 9 1 11 2 16 11 7 11 13 1 13 7 13 9 1 11 2 7 9 1 11 3 13 1 11 11 2
25 1 9 9 15 13 13 12 9 1 12 9 9 1 11 11 7 13 11 13 9 9 11 11 11 2
10 9 9 11 13 9 9 9 2 9 2
54 15 13 2 11 13 1 12 9 0 1 11 2 16 11 5 11 12 2 12 11 2 11 5 11 12 2 12 11 7 13 1 11 5 11 12 2 12 11 2 10 9 9 11 11 3 13 1 9 12 1 1 12 9 2
11 10 0 9 13 7 3 3 13 9 9 2
22 11 11 13 10 9 1 9 15 13 9 9 12 12 2 7 9 12 9 2 12 2 2
20 9 0 11 11 2 2 13 9 0 1 11 11 2 13 9 11 11 7 9 2
26 10 9 13 9 9 15 3 2 3 13 9 16 3 13 9 7 13 9 9 7 13 9 9 1 9 2
70 16 1 9 15 13 13 3 2 16 13 3 3 9 0 0 7 9 15 3 0 15 13 1 9 9 7 9 15 13 2 16 9 0 13 1 12 5 2 1 9 9 3 0 1 15 13 1 11 11 2 16 3 13 1 0 2 3 1 9 13 15 13 9 14 13 1 9 9 9 2
27 11 11 15 13 1 12 9 7 9 11 15 13 1 12 9 3 13 7 3 13 1 3 13 9 14 3 2
25 11 7 11 3 3 0 2 11 13 9 9 2 9 1 9 9 2 16 11 13 9 10 9 0 2
11 11 11 3 13 9 12 11 11 11 11 2
9 10 12 9 13 1 9 9 10 2
39 10 1 9 2 9 10 13 1 12 11 0 2 9 11 2 9 11 2 9 11 2 7 9 11 2 2 16 9 2 9 15 0 14 13 1 9 9 10 2
22 11 7 11 13 9 1 9 11 12 0 1 9 9 2 9 11 11 2 12 5 12 2
19 1 1 9 2 9 0 13 9 9 2 9 0 15 0 1 9 9 0 2
18 13 1 11 2 11 3 13 1 9 11 2 15 13 9 1 11 11 2
15 13 10 9 9 0 0 15 13 1 13 9 2 9 10 2
17 11 11 10 13 16 9 13 9 9 13 9 15 13 1 12 9 2
12 3 15 13 3 15 14 0 1 1 9 10 2
15 11 11 2 9 13 9 1 9 9 9 1 9 15 0 2
75 9 10 3 13 9 1 9 9 9 11 1 12 9 11 2 11 11 11 2 2 11 11 11 11 2 2 11 11 11 11 2 2 11 11 11 7 11 11 11 2 11 2 1 9 12 11 12 15 13 1 2 11 12 11 2 2 12 11 12 2 13 9 11 11 11 1 13 9 13 9 2 11 7 11 2
15 9 10 13 1 12 9 15 1 10 9 13 1 9 9 2
9 11 13 9 1 9 0 9 11 2
30 10 9 1 9 13 1 9 9 11 2 16 9 0 13 1 9 9 7 9 2 9 0 9 3 7 3 9 1 12 2
35 11 12 1 11 11 15 0 3 13 13 1 12 2 1 12 9 7 12 9 1 9 9 2 9 2 9 2 7 9 1 9 9 11 11 2
20 9 10 3 3 13 9 2 9 2 7 9 2 7 3 3 9 9 7 9 2
11 1 9 0 3 10 9 3 13 1 3 2
11 11 10 13 9 9 0 1 12 9 10 2
25 10 9 1 12 13 1 11 11 2 9 10 3 13 9 13 11 2 11 11 11 11 11 11 2 2
20 10 9 11 1 9 13 11 15 3 14 13 9 13 13 1 9 9 9 0 2
26 9 9 11 13 9 9 9 9 9 15 13 9 11 2 11 2 13 12 9 9 2 9 7 9 2 2
28 16 11 3 3 13 9 9 1 11 11 11 7 3 13 1 9 2 9 2 1 9 0 15 7 1 9 0 2
14 15 13 11 11 11 1 12 11 12 1 12 11 12 2
29 11 11 11 2 13 1 11 11 2 2 13 9 11 15 13 1 9 9 11 11 11 9 9 11 9 12 11 11 2
17 9 1 11 13 11 11 2 16 9 1 9 13 11 11 2 11 2
33 11 15 13 1 11 11 11 2 11 11 11 11 2 7 3 9 1 11 2 11 2 11 2 11 2 11 2 11 2 11 7 11 2
20 11 11 13 10 10 9 1 11 11 11 2 11 11 11 2 11 11 2 11 2
10 9 12 11 12 13 9 13 9 9 2
40 3 9 9 9 15 13 13 9 9 7 9 2 7 16 9 1 13 9 13 9 10 13 1 9 9 2 7 3 13 1 9 2 9 1 9 11 9 9 2 2
21 9 11 13 1 9 9 15 13 9 0 1 9 2 11 1 11 13 2 9 2 2
23 11 11 13 10 10 9 15 13 1 11 9 11 11 2 11 11 11 2 11 11 2 11 2
4 9 9 13 2
26 11 2 11 11 7 11 13 1 9 2 7 1 3 15 13 9 9 2 9 11 2 7 9 11 11 2
25 9 11 13 1 9 9 9 1 13 9 7 9 9 7 13 1 9 13 9 1 13 9 3 0 2
20 1 10 1 3 13 9 1 9 9 2 9 9 3 15 3 13 9 1 9 2
20 11 11 13 10 9 9 9 1 11 2 11 11 2 11 10 13 1 9 12 2
13 11 11 13 12 9 2 9 0 2 0 7 0 2
24 11 0 3 13 9 7 13 1 0 2 1 13 9 9 1 1 9 2 1 13 10 9 9 2
16 11 3 0 1 9 9 1 12 9 1 13 9 9 1 9 2
20 1 12 9 11 13 9 9 1 11 2 1 9 15 13 1 9 1 13 9 2
30 11 2 11 13 9 11 11 2 9 16 13 9 11 2 9 16 13 9 9 10 1 9 9 2 9 9 11 2 9 2
28 1 1 9 9 9 9 13 2 11 2 11 11 7 11 2 11 2 11 11 7 11 11 11 2 7 11 2 2
33 1 9 12 11 13 1 12 0 1 9 12 2 16 13 13 1 9 12 1 9 0 7 3 13 13 9 12 1 9 12 11 12 2
132 11 11 11 13 9 11 11 11 1 9 10 13 9 2 16 1 9 2 9 11 11 11 11 5 11 11 2 15 13 2 16 0 9 9 11 11 11 7 11 11 11 13 1 9 3 7 11 11 9 13 13 11 11 15 13 11 11 11 11 13 9 11 11 0 1 9 12 2 12 1 9 9 8 2 12 2 16 13 9 11 11 12 11 13 9 9 7 13 9 1 9 11 2 7 13 11 11 1 11 11 1 9 12 13 1 11 11 10 9 9 11 1 9 7 9 3 13 9 2 9 1 11 11 3 13 9 0 3 13 9 11 2
14 11 11 2 2 13 10 9 2 9 2 7 9 11 2
37 1 9 12 2 13 9 9 1 9 9 2 11 2 11 11 2 10 9 9 9 9 2 13 1 13 9 1 9 9 1 13 9 9 0 15 0 2
11 11 10 13 9 1 9 9 9 2 9 2
9 11 2 1 0 13 1 10 9 2
25 1 1 9 9 15 0 3 13 9 9 2 3 13 9 15 13 13 9 1 9 9 1 9 11 2
15 15 3 13 9 1 9 1 14 13 9 2 13 10 9 2
14 9 0 9 10 3 13 9 2 13 12 9 12 9 2
33 11 15 13 9 7 9 7 9 10 13 10 9 13 7 13 9 9 1 11 11 2 11 11 2 1 9 12 1 11 2 11 2 2
19 11 13 1 11 2 7 14 0 3 2 11 13 9 15 13 11 7 11 2
15 9 9 10 13 11 11 1 13 13 11 11 1 9 12 2
34 9 13 16 9 11 11 11 3 13 1 11 11 11 2 11 2 7 16 9 9 14 3 13 1 9 2 9 9 11 7 1 9 0 2
23 1 9 12 2 15 13 1 11 1 1 15 13 9 9 1 9 0 7 0 1 11 11 2
16 11 13 10 9 1 9 11 11 2 11 11 2 11 11 11 2
16 9 10 13 11 11 11 2 11 11 7 9 0 9 9 11 2
10 11 9 10 13 11 16 15 13 9 2
11 11 13 13 2 13 7 13 16 15 13 2
35 11 11 11 11 13 1 9 11 11 16 9 3 13 1 11 2 11 11 11 13 1 15 7 13 10 9 1 11 2 10 11 11 1 15 2
16 10 9 3 13 1 13 9 15 15 2 7 13 9 0 9 2
35 1 9 15 13 9 7 9 15 13 0 2 15 13 9 15 13 9 15 3 13 10 13 1 11 2 10 9 10 13 1 9 7 9 13 2
19 15 13 9 9 0 9 11 2 3 9 9 15 3 13 1 14 13 3 2
10 11 3 13 11 2 16 11 14 13 2
9 15 13 1 9 15 0 7 0 2
18 9 9 1 12 9 11 2 1 12 5 2 2 13 9 7 13 9 2
39 9 9 0 11 11 11 7 2 11 11 11 11 11 2 1 9 11 2 9 13 1 9 9 0 11 2 13 10 9 9 15 13 1 11 2 9 11 11 2
16 9 9 10 13 1 9 11 11 2 11 0 13 1 11 11 2
30 9 0 11 3 13 1 9 0 2 9 2 9 7 9 2 9 9 2 7 9 7 9 2 2 9 2 7 9 9 2
11 3 11 13 9 1 13 9 10 1 9 2
32 9 2 7 1 3 2 3 13 1 9 9 7 9 9 2 13 9 15 13 9 2 9 9 15 13 1 9 2 9 9 9 2
24 1 10 2 15 3 13 9 11 11 11 11 11 2 11 2 7 13 9 0 1 10 9 9 2
26 15 13 13 9 15 14 3 13 16 3 13 13 9 2 1 0 1 9 9 2 9 9 7 9 9 2
6 9 1 9 9 11 2
26 11 13 9 1 9 0 11 11 2 11 12 3 13 1 9 2 9 11 11 9 2 11 11 11 2 2
29 9 0 11 13 1 9 9 9 2 9 9 2 7 3 9 2 7 3 9 9 15 1 9 9 2 9 9 13 2
27 1 11 11 12 2 11 11 11 11 13 9 9 11 1 9 11 2 11 2 11 2 11 2 11 2 11 2
28 16 9 14 13 9 2 9 9 9 7 13 1 1 10 9 10 2 10 9 9 14 13 7 3 3 13 9 2
30 3 3 15 13 1 9 1 9 2 9 2 9 7 9 0 2 16 3 0 9 7 9 10 0 1 15 13 1 9 2
5 9 15 3 13 2
15 13 3 9 5 9 15 3 13 9 1 13 1 9 0 2
20 13 1 10 9 11 2 15 13 9 7 9 15 0 13 1 9 7 9 11 2
23 1 11 11 12 2 9 0 13 1 9 7 9 2 1 9 13 11 13 1 12 1 11 2
10 11 11 13 1 12 7 13 13 12 2
21 1 9 12 2 11 13 9 0 1 9 9 5 9 1 11 1 9 11 2 12 2
35 1 11 11 11 11 2 11 13 1 2 9 9 2 2 7 13 1 9 12 15 1 9 0 13 9 2 1 9 2 11 1 9 9 2 2
14 11 13 9 1 9 11 2 11 2 11 11 2 11 2
10 11 13 1 12 12 1 1 9 9 2
26 9 0 11 1 3 3 13 11 11 11 2 7 3 3 13 1 11 2 11 15 13 1 11 11 11 2
12 14 2 9 10 2 2 9 15 13 1 9 2
28 9 2 9 2 15 13 9 1 9 11 7 9 2 13 9 9 1 9 9 0 1 11 11 11 7 9 11 2
18 11 13 9 11 11 15 12 1 9 9 11 11 15 13 0 1 9 2
12 11 11 13 9 1 11 11 2 9 9 11 2
14 9 13 9 12 14 2 2 3 0 9 13 9 12 2
23 11 13 9 1 9 0 1 9 9 7 9 9 1 0 13 1 11 2 11 1 9 12 2
26 16 11 0 13 9 1 13 9 10 16 15 14 3 13 9 0 2 16 3 3 13 9 11 1 9 2
19 3 10 9 0 15 3 13 3 3 13 15 12 9 15 13 13 9 9 2
12 9 0 13 2 3 11 11 11 13 1 9 2
25 9 10 13 9 9 11 15 13 1 12 9 2 15 3 13 2 13 1 11 1 9 12 11 12 2
20 11 11 13 9 9 11 11 15 13 3 1 9 9 15 13 9 1 9 0 2
19 1 9 9 15 0 10 9 11 11 14 13 1 9 9 16 13 1 9 2
22 11 11 13 10 10 9 15 13 1 11 11 11 2 11 11 11 2 9 11 2 11 2
8 16 11 13 1 9 1 11 2
35 11 11 11 11 2 2 2 13 3 1 11 11 7 11 11 2 2 13 10 9 9 9 13 9 15 13 1 9 11 3 13 1 9 9 2
11 9 13 0 9 9 9 7 3 14 13 2
27 11 13 9 12 5 1 11 11 9 1 9 3 2 3 1 12 5 12 2 7 12 5 1 1 9 9 2
30 9 9 14 3 13 2 16 10 9 2 13 11 2 11 11 2 2 13 16 9 13 1 9 9 1 9 12 11 11 2
28 11 11 2 1 9 15 0 2 13 1 9 13 1 9 10 13 1 15 13 2 7 13 14 0 1 9 10 2
29 1 11 11 12 2 11 11 11 3 13 9 1 11 3 9 11 13 13 9 15 13 11 11 1 9 0 1 11 2
52 9 14 3 3 0 1 9 2 3 13 11 11 1 9 9 2 16 13 9 15 0 7 13 9 1 10 2 3 1 9 0 2 15 13 9 3 13 1 9 0 2 7 0 10 9 15 14 13 1 9 9 2
33 9 13 12 9 1 13 9 9 12 2 12 12 2 2 9 9 12 2 12 9 5 12 2 2 9 10 13 9 9 0 13 9 2
54 11 13 9 11 1 9 3 13 1 9 11 11 15 3 13 0 9 9 13 0 9 2 16 9 11 11 2 13 9 11 2 11 13 1 9 9 2 9 12 2 12 2 12 2 2 16 1 11 11 13 11 11 11 2
23 1 9 12 7 12 2 1 9 11 11 11 2 2 9 2 11 11 11 11 13 9 11 2
19 16 1 9 12 15 3 0 13 11 11 11 1 9 11 11 11 1 11 2
14 3 13 3 9 9 7 13 9 9 1 13 9 9 2
52 1 11 12 2 13 9 9 11 7 11 1 11 7 11 7 11 11 1 11 2 10 9 1 12 9 10 13 1 11 7 13 1 13 12 9 10 7 13 10 9 15 3 0 1 9 2 9 15 13 13 13 2
13 1 9 2 9 9 9 9 10 13 13 7 13 2
11 11 13 9 0 1 12 11 12 1 11 2
36 11 2 11 2 11 2 9 2 11 11 2 2 13 2 13 2 13 7 13 10 2 9 9 2 12 9 13 11 11 9 2 11 11 11 2 2
14 15 3 13 16 10 9 11 3 13 15 1 9 0 2
19 16 3 12 9 10 14 3 13 15 2 15 2 16 13 1 10 9 0 2
6 9 10 13 9 12 2
11 11 13 9 9 0 1 9 9 11 11 2
14 1 9 12 2 9 9 9 15 13 11 13 12 9 2
35 11 11 3 13 16 9 9 11 2 9 9 2 9 9 9 2 9 2 2 13 9 15 13 0 7 13 1 9 2 7 7 16 9 0 2
3 15 14 2
8 13 1 11 2 13 9 9 2
11 1 9 10 15 13 1 9 11 11 11 2
8 9 15 13 13 0 7 0 2
11 9 10 3 13 1 9 1 9 11 12 2
8 3 9 9 9 11 1 11 2
21 9 12 13 1 9 12 11 12 1 12 9 12 2 1 11 11 11 1 9 9 2
16 11 13 10 9 1 9 11 11 2 11 11 2 11 11 11 2
21 9 9 13 2 2 1 12 12 9 9 14 13 2 16 13 1 9 15 13 2 2
17 11 11 13 9 0 1 9 9 1 11 11 13 9 1 9 9 2
14 1 11 2 9 11 0 1 9 13 9 2 11 2 2
14 11 3 13 1 9 9 1 9 9 7 9 9 0 2
81 15 13 11 11 2 7 13 1 11 11 0 11 11 2 15 2 11 12 2 11 10 11 2 13 11 2 13 1 9 2 9 13 2 13 9 2 9 2 7 13 9 0 11 0 7 13 11 0 7 1 9 2 3 1 9 15 7 0 2 0 1 9 2 9 2 9 2 9 2 9 7 13 9 2 9 2 7 0 2 0 2
18 1 9 9 9 11 12 2 13 9 10 13 9 9 9 1 12 9 2
16 11 11 13 9 9 1 9 11 3 13 9 9 1 9 10 2
12 3 9 10 2 9 9 9 1 9 9 13 2
19 11 9 3 3 3 0 1 9 9 1 1 9 12 2 2 12 2 12 2
14 1 13 9 9 9 11 2 11 3 13 9 13 9 2
10 3 11 15 14 9 11 11 13 11 2
45 11 13 1 10 9 9 13 11 11 11 11 11 13 1 9 0 1 11 11 1 9 11 12 2 1 9 10 11 10 2 11 11 11 2 13 1 11 11 7 2 11 11 2 2 2
27 9 2 9 15 3 0 13 1 9 9 13 2 9 15 3 13 1 9 9 16 2 1 9 0 2 9 9
33 11 11 2 11 5 11 7 11 5 11 16 13 10 13 1 9 9 10 2 11 13 3 1 13 13 11 5 11 1 9 11 11 2
44 11 11 11 13 10 9 9 9 9 11 11 15 13 1 9 2 9 11 2 1 9 12 2 11 11 3 13 10 9 7 9 1 10 9 9 1 13 9 1 9 1 9 0 2
35 16 9 1 9 9 9 9 10 3 0 2 7 0 1 9 2 7 9 15 3 0 1 9 10 13 9 10 9 1 9 0 1 11 11 2
28 1 9 1 11 11 11 2 15 13 1 12 9 1 9 9 11 9 9 2 7 1 9 9 11 11 11 11 2
29 1 9 9 7 9 0 2 9 9 0 13 1 11 7 3 2 3 1 9 11 2 1 1 11 11 11 11 2 2
13 9 10 13 1 11 11 11 7 11 1 11 11 2
19 3 1 9 12 1 12 2 9 9 0 13 13 9 0 1 13 9 9 2
25 16 9 10 13 1 9 9 9 2 16 3 13 1 9 9 0 7 0 2 7 13 1 9 0 2
42 11 11 13 1 9 2 9 11 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 16 9 12 11 13 1 9 0 11 11 9 0 2
20 15 13 1 9 0 11 11 11 1 11 2 11 2 11 2 11 2 7 11 2
14 14 15 13 2 15 13 9 11 13 13 15 1 9 2
19 15 3 13 1 11 11 2 11 2 11 11 2 7 13 9 9 1 12 2
16 11 13 9 1 9 11 2 11 11 2 11 11 11 2 11 2
6 13 1 9 1 9 2
16 9 9 9 11 11 13 1 5 12 2 12 12 1 9 12 2
36 9 9 10 13 10 9 15 13 1 9 2 9 7 9 16 15 13 9 2 9 9 1 9 7 9 13 9 2 9 9 2 9 9 7 9 2
21 9 9 9 1 9 1 9 3 3 13 1 9 1 1 10 9 0 1 9 11 2
23 11 9 9 1 11 11 2 2 11 11 2 13 9 9 1 2 11 2 2 9 0 9 2
17 11 15 13 1 11 2 3 13 9 11 1 9 9 9 9 10 2
21 11 11 11 2 13 9 15 3 0 3 13 1 11 11 11 2 3 1 11 11 2
19 1 15 13 9 2 13 9 15 15 13 1 11 11 13 11 15 3 13 2
79 11 13 9 7 13 1 13 9 1 13 1 1 9 1 1 11 11 2 11 15 3 13 9 10 3 13 9 1 13 9 15 13 9 11 13 9 1 9 11 14 13 3 13 15 2 16 13 9 10 9 11 3 13 1 13 11 7 3 13 16 11 3 13 0 9 10 2 16 11 7 11 13 1 9 15 10 2 10 2
8 9 15 13 9 11 1 11 2
18 11 11 11 13 0 1 11 11 11 1 9 11 2 11 2 11 11 2
25 11 1 9 11 11 11 11 11 13 1 9 9 1 10 9 11 11 11 11 16 9 13 1 0 2
6 16 9 15 3 13 2
19 11 11 11 13 9 9 9 12 11 2 9 10 13 1 9 12 11 12 2
27 16 15 13 16 2 9 2 9 1 9 15 0 3 13 2 13 7 9 2 9 14 0 2 13 2 13 2
7 11 11 13 9 10 9 2
17 11 13 13 0 3 13 9 1 11 11 2 11 11 7 11 11 2
14 11 13 9 9 2 9 2 1 12 1 9 9 10 2
16 11 13 10 10 9 1 11 11 2 11 2 11 11 2 11 2
19 9 10 3 13 1 11 11 2 15 12 9 13 1 9 12 11 12 2 2
18 11 11 11 11 7 11 11 13 9 9 11 11 1 9 11 11 11 2
24 11 11 2 2 13 9 15 13 1 13 9 1 1 9 2 9 9 2 1 13 3 9 9 2
31 9 3 13 9 9 15 0 7 13 9 15 0 2 9 3 13 1 9 9 9 9 7 3 9 1 9 13 9 3 9 2
40 1 9 15 0 10 13 9 3 9 10 3 0 1 1 9 2 9 15 3 0 7 9 2 15 13 9 9 2 16 1 9 10 14 13 9 7 9 15 3 2
34 2 9 2 12 2 12 2 9 9 9 11 11 11 7 11 13 16 9 11 11 13 1 10 9 15 13 1 9 9 2 9 9 2 2
28 1 13 1 10 9 11 2 11 13 10 9 0 15 13 11 11 2 2 11 11 2 2 1 10 9 11 11 2
22 9 9 9 15 14 13 9 10 2 7 13 9 9 1 1 9 16 13 9 9 9 2
21 1 9 11 11 11 11 11 11 11 1 1 9 12 13 13 9 11 0 7 0 2
12 11 11 13 10 9 9 11 1 9 11 11 2
13 1 9 10 2 9 9 13 1 9 2 9 9 2
50 9 9 2 11 2 11 2 11 11 2 9 2 11 2 11 2 11 11 1 11 9 12 11 2 11 2 11 11 11 2 9 9 9 1 9 9 11 2 9 1 9 0 0 1 9 9 1 11 11 2
11 15 3 13 16 13 10 9 13 3 0 2
21 1 9 9 11 11 3 0 7 0 1 9 9 9 13 9 7 9 9 15 0 2
18 11 9 10 13 11 13 9 9 0 7 3 13 9 1 13 9 9 2
11 1 9 11 2 9 11 13 1 11 11 2
16 11 13 12 9 0 1 13 11 11 12 1 9 12 9 12 2
59 11 10 13 9 9 11 11 11 15 2 1 12 2 13 1 9 9 9 1 11 2 11 2 11 2 7 11 3 13 1 15 13 1 9 11 11 2 11 11 13 9 9 15 13 1 11 11 2 11 11 2 7 13 1 9 9 11 9 2
12 11 11 13 9 9 12 9 1 11 2 11 2
21 9 10 13 3 1 9 9 12 2 12 2 1 9 12 7 1 9 12 2 12 2
14 11 11 13 9 9 11 11 11 1 2 11 11 2 2
16 11 11 3 3 13 9 2 1 3 9 1 9 9 9 9 2
18 11 11 3 3 13 9 15 0 1 9 9 1 11 2 11 7 11 2
13 12 2 1 9 12 11 12 9 0 9 11 13 2
16 1 9 10 9 9 3 13 7 3 13 9 9 15 3 13 2
20 9 2 12 13 9 9 3 3 2 13 10 12 9 9 15 3 0 7 9 2
8 3 15 10 3 3 3 13 2
26 15 15 13 9 7 9 2 9 10 13 1 11 11 2 11 11 7 10 9 9 11 3 1 9 12 2
8 0 16 9 0 1 9 1 2
18 9 11 11 11 13 9 9 15 13 1 11 2 11 11 2 11 11 2
19 16 1 0 13 0 1 9 9 1 9 9 2 11 11 13 1 9 9 2
6 9 3 13 1 9 2
38 15 3 13 9 11 2 3 9 13 9 9 10 2 16 15 14 3 13 2 7 13 1 11 2 3 9 11 7 9 0 1 11 13 1 9 12 9 2
14 11 7 9 9 1 3 13 1 9 1 12 9 1 2
26 1 12 11 12 2 9 11 11 13 9 1 12 9 11 2 12 9 0 7 12 9 2 9 9 9 2
13 11 11 11 2 2 13 10 9 7 9 13 11 2
22 1 9 9 9 9 9 13 1 9 2 11 9 9 9 13 1 13 9 10 1 9 2
7 0 9 9 9 9 2 2
31 9 9 10 13 12 9 16 11 2 9 2 2 11 2 9 2 2 11 2 9 5 9 2 7 11 2 9 5 9 2 2
23 9 3 1 0 13 13 11 15 13 2 7 1 11 11 1 9 11 2 7 0 11 11 2
84 11 2 2 13 9 9 1 9 12 9 7 9 11 2 11 2 15 3 13 1 9 11 1 11 11 2 9 11 2 9 11 2 11 2 7 9 9 2 11 11 3 13 1 9 11 1 11 2 11 2 2 15 13 3 14 1 13 9 0 2 16 9 0 2 11 2 2 7 0 1 11 11 7 9 11 11 2 11 11 1 11 13 11 2
85 11 13 9 16 12 13 1 9 15 13 1 9 9 3 2 3 9 13 9 13 9 1 9 13 9 13 1 9 9 3 9 13 9 13 1 9 9 3 9 13 9 2 16 3 13 13 9 1 9 10 1 9 1 12 1 9 1 9 9 9 1 12 2 11 1 2 9 9 2 13 9 1 9 9 1 9 10 13 9 9 1 9 15 13 2
31 1 12 9 11 2 12 5 13 9 9 1 9 9 2 3 2 13 1 9 0 2 0 1 9 9 0 2 1 9 9 2
53 9 11 2 11 7 11 2 11 3 13 9 13 14 1 12 9 0 2 13 9 16 9 9 11 11 11 1 11 13 1 9 12 2 9 9 11 1 11 2 7 9 9 11 2 13 9 10 2 13 1 9 12 2
13 11 11 13 10 9 9 12 9 9 11 11 12 2
54 9 12 12 9 9 9 13 1 11 1 9 1 13 9 1 9 9 15 3 0 1 11 11 2 11 15 13 9 10 13 3 11 11 11 2 11 11 11 2 11 11 11 2 11 11 11 11 11 2 7 11 11 11 2
66 11 11 1 9 13 1 9 9 9 11 11 1 9 2 9 9 9 11 12 2 12 9 7 12 2 12 5 1 9 11 11 11 2 1 0 13 1 12 9 2 12 9 2 12 9 7 12 9 2 16 13 9 9 9 10 13 9 9 0 7 9 1 9 12 9 2
17 10 9 9 5 9 13 13 9 16 9 13 13 1 12 2 12 2
11 11 13 9 9 15 13 9 1 11 11 2
21 9 2 9 15 13 13 9 2 9 2 9 2 9 2 9 2 9 2 7 9 2
10 11 11 11 13 9 9 9 11 11 2
21 9 12 9 12 9 2 9 12 13 12 9 2 7 9 1 9 12 13 12 9 2
22 9 1 9 15 0 2 7 9 15 13 9 2 7 9 1 9 15 0 1 9 0 2
12 12 2 9 13 1 9 7 9 2 9 0 2
29 1 9 9 2 9 2 9 9 11 13 2 12 5 9 1 11 11 2 12 5 1 11 2 7 12 5 1 11 2
27 9 13 9 9 9 11 2 11 11 2 9 11 11 11 15 13 9 1 9 9 7 9 9 11 11 11 2
3 9 9 2
8 3 15 13 0 7 9 15 2
20 3 15 13 3 9 11 2 14 13 9 11 15 9 10 3 13 1 9 11 2
18 9 9 9 13 13 1 12 9 2 3 2 9 15 0 13 13 9 2
13 9 10 11 11 13 1 11 11 11 11 15 0 2
18 11 5 9 11 13 9 1 9 11 2 11 11 2 11 11 2 11 2
28 11 11 11 11 11 11 11 2 11 2 11 2 7 11 13 9 2 9 13 1 12 2 12 15 13 9 9 2
13 11 11 2 2 13 10 9 9 9 0 13 11 2
44 9 2 9 10 13 2 13 9 9 11 11 11 2 2 7 3 3 13 11 2 11 11 2 2 2 9 9 3 13 1 9 9 9 2 9 9 2 9 9 7 9 2 9 2
4 9 1 11 2
25 1 13 9 1 11 2 11 3 13 9 1 9 9 9 1 10 9 15 13 1 9 9 9 10 2
21 11 3 13 1 9 9 2 1 9 9 9 1 9 13 3 13 1 9 11 11 2
21 11 10 13 1 9 0 3 2 14 15 13 2 3 9 9 3 3 13 1 11 2
23 11 13 9 0 11 1 12 11 12 1 9 11 5 12 7 3 13 1 9 12 12 9 2
16 1 13 9 9 7 9 2 9 10 3 13 1 10 9 9 2
13 9 1 11 11 11 13 9 13 1 9 1 9 2
43 1 9 12 12 9 0 13 9 0 9 11 2 15 13 1 1 12 3 13 9 9 11 11 2 9 0 9 7 9 11 1 9 12 7 9 9 11 11 11 1 9 12 2
18 1 11 11 13 1 9 10 3 13 9 9 15 9 13 9 1 9 2
30 11 13 9 15 13 1 9 9 15 14 0 2 9 13 1 9 12 2 12 9 15 13 1 9 1 13 2 13 9 2
14 11 11 11 13 9 10 9 0 9 1 11 11 11 2
32 12 11 12 2 7 12 11 12 2 13 9 12 2 13 9 1 9 9 11 15 12 1 9 1 11 1 11 11 1 9 11 2
34 11 13 1 9 0 10 3 1 11 11 2 3 15 13 3 1 11 11 1 9 11 11 2 7 13 3 0 1 11 7 1 11 11 2
17 11 3 13 1 11 2 9 9 11 15 0 2 1 13 11 11 2
44 3 15 13 13 9 15 7 3 3 13 10 1 10 15 15 13 2 13 1 9 11 2 11 2 7 11 2 11 11 2 2 15 1 10 3 3 13 9 1 9 11 7 11 2
9 3 15 3 13 10 9 10 10 2
16 11 13 10 9 1 9 11 11 2 11 11 2 11 11 11 2
23 11 11 13 9 10 9 11 9 15 13 1 9 9 12 2 12 2 15 13 9 11 11 2
15 9 10 3 13 11 11 11 1 12 7 11 11 1 12 2
25 11 15 13 9 0 13 2 11 11 2 2 15 13 1 11 2 11 11 2 16 9 11 13 9 2
7 16 11 0 2 11 13 2
10 15 13 9 9 1 9 7 9 0 2
36 11 11 11 12 13 9 9 15 13 11 2 11 1 9 12 11 12 1 9 12 2 12 2 12 11 2 12 2 12 2 12 1 9 0 2 2
10 9 10 13 1 9 9 1 9 10 2
20 3 10 13 16 11 13 10 9 9 10 2 9 15 3 13 9 15 15 13 2
46 1 13 11 11 2 11 11 11 15 3 13 9 1 11 2 13 9 11 11 7 9 9 2 10 9 9 15 13 11 1 15 15 13 0 2 1 13 10 9 7 9 1 9 9 2 2
16 11 13 9 9 15 13 1 12 9 11 15 13 11 9 9 2
42 11 11 11 13 1 10 9 2 13 9 9 0 2 9 2 9 9 2 7 9 0 1 9 0 15 13 11 2 3 13 1 11 11 11 2 1 13 9 11 11 11 2
29 9 9 11 9 9 9 13 1 9 1 9 0 2 9 9 9 2 2 1 9 9 9 0 3 0 1 9 9 2
16 11 13 9 1 9 11 2 11 11 11 2 11 11 2 11 2
7 11 14 13 2 15 11 2
35 11 9 3 13 1 11 11 7 9 11 1 9 2 16 9 9 3 13 1 9 11 1 11 0 2 9 2 7 9 9 2 9 11 11 2
17 9 0 3 3 3 13 1 9 2 9 7 9 13 1 9 13 2
83 3 16 2 1 9 13 1 9 12 9 7 0 0 9 2 16 15 0 2 15 13 1 11 11 2 16 1 9 10 9 1 9 11 2 11 2 12 2 12 2 12 2 2 12 2 12 9 2 2 11 2 12 2 12 2 12 2 2 11 11 15 13 1 11 2 11 2 12 2 12 2 12 2 2 11 15 9 2 11 2 12 2 2
19 9 10 3 13 1 9 1 9 9 12 2 15 13 9 7 9 1 13 2
27 9 2 11 2 13 1 13 9 10 1 9 2 1 11 2 2 15 13 1 11 11 1 9 12 2 12 2
20 9 0 11 13 9 11 2 1 9 12 2 12 11 7 12 2 12 9 9 2
27 9 1 11 11 11 11 3 13 1 11 11 2 16 13 11 1 11 16 9 0 1 9 0 1 9 13 2
15 16 13 1 9 12 2 1 0 13 9 13 11 11 11 2
13 3 13 9 9 1 11 11 2 11 11 1 11 2
27 11 14 3 13 1 9 9 7 9 9 2 16 9 9 15 13 1 1 9 7 9 15 0 2 11 2 2
16 11 13 9 11 2 16 13 11 11 2 9 9 12 10 11 2
21 16 9 12 13 9 1 11 11 1 0 2 0 1 9 1 9 9 9 11 11 2
12 11 11 13 1 9 9 2 9 2 7 9 2
23 11 2 9 15 13 1 9 0 1 9 0 9 13 0 9 10 3 3 14 13 9 9 2
25 9 9 5 9 9 3 3 0 15 13 9 2 9 11 11 2 11 9 2 9 9 9 2 9 2
28 1 9 12 2 16 11 12 9 2 11 13 1 9 9 2 13 11 11 7 9 1 12 9 1 9 0 9 2
46 9 9 9 11 11 11 3 13 12 9 0 3 11 11 7 11 11 2 16 1 9 13 9 12 11 12 2 11 11 11 13 12 9 3 9 11 2 11 11 2 11 11 7 11 11 2
11 11 1 9 15 0 13 1 13 9 10 2
6 2 9 2 12 2 2
29 11 11 11 13 10 9 0 9 15 13 1 11 2 11 11 11 11 11 12 11 11 12 2 12 9 11 11 11 2
38 11 11 11 2 11 13 2 9 9 2 7 2 9 0 2 1 11 2 13 1 9 12 11 12 1 9 2 9 11 2 9 11 2 11 11 11 2 2
11 9 10 1 9 13 0 1 9 9 9 2
46 9 1 9 11 2 11 7 11 11 2 9 11 11 15 15 14 0 7 14 13 13 13 1 11 11 2 11 13 13 11 1 9 9 1 12 9 1 11 11 2 7 13 9 1 9 2
17 11 13 9 1 9 11 11 2 11 11 11 2 11 11 2 11 2
13 11 13 16 13 9 3 13 9 0 1 9 11 2
9 15 15 13 1 9 10 14 13 2
28 1 10 13 9 16 9 10 13 9 0 11 15 9 10 3 13 9 2 1 1 9 13 11 11 1 11 11 2
26 9 3 0 13 1 11 11 11 12 2 15 13 1 11 1 12 11 12 1 9 9 2 13 12 9 2
19 11 11 15 3 0 1 11 11 1 0 11 2 11 2 11 2 7 11 2
4 0 9 13 11
12 9 9 9 13 1 9 15 13 1 9 9 2
35 11 11 11 2 2 2 3 13 1 11 11 11 11 11 11 2 2 2 13 10 10 9 15 13 1 11 11 2 11 1 9 0 7 0 2
7 9 10 13 9 9 12 2
10 3 15 13 2 16 10 9 3 13 2
52 11 13 9 9 1 9 12 1 9 15 15 13 2 11 11 11 11 11 7 11 11 11 11 2 16 2 15 3 13 9 15 1 11 11 16 11 13 16 9 15 1 11 11 0 3 13 1 9 0 1 11 2
14 10 9 13 1 9 9 2 3 9 9 1 9 9 2
15 1 12 9 9 9 9 13 9 2 9 2 9 9 13 2
12 9 3 1 9 9 7 1 9 9 7 9 2
37 9 13 3 1 9 2 9 9 9 2 9 2 9 9 2 9 9 9 2 9 9 7 13 9 2 1 3 9 2 9 7 9 2 9 10 9 2
37 16 16 3 3 13 2 15 9 2 9 0 2 1 0 0 16 9 13 10 9 1 9 0 7 1 9 13 9 15 0 1 9 15 0 0 3 2
26 16 9 9 15 0 13 2 9 10 13 16 9 10 13 1 9 9 9 15 0 7 0 15 13 11 2
12 16 12 9 3 2 9 10 3 2 3 13 2
7 7 15 9 1 9 9 2
34 9 10 13 9 1 9 1 9 0 11 11 7 11 11 11 2 11 2 1 13 1 9 1 13 9 9 2 7 13 1 9 2 0 2
14 11 13 9 1 9 11 2 11 11 2 11 2 11 2
8 9 13 1 12 9 1 9 2
30 11 9 10 13 9 0 0 11 2 11 2 11 2 10 9 10 13 2 7 3 13 1 10 9 2 1 9 9 11 2
47 1 10 13 1 9 13 11 5 11 2 1 9 12 11 12 13 3 1 12 9 2 3 2 3 3 13 12 9 11 10 1 9 13 3 9 2 16 0 13 12 11 11 7 12 11 11 2
10 9 10 2 11 13 1 9 11 11 2
26 9 10 15 13 1 9 11 2 15 0 13 1 11 1 9 11 12 1 9 12 11 11 11 9 10 2
6 11 13 13 11 11 2
14 9 9 9 2 1 9 13 9 7 9 1 9 9 2
28 11 11 11 11 11 11 7 9 13 11 7 13 1 11 1 9 12 1 11 13 9 1 15 11 11 11 11 2
33 9 10 13 9 9 15 1 15 13 1 9 9 2 11 11 2 15 13 1 10 9 9 9 1 3 3 13 10 10 10 1 11 2
38 11 11 13 16 15 3 13 9 9 11 1 2 11 11 2 2 16 13 9 9 11 7 9 13 1 9 2 1 13 1 10 3 13 9 1 9 12 2
12 9 10 3 11 11 11 13 1 0 9 12 2
9 1 11 11 3 13 1 9 9 2
19 2 11 11 11 2 15 0 13 13 1 9 0 2 9 2 1 9 11 2
11 11 10 3 13 1 9 11 0 1 9 2
18 11 11 13 9 15 13 1 11 11 11 2 11 11 2 11 2 11 2
10 11 2 11 13 10 9 15 3 13 2
11 11 9 10 3 13 10 9 9 1 0 2
9 16 11 13 15 13 9 1 9 2
18 3 0 3 15 3 13 1 9 11 11 2 3 3 1 0 9 13 2
21 9 15 13 2 13 9 16 3 1 9 9 7 9 9 0 2 13 1 9 9 2
10 9 12 7 9 13 1 12 11 12 2
10 11 11 13 9 15 3 0 1 11 2
27 1 0 9 2 11 2 13 10 9 15 13 9 10 1 13 9 2 9 15 13 1 13 10 9 11 0 2
21 9 2 9 9 1 9 13 1 11 11 2 16 13 9 2 9 0 7 13 9 2
28 1 10 9 9 15 0 2 11 11 13 9 0 1 13 7 13 10 9 7 9 16 13 1 9 2 9 10 2
29 9 9 9 1 9 2 13 1 9 2 9 9 2 16 9 9 3 13 2 13 9 9 2 9 15 3 13 9 2
15 11 9 9 12 9 3 13 9 2 9 1 1 9 9 2
5 2 15 13 9 2
17 11 7 9 2 9 9 3 13 1 9 11 11 11 1 13 9 2
18 11 11 1 11 3 13 1 11 3 10 1 3 13 7 13 11 11 2
6 11 13 10 9 15 2
22 11 11 13 1 12 9 16 2 11 11 2 11 11 2 11 11 2 11 2 7 11 2
21 9 10 14 13 9 9 15 3 3 16 3 13 0 1 9 2 9 15 3 0 2
23 1 12 2 11 11 12 13 12 9 0 7 12 9 0 2 13 9 9 9 1 12 9 2
20 9 11 13 9 13 9 15 13 1 11 7 13 1 9 1 9 12 1 12 2
29 9 11 11 11 13 1 9 12 2 3 1 9 11 13 9 9 11 11 11 11 11 15 0 13 1 11 11 11 2
14 9 10 13 9 9 1 9 15 3 0 1 10 9 2
12 11 9 1 9 11 13 2 9 15 0 2 2
16 9 16 12 9 15 13 1 11 3 13 9 7 9 15 0 2
30 9 10 13 1 9 0 11 11 11 11 11 2 12 9 2 1 9 0 15 13 1 10 9 3 1 9 11 2 11 2
8 13 1 9 11 2 11 11 2
13 1 1 2 15 3 13 9 9 0 1 10 11 2
8 11 13 10 10 9 15 13 2
10 9 12 13 9 9 11 11 1 9 2
39 7 11 13 10 9 15 13 1 9 9 2 15 13 9 1 9 9 1 11 7 13 9 1 9 11 2 13 9 9 12 5 12 9 15 3 13 1 11 2
23 15 15 3 13 3 13 13 9 0 1 11 13 13 1 13 9 0 2 11 2 9 11 2
14 11 13 9 1 11 11 2 11 2 11 11 2 11 2
42 1 9 10 2 11 11 3 13 1 11 11 11 2 1 3 9 11 11 3 13 15 1 11 11 11 1 9 11 11 7 13 9 9 11 13 11 16 15 13 9 11 2
14 11 13 1 11 1 10 9 1 11 7 11 1 11 2
12 13 12 5 2 12 9 2 1 9 9 11 2
25 11 13 1 11 9 1 9 11 11 2 2 1 9 11 11 2 15 13 9 9 1 9 9 11 2
26 11 11 11 2 11 2 2 2 13 9 11 11 13 11 11 2 9 11 1 9 9 9 0 7 9 2
17 11 13 9 9 1 9 11 11 2 3 13 9 9 1 9 10 2
19 9 10 3 13 1 9 1 13 9 0 7 13 9 0 1 9 2 9 2
16 9 2 9 0 1 1 9 2 9 2 9 2 9 2 9 2
13 1 10 2 12 13 3 3 13 9 9 1 9 2
69 7 9 9 0 1 9 9 12 9 1 1 11 11 2 11 11 11 2 11 11 11 2 11 2 2 11 11 2 11 9 11 2 11 11 11 2 11 11 11 2 7 11 11 2 11 11 11 2 11 11 11 2 11 13 10 10 9 9 0 1 11 15 3 13 9 9 9 0 2
21 1 9 12 2 11 13 9 12 11 11 2 10 13 15 13 3 9 13 9 1 2
11 16 2 3 10 9 13 9 2 11 2 2
10 1 9 11 2 15 13 1 9 0 2
126 9 9 13 9 13 0 1 9 3 11 2 11 11 2 11 2 11 2 11 2 11 2 11 11 11 11 11 2 11 2 11 2 9 2 11 2 11 2 11 2 11 2 11 11 2 11 2 11 2 11 11 7 11 13 9 11 11 7 11 11 11 11 11 2 9 9 10 13 1 12 11 12 2 9 10 9 10 13 9 9 11 2 11 0 1 9 11 7 11 13 1 9 1 9 9 2 9 0 1 9 2 9 9 1 13 9 7 9 9 1 9 7 9 11 11 11 11 13 9 1 13 9 11 15 13 2
19 15 13 1 11 2 2 9 9 2 9 9 2 16 15 13 15 0 10 2
7 9 0 3 3 12 9 2
22 11 11 11 2 9 9 9 15 0 13 10 9 9 9 0 15 14 0 13 2 8 2
41 9 10 13 1 9 2 9 15 13 9 2 9 9 11 7 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 7 3 10 3 2
38 11 2 9 10 13 1 9 9 1 13 9 15 0 2 9 9 0 2 9 9 9 7 9 9 9 2 9 0 2 7 9 0 9 11 1 13 9 2
50 1 13 10 11 1 10 9 2 10 9 9 13 1 11 11 11 2 11 1 11 11 2 1 11 11 11 2 11 2 15 13 9 11 1 9 10 7 10 9 0 15 13 1 13 9 0 1 9 9 2
16 9 10 13 0 3 1 11 11 2 15 3 13 9 9 9 2
8 11 9 15 0 7 0 9 2
32 11 11 13 9 2 9 0 1 10 9 1 11 11 2 1 12 2 7 13 12 1 1 12 2 11 11 2 1 1 11 11 2
18 3 11 7 11 3 13 9 15 15 13 9 9 0 15 13 1 10 2
13 16 3 2 3 13 2 11 13 1 11 7 11 2
27 11 12 5 3 13 1 9 12 5 16 10 9 0 9 13 9 1 9 2 3 3 13 7 13 1 11 2
19 1 9 2 9 9 9 2 9 9 1 9 9 2 9 9 7 9 13 2
6 11 1 10 9 2 2
29 11 11 11 13 9 9 2 1 9 1 11 11 7 9 2 9 11 1 1 11 11 2 11 2 11 2 7 11 2
43 11 11 13 9 0 1 9 9 1 9 11 1 1 11 7 11 2 13 9 9 11 11 15 13 1 11 1 12 2 1 9 11 3 15 13 1 11 16 3 13 1 9 2
11 11 13 9 9 0 15 13 0 7 0 2
26 2 11 11 2 1 9 11 2 13 9 9 15 13 1 9 9 11 2 9 11 2 11 1 9 12 2
14 11 11 13 9 1 11 11 2 11 2 11 2 11 2
25 11 0 15 13 9 2 11 11 11 11 2 11 2 2 2 7 9 13 1 0 1 12 11 12 2
17 11 11 11 13 13 7 13 1 9 11 11 11 11 2 11 2 2
20 9 9 13 9 9 9 15 13 1 9 1 9 2 9 2 9 7 9 0 2
9 9 10 13 1 9 9 1 12 2
31 1 10 2 11 11 3 13 11 12 9 2 2 7 11 11 2 1 12 11 12 2 15 3 13 13 11 2 13 11 11 11
18 9 12 11 11 13 9 11 1 9 11 16 9 7 9 1 9 9 2
13 11 11 11 12 9 13 9 12 1 9 12 9 2
14 11 13 9 1 9 11 2 11 2 11 11 2 11 2
14 11 11 13 1 10 9 15 13 9 2 9 1 9 2
57 11 11 2 11 11 11 11 11 2 11 11 11 11 2 11 11 11 11 11 2 11 11 11 2 11 11 11 2 11 11 11 11 11 12 2 12 5 11 11 11 12 2 12 5 11 11 11 11 12 2 12 5 11 12 2 12 5
49 3 13 1 9 11 2 11 11 1 9 9 12 2 12 1 12 2 12 15 13 1 11 11 2 1 9 11 11 2 11 11 2 15 13 1 11 11 13 1 9 9 12 2 12 1 12 2 12 2
47 1 12 11 12 2 11 13 9 9 9 1 11 15 13 1 9 12 9 9 9 11 11 2 16 9 13 7 9 3 13 9 9 9 2 11 13 9 16 11 11 11 2 11 13 9 9 2
7 9 9 11 10 3 13 2
11 15 14 13 7 13 16 13 9 13 0 2
77 9 13 10 9 9 9 11 3 0 11 13 9 1 13 2 1 0 2 2 9 2 5 5 8 2 8 2 8 5 8 5 8 5 8 5 8 2 8 11 3 13 12 9 7 9 9 11 11 13 1 9 9 9 9 9 2 15 9 9 13 9 11 2 11 2 1 10 9 9 9 9 0 1 12 9 12 2
18 1 16 10 13 15 13 1 1 2 13 15 1 7 13 15 13 1 2
65 9 9 9 0 1 12 13 12 2 12 5 2 13 1 11 1 12 16 9 13 1 12 2 12 5 1 11 11 2 9 7 9 1 12 2 12 5 7 9 1 12 2 12 5 2 9 0 2 0 9 1 12 1 9 9 2 10 9 15 3 13 1 9 0 2
29 1 0 9 15 13 9 1 9 9 2 1 11 2 7 15 13 9 7 13 1 9 0 2 1 9 1 9 9 2
23 10 9 13 12 9 10 2 11 11 11 11 2 2 2 11 11 11 2 7 2 11 2 2
7 11 2 11 3 13 9 2
8 7 3 3 3 0 1 11 2
35 11 16 13 9 9 9 0 11 7 11 11 13 13 10 10 1 9 13 9 0 0 9 9 15 3 13 1 11 11 13 1 9 9 9 2
33 16 13 9 9 9 9 2 11 2 11 11 7 13 1 11 11 12 2 0 9 11 11 2 11 2 10 3 13 1 11 11 12 2
35 10 9 9 15 0 7 10 16 7 2 11 11 2 11 11 9 2 11 12 2 2 11 11 11 2 9 9 9 11 2 2 7 11 11 2
14 11 13 9 0 15 3 0 2 3 11 11 11 11 2
24 1 9 12 2 15 13 12 9 9 0 7 15 3 0 1 9 11 0 15 3 13 9 9 2
24 11 11 13 10 10 9 15 13 1 11 11 11 11 2 9 11 11 2 11 11 11 2 11 2
30 11 11 11 13 2 9 9 2 2 7 9 13 12 9 9 7 10 9 15 16 15 13 9 1 11 1 9 3 13 2
19 9 0 13 9 1 11 11 11 2 9 10 1 9 13 9 9 11 11 2
24 11 11 13 10 9 9 11 11 2 1 9 11 11 11 2 1 11 11 1 9 12 2 12 2
14 14 15 10 13 1 9 0 2 16 15 3 13 15 2
35 11 10 13 1 9 0 11 12 2 11 2 1 9 9 2 11 13 1 13 11 7 3 2 9 2 11 11 13 1 11 7 11 13 0 2
26 16 9 0 13 1 11 1 11 2 11 13 1 11 1 9 9 15 3 13 1 15 3 13 1 9 2
16 14 9 9 11 7 11 0 9 2 9 7 9 9 3 3 2
11 9 9 10 13 9 1 2 11 11 2 2
14 11 15 13 9 12 11 11 3 2 3 13 1 9 2
31 1 9 2 9 2 9 7 9 1 9 1 10 9 7 9 2 16 9 11 11 12 13 10 9 9 9 11 11 9 11 2
9 16 14 0 13 2 13 11 11 2
11 11 11 14 13 9 2 9 15 13 9 2
11 11 13 9 15 13 1 11 11 2 11 2
14 9 10 13 9 0 1 10 9 7 9 1 9 9 2
20 11 2 9 2 13 1 9 9 9 2 9 9 15 13 2 13 1 9 2 2
23 9 10 13 9 1 11 2 10 9 1 12 9 1 0 11 2 15 3 13 13 1 11 2
11 14 15 9 0 2 2 0 15 9 0 2
63 1 9 16 9 3 13 1 9 2 11 2 11 11 9 2 13 9 9 9 9 1 13 9 1 10 11 11 2 11 1 9 5 9 9 13 9 0 1 9 10 11 16 13 9 0 3 13 9 9 5 9 9 15 3 13 2 13 9 2 1 9 10 2
17 11 13 10 9 9 1 9 11 11 2 9 11 2 11 11 11 2
12 9 12 13 12 9 3 2 3 1 9 12 2
37 9 10 1 13 1 9 11 11 11 2 16 13 3 13 9 2 9 7 9 2 3 1 13 9 9 9 9 15 3 1 13 1 9 2 9 0 2
47 11 11 12 13 11 11 11 9 11 11 11 2 9 11 11 2 1 11 11 2 9 2 7 13 12 9 9 2 3 2 12 2 11 11 12 2 12 2 11 11 2 7 12 2 11 11 2
15 11 3 3 13 9 9 9 15 13 7 13 1 9 9 2
40 9 9 13 9 9 9 1 9 11 15 13 1 9 9 12 12 15 13 1 13 9 11 1 9 11 2 13 9 10 9 2 3 13 1 9 0 7 9 0 2
23 3 2 11 10 13 1 13 9 1 13 16 14 3 13 11 10 7 15 13 9 1 9 2
21 11 9 1 9 2 12 2 12 5 9 2 1 9 9 13 0 2 0 2 9 2
44 15 13 11 11 11 2 11 11 11 2 11 11 11 2 7 11 11 11 11 11 2 1 10 2 13 10 9 3 13 11 15 3 13 2 13 0 2 3 11 11 11 2 11 2
25 16 1 9 9 2 9 0 2 0 13 9 0 2 7 13 1 1 9 9 9 2 9 0 2 2
16 11 11 2 9 11 11 11 2 7 11 11 3 13 9 10 2
21 16 9 0 16 9 3 13 2 16 9 10 3 13 9 7 9 15 3 13 9 2
21 15 13 9 9 9 11 15 13 1 11 11 1 9 1 9 1 9 12 11 12 2
7 3 9 3 13 9 0 2
41 11 11 11 2 2 12 11 12 2 12 11 12 2 13 9 9 11 11 15 0 15 0 1 9 11 2 11 11 11 7 11 2 7 3 11 11 7 11 11 11 2
55 11 11 2 2 13 10 9 9 9 11 11 15 13 3 1 9 9 1 9 2 9 9 9 2 7 9 10 15 3 13 9 1 12 9 11 11 2 1 11 11 15 3 13 9 1 9 11 11 2 1 9 11 11 11 2
14 9 9 11 11 15 0 10 13 5 13 1 11 11 2
18 13 3 2 3 1 13 9 2 16 13 1 9 3 3 9 15 13 2
14 11 13 9 1 11 11 2 7 2 11 11 2 11 2
5 13 15 13 0 2
15 9 9 13 1 9 9 7 9 12 3 13 0 7 0 2
11 11 16 15 13 12 9 1 9 0 11 2
10 9 9 13 1 12 11 12 1 11 2
19 11 13 10 10 9 1 11 11 2 11 11 11 2 11 11 11 2 11 2
14 11 13 9 1 9 11 2 11 2 11 11 2 11 2
9 9 10 13 1 11 11 2 11 2
12 9 9 1 9 2 9 7 9 0 13 0 2
8 16 9 3 14 13 9 0 2
13 1 9 9 9 13 1 13 1 9 12 1 9 2
35 16 13 1 11 11 11 11 2 11 13 9 1 13 9 1 11 11 2 15 13 9 7 13 11 11 2 11 11 2 7 11 11 1 13 2
11 11 0 1 9 10 13 11 11 7 11 2
24 1 11 11 3 2 11 11 12 2 15 13 9 12 7 13 1 11 2 11 11 1 9 0 2
8 15 3 3 13 9 10 9 2
12 9 10 13 0 7 0 13 1 9 2 9 2
16 9 10 12 9 13 1 9 9 9 1 11 11 1 9 12 2
7 9 13 3 0 1 11 2
13 10 9 9 13 11 11 11 11 11 13 9 10 2
63 10 9 11 3 13 9 11 2 11 7 11 1 9 2 7 9 11 3 3 13 9 11 11 11 2 11 2 1 9 9 1 9 9 1 9 12 2 7 0 9 9 10 9 15 3 0 2 9 9 9 0 1 11 3 13 2 3 1 9 2 9 0 2
14 11 13 7 13 9 9 16 9 9 13 13 9 9 2
16 1 3 9 2 10 9 9 13 1 11 7 13 1 9 11 2
15 11 2 11 2 3 13 15 9 9 13 9 1 3 0 2
10 15 3 13 9 9 13 0 0 0 2
10 9 15 13 9 10 2 11 3 13 2
43 1 9 9 10 13 1 12 9 0 2 16 9 7 9 15 13 9 0 1 13 3 1 13 9 0 15 13 9 1 9 2 9 7 9 9 0 1 13 9 3 3 3 2
23 11 13 10 10 9 15 13 1 11 11 11 2 11 11 11 2 11 11 11 11 2 11 2
12 9 9 0 0 13 1 9 9 9 11 11 2
18 11 1 11 11 13 9 15 3 13 3 13 1 9 15 13 13 9 2
10 13 1 9 13 13 9 1 9 12 2
10 1 9 13 2 9 13 1 9 0 2
24 11 13 10 10 9 15 13 1 11 11 2 11 11 11 2 11 11 11 2 11 11 2 11 2
22 9 9 13 9 9 9 11 9 12 2 7 3 13 12 5 9 9 10 1 9 12 2
17 15 13 12 9 1 9 0 7 13 9 2 9 2 7 9 9 2
16 3 13 15 1 9 9 9 0 2 3 13 15 1 1 9 2
53 1 10 3 11 11 7 9 9 10 2 1 2 11 11 11 11 2 11 2 11 11 11 2 11 11 11 11 2 11 2 11 11 11 11 2 11 2 11 11 11 11 11 2 7 3 3 9 9 0 15 3 10 2
23 11 9 11 11 11 11 2 11 13 16 10 9 11 15 13 1 12 14 13 3 9 9 2
13 1 9 10 15 13 1 9 11 11 11 1 9 2
58 11 13 10 9 1 9 7 9 2 9 2 10 9 9 2 7 0 1 9 15 3 15 13 1 9 1 10 9 15 0 13 2 16 15 13 9 1 1 10 9 15 3 0 2 1 9 11 1 11 2 15 13 2 7 11 1 11 2
38 1 13 9 2 11 2 11 7 11 3 13 7 13 1 11 2 1 11 2 11 15 0 13 10 9 9 1 1 9 0 2 9 2 11 2 3 13 2
7 15 13 13 10 9 0 2
153 1 1 9 0 9 11 11 13 9 9 11 2 11 2 1 11 2 11 2 13 2 7 9 9 11 2 11 2 7 11 2 11 2 7 14 11 2 11 2 2 9 9 9 13 2 9 2 11 11 2 1 1 11 2 11 11 2 14 13 2 2 7 14 2 11 2 11 11 2 1 1 11 2 11 2 2 9 2 9 0 10 3 13 1 9 11 11 2 9 2 9 9 11 2 11 2 11 5 2 11 2 12 12 12 12 12 9 2 9 2 9 2 5 12 2 2 2 2 11 5 2 11 2 12 5 5 2 9 2 9 2 0 2 9 2 9 0 5 12 2 11 2 11 2 5 11 2 2 2 11 11 9 2
19 11 11 13 10 10 9 1 11 11 11 2 11 11 2 11 11 2 11 2
11 11 13 3 11 3 13 9 1 13 1 2
20 11 13 1 9 15 3 3 13 1 9 2 1 9 12 9 9 11 13 9 2
10 9 3 13 2 3 13 1 9 9 2
16 9 12 11 12 2 11 13 9 1 9 9 11 11 2 15 2
11 9 10 13 9 11 11 7 11 11 11 2
22 9 9 7 15 0 15 3 13 9 1 11 2 3 13 9 0 15 13 1 9 0 2
18 9 9 9 15 13 11 1 9 13 9 9 0 15 13 0 7 0 2
8 10 9 9 11 13 1 12 2
14 9 2 15 13 2 9 9 1 9 15 13 9 0 2
16 10 9 3 13 15 13 9 2 9 2 1 9 7 9 0 2
21 11 11 13 9 9 9 1 9 11 11 2 11 11 11 2 11 11 11 2 11 2
23 11 11 13 1 9 2 9 15 3 13 9 1 9 11 2 7 3 13 9 0 16 10 2
21 1 9 10 15 13 9 1 10 9 0 1 11 7 13 9 10 9 11 11 12 2
14 9 9 15 13 1 11 11 13 9 1 11 7 9 2
11 11 13 11 1 10 9 9 1 9 0 2
10 3 9 11 16 15 13 9 0 9 2
13 11 11 12 11 13 9 0 1 11 11 12 11 2
9 3 11 11 13 3 1 9 11 2
14 1 9 9 10 2 11 11 11 3 10 9 13 9 2
37 11 3 3 13 1 9 0 2 7 3 2 3 13 1 9 0 1 9 9 11 11 7 1 9 2 1 1 9 2 11 2 7 2 11 2 2 2
41 9 9 13 16 9 10 13 16 10 9 9 2 9 11 10 13 1 9 9 15 0 1 1 9 9 1 9 1 2 11 11 2 2 9 2 15 13 9 9 9 2
13 11 13 1 9 0 9 7 9 12 2 11 11 2
26 1 9 1 9 0 2 9 13 1 10 9 9 9 9 2 7 1 9 7 1 9 9 11 1 11 2
38 11 2 11 11 11 7 11 2 9 11 2 11 11 11 7 9 9 2 13 9 9 7 9 0 11 2 7 9 9 0 9 10 1 9 9 7 9 2
22 3 9 0 2 12 5 2 15 13 1 9 11 2 11 2 7 9 9 2 13 9 2
50 9 9 9 10 13 1 11 11 11 15 0 1 2 11 11 11 2 1 11 11 11 2 11 11 7 11 11 11 2 9 12 13 2 11 11 11 2 16 1 9 9 2 9 10 15 3 13 12 9 2
12 1 1 9 3 2 15 13 1 11 2 11 2
28 11 11 2 9 11 2 11 11 2 13 9 12 0 1 9 10 9 9 1 11 15 13 1 10 11 7 11 2
23 9 10 13 9 1 9 11 7 9 11 2 15 13 16 9 13 1 9 9 7 9 9 2
52 11 7 9 9 15 3 13 13 9 9 9 15 13 9 9 2 1 11 2 9 9 1 9 14 13 13 9 7 13 1 10 9 2 7 9 9 9 15 0 1 9 9 7 9 9 3 13 7 13 1 9 2
18 11 13 1 9 0 2 2 2 2 11 11 13 12 2 12 1 0 2
25 3 13 9 11 15 0 13 16 13 1 11 2 11 11 2 11 13 1 9 9 9 11 11 11 2
22 9 11 12 2 11 13 1 9 9 1 11 11 5 11 2 9 9 1 11 2 11 2
9 10 9 3 15 13 0 1 0 2
6 10 9 11 13 9 2
28 9 9 13 10 13 1 9 15 7 3 13 1 9 9 15 13 9 9 10 9 7 2 9 10 9 9 2 2
25 16 10 9 13 2 10 9 13 14 9 1 13 9 15 2 3 13 9 9 11 1 9 0 11 2
29 11 9 10 13 1 9 9 11 11 11 11 11 15 7 1 9 11 11 11 11 11 11 11 3 1 11 11 11 2
41 16 11 7 11 3 13 13 2 16 2 9 15 3 13 16 11 3 13 9 1 9 9 9 11 13 9 9 15 13 10 9 9 9 16 3 13 1 9 9 9 2
10 9 9 10 13 7 13 1 11 11 2
29 10 9 2 9 1 9 9 2 15 13 1 9 11 13 13 9 9 1 9 9 0 7 9 9 15 13 1 11 2
10 10 2 10 9 3 13 9 15 0 2
13 15 13 9 9 15 14 13 2 13 1 9 11 2
16 9 11 13 1 9 9 15 3 0 1 13 9 9 9 13 2
16 12 12 9 3 13 3 13 9 0 15 13 1 9 11 11 2
10 13 13 3 2 9 13 9 9 9 2
18 11 11 3 13 1 11 11 2 9 15 13 1 11 11 11 1 12 2
15 11 11 12 13 10 9 1 11 11 2 11 11 2 11 2
11 1 9 0 1 9 7 9 2 13 11 2
22 11 11 13 10 10 9 15 13 1 11 11 11 2 11 9 2 11 11 11 2 11 2
24 9 1 9 9 13 1 9 9 9 12 3 9 0 15 13 12 9 7 12 9 7 12 9 2
29 9 10 13 1 11 11 12 1 13 9 11 2 7 1 9 12 1 9 11 2 15 3 13 1 11 11 9 12 2
13 11 13 9 15 13 1 9 11 1 11 2 11 2
28 11 11 11 11 2 9 11 11 2 13 9 15 13 9 9 7 9 9 15 13 11 11 1 11 2 11 11 2
20 11 11 13 10 10 9 1 11 11 11 2 11 11 2 11 11 11 2 11 2
28 0 9 11 2 3 15 13 0 2 13 9 11 0 0 1 9 11 7 11 7 9 11 0 1 9 11 11 2
12 11 3 3 13 9 9 1 11 7 9 9 2
47 1 13 9 10 2 11 13 1 9 0 1 11 11 2 11 11 11 2 9 9 1 11 11 11 11 2 2 11 11 11 11 2 7 3 9 0 0 15 13 1 11 11 11 2 11 2 2
21 13 3 12 12 9 1 9 11 11 9 12 2 9 0 9 10 13 9 9 10 2
15 11 13 1 9 15 13 0 1 0 9 9 9 11 10 2
16 11 0 10 13 3 1 12 9 9 2 1 1 13 9 9 2
30 9 9 9 15 3 0 13 12 2 12 11 2 1 15 13 1 9 9 2 2 16 9 0 13 1 12 2 12 11 2
15 13 11 11 15 13 1 11 11 9 11 1 11 7 11 2
27 1 9 10 13 1 9 9 9 11 13 11 11 13 1 9 9 11 1 9 11 2 11 11 1 9 12 2
23 9 9 7 9 9 10 13 13 1 9 11 11 11 2 15 13 1 9 9 12 2 12 2
7 11 11 13 9 12 1 11
22 7 3 13 9 1 11 11 2 15 14 3 13 9 1 9 9 16 3 13 9 9 2
31 1 7 10 2 9 9 9 14 3 13 7 16 9 10 9 13 16 10 0 1 13 9 9 7 15 14 13 1 13 9 2
15 16 12 9 15 13 10 9 13 9 2 15 13 1 0 2
10 11 11 1 13 9 11 13 1 0 2
12 1 9 0 9 2 9 14 13 9 15 0 2
22 11 9 13 1 12 9 12 15 3 13 7 13 9 9 15 13 1 1 9 9 9 2
8 3 11 7 11 13 9 15 2
15 12 13 1 9 12 2 3 13 12 9 2 1 12 9 2
39 16 2 1 9 0 2 13 1 11 11 2 1 0 15 13 11 11 7 11 11 1 9 12 2 12 2 12 2 12 2 12 2 12 7 13 9 1 11 2
10 11 11 3 13 9 1 9 15 0 2
30 15 0 13 11 11 7 9 11 1 1 9 3 13 1 0 2 9 9 13 7 9 7 9 7 9 1 3 13 9 2
18 11 11 13 10 10 9 1 11 11 2 11 11 2 11 11 2 11 2
30 1 9 9 7 0 2 9 0 9 7 9 3 3 13 1 13 1 9 9 0 1 13 9 9 7 9 7 9 0 2
14 11 13 9 1 11 11 2 11 2 11 11 2 11 2
31 9 10 13 9 9 9 13 3 0 2 1 9 9 9 2 9 15 13 3 13 1 3 0 7 0 1 13 9 9 9 2
10 3 11 11 3 3 3 13 9 9 2
15 9 0 9 13 9 16 10 9 15 13 13 10 9 9 2
25 11 11 2 9 9 9 1 9 2 13 16 7 9 11 2 11 3 13 9 9 9 1 13 9 2
20 9 9 11 9 13 9 2 2 9 9 0 2 2 1 10 9 9 13 0 2
23 9 11 11 13 10 10 9 15 13 1 11 11 11 2 11 9 11 2 11 11 2 11 2
5 15 3 3 13 2
18 1 0 2 11 11 3 13 0 1 11 1 9 0 7 9 9 9 2
12 9 9 3 1 9 9 8 5 8 9 11 2
10 11 13 12 9 15 13 1 9 10 2
16 1 9 9 9 9 9 2 9 9 9 3 13 7 13 9 2
15 11 11 13 13 11 11 7 9 7 9 15 0 7 0 2
10 9 11 13 9 1 3 13 1 9 2
45 9 10 3 13 9 9 9 7 9 2 9 0 1 13 1 9 2 9 11 11 11 2 1 16 10 1 1 9 10 13 3 9 2 9 11 2 11 7 9 15 13 1 9 9 2
10 16 0 2 9 11 3 13 9 0 2
13 10 9 9 11 13 9 10 2 3 14 1 13 2
22 11 2 9 11 2 11 2 7 9 13 9 0 16 3 0 1 9 9 2 9 2 2
21 1 9 9 2 7 3 3 13 9 9 2 13 9 11 11 2 15 9 11 13 2
11 11 13 13 9 1 13 7 13 9 10 2
53 9 15 3 13 1 9 11 1 9 1 10 13 9 9 11 11 11 16 11 2 11 11 11 2 15 13 10 10 9 9 11 11 7 3 13 1 9 1 9 12 2 12 2 7 10 10 9 0 14 11 11 11 2
28 11 2 12 2 12 3 13 3 9 9 1 9 11 11 2 9 9 9 11 15 3 3 13 9 11 1 9 2
15 15 3 13 1 9 11 2 12 7 11 2 12 1 11 2
30 11 15 3 2 13 1 9 0 13 9 11 0 13 9 1 13 1 9 9 7 13 1 10 9 1 11 7 9 9 2
11 15 13 1 11 11 11 1 11 11 11 2
42 11 3 13 9 9 15 3 3 2 12 2 12 9 2 13 9 15 3 0 2 11 11 2 2 9 0 12 12 15 3 13 2 9 3 0 2 9 3 0 7 0 2
6 11 11 13 12 9 2
10 16 10 9 10 9 9 13 9 11 2
25 9 9 11 13 1 9 12 11 12 1 11 11 2 11 2 9 10 15 3 13 11 2 11 2 2
8 11 10 13 1 9 11 11 2
74 11 11 1 11 7 11 11 2 9 1 11 11 11 11 2 13 9 1 9 9 11 15 3 0 13 11 11 11 2 9 11 11 1 11 3 13 1 9 12 11 2 12 9 1 9 11 2 15 13 9 0 3 13 9 11 2 7 9 12 11 12 2 9 0 9 11 1 1 9 9 11 11 2 2
27 9 15 0 2 3 13 1 11 11 11 2 3 3 14 9 1 0 15 3 0 1 9 9 7 9 0 2
15 9 2 11 11 5 10 9 3 2 11 13 9 9 0 2
27 11 11 2 13 12 9 12 7 11 11 2 13 9 11 7 9 11 11 11 2 11 11 11 2 1 12 2
19 11 10 13 13 12 9 1 9 12 7 13 3 13 1 12 1 9 0 2
9 16 0 9 1 9 9 11 11 2
32 11 11 11 3 13 9 3 13 11 11 16 13 9 11 12 11 11 9 12 1 0 13 1 9 11 11 11 11 1 9 12 2
15 1 12 9 13 1 1 11 11 2 12 9 3 13 13 2
13 3 2 9 15 13 1 15 15 3 0 1 9 2
55 7 3 10 11 3 13 1 13 9 10 9 1 9 9 15 0 2 1 9 2 9 7 9 7 9 2 1 9 15 0 7 9 15 13 7 1 9 15 0 2 1 15 13 11 2 11 2 9 1 11 2 1 9 9 2
47 1 15 13 1 9 2 11 11 13 9 1 9 2 9 10 15 13 9 0 7 13 1 9 11 2 15 3 13 1 2 9 9 2 1 9 9 2 7 1 0 1 9 2 11 11 11 2
14 11 11 13 9 1 10 10 9 9 9 1 9 11 2
17 15 13 9 11 7 9 9 2 11 11 2 13 9 1 9 11 2
14 9 15 3 13 1 2 10 9 11 2 7 3 9 2
12 11 11 11 11 11 2 2 13 9 0 11 2
18 11 11 11 13 9 0 7 9 0 1 12 9 2 9 2 5 2 2
25 11 3 3 14 3 3 13 9 1 9 11 11 7 11 11 2 7 3 13 9 1 11 7 11 2
31 9 0 2 12 2 2 11 7 9 9 11 11 13 9 9 1 11 13 1 11 11 2 7 9 11 11 13 1 11 11 2
21 11 11 13 10 12 9 15 13 1 11 11 2 11 11 11 2 9 11 2 11 2
11 11 11 13 3 2 16 13 9 9 11 2
17 9 10 3 13 1 13 9 9 9 9 2 9 13 1 9 11 2
11 11 10 3 3 13 13 9 0 7 9 2
12 9 10 13 1 11 11 7 9 9 11 11 2
30 0 9 15 3 13 0 1 3 9 13 11 11 2 11 11 11 2 11 11 2 9 2 7 11 11 2 9 9 2 2
5 9 9 9 9 2
23 11 10 13 9 7 11 11 13 9 10 1 13 9 9 0 3 0 9 10 2 11 11 2
14 11 13 9 1 11 11 2 11 2 11 11 2 11 2
12 1 9 12 2 9 10 13 9 1 12 9 2
26 3 15 13 9 15 7 9 9 15 3 0 2 11 13 12 9 12 2 16 11 13 12 11 12 2 2
16 11 2 2 13 9 9 9 11 1 11 15 3 13 9 11 2
6 9 15 13 9 10 2
8 11 0 13 9 9 9 9 2
17 11 9 0 15 3 0 13 9 9 2 9 9 1 9 3 0 2
15 11 9 3 13 1 13 9 0 7 15 9 0 7 0 2
13 11 11 7 11 13 9 15 1 13 3 9 9 2
39 9 10 1 13 11 7 11 11 3 13 9 11 11 15 3 13 1 11 1 13 9 9 11 11 15 13 1 9 7 9 1 9 0 1 11 2 11 2 2
30 2 12 9 15 0 0 7 0 3 1 9 13 9 0 11 2 15 3 13 1 9 0 1 11 11 7 11 11 11 2
50 3 10 9 13 1 9 9 2 16 9 2 9 15 13 9 10 2 9 10 13 9 1 9 9 15 13 10 9 2 11 11 3 13 1 9 9 7 3 13 12 9 2 7 13 9 13 0 1 11 2
16 15 14 3 13 9 2 16 3 13 13 1 12 9 1 12 2
10 11 11 3 2 3 3 13 1 11 2
15 10 9 1 9 10 13 9 11 2 11 1 9 9 15 2
22 9 1 9 15 13 1 9 11 11 2 7 13 1 9 12 1 9 11 1 9 0 2
13 9 0 15 2 11 11 10 2 13 1 9 12 2
12 15 3 13 9 9 14 2 2 3 9 11 2
16 9 10 13 1 9 9 0 11 0 15 3 13 1 11 11 2
15 9 11 11 11 3 13 9 9 1 11 11 7 11 11 2
35 11 11 11 11 11 11 1 9 10 2 11 11 15 13 1 12 3 13 9 11 2 11 11 13 10 10 9 15 3 13 1 11 11 11 2
14 1 13 9 2 15 13 1 9 10 13 9 15 13 2
34 9 10 1 12 9 13 16 13 9 9 9 9 2 16 1 9 0 16 14 13 1 0 3 13 9 15 0 1 9 9 7 9 9 2
14 9 1 9 2 9 2 9 2 9 0 7 9 9 2
105 1 9 12 11 7 11 13 13 11 1 0 1 11 2 1 9 12 2 11 13 1 11 11 2 10 9 0 11 11 11 2 1 13 7 13 9 9 11 1 11 5 11 2 1 9 3 0 9 11 13 1 11 2 7 9 0 15 0 2 14 0 1 11 2 1 9 12 2 9 11 11 11 7 11 11 13 9 1 9 11 2 15 13 1 2 9 2 2 7 9 1 9 9 9 0 3 13 2 13 1 2 9 9 2 2
33 11 11 13 9 3 12 11 2 1 9 10 13 9 0 2 14 13 9 9 2 2 11 11 10 13 1 12 9 9 3 2 12 2
64 9 10 3 13 9 9 0 0 15 13 3 1 13 9 0 1 9 1 13 9 9 2 13 3 9 1 9 2 11 11 2 11 13 13 1 9 9 15 13 9 2 9 1 3 2 11 2 9 15 3 0 13 3 13 0 7 13 9 1 9 7 9 0 2
20 11 11 13 12 9 9 10 9 2 1 9 1 12 5 2 15 13 9 0 2
29 11 11 11 12 2 12 13 9 0 11 11 11 2 1 9 9 3 13 1 9 11 11 15 3 13 1 12 9 2
21 11 11 13 3 12 9 1 9 9 11 2 11 11 11 2 11 11 11 2 11 2
3 1 9 2
20 16 1 9 10 15 13 1 9 9 2 11 11 2 11 11 15 13 11 11 2
18 11 7 11 11 13 2 11 11 2 1 11 11 11 1 9 11 12 2
6 9 9 11 10 9 2
29 1 9 12 2 9 11 2 12 2 13 9 11 1 11 11 1 11 11 11 2 11 11 11 11 11 11 11 2 2
29 11 11 3 3 13 3 13 3 3 3 11 11 7 13 13 10 9 1 9 1 9 9 0 15 3 3 15 9 2
25 3 2 9 15 13 11 2 11 2 9 0 15 13 13 9 2 13 9 1 9 9 9 15 13 2
6 10 0 9 13 9 2
5 9 9 13 11 2
40 1 9 9 9 9 3 0 13 1 9 9 1 12 9 2 9 9 12 9 9 9 12 9 9 9 12 9 9 12 9 2 9 12 9 7 0 1 12 9 2
10 7 3 11 11 15 3 13 9 11 2
61 1 9 12 11 12 11 11 11 11 13 9 0 15 13 1 11 11 2 11 2 16 15 13 1 11 11 11 12 0 11 11 11 1 11 11 11 2 9 10 13 1 13 11 11 12 2 9 0 11 2 1 9 1 11 2 1 9 12 2 12 2
45 9 9 0 0 2 13 2 0 3 2 3 13 1 9 2 0 7 13 2 12 2 12 5 9 12 2 12 2 12 5 2 1 9 2 9 15 13 13 9 2 13 1 12 9 2
19 9 13 2 9 10 9 13 1 11 11 7 1 9 12 13 9 12 9 2
13 3 3 13 9 2 13 9 7 9 2 9 0 2
22 11 2 11 11 13 10 9 1 9 7 9 1 11 11 16 11 11 11 11 11 11 2
15 10 13 9 10 13 0 2 3 13 1 12 9 15 13 2
11 13 13 11 11 12 2 12 2 12 2 2
26 9 13 1 11 11 2 9 10 3 13 1 11 11 11 2 11 2 2 16 9 13 9 1 11 12 2
38 9 9 1 9 10 3 13 9 15 3 0 7 3 13 9 15 0 2 0 0 2 16 1 12 12 9 3 13 1 9 12 1 9 12 9 9 0 2
38 16 9 0 11 13 1 9 0 11 2 7 16 11 13 9 9 11 11 3 10 9 1 11 2 3 11 3 13 2 13 1 9 11 7 11 1 9 2
54 1 15 13 15 13 1 11 11 15 13 2 11 11 11 11 2 2 11 11 1 9 7 3 11 11 11 2 11 2 11 11 9 2 11 2 3 13 11 2 11 1 12 9 1 9 7 9 15 13 1 9 9 11 2
38 1 9 15 13 1 9 11 2 15 13 13 16 1 13 9 7 9 15 13 1 0 7 0 1 13 9 2 9 9 2 9 15 13 1 11 3 13 2
21 11 9 1 9 13 12 2 12 9 9 9 1 9 2 0 12 2 12 1 9 2
28 1 13 1 11 2 11 11 2 12 9 10 13 15 3 0 2 1 9 9 9 2 1 1 9 9 9 9 2
26 11 2 9 15 13 9 10 13 16 11 11 3 13 15 13 1 9 15 14 0 1 9 2 9 0 2
15 9 9 13 10 9 9 15 13 1 9 1 9 1 9 2
14 9 9 11 3 13 1 12 11 12 1 12 11 12 2
47 9 9 9 7 3 3 13 1 9 9 0 13 9 1 9 15 3 0 7 0 2 15 3 13 1 9 1 9 2 16 3 3 1 9 12 5 12 12 5 1 9 7 1 9 9 9 2
18 13 9 1 12 9 1 13 10 9 15 13 1 9 10 1 9 0 2
23 11 11 1 9 10 0 13 1 10 9 15 9 10 13 11 1 1 9 9 11 7 11 2
14 16 1 11 2 11 13 1 9 7 9 11 7 11 2
28 1 9 10 9 15 0 7 13 3 13 7 9 13 1 9 9 11 1 9 9 0 2 9 3 13 0 3 2
19 9 11 11 13 0 1 9 9 9 15 13 9 7 1 1 9 9 9 2
135 11 11 11 11 2 11 2 1 11 11 11 11 11 11 2 11 2 1 11 11 2 11 11 7 11 11 11 11 11 11 2 11 2 1 11 11 11 11 11 11 2 11 2 1 11 11 2 11 11 2 11 11 2 11 11 11 11 11 2 11 11 11 2 1 11 11 11 11 11 2 11 5 11 2 11 11 2 1 11 11 11 11 11 11 2 11 11 2 1 11 11 11 11 11 11 2 11 11 2 1 11 11 2 11 11 7 11 11 2 11 11 11 11 2 11 11 2 1 11 11 11 11 11 11 2 11 2 11 11 2 1 11 11 11 11
16 16 3 2 9 3 13 1 9 7 9 9 11 13 0 9 2
22 3 3 10 9 15 13 3 3 0 1 0 3 13 9 1 13 9 9 9 15 13 2
12 2 11 2 13 13 0 2 11 1 9 10 2
13 11 13 10 11 1 1 9 11 2 11 2 11 2
14 15 13 9 10 1 2 11 11 2 2 9 9 2 2
16 11 11 11 2 9 0 11 11 12 1 11 2 13 1 1 2
26 9 11 11 11 2 2 13 10 9 1 11 15 13 9 9 12 12 2 7 9 12 9 2 12 2 2
6 3 11 13 1 9 2
11 9 10 0 13 1 9 1 0 2 0 2
25 11 11 11 11 11 2 11 11 11 11 11 11 11 2 13 9 11 9 12 15 13 1 11 11 2
16 16 9 1 9 2 11 13 13 1 11 11 2 9 11 11 2
4 3 9 13 2
15 15 13 1 9 1 9 12 11 12 1 13 9 1 9 2
11 9 11 13 1 9 10 9 1 9 9 2
20 11 11 1 9 13 1 13 3 1 9 12 2 10 2 7 3 13 1 9 2
25 9 9 3 13 12 0 2 9 1 9 11 2 9 10 13 10 9 1 13 9 7 9 0 15 2
6 9 9 9 0 10 2
15 3 12 9 12 9 2 2 2 2 2 2 2 2 2 2
78 9 15 13 14 13 1 12 9 1 10 9 15 13 9 9 2 11 2 7 9 15 3 13 1 9 9 11 2 16 9 1 9 11 9 0 2 1 13 9 2 9 9 1 9 9 11 2 9 15 13 1 9 1 11 2 11 2 11 7 9 0 15 13 9 9 3 13 1 11 11 15 9 3 13 1 11 11 2
10 11 10 13 9 15 3 13 1 11 2
27 9 9 13 13 12 9 9 9 15 13 1 11 7 11 1 9 11 11 11 2 9 11 13 9 9 0 2
18 11 11 15 13 9 13 0 3 13 9 2 16 9 11 11 3 0 2
26 9 0 3 13 3 10 9 15 13 1 9 2 9 1 13 3 13 1 9 9 16 9 10 14 13 2
70 11 11 13 3 9 9 2 1 11 13 11 15 13 9 9 11 1 3 1 9 9 1 9 1 11 9 1 11 2 11 11 3 13 1 13 10 9 15 13 9 9 2 1 9 15 0 2 11 1 11 11 2 9 9 9 1 13 11 2 9 9 1 11 11 2 7 9 9 9 2
36 3 1 0 13 9 2 9 15 13 1 3 7 9 9 9 15 13 1 9 2 7 13 10 12 9 1 9 9 2 15 0 9 1 9 9 2
32 15 13 1 11 13 9 9 11 11 11 2 7 13 9 11 12 1 11 15 13 1 13 1 9 9 13 9 15 13 9 11 2
17 9 10 12 13 1 9 12 11 12 7 13 1 9 12 11 12 2
21 11 2 11 11 13 9 15 0 7 0 1 13 9 3 15 13 1 10 11 11 2
26 11 3 13 2 14 2 16 9 2 9 15 0 13 1 13 7 3 13 16 15 9 11 2 7 11 2
34 15 13 9 10 9 3 2 13 1 9 9 9 0 2 9 9 2 2 16 15 13 9 11 2 15 9 10 13 9 9 1 9 9 2
14 7 9 15 3 13 1 11 7 11 1 13 9 15 2
8 3 9 9 9 11 7 11 2
10 11 2 11 3 3 0 1 13 9 2
39 1 13 2 13 1 9 9 2 16 9 3 2 3 13 9 2 7 9 2 16 11 13 10 9 15 13 11 2 2 11 13 13 3 0 1 9 9 11 2
15 1 9 0 13 9 3 3 2 3 3 3 13 9 0 2
24 11 13 9 2 9 1 9 1 1 11 7 11 13 1 13 11 2 11 13 3 1 9 9 2
27 1 0 13 2 11 11 2 2 11 13 1 11 7 11 1 10 9 9 1 13 9 11 15 3 1 11 2
25 3 3 2 3 13 3 12 9 0 1 9 15 0 2 3 11 11 11 2 11 7 11 11 11 2
40 11 11 2 2 13 0 9 1 11 11 11 15 13 9 13 9 7 13 1 9 9 7 9 9 2 9 10 3 13 9 1 13 9 1 9 1 13 9 0 2
27 7 3 13 1 11 2 15 3 13 9 1 9 0 2 16 3 2 3 3 15 13 9 9 1 13 9 2
18 11 2 9 10 1 0 13 15 13 9 2 9 2 9 2 7 9 2
17 9 11 13 11 2 11 13 1 9 0 1 9 1 12 9 9 2
21 9 15 14 13 1 9 11 2 16 15 3 13 11 1 9 1 10 9 1 11 2
15 11 9 1 11 11 13 11 11 11 11 11 1 9 0 2
33 11 11 14 13 16 12 9 3 2 9 10 13 7 13 16 15 13 9 11 11 11 1 9 9 9 9 2 7 1 9 10 9 2
8 11 11 13 9 1 12 9 2
27 9 11 11 2 3 13 1 1 1 11 11 7 9 13 11 11 11 3 13 1 9 9 9 11 11 11 2
5 15 9 11 11 2
17 3 13 9 9 0 1 11 15 15 13 16 1 9 10 13 9 2
11 0 9 9 10 2 3 11 13 13 9 2
20 16 11 13 1 12 9 9 1 11 11 12 2 11 13 12 5 1 9 10 2
19 1 9 10 14 11 0 15 13 15 1 13 9 2 9 2 1 9 15 2
15 7 9 2 9 13 13 1 15 7 13 9 0 1 0 2
16 1 9 11 11 15 13 13 1 13 11 3 1 11 11 11 2
23 13 1 9 12 2 9 0 1 9 9 9 13 13 9 9 1 11 0 16 13 11 11 2
20 11 13 1 11 1 11 11 2 11 2 10 9 11 1 9 9 10 2 12 2
23 1 12 9 3 1 11 7 11 2 15 13 11 7 11 1 9 12 2 12 1 9 13 2
5 15 15 13 9 2
22 11 3 13 0 2 0 1 10 9 1 9 9 9 2 9 2 1 9 9 13 0 2
25 11 11 11 13 9 10 10 9 15 13 1 9 11 11 11 2 11 11 2 11 11 11 2 11 2
7 11 13 9 9 1 11 2
16 1 9 2 11 13 9 1 11 11 11 7 13 9 9 9 2
15 9 15 3 3 13 13 1 12 2 12 9 1 9 0 2
15 16 9 9 3 13 13 9 2 7 9 9 13 9 11 2
8 11 2 11 11 11 2 11 11
9 11 3 13 1 11 2 11 11 2
13 11 11 2 3 15 13 1 11 11 13 1 9 2
17 11 13 9 15 13 1 11 11 2 11 11 2 11 11 2 11 2
18 11 9 9 11 2 11 13 9 9 9 15 13 11 11 7 11 11 2
6 11 13 9 1 15 2
25 3 1 9 12 2 11 13 13 9 11 7 3 13 9 3 12 9 2 12 9 3 13 9 0 2
23 11 11 13 10 9 11 13 9 12 15 13 1 11 11 7 13 1 11 11 7 11 11 2
23 13 1 9 12 2 11 3 13 1 2 11 11 11 2 16 13 10 9 15 13 9 10 2
20 12 11 13 9 12 2 12 2 9 12 2 12 1 9 0 2 1 11 11 2
29 9 9 9 9 9 1 13 9 1 9 9 13 1 9 2 9 1 9 13 9 9 2 16 9 10 13 9 13 2
7 9 9 11 13 12 9 2
11 15 3 3 13 9 2 16 0 1 13 2
18 1 9 9 9 10 13 3 0 13 1 9 1 9 9 7 9 0 2
7 3 11 11 13 7 13 2
20 9 10 13 9 1 11 11 11 2 11 7 11 11 2 1 11 2 11 12 2
26 3 9 13 0 2 15 13 13 9 2 9 9 2 15 13 9 2 7 9 9 2 15 13 9 9 2
92 9 0 2 1 9 9 7 9 9 0 2 13 10 9 9 2 15 3 13 1 13 2 9 0 2 9 2 9 7 13 9 0 7 13 0 2 15 3 13 1 9 0 1 9 9 2 9 9 0 1 9 9 0 7 9 0 13 1 10 9 2 16 13 1 9 9 2 9 9 0 2 1 13 9 0 15 0 3 13 1 9 2 9 2 7 9 2 9 2 10 9 2
14 16 15 3 13 16 11 14 3 13 1 9 1 10 2
27 10 9 9 10 3 13 11 2 16 15 3 13 1 13 9 15 1 11 7 11 15 13 2 12 9 2 2
11 3 9 14 13 9 11 2 11 5 9 2
189 9 9 11 2 11 11 3 1 9 12 2 15 3 9 1 11 2 11 2 11 2 15 3 13 1 11 11 11 12 11 2 7 1 9 12 3 13 9 9 11 12 1 13 11 2 11 9 13 11 2 11 2 11 2 1 9 12 13 9 9 11 12 1 13 9 2 9 2 11 11 11 9 12 2 12 2 1 9 12 13 9 9 11 12 1 13 11 2 11 2 11 2 11 2 11 1 9 12 2 12 2 1 9 12 13 9 9 11 11 12 1 13 11 2 11 2 11 9 9 12 2 12 2 1 9 12 13 9 9 11 11 12 1 13 11 2 11 2 11 11 11 2 11 2 11 9 9 12 2 12 2 1 9 12 13 9 9 11 12 1 13 11 2 11 11 9 9 12 2 12 2 1 9 12 13 9 9 11 12 1 13 11 2 11 11 11 1 12 2
34 11 5 11 11 11 11 2 11 5 11 11 2 11 5 11 11 11 11 2 11 5 11 2 11 5 11 2 11 2 11 5 11 11 2
11 9 9 15 0 13 7 13 13 11 11 2
18 11 13 9 15 13 1 11 11 11 2 11 11 11 2 11 2 11 2
26 11 11 13 9 2 11 11 2 1 9 9 9 2 7 13 9 2 11 11 2 9 0 1 11 11 2
21 9 10 13 10 10 9 15 0 1 11 7 13 1 9 9 15 13 11 11 11 2
20 11 11 2 9 11 2 2 11 11 2 11 11 2 7 11 11 2 11 2 2
12 9 9 1 9 10 1 9 12 3 12 9 2
12 11 13 9 3 2 3 13 11 13 1 11 2
42 9 9 11 2 0 9 10 1 0 9 0 2 3 9 13 9 0 7 0 9 9 2 11 2 15 13 1 13 9 7 3 13 13 9 15 0 1 9 2 0 9 2
18 11 13 9 1 11 11 11 11 2 2 11 2 2 2 2 11 2 2
12 11 13 11 16 9 15 13 1 11 9 12 2
12 9 15 3 11 13 1 13 10 9 0 11 2
15 13 9 11 1 9 0 15 13 9 1 13 9 9 10 2
10 15 3 13 9 15 13 1 9 0 2
17 1 10 9 0 3 13 1 9 13 9 11 2 3 11 2 11 2
11 1 11 2 15 13 10 9 1 9 11 2
15 11 10 3 13 2 7 3 15 13 1 9 1 9 9 2
4 3 13 9 2
14 9 9 1 9 13 12 2 12 2 2 12 2 9 2
9 13 11 11 2 9 9 13 15 2
9 11 13 9 1 11 2 11 2 2
18 7 10 2 12 12 9 0 13 3 7 9 2 9 15 0 2 0 2
21 9 9 9 1 9 0 3 3 0 16 13 1 9 15 13 1 10 9 3 3 2
9 15 15 13 1 9 10 13 9 2
31 9 9 9 10 16 9 1 10 9 1 10 9 15 13 9 15 0 13 1 10 9 15 9 0 7 3 3 3 14 13 2
34 11 11 2 2 11 11 2 2 13 9 9 9 15 13 1 11 15 13 1 9 11 11 2 1 10 10 9 9 13 1 9 15 0 2
15 1 9 0 2 9 2 9 0 11 13 9 13 9 9 2
22 13 11 11 3 13 9 11 7 13 9 11 11 11 11 2 16 1 0 15 3 13 2
25 9 10 3 13 1 9 12 2 12 1 11 2 11 5 11 2 7 3 13 1 13 10 9 9 2
14 13 3 3 1 13 1 9 7 9 13 10 9 13 2
9 11 11 13 9 1 13 10 9 2
14 11 13 10 9 1 11 11 2 11 11 11 2 11 2
11 1 9 13 12 9 0 9 9 1 9 2
9 1 9 2 15 13 0 1 11 2
14 16 13 9 9 13 9 2 16 9 12 1 1 9 2
16 9 10 13 1 13 9 11 1 12 1 12 9 13 9 12 2
15 1 9 12 11 13 1 11 2 1 9 3 13 3 9 2
18 11 11 3 13 9 1 9 11 2 15 3 13 1 9 1 11 12 2
68 11 2 9 15 13 11 1 9 15 0 13 16 1 9 0 9 1 11 11 2 11 13 9 1 9 2 11 3 13 9 1 0 16 9 1 11 13 9 11 2 16 15 3 0 2 7 11 3 13 16 13 11 13 9 1 9 0 2 16 9 15 1 9 0 13 11 11 2
5 2 13 9 15 2
41 13 1 9 12 11 12 2 1 11 2 11 2 9 9 11 11 2 11 13 10 9 1 9 12 12 9 2 1 9 11 11 2 11 2 15 3 13 1 12 9 2
17 9 0 10 3 0 1 13 1 9 2 16 3 13 9 0 2 2
35 1 10 9 15 13 11 3 13 9 1 11 2 16 15 13 9 2 9 9 15 13 1 9 9 12 2 7 10 9 1 13 9 1 11 2
9 9 1 11 11 14 3 1 9 2
28 3 13 1 9 10 9 9 1 10 9 0 1 12 9 7 9 0 3 13 10 9 3 9 9 9 0 0 2
84 3 3 1 9 9 9 12 1 1 9 12 9 10 3 13 9 0 1 11 11 7 9 15 13 1 9 0 7 13 1 9 0 15 13 1 9 11 11 13 1 9 11 13 1 11 11 7 11 11 15 13 1 9 11 1 13 1 11 11 15 13 11 11 1 9 9 10 2 10 9 2 2 11 11 11 13 3 13 9 1 11 11 2 2
14 9 9 0 15 13 9 3 13 9 1 13 9 9 2
23 11 13 1 10 9 15 13 9 2 9 9 2 2 7 9 0 15 13 1 9 7 9 2
21 9 9 9 10 13 9 15 13 1 9 9 9 7 9 9 10 15 13 9 0 2
22 11 13 10 10 9 1 11 11 11 2 11 11 11 2 11 2 11 11 11 2 11 2
20 3 11 3 3 13 11 9 15 13 16 9 2 11 2 3 13 16 11 2 2
16 1 10 9 7 9 2 3 11 3 13 7 9 11 3 13 2
14 11 13 13 10 9 15 13 9 1 13 7 13 15 2
17 11 13 9 15 13 1 11 2 7 3 14 13 1 9 9 9 2
22 11 11 1 0 1 9 9 9 9 0 2 9 2 9 11 2 7 9 0 1 9 2
42 9 0 2 13 7 9 13 2 13 9 0 2 1 9 12 2 12 2 12 2 12 5 2 9 12 5 2 13 13 12 2 12 2 9 13 9 2 7 9 0 0 2
52 1 11 11 2 9 11 11 13 1 9 9 2 16 1 11 11 2 9 11 11 13 1 9 1 11 2 1 9 10 3 3 13 9 1 2 3 12 9 1 9 15 0 1 1 11 11 13 12 1 15 0 2
16 11 13 1 9 0 9 2 13 1 9 9 16 13 1 9 2
33 11 2 3 13 1 11 1 9 0 2 13 9 9 15 13 1 11 11 7 0 1 9 0 2 3 1 9 2 9 7 9 9 2
24 13 11 1 9 2 9 9 9 13 1 9 9 9 0 2 13 9 0 2 0 2 13 9 2
26 16 2 3 11 11 3 13 9 9 0 1 12 9 9 2 16 9 9 9 1 9 10 3 0 3 2
21 9 10 13 1 12 7 13 3 1 12 2 3 9 0 15 13 11 11 11 13 2
23 9 10 2 3 13 1 9 9 9 11 2 9 10 3 13 1 9 9 9 1 9 0 2
9 7 9 15 13 1 2 9 2 2
20 11 13 2 9 11 2 2 11 11 2 2 7 9 2 9 13 2 9 2 2
12 9 9 13 1 9 15 13 9 16 13 9 2
17 11 13 1 9 10 2 9 9 15 15 13 16 3 13 9 0 2
19 11 11 13 9 9 11 11 2 9 11 11 2 9 11 2 7 9 11 2
24 1 12 9 10 13 1 1 12 9 9 1 11 15 0 3 13 11 11 1 13 1 12 9 2
18 9 10 13 1 9 9 7 9 9 9 1 11 11 15 13 1 13 2
37 1 9 2 15 13 9 1 13 9 11 15 13 7 13 12 12 11 2 1 11 2 13 12 11 11 2 11 15 13 9 10 13 7 13 1 11 2
5 9 9 13 9 2
17 11 9 0 1 11 13 10 9 9 15 13 1 11 13 9 12 2
18 11 11 11 11 2 11 2 1 0 13 9 9 1 9 0 9 9 2
18 10 9 9 9 15 3 13 1 11 11 2 0 1 11 11 11 2 2
14 1 9 10 2 11 13 15 3 13 1 9 9 0 2
45 11 13 9 1 9 11 7 3 13 1 10 9 1 11 11 2 11 11 11 7 9 9 2 1 0 9 12 2 11 13 1 11 11 1 9 9 11 7 13 9 13 11 5 11 2
18 9 3 13 2 13 2 13 2 7 13 9 7 9 1 12 0 0 2
18 11 13 9 9 1 9 11 3 13 9 9 1 9 10 1 9 12 2
22 10 11 11 13 1 9 0 15 13 9 9 9 0 7 9 9 2 1 11 11 11 2
25 11 3 13 9 1 13 9 15 0 2 15 3 13 9 0 7 0 1 9 1 12 2 12 12 2
34 9 15 13 9 12 10 13 1 9 12 11 2 16 13 9 2 12 11 10 3 13 9 9 9 1 9 13 9 0 9 11 7 11 2
17 16 2 9 13 13 9 0 7 13 9 2 9 10 1 9 15 2
11 11 13 10 9 11 15 13 1 9 12 2
17 11 11 11 12 13 11 11 11 12 2 12 2 15 13 1 11 2
23 1 9 11 12 2 11 13 12 9 1 11 1 9 9 3 1 12 2 12 9 1 11 2
13 11 11 11 2 2 2 13 9 9 9 1 11 2
44 1 9 9 11 10 11 3 13 13 9 11 9 11 2 16 11 11 2 11 2 11 11 10 13 1 11 11 1 9 12 2 10 2 7 9 11 13 9 9 1 9 9 11 2
22 1 9 9 9 10 13 1 9 9 15 3 13 1 13 11 11 1 9 11 11 11 2
9 9 9 11 11 13 9 0 11 2
54 1 13 9 9 9 9 15 13 2 11 13 9 0 15 13 9 1 11 11 2 11 9 7 9 10 0 2 3 1 13 11 15 13 1 9 2 9 13 7 9 2 9 13 9 1 9 11 2 11 7 11 5 11 2
13 11 2 11 2 11 13 10 9 0 1 9 11 2
28 9 10 13 9 15 0 1 9 9 7 9 9 11 2 3 9 9 9 15 13 7 9 7 13 13 1 9 2
22 11 3 3 13 9 1 2 3 13 9 9 2 11 3 0 1 9 2 9 9 9 2
29 10 9 10 13 13 9 9 7 14 3 13 2 10 9 15 0 3 3 13 1 10 9 7 13 1 9 15 13 2
6 7 1 9 15 13 2
24 11 11 2 11 2 12 11 11 2 13 9 9 11 11 11 11 15 13 1 11 11 2 11 2
28 16 9 11 7 11 1 9 0 2 0 1 11 11 15 13 1 11 1 3 13 7 13 1 3 1 12 9 2
13 16 3 13 9 0 9 11 1 13 9 11 10 2
9 3 9 9 9 9 14 13 9 2
15 11 11 13 10 9 1 11 11 2 11 11 11 2 11 2
21 11 11 11 9 10 3 13 11 11 2 16 11 11 13 9 1 9 1 11 11 2
24 9 10 11 12 2 13 2 11 12 2 2 13 9 9 9 11 11 1 11 11 1 11 11 2
18 11 9 10 13 12 9 2 3 11 11 2 11 11 2 7 11 11 2
22 1 9 9 11 12 2 11 11 11 11 13 9 1 9 11 11 7 11 1 9 11 2
34 1 9 12 2 11 11 11 13 9 9 15 13 1 9 9 2 9 0 7 0 7 9 2 9 15 13 1 9 13 7 13 9 9 2
19 16 9 1 11 2 9 11 2 15 0 13 1 13 9 1 9 12 11 2
55 1 9 12 2 12 11 13 1 11 11 11 11 11 2 3 1 9 12 2 12 15 13 1 9 11 11 11 11 7 3 13 11 11 11 11 11 2 12 2 12 2 7 9 9 9 9 7 11 11 2 12 2 12 2 2
90 1 13 9 9 7 9 0 2 1 9 2 12 5 9 5 11 5 12 5 12 9 12 11 12 2 11 13 9 9 13 11 11 11 2 11 2 1 11 11 12 2 1 9 9 2 12 5 11 2 12 5 11 2 12 5 12 15 13 1 11 2 11 2 11 11 2 9 2 2 1 9 12 11 12 2 11 11 12 13 7 13 9 2 11 2 1 11 11 11 2
22 1 9 12 11 13 1 11 1 10 9 7 9 15 3 14 13 0 16 9 10 13 2
19 1 9 10 10 9 1 13 3 13 13 1 13 9 7 13 9 10 9 2
29 1 9 2 9 13 13 9 15 3 15 13 1 10 1 9 2 9 11 2 9 11 2 9 9 7 0 2 0 2
18 11 11 11 1 9 11 13 1 2 10 9 9 2 2 16 9 0 2
23 3 1 9 2 11 7 11 3 13 10 9 2 7 3 9 2 13 9 15 0 1 15 2
25 11 11 11 13 9 9 9 11 2 11 2 11 2 11 15 13 9 9 15 13 1 11 7 11 2
13 16 9 13 2 9 9 9 12 3 13 1 11 2
7 3 15 13 13 9 15 2
18 11 0 13 2 11 11 2 13 9 12 2 12 5 1 1 9 9 2
12 9 7 9 13 9 0 1 9 9 11 9 2
15 11 3 13 9 9 9 9 15 0 1 9 0 1 0 2
10 16 11 13 2 15 15 3 13 9 2
66 11 13 9 2 9 1 9 9 11 11 11 11 11 11 15 13 1 11 11 2 9 11 11 7 9 9 9 11 11 1 11 15 13 1 11 1 12 11 2 7 9 2 9 9 9 2 12 11 11 1 11 11 0 12 11 9 9 11 11 11 15 13 1 11 11 2
22 1 9 1 11 11 2 11 13 9 2 9 2 12 9 9 2 9 2 9 7 9 2
14 11 13 9 1 11 11 2 11 2 11 11 2 11 2
20 3 3 15 3 1 9 0 16 13 2 10 9 11 13 15 13 1 1 11 2
16 9 10 13 9 9 9 15 13 11 12 9 1 9 12 13 2
28 1 11 12 2 15 13 1 13 1 11 11 11 11 2 15 13 9 1 11 11 1 9 12 11 12 1 11 2
17 3 11 9 13 9 1 9 11 7 10 9 15 13 1 11 11 2
25 11 3 13 10 9 1 9 9 2 1 1 12 11 11 2 12 11 11 2 12 11 11 2 11 2
12 11 13 10 9 1 11 2 9 9 1 11 2
28 1 9 9 10 2 9 10 9 0 7 9 15 13 9 9 13 1 9 13 13 9 11 11 9 12 11 12 2
18 11 13 10 9 9 1 9 11 2 11 11 2 11 11 11 2 11 2
17 9 9 9 7 15 3 3 13 1 9 9 13 9 10 2 9 2
31 1 12 13 12 9 9 2 10 9 0 2 2 7 3 1 12 11 12 2 16 11 11 13 1 11 11 2 13 9 11 2
25 1 9 2 11 11 13 1 9 11 11 11 2 11 15 0 13 1 9 7 13 3 13 1 9 2
41 16 13 9 9 0 2 9 9 2 2 9 11 11 13 1 10 9 11 15 13 1 11 11 2 11 11 2 7 11 11 11 2 11 11 2 7 13 1 11 11 2
16 9 0 9 11 11 11 13 1 9 0 2 12 2 12 2 2
38 11 13 9 0 1 11 11 1 9 12 11 12 2 15 13 9 12 1 11 1 11 11 2 13 1 11 1 12 2 12 2 12 2 12 9 11 2 2
15 11 11 2 11 1 9 9 0 11 13 9 1 9 11 2
16 9 9 9 7 9 15 0 13 1 10 9 9 1 9 9 2
17 11 11 11 11 11 11 13 10 9 15 13 1 9 9 15 0 2
9 1 9 11 11 15 13 1 11 2
10 9 15 0 10 13 1 11 11 11 2
51 11 10 13 2 11 1 11 2 7 15 15 13 9 10 9 1 9 1 11 2 1 11 2 11 2 11 11 2 2 9 2 9 2 9 7 3 13 1 9 9 1 11 2 9 2 7 9 16 1 11 2
23 1 13 10 9 15 0 1 11 11 11 2 11 13 1 11 11 11 11 15 12 2 12 2
20 11 3 3 13 11 11 11 2 2 11 2 2 15 13 9 9 1 9 0 2
6 10 9 13 10 9 2
32 10 9 3 13 10 9 1 9 9 0 7 0 1 9 9 9 0 2 16 15 13 9 13 0 7 0 1 9 9 9 0 2
25 9 0 9 9 9 9 15 13 1 11 2 13 11 12 7 11 12 2 13 9 1 13 9 9 2
35 9 15 3 0 1 9 11 13 1 0 15 13 1 12 9 1 11 7 11 11 2 9 12 2 11 7 11 11 2 9 12 2 12 2 2
18 1 9 9 11 9 2 2 9 2 13 1 9 9 15 0 7 0 2
23 15 3 13 11 11 2 1 13 9 9 10 2 11 13 9 0 15 13 1 3 13 9 2
39 15 3 3 14 3 13 9 9 9 2 15 3 13 9 2 9 0 1 13 9 2 1 9 9 0 1 9 2 9 10 2 9 9 2 7 9 9 9 2
18 11 3 0 1 11 11 11 13 2 11 11 11 11 2 1 9 12 2
16 1 9 0 2 9 10 3 13 9 7 9 7 16 13 9 2
35 10 9 16 9 12 9 2 15 13 1 9 9 2 11 11 2 15 13 12 9 15 13 1 13 9 15 3 12 9 9 9 9 3 13 2
7 11 15 0 15 3 13 2
32 11 13 9 15 13 1 13 9 7 9 9 1 10 9 1 10 9 0 2 9 1 9 9 2 9 2 9 9 2 7 9 2
25 11 11 2 2 13 9 11 11 11 11 11 2 5 5 8 2 8 2 8 2 8 2 11 2 2
21 11 13 9 9 9 11 13 1 10 9 0 11 11 2 1 1 9 1 9 13 2
15 11 13 1 13 9 9 15 13 7 15 14 0 1 9 2
17 9 13 9 11 11 11 11 1 9 9 11 15 10 3 13 3 2
37 9 9 9 9 15 13 1 9 2 9 2 9 9 2 9 9 0 2 9 9 9 2 9 2 9 2 7 9 9 0 9 13 12 2 12 9 2
8 3 11 13 0 9 13 15 2
18 15 13 13 9 9 1 11 2 1 13 9 9 9 1 9 9 9 2
59 13 9 9 15 3 13 11 11 11 2 11 2 3 3 13 10 9 9 15 13 9 9 2 9 2 9 9 2 9 7 9 9 15 0 0 2 3 10 9 9 9 2 13 11 11 2 15 13 10 9 9 1 9 9 9 2 11 2 2
19 3 3 3 13 9 9 1 13 9 9 2 9 0 2 7 9 1 13 2
11 15 3 13 9 11 1 11 11 2 11 2
9 16 9 14 9 15 0 1 13 9
48 11 11 1 11 13 9 15 0 1 10 9 13 2 16 15 3 13 9 0 1 13 1 11 7 9 1 2 11 2 9 9 0 2 11 11 7 11 2 9 11 2 13 9 0 1 9 10 2
13 11 15 13 1 11 13 9 15 0 1 11 11 2
28 9 9 13 16 9 13 9 0 0 1 9 9 0 2 15 13 1 9 15 14 9 0 1 9 0 15 0 2
24 1 13 13 2 11 13 9 11 11 11 1 11 1 11 11 1 9 11 11 1 13 1 11 2
8 13 9 15 13 9 1 11 2
22 9 2 9 0 9 11 13 3 0 0 1 9 9 2 9 2 7 0 1 10 9 2
35 16 3 0 16 15 0 13 9 1 11 13 11 11 1 9 9 12 2 16 3 1 9 12 9 13 9 2 9 0 1 11 11 11 10 2
23 9 3 13 1 9 1 9 0 2 9 0 2 7 9 9 1 9 2 9 2 9 2 2
13 11 13 10 9 1 11 11 2 11 11 2 11 2
32 3 2 1 3 13 2 11 11 13 1 9 9 2 13 9 15 13 13 11 2 7 9 13 13 9 13 11 1 10 9 9 2
16 11 11 11 2 2 13 10 9 2 9 2 7 9 9 11 2
19 11 13 9 9 1 9 12 2 1 9 11 2 11 2 11 11 2 11 2
3 9 9 2
17 3 13 1 11 11 7 11 11 3 13 1 11 11 1 9 12 2
23 9 9 13 1 12 9 2 16 2 1 9 0 9 13 1 10 9 0 15 13 1 9 2
32 11 13 10 11 11 1 13 11 11 2 11 13 1 11 11 11 1 9 13 2 11 11 11 2 13 1 9 1 9 9 9 2
19 11 13 9 9 1 9 11 11 11 2 11 11 2 11 11 11 2 11 2
13 9 3 13 9 9 9 15 0 1 13 7 13 2
10 9 10 13 9 9 9 2 12 11 2
78 9 9 11 11 13 1 9 9 1 9 9 0 2 9 11 2 11 2 11 2 11 2 11 2 11 11 2 11 7 11 2 10 9 9 0 1 11 11 11 7 10 1 11 11 14 3 13 9 9 1 11 7 11 2 16 3 13 1 2 11 2 2 7 9 15 1 2 11 2 2 9 11 11 1 11 11 11 2
10 11 13 9 2 1 9 3 13 9 2
22 1 9 9 2 15 3 13 10 1 9 1 13 9 1 9 15 13 1 11 11 15 2
20 16 11 13 11 11 11 2 12 2 12 2 2 9 11 3 13 9 9 11 2
27 11 11 11 11 2 11 2 13 10 9 0 15 13 1 11 11 2 11 11 2 1 12 9 9 1 11 2
15 11 9 11 2 15 13 11 2 13 9 0 1 9 10 2
21 14 3 10 3 2 11 3 13 1 11 11 11 2 0 1 9 2 7 13 0 2
14 9 10 13 0 1 9 11 11 1 11 11 11 11 2
18 1 9 12 2 15 13 1 11 11 11 11 11 2 11 2 1 9 2
24 11 13 10 10 9 1 11 2 13 1 11 11 2 9 10 3 13 1 10 9 1 9 10 2
24 11 13 9 0 15 13 12 11 12 2 13 12 1 12 9 7 13 11 2 11 11 11 2 2
34 16 9 3 0 7 9 9 9 9 3 0 1 13 7 13 9 2 16 9 15 13 13 1 9 1 9 9 13 9 15 0 7 0 2
48 11 13 1 0 11 7 1 1 9 1 11 11 2 9 11 11 10 13 11 2 11 9 3 2 3 9 11 1 9 9 1 9 7 13 2 9 1 11 13 9 9 15 3 0 16 11 11 2
13 9 13 12 9 10 13 13 1 9 12 11 12 2
32 11 11 11 7 9 9 11 11 11 11 11 13 10 9 9 9 9 15 13 1 11 2 11 9 2 12 2 11 11 2 11 2
64 11 11 3 13 1 9 12 7 13 9 0 15 13 1 11 1 9 9 1 9 5 12 9 2 9 0 7 0 2 10 9 13 1 9 1 9 1 9 2 16 9 3 13 0 1 9 16 13 1 9 9 9 1 12 9 2 16 15 13 13 9 3 3 2
34 1 9 11 2 10 0 9 11 1 11 11 11 7 13 11 13 13 1 11 11 1 9 9 9 11 2 15 13 1 9 9 11 11 2
26 9 9 1 11 2 11 2 7 11 2 11 7 10 9 15 3 13 1 0 1 11 2 13 7 13 2
14 9 9 9 13 2 13 13 1 9 9 9 15 13 2
14 11 13 9 1 11 11 2 11 11 2 11 2 11 2
20 9 9 9 7 9 15 13 1 11 1 3 0 13 9 9 9 9 10 1 9
13 11 11 11 11 2 2 2 2 13 10 9 11 2
6 11 11 3 3 0 2
23 1 9 2 9 9 2 9 9 2 7 3 9 13 1 9 9 9 15 13 1 9 9 2
25 9 10 13 9 1 12 2 12 12 1 9 9 13 1 9 7 13 9 9 15 9 13 12 12 2
13 11 11 11 13 10 10 9 1 11 11 2 11 2
28 1 9 12 11 11 3 13 9 9 9 9 2 1 9 9 9 3 0 1 9 9 9 9 0 10 2 11 2
5 9 15 3 13 2
13 11 13 9 1 11 11 1 13 9 1 9 9 2
8 16 15 3 13 13 10 9 2
10 3 3 2 11 3 13 1 11 11 2
6 1 1 9 13 0 2
19 13 15 13 1 9 15 13 9 16 9 13 13 9 7 3 13 9 9 2
23 9 10 3 3 13 1 10 9 9 1 9 2 9 0 1 11 2 1 9 13 7 13 2
5 9 13 11 11 2
9 11 2 11 2 15 15 13 15 2
46 16 9 0 13 1 9 9 11 2 9 10 13 9 1 0 1 9 11 1 9 11 1 9 12 11 2 7 3 13 1 9 1 9 11 1 9 1 9 11 11 15 13 1 9 12 2
20 1 13 1 11 12 1 1 9 12 2 11 13 1 11 2 9 9 11 11 2
14 10 13 13 9 0 9 12 1 9 9 10 1 11 2
121 1 9 9 13 1 13 9 2 16 3 2 9 2 0 13 9 2 1 9 0 15 13 2 9 2 2 9 10 13 9 9 15 0 2 0 2 3 1 9 9 1 13 9 9 2 2 9 11 11 11 11 11 11 11 11 11 2 11 11 2 2 2 9 1 2 9 2 3 13 1 10 9 1 13 9 7 9 2 1 2 9 2 7 2 11 2 1 7 1 9 11 2 2 9 2 1 1 9 11 2 7 2 9 2 1 1 9 11 2 1 9 11 2 1 9 11 2 1 9 11 2
22 11 11 2 1 1 10 9 0 1 1 2 13 10 9 9 1 9 2 9 2 9 2
5 3 15 13 9 2
15 3 13 1 11 7 11 2 3 13 1 11 1 9 12 2
19 9 3 2 13 12 9 9 9 2 16 9 0 2 0 0 2 7 0 2
26 16 9 9 2 7 13 13 9 1 9 2 11 11 11 3 13 13 9 2 7 13 9 0 1 11 2
13 15 13 1 9 16 9 13 11 1 9 13 11 2
17 11 13 12 9 1 11 11 11 1 9 12 1 9 1 9 9 2
10 16 15 14 0 1 2 16 9 3 2
23 3 15 13 9 0 15 13 2 0 2 7 9 9 1 9 0 2 7 16 15 13 9 2
15 1 9 2 9 9 10 13 10 9 9 15 3 13 13 2
5 15 15 13 0 2
13 16 11 13 2 11 13 1 9 7 3 13 11 2
10 13 10 9 1 9 11 11 1 11 2
55 9 10 9 2 9 9 13 11 2 11 2 11 2 3 13 0 1 9 7 9 15 0 1 2 11 2 2 9 14 3 1 9 7 9 2 16 3 3 9 2 9 9 2 13 1 9 9 2 9 2 9 7 0 9 2
6 9 10 13 9 9 12
12 3 2 9 9 11 11 13 1 9 11 11 2
55 16 1 9 9 2 9 9 15 3 13 2 9 13 9 9 2 9 2 1 2 11 11 2 11 11 11 11 2 11 11 2 11 11 2 11 11 2 11 11 11 2 11 11 2 11 11 11 11 2 11 11 9 11 11 2
14 3 9 9 9 1 10 9 15 13 9 9 12 9 2
5 9 9 11 10 2
36 11 3 13 3 9 11 1 13 13 11 11 1 13 11 2 15 3 13 1 11 11 11 2 16 13 16 11 3 13 1 9 10 1 13 9 2
48 9 2 9 9 7 9 2 1 15 14 13 1 9 9 2 16 13 1 9 1 9 0 2 3 9 0 2 9 7 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 7 9 2
20 1 9 9 9 10 13 11 11 2 1 13 11 15 13 1 9 9 9 10 2
39 11 11 12 11 7 13 3 1 9 11 13 10 9 11 1 11 1 11 15 13 1 11 2 9 2 11 11 2 11 11 11 2 11 11 11 2 11 11 2
14 1 9 0 1 9 10 2 11 13 9 11 15 13 2
17 11 11 13 9 15 13 9 2 13 0 2 7 13 1 9 13 2
8 15 13 1 9 12 11 12 2
19 9 15 13 9 1 9 10 13 11 11 2 15 13 9 1 12 1 12 2
16 1 9 12 2 9 10 13 9 1 12 9 7 12 9 9 2
9 10 9 11 13 9 1 9 15 2
15 1 9 9 12 2 9 11 13 3 13 1 9 9 9 2
31 1 9 9 15 13 1 9 1 11 2 11 1 9 12 1 12 1 13 13 9 2 11 2 9 1 9 15 1 9 12 2
5 11 11 2 11 2
13 16 13 13 0 2 15 3 13 9 2 3 11 2
27 11 13 9 1 2 9 9 2 2 16 3 15 14 13 9 1 9 2 9 3 2 15 3 0 15 0 2
16 9 2 11 2 13 1 9 11 11 2 15 13 2 9 2 2
32 15 13 13 1 9 2 9 1 11 11 9 1 9 10 9 9 14 0 2 1 13 9 2 11 5 11 11 2 1 9 12 2
14 13 3 9 2 9 15 0 1 9 9 10 3 13 2
34 1 16 10 2 16 13 9 9 15 13 1 9 9 3 1 9 15 0 2 3 3 3 13 9 1 9 9 9 15 0 1 3 13 2
35 11 14 13 0 1 13 9 9 2 16 1 9 0 1 11 12 10 2 12 2 12 2 2 11 0 13 11 12 7 13 3 12 9 3 2
24 1 10 2 11 3 3 13 9 9 2 9 1 12 9 7 13 9 9 0 1 12 12 9 2
7 9 15 13 1 9 15 2
19 9 9 15 13 9 15 3 0 1 9 11 13 9 9 2 9 7 9 2
45 9 10 13 12 9 2 11 11 1 11 2 11 2 11 11 1 11 11 7 11 11 1 9 2 9 2 7 9 15 13 1 9 9 1 11 11 3 0 1 11 11 1 11 11 2
11 11 1 9 12 2 13 9 1 12 9 2
16 11 13 10 9 1 9 11 11 2 11 11 2 11 11 11 2
33 11 13 1 9 1 10 9 9 0 10 7 1 1 9 9 1 15 13 1 9 2 1 9 9 2 7 7 9 9 13 10 9 2
33 9 10 13 9 1 9 11 3 13 2 11 11 11 13 7 13 11 7 11 11 15 13 1 9 2 11 11 1 9 13 1 11 2
19 16 1 9 9 9 2 9 13 10 2 10 9 15 13 1 13 0 9 2
39 9 12 9 15 3 13 9 9 9 2 11 11 2 2 16 10 9 9 10 15 3 3 13 1 10 9 11 2 7 14 13 3 10 9 1 11 7 11 2
11 11 7 11 13 11 16 11 13 15 10 2
22 1 12 11 12 2 13 9 9 1 11 11 15 13 9 10 1 11 11 11 10 11 2
25 9 2 11 3 13 1 11 2 15 11 2 2 15 13 9 9 0 9 11 11 11 1 9 10 2
23 16 10 9 11 13 9 10 1 11 2 16 11 13 2 2 11 0 1 9 13 13 9 2
26 1 9 12 2 11 11 11 2 9 10 9 1 9 9 2 13 9 15 13 9 9 9 16 9 13 2
20 3 2 9 13 1 9 2 9 9 2 9 0 15 13 1 0 2 7 9 2
19 10 9 9 3 3 13 9 15 0 2 9 9 2 1 13 9 15 0 2
40 1 9 9 2 9 10 13 9 0 2 11 11 2 2 9 9 13 2 11 11 5 10 2 9 9 10 15 13 15 9 2 2 2 1 9 15 3 0 13 2
70 16 7 2 11 11 15 13 1 9 13 0 11 2 9 9 13 11 11 2 9 11 2 11 11 11 2 7 11 13 9 11 11 2 11 11 2 11 2 7 10 0 9 11 12 1 11 2 9 9 11 13 1 9 11 15 13 9 1 11 11 2 16 9 3 13 1 1 9 11 2
8 11 11 13 0 1 12 9 2
71 11 3 13 9 0 2 16 2 3 13 2 2 9 9 9 2 9 1 9 9 15 13 2 9 9 7 9 9 2 9 1 9 9 15 13 1 9 9 13 9 9 9 0 1 1 9 9 15 3 2 9 11 2 7 11 11 2 10 13 7 11 13 9 2 9 0 1 9 9 2 2
12 1 9 0 2 11 13 9 11 7 11 2 2
35 11 13 11 1 9 12 11 12 1 9 12 9 7 12 2 12 12 9 9 11 2 7 10 0 9 11 11 11 9 10 13 1 9 9 2
18 3 9 9 13 2 12 2 10 9 9 13 9 12 9 1 9 0 2
15 11 1 0 13 13 11 1 11 1 9 3 12 9 3 2
34 1 11 12 2 11 11 11 11 11 7 11 11 11 11 11 13 9 0 1 13 9 0 1 9 9 9 11 7 11 11 11 11 11 2
29 9 10 13 9 1 11 11 11 11 2 11 2 11 11 2 11 10 13 10 9 1 11 2 11 2 1 9 12 2
24 9 11 2 11 11 11 1 11 11 11 2 11 11 7 11 11 11 2 2 13 16 10 9 2
14 11 13 9 1 11 11 2 11 2 11 11 2 11 2
25 11 11 2 11 2 11 2 2 13 10 9 9 9 13 11 11 15 13 1 9 11 1 9 9 2
10 9 13 12 5 2 9 1 12 9 2
10 1 9 11 11 2 11 13 9 13 2
12 11 11 2 2 13 9 9 11 11 9 11 2
24 1 9 10 9 11 2 12 13 1 13 9 1 9 0 2 7 9 1 13 9 1 9 9 2
25 11 2 11 11 11 9 1 9 2 9 15 13 9 0 11 11 10 13 10 9 9 9 2 9 2
19 3 11 11 1 12 2 9 10 13 9 0 11 11 2 16 9 3 0 2
17 11 3 13 15 1 9 0 7 3 3 13 1 13 1 1 9 2
20 16 3 13 9 0 2 9 2 7 9 9 15 0 2 9 3 13 11 11 2
16 11 2 13 2 2 13 9 9 15 3 13 9 1 11 11 2
62 15 3 13 1 9 1 11 11 11 11 2 9 1 9 12 2 12 13 9 1 9 0 2 1 9 15 0 2 11 1 11 2 13 10 9 2 13 16 9 0 11 2 1 9 12 11 2 2 11 2 13 0 1 9 9 11 11 2 15 13 2 2
46 9 9 1 9 0 13 9 15 13 3 2 3 10 2 13 1 9 12 1 11 11 2 15 3 13 11 11 7 11 2 9 15 13 9 1 9 7 9 0 1 13 9 1 10 9 2
20 1 9 2 9 10 3 13 1 9 15 13 9 2 3 13 9 9 9 2 2
10 10 9 15 0 13 1 10 9 10 2
16 11 2 11 13 10 9 1 11 11 11 2 11 11 2 11 2
11 11 13 1 13 11 2 3 15 13 11 2
34 1 9 12 9 2 9 10 13 16 2 11 11 13 9 9 1 9 13 1 15 13 1 14 13 0 1 9 2 9 1 9 7 9 2
18 15 13 9 0 1 15 11 2 7 15 15 1 9 0 3 13 11 2
37 1 9 13 9 7 9 9 9 10 2 10 9 3 13 1 9 9 10 7 3 13 9 15 13 7 13 0 1 9 9 15 13 2 11 11 2 2
15 9 9 9 1 9 11 11 3 13 1 13 1 9 10 2
28 1 9 0 1 9 11 11 11 2 9 7 9 1 9 7 9 3 13 9 7 13 3 9 1 0 9 9 2
7 9 12 9 1 9 9 2
17 15 13 9 15 3 0 9 15 3 15 13 2 1 10 2 2 2
5 0 9 9 15 2
14 16 9 0 2 11 11 2 11 2 13 10 9 11 2
8 3 15 13 3 7 13 15 2
11 11 13 9 15 13 1 11 11 2 11 2
35 11 9 1 9 11 13 9 2 1 13 2 2 16 10 9 2 9 13 9 2 15 3 13 10 9 1 9 7 15 13 9 1 9 13 2
14 11 3 13 1 9 9 2 0 2 0 2 0 2 2
35 1 10 9 11 1 9 9 11 1 11 2 11 11 2 9 2 9 9 11 15 13 3 12 9 9 2 12 9 9 2 7 12 9 9 2
34 1 9 9 11 11 2 11 11 11 13 1 11 1 11 11 12 2 13 9 9 10 15 13 3 9 11 2 1 9 9 12 1 12 2
30 3 10 9 15 3 3 15 13 2 1 9 15 0 7 9 9 2 15 0 1 12 2 12 9 1 2 11 3 13 2
14 11 2 11 2 13 9 9 9 0 7 9 1 12 2
11 16 10 3 15 3 15 13 1 9 10 2
45 11 1 9 11 11 7 11 11 11 1 13 9 1 13 10 9 0 7 13 0 1 11 2 13 1 13 9 2 9 9 2 9 2 9 9 2 9 9 7 9 2 9 9 0 2
13 11 13 3 13 1 13 9 9 1 0 16 13 2
13 11 13 1 9 12 15 13 11 1 9 11 11 2
17 11 11 11 13 9 0 0 1 11 7 13 9 0 12 1 11 2
24 9 9 15 0 1 9 13 9 1 11 11 3 13 2 3 0 2 7 3 13 1 9 11 2
4 3 9 13 2
23 16 9 9 13 1 13 13 10 9 0 15 3 13 3 9 11 11 11 15 13 1 12 2
11 11 2 9 0 3 3 13 9 9 0 2
24 11 13 10 10 9 9 9 15 9 2 9 1 9 0 3 13 1 13 9 0 7 10 9 2
22 11 11 13 10 10 9 15 13 1 11 11 11 2 11 11 11 2 11 11 2 11 2
29 11 3 13 9 16 9 11 3 13 1 9 2 16 14 13 9 3 13 1 9 15 0 16 9 11 13 1 9 2
10 9 2 11 11 2 3 3 3 13 2
24 11 10 13 9 15 13 1 9 0 7 13 1 9 9 1 13 9 0 1 9 2 9 0 2
16 11 13 10 9 1 9 11 11 2 11 11 2 11 11 11 2
37 16 2 1 0 9 15 13 9 10 16 13 16 9 3 0 7 3 13 1 9 11 11 2 1 9 15 0 15 13 11 11 2 10 9 1 11 2
24 11 0 9 10 13 9 11 15 0 7 9 1 9 3 13 3 13 9 10 3 0 1 11 2
21 9 13 1 13 9 9 15 0 2 16 9 13 1 13 9 13 9 16 13 9 2
16 11 9 3 13 9 9 3 3 1 12 2 12 2 12 9 2
11 9 3 15 13 9 9 9 7 9 10 2
12 11 11 1 9 12 2 13 9 1 12 9 2
16 9 9 13 3 1 9 10 9 2 13 1 9 9 9 0 2
139 1 10 2 11 2 11 3 13 13 9 1 13 9 9 9 7 11 2 1 9 9 1 11 7 11 2 9 11 11 11 11 11 2 16 11 15 13 10 11 1 9 9 3 13 9 9 9 2 11 11 11 2 1 9 1 13 9 9 9 2 9 9 2 7 9 9 9 2 11 2 9 0 2 15 13 1 11 2 11 13 9 9 9 2 9 9 11 12 2 9 11 0 9 2 7 9 9 9 2 1 10 9 0 1 2 9 12 9 9 2 9 11 12 2 9 9 12 2 9 9 12 2 7 10 9 0 15 13 2 13 1 10 9 9 1 9 11 11 2
14 1 12 9 0 2 11 11 13 9 1 9 9 9 2
16 11 2 2 2 13 9 15 13 1 11 11 2 11 2 11 2
12 9 2 9 10 1 9 13 13 12 11 12 2
9 15 13 1 9 9 1 9 12 2
28 11 2 9 9 2 9 15 13 9 0 1 9 2 13 9 0 1 9 9 0 7 0 15 13 11 11 0 2
26 16 1 0 13 2 11 11 3 13 9 0 0 1 13 9 9 9 0 1 9 9 9 1 11 11 2
14 3 3 11 11 13 9 13 11 9 11 1 9 0 2
34 1 13 1 9 2 9 9 0 15 13 13 9 13 12 5 12 2 7 9 9 12 12 15 13 13 9 3 13 12 5 12 2 9 2
6 11 0 13 11 11 2
15 11 13 9 1 9 11 11 2 11 11 2 11 2 11 2
100 1 9 12 11 12 3 13 11 11 7 1 11 11 11 13 12 9 11 11 11 11 15 13 1 9 12 11 12 1 13 9 9 0 16 11 11 1 9 2 11 11 7 11 11 11 1 9 9 7 1 9 12 11 12 15 0 3 13 13 9 11 11 11 11 0 1 9 9 9 12 2 12 1 9 11 11 11 9 2 12 5 12 5 11 5 12 1 9 9 9 11 11 11 11 9 9 12 2 12 2
8 1 12 10 9 15 3 0 2
83 9 11 11 7 13 1 11 11 11 13 9 12 9 13 1 12 9 7 12 9 2 11 11 13 12 5 12 12 2 12 5 12 12 9 9 7 12 5 12 12 2 12 5 12 12 9 9 1 9 0 2 0 1 9 9 9 12 2 12 9 9 9 9 13 9 9 9 11 11 15 13 1 9 13 9 9 9 1 9 9 7 9 2
17 14 3 10 2 3 3 9 0 15 14 13 1 9 11 1 11 2
16 1 9 12 2 10 2 10 11 7 10 11 13 0 1 11 2
13 11 11 2 2 13 10 9 7 9 9 9 11 2
11 9 13 1 13 12 9 13 11 7 11 2
23 2 11 11 11 2 13 9 1 9 9 0 11 15 14 13 2 2 9 1 10 9 2 2
11 11 10 2 11 13 13 9 12 9 9 2
20 11 13 10 10 9 15 13 1 9 11 11 2 11 11 2 11 11 2 11 2
17 15 13 9 9 1 9 9 15 3 13 12 9 12 1 9 10 2
29 9 3 3 0 13 1 9 10 2 9 7 9 9 15 13 1 9 10 13 9 0 13 9 15 13 1 9 0 2
31 11 2 11 11 13 16 9 2 11 2 11 11 2 13 1 9 0 15 13 9 15 3 13 9 15 13 9 1 10 9 2
20 11 11 10 13 11 11 12 1 9 9 9 3 13 9 1 13 1 9 9 2
41 11 11 11 11 2 2 13 9 9 9 9 9 11 2 11 3 13 1 9 0 1 11 11 2 11 11 2 11 11 2 11 11 2 11 11 11 2 7 11 11 11
33 11 11 11 2 15 13 1 9 0 11 2 3 0 1 11 11 1 9 12 2 10 16 15 1 9 11 7 11 3 13 1 9 2
34 15 13 9 13 0 9 10 14 3 9 9 2 7 3 7 0 9 15 13 9 7 9 9 7 9 11 3 13 9 7 9 11 11 2
32 11 10 13 1 9 9 7 13 9 12 2 1 13 9 12 5 2 9 12 5 7 9 12 5 1 9 0 13 1 9 9 2
9 15 13 3 3 13 12 0 0 2
28 11 13 9 15 14 13 1 11 11 16 11 13 9 2 11 11 11 2 16 9 15 13 1 11 14 13 12 2
27 1 1 11 2 9 11 13 10 9 0 1 1 11 2 11 2 11 2 11 2 7 9 0 1 11 11 2
12 11 7 11 13 9 1 11 11 12 11 11 2
20 11 11 13 10 12 9 1 9 11 15 13 9 0 1 12 11 1 11 11 2
11 9 9 15 13 1 9 9 3 13 9 2
22 14 3 9 14 2 1 1 9 13 9 11 15 13 0 2 13 1 9 15 3 13 2
15 9 1 9 9 9 9 9 15 13 0 1 9 9 9 2
13 1 10 9 10 13 10 10 9 1 11 1 11 2
26 10 9 15 13 1 11 11 11 11 1 11 11 12 13 9 9 7 9 9 2 9 13 9 9 0 2
10 11 11 3 13 9 9 3 2 3 2
26 9 10 14 13 0 2 16 3 13 3 1 9 9 3 2 3 2 3 13 7 9 0 2 0 2 2
19 15 13 16 3 13 9 1 11 1 11 11 11 2 7 1 9 11 11 2
9 9 9 9 13 12 2 2 12 2
23 3 10 9 13 1 9 11 11 2 15 13 0 7 13 12 9 2 12 0 7 12 0 2
38 16 0 13 2 11 11 12 11 2 15 13 1 11 11 2 11 11 2 11 2 13 9 13 12 11 3 9 11 11 2 11 11 2 7 11 11 11 2
15 11 11 2 7 13 11 11 2 2 13 9 9 1 11 2
22 11 11 7 3 13 1 11 11 2 2 13 9 9 9 7 9 7 9 9 1 9 2
14 9 3 3 13 2 16 11 11 0 9 1 12 9 2
18 16 9 9 7 9 13 1 9 0 2 16 9 15 3 1 9 0 2
20 9 13 11 11 11 10 13 9 10 9 9 1 11 11 2 11 2 7 11 2
27 1 9 2 9 15 0 2 9 9 13 9 9 3 2 9 2 2 9 9 2 2 16 3 13 9 9 2
33 11 9 11 11 12 13 12 11 12 1 9 12 2 12 9 0 2 12 11 12 1 9 12 2 12 11 2 0 11 11 2 11 2
45 9 9 11 11 11 1 11 2 11 11 11 2 11 11 2 11 11 2 7 11 11 13 11 11 11 1 13 9 2 13 9 9 15 3 0 2 7 9 9 7 9 15 3 9 2
40 9 10 13 9 0 11 11 11 11 12 5 11 11 11 11 11 11 5 11 11 11 15 13 1 9 9 7 13 1 9 11 15 13 2 9 1 9 12 2 2
18 9 9 13 1 11 11 11 3 13 1 9 2 9 15 13 9 9 2
13 11 11 11 3 13 0 2 16 9 11 3 13 2
17 11 11 13 12 9 15 13 1 9 9 11 11 1 9 13 9 2
13 11 11 13 10 9 11 11 15 13 1 9 12 2
51 16 10 2 11 15 13 3 2 3 1 9 11 2 2 13 12 9 9 11 12 1 9 12 1 9 9 9 2 9 11 2 11 13 9 2 9 11 13 1 9 7 13 11 1 13 9 9 1 9 10 2
19 15 13 10 9 0 2 11 11 2 11 2 7 12 9 13 11 7 11 2
20 11 11 9 11 2 11 7 11 11 2 13 9 9 9 9 9 0 1 11 2
6 11 10 13 9 12 2
31 1 9 12 11 12 9 9 12 1 9 9 11 2 11 2 11 13 1 9 9 1 11 7 9 9 9 9 1 11 11 2
16 13 9 16 15 3 13 1 1 9 2 11 3 3 12 9 2
23 11 13 10 10 9 1 9 11 11 11 11 2 11 11 11 11 2 11 11 11 2 11 2
164 1 13 9 9 10 11 9 11 11 11 11 11 11 11 13 13 9 9 9 11 7 13 9 0 0 1 9 9 2 15 13 13 1 9 1 11 11 11 11 2 11 10 13 1 7 13 9 0 1 9 11 11 11 2 9 7 9 9 11 11 11 11 11 11 11 11 11 2 16 13 1 9 11 11 11 11 11 2 9 12 9 12 3 2 11 2 16 1 13 7 13 9 11 15 3 13 1 11 11 11 11 2 3 13 11 11 11 11 11 11 11 11 11 2 11 2 16 1 11 11 11 11 11 11 11 11 11 3 13 9 1 13 9 7 13 13 3 1 13 9 11 7 11 11 11 9 11 11 11 11 11 11 11 2 12 2 9 2 11 11 2 7 9 2
19 11 12 10 13 1 12 9 12 2 1 1 11 12 2 12 11 3 13 2
27 1 9 0 12 2 15 13 1 11 11 2 16 1 12 11 12 15 13 1 11 11 1 9 9 12 9 2
29 1 11 9 15 13 9 9 9 0 1 0 10 3 13 12 9 9 2 12 13 9 5 12 5 12 5 2 9 2
15 1 11 2 11 13 1 11 7 3 13 11 2 11 11 2
5 9 10 9 0 2
21 11 13 9 11 11 11 2 9 2 11 11 15 0 2 7 11 11 11 11 11 2
22 11 11 11 5 11 2 11 2 13 12 12 2 12 5 2 9 11 2 11 2 11 2
16 16 3 0 0 2 9 11 7 11 13 1 13 3 12 9 2
46 11 9 0 11 15 13 1 11 2 9 7 9 2 13 9 11 1 11 15 13 12 9 11 11 0 1 9 11 7 9 11 2 11 7 11 13 9 1 1 11 1 9 9 9 11 2
7 9 3 11 2 3 14 2
18 11 15 13 9 0 1 13 9 0 11 10 13 13 9 9 9 0 2
20 3 11 7 9 3 13 9 15 3 13 7 3 0 3 13 9 1 9 15 2
11 9 10 9 11 7 3 9 0 11 11 2
25 11 11 2 11 2 11 11 2 13 9 15 13 1 1 9 11 2 9 13 12 9 2 12 2 2
3 0 3 2
38 11 9 5 9 3 13 9 1 9 2 9 9 7 3 10 9 13 16 0 9 13 10 9 9 9 2 1 0 9 9 2 9 2 7 9 7 9 2
34 16 3 15 13 13 9 11 2 12 9 13 9 15 1 1 9 11 11 2 15 3 15 13 1 9 9 11 1 9 9 2 13 9 2
7 15 13 1 11 11 11 2
23 11 11 11 13 9 1 1 11 11 2 11 11 7 10 11 11 7 11 11 1 11 11 2
19 11 11 11 13 1 0 11 2 11 11 11 2 11 2 1 12 11 12 2
32 1 9 15 0 15 3 13 11 11 7 1 9 12 13 9 9 11 15 13 1 9 10 3 3 1 11 11 11 2 11 2 2
19 11 11 12 13 16 11 5 11 3 13 9 10 9 1 11 11 11 11 2
37 16 9 9 13 9 9 15 3 3 2 16 9 3 13 1 9 12 15 13 1 10 9 9 9 7 9 1 9 9 15 0 7 9 9 15 13 2
15 9 11 3 13 9 13 9 16 13 7 3 13 9 0 2
15 11 3 13 10 9 2 13 9 1 11 11 1 11 11 2
15 11 11 13 10 9 9 9 9 7 9 11 2 11 11 2
21 11 12 9 0 13 11 3 1 9 1 9 0 1 0 2 0 9 9 9 9 2
20 11 11 3 3 3 0 13 1 11 7 9 9 9 10 13 9 9 1 1 2
18 11 13 9 1 9 2 0 9 9 2 0 9 2 7 9 0 9 2
23 2 11 11 11 2 13 9 1 13 9 9 15 13 1 11 7 11 2 9 1 11 2 2
21 11 11 12 2 9 13 9 9 2 10 2 9 13 1 11 11 11 2 11 2 2
16 15 1 9 9 2 3 15 3 13 1 9 15 0 1 10 2
33 11 13 9 15 13 1 11 11 15 13 1 11 11 2 9 9 7 9 15 13 9 10 1 1 9 12 9 1 9 12 2 12 2
25 9 13 10 9 9 0 13 11 11 2 15 3 3 13 1 11 2 11 9 13 1 11 1 9 2
34 9 2 9 2 3 13 1 9 15 13 1 9 2 9 2 9 7 9 9 0 15 13 2 9 2 9 11 2 11 2 9 7 11 2
19 1 9 10 3 13 13 13 10 9 13 11 2 16 9 1 11 14 13 2
11 3 2 3 13 11 11 1 11 11 11 2
14 11 13 9 1 11 11 2 11 2 11 11 2 11 2
30 11 10 13 9 15 3 0 2 9 9 11 2 2 16 9 10 1 11 11 3 1 9 9 9 2 9 9 0 2 2
6 10 0 9 13 9 2
37 1 9 12 11 12 2 1 9 9 9 1 11 11 2 11 13 1 9 9 12 2 16 13 1 9 1 12 9 9 1 11 11 13 12 2 12 2
11 9 10 13 9 1 0 9 9 11 11 2
15 11 3 13 9 1 13 1 11 11 11 11 1 9 12 2
25 9 10 13 9 9 9 0 1 9 11 7 9 11 15 13 1 9 11 2 11 2 11 2 11 2
20 11 13 10 10 9 1 9 9 11 2 9 11 11 2 9 11 11 2 11 2
24 1 9 11 11 11 2 11 11 2 13 2 16 11 13 10 9 15 0 1 13 1 9 9 2
15 7 14 13 9 11 11 15 13 11 1 11 1 9 12 2
59 9 10 11 11 11 11 3 13 9 15 13 11 1 9 9 11 2 1 13 9 9 7 13 9 9 9 11 11 11 11 2 16 13 9 9 11 11 7 15 3 13 1 11 2 9 9 11 11 11 11 11 13 1 12 2 12 2 9 2
38 9 2 9 9 9 9 10 1 1 2 7 7 2 11 13 9 9 15 0 7 0 2 0 2 1 9 0 2 13 1 9 2 9 9 7 9 0 2
10 9 9 9 1 9 13 9 1 9 2
18 9 15 0 1 9 9 1 9 9 0 13 1 9 9 9 9 0 2
12 9 9 15 3 13 1 9 1 12 9 10 2
16 11 7 13 10 2 10 9 15 13 1 9 11 2 1 9 2
20 9 10 13 1 11 11 7 9 10 2 16 0 1 13 9 1 9 0 10 2
20 1 12 2 11 13 1 11 11 15 9 0 11 2 7 13 0 1 9 9 2
13 1 9 9 11 13 13 2 11 11 3 3 13 2
43 1 9 2 1 9 9 11 9 3 13 13 11 11 2 11 11 11 2 2 1 9 9 11 2 11 11 2 11 11 2 2 9 9 11 2 7 11 11 2 11 11 2 2
12 11 11 11 11 12 2 11 11 11 2 11 2
17 11 13 9 15 13 1 11 11 2 11 11 2 11 11 2 11 2
13 2 7 15 15 13 13 3 1 10 9 11 11 2
9 11 2 9 9 13 1 9 9 2
120 1 10 9 2 9 13 11 11 2 11 2 12 2 2 11 11 9 1 9 9 1 11 11 11 11 2 11 2 11 9 11 11 11 11 11 11 2 9 11 11 2 11 2 12 2 2 9 9 9 11 11 2 11 11 2 11 2 12 2 2 11 11 11 12 2 9 1 9 9 1 11 11 11 11 9 11 11 2 11 2 12 2 2 11 11 11 11 11 12 2 12 2 11 2 12 2 2 9 9 11 2 11 2 12 2 2 9 9 11 2 11 7 11 11 2 11 2 12 2 2
52 9 7 9 13 10 9 15 13 1 11 11 11 1 13 9 9 3 2 3 10 9 0 15 3 0 7 3 13 15 13 10 9 0 15 0 2 11 2 13 9 2 9 7 9 2 9 15 13 1 9 9 2
24 9 1 9 9 1 9 11 11 7 9 2 13 10 10 9 1 11 7 9 15 14 13 9 2
22 10 15 9 14 9 9 9 2 13 3 9 2 9 9 2 16 3 9 9 16 9 2
23 11 2 9 9 2 9 14 3 13 1 7 13 12 0 0 16 15 13 1 9 9 0 2
6 3 11 3 13 11 2
20 16 9 13 2 11 11 0 13 9 11 11 2 9 10 15 3 13 12 9 2
51 2 15 14 13 9 2 16 9 9 2 9 11 3 1 9 2 9 0 15 2 2 13 11 2 9 3 2 11 13 1 11 11 2 1 9 9 0 11 11 11 11 11 11 8 2 11 2 1 11 11 2
9 16 3 9 0 13 1 9 11 2
18 11 9 0 13 1 12 7 12 2 9 2 9 1 11 11 7 11 2
12 9 10 13 1 9 9 9 9 7 9 9 2
8 10 9 3 3 13 9 10 2
35 11 14 13 9 11 11 1 10 9 0 2 9 11 13 9 10 1 9 0 2 11 2 7 3 2 9 11 2 13 9 9 9 10 2 2
20 11 13 1 9 0 2 1 9 12 9 13 1 9 2 9 15 13 9 11 2
9 14 15 0 2 2 3 15 0 2
22 3 1 13 11 11 11 2 11 2 1 9 16 9 9 13 0 1 9 9 7 9 2
14 11 13 16 14 13 9 1 9 15 13 9 9 9 2
21 12 9 13 1 10 9 15 13 9 3 13 7 14 3 13 2 7 1 9 9 2
4 15 15 9 2
9 1 11 2 11 13 9 9 11 2
32 16 3 1 11 2 11 13 1 9 7 3 0 1 9 11 11 7 11 11 2 11 15 0 13 3 1 11 15 13 1 11 2
15 9 11 10 13 9 1 9 9 11 11 11 2 11 11 2
30 11 13 9 1 9 9 9 10 0 7 3 13 9 9 2 9 7 9 9 15 13 1 13 9 9 7 13 1 9 2
34 15 13 9 0 12 1 9 11 11 9 12 1 2 1 12 11 12 9 9 11 11 13 1 9 1 9 2 16 11 13 9 0 0 2
24 9 9 10 13 1 9 15 13 1 9 9 2 11 2 2 9 9 15 13 0 1 9 9 2
11 11 13 1 11 1 11 1 13 9 9 2
15 1 9 12 9 2 15 3 13 11 11 11 12 1 11 2
21 11 13 1 9 15 13 9 9 10 9 9 0 1 11 11 1 9 2 11 11 2
18 11 13 9 15 13 1 11 11 11 2 11 11 2 11 11 2 11 2
33 1 9 2 15 13 3 9 13 1 10 9 11 2 15 3 0 1 9 15 13 11 11 2 11 2 15 3 13 9 1 11 11 2
33 11 11 2 11 2 9 9 9 11 2 15 9 13 9 9 7 9 9 11 11 2 13 1 9 9 7 7 11 11 1 11 12 2
16 13 1 9 9 11 2 9 10 9 1 13 1 11 11 13 2
12 1 9 10 3 13 9 2 9 15 3 13 2
23 9 12 5 9 1 9 9 13 1 9 0 2 1 9 9 2 9 0 2 7 9 0 2
19 11 11 2 13 12 11 12 2 13 10 9 13 11 15 13 12 11 11 2
31 13 1 11 2 11 7 11 2 11 11 2 15 13 9 9 1 11 2 7 3 1 11 2 7 16 15 13 10 9 9 2
5 15 13 1 11 2
35 1 9 2 9 10 0 16 9 9 2 9 7 9 9 2 3 13 0 1 9 9 0 7 3 13 1 9 9 1 9 0 15 3 13 2
10 9 10 3 13 9 15 13 2 3 2
18 11 11 2 2 13 9 9 11 11 11 9 12 13 1 11 11 11 2
24 10 9 13 9 10 1 10 9 0 2 16 13 1 10 9 15 3 3 13 9 2 9 0 2
14 16 2 15 3 9 9 9 0 1 11 11 11 11 2
5 15 9 13 0 2
8 11 0 10 3 13 9 9 2
27 11 13 9 9 1 9 11 2 11 11 2 11 7 11 2 11 16 13 9 9 1 9 10 1 9 12 2
5 3 15 13 3 2
15 11 11 13 9 1 9 11 2 11 2 11 11 2 11 2
14 16 9 11 1 9 12 13 11 2 11 11 13 9 2
27 11 9 3 13 11 11 2 15 0 7 13 2 13 0 9 2 7 11 11 13 7 3 13 13 11 11 2
12 9 15 3 13 11 16 13 11 7 11 0 2
11 11 11 11 2 11 13 9 1 12 9 2
32 9 11 9 10 13 1 13 9 15 13 1 9 2 16 7 1 9 9 11 3 3 9 15 13 2 13 10 9 15 13 9 2
17 11 13 9 15 13 1 9 11 2 11 11 2 11 11 2 11 2
37 9 15 3 13 1 9 9 9 1 9 12 12 2 15 3 3 13 9 2 13 13 1 13 10 11 11 11 1 9 1 9 12 1 11 2 11 2
21 9 10 15 13 1 11 7 3 13 1 9 9 9 2 9 9 2 7 9 9 2
11 9 11 15 3 0 13 9 7 9 0 2
31 1 9 13 12 5 11 2 12 5 12 9 12 11 12 1 9 9 9 2 11 11 11 11 13 16 9 9 13 1 11 2
13 11 9 13 9 15 0 7 0 1 12 11 12 2
12 1 9 10 2 9 3 13 9 9 1 11 2
18 11 13 9 9 11 11 11 9 9 11 11 11 2 13 1 9 12 2
8 16 12 9 11 13 1 9 2
14 1 9 12 15 13 1 11 11 11 1 11 11 11 2
23 10 9 15 3 13 13 13 9 1 13 9 7 10 0 13 9 0 1 10 0 9 11 2
30 11 11 11 2 13 1 9 9 0 7 9 11 11 2 3 9 0 2 2 11 2 11 11 2 11 11 7 11 11 2
26 1 9 2 9 2 9 0 1 13 9 9 0 2 0 1 11 13 1 3 3 13 1 9 1 11 2
7 3 15 13 9 12 5 2
18 9 9 9 10 14 13 1 9 1 9 9 9 10 13 1 9 9 2
17 3 2 9 3 1 13 9 7 9 15 13 1 13 10 9 0 2
20 15 3 13 9 2 11 11 2 7 9 3 13 12 9 3 0 13 9 9 2
13 2 11 11 11 2 9 9 15 13 0 1 15 2
57 1 11 11 11 2 11 2 9 10 2 15 15 13 1 9 9 2 9 2 13 9 15 0 2 15 13 13 9 9 2 9 11 2 11 2 11 1 10 9 1 13 9 9 11 2 11 2 11 1 9 1 11 2 11 2 11 2
16 1 9 10 2 1 9 11 13 12 9 15 3 13 7 13 2
27 11 15 13 1 9 10 14 3 13 3 16 3 13 9 2 9 9 2 15 1 9 13 3 13 9 2 2
14 1 0 9 10 2 12 2 11 3 13 13 12 9 2
24 1 9 0 2 11 7 9 2 11 2 13 1 11 16 13 1 9 2 11 2 1 13 9 2
31 10 2 10 3 13 1 9 15 13 1 11 11 11 1 11 11 1 9 11 9 11 2 11 11 9 11 2 11 2 11 2
16 1 11 2 11 13 9 15 0 7 3 13 9 15 3 0 2
19 11 13 12 2 12 9 1 11 11 15 10 9 13 1 9 11 11 11 2
12 16 11 1 9 15 2 15 15 3 13 15 2
7 2 3 14 11 11 11 2
19 1 9 12 2 12 2 11 9 10 13 1 13 9 9 1 13 9 9 2
18 9 10 13 9 9 2 7 9 9 9 1 13 1 9 1 9 9 2
26 9 15 13 1 10 9 9 11 11 13 9 1 9 1 9 2 15 1 10 9 13 16 9 1 9 2
41 11 11 11 11 2 2 13 9 0 11 2 9 1 9 11 11 2 11 11 11 11 13 1 12 9 2 1 9 12 2 12 7 12 3 13 1 9 11 7 11 2
17 11 11 13 16 11 13 9 9 9 15 14 13 1 1 9 9 2
10 11 11 11 11 13 1 9 11 11 2
22 1 9 13 9 2 9 13 13 12 9 2 1 11 7 11 3 10 9 0 1 11 2
23 15 13 9 2 9 9 7 13 1 9 0 9 3 9 9 7 9 9 9 2 9 2 2
22 11 11 13 10 10 9 15 13 1 9 11 11 2 11 9 11 2 11 11 2 11 2
6 9 11 3 13 13 2
6 1 9 3 15 13 2
14 11 13 9 1 9 11 2 11 2 11 11 2 11 2
5 3 10 3 13 2
10 9 10 2 9 9 11 13 9 11 2
13 1 9 12 11 11 13 0 7 13 1 9 0 2
17 11 2 9 15 3 13 11 3 13 7 13 0 1 9 11 13 2
16 1 9 10 15 13 1 9 11 11 12 2 15 13 1 9 2
7 2 3 15 13 9 11 2
10 16 3 2 9 10 3 13 9 3 2
30 11 15 14 13 9 2 9 10 13 11 1 12 9 2 9 9 15 3 13 1 9 9 3 13 1 0 16 13 11 2
16 9 10 13 1 9 9 9 9 9 9 12 1 5 1 12 2
21 11 11 13 9 9 0 2 13 9 9 9 11 11 11 11 7 9 9 11 11 2
17 12 2 11 11 11 7 11 11 11 2 13 9 9 13 10 9 2
24 14 11 11 3 13 10 9 0 2 16 15 13 11 10 2 9 9 9 0 7 13 15 13 2
21 11 0 11 13 2 13 1 10 10 9 9 9 15 13 1 9 9 1 9 0 2
19 11 3 13 13 9 1 9 7 9 1 9 1 9 7 10 9 1 9 2
34 10 0 9 11 11 3 15 15 3 1 11 11 11 9 9 2 11 2 1 9 2 9 9 3 11 2 9 13 9 15 13 1 9 2
8 13 11 13 9 9 1 11 2
4 1 1 11 2
30 1 9 12 11 13 9 9 11 2 11 11 7 3 13 9 9 2 9 9 9 2 9 7 9 2 1 9 11 11 2
10 1 13 9 3 13 9 7 3 9 2
15 11 3 13 1 9 9 11 2 11 11 0 11 2 11 2
63 11 11 11 11 2 7 11 11 11 2 11 2 13 9 0 11 11 11 15 13 1 9 12 2 15 13 9 7 9 1 11 11 2 11 11 13 10 9 1 10 9 0 15 13 1 9 0 2 9 7 9 9 15 13 9 1 11 7 9 2 9 9 2
22 11 11 2 13 11 11 11 12 2 2 13 10 9 2 9 9 11 11 1 11 11 2
16 1 12 2 9 11 11 11 13 9 11 12 15 13 9 9 2
12 10 9 2 9 14 3 13 0 1 9 9 2
14 11 11 11 3 13 9 15 3 0 1 10 9 9 2
14 11 13 9 1 11 11 2 11 2 11 11 2 11 2
17 11 13 10 10 9 1 9 11 2 9 11 2 11 11 2 11 2
12 11 11 7 11 11 13 9 0 1 9 11 2
33 11 11 13 0 1 11 11 11 11 2 11 2 2 11 11 11 3 13 13 1 11 2 11 11 2 7 11 2 11 11 11 2 2
8 11 10 13 1 11 2 11 2
10 14 1 9 0 2 9 10 14 13 2
8 9 10 13 1 9 10 9 2
14 11 2 9 13 9 15 13 11 13 11 11 11 0 2
3 2 7 2
23 1 13 9 0 15 9 11 0 7 13 11 11 2 11 13 1 10 9 11 13 11 11 2
8 9 13 13 12 12 2 12 2
31 13 1 9 9 11 2 11 11 11 13 15 1 11 2 11 12 12 2 9 0 2 0 9 2 9 9 1 9 11 11 2
12 1 9 12 2 9 10 13 9 1 12 9 2
40 9 9 0 13 10 9 15 3 13 13 9 9 15 3 0 7 0 1 9 0 7 9 9 13 9 9 9 2 3 13 3 0 1 12 5 2 12 12 2 2
33 16 13 1 11 2 11 11 11 11 1 12 11 12 13 1 11 11 2 16 9 9 11 15 13 1 9 11 2 3 13 1 11 2
7 2 3 9 13 9 10 2
31 11 2 9 9 9 1 0 1 9 9 2 9 15 0 2 9 9 15 13 9 2 9 12 7 9 3 2 3 9 0 2
33 11 13 13 9 10 1 11 2 12 11 12 2 7 11 1 9 12 11 12 2 9 1 9 12 2 12 11 2 11 5 12 2 2
28 16 15 3 13 1 9 12 2 7 15 14 13 10 9 1 9 2 11 2 2 15 1 9 0 13 9 12 2
63 11 11 2 12 2 7 3 13 11 11 2 13 10 9 9 9 0 2 13 0 15 13 1 9 9 11 11 7 3 13 3 1 11 2 11 10 3 13 9 9 1 9 0 2 12 9 2 3 12 9 2 1 9 0 7 0 2 7 1 10 9 9 2
27 11 13 9 3 13 13 11 9 9 9 9 11 11 2 11 11 2 1 9 11 11 11 5 11 9 12 2
50 1 9 12 3 13 9 12 2 12 12 12 2 9 2 16 1 9 10 9 9 9 11 11 11 13 1 12 2 12 12 2 9 2 12 2 12 12 2 9 7 12 2 12 12 12 12 12 2 9 2
9 3 13 9 1 9 15 3 0 2
21 11 11 13 3 13 9 15 0 1 9 9 12 11 2 15 13 1 12 11 12 2
7 9 0 7 9 9 9 2
24 11 11 15 13 0 1 9 9 15 13 13 9 10 1 9 0 13 7 13 10 9 10 9 2
34 1 9 2 9 0 15 13 1 1 9 2 1 9 10 11 2 13 3 2 3 12 9 9 2 2 12 2 0 1 13 9 1 9 2
31 12 9 10 13 11 11 2 0 2 2 11 2 11 2 11 2 11 2 11 2 11 11 2 11 11 2 7 11 2 11 2
21 11 9 13 10 9 1 11 11 11 2 11 11 11 2 11 11 11 11 2 11 2
14 16 15 13 9 0 13 2 3 11 13 1 9 9 2
17 15 3 15 3 13 11 1 11 11 2 11 11 2 7 11 11 2
9 1 9 10 13 11 2 11 2 2
29 1 9 11 11 2 12 2 7 11 2 12 2 2 11 13 9 13 11 2 7 13 11 11 11 1 11 11 11 2
9 9 13 9 11 7 9 9 11 2
6 9 13 3 13 9 2
14 1 9 2 9 1 9 10 3 13 9 10 1 15 2
17 11 13 16 9 2 3 9 2 9 2 13 1 9 2 9 9 2
11 1 9 2 11 11 11 13 9 9 9 2
23 9 10 9 9 0 3 13 1 9 11 2 11 2 7 11 2 16 9 3 13 1 9 2
59 9 1 11 2 9 7 11 13 1 1 9 9 2 11 2 12 2 2 16 9 9 15 13 1 11 1 9 12 13 1 11 2 11 7 11 2 11 9 13 3 1 9 0 2 16 3 3 13 1 9 9 1 12 12 1 1 9 9 2
22 11 2 11 11 2 2 11 2 11 11 2 7 11 2 11 11 2 3 13 1 0 2
14 11 11 11 11 13 3 13 1 9 10 9 11 11 2
24 2 1 9 15 13 13 7 3 13 1 9 15 0 7 2 13 2 14 13 9 9 1 13 2
8 11 0 13 1 9 11 11 2
7 3 16 9 11 7 11 2
49 11 11 1 11 2 11 2 11 13 9 0 1 9 9 9 11 11 11 11 11 2 15 3 13 9 15 13 1 9 11 11 15 14 0 1 9 16 11 11 11 11 11 7 11 2 11 11 11 2
27 1 9 11 2 11 13 1 12 9 2 3 2 13 9 7 9 1 9 15 3 9 7 0 1 9 9 2
28 9 9 10 13 9 2 9 7 9 2 2 11 2 11 11 2 3 13 11 2 2 11 11 2 7 11 11 2
14 1 9 9 1 9 10 2 15 15 14 13 11 11 2
41 11 11 11 13 9 2 9 2 9 10 9 13 1 9 0 1 11 2 9 10 9 9 11 2 11 2 3 13 12 9 2 11 7 11 2 3 13 1 9 9 2
11 9 15 3 1 13 9 9 15 3 0 2
24 11 15 13 3 13 11 11 2 7 1 10 9 7 9 2 9 13 9 16 0 1 9 11 2
20 11 13 13 2 13 9 1 11 2 15 3 13 1 11 11 11 2 11 2 2
12 3 9 7 9 13 9 15 0 9 14 13 2
18 1 9 2 1 9 2 3 1 12 5 9 9 2 11 2 13 9 2
17 11 15 13 9 10 13 1 12 12 11 5 1 9 9 9 10 2
17 3 0 3 2 9 10 15 0 1 10 9 11 3 13 1 11 2
19 9 10 10 3 13 1 9 12 9 2 7 9 13 1 9 12 9 9 2
16 11 1 9 10 3 13 1 10 9 13 11 7 11 15 13 2
27 1 9 12 2 11 13 3 10 9 15 3 13 9 9 7 10 9 0 7 13 9 1 9 9 15 0 2
10 9 10 13 9 12 9 1 9 12 2
50 13 9 9 12 5 12 2 9 9 1 11 1 9 9 7 14 2 9 13 1 13 1 11 11 0 1 9 12 9 15 13 2 9 11 11 11 11 11 7 11 2 15 3 13 1 11 12 5 12 2
14 11 11 13 12 9 1 9 1 1 10 9 1 11 2
31 13 12 9 7 2 11 1 11 2 2 10 9 0 1 9 11 7 9 11 2 13 1 10 9 9 0 13 9 9 2 2
18 9 10 2 9 1 9 14 3 13 5 13 7 3 13 9 9 10 2
15 15 13 9 10 13 9 9 9 0 1 9 13 9 9 2
17 1 9 10 2 9 9 3 13 9 13 7 13 9 15 13 9 2
38 3 13 1 9 9 9 9 11 2 9 9 0 3 13 2 1 9 11 11 2 9 9 2 9 2 9 2 11 11 2 11 11 9 2 7 0 9 2
24 16 11 14 13 1 9 9 10 3 13 2 9 9 9 15 0 1 9 9 9 15 7 14 2
16 13 9 9 11 1 9 15 13 9 16 9 13 9 9 9 2
21 11 13 9 0 12 9 15 13 1 9 9 1 12 9 7 9 3 9 12 9 2
25 9 15 13 13 9 2 9 11 2 7 9 9 3 11 2 7 2 3 10 13 3 0 2 0 2
31 0 1 9 1 9 1 9 9 9 9 1 9 9 11 11 11 13 1 9 12 9 9 2 13 1 11 12 1 11 12 2
26 13 0 0 1 11 7 11 2 9 9 9 11 11 13 1 11 11 11 2 11 11 11 2 11 11 2
4 11 9 12 2
10 16 9 14 3 13 1 9 15 13 2
24 1 11 13 9 9 0 1 11 3 11 11 2 0 11 11 2 7 11 11 7 11 11 11 2
37 3 2 9 10 13 1 9 13 12 7 12 9 2 16 1 9 12 9 13 7 9 10 13 16 9 3 13 12 7 12 9 1 3 13 9 10 2
33 1 9 11 13 10 9 1 11 11 2 12 9 15 13 1 11 13 1 9 10 11 1 11 7 13 12 9 11 7 13 10 9 2
26 11 10 13 13 1 9 12 2 12 2 11 11 11 13 9 9 15 0 7 15 3 13 1 9 11 2
13 11 9 10 3 3 13 1 11 2 3 1 11 2
15 12 10 9 13 1 9 0 2 7 3 12 10 9 13 2
40 12 9 0 9 11 13 1 9 11 1 13 9 2 9 9 1 13 9 9 11 11 15 0 7 9 9 11 11 11 2 15 3 13 1 9 10 1 12 11 2
26 9 10 3 13 1 0 1 9 9 2 11 11 2 11 11 2 11 11 2 11 11 2 7 11 11 2
13 9 13 1 9 9 7 1 9 10 2 12 9 2
20 1 9 0 10 16 11 11 11 14 13 0 2 1 13 11 11 1 11 11 2
58 11 10 13 10 9 2 1 1 13 3 13 9 15 13 9 15 14 3 13 11 2 7 14 13 9 1 9 2 16 9 10 13 9 2 3 9 3 0 7 3 13 1 11 7 11 2 16 1 9 10 9 3 3 13 1 10 9 2
4 0 9 11 2
10 9 10 13 0 2 7 15 13 0 2
19 9 10 13 1 13 9 2 9 15 3 13 9 9 15 13 1 0 9 2
25 11 2 11 11 2 2 13 9 9 9 0 1 11 11 1 11 11 2 12 13 1 12 11 12 2
24 9 10 3 13 1 9 10 9 1 11 2 11 2 11 2 11 9 9 2 9 9 1 9 2
10 7 12 9 14 13 16 10 3 9 2
16 9 7 9 13 9 15 13 3 0 16 1 9 13 9 9 2
18 3 10 9 10 0 13 1 9 9 2 9 13 9 0 15 0 13 2
12 1 9 12 7 12 2 15 13 11 11 11 2
31 1 9 1 9 12 2 9 11 11 13 2 16 10 9 0 15 13 13 1 11 11 2 3 9 1 9 9 14 3 13 2
12 12 2 1 9 13 13 1 9 1 10 9 2
2 13 2
16 11 13 9 1 9 11 11 2 11 11 2 11 11 2 11 2
13 11 1 9 12 13 11 2 11 2 11 11 9 2
19 15 13 1 12 9 12 9 9 9 7 13 9 9 1 11 11 2 11 2
10 9 10 15 13 9 9 3 9 10 2
18 9 9 10 3 13 9 9 9 9 9 9 7 9 7 9 9 0 2
36 10 9 15 13 13 9 1 9 15 0 1 9 2 9 11 7 11 11 11 2 7 9 9 1 9 10 0 1 9 9 1 9 11 7 11 2
22 10 9 13 16 15 13 9 1 11 2 16 13 7 3 13 10 9 1 13 1 11 2
23 9 1 9 11 3 13 16 9 9 3 0 7 3 3 13 1 9 13 1 9 13 3 2
53 10 9 1 9 15 3 0 2 3 9 1 10 9 1 9 13 0 1 9 9 15 13 2 7 3 9 1 9 9 13 2 16 9 13 1 13 13 9 10 2 7 7 9 10 9 9 13 9 10 1 9 9 2
33 16 9 15 13 13 1 9 2 9 11 13 0 2 9 11 11 13 9 9 2 9 11 2 1 9 10 1 9 11 1 9 12 2
7 13 9 0 16 11 11 2
20 16 12 9 9 11 2 11 2 11 9 2 7 11 2 11 11 2 2 13 2
19 11 15 13 9 2 9 12 2 13 13 1 9 0 2 0 2 7 0 2
11 9 9 9 15 3 0 3 13 9 10 2
18 9 9 9 13 9 2 16 9 0 3 13 12 12 9 9 1 9 2
8 0 9 15 13 10 14 13 2
37 3 9 2 9 13 2 1 9 12 2 11 13 1 9 11 7 1 13 1 11 2 11 2 16 2 1 9 15 13 9 9 9 1 11 11 11 2
17 11 13 9 15 13 1 11 11 2 11 11 2 11 11 2 11 2
14 16 15 13 9 0 2 15 13 13 9 7 13 9 2
22 11 11 2 11 11 2 13 13 11 13 1 10 9 1 13 9 1 11 13 12 9 2
12 9 10 13 0 9 9 9 15 13 9 12 2
21 11 13 10 10 9 15 13 1 11 11 11 2 11 11 2 11 11 11 2 11 2
7 3 11 1 11 3 13 2
13 11 9 3 13 1 11 1 11 2 11 7 11 2
16 11 13 10 9 1 9 11 11 2 11 11 2 11 11 11 2
27 9 10 15 3 13 12 9 16 11 7 11 2 10 3 13 9 1 9 2 9 15 3 3 13 1 11 2
15 16 9 15 13 1 9 2 11 2 13 1 9 11 11 2
10 15 13 9 15 3 13 1 9 10 2
23 11 11 13 1 12 11 12 1 11 2 11 11 11 11 11 15 13 9 11 11 7 11 2
22 15 3 13 1 9 9 2 11 11 2 1 11 11 11 2 11 13 9 12 1 11 2
10 11 3 13 1 1 9 12 1 12 2
36 9 1 9 2 9 10 3 2 3 13 2 7 9 0 13 1 11 11 15 13 9 9 2 9 10 3 13 9 1 9 2 9 0 1 12 2
25 9 10 3 13 9 9 11 2 13 13 12 9 9 9 9 15 13 1 9 1 13 9 15 13 2
17 1 9 9 2 11 13 9 1 11 11 1 11 2 11 2 11 2
44 3 13 9 9 1 9 11 2 11 1 11 2 3 11 2 1 9 12 2 7 13 1 9 9 0 1 11 11 1 9 12 2 15 3 13 9 1 9 15 0 1 9 12 2
11 3 15 15 13 9 1 13 9 11 11 2
25 11 3 3 13 1 9 0 1 13 9 7 9 9 7 9 10 9 2 3 1 9 15 13 3 2
20 16 15 15 13 1 9 13 1 9 10 2 15 14 13 13 16 9 13 11 2
17 7 16 11 11 13 12 2 12 9 1 11 15 13 9 1 9 2
10 10 9 9 3 13 13 13 1 9 2
25 9 9 10 13 0 13 9 9 3 0 15 13 1 9 9 15 3 0 1 9 9 7 9 9 2
36 9 9 11 9 1 9 9 9 9 13 1 13 9 11 2 1 1 3 13 9 1 9 9 1 11 11 7 9 10 15 3 13 1 9 9 2
11 9 10 15 13 1 13 9 11 1 9 2
28 11 11 13 13 9 2 13 9 9 9 2 9 9 9 2 9 2 1 13 9 2 9 0 2 1 9 0 2
15 11 9 11 2 11 13 9 9 1 11 11 11 2 11 2
18 11 13 13 9 2 15 13 9 1 10 9 9 2 0 9 1 9 2
2 3 2
11 11 1 9 12 2 13 9 1 12 9 2
31 16 11 11 3 13 9 1 13 9 7 13 9 2 9 15 2 11 2 11 11 2 2 11 3 13 1 3 13 1 11 2
39 9 9 10 13 1 11 11 2 12 2 12 2 2 15 3 9 1 9 10 12 9 13 1 10 9 0 1 11 7 3 1 10 11 11 2 11 11 2 2
15 11 11 13 10 9 1 11 11 11 2 11 11 2 11 2
14 11 13 9 1 9 11 2 11 2 11 11 2 11 2
7 7 9 9 15 3 13 2
44 7 13 1 9 15 13 1 11 2 11 2 9 10 13 11 2 1 13 9 11 2 11 2 11 13 11 11 11 2 11 12 2 2 11 11 7 11 11 1 13 11 11 11 2
13 3 11 11 13 11 11 11 5 11 11 11 11 2
10 11 9 13 12 5 1 9 12 9 2
33 9 9 0 9 10 13 9 11 2 12 5 2 2 9 11 2 12 5 2 2 9 11 2 12 5 2 7 11 2 12 5 2 2
18 11 11 11 13 9 9 9 0 15 13 1 9 11 11 7 11 11 2
7 0 7 14 9 15 10 2
22 1 9 9 2 9 9 9 3 3 0 1 9 2 1 3 9 15 13 1 9 9 2
18 16 11 3 13 9 11 2 7 7 11 1 11 2 7 11 1 11 2
16 12 9 0 10 3 3 3 0 13 1 11 11 11 11 11 2
7 11 10 13 1 11 11 2
7 11 2 15 15 3 13 2
8 11 11 13 9 1 9 11 2
10 2 11 2 14 15 0 1 9 11 2
74 9 2 9 11 15 13 9 1 0 2 11 11 2 2 2 11 2 2 2 11 11 2 2 2 9 11 2 2 11 2 2 2 11 2 2 2 9 11 2 2 2 11 2 2 2 9 2 2 2 11 1 11 2 2 2 11 11 2 2 2 11 2 2 7 3 9 2 9 9 11 2 11 0 2
20 15 12 1 11 11 2 9 9 1 9 11 15 3 13 1 11 11 1 0 2
9 2 11 2 1 9 15 9 10 2
12 9 9 9 7 15 13 15 14 13 1 9 2
6 2 3 14 13 9 2
10 3 9 11 11 7 11 13 1 0 2
28 9 10 1 9 2 9 10 13 9 9 9 9 9 13 1 9 9 0 9 15 13 1 9 9 12 11 12 2
33 2 2 9 11 2 2 10 9 0 1 11 2 3 13 0 1 9 2 10 9 0 1 9 11 2 3 13 0 1 9 9 2 2
22 1 12 11 12 2 11 11 13 13 9 1 9 0 2 1 11 11 11 1 0 9 2
15 11 10 13 12 1 12 9 7 9 15 13 1 11 11 2
34 3 9 9 15 13 9 15 0 2 9 0 2 9 2 15 13 1 0 1 9 2 9 2 9 9 2 9 2 9 0 2 7 9 2
20 1 9 11 11 9 12 2 11 11 13 13 12 2 1 11 11 7 11 11 2
17 16 13 9 2 15 13 11 13 11 11 11 7 13 2 11 2 2
26 1 9 11 12 2 11 13 9 1 13 9 2 9 9 1 9 0 1 10 9 1 9 9 11 11 2
15 11 10 13 12 1 12 9 7 9 15 13 1 11 11 2
11 16 2 9 11 13 1 11 2 7 9 2
8 9 9 13 9 13 9 11 2
13 1 3 13 11 2 10 9 9 3 13 3 3 2
14 3 11 13 9 9 0 10 9 1 3 1 12 9 2
14 13 13 11 10 2 2 3 15 13 9 15 0 10 2
9 9 15 3 13 1 9 9 9 2
7 3 15 13 11 1 11 2
10 14 15 10 11 7 15 13 9 11 2
19 3 1 12 9 2 12 9 9 10 13 2 3 9 15 3 3 3 0 2
14 1 3 2 9 1 12 9 3 13 1 9 15 0 2
21 11 11 13 10 10 9 1 9 11 11 11 2 11 11 11 2 11 11 2 11 2
23 15 14 13 16 15 3 13 9 2 9 1 12 9 15 0 11 0 7 3 13 1 13 2
32 11 11 11 13 9 15 13 13 1 11 11 2 11 10 3 13 1 9 15 13 1 9 2 9 9 15 13 13 7 14 13 2
32 11 15 13 3 13 9 1 11 7 11 7 11 13 13 9 1 9 0 7 13 9 11 11 11 11 15 3 13 11 7 11 2
14 11 0 13 9 13 0 0 1 9 7 9 13 0 2
14 10 9 0 15 9 1 13 9 15 13 1 9 10 2
38 9 10 13 9 9 9 16 11 2 11 2 11 2 15 13 9 9 7 9 16 13 1 9 0 2 15 3 13 1 9 15 13 1 9 12 9 10 2
42 3 13 9 0 9 11 2 11 1 9 11 11 11 11 2 11 11 2 11 2 9 12 2 11 2 11 13 13 1 10 9 1 13 9 10 9 2 3 13 9 2 2
16 15 13 9 2 9 1 9 2 16 15 14 3 13 15 0 2
22 1 9 12 2 9 10 13 9 9 1 12 9 7 13 9 9 12 2 12 12 2 2
38 11 15 13 10 9 13 1 9 11 11 11 11 2 10 9 13 9 0 2 16 9 9 13 9 9 2 9 2 9 2 7 9 13 1 9 15 13 2
47 11 13 0 10 13 3 1 10 9 0 1 9 2 9 2 11 2 2 2 11 2 11 2 11 2 2 9 2 9 2 2 2 9 2 9 2 9 2 9 2 10 9 1 11 0 2 2
22 11 11 13 9 15 13 1 11 11 2 11 11 2 11 7 13 9 0 1 9 11 2
18 11 11 11 11 2 2 2 3 13 1 11 2 13 9 9 0 11 2
11 11 12 3 9 0 2 0 7 0 2 2
72 11 11 1 9 15 13 11 11 2 11 13 16 2 9 15 0 3 13 13 11 2 11 2 2 11 2 11 2 11 7 11 2 15 13 10 9 15 0 1 9 1 11 7 11 2 15 10 13 9 1 11 2 11 9 0 7 3 13 1 11 2 9 0 1 9 9 13 1 9 7 9 2
20 7 14 3 13 15 13 7 13 1 9 15 13 11 11 2 12 2 12 2 2
26 15 13 2 11 11 2 2 10 9 13 9 1 11 2 10 9 9 11 15 0 2 13 1 9 12 2
7 11 9 10 13 1 11 2
26 16 13 9 9 15 15 13 16 15 13 11 2 11 3 13 2 2 16 9 0 14 3 13 2 2 2
25 9 10 11 11 13 9 9 9 0 1 9 0 7 9 7 9 15 0 1 0 9 9 1 9 2
15 11 11 7 9 11 13 9 15 13 9 11 7 11 11 2
11 11 13 9 1 9 0 15 13 9 0 2
55 9 1 13 9 1 10 9 9 13 1 9 12 2 9 9 9 1 13 13 9 15 3 13 1 2 9 11 11 11 2 1 9 2 9 10 13 1 9 9 9 7 9 9 9 15 3 13 7 3 3 9 13 9 9 2
21 9 15 13 1 11 13 13 11 2 11 11 11 13 16 3 13 9 9 11 15 2
31 16 11 13 9 2 3 9 0 9 9 11 11 3 13 9 2 16 15 13 1 13 9 2 9 0 10 1 1 9 11 2
39 3 2 11 11 2 13 11 2 11 9 1 9 0 13 1 13 9 1 9 1 9 9 0 1 9 13 1 9 0 2 13 9 1 9 0 7 9 9 2
14 11 13 9 15 13 1 13 1 12 9 9 15 13 2
10 9 10 3 13 1 11 7 1 11 2
10 11 13 1 11 13 14 13 9 0 2
36 11 11 11 7 11 13 9 1 11 7 13 9 15 15 13 9 11 12 2 11 10 13 9 15 1 13 10 10 9 9 2 11 2 1 11 2
40 1 13 9 0 9 10 2 11 11 11 11 3 13 9 1 12 9 0 2 16 2 11 11 2 11 2 2 2 2 11 11 11 2 7 2 11 11 11 2 2
16 12 9 10 13 16 9 11 3 13 9 9 0 11 11 11 2
54 3 1 13 9 2 9 11 2 12 9 12 9 12 11 12 1 9 2 9 9 3 13 9 9 9 1 9 9 9 12 9 12 2 1 9 15 0 9 9 9 1 9 11 11 1 9 0 13 13 11 2 12 9 2
15 1 9 9 9 14 13 9 2 16 13 1 10 9 9 2
19 9 2 9 11 2 11 2 13 10 9 1 11 15 13 0 9 1 11 2
13 11 11 11 2 2 2 13 9 9 9 1 11 2
24 1 11 11 11 9 11 13 3 1 12 9 1 12 9 1 9 9 10 13 7 13 1 12 2
33 16 14 13 9 2 16 9 13 1 0 1 11 11 12 2 15 3 13 9 9 1 9 11 15 13 1 9 12 11 1 9 10 2
18 15 3 13 9 15 2 13 9 15 3 9 7 13 9 15 2 2 2
44 11 2 11 2 11 2 13 10 9 9 9 15 13 1 9 9 9 11 2 11 2 13 1 9 11 11 2 11 13 1 11 1 9 9 2 11 1 9 2 7 11 1 9 2
34 11 2 9 9 9 11 15 0 13 11 11 15 13 1 11 7 13 9 11 0 1 9 7 13 1 9 11 11 11 11 1 9 12 2
14 14 0 13 9 2 9 13 1 9 11 1 13 9 2
14 11 2 11 11 11 2 13 1 9 9 11 11 11 2
65 11 9 11 11 1 9 11 11 11 1 9 11 11 7 11 2 11 2 3 0 2 3 1 9 12 3 13 9 1 11 2 12 2 12 2 2 2 12 11 12 12 12 12 12 12 12 12 12 9 9 2 1 12 9 11 2 2 3 0 13 0 9 15 13 2
34 11 11 11 12 13 9 12 2 12 9 9 9 11 11 9 12 15 13 1 11 11 11 2 11 2 11 2 11 1 9 12 11 12 2
17 11 9 0 1 9 13 1 12 9 12 1 9 9 9 9 12 2
25 1 13 11 2 9 0 9 9 9 3 13 1 9 7 9 1 9 13 3 13 9 15 0 0 2
29 11 1 9 10 13 2 9 9 15 0 13 1 9 11 11 2 2 7 3 2 13 1 9 2 9 9 11 2 2
36 7 3 0 3 2 1 13 10 9 9 0 1 9 7 9 2 3 13 2 13 10 2 9 9 9 9 9 1 9 15 3 13 1 10 9 2
20 9 9 9 3 0 3 3 13 2 2 15 0 3 0 7 15 0 3 0 2
26 9 11 11 13 10 9 0 11 15 13 9 0 13 9 10 10 9 7 9 9 11 15 13 1 11 2
18 1 9 2 15 13 11 11 11 1 9 12 2 15 13 9 9 9 2
29 1 9 12 11 12 1 9 9 11 11 9 12 9 12 9 2 12 5 12 5 12 2 11 13 13 11 11 11 2
13 9 12 13 1 11 12 2 11 12 1 12 9 2
8 11 11 13 9 0 3 11 2
22 11 15 13 13 10 9 15 10 2 10 13 1 12 9 16 2 11 2 11 7 11 2
18 11 9 10 13 0 1 9 9 15 13 1 10 9 1 9 0 9 2
43 15 12 9 15 13 9 1 9 1 9 12 9 2 16 15 13 16 10 11 2 11 11 2 16 14 13 1 9 15 0 2 3 9 3 13 2 16 1 9 12 13 9 2
19 11 11 2 15 3 13 1 11 2 13 10 9 9 0 1 9 11 11 2
3 0 3 2
4 13 9 11 2
53 3 1 9 12 11 12 9 9 2 9 9 12 11 2 11 13 13 9 11 11 7 3 13 11 1 9 12 2 12 2 9 10 13 12 2 12 9 7 1 12 12 1 9 0 1 12 9 5 9 1 11 11 2
28 16 9 7 9 9 0 3 13 9 1 9 2 9 9 15 13 9 1 9 0 3 0 1 9 0 1 13 2
44 11 11 2 11 13 13 1 9 12 16 10 9 3 2 9 11 13 7 9 10 13 9 1 9 0 2 0 1 11 11 2 9 12 7 9 15 3 0 1 10 11 11 13 2
23 9 9 10 13 9 9 12 11 2 2 16 13 9 9 1 12 2 12 9 2 12 2 2
24 16 9 1 13 11 11 3 3 3 13 16 15 3 3 13 16 13 9 13 9 15 13 0 2
12 11 11 13 9 15 13 1 11 11 2 11 2
9 15 13 1 9 1 11 13 11 2
7 9 9 11 1 9 10 2
16 15 13 10 9 9 2 11 11 11 2 13 12 11 12 2 2
27 11 15 13 1 9 11 2 11 13 2 11 15 13 1 9 11 2 11 2 7 9 11 2 15 2 13 2
10 9 10 13 9 0 1 9 11 11 2
31 10 9 3 13 9 1 0 2 16 10 9 3 13 16 14 3 13 9 2 16 16 3 0 2 7 3 13 12 9 9 2
28 15 13 11 9 2 11 11 2 11 2 12 2 12 2 7 11 11 11 2 11 2 11 2 12 2 9 2 2
12 9 15 13 1 13 9 12 11 2 12 9 2
29 11 13 1 11 11 7 13 1 9 1 13 11 11 7 11 11 1 9 12 2 12 2 12 2 2 12 2 12 2
23 1 9 13 3 13 2 2 11 11 2 11 11 11 11 11 11 11 11 11 11 11 2 2
32 1 9 12 2 9 10 13 9 9 1 12 9 7 13 9 9 12 9 2 2 9 10 13 9 9 9 12 9 5 9 2 2
25 11 11 11 2 2 13 10 9 9 9 13 9 15 13 1 9 12 2 11 3 13 1 9 9 2
11 11 13 10 9 1 2 11 11 2 11 2
21 11 13 9 0 1 9 1 7 1 9 1 10 9 11 2 7 0 1 9 9 2
19 12 9 10 13 1 9 11 0 1 10 2 13 9 9 7 9 9 9 2
5 9 10 3 0 2
26 9 12 2 11 13 1 11 11 11 2 12 2 1 11 11 2 7 9 0 11 11 11 2 12 2 2
7 11 13 9 1 12 9 2
18 11 11 13 10 10 9 1 11 11 2 11 11 2 11 11 2 11 2
25 16 9 15 0 10 15 13 9 15 0 0 2 16 3 3 13 10 9 9 2 1 12 9 0 2
44 9 15 3 0 1 11 1 9 3 13 1 9 10 2 15 3 13 9 1 9 9 11 2 13 9 9 11 11 2 9 9 9 2 9 9 2 11 13 7 9 9 1 11 2
17 16 13 1 1 11 11 13 1 9 0 1 9 7 9 1 9 2
28 9 10 13 1 11 11 2 7 13 11 11 2 11 11 2 11 2 11 2 11 2 11 11 2 7 11 11 2
10 9 3 13 1 9 9 11 2 12 2
27 15 13 9 9 1 11 11 11 1 9 11 11 2 12 11 1 9 12 11 12 1 9 1 11 11 11 2
17 11 15 13 1 11 2 11 13 3 13 1 9 0 7 9 0 2
14 9 15 3 15 13 1 9 0 13 9 1 9 10 2
20 11 11 2 2 13 10 9 9 9 9 2 9 11 11 15 13 1 11 11 2
21 9 1 1 9 11 11 2 3 2 3 12 2 12 5 2 16 1 9 11 11 2
28 11 13 10 1 9 7 13 9 15 13 1 9 0 1 9 7 13 1 1 9 9 0 7 9 2 9 9 2
7 9 3 13 1 13 9 2
17 11 13 1 10 10 9 9 1 11 1 13 11 11 1 9 12 2
16 1 9 12 9 9 10 13 9 13 9 1 9 11 11 11 2
28 11 13 0 2 9 9 0 12 12 11 2 9 2 9 9 2 9 9 1 11 2 2 9 9 0 12 12 2
7 9 15 14 13 11 11 2
16 11 11 1 9 11 0 2 11 11 2 2 13 0 1 11 2
11 3 2 9 9 11 13 3 1 12 9 2
13 11 13 10 9 9 1 11 15 13 1 9 12 2
9 9 10 13 9 9 11 2 11 2
7 9 0 1 9 7 14 2
16 15 13 9 11 12 1 11 2 15 13 9 1 9 12 1 2
24 1 9 10 9 3 13 1 10 9 11 2 15 13 9 11 2 9 15 13 2 1 10 9 2
29 11 11 15 13 1 9 0 13 9 13 3 0 1 10 9 7 13 13 1 10 9 2 13 1 11 11 9 12 2
22 1 16 11 3 13 9 7 14 1 9 2 15 13 1 9 1 10 9 9 15 0 2
38 16 9 10 13 1 9 15 3 13 1 9 9 9 13 2 16 1 9 9 10 3 13 10 9 0 1 0 2 0 16 3 13 9 9 1 10 9 2
11 9 0 9 10 13 1 9 12 11 12 2
34 1 9 7 9 9 10 0 13 9 1 13 2 1 9 11 2 9 0 11 7 11 2 7 9 9 9 9 7 9 13 0 11 11 2
58 15 3 13 1 10 9 2 1 11 11 2 11 11 9 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 2 11 11 2 7 11 11 2
23 3 2 16 10 11 11 10 13 14 0 16 9 9 15 3 2 2 11 13 9 1 11 2
21 11 13 9 0 1 9 12 12 11 2 7 9 11 12 11 7 9 9 12 11 2
14 1 15 2 12 9 10 3 13 13 1 12 11 12 2
19 9 11 11 13 9 12 9 1 11 11 11 2 11 2 11 11 2 11 2
23 1 11 2 11 13 9 1 9 2 9 9 9 2 9 0 2 7 9 0 15 3 0 2
19 9 9 15 0 13 9 15 13 13 1 10 9 15 13 7 13 1 9 2
76 1 9 12 9 13 1 13 9 9 13 9 9 11 2 3 9 11 15 13 1 10 11 11 2 10 9 7 11 13 1 13 10 9 13 11 11 11 11 11 15 13 1 13 9 9 2 9 9 2 9 2 2 7 9 1 9 11 2 15 13 9 1 12 9 12 2 13 1 10 9 9 0 2 9 2 2
6 3 15 13 1 9 2
40 1 9 12 9 11 15 13 9 11 13 12 9 2 16 2 1 11 2 9 9 0 15 13 1 9 12 2 16 9 9 1 12 9 7 9 9 1 12 9 2
21 3 2 1 9 15 13 1 11 11 2 11 10 13 9 16 15 13 11 1 9 2
22 11 11 13 10 10 9 15 13 1 11 11 11 2 11 11 11 2 11 11 2 11 2
12 16 3 13 1 9 9 10 11 13 13 9 2
3 1 1 2
3 15 9 2
48 11 2 2 13 9 0 15 13 15 13 1 9 11 2 9 10 3 13 1 11 9 1 9 9 2 1 9 11 1 9 11 7 1 11 0 2 7 3 3 13 1 9 9 0 7 11 9 2
21 9 2 9 10 13 0 2 3 2 1 13 9 3 0 2 1 1 9 7 9 2
17 1 9 9 7 13 9 9 2 13 9 10 9 1 1 9 9 2
17 11 10 13 9 9 12 9 2 2 1 13 9 9 1 12 9 2
27 11 2 1 2 13 10 9 13 15 13 1 1 9 7 9 0 2 7 9 9 9 15 13 1 9 0 2
8 9 3 2 9 10 13 3 2
15 9 10 13 1 1 11 11 11 7 10 9 1 11 11 2
12 15 3 3 13 11 11 11 1 12 11 12 2
13 9 9 3 13 1 9 11 1 9 11 1 11 2
32 1 9 2 9 15 13 9 10 13 9 16 13 9 9 7 9 2 9 0 15 13 1 9 3 13 12 1 12 9 11 10 2
34 1 9 15 3 0 1 11 11 11 2 11 13 11 1 13 11 11 2 11 2 7 11 11 13 1 11 11 1 11 1 9 13 11 2
4 15 14 13 2
20 9 9 3 13 1 9 9 9 1 13 9 9 11 11 15 13 9 9 9 2
21 11 11 3 13 12 9 0 11 11 1 9 12 7 1 9 12 1 11 11 11 2
24 9 11 3 13 1 9 1 11 1 9 11 15 13 1 11 2 16 9 9 10 3 3 13 2
17 10 9 1 9 3 13 1 9 9 7 9 1 13 16 14 13 2
7 9 0 13 9 1 11 2
14 9 10 13 1 9 11 11 2 11 11 2 12 2 2
20 9 10 13 9 1 9 9 12 11 11 11 11 1 9 9 13 7 9 0 2
21 1 9 2 13 12 9 9 2 9 0 13 1 13 9 7 9 15 13 9 9 2
18 3 13 13 9 10 2 10 9 9 7 10 2 10 13 10 9 9 2
13 9 9 13 1 9 0 1 9 15 14 13 9 2
10 9 9 9 11 12 13 9 11 12 2
82 16 9 0 1 9 9 9 13 1 9 12 1 9 3 1 2 12 2 12 5 2 16 13 2 13 9 9 9 1 12 9 10 13 1 12 2 12 5 16 16 13 1 12 9 0 9 0 2 0 9 3 1 12 2 12 5 2 1 13 10 9 9 1 0 2 0 7 1 9 15 13 1 9 9 12 13 9 9 13 3 0 2
16 11 3 13 9 1 9 9 10 2 16 9 3 13 9 9 2
39 10 13 9 1 11 11 11 2 11 9 11 9 1 9 11 11 2 11 9 0 2 11 11 2 11 11 2 11 11 2 11 2 11 11 7 11 9 0 2
14 16 10 9 11 0 13 10 9 1 9 9 1 13 2
22 1 9 12 11 12 2 9 10 13 9 16 9 9 13 9 13 15 1 9 9 0 2
28 1 12 9 2 9 2 9 11 13 9 10 1 13 1 10 9 15 13 11 11 7 13 11 2 9 9 2 2
18 1 9 15 0 7 14 13 9 2 9 0 3 13 1 9 0 0 2
15 1 13 2 9 15 13 1 9 12 10 0 0 1 9 2
19 3 15 14 13 1 2 16 15 13 15 1 9 7 9 1 9 7 9 2
14 11 13 9 1 9 11 2 9 2 11 11 2 11 2
16 11 13 9 9 12 1 9 9 11 2 10 9 9 1 11 2
14 2 11 2 15 1 13 7 9 10 13 9 9 13 2
17 9 0 13 11 11 11 2 11 11 2 11 11 2 7 11 11 2
20 10 9 15 14 13 1 9 9 13 1 9 15 13 9 9 1 11 11 11 2
10 11 11 2 2 13 10 9 1 11 2
25 16 7 11 11 7 9 11 13 1 11 2 11 11 2 3 15 13 0 9 1 9 9 9 9 2
26 9 9 1 11 11 3 13 1 9 9 7 3 13 2 13 1 10 2 9 0 9 9 13 9 11 2
26 9 11 1 13 9 9 3 13 9 2 16 14 3 13 16 13 10 9 15 3 13 1 9 11 11 2
14 11 3 13 9 9 2 1 9 11 2 7 11 2 2
7 3 11 3 3 13 9 2
8 1 9 10 13 9 11 11 2
12 11 12 3 13 9 9 1 0 1 11 11 2
33 11 11 11 12 7 9 9 11 11 11 11 11 12 13 10 9 11 11 11 15 13 1 11 2 11 11 12 2 11 11 2 11 2
16 11 11 13 9 1 9 11 1 11 15 13 1 13 9 9 2
7 9 10 13 1 9 12 2
34 11 13 9 9 9 15 0 7 0 15 13 11 11 2 13 1 9 1 11 11 7 11 2 7 1 13 9 1 13 9 2 9 0 2
15 9 10 13 1 11 11 2 7 1 11 11 1 9 11 2
22 7 9 10 3 13 9 0 15 14 13 11 13 15 3 14 13 9 9 1 11 11 2
11 11 9 3 13 9 2 9 2 7 9 2
20 9 9 13 3 3 3 2 3 1 13 16 11 3 13 9 0 1 3 9 2
21 1 10 9 11 13 13 1 9 0 13 9 2 11 2 15 15 3 13 1 11 2
14 1 9 2 11 13 1 9 15 0 2 0 7 0 2
29 9 9 10 14 13 13 11 11 7 13 12 9 1 9 12 1 12 2 16 7 9 0 9 13 13 1 11 11 2
22 9 10 1 9 2 9 2 9 2 9 2 9 9 7 9 2 9 9 13 1 9 2
17 9 2 9 0 15 13 13 9 11 1 11 3 13 9 15 0 2
22 1 12 9 0 2 9 11 3 0 0 2 16 15 3 13 0 13 9 1 9 9 2
20 3 10 9 15 13 2 3 3 13 1 9 9 1 9 9 9 9 15 0 2
15 9 9 13 10 10 9 9 15 13 1 11 12 1 11 2
21 11 11 13 9 11 11 1 11 1 9 12 7 9 3 2 15 13 9 11 11 2
10 9 9 13 11 2 16 9 13 11 2
52 7 2 1 9 2 11 11 13 10 9 2 9 2 12 1 12 9 7 12 1 12 9 2 7 9 9 2 12 1 12 9 2 2 9 9 2 10 9 2 7 10 9 9 7 9 9 15 9 10 3 13 2
26 11 15 13 1 10 9 0 1 12 9 2 9 11 12 9 1 9 2 7 10 0 9 2 9 0 2
17 11 13 10 9 7 13 1 11 11 11 2 11 11 2 11 11 2
25 9 9 15 13 2 16 11 2 11 0 1 9 2 3 3 13 1 9 9 9 1 9 9 10 2
25 11 2 9 1 11 11 11 9 7 11 11 11 1 9 11 13 0 9 0 11 1 9 9 11 2
24 9 9 9 10 1 13 9 9 1 9 9 1 9 9 7 13 1 9 9 1 9 3 0 2
14 11 13 0 7 9 15 13 9 7 13 10 9 0 2
11 11 10 13 9 9 10 0 13 9 11 2
13 15 13 16 9 11 13 9 9 7 3 13 15 2
41 1 9 2 9 2 9 9 15 13 13 0 10 3 13 2 1 9 11 11 2 11 11 2 11 11 2 11 11 11 2 11 11 11 2 11 11 2 11 11 9 2
20 10 9 3 3 13 11 15 13 9 9 15 9 2 9 3 13 13 1 9 2
19 11 11 11 2 2 2 13 9 9 9 9 1 9 15 13 1 9 0 2
8 11 13 3 11 14 13 3 2
18 1 9 15 0 2 11 13 9 0 15 13 9 15 13 9 9 11 2
4 13 9 11 2
12 9 7 9 10 9 9 10 15 13 9 9 2
12 13 3 1 10 11 0 15 3 13 9 0 2
14 9 9 13 9 15 13 9 1 13 7 13 9 9 2
23 0 9 12 11 12 2 11 11 13 13 1 11 2 11 2 11 7 11 2 11 2 11 2
10 2 2 9 15 3 13 9 1 9 2
16 9 0 15 0 1 9 9 9 10 13 1 9 9 3 13 2
29 16 9 10 3 13 9 2 16 9 15 0 1 9 9 14 13 9 7 9 15 13 1 9 2 9 15 3 0 2
16 3 2 15 3 13 1 11 11 7 13 12 9 7 12 9 2
20 1 9 12 1 12 2 11 13 3 13 1 11 13 15 13 1 11 11 11 2
10 9 0 15 13 11 7 13 1 11 2
17 9 10 13 1 9 9 9 15 0 2 13 1 9 9 9 11 2
36 11 11 11 2 11 11 11 2 12 11 12 2 12 11 12 2 13 10 9 11 11 2 7 3 10 9 2 9 2 9 9 2 9 7 9 2
24 9 9 10 1 12 9 1 9 9 9 2 15 13 1 12 9 1 1 9 15 13 9 10 2
29 11 11 11 13 10 10 9 9 2 9 9 11 11 15 13 1 9 11 7 11 11 2 11 11 2 11 11 11 2
15 11 11 13 10 9 9 1 9 9 11 11 2 9 11 2
70 9 0 15 13 1 11 11 7 11 11 13 0 1 11 1 13 9 7 13 1 9 0 11 2 16 9 0 1 11 11 2 11 11 2 7 11 11 3 13 9 15 1 10 9 15 1 11 7 9 0 11 2 9 9 9 15 13 1 9 12 13 9 9 11 11 1 9 9 12 2
22 7 9 2 7 9 2 0 13 9 11 2 16 15 13 13 15 7 13 1 9 15 2
32 11 10 13 1 7 13 1 11 11 2 10 9 0 15 13 1 9 11 11 11 2 11 11 11 7 11 11 11 1 9 9 2
12 7 9 0 13 2 15 15 3 0 1 15 2
20 11 11 2 11 11 13 9 9 12 11 10 13 1 9 11 11 2 11 11 2
15 7 3 9 11 3 0 13 11 15 3 3 13 10 9 2
10 11 7 9 13 10 9 9 15 13 2
22 1 9 10 2 15 13 1 9 9 7 13 9 9 2 3 13 9 15 0 1 15 2
8 11 10 13 1 11 9 12 2
12 11 2 2 13 10 9 1 9 11 1 11 2
41 11 3 13 1 10 9 9 9 2 15 13 1 9 2 9 2 9 2 9 2 7 9 2 11 9 2 3 0 1 9 9 15 0 1 9 2 9 2 7 9 2
14 10 9 3 9 9 13 2 3 9 9 7 9 13 2
25 1 9 2 11 14 3 13 1 11 2 16 0 1 13 1 9 11 11 15 13 1 11 9 12 2
36 9 10 3 13 0 1 12 9 0 2 1 9 15 13 1 12 9 1 12 2 8 13 12 10 9 3 2 7 1 9 13 9 9 2 9 2
35 1 1 13 9 9 1 9 15 13 7 13 9 9 2 9 2 1 9 1 13 1 9 0 2 13 1 9 15 3 3 13 2 9 2 2
47 9 10 13 1 12 11 12 11 11 9 10 13 11 11 11 9 12 2 12 1 11 11 5 11 11 11 11 2 11 11 11 13 9 9 11 11 11 11 11 1 11 15 13 1 11 11 2
27 1 9 12 7 3 11 13 9 1 9 0 1 9 2 9 2 9 9 7 9 9 1 9 12 2 12 2
28 11 9 10 13 1 13 10 9 0 15 13 9 11 16 10 9 10 13 2 13 10 9 1 10 9 15 13 2
20 1 10 9 9 9 14 13 13 9 11 11 11 2 16 3 1 13 9 0 2
9 11 11 13 9 11 1 9 11 2
10 9 10 13 9 3 0 9 1 9 2
24 15 13 9 1 11 11 11 1 9 11 11 11 1 9 12 11 12 1 9 13 11 11 11 2
11 11 11 13 9 9 15 0 1 11 11 2
22 11 13 9 13 1 9 7 9 15 13 12 9 15 3 0 1 9 9 12 2 9 2
23 11 11 13 10 10 9 15 13 1 11 11 11 2 11 11 11 2 11 11 11 2 11 2
25 1 9 12 2 15 13 1 11 1 13 9 9 9 1 11 11 12 1 9 9 0 1 12 9 2
13 11 13 9 9 9 1 9 12 9 12 2 12 2
24 11 11 13 9 9 2 9 15 13 1 11 11 2 11 2 11 2 11 2 11 2 7 11 2
22 11 15 0 2 15 3 9 1 13 2 14 3 3 3 1 0 13 9 1 15 0 2
51 11 11 2 15 13 9 2 9 9 7 10 9 9 9 2 13 10 9 2 9 12 2 12 2 1 9 9 10 1 9 9 2 5 5 8 2 9 2 9 2 9 5 9 2 9 2 9 15 15 13 2
33 1 11 11 11 15 10 9 15 3 0 13 12 9 1 11 2 9 9 0 15 3 13 9 9 2 7 11 2 9 1 9 2 2
23 11 11 13 9 9 9 15 13 1 11 11 11 11 2 11 11 11 2 11 11 2 11 2
15 3 11 13 9 2 13 9 9 7 3 13 9 1 9 2
45 10 9 13 16 9 1 2 9 10 3 0 2 7 12 9 9 9 0 15 13 1 9 12 1 13 11 7 11 2 11 11 11 7 11 11 2 14 3 13 13 9 12 9 10 2
19 11 13 9 9 9 0 1 9 1 11 15 13 13 1 9 12 2 10 2
66 11 11 11 1 11 11 2 11 11 11 13 10 9 15 13 3 1 9 10 13 10 9 0 15 3 0 2 7 13 1 9 15 13 9 0 15 1 2 11 11 11 11 1 9 12 2 12 1 9 2 9 10 3 13 10 9 9 2 9 10 3 13 9 13 9 2
18 10 10 9 0 13 1 13 9 0 2 11 1 9 1 9 9 11 2
12 16 9 10 3 13 2 9 3 3 13 15 2
20 9 13 11 10 10 16 15 3 13 9 1 9 2 14 13 9 1 9 9 2
77 10 13 9 0 1 9 11 1 11 7 13 9 1 9 15 3 0 1 9 9 9 1 3 2 9 13 9 1 9 1 9 2 2 3 9 9 0 15 1 11 14 13 1 13 0 1 9 2 7 1 15 13 1 12 11 1 9 15 15 0 7 3 14 3 3 9 1 15 1 9 15 3 13 7 9 9 2
43 11 11 11 11 2 11 13 9 0 11 11 11 11 2 11 11 11 11 11 11 11 11 11 11 11 11 11 11 11 11 10 2 11 11 2 11 11 2 11 11 2 11 2
23 1 9 2 9 9 1 9 2 14 13 9 9 2 9 1 9 15 13 1 9 10 0 2
12 1 10 2 15 13 16 0 3 13 10 9 2
21 16 2 3 9 9 13 16 9 0 1 0 2 7 3 1 0 2 1 9 9 2
17 11 14 13 9 9 2 16 13 9 7 9 1 11 11 2 11 2
15 11 3 13 9 15 3 13 1 9 14 9 1 1 9 2
72 9 9 2 9 2 16 14 9 1 11 15 10 2 3 13 1 1 9 10 2 15 13 1 11 11 2 13 1 11 11 7 11 11 11 2 7 13 9 11 2 11 2 11 2 11 2 7 11 11 2 10 3 13 9 15 0 2 0 1 11 11 2 11 11 2 11 2 11 11 7 11 2
11 11 10 13 9 9 10 0 13 9 11 2
12 15 3 13 9 11 1 9 9 2 9 9 2
14 11 3 13 1 13 9 0 1 9 9 9 13 0 2
12 11 13 10 9 2 11 2 1 11 2 11 2
42 1 10 10 9 0 11 2 11 11 11 2 15 13 3 13 1 9 12 9 2 14 3 13 16 16 10 9 13 1 1 9 0 2 9 15 0 7 3 13 9 13 2
22 9 1 9 10 15 3 13 1 10 9 9 11 11 13 10 9 7 1 9 3 13 2
18 13 0 1 9 15 9 9 0 2 14 13 2 1 9 9 15 0 2
23 9 0 3 0 9 13 1 13 9 2 9 0 2 1 9 10 2 3 9 1 9 9 2
14 13 12 9 9 0 7 0 1 11 11 1 9 9 2
35 11 2 11 2 11 11 2 2 13 9 9 9 11 15 9 10 13 1 11 11 11 2 1 9 9 1 11 11 2 15 13 10 9 9 2
22 11 11 13 10 10 9 15 13 1 11 11 11 2 11 11 11 2 11 11 2 11 2
6 9 12 9 1 9 2
17 11 11 1 11 11 13 11 1 13 2 2 11 11 11 2 2 2
51 1 1 9 0 10 13 9 11 2 11 2 9 11 11 2 2 11 11 2 9 11 2 2 11 2 11 11 2 9 11 2 2 11 11 11 2 9 11 2 2 7 11 2 11 2 9 11 5 11 2 2
30 1 9 9 1 13 9 2 10 9 9 1 11 2 15 13 1 11 2 11 2 11 2 11 2 7 13 11 12 11 2
35 16 11 11 13 1 13 1 11 2 9 9 13 1 14 13 15 3 2 15 3 13 1 13 1 15 2 15 13 16 15 13 10 9 9 2
15 11 11 13 9 11 15 13 1 0 1 11 7 11 11 2
18 1 9 0 2 9 9 3 13 3 1 9 1 9 9 9 15 0 2
7 9 9 7 9 9 9 2
5 3 9 13 11 2
11 15 13 3 1 12 2 12 12 9 9 2
16 7 1 9 15 0 13 12 9 9 9 3 11 7 11 11 2
109 9 9 11 11 16 13 1 9 0 9 9 9 3 13 16 9 9 0 1 9 9 7 9 3 13 9 0 1 11 2 1 9 0 1 9 9 9 9 7 9 2 9 9 7 9 9 7 9 9 15 3 13 9 0 7 9 9 15 3 0 9 9 9 9 1 11 13 1 12 9 2 1 9 9 9 9 2 7 9 9 9 7 9 1 11 11 13 2 11 11 13 1 11 11 2 11 11 2 1 11 11 11 12 1 9 11 11 12 2
26 9 0 9 10 13 1 13 9 0 2 9 0 9 2 7 13 9 9 1 9 9 9 7 9 0 2
33 9 11 11 13 9 9 1 11 11 1 11 11 12 1 11 11 2 9 11 7 10 9 13 9 11 1 11 11 12 1 11 12 2
16 9 9 9 10 13 3 1 13 9 9 1 9 9 9 0 2
6 11 2 9 10 9 2
33 11 13 9 0 11 15 13 1 9 2 9 11 2 7 13 16 15 13 9 0 7 0 1 10 9 15 9 1 9 10 9 11 2
17 16 3 2 9 2 9 9 13 13 9 9 1 7 1 10 9 2
51 9 0 15 15 13 13 9 9 2 15 13 10 9 15 14 0 7 13 9 9 0 2 1 15 3 15 13 16 13 9 11 1 9 15 15 13 16 13 10 9 9 9 0 1 13 9 9 1 9 15 2
32 16 3 13 3 9 15 13 1 9 2 13 11 11 11 2 3 13 9 15 0 2 0 13 9 2 9 9 9 10 1 11 2
35 1 13 9 2 9 1 9 15 13 9 7 3 3 13 0 1 9 9 11 2 9 1 9 12 11 12 13 9 1 9 0 9 9 10 2
35 11 2 12 11 13 1 9 9 0 1 9 11 1 9 12 11 2 12 2 1 13 9 13 1 9 0 1 12 9 1 9 9 9 12 2
22 9 0 9 13 1 9 0 15 0 13 9 9 15 0 0 7 9 9 11 11 11 2
7 1 10 9 9 10 3 2
15 15 13 1 2 11 13 9 1 11 7 11 1 11 11 2
34 9 10 3 13 1 11 11 2 11 2 11 11 2 7 9 11 11 11 1 11 11 11 1 9 11 2 12 9 12 10 9 12 9 2
21 11 11 2 11 2 11 11 15 0 3 13 1 9 2 9 9 11 15 3 13 2
33 1 12 11 12 2 12 11 12 2 15 13 11 11 11 11 11 11 2 15 3 13 11 11 11 1 12 11 12 1 12 11 12 2
14 11 3 11 14 13 14 0 3 1 9 7 9 15 2
13 1 12 9 12 11 2 11 11 13 9 11 11 2
37 16 9 10 9 0 2 9 2 9 0 7 9 1 9 10 3 13 1 9 9 2 9 2 9 9 2 9 9 2 9 2 9 2 9 7 9 2
13 9 10 13 1 11 11 2 11 2 12 11 12 2
2 11 11
45 9 10 13 1 9 9 9 1 11 11 7 11 11 11 13 9 9 11 9 12 11 12 1 11 11 11 2 16 11 13 0 9 16 13 9 1 12 9 3 2 3 1 9 0 2
28 11 11 11 11 11 13 1 11 11 2 2 13 10 9 9 9 13 11 15 13 1 9 11 11 1 9 9 2
11 9 10 13 1 9 11 1 12 11 12 2
27 16 3 1 9 12 11 12 2 11 11 11 12 13 9 13 9 11 11 1 11 11 9 12 2 12 2 2
20 11 11 13 9 0 1 9 0 11 2 9 9 9 9 9 11 1 11 11 2
23 1 13 12 9 2 9 13 9 0 1 11 11 7 11 11 11 11 11 1 12 11 12 2
31 11 11 11 13 9 9 2 3 1 11 11 2 11 2 11 2 1 9 9 11 11 11 2 11 2 11 7 0 9 2 2
7 11 0 11 13 9 0 2
10 3 15 13 9 15 1 10 15 13 2
13 1 9 1 9 3 13 16 2 9 2 13 9 2
43 9 9 0 1 9 9 10 13 12 9 15 13 1 12 9 0 13 7 12 9 0 0 0 1 2 1 9 9 12 9 7 9 9 0 2 9 5 12 2 12 2 12 2
25 9 1 9 15 13 11 7 11 13 15 0 2 7 1 15 13 2 13 9 9 3 13 9 15 2
19 9 15 14 0 1 11 11 11 7 11 11 11 2 13 9 10 3 0 2
28 10 9 9 13 9 9 9 15 0 1 9 2 9 2 2 13 1 9 12 1 9 15 0 2 1 9 12 2
17 9 11 16 3 13 7 9 1 15 1 2 9 0 2 15 13 2
116 9 10 13 1 9 9 9 11 2 1 12 9 1 9 1 11 2 11 11 11 7 12 9 1 9 1 11 2 11 2 11 11 11 11 2 11 11 11 2 11 2 9 9 7 9 9 1 11 11 2 11 11 11 11 11 2 11 11 11 2 11 2 11 9 9 9 1 11 11 2 11 11 11 2 11 2 11 11 11 2 11 2 2 11 11 11 11 2 2 11 11 11 11 1 11 11 2 11 11 2 11 2 11 11 11 2 11 2 11 11 11 11 1 9 9 11
13 9 0 13 1 10 2 10 9 9 9 7 0 2
34 15 13 11 11 11 2 11 2 11 11 2 7 11 11 2 1 11 11 12 2 9 12 9 2 15 13 1 11 11 15 13 12 9 2
26 9 1 11 2 3 12 1 12 9 15 13 13 9 3 13 9 9 1 9 9 11 11 2 11 12 2
10 9 10 3 13 0 1 9 11 11 2
25 1 9 0 2 9 9 2 9 2 9 1 9 2 13 1 9 9 9 15 3 13 1 9 10 2
23 11 13 1 9 11 11 11 11 15 13 1 2 9 9 2 1 9 2 9 7 9 10 2
14 9 9 12 2 12 12 2 1 9 9 5 12 9 2
12 1 9 0 2 15 13 1 11 11 7 11 2
13 11 12 13 10 10 9 9 9 9 11 11 11 2
15 1 9 9 9 3 13 1 9 9 9 15 3 13 1 2
27 12 2 11 13 9 1 11 2 11 13 1 11 2 12 2 9 0 11 11 1 11 1 10 9 15 13 2
84 11 2 11 5 11 5 11 5 11 2 9 5 9 2 8 5 9 2 13 10 9 2 9 5 9 2 11 1 13 9 15 13 9 2 13 1 2 9 9 9 9 1 9 9 2 9 2 9 2 2 1 9 2 9 2 9 0 2 13 9 2 9 9 2 9 9 2 7 9 2 9 9 9 2 9 2 7 2 9 2 13 7 13 2
17 16 2 9 0 1 9 10 14 13 9 1 11 11 1 9 12 2
25 11 11 13 9 1 13 1 9 9 9 9 10 13 9 9 7 9 9 9 9 11 15 3 0 2
8 9 10 14 13 1 9 10 2
24 3 9 2 15 13 10 9 9 1 12 2 12 9 0 9 2 15 14 13 9 9 13 9 2
24 15 3 13 11 11 2 11 11 2 9 11 7 2 1 9 12 2 9 0 11 1 9 12 2
29 11 2 12 11 11 13 9 1 11 2 12 11 15 3 13 12 9 1 12 9 1 11 1 9 0 13 12 9 2
9 1 10 15 13 9 0 1 11 2
19 16 2 1 12 2 13 9 0 10 11 9 0 11 15 13 9 1 12 2
25 13 3 1 12 3 9 15 13 1 2 2 9 15 13 0 1 11 2 14 13 15 13 0 2 2
6 9 10 13 9 12 2
31 11 13 12 10 13 9 9 11 2 9 10 13 1 11 11 2 11 13 9 1 11 11 7 11 2 0 9 0 1 11 2
17 11 11 13 11 1 13 9 11 2 11 15 13 1 9 9 11 2
19 11 13 9 9 1 9 1 9 2 2 11 2 7 9 1 9 12 5 2
18 9 10 13 1 11 11 2 11 11 2 11 11 2 7 3 3 3 2
34 16 15 13 9 2 16 13 9 10 1 9 0 2 9 2 9 2 9 2 7 1 15 15 13 9 15 3 0 7 3 0 1 9 2
16 13 1 11 2 11 7 11 16 13 1 11 11 1 9 12 2
11 9 9 15 3 13 1 11 11 11 11 2
13 11 13 9 11 11 2 11 2 11 11 2 11 2
17 11 13 1 9 11 11 11 2 15 1 9 11 1 0 13 9 2
13 3 11 13 9 3 1 13 9 7 9 1 9 2
12 14 11 15 13 2 2 14 9 15 13 3 2
19 11 13 1 10 9 1 2 0 2 0 12 7 1 2 11 11 11 2 2
6 9 10 13 12 9 2
54 2 11 11 11 9 9 9 9 2 11 2 9 2 11 2 2 7 2 11 2 2 13 9 9 9 1 9 0 0 2 2 15 2 2 15 13 1 9 0 2 9 2 13 2 7 2 13 2 1 9 2 9 2 2
36 1 9 12 2 12 2 11 13 9 9 11 1 11 11 2 11 13 1 11 11 10 2 12 2 13 11 11 11 2 1 11 12 1 9 12 2
20 11 10 13 9 9 12 12 2 2 1 13 9 9 1 12 9 2 12 2 2
16 11 2 9 15 13 13 1 1 9 9 11 11 11 11 11 2
54 11 2 11 11 7 11 11 2 13 10 9 0 9 2 11 11 11 2 15 13 1 9 12 11 12 1 11 2 15 13 9 1 9 13 9 9 15 0 2 11 11 2 7 9 9 9 1 11 2 3 1 9 0 2
23 1 10 11 11 10 3 13 1 9 9 7 9 11 15 13 1 11 15 13 1 11 11 2
18 11 11 1 9 11 3 13 9 9 7 9 15 0 1 9 9 9 2
24 9 9 3 13 9 0 1 9 16 3 13 1 9 2 9 9 2 9 15 13 9 7 9 2
6 9 0 13 9 9 2
7 11 11 13 9 9 9 2
37 16 15 3 13 9 9 9 9 0 9 11 2 11 7 11 2 7 3 13 10 9 9 1 9 9 11 2 11 13 13 9 15 3 13 9 9 2
17 9 0 2 9 9 0 2 9 9 0 2 0 2 9 0 0 2
15 11 11 13 10 9 15 13 9 12 15 13 9 11 11 2
26 11 11 13 1 9 12 11 12 1 0 9 11 1 12 5 9 9 11 2 11 2 13 9 0 11 2
8 7 15 15 13 9 9 10 2
29 9 10 3 13 2 7 1 9 9 11 11 11 11 11 2 3 13 9 1 11 15 13 9 3 1 9 9 15 2
10 11 11 13 9 9 9 15 3 0 2
11 11 12 1 0 13 1 2 11 11 2 2
18 9 10 13 9 1 12 9 7 13 9 9 1 12 9 1 9 12 2
24 11 2 9 13 10 9 9 9 9 0 7 9 0 2 1 9 11 1 1 0 13 1 9 2
16 9 15 3 13 2 3 15 14 13 15 13 1 9 1 9 2
16 11 13 9 11 1 9 9 13 0 2 0 9 7 9 9 2
18 1 9 12 2 11 13 1 9 1 9 1 11 7 13 1 11 11 2
36 9 11 12 13 9 9 9 9 1 11 11 12 1 11 1 11 2 9 2 9 9 11 11 12 2 12 13 11 1 11 2 9 11 11 12 2
16 11 3 13 12 9 11 2 3 11 2 11 2 11 7 11 2
31 9 3 3 3 1 13 9 9 10 16 13 3 13 10 9 9 15 0 2 3 13 7 13 1 9 11 1 9 9 11 2
6 9 13 1 0 9 2
20 13 2 11 2 16 9 11 11 11 11 13 11 11 11 15 13 1 9 11 2
11 9 9 1 11 13 13 9 9 1 9 2
17 1 12 11 12 13 9 1 9 11 15 13 13 9 7 9 0 2
22 10 9 13 11 1 11 5 11 11 2 11 2 13 9 0 15 13 9 9 9 10 2
8 16 3 13 10 9 1 11 2
9 9 0 16 9 9 3 3 13 2
15 1 10 3 2 15 14 13 1 9 9 2 9 9 0 2
5 11 11 11 12 2
12 16 9 13 1 11 11 2 11 2 11 11 2
24 11 13 10 9 1 9 11 2 11 2 11 1 9 11 2 11 2 11 1 9 2 9 11 2
23 11 15 13 1 9 13 13 9 9 1 9 11 15 0 1 13 1 9 9 15 3 13 2
6 9 9 9 1 9 2
13 11 13 9 9 15 13 0 15 13 1 11 11 2
13 1 12 2 12 15 13 9 9 1 11 11 11 2
19 16 13 9 11 11 11 11 2 15 3 13 13 9 11 1 11 1 12 2
13 16 9 13 7 13 1 10 9 0 9 7 9 2
14 11 13 16 11 11 13 9 2 16 11 13 11 2 2
19 1 9 9 2 11 2 11 12 2 11 2 7 11 2 11 11 2 13 2
54 11 14 13 13 9 1 9 9 9 15 13 1 11 11 2 9 9 0 1 11 11 2 9 0 2 0 1 9 11 11 11 2 9 0 2 0 1 9 11 7 11 7 9 9 13 9 0 1 9 9 15 13 9 2
13 11 11 10 13 9 1 3 1 12 9 9 0 2
14 1 9 3 2 9 3 13 9 0 1 9 9 11 2
102 16 1 9 1 13 1 9 9 2 9 9 2 9 11 2 9 9 2 7 9 9 2 3 13 9 2 9 1 11 11 11 11 2 13 2 9 12 9 2 12 2 2 9 12 9 2 12 2 7 13 2 12 2 2 9 9 9 2 12 2 2 9 12 2 7 9 11 11 2 11 9 11 11 11 11 12 2 1 9 0 11 11 11 11 11 7 11 11 11 13 2 13 2 11 2 11 1 11 11 11 11 2
4 3 9 0 2
9 11 11 7 11 13 1 9 12 2
26 11 13 1 13 12 11 12 1 9 9 1 11 11 11 1 11 11 1 9 9 15 3 9 9 11 2
22 11 13 9 9 9 9 11 7 10 0 13 2 13 15 0 2 0 7 15 14 13 2
33 11 9 1 9 3 13 1 9 1 12 9 1 11 11 7 10 9 1 11 11 3 9 9 11 2 11 11 11 11 11 5 11 2
38 1 9 9 9 9 11 11 10 14 3 13 1 0 1 9 15 13 16 13 1 9 15 14 0 7 9 9 15 0 13 1 13 7 13 9 11 11 2
14 11 11 3 13 12 9 1 2 7 3 13 12 9 2
5 9 9 13 11 2
18 0 10 9 9 9 13 9 2 9 9 2 9 2 9 9 7 9 2
16 7 9 12 15 13 9 11 11 9 11 2 11 11 11 11 2
21 3 3 2 15 9 12 13 1 11 1 9 10 7 1 0 13 1 10 9 0 2
39 16 3 2 9 10 13 9 15 3 0 13 1 9 9 0 1 11 11 11 11 7 11 11 11 2 16 14 3 0 1 9 9 0 1 9 12 3 11 2
43 11 0 0 13 1 9 9 0 11 11 11 2 9 12 2 11 13 9 15 3 0 1 0 0 1 9 13 11 11 12 2 11 2 15 0 1 11 15 13 1 9 9 2
3 0 9 2
22 9 9 9 0 1 12 9 0 2 11 2 11 2 7 11 2 3 3 13 12 12 2
34 9 13 2 1 9 13 9 9 1 0 2 7 9 15 13 9 13 1 9 9 2 13 1 9 11 2 2 1 13 9 9 7 9 2
42 1 9 11 9 10 13 1 9 2 9 9 9 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 7 0 2 0 2
43 1 9 9 11 0 2 11 2 11 3 13 9 15 3 3 0 2 12 11 12 2 12 2 12 2 9 2 2 16 1 3 9 3 9 3 13 2 3 16 9 3 13 2
32 11 3 13 1 9 9 2 11 2 2 13 9 2 2 15 3 13 1 9 9 1 9 1 11 2 16 13 9 0 1 9 2
43 11 2 9 1 9 13 9 16 13 1 9 9 9 2 7 9 3 2 3 15 3 13 10 9 3 13 9 0 2 7 1 9 7 1 9 15 13 1 9 1 9 15 2
26 11 13 7 13 1 11 7 11 2 16 11 2 13 1 9 2 9 2 13 1 13 7 11 3 13 2
22 1 9 15 0 2 16 11 11 11 13 1 10 9 2 15 3 13 9 1 9 10 2
21 1 9 12 11 12 2 11 11 13 1 9 11 11 2 16 3 13 1 9 12 2
20 13 1 11 11 2 7 13 1 11 11 11 1 9 11 1 11 7 1 11 2
17 11 11 2 2 13 10 9 2 9 2 9 2 7 9 13 11 2
16 11 7 11 11 1 0 13 9 9 10 9 1 12 7 12 2
20 9 1 2 9 2 13 2 9 2 3 13 1 9 9 2 7 1 9 11 2
25 9 2 9 11 12 9 13 11 1 9 12 16 11 9 11 13 9 0 1 9 2 9 1 13 2
19 11 9 13 1 9 9 9 7 9 1 9 9 2 9 9 2 7 9 2
16 16 13 9 0 1 9 10 2 11 3 13 1 9 11 12 2
17 10 9 13 9 1 9 9 9 11 7 10 9 3 13 9 9 2
9 15 13 11 9 1 9 7 9 2
15 3 2 3 15 10 13 9 15 0 7 13 9 7 14 2
36 16 1 9 9 9 12 13 12 7 3 9 0 3 13 9 9 2 16 9 9 10 13 13 9 9 9 15 13 1 13 12 9 11 3 13 2
40 9 11 11 13 13 1 9 9 7 1 13 11 11 11 11 2 15 13 1 11 11 11 1 10 11 5 11 7 13 1 9 9 7 9 1 11 11 11 11 2
37 11 3 13 10 9 0 15 13 1 9 15 0 15 14 3 13 1 13 9 0 10 1 1 9 1 13 9 9 1 9 9 0 10 15 3 0 2
22 11 11 13 10 9 1 11 15 13 9 9 12 12 2 7 9 12 9 2 12 2 2
11 11 1 9 12 2 13 9 1 12 9 2
22 16 1 13 9 10 9 2 11 2 11 13 10 9 1 3 13 7 3 13 9 0 2
21 1 9 15 13 1 9 9 2 9 10 13 1 9 0 1 13 9 1 9 10 2
14 16 2 1 11 11 2 9 9 9 0 13 9 10 2
28 3 9 7 10 2 3 1 9 12 11 12 11 11 13 13 9 11 1 9 9 0 2 9 2 9 9 0 2
8 13 9 1 9 2 9 0 2
45 11 9 1 0 13 9 9 0 2 11 2 2 7 16 11 11 3 13 9 7 9 1 9 9 2 13 3 9 9 9 2 7 7 16 1 11 10 3 13 9 0 2 11 2 2
15 11 11 13 9 9 12 2 7 9 3 13 1 11 12 2
8 11 0 13 9 7 9 9 2
16 16 13 9 1 9 9 11 7 11 2 11 13 1 9 9 2
26 1 12 11 12 2 11 13 9 12 1 11 1 9 12 2 12 1 11 11 1 9 11 11 11 12 2
8 11 11 11 13 1 11 11 2
20 11 11 11 7 11 11 2 2 13 9 9 9 1 9 1 9 0 1 11 2
11 11 10 9 10 11 1 9 9 13 9 2
5 15 3 11 11 2
14 1 12 11 13 13 1 11 11 11 11 2 11 2 2
32 1 9 12 15 1 13 13 1 13 13 1 9 9 11 9 12 2 12 2 1 9 9 2 13 1 11 11 2 1 9 0 2
44 11 13 9 10 9 9 1 11 2 11 15 13 1 9 12 11 12 15 9 10 13 1 11 11 2 9 2 2 11 2 11 2 2 11 2 11 2 2 7 11 2 11 2 2
34 16 10 9 13 16 9 3 13 9 15 13 15 13 9 1 9 0 2 13 9 2 9 7 9 0 2 1 9 2 9 9 7 9 2
10 16 9 10 13 1 9 1 9 11 2
87 11 11 11 2 11 2 7 9 11 11 1 14 3 3 13 13 1 1 9 9 11 11 1 11 2 11 11 12 3 13 1 9 11 11 3 13 15 10 9 2 7 3 3 13 1 10 9 1 9 11 2 1 3 2 9 11 1 11 2 12 2 2 9 11 1 11 2 12 2 2 9 11 2 12 2 7 11 2 12 2 7 9 11 2 12 2 2
16 11 11 14 3 13 1 11 2 16 3 1 9 9 1 11 2
16 1 11 2 15 13 1 10 10 9 15 3 13 1 9 10 2
10 9 10 3 13 12 9 1 9 12 2
21 16 3 2 11 3 13 9 9 1 11 1 13 1 9 11 11 3 13 1 11 2
11 3 10 9 3 13 9 1 13 9 10 2
16 11 1 12 9 15 13 9 2 9 13 9 13 1 9 9 2
8 3 11 13 11 7 11 3 2
10 9 3 15 3 13 1 9 9 15 2
14 12 9 13 2 13 1 12 9 2 1 12 9 9 2
38 1 9 9 11 1 9 9 2 12 5 12 9 12 11 12 1 9 9 13 9 2 16 1 9 10 11 11 9 3 13 11 11 11 9 11 11 11 2
54 9 11 11 11 3 13 13 11 11 2 11 2 7 11 2 0 9 1 9 0 1 11 2 11 14 14 13 1 9 9 9 2 3 1 9 12 11 12 13 9 9 15 13 13 10 9 11 2 3 1 9 11 11 2
16 1 9 2 9 11 10 2 10 9 13 1 9 10 2 10 2
11 9 10 13 9 1 13 9 1 9 12 2
8 15 13 10 9 7 12 9 2
16 3 10 11 11 3 13 1 9 11 11 2 13 11 11 11 2
17 10 9 13 1 11 11 11 2 7 9 13 11 11 7 11 11 2
10 9 10 3 13 7 13 0 7 0 2
13 1 9 12 2 9 10 13 9 9 0 12 9 2
21 9 12 11 7 11 12 11 1 11 13 10 9 1 9 11 1 11 1 11 11 2
10 9 10 13 12 9 1 9 9 11 2
8 11 11 3 13 9 9 9 2
115 9 9 9 13 11 11 11 15 3 13 9 2 9 1 10 9 9 11 5 11 2 11 11 11 7 9 9 13 1 11 5 11 1 7 1 9 11 11 11 1 11 11 2 11 11 11 11 13 1 9 9 1 0 9 9 2 11 11 11 13 11 11 11 15 3 13 1 9 9 11 7 11 11 11 11 3 13 1 10 9 3 13 9 11 5 11 2 11 14 3 13 1 9 9 9 16 3 13 11 1 13 9 1 10 9 15 0 1 9 9 9 11 13 0 2
8 9 10 13 13 1 9 12 2
24 9 10 13 9 9 9 9 2 9 2 11 2 9 15 13 9 1 9 0 2 9 2 9 2
16 11 9 3 13 0 1 9 7 1 11 0 1 9 11 11 2
17 3 12 9 0 10 13 13 9 9 13 11 2 3 13 11 2 2
19 2 7 10 11 13 1 15 10 9 1 9 11 2 2 11 11 11 11 2
34 16 11 3 13 1 9 2 9 15 3 0 13 9 9 15 2 3 2 3 1 9 3 1 12 9 2 1 1 11 11 2 11 2 2
25 1 11 11 13 1 9 1 11 11 12 2 9 13 9 0 11 1 12 9 0 1 9 2 9 2
90 11 11 11 15 13 1 11 2 9 1 12 9 1 12 9 0 3 11 11 2 11 11 7 11 13 12 9 3 11 1 11 2 9 9 1 11 2 9 9 1 11 11 2 9 9 9 1 11 2 9 9 11 1 11 7 9 9 1 11 11 13 9 1 10 9 9 9 0 1 9 2 11 11 2 13 13 9 15 0 2 0 13 1 9 9 13 0 13 9 2
35 7 1 9 11 11 11 2 11 11 2 2 11 11 13 11 15 3 13 7 13 9 15 3 13 1 9 11 15 11 11 13 9 1 11 2
18 9 9 1 9 9 11 11 9 9 0 13 9 9 9 7 9 11 2
14 11 13 9 11 7 11 1 11 12 1 11 1 9 2
8 9 10 3 13 1 9 12 2
19 1 9 9 9 9 2 9 0 13 1 13 9 9 7 13 9 9 9 2
49 9 9 9 10 13 1 11 11 2 16 9 9 9 15 13 1 9 9 9 13 1 10 10 9 9 0 15 13 1 9 2 9 9 9 11 2 11 12 2 11 11 12 2 12 11 11 12 2 2
4 3 15 13 2
23 3 3 10 9 9 15 3 13 9 1 1 9 9 2 9 2 9 2 9 0 7 9 2
12 9 0 10 12 9 13 11 1 12 9 12 2
19 9 11 13 3 0 13 9 0 9 15 14 3 13 10 9 1 9 9 2
26 1 9 10 3 13 9 11 15 12 9 2 16 3 1 12 7 12 15 13 1 11 11 7 11 11 2
28 11 10 13 9 0 9 0 15 13 1 9 1 12 1 12 9 9 0 2 3 9 2 9 2 9 7 9 2
32 11 13 1 0 2 15 13 9 9 11 2 13 15 1 9 15 2 13 1 9 2 9 11 2 7 13 9 15 15 13 11 2
45 3 13 1 9 9 7 9 2 11 11 2 13 9 2 2 11 11 2 11 11 2 2 13 1 9 2 9 11 2 1 11 11 11 2 7 0 11 11 2 9 11 11 11 2 2
32 1 9 0 2 9 9 3 13 3 0 16 15 13 9 15 13 10 0 15 3 13 16 9 13 1 9 1 2 9 1 9 2
42 1 1 9 9 11 2 9 11 1 11 13 2 16 9 13 13 9 9 9 2 1 0 13 11 2 11 2 11 2 2 11 2 11 2 11 2 7 11 2 11 2 2
20 9 9 0 11 11 13 10 9 9 0 15 13 1 11 11 2 11 2 11 2
14 9 11 11 14 13 1 11 7 9 2 9 11 11 2
10 9 12 11 13 1 1 9 11 11 2
12 11 3 13 9 15 13 9 9 13 14 0 2
28 11 15 13 9 2 16 13 1 13 10 9 2 9 12 9 9 15 13 1 10 9 2 1 9 2 1 9 2
5 0 9 9 10 2
57 11 13 2 11 11 2 10 9 15 13 1 9 1 9 15 3 13 2 15 3 2 3 14 3 13 2 7 1 9 15 3 13 1 0 2 16 9 15 3 3 13 2 9 9 2 2 9 10 13 9 2 9 0 1 9 9 2
18 11 10 13 9 0 15 13 9 15 13 9 11 2 7 3 13 9 2
10 9 15 3 13 1 9 2 7 13 2
15 11 13 9 1 11 11 2 11 11 2 11 11 2 11 2
19 11 11 11 11 13 9 11 15 13 1 9 12 1 13 1 11 2 11 2
13 11 0 11 11 13 10 0 3 15 3 13 11 2
37 1 11 2 9 11 1 9 2 9 9 12 11 12 13 9 9 15 10 7 10 0 9 13 1 9 1 9 1 0 15 13 1 9 9 15 13 2
24 12 9 3 13 2 13 2 7 3 13 1 13 9 1 9 9 0 15 9 13 1 11 11 2
23 13 1 10 9 1 11 11 11 16 9 10 2 13 9 1 0 1 10 9 9 11 2 2
14 11 13 9 2 9 2 9 9 2 7 9 9 9 2
32 9 10 10 14 9 1 9 11 11 2 7 9 9 15 13 1 9 10 15 13 10 9 2 9 15 3 13 9 0 9 10 2
31 11 9 12 13 2 2 1 9 9 11 10 2 16 10 9 9 2 9 15 1 9 0 13 11 2 13 14 0 3 2 2
21 1 9 10 11 11 11 13 9 1 9 11 11 11 15 13 1 9 12 11 12 2
2 3 2
56 9 0 10 13 1 11 1 10 9 0 2 7 13 1 9 9 0 9 9 9 0 15 3 13 11 2 3 9 1 9 13 1 2 11 11 2 7 11 11 2 2 7 13 13 15 3 0 1 9 2 9 9 9 0 10 2
7 9 9 9 10 13 12 2
41 9 11 2 13 9 15 13 1 11 11 11 16 13 1 9 9 7 9 7 16 9 11 13 1 9 11 11 2 15 13 9 11 1 9 11 11 11 1 9 9 2
13 14 13 9 15 3 13 9 9 1 0 2 14 2
28 11 11 7 3 13 9 9 1 9 11 13 10 9 9 0 15 13 1 9 9 11 2 11 11 11 2 11 2
15 10 0 3 13 1 9 13 7 9 9 2 9 9 2 2
31 16 9 10 9 13 9 11 2 16 9 9 9 10 2 16 9 11 13 1 13 1 0 9 11 15 0 1 10 9 0 2
24 3 9 0 15 13 1 11 2 3 1 12 2 12 9 0 2 11 11 13 9 1 9 11 2
12 3 3 13 9 14 13 2 1 9 0 13 2
33 11 11 11 10 0 13 1 9 11 7 13 10 9 13 1 9 11 2 10 0 15 13 1 9 11 10 13 1 9 11 7 11 2
24 9 2 9 15 3 0 9 3 13 13 1 9 15 13 1 10 9 7 13 9 15 3 0 2
25 16 11 14 13 9 9 13 11 2 7 7 13 10 9 0 15 13 1 11 11 2 1 11 13 2
17 9 9 15 2 9 9 2 9 0 9 2 9 13 7 11 11 2
11 3 9 11 11 3 13 1 9 9 11 2
15 1 11 2 11 13 13 11 2 7 11 13 13 9 11 2
13 9 0 9 9 11 11 1 0 9 12 2 12 2
10 7 11 2 11 11 2 9 0 11 2
36 11 11 11 11 11 1 0 13 9 15 3 13 1 9 2 1 3 12 9 9 1 9 9 2 11 15 13 2 10 13 1 9 9 11 11 2
20 11 11 13 10 10 11 15 13 1 11 9 2 11 11 2 11 11 2 11 2
18 1 9 9 13 11 11 7 15 3 13 1 11 11 2 11 11 2 2
38 11 13 9 0 1 9 12 1 9 12 9 11 11 1 11 11 2 15 13 9 1 10 9 7 13 2 13 1 9 9 9 0 1 9 9 9 11 2
11 11 2 11 2 11 13 10 9 1 11 2
14 11 13 9 1 11 11 2 11 11 2 11 2 9 2
18 9 9 10 13 15 12 1 11 2 12 1 11 7 15 12 1 9 2
18 3 9 10 13 9 11 11 7 3 10 9 0 15 13 9 11 11 2
12 9 15 13 13 9 9 15 0 1 9 0 2
72 3 11 11 11 2 9 9 11 11 13 9 2 12 5 2 2 9 12 2 12 9 2 12 5 2 2 9 12 2 12 9 2 12 5 2 2 11 11 2 11 2 12 5 2 2 11 11 2 12 5 2 2 11 11 2 12 5 2 2 9 11 2 12 5 2 7 11 2 12 5 2 2
18 10 2 10 9 13 13 1 10 9 16 15 13 7 13 1 10 9 2
12 11 3 13 1 10 9 2 7 3 13 9 2
12 1 9 11 2 11 11 1 0 13 13 11 2
14 16 10 1 11 2 15 13 13 5 13 10 9 9 2
15 16 10 9 13 13 7 11 13 13 2 9 1 9 0 2
10 9 10 13 12 11 11 2 13 11 11
15 3 15 9 9 13 9 15 0 13 9 10 13 1 15 2
13 1 9 2 9 0 15 13 9 0 7 13 9 2
18 10 0 11 13 0 1 9 1 9 9 7 0 1 11 0 7 0 2
2 3 2
11 11 11 2 13 10 9 9 1 9 9 2
10 11 3 13 1 13 9 7 9 9 2
9 16 13 2 16 9 11 3 13 2
21 9 9 11 13 1 9 9 7 9 11 2 11 11 2 9 9 10 13 9 0 2
16 9 13 1 10 10 9 9 9 9 11 11 2 11 11 11 2
22 1 1 9 13 13 12 9 2 7 11 2 11 11 2 11 2 9 9 9 11 11 2
13 11 11 13 10 9 1 11 11 2 11 2 11 2
12 9 10 3 2 3 13 9 9 15 13 9 2
15 11 11 13 10 9 1 11 11 2 11 11 11 2 11 2
12 7 11 7 11 2 9 11 2 13 9 15 2
29 1 9 9 2 9 2 9 15 13 1 13 9 13 0 2 3 10 9 13 9 9 15 13 2 1 13 1 9 2
22 11 11 13 1 11 11 11 11 11 11 1 9 12 2 16 9 11 11 13 9 10 2
7 2 3 9 14 3 13 2
11 11 1 11 0 9 13 1 12 11 12 2
15 15 3 13 9 1 13 9 11 1 13 15 16 14 13 2
50 1 9 9 0 12 2 13 1 9 0 12 2 5 2 2 15 9 13 12 9 9 9 2 9 1 9 0 12 1 9 11 2 11 11 13 12 9 1 9 11 2 16 11 9 0 7 9 9 0 2
5 9 13 1 11 2
16 11 13 10 9 1 9 11 2 9 9 11 2 11 2 11 2
51 1 9 9 11 11 13 10 9 15 13 9 11 11 5 9 11 1 11 11 15 13 2 11 11 11 11 2 1 9 9 9 11 11 1 13 9 7 9 13 1 12 9 9 9 15 13 1 9 9 9 2
16 1 10 2 13 3 1 9 1 10 9 9 1 9 1 11 2
20 9 10 13 1 9 12 2 12 9 9 11 11 1 11 11 2 9 12 2 2
13 11 11 12 13 1 12 9 15 13 1 12 9 2
29 11 11 11 2 11 11 2 11 11 2 7 11 2 11 11 13 9 11 11 9 12 15 13 1 11 11 2 11 2
13 11 11 13 10 9 9 15 13 1 11 2 11 2
21 1 10 2 1 9 9 9 11 3 13 1 15 3 0 1 9 10 9 15 13 2
18 1 9 2 11 13 1 9 9 9 11 11 11 2 3 11 7 11 2
11 1 0 2 9 13 1 9 9 10 9 2
10 9 10 13 9 1 12 11 12 9 2
31 1 9 10 13 9 9 15 3 13 2 11 11 2 2 9 10 13 11 11 1 9 7 11 11 2 9 11 2 1 9 2
16 11 13 9 1 11 11 2 11 11 2 11 11 11 2 11 2
11 15 13 9 0 1 11 0 13 9 9 2
7 9 0 13 13 9 10 2
45 1 10 3 9 9 10 3 13 16 13 9 15 0 2 16 3 13 3 3 2 3 9 15 3 13 16 9 9 7 9 9 2 7 3 3 13 9 0 1 13 7 13 1 0 2
19 11 11 13 10 9 15 13 1 11 11 11 2 11 11 2 11 2 11 2
43 11 13 9 1 9 11 9 12 2 11 2 11 2 11 2 2 2 16 9 9 0 1 11 11 11 2 11 11 3 13 1 9 11 11 2 11 11 11 11 11 11 2 2
20 9 9 2 9 9 2 13 9 9 1 9 9 13 9 9 1 9 1 9 2
17 9 10 13 9 1 11 11 10 2 12 1 9 9 11 1 11 2
9 3 15 13 9 0 9 11 11 2
6 13 1 11 2 11 2
16 9 0 2 11 9 11 11 11 11 2 11 9 0 2 11 11
7 13 9 12 1 12 9 2
41 9 9 13 1 9 9 2 9 2 9 0 15 13 9 1 9 2 1 13 1 9 2 16 9 0 13 1 9 9 2 9 2 9 0 15 13 9 13 9 2 2
17 3 1 9 9 9 10 2 1 9 3 9 13 9 15 0 10 2
15 16 3 9 10 13 9 9 1 1 9 7 9 15 3 2
18 11 0 9 10 13 9 9 11 11 11 2 11 2 11 2 11 2 2
30 9 10 13 1 0 1 13 10 9 7 9 2 13 9 15 13 9 2 13 10 9 9 2 7 13 9 11 11 11 2
25 11 11 11 11 11 13 1 9 10 1 9 12 2 7 1 9 12 9 1 11 13 1 11 11 2
9 1 12 12 9 2 15 13 13 2
44 16 13 3 0 2 11 13 9 9 12 12 1 11 12 2 11 13 1 11 2 11 2 11 2 11 0 1 9 11 11 2 11 11 11 2 15 3 13 12 9 1 9 12 2
25 9 10 13 9 0 9 9 1 11 1 9 12 7 13 1 11 2 9 15 3 0 1 9 9 2
19 15 13 9 9 15 13 1 11 11 2 11 11 2 11 2 7 11 11 2
28 3 2 11 3 13 15 1 9 9 1 11 2 11 2 7 13 1 9 9 0 1 13 9 15 13 1 9 2
15 10 9 10 3 13 1 9 11 7 13 1 13 9 9 2
7 3 9 9 11 7 11 2
18 11 13 9 9 0 15 9 13 13 9 2 12 1 9 9 9 9 2
16 9 13 1 9 11 12 9 1 11 11 11 2 11 11 2 2
24 11 13 9 9 9 11 11 7 13 9 9 15 13 1 0 15 3 3 13 1 11 7 11 2
28 16 13 15 13 11 11 1 11 11 2 11 11 11 2 11 11 11 11 2 11 11 11 2 7 11 11 11 2
14 13 1 3 0 1 9 0 7 1 13 1 13 9 2
30 11 11 2 11 11 2 12 11 12 2 12 11 12 2 13 10 9 2 0 2 0 2 7 9 1 9 0 1 11 2
14 11 11 13 12 9 3 2 11 2 11 2 7 11 2
13 11 13 10 10 9 9 15 13 9 9 15 13 2
29 3 11 11 13 12 9 7 12 9 9 2 15 9 10 9 13 0 1 10 11 2 13 11 2 11 2 7 11 2
34 15 13 13 2 13 1 11 2 11 11 2 11 2 10 11 15 3 13 11 7 13 13 1 1 11 2 1 9 0 1 13 10 9 2
17 1 9 12 2 1 11 7 11 13 11 2 11 11 11 11 2 2
16 16 9 0 3 13 2 7 9 10 9 10 9 0 2 2 2
16 11 3 13 1 9 1 11 2 11 3 13 1 9 9 13 2
34 10 9 10 13 11 1 12 11 12 1 9 0 11 15 0 2 11 11 11 11 2 13 1 11 11 11 7 10 9 2 11 11 11 2
35 9 10 13 9 11 1 2 0 1 11 1 11 1 9 2 9 9 1 11 10 13 1 9 12 9 9 2 13 1 9 11 1 9 12 2
19 14 11 2 9 9 10 2 16 11 13 2 7 9 9 2 16 11 13 2
12 11 11 13 11 2 11 15 13 1 9 11 2
25 1 9 0 1 9 10 2 9 13 9 10 1 9 0 1 13 9 1 9 1 13 1 9 9 2
8 11 2 9 13 1 9 12 2
9 9 0 9 1 9 10 13 11 2
19 11 13 10 10 9 1 11 11 11 11 2 11 11 2 11 11 2 11 2
41 11 1 9 10 13 1 1 12 7 12 2 12 15 3 13 12 9 9 1 15 0 2 3 11 2 1 9 12 2 7 12 2 12 2 7 11 12 2 12 2 2
7 11 12 13 1 9 12 2
18 1 10 9 7 9 2 9 13 9 15 14 0 2 0 2 1 9 2
14 11 11 2 11 13 9 15 13 1 11 11 2 11 2
10 11 13 13 11 7 3 13 9 0 2
21 14 9 1 9 9 7 9 11 11 13 11 11 10 13 9 11 15 13 1 11 2
12 9 0 15 3 13 1 9 3 13 1 9 2
11 11 11 3 0 7 13 2 3 9 13 2
9 11 9 13 9 0 9 9 10 2
11 11 3 13 1 9 11 11 1 9 12 2
8 9 11 1 9 10 13 11 2
15 1 9 12 2 9 11 13 12 9 11 16 14 13 9 2
10 11 10 3 13 1 9 15 3 0 2
45 9 9 9 13 9 1 9 9 1 14 2 3 0 2 12 0 0 2 7 13 3 13 9 1 2 9 2 9 2 7 9 10 3 13 1 9 9 15 13 9 2 9 10 9 2
7 16 15 3 13 1 11 2
7 0 13 9 3 3 0 2
10 11 2 14 11 2 3 11 13 15 2
10 15 13 9 0 1 13 9 9 10 2
9 16 15 13 13 9 10 9 9 2
16 13 1 9 9 0 2 9 10 13 9 9 0 12 9 11 2
33 11 2 9 13 1 13 9 9 10 3 13 1 9 11 1 2 9 9 2 2 11 11 2 2 7 13 1 9 11 1 11 11 2
31 16 2 11 2 15 13 3 14 13 1 9 0 1 9 10 9 0 2 9 10 3 13 1 9 11 1 13 1 9 11 2
23 15 13 9 1 13 9 7 13 9 1 1 9 2 1 13 9 1 9 9 15 0 2 2
14 2 11 11 2 3 15 13 9 15 3 15 13 9 2
9 1 12 9 10 13 2 11 2 2
5 9 9 1 11 2
11 9 10 13 9 0 11 11 7 11 11 2
15 11 13 10 9 1 9 9 11 2 11 11 2 11 11 2
24 1 0 9 2 15 13 9 11 13 9 0 11 11 7 13 9 2 9 0 7 9 2 0 2
18 16 2 11 11 15 15 13 13 10 10 15 13 3 1 11 7 11 2
8 11 11 11 13 3 9 13 2
4 2 2 2 2
21 16 16 9 0 9 9 14 13 2 9 2 9 2 15 13 9 9 10 3 13 2
24 11 11 13 10 9 9 0 11 11 2 13 1 11 11 11 2 11 7 9 11 11 11 11 2
16 9 9 10 13 11 2 11 13 9 0 9 11 2 1 11 2
19 11 13 10 10 9 1 11 11 2 11 11 11 2 11 11 11 2 11 2
37 9 10 2 13 1 11 11 13 10 9 1 12 9 2 9 3 2 3 12 5 2 1 9 13 1 12 1 12 5 7 1 9 3 1 12 9 2
10 11 11 11 13 1 9 1 12 5 2
32 1 9 9 9 2 1 9 9 9 15 13 1 9 2 9 13 1 9 9 9 2 9 15 13 9 13 9 1 9 9 2 2
24 1 13 9 11 11 2 11 3 3 13 10 9 0 11 11 1 9 9 15 13 1 9 9 2
34 9 9 9 0 1 9 12 13 1 9 9 15 13 12 9 7 1 9 11 15 13 12 9 1 9 9 9 3 2 3 12 7 12 2
24 13 1 9 2 9 0 2 13 1 9 0 1 1 9 9 2 13 7 1 9 2 9 0 2
15 9 11 3 3 0 2 16 13 9 1 9 11 7 9 2
9 15 13 11 11 11 2 12 2 2
32 1 3 13 9 9 7 9 1 1 13 9 1 9 9 9 2 9 9 15 0 2 7 9 9 0 2 0 13 15 1 13 2
12 1 9 12 2 9 10 13 9 1 12 9 2
24 9 9 15 3 13 9 9 9 0 9 1 9 9 9 11 0 13 9 15 13 1 9 11 2
25 1 9 11 12 2 9 11 13 1 11 2 11 2 11 7 14 3 3 13 3 1 11 2 11 2
6 15 13 11 13 9 2
16 12 9 9 16 11 7 11 3 9 10 13 1 9 9 9 2
12 3 3 15 14 13 9 7 9 9 0 15 2
17 9 10 13 1 0 1 9 9 2 16 3 0 9 7 3 13 2
10 11 11 13 9 0 16 11 11 11 2
23 11 11 13 10 10 9 15 13 1 11 11 2 9 11 11 11 2 11 11 11 2 11 2
13 11 11 13 10 9 1 11 15 13 9 1 11 2
17 11 2 9 9 9 11 15 3 13 13 11 11 11 9 11 11 2
27 12 9 13 13 9 0 12 12 2 12 1 2 1 12 12 9 9 2 15 13 0 9 9 9 1 9 2
12 3 11 13 9 11 1 11 11 1 9 12 2
22 11 11 11 13 10 10 9 15 13 1 11 11 2 11 11 11 2 11 11 2 11 2
21 9 1 9 0 3 13 1 9 7 9 2 1 3 2 3 13 12 5 9 9 2
30 16 1 9 10 0 2 11 9 10 13 1 11 13 9 2 13 9 1 9 2 9 2 3 15 13 9 7 13 1 2
39 11 11 13 1 9 12 2 1 12 9 13 13 11 11 7 1 9 0 3 13 11 11 2 9 2 11 13 0 9 1 9 1 9 1 9 11 2 11 2
48 1 9 2 9 9 15 13 9 2 16 3 9 9 13 1 9 15 0 13 9 7 13 10 10 9 9 1 11 1 13 2 11 2 1 1 9 9 9 2 11 2 1 11 2 11 7 11 2
22 11 11 13 10 10 9 15 13 1 11 11 2 9 11 11 2 11 11 11 2 11 2
35 9 1 9 9 13 1 0 1 9 11 11 7 11 1 9 7 1 9 9 12 15 13 1 3 9 1 9 2 9 1 13 9 11 11 2
22 9 2 9 1 9 1 9 0 1 9 9 9 0 15 14 3 13 9 2 9 2 2
23 1 12 11 12 2 11 11 11 7 11 11 13 9 9 2 15 13 9 1 9 9 10 2
21 9 10 3 0 1 9 15 13 3 10 0 2 9 0 15 14 0 1 11 11 2
8 15 13 9 12 1 12 9 2
6 11 9 10 13 0 2
34 1 13 9 11 2 11 11 2 9 16 11 1 10 2 10 9 5 9 9 3 13 9 1 0 2 9 11 2 3 14 13 11 11 2
16 9 10 3 13 9 2 13 2 7 9 9 9 15 3 0 2
9 9 10 3 13 9 12 2 12 2
36 11 11 3 13 12 9 0 2 3 11 11 1 11 11 2 11 11 1 11 11 2 11 11 1 11 11 2 11 11 11 2 7 11 11 11 2
24 9 9 15 0 13 9 9 2 9 13 10 9 2 7 9 15 3 0 1 11 9 2 12 2
20 1 12 11 12 2 11 13 3 13 9 1 11 1 9 11 14 13 9 10 2
12 3 10 9 0 2 16 11 2 11 2 13 2
9 16 9 12 13 9 0 11 11 2
14 3 13 1 12 9 1 9 0 1 9 9 9 11 2
13 11 11 13 10 9 9 11 15 13 1 9 12 2
23 9 13 7 13 9 9 2 9 9 15 3 0 1 9 2 9 15 15 13 1 11 12 2
26 11 2 11 2 11 2 11 11 11 11 11 11 11 2 11 11 11 13 9 9 9 11 11 11 11 2
17 11 9 10 13 10 11 7 9 0 15 13 13 13 9 11 11 2
55 10 10 9 2 2 11 11 11 11 2 13 1 1 9 9 15 3 13 1 9 11 11 11 2 1 11 11 12 2 9 2 11 11 11 11 11 2 13 1 9 12 1 9 9 11 1 13 9 9 12 1 12 9 12 2
24 1 9 0 2 9 10 13 9 9 9 2 11 2 9 9 11 11 7 9 9 11 11 11 2
20 1 9 9 11 2 3 11 2 11 13 1 9 0 7 3 13 9 1 11 2
25 11 11 13 10 10 9 15 13 1 11 11 2 11 11 11 2 11 11 11 2 11 11 2 11 2
13 11 11 2 2 13 10 9 0 9 9 1 11 2
21 11 13 9 11 11 15 13 0 9 11 1 11 2 1 12 5 1 0 11 2 2
34 10 9 9 0 11 3 9 3 13 1 10 9 1 9 11 2 11 11 15 0 1 9 2 9 2 7 9 3 13 1 11 7 11 2
22 11 11 11 11 13 1 9 12 11 12 1 11 11 2 10 9 1 11 2 9 11 2
15 11 3 13 1 9 2 9 1 13 13 9 2 9 0 2
15 9 11 13 13 1 9 9 15 13 9 10 9 9 11 2
10 9 9 13 3 9 9 1 13 9 2
33 1 9 12 2 11 11 11 11 11 2 3 13 1 9 12 9 9 2 7 0 12 3 13 1 0 1 12 9 9 1 9 12 2
21 1 13 9 15 3 0 2 9 10 9 2 7 9 2 9 10 14 0 13 9 2
17 16 11 13 1 11 2 3 13 11 0 1 0 13 9 1 11 2
11 9 10 3 13 3 1 9 9 9 11 2
39 9 3 13 1 11 11 11 11 1 9 12 11 12 7 13 1 12 9 3 11 2 11 2 11 2 11 2 11 2 11 7 11 1 12 9 9 13 9 2
9 9 0 13 1 9 12 11 12 2
25 1 12 2 9 11 11 13 2 1 12 12 2 9 11 7 9 2 9 15 13 13 1 11 13 2
29 1 9 9 11 11 12 11 2 11 11 11 2 15 13 12 11 12 2 15 13 9 9 1 11 11 7 11 11 2
28 11 2 9 1 9 11 11 13 9 2 9 9 0 11 2 1 1 9 2 11 13 9 2 15 13 11 11 2
18 9 0 10 13 1 0 16 15 13 11 11 1 11 11 1 11 11 2
32 11 11 11 2 9 11 2 11 11 11 2 2 12 11 12 2 12 11 12 2 13 11 11 12 1 9 12 1 13 1 12 2
14 11 9 9 13 7 9 10 13 1 2 11 11 2 2
25 1 1 9 10 1 9 2 13 10 9 7 0 0 9 15 14 3 13 1 11 11 7 9 11 2
38 11 2 9 9 2 9 11 13 2 1 1 9 11 2 11 2 1 9 11 2 11 11 15 13 13 9 11 2 10 9 9 3 13 12 9 15 0 2
24 1 9 11 2 11 11 2 2 10 9 11 13 0 2 15 3 13 1 9 15 0 3 0 2
32 11 3 13 1 9 9 11 11 11 1 13 9 11 2 12 2 1 9 9 1 0 2 2 11 2 7 2 11 11 11 2 2
15 11 3 13 9 13 11 11 7 13 11 11 1 9 12 2
84 9 10 13 9 9 15 0 7 9 0 7 0 1 9 1 11 11 11 2 13 1 9 11 11 7 11 11 2 9 9 2 11 2 3 13 9 9 9 2 16 11 11 11 7 11 1 11 2 11 11 11 1 11 7 9 0 1 11 2 7 11 11 7 11 11 11 2 11 3 13 9 0 9 9 1 9 9 0 0 11 2 11 11 2
35 13 9 2 9 2 9 9 15 0 9 13 9 2 9 11 15 13 1 9 10 13 16 15 15 14 3 13 1 0 16 9 10 14 13 2
8 11 2 15 3 13 1 9 2
17 11 13 9 15 13 1 9 11 2 11 11 2 11 11 2 11 2
8 11 9 0 9 9 1 9 12
10 9 11 11 10 13 9 15 13 11 2
8 11 2 11 2 7 11 11 2
19 16 9 10 13 10 9 1 9 15 1 13 9 2 9 15 13 11 11 2
8 11 13 9 15 0 1 9 2
6 9 15 3 15 13 2
12 11 13 9 11 11 0 13 12 11 12 9 2
40 1 9 12 2 11 9 1 11 2 11 11 11 11 11 11 13 9 15 13 10 9 0 1 9 10 2 9 9 7 9 9 15 13 1 11 11 1 9 10 2
15 11 2 11 2 11 13 9 1 9 11 1 9 9 11 2
6 9 9 3 1 10 2
17 14 11 3 13 16 11 11 2 9 10 3 13 12 12 12 9 2
24 9 9 15 0 3 13 11 13 1 11 2 1 11 11 13 13 9 1 0 9 0 11 11 2
18 9 2 11 3 13 9 11 2 16 15 3 13 1 9 9 15 0 2
32 1 9 1 11 2 1 0 13 1 9 12 9 2 12 2 11 2 11 11 12 1 10 9 1 9 9 13 13 9 2 9 2
26 1 9 2 9 10 13 9 7 9 9 15 0 1 9 9 2 1 9 9 9 7 9 15 3 0 2
15 11 11 2 15 13 1 12 9 7 1 9 13 12 9 2
6 11 14 13 9 0 2
31 1 11 11 11 2 11 13 16 15 13 9 3 3 1 10 9 11 11 2 7 3 9 9 7 9 7 3 9 15 13 2
18 16 9 11 3 0 1 12 11 5 11 11 2 9 3 13 1 9 2
27 3 13 9 9 12 9 2 9 9 10 3 13 12 10 9 9 1 10 9 15 12 1 1 13 9 0 2
12 0 11 10 2 9 2 7 2 9 2 11 2
21 11 11 13 10 10 9 15 13 1 11 11 11 2 11 11 2 11 11 2 11 2
44 9 10 13 9 12 16 3 2 3 13 1 9 7 9 13 9 13 2 2 11 3 13 9 13 0 11 12 9 12 2 7 3 11 11 2 11 2 9 13 0 0 9 12 2
27 11 13 9 15 13 1 3 13 2 3 13 1 9 1 9 9 2 9 9 9 2 7 1 9 2 9 2
21 11 10 13 12 1 12 9 7 9 15 13 1 11 11 2 11 10 13 9 12 2
12 16 14 3 13 9 2 3 15 13 9 9 2
15 11 15 13 9 11 2 13 13 9 16 11 13 13 9 2
16 1 13 2 9 3 3 13 16 15 13 7 3 3 13 13 2
24 9 11 11 2 11 11 2 1 9 13 3 13 1 9 9 12 2 12 2 3 0 1 11 2
16 16 1 10 9 11 2 15 3 13 9 2 9 11 15 0 2
21 14 3 0 1 11 5 11 11 11 2 13 3 9 9 9 7 11 3 11 11 2
24 11 11 11 11 2 2 13 10 10 11 9 1 11 11 2 11 11 2 11 11 2 11 2 2
4 15 13 0 2
19 15 13 13 1 13 1 2 11 11 2 2 11 11 2 11 7 11 2 2
25 9 9 3 13 9 0 15 13 9 3 13 2 13 2 13 9 9 9 2 9 15 13 2 13 2
12 9 15 13 9 13 3 3 11 1 9 9 2
11 9 9 0 13 1 9 9 0 15 0 2
5 9 10 1 9 2
31 11 0 13 9 9 9 1 11 11 11 11 3 11 11 11 11 2 9 2 11 11 11 11 2 11 11 13 9 9 10 2
19 11 11 11 10 13 9 16 13 1 9 9 15 13 1 9 9 7 9 2
29 9 9 1 9 11 13 9 2 9 9 9 1 9 10 1 9 9 9 1 9 9 12 2 12 1 12 2 12 2
38 10 9 11 11 3 13 9 13 11 15 13 1 11 11 11 2 9 11 7 11 2 9 9 1 9 0 2 1 11 11 11 2 3 13 9 9 10 2
20 11 11 13 10 10 9 1 11 11 2 11 11 11 2 11 11 11 2 11 2
35 1 13 9 9 3 9 15 3 0 2 11 11 9 13 11 11 2 9 9 0 10 2 13 1 9 9 1 9 0 2 13 13 1 12 2
8 9 10 13 11 11 11 11 2
37 1 9 9 12 2 11 11 3 9 1 9 9 9 1 9 11 11 11 11 1 13 9 9 9 15 9 14 9 1 9 12 11 12 2 9 2 2
11 11 13 1 13 1 13 0 1 11 11 2
15 1 9 9 1 9 9 2 11 13 13 13 9 13 11 2
20 16 11 11 13 0 2 15 14 3 13 10 10 9 2 16 11 11 1 13 2
36 9 3 0 7 0 12 1 11 11 11 11 11 11 1 9 9 9 9 12 13 2 11 11 5 12 11 2 11 5 12 11 2 9 9 12 2
23 11 11 13 10 10 9 15 13 1 9 9 11 2 9 11 2 11 11 2 11 2 11 2
25 1 11 11 11 12 5 12 2 11 13 3 13 11 11 1 13 9 16 13 11 11 1 9 12 2
8 9 10 13 9 1 12 9 2
70 11 2 1 9 12 9 1 11 2 13 9 0 1 11 11 9 2 11 11 2 11 11 2 10 9 0 1 9 2 1 15 15 13 9 0 2 16 11 11 2 11 7 10 11 11 2 2 11 11 2 10 9 0 1 11 2 2 1 11 11 11 2 7 11 11 1 9 1 12 2
26 13 9 0 15 13 1 9 1 9 9 9 2 11 11 11 2 2 15 3 2 3 13 1 9 9 2
7 15 0 7 13 1 11 2
14 11 13 9 1 11 11 2 11 2 11 11 2 11 2
15 11 13 7 13 13 10 9 1 9 9 2 3 11 11 2
19 11 13 9 15 13 1 9 11 2 11 11 11 2 11 11 11 2 11 2
22 11 11 11 2 2 13 9 9 9 13 9 12 5 1 11 15 13 1 9 11 11 2
18 11 2 2 13 9 11 7 9 1 9 11 2 11 2 11 2 9 2
14 11 11 11 11 13 11 11 11 12 15 13 1 12 2
19 11 11 3 13 9 1 12 9 2 16 9 9 3 3 13 12 3 12 2
29 1 11 1 9 10 9 3 13 9 1 13 1 9 2 9 0 1 11 11 2 11 11 2 11 11 7 11 11 2
5 9 9 13 12 2
26 9 10 3 13 16 9 15 13 1 0 1 9 9 9 1 9 1 9 0 3 13 13 9 9 11 2
17 11 13 1 9 11 7 13 9 2 9 1 9 9 1 12 9 2
20 9 9 7 9 9 13 10 10 9 9 1 9 9 15 13 1 3 7 0 2
9 9 10 13 12 5 1 9 0 2
15 11 11 13 9 1 11 11 2 11 2 11 11 2 11 2
21 1 9 9 0 7 9 9 2 9 10 13 1 9 0 1 9 11 2 11 2 2
13 9 10 13 1 11 11 15 14 0 13 11 11 2
16 7 3 9 9 1 11 2 14 11 7 11 7 10 9 11 2
36 9 0 13 9 0 9 3 9 9 2 14 3 13 9 2 16 9 9 2 9 13 9 1 9 2 9 15 13 7 9 1 9 7 9 0 2
23 11 11 3 13 9 7 9 9 1 12 9 1 10 9 1 11 11 16 13 11 11 11 2
12 3 9 9 1 10 9 13 16 13 9 9 2
49 10 9 2 9 0 9 9 1 9 0 13 9 9 2 13 1 9 10 2 11 3 3 13 9 7 9 0 16 3 13 9 10 2 13 13 9 2 9 0 2 3 13 1 9 2 9 9 0 2
16 9 11 11 13 14 0 1 9 9 11 15 0 2 11 11 2
44 9 9 11 11 1 11 2 7 9 16 15 13 9 9 2 9 0 2 7 9 0 13 1 10 9 1 12 9 2 16 9 11 9 9 7 9 13 3 3 16 13 11 11 2
25 11 12 11 13 9 9 9 11 11 1 11 2 11 2 1 9 13 9 9 9 11 11 9 12 2
13 9 2 9 11 13 9 9 9 15 0 7 0 2
26 11 11 3 13 9 0 9 15 13 10 9 1 9 12 11 13 1 9 11 11 11 11 7 11 11 2
36 16 13 11 11 11 11 11 11 11 3 3 13 12 5 1 9 9 1 9 9 12 5 12 7 3 13 13 12 5 1 9 9 12 5 12 2
33 1 9 11 12 2 9 11 13 12 9 7 9 11 11 2 9 13 12 9 2 1 9 12 2 11 11 13 1 9 9 0 9 2
28 9 15 13 2 11 11 11 11 11 11 2 15 13 1 1 9 11 11 2 13 1 11 1 13 11 11 15 2
12 11 13 9 9 0 1 9 9 11 2 11 2
9 16 2 9 9 0 13 1 0 2
17 9 9 0 15 13 11 2 12 13 11 11 11 1 12 11 12 2
25 16 11 13 9 10 9 11 1 11 1 13 9 1 9 11 2 11 13 13 9 9 2 9 10 2
8 11 13 1 9 15 14 0 2
20 16 11 1 12 7 11 1 9 12 11 12 2 16 13 9 0 11 11 11 2
14 11 13 9 1 11 11 2 11 11 2 11 2 11 2
16 16 13 1 9 2 11 7 9 13 9 9 1 9 15 0 2
42 1 9 9 2 11 11 13 9 11 11 13 9 9 5 9 15 3 13 10 10 2 13 10 10 9 1 9 11 11 2 2 1 9 1 9 16 14 3 13 11 11 2
23 11 15 13 13 9 7 9 9 9 1 9 9 2 11 2 11 11 11 11 11 11 2 2
12 1 11 14 1 13 9 10 13 9 10 9 2
8 7 3 3 15 3 15 13 2
59 1 9 12 2 11 13 1 9 9 9 11 11 2 15 10 9 3 13 9 9 1 9 11 11 11 11 2 12 2 2 13 1 9 11 11 11 2 1 9 12 2 11 11 13 9 11 11 2 10 9 11 11 11 1 9 11 11 11 2
30 1 1 9 11 11 0 2 11 11 11 5 11 11 13 10 9 11 2 1 11 11 2 11 11 2 11 2 7 9 2
14 9 3 13 9 2 15 3 2 3 13 12 9 9 2
16 1 9 11 2 11 13 11 10 9 9 7 13 9 13 11 2
9 11 13 10 9 9 15 3 13 2
41 11 9 9 11 13 15 0 2 7 16 13 9 9 9 11 2 11 2 11 11 2 2 11 2 11 2 11 11 2 2 7 9 9 0 11 2 11 2 11 2 2
20 9 10 13 9 15 3 0 15 13 11 11 2 11 1 0 12 7 12 9 2
7 9 15 3 13 1 11 2
12 9 10 13 9 0 15 13 10 9 1 9 2
31 1 9 2 12 1 12 9 9 15 13 10 3 13 1 9 11 1 9 9 9 9 11 15 12 2 12 1 12 11 12 2
8 15 9 15 13 9 0 11 2
34 1 9 1 9 13 12 9 1 9 9 7 9 7 12 9 1 9 9 1 9 9 9 9 2 9 11 11 2 11 11 7 9 9 2
23 11 9 13 9 10 1 10 9 2 9 2 9 9 2 9 9 9 2 7 10 9 9 2
12 10 9 10 2 10 13 12 9 1 12 9 2
16 9 9 16 15 13 15 9 11 13 16 15 13 10 9 9 2
16 11 9 10 13 1 9 9 9 15 3 3 13 9 0 11 2
4 3 15 13 2
13 11 11 11 2 2 2 13 9 9 9 1 11 2
12 0 9 9 9 13 1 10 9 1 9 0 2
29 9 10 3 13 16 1 9 15 13 11 2 15 13 16 1 9 2 9 13 2 9 2 9 15 13 3 3 13 2
14 3 13 1 13 9 1 9 9 15 13 13 1 9 2
7 11 3 13 9 10 11 2
4 15 1 11 2
11 11 13 10 1 11 2 11 2 11 11 2
