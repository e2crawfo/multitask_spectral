799 17
6 11 13 10 0 9 2
9 15 13 9 10 15 9 14 13 2
9 15 13 1 15 9 1 10 9 2
13 1 10 12 9 13 15 10 0 9 1 10 9 2
4 15 13 0 2
16 3 15 9 13 3 0 9 2 15 4 15 3 3 3 13 2
23 7 15 0 13 16 10 9 14 3 1 10 9 13 7 3 1 15 9 1 10 9 13 2
7 15 13 15 3 3 0 2
15 7 9 7 9 2 15 13 0 1 10 9 7 10 9 2
7 4 10 0 9 3 13 2
3 0 9 2
3 0 9 2
15 3 1 10 0 9 1 11 11 2 15 4 15 3 13 2
19 12 9 9 1 10 9 1 10 11 11 1 10 0 9 1 10 11 11 2
15 15 13 0 9 7 10 9 10 9 1 15 9 13 0 2
19 15 1 9 13 15 9 1 9 7 9 10 9 7 4 15 1 9 13 2
10 9 2 9 2 0 9 7 0 9 2
6 15 4 15 14 13 2
8 4 3 9 7 9 3 13 2
8 15 4 15 9 3 3 13 2
17 16 15 3 0 7 0 1 9 13 4 15 1 11 3 14 13 2
9 0 9 4 15 10 15 9 13 2
22 15 13 15 2 15 9 13 1 15 9 0 2 3 13 15 0 9 1 10 0 9 2
9 3 12 11 4 3 10 9 13 2
13 15 13 1 10 9 3 7 10 0 9 1 15 2
15 15 4 3 13 2 16 15 15 14 3 1 10 9 13 2
12 3 10 3 0 9 7 10 0 9 4 13 2
7 10 9 13 0 7 0 2
16 1 10 11 12 4 15 10 9 1 10 12 2 15 9 13 2
6 10 9 13 3 0 2
15 15 13 10 0 9 1 9 2 13 15 1 9 3 13 2
9 3 2 4 2 15 3 3 13 2
14 15 13 10 0 9 1 0 9 2 9 1 9 1 2
11 15 9 4 15 9 3 14 3 13 4 2
11 10 9 10 0 9 13 3 0 7 0 2
16 15 13 1 15 1 10 9 1 7 15 9 4 3 14 13 2
18 10 9 13 3 1 2 15 1 9 1 10 9 1 10 9 14 13 2
12 1 12 11 13 15 1 15 3 15 0 9 2
14 10 9 13 3 1 10 9 3 2 12 2 2 11 2
10 1 0 9 13 3 15 9 10 9 2
23 10 0 9 13 1 15 1 1 15 9 1 9 1 7 13 10 9 10 9 10 9 3 2
25 3 13 3 2 16 15 1 9 10 9 10 9 1 12 2 2 11 1 10 9 15 9 13 4 2
8 15 9 4 3 14 13 4 2
16 1 10 9 13 15 3 2 16 10 9 10 9 3 0 13 2
10 1 10 9 10 0 9 2 3 3 2
23 11 7 11 11 13 10 11 1 0 9 7 13 15 9 1 12 9 1 10 9 7 10 9
12 1 15 0 9 2 13 15 1 10 9 0 2
9 0 0 9 15 3 3 0 13 2
7 0 9 1 0 9 11 2
12 3 0 9 7 0 9 9 9 13 3 0 2
3 3 14 13
15 1 12 13 15 9 3 12 3 1 9 9 1 15 9 2
22 1 12 13 3 15 3 7 1 7 1 13 15 9 7 3 3 15 7 15 9 1 2
15 10 9 10 9 1 15 9 13 0 7 3 14 1 9 2
30 15 13 2 16 10 9 10 9 1 11 15 3 0 13 4 16 3 9 1 12 9 1 15 9 7 9 13 4 4 2
15 15 13 0 7 13 14 3 1 10 0 0 9 0 9 2
17 13 15 3 1 10 9 10 0 9 1 15 11 9 1 11 13 2
23 3 4 3 10 15 9 1 12 9 10 9 13 4 1 10 9 1 10 0 9 14 13 2
12 1 15 13 1 15 10 9 10 9 15 9 2
16 15 9 13 0 7 15 13 3 1 15 9 1 15 1 9 2
11 4 2 15 3 3 1 15 9 13 13 2
20 15 3 13 3 10 9 15 3 0 9 1 10 9 13 2 4 3 3 13 2
11 9 13 0 2 7 3 3 0 7 0 2
15 10 9 4 15 3 1 9 13 2 3 16 15 0 13 2
28 1 10 9 1 0 9 4 15 3 13 7 13 1 0 9 12 0 9 13 2 15 3 1 15 9 13 4 2
12 15 4 3 10 0 9 1 0 9 3 13 2
11 4 3 3 1 10 9 11 13 7 13 2
11 0 9 1 10 0 9 1 15 0 9 2
9 1 15 10 9 9 9 1 11 2
14 3 4 15 3 13 2 16 15 1 10 0 9 13 2
13 15 13 10 9 2 16 15 1 15 9 13 4 2
7 13 15 1 0 9 2 2
25 15 9 7 15 15 9 13 15 2 16 15 15 9 14 3 13 4 2 1 9 1 10 9 2 2
14 9 11 13 3 3 0 7 10 9 4 14 13 3 2
26 1 0 9 4 15 3 15 9 13 2 7 15 4 3 3 3 12 12 9 3 13 7 15 9 13 2
9 1 15 3 15 0 9 1 11 2
22 1 15 9 13 15 15 9 1 9 11 1 10 9 2 4 15 3 3 3 3 13 2
13 3 13 10 0 9 3 2 15 15 3 0 13 2
18 15 1 10 9 13 15 3 1 0 2 3 4 15 9 14 13 4 2
6 3 3 7 1 11 2
14 15 4 15 3 0 13 3 16 15 3 3 0 13 2
9 4 15 13 13 7 13 3 0 2
8 3 13 15 10 0 9 3 2
11 3 3 10 0 9 13 15 15 0 9 2
11 15 13 14 3 9 7 3 9 7 9 2
16 15 9 2 9 13 3 0 2 3 4 15 15 7 3 13 2
29 15 13 3 3 3 3 2 15 3 1 10 9 2 9 2 7 15 4 15 3 1 10 0 9 10 0 9 13 2
42 15 13 14 2 16 15 15 13 2 16 15 0 13 2 7 15 13 3 0 2 13 15 3 1 2 3 16 15 1 15 13 2 7 10 9 13 15 3 3 13 1 2
18 15 4 12 9 1 10 9 2 11 2 13 7 13 3 1 3 0 2
20 10 9 0 7 0 2 10 9 7 10 9 0 7 0 2 9 2 15 9 2
16 10 9 4 3 1 10 9 2 9 13 2 10 9 13 0 2
22 10 9 1 10 9 2 0 9 2 9 1 9 1 3 12 2 2 8 2 10 9 2
10 10 9 1 3 1 3 1 10 9 2
11 15 13 15 1 15 0 9 1 10 9 2
27 15 4 15 13 15 13 3 1 10 0 0 9 14 13 2 16 3 3 9 4 1 0 9 1 11 13 2
16 7 15 13 10 9 1 10 9 10 9 7 15 13 11 11 2
30 15 13 15 1 12 9 1 9 2 7 16 15 15 1 10 9 11 13 13 15 3 3 15 3 7 13 1 0 9 2
12 15 13 3 3 10 0 7 0 9 7 15 2
18 15 13 3 14 2 16 3 3 13 15 3 1 9 1 10 0 9 2
5 4 15 3 13 2
23 1 10 0 9 2 4 15 1 10 9 1 9 11 13 7 4 3 3 3 10 9 13 2
19 3 13 15 3 3 12 9 3 2 4 0 9 13 7 13 3 3 0 2
15 15 4 3 1 0 9 13 7 7 1 9 7 9 13 2
16 3 4 10 9 3 3 13 2 16 15 14 1 0 9 13 2
12 15 3 10 0 9 13 15 13 3 3 0 2
14 3 15 13 3 3 2 16 15 15 3 3 3 13 2
16 16 3 9 13 2 13 10 2 11 11 2 3 15 0 9 2
15 10 9 13 1 3 3 0 9 7 10 9 13 3 0 2
14 3 4 15 3 10 9 10 9 13 7 13 3 0 2
7 15 4 10 9 3 13 2
12 15 13 10 9 3 2 7 15 1 0 9 2
14 10 9 13 3 3 2 10 9 13 0 7 3 0 2
17 10 9 4 3 3 13 2 7 13 1 0 9 1 10 9 3 2
5 15 13 3 3 2
5 0 9 11 7 11
5 15 4 14 13 2
17 3 4 15 15 1 15 0 9 13 2 7 15 4 15 13 4 2
19 15 13 3 3 10 9 2 15 3 3 3 13 4 2 16 15 13 4 2
20 1 0 7 0 9 4 15 1 15 9 15 9 13 2 3 1 3 12 11 2
14 1 10 9 1 10 9 4 10 9 7 9 3 13 2
15 15 9 4 13 7 3 1 10 9 4 15 15 9 13 2
14 15 4 3 15 12 9 13 2 15 15 0 9 13 2
13 15 13 15 9 3 1 11 12 7 13 3 0 2
10 9 2 9 2 9 7 9 13 0 2
31 10 9 13 0 2 10 9 4 3 13 2 10 9 13 0 7 4 3 14 13 2 16 10 9 3 0 7 0 13 4 2
15 10 0 9 4 3 13 2 13 10 9 2 4 3 13 2
9 0 9 2 0 9 1 0 9 2
6 4 15 9 3 13 2
17 15 13 1 10 11 1 11 11 7 4 1 10 9 11 11 13 2
23 10 9 15 9 1 10 10 9 13 3 0 2 7 9 11 13 3 10 9 1 15 9 2
4 15 13 0 2
18 1 10 3 12 0 9 13 15 3 15 9 2 15 3 15 9 13 2
15 3 4 3 3 3 3 1 11 11 7 3 1 11 13 2
13 7 7 1 10 9 7 1 10 9 4 15 13 2
16 3 1 10 9 2 7 15 15 13 4 2 13 15 3 0 2
3 9 3 2
16 10 9 11 4 1 10 0 12 9 15 9 1 15 9 13 2
27 1 0 9 4 15 15 3 3 1 15 9 13 2 16 15 0 9 3 3 7 3 1 15 9 13 4 2
13 10 9 13 0 7 3 1 9 1 10 9 0 2
21 15 4 15 1 10 11 1 10 9 13 7 13 10 0 9 7 0 9 3 0 2
11 15 4 3 3 7 3 13 1 10 9 2
11 1 10 9 13 15 15 1 10 9 3 2
12 12 9 7 10 0 9 1 10 0 9 11 2
4 15 9 1 11
23 3 15 9 2 7 10 9 1 9 13 15 1 15 9 2 15 1 10 9 11 13 4 2
18 15 4 15 3 13 4 2 3 15 10 0 9 1 9 1 3 13 2
25 7 1 15 10 0 9 13 4 2 13 10 3 3 0 9 10 9 7 9 3 1 10 0 9 2
10 15 9 7 15 9 2 1 10 9 2
24 3 13 10 9 10 9 1 3 2 12 9 14 13 7 1 12 9 4 3 3 15 9 13 2
19 15 13 3 3 3 2 16 15 3 15 13 7 10 9 0 7 0 13 2
17 3 4 15 3 3 13 15 10 9 15 9 13 2 3 13 4 2
16 10 9 11 13 1 0 9 1 10 9 10 9 7 9 9 2
14 15 13 15 3 3 0 7 13 1 10 9 3 0 2
10 9 1 15 9 1 10 0 9 3 2
24 10 9 13 3 3 0 2 7 15 13 3 1 10 0 9 15 0 9 1 10 13 9 3 2
18 9 1 15 9 13 3 1 9 3 16 10 9 3 10 15 0 13 2
14 3 13 15 3 1 10 1 10 9 13 9 1 15 2
10 15 13 15 3 9 7 13 15 9 2
11 15 9 13 10 9 3 3 3 0 1 2
23 1 10 9 1 15 13 4 2 16 10 0 9 15 13 2 13 15 15 10 9 3 3 2
20 10 9 10 0 9 13 3 3 0 7 3 13 15 9 3 1 10 0 9 2
12 10 11 13 10 0 9 1 0 9 2 9 2
3 0 9 2
13 1 10 9 10 9 13 10 9 10 9 15 9 2
18 3 1 10 0 9 4 15 14 13 2 16 15 3 1 10 9 13 2
11 10 9 10 9 13 3 1 10 9 0 2
11 9 15 9 13 10 9 10 11 14 13 2
34 15 4 15 3 1 10 11 3 1 9 13 7 15 9 13 15 2 15 4 3 3 13 1 10 11 3 7 15 4 3 3 9 13 2
11 1 10 9 13 3 3 15 11 3 3 2
11 7 3 3 10 0 0 9 1 0 9 2
25 1 3 10 9 1 10 9 7 1 9 13 15 15 3 2 16 3 10 9 3 3 9 13 4 2
5 15 13 3 0 2
7 0 9 2 9 1 9 2
14 0 7 0 9 2 1 0 9 2 2 7 0 9 2
20 3 13 4 15 16 15 0 9 1 9 7 10 9 1 10 9 2 9 13 2
9 9 4 3 3 1 0 9 13 2
7 15 4 3 15 9 13 2
10 7 10 9 2 9 2 9 13 3 2
16 15 4 3 14 3 13 2 16 15 1 15 9 0 9 13 2
6 10 9 1 10 9 2
9 15 13 2 13 7 13 3 3 2
20 15 13 3 1 15 9 1 10 11 11 2 16 10 9 3 10 9 3 13 2
24 15 9 4 3 14 3 1 9 13 2 7 1 10 0 9 13 15 15 3 1 0 9 3 2
4 13 12 9 2
21 4 3 15 9 14 13 2 16 10 11 1 13 9 7 9 10 9 14 13 4 2
11 4 9 3 3 13 4 16 15 13 4 2
13 1 3 12 8 8 13 15 3 3 14 3 0 2
5 2 3 0 9 2
12 15 13 3 1 10 9 10 11 11 1 11 2
8 15 4 3 3 3 3 13 2
31 10 9 13 3 0 1 10 0 11 2 9 7 13 1 0 9 2 9 2 9 2 9 7 9 2 10 0 9 7 9 2
30 3 16 15 10 9 13 13 15 10 0 9 1 0 9 2 10 0 9 2 0 9 1 0 9 7 0 0 9 1 2
12 10 9 13 3 0 7 15 13 1 0 9 2
15 15 4 15 15 3 1 10 9 13 2 15 4 15 13 2
14 0 9 7 10 9 13 3 2 3 15 13 10 3 0
10 15 13 3 0 2 16 15 15 13 2
7 4 3 14 15 13 4 2
40 15 13 1 15 9 10 9 2 15 15 1 0 9 1 10 9 2 10 9 2 10 9 10 9 2 10 9 1 10 9 7 3 10 9 10 9 2 9 13 2
8 3 13 11 11 15 0 9 2
26 15 13 1 15 2 16 11 11 10 9 15 9 2 9 1 10 0 9 1 10 0 9 3 13 4 2
18 1 15 13 11 11 1 10 0 9 4 2 15 15 14 3 13 4 2
11 15 13 10 0 9 10 9 15 9 13 2
12 3 4 15 3 3 3 13 7 15 4 13 2
11 3 13 15 1 15 1 12 9 3 0 2
9 9 11 4 3 3 1 15 13 2
22 15 4 15 1 15 9 13 7 13 15 15 14 13 2 15 1 10 9 3 13 4 2
5 15 13 3 0 2
13 1 15 9 4 15 3 3 1 9 11 13 2 2
22 15 4 15 10 9 13 13 7 13 3 1 12 9 2 15 15 0 9 3 13 4 2
33 10 9 13 15 3 9 9 11 7 7 15 13 2 13 10 9 2 15 15 3 13 12 8 1 15 10 0 15 9 2 2 2 2
10 7 10 9 13 3 0 1 2 2 2
19 13 3 3 1 15 9 1 9 9 11 1 9 7 15 4 3 13 4 2
12 9 9 11 13 10 3 0 7 3 0 9 2
19 10 9 13 3 3 0 2 0 9 2 0 7 0 9 2 15 0 2 2
6 4 15 3 3 13 2
15 3 3 13 15 10 3 9 1 10 9 1 9 9 11 2
17 3 4 15 3 13 7 4 3 12 9 13 2 3 1 9 2 2
14 10 9 1 10 9 13 3 0 3 3 10 9 9 2
9 4 1 15 9 15 0 9 13 2
4 3 14 13 2
9 0 7 0 9 3 1 10 9 2
5 0 9 1 9 2
18 15 13 0 9 1 10 11 7 13 3 1 10 9 15 3 13 4 2
15 15 13 12 0 9 2 15 3 3 1 15 9 13 4 2
19 3 13 15 10 11 10 0 9 13 2 3 16 15 15 9 14 13 4 2
17 3 13 15 2 13 10 11 3 2 16 10 9 1 9 13 4 2
17 3 15 13 3 0 9 15 15 9 13 4 7 15 3 0 13 2
6 9 10 9 1 10 9
14 10 9 11 13 10 3 0 9 2 3 3 14 13 2
13 4 3 3 13 2 3 13 3 10 9 3 0 2
23 10 9 13 3 3 1 10 0 9 3 10 0 9 9 13 4 16 15 10 9 14 13 2
19 10 9 4 1 9 13 7 10 9 15 1 15 1 9 7 2 9 13 2
6 3 0 9 7 9 2
5 4 15 3 13 2
16 9 11 13 3 0 2 3 1 10 9 13 7 13 3 0 2
9 10 9 8 9 13 3 3 0 2
14 15 9 1 10 9 1 15 15 3 13 1 15 9 2
19 9 11 13 15 3 3 1 10 9 8 9 3 7 4 15 3 3 13 2
3 15 0 2
13 0 9 7 10 9 13 1 3 3 3 0 9 2
10 1 10 11 11 4 9 3 0 13 2
15 10 9 2 9 2 9 7 3 10 9 13 3 0 2 2
12 3 11 11 7 10 11 11 4 0 9 13 2
22 10 9 13 3 3 1 15 9 1 10 9 9 2 9 8 2 2 1 10 9 9 2
15 1 10 9 13 3 3 9 2 11 2 16 15 15 13 2
12 15 4 14 3 1 10 9 9 10 9 13 2
3 3 0 2
11 3 0 11 11 13 3 7 15 13 2 2
13 15 8 15 13 15 3 3 1 10 0 9 2 2
9 10 9 7 10 9 13 3 0 2
15 10 9 1 10 11 11 2 11 4 15 1 15 9 13 2
14 15 13 15 1 9 1 10 0 9 1 11 7 11 2
34 1 10 0 9 13 15 3 0 7 3 10 9 13 0 7 13 15 10 9 1 10 0 9 2 15 3 3 3 13 2 16 9 13 2
29 15 4 15 1 10 0 9 1 9 2 7 9 3 3 3 13 2 16 15 1 9 12 9 1 0 9 13 4 2
13 1 10 9 1 9 1 11 13 15 3 14 3 2
9 15 1 15 3 14 13 2 2 2
12 16 15 3 9 4 13 2 3 1 11 11 2
15 0 0 9 2 3 7 1 10 9 2 9 11 2 11 2
12 15 9 1 9 2 15 15 9 1 9 13 2
14 3 13 15 0 9 2 10 0 9 1 3 12 9 2
11 10 9 11 13 1 9 3 1 15 9 2
13 1 11 11 13 15 0 0 9 1 3 0 9 2
14 10 9 7 10 9 13 3 0 7 10 9 13 0 2
21 15 13 3 10 0 9 9 7 3 13 15 3 3 10 0 9 7 10 0 9 2
13 10 9 13 3 0 7 10 0 9 13 3 0 2
10 1 15 15 10 0 9 9 1 11 2
11 13 10 9 1 10 9 2 13 3 0 2
19 10 9 3 1 10 11 2 15 3 1 10 15 3 13 2 13 3 0 2
28 10 9 13 0 7 13 9 7 10 0 2 0 9 2 9 2 15 15 3 1 12 2 9 2 9 14 13 2
10 10 9 13 3 0 2 0 7 0 2
7 1 10 9 3 14 13 2
7 0 9 15 3 13 4 2
11 1 10 0 9 8 4 10 9 3 13 2
31 10 9 4 15 1 15 0 9 3 13 7 13 10 0 9 1 9 2 9 2 9 8 10 9 13 0 2 0 7 0 2
5 0 9 1 15 9
16 1 10 11 11 9 4 15 1 10 9 1 9 11 0 13 2
12 15 13 3 3 3 2 12 9 9 1 11 2
14 1 10 9 7 9 15 9 11 11 13 15 3 0 2
26 1 15 9 4 15 3 3 15 9 13 7 3 13 1 10 9 1 0 0 9 1 0 9 2 9 2
15 3 4 15 1 10 0 9 1 10 9 11 1 9 13 2
13 15 4 15 3 13 2 7 4 3 3 9 13 2
4 0 0 9 2
4 9 13 0 2
3 0 9 2
7 9 3 0 2 11 11 2
4 13 3 0 2
6 13 15 3 14 3 2
5 15 13 15 0 2
6 3 13 0 9 9 2
7 0 9 9 1 9 2 11
12 13 0 9 1 11 7 4 10 9 3 13 2
10 9 4 3 3 7 1 0 9 13 2
14 4 15 3 1 10 9 13 7 3 1 10 9 13 2
23 13 3 1 10 11 7 1 10 11 2 9 13 0 7 13 9 2 1 15 15 15 13 2
9 4 15 10 0 9 3 14 13 2
14 13 10 9 3 15 9 7 4 3 3 0 9 13 2
3 13 3 2
15 15 4 13 7 13 3 1 9 15 9 15 15 3 13 2
6 3 3 0 7 0 2
19 10 9 10 9 13 3 11 2 9 7 13 15 11 2 13 11 2 9 2
11 3 13 15 1 10 9 2 11 1 11 2
13 16 15 15 3 14 13 13 2 13 15 15 3 2
21 3 1 10 0 9 2 15 13 3 12 9 2 4 15 3 3 1 15 9 13 2
14 15 13 3 3 14 1 9 2 7 10 9 13 1 2
24 12 9 3 13 15 9 1 7 1 9 1 9 2 9 7 9 1 10 9 3 13 15 9 2
24 15 4 15 13 3 4 15 12 9 7 12 9 13 16 15 9 13 2 15 15 1 15 13 2
16 1 10 9 13 15 15 2 9 2 10 9 13 3 12 9 2
18 7 3 3 2 10 9 1 10 9 3 1 9 2 3 1 10 9 2
6 15 13 15 9 13 2
23 4 15 10 9 3 1 12 9 13 2 4 15 15 15 9 2 9 2 9 7 9 13 2
12 3 1 15 9 2 9 3 2 9 15 13 2
9 1 3 13 15 10 9 15 9 2
12 7 16 15 1 10 9 13 13 15 15 8 2
11 3 4 15 1 15 2 0 2 9 13 2
7 15 9 13 15 15 13 2
13 3 10 9 3 15 15 9 1 10 0 9 13 2
10 3 13 9 9 9 7 13 3 0 2
16 15 13 1 12 9 10 11 11 7 13 15 3 3 3 0 2
16 4 1 10 12 9 10 9 2 1 9 0 9 2 3 13 2
20 7 3 3 4 15 3 3 2 3 3 7 3 3 7 1 9 11 13 4 2
12 9 13 3 3 1 15 10 0 9 14 13 2
20 7 16 15 15 3 10 0 9 13 2 4 15 3 9 1 10 0 9 13 2
9 10 9 13 1 15 3 10 9 2
9 7 15 4 1 9 11 3 13 2
7 15 13 3 9 1 15 2
27 3 13 15 16 15 14 3 12 9 2 9 1 9 13 1 15 1 9 11 3 7 3 2 13 14 13 2
17 15 13 1 15 9 3 0 0 9 15 10 9 10 9 3 13 2
11 9 1 0 9 1 9 11 1 10 9 2
6 15 4 10 9 13 2
6 3 0 7 1 9 2
12 9 3 0 2 16 15 10 9 14 13 4 2
15 16 15 3 1 11 9 13 4 2 13 15 3 3 3 2
8 10 9 10 9 13 3 0 2
17 15 13 3 3 2 1 0 2 9 2 3 13 15 3 0 9 2
11 3 13 15 0 0 9 1 10 9 8 2
5 10 9 13 0 2
7 3 13 15 15 9 3 2
5 15 13 3 3 2
13 10 9 13 0 16 15 13 7 10 9 13 0 2
13 10 9 13 0 7 3 3 15 15 10 9 13 2
7 3 1 15 3 14 13 2
20 15 9 13 3 3 14 3 1 11 2 11 0 7 10 9 13 14 10 0 2
5 15 4 13 4 2
3 11 13 2
26 10 11 13 10 0 9 2 1 15 1 9 14 13 2 1 10 9 14 13 7 10 9 13 14 13 2
8 15 13 3 3 1 10 11 2
11 1 10 0 9 13 15 3 3 15 9 2
12 10 9 13 3 13 9 1 10 11 2 9 2
25 9 7 9 4 1 15 9 3 0 13 7 15 4 15 1 10 9 1 9 7 15 9 3 13 2
13 3 13 15 7 10 9 7 3 10 9 10 11 2
16 15 4 11 1 11 1 0 9 10 9 7 9 1 9 13 2
12 1 11 13 15 3 9 7 9 1 10 9 2
14 11 11 13 15 10 0 2 7 3 14 15 10 9 2
16 10 9 1 10 9 10 9 7 3 1 10 11 13 3 0 2
19 3 4 15 13 2 3 0 9 13 2 15 10 9 10 9 3 0 13 2
39 15 4 14 3 3 1 15 9 13 2 12 1 12 9 2 2 7 3 1 10 9 2 1 10 9 0 9 3 1 10 9 13 2 16 15 14 0 13 2
11 0 7 0 13 10 9 2 7 3 0 2
14 16 15 3 1 9 13 2 4 15 3 0 9 13 2
19 10 3 1 10 9 13 9 13 3 0 2 16 15 15 3 3 13 4 2
33 10 9 1 10 9 10 0 9 13 2 7 15 14 10 0 9 2 12 9 2 13 2 15 1 10 2 9 2 2 9 0 13 2
9 0 9 1 10 9 13 0 1 2
7 3 13 10 9 3 9 2
14 3 4 3 3 13 2 0 7 0 7 1 0 9 2
6 3 13 15 3 0 2
10 4 0 9 10 11 9 1 11 13 2
14 10 9 11 9 2 9 2 13 3 0 7 3 13 2
15 1 15 11 9 1 7 1 11 4 15 15 9 3 13 2
8 15 4 1 15 9 3 13 2
11 15 0 9 16 15 1 9 7 9 13 2
12 4 3 3 3 13 7 4 15 3 3 13 2
14 4 3 3 3 3 13 7 15 4 3 15 3 13 2
18 1 10 9 13 15 3 0 2 7 3 1 10 9 13 15 15 13 2
6 0 9 7 0 9 2
13 15 13 1 9 3 15 9 7 4 3 3 13 2
12 15 13 15 9 15 1 15 14 13 4 4 2
9 3 0 9 2 0 9 7 9 2
5 15 13 15 3 2
12 3 0 9 7 10 9 13 3 3 12 9 2
14 15 13 3 0 1 11 7 4 3 3 3 3 13 2
10 2 10 9 11 13 3 3 0 2 2
21 10 9 11 13 14 3 10 0 9 1 0 9 2 15 13 3 3 10 0 9 2
6 12 9 4 15 13 2
19 12 9 13 10 9 3 0 7 12 9 3 13 15 10 0 9 1 9 2
6 3 13 9 9 9 2
16 1 9 1 9 7 9 13 10 9 11 11 11 15 0 9 2
7 15 4 1 10 9 13 2
11 1 10 9 4 15 3 1 10 9 13 2
11 9 11 13 15 10 9 13 7 14 13 2
12 1 10 9 4 15 1 15 3 10 9 13 2
14 10 9 13 14 1 9 7 4 3 1 10 9 13 2
5 15 4 15 13 2
6 10 9 4 3 13 2
8 10 9 1 10 9 13 0 2
8 1 10 9 13 15 7 13 2
16 13 3 3 3 2 16 15 1 12 1 11 1 9 13 4 2
25 15 9 2 9 4 3 13 7 1 10 0 9 1 10 9 4 15 3 15 9 1 10 9 13 2
5 10 9 13 0 2
24 16 15 10 9 13 4 7 15 3 3 3 13 4 2 13 15 15 1 9 2 9 7 9 2
34 1 12 9 13 15 1 10 0 9 1 10 9 1 9 11 2 15 15 3 10 9 15 9 3 13 1 9 2 9 1 9 13 4 2
8 10 9 13 1 15 0 9 2
5 10 9 13 3 2
6 4 15 1 9 13 2
14 10 9 13 3 1 10 13 9 0 7 13 0 9 2
6 15 1 15 3 13 2
20 16 15 9 3 14 1 9 13 2 13 15 15 3 3 15 10 3 13 9 2
22 3 15 1 9 2 7 15 15 3 0 7 0 13 2 15 13 3 3 1 15 9 2
8 15 3 4 3 3 3 13 2
8 10 9 13 0 2 3 0 2
12 3 4 15 15 1 10 9 13 7 3 13 2
9 3 13 15 9 1 10 11 14 2
6 15 4 3 15 13 2
8 10 9 3 13 3 3 0 2
12 15 13 3 3 1 9 15 1 9 13 4 2
16 15 13 9 2 15 1 10 9 13 4 2 15 14 0 13 2
8 10 9 15 9 13 3 0 2
14 13 9 2 1 9 2 1 0 9 7 10 0 9 2
18 3 13 10 9 1 10 9 9 2 16 10 9 13 1 10 9 0 2
10 9 4 10 9 1 10 9 13 13 2
7 15 4 15 10 11 13 2
15 15 13 1 10 9 1 11 1 15 9 1 11 7 11 2
11 15 4 3 1 15 9 10 0 9 13 2
10 3 4 15 15 1 0 9 3 13 2
19 15 13 15 9 1 9 7 15 15 3 13 4 1 15 10 0 9 13 2
8 10 9 13 3 0 7 0 2
18 15 4 8 9 13 7 15 10 9 1 10 9 11 1 10 11 13 2
7 15 4 10 9 3 13 2
7 15 13 3 3 0 1 2
17 16 10 9 7 10 9 1 10 11 13 4 15 10 9 3 13 2
6 10 9 13 3 0 2
6 15 13 15 3 3 2
13 1 15 10 0 9 7 10 0 9 13 3 0 2
14 1 15 9 13 15 3 0 10 0 9 13 14 4 2
37 10 9 1 10 11 13 3 0 2 15 13 1 10 0 9 1 2 15 9 4 3 13 2 15 9 2 11 2 13 10 9 1 10 0 9 1 2
9 15 1 15 0 9 3 15 13 2
21 3 1 10 15 9 13 15 10 9 1 10 9 10 9 7 10 9 10 0 9 2
7 1 15 9 4 15 13 2
10 15 9 13 10 0 9 9 2 2 2
17 15 4 3 14 13 2 4 3 3 13 7 4 10 9 3 13 2
13 15 4 3 15 9 13 7 15 13 0 7 0 2
13 1 15 9 4 15 3 10 9 7 10 9 13 2
5 15 13 3 0 2
14 15 13 10 0 2 0 9 2 3 3 10 9 3 2
7 10 0 9 13 15 14 2
21 10 9 4 14 13 2 13 1 10 9 7 15 13 15 9 2 9 7 9 8 8
23 10 9 13 3 0 2 10 9 13 3 3 3 15 9 1 7 4 3 1 10 9 13 2
13 0 2 7 15 4 15 9 3 14 13 2 2 2
24 3 2 10 9 13 3 3 1 10 9 7 15 4 15 1 10 9 7 9 14 3 3 13 2
10 10 9 13 0 7 13 14 3 0 2
13 1 10 9 13 1 15 10 0 0 7 0 9 2
15 10 11 13 0 2 10 9 3 13 15 3 14 3 0 2
18 10 9 2 13 3 3 0 2 15 13 15 3 0 1 10 10 9 2
12 3 4 15 3 3 15 15 9 1 11 13 2
9 15 13 0 1 15 3 14 13 2
9 3 4 15 3 13 2 2 2 2
5 15 13 3 0 2
15 10 9 10 9 11 1 10 9 11 13 0 1 10 9 2
13 10 9 0 2 0 1 10 9 7 3 3 13 2
14 10 9 14 15 2 7 1 10 9 7 9 3 0 2
9 4 1 3 15 3 3 15 13 2
8 15 4 10 9 1 9 13 2
19 10 9 1 10 12 2 9 10 11 11 11 14 9 1 11 4 3 13 2
16 9 13 10 0 9 3 1 10 9 2 15 1 0 9 13 2
16 1 10 0 9 13 10 9 2 16 15 13 2 15 9 1 2
9 10 9 13 0 9 1 0 9 2
21 10 1 11 0 9 1 10 9 7 10 9 4 13 7 13 10 9 1 10 3 2
7 10 9 13 0 2 2 2
13 0 13 2 10 9 12 2 9 2 13 3 0 2
9 10 0 9 13 3 1 10 9 2
15 10 9 13 3 0 7 9 4 15 1 12 9 3 13 2
6 10 9 13 3 0 2
15 3 4 15 1 2 3 2 15 9 2 7 9 3 13 2
9 15 13 0 9 1 10 11 13 2
4 15 13 0 2
10 3 13 15 1 9 14 10 0 9 2
7 15 4 15 3 0 13 2
11 3 3 1 10 9 13 10 9 3 0 2
9 1 15 9 13 15 10 15 9 2
7 15 9 13 3 3 0 2
10 1 10 9 13 16 15 3 0 13 2
14 1 10 9 15 9 4 15 1 9 3 12 8 13 2
13 3 13 10 9 3 0 7 10 9 13 3 0 2
17 1 0 9 4 15 13 14 13 2 16 15 9 3 13 4 4 2
12 15 4 15 3 3 13 1 3 15 14 13 2
15 3 13 10 9 9 1 9 7 2 7 1 0 9 1 2
8 15 13 10 9 3 10 9 2
5 3 3 3 0 2
6 10 9 13 3 0 2
17 3 4 10 9 1 15 9 3 3 1 10 9 1 10 15 13 2
13 10 9 13 0 7 0 2 7 15 13 14 1 2
20 15 4 10 9 1 0 9 13 7 10 9 1 0 9 1 10 9 3 13 2
17 15 0 9 4 12 0 9 13 7 15 4 3 3 10 9 13 2
25 3 3 4 3 3 10 9 13 4 2 15 4 14 13 2 16 10 9 12 9 1 10 9 13 2
16 3 13 15 3 3 2 16 15 9 1 0 9 13 4 4 2
12 3 4 15 15 1 15 0 9 12 8 13 2
11 1 10 9 13 15 3 3 3 12 8 2
4 11 13 0 2
20 3 1 15 10 0 9 1 10 9 2 16 14 3 3 10 11 11 3 13 2
6 10 9 13 3 15 2
11 3 13 15 3 0 0 9 1 10 9 2
18 7 15 4 13 15 15 14 3 1 10 9 3 1 10 15 9 13 2
33 10 9 13 3 10 9 10 0 0 9 2 15 15 0 9 1 10 9 1 9 2 7 9 7 10 9 1 9 2 7 9 13 2
40 11 2 11 2 9 1 11 0 9 11 2 11 2 13 2 7 10 11 1 10 9 10 0 0 9 2 10 9 1 9 7 9 3 14 10 0 9 13 4 2
11 10 9 13 15 3 2 10 15 13 15 2
16 15 13 3 2 16 15 10 9 10 0 12 9 1 9 13 2
20 11 13 3 9 1 10 0 9 2 16 10 0 9 4 15 1 10 15 13 2
13 11 13 0 7 13 15 3 1 10 0 9 3 2
36 11 2 9 2 10 11 7 11 4 11 9 11 11 3 1 10 11 13 2 10 9 1 10 9 11 11 2 11 7 12 0 9 0 14 13 2
15 1 10 9 13 10 9 1 10 9 1 1 9 12 9 2
13 12 9 13 3 0 2 16 10 9 1 9 13 2
26 10 9 1 11 13 10 0 0 9 1 10 9 7 9 10 0 9 1 10 0 9 2 2 13 9 2
25 1 10 11 4 10 11 1 10 9 10 1 10 12 2 11 12 0 9 10 11 1 10 11 13 2
9 10 9 13 3 9 1 9 11 2
14 9 10 9 4 3 10 2 0 9 1 11 13 2 2
4 11 13 11 2
7 10 9 13 1 10 9 2
22 10 0 9 13 2 10 0 9 7 15 12 9 0 9 4 1 9 13 2 11 13 2
26 10 9 10 11 11 2 11 11 2 13 2 10 11 4 3 13 2 2 15 0 9 15 13 4 2 2
13 3 4 3 12 9 0 2 3 0 9 13 4 2
12 10 9 4 10 9 10 0 0 9 1 12 13
7 9 13 7 13 10 15 2
9 10 0 9 13 9 1 10 9 2
15 10 9 13 3 14 1 15 9 2 15 1 9 0 13 2
7 7 15 13 15 14 13 2
12 10 9 10 9 2 7 9 13 10 11 14 2
14 10 9 4 15 1 10 0 2 0 2 9 2 13 2
10 10 9 1 13 10 9 10 0 9 2
41 10 9 10 9 1 9 10 9 13 1 10 9 3 10 9 2 13 10 11 2 11 2 1 10 1 10 11 1 11 0 9 2 8 2 12 8 12 2 12 2 2
15 0 9 7 9 4 13 2 1 10 9 15 9 14 13 2
15 10 9 1 10 0 2 9 2 13 3 10 0 9 3 2
13 3 4 15 10 9 10 9 3 13 2 13 15 2
18 1 0 9 4 10 9 15 9 1 9 1 10 9 1 10 9 13 2
24 10 9 1 10 9 2 15 1 10 0 9 1 11 1 10 0 9 13 4 2 13 15 14 2
19 10 0 9 4 1 10 11 12 0 11 2 9 1 10 9 10 9 13 2
20 10 9 10 1 0 9 1 15 9 4 15 1 12 1 12 1 12 12 13 2
13 10 2 9 2 4 15 9 1 10 0 11 13 2
30 10 9 4 3 3 14 3 7 1 0 9 1 3 0 9 13 4 2 7 1 3 0 9 2 15 1 0 9 13 2
24 10 0 9 2 10 9 10 9 14 13 2 13 3 10 0 9 2 2 13 11 11 1 11 2
13 10 9 10 9 1 9 1 10 9 13 10 9 2
16 10 9 0 9 4 15 1 0 9 3 3 1 10 9 13 2
32 10 9 4 15 13 2 16 15 10 9 3 13 4 7 10 9 10 9 13 4 2 1 15 10 0 9 2 15 3 13 2 2
28 10 9 11 2 8 12 2 2 11 2 8 12 2 7 11 2 11 2 8 2 9 2 13 3 3 0 9 2
23 10 11 4 10 0 9 10 9 2 1 9 2 9 2 9 2 9 2 7 9 13 2 2
13 10 11 13 1 15 3 1 10 9 1 11 11 2
16 9 11 11 2 9 2 13 15 1 0 9 1 11 2 9 2
18 10 9 1 10 11 2 9 1 15 9 1 11 4 1 10 11 13 2
22 11 13 15 1 15 9 2 4 7 3 1 11 3 13 2 16 15 1 10 9 13 2
9 10 9 4 1 10 11 13 4 2
7 9 13 10 9 15 9 2
10 9 13 15 14 3 1 10 0 9 2
7 12 13 15 3 10 9 2
18 15 13 10 9 2 16 10 0 9 1 10 9 1 3 0 13 4 2
23 9 1 10 9 2 13 7 1 10 9 1 0 9 7 3 1 10 9 2 7 0 9 2
33 10 9 10 9 13 15 0 9 1 10 0 9 10 9 1 10 9 0 7 13 10 9 0 9 1 10 11 15 9 1 0 9 2
29 10 9 13 1 9 0 2 4 7 2 7 1 15 3 0 9 10 0 9 2 3 3 3 1 10 9 13 4 2
39 15 13 3 2 16 7 15 10 9 13 7 13 2 3 15 13 2 15 1 9 14 13 13 2 2 13 10 9 2 16 15 1 10 9 9 14 13 13 2
21 15 1 11 3 1 10 9 13 4 2 4 15 1 10 9 14 1 10 9 13 2
9 10 9 13 3 3 1 10 9 2
8 1 11 13 9 10 9 3 2
35 10 9 7 9 2 15 11 13 2 13 1 10 9 10 9 13 2 15 2 3 1 15 11 2 9 2 10 9 2 0 9 2 13 4 2
8 3 0 2 13 11 11 15 2
7 9 2 15 15 13 4 2
17 15 13 1 10 0 0 9 1 0 0 9 2 2 13 15 3 2
16 3 13 15 10 9 2 7 10 0 9 13 15 3 14 0 2
13 10 9 10 9 9 12 13 1 10 9 11 11 2
22 10 9 2 3 10 9 12 10 11 2 13 0 9 1 10 9 1 10 0 9 3 2
26 0 9 13 15 9 3 3 1 2 7 9 14 0 13 2 9 1 10 0 9 1 15 0 14 13 2
22 10 9 10 9 13 1 10 0 9 1 2 1 15 10 9 0 13 2 10 9 13 2
16 11 2 11 11 2 11 11 2 11 11 7 15 15 13 0 2
19 15 4 14 13 2 16 15 15 9 13 4 2 15 4 15 9 3 13 2
19 11 2 15 1 10 0 11 11 1 10 0 11 2 11 13 2 13 9 2
18 10 0 9 10 9 13 10 9 10 0 9 2 10 9 7 10 9 2
21 10 9 13 3 1 9 2 16 11 10 9 3 1 10 9 1 10 9 13 4 2
23 10 1 3 12 9 0 9 1 10 9 11 2 11 13 1 10 0 11 10 0 9 3 2
12 10 0 9 13 1 11 7 13 15 10 9 2
16 10 9 4 3 1 0 9 1 10 9 15 11 2 9 13 2
32 11 11 7 11 2 9 11 11 13 1 15 9 1 10 12 2 9 1 10 11 1 11 10 9 1 2 10 0 9 10 11 2
26 1 9 1 9 11 11 4 10 9 3 1 10 9 13 2 2 16 15 9 1 15 9 13 4 2 2
25 10 9 1 11 2 11 7 11 13 15 3 1 9 3 2 10 9 1 10 9 10 9 14 13 2
21 9 4 15 9 3 15 2 0 2 2 2 0 2 7 2 0 2 9 3 13 2
20 10 9 10 9 1 10 9 1 9 2 11 11 2 13 10 0 9 10 9 2
14 12 12 9 13 1 12 9 7 4 1 12 9 13 2
23 9 11 11 4 10 9 1 10 9 1 15 0 9 11 11 1 2 0 9 3 2 13 2
16 1 1 10 15 4 0 12 9 15 9 13 2 2 13 9 2
11 3 4 15 3 7 3 13 7 9 13 2
8 1 10 12 2 11 13 9 2
16 11 13 1 11 7 11 1 2 9 2 9 7 9 2 3 2
32 10 11 2 11 2 4 9 1 10 9 10 0 9 13 2 1 15 9 1 10 9 1 3 12 9 15 9 1 9 13 4 2
12 12 9 13 10 9 1 1 10 9 12 1 2
26 9 13 15 1 10 0 9 1 2 7 1 10 11 13 10 9 1 11 1 10 9 1 9 7 9 2
18 11 11 13 1 10 0 12 9 1 10 9 1 10 11 1 10 11 2
22 10 9 2 7 9 11 4 3 3 3 1 10 9 1 9 13 2 13 9 11 11 2
12 0 9 13 1 3 1 10 9 9 7 9 2
8 1 11 13 15 1 10 9 2
12 15 13 9 2 3 0 9 2 2 13 15 2
20 9 11 11 13 1 10 11 10 9 1 10 11 2 11 2 9 1 11 1 2
13 11 11 4 15 10 9 13 2 2 13 10 9 2
7 10 9 10 9 13 0 2
31 3 13 15 1 10 9 10 9 1 9 2 15 1 9 1 0 9 13 4 2 2 13 15 1 10 1 10 11 0 9 2
27 10 11 2 9 11 11 13 10 9 2 16 10 9 3 10 9 1 10 9 1 10 9 1 10 11 13 2
25 10 9 13 1 10 9 11 10 9 2 16 15 10 11 1 10 0 9 3 1 10 9 13 4 2
28 10 9 13 3 1 12 9 8 1 10 9 1 11 2 11 2 11 2 1 7 13 12 9 3 10 9 3 2
15 11 13 10 9 1 2 15 4 1 10 9 0 9 13 2
19 10 9 10 9 13 15 3 0 2 16 1 15 9 7 9 13 4 4 2
14 10 11 2 11 4 15 0 9 1 9 1 9 13 2
6 11 7 11 13 9 2
23 9 2 10 15 3 2 13 1 10 12 9 9 11 2 9 11 2 9 11 7 9 11 2
18 9 1 9 7 0 9 1 10 12 2 9 13 10 9 2 9 0 2
13 9 1 9 7 9 13 3 9 1 9 7 9 2
13 10 9 13 1 10 12 2 11 1 12 2 11 2
17 10 11 11 13 1 15 9 10 9 1 10 12 2 11 12 1 2
42 3 4 15 3 3 13 2 2 13 10 0 9 15 9 2 15 15 1 9 1 9 2 7 9 13 2 16 11 7 11 1 10 12 2 11 1 0 9 15 9 13 2
17 9 11 11 13 11 1 10 11 3 1 2 15 9 1 11 13 2
19 9 13 1 10 0 2 0 9 2 10 9 7 10 0 9 1 10 9 2
14 15 13 3 1 10 0 9 1 2 1 9 10 9 2
11 10 9 11 13 10 0 9 2 0 2 2
20 15 13 15 2 16 10 9 3 13 7 15 0 9 2 2 13 9 11 11 2
21 3 13 10 9 10 9 1 2 0 9 2 1 10 9 2 15 15 1 11 13 2
21 9 2 16 3 0 0 9 1 10 11 13 7 15 0 13 2 4 10 9 13 2
10 10 9 4 3 1 10 9 13 4 2
20 1 10 11 4 10 0 9 12 0 0 9 13 2 15 1 10 9 13 4 2
22 10 0 9 2 9 7 9 13 7 3 0 2 16 0 10 9 13 2 4 13 4 2
17 9 10 9 7 14 3 10 9 10 9 7 9 13 3 10 9 2
13 10 9 13 15 2 16 9 0 7 14 0 13 2
13 10 9 13 2 16 3 12 9 1 10 9 13 2
12 10 9 13 3 3 1 9 1 9 10 9 2
12 12 12 9 4 13 2 10 9 1 9 13 2
23 11 13 1 10 0 9 0 9 1 10 0 9 1 10 9 2 1 15 1 9 7 9 2
11 2 8 8 2 4 3 1 10 9 13 2
10 11 4 1 10 9 12 1 11 13 2
13 0 9 13 3 3 1 10 9 10 9 7 9 2
6 3 13 15 15 3 2
15 10 9 4 1 12 9 9 1 10 9 1 12 9 13 2
28 15 13 3 0 2 4 15 15 15 9 1 10 9 13 2 2 13 10 3 1 10 9 10 0 9 0 9 2
13 10 9 4 1 10 0 12 9 12 9 9 13 2
19 11 4 1 10 0 9 10 0 9 1 9 11 3 1 10 0 9 13 2
35 3 13 10 9 9 1 10 9 2 16 15 13 4 2 3 13 2 15 3 13 4 2 2 13 11 11 2 9 2 9 1 10 9 11 2
20 10 9 4 1 10 12 2 11 1 12 3 3 12 9 1 10 9 0 13 2
15 9 13 15 2 10 9 14 13 7 10 9 1 9 13 2
20 10 9 1 11 2 11 13 14 3 15 2 15 15 3 13 2 2 13 11 2
38 9 10 0 9 13 10 9 10 2 9 2 1 0 9 2 10 9 7 9 10 9 1 0 9 1 15 1 9 10 9 7 11 2 9 7 0 9 2
25 10 9 13 1 10 9 10 9 1 9 2 13 10 9 15 9 2 3 13 10 9 3 0 9 2
16 15 13 2 3 1 10 9 10 11 10 9 13 14 4 2 2
27 10 0 9 11 11 4 10 9 13 7 13 9 1 10 9 2 9 7 13 15 3 3 1 15 9 1 2
42 9 0 9 13 3 10 9 9 10 0 9 2 11 2 1 11 1 11 2 1 10 0 9 1 10 9 10 9 2 9 7 9 10 0 9 1 9 12 8 9 13 2
11 10 9 13 9 2 16 15 15 9 13 2
31 15 13 9 2 7 13 15 15 15 0 9 2 15 13 9 2 7 15 9 2 15 13 15 9 2 7 3 10 9 2 2
15 1 9 4 15 3 9 1 10 9 1 11 1 0 13 2
20 10 9 1 11 13 1 9 10 0 11 2 11 1 9 1 10 0 9 1 2
14 10 9 4 10 1 10 9 0 9 7 13 7 13 2
28 1 11 13 15 9 1 10 0 9 2 7 9 1 2 1 15 1 15 9 1 10 9 1 10 0 0 9 2
26 9 13 10 9 10 9 1 11 1 10 0 9 2 3 7 1 0 9 2 13 15 1 10 0 9 2
47 10 11 2 9 11 11 2 12 9 0 2 1 0 9 3 9 10 0 11 11 11 2 4 1 10 9 15 0 9 3 1 2 9 2 10 11 11 2 9 2 9 7 9 1 9 13 2
12 11 7 10 15 0 0 9 11 11 13 0 2
36 9 11 11 2 11 2 2 11 11 2 10 11 7 9 13 10 9 7 10 2 0 9 2 7 2 3 0 2 7 1 10 9 2 0 2 2
17 0 9 4 1 12 9 7 10 0 9 4 1 12 9 3 13 2
21 11 11 13 1 10 11 1 10 9 1 2 15 13 2 15 9 2 1 10 9 2
21 9 13 1 10 9 1 12 9 3 7 4 1 0 9 13 7 1 0 9 13 2
21 15 13 14 15 9 2 2 13 9 11 11 1 10 9 1 10 0 9 11 11 2
33 10 9 10 9 1 9 13 9 10 9 10 9 11 2 15 1 10 9 3 10 0 9 10 3 0 3 12 12 11 2 9 13 2
22 10 9 13 15 1 10 11 2 2 13 10 9 2 2 7 15 4 15 9 3 13 2
24 10 0 9 1 0 2 9 2 9 1 10 9 2 9 13 2 15 9 4 2 0 2 13 2
19 15 4 3 0 9 1 10 9 14 13 13 2 2 13 11 11 10 9 2
11 15 13 15 1 9 1 10 9 1 11 2
40 15 9 13 11 0 9 2 3 4 15 11 14 3 13 2 2 13 11 11 2 2 11 13 3 2 16 15 3 1 10 9 13 2 16 15 15 3 0 13 2
18 1 9 13 15 15 9 1 10 9 2 2 13 10 11 2 9 3 2
11 1 10 9 10 9 4 15 14 13 2 2
12 11 13 3 1 10 0 0 9 10 0 9 2
23 12 4 9 2 15 1 3 12 9 1 11 13 2 10 9 13 2 7 15 0 9 13 2
33 9 4 15 14 3 13 2 0 9 14 13 2 7 2 4 10 9 10 0 9 13 2 2 13 11 11 2 9 1 10 11 11 2
9 13 3 1 2 16 15 15 13 2
29 10 9 1 11 7 15 9 4 10 3 0 2 3 3 10 0 9 1 10 0 9 10 9 1 9 7 9 13 2
6 11 13 15 1 9 2
21 15 9 13 0 2 1 3 15 14 13 2 3 1 9 2 7 9 7 1 9 2
8 15 13 3 0 9 1 11 2
12 10 9 13 1 10 11 1 11 9 1 11 2
13 15 9 4 3 1 10 9 1 10 11 3 13 2
13 9 1 13 10 9 3 1 9 1 10 0 9 2
7 10 0 9 4 15 13 2
18 10 9 7 15 9 13 3 3 7 4 3 1 10 11 1 11 13 2
15 3 10 12 11 4 15 1 9 3 13 2 2 13 11 2
17 10 11 11 11 13 0 9 7 13 1 9 1 10 9 1 11 2
18 10 11 13 1 12 9 7 13 3 12 9 1 15 9 1 10 11 2
9 10 0 9 4 10 0 9 13 2
37 11 11 2 11 2 13 1 10 11 1 10 11 2 10 0 9 1 9 7 9 2 1 2 15 0 9 13 7 9 12 1 10 9 13 4 4 2
20 11 11 4 3 1 15 9 13 2 13 7 3 1 10 0 9 1 10 9 2
18 10 9 1 10 9 13 15 1 3 3 3 12 12 7 12 12 9 2
17 15 13 3 3 15 1 10 9 10 9 2 2 2 13 11 1 2
24 2 3 13 15 10 0 9 1 9 7 1 10 0 9 7 3 1 0 9 7 9 13 2 2
13 11 2 11 2 13 1 12 9 1 11 2 11 2
23 12 7 12 13 11 9 1 11 0 9 2 13 3 7 10 9 1 7 13 1 10 9 2
14 10 11 13 1 3 3 15 0 9 3 1 9 1 2
25 10 0 9 13 2 10 11 2 9 3 14 13 2 15 11 2 9 7 14 11 2 9 14 13 2
20 10 9 4 1 10 9 13 2 16 15 1 10 9 3 1 10 9 13 4 2
9 12 12 9 4 3 1 9 13 2
27 10 9 7 10 9 11 7 11 4 1 10 11 1 11 15 0 9 1 10 0 9 2 11 2 3 13 2
25 9 4 13 4 4 2 0 9 1 15 9 14 13 7 13 2 16 10 0 9 3 9 13 4 2
12 11 13 3 10 9 2 15 9 13 10 9 2
36 10 9 13 1 15 9 3 2 16 15 9 3 1 10 9 13 10 9 3 1 9 7 10 9 2 1 3 0 9 1 10 0 7 0 9 2
14 1 10 0 9 4 10 9 9 1 10 0 9 13 2
26 12 9 10 0 9 13 12 1 0 7 0 9 2 12 9 1 9 7 3 10 9 1 9 7 9 2
11 10 0 9 4 3 10 11 10 9 13 2
11 10 9 13 14 1 10 9 10 9 13 2
29 15 4 14 13 13 2 7 10 0 9 3 1 10 9 10 0 9 14 1 15 9 13 2 2 13 10 9 3 2
16 11 13 15 3 3 1 10 9 1 10 0 9 10 9 1 2
36 15 1 0 9 13 4 2 13 15 3 1 15 15 1 11 14 0 9 2 15 3 15 0 9 13 4 2 2 13 11 11 2 11 2 9 2
23 15 13 9 1 7 13 3 15 9 2 2 13 9 11 11 1 10 11 1 11 1 11 2
28 11 11 4 15 3 13 2 10 3 12 12 9 1 10 0 9 11 1 9 1 10 9 1 10 9 14 13 2
17 3 13 11 10 0 9 2 15 13 1 10 9 2 1 10 9 2
9 9 4 11 1 11 14 3 13 2
25 11 13 1 0 9 7 3 0 9 2 10 0 9 10 0 9 4 15 1 15 0 9 14 13 2
11 13 15 10 9 1 2 3 13 10 9 2
14 10 11 2 9 11 11 13 15 1 10 0 9 0 2
18 9 10 9 13 3 12 9 10 9 7 12 9 10 9 1 10 9 2
27 9 4 1 10 9 1 10 0 9 10 9 10 9 14 3 1 0 9 13 7 13 3 3 2 9 2 2
9 12 9 4 1 9 0 9 13 2
32 11 13 12 9 9 1 2 0 9 2 1 10 9 2 16 10 9 0 13 7 10 9 3 14 13 2 7 1 9 13 4 2
14 15 4 3 9 11 13 2 16 15 0 13 14 13 2
8 9 1 15 0 9 13 0 2
4 15 13 15 2
23 15 4 13 13 2 16 10 0 9 14 3 13 4 2 2 13 1 10 9 11 10 15 2
24 9 1 10 9 1 11 11 2 11 11 7 11 11 7 15 15 13 15 3 3 1 12 11 2
11 15 13 2 16 15 3 3 10 9 13 2
22 10 9 4 15 1 0 9 1 10 11 2 11 7 10 11 13 2 13 10 9 1 2
19 3 13 10 9 11 3 2 7 15 4 3 10 9 13 2 2 3 11 2
10 10 9 4 15 13 2 2 13 11 2
18 7 14 10 9 13 3 2 7 9 2 9 2 9 2 2 13 11 2
11 10 9 13 10 0 2 7 3 0 9 2
8 10 11 4 3 0 9 13 2
16 15 4 15 13 2 15 15 13 2 2 13 11 9 11 11 2
25 9 1 10 9 4 11 11 2 15 10 9 10 9 7 10 0 9 13 2 10 0 0 9 13 2
22 10 9 4 13 2 10 3 2 9 11 15 9 14 13 7 1 10 9 11 14 13 2
19 10 9 4 1 12 9 2 10 9 1 0 9 7 3 1 12 9 13 2
7 10 9 13 3 12 9 2
12 10 9 4 12 3 1 3 12 9 11 13 2
9 10 9 4 1 11 12 9 13 2
20 10 9 13 1 10 9 10 9 1 9 1 12 12 7 12 12 11 1 9 2
7 15 13 1 9 10 9 2
11 3 13 10 0 9 0 2 14 10 9 2
18 10 9 13 15 14 3 13 2 1 9 13 2 2 13 9 11 11 2
9 7 15 13 10 0 9 3 2 2
24 10 9 4 15 0 9 1 10 0 9 13 2 1 15 1 10 9 10 9 13 10 9 0 2
12 11 9 11 13 9 1 0 9 1 10 9 2
17 3 13 15 9 10 0 2 2 13 11 2 2 7 3 0 2 2
19 15 13 3 3 2 16 10 9 15 13 4 2 16 15 14 3 13 2 2
11 3 13 15 15 9 3 10 0 0 9 2
20 10 9 13 3 3 3 10 9 1 10 9 2 15 13 4 1 10 0 9 2
16 3 3 1 0 9 2 2 7 11 11 1 10 0 9 13 2
13 10 9 4 1 10 0 9 1 3 12 9 13 2
34 1 9 10 9 1 10 11 13 10 0 9 1 10 9 11 1 2 15 9 1 10 11 1 10 9 2 9 13 7 3 12 9 13 2
14 3 4 15 10 9 13 2 10 9 1 11 14 13 2
19 12 9 13 15 2 10 9 10 9 14 13 7 1 1 10 0 9 13 2
27 1 9 4 15 13 2 1 1 15 9 15 3 13 4 2 1 10 9 1 11 3 3 3 14 13 2 2
17 9 11 11 13 15 0 1 10 9 10 11 2 9 1 10 11 2
23 9 11 11 2 11 4 10 0 9 1 0 9 1 10 3 12 12 9 1 11 11 13 2
11 12 12 9 13 1 10 9 7 4 13 2
30 11 11 13 2 10 0 9 4 10 9 13 2 10 1 0 9 7 0 9 15 9 10 9 1 10 11 11 13 4 2
15 11 7 15 9 11 11 4 3 2 9 11 11 3 13 2
18 10 11 2 9 4 13 2 10 9 1 10 9 10 9 12 14 13 2
25 10 9 4 12 9 3 1 12 12 9 3 10 9 1 10 11 11 7 10 0 2 0 11 13 2
15 9 13 9 2 7 10 9 13 10 9 3 3 3 0 2
15 10 9 13 1 3 14 3 0 9 2 2 13 11 3 2
15 15 13 1 10 9 1 10 9 2 2 13 9 11 11 2
10 10 9 13 3 1 9 2 1 9 2
42 10 9 11 13 1 0 9 10 9 10 9 7 9 11 11 3 2 15 3 1 10 9 1 11 11 13 4 2 2 13 10 9 1 10 9 9 7 3 0 9 1 2
10 15 13 0 2 16 15 13 4 4 2
14 7 15 13 3 10 15 9 2 1 15 3 3 13 2
11 15 13 2 16 15 14 3 0 9 13 2
9 15 4 15 3 3 1 9 13 2
11 1 10 9 13 10 0 9 14 14 13 2
18 10 9 13 1 9 2 0 2 2 1 10 9 13 15 9 7 9 2
36 9 13 1 15 9 1 10 0 9 2 15 15 1 9 2 9 7 9 13 7 3 9 1 10 0 9 7 9 7 10 15 0 0 9 13 2
31 11 11 2 11 2 13 1 10 11 1 2 15 4 10 1 10 11 2 11 2 9 11 11 0 2 11 1 9 2 13 2
16 11 13 15 10 9 2 16 15 1 10 0 11 15 9 13 2
24 15 4 10 9 13 2 7 15 4 15 14 13 2 2 13 10 9 2 10 10 9 3 13 2
17 10 9 13 15 1 10 0 9 10 9 1 10 0 9 1 9 2
41 10 0 9 2 15 1 10 9 7 9 0 9 10 0 9 1 9 13 2 13 10 0 9 3 0 1 10 0 9 2 15 1 10 0 9 1 9 10 9 13 2
32 15 13 15 9 3 2 3 13 3 10 9 1 10 9 2 2 2 13 10 9 10 9 2 11 11 2 1 10 11 1 11 2
12 15 4 3 3 13 2 2 13 10 9 1 2
7 15 4 10 9 13 2 2
16 10 0 0 9 13 3 3 1 0 9 1 10 9 1 11 2
30 16 11 10 9 3 13 2 3 4 10 9 10 9 2 3 1 10 0 7 0 9 3 13 2 2 13 9 11 11 2
18 7 10 11 13 3 3 1 10 9 0 2 2 13 15 1 10 9 2
21 15 13 2 16 9 14 3 3 14 13 13 2 16 15 15 1 12 9 13 4 2
22 10 9 4 13 2 7 9 2 15 0 9 1 10 9 13 4 2 10 0 9 13 2
5 11 13 3 0 2
22 9 11 11 13 2 10 9 1 10 11 2 9 13 2 10 0 7 0 9 3 2 2
35 11 0 9 11 11 2 10 3 1 11 11 1 9 13 4 2 13 10 2 11 11 2 10 0 9 2 15 3 1 0 9 1 9 13 2
13 10 9 2 9 13 12 3 1 9 1 10 9 2
20 1 10 0 11 9 4 15 10 9 1 10 9 1 10 9 1 9 3 13 2
17 3 13 15 0 9 2 15 13 1 11 10 11 3 14 3 2 2
16 9 11 11 2 11 2 13 11 1 2 3 3 1 11 13 2
8 15 13 10 9 0 0 9 2
7 10 9 4 3 13 4 2
13 3 3 12 9 9 4 3 1 9 10 9 13 2
17 10 9 4 1 9 10 9 1 10 0 9 10 9 1 11 13 2
31 1 11 13 1 10 11 12 9 10 9 2 1 12 9 13 10 0 9 11 11 1 10 0 9 2 12 9 13 11 11 2
21 10 9 4 1 10 9 10 9 0 13 2 15 1 12 9 1 11 13 4 4 2
13 12 9 7 9 4 1 9 10 9 13 4 4 2
26 10 0 0 9 4 1 10 11 3 13 2 10 9 15 9 1 12 9 1 10 11 1 12 14 13 2
