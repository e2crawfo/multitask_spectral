564 11
13 7 16 0 15 9 13 15 13 15 7 13 1 15
9 13 3 9 15 6 6 7 6 6
7 13 0 15 7 13 9 15
11 13 3 15 0 3 3 9 15 0 0 13
13 15 3 3 13 15 13 1 9 15 7 13 9 15
7 9 15 13 9 13 15 3
16 3 13 15 9 1 9 3 9 7 9 13 3 9 13 7 13
4 0 1 13 15
6 3 13 16 3 13 13
11 0 3 13 13 7 13 13 7 13 13 15
7 7 3 15 13 15 15 13
7 0 3 13 15 1 0 9
14 7 13 9 7 13 9 7 13 9 7 13 15 9 0
6 7 3 13 15 1 9
8 7 3 13 9 7 13 9 15
6 3 13 9 7 9 9
4 11 3 13 15
10 3 13 13 9 7 9 7 13 9 0
3 7 13 15
5 9 13 15 9 15
12 13 3 9 13 15 7 13 9 13 9 0 9
5 9 13 7 3 9
14 16 3 3 3 13 15 9 7 9 13 15 7 9 13
5 9 9 15 13 15
5 7 13 9 13 0
7 7 13 12 1 12 9 15
2 0 13
12 16 3 3 3 13 0 9 15 1 15 13 15
12 3 15 3 13 13 7 9 9 15 13 1 15
14 15 3 13 13 15 3 13 13 7 0 15 3 13 13
18 0 3 15 13 15 1 9 13 15 3 15 1 9 15 15 13 1 9
22 7 15 3 13 12 1 0 0 9 0 9 3 1 9 9 6 13 15 3 13 9 15
14 6 15 13 9 15 1 9 15 7 13 9 15 1 15
5 13 15 7 3 13
10 11 7 11 3 13 1 9 0 3 15
21 13 9 15 1 15 7 13 15 1 15 16 0 13 7 13 9 7 13 9 9 15
8 13 15 16 9 3 0 13 3
3 3 13 9
9 13 9 15 1 15 7 9 9 13
18 0 9 13 15 1 15 13 7 0 9 7 9 13 15 1 15 3 13
6 9 13 1 15 9 13
6 3 13 7 9 0 0
19 7 13 15 1 15 9 0 7 16 13 1 9 13 7 15 9 1 9 13
5 1 15 9 13 15
29 13 3 9 9 0 7 9 3 13 7 9 15 13 16 3 13 9 7 9 13 7 9 13 7 13 15 7 13 15
25 7 13 1 0 9 0 13 13 9 7 13 15 7 13 9 3 13 7 13 0 12 0 12 0 12
4 9 3 13 15
4 15 9 13 15
14 7 1 9 15 13 7 15 15 13 13 7 13 9 0
4 13 15 6 9
9 7 9 15 3 15 3 1 15 13
4 13 3 15 11
11 7 13 11 13 3 1 9 1 0 9 12
4 0 3 13 15
9 9 3 13 1 9 9 13 15 9
11 9 16 15 13 13 15 13 1 15 1 9
9 1 15 15 13 9 0 1 9 15
5 7 13 9 13 15
5 13 3 11 13 15
10 7 6 9 0 1 9 0 13 13 13
4 0 3 13 13
17 7 13 15 16 9 13 15 13 0 13 0 0 7 0 13 0 13
4 12 7 3 9
2 7 3
11 13 3 11 1 9 11 0 13 9 15 13
5 7 13 11 13 15
6 0 3 13 15 13 11
3 6 13 15
9 7 13 9 13 0 7 13 15 3
7 11 3 13 3 7 13 15
3 3 13 15
2 7 13
7 15 3 0 13 1 9 0
15 16 3 9 15 7 9 15 13 15 13 15 7 13 1 15
13 3 13 9 1 9 15 0 16 13 12 1 0 0
6 3 13 1 15 11 13
11 13 3 9 9 0 13 15 7 9 13 15
13 7 13 15 9 15 13 15 9 16 13 15 9 15
11 7 13 15 9 15 7 13 12 1 9 12
12 16 3 13 9 9 1 9 0 13 3 13 15
22 10 3 13 3 9 13 3 13 3 9 13 13 9 7 9 7 13 0 15 3 0 15
17 3 13 15 16 0 13 9 1 9 0 13 3 0 1 9 0 13
28 15 13 1 15 1 9 3 13 9 0 1 9 9 15 13 3 15 1 12 1 12 9 13 12 1 12 9 0
11 1 12 3 1 12 9 13 13 0 13 0
9 7 13 15 9 13 1 0 1 0
8 13 3 0 0 13 3 3 15
2 15 13
9 3 3 9 15 15 13 15 13 15
16 13 3 11 13 15 9 15 7 3 13 15 9 7 1 15 13
22 13 3 9 7 13 15 13 15 11 13 9 7 9 7 13 1 9 15 7 13 1 15
2 13 13
7 3 3 13 15 1 9 13
14 7 3 13 1 9 13 1 15 13 9 7 9 0 13
2 3 13
5 3 3 13 15 13
11 13 3 11 9 9 0 7 3 13 15 9
10 9 15 9 13 13 0 13 1 9 9
4 6 9 15 13
18 7 13 9 0 1 9 13 15 15 13 0 3 7 0 7 13 9 13
9 7 13 1 15 9 15 1 9 13
4 0 3 13 15
21 13 3 1 15 12 9 7 0 13 15 13 7 3 13 9 13 3 9 15 9 15
5 13 9 0 7 0
7 13 3 9 13 15 11 13
4 13 3 9 15
11 7 15 13 15 13 15 7 13 15 13 15
6 0 7 0 15 0 13
8 0 3 13 13 7 0 3 13
6 7 15 13 9 9 15
6 3 13 13 15 16 13
2 13 15
18 13 3 9 1 9 7 9 1 9 7 13 9 7 9 7 9 1 9
17 3 3 9 13 1 9 7 13 15 1 9 3 13 3 9 9 0
17 7 1 9 0 7 1 9 0 15 3 13 7 9 0 3 9 12
15 0 1 3 15 13 0 16 1 15 3 13 9 9 0 13
8 13 3 9 13 15 15 7 13
17 13 3 15 13 13 9 7 0 13 1 15 1 9 7 13 13 9
11 7 13 12 13 13 9 7 13 9 9 15
6 9 12 9 15 13 13
6 13 3 9 15 13 15
7 9 3 15 13 13 7 13
8 13 3 15 7 3 13 15 13
11 7 13 0 1 9 0 7 9 1 9 0
5 13 3 11 13 15
6 0 3 13 15 12 9
9 9 3 13 13 1 12 1 12 9
6 13 3 11 13 15 13
9 7 13 9 7 9 13 13 15 13
11 7 13 11 7 12 9 0 13 13 7 13
6 9 3 0 7 9 0
1 13
4 11 3 13 15
11 3 1 9 3 13 1 9 7 9 13 15
5 7 13 9 13 15
7 3 9 13 9 15 13 16
5 11 15 13 13 15
10 7 13 15 13 7 13 15 0 11 9
11 0 3 13 15 9 0 9 9 1 0 9
4 3 13 15 11
8 3 3 13 3 1 9 15 1
3 9 13 15
8 11 3 13 13 15 16 15 13
13 13 3 15 13 9 15 13 9 7 13 13 15 3
9 3 13 3 1 9 7 9 13 15
6 1 9 0 9 0 13
4 1 12 9 13
5 7 6 9 13 0
5 13 9 3 13 11
4 3 13 15 11
10 7 13 15 9 0 1 9 1 0 9
3 13 9 0
17 7 3 13 1 9 7 13 13 15 9 7 9 3 9 13 1 15
1 13
4 15 3 13 0
16 7 3 9 3 13 13 11 7 13 1 0 9 7 3 9 13
1 13
9 7 13 1 15 13 13 9 13 12
17 7 16 13 16 9 13 9 0 13 1 9 9 7 13 13 15 13
6 7 13 1 9 15 13
14 1 15 9 0 7 9 13 15 7 15 9 3 13 15
12 7 13 15 16 1 9 13 15 16 1 15 13
14 7 3 13 9 1 9 9 13 1 15 3 15 13 13
16 7 11 0 7 11 9 0 3 13 15 9 11 15 13 9 0
12 7 16 9 1 15 13 15 3 13 13 9 0
4 7 13 15 13
4 7 13 3 13
7 15 13 13 13 0 9 0
18 7 9 9 0 7 9 9 7 1 0 9 13 13 9 7 1 9 13
10 7 0 9 0 13 15 9 3 13 13
3 7 13 15
11 15 3 13 0 16 7 9 7 9 13 15
4 15 15 13 9
6 7 13 13 15 13 13
5 9 15 1 9 13
6 13 9 13 15 7 13
3 15 13 9
9 3 0 13 0 7 15 9 13 15
50 7 13 12 1 12 7 13 15 13 12 7 12 7 13 15 9 1 9 0 7 13 15 16 15 3 13 1 9 3 9 12 7 9 7 9 7 1 9 9 7 13 1 9 7 3 13 15 1 12 9
6 15 15 13 11 0 13
9 15 3 13 13 15 1 9 9 15
23 0 3 13 13 15 1 9 7 13 9 15 1 9 7 13 15 9 7 9 13 15 9 15
19 7 3 9 0 13 13 1 15 9 15 13 16 0 13 9 7 3 9 13
3 7 13 13
13 7 9 13 13 9 1 9 9 7 0 12 1 9
8 1 0 3 13 15 9 7 9
6 13 9 15 7 9 15
13 7 3 13 1 9 1 9 13 15 9 15 1 9
9 7 13 15 16 13 9 1 9 15
16 7 3 13 11 1 9 0 7 0 13 1 9 0 1 9 0
18 1 0 9 3 0 13 9 7 3 13 15 13 13 9 15 11 13 15
20 7 13 9 13 1 9 7 13 12 10 9 9 13 13 7 13 9 15 16 13
5 7 13 9 15 13
1 12
7 7 13 15 1 9 15 13
3 15 13 11
13 15 3 3 13 9 15 15 1 7 9 0 13 15
3 0 3 13
6 11 3 13 3 13 15
9 7 9 13 7 13 9 15 7 13
3 0 3 13
10 0 3 3 13 9 7 13 15 13 15
4 13 15 11 13
8 7 16 9 15 13 15 13 15
5 0 3 13 13 15
3 7 13 15
13 15 3 3 13 9 0 3 9 3 13 13 1 15
2 3 13
5 13 3 13 9 0
11 7 1 15 13 11 7 11 9 0 13 15
1 13
17 3 9 0 3 13 16 13 15 7 13 7 13 9 15 9 1 0
1 13
4 9 15 13 15
2 13 15
24 7 13 9 3 13 9 13 16 3 13 1 15 15 7 13 1 15 15 3 13 1 15 3 9
11 7 13 9 7 9 7 13 3 15 13 13
10 9 0 3 13 1 9 3 7 1 9
5 7 13 15 9 13
4 13 15 9 15
10 9 15 9 13 13 0 13 1 9 9
5 13 3 7 3 13
5 7 13 15 1 15
6 12 3 15 13 15 9
5 11 3 13 15 16
6 0 3 11 13 15 9
18 15 3 1 9 15 13 7 0 1 9 15 15 15 13 13 15 9 15
13 0 3 13 1 15 9 13 16 15 13 7 0 13
8 3 15 3 13 13 7 9 0
14 7 3 16 13 15 15 6 3 11 6 3 3 13 9
13 6 13 15 16 3 13 13 9 0 16 15 0 13
8 13 3 9 7 9 1 12 9
3 7 13 15
2 9 13
2 7 0
4 0 13 9 15
9 7 1 0 3 13 13 15 1 11
6 13 3 16 13 13 15
5 3 13 12 9 13
2 13 9
2 9 9
5 15 0 1 15 13
4 15 15 15 13
10 7 13 15 9 3 13 13 1 13 16
12 3 16 9 3 13 12 9 13 15 15 12 9
4 3 13 3 15
6 11 3 3 13 13 15
12 7 13 15 1 9 7 13 1 15 13 0 9
13 7 13 7 13 9 15 13 9 1 15 15 15 13
9 3 13 16 13 16 13 11 13 15
25 7 13 9 7 13 15 13 15 1 9 7 13 1 9 15 13 13 1 9 7 13 9 1 9 9
3 3 13 15
17 13 3 11 3 1 0 9 13 15 1 11 9 1 15 13 12 9
5 9 3 13 0 13
11 13 3 15 15 9 0 13 1 0 9 0
5 7 13 9 13 15
30 1 0 3 9 13 13 9 11 1 9 1 9 0 15 9 11 1 9 13 9 15 9 11 1 9 0 7 9 9 11
3 6 9 0
11 7 0 15 9 13 16 13 9 13 1 9
8 13 13 0 7 13 15 13 0
9 13 3 9 15 3 13 13 13 15
7 7 15 9 9 0 13 15
4 7 13 15 9
10 13 3 13 1 9 13 15 1 9 0
32 3 13 9 15 9 1 9 15 1 9 16 13 9 15 9 15 15 13 13 1 9 15 9 9 1 9 9 7 9 9 15 11
4 15 16 13 15
4 0 13 9 15
7 3 3 9 1 9 9 13
5 15 0 13 15 13
27 11 3 9 13 15 1 11 9 9 15 7 1 15 0 15 13 11 13 3 0 1 15 7 13 11 1 9
7 7 13 15 9 1 9 0
8 16 9 13 0 13 15 3 3
10 9 0 1 15 15 1 13 15 13 0
12 7 13 15 1 9 15 16 1 9 13 9 15
13 7 13 15 9 1 9 13 1 15 3 3 13 15
10 13 3 3 9 1 0 13 7 13 16
21 13 3 1 12 1 9 15 13 0 13 15 1 9 13 3 7 13 13 1 9 9
8 13 1 15 16 9 0 13 9
1 13
6 7 13 9 15 13 15
2 15 13
9 13 3 9 3 13 13 1 15 9
18 13 3 1 9 0 13 15 1 9 7 13 9 15 9 7 13 13 9
6 7 13 9 13 0 9
14 0 3 13 15 9 7 13 15 1 15 15 13 13 11
7 13 15 1 0 9 7 13
4 0 13 13 15
13 7 16 1 9 13 1 15 13 13 15 15 9 13
8 0 3 9 15 13 13 15 15
4 7 3 13 15
4 9 3 13 15
7 3 1 11 0 9 3 13
3 9 15 13
7 15 3 13 13 7 15 13
11 6 10 1 9 0 7 9 13 1 0 13
12 7 15 9 13 3 9 13 9 13 15 9 0
9 6 9 9 7 9 9 9 7 9
4 13 3 0 9
3 13 3 15
15 7 3 13 0 13 1 9 7 13 13 7 9 0 13 15
4 13 3 9 0
19 15 3 13 13 15 15 7 15 3 13 3 15 13 15 13 13 15 1 15
4 13 3 15 13
13 15 3 0 13 16 7 9 13 7 9 7 13 15
5 13 3 15 11 13
21 7 13 1 9 0 13 15 13 1 9 15 16 9 0 13 15 16 12 1 12 9
4 13 15 15 15
6 11 3 13 13 15 13
12 0 3 13 15 3 7 13 15 1 9 13 13
9 13 3 13 1 9 13 7 13 3
7 13 3 12 1 12 13 15
19 13 3 12 9 7 12 9 13 1 9 13 15 7 13 7 13 9 13 9
32 0 3 13 15 13 15 3 13 0 13 16 13 9 0 3 13 7 13 13 1 9 7 9 7 9 7 13 13 7 0 9 13
11 7 3 13 9 13 15 11 12 7 0 13
5 13 15 9 15 3
15 11 3 13 9 9 15 13 9 13 15 1 15 7 13 15
9 7 13 13 1 9 0 16 13 15
4 13 3 1 0
5 13 3 1 15 11
3 9 9 0
10 3 0 13 16 13 15 1 15 9 0
7 7 13 15 1 9 12 13
3 13 3 15
13 13 3 15 1 15 9 13 15 1 9 7 13 15
9 9 15 9 11 13 15 1 9 15
17 7 13 13 15 1 9 15 13 15 16 13 13 15 9 15 1 15
11 7 3 13 15 1 9 7 13 15 1 9
19 16 3 3 13 15 13 16 13 9 15 7 1 9 15 13 13 15 15 13
8 7 13 13 9 7 0 13 0
13 13 3 3 13 0 13 9 15 9 1 9 13 15
8 9 0 13 1 9 1 9 0
12 9 3 13 13 15 16 3 3 13 15 1 9
6 9 0 13 3 15 13
6 0 3 13 7 13 13
3 6 13 15
11 7 0 15 13 9 1 9 0 13 15 15
6 13 3 9 1 15 13
4 0 1 13 15
20 16 3 3 9 3 1 9 13 7 3 1 9 13 9 3 13 3 3 15 0
20 7 15 0 9 13 9 15 3 13 15 1 9 16 13 7 13 3 13 15 15
17 15 3 13 0 9 7 0 15 13 9 1 9 15 13 1 9 9
8 13 3 16 9 13 13 1 9
2 13 15
4 13 3 0 9
9 16 3 3 3 1 13 9 13 15
4 15 13 9 0
4 7 13 13 15
13 7 6 13 0 15 13 0 7 13 0 15 13 0
5 0 13 1 9 0
12 13 3 1 13 9 13 3 9 13 13 1 15
19 7 3 13 9 13 0 9 0 0 7 0 13 16 3 13 0 15 13 15
2 13 15
8 3 13 15 9 9 13 9 15
5 13 9 13 3 13
9 13 15 1 15 16 13 9 15 13
15 7 13 13 9 15 1 9 15 13 9 7 15 3 13 15
22 3 3 15 3 13 13 15 9 15 7 0 15 13 7 13 13 1 9 15 7 13 15
6 7 13 12 1 9 13
11 9 15 3 1 15 13 7 15 15 15 13
3 13 3 13
6 7 1 0 3 0 13
10 3 15 13 1 9 0 9 1 9 13
17 7 1 9 13 9 15 13 1 9 13 11 3 7 11 1 9 15
4 13 3 15 11
22 0 15 13 13 16 13 9 0 13 1 9 15 7 13 1 9 3 16 13 0 0 12
14 15 3 1 15 9 13 13 7 13 15 13 1 9 13
4 11 9 13 15
2 13 13
2 6 3
4 13 12 3 13
11 9 3 13 1 9 0 7 13 1 15 13
17 13 3 7 1 15 13 15 1 15 16 13 9 7 13 0 9 0
2 13 15
6 7 13 15 15 9 13
6 13 9 15 7 9 15
13 0 3 13 9 1 0 9 13 3 0 1 9 13
8 13 3 12 1 12 13 1 15
4 9 15 13 15
8 3 3 13 15 1 9 15 13
14 9 15 0 9 13 1 9 3 13 15 9 7 13 15
11 16 1 0 0 13 13 9 13 1 12 9
7 1 9 15 13 15 0 9
20 3 9 15 0 3 13 15 16 9 13 13 1 15 13 3 7 13 15 1 15
7 0 3 13 16 9 13 15
12 7 16 13 15 13 9 13 15 1 15 13 16
10 16 3 13 1 9 9 15 9 13 15
5 7 13 0 13 9
1 13
7 0 13 1 9 0 13 15
3 13 15 9
6 7 0 13 9 13 0
20 7 16 13 0 3 11 13 1 9 3 13 9 9 0 7 9 0 7 9 0
11 13 1 0 15 16 13 9 15 9 9 15
6 3 13 3 1 9 15
18 15 3 13 15 9 7 9 15 3 13 13 15 7 13 15 13 15 15
12 7 3 13 9 0 1 9 1 9 7 9 0
20 13 3 1 0 9 13 15 16 13 15 13 15 0 13 13 7 13 1 9 0
6 13 13 15 9 16 13
3 7 3 13
10 7 13 9 9 13 13 7 13 15 13
10 9 9 13 15 7 13 15 9 13 15
3 13 3 15
8 7 13 13 1 9 1 9 0
11 7 13 9 15 3 3 9 9 13 1 9
10 13 3 3 15 13 1 15 13 13 15
10 13 3 15 13 7 13 15 1 9 0
2 9 13
8 7 9 13 11 13 15 15 13
9 3 13 9 0 13 1 0 9 0
21 13 3 13 1 0 9 13 16 13 0 1 15 7 13 15 9 15 13 1 15 13
3 7 7 11
1 13
19 13 3 1 9 15 0 9 9 9 7 9 15 7 13 15 7 13 15 15
11 13 3 1 11 3 15 12 9 1 15 13
13 13 3 15 15 3 9 13 7 9 13 15 7 13
6 7 0 15 0 3 13
4 7 0 13 13
18 7 13 9 15 7 13 15 1 9 13 15 0 12 1 12 7 15 0
9 13 3 15 15 9 11 13 1 15
18 7 13 15 1 15 1 9 7 13 3 3 7 9 13 0 3 3 13
8 0 3 13 15 9 7 13 15
2 15 13
5 13 3 15 0 3
12 15 3 13 1 9 0 16 13 15 9 1 3
4 15 13 1 9
2 15 13
6 13 11 15 13 13 11
14 15 13 11 1 9 7 9 13 11 9 0 15 1 11
5 13 11 7 13 15
13 3 13 9 13 7 9 0 13 7 13 1 9 0
16 13 3 3 9 0 12 13 1 9 0 13 1 12 7 12 9
17 13 9 9 11 1 11 0 7 13 9 15 7 13 1 15 9 15
5 13 11 7 13 15
2 13 11
5 13 11 7 13 15
14 7 3 13 3 13 13 16 3 13 1 9 0 9 0
7 7 13 1 11 7 13 15
5 13 3 1 15 13
6 13 3 15 13 1 11
11 3 15 9 13 1 15 13 13 9 9 13
5 13 11 7 13 15
18 9 9 13 15 16 13 9 3 7 1 9 0 7 1 11 13 15 9
5 15 13 13 1 15
5 0 3 13 1 15
14 1 0 3 13 9 0 16 15 13 13 7 15 13 13
13 0 3 13 7 13 16 0 13 1 9 9 9 11
10 16 9 7 9 3 13 3 13 9 13
7 3 1 9 0 13 15 9
13 0 13 11 13 7 13 16 0 9 3 13 13 15
8 1 0 3 13 15 11 1 9
4 6 6 13 15
11 7 9 13 15 3 9 13 16 9 0 13
6 15 3 13 9 0 0
8 16 15 13 1 9 15 0 13
6 13 3 1 9 9 0
3 13 3 11
18 11 3 13 16 13 13 16 13 15 7 13 9 13 3 1 9 0 12
6 15 13 16 13 9 0
16 3 11 13 15 9 1 9 7 9 15 13 15 9 0 1 9
24 0 3 13 9 9 15 16 0 13 9 7 13 1 15 13 9 0 7 13 15 15 1 0 9
4 13 13 1 9
14 0 13 9 13 1 9 16 16 1 15 15 13 3 13
12 9 3 15 0 13 9 7 9 15 0 13 9
4 0 3 15 13
6 13 3 11 12 1 12
11 9 15 3 3 13 7 9 15 3 13 0
8 7 9 0 13 1 15 1 9
18 16 15 13 9 15 13 13 1 9 15 1 9 13 7 15 1 15 13
7 12 9 13 7 15 13 15
8 13 3 1 9 13 11 7 13
13 13 15 7 3 13 7 3 13 15 15 3 13 13
13 3 3 3 13 9 0 13 16 11 3 3 13 13
11 13 3 9 1 9 7 9 7 13 15 0
4 15 3 15 13
5 15 3 15 3 13
5 15 1 15 0 13
3 13 3 15
3 13 3 9
3 13 3 15
11 3 13 15 12 9 16 15 0 13 15 3
5 6 6 13 15 16
7 15 3 1 9 13 7 13
11 16 3 9 13 1 15 15 3 13 9 15
4 6 6 13 15
9 16 15 13 15 0 9 15 15 13
4 6 6 13 15
7 13 9 3 15 3 13 13
2 15 13
1 13
14 3 3 3 13 3 13 7 15 15 13 9 15 3 13
3 13 9 9
7 3 3 15 13 9 15 13
12 16 3 13 1 9 13 0 3 13 13 13 15
3 0 3 13
1 13
5 13 3 15 3 11
25 7 9 15 13 9 15 3 13 9 15 13 9 13 7 13 9 7 13 7 9 13 15 7 13 9
4 3 9 15 13
8 13 3 3 9 9 16 15 13
32 16 0 13 0 1 15 13 9 0 7 3 13 15 9 13 15 9 13 7 13 1 9 15 13 16 13 16 13 16 9 0 13
15 13 3 11 13 9 9 7 13 9 9 15 15 9 11 13
12 9 3 13 15 9 13 9 7 3 3 13 3
6 11 3 13 1 9 15
9 11 3 3 13 16 11 13 13 15
5 15 13 9 7 9
3 13 3 9
3 0 3 13
8 7 13 13 13 9 7 9 9
21 15 3 13 15 7 13 16 0 13 15 16 12 9 13 1 9 7 3 15 9 13
8 11 3 12 13 1 13 1 15
11 0 3 1 15 3 13 7 15 3 3 13
17 13 3 9 15 13 1 15 3 11 13 1 9 7 13 15 1 0
7 7 3 11 7 11 13 11
9 3 15 1 9 0 13 7 15 1
8 3 1 0 9 9 1 15 13
11 0 13 11 3 13 9 15 7 13 1 15
9 9 15 13 0 13 15 1 0 9
5 13 11 7 13 15
6 13 3 13 3 9 13
17 16 3 15 13 15 9 9 7 9 3 15 0 13 15 15 13 9
4 6 6 13 15
5 3 13 13 3 11
3 9 3 13
6 3 3 13 15 15 9
7 15 13 9 7 9 7 9
3 13 15 9
9 7 16 15 13 1 9 15 15 13
10 13 9 15 7 13 15 0 13 13 15
3 9 13 15
18 15 13 1 15 7 15 1 15 13 9 0 16 1 15 3 13 13 15
10 15 9 15 13 16 13 15 15 13 15
5 13 9 0 9 15
3 13 15 3
2 3 13
10 3 0 13 13 15 7 3 13 13 3
2 13 3
17 3 3 13 9 1 0 3 13 9 1 9 16 13 15 9 1 9
12 7 15 12 13 7 13 12 16 9 1 15 13
19 7 3 13 15 15 9 1 15 0 9 15 13 3 16 3 13 9 1 15
30 3 13 1 15 1 9 15 13 15 1 9 15 15 13 13 15 13 7 15 1 15 3 13 3 9 0 16 13 15 9
16 7 15 9 15 13 13 15 13 15 16 13 12 3 3 15 12
2 15 13
2 11 9
4 13 9 1 9
9 13 15 15 7 1 9 15 13 15
16 15 1 0 13 15 7 1 0 13 1 15 9 16 13 1 9
4 13 3 11 9
2 6 9
3 3 13 15
6 16 0 13 13 9 9
2 13 15
3 13 3 13
9 13 3 9 3 0 1 9 13 15
5 7 13 9 13 9
3 7 13 11
10 13 3 11 7 0 9 7 13 1 9
7 16 3 13 15 13 1 9
8 0 3 13 16 9 13 13 15
13 13 1 9 15 7 9 15 7 9 15 7 9 15
7 7 0 13 13 7 13 15
2 9 15
7 3 13 3 9 16 11 13
18 11 3 11 13 16 9 13 9 13 15 13 3 0 7 13 15 1 9
1 13
4 13 15 3 3
