600 11
12 9 13 16 1 9 12 9 15 14 9 13 2
26 9 15 13 16 9 1 10 9 9 13 2 10 9 13 16 1 9 16 1 9 15 13 2 9 13 2
12 9 2 1 9 9 1 9 9 9 9 13 2
21 9 12 9 1 12 9 9 7 9 9 13 16 1 9 9 15 1 9 9 13 2
43 9 16 9 9 1 9 13 16 15 14 1 9 13 2 1 9 9 9 7 9 9 7 9 2 10 9 1 9 15 14 0 13 2 16 0 13 9 9 9 9 13 13 2
53 10 9 14 4 13 16 9 9 0 13 2 7 9 1 9 9 15 7 9 1 9 2 9 1 9 1 9 0 13 2 7 1 12 12 9 10 0 16 9 9 13 9 13 2 7 9 9 14 1 3 13 13 2
16 10 9 1 9 9 0 1 9 1 9 7 9 14 9 13 2
43 1 9 9 7 9 1 9 9 13 16 9 15 13 13 2 13 7 13 1 15 9 13 9 7 13 1 9 2 16 15 10 9 13 16 15 1 15 1 9 13 13 13 2
2 13 2
56 15 16 9 9 1 15 13 16 9 0 13 7 1 9 15 9 13 2 16 9 7 9 7 9 2 7 15 9 16 9 13 16 1 9 7 9 1 9 7 9 1 9 13 2 9 13 1 15 16 9 0 1 9 15 13 2
11 1 9 9 9 7 9 16 10 9 13 2
9 13 2 13 7 13 1 15 9 2
22 3 9 0 13 7 9 0 15 9 0 1 15 13 16 4 13 7 15 14 9 13 2
8 9 1 9 9 0 9 13 2
30 9 16 1 9 9 7 9 13 2 1 9 9 0 9 13 2 3 13 4 9 0 2 16 9 9 9 13 1 9 2
17 9 0 7 9 0 1 9 2 0 15 16 9 0 13 1 9 2
15 15 9 1 9 9 13 2 15 9 0 9 7 9 13 2
13 1 9 9 13 3 2 9 1 9 15 13 3 2
14 9 0 9 13 3 2 9 1 9 7 9 13 3 2
15 13 16 0 9 13 16 9 2 3 1 9 13 9 9 2
13 13 3 9 9 15 2 0 13 9 1 9 15 2
16 3 13 16 9 3 13 3 2 1 1 9 1 3 13 3 2
11 16 15 2 9 1 9 9 15 15 13 2
35 1 12 9 9 0 9 2 16 9 0 14 10 9 9 9 13 2 4 1 9 9 0 1 9 7 9 14 1 9 15 1 9 0 13 2
29 9 9 9 0 1 15 13 16 9 9 9 1 9 13 13 16 9 0 1 7 2 3 9 12 9 14 9 13 2
10 9 9 7 9 9 1 9 13 13 2
19 10 9 0 9 1 9 9 0 13 7 15 9 13 16 1 15 9 13 2
33 9 7 9 16 3 9 0 1 9 9 13 2 7 9 3 9 7 9 7 9 9 0 15 13 2 9 15 14 1 9 4 13 2
25 9 16 9 1 9 1 9 13 2 1 9 9 13 16 1 9 9 7 10 9 0 9 13 13 2
17 16 1 9 15 3 9 13 2 1 9 1 15 9 7 9 13 2
15 9 0 7 9 0 2 1 9 7 1 9 15 3 9 2
12 9 9 1 9 9 2 9 9 1 9 9 2
16 9 13 3 1 9 15 0 2 3 0 13 1 9 15 0 2
15 9 7 9 7 9 7 9 2 3 0 1 9 13 9 2
39 2 9 9 9 9 2 9 12 2 16 9 9 9 16 12 9 0 13 2 0 13 1 9 0 2 13 9 3 9 2 1 9 9 7 9 7 9 13 2
36 7 2 3 9 7 9 7 9 0 2 13 13 9 1 9 2 9 9 9 12 7 12 2 9 9 9 1 9 1 9 9 9 15 14 13 2
41 15 9 13 16 1 9 9 0 2 1 3 7 3 2 10 9 9 1 9 13 2 7 9 9 13 1 9 9 2 10 9 16 0 9 0 7 9 0 15 13 2
38 0 1 9 9 13 16 3 9 9 9 1 9 0 9 14 0 13 7 9 9 9 9 0 13 13 2 16 9 9 9 14 1 9 9 9 0 13 2
14 7 3 9 9 9 1 9 9 12 1 12 9 13 2
5 9 7 9 2 2
23 9 9 9 9 9 9 1 9 9 0 9 1 9 9 9 7 9 1 13 7 13 13 2
23 9 15 14 13 2 9 9 9 0 13 16 0 1 9 9 0 9 1 1 9 9 13 2
38 10 9 0 1 0 9 0 1 9 12 1 3 9 13 1 7 1 0 9 2 9 0 9 12 9 9 0 15 2 0 1 9 9 1 9 9 13 2
24 9 0 9 9 7 1 1 15 9 0 7 9 0 1 9 1 9 9 9 9 0 13 13 2
21 9 9 9 9 15 13 16 9 0 7 9 3 1 0 0 16 9 9 0 13 2
36 9 9 9 9 1 0 0 0 1 9 9 7 9 7 3 9 0 9 0 13 1 7 9 13 9 0 0 15 14 1 12 9 0 9 13 2
19 9 9 9 1 9 9 3 9 13 16 9 9 9 9 14 0 9 13 2
30 9 9 9 9 9 14 1 9 10 9 0 7 9 0 0 13 7 9 9 1 9 0 9 7 9 0 9 0 13 2
12 9 0 9 12 9 0 1 9 9 9 13 2
28 9 0 9 9 9 1 9 9 0 1 9 7 9 1 9 0 9 1 9 9 9 14 1 9 0 0 13 2
25 15 16 9 9 9 1 9 0 9 13 9 0 9 1 9 0 0 3 9 7 10 9 0 13 2
18 9 10 9 1 9 0 9 0 0 13 16 3 15 9 0 9 13 2
10 3 9 0 1 10 9 0 13 13 2
31 9 9 13 9 9 9 9 1 9 9 9 1 1 9 9 7 9 9 0 0 15 1 9 15 2 9 7 9 2 13 2
39 1 9 15 7 9 0 0 9 13 7 9 9 13 7 9 16 1 0 9 9 0 13 2 16 10 12 9 1 1 9 1 9 9 9 2 9 0 13 2
57 9 0 13 16 9 9 9 1 9 12 16 1 9 9 9 7 9 0 13 12 9 0 0 1 9 13 16 1 9 9 9 16 9 0 9 7 9 16 1 9 13 9 9 0 14 1 9 0 1 9 9 9 13 2 9 13 2
28 16 9 0 9 7 9 1 10 9 1 9 9 7 9 7 9 3 13 7 9 0 15 1 1 9 9 13 2
25 9 9 9 1 9 9 0 3 9 7 9 16 1 9 0 7 0 1 9 0 13 3 9 13 2
27 16 0 9 0 2 0 9 9 0 7 9 0 7 9 0 13 7 3 1 10 9 1 9 9 1 13 2
11 16 0 0 10 9 9 2 9 4 13 2
54 1 1 9 9 7 9 9 1 9 2 9 0 13 16 12 1 9 9 9 7 9 0 9 1 9 16 9 0 13 16 9 13 1 9 9 9 7 1 9 1 9 9 9 0 1 9 7 15 1 9 9 0 13 2
38 1 1 10 9 2 9 9 9 7 9 15 1 9 1 9 9 7 9 9 12 9 0 1 9 13 7 9 13 16 3 1 12 9 1 9 9 13 2
14 16 1 12 9 0 7 0 9 0 1 15 9 13 2
16 9 9 9 1 9 9 1 9 0 9 9 1 9 0 13 2
54 16 9 9 9 9 14 1 9 9 0 9 9 0 7 9 0 7 9 9 1 9 0 7 9 15 13 2 9 0 9 13 7 3 16 9 9 9 9 9 9 9 0 7 0 7 0 13 2 0 9 14 9 13 2
13 16 4 12 9 0 7 0 1 15 9 0 13 2
14 15 9 1 9 7 9 9 9 0 7 9 15 13 2
19 9 15 13 2 10 9 9 1 9 0 7 9 9 1 1 9 9 13 2
23 16 9 9 9 0 1 9 13 2 16 9 9 0 13 9 9 9 13 0 7 0 13 2
23 3 1 3 9 0 9 9 9 3 3 9 2 12 9 0 13 16 9 9 14 0 13 2
29 1 9 9 9 16 9 0 7 7 0 13 0 13 9 13 7 7 9 9 0 13 9 14 1 0 0 9 13 2
21 16 1 9 9 9 7 9 9 2 0 9 1 9 9 0 2 0 7 0 13 2
22 9 1 1 0 9 1 9 9 9 3 9 9 0 1 1 9 9 0 9 13 13 2
20 0 13 16 9 1 1 9 9 0 7 9 15 16 0 15 9 13 0 13 2
25 9 0 3 9 9 16 1 9 9 7 7 9 0 0 15 2 12 9 0 1 9 0 9 13 2
51 16 15 1 10 9 1 12 12 9 0 1 10 9 9 13 7 9 0 9 1 9 15 14 9 9 7 9 13 2 9 0 7 9 14 16 1 9 0 0 1 12 1 12 9 9 9 0 13 9 13 2
30 1 1 9 1 9 9 9 0 9 13 9 9 14 1 9 3 13 7 1 9 9 9 9 9 7 9 14 9 13 2
20 16 3 0 7 0 13 16 9 1 9 16 3 1 9 12 9 13 0 13 2
15 1 9 12 0 0 13 16 10 9 1 12 9 13 13 2
23 10 9 4 9 13 13 1 7 9 1 9 13 16 9 9 1 9 7 9 0 0 13 2
18 1 0 9 1 9 9 9 7 9 9 9 9 1 9 15 9 13 2
15 9 9 9 1 9 7 9 2 9 15 15 14 9 13 2
12 7 1 9 0 15 2 9 9 7 9 13 2
16 1 9 0 9 15 9 13 2 3 15 14 9 9 9 13 2
19 9 13 1 15 6 9 0 2 9 15 1 9 9 15 2 3 0 13 2
14 9 9 9 15 13 2 9 1 3 9 9 9 13 2
21 6 0 9 2 9 15 9 16 3 2 9 7 9 2 1 9 15 1 9 13 2
21 1 9 15 7 15 13 9 1 9 9 2 9 15 1 9 9 7 9 9 13 2
16 9 15 9 9 13 2 16 1 9 9 13 9 2 0 13 2
15 1 9 9 9 15 9 13 2 9 9 9 9 9 13 2
13 9 0 9 9 13 9 9 14 1 9 3 13 2
14 0 9 9 1 9 0 9 9 1 1 9 0 13 2
24 9 1 9 0 9 16 1 9 1 9 9 13 13 2 9 0 1 9 9 0 1 9 13 2
24 1 10 9 2 9 9 9 1 9 9 13 7 9 9 2 9 1 9 9 1 9 0 13 2
25 1 9 15 2 9 7 9 0 3 0 7 0 13 16 3 0 9 9 9 14 16 0 13 13 2
24 9 9 15 16 16 9 16 0 1 9 1 9 9 7 9 0 3 13 7 7 3 0 13 2
10 9 1 10 9 1 9 0 0 13 2
22 9 9 9 0 13 7 1 9 9 12 1 3 3 9 0 1 9 1 15 9 13 2
23 9 10 9 9 13 2 7 9 7 9 9 1 9 13 16 3 9 14 16 1 9 13 2
30 9 10 9 9 9 1 9 0 7 9 1 9 0 1 9 9 13 2 7 9 0 9 9 1 9 7 9 0 13 2
36 9 0 1 9 9 9 9 1 9 0 1 15 13 2 1 9 7 10 9 1 9 12 9 0 3 12 9 15 1 9 9 0 9 13 13 2
9 10 9 3 0 16 1 9 13 2
35 9 9 1 9 0 9 10 9 16 0 1 9 12 9 1 9 9 12 13 2 3 9 9 0 9 14 1 9 12 9 0 9 13 13 2
30 9 1 9 1 10 9 13 1 9 1 9 7 9 9 9 13 2 1 9 1 9 9 13 7 9 9 14 0 13 2
34 15 3 9 1 9 0 9 0 1 9 13 16 9 0 9 2 9 9 1 9 7 9 0 7 9 0 1 9 0 14 16 0 13 2
23 1 10 10 9 2 9 9 9 13 13 16 9 0 9 9 10 9 0 1 9 0 13 2
48 3 1 9 1 9 9 0 16 12 9 1 9 9 14 1 9 9 0 9 9 9 13 2 12 9 1 9 13 7 9 1 9 0 14 1 9 1 9 9 1 9 13 2 9 3 0 13 2
37 9 9 1 9 0 2 9 0 14 1 9 9 0 9 9 9 13 16 1 9 15 4 1 0 9 0 7 9 12 0 15 2 9 2 9 13 2
40 1 9 15 2 9 9 9 9 3 1 9 9 9 9 9 0 1 9 9 9 0 7 9 9 0 16 9 0 1 12 9 0 9 10 9 13 2 9 13 2
53 9 9 1 9 16 1 9 9 9 9 9 13 2 1 9 12 1 3 1 9 9 0 1 9 0 9 13 13 2 3 1 9 9 9 0 16 9 9 1 9 1 9 0 1 9 0 9 9 9 10 9 13 2
20 9 16 9 9 14 0 13 9 0 7 0 9 1 9 1 9 9 9 13 2
34 9 9 9 1 9 9 0 12 9 0 14 16 10 9 1 9 0 0 13 13 9 13 7 1 10 9 9 1 9 9 0 9 13 2
21 1 9 15 2 3 9 12 9 1 9 0 9 9 0 1 9 0 9 9 13 2
29 9 0 10 9 16 3 1 9 9 0 9 12 9 13 13 16 3 10 9 1 9 9 9 1 9 9 0 13 2
26 0 9 9 0 9 0 3 9 0 0 7 0 9 13 16 3 9 1 9 9 1 9 0 9 13 2
20 7 15 16 3 9 9 15 1 9 13 13 9 0 7 0 9 0 9 13 2
28 9 9 9 15 1 1 9 9 1 0 9 9 0 14 0 13 7 1 3 9 0 16 1 10 9 13 13 2
27 9 9 0 1 9 0 9 9 9 9 9 1 12 9 13 7 9 9 1 9 1 9 1 9 13 13 2
39 1 9 15 2 9 9 3 1 9 10 9 16 9 0 9 9 0 1 9 0 9 14 1 9 13 3 9 9 9 0 14 0 13 7 9 9 9 13 2
40 1 10 9 2 9 9 9 3 1 0 9 9 9 0 1 9 9 0 7 0 9 13 16 10 9 1 9 9 0 0 13 7 1 9 0 9 0 4 13 2
38 9 0 1 9 9 1 1 9 0 1 9 9 9 7 9 9 9 9 9 1 10 9 9 9 9 9 9 7 9 7 9 9 0 1 9 13 13 2
19 15 1 9 0 9 0 9 14 9 1 9 9 1 9 7 9 9 13 2
39 9 0 13 16 9 1 10 9 0 1 9 13 7 15 0 9 13 16 9 0 0 7 0 1 9 0 3 1 9 9 13 7 3 9 15 14 9 13 2
28 1 9 15 2 9 0 7 0 9 9 1 9 9 1 9 9 9 0 9 13 16 3 1 3 9 0 13 2
20 9 9 3 12 9 13 7 12 9 0 14 1 9 0 1 9 9 13 13 2
29 16 15 1 9 0 1 9 15 9 9 9 13 1 9 13 2 7 3 9 1 9 7 9 0 1 15 13 13 2
15 1 9 15 2 9 9 15 3 1 9 0 9 0 13 2
9 12 9 0 1 9 1 9 13 2
22 9 9 7 9 0 9 9 9 9 3 1 9 9 9 9 13 7 1 9 9 13 2
43 1 9 16 1 10 9 1 9 9 9 2 9 1 9 9 0 9 9 2 9 9 7 9 0 10 9 0 13 2 9 9 9 12 0 10 12 9 14 1 9 9 13 2
32 1 9 12 9 9 9 12 9 9 1 9 9 9 2 9 2 9 2 9 2 9 9 2 9 9 7 9 9 13 13 13 2
51 7 1 9 12 9 9 0 9 9 9 2 12 9 1 9 9 9 2 9 2 9 9 2 9 0 7 9 0 9 13 16 9 1 9 1 10 9 7 9 9 10 9 9 9 1 9 15 9 4 13 2
67 3 1 9 9 9 9 9 1 9 9 1 9 0 2 9 9 7 9 7 3 1 9 9 0 13 7 0 9 0 2 0 9 0 9 9 1 9 7 9 9 9 1 9 9 0 2 9 9 2 9 2 9 7 9 9 13 7 9 0 9 9 1 12 9 9 13 2
23 9 9 9 9 9 7 9 0 2 9 1 1 9 7 9 0 14 9 0 9 9 13 2
47 9 9 16 9 9 1 9 9 9 0 9 7 9 9 9 0 1 9 9 7 9 9 9 0 9 13 13 2 12 1 9 16 3 9 15 13 2 9 9 7 9 9 1 9 9 13 2
45 9 9 7 9 13 2 9 9 16 3 9 15 13 2 9 13 13 16 0 7 0 13 2 3 16 9 1 9 15 0 13 2 4 1 9 2 9 7 9 1 9 0 9 13 2
38 9 9 9 13 2 1 9 15 9 13 2 9 15 3 9 0 13 7 9 9 0 13 16 9 0 9 14 1 9 7 9 7 1 0 1 9 13 2
47 15 13 2 16 9 9 15 14 13 2 10 9 3 1 9 15 0 13 7 9 13 0 1 9 2 9 7 9 15 2 3 16 4 13 2 9 13 7 3 9 15 1 9 15 3 13 2
17 9 9 7 9 0 13 2 0 9 15 4 15 13 16 9 13 2
19 16 15 15 10 9 14 0 13 9 0 7 0 1 9 9 0 9 13 2
20 9 9 13 2 3 9 9 2 9 2 9 7 9 13 2 9 9 9 13 2
55 15 0 13 2 1 9 0 3 9 0 12 9 9 9 9 1 12 9 0 9 13 7 9 9 16 9 14 9 13 2 7 3 9 12 9 13 7 9 0 9 3 9 9 14 9 13 16 9 13 2 3 3 9 13 2
15 9 13 2 4 13 16 3 9 0 9 7 9 0 13 2
34 9 9 13 2 9 9 9 15 15 13 16 15 14 1 9 9 13 2 3 9 15 9 13 7 3 4 0 13 16 1 9 9 13 2
41 15 13 2 0 13 1 9 9 13 16 1 9 9 2 9 7 9 1 9 0 15 16 9 13 7 10 9 3 1 9 9 0 2 0 9 7 12 9 0 13 2
30 15 13 2 15 1 10 9 2 9 9 7 9 13 7 10 9 16 1 9 9 15 0 13 2 4 1 9 9 13 2
28 15 9 15 14 1 10 9 9 13 16 3 1 9 0 9 16 1 9 0 13 1 9 9 13 16 0 13 2
34 9 13 2 4 3 1 9 9 7 9 13 2 3 7 9 0 1 9 7 9 2 12 1 0 9 13 16 3 1 9 15 0 13 2
46 9 9 7 9 0 13 2 1 9 7 15 1 9 9 9 13 1 9 3 9 16 12 9 9 15 9 7 9 1 9 9 13 9 0 1 9 9 2 3 0 9 1 9 15 13 2
28 9 16 3 1 9 9 1 13 13 2 13 2 9 15 12 9 9 13 7 9 9 2 3 9 0 16 13 2
37 9 9 9 9 9 9 9 9 13 9 0 9 1 9 0 1 10 9 2 1 9 9 0 7 9 9 1 9 0 15 7 9 9 0 9 13 2
49 9 9 1 9 9 9 9 9 0 9 9 13 2 15 1 9 9 9 7 9 7 9 1 9 9 2 3 9 0 14 9 13 2 7 9 0 15 9 7 9 9 12 7 0 1 10 9 13 2
32 9 9 9 9 9 0 2 0 7 3 0 1 12 9 14 1 9 9 9 0 13 7 9 9 9 12 9 1 10 9 13 2
27 15 9 9 1 9 9 7 9 14 1 9 9 9 12 9 9 13 7 15 14 9 1 9 9 9 13 2
25 9 9 9 9 0 9 9 1 10 9 13 2 15 9 0 1 9 9 0 7 0 12 9 13 2
19 15 9 9 13 16 9 9 7 9 9 1 9 0 0 7 0 4 13 2
44 9 9 0 9 9 16 9 0 1 9 14 1 9 9 15 0 7 0 9 13 2 7 1 9 1 9 7 9 0 1 12 9 2 9 9 9 0 1 0 1 9 0 13 2
33 9 9 12 9 0 9 9 13 2 1 15 7 9 9 7 9 1 9 9 1 9 9 9 1 9 9 9 13 13 2 9 13 2
37 15 16 1 9 9 9 9 1 9 9 7 7 9 9 10 9 1 9 1 9 9 13 2 13 2 9 9 4 3 9 14 1 9 15 9 13 2
49 9 16 1 9 9 12 1 12 9 13 2 9 13 9 15 2 9 0 15 9 13 7 13 2 1 9 9 16 12 9 14 9 13 4 15 14 1 9 0 13 7 1 3 3 0 9 13 13 2
61 9 0 9 9 1 15 16 3 9 9 9 9 1 10 9 3 0 13 13 2 0 9 9 9 9 9 9 9 0 1 9 9 9 13 2 7 4 9 13 16 12 9 9 16 9 9 9 7 9 13 7 3 9 9 1 10 9 0 13 13 2
55 9 1 9 1 10 9 16 16 1 9 15 9 3 0 9 1 9 9 9 13 13 16 15 1 9 15 16 9 0 9 13 2 9 13 2 3 0 13 2 9 9 9 0 7 0 1 9 13 2 16 9 9 9 13 2
30 15 13 2 12 9 9 13 2 0 13 15 13 16 1 9 10 10 9 13 7 9 1 9 9 0 7 9 13 13 2
27 1 10 9 0 9 9 13 16 1 9 15 9 1 9 9 9 13 2 3 9 9 9 15 14 9 13 2
16 13 2 9 1 9 9 9 13 13 10 9 9 0 14 13 2
30 1 9 1 9 9 9 9 13 16 13 2 1 9 0 9 9 9 9 13 7 9 13 9 1 9 9 1 9 13 2
27 9 16 9 9 1 9 9 13 13 2 9 9 9 3 0 13 7 9 9 1 9 0 9 9 9 13 2
31 9 0 9 0 9 13 2 9 9 0 1 12 12 9 9 0 0 0 9 13 16 10 9 1 1 9 12 2 9 13 2
62 9 9 9 3 1 9 0 9 9 0 7 0 1 9 1 9 13 2 9 0 0 9 1 9 0 9 13 16 9 0 1 9 1 9 9 0 9 2 9 0 0 2 0 7 9 0 2 9 2 1 9 9 13 16 1 0 1 9 0 9 13 2
52 15 1 1 9 0 9 0 1 1 9 9 1 9 1 9 0 9 13 2 1 9 10 9 2 9 1 9 0 7 9 0 9 0 9 0 9 1 9 13 7 9 0 13 10 9 14 1 9 0 9 13 2
25 15 13 2 9 10 9 1 9 0 3 1 9 7 9 16 9 0 13 2 1 9 0 9 13 2
20 7 16 0 13 2 9 13 9 9 15 1 9 0 16 1 9 0 13 13 2
31 9 0 9 9 3 1 9 9 9 9 13 2 9 12 9 9 0 9 9 15 14 1 1 9 9 9 9 0 13 13 2
47 1 9 9 10 9 9 9 0 10 9 1 9 9 9 9 9 2 9 12 0 1 9 9 1 9 9 1 9 9 1 9 9 9 7 9 9 1 9 12 9 9 1 9 9 0 13 2
39 9 9 0 9 9 9 0 1 9 9 9 12 0 1 9 9 1 9 9 1 9 9 1 9 9 2 9 7 9 1 12 9 9 1 9 9 0 13 2
34 9 9 0 9 9 9 9 2 12 0 2 0 1 9 9 1 9 9 1 9 9 1 9 9 1 12 9 9 1 9 9 0 13 2
25 9 9 0 9 9 9 9 2 0 12 0 2 1 9 9 7 9 9 1 12 9 9 0 13 2
29 9 9 0 9 9 9 9 2 9 0 2 12 0 2 1 9 9 7 9 1 9 9 1 12 9 9 0 13 2
41 1 1 9 9 2 9 9 9 9 9 9 9 0 1 0 1 9 1 15 16 9 15 1 9 7 9 1 15 9 9 13 9 0 9 9 1 9 9 13 13 2
34 9 9 9 16 9 13 2 12 9 0 9 1 9 9 9 2 9 9 7 9 9 1 9 1 9 9 7 9 9 0 2 9 13 2
8 9 0 9 3 1 9 13 2
40 9 9 2 9 9 9 9 9 0 10 9 1 9 0 9 14 16 3 0 9 13 2 1 9 3 0 9 9 12 9 1 9 0 7 0 2 3 9 13 2
41 9 9 9 9 9 9 0 9 1 9 1 9 9 12 9 1 9 0 0 7 0 13 2 9 9 9 9 9 0 9 1 9 12 9 14 1 15 0 4 13 2
37 15 13 2 9 9 1 9 1 9 1 0 9 9 9 0 12 9 16 1 9 12 9 7 0 9 15 1 9 12 1 9 0 13 2 9 13 2
38 9 13 2 9 14 16 9 1 9 0 9 0 13 1 10 9 4 9 13 16 9 9 0 9 1 12 9 0 12 9 1 9 0 15 9 13 13 2
50 15 1 9 0 9 7 9 13 2 12 9 1 9 0 1 9 9 0 1 9 7 9 0 9 0 13 7 9 9 1 9 9 9 9 9 1 9 9 9 9 7 9 9 12 9 9 0 4 13 2
47 9 9 9 0 9 13 2 1 1 9 0 9 9 7 9 2 12 9 12 9 0 0 16 9 0 2 9 0 2 9 0 7 9 0 1 9 1 9 9 14 9 13 2 16 9 13 2
37 15 9 9 9 7 9 14 1 9 9 9 13 7 13 2 1 9 12 9 9 1 9 1 12 12 9 7 9 1 9 1 12 12 9 0 13 2
28 15 13 2 9 9 0 9 1 9 1 9 12 0 12 12 9 7 9 0 1 9 12 12 9 9 13 13 2
28 9 13 2 9 0 2 0 2 9 0 2 9 2 9 2 9 0 7 9 2 9 0 0 9 1 9 13 2
10 9 0 13 1 9 9 9 9 13 2
28 1 10 9 9 2 9 7 9 0 1 10 9 0 9 9 13 7 9 9 0 9 1 9 0 9 0 13 2
27 7 1 9 2 12 9 0 1 9 7 9 9 13 1 9 12 7 7 12 9 9 1 9 13 13 2 2
77 9 9 1 9 1 9 12 9 9 0 9 9 0 9 1 9 9 0 9 1 9 14 0 13 7 3 13 13 2 9 0 9 0 9 1 9 15 13 16 9 14 1 9 9 7 9 9 9 13 7 1 15 9 13 2 15 14 0 9 0 13 7 13 16 15 13 9 15 14 13 7 9 15 14 9 13 2
23 3 3 9 9 0 0 13 2 16 1 10 9 16 9 0 0 1 12 9 1 3 13 2
64 4 9 13 16 10 9 0 4 3 9 0 0 14 1 9 1 9 7 9 9 9 7 7 0 1 9 0 9 9 13 16 1 9 9 0 7 1 9 9 0 0 9 13 7 15 1 9 15 13 16 9 0 15 15 9 13 16 15 7 9 14 9 13 2
47 0 1 9 9 0 9 0 1 10 9 13 16 16 9 7 9 1 15 1 9 0 1 9 1 9 9 0 13 7 9 15 15 1 9 9 0 9 13 1 10 9 9 0 9 0 13 2
62 4 9 13 9 16 1 9 9 13 2 0 9 9 1 9 0 9 13 2 16 3 9 1 0 9 9 0 13 2 0 3 9 13 16 1 9 4 9 15 13 7 1 9 9 0 0 13 16 9 1 9 13 7 9 14 1 9 15 15 0 13 2
66 4 1 10 9 16 9 13 16 9 9 13 7 9 1 1 9 1 9 13 7 10 9 1 12 3 0 7 0 9 13 2 7 9 9 9 7 9 9 1 9 9 15 13 16 9 0 1 9 0 9 9 13 13 7 4 9 0 14 1 9 1 9 0 9 13 2
67 0 13 16 1 10 9 9 9 9 9 7 7 9 9 9 16 9 0 14 1 9 9 13 9 9 9 13 7 12 9 0 1 9 9 0 1 9 0 9 13 0 1 15 7 1 9 0 7 9 0 1 9 0 1 15 13 7 4 9 9 14 1 9 9 0 13 2
55 9 9 0 1 9 15 2 1 9 9 13 2 13 13 2 9 9 0 7 9 1 9 0 7 1 9 9 0 9 2 9 9 0 1 9 14 1 9 9 7 9 9 0 1 1 9 9 14 0 1 9 9 13 13 2
54 16 10 9 7 9 16 3 9 1 9 9 15 0 13 2 9 13 3 7 3 1 10 9 9 0 13 7 1 1 9 9 0 13 16 9 0 9 13 2 7 1 10 9 15 9 13 16 1 9 0 9 0 13 2
33 1 9 0 10 9 7 9 16 2 9 0 1 9 9 0 1 9 0 1 9 0 1 9 9 9 9 7 9 2 9 4 13 2
37 15 1 9 13 16 15 1 10 9 7 9 1 1 9 3 0 2 7 9 9 15 2 3 9 0 13 7 3 9 7 9 14 16 1 9 13 2
40 3 3 16 0 13 13 7 3 9 10 9 9 7 9 1 9 0 0 16 1 9 9 15 1 9 7 9 2 9 13 2 0 1 9 3 13 1 9 0 2
56 3 7 10 9 7 9 1 12 9 0 0 13 7 3 0 13 16 16 9 9 0 15 9 14 1 9 0 13 2 3 9 1 9 9 0 9 13 2 7 15 0 9 13 16 0 13 9 7 9 9 0 1 15 9 13 2
22 9 0 4 13 16 16 15 1 10 9 3 9 13 7 10 9 1 9 0 9 13 2
25 16 10 9 2 1 9 0 0 13 7 16 9 0 9 13 2 3 1 10 9 2 9 0 13 2
29 3 7 1 10 9 2 9 10 9 0 7 0 14 1 9 0 15 9 13 7 1 9 15 2 15 9 4 13 2
120 1 9 7 9 1 9 0 7 0 1 9 9 9 7 9 2 9 13 16 3 10 9 7 9 0 7 0 1 1 9 9 2 3 1 15 1 9 0 7 0 1 9 15 1 9 9 0 9 9 13 2 9 13 7 15 9 9 15 16 13 2 7 9 0 1 10 9 15 13 16 10 9 9 7 9 7 10 9 1 9 9 2 0 9 0 7 0 0 16 13 7 1 3 1 9 0 9 13 16 9 9 7 9 1 9 9 1 9 9 2 1 9 9 0 9 13 7 9 13 2
36 10 9 0 13 16 3 9 1 9 9 1 9 9 13 7 3 0 2 9 13 13 7 9 0 0 1 10 9 7 9 2 1 9 13 13 2
59 3 1 9 9 4 13 16 16 10 9 9 1 9 9 7 9 9 9 0 1 10 9 12 9 0 1 9 1 9 7 9 9 1 9 0 13 13 7 15 7 15 1 9 10 9 2 1 9 0 7 0 1 1 10 9 9 9 13 2
15 9 1 9 0 1 10 9 1 9 3 9 2 9 13 2
30 16 1 9 13 16 0 1 9 7 9 16 1 9 9 9 13 2 0 1 9 9 7 9 13 16 1 10 9 13 2
15 1 9 9 2 9 0 7 3 0 1 10 9 4 13 2
12 4 9 13 16 6 9 0 7 0 9 13 2
17 9 1 9 9 14 1 9 10 9 1 9 0 2 0 4 13 2
25 12 2 9 0 13 2 16 3 1 9 9 9 9 0 7 9 9 12 9 9 7 9 0 13 2
8 1 9 2 4 9 0 13 2
14 12 2 9 0 13 2 15 14 1 9 9 4 13 2
53 9 9 16 3 1 9 0 9 2 12 2 12 9 9 9 14 1 9 9 1 15 9 13 7 9 12 9 0 0 13 2 3 1 9 9 9 3 1 0 9 0 9 9 7 1 12 2 12 9 9 0 13 2
21 1 9 0 4 1 9 0 2 9 0 13 7 9 13 16 6 2 9 0 13 2
2 3 2
21 3 1 10 9 16 1 9 0 7 0 16 4 9 0 3 0 9 14 9 13 2
70 9 9 0 13 1 9 16 9 0 1 9 9 0 13 7 9 0 16 3 1 9 9 12 9 0 9 13 13 2 9 13 9 14 1 9 15 9 2 9 2 9 2 9 7 9 2 13 7 1 9 16 3 16 13 9 13 2 9 13 2 16 9 16 13 15 1 9 9 13 2
19 1 10 9 3 9 9 9 16 3 0 9 0 1 9 13 3 9 13 2
18 1 9 13 16 12 9 1 9 9 9 7 9 7 9 0 9 13 2
29 9 0 1 1 9 9 0 7 9 9 1 9 9 9 7 9 7 9 9 0 1 9 9 7 9 7 9 13 2
29 1 10 9 2 9 9 9 2 9 2 9 9 7 2 9 13 7 9 9 9 2 9 2 9 7 9 9 13 2
20 1 9 0 9 0 2 9 13 16 1 1 9 9 0 0 7 9 0 13 2
20 10 9 9 1 9 9 9 7 1 9 9 9 9 2 1 9 2 0 13 2
15 7 3 1 9 13 1 9 0 2 9 7 9 13 13 2
15 9 7 9 9 9 2 1 9 0 0 9 0 13 13 2
14 9 9 9 14 4 9 9 1 9 9 9 0 13 2
39 9 9 1 10 9 16 9 7 9 10 9 9 0 9 0 1 9 7 9 0 1 9 0 13 7 15 14 1 1 9 9 7 9 9 0 3 0 13 2
16 10 9 0 16 1 9 9 0 13 13 2 9 10 9 13 2
41 16 9 9 9 1 9 9 9 0 14 1 9 9 13 7 9 7 9 15 14 9 1 9 9 9 9 0 9 13 2 9 9 3 9 0 1 9 0 4 13 2
19 9 7 9 16 1 9 9 9 13 2 3 9 0 14 1 9 4 13 2
51 9 9 1 9 1 9 9 9 9 7 9 7 9 1 9 16 1 9 9 0 7 9 0 9 13 13 2 0 13 9 0 15 14 1 9 9 13 7 9 9 13 16 1 9 9 0 0 9 0 13 2
30 9 9 1 9 15 9 9 0 9 14 1 9 0 7 0 9 16 3 9 13 1 0 9 13 7 3 13 13 2 2
42 9 9 0 9 7 9 1 9 9 7 9 9 9 7 9 9 1 10 12 9 9 1 15 13 16 15 1 9 0 9 7 9 0 9 3 1 9 0 15 9 13 2
41 9 9 9 1 10 9 9 13 13 16 9 9 9 1 9 9 9 0 2 9 0 13 7 9 9 10 9 1 10 9 2 9 9 0 9 9 7 9 9 13 2
29 16 16 3 9 9 9 2 9 2 3 9 1 9 9 3 9 9 9 14 13 2 7 9 0 16 0 13 13 2
19 1 1 9 9 9 2 9 9 9 9 9 0 0 14 1 9 13 13 2
64 9 0 9 16 9 9 1 15 9 13 15 13 16 16 9 0 15 1 9 9 9 9 2 7 1 3 9 9 9 0 1 9 1 12 12 9 7 0 15 15 14 1 9 1 9 15 13 13 2 16 4 10 9 9 0 14 3 1 9 1 10 9 13 2
51 16 1 9 9 9 0 2 9 9 14 1 9 0 7 1 9 9 0 1 9 12 9 13 2 3 16 0 13 2 9 0 1 9 0 9 15 9 13 2 3 9 13 16 3 1 10 9 0 9 13 2
22 16 1 9 1 9 0 9 2 3 4 1 9 9 1 9 9 7 9 0 9 13 2
44 1 9 3 2 9 9 0 7 9 9 7 9 16 9 14 0 13 16 0 0 9 7 9 1 9 9 9 0 9 13 7 3 0 1 9 9 9 0 1 9 7 9 0 2
37 1 9 9 9 3 1 13 16 9 0 15 7 9 15 1 9 9 9 13 7 0 9 9 0 0 1 9 9 13 16 1 9 15 9 13 13 2
29 15 3 1 15 7 9 0 13 16 1 9 9 9 0 1 9 9 7 9 0 9 0 3 4 9 14 9 13 2
38 12 9 0 1 9 1 0 9 9 9 9 1 1 1 9 1 12 12 9 0 2 13 2 9 0 9 3 1 9 9 15 1 9 0 15 9 13 2
60 9 9 9 0 1 9 16 1 9 0 9 9 1 9 9 1 9 0 9 13 2 13 2 0 1 9 0 2 3 1 0 9 16 1 9 15 3 13 2 1 9 9 2 1 0 1 9 2 1 9 9 15 2 1 9 0 15 1 13 2
30 9 13 2 0 1 10 9 2 1 9 9 0 1 9 0 7 9 0 15 2 1 9 0 15 1 9 2 9 13 2
14 7 10 0 9 1 10 12 9 9 15 2 9 13 2
17 9 0 9 12 9 0 7 0 14 9 13 7 15 13 9 15 2
37 9 9 1 9 16 1 9 0 0 16 1 9 7 9 0 13 7 1 9 9 0 7 0 1 9 15 1 13 1 9 10 9 9 13 13 13 2
33 9 9 3 1 12 9 9 1 9 2 1 9 3 0 15 1 9 12 9 9 1 9 2 9 13 16 1 9 2 1 9 13 2
32 9 1 12 9 0 0 2 2 12 9 0 2 14 0 13 16 3 0 9 0 1 12 9 13 16 1 9 1 9 9 13 2
16 15 13 2 0 1 9 0 9 2 9 0 1 9 3 13 2
17 15 9 13 16 16 1 9 13 2 1 10 9 1 9 9 13 2
22 1 9 7 15 0 13 7 15 4 9 13 9 15 14 1 10 9 9 2 0 13 2
33 9 13 2 1 9 15 1 9 1 9 9 13 2 7 3 9 0 0 13 2 15 4 1 9 2 1 9 0 7 0 9 13 2
9 1 9 15 9 0 1 9 13 2
8 15 0 12 9 3 0 13 2
29 9 9 15 1 1 15 0 13 2 7 9 0 0 0 9 13 16 16 1 15 9 13 13 2 3 1 4 13 2
18 9 0 13 16 1 9 2 3 3 4 1 12 9 9 0 9 13 2
20 7 1 9 15 1 9 15 9 13 2 9 16 1 10 9 9 2 0 13 2
11 9 9 16 1 9 15 2 9 0 13 2
20 15 13 2 9 1 9 9 1 9 0 13 7 3 9 1 9 2 0 13 2
8 1 9 0 9 10 9 13 2
6 7 9 1 15 13 2
7 15 0 1 9 9 13 2
11 1 9 15 9 9 7 9 9 9 13 2
40 9 9 9 9 1 9 9 15 1 9 0 1 9 9 9 2 9 12 9 0 9 13 16 12 9 3 9 0 15 1 9 14 3 13 16 1 9 15 13 2
20 15 3 1 9 9 15 1 9 13 13 9 1 9 1 9 9 15 0 13 2
18 9 1 9 1 9 9 9 13 7 13 16 1 3 1 9 4 13 2
10 15 1 9 0 1 9 2 0 13 2
16 1 9 9 2 9 1 9 0 2 16 0 13 7 7 0 2
17 15 16 12 1 9 12 9 0 13 16 1 9 9 9 13 13 2
22 15 16 3 1 9 9 9 0 13 13 7 1 15 2 9 15 1 9 7 9 13 2
15 7 9 9 15 13 2 15 1 9 9 0 1 9 13 2
5 3 15 14 13 2
13 15 1 9 9 1 9 2 1 9 0 9 13 2
16 9 9 9 9 13 7 9 0 1 9 9 7 9 0 13 2
8 7 9 14 13 3 9 13 2
49 9 13 2 9 1 0 1 9 9 0 7 0 13 16 16 15 9 14 9 13 7 1 9 13 2 1 9 9 9 9 1 9 2 9 3 0 9 13 7 10 9 1 9 15 1 9 9 13 2
21 9 9 3 1 12 9 9 1 9 2 3 12 9 13 16 1 9 1 13 13 2
14 15 1 9 9 1 9 2 1 9 9 12 9 13 2
15 15 12 9 1 9 12 9 0 1 9 9 0 9 13 2
26 7 1 9 9 1 9 13 2 15 3 1 9 15 9 9 13 7 3 16 4 10 9 14 0 13 2
25 9 9 2 1 9 9 9 7 9 9 13 13 2 1 9 9 2 9 0 13 7 9 9 13 2
50 9 1 15 13 16 9 13 7 3 1 9 7 9 2 7 1 3 10 9 9 9 1 9 13 7 16 9 15 3 0 13 16 15 13 1 9 0 13 3 1 9 7 9 2 9 7 9 0 13 2
16 9 7 9 7 9 7 9 0 1 15 0 9 9 9 13 2
21 9 9 9 2 9 2 3 9 9 7 9 9 1 10 9 0 7 9 0 13 2
36 9 9 2 9 2 3 13 13 16 0 9 1 9 13 2 7 10 9 7 9 9 15 13 16 9 1 9 14 0 0 9 7 9 9 13 2
25 16 1 9 9 2 9 2 9 13 16 0 9 15 13 2 9 15 1 9 10 9 1 9 13 2
27 9 9 9 2 9 2 12 9 0 13 2 12 2 3 1 9 9 9 16 9 0 1 9 13 9 13 2
21 12 2 9 14 1 9 12 9 16 9 0 7 0 14 1 9 13 13 9 13 2
19 12 2 9 9 1 9 7 9 1 10 9 16 9 9 14 0 13 13 2
5 9 0 15 13 2
23 9 1 9 9 2 9 2 13 1 9 9 7 9 9 2 9 2 13 2 7 9 13 2
30 9 9 2 9 2 1 9 13 2 9 15 16 9 14 0 13 0 9 1 9 13 7 3 3 15 1 10 9 13 2
14 9 7 9 16 9 0 1 9 13 2 0 7 0 2
12 9 13 2 15 16 13 1 15 9 4 13 2
12 1 9 9 6 9 15 3 1 15 9 13 2
15 9 14 1 9 9 9 13 15 16 1 9 15 9 13 2
29 1 9 9 16 15 14 1 9 13 1 9 9 4 13 7 9 2 9 2 16 9 9 1 15 13 9 15 13 2
37 9 13 2 15 16 13 15 14 1 9 1 9 0 4 13 2 16 15 14 1 9 0 13 2 15 16 15 7 9 15 14 1 9 9 0 13 2
17 7 15 14 1 0 1 9 0 13 1 15 7 1 9 9 13 2
10 9 16 1 9 9 9 13 7 13 2
14 15 0 13 7 9 13 2 15 15 14 0 0 13 2
13 16 0 13 7 9 13 9 15 14 9 4 13 2
11 9 9 1 9 13 16 1 9 0 13 2
5 15 4 9 13 2
4 15 9 13 2
22 9 1 9 13 2 9 1 10 0 9 2 9 8 9 2 9 2 7 2 9 13 2
11 16 15 9 13 2 15 9 9 4 13 2
9 9 13 16 3 1 9 4 13 2
14 9 1 9 9 13 13 2 15 14 1 9 13 13 2
11 9 7 9 7 9 7 9 0 9 13 2
21 13 2 3 15 0 9 15 9 13 7 9 9 14 1 9 9 9 15 9 13 2
18 1 9 8 9 2 9 2 7 9 7 9 7 9 7 9 9 13 2
6 9 14 3 9 13 2
20 1 10 9 13 2 15 9 0 9 13 1 15 12 9 1 9 16 9 13 2
18 1 9 9 2 9 2 13 13 9 10 12 9 0 1 9 15 13 2
11 10 9 14 1 12 9 0 16 13 13 2
29 16 9 3 9 14 9 7 9 13 13 16 10 12 9 9 13 1 9 9 13 7 9 3 1 15 9 13 13 2
10 9 9 8 9 2 9 2 0 13 2
12 7 0 13 10 9 3 9 1 15 4 13 2
13 1 9 9 2 9 2 9 2 2 9 9 13 2
13 1 9 9 13 13 2 0 9 9 7 9 13 2
20 9 9 2 9 2 7 9 9 0 9 2 9 7 2 16 1 9 0 13 2
9 9 14 16 1 9 9 13 13 2
16 9 9 13 1 9 0 7 9 9 7 9 9 9 9 9 2
14 3 13 2 6 9 9 2 1 9 1 9 0 13 2
25 3 9 7 9 2 9 7 9 14 0 13 3 15 7 9 14 9 13 7 15 1 9 9 13 2
8 9 14 1 0 9 9 13 2
5 9 9 0 13 2
5 0 9 9 13 2
17 9 16 1 9 1 9 9 13 2 0 9 1 9 1 9 13 2
17 1 9 9 16 1 9 9 9 0 1 9 13 1 15 9 13 2
30 9 9 2 9 2 1 13 7 13 2 1 9 9 9 16 1 9 9 7 9 7 9 0 1 9 13 14 9 13 2
13 9 13 2 16 9 15 1 10 9 15 15 13 2
8 9 2 9 2 13 2 6 2
8 9 13 2 1 15 9 13 2
11 15 16 13 9 15 1 9 15 0 13 2
7 9 15 9 9 9 13 2
9 9 15 7 9 15 0 9 13 2
17 7 1 9 15 2 9 15 7 9 15 9 14 1 9 0 13 2
9 9 1 9 15 9 14 9 13 2
19 2 9 1 9 2 9 9 2 9 2 13 2 9 15 1 15 0 13 2
15 15 9 0 14 1 9 13 2 9 14 1 9 9 13 2
14 9 13 2 1 9 2 16 13 15 1 15 0 13 2
12 1 9 9 9 0 9 9 2 9 2 13 2
14 9 2 9 2 13 2 10 9 0 7 9 0 13 2
12 9 0 7 9 9 7 9 1 15 0 13 2
26 9 13 2 0 13 1 9 15 9 13 2 16 10 9 14 1 9 15 16 13 15 15 14 9 13 2
27 9 9 1 9 13 7 13 2 9 2 9 2 9 2 13 7 3 1 15 9 14 1 9 9 0 13 2
8 9 9 14 1 9 9 13 2
15 16 3 9 9 13 2 15 9 14 1 9 9 15 13 2
17 9 16 1 3 9 2 9 0 14 9 13 16 9 14 9 13 2
14 9 9 14 9 13 16 9 2 9 2 9 13 13 2
13 9 16 1 9 9 13 16 9 3 9 13 13 2
9 10 9 1 9 9 15 9 13 2
22 15 16 1 9 15 13 16 1 9 1 9 1 9 9 7 9 9 1 9 9 13 2
11 9 1 13 7 9 9 0 14 9 13 2
19 13 2 9 2 9 14 1 9 9 0 13 16 0 9 14 1 9 13 2
10 9 16 12 9 14 1 9 9 13 2
12 1 9 7 9 15 9 16 1 9 9 13 2
7 9 3 1 9 9 13 2
9 1 9 3 13 7 1 9 13 2
24 10 9 13 13 1 9 7 1 9 9 0 7 0 13 2 1 9 0 1 9 7 9 13 2
13 9 13 9 14 16 9 13 13 1 9 15 13 2
27 9 8 9 2 9 2 7 2 9 13 2 15 3 1 9 9 13 7 13 16 10 0 9 16 9 13 2
32 16 12 9 1 15 9 0 13 16 13 9 13 2 15 14 9 7 9 13 2 9 15 13 13 7 9 15 1 9 1 13 2
17 9 1 9 9 9 13 2 6 9 9 10 0 9 16 9 13 2
25 9 1 9 9 13 2 6 9 9 2 16 1 1 15 9 13 2 9 13 16 9 15 14 13 2
5 9 13 2 6 2
11 3 9 9 9 1 15 9 9 0 13 2
20 9 9 2 9 9 0 9 14 3 9 13 13 2 9 1 9 9 13 13 2
10 1 9 9 1 9 0 9 13 13 2
5 9 13 2 9 2
26 15 1 9 15 7 9 15 2 9 14 1 9 9 9 13 2 8 8 8 2 1 9 9 9 13 2
30 1 9 9 8 9 2 9 2 7 9 2 9 9 13 13 2 15 9 13 1 9 0 9 9 2 9 14 9 13 2
37 10 9 2 12 1 0 7 0 9 9 7 9 9 13 7 9 10 9 16 9 9 7 9 9 1 12 9 1 9 0 7 9 7 9 0 13 2
17 10 9 2 1 12 9 2 9 0 7 0 7 0 9 9 13 2
15 1 1 15 15 10 9 7 9 14 16 3 9 9 13 2
22 9 9 9 9 13 2 9 9 14 3 9 13 13 16 9 9 14 9 1 9 13 2
46 12 1 9 9 1 15 16 3 9 13 9 13 1 3 0 13 16 10 9 16 1 9 9 3 12 9 1 9 9 9 13 2 3 1 9 1 9 1 9 2 9 14 1 9 13 2
25 1 9 0 9 9 2 9 9 9 13 7 9 9 1 9 12 9 3 13 1 9 9 9 13 2
43 9 9 9 3 1 9 1 9 7 9 1 9 9 1 9 1 9 2 1 9 13 13 16 15 9 9 9 14 1 9 9 9 9 13 7 1 10 9 1 9 9 13 2
23 1 9 9 0 9 7 9 0 2 12 9 12 0 1 9 9 9 9 1 9 13 13 2
23 9 9 0 9 9 13 2 10 9 12 1 0 9 0 1 9 9 1 9 0 9 13 2
26 9 9 13 2 10 9 0 1 9 13 16 1 3 9 12 1 12 9 9 13 7 12 9 9 13 2
28 15 13 2 9 9 0 9 0 0 7 0 1 9 7 9 9 0 13 16 9 9 0 15 1 9 9 13 2
29 15 13 2 12 9 9 2 9 2 9 2 9 2 9 2 9 7 9 16 1 9 10 9 1 9 9 13 13 2
25 9 9 13 2 9 10 9 1 9 9 9 9 9 7 9 9 9 1 9 9 1 10 9 13 2
27 1 9 9 9 9 0 1 9 9 9 9 0 9 1 9 9 0 9 9 9 1 9 9 1 9 13 2
37 1 10 9 0 16 9 9 9 9 13 7 1 9 9 9 0 9 7 9 9 13 13 2 12 9 0 0 1 9 9 9 1 9 9 9 13 2
52 9 0 9 2 9 9 1 9 0 7 9 0 15 2 9 9 1 9 9 7 9 2 9 0 1 9 9 2 9 9 0 0 7 9 0 15 2 1 9 9 9 13 16 1 10 9 1 9 0 9 13 2
29 0 1 9 10 9 2 9 9 0 7 9 7 9 9 9 10 9 1 9 9 9 0 1 9 1 9 9 13 2
21 0 1 9 9 0 9 9 9 9 9 9 9 9 9 1 9 1 9 9 13 2
22 9 9 2 9 7 9 1 10 9 13 2 10 9 1 9 9 0 9 9 13 13 2
21 9 9 9 13 2 9 9 0 9 9 2 9 7 9 0 7 0 7 9 13 2
17 1 10 9 1 9 9 9 9 9 9 16 1 9 9 9 13 2
19 1 9 10 9 1 12 9 9 2 12 12 9 9 1 9 13 13 13 2
19 9 9 0 9 9 13 2 3 12 12 9 1 9 9 10 9 9 13 2
33 9 9 13 2 1 10 9 9 12 12 7 12 12 9 1 9 9 9 7 9 7 9 1 9 9 0 7 9 9 13 13 13 2
22 15 13 2 10 9 9 9 12 9 0 9 0 1 9 9 9 1 12 9 0 13 2
21 9 9 0 0 9 1 9 9 9 1 9 9 1 9 9 7 9 0 9 13 2
29 10 9 16 0 12 12 7 12 9 9 13 1 9 1 9 12 12 7 12 9 2 9 9 9 9 9 13 13 2
40 1 10 9 1 12 9 2 9 9 9 9 2 9 9 2 9 9 2 9 0 2 9 9 7 0 2 9 9 7 9 9 7 9 9 1 9 9 13 13 2
29 1 1 9 9 9 0 7 0 9 9 2 3 12 7 12 9 9 1 9 0 13 1 10 9 9 0 14 13 2
16 9 9 9 9 10 9 14 12 12 7 12 12 9 9 13 2
43 9 13 2 1 9 0 0 1 12 12 7 12 9 9 1 9 0 1 9 9 9 0 7 0 9 9 0 14 13 16 10 9 1 1 9 12 9 0 1 9 13 13 2
20 9 9 7 9 9 9 0 3 10 9 14 12 12 7 12 12 9 9 13 2
17 9 9 9 13 2 10 9 1 9 9 1 10 9 9 4 13 2
26 15 13 2 9 9 9 1 9 7 9 1 9 0 7 0 10 9 1 9 9 9 3 0 4 13 2
37 9 13 1 9 10 9 1 9 10 9 9 0 2 12 2 12 9 1 9 0 7 7 0 9 13 16 9 10 9 1 0 9 9 12 9 13 2
35 1 1 9 15 2 9 0 1 9 9 9 1 9 0 16 12 1 12 13 16 9 9 9 7 9 9 12 9 1 0 9 0 9 13 2
15 9 9 9 1 9 0 1 9 9 9 7 9 9 13 2
26 1 9 9 0 12 12 9 9 9 1 9 9 13 16 1 10 9 12 12 9 0 7 9 0 13 2
31 1 9 1 9 0 1 9 9 0 1 9 9 9 9 1 10 9 0 1 9 13 7 1 9 9 9 1 9 9 13 2
34 9 9 9 1 9 9 2 9 2 9 2 9 2 9 2 9 7 9 1 9 0 10 9 2 1 12 9 9 1 9 0 9 13 2
21 9 9 1 9 9 9 9 1 9 0 10 9 2 1 12 9 9 9 4 13 2
20 9 9 9 13 2 3 9 0 10 9 1 12 9 9 1 12 12 9 13 2
34 9 9 13 2 1 9 0 9 12 9 0 1 9 9 2 9 0 7 0 9 2 9 9 1 12 9 9 7 12 9 9 9 13 2
18 1 9 15 3 1 9 12 9 0 1 10 9 12 12 9 9 13 2
36 15 13 2 9 3 9 12 9 7 9 2 9 9 2 9 2 9 2 9 2 9 0 2 9 9 1 9 0 1 10 9 1 9 9 13 2
22 0 9 9 0 9 9 7 9 9 2 1 9 9 9 9 7 9 9 9 0 13 2
44 9 1 9 10 9 0 9 9 9 9 7 9 9 1 9 0 9 0 2 9 9 0 1 9 9 9 7 9 9 7 9 9 1 9 7 9 15 1 9 0 9 9 13 2
26 9 9 7 9 9 9 9 9 9 13 2 3 12 12 9 1 9 9 10 9 1 9 9 13 13 2
30 9 9 13 2 9 9 1 9 1 9 9 9 0 1 9 9 9 7 9 9 0 1 1 9 0 1 9 9 13 2
49 15 9 13 2 1 0 9 1 9 12 9 9 0 0 1 9 9 9 7 9 9 0 7 1 1 15 9 12 9 9 0 0 1 9 9 2 9 7 9 1 9 0 1 1 9 9 13 13 2
34 9 9 7 9 9 9 9 9 13 2 9 0 9 1 9 9 9 9 9 12 9 0 2 0 1 9 7 0 1 9 0 9 13 2
21 9 9 9 9 13 2 0 1 12 12 9 9 9 7 9 1 9 9 9 13 2
26 9 9 13 2 10 9 9 1 12 12 7 12 9 9 9 9 1 9 9 0 1 9 1 9 13 2
27 9 9 1 9 9 9 1 9 9 7 9 9 1 9 9 2 9 7 9 2 1 9 0 9 9 13 2
25 15 9 13 2 12 12 7 12 9 1 9 9 1 9 9 7 12 9 1 9 9 9 13 13 2
27 9 13 2 10 9 9 1 9 12 9 7 9 1 9 12 12 7 12 9 1 9 9 1 9 9 13 2
27 15 13 2 1 3 0 1 12 12 9 9 0 9 1 9 1 9 9 9 13 7 9 9 9 9 13 2
34 1 9 9 9 1 9 9 0 1 9 9 9 9 0 2 9 9 0 10 9 1 9 0 1 12 9 1 12 2 12 9 9 13 2
24 9 9 9 1 9 9 0 9 9 13 2 1 10 9 9 9 9 1 9 10 9 9 13 2
25 15 9 9 9 0 0 9 1 9 9 9 14 9 1 9 9 0 0 7 9 9 0 9 13 2
25 9 0 9 0 9 1 9 0 0 1 9 0 13 16 9 9 9 14 1 10 9 9 13 13 2
40 9 1 9 0 7 0 0 1 9 9 16 1 12 9 3 9 13 2 0 1 9 0 9 7 9 9 0 1 0 9 1 9 9 1 9 9 9 9 13 2
66 1 9 9 0 9 9 0 9 2 10 9 16 0 9 9 0 2 0 2 9 0 2 9 9 2 9 2 9 2 9 2 9 0 2 9 0 2 9 0 7 9 0 7 2 13 2 12 9 3 1 9 9 1 9 13 16 0 1 9 7 9 0 10 9 13 2
31 10 9 16 1 12 0 9 9 9 7 1 9 9 0 3 13 2 1 9 9 12 1 9 9 9 9 1 9 9 13 2
38 9 1 9 3 1 9 1 9 9 9 1 10 9 9 13 13 16 15 1 1 9 15 9 14 16 1 9 1 9 1 9 9 13 1 9 9 13 2
34 9 9 0 1 9 9 0 9 9 1 9 13 16 1 9 9 0 0 1 9 0 16 9 15 3 1 9 0 1 13 13 13 13 2
24 9 9 9 1 9 0 7 0 13 16 3 1 9 12 1 12 3 1 9 1 10 9 13 2
29 10 9 3 1 9 0 9 9 9 9 1 15 14 9 13 7 1 9 9 9 1 9 0 3 1 9 9 13 2
11 9 9 9 2 9 9 9 9 9 13 2
6 9 2 9 0 9 2
23 9 9 9 9 0 9 9 9 9 2 9 9 9 1 9 12 0 9 0 14 9 13 2
34 9 9 9 9 9 0 7 9 0 9 7 9 9 1 9 12 0 0 1 9 9 9 9 7 1 9 9 9 7 9 1 9 13 2
13 9 15 9 9 9 9 1 9 0 9 9 13 2
49 9 9 0 15 14 1 9 0 1 9 9 9 7 9 0 14 1 9 9 7 9 9 1 9 13 7 3 1 1 9 9 1 9 9 7 9 9 9 9 1 9 9 9 1 9 9 0 13 2
16 10 9 16 0 9 0 1 9 0 9 9 1 9 9 13 2
48 9 3 1 9 9 1 9 9 9 9 9 9 1 9 13 7 1 9 3 1 9 7 9 0 1 9 9 2 9 9 7 9 9 9 13 7 1 9 12 1 9 1 9 9 9 0 13 2
32 9 9 9 1 9 9 9 0 7 0 7 12 9 9 1 9 9 2 9 9 0 7 9 1 9 0 0 14 1 9 13 2
15 0 9 0 9 2 9 0 2 9 9 2 1 9 13 2
12 9 1 9 0 9 9 1 9 15 9 13 2
4 9 2 9 2
37 0 1 9 9 9 0 7 9 0 9 2 12 9 9 16 1 9 9 1 9 13 13 2 9 9 1 9 0 15 1 9 9 9 9 9 13 2
28 1 12 9 10 9 9 12 9 0 1 9 7 9 7 1 9 0 15 9 12 9 0 1 9 9 13 13 2
23 10 9 1 9 9 12 1 9 0 13 13 7 3 1 12 9 9 7 0 1 13 13 2
32 10 9 9 1 9 0 1 9 9 0 7 9 0 3 1 9 0 9 9 13 16 9 1 9 9 9 16 1 15 9 13 2
32 9 1 9 9 9 9 1 9 0 1 9 2 9 9 2 9 2 1 9 9 0 9 2 1 9 9 7 9 9 9 13 2
61 10 9 16 1 9 9 0 9 7 9 9 0 1 9 9 9 9 9 2 9 2 0 13 2 12 9 9 14 1 9 9 2 9 2 0 2 9 0 2 9 7 9 7 9 1 9 9 2 9 2 9 2 9 7 9 1 15 9 13 13 2
12 9 9 9 9 1 12 9 0 14 9 13 2
64 1 9 9 9 9 9 9 9 1 9 9 9 9 12 9 0 2 0 1 9 9 9 16 1 9 9 9 0 15 13 1 9 9 9 13 13 16 1 9 15 1 9 9 9 9 13 2 7 9 9 10 9 14 9 13 7 9 13 1 1 9 9 13 2
23 7 3 1 9 0 9 1 12 9 0 9 13 16 1 12 9 1 9 9 9 9 13 2
14 9 0 3 2 9 0 7 0 0 9 9 9 13 2
34 10 9 3 9 0 0 1 9 9 0 9 14 1 9 9 2 1 9 13 13 7 3 16 9 9 9 14 1 9 15 9 13 13 2
30 15 16 9 13 3 3 1 9 1 9 9 1 9 13 7 9 13 1 9 9 9 9 2 12 9 14 1 15 13 2
30 9 9 9 1 9 9 9 0 13 7 9 14 1 9 1 9 9 13 16 10 9 14 1 9 1 9 1 9 13 2
34 9 9 9 13 2 9 9 0 9 9 1 0 9 9 9 0 9 9 9 1 9 12 16 1 9 9 9 0 4 13 2 9 13 2
19 10 9 9 13 1 9 12 1 12 9 9 9 0 1 9 9 0 13 2
45 9 9 0 9 9 16 1 9 3 10 9 3 9 9 7 9 9 0 14 1 15 9 13 13 2 9 3 1 9 0 9 16 1 9 9 9 9 0 13 2 1 9 9 13 2
33 9 0 9 9 0 9 9 1 9 9 1 9 0 1 9 2 1 9 12 7 12 9 9 1 9 9 0 9 9 0 4 13 2
14 9 9 9 1 12 9 9 7 1 12 9 0 13 2
55 9 9 9 13 2 1 9 0 9 9 0 9 9 1 9 1 9 0 1 9 2 9 16 1 9 3 9 0 9 9 13 7 7 9 16 9 9 1 9 0 9 0 7 0 9 14 1 9 3 13 2 13 9 13 2
16 9 9 9 0 9 9 1 9 9 12 9 9 0 9 13 2
45 1 10 9 12 9 9 9 9 2 9 9 2 9 9 2 9 9 2 9 9 2 9 9 9 2 9 9 2 9 9 2 9 9 2 9 9 2 9 9 7 9 9 9 13 2
49 1 0 9 10 9 12 9 1 9 9 1 9 9 7 9 0 13 16 9 0 1 9 0 9 4 13 2 9 9 1 9 9 9 2 16 9 10 9 1 9 9 9 1 9 0 9 4 13 2
28 1 9 0 10 9 9 9 9 2 9 9 2 9 9 7 9 9 1 9 9 13 7 1 9 0 9 13 2
25 9 9 9 0 9 9 0 9 9 14 16 1 9 12 9 0 13 2 9 9 9 1 9 13 2
4 9 2 9 2
28 0 9 9 13 16 9 9 1 9 9 12 2 12 9 9 13 7 1 10 9 9 9 0 9 9 9 13 2
28 9 9 0 9 9 9 9 13 2 9 1 9 2 1 9 12 1 9 9 9 9 1 1 9 9 13 13 2
36 10 9 13 2 9 9 1 9 1 1 9 9 7 9 16 1 9 0 1 9 12 2 12 7 12 2 12 9 13 13 16 9 9 0 13 2
4 9 2 9 2
41 12 9 0 9 9 13 2 1 9 7 1 9 12 0 2 12 2 12 9 9 9 10 9 1 9 9 13 2 10 9 1 9 12 1 12 2 12 9 9 13 2
25 9 9 1 9 9 1 10 9 13 2 1 9 0 1 9 0 12 9 9 0 1 9 9 13 2
12 1 9 7 0 10 9 1 9 12 9 13 2
6 9 2 9 0 9 2
23 9 9 9 4 1 12 9 9 9 9 0 9 9 0 9 0 7 9 1 9 0 13 2
30 1 9 9 9 9 9 2 9 1 9 16 1 9 9 9 13 7 7 3 0 1 9 13 2 1 10 9 9 13 2
18 15 13 9 9 1 9 9 0 1 9 9 7 0 10 9 9 13 2
8 9 10 9 14 9 13 13 2
16 9 0 9 9 1 9 9 1 9 9 0 9 9 9 13 2
26 10 9 1 9 12 9 1 9 12 9 1 9 9 2 9 2 9 7 9 1 9 12 9 0 13 2
21 9 1 10 9 1 12 9 7 1 9 9 12 1 12 9 1 9 1 15 13 2
38 9 9 9 0 1 9 9 10 9 1 9 9 9 0 13 2 9 1 9 10 9 9 7 9 9 1 9 9 0 7 0 9 9 1 9 9 13 2
42 9 9 13 2 1 9 16 9 9 9 0 1 9 9 1 9 9 13 0 13 16 1 10 9 7 10 9 1 9 16 9 9 1 9 7 9 14 13 2 9 13 2
23 9 9 9 0 0 9 13 2 1 9 9 9 9 9 0 9 15 9 9 9 15 13 2
35 10 9 1 9 0 16 9 9 0 13 13 2 9 9 9 3 9 9 9 9 9 1 9 9 0 9 9 9 9 1 9 9 9 13 2
21 9 9 16 1 9 0 9 9 1 1 9 9 9 9 13 2 1 9 9 13 2
29 9 9 9 1 9 12 9 13 7 9 9 15 1 0 9 9 9 9 1 9 9 9 9 9 9 9 13 13 2
30 0 13 9 9 16 1 9 9 1 9 9 9 9 13 7 1 0 9 0 1 10 9 9 9 9 7 9 9 13 2
4 9 14 13 2
25 9 1 9 1 12 9 9 0 7 0 1 9 9 13 7 12 9 0 0 7 12 9 14 13 2
32 9 10 9 9 13 16 9 10 9 3 0 13 7 16 9 14 9 13 1 9 0 0 9 0 13 7 0 1 9 9 13 2
10 3 0 13 9 15 14 1 9 13 2
38 9 10 9 9 13 16 10 9 0 14 3 1 9 9 1 9 9 13 13 7 1 9 9 13 16 15 14 3 1 15 7 9 9 13 1 15 13 2
30 10 9 0 12 0 9 12 0 13 7 1 9 12 0 15 16 9 0 7 9 15 13 9 15 14 0 9 9 13 2
7 9 0 1 9 0 13 2
4 9 2 9 2
27 0 1 12 12 9 1 9 9 1 9 9 9 16 9 9 9 0 15 13 2 9 9 1 9 0 13 2
44 9 9 9 9 9 9 9 9 9 1 9 1 9 10 9 13 2 9 9 9 13 16 12 9 1 9 9 0 9 9 9 9 9 10 9 9 9 2 9 2 14 0 13 2
27 1 9 12 1 9 9 2 3 12 9 1 9 10 9 0 7 0 9 1 15 1 9 1 9 0 13 2
25 9 16 9 9 9 9 0 9 9 14 1 9 1 13 7 1 9 13 16 9 15 14 9 13 2
8 9 0 9 0 1 9 0 9
4 9 2 9 2
26 9 0 9 0 1 9 0 9 1 9 9 9 3 9 13 7 9 0 1 10 9 9 0 9 13 2
37 1 9 9 0 9 2 9 9 0 1 12 9 1 9 9 9 1 9 9 2 1 12 9 3 9 13 7 9 0 1 10 9 3 9 13 13 2
25 9 0 9 9 13 2 1 9 0 9 0 1 12 12 9 0 9 2 13 7 7 9 13 13 2
22 1 9 0 9 0 7 9 9 15 9 1 9 13 7 9 15 14 12 9 0 13 2
18 15 1 9 3 9 9 7 9 9 14 1 9 9 9 0 13 13 2
20 10 9 0 1 0 9 0 9 1 9 0 1 12 0 9 0 9 13 13 2
17 1 9 9 10 9 0 2 9 9 14 1 9 12 9 9 13 2
9 9 1 9 12 0 1 9 13 2
4 9 2 9 2
26 9 1 9 12 2 12 9 1 9 9 9 9 1 9 9 1 9 13 7 3 12 0 1 9 13 2
41 1 9 9 9 7 9 9 9 9 9 9 9 1 9 1 9 9 9 2 10 9 9 12 2 12 9 9 9 1 9 9 1 9 9 1 9 9 1 9 13 2
29 9 9 1 9 13 16 10 9 3 1 10 9 9 13 13 16 9 9 0 9 0 9 9 1 12 9 0 13 2
18 1 9 9 0 0 7 9 9 2 3 12 9 1 10 9 0 13 2
21 9 1 1 9 10 9 7 9 2 9 0 16 1 9 0 1 9 0 13 13 2
34 1 9 12 9 9 9 9 1 9 2 9 10 9 9 16 0 1 9 9 0 13 2 3 0 13 7 9 4 9 1 15 9 13 2
30 9 9 9 9 9 9 9 9 7 9 0 9 9 14 9 13 7 9 9 9 0 9 0 1 10 9 14 0 13 2
40 1 9 9 9 9 9 9 1 9 1 9 0 4 1 9 9 9 1 9 13 7 1 9 9 9 9 9 9 2 9 9 1 9 9 0 0 9 4 13 2
10 9 9 9 9 0 3 9 4 13 2
40 9 14 9 13 7 16 1 9 1 10 12 9 0 2 16 0 13 16 9 0 7 9 13 12 9 0 2 1 9 13 13 7 9 0 0 1 9 9 13 2
52 3 9 0 7 0 16 1 9 0 1 9 9 13 13 9 1 15 13 16 1 9 9 1 10 12 9 0 2 15 16 9 13 9 13 2 10 9 0 0 13 16 13 4 1 9 12 9 0 9 0 13 2
60 9 3 15 3 9 9 0 9 13 16 1 9 0 9 9 7 9 1 9 9 2 9 0 9 14 0 1 9 13 7 16 9 9 1 9 0 15 2 9 13 16 4 9 9 14 0 7 0 13 3 15 7 15 14 1 9 2 9 13 2
50 3 15 16 10 9 1 9 9 13 2 9 10 9 0 14 16 1 15 0 13 7 1 9 9 13 16 9 0 15 9 13 3 7 3 9 1 1 0 9 9 16 9 0 9 7 9 9 15 13 2
19 9 9 0 9 9 9 13 16 9 9 9 0 1 9 9 0 9 13 2
33 10 9 13 13 2 9 9 9 13 2 1 0 9 9 9 0 1 9 0 9 13 9 9 9 9 1 9 9 9 0 9 13 2
37 1 9 9 9 9 2 9 16 1 9 9 9 9 13 13 2 3 12 1 12 9 1 9 1 10 9 9 13 7 1 9 16 9 9 9 13 2
43 15 13 2 3 9 9 0 1 9 0 1 9 0 9 13 16 10 9 1 9 15 13 16 16 9 9 1 10 9 9 13 7 7 9 9 9 0 14 1 9 4 13 2
36 9 0 13 2 16 10 9 9 0 2 9 9 7 9 16 9 15 1 12 1 12 9 4 13 13 1 9 9 9 13 2 15 9 9 13 2
35 9 9 9 16 1 9 9 0 15 13 2 3 9 0 1 9 15 16 3 9 9 9 9 1 9 0 14 1 9 4 13 2 0 13 2
27 9 15 0 13 16 9 9 0 9 13 9 9 9 9 13 7 1 9 9 0 1 9 7 9 9 13 2
43 12 9 0 1 9 15 13 2 1 9 9 10 9 9 0 3 9 9 9 2 9 7 9 9 0 13 7 3 1 9 9 13 16 1 1 9 7 9 12 9 9 13 2
20 12 9 0 9 16 9 9 13 2 9 9 1 9 9 0 9 9 9 13 2
58 1 10 9 16 1 9 9 0 9 9 13 2 9 9 9 10 9 2 1 10 9 16 9 9 9 1 9 0 9 9 9 9 9 13 2 10 9 14 1 15 9 13 7 13 2 9 0 9 1 1 1 9 9 9 15 9 13 2
51 9 9 1 9 9 13 2 0 9 0 15 14 1 9 9 0 13 16 9 13 9 9 9 9 2 9 9 1 9 1 9 9 0 9 2 9 0 14 1 9 0 9 0 0 3 1 9 9 9 13 2
36 1 10 9 2 9 1 9 1 9 9 9 9 9 1 9 13 2 10 9 16 1 9 9 1 9 13 2 9 9 7 9 15 9 4 13 2
26 15 13 2 9 0 9 1 9 7 9 9 9 9 13 7 9 9 16 4 1 1 9 9 9 13 2
30 9 9 16 13 2 0 9 9 1 9 9 9 9 9 13 7 1 9 0 12 12 9 0 1 9 9 0 9 13 2
35 9 0 0 9 9 9 9 9 9 9 9 1 9 9 9 0 13 7 1 15 9 9 9 2 9 9 7 9 9 1 9 15 0 13 2
31 1 0 9 9 9 9 1 9 9 9 1 9 12 1 12 9 13 7 1 9 9 9 9 1 9 0 10 9 9 13 2
48 3 7 1 9 0 9 9 9 1 9 1 9 9 9 1 9 12 1 12 0 13 7 9 1 9 0 13 7 1 10 9 10 9 9 9 9 1 9 12 1 12 1 9 9 9 0 13 2
20 9 9 9 9 9 1 10 9 0 9 15 14 1 9 9 9 9 4 13 2
18 9 9 3 1 15 1 9 9 9 7 9 9 9 14 0 13 13 2
26 1 9 9 1 9 0 16 15 9 1 9 9 13 13 7 9 9 1 9 13 13 2 9 13 13 2
22 9 1 9 0 7 0 16 1 9 9 1 9 9 0 7 1 1 9 0 13 13 2
9 9 7 9 7 9 15 0 13 2
16 3 9 15 9 9 13 16 9 7 9 14 1 9 9 13 2
19 7 16 1 9 9 12 9 9 13 16 3 9 1 1 15 1 9 13 2
47 7 16 1 9 9 9 9 7 9 9 13 3 9 13 9 3 0 7 0 1 9 14 13 16 9 0 9 7 9 15 14 1 9 9 7 9 9 1 9 1 9 9 1 9 15 13 2
35 9 16 15 14 1 9 12 9 1 9 9 7 9 1 9 9 9 9 13 7 9 15 14 13 7 1 9 9 9 9 1 9 9 13 2
29 1 10 9 16 16 13 9 0 9 1 9 9 13 13 1 9 0 9 7 1 9 0 1 9 7 9 15 13 2
16 3 15 12 9 0 13 16 1 1 9 1 3 1 9 13 2
65 15 9 1 9 15 10 9 13 2 1 9 9 9 9 0 13 0 1 9 0 7 12 12 9 3 0 0 7 1 1 9 9 16 9 1 9 13 1 9 9 9 0 9 9 0 13 2 9 9 1 0 13 13 7 0 9 9 9 0 1 9 9 13 13 2
76 15 0 9 1 15 1 0 9 9 9 9 13 7 3 3 9 9 13 7 0 13 13 10 9 14 1 9 13 7 1 13 2 7 9 13 15 13 1 9 9 9 0 9 4 13 7 9 0 13 16 10 9 1 9 10 9 13 16 9 9 3 9 13 7 1 9 9 7 9 9 1 9 15 13 13 2
35 12 2 13 3 10 9 9 0 1 9 9 9 13 7 16 3 13 3 0 13 9 1 15 14 13 7 1 9 9 9 1 13 7 13 2
26 1 9 12 1 9 9 9 13 1 9 9 9 9 7 9 15 1 9 7 9 7 15 9 9 13 2
25 1 9 12 9 0 1 9 7 9 0 12 9 9 9 0 1 9 9 9 2 9 9 9 13 2
58 9 1 3 9 13 16 1 1 15 13 13 2 10 9 9 0 16 1 9 9 0 13 7 9 15 14 9 9 1 9 9 9 9 1 9 13 13 1 9 0 9 1 9 9 9 1 9 9 9 9 9 13 2 1 12 9 12 2
43 12 2 1 9 1 9 9 16 1 9 2 1 9 1 9 9 9 2 9 9 2 9 9 9 9 2 9 13 13 9 15 14 1 9 9 13 16 1 9 0 13 13 2
34 3 10 9 16 1 12 13 13 13 9 9 14 1 10 9 9 13 16 9 9 15 14 13 7 9 15 14 13 7 1 9 13 13 2
14 9 1 12 1 9 1 9 13 7 1 3 1 9 2
9 9 10 9 9 0 1 3 13 2
19 9 15 1 9 0 9 1 12 9 0 1 9 0 15 3 7 0 13 2
65 16 9 9 2 1 9 9 9 2 3 1 9 0 13 2 7 3 1 9 9 9 13 9 16 1 9 3 9 7 9 3 1 9 7 9 9 0 9 13 2 7 9 15 16 9 13 7 7 1 9 9 0 16 1 9 1 9 9 9 0 9 13 2 13 2
37 10 9 9 9 9 0 16 1 9 9 0 3 0 13 7 1 9 0 16 3 1 9 0 9 10 9 1 9 0 9 13 2 15 14 9 13 2
28 3 10 9 16 9 15 3 1 1 9 0 0 13 13 2 3 16 1 9 15 7 1 9 9 0 9 13 2
70 10 9 9 0 16 13 2 1 1 9 1 10 9 16 9 3 9 9 13 2 9 16 13 16 1 9 9 0 16 1 3 7 3 1 1 9 9 1 9 7 9 9 13 9 13 16 9 15 9 15 14 1 15 13 7 4 1 9 9 0 15 3 1 9 9 15 15 9 13 2
27 16 10 9 7 7 10 9 0 13 7 10 12 9 13 16 9 7 9 15 15 14 1 9 9 0 13 2
19 1 3 4 1 12 9 0 0 9 9 13 16 1 9 9 9 9 13 2
23 9 9 9 9 2 9 9 9 14 1 9 9 9 1 9 9 7 1 9 12 9 13 2
36 10 9 16 1 9 1 9 9 1 9 7 9 1 9 9 9 13 2 12 1 0 9 13 16 1 3 1 9 1 9 9 0 0 13 13 2
33 9 9 9 16 9 9 14 16 1 9 15 1 9 0 1 9 13 13 2 9 7 1 9 9 7 9 9 9 15 0 13 12 2
52 9 9 9 1 9 9 9 9 9 1 10 9 0 13 16 9 9 9 1 9 9 0 16 9 1 9 9 13 13 7 10 9 1 9 16 1 9 0 13 3 13 13 9 9 9 14 1 10 9 0 13 2
32 16 9 0 9 0 1 15 1 9 9 0 15 9 13 2 9 9 0 9 7 9 1 1 1 9 0 1 15 0 9 13 2
33 1 0 16 1 9 3 1 9 0 1 0 1 9 0 13 2 3 7 3 9 9 7 9 0 9 0 7 1 0 9 9 13 2
49 1 10 9 7 1 9 0 9 7 9 2 9 7 9 9 0 9 1 9 0 1 9 9 2 9 9 1 1 9 9 9 15 2 7 9 1 9 9 9 0 15 1 9 9 9 3 0 13 2
18 1 3 9 9 1 9 7 9 13 16 15 14 1 9 15 13 13 2
