1957 11
20 7 13 16 13 9 0 1 12 9 7 13 0 1 12 9 13 3 9 9 13
23 7 13 7 3 9 0 7 15 13 1 15 13 9 7 13 13 15 9 7 13 13 16 13
10 7 16 13 9 0 13 0 9 13 13
29 7 13 0 9 0 7 15 13 1 15 13 13 15 16 13 9 1 9 7 16 3 15 13 7 13 13 15 9 0
26 7 16 13 9 0 13 0 9 13 13 7 13 7 3 9 0 7 15 13 1 15 13 9 1 9 0
23 7 13 3 9 1 9 12 9 13 9 9 9 7 12 9 9 9 7 9 7 9 3 13
13 7 16 13 9 0 13 9 0 9 13 13 7 13
32 7 3 9 0 7 15 13 3 9 15 9 7 0 13 15 7 13 13 15 9 1 12 9 9 13 9 9 7 9 7 9 9
18 7 16 13 0 9 13 1 9 9 9 1 9 9 7 1 9 15 13
29 7 13 13 15 0 9 0 7 13 13 15 16 13 9 3 0 16 13 9 15 7 9 15 15 13 13 16 7 15
26 7 13 16 13 9 0 7 9 13 13 0 7 9 13 13 0 3 9 0 7 9 0 13 13 16 9
15 7 9 9 13 1 9 16 9 13 9 0 16 9 0 13
16 7 9 13 16 9 13 7 0 9 7 9 1 9 0 13 13
23 7 9 9 7 9 7 9 7 9 7 9 7 0 9 7 9 13 15 1 9 7 9 9
20 7 13 9 7 9 13 1 15 7 13 15 1 9 13 1 9 7 1 9 9
28 1 15 13 12 9 13 1 12 9 9 13 12 9 9 16 13 9 1 9 7 3 1 9 7 3 1 0 9
25 7 13 0 9 13 1 9 9 13 9 9 0 7 13 9 0 12 9 15 13 13 13 9 7 9
14 7 13 9 0 13 9 9 0 15 13 1 9 7 9
23 7 0 9 13 1 9 9 7 9 7 12 9 7 13 1 9 9 1 9 0 7 13 9
18 7 13 0 1 9 13 15 15 15 13 13 9 0 15 13 7 3 13
27 7 13 15 9 0 15 13 7 13 15 15 13 15 13 1 9 0 7 13 9 0 7 13 15 1 9 9
22 3 13 1 9 9 7 13 15 9 7 9 1 9 15 7 15 13 1 9 13 1 15
16 3 13 7 3 13 3 7 3 13 1 15 9 7 3 0 9
13 7 16 13 9 0 13 13 9 1 9 3 0 9
14 7 13 12 9 13 1 9 9 7 13 13 15 12 9
29 7 0 9 13 7 13 1 9 13 9 0 7 13 13 15 9 0 16 13 9 9 0 1 9 0 15 13 1 9
12 7 13 9 9 1 9 9 1 9 9 1 9
24 7 13 9 9 7 13 15 1 9 9 7 13 1 9 7 13 13 9 7 9 7 9 7 9
12 7 12 9 15 13 12 9 13 15 16 9 13
36 7 0 9 13 7 13 13 9 7 9 13 1 9 7 13 13 1 9 7 0 9 9 13 13 7 0 9 9 13 13 7 0 9 0 13 13
22 7 0 9 9 13 7 3 9 0 9 13 13 13 1 9 7 13 13 0 9 9 9
14 7 13 13 0 9 9 15 13 9 7 0 3 9 13
24 7 0 9 9 13 7 13 1 9 9 0 13 3 9 7 13 1 0 9 9 7 1 9 9
24 7 9 9 13 9 7 13 13 0 9 9 1 9 7 0 9 13 13 1 9 16 0 13 13
33 7 0 9 9 13 7 13 13 0 9 9 7 0 9 9 7 0 9 9 16 13 0 9 15 7 9 3 13 9 0 7 9 3
30 7 13 7 13 9 0 9 13 1 0 9 13 9 0 6 6 6 13 1 9 1 0 9 9 12 9 15 13 9 13
20 7 0 9 9 13 7 13 9 1 9 13 1 9 7 13 13 15 9 9 9
21 7 13 9 9 7 13 9 9 16 9 9 0 7 13 13 9 7 9 1 9 9
17 7 1 9 13 8 1 9 7 13 13 15 9 16 13 9 9 9
26 7 13 13 15 3 13 9 9 7 3 0 9 7 3 0 9 16 3 9 15 3 13 9 9 1 9
21 7 13 13 15 16 13 15 7 16 13 9 8 7 9 15 16 9 9 16 13 9
19 7 1 9 15 13 9 9 7 3 13 15 7 13 13 7 13 9 1 15
12 7 13 9 16 9 9 7 9 15 16 9 13
18 7 13 9 16 9 0 7 9 9 15 16 9 9 9 0 13 1 9
16 7 13 9 0 8 7 9 1 9 15 9 15 13 9 9 8
18 7 0 9 9 13 7 13 9 0 1 9 9 0 15 13 1 9 9
21 7 13 13 12 9 15 13 13 1 9 7 9 7 9 7 9 16 13 0 9 9
35 7 3 13 9 1 9 7 15 13 1 15 13 9 0 7 0 7 0 7 9 9 13 3 9 9 7 1 9 15 13 9 7 9 7 9
22 9 7 9 1 9 15 13 7 1 9 15 16 9 15 0 9 13 9 7 1 15 13
44 7 0 9 15 3 13 13 1 15 9 7 3 9 13 1 9 9 0 16 3 13 9 7 9 0 7 0 7 0 7 0 7 0 8 7 3 13 13 7 3 13 7 3 13
22 7 3 13 9 1 9 0 7 3 1 9 0 7 3 1 9 0 7 3 1 9 0
18 7 13 1 9 0 9 13 7 13 9 0 0 1 9 0 7 1 9
17 7 13 9 0 3 16 9 13 7 16 13 13 13 12 9 9 0
24 7 16 13 13 12 9 13 13 7 13 9 1 9 13 13 15 13 13 12 9 7 13 15 13
15 7 9 15 13 13 1 9 7 1 9 13 9 0 1 9
36 7 13 1 13 1 9 9 15 13 9 7 15 15 1 15 13 7 9 7 15 15 1 15 13 7 9 7 15 1 3 13 16 9 3 3 13
30 7 13 1 9 13 15 16 13 15 9 7 13 15 13 7 13 15 7 13 13 9 0 7 1 9 0 13 0 3 9
25 7 13 9 1 9 9 7 13 15 7 13 1 9 0 3 9 0 7 16 13 15 13 13 9 0
15 7 13 15 13 15 3 13 9 7 9 7 9 7 9 0
19 7 13 13 15 9 0 9 13 13 7 13 9 9 7 9 7 13 1 15
23 9 7 15 13 3 9 13 3 7 3 13 15 16 13 13 9 7 9 13 13 9 12 0
13 7 13 0 9 0 7 13 9 12 0 12 13 9
12 15 13 0 9 7 0 9 1 9 9 9 13
25 7 16 15 15 13 13 9 13 1 9 15 7 13 9 15 7 16 15 13 15 13 3 13 15 13
26 15 13 9 13 9 16 13 9 9 15 7 9 13 1 9 13 15 1 9 7 13 9 0 9 3 13
20 7 16 13 9 0 9 15 13 1 9 13 1 15 9 7 13 15 7 13 15
25 7 13 1 9 7 9 7 9 7 9 9 15 1 12 9 7 9 7 9 15 3 13 13 1 9
22 7 13 9 13 1 15 7 13 7 9 13 3 16 15 0 9 13 15 15 13 1 9
27 7 1 9 12 7 9 9 9 1 9 13 1 15 7 13 1 9 0 7 9 0 13 1 15 15 13 15
21 7 13 9 0 1 9 13 15 13 3 7 13 1 9 1 9 7 13 15 9 15
33 7 1 15 9 13 13 9 0 7 0 9 9 13 7 13 13 1 9 9 9 12 12 7 0 1 9 13 13 7 13 9 9 9
28 7 0 9 9 13 7 13 13 9 0 1 9 13 13 13 9 15 9 9 0 7 9 15 7 13 1 9 9
19 7 12 12 9 15 1 9 9 13 1 9 0 13 1 9 0 7 13 9
11 7 1 9 13 7 13 13 7 13 16 13
24 7 13 13 0 9 1 9 7 3 9 0 0 13 9 12 7 9 12 7 1 9 0 12 9
27 7 9 15 13 0 9 9 9 7 13 15 1 9 7 9 13 1 9 15 13 13 16 16 13 9 15 13
23 7 13 9 0 15 13 13 0 9 1 9 0 7 13 13 9 15 1 9 7 1 9 15
19 7 9 13 1 9 3 13 9 13 1 9 16 3 13 15 9 12 0 12
19 7 13 13 9 1 9 9 7 9 15 13 1 9 7 9 13 7 9 15
12 7 3 13 7 3 9 13 13 15 3 1 9
37 7 13 9 0 1 9 13 3 13 13 9 7 9 7 9 9 0 7 9 9 15 16 13 13 9 9 0 15 13 15 1 9 9 0 9 7 9
20 7 15 13 15 1 9 9 7 1 9 9 0 7 3 13 9 0 3 1 9
25 3 13 9 7 15 13 1 15 6 9 7 9 16 13 9 1 15 13 9 0 13 16 0 9 13
15 7 16 13 9 16 13 13 1 9 13 13 9 15 13 0
27 7 13 13 9 0 9 9 0 16 13 1 9 1 9 0 3 13 1 9 7 9 7 0 9 1 9 9
17 7 13 9 1 9 0 1 9 9 3 9 16 15 13 13 1 9
18 7 13 9 9 7 13 9 9 0 7 13 9 15 13 9 1 9 0
23 7 13 13 9 1 9 7 13 13 9 1 0 1 9 15 15 13 9 9 7 13 9 9
5 7 13 1 9 9
24 7 13 1 9 9 13 13 9 12 7 9 12 7 1 9 15 12 9 7 1 9 15 9 9
22 7 0 1 9 0 3 13 1 9 7 9 9 15 13 13 7 13 13 0 9 1 9
20 7 13 9 16 13 9 9 7 13 9 13 15 0 9 7 15 13 13 1 15
18 7 13 13 15 9 13 0 7 9 7 13 13 15 9 13 9 12 9
20 7 13 9 0 1 9 1 9 13 9 15 7 9 15 7 15 15 1 9 13
25 7 13 13 15 9 13 1 9 7 13 15 7 13 13 15 9 1 0 9 7 9 7 9 7 9
22 7 13 15 0 15 13 9 15 3 13 13 9 1 9 9 9 15 13 13 1 9 9
5 16 15 13 9 13
17 7 13 0 9 13 1 9 7 13 9 0 0 9 7 13 16 9
24 7 9 0 9 0 13 1 9 15 7 13 9 7 13 1 15 13 9 0 15 13 13 9 9
16 7 13 9 0 16 3 9 13 1 9 13 1 9 1 9 9
28 7 13 13 9 1 9 15 13 13 15 13 1 9 9 13 13 1 9 16 13 9 9 15 13 9 9 7 13
22 7 13 13 15 16 13 9 9 9 16 7 13 9 9 7 13 15 3 13 9 9 13
23 7 13 0 0 7 0 7 0 7 0 7 0 7 0 13 9 1 0 9 7 1 9 0
20 15 9 13 15 13 9 13 9 9 9 7 9 13 7 9 15 13 0 12 12
27 7 13 7 3 9 13 1 9 9 7 1 15 12 12 12 12 13 9 15 7 9 9 15 13 1 9 0
24 7 13 9 1 9 3 9 9 0 7 3 9 9 0 7 9 15 13 16 9 13 1 9 0
29 7 13 3 9 0 1 9 7 1 12 9 7 9 7 9 13 13 9 16 15 12 12 12 0 15 13 13 1 9
11 7 1 9 15 3 13 13 9 1 9 13
26 7 13 0 9 13 1 0 9 13 9 0 16 13 13 1 9 7 1 0 9 7 9 7 9 7 9
20 7 0 9 13 13 13 13 13 9 15 0 15 1 9 9 9 0 13 0 9
27 7 0 9 0 13 13 15 13 9 0 16 15 13 9 7 9 15 7 13 9 1 9 0 7 1 9 0
28 7 15 13 1 9 9 9 15 13 13 9 1 9 9 15 7 13 9 7 9 1 9 9 13 7 1 9 9
27 7 9 9 15 1 9 9 13 7 13 9 9 7 9 15 13 9 7 9 15 7 16 15 13 9 9 15
11 15 9 9 13 15 13 9 9 7 9 9
27 7 13 9 1 9 13 13 0 0 15 1 9 13 3 3 13 9 16 13 1 9 0 9 16 15 13 15
25 7 13 7 3 9 0 7 1 9 13 0 9 9 13 1 9 0 9 0 7 1 9 0 9 0
27 7 0 9 13 1 9 13 9 0 1 13 1 9 13 9 0 7 13 16 13 9 16 13 16 13 9 9
14 7 13 15 13 1 9 9 0 1 9 7 13 13 9
15 7 0 9 13 1 9 15 13 1 9 13 7 15 9 0
18 7 13 9 9 0 1 9 7 13 9 9 7 13 1 9 9 9 0
19 7 13 13 9 1 9 7 13 9 1 9 3 1 9 9 1 9 12 0
26 7 13 3 9 0 13 9 7 15 15 13 9 7 9 15 7 9 9 15 13 1 9 9 13 9 9
25 15 3 13 9 7 13 9 0 16 0 0 16 0 9 13 7 13 1 9 0 16 9 0 13 13
13 7 1 15 13 7 3 13 13 9 9 9 1 9
19 7 13 12 9 13 12 9 1 9 13 9 0 0 7 13 1 9 9 0
18 7 0 1 12 9 13 12 9 12 9 0 0 9 9 13 1 9 9
24 7 13 13 9 9 1 9 9 7 1 9 15 7 9 13 13 1 9 16 13 12 9 12 9
18 7 13 9 0 1 9 13 12 9 13 7 13 12 9 9 9 1 9
28 7 13 0 7 13 9 0 1 9 7 13 13 9 0 7 0 1 9 15 13 9 9 7 15 15 13 9 15
21 7 0 13 9 0 1 9 7 13 13 9 3 0 7 0 9 13 13 13 1 9
15 7 0 13 9 0 1 9 7 1 9 9 7 13 13 9
16 7 13 9 9 13 0 13 15 13 7 15 13 0 16 15 13
13 16 9 9 7 9 13 7 9 15 13 13 0 13
13 7 13 9 13 3 9 9 0 0 7 0 9 0
16 7 0 13 9 0 1 9 7 13 13 15 9 13 9 7 9
22 7 13 9 9 0 7 13 9 9 13 9 1 15 9 7 3 13 9 16 13 15 9
20 7 0 13 9 0 1 9 9 7 13 13 9 15 0 7 13 9 0 1 9
16 7 13 9 9 1 9 7 9 0 7 3 13 9 1 9 0
21 7 0 13 9 0 1 9 15 0 9 7 13 9 15 16 13 9 9 1 9 9
19 7 13 1 9 9 7 1 9 9 7 1 9 9 9 12 0 1 9 9
9 7 13 15 1 9 15 13 9 9
18 7 0 13 9 0 1 9 7 13 9 0 1 9 1 9 13 13 13
26 7 13 13 9 7 9 7 9 7 9 13 13 0 0 3 13 1 3 9 13 1 9 0 9 3 0
27 7 13 13 9 0 1 12 9 7 9 9 13 7 9 0 13 1 9 1 9 13 15 9 9 9 9 15
9 7 0 9 13 7 9 3 13 13
22 7 9 0 16 9 13 1 9 1 9 7 13 9 9 1 9 9 3 0 13 13 3
26 7 13 0 1 12 9 15 13 12 9 7 13 13 15 13 13 13 15 9 9 0 15 13 1 9 0
16 1 15 13 13 9 9 7 13 13 15 13 9 1 9 9 15
23 7 13 15 1 9 1 9 7 13 9 13 1 9 0 0 9 9 13 9 12 7 9 12
27 7 9 13 13 9 7 9 7 13 9 7 9 0 7 9 13 9 0 1 9 0 0 9 7 9 9 15
20 7 13 9 0 1 9 9 7 1 9 9 9 7 13 13 16 13 15 9 0
23 7 13 15 9 3 13 15 15 13 9 9 7 9 15 13 15 15 13 9 12 7 12 9
38 9 15 13 13 7 3 13 7 13 13 1 9 7 1 9 13 7 13 13 9 15 3 13 13 9 1 9 9 1 9 9 13 9 16 13 7 3 13
20 7 15 13 9 15 13 9 12 9 12 9 13 1 15 9 13 7 9 12 13
15 12 13 0 13 0 3 13 7 16 13 13 15 0 9 13
19 7 9 15 13 7 3 13 7 15 0 13 7 1 12 13 7 1 9 13
21 7 12 9 15 13 12 9 13 15 9 3 13 7 9 3 9 0 9 13 1 9
11 15 0 9 13 7 9 7 9 0 9 13
25 15 1 9 13 7 9 13 15 3 9 9 13 7 9 9 7 15 1 15 13 13 7 13 7 0
15 7 13 15 9 15 13 3 9 13 9 13 7 9 7 9
13 7 9 15 13 13 9 0 15 13 9 1 9 9
19 7 1 15 13 0 9 13 1 9 13 9 0 7 9 13 13 1 9 15
25 7 13 1 0 9 13 13 13 9 0 7 13 13 9 9 7 9 0 9 0 7 9 0 9 0
24 7 13 0 9 1 9 13 13 1 15 9 0 16 3 9 13 9 15 7 1 9 15 3 13
18 13 15 16 15 13 7 13 9 1 9 15 1 9 15 13 13 15 3
28 3 13 15 7 1 9 13 3 13 15 9 7 9 16 1 9 0 13 13 9 7 9 3 13 7 9 3 13
23 7 13 7 13 15 1 15 9 9 15 1 15 13 13 7 1 9 13 16 13 9 9 15
14 7 9 9 13 7 13 1 15 3 9 15 9 13 3
22 7 9 0 9 9 13 1 15 7 9 0 7 0 13 1 15 7 3 15 3 3 13
17 9 15 15 0 13 13 1 15 3 13 1 9 9 15 13 7 13
24 3 0 9 13 13 0 9 7 0 9 7 9 15 1 9 13 7 9 7 15 9 13 3 13
12 7 13 13 9 9 15 13 15 0 9 15 0
35 7 13 9 1 9 0 7 13 13 7 13 13 6 6 9 0 1 15 0 13 13 9 15 13 9 1 9 1 9 15 16 0 9 13 13
17 13 1 15 9 7 9 7 9 7 9 3 13 9 9 0 1 15
33 7 9 9 7 9 7 9 13 7 9 3 13 1 15 3 7 0 9 0 9 3 13 1 15 15 7 9 9 3 13 1 15 15
30 7 9 9 3 13 15 3 7 9 9 7 9 3 13 3 1 15 16 9 0 13 9 9 16 1 9 0 13 0 9
16 7 1 15 9 9 7 9 13 13 7 9 15 13 13 1 9
20 1 15 13 3 9 0 9 0 1 9 13 6 9 7 9 7 9 9 0 13
11 7 3 13 6 7 9 15 13 1 9 9
17 7 13 9 12 12 7 12 9 7 13 9 13 1 9 13 3 6
24 7 13 3 9 9 0 7 16 9 9 0 7 16 9 9 0 13 6 16 13 9 9 0 0
16 13 7 13 7 13 9 15 16 13 9 9 7 9 15 13 15
15 7 13 13 15 16 13 15 9 13 0 9 16 9 13 9
20 7 13 15 13 9 8 1 9 9 9 13 13 7 13 15 15 9 0 9 13
31 7 13 1 9 15 16 13 15 7 13 15 13 16 13 9 0 13 7 9 0 13 9 9 9 13 9 16 9 13 9 9
23 7 13 9 13 7 6 9 0 7 15 13 1 15 13 9 7 0 13 7 9 13 7 13
12 7 13 13 9 13 9 7 13 9 15 9 9
15 7 9 15 13 1 9 13 15 1 9 0 13 9 0 0
28 7 1 9 15 13 9 0 16 1 15 13 9 7 15 13 15 1 9 0 7 15 13 9 9 9 9 9 0
14 7 13 1 9 7 1 9 0 13 9 9 7 9 13
25 7 13 0 9 13 1 9 7 13 9 0 13 0 9 15 13 1 9 9 13 13 1 9 0 9
23 7 13 9 7 9 9 7 9 15 13 1 13 9 1 15 15 13 1 9 7 1 9 15
35 7 13 13 9 7 1 15 9 15 13 9 1 15 15 13 15 15 13 9 9 15 7 13 9 15 0 13 13 15 0 1 9 9 13 9
21 7 9 13 13 1 9 13 1 9 15 13 1 9 15 7 0 9 13 13 9 15
15 7 13 9 13 1 9 13 9 9 7 9 0 1 9 0
28 0 7 0 15 13 9 1 9 0 1 15 0 9 3 13 9 7 13 9 9 7 9 7 13 1 15 12 9
12 7 13 1 9 9 7 13 9 9 7 9 13
25 7 13 9 1 9 1 9 7 13 15 7 9 15 13 15 13 13 1 9 9 7 9 3 3 9
23 7 13 9 0 0 7 13 1 15 1 15 9 13 9 7 9 7 9 3 13 13 1 15
36 7 13 9 0 7 0 13 1 9 9 7 9 13 13 7 0 9 13 13 15 13 9 7 13 13 9 1 15 15 13 13 1 9 1 9 15
26 7 13 9 9 15 1 15 13 7 9 7 0 13 9 15 1 15 13 7 13 13 1 9 1 9 15
14 7 15 3 13 13 1 9 9 13 13 13 1 9 9
19 7 13 9 0 7 9 0 0 16 9 7 0 9 13 7 9 3 3 13
17 7 9 0 9 0 13 13 1 9 1 9 13 16 9 13 9 0
29 7 13 9 0 1 9 13 3 9 9 1 9 7 13 1 15 7 15 9 15 13 7 15 9 1 15 13 15 9
27 7 13 9 0 9 1 9 15 7 9 3 3 13 7 3 9 7 3 9 7 3 9 13 3 15 0 13
20 7 13 15 13 1 9 3 0 13 9 7 13 13 16 0 9 0 13 7 0
13 15 13 13 15 7 13 15 9 7 15 13 15 9
30 0 7 7 0 7 9 7 9 7 9 7 9 7 9 7 0 9 9 15 13 1 9 13 9 7 9 15 13 9 0
24 7 13 9 0 7 0 13 9 12 7 1 9 9 12 7 9 13 15 13 9 12 9 9 9
32 7 9 1 9 13 13 7 9 15 0 13 0 7 9 7 13 13 9 1 9 1 9 12 12 9 7 9 7 9 15 0 13
14 7 13 13 9 15 12 12 12 9 9 9 15 13 9
23 7 12 9 12 9 13 1 0 7 0 9 13 1 0 9 7 9 9 9 0 3 9 0
15 7 9 3 13 1 15 9 16 9 0 9 15 13 7 9
22 7 9 3 13 9 7 3 9 16 13 1 15 16 9 9 13 15 7 9 15 13 9
16 7 13 9 1 9 15 7 9 9 13 9 0 7 9 1 15
12 7 9 15 3 13 1 9 9 16 3 13 3
8 7 13 9 7 9 9 1 15
20 7 3 13 1 15 15 9 7 13 9 7 9 16 15 13 13 1 9 9 9
15 7 13 15 9 9 9 0 3 9 13 1 9 9 7 9
19 7 0 9 3 13 3 7 9 9 7 9 1 15 13 7 9 15 13 15
10 7 13 9 15 7 9 15 1 9 15
24 7 9 3 3 13 7 3 13 9 9 7 3 9 9 3 9 9 13 15 7 13 1 9 9
24 7 13 15 15 9 0 7 0 13 7 9 9 9 9 13 9 0 13 9 0 15 13 13 3
11 7 3 13 3 0 15 13 9 9 9 15
13 7 13 15 3 13 9 9 9 15 9 16 3 13
20 15 13 13 3 7 15 1 9 13 13 3 7 0 9 13 3 7 9 13 3
21 7 9 7 9 13 13 7 15 13 13 13 7 15 13 13 15 13 13 9 9 3
22 13 15 0 13 9 9 9 15 16 15 13 1 15 13 9 1 15 9 13 1 9 0
29 7 16 15 13 1 9 9 9 15 13 9 9 15 1 9 9 7 1 9 0 7 1 15 15 13 13 1 9 0
14 16 9 0 3 13 1 9 9 15 0 13 1 0 2
13 13 7 13 1 15 9 9 0 9 9 0 13 2
15 13 3 15 0 7 13 9 9 2 15 3 10 9 13 2
48 7 15 13 1 15 16 9 13 13 1 15 13 2 16 15 9 9 2 16 15 13 2 16 1 0 9 13 4 2 7 2 15 3 0 13 2 16 0 9 3 9 1 0 9 9 13 13 2
30 13 3 9 9 0 1 9 0 13 2 1 9 1 9 3 13 2 13 2 16 1 0 2 15 13 9 9 15 13 2
22 15 7 2 7 15 2 7 16 12 3 13 9 9 2 3 3 1 15 0 9 13 2
47 16 2 1 13 9 13 7 15 9 13 2 13 15 13 15 9 15 9 15 15 9 3 13 2 7 15 9 9 13 2 3 3 13 15 13 9 2 16 13 9 2 7 15 9 13 13 2
11 3 13 7 0 15 9 9 1 9 13 2
8 0 3 9 13 13 1 9 2
9 15 7 9 13 0 9 9 13 2
13 15 3 9 0 3 15 9 13 13 16 9 0 2
7 3 9 0 9 13 13 2
33 15 0 0 15 9 7 15 1 15 13 2 3 13 9 7 9 0 15 13 2 3 1 15 9 15 13 2 7 1 15 15 13 2
22 15 0 2 0 9 3 15 9 13 13 16 0 2 9 15 15 13 2 9 13 13 2
9 15 3 9 9 3 13 1 9 2
2 0 2
6 9 13 9 0 9 2
12 1 13 7 9 3 13 0 9 16 1 9 2
8 3 3 3 1 9 10 13 2
9 3 3 1 15 9 9 9 13 2
2 3 2
9 15 1 15 0 13 16 9 13 2
9 3 13 15 7 1 15 13 13 2
14 1 15 7 16 13 9 9 15 13 2 0 0 13 2
30 13 3 1 15 0 9 9 2 16 3 0 9 9 3 13 2 16 0 13 15 2 9 13 2 15 13 9 3 13 2
6 3 7 1 9 13 2
6 13 0 1 9 10 2
4 3 13 9 2
11 3 13 3 15 9 9 15 1 9 13 2
2 0 2
29 9 15 13 1 9 3 1 0 2 3 1 15 15 0 2 13 0 2 16 9 15 13 1 9 1 15 16 13 2
12 13 3 3 9 1 15 9 13 1 9 3 2
7 0 3 1 0 9 13 2
26 9 7 13 9 9 2 7 0 9 9 13 13 1 15 15 13 9 2 7 3 1 16 13 9 3 2
9 3 9 1 9 9 13 9 9 2
11 3 13 3 13 9 9 1 9 10 0 2
13 16 9 0 3 13 1 9 9 15 13 1 9 2
44 3 2 13 15 15 9 9 2 9 16 13 2 15 1 9 1 9 13 2 1 15 3 1 0 15 9 13 2 1 1 9 13 1 15 0 2 1 15 9 1 15 13 13 2
28 13 3 9 9 13 0 2 0 2 0 2 3 0 2 12 2 7 15 3 2 15 1 9 0 1 9 13 2
17 1 0 7 15 9 9 13 3 0 1 9 2 7 3 1 9 2
19 16 3 0 9 13 13 9 0 2 3 0 15 13 3 13 0 7 0 2
30 7 15 13 1 15 9 0 9 2 16 2 1 9 0 9 1 9 13 2 13 15 13 9 2 7 3 1 15 13 2
22 1 9 7 13 0 9 1 9 2 13 16 13 1 15 13 2 3 15 13 13 0 2
12 15 7 13 0 9 15 1 9 13 1 9 2
11 3 13 7 7 15 1 0 9 9 0 2
16 15 3 15 13 15 9 2 13 1 9 15 9 16 1 0 2
21 15 3 15 13 1 9 2 13 3 7 1 0 2 13 7 1 0 1 15 9 2
14 9 7 13 9 0 9 2 1 10 9 15 0 13 2
19 9 3 13 15 0 9 0 13 10 9 2 16 13 15 9 15 4 13 2
24 1 13 7 9 1 9 13 1 9 9 0 13 2 1 9 15 9 2 15 1 9 9 13 2
11 3 13 3 15 9 9 0 15 0 9 2
2 3 2
14 13 1 9 13 9 13 1 9 2 16 1 13 13 2
18 9 3 2 15 13 0 9 2 13 9 15 3 13 9 1 0 9 2
25 15 7 9 1 9 9 1 9 13 13 3 1 9 1 15 0 1 9 13 2 7 15 0 9 2
17 0 3 13 4 15 1 0 9 13 13 15 15 1 0 13 13 2
9 3 13 3 15 9 0 0 9 2
2 0 2
5 9 10 9 13 2
9 15 3 3 0 7 0 13 13 2
9 9 7 7 9 0 9 9 13 2
8 15 13 3 15 10 0 13 2
13 13 7 9 15 1 9 13 2 0 9 13 13 2
30 15 13 1 0 15 15 0 1 9 1 9 9 13 2 15 2 10 9 13 2 16 9 15 13 2 1 9 0 13 2
24 16 7 15 13 15 3 1 0 9 13 9 9 16 15 9 15 9 13 2 13 15 13 0 2
10 15 3 13 9 2 15 13 0 9 2
12 3 3 13 1 15 9 1 9 0 9 9 2
2 3 2
6 9 1 9 9 13 2
7 1 9 7 9 13 9 2
20 3 13 15 3 13 16 13 16 0 13 15 15 13 2 16 13 1 12 0 2
23 9 7 13 0 9 13 2 15 13 9 9 1 0 15 15 15 1 9 9 13 13 4 2
9 3 13 3 1 15 9 0 9 2
2 3 2
11 9 1 13 4 0 9 2 13 15 9 2
9 0 7 9 10 9 0 13 9 2
18 15 3 9 9 0 13 15 9 2 15 13 3 13 15 0 13 9 2
32 15 7 3 13 9 15 9 1 9 1 9 13 13 2 16 3 2 15 9 13 2 15 13 13 2 15 1 15 9 3 13 2
9 3 13 3 1 15 9 9 9 2
2 3 2
11 9 15 13 1 9 13 16 13 1 9 2
12 1 15 3 13 1 9 2 15 13 1 9 2
16 13 7 15 9 1 9 1 15 16 13 9 1 16 13 0 2
14 15 3 13 13 1 9 15 15 9 13 13 1 9 2
24 3 15 9 13 16 0 1 9 13 2 16 0 2 1 0 13 2 13 1 9 1 0 3 2
18 15 0 15 9 15 3 13 3 1 9 13 2 16 13 1 9 0 2
24 3 1 10 9 13 0 1 9 0 9 13 2 15 15 2 1 15 9 2 3 13 3 13 2
16 9 7 10 13 1 9 1 10 0 2 16 1 0 13 4 2
28 12 7 0 13 3 1 9 0 13 1 9 0 2 15 13 9 2 16 9 3 1 9 0 2 15 13 9 2
14 1 15 13 16 15 9 9 0 13 13 3 1 9 2
12 15 3 13 1 15 0 9 2 15 13 9 2
23 15 7 3 13 13 9 15 1 9 1 9 13 13 2 16 2 15 13 2 3 0 13 2
11 3 13 3 15 9 9 0 1 0 9 2
13 16 9 0 3 13 1 9 9 15 13 1 9 2
23 13 7 7 15 9 9 2 3 1 15 0 9 13 2 15 3 9 1 9 1 9 13 2
43 15 3 3 1 15 9 15 1 9 1 9 13 2 13 2 16 15 1 9 1 9 13 1 15 2 1 15 9 2 9 13 13 3 13 2 16 1 9 15 9 13 4 2
14 3 13 7 0 7 1 15 9 9 0 9 9 13 2
12 9 3 13 9 9 9 2 16 1 13 13 2
25 1 9 7 9 13 9 9 0 3 1 15 15 13 1 9 9 2 16 0 9 13 1 9 9 2
9 3 3 9 13 15 15 13 13 2
12 3 13 3 7 1 15 9 9 0 9 9 2
2 3 2
13 13 4 1 16 0 9 3 13 0 1 9 9 2
8 1 9 7 9 9 13 9 2
22 9 3 13 1 9 15 15 15 13 2 16 13 2 3 7 1 15 9 9 0 13 2
10 3 13 3 1 15 9 0 9 9 2
2 3 2
17 15 13 2 9 13 15 15 15 1 15 13 2 15 15 3 13 2
10 3 9 3 13 9 9 0 16 9 2
24 3 7 13 15 3 13 1 15 13 16 13 15 9 9 13 1 13 16 15 13 15 3 13 2
16 7 3 9 13 13 0 2 7 13 16 13 13 9 9 13 2
19 16 7 16 15 0 13 15 3 1 15 13 2 3 13 15 1 0 13 2
9 13 3 0 7 1 9 9 9 2
15 3 3 13 15 0 1 15 0 2 15 9 9 13 13 2
19 3 13 7 0 9 9 13 0 7 0 2 16 1 13 13 1 9 9 2
17 7 3 2 16 13 0 7 0 2 1 15 9 9 3 13 13 2
11 13 3 15 9 9 1 9 9 9 9 2
25 7 15 9 13 9 0 13 9 2 16 0 13 2 7 1 13 0 13 2 16 13 9 7 9 2
18 1 3 1 0 9 9 9 9 13 2 0 13 16 13 1 9 9 2
2 0 2
12 1 9 2 1 13 0 9 2 0 9 13 2
12 9 7 9 3 13 9 2 7 3 15 13 2
7 16 15 13 13 15 13 2
10 3 13 3 1 9 9 0 9 9 2
2 3 2
16 9 1 9 13 4 9 16 0 9 9 2 3 9 2 13 2
22 1 9 7 9 3 13 9 13 9 13 9 2 16 9 1 13 13 2 3 1 13 2
18 3 7 9 13 12 8 12 2 16 16 1 9 13 2 13 1 9 2
14 13 3 1 9 9 13 9 2 1 0 13 9 13 2
14 1 16 13 8 12 2 13 0 1 9 1 9 10 2
13 3 13 3 0 16 1 9 9 0 9 0 13 2
16 3 1 15 9 9 13 13 9 13 1 9 7 9 9 0 2
11 13 7 7 3 15 9 1 9 0 9 2
32 13 4 3 1 0 9 16 0 9 13 2 13 9 10 2 13 7 15 13 1 15 2 7 15 13 1 15 1 9 10 9 2
23 15 0 0 13 16 15 15 13 1 15 2 13 9 15 2 1 13 1 9 9 13 9 2
35 3 2 1 9 13 9 10 9 0 13 2 16 1 0 13 2 0 13 16 0 9 13 2 13 10 9 2 13 1 9 9 15 15 9 2
26 9 3 15 1 9 9 9 13 2 15 9 1 9 13 2 16 7 9 9 0 13 13 1 9 13 2
22 15 3 9 13 9 13 13 1 15 15 13 2 13 9 9 9 16 15 13 9 13 2
30 16 3 15 13 0 9 9 13 1 15 9 1 15 16 13 9 13 2 13 13 3 9 1 15 9 13 9 13 13 2
5 15 7 9 13 2
41 9 3 10 2 1 9 0 2 15 13 1 9 2 15 3 15 13 1 9 0 2 15 13 2 16 15 13 9 1 9 2 16 13 1 15 15 1 0 13 4 2
31 16 3 1 9 0 15 13 1 9 2 13 13 15 10 1 13 9 13 2 0 13 16 15 1 15 9 13 15 9 13 2
23 7 1 13 2 13 15 9 13 2 13 9 15 9 15 9 13 2 13 15 2 13 9 2
33 16 7 1 9 15 13 1 9 2 15 9 13 13 1 13 9 13 2 3 13 0 16 9 1 9 15 9 13 9 0 9 13 2
19 16 7 1 9 15 13 1 9 2 1 13 9 13 13 2 15 9 13 2
24 9 3 13 16 1 9 0 9 13 2 1 15 13 15 1 9 13 2 13 1 13 9 13 2
16 13 3 9 9 13 9 9 15 13 9 15 3 13 10 9 2
20 4 3 9 13 13 15 9 16 13 9 2 1 9 0 9 13 15 15 13 2
25 16 7 15 15 0 1 9 0 13 2 13 15 13 9 2 13 1 9 0 13 9 15 0 13 2
15 7 16 15 9 13 9 2 0 13 3 13 9 15 9 2
13 7 1 3 13 13 1 0 2 13 16 13 3 2
15 13 3 9 10 13 9 9 1 13 9 3 13 15 9 2
7 15 7 13 9 9 13 2
20 13 3 9 10 2 1 9 15 0 15 1 9 13 2 13 1 13 9 13 2
10 13 7 1 15 13 1 15 0 9 2
32 13 3 16 13 12 9 2 16 13 9 2 1 15 7 1 15 13 0 1 9 9 0 2 15 13 0 1 15 7 1 15 2
20 13 3 16 13 15 3 13 1 15 3 9 2 13 15 1 15 7 1 15 2
45 7 9 13 15 9 10 13 4 13 2 16 13 4 2 3 13 15 9 0 7 0 2 1 9 13 3 13 9 9 2 7 0 7 0 2 1 13 2 16 13 3 2 13 0 2
14 9 3 10 13 4 13 9 15 9 13 12 1 10 2
7 15 7 13 9 9 13 2
9 4 3 9 10 13 13 9 13 2
10 16 7 13 13 2 9 15 0 13 2
24 1 3 13 2 16 3 2 13 0 2 13 16 9 13 13 9 15 0 2 3 9 7 9 2
22 9 7 9 7 9 15 0 2 15 9 0 1 9 13 2 13 1 15 9 7 9 2
14 13 3 3 0 9 9 13 2 15 13 0 7 0 2
20 3 13 3 0 16 1 15 16 13 9 9 0 1 9 2 13 9 9 13 2
2 3 2
34 3 13 15 9 9 15 1 9 3 13 13 1 15 9 2 1 15 15 13 1 9 1 15 9 2 16 15 1 9 13 1 15 9 2
26 3 3 13 15 9 9 2 7 9 13 2 16 13 9 13 0 1 9 7 0 2 16 15 0 13 2
34 9 7 9 7 9 9 0 3 13 13 1 9 1 15 0 9 2 16 9 2 1 0 2 13 9 9 13 2 15 4 1 9 13 2
16 13 3 3 0 9 13 9 13 2 15 15 9 13 1 9 2
14 3 3 1 15 16 15 9 13 2 9 13 13 13 2
2 3 2
40 16 9 9 13 13 13 15 9 1 9 9 7 9 15 0 2 3 13 13 16 13 15 9 1 9 16 13 16 9 15 0 13 15 9 13 2 16 0 13 2
16 13 3 16 3 13 15 9 16 3 1 9 9 16 13 9 2
11 15 7 13 9 0 2 9 3 7 9 2
16 3 3 1 15 9 1 9 13 15 13 13 16 13 9 15 2
13 13 7 9 2 3 1 15 13 9 16 1 9 2
12 3 13 3 13 9 13 1 9 9 15 0 2
2 0 2
13 0 13 9 9 13 1 0 16 12 0 1 15 2
13 7 13 9 12 0 3 13 1 13 9 15 0 2
20 0 3 13 2 1 15 16 13 9 0 2 15 9 13 13 1 13 9 9 2
18 0 3 8 1 15 16 13 15 9 0 9 2 13 13 9 9 13 2
2 3 2
30 16 3 13 16 9 13 9 13 2 1 15 9 13 9 0 2 15 9 9 9 13 1 0 3 13 1 13 9 15 2
22 3 1 9 13 9 7 9 9 15 13 1 9 7 9 2 7 16 9 13 9 9 2
20 9 7 9 2 1 9 3 13 13 1 9 15 13 2 16 13 9 12 9 2
10 3 7 3 15 13 9 13 1 0 2
16 9 7 9 2 15 3 3 13 13 16 16 9 13 9 9 2
9 3 3 1 9 15 9 9 13 2
7 9 7 9 13 9 15 2
8 15 7 1 13 13 3 13 2
18 3 9 9 13 13 9 0 10 15 9 13 2 16 9 0 9 0 2
15 3 13 3 0 16 1 0 9 13 13 1 13 9 13 2
2 3 2
17 10 0 1 15 9 13 1 9 7 9 2 1 15 9 0 13 2
29 16 3 1 15 16 13 9 7 9 15 0 2 13 1 13 9 13 2 13 16 13 9 13 13 1 15 9 0 2
5 15 7 3 13 2
20 3 13 3 15 0 9 15 13 1 15 9 13 15 13 2 7 0 16 13 2
18 3 13 3 0 16 1 15 16 13 9 0 2 13 1 13 9 13 2
36 16 7 13 16 13 0 13 15 15 0 9 16 3 3 4 13 2 15 15 13 2 16 3 13 0 1 15 9 15 13 1 13 9 13 13 2
27 10 3 0 9 15 9 13 1 9 0 0 1 15 13 2 15 9 1 0 13 2 16 13 1 9 0 2
17 0 7 3 13 13 1 9 9 0 2 16 1 0 9 4 13 2
16 3 13 3 0 15 9 13 1 15 1 13 9 13 13 13 2
13 16 3 13 1 15 9 13 9 13 16 13 9 2
51 16 0 9 13 16 9 0 13 0 7 0 2 3 15 9 9 0 13 9 9 2 16 1 0 13 4 2 3 13 7 0 16 15 9 1 0 13 2 13 16 9 0 10 3 13 13 1 13 9 13 2
15 13 3 16 15 2 1 9 0 9 2 13 9 13 13 2
7 15 3 13 13 15 9 2
26 15 16 13 1 9 1 10 9 2 7 1 0 9 10 9 2 13 9 10 0 2 7 9 7 9 2
12 16 3 9 9 13 2 3 9 9 9 9 2
14 3 9 2 1 13 1 15 9 2 13 1 15 13 2
24 9 7 0 2 15 15 13 15 16 9 0 13 1 9 13 13 1 9 0 2 9 13 0 2
18 12 16 13 13 1 9 4 13 1 9 2 15 13 1 9 9 13 2
7 0 13 13 13 1 9 2
10 15 3 12 9 13 13 1 9 0 2
15 16 3 13 9 9 1 9 2 13 1 15 15 13 9 2
14 3 7 13 1 9 10 9 2 16 0 9 13 13 2
22 7 3 0 13 16 3 10 9 13 2 16 13 9 2 16 15 9 13 1 0 13 2
40 13 3 3 15 9 9 1 9 2 1 15 16 10 13 1 9 13 1 9 2 15 13 9 0 9 2 7 1 15 16 13 10 0 2 7 13 7 3 13 2
49 1 7 9 0 3 13 13 9 13 2 1 15 9 2 16 3 13 4 2 13 16 13 1 9 1 9 9 13 2 16 9 13 2 15 1 15 13 9 13 2 13 9 9 1 9 7 15 15 2
12 3 16 1 15 13 16 3 13 1 9 0 2
36 7 2 1 1 9 9 13 13 13 10 13 1 9 15 13 0 9 2 7 13 9 13 2 1 9 15 13 9 13 2 7 10 0 3 13 2
63 7 1 15 2 1 15 9 15 13 1 9 2 13 1 9 9 13 2 3 16 7 15 9 7 13 1 15 13 0 15 1 13 9 13 2 16 13 1 9 0 2 16 13 9 0 2 7 16 9 0 13 15 9 1 15 1 15 9 15 13 9 13 2
11 7 15 13 0 1 15 13 15 12 9 2
30 3 2 16 9 1 9 13 9 1 3 9 0 1 15 13 1 9 13 2 13 15 9 13 15 9 2 16 13 4 2
16 7 13 15 9 13 2 1 15 13 9 13 16 13 1 0 2
28 7 3 2 16 1 9 0 3 13 9 0 0 2 16 0 13 9 2 1 15 3 9 13 1 0 9 13 2
12 7 15 13 0 1 15 13 0 9 1 0 2
20 0 7 13 1 15 16 2 1 0 9 2 13 9 13 13 9 16 13 15 2
10 1 0 15 0 9 2 13 1 13 2
16 3 1 15 16 15 13 16 9 2 13 15 7 15 9 13 2
5 15 7 0 13 2
17 9 3 1 9 2 16 9 0 2 13 1 9 13 0 7 0 2
13 0 7 3 13 13 9 0 7 0 2 1 15 2
30 1 15 3 13 9 0 2 15 13 15 16 9 2 13 0 7 0 2 9 0 13 2 15 13 0 2 13 9 13 2
26 1 3 9 13 2 1 9 2 13 13 15 9 13 0 2 0 13 16 9 13 13 9 9 1 9 2
2 3 2
16 9 9 2 16 13 9 2 13 0 2 16 9 9 13 0 2
18 3 3 13 15 9 2 1 15 13 2 16 0 16 7 9 16 0 2
20 16 3 3 13 9 13 13 0 1 9 1 9 2 0 13 16 13 9 15 2
2 3 2
5 13 15 0 13 2
16 12 9 2 16 13 9 2 15 13 9 1 15 13 15 9 2
15 3 7 15 9 13 13 2 7 15 13 9 13 13 10 2
7 15 9 2 16 9 0 2
27 15 3 13 13 2 3 16 15 13 2 7 16 9 0 1 15 13 1 9 2 16 9 0 1 9 9 2
13 0 9 2 16 0 1 15 9 13 1 9 15 2
18 16 3 9 3 1 9 13 13 9 13 2 13 15 9 13 15 13 2
24 3 7 13 15 9 0 2 16 3 13 9 16 13 9 13 7 9 0 2 7 9 1 9 2
20 7 3 0 9 2 16 13 1 9 0 13 9 0 15 15 9 0 13 9 2
17 3 7 13 9 16 9 0 2 7 9 1 9 2 13 9 13 2
19 3 3 13 13 16 3 13 9 13 1 9 13 16 13 15 1 9 0 2
17 16 7 16 1 9 0 2 13 16 15 13 9 13 13 13 9 2
18 15 7 13 3 13 16 1 9 9 13 7 9 9 13 12 1 9 2
19 0 3 13 2 16 13 12 9 1 9 0 2 16 9 12 13 9 15 2
10 13 3 9 13 12 1 9 1 9 2
17 3 7 1 9 0 2 16 3 3 13 9 13 9 2 7 9 2
12 3 3 1 9 7 9 13 12 1 9 0 2
13 13 3 16 9 13 13 1 9 12 1 9 0 2
20 13 3 7 9 0 2 7 9 15 2 7 3 15 9 13 2 16 9 13 2
13 3 3 1 9 9 13 13 16 9 13 9 13 2
2 0 2
28 16 9 13 3 13 9 15 9 2 3 16 1 15 13 13 2 15 9 13 13 9 15 9 1 15 0 13 2
15 13 3 16 12 9 3 1 9 13 13 16 1 9 10 2
20 15 7 13 3 16 15 13 9 13 13 13 13 1 15 2 16 3 13 4 2
7 13 3 15 13 12 13 2
4 15 13 0 2
7 9 3 10 0 3 13 2
30 0 3 16 2 16 13 9 15 9 2 13 16 13 10 9 2 7 3 1 9 10 9 2 3 7 1 9 9 9 2
21 1 3 13 9 9 2 13 9 7 9 13 3 2 3 3 16 13 1 9 9 2
37 0 7 2 1 13 9 9 1 9 2 13 15 9 2 15 13 13 2 1 10 9 2 3 7 1 9 15 13 9 13 2 16 3 13 9 13 2
16 3 1 9 9 1 9 3 13 13 16 9 3 13 9 13 2
13 0 2 16 15 9 13 9 9 15 13 9 15 2
22 16 3 13 9 13 13 9 9 9 1 9 2 13 16 9 1 9 13 3 9 13 2
5 15 9 3 13 2
18 13 3 16 13 9 13 13 1 9 0 2 15 1 9 1 9 13 2
34 0 2 16 15 15 13 13 2 13 9 16 1 0 2 1 10 9 9 13 1 9 13 2 15 13 9 10 7 3 7 1 0 9 2
27 16 3 1 9 9 13 3 9 9 2 13 3 16 9 13 13 15 15 13 7 3 2 7 1 0 9 2
20 13 7 9 13 3 13 15 1 9 9 1 9 13 2 7 1 0 7 3 2
10 3 15 13 4 15 1 15 9 13 2
12 3 13 3 9 9 9 1 9 13 9 13 2
13 16 3 13 1 15 9 13 9 13 16 13 9 2
53 16 0 0 9 13 1 9 9 1 15 16 13 9 0 1 9 0 0 2 9 0 9 15 13 13 1 13 16 3 13 9 13 2 1 15 16 13 9 0 0 2 7 1 15 1 9 13 2 16 7 9 13 2
31 13 3 0 2 16 0 13 13 16 9 13 15 13 1 9 0 13 1 15 7 16 13 1 9 2 7 16 9 1 9 2
27 9 3 1 9 2 15 13 2 3 0 13 15 9 15 13 13 2 7 3 15 15 13 13 13 1 9 2
8 15 3 13 1 10 9 13 2
27 15 7 15 13 13 13 1 9 3 0 13 9 1 9 16 13 2 16 0 13 13 13 1 9 16 13 2
23 13 7 15 1 15 13 13 1 9 0 2 3 1 9 7 1 10 9 2 16 0 0 2
32 15 7 13 13 9 3 13 1 9 1 9 2 1 15 13 13 1 9 15 15 13 1 9 2 7 3 13 9 9 1 9 2
15 3 7 9 15 0 1 9 2 1 12 9 2 9 13 2
10 13 7 13 1 9 1 0 9 13 2
14 1 15 7 13 13 1 9 15 2 15 1 9 13 2
24 13 3 15 13 13 1 9 13 9 7 9 1 9 2 3 1 0 9 2 7 15 9 13 2
23 12 7 9 3 13 12 16 12 15 13 1 15 16 9 1 9 2 7 16 9 1 9 2
24 13 3 16 9 13 13 1 0 9 9 1 9 7 16 9 1 9 2 7 16 9 1 9 2
8 15 3 15 13 13 3 13 2
28 9 0 2 1 13 2 1 15 9 2 15 9 13 2 13 9 13 7 15 9 13 2 7 3 0 13 0 2
5 13 3 9 15 2
10 3 15 9 3 13 13 1 9 15 2
5 3 7 15 9 2
38 7 9 9 2 1 15 9 7 9 13 9 2 7 1 9 0 13 9 3 0 2 16 9 13 2 7 3 1 13 9 7 9 2 16 15 0 13 2
18 16 9 13 1 0 9 7 9 2 13 7 1 9 2 7 15 3 2
22 3 3 13 9 9 1 15 9 2 7 3 3 13 13 16 9 9 13 1 15 9 2
20 7 0 13 0 2 7 3 13 2 3 3 9 0 2 7 1 9 13 9 2
8 3 2 0 9 0 13 9 2
5 3 13 0 9 2
32 0 7 9 13 9 2 15 13 9 9 2 16 2 16 9 13 1 9 1 0 8 2 15 9 13 9 9 13 9 3 13 2
38 1 15 7 9 9 2 16 9 15 13 2 13 13 16 13 9 7 9 3 13 1 9 2 7 1 9 2 3 3 9 13 1 9 2 7 1 0 2
14 1 15 7 16 13 2 3 13 16 13 15 16 9 2
36 9 3 0 9 2 16 3 13 0 0 9 9 2 13 3 0 3 1 9 9 2 13 3 0 10 9 2 16 3 13 1 9 1 15 9 2
32 1 0 13 16 9 13 13 15 2 16 13 1 9 7 0 2 3 16 1 9 7 9 2 7 1 9 9 2 16 13 4 2
13 15 3 9 13 9 15 2 15 1 9 9 13 2
13 0 7 9 13 9 0 2 16 9 13 9 9 2
38 0 3 2 16 9 1 9 7 9 0 13 2 13 9 0 0 0 2 1 9 7 9 2 7 9 9 2 7 9 0 2 13 9 9 1 9 0 2
37 15 0 0 1 9 7 9 0 13 2 13 15 9 9 2 1 0 9 13 2 1 13 7 9 2 15 9 1 9 0 13 2 16 1 13 4 2
31 3 1 15 2 1 0 9 9 9 13 1 9 0 9 2 7 1 15 2 1 0 9 9 3 13 9 7 9 1 9 2
30 16 7 9 9 13 1 9 9 15 13 1 9 9 2 15 13 13 0 9 15 2 3 9 15 9 13 1 9 9 2
17 1 0 15 2 15 13 0 13 9 1 0 9 2 13 15 13 2
10 0 2 3 13 13 1 9 7 9 2
18 0 9 2 13 9 9 7 9 0 2 0 9 2 13 3 9 9 2
24 7 1 15 13 3 13 13 15 16 3 13 0 16 9 7 16 9 0 2 3 16 13 9 2
27 1 0 3 13 16 9 2 16 13 1 9 1 15 9 2 9 3 13 2 9 7 9 13 1 9 9 2
10 7 13 16 10 9 9 13 9 9 2
24 15 3 13 2 16 15 13 0 9 13 1 9 9 2 9 0 13 9 9 2 7 3 9 2
15 9 7 1 9 0 3 13 9 3 2 7 9 7 9 2
10 13 16 9 13 13 1 9 7 9 2
18 3 2 15 3 13 9 2 7 13 9 3 2 13 9 0 7 0 2
12 13 3 1 9 9 2 16 13 9 15 9 2
14 7 3 13 9 1 15 15 2 7 1 15 9 15 2
31 16 1 15 15 2 0 13 16 9 15 13 9 2 16 13 9 15 9 1 9 3 2 16 9 2 16 9 2 13 9 2
29 16 7 13 9 1 15 9 15 2 15 9 2 13 13 9 2 7 15 9 15 0 13 9 2 13 13 0 13 2
29 3 7 13 15 2 16 9 15 13 1 13 9 7 0 13 9 15 1 10 9 0 2 13 9 16 13 9 0 2
15 13 3 9 9 0 2 1 0 9 0 2 1 9 0 2
16 9 3 0 13 9 0 2 3 7 15 13 1 9 7 9 2
47 16 3 9 0 13 13 1 9 7 9 2 9 9 13 1 15 16 0 2 7 3 3 13 16 0 2 16 13 1 9 0 2 15 13 9 9 1 9 0 2 9 3 13 9 9 9 2
20 13 3 16 9 0 2 7 10 0 9 13 9 0 2 13 9 9 7 9 2
34 13 7 15 9 0 1 9 0 2 1 9 0 9 0 2 16 13 1 9 13 2 3 9 0 13 9 0 2 9 7 13 9 0 2
19 3 15 9 1 9 0 13 2 3 13 16 9 13 13 1 9 7 9 2
29 1 0 13 16 9 13 9 13 9 2 7 9 2 3 9 2 16 13 9 1 9 9 13 2 13 15 9 13 2
24 16 15 7 13 9 0 2 3 13 9 1 15 0 9 2 7 13 9 13 1 9 1 9 2
43 3 1 9 13 2 9 13 16 1 15 15 13 13 1 9 7 9 2 15 13 15 9 16 13 1 9 1 9 2 15 0 3 13 9 2 10 0 13 16 0 9 15 2
38 15 7 9 13 1 15 0 13 2 13 16 13 9 2 16 3 15 9 2 7 15 3 13 2 13 15 9 2 16 13 9 2 12 8 1 8 8 2
25 1 9 0 0 13 9 1 9 7 9 2 3 3 1 9 7 9 2 7 1 9 7 9 13 2
37 3 15 1 15 13 9 2 3 13 13 7 13 16 1 15 2 15 0 3 13 2 16 9 7 9 0 2 13 13 7 13 1 9 7 9 9 2
19 15 3 3 13 0 3 0 1 15 2 7 1 15 0 15 13 9 3 2
11 9 7 1 15 13 9 2 15 13 9 2
27 3 9 1 15 13 13 1 9 2 16 13 9 2 1 15 7 13 1 15 9 2 16 13 9 1 15 2
9 0 13 7 16 9 13 1 15 2
9 3 0 13 16 9 0 13 13 2
21 13 3 16 9 13 1 9 7 9 13 2 16 15 13 2 3 13 13 15 0 2
27 16 16 3 13 13 1 9 7 9 2 7 13 9 0 2 0 13 16 0 13 1 15 13 9 1 9 2
27 3 3 13 13 16 15 9 13 13 16 12 12 9 2 16 16 13 9 13 2 3 13 13 16 12 3 2
14 15 3 13 2 16 3 9 13 13 1 9 7 9 2
41 16 3 9 15 13 1 9 15 2 0 13 16 7 9 13 9 9 9 2 16 3 9 13 0 1 9 1 0 9 2 7 3 13 3 9 1 9 7 9 0 2
7 7 9 13 9 9 9 2
10 0 2 3 0 9 13 9 16 9 2
16 0 2 3 1 9 15 9 13 9 0 2 13 15 15 9 2
11 0 2 3 13 1 15 15 15 9 0 2
12 0 2 15 13 13 9 15 0 9 13 9 2
10 13 16 0 9 3 13 9 16 9 2
7 3 3 13 9 16 9 2
21 3 2 10 9 13 1 9 9 15 13 9 2 3 3 13 9 1 9 7 9 2
22 16 3 9 13 9 16 9 2 1 10 9 13 13 9 2 13 16 9 13 13 9 2
8 3 3 9 13 9 16 9 2
25 3 2 15 9 0 13 9 15 9 2 13 9 0 7 0 2 16 13 13 1 13 1 9 13 2
35 7 9 9 13 3 13 1 9 0 7 0 2 7 3 0 7 0 2 3 9 3 13 0 0 7 0 2 7 0 3 2 16 7 9 2
8 3 7 9 9 13 9 9 2
22 3 2 15 15 1 15 13 9 2 3 13 9 16 9 2 16 9 13 15 15 13 2
12 7 3 15 9 9 3 13 15 9 1 15 2
7 3 3 13 9 16 9 2
22 7 9 1 15 13 13 9 2 3 3 1 9 15 2 7 1 9 10 13 9 9 2
13 3 1 9 7 9 3 13 12 0 2 7 0 2
9 9 3 3 13 13 1 0 9 2
9 3 0 9 3 13 9 16 9 2
16 7 1 2 1 9 2 1 12 8 2 9 13 1 9 9 2
7 0 3 9 13 9 9 2
20 13 13 16 0 13 13 16 9 2 15 13 0 9 9 2 13 0 9 9 2
32 15 3 15 0 15 13 2 13 9 15 15 9 13 2 16 15 0 13 9 2 13 9 2 7 15 0 13 9 2 13 9 2
10 3 9 13 9 9 2 7 9 9 2
18 15 3 9 15 0 13 2 7 13 9 7 9 0 2 13 9 9 2
36 16 15 7 13 13 9 0 3 13 9 9 2 13 16 13 9 15 15 9 15 13 13 2 13 15 9 9 2 13 3 15 15 13 15 13 2
21 0 16 2 1 9 13 15 9 1 9 15 9 13 12 2 13 1 9 7 9 2
14 16 9 3 13 9 15 2 13 16 13 1 9 15 2
20 13 3 0 9 15 9 13 2 16 15 9 13 2 16 9 0 13 9 15 2
15 3 3 1 15 9 9 13 16 0 9 13 9 16 9 2
8 13 7 15 9 1 0 9 2
10 13 3 16 0 9 13 0 9 9 2
30 7 13 13 16 2 3 9 13 0 2 3 3 13 9 0 2 7 0 15 13 2 7 3 10 9 7 9 13 15 2
16 3 13 16 9 13 9 13 15 9 15 3 13 1 9 0 2
33 7 3 3 13 1 9 9 2 3 3 13 9 9 9 0 13 2 16 9 0 0 16 9 9 2 7 9 0 0 16 9 0 2
9 9 7 0 13 0 1 9 9 2
24 13 7 13 16 2 16 15 13 9 13 1 9 7 9 2 15 9 13 13 9 13 9 9 2
33 1 3 9 13 9 2 9 0 13 9 1 9 3 2 15 9 15 15 13 1 9 7 9 13 2 13 13 15 9 1 15 15 2
29 16 7 1 15 15 13 9 2 15 15 13 9 13 9 2 7 15 15 13 9 13 0 13 2 16 1 13 4 2
15 0 9 13 16 7 3 3 13 7 3 3 0 9 13 13
24 0 13 13 0 13 9 13 3 16 15 15 9 9 13 13 3 13 0 16 0 11 0 9 13
15 1 15 9 3 9 15 15 13 13 13 16 1 9 15 13
7 1 0 9 9 1 9 13
7 16 15 13 1 9 0 13
28 11 13 9 13 1 9 1 9 9 7 9 9 1 9 9 13 15 3 3 1 9 9 13 15 9 13 1 9
16 9 16 15 15 7 1 15 13 3 13 9 1 11 13 13 9
4 0 9 13 11
25 13 3 9 0 16 3 9 1 9 9 13 15 1 9 15 13 13 0 0 3 9 7 0 9 13
22 3 9 3 12 9 13 16 1 0 9 9 7 15 0 3 3 0 7 0 12 9 13
29 13 16 3 9 11 13 3 13 9 3 9 9 13 3 7 13 16 16 9 13 9 3 1 0 11 9 9 13 13
20 0 9 9 0 7 15 9 9 0 9 13 13 3 16 0 13 3 13 13 15
8 3 16 15 9 11 9 13 13
12 0 16 0 9 13 1 11 13 11 15 9 13
28 0 9 1 9 0 13 9 1 9 13 12 9 1 0 9 12 15 13 9 9 7 15 1 9 9 15 13 13
33 11 3 13 15 13 1 11 16 9 13 16 15 9 3 9 9 13 13 16 3 12 9 1 9 9 13 9 13 15 13 9 7 13
8 3 0 9 3 7 3 13 13
9 15 16 13 15 0 9 15 9 13
8 15 9 9 7 15 13 13 13
64 13 15 16 1 0 9 9 9 0 1 0 9 9 13 3 0 9 3 3 1 9 11 3 9 0 13 3 16 0 9 0 9 9 15 9 13 16 0 11 9 13 9 7 13 9 7 9 1 0 9 13 15 1 15 11 0 7 0 13 0 7 9 0 13
20 0 16 3 1 9 1 15 0 9 13 13 13 16 1 9 9 7 9 9 13
15 13 13 0 9 16 15 1 11 9 13 7 15 9 11 13
9 0 9 15 9 13 13 1 15 13
19 3 13 15 16 1 11 9 13 15 1 15 13 16 15 9 0 15 9 13
16 16 15 11 13 15 9 9 3 13 15 15 1 1 15 9 13
21 16 9 9 13 13 13 15 11 1 15 15 9 1 13 11 15 13 9 0 9 13
11 0 3 7 9 13 3 7 3 9 13 13
11 3 16 9 7 9 13 9 13 15 3 13
12 9 9 9 9 13 3 7 13 1 9 9 0
19 15 3 7 3 13 3 7 13 3 7 1 9 9 15 9 7 9 13 13
6 15 9 15 3 13 13
26 3 3 13 13 11 9 9 15 9 7 1 15 9 13 16 9 13 13 1 9 16 9 16 9 3 13
15 16 9 9 1 11 13 15 15 15 13 3 11 13 9 13
18 15 16 13 7 9 13 1 0 9 15 0 3 1 9 7 1 9 13
29 3 16 1 15 9 9 13 1 9 9 13 13 3 13 3 13 16 13 9 13 13 15 1 15 1 9 1 9 13
3 7 13 9
5 1 0 1 9 13
7 12 0 9 1 9 0 13
9 15 0 13 9 3 1 9 9 13
24 15 16 13 11 11 9 15 9 13 16 0 13 3 15 15 1 9 13 0 9 13 15 9 13
12 3 16 13 3 15 13 11 1 15 9 15 13
69 3 16 1 0 3 7 15 9 13 9 15 0 11 1 9 13 1 15 9 11 7 11 0 9 13 15 13 15 15 7 15 1 9 7 9 9 0 13 3 7 15 1 0 9 13 3 7 1 9 0 13 0 7 13 7 9 13 7 13 13 7 9 13 7 9 0 7 9 13
22 1 15 13 9 15 3 9 11 0 11 0 15 3 0 9 0 9 3 3 11 9 13
7 0 13 9 15 1 15 13
25 3 13 9 9 0 9 3 1 9 9 13 13 13 9 7 9 13 13 9 13 9 13 9 7 13
13 3 3 0 9 15 9 9 13 7 15 15 13 13
42 3 9 13 9 15 9 13 13 13 0 9 16 16 13 9 15 13 11 11 9 13 9 7 13 16 0 13 9 9 13 15 0 15 9 1 9 13 13 9 7 15 13
21 0 9 3 11 1 9 13 9 13 16 15 1 9 13 3 13 9 9 7 9 13
17 13 3 3 9 7 3 1 0 9 16 15 9 7 9 1 15 13
14 13 7 13 0 9 15 15 9 0 13 0 7 9 13
72 13 3 15 9 15 9 13 16 9 3 16 9 15 13 3 3 1 0 9 0 9 13 7 15 13 0 13 9 16 3 0 9 16 13 9 1 15 13 13 0 9 13 7 13 0 7 1 9 9 13 9 9 7 13 13 16 9 9 0 9 9 13 15 3 3 3 13 7 3 13 3 13
11 3 16 9 13 9 15 11 12 9 13 13
3 9 9 13
35 9 3 0 9 13 3 16 15 0 9 9 13 3 7 13 9 9 7 9 3 13 16 3 3 9 13 3 3 9 13 13 9 13 9 13
13 15 9 1 0 9 9 13 9 0 9 9 13 13
43 3 9 9 12 15 1 0 9 9 9 13 9 13 9 13 1 0 9 1 9 13 7 11 11 9 9 13 7 1 9 0 15 9 1 15 9 13 13 0 9 9 15 13
24 12 13 7 13 16 3 1 15 9 7 9 15 15 1 15 13 13 9 13 13 16 15 9 13
49 3 3 1 11 13 9 9 13 1 0 9 3 13 13 13 7 1 9 3 3 13 3 1 9 0 1 0 9 9 0 9 1 15 15 1 9 9 7 9 13 13 13 16 1 12 9 15 9 13
20 9 13 13 16 9 1 11 15 0 1 9 0 7 1 9 9 13 13 13 13
54 15 1 9 16 0 0 9 1 9 13 7 3 15 3 0 9 9 9 13 13 3 7 9 13 3 7 9 13 13 9 13 3 3 13 9 3 15 15 9 9 13 16 9 13 9 13 0 9 15 3 13 1 9 13
13 3 15 9 9 13 9 7 13 15 1 9 15 13
21 15 9 0 3 1 15 9 13 0 9 1 11 11 13 16 13 15 13 9 15 13
37 3 16 13 15 3 9 0 9 13 7 1 9 3 3 7 13 15 3 9 9 9 13 7 9 9 13 16 0 9 13 13 15 7 3 13 9 13
7 3 15 3 0 9 9 13
24 15 13 9 3 13 16 16 15 0 9 9 1 9 9 7 13 0 13 15 9 9 12 9 13
14 15 13 0 3 7 3 15 13 3 7 3 9 13 13
28 0 0 1 9 13 16 1 0 9 9 3 15 0 15 9 9 13 3 0 9 7 9 15 13 9 13 3 13
18 3 0 9 13 16 3 0 9 1 15 13 13 7 9 13 13 7 13
21 15 9 13 9 0 9 13 9 7 15 3 13 1 9 9 15 13 3 0 9 13
32 15 0 13 9 16 15 1 9 9 3 1 15 13 15 15 9 13 16 15 0 1 9 13 7 0 9 3 13 7 15 9 13
43 15 3 11 13 15 9 1 9 3 3 13 9 7 13 7 9 13 7 9 3 9 13 1 0 9 3 3 9 9 7 15 13 1 9 9 9 13 3 13 13 16 9 13
15 9 3 13 13 15 9 15 1 9 13 7 9 9 13 13
12 3 3 7 9 9 3 7 9 7 9 9 13
18 9 3 1 15 13 3 13 16 0 9 1 9 13 13 9 7 13 13
21 7 0 9 9 13 1 0 9 15 1 9 13 13 7 1 11 13 9 9 13 13
24 9 11 13 11 0 15 13 13 15 13 15 7 9 13 7 13 9 7 13 9 1 9 13 13
4 7 9 13 9
10 0 13 9 7 0 9 9 9 13 13
54 3 9 3 3 15 9 13 15 13 12 12 9 16 0 3 3 12 9 13 16 15 15 13 9 13 1 11 13 3 13 15 13 15 16 9 15 3 3 1 11 13 7 0 9 9 13 1 0 13 9 13 3 15 13
68 0 13 9 7 9 1 9 7 9 13 16 15 9 9 13 0 9 13 16 3 0 9 3 0 7 9 7 9 13 9 0 15 9 0 7 3 13 1 15 1 9 13 3 3 13 15 13 9 16 3 3 13 13 7 0 13 9 3 13 3 16 16 15 13 1 9 13 13
12 7 16 0 13 9 9 0 13 9 3 11 13
18 0 15 3 0 9 13 3 0 9 9 13 0 3 9 1 0 9 13
38 9 16 1 9 9 13 13 9 15 9 13 9 1 15 9 13 16 1 9 13 9 9 15 7 15 1 9 13 7 15 15 9 13 13 12 1 9 13
14 0 1 15 9 1 9 13 16 3 13 0 1 11 9
21 3 13 12 0 9 15 1 0 9 1 12 9 12 9 13 16 1 0 9 13 13
23 3 9 9 9 13 13 9 7 9 15 3 9 1 9 13 13 0 9 13 15 9 13 13
11 0 3 1 0 0 9 16 13 13 9 13
16 9 9 13 16 3 15 1 9 13 3 1 11 9 1 9 13
34 3 7 9 1 9 3 1 9 13 7 15 3 13 13 9 0 9 7 9 1 0 13 13 7 15 1 0 9 13 9 1 9 13 13
45 3 9 9 9 9 1 9 13 7 0 9 0 7 9 13 16 1 0 7 0 9 13 9 13 7 3 13 7 13 7 1 9 13 7 1 9 13 7 15 3 1 9 3 13 13
13 13 9 3 15 9 9 9 13 3 13 7 9 13
20 3 15 9 9 9 13 7 3 9 12 3 13 7 0 9 13 0 1 15 13
5 0 9 9 7 13
16 15 1 9 13 3 13 9 1 9 13 15 9 13 9 7 13
37 3 11 9 9 7 13 15 7 15 1 9 1 9 13 3 13 1 9 11 13 15 0 9 1 0 9 9 1 9 11 1 9 9 13 9 13 13
9 0 0 1 13 7 15 9 13 13
20 16 9 13 3 7 13 13 13 15 0 15 0 1 0 13 13 15 0 9 13
8 16 1 0 13 3 13 0 13
8 13 16 15 13 13 13 9 13
17 0 9 13 16 1 13 13 11 9 3 13 13 0 15 9 9 13
6 0 9 7 9 9 13
4 13 9 3 9
18 13 0 15 9 9 15 3 9 9 13 7 0 13 7 0 1 13 13
7 0 16 1 15 11 9 13
42 1 11 3 3 1 15 9 7 1 15 9 7 3 3 1 0 9 9 13 15 7 9 9 13 15 0 9 15 9 13 13 15 1 9 9 7 9 15 9 9 7 13
5 1 15 9 9 13
11 0 9 0 13 9 0 7 0 13 9 13
12 0 3 15 9 13 12 15 0 1 15 13 9
20 3 7 9 13 13 15 9 13 16 1 0 3 9 0 0 7 9 0 9 13
6 15 13 13 9 13 9
16 11 9 13 11 9 7 9 9 13 11 9 0 3 11 9 13
9 0 15 9 3 9 13 9 7 13
13 9 3 13 0 7 9 15 9 1 9 9 9 13
31 7 3 15 1 9 1 9 13 15 9 13 15 13 13 13 13 15 15 7 9 7 9 13 15 7 9 13 7 1 9 13
14 9 3 9 9 7 0 9 9 0 1 9 7 9 13
9 1 15 0 3 9 9 7 3 13
6 15 13 9 3 1 9
9 0 9 9 7 11 11 11 9 13
9 0 13 0 1 9 15 1 15 13
9 15 15 1 9 13 15 11 9 13
30 16 13 1 9 9 13 3 13 9 7 9 9 0 13 9 0 13 9 9 3 7 1 0 13 7 13 13 0 13 9
20 13 11 9 9 7 12 12 9 1 15 9 3 9 13 13 9 7 1 11 13
7 3 15 15 9 9 9 13
4 3 9 15 13
10 0 13 15 7 15 9 0 1 9 13
6 15 9 13 1 9 13
5 0 3 0 13 9
5 9 1 9 13 13
7 1 9 7 9 9 0 13
11 1 11 7 1 11 3 13 15 13 16 13
13 0 9 15 15 13 16 13 16 3 13 11 15 9
4 13 11 11 3
15 15 3 13 3 16 15 13 15 13 13 8 8 8 8 8
7 9 13 15 13 0 9 9
7 3 1 15 1 15 15 13
17 1 15 13 13 0 13 3 0 15 9 3 7 15 3 7 15 13
11 9 15 13 7 13 13 15 15 15 13 13
19 3 3 3 7 15 13 16 13 15 1 11 13 3 7 3 15 11 13 13
16 15 13 15 13 1 9 0 1 15 13 13 9 15 9 13 13
15 9 0 11 15 15 3 13 7 13 9 13 11 11 13 3
29 15 13 15 15 15 13 15 7 13 13 13 9 16 3 3 13 7 13 13 15 15 15 13 13 3 9 15 13 13
16 9 15 0 1 9 0 1 15 1 15 13 3 3 15 3 13
5 9 0 13 9 15
18 7 16 15 13 0 13 9 0 9 13 0 13 1 9 7 1 15 9
29 16 1 9 15 13 13 15 3 13 13 13 13 15 3 13 13 3 11 3 9 15 9 3 7 3 13 13 9 13
10 3 1 11 9 0 0 9 13 3 13
34 1 15 15 11 9 13 11 7 15 13 13 0 13 9 1 11 11 3 1 13 9 13 9 15 13 7 1 15 9 0 9 9 13 13
4 9 13 0 9
9 0 15 3 13 9 13 1 9 13
3 0 13 11
28 13 3 15 13 16 1 11 1 9 13 13 3 0 9 9 0 7 9 16 9 13 9 1 11 11 1 9 13
4 13 7 13 11
14 15 13 1 9 15 13 3 15 13 7 3 13 3 13
23 3 16 0 9 7 15 3 13 13 13 7 9 13 13 13 9 9 1 13 1 9 15 13
3 0 3 0
2 15 0
13 0 13 16 15 3 0 13 16 15 3 3 13 13
6 3 15 1 9 11 13
14 11 9 0 13 1 15 11 11 11 11 11 9 3 13
7 0 13 9 9 11 3 9
23 15 3 16 9 9 15 13 13 3 3 7 3 13 13 16 9 9 7 0 1 15 9 13
24 7 9 16 13 15 13 0 9 3 16 3 1 9 1 15 1 15 3 1 0 9 9 11 13
29 15 3 9 13 13 15 1 9 11 9 13 15 9 9 13 13 16 15 13 16 3 9 15 1 15 9 11 11 13
2 13 9
21 3 3 6 9 0 9 0 3 9 0 9 7 9 0 9 0 9 1 9 9 13
33 0 15 0 3 3 15 13 3 13 16 1 15 1 15 13 1 15 3 9 15 13 15 13 0 13 15 13 13 9 0 15 13 13
16 3 13 13 11 3 11 0 0 3 13 1 9 1 9 0 13
3 7 15 13
6 1 0 0 13 15 13
25 11 3 9 9 15 9 13 13 13 7 0 7 0 16 9 1 9 13 15 0 0 9 0 9 13
20 9 15 15 1 11 13 0 13 3 16 7 11 15 13 7 11 15 1 15 13
25 13 1 15 13 15 9 13 8 15 15 9 15 8 7 15 9 15 7 0 1 8 13 1 15 13
7 7 13 3 16 15 3 13
10 15 3 13 13 7 9 7 9 9 15
9 7 0 9 9 9 3 13 15 15
15 11 15 1 9 13 13 13 1 9 15 9 13 3 0 13
4 3 13 0 0
9 3 9 7 9 7 9 7 9 0
11 15 15 13 9 13 15 12 9 9 13 13
10 13 9 9 1 9 1 9 15 9 13
13 13 3 11 11 15 9 9 15 15 3 3 13 3
18 15 13 9 15 3 13 3 13 15 0 13 11 9 0 13 9 13 15
7 1 9 3 13 0 9 13
29 9 13 16 9 12 9 13 9 13 9 16 13 9 1 9 13 15 13 11 9 13 7 9 16 0 15 1 9 13
10 0 0 15 3 13 16 3 15 13 13
8 1 15 3 9 3 1 15 13
6 0 16 13 1 15 13
1 3
12 3 16 1 15 9 15 13 13 15 9 0 13
6 15 13 3 0 15 13
16 11 9 3 3 15 13 16 15 9 3 9 13 7 11 15 8
15 15 3 3 3 15 15 1 0 9 9 13 1 0 9 13
3 0 1 11
3 7 3 13
10 0 3 3 13 7 3 9 9 13 13
14 9 0 0 13 3 3 0 9 9 7 3 0 9 9
4 15 13 3 0
16 16 3 11 15 3 9 3 13 0 13 0 3 3 13 9 0
3 3 15 13
7 11 15 9 13 3 3 15
10 16 15 13 13 16 13 7 1 15 13
13 8 1 9 13 7 6 0 9 11 15 1 9 13
10 7 6 15 3 13 9 13 11 3 13
5 15 13 13 16 13
19 15 13 0 15 1 9 15 7 11 9 13 13 7 9 16 1 11 11 13
12 1 15 15 0 9 13 13 16 15 9 9 13
7 1 9 13 9 16 15 13
12 15 16 1 0 3 13 16 15 13 1 0 13
3 13 1 9
12 3 3 11 15 15 13 1 11 7 1 11 13
12 7 16 1 9 13 1 9 0 1 11 9 9
4 7 0 3 13
5 3 15 9 13 13
5 13 3 0 9 9
17 11 15 13 16 11 0 1 15 13 15 1 9 15 9 15 9 13
12 13 9 7 9 13 13 15 13 7 13 1 9
2 11 1
3 3 3 13
11 3 13 13 15 13 3 3 0 9 3 13
8 3 3 1 3 15 1 0 13
8 15 1 0 13 13 3 1 3
5 15 8 15 13 13
2 15 11
21 16 15 16 13 15 13 13 15 3 9 3 13 7 0 9 3 3 13 8 8 8
7 13 15 13 13 15 13 0
8 6 1 0 9 11 0 11 9
19 11 3 13 13 16 15 9 13 7 3 13 1 0 9 3 0 3 0 13
3 3 3 13
4 0 3 15 13
35 3 16 15 9 13 15 0 9 15 3 13 13 13 3 13 13 0 3 13 7 3 3 16 9 11 13 9 0 13 15 9 13 0 1 0
13 15 13 13 16 11 3 1 9 13 15 13 3 13
18 13 3 1 0 9 15 15 3 3 16 13 13 7 13 16 3 3 13
6 15 13 15 3 13 13
20 3 3 15 13 0 1 15 7 3 8 0 13 3 15 9 13 15 13 15 9
17 13 15 9 15 1 15 13 3 13 9 7 0 13 13 15 13 0
11 13 13 9 9 7 3 16 15 13 0 9
8 0 15 13 7 13 15 3 13
8 7 3 15 13 16 16 13 13
2 13 3
11 11 15 9 15 15 0 9 13 0 15 13
2 9 15
9 0 13 9 1 15 0 3 13 13
3 15 3 13
5 15 3 8 3 3
6 11 15 9 13 13 3
1 13
18 3 7 3 13 1 9 13 13 3 7 13 15 9 13 1 9 13 13
25 15 13 11 7 15 11 3 7 13 15 9 3 7 9 16 3 13 0 9 9 15 1 0 13 13
11 3 13 9 16 0 3 13 1 9 11 13
6 11 15 13 9 13 13
4 1 13 15 13
12 3 11 15 3 13 7 3 15 13 13 13 13
41 1 0 11 13 7 3 1 15 0 13 15 3 13 15 9 3 13 16 13 1 9 15 9 7 9 9 13 16 15 9 13 1 15 15 0 13 16 0 13 13 13
2 9 13
12 12 0 15 13 13 15 15 13 13 16 15 13
16 11 11 3 13 1 9 7 9 0 7 0 7 0 15 9 13
4 7 3 13 13
23 3 13 9 13 9 9 11 1 15 11 9 13 7 11 11 0 11 7 11 9 9 0 9
33 0 3 9 11 15 15 3 9 16 13 11 11 1 0 9 13 13 11 1 9 13 15 7 1 0 9 13 3 11 9 13 3 13
6 3 13 15 15 9 0
15 16 15 1 15 13 15 9 13 0 13 1 15 15 15 13
7 15 3 15 13 7 13 13
13 3 13 0 16 3 13 3 0 9 13 15 13 13
4 0 13 3 13
7 15 13 0 7 0 9 13
12 16 15 3 13 13 0 3 1 0 9 15 9
2 13 9
30 3 7 15 9 3 13 7 15 3 13 7 13 16 13 0 3 9 1 11 3 3 13 3 7 13 15 1 9 15 13
6 15 3 16 13 15 13
18 13 16 11 13 16 12 9 13 12 9 9 11 11 0 9 1 11 13
27 0 3 15 13 13 13 3 7 15 13 13 7 15 13 3 7 3 0 13 15 15 3 1 15 9 13 13
21 16 13 16 3 13 16 9 9 11 1 15 13 13 15 3 13 13 7 3 3 13
7 3 11 13 7 0 9 9
11 16 15 13 0 13 13 1 0 15 13 13
12 15 3 1 15 1 15 3 9 13 3 1 15
9 15 16 13 13 13 15 9 15 0
13 15 3 13 15 9 13 13 16 15 0 13 15 13
8 15 9 3 13 13 16 15 13
3 15 3 13
20 7 3 3 1 9 13 16 15 15 15 15 9 0 13 13 0 0 7 13 13
30 1 0 15 0 13 15 3 13 16 3 3 1 9 3 13 7 15 0 13 15 3 0 9 3 13 7 15 1 3 13
15 7 3 13 16 7 15 9 13 9 7 15 9 3 9 13
5 3 13 0 15 13
23 15 9 15 13 13 16 9 7 9 15 15 13 13 13 15 1 15 15 3 15 9 13 13
6 3 0 9 15 15 13
20 3 15 3 13 1 15 15 9 9 11 1 9 9 13 16 13 16 7 13 13
43 3 13 11 9 3 1 15 13 1 15 3 9 13 16 3 7 13 9 15 13 7 15 3 13 13 7 3 13 16 15 13 15 7 13 3 15 3 11 9 13 7 13 11
13 15 3 9 15 3 1 15 13 0 9 13 15 0
1 13
3 13 1 0
2 15 0
13 16 15 1 0 9 1 15 9 13 3 15 0 13
28 15 13 16 16 15 13 15 13 15 1 9 3 3 1 15 13 7 15 9 3 13 9 15 13 9 13 16 13
12 1 11 13 1 15 9 15 13 13 13 1 15
26 9 3 1 12 9 9 13 13 15 0 9 0 0 9 13 15 13 3 7 15 13 9 0 9 13 13
11 3 3 15 13 15 3 0 15 13 9 9
29 3 13 15 16 16 15 9 13 13 9 0 9 9 13 9 13 13 9 16 12 9 13 1 0 9 13 0 7 13
8 16 13 15 9 15 13 15 0
2 13 3
6 15 15 3 13 3 13
10 15 9 13 1 9 0 9 9 13 13
11 15 9 0 1 12 9 7 12 9 9 13
4 16 3 9 13
25 16 3 3 15 1 15 3 1 0 9 13 13 1 15 16 15 3 3 9 15 7 3 9 3 13
29 16 1 11 13 13 13 9 13 3 7 15 9 13 13 7 3 16 9 12 3 13 9 7 9 9 13 13 3 13
6 3 9 9 11 13 13
5 7 3 13 3 13
7 9 13 13 15 9 15 9
62 13 15 3 13 3 13 15 3 13 3 15 1 15 13 3 16 0 13 15 15 1 9 15 13 16 1 15 13 3 16 1 15 7 13 15 7 13 7 16 13 1 15 9 15 9 15 13 15 13 7 15 13 0 9 7 9 15 9 7 3 9 9
4 13 1 15 13
8 0 13 13 7 15 9 13 13
2 0 11
11 11 1 0 9 3 1 9 9 3 0 13
2 0 0
5 9 0 15 3 13
12 3 13 1 15 0 9 16 15 13 15 13 13
7 6 11 3 15 13 3 9
12 3 3 3 13 15 13 13 0 15 13 13 8
7 7 3 0 13 3 3 13
8 13 15 13 7 15 9 0 13
7 3 3 1 9 7 1 9
6 15 9 3 13 9 15
6 3 3 13 1 15 0
7 3 1 0 9 0 3 13
12 0 15 1 9 15 13 7 15 3 3 9 9
11 15 3 1 9 0 9 11 7 11 15 13
10 3 3 13 16 13 16 3 15 13 0
8 1 9 16 13 15 16 13 13
14 7 13 3 15 1 0 16 13 13 0 3 8 8 8
8 3 13 1 0 3 3 0 13
7 13 1 15 3 15 9 13
3 13 16 13
13 11 0 15 13 3 16 13 15 1 15 15 9 13
9 9 13 1 9 11 3 1 9 13
3 3 3 13
6 3 3 7 1 9 13
9 1 0 3 16 0 13 11 13 13
2 13 12
4 15 0 15 13
4 9 0 7 9
5 11 11 15 9 13
15 1 15 3 13 16 15 1 11 13 13 15 13 7 9 13
8 3 15 13 1 11 3 1 11
13 15 1 9 3 13 12 3 0 9 1 15 11 13
10 3 13 0 9 9 3 0 1 11 9
8 3 1 15 15 13 1 11 11
6 3 15 13 3 0 9
8 7 0 13 0 9 15 1 13
14 15 3 13 9 16 15 3 9 3 3 13 0 16 13
20 3 9 13 16 0 9 1 9 13 1 0 9 15 13 1 15 13 1 0 9
4 3 15 3 13
33 11 15 13 0 9 0 13 16 15 9 15 3 13 9 1 11 13 0 9 3 1 3 15 15 0 9 13 13 9 3 9 15 13
18 1 9 9 0 1 11 1 15 9 13 15 7 13 0 11 0 9 13
28 3 11 9 15 13 7 11 13 13 1 9 0 15 15 13 9 13 16 9 13 7 3 1 9 11 13 13 3
3 3 7 3
2 12 13
14 13 3 3 0 3 15 13 9 13 15 15 9 13 13
6 0 3 7 0 15 13
4 0 3 13 3
10 13 3 13 1 9 7 13 13 6 3
8 15 16 3 13 15 15 11 13
8 3 13 0 16 15 3 15 13
11 1 11 13 13 3 13 7 3 16 12 13
6 15 11 7 13 1 11
1 0
3 15 3 11
13 1 0 16 13 13 1 15 15 15 0 13 15 11
1 13
8 15 1 0 13 7 3 13 13
6 3 13 15 13 7 13
11 3 13 0 7 15 13 7 15 0 9 13
3 1 11 3
28 1 11 3 13 16 15 1 12 13 15 7 16 11 13 13 7 13 9 7 16 13 3 16 15 13 16 13 13
22 3 3 7 15 13 13 15 3 13 13 3 7 15 13 0 3 15 3 7 13 9 13
17 0 13 1 0 9 7 3 0 13 16 15 9 15 13 13 9 13
6 15 3 15 3 13 13
6 16 0 0 13 15 13
2 15 13
2 15 13
7 7 0 3 13 3 13 13
11 15 3 16 15 13 3 13 7 16 8 13
19 3 15 11 13 9 3 7 9 9 7 9 9 1 15 7 1 15 15 9
4 7 0 0 13
9 9 0 7 9 0 13 7 15 8
9 11 3 13 9 13 7 13 11 13
4 3 13 13 8
6 3 3 3 13 9 13
10 15 15 3 15 9 3 15 9 13 0
12 7 3 3 16 13 15 13 11 15 1 9 13
39 7 16 13 3 15 13 13 7 13 15 1 9 0 13 13 3 3 3 3 15 13 13 13 1 15 15 7 3 3 7 3 9 9 7 13 7 13 3 13
8 9 15 15 3 0 3 13 9
6 1 0 9 9 9 13
11 3 0 13 16 3 3 15 0 13 0 15
38 13 3 3 15 9 7 15 1 9 0 13 13 3 13 7 3 9 3 3 7 1 12 9 7 9 15 13 15 0 9 3 9 3 7 1 9 13 3
7 13 11 1 9 15 9 9
6 13 1 15 0 9 15
11 11 15 16 15 13 13 13 13 11 3 11
27 11 1 9 11 13 1 15 9 15 1 11 1 11 1 9 1 11 9 1 11 15 11 9 0 13 9 15
10 15 15 11 9 1 15 15 9 13 13
3 9 13 0
2 3 13
15 0 3 3 13 3 7 0 9 3 7 3 0 9 13 13
5 3 1 9 13 3
1 13
8 1 0 11 13 9 1 9 13
4 15 15 11 13
3 15 13 0
6 3 3 9 11 13 13
3 11 13 8
5 0 15 3 13 12
6 15 3 13 0 9 13
10 3 13 16 15 3 15 1 15 13 13
24 15 3 7 15 9 3 0 7 6 9 15 13 13 15 0 15 3 13 3 9 3 9 9 9
10 0 3 9 3 1 15 13 1 0 9
26 3 9 13 15 9 15 9 15 9 9 7 9 13 16 7 0 7 9 0 15 9 13 0 9 9 13
16 7 3 3 13 3 13 3 16 9 0 11 3 3 3 13 13
6 15 9 1 11 13 13
27 15 3 9 13 13 16 15 3 13 15 1 15 15 9 13 7 3 0 13 3 1 11 9 3 1 9 0
12 9 16 11 9 13 13 3 13 16 9 0 13
1 13
1 13
3 15 15 0
4 7 1 9 13
5 13 15 9 3 11
13 9 3 15 9 13 0 7 1 9 15 15 1 13
9 15 3 7 13 15 3 7 13 13
19 15 3 15 1 15 11 13 9 11 11 11 11 15 1 9 9 11 13 13
10 13 16 13 0 9 13 1 9 0 9
5 7 3 0 13 9
14 15 3 13 1 15 13 1 0 9 16 13 3 0 13
4 3 13 15 13
3 15 8 13
12 0 3 13 11 1 11 7 11 9 13 0 9
6 3 11 13 13 3 13
5 7 6 15 15 13
13 16 3 13 3 13 15 9 13 0 7 0 1 9
5 13 1 15 9 9
26 0 15 1 9 3 3 13 3 13 1 9 9 1 9 13 13 9 13 15 1 9 7 13 7 13 13
6 1 9 15 13 13 13
21 3 7 9 13 0 9 7 9 9 13 0 16 0 3 13 0 9 9 9 9 0
15 16 1 11 7 1 9 3 13 11 1 3 1 11 13 13
5 3 15 0 9 13
12 3 13 3 13 15 7 1 15 0 1 9 13
8 11 3 15 15 1 0 13 13
8 1 15 3 13 0 9 11 13
7 15 9 1 11 11 13 13
1 13
8 9 9 11 11 9 11 9 11
4 11 3 13 11
4 11 3 13 11
10 15 3 9 1 11 3 1 11 9 12
5 7 13 9 15 11
10 13 3 9 15 1 9 7 13 13 15
6 13 7 13 3 1 9
12 15 13 13 9 7 9 15 9 7 13 1 11
7 13 13 3 15 13 9 9
12 13 3 15 16 13 9 1 9 0 13 9 11
13 3 13 11 1 11 1 11 1 11 16 13 1 15
9 0 13 9 15 13 1 15 15 13
21 13 13 3 16 9 15 13 1 15 7 1 9 13 15 16 3 13 1 9 9 15
8 9 9 15 13 7 0 0 13
26 13 3 1 9 11 13 12 9 11 15 13 11 7 11 9 15 13 9 1 9 13 3 9 7 13 0
8 0 0 9 16 15 13 9 9
9 3 3 13 13 9 15 13 1 15
30 16 3 13 9 15 1 9 7 3 13 13 16 9 15 13 15 1 15 13 3 9 15 1 9 7 13 3 13 9 15
15 13 3 15 16 13 12 9 15 3 0 9 15 13 1 9
5 13 3 9 9 15
6 15 13 1 15 13 15
9 7 16 13 9 15 3 15 0 13
3 6 13 15
3 13 9 15
9 7 9 15 15 13 1 0 13 15
16 13 3 15 16 3 11 1 15 9 15 13 13 3 12 1 0
4 13 9 9 15
17 3 7 13 9 15 1 9 16 3 13 15 9 15 7 13 13 15
12 15 3 15 13 16 13 15 9 3 15 13 15
6 0 3 9 9 0 13
6 13 1 15 15 13 9
7 7 6 0 13 13 15 13
4 7 13 0 11
8 9 3 13 13 15 0 9 13
9 9 13 15 3 13 7 13 9 15
5 15 0 13 0 9
8 16 13 15 13 15 1 9 9
8 7 6 13 15 9 13 1 9
12 16 13 3 16 9 9 13 9 1 9 13 9
19 7 13 13 13 15 1 9 6 0 9 7 9 13 13 1 11 7 9 15
4 7 13 0 11
14 7 16 13 11 1 9 9 7 13 9 7 9 13 13
6 13 16 13 0 13 15
11 7 13 9 13 13 0 7 13 13 9 13
20 7 13 12 9 15 13 0 9 9 0 16 13 15 7 13 15 9 7 15 9
2 0 13
10 16 3 3 13 0 9 15 1 15 13
8 13 3 15 1 0 9 15 13
12 13 9 16 13 3 9 15 7 9 3 9 15
12 7 15 13 9 7 9 1 15 3 13 15 0
9 13 3 16 13 7 13 1 9 15
2 0 13
7 3 13 15 3 0 3 9
6 15 3 0 13 9 0
15 3 13 13 9 1 15 13 13 0 9 15 16 3 13 9
8 3 9 3 3 13 13 1 15
5 9 3 13 13 15
5 11 3 13 13 3
6 7 13 15 9 7 13
5 3 15 9 13 15
21 7 13 9 0 7 9 15 0 7 13 9 0 7 9 15 0 16 1 9 9 13
6 9 0 7 0 9 13
8 7 13 13 13 9 13 7 13
6 6 9 15 7 9 15
10 9 3 13 13 7 16 3 13 9 13
18 15 15 13 9 9 7 3 13 13 0 7 13 15 13 13 1 9 15
11 16 3 13 9 7 9 13 3 13 3 9
12 13 15 13 3 1 9 7 1 9 9 13 9
5 13 1 9 9 15
7 9 3 15 13 15 13 9
14 7 1 9 0 13 7 13 0 15 13 7 13 9 0
2 13 15
5 3 3 0 15 0
15 7 13 13 9 15 1 9 7 13 13 9 7 13 9 15
4 3 13 3 13
15 7 3 13 9 13 1 9 7 13 15 1 9 16 13 9
2 13 9
4 9 0 15 13
6 7 15 13 0 13 13
5 15 13 9 7 9
7 3 15 13 1 9 13 9
5 13 15 9 9 11
9 3 13 0 13 9 9 7 13 9
16 7 13 1 15 9 0 13 15 1 0 0 0 0 7 15 0
3 3 9 13
8 7 13 1 15 9 7 9 13
5 9 3 9 3 13
10 15 13 1 15 0 9 16 9 3 13
13 15 11 9 15 3 11 15 3 11 7 12 1 9
11 3 3 13 15 15 9 13 7 15 15 9
17 13 15 1 3 13 15 3 13 9 16 13 9 9 13 1 9 15
6 7 6 9 1 9 13
5 7 13 15 9 13
9 6 9 0 7 0 3 13 15 1
10 0 3 9 3 13 3 1 9 7 9
4 15 15 13 11
8 0 13 13 15 1 15 7 15
22 16 13 15 12 9 7 13 12 1 15 3 13 12 12 1 9 7 13 13 15 15 13
10 7 15 13 1 9 13 13 3 1 9
21 16 3 3 13 3 13 13 15 9 13 7 9 15 7 9 7 15 15 13 7 13
10 7 13 7 13 15 1 9 16 13 13
18 7 13 1 15 9 13 15 7 13 16 13 9 13 9 15 15 1 9
10 11 1 9 9 15 13 15 13 9 15
10 7 13 9 15 15 0 13 1 9 9
3 15 13 15
7 13 3 0 9 13 3 13
28 7 15 15 13 9 7 9 7 9 7 9 7 9 7 9 7 9 7 9 1 9 15 9 13 7 9 0 13
6 15 3 13 0 9 0
7 7 13 13 1 9 9 13
7 0 13 3 13 0 3 13
7 13 13 9 15 15 13 13
5 3 3 13 1 15
8 7 13 11 7 13 15 7 13
3 6 9 11
5 9 15 9 9 13
9 7 13 0 13 3 1 9 1 11
3 6 13 15
6 3 0 13 1 15 13
9 9 13 12 9 7 13 1 0 13
1 13
12 7 9 13 9 15 15 13 15 13 15 3 13
14 7 16 13 9 9 7 9 9 15 13 16 1 15 13
9 0 3 13 9 15 7 9 13 13
8 9 3 3 13 3 13 9 0
6 13 3 15 15 15 13
3 3 13 0
9 7 3 13 9 13 9 15 9 15
10 15 13 9 11 7 9 11 7 9 11
6 13 9 15 3 15 0
6 9 3 15 13 15 13
6 3 9 15 12 13 11
13 0 7 0 15 3 0 13 9 7 9 15 13 9
22 6 15 9 7 9 9 16 13 15 1 3 13 9 7 9 3 3 0 13 9 7 9
11 3 6 15 13 1 15 9 7 9 7 9
6 7 13 11 1 9 13
3 15 13 11
7 7 0 9 13 7 13 0
6 3 13 9 3 13 9
12 6 13 15 16 3 13 0 9 16 15 0 13
10 13 3 16 13 15 9 9 15 13 13
9 12 3 1 15 13 0 7 12 0
3 13 0 13
31 3 3 9 13 13 9 15 7 13 0 0 15 7 12 13 12 9 15 3 12 15 3 12 15 1 0 9 7 13 13 3
9 16 1 0 13 0 1 0 15 13
6 9 13 16 9 0 13
5 9 13 7 13 15
3 6 13 15
20 9 3 15 13 13 7 13 7 9 7 0 7 0 7 1 9 7 3 13 15
2 13 3
5 15 3 3 3 13
6 3 13 13 15 13 9
6 7 13 3 13 0 13
16 13 3 15 13 11 9 7 13 7 13 13 7 9 15 7 13
10 3 16 13 15 13 15 1 3 15 13
8 3 3 3 15 13 7 3 15
8 3 13 1 9 15 7 13 0
6 7 3 13 1 11 13
17 3 13 16 3 13 13 9 15 7 13 15 3 0 3 12 9 9
15 9 3 9 7 15 9 13 0 9 1 11 16 15 9 13
3 13 0 11
3 9 13 9
6 16 9 13 3 15 13
5 7 13 9 15 13
3 13 15 11
7 13 3 16 1 9 13 15
8 15 3 13 1 11 15 13 11
5 7 13 0 9 13
7 13 3 13 9 0 9 11
12 15 13 9 7 1 9 0 13 13 15 3 0
1 13
15 1 15 13 11 11 7 11 11 7 11 9 7 9 9 11
19 13 3 13 9 3 1 9 0 16 3 13 9 15 7 13 15 7 13 9
6 9 3 9 13 1 9
1 13
4 3 13 0 11
11 7 13 13 9 0 1 9 3 1 0 9
11 6 13 9 15 1 9 15 15 13 9 15
7 13 13 9 7 13 9 9
5 7 13 1 9 15
12 7 13 15 9 0 7 13 9 0 13 1 15
15 9 3 13 16 13 9 13 1 15 15 3 13 7 9 13
12 7 13 13 1 9 15 7 15 11 7 9 13
3 13 15 13
12 13 3 3 15 1 9 13 7 13 1 9 15
8 13 9 15 7 13 1 9 15
10 3 13 9 9 3 9 1 0 13 13
4 9 3 13 15
9 7 13 15 16 9 13 16 13 0
13 13 3 3 9 1 9 9 13 1 15 3 15 13
10 7 13 1 9 13 1 15 15 13 15
17 7 9 15 1 11 13 13 16 11 13 7 16 1 9 9 13 9
3 9 0 13
6 7 3 13 13 1 9
3 7 13 0
24 7 0 13 15 1 9 0 13 13 15 13 9 7 13 7 13 12 12 7 12 12 7 12 12
5 15 3 13 13 0
23 7 16 13 13 13 7 13 0 15 9 7 13 9 0 3 16 13 1 9 15 9 9 13
6 7 13 15 7 13 15
8 7 13 0 9 7 13 1 15
3 3 15 13
8 13 15 1 9 16 1 15 13
40 7 9 15 13 1 9 9 9 12 7 13 0 13 1 0 9 7 13 15 15 3 7 15 13 7 3 3 13 16 13 1 11 13 1 9 3 7 13 9 15
21 9 3 13 7 13 13 15 13 13 1 15 13 7 13 1 15 7 13 15 15 9
13 7 13 1 9 9 7 13 9 7 13 7 13 3
6 7 3 13 9 7 13
16 7 15 13 9 15 13 13 0 7 9 0 15 1 9 15 13
28 7 13 15 16 15 13 1 9 3 9 3 3 9 3 9 3 7 1 9 9 7 0 9 7 16 13 12 9
2 11 13
10 11 3 13 11 13 15 9 0 7 0
3 7 13 0
8 0 13 9 0 7 3 9 13
4 12 7 12 9
14 7 16 3 13 13 9 1 0 9 7 15 0 1 9
6 7 3 3 1 15 13
7 7 1 9 16 13 3 13
6 7 15 0 0 13 0
5 13 15 15 7 13
11 3 9 3 3 9 1 9 13 1 9 9
4 8 15 13 13
11 7 16 13 15 0 1 9 15 13 1 9
7 13 3 15 13 3 12 12
4 7 13 15 13
5 7 9 13 3 13
8 7 13 9 0 13 15 1 9
11 7 13 13 11 7 9 15 1 9 11 11
13 15 3 13 9 16 13 9 0 7 9 13 9 15
6 9 0 13 3 15 13
12 7 9 13 1 15 13 15 13 16 1 0 13
4 15 1 15 13
8 7 16 13 0 3 9 13 15
1 13
3 7 13 0
4 15 1 9 13
8 15 16 9 15 13 15 13 15
5 3 0 13 13 15
7 15 3 9 13 9 3 13
3 6 13 15
7 9 15 0 13 1 9 15
9 3 0 15 9 13 1 9 9 13
4 13 11 15 13
23 3 6 13 1 11 7 9 9 13 9 9 7 9 7 0 7 13 15 9 7 13 15 9
6 7 9 15 9 13 15
4 9 11 13 15
3 9 16 13
3 7 13 15
6 0 15 13 1 9 9
10 3 3 3 1 0 15 9 1 15 13
10 13 3 15 16 0 9 13 1 9 15
10 15 15 13 13 13 16 13 7 13 15
4 13 11 13 0
3 13 9 15
10 9 15 13 13 0 13 13 1 9 9
7 13 13 9 11 7 3 13
11 13 3 15 13 11 11 7 15 13 9 9
5 7 13 15 3 12
6 3 13 9 0 7 0
6 13 9 15 3 15 0
6 7 13 9 15 13 0
5 13 15 3 0 13
3 9 9 0
8 15 3 13 1 9 0 0 13
17 13 3 9 7 9 7 13 9 7 9 1 13 16 13 13 3 13
12 6 13 15 16 3 13 9 0 16 15 0 13
6 15 3 15 13 15 13
12 13 3 9 0 13 3 3 12 9 7 13 0
10 13 1 9 7 13 15 9 9 9 13
8 3 0 13 13 7 13 15 3
7 7 13 9 9 13 13 15
7 7 16 13 13 15 1 11
4 13 3 16 13
8 7 3 15 15 13 7 15 15
10 13 3 9 0 13 7 13 15 13 15
7 13 3 9 15 9 15 13
14 0 3 9 7 15 9 13 1 11 9 16 15 9 13
6 0 3 13 7 15 13
7 15 15 13 15 13 9 9
14 3 3 16 13 0 9 13 13 13 16 0 1 0 13
3 7 13 13
9 11 3 3 15 13 3 16 13 11
4 3 0 3 13
5 7 13 9 15 9
6 15 0 3 13 0 13
14 13 3 12 7 13 9 9 13 7 9 9 13 15 13
35 7 16 3 3 13 13 16 13 9 15 13 1 9 13 11 1 11 0 9 15 3 0 13 13 9 9 7 3 13 1 11 7 13 9 11
5 7 13 13 13 9
6 3 15 13 3 13 15
3 3 0 13
2 9 13
24 13 13 3 16 9 13 1 9 9 15 1 9 1 9 9 9 13 16 9 13 13 1 9 9
7 7 13 16 13 15 1 9
3 9 15 1
7 3 13 0 16 9 3 13
14 13 3 11 1 9 0 13 1 0 1 9 1 9 11
4 13 9 15 9
8 13 3 11 1 0 3 9 12
8 13 3 9 15 15 13 13 15
8 7 11 9 15 13 13 9 0
4 7 0 15 9
16 7 15 15 13 13 13 3 1 0 15 13 13 1 9 1 15
5 7 13 9 7 13
9 7 13 1 0 15 15 13 9 11
4 7 13 13 13
10 7 9 15 13 15 9 0 1 9 15
10 13 3 1 9 15 13 16 13 1 15
7 15 13 12 9 13 3 13
10 7 13 9 0 0 9 3 9 1 15
10 16 9 9 13 13 9 0 16 9 13
14 7 13 0 1 11 7 13 15 1 9 9 7 13 0
7 7 13 13 0 9 9 11
5 3 0 9 13 11
9 7 0 0 13 1 11 1 11 9
6 15 15 7 15 11 9
8 13 3 1 9 13 1 9 11
6 7 13 13 1 9 9
10 15 16 13 11 11 13 1 9 11 13
1 13
17 7 13 9 13 7 9 9 15 13 1 15 9 11 7 11 7 11
7 15 13 13 9 3 0 9
7 7 13 1 9 15 13 9
8 3 1 9 7 9 13 7 13
7 13 3 3 9 1 0 16
5 15 3 13 9 15
12 15 3 13 13 9 7 13 1 3 15 13 11
6 0 15 3 13 16 13
6 1 0 13 9 9 15
11 7 16 13 15 15 15 13 15 15 13 9
3 13 7 13
9 9 3 15 1 9 15 13 3 13
11 15 3 13 15 9 9 7 3 13 15 13
7 7 13 9 7 13 9 15
6 13 1 9 15 13 9
3 9 15 13
7 11 9 13 15 1 15 13
4 9 0 9 13
10 15 3 0 13 1 9 9 0 13 0
10 6 9 9 7 13 9 9 9 7 9
3 3 0 13
7 13 15 9 0 16 13 3
54 7 15 9 13 1 9 7 9 13 7 13 9 9 7 12 1 0 7 9 15 15 13 13 1 9 0 7 9 11 15 13 11 1 15 9 12 13 7 11 9 11 9 11 7 11 7 15 0 15 13 15 1 9 15
5 15 13 9 13 13
5 7 0 9 3 13
10 9 15 7 9 15 13 3 13 15 13
10 3 0 13 13 9 7 9 9 7 13
9 15 15 7 15 13 11 9 9 0
9 13 3 3 9 9 0 13 1 9
7 13 3 7 13 9 9 15
28 13 3 9 16 3 13 13 13 7 13 1 9 0 7 1 15 9 13 15 13 1 15 9 7 3 3 13 13
21 7 16 13 9 3 13 13 15 1 15 3 11 7 11 7 11 7 9 7 9 9
12 7 13 9 15 15 13 16 15 13 15 13 13
3 7 13 11
4 13 3 1 0
10 7 13 7 13 9 15 16 13 1 9
4 13 11 11 13
6 7 13 13 0 1 9
20 7 6 9 13 0 7 3 13 7 13 7 13 15 1 9 7 3 13 13 15
10 9 3 9 13 13 16 13 1 9 9
5 7 13 1 0 11
5 7 13 1 15 9
4 13 7 15 11
3 7 13 0
5 3 3 1 15 13
3 7 13 0
19 7 15 13 15 13 9 3 9 7 15 13 9 3 9 7 15 13 9 13
29 13 9 9 15 1 0 9 15 7 1 0 9 15 7 1 15 9 15 7 1 15 9 15 7 9 15 3 15 0
4 7 13 0 13
3 3 0 13
5 7 13 13 0 9
6 9 15 0 13 15 3
2 13 15
13 16 3 3 11 1 15 0 13 13 3 13 9 15
4 7 3 13 13
5 9 0 9 0 13
9 16 3 0 13 3 9 15 0 13
5 3 15 13 13 9
6 6 15 16 13 9 9
14 0 3 9 13 3 16 15 3 13 13 13 1 9 15
15 3 12 9 13 9 7 12 1 0 3 13 1 9 1 9
9 15 13 16 3 13 3 13 9 15
4 13 3 0 9
11 15 3 15 13 13 13 1 9 15 9 12
6 0 3 15 9 9 13
14 6 13 15 16 13 15 7 13 0 13 7 13 13 0
47 3 16 13 9 0 1 9 15 9 13 9 15 13 7 13 13 9 7 9 7 13 7 13 7 13 13 9 9 0 1 9 15 3 13 7 9 15 13 7 13 15 9 7 15 1 0 13
16 13 3 1 0 12 1 9 12 13 12 1 12 7 12 1 12
32 16 3 13 1 0 15 1 9 1 9 13 9 13 1 0 16 3 13 15 1 9 7 9 13 15 9 7 9 13 15 1 9
6 3 3 1 13 13 15
7 13 3 1 0 9 7 13
5 15 0 13 9 9
4 13 15 3 13
9 13 7 13 3 16 11 13 15 13
17 7 13 13 16 13 1 9 15 9 9 9 13 9 7 15 13 15
18 16 13 13 1 9 3 13 1 0 9 16 3 0 15 13 13 1 15
47 16 13 9 7 9 13 13 9 15 3 7 9 15 3 7 0 3 7 9 0 16 3 3 15 15 13 7 13 15 9 7 16 13 9 13 0 0 0 0 7 0 13 16 3 13 13 15
7 13 3 1 9 7 9 9
30 16 15 13 1 15 7 3 13 9 15 7 9 7 9 7 9 7 9 7 9 3 3 3 9 15 3 13 13 15 9
5 15 13 9 13 13
21 7 15 9 13 9 12 16 13 9 12 3 13 9 7 13 9 7 13 3 16 13
15 7 16 15 13 13 13 9 0 1 9 0 7 15 13 13
7 13 15 3 12 1 9 15
7 13 3 9 15 0 1 9
16 7 16 9 15 0 15 13 9 15 1 9 13 13 0 9 13
3 13 7 0
8 7 13 9 9 9 16 3 13
6 3 13 9 13 7 9
9 15 15 13 9 15 7 13 0 13
4 7 13 0 11
3 3 0 13
6 16 13 9 15 13 0
4 7 3 13 15
12 3 13 13 15 13 7 13 9 9 3 0 9
12 13 9 3 13 13 12 9 9 9 7 3 13
6 7 13 9 7 13 15
4 0 13 9 11
3 13 13 0
24 3 16 9 3 13 3 7 9 13 3 16 0 13 15 0 9 13 0 16 1 0 13 13 15
18 9 9 13 15 16 3 13 3 0 9 9 0 9 7 3 3 0 9
6 15 16 13 9 13 0
4 3 12 15 13
2 13 0
9 7 16 13 13 15 7 9 0 13
8 13 3 11 13 0 13 1 15
4 7 13 13 11
6 13 3 11 13 1 9
3 13 16 13
4 7 0 13 13
4 7 13 1 15
9 13 3 0 9 13 9 15 1 0
8 7 15 9 1 9 13 1 0
13 7 13 1 9 13 13 13 1 0 7 13 13 0
8 7 15 13 15 13 15 0 9
6 7 13 15 13 3 13
4 7 13 0 13
9 13 7 13 9 0 7 13 9 15
1 11
4 7 0 13 0
20 16 3 13 0 3 11 13 1 9 3 13 9 9 11 7 9 11 7 9 11
11 13 1 0 15 16 13 9 15 9 9 15
10 3 15 0 1 13 15 13 1 9 9
3 7 9 13
16 15 3 13 15 9 7 9 15 3 13 13 7 13 15 0 15
20 7 13 1 9 9 7 9 13 1 15 9 7 11 13 1 9 16 13 9 9
3 13 3 9
4 7 13 1 15
14 13 3 15 16 1 0 3 13 0 16 13 1 9 9
9 7 3 9 9 1 15 13 13 13
9 3 15 0 13 15 13 7 15 13
12 9 15 1 0 13 7 1 9 7 1 9 13
10 7 15 3 13 13 9 15 7 13 9
7 7 16 13 1 9 13 0
13 7 13 12 1 0 9 9 9 7 13 9 15 0
14 13 3 9 1 0 9 7 13 0 13 11 1 0 15
6 3 3 0 1 0 13
4 7 13 15 13
5 15 3 13 9 9
4 15 13 9 9
22 13 3 13 1 0 9 13 15 3 16 13 0 1 0 7 13 9 15 13 1 15 13
4 7 3 7 11
11 7 16 13 15 13 11 15 0 13 1 9
11 3 16 1 0 9 0 13 1 0 15 13
11 13 3 15 3 9 13 7 9 13 0 13
5 0 3 15 0 13
4 7 0 13 13
17 13 3 9 15 1 15 13 1 11 13 9 7 3 13 13 9 15
26 13 3 13 13 15 16 3 1 11 13 13 16 13 9 9 13 1 9 9 9 7 13 7 9 0 13
7 7 0 11 13 13 1 0
5 7 13 9 3 13
8 7 13 0 9 13 13 1 11
9 15 13 13 7 9 13 1 9 15
40 3 13 0 9 16 13 9 7 13 15 16 3 13 13 7 3 13 11 13 7 13 1 0 9 0 7 13 1 9 15 9 7 9 9 1 15 9 13 1 11
6 0 13 1 9 1 9
8 1 0 13 7 15 15 3 13
8 9 7 9 1 11 11 13 13
2 7 13
10 0 9 13 11 11 13 1 15 7 13
3 7 15 13
2 13 15
6 15 13 11 15 13 11
3 13 7 13
5 13 11 7 13 15
4 7 13 15 11
5 13 3 7 13 9
3 13 3 9
14 15 3 13 0 9 13 15 15 13 16 13 9 1 15
7 15 13 13 1 9 9 13
17 6 6 13 15 16 15 13 13 7 15 13 13 7 9 15 3 13
17 15 3 15 0 13 13 9 7 3 13 1 9 16 3 13 9 15
11 3 13 9 13 15 16 13 15 13 1 9
7 7 15 13 7 13 0 13
16 13 3 1 9 11 15 13 11 1 9 15 13 11 11 9 15
14 7 9 15 13 15 13 1 15 9 9 13 1 9 0
12 12 3 9 13 7 3 15 13 3 13 15 9
8 3 7 9 0 13 15 13 15
4 15 13 1 15
5 13 3 9 1 3
8 15 13 7 15 1 9 15 13
13 0 3 11 9 13 16 9 1 15 9 9 3 13
6 9 13 16 13 9 15
8 16 13 3 15 15 1 15 13
7 15 15 13 0 0 15 13
13 13 0 9 7 13 9 16 11 13 15 13 15 0
9 7 0 0 13 15 9 16 15 13
16 13 13 0 16 13 9 1 15 15 15 1 9 13 13 9 15
6 0 13 9 13 7 13
5 9 1 9 3 13
10 1 0 13 11 1 9 11 15 13 11
6 13 15 13 9 16 13
4 0 3 13 15
4 6 6 13 15
2 15 13
4 15 13 9 9
2 7 13
11 3 3 9 13 15 3 15 15 13 1 9
6 13 3 9 1 3 13
4 9 13 15 13
5 3 3 15 13 13
6 1 0 13 11 1 11
6 9 3 15 3 13 13
4 15 3 13 16
19 16 15 13 9 15 13 13 1 9 3 1 9 13 7 15 1 15 0 13
6 12 9 13 7 15 13
8 13 3 13 1 9 11 7 13
7 7 3 13 15 3 13 13
3 15 3 13
2 13 9
9 13 7 13 16 9 1 11 3 13
9 11 3 13 15 3 9 13 1 9
2 15 9
5 13 11 7 13 15
4 3 13 9 15
3 15 15 13
7 0 0 13 0 13 1 15
8 9 3 3 13 1 9 1 0
7 16 9 11 13 9 11 13
11 3 7 3 1 15 0 13 7 0 15 13
7 15 13 1 9 9 9 13
10 16 15 9 15 13 9 3 13 1 0
13 13 9 15 15 13 15 15 15 13 16 9 15 13
6 13 9 3 15 13 13
2 15 3
6 7 13 7 13 7 13
5 13 3 1 9 15
4 7 13 15 13
7 0 13 9 15 16 13 9
8 12 13 16 0 16 13 3 13
5 15 3 11 9 13
2 13 9
3 9 15 13
5 13 3 15 3 11
7 0 9 9 15 13 1 9
13 3 15 9 13 16 15 13 9 15 16 3 13 15
6 0 9 3 13 9 13
10 7 15 3 13 16 3 13 1 9 15
3 13 15 9
10 13 3 11 11 7 9 15 11 7 11
7 0 13 7 1 0 13 15
8 13 3 11 15 13 11 1 9
12 7 3 3 13 16 15 13 1 9 13 15 9
2 13 0
9 9 16 13 3 3 13 13 9 15
11 11 3 3 13 1 15 3 0 13 1 9
6 11 3 13 3 9 13
10 13 3 11 7 13 1 3 1 9 13
9 13 0 16 1 9 9 15 13 0
6 0 3 13 9 15 3
5 13 11 7 13 11
5 3 9 15 13 13
4 13 11 7 13
5 15 13 0 9 9
19 13 9 15 7 13 15 9 16 3 13 9 7 13 9 7 13 7 13 15
4 7 13 15 11
10 9 3 3 9 15 7 7 9 7 9
3 9 7 9
4 15 13 15 13
9 13 3 1 3 9 13 1 15 13
3 13 15 11
6 9 3 0 15 1 13
3 13 15 11
7 7 3 13 15 7 13 15
8 9 3 1 15 13 15 13 9
4 3 13 15 9
5 13 11 7 13 15
5 13 16 15 13 15
5 7 9 15 9 13
8 3 13 15 9 3 15 13 15
6 0 13 15 16 13 3
10 7 0 13 16 3 13 9 3 7 15
14 7 16 13 0 13 9 1 9 7 1 9 7 1 9
6 1 15 13 7 13 15
11 0 7 3 13 15 7 3 0 7 13 15
4 6 6 13 15
7 3 13 9 7 13 1 9
9 0 13 13 15 16 1 15 9 13
7 9 13 15 13 15 16 13
13 3 13 16 13 15 1 9 7 16 13 15 1 0
7 9 0 7 9 15 3 13
2 11 9
5 13 15 16 15 13
12 9 3 7 9 7 9 9 13 11 7 13 15
8 3 3 15 1 9 13 9 0
8 13 15 15 13 15 13 13 15
7 3 3 15 1 9 15 13
6 7 13 11 7 13 15
14 16 1 0 9 13 9 15 9 15 13 16 3 13 9
11 7 16 0 13 3 13 1 9 7 13 15
6 7 13 1 15 7 13
1 13
6 11 3 9 3 13 15
7 15 15 15 9 13 13 11
2 13 15
9 3 13 15 7 13 1 0 15 13
9 7 1 0 9 13 15 9 1 15
12 7 0 3 13 9 7 0 15 13 13 1 15
3 7 13 11
9 13 9 1 9 7 13 3 13 15
7 11 3 13 1 9 3 13
3 13 15 11
3 13 15 11
5 13 3 15 15 9
5 13 11 7 13 15
4 13 15 11 11
2 13 15
14 3 3 3 13 1 9 7 3 1 9 12 13 9 9
12 7 13 11 7 13 9 7 13 15 7 9 3
2 13 0
5 15 13 16 13 15
7 7 13 16 0 13 9 15
8 9 3 1 9 0 13 9 11
28 7 16 13 1 9 13 3 13 11 7 11 11 7 11 11 7 11 11 7 11 11 11 7 11 11 7 11 11
6 13 13 3 1 9 9
18 7 13 13 3 1 9 9 3 13 9 0 7 13 0 9 3 13 13
4 15 0 13 13
18 3 3 1 9 15 7 1 9 15 1 9 0 13 1 9 15 7 13
17 1 0 13 13 9 15 7 13 9 15 3 3 9 15 13 1 9
5 13 1 9 0 0
11 11 3 7 11 13 1 9 1 9 9 0
8 1 9 11 11 9 13 7 13
27 9 11 7 9 11 7 9 11 9 9 15 13 9 15 11 15 15 3 13 7 13 1 9 11 13 0 13
8 15 13 1 15 15 13 13 15
7 0 3 15 15 13 9 13
22 13 3 11 9 7 11 13 16 9 13 1 9 7 9 13 7 13 15 16 1 11 13
9 3 3 13 15 13 7 13 3 13
19 9 3 15 9 11 1 11 9 15 13 9 7 13 1 9 9 0 9 15
15 13 13 3 3 9 12 9 7 9 15 13 15 13 13 13
7 7 13 7 13 1 9 15
11 7 13 9 1 9 7 13 0 1 9 0
6 13 3 15 13 15 16
11 9 9 15 13 11 15 15 13 13 1 9
5 7 3 3 13 15
10 3 13 0 15 13 9 9 7 13 9
5 9 9 7 9 13
5 7 13 0 9 9
14 13 3 11 13 11 9 15 7 15 9 1 9 12 12
17 16 3 13 15 12 9 9 13 1 9 15 16 13 9 15 9 11
9 3 13 15 15 13 3 13 3 9
8 9 3 1 15 13 9 0 13
6 13 15 9 15 13 15
5 11 3 13 0 9
5 9 11 13 9 15
15 13 3 9 0 15 1 11 13 3 13 7 13 9 15 13
6 7 16 13 13 13 11
10 3 13 15 9 3 7 9 1 9 0
3 0 13 0
9 13 7 11 16 13 7 13 15 1
13 13 3 11 9 15 7 13 1 9 0 13 0 11
36 11 3 3 13 9 7 9 1 9 9 13 1 9 9 7 13 1 15 9 1 11 1 9 16 16 15 13 0 9 9 7 9 13 13 1 11
7 13 13 1 9 15 13 0
7 7 13 11 7 13 1 9
12 7 3 1 0 13 16 13 0 13 1 9 9
6 13 3 7 13 1 9
9 7 13 0 15 15 13 11 7 11
15 7 13 0 15 9 13 7 13 9 7 9 15 13 0 11
13 13 13 3 16 9 0 13 1 11 1 15 11 9
20 7 16 13 9 15 13 0 13 12 9 15 7 9 13 9 1 0 15 0 13
6 13 3 11 1 9 13
11 16 13 11 0 15 11 7 13 1 9 13
5 15 1 9 13 15
22 1 9 13 16 3 13 9 9 9 7 1 15 9 15 13 15 7 13 9 0 13 0
13 3 13 11 9 0 13 9 0 1 15 15 13 9
7 13 3 11 13 0 9 13
7 7 13 13 3 15 1 9
23 16 3 0 9 13 0 9 3 3 15 15 13 1 9 11 11 15 15 13 15 13 13 9
11 15 7 13 13 1 0 1 9 11 7 11
10 7 6 9 9 13 7 9 13 1 9
5 13 3 15 9 13
5 3 0 13 1 15
14 13 3 9 13 3 0 9 1 9 15 1 11 13 13
6 9 3 9 13 7 13
25 7 16 13 0 9 3 11 13 15 9 9 9 0 15 9 13 11 15 13 1 9 11 11 9 0
8 11 3 13 1 15 13 13 11
32 15 3 13 11 7 9 15 0 13 7 9 9 15 1 15 9 13 13 13 7 15 9 9 13 1 15 13 1 11 16 13 15
5 13 15 0 11 0
11 13 3 0 13 16 0 9 13 15 9 0
9 13 3 9 13 13 7 13 9 9
5 13 13 3 9 9
7 9 0 13 9 13 1 15
9 7 0 13 3 13 9 16 15 13
8 13 13 3 9 3 0 1 9
5 7 0 13 9 9
44 16 13 16 15 1 15 13 13 15 9 13 9 15 15 3 13 13 15 13 1 12 13 9 7 13 1 15 1 0 15 11 7 11 9 15 13 9 15 1 9 9 15 11 11
14 11 3 7 11 13 11 13 7 13 1 15 0 9 9
10 0 9 13 15 1 11 13 7 11 9
7 7 9 1 9 11 13 13
10 15 9 13 9 13 0 15 13 1 11
4 7 13 0 9
7 7 13 15 15 1 9 13
8 13 3 9 9 9 0 11 16
11 7 13 13 13 15 7 13 13 16 13 9
10 0 15 9 13 3 3 13 15 13 11
6 11 3 7 11 13 3
11 13 13 15 13 0 0 15 1 15 13 9
34 13 7 1 12 15 9 9 13 1 0 9 9 13 13 9 7 9 9 15 13 9 16 3 13 15 7 13 16 3 3 13 1 15 15
6 15 3 9 13 15 13
5 1 0 1 9 13
23 13 3 15 16 0 9 13 3 13 7 13 7 13 3 13 1 15 9 13 13 13 1 11
11 3 3 9 13 3 13 1 9 13 11 11
3 13 3 11
7 13 15 1 11 15 11 13
9 7 13 9 0 13 9 9 12 12
31 3 3 3 0 13 15 9 1 9 13 7 3 0 9 11 9 1 9 13 7 3 13 13 9 15 15 0 11 7 9 13
9 11 3 9 9 13 13 9 13 9
18 3 3 13 13 9 0 16 15 0 13 1 15 3 13 13 9 9 0
10 16 3 13 15 1 11 13 15 13 11
22 3 7 13 9 0 3 15 16 13 9 15 7 9 15 13 1 9 11 13 9 9 9
18 0 13 16 1 15 15 15 9 13 7 0 15 15 1 13 13 9 0
6 3 3 9 13 13 9
13 7 13 1 9 11 9 15 13 1 12 13 1 15
16 15 3 3 3 13 7 3 13 1 11 0 13 1 9 9 11
5 7 15 9 13 9
24 16 3 12 9 13 0 15 1 11 13 9 16 13 15 1 9 13 15 9 7 13 15 9 13
5 7 13 1 15 11
17 1 15 3 9 13 1 9 11 13 16 13 3 13 1 11 16 13
2 7 13
18 9 9 15 13 15 16 13 9 15 7 13 0 7 13 9 1 9 15
12 13 3 15 3 1 0 9 7 13 9 15 13
2 13 15
21 0 3 9 13 13 3 15 1 9 13 1 9 13 15 7 13 9 13 7 15 9
3 13 3 11
18 7 16 0 9 13 13 15 1 11 1 0 9 13 9 13 15 15 9
1 3
7 16 9 1 15 15 1 15
6 16 7 3 13 9 13
5 9 3 13 1 0
9 3 1 11 11 1 9 15 15 13
8 9 13 13 15 9 9 15 13
19 3 1 12 9 15 15 1 12 9 13 13 7 9 7 9 7 9 7 0
10 13 16 3 9 9 13 3 13 7 9
8 16 0 3 13 3 9 13 13
12 13 0 15 0 9 13 9 0 15 13 1 0
13 7 13 15 1 9 7 15 13 15 1 9 7 9
11 3 9 9 15 13 1 11 16 1 9 13
9 7 13 7 13 15 3 3 11 9
9 1 15 13 15 9 9 7 9 0
9 7 13 3 9 13 7 13 3 9
19 3 7 13 13 13 7 9 0 15 1 9 13 13 15 13 0 7 13 9
4 13 1 0 9
10 13 15 9 16 13 15 15 1 9 13
19 13 15 1 9 9 9 1 9 9 7 1 11 11 9 9 1 9 7 9
4 9 3 3 13
13 13 9 9 15 13 7 15 13 7 15 13 13 0
9 7 9 15 3 9 13 1 9 15
16 0 13 15 13 12 9 1 9 15 15 13 1 0 12 9 0
7 15 13 3 13 1 9 0
8 15 13 9 13 15 9 13 9
7 7 3 13 13 1 9 15
7 3 7 15 13 1 9 15
11 7 13 0 9 1 11 15 3 13 9 15
10 6 13 0 16 13 7 13 1 9 15
7 3 7 0 13 3 7 0
10 15 13 13 15 13 15 1 1 9 15
9 15 13 0 13 9 7 13 9 15
14 7 13 7 13 9 9 0 1 9 9 7 0 7 0
21 7 6 9 0 7 15 13 1 0 13 9 7 13 13 15 9 7 13 13 16 13
10 7 16 13 9 0 13 9 0 9 13
13 7 9 13 13 0 7 9 13 13 0 3 9 0
14 7 13 9 0 12 9 15 13 13 13 9 7 9 13
5 1 9 11 12 12
19 9 7 9 7 9 7 9 9 7 9 7 9 7 9 9 15 1 9 9
36 7 0 9 13 7 13 13 9 7 9 13 1 9 7 13 13 1 9 7 0 9 9 13 13 7 0 9 9 13 13 7 15 9 0 13 13
5 7 0 9 9 13
6 7 9 15 3 9 13
7 7 9 0 9 3 0 12
27 7 13 15 9 0 13 1 9 13 9 7 9 1 9 15 7 9 15 13 3 9 7 9 15 3 9 9
16 7 13 1 13 1 9 9 15 13 9 7 15 15 1 0 13
16 7 13 1 9 15 3 9 0 7 16 13 15 13 13 9 15
10 0 13 9 13 9 16 13 9 9 15
8 7 13 13 9 0 1 9 13
11 7 6 9 0 0 13 9 12 7 9 12
7 7 13 9 0 1 9 13
5 7 13 1 9 9
6 7 15 13 13 1 15
17 7 13 15 9 13 1 9 7 13 9 12 0 9 7 13 3 9
4 9 3 9 13
6 0 15 13 9 3 13
14 13 9 15 7 13 16 13 9 16 13 16 13 9 9
7 0 7 0 9 15 9 9
8 7 15 9 13 13 13 1 9
16 7 13 9 9 1 9 7 9 15 7 3 13 9 1 9 15
8 7 13 13 9 0 1 12 9
27 7 9 13 13 9 7 9 7 13 9 7 9 0 7 9 13 9 0 1 9 15 0 9 7 9 9 15
7 7 0 13 9 15 13 9
7 7 9 9 1 0 13 13
6 7 13 15 13 1 9
15 7 16 13 7 13 13 16 13 1 9 9 15 15 0 13
34 9 3 10 0 13 3 13 1 9 9 9 15 13 3 3 13 13 13 7 15 13 1 0 12 13 3 12 1 0 3 12 12 13 13
6 3 3 16 13 0 13
48 15 9 1 0 9 13 16 3 15 13 3 7 3 1 9 3 13 1 9 7 3 1 0 13 7 16 1 9 7 1 0 13 3 13 0 10 9 16 13 1 9 0 10 0 15 13 0 11
37 13 3 0 9 15 1 9 11 7 13 9 9 15 7 3 13 15 3 16 13 1 9 13 15 9 9 0 9 15 13 1 9 15 1 0 9 13
4 3 3 13 9
6 7 3 13 9 13 3
8 13 3 9 3 13 13 9 0
24 3 13 15 3 3 10 9 15 13 13 9 16 13 13 15 9 9 3 3 13 0 11 13 9
41 7 3 3 13 9 0 15 15 13 3 7 3 3 7 15 9 15 9 11 13 13 7 13 1 9 9 13 3 3 0 9 15 3 13 1 9 9 13 13 1 11
3 7 15 0
19 3 15 1 0 15 1 0 1 9 15 13 15 3 3 1 9 15 1 0
15 11 3 13 9 0 1 0 9 1 15 9 13 9 9 11
25 7 3 3 13 1 11 13 1 9 15 13 11 15 13 9 1 9 11 3 13 13 13 11 1 11
13 3 3 0 13 7 3 0 13 16 3 3 9 13
10 0 13 3 9 11 15 13 3 9 11
21 13 3 9 13 1 9 15 13 11 15 13 1 0 9 1 15 3 9 11 9 13
16 15 3 16 13 1 0 9 13 1 9 0 7 13 13 3 9
14 1 0 3 9 9 13 0 1 9 3 11 7 0 0
34 13 13 3 1 9 3 9 7 9 0 1 9 11 13 13 3 9 12 7 3 3 1 10 0 9 7 9 15 15 1 13 13 1 9
16 3 3 15 1 0 15 3 13 3 13 13 3 3 15 15 13
23 0 3 9 11 15 13 9 9 3 13 3 7 3 3 15 9 11 1 3 3 13 9 13
18 3 1 11 3 0 9 0 9 13 3 13 9 0 15 3 3 13 9
4 3 13 13 15
15 6 0 9 1 9 9 0 15 13 0 13 1 9 9 11
15 13 3 1 15 0 9 3 9 3 13 13 13 0 11 9
21 3 13 1 0 9 13 9 1 0 15 13 0 15 9 13 0 13 9 1 11 0
24 15 13 1 0 9 15 13 13 13 9 15 13 13 3 1 9 12 3 1 3 13 0 13 9
44 3 3 1 9 11 9 15 13 13 1 11 1 11 13 9 1 9 7 9 15 9 11 11 15 13 11 7 3 13 9 9 11 13 1 9 11 15 13 9 0 9 15 13 11
12 3 16 13 3 13 1 9 7 1 9 0 11
28 3 13 1 0 9 9 7 3 13 9 9 0 15 15 3 3 13 15 13 0 9 7 3 0 7 3 0 9
20 0 3 13 0 9 3 16 0 9 3 13 3 3 13 9 1 9 13 9 11
28 0 3 3 15 0 13 16 9 10 7 11 1 9 7 9 1 11 15 15 3 13 0 9 13 15 1 10 0
32 3 13 15 3 1 9 15 13 1 9 1 0 9 3 13 9 0 11 15 13 1 0 9 7 1 0 9 3 3 13 0 9
26 3 3 15 3 1 9 9 3 13 13 3 7 3 1 9 13 9 7 12 15 15 9 15 15 3 13
5 3 13 15 0 9
6 3 13 15 10 0 9
28 1 15 9 16 13 13 13 1 9 9 13 3 9 10 1 11 13 3 12 9 0 9 7 13 9 13 15 9
15 11 3 16 13 13 13 3 9 16 15 15 0 13 9 13
35 3 16 13 1 0 9 7 9 3 7 3 3 1 0 9 15 3 0 13 3 13 9 15 11 9 13 15 3 1 15 9 15 13 13 13
20 6 7 13 9 1 9 7 3 13 3 9 7 1 3 9 3 13 9 1 15
23 9 3 1 3 3 13 7 1 9 0 13 3 3 7 9 3 9 13 15 13 1 1 9
27 7 3 3 9 13 15 15 13 13 13 9 3 9 7 13 1 15 7 3 13 15 3 0 3 3 9 3
3 3 13 0
12 9 3 0 13 16 1 9 9 9 0 3 13
8 3 3 13 12 9 7 13 9
21 15 9 16 13 0 9 13 16 13 9 9 7 3 1 0 9 7 3 0 9 13
5 13 1 9 3 9
19 9 3 7 9 1 9 7 9 7 9 7 0 9 3 7 13 7 13 13
4 0 9 1 11
7 3 9 0 16 13 13 3
5 0 3 9 0 13
28 9 3 0 3 0 13 0 9 1 0 1 11 13 1 9 0 9 7 15 13 15 9 13 1 0 13 1 9
7 0 3 9 9 13 9 0
13 1 15 3 16 3 13 1 9 13 9 1 11 9
8 15 3 9 0 1 11 13 13
9 13 3 0 9 7 13 9 13 9
65 13 3 9 1 9 0 15 13 1 9 13 9 1 9 1 11 7 3 13 15 9 13 9 0 13 1 11 1 9 9 7 3 15 13 1 9 15 13 13 16 9 13 0 15 1 9 13 13 15 13 1 11 15 13 1 9 9 3 13 9 10 1 15 13 9
8 7 3 13 15 9 7 15 9
25 1 0 3 15 1 9 0 15 13 1 9 13 15 7 3 3 1 9 0 9 3 9 7 9 13
5 13 16 15 15 13
12 3 3 3 3 0 9 16 3 9 13 3 13
4 3 3 9 13
10 3 0 9 15 13 1 9 3 1 3
48 7 3 13 9 9 1 11 1 9 15 13 3 13 9 1 9 13 1 15 9 0 13 1 9 9 9 7 13 9 0 13 1 15 13 9 0 9 13 7 13 13 1 9 3 9 9 3 9
3 13 3 9
7 3 13 1 9 3 9 13
22 7 3 16 13 13 13 10 9 1 9 3 13 9 9 11 1 11 13 0 1 9 0
4 3 13 1 0
33 13 3 10 9 0 0 1 9 0 15 13 1 9 7 0 9 7 0 9 3 3 3 16 3 9 13 1 9 1 11 13 1 9
6 0 1 0 12 9 13
19 13 9 3 0 1 9 13 15 1 9 15 3 3 9 0 9 9 9 0
15 16 3 3 13 13 13 15 9 1 9 0 15 13 1 9
11 3 3 1 0 15 1 11 13 13 1 11
21 7 3 3 13 1 9 15 9 3 1 12 0 1 9 9 13 7 9 0 9 10
5 3 13 3 1 9
7 1 9 3 15 3 13 13
38 16 3 13 15 9 9 3 15 9 1 0 15 13 15 13 12 9 13 9 9 0 9 0 15 13 1 9 13 3 7 3 9 1 9 7 13 9 15
10 16 3 1 15 13 13 0 3 13 13
10 3 3 13 9 3 1 9 0 1 9
11 3 0 7 0 15 13 13 9 1 11 13
29 7 3 1 0 3 13 13 16 3 3 0 9 0 13 0 9 13 15 9 9 13 13 16 3 15 9 0 9 13
12 3 0 7 0 9 1 9 0 15 13 9 13
