386 17
4 1 11 12 11
27 3 4 4 16 9 1 9 10 0 9 13 4 1 10 0 9 7 9 1 9 7 0 1 10 15 9 2
18 3 13 9 9 4 1 10 9 16 3 1 9 7 0 9 3 4 2
21 3 4 1 9 16 9 9 13 1 0 9 7 15 9 7 9 4 4 7 4 2
22 3 10 9 0 9 13 2 13 1 9 4 7 4 0 1 10 0 9 1 10 9 2
33 1 10 9 13 10 13 9 0 1 15 16 10 9 4 7 9 4 2 3 10 9 2 10 9 2 9 2 9 2 9 7 9 2
8 10 9 1 15 8 1 10 9
19 10 9 9 1 10 11 13 1 0 11 1 15 9 1 15 9 4 4 2
15 3 13 3 0 0 9 4 1 9 15 1 10 9 13 2
18 15 4 0 1 10 9 1 10 13 9 1 15 13 7 13 1 9 2
34 8 10 9 1 15 9 2 13 3 4 4 16 10 9 9 10 15 9 4 7 7 10 9 1 10 9 9 0 9 7 15 9 4 2
1 9
11 9 1 10 9 1 10 15 9 4 4 2
21 10 9 1 10 11 13 0 4 4 16 10 9 9 4 1 10 9 1 15 8 2
16 3 1 10 9 1 10 9 7 9 13 15 10 0 9 4 2
9 10 9 13 9 4 7 9 4 2
25 0 13 10 9 3 3 15 0 4 1 10 9 1 10 11 7 15 4 0 1 9 1 10 9 2
16 3 13 10 9 3 3 1 10 9 4 15 9 4 4 4 2
32 3 13 10 9 1 10 11 15 9 1 10 9 15 3 16 1 3 1 15 9 8 9 7 9 4 4 7 15 0 4 4 2
16 15 13 3 0 7 0 16 1 3 1 4 4 1 15 9 2
22 9 13 3 3 0 4 15 15 9 4 7 10 0 2 0 9 4 1 10 15 9 2
12 3 4 13 9 4 8 9 2 9 7 9 2
4 9 1 10 9
1 8
10 15 13 8 15 0 8 3 1 13 2
9 1 15 9 13 15 9 13 4 2
18 10 9 13 8 10 9 1 10 9 4 7 0 10 11 1 9 4 2
23 9 1 10 9 15 9 1 10 9 7 10 9 1 9 7 0 1 12 7 10 0 9 2
20 10 9 4 3 0 4 1 15 8 2 10 0 9 1 15 1 11 13 9 2
14 3 13 9 4 16 10 9 1 10 0 9 4 4 2
3 1 9 11
32 10 9 1 15 8 7 15 13 1 10 0 9 13 0 4 1 13 0 9 1 9 1 9 7 0 1 12 1 12 9 11 2
14 3 10 9 4 4 2 4 3 3 3 0 1 4 2
2 11 15
33 1 15 9 13 10 9 7 10 9 8 10 9 1 10 11 7 0 9 1 9 7 0 3 0 4 4 7 0 13 0 4 4 2
22 10 9 1 15 8 4 3 3 3 15 9 1 10 0 9 3 13 2 13 7 13 2
28 15 4 3 10 0 9 1 10 0 9 9 13 2 0 0 9 1 9 7 0 1 12 1 12 9 11 11 2
16 3 13 15 10 0 9 3 1 10 0 2 0 7 0 9 2
4 3 1 10 9
23 10 0 9 13 1 12 9 2 3 3 12 4 4 1 10 9 9 7 12 1 10 9 2
19 12 9 4 0 4 7 12 9 13 10 9 5 13 9 2 9 12 2 2
8 9 1 10 12 9 1 15 8
6 11 12 2 9 7 9
6 9 12 2 9 7 9
22 1 9 7 13 13 15 1 15 0 13 1 9 1 10 9 1 10 9 7 9 9 2
12 3 4 10 9 4 15 10 9 13 7 13 2
5 9 12 2 9 13
5 10 9 4 0 2
28 3 1 0 9 0 10 0 13 9 13 7 8 13 2 3 1 9 7 9 13 13 16 8 13 13 4 4 2
6 9 12 2 9 7 9
10 9 12 2 9 2 9 2 9 7 9
10 9 12 2 9 2 13 2 9 7 9
1 11
21 8 2 12 9 2 13 7 1 9 16 9 10 9 2 3 10 9 1 10 9 2
1 11
13 15 13 1 10 9 1 11 9 10 9 1 4 2
11 3 13 15 0 9 1 15 9 4 4 2
22 10 9 13 10 9 3 3 1 10 9 7 13 16 0 9 1 10 9 1 11 9 2
5 11 12 2 13 13
31 1 15 13 1 10 9 4 4 1 15 9 10 9 7 10 9 4 4 7 16 10 9 10 9 7 9 1 15 9 4 2
26 15 13 3 3 4 1 10 0 9 1 0 0 9 2 16 10 0 1 9 7 1 10 9 13 9 2
15 3 4 4 1 15 9 0 7 9 1 9 4 1 9 2
5 9 12 2 9 13
10 9 12 2 9 2 9 2 9 7 9
1 11
5 8 4 12 9 2
10 15 4 0 0 7 13 3 0 9 2
18 15 9 13 10 11 16 15 15 0 4 16 0 1 11 16 1 4 2
6 9 12 2 9 1 9
19 10 0 13 3 10 0 9 1 4 1 11 9 7 0 9 1 10 9 2
10 8 13 15 10 9 1 10 9 3 2
10 9 12 2 9 2 13 2 9 7 9
34 10 9 1 10 9 13 15 3 1 13 3 10 9 1 10 9 1 15 9 4 7 1 10 9 15 10 9 1 10 9 13 1 13 2
14 8 13 15 10 9 1 10 9 1 11 7 15 9 2
1 13
14 11 0 1 10 9 4 8 10 9 3 4 1 9 2
7 3 4 0 3 9 4 2
6 11 12 2 9 7 9
9 13 7 9 4 1 15 9 4 2
18 0 15 9 13 3 10 9 2 9 1 9 2 9 2 9 7 9 2
8 10 0 9 4 10 0 9 2
8 0 13 3 3 9 7 9 2
1 11
1 11
16 8 4 12 9 0 16 10 0 9 1 15 8 8 10 9 2
13 3 4 10 9 9 1 10 9 1 10 9 4 2
13 15 4 3 4 1 10 9 1 10 12 13 9 2
9 1 11 4 3 15 9 1 4 2
15 4 15 3 10 9 2 3 13 15 3 0 9 4 4 2
10 11 12 2 9 2 11 2 15 7 9
15 7 9 16 0 15 13 0 7 1 9 9 7 9 4 2
31 3 4 9 9 4 1 15 13 7 1 15 13 1 0 9 1 15 9 1 3 9 1 15 13 1 9 7 1 0 9 2
3 9 1 9
14 9 13 9 4 1 9 16 13 2 9 7 0 13 2
1 11
14 8 2 12 9 2 4 1 10 9 3 0 7 0 2
27 16 10 0 11 7 15 9 3 13 2 13 16 10 9 0 13 1 9 7 9 15 1 9 1 13 13 2
9 3 13 3 15 9 1 0 9 2
22 10 9 1 11 13 15 3 3 7 13 1 3 0 1 4 3 15 1 9 4 4 2
13 15 13 0 9 3 0 9 7 0 9 7 9 2
21 11 9 13 1 10 9 9 3 15 13 9 1 11 4 4 7 0 9 4 4 2
28 3 13 10 0 9 1 10 0 9 2 16 15 15 9 13 4 4 7 1 15 13 4 1 10 9 1 11 2
6 11 12 2 15 1 11
13 10 9 15 10 9 1 10 9 13 4 4 4 2
25 15 13 3 10 0 9 4 7 15 13 3 4 1 9 15 9 13 1 13 7 15 9 9 13 2
25 3 4 3 1 15 9 9 1 10 0 9 2 4 3 15 9 7 3 4 10 9 1 10 9 2
27 16 9 1 15 9 3 1 13 13 10 11 0 4 1 3 10 9 2 10 9 2 10 9 2 8 3 2
1 9
1 11
22 10 0 13 10 0 9 1 10 0 9 16 12 9 3 10 0 9 2 11 2 13 2
9 10 9 13 0 10 0 13 9 2
33 15 13 10 0 1 16 10 9 0 4 0 3 4 15 3 3 0 1 10 9 2 13 10 9 12 7 16 3 10 13 9 13 2
11 1 10 9 1 15 13 13 10 13 9 2
27 15 13 3 3 0 1 10 9 7 9 1 16 15 3 2 3 13 3 10 0 3 4 2 3 13 4 2
10 11 12 2 11 2 9 2 11 7 9
17 1 15 9 13 15 16 10 9 15 10 9 7 9 1 9 13 2
13 10 9 2 11 2 4 10 0 9 0 1 9 2
15 9 2 13 7 13 4 0 1 0 2 0 9 1 9 2
9 1 0 9 4 3 9 1 9 2
13 1 9 1 9 4 9 7 9 3 9 10 9 2
1 11
15 8 2 12 9 2 13 15 0 16 10 15 1 15 9 2
24 15 9 4 13 1 10 9 1 10 0 13 0 9 2 15 1 12 1 0 9 13 4 4 2
30 3 1 15 0 9 4 11 7 15 9 4 1 10 11 2 10 9 15 0 9 1 10 9 1 9 13 3 1 4 2
15 15 13 3 9 1 13 9 1 10 9 7 0 0 9 2
24 10 9 13 1 3 12 0 1 10 9 2 15 0 13 2 10 9 2 10 9 7 10 9 2
24 1 10 9 1 10 11 13 10 9 1 11 3 15 11 4 4 7 3 15 15 9 4 4 2
9 15 13 15 1 10 9 0 13 2
2 15 9
6 9 12 2 9 7 9
4 11 12 0 0
23 10 9 13 3 1 10 0 9 11 1 12 2 3 10 9 1 10 9 0 4 13 4 2
1 9
19 10 9 1 15 8 1 12 13 10 9 9 2 11 2 0 9 7 11 2
23 15 12 9 4 1 15 9 3 15 13 7 4 3 3 16 9 4 1 10 9 0 9 2
23 16 3 15 0 9 7 9 13 1 15 13 1 10 0 9 2 4 15 8 16 15 4 2
23 1 10 9 4 4 3 13 4 4 4 15 9 1 9 2 0 9 7 9 4 13 4 2
39 1 9 13 10 0 9 4 4 4 1 0 9 15 0 1 10 0 9 4 13 4 2 3 9 2 7 9 15 1 13 9 13 13 4 2 3 0 2 2
25 10 9 1 9 13 10 0 9 1 15 2 8 2 13 1 10 11 7 13 3 3 1 10 9 2
4 11 12 0 9
1 9
19 10 9 2 0 9 2 13 15 15 9 1 2 9 2 13 4 4 4 2
8 15 4 10 9 1 15 9 2
26 3 13 15 0 9 7 9 1 15 13 1 10 2 0 9 2 2 7 15 8 13 16 15 4 4 2
23 10 13 9 1 10 9 4 15 13 2 15 0 13 1 10 9 1 10 9 1 10 9 2
21 3 13 3 10 9 15 16 9 13 4 2 7 15 9 4 1 15 9 13 12 2
6 12 1 9 13 9 12
3 11 11 12
16 10 9 4 10 0 9 1 10 9 1 10 0 9 12 9 2
1 9
24 9 2 9 7 15 9 1 15 7 1 10 9 15 0 9 1 10 0 9 1 10 13 9 2
16 1 9 1 15 9 13 15 8 13 9 2 9 7 9 8 2
12 1 15 13 1 10 9 13 15 13 9 8 2
18 3 13 10 0 9 2 15 10 9 13 3 13 9 4 13 4 12 2
3 11 12 9
15 1 10 9 4 10 9 4 1 10 9 9 7 10 9 2
1 9
18 15 13 1 10 9 1 9 7 0 13 1 10 0 9 1 10 9 2
15 1 15 13 1 9 7 9 1 9 13 10 0 13 9 2
9 15 9 4 4 1 2 8 2 2
24 1 10 0 9 2 9 7 9 2 13 15 8 0 16 0 9 15 1 15 9 4 4 12 2
14 15 8 13 10 9 11 8 11 7 1 0 9 11 2
31 1 9 4 10 9 1 10 9 1 9 7 9 4 2 7 15 4 3 3 0 4 2 3 3 13 4 4 1 15 8 2
29 15 13 3 10 9 1 0 9 1 10 9 1 10 9 12 9 2 7 13 3 9 1 10 13 9 1 9 9 2
47 1 9 7 0 1 10 9 15 0 8 13 9 5 9 4 7 1 9 2 16 15 8 2 11 2 12 7 12 2 15 8 2 11 2 2 15 8 2 11 2 7 15 8 2 11 2 2
15 3 13 3 15 9 1 10 0 9 1 15 13 5 9 2
35 3 13 16 15 9 3 4 4 4 1 10 9 3 10 11 8 4 2 4 3 10 9 1 9 0 16 12 9 3 1 10 9 9 4 2
13 10 0 9 4 4 8 10 1 10 9 13 9 2
10 3 13 15 8 1 15 9 16 9 2
3 11 11 12
1 8
21 10 9 1 10 9 13 3 3 16 10 9 3 1 10 9 1 9 0 4 4 2
1 9
32 1 10 9 2 9 2 13 15 8 1 8 10 9 9 1 15 9 4 2 15 15 0 2 0 2 0 7 0 13 8 13 2
19 10 9 4 3 0 3 0 7 3 3 0 16 16 9 0 1 4 4 2
13 10 10 9 4 1 10 16 9 9 3 1 4 2
8 1 9 13 15 3 4 3 2
3 13 7 9
7 13 7 9 2 9 7 9
13 13 2 15 13 13 2 13 2 13 2 13 2 9
10 9 7 9 2 9 2 0 9 2 9
7 13 2 9 2 9 2 13
5 9 2 9 2 9
20 10 1 11 13 9 13 1 10 0 9 7 3 1 10 9 9 1 15 8 2
12 3 13 15 0 9 1 15 13 1 15 9 2
25 3 4 3 10 0 9 15 3 10 9 13 4 12 7 3 3 13 15 8 16 0 9 4 4 2
26 0 9 1 10 9 7 10 9 1 9 1 9 7 9 1 11 13 4 1 10 0 9 1 10 9 2
3 11 12 8
1 9
3 1 11 11
23 15 13 1 10 0 9 1 10 9 4 1 10 9 9 1 15 8 4 2 9 12 2 2
11 15 13 3 1 10 9 1 9 1 9 2
12 10 0 13 3 1 10 13 9 1 10 9 2
30 15 13 3 1 10 9 1 10 0 9 2 3 1 10 9 1 0 9 15 1 12 12 9 4 4 2 8 1 12 2
21 16 10 9 1 15 9 0 4 2 4 15 3 1 10 9 9 1 15 8 4 2
28 1 9 1 10 0 9 4 10 0 9 0 12 7 4 10 9 2 15 4 4 1 15 8 1 0 9 4 2
16 10 9 13 10 0 9 1 10 9 1 10 3 0 0 9 2
17 3 13 15 8 10 0 9 1 15 13 1 10 9 1 0 9 2
23 1 9 1 10 9 1 10 0 9 13 10 9 1 10 0 10 9 4 1 10 0 12 2
3 1 11 11
17 10 9 1 10 9 13 1 10 9 1 9 1 8 2 11 2 2
11 15 13 0 10 9 13 3 1 15 8 2
15 0 9 13 9 1 0 2 0 7 0 9 1 10 9 2
31 1 9 1 10 9 1 10 0 9 16 10 9 2 9 2 9 2 9 2 4 10 9 4 1 9 7 1 9 1 9 2
19 15 4 10 0 9 1 10 0 9 1 10 9 1 10 9 1 15 9 2
10 1 11 11 7 11 11 1 9 7 9
34 15 13 1 9 7 15 13 1 9 7 9 1 0 7 9 9 4 0 16 9 1 4 4 7 13 9 1 10 9 9 1 15 8 2
26 16 10 0 9 1 15 8 0 13 2 13 15 9 9 1 9 7 9 0 1 10 0 9 4 4 2
3 11 12 9
1 8
1 9
28 16 1 10 9 2 8 2 2 12 2 4 9 15 9 1 2 8 2 13 0 1 15 0 13 1 0 9 2
15 10 0 9 1 15 2 3 7 15 2 4 3 3 0 2
22 3 13 15 9 8 2 9 13 2 7 0 9 1 9 7 9 3 13 2 3 2 2
20 16 10 0 9 1 15 8 0 13 2 13 15 9 1 10 0 9 4 4 2
3 9 1 8
4 11 11 11 11
1 9
16 15 13 1 10 0 9 4 0 1 15 0 13 1 0 9 2
15 10 0 9 1 15 2 3 7 15 2 4 3 3 0 2
22 3 13 15 9 8 2 9 13 2 7 0 9 1 9 7 9 3 13 2 3 2 2
20 16 10 0 9 1 15 8 0 13 2 13 15 9 1 10 0 9 4 4 2
4 11 11 11 11
1 9
1 9
19 15 8 13 1 15 9 1 12 10 3 0 9 1 9 1 15 9 4 2
17 8 13 15 3 13 1 13 7 13 9 1 10 0 7 0 9 2
6 1 4 13 8 3 2
1 9
9 9 7 0 9 2 9 7 9 2
3 9 7 9
1 9
1 0
16 15 13 1 10 0 9 4 0 1 15 0 13 1 0 9 2
15 10 0 9 1 15 2 3 7 15 2 4 3 3 0 2
22 3 13 15 9 8 2 9 13 2 7 0 9 1 9 7 9 3 13 2 3 2 2
20 3 13 15 10 9 2 11 2 3 9 16 9 10 9 13 15 15 0 13 2
20 16 10 0 9 1 15 8 0 13 2 13 15 9 1 10 0 9 4 4 2
3 11 11 11
1 9
34 15 13 1 15 9 3 1 10 9 1 10 9 15 2 7 1 10 9 1 9 1 9 7 0 2 16 15 10 9 3 0 13 4 2
10 7 3 13 15 10 9 1 15 9 2
22 10 9 2 0 9 2 13 3 15 8 13 1 15 9 1 9 15 9 16 9 13 2
35 16 10 0 9 0 0 9 13 4 2 13 10 9 3 1 10 9 9 1 15 8 2 16 15 1 9 13 1 10 0 9 3 0 4 2
5 9 12 2 9 13
7 11 12 13 9 11 5 11
13 3 13 15 10 9 1 9 7 9 7 1 9 2
22 15 13 1 10 9 1 9 7 9 4 10 9 1 15 13 1 10 9 1 10 9 2
10 15 9 4 8 1 15 9 3 4 2
14 15 9 4 3 3 1 10 9 9 1 15 8 4 2
4 11 12 13 13
17 15 13 1 10 9 13 3 15 13 1 10 9 1 9 7 9 2
4 1 11 12 11
16 15 9 13 10 9 1 10 9 7 10 9 3 0 9 0 2
13 15 9 4 3 16 15 4 1 10 9 1 12 2
20 15 13 1 10 9 13 3 3 9 3 1 4 1 10 9 9 1 15 8 2
8 11 12 15 10 9 7 9 11
22 1 10 9 2 9 7 9 13 10 9 7 15 8 1 8 1 15 13 1 10 9 2
25 1 15 0 13 1 10 9 1 10 9 4 15 0 1 15 9 1 13 15 9 4 7 4 4 2
22 3 13 15 0 9 1 9 2 16 9 2 9 2 9 2 9 7 9 8 4 4 2
4 11 12 15 9
12 15 13 10 0 9 2 8 10 9 1 9 2
15 7 1 10 15 9 4 10 9 3 0 16 1 10 15 2
32 1 15 9 4 10 9 11 4 2 4 10 9 1 10 9 4 7 13 10 13 9 8 10 11 2 9 7 9 2 0 4 2
24 15 13 1 10 9 1 10 13 9 2 10 9 2 4 1 9 16 8 0 9 13 1 13 2
13 15 13 1 15 13 1 9 13 1 0 9 4 2
30 3 13 15 9 8 15 13 1 9 13 2 7 10 0 9 1 15 0 0 13 4 16 1 4 2 13 2 3 2 2
43 10 1 15 8 1 12 13 9 4 3 4 2 16 0 4 13 4 1 10 9 7 10 9 1 15 3 2 8 16 9 4 13 4 4 8 9 9 2 9 7 0 9 2
8 9 13 8 4 4 4 8 2
11 13 9 2 3 15 13 1 10 15 9 2
10 13 9 2 3 15 13 1 10 9 2
21 1 10 0 9 13 15 13 1 10 15 9 7 9 16 10 9 1 10 9 4 2
8 1 10 0 9 13 9 15 2
21 15 13 4 16 15 1 10 15 0 9 4 3 0 4 15 3 15 9 3 13 2
6 9 12 2 9 7 9
3 11 12 11
2 10 9
21 10 0 9 1 9 1 12 1 12 9 4 0 4 1 3 12 9 1 12 9 2
1 9
1 0
31 16 10 9 2 9 2 4 2 13 3 15 1 10 9 0 1 10 9 1 11 7 11 7 4 15 1 0 9 15 9 2
12 3 4 1 10 13 9 10 15 13 9 0 2
9 1 11 8 11 11 2 11 7 11
17 1 12 13 10 0 9 1 9 10 9 1 11 2 11 7 11 2
3 1 11 11
26 13 9 1 10 9 13 1 10 9 7 9 1 10 0 9 11 2 8 13 1 0 9 1 9 2 2
23 10 0 9 1 9 7 0 1 12 1 12 9 4 1 9 1 12 0 9 2 11 2 2
13 13 9 1 10 9 13 1 10 9 7 0 9 2
15 10 13 9 1 10 9 1 15 13 4 4 1 15 8 2
17 11 11 5 0 9 1 0 9 2 13 1 10 0 9 1 11 2
2 1 11
1 8
13 1 9 13 13 9 9 1 10 9 1 10 9 2
15 10 13 9 1 10 9 1 15 9 4 4 1 15 8 2
4 1 11 11 13
14 1 3 1 9 10 12 9 15 9 3 1 15 3 2
17 15 0 9 13 1 10 0 9 1 10 9 4 4 1 0 9 2
5 1 11 11 7 9
15 1 15 13 1 9 7 9 1 9 13 10 0 13 9 2
31 1 9 4 10 9 1 10 9 1 9 7 9 4 2 7 15 13 3 3 3 3 16 15 1 0 9 0 13 4 4 2
19 0 13 3 9 4 4 1 15 8 2 3 10 9 4 4 1 15 8 2
4 1 11 11 9
29 1 3 12 4 0 10 11 7 10 3 13 13 9 11 4 1 15 13 1 12 9 0 9 1 10 9 1 9 2
15 10 13 9 1 10 9 1 15 9 4 4 1 15 8 2
17 10 9 4 15 1 0 9 10 9 4 13 4 1 10 0 9 2
17 11 11 5 0 0 0 9 2 13 1 8 2 11 2 1 11 2
9 3 13 3 15 0 9 1 9 2
3 11 12 9
1 9
18 10 9 2 11 2 4 8 12 4 1 10 9 1 9 1 0 9 2
15 3 13 3 15 9 0 9 7 4 15 9 3 3 4 2
8 3 4 10 0 9 9 4 2
10 10 11 13 3 16 1 10 13 9 2
19 10 9 7 10 9 1 9 11 4 4 4 1 10 11 4 3 3 4 2
19 16 10 9 9 1 9 2 4 10 9 1 9 11 0 3 1 9 4 2
17 8 15 0 13 10 9 11 9 0 13 1 10 9 4 4 4 2
20 3 2 10 3 13 9 1 9 4 0 2 16 15 13 4 4 1 0 9 2
25 1 10 9 1 9 2 7 8 10 11 16 3 2 13 10 1 15 8 13 9 16 0 9 12 2
17 0 9 1 10 11 13 8 1 10 9 9 1 15 8 4 4 2
6 13 3 9 11 11 2
5 15 13 4 4 2
57 11 10 9 13 10 9 1 10 9 3 10 9 1 10 9 9 13 2 11 5 9 2 11 5 9 2 9 5 9 2 12 5 9 2 9 5 6 2 9 5 9 2 9 5 9 2 11 5 8 9 9 2 8 5 9 11 2
5 2 8 5 8 2
10 9 12 2 9 2 9 2 9 7 9
5 11 12 9 13 9
27 0 13 15 9 1 10 9 3 9 1 15 0 1 15 13 1 10 11 1 12 1 9 7 12 1 9 2
1 9
26 1 15 8 2 11 2 4 10 9 4 1 10 9 9 9 13 2 0 0 16 15 8 2 11 2 2
22 1 10 0 9 16 15 13 1 10 9 7 1 9 13 15 10 9 13 1 10 9 2
17 0 13 3 0 9 8 15 13 1 9 1 9 2 9 7 9 2
16 15 9 13 3 1 10 9 7 3 1 10 13 9 7 0 2
10 9 12 2 9 2 13 2 9 7 9
3 11 11 9
22 10 9 1 15 0 9 4 3 4 1 10 9 1 10 9 1 12 1 9 1 12 2
1 9
19 1 15 8 2 11 2 4 15 13 1 15 9 10 0 9 3 1 4 2
11 1 10 9 13 15 3 13 8 16 15 2
24 1 15 0 9 13 3 10 9 9 3 8 10 9 2 13 1 9 12 1 10 0 9 2 2
29 15 8 13 10 9 3 1 10 9 15 10 9 1 15 9 13 4 7 4 3 10 3 0 0 9 1 15 8 2
25 10 9 13 3 10 9 16 1 13 9 15 1 10 9 9 13 1 4 2 13 1 9 11 2 2
15 1 9 2 3 8 9 2 13 9 1 10 13 9 9 2
21 3 13 10 9 1 15 9 1 15 13 1 10 9 1 10 9 1 10 0 9 2
1 0
5 9 12 2 9 13
5 11 12 9 1 13
22 15 8 13 3 1 15 9 3 4 16 3 9 1 9 1 4 1 10 9 11 13 2
26 10 0 9 1 10 9 13 4 4 1 0 0 9 1 10 0 9 9 7 0 1 12 1 12 9 2
36 1 15 9 13 9 1 9 1 15 13 1 15 13 1 10 9 2 7 8 10 9 1 10 9 11 1 11 7 11 1 11 13 9 4 4 2
16 8 15 9 3 1 10 9 9 13 2 4 15 3 1 9 2
22 1 15 9 4 3 15 13 1 10 9 2 9 12 2 8 9 2 9 12 2 0 2
5 11 11 4 13 9
1 9
20 15 13 1 9 1 9 5 9 13 1 15 13 1 9 2 13 9 12 2 2
13 3 13 1 10 9 1 15 9 13 9 4 4 2
7 3 13 15 9 7 9 2
10 9 12 2 9 2 9 2 9 7 9
3 11 12 9
1 9
11 9 4 0 4 1 10 9 1 10 9 2
15 15 13 1 15 9 2 9 12 2 13 3 3 4 4 2
20 15 13 16 9 16 15 8 1 12 0 10 0 9 1 12 1 9 4 4 2
26 10 9 1 9 2 9 2 9 7 9 4 13 2 7 1 15 9 13 10 0 9 1 10 9 3 2
13 15 13 16 8 9 1 13 9 7 9 4 4 2
13 1 10 9 1 10 9 13 10 9 4 4 3 2
2 13 9
2 13 9
2 0 9
34 13 9 13 1 10 0 13 9 4 2 8 16 10 9 10 0 0 9 13 7 13 1 0 9 15 0 4 1 10 9 1 10 9 2
42 16 10 9 1 0 9 13 2 13 10 13 9 1 10 13 9 4 4 2 16 3 9 2 8 5 11 2 2 9 2 8 7 8 2 7 9 1 9 2 8 2 2
13 3 13 15 9 1 9 3 10 9 9 13 4 2
1 9
1 9
1 9
1 9
1 11
10 9 2 13 2 9 2 9 2 13 2
28 13 9 4 3 13 1 15 13 1 10 0 9 1 10 9 7 1 10 9 1 10 9 7 9 1 10 9 2
19 15 9 13 3 1 9 4 2 7 3 0 0 4 4 8 9 7 9 2
17 1 15 9 13 15 1 9 2 16 10 9 1 15 0 13 4 2
8 15 9 4 4 1 15 8 2
9 10 9 1 9 7 9 4 13 2
38 16 10 9 1 9 13 2 15 13 3 4 4 1 10 9 7 9 1 10 9 2 13 1 10 9 16 15 3 0 13 4 1 9 2 9 7 9 2
18 8 9 13 3 10 9 1 9 3 10 0 9 1 15 9 13 4 2
1 9
32 0 9 4 3 4 1 10 9 13 1 10 9 7 9 1 10 9 1 9 7 1 15 13 1 9 7 9 1 9 7 9 2
20 15 9 4 3 3 4 8 9 7 13 7 3 2 13 2 9 1 10 9 2
