481 11
18 2 4 13 2 13 11 2 14 13 9 9 1 9 1 9 0 2 2
20 9 9 4 13 13 1 9 9 2 13 1 9 10 11 9 2 9 0 9 2
23 2 15 13 3 2 13 3 1 9 1 9 2 14 13 9 0 0 1 9 1 9 2 2
24 1 3 2 10 9 4 4 13 9 1 11 15 15 13 1 9 7 3 9 1 9 10 9 2
21 4 13 10 9 2 9 0 7 9 1 9 0 2 13 0 9 1 9 1 9 2
21 15 4 13 16 9 15 13 9 1 9 4 13 10 9 1 9 0 2 13 9 2
16 1 9 10 9 4 13 9 1 15 0 2 13 9 9 9 2
34 1 9 2 1 9 11 4 13 9 3 12 12 1 9 2 9 1 11 0 13 15 3 1 10 9 1 9 1 9 11 0 7 11 2
29 3 2 16 1 9 4 13 12 12 9 2 10 9 3 3 9 15 13 1 12 12 2 1 9 13 1 12 12 2
24 9 0 13 14 13 1 9 11 2 1 9 9 9 2 10 9 0 13 1 9 1 9 0 2
35 9 9 0 2 11 2 9 2 13 1 11 1 9 11 11 9 12 2 13 9 0 1 9 1 10 9 15 13 10 3 1 9 1 9 2
35 9 9 12 5 9 13 1 9 12 1 9 9 12 16 2 9 1 9 2 1 9 9 9 2 13 13 9 13 9 9 7 10 9 9 2
21 6 2 14 13 2 14 13 1 9 14 13 9 9 1 9 15 15 13 9 10 2
23 9 9 4 13 7 15 14 13 13 15 4 13 9 0 1 15 1 15 7 1 9 0 2
25 15 15 13 13 1 0 9 2 15 15 15 15 13 2 3 10 3 0 9 2 14 15 13 13 2
22 9 9 13 14 15 13 9 0 1 9 1 14 13 1 11 7 4 13 1 9 11 2
21 1 10 9 2 11 9 4 13 1 9 10 9 7 15 4 13 9 1 9 0 2
23 1 9 9 2 9 15 4 4 13 1 3 12 1 12 1 9 7 13 1 12 1 9 2
23 3 4 13 16 15 15 4 13 3 13 9 1 9 2 9 1 9 9 2 9 1 9 2
17 1 15 15 14 13 15 1 9 13 1 11 14 4 13 0 9 2
17 1 9 0 15 4 4 13 15 4 13 9 1 9 1 12 9 2
25 3 15 15 4 13 0 2 11 15 4 13 1 9 10 1 9 1 15 13 7 4 4 13 9 2
14 1 12 9 2 9 1 9 15 13 9 13 1 3 2
15 7 15 3 4 13 2 7 15 13 3 14 4 13 0 2
22 3 15 4 13 3 2 0 1 9 2 9 0 4 13 9 1 14 15 13 1 9 2
28 3 2 15 15 15 4 13 1 9 0 1 9 1 9 4 13 9 14 13 10 9 1 9 13 1 9 0 2
31 3 2 1 12 9 2 9 11 4 13 9 9 9 3 1 11 10 12 9 1 9 10 9 0 14 13 9 9 7 9 2
34 1 9 1 9 0 10 9 13 1 9 2 9 1 9 4 13 10 9 10 9 2 0 13 11 11 2 9 9 0 10 10 9 0 2
26 1 11 15 4 13 12 9 10 9 0 7 10 9 13 9 1 9 0 0 2 15 14 4 4 13 2
28 9 4 4 13 1 9 1 9 2 1 15 13 10 9 1 9 13 1 9 1 15 15 4 13 1 9 0 2
32 9 1 9 9 7 9 13 16 4 13 14 13 12 0 9 2 0 2 2 0 11 7 11 2 1 9 0 12 2 3 12 2
11 13 9 1 11 10 9 1 9 11 0 2
32 9 1 9 0 11 11 2 15 4 4 13 7 1 9 1 9 2 4 4 13 10 12 0 9 1 9 1 11 2 11 7 11
16 9 1 9 9 0 4 13 10 9 13 9 9 1 10 9 2
25 9 15 12 1 9 9 10 9 4 13 3 12 9 0 2 7 4 13 9 0 9 10 9 0 2
19 9 0 4 13 9 10 9 13 1 9 13 1 9 7 9 1 9 0 2
12 11 4 13 11 10 9 0 1 9 10 0 2
22 9 0 9 13 16 9 0 9 4 13 7 15 9 1 15 4 13 9 1 9 11 2
21 3 1 9 2 15 4 13 10 9 10 10 11 11 2 9 9 1 9 10 11 2
25 11 2 10 9 13 1 9 2 13 9 1 9 9 9 1 2 9 2 0 1 10 9 10 9 2
25 3 1 9 9 13 1 9 2 9 14 4 13 1 9 13 9 10 7 3 14 4 13 9 0 2
21 0 9 1 9 9 7 10 9 4 13 1 9 7 9 1 9 0 10 9 0 2
22 3 9 9 0 4 10 9 2 7 9 15 2 7 0 2 7 0 2 13 3 0 2
25 0 9 0 0 1 9 15 13 9 10 11 11 1 9 0 0 1 9 12 10 9 10 12 10 2
25 9 0 1 15 15 13 11 11 1 9 1 9 15 13 3 1 9 7 15 13 1 10 9 0 2
22 1 14 13 1 9 2 9 13 9 15 2 0 7 1 9 2 15 15 13 1 11 2
22 1 9 2 9 13 9 0 2 0 2 15 15 13 9 0 13 1 10 0 9 0 2
22 9 10 11 2 9 13 1 9 0 2 0 2 15 13 1 11 9 10 9 1 9 2
13 1 10 9 15 13 9 10 11 11 7 11 11 2
23 11 11 0 1 9 11 11 11 11 2 3 11 11 11 2 1 9 2 9 1 13 0 2
24 10 13 1 11 9 11 1 11 1 11 7 15 13 1 11 11 1 11 11 7 1 11 11 2
15 13 9 1 9 2 9 6 11 13 10 9 0 2 0 2
17 9 13 1 9 0 1 9 0 0 1 9 2 9 2 7 9 2
15 9 9 0 13 1 10 9 3 0 2 12 5 9 2 2
18 1 9 2 9 2 15 13 9 12 12 9 1 11 13 1 11 11 2
16 11 9 11 13 9 10 11 2 13 15 1 9 9 1 9 2
25 1 10 9 2 9 2 9 2 15 13 7 0 1 9 2 9 0 2 1 9 9 2 9 2 2
15 3 2 9 13 9 10 9 3 0 2 9 11 9 2 2
25 9 13 1 9 7 9 9 1 9 2 13 1 9 10 9 1 9 0 1 9 0 7 9 0 2
18 1 10 9 3 0 2 15 13 9 9 0 10 9 0 7 0 0 2
22 9 0 2 9 13 1 9 2 9 0 2 2 13 1 11 1 9 9 2 9 9 2
24 9 0 2 3 3 0 3 0 2 9 2 2 9 0 15 13 9 2 2 13 1 9 0 2
25 13 15 9 1 9 7 2 15 13 13 2 9 2 15 13 10 9 0 10 9 2 0 0 2 2
14 10 3 1 9 10 9 13 3 1 10 9 3 0 2
19 9 13 1 10 12 1 9 10 9 1 9 10 9 13 1 10 9 0 2
23 1 9 10 13 12 1 9 0 1 12 1 9 2 1 14 13 9 15 13 1 9 11 2
25 1 9 9 2 1 12 1 9 1 9 2 15 15 4 13 9 0 10 9 9 1 0 9 0 2
25 13 9 9 11 2 9 1 9 2 9 2 2 11 11 7 9 11 11 2 1 9 10 11 2 2
16 9 0 13 1 9 15 13 14 13 1 9 9 0 1 9 2
23 16 13 1 9 7 9 0 1 9 2 14 13 1 13 3 9 9 10 9 2 9 2 2
23 13 1 9 2 4 13 2 3 12 9 2 3 9 1 9 1 9 1 11 2 13 1 9
26 0 3 2 7 14 0 3 2 9 10 1 2 9 2 0 1 9 13 9 2 9 2 9 10 11 2
21 13 1 10 0 9 7 13 2 3 2 1 9 2 9 15 13 3 1 9 0 2
23 13 9 10 9 0 3 9 4 13 1 9 10 9 10 9 7 13 1 10 9 0 0 2
23 1 9 4 13 1 9 2 11 11 2 1 11 2 3 1 9 13 9 1 9 1 9 2
15 10 9 13 14 15 15 13 9 9 9 0 1 9 0 2
19 13 14 13 9 7 9 0 1 15 13 14 15 13 2 3 9 13 11 2
27 16 9 15 15 4 13 16 13 10 9 1 10 9 1 9 2 15 13 14 15 13 1 14 13 10 9 2
22 16 13 1 9 7 16 15 15 13 10 0 9 2 13 14 15 13 9 16 13 11 2
26 11 4 4 13 14 15 13 1 10 9 0 1 9 13 9 1 9 0 2 11 2 0 11 9 2 2
28 1 10 9 1 11 13 12 7 12 9 0 2 13 1 9 2 15 13 12 2 12 9 1 9 0 2 0 2
30 11 12 9 5 9 9 0 13 0 1 9 1 0 11 13 1 9 1 9 1 9 13 1 9 2 1 9 1 9 2
17 9 11 4 13 3 13 1 9 0 1 14 4 13 1 9 0 2
30 13 9 0 3 0 11 4 4 13 3 1 14 13 9 10 9 0 1 9 10 9 13 9 1 11 9 2 11 2 2
16 0 9 13 9 0 1 15 1 9 0 2 9 7 9 2 2
24 1 9 9 0 1 9 9 0 0 2 15 13 13 16 9 9 13 3 9 7 14 13 9 2
25 1 9 9 1 9 4 4 13 10 9 1 9 11 12 2 13 9 0 1 9 1 3 12 9 2
23 2 9 12 2 5 1 9 11 2 13 1 10 9 9 9 2 1 9 2 9 12 2 2
29 16 4 13 10 9 1 11 16 15 13 9 16 13 3 14 4 13 10 9 2 0 3 1 9 9 7 9 0 2
30 9 1 9 1 15 9 4 4 13 1 9 7 4 4 13 1 14 13 3 1 9 2 13 14 15 4 13 3 3 2
15 13 14 13 1 9 15 16 13 14 13 7 14 13 11 2
13 9 0 10 9 13 3 12 7 13 1 12 9 2
18 9 1 9 13 3 1 13 1 9 0 7 4 13 1 3 12 9 2
24 13 9 15 16 13 2 13 16 4 13 13 7 13 14 13 0 7 16 13 14 15 13 9 2
25 14 13 9 1 11 7 1 15 10 9 0 1 14 15 13 9 16 15 4 13 13 9 1 11 2
16 15 4 13 16 9 13 9 13 0 7 13 0 1 9 0 2
30 9 9 1 9 15 13 0 1 10 9 15 15 13 9 2 3 13 9 9 0 2 13 13 9 3 13 14 13 11 2
14 9 4 4 13 1 12 1 12 1 9 13 1 9 2
18 3 1 9 2 9 13 9 14 13 1 3 12 9 1 12 1 9 2
27 3 1 9 13 14 13 3 16 9 4 13 1 9 0 7 16 4 13 1 9 1 9 0 1 9 9 2
20 1 16 9 9 13 0 2 9 0 15 13 1 10 9 1 9 10 9 0 2
17 1 0 2 13 14 13 9 15 16 9 9 15 13 7 9 13 2
16 9 4 13 9 1 9 12 5 12 7 15 4 13 1 9 2
19 9 9 13 13 1 9 0 16 15 13 10 9 0 7 3 1 9 0 2
28 9 0 9 0 2 0 2 1 9 9 0 2 13 1 2 11 2 1 10 9 7 1 2 11 2 1 15 2
21 16 15 13 10 9 7 13 16 13 3 14 4 13 10 9 2 13 3 9 15 2
20 16 9 13 14 13 9 7 1 9 1 15 13 9 2 9 1 11 13 0 2
17 0 10 9 1 9 2 13 9 13 9 16 9 4 13 13 9 9
13 14 15 13 16 9 1 9 4 13 9 1 9 2
11 10 9 4 4 13 9 1 1 12 9 2
18 9 14 13 1 10 9 3 13 9 2 9 0 7 9 0 10 9 2
17 12 9 0 1 9 15 13 13 1 9 2 9 0 0 7 9 2
15 1 9 2 13 0 10 9 13 1 9 13 9 1 9 2
16 9 9 15 13 16 9 7 9 13 1 9 12 15 4 13 2
26 12 2 15 13 9 1 9 0 1 12 12 1 10 9 1 9 7 15 13 12 9 1 10 9 9 2
32 2 12 2 10 10 12 9 10 9 0 0 1 12 11 1 9 13 0 9 9 1 15 15 13 9 1 9 12 1 0 9 2
32 2 12 2 0 9 13 3 1 12 9 10 12 9 15 13 9 1 15 9 15 4 13 15 15 9 9 0 0 1 10 9 2
21 2 9 2 9 9 0 10 9 2 13 1 9 12 2 11 11 2 9 12 2 2
17 1 10 9 2 9 13 9 0 1 14 13 9 14 15 13 9 2
25 2 12 2 9 9 13 1 0 9 13 9 9 1 9 1 11 15 7 10 9 0 1 9 10 2
21 9 1 9 10 0 9 13 9 9 11 2 3 3 4 13 1 9 12 1 9 2
22 2 12 2 9 1 13 14 4 13 9 7 9 15 14 4 13 9 9 0 1 9 2
25 2 12 2 9 1 9 13 13 14 13 0 0 7 3 14 14 13 9 9 0 1 9 1 9 2
22 2 12 2 9 13 1 9 0 15 13 9 7 15 13 3 1 9 11 2 0 2 2
26 1 9 10 2 9 14 4 13 1 9 2 1 12 12 9 2 1 9 15 13 1 9 0 7 0 2
11 9 15 13 9 1 9 9 1 9 0 2
23 9 1 9 1 9 1 9 15 13 9 0 1 9 1 12 1 9 1 10 9 1 9 2
25 9 9 1 9 4 13 1 10 9 3 1 0 7 0 3 1 14 13 9 1 9 9 0 0 2
23 2 9 2 1 9 9 1 9 0 7 3 0 1 12 1 9 2 9 0 13 1 12 2
29 12 2 1 9 1 15 1 9 4 13 10 0 9 2 15 15 13 9 0 1 9 12 2 12 2 12 7 12 2
22 2 12 2 9 13 3 9 13 1 0 9 14 15 13 1 9 9 1 9 10 9 2
24 12 9 2 15 2 13 2 13 2 2 9 15 7 9 13 13 1 9 1 9 2 9 2 2
13 15 13 14 13 2 0 9 2 9 0 10 9 2
15 10 9 4 13 1 0 9 2 9 1 9 10 9 2 2
30 2 12 2 13 1 12 9 12 2 9 13 1 9 2 12 2 9 2 9 2 7 1 9 2 12 2 13 1 12 2
20 9 1 14 13 3 9 1 9 13 14 13 0 1 9 1 9 7 9 10 2
16 1 15 2 9 2 0 3 1 10 9 2 4 13 0 9 2
22 10 9 7 9 1 15 4 4 13 14 4 13 7 13 1 3 1 10 9 0 3 2
24 1 14 13 1 9 9 9 0 10 10 3 1 9 2 15 13 13 10 9 0 1 9 0 2
12 12 2 9 4 13 3 1 9 0 1 9 2
14 12 2 9 15 13 1 9 9 0 10 9 1 9 2
14 11 2 9 0 13 9 9 10 9 0 7 9 15 2
17 12 2 2 9 1 9 2 13 10 9 0 1 9 13 1 9 2
20 2 12 2 9 9 0 1 9 4 13 13 1 14 13 9 9 1 9 9 2
14 9 9 2 9 2 15 13 14 4 13 2 9 2 2
18 1 9 9 13 1 9 2 9 0 13 13 9 1 9 13 1 10 9
30 2 12 2 9 1 9 7 9 0 13 1 9 9 12 1 9 15 13 13 9 1 0 9 2 16 9 14 13 3 2
21 9 3 13 2 13 1 10 9 0 1 9 0 15 14 13 10 9 15 15 13 2
23 2 12 2 9 0 10 9 15 13 9 9 13 1 9 15 13 1 9 9 7 10 9 2
18 2 12 2 9 1 9 1 12 9 1 9 13 4 13 1 9 9 2
13 13 3 14 4 13 7 1 10 9 7 1 15 2
13 15 13 9 9 10 0 9 0 13 1 9 10 2
14 1 10 12 9 2 11 11 13 2 11 11 9 2 2
15 2 0 2 2 2 0 2 15 13 1 0 9 8 9 2
16 11 11 15 13 9 2 13 3 0 7 3 13 1 9 0 2
15 9 15 13 9 11 11 7 9 15 13 1 0 10 9 2
13 15 2 1 9 10 2 14 15 3 13 1 0 2
11 2 14 13 1 3 0 2 15 4 13 2
25 7 3 9 1 3 15 13 2 4 13 16 14 4 13 3 0 14 13 2 9 9 1 9 2 2
25 16 1 12 2 3 13 14 15 13 2 3 4 9 14 15 13 9 7 9 1 9 10 1 9 2
26 9 13 2 13 15 2 0 9 1 14 14 13 1 9 10 9 15 14 15 13 10 9 1 9 0 2
30 2 3 2 13 11 9 1 9 10 3 0 2 1 14 14 13 1 11 2 13 10 9 0 2 15 13 1 9 9 2
16 16 13 9 10 9 2 9 4 4 13 3 1 9 1 9 2
13 9 10 9 15 13 1 15 13 1 14 13 9 2
20 9 10 15 13 1 10 0 9 1 0 10 1 9 2 15 15 13 1 9 2
18 9 2 13 3 1 3 4 13 9 2 3 14 15 13 14 15 13 2
23 15 3 15 13 1 9 10 2 15 15 13 3 1 0 16 13 14 15 13 9 1 3 2
28 9 1 9 15 13 9 1 9 7 13 1 9 9 0 1 0 9 0 16 13 10 9 3 1 0 1 9 2
21 15 4 13 9 2 15 9 2 15 9 0 2 15 1 9 2 14 15 3 13 2
14 11 13 0 15 9 2 3 3 11 2 1 10 9 2
13 7 14 15 4 13 14 13 7 15 1 9 9 2
23 13 1 9 1 9 1 9 2 1 15 7 15 13 9 2 14 9 2 3 4 4 13 2
26 7 14 13 14 13 9 2 16 10 9 1 9 15 13 3 1 9 2 13 15 14 13 3 12 9 2
16 13 10 9 2 10 9 1 15 1 0 4 13 15 14 13 2
19 15 13 9 1 9 2 13 9 1 15 13 9 7 15 13 14 15 13 2
16 7 15 13 10 3 0 2 1 14 4 13 1 9 1 9 2
19 15 13 9 2 0 15 2 13 9 9 2 7 15 13 1 9 10 0 2
18 3 15 13 13 1 9 2 13 2 15 1 9 7 9 13 1 9 2
19 2 11 2 9 2 13 15 10 11 14 15 13 7 1 2 13 9 2 2
13 2 9 2 14 13 7 15 16 9 13 9 0 2
12 2 15 13 2 9 11 2 15 13 9 0 2
18 4 4 13 1 9 7 15 15 4 13 10 9 1 9 1 10 9 2
28 2 3 3 2 9 9 2 13 15 2 0 16 15 15 13 9 14 13 15 3 3 1 9 1 10 0 9 0
25 1 9 2 3 1 10 9 1 9 9 9 10 12 10 2 15 13 7 9 1 9 1 9 0 2
22 15 13 7 3 9 16 4 14 15 13 7 13 3 1 9 14 15 13 9 1 9 2
28 3 13 10 9 2 13 14 15 13 1 9 3 10 9 1 9 3 0 7 15 3 13 7 13 7 10 9 2
23 9 4 13 9 1 9 10 7 10 9 15 4 13 3 10 2 6 2 13 1 0 9 2
26 15 4 13 1 10 9 1 9 1 3 15 1 9 1 9 15 15 13 9 12 9 1 9 9 0 2
11 4 13 14 13 1 3 9 7 9 9 2
13 4 4 13 14 15 13 10 9 1 9 10 12 2
12 1 9 0 2 1 3 13 2 9 13 9 2
22 9 2 10 9 1 9 0 2 13 3 14 15 13 9 16 14 15 13 13 10 9 2
20 4 13 9 3 1 10 9 2 13 2 16 14 15 4 13 13 3 1 9 2
19 1 12 9 1 15 4 13 15 13 10 9 0 2 11 11 13 9 9 2
15 13 9 1 15 13 2 1 14 13 1 10 9 3 0 2
10 14 13 13 1 9 9 1 10 9 2
10 9 10 9 13 14 15 13 1 9 2
18 15 13 16 4 13 14 13 3 3 9 1 15 15 4 13 1 9 2
26 13 1 9 9 7 3 13 2 10 9 3 10 0 2 1 15 13 14 15 13 9 3 16 15 13 2
14 15 15 4 13 14 13 15 15 4 13 3 1 0 2
21 1 15 13 13 1 9 2 1 15 3 13 2 13 14 15 13 10 9 1 9 2
8 11 4 13 14 13 9 15 2
15 14 15 13 1 10 9 4 13 14 15 13 1 9 10 2
14 4 13 14 13 3 1 9 14 13 15 13 14 13 2
13 16 0 15 13 2 14 13 14 13 1 10 9 2
15 9 0 2 0 7 0 4 13 2 14 15 3 13 13 2
21 10 9 0 13 1 9 7 1 9 15 14 15 4 13 13 9 1 10 9 0 2
17 15 15 13 9 1 9 16 15 4 4 13 13 3 1 15 9 2
13 11 0 14 15 13 13 1 9 1 15 13 9 2
15 13 14 13 2 3 4 13 1 15 2 10 12 1 9 2
7 15 15 13 13 9 0 2
14 15 4 13 9 1 9 2 13 14 13 15 1 15 2
22 10 11 15 15 13 3 13 14 13 3 3 3 15 15 15 13 1 10 9 1 9 2
9 9 10 1 3 13 14 13 0 2
18 15 13 16 1 10 9 3 1 0 1 9 9 10 15 3 13 13 2
13 9 15 13 13 7 15 4 13 2 3 2 3 2
7 3 13 13 9 1 9 2
20 15 13 7 0 2 7 0 2 7 0 2 13 14 13 1 15 10 9 0 2
22 3 13 3 15 16 14 13 3 14 13 9 10 13 13 3 1 10 9 15 3 0 2
16 1 3 13 15 2 3 2 14 13 16 3 13 14 13 11 2
14 13 13 15 1 15 1 10 9 15 14 13 4 13 2
14 14 13 3 9 15 15 4 4 13 13 9 1 9 2
14 9 13 4 13 4 13 3 1 10 12 9 0 0 2
13 15 4 13 13 1 9 9 9 3 0 1 9 2
12 15 13 13 0 9 1 9 15 13 9 13 2
20 9 0 13 4 13 1 10 9 1 10 9 0 2 10 9 0 7 10 9 2
21 9 4 13 10 0 9 7 9 13 4 13 1 9 9 9 3 3 15 13 3 2
20 15 4 13 13 16 2 1 11 11 2 13 7 9 1 11 10 9 9 9 2
14 11 4 13 9 10 3 0 1 15 15 13 13 9 2
28 15 4 13 3 3 10 9 14 15 13 3 1 9 15 7 13 2 7 14 15 3 13 1 15 15 4 0 2
14 14 13 1 9 2 7 15 13 13 14 13 1 15 2
10 1 9 14 15 13 13 9 1 9 2
14 15 13 14 13 1 9 7 14 14 15 13 1 9 2
10 7 0 7 1 9 0 14 15 13 2
17 13 10 0 9 2 0 7 0 1 9 2 7 0 3 15 13 2
14 13 10 9 0 2 0 7 0 16 14 15 3 13 2
15 15 4 13 9 0 2 13 7 13 3 15 13 1 3 2
17 4 13 13 1 9 2 1 9 0 2 3 14 15 13 3 3 2
13 4 14 15 13 2 13 2 1 15 14 4 13 2
11 9 13 3 14 4 3 13 3 3 0 2
12 9 15 13 9 2 9 2 13 3 10 9 2
19 13 7 13 12 9 3 15 13 1 10 9 3 0 9 0 10 9 0 2
11 13 1 3 3 13 3 14 13 10 9 2
17 13 14 13 9 0 13 1 3 10 9 1 9 10 11 3 9 2
12 13 4 13 1 10 9 2 1 9 10 9 2
12 13 7 13 15 14 13 1 9 7 1 15 2
15 9 9 2 13 11 2 13 15 2 13 9 1 9 13 2
7 1 15 13 4 13 13 2
13 10 12 9 1 9 13 3 13 14 13 12 9 2
12 13 1 10 9 0 7 0 7 13 3 13 2
19 13 1 15 9 0 2 13 2 7 13 13 2 1 9 2 10 9 0 2
9 13 9 15 2 15 13 13 9 2
21 9 14 15 13 13 2 1 9 2 9 1 9 1 15 4 13 15 1 9 9 2
17 7 3 4 13 1 3 2 13 14 15 13 1 15 10 9 0 2
10 13 14 15 13 3 3 2 13 0 2
18 15 14 15 13 13 14 13 3 2 16 13 9 7 9 15 1 9 2
8 13 3 14 13 1 3 3 2
12 4 13 13 3 15 4 13 1 9 9 0 2
20 14 13 0 2 7 15 13 2 13 15 15 2 7 14 13 10 9 1 9 2
9 15 4 13 2 3 3 4 13 2
10 11 15 13 15 13 1 9 14 13 2
24 1 9 10 2 9 9 15 13 2 7 14 13 15 13 2 7 3 9 14 4 13 1 9 2
16 13 15 3 9 7 9 2 14 13 15 13 2 7 15 13 2
15 16 4 13 3 4 13 2 14 13 14 15 13 1 9 2
9 13 7 1 9 9 15 13 9 2
15 13 14 15 13 1 10 2 3 2 1 11 13 1 13 2
17 1 15 13 13 3 15 3 15 2 14 15 13 7 14 15 13 2
13 15 4 13 9 15 4 13 3 10 9 10 9 2
14 9 15 15 4 13 15 13 3 1 9 10 9 13 2
14 15 3 4 13 9 15 15 13 7 1 15 15 13 2
24 9 7 9 15 13 3 3 1 9 1 9 0 2 3 3 13 9 1 9 15 14 13 9 2
24 15 13 3 10 9 7 15 4 13 9 10 2 4 13 15 3 3 7 4 13 9 7 9 2
11 7 9 2 3 13 2 3 3 15 13 2
14 9 3 15 13 1 9 14 13 15 15 4 13 9 2
6 9 15 4 13 3 2
9 15 4 13 14 13 1 9 15 2
18 3 4 13 11 9 1 9 11 0 1 9 2 4 13 9 1 11 2
18 7 15 4 4 13 15 1 15 2 1 15 4 4 13 1 9 10 2
6 9 7 9 15 13 2
27 13 2 9 2 15 4 3 13 2 7 16 4 13 15 14 4 3 13 2 15 4 13 15 15 4 13 2
12 15 13 1 15 7 13 14 13 15 3 0 2
6 9 13 9 9 11 2
17 3 15 4 13 15 3 7 3 2 3 14 4 13 9 7 9 2
30 3 15 13 9 1 9 2 15 13 1 9 3 1 9 2 3 15 13 9 1 9 2 15 13 1 9 3 1 9 2
17 9 9 15 13 1 9 10 1 9 7 13 9 0 1 9 0 2
20 16 15 13 1 9 2 13 9 2 3 14 15 13 1 9 1 9 1 9 2
11 9 9 13 1 9 0 7 1 9 0 2
11 11 4 9 2 11 9 2 7 11 9 2
6 11 15 13 1 9 2
9 14 13 10 9 14 13 1 9 2
19 1 10 9 2 0 3 1 9 9 2 9 10 0 15 13 3 1 9 2
18 13 15 1 10 9 1 0 9 0 2 16 9 15 13 1 10 9 2
14 9 1 3 13 2 9 10 0 13 1 9 1 15 2
19 3 2 1 9 2 10 9 0 13 10 9 1 9 0 1 9 1 9 2
23 9 13 1 10 9 1 9 0 2 3 10 9 0 2 15 13 9 0 1 9 9 3 2
16 11 13 10 9 7 9 13 3 2 16 9 3 15 3 13 2
22 9 15 15 13 9 2 13 13 0 3 3 2 7 14 13 3 14 15 13 1 15 2
13 3 2 3 1 9 0 1 3 2 9 13 0 2
10 9 4 13 0 1 10 9 1 12 2
15 9 13 0 1 9 7 9 0 1 9 1 9 10 11 2
28 11 15 13 9 0 2 11 15 13 9 0 7 13 14 13 9 14 15 13 1 9 14 13 15 3 13 11 2
24 9 7 9 15 13 1 9 2 13 9 7 13 13 14 13 2 14 13 7 14 13 9 3 2
28 11 4 13 10 9 3 0 1 10 9 1 11 2 11 2 3 11 2 12 1 9 2 7 11 4 13 9 2
30 15 14 15 13 13 10 9 10 9 13 1 9 15 14 14 13 10 9 1 9 3 13 9 9 10 1 10 9 0 2
11 13 15 1 9 2 11 15 13 9 0 2
22 3 3 4 13 10 9 0 7 10 9 0 1 9 13 3 9 4 13 14 13 9 2
21 16 9 9 4 13 0 16 9 9 15 13 2 12 9 7 9 4 13 3 0 2
13 11 13 9 1 9 13 11 9 7 9 0 0 2
13 11 13 9 1 9 2 11 9 7 9 0 0 2
23 9 1 9 10 13 0 7 0 13 15 1 9 0 7 0 13 7 10 9 1 9 0 2
23 9 1 9 10 13 0 7 0 2 15 1 9 0 7 0 2 7 10 9 1 9 0 2
14 0 9 1 9 10 13 10 9 0 10 10 9 0 2
16 3 3 1 10 12 1 9 1 9 11 13 1 9 1 9 2
25 9 9 7 9 13 3 12 13 9 9 1 9 12 2 7 9 7 9 9 2 3 9 13 12 2
25 9 9 7 9 13 3 12 2 9 9 1 9 12 2 7 9 7 9 9 2 3 9 2 12 2
29 3 10 9 1 15 15 13 13 13 7 9 0 7 0 1 0 2 7 13 13 9 1 11 1 9 1 9 0 2
56 13 0 16 12 7 0 9 1 9 10 10 11 12 4 13 1 9 1 10 9 0 4 13 2 3 4 13 15 10 10 11 12 7 11 12 2 11 12 2 9 11 2 11 7 11 12 2 11 12 2 11 12 7 11 12 2
15 12 12 1 9 2 9 7 9 13 9 1 9 1 11 2
35 13 10 9 0 2 0 2 1 9 0 0 2 0 2 1 9 1 9 2 15 15 13 2 9 1 9 2 1 12 12 1 9 1 9 2
29 3 16 13 10 9 0 1 15 1 9 1 13 9 2 16 15 13 3 1 9 0 7 1 10 9 0 1 9 2
51 7 13 10 9 3 1 9 2 3 1 0 7 13 1 10 9 0 2 1 9 0 1 0 7 1 0 0 2 16 15 13 9 1 9 2 15 13 9 9 2 15 13 1 9 7 15 13 0 7 0 2
17 9 0 11 4 9 0 4 13 9 1 12 10 9 9 1 11 2
34 10 9 2 13 1 9 12 1 9 2 13 10 9 0 2 3 10 9 1 9 0 2 15 13 9 7 9 0 4 9 0 10 9 2
19 9 4 13 1 9 9 0 13 1 9 9 1 9 0 13 1 9 0 2
15 9 9 13 9 1 11 13 0 3 1 10 15 1 9 2
11 11 13 10 3 0 9 7 3 9 11 2
10 11 2 11 2 11 2 11 7 11 2
9 10 9 1 10 9 15 13 12 2
10 11 2 11 2 11 2 11 7 11 2
14 9 11 15 13 1 9 9 10 1 10 12 9 0 2
5 9 11 13 0 2
18 9 9 15 13 1 9 11 2 1 9 9 1 9 0 9 1 9 2
29 1 9 9 9 1 9 2 9 0 1 11 13 0 1 10 9 10 9 7 13 0 1 10 9 1 9 13 0 2
26 9 2 0 1 12 2 13 4 13 3 1 10 9 0 2 3 12 9 1 9 4 4 13 1 12 2
26 3 2 11 2 1 9 9 12 5 12 1 12 9 12 4 13 12 2 12 5 1 9 1 9 11 2
5 11 15 13 12 2
14 10 10 9 1 10 12 9 13 15 10 9 9 11 2
11 11 13 0 1 3 10 9 0 0 9 2
34 1 14 13 4 13 9 1 9 0 2 1 9 11 15 4 13 12 9 1 9 3 10 9 10 10 9 0 1 9 0 7 15 0 2
19 1 9 2 9 11 4 13 2 1 9 0 2 1 9 2 9 7 9 2
28 9 2 9 0 1 9 0 2 4 13 1 15 7 3 10 9 7 4 13 1 10 9 0 7 10 9 0 2
8 9 3 0 13 4 13 9 2
12 11 13 12 1 9 2 1 15 12 13 9 2
13 9 1 9 15 13 1 9 0 10 11 13 1 12
27 9 11 1 9 4 13 3 1 12 9 12 2 3 9 11 15 0 1 10 9 13 2 9 9 2 9 2
43 1 12 2 1 9 0 1 9 2 9 10 4 13 10 9 1 9 0 1 12 2 12 5 2 15 1 10 3 0 1 11 7 4 13 9 1 9 13 1 11 1 12 2
16 10 9 0 15 13 9 0 2 10 9 0 7 10 9 0 2
12 15 13 15 1 10 3 0 9 0 10 11 2
8 1 9 9 1 11 15 13 2
16 9 0 0 1 11 2 1 9 9 12 2 4 13 1 12 2
30 1 9 10 0 2 11 13 10 9 1 9 4 3 10 9 1 9 2 15 13 9 1 9 11 7 9 1 9 15 2
20 1 12 9 15 13 9 1 14 13 0 9 1 11 1 9 9 1 9 0 2
31 9 0 0 15 13 3 1 10 9 3 0 2 1 10 9 2 7 13 0 1 9 0 0 9 0 7 3 10 9 11 2
8 1 12 2 1 11 13 12 2
6 12 9 1 9 0 2
4 11 13 12 2
35 12 1 9 0 1 9 12 2 15 13 13 9 0 1 9 0 0 7 3 12 2 15 13 13 3 1 9 0 10 9 7 1 9 0 2
12 0 9 15 13 1 10 9 1 9 13 11 2
17 11 15 13 1 10 9 10 9 0 7 13 10 9 0 7 9 2
12 1 10 3 0 9 0 10 9 11 15 13 2
58 9 0 2 9 1 9 2 9 9 0 2 9 0 2 9 11 2 9 11 2 9 0 2 9 9 2 9 9 2 9 0 1 9 10 11 2 9 0 1 9 10 11 2 9 0 1 9 0 11 11 2 9 11 2 9 10 9 2
14 11 4 13 1 9 1 9 10 11 2 1 9 11 2
24 10 12 9 1 9 0 2 13 1 9 0 0 2 15 13 9 1 3 3 1 12 1 9 2
15 11 13 10 9 0 1 9 10 0 7 10 9 0 0 2
20 9 0 4 4 13 1 10 9 1 9 9 0 7 0 2 1 15 10 9 2
30 12 9 10 9 10 12 10 13 10 9 0 1 9 0 2 15 13 9 10 0 1 9 0 1 9 1 9 0 0 2
25 1 9 2 10 9 3 4 13 11 11 2 3 11 11 11 4 13 9 10 3 0 1 10 9 2
12 9 0 4 13 14 15 13 1 0 9 0 2
9 10 3 0 9 1 10 9 13 2
30 1 10 1 10 12 9 0 2 9 0 4 13 10 9 0 7 4 13 9 3 1 10 9 1 9 7 9 10 9 2
11 9 1 9 4 13 3 0 1 0 9 2
12 1 10 9 2 9 1 10 3 0 4 4 2
16 10 9 10 9 2 4 13 11 11 7 11 11 2 13 9 2
24 13 1 9 0 2 9 1 9 1 9 7 9 4 13 10 9 1 9 0 1 12 9 0 2
32 10 9 4 13 3 1 9 0 2 3 7 10 9 0 2 9 0 2 0 1 9 7 9 1 9 2 7 9 0 0 2 2
12 11 4 13 10 3 0 9 0 1 10 9 2
28 9 4 13 1 11 1 12 3 12 3 12 9 4 13 9 1 11 1 9 9 1 9 0 15 2 11 11 2
10 1 10 3 0 9 0 2 15 13 2
10 9 0 13 0 1 12 9 1 9 2
22 9 0 2 9 0 7 9 0 2 13 1 9 9 0 0 2 3 0 9 9 0 2
14 1 9 1 9 2 9 11 4 0 0 10 9 9 2
8 12 9 4 13 13 1 12 2
4 12 1 9 2
10 0 9 4 13 14 13 13 1 12 2
24 1 10 9 13 1 9 9 0 2 9 2 2 9 1 9 9 1 9 0 10 13 9 0 2
24 9 0 10 9 0 10 9 0 4 13 7 13 9 2 9 7 9 9 9 11 7 9 11 2
47 9 0 0 4 13 9 1 9 12 1 9 9 0 1 9 1 9 2 3 12 9 0 1 9 7 9 0 2 0 1 9 9 0 11 7 13 1 9 9 2 4 13 1 12 9 12 2
32 1 9 9 0 2 1 9 12 2 15 4 13 1 9 9 1 11 7 11 7 9 10 9 0 0 15 15 4 13 9 9 2
33 12 9 0 10 9 0 4 13 1 9 12 9 7 4 13 1 12 9 2 1 9 11 2 11 2 11 2 11 2 11 7 9 2
12 1 9 11 2 9 0 4 13 1 10 9 2
31 9 0 10 9 2 9 2 4 4 13 1 12 9 12 2 1 14 13 1 10 9 0 0 9 10 9 9 1 9 11 2
22 1 10 12 1 9 1 9 2 9 9 15 4 13 1 9 1 9 9 0 7 0 2
17 1 9 1 10 12 9 0 9 0 4 13 12 9 1 9 0 2
10 1 9 2 1 9 2 1 9 9 2
13 9 1 9 13 1 10 0 9 10 0 2 9 2
12 9 0 1 9 13 9 0 1 9 1 12 2
24 1 9 12 2 9 4 13 9 0 1 9 10 9 0 1 11 2 12 9 0 4 11 11 2
20 1 9 0 2 0 1 9 10 11 4 13 1 3 1 12 9 0 1 9 2
33 10 3 0 9 1 9 1 11 13 9 11 2 15 1 12 4 13 12 9 1 9 11 7 0 1 11 15 4 13 9 9 0 2
20 12 9 10 11 10 9 0 4 13 1 12 3 4 13 3 1 10 0 9 2
39 3 3 2 9 11 4 13 0 1 10 9 9 0 13 1 9 12 2 9 13 12 9 1 9 2 15 1 12 7 12 7 15 1 9 2 15 1 12 2
20 9 0 4 13 10 9 0 1 9 9 1 15 11 4 13 0 1 0 9 2
29 11 11 2 1 9 10 0 13 1 9 9 3 9 10 9 4 13 1 9 1 9 0 3 9 9 10 12 10 2
17 1 12 9 12 15 13 9 0 2 9 9 11 2 2 9 2 2
6 15 13 3 10 9 2
30 9 0 2 9 2 9 2 9 0 10 9 10 2 2 9 2 9 2 9 2 9 1 9 2 9 2 9 7 9 2
16 9 0 9 13 0 9 0 2 3 9 9 15 13 1 12 2
13 1 12 15 13 9 0 1 9 0 2 9 9 2
19 1 12 15 13 9 0 2 1 15 4 13 3 10 9 1 10 9 2 2
13 1 11 2 12 9 1 9 4 4 13 1 12 2
11 9 0 1 9 7 9 13 9 1 12 2
41 1 9 11 1 9 0 13 9 1 12 9 1 9 12 1 9 0 0 2 12 2 12 2 12 2 7 1 12 9 1 9 12 1 15 0 2 12 2 12 2 2
32 1 12 2 1 9 0 0 9 1 9 4 11 15 4 13 1 9 12 2 13 9 1 9 2 3 9 0 4 13 9 12 2
36 1 11 11 7 11 11 2 12 13 9 0 9 11 1 12 7 12 2 11 4 13 1 12 9 0 1 9 11 2 1 3 4 15 13 3 2
13 1 9 9 10 9 15 4 13 1 12 9 0 2
23 12 9 0 1 10 9 0 1 9 13 9 1 12 2 1 11 2 11 11 13 9 12 2
19 1 12 2 1 11 2 9 11 11 13 12 9 1 10 9 0 1 9 2
10 9 9 9 13 3 9 0 1 9 2
20 9 13 1 11 1 9 9 10 12 10 2 1 9 9 15 13 1 9 0 2
20 12 9 0 10 11 4 13 1 12 2 1 12 9 2 7 15 13 3 9 2
25 10 9 3 3 2 1 12 2 15 13 1 11 12 9 1 9 2 1 9 15 13 3 9 9 2
10 9 4 13 9 0 1 9 9 11 2
15 10 10 9 4 4 16 9 13 9 1 9 0 10 9 2
21 13 0 3 16 9 7 9 13 12 9 1 10 12 10 9 2 10 12 4 9 2
21 1 12 2 11 11 4 13 3 12 9 1 9 0 7 10 9 1 9 12 9 2
13 1 12 2 12 9 0 1 11 4 13 1 11 2
20 9 4 4 13 1 9 1 12 2 1 9 1 12 2 7 1 9 1 12 2
10 1 12 2 4 4 13 1 10 9 2
23 1 12 2 9 4 13 1 9 9 2 1 14 13 9 0 10 9 2 13 1 11 11 2
36 1 12 7 12 2 9 4 13 9 11 2 3 2 1 12 7 12 2 3 11 3 7 11 4 13 9 1 3 10 9 0 10 11 7 11 2
25 1 12 2 3 9 10 12 9 4 13 0 2 1 9 1 11 2 9 9 4 4 13 1 11 2
21 1 14 13 9 13 9 1 12 2 1 9 9 9 2 15 4 13 9 10 12 2
25 1 12 2 9 1 9 7 9 4 4 13 3 1 15 1 9 7 9 2 7 9 1 9 0 2
16 4 4 13 9 0 2 1 9 9 2 9 0 7 9 9 2
10 1 9 12 2 0 14 13 9 11 2
13 10 12 9 0 4 13 10 9 0 1 9 0 2
33 1 9 12 2 9 4 13 9 10 9 0 1 9 0 7 9 0 2 9 1 15 10 0 9 1 9 0 10 9 4 4 13 2
10 1 9 2 9 13 0 1 9 0 2
10 9 9 13 14 4 13 1 9 9 2
9 9 9 4 13 3 13 1 9 2
30 1 9 0 2 9 9 4 3 13 1 9 7 9 1 0 2 15 4 13 10 9 2 3 9 9 0 4 4 13 2
14 15 4 4 13 10 9 3 3 2 1 12 9 12 2
19 9 15 13 1 9 11 2 10 9 10 9 2 15 15 13 1 9 11 2
45 1 9 10 2 9 13 0 9 10 10 12 9 9 2 11 2 11 2 11 2 11 2 11 7 11 2 1 9 13 1 12 9 1 9 9 7 12 9 1 9 11 7 9 11 2
11 0 9 13 11 2 9 2 9 7 9 2
46 9 3 13 13 1 9 11 7 1 9 9 2 0 1 9 0 9 2 16 3 15 13 9 2 2 1 9 1 9 2 13 9 0 2 1 15 4 13 3 12 9 1 9 1 9 2
69 9 0 15 4 13 1 10 9 2 13 1 12 9 2 9 12 2 9 11 2 9 2 9 2 9 2 9 2 9 7 3 11 7 9 2 1 10 12 9 2 9 12 2 2 4 4 13 9 9 2 9 0 2 1 9 2 2 11 2 9 0 2 1 9 2 3 0 9 2
34 9 13 3 9 10 9 15 2 1 9 1 9 0 2 4 13 3 9 0 2 7 2 1 9 1 9 0 2 15 13 3 9 0 2
9 11 2 11 2 11 7 9 9 2
25 9 13 10 9 0 0 2 13 13 1 9 1 9 1 9 0 2 9 13 0 2 3 9 0 2
23 1 9 9 1 12 2 9 4 3 9 1 9 10 12 9 10 11 1 11 2 13 12 2
4 12 1 9 2
3 12 9 2
22 1 12 9 0 10 9 0 1 9 2 9 9 11 13 2 1 9 12 2 1 12 2
31 9 13 9 0 9 2 10 12 0 9 2 10 9 9 1 9 1 9 0 7 10 12 9 0 0 2 9 1 9 2 2
4 12 1 9 2
13 9 0 2 9 1 9 2 4 4 13 1 12 2
9 11 13 10 9 0 0 10 11 2
24 9 0 7 15 10 9 4 13 9 1 12 9 2 0 9 7 9 1 9 4 0 1 9 2
20 10 9 13 1 9 1 9 2 9 9 9 2 11 2 11 9 11 3 2 2
8 10 9 0 1 9 0 13 2
11 12 9 1 9 4 4 13 1 9 9 2
11 9 9 11 13 10 3 0 1 9 11 2
11 1 9 1 9 10 9 2 1 9 9 2
32 1 9 1 9 0 2 11 1 3 15 13 3 10 0 9 1 11 7 11 2 1 9 7 9 2 1 9 2 9 7 9 2
22 1 9 0 9 0 15 4 13 1 9 0 9 0 1 9 9 12 9 7 9 11 2
38 7 0 9 9 15 4 13 1 9 0 2 3 15 4 13 10 0 9 10 9 0 2 1 14 15 13 9 1 9 16 15 1 9 0 13 9 9 2
12 10 12 9 1 9 9 13 1 9 1 9 2
6 1 9 13 12 9 2
23 9 11 2 12 2 2 9 0 11 2 9 11 2 9 11 7 10 9 1 9 1 11 2
12 1 9 12 9 13 12 9 1 9 0 9 2
13 9 1 9 13 9 1 9 9 9 2 12 2 2
24 1 12 2 9 0 1 9 1 11 4 13 0 9 2 13 12 9 1 9 0 0 1 9 2
17 9 0 9 12 13 0 7 0 2 13 13 1 10 9 1 9 2
8 10 9 1 11 13 9 0 2
16 1 12 9 9 4 13 13 2 16 13 3 10 9 3 0 2
16 9 4 13 1 9 2 7 1 10 9 15 4 13 9 15 2
33 9 1 9 11 11 4 13 1 12 9 0 9 9 2 12 9 1 9 11 11 0 1 11 7 12 9 11 8 0 1 9 11 2
13 14 13 9 1 14 12 4 7 10 12 1 9 2
10 9 0 1 9 2 1 9 7 9 2
9 12 12 1 9 4 13 1 9 2
