790 17
24 1 0 0 9 0 9 1 9 11 4 13 12 9 7 9 1 12 9 11 2 11 7 11 2
17 11 4 13 9 0 9 2 7 15 15 4 13 13 1 0 9 2
8 9 9 9 9 13 0 0 2
18 0 9 13 0 9 2 0 2 0 7 0 13 0 7 0 1 0 2
22 13 15 3 16 0 9 2 1 9 2 9 2 9 2 1 9 7 13 3 0 9 2
18 1 9 9 15 3 13 9 1 9 2 9 2 9 2 9 7 9 2
10 7 0 9 11 13 14 3 0 9 2
20 9 0 12 9 13 0 1 10 9 7 14 3 15 1 11 10 9 13 3 2
20 3 14 13 9 1 0 9 2 7 4 10 9 1 9 13 3 0 0 9 2
24 1 0 9 15 3 13 9 2 13 9 0 7 3 3 0 2 14 3 7 3 13 0 9 2
29 1 12 1 2 9 2 11 13 14 3 0 9 2 13 7 3 16 9 0 9 2 16 13 1 9 1 10 9 2
12 1 10 9 13 1 9 0 9 0 9 11 2
39 1 0 9 4 10 9 13 1 15 2 16 13 11 0 0 9 1 9 9 2 9 7 9 2 7 14 13 2 16 15 1 15 13 14 9 1 0 9 2
37 9 14 13 2 16 4 13 1 10 9 11 1 10 9 0 11 16 1 9 1 11 2 7 15 14 1 0 9 3 3 3 13 9 9 1 9 2
17 1 11 13 3 9 1 9 7 9 2 7 9 13 1 10 9 2
6 3 15 9 3 13 2
22 1 9 13 9 2 13 1 9 9 7 0 0 9 7 13 1 0 9 1 15 9 2
10 3 15 10 9 14 14 13 1 9 2
31 3 0 4 13 1 9 10 9 2 16 15 4 13 12 1 9 1 9 0 9 2 16 15 4 13 12 1 0 0 9 2
23 9 13 7 2 16 1 9 1 10 9 3 13 14 9 2 7 14 13 13 1 0 9 2
16 1 9 9 9 13 3 0 13 2 3 0 9 13 0 9 2
18 1 0 9 7 14 13 13 10 0 9 2 16 4 2 13 2 9 2
11 9 13 3 3 1 0 9 9 7 9 2
20 16 15 9 13 1 9 2 13 9 3 1 15 2 16 0 9 13 0 13 2
15 14 9 7 9 13 3 7 3 2 3 13 0 0 9 2
32 10 9 1 12 9 13 0 9 1 9 9 2 1 0 9 7 13 0 9 2 1 15 14 14 4 13 0 13 1 0 9 2
16 11 13 0 9 2 1 15 11 13 10 0 9 1 0 9 2
7 15 3 0 3 14 13 2
38 3 13 14 1 10 2 3 0 2 9 9 0 0 9 2 7 13 1 9 1 2 0 9 2 1 0 9 9 7 2 0 9 2 1 0 9 9 2
45 0 9 4 13 14 14 0 1 0 9 2 16 4 9 13 16 9 1 0 9 0 9 7 0 9 0 2 0 9 2 7 9 13 1 11 3 3 2 0 2 9 16 0 9 2
45 16 15 14 13 1 9 2 4 13 3 0 9 13 16 9 2 0 14 1 10 0 9 2 3 4 15 3 13 1 0 9 2 16 4 13 0 0 9 9 1 0 9 0 9 2
14 0 9 4 3 13 0 9 14 1 10 9 1 15 2
10 0 9 15 13 1 0 9 7 9 2
20 16 13 14 10 9 1 9 2 3 3 1 9 13 1 9 2 16 13 9 2
5 1 9 13 9 2
24 11 13 1 9 0 9 1 9 0 9 11 11 12 1 0 9 1 0 9 9 1 0 9 2
7 0 9 13 1 0 9 2
5 9 9 1 0 9
25 16 13 1 0 9 2 16 15 1 10 9 13 1 9 2 3 13 0 9 2 16 13 15 0 2
30 10 12 9 1 9 13 7 0 1 9 2 9 2 9 7 1 9 9 0 9 2 1 9 7 3 13 3 1 9 2
47 16 7 15 0 9 14 13 13 1 9 2 15 3 13 1 9 1 0 0 0 0 9 11 11 7 1 11 7 7 15 1 0 9 13 0 9 0 2 0 2 0 2 0 7 0 9 2
23 1 9 2 15 13 1 0 9 2 4 11 13 2 16 13 0 1 15 2 15 9 13 2
4 0 13 0 2
10 11 4 13 2 16 13 0 9 0 2
35 1 9 1 9 0 9 4 11 13 2 16 4 13 0 9 14 1 9 1 15 2 15 4 13 9 1 0 9 2 16 4 3 13 9 2
6 11 4 13 0 9 2
17 1 9 13 1 0 9 2 1 15 13 0 2 16 9 14 13 2
12 3 4 9 13 9 2 7 14 13 10 9 2
10 9 13 3 13 3 2 1 0 9 2
24 11 4 13 2 16 4 0 9 13 2 0 15 13 13 2 15 13 0 1 9 1 0 9 2
5 9 9 13 9 2
29 16 3 13 2 13 1 9 13 3 3 2 13 7 15 13 14 9 2 16 15 1 15 3 3 13 1 10 9 2
11 9 13 12 1 0 9 2 16 13 9 2
28 9 15 1 9 13 2 16 13 1 9 7 16 15 3 0 9 13 10 9 2 7 15 13 1 10 9 9 2
20 3 15 15 13 0 13 2 16 4 13 9 7 0 9 2 16 15 15 13 2
19 14 13 2 16 15 9 7 9 3 13 2 16 15 13 9 7 0 9 2
13 14 15 13 0 13 1 9 7 9 13 9 9 2
21 14 15 16 9 9 14 13 15 7 7 14 3 3 1 10 9 2 16 4 13 2
7 9 13 0 2 0 9 2
12 16 15 13 15 2 15 15 13 1 0 9 2
17 13 7 3 13 15 13 0 9 7 13 9 2 16 15 15 13 2
29 1 15 13 10 9 2 7 16 13 15 0 9 2 9 0 9 7 9 15 7 15 0 1 9 2 16 13 0 2
24 13 2 16 9 1 10 0 9 13 9 2 7 16 13 10 0 9 2 1 15 15 13 15 2
10 10 0 9 13 12 3 0 9 9 2
34 13 15 1 0 9 7 0 9 2 1 9 9 2 1 9 9 7 1 0 2 0 9 2 16 15 13 2 9 2 7 2 9 2 2
9 9 3 13 10 9 15 16 9 2
11 10 9 9 13 3 0 9 2 16 13 2
8 10 9 15 13 0 9 9 2
15 9 9 7 9 3 13 9 9 2 16 4 15 13 13 2
18 9 9 7 9 12 9 9 13 1 0 9 2 1 15 3 13 9 2
19 0 9 2 16 15 13 13 2 14 13 9 2 9 2 9 7 0 9 2
30 16 15 13 1 9 7 13 10 9 1 0 9 2 15 13 2 15 9 13 7 10 4 13 10 9 1 0 0 9 2
27 3 13 10 9 2 15 9 13 13 7 13 1 9 2 1 15 7 14 13 14 0 9 1 10 9 9 2
18 15 4 3 13 0 9 9 2 16 13 2 16 9 13 15 1 15 2
19 14 3 4 13 9 7 7 4 1 9 13 10 9 7 9 1 0 9 2
30 15 13 9 2 16 15 13 3 13 2 16 4 3 13 2 3 15 4 9 13 7 3 3 16 1 9 1 0 9 2
17 9 13 0 9 2 16 15 9 13 2 16 4 15 13 1 9 2
20 9 1 9 3 13 2 7 16 13 1 0 7 0 9 9 2 0 1 9 2
18 16 4 3 13 1 10 9 2 15 4 10 9 13 10 9 1 9 2
8 13 4 2 16 4 9 13 2
17 1 9 1 10 9 4 13 13 2 16 4 15 9 13 1 9 2
18 16 4 10 9 13 3 2 15 4 13 2 16 15 9 13 1 9 2
16 1 10 9 15 4 13 1 9 2 16 13 2 16 4 13 2
16 0 9 15 4 1 10 9 13 2 16 2 4 13 9 2 2
20 10 9 4 3 13 2 1 15 4 9 3 13 2 16 2 4 13 9 2 2
10 3 4 10 9 13 2 1 15 13 2
12 2 9 4 13 2 16 4 1 9 13 9 2
10 2 7 4 13 2 2 4 14 13 2
11 0 9 13 3 3 0 9 1 10 9 2
22 3 13 10 9 7 1 9 15 1 0 2 0 7 0 0 9 13 3 3 7 3 2
14 1 11 7 14 14 1 15 13 13 9 9 7 9 2
8 3 13 1 9 0 1 15 2
23 1 10 9 7 15 4 13 2 3 15 13 9 1 10 9 2 7 1 9 4 15 13 2
14 13 4 15 1 9 0 9 1 9 7 13 10 9 2
8 9 15 3 13 3 16 9 2
17 3 4 13 1 9 1 9 2 13 9 7 15 13 13 10 9 2
22 2 9 2 16 13 1 9 2 16 13 9 2 13 1 9 9 1 9 1 9 9 2
20 9 12 9 8 13 1 9 9 1 0 9 2 16 13 0 1 9 0 9 2
11 1 9 2 9 2 9 7 13 0 9 2
7 1 9 9 13 0 9 2
17 15 13 10 0 9 2 16 13 1 0 9 2 7 9 1 9 2
9 9 10 9 13 1 3 0 9 2
9 1 0 9 13 9 0 1 9 2
8 1 11 13 12 0 0 9 2
6 10 9 13 0 9 2
17 9 1 9 13 0 7 0 1 9 7 9 1 9 7 0 9 2
8 9 13 0 1 0 9 11 2
16 9 1 0 9 13 1 10 9 2 16 13 9 1 9 11 2
24 14 2 7 13 2 16 13 0 2 16 4 15 13 1 10 9 2 16 15 13 13 0 9 2
19 9 7 12 12 9 4 13 1 0 0 9 2 16 4 15 3 13 9 2
12 15 13 0 9 10 9 2 0 9 15 15 2
6 0 9 13 10 9 2
30 9 11 13 2 16 4 11 3 13 3 12 2 0 0 9 2 16 4 0 9 1 9 0 0 9 13 1 12 9 2
36 9 12 4 0 0 9 13 12 9 9 2 1 12 9 3 16 9 12 2 7 1 15 13 1 0 9 11 2 1 15 15 11 13 1 9 2
49 9 9 1 0 9 7 0 9 1 12 9 2 15 4 13 0 9 9 2 16 4 13 9 1 9 1 9 14 1 9 9 2 14 3 13 12 9 0 9 2 11 2 11 2 11 7 11 2 2
39 1 10 9 13 11 11 1 0 9 13 1 3 0 7 0 0 9 2 16 13 0 7 1 9 9 16 14 1 0 0 9 7 9 0 9 7 0 9 2
26 7 15 13 15 2 16 15 4 13 1 3 13 1 2 9 2 0 9 2 0 9 7 0 9 2 2
9 1 9 0 9 13 10 9 0 2
28 15 13 2 16 15 4 0 9 9 13 1 0 0 9 2 12 9 2 2 16 4 13 14 0 9 10 9 2
30 9 9 0 9 13 9 9 1 9 1 10 0 9 2 9 9 1 0 9 1 9 7 9 9 7 0 9 1 9 2
19 9 4 13 9 1 9 11 1 11 2 1 10 9 7 4 15 13 11 2
19 0 13 0 7 0 2 14 0 7 13 3 2 16 15 13 1 0 9 2
15 15 13 14 1 11 2 16 4 3 13 9 7 13 9 2
15 2 0 9 15 3 3 13 2 7 13 9 2 16 13 2
19 1 15 13 3 10 0 9 1 9 2 3 7 4 13 14 1 9 3 2
29 1 9 4 13 2 16 4 9 2 16 4 3 1 9 3 13 1 0 9 1 0 11 2 13 0 9 0 9 2
11 9 1 11 13 1 3 12 12 9 9 2
12 16 13 1 10 9 1 9 2 13 0 9 2
22 10 9 13 9 2 16 15 1 3 9 10 0 9 13 0 9 2 0 9 9 8 2
24 16 13 10 9 1 0 8 2 15 13 9 2 16 15 14 3 13 2 16 13 10 9 9 2
12 15 3 13 1 0 9 7 9 1 0 9 2
9 9 15 3 13 7 3 13 9 2
23 1 10 9 13 10 9 1 0 8 7 9 10 9 9 13 1 9 2 16 13 1 9 2
13 1 0 9 7 8 13 0 9 2 1 9 9 2
14 9 13 9 2 16 9 14 13 2 7 13 3 9 2
5 2 15 14 13 2
19 9 15 4 13 0 2 7 4 13 1 9 12 0 0 9 2 9 11 2
43 11 11 2 9 9 1 11 11 2 16 13 1 9 0 11 7 9 0 9 2 7 15 4 1 9 3 13 2 16 4 0 9 13 13 0 9 1 9 1 12 9 3 2
31 3 4 13 1 9 0 11 2 16 4 13 3 13 9 2 7 9 1 11 2 16 4 13 10 9 2 14 3 13 0 2
51 9 11 13 14 3 1 9 7 4 13 3 1 9 14 12 0 9 1 10 9 2 3 7 4 3 13 1 9 14 1 12 9 1 9 0 9 7 1 12 1 9 1 0 11 1 11 8 11 1 11 2
7 9 4 13 1 10 9 2
32 2 1 3 0 7 0 9 9 7 14 4 13 14 2 16 4 0 9 15 13 1 9 7 9 0 9 2 2 13 11 11 2
8 2 0 9 13 0 1 9 2
29 11 13 3 0 1 0 9 1 9 2 16 14 3 13 0 9 2 16 13 1 9 10 9 3 10 16 12 9 2
27 14 9 1 9 4 13 1 9 1 10 16 12 9 2 16 15 4 0 0 9 1 0 9 13 1 11 2
9 2 14 13 3 2 3 13 0 2
15 10 9 4 13 0 1 12 9 2 7 4 13 0 9 2
7 0 9 4 13 0 9 2
29 0 9 1 9 15 15 14 13 3 15 0 2 13 7 1 9 2 1 15 4 3 2 13 2 9 1 0 9 2
11 0 9 13 14 9 2 16 13 1 9 2
29 1 3 12 9 15 4 13 9 7 0 9 11 4 1 11 13 0 9 0 9 2 16 15 1 9 4 14 13 2
24 16 7 13 3 9 14 0 2 3 3 13 1 9 2 16 15 13 15 2 15 4 3 13 2
14 16 15 1 15 14 4 13 2 13 1 9 0 9 2
13 9 13 15 2 16 1 15 3 13 1 0 9 2
3 2 11 2
10 9 11 15 4 13 9 1 9 11 2
43 0 9 2 9 11 2 9 2 1 15 4 0 0 9 13 14 3 2 16 4 15 1 0 9 13 1 0 9 1 0 9 2 0 9 3 13 9 1 9 0 9 11 2
31 0 4 1 9 9 1 12 9 13 2 16 14 13 1 10 9 2 7 13 1 9 10 9 1 10 9 7 1 10 9 2
8 13 4 2 16 13 3 0 2
18 13 4 15 13 0 14 2 16 4 13 9 2 16 4 0 13 9 2
14 12 9 15 14 13 2 3 4 1 9 13 0 9 2
28 10 9 7 4 13 14 15 2 16 4 9 1 9 13 1 9 11 7 11 7 13 2 16 13 0 1 15 2
11 1 0 0 9 15 1 9 3 13 9 2
18 7 13 3 2 16 1 0 9 1 9 13 9 2 9 9 12 2 2
19 1 10 9 13 0 9 2 16 14 1 9 14 13 1 9 9 1 9 2
18 11 4 13 1 9 2 7 15 4 9 13 2 3 4 13 1 9 2
24 1 9 9 1 0 9 4 11 13 2 16 4 0 9 9 13 1 9 0 9 7 0 9 2
31 1 0 9 2 16 15 13 1 0 9 2 4 13 9 7 9 9 1 0 9 0 9 7 9 1 0 9 7 0 9 2
78 0 9 1 11 2 1 9 0 0 9 4 13 1 9 2 12 9 2 0 9 2 1 15 4 15 13 0 0 9 9 1 11 2 0 0 9 2 1 9 2 2 16 13 1 9 9 1 9 11 11 2 0 9 9 7 4 13 0 0 9 9 11 2 16 4 1 10 0 9 0 9 12 9 13 0 0 9 2
23 0 0 9 4 13 0 9 3 0 0 9 2 0 7 15 13 14 1 9 1 0 9 2
68 16 13 9 14 9 0 9 7 0 9 9 0 9 11 1 9 7 9 2 13 3 13 11 11 2 16 4 10 9 13 1 9 2 15 1 9 7 15 4 13 11 11 2 16 4 1 9 3 13 11 7 3 13 1 0 9 1 0 9 13 9 7 9 13 1 0 9 2
21 11 11 2 16 4 15 0 0 9 13 10 9 2 4 1 15 3 13 10 9 2
47 0 9 11 11 2 16 4 13 14 1 0 9 12 0 9 2 4 1 0 7 0 9 13 1 9 1 9 9 7 3 13 9 1 9 2 16 15 4 3 13 14 14 3 0 11 11 2
17 3 15 15 13 2 16 15 4 9 13 3 1 10 9 10 9 2
46 1 15 11 13 2 16 15 13 3 0 13 9 9 2 1 15 15 4 12 9 13 1 9 2 7 4 13 0 9 2 16 9 2 16 13 0 7 3 0 9 1 0 9 2 13 2
8 0 9 15 15 3 14 13 2
10 9 4 13 1 9 12 1 0 9 2
30 10 9 4 13 12 0 9 1 9 9 7 9 0 0 9 2 16 15 4 1 9 1 9 1 10 9 13 0 9 2
11 14 9 9 7 9 13 0 7 0 9 2
21 13 2 16 13 10 9 3 0 2 7 16 13 0 2 13 13 10 9 1 15 2
10 14 0 9 15 15 4 13 1 9 2
15 16 0 9 13 9 0 2 4 3 13 1 10 0 9 2
7 14 4 13 13 0 9 2
25 11 4 13 15 2 16 4 13 7 1 9 13 2 16 9 13 9 2 7 1 9 15 13 9 2
33 0 13 2 16 4 15 13 14 1 9 2 16 4 3 7 3 0 2 1 9 0 9 13 1 0 0 7 3 0 2 0 9 2
25 10 9 9 4 13 9 9 1 9 0 9 2 9 3 2 16 4 10 9 13 0 9 7 9 2
4 13 0 9 2
41 0 0 9 10 9 1 9 0 9 4 1 0 13 2 16 4 13 9 15 2 16 4 13 3 0 2 1 15 16 15 4 13 0 2 15 0 9 7 0 9 2
16 9 10 9 13 9 9 2 15 13 0 1 0 9 10 9 2
13 1 0 9 9 9 12 9 0 9 9 4 13 2
28 9 3 7 3 13 10 9 2 7 15 9 3 14 13 14 1 9 2 16 4 13 0 7 3 0 11 9 2
20 9 9 0 9 13 1 9 1 9 0 2 7 13 1 9 10 9 3 9 2
29 7 4 15 1 0 9 1 9 1 0 9 14 1 9 13 2 16 13 9 1 9 12 0 9 1 0 0 9 2
11 0 13 9 9 1 0 9 7 9 9 2
22 15 1 11 3 13 1 9 9 0 9 2 7 7 15 14 13 1 9 0 0 9 2
24 12 9 0 9 2 9 10 9 4 1 9 15 0 13 12 9 9 11 7 11 11 1 11 2
16 7 16 4 15 9 12 13 2 4 13 1 15 14 9 11 2
16 9 12 4 1 9 11 13 10 9 7 15 13 14 0 9 2
24 1 9 4 3 12 2 0 11 13 1 0 0 9 2 9 7 4 1 12 9 13 16 9 2
8 15 7 14 4 15 4 13 2
5 3 13 0 13 2
9 13 13 0 7 14 3 15 13 2
26 3 7 14 13 2 3 14 13 9 7 13 2 16 13 9 2 16 4 2 13 9 2 3 14 3 2
7 15 13 2 1 15 13 2
5 7 9 16 9 2
13 1 11 4 15 3 13 9 7 9 0 9 11 2
19 13 4 0 2 16 13 1 9 1 9 2 16 13 1 9 3 3 0 2
10 3 7 4 13 13 2 4 13 9 2
4 13 4 9 2
7 13 4 13 3 16 3 2
5 13 4 13 0 2
8 11 4 13 1 9 0 9 2
13 16 4 15 13 9 2 4 14 3 13 10 9 2
11 1 10 9 15 4 13 10 9 1 9 2
11 9 15 4 13 9 2 16 13 3 0 2
15 3 1 9 4 13 2 16 13 15 2 15 14 4 13 2
16 3 4 13 15 15 2 14 16 4 10 0 9 13 0 0 2
13 3 15 4 13 13 1 10 9 2 1 10 9 2
8 0 9 4 3 3 13 0 2
15 11 4 13 2 11 7 15 4 13 16 9 1 0 9 2
8 9 9 12 4 13 3 9 2
18 1 10 9 4 15 13 2 16 4 13 1 9 9 2 16 13 3 2
18 12 9 3 2 16 4 13 1 0 9 2 4 13 10 0 9 9 2
22 13 4 2 16 4 13 0 7 0 2 16 4 15 13 1 10 9 2 1 10 9 2
16 14 0 4 13 2 16 4 15 13 1 11 2 1 10 9 2
12 13 4 0 0 2 14 16 4 13 1 9 2
10 1 12 9 0 9 4 13 1 11 2
19 13 15 4 1 0 9 7 1 9 13 11 2 9 7 9 1 0 9 2
11 11 4 13 0 1 10 2 0 9 2 2
19 3 3 4 13 1 9 1 0 9 2 7 3 4 13 10 9 7 9 2
13 2 15 4 3 13 1 9 2 2 13 3 11 2
15 13 15 4 9 7 15 3 13 2 16 4 13 3 0 2
16 9 2 0 0 9 9 2 2 9 1 0 9 13 0 9 2
9 14 0 9 10 9 13 9 9 2
16 13 0 9 1 9 2 16 13 0 0 9 7 0 9 9 2
13 9 9 9 15 13 13 1 9 9 7 0 9 2
19 2 9 9 14 13 1 0 2 7 1 15 13 9 1 9 7 13 9 9
5 9 13 3 0 2
10 0 0 0 9 9 7 13 0 9 2
6 9 3 14 13 3 2
5 14 15 14 13 2
5 1 9 9 9 2
5 1 9 1 9 2
28 14 4 7 15 13 13 2 16 4 15 3 13 1 10 3 0 0 9 2 16 4 14 3 13 1 0 9 2
13 1 9 13 14 9 9 2 16 13 1 9 9 2
28 3 13 3 13 9 9 0 9 1 9 0 9 2 16 13 1 15 0 9 7 9 15 13 14 1 0 9 2
26 9 0 9 11 11 4 13 2 16 0 9 9 13 3 0 2 7 9 1 9 9 14 13 3 0 2
19 1 15 9 1 0 9 12 1 11 13 12 9 2 16 13 1 9 9 2
21 13 4 2 16 9 0 9 14 4 13 9 1 9 7 0 9 0 1 0 9 2
34 14 2 3 15 3 13 1 15 13 2 7 16 9 1 0 7 0 9 14 0 10 9 13 9 9 2 13 10 10 9 14 3 0 2
35 1 0 9 11 11 1 0 9 15 13 12 9 0 7 0 9 2 10 0 9 7 4 3 13 10 9 0 9 2 15 4 11 3 13 2
6 9 4 13 14 0 2
20 1 0 9 1 9 4 13 3 7 14 1 0 9 4 1 9 1 9 13 2
21 9 2 1 15 15 4 13 0 0 9 2 13 12 0 7 3 0 1 0 9 2
12 10 9 4 13 1 10 9 0 9 7 9 2
7 0 9 14 4 13 9 2
17 4 13 13 10 9 2 7 4 13 1 9 0 1 9 7 9 2
31 3 16 0 9 7 9 2 16 4 15 13 2 16 4 13 9 7 13 10 9 2 4 13 1 10 9 0 9 14 9 2
48 16 3 16 9 9 0 0 9 4 1 15 13 10 9 10 9 2 4 13 10 9 3 0 1 10 9 0 9 7 9 2 1 15 4 13 2 16 4 15 1 9 13 1 9 0 0 9 2
37 1 9 7 9 10 9 15 3 3 13 14 1 0 9 2 16 13 11 7 0 9 2 16 3 16 0 9 13 16 9 7 14 4 13 0 9 2
11 0 9 4 13 2 16 0 9 13 9 2
11 1 0 0 9 13 9 9 9 0 9 2
37 1 11 4 13 0 9 1 0 9 1 9 11 11 2 16 4 12 12 9 3 13 2 16 4 13 1 9 0 9 7 3 13 0 1 0 9 2
11 10 9 13 14 1 0 9 1 0 9 2
15 11 2 11 7 11 13 0 2 7 14 13 10 0 9 2
14 16 4 1 9 13 0 9 2 13 13 9 7 9 2
13 9 7 0 9 4 13 0 1 9 7 9 0 2
19 7 9 7 9 4 13 13 3 0 2 14 16 4 13 0 13 0 9 2
8 9 13 9 9 1 9 12 2
10 1 10 9 13 9 9 3 0 9 2
13 16 9 4 14 9 13 1 9 7 13 1 9 2
12 0 1 10 9 1 9 13 9 7 9 13 2
12 9 2 16 13 10 9 2 9 13 1 9 2
34 15 13 14 0 9 9 2 16 9 2 16 4 13 1 9 2 4 9 13 9 2 16 15 14 13 13 7 16 4 3 13 10 9 2
10 11 4 1 0 9 13 1 0 9 2
7 7 9 16 15 13 0 2
18 1 15 13 0 9 2 7 1 15 13 9 2 9 7 0 9 9 2
14 1 9 4 12 2 9 13 3 1 12 2 0 9 2
15 9 11 2 11 11 11 2 4 9 12 13 11 7 11 2
13 1 9 11 13 0 9 3 0 3 1 9 9 2
11 16 9 13 1 0 9 2 13 0 9 2
8 0 9 13 3 0 9 9 2
14 9 11 15 3 3 13 9 1 0 7 0 9 9 2
10 3 13 0 9 11 0 9 12 9 2
13 9 9 11 15 13 14 2 16 9 1 9 13 2
24 3 16 13 0 9 1 9 11 3 0 9 2 13 0 9 1 9 11 0 7 3 3 0 2
12 13 1 9 9 9 7 0 9 1 0 9 2
11 9 4 1 9 11 13 1 9 7 9 2
22 1 9 1 9 13 0 9 7 15 15 4 13 9 2 16 15 4 13 1 0 9 2
25 1 15 3 9 1 0 9 1 9 13 1 0 9 2 1 15 7 1 9 14 13 14 9 9 2
21 11 4 1 0 9 7 3 1 9 11 13 9 9 11 1 9 11 2 11 9 2
30 9 2 16 4 9 1 11 9 9 1 11 3 13 2 15 4 13 2 11 13 14 11 9 7 11 9 1 11 2 2
20 16 13 13 9 11 2 3 13 0 9 1 10 0 9 7 0 9 1 9 2
15 1 0 9 15 13 1 3 10 9 2 16 4 15 13 2
12 3 4 10 9 13 2 3 4 0 9 13 2
24 7 3 2 16 4 3 0 13 1 10 9 2 15 15 4 3 13 2 3 15 13 1 9 2
10 3 15 4 13 1 0 9 7 13 2
8 14 7 3 13 3 0 9 2
8 0 7 13 14 1 0 9 2
8 3 13 14 10 16 12 9 2
15 14 13 2 3 13 14 10 0 9 3 0 9 1 9 2
31 1 15 13 14 0 0 9 7 9 2 7 16 15 3 3 13 1 10 16 12 0 9 2 1 15 0 13 14 12 9 2
13 1 15 15 4 15 13 2 15 4 13 0 13 2
17 7 3 4 1 0 0 9 2 16 15 3 13 2 3 13 0 2
12 0 13 1 11 2 13 15 14 1 0 9 2
11 0 9 11 11 13 14 3 3 1 9 2
13 1 0 9 1 9 1 9 1 11 4 13 9 2
7 9 4 13 0 7 0 2
18 13 15 4 1 10 0 9 2 15 15 13 1 9 7 13 1 9 2
21 11 4 13 1 9 16 9 9 2 7 15 4 1 9 13 7 13 0 0 9 2
27 9 4 1 15 13 1 9 2 15 7 14 13 13 1 0 9 2 15 0 9 4 1 9 13 1 9 2
14 9 2 16 13 9 0 9 2 13 0 7 14 0 2
10 3 1 11 15 13 0 7 0 9 2
13 0 9 13 13 11 11 1 9 1 9 0 9 2
23 10 9 1 9 13 14 0 2 7 14 0 2 7 4 1 9 13 9 7 14 0 9 2
23 1 0 9 7 4 13 0 2 7 15 4 13 3 3 2 16 4 3 7 3 3 13 2
24 15 3 15 4 3 13 1 10 0 0 9 2 7 4 14 1 0 9 13 1 9 15 0 2
33 16 9 1 0 9 14 4 13 13 1 10 9 2 13 9 14 1 0 9 3 0 2 15 13 2 16 13 13 0 14 10 9 2
25 7 1 10 9 14 14 4 13 1 9 2 1 15 15 13 1 9 2 14 7 4 13 0 9 2
6 0 9 4 13 9 2
16 9 2 16 4 14 3 13 2 13 0 1 9 1 0 9 2
15 0 9 2 1 15 9 9 14 13 13 2 7 13 9 2
15 11 4 13 0 2 16 11 3 14 4 13 9 1 9 2
20 9 1 9 13 3 0 0 9 3 1 9 7 1 2 3 7 3 15 13 2
6 3 15 4 13 15 2
12 16 16 14 4 14 13 9 2 1 15 13 2
21 10 9 9 4 13 1 9 1 11 2 9 7 4 13 1 0 9 1 9 9 2
7 3 15 4 3 13 9 2
13 9 4 3 13 0 2 16 16 4 13 0 9 2
5 11 4 14 13 2
7 3 15 4 13 0 9 2
9 15 13 9 2 16 13 1 11 2
10 11 11 4 1 0 9 3 13 9 2
11 1 9 4 15 13 0 9 2 3 13 2
4 15 13 9 2
10 13 4 1 9 7 13 1 0 9 2
10 11 15 4 13 1 9 9 1 9 2
10 1 10 9 4 13 0 9 9 11 2
13 1 10 9 4 13 1 9 3 0 9 0 9 2
16 1 9 4 13 9 2 16 15 4 3 13 1 9 0 9 2
24 11 4 10 9 13 2 16 13 2 7 15 4 13 11 2 14 16 4 3 13 1 0 9 2
12 4 15 13 13 2 16 4 13 3 14 14 2
14 13 4 2 15 15 15 13 13 2 16 4 13 13 2
7 1 9 15 4 11 13 2
7 13 4 1 10 9 9 2
11 11 4 13 0 15 2 16 4 13 9 2
21 11 4 13 9 7 13 11 11 2 16 13 1 15 7 15 1 9 13 1 9 2
6 11 15 4 3 13 2
7 2 14 2 2 4 13 2
6 10 9 4 13 9 2
9 14 7 15 13 3 3 11 11 2
3 13 15 2
6 13 4 0 7 0 2
9 13 15 4 2 16 15 15 13 2
15 9 4 13 1 11 2 16 4 13 9 0 1 0 9 2
5 9 4 13 14 2
8 10 9 4 15 13 1 11 2
14 11 4 3 13 7 9 9 15 15 4 13 1 9 2
17 13 15 4 1 11 11 2 7 15 15 4 14 13 1 0 9 2
9 9 1 15 4 13 9 11 11 2
17 0 13 3 0 7 13 14 0 2 7 14 1 15 13 0 9 2
7 0 1 15 13 11 11 2
14 9 13 0 9 7 4 13 1 9 0 9 7 9 2
15 1 0 9 1 9 0 9 0 0 9 4 13 13 9 2
26 13 4 15 15 14 9 7 9 2 16 4 1 10 9 13 1 0 0 9 7 13 13 9 7 9 2
24 16 4 9 13 1 9 2 4 15 1 0 9 13 9 2 0 9 2 9 7 0 0 9 2
16 0 0 0 9 13 0 1 0 2 0 9 1 9 1 9 2
32 0 0 9 2 9 2 0 1 0 9 2 0 1 9 2 9 2 9 2 9 2 9 2 9 7 9 2 13 0 0 9 2
11 10 9 4 1 9 13 9 7 13 9 2
29 9 15 4 3 13 1 9 2 7 9 15 4 13 7 9 15 4 1 10 9 2 1 9 7 9 13 1 9 2
24 9 9 14 4 13 1 10 10 0 9 2 7 4 3 13 0 7 3 13 10 9 1 9 2
19 1 11 7 1 9 4 1 0 9 1 0 9 13 14 0 9 7 9 2
33 9 14 1 10 9 14 4 13 15 16 3 2 7 4 1 9 13 9 2 9 2 0 0 9 2 16 4 15 15 13 1 9 2
28 15 15 4 13 1 0 9 2 4 13 13 14 0 9 7 9 2 16 4 1 0 9 9 13 1 0 9 2
12 1 9 4 9 1 0 9 13 12 9 9 2
30 9 13 9 2 16 4 10 0 9 1 0 9 13 0 9 0 9 7 13 9 2 16 4 15 13 1 10 0 9 2
14 1 0 9 13 3 9 9 2 16 13 9 7 9 2
8 11 9 4 14 14 3 13 2
19 7 7 4 1 0 9 9 13 13 2 7 4 13 9 0 9 7 9 2
20 13 4 2 16 4 9 13 0 0 9 2 16 13 3 1 9 1 0 9 2
19 16 9 4 13 2 16 4 15 13 1 0 9 2 4 15 13 14 9 2
24 16 1 0 9 9 4 13 9 1 9 2 4 9 13 3 13 1 10 9 7 13 10 9 2
11 0 9 11 9 4 3 13 9 0 9 2
13 1 0 9 4 13 0 14 13 9 7 13 9 2
14 9 4 15 13 13 1 9 2 16 15 4 9 13 2
12 3 4 0 9 13 14 9 0 9 7 9 2
10 3 7 15 4 9 13 3 1 9 2
17 13 4 1 9 7 1 9 7 3 4 13 1 9 3 0 9 2
15 1 0 0 9 13 9 9 2 9 2 9 7 0 9 2
6 3 4 13 3 3 2
12 13 15 4 2 3 7 15 3 13 1 9 2
25 11 4 13 10 9 1 9 2 16 4 13 14 0 2 3 16 4 0 11 13 12 9 1 11 2
18 9 1 9 15 4 3 13 2 7 4 13 11 13 1 9 7 9 2
10 1 9 4 13 1 9 14 1 9 2
19 2 13 15 2 15 15 4 13 2 16 4 15 13 3 2 2 4 13 2
8 13 2 15 15 13 1 9 2
3 13 9 2
11 3 4 13 2 16 15 14 4 13 3 2
17 1 9 4 13 9 2 16 4 3 13 7 13 9 9 1 15 2
13 3 15 14 13 13 2 11 9 13 3 1 9 2
26 3 15 13 13 1 0 9 2 7 0 9 9 2 16 4 13 0 9 10 9 2 4 15 3 13 2
7 16 1 9 15 14 13 2
15 11 4 14 13 1 9 7 9 4 3 13 9 1 9 2
12 9 4 14 3 13 9 2 3 15 4 13 2
6 13 4 7 15 13 2
8 9 13 13 3 2 1 9 2
14 13 4 11 1 0 9 1 9 2 13 9 7 13 2
34 7 9 13 3 0 7 0 2 10 0 9 2 9 9 11 1 0 0 9 7 10 9 1 3 0 11 2 3 13 14 1 0 9 2
23 0 9 1 0 9 9 7 0 9 4 13 1 9 9 2 4 7 3 13 1 10 9 2
27 9 1 9 11 11 4 13 3 2 0 9 9 7 4 13 0 7 0 9 11 11 1 9 0 9 11 2
18 11 11 4 13 0 7 0 11 2 11 11 11 7 4 13 10 11 2
16 1 9 11 7 9 11 4 15 13 9 11 11 7 11 11 2
28 1 9 14 3 13 0 9 2 9 7 0 9 2 7 13 3 0 14 9 0 9 7 9 1 10 0 9 2
10 7 0 16 0 13 1 3 0 9 2
30 3 14 13 1 0 14 12 9 0 0 9 11 11 2 0 1 0 0 9 1 9 2 9 1 15 13 9 0 9 2
40 3 13 1 0 9 3 0 9 2 3 16 9 1 9 9 1 0 0 9 13 0 9 2 16 15 3 13 7 0 0 9 16 9 9 2 9 7 0 9 2
36 15 13 0 9 2 15 15 4 3 13 1 9 14 3 0 9 9 1 12 7 12 9 11 11 7 0 9 1 9 9 9 1 9 11 11 2
23 14 11 11 4 13 2 16 4 10 9 14 13 3 3 1 11 2 3 1 3 0 9 2
14 11 4 10 9 3 3 13 2 16 4 13 0 9 2
15 9 4 13 14 14 12 2 16 15 4 9 13 1 9 2
7 14 3 15 4 11 13 2
18 15 15 4 13 7 7 15 15 4 3 1 10 9 3 13 15 0 2
6 13 15 4 7 13 2
6 3 7 13 15 0 2
18 9 1 9 13 14 1 11 0 2 7 16 13 10 9 0 7 0 2
9 3 9 13 9 9 1 0 9 2
31 1 3 0 9 4 15 13 3 13 14 0 9 9 9 2 7 7 10 9 13 0 1 9 9 9 1 0 9 11 11 2
18 13 10 9 2 16 4 10 12 9 3 13 2 15 15 1 15 13 2
20 14 2 15 4 1 0 13 11 2 13 1 10 9 7 16 13 0 2 2 2
3 2 8 2
22 1 15 15 1 10 0 9 13 11 11 2 9 12 9 0 0 9 11 11 1 11 2
25 1 11 13 0 2 16 15 9 14 4 3 13 2 7 0 9 9 13 3 0 1 9 1 9 2
20 11 4 1 9 1 11 13 2 16 11 0 7 0 9 1 11 13 0 9 2
43 7 13 13 14 2 16 15 4 11 13 10 0 9 2 16 14 3 13 9 1 11 2 7 3 14 13 13 0 9 1 9 1 9 2 15 4 13 0 0 9 11 11 2
10 15 2 15 13 2 14 3 14 13 2
13 9 14 14 13 7 15 1 0 9 4 3 13 2
6 15 15 14 4 13 2
20 13 4 14 12 15 2 16 4 15 13 1 9 12 9 2 16 4 13 9 2
7 15 4 1 9 13 3 2
22 1 11 4 1 0 9 0 14 13 9 2 7 4 15 3 13 2 16 15 13 11 2
15 1 10 9 14 4 13 13 1 9 14 1 0 0 9 2
12 3 15 15 4 13 2 7 13 3 0 9 2
9 9 1 9 13 1 15 0 9 2
15 1 15 7 13 14 9 15 2 16 1 9 3 3 13 2
21 9 4 3 13 0 9 2 1 15 3 15 13 2 3 13 1 15 9 10 9 2
18 16 4 1 10 0 9 13 1 14 2 3 13 3 1 9 1 9 2
10 1 11 11 4 1 11 11 13 0 9
25 9 2 10 13 11 2 15 3 1 9 10 9 1 0 9 3 0 9 13 14 3 0 9 9 2
27 1 9 10 9 0 0 9 1 11 4 13 0 9 9 2 16 14 3 13 10 14 9 7 0 0 9 2
19 0 9 11 2 15 9 14 15 14 13 2 13 0 1 9 7 0 9 2
38 10 0 2 9 9 2 4 11 1 9 13 1 0 9 2 1 15 15 4 13 1 0 9 1 14 3 0 9 1 9 9 11 2 9 1 9 2 2
38 0 1 9 7 0 9 1 11 4 13 3 13 2 16 13 9 14 2 1 9 2 2 16 15 13 1 0 9 2 13 7 16 15 15 0 14 4 2
12 9 0 9 13 1 9 1 9 0 9 9 2
24 1 0 9 15 1 0 9 2 0 9 2 13 0 9 2 16 15 0 0 9 13 0 9 2
29 9 13 3 3 14 1 9 0 9 2 7 7 13 1 9 1 0 9 2 16 13 9 7 9 9 1 0 9 2
27 9 0 9 13 3 9 0 0 9 1 0 9 2 9 7 9 0 9 2 9 0 9 2 0 0 9 2
12 12 3 0 9 1 9 1 9 13 0 9 2
23 3 3 1 9 15 9 13 1 0 7 0 9 7 13 9 2 16 15 1 9 9 13 2
17 3 7 3 13 3 0 15 2 3 0 9 0 9 9 1 15 2
24 3 0 7 0 13 9 2 16 15 3 13 9 1 9 7 14 9 2 16 13 9 1 9 2
16 1 9 13 9 2 9 2 1 9 2 3 15 13 14 9 2
7 0 9 3 13 7 13 2
14 10 10 9 3 13 1 9 1 9 2 3 0 9 2
19 9 1 0 9 13 0 9 9 7 0 9 2 9 7 0 9 9 2 2
26 9 10 9 1 9 13 0 1 0 9 2 9 2 8 8 13 10 9 16 8 8 2 7 1 9 2
10 0 9 7 9 13 9 9 1 9 2
17 0 0 9 13 0 9 1 9 9 9 9 7 9 7 0 9 2
8 9 10 9 13 3 10 9 2
44 0 0 9 13 2 16 14 4 0 0 9 13 12 1 12 9 0 0 9 9 2 16 15 13 1 12 9 2 1 9 2 9 7 0 9 7 14 4 13 10 9 12 9 2
20 0 9 7 9 2 8 8 2 13 0 9 2 16 15 3 13 1 9 9 2
17 1 9 13 9 2 8 8 2 2 9 7 13 0 14 10 9 2
11 9 13 14 3 0 2 1 15 0 9 2
9 9 13 1 9 1 3 0 9 2
20 0 9 13 0 9 2 1 9 7 1 0 9 13 0 9 2 16 3 13 2
8 3 4 10 9 14 13 9 2
17 3 13 2 16 1 9 3 13 9 1 9 1 9 1 0 9 2
10 0 9 4 13 14 1 10 0 9 2
18 13 4 2 16 9 1 9 1 9 2 9 1 9 2 13 9 9 2
13 1 15 7 15 4 1 0 9 13 14 0 9 2
17 1 0 9 4 13 14 9 2 9 1 0 9 2 7 0 9 2
11 1 0 9 3 13 0 9 9 1 9 2
28 13 4 14 2 16 4 9 9 13 9 9 2 3 3 0 7 0 9 9 2 2 7 13 2 16 13 3 2
9 9 1 9 3 13 1 12 9 2
22 0 9 2 0 9 2 9 7 0 9 13 3 0 7 3 13 0 9 9 1 9 2
13 13 15 13 14 0 9 7 1 0 2 0 9 2
23 13 2 16 13 10 9 13 3 7 16 13 1 9 7 9 0 2 7 16 9 13 3 2
19 9 13 14 1 0 9 2 7 1 3 14 4 13 0 0 9 1 9 2
7 13 14 0 7 0 9 2
7 9 13 1 9 1 9 2
26 1 9 0 9 0 9 7 9 3 1 9 9 3 13 7 13 9 2 16 4 3 13 9 9 9 2
6 7 9 13 0 9 2
19 3 13 0 2 16 9 13 9 2 16 13 14 0 2 0 9 1 9 2
11 1 9 9 13 3 12 1 12 9 9 2
14 1 11 15 13 1 0 9 7 0 9 10 12 9 2
16 10 9 13 9 2 7 0 9 14 13 13 9 1 0 9 2
27 9 2 16 13 9 1 15 13 2 15 3 13 9 7 13 9 1 0 9 2 16 15 15 13 1 9 2
26 9 2 16 15 13 1 9 2 13 1 9 0 9 2 16 13 9 1 0 9 7 13 9 9 15 2
9 10 9 13 0 13 1 0 9 2
13 16 13 9 14 3 1 9 2 13 0 9 9 2
17 16 13 1 0 9 2 13 9 13 13 9 2 16 4 13 9 2
7 13 9 1 0 9 0 2
21 7 1 10 0 0 9 3 13 9 0 9 9 1 9 7 1 15 9 0 9 2
23 10 9 14 3 13 0 2 7 4 3 13 2 16 0 9 13 9 9 2 0 9 2 2
20 0 9 1 3 0 9 7 13 9 9 2 3 16 3 3 13 1 9 9 2
26 13 2 16 3 13 1 10 9 0 9 1 0 9 2 1 15 7 14 13 13 1 9 0 9 9 2
53 1 9 1 9 9 7 9 9 1 9 0 9 7 15 9 9 13 1 9 9 9 12 2 0 9 2 7 9 12 2 0 9 2 9 7 0 9 3 0 9 12 9 2 0 9 2 7 0 9 2 9 2 2
23 16 0 9 7 13 0 2 4 13 0 9 1 9 1 9 9 1 9 2 9 7 9 2
20 9 1 9 0 9 4 0 9 1 10 9 13 2 16 4 3 13 0 9 2
20 3 13 9 1 9 0 0 9 4 1 9 0 0 9 0 9 3 13 9 2
24 0 9 4 13 1 0 9 2 1 15 4 0 9 13 3 2 3 7 4 13 14 10 9 2
30 16 4 15 1 0 9 13 2 16 13 0 3 13 14 0 0 9 9 2 4 15 13 0 9 1 9 9 0 9 2
25 9 2 16 15 1 9 13 1 9 2 4 1 9 9 13 0 9 7 15 3 13 3 1 9 2
22 9 4 13 14 0 1 9 1 0 9 9 2 7 9 2 16 14 4 13 13 9 2
8 9 9 13 14 0 9 0 2
11 16 9 13 2 13 9 10 9 7 15 2
22 9 4 13 9 7 9 10 9 2 16 4 15 13 1 9 9 1 9 1 11 11 2
11 9 13 12 9 0 9 1 0 0 9 2
17 1 0 9 13 0 9 1 0 9 2 16 16 9 13 9 3 2
10 9 1 12 0 9 13 3 0 9 2
31 14 16 4 15 15 13 2 4 15 13 1 0 9 2 0 9 2 16 13 9 1 0 9 2 15 14 4 13 3 13 2
17 15 13 3 3 2 16 16 4 15 3 1 3 13 9 0 9 2
17 9 2 16 15 13 1 12 0 0 9 2 13 1 9 0 9 2
6 10 9 13 9 12 2
22 15 13 2 16 4 13 13 0 9 9 2 16 13 0 9 2 0 9 7 9 9 2
19 14 3 7 9 9 13 1 0 9 2 16 13 9 2 9 7 0 9 2
26 0 9 13 0 9 9 2 7 13 1 10 0 9 0 9 0 9 9 12 7 9 12 7 0 9 2
28 16 13 9 9 9 7 9 14 1 9 9 9 2 13 14 9 1 9 1 9 7 0 9 7 9 16 9 2
22 1 15 15 13 0 9 9 1 9 7 0 9 2 16 13 15 9 1 0 10 9 2
3 2 13 2
15 13 2 2 15 4 14 3 13 11 7 13 9 1 9 2
9 9 4 13 0 1 0 0 9 2
10 9 4 1 10 9 14 3 13 9 2
5 0 2 0 9 2
9 9 1 15 4 13 3 0 9 2
10 0 9 9 4 13 7 3 1 9 2
18 1 9 0 9 4 9 9 13 7 1 9 16 1 9 7 0 9 2
25 9 4 1 10 9 14 13 0 9 2 7 7 4 13 3 10 9 2 16 4 15 14 3 13 2
6 0 9 4 13 0 2
7 0 9 4 13 14 0 2
19 1 15 1 0 9 14 4 13 15 14 2 16 4 3 13 14 10 9 2
23 2 13 14 12 9 2 2 4 13 9 2 16 15 4 3 13 7 3 3 13 1 9 2
23 11 15 4 13 2 3 4 13 9 14 3 0 2 16 4 13 2 16 13 10 9 0 2
15 2 15 13 3 3 2 2 4 1 0 9 13 11 11 2
22 0 9 4 3 13 9 0 9 7 3 13 10 9 3 1 9 0 0 7 0 9 2
40 1 15 4 13 9 1 9 9 7 1 0 0 9 2 16 4 13 0 1 10 9 2 0 7 0 2 7 9 2 1 0 9 2 3 4 13 10 0 9 2
11 3 4 9 0 9 1 0 9 3 13 2
18 1 9 12 9 4 0 9 13 9 0 9 2 9 0 9 7 0 2
20 3 15 4 0 9 1 9 0 9 13 7 13 15 4 9 0 9 10 9 2
17 1 12 9 15 13 0 1 12 9 2 16 15 13 1 0 9 2
23 16 15 13 1 11 11 11 9 2 13 14 9 1 12 7 12 9 2 16 13 1 9 2
12 14 0 9 15 13 14 1 0 9 1 9 2
30 9 11 11 13 1 10 0 9 0 2 7 14 13 0 9 9 1 9 11 2 16 15 13 0 13 12 9 2 9 2
27 1 9 2 16 4 13 0 2 4 13 14 0 13 3 0 9 2 7 4 13 9 0 1 3 0 9 2
28 16 4 11 13 0 9 7 13 0 0 9 2 4 10 9 2 9 7 14 9 3 1 9 13 9 10 9 2
12 3 4 15 14 1 0 9 13 13 0 9 2
12 0 9 13 0 9 2 16 4 13 1 15 2
22 10 9 13 3 0 2 16 4 13 10 9 1 9 2 7 7 4 15 3 3 13 2
44 3 1 9 9 1 11 7 1 9 9 11 13 10 9 1 0 9 2 16 13 9 2 16 13 9 2 0 2 1 15 15 0 9 13 2 14 16 13 9 2 9 7 9 2
24 0 9 4 13 2 16 9 3 3 13 0 9 2 15 13 0 9 0 7 0 9 0 9 2
21 2 15 2 16 9 1 10 9 13 3 2 13 0 1 10 9 2 2 13 11 2
16 0 9 1 9 13 9 2 16 13 9 1 0 7 0 9 2
15 14 9 13 13 9 1 0 9 2 2 7 9 14 13 2
15 11 13 2 16 13 0 9 0 14 1 9 0 9 9 2
41 1 0 9 2 1 15 15 13 1 9 2 0 9 13 9 0 9 2 16 0 9 13 9 7 9 2 7 9 2 0 9 2 16 1 9 1 0 13 0 9 2
6 15 14 13 3 3 2
22 3 1 11 4 13 13 9 9 1 9 2 7 15 0 0 9 1 15 4 3 13 2
15 1 0 9 4 0 9 3 13 7 9 4 13 14 0 2
6 7 4 9 3 13 2
15 1 0 9 4 13 8 11 2 16 4 13 9 1 11 2
30 13 2 16 1 9 1 9 4 13 0 9 1 9 2 7 1 10 9 13 1 0 10 0 9 2 16 13 9 9 2
16 3 15 14 13 0 9 14 0 9 2 16 14 13 0 9 2
14 9 9 1 0 0 9 4 1 9 13 0 9 9 2
8 0 9 13 7 3 0 9 2
12 3 0 0 9 9 13 9 2 9 7 9 2
11 1 9 9 11 12 4 13 14 12 9 2
17 1 15 15 10 0 0 0 0 9 14 3 13 1 9 1 11 2
32 1 9 9 12 4 11 1 9 9 1 9 12 9 1 0 9 11 13 9 0 9 2 16 15 13 10 12 9 9 1 11 2
15 3 4 13 0 2 16 4 11 12 13 1 3 0 9 2
35 1 9 10 9 4 13 2 16 4 14 10 12 9 13 9 11 2 1 9 1 9 7 4 9 13 9 2 16 15 1 0 9 13 9 2
11 10 0 9 1 15 14 3 9 14 13 2
19 16 1 9 4 0 9 1 9 7 11 13 9 1 9 9 1 0 11 2
31 11 13 0 1 9 2 16 4 13 9 9 7 9 9 1 9 1 9 2 1 15 7 4 0 13 0 9 9 7 9 2
15 13 4 14 2 16 9 1 0 9 13 14 0 9 9 2
8 9 9 13 7 0 7 0 2
45 0 9 15 13 9 2 16 4 1 9 12 10 9 3 3 13 1 0 9 2 3 4 7 11 1 9 10 0 9 2 0 9 7 1 0 9 9 3 0 9 13 10 0 9 2
34 3 7 15 13 3 2 16 1 10 9 1 12 9 2 16 13 2 4 9 3 13 10 2 0 9 2 10 9 2 7 9 0 9 2
16 1 9 15 9 14 14 3 13 2 10 0 9 7 13 0 2
12 9 1 9 1 9 0 9 13 0 0 9 2
21 13 15 2 16 3 9 1 9 3 13 1 9 2 16 4 13 14 1 0 0 2
30 0 9 15 13 1 0 0 9 1 0 9 2 0 1 9 1 9 3 0 9 0 0 0 9 7 0 0 9 9 2
18 9 4 13 0 9 1 10 9 2 16 15 13 9 12 0 9 9 2
12 10 0 9 4 13 16 0 0 1 0 9 2
8 3 15 4 13 14 10 9 2
11 15 4 13 7 15 4 13 9 1 9 2
13 1 10 9 13 9 0 9 12 9 7 12 9 2
19 15 13 3 15 9 2 16 15 13 0 9 2 16 13 1 9 12 9 2
28 0 9 1 9 13 13 1 12 7 1 12 0 9 0 9 7 12 2 2 12 9 9 1 9 0 0 9 2
29 13 13 14 3 0 0 9 2 16 13 0 9 9 2 16 15 13 1 0 9 9 13 1 12 2 2 12 9 2
22 3 16 1 0 9 13 0 9 2 13 1 0 9 0 9 1 0 9 2 0 9 2
7 9 10 9 13 12 9 2
26 0 9 2 16 13 3 0 1 9 1 9 0 9 2 13 3 12 0 0 9 1 0 7 0 9 2
13 1 10 9 13 1 0 0 9 0 3 9 9 2
18 2 3 2 16 4 1 10 9 1 9 13 9 2 2 4 13 11 2
21 16 0 9 1 0 9 13 2 10 0 9 3 1 0 0 9 13 9 0 9 2
21 9 9 13 1 0 0 9 0 9 2 16 15 13 1 9 1 0 9 0 9 2
21 9 2 16 15 1 0 9 13 0 0 9 2 13 16 0 9 1 0 9 9 2
27 16 13 0 0 9 0 2 0 9 14 13 13 0 9 0 9 1 0 9 2 15 15 3 13 16 9 2
15 0 13 9 0 9 9 2 0 0 9 2 8 11 2 2
26 3 4 9 13 9 1 15 2 15 4 15 13 1 9 2 13 9 7 9 2 16 4 14 15 13 2
10 0 9 13 14 0 7 15 14 13 2
13 0 9 2 3 3 15 13 7 14 13 13 9 2
8 10 0 9 13 0 7 0 2
7 13 4 15 14 0 9 2
32 14 1 0 9 4 11 1 11 13 10 9 2 0 0 9 0 9 3 3 1 9 13 1 15 2 16 15 1 15 13 11 2
8 11 1 11 4 13 14 3 2
10 1 15 14 4 14 13 14 0 9 2
36 10 9 1 0 9 15 15 3 13 3 0 2 1 9 9 7 4 13 0 0 9 10 0 7 0 9 2 16 15 3 4 13 3 3 13 2
25 14 3 4 11 1 10 0 9 13 15 2 15 13 0 7 0 2 1 9 9 9 13 1 15 2
21 9 3 3 13 3 3 1 10 9 2 7 14 15 4 0 15 11 13 1 15 2
10 0 9 15 4 13 0 1 0 9 2
26 16 11 2 16 13 3 0 14 1 0 9 2 13 1 9 2 4 3 3 0 1 15 13 3 15 2
8 9 15 15 14 4 13 13 2
12 2 14 2 3 13 2 2 4 13 11 11 2
19 3 4 13 1 0 9 7 11 4 13 0 0 9 1 9 7 13 13 2
47 11 15 4 14 3 13 3 7 1 15 2 16 15 4 9 13 9 2 1 9 13 0 0 9 2 0 9 2 0 2 0 9 7 0 2 0 9 2 16 15 4 13 1 0 0 9 2
18 13 4 0 9 7 13 4 13 14 9 9 2 16 15 4 13 11 2
22 1 0 9 4 13 0 9 2 1 9 7 15 4 13 9 2 16 15 4 13 9 2
4 11 4 13 2
10 3 3 7 3 15 4 13 9 9 2
8 9 13 14 3 0 9 9 2
29 0 9 1 15 13 1 15 2 16 13 1 9 0 9 2 16 13 0 7 0 9 2 9 1 0 0 9 2 2
6 15 13 9 7 9 2
11 16 13 2 13 0 9 0 9 3 0 2
24 1 9 13 2 16 13 0 0 9 3 3 16 0 1 9 0 9 9 7 9 1 0 9 2
7 9 7 13 3 0 9 2
18 13 15 9 0 9 7 13 15 0 9 7 9 2 16 13 10 9 2
22 15 13 2 16 3 0 9 3 13 1 10 9 7 16 15 1 15 1 0 13 9 2
21 1 3 0 0 9 13 14 3 0 13 2 16 15 4 10 9 3 13 3 3 2
14 0 9 1 0 9 13 14 1 9 7 9 1 9 2
20 15 7 13 1 0 9 2 16 13 9 1 0 9 3 0 2 3 0 9 2
15 15 1 0 9 3 13 7 1 9 9 13 2 16 13 2
19 4 14 13 0 9 0 9 7 9 1 9 1 0 9 13 3 0 9 2
16 0 9 11 11 13 0 2 16 1 0 9 13 9 0 9 2
22 1 15 4 14 0 0 9 11 11 13 2 16 15 4 9 1 0 9 1 11 13 2
15 0 11 13 3 13 14 10 9 2 16 4 3 13 9 2
26 11 1 9 9 9 2 16 4 13 1 9 1 9 1 9 9 9 2 4 3 13 1 0 9 9 2
51 1 0 9 7 9 2 15 9 13 10 9 1 9 9 1 9 0 9 7 9 9 1 0 9 2 4 15 9 1 9 0 9 13 14 1 9 2 4 1 0 9 13 11 11 2 9 0 9 1 9 2
15 1 0 9 13 1 9 1 9 0 9 0 12 9 9 2
16 15 13 3 14 1 9 9 0 9 2 1 15 4 13 9 2
11 1 0 9 9 13 3 10 16 9 9 2
19 3 0 9 9 9 13 1 3 0 0 9 2 16 4 15 16 14 13 2
8 14 0 9 15 14 13 13 2
6 9 13 14 1 9 2
7 0 9 13 0 1 9 2
34 10 0 9 11 11 4 13 10 0 9 14 1 0 9 11 11 2 16 15 4 13 13 9 2 1 15 4 0 9 13 14 10 9 2
26 3 4 1 10 0 9 13 9 9 11 11 2 3 16 15 4 3 13 1 9 0 0 7 0 9 2
18 11 11 13 2 16 4 13 3 13 9 1 9 1 0 7 0 9 2
16 9 1 15 15 1 15 13 1 9 7 9 0 9 1 0 2
31 10 9 4 1 9 0 0 9 0 9 4 13 0 9 9 11 11 2 16 4 1 11 13 9 1 9 9 1 0 9 2
21 13 4 2 16 2 13 15 13 9 2 7 9 14 13 13 1 9 0 9 2 2
39 2 16 3 14 13 9 1 9 0 9 2 4 10 9 13 13 0 9 2 2 4 13 0 9 2 0 2 16 15 4 13 0 9 1 0 9 11 11 2
9 2 14 2 2 4 13 1 9 2
14 2 9 15 13 1 9 1 9 2 16 13 1 9 2
12 3 13 10 0 9 1 10 9 7 13 9 2
16 16 13 1 15 2 3 13 9 2 13 10 9 7 0 9 2
8 13 15 0 9 7 15 13 2
26 1 9 9 4 13 2 16 13 9 0 0 9 2 16 2 13 11 1 15 2 16 15 13 13 2 2
24 1 0 9 2 1 15 4 13 14 9 9 9 2 4 3 1 12 9 9 13 1 9 9 2
28 14 1 0 0 9 15 1 9 11 3 14 3 13 2 0 9 7 15 4 13 14 9 0 9 1 0 9 2
33 1 9 0 9 7 0 9 4 0 9 13 14 1 9 2 1 12 9 9 2 1 15 7 4 9 13 14 1 9 7 9 9 2
20 3 4 13 1 9 11 7 11 1 11 2 16 4 13 9 12 0 0 9 2
12 13 4 0 9 9 7 4 10 9 13 9 2
16 11 4 13 1 0 9 13 9 7 9 2 16 15 3 13 2
13 16 4 15 13 1 15 2 4 9 13 0 9 2
34 9 4 13 1 9 0 9 2 16 4 13 1 9 2 7 16 4 13 2 16 4 13 1 9 7 15 13 2 1 0 9 1 9 2
14 16 13 15 9 1 9 2 4 13 15 15 3 0 2
9 7 4 15 13 0 9 1 9 2
20 16 1 0 9 15 4 13 0 13 2 15 4 11 13 2 16 15 4 13 2
15 7 14 15 15 13 2 16 0 9 1 9 14 13 13 2
9 1 0 15 13 2 9 13 9 2
18 7 1 9 3 14 13 9 2 0 9 2 7 14 13 14 0 9 2
19 16 15 4 13 0 7 0 0 9 7 10 9 9 2 15 4 9 13 2
32 16 13 3 1 10 0 9 2 15 4 13 15 2 16 14 4 13 1 9 2 16 4 15 1 0 9 13 3 1 10 9 2
6 13 15 4 1 9 2
25 1 0 0 9 13 0 9 9 1 9 2 7 4 9 1 10 9 13 9 14 1 0 9 9 2
22 3 1 9 0 9 7 15 4 14 1 9 9 13 13 1 9 9 1 9 9 9 2
27 1 15 4 1 0 9 3 13 14 1 9 10 9 2 16 1 0 9 13 10 0 9 16 15 13 9 2
29 14 13 14 15 0 2 16 1 10 9 13 0 14 10 9 2 16 4 13 1 10 9 14 0 2 0 7 0 2
20 7 3 13 1 0 9 2 9 13 9 2 16 4 15 0 9 13 1 9 2
12 0 0 9 4 13 1 9 12 9 7 12 9
9 2 3 13 2 16 15 13 3 2
56 11 13 3 14 3 0 2 16 3 13 2 3 9 13 7 15 13 1 9 2 2 13 11 11 2 16 4 13 14 2 16 4 13 9 2 16 11 4 13 7 16 4 13 9 9 7 0 9 0 2 1 15 0 0 9 2
10 2 13 15 3 2 16 4 3 13 2
21 0 4 13 14 0 9 1 9 1 9 12 2 3 16 4 1 0 9 13 3 2
25 1 11 4 13 14 1 0 9 2 1 11 2 16 4 13 0 9 2 15 4 13 1 0 9 2
18 15 13 14 0 9 0 1 2 9 9 2 1 11 7 9 0 9 2
18 11 4 13 14 0 9 1 11 7 10 10 9 2 16 13 0 9 2
8 13 1 10 10 9 1 9 2
19 13 13 1 9 7 0 9 2 7 13 1 9 7 15 1 0 9 13 2
11 13 2 16 4 9 9 3 13 10 9 2
8 3 15 4 13 1 0 13 2
4 13 1 3 2
5 15 15 3 13 2
9 3 4 15 13 1 11 2 11 2
16 13 9 0 0 9 2 1 9 12 4 13 10 9 11 11 2
10 3 15 4 13 13 9 1 9 9 2
13 14 2 15 13 9 2 16 4 13 0 1 11 2
12 13 4 0 9 1 0 9 7 1 10 9 2
15 3 4 13 1 9 9 2 9 2 9 2 9 2 2 2
9 10 9 4 13 0 9 7 9 2
16 3 4 13 2 3 15 3 13 2 7 4 15 13 3 13 2
21 13 15 2 3 4 13 1 9 1 11 7 11 1 10 9 2 0 1 10 9 2
9 2 15 13 9 7 9 1 9 2
9 1 11 13 13 2 2 4 13 2
21 3 15 4 13 2 16 4 13 9 2 16 4 0 9 11 13 9 1 9 9 2
10 13 4 3 0 2 7 13 4 15 2
9 0 0 9 4 13 1 12 9 2
33 0 0 9 11 2 16 13 1 0 0 0 9 0 9 7 15 13 1 9 0 2 14 12 2 0 9 2 13 14 1 0 9 2
18 9 13 0 13 1 9 1 9 7 0 9 2 15 3 14 3 13 2
13 7 15 3 14 3 13 14 1 3 0 0 9 2
17 15 15 13 1 0 9 2 10 9 7 13 1 9 0 0 9 2
13 14 13 0 2 16 15 2 15 9 13 2 13 2
35 3 13 9 1 9 10 0 9 7 14 1 15 2 10 9 13 1 15 1 10 0 9 2 0 9 1 9 1 15 2 15 13 0 9 2
26 9 3 13 14 2 16 13 14 3 3 13 1 9 9 7 1 15 2 15 3 13 1 9 0 9 2
17 14 1 0 9 0 9 14 3 15 1 12 9 4 13 1 0 2
37 0 9 15 4 3 13 1 9 0 9 2 3 7 4 13 9 0 9 2 16 4 3 13 0 9 0 9 2 16 4 13 0 1 10 10 9 2
24 1 15 4 15 1 9 13 3 0 9 9 1 9 7 4 13 9 1 10 9 13 10 9 2
9 7 3 4 13 0 9 1 9 2
11 3 15 13 13 1 0 9 1 9 9 2
30 16 13 13 10 9 2 15 15 15 13 10 0 7 0 9 2 13 3 13 2 15 10 9 13 7 1 15 13 0 2
26 1 15 7 13 13 9 9 2 7 16 4 3 13 9 10 0 9 7 3 10 0 9 1 12 9 2
25 16 4 13 2 10 13 0 9 2 15 13 13 1 9 2 14 16 4 13 9 2 16 4 13 2
14 15 13 0 9 2 16 9 13 14 9 7 3 13 2
26 13 15 13 0 9 7 13 1 3 0 9 9 2 16 13 15 10 9 7 9 7 9 7 14 9 2
10 15 15 4 14 13 16 9 1 9 2
32 7 13 0 2 16 13 3 9 1 15 2 16 13 2 16 4 13 3 3 0 7 0 9 2 16 13 15 2 1 15 13 2
7 13 15 9 10 9 9 2
20 16 15 13 2 16 15 9 13 9 2 7 15 13 2 16 13 1 0 9 2
9 15 13 9 1 15 1 10 9 2
17 7 7 13 15 3 0 9 1 9 9 7 15 14 13 13 0 2
11 3 3 13 15 15 2 16 13 0 9 2
17 3 13 0 9 0 2 0 9 1 9 2 16 15 13 13 3 2
17 3 9 0 0 9 13 1 15 2 16 13 10 9 7 10 9 2
17 1 10 9 15 0 9 7 9 9 13 2 16 3 13 0 9 2
21 0 0 9 2 1 15 13 9 2 13 14 9 0 9 7 0 9 0 0 9 2
25 16 10 0 9 13 7 14 15 10 0 9 2 9 2 2 9 2 9 2 7 9 2 9 2 2
51 10 9 4 1 9 1 3 0 0 12 9 7 1 9 2 16 4 13 0 12 9 2 13 1 0 9 2 1 15 13 14 3 2 7 1 15 4 13 1 1 9 12 2 16 3 13 9 0 0 9 2
5 3 15 13 13 2
7 9 13 3 13 16 13 2
20 7 14 9 1 9 2 1 9 13 10 9 0 9 0 1 12 1 12 9 2
25 3 4 14 13 1 9 1 9 10 0 9 2 7 9 15 15 7 13 3 0 2 0 2 0 2
39 13 7 15 2 16 15 1 10 9 3 3 13 10 9 7 10 10 9 1 9 2 16 13 0 1 9 7 9 15 2 15 4 3 3 14 1 3 13 2
18 0 13 11 11 2 0 9 7 9 1 9 1 9 2 1 0 9 2
12 9 4 13 14 0 2 15 4 11 3 13 2
29 1 9 4 13 3 0 9 2 10 9 1 9 0 9 7 0 9 2 1 15 15 4 13 13 15 1 10 9 2
9 9 4 13 2 14 16 4 13 2
8 13 1 11 4 13 0 9 2
10 3 4 13 1 0 9 7 13 9 2
18 0 4 13 2 16 15 9 3 13 9 2 7 13 4 0 0 9 2
12 14 16 15 4 2 13 2 9 1 0 9 2
15 8 11 11 4 13 11 1 0 0 9 1 10 0 9 2
21 3 15 4 13 2 15 4 13 1 11 11 0 2 0 2 3 3 0 0 9 2
9 11 11 4 13 9 7 15 13 2
9 0 13 2 16 4 13 14 0 2
6 13 13 2 4 13 2
9 3 3 4 13 9 1 10 9 2
10 3 3 4 13 10 9 1 11 9 2
26 1 12 9 4 13 10 9 3 0 2 4 13 11 11 2 16 4 13 0 9 2 16 4 13 3 2
18 16 15 4 11 11 1 9 3 13 2 15 4 13 2 16 13 0 2
24 3 15 4 13 10 9 7 13 4 13 2 16 11 14 13 1 9 2 16 4 13 11 11 2
26 14 10 9 4 13 0 2 7 16 4 13 11 1 9 2 4 3 3 13 2 16 4 15 3 13 2
19 3 15 4 13 2 16 14 4 13 1 9 2 16 4 3 13 0 9 2
28 9 2 16 15 4 0 9 13 1 0 9 2 10 4 13 11 2 4 13 12 10 0 9 2 16 4 13 2
39 13 15 4 2 16 4 13 9 2 16 4 15 13 1 9 1 9 2 7 9 2 16 4 13 1 10 9 2 7 13 15 4 2 16 4 13 10 9 2
5 13 4 1 9 2
25 9 1 0 4 13 1 0 9 2 7 11 4 13 0 0 9 7 13 9 2 16 15 4 13 2
16 11 4 1 9 13 9 2 16 4 13 1 9 1 9 9 2
15 3 16 4 13 2 16 13 11 0 2 15 4 13 9 2
26 9 4 13 3 0 7 9 4 13 1 9 2 7 4 13 0 9 1 15 2 16 4 13 13 0 2
10 15 15 4 13 2 15 4 13 11 2
11 13 2 16 13 3 3 2 4 13 11 2
10 3 4 13 1 15 2 16 4 13 2
24 3 4 15 13 2 16 14 13 13 7 13 2 15 15 13 2 7 3 4 13 0 1 15 2
15 16 4 13 9 2 13 2 16 13 2 16 13 1 15 2
10 13 15 13 1 9 2 16 4 13 2
19 3 15 4 13 2 3 16 4 13 2 16 13 3 0 7 14 3 0 2
15 13 4 1 9 1 0 9 2 16 15 4 13 10 9 2
15 3 4 15 13 14 13 2 16 13 10 0 9 3 9 2
38 11 4 3 13 1 11 11 7 15 13 2 16 4 13 0 9 2 16 15 4 13 1 15 2 16 15 4 13 1 9 9 2 10 0 9 1 11 2
9 2 13 15 2 2 4 3 13 2
