1798 11
10 11 7 2 10 12 9 10 13 4 2
8 11 9 9 3 13 4 11 2
13 15 9 2 9 12 2 9 10 2 3 13 4 2
7 12 9 13 4 9 13 2
11 3 13 4 9 0 3 13 4 9 13 2
7 11 9 0 13 13 4 2
7 0 9 9 0 13 4 2
10 7 2 13 7 3 13 4 13 4 2
19 9 10 2 11 7 11 9 13 4 13 4 2 7 3 9 13 4 11 2
10 9 13 2 11 14 13 10 0 0 2
12 3 2 11 3 13 11 9 7 13 4 11 2
15 12 9 10 11 7 11 9 0 7 0 13 4 9 9 2
23 15 9 9 13 2 7 10 13 13 9 2 7 9 0 12 7 13 2 9 13 4 13 2
15 10 2 7 2 9 13 4 9 11 11 13 4 9 0 2
5 7 2 13 9 2
6 3 14 4 13 9 2
11 9 9 2 0 7 0 13 13 4 9 2
8 3 9 9 13 4 9 9 2
7 9 13 3 13 4 9 2
19 12 2 7 2 11 9 13 4 2 11 9 2 11 13 9 9 9 13 2
14 7 2 13 13 4 15 13 9 2 3 0 2 13 2
20 9 2 9 0 9 9 9 0 13 7 0 13 4 3 13 2 3 13 13 2
13 11 10 9 13 9 9 13 4 9 0 13 4 2
5 10 9 13 4 2
17 9 0 13 2 7 9 12 13 9 4 9 12 13 13 9 13 2
21 10 3 3 13 4 2 10 10 9 13 7 0 2 15 9 13 2 3 13 4 2
15 9 0 11 9 9 9 13 4 9 7 9 0 13 4 2
10 11 9 13 9 13 11 9 11 9 2
16 11 2 8 11 2 11 2 11 7 11 7 9 13 13 3 2
13 14 4 13 13 4 2 7 3 13 13 4 9 2
10 2 9 9 13 4 7 9 0 13 2
12 9 10 9 0 13 7 13 3 0 13 4 2
8 11 7 14 13 3 9 13 2
5 13 4 13 4 2
10 9 13 7 14 2 9 0 13 4 2
8 9 0 13 4 9 0 7 2
8 3 2 11 7 11 13 4 2
16 11 13 13 9 0 13 4 9 2 2 15 9 14 13 2 2
11 3 12 9 0 13 4 9 11 7 11 2
6 2 9 0 13 3 2
7 2 9 10 13 9 13 2
25 3 13 7 9 13 9 14 4 13 2 13 3 2 10 10 13 4 10 9 11 9 0 7 0 2
11 9 10 13 4 2 14 4 15 9 13 2
8 9 0 13 4 9 7 9 2
11 11 9 13 13 7 13 13 9 13 4 2
23 7 2 9 13 9 13 9 11 10 9 13 4 2 11 9 14 4 10 13 9 10 13 2
6 9 9 13 13 4 2
16 9 9 13 2 9 9 13 3 11 2 12 2 11 11 9 2
11 2 11 13 13 4 2 9 13 3 2 2
3 9 13 2
11 12 9 9 13 2 7 3 9 10 13 2
5 11 13 4 12 2
16 3 2 3 2 3 7 3 13 4 7 2 9 12 13 9 2
11 0 13 4 11 7 11 9 10 10 9 2
13 9 0 13 2 7 9 3 13 10 13 9 13 2
8 3 3 13 9 2 9 13 2
9 11 12 9 9 13 4 9 0 2
6 11 7 3 13 4 2
14 2 7 9 10 0 13 9 9 9 13 9 13 2 2
13 11 9 10 9 13 4 11 9 7 9 13 4 2
11 9 13 4 12 9 9 13 3 2 0 2
15 7 15 9 13 10 14 13 9 2 7 13 9 13 4 2
5 2 14 13 9 2
12 12 9 3 13 4 2 7 14 4 9 13 2
5 9 0 13 4 2
11 11 7 11 13 13 3 2 11 13 4 2
13 7 2 9 2 9 7 9 9 0 0 13 3 2
9 0 2 10 9 13 9 13 13 2
8 10 13 9 3 13 4 9 2
10 9 0 9 7 9 13 4 9 10 2
9 12 9 9 2 9 0 13 4 2
13 2 11 2 9 9 9 9 13 3 10 12 9 2
14 15 9 9 7 9 9 13 13 2 0 13 13 4 2
7 9 9 9 13 4 3 2
12 15 9 13 4 7 13 10 13 4 9 2 2
9 7 10 13 9 0 7 9 0 2
17 9 10 9 13 2 11 13 4 12 9 0 13 7 10 13 9 2
10 12 9 13 13 4 2 9 2 9 2
10 12 11 9 13 4 3 2 12 2 2
13 9 0 2 11 2 11 2 11 7 11 13 4 2
10 15 9 13 13 4 9 10 0 13 2
6 10 9 13 9 10 2
13 9 9 9 13 9 15 9 9 13 9 13 4 2
6 9 9 13 9 13 2
7 10 9 12 13 4 3 2
12 3 9 7 3 13 4 0 9 13 12 9 2
17 11 9 9 13 4 9 13 2 13 4 10 9 9 13 4 13 2
17 12 11 11 11 9 13 4 9 2 9 12 9 9 13 13 4 2
4 9 13 9 2
8 14 2 14 4 3 13 9 2
9 9 7 3 13 2 9 9 13 2
6 9 9 12 13 4 2
14 13 4 9 9 7 9 10 9 7 9 13 4 9 2
7 10 9 10 7 13 4 2
13 11 9 13 4 12 9 10 2 9 13 4 3 2
15 9 9 13 4 2 11 9 0 9 9 13 13 4 9 2
9 9 2 7 2 14 4 9 13 2
4 9 0 13 2
9 12 9 2 7 2 0 13 9 2
9 9 9 13 13 4 11 12 13 2
6 9 15 9 13 13 2
8 9 4 9 3 15 13 4 2
16 9 9 7 0 13 9 9 3 13 4 2 13 0 9 2 2
9 15 9 13 4 2 13 4 11 2
6 9 13 11 9 0 2
12 11 13 14 4 3 13 2 7 0 11 13 2
11 7 9 9 13 4 2 14 9 13 9 2
6 9 12 9 13 4 2
7 11 13 13 4 9 2 2
19 12 13 4 11 11 11 12 9 9 13 2 7 9 0 7 0 13 4 2
26 10 2 13 13 11 13 10 13 2 7 3 2 15 9 9 12 0 13 4 2 2 13 11 11 9 2
16 3 11 9 13 4 9 9 10 13 4 9 10 9 3 13 2
11 11 2 7 2 11 13 4 2 12 2 2
10 2 15 9 13 4 10 13 4 2 2
11 0 13 13 2 7 3 13 4 9 13 2
17 13 13 4 11 15 9 13 7 11 9 2 9 2 13 13 4 2
15 9 10 2 11 9 12 9 0 7 12 0 13 9 13 2
19 7 2 11 12 9 9 13 4 3 11 13 2 7 10 9 13 4 3 2
9 11 9 0 9 9 13 4 11 2
12 13 0 13 4 9 13 7 14 4 9 13 2
10 3 9 9 9 0 13 4 9 12 2
7 3 13 9 13 9 13 2
13 3 2 0 9 13 9 0 9 13 14 13 3 2
6 9 0 10 9 13 2
4 9 13 4 2
8 9 12 9 13 12 9 9 2
9 12 9 13 4 9 13 9 9 2
4 2 9 13 2
6 7 9 12 13 10 2
11 9 14 13 7 9 14 13 14 13 9 2
11 9 10 9 3 12 9 7 9 13 0 2
17 11 9 9 13 4 7 3 11 2 0 2 9 9 12 13 4 2
18 9 12 13 13 4 2 9 13 7 9 12 9 13 4 13 13 3 2
7 9 9 9 9 13 4 2
11 9 12 9 7 12 9 13 4 9 10 2
13 11 0 2 13 9 2 13 4 11 2 9 0 2
9 13 13 4 2 3 9 13 13 2
13 3 2 9 15 13 4 10 9 13 4 9 13 2
17 9 9 10 9 10 10 13 3 13 3 2 13 4 0 9 10 2
14 11 9 13 2 11 7 11 13 7 11 11 13 4 2
29 7 9 2 7 9 12 13 4 2 9 9 10 9 13 2 9 13 2 7 9 13 4 3 3 2 0 9 13 2
13 9 9 13 4 2 7 3 13 4 9 10 2 2
11 2 9 13 4 2 7 13 13 4 9 2
13 2 11 10 9 0 7 9 9 15 9 13 4 2
10 9 9 13 10 2 9 0 13 4 2
11 9 7 9 13 7 9 0 13 9 13 2
13 10 9 9 13 7 9 0 7 0 9 13 4 2
8 9 9 9 9 9 13 4 2
16 13 4 9 0 9 2 9 10 13 2 11 13 3 2 0 2
4 12 13 4 2
21 7 2 13 4 0 13 4 9 10 3 13 2 2 10 9 0 10 13 4 2 2
20 7 2 9 9 13 4 9 3 13 4 7 9 3 0 13 2 9 9 13 2
16 3 14 4 13 3 9 9 10 9 13 9 13 4 3 0 2
18 11 9 11 2 11 2 11 2 11 2 11 2 11 7 11 13 4 2
10 3 2 10 10 13 4 9 13 9 2
10 10 9 7 9 13 4 2 7 10 2
18 3 9 9 13 4 2 9 9 13 7 9 12 13 9 7 9 0 2
8 9 9 9 0 9 13 4 2
19 2 0 9 3 0 13 4 2 11 3 0 13 4 2 7 4 9 13 2
18 7 2 11 13 4 10 9 11 9 7 9 13 13 2 7 14 9 2
11 7 2 9 9 0 9 13 13 4 13 2
14 11 9 0 2 11 2 3 9 0 13 13 4 3 2
11 3 13 13 2 7 11 14 13 3 9 2
9 9 0 9 7 13 13 9 10 2
3 9 13 2
8 9 10 2 9 2 13 4 2
16 9 7 9 13 4 9 13 4 9 13 13 4 7 9 13 2
8 3 9 12 9 0 13 4 2
13 11 12 9 13 4 9 2 9 0 13 4 3 2
4 0 13 4 2
6 11 12 9 13 4 2
8 2 15 13 4 9 4 13 2
11 9 10 12 9 13 7 12 9 13 0 2
8 7 9 12 13 2 15 9 2
9 2 9 7 0 9 9 13 3 2
13 9 12 12 9 13 4 2 7 9 13 13 9 2
9 9 9 12 7 11 9 12 13 2
9 7 2 9 13 2 13 2 4 2
5 10 9 0 13 2
6 3 13 4 0 13 2
17 3 2 9 10 9 13 9 9 13 4 2 13 4 9 13 3 2
9 3 3 3 13 10 13 4 9 2
5 3 14 4 13 2
6 3 13 4 9 9 2
15 11 13 9 9 13 4 11 2 11 10 9 12 9 13 2
17 11 2 11 9 2 13 4 9 0 2 3 13 4 3 12 9 2
10 11 2 11 9 9 9 13 4 3 2
11 9 13 9 2 10 13 13 4 9 0 2
10 13 12 9 2 7 2 3 0 13 2
10 3 12 13 4 11 2 7 12 11 2
6 9 0 13 4 9 2
19 3 9 0 13 4 2 7 9 0 14 4 3 13 13 2 9 0 13 2
12 11 11 13 4 12 9 9 9 13 13 4 2
5 9 2 9 13 2
6 13 13 13 4 9 2
17 2 9 9 13 13 4 2 7 10 9 13 7 9 13 13 4 2
3 13 4 2
12 11 9 14 4 13 11 9 9 2 9 9 2
13 11 10 9 7 2 11 7 11 0 9 13 4 2
6 11 9 13 4 9 2
15 2 12 9 13 4 9 2 7 3 9 0 13 4 0 2
6 15 9 9 13 4 2
12 12 9 2 11 2 11 7 11 13 4 9 2
10 11 9 12 13 4 2 10 9 13 2
5 13 9 13 9 2
8 9 2 15 9 9 10 13 2
7 10 13 12 9 9 0 2
5 0 9 12 13 2
7 9 0 13 4 9 13 2
17 9 9 13 13 4 11 9 0 13 3 7 9 9 9 13 4 2
9 9 9 13 4 9 13 13 3 2
20 11 11 9 11 9 2 0 2 13 7 11 13 13 13 13 13 4 3 9 2
6 7 11 9 0 13 2
10 7 2 15 14 4 13 12 11 13 2
8 9 13 2 9 13 13 4 2
22 12 12 9 0 9 10 13 4 11 2 9 9 0 7 9 13 10 13 4 9 9 2
6 9 3 13 4 9 2
9 11 2 9 2 13 4 13 9 2
18 10 12 9 13 11 2 7 3 13 13 4 2 6 10 13 4 2 2
8 11 2 11 2 13 4 11 2
7 13 2 9 0 13 11 2
13 11 11 0 13 4 11 9 13 13 4 9 0 2
12 15 3 13 9 3 0 13 13 4 11 9 2
6 10 13 4 11 9 2
18 13 9 2 11 2 12 9 9 0 9 2 13 4 7 13 4 11 2
15 9 2 13 9 9 13 9 9 2 3 9 13 4 13 2
14 0 13 2 10 10 13 4 9 9 9 9 0 13 2
28 11 11 11 9 3 13 4 9 0 12 9 2 13 2 4 7 13 9 13 4 2 9 0 9 9 13 3 2
8 15 9 9 9 13 13 4 2
12 11 2 7 2 2 9 13 2 13 4 13 2
13 9 13 4 9 2 12 9 9 13 9 12 9 2
5 12 9 13 13 2
9 11 2 11 7 10 0 9 13 2
11 3 3 2 3 3 2 11 13 4 13 2
15 9 0 9 0 13 4 9 0 2 9 9 9 13 4 2
10 9 13 9 2 11 13 4 13 12 2
9 3 13 2 3 2 9 10 9 2
19 9 3 13 4 12 9 2 12 9 2 7 3 13 4 12 9 13 4 2
9 0 9 2 7 2 3 0 13 2
13 2 9 14 4 3 13 2 7 9 10 13 4 2
12 2 9 13 4 2 7 10 3 0 13 15 2
12 9 9 9 9 10 9 13 9 9 13 3 2
8 9 13 14 13 9 0 11 2
15 11 13 4 2 3 11 9 13 4 9 9 9 12 13 2
13 9 9 13 9 13 4 7 9 13 4 9 9 2
19 2 11 9 13 9 13 4 7 15 7 9 13 4 3 9 0 13 13 2
12 10 9 9 13 4 12 9 9 0 9 9 2
9 9 12 13 7 12 9 13 4 2
7 9 2 9 2 13 4 2
14 3 2 13 4 12 9 7 12 9 2 3 10 13 2
21 12 9 9 9 13 2 14 13 9 0 2 7 9 3 3 13 3 9 13 3 2
14 11 3 13 4 14 4 0 13 2 9 10 13 4 2
8 9 13 4 9 9 9 13 2
19 2 15 9 10 13 2 9 10 13 9 13 4 9 9 12 13 9 2 2
5 12 9 13 4 2
7 2 9 7 9 9 13 2
13 9 10 9 9 9 13 4 2 7 9 13 4 2
7 9 11 13 4 2 12 2
7 9 13 13 4 11 9 2
14 11 9 11 13 9 12 12 9 13 7 12 13 4 2
24 10 13 4 13 12 2 7 9 9 14 13 13 9 2 10 13 13 4 11 13 4 12 9 2
8 0 14 13 9 9 13 4 2
12 7 2 9 9 10 13 4 9 9 13 4 2
10 9 13 13 13 4 9 0 12 9 2
8 10 9 2 9 13 13 4 2
9 9 2 7 2 9 0 13 4 2
12 12 9 13 4 11 2 7 12 13 4 9 2
7 11 9 13 4 9 9 2
6 10 13 9 0 9 2
6 2 10 9 13 4 2
5 9 9 10 13 2
6 11 9 0 13 10 2
12 11 9 0 2 9 3 13 4 9 13 13 2
12 10 13 7 9 10 9 13 0 13 4 9 2
16 3 14 13 9 13 7 9 13 9 13 11 2 13 2 13 2
22 11 2 9 13 4 2 3 13 4 14 13 10 9 10 13 2 9 10 3 13 7 2
16 9 13 11 9 2 11 9 7 13 4 2 12 13 4 13 2
17 2 9 10 0 13 9 13 7 0 13 9 9 3 3 13 2 2
22 13 2 11 2 9 10 9 2 13 4 2 2 11 9 13 4 9 7 9 13 2 2
17 9 3 13 4 9 9 13 2 7 9 13 3 9 9 9 13 2
29 11 13 13 3 2 11 9 11 9 13 10 3 7 3 9 7 9 13 4 2 7 9 0 13 7 13 4 3 2
11 12 12 9 11 13 4 2 11 7 11 2
7 11 9 9 12 13 4 2
9 9 13 4 12 9 0 9 13 2
19 9 10 12 9 9 7 9 9 13 4 2 7 0 9 0 7 0 13 2
19 12 9 13 4 9 2 11 11 0 13 4 12 2 7 11 7 11 12 2
7 11 9 9 7 3 13 2
7 13 4 10 9 12 9 2
15 12 9 9 10 8 0 13 2 10 9 12 9 13 4 2
11 11 9 9 12 13 4 7 9 0 13 2
4 10 13 4 2
6 7 14 13 10 14 2
9 9 2 7 2 0 9 13 4 2
13 9 9 11 11 9 13 7 14 4 9 0 13 2
11 9 0 12 7 9 0 13 13 15 9 2
9 9 9 10 2 9 9 13 4 2
14 7 2 11 9 13 4 12 9 14 4 13 9 13 2
6 11 7 11 13 4 2
13 12 3 11 13 9 13 7 12 0 9 13 4 2
11 9 9 2 11 9 9 0 13 4 3 2
10 3 9 0 13 4 13 4 11 9 2
7 11 12 9 13 4 9 2
16 9 9 13 4 13 4 2 7 2 9 13 13 9 13 13 2
15 10 12 9 13 4 11 11 11 9 9 11 11 11 9 2
20 14 4 9 10 13 13 2 7 9 10 13 9 13 0 3 13 2 2 13 2
5 11 9 13 4 2
16 11 9 13 2 9 12 9 9 9 13 4 9 9 11 9 2
9 3 9 13 13 4 13 15 9 2
10 12 9 11 11 13 4 2 12 2 2
30 13 13 11 7 11 9 14 13 9 10 2 7 9 7 9 7 0 13 9 13 2 7 9 9 10 0 13 9 10 2
7 7 12 9 0 13 4 2
22 0 9 10 2 9 9 13 9 13 2 9 0 2 9 0 7 9 0 13 9 4 2
31 9 11 2 11 2 11 7 11 2 2 11 2 11 2 11 7 11 2 7 11 2 11 2 11 2 11 2 13 10 9 2
5 9 7 13 4 2
15 9 12 12 9 9 13 4 2 7 12 9 13 4 9 2
10 13 2 9 0 13 4 9 13 0 2
8 11 9 0 13 4 3 7 2
15 2 9 2 9 2 9 2 9 2 9 10 13 4 9 2
12 0 13 4 2 11 9 0 7 9 13 4 2
17 2 7 3 13 4 12 9 10 9 7 9 14 4 9 13 2 2
14 11 10 9 9 13 4 9 10 13 9 13 13 4 2
15 11 0 9 0 13 4 13 9 9 0 13 4 13 4 2
13 10 13 4 9 13 13 4 2 9 0 13 4 2
11 9 12 11 9 7 9 13 9 13 4 2
11 11 9 13 9 2 11 9 12 13 4 2
10 11 9 0 2 11 9 13 13 13 2
20 3 2 12 11 3 13 9 2 12 9 9 13 11 2 7 11 12 10 14 2
6 12 9 0 13 4 2
19 9 12 14 13 0 0 9 13 2 7 11 9 9 10 13 4 11 9 2
14 2 9 9 9 13 9 13 9 2 9 0 13 2 2
6 9 9 13 13 4 2
11 9 9 12 13 7 13 4 3 13 9 2
11 11 9 13 2 7 9 13 9 13 4 2
6 12 13 7 9 13 2
7 0 13 4 12 9 2 2
13 11 2 11 2 11 7 11 7 13 9 13 4 2
12 9 9 13 4 2 9 13 9 13 2 2 2
5 9 11 9 13 2
7 3 11 13 4 9 10 2
21 2 14 2 13 3 2 11 2 11 2 11 7 12 13 4 2 7 15 9 0 2
8 13 3 7 13 13 4 10 2
13 11 3 13 4 9 2 9 9 7 9 9 13 2
9 12 9 13 2 7 9 9 13 2
21 11 0 13 4 12 9 13 2 7 2 9 9 7 9 0 2 13 4 13 4 2
7 9 13 9 13 9 10 2
12 2 15 9 14 4 3 13 2 7 9 13 2
7 9 9 13 4 2 0 2
17 11 0 9 13 4 12 9 7 9 10 9 9 13 4 12 9 2
5 10 9 10 13 2
8 10 7 11 9 10 13 4 2
9 9 10 15 9 13 15 9 13 2
18 9 9 9 0 13 4 2 12 9 9 13 9 13 4 11 11 9 2
6 13 4 9 2 13 2
12 9 9 12 13 4 2 15 9 9 13 9 2
5 15 13 4 9 2
10 7 12 13 4 2 9 9 12 9 2
13 2 0 10 9 13 9 13 15 9 9 9 2 2
8 13 7 9 13 13 4 3 2
8 10 9 13 4 13 4 11 2
9 9 2 0 2 13 13 3 11 2
8 9 0 9 0 13 13 4 2
12 9 13 4 9 2 9 9 2 13 4 9 2
43 2 9 9 2 9 9 2 9 0 2 9 2 9 7 9 0 9 2 9 7 9 0 2 9 0 2 9 9 9 2 9 0 9 7 9 0 0 2 13 13 4 11 2
14 9 7 9 13 9 0 7 9 3 13 9 0 13 2
9 12 9 13 4 2 12 9 9 2
25 10 9 9 0 10 13 2 11 9 9 13 9 13 2 0 10 13 7 9 0 9 9 0 13 2
5 0 9 0 13 2
12 9 0 0 10 7 13 4 9 0 13 2 2
9 11 9 13 7 12 9 0 13 2
10 11 7 11 9 0 13 4 12 9 2
6 2 13 4 11 2 2
6 7 3 10 13 13 2
5 3 13 4 9 2
16 0 9 13 9 13 4 9 9 0 13 2 11 13 7 14 2
7 0 9 9 12 13 4 2
10 11 7 11 9 9 9 13 4 9 2
8 12 13 4 11 12 9 0 2
15 9 9 10 3 13 4 11 11 11 9 2 11 13 4 2
10 3 3 11 9 9 13 4 9 12 2
11 3 8 11 9 0 13 4 9 13 9 2
26 11 11 11 9 9 11 11 8 11 12 13 4 3 2 9 10 13 9 10 9 0 13 11 11 9 2
16 0 9 14 4 9 0 7 0 9 13 2 9 0 9 7 2
21 11 2 3 2 13 13 9 9 7 11 12 9 9 13 9 13 7 10 13 4 2
9 14 4 10 13 9 13 4 9 2
11 9 0 9 13 11 9 0 7 9 9 2
8 9 10 12 13 13 11 9 2
12 11 13 4 12 12 9 2 11 9 12 9 2
12 11 9 10 13 4 9 13 2 11 13 4 2
27 11 11 2 11 11 7 11 11 2 7 2 3 13 4 2 10 0 8 3 2 7 10 9 9 13 3 2
12 9 0 13 4 2 7 9 7 9 13 4 2
8 7 3 13 4 10 9 12 2
3 3 13 2
15 9 9 13 4 2 12 12 9 13 12 12 13 13 4 2
18 11 9 9 3 13 4 2 0 12 12 9 12 13 4 9 13 9 2
9 12 9 7 2 9 13 13 4 2
17 2 0 13 9 0 0 12 13 2 9 7 9 0 0 13 4 2
14 11 9 0 13 7 10 13 4 11 9 9 9 10 2
13 11 13 2 11 9 9 0 13 4 12 12 9 2
5 10 9 13 4 2
18 9 9 13 4 11 2 7 11 9 9 3 13 13 13 4 12 9 2
6 9 10 0 0 13 2
7 9 0 13 4 2 7 2
4 13 4 9 2
11 11 2 7 2 14 4 9 10 3 13 2
4 13 4 11 2
17 9 11 11 11 13 4 3 9 11 11 9 2 11 9 0 9 2
14 11 13 4 9 9 0 7 9 13 4 9 13 9 2
8 2 13 4 11 9 13 9 2
8 12 9 9 9 9 13 4 2
28 11 9 9 12 9 13 13 3 2 0 9 9 13 4 7 9 0 13 4 9 9 12 9 9 13 4 9 2
3 3 13 2
8 12 9 9 0 13 4 3 2
5 9 0 13 4 2
19 7 0 9 0 9 3 13 9 9 13 4 0 9 10 7 9 0 12 2
9 11 13 2 0 9 10 13 4 2
6 9 12 9 13 4 2
20 11 11 11 0 12 9 7 13 11 0 12 9 2 0 0 13 0 9 13 2
8 0 2 0 7 0 13 4 2
14 12 9 13 13 9 7 12 9 13 9 9 13 4 2
7 9 9 11 9 13 4 2
14 9 9 10 11 13 4 12 9 13 4 9 0 9 2
26 11 9 13 9 9 0 9 0 13 4 2 7 9 0 9 0 7 9 13 7 9 9 13 13 13 2
6 9 0 12 13 4 2
12 2 9 13 9 0 13 2 10 9 13 4 2
15 9 9 0 9 13 4 3 2 7 11 14 4 9 13 2
6 9 7 2 0 13 2
10 0 9 3 13 13 4 9 13 4 2
10 14 4 13 10 13 4 9 12 13 2
37 11 9 12 9 0 0 2 0 7 0 13 13 4 2 7 10 7 10 2 11 2 2 9 2 9 2 9 9 7 9 9 10 2 13 13 4 2
18 3 2 3 9 0 13 4 10 9 2 9 7 9 12 9 2 3 2
9 9 9 13 10 9 14 13 11 2
11 12 9 13 7 2 9 13 14 4 9 2
16 9 13 9 9 13 4 9 2 7 11 9 13 4 0 9 2
5 13 13 2 3 2
7 9 10 9 12 13 4 2
11 9 13 9 0 10 3 13 13 4 13 2
9 2 6 14 4 9 10 9 13 2
6 2 13 4 9 2 2
5 3 13 4 0 2
15 2 13 9 10 9 0 12 13 2 15 2 3 13 9 2
14 0 9 9 2 9 7 9 9 9 0 13 4 9 2
4 9 3 13 2
10 9 10 9 13 9 13 9 0 9 2
6 11 9 10 13 4 2
14 14 4 13 9 3 10 13 14 4 2 9 13 3 2
12 9 13 4 11 9 2 7 13 4 9 9 2
11 9 0 9 13 4 9 0 9 9 13 2
7 12 9 12 13 4 9 2
19 3 9 0 13 7 2 9 9 10 13 4 9 12 12 9 7 9 13 2
11 11 14 4 13 2 15 15 9 13 7 2
22 2 3 3 7 9 0 13 4 13 4 15 9 9 0 13 11 10 13 9 0 2 2
4 11 13 0 2
4 3 13 4 2
19 3 2 9 9 13 4 7 9 9 9 13 13 4 9 9 9 13 4 2
5 12 9 13 4 2
9 2 10 9 14 4 9 9 13 2
7 12 9 9 13 9 3 2
9 11 13 4 9 9 13 4 12 2
16 15 9 13 11 9 13 4 10 9 9 9 0 0 12 13 2
10 9 9 9 0 13 4 10 13 13 2
12 9 13 13 4 13 2 7 3 13 4 13 2
16 9 0 9 9 3 0 13 2 9 3 9 13 9 13 4 2
20 11 2 11 2 13 4 3 11 9 9 2 7 11 11 0 13 4 9 9 2
16 15 13 13 3 2 9 0 13 4 2 7 9 12 13 13 2
8 7 11 9 9 13 4 9 2
22 11 9 9 2 11 13 13 9 13 2 9 9 13 4 3 2 9 7 9 9 13 2
14 9 2 9 2 9 12 2 7 9 0 13 9 10 2
5 2 14 4 13 2
8 3 2 10 9 9 13 4 2
17 2 14 13 10 9 13 15 13 2 10 9 2 11 0 9 13 2
8 9 13 4 9 2 14 0 2
16 2 9 13 9 12 7 0 13 2 7 9 13 13 4 2 2
5 13 4 9 2 2
5 12 9 13 11 2
7 9 9 13 9 13 4 2
18 7 11 13 4 9 2 7 15 13 4 2 13 4 9 10 9 13 2
13 11 7 13 4 11 13 9 0 10 14 4 0 2
26 2 15 13 4 12 9 13 4 10 2 7 3 13 4 12 13 2 2 13 3 2 3 2 9 11 2
8 11 9 9 13 4 11 11 2
8 10 13 2 9 10 13 4 2
12 9 9 13 4 9 2 9 9 13 13 4 2
21 12 9 2 11 2 12 13 13 4 9 9 9 2 7 9 13 11 13 3 13 2
7 2 3 13 4 9 10 2
11 9 0 9 13 7 2 9 2 13 4 2
9 3 13 9 13 9 13 9 13 2
11 9 9 13 4 9 0 9 7 9 13 2
15 7 2 9 7 9 3 13 4 9 14 4 0 9 13 2
22 9 3 13 4 9 7 2 7 11 9 9 13 4 11 11 7 11 14 4 11 13 2
4 12 13 4 2
8 9 12 13 4 11 9 0 2
6 12 9 13 4 9 2
4 9 3 13 2
14 7 3 7 9 0 13 4 2 7 9 0 13 13 2
10 9 13 3 2 9 0 13 9 13 2
10 7 9 13 10 13 9 13 3 2 2
8 9 0 12 12 9 13 4 2
5 13 4 9 10 2
8 3 3 2 9 13 4 10 2
24 9 9 9 9 9 9 9 9 13 9 13 4 2 7 9 2 9 13 4 9 2 13 4 2
8 9 2 11 9 9 13 4 2
8 11 9 3 9 9 13 4 2
11 3 3 13 7 2 7 9 0 12 13 2
14 9 9 0 13 2 7 3 9 10 13 13 4 13 2
17 11 9 0 9 9 7 9 10 9 13 9 9 13 13 4 11 2
18 9 2 13 4 9 0 3 13 7 8 9 9 9 15 0 13 4 2
15 11 7 11 15 13 13 11 9 9 13 14 13 9 12 2
7 2 9 9 0 13 9 2
9 9 0 2 0 7 9 13 13 2
9 9 3 13 4 12 11 11 9 2
5 15 9 9 13 2
9 3 10 13 11 9 7 9 9 2
6 2 15 0 9 13 2
7 9 10 0 9 13 13 2
9 3 13 4 13 2 3 13 7 2
13 11 2 11 7 11 2 7 2 14 13 13 9 2
8 11 2 7 2 12 13 4 2
8 11 10 9 13 4 9 10 2
5 9 3 13 4 2
8 2 9 9 13 9 13 2 2
10 9 0 10 13 4 7 9 13 4 2
10 7 2 11 11 9 9 13 4 9 2
9 9 12 13 4 9 10 0 13 2
21 9 0 9 2 9 12 9 13 14 4 13 2 13 2 9 0 13 4 10 9 2
9 9 10 13 9 10 13 9 13 2
19 3 2 7 2 11 9 11 11 0 9 13 4 12 9 13 4 2 9 2
13 11 7 3 13 2 7 10 9 13 4 11 3 2
6 7 13 13 4 9 2
12 7 2 11 9 13 4 0 9 0 13 4 2
14 2 9 9 13 7 3 10 9 12 9 9 7 9 2
6 9 2 12 9 13 2
12 9 0 9 3 13 13 4 11 11 11 11 2
6 13 13 9 9 13 2
6 3 13 9 13 9 2
18 9 2 9 2 9 9 2 9 2 9 2 9 2 13 4 9 9 2
4 0 13 9 2
5 7 14 13 10 2
6 9 12 14 13 0 2
6 12 12 13 4 9 2
6 12 9 3 0 13 2
5 11 9 13 4 2
12 9 2 7 2 14 13 2 7 9 9 13 2
7 9 9 9 0 13 4 2
11 14 4 11 3 13 4 8 10 13 3 2
6 10 13 9 0 9 2
11 3 2 7 2 11 14 4 9 9 13 2
13 11 9 13 4 3 2 0 13 7 9 0 13 2
13 14 4 9 13 2 14 4 3 9 0 10 13 2
13 9 12 9 9 14 13 13 9 9 9 13 13 2
14 2 9 10 2 7 2 0 14 13 15 2 9 7 2
20 9 2 12 12 9 7 9 13 4 7 12 9 13 4 2 12 9 9 2 2
12 2 9 13 4 11 13 2 11 9 13 2 2
5 9 9 13 11 2
13 2 3 14 13 9 9 13 9 2 9 13 4 2
11 9 0 13 9 2 0 9 13 13 3 2
9 0 9 9 0 13 13 4 2 2
19 2 9 9 0 13 4 2 7 14 4 9 13 7 0 9 0 13 10 2
6 2 9 12 13 9 2
7 11 12 9 13 0 4 2
19 9 11 11 0 13 4 2 14 13 9 2 12 9 0 13 9 0 7 2
7 2 9 10 13 4 2 2
7 3 2 3 13 13 4 2
6 15 10 9 13 4 2
12 9 2 11 7 11 13 4 9 2 12 9 2
8 3 9 13 4 11 9 13 2
8 14 13 0 9 9 13 9 2
17 2 11 0 9 9 13 4 7 9 0 13 4 13 4 9 9 2
7 2 13 2 9 2 13 2
14 15 13 4 9 10 9 13 7 13 4 2 7 14 2
22 11 2 7 2 14 4 13 9 13 9 13 2 10 9 9 9 14 13 9 9 2 2
8 9 9 9 13 4 13 4 2
18 2 9 3 3 13 4 2 7 10 13 4 9 2 2 13 4 11 2
9 3 2 7 2 9 9 13 13 2
13 10 13 11 12 9 9 9 13 4 3 7 3 2
13 9 9 10 9 7 9 10 9 7 9 13 13 2
30 11 3 13 12 9 13 9 2 11 9 13 9 4 3 12 9 2 12 2 2 7 10 13 4 2 11 2 11 2 2
7 9 9 9 9 0 13 2
19 7 2 9 9 10 11 9 13 9 2 11 9 9 12 13 4 13 11 2
12 11 11 0 10 12 9 9 13 4 3 11 2
15 9 12 9 2 9 7 9 10 2 13 4 13 4 11 2
12 3 13 4 9 10 13 9 12 13 13 4 2
5 9 0 10 13 2
5 9 0 0 13 2
16 3 7 9 13 9 13 9 13 4 2 7 3 14 4 13 2
30 9 2 11 9 13 4 9 13 2 7 2 9 2 7 2 11 9 13 4 0 2 7 2 3 2 9 13 4 9 2
6 11 9 7 13 9 2
5 15 9 9 13 2
13 9 13 12 9 13 4 7 3 9 0 13 4 2
6 9 3 0 13 4 2
18 9 9 9 9 13 3 2 3 10 9 0 7 0 9 13 9 13 2
14 2 9 9 13 7 3 10 9 12 9 9 7 9 2
13 13 9 9 12 9 13 11 13 4 9 13 4 2
10 9 9 2 7 2 14 4 10 13 2
13 11 9 13 4 9 13 2 12 9 9 13 13 2
12 12 9 2 3 13 9 10 12 9 13 4 2
7 9 7 13 4 9 9 2
13 9 13 7 2 10 9 13 4 11 9 10 9 2
3 13 4 2
6 14 13 10 9 13 2
10 13 4 13 14 4 9 10 10 13 2
21 14 11 14 11 9 0 13 4 2 7 11 11 11 9 9 0 13 4 13 4 2
12 0 13 2 7 9 13 4 3 13 4 9 2
4 9 9 13 2
7 3 9 9 9 13 4 2
14 9 10 9 0 0 2 0 11 0 2 13 4 11 2
8 11 9 12 9 9 13 11 2
5 7 15 10 13 2
10 11 7 11 9 3 13 4 3 7 2
7 9 10 9 12 13 4 2
11 9 10 9 13 4 9 10 9 9 13 2
6 12 9 13 4 9 2
4 14 13 3 2
7 9 13 9 12 2 6 2
8 10 12 9 13 4 9 13 2
14 9 10 2 9 13 2 9 0 0 7 0 13 4 2
14 2 15 11 12 13 7 11 11 13 2 13 13 2 2
9 0 13 2 7 13 13 15 9 2
15 2 9 0 13 4 3 2 7 13 13 4 9 0 9 2
22 13 12 9 13 4 12 9 11 11 11 11 9 2 7 3 13 4 12 9 10 9 2
22 11 9 9 12 2 9 12 7 9 12 9 2 2 10 9 0 2 2 9 13 4 2
21 9 9 9 9 9 13 9 13 4 2 7 9 10 13 13 4 14 9 14 9 2
5 3 13 9 13 2
6 2 9 13 4 2 2
9 11 10 14 4 13 11 9 9 2
15 11 9 2 9 9 0 0 14 13 9 9 13 4 9 2
11 2 3 13 9 0 15 9 13 7 13 2
7 9 0 10 13 4 15 2
11 11 11 9 9 0 13 9 13 4 3 2
12 9 9 2 11 13 4 12 12 2 12 2 2
7 9 7 0 13 9 13 2
13 11 9 13 4 11 9 2 12 9 10 13 3 2
7 9 9 13 4 9 9 2
9 12 9 10 3 13 4 14 13 2
10 3 2 9 9 13 9 13 4 11 2
6 2 11 9 13 2 2
15 2 7 9 10 9 2 9 13 4 2 9 13 9 13 2
21 9 12 9 9 13 4 9 9 9 2 7 13 9 10 3 13 4 9 15 13 2
6 2 13 2 9 9 2
7 14 13 7 3 9 10 2
17 9 10 13 4 0 7 9 9 9 13 0 10 9 13 9 13 2
7 15 11 11 13 4 9 2
14 9 10 13 3 2 12 9 9 12 13 4 13 4 2
12 13 13 4 2 7 2 12 9 9 9 13 2
10 9 0 10 12 12 9 13 4 0 2
13 3 13 4 9 2 9 2 9 0 10 9 13 2
28 9 13 2 11 9 12 12 9 9 12 13 9 2 9 12 9 9 13 4 12 9 9 0 2 11 13 4 2
5 3 13 13 4 2
7 9 0 13 13 4 3 2
8 14 13 3 7 9 13 9 2
20 11 11 9 12 9 13 4 9 9 9 12 9 2 12 2 12 7 12 2 2
10 9 9 2 11 9 9 0 13 4 2
8 11 13 4 2 3 13 4 2
5 11 0 9 13 2
13 14 13 14 13 10 13 2 9 13 13 4 7 2
14 2 9 13 9 13 2 3 13 4 13 4 7 14 2
6 7 2 0 13 9 2
13 9 0 13 4 2 7 9 0 14 4 10 13 2
14 9 9 9 14 13 7 2 9 0 13 4 10 9 2
5 10 9 13 4 2
15 0 9 7 9 0 13 4 9 7 11 13 4 9 0 2
7 9 9 13 13 9 13 2
5 2 2 0 13 2
5 9 0 9 13 2
5 3 13 11 12 2
7 9 9 9 13 9 11 2
3 13 4 2
8 3 13 4 9 12 9 12 2
9 3 11 11 0 13 4 9 9 2
15 9 13 9 13 9 2 13 7 13 13 9 13 4 9 2
28 11 2 11 2 9 2 9 13 13 4 2 7 9 12 12 9 10 13 3 11 2 13 7 13 2 13 4 2
23 11 9 11 11 9 0 13 4 3 0 9 2 11 11 9 13 7 13 9 11 9 9 2
9 11 11 11 9 3 13 9 13 2
8 3 2 9 10 9 13 4 2
15 11 0 12 13 4 9 2 7 3 14 13 9 9 9 2
13 9 7 9 9 13 2 2 10 9 10 14 13 2
16 15 9 2 15 9 2 15 9 2 9 10 9 10 13 4 2
8 11 11 7 13 9 13 4 2
7 2 10 13 4 2 11 2
16 7 13 14 4 9 9 13 2 7 2 9 9 0 13 9 2
17 10 13 7 2 7 2 3 13 4 9 9 9 3 13 4 9 2
12 12 9 14 4 9 13 11 2 11 7 11 2
12 9 9 9 13 4 2 7 14 4 9 13 2
13 9 9 11 13 4 2 7 9 13 4 3 9 2
10 9 2 3 9 0 13 7 13 4 2
5 2 3 9 13 2
6 9 9 12 13 4 2
17 9 2 3 2 12 9 13 4 2 9 12 13 7 12 13 4 2
16 11 7 11 3 13 2 7 11 12 13 9 13 4 13 4 2
7 15 9 0 13 4 10 2
15 11 13 4 3 9 0 12 13 2 9 0 12 13 3 2
21 2 9 0 13 2 15 9 12 13 4 9 10 9 7 9 10 9 9 13 2 2
8 2 3 9 0 13 4 2 2
14 11 11 9 12 11 13 4 9 13 11 13 14 4 2
9 3 13 13 4 10 13 9 9 2
18 9 0 9 10 13 13 4 2 11 9 13 4 13 2 9 2 13 2
9 13 4 13 9 9 13 4 13 2
6 11 9 10 13 4 2
15 15 0 13 12 7 12 9 13 7 10 7 10 13 9 2
15 15 9 13 4 3 13 4 2 7 3 13 4 9 9 2
15 12 3 13 4 3 13 4 2 7 12 13 4 9 13 2
23 9 7 9 2 11 2 11 2 7 11 2 11 2 2 13 4 11 11 9 9 12 9 2
7 13 13 9 13 9 9 2
10 2 3 2 7 13 4 9 9 2 2
5 15 13 4 9 2
22 2 0 9 14 13 13 4 7 3 2 0 2 9 7 9 13 4 9 13 4 2 2
9 10 13 3 13 13 4 2 7 2
12 3 2 9 13 4 2 9 15 13 14 4 2
10 11 11 12 9 7 13 4 11 9 2
11 9 9 13 4 2 10 13 9 0 4 2
8 2 12 9 9 13 4 2 2
4 2 14 13 2
10 12 9 9 13 4 12 9 13 4 2
22 11 9 11 9 13 4 0 9 2 12 9 2 9 0 2 9 13 7 13 9 13 2
8 11 13 11 9 12 13 4 2
11 9 9 13 4 2 9 9 13 13 3 2
13 9 12 9 13 4 2 7 13 13 9 13 4 2
8 15 3 10 9 13 4 3 2
11 9 0 9 13 4 2 9 0 13 3 2
7 3 13 4 9 9 9 2
6 2 13 9 9 9 2
7 9 9 0 9 13 4 2
6 2 13 4 9 2 2
5 9 2 0 13 2
24 13 4 14 4 10 13 2 9 12 9 12 13 13 4 2 7 9 9 3 13 4 10 2 2
19 7 2 11 9 9 13 13 9 2 7 2 3 2 11 9 9 9 13 2
8 12 9 13 4 11 9 12 2
7 7 11 3 13 4 9 2
17 9 9 13 4 12 9 7 2 7 14 4 13 9 13 9 10 2
10 7 11 13 4 10 3 14 4 13 2
5 7 2 10 13 2
9 3 2 12 9 9 13 4 11 2
17 13 4 11 7 9 0 9 0 13 4 9 9 9 13 4 3 2
16 12 9 9 0 13 9 2 12 13 4 11 9 9 9 9 2
9 12 9 7 2 9 13 13 4 2
13 14 13 10 9 13 2 10 9 13 4 9 13 2
7 9 9 7 13 13 4 2
8 9 9 2 9 9 13 4 2
7 11 9 15 13 4 3 2
6 3 13 15 9 0 2
14 9 12 13 4 9 2 11 11 11 9 9 9 13 2
11 11 0 13 2 11 13 4 7 0 13 2
12 11 9 0 9 13 2 11 9 7 0 13 2
5 9 12 9 13 2
5 9 0 13 10 2
5 12 9 13 4 2
9 2 0 13 9 3 0 13 2 2
16 14 4 9 0 13 2 7 3 2 3 13 4 12 9 13 2
8 9 10 13 9 13 13 4 2
20 11 11 9 9 12 9 3 9 7 9 9 13 4 13 4 3 11 11 9 2
8 9 9 0 13 4 12 9 2
7 10 13 4 9 10 13 2
11 10 0 9 10 9 0 12 13 9 13 2
20 11 3 13 4 9 2 13 2 10 13 4 2 3 9 13 7 9 13 4 2
24 9 2 7 2 14 4 0 13 2 7 14 4 0 9 13 13 2 9 14 13 3 13 2 2
13 11 13 3 13 0 13 4 9 12 13 9 13 2
7 13 4 9 13 13 4 2
7 2 10 13 13 13 10 2
9 9 13 7 9 11 13 4 3 2
6 8 2 10 13 9 2
10 2 9 14 4 9 9 13 9 13 2
5 11 12 9 13 2
8 3 9 0 7 0 13 4 2
9 0 12 9 3 13 13 9 9 2
7 9 2 10 13 0 13 2
8 11 9 9 9 13 9 13 2
6 13 7 9 13 9 2
11 3 2 9 9 9 13 9 9 7 9 2
9 9 9 11 11 0 9 13 4 2
9 10 9 13 2 7 3 3 13 2
4 9 13 13 2
16 2 12 9 13 7 2 9 13 14 4 9 13 4 11 13 2
10 9 0 13 15 9 0 13 9 13 2
20 11 0 9 2 9 9 13 2 12 9 9 13 7 9 0 9 0 13 4 2
9 11 9 3 13 4 9 0 9 2
6 2 9 10 13 4 2
16 11 11 7 11 11 0 9 9 13 9 13 4 9 10 9 2
9 7 13 4 13 2 9 13 4 2
8 0 7 0 13 4 3 9 2
21 11 11 9 13 4 9 9 2 12 9 2 9 0 2 9 13 7 13 9 13 2
12 10 12 9 9 13 4 7 12 9 7 12 2
24 10 13 4 2 13 4 14 13 2 15 13 4 9 2 2 7 9 8 2 0 13 2 13 2
7 3 7 3 10 13 4 2
9 11 9 12 12 3 13 4 9 2
7 11 10 10 0 3 13 2
20 11 11 11 9 0 9 10 9 7 11 13 9 13 9 10 9 13 4 3 2
7 7 2 9 10 13 4 2
5 7 9 0 13 2
12 9 9 9 2 11 2 9 9 13 4 9 2
27 9 9 9 2 9 9 2 11 9 13 13 4 11 9 9 9 9 13 4 10 7 10 9 13 13 9 2
5 13 13 15 13 2
21 9 13 2 9 9 2 9 2 9 9 2 9 9 7 9 9 13 0 13 4 2
10 3 13 10 13 4 11 9 13 2 2
4 9 0 13 2
7 12 11 9 13 4 9 2
8 10 10 13 4 0 9 10 2
4 13 13 4 2
21 0 2 9 13 13 4 2 14 4 12 9 9 13 9 13 7 10 13 4 9 2
25 11 11 14 4 13 11 7 11 9 9 2 7 3 9 3 0 13 2 7 10 9 0 13 4 2
8 11 9 0 12 9 13 4 2
15 11 2 7 2 0 13 4 7 11 3 3 13 4 7 2
12 3 9 2 9 2 7 3 9 13 13 4 2
10 2 9 13 3 7 13 13 4 3 2
17 13 14 4 9 13 4 9 9 9 9 4 2 7 9 9 14 2
24 9 9 10 9 12 13 7 9 0 0 13 4 2 13 2 7 12 5 9 9 13 4 9 2
20 9 9 0 13 13 9 13 11 11 0 3 2 11 9 2 9 0 13 9 2
6 11 9 9 13 4 2
16 9 10 11 0 9 13 13 4 13 4 9 0 12 9 13 2
25 11 13 3 9 12 2 7 3 13 12 9 7 9 13 2 7 11 13 4 9 2 12 9 9 2
20 3 9 0 9 13 13 9 13 2 7 9 2 9 0 13 2 13 4 11 2
18 12 2 11 9 9 9 12 9 11 11 0 13 4 2 11 12 9 2
6 3 9 9 13 4 2
7 9 3 13 9 4 9 2
14 13 7 3 9 13 4 2 9 9 13 7 13 4 2
12 11 13 2 9 0 2 9 13 4 13 4 2
9 9 2 7 2 9 13 13 4 2
5 11 13 4 9 2
14 9 2 9 7 10 10 9 9 13 4 9 9 10 2
16 9 7 9 9 2 3 9 9 13 3 2 13 13 4 3 2
6 9 9 13 4 9 2
6 0 13 4 9 13 2
19 11 9 13 3 2 9 12 9 13 9 12 13 4 7 9 12 13 4 2
6 9 10 9 9 13 2
8 11 9 0 13 4 13 11 2
11 12 9 9 0 13 9 13 12 9 12 2
12 9 12 9 13 4 9 12 0 9 13 4 2
13 11 9 13 9 4 9 10 13 13 4 10 9 2
5 15 7 9 13 2
21 9 13 4 9 0 0 9 13 4 3 11 2 3 10 12 9 13 4 13 4 2
12 7 12 12 13 4 3 14 4 10 9 13 2
8 2 15 10 13 9 13 2 2
23 11 2 12 9 12 9 9 13 4 7 9 12 13 10 9 9 9 2 9 7 9 13 2
5 7 10 9 13 2
26 9 9 13 10 9 12 13 2 7 13 9 0 13 9 9 10 13 9 2 7 10 13 9 13 4 2
15 3 13 4 11 11 9 9 0 13 7 9 3 13 9 2
6 7 9 13 9 13 2
13 9 0 13 7 2 14 4 9 9 13 9 13 2
6 2 10 13 2 11 2
6 12 9 13 4 11 2
7 11 9 13 3 13 4 2
4 9 3 13 2
12 10 13 7 2 11 13 13 13 4 11 9 2
10 9 12 9 9 9 13 13 4 11 2
24 9 9 0 13 4 12 9 7 3 13 4 9 13 2 9 13 7 9 9 9 9 13 2 2
6 9 10 9 13 4 2
28 11 10 14 4 10 9 0 13 2 9 13 13 2 9 9 0 12 9 13 13 4 2 15 9 9 13 13 2
8 9 13 4 7 13 9 9 2
7 3 13 9 13 3 13 2
23 9 9 13 9 13 4 3 9 13 9 2 7 3 3 13 4 14 13 15 2 0 13 2
9 10 9 2 0 7 9 13 4 2
10 12 9 13 4 11 9 10 9 12 2
21 9 0 0 9 0 9 11 9 13 9 13 13 4 2 7 14 4 9 0 13 2
10 11 13 9 14 4 10 9 9 13 2
7 3 9 0 13 9 9 2
7 11 9 2 7 2 13 2
10 2 11 9 0 7 13 13 4 2 2
13 9 9 10 13 4 9 2 15 9 13 4 3 2
8 2 3 9 13 15 9 2 2
16 11 13 13 4 9 12 9 2 7 12 9 12 13 12 9 2
6 2 10 13 4 9 2
31 9 12 5 9 13 4 2 9 0 13 7 3 13 7 13 13 4 7 3 9 15 13 13 4 2 9 0 7 13 4 2
11 11 9 0 13 7 11 13 3 0 13 2
5 11 9 7 13 2
13 7 9 13 4 10 9 2 3 0 13 9 13 2
14 9 9 9 9 13 9 0 13 9 9 9 9 12 2
15 3 2 11 9 13 4 2 7 9 13 4 15 9 13 2
8 12 9 13 9 13 0 10 2
17 2 6 2 6 2 7 11 9 13 2 9 9 13 4 2 10 2
15 3 9 13 4 11 9 2 7 3 9 2 11 13 4 2
9 0 14 13 13 4 11 9 0 2
10 9 13 4 10 9 11 9 3 13 2
5 3 13 4 9 2
10 11 13 4 11 12 9 9 2 3 2
17 10 9 2 9 2 12 9 7 12 9 7 13 4 13 4 11 2
17 9 13 13 2 13 9 0 9 9 0 12 8 0 13 13 13 2
5 9 3 0 13 2
19 11 11 9 0 0 9 10 9 9 12 13 4 13 4 3 9 9 9 2
15 11 9 14 13 13 2 9 14 4 9 13 12 12 9 2
13 3 13 4 3 2 3 13 4 12 9 13 9 2
20 10 13 2 9 9 13 4 3 2 7 11 13 13 4 2 0 9 13 4 2
11 9 0 2 9 9 9 9 9 13 4 2
4 13 13 4 2
9 12 9 13 13 4 11 13 9 2
9 13 13 4 7 14 4 13 13 2
14 11 11 11 9 11 9 13 4 3 9 9 0 13 2
15 7 2 3 2 9 7 9 13 4 2 9 12 2 11 2
14 3 2 11 9 10 13 4 9 11 11 13 13 9 2
8 0 13 4 12 9 13 9 2
12 7 2 9 0 9 3 9 13 4 11 9 2
16 3 9 3 13 4 13 13 4 2 7 9 10 13 9 0 2
4 9 10 13 2
8 9 3 14 13 13 4 3 2
11 9 12 13 13 13 4 2 9 13 4 2
6 12 9 13 4 9 2
16 11 12 9 13 9 0 13 13 4 3 13 4 15 9 11 2
8 3 13 14 4 9 0 13 2
8 2 3 13 4 2 3 2 2
10 2 9 9 9 7 10 9 13 4 2
8 11 9 13 7 9 13 4 2
12 9 9 9 13 4 9 9 10 13 4 9 2
6 11 9 3 13 4 2
9 3 7 12 9 9 12 13 4 2
21 11 9 13 9 13 4 2 7 11 9 0 13 9 0 12 13 7 3 13 4 2
11 9 9 7 9 9 9 13 7 13 4 2
6 11 9 13 4 3 2
4 9 9 13 2
10 13 4 2 11 9 9 2 2 9 2
9 9 10 2 9 9 3 0 13 2
8 11 7 11 7 9 13 4 2
10 10 9 2 11 7 11 13 4 9 2
10 7 2 3 2 15 9 13 13 4 2
12 2 14 13 10 9 2 9 9 13 9 13 2
9 11 7 0 13 4 9 10 9 2
6 14 13 10 13 4 2
8 2 10 13 2 13 13 4 2
6 10 13 0 9 9 2
4 10 9 13 2
13 14 12 2 14 10 2 0 9 13 9 13 4 2
11 9 9 7 9 9 9 0 13 4 10 2
9 11 7 11 9 11 9 13 4 2
8 9 9 11 13 4 12 9 2
9 2 15 10 7 13 4 9 10 2
9 9 0 7 9 0 9 13 4 2
15 3 11 13 9 0 9 2 7 3 14 13 9 9 0 2
6 3 14 13 0 0 2
8 11 0 13 3 9 3 13 2
7 11 13 4 11 12 9 2
8 2 0 2 3 9 13 13 2
7 10 10 13 4 11 3 2
29 7 9 9 13 13 9 2 7 9 2 7 0 9 3 13 13 4 2 9 13 4 2 7 3 9 0 13 4 2
6 9 12 13 4 0 2
14 9 13 4 9 9 13 2 11 9 0 9 13 4 2
16 2 7 3 11 11 13 2 3 2 13 4 9 10 9 13 2
6 9 0 9 9 13 2
5 12 12 9 13 2
9 2 0 9 13 13 7 13 4 2
11 9 3 13 13 4 2 9 0 13 4 2
7 3 2 0 0 13 9 2
8 2 7 2 14 4 15 13 2
4 15 13 3 2
7 11 9 0 9 13 4 2
25 2 9 0 3 13 13 4 2 10 13 9 0 13 4 9 2 7 10 13 9 13 9 0 2 2
6 11 9 13 4 11 2
7 9 9 0 13 9 13 2
13 11 9 13 9 2 11 2 11 7 11 13 4 2
7 2 14 2 14 13 10 2
5 2 0 13 4 2
11 9 9 7 14 4 0 9 13 12 9 2
8 9 0 13 4 9 0 0 2
13 13 13 11 11 11 9 11 9 13 4 9 0 2
19 9 2 9 13 2 13 7 13 7 9 0 13 13 4 9 13 7 13 2
8 2 14 4 3 10 13 2 2
8 9 7 13 4 3 2 9 2
11 9 0 12 13 13 9 12 7 13 4 2
10 0 9 11 13 4 9 2 10 13 2
9 14 4 13 9 9 0 13 4 2
16 10 13 0 13 2 7 0 13 4 9 9 0 10 13 4 2
15 3 9 13 4 2 10 9 9 9 9 13 4 3 9 2
11 11 9 0 2 15 13 4 9 9 13 2
8 9 0 9 13 4 3 7 2
13 11 2 13 9 12 9 9 13 4 11 9 13 2
16 9 2 9 2 2 9 10 13 7 9 13 9 13 4 13 2
11 9 9 9 0 12 9 13 4 9 9 2
15 11 9 0 2 11 13 9 13 9 2 11 13 13 4 2
17 2 15 9 10 13 3 2 14 13 0 2 14 13 9 9 12 2
31 9 14 4 9 13 2 7 9 13 9 13 4 9 2 3 13 4 13 4 2 7 9 9 12 13 4 13 2 12 9 2
7 9 0 9 9 13 4 2
18 9 10 2 9 9 12 13 9 13 9 2 2 9 9 0 13 2 2
11 13 10 9 12 7 9 10 4 9 7 2
19 9 11 11 9 14 4 9 0 13 2 9 13 7 9 12 9 13 4 2
6 2 9 10 13 4 2
10 9 14 4 9 9 13 9 9 13 2
10 13 13 4 2 9 9 10 13 4 2
8 9 0 13 2 9 0 13 2
12 10 13 4 9 12 9 13 4 11 9 13 2
7 3 2 9 10 13 4 2
17 11 7 9 12 13 4 3 13 12 9 2 7 14 4 9 13 2
5 3 0 13 10 2
13 10 9 2 13 2 13 9 13 13 4 13 4 2
13 3 13 14 4 7 2 9 10 13 9 9 13 2
11 11 9 9 2 7 2 13 13 4 9 2
11 0 9 13 13 4 11 11 13 12 9 2
7 12 9 13 4 11 11 2
6 7 9 9 13 4 2
20 7 2 9 0 12 13 13 2 9 3 13 13 3 10 13 4 13 4 2 2
7 10 13 4 9 10 13 2
7 7 0 10 9 13 4 2
6 9 3 13 4 9 2
5 11 9 13 4 2
5 14 13 13 13 2
26 9 0 10 13 4 2 9 13 9 13 4 2 7 12 9 0 13 2 9 9 9 13 13 13 4 2
7 0 13 4 9 3 13 2
9 9 0 9 13 13 9 13 11 2
9 3 11 13 9 9 10 13 4 2
25 7 2 9 0 9 13 11 7 9 9 9 13 14 4 7 2 3 7 3 9 9 13 4 13 2
15 11 9 9 2 9 0 12 3 13 2 13 4 13 4 2
15 2 9 9 3 13 4 2 9 13 2 9 9 13 13 2
4 14 13 9 2
5 2 13 4 2 2
9 9 9 0 13 2 7 9 13 2
13 9 13 9 2 9 7 9 9 13 4 11 9 2
5 9 0 13 4 2
9 11 14 4 9 0 13 3 9 2
5 2 9 13 4 2
23 10 14 4 13 10 9 10 13 9 9 9 10 13 15 9 13 14 4 9 12 13 7 2
3 9 13 2
8 3 12 9 13 4 9 9 2
12 11 9 0 12 9 9 13 13 2 9 12 2
5 9 10 9 13 2
17 11 11 13 4 9 9 13 7 15 12 13 2 7 15 13 4 2
7 9 9 13 4 0 9 2
5 11 12 13 4 2
3 0 13 2
5 9 9 0 13 2
18 11 9 9 0 9 10 13 13 2 2 12 9 13 9 14 13 2 2
15 11 11 2 7 2 12 9 13 4 9 13 13 13 4 2
5 9 13 4 10 2
7 9 11 9 13 4 9 2
4 14 13 10 2
9 9 9 11 9 12 9 13 4 2
6 9 9 13 4 9 2
10 10 12 13 13 11 9 13 4 9 2
8 2 13 9 9 13 4 9 2
17 3 7 3 13 9 3 13 4 9 13 9 0 7 10 13 4 2
9 9 9 9 12 9 9 0 13 2
18 11 9 9 0 13 4 9 7 9 9 3 13 4 9 13 13 9 2
10 3 2 12 9 11 9 13 13 4 2
9 11 2 7 2 9 9 13 4 2
11 10 11 3 13 4 2 3 13 4 7 2
17 9 9 10 9 10 13 4 7 9 9 10 2 9 9 13 4 2
7 9 9 9 9 13 4 2
14 9 9 9 9 0 13 4 12 9 2 9 9 13 2
14 11 9 13 4 12 9 2 11 9 12 9 13 3 2
5 10 9 13 4 2
9 9 0 9 9 13 4 9 0 2
11 2 9 7 9 13 13 4 13 9 2 2
5 3 13 4 9 2
13 9 13 9 10 9 13 2 7 3 13 0 13 2
6 3 13 4 3 9 2
8 2 15 14 4 3 9 13 2
15 10 9 13 4 2 7 9 9 7 0 9 13 4 3 2
10 10 13 4 11 9 0 9 13 13 2
14 9 2 7 2 2 0 9 13 4 9 2 13 4 2
12 10 2 9 13 4 9 2 9 0 13 4 2
17 0 9 13 13 2 7 10 9 13 2 9 13 9 0 13 11 2
20 9 0 11 9 13 9 13 7 9 9 0 9 0 9 0 13 4 13 4 2
14 9 13 9 4 2 7 9 13 13 2 9 9 13 2
20 9 9 14 13 7 2 11 10 10 9 13 4 9 7 9 9 11 7 11 2
12 2 9 13 13 9 7 10 10 9 0 13 2
12 9 0 7 9 9 13 4 3 11 13 4 2
17 0 9 7 9 13 4 3 7 3 11 2 7 9 11 13 4 2
14 11 9 0 13 2 7 9 10 9 13 13 4 11 2
9 2 9 0 2 13 4 11 11 2
17 9 9 0 13 2 11 7 11 11 0 9 10 13 9 13 4 2
9 7 2 3 9 10 13 9 13 2
10 12 9 13 4 2 9 0 12 13 2
11 11 9 1 2 7 2 15 10 7 13 2
11 0 9 13 4 9 10 13 4 15 1 2
36 11 11 9 0 7 11 11 10 9 9 9 3 9 12 13 4 2 9 0 3 2 11 11 1 9 2 7 2 11 9 13 4 2 9 12 2
12 9 13 4 7 2 3 13 9 10 13 4 2
23 3 2 0 9 11 9 13 4 10 13 4 11 9 2 7 0 13 14 4 7 0 13 2
12 7 13 4 9 0 13 4 9 9 9 1 2
15 9 11 9 9 13 2 7 2 9 10 2 9 0 13 2
19 11 9 12 2 12 13 4 12 9 9 9 2 11 8 11 3 0 7 2
18 9 12 3 2 9 12 2 13 4 11 9 11 9 3 2 12 2 2
10 10 12 2 11 11 13 4 9 10 2
16 13 9 12 13 4 3 11 11 11 11 12 9 9 9 9 2
21 7 11 9 13 3 2 3 13 4 11 2 3 7 3 2 0 7 2 9 1 2
16 11 3 0 13 2 13 2 13 10 9 11 2 11 7 11 2
10 11 12 9 13 4 9 9 12 13 2
16 11 1 2 11 11 13 12 9 0 9 9 11 1 13 4 2
31 11 13 9 2 11 13 4 9 1 13 2 9 12 2 2 9 12 11 13 4 9 2 12 3 11 11 2 7 12 11 2
33 11 11 11 8 11 11 9 9 9 9 12 9 0 13 4 11 9 0 9 11 11 2 11 11 11 7 11 11 11 11 9 1 2
22 9 9 2 3 2 9 1 9 2 2 13 2 13 4 9 2 9 13 0 13 9 2
16 2 2 13 4 2 7 9 9 10 1 9 14 4 13 13 2
27 11 11 11 9 10 13 4 9 2 7 2 11 11 9 0 12 9 13 13 12 9 0 3 13 4 3 2
7 13 4 9 14 13 9 2
24 9 10 2 12 9 12 13 3 2 12 9 13 4 9 10 2 3 0 0 9 13 9 13 2
12 3 9 1 2 12 9 13 4 2 12 2 2
18 12 9 3 2 11 2 11 0 9 12 13 4 2 11 11 9 9 2
22 13 13 9 13 2 11 9 11 11 9 13 13 4 2 9 3 2 13 13 11 9 2
22 11 9 3 14 4 9 13 11 9 2 7 2 7 2 3 13 4 9 1 11 9 2
10 11 11 12 9 12 9 9 13 4 2
9 10 9 9 9 9 13 13 2 2
24 10 1 2 9 12 9 9 13 4 12 9 11 2 11 11 9 9 7 11 11 12 9 13 2
14 9 9 13 4 9 10 13 4 13 9 9 11 11 2
12 11 8 11 9 1 13 13 4 9 7 9 2
23 13 13 2 7 2 9 12 9 15 13 2 7 10 10 2 3 2 9 13 9 4 13 2
8 11 11 7 9 13 4 11 2
10 7 2 9 1 9 0 13 4 2 2
20 9 13 9 0 13 4 11 2 7 12 9 13 9 13 13 4 9 9 0 2
25 9 13 4 2 12 9 0 13 2 12 9 1 13 2 7 3 11 11 0 13 4 9 14 13 2
29 10 10 1 9 0 2 9 13 2 7 9 0 9 12 8 3 13 4 0 13 2 14 9 2 14 10 10 9 2
18 11 7 11 11 13 4 9 7 10 1 11 2 11 7 11 13 4 2
15 7 2 11 11 11 9 9 13 4 2 7 11 11 13 2
9 3 9 12 9 9 13 4 11 2
16 9 9 9 13 4 9 2 12 9 11 11 13 4 9 0 2
23 0 9 13 2 11 2 11 9 9 2 2 7 9 9 11 7 11 9 9 9 13 4 2
14 14 4 3 11 11 13 2 14 4 3 9 9 13 2
22 9 3 12 9 11 13 4 9 1 9 9 2 15 3 2 13 4 13 2 11 9 2
14 9 11 13 4 14 2 9 12 9 13 4 13 9 2
7 9 13 4 9 1 9 2
16 2 15 13 4 2 7 2 11 9 9 10 1 15 2 7 2
26 9 10 1 2 9 7 9 9 9 2 13 9 2 9 7 10 9 9 7 9 9 9 9 13 4 2
14 11 9 9 9 13 4 3 13 4 9 2 9 13 2
11 11 12 9 1 9 13 4 12 9 13 2
18 0 9 9 9 12 4 2 7 9 10 2 9 11 9 13 4 12 2
22 11 9 9 13 4 9 12 2 10 12 9 9 1 13 4 2 3 9 13 4 3 2
13 9 10 9 12 2 10 12 2 2 13 10 1 2
21 9 9 7 11 11 9 0 13 4 9 1 13 4 2 9 13 13 9 13 3 2
30 9 2 9 2 9 10 2 12 7 12 13 4 2 7 3 13 4 9 2 3 0 7 2 9 9 9 12 7 9 2
27 9 9 13 9 12 13 4 3 3 9 0 11 2 11 13 4 11 7 11 2 7 3 12 9 13 4 2
21 3 7 10 9 0 13 9 13 2 9 1 9 9 0 13 4 9 0 1 2 2
28 7 12 13 2 7 14 13 10 2 11 11 0 7 11 11 0 3 13 4 9 0 9 10 13 9 9 1 2
16 3 2 9 13 9 9 0 9 13 4 7 9 0 9 9 2
6 11 11 11 9 13 2
7 10 9 13 4 9 1 2
8 10 10 1 9 0 12 13 2
18 3 1 2 9 9 2 9 0 13 4 2 7 9 9 13 4 9 2
21 13 4 9 10 13 9 2 10 14 13 11 13 4 9 0 2 0 1 9 13 2
20 11 9 9 0 0 13 13 4 12 9 9 9 13 7 2 12 7 2 13 2
16 12 9 11 9 9 13 13 4 11 11 1 11 13 13 4 2
23 7 2 11 9 13 13 4 13 0 0 9 13 13 2 7 2 7 2 11 9 9 13 2
9 2 9 1 2 9 13 4 2 2
7 11 11 13 4 11 9 2
15 11 9 9 11 9 9 9 0 13 13 4 3 11 9 2
19 11 13 9 1 2 11 13 4 9 0 0 12 13 11 9 13 13 4 2
15 15 12 9 12 10 1 13 9 14 4 3 13 9 9 2
22 9 1 2 9 10 13 4 12 9 11 11 11 9 9 12 9 7 9 0 9 13 2
13 9 9 12 9 9 13 4 14 4 10 13 13 2
28 9 10 1 0 9 14 13 7 2 9 9 13 4 2 2 9 9 7 9 3 9 0 1 13 4 13 4 2
18 2 9 3 13 4 2 7 3 8 9 0 13 4 2 12 9 0 2
18 13 4 9 11 2 11 2 9 13 12 9 0 9 1 3 13 4 2
27 9 1 2 9 13 4 11 11 2 11 2 11 2 11 2 11 2 11 11 9 2 11 7 11 9 9 2
26 3 3 2 11 9 10 13 4 0 9 9 0 13 2 7 13 13 9 10 13 3 0 13 4 10 2
28 7 2 11 11 7 11 11 11 7 11 9 9 13 4 11 14 13 3 11 9 9 2 11 9 9 9 7 2
19 13 9 1 13 4 9 0 9 9 2 9 2 9 7 9 0 13 3 2
27 11 11 9 7 2 0 13 4 2 9 12 9 13 4 13 3 11 7 3 10 9 0 14 13 13 4 2
12 15 9 11 1 13 4 9 9 10 0 13 2
17 9 13 4 9 13 9 13 2 3 4 13 9 9 11 9 13 2
11 9 0 9 0 9 9 9 13 9 13 2
19 7 2 11 9 0 11 11 9 9 9 9 1 15 9 13 4 13 4 2
18 10 9 9 13 2 3 2 9 12 1 13 2 9 13 4 13 4 2
16 9 9 10 11 1 9 1 13 4 2 7 9 10 9 13 2
20 9 9 12 9 14 4 9 0 13 2 11 7 11 1 3 13 4 9 9 2
16 9 9 2 0 13 9 13 10 2 3 1 3 3 13 4 2
12 9 13 14 4 3 13 2 3 13 3 10 2
12 9 9 9 14 13 9 13 4 2 12 12 2
5 11 14 2 13 2
12 9 9 9 2 7 2 9 9 9 13 4 2
23 11 2 7 2 9 13 7 9 13 13 2 2 11 9 9 10 13 2 13 4 13 9 2
20 15 9 0 3 13 9 13 9 13 4 2 7 10 14 4 13 15 13 9 2
24 7 2 3 3 2 9 0 9 0 13 2 11 9 11 9 9 13 4 9 3 13 4 3 2
9 9 13 13 9 0 13 4 11 2
18 12 9 1 13 12 9 9 0 9 2 10 12 9 0 13 13 4 2
7 11 1 13 4 3 11 2
24 11 9 12 1 13 4 13 4 3 2 3 2 9 13 4 7 15 10 9 9 13 13 4 2
11 3 3 2 9 10 3 7 13 4 9 2
12 9 10 2 9 1 9 9 14 13 13 4 2
19 11 11 9 9 13 7 12 9 9 0 1 12 9 13 4 9 11 0 2
12 12 9 0 7 12 9 13 4 9 0 9 2
17 9 9 9 9 9 13 13 13 4 2 9 2 9 9 9 9 2
7 9 1 9 0 13 13 2
17 11 9 11 11 1 2 7 11 9 11 11 1 2 9 13 4 2
9 9 11 1 13 13 4 0 9 2
9 11 9 12 12 9 9 13 4 2
19 12 9 1 2 11 9 9 7 9 10 13 13 9 12 9 13 9 12 2
10 9 0 11 9 13 4 0 9 1 2
20 10 10 1 2 9 13 9 13 9 9 9 2 9 7 9 0 13 4 13 2
19 3 2 14 4 13 11 11 3 13 4 2 9 7 3 2 9 0 12 2
39 13 4 2 9 10 2 9 2 9 13 9 9 7 2 10 9 2 9 9 13 4 10 2 9 12 9 1 13 14 13 7 2 7 2 9 14 13 2 2
12 11 11 11 9 9 9 13 4 11 9 10 2
19 9 10 11 9 11 9 11 9 11 9 9 13 7 13 9 13 13 4 2
8 11 15 13 4 3 13 4 2
21 9 11 9 9 9 13 4 7 2 11 9 14 7 2 9 13 10 12 13 4 2
12 9 1 2 9 13 4 3 7 9 9 0 2
11 9 1 0 13 2 7 9 0 13 2 2
10 3 9 10 11 9 12 9 13 4 2
18 11 11 11 9 9 3 13 13 4 3 9 9 9 13 4 9 0 2
7 2 9 9 12 13 2 2
9 12 11 11 13 4 2 12 5 2
16 11 0 9 0 13 4 11 1 2 7 11 9 13 13 9 2
9 3 2 12 1 9 10 13 4 2
10 9 9 13 11 11 11 13 3 13 2
17 11 11 7 11 9 11 11 11 13 11 9 9 13 4 12 9 2
9 11 11 11 9 0 13 4 11 2
13 11 9 2 9 1 4 13 2 15 13 4 9 2
16 12 9 1 13 4 9 9 9 7 8 9 13 4 11 9 2
22 2 3 2 0 13 4 11 13 7 11 2 11 7 11 1 9 0 13 2 3 13 2
17 2 3 7 3 13 9 13 10 9 13 2 11 9 9 1 2 2
26 9 9 13 4 2 10 9 13 4 3 3 2 9 10 13 4 9 2 9 0 9 3 13 4 9 2
13 9 14 4 13 9 3 1 9 11 13 12 9 2
13 9 10 2 11 11 9 12 9 9 13 4 10 2
15 9 7 2 9 13 2 15 9 8 0 13 4 9 10 2
8 9 10 13 4 11 11 11 2
14 15 3 9 0 13 4 2 12 7 9 9 9 2 2
21 11 11 9 9 9 7 9 1 9 13 4 2 11 13 9 9 9 0 13 4 2
15 9 9 9 2 3 9 0 7 9 0 9 10 13 4 2
24 11 9 3 2 9 13 9 14 4 13 2 7 9 15 10 13 7 9 0 13 4 9 2 2
19 11 13 4 9 2 11 9 10 0 1 13 9 13 9 13 9 13 4 2
12 11 0 11 13 4 3 9 13 2 9 1 2
6 9 9 1 13 4 2
35 11 11 9 0 7 14 4 3 0 9 13 2 7 4 12 9 13 9 2 11 11 2 11 11 2 11 11 2 2 12 11 9 9 13 2
12 11 11 9 0 9 13 4 9 9 13 9 2
5 7 10 9 13 2
26 11 9 9 12 13 13 3 2 12 9 0 13 4 13 4 9 2 11 9 1 2 11 12 9 9 2
19 9 10 13 4 9 0 2 11 9 12 13 4 2 9 0 13 9 13 2
10 7 2 0 13 13 10 9 13 4 2
17 9 12 2 11 11 9 12 9 2 12 9 13 4 9 12 9 2
11 9 10 13 9 1 13 9 13 13 4 2
6 13 15 1 13 4 2
16 9 10 9 0 11 7 11 9 9 1 13 9 3 13 4 2
25 9 13 9 14 4 13 10 9 2 7 3 9 12 1 2 13 13 4 12 10 13 9 7 9 2
7 9 9 1 13 4 11 2
10 13 11 13 4 3 9 9 0 13 2
20 12 9 10 15 3 13 4 15 2 7 9 10 2 15 7 3 13 4 15 2
7 7 11 11 9 13 9 2
10 11 11 13 13 4 10 9 13 3 2
6 9 2 13 4 13 2
16 9 1 2 13 2 13 4 11 11 9 0 13 0 4 9 2
16 9 1 9 7 9 9 1 13 11 9 13 4 9 13 11 2
24 9 10 12 9 13 12 9 13 4 2 7 9 10 14 4 11 11 9 13 2 11 11 7 2
11 11 11 7 11 11 13 4 11 13 9 2
6 9 1 13 4 9 2
14 3 1 12 7 9 13 13 4 9 10 3 13 4 2
28 2 9 13 4 2 10 13 4 2 10 2 3 2 15 9 13 2 2 9 1 2 11 2 13 4 3 2 2
13 9 11 2 9 12 2 11 12 9 13 4 3 2
24 11 9 13 2 7 2 11 0 4 2 7 9 9 1 13 2 9 13 4 9 12 9 9 2
8 11 11 14 4 9 1 13 2
24 11 9 11 13 4 9 9 0 13 4 11 9 2 7 3 9 11 13 4 2 12 9 9 2
27 9 10 1 7 11 9 13 4 11 9 0 7 0 13 4 9 9 14 4 10 13 11 9 12 9 9 2
23 13 4 9 10 13 4 2 7 3 13 4 2 9 13 2 9 1 9 0 10 9 13 2
39 11 11 11 3 9 0 13 4 11 13 12 9 2 12 9 9 1 2 2 7 14 4 3 13 12 9 13 9 2 7 2 9 2 9 9 13 4 9 2
38 3 2 11 9 12 2 9 2 11 1 13 4 2 11 2 9 12 2 9 2 11 1 13 4 2 12 9 2 7 12 2 9 2 11 1 2 9 2
16 9 10 2 11 0 9 0 2 11 11 2 9 0 13 4 2
17 9 3 13 13 11 9 9 12 2 7 15 0 9 13 9 13 2
8 11 11 11 9 13 4 3 2
30 9 13 0 7 11 9 9 13 11 11 9 13 4 2 3 13 9 13 14 4 2 9 7 9 13 13 4 13 9 2
32 11 11 11 11 9 1 9 13 4 2 9 0 2 0 7 0 2 9 0 2 13 7 9 0 8 9 2 0 2 13 4 2
19 9 14 4 9 9 13 2 3 3 4 13 3 2 7 3 2 3 9 2
12 10 9 13 11 11 2 3 2 0 9 9 2
15 3 2 11 11 11 9 9 13 13 4 11 9 0 13 2
20 11 12 7 11 12 13 4 3 2 7 9 11 0 1 13 13 4 0 9 2
22 13 9 13 9 9 13 4 13 9 9 2 3 3 11 2 11 2 11 11 7 11 2
12 12 9 3 13 4 12 9 1 13 4 9 2
5 3 9 13 4 2
13 9 11 11 9 9 9 9 13 14 4 13 4 2
18 9 9 0 9 13 13 4 2 11 9 9 0 11 11 13 4 9 2
19 2 10 2 3 0 2 9 7 9 3 13 4 9 0 7 0 9 2 2
24 11 11 12 9 12 11 9 13 4 9 13 9 13 4 9 2 7 12 9 10 13 4 9 2
25 7 10 9 2 11 2 9 2 13 4 10 9 13 4 2 9 9 7 9 2 13 2 9 3 2
8 2 0 13 4 2 9 1 2
20 7 2 3 13 4 3 11 11 11 13 4 2 12 9 3 2 11 9 9 2
13 9 7 9 10 9 13 4 13 12 9 0 9 2
16 12 12 9 2 9 0 1 13 4 9 1 2 9 13 9 2
16 9 0 13 2 7 12 1 13 4 9 2 3 12 9 13 2
7 11 11 12 9 13 4 2
15 12 9 9 7 2 12 9 13 12 9 0 9 13 9 2
14 9 9 7 9 10 2 9 0 1 2 13 13 4 2
8 12 7 12 9 13 9 13 2
11 3 7 14 13 0 11 9 11 9 13 2
13 3 9 13 11 13 7 2 9 10 13 4 11 2
7 15 13 10 13 7 13 2
9 11 12 13 4 11 1 2 9 2
11 2 9 0 1 9 0 13 4 9 13 2
8 9 11 9 0 4 13 13 2
11 2 10 13 9 13 10 12 1 13 4 2
9 9 3 2 12 9 9 13 9 2
15 10 3 14 13 13 4 11 9 7 13 4 3 9 2 2
19 11 11 9 11 11 13 4 11 11 9 2 7 10 9 9 9 12 13 2
16 9 13 4 11 9 0 2 7 3 13 4 12 9 9 0 2
14 9 9 0 9 9 0 13 4 9 9 2 9 1 2
10 3 9 0 13 4 2 10 14 10 2
15 0 3 2 9 13 4 10 9 8 9 10 10 13 4 2
11 3 2 11 11 11 13 4 11 11 0 2
22 2 9 2 13 4 11 11 11 2 7 11 9 2 9 9 3 0 2 13 13 4 2
27 11 12 7 11 0 9 13 4 9 11 12 7 11 1 2 9 10 13 13 7 2 12 2 12 9 2 2
12 9 13 9 1 9 13 7 9 13 13 4 2
14 9 0 1 2 9 9 10 9 7 9 0 13 13 2
11 3 0 13 7 9 9 13 4 10 1 2
20 9 0 13 4 2 9 9 9 9 3 13 7 9 3 2 13 9 13 4 2
17 7 2 11 11 11 13 4 7 3 7 3 13 11 11 11 13 2
17 2 9 0 12 1 13 7 13 13 9 13 11 11 15 13 9 2
12 13 4 9 9 13 2 9 2 9 7 9 2
6 15 1 13 3 13 2
16 7 9 10 13 4 11 13 7 11 11 13 4 9 10 13 2
10 9 9 13 4 11 12 9 12 9 2
13 13 4 9 13 4 9 9 0 7 9 0 1 2
23 11 11 0 2 7 2 3 3 13 4 9 11 13 9 7 3 3 0 9 1 13 4 2
26 11 9 9 0 9 1 2 11 9 7 12 9 9 9 14 4 11 9 3 3 9 0 7 0 13 2
18 3 3 9 10 9 10 13 4 2 7 9 9 7 14 13 13 9 2
13 9 0 13 15 1 7 9 3 13 4 9 9 2
13 13 9 1 7 12 9 7 3 13 4 9 9 2
16 9 9 3 13 7 9 3 13 9 13 2 7 9 10 3 2
25 11 9 9 1 9 13 4 2 7 9 10 2 9 0 12 2 11 1 13 9 0 13 13 4 2
13 10 1 2 14 13 13 9 9 13 13 0 9 2
13 9 1 13 4 11 7 11 2 12 9 13 13 2
17 9 2 11 11 7 11 11 9 9 12 9 13 3 13 4 9 2
15 11 2 11 2 11 7 9 11 7 3 9 13 13 4 2
20 7 2 9 3 13 4 13 2 9 9 0 13 7 9 0 13 13 11 2 2
11 7 2 9 2 3 7 13 9 13 11 2
12 11 9 13 7 9 1 9 0 13 13 3 2
18 11 11 9 1 2 12 9 9 0 4 9 9 9 13 3 9 13 2
8 13 9 13 2 10 9 1 2
13 9 0 13 4 13 11 2 12 12 9 0 7 2
21 11 1 2 11 11 11 9 7 0 13 4 9 11 9 9 13 2 9 0 13 2
16 3 11 11 13 4 2 9 1 2 7 11 9 12 13 4 2
14 11 11 9 7 9 1 13 4 2 2 0 2 13 2
23 3 11 11 7 11 11 9 13 4 2 7 3 7 12 9 13 4 3 13 4 10 9 2
25 11 2 9 9 2 11 2 11 2 9 11 2 11 2 11 2 11 2 11 7 11 13 4 9 2
11 9 0 13 2 9 9 0 13 13 4 2
22 9 9 9 2 11 9 13 4 9 2 7 12 9 9 13 3 9 9 9 3 13 2
20 9 13 4 3 7 3 2 7 12 9 13 4 11 2 11 2 11 7 11 2
5 14 3 13 7 2
18 3 2 9 9 10 2 9 10 2 13 2 4 0 9 3 13 4 2
7 9 3 13 7 9 0 2
16 9 10 9 0 13 11 2 7 14 13 9 9 0 7 9 2
24 15 9 0 2 9 13 4 2 9 13 9 13 4 2 3 9 9 2 7 3 7 9 13 2
8 12 0 9 9 0 9 13 2
30 11 9 1 2 9 12 9 0 2 11 11 11 2 11 11 11 7 11 11 2 13 13 4 13 12 9 11 13 4 2
13 11 9 11 11 2 7 2 3 13 4 9 9 2
17 12 1 2 7 2 9 13 13 13 7 9 9 9 0 13 0 2
11 11 11 7 13 13 4 11 2 10 9 2
21 9 9 2 7 9 9 9 2 11 2 9 13 9 13 4 12 11 9 9 11 2
12 11 9 9 12 9 0 13 4 11 0 9 2
8 13 4 13 13 9 9 1 2
21 9 9 9 11 13 4 12 9 4 7 2 11 11 2 3 12 9 7 13 4 2
25 11 9 9 9 11 11 11 9 11 11 11 9 9 13 4 9 2 7 10 1 11 11 13 4 2
16 13 2 9 9 13 9 2 9 9 13 4 7 9 13 4 2
16 13 7 2 14 13 10 2 13 4 9 0 2 9 13 4 2
11 11 9 9 13 13 4 11 1 9 9 2
22 3 13 12 9 9 13 4 2 7 7 2 9 13 13 4 9 0 9 13 4 9 2
15 11 7 11 11 9 9 9 9 11 11 9 9 13 4 2
6 9 9 9 13 4 2
14 11 11 11 11 11 13 4 2 3 0 2 11 13 2
9 3 13 4 11 12 9 9 9 2
19 10 2 11 13 4 9 11 9 14 7 2 11 9 13 7 13 9 13 2
21 9 13 4 9 3 13 4 9 2 9 2 9 2 9 2 9 7 9 1 9 2
18 3 13 4 9 12 9 1 12 9 2 7 11 13 4 9 7 0 2
14 11 9 0 9 13 4 2 7 11 9 13 4 13 2
31 11 9 13 2 9 9 12 9 0 10 13 13 4 7 10 15 9 3 13 4 2 9 13 2 3 15 13 4 13 3 2
10 15 13 9 1 13 2 9 11 1 2
10 11 9 13 13 9 0 9 0 9 2
16 10 2 3 13 4 9 9 3 13 12 9 2 11 9 1 2
17 11 9 14 4 3 0 13 11 2 14 4 3 11 11 9 13 2
27 9 9 2 11 9 13 9 11 0 13 13 4 11 11 9 9 9 7 9 0 9 9 13 13 4 9 2
7 11 11 11 13 4 9 2
16 11 11 9 9 13 4 9 10 13 4 11 11 12 9 11 2
15 7 9 13 7 15 1 13 13 13 2 3 13 4 9 2
24 9 11 10 9 10 9 13 13 4 10 9 13 4 2 3 3 2 9 13 7 9 0 13 2
12 12 11 11 11 13 4 9 2 10 9 1 2
10 11 11 9 13 11 11 13 4 11 2
7 3 7 3 11 13 4 2
10 9 9 9 9 0 12 13 4 9 2
14 9 12 9 13 9 2 7 9 1 13 3 9 9 2
10 12 9 9 14 13 9 2 9 1 2
30 2 9 0 2 9 0 11 11 11 0 9 7 11 11 9 0 9 13 4 7 2 15 9 3 13 2 4 13 4 2
8 15 1 13 9 0 7 0 2
35 11 9 2 12 2 7 9 2 12 2 3 13 13 2 7 11 9 2 12 2 2 11 9 2 12 2 2 9 9 7 2 12 2 13 2
24 9 10 13 4 13 11 11 9 0 9 9 0 9 9 12 9 13 4 13 4 13 4 9 2
15 9 9 7 9 1 9 0 7 0 2 9 9 13 13 2
12 9 9 10 13 13 4 7 3 3 13 4 2
12 9 10 2 9 14 7 2 9 7 13 4 2
13 14 4 11 11 9 13 12 7 9 11 9 9 2
6 11 11 9 13 4 2
15 3 13 4 9 0 10 2 7 13 13 2 15 9 1 2
13 11 11 7 11 11 9 13 4 11 12 9 13 2
17 2 9 13 2 9 3 8 3 13 13 4 9 9 13 2 2 2
39 3 9 11 9 12 13 4 0 9 13 2 7 9 12 9 9 9 13 13 4 10 9 2 9 2 9 0 2 9 2 2 13 4 3 9 13 4 9 2
23 9 11 9 11 9 9 13 11 9 9 2 10 9 7 9 9 1 0 9 12 13 4 2
16 3 2 11 12 9 1 2 9 13 9 1 13 4 9 10 2
25 3 2 11 11 11 2 9 13 9 9 2 13 13 4 3 2 2 10 13 13 4 9 0 2 2
23 2 9 9 9 2 9 2 7 2 9 0 2 9 2 9 2 6 9 7 9 13 4 2
8 3 7 9 0 13 4 13 2
5 9 13 0 4 2
20 0 11 14 13 9 3 9 2 9 9 9 10 15 13 4 2 9 9 12 2
13 9 0 12 2 7 9 12 13 4 9 9 12 2
20 11 11 9 9 13 4 13 9 10 11 2 7 11 9 0 13 4 12 9 2
17 9 13 9 1 2 12 9 9 12 9 9 13 4 11 9 9 2
13 11 9 9 0 1 13 2 11 10 13 3 13 2
30 9 0 13 11 1 9 12 9 9 13 2 7 2 10 1 2 9 7 9 9 13 2 7 3 0 9 0 13 4 2
15 12 9 1 13 9 13 9 11 11 9 9 9 12 1 2
10 11 9 13 4 11 9 1 9 10 2
14 9 0 9 11 11 7 11 11 3 13 4 12 9 2
15 2 9 9 2 13 4 3 11 9 2 9 0 12 1 2
9 3 13 12 9 11 13 2 13 2
19 3 2 11 7 11 7 9 13 4 13 11 9 13 4 12 9 13 3 2
26 10 9 2 0 9 9 1 2 10 9 13 4 2 3 3 9 2 9 7 10 1 13 4 9 0 2
17 3 2 13 9 13 2 11 1 13 4 3 11 9 11 9 0 2
8 2 13 9 3 13 12 13 2
14 9 3 2 7 2 3 9 0 13 4 0 1 9 2
25 9 13 4 9 9 9 0 13 2 7 2 7 2 14 13 9 11 9 11 9 13 4 9 0 2
25 11 11 0 2 7 2 9 13 4 9 3 9 10 9 13 4 7 3 3 13 4 2 9 1 2
7 12 9 9 11 13 4 2
21 13 7 9 13 13 4 9 0 13 3 15 9 13 7 9 12 9 9 9 13 2
8 11 11 11 12 9 13 4 2
10 11 11 2 0 2 13 4 11 9 2
19 9 13 4 2 0 9 2 9 9 12 2 9 0 13 9 10 13 4 2
8 11 11 11 3 13 4 11 2
16 7 2 11 7 11 9 9 9 13 7 3 9 1 13 4 2
28 11 9 1 13 4 9 9 7 9 2 7 11 9 1 13 9 3 13 4 9 2 7 0 9 14 4 13 2
17 11 11 13 4 9 9 1 2 7 11 7 11 0 1 9 9 2
17 3 2 9 1 10 9 13 4 2 7 9 3 3 13 9 13 2
30 11 13 4 9 12 9 13 9 9 1 2 7 12 9 13 4 9 2 11 0 9 13 2 11 9 13 4 9 13 2
15 12 9 0 13 9 13 13 4 9 11 9 9 11 11 2
18 3 2 9 13 2 9 0 1 13 12 12 9 9 13 9 13 4 2
29 11 2 7 2 2 13 4 12 7 12 9 9 13 2 13 4 13 4 2 9 10 1 9 12 13 4 9 13 2
18 2 11 11 2 11 11 8 11 2 11 11 7 11 11 9 0 13 2
18 11 9 7 9 13 4 11 7 11 9 2 9 9 1 2 13 4 2
15 3 0 13 4 11 11 2 3 2 11 11 0 9 13 2
13 9 9 9 9 4 13 9 9 13 3 2 11 2
13 9 13 3 13 11 11 9 2 12 9 13 4 2
18 7 2 9 13 3 2 13 4 3 13 9 9 3 9 12 13 4 2
19 9 9 9 9 9 2 12 9 13 4 3 9 1 13 7 0 13 9 2
10 2 9 9 13 7 9 13 9 13 2
21 11 11 9 3 13 7 3 9 7 9 9 0 9 12 13 9 13 11 9 11 2
30 11 9 14 4 9 0 13 9 13 11 9 11 11 9 0 1 13 9 1 2 3 9 0 9 12 13 4 9 13 2
15 9 0 13 4 9 13 2 7 9 0 15 10 13 4 2
13 3 13 3 13 9 9 0 1 13 9 13 4 2
23 12 9 1 2 9 0 12 13 4 2 7 11 11 9 9 1 13 4 9 0 13 4 2
12 11 9 13 4 2 12 9 11 11 13 13 2
25 9 12 12 7 12 9 13 4 13 4 9 0 2 7 9 0 13 4 11 9 12 13 4 9 2
15 2 9 10 13 4 2 9 10 13 7 15 7 14 2 2
18 9 12 2 9 2 11 7 11 9 2 9 7 9 0 13 9 13 2
11 9 7 9 0 1 2 12 9 9 13 2
22 9 0 9 11 11 9 1 9 9 13 13 4 2 3 7 2 9 0 2 13 13 2
22 11 9 13 2 7 2 11 9 13 9 13 2 7 10 9 13 4 3 11 11 9 2
21 7 10 9 0 13 4 2 9 1 13 9 13 7 9 9 9 0 13 9 2 2
20 3 13 9 13 13 4 2 7 3 3 1 10 12 13 4 9 1 13 9 2
14 9 13 3 2 3 13 7 3 13 9 13 9 9 2
10 11 9 9 7 13 4 9 9 10 2
12 9 13 2 11 11 11 9 13 4 3 9 2
16 11 9 0 0 12 9 9 13 3 2 9 9 13 4 11 2
12 0 9 9 1 13 4 2 11 12 13 4 2
14 9 13 9 9 8 0 13 4 9 13 9 0 9 2
7 9 9 12 1 13 4 2
12 9 10 9 13 13 12 9 11 11 9 9 2
15 2 3 3 2 9 0 12 9 10 9 12 13 4 2 2
10 2 12 7 2 9 9 14 4 13 2
7 11 11 13 10 9 9 2
15 9 11 9 9 0 12 7 0 9 13 11 11 13 4 2
26 11 11 9 9 13 4 9 1 13 9 2 7 2 11 7 11 11 3 9 0 2 13 4 13 4 2
15 9 13 3 13 13 4 2 9 12 11 11 1 3 0 2
16 11 1 13 9 0 9 0 13 13 2 7 2 11 9 11 2
12 11 11 13 4 9 0 13 4 11 1 9 2
9 12 9 4 13 13 11 11 11 2
13 11 3 13 4 11 9 1 7 14 4 9 13 2
14 11 1 2 11 9 11 4 9 12 9 13 4 13 2
19 9 9 13 4 11 11 11 12 9 9 13 2 7 9 9 13 4 3 2
21 11 11 0 13 4 3 2 3 13 15 9 0 0 13 2 7 9 9 9 0 2
20 3 13 4 2 11 0 9 0 9 12 13 4 2 11 11 9 2 9 12 2
36 9 0 9 9 0 2 9 14 4 3 9 0 13 9 13 2 9 0 10 9 13 3 13 4 2 9 3 13 7 2 9 13 4 3 9 2
11 12 9 13 4 2 9 9 0 0 12 2
23 9 2 11 2 13 10 2 13 0 13 9 9 13 7 9 1 10 9 0 9 13 4 2
21 9 1 2 7 2 9 9 9 13 4 13 11 2 7 2 9 2 9 13 4 2
9 10 1 2 9 12 13 4 9 2
9 9 2 11 11 13 4 9 9 2
13 14 4 3 13 9 13 10 9 13 9 7 9 2
11 3 2 11 11 9 12 9 13 4 11 2
10 2 15 9 3 1 13 4 13 13 2
11 12 9 1 2 9 7 13 4 2 3 2
16 3 2 13 13 4 2 12 7 9 13 9 13 13 4 9 2
15 14 9 13 2 9 13 4 2 7 10 3 13 4 13 2
11 9 10 13 4 9 9 9 9 12 9 2
13 9 10 2 11 1 9 10 7 13 4 13 9 2
15 11 11 9 12 2 9 7 9 1 13 4 11 9 9 2
10 11 2 9 2 13 4 11 1 9 2
31 3 2 9 0 3 3 0 2 9 13 7 13 3 13 4 2 7 15 2 12 9 2 14 4 10 9 13 13 9 13 2
19 11 10 12 9 13 4 12 9 2 9 1 3 7 3 13 4 9 13 2
11 9 13 4 2 7 14 9 1 2 9 2
26 0 10 9 9 9 14 13 2 9 13 0 9 9 7 2 9 0 2 9 0 1 9 0 9 13 2
14 9 1 2 13 9 12 13 4 3 3 11 9 0 2
25 11 9 14 13 9 2 15 13 4 9 12 9 13 2 3 7 2 9 0 7 0 13 4 13 2
16 9 0 9 9 12 13 4 3 9 2 7 14 4 9 13 2
16 9 13 11 9 0 13 4 9 2 11 9 7 11 9 9 2
12 9 0 9 13 9 7 0 13 4 12 9 2
28 9 10 10 9 13 4 9 10 11 9 2 12 2 9 1 13 4 11 9 12 9 9 2 13 4 9 9 2
17 11 11 9 3 13 4 9 7 9 0 9 0 9 13 9 13 2
8 10 9 2 10 9 13 4 2
23 9 2 15 9 2 9 0 10 13 13 7 9 10 2 10 9 1 2 9 0 13 13 2
9 2 9 13 3 13 13 9 13 2
23 7 9 14 4 3 13 7 9 12 2 3 1 13 3 2 9 0 13 13 4 2 7 2
18 9 10 9 1 13 9 12 9 9 13 4 9 2 13 3 4 13 2
18 0 9 2 9 9 1 2 0 11 13 9 13 4 2 11 9 0 2
13 11 0 7 11 8 12 9 9 0 13 13 4 2
25 9 0 9 10 2 0 2 3 7 3 9 9 0 13 9 13 2 7 2 9 2 9 9 13 2
17 12 9 9 7 9 9 9 13 13 9 3 11 2 11 1 9 2
14 12 3 2 11 9 9 9 0 12 9 13 4 3 2
19 11 1 11 0 4 13 2 7 15 9 11 7 11 10 9 0 13 4 2
23 11 13 9 2 11 9 2 9 12 2 7 0 9 0 2 9 12 2 13 13 11 11 2
12 13 13 3 11 9 9 11 13 4 9 0 2
17 7 11 9 11 13 7 11 9 13 4 2 9 1 13 4 3 2
6 9 0 13 4 7 2
8 7 9 1 13 9 13 4 2
18 9 1 2 9 10 3 11 9 9 12 12 9 9 13 9 13 4 2
9 9 13 4 11 11 12 12 9 2
26 11 11 13 9 13 4 11 9 12 9 0 0 13 13 2 7 9 0 3 13 7 0 12 13 4 2
10 10 1 9 7 11 13 13 4 3 2
27 7 15 10 9 9 13 13 9 13 2 9 13 9 13 4 9 2 9 8 0 13 7 10 9 0 13 2
27 9 9 0 9 13 13 4 3 2 7 9 1 7 2 14 4 0 9 13 2 7 14 13 11 1 9 2
21 0 10 2 9 9 9 0 13 9 9 9 1 2 7 3 0 2 13 4 9 2
16 7 0 14 4 9 13 2 9 13 2 9 12 1 13 9 2
8 11 11 13 9 13 4 9 2
21 11 11 11 13 4 9 10 13 12 9 9 0 2 11 9 13 4 9 0 2 2
11 11 11 9 13 4 3 9 2 9 13 2
21 11 9 2 11 9 2 3 0 13 2 7 11 13 4 9 1 13 13 4 2 2
21 11 9 9 10 12 12 9 0 13 2 7 9 10 9 0 13 11 9 13 9 2
7 9 10 13 4 11 11 2
23 11 9 9 13 9 13 4 2 7 3 7 2 13 13 4 3 10 9 13 9 13 4 2
28 11 7 11 9 1 9 13 9 13 2 3 9 10 11 11 9 11 9 7 11 11 9 11 9 9 13 4 2
20 3 2 9 11 9 1 13 3 13 13 4 9 2 7 3 2 13 13 4 2
23 9 10 0 13 4 13 4 11 2 7 11 7 3 13 0 13 9 0 0 7 0 13 2
30 9 11 0 11 11 9 2 11 11 11 0 2 11 11 0 7 11 11 0 13 13 4 0 9 12 9 9 9 0 2
14 9 9 13 3 2 12 9 1 9 13 4 9 11 2
10 9 10 2 9 9 9 3 13 4 2
15 14 13 2 3 3 2 0 9 0 7 0 13 9 0 2
18 9 0 2 7 2 13 13 4 9 9 9 9 13 4 13 9 9 2
21 11 9 13 7 13 2 9 1 2 9 2 9 0 10 1 2 9 0 10 1 2
13 3 7 3 13 4 9 10 13 13 9 12 9 2
6 9 13 9 9 13 2
12 10 1 2 9 9 9 12 9 9 13 4 2
15 11 11 11 9 9 7 9 13 4 11 11 9 3 13 2
18 7 2 9 13 4 0 10 0 13 2 12 12 7 12 9 1 13 2
21 7 13 4 9 0 12 9 9 0 10 1 2 9 0 7 9 0 1 2 7 2
12 3 13 2 7 2 9 2 11 2 9 12 2
19 9 0 1 10 9 10 13 9 0 2 7 2 9 0 3 13 9 13 2
10 10 10 9 9 13 2 7 11 14 2
22 12 9 9 12 13 4 2 7 3 9 13 4 11 12 7 11 2 7 11 7 11 2
28 13 4 9 9 2 9 2 9 2 9 9 2 9 9 7 9 2 9 9 2 9 2 9 2 9 7 9 2
34 9 10 2 9 9 7 9 9 2 9 9 9 1 9 13 9 13 7 10 13 4 2 9 0 13 4 2 3 13 4 13 7 13 2
15 9 10 1 11 10 9 13 4 2 9 9 0 13 4 2
16 14 13 3 0 2 9 9 12 15 13 4 3 3 13 9 2
16 9 12 12 0 13 4 2 10 0 11 9 2 9 13 13 2
9 12 9 9 9 13 4 13 4 2
16 9 10 9 3 2 11 11 9 9 9 3 13 9 13 4 2
14 11 9 10 9 13 4 13 7 13 9 12 9 13 2
21 7 2 2 9 1 9 2 13 4 7 2 9 3 7 3 13 4 13 11 9 2
12 0 9 13 9 2 11 11 9 9 13 4 2
29 11 9 9 1 9 13 4 2 9 13 2 7 11 2 11 11 9 1 2 13 4 2 9 7 9 0 2 13 2
16 9 13 4 9 10 9 2 9 13 2 9 1 13 9 13 2
18 9 9 1 13 4 9 13 13 13 4 9 9 0 9 0 13 4 2
10 9 7 9 10 10 13 4 3 11 2
35 9 1 9 13 9 11 11 13 13 9 13 11 2 7 0 2 9 9 0 2 13 13 4 2 2 3 2 11 0 13 4 9 13 2 2
38 11 11 11 9 1 9 10 9 7 9 13 4 9 13 4 2 9 9 10 13 4 13 9 9 1 13 2 7 10 9 10 9 13 14 4 13 4 2
19 11 11 9 13 4 2 2 11 11 7 11 11 9 0 9 2 13 13 2
15 3 1 9 9 4 13 12 9 13 13 4 9 10 13 2
16 11 9 9 1 2 9 12 9 13 4 9 7 10 12 9 2
17 11 9 9 13 4 11 9 11 9 0 1 13 12 9 9 9 2
21 11 13 4 2 12 9 9 0 13 9 13 9 12 11 9 13 13 4 9 10 2
16 9 9 15 3 13 13 2 7 9 3 13 4 9 7 9 2
12 14 2 7 10 9 0 13 0 9 9 3 2
35 0 9 9 13 4 13 9 1 13 4 10 9 2 0 7 9 9 2 13 4 9 14 4 9 9 0 13 7 3 9 0 10 13 4 2
36 9 2 0 9 1 2 9 9 13 9 2 9 1 3 11 9 13 4 3 11 8 8 11 2 11 11 13 2 13 4 9 11 13 4 9 2
20 13 4 9 11 11 9 13 4 9 2 9 3 13 0 9 13 14 4 7 2
10 9 9 10 14 13 3 0 15 1 2
33 9 13 14 13 9 10 9 12 12 13 2 11 7 11 14 4 13 3 2 7 2 11 11 7 11 11 11 12 13 4 12 13 2
8 10 9 12 13 11 11 7 2
13 12 12 9 9 3 13 4 9 12 1 13 4 2
30 11 1 2 9 12 1 9 2 14 4 0 13 2 2 7 12 13 4 2 9 13 9 7 11 9 2 13 13 4 2
14 11 11 11 9 9 9 1 2 0 13 4 3 13 2
17 9 13 9 9 7 9 9 12 13 9 13 9 1 13 9 13 2
6 7 7 10 13 4 2
19 0 13 9 7 9 0 13 2 9 9 10 11 2 9 10 11 7 11 2
22 9 10 13 4 9 10 2 7 2 9 7 9 1 13 7 2 0 13 3 13 13 2
16 2 11 11 2 11 11 13 4 2 11 7 11 13 4 11 2
11 11 2 9 1 9 2 13 4 9 9 2
10 10 3 13 4 11 11 0 9 13 2
11 9 13 4 13 9 9 13 9 0 12 2
12 3 3 2 9 10 12 12 9 13 11 9 2
28 7 2 12 12 9 9 7 9 1 9 9 13 4 11 9 10 9 2 11 9 2 14 4 3 9 1 13 2
21 11 9 9 2 11 2 11 7 11 9 9 13 4 2 3 11 9 13 9 1 2
14 2 13 9 10 2 7 12 7 2 14 13 0 2 2
18 3 2 11 11 11 9 13 4 9 10 13 2 7 10 9 13 4 2
20 11 11 11 9 7 9 9 2 9 11 13 2 13 4 3 9 13 13 4 2
25 13 7 12 9 2 11 2 0 11 2 9 2 12 9 13 4 2 11 9 2 2 9 10 1 2
14 7 2 9 10 9 13 4 13 4 2 7 9 3 2
16 0 0 0 9 13 9 13 4 12 9 9 2 13 9 1 2
25 9 0 13 3 13 13 4 3 11 11 11 12 9 2 7 10 11 9 10 12 12 13 4 9 2
10 12 13 9 2 3 0 13 9 1 2
13 10 0 3 2 13 13 9 10 9 13 4 9 2
19 11 9 9 13 4 2 7 14 4 3 13 2 7 14 2 7 2 9 2
24 11 11 9 0 9 7 9 11 9 9 11 11 13 13 4 9 2 7 9 13 9 13 4 2
16 2 11 11 3 13 13 4 9 0 13 9 7 9 0 13 2
18 9 10 13 4 9 11 11 1 13 4 12 9 10 14 4 9 13 2
18 11 1 11 11 0 13 11 1 3 2 7 11 13 4 9 13 4 2
15 12 7 13 4 13 2 12 9 13 4 0 9 10 1 2
14 9 13 9 9 9 1 2 9 12 9 12 13 4 2
14 9 0 9 0 11 11 13 4 2 7 9 13 4 2
11 11 11 14 13 9 12 9 13 9 0 2
10 15 13 4 2 14 4 15 7 13 2
22 9 9 7 9 9 7 9 0 13 4 10 1 2 7 10 9 9 0 13 13 4 2
18 13 4 2 3 2 9 0 10 13 4 14 9 2 7 9 9 9 2
24 9 10 1 2 9 13 4 9 15 9 13 9 13 4 2 9 9 14 4 0 1 13 7 2
20 12 9 11 0 13 4 11 1 2 7 9 12 13 4 11 7 12 13 4 2
20 12 9 9 9 13 4 12 11 9 2 11 7 9 9 0 3 13 14 4 2
15 11 11 2 12 9 9 9 0 3 2 11 13 4 12 2
17 9 1 13 9 10 2 9 0 2 13 4 7 9 13 13 4 2
16 3 9 14 4 3 3 13 2 7 9 10 13 9 13 9 2
16 12 9 2 3 7 3 13 4 11 2 7 13 4 9 13 2
12 11 13 4 12 9 0 2 7 11 12 9 2
13 9 0 3 0 3 13 4 13 4 10 2 9 2
8 14 13 11 9 9 13 4 2
13 11 2 9 10 13 9 0 1 13 4 12 9 2
19 11 9 8 3 13 4 3 2 7 11 7 11 11 7 14 4 3 13 2
22 7 2 3 13 7 9 13 4 9 9 9 0 9 13 4 2 9 10 13 9 0 2
21 9 13 13 13 4 9 11 9 2 11 9 12 13 4 2 7 11 7 13 13 2
9 3 9 13 4 11 11 13 9 2
9 9 1 13 9 9 0 0 13 2
11 12 15 13 4 9 2 9 12 13 4 2
9 9 9 13 4 12 11 4 13 2
8 3 7 3 9 10 13 4 2
21 3 2 7 2 11 7 11 11 11 11 9 0 9 11 9 13 11 2 9 13 2
11 7 2 9 2 11 13 4 3 9 10 2
10 0 7 9 10 9 3 13 4 2 2
9 9 1 13 7 9 9 13 2 2
25 9 11 11 9 13 4 9 10 13 4 11 9 2 11 11 9 9 0 7 3 9 9 9 13 2
41 11 0 13 11 3 0 13 9 2 3 13 3 11 9 14 13 3 0 7 2 7 2 11 9 0 0 9 2 0 13 0 13 11 2 2 9 0 9 13 2 2
14 9 3 2 11 9 10 9 0 0 13 4 9 0 2
20 10 1 10 12 13 7 0 13 2 15 0 13 15 0 14 13 0 13 3 2
9 9 1 13 9 13 0 12 9 2
15 9 10 9 0 13 4 7 9 1 13 4 9 9 13 2
20 11 12 7 11 3 14 4 0 9 13 11 9 7 11 11 11 13 9 0 2
12 12 9 10 9 13 13 4 13 4 9 0 2
17 2 0 9 9 10 13 4 2 7 3 1 14 4 3 13 13 2
12 11 11 9 13 9 0 12 9 12 13 11 2
14 3 2 12 9 9 9 0 9 13 11 9 9 13 2
24 11 12 9 11 11 2 7 2 9 0 13 7 9 13 4 11 9 2 12 9 13 4 7 2
15 13 9 2 9 12 9 13 4 11 2 7 12 9 9 2
10 9 1 13 3 2 15 9 13 4 2
12 9 10 11 11 11 11 13 9 12 9 13 2
7 3 13 4 11 11 9 2
8 9 1 13 7 9 13 4 2
23 9 2 9 9 2 11 11 12 9 9 12 13 4 9 7 9 2 0 2 9 9 13 2
12 12 9 13 4 11 11 9 2 12 9 9 2
9 12 9 0 13 2 11 11 0 2
19 0 2 12 12 9 9 9 0 13 4 2 7 3 0 13 4 9 1 2
15 10 10 3 13 2 7 10 9 0 13 7 9 1 13 2
5 2 11 11 13 2
22 11 11 7 2 11 11 9 0 9 13 4 2 7 13 12 9 11 9 13 4 9 2
10 12 9 3 2 11 11 11 13 4 2
27 9 9 9 7 9 9 14 4 9 9 3 13 2 9 7 9 13 4 2 12 9 9 7 12 9 9 2
18 9 9 13 4 2 9 13 2 13 13 4 11 11 2 11 11 9 2
12 9 2 9 9 9 13 13 2 14 9 0 2
13 11 1 2 9 10 10 14 13 9 13 9 9 2
16 11 11 3 9 0 13 4 11 1 2 7 0 13 4 9 2
19 9 10 7 9 9 1 10 10 3 13 2 0 9 9 3 13 13 4 2
20 11 9 9 0 12 9 13 4 11 13 11 9 0 9 11 11 13 9 13 2
28 12 9 1 2 11 13 4 10 9 9 1 13 9 13 7 9 10 3 9 11 9 3 13 9 13 4 11 2
12 11 13 12 9 1 13 4 11 12 9 9 2
19 9 7 9 13 9 13 11 11 3 2 11 9 7 9 11 13 9 1 2
11 9 2 13 4 15 7 12 9 10 1 2
17 11 11 9 11 11 11 9 13 4 2 7 14 13 10 13 9 2
8 12 9 13 9 11 9 0 2
30 0 13 4 12 2 9 14 13 0 2 7 9 12 13 4 13 9 9 13 4 9 1 2 7 9 3 13 13 4 2
11 15 13 9 3 10 9 1 2 9 13 2
17 11 11 9 1 2 12 9 9 2 12 9 9 2 13 4 11 2
14 11 13 4 3 11 11 2 11 11 11 9 9 9 2
21 12 9 9 9 13 4 2 11 2 11 2 2 7 9 0 9 11 9 13 4 2
23 11 11 11 9 9 9 13 4 3 11 11 13 9 1 2 7 9 3 13 4 13 4 2
15 11 11 9 0 13 4 11 9 7 11 12 9 13 4 2
12 12 9 2 9 10 13 4 7 10 0 9 2
22 9 9 10 2 9 1 2 9 13 4 13 11 2 7 13 9 9 13 4 9 10 2
3 9 13 2
16 9 0 12 9 9 13 4 9 9 9 9 1 9 9 13 2
11 11 9 9 13 4 2 0 3 2 0 2
15 0 9 10 2 11 9 0 13 2 7 9 0 9 0 2
9 9 10 9 9 13 4 9 9 2
23 13 4 9 1 2 9 9 11 11 9 12 12 7 12 9 9 13 4 0 2 13 4 2
10 9 0 13 2 9 0 13 9 1 2
17 11 9 9 10 9 13 13 4 3 2 7 15 14 4 3 13 2
16 11 10 3 1 9 0 3 13 4 10 9 13 4 9 1 2
9 9 12 9 13 4 12 0 1 2
11 11 7 11 11 13 4 14 4 9 13 2
6 13 11 0 1 13 2
14 9 1 13 9 0 3 13 13 4 3 11 9 11 2
27 13 4 2 15 9 0 13 2 7 0 13 2 9 0 9 12 13 2 7 2 9 10 11 9 9 13 2
24 13 4 9 11 11 11 3 13 9 2 3 12 9 13 4 11 7 11 11 11 2 12 2 2
10 9 13 2 11 9 13 4 13 9 2
23 3 9 0 1 13 4 12 9 13 9 2 7 3 2 0 9 14 2 13 13 4 11 2
23 11 9 11 12 9 13 4 12 9 1 2 11 11 11 13 4 9 0 7 11 11 9 2
28 11 9 13 9 0 9 2 3 12 9 13 4 7 10 9 9 1 13 4 2 3 9 10 9 0 13 4 2
12 11 9 12 9 0 13 13 4 2 13 13 2
9 11 11 9 7 9 13 4 13 2
15 11 3 13 12 9 9 2 11 1 2 7 14 4 13 2
7 9 1 9 0 13 4 2
9 9 9 3 12 7 3 9 13 2
12 11 9 9 0 13 4 9 11 1 13 9 2
11 11 11 13 9 9 0 13 4 13 4 2
12 9 10 11 11 13 4 11 11 2 12 2 2
17 9 0 9 0 13 4 2 7 11 9 9 1 10 9 13 4 2
14 3 2 15 9 13 13 4 2 11 12 2 11 12 2
20 2 9 13 3 7 12 9 13 4 2 9 10 11 9 0 13 4 9 13 2
28 10 2 13 9 9 13 4 9 9 0 9 7 9 2 11 2 9 11 7 11 2 11 11 9 9 13 4 2
20 11 11 7 2 12 13 4 11 9 9 13 9 2 11 9 13 9 13 4 2
26 11 11 9 9 2 9 13 13 4 7 0 9 2 11 9 2 13 2 7 13 9 13 4 13 13 2
12 11 11 9 9 0 13 4 13 4 3 9 2
17 9 2 9 2 9 2 9 2 9 7 9 9 9 1 13 9 2
10 11 11 9 12 11 9 13 4 9 2
10 9 12 9 1 13 4 7 12 9 2
31 11 11 11 9 10 2 11 9 9 2 0 9 3 13 13 4 2 13 13 4 11 11 9 0 9 7 11 11 11 9 2
17 11 11 2 7 2 14 4 13 2 7 9 10 13 3 13 4 2
15 2 0 1 9 9 13 2 7 9 13 9 10 9 13 2
15 3 0 7 2 9 10 1 9 13 0 13 13 4 11 2
22 11 9 2 13 12 9 11 11 1 13 12 7 9 14 4 2 9 0 2 12 13 2
6 9 11 11 13 4 2
8 9 1 2 9 0 13 4 2
18 0 9 9 11 0 9 9 13 14 4 10 9 9 13 13 4 13 2
8 9 0 9 9 13 4 9 2
12 9 10 13 13 9 1 10 9 13 13 4 2
10 9 0 9 13 4 11 7 11 1 2
10 9 12 12 1 13 4 3 0 9 2
11 2 9 1 0 9 12 13 4 9 2 2
15 11 9 1 11 7 11 13 4 9 12 9 13 13 4 2
16 11 9 2 11 2 9 9 13 4 11 9 13 4 12 9 2
9 3 9 12 9 3 13 4 13 2
17 9 12 9 13 9 11 11 2 12 2 11 2 2 7 9 12 2
20 9 9 2 2 0 8 3 13 2 9 0 3 3 13 10 13 10 9 2 2
25 11 11 2 11 2 11 11 2 11 7 10 1 9 13 4 12 9 7 10 11 9 13 13 4 2
7 11 9 13 13 10 1 2
20 9 0 13 4 11 2 7 10 0 9 9 13 0 13 2 9 0 13 4 2
9 9 1 9 10 7 10 13 4 2
6 10 13 4 11 11 2
10 11 13 4 2 3 1 2 12 9 2
10 3 2 9 9 13 9 9 13 4 2
13 9 1 11 2 9 2 13 4 11 9 13 9 2
11 12 9 9 9 13 4 11 9 1 9 2
11 11 9 11 9 9 13 4 9 9 13 2
6 9 9 1 13 4 2
12 9 9 9 0 2 7 2 11 11 13 4 2
14 12 9 2 9 13 4 11 7 9 1 13 4 9 2
15 11 3 13 2 9 9 9 10 13 11 1 9 13 4 2
12 11 11 0 9 13 4 2 12 9 13 4 2
11 9 9 7 2 11 11 13 4 2 9 2
23 9 9 0 13 4 11 1 13 11 9 9 7 11 1 9 13 9 7 14 4 13 3 2
12 11 9 13 4 9 2 9 13 13 13 13 2
9 9 9 13 13 4 2 10 13 2
6 11 11 13 4 9 2
11 12 10 2 9 12 3 13 4 9 1 2
26 9 9 11 11 3 13 4 2 11 9 13 4 9 9 9 2 2 11 11 9 3 13 9 13 2 2
19 9 7 9 10 9 9 0 13 11 9 11 12 13 4 9 2 12 9 2
20 9 10 9 0 13 13 9 9 9 13 4 9 13 12 9 9 1 13 4 2
22 9 1 2 11 11 7 11 9 7 13 4 10 9 2 7 10 12 9 9 13 13 2
15 2 15 3 13 9 7 15 9 1 13 4 9 0 13 2
11 2 12 9 11 3 13 9 0 13 2 2
17 11 11 9 2 0 9 0 13 4 2 7 9 9 9 13 3 2
8 11 11 11 13 2 12 2 2
11 2 2 3 7 3 9 1 9 13 4 2
6 13 13 4 9 1 2
22 9 0 9 3 13 4 2 7 11 11 11 9 1 10 13 12 9 0 13 13 4 2
25 15 9 10 0 1 9 13 4 7 7 9 12 12 9 13 7 9 3 13 7 9 3 0 13 2
16 3 2 14 13 9 0 9 13 2 9 1 13 14 4 7 2
15 7 9 10 13 4 9 9 13 2 11 10 9 13 4 2
29 11 9 2 7 2 9 9 13 9 13 3 7 0 9 3 13 4 0 9 9 0 2 9 9 13 11 9 1 2
26 10 1 2 9 0 9 13 4 9 12 7 9 10 3 13 4 9 9 11 9 2 12 11 1 9 2
19 9 10 13 11 2 7 13 4 9 11 13 4 12 0 13 9 13 9 2
11 11 2 3 13 4 9 9 9 9 9 2
13 9 10 9 13 4 2 9 13 7 9 13 13 2
19 9 12 9 9 10 13 7 10 9 10 9 4 13 2 13 13 9 13 2
8 10 9 1 13 4 10 9 2
23 11 11 9 12 9 9 13 4 3 9 13 9 9 2 9 0 9 10 10 13 13 4 2
26 11 11 2 11 11 7 11 11 13 13 7 13 13 11 11 2 11 11 7 11 11 9 13 11 1 2
16 3 13 10 1 2 7 10 10 9 9 13 14 4 9 13 2
16 10 10 2 7 2 9 0 13 4 11 9 9 3 13 3 2
15 12 9 9 2 11 11 11 13 4 11 9 9 13 9 2
26 2 9 0 10 9 9 9 9 9 10 13 9 13 4 2 7 2 3 7 3 11 9 13 4 2 2
12 11 11 13 4 2 3 2 9 0 9 0 2
9 11 11 0 13 9 9 10 9 2
10 9 11 9 2 13 9 0 13 4 2
10 9 0 13 4 11 11 11 9 0 2
14 11 9 13 13 4 13 7 9 10 13 4 0 9 2
16 9 9 0 11 7 11 1 9 12 9 13 4 2 9 9 2
20 9 0 9 2 11 2 9 9 13 0 4 2 7 11 11 12 9 13 13 2
22 13 2 2 9 9 2 7 2 9 8 9 1 2 9 13 9 10 13 9 13 4 2
16 2 14 13 15 0 9 1 2 7 3 0 13 9 0 13 2
9 11 7 11 11 11 13 4 3 2
26 12 9 11 13 2 11 13 7 12 9 13 3 9 11 13 7 2 3 2 9 13 11 11 2 13 2
10 7 13 4 11 11 11 9 9 0 2
15 10 1 10 2 9 2 13 4 13 4 11 9 9 9 2
19 3 2 10 10 15 1 13 13 2 7 0 9 13 9 0 0 13 4 2
20 11 11 11 2 9 10 1 11 9 13 2 9 0 9 9 0 0 13 4 2
22 13 13 9 14 13 11 9 2 9 7 9 2 13 2 7 7 9 13 9 9 13 2
12 11 11 13 4 2 13 2 13 11 13 9 2
12 12 9 1 13 4 2 3 9 10 13 13 2
11 2 9 9 0 13 7 9 13 9 13 2
16 9 13 7 10 13 4 9 9 9 13 4 9 1 9 0 2
18 11 2 9 13 4 9 9 1 2 9 1 9 13 9 13 13 4 2
9 7 2 3 3 9 0 13 9 2
8 9 11 9 2 13 2 13 2
41 7 12 9 0 1 11 9 9 0 13 4 2 9 12 9 12 9 13 4 2 3 12 9 0 13 4 2 9 11 13 4 7 11 2 9 3 0 2 9 13 2
18 2 11 9 0 12 13 2 7 2 3 2 7 9 9 13 4 13 2
17 3 9 13 9 11 9 13 9 11 12 13 13 4 10 9 9 2
19 9 13 9 3 9 13 4 2 7 11 1 14 4 10 15 9 10 13 2
46 11 7 11 13 2 0 9 1 2 3 13 9 13 14 13 0 2 7 13 9 13 2 7 2 9 10 2 0 13 9 13 2 7 9 12 9 1 10 9 13 4 13 9 13 4 2
14 9 9 1 2 3 3 13 7 3 9 0 13 4 2
28 12 9 3 13 9 13 4 9 0 14 4 9 13 9 2 2 9 9 10 13 2 13 4 9 0 9 13 2
12 11 9 1 13 9 13 9 13 13 4 2 2
8 11 9 1 9 0 13 11 2
10 11 9 12 9 13 4 11 12 7 2
19 9 9 1 2 11 11 9 7 9 12 9 9 9 13 4 9 13 4 2
25 3 9 3 13 14 4 9 9 13 4 11 13 10 9 2 7 3 9 10 9 13 4 9 10 2
