15696 17
6 9 7 9 1 9 5
13 9 2 9 7 9 13 1 9 1 10 0 9 2
9 7 1 9 2 11 8 8 11 2
28 9 13 9 2 11 11 11 11 8 11 2 2 15 13 0 9 1 0 9 2 1 9 2 9 7 0 9 2
12 3 13 2 11 8 11 2 8 8 8 2 2
23 15 13 0 9 13 1 0 9 2 9 13 1 0 9 2 7 0 9 1 9 7 9 2
12 9 13 2 11 8 2 8 8 8 8 2 2
20 9 1 0 9 2 0 9 1 9 2 0 9 2 0 9 2 9 7 9 2
33 7 9 2 2 11 8 8 11 2 8 8 8 8 2 13 1 11 7 9 1 0 0 9 2 9 7 9 2 7 9 1 9 2
4 13 1 9 5
18 0 0 2 9 12 2 13 9 15 1 9 1 14 13 9 1 11 2
28 1 9 7 0 9 13 15 1 9 2 0 2 9 2 9 2 9 7 9 1 9 2 9 7 0 0 9 2
17 15 4 13 0 1 9 11 2 9 11 2 9 11 7 9 11 2
12 10 0 9 13 1 0 9 3 10 0 9 2
12 15 13 9 1 9 1 11 7 9 1 9 2
13 3 1 9 13 9 11 7 9 9 2 11 11 2
15 1 13 9 9 2 11 11 11 2 1 9 11 1 9 2
16 3 1 0 9 13 9 2 11 11 2 7 9 11 1 11 2
17 15 13 3 9 16 9 1 10 12 9 4 13 1 0 0 9 2
13 7 3 13 3 9 1 11 7 11 9 15 3 2
4 9 7 9 5
16 1 10 9 9 13 11 9 11 11 11 1 9 11 1 11 2
39 3 9 11 1 11 1 11 0 9 2 11 11 2 3 9 11 1 11 1 10 0 9 11 7 3 3 1 9 10 0 9 2 11 1 10 9 11 11 2
16 0 9 13 3 1 10 0 9 2 3 3 1 10 0 9 2
22 9 4 13 1 10 12 9 0 9 11 11 15 13 9 9 2 11 11 2 1 9 2
20 9 13 0 9 1 11 11 9 2 9 11 2 15 3 13 14 13 0 9 2
11 7 1 9 13 9 9 2 11 7 11 2
6 9 2 0 7 9 5
18 1 9 4 9 1 10 12 9 2 9 9 7 10 0 0 0 13 2
32 0 9 13 9 11 7 11 11 11 10 9 1 9 2 16 9 13 11 9 1 9 7 10 0 9 13 9 11 1 10 9 2
28 9 11 11 13 3 10 11 1 9 11 11 1 9 2 7 9 11 11 11 13 0 3 0 1 9 1 11 2
31 9 11 11 13 9 11 1 11 1 10 9 2 16 9 11 4 13 10 2 9 11 2 2 10 12 9 0 9 11 11 2
29 1 10 0 9 4 9 11 7 11 13 1 9 2 16 11 11 7 11 11 11 1 9 9 13 1 10 12 0 2
5 11 4 13 9 5
20 11 13 9 1 10 0 0 9 1 11 2 16 11 13 15 1 10 0 9 2
6 11 11 4 13 9 2
21 10 0 9 1 11 13 9 9 0 1 10 9 15 4 13 9 1 10 0 9 2
23 1 1 13 15 0 16 11 4 13 9 1 9 7 9 2 1 3 11 11 7 11 11 2
16 11 13 9 3 1 10 9 2 16 11 13 0 9 1 9 2
18 16 11 13 9 1 9 2 13 10 9 1 16 9 13 15 1 9 2
10 10 9 13 0 1 10 9 1 9 2
19 1 9 4 9 13 1 11 11 11 2 16 11 11 11 13 9 1 9 2
9 11 11 4 3 13 9 1 11 2
9 11 13 3 9 1 9 7 9 2
17 11 13 9 1 12 9 2 9 2 9 7 9 2 9 7 9 2
12 1 10 12 0 13 11 9 3 1 10 9 2
12 11 4 13 9 7 9 2 16 11 13 9 2
7 11 4 3 13 10 9 2
21 11 11 4 13 9 1 9 2 9 7 9 2 16 15 13 0 9 1 10 9 2
10 11 11 13 0 9 1 9 7 9 2
7 0 9 1 11 1 9 5
2 0 5
3 0 9 2
12 11 13 1 10 0 9 1 10 12 0 9 2
12 3 1 9 13 9 0 9 2 1 1 9 2
9 0 13 0 9 1 10 0 9 2
4 13 9 1 2
23 1 9 9 13 9 11 11 11 1 1 9 11 11 11 9 2 9 1 9 1 10 10 2
19 3 13 15 10 12 9 9 1 12 9 15 0 9 4 13 1 11 9 2
14 1 9 4 9 13 9 7 9 1 10 0 9 11 2
34 1 16 12 1 12 9 1 11 4 13 10 10 9 2 7 1 16 11 4 4 13 10 9 1 9 1 11 2 13 9 3 0 0 2
12 7 11 4 1 9 3 13 9 1 11 9 2
16 1 10 9 4 15 3 3 13 15 15 13 10 9 1 9 2
17 2 15 1 9 13 0 2 15 0 13 1 10 9 2 13 15 2
19 11 13 1 9 14 13 9 1 9 2 7 3 13 15 3 10 9 9 2
32 15 7 10 9 4 13 1 9 0 16 9 0 9 13 14 13 9 1 9 2 13 10 9 1 9 7 13 9 1 12 9 2
31 3 16 11 2 9 11 11 7 9 11 11 15 13 13 10 9 0 9 2 7 3 10 0 2 13 9 1 9 0 0 2
15 1 0 9 13 0 9 1 0 9 1 10 9 11 13 2
19 10 9 13 15 15 3 0 15 13 2 1 14 13 10 0 9 1 9 2
18 11 13 16 10 0 9 3 4 13 0 1 14 13 1 9 1 11 2
29 2 15 13 0 3 1 14 13 16 10 0 9 4 15 13 9 1 11 1 2 0 7 0 2 13 15 1 9 2
12 7 11 4 13 1 16 9 1 11 3 13 2
38 1 9 1 9 4 15 13 16 10 12 9 13 9 1 11 1 0 9 2 1 9 1 10 9 1 9 15 11 2 11 7 9 13 1 12 9 3 2
13 11 13 0 0 1 0 9 1 9 7 1 9 2
28 1 9 13 15 16 10 0 4 13 1 14 13 9 1 9 2 3 16 9 3 13 0 1 10 9 15 13 2
31 7 11 7 11 13 3 10 9 16 10 9 1 9 1 10 4 13 15 0 14 13 9 1 10 9 1 11 7 3 11 2
14 7 11 9 13 1 1 14 13 9 0 0 1 11 2
25 1 10 9 7 12 4 15 0 13 16 9 13 1 1 14 13 1 10 0 9 1 10 12 9 2
14 15 13 3 3 0 16 11 3 4 13 9 1 9 2
27 1 9 13 15 3 0 10 9 2 1 14 13 16 15 13 2 10 3 0 2 14 13 1 10 0 9 2
12 2 15 4 13 3 0 9 13 2 13 15 2
15 16 11 13 14 13 15 1 14 13 9 2 13 11 3 2
12 2 15 13 10 9 0 14 13 1 15 3 2
7 11 13 9 1 11 10 5
29 1 9 9 1 11 7 9 1 11 2 11 11 7 11 1 11 12 9 1 9 9 2 13 15 3 0 10 9 2
25 1 9 13 11 9 1 14 13 1 16 9 13 10 9 1 9 1 11 11 11 1 10 0 9 2
49 11 11 11 4 13 14 13 15 0 16 9 4 13 2 7 16 15 13 16 9 2 7 3 15 10 2 4 13 10 0 9 7 16 15 13 16 10 12 9 4 13 16 9 0 3 13 10 9 2
33 7 1 9 13 3 11 1 9 9 16 10 12 0 9 13 0 1 14 13 9 0 9 11 11 10 0 9 1 9 1 11 9 2
11 10 9 4 0 13 10 9 1 10 9 2
14 1 15 13 10 9 15 0 1 9 13 11 0 9 2
25 7 9 4 0 13 1 16 9 0 9 11 11 4 13 1 9 1 9 1 10 0 9 15 13 2
44 9 1 11 9 13 10 0 9 1 9 7 0 9 2 9 1 16 10 0 9 13 9 1 14 13 3 15 4 13 0 0 7 0 0 9 7 10 0 0 9 1 11 9 2
28 7 9 1 9 4 13 1 16 10 12 9 3 3 4 13 16 15 13 0 1 11 9 1 14 13 1 9 2
22 15 4 3 13 10 0 0 9 1 11 1 14 13 0 10 0 9 2 3 0 9 2
33 3 16 0 1 11 7 11 13 1 1 14 13 0 1 14 13 15 2 13 15 10 9 16 11 13 10 0 9 1 11 0 9 2
47 10 12 9 4 3 13 1 11 7 11 1 10 9 15 4 13 0 1 9 1 9 2 7 15 4 4 13 1 14 13 1 11 1 9 3 3 1 10 9 2 7 3 1 9 1 9 2
15 7 15 13 9 15 0 1 10 10 9 13 10 0 9 2
22 10 9 1 11 0 13 3 16 15 4 13 10 9 1 16 11 4 13 1 11 9 2
9 1 15 13 15 0 9 1 11 2
22 10 12 9 13 3 16 10 9 4 13 0 1 0 9 16 15 7 11 13 0 9 2
19 10 9 13 0 1 11 1 16 15 3 13 14 13 0 1 10 12 9 2
36 11 2 11 7 11 4 3 13 0 1 16 9 1 11 4 13 15 0 0 9 1 9 1 10 12 9 15 4 13 1 14 13 1 1 9 2
19 11 4 13 15 0 10 9 15 13 1 14 4 13 9 1 10 0 9 2
33 3 16 15 1 9 13 1 16 10 9 13 16 10 9 13 0 2 4 15 0 4 13 3 0 9 1 14 13 0 1 10 9 2
8 9 11 13 9 1 0 9 5
19 11 0 9 2 9 11 11 2 13 9 1 14 13 10 9 7 3 13 2
22 11 13 15 1 10 0 9 11 3 1 11 2 1 1 11 2 16 9 13 10 9 2
12 15 4 13 9 9 1 14 13 2 7 13 2
11 11 1 9 7 9 2 1 10 0 9 5
3 0 9 5
3 0 9 5
22 11 11 4 13 1 9 2 7 13 0 2 10 0 9 2 15 13 10 15 15 13 2
10 0 10 15 15 13 16 15 13 0 2
8 11 4 13 1 14 13 9 2
33 1 11 11 2 15 4 13 1 9 1 0 12 9 3 2 4 11 13 10 0 0 9 15 4 13 0 9 1 9 7 10 9 2
21 11 4 13 1 9 2 7 13 0 2 10 0 9 2 15 13 10 15 15 13 2
10 0 10 15 15 13 16 15 13 0 2
7 16 15 3 4 13 9 2
6 16 15 3 13 9 2
5 16 15 13 9 2
5 16 15 13 0 2
5 16 15 13 9 2
5 16 15 13 9 2
13 0 16 15 13 2 4 11 11 13 10 0 9 2
17 4 15 13 11 10 9 2 13 15 1 0 9 1 12 9 9 2
21 15 13 0 1 10 9 2 7 15 13 0 0 9 1 0 9 11 13 15 1 2
18 11 5 9 2 15 11 3 4 13 1 1 11 9 2 13 12 9 2
2 9 2
17 0 4 13 16 15 3 13 3 15 13 7 16 15 4 13 15 2
2 9 2
28 0 0 1 0 9 13 3 9 15 4 13 15 10 0 7 0 9 16 15 3 13 9 2 7 0 7 0 2
2 0 2
14 11 2 0 1 11 2 13 15 0 9 1 0 9 2
12 15 4 13 1 9 7 4 3 13 1 9 2
13 1 9 4 15 13 1 14 13 0 9 1 9 2
8 10 0 9 2 15 4 13 2
12 10 9 1 9 1 10 0 9 13 1 9 2
20 11 4 13 10 10 9 2 11 2 1 9 1 11 2 15 3 13 1 15 2
16 9 9 2 15 13 1 11 11 11 2 13 0 1 1 9 2
14 3 11 9 2 11 2 13 11 5 9 0 1 9 2
41 11 13 1 12 9 2 7 0 9 13 0 9 9 7 9 2 9 2 0 1 9 2 11 5 11 7 9 1 14 13 9 1 9 0 2 1 9 7 1 9 2
27 11 9 2 1 9 11 2 13 9 1 3 12 9 9 9 1 2 7 13 0 9 1 12 9 1 15 2
26 10 0 9 13 1 9 1 11 2 7 3 1 11 2 11 2 11 7 11 1 11 13 0 9 9 2
12 1 9 13 9 11 9 1 12 9 0 9 2
30 9 9 2 11 2 13 1 9 1 0 9 2 1 1 9 2 7 3 0 2 0 2 9 1 9 1 9 1 9 2
8 10 0 9 13 9 1 11 2
19 11 13 3 9 1 10 0 11 1 10 9 7 1 11 1 11 1 11 2
11 9 13 3 1 14 4 13 10 0 9 2
7 9 13 0 1 11 9 2
49 7 9 13 9 1 10 9 9 1 10 9 1 9 15 13 9 1 15 2 1 10 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 0 2 9 2 9 7 9 2
35 10 1 11 0 9 13 3 1 9 1 9 7 9 1 9 1 0 9 2 3 3 1 9 1 11 11 1 1 10 0 9 9 9 1 2
13 10 0 0 9 13 1 9 1 11 0 1 9 2
23 15 4 3 0 13 1 9 2 0 1 16 11 4 13 10 0 9 15 13 0 1 9 2
7 13 1 9 7 1 11 5
5 13 9 10 9 5
2 9 5
21 11 2 3 1 9 7 9 13 9 1 9 9 1 9 1 9 11 11 7 11 2
6 1 12 13 15 1 2
2 9 2
23 9 13 2 9 13 7 9 13 15 9 9 3 1 9 9 2 11 7 11 9 11 11 2
6 7 15 1 10 9 2
6 9 13 9 7 9 2
25 9 13 9 1 9 9 1 11 9 13 1 2 7 0 9 13 1 7 13 9 1 11 1 11 2
8 11 11 7 11 11 13 9 2
22 11 11 2 15 13 11 9 1 12 2 13 3 10 9 1 10 0 9 9 1 11 2
21 7 10 9 13 15 15 1 9 2 15 15 4 13 15 1 0 15 13 1 11 2
34 11 11 1 11 2 9 1 12 2 13 3 10 0 9 11 13 1 9 2 2 7 9 13 3 9 1 9 1 9 2 1 0 9 2
12 15 13 3 3 9 7 9 2 13 15 1 2
22 0 9 1 11 11 11 2 7 11 9 1 11 2 11 11 2 13 1 9 1 11 2
39 2 11 13 12 0 9 15 13 1 9 7 13 9 2 7 15 13 9 15 4 13 0 1 10 1 10 9 2 13 2 11 11 2 2 13 1 10 11 2
41 9 2 11 2 11 1 11 2 11 11 2 9 2 11 11 7 11 11 11 13 16 9 9 4 13 3 0 0 1 9 1 9 7 9 1 10 0 9 1 9 2
42 15 13 3 16 9 4 13 0 1 10 9 1 0 9 2 15 4 3 13 10 9 1 11 1 14 13 0 1 1 14 13 9 15 4 13 1 9 7 11 1 9 2
18 9 1 9 13 15 3 2 16 9 13 15 1 9 1 1 11 11 2
34 9 11 11 2 1 10 9 1 11 13 1 9 7 9 2 7 9 11 11 13 10 9 1 16 0 9 4 13 3 1 9 7 9 2
7 1 11 11 13 9 1 2
13 7 9 0 13 9 1 1 11 0 0 0 9 2
22 0 2 0 9 4 13 3 1 2 15 0 1 9 1 10 0 9 1 10 0 11 2
19 11 11 13 3 1 10 9 11 7 9 1 11 9 11 11 7 10 9 2
19 15 13 0 2 13 2 13 7 4 3 3 13 9 1 7 13 1 3 2
4 7 9 13 2
11 1 11 11 0 9 4 15 13 1 9 2
6 13 9 0 1 9 5
4 11 1 9 5
28 0 9 1 0 9 9 1 10 9 7 1 10 9 13 11 7 11 9 16 11 9 4 13 1 11 9 9 2
4 10 3 0 2
38 0 2 7 0 3 2 13 11 9 11 11 9 1 10 0 0 15 4 13 15 1 9 9 16 15 9 1 11 7 10 9 13 9 9 1 11 9 2
13 2 1 9 4 15 4 13 10 9 1 11 2 2
31 0 7 0 13 15 3 2 1 9 11 2 9 7 9 11 11 2 1 9 1 9 2 1 9 2 9 2 11 7 11 2
44 7 1 0 0 9 7 9 1 10 0 9 9 2 15 1 0 7 0 2 1 9 7 9 2 9 7 9 1 0 9 13 10 9 1 12 9 1 10 9 1 10 0 9 2
34 1 9 0 9 1 10 0 9 1 0 9 1 10 0 9 16 9 13 1 2 13 11 11 15 1 3 14 13 10 0 9 1 11 2
14 10 0 9 13 1 10 0 9 16 9 3 13 9 2
16 7 3 10 9 16 9 1 10 0 9 13 3 0 7 0 2
28 11 2 15 3 1 11 4 13 1 11 9 1 9 1 9 2 4 3 13 9 0 7 0 1 10 0 9 2
9 15 13 15 3 1 9 2 3 2
18 2 15 13 1 9 0 1 10 9 1 10 0 7 10 0 1 9 2
49 15 4 1 9 13 16 15 3 13 1 10 9 15 10 0 7 0 4 13 2 3 16 15 1 3 0 9 1 15 13 14 13 9 1 9 2 0 9 2 9 2 9 7 9 2 2 13 15 2
15 1 9 1 15 1 0 13 9 7 13 9 1 1 9 2
27 2 15 4 13 1 10 0 0 9 7 13 16 1 14 13 10 12 9 2 13 15 10 9 15 13 2 2
18 2 10 9 13 1 16 15 13 9 1 12 9 2 2 13 15 0 2
19 2 10 9 1 2 0 9 2 13 1 16 12 9 13 15 1 10 10 2
16 9 13 1 16 12 12 9 3 4 13 10 0 9 1 9 2
30 15 15 13 1 10 0 9 1 14 13 12 9 9 2 13 3 3 0 1 10 9 1 0 9 2 2 13 11 11 2
23 9 9 2 11 11 2 13 10 9 1 12 2 10 12 1 11 2 10 0 1 11 9 2
30 15 13 1 10 16 2 1 10 0 0 9 2 14 13 9 7 13 9 2 13 11 3 3 15 10 9 4 13 1 2
20 1 0 0 9 13 9 0 1 9 7 13 1 10 9 1 10 12 9 2 2
34 3 13 15 0 1 10 12 9 9 15 2 13 3 0 0 1 10 0 9 1 0 9 2 1 2 10 0 9 1 11 0 9 2 2
22 1 9 9 13 15 3 0 16 2 15 4 13 0 1 11 11 1 14 13 11 2 2
32 2 3 12 1 11 12 0 9 4 13 1 11 1 0 9 7 0 9 2 3 11 11 2 9 10 9 2 2 13 11 0 2
19 11 13 3 10 12 9 1 11 15 4 13 9 2 3 1 16 15 13 2
42 2 10 0 11 13 7 14 13 10 9 15 11 7 10 9 11 11 3 4 13 2 7 14 13 15 1 14 13 0 1 9 1 10 3 0 0 11 2 2 13 11 2
5 13 10 0 9 5
5 2 11 11 2 5
7 10 0 9 13 1 9 2
27 9 9 2 13 1 9 1 11 11 2 11 7 11 2 13 9 15 1 11 11 1 14 13 10 0 9 2
32 2 8 8 8 8 8 2 13 11 11 1 11 7 13 1 1 11 11 2 15 4 13 1 1 9 1 0 9 1 12 9 2
15 1 15 13 12 9 1 12 0 9 1 11 11 11 11 2
10 1 12 9 4 11 11 4 13 1 2
10 1 12 1 15 4 11 13 1 9 2
25 9 4 11 2 10 9 11 11 7 9 0 13 1 11 11 1 0 9 7 1 10 0 9 9 2
20 10 0 2 11 11 2 11 7 11 2 13 1 9 3 1 0 9 1 11 2
42 2 15 13 1 10 0 9 2 7 3 0 15 13 9 1 9 15 4 13 1 9 2 13 15 9 1 10 0 9 2 13 9 11 16 15 13 9 1 9 9 12 2
19 1 9 11 11 13 15 10 0 9 16 15 4 13 15 1 10 0 9 2
26 15 13 11 11 2 11 11 2 1 0 9 1 2 8 11 2 7 13 12 9 1 0 14 13 9 2
5 2 4 13 9 2
3 13 3 2
12 2 8 8 8 8 8 2 13 11 1 9 2
13 2 15 13 3 1 14 13 9 2 7 13 9 2
28 10 9 1 9 13 9 2 9 2 9 7 9 2 13 9 11 11 2 15 13 9 9 3 1 9 11 11 2
24 16 9 13 0 2 3 1 9 15 13 11 11 1 9 2 13 9 11 11 10 0 9 1 2
22 2 15 13 0 0 1 14 13 3 1 9 2 16 15 4 13 11 13 1 0 9 2
38 11 4 4 13 2 7 15 4 13 9 2 7 11 13 10 0 9 16 15 13 1 9 2 7 15 13 3 0 2 13 15 1 10 9 1 9 11 2
22 11 13 9 1 11 11 1 16 15 13 10 9 2 1 9 2 7 3 1 10 9 2
15 10 0 9 4 1 0 1 12 9 13 1 11 1 9 2
10 11 13 15 1 14 13 9 1 9 2
12 7 16 9 13 10 0 9 2 13 15 3 2
12 2 15 13 3 10 0 9 1 9 7 9 2
8 15 13 10 9 7 13 15 2
10 15 4 13 10 0 9 2 13 11 2
33 9 11 11 13 16 9 2 9 7 9 2 1 0 9 7 9 1 11 11 2 13 0 1 3 2 1 10 9 7 9 1 9 2
23 2 15 4 13 1 14 13 9 0 0 2 13 9 2 13 1 1 10 2 11 9 2 2
23 2 16 15 13 9 1 9 4 15 13 10 0 9 1 14 13 1 1 0 9 1 9 2
55 7 1 10 10 9 2 10 0 9 14 13 9 7 9 1 2 13 15 9 7 9 1 10 10 9 1 1 10 0 9 2 13 11 9 11 11 1 9 9 7 13 1 9 7 9 15 4 13 1 1 14 13 11 11 2
5 9 11 13 9 5
18 1 9 1 11 9 1 9 13 15 0 1 2 11 11 2 1 11 2
19 9 11 7 9 1 9 13 9 1 9 2 7 13 0 9 1 9 3 2
19 9 13 9 11 7 9 1 9 16 10 9 13 1 9 2 11 11 2 2
15 7 3 13 15 0 0 9 1 11 9 7 1 1 11 2
20 9 9 13 9 2 11 2 2 7 3 13 15 9 1 9 1 11 11 11 2
9 3 13 11 11 0 12 9 9 2
26 7 9 1 9 11 11 13 15 3 3 2 3 13 10 0 9 1 1 0 9 2 1 10 0 9 2
11 13 0 9 3 2 7 13 0 1 11 2
7 11 11 13 15 1 11 5
19 11 11 11 13 14 13 15 1 14 13 3 2 7 3 13 9 3 0 2
8 1 11 13 15 0 9 9 2
13 11 0 9 2 11 11 11 2 13 15 9 3 2
21 10 0 9 1 9 1 11 4 3 13 14 13 1 9 3 1 9 1 9 9 2
17 1 12 9 9 13 15 9 7 9 12 1 11 9 1 11 11 2
13 2 15 13 10 9 15 15 13 0 0 0 1 2
11 15 13 16 15 4 13 14 13 1 9 2
29 15 13 0 0 16 15 13 14 13 9 10 1 9 1 9 15 13 1 11 7 11 2 13 9 11 11 1 11 2
29 11 11 13 9 1 9 1 9 12 9 9 2 1 9 4 15 13 10 9 16 10 12 0 1 9 9 4 13 2
13 2 15 13 0 14 13 3 15 13 15 1 9 2
14 15 13 3 10 9 15 13 0 0 1 2 13 11 2
10 11 11 4 3 13 2 9 2 9 2
19 15 13 9 12 1 12 9 9 2 12 2 7 12 1 9 2 12 2 2
16 11 11 13 3 9 9 2 7 13 9 12 1 12 9 0 2
9 11 11 13 9 1 12 9 9 2
10 10 9 2 12 9 9 2 13 9 2
17 2 15 13 0 10 0 9 1 10 1 9 2 13 11 1 11 2
5 9 13 11 11 5
4 2 13 0 5
4 2 0 0 5
6 2 4 3 13 0 5
10 9 13 9 2 7 9 13 1 9 2
18 7 11 11 13 3 1 1 11 11 2 7 15 13 3 0 9 1 2
13 11 11 7 11 11 13 0 0 3 1 11 11 2
9 3 13 15 9 1 10 11 11 2
6 7 15 13 3 3 2
33 1 14 4 13 1 10 0 9 1 9 1 1 10 9 1 9 2 7 13 1 9 1 10 9 2 13 11 15 1 14 13 9 2
9 2 15 13 3 0 9 1 9 2
13 15 13 3 14 13 2 7 4 3 3 13 15 2
13 15 13 0 16 15 13 1 9 1 10 0 13 2
15 7 15 13 3 1 14 3 13 15 2 13 11 1 11 2
11 15 4 1 13 10 9 1 10 10 9 2
28 3 3 13 15 0 1 9 2 7 16 15 13 14 13 9 7 13 1 9 2 13 0 1 14 13 1 9 2
18 7 15 13 0 1 16 0 9 13 1 9 1 9 9 1 0 9 2
14 9 13 3 0 16 9 11 11 13 14 13 1 9 2
10 2 9 13 3 3 15 14 13 1 2
7 7 15 13 0 7 3 2
10 3 13 15 1 11 16 15 4 13 2
17 1 14 4 4 13 1 9 15 2 13 15 12 9 1 10 9 2
14 15 13 3 14 13 9 2 7 13 9 2 13 11 2
6 7 3 13 15 3 2
6 10 0 9 13 3 2
12 7 9 13 1 9 2 7 13 1 9 0 2
8 3 13 15 15 1 14 13 2
9 2 15 13 3 0 9 1 9 2
9 15 13 3 0 15 0 7 0 2
13 15 13 9 1 0 12 9 2 13 11 1 11 2
29 16 15 13 3 12 9 10 9 13 15 14 3 13 0 1 14 13 9 0 1 11 11 2 15 13 1 12 9 2
6 7 1 1 1 9 2
9 9 1 11 13 11 10 0 9 2
19 1 9 2 12 9 1 10 0 9 1 10 9 2 13 15 0 1 9 2
7 15 4 3 4 13 0 2
8 2 6 2 15 13 15 3 2
17 15 4 4 13 1 0 1 9 1 15 3 2 15 13 15 3 2
20 7 15 13 0 0 0 14 13 1 1 14 13 1 10 9 3 2 13 11 2
13 1 16 0 0 9 4 13 2 13 15 1 9 2
17 11 13 0 11 11 0 2 7 4 3 13 1 9 1 10 9 2
10 2 11 13 3 16 15 4 13 15 2
20 15 13 15 3 1 9 2 7 3 13 15 0 7 15 13 1 9 1 9 2
5 15 13 0 0 2
10 15 4 3 13 0 3 2 13 11 2
15 9 1 12 13 1 10 0 9 1 10 0 9 1 9 2
13 1 9 4 15 13 0 1 9 1 0 0 9 2
17 2 7 15 15 13 3 13 3 9 0 2 13 15 1 11 9 2
18 3 0 9 11 11 2 11 11 7 11 11 13 0 9 1 11 11 2
3 13 9 5
4 9 9 12 5
6 9 13 0 0 9 2
4 13 15 3 2
8 13 1 10 9 3 1 9 2
11 9 1 9 13 14 13 16 9 13 0 2
14 3 13 15 16 0 9 3 13 1 9 1 10 9 2
20 7 15 15 4 13 9 2 13 16 9 1 12 9 1 10 9 13 0 0 2
20 1 7 1 13 3 9 16 9 3 13 10 9 15 15 13 0 4 13 1 2
17 7 15 15 4 13 9 2 13 16 1 9 13 0 9 0 0 2
23 0 0 9 1 10 0 7 0 9 2 0 9 2 16 0 9 2 8 2 2 13 0 2
22 10 9 1 9 13 16 2 15 2 4 13 0 7 10 9 4 13 16 15 4 13 2
15 7 15 13 3 0 1 9 2 3 16 9 4 13 3 2
7 3 4 15 13 0 3 2
14 10 0 1 10 9 13 0 1 16 0 9 13 0 2
15 7 3 13 15 3 16 10 0 0 13 1 0 9 3 2
12 9 13 3 1 9 2 13 15 1 7 1 2
11 7 13 3 9 1 0 9 1 9 3 2
13 15 4 13 9 1 10 0 9 1 14 13 9 2
17 15 13 0 9 15 13 1 16 0 13 3 0 0 9 1 0 2
19 10 0 13 3 0 1 16 7 13 15 0 2 7 3 13 15 15 3 2
6 7 9 13 0 0 2
15 0 13 15 0 16 15 4 13 3 0 1 10 10 9 2
26 1 0 7 0 9 3 2 7 1 9 7 9 13 15 1 10 0 9 1 14 4 13 1 10 9 2
9 10 0 9 4 15 13 1 15 2
17 1 9 1 14 13 1 9 2 4 15 13 1 7 13 15 10 2
10 15 13 3 3 9 13 3 0 9 2
5 9 13 0 9 2
18 7 1 9 1 14 13 1 9 2 4 15 13 1 7 13 15 10 2
5 2 9 13 0 5
2 9 5
9 10 9 4 13 1 10 0 9 2
12 9 13 1 9 1 9 1 11 9 11 9 2
13 11 13 9 1 10 0 9 1 11 2 13 11 2
39 2 1 0 9 13 15 9 1 0 9 2 7 15 13 0 1 16 0 0 9 0 13 2 7 16 0 9 13 2 13 9 11 11 11 1 11 1 11 2
20 9 1 11 2 15 3 13 11 2 13 1 9 10 0 9 1 11 9 11 2
21 7 9 1 9 3 0 9 2 11 11 11 2 4 13 1 15 12 9 1 9 2
39 2 15 4 13 9 1 10 9 3 2 7 16 15 3 4 13 13 15 10 0 9 1 10 9 1 9 7 11 1 1 11 2 13 9 11 11 1 11 2
13 9 4 13 1 9 1 16 10 9 4 13 9 2
15 1 11 13 9 3 3 2 7 9 7 9 4 4 13 2
12 3 13 9 15 3 0 16 9 0 4 13 2
12 2 10 9 1 9 4 13 10 0 1 0 2
16 15 4 13 10 0 9 9 7 0 9 1 9 2 13 11 2
5 13 9 1 11 5
2 9 2
4 13 14 13 2
23 9 13 9 2 7 9 11 11 11 13 0 11 9 15 3 4 13 1 11 1 12 9 2
11 2 10 9 13 0 1 11 7 11 11 2
35 3 7 0 2 7 1 14 13 15 3 2 11 13 10 0 9 14 13 2 7 3 4 15 0 13 9 1 9 9 2 13 11 11 11 2
26 15 13 16 15 1 9 7 13 7 4 13 15 1 1 9 9 2 7 1 9 4 15 3 13 15 2
14 9 13 1 9 1 9 11 7 9 11 9 1 11 2
8 15 4 13 1 11 1 9 2
23 11 13 9 0 9 2 7 11 13 10 0 0 9 1 10 9 15 13 10 9 1 9 2
27 2 10 0 9 13 0 9 1 14 13 3 15 13 1 11 2 7 15 13 15 9 0 4 13 15 1 2
23 15 4 3 13 3 1 9 1 9 2 13 11 2 15 13 9 1 14 13 0 7 0 2
20 16 15 13 0 14 13 1 11 2 4 1 10 9 9 11 7 9 11 13 2
19 1 9 13 0 10 12 9 0 9 1 11 2 7 15 13 9 1 11 2
24 3 13 15 1 10 1 9 1 11 11 2 11 2 7 13 11 11 11 9 2 9 11 11 2
15 11 7 11 13 1 10 1 9 2 15 13 11 0 9 2
8 1 10 9 13 9 9 0 2
15 2 9 1 10 9 4 13 3 15 13 15 1 0 9 2
22 0 13 3 10 9 0 2 3 4 15 13 15 1 10 0 10 9 2 13 9 11 2
12 9 11 13 0 1 7 9 7 11 11 11 2
24 2 15 13 0 9 2 7 15 4 13 15 13 0 14 13 9 1 15 2 13 11 1 11 2
18 9 11 7 9 11 13 3 9 1 14 13 10 9 1 9 1 11 2
11 9 13 10 0 9 16 9 13 1 9 2
12 1 9 1 9 13 11 11 11 1 11 9 2
6 15 13 9 1 11 2
15 3 13 15 11 9 1 9 2 11 2 2 1 12 0 2
11 11 13 1 9 1 12 9 9 1 11 2
14 11 13 10 9 15 13 0 1 9 1 9 1 9 2
17 2 3 1 13 15 3 16 15 13 10 0 9 2 13 9 11 2
12 7 15 7 11 13 0 1 16 11 13 0 2
35 7 9 11 13 16 15 1 0 9 13 1 10 10 9 1 1 12 2 12 9 3 16 15 10 13 7 13 9 1 9 1 11 7 11 2
6 2 13 15 14 13 2
13 2 15 13 15 2 7 15 4 3 13 1 15 2
6 15 4 3 13 1 2
21 8 8 8 13 15 15 15 13 2 7 15 13 0 9 1 15 2 13 9 11 2
4 11 4 13 5
6 3 0 0 2 7 2
4 13 1 9 5
4 9 1 9 2
5 15 13 1 11 2
4 10 0 9 2
10 9 1 9 3 15 13 0 1 9 2
8 15 4 15 0 13 1 11 2
7 14 13 15 0 13 0 2
10 10 0 9 13 10 9 1 9 10 2
28 15 13 3 9 1 0 9 15 3 13 1 1 11 2 7 9 1 9 1 9 16 15 1 9 13 15 1 2
14 9 7 0 9 10 4 13 1 1 15 13 3 9 2
19 1 3 4 15 0 13 0 14 13 9 1 9 15 3 3 4 13 15 2
17 11 13 1 9 1 0 9 1 0 10 10 1 12 9 0 9 2
5 15 13 12 9 2
10 1 9 4 9 13 12 9 1 9 2
19 3 4 9 13 1 14 4 13 10 0 9 0 1 2 9 7 9 2 2
31 15 4 3 13 9 1 11 9 1 11 7 1 11 1 11 7 13 10 9 2 1 9 0 9 2 1 14 13 1 9 2
18 1 0 9 2 7 0 3 1 9 2 4 3 9 13 0 1 9 2
17 15 13 10 0 9 16 9 3 0 13 9 1 14 13 9 10 2
23 16 10 0 15 13 1 1 9 13 10 9 1 9 0 1 10 9 2 4 15 13 9 2
17 1 11 9 4 3 15 15 4 13 14 4 13 1 9 13 13 2
14 1 9 13 10 0 2 0 9 10 9 9 13 9 2
10 9 2 3 2 4 13 9 1 9 2
29 2 15 13 16 10 0 9 13 1 7 13 0 9 15 3 4 4 13 16 15 13 9 1 14 13 1 0 9 2
27 15 13 3 3 1 9 2 7 15 13 9 15 13 0 1 9 1 10 10 2 13 9 11 11 1 11 2
11 15 13 1 16 11 9 13 10 0 9 2
28 2 15 13 3 9 1 16 9 4 13 0 1 9 2 7 3 16 15 13 10 0 9 1 9 2 13 15 2
18 3 9 15 1 9 13 0 1 9 4 13 7 13 1 11 0 9 2
23 9 15 3 13 9 10 0 1 9 4 13 1 15 1 10 10 9 1 10 9 13 8 2
15 15 13 1 10 10 0 9 2 7 11 13 3 10 9 2
6 15 13 0 1 9 2
18 14 13 15 13 1 11 9 13 1 15 14 13 1 14 13 3 0 2
8 15 13 15 1 9 1 9 2
7 0 9 4 3 4 13 2
19 15 4 13 16 9 4 13 1 9 3 0 0 9 1 9 13 1 9 2
32 7 1 16 9 4 13 3 0 2 4 15 13 10 0 9 1 16 9 1 9 13 0 2 7 16 9 4 13 0 7 0 2
23 9 4 1 9 9 13 9 1 10 9 15 4 13 2 3 15 15 13 15 14 13 0 2
13 9 7 9 11 11 1 11 4 3 13 1 9 2
17 2 15 13 3 10 9 1 15 1 16 9 15 13 4 13 0 2
30 16 15 13 1 9 13 0 10 9 1 16 15 13 9 1 9 2 7 15 13 15 16 15 13 10 9 1 10 9 2
24 1 3 4 15 3 13 1 9 2 7 3 1 10 0 0 9 13 15 3 1 14 4 13 2
29 16 0 9 4 13 7 13 2 4 15 3 13 10 0 9 1 15 15 13 1 11 1 10 0 9 2 13 15 2
7 11 2 13 2 1 11 5
6 2 15 4 13 9 5
3 10 9 5
6 2 13 1 1 9 5
8 11 13 3 9 1 14 13 2
18 9 13 11 1 0 2 7 13 16 15 13 15 16 15 13 10 9 2
2 11 2
24 10 0 9 11 10 9 1 11 4 13 1 10 0 9 2 16 9 7 9 3 13 0 9 2
17 10 9 13 15 10 0 9 11 11 11 15 13 0 9 1 9 2
22 1 9 9 4 10 9 13 0 1 1 10 9 15 13 10 0 9 2 13 9 11 2
34 9 13 11 2 7 13 15 1 14 4 13 9 9 1 11 2 10 9 1 11 2 7 10 9 7 9 1 11 2 1 9 1 11 2
5 2 15 13 0 2
6 15 13 1 15 15 2
13 15 4 13 9 1 9 9 2 13 9 1 9 2
16 9 13 3 1 9 1 9 2 7 13 15 0 9 1 9 2
19 11 13 9 1 14 13 9 10 2 7 9 13 1 14 13 15 1 9 2
4 13 9 3 2
11 7 11 7 11 13 9 11 1 10 9 2
10 9 2 9 9 2 13 0 1 11 2
21 1 10 9 3 13 10 11 0 9 0 9 1 14 13 1 9 1 11 7 11 2
12 1 9 13 9 9 1 9 7 9 1 9 2
6 1 9 13 9 9 2
14 2 9 13 1 1 9 2 13 9 1 9 10 9 2
14 15 4 13 1 1 16 9 13 1 1 9 2 3 2
5 9 1 11 9 5
3 13 9 2
5 13 3 1 9 2
9 0 9 4 13 1 1 0 9 2
4 11 13 9 2
44 9 11 13 1 10 9 11 10 3 16 11 11 2 3 2 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 7 11 11 2 0 1 2 4 13 14 13 0 9 2
18 9 1 11 11 2 11 11 11 2 1 0 2 13 0 2 9 2 2
6 1 9 13 15 11 2
20 1 10 9 13 15 3 9 1 9 1 10 1 10 0 9 1 10 0 9 2
10 9 1 11 11 13 14 13 0 9 2
20 7 1 1 9 13 11 11 2 15 4 13 10 11 10 1 9 1 12 9 2
12 2 15 13 0 16 11 4 13 9 1 9 2
16 15 13 1 10 9 2 13 9 1 11 11 2 11 11 11 2
32 11 4 13 1 1 10 0 9 1 9 9 2 3 1 10 12 9 15 4 13 1 1 14 13 1 1 11 2 9 1 9 2
34 2 11 13 0 0 9 2 7 9 13 10 10 9 14 13 1 2 0 9 2 7 15 4 3 13 0 9 3 3 2 13 11 11 2
37 9 11 11 2 11 11 11 2 9 2 2 11 11 2 9 2 2 11 11 11 2 9 2 7 11 11 2 9 2 4 13 1 11 1 10 9 2
11 2 9 15 4 13 1 9 13 0 9 2
11 3 4 15 13 15 9 1 10 0 9 2
25 15 13 11 1 14 13 2 7 15 13 3 9 1 9 2 7 10 0 9 13 14 13 10 9 2
14 7 15 4 3 13 1 9 1 12 11 2 13 11 2
25 12 9 1 12 7 12 9 4 1 0 4 13 1 1 14 13 10 0 9 3 1 9 1 9 2
23 10 0 0 1 15 13 11 11 2 12 2 1 11 2 3 0 1 9 3 1 11 11 2
62 2 15 13 15 0 7 1 11 7 9 2 13 11 2 15 3 1 11 11 2 12 2 11 2 11 11 2 12 2 11 2 11 11 2 12 2 11 2 11 11 2 12 2 11 7 11 11 2 12 2 11 13 10 0 9 1 9 1 9 11 10 2
34 1 15 15 4 13 11 9 2 13 15 1 11 11 9 12 1 9 2 3 1 12 10 1 10 9 2 7 3 12 9 1 10 9 2
34 2 15 13 0 1 16 15 13 3 1 9 2 7 15 13 1 10 9 2 3 16 15 3 13 0 9 13 10 10 9 2 13 11 2
8 1 9 13 15 0 0 9 2
15 3 13 9 3 0 1 16 9 13 1 1 9 7 9 2
26 14 13 1 1 9 1 11 11 1 9 2 13 3 9 1 9 10 0 9 1 10 0 0 0 9 2
5 2 10 0 9 5
22 9 11 11 7 11 11 4 3 13 10 0 9 2 13 9 11 11 1 11 1 11 2
15 2 11 11 13 0 9 2 7 15 13 9 4 13 15 2
9 11 13 0 1 9 2 13 11 2
29 2 15 13 0 1 10 9 14 13 0 9 2 1 11 2 11 7 11 1 9 7 11 2 11 7 11 1 9 2
11 11 13 3 10 10 0 9 2 13 9 2
7 1 11 13 11 11 9 2
14 7 15 13 3 9 1 11 2 9 11 0 4 13 2
26 2 15 13 0 14 13 9 1 9 1 9 3 1 9 2 7 15 13 3 0 0 2 13 11 0 2
19 2 15 13 3 10 9 16 15 13 1 0 1 0 9 2 13 11 11 2
11 11 13 10 9 13 1 10 0 9 11 2
23 0 9 13 1 9 11 2 15 13 10 0 9 2 7 15 3 4 13 1 10 0 11 2
7 11 13 0 7 13 9 2
7 11 13 3 2 9 2 2
17 15 4 3 13 0 0 14 13 9 9 1 0 9 2 13 11 2
18 2 11 13 10 0 0 9 2 7 15 13 3 9 9 2 13 15 2
17 2 9 15 13 13 9 15 13 0 2 7 15 13 0 0 9 2
20 9 13 9 4 4 13 1 9 11 7 11 1 9 2 1 9 1 3 11 2
20 2 15 4 3 13 14 13 0 0 2 7 15 4 13 0 0 2 13 9 2
7 2 0 14 13 9 3 5
12 11 11 11 13 15 1 14 4 13 9 3 2
16 0 4 13 11 7 11 1 9 1 16 9 0 9 4 13 2
16 11 11 13 10 0 9 0 9 1 16 9 11 11 4 13 2
21 2 15 13 0 0 14 13 9 7 10 9 2 0 2 13 11 11 11 1 11 2
21 10 0 9 7 9 1 11 11 4 13 14 13 1 9 11 11 0 9 9 9 2
29 9 11 11 11 2 11 2 4 13 9 1 10 9 15 4 13 1 1 9 9 16 11 13 1 9 9 1 11 2
9 15 13 10 9 1 10 0 9 2
26 2 15 13 11 7 11 11 1 10 0 9 2 7 9 7 9 1 10 0 9 2 13 11 1 11 2
19 9 13 15 13 10 0 9 14 13 1 10 9 16 10 0 9 4 13 2
24 9 11 11 13 10 9 1 9 7 9 1 9 1 9 1 9 11 11 7 11 11 0 9 2
7 2 10 0 7 0 9 2
25 15 13 9 7 15 13 9 7 9 15 3 4 13 9 2 13 11 9 7 9 11 11 1 11 2
18 11 4 13 1 9 7 9 9 2 11 11 2 1 9 1 9 9 2
25 1 9 1 1 9 13 15 16 15 13 11 11 7 11 11 4 13 2 10 0 7 0 9 2 2
8 9 9 4 13 1 11 11 2
33 11 13 0 9 16 15 4 13 9 16 15 2 1 9 1 14 13 9 2 4 13 10 9 1 9 11 2 16 15 13 15 13 2
28 2 15 13 1 0 9 15 4 13 16 10 9 2 9 11 11 7 10 9 2 11 11 2 4 13 10 9 2
8 9 4 13 11 11 11 2 2
16 9 11 11 11 13 10 0 9 1 11 7 11 7 0 9 2
19 2 15 13 10 9 10 9 10 9 4 13 7 10 0 9 1 10 9 2
20 15 4 13 9 3 0 7 13 11 9 1 11 11 2 13 9 11 1 11 2
5 2 0 1 9 5
16 9 11 13 0 0 1 9 11 11 2 11 2 13 1 9 2
10 1 9 13 15 7 9 11 1 9 2
15 2 15 13 0 14 13 3 11 9 13 1 9 1 9 2
26 1 1 9 13 3 10 9 0 2 7 3 4 9 3 13 15 1 10 0 10 9 2 13 9 11 2
13 9 13 1 11 2 7 9 13 1 11 1 9 2
19 1 9 13 9 1 11 2 15 13 9 1 7 11 7 0 10 0 9 2
12 9 13 1 10 0 9 15 13 11 0 9 2
8 1 10 9 13 9 9 0 2
10 9 13 11 9 9 10 1 10 9 2
23 9 11 7 9 11 4 3 13 11 9 11 11 2 15 13 1 1 11 11 11 1 12 2
12 2 9 13 0 9 2 7 15 13 3 11 2
13 15 13 0 14 13 10 9 2 13 11 1 11 2
9 2 13 9 16 9 1 11 13 5
21 9 1 9 11 2 11 11 2 13 15 13 9 1 11 1 9 1 9 1 11 2
8 9 1 11 13 2 13 11 2
14 2 0 1 9 13 10 9 1 14 13 15 1 15 2
26 13 15 10 0 9 1 10 0 9 1 10 0 9 1 9 1 2 7 15 15 13 15 13 10 9 2
9 0 1 9 1 9 13 1 9 2
19 15 13 0 14 4 9 13 1 10 9 2 13 11 1 10 9 1 11 2
7 11 13 9 1 9 11 2
27 1 9 1 3 15 13 15 1 10 0 9 2 13 15 16 15 4 13 0 1 14 13 9 1 10 9 2
18 9 11 4 13 1 11 1 11 1 9 2 7 13 1 0 9 9 2
15 9 11 11 13 0 1 11 9 1 16 9 13 1 11 2
19 2 15 13 10 0 15 4 13 2 7 15 13 0 9 1 10 0 9 2
23 15 13 10 9 1 0 1 16 9 4 13 15 0 2 7 15 13 15 0 2 13 11 2
22 10 0 9 1 9 13 11 11 1 11 1 11 2 15 0 9 4 13 9 1 11 2
18 2 11 13 16 15 4 13 9 1 12 9 16 9 13 15 3 0 2
16 15 13 10 1 9 0 9 2 7 10 9 16 15 13 9 2
11 15 13 0 9 16 9 13 2 13 11 2
11 11 4 3 13 9 1 14 13 0 9 2
6 0 9 1 11 11 5
14 9 11 11 4 13 10 0 9 1 0 9 1 9 2
9 9 13 1 9 2 13 10 9 2
20 9 11 11 13 9 16 11 13 1 9 1 10 12 7 10 0 9 0 9 2
13 10 12 9 0 0 9 4 3 13 9 7 9 2
33 2 15 13 15 14 4 13 16 9 11 9 13 0 7 16 15 13 10 9 15 4 13 15 2 13 15 1 10 0 9 1 11 2
10 9 4 13 1 11 1 9 11 11 2
26 10 9 1 11 13 16 15 13 1 10 9 11 0 1 16 9 13 1 7 16 15 13 1 0 9 2
21 2 15 13 15 1 9 2 15 13 15 4 13 15 1 3 1 9 2 13 15 2
21 15 4 0 13 14 13 1 1 0 0 9 7 13 9 1 10 0 9 11 11 2
9 11 11 4 13 1 11 1 12 2
4 9 1 9 5
20 11 11 7 0 13 0 1 10 9 2 9 13 0 7 15 13 0 9 0 2
4 10 9 13 2
13 9 1 11 1 14 13 1 0 9 1 10 9 2
14 1 10 9 1 9 2 13 11 11 3 10 0 9 2
9 1 1 12 9 9 4 15 13 2
23 15 13 10 1 9 1 12 15 3 13 0 2 7 0 2 3 11 7 10 0 10 9 2
13 11 4 13 10 0 9 1 12 13 1 0 9 2
11 10 0 9 1 0 9 2 1 9 9 2
16 0 0 9 1 9 1 0 0 9 1 3 9 1 1 12 2
11 10 9 1 0 9 15 13 1 0 9 2
20 9 1 9 1 9 13 1 9 1 14 13 9 1 1 9 2 0 9 3 2
8 15 13 0 9 2 11 11 2
2 11 2
14 11 11 13 0 1 9 1 11 1 9 9 1 11 2
10 7 15 13 3 2 0 2 1 9 2
17 2 15 4 13 15 0 1 1 9 2 7 13 3 3 0 0 2
22 15 13 1 11 1 14 13 15 2 7 15 13 15 3 16 15 3 13 9 1 9 2
21 15 4 13 3 0 9 1 1 9 2 13 15 13 10 9 2 13 9 1 11 2
8 2 0 3 1 14 13 0 5
17 9 9 13 16 15 3 13 2 0 2 1 9 1 11 1 3 2
16 2 15 13 15 13 0 3 1 14 13 0 1 9 1 9 2
17 15 4 13 11 11 2 7 4 0 13 1 15 9 3 1 11 2
13 9 16 15 3 13 14 13 0 9 2 13 11 2
14 16 11 3 13 1 11 11 2 13 11 3 3 0 2
6 2 0 9 1 9 5
15 2 15 13 3 3 0 16 15 3 13 1 1 11 11 2
14 15 13 16 10 9 13 0 0 1 0 2 13 11 2
11 15 4 13 15 0 1 0 1 9 3 2
11 2 1 15 0 4 15 13 10 0 9 2
22 15 7 10 9 13 1 9 1 10 0 9 1 10 10 9 2 7 15 4 15 13 2
16 11 13 10 0 9 2 15 13 0 0 2 13 11 1 11 2
2 11 2
13 11 11 4 3 3 13 15 15 13 10 0 9 2
25 11 13 10 0 9 1 11 1 11 11 9 2 7 13 16 15 3 13 10 0 1 0 9 3 2
12 2 6 2 15 13 3 10 0 2 13 11 2
7 2 3 13 15 10 9 2
12 2 15 13 15 3 2 13 9 1 10 9 2
14 9 13 15 0 3 0 9 2 16 9 13 1 9 2
13 3 13 9 1 1 10 0 9 1 9 1 11 2
2 11 2
8 11 11 2 11 12 2 12 2
19 1 0 9 13 11 11 1 9 2 13 0 1 9 7 13 0 10 9 2
6 2 10 9 13 10 2
13 2 9 13 0 2 10 0 9 1 10 0 9 2
18 0 13 15 1 1 9 15 13 1 10 9 7 13 3 13 1 15 2
9 3 4 15 13 1 9 1 9 2
7 15 13 10 9 14 13 2
19 3 13 15 10 0 9 7 15 13 15 12 2 12 2 13 9 1 11 2
17 15 13 9 1 0 9 2 13 0 1 2 7 13 16 9 13 2
9 2 15 13 15 3 0 1 15 2
11 14 13 0 1 10 10 0 9 13 0 2
12 16 15 13 1 9 13 15 0 9 1 9 2
21 1 9 7 9 13 15 16 15 4 13 2 7 13 15 1 16 10 9 4 13 2
15 15 13 3 2 3 13 15 3 14 13 9 2 13 9 2
4 2 10 9 5
8 10 9 4 15 3 13 0 2
18 10 9 13 9 1 11 2 7 13 16 11 13 7 13 1 10 9 2
8 10 9 4 13 15 1 9 2
15 2 15 15 13 10 9 4 13 16 9 13 10 0 9 2
7 15 13 0 7 0 0 2
22 9 13 15 1 2 1 16 11 2 11 2 13 1 9 1 15 2 13 9 11 11 2
3 2 0 2
23 7 15 13 0 0 1 14 13 3 11 4 13 1 9 1 3 0 9 1 9 1 15 2
12 1 11 13 15 10 9 15 3 13 10 9 2
21 3 13 11 3 0 16 15 4 13 1 2 7 1 9 13 9 0 9 1 9 2
11 15 13 3 0 9 2 13 0 11 11 2
3 11 0 5
10 9 11 11 4 3 13 9 11 11 2
28 2 15 13 10 9 1 9 2 7 0 13 15 15 1 9 13 1 9 3 0 2 3 16 15 13 15 0 2
22 1 0 9 13 15 0 0 2 13 1 10 9 9 7 4 3 13 10 9 7 12 2
9 15 13 11 3 13 1 1 9 2
24 3 10 9 1 11 1 11 11 2 0 12 2 12 2 7 9 1 11 13 11 9 1 9 2
4 0 1 9 5
12 2 15 13 15 0 1 1 9 1 0 9 2
24 3 13 15 1 10 9 1 16 11 13 12 2 12 2 7 15 13 3 9 13 0 3 0 2
11 15 13 15 10 0 9 2 13 11 11 2
16 11 11 13 1 16 15 3 4 13 1 9 1 10 0 9 2
20 2 15 13 3 3 0 1 16 15 13 10 3 0 9 15 13 1 0 9 2
7 15 13 3 3 0 0 2
13 15 13 9 15 13 15 4 13 15 1 0 9 2
3 11 11 2
11 11 13 12 2 12 1 11 11 1 9 2
6 13 9 1 9 3 2
10 10 9 4 13 2 9 0 1 9 5
5 9 0 1 9 5
4 11 13 0 5
4 9 1 9 5
7 9 11 13 10 9 9 2
9 10 0 9 13 9 12 1 9 2
7 9 4 0 13 1 9 2
10 9 4 13 1 11 9 12 9 9 2
19 2 15 13 15 3 1 9 7 9 2 2 13 15 1 10 9 1 11 2
39 11 4 3 13 9 1 0 9 2 7 1 15 11 13 2 13 15 10 9 1 10 9 15 13 16 15 13 14 13 1 1 11 1 11 3 0 1 0 2
10 9 7 9 13 11 1 9 9 9 2
9 9 11 4 13 10 9 0 9 2
13 3 4 15 13 1 3 9 13 7 9 0 9 2
11 9 11 13 1 0 9 1 9 11 9 2
30 9 13 1 9 1 11 1 0 9 2 7 3 4 9 13 9 1 14 13 0 9 2 7 13 9 9 2 1 9 2
18 11 13 15 1 16 9 11 11 4 13 1 7 1 16 11 13 0 2
19 7 9 13 15 0 16 9 11 3 0 13 1 3 1 14 13 9 3 2
19 9 4 0 13 9 9 0 0 2 7 15 4 13 1 9 1 9 11 2
12 0 9 13 11 2 11 7 11 2 1 11 2
10 3 0 9 1 11 7 11 13 0 2
19 7 9 4 3 3 13 10 0 10 9 1 10 0 9 2 0 0 9 2
14 1 10 0 9 13 15 3 9 15 3 13 12 9 2
24 10 0 9 4 3 13 1 9 0 2 9 11 11 2 12 2 2 9 1 9 1 10 9 2
12 3 1 9 12 9 13 9 1 9 1 11 2
18 9 13 15 0 9 1 0 9 1 11 7 10 0 9 2 1 11 2
14 10 9 4 15 4 13 9 1 11 0 9 9 12 2
16 13 1 10 9 1 11 7 11 1 9 1 9 1 10 9 2
6 11 13 1 1 11 5
3 9 12 5
3 0 9 5
12 9 11 4 13 1 1 11 1 9 9 9 2
6 3 13 9 1 9 2
8 9 13 11 1 9 9 9 2
28 0 9 1 13 9 7 9 1 9 1 9 9 2 16 15 1 9 4 4 13 10 9 1 9 9 7 9 2
13 10 0 0 13 16 9 11 4 13 1 10 9 2
30 7 9 4 13 3 1 16 1 10 9 2 9 7 11 0 9 4 13 1 9 9 7 9 2 1 10 9 1 11 2
10 9 4 13 9 12 1 9 1 9 2
15 1 1 13 9 9 11 11 2 15 13 12 9 0 9 2
10 11 13 3 9 11 1 10 0 9 2
10 9 11 4 3 13 1 9 1 9 2
13 16 9 13 11 1 9 1 9 2 13 15 1 2
30 15 4 4 13 1 16 9 11 4 13 9 2 3 15 9 9 11 11 13 16 9 11 11 4 13 1 9 1 9 2
32 7 16 10 0 9 4 13 0 0 1 10 12 0 2 4 9 13 15 1 16 9 4 13 1 0 9 1 9 2 1 11 2
41 16 9 7 9 13 1 11 10 9 1 9 2 3 15 13 16 11 11 4 13 0 9 1 9 2 13 0 16 9 1 9 7 10 0 9 13 3 0 1 3 2
5 9 4 0 13 2
5 11 13 1 9 5
14 11 11 13 0 0 1 14 4 13 10 9 9 9 2
11 15 13 9 1 11 15 13 15 1 9 2
28 10 9 1 9 13 9 7 13 16 9 15 10 9 13 10 1 11 3 0 7 0 9 2 4 13 1 9 2
25 15 13 3 10 9 1 2 11 2 15 10 9 13 10 0 9 1 0 9 1 11 7 11 11 2
23 10 0 9 4 15 13 1 9 9 0 1 9 1 9 7 9 1 9 1 10 0 9 2
26 9 0 9 9 13 1 16 15 4 13 9 1 9 1 10 0 9 11 11 1 3 12 9 1 9 2
12 2 15 4 13 9 7 9 1 9 1 9 2
18 11 11 13 3 1 9 1 14 13 10 9 15 13 1 9 1 9 2
4 2 12 9 5
3 0 9 5
4 0 1 11 5
3 12 9 5
20 11 11 13 3 16 15 13 1 14 4 13 11 16 15 13 15 1 9 12 2
11 2 15 13 9 1 9 3 1 10 9 2
22 16 15 4 13 2 3 0 9 13 2 13 15 0 1 16 11 3 4 4 13 9 2
27 3 13 15 9 9 0 1 9 7 3 10 10 9 0 1 9 2 13 11 1 10 9 1 11 9 9 2
15 2 3 13 15 1 7 13 7 13 10 9 2 13 11 2
7 9 4 13 10 0 9 2
21 2 1 11 2 11 2 11 7 11 4 15 13 10 0 15 13 1 10 0 9 2
9 15 4 13 10 9 15 13 0 2
17 1 14 13 15 13 15 10 9 15 3 13 1 9 2 13 11 2
37 11 13 0 0 1 9 16 15 13 0 1 16 15 13 1 9 1 11 11 11 2 0 15 9 11 11 11 13 9 1 10 9 16 11 13 9 2
12 1 9 4 11 4 13 1 11 9 11 11 2
17 2 15 13 10 0 9 1 11 1 16 15 4 13 14 13 3 2
20 15 13 2 15 13 3 15 1 15 2 7 10 9 1 10 9 2 13 11 2
19 9 13 16 9 13 10 0 9 1 16 11 4 13 14 13 15 15 13 2
9 2 1 9 4 15 13 12 9 2
17 15 13 1 14 13 1 9 1 9 1 16 15 0 13 0 0 2
13 11 4 13 1 9 1 15 15 13 0 0 1 2
36 2 15 13 3 9 1 14 13 1 10 9 2 7 10 1 15 15 4 13 13 16 15 13 9 1 11 7 15 13 9 1 11 3 1 12 2
12 9 15 4 13 1 11 13 15 3 0 1 2
14 15 4 13 0 9 1 9 15 4 13 2 13 11 2
4 10 9 9 5
4 0 0 9 2
5 13 1 10 9 2
5 1 0 13 0 2
3 0 9 2
5 0 9 1 11 2
3 0 9 2
4 9 1 9 2
5 9 4 13 9 2
9 1 0 9 13 3 10 9 1 2
10 1 0 9 13 0 1 9 9 9 2
13 9 13 1 1 14 13 10 0 9 9 7 9 2
12 1 10 9 13 9 1 9 1 15 7 15 2
14 1 9 2 10 9 2 7 9 15 4 15 13 1 2
14 7 15 16 9 13 15 1 15 7 13 10 0 9 2
14 9 15 15 10 13 7 13 2 4 13 10 10 9 2
13 15 4 10 13 9 15 4 13 16 9 13 9 2
11 11 13 15 9 1 0 9 7 0 9 2
10 9 1 9 4 13 10 9 1 9 2
6 10 10 13 0 9 2
19 9 1 9 2 9 7 9 13 1 15 0 9 2 3 1 10 0 9 2
10 1 10 9 13 10 0 9 1 0 2
19 15 4 13 1 9 7 13 9 2 7 1 9 0 9 2 1 10 9 2
20 9 13 10 9 9 2 7 15 4 3 3 13 3 15 4 13 15 1 15 2
7 1 10 9 2 15 13 2
17 10 0 0 7 0 9 13 3 3 3 0 15 15 3 4 13 2
26 15 13 15 3 1 9 3 2 3 16 9 1 9 13 1 0 9 0 1 10 9 15 13 1 9 2
15 1 13 9 1 9 7 9 1 9 2 7 15 13 0 2
14 1 11 13 15 1 12 9 9 7 1 12 12 9 2
22 9 4 13 1 1 10 0 0 9 1 0 2 0 15 0 0 9 13 1 1 9 2
19 12 9 1 10 9 1 9 7 12 9 1 9 1 9 13 1 9 9 2
14 15 4 4 13 1 10 0 7 0 9 1 10 9 2
27 9 7 11 9 13 9 7 9 1 10 1 9 1 9 1 9 2 7 9 10 4 13 9 1 10 9 2
5 7 3 13 9 2
8 13 1 9 3 9 1 9 2
10 10 0 0 9 13 3 0 14 13 2
18 9 1 9 1 11 1 11 13 15 9 1 15 2 11 0 9 2 2
28 15 13 3 0 9 1 0 9 2 16 0 0 9 13 0 9 7 13 9 7 9 1 9 1 1 9 9 2
30 10 9 9 1 11 1 11 2 12 2 13 15 10 9 1 9 1 15 15 13 10 9 0 1 9 2 10 0 9 2
32 1 10 9 0 13 9 10 0 9 2 7 15 13 0 9 1 10 0 9 3 15 4 13 9 2 3 1 14 13 10 9 2
26 1 11 4 15 13 10 0 9 1 12 9 5 9 2 9 2 1 9 2 15 15 13 11 0 9 2
14 10 0 9 13 1 12 9 5 9 7 3 0 0 2
24 1 0 9 4 3 10 9 2 13 2 2 16 10 0 9 13 0 1 9 9 13 1 9 2
25 10 0 9 11 11 13 3 0 7 13 12 9 5 9 2 7 10 9 2 1 14 13 9 13 2
10 7 15 13 16 9 13 10 0 9 2
9 4 3 15 3 0 13 1 9 2
15 7 4 15 13 9 1 16 9 1 10 0 13 13 15 2
23 16 9 13 15 13 9 15 13 9 2 3 4 15 3 3 4 13 9 0 0 0 9 2
14 9 9 1 10 9 13 16 9 13 1 9 7 9 2
9 9 13 16 9 1 9 13 9 2
14 3 13 9 1 16 15 4 13 0 1 14 13 9 2
13 15 1 9 7 9 1 9 16 9 13 1 9 2
6 3 13 15 3 3 2
11 9 13 15 0 2 0 7 13 9 10 2
18 15 13 3 14 13 1 10 9 1 16 9 13 0 7 13 1 9 2
4 3 2 0 2
16 11 9 7 11 13 16 15 3 13 10 9 1 9 7 9 2
30 10 9 13 15 0 14 13 15 1 1 10 0 2 16 9 13 0 9 1 9 1 9 1 14 13 9 7 13 9 2
46 0 9 4 3 13 16 15 4 13 9 2 13 11 7 9 2 13 9 1 1 9 2 3 13 1 9 2 13 1 0 9 2 0 9 13 0 9 2 2 7 13 9 1 0 9 2
19 10 9 13 0 16 9 7 9 13 0 2 16 9 1 0 9 13 0 2
17 16 9 13 9 2 4 9 13 0 0 9 1 14 13 0 9 2
17 3 0 13 9 2 3 13 15 9 2 7 1 10 9 13 9 2
32 11 9 2 11 2 2 11 9 2 11 2 7 10 0 11 2 11 2 13 9 14 13 2 7 15 4 13 1 0 0 9 2
13 3 4 9 7 9 13 1 11 7 9 9 11 2
19 9 13 16 10 9 13 0 0 1 0 10 9 16 15 13 0 9 0 2
9 15 13 15 3 0 14 13 9 2
21 13 15 3 9 2 7 3 13 15 16 1 9 13 2 16 9 13 9 14 13 2
27 10 0 0 9 1 0 9 1 9 1 9 4 13 16 9 0 9 4 13 1 1 0 9 1 10 9 2
9 15 4 13 1 9 1 12 9 2
14 13 15 13 14 13 3 0 0 9 1 10 0 9 2
2 11 2
8 15 4 13 1 9 7 9 5
2 9 5
2 9 5
10 9 11 13 12 0 9 1 0 9 2
16 2 10 1 15 4 13 1 9 7 9 2 13 9 11 11 2
20 11 13 1 11 16 9 3 13 1 16 11 10 4 13 10 0 7 0 9 2
16 2 15 13 3 9 4 13 10 0 9 15 10 9 3 13 2
12 4 11 10 13 15 2 13 15 9 7 9 2
13 3 3 10 0 9 13 3 2 13 11 1 11 2
18 15 4 9 9 13 1 1 9 1 11 1 10 9 1 9 1 15 2
17 9 13 3 10 3 0 9 2 7 15 1 11 9 4 13 1 2
24 11 13 1 11 9 2 16 12 0 0 9 4 13 1 1 9 1 0 9 1 9 1 11 2
23 2 7 15 13 16 10 10 12 9 15 13 10 9 1 9 12 2 12 2 4 4 13 2
17 15 4 13 0 9 1 0 9 2 1 3 9 13 15 0 9 2
30 1 10 9 4 15 4 4 13 3 0 9 2 7 3 13 15 9 1 0 9 1 10 9 1 12 9 2 13 9 2
29 11 13 16 15 10 7 9 4 13 10 9 1 9 1 0 9 15 3 4 4 13 1 9 1 0 9 1 9 2
7 2 9 13 0 7 0 2
12 15 4 0 13 0 1 0 9 2 13 9 2
16 11 9 13 3 9 9 12 1 14 13 10 0 9 1 9 2
20 15 13 0 16 9 1 11 9 4 4 13 1 1 0 9 1 9 7 9 2
4 0 1 9 5
3 0 9 2
2 9 2
4 13 1 9 2
2 0 2
2 9 2
9 9 13 9 10 9 9 1 9 2
14 15 13 0 9 7 0 9 15 13 1 14 13 0 2
11 15 13 1 10 0 9 1 10 9 9 2
11 9 13 0 9 1 16 9 13 1 15 2
7 9 13 15 15 13 1 2
22 9 13 1 10 9 1 16 9 1 9 9 4 13 2 7 16 15 13 15 1 9 2
9 7 15 13 3 10 0 0 9 2
28 1 9 4 15 13 9 1 9 1 11 11 1 11 11 2 0 10 1 2 9 0 9 1 9 7 9 2 2
9 15 4 3 13 3 0 15 13 2
25 11 13 10 0 9 14 4 13 1 2 11 11 2 1 10 0 9 2 11 8 11 2 1 12 2
28 9 13 15 16 15 1 14 13 9 7 9 1 10 9 4 13 9 1 9 1 14 13 0 9 1 0 9 2
19 15 13 16 11 4 13 0 0 7 0 1 10 9 1 10 3 0 9 2
27 15 0 0 9 1 0 9 1 9 2 9 11 11 1 11 1 11 2 13 0 0 0 16 15 13 15 2
14 15 13 1 11 1 9 2 1 10 9 1 11 9 2
13 2 15 13 0 1 16 10 10 9 9 13 9 2
13 15 4 13 10 9 1 9 1 10 10 0 9 2
18 13 15 3 15 2 13 15 10 0 9 15 0 4 13 0 9 2 2
14 12 9 13 10 0 9 2 13 1 14 13 10 0 2
23 15 13 1 9 1 11 9 2 15 13 15 13 0 1 9 9 1 12 9 9 1 9 2
9 7 15 13 3 9 1 12 9 2
32 3 9 4 13 1 1 3 14 13 1 10 9 1 14 13 9 9 2 1 3 14 13 1 10 9 2 4 15 13 15 1 2
24 10 10 0 9 13 10 9 9 1 9 2 15 13 10 9 9 9 13 15 1 10 0 9 2
10 7 10 9 2 15 0 4 13 15 2
22 10 9 1 10 9 14 13 9 1 2 13 14 13 16 15 14 13 1 9 13 0 2
2 9 2
16 16 15 13 1 10 9 1 12 9 2 4 3 15 13 0 2
8 3 2 15 13 3 10 9 2
18 7 15 13 3 16 14 13 1 10 9 1 12 9 2 15 13 0 2
18 1 9 7 0 9 1 11 13 15 0 0 9 1 0 7 0 9 2
15 13 1 9 1 0 9 2 7 13 14 13 10 0 9 2
4 13 1 9 5
4 13 1 9 5
3 0 9 5
3 11 9 5
2 11 2
5 2 11 1 11 2
10 13 15 13 16 15 13 2 13 9 2
10 11 11 13 11 0 9 2 7 9 2
7 15 13 11 13 9 9 2
6 2 9 2 11 2 5
12 11 0 9 13 10 0 9 1 9 1 11 2
24 9 13 9 1 10 0 12 9 1 2 9 2 2 7 0 13 15 16 11 9 13 0 9 2
9 7 11 4 3 13 1 10 9 2
18 2 15 4 13 1 0 9 2 10 9 1 15 2 13 11 1 11 5
29 10 0 9 13 10 0 9 1 3 10 0 9 1 10 0 9 3 13 14 13 3 10 9 15 13 0 1 9 2
16 2 15 4 13 3 2 7 9 1 13 0 9 2 13 15 2
9 2 4 11 13 9 1 11 11 2
18 2 15 4 3 13 15 1 14 13 1 1 10 12 0 1 9 3 2
12 13 15 13 16 15 13 2 13 11 7 13 2
20 15 13 11 13 0 9 9 2 7 13 16 11 13 3 14 13 15 1 9 2
20 2 15 13 2 9 2 2 7 15 13 3 15 1 11 7 15 4 13 0 2
12 15 13 0 0 2 0 7 13 10 0 9 2
19 15 4 13 15 1 10 10 12 15 13 2 7 10 12 15 0 13 1 2
29 10 9 4 13 0 2 7 15 13 1 11 1 14 13 1 10 12 2 13 9 15 13 9 9 1 10 0 9 2
8 15 13 9 1 9 11 11 2
10 9 13 11 3 4 13 16 15 13 2
20 2 15 13 9 1 10 0 9 2 7 15 13 0 0 1 14 13 1 11 2
16 7 15 4 15 3 13 14 13 1 10 0 9 2 13 9 2
14 15 13 11 0 9 4 13 9 1 0 2 0 9 2
20 2 15 4 13 10 9 2 7 3 4 15 13 1 9 1 9 15 4 13 2
16 3 13 15 10 0 9 2 7 15 4 15 13 2 13 15 2
12 9 13 0 1 16 11 13 9 1 11 9 2
21 2 11 7 11 13 1 9 1 2 7 3 4 11 7 15 13 0 1 14 13 2
13 1 15 4 10 0 9 1 11 13 14 13 9 2
25 15 4 13 0 0 1 10 9 2 7 15 4 3 13 0 3 1 14 13 15 1 2 13 11 2
8 0 12 13 1 9 1 11 5
4 9 1 11 5
5 13 11 1 9 5
4 0 14 13 5
7 1 10 0 13 12 9 2
23 10 0 9 1 9 1 11 1 11 4 3 13 1 1 1 12 2 13 9 1 11 9 2
24 15 13 3 3 9 1 0 1 10 0 0 9 2 16 0 9 13 15 0 14 13 1 9 2
32 10 9 15 13 9 11 1 11 9 11 2 13 3 1 9 1 9 2 7 13 3 10 0 0 9 1 1 11 0 1 9 2
17 10 9 1 9 1 9 1 9 4 13 9 1 9 1 10 9 2
3 13 3 2
7 0 9 1 9 1 11 5
30 9 4 12 9 1 9 13 1 11 11 11 11 2 10 0 0 9 1 11 16 10 12 0 9 13 11 2 13 11 2
22 11 9 11 11 13 9 9 16 9 1 9 7 9 13 1 9 3 1 11 1 11 2
16 3 9 7 9 4 4 13 1 11 2 9 13 10 0 9 2
25 11 0 9 13 15 0 2 7 9 12 9 9 0 9 13 9 3 1 1 11 11 11 1 11 2
35 15 13 3 0 16 15 4 13 15 1 11 2 7 13 9 1 10 0 11 1 9 2 7 10 0 11 9 2 13 11 11 2 11 2 2
29 9 2 15 1 9 13 10 9 0 9 12 1 11 2 13 9 1 0 2 2 4 13 1 9 16 15 13 11 2
29 1 11 11 2 13 9 2 4 15 13 9 1 0 1 10 0 9 1 16 9 4 13 1 14 13 9 3 9 2
17 2 15 13 9 1 9 1 9 7 9 2 7 10 9 13 9 2
28 10 2 9 2 13 0 7 0 3 0 1 16 15 4 13 13 14 13 2 13 9 1 11 11 2 11 11 2
26 1 0 1 9 1 11 13 10 0 1 11 1 9 1 1 9 10 16 9 0 13 16 11 13 0 5
17 2 10 9 13 0 7 15 4 13 0 9 1 9 2 1 11 2
27 10 9 13 16 15 13 0 14 13 10 3 0 9 1 1 9 10 9 2 13 9 11 11 1 11 11 2
6 13 9 1 10 9 5
7 9 13 1 9 1 9 5
31 10 0 9 4 13 9 2 9 7 9 1 10 9 1 9 15 13 3 0 1 15 15 13 1 1 9 2 13 9 11 2
16 0 1 12 9 13 1 16 9 13 9 1 11 1 11 9 2
17 0 0 9 13 1 0 9 1 14 13 15 10 0 9 1 9 2
22 2 4 3 10 0 9 13 10 10 9 2 13 9 16 15 13 1 9 1 0 9 2
31 2 4 15 3 13 2 3 1 9 7 9 2 9 9 1 14 13 9 1 10 0 9 2 1 9 1 0 9 1 11 2
23 9 11 13 11 2 15 1 10 0 9 1 11 13 16 9 1 9 13 9 1 10 0 2
28 2 4 3 9 1 9 2 1 9 2 1 9 7 1 7 1 1 9 13 9 1 10 0 9 2 13 15 2
14 1 10 9 1 11 13 9 1 10 9 1 12 9 2
26 15 4 3 13 1 9 1 11 11 2 10 0 9 15 9 11 4 4 13 15 1 12 9 1 12 2
4 4 4 13 5
3 0 9 2
6 0 9 2 0 9 2
4 9 7 9 2
3 1 0 2
13 9 7 9 13 3 7 0 2 7 3 0 3 2
18 15 13 16 9 1 9 4 13 1 0 9 0 16 9 13 1 9 2
2 9 2
7 2 0 1 11 2 2 2
17 9 4 4 13 2 2 13 9 11 11 1 9 1 9 1 11 2
18 9 0 9 4 0 13 1 1 9 1 9 1 9 2 9 7 9 2
15 9 1 9 2 9 7 10 9 13 1 1 9 1 9 2
16 1 3 4 9 0 13 13 1 9 7 9 1 15 1 9 2
22 15 13 3 10 9 16 15 3 13 0 9 1 9 1 16 15 2 4 4 13 2 2
18 15 13 1 10 0 16 9 1 0 9 13 0 0 1 9 7 9 2
15 3 13 15 0 16 9 13 0 0 1 9 9 7 9 2
11 3 0 4 9 13 0 1 0 0 9 2
14 15 13 3 14 13 1 10 9 15 13 1 0 9 2
32 16 15 13 1 0 9 13 15 0 14 13 16 9 3 0 13 15 1 9 1 0 9 1 1 9 1 16 10 0 4 13 2
11 15 13 10 0 9 1 9 1 0 9 2
11 15 13 0 16 10 9 13 0 1 9 2
34 9 4 13 3 2 1 9 1 9 1 1 9 11 2 0 9 1 0 9 2 1 10 0 11 11 2 7 0 9 1 9 7 9 2
31 0 9 4 13 15 3 16 9 3 0 4 13 0 1 9 1 9 2 7 4 13 1 9 1 9 1 14 13 0 9 2
17 0 7 0 9 13 16 9 3 4 13 1 9 7 9 15 13 2
18 3 13 15 14 13 1 0 9 1 9 1 10 0 9 1 0 9 2
34 1 10 10 9 13 7 9 7 9 1 0 9 1 9 1 10 9 1 9 1 0 0 9 2 7 3 3 1 10 9 15 4 13 2
29 1 14 4 13 10 9 1 9 2 4 3 9 3 13 15 15 13 0 1 2 3 13 0 9 1 9 7 9 2
15 1 14 13 0 13 15 0 16 0 9 13 0 1 9 2
13 15 4 13 1 0 1 16 0 9 13 0 9 2
38 1 10 1 9 0 0 9 1 11 11 11 8 11 11 2 11 2 2 13 9 10 9 1 3 0 15 13 9 1 9 2 3 10 9 1 15 10 2
31 15 13 3 16 0 0 9 13 9 1 0 0 9 2 7 16 9 7 10 15 3 13 0 9 1 0 9 4 4 13 2
20 9 13 16 0 9 3 13 0 9 1 15 15 3 13 9 1 9 7 9 2
22 13 15 3 13 10 9 1 0 9 1 0 9 1 0 0 9 7 1 9 7 9 2
10 15 4 13 1 14 13 10 1 9 2
30 1 0 9 1 9 7 9 13 15 9 9 1 14 13 0 7 0 7 1 14 13 1 9 1 10 1 9 0 9 2
28 9 1 0 9 4 3 13 16 9 13 15 1 14 13 0 1 10 9 7 9 15 13 1 9 1 0 9 2
4 15 13 0 2
19 15 13 0 14 13 0 9 7 9 1 9 1 14 13 9 1 0 9 2
19 0 13 15 0 13 9 1 9 1 14 13 16 15 13 7 13 0 0 2
22 1 9 1 15 13 15 3 0 14 13 0 1 16 9 7 9 3 4 13 10 9 2
8 15 4 13 9 1 0 9 2
22 1 9 7 9 4 9 13 10 0 9 3 16 15 4 13 0 9 14 13 1 9 2
19 15 4 1 9 13 0 9 1 14 13 9 9 1 14 13 9 7 9 2
20 0 9 13 0 2 7 10 9 15 13 14 13 9 2 4 13 1 14 13 2
11 15 4 3 13 10 0 13 10 0 9 2
5 11 13 1 9 5
3 2 6 2
4 13 9 9 5
3 9 13 5
5 11 12 2 12 2
10 7 9 13 3 10 0 9 1 9 2
4 13 1 9 2
24 11 11 11 13 16 9 4 13 1 1 15 2 3 16 15 13 1 10 0 9 1 12 9 2
16 10 0 12 9 13 11 10 9 7 0 0 9 1 11 11 2
6 3 13 15 0 9 2
5 1 9 2 3 2
4 11 11 11 2
21 3 13 15 1 9 15 13 1 11 11 9 2 1 10 9 16 15 3 13 9 2
21 2 15 13 3 1 9 2 7 13 15 1 16 15 3 0 13 1 2 13 11 2
14 9 11 11 13 0 0 2 7 13 0 9 1 11 2
14 9 13 1 9 2 7 3 13 11 1 9 1 11 2
4 1 9 3 2
3 0 9 2
17 11 10 4 3 13 0 1 14 13 3 0 1 1 11 0 9 2
8 2 15 13 15 16 11 13 2
5 2 3 13 15 2
6 6 2 2 13 9 2
25 2 3 13 15 0 2 7 13 1 1 14 13 1 2 13 11 2 15 13 11 13 1 9 1 2
29 9 13 3 1 9 1 11 9 2 7 13 3 16 11 9 13 0 1 10 9 15 4 13 1 0 9 9 12 2
15 15 13 3 15 7 10 1 0 7 0 15 13 10 0 2
12 1 10 9 13 9 9 0 9 1 0 9 2
22 2 11 2 3 13 15 2 13 9 1 0 9 10 9 11 11 11 13 9 1 1 2
12 15 4 13 15 9 7 9 1 11 9 13 2
27 1 12 9 13 11 11 10 9 1 9 2 7 13 1 16 9 13 10 9 2 1 10 9 0 1 9 2
16 15 13 9 1 1 10 0 9 1 11 2 3 11 13 9 2
22 15 13 3 9 1 1 10 9 15 4 13 0 9 1 15 7 10 9 10 0 9 2
10 11 13 16 9 4 13 1 1 15 2
5 2 3 13 15 2
19 15 4 13 1 15 10 9 15 4 13 3 2 15 13 3 0 2 15 2
15 15 13 3 10 9 1 16 15 4 13 0 1 10 0 2
13 2 15 4 3 13 9 10 0 9 2 13 11 2
6 2 7 9 13 3 2
13 15 15 13 14 13 0 1 1 9 2 13 9 2
18 11 4 13 0 1 9 1 0 9 2 7 1 0 9 13 15 0 2
8 15 4 3 13 9 1 9 2
13 2 10 9 1 14 13 15 1 2 13 11 11 2
18 9 13 16 15 2 3 2 13 9 2 7 3 15 15 4 13 9 2
11 15 13 9 1 9 0 9 2 11 11 2
13 2 15 4 3 13 10 9 1 9 2 13 11 2
8 11 11 5 11 11 5 11 5
3 0 9 5
3 2 9 5
5 2 9 1 11 5
27 10 0 9 1 9 1 11 1 9 12 13 1 9 16 15 13 15 11 11 1 0 9 1 11 10 9 2
6 9 13 1 0 9 2
24 15 13 2 0 11 2 1 10 9 13 7 1 9 2 11 2 7 9 2 11 2 1 9 2
11 2 11 11 13 1 10 10 9 1 15 2
23 15 13 1 9 2 7 4 3 13 1 10 0 9 2 7 15 4 15 13 2 13 11 2
25 15 13 3 9 1 11 1 11 11 1 11 2 7 10 9 4 15 13 1 10 0 9 1 11 2
5 15 13 0 9 2
22 15 13 3 11 11 2 15 3 4 13 1 9 1 10 0 9 3 16 15 13 0 2
22 7 11 9 13 10 0 9 2 7 3 4 11 13 1 9 1 9 11 2 11 11 2
14 1 10 9 3 13 15 1 9 1 11 9 1 11 2
46 2 3 0 15 13 2 3 0 0 13 15 1 16 11 13 10 0 9 15 13 2 7 16 15 4 13 0 14 13 11 10 0 0 9 2 13 11 11 1 11 3 1 9 1 9 2
20 2 15 13 11 1 10 9 1 14 13 1 15 15 13 15 2 13 15 1 2
18 15 13 1 10 9 11 9 11 11 1 10 9 15 0 4 13 15 2
18 1 9 4 15 13 9 2 7 13 3 1 1 0 9 2 1 11 2
17 1 9 11 11 13 15 10 0 9 15 4 13 1 10 0 9 2
6 2 15 13 0 9 2
27 15 13 9 7 11 4 13 10 0 9 15 4 13 0 1 0 9 2 13 11 11 2 0 9 1 11 2
9 9 1 11 11 4 13 0 3 2
14 11 4 1 11 11 4 13 15 14 13 9 1 11 2
13 7 15 4 3 13 1 11 2 16 15 13 9 2
9 11 11 13 1 9 9 1 11 2
29 15 13 1 0 9 11 0 0 9 2 0 1 10 0 9 2 7 4 13 1 11 1 0 9 11 11 1 12 2
9 15 4 13 0 9 1 12 9 2
12 2 15 13 0 1 11 2 7 9 1 11 2
16 1 9 13 15 10 9 15 13 2 13 15 1 11 1 9 2
9 1 9 13 15 3 0 1 9 2
4 9 1 11 5
5 2 11 11 2 2
13 15 13 15 15 13 10 0 9 1 11 11 9 2
13 10 9 13 15 0 1 0 9 1 10 0 9 2
26 1 9 13 11 11 9 1 12 10 0 9 16 10 0 9 4 13 15 1 0 9 7 9 1 9 2
11 15 13 10 9 1 9 11 9 1 9 2
10 15 13 0 2 9 1 11 2 3 2
13 15 13 16 9 4 13 1 9 1 9 10 9 2
10 3 4 9 13 10 9 10 10 9 2
8 15 13 14 13 10 0 9 2
15 7 3 4 15 1 9 7 9 13 1 10 9 1 11 2
26 11 13 10 0 9 16 9 13 1 9 7 9 0 9 2 1 9 2 1 9 2 1 9 1 9 2
14 3 3 2 0 1 11 2 4 3 9 13 10 9 2
6 7 11 9 13 9 2
8 13 9 13 15 15 15 13 2
4 1 10 9 2
20 3 4 3 0 9 13 0 3 1 14 13 9 10 9 1 10 0 0 9 2
6 10 0 11 1 9 2
25 3 15 10 0 9 3 13 3 10 9 1 9 2 4 10 0 9 13 1 10 0 9 1 11 2
9 10 0 11 4 0 13 1 9 2
15 9 11 11 11 4 3 13 16 10 0 9 13 3 0 2
5 15 13 10 9 2
8 7 9 4 13 10 9 1 2
7 0 9 4 3 13 9 2
18 15 13 0 16 9 1 11 3 13 16 15 4 13 1 11 11 9 2
21 3 15 15 13 3 0 0 2 4 15 3 4 13 3 14 13 9 0 3 3 2
25 15 13 3 10 9 13 1 16 10 0 0 0 9 1 11 13 0 1 11 11 1 9 1 9 2
6 15 4 13 1 9 2
19 0 4 10 0 2 0 9 1 9 1 0 9 13 1 0 9 7 9 2
4 9 13 0 2
16 7 15 13 3 1 10 9 3 10 0 9 1 11 3 13 2
19 7 9 1 11 4 13 15 0 1 9 0 1 10 0 0 9 0 9 2
4 9 1 11 2
7 7 11 13 0 10 10 2
9 11 13 0 10 0 9 1 11 2
15 15 4 3 13 0 1 9 14 13 15 1 9 1 11 2
7 15 4 15 3 13 1 2
21 15 13 3 0 1 9 14 13 1 1 10 9 3 15 15 13 1 11 11 9 2
5 7 3 3 0 2
6 9 13 10 0 9 2
18 7 15 13 3 3 0 14 13 9 1 16 11 9 4 13 1 11 2
19 11 11 2 0 9 1 11 1 11 9 2 13 3 1 9 0 1 11 2
13 10 0 9 13 3 16 11 13 10 9 1 9 2
35 9 1 0 9 1 9 2 9 2 7 9 1 9 7 10 0 0 9 2 4 13 11 9 1 10 0 9 3 16 9 10 13 0 0 2
19 4 0 9 1 9 1 9 13 1 9 1 9 2 4 11 3 4 13 2
8 10 9 13 0 9 1 15 2
18 7 15 13 3 1 14 4 13 0 9 1 9 1 9 3 1 9 2
14 15 4 13 1 16 10 0 9 4 13 1 10 9 2
9 15 13 3 14 13 15 1 3 2
8 3 4 15 13 9 7 9 2
5 11 1 0 9 5
3 12 9 2
3 13 9 2
44 11 4 13 10 9 1 9 7 9 2 15 4 13 9 1 14 13 10 9 10 9 1 0 9 1 9 13 1 9 2 7 10 9 15 4 13 1 10 0 0 9 1 9 2
11 0 9 1 9 4 13 0 1 10 9 2
19 0 13 4 10 1 10 0 9 1 0 9 7 0 9 13 9 1 9 2
19 15 13 12 9 15 4 13 16 9 4 13 0 0 9 1 9 7 9 2
10 3 4 9 13 1 0 9 7 9 2
17 3 4 15 13 1 16 10 0 0 9 1 9 13 3 1 9 2
29 15 4 13 1 7 0 9 1 9 2 3 1 9 7 9 2 7 1 9 1 0 9 7 9 15 13 0 9 2
15 3 13 15 0 16 9 1 9 1 9 13 1 0 9 2
15 0 9 13 3 10 0 9 1 9 1 9 13 1 12 2
22 0 13 15 16 10 0 0 9 2 11 2 2 0 1 11 1 1 11 2 13 1 2
23 10 9 13 3 10 9 1 9 15 0 9 13 2 7 9 13 3 10 0 0 0 9 2
22 9 13 3 7 14 13 9 1 9 1 9 2 7 13 16 15 13 0 0 1 9 2
28 13 1 9 0 9 1 9 2 4 11 11 2 11 2 11 2 13 1 10 9 15 13 12 9 1 9 9 2
25 9 1 9 13 14 13 0 9 1 0 9 2 7 9 4 0 13 13 1 0 9 1 0 9 2
24 1 9 1 11 9 1 9 7 9 13 15 0 1 10 9 11 9 13 1 9 1 0 9 2
42 1 9 1 16 15 13 9 1 9 1 0 0 9 7 0 9 2 13 9 9 16 15 13 0 14 13 1 3 9 1 0 9 4 13 1 0 9 1 10 0 9 2
35 1 9 1 15 2 13 11 16 15 1 9 1 10 9 13 1 10 9 1 1 12 9 9 1 9 1 9 1 0 9 1 11 7 11 2
6 9 4 13 1 11 2
25 9 1 0 7 0 0 9 13 0 2 7 15 4 13 9 1 14 13 9 2 0 9 7 9 2
13 9 4 13 0 1 10 0 9 7 13 1 11 2
26 9 1 9 4 13 10 0 9 1 14 13 9 1 11 7 9 2 16 10 9 4 13 10 0 9 2
10 11 13 3 0 0 1 9 1 9 2
19 1 14 13 1 0 1 10 9 1 9 1 0 9 4 15 13 3 0 2
6 2 11 13 10 9 5
3 0 11 5
2 9 5
7 11 2 11 12 2 12 2
7 9 1 11 11 1 9 2
2 0 2
23 2 11 13 0 7 0 10 9 15 15 3 4 13 1 2 13 11 11 1 9 1 11 2
2 11 2
32 2 11 13 0 7 0 10 9 15 15 3 4 13 1 2 13 10 0 7 0 9 11 11 1 11 1 14 4 13 1 9 2
6 2 13 15 15 6 2
21 3 13 15 11 13 10 9 2 13 9 11 11 16 15 4 13 15 9 4 13 2
9 9 11 11 13 14 13 9 9 2
19 2 10 9 2 13 9 15 13 2 1 2 7 13 15 15 13 1 9 2
7 13 12 9 1 11 11 2
5 2 15 13 15 2
13 15 4 13 0 9 1 15 1 9 2 13 11 2
2 9 2
5 13 11 9 3 5
7 2 0 0 14 13 11 5
8 2 13 11 12 1 12 9 5
11 15 13 15 0 3 1 11 11 9 9 2
24 1 16 11 4 13 1 1 12 2 12 1 11 11 2 13 11 0 0 9 15 4 13 9 2
16 0 11 11 2 15 4 13 1 9 1 0 9 2 4 13 2
7 2 15 13 0 1 15 2
15 15 4 13 0 2 13 9 15 13 3 1 9 12 9 2
11 16 11 3 13 9 13 11 11 1 9 2
16 2 15 13 0 0 16 15 3 13 16 15 13 10 0 9 2
24 3 13 15 3 0 16 11 13 2 13 11 2 15 3 13 0 0 1 9 15 13 11 9 2
13 2 15 13 10 9 2 7 0 7 0 3 0 2
30 9 13 3 1 9 1 1 9 2 13 11 2 15 13 16 15 13 1 11 11 15 13 0 1 9 1 9 1 9 2
12 11 13 9 1 9 16 15 13 15 1 9 2
18 11 13 11 13 9 15 13 1 9 2 7 13 3 0 1 9 10 2
13 2 9 13 1 9 1 15 2 7 15 13 0 2
18 15 13 16 15 3 4 13 10 9 1 9 1 10 9 2 13 9 2
8 0 0 0 1 9 1 9 5
12 0 4 13 0 7 0 0 1 9 1 9 2
10 11 13 9 1 9 9 13 3 0 2
2 11 2
5 13 15 9 9 5
16 3 10 0 9 4 11 13 12 9 15 13 9 2 13 11 2
11 1 0 9 13 15 12 9 1 0 9 2
15 2 0 9 13 3 0 9 2 13 9 11 11 1 11 2
15 7 9 13 1 0 2 7 3 0 0 0 7 0 9 2
23 13 15 3 12 9 0 1 16 9 13 0 2 4 15 13 15 1 2 13 10 0 9 2
17 2 1 0 9 4 15 13 0 16 15 13 0 9 2 13 11 2
24 15 13 16 15 3 4 13 0 9 1 9 1 0 0 9 2 1 9 1 9 7 0 9 2
5 4 11 13 15 5
3 13 9 2
2 9 2
2 9 2
20 1 0 9 1 11 2 4 3 9 11 7 11 11 13 14 13 1 10 9 2
10 2 15 4 13 10 0 9 1 11 2
21 15 13 15 13 10 0 9 1 14 13 1 15 15 4 13 0 1 9 1 11 2
14 3 4 15 3 13 9 1 3 11 11 13 10 9 2
8 15 13 3 15 13 1 9 2
24 16 15 13 0 9 1 9 2 4 15 1 0 9 13 1 9 2 13 9 11 11 1 11 2
25 2 7 16 3 11 11 4 13 1 9 2 13 3 3 15 15 15 4 13 1 10 9 1 15 2
37 2 3 3 2 7 3 13 9 14 13 16 15 13 9 1 15 2 15 4 13 15 1 16 15 13 0 1 9 7 9 1 9 2 9 7 9 2
19 7 15 13 10 9 1 14 13 10 9 1 11 11 1 1 11 1 9 2
13 1 11 4 9 1 11 7 11 13 10 0 9 2
37 10 1 10 0 13 16 9 13 11 1 9 2 7 4 13 11 1 14 13 10 9 1 12 9 9 15 11 4 13 1 11 1 0 9 1 9 2
21 11 13 3 1 1 10 0 9 1 14 13 9 1 9 0 16 15 13 9 1 2
20 15 13 0 3 1 1 14 13 9 1 14 13 0 0 7 0 9 1 9 2
23 16 9 1 9 13 14 13 3 0 2 4 15 13 15 1 7 15 4 13 10 0 0 2
12 2 15 13 1 9 15 13 0 0 1 11 2
17 15 4 13 1 9 2 7 13 16 0 9 3 13 1 9 12 2
10 10 9 4 13 0 0 2 13 11 2
9 2 15 13 1 9 0 1 9 2
13 0 9 15 13 9 1 9 13 3 3 0 9 2
14 1 0 9 13 15 0 14 13 15 1 1 9 9 2
23 16 0 9 7 9 3 13 9 1 14 13 15 1 9 2 4 15 13 0 2 13 15 2
19 15 13 16 15 13 0 9 15 13 10 9 1 9 16 9 13 3 0 2
7 2 9 4 13 1 9 2
60 7 16 11 13 1 1 10 9 1 11 1 1 9 0 9 1 9 7 0 0 9 16 15 13 0 14 13 15 1 9 2 7 15 3 13 10 9 2 13 15 10 9 15 1 0 9 4 13 0 0 9 1 14 13 1 9 2 13 11 2
6 0 9 0 1 9 5
4 0 1 9 2
4 3 3 0 2
3 13 9 2
10 0 9 13 0 9 7 9 1 9 2
12 12 9 1 10 0 9 1 11 13 1 9 2
20 15 13 0 1 9 1 9 1 11 16 9 1 10 0 9 15 13 13 0 2
4 9 2 11 5
27 11 11 2 0 9 1 11 11 2 7 9 11 11 13 9 13 0 0 1 9 16 15 4 13 0 9 2
13 16 15 13 1 9 13 15 9 15 13 0 1 2
17 2 9 13 10 9 15 13 0 1 1 9 2 16 15 13 1 2
13 3 13 9 1 9 9 7 9 2 13 11 11 2
17 10 0 9 4 13 15 1 15 15 4 13 16 15 13 1 9 2
12 12 9 1 9 15 13 1 11 2 13 9 2
23 11 11 1 11 13 16 3 16 0 9 3 13 3 0 9 1 9 2 13 15 3 0 2
14 0 1 10 0 9 13 9 1 9 7 11 10 9 2
24 2 15 13 0 9 13 1 9 1 9 1 9 2 13 11 2 7 13 9 7 9 7 9 2
10 2 0 4 13 1 9 10 0 9 2
15 4 3 10 9 13 0 0 1 9 7 9 13 1 9 2
27 2 0 9 13 1 0 0 9 1 0 2 7 15 4 3 13 10 9 1 10 0 9 3 2 13 11 2
14 15 13 1 16 16 15 13 9 2 4 9 13 0 2
23 9 1 9 15 13 1 12 2 13 12 9 0 1 9 1 9 15 4 13 0 1 12 2
14 16 9 1 11 4 13 9 1 9 2 13 9 0 2
18 2 0 9 7 11 9 1 9 2 13 9 2 13 0 9 11 11 2
3 13 9 5
3 0 9 5
4 9 1 9 5
3 11 9 5
2 9 5
5 12 9 1 9 5
7 11 2 11 12 2 12 2
16 11 11 13 15 13 10 9 14 13 1 9 1 11 11 9 2
32 2 15 13 10 9 15 13 11 2 7 15 3 13 1 11 1 9 2 13 11 1 16 15 4 4 10 9 13 12 2 12 2
15 15 13 0 1 9 2 7 3 13 15 9 13 1 9 2
13 2 15 13 3 3 14 13 9 1 10 10 9 2
12 13 15 1 9 1 12 9 13 9 0 0 2
17 7 9 2 15 13 10 0 9 1 9 2 13 0 14 13 3 2
8 9 13 3 1 2 13 11 2
19 15 13 10 0 9 1 9 1 9 2 7 13 9 1 10 7 11 9 2
10 3 11 13 10 9 15 4 13 1 2
10 2 15 13 10 9 15 13 0 0 2
12 3 13 15 10 0 9 2 0 9 7 15 2
5 7 9 13 15 2
16 15 13 10 9 16 15 13 9 1 10 10 9 2 13 15 2
26 15 13 0 1 16 9 3 13 9 1 0 9 13 9 2 7 13 15 15 1 15 13 10 0 9 2
14 2 15 13 15 1 9 2 2 7 15 13 15 0 2
17 9 13 16 15 4 13 2 7 15 13 15 0 1 16 15 13 2
13 2 12 9 1 1 9 2 15 13 15 1 15 2
16 2 15 13 9 15 13 9 2 7 15 13 10 9 1 9 2
10 15 13 0 2 0 7 0 1 11 2
16 11 13 10 0 9 2 7 13 1 10 0 7 0 0 9 2
24 7 10 0 0 9 13 0 1 9 16 9 13 15 2 7 4 1 10 9 13 1 1 11 2
30 10 0 9 13 1 0 9 10 9 2 16 11 13 0 0 1 2 7 10 1 10 12 9 13 14 13 0 1 9 2
14 16 9 13 12 9 4 9 3 13 10 12 9 10 2
38 11 11 13 1 11 12 9 16 15 13 15 0 7 4 13 1 10 9 3 0 1 12 9 1 1 9 10 9 9 2 7 9 11 11 13 3 0 2
41 11 12 9 16 0 9 1 0 9 4 13 13 11 11 1 16 15 4 13 3 1 0 9 1 12 9 9 12 9 1 9 2 7 9 13 0 7 13 1 9 2
11 3 2 1 9 1 0 9 2 13 9 2
15 11 13 10 1 0 9 1 11 11 11 1 1 11 9 2
22 11 11 13 1 9 7 13 9 0 2 7 1 3 0 0 0 2 1 10 0 9 2
12 9 11 11 13 9 2 1 0 9 1 9 2
10 11 11 13 9 1 9 1 0 9 2
17 9 13 1 9 1 0 9 1 9 1 9 12 2 12 1 11 2
17 1 9 13 11 0 2 7 13 1 0 9 1 9 10 0 9 2
7 7 15 13 3 12 9 2
7 11 11 1 9 1 0 2
6 9 13 1 12 9 2
20 11 11 13 1 9 2 7 13 3 14 13 9 1 9 1 9 1 11 9 2
24 7 9 13 0 1 11 11 11 1 0 9 2 15 0 4 13 9 1 9 1 11 1 9 2
17 11 13 1 10 0 1 9 2 7 13 3 1 14 13 0 9 2
16 7 10 0 9 13 3 0 7 0 1 10 0 7 0 9 2
15 12 9 1 9 13 3 0 9 14 13 1 10 0 9 2
19 11 11 11 13 9 1 9 1 11 9 7 13 15 1 14 13 15 3 2
35 15 13 0 2 1 1 15 0 2 1 7 11 11 2 11 11 7 11 11 2 16 15 0 13 9 1 1 9 1 9 1 10 0 9 2
6 0 9 1 11 11 2
41 11 9 1 9 9 11 11 4 3 13 1 1 9 2 7 13 3 0 1 16 15 13 1 12 9 1 10 9 1 11 0 12 9 1 9 2 7 9 13 1 2
30 11 13 1 1 9 0 9 1 9 1 9 2 7 13 0 9 1 9 9 1 3 12 9 1 1 7 9 7 9 2
16 11 13 3 1 9 9 7 13 12 9 1 1 11 1 9 2
4 9 13 9 5
11 9 1 11 13 0 9 0 1 0 9 2
10 9 13 3 0 0 1 9 1 11 2
11 3 13 11 11 1 9 1 11 11 11 2
7 2 9 2 11 11 2 5
11 9 4 4 13 1 0 0 9 10 9 2
33 9 11 11 13 1 10 16 9 1 11 7 1 11 11 9 1 11 13 2 10 9 2 7 2 3 13 3 14 13 9 1 2 2
9 9 4 13 1 1 9 1 11 2
9 9 13 0 14 13 1 0 11 2
2 9 2
7 13 7 13 11 11 9 5
19 9 11 1 11 4 13 1 10 9 1 9 2 7 15 13 0 14 13 2
3 11 11 2
12 2 9 13 15 15 13 1 15 1 2 6 2
26 15 4 3 13 1 9 16 9 13 0 1 9 1 11 13 1 1 9 11 2 16 15 13 10 9 2
9 1 11 13 15 1 9 0 0 2
16 7 1 9 13 9 0 1 9 1 15 9 1 9 7 9 2
3 11 11 2
14 2 9 15 13 13 0 1 1 10 10 9 1 11 2
21 1 10 9 13 15 1 9 1 11 7 3 13 9 0 2 15 13 10 0 9 2
14 1 11 13 15 0 9 2 7 13 15 0 1 9 2
2 9 2
5 2 0 1 11 5
5 11 13 10 9 5
3 11 11 2
13 2 3 13 9 9 2 15 13 3 1 9 1 2
13 7 1 9 1 11 13 15 0 0 1 9 3 2
7 9 13 2 1 10 9 2
8 7 9 13 15 3 0 0 2
3 11 11 2
27 2 9 1 11 13 0 1 15 2 7 1 9 1 15 4 15 13 0 0 9 16 15 0 4 4 13 2
8 15 4 13 0 3 1 9 2
5 11 1 0 9 5
7 15 13 2 13 7 13 2
10 9 13 15 12 9 1 9 1 11 2
16 7 15 13 15 7 3 2 13 15 10 1 9 1 0 9 2
5 10 9 13 0 2
19 2 15 4 3 13 16 15 13 10 9 2 10 9 1 11 11 11 2 2
4 15 13 0 2
5 15 13 0 9 2
25 15 13 2 10 12 2 3 12 9 1 11 9 3 12 7 10 9 1 10 9 2 11 11 11 2
53 15 4 13 0 1 9 11 13 10 0 9 1 12 9 3 2 15 4 13 3 1 9 2 3 0 15 4 13 1 9 9 2 7 4 13 1 9 1 15 1 11 11 3 9 7 9 1 15 13 1 14 13 2
12 2 6 2 15 13 15 3 2 2 13 15 2
10 2 15 13 3 3 9 1 15 2 2
54 7 3 13 15 15 1 9 16 15 13 0 14 13 16 15 3 13 0 9 1 10 9 2 1 0 16 15 3 13 9 2 3 16 15 13 0 0 1 11 9 7 10 0 9 10 9 7 9 13 1 10 0 9 2
11 1 9 13 15 10 0 9 1 12 9 2
30 0 9 1 9 1 10 12 9 15 13 1 10 9 16 11 9 13 10 9 9 7 4 13 9 1 11 11 1 9 2
4 9 4 13 2
34 3 13 15 2 3 1 9 2 7 13 1 1 9 1 10 9 2 1 10 10 0 9 2 15 4 13 12 9 0 3 1 11 9 2
33 15 13 3 9 1 9 11 2 10 9 15 0 1 10 9 4 13 10 0 9 2 15 13 9 1 0 9 7 15 13 15 9 2
23 15 13 1 9 9 11 13 1 10 0 7 0 9 1 1 9 2 0 9 12 1 9 2
19 15 13 0 16 15 13 0 3 3 2 7 16 15 13 1 9 1 9 2
45 9 1 0 9 13 0 9 2 3 0 9 11 1 9 2 7 15 13 0 11 10 9 15 4 13 1 16 9 9 7 9 13 10 9 0 1 10 0 9 3 1 1 10 9 2
21 11 13 1 9 1 10 9 15 3 4 13 1 9 1 11 2 15 13 1 9 2
39 9 4 3 0 13 1 10 0 0 9 15 11 2 10 0 0 2 7 3 9 1 11 2 4 13 9 1 0 9 7 9 2 0 10 9 1 10 9 2
36 15 13 1 10 9 2 3 0 1 9 4 13 14 13 0 1 9 1 9 1 15 2 16 11 11 11 4 13 1 10 1 9 0 0 9 2
12 16 10 0 1 12 9 13 15 2 13 15 2
8 2 7 15 13 3 9 2 2
7 0 9 2 13 1 9 2
20 7 10 9 1 9 2 15 13 14 4 13 9 2 13 15 4 13 3 0 2
5 0 13 15 10 2
25 7 15 4 3 13 0 9 1 9 2 15 4 13 15 13 1 0 9 2 1 9 7 1 9 2
17 0 2 0 7 0 1 10 3 0 2 4 15 13 1 10 9 2
11 11 11 11 4 13 10 12 9 1 9 2
12 15 13 0 1 9 7 9 2 9 7 9 2
4 15 13 0 2
30 15 4 13 15 11 7 11 2 13 9 1 9 1 9 1 9 2 0 3 10 0 2 7 3 1 0 9 1 11 2
20 3 4 15 13 1 11 1 10 9 2 7 3 1 14 13 1 1 9 9 2
26 3 1 4 15 13 1 10 9 2 13 9 1 0 9 2 13 12 9 9 2 7 13 9 1 9 2
12 9 13 1 0 0 9 3 3 1 10 9 2
28 15 4 13 14 13 0 9 2 4 13 1 9 10 9 1 9 5 9 2 7 13 0 9 1 10 0 9 2
45 9 16 15 4 13 1 7 13 2 4 15 13 10 0 9 2 3 16 10 0 9 3 13 0 2 7 16 9 13 12 9 2 16 9 13 0 0 9 2 7 16 15 13 9 2
35 1 10 9 9 11 10 13 1 12 2 7 15 11 7 11 3 13 15 1 1 1 12 2 2 2 13 15 3 10 0 9 15 13 1 2
24 9 9 13 11 13 1 15 10 2 15 4 13 9 0 9 3 0 9 13 10 0 9 0 2
15 16 15 13 0 1 2 4 9 13 0 9 3 9 1 2
39 11 7 10 10 15 4 13 15 1 15 2 4 3 13 1 1 11 11 7 11 2 11 9 2 15 13 15 14 4 13 1 9 7 9 1 9 1 11 2
28 15 13 1 10 9 3 11 11 1 9 2 7 4 1 9 13 1 11 2 10 0 2 3 3 9 0 9 2
22 7 9 9 7 9 4 13 1 11 2 9 11 13 1 9 2 7 15 10 9 13 2
13 3 13 0 9 10 9 1 9 1 9 1 9 2
9 10 9 4 13 9 1 0 9 2
8 0 7 0 9 13 0 9 2
15 7 3 9 9 7 9 4 13 9 1 0 7 0 9 2
7 10 0 9 13 0 1 2
30 16 15 1 9 13 1 10 0 9 2 13 1 9 1 9 1 7 1 11 2 13 15 9 15 13 10 9 14 13 2
5 3 0 0 3 5
12 0 0 13 14 13 9 2 3 1 11 9 2
10 10 9 1 11 4 15 3 13 0 2
8 13 15 15 14 13 9 1 2
15 15 13 12 9 1 1 9 1 9 1 11 2 13 15 2
31 0 4 15 13 10 9 1 12 9 9 1 9 2 12 9 15 3 3 13 2 7 15 13 1 10 9 1 9 0 9 2
3 1 13 2
3 0 0 2
8 15 13 10 3 3 0 9 2
31 15 15 1 10 9 13 9 2 1 10 9 1 11 9 2 4 13 12 9 1 9 2 7 10 9 7 9 13 0 0 2
18 15 12 15 13 3 0 2 13 1 7 1 1 1 9 0 1 9 2
16 3 10 9 13 15 1 3 15 4 13 14 13 10 0 9 2
21 10 9 9 13 1 9 2 7 15 13 3 0 2 13 15 0 16 9 13 0 2
16 3 13 9 14 13 10 9 1 9 2 1 10 0 9 9 2
8 7 4 15 13 16 15 13 2
43 1 9 9 13 15 3 10 0 9 15 13 16 9 4 13 1 10 9 2 7 3 1 10 0 0 9 1 9 1 16 9 13 10 0 9 15 0 0 9 13 15 1 2
10 9 2 9 2 9 2 9 2 9 2
17 0 13 9 7 13 0 9 1 9 0 9 2 7 0 7 0 2
12 3 13 10 0 2 9 11 2 11 2 11 2
36 9 13 3 9 1 0 7 0 9 2 9 9 4 0 3 13 1 3 1 9 2 7 10 9 1 9 13 9 9 7 9 1 10 0 9 2
23 1 9 13 9 1 0 9 3 0 1 1 9 2 10 0 9 4 13 10 9 1 9 2
32 3 16 11 11 1 11 13 10 0 9 9 1 9 11 2 13 15 1 9 10 0 9 7 9 13 0 1 10 9 7 9 2
6 7 3 13 11 11 2
34 10 0 0 9 13 1 1 0 11 2 9 2 15 3 13 10 0 9 1 9 2 7 15 13 1 1 9 7 13 3 1 10 9 2
30 3 13 0 0 9 16 2 8 8 2 13 2 10 0 9 2 2 7 10 13 0 11 1 9 2 11 2 7 13 2
39 11 13 10 0 9 1 10 9 1 10 9 3 12 2 15 13 9 1 9 7 13 1 1 11 9 10 0 9 1 9 7 9 2 1 9 7 10 9 2
20 7 15 13 10 9 16 11 3 13 1 9 1 14 13 9 1 0 0 9 2
16 3 13 15 1 0 9 10 0 9 1 9 1 9 7 9 2
28 10 9 1 9 9 13 0 7 0 2 7 1 9 1 10 9 4 15 13 0 0 9 1 9 1 0 9 2
31 7 9 2 15 1 15 10 3 13 0 1 9 7 9 2 13 0 7 0 1 9 2 1 9 1 10 9 7 0 9 2
27 1 10 0 9 4 3 9 13 9 1 0 9 2 7 15 13 9 1 9 2 16 15 3 4 13 9 2
10 9 13 3 1 3 0 7 0 9 2
6 9 13 15 1 1 2
13 3 13 9 1 9 2 7 3 0 1 0 9 2
43 9 10 0 13 1 0 9 2 16 15 4 13 10 9 9 16 15 13 0 2 7 4 13 9 1 9 2 13 16 15 3 13 0 1 9 1 9 2 9 7 10 9 2
13 3 3 1 9 4 15 13 0 1 10 9 9 2
19 9 13 3 13 10 0 0 9 2 7 9 4 15 3 3 13 7 13 2
22 3 13 9 1 14 13 10 0 9 2 1 0 0 0 7 0 9 2 0 3 0 2
29 14 13 9 2 0 9 2 1 0 9 13 14 13 1 9 1 9 2 13 15 1 2 13 10 0 10 0 9 2
16 15 13 9 1 9 2 7 3 1 0 9 2 9 2 9 2
47 9 4 13 3 0 15 13 2 7 3 0 15 13 16 15 4 13 2 7 9 1 14 13 2 9 1 14 13 0 9 7 9 1 9 1 10 9 15 13 9 2 13 1 10 9 9 2
18 3 1 11 13 15 3 3 16 9 4 13 0 9 1 9 7 9 2
25 1 9 1 10 9 13 10 0 9 0 9 2 3 0 13 15 3 2 7 13 0 9 1 9 2
21 15 13 1 10 0 13 3 0 15 13 9 1 10 2 0 2 9 9 1 9 2
15 7 15 13 3 15 13 16 15 3 4 13 2 11 2 2
38 15 13 10 0 0 9 2 9 13 15 3 2 11 11 11 2 15 4 13 1 11 11 1 9 2 7 15 3 13 14 13 10 9 7 9 1 9 2
31 10 9 13 15 1 15 1 10 0 9 2 10 0 9 1 9 7 9 2 0 10 9 2 4 13 1 1 10 0 9 2
9 10 9 4 13 1 9 1 9 2
3 15 13 2
12 2 15 13 3 10 0 9 15 13 1 2 2
5 11 11 11 13 2
15 2 6 6 2 15 4 13 10 0 9 1 1 12 9 2
18 13 15 13 15 4 13 14 13 10 0 9 1 0 12 9 1 2 2
6 10 0 9 13 0 5
3 11 9 2
4 9 1 9 2
2 9 2
10 11 11 13 3 1 9 1 10 9 2
10 16 15 3 13 9 14 13 10 9 2
23 11 9 1 14 13 10 9 7 10 9 1 0 9 4 3 13 9 1 0 9 1 9 2
20 0 15 10 9 4 13 1 9 2 13 11 0 9 1 9 10 9 1 11 2
13 11 13 0 1 16 9 4 13 15 1 9 1 2
18 3 13 15 3 12 9 1 10 0 9 16 15 13 11 11 0 9 2
11 15 13 0 3 1 9 1 10 0 13 2
13 11 13 1 10 9 0 9 15 13 0 1 9 2
38 1 9 11 11 0 9 1 11 7 11 9 2 1 9 2 7 10 0 0 9 1 15 15 4 13 1 14 13 9 9 2 13 9 1 0 9 0 2
9 11 4 3 13 0 9 14 13 2
34 1 1 10 0 10 9 3 4 15 13 1 0 9 16 15 4 13 1 10 1 9 0 9 2 9 9 1 9 7 9 1 0 9 2
10 0 9 13 0 7 0 9 13 9 2
19 9 1 11 4 1 0 13 1 10 0 9 16 15 4 13 12 9 1 2
32 15 4 13 0 16 15 3 4 13 9 1 14 13 10 9 16 9 7 9 3 4 13 1 0 7 0 9 1 10 0 9 2
5 11 13 15 13 2
10 1 9 13 15 1 10 9 0 9 2
8 1 9 1 14 3 13 0 2
17 1 15 15 4 13 14 13 9 1 15 15 13 1 10 0 9 2
4 9 13 0 2
5 15 13 0 0 2
39 15 13 10 9 1 10 9 15 13 1 10 0 9 1 14 13 0 7 0 0 2 7 10 9 15 13 14 13 15 1 1 10 9 1 13 10 10 9 2
20 9 4 3 3 13 1 10 0 9 1 10 0 9 15 13 1 10 0 9 2
9 13 1 9 15 13 10 10 9 2
25 16 13 7 13 9 2 15 13 1 10 0 9 2 7 13 3 9 7 9 1 11 4 13 9 2
23 15 15 13 9 1 9 1 10 9 1 1 0 0 9 14 13 10 9 2 10 10 9 2
40 2 7 10 9 15 15 1 10 9 4 13 1 1 3 0 9 15 13 1 14 13 10 9 1 9 2 13 3 1 15 1 0 1 10 10 2 2 13 11 2
30 1 11 9 13 15 16 9 13 1 11 2 15 1 9 1 10 9 0 9 4 13 0 9 1 9 9 7 9 2 2
19 15 15 13 2 13 11 1 9 1 10 9 1 9 7 10 3 0 9 2
6 10 0 2 9 2 5
3 9 9 2
3 0 9 2
3 9 9 2
3 11 11 2
4 9 13 15 2
4 9 1 9 2
26 16 9 11 11 13 16 15 3 13 9 2 13 15 16 15 3 13 9 1 10 9 1 10 0 9 2
3 0 0 2
33 1 9 11 11 13 11 9 1 10 0 9 15 13 9 1 0 9 2 7 15 0 0 13 1 9 1 9 1 14 13 15 0 2
19 3 13 11 10 9 1 9 2 7 0 3 15 4 13 2 13 15 1 2
8 11 13 11 1 12 1 9 2
46 11 11 13 1 11 7 11 9 16 16 11 13 2 13 11 0 1 12 0 0 9 2 10 12 1 11 11 16 15 13 9 1 0 9 5 9 2 10 0 1 16 9 4 13 9 2
14 10 9 13 0 2 0 9 2 16 11 9 13 11 2
14 0 1 9 7 9 9 13 9 1 9 9 10 9 2
23 9 3 1 11 11 11 13 0 9 15 13 9 3 3 4 13 2 7 3 13 0 9 2
20 3 13 10 0 9 1 9 11 11 15 13 10 0 9 1 10 0 9 9 2
13 9 13 16 9 15 13 1 0 2 3 13 3 2
5 9 13 10 9 2
8 15 13 1 9 0 9 1 2
31 9 7 9 13 1 0 9 0 0 0 16 9 0 13 2 0 1 9 2 13 0 11 11 2 3 13 1 11 0 0 2
17 1 11 8 2 11 8 8 8 8 13 15 3 0 9 0 13 2
40 15 13 16 9 1 0 9 13 10 9 1 0 9 7 13 1 9 1 10 9 16 9 2 3 1 9 2 13 1 10 0 9 1 0 9 1 14 13 9 2
4 9 13 0 2
12 1 9 1 9 13 15 9 15 13 0 9 2
7 9 1 9 13 3 0 2
19 3 10 9 1 14 13 10 0 9 7 9 1 9 13 1 9 1 12 2
24 7 10 10 15 1 10 0 9 13 9 9 2 4 10 9 0 13 1 0 1 9 15 13 2
17 11 4 0 13 10 0 2 9 2 1 10 10 0 7 0 9 2
15 15 13 3 0 14 13 10 0 9 9 2 11 1 9 2
21 15 15 10 9 13 1 9 1 9 2 13 10 10 15 1 9 13 1 9 9 2
4 9 4 13 2
8 11 11 4 13 9 1 11 2
21 15 13 1 15 15 13 2 1 2 7 13 0 3 1 15 15 13 2 1 2 2
22 15 15 1 13 0 4 3 13 9 2 1 0 10 10 9 1 9 1 9 1 15 2
13 16 11 11 13 9 1 9 2 13 15 10 0 2
4 9 13 0 2
12 15 13 11 7 9 0 1 9 0 1 9 2
5 7 9 4 13 2
9 9 4 13 7 0 13 9 9 2
6 9 7 9 13 0 2
17 1 9 13 0 15 0 9 2 16 9 7 10 9 0 4 13 2
24 11 2 11 2 13 1 10 9 9 1 9 1 0 1 9 15 13 9 2 7 12 1 9 2
17 15 4 13 1 9 3 0 16 15 4 13 2 10 0 9 2 2
17 9 13 0 15 7 13 9 1 14 13 10 0 0 1 0 9 2
22 1 9 3 4 9 9 13 1 12 9 1 12 1 12 9 1 12 2 1 1 11 2
9 9 4 13 9 2 9 1 9 2
10 9 13 1 10 9 1 10 0 9 2
45 9 7 9 11 11 13 1 11 11 11 16 10 0 9 3 4 4 13 1 10 9 1 9 16 9 1 0 9 13 0 0 1 10 9 2 3 10 9 16 10 0 1 9 13 2
7 1 14 13 11 1 12 2
18 2 13 15 10 9 1 9 0 9 16 9 13 1 0 9 2 2 2
20 1 10 9 9 13 7 9 0 9 1 9 0 13 2 13 9 3 1 9 2
24 9 13 10 9 2 16 10 0 9 13 0 9 13 1 9 15 13 2 9 2 0 1 9 2
25 11 11 11 12 13 3 0 16 9 13 9 9 16 9 1 12 4 13 15 1 9 1 0 9 2
8 9 1 9 13 1 0 9 2
20 1 10 4 9 13 15 0 0 1 10 9 1 14 13 15 10 0 0 9 2
6 7 9 4 3 13 2
13 11 4 13 1 12 9 1 9 1 12 1 9 2
14 9 1 15 9 13 7 15 9 13 1 13 3 0 2
9 16 10 9 1 11 3 13 15 2
12 2 15 13 16 15 4 13 10 12 9 2 2
7 15 13 15 0 9 1 2
16 15 4 15 13 9 1 16 15 3 13 2 13 15 1 11 2
8 4 9 3 13 1 1 9 2
8 4 11 11 13 1 1 9 2
8 9 1 0 9 13 3 0 2
6 3 11 11 13 15 2
15 15 13 0 10 1 9 1 16 9 11 13 10 0 9 2
20 11 4 13 10 9 9 11 11 13 1 1 0 9 16 10 0 9 13 15 2
18 9 1 9 13 1 9 0 1 10 9 2 7 15 13 0 0 0 2
22 9 11 13 0 9 1 15 15 4 13 16 10 9 13 15 1 9 1 10 0 0 2
14 9 2 9 1 9 2 9 1 9 7 14 13 9 2
21 10 0 9 11 11 2 0 1 10 9 1 10 0 9 2 13 0 9 1 9 2
9 11 11 13 0 1 9 9 1 2
27 2 15 13 14 13 10 9 1 14 13 0 9 1 9 2 3 3 1 0 9 2 7 3 1 11 2 2
20 9 9 13 0 14 13 1 10 0 9 0 9 1 14 13 7 13 10 9 2
5 3 13 15 10 2
8 13 9 2 0 9 1 9 5
3 1 9 2
3 9 13 2
2 11 2
4 1 9 1 2
16 0 9 13 1 2 16 15 1 10 0 13 1 10 0 9 2
10 1 9 9 4 11 1 9 13 0 2
17 0 4 15 13 1 1 10 0 9 7 13 1 15 10 9 13 2
13 11 7 11 1 0 7 0 9 13 1 9 11 2
18 9 15 0 3 13 1 9 2 4 13 10 9 1 9 1 0 9 2
22 1 9 13 7 0 7 0 9 10 0 9 2 13 11 11 2 9 1 11 1 11 2
12 11 7 11 1 0 7 0 9 13 1 9 2
11 1 9 4 11 13 15 1 1 9 9 2
13 1 9 1 9 15 4 13 2 13 2 9 2 2
15 2 15 13 1 9 2 1 10 9 1 14 13 1 9 2
18 15 13 16 3 9 3 4 13 1 9 1 10 9 1 14 13 9 2
7 2 15 13 2 13 11 2
10 2 9 4 3 13 3 10 0 9 2
7 0 15 13 15 1 15 2
38 10 1 9 13 3 16 0 10 9 4 13 15 1 0 9 2 3 10 0 2 7 9 1 9 16 0 0 13 2 16 15 3 13 0 1 0 10 2
11 10 9 10 10 9 13 2 13 1 12 2
10 10 9 4 15 13 1 1 0 9 2
7 3 13 0 0 7 0 2
21 10 9 1 9 9 1 9 1 11 13 1 15 15 15 13 1 10 9 0 9 2
11 10 0 9 4 13 1 9 1 0 9 2
16 2 3 13 15 1 9 7 13 1 9 1 9 2 13 11 2
9 0 0 1 9 4 13 1 9 2
8 9 2 9 2 13 2 9 2
8 10 0 9 13 10 0 9 2
24 9 13 9 2 9 13 9 2 9 13 9 2 7 2 1 10 10 9 1 10 10 2 9 2
13 10 9 13 1 9 7 13 1 1 9 1 9 2
8 9 2 9 2 9 2 9 2
17 2 15 13 9 1 16 10 9 4 4 13 1 10 9 1 9 2
12 2 12 9 1 11 13 10 9 2 13 11 2
31 10 1 9 0 9 13 15 14 13 11 2 11 0 9 2 15 13 1 1 12 7 1 10 4 13 1 10 9 10 9 2
11 3 13 15 3 11 1 9 3 1 12 2
31 2 11 13 3 0 1 15 2 16 15 13 3 0 1 16 15 13 10 0 9 1 9 1 9 1 10 9 2 13 11 2
13 3 13 15 10 9 1 11 2 9 0 1 11 2
10 3 4 15 13 9 1 10 0 9 2
16 9 0 9 4 13 0 9 1 3 0 1 1 9 15 13 2
4 2 10 9 2
32 1 15 15 4 13 1 12 2 13 9 0 0 2 7 1 10 0 1 9 1 9 13 10 9 1 0 9 1 2 13 15 2
25 15 13 10 0 9 15 13 16 10 0 4 13 9 1 9 16 15 3 0 4 13 9 1 9 2
12 1 9 13 10 0 1 15 10 10 0 9 2
21 2 15 13 1 10 9 2 7 13 3 10 9 1 14 13 15 0 2 13 11 2
6 4 13 9 1 9 5
7 11 13 1 9 1 11 2
18 11 0 9 13 9 16 10 0 9 11 4 13 1 9 1 0 9 2
22 2 15 4 3 13 9 1 9 1 9 0 2 13 9 1 9 2 11 11 1 11 2
14 15 13 0 9 9 4 13 9 1 9 1 10 9 2
16 1 11 13 15 3 9 1 9 2 7 9 4 13 1 0 2
26 2 10 0 9 11 4 3 13 1 9 1 2 7 15 4 3 4 13 1 14 13 9 2 13 15 2
15 9 1 11 2 11 11 2 13 15 13 0 1 9 1 2
30 2 15 13 3 1 1 16 15 13 0 9 7 9 1 9 2 7 15 13 3 15 13 1 14 13 9 2 13 11 2
9 11 13 3 1 9 1 11 9 2
6 9 1 12 9 13 5
18 9 1 9 4 15 13 12 9 1 10 9 1 11 12 9 1 11 2
18 0 4 15 13 10 9 11 12 15 0 13 1 9 1 10 12 9 2
11 10 10 9 4 9 0 13 10 9 1 2
19 9 1 11 4 13 10 9 2 7 13 0 0 1 9 1 10 12 9 2
4 1 0 9 5
2 9 2
2 0 2
2 9 2
27 10 12 0 9 4 13 10 9 15 3 7 0 13 10 9 1 15 15 3 13 1 9 1 9 1 9 2
26 9 2 15 13 0 9 1 9 2 4 13 1 16 0 9 13 1 9 7 4 13 0 15 15 13 2
38 10 12 0 9 11 11 7 11 11 15 13 3 1 9 1 11 2 11 11 11 2 2 13 3 10 0 0 9 1 9 2 7 1 0 7 0 9 2
18 9 4 13 1 15 2 16 10 12 4 13 15 1 9 1 9 9 2
13 1 9 15 3 13 2 13 15 3 9 1 15 2
21 9 15 13 2 1 2 9 2 7 2 0 11 2 7 2 11 2 2 13 15 2
30 0 9 10 1 10 12 9 1 9 1 11 2 7 10 0 7 0 9 15 13 15 2 13 10 9 1 3 9 13 2
12 3 4 15 13 9 1 10 9 9 4 13 2
22 9 13 14 13 10 3 0 9 1 0 1 15 15 13 10 9 15 13 15 1 11 2
9 7 15 4 13 9 1 9 9 2
37 13 9 1 16 10 0 9 13 0 2 16 15 4 13 1 9 1 0 9 7 16 15 2 15 15 13 1 11 9 2 13 9 1 2 9 2 2
21 10 0 15 13 15 1 9 1 10 9 2 13 3 13 15 15 3 13 9 9 2
25 15 15 13 11 9 1 10 9 2 4 0 13 15 1 9 1 10 9 15 3 13 10 9 1 2
27 15 4 3 13 9 1 0 1 15 15 13 1 9 1 1 10 9 2 1 10 9 16 15 13 0 9 2
21 16 15 4 13 2 13 15 3 9 1 16 10 12 13 10 0 9 1 10 9 2
14 15 13 0 16 9 13 2 7 15 13 10 9 3 2
14 10 12 4 13 0 9 2 7 15 13 9 1 9 2
12 11 13 0 0 7 1 9 0 1 10 9 2
6 11 0 0 7 0 2
28 3 13 15 10 9 1 10 9 15 3 3 0 2 7 0 4 4 13 10 9 2 1 9 1 10 0 9 2
11 1 9 1 10 9 1 9 13 15 9 2
28 1 10 12 9 0 9 15 13 15 1 10 0 0 9 2 7 16 11 9 1 0 0 9 13 1 10 9 2
9 10 12 9 0 9 13 1 0 2
9 9 7 9 1 9 4 13 1 2
6 9 13 10 0 9 2
15 15 13 9 1 10 9 1 9 15 3 7 0 13 9 2
16 1 9 4 9 3 3 13 10 0 9 10 12 0 4 13 2
43 7 13 1 9 1 9 9 2 7 9 9 2 13 15 3 14 13 16 15 4 2 13 2 10 9 1 1 10 9 7 9 15 4 13 11 1 11 0 9 7 0 9 2
4 9 1 9 5
4 10 0 9 2
4 11 9 10 2
4 11 9 10 2
3 11 9 2
4 0 9 10 2
2 9 2
17 9 4 13 10 0 9 1 11 2 9 0 9 1 9 7 9 2
10 7 11 0 9 1 0 9 4 13 2
47 2 11 1 10 0 2 13 9 1 10 9 1 10 0 9 11 11 1 9 1 9 1 11 0 9 2 11 2 15 3 13 3 1 11 2 9 1 10 9 1 11 7 10 9 1 11 2
30 9 1 9 11 7 11 13 10 9 1 12 9 7 9 2 10 9 9 7 10 3 0 9 1 0 9 7 0 9 2
37 11 7 11 2 15 1 9 1 11 2 4 1 9 1 12 5 12 13 10 0 9 15 13 1 1 9 1 11 10 9 2 0 1 11 7 11 2
32 10 0 9 4 9 13 10 0 9 1 9 2 0 1 9 1 10 12 0 9 1 9 2 11 2 1 11 1 12 9 3 2
10 0 13 16 15 0 4 13 1 9 2
21 11 13 1 11 13 9 1 9 15 0 9 2 7 10 9 11 3 2 0 13 2
32 11 2 0 13 1 11 7 1 9 3 1 11 2 13 1 0 9 0 1 14 13 7 10 0 9 7 10 0 9 1 9 2
17 3 13 10 0 9 0 1 9 11 1 12 9 1 16 11 13 2
34 10 0 12 9 13 11 9 1 10 0 9 2 16 10 0 9 2 9 11 11 1 12 13 9 1 10 0 9 1 10 0 0 9 2
17 9 7 10 9 4 13 11 7 11 3 3 0 2 7 3 0 2
37 3 0 4 15 13 1 1 11 2 0 10 0 9 2 15 1 12 13 1 9 1 14 13 9 1 11 2 7 11 2 15 4 13 0 0 0 2
25 3 3 1 11 2 9 1 1 12 9 9 2 13 15 0 13 3 0 9 4 13 10 0 9 2
17 9 13 16 9 4 13 11 2 7 1 10 9 13 11 0 9 2
28 15 13 1 1 1 16 11 1 0 13 1 10 9 0 9 1 0 2 0 9 7 9 1 10 3 0 9 2
22 1 10 10 0 9 4 11 13 1 9 1 11 2 1 9 3 13 1 10 0 9 2
17 10 0 9 13 9 1 12 2 16 11 13 9 3 9 4 13 2
24 9 2 13 1 9 1 0 9 15 13 14 13 0 1 10 0 9 2 13 10 9 1 11 2
26 11 13 16 10 0 9 13 1 0 9 1 9 1 9 2 7 13 9 1 9 1 0 9 7 9 2
15 15 13 3 10 9 1 11 1 10 10 2 0 0 9 2
23 9 1 9 13 3 0 16 11 9 13 15 3 0 16 9 4 13 10 9 15 4 13 2
9 15 13 10 9 0 9 13 15 2
6 11 13 15 0 9 2
18 15 13 16 9 13 9 9 2 3 16 15 13 10 0 9 1 9 2
20 15 13 0 9 2 15 3 4 13 1 1 11 2 7 1 9 1 0 9 2
13 10 9 15 3 13 3 2 4 3 13 10 9 2
22 9 1 0 9 2 15 11 4 13 10 0 9 1 2 13 1 1 14 13 9 0 2
13 3 13 11 3 10 10 9 2 7 3 10 9 2
8 9 4 13 10 15 1 9 2
10 0 13 9 1 9 1 14 13 9 2
46 7 16 9 1 10 9 1 11 1 9 13 1 14 13 0 1 0 9 1 9 2 13 15 3 0 14 13 9 1 11 9 1 14 13 9 9 12 9 9 2 10 9 1 11 9 2
9 10 9 13 3 0 1 10 9 2
21 11 0 9 7 9 2 10 0 0 9 11 11 2 13 9 7 10 0 0 9 2
20 11 13 3 16 11 0 2 0 9 4 13 11 1 9 1 10 0 0 9 2
14 1 9 1 14 13 1 13 15 9 2 1 10 9 2
9 15 13 11 9 1 9 1 11 2
36 3 1 11 4 15 1 9 2 1 11 9 7 11 7 11 9 2 13 16 10 0 9 0 7 0 0 0 9 2 11 2 0 4 4 13 2
29 3 4 10 0 9 1 9 13 1 16 11 13 10 9 2 1 1 0 0 2 1 9 1 10 0 0 0 9 2
17 7 15 13 16 11 0 13 9 0 1 9 2 1 9 1 11 2
14 7 9 4 13 15 1 14 4 13 0 0 1 9 2
17 10 9 16 12 1 10 12 9 1 11 13 0 2 13 15 9 2
18 9 4 3 13 1 9 1 15 2 7 10 0 9 1 9 13 0 2
9 15 13 1 9 1 1 11 9 2
13 15 13 3 3 10 0 12 9 9 15 4 13 2
7 15 13 10 3 0 9 2
20 10 0 10 12 9 4 13 0 1 10 0 9 1 10 0 9 9 0 9 2
9 15 13 11 15 13 9 0 9 2
3 0 9 5
12 15 13 3 9 9 16 9 13 10 0 9 2
11 15 13 0 9 15 13 15 2 13 9 2
8 1 11 11 11 2 12 2 2
18 15 15 13 0 1 9 2 13 3 3 0 1 9 4 13 15 0 2
4 13 9 3 2
44 11 13 10 1 11 0 9 2 15 4 13 9 9 1 11 2 7 15 13 3 1 1 9 16 0 9 13 15 10 0 9 7 10 9 1 14 13 1 14 13 0 1 9 2
27 0 0 9 15 13 9 1 9 2 15 15 13 1 1 11 2 2 13 2 3 1 10 9 1 0 9 2
13 7 15 13 3 9 9 16 9 13 10 0 9 2
8 15 13 0 9 15 13 15 2
13 7 1 15 10 13 3 0 9 7 0 7 0 2
5 15 4 3 13 2
5 1 9 1 9 5
11 11 11 11 13 10 1 11 0 0 9 2
27 1 10 0 9 1 9 2 9 7 9 4 15 13 9 1 15 1 10 0 1 10 9 15 4 4 13 2
25 1 9 1 11 11 0 9 13 15 15 0 3 0 0 1 9 1 1 9 2 15 13 1 9 2
18 1 9 1 11 9 13 15 9 1 10 9 15 4 13 0 0 9 2
23 10 0 9 11 13 1 10 9 2 13 0 1 16 15 13 10 1 9 11 0 0 9 2
18 1 9 7 9 13 15 10 0 9 1 9 1 9 1 10 0 9 2
33 7 1 10 10 0 9 2 9 1 10 0 9 7 9 2 9 2 2 13 9 1 11 1 9 0 0 16 15 3 4 13 15 2
17 10 9 13 15 3 14 13 16 9 13 15 1 1 11 7 9 2
13 9 1 9 13 16 11 3 13 0 1 0 9 2
28 15 13 9 16 15 1 0 9 1 10 0 9 13 1 9 1 9 2 16 9 4 13 0 1 9 1 9 2
14 7 9 1 14 13 9 1 9 4 3 13 1 10 2
11 11 4 13 9 10 0 0 9 1 9 2
24 10 0 1 11 0 9 13 3 16 15 13 14 13 10 0 9 1 14 13 1 10 0 9 2
31 12 9 1 16 15 4 13 11 16 15 13 14 13 1 2 13 15 1 11 7 10 9 16 15 13 1 14 13 1 9 2
24 9 13 14 13 9 1 9 1 9 1 10 0 9 2 7 11 4 4 13 11 9 1 9 2
16 15 13 9 1 16 10 9 3 4 13 0 1 10 0 9 2
15 7 15 4 13 9 14 13 0 1 9 9 1 10 9 2
12 7 15 13 10 0 9 16 10 9 3 13 2
8 3 13 11 1 10 0 9 2
26 15 13 0 16 10 3 0 9 13 3 0 1 1 10 9 1 16 9 9 3 13 1 14 13 1 2
17 7 15 13 0 16 9 3 4 13 10 9 11 4 13 9 9 2
10 15 13 9 1 3 11 10 9 13 2
3 9 9 5
18 15 13 0 3 0 16 0 9 13 14 13 15 1 1 10 0 9 2
30 3 4 11 13 9 1 14 13 1 9 1 10 0 9 1 11 2 16 0 0 9 1 12 0 9 4 4 13 9 2
28 9 4 4 13 1 12 9 2 7 1 9 4 9 4 13 15 1 9 1 9 2 0 13 1 12 0 9 2
9 11 13 0 1 16 9 13 0 2
32 9 4 4 13 1 16 9 4 13 9 2 7 1 9 1 11 4 9 4 13 1 16 10 0 9 4 4 13 1 0 9 2
26 10 0 7 0 9 4 13 16 9 4 13 10 9 0 9 1 10 9 2 9 15 9 3 3 13 2
35 7 1 9 1 14 13 0 9 2 13 10 0 9 16 15 3 4 13 9 2 7 16 15 2 0 1 10 9 2 3 13 9 1 9 2
14 1 14 13 9 13 10 9 0 1 0 9 1 9 2
25 16 11 13 9 1 10 0 9 1 16 9 13 16 9 3 4 13 2 13 15 10 9 1 15 2
35 7 16 11 1 10 9 13 16 2 15 13 3 0 15 13 1 16 9 4 4 13 1 0 9 2 2 13 9 9 1 9 1 10 9 2
9 10 9 1 9 2 9 7 9 5
11 9 11 11 13 10 0 9 1 11 9 2
11 0 13 9 10 1 10 0 1 9 9 2
12 11 4 13 9 0 0 9 3 1 0 9 2
35 1 9 1 0 1 12 9 1 11 0 9 4 15 13 10 9 0 9 2 7 4 3 13 14 13 9 1 10 0 9 15 15 13 1 2
17 9 1 9 13 3 0 9 0 2 16 10 9 4 13 1 9 2
18 3 16 15 13 9 2 13 15 16 15 13 14 13 3 0 1 9 2
25 9 9 13 1 15 10 9 1 10 0 9 16 11 3 13 15 1 10 0 9 1 10 0 9 2
17 15 13 16 9 0 9 3 3 13 9 2 7 3 9 1 9 2
27 10 10 9 13 0 0 2 16 9 4 13 7 10 0 9 1 9 2 9 7 9 4 13 0 10 9 2
32 3 4 11 3 13 10 0 9 1 14 13 1 10 0 9 1 0 9 15 13 11 9 1 9 11 11 11 7 9 11 11 2
13 9 1 9 1 10 0 1 10 0 4 0 13 2
25 11 13 1 9 1 1 10 9 15 3 3 13 9 0 0 2 7 15 3 13 9 9 7 9 2
24 9 1 11 0 9 13 3 3 16 0 0 9 1 12 9 13 16 10 9 13 0 1 9 2
41 3 16 9 1 11 9 13 0 1 14 13 10 9 2 4 11 1 10 9 13 1 14 13 9 1 10 0 9 1 16 9 3 13 10 1 10 0 9 1 11 2
25 9 13 0 1 11 0 9 1 10 9 1 9 2 15 4 13 9 1 10 0 9 1 0 9 2
13 10 9 13 3 9 10 0 9 1 11 11 9 2
17 9 9 13 10 0 1 16 11 11 13 1 9 1 11 11 11 2
22 9 1 11 13 15 1 0 1 10 0 9 9 2 16 9 4 13 1 0 0 9 2
26 15 13 3 14 13 1 10 0 9 11 11 1 12 7 11 11 2 9 1 9 1 11 2 1 12 2
25 9 1 11 13 3 0 1 9 1 11 0 9 11 11 1 9 7 11 0 9 11 11 1 12 2
17 1 10 9 13 9 1 10 9 1 0 9 1 9 1 0 9 2
19 15 13 0 3 10 0 16 9 13 14 13 0 9 15 13 1 0 9 2
27 10 0 9 1 10 0 9 11 11 11 1 12 13 1 10 0 9 14 13 9 1 9 0 0 0 9 2
28 9 4 1 9 3 13 1 9 1 9 1 11 2 9 1 9 1 10 0 11 7 9 1 10 9 1 11 2
13 1 10 0 9 13 3 9 15 13 1 9 9 2
8 11 13 12 9 1 10 9 2
30 10 0 9 1 11 13 3 1 9 2 16 9 7 10 9 13 3 1 1 10 0 9 1 15 15 4 13 1 11 2
23 1 9 13 10 0 0 9 1 9 1 14 13 10 9 15 11 7 10 9 13 1 9 2
18 9 13 0 2 3 0 16 9 4 13 9 7 9 1 10 0 9 2
12 16 9 13 2 4 10 0 13 1 0 9 2
16 11 13 10 0 9 1 10 9 2 7 4 13 9 1 15 2
23 7 15 13 9 1 16 9 1 11 9 13 9 1 14 13 10 10 1 10 0 7 0 2
13 11 13 9 1 14 13 0 9 1 10 9 1 2
3 9 9 5
41 10 0 9 1 10 0 11 4 13 1 10 9 15 13 14 13 0 2 0 9 7 10 9 15 2 1 9 1 11 2 13 0 3 0 0 1 9 1 1 9 2
21 15 13 0 1 10 0 9 1 9 1 0 9 2 7 13 3 1 0 0 9 2
21 11 13 3 0 16 15 13 0 9 1 14 13 0 9 1 10 9 1 1 10 2
17 0 13 9 16 15 13 3 0 1 10 0 9 1 9 1 1 2
16 15 13 0 7 0 9 15 13 0 1 14 13 9 1 9 2
45 11 0 0 9 2 11 11 2 13 3 3 0 9 16 15 1 10 9 1 7 9 11 11 7 9 11 11 13 14 13 9 1 9 1 9 16 9 13 0 9 1 9 1 9 2
41 15 13 11 13 10 0 9 16 15 13 9 3 13 0 0 1 10 9 9 7 1 9 7 9 4 13 1 9 9 2 1 1 10 9 1 10 9 1 12 9 2
27 15 13 3 0 1 9 1 16 9 1 10 0 9 1 9 13 16 9 3 13 0 9 7 9 1 0 2
11 11 11 13 3 1 1 14 13 10 9 2
50 10 9 1 16 11 9 1 9 3 13 10 0 9 2 13 12 1 0 9 15 13 1 16 11 3 13 0 0 1 3 15 3 4 13 0 1 3 15 4 13 0 9 1 14 13 0 1 10 9 2
27 10 0 9 1 9 13 3 16 11 3 4 13 1 9 16 15 3 4 13 0 3 1 10 12 0 9 2
38 15 13 0 9 16 9 1 9 7 4 13 1 9 7 1 9 11 9 1 9 1 9 9 2 7 16 15 4 13 3 0 9 1 14 13 0 9 2
19 9 13 10 9 16 15 13 16 9 13 10 9 1 0 9 1 0 9 2
35 7 15 13 0 1 14 13 0 1 10 9 1 9 9 15 13 15 1 3 0 9 4 13 1 14 13 9 7 13 9 1 9 1 9 2
19 1 0 9 13 15 16 10 9 1 9 3 4 13 1 10 9 15 13 2
4 9 13 0 5
18 11 9 11 11 4 13 0 9 1 10 9 1 9 1 11 0 9 2
21 10 0 9 2 10 0 9 11 11 2 4 0 13 10 0 9 1 10 0 9 2
15 1 11 4 11 13 3 0 1 9 1 0 9 1 9 2
11 15 4 3 4 13 9 1 9 11 11 2
13 11 13 9 10 9 1 11 1 14 13 1 9 2
25 15 4 13 1 9 1 11 2 11 2 11 7 11 2 1 9 1 16 11 7 9 3 13 0 2
15 15 13 10 0 9 1 9 1 16 15 13 1 0 9 2
8 11 13 0 1 14 13 9 2
11 15 13 1 2 0 9 2 1 0 9 2
17 15 13 3 0 1 1 7 1 2 16 11 13 0 1 10 9 2
24 11 0 9 1 11 13 0 9 1 10 9 2 7 13 3 14 13 0 0 16 9 4 13 2
12 0 9 13 16 11 4 13 1 12 9 9 2
16 7 9 1 0 9 4 13 3 0 16 15 13 1 12 9 2
17 3 4 11 13 15 1 10 0 9 1 10 0 9 2 11 11 2
8 3 13 15 0 1 10 9 2
16 11 13 3 9 1 0 9 1 9 1 9 15 4 13 9 2
6 9 4 13 0 1 5
20 1 9 13 9 11 11 1 11 9 1 14 13 10 0 9 1 10 0 9 2
3 9 13 2
7 13 9 3 2 13 0 2
11 15 13 10 0 9 2 3 0 15 13 2
19 1 0 9 13 15 3 0 14 13 3 9 1 14 13 0 9 1 9 2
23 9 13 3 16 15 13 3 0 14 13 15 15 13 1 1 14 13 10 0 9 1 9 2
23 1 0 9 13 15 9 1 10 9 2 3 16 15 3 1 9 13 9 1 10 0 9 2
16 16 15 13 15 9 4 13 2 3 13 15 3 0 15 13 2
18 11 13 1 10 9 1 10 0 9 2 7 3 1 10 0 0 9 2
15 3 4 15 13 9 1 14 13 0 1 9 1 11 9 2
23 0 13 4 11 1 9 1 10 0 12 9 4 13 15 14 13 9 0 1 10 10 9 2
24 3 13 10 9 15 0 4 13 3 1 11 2 3 9 1 10 9 15 13 10 0 0 9 2
23 1 1 9 1 1 9 4 9 1 9 1 9 4 13 1 3 12 1 0 12 9 9 2
12 3 10 9 1 9 1 9 4 13 1 9 2
14 15 13 12 9 1 10 9 2 1 9 1 10 0 2
19 1 9 13 10 2 0 2 9 1 9 1 9 15 13 1 10 0 9 2
14 9 1 9 2 13 1 12 9 2 4 13 1 9 2
12 7 1 9 13 9 1 3 12 9 0 9 2
22 0 0 13 15 16 11 4 13 1 0 9 1 14 13 1 12 9 0 9 1 15 2
13 1 9 13 10 3 0 7 3 0 9 1 9 2
22 9 13 1 0 9 7 9 1 14 13 10 0 9 1 9 7 9 1 9 1 9 2
11 15 13 15 3 1 9 2 12 9 9 2
23 1 9 4 9 13 1 9 1 9 1 9 2 15 1 12 3 4 13 1 12 9 9 2
15 3 0 4 11 13 9 1 9 1 14 13 9 1 9 2
14 3 0 1 9 11 13 1 9 2 13 15 15 13 2
24 3 0 9 9 4 13 10 9 2 3 0 4 15 13 11 7 9 1 10 0 9 15 13 2
3 11 9 5
18 15 13 15 1 9 1 10 9 16 11 9 1 11 0 9 13 9 2
11 9 9 13 3 0 10 0 9 1 9 2
33 0 13 15 0 9 1 16 11 9 1 11 0 9 13 10 9 15 4 13 0 1 2 9 2 1 9 9 7 9 10 0 9 2
13 0 10 0 9 4 3 13 2 9 4 13 9 2
13 3 13 13 9 10 9 1 9 1 11 11 9 2
13 1 9 1 9 4 15 13 9 1 11 11 9 2
25 15 13 0 9 1 11 2 7 7 11 11 7 11 11 13 15 13 1 9 1 14 13 11 9 2
4 15 13 0 2
28 1 10 0 4 15 13 9 7 9 3 1 14 13 10 9 1 9 9 2 7 3 13 15 1 10 0 9 2
25 1 10 0 4 15 13 16 1 9 4 11 13 1 11 9 2 3 1 10 0 0 9 0 9 2
23 7 1 10 0 13 10 0 9 3 3 1 14 13 11 9 3 16 15 13 1 1 15 2
24 3 13 15 3 3 1 10 0 9 1 10 0 9 16 9 13 9 1 10 0 9 1 9 2
15 1 10 9 4 10 12 9 13 0 0 2 7 0 0 2
6 15 4 13 9 0 2
5 13 9 1 15 5
8 11 4 13 1 10 0 9 2
24 1 9 1 3 0 9 1 9 13 15 1 1 14 13 3 0 9 10 9 1 1 9 12 2
13 15 4 3 4 13 10 0 9 1 9 11 11 2
30 1 11 9 4 15 13 16 10 9 16 9 13 3 0 1 9 2 13 15 15 13 0 1 14 13 9 9 1 15 2
29 1 9 2 7 3 0 1 9 9 2 13 15 16 9 1 1 10 0 0 9 1 9 1 0 9 13 0 0 2
22 14 13 9 1 9 1 4 13 0 9 15 3 10 9 4 13 0 9 1 14 13 2
34 9 1 10 0 9 1 9 4 3 13 1 3 1 10 0 9 1 9 7 9 2 9 2 9 7 10 9 15 13 1 9 1 12 2
34 7 15 13 3 1 14 13 1 16 10 9 0 13 10 0 9 1 16 11 13 3 0 0 9 1 9 1 11 11 9 3 10 9 2
20 1 9 1 0 9 1 9 1 9 4 11 13 3 0 9 1 9 7 9 2
30 16 0 9 1 0 9 3 4 13 9 2 16 10 9 1 10 0 9 4 13 0 2 13 0 1 14 13 9 9 2
44 9 0 9 1 9 1 9 1 9 4 3 3 0 13 1 16 15 13 0 1 10 0 9 1 9 2 7 16 10 9 1 11 2 1 15 2 4 13 10 0 9 1 11 2
12 9 1 9 13 1 10 0 13 0 1 0 2
4 9 13 0 2
30 9 15 13 14 13 1 9 1 0 9 2 13 10 9 15 13 1 10 0 9 15 13 1 9 14 13 9 1 9 2
20 1 10 9 4 15 13 0 1 14 13 9 1 10 12 7 10 0 0 9 2
18 7 1 12 9 13 15 15 13 9 1 14 13 0 9 1 11 9 2
25 9 1 0 9 13 3 0 1 9 1 10 0 0 9 9 7 10 0 9 1 0 9 1 9 2
15 15 13 0 16 9 11 11 3 4 13 0 9 1 9 2
8 3 3 13 11 9 1 15 2
2 9 5
6 9 13 0 1 11 2
21 15 13 0 1 9 9 1 0 9 1 9 16 15 13 10 0 7 0 9 0 2
27 1 10 9 13 15 3 0 16 11 13 9 1 9 15 4 13 9 2 1 16 0 9 1 9 4 13 2
16 9 1 9 15 3 4 13 2 13 15 0 1 11 10 9 2
47 1 10 9 16 9 1 0 0 9 13 1 0 2 13 15 0 9 1 9 1 10 9 16 3 11 2 15 4 13 1 10 9 1 0 9 1 9 1 12 2 3 13 15 0 1 9 2
14 3 0 0 13 15 1 9 15 13 7 4 13 9 2
13 9 13 10 9 1 14 13 9 3 0 1 0 2
8 9 13 0 0 0 9 9 2
14 15 4 3 13 0 1 16 11 13 1 7 13 9 2
27 0 9 1 9 7 0 0 9 1 9 15 13 2 13 0 7 1 10 0 9 2 7 1 0 9 9 2
11 16 11 3 13 1 2 13 9 1 9 2
4 9 13 0 2
10 11 4 13 9 9 3 0 1 0 2
28 16 15 13 9 2 13 10 0 9 9 1 9 4 13 1 2 16 15 4 13 3 0 1 10 9 1 9 2
2 9 5
9 9 1 9 2 15 13 0 15 2
10 15 13 9 1 9 1 9 1 9 2
17 9 1 10 0 9 13 0 3 0 2 10 9 13 1 0 9 2
7 0 13 3 10 0 9 2
22 10 9 1 11 13 1 10 9 15 15 1 15 13 10 9 1 9 1 12 9 9 2
21 4 9 13 1 11 2 4 11 11 3 4 13 15 10 9 2 10 9 1 9 2
25 7 9 13 16 10 9 15 4 13 9 1 9 1 9 2 13 0 1 14 13 10 9 1 9 2
28 9 1 16 10 0 13 0 9 1 10 0 0 9 1 9 2 13 3 1 1 9 0 2 15 3 13 9 2
16 11 9 13 0 9 1 15 15 13 1 0 9 1 0 9 2
8 7 0 9 4 13 10 0 2
13 9 1 15 15 1 9 13 9 2 4 13 9 2
13 9 4 13 1 9 1 3 0 7 0 0 9 2
15 10 0 9 13 10 0 9 7 13 3 10 9 0 9 2
8 7 9 13 3 0 1 9 2
20 0 1 10 3 0 3 1 9 4 0 4 13 9 1 10 0 13 1 9 2
8 3 4 15 13 0 0 0 2
5 3 13 11 9 2
7 10 0 0 9 1 11 5
29 9 11 11 4 13 10 9 9 1 16 11 9 1 12 1 12 9 13 10 9 1 10 0 9 1 10 0 9 2
12 11 4 0 9 13 15 1 10 0 0 9 2
41 15 13 3 0 3 1 10 0 9 2 7 15 13 3 0 16 11 13 14 13 10 10 1 11 11 1 12 2 12 2 16 9 0 9 13 15 0 0 1 11 2
24 15 4 13 12 9 16 15 3 13 14 13 10 9 1 9 1 10 2 7 3 10 2 9 2
22 1 0 9 2 7 1 9 7 9 1 10 10 0 9 2 13 11 9 1 10 9 2
8 9 13 14 13 1 10 9 2
24 15 13 3 3 1 14 13 9 16 11 9 13 9 1 16 9 3 13 9 1 9 1 11 2
26 1 16 11 13 10 0 9 1 11 1 9 2 4 11 13 16 11 4 13 1 14 13 9 1 11 2
33 11 4 13 15 1 15 15 1 15 13 1 0 9 2 7 3 4 15 13 1 16 9 13 1 1 9 1 7 11 7 11 9 2
17 11 0 9 13 9 7 4 1 0 13 10 9 1 9 1 9 2
19 11 4 3 13 10 10 9 2 7 4 13 0 1 14 13 15 0 9 2
20 1 9 13 10 1 10 0 9 1 9 2 11 11 1 11 2 3 1 9 2
18 15 13 3 16 15 3 4 13 9 1 16 10 3 0 9 13 0 2
19 3 13 11 10 12 9 15 13 1 14 4 13 16 9 13 10 0 9 2
8 0 9 4 13 1 9 1 2
15 0 2 7 0 3 3 9 2 13 16 9 13 0 0 2
18 9 13 12 9 9 1 10 9 1 12 9 2 1 11 9 1 9 2
21 10 0 9 13 1 14 13 9 1 9 15 3 13 9 1 14 13 10 10 9 2
15 15 4 13 16 9 1 9 1 9 4 13 1 12 9 2
10 7 9 13 3 1 14 13 1 15 2
12 1 12 9 4 3 12 9 9 13 1 9 2
18 3 13 9 1 14 13 9 1 14 13 0 1 15 15 4 13 9 2
25 11 4 1 15 14 13 13 10 9 2 7 15 13 3 3 0 14 13 15 15 1 9 4 13 2
4 9 0 9 2
29 11 9 4 1 3 0 9 13 10 9 1 11 1 3 14 13 15 9 13 14 13 1 14 13 0 1 9 10 2
12 15 4 0 13 14 13 1 9 7 13 9 2
14 4 3 9 0 9 14 13 1 3 13 10 0 9 2
5 0 13 15 15 2
29 10 9 15 13 0 0 9 2 7 15 4 13 10 9 0 1 12 2 4 13 0 1 9 2 3 1 10 9 2
17 7 1 9 1 9 1 0 0 10 9 2 13 0 9 0 0 2
11 10 3 0 9 4 13 2 13 7 13 2
22 7 15 13 3 0 16 15 0 13 10 0 0 9 2 3 16 15 13 0 1 9 2
29 1 9 1 9 15 4 13 0 1 9 2 13 15 1 16 16 11 13 0 2 13 0 0 1 10 9 1 9 2
11 3 0 13 9 1 9 15 13 0 9 2
19 1 0 9 4 11 9 13 11 1 3 14 13 9 1 0 9 1 9 2
18 10 9 4 9 11 11 1 10 0 9 13 0 9 1 9 1 9 2
24 16 15 1 9 13 9 9 1 9 2 13 15 3 9 1 9 2 7 9 1 9 1 9 2
4 15 0 0 2
26 1 9 13 11 9 1 11 9 1 14 13 0 0 9 4 13 1 11 2 16 15 3 4 13 9 2
19 15 13 0 1 9 1 9 0 9 1 16 9 0 13 0 1 0 9 2
34 3 13 7 0 9 11 11 11 2 11 0 9 11 11 7 11 9 11 11 11 0 9 1 16 10 9 3 4 4 13 9 1 11 2
23 3 10 0 9 2 15 13 10 10 9 1 11 2 4 13 0 1 9 1 9 1 9 2
15 10 9 4 13 0 16 11 4 13 10 0 9 1 9 2
17 1 9 4 0 9 13 9 1 11 1 14 13 9 3 1 9 2
26 4 11 13 16 15 13 10 0 9 9 0 2 13 15 16 9 3 13 10 0 2 7 3 13 1 2
16 15 4 1 3 9 13 0 9 10 0 9 13 15 10 9 2
2 0 5
12 11 13 9 9 1 12 0 9 1 0 9 2
19 9 11 11 11 13 9 9 1 0 9 2 16 9 11 11 13 11 9 2
7 15 13 15 1 0 9 2
23 11 4 1 0 9 13 10 1 11 0 9 2 1 0 9 1 0 9 7 1 0 9 2
36 1 0 13 9 16 10 9 3 4 13 10 9 15 4 13 0 1 10 0 0 9 2 1 9 2 0 9 2 9 7 10 0 9 2 9 2
32 11 11 13 9 1 10 9 1 10 9 2 7 4 1 9 13 1 9 1 9 16 15 13 14 13 1 9 10 9 1 9 2
16 9 2 0 9 2 9 7 9 13 9 11 0 1 0 9 2
22 11 4 13 1 14 13 9 7 1 14 13 9 1 9 15 15 3 13 0 9 1 2
29 9 13 3 0 2 7 4 3 13 1 15 1 9 2 15 3 13 0 1 14 13 10 3 0 9 1 0 9 2
25 1 13 3 9 10 9 7 9 11 13 1 1 2 7 10 9 1 14 13 1 1 10 0 9 2
13 15 13 14 13 9 7 9 1 10 0 0 9 2
7 15 13 0 10 9 0 2
3 9 9 5
24 3 1 11 2 11 2 11 7 11 13 11 9 1 10 0 9 1 9 1 9 11 1 9 2
51 1 9 1 9 1 10 9 15 13 0 14 13 1 2 13 9 10 9 1 16 11 4 13 1 10 0 2 0 7 0 9 1 9 2 1 0 9 7 9 2 7 1 0 9 1 9 1 9 7 9 2
16 15 13 1 10 9 9 13 2 16 9 1 0 9 13 9 2
22 9 13 1 1 9 1 9 2 9 1 9 2 7 1 9 1 0 9 1 9 9 2
16 9 13 2 7 9 13 0 10 0 9 1 9 1 0 9 2
47 10 0 12 9 1 9 13 10 0 2 7 15 13 15 16 11 11 11 2 10 1 11 0 9 2 3 4 13 0 1 1 0 9 7 4 13 0 9 1 11 2 11 7 11 1 15 2
30 11 13 0 1 9 1 9 1 9 1 11 2 1 0 1 0 9 2 7 13 3 0 10 9 1 11 1 0 9 2
12 7 11 2 11 7 11 0 0 9 13 0 2
19 3 10 9 4 15 13 16 9 3 3 13 1 0 2 0 7 0 9 2
11 9 9 13 3 9 1 14 13 1 15 2
5 9 4 13 0 5
29 2 9 7 9 2 13 9 1 11 2 11 11 2 1 9 1 10 0 9 15 3 13 7 13 1 0 0 9 2
13 9 1 9 13 3 9 1 9 1 11 1 9 2
17 15 13 3 0 9 7 9 1 10 0 9 1 16 9 4 13 2
16 10 0 9 13 1 0 0 9 2 15 9 13 1 0 9 2
14 9 1 11 13 3 0 9 1 10 9 15 4 13 2
19 10 0 9 13 1 10 10 9 2 1 9 1 14 13 9 1 10 9 2
22 15 15 0 13 1 2 13 10 0 9 1 9 7 9 2 12 9 15 15 13 0 2
32 15 4 13 9 1 10 9 3 3 3 9 2 7 3 9 10 7 0 9 13 7 13 9 1 10 2 1 7 9 7 9 2
11 9 1 9 7 9 4 13 10 10 9 2
28 15 13 3 10 9 1 16 10 0 9 10 1 15 7 13 9 1 7 0 9 1 15 10 0 9 4 13 2
28 0 9 15 13 9 1 9 7 9 0 2 13 15 0 0 14 13 1 9 1 0 9 1 9 1 9 9 2
11 3 4 15 13 1 14 13 9 1 9 2
13 9 1 0 9 13 10 0 9 15 13 0 9 2
27 15 13 3 0 14 13 9 1 16 3 9 1 10 0 9 1 9 13 1 1 9 7 13 1 0 9 2
9 15 13 0 9 1 9 7 9 2
27 9 1 16 15 13 10 0 9 1 9 2 9 7 9 4 3 13 3 0 16 9 4 13 1 0 9 2
27 9 15 15 4 13 1 11 1 10 9 2 4 3 13 1 9 1 10 0 9 15 13 9 1 0 9 2
24 0 4 15 13 15 0 16 10 0 9 13 16 15 4 13 15 0 0 9 1 9 1 9 2
6 15 13 3 3 9 2
21 10 9 4 13 0 2 1 9 1 13 1 1 9 15 13 0 0 0 7 0 2
11 3 4 9 1 9 7 9 13 0 0 2
3 0 9 5
23 9 2 9 7 9 4 13 12 9 9 1 9 1 11 1 9 1 9 2 9 7 9 2
17 9 4 3 1 9 13 12 9 2 10 9 1 9 1 1 9 2
13 10 10 13 9 2 9 1 9 1 0 9 2 2
12 9 1 9 9 1 9 11 13 0 12 9 2
20 9 1 9 0 2 3 12 9 2 7 9 2 7 3 0 1 9 9 12 2
17 0 9 13 9 1 10 12 9 9 9 4 4 13 1 1 9 2
16 9 4 1 0 9 13 1 9 15 13 9 1 9 1 9 2
22 7 9 9 2 9 7 9 0 9 1 10 9 1 0 9 13 9 11 9 13 1 2
9 11 4 13 0 9 1 0 9 2
13 10 1 15 4 13 0 9 1 0 9 1 9 2
7 9 13 0 10 12 9 2
16 1 0 1 11 2 11 11 11 2 13 9 0 0 1 9 2
13 7 1 9 1 9 2 9 1 9 7 9 9 2
28 15 13 0 16 9 1 1 12 9 9 1 9 1 9 15 13 1 9 1 10 0 2 4 13 9 1 9 2
8 9 4 1 10 13 1 9 2
27 7 10 0 9 9 7 10 0 9 1 12 9 9 2 13 16 9 1 10 0 9 9 0 1 13 0 2
10 9 1 9 4 13 0 10 0 9 2
17 7 15 13 0 16 9 0 9 13 0 1 14 13 7 13 9 2
13 9 4 13 10 0 9 15 4 13 1 1 9 2
6 3 13 15 0 1 2
3 0 9 5
34 11 9 1 11 7 9 2 11 2 1 9 1 9 1 12 13 10 1 10 0 15 10 9 4 13 1 10 9 1 9 1 0 9 2
39 16 11 13 16 15 3 4 2 13 11 7 9 9 1 12 2 2 13 15 1 9 16 11 10 9 3 4 13 16 9 9 13 10 9 1 9 1 9 2
16 15 13 10 0 9 1 9 1 10 1 9 1 10 0 9 2
11 15 4 7 11 7 11 13 1 1 9 2
20 9 1 11 13 3 3 0 16 10 3 0 9 1 9 9 13 1 0 9 2
27 15 13 3 0 0 16 9 13 0 1 1 9 1 9 15 13 0 0 1 16 10 0 9 13 1 9 2
14 1 11 4 10 9 9 13 0 9 1 9 1 9 2
28 15 13 1 10 16 9 1 11 9 3 4 13 10 9 15 13 9 1 2 7 16 11 9 3 4 13 9 2
16 11 13 3 0 9 1 9 1 0 7 9 1 10 0 9 2
45 16 0 1 9 13 16 11 9 3 13 0 2 7 16 0 9 1 9 9 3 4 13 0 9 2 13 15 10 9 1 14 13 16 15 4 13 0 9 14 13 1 10 0 9 2
23 15 13 0 16 9 1 11 9 1 9 1 3 0 9 13 9 15 3 13 10 0 9 2
16 9 11 11 13 16 9 3 3 7 0 13 11 9 7 0 2
21 9 13 1 9 15 4 13 9 1 14 13 10 9 15 1 10 9 4 0 13 2
30 3 13 15 3 9 9 2 7 1 0 9 11 9 2 14 4 13 1 1 10 9 10 0 9 3 4 13 0 1 2
7 9 13 0 0 1 11 2
16 10 9 15 13 9 1 10 9 9 13 2 4 3 13 1 2
40 16 15 4 13 15 10 9 15 4 13 1 3 0 9 2 13 9 9 1 14 13 10 0 9 13 1 12 9 1 14 13 2 1 10 3 0 9 1 0 2
19 11 13 3 9 1 14 4 13 1 16 15 3 13 9 1 11 0 0 2
3 0 0 5
6 11 13 15 0 0 2
21 1 9 13 9 10 0 9 3 2 1 10 9 1 0 9 1 10 0 9 9 2
10 9 13 1 9 1 9 7 13 9 2
9 9 1 11 4 3 3 13 0 2
12 9 0 9 13 10 9 1 3 10 9 9 2
16 15 13 0 1 0 16 9 13 9 1 14 13 9 1 9 2
16 9 1 11 4 13 1 10 9 15 0 1 9 13 1 11 2
11 11 9 13 16 9 4 13 0 1 9 2
25 9 13 0 3 0 16 10 0 4 13 15 14 13 15 1 0 12 9 15 0 4 13 1 15 2
14 7 9 2 9 7 9 4 13 9 16 9 4 13 2
22 3 4 11 9 3 13 1 10 9 11 13 14 13 9 1 9 0 10 9 1 11 2
9 0 9 13 9 1 14 13 0 2
12 7 3 13 15 3 0 11 15 4 13 1 2
11 3 13 15 3 11 15 4 13 9 1 2
12 7 16 11 4 13 2 4 10 9 13 1 2
11 11 13 10 1 10 0 0 9 1 11 2
10 15 13 3 16 9 3 13 0 9 2
13 7 9 1 0 9 1 9 4 13 1 1 9 2
8 9 4 3 13 9 1 11 2
4 0 0 9 5
4 0 0 0 2
3 0 9 2
4 4 4 13 2
2 9 2
3 0 9 2
2 9 2
3 0 0 2
4 10 0 9 2
3 13 9 2
25 10 9 4 13 9 1 14 13 9 1 10 9 1 14 13 9 10 9 1 14 13 0 7 0 2
10 9 13 1 0 9 2 13 11 11 2
21 0 0 13 0 7 0 1 9 1 0 9 2 7 13 0 1 9 7 0 9 2
17 11 13 1 9 0 9 1 9 16 9 7 9 13 10 0 9 2
9 11 13 3 0 9 1 0 9 2
16 9 1 10 9 4 13 0 0 9 1 9 1 9 1 11 2
24 9 13 1 11 0 9 0 9 1 9 1 9 9 2 7 13 0 16 11 3 13 0 9 2
16 15 13 0 9 1 9 0 7 9 1 9 1 9 15 13 2
17 9 13 1 0 9 0 9 2 7 0 13 1 0 9 1 1 2
13 9 13 16 9 13 9 1 14 13 0 7 0 2
21 15 13 16 10 0 9 13 0 9 2 15 13 16 15 3 13 15 0 7 0 2
16 0 9 2 9 2 9 2 10 0 9 7 9 13 0 3 2
12 15 13 10 9 0 9 14 13 7 13 15 2
17 0 9 13 9 1 9 2 9 2 9 2 9 2 9 7 9 2
25 9 1 0 9 13 9 1 9 2 7 13 3 3 3 9 1 15 10 2 7 3 9 1 10 2
21 15 13 3 9 1 9 2 9 1 14 4 13 7 13 15 1 1 10 9 9 2
22 1 12 9 1 10 9 4 13 1 0 9 7 9 2 7 15 13 15 3 0 1 2
12 15 13 3 3 15 15 13 7 13 10 9 2
23 9 1 15 13 1 3 15 4 13 9 7 10 9 15 0 4 13 1 15 10 7 9 2
20 15 13 1 9 15 13 10 9 2 13 9 10 7 0 13 9 1 14 13 2
31 9 13 9 2 9 15 13 9 2 0 9 7 10 9 16 15 4 13 2 13 7 13 2 1 14 4 13 2 7 13 2
18 15 4 13 9 2 9 7 9 7 4 3 13 9 7 9 5 9 2
30 9 1 0 9 4 1 14 4 13 1 9 7 9 2 4 13 16 15 3 13 0 3 7 13 15 9 1 10 9 2
17 15 4 3 0 13 9 1 14 13 2 15 4 13 10 0 9 2
7 16 15 4 4 13 1 2
12 15 4 13 14 13 15 9 2 9 7 9 2
14 9 13 9 7 13 15 15 2 4 13 15 0 2 2
13 3 13 15 9 2 9 2 9 7 10 0 9 2
24 7 1 10 9 13 15 0 2 15 13 3 0 2 15 4 13 0 2 7 9 4 13 15 2
32 15 13 9 1 14 13 15 1 15 15 13 7 13 9 1 9 2 14 13 1 14 13 2 0 15 15 13 15 0 7 0 2
17 15 13 9 10 2 15 13 9 1 9 7 9 1 14 13 15 2
7 0 13 9 9 1 15 2
33 15 13 9 1 14 13 15 15 13 2 1 3 14 13 0 3 2 1 3 14 4 13 2 1 14 13 9 7 1 14 4 13 2
7 9 13 15 3 0 9 2
12 0 0 9 13 9 7 4 3 13 1 9 2
14 9 2 9 7 9 13 15 1 10 1 14 13 9 2
9 9 13 9 1 9 7 13 9 2
11 9 13 9 2 13 9 7 13 15 0 2
6 9 13 1 0 9 2
29 2 15 13 10 9 2 7 2 15 13 3 0 3 2 7 2 15 13 15 3 2 15 13 1 14 13 0 2 2
22 9 13 1 0 9 1 10 0 2 7 15 4 13 9 1 10 0 1 14 13 15 2
28 10 0 1 15 13 3 9 2 16 15 13 1 9 1 9 7 9 1 14 13 2 7 1 9 1 10 9 2
11 10 0 2 0 9 7 9 13 10 9 2
18 0 9 13 9 2 9 1 14 13 15 7 9 1 0 9 1 10 2
25 15 13 1 15 10 1 0 2 9 1 0 7 0 2 7 1 9 1 0 2 0 7 1 9 2
8 13 15 10 9 9 4 13 2
7 10 9 15 4 13 9 2
25 3 13 15 3 2 3 4 15 13 1 9 7 13 9 1 9 2 9 2 9 2 9 7 9 2
19 15 13 1 9 0 9 2 7 15 13 3 9 1 9 2 9 7 9 2
12 3 13 15 16 15 4 13 2 13 7 13 2
19 15 4 13 1 9 1 14 4 13 2 7 3 1 9 1 14 13 9 2
12 7 15 4 13 1 9 2 1 9 7 9 2
22 13 15 0 16 15 13 0 7 0 2 0 1 3 14 13 15 7 3 13 0 3 2
13 10 9 13 3 9 1 16 9 7 9 0 13 2
6 3 13 15 3 9 2
14 15 15 13 9 1 9 7 0 9 2 9 7 9 2
10 9 9 13 14 13 9 1 1 9 2
11 3 14 13 9 0 2 7 13 1 9 2
18 16 9 2 0 1 0 9 2 13 9 1 9 13 15 0 0 0 2
27 1 2 16 0 7 0 9 13 0 2 7 2 16 15 13 1 10 9 16 15 13 0 1 10 0 2 2
14 15 4 13 0 0 2 7 3 4 15 3 4 13 2
22 16 15 13 10 9 1 10 9 2 13 15 3 3 9 2 7 15 13 3 15 10 2
11 14 13 1 1 15 15 13 2 13 0 2
4 15 13 9 2
17 9 4 4 13 2 0 4 3 13 16 9 13 0 16 15 13 2
9 9 1 0 9 2 13 0 9 2
13 15 13 9 2 7 15 13 3 1 9 7 9 2
21 15 13 3 9 2 15 13 3 2 15 13 3 2 7 15 13 15 9 7 9 2
18 15 13 15 2 15 13 1 9 7 9 7 15 13 0 7 0 9 2
12 15 13 10 2 7 13 0 1 9 7 9 2
17 15 4 13 16 10 9 13 0 7 16 15 13 0 0 1 10 2
12 13 15 3 10 9 7 10 9 15 4 13 2
9 4 15 3 3 13 10 0 9 2
30 10 9 1 0 9 2 9 7 9 2 0 9 2 9 2 0 0 7 0 2 7 9 15 13 1 0 9 1 15 2
16 10 9 13 1 10 0 9 2 10 9 15 4 13 0 9 2
21 9 1 14 13 9 1 10 9 1 14 13 9 10 9 1 14 13 0 7 13 2
21 15 13 3 3 14 13 16 15 13 0 2 9 4 3 13 9 1 14 13 15 2
22 15 4 13 10 10 9 2 10 10 9 1 9 2 9 1 10 9 7 0 0 9 2
4 13 15 9 2
6 15 13 9 14 13 2
7 1 9 1 10 10 9 2
4 1 0 9 5
17 10 9 15 13 1 11 2 13 15 15 14 13 1 9 3 1 2
16 3 4 15 13 15 1 14 4 0 13 1 10 0 0 9 2
10 13 9 1 11 11 11 1 9 12 2
6 10 9 13 3 0 2
11 2 15 15 13 0 2 9 13 10 9 2
16 3 13 15 0 14 13 16 9 9 13 9 1 10 0 9 2
6 3 13 15 3 15 2
21 11 7 11 13 9 15 13 1 0 2 13 0 7 13 15 7 10 9 1 0 2
10 0 13 3 1 9 1 11 7 11 2
18 3 11 4 13 15 1 9 9 16 15 13 10 9 7 13 1 9 2
14 10 0 9 1 11 1 9 13 15 15 15 13 1 2
16 3 1 13 15 3 1 16 15 13 16 15 13 3 0 9 2
21 11 13 10 9 1 10 1 3 9 1 9 2 7 13 0 10 0 1 10 9 2
8 10 0 9 13 14 13 11 2
6 15 13 3 10 9 2
10 7 3 11 13 10 9 1 0 9 2
21 9 1 14 13 9 13 3 0 2 7 3 13 15 0 1 9 1 10 0 9 2
16 15 13 3 11 9 1 14 13 9 1 11 0 2 9 13 2
10 1 9 13 15 0 9 1 0 9 2
12 15 13 10 0 9 1 9 7 10 0 9 2
28 4 11 13 10 9 1 9 1 10 0 9 1 10 9 2 4 11 9 13 1 0 0 0 9 2 3 9 2
20 1 9 13 0 9 1 9 2 15 4 13 0 1 10 2 9 2 1 11 2
12 3 13 11 0 10 9 1 9 1 0 9 2
10 1 10 0 9 13 15 1 10 9 2
23 10 0 9 13 3 1 0 9 2 15 15 13 10 0 9 14 13 10 3 0 9 1 2
20 15 13 3 11 15 4 13 11 2 16 15 3 13 10 9 15 4 13 15 2
8 11 4 3 13 2 9 2 2
19 1 12 1 11 13 15 0 0 9 1 0 9 2 7 9 1 10 9 2
5 10 10 13 3 2
12 15 13 3 1 1 16 11 13 15 1 15 2
7 0 2 9 2 13 0 2
12 15 13 10 9 1 16 9 13 10 0 9 2
6 3 13 3 0 9 2
29 15 13 3 0 14 13 10 9 1 0 9 16 10 0 3 4 13 1 7 13 2 7 9 13 15 3 1 9 2
12 10 9 15 13 1 9 2 4 0 13 9 2
17 10 9 13 1 2 9 7 9 2 7 1 0 9 1 9 9 2
6 11 13 9 1 9 2
6 11 4 3 13 9 2
21 10 9 4 1 0 9 13 1 10 9 0 9 2 7 15 3 3 1 10 9 2
23 7 10 0 9 13 2 8 8 8 8 2 2 7 15 13 3 0 16 11 13 11 9 2
9 15 4 13 11 1 9 1 11 2
6 11 13 0 1 9 2
11 11 13 12 9 2 0 9 1 0 9 2
31 7 10 10 9 13 10 0 9 2 16 9 3 4 13 1 0 9 10 1 0 2 7 3 1 10 0 9 16 9 13 2
8 9 13 1 9 1 11 9 2
20 15 13 3 11 15 4 13 11 2 16 15 3 13 10 9 15 4 13 15 2
11 9 9 13 0 3 16 15 13 3 0 2
10 13 9 1 11 11 11 1 9 12 2
4 9 1 9 5
3 0 0 2
14 11 11 4 13 0 2 9 2 1 0 9 1 9 2
11 15 13 10 9 16 15 4 13 0 9 2
23 9 1 9 3 13 15 14 13 10 9 1 9 2 3 16 15 13 10 0 7 0 9 2
34 10 9 11 11 11 13 15 2 7 13 1 9 1 11 11 16 15 4 13 16 10 0 9 1 9 13 3 0 1 9 1 1 9 2
21 7 15 13 3 3 0 15 10 0 9 13 2 3 15 10 0 9 13 15 1 2
13 16 15 13 9 0 9 2 13 15 3 0 0 2
13 11 4 13 0 2 9 2 1 0 9 1 9 2
19 16 15 13 10 9 1 0 9 7 0 0 7 0 2 13 15 10 9 2
17 9 1 9 13 16 15 3 13 10 0 2 3 0 9 1 9 2
13 15 4 3 7 13 9 1 0 9 7 0 9 2
19 15 13 3 15 15 0 1 10 10 2 15 13 10 9 1 15 15 13 2
22 7 15 13 3 3 15 15 13 9 2 7 3 16 9 0 13 0 1 15 9 13 2
30 7 16 15 3 13 10 1 2 9 2 7 10 0 9 2 13 9 3 0 2 1 2 10 9 2 13 10 9 0 2
48 0 9 2 1 10 9 7 10 9 2 13 3 3 9 1 16 15 15 13 1 2 7 15 3 13 9 1 10 0 7 0 9 2 7 3 13 15 13 10 0 0 7 0 2 4 13 1 2
8 10 0 9 13 0 14 13 2
31 10 0 9 4 3 3 3 4 13 16 10 12 13 3 0 1 10 0 2 7 15 13 10 9 1 14 13 2 9 2 2
28 15 4 3 3 4 13 16 2 16 15 13 1 9 2 4 3 15 13 16 15 13 10 0 0 1 15 2 2
8 10 0 9 4 0 1 9 2
16 10 0 0 1 9 13 9 15 13 0 2 7 0 7 0 2
12 10 10 4 15 13 1 9 2 0 1 11 2
18 15 13 3 0 13 0 0 14 13 10 0 9 2 10 9 1 3 2
12 9 1 0 2 9 7 9 2 4 3 13 2
25 10 0 9 1 9 7 9 13 15 0 13 16 3 13 10 9 2 7 10 0 9 13 15 10 2
14 15 13 0 1 10 0 9 15 3 13 10 0 9 2
17 11 13 3 9 1 9 1 9 1 11 7 9 1 9 1 9 2
35 15 13 0 2 7 0 7 0 2 3 10 9 1 9 7 9 2 7 15 13 3 0 13 9 1 14 13 16 2 3 13 15 3 2 2
27 15 13 10 9 13 1 0 9 3 15 13 1 9 2 7 10 9 15 4 13 1 9 13 10 10 9 2
17 15 13 3 10 9 1 9 0 9 7 10 0 9 13 15 1 2
9 1 11 1 11 13 11 1 11 2
17 2 16 15 13 10 9 1 15 2 13 15 15 15 13 15 2 2
10 15 13 9 9 2 7 15 13 0 2
15 10 0 0 13 0 13 2 7 9 0 13 15 15 13 2
18 9 1 2 9 2 13 0 1 10 1 15 15 13 1 10 10 9 2
7 4 11 13 9 0 9 2
3 10 9 2
3 13 0 2
4 9 7 9 2
4 9 13 0 2
2 9 2
4 11 13 9 2
23 1 16 11 11 13 9 2 4 15 13 1 9 1 9 1 10 10 9 11 1 14 13 2
10 15 4 3 13 0 9 1 10 9 2
2 9 2
40 3 16 9 1 9 13 0 0 1 9 2 13 15 9 15 13 1 0 7 0 9 1 9 1 0 9 2 16 9 13 0 1 14 13 9 1 0 0 9 2
15 15 13 2 16 11 7 11 13 1 10 10 9 1 9 2
49 15 13 3 0 2 7 10 0 9 11 13 14 13 15 16 11 13 1 1 9 2 7 11 13 16 10 0 9 3 7 0 11 2 4 13 7 16 15 13 0 7 16 15 4 13 1 12 9 2
4 3 13 15 2
24 11 13 1 9 1 10 0 0 9 1 16 10 0 9 1 11 4 13 1 16 10 13 1 2
34 9 1 11 7 11 1 9 1 9 1 11 1 9 4 13 0 1 9 7 9 1 16 9 13 10 0 9 2 7 3 0 1 9 2
28 0 9 13 16 12 9 1 10 9 1 11 13 1 12 9 16 10 9 4 13 1 10 9 1 9 1 11 2
17 1 1 10 0 9 4 15 3 13 9 1 11 1 0 0 9 2
33 10 9 13 0 0 2 7 9 13 0 2 7 1 0 9 1 11 1 9 1 11 2 13 0 9 3 14 13 3 10 0 9 2
13 9 4 3 13 16 11 1 9 4 4 13 9 2
49 15 4 3 13 1 1 9 1 11 7 11 1 9 1 10 9 1 14 13 16 15 13 10 9 1 11 2 7 16 9 13 1 1 10 0 9 7 10 0 9 1 12 9 1 10 9 1 11 2
5 11 9 13 0 2
47 1 9 11 1 14 13 2 15 15 0 13 3 16 15 13 10 0 9 1 10 0 9 2 13 15 3 3 0 9 1 10 0 9 1 10 9 2 7 3 11 9 1 14 13 1 9 2
21 10 9 1 9 7 9 13 0 7 3 0 1 11 2 15 15 0 13 1 9 2
16 1 16 15 13 9 2 4 15 0 13 1 9 1 10 9 2
9 15 4 13 0 9 1 10 9 2
20 10 0 9 7 9 11 11 13 0 3 0 1 10 9 1 11 11 3 1 2
25 15 13 3 0 3 0 9 1 10 0 9 1 14 13 0 9 1 1 0 2 7 3 0 9 2
9 10 9 1 9 13 3 10 9 2
22 9 1 16 3 4 9 13 10 0 9 2 13 10 0 9 1 9 1 9 1 9 2
22 3 0 13 10 9 1 16 9 15 13 9 1 13 9 1 10 9 7 13 10 9 2
23 9 1 10 10 9 1 9 13 10 9 1 12 9 9 2 7 10 0 0 9 1 9 2
10 9 9 1 9 1 12 9 4 13 2
26 11 13 0 7 1 9 7 9 2 7 15 13 3 10 9 1 9 1 9 2 11 13 3 10 9 2
45 11 13 3 10 12 9 1 9 15 13 1 1 14 13 1 10 9 2 7 15 4 1 10 9 3 13 16 12 9 13 1 9 2 7 15 13 3 1 11 0 9 1 9 9 2
37 10 9 2 1 11 2 4 13 0 1 9 1 11 2 7 11 13 1 9 1 0 9 2 7 3 4 15 13 1 0 16 15 4 13 1 9 2
33 3 16 0 0 9 13 1 0 9 7 9 1 11 9 2 13 10 10 9 10 10 16 15 13 1 9 1 9 2 7 4 13 2
24 11 13 15 16 15 13 9 2 7 4 13 1 9 1 9 1 9 1 16 9 13 10 9 2
25 11 4 0 3 13 0 9 1 14 13 10 9 1 11 1 16 15 1 13 9 1 9 1 9 2
40 12 9 1 11 13 9 1 10 9 2 7 1 9 1 9 1 0 9 7 14 13 9 10 9 1 9 2 13 15 10 9 1 16 9 1 0 9 4 13 2
27 0 9 1 9 7 9 1 0 9 1 9 2 13 10 0 9 1 14 4 13 14 13 9 1 10 9 2
31 9 1 9 13 3 3 0 1 11 15 0 9 1 9 13 1 11 2 7 10 9 13 3 0 9 1 9 7 0 9 2
26 9 13 0 9 1 0 9 1 0 9 1 9 2 9 7 10 9 15 13 9 1 16 9 13 9 2
16 9 1 9 1 10 0 7 0 9 1 11 1 11 13 3 2
21 3 4 15 2 11 2 13 0 1 10 9 16 11 13 1 2 7 13 3 0 2
37 11 13 0 1 0 1 11 1 9 2 7 13 1 10 9 16 11 7 4 13 1 3 12 9 2 7 16 15 13 1 12 9 3 0 1 9 2
39 3 4 13 3 0 11 13 1 9 3 1 11 2 7 1 14 13 1 1 0 9 2 7 16 10 9 13 10 9 3 3 1 11 2 7 1 0 9 2
30 16 11 4 13 14 13 10 0 0 9 1 11 1 9 1 11 3 3 9 13 10 9 1 9 2 13 9 10 9 2
24 11 4 3 3 13 0 9 1 10 9 1 9 1 10 0 9 7 1 9 2 9 7 9 2
15 1 0 9 1 10 9 4 15 13 1 10 9 1 9 2
4 10 0 9 5
14 15 13 0 7 0 16 15 13 0 0 1 0 9 2
16 7 10 1 10 0 0 9 1 11 13 10 9 1 12 9 2
19 15 13 3 10 9 1 11 2 0 1 9 11 2 7 13 15 10 9 2
7 10 0 13 11 11 1 2
7 11 13 12 9 7 9 2
11 9 10 13 9 1 11 1 12 1 12 2
18 3 4 11 13 0 0 9 7 13 0 1 10 9 1 9 1 9 2
11 1 10 9 3 13 15 3 9 1 11 2
11 3 13 15 9 1 9 15 13 10 9 2
25 11 11 11 11 13 11 0 9 2 13 1 11 2 7 4 1 0 9 13 1 15 7 10 9 2
24 3 13 15 1 10 9 1 9 2 10 0 9 1 9 16 15 13 10 0 1 10 0 9 2
9 15 4 13 16 9 1 11 13 2
23 0 4 4 13 7 13 1 10 0 9 1 0 9 2 0 1 11 11 1 11 0 9 2
39 15 13 3 16 15 15 13 13 0 2 7 11 13 1 10 9 10 9 1 16 10 9 4 13 0 9 7 9 3 1 10 9 16 9 13 1 0 9 2
13 14 13 1 1 11 1 9 1 0 9 13 0 2
25 0 9 4 15 13 1 9 15 4 13 15 16 15 13 0 7 15 13 1 11 9 1 11 9 2
17 9 15 13 9 1 9 1 9 4 13 7 13 0 9 1 9 2
11 15 13 0 0 14 13 1 0 0 9 2
13 0 1 11 4 3 13 9 7 13 0 0 9 2
25 3 16 11 0 4 13 10 9 1 11 1 12 2 13 9 1 9 1 10 0 7 3 0 9 2
19 9 9 13 3 0 1 9 0 9 2 16 10 0 11 0 13 0 9 2
21 1 11 13 9 14 4 13 1 10 0 9 2 15 1 15 13 1 9 0 1 2
29 16 9 3 13 1 11 2 4 15 13 16 10 0 9 13 0 2 7 0 13 9 2 9 15 13 15 1 9 2
18 10 0 13 16 3 10 9 0 13 13 3 1 9 15 13 0 0 2
10 15 4 3 3 13 9 1 0 9 2
10 3 4 15 13 9 15 3 13 0 2
5 15 13 3 9 2
12 7 3 1 11 13 9 2 1 9 1 11 2
15 16 15 13 9 16 15 3 13 15 1 2 13 15 3 2
13 11 13 0 0 0 7 0 16 15 4 13 15 2
22 9 13 0 0 9 2 15 15 13 4 13 1 9 1 9 15 13 1 14 13 1 2
7 7 9 13 0 3 0 2
8 15 13 9 2 9 7 9 2
4 9 13 0 2
16 13 15 10 9 1 10 0 9 2 13 15 3 9 1 9 2
8 3 10 12 9 13 1 11 2
13 4 15 13 9 1 9 2 13 11 11 12 9 2
18 3 4 15 13 1 9 1 0 0 9 1 0 9 2 9 7 9 2
5 7 1 13 15 2
7 1 12 0 9 2 11 2
4 9 13 1 5
2 9 5
4 0 7 0 5
4 0 7 0 5
2 9 5
16 3 10 0 9 1 9 2 9 2 13 0 13 1 1 11 2
3 0 9 2
15 11 1 12 4 13 10 9 16 9 13 10 3 0 9 2
10 9 13 10 10 9 1 9 7 9 2
15 9 13 3 0 1 1 9 2 1 15 15 4 13 1 2
21 1 13 15 10 9 2 0 0 15 15 4 13 1 9 1 9 1 9 7 9 2
28 10 0 9 13 9 1 10 9 2 15 15 13 1 9 2 9 2 9 1 10 10 2 9 1 9 7 9 2
14 15 13 15 3 1 0 9 15 3 13 1 0 9 2
15 7 3 16 10 0 9 13 2 13 9 0 1 10 9 2
12 9 1 9 13 0 0 2 13 0 9 9 2
36 9 13 15 1 1 9 1 14 13 9 13 1 9 7 9 2 15 13 0 2 15 13 3 0 1 10 9 7 13 0 1 9 1 10 9 2
24 0 9 13 15 10 10 0 9 1 2 7 15 14 13 3 15 13 1 10 9 13 10 9 2
22 15 13 9 0 13 13 14 13 1 10 9 1 15 15 13 1 9 7 9 14 13 2
4 9 13 15 2
16 16 0 9 3 13 2 0 2 2 13 15 0 9 1 15 2
29 2 9 2 1 9 13 14 13 15 10 7 3 15 4 13 2 1 14 13 0 9 2 1 11 1 1 9 11 2
12 13 9 10 9 15 13 1 9 1 9 3 2
15 7 13 15 10 9 15 4 13 15 1 15 15 13 9 2
13 1 9 13 9 1 9 3 0 1 9 7 9 2
19 15 4 13 15 0 14 4 13 15 15 13 0 7 0 1 0 7 0 2
15 15 13 15 15 4 13 16 11 13 1 0 9 1 9 2
10 2 9 2 4 15 3 13 15 1 2
27 3 9 13 9 1 9 2 7 3 16 2 15 2 13 9 2 4 15 13 10 0 9 1 2 9 2 2
8 7 13 9 9 3 11 13 2
22 15 4 13 16 9 13 9 2 7 4 3 13 9 16 15 13 15 2 10 10 10 2
27 10 9 1 16 2 11 13 9 2 4 3 4 13 1 15 15 13 16 2 9 2 3 13 10 0 9 2
28 16 15 13 15 9 2 9 2 15 15 13 1 11 7 9 9 2 13 15 0 1 15 15 3 4 13 15 2
33 15 13 9 1 0 9 1 9 7 9 2 15 13 0 9 7 0 9 2 7 15 4 13 15 9 13 1 1 1 14 13 9 2
16 13 15 1 1 9 11 9 2 13 15 10 9 1 0 9 2
9 10 0 9 13 1 9 7 9 2
23 9 4 13 0 2 7 3 0 13 2 1 14 13 1 1 9 2 15 15 3 0 13 2
12 10 0 9 1 9 7 9 13 15 12 9 2
35 10 12 13 16 9 4 13 0 7 9 1 14 13 10 0 9 3 2 10 10 13 16 9 15 13 1 10 9 13 10 10 1 10 9 2
28 15 4 1 9 13 9 16 15 13 15 3 15 4 13 9 15 13 2 9 2 2 10 9 7 9 1 9 2
30 15 4 13 9 0 9 16 15 4 13 11 1 9 1 9 7 15 4 13 11 16 15 13 0 1 7 9 7 9 2
36 7 1 9 11 13 15 9 1 15 4 13 0 0 1 15 15 13 15 1 9 2 7 15 13 10 9 1 16 9 9 13 0 7 3 0 2
14 3 10 0 9 1 9 2 9 2 13 0 13 1 2
7 10 9 13 0 1 10 5
3 0 9 2
7 13 15 15 13 9 1 2
5 9 2 3 9 2
2 9 2
21 11 11 11 4 1 9 4 13 16 15 13 9 7 9 1 11 1 10 0 9 2
2 9 2
21 0 13 11 11 7 11 11 16 15 13 10 9 1 11 3 9 13 0 3 0 2
15 10 12 4 13 10 9 15 3 11 7 11 4 13 1 2
24 10 12 0 9 13 16 11 9 2 1 9 1 11 7 11 2 13 0 9 1 9 1 11 2
17 16 10 12 9 13 1 0 16 15 7 13 9 7 9 1 11 2
32 9 13 10 0 9 1 0 9 1 9 1 9 7 9 2 7 0 9 1 9 1 0 0 9 7 0 0 9 1 9 9 2
25 11 13 10 9 0 1 10 0 0 9 2 0 15 9 13 0 9 1 9 7 9 1 9 13 2
18 7 9 13 3 10 9 1 9 1 15 1 15 15 13 15 4 13 2
16 7 9 2 11 11 9 7 9 4 13 0 9 1 10 9 2
12 16 11 4 4 13 2 4 11 7 11 13 2
15 9 11 11 4 13 0 9 0 1 14 13 11 9 1 2
27 9 4 13 2 3 16 15 13 0 9 1 14 13 1 9 2 7 16 9 1 0 9 1 9 13 0 2
13 10 0 4 13 9 1 11 9 1 10 0 9 2
32 15 13 1 14 13 0 9 1 11 1 10 0 9 15 13 1 2 1 1 15 15 0 4 13 1 0 9 1 10 0 9 2
16 3 16 10 0 9 3 13 10 9 2 13 10 0 9 0 2
9 9 1 1 2 9 13 15 3 2
9 10 0 9 4 3 13 1 9 2
10 16 9 11 11 1 10 0 9 13 2
15 2 15 13 10 9 1 9 2 1 15 13 15 9 2 2
15 10 9 1 3 0 9 13 3 0 16 15 13 1 9 2
23 7 9 4 3 3 13 1 2 15 4 3 13 2 7 3 4 15 3 13 9 1 9 2
24 10 0 0 9 13 9 1 0 9 16 10 9 1 9 3 4 13 15 3 3 9 13 0 2
15 15 13 1 0 9 9 2 3 13 7 4 15 13 0 2
18 0 9 4 1 9 3 13 2 3 4 15 0 13 1 10 0 9 2
23 0 3 13 11 0 9 2 0 9 4 3 0 13 16 15 0 13 1 14 13 0 9 2
20 9 7 9 13 3 0 0 2 7 4 3 0 0 13 1 10 0 0 9 2
17 9 4 3 13 3 2 15 13 15 3 0 1 9 1 12 9 2
14 1 10 9 13 9 1 9 0 2 3 1 0 9 2
21 1 9 13 9 9 0 1 10 9 2 16 1 9 13 10 9 3 0 1 9 2
29 9 1 9 7 9 1 11 1 9 13 0 1 10 0 0 9 2 7 13 1 9 0 1 10 9 1 0 9 2
14 1 9 4 10 0 9 13 0 1 9 1 10 9 2
28 15 4 13 1 9 1 9 2 13 9 1 10 9 1 9 1 0 2 3 0 9 2 7 13 0 1 9 2
8 0 9 1 0 9 1 9 2
45 1 9 13 15 3 15 15 3 4 13 2 15 13 1 9 2 1 12 9 9 14 1 9 2 12 9 9 1 9 7 10 9 1 12 9 13 10 12 0 16 9 13 1 9 2
9 9 4 13 16 9 13 0 9 2
33 1 9 1 9 1 9 1 9 7 9 4 9 1 9 1 0 9 13 2 0 15 15 13 1 9 1 9 2 7 1 15 9 2
22 0 9 1 9 1 9 1 14 13 9 7 9 3 9 1 0 9 13 1 12 9 2
32 1 9 13 10 9 9 1 12 9 9 1 9 16 15 13 14 13 2 16 9 13 0 1 9 1 9 16 15 13 1 9 2
20 15 13 3 3 10 0 9 2 7 13 3 10 9 1 9 1 0 0 9 2
11 13 9 9 1 14 13 10 9 1 9 2
15 1 9 13 9 1 9 7 9 0 2 16 9 13 0 2
17 15 4 3 13 10 9 15 13 16 9 4 13 1 10 9 0 2
14 10 0 13 9 11 1 0 12 9 9 1 0 9 2
29 10 10 9 4 1 10 9 13 1 16 10 0 9 13 15 15 13 9 2 16 15 3 3 13 14 13 15 0 2
6 9 15 4 13 1 5
4 4 3 13 2
2 9 2
4 9 1 9 2
21 9 13 1 14 13 0 1 16 15 13 0 16 0 13 1 9 1 11 0 9 2
11 7 9 4 13 16 9 13 9 1 9 2
23 15 15 4 13 9 7 9 7 9 1 11 0 9 4 13 15 1 11 7 10 0 9 2
13 16 15 13 0 13 10 10 9 15 4 13 3 2
30 7 1 14 4 13 1 1 10 9 2 10 9 7 2 1 0 9 2 9 2 13 10 0 9 1 9 1 9 9 2
13 15 13 3 14 4 13 7 9 1 11 0 9 2
12 1 0 13 15 1 12 9 1 9 1 11 2
22 10 9 1 12 13 16 3 12 9 1 11 9 13 16 11 11 13 1 1 10 0 2
11 10 9 13 0 2 16 12 9 13 9 2
18 15 13 16 9 1 9 1 11 0 9 13 7 13 0 1 10 9 2
28 7 10 15 15 3 13 1 9 13 0 1 14 13 9 1 9 2 7 3 13 10 0 9 1 11 0 9 2
11 15 15 13 2 13 10 0 9 1 9 2
22 9 1 11 11 1 11 11 7 11 11 1 9 1 9 13 1 10 1 9 1 9 2
25 9 13 1 16 9 13 15 1 1 9 2 7 13 9 2 3 16 15 3 13 15 11 13 1 2
18 15 13 0 9 1 10 9 2 1 11 0 9 2 7 10 0 9 2
7 0 13 15 10 0 9 2
11 7 9 7 9 13 10 0 7 0 9 2
12 11 13 1 9 10 9 15 13 0 7 0 2
14 7 15 15 13 11 13 10 9 1 15 15 13 11 2
8 1 11 0 9 13 15 0 2
22 3 4 1 7 1 15 15 13 14 13 9 13 10 9 0 2 3 0 0 13 9 2
13 7 15 4 13 1 9 2 3 3 1 0 9 2
24 1 0 11 13 11 11 1 9 1 16 11 8 3 13 1 9 1 14 13 15 1 1 9 2
15 2 15 13 0 1 14 13 9 1 10 2 15 13 9 2
9 9 13 16 11 8 3 13 15 2
22 13 15 16 15 13 0 2 10 9 15 0 13 1 14 13 3 0 10 9 13 2 2
30 9 1 11 0 9 4 13 2 7 4 0 13 2 16 15 3 7 0 13 15 15 13 1 10 0 9 15 13 15 2
15 3 4 15 3 13 1 3 0 9 1 9 1 10 0 2
19 15 4 3 3 13 10 9 1 15 15 1 9 1 9 4 13 1 9 2
11 1 9 4 9 0 13 9 1 10 9 2
7 7 9 4 3 13 0 2
29 0 9 1 9 4 1 9 13 1 10 9 15 13 16 0 9 13 0 3 0 9 1 9 1 9 1 0 9 2
27 0 1 15 4 13 1 16 9 2 0 1 10 0 9 1 0 9 2 13 10 0 9 1 10 0 9 2
12 7 3 0 0 13 15 16 9 13 9 9 2
6 0 2 7 0 0 5
3 9 3 5
2 9 5
11 13 1 13 9 7 9 15 1 3 0 2
5 15 13 10 9 2
14 13 1 13 15 3 0 0 2 7 9 13 3 0 2
14 1 9 1 11 11 11 4 15 13 1 0 0 9 2
18 1 10 1 10 3 0 13 9 1 10 0 9 9 1 11 9 1 2
12 9 13 16 9 9 4 13 1 12 1 10 2
15 1 0 9 13 15 0 9 1 16 10 0 9 13 12 2
8 15 13 9 1 10 0 9 2
29 1 9 1 9 13 0 9 1 1 15 7 13 16 15 1 11 0 13 0 9 1 9 15 9 4 13 1 1 2
8 15 4 13 16 15 3 13 2
27 15 13 0 14 13 1 9 15 13 1 9 1 9 2 7 9 13 0 13 0 7 0 0 1 15 9 2
9 15 13 3 0 0 0 7 0 2
15 9 13 0 0 7 0 1 14 13 9 7 9 0 0 2
8 9 13 0 10 0 0 9 2
21 16 12 9 13 2 13 15 3 1 9 2 3 0 1 3 1 9 15 13 1 2
22 12 9 4 3 3 13 1 9 3 2 7 4 3 3 13 1 15 10 10 13 1 2
11 15 13 3 3 0 1 10 0 0 11 2
12 14 13 9 13 0 10 0 1 15 1 9 2
22 15 13 3 0 1 15 13 3 0 1 10 9 15 4 13 3 1 14 13 1 9 2
30 10 0 0 9 13 11 11 1 11 11 11 1 9 1 11 1 12 1 16 15 4 13 1 7 2 13 2 10 9 2
6 15 13 15 3 0 2
5 15 13 3 3 2
11 1 11 13 9 14 13 7 15 13 15 2
32 3 16 10 0 9 13 0 9 2 15 15 13 1 7 9 7 9 2 4 10 9 3 4 13 2 1 16 15 13 0 9 2
23 15 13 1 9 0 0 16 15 4 13 3 0 15 15 13 2 16 10 9 13 3 0 2
8 1 11 13 0 10 0 9 2
18 1 11 13 15 3 0 9 2 7 10 0 15 13 4 13 1 12 2
18 11 13 10 3 0 9 16 15 10 9 4 13 10 9 1 0 9 2
7 1 11 13 9 0 0 2
13 15 13 3 10 9 7 9 15 4 13 0 0 2
12 1 11 4 10 0 9 13 1 0 7 9 2
15 11 13 1 9 0 7 9 7 9 13 10 0 0 9 2
13 1 11 4 15 3 13 1 9 1 9 7 9 2
8 3 0 13 15 3 1 11 2
11 0 9 13 1 0 0 1 10 0 9 2
12 1 10 0 0 7 0 9 13 15 0 0 2
16 15 13 3 10 0 9 2 0 9 13 3 1 10 0 9 2
11 15 13 15 15 15 13 1 11 7 11 2
31 9 13 10 0 9 1 16 15 13 15 0 1 11 2 3 3 3 0 16 15 13 10 9 3 0 1 11 7 11 3 2
20 9 4 13 1 10 9 15 1 10 0 9 4 13 1 1 10 0 0 9 2
13 15 13 3 3 3 0 2 3 1 9 7 9 2
7 4 11 7 11 13 9 2
3 3 12 2
23 0 0 13 1 16 15 3 13 11 7 11 15 4 13 9 2 7 11 2 11 7 11 2
16 9 1 10 12 13 0 0 2 7 15 4 3 13 9 3 2
34 16 11 11 13 1 9 1 11 0 1 9 2 13 15 0 1 10 9 15 4 13 3 0 1 10 0 9 2 9 2 11 7 11 2
19 2 10 9 4 3 4 13 10 0 0 9 2 10 0 9 7 9 2 2
19 0 0 4 15 3 13 16 3 4 11 13 15 1 9 2 9 7 9 2
8 10 9 4 15 3 13 13 2
9 7 1 10 10 9 13 11 0 2
9 9 10 4 0 13 1 10 9 2
16 10 0 9 13 14 13 1 11 1 10 9 1 0 9 9 2
20 3 13 11 9 1 9 0 2 16 9 13 1 11 0 7 0 0 0 9 2
23 3 13 15 0 9 1 11 1 9 2 7 10 0 9 13 15 3 3 0 1 10 9 2
35 0 13 15 0 9 1 10 9 1 11 2 7 15 4 13 0 16 15 3 0 13 10 0 9 1 16 11 3 13 1 10 3 0 9 2
11 11 7 11 4 13 3 1 10 0 9 2
12 10 0 9 4 4 13 1 10 0 0 9 2
16 1 12 13 10 0 9 1 11 3 12 9 1 11 3 9 2
17 11 2 3 9 0 9 2 13 10 0 9 1 10 9 1 11 2
19 10 9 4 1 0 9 13 1 14 13 10 0 9 11 13 1 10 9 2
9 0 9 13 3 10 0 0 9 2
23 10 0 0 7 0 9 1 11 13 10 0 9 1 9 1 10 0 9 1 12 2 12 2
13 0 4 13 1 3 9 4 13 1 10 0 9 2
17 1 9 13 10 0 9 0 0 2 9 1 11 13 10 12 0 2
20 16 9 3 13 1 11 2 13 3 9 1 10 0 0 0 9 10 0 9 2
30 0 13 15 3 16 11 3 4 13 3 0 1 10 0 9 7 1 9 2 16 10 9 1 11 3 4 13 11 0 2
15 10 0 9 1 10 0 9 1 0 9 2 13 3 0 2
26 3 4 9 13 14 13 1 0 9 1 16 9 3 0 4 13 10 0 9 15 4 13 1 0 9 2
14 10 0 9 13 3 1 9 1 14 13 10 0 9 2
22 15 13 0 1 10 9 16 9 4 13 9 1 9 1 3 15 4 13 1 0 9 2
9 3 4 11 13 15 0 1 11 2
16 4 11 0 13 10 0 9 2 4 10 0 9 3 13 0 2
19 15 4 13 16 15 13 1 9 7 16 9 4 13 10 0 9 1 9 2
9 0 9 4 3 13 1 1 9 2
14 0 13 1 16 11 13 0 1 14 13 10 10 9 2
7 15 13 10 9 1 9 2
11 11 13 0 0 2 7 9 4 0 13 2
13 9 13 3 3 0 1 16 12 9 3 4 13 2
4 11 1 9 5
3 13 3 2
2 9 2
4 10 0 9 2
2 0 2
5 1 9 1 9 2
3 11 13 2
3 0 9 2
10 0 9 4 9 9 4 13 1 11 2
29 12 9 1 9 1 9 13 9 14 13 10 0 2 0 7 0 9 15 13 15 10 1 10 0 9 1 10 9 2
22 3 13 15 1 16 3 1 10 0 0 9 9 2 4 15 13 9 15 13 10 9 2
26 10 0 9 1 14 13 0 2 7 1 9 2 4 4 13 1 10 9 2 7 13 1 9 10 9 2
25 11 4 13 0 1 9 2 10 0 9 13 11 2 16 11 4 4 13 1 0 9 1 10 9 2
14 15 13 10 0 1 15 9 13 3 0 1 1 9 2
9 9 11 11 13 0 10 0 9 2
7 9 13 0 1 10 9 2
9 9 9 4 3 13 9 1 9 2
16 11 9 13 1 9 10 9 1 12 9 9 1 9 1 12 2
7 7 15 13 9 1 11 2
18 3 4 9 11 11 13 1 10 9 15 3 13 9 1 14 13 9 2
21 11 4 13 1 10 0 9 1 9 2 7 9 4 13 15 1 1 9 1 9 2
14 15 13 3 3 3 1 14 13 9 1 14 4 13 2
15 11 4 0 1 10 9 13 10 0 9 16 15 13 3 2
8 7 12 0 9 13 1 9 2
11 15 13 3 0 1 14 13 9 1 9 2
19 10 9 4 3 13 1 9 16 9 4 13 1 9 2 7 3 0 3 2
17 9 4 13 10 9 1 16 11 13 10 0 9 15 11 4 13 2
21 1 10 9 1 9 4 9 13 14 13 9 1 0 9 15 3 13 0 0 9 2
10 16 9 4 13 2 4 9 13 1 2
15 15 4 13 10 9 2 7 1 10 9 4 9 13 9 2
17 11 4 13 15 2 7 0 3 0 1 14 13 0 9 1 11 2
14 1 11 13 11 11 1 9 15 3 4 13 1 11 2
7 11 4 3 13 10 9 2
18 15 13 3 1 11 1 0 9 2 16 15 3 1 10 0 13 13 2
27 10 9 1 14 13 3 1 0 9 1 10 9 2 1 11 9 1 9 1 9 12 2 13 3 3 0 2
26 1 11 13 15 10 0 9 2 7 3 4 11 3 10 9 13 10 0 2 0 9 10 9 1 9 2
19 11 4 3 13 10 0 9 1 14 4 13 11 1 9 0 9 1 9 2
20 3 16 15 13 10 9 1 9 1 12 9 1 11 12 2 13 15 3 0 2
16 9 4 13 14 13 9 1 9 1 0 9 2 9 7 9 2
16 1 0 9 4 9 13 9 2 13 10 9 7 13 10 9 2
9 10 15 1 9 1 10 0 9 2
19 9 13 3 3 0 2 9 4 3 13 2 7 1 11 13 9 9 9 2
9 0 9 4 13 1 9 7 9 2
33 0 9 4 13 1 12 9 1 0 9 1 12 1 12 9 1 12 2 9 4 13 10 10 12 9 7 9 13 1 11 11 13 2
12 3 1 9 13 11 9 0 1 14 13 9 2
26 15 13 3 0 9 1 10 9 15 1 9 13 10 9 1 12 9 2 7 3 9 13 10 0 9 2
13 3 13 9 0 0 1 16 11 13 10 0 9 2
43 15 13 10 0 0 16 10 0 0 9 1 11 2 9 1 9 13 10 9 1 11 2 13 0 9 1 14 13 1 0 9 2 7 13 9 16 15 4 13 1 10 9 2
8 10 0 9 4 3 13 9 2
16 0 13 16 9 11 11 7 10 9 0 13 3 0 1 9 2
15 15 13 15 1 0 1 0 9 1 10 0 7 0 9 2
29 10 0 9 13 16 1 11 13 15 1 9 2 16 10 0 9 3 4 13 9 2 15 0 13 0 9 1 15 2
14 15 4 13 0 14 13 9 1 11 0 9 1 12 2
21 15 15 3 13 1 1 14 13 9 2 4 0 13 1 1 9 16 9 9 13 2
10 7 3 3 1 9 4 11 13 9 2
15 1 9 9 4 15 13 0 9 1 9 1 10 0 9 2
29 9 13 0 7 0 2 1 12 4 9 13 1 12 9 2 9 1 1 12 9 7 12 9 1 9 4 13 0 2
19 1 0 9 10 9 4 10 9 13 10 10 9 1 14 13 10 0 9 2
11 11 4 3 3 13 16 15 4 13 9 2
14 10 9 4 13 15 10 16 11 10 13 9 1 9 2
35 0 4 15 1 14 13 9 1 15 2 7 14 13 1 16 10 9 7 9 13 1 10 9 2 13 1 1 14 13 14 13 10 0 9 2
11 3 9 11 4 13 9 1 9 1 11 2
14 1 9 13 15 10 9 16 10 0 9 13 1 9 2
19 16 11 9 3 4 13 9 2 4 15 13 10 0 9 1 0 0 9 2
17 11 2 3 7 9 7 0 9 13 2 13 1 10 3 0 9 2
20 13 15 13 15 4 13 3 0 7 0 1 9 15 15 3 4 13 1 9 2
6 11 4 13 0 9 5
5 13 15 1 11 2
16 9 1 0 9 1 9 1 11 4 13 10 9 1 0 9 2
38 16 10 0 9 13 14 13 15 1 2 0 9 2 1 10 0 2 9 2 2 13 0 9 14 13 0 1 1 9 1 14 13 0 9 1 0 9 2
28 1 11 13 15 2 2 2 1 0 9 2 2 15 13 16 15 13 9 1 11 2 7 15 13 15 3 2 2
8 15 15 4 13 2 13 3 2
7 15 13 0 9 1 9 2
15 9 2 9 2 13 10 2 0 9 2 1 0 0 9 2
31 15 13 3 16 15 13 10 0 9 15 3 13 1 9 2 9 7 9 2 0 11 2 11 2 2 7 3 3 3 11 2
30 9 13 3 3 16 15 4 13 9 1 11 1 10 9 1 10 0 9 2 7 16 15 13 13 9 1 10 0 9 2
36 15 13 0 0 2 16 10 9 15 13 9 1 15 15 13 1 1 10 0 9 2 13 0 0 1 9 15 4 13 1 7 13 9 1 9 2
14 9 1 0 9 1 9 4 13 10 9 1 0 9 2
16 0 0 9 13 0 1 3 15 15 13 2 3 13 7 13 2
14 10 9 7 10 9 15 3 13 0 2 4 13 0 2
5 15 13 11 9 2
32 7 9 1 16 11 4 13 0 9 2 13 0 3 0 7 1 9 1 9 2 15 15 4 13 1 9 1 9 9 1 9 2
14 9 1 9 1 9 13 3 16 15 4 13 1 9 2
5 15 13 1 9 2
32 14 13 13 3 14 13 9 7 14 13 10 9 2 7 14 13 0 2 3 16 15 4 13 1 9 1 0 9 1 10 9 2
10 10 2 15 2 4 13 0 9 1 2
29 15 15 13 1 10 0 0 9 2 4 13 1 10 11 2 7 15 4 13 1 9 1 14 13 2 13 9 11 2
9 3 13 15 3 0 1 10 9 2
17 15 13 0 16 9 4 13 0 9 7 13 0 0 1 14 13 2
15 15 13 0 9 15 13 0 9 16 15 13 9 1 9 2
8 7 13 3 10 9 3 0 2
8 15 13 15 3 15 15 13 2
13 10 0 9 2 9 11 2 13 10 0 9 0 2
14 13 9 11 2 13 15 0 9 7 13 0 9 0 2
11 16 15 13 0 2 13 3 9 3 0 2
23 3 13 3 10 9 3 0 2 0 1 10 9 1 11 2 15 13 0 10 9 1 9 2
22 7 16 15 13 16 11 0 13 10 0 9 1 9 1 9 2 13 3 9 3 0 2
8 15 13 3 3 1 10 9 2
26 16 15 13 10 0 2 13 15 10 9 1 14 13 9 1 3 15 4 13 10 9 1 10 3 0 2
18 7 16 9 13 9 2 3 13 3 0 9 0 0 1 16 9 13 2
21 15 13 3 1 10 9 7 9 1 9 2 7 1 0 9 7 1 9 1 9 2
9 11 9 2 15 0 1 15 10 5
3 13 3 2
4 9 13 1 2
28 16 0 0 4 13 0 7 0 0 1 14 13 9 1 9 2 13 11 9 3 0 1 16 15 3 13 9 2
10 15 4 13 10 9 9 1 11 9 2
14 10 0 4 13 15 1 9 9 2 7 13 0 0 2
14 10 0 0 9 11 9 13 10 0 7 0 0 9 2
13 1 9 13 12 0 9 9 1 10 9 0 9 2
5 0 13 0 0 2
18 1 10 13 15 0 14 13 9 1 10 9 9 4 13 1 10 9 2
20 1 10 9 13 9 1 9 1 11 9 16 15 13 9 7 13 14 13 9 2
26 9 1 9 4 3 13 1 0 9 2 7 9 13 0 9 1 0 9 1 3 15 4 13 11 9 2
14 1 10 0 13 13 9 0 9 1 14 13 9 9 2
17 1 10 0 13 11 9 15 0 1 10 0 16 15 3 13 9 2
11 1 9 7 9 13 15 9 10 0 9 2
16 9 9 13 16 11 13 9 2 7 3 3 9 1 11 9 2
16 7 10 0 9 1 11 9 7 10 9 13 1 9 1 11 2
17 10 3 0 9 13 3 1 14 13 16 11 7 13 11 7 9 2
38 10 0 9 1 11 1 12 2 15 7 13 16 9 13 9 2 2 2 7 13 10 9 0 9 2 13 16 11 11 13 2 1 10 9 1 11 2 2
11 15 13 7 9 7 9 2 0 7 9 2
5 11 9 13 0 2
12 15 13 9 7 13 10 10 0 13 1 9 2
14 9 13 11 1 11 9 2 7 13 16 15 13 0 2
12 3 13 4 15 3 13 16 9 13 0 0 2
25 7 11 11 2 1 11 9 2 7 9 0 9 4 13 1 16 11 3 13 10 10 1 10 9 2
10 7 11 9 13 10 9 1 10 9 2
20 15 13 1 1 10 9 10 0 13 2 3 16 15 3 4 13 10 10 9 2
26 11 11 13 3 16 10 0 0 2 7 3 11 0 9 2 13 11 0 0 16 15 10 13 9 1 2
14 0 13 16 11 9 13 10 0 0 9 1 9 12 2
18 1 9 13 15 16 11 3 13 1 0 7 2 10 0 9 2 13 2
20 15 13 0 16 9 1 9 13 3 9 9 13 1 11 11 7 13 9 12 2
8 7 3 12 13 10 0 9 2
13 9 9 13 3 1 16 10 0 9 3 4 13 2
19 9 15 4 13 2 13 0 2 15 15 3 4 13 1 9 1 11 9 2
17 0 1 12 13 9 2 0 1 9 1 16 9 13 10 0 9 2
10 7 1 10 9 4 11 9 13 0 2
17 1 11 13 15 1 0 3 0 9 3 1 1 12 2 1 12 2
16 15 13 10 0 0 9 7 13 0 7 10 9 1 10 0 2
5 11 13 1 9 5
4 9 1 11 2
3 0 9 2
15 11 13 0 0 9 1 9 7 1 9 1 9 7 9 2
11 7 14 13 9 9 3 1 9 13 0 2
20 1 12 13 9 1 10 0 9 11 11 9 1 9 1 9 11 11 9 1 2
14 1 12 9 9 13 11 15 0 0 11 9 1 9 2
27 10 9 13 10 1 0 9 1 16 11 13 9 1 14 13 10 0 0 9 15 3 13 0 1 0 9 2
30 1 9 11 11 11 2 9 1 11 1 11 2 4 11 1 12 3 0 13 1 9 1 14 13 10 9 7 11 9 2
17 9 13 10 9 1 9 1 12 2 9 9 1 7 9 1 11 2
10 11 4 3 13 9 16 15 13 9 2
19 10 9 4 13 10 0 9 1 11 9 7 4 13 1 9 12 0 9 2
19 7 9 4 13 0 1 1 11 2 1 9 11 11 2 0 13 11 11 2
15 1 12 13 3 9 14 13 9 7 13 1 0 0 9 2
24 10 0 9 11 11 1 11 9 4 1 9 13 16 11 0 4 13 9 1 0 9 1 11 2
22 10 10 9 16 10 0 9 0 13 9 1 9 2 13 9 9 2 15 3 13 0 2
8 11 4 13 9 9 1 9 2
20 1 10 0 9 11 11 4 15 13 10 9 1 9 1 14 13 10 0 9 2
30 11 3 0 9 2 11 11 2 13 16 10 0 9 15 13 11 1 9 1 9 1 9 12 2 13 10 9 1 15 2
38 10 0 1 11 9 13 16 9 1 11 4 13 1 0 9 10 0 9 16 10 0 9 2 1 11 1 9 2 13 9 1 11 3 1 9 1 12 2
25 9 13 1 9 1 11 7 11 7 4 1 9 13 1 14 13 10 0 9 1 16 11 13 11 2
17 11 13 16 11 0 9 4 13 10 0 1 11 7 13 10 0 2
15 10 0 9 1 11 4 13 10 0 9 0 9 1 9 2
5 9 4 3 13 2
32 3 4 9 11 11 11 7 10 0 0 9 11 11 13 1 16 15 13 16 7 11 7 9 13 9 1 14 13 11 1 9 2
20 7 11 13 10 9 2 3 3 10 0 9 2 7 4 3 3 13 1 9 2
33 10 0 11 4 1 9 13 9 2 9 7 9 1 0 2 7 13 1 10 0 9 11 8 11 11 12 9 1 9 1 0 9 2
10 9 13 0 1 10 0 2 0 11 2
21 9 11 11 4 1 11 11 2 9 1 11 9 1 9 2 13 10 9 1 9 2
9 15 13 16 15 10 13 1 11 5
3 0 9 2
14 15 13 3 0 1 11 2 11 11 2 11 7 11 2
11 15 13 3 10 0 9 15 13 1 11 2
16 1 9 13 15 10 10 0 9 1 11 9 1 9 1 11 2
17 1 10 10 9 4 12 9 0 0 13 1 11 1 9 1 11 2
35 10 9 13 9 1 10 0 9 1 9 1 11 2 11 7 11 11 7 10 0 2 11 11 2 15 13 1 9 1 10 0 9 1 0 2
12 15 4 13 0 9 1 9 1 10 0 9 2
15 10 0 9 4 10 9 7 9 13 1 7 1 0 11 2
27 3 13 10 0 9 14 13 16 11 11 9 0 13 9 1 10 0 9 15 4 13 1 0 9 1 12 2
18 0 13 10 0 9 0 1 0 9 1 0 9 1 10 3 0 9 2
27 1 11 2 1 1 11 11 2 13 0 9 14 13 9 15 4 13 0 9 2 7 15 3 13 0 9 2
7 10 9 13 9 0 9 2
13 10 9 13 15 14 13 0 9 7 10 9 1 2
6 7 3 13 3 9 2
16 10 9 1 9 1 11 7 1 10 9 1 11 13 0 9 2
15 0 9 15 13 1 0 7 0 9 1 11 11 13 3 2
36 10 0 9 13 15 0 9 1 3 0 9 2 1 9 1 10 9 7 10 9 2 13 9 1 1 10 11 9 13 1 9 2 9 7 9 2
21 10 9 4 10 0 9 2 0 11 11 2 13 1 11 1 10 0 9 1 11 2
15 7 11 2 15 13 11 11 2 7 9 11 13 9 0 2
17 7 1 10 9 1 9 2 1 9 7 1 9 4 15 3 13 2
19 10 0 9 13 15 10 0 9 1 10 0 7 0 9 1 9 1 11 2
31 10 9 13 0 9 15 1 1 11 9 1 10 0 9 1 14 13 10 0 9 15 3 3 13 1 9 1 9 7 9 2
17 1 9 13 15 1 1 0 0 9 7 10 9 1 9 7 9 2
18 12 0 4 0 13 1 11 16 11 1 11 9 13 9 0 1 12 2
19 15 13 1 9 9 1 9 2 1 9 2 1 0 9 2 7 1 9 2
6 9 4 13 0 0 2
17 16 15 10 13 1 11 7 11 11 4 9 13 10 9 1 11 2
22 15 13 0 16 0 9 13 0 9 1 10 0 9 1 9 1 12 7 9 1 12 2
15 9 13 1 1 9 16 15 13 1 15 15 13 1 11 2
35 9 1 9 2 9 7 11 9 1 0 13 16 0 9 4 13 2 1 9 2 10 0 9 1 9 15 13 9 1 15 10 7 10 9 2
10 7 2 10 0 9 13 3 10 9 2
5 16 9 13 9 5
2 9 2
2 9 2
4 10 0 0 2
4 11 11 11 2
2 9 2
7 11 11 13 10 0 9 2
25 7 4 15 4 13 1 10 10 1 2 8 2 8 8 2 7 16 15 13 11 0 2 0 9 2
8 3 3 1 4 9 13 9 2
13 7 15 13 15 15 13 3 2 15 0 13 0 2
26 2 11 11 8 8 2 1 10 9 1 11 11 1 11 11 9 2 9 16 11 13 1 9 1 11 2
19 9 2 11 11 11 11 2 4 13 1 11 9 2 11 11 11 11 2 2
12 15 13 10 9 14 13 0 9 13 1 9 2
19 7 15 13 15 0 7 1 9 13 3 0 9 1 15 15 0 4 13 2
18 3 0 13 3 10 9 1 10 0 9 2 7 1 15 15 13 3 2
22 4 15 13 11 11 2 8 8 8 8 2 16 3 11 4 13 1 1 11 0 3 2
42 3 11 11 2 8 2 8 8 2 4 13 10 0 9 1 9 9 16 15 4 13 15 16 11 3 13 14 13 1 1 10 0 9 7 11 7 9 3 13 1 15 2
12 10 0 9 4 13 11 9 0 2 3 0 2
13 7 10 9 0 9 13 1 15 15 13 1 9 2
9 11 13 0 9 1 11 0 9 2
24 11 2 13 3 15 11 4 13 1 15 2 7 15 15 4 13 1 11 2 4 13 0 3 2
21 10 10 13 2 11 8 8 11 2 1 9 9 1 10 0 9 1 11 1 12 2
39 11 11 11 13 3 16 11 1 10 9 13 2 15 13 10 9 2 7 16 15 4 13 15 1 2 8 8 8 2 2 7 3 13 11 1 10 9 9 2
21 1 11 9 4 3 11 13 1 11 2 7 15 4 3 13 1 11 9 7 9 2
5 7 9 13 15 2
30 1 10 9 4 11 11 11 13 1 10 2 15 13 15 14 13 0 1 9 10 2 7 15 13 10 9 14 13 2 2
39 9 13 3 1 10 0 9 1 9 7 4 13 0 1 10 9 1 11 9 7 9 2 1 1 1 16 9 3 4 13 16 9 13 11 1 1 9 2 2
19 10 0 2 9 1 9 2 13 3 11 0 9 1 14 13 9 9 1 2
32 15 13 10 10 2 9 2 2 1 16 9 1 3 4 13 9 1 9 2 15 13 9 1 14 13 9 1 1 9 10 9 2
21 15 4 13 10 3 0 9 3 1 16 15 13 1 9 1 11 11 9 1 9 2
10 11 11 4 3 13 1 1 9 9 2
27 1 11 11 1 11 7 11 11 1 11 13 11 9 1 10 0 0 9 15 13 1 9 1 10 0 9 2
6 9 9 13 15 3 2
23 7 1 10 9 1 12 13 15 0 0 16 2 9 13 9 7 3 9 2 1 11 9 2
17 7 1 10 0 13 15 11 11 10 0 2 1 1 0 2 9 2
14 2 9 4 13 15 7 15 4 13 15 1 10 2 2
12 1 9 13 15 1 1 16 9 3 13 9 2
17 11 4 3 4 13 1 2 10 0 9 2 7 2 9 9 2 2
19 7 1 10 0 9 2 1 10 15 1 9 1 16 15 4 4 13 1 2
8 2 15 13 15 13 9 2 2
18 1 11 13 0 11 11 1 10 0 1 10 10 0 9 9 4 13 2
24 3 1 10 0 9 1 9 1 12 13 9 15 1 9 2 12 9 1 2 13 1 10 9 2
17 2 15 13 10 10 14 13 1 9 2 9 2 9 7 9 2 2
48 0 13 2 2 4 3 0 13 3 0 14 13 1 3 0 2 7 3 0 2 1 11 1 11 1 12 2 9 15 13 9 9 2 8 8 2 2 2 9 2 15 13 11 1 12 1 9 2
10 15 13 3 1 0 9 3 1 3 2
25 12 9 1 16 11 13 10 9 2 13 11 11 1 9 12 1 9 1 11 9 1 11 1 11 2
10 12 9 0 4 9 13 9 1 11 2
19 1 10 0 9 13 11 0 9 1 9 15 13 0 1 14 13 11 9 2
7 1 15 13 9 1 11 2
11 9 1 13 12 1 9 1 9 1 11 2
20 0 13 10 0 9 2 0 9 2 9 4 1 0 9 1 0 1 0 9 2
14 7 16 3 9 13 1 11 0 2 13 15 10 9 2
15 11 13 1 1 9 7 9 4 0 1 0 9 1 9 2
18 7 1 10 0 1 10 9 13 15 3 9 11 13 1 2 7 9 2
25 15 13 3 1 10 9 2 7 1 15 2 9 13 0 7 0 2 0 7 0 2 13 11 9 2
7 0 0 2 13 10 9 2
16 15 13 0 0 1 10 2 1 11 11 1 10 9 1 11 2
28 15 13 1 3 15 13 2 15 11 11 13 15 16 15 1 10 0 9 1 12 13 9 2 9 1 9 2 2
27 9 4 13 1 10 0 9 1 16 0 9 4 13 14 13 15 9 1 9 1 14 13 10 9 1 9 2
9 9 13 1 9 7 9 1 9 2
11 7 1 7 1 9 4 11 13 0 9 2
26 10 0 4 13 11 11 11 7 10 2 11 13 9 10 16 15 13 2 7 10 9 1 10 0 9 2
7 7 15 13 15 15 13 2
14 0 2 0 2 3 0 2 0 0 2 7 3 0 2
6 0 13 15 1 9 2
28 7 11 11 2 7 0 7 0 2 15 1 9 9 1 9 1 9 3 4 2 13 9 1 10 0 9 2 2
27 1 11 11 4 15 13 0 16 15 13 15 14 13 1 11 11 11 14 13 11 1 10 0 2 0 9 2
25 11 11 11 7 11 11 13 10 12 15 4 13 15 13 14 13 3 11 9 1 14 13 1 9 2
20 4 15 13 1 14 13 11 0 9 1 0 9 2 4 15 13 11 11 11 2
19 10 0 1 10 9 4 15 3 13 2 15 0 1 15 3 13 1 9 2
37 15 13 0 2 0 0 2 4 13 15 1 1 10 0 9 7 9 2 7 13 3 1 0 3 15 4 13 9 3 1 3 14 13 15 0 0 2
19 3 13 15 1 9 0 2 7 15 13 1 10 9 3 1 9 7 9 2
11 1 11 7 9 13 9 0 0 1 11 2
7 0 13 11 13 11 9 2
14 11 13 9 2 10 9 1 9 1 10 0 9 2 2
10 1 10 9 13 15 11 7 11 9 2
19 10 0 7 0 0 9 13 15 1 10 0 9 1 9 1 11 9 12 2
22 12 9 13 2 15 1 1 9 0 9 1 11 9 1 9 1 7 3 3 1 9 2
9 1 11 9 4 10 12 13 1 2
6 11 13 10 9 3 2
9 2 15 13 15 3 0 15 13 2
12 3 13 10 9 2 7 3 13 10 9 2 2
5 0 2 7 0 2
28 15 13 0 1 10 10 11 15 13 16 9 4 13 0 1 10 0 9 1 10 0 9 1 11 1 9 1 2
15 15 13 1 11 16 11 11 13 10 9 1 9 3 1 2
6 7 1 11 0 9 2
12 2 8 8 8 8 2 8 8 8 8 2 2
8 11 11 13 3 3 11 9 2
5 15 13 3 11 2
5 13 10 0 9 2
4 9 0 9 2
4 1 9 9 2
5 1 0 1 0 2
3 0 0 2
3 9 0 2
3 9 13 2
3 0 9 2
3 9 0 2
4 0 1 9 2
24 15 13 0 3 9 16 11 9 2 11 11 2 13 16 10 0 9 4 13 0 1 12 9 2
9 15 13 3 10 0 15 13 15 2
5 3 3 10 0 2
11 10 0 4 0 4 13 1 12 9 3 2
12 11 0 9 13 1 9 0 0 1 9 9 2
19 7 9 1 13 15 0 0 1 9 1 0 2 0 9 1 10 0 9 2
21 0 13 15 10 9 1 12 1 9 9 2 11 7 11 2 15 13 1 1 9 2
2 11 2
10 10 9 13 1 2 7 15 13 1 2
2 11 2
5 7 15 13 0 2
2 11 2
10 6 2 15 13 1 7 15 13 1 2
12 7 10 9 15 13 1 2 15 13 3 1 2
30 15 13 1 10 9 1 10 0 9 2 15 13 7 13 2 16 15 3 13 10 0 9 10 1 9 2 15 13 3 2
8 9 13 2 15 13 7 13 2
9 11 11 13 10 9 3 1 12 2
16 1 10 12 9 15 4 13 1 10 9 2 4 9 13 9 2
13 7 0 13 15 0 1 1 0 9 1 9 9 2
28 0 13 15 3 16 9 0 9 2 11 11 2 13 1 11 9 7 13 16 10 0 9 4 13 1 12 9 2
19 0 1 11 2 15 1 9 1 11 13 1 11 2 13 9 1 0 9 2
17 15 13 1 9 16 10 9 1 9 13 0 1 1 10 10 9 2
17 7 1 9 13 9 1 9 2 15 3 13 0 0 1 11 9 2
18 7 16 11 13 9 2 4 15 1 10 0 13 9 1 10 11 9 2
10 3 13 15 10 9 15 4 13 0 2
18 16 3 9 13 9 1 9 2 13 15 1 14 13 1 0 1 0 2
21 16 3 15 4 13 2 13 15 0 13 3 11 7 11 15 13 0 0 0 0 2
20 16 3 9 7 0 9 13 1 9 2 13 15 1 0 9 10 9 7 9 2
13 9 0 9 13 10 0 0 9 1 10 0 9 2
10 9 0 9 13 9 1 10 10 9 2
10 15 13 0 0 3 15 9 13 15 2
15 1 15 15 13 14 13 15 0 0 2 13 9 0 1 2
17 9 13 3 0 1 16 9 2 9 2 9 7 9 4 13 9 2
9 9 1 9 13 1 3 9 0 2
16 16 11 11 0 9 13 1 2 13 9 1 14 13 9 3 2
7 7 15 13 3 0 9 2
35 10 10 9 13 16 9 0 3 13 1 14 13 15 1 9 1 9 1 14 13 2 9 2 10 9 1 16 15 13 15 1 9 7 9 2
28 1 10 9 2 1 1 1 16 10 0 9 4 13 15 10 10 9 2 3 3 9 2 2 13 3 9 0 2
11 3 13 9 3 10 9 1 9 1 9 2
20 15 13 1 3 9 3 12 1 9 1 16 9 7 9 3 13 9 1 9 2
26 10 10 2 3 3 0 2 13 16 15 0 13 13 9 15 13 10 0 0 9 2 10 0 9 2 2
12 7 3 0 15 4 13 2 13 10 0 9 2
25 10 9 9 13 3 0 0 9 1 9 7 1 9 4 13 10 0 9 2 4 0 9 4 13 2
13 7 3 4 9 1 9 13 10 0 9 1 15 2
31 1 9 9 13 15 0 1 15 16 9 1 7 0 4 13 14 13 9 1 9 1 14 13 9 1 14 13 10 0 9 2
5 15 13 15 0 2
25 11 11 11 11 7 11 11 11 2 12 1 10 0 9 1 10 0 9 7 9 2 13 1 9 2
24 15 13 15 0 0 14 13 9 1 14 13 1 9 9 1 14 13 9 1 14 13 1 9 2
12 10 0 9 4 13 10 10 2 7 13 1 2
22 10 0 15 4 13 15 2 13 3 0 0 9 16 15 3 13 10 0 9 1 9 2
4 3 13 9 2
15 9 13 1 9 2 9 1 9 7 10 0 2 0 9 2
17 0 13 9 1 9 7 9 3 0 16 9 4 13 10 9 0 2
9 15 13 3 15 3 13 15 1 2
16 9 4 13 9 0 9 0 15 9 1 9 3 4 0 13 2
24 10 0 9 4 0 3 13 1 9 2 7 15 13 1 0 9 9 15 4 13 10 0 9 2
24 1 10 0 9 1 9 13 0 9 3 1 10 0 9 2 7 3 13 9 9 1 9 0 2
24 4 10 0 9 15 13 1 13 0 2 4 10 9 9 1 9 13 1 2 13 0 1 9 2
7 9 13 0 1 14 13 2
10 0 9 7 3 10 9 1 9 9 2
8 7 1 14 13 15 0 0 2
4 1 9 9 2
20 0 9 2 7 0 10 0 2 13 15 0 1 10 9 15 13 10 9 1 2
19 9 13 3 0 2 16 9 13 9 2 7 15 13 1 9 7 1 9 2
12 3 13 10 9 3 15 4 13 1 1 15 2
18 1 9 1 0 1 0 9 13 9 1 9 3 1 1 9 1 9 2
7 7 9 13 3 1 9 2
7 15 4 13 9 1 9 2
48 15 13 3 10 9 1 9 1 16 15 13 1 14 13 0 14 13 0 9 7 0 9 1 10 9 3 15 13 9 15 13 9 7 9 9 2 16 15 13 1 10 9 3 9 13 0 9 2
14 16 15 4 4 13 2 13 10 9 0 0 1 9 2
24 7 15 13 16 15 13 0 0 14 13 10 9 1 11 11 2 7 15 0 3 1 10 9 2
8 15 13 3 0 9 1 15 2
15 9 9 4 4 13 3 0 9 16 9 4 13 10 9 2
8 10 0 0 9 4 3 13 2
26 15 13 15 13 0 0 14 13 10 9 15 13 10 0 9 9 1 9 1 9 3 0 1 12 9 2
5 13 10 0 9 2
4 0 9 13 5
3 0 9 2
2 13 2
2 9 2
4 15 1 3 2
4 0 1 11 2
10 15 13 3 3 11 15 13 1 9 2
12 9 1 11 13 1 10 9 2 16 9 13 2
7 7 10 0 13 1 9 2
7 9 1 10 9 13 1 2
13 15 4 13 0 14 13 10 0 11 1 9 9 2
18 9 12 13 1 12 7 13 10 9 1 15 15 4 13 9 10 9 2
7 3 4 9 13 0 9 2
16 15 4 13 0 16 9 1 11 4 13 3 0 9 1 11 2
18 9 13 1 15 10 1 9 0 9 2 15 3 13 12 9 1 9 2
20 3 11 2 15 3 13 3 0 1 14 13 0 9 2 13 12 9 3 0 2
6 7 15 13 10 9 2
42 0 16 10 0 9 2 11 12 2 13 0 9 1 9 1 10 0 9 2 10 0 9 7 9 2 15 13 16 9 4 13 10 9 9 4 13 2 13 11 9 9 2
21 15 13 3 10 0 2 0 9 2 15 9 13 0 9 1 14 13 1 10 9 2
8 1 10 0 9 2 13 15 2
21 1 9 7 9 1 0 9 7 5 7 0 9 1 0 9 1 9 2 13 10 2
31 9 1 11 13 0 0 2 7 15 4 13 1 0 9 16 9 2 11 11 2 13 1 9 7 9 16 11 4 4 13 2
23 9 0 0 9 2 3 13 1 11 2 13 1 9 1 9 7 13 3 3 0 1 9 2
12 15 4 0 13 10 0 15 4 13 10 0 2
15 16 3 15 4 13 2 13 9 1 0 9 1 0 9 2
16 7 11 2 1 0 11 1 12 9 2 13 10 14 13 1 2
19 1 1 0 9 4 9 3 13 12 0 9 1 12 1 10 9 1 9 2
8 15 13 10 9 1 12 9 2
25 3 13 9 0 2 3 16 9 1 9 3 13 10 9 1 12 9 0 15 9 13 0 1 13 2
41 15 13 0 1 9 2 15 1 10 0 4 4 13 10 0 9 2 7 3 0 1 9 1 10 9 15 1 1 13 1 10 1 10 0 9 0 7 0 0 9 2
11 10 0 4 13 9 2 7 13 15 3 2
33 10 0 9 1 9 4 15 13 1 16 9 13 3 0 0 16 15 2 3 13 1 9 1 15 16 15 4 13 10 0 9 2 2
32 14 13 9 1 0 9 13 10 0 10 9 4 13 2 3 16 3 15 14 13 9 4 13 0 7 3 13 11 11 12 9 2
12 15 4 0 13 9 1 1 9 1 0 9 2
10 3 4 15 13 0 0 1 10 9 2
16 9 1 11 13 0 16 10 0 13 7 13 0 1 12 9 2
58 1 0 9 3 1 9 13 15 3 1 14 13 1 16 9 13 15 2 3 16 15 13 0 9 1 9 1 10 9 9 13 2 3 3 1 11 7 3 1 11 2 1 3 14 13 9 15 4 13 10 12 0 9 2 11 7 11 2
14 10 0 9 4 13 1 9 1 7 4 13 1 15 2
20 7 15 13 1 9 1 16 9 4 13 3 0 1 16 10 0 9 13 1 2
11 9 4 1 13 9 2 13 9 15 1 2
7 15 13 9 0 9 1 2
24 7 0 9 1 10 0 9 13 16 7 9 2 9 7 9 13 1 14 13 10 0 0 9 2
39 10 0 0 9 2 10 9 15 4 13 10 0 9 1 10 9 7 15 0 2 16 10 0 9 4 13 2 4 13 10 0 9 1 9 1 10 0 9 2
15 10 0 4 13 2 9 1 9 2 0 1 10 0 9 2
11 7 3 13 15 1 3 0 9 15 9 2
10 10 0 9 13 0 1 9 1 9 2
15 15 13 0 9 16 9 3 13 1 1 10 0 0 9 2
17 15 4 13 7 13 7 13 10 9 9 0 0 1 9 1 9 2
18 1 10 0 9 13 2 15 2 11 2 11 2 11 2 11 7 11 2
24 0 13 9 0 0 2 11 2 11 2 11 7 9 13 1 2 7 9 13 1 9 10 9 2
14 3 13 3 10 9 1 9 2 7 13 3 1 9 2
30 1 10 0 9 4 9 13 10 11 1 9 1 2 1 14 13 9 16 15 4 13 10 0 9 16 15 0 13 13 2
17 0 4 9 13 2 16 9 3 4 13 3 0 9 15 4 13 2
32 1 9 2 13 11 11 2 10 1 0 9 9 2 13 9 15 1 3 1 14 13 16 15 13 0 9 1 10 9 15 13 2
24 9 13 0 7 0 0 1 9 1 14 13 10 0 9 1 9 1 10 9 1 15 1 3 2
15 1 10 9 4 15 13 16 15 13 0 1 15 1 9 2
9 3 3 9 13 0 1 0 9 2
7 15 13 1 9 1 9 2
9 7 15 13 9 0 1 9 3 2
9 15 13 1 10 0 9 7 9 2
10 3 10 9 4 9 13 1 9 1 2
24 1 9 1 9 15 9 1 11 13 1 2 13 9 9 3 1 3 1 10 0 9 14 13 2
11 10 0 9 13 0 14 13 9 1 9 2
37 1 11 13 9 2 15 3 13 7 11 7 11 11 2 1 1 0 13 9 1 0 2 0 0 9 2 0 15 7 10 0 7 9 1 13 3 2
8 11 13 3 0 9 0 9 2
27 1 0 9 4 15 1 9 13 0 9 1 11 1 1 11 2 7 11 9 13 0 1 1 10 10 9 2
32 1 11 13 9 2 0 0 2 14 13 10 0 9 1 1 11 7 1 1 11 2 1 11 4 9 13 12 9 9 1 9 2
34 10 0 9 9 13 1 9 1 11 11 1 11 1 9 9 1 14 13 10 9 1 9 1 9 2 13 3 16 9 4 13 3 1 2
11 16 9 13 1 2 13 15 15 10 3 2
10 15 13 1 10 9 9 9 4 13 2
36 9 1 14 13 10 9 15 3 4 13 9 1 10 0 9 2 15 13 0 1 1 9 1 0 9 7 15 3 13 3 0 2 13 3 0 2
18 16 0 4 13 15 2 3 0 1 11 2 13 0 1 9 0 9 2
10 0 9 13 10 0 9 16 9 13 2
5 13 10 0 9 2
5 9 4 3 13 5
3 13 9 2
2 9 2
19 11 13 9 7 9 1 9 2 7 13 1 9 1 10 0 9 1 9 2
9 14 13 1 15 13 14 13 9 2
2 9 2
8 9 13 9 2 7 1 0 2
15 10 0 13 3 16 1 10 9 4 9 13 1 10 0 2
34 9 15 13 9 0 2 10 0 9 11 11 2 13 3 2 10 0 9 2 2 15 0 13 14 13 1 10 0 9 1 10 0 9 2
22 15 13 15 16 15 13 11 11 9 2 2 11 1 10 9 2 2 1 11 0 9 2
14 3 13 15 1 9 7 13 15 1 9 1 0 9 2
30 10 9 4 0 13 1 10 10 1 10 9 1 9 1 9 7 10 9 2 6 9 2 1 14 13 9 1 14 13 2
48 9 11 13 4 13 1 10 10 9 2 7 15 4 13 16 9 1 9 9 3 13 9 1 10 0 9 7 10 0 9 2 7 16 15 3 4 13 15 1 2 0 2 2 3 11 0 13 2
19 3 4 15 13 9 1 10 0 7 0 9 2 7 1 9 9 13 0 2
28 9 9 13 9 2 9 7 9 1 9 2 1 9 11 11 9 1 9 15 4 13 1 10 0 9 1 12 2
24 9 4 3 13 9 1 2 11 11 11 8 11 11 2 1 0 9 1 10 0 9 1 9 2
11 11 13 10 0 7 0 9 1 10 9 2
11 15 4 3 13 16 9 1 9 13 9 2
24 15 4 13 9 7 9 1 1 14 13 9 1 9 1 11 11 11 2 11 11 7 11 11 2
27 11 2 1 0 2 13 14 13 15 3 14 13 0 1 10 9 1 14 13 16 15 13 7 13 10 9 2
14 11 13 3 10 9 1 0 9 15 3 4 13 0 2
16 10 9 1 10 0 9 1 11 13 16 15 3 13 0 9 2
17 1 12 0 4 15 13 1 10 0 7 1 10 0 0 0 9 2
6 10 9 13 3 0 2
26 3 2 15 13 0 0 9 1 10 0 9 2 1 9 1 15 2 7 13 11 1 9 1 0 9 2
11 10 9 13 11 1 9 1 9 1 9 2
28 9 15 4 13 1 9 4 3 13 15 1 2 9 2 9 1 11 9 14 13 2 7 15 4 0 3 13 2
30 16 9 13 14 13 9 1 15 1 9 7 9 2 13 15 3 10 0 9 1 11 1 10 9 15 13 1 0 9 2
19 1 11 4 10 0 9 1 11 11 2 11 11 2 13 9 1 9 10 2
11 3 13 15 3 16 0 9 13 1 9 2
24 15 13 0 16 11 3 13 9 1 15 2 7 3 13 15 1 9 1 16 15 13 9 0 2
3 9 13 2
2 7 2
2 0 2
4 10 0 9 2
13 13 15 0 14 13 9 2 9 2 7 0 9 2
7 4 15 13 10 0 9 2
9 7 15 13 15 0 1 10 9 2
19 10 9 13 15 9 1 14 13 1 1 0 9 7 13 0 9 1 11 2
20 1 10 9 10 12 9 15 13 1 10 9 2 3 15 13 2 9 13 2 2
18 1 9 13 15 2 0 9 2 2 10 9 1 9 15 13 12 9 2
20 16 12 0 9 7 9 13 3 2 13 15 2 1 10 9 1 15 2 0 2
26 15 13 15 1 9 1 9 2 0 9 2 0 9 2 0 0 2 0 0 2 0 9 7 0 9 2
16 9 11 11 13 0 9 10 1 14 13 1 10 2 9 2 2
13 15 13 16 10 0 9 1 9 13 9 10 0 2
12 7 15 13 0 0 1 16 15 13 3 9 2
36 15 13 0 0 0 16 15 4 13 10 0 9 2 16 15 4 13 10 0 9 7 16 15 4 13 10 0 9 2 1 9 2 14 13 9 2
25 9 13 1 16 15 13 1 0 9 2 9 13 9 2 7 9 13 16 10 9 1 15 13 0 2
31 1 10 0 9 1 9 1 9 13 0 1 15 14 13 10 0 9 2 1 9 1 16 11 11 11 11 13 10 0 9 2
13 9 13 9 7 13 1 9 15 15 13 13 0 2
24 9 13 9 1 14 13 2 0 0 2 2 7 1 9 13 15 1 9 2 3 1 9 2 2
15 10 9 1 15 13 3 10 9 1 0 9 1 9 10 2
32 15 13 16 15 3 13 0 0 14 13 1 0 9 1 9 2 16 15 13 2 10 0 2 16 9 0 3 13 1 0 9 2
15 9 4 3 13 1 16 15 13 1 2 0 0 9 2 2
12 10 12 10 9 4 13 0 1 2 13 11 2
15 15 13 10 0 9 3 0 16 15 3 13 1 15 0 2
8 7 3 4 10 9 13 0 2
7 13 15 0 10 0 9 2
13 7 13 15 0 1 9 1 0 9 14 13 0 2
11 2 10 0 9 13 1 0 3 0 2 2
23 15 13 15 13 9 16 15 13 14 13 0 0 2 16 15 13 15 0 7 13 0 9 2
26 15 13 9 1 0 9 2 7 13 16 9 13 9 2 3 16 9 3 4 0 13 3 1 0 9 2
8 9 13 10 0 9 1 9 2
12 7 13 15 0 0 0 14 13 10 0 9 2
6 4 15 13 3 0 2
6 4 15 13 1 9 2
13 13 15 3 0 1 15 9 14 13 1 0 9 2
7 13 15 0 10 0 9 2
17 7 4 15 13 15 9 1 0 9 1 9 2 0 9 7 9 2
4 9 4 13 2
44 15 13 14 13 1 2 13 10 9 1 9 2 3 15 4 13 10 0 9 2 13 15 1 10 0 9 2 7 13 10 0 9 2 13 0 9 7 13 0 9 1 10 9 2
8 15 13 1 14 13 0 0 2
6 13 15 2 11 11 2
4 15 13 15 2
2 9 2
2 9 2
3 0 9 2
4 15 4 13 2
5 12 9 1 9 2
5 1 9 1 9 2
6 1 10 0 9 9 2
5 1 10 10 9 2
12 15 13 10 0 1 15 2 7 15 13 15 2
13 13 15 0 3 3 14 4 13 1 10 0 9 2
8 3 13 10 9 1 1 11 2
10 11 11 13 15 7 13 9 1 11 2
31 1 0 12 9 4 15 13 10 0 1 14 13 10 9 2 10 9 1 14 13 15 1 15 10 2 10 0 1 0 9 2
33 11 13 0 1 9 0 9 2 0 16 15 13 2 0 15 15 13 15 7 13 15 4 13 14 13 0 1 10 0 1 10 9 2
24 15 1 1 2 4 15 13 1 15 15 13 1 10 0 9 2 7 15 13 1 15 2 0 2
35 3 13 15 14 13 10 0 9 1 10 9 7 9 2 7 10 1 10 9 2 15 4 13 11 9 1 0 9 2 4 13 15 10 10 2
9 11 11 13 1 9 1 14 13 2
12 16 15 10 13 9 2 13 15 9 1 9 2
31 16 11 13 2 15 4 3 13 15 1 10 9 15 3 11 9 1 9 2 11 2 2 11 11 2 4 13 15 1 1 2
12 11 11 13 1 15 15 3 4 13 15 13 2
12 15 13 15 4 13 7 4 13 15 1 15 2
8 7 15 4 3 13 1 15 2
14 15 13 10 9 2 7 13 3 3 0 15 4 13 2
10 15 13 15 11 11 3 4 13 1 2
28 3 0 2 10 0 9 1 9 2 3 10 0 9 1 11 11 2 15 1 10 9 13 1 10 9 1 9 2
22 7 15 13 2 7 1 9 4 15 13 1 11 1 11 1 14 13 15 12 9 9 2
7 15 13 3 14 13 9 2
7 9 13 16 9 13 15 2
15 15 4 13 10 0 9 1 16 15 3 4 13 1 9 2
10 15 13 3 3 16 15 3 4 13 2
6 7 0 4 15 13 2
6 11 9 13 1 9 2
49 10 9 15 13 10 9 2 9 7 9 2 4 9 1 15 15 13 11 7 9 1 2 16 15 13 15 2 3 15 13 16 15 13 15 7 3 7 15 15 13 9 13 1 9 1 0 12 9 2
25 0 4 11 13 9 1 14 13 9 2 7 15 13 10 9 2 10 9 1 0 9 1 11 12 2
42 16 11 3 4 13 1 9 2 13 15 3 3 9 1 15 2 15 15 1 0 9 4 13 1 16 15 1 9 13 0 0 1 9 1 9 7 10 9 1 10 9 2
11 15 13 10 9 1 10 9 15 13 9 2
11 10 0 1 9 13 3 0 2 3 0 2
6 15 13 0 1 15 2
18 7 10 9 15 13 1 10 9 2 13 1 16 9 1 0 9 13 2
8 15 3 1 13 15 1 15 2
19 7 15 13 3 0 15 2 7 15 13 3 3 16 9 4 13 7 3 2
11 7 0 3 1 15 2 16 3 13 9 2
11 1 9 13 11 1 10 9 10 0 9 2
5 3 15 13 0 2
33 4 15 13 1 9 2 4 9 1 10 9 13 1 10 9 15 13 2 10 9 15 13 1 7 10 9 15 0 4 4 13 0 2
10 9 1 15 4 13 9 16 9 13 2
5 0 2 1 13 2
7 15 4 13 0 1 15 2
10 7 15 15 4 13 2 4 3 13 2
9 7 4 13 2 13 15 1 1 2
7 10 9 13 10 10 9 2
15 15 13 0 3 9 16 11 9 4 13 0 1 11 3 2
17 9 13 3 1 16 15 4 4 13 2 3 13 15 15 3 13 2
12 1 0 9 4 9 1 0 0 9 3 13 2
6 1 9 2 1 9 2
13 7 1 14 13 15 9 1 9 2 0 9 7 2
7 9 1 9 13 0 0 2
26 15 4 3 10 9 13 0 1 14 13 1 9 1 16 10 0 9 3 4 4 13 1 0 0 9 2
30 7 16 15 13 11 9 2 1 14 4 13 15 15 13 1 9 1 11 11 7 11 11 1 10 0 9 1 9 9 2
12 7 11 11 13 0 11 9 2 4 15 13 2
3 0 15 2
13 7 1 11 9 13 10 9 15 13 1 0 9 2
9 3 3 13 11 11 9 1 9 2
9 15 4 1 15 13 1 1 9 2
17 3 13 15 1 1 9 16 9 0 3 4 13 0 1 1 9 2
16 3 4 15 13 9 1 10 9 15 4 13 0 1 10 9 2
6 7 15 4 3 13 2
10 7 4 15 13 0 1 16 9 13 2
23 1 9 9 13 15 3 0 1 16 10 9 13 16 10 2 9 2 13 14 13 0 3 2
11 7 15 13 16 2 9 2 13 0 3 2
4 10 0 9 2
11 15 13 10 9 1 10 0 9 1 11 2
19 9 13 2 9 13 9 1 0 9 2 9 13 15 0 7 0 1 9 2
5 7 11 13 15 2
14 10 9 7 9 4 1 10 9 13 9 10 1 9 2
34 15 3 1 13 3 10 9 16 15 0 13 15 1 14 13 1 10 0 9 7 16 15 10 9 13 3 0 1 9 16 15 13 3 2
3 7 15 2
18 1 9 1 11 4 15 1 9 13 1 9 11 7 3 3 1 11 2
2 0 2
11 15 13 16 15 4 13 0 0 1 9 2
10 3 13 15 9 1 9 15 4 13 2
8 15 4 13 9 2 13 15 2
8 15 4 13 0 1 15 3 2
37 13 15 9 1 2 13 15 2 13 15 1 9 2 13 11 3 7 3 2 3 16 15 13 9 7 16 15 4 13 10 12 9 0 1 10 9 2
12 15 13 0 16 15 13 1 16 9 4 13 2
8 15 13 0 1 10 15 3 2
7 7 3 3 13 15 3 2
17 9 1 9 13 15 1 1 10 9 3 15 3 13 9 15 13 2
26 13 11 0 2 4 15 3 13 1 16 15 13 10 9 9 1 11 16 15 4 13 1 9 1 11 2
5 0 2 1 13 2
9 7 13 15 3 15 4 13 15 2
14 13 15 16 2 15 3 1 2 4 13 15 1 15 2
7 15 13 1 3 9 0 2
8 15 13 10 9 1 11 11 2
3 3 13 2
3 3 13 2
14 13 1 3 10 0 9 7 9 7 13 15 1 9 2
50 15 4 0 13 15 13 9 2 7 1 3 9 13 15 15 3 1 12 9 9 2 15 10 4 13 1 10 0 9 9 2 7 15 3 4 13 9 9 7 3 3 3 13 10 9 15 4 13 1 2
7 13 15 1 15 2 11 2
8 13 15 2 3 13 15 3 2
8 15 13 10 9 0 14 13 2
5 13 10 0 9 2
4 9 1 9 2
4 13 15 0 5
4 13 3 1 5
4 4 13 9 5
13 15 4 0 13 16 11 11 11 13 10 0 9 2
17 15 13 3 3 0 0 1 9 7 13 0 1 0 9 1 9 2
11 7 15 13 3 16 15 13 9 1 9 2
13 15 13 3 3 10 0 15 13 9 1 1 9 2
29 15 13 0 14 13 15 13 3 16 11 11 11 1 12 9 3 13 1 9 1 11 9 1 14 13 9 3 1 2
13 0 13 13 15 0 14 13 1 9 1 15 10 2
5 15 13 0 0 2
38 7 16 10 9 3 13 14 13 1 9 1 10 9 2 4 15 13 0 1 16 15 0 13 10 9 1 15 10 15 15 4 13 3 0 14 13 1 2
31 0 16 15 13 0 9 2 3 0 9 7 9 7 3 13 15 1 16 15 3 13 16 9 1 11 4 13 3 1 12 2
9 11 11 11 0 9 13 11 11 2
29 15 13 0 9 3 0 1 11 2 13 10 9 3 1 11 15 13 11 9 1 11 9 1 14 13 10 0 9 2
39 7 15 13 3 1 9 1 11 9 2 15 13 3 3 1 9 1 11 2 7 3 0 15 13 4 15 3 3 13 16 11 3 13 10 9 1 0 11 2
21 3 4 15 13 7 0 1 11 7 13 15 1 12 7 15 1 10 9 15 13 2
23 1 9 1 10 0 4 15 0 13 9 1 11 1 16 15 4 13 10 0 9 1 15 2
8 0 13 4 15 13 10 10 2
3 7 9 2
3 13 3 2
14 16 11 13 9 2 13 15 1 9 7 9 1 11 2
6 15 13 1 1 9 2
18 15 13 0 1 10 9 15 4 13 1 11 7 13 15 13 1 9 2
15 3 4 15 13 3 7 4 13 1 11 1 9 7 9 2
56 9 1 13 15 0 16 15 3 3 13 15 10 15 4 13 2 7 9 2 15 13 1 15 12 9 1 9 7 3 9 2 16 9 2 7 0 9 2 11 11 11 2 13 0 3 1 11 1 9 7 10 0 9 1 9 2
28 11 13 1 10 9 1 9 1 9 2 0 1 15 15 13 1 11 2 3 9 13 9 1 9 1 9 3 2
7 9 13 3 13 1 15 2
18 10 9 1 9 13 10 9 1 16 11 13 0 9 1 9 0 9 2
10 10 9 2 3 2 1 10 9 9 2
5 9 13 3 15 2
13 7 0 13 11 11 1 9 1 10 0 9 9 2
4 2 9 2 2
16 2 13 1 9 2 3 2 3 15 15 13 2 1 10 9 2
10 1 10 9 13 15 0 1 11 9 2
27 0 1 10 10 9 4 15 13 16 10 9 2 9 7 3 2 13 1 1 10 0 9 9 1 0 9 2
35 15 13 11 11 11 1 11 2 1 0 1 16 15 10 4 13 1 12 9 1 0 9 2 2 15 13 11 1 0 9 1 10 0 9 2
9 15 13 3 11 11 9 1 11 2
12 2 15 4 13 16 11 4 13 1 10 0 2
43 15 13 0 3 1 14 13 10 9 2 2 7 15 13 10 10 11 15 1 9 1 11 13 1 10 0 9 1 9 1 14 4 13 11 1 0 9 1 10 9 1 11 2
17 1 10 10 2 3 3 3 0 9 2 13 11 3 0 9 1 2
20 7 15 4 13 16 15 1 9 4 13 15 1 10 9 1 0 9 1 9 2
11 15 13 3 14 13 16 15 13 0 3 2
13 10 0 9 1 10 0 9 2 9 7 3 9 2
9 0 9 13 15 1 10 9 3 2
46 16 11 2 1 0 2 2 3 13 1 14 13 1 11 2 15 4 3 13 9 1 11 7 11 11 2 15 13 0 9 14 13 2 2 13 15 0 1 10 9 1 9 1 10 0 2
8 9 13 10 0 9 1 11 2
23 15 4 11 4 13 1 16 15 13 14 13 9 1 11 2 1 0 10 1 11 0 9 2
18 3 13 15 14 13 15 1 16 9 1 10 3 0 9 0 13 9 2
10 7 3 4 15 13 11 11 11 0 2
27 11 13 10 12 9 1 11 2 0 1 11 2 3 9 13 0 2 7 11 2 15 1 9 13 1 9 2
23 7 15 13 0 3 2 3 9 13 14 13 9 1 2 3 2 9 2 15 13 1 15 2
4 0 3 1 2
37 9 13 0 12 9 2 15 4 13 16 15 3 13 9 1 11 11 11 2 7 3 1 10 0 9 15 13 9 1 10 12 0 9 9 13 9 2
7 11 4 3 3 13 9 2
11 15 13 3 3 16 9 13 0 7 0 2
19 9 2 3 9 1 9 1 0 9 2 13 12 9 1 10 9 9 13 2
16 3 13 15 0 0 12 9 1 10 9 15 13 1 1 9 2
3 7 9 2
23 1 10 9 1 1 12 2 3 9 13 7 9 3 13 10 0 9 2 4 9 1 13 2
16 15 13 9 15 13 10 9 1 14 13 9 1 14 13 15 2
11 10 0 9 4 13 10 9 7 13 9 2
24 1 11 4 10 0 13 15 2 1 10 1 14 13 10 0 9 7 9 1 9 1 0 9 2
35 15 13 10 9 11 13 1 1 2 10 9 15 1 9 13 12 2 12 9 1 10 9 3 9 1 9 1 10 0 9 4 13 0 9 2
8 13 3 9 7 9 1 15 2
5 3 1 10 9 2
14 10 0 0 1 0 9 13 16 15 3 13 10 9 2
41 10 0 13 0 14 4 13 15 0 9 1 2 14 13 10 0 2 0 15 9 13 15 13 0 14 13 1 1 9 1 10 3 0 2 9 2 1 11 11 11 2
7 15 13 9 1 15 1 2
43 7 3 13 15 3 0 16 10 12 15 0 2 1 1 0 2 4 13 15 0 13 10 9 3 0 7 0 9 1 15 10 2 11 11 11 2 11 11 2 11 11 3 2
9 7 15 1 15 4 13 1 11 2
12 11 11 11 4 13 1 10 9 1 11 9 2
41 15 4 4 13 10 9 1 9 1 11 1 10 0 2 7 15 4 2 1 15 2 13 10 9 7 9 1 1 9 1 14 13 1 1 9 1 0 9 1 9 2
10 15 13 3 15 13 1 9 1 11 2
10 3 3 9 16 9 1 9 13 9 2
5 13 10 0 9 2
5 11 11 1 9 5
2 13 5
4 4 3 13 5
4 13 3 1 5
4 13 1 9 5
2 0 5
21 15 4 10 9 13 2 10 11 2 16 9 13 0 1 14 13 1 9 10 9 2
21 1 9 4 15 13 10 0 9 1 2 9 2 2 9 7 2 10 0 9 2 2
24 11 11 4 13 15 14 13 9 11 11 7 11 11 0 9 1 10 9 1 2 9 11 2 2
6 15 1 15 13 1 2
7 15 13 3 3 1 9 2
25 1 9 13 15 0 16 10 0 9 13 1 16 9 4 13 10 0 9 16 0 9 4 13 1 2
11 15 13 3 14 13 16 15 13 15 0 2
16 1 11 0 4 15 13 1 1 16 10 0 9 13 1 9 2
15 1 0 9 13 10 0 16 11 7 11 4 13 9 0 2
51 1 9 4 9 1 9 13 0 9 2 9 13 0 2 9 3 0 2 9 13 0 1 9 3 2 1 10 9 1 9 2 2 7 1 9 9 4 9 13 15 1 1 9 1 16 9 13 1 1 11 2
14 7 15 13 10 0 9 1 0 9 1 9 15 13 2
33 16 15 3 13 3 2 13 15 1 0 9 10 0 9 1 14 13 15 10 1 1 1 16 9 9 1 10 9 9 13 1 9 2
14 1 9 13 11 0 7 0 16 9 4 13 0 1 2
28 3 13 2 11 11 2 7 13 9 1 11 1 11 1 16 9 13 10 0 9 1 16 15 13 16 9 13 2
24 15 13 3 15 16 9 13 2 7 15 13 3 3 1 11 2 3 11 13 14 13 1 9 2
14 16 11 4 13 9 0 16 0 9 13 2 13 0 2
17 9 13 3 16 9 1 15 14 13 13 1 16 9 3 4 13 2
26 0 13 15 1 1 16 9 0 13 1 1 9 7 16 11 13 1 0 0 9 16 10 0 9 13 2
5 10 10 13 9 2
16 7 6 2 15 13 15 0 1 11 1 1 10 0 10 9 2
6 15 13 0 1 15 2
12 7 1 9 9 1 9 4 15 3 3 13 2
19 15 13 11 9 1 16 10 0 9 4 13 2 10 0 9 3 13 1 2
13 9 13 0 7 0 3 1 10 9 15 4 13 2
20 10 0 13 16 9 4 13 1 10 0 9 1 0 9 2 3 0 1 9 2
20 3 4 3 11 7 11 11 13 15 3 1 1 9 15 15 0 3 4 13 2
26 15 4 3 13 1 1 9 7 11 11 11 9 1 9 1 11 2 7 15 1 9 13 11 0 1 2
23 15 1 10 9 1 12 9 13 16 15 0 3 3 13 9 1 11 15 13 9 1 11 2
24 15 13 3 16 12 9 1 0 9 3 13 9 1 9 2 3 11 4 13 15 1 14 13 2
27 9 11 5 11 4 3 13 15 14 13 9 11 11 7 11 11 0 9 1 10 9 1 2 9 11 2 2
6 15 1 15 13 1 2
7 15 13 3 3 1 9 2
23 15 13 3 1 0 9 2 10 3 13 10 1 16 15 3 13 0 0 2 12 9 2 2
10 9 4 15 3 13 15 0 1 1 2
25 0 0 13 15 16 11 13 16 2 9 2 4 13 0 9 1 0 9 7 0 0 9 1 9 2
29 15 4 3 13 10 0 9 7 10 9 15 13 14 13 0 9 7 13 0 9 3 16 9 13 9 3 1 11 2
11 16 11 0 13 15 2 3 13 3 0 2
3 8 8 2
11 10 0 9 1 10 0 9 13 15 3 2
12 0 1 9 13 11 11 1 11 11 1 9 2
41 0 0 1 10 9 0 9 2 1 11 11 1 9 2 15 4 13 10 9 9 1 9 1 11 2 13 15 16 9 13 2 0 9 7 9 2 1 10 0 9 2
9 15 13 10 9 1 14 13 1 2
18 9 13 3 16 11 0 13 9 1 10 0 9 2 1 10 0 9 2
6 3 13 15 1 15 2
29 16 15 13 15 15 13 10 9 1 0 10 0 11 2 3 13 15 10 0 9 2 1 10 10 0 7 0 9 2
55 0 1 9 2 3 11 13 15 0 1 7 13 9 1 11 11 7 11 2 16 11 4 13 15 1 11 11 11 2 4 11 7 10 0 9 13 1 14 13 1 16 15 1 15 1 0 9 4 13 1 1 10 9 9 2
5 1 9 2 6 2
26 7 3 4 10 9 1 11 13 10 10 1 14 13 1 9 1 10 10 16 10 0 9 4 13 1 2
11 15 13 15 15 13 2 10 0 9 2 2
6 3 15 13 9 0 2
41 9 0 13 3 16 11 13 10 9 9 9 1 11 2 15 1 10 9 4 13 0 0 2 7 15 1 1 1 16 10 0 9 1 9 13 3 10 9 1 11 2
31 16 15 4 13 10 9 1 0 1 10 0 2 4 15 3 13 9 1 16 9 9 1 15 4 13 0 0 1 10 10 2
19 10 9 13 11 11 10 0 0 9 1 14 13 16 11 3 4 4 13 2
24 9 2 15 13 16 9 4 13 0 1 9 2 4 13 1 10 0 9 1 10 9 0 9 2
25 10 9 13 1 0 11 1 14 13 9 2 7 15 2 3 0 11 10 2 13 16 9 4 13 2
31 11 4 13 2 7 16 15 13 2 13 15 0 10 9 1 9 15 13 9 2 0 0 10 9 2 1 14 13 10 9 2
24 10 9 4 15 1 10 0 13 10 9 15 10 9 1 9 4 13 15 1 9 7 0 9 2
27 7 15 13 0 16 9 13 16 15 13 10 0 9 15 4 13 9 7 3 9 15 4 13 10 0 9 2
7 3 0 13 15 11 9 2
5 13 10 0 9 2
4 9 1 9 5
3 10 9 2
3 0 0 2
17 9 11 11 13 1 10 9 16 9 3 4 13 10 9 1 11 2
18 1 0 9 1 9 4 15 13 14 13 9 1 15 15 3 13 9 2
21 3 0 9 1 9 1 11 8 11 2 11 1 11 11 2 13 10 9 10 9 2
19 10 0 9 1 9 1 9 7 9 13 9 1 15 1 9 1 9 10 2
24 15 13 1 16 15 4 13 1 9 1 9 2 9 7 13 15 1 9 1 10 9 1 9 2
18 1 16 15 4 13 1 9 14 13 10 9 1 9 1 11 3 0 2
9 7 15 13 3 0 9 1 9 2
19 7 9 2 9 7 9 1 0 0 9 13 10 9 1 10 0 0 9 2
21 16 9 11 13 1 10 9 2 13 0 9 0 7 4 0 13 1 10 0 9 2
23 3 13 10 0 9 1 9 10 9 1 0 9 2 10 0 9 7 10 9 1 0 9 2
22 10 9 13 10 9 1 16 9 13 10 9 2 3 10 0 0 9 3 1 13 1 2
17 10 12 1 12 9 9 1 11 13 10 0 9 1 10 0 9 2
30 11 13 10 9 1 10 0 9 1 9 1 10 0 9 1 0 14 13 0 9 15 13 9 0 9 1 9 1 9 2
23 11 4 3 3 13 9 1 14 13 10 0 11 11 1 10 0 9 1 10 9 1 9 2
22 3 0 13 10 0 9 7 0 9 1 10 9 16 9 4 0 13 1 10 0 9 2
41 10 1 9 0 9 13 15 10 0 9 16 9 13 3 0 16 15 4 13 1 9 7 9 1 2 7 9 13 1 1 10 0 9 1 0 9 1 9 1 9 2
30 15 4 13 10 9 1 2 7 1 11 9 7 0 9 13 15 10 0 7 0 0 9 2 3 3 0 9 1 11 2
11 0 9 13 0 14 13 1 10 0 9 2
27 9 13 0 0 1 9 1 9 7 9 13 0 0 0 2 13 9 1 11 9 7 13 1 9 1 9 2
21 1 10 0 9 13 3 9 0 0 9 1 9 7 10 9 1 0 9 1 11 2
29 10 1 10 0 0 1 10 9 1 0 9 13 10 0 9 1 11 2 15 13 10 0 9 0 1 9 1 9 2
21 15 13 10 9 1 3 9 1 9 13 2 7 15 13 3 0 1 14 13 15 2
22 16 9 2 11 2 13 11 4 15 13 9 1 9 1 15 9 13 2 10 9 2 2
11 15 13 15 9 1 11 4 13 9 1 2
29 7 16 9 1 11 13 14 4 13 1 0 9 2 13 3 9 7 9 1 11 1 9 2 9 7 9 10 9 2
19 15 13 3 3 16 9 1 14 13 0 13 15 9 1 15 14 13 0 2
4 13 0 9 5
2 0 2
3 0 9 2
2 9 2
10 1 9 13 11 0 1 0 7 0 2
7 9 1 9 13 11 9 2
7 15 13 15 1 0 9 2
17 15 13 3 3 9 1 11 15 13 1 0 9 1 11 1 9 2
24 9 13 3 0 10 9 1 10 0 9 9 1 15 10 7 10 0 9 15 13 1 1 9 2
22 10 0 9 15 13 0 1 11 2 4 3 13 14 13 1 1 9 9 7 9 9 2
10 15 13 1 9 7 1 9 7 9 2
26 10 3 0 0 9 1 0 9 2 11 11 2 11 2 1 11 2 13 16 9 4 13 1 0 9 2
42 11 4 13 1 12 0 1 14 13 9 1 14 13 0 9 2 7 16 15 13 9 1 12 9 3 2 13 9 0 10 2 14 13 9 1 10 0 0 9 7 9 2
10 15 13 3 0 9 15 13 10 9 2
32 10 0 9 1 9 1 11 1 11 2 11 11 2 13 9 1 10 0 9 3 0 1 9 3 13 10 0 9 1 0 9 2
18 11 11 2 9 7 9 2 13 10 3 0 15 4 13 9 1 9 2
26 7 1 9 4 10 0 9 13 1 11 2 10 0 9 11 11 2 15 4 13 12 9 1 0 9 2
13 1 9 9 4 3 10 0 9 1 9 13 15 2
17 0 9 7 9 13 0 1 9 7 9 1 11 11 11 2 11 2
18 3 0 4 0 11 4 13 1 9 11 11 2 15 13 9 1 9 2
13 0 9 13 0 0 1 14 13 10 0 0 9 2
36 9 11 11 13 3 11 9 1 9 1 16 9 13 0 1 15 1 14 13 0 9 7 16 15 1 0 9 1 9 1 0 9 13 0 9 2
16 10 9 1 10 0 0 9 13 3 16 15 13 10 0 9 2
28 11 13 1 1 10 0 9 2 7 0 3 4 15 1 0 9 4 13 0 0 9 2 13 1 11 11 11 2
32 3 4 11 13 0 9 7 13 0 0 0 9 1 16 15 1 9 13 10 0 9 1 10 0 11 0 9 2 11 11 11 2
37 15 13 10 0 7 0 9 1 10 0 0 9 16 0 9 2 1 9 1 9 2 13 1 0 1 9 2 7 13 0 2 0 7 0 0 9 2
23 7 0 9 4 13 1 2 7 9 10 0 9 13 1 10 10 9 2 4 13 1 9 2
13 1 9 13 10 0 9 1 9 1 0 7 0 2
5 10 9 0 9 5
2 9 2
3 4 13 2
7 15 13 10 9 0 9 2
13 15 15 13 0 1 14 13 9 13 3 7 0 2
21 15 15 13 0 1 14 13 9 2 13 0 9 7 0 9 4 3 7 0 13 2
12 9 1 9 13 3 0 9 1 9 0 9 2
16 9 13 12 9 1 15 15 13 9 7 9 1 9 1 9 2
14 12 9 1 15 15 13 1 9 2 13 1 0 9 2
13 10 12 0 0 9 13 1 12 9 1 9 9 2
8 11 3 13 1 12 9 0 2
33 10 12 0 0 9 1 9 9 13 1 3 12 9 1 9 9 2 16 10 12 0 0 9 13 1 0 1 12 9 1 9 9 2
15 15 13 1 10 9 1 9 15 11 11 3 4 13 1 2
38 10 0 4 13 1 9 2 11 11 8 8 11 11 2 2 15 11 11 13 1 1 9 1 9 1 10 0 0 9 15 13 9 1 14 13 9 1 2
33 1 10 9 1 9 13 15 0 16 9 2 9 7 9 4 13 1 9 15 4 13 10 0 9 16 15 13 3 0 1 15 10 2
36 1 10 9 9 0 9 4 15 7 10 9 3 4 13 2 3 16 9 7 9 13 0 7 0 2 7 15 13 0 9 7 0 9 7 9 2
28 7 0 9 2 0 9 2 0 9 7 0 2 0 9 13 0 0 1 16 15 4 13 14 13 9 1 12 2
15 1 15 4 15 13 16 15 3 13 0 9 3 7 3 2
20 2 9 2 13 9 15 4 13 0 9 1 9 1 14 13 0 9 7 9 2
9 9 13 10 9 7 9 0 0 2
17 0 9 13 9 2 9 7 0 0 9 2 9 2 9 7 9 2
10 11 4 13 7 13 0 1 10 9 2
20 16 9 11 13 10 0 9 1 12 2 13 15 12 7 13 1 12 9 9 2
24 16 10 0 9 11 13 10 0 11 9 1 2 13 9 12 9 0 2 7 10 0 9 0 2
22 1 10 0 0 9 1 9 1 11 4 15 13 14 13 10 2 0 9 1 9 2 2
27 1 9 0 9 1 9 4 9 1 9 2 9 7 9 1 9 1 9 13 10 0 9 1 10 0 9 2
16 3 4 15 13 1 9 1 2 7 13 0 0 1 2 9 2
25 1 12 13 15 0 14 13 9 1 11 11 13 16 9 3 13 9 7 9 1 10 0 0 9 2
17 15 4 3 13 7 13 9 16 15 13 3 7 9 13 10 9 2
11 16 9 13 1 13 0 9 1 0 9 2
24 1 9 1 11 1 9 13 15 15 15 13 0 2 7 3 13 0 0 2 15 13 15 0 2
35 10 9 15 13 1 9 1 9 13 0 9 7 9 1 14 13 9 7 13 1 0 9 1 9 1 9 1 16 2 9 13 1 9 2 2
12 3 4 15 13 9 2 16 15 13 3 0 2
4 10 0 0 5
2 13 2
2 9 2
6 4 0 9 13 1 2
5 13 9 0 0 2
17 1 10 0 9 13 12 0 9 1 14 13 9 1 10 0 9 2
25 11 0 9 4 13 1 9 1 11 11 2 9 3 0 9 1 0 9 7 0 9 3 1 9 2
36 16 0 0 0 4 13 9 0 2 0 9 7 13 15 1 1 9 2 4 11 11 1 10 0 9 13 15 1 10 0 9 1 0 0 9 2
44 16 9 1 11 1 10 0 9 3 13 10 0 0 9 1 10 12 9 1 0 9 15 3 13 10 13 9 2 4 10 9 3 13 14 13 9 9 1 14 13 11 0 9 2
19 16 11 13 10 9 15 0 11 11 13 1 1 2 13 3 9 1 9 2
27 3 4 15 3 13 0 9 1 9 16 15 13 16 11 4 13 9 9 1 10 0 2 0 7 0 9 2
14 15 4 13 3 0 14 13 9 1 10 0 0 9 2
15 7 3 16 11 3 13 0 9 1 9 2 13 9 0 2
13 15 4 13 10 9 1 0 9 1 10 0 9 2
35 10 9 13 10 0 9 1 9 2 9 1 10 0 9 7 10 0 9 1 14 13 1 14 13 9 1 9 1 0 9 7 9 1 0 2
13 10 0 0 9 1 14 13 10 9 13 3 3 2
11 11 13 0 9 1 9 10 12 4 13 2
19 10 1 9 10 13 1 9 16 10 13 1 0 9 2 0 13 1 9 2
31 10 0 9 13 1 9 1 0 9 2 3 15 13 16 7 13 15 1 9 7 13 0 7 15 13 15 7 15 13 0 2
15 3 13 15 0 1 14 13 11 9 2 7 13 15 9 2
12 13 10 0 9 14 13 11 9 7 10 9 2
15 1 9 13 10 9 0 9 15 3 13 9 1 0 9 2
16 10 9 1 0 1 11 0 9 9 13 0 9 7 0 9 2
18 15 13 9 1 9 11 11 11 9 1 9 1 14 13 10 0 9 2
17 3 13 11 9 15 13 16 0 9 13 10 0 9 7 3 0 2
18 1 3 13 15 3 9 1 10 0 9 16 0 9 13 0 7 3 2
21 11 13 3 9 1 14 13 10 0 7 0 0 9 1 9 15 4 13 0 9 2
35 15 13 0 14 13 3 9 9 1 9 1 7 9 7 9 4 13 1 10 11 3 0 2 0 7 0 9 13 7 13 1 9 1 0 2
26 11 0 9 13 1 10 0 7 0 9 9 1 14 13 10 9 3 3 1 9 2 7 1 9 0 2
6 9 1 9 1 9 5
2 0 2
5 2 9 2 11 2
2 9 2
18 9 16 9 13 0 1 0 9 2 0 9 7 9 13 10 9 0 2
15 9 1 9 9 13 0 13 9 1 0 0 9 1 15 2
40 14 13 9 13 0 0 2 1 10 12 9 4 15 13 1 0 9 1 2 10 10 2 2 16 9 1 11 7 9 1 10 10 9 0 13 15 1 1 9 2
8 15 4 13 1 10 0 9 2
22 11 3 0 9 2 11 11 2 13 9 15 13 0 9 1 14 13 1 9 12 0 2
24 11 11 0 9 13 11 9 2 7 15 13 10 9 14 13 16 11 3 13 0 9 14 13 2
12 7 11 11 13 15 13 1 14 13 10 9 2
22 15 13 0 16 11 11 4 13 11 1 9 1 9 15 13 11 0 9 0 1 9 2
49 11 13 3 0 3 1 3 14 13 1 11 9 2 7 3 4 15 13 15 10 0 1 14 13 15 1 9 2 3 16 15 13 10 0 9 16 15 1 11 13 16 15 4 13 10 9 1 15 2
22 0 4 15 13 15 0 1 10 0 9 15 0 13 15 1 9 14 13 15 1 15 2
13 11 0 9 2 11 11 11 2 13 10 10 9 2
15 15 13 3 1 1 9 7 4 13 10 9 9 1 9 2
43 11 4 13 0 1 10 9 1 10 9 2 7 13 9 1 10 0 9 2 7 1 16 15 13 9 1 9 9 0 15 15 3 13 0 1 15 15 13 14 13 9 9 2
37 1 9 1 10 9 13 15 1 9 0 14 13 15 3 1 2 9 2 11 2 1 10 9 1 9 2 0 9 2 0 9 7 9 1 11 11 2
12 3 4 10 0 9 13 15 0 1 0 9 2
22 1 10 10 9 4 9 1 11 1 0 9 3 1 9 7 9 2 13 0 1 9 2
14 11 11 11 13 3 3 0 2 7 13 0 1 9 2
25 15 4 13 0 1 9 2 7 4 13 0 1 9 1 9 1 9 1 0 9 1 9 7 9 2
18 11 0 9 2 11 11 2 13 9 7 13 15 3 1 10 10 9 2
37 11 13 1 9 2 7 10 9 13 9 15 13 0 9 2 7 15 13 16 9 1 11 7 11 13 1 0 9 2 3 16 11 0 0 9 13 2
26 10 1 10 9 4 13 0 0 9 1 9 9 2 7 9 9 4 0 13 1 9 1 9 1 9 2
5 9 13 10 9 5
2 9 2
2 0 2
4 15 13 9 2
11 15 13 10 9 16 15 13 9 1 11 2
26 10 0 1 9 4 13 12 2 7 15 13 0 3 15 9 13 1 9 2 7 9 13 0 0 0 2
21 10 12 15 13 2 13 10 9 15 13 1 9 1 11 9 15 4 13 1 11 2
24 1 7 1 16 15 0 3 13 9 1 11 2 15 13 1 9 2 2 4 15 13 9 3 2
5 15 13 9 0 2
20 15 4 3 13 15 14 13 10 3 0 9 14 13 10 0 9 10 0 9 2
22 11 7 11 13 0 2 13 9 2 15 13 1 14 4 13 2 9 2 1 9 10 2
11 11 13 0 16 15 13 9 2 13 9 2
20 15 13 9 1 7 9 1 2 16 15 13 0 1 14 13 9 11 7 11 2
9 15 13 16 15 13 0 7 0 2
7 3 13 15 0 7 0 2
22 15 13 10 0 9 1 10 0 9 15 13 1 16 9 4 13 9 1 10 0 9 2
26 15 13 3 3 0 1 14 13 10 10 9 2 13 15 2 16 15 4 13 9 1 10 9 1 9 2
16 3 13 15 10 9 16 15 4 13 1 9 1 2 9 2 2
17 9 13 1 9 1 9 2 1 9 7 2 3 0 2 1 11 2
36 15 13 1 9 1 9 2 13 0 9 2 7 13 16 15 15 13 11 13 9 1 12 9 2 0 3 4 13 14 13 3 10 9 1 11 2
23 9 13 15 1 14 13 1 9 2 13 1 1 9 7 13 16 15 13 0 1 1 9 2
36 9 10 2 13 2 9 2 2 15 13 0 1 0 9 1 9 2 13 0 1 16 15 4 13 1 16 15 13 3 14 13 0 9 1 9 2
23 15 13 9 7 9 2 7 10 0 9 13 2 1 9 2 16 15 13 9 9 7 9 2
24 9 13 16 15 13 9 9 16 15 13 12 9 0 2 7 13 15 13 11 16 15 13 12 2
29 0 1 13 9 7 9 0 0 1 16 9 4 13 10 9 16 15 13 10 9 2 7 3 13 9 1 11 11 2
18 10 0 9 1 10 0 9 13 16 10 0 13 9 1 10 0 9 2
6 15 13 10 0 9 2
6 15 13 10 0 9 2
8 15 13 9 1 10 0 9 2
26 3 0 13 15 1 10 10 9 2 16 15 13 16 9 13 0 9 1 10 0 11 9 15 13 1 2
9 10 0 9 13 16 9 13 9 2
8 3 13 9 7 13 1 9 2
20 7 15 4 13 10 9 1 3 14 13 16 9 4 2 13 10 0 9 2 2
19 6 2 3 0 13 15 1 9 9 1 9 2 16 15 13 15 0 9 2
35 9 13 1 0 9 1 14 13 15 1 9 2 16 9 13 1 9 1 14 13 16 15 13 16 9 15 13 1 9 1 9 2 13 0 2
12 15 13 0 1 10 0 9 1 10 0 9 2
21 16 9 3 13 1 1 9 1 9 1 11 2 13 9 9 1 1 9 7 9 2
5 9 13 1 9 2
6 7 9 13 1 9 2
33 1 1 9 1 10 0 2 0 9 13 10 0 9 14 13 15 1 0 9 2 10 0 9 15 4 13 1 10 9 10 0 9 2
13 2 15 4 13 14 13 2 2 13 10 0 9 2
8 2 3 0 1 3 0 2 2
5 9 1 0 11 5
3 0 9 2
6 11 9 13 0 0 2
10 3 4 11 13 11 11 14 13 9 2
19 11 9 1 11 13 10 0 9 1 16 11 4 13 1 3 1 0 9 2
23 11 7 9 11 11 4 13 1 0 9 1 9 9 1 9 1 9 2 9 1 9 2 2
24 0 1 11 11 2 15 13 10 0 0 9 1 11 11 11 2 13 15 3 1 9 10 9 2
21 2 15 4 13 0 1 1 11 11 2 13 10 0 9 1 9 1 10 0 9 2
19 9 3 13 16 10 0 9 11 4 13 1 1 2 3 13 1 1 9 2
19 16 11 1 12 4 13 0 9 2 13 3 9 10 0 2 0 11 11 2
20 2 15 13 10 9 15 13 9 0 1 9 2 2 13 11 0 9 11 11 2
12 9 7 9 13 10 9 2 7 13 10 10 2
22 1 12 13 11 15 0 0 1 15 9 9 10 9 1 9 13 15 1 9 1 11 2
38 16 9 7 10 0 13 0 1 11 11 7 10 0 9 1 7 1 9 2 13 15 0 3 0 0 2 3 16 9 13 1 9 1 10 9 7 9 2
18 15 13 10 0 11 11 15 13 9 1 10 0 9 1 9 7 9 2
13 10 0 9 13 0 0 9 1 11 1 10 9 2
13 1 9 1 10 0 9 13 0 9 1 11 9 2
7 15 13 10 12 0 9 2
22 15 13 10 0 0 9 1 14 13 11 9 7 13 1 9 1 10 0 7 0 9 2
41 15 4 13 1 16 9 13 10 3 0 9 1 14 13 0 9 1 11 11 2 11 2 11 2 11 2 11 7 11 1 9 1 9 15 13 10 0 7 0 11 2
20 11 13 1 10 0 7 0 9 1 11 16 3 11 7 11 13 9 1 12 2
40 11 13 10 0 9 1 11 0 9 2 7 10 0 9 13 2 1 10 10 2 16 11 13 3 0 2 0 2 0 7 0 1 14 13 0 1 0 0 9 2
6 11 13 3 0 3 2
35 16 11 1 11 9 13 16 10 10 9 13 0 1 14 13 1 10 0 0 9 1 7 1 11 2 4 15 3 13 16 11 13 1 11 2
24 10 9 1 9 1 11 13 3 16 11 4 13 3 0 10 0 9 1 11 7 11 4 13 2
21 1 12 4 11 3 13 1 12 9 9 2 1 12 9 9 2 1 11 7 11 2
11 10 10 9 4 0 13 0 10 9 1 2
23 15 13 0 1 12 9 10 0 9 11 4 13 1 9 1 1 12 9 1 10 10 9 2
43 3 13 3 11 0 9 1 11 16 3 10 2 0 2 9 7 3 0 0 9 4 13 10 2 9 2 1 11 1 12 9 1 9 7 9 16 11 7 9 4 13 9 2
41 1 10 10 12 9 4 11 1 10 0 9 13 1 9 7 9 1 1 10 11 2 11 2 11 11 2 11 2 11 11 2 11 2 11 2 11 2 11 7 11 2
11 11 13 2 1 15 2 0 1 10 9 2
6 9 1 1 11 13 5
2 9 2
15 0 11 4 13 12 9 9 1 9 1 14 13 0 11 2
21 13 15 10 9 15 13 16 0 9 13 1 1 11 3 0 15 4 13 10 9 2
5 0 9 13 0 5
4 0 1 9 2
12 15 13 3 0 14 13 16 9 13 15 0 2
16 15 3 1 10 0 9 15 13 9 10 16 15 13 0 0 2
4 13 15 0 2
15 0 3 13 9 1 9 1 9 3 1 16 9 4 13 2
11 10 9 4 13 16 0 4 13 14 13 2
7 15 13 0 14 13 9 2
5 7 0 13 15 2
11 7 9 1 10 0 0 13 3 10 9 2
18 15 13 15 15 1 0 9 13 10 0 3 13 9 14 13 10 9 2
19 11 11 13 10 9 1 9 2 7 13 0 16 10 0 0 13 9 0 2
5 3 13 15 15 2
5 7 15 13 0 2
8 9 13 0 16 15 13 9 2
24 0 13 15 7 9 2 9 7 9 15 13 0 1 14 13 16 15 13 1 9 12 9 0 2
5 9 13 0 9 2
7 3 4 10 9 13 0 2
18 15 4 3 13 10 12 9 10 2 0 2 2 16 9 13 3 9 2
13 7 1 11 13 15 16 15 13 0 14 13 9 2
5 15 4 13 1 2
5 3 13 15 9 2
9 1 10 9 13 15 10 1 9 2
15 3 0 15 9 4 13 1 10 9 2 4 9 13 3 2
15 3 13 15 1 9 16 11 11 0 13 1 10 0 9 2
8 1 11 13 9 3 0 9 2
24 3 13 3 0 9 9 1 9 2 0 7 0 16 2 0 9 13 10 9 9 13 1 2 2
10 10 0 13 16 3 0 13 11 9 2
24 11 11 13 11 7 13 3 9 3 13 2 3 9 1 14 13 9 9 2 2 0 9 2 2
7 3 15 13 15 1 9 2
20 11 11 2 0 9 2 13 3 3 9 4 2 13 10 9 1 10 9 2 2
4 15 13 0 2
12 3 13 15 2 3 14 13 9 1 9 2 2
2 6 2
19 9 13 3 9 1 14 13 16 15 3 13 0 7 3 13 9 1 9 2
21 13 16 15 1 9 13 10 0 3 1 15 13 16 10 0 9 13 9 1 9 2
19 7 1 0 7 1 0 9 4 15 13 1 14 13 9 1 10 0 9 2
25 15 13 0 9 2 7 3 3 0 9 2 13 14 13 3 9 1 9 2 1 9 7 1 9 2
9 3 13 15 0 14 13 1 9 2
11 15 13 3 14 13 0 1 9 0 9 2
23 3 4 3 9 10 13 16 9 13 1 9 2 1 9 15 4 13 7 9 15 4 13 2
15 9 2 13 15 9 2 13 15 9 2 13 0 7 0 2
13 15 13 15 1 10 9 9 4 13 9 7 9 2
28 10 9 13 16 9 4 13 0 9 2 0 0 9 7 0 9 1 14 13 10 9 1 10 0 7 0 9 2
21 1 9 4 15 1 9 13 1 9 1 3 0 9 15 13 0 1 9 1 9 2
11 15 13 0 16 10 0 1 9 13 0 2
7 9 2 9 2 0 9 2
8 15 13 10 10 13 1 9 2
14 10 0 9 2 15 13 9 7 9 2 13 3 9 2
3 3 9 2
6 13 15 0 1 9 2
2 9 2
2 9 2
9 0 1 10 0 9 13 1 9 2
11 7 13 15 3 0 1 14 13 1 15 2
10 0 9 15 13 1 1 9 1 15 2
8 9 15 2 13 2 1 9 2
7 9 15 13 1 0 9 2
6 9 15 13 1 9 2
9 9 15 3 13 15 1 9 10 2
6 9 15 13 1 9 2
6 0 9 13 1 9 2
5 0 9 13 9 2
16 0 9 15 3 13 14 13 1 9 2 13 9 1 1 0 2
13 9 1 9 1 9 7 9 13 0 9 1 9 2
16 9 13 1 9 1 1 9 1 14 13 0 9 1 10 0 2
12 15 13 0 3 0 9 2 7 1 7 1 2
10 15 13 3 0 16 15 3 13 0 2
14 0 13 1 1 9 2 7 0 9 4 13 1 9 2
11 16 11 11 4 13 15 1 9 1 9 2
3 15 13 2
18 9 13 3 16 10 0 9 15 13 1 2 0 0 13 1 0 9 2
6 7 13 1 10 9 2
5 15 13 1 9 2
11 3 13 0 15 13 0 14 13 1 9 2
6 9 1 15 13 0 2
14 1 10 0 13 15 0 1 16 9 4 13 1 9 2
17 0 9 1 16 10 3 13 0 3 2 7 16 15 13 0 1 2
4 9 13 0 2
16 3 0 15 9 13 9 1 9 2 0 0 1 10 0 9 2
32 1 10 0 13 0 1 9 7 9 15 13 1 10 0 9 2 3 9 1 10 9 16 9 7 9 4 4 13 1 0 9 2
9 3 13 15 0 14 13 0 9 2
19 7 1 10 0 13 15 16 0 9 4 13 0 2 7 1 10 9 0 2
28 15 15 13 0 1 9 7 9 2 13 0 9 15 3 13 0 1 14 4 13 3 9 2 0 2 4 13 2
29 10 15 4 15 13 1 15 16 15 4 13 1 9 7 9 2 1 10 9 7 9 15 13 10 0 7 0 9 2
7 9 4 3 13 1 9 2
15 7 15 4 3 13 15 1 14 13 10 9 1 10 9 2
15 15 15 13 9 2 4 13 1 0 9 1 9 7 9 2
13 7 13 15 3 2 13 15 15 1 9 7 11 2
22 15 15 13 1 0 9 2 4 13 0 1 9 1 0 7 0 9 1 9 1 9 2
10 7 15 4 13 16 9 1 9 13 2
30 16 15 0 13 16 9 13 10 9 1 15 10 2 4 15 13 0 1 14 13 1 15 2 3 16 15 13 0 1 2
41 7 2 3 0 2 15 15 13 1 9 1 10 9 2 7 15 13 15 10 3 2 4 3 13 0 1 14 13 1 16 15 4 9 4 13 2 7 16 9 13 2
13 7 15 4 3 13 9 3 1 2 10 10 2 2
29 16 0 9 13 0 9 13 0 2 13 0 9 1 15 7 13 0 9 1 10 0 9 2 15 13 15 15 1 2
16 16 9 13 9 7 13 9 1 9 2 15 13 15 15 13 2
3 0 13 2
26 15 9 9 13 15 0 0 1 10 9 7 1 9 1 15 2 15 15 13 1 9 1 10 0 9 2
6 1 9 1 0 9 5
5 9 7 0 9 2
3 0 9 2
3 0 0 2
9 9 1 9 1 11 13 3 0 2
19 3 4 10 0 9 1 10 0 9 13 1 10 10 2 3 0 0 9 2
23 11 13 1 9 2 9 2 7 2 9 1 0 9 2 2 2 8 8 8 8 2 2 2
13 0 13 15 3 4 13 2 7 15 13 10 0 2
21 1 11 13 15 10 9 1 0 9 1 9 1 0 9 7 9 1 10 0 9 2
20 1 0 13 11 9 1 9 2 10 0 9 7 9 1 9 1 10 0 9 2
21 11 0 9 13 2 9 1 9 2 2 2 8 8 8 2 2 1 10 0 9 2
12 3 13 9 10 9 1 9 1 9 7 9 2
19 9 13 9 1 9 9 16 15 13 9 7 10 0 0 9 0 1 9 2
7 9 13 16 9 4 13 2
21 0 13 9 9 15 3 3 13 0 9 1 9 1 0 9 1 14 13 1 15 2
6 9 4 15 13 0 2
24 9 13 16 0 9 2 1 10 9 2 4 13 16 10 13 10 9 7 9 2 9 7 9 2
22 9 4 13 14 13 9 1 9 7 9 1 9 1 9 2 3 14 13 9 1 9 2
16 9 1 10 0 11 13 9 1 10 0 0 9 1 10 9 2
8 9 1 9 1 9 13 0 2
8 3 13 15 10 9 1 9 2
10 3 13 15 9 1 9 1 0 9 2
28 1 10 0 9 3 0 13 15 1 16 0 13 10 9 1 16 9 4 13 0 2 7 16 10 9 13 9 2
14 15 4 2 1 9 2 13 0 15 13 1 9 9 2
15 3 13 15 16 0 9 13 0 0 1 9 1 0 9 2
34 7 11 9 13 9 1 9 1 10 9 3 16 2 9 2 13 15 15 4 13 1 7 9 15 15 4 2 1 9 2 2 13 2 2
12 1 2 9 2 13 10 0 1 2 9 2 2
18 1 0 9 13 15 0 14 13 9 1 9 7 3 9 1 0 9 2
15 10 9 1 9 1 9 13 3 13 1 10 9 1 9 2
33 1 11 9 1 0 9 1 0 9 0 1 9 13 10 9 0 2 3 13 2 1 9 1 9 2 9 1 3 9 1 0 9 2
34 3 13 15 10 9 1 0 9 1 9 1 0 9 2 15 13 1 11 2 1 10 12 9 2 7 9 2 9 7 9 1 10 0 2
14 1 0 7 3 13 9 3 3 0 1 14 13 9 2
9 9 13 1 15 7 9 7 9 2
11 0 9 4 13 10 0 9 1 10 9 2
5 0 9 1 11 5
6 11 4 13 0 9 2
18 9 4 3 13 1 9 2 7 15 13 3 0 3 10 0 9 13 2
23 0 1 10 0 9 2 11 7 11 2 4 11 3 13 3 1 9 16 15 13 0 9 2
22 1 11 4 0 9 13 1 9 2 7 0 9 4 0 9 4 2 13 2 1 9 2
23 1 11 13 15 0 0 7 0 1 15 2 7 3 13 15 3 16 9 0 13 10 9 2
8 1 11 4 15 3 13 9 2
19 11 11 11 11 4 13 9 0 1 11 11 11 11 2 15 13 0 9 2
35 15 13 10 0 9 1 15 15 4 13 1 10 2 0 9 2 1 9 2 16 9 2 1 0 9 2 13 0 1 12 0 9 1 9 2
16 11 13 0 0 1 9 16 15 13 1 9 1 12 9 3 2
28 0 13 0 1 9 2 9 11 11 2 2 9 11 2 2 2 15 4 13 9 1 0 0 9 1 12 9 2
54 1 9 1 14 13 1 1 10 9 1 0 9 2 7 1 2 0 2 9 1 9 2 13 2 9 11 2 3 9 1 11 9 1 14 13 9 2 9 2 1 10 0 9 2 1 9 1 9 2 0 9 7 9 2
14 11 4 4 13 16 15 13 0 9 1 2 9 11 2
16 15 13 3 1 11 9 16 9 1 11 13 14 13 15 0 2
21 7 9 0 9 13 3 1 0 9 1 11 9 2 7 13 10 10 9 1 9 2
13 11 13 9 1 14 13 0 9 7 14 13 9 2
13 15 13 3 9 1 14 13 9 7 10 0 9 2
15 3 1 10 1 10 9 4 15 13 0 9 1 0 9 2
25 11 0 9 1 10 10 9 13 10 9 2 7 3 3 10 9 1 15 15 4 13 15 1 11 2
19 11 13 3 1 9 1 0 9 7 9 1 0 9 1 14 13 0 9 2
16 10 0 9 2 11 2 4 13 7 13 9 1 10 0 9 2
28 1 9 1 14 4 13 1 9 16 15 13 12 9 2 13 15 3 9 1 11 10 9 7 9 1 10 0 2
13 0 0 9 4 15 3 13 0 14 13 9 1 2
14 11 13 3 1 10 0 9 1 0 9 7 0 9 2
10 15 13 9 1 16 15 4 13 9 2
16 1 9 4 15 4 13 1 10 9 15 13 10 9 1 9 2
12 9 2 10 0 9 7 0 9 13 1 9 2
6 11 4 13 10 9 2
10 11 4 13 11 1 9 7 0 9 2
16 15 13 1 9 0 15 13 15 16 15 13 0 9 1 9 2
13 15 4 13 0 1 3 11 4 13 3 10 9 2
17 15 4 3 4 13 16 2 9 11 2 9 9 13 1 1 9 2
6 15 4 13 10 9 2
12 0 9 13 16 2 9 11 2 3 13 0 2
5 3 13 15 3 2
3 0 9 2
3 13 9 2
21 1 14 13 1 9 1 11 4 15 13 1 9 0 9 1 15 15 13 1 9 2
25 9 15 13 1 11 13 0 0 0 1 0 9 2 0 13 0 13 1 10 0 9 1 0 9 2
16 13 15 0 3 1 9 2 13 0 9 1 10 9 1 9 2
19 3 13 15 1 0 9 7 13 15 13 0 16 0 7 0 0 13 15 2
38 3 13 15 15 16 15 13 9 1 15 14 13 2 1 9 2 1 0 9 2 0 2 0 2 0 2 0 7 0 2 0 2 0 7 2 0 2 2
24 9 13 10 0 0 9 2 15 13 1 14 13 15 1 15 15 13 2 7 15 15 3 13 2
17 15 13 3 0 9 2 0 1 0 9 7 9 1 11 1 9 2
30 3 13 15 0 14 13 2 16 15 13 1 0 9 2 16 9 13 10 0 10 2 7 0 2 9 1 10 0 9 2
19 10 9 1 0 9 2 13 1 2 13 3 0 15 13 3 1 0 9 2
31 1 9 4 9 13 0 9 2 15 4 13 0 2 2 13 1 9 2 2 7 13 9 1 14 13 15 15 13 15 1 2
28 3 15 13 1 2 1 11 2 13 9 7 0 9 2 9 7 10 0 9 0 9 1 10 9 2 3 9 2
25 16 15 4 13 3 0 1 11 2 7 13 7 13 10 9 15 3 4 4 13 1 1 0 9 2
12 10 9 4 4 13 7 13 1 0 9 0 2
35 7 16 15 13 0 1 10 0 9 2 4 10 0 13 16 15 13 7 0 7 0 2 9 10 4 13 16 9 4 13 1 9 0 0 2
7 9 0 9 13 3 0 2
29 1 9 13 15 3 3 0 0 2 7 0 16 15 4 13 15 0 2 3 4 10 13 16 15 13 15 14 13 2
15 1 0 9 13 3 0 2 0 2 9 1 9 1 9 2
13 1 9 4 3 9 13 14 13 2 1 9 2 2
7 0 9 13 1 9 1 2
28 9 1 11 13 0 2 7 4 13 1 12 9 1 9 1 12 1 12 9 1 12 2 10 9 1 12 9 2
9 9 13 3 10 1 15 15 13 2
30 1 11 13 15 1 16 12 0 1 9 13 0 1 9 1 9 9 2 7 16 0 12 9 9 13 1 9 1 9 2
17 1 9 13 15 16 9 13 12 2 0 2 9 10 9 1 9 2
17 16 9 13 10 9 1 9 7 10 9 13 15 3 1 0 9 2
22 10 9 1 12 13 1 10 0 9 1 9 2 0 9 7 14 13 9 3 0 0 2
19 9 0 9 1 14 13 0 7 13 0 2 13 3 0 16 15 13 9 2
10 15 13 14 13 1 9 1 12 9 2
18 9 4 0 13 14 13 9 1 9 1 9 1 9 7 1 0 9 2
9 15 4 13 0 9 2 7 9 2
12 7 15 13 0 1 1 0 7 0 0 9 2
14 0 4 9 3 13 1 0 9 7 13 1 0 9 2
5 14 13 9 0 5
3 0 0 2
5 0 2 3 0 2
12 1 14 13 0 1 9 4 15 13 9 0 2
13 15 4 3 13 14 13 15 1 1 3 10 0 2
28 0 13 10 9 15 13 3 0 16 9 9 1 11 13 1 10 9 2 15 2 13 2 3 15 10 1 9 2
24 10 13 10 0 9 3 2 15 2 13 9 7 2 3 15 13 10 9 1 10 1 15 2 2
15 15 13 0 9 1 14 13 0 9 0 9 1 10 0 2
45 1 10 9 13 15 0 14 4 13 1 16 11 9 7 0 9 13 1 0 9 2 3 0 9 13 15 15 13 14 13 2 7 0 9 2 3 0 9 13 10 0 9 1 9 2
10 7 0 7 0 9 13 0 1 11 2
10 9 13 16 3 15 13 0 1 15 2
14 15 13 3 3 16 15 15 0 13 2 0 13 9 2
29 11 13 10 9 9 1 14 13 0 1 9 7 10 0 9 1 10 9 7 9 1 9 1 2 10 0 11 2 2
12 9 13 1 9 3 16 9 7 9 4 13 2
12 10 2 0 0 0 9 2 13 10 0 9 2
6 15 13 0 1 9 2
9 2 0 2 9 13 3 1 15 2
20 15 13 3 7 0 9 1 9 2 9 9 15 4 13 1 0 2 4 13 2
26 1 9 4 15 13 10 0 9 1 10 0 2 7 10 1 15 13 0 1 14 13 10 9 1 9 2
13 9 13 1 15 2 1 16 15 13 9 7 9 2
9 9 13 15 1 15 2 1 9 2
56 16 15 13 1 9 16 11 1 9 13 10 0 7 0 9 2 4 15 13 0 1 7 9 7 9 16 0 13 10 0 9 12 9 1 9 2 3 3 16 15 4 13 2 13 15 7 13 2 7 15 13 9 3 1 9 2
17 0 2 9 13 1 10 9 16 9 1 11 13 10 0 7 0 2
19 15 13 16 10 9 3 4 13 0 9 1 2 3 9 2 9 7 9 2
31 3 4 9 1 9 11 11 11 1 10 0 0 9 1 9 2 16 9 4 13 3 16 15 3 13 10 2 13 1 0 2
20 16 15 13 9 1 15 1 9 2 13 15 3 3 9 1 9 1 10 9 2
30 7 16 15 3 2 1 9 1 9 2 4 13 1 9 7 9 15 4 13 1 9 1 9 2 4 9 13 3 0 2
9 10 1 15 15 4 13 1 13 2
24 3 13 9 15 13 0 1 2 9 0 2 2 1 9 15 14 13 0 7 9 1 10 9 2
18 3 4 15 13 0 7 0 9 1 10 9 15 13 0 7 3 0 2
37 9 2 9 1 9 2 9 15 13 13 1 1 10 0 9 2 7 0 9 1 15 15 13 0 2 13 10 1 15 15 4 13 10 9 1 9 2
7 3 13 15 10 10 9 2
2 9 5
4 10 9 9 2
4 9 7 9 2
4 9 7 9 2
4 13 1 9 2
13 9 11 11 4 13 16 9 11 11 13 9 0 2
9 3 4 0 9 13 14 13 9 2
13 1 10 0 9 4 11 9 3 13 10 10 9 2
15 3 13 15 7 15 3 0 1 10 9 1 10 0 9 2
23 10 0 0 9 4 13 1 16 9 4 13 15 15 13 1 1 14 13 0 9 1 9 2
26 3 13 11 11 1 11 3 15 13 10 9 15 13 2 3 10 9 2 16 15 13 10 9 1 9 2
21 11 13 3 0 16 15 2 1 9 2 13 11 1 2 9 1 11 0 9 2 2
4 15 13 9 2
11 9 13 16 15 13 7 1 9 7 9 2
19 9 9 13 9 2 9 2 2 9 2 9 2 7 9 2 0 9 2 2
16 10 9 13 1 11 9 2 7 9 13 2 11 13 0 9 2
15 11 13 1 10 9 9 1 9 7 10 0 9 1 11 2
33 15 13 1 1 14 13 16 9 1 16 15 4 13 1 14 13 1 15 2 13 16 15 13 10 10 9 1 9 7 10 0 9 2
34 1 9 1 10 0 9 4 15 13 14 13 9 1 10 12 9 1 9 7 13 1 10 0 2 0 9 15 15 13 0 14 13 1 2
25 11 13 3 1 1 10 0 9 1 9 1 12 16 10 9 13 0 1 14 13 9 9 1 11 2
17 9 13 2 7 9 13 0 2 7 2 9 13 14 13 1 2 2
19 1 10 9 13 9 10 9 2 9 1 10 0 9 7 9 13 10 9 2
26 1 11 4 3 15 1 9 2 13 1 9 2 1 14 13 2 1 9 2 3 10 9 4 13 1 2
28 11 13 0 9 1 10 9 1 0 9 7 9 1 10 9 2 1 14 13 10 0 9 1 16 9 13 0 2
11 1 10 9 13 11 10 9 0 1 9 2
16 15 13 15 1 14 13 15 0 0 2 0 0 7 0 0 2
17 11 13 15 1 16 9 1 9 13 0 9 7 13 1 10 9 2
13 0 13 15 16 11 7 11 4 13 0 1 15 2
40 15 13 16 9 1 14 13 9 4 13 2 7 16 10 0 9 4 13 15 1 15 2 7 3 13 15 9 1 0 9 1 11 2 10 0 9 3 1 11 2
6 11 13 3 0 9 2
12 15 13 0 15 9 1 10 0 9 4 13 2
19 15 13 1 9 1 14 13 10 0 9 7 13 9 7 9 1 11 9 2
12 15 13 1 16 15 13 15 15 13 0 0 2
17 0 9 15 1 9 13 9 1 9 13 0 1 9 9 7 9 2
7 7 0 9 13 3 9 2
39 13 9 14 13 15 2 4 15 13 1 0 9 15 13 9 2 15 13 1 9 7 15 13 15 10 9 1 14 13 1 1 10 0 7 0 1 15 10 2
5 15 4 13 9 5
3 3 0 2
2 0 2
24 3 13 9 1 9 0 0 1 16 9 1 10 0 9 4 13 16 9 3 4 13 3 0 2
27 9 1 10 0 9 2 9 2 4 13 9 2 13 9 1 9 7 13 9 1 9 1 0 9 1 9 2
24 9 13 1 1 9 2 7 9 1 9 13 0 1 14 13 9 1 1 1 0 9 3 0 2
41 16 15 13 14 13 10 0 0 9 2 0 15 10 0 9 13 0 7 1 10 9 2 4 15 13 16 15 13 14 13 10 0 9 1 9 15 0 4 13 9 2
9 11 7 11 0 9 4 13 9 2
28 10 0 9 1 12 9 9 1 9 4 3 13 2 9 13 3 12 9 0 1 12 1 1 10 0 9 12 2
37 9 1 14 13 9 1 9 4 13 1 16 15 4 13 15 2 12 9 2 2 7 9 13 1 16 9 1 14 13 1 9 1 0 9 4 13 2
15 15 15 13 0 3 13 14 13 1 9 15 3 13 9 2
12 0 13 13 14 13 16 15 3 13 10 9 2
19 0 0 13 15 14 13 1 15 15 13 10 9 2 7 13 13 14 13 2
21 10 0 9 15 13 2 13 14 13 1 9 1 12 9 1 12 9 1 0 9 2
13 9 13 14 13 9 1 9 1 10 9 1 9 2
8 9 4 13 0 7 0 13 2
22 10 9 9 4 13 3 15 13 0 0 2 7 9 1 10 9 4 13 0 1 9 2
16 10 9 13 16 1 9 2 9 7 9 4 10 9 13 9 2
20 9 13 0 1 10 0 9 2 15 15 13 1 9 13 3 3 1 10 9 2
27 9 2 3 15 13 1 9 2 13 3 0 1 14 13 0 1 0 9 2 0 1 9 7 0 1 9 2
16 16 9 9 13 3 0 1 14 13 9 13 3 15 10 9 2
18 10 0 0 13 16 7 9 7 9 13 14 13 9 1 9 1 9 2
14 11 13 9 1 10 0 9 1 9 7 9 1 9 2
13 15 13 16 7 9 7 9 1 0 9 4 13 2
28 9 4 13 1 10 9 1 12 9 0 9 1 9 1 9 2 12 9 2 2 7 15 1 7 1 0 9 2
26 9 4 13 10 9 1 12 9 1 9 1 9 1 7 1 0 9 7 1 0 9 2 12 9 2 2
18 15 4 13 10 0 9 2 7 15 13 0 16 15 13 10 9 1 2
6 15 13 15 9 13 2
10 7 9 1 9 13 3 14 13 9 2
16 7 10 0 9 13 10 9 1 14 13 15 1 14 13 15 2
8 9 13 3 3 3 0 3 2
13 7 9 13 10 9 7 15 13 1 15 7 15 2
5 13 9 10 9 5
3 0 9 2
3 0 9 2
20 11 11 4 3 1 10 9 13 1 14 13 1 10 0 9 1 11 7 11 2
14 9 4 3 13 0 1 14 13 9 10 10 0 9 2
19 10 0 9 1 11 13 1 11 1 14 13 10 0 0 9 11 11 9 2
20 15 13 3 0 9 11 11 1 0 9 16 15 13 1 9 1 11 1 9 2
23 10 9 9 1 11 10 0 9 4 13 1 10 9 1 14 13 9 1 9 10 0 9 2
9 15 4 13 9 1 11 0 9 2
15 9 11 13 16 3 10 0 9 13 15 13 1 0 9 2
16 3 1 13 15 1 9 1 9 16 9 4 13 2 13 15 2
11 15 13 1 9 1 10 0 9 1 11 2
25 15 13 14 13 1 9 1 9 7 9 2 0 9 7 9 7 9 1 9 1 10 0 0 9 2
25 15 13 11 9 1 10 9 1 12 2 7 4 3 13 16 10 0 9 1 10 0 9 4 13 2
10 10 0 7 0 9 1 11 13 0 2
22 11 13 16 0 10 9 9 13 1 9 1 9 2 16 9 13 9 1 9 7 9 2
17 3 16 9 4 10 13 10 0 9 2 13 9 10 0 0 9 2
11 1 12 9 1 9 1 9 13 0 0 2
21 15 4 3 13 16 11 13 1 12 9 1 0 9 1 0 9 7 1 0 9 2
11 3 3 4 0 13 2 7 3 10 9 2
17 7 0 7 9 13 1 9 1 10 9 1 0 9 1 12 9 2
10 9 13 1 9 15 0 4 13 15 2
23 9 11 11 4 10 0 9 13 1 14 13 9 1 1 9 9 7 1 1 10 0 9 2
25 16 11 1 0 9 13 10 9 1 12 2 13 9 0 1 10 9 7 9 4 13 1 11 9 2
11 10 9 1 9 4 13 1 10 0 9 2
21 15 13 1 15 15 13 16 15 3 4 13 10 9 1 14 13 0 7 0 9 2
18 15 13 15 14 13 10 0 9 15 1 9 13 3 1 9 1 9 2
16 11 4 1 10 9 13 2 13 7 13 9 1 9 7 9 2
7 3 13 9 0 1 9 2
31 15 4 10 0 9 13 10 9 9 1 11 15 4 13 1 16 9 3 13 1 10 0 0 9 2 1 10 9 1 11 2
16 3 4 10 0 9 13 1 16 11 11 3 13 9 1 9 2
21 3 4 9 13 0 7 0 1 14 13 9 0 9 1 9 7 9 10 0 9 2
25 7 9 1 11 4 13 1 0 1 9 2 9 4 3 13 14 13 9 7 9 1 9 1 9 2
18 15 4 3 13 16 10 0 9 9 3 10 9 13 1 9 1 9 2
5 9 3 1 9 5
2 9 2
14 10 0 9 13 1 9 2 7 9 1 9 13 0 2
5 15 13 11 1 2
15 1 9 13 11 11 1 9 1 12 0 9 1 9 9 2
24 3 13 9 12 9 1 0 9 2 12 9 9 2 12 9 0 0 7 12 9 1 0 9 2
18 1 9 13 15 16 1 12 0 9 13 3 12 1 9 1 0 9 2
16 9 4 0 13 16 11 13 9 1 0 9 1 10 0 9 2
13 15 13 0 16 3 0 9 13 9 1 0 9 2
18 9 13 16 9 9 0 4 13 1 1 9 1 10 9 9 13 1 2
6 0 9 13 3 12 2
12 1 9 13 15 3 0 9 15 13 0 9 2
14 0 7 0 9 13 0 1 9 2 7 1 9 9 2
19 0 7 0 9 13 1 3 12 9 1 9 1 9 7 12 9 1 9 2
15 1 12 13 9 9 1 1 12 9 1 9 1 9 1 2
17 9 1 9 13 2 0 15 15 15 13 0 4 13 9 1 9 2
24 1 9 4 12 0 0 13 1 11 0 9 16 9 13 14 13 9 1 10 0 9 7 9 2
24 15 0 13 13 3 3 7 0 9 7 0 9 1 9 2 7 0 9 1 14 13 10 9 2
8 10 9 1 9 1 0 0 2
13 1 0 4 9 1 9 13 0 7 3 1 9 2
19 1 12 13 9 0 12 9 2 1 12 4 15 3 13 2 1 12 9 2
15 1 10 9 4 9 13 1 9 7 14 13 1 0 9 2
9 0 0 4 3 13 1 0 9 2
26 10 10 9 1 0 9 13 15 1 11 0 9 1 14 13 10 0 0 9 2 9 2 1 0 9 2
18 1 9 4 9 1 0 9 4 13 11 1 9 1 16 9 4 13 2
38 15 13 0 9 7 9 1 9 15 13 1 0 9 2 1 0 15 13 0 0 7 1 10 9 13 10 9 1 0 9 15 3 4 13 1 10 9 2
17 15 13 0 14 13 3 9 7 9 0 13 0 0 7 10 9 2
24 9 4 0 13 1 16 9 1 10 9 13 0 9 1 9 1 10 9 2 0 0 7 9 2
39 0 0 4 13 9 1 2 9 2 1 9 1 9 1 9 2 7 9 1 9 2 1 9 1 14 13 0 9 2 7 1 11 2 4 3 13 10 9 2
18 1 0 9 1 9 2 4 15 13 9 1 10 9 3 1 11 9 2
5 1 9 1 9 5
4 9 1 9 2
4 9 1 9 2
13 0 9 13 11 11 1 10 3 0 0 0 9 2
6 7 1 9 13 15 2
7 4 15 3 13 10 9 2
10 11 11 13 10 9 1 10 0 9 2
26 0 0 0 13 15 10 0 9 1 11 0 9 1 1 10 9 9 7 9 15 13 0 2 0 9 2
30 9 1 11 2 9 1 11 2 0 9 1 11 2 9 1 9 2 9 1 9 1 11 2 9 7 0 9 1 9 2
7 15 4 13 9 1 0 2
28 1 9 1 11 9 1 14 13 0 0 1 0 9 1 11 2 13 15 11 0 9 1 14 13 9 1 11 2
20 11 4 3 13 10 0 0 9 2 3 0 1 10 0 9 1 10 0 9 2
11 7 9 1 15 9 4 13 13 3 0 2
18 9 4 13 0 0 16 15 3 13 2 3 16 15 3 13 1 10 2
20 10 0 9 1 11 3 13 15 10 0 9 1 16 9 1 9 4 13 9 2
12 3 16 9 3 13 15 1 2 3 13 9 2
12 7 15 4 13 1 9 2 7 4 13 9 2
18 0 13 15 16 11 13 0 9 1 14 13 1 1 11 10 0 9 2
8 15 13 3 16 11 13 9 2
17 3 10 11 9 13 0 1 2 7 15 4 3 13 9 1 9 2
14 15 13 9 2 15 3 4 13 9 1 9 1 9 2
22 1 3 0 4 11 3 13 15 9 1 14 13 1 0 9 1 9 1 11 1 9 2
22 15 13 3 3 0 1 10 9 3 7 9 7 9 7 9 13 0 9 1 10 9 2
10 7 3 0 1 9 13 9 1 11 2
11 15 13 0 9 1 9 1 0 9 9 2
11 9 4 13 0 2 7 4 13 10 9 2
11 9 13 2 7 0 13 14 13 1 11 2
11 11 13 3 1 9 10 9 1 0 9 2
13 0 13 15 3 13 10 9 1 9 15 13 1 2
12 3 9 11 11 4 13 9 1 10 0 9 2
23 9 4 13 0 9 1 11 0 9 1 14 13 10 9 2 7 0 13 15 13 1 15 2
20 4 9 1 11 9 13 1 9 1 11 1 10 9 1 14 13 0 0 9 2
2 3 2
15 3 4 10 10 9 1 0 13 0 9 0 1 10 9 2
13 7 9 4 3 13 1 0 9 2 0 1 9 2
11 15 4 13 9 1 9 7 13 9 0 2
36 9 13 1 10 9 10 9 1 11 1 10 3 0 0 9 2 7 15 13 2 15 15 10 13 2 10 9 1 9 1 10 9 15 4 13 2
18 3 4 15 13 16 10 0 9 1 9 3 13 10 10 9 7 9 2
7 9 1 11 7 1 11 2
3 0 9 2
7 11 9 1 9 13 0 2
24 1 14 13 14 13 0 9 1 10 0 2 4 15 4 13 15 1 14 13 9 1 1 9 2
16 9 11 11 13 1 9 9 1 10 0 9 1 9 1 9 2
18 15 13 10 0 9 13 1 0 9 1 11 2 13 1 9 1 11 2
23 9 13 16 9 7 0 9 4 13 12 9 9 7 9 1 11 1 14 13 9 1 9 2
18 1 2 9 2 13 2 9 15 4 13 1 9 1 9 1 9 2 2
8 11 0 9 1 9 13 0 2
13 9 1 9 2 7 9 1 14 13 9 7 9 2
9 1 1 4 9 13 9 1 9 2
14 14 13 9 13 3 0 1 9 1 0 9 4 13 2
14 1 9 13 9 9 1 9 15 13 1 9 1 9 2
55 16 9 13 9 1 14 13 10 9 1 11 1 9 1 9 2 13 9 1 9 16 7 13 9 1 16 10 9 13 14 13 9 1 11 1 0 9 2 7 9 4 13 9 1 9 3 15 0 13 0 14 13 0 9 2
25 1 1 13 15 16 9 1 11 7 2 0 2 9 2 7 9 9 13 10 12 9 15 13 9 2
6 3 13 0 9 9 2
30 16 9 13 3 0 16 9 13 14 13 2 13 15 3 7 0 14 13 1 9 15 13 0 2 3 0 9 1 9 2
32 16 9 1 9 2 1 9 1 10 9 15 13 2 3 13 9 2 4 15 13 9 1 10 3 0 9 2 15 4 13 0 2
32 3 2 16 9 1 9 13 1 14 13 9 1 2 4 9 13 1 0 9 2 0 9 2 1 10 9 3 9 3 13 0 2
27 9 13 1 9 16 9 2 7 9 2 13 0 2 3 3 1 9 2 7 3 1 9 1 9 1 9 2
8 9 1 9 4 13 0 9 2
13 9 4 3 13 1 0 9 15 4 13 1 11 2
33 3 4 11 9 1 11 13 1 15 15 0 13 1 0 9 2 13 7 13 1 10 10 0 9 2 9 1 9 15 13 1 9 2
8 7 11 7 11 13 10 0 2
8 10 0 0 9 13 0 9 2
14 11 13 16 9 3 1 0 9 4 13 9 7 9 2
30 9 1 11 1 9 4 3 13 1 0 9 1 11 2 15 4 13 3 7 0 1 0 9 2 3 1 9 1 11 2
16 10 0 9 1 0 9 4 13 0 9 15 3 4 0 13 2
8 9 11 11 4 13 1 9 2
5 9 13 10 9 5
4 9 13 3 2
4 0 1 9 2
4 4 4 13 2
4 9 1 9 2
2 9 2
3 13 9 2
20 3 4 3 0 0 9 2 9 7 9 13 3 0 9 15 13 3 0 9 2
34 1 9 13 0 9 1 9 3 12 7 12 9 2 16 9 2 1 11 11 2 13 10 0 9 15 13 0 9 2 13 11 11 11 2
3 0 9 2
6 0 9 13 0 9 2
10 7 9 1 0 9 13 3 0 9 2
34 9 15 3 13 9 1 10 9 2 13 14 13 0 9 15 13 3 0 1 9 1 9 2 9 7 9 16 9 13 9 1 14 13 2
9 16 9 3 13 2 13 10 9 2
17 7 15 13 10 9 15 3 13 0 1 1 0 1 9 1 9 2
29 3 4 9 13 16 11 11 13 3 0 2 7 16 0 9 4 13 0 2 0 1 11 11 9 1 11 0 9 2
12 1 12 9 3 13 9 10 0 9 1 11 2
34 11 11 7 11 11 2 11 11 7 11 11 13 9 15 13 7 13 0 1 2 15 13 9 2 15 4 13 1 0 7 1 0 9 2
23 9 4 13 0 3 2 1 9 1 0 9 7 1 14 13 9 1 10 0 9 1 9 2
12 13 10 1 9 0 9 1 14 13 10 9 2
7 3 13 15 3 1 9 2
16 9 4 3 13 0 9 16 15 3 13 15 13 0 1 15 2
5 7 15 13 15 2
24 7 3 16 9 3 3 13 1 1 9 2 13 9 3 10 9 1 9 15 13 1 1 9 2
6 1 9 13 3 0 2
10 15 13 3 16 15 3 13 0 9 2
24 11 11 2 11 11 11 2 11 11 2 0 0 9 2 15 13 3 15 15 13 9 7 9 2
15 15 13 0 1 9 2 7 15 13 15 10 0 0 9 2
20 11 2 15 13 1 12 2 13 3 1 0 1 11 16 9 1 9 4 13 2
11 15 13 0 2 7 9 13 0 1 9 2
4 9 13 0 2
24 0 9 2 0 9 2 0 9 13 0 2 7 15 13 11 11 11 2 11 11 7 11 11 2
24 15 4 13 1 9 2 15 3 3 4 13 9 2 7 15 4 13 10 9 1 14 13 9 2
13 10 2 15 2 4 3 1 10 9 13 1 9 2
28 10 2 15 2 13 1 10 9 14 13 15 14 13 1 10 0 9 1 9 2 1 9 2 1 9 7 9 2
23 9 1 9 4 0 3 13 15 2 7 1 10 9 15 3 4 13 15 3 0 1 9 2
8 15 13 10 10 1 10 9 2
13 1 9 13 0 9 1 9 3 12 7 12 9 2
15 9 13 3 1 1 9 2 9 13 3 1 2 9 2 2
43 16 0 9 13 9 7 9 4 13 0 0 2 7 1 9 13 9 2 9 2 15 15 13 9 7 3 13 9 2 13 9 1 3 14 13 16 3 9 7 9 13 0 2
22 2 4 10 0 1 0 9 13 16 9 13 9 1 9 1 14 13 10 0 9 2 2
17 3 13 15 0 16 15 13 9 1 9 15 1 0 9 13 15 2
5 10 9 13 9 2
33 0 9 15 4 13 0 9 1 10 9 0 1 9 7 9 2 13 10 0 9 15 13 0 9 1 9 15 13 10 9 1 9 2
16 11 11 2 11 11 2 11 11 7 11 11 4 13 1 9 2
27 3 13 10 0 9 1 9 1 9 7 10 9 7 9 2 7 1 14 13 9 1 10 0 9 1 9 2
23 10 0 9 13 0 3 0 2 15 13 10 9 1 9 1 11 7 11 2 11 7 11 2
16 7 9 4 13 1 9 1 10 2 0 3 3 0 2 9 2
46 0 13 15 0 9 1 0 9 1 9 15 1 9 13 9 15 4 13 2 3 2 1 9 2 7 1 15 15 1 9 13 9 7 9 15 4 13 1 10 10 9 9 15 13 15 2
34 1 1 9 4 9 1 0 9 13 9 1 0 9 2 1 9 2 1 9 7 9 2 7 3 1 9 1 10 9 1 9 7 9 2
29 2 9 2 13 1 10 9 0 3 2 0 9 2 2 15 13 0 10 15 1 2 10 0 0 9 1 9 2 2
23 15 13 10 0 9 16 10 9 13 1 16 9 1 9 7 9 3 13 3 0 1 15 2
25 9 13 15 13 1 9 2 7 9 13 3 9 9 0 2 15 13 15 2 7 9 13 10 9 2
14 1 9 4 9 1 9 13 10 10 9 1 10 9 2
15 1 9 9 4 9 9 13 3 0 0 1 0 9 9 2
18 15 13 1 0 9 9 2 9 2 7 15 15 0 0 4 13 9 2
25 9 1 0 9 4 3 3 4 13 15 0 2 1 10 9 3 9 0 9 1 0 9 13 0 2
45 16 1 10 9 15 3 13 15 0 1 9 2 7 1 0 9 13 15 1 10 9 0 1 9 2 9 2 9 2 9 1 10 9 2 13 0 9 15 1 0 9 13 14 13 2
7 15 13 3 15 13 0 2
11 9 13 3 3 16 9 13 0 7 0 2
24 7 0 3 16 0 9 4 13 1 10 0 9 3 2 7 1 16 9 0 13 9 0 9 2
5 3 4 9 13 2
19 9 4 13 9 1 3 14 13 15 1 9 2 13 15 15 3 13 10 2
17 10 0 7 0 9 1 11 1 9 4 3 13 1 0 0 9 2
17 7 3 3 9 2 9 7 9 4 13 1 0 9 1 0 9 2
15 7 15 13 0 3 10 9 16 10 9 4 13 1 15 2
22 7 15 13 0 2 7 0 2 16 0 9 4 13 9 1 14 13 10 0 0 9 2
6 15 13 10 0 9 2
10 0 2 9 2 4 13 0 1 9 2
19 7 9 4 3 13 2 7 7 9 7 10 10 4 13 9 10 0 9 2
13 7 10 9 14 13 9 13 2 13 10 9 2 2
17 15 13 0 3 1 14 13 10 0 9 2 7 9 13 3 0 2
30 7 4 0 1 10 0 9 15 13 0 9 2 13 0 1 1 9 2 1 9 7 9 2 7 9 2 9 7 9 2
20 4 10 0 1 0 9 13 16 9 13 9 1 9 1 14 13 10 0 9 2
13 2 8 8 8 2 8 8 8 8 8 8 2 2
25 1 9 13 9 16 3 4 3 0 0 9 2 9 7 9 13 3 0 9 15 13 3 0 9 2
6 14 13 13 14 13 5
3 0 9 2
4 9 7 9 2
2 9 2
2 9 2
4 10 0 9 2
3 9 9 2
5 1 9 1 9 2
3 0 9 2
10 11 11 13 3 0 9 13 9 9 2
21 11 11 4 13 16 9 13 1 15 15 15 13 9 1 10 9 2 13 11 11 2
6 14 13 13 14 13 2
9 10 9 4 13 1 9 11 11 2
33 1 10 0 0 9 7 9 1 9 0 11 13 11 0 10 9 2 7 15 13 1 1 9 9 7 13 0 1 0 9 1 11 2
19 7 15 13 16 15 2 12 9 3 0 2 13 16 15 10 4 13 11 2
16 14 13 13 14 13 2 10 9 4 3 13 1 11 11 9 2
19 9 9 1 9 4 1 9 0 13 16 15 3 4 13 1 14 13 9 2
20 9 13 1 15 10 9 2 10 9 1 10 0 0 9 9 1 14 13 15 2
35 10 0 9 2 15 13 9 1 9 7 9 2 4 3 13 1 10 0 9 1 14 13 1 9 9 9 1 14 13 3 3 1 14 13 2
11 11 11 13 10 0 9 1 9 0 9 2
20 10 0 9 1 1 1 16 15 3 13 9 1 14 13 2 0 1 14 13 2
9 9 10 13 0 2 0 2 0 2
13 15 13 0 9 7 0 0 9 3 1 11 11 2
15 9 7 9 13 3 9 10 2 7 15 13 3 10 9 2
15 9 13 15 1 10 0 9 7 13 1 9 7 0 9 2
21 15 13 1 10 9 1 9 9 2 9 9 2 9 9 2 9 9 7 9 9 2
14 10 0 9 1 0 9 2 9 7 9 13 11 11 2
31 15 13 1 10 0 2 7 0 9 2 1 9 4 15 13 0 2 13 14 13 2 13 2 13 2 13 2 13 2 13 2
20 10 9 13 0 9 2 3 1 10 9 7 9 2 3 1 10 9 7 9 2
28 13 1 12 1 10 0 9 1 11 1 1 11 13 15 1 1 10 0 9 15 13 10 1 9 0 0 9 2
29 15 4 13 0 9 1 9 7 13 10 9 0 9 1 10 9 0 0 9 15 1 9 1 10 0 9 13 9 2
26 1 9 13 15 1 9 1 10 9 2 7 13 9 16 15 13 14 13 1 10 0 9 7 13 9 2
10 3 4 15 1 0 9 13 1 11 2
18 9 13 1 12 1 10 9 15 4 0 13 1 9 16 15 4 13 2
30 1 10 0 9 10 13 15 9 1 10 0 9 2 1 10 9 2 9 7 9 2 10 9 7 9 15 15 13 3 2
12 3 13 0 9 7 0 9 1 10 0 9 2
16 11 11 13 0 9 1 0 9 2 0 4 15 13 1 11 2
22 16 15 0 13 9 1 11 2 4 15 13 9 2 7 1 12 4 15 13 1 11 2
15 1 10 0 9 4 11 11 3 13 1 14 13 10 9 2
24 9 10 13 0 1 9 1 14 13 1 7 9 1 9 2 15 0 13 15 15 13 1 9 2
18 15 13 0 7 0 1 10 0 9 7 10 0 9 15 13 1 11 2
21 15 13 10 9 1 9 7 9 1 10 0 9 15 15 13 1 10 0 0 9 2
36 9 13 0 7 0 0 2 15 13 1 9 2 7 15 13 3 11 11 13 15 2 0 2 0 2 0 1 9 15 7 13 0 7 9 0 2
9 15 13 1 10 0 0 2 0 2
26 1 4 15 3 13 0 0 2 10 0 9 7 10 0 9 13 3 10 9 14 13 10 0 9 1 2
25 1 15 13 15 10 0 9 2 1 0 9 16 15 13 9 15 13 15 1 14 13 0 7 0 2
31 15 15 13 1 11 11 2 13 16 15 1 9 10 3 13 1 10 0 2 3 13 1 9 7 3 13 1 10 0 9 2
10 15 13 10 9 16 15 13 9 9 2
23 1 10 3 0 0 9 2 10 3 0 9 11 2 11 11 11 2 2 13 15 9 9 2
39 1 11 0 9 9 1 11 1 12 4 10 9 7 9 1 12 7 12 9 1 10 0 9 13 1 11 2 16 15 4 13 1 14 4 13 1 11 9 2
9 9 13 12 9 1 10 0 9 2
25 15 13 1 9 1 11 11 2 3 15 0 9 1 9 2 16 9 13 15 1 14 13 1 9 2
16 11 4 13 15 1 10 1 10 9 1 11 1 12 7 12 2
16 15 13 3 3 2 7 11 11 13 1 11 7 10 9 9 2
12 1 12 13 11 2 7 9 13 3 1 9 2
8 15 13 11 1 9 1 9 2
26 11 11 13 15 9 9 1 14 13 0 9 7 13 2 1 9 1 9 2 3 1 10 0 0 9 2
15 0 7 1 14 13 13 15 1 9 10 1 10 9 9 2
38 15 13 3 1 10 0 9 1 3 15 1 9 2 0 1 9 7 0 1 16 10 0 9 4 13 2 1 9 13 1 14 13 9 1 10 0 9 2
18 7 9 13 3 1 14 13 9 1 9 2 3 1 14 13 9 1 2
13 1 9 2 12 9 0 2 13 10 0 9 9 2
26 3 13 15 15 0 16 1 10 9 15 4 13 1 11 11 2 13 15 3 10 9 1 10 9 9 2
26 15 15 7 10 9 9 1 11 4 13 1 1 1 9 2 13 3 1 9 2 3 1 9 2 0 2
9 4 15 4 13 0 9 1 15 2
13 7 13 15 15 15 3 4 13 0 0 1 9 2
23 2 9 4 1 10 9 13 1 11 2 2 13 11 0 9 0 1 10 9 1 11 11 2
16 15 13 3 0 2 1 16 15 4 13 9 1 10 0 9 2
21 7 11 13 1 0 0 7 0 0 9 2 15 4 13 1 14 13 2 9 2 2
21 11 11 11 11 2 16 9 1 11 13 2 4 13 1 1 9 1 10 0 9 2
6 10 9 13 3 0 2
8 10 0 13 9 0 0 9 2
9 9 1 0 9 13 1 10 9 2
35 11 11 4 13 16 10 9 13 10 9 1 14 13 3 0 9 13 9 9 7 14 13 16 9 13 1 15 15 15 13 9 1 10 9 2
32 1 10 9 13 15 0 16 10 9 1 9 7 10 9 9 1 11 13 3 0 9 1 9 13 1 9 9 1 11 1 9 2
11 3 13 15 0 14 13 1 11 11 9 2
5 4 15 4 13 2
4 9 1 9 2
4 13 1 9 2
5 13 15 1 11 2
4 4 13 3 2
5 9 9 1 9 2
18 11 4 3 3 13 9 9 2 9 4 13 10 0 9 1 9 9 2
29 1 9 13 3 11 3 10 0 9 1 15 16 15 13 9 2 7 15 4 3 3 13 0 0 2 13 11 11 2
5 1 9 1 11 2
17 10 9 15 11 13 9 2 13 15 1 1 10 0 9 1 11 2
18 9 13 10 9 1 9 11 11 1 9 2 15 13 1 9 1 9 2
13 1 11 13 15 9 1 15 1 9 7 1 9 2
5 9 13 10 9 2
34 11 9 13 1 11 2 10 0 9 2 2 0 1 1 11 2 15 13 11 12 9 2 16 9 13 1 9 1 14 13 9 0 9 2
22 9 13 12 9 9 1 10 9 15 13 10 0 1 9 2 10 9 1 9 1 11 2
23 9 13 12 9 2 10 0 1 9 2 7 15 13 0 1 12 0 9 7 3 0 0 2
4 9 13 0 2
27 10 0 9 1 12 9 1 9 0 9 2 9 1 4 0 12 13 1 10 9 1 10 1 9 1 9 2
25 10 0 9 1 9 13 9 1 15 9 4 13 1 1 9 1 9 7 9 2 9 1 0 9 2
9 11 13 3 0 1 9 7 9 2
6 9 12 13 1 12 2
25 15 13 10 9 1 0 9 1 11 2 7 13 1 9 14 13 12 9 1 9 1 11 1 12 2
13 11 13 1 10 0 9 15 4 13 2 1 12 2
14 1 9 13 12 1 0 9 7 12 1 10 12 9 2
10 16 15 13 9 2 4 13 1 0 2
9 1 10 9 1 9 13 11 9 2
17 15 13 9 1 10 0 9 2 15 4 13 12 9 9 1 9 2
8 0 9 4 13 0 9 12 2
17 1 9 13 9 12 9 2 7 1 9 1 12 4 9 13 0 2
15 3 13 15 9 2 9 7 9 1 12 9 7 12 0 2
28 3 3 13 15 1 9 9 1 9 1 10 0 9 2 12 0 9 2 12 9 2 12 9 7 10 0 9 2
21 9 13 0 7 0 2 1 9 2 12 0 9 2 1 10 1 15 10 0 9 2
10 9 15 13 15 1 2 13 0 0 2
18 2 15 13 15 2 9 2 13 15 2 16 15 13 16 15 13 3 2
22 2 4 11 13 9 7 13 14 13 10 1 10 9 15 1 15 3 13 1 9 2 2
14 0 9 1 9 7 9 13 1 0 0 9 1 9 2
9 11 13 0 1 14 13 10 9 2
9 15 13 10 9 1 10 0 9 2
12 0 9 13 1 0 9 2 10 10 13 9 2
11 9 1 9 1 9 13 0 1 0 9 2
19 10 0 9 13 15 3 16 15 13 1 14 4 13 9 0 1 1 11 2
26 10 0 9 1 9 13 0 0 2 7 4 13 10 9 1 9 1 9 1 16 15 13 15 11 13 2
26 15 13 3 3 2 7 3 13 15 1 9 1 9 10 7 13 11 1 0 0 9 2 7 13 0 2
6 2 13 15 1 11 2
23 1 10 0 9 1 15 2 13 15 0 10 0 9 1 9 2 7 9 13 1 1 9 2
18 1 11 13 9 1 9 15 15 15 13 1 9 1 10 9 1 9 2
25 1 9 13 3 11 3 10 0 9 1 15 16 15 13 9 2 7 15 4 3 3 13 0 0 2
14 10 9 13 9 2 3 3 1 14 13 9 0 9 2
30 10 9 13 15 15 12 9 14 13 2 16 9 0 9 13 0 0 1 9 1 12 2 7 1 1 0 1 10 9 2
11 15 4 15 1 11 13 0 1 12 9 2
20 15 4 13 0 1 0 9 2 15 4 13 1 0 9 7 0 9 3 1 2
11 7 3 4 9 1 10 9 13 1 9 2
32 11 9 1 9 7 0 9 13 16 15 3 4 13 14 13 1 15 14 13 9 9 2 15 4 13 10 0 9 1 9 9 2
9 9 1 9 1 11 13 3 0 2
6 10 9 13 0 0 2
11 11 13 1 2 9 2 1 9 1 9 2
30 15 13 0 1 15 3 1 10 0 9 2 15 1 10 9 10 9 13 13 1 11 2 2 14 13 1 1 15 15 2
44 4 15 3 13 0 1 1 9 1 10 9 3 16 15 3 4 13 16 15 13 1 1 2 7 4 15 13 9 7 13 14 13 10 1 10 9 15 1 15 3 13 1 9 2
16 3 13 10 9 15 13 1 1 9 9 2 3 10 0 9 2
12 15 4 1 0 9 13 10 9 9 1 9 2
27 7 0 13 15 10 9 1 10 9 1 14 13 11 1 10 0 9 1 9 1 14 13 9 7 9 1 2
19 15 13 3 1 9 1 10 9 1 9 9 1 14 13 3 0 9 9 2
15 15 13 3 9 1 9 1 9 2 9 1 9 7 9 2
12 9 13 0 2 7 13 0 9 1 0 9 2
33 7 11 13 3 3 10 9 16 1 10 9 7 10 0 9 1 0 9 2 4 15 13 1 14 13 15 1 10 0 9 1 9 2
10 15 13 3 0 16 9 1 9 13 2
11 10 9 4 13 10 0 9 1 1 15 2
14 11 2 11 7 11 4 10 13 9 1 1 10 9 2
13 9 7 9 4 13 1 10 9 15 4 13 1 2
7 13 11 15 1 12 9 2
25 15 13 0 15 3 4 13 0 3 1 10 10 0 9 15 4 13 9 1 10 9 1 9 9 2
4 9 1 11 5
4 9 7 9 2
2 9 2
4 9 7 9 2
4 0 0 9 2
2 11 2
3 0 9 2
2 9 2
3 0 9 2
17 11 9 13 0 9 15 0 9 0 13 1 9 1 10 0 9 2
17 11 11 11 4 13 0 1 10 9 1 11 10 0 9 1 12 2
8 11 11 13 12 0 1 9 2
14 15 13 15 1 10 9 7 4 3 4 13 1 9 2
8 15 13 16 9 9 13 0 2
35 1 16 11 13 9 2 11 1 10 0 2 0 9 2 4 12 9 13 15 1 1 9 2 13 9 1 9 1 9 1 11 11 11 2 2
15 11 4 13 0 1 10 9 1 11 10 0 9 1 12 2
6 15 4 13 10 9 2
6 15 4 13 10 9 2
8 11 11 13 12 0 1 9 2
14 15 13 15 1 10 9 7 4 3 4 13 1 9 2
19 9 2 15 4 13 1 11 9 2 13 10 9 1 9 9 1 0 9 2
32 15 13 16 0 9 4 13 10 0 9 1 14 13 11 13 1 9 1 11 2 7 16 15 4 4 4 13 1 9 1 3 2
10 1 1 9 13 15 12 9 1 9 2
18 15 13 15 2 1 15 2 13 10 9 1 10 0 9 1 0 9 2
20 11 1 2 0 9 2 13 3 0 9 1 10 2 7 4 3 13 15 3 2
7 9 7 9 13 3 3 2
20 9 1 9 1 11 13 3 1 10 9 1 1 9 1 9 10 2 9 2 2
28 15 4 0 13 11 12 2 12 2 2 7 9 1 15 4 1 13 1 9 11 11 11 1 10 9 1 9 2
18 9 13 0 9 1 3 11 4 13 10 0 9 1 0 7 0 9 2
20 15 13 16 11 13 10 0 0 9 2 7 10 0 9 7 9 1 0 9 2
23 10 9 1 15 4 13 11 9 1 9 1 14 13 1 10 0 9 1 9 2 9 2 2
13 2 9 13 16 9 3 4 13 1 1 10 9 2
43 1 9 1 0 9 2 0 9 2 0 9 2 0 9 1 0 9 1 1 2 13 11 1 10 0 9 1 9 15 13 1 16 0 12 9 13 9 1 11 1 9 2 2
25 15 13 3 9 7 9 2 3 11 2 11 2 2 15 13 14 13 10 9 15 13 1 10 9 2
22 1 10 4 10 0 0 9 1 11 13 14 13 9 1 10 0 9 1 11 1 11 2
27 15 13 10 9 15 7 13 9 9 7 16 15 4 13 1 0 9 1 0 2 1 9 1 9 7 9 2
38 10 0 9 0 9 1 11 2 3 10 1 11 0 9 1 0 2 0 7 0 9 13 2 13 3 3 1 16 15 13 0 9 1 0 9 1 9 2
13 16 0 9 3 13 10 0 2 13 1 15 0 2
24 11 13 1 9 10 0 9 1 9 1 10 0 0 2 16 15 13 9 7 9 1 14 13 2
23 0 7 0 9 4 13 15 1 10 9 2 16 0 9 13 0 0 1 0 7 10 9 2
25 0 9 0 9 1 10 9 13 0 16 11 9 13 0 9 9 0 13 1 9 1 10 0 9 2
30 14 13 15 1 9 1 9 9 13 0 9 1 15 9 13 7 1 9 15 1 4 13 9 1 10 10 2 9 2 2
16 1 0 9 2 13 3 9 1 0 9 2 0 9 7 9 2
14 3 3 10 0 9 2 9 2 4 13 1 10 9 2
32 15 4 13 1 9 1 0 9 15 2 1 9 1 15 2 1 9 13 16 0 9 3 13 15 1 15 0 9 13 1 9 2
49 16 15 1 11 9 13 16 2 15 4 13 15 7 3 4 13 0 2 1 10 0 9 1 15 2 7 3 3 11 9 1 0 9 4 4 13 2 3 13 0 1 9 1 10 9 1 15 10 2
21 10 0 9 4 1 10 0 13 14 13 15 0 9 1 0 7 0 9 7 9 2
45 11 11 11 2 11 9 1 11 11 5 9 1 10 0 9 1 11 7 11 9 1 11 2 2 13 9 0 1 9 13 0 7 0 1 0 9 1 10 9 15 13 1 10 9 2
18 11 13 10 9 1 15 10 0 13 2 0 2 1 3 12 9 3 2
35 10 9 13 16 9 13 0 16 15 0 13 9 1 14 13 9 7 0 9 2 7 15 13 9 1 3 15 0 4 13 1 1 10 9 2
28 15 4 3 13 0 1 16 9 9 1 10 9 13 0 9 5 9 7 16 15 13 0 9 15 13 1 9 2
25 7 11 0 9 2 9 7 9 15 1 13 1 9 1 11 9 1 9 0 1 9 2 13 0 2
27 10 9 15 4 13 1 0 9 1 0 9 1 11 3 2 13 16 9 1 9 3 13 0 1 0 9 2
23 1 0 4 3 9 3 13 1 9 2 0 9 7 9 1 9 1 9 2 7 1 9 2
10 1 0 0 9 7 9 13 15 0 2
10 10 9 1 15 4 10 0 9 13 2
40 1 10 9 1 10 0 9 1 12 9 3 13 10 0 9 9 1 14 13 9 1 10 9 2 3 13 10 0 9 1 1 9 7 13 15 14 13 1 15 2
22 10 9 13 1 9 9 1 11 2 7 13 1 0 9 1 11 1 14 13 11 9 2
14 0 10 9 1 9 13 11 10 9 1 0 0 9 2
4 9 7 9 2
17 9 15 13 9 1 9 3 1 9 2 1 9 2 9 7 9 2
31 1 10 0 9 1 10 4 15 3 13 1 12 2 9 2 2 12 1 9 1 9 1 0 9 2 7 12 1 10 10 2
20 16 12 0 2 1 0 9 2 4 13 15 9 7 9 13 0 9 7 9 2
26 11 13 0 0 0 7 0 9 1 10 9 2 7 1 0 13 10 9 10 9 1 0 9 0 9 2
8 2 15 4 13 9 1 9 5
4 0 1 9 2
2 0 5
4 13 9 1 2
5 15 13 12 9 2
3 1 9 2
4 4 13 1 2
17 15 4 13 9 1 9 15 4 13 1 9 1 11 2 1 9 2
10 15 4 13 1 16 15 4 13 9 2
5 11 13 1 9 2
6 2 13 9 7 9 5
3 0 9 2
6 13 15 13 15 11 2
7 15 13 0 9 1 9 2
17 3 13 15 15 12 2 7 15 13 3 1 10 0 9 1 11 2
20 15 13 0 0 2 13 15 1 9 1 10 9 7 4 13 1 9 7 9 2
4 11 13 0 2
19 1 10 9 9 3 4 15 13 1 16 9 3 4 13 1 9 15 13 2
8 15 13 7 13 16 15 13 2
17 9 13 0 0 1 10 9 15 3 4 13 2 7 9 13 0 2
9 7 3 4 15 13 9 1 9 2
8 15 13 0 1 14 13 15 2
16 15 13 0 1 16 15 13 10 9 0 1 9 15 13 9 2
14 15 13 3 10 12 9 1 9 2 7 1 0 9 2
7 15 13 3 15 15 13 2
4 15 13 0 2
9 15 13 10 1 15 4 13 0 2
6 13 15 13 15 11 2
5 15 13 11 9 2
8 15 13 0 2 13 0 9 2
10 10 9 13 15 1 2 0 0 2 2
21 11 13 0 2 7 3 11 13 16 9 13 1 0 9 1 10 9 15 13 1 2
7 11 13 10 0 0 9 2
18 3 15 13 3 9 13 0 1 10 9 15 3 4 13 1 10 9 2
10 10 1 15 13 0 2 0 9 2 2
21 11 13 9 7 9 7 1 0 9 4 15 13 1 14 4 13 10 9 1 9 2
12 15 4 13 9 2 15 13 10 0 9 9 2
6 15 13 9 1 11 2
24 1 9 13 15 15 16 15 4 13 12 0 9 2 15 1 10 9 7 15 1 10 0 9 2
5 15 13 10 9 2
4 9 1 0 2
25 11 13 3 13 9 1 0 2 7 15 13 1 9 10 9 1 10 9 15 13 0 1 0 9 2
17 9 13 2 13 11 2 16 9 4 13 15 0 9 9 1 9 2
14 15 13 1 10 0 9 2 7 15 4 15 3 13 2
4 11 13 0 2
11 15 13 9 1 7 11 7 11 1 0 2
10 15 13 10 9 9 1 11 7 13 2
6 3 13 15 10 0 2
5 3 13 0 9 2
7 15 13 0 7 0 9 2
9 1 9 13 15 10 9 7 13 2
18 2 12 2 13 15 15 3 1 9 15 0 13 9 1 9 1 9 2
23 2 12 2 4 15 13 2 15 11 13 2 16 10 9 4 13 15 0 9 9 1 9 2
6 9 13 0 7 0 2
10 2 12 2 9 1 15 4 13 9 2
7 15 4 3 13 15 0 2
14 2 12 2 15 13 3 9 1 15 15 4 4 13 2
2 0 2
16 15 13 7 13 10 9 2 10 9 1 9 15 13 1 9 2
10 2 15 11 13 13 0 2 13 15 2
25 15 13 3 0 9 1 15 2 7 16 15 13 1 9 13 15 15 1 1 10 0 11 0 9 2
15 1 12 4 15 13 0 9 2 0 9 2 1 12 9 2
11 15 13 3 15 13 2 10 9 7 9 2
10 7 11 7 11 13 1 10 0 9 2
27 11 13 1 10 0 9 1 14 13 9 1 15 15 13 1 10 0 0 9 1 10 9 15 13 10 9 2
27 11 13 10 0 1 10 9 1 14 13 9 1 10 9 1 10 9 15 1 9 4 13 0 1 0 9 2
19 15 4 13 0 9 1 0 9 2 7 1 9 13 3 9 0 1 15 2
11 3 13 10 0 1 11 0 1 10 9 2
18 15 3 4 13 16 1 10 9 12 9 1 9 13 10 9 1 9 2
4 13 15 0 2
4 13 15 0 2
17 0 0 13 15 14 13 16 15 13 9 1 2 15 13 0 0 2
12 7 4 15 3 13 16 11 7 11 4 13 2
19 4 15 3 13 16 9 3 13 0 9 1 9 1 0 9 7 11 9 2
10 15 4 13 15 1 1 10 0 9 2
23 10 0 9 9 13 9 1 9 1 9 1 9 2 1 9 7 9 2 7 1 0 9 2
6 15 13 3 10 9 2
12 7 10 0 4 13 16 10 9 3 4 13 2
30 9 13 1 9 1 0 9 2 7 11 2 11 7 11 13 1 10 9 3 9 13 1 9 4 13 1 10 0 9 2
5 15 4 13 9 2
17 15 4 13 9 1 9 15 4 13 1 9 1 11 2 1 9 2
22 15 4 13 1 16 15 4 13 9 2 7 1 10 9 1 11 0 9 13 15 3 2
12 2 12 2 9 13 14 13 0 9 1 9 2
28 2 12 2 10 0 9 13 0 9 1 10 0 0 9 2 7 13 1 14 13 10 0 0 0 9 15 13 2
41 2 12 2 1 9 13 10 0 0 0 9 0 9 2 15 3 3 13 16 15 13 15 15 13 0 0 1 14 13 9 2 7 3 13 15 0 9 1 9 2 2
11 2 12 2 10 0 9 13 3 1 15 2
15 15 15 13 3 13 0 9 1 0 9 1 9 7 9 2
20 1 0 9 13 15 3 0 9 2 1 10 0 0 9 1 10 0 9 11 2
7 15 13 1 9 1 9 2
10 15 13 15 4 13 1 9 7 9 2
19 3 13 15 10 0 9 7 0 0 9 1 9 15 3 13 3 3 0 2
8 15 13 10 9 14 13 9 2
5 15 13 3 0 2
9 10 10 9 13 15 3 1 9 2
23 15 13 15 16 15 1 12 2 12 9 4 13 7 0 9 7 9 13 1 9 1 9 2
5 10 9 13 0 2
13 7 7 9 7 9 4 2 1 9 2 13 0 2
11 9 4 13 0 2 15 4 13 0 9 2
10 10 10 9 4 3 13 9 1 9 2
14 0 4 3 9 13 14 13 0 9 1 9 7 9 2
19 3 4 15 3 13 10 0 9 2 7 15 4 13 0 0 1 1 9 2
11 3 4 15 13 10 0 9 13 1 9 2
6 3 4 15 13 9 2
6 15 13 10 0 9 2
13 1 0 9 4 10 0 9 7 9 13 15 3 2
10 15 4 13 9 11 1 14 13 1 2
7 11 7 11 13 3 3 2
15 10 0 9 4 15 13 9 1 7 13 0 9 1 9 2
19 1 15 13 15 15 13 2 0 9 2 10 9 1 9 1 9 1 9 2
17 7 0 16 15 13 2 4 13 1 0 9 7 13 16 9 13 2
3 1 9 2
11 11 11 4 13 1 14 13 10 0 9 2
9 15 4 3 13 1 9 1 9 2
9 15 4 13 0 1 10 0 9 2
14 15 4 13 10 0 9 14 13 1 7 11 7 11 2
6 15 4 3 13 9 2
51 1 9 1 9 13 9 11 9 1 3 15 4 13 0 9 1 9 1 0 9 2 1 14 13 9 1 10 0 2 0 9 1 10 9 1 1 0 9 9 9 2 1 10 9 1 10 0 0 11 9 2
27 10 9 15 13 0 2 3 1 16 9 4 13 1 9 2 13 9 1 3 15 4 13 14 13 10 9 2
38 15 13 0 0 9 2 0 1 10 0 0 9 2 1 14 13 9 0 1 9 2 7 15 13 1 10 3 0 1 9 7 9 13 1 9 1 9 2
20 7 12 9 13 16 15 13 0 14 13 10 0 9 1 9 0 9 1 11 2
24 16 11 2 11 7 11 13 0 0 0 9 1 9 1 11 2 13 3 0 10 0 9 13 2
6 15 13 3 3 0 2
18 11 13 0 0 9 7 9 1 0 9 3 11 2 11 7 11 13 2
26 9 7 9 1 9 7 9 1 11 13 3 14 13 3 9 1 9 1 2 8 8 8 8 8 2 2
40 15 13 3 16 15 0 13 10 9 1 16 15 13 9 15 4 13 10 0 9 1 9 2 1 1 0 10 9 2 7 16 15 1 9 13 1 15 15 13 2
32 11 13 3 0 9 9 9 1 0 2 0 2 9 2 7 0 9 1 0 9 2 9 7 9 15 13 0 9 1 0 9 2
19 15 13 15 0 14 13 9 1 0 9 1 11 13 1 1 0 10 9 2
17 9 13 1 11 2 15 15 13 10 9 1 16 9 1 9 13 2
5 7 9 7 9 2
37 15 13 3 3 16 7 10 0 7 0 9 4 13 0 10 0 9 2 7 10 0 9 13 16 0 12 9 1 0 9 13 9 1 9 1 12 2
12 7 1 11 13 15 9 15 13 9 0 9 2
27 11 9 7 9 2 11 2 13 1 9 9 1 12 1 10 9 2 3 10 0 0 9 7 9 1 11 2
27 15 13 16 1 9 1 9 13 9 0 1 10 9 1 10 0 9 2 7 9 1 10 9 13 12 9 2
9 9 4 13 9 0 0 7 0 2
15 0 13 15 15 1 15 2 7 1 9 13 15 0 0 2
50 1 10 9 13 15 1 0 9 3 10 9 1 14 13 9 11 11 0 2 1 9 1 16 15 4 13 1 0 9 2 1 10 9 16 0 13 10 9 1 14 4 13 10 0 9 1 10 0 9 2
11 7 15 13 0 14 13 16 9 13 0 2
25 7 0 13 15 1 10 9 3 16 0 9 13 0 0 2 7 4 13 0 9 2 1 0 9 2
18 1 9 13 15 0 0 0 16 11 4 13 10 0 9 1 0 9 2
17 3 13 0 1 10 0 9 1 11 1 10 0 9 1 10 9 2
33 16 0 9 13 1 10 0 9 2 13 15 3 0 3 3 16 15 13 7 13 1 1 9 16 15 3 4 13 10 0 9 3 2
20 6 2 15 4 0 1 7 1 13 1 9 1 16 0 9 4 13 3 0 2
8 9 4 13 9 1 11 0 2
5 15 13 0 0 2
24 3 4 9 1 9 1 9 13 16 10 9 0 9 4 13 10 0 9 1 14 13 1 9 2
28 7 1 11 1 11 7 11 13 15 3 0 0 16 9 4 13 15 1 9 1 10 0 9 7 10 0 9 2
14 3 13 15 0 0 9 15 3 3 13 9 1 9 2
27 1 10 3 0 9 15 15 1 15 13 1 11 2 4 15 13 0 0 9 1 16 15 13 1 10 9 2
21 9 1 16 9 3 13 14 13 0 0 9 13 16 15 3 13 0 3 1 15 2
2 6 2
25 9 4 3 13 0 16 15 13 1 9 2 7 3 0 4 15 1 9 13 9 9 1 10 9 2
18 7 15 13 3 3 1 10 0 9 9 2 7 15 13 10 0 9 2
21 3 13 15 1 15 9 1 3 0 9 15 4 13 16 15 13 9 1 1 9 2
17 15 4 13 16 10 0 9 1 9 4 13 0 1 0 0 9 2
24 11 9 1 9 13 16 12 9 1 10 0 9 1 10 9 13 0 1 10 12 0 0 9 2
21 9 13 10 10 9 2 7 15 13 0 0 9 15 15 3 4 13 0 14 13 2
14 16 9 1 9 13 2 4 15 4 13 10 0 9 2
7 15 13 3 3 3 0 2
13 0 9 13 0 0 9 2 1 0 9 1 9 2
21 16 9 9 13 1 9 1 0 9 2 13 15 0 9 1 14 13 15 1 0 2
62 0 13 15 3 16 16 11 0 13 9 3 1 14 13 9 7 9 2 4 15 1 9 2 16 0 9 7 9 7 0 9 3 4 13 1 1 0 9 1 0 9 2 13 10 0 9 1 9 1 0 9 2 1 14 13 14 13 9 1 9 0 2
49 1 16 9 4 13 9 1 0 0 9 2 4 15 13 1 1 16 15 4 13 10 0 0 0 9 7 9 2 15 13 16 15 2 7 3 0 9 2 0 13 9 1 15 15 13 10 0 9 2
14 16 15 13 4 15 13 0 7 0 1 9 1 9 2
30 9 7 0 9 4 13 9 14 13 2 7 10 0 9 4 3 13 1 1 9 11 2 13 1 10 0 9 1 9 2
22 1 10 0 9 15 9 13 14 13 2 4 10 0 13 15 1 14 13 1 12 9 2
30 10 9 13 3 3 3 0 2 7 4 1 9 1 0 10 0 9 2 1 10 9 13 1 9 1 0 7 0 9 2
8 15 15 4 13 14 13 9 5
3 11 9 2
2 9 2
3 0 9 2
3 9 9 2
3 0 9 2
3 9 13 2
3 0 9 2
11 11 4 13 10 0 0 9 2 11 11 2
11 10 0 7 0 9 11 4 13 10 9 2
15 3 13 15 1 9 2 7 1 10 9 13 9 1 11 2
13 13 10 9 1 10 0 2 0 9 1 0 9 2
15 15 4 13 1 12 7 13 12 9 1 10 0 9 9 2
21 10 0 9 1 9 2 15 13 1 0 9 2 13 11 11 2 13 11 1 9 2
12 1 9 0 0 1 9 13 15 9 1 9 2
9 15 4 13 10 9 1 9 10 2
7 7 3 13 15 3 9 2
28 12 9 0 2 16 9 11 13 1 0 9 1 11 7 0 11 13 1 1 9 2 13 9 7 13 1 9 2
12 2 8 2 8 8 8 8 8 8 8 2 2
10 2 6 2 15 13 3 0 11 2 2
19 11 13 0 1 12 9 7 9 1 9 2 15 13 1 11 11 1 12 2
25 15 13 3 3 1 10 0 9 2 7 3 1 12 9 13 15 1 1 11 2 10 9 1 11 2
17 11 13 9 1 0 9 2 13 15 3 7 13 1 10 0 9 2
5 15 13 12 9 2
13 11 13 0 9 1 9 1 10 10 9 1 11 2
26 10 0 9 2 13 12 2 16 15 13 9 0 9 1 11 11 2 13 15 1 10 0 9 1 9 2
6 9 9 13 3 0 2
9 10 0 9 13 1 9 11 9 2
9 1 9 13 15 0 1 0 9 2
3 2 11 2
5 13 1 9 2 2
14 7 15 13 0 1 11 2 10 9 7 10 12 9 2
28 1 9 13 15 3 10 1 14 13 15 1 16 11 11 2 12 2 13 0 12 9 1 14 13 9 1 9 2
21 3 0 13 15 16 15 3 13 10 0 9 1 10 12 9 9 1 12 9 0 2
25 11 13 10 0 9 7 0 9 15 0 13 2 13 2 13 7 13 9 0 1 14 13 15 0 2
14 1 10 9 13 9 15 0 1 10 0 9 1 9 2
27 15 13 3 10 9 16 9 9 4 13 1 11 11 2 7 15 13 1 14 13 1 10 9 15 13 1 2
16 1 11 9 13 11 10 0 7 13 10 0 9 1 12 9 2
31 7 3 10 0 9 0 9 13 1 9 7 9 1 10 9 2 13 15 9 1 11 15 13 1 9 9 9 1 10 0 2
7 9 13 11 1 0 9 2
40 3 1 9 2 9 11 2 13 15 1 12 9 1 1 12 9 1 9 1 0 2 9 15 4 13 15 1 14 13 9 1 15 15 4 13 1 10 0 9 2
15 11 13 3 0 1 16 11 13 10 0 1 10 0 9 2
23 7 10 9 1 9 13 1 0 4 13 10 0 9 1 9 1 9 1 10 0 10 9 2
24 7 15 4 13 1 14 13 10 0 0 9 15 13 9 10 0 9 7 10 0 9 1 9 2
12 9 13 1 12 9 2 1 11 9 1 9 2
46 15 13 10 0 9 15 13 15 1 10 0 2 7 0 9 1 9 2 9 1 9 2 9 2 9 2 9 2 9 7 0 9 2 13 1 9 1 9 15 13 1 1 10 0 9 2
45 1 10 9 13 9 0 1 10 0 9 9 1 9 2 0 15 15 13 10 9 1 10 0 9 1 11 0 2 0 7 0 0 9 2 15 13 1 9 7 13 14 13 1 9 2
20 11 0 9 13 10 9 1 1 9 2 1 10 0 0 2 7 0 0 9 2
30 0 15 15 1 10 0 9 13 9 7 9 1 10 0 9 2 13 15 1 10 0 9 3 0 1 10 9 1 11 2
27 15 13 10 0 9 14 13 1 1 10 0 0 9 2 15 13 10 0 9 9 1 10 1 9 0 9 2
26 11 13 1 0 0 2 13 15 10 9 7 10 9 2 13 1 1 9 10 0 9 1 9 0 9 2
14 7 10 0 9 13 11 2 10 9 7 10 12 9 2
45 0 1 9 7 0 1 10 0 2 0 1 10 0 9 7 11 0 9 2 1 10 0 0 9 7 0 0 9 2 13 9 9 1 10 0 9 1 15 15 4 13 14 13 9 2
34 15 4 13 1 16 11 11 2 10 12 15 1 10 9 4 13 1 14 13 0 0 9 1 10 9 1 11 2 13 0 1 10 9 2
23 11 13 10 0 9 1 15 9 13 1 1 2 7 13 10 0 9 1 9 1 0 9 2
17 9 9 13 16 15 3 0 13 10 0 9 9 13 1 0 9 2
19 1 0 9 13 11 10 9 15 13 1 1 9 1 0 9 1 11 11 2
12 9 13 10 0 9 1 9 1 9 0 9 2
18 15 13 10 9 1 9 16 10 9 13 7 13 10 9 1 1 9 2
18 1 11 4 15 13 10 9 1 9 0 9 7 0 9 1 1 11 2
12 7 1 9 13 3 10 0 9 1 9 9 2
16 1 7 0 13 10 0 0 2 0 0 9 1 9 0 9 2
14 1 3 9 4 9 13 9 1 9 11 11 11 9 2
23 15 15 13 9 2 1 10 0 9 7 10 0 0 9 2 13 16 9 10 13 10 9 2
28 15 13 10 0 9 9 2 9 15 13 1 1 10 0 9 2 9 15 9 13 7 13 1 9 1 10 9 2
27 14 13 1 10 0 9 14 13 10 9 0 9 2 9 7 0 9 9 2 13 0 7 0 1 14 13 2
17 7 0 13 15 1 16 0 2 0 9 13 1 9 7 9 3 2
2 9 2
2 0 2
2 0 2
2 0 2
12 11 10 4 3 4 13 15 1 10 9 9 2
8 15 13 10 0 9 1 9 2
37 7 15 13 0 16 15 1 9 13 1 9 7 10 9 15 15 13 13 9 1 2 7 3 0 2 13 14 13 9 1 9 9 7 9 0 9 2
24 9 13 3 10 0 9 1 11 9 2 11 11 11 2 11 8 8 11 8 11 2 12 2 2
29 3 13 9 9 10 0 9 1 9 9 2 15 0 13 10 0 9 2 7 9 9 2 15 13 9 7 9 9 2
17 15 13 9 1 7 9 7 9 1 10 3 0 1 0 0 9 2
7 11 0 9 13 0 9 2
26 1 0 9 13 15 0 9 1 9 7 9 2 1 0 9 7 0 9 2 1 9 9 7 10 9 2
19 11 8 8 11 8 11 11 11 2 12 2 13 10 0 9 1 0 9 2
29 1 11 11 11 11 8 11 11 11 11 11 11 2 12 2 4 15 13 10 9 0 9 1 9 2 9 7 9 2
22 7 1 10 0 9 13 3 0 9 1 10 0 9 11 11 11 10 9 2 12 2 2
20 11 13 10 9 9 15 0 13 2 7 15 4 3 13 15 1 14 13 15 2
18 0 0 13 15 3 2 3 16 10 9 2 0 1 9 2 13 0 2
16 10 12 9 15 13 1 9 10 2 13 9 7 10 0 9 2
9 3 0 13 11 10 2 9 2 2
19 15 13 10 9 15 13 0 1 14 13 15 1 1 9 1 10 12 9 2
14 15 13 10 1 10 0 9 15 4 13 1 0 9 2
6 0 1 11 11 11 5
5 14 13 10 9 5
2 9 2
2 9 2
2 9 2
2 9 2
4 9 1 9 2
3 0 9 2
2 0 2
18 15 13 10 9 1 9 1 11 12 1 9 1 11 9 0 9 12 2
21 15 13 10 9 1 9 1 12 1 9 1 11 9 0 9 12 2 13 11 11 2
9 3 1 11 11 11 9 1 9 2
6 9 2 11 11 11 5
4 9 13 9 2
15 11 4 10 0 12 9 13 15 10 0 9 1 11 12 2
26 9 13 0 3 9 13 15 1 9 2 7 13 1 10 0 9 14 13 9 1 9 11 7 9 11 2
17 9 13 1 14 13 12 1 9 2 11 11 7 11 11 1 12 2
13 9 7 9 12 2 12 13 3 0 1 0 9 2
17 14 13 1 9 13 3 0 1 10 9 1 9 1 10 0 9 2
16 7 9 4 1 9 13 3 16 15 4 13 3 9 13 9 2
19 16 15 13 2 4 9 13 1 10 0 9 1 0 2 0 7 0 9 2
20 1 10 15 15 13 2 13 15 15 15 13 16 9 3 4 13 1 0 9 2
31 15 13 9 11 11 11 2 12 2 12 2 15 4 13 9 0 9 1 14 13 9 9 2 13 10 9 7 13 1 9 2
21 1 16 9 1 9 13 0 1 9 2 13 15 10 10 9 1 10 0 1 9 2
25 10 9 9 1 11 11 1 9 13 3 3 10 0 9 2 15 0 9 2 11 7 9 12 2 2
27 9 1 9 13 10 0 9 2 7 0 9 4 1 9 13 9 1 1 14 13 16 10 0 9 4 13 2
23 15 13 0 1 9 1 11 16 15 0 11 1 9 1 9 9 11 11 4 13 1 12 2
41 1 9 12 13 3 9 9 2 11 1 9 1 9 1 11 2 2 11 12 2 15 13 9 7 10 0 1 9 1 9 1 9 7 1 1 12 0 9 1 9 2
23 9 4 13 1 1 10 0 9 1 0 9 2 7 3 13 1 1 10 0 9 1 9 2
20 0 13 1 15 1 10 9 1 10 9 15 4 13 1 15 15 13 1 9 2
18 9 13 3 1 0 8 15 13 2 9 2 7 13 1 9 2 8 2
13 15 15 13 10 10 2 13 10 10 9 1 9 2
11 1 10 0 9 3 13 15 15 1 11 2
21 7 15 13 3 3 1 0 0 9 2 15 13 3 0 7 0 0 2 0 9 2
29 14 13 9 9 1 10 9 2 3 15 13 1 12 7 4 13 1 9 1 1 12 2 4 13 1 9 7 9 2
21 9 13 16 9 4 13 9 1 12 9 2 10 0 2 10 0 2 13 1 9 2
6 10 0 9 13 0 2
24 10 0 9 1 9 13 15 1 11 11 11 7 11 11 9 11 0 9 11 12 2 12 2 5
31 4 15 13 9 1 9 4 15 13 1 9 7 9 11 11 11 15 4 13 0 7 13 0 1 10 0 2 7 0 9 2
32 7 2 11 11 13 1 11 11 8 11 2 12 2 3 10 9 2 9 2 4 13 1 9 1 16 10 0 4 13 1 9 2
18 11 13 9 1 10 0 9 1 9 16 15 13 9 3 7 3 9 2
35 1 11 9 2 11 8 11 11 2 12 2 7 11 8 11 2 12 2 2 13 15 3 9 1 9 7 9 4 13 1 9 1 0 9 2
20 2 11 1 9 2 13 10 9 1 11 11 7 11 11 13 1 11 0 9 2
18 15 13 3 10 0 9 1 0 9 4 13 9 9 1 9 1 11 2
8 3 0 4 15 13 1 9 2
28 9 13 3 9 7 9 2 13 1 9 2 4 13 9 1 1 10 0 9 2 1 9 1 9 7 11 9 2
16 15 13 15 11 4 13 1 1 1 14 13 1 2 9 2 2
14 7 11 11 13 0 9 12 1 10 9 0 4 13 2
27 9 2 9 11 11 2 13 0 9 12 10 9 2 2 11 2 11 0 9 2 2 16 15 13 0 9 2
48 2 15 13 3 1 10 0 1 0 9 15 13 1 9 1 9 2 7 3 0 9 1 11 1 12 2 15 13 9 1 14 13 9 1 9 1 11 1 15 15 3 13 7 13 9 1 0 2
33 2 2 2 1 12 4 0 1 9 1 15 15 4 0 13 1 10 9 2 13 9 1 14 13 1 10 9 15 13 1 9 2 2
19 9 13 10 9 15 9 7 9 1 11 4 4 13 1 10 0 12 9 2
16 9 1 11 11 2 11 11 2 4 0 4 13 1 10 9 2
7 9 13 14 13 1 0 2
10 15 13 10 9 3 1 11 7 11 2
17 9 11 2 11 11 7 10 13 0 9 1 10 0 7 0 9 2
18 9 13 9 1 10 9 2 7 3 0 9 1 9 9 4 13 9 2
17 9 1 9 11 2 11 11 11 2 13 1 11 0 9 10 9 2
7 2 0 9 4 3 13 2
6 3 13 15 15 3 5
5 9 1 14 13 5
5 0 14 13 1 5
4 9 1 9 5
3 9 0 5
4 9 7 9 5
3 13 9 5
2 13 5
4 13 1 9 5
19 15 13 9 7 9 2 13 1 9 1 9 1 9 2 13 9 1 9 2
7 3 4 15 3 13 15 2
31 13 15 15 15 13 9 3 1 14 13 16 15 13 10 0 0 1 7 9 7 9 9 1 9 1 9 2 13 11 11 2
7 9 2 11 11 5 11 5
4 9 7 9 2
25 9 1 9 7 9 1 10 1 9 0 2 0 7 0 0 9 4 1 3 0 13 0 1 9 2
13 4 9 13 10 9 2 4 15 4 13 1 9 2
13 15 4 3 2 1 0 9 1 9 2 13 15 2
24 15 4 3 13 1 16 10 9 0 13 14 13 9 1 2 9 2 2 3 16 15 13 0 2
17 9 7 9 1 15 15 13 15 0 4 3 13 3 0 1 9 2
40 10 12 9 15 4 13 14 13 9 1 9 13 11 11 11 2 15 3 13 15 1 1 9 2 0 15 11 3 4 13 1 2 9 0 9 14 13 1 2 2
5 11 13 1 9 2
6 13 15 15 13 9 5
15 9 7 9 9 1 14 13 10 0 1 9 9 13 0 2
43 3 3 3 0 2 16 3 0 9 1 16 9 1 14 13 15 0 3 13 10 0 3 1 9 2 4 13 1 16 15 13 10 0 9 1 9 2 9 2 9 7 9 2
33 13 15 0 1 9 2 13 9 1 2 16 9 4 4 13 9 2 1 0 9 1 10 0 9 1 9 2 9 2 9 7 9 2
10 13 15 3 13 3 0 9 1 9 2
18 10 3 0 1 15 13 0 2 0 7 0 1 10 10 3 1 9 2
16 15 13 3 16 15 3 13 0 2 0 7 0 9 1 11 2
33 7 15 15 13 0 2 15 15 13 0 7 15 3 0 13 1 9 1 14 13 1 9 2 13 10 9 15 13 7 3 3 15 2
10 15 13 3 3 15 9 3 13 1 2
17 15 13 1 10 15 10 15 3 13 1 9 1 14 13 9 10 2
29 15 13 10 9 15 13 9 1 9 1 12 7 15 1 9 7 9 4 13 10 9 13 1 16 15 13 1 15 2
29 15 13 15 15 1 12 2 12 9 4 13 1 15 1 9 0 0 9 2 7 3 13 1 1 10 9 1 9 2
16 15 13 15 15 4 13 10 9 1 10 9 7 13 0 0 2
12 15 15 13 0 7 3 3 4 13 0 0 2
15 15 15 13 16 9 4 13 0 14 13 1 1 3 9 2
17 15 1 15 15 3 4 4 13 1 9 7 4 13 1 1 9 2
34 15 13 3 1 10 9 15 1 12 9 3 13 0 1 9 2 13 9 7 15 1 12 9 3 4 4 13 16 9 3 13 3 0 2
25 1 10 9 13 10 9 1 0 9 0 16 15 13 0 1 9 2 1 16 15 13 12 9 0 2
32 10 9 1 9 3 15 3 13 1 9 2 13 3 10 0 0 2 1 1 9 9 1 9 7 9 2 9 2 9 7 9 2
20 15 4 13 1 14 13 1 0 0 9 1 10 0 9 2 0 1 10 9 2
25 9 13 1 9 7 9 2 7 15 4 10 13 0 1 16 15 13 0 1 10 9 1 3 15 2
8 15 3 1 9 1 10 9 2
20 10 9 15 13 11 1 14 13 9 7 13 16 15 13 9 0 9 7 9 2
18 16 12 1 12 9 1 12 7 12 13 1 10 7 10 9 1 9 2
15 15 13 10 9 16 12 9 1 15 4 13 1 10 9 2
27 13 15 15 15 13 9 3 1 14 13 16 15 13 10 0 0 1 7 9 7 9 9 1 9 1 9 2
11 4 15 13 16 9 13 0 2 7 0 2
18 4 15 13 0 16 9 7 9 10 13 1 9 1 14 13 0 9 2
27 3 3 10 0 9 4 4 13 15 16 15 13 10 0 9 1 16 10 0 9 13 0 1 10 0 9 2
31 10 0 9 1 9 2 11 11 11 2 4 12 9 13 16 12 9 1 15 13 9 0 2 16 9 1 11 13 10 0 2
24 13 15 16 15 4 13 11 0 1 14 13 1 16 15 13 0 0 2 7 13 15 0 0 2
22 1 12 13 15 3 12 9 1 12 9 1 11 2 3 13 15 15 12 9 1 12 2
18 1 9 13 15 1 9 1 14 13 12 2 12 0 9 1 1 9 2
6 4 15 13 15 0 2
2 3 2
7 4 15 13 9 9 0 2
2 3 2
21 6 2 9 4 13 0 2 0 0 1 2 7 15 4 13 9 2 9 7 9 2
18 15 13 15 15 9 4 13 1 2 7 15 13 0 0 1 9 10 2
12 3 3 0 15 10 9 13 1 14 13 9 2
8 15 4 3 13 10 0 9 2
10 15 13 9 7 9 1 10 0 9 2
33 15 13 1 9 12 9 1 9 2 9 1 15 13 1 9 2 7 15 13 1 12 9 1 0 9 15 13 10 9 9 1 9 2
9 15 13 0 9 7 9 1 9 2
18 15 13 9 1 0 9 1 9 7 0 9 15 9 3 3 4 13 2
16 15 13 9 7 9 1 9 13 1 11 7 13 1 11 11 2
24 15 13 9 2 13 9 2 13 1 9 2 9 2 9 7 9 2 7 3 13 15 3 0 2
32 15 13 0 9 2 0 9 2 9 7 9 2 15 9 1 10 0 9 15 4 13 15 0 2 7 15 0 13 1 10 9 2
15 15 13 3 10 0 9 15 13 1 9 1 9 1 9 2
14 15 13 9 1 9 2 1 14 13 1 9 7 9 2
29 1 10 9 13 15 15 0 9 16 15 3 0 13 1 1 14 13 10 9 1 9 1 14 13 1 10 0 9 2
5 4 15 3 13 2
33 2 13 15 1 1 9 2 13 1 9 7 9 10 2 13 10 9 9 2 13 0 9 2 13 10 9 7 13 1 9 13 2 2
19 3 13 10 0 3 1 10 9 1 9 10 1 9 2 9 1 9 1 2
13 9 13 1 9 2 9 7 9 1 10 0 9 2
9 10 0 9 13 1 9 1 9 2
15 0 13 15 0 2 3 16 15 4 13 2 8 8 2 2
14 15 13 10 9 1 0 9 2 15 9 13 10 9 2
21 3 13 15 7 13 1 15 16 15 13 1 3 0 15 13 7 3 0 15 13 2
39 7 3 13 15 1 14 13 0 2 16 15 3 0 13 14 13 9 1 3 15 2 1 15 2 13 10 0 9 1 11 1 16 15 13 1 9 1 9 2
17 9 13 1 10 0 0 9 1 15 10 2 3 1 15 12 9 2
15 15 13 1 9 1 9 9 7 9 9 1 9 7 9 2
43 10 9 13 0 2 16 10 0 3 13 7 13 14 13 9 2 13 0 9 2 13 9 7 13 9 1 0 14 13 1 9 7 9 1 9 1 1 9 2 9 7 9 2
41 15 4 0 13 1 9 1 10 9 2 7 15 4 10 9 13 0 1 14 13 0 9 1 9 2 3 3 10 0 9 1 9 2 9 2 9 2 9 7 9 2
4 10 0 9 5
2 9 2
6 3 1 14 13 1 2
3 10 9 2
4 10 0 9 2
3 10 9 2
2 9 2
3 13 1 2
3 0 9 2
2 9 2
4 9 1 9 2
17 11 9 1 10 9 1 9 13 3 0 9 2 15 13 0 9 2
16 11 9 13 9 0 9 9 1 10 0 9 15 11 4 13 2
5 9 13 3 0 2
18 15 13 3 1 1 9 0 9 2 3 9 9 1 9 7 0 9 2
8 1 0 9 13 9 1 0 2
10 0 7 0 0 1 2 0 2 0 2
6 7 1 10 0 9 2
2 11 2
3 7 9 2
3 6 11 2
10 15 13 16 15 13 1 9 1 9 2
15 15 13 3 0 1 11 2 15 13 16 15 3 13 9 2
18 2 15 13 3 10 15 15 13 16 15 13 0 12 9 1 9 2 2
40 9 13 7 13 16 11 4 13 10 0 9 1 1 9 2 7 3 2 13 2 1 14 13 9 1 9 1 1 9 2 7 15 4 3 3 13 1 10 9 2
20 15 13 3 10 16 11 13 10 9 2 7 15 13 3 3 10 0 1 15 2
31 9 13 16 11 4 13 1 9 1 9 2 7 11 13 16 15 3 4 13 10 0 9 7 3 13 15 0 0 1 9 2
12 3 13 15 16 15 13 9 0 1 1 9 2
22 15 16 11 13 0 9 1 1 9 13 3 10 9 1 10 9 16 15 3 13 1 2
19 16 11 13 0 1 2 4 15 13 15 1 11 1 0 9 7 9 9 2
14 14 0 13 15 1 14 13 1 0 9 13 1 0 2
13 1 9 1 9 4 11 0 13 1 9 7 9 2
7 15 4 9 4 13 1 2
18 16 9 1 9 13 0 1 9 7 9 2 4 3 3 11 13 1 2
23 15 4 3 13 10 9 1 15 15 13 16 15 13 14 13 11 2 1 14 13 15 3 2
14 10 0 2 0 2 9 13 3 3 0 0 1 15 2
24 9 4 13 16 11 4 13 9 1 1 10 0 9 2 7 15 4 3 13 11 1 0 9 2
17 4 15 4 13 10 9 2 4 15 13 1 9 15 4 13 15 2
12 7 13 15 0 10 9 13 1 9 1 9 2
5 15 13 3 0 2
38 3 3 0 16 10 0 9 13 1 16 15 4 13 10 10 9 1 9 2 16 15 13 3 0 9 1 9 2 13 15 3 3 15 1 9 14 13 2
21 16 11 4 4 13 10 9 1 1 9 1 9 9 2 13 3 1 10 10 9 2
25 15 13 3 10 16 11 13 0 1 7 9 7 9 2 7 9 9 7 9 4 13 0 1 11 2
12 15 13 3 9 4 13 1 10 10 9 3 2
26 15 13 16 15 3 13 10 0 9 1 15 10 9 2 4 15 3 13 10 1 9 10 1 10 9 2
3 3 11 5
2 3 2
29 15 13 7 9 7 9 1 14 13 9 1 11 0 9 2 15 13 0 1 9 10 12 2 7 15 13 0 9 2
32 15 13 1 9 16 9 13 9 0 12 1 9 2 15 13 16 15 13 0 1 3 9 3 1 14 13 9 1 10 9 9 2
15 13 1 9 15 15 4 13 1 9 7 11 9 1 9 2
3 0 13 2
17 16 15 13 10 9 2 13 15 16 11 11 0 13 3 15 13 2
15 7 16 15 13 15 13 10 9 2 13 15 0 14 13 2
3 15 13 2
8 9 7 9 1 10 0 9 2
13 7 15 13 9 14 13 12 0 9 0 1 9 2
12 15 13 9 14 13 1 7 13 1 10 9 2
4 0 13 0 2
8 7 15 13 0 0 1 15 2
2 9 2
2 9 2
4 15 13 0 2
15 15 15 4 13 0 9 1 15 2 13 14 13 0 9 2
3 13 9 2
18 15 4 13 0 9 2 7 15 4 13 15 15 13 1 14 13 9 2
14 14 13 1 1 9 1 9 4 0 13 0 0 0 2
11 15 4 3 13 0 14 13 1 0 9 2
8 15 4 13 16 15 13 9 2
16 7 15 4 13 16 9 3 13 9 7 15 13 3 10 9 2
18 15 4 13 3 9 1 15 10 2 7 15 4 13 0 2 0 9 2
12 1 9 1 11 11 9 2 4 15 13 11 2
9 15 4 13 9 1 9 7 9 2
3 0 9 2
10 9 13 16 15 3 13 15 15 13 2
12 15 4 3 13 10 9 15 4 13 10 9 2
27 16 9 4 13 1 15 10 9 1 2 7 15 13 9 1 9 7 10 9 2 13 15 15 0 2 0 2
16 7 3 4 15 13 0 1 16 10 9 0 4 13 10 9 2
13 13 15 9 3 2 13 15 1 1 10 0 9 2
13 15 13 0 9 7 9 2 1 14 13 15 3 2
22 3 4 15 13 0 9 7 10 9 9 1 9 2 7 3 4 15 13 15 1 9 2
6 7 9 4 13 0 2
13 3 15 13 0 1 0 9 7 9 1 10 9 2
7 7 15 13 3 3 0 2
17 7 16 15 13 2 13 15 3 3 10 9 9 2 9 7 9 2
5 7 3 13 9 2
7 3 13 15 10 9 9 2
8 15 13 0 3 0 9 0 2
9 16 3 13 1 9 1 10 9 2
12 9 1 11 13 4 13 0 1 10 15 12 2
13 15 4 10 9 9 13 1 0 0 9 7 9 2
19 10 1 9 15 4 13 2 4 13 3 9 16 15 4 13 15 1 0 2
6 9 1 9 13 0 2
2 9 5
22 3 1 14 13 3 1 10 9 2 7 1 9 13 15 0 9 1 14 13 15 1 2
8 15 13 0 9 1 0 9 2
12 7 3 4 15 3 13 3 3 0 15 13 2
33 11 4 0 13 10 9 1 10 9 7 0 9 7 9 7 15 2 7 15 4 3 13 9 7 13 1 3 9 7 10 9 3 2
18 7 1 15 15 4 13 9 2 13 15 0 0 14 13 10 0 9 2
10 7 13 15 1 16 15 13 3 0 2
21 7 6 2 15 13 0 0 9 15 4 13 15 1 2 7 15 4 13 3 0 2
2 6 2
7 15 13 0 1 10 9 2
19 7 1 9 1 9 9 2 4 15 3 13 15 1 3 15 4 13 1 2
15 15 4 0 13 1 11 2 7 4 3 13 1 9 10 2
19 6 2 3 3 15 15 13 7 13 2 13 15 16 15 13 0 1 9 2
17 15 4 13 10 10 9 1 11 2 7 15 13 0 14 13 1 2
9 15 4 3 13 9 1 0 9 2
4 7 15 9 2
16 4 15 13 0 1 3 10 9 2 7 4 15 13 0 0 2
11 0 9 13 3 1 16 15 4 13 9 2
13 9 10 13 10 9 13 10 0 1 1 11 9 2
6 7 15 4 15 13 2
9 13 15 9 2 13 15 3 1 2
21 15 13 10 0 7 0 9 15 4 13 1 10 9 2 7 15 4 3 13 9 2
22 7 6 2 10 9 1 15 13 0 3 0 2 7 15 13 3 9 1 10 0 9 2
9 10 0 9 1 15 2 1 9 2
17 2 7 16 15 13 1 9 2 1 9 13 15 10 0 0 9 2
8 1 9 1 10 1 15 2 2
9 13 10 0 9 1 7 1 9 2
2 9 2
4 7 0 9 5
10 15 13 3 10 9 1 9 10 9 2
10 7 15 4 3 3 13 9 9 1 2
16 15 4 13 1 9 2 9 7 9 2 15 1 10 10 9 2
3 2 11 2
11 3 13 15 3 0 1 10 9 1 15 2
19 13 1 3 15 13 9 2 10 9 13 1 10 9 1 10 0 9 2 2
5 6 3 2 3 2
9 9 4 13 1 0 9 1 9 2
24 9 13 10 0 9 2 3 15 3 13 2 7 13 15 10 0 9 2 3 15 3 13 2 2
6 7 1 9 13 9 2
23 0 9 1 0 9 4 13 1 1 0 9 7 13 0 1 1 9 0 2 3 0 9 2
17 2 9 13 15 1 3 2 3 2 15 13 3 3 0 0 2 2
27 3 13 15 1 1 9 2 16 9 4 13 2 13 2 13 7 13 10 15 15 13 1 9 2 9 2 2
34 1 10 12 9 10 13 15 14 13 1 10 9 1 9 2 8 2 8 8 8 2 2 2 7 9 0 13 15 1 15 1 9 3 2
24 2 15 13 3 15 15 13 10 0 1 9 2 15 4 13 1 7 1 15 15 13 15 2 5
37 1 9 4 15 13 1 10 9 1 9 2 7 13 16 9 13 0 16 15 13 2 0 9 3 2 3 3 0 9 7 9 3 3 3 0 9 2
7 15 13 15 7 13 15 2
5 13 10 0 9 2
15 9 7 9 7 9 1 9 10 2 7 1 9 10 11 2
5 11 13 3 2 2
23 2 11 13 3 15 15 3 4 13 1 3 1 9 2 15 13 1 1 10 10 9 2 5
16 1 9 13 15 7 10 0 3 14 13 15 10 9 1 9 2
16 15 13 15 13 0 1 10 0 9 14 4 13 10 0 3 2
17 1 9 13 15 9 1 15 2 3 0 2 3 0 9 7 9 2
62 1 10 0 9 2 0 1 9 7 9 2 9 13 10 10 9 3 2 15 4 3 3 13 9 9 2 2 6 2 3 2 2 2 13 15 9 1 11 7 13 15 1 9 2 16 15 7 10 0 13 0 1 9 7 13 1 15 1 9 1 9 2
34 16 15 4 13 16 15 0 13 10 3 0 9 7 16 9 13 1 11 1 9 16 15 13 1 9 2 6 2 3 13 15 0 9 2
10 13 10 0 9 2 1 7 1 9 2
4 10 0 9 5
8 9 12 13 10 9 1 9 2
26 15 13 15 1 1 9 1 10 0 9 1 11 7 13 2 15 0 2 10 0 9 1 9 1 11 2
25 10 9 0 13 15 10 0 9 1 1 14 13 10 2 3 2 0 0 7 0 0 9 1 11 2
49 1 9 4 15 3 4 13 2 6 2 0 1 15 0 2 1 9 10 7 3 13 15 9 1 14 13 1 10 0 9 1 9 2 15 0 13 15 10 0 7 13 15 1 14 13 1 10 9 2
6 3 3 1 10 9 2
18 15 13 0 15 13 13 0 1 9 2 1 10 15 15 13 9 1 2
16 9 10 1 11 13 3 1 2 9 2 9 9 1 10 9 2
58 15 13 10 0 9 1 15 2 1 10 13 11 1 16 15 13 15 9 7 11 13 1 9 3 15 0 10 3 4 13 10 9 2 15 4 13 9 1 15 10 2 16 15 13 0 9 1 14 13 1 10 9 13 15 10 10 9 2
7 6 2 3 13 15 15 2
29 7 3 13 15 0 3 15 0 4 13 10 9 2 16 16 15 3 13 10 9 4 15 3 13 13 14 13 15 2
13 10 9 4 15 3 3 13 2 15 13 0 0 2
12 7 9 13 1 0 9 2 0 0 3 0 2
10 7 3 13 15 3 15 1 10 9 2
18 0 13 15 0 1 11 7 11 2 15 1 9 13 16 9 13 0 2
18 10 9 4 3 3 13 10 0 9 1 11 11 0 9 1 10 9 2
6 1 9 3 2 0 2
15 7 9 13 2 15 11 13 2 10 9 1 0 7 0 2
16 10 9 13 1 2 1 10 0 9 1 14 13 15 15 13 2
16 7 15 15 13 13 3 0 7 13 9 1 14 13 0 0 2
15 11 13 1 2 9 2 2 10 9 1 15 15 13 1 2
7 3 15 13 15 15 13 2
17 7 3 13 15 3 10 9 2 3 0 9 3 13 10 0 9 2
26 15 4 3 13 10 9 1 10 9 7 15 13 9 15 0 13 9 1 16 15 13 0 9 7 9 2
27 7 1 16 15 4 13 3 0 0 1 15 2 13 15 1 16 10 9 13 0 1 15 15 13 14 13 2
21 3 13 15 2 3 15 4 13 2 1 10 9 1 10 9 15 4 13 1 1 2
23 4 15 13 3 16 12 9 9 13 10 9 15 0 1 15 13 0 1 10 10 9 9 2
7 15 13 15 0 15 13 2
18 1 10 0 13 13 15 0 0 14 13 16 15 13 9 1 15 10 2
20 2 15 13 3 0 1 14 13 1 10 9 2 3 13 15 3 10 9 2 2
14 16 15 13 9 2 13 15 0 13 10 0 0 9 2
26 1 9 13 15 0 2 0 1 15 10 10 0 9 13 2 10 0 9 15 3 13 3 10 12 9 2
14 13 15 0 1 15 10 10 13 2 7 13 15 3 2
22 15 13 14 13 9 10 1 14 13 2 13 2 13 7 13 1 9 15 13 13 0 2
14 7 15 13 3 3 16 10 10 13 14 13 10 10 2
22 1 14 4 13 3 0 1 9 1 9 1 1 2 13 15 3 0 0 1 15 10 2
24 7 1 10 12 9 13 15 1 16 2 3 2 15 15 13 15 1 9 13 15 13 10 9 2
16 0 13 15 0 0 9 1 9 1 10 10 9 9 2 9 2
28 7 0 1 10 0 9 4 13 1 9 16 15 13 0 10 9 1 9 7 16 15 1 9 13 9 1 15 2
18 9 1 9 13 14 13 16 9 1 0 7 0 9 3 13 10 9 2
12 7 15 1 15 13 16 15 3 13 15 3 2
11 15 13 3 3 0 0 1 15 10 3 2
21 0 9 2 3 0 1 15 15 4 13 15 0 1 1 3 2 13 1 0 9 2
5 3 13 9 9 2
22 10 0 9 4 13 15 16 15 13 9 0 9 1 9 7 9 13 0 1 10 9 2
11 15 4 3 13 9 2 7 15 13 0 2
13 1 10 7 10 9 13 15 14 13 9 1 9 2
7 15 13 14 13 1 15 2
6 15 13 14 13 9 2
30 1 10 7 10 9 13 15 14 13 2 15 15 13 13 2 9 2 9 2 2 15 13 0 1 1 2 8 2 2 2
53 15 13 14 13 1 9 15 13 1 2 15 13 1 9 7 13 0 1 1 9 1 9 0 11 16 9 1 9 13 0 1 10 9 9 2 16 9 13 0 2 9 13 1 7 10 9 13 1 9 2 6 2 2
19 7 1 10 7 10 9 13 15 14 13 16 15 13 3 0 1 10 9 2
20 7 3 13 15 3 0 3 0 15 13 14 13 15 0 1 14 13 3 15 2
14 15 13 9 1 9 1 9 1 2 15 13 15 2 2
13 9 13 9 7 13 1 9 1 16 9 13 0 2
6 9 13 10 9 9 2
6 9 13 10 0 9 2
25 1 9 13 15 10 9 1 9 7 10 0 9 1 16 2 9 13 9 2 3 13 15 3 2 2
8 9 13 1 11 11 1 9 2
18 15 13 1 9 2 13 1 9 7 13 15 13 0 16 15 13 9 2
25 10 9 9 13 0 7 15 13 0 7 0 2 13 15 15 1 1 10 9 0 9 2 0 0 2
16 0 9 7 0 9 16 15 13 6 1 9 7 13 1 2 2
9 3 13 13 15 3 0 1 15 2
7 7 15 13 3 10 9 2
48 9 13 16 15 1 9 13 3 0 9 1 10 10 2 0 0 1 15 2 7 15 13 9 1 16 15 3 13 1 9 2 15 4 13 2 2 7 16 15 13 9 15 13 0 0 9 1 2
7 3 16 15 13 0 0 2
5 3 15 13 0 2
10 3 15 13 10 12 15 13 15 1 2
8 0 3 13 15 3 0 9 2
23 15 4 3 13 9 10 2 15 13 3 16 15 13 9 1 0 9 7 15 4 3 13 2
9 3 9 13 0 1 10 10 9 2
14 7 2 3 15 4 13 1 10 0 9 1 0 9 2
6 10 9 13 3 0 2
7 1 9 4 15 13 9 2
2 0 2
6 13 11 10 0 0 2
24 11 11 0 9 4 13 14 13 10 0 9 2 7 1 9 13 11 1 10 3 0 0 9 2
3 0 9 2
66 15 0 13 3 0 0 1 16 9 15 13 9 1 9 9 2 13 0 0 1 9 2 0 7 0 2 2 6 6 2 3 13 15 3 1 0 16 15 13 12 2 7 15 13 15 1 14 0 3 13 15 1 9 15 15 13 1 10 10 9 7 10 0 9 2 2
17 10 9 13 3 3 10 7 0 7 0 9 1 15 14 13 9 2
30 0 0 0 2 15 13 15 16 7 11 11 7 15 10 9 4 4 13 1 9 2 1 1 10 0 0 7 0 9 2
4 3 2 11 2
9 15 1 10 9 4 13 1 9 2
45 3 15 13 13 11 9 10 0 0 7 0 0 15 0 9 13 1 1 16 15 1 3 13 9 2 0 1 2 9 13 3 3 15 15 0 13 1 1 0 9 2 7 2 2 2
30 4 15 0 13 3 3 2 16 0 7 0 9 1 10 10 9 13 15 13 3 0 14 13 9 2 0 1 0 9 2
11 7 1 3 9 2 3 2 3 2 3 2
8 4 15 13 9 1 15 3 2
8 13 11 0 0 0 7 0 2
31 7 4 15 0 7 0 13 3 0 16 9 13 10 0 0 9 2 1 9 1 9 7 0 9 1 14 13 1 0 9 2
42 7 3 2 15 13 3 14 13 15 0 3 3 2 7 4 9 0 13 3 0 16 15 1 9 4 13 9 1 0 9 1 9 1 9 1 9 1 14 13 1 9 2
8 4 15 13 0 1 0 9 2
2 9 2
14 0 15 2 16 15 13 2 15 13 15 0 1 9 2
11 13 16 15 3 4 13 15 1 14 13 2
6 15 13 3 0 0 2
9 7 3 13 15 0 13 0 0 2
6 10 9 1 15 2 2
16 7 3 13 15 3 0 10 15 13 16 9 10 3 4 13 2
2 13 2
32 7 1 15 15 13 0 2 15 13 0 1 16 15 13 10 0 9 2 3 16 15 13 15 9 1 14 13 0 0 1 9 2
6 0 9 7 0 9 5
6 3 13 10 0 9 2
27 1 16 15 13 0 1 0 13 15 3 0 16 15 13 9 0 1 14 13 1 1 10 0 2 9 2 2
44 1 9 13 15 1 9 16 15 13 1 1 10 0 9 16 15 13 1 1 10 9 1 11 2 13 15 0 1 0 9 1 11 16 15 13 10 9 1 11 11 1 9 1 2
19 14 13 15 9 1 13 2 1 15 15 4 13 10 9 2 10 0 9 2
20 7 0 3 2 13 15 15 15 13 3 4 15 3 13 9 1 15 1 15 2
39 15 15 13 15 0 13 16 10 9 13 1 7 13 15 16 15 0 4 13 15 1 9 15 15 15 3 4 13 9 1 10 9 1 11 2 3 4 13 2
30 15 13 0 0 0 1 9 7 9 1 14 13 12 9 1 9 16 15 4 13 15 10 0 7 0 9 1 0 9 2
25 15 13 1 9 10 0 9 16 15 0 4 13 1 10 1 15 15 13 1 10 9 15 4 13 2
8 10 9 1 0 9 13 15 2
16 15 13 1 10 9 10 9 1 11 2 3 1 9 10 9 2
41 7 9 10 13 16 15 13 0 1 9 1 10 0 9 2 3 16 15 3 13 0 14 13 1 16 10 0 9 1 9 3 13 9 1 0 1 10 9 0 9 2
29 7 1 9 1 10 0 9 5 0 9 4 15 1 3 13 3 15 1 3 1 11 1 16 15 13 15 1 15 2
20 3 3 13 15 3 0 1 0 9 14 13 10 0 0 9 1 9 3 1 2
5 7 15 13 15 2
32 16 10 7 10 9 15 4 13 10 9 1 11 13 1 7 13 1 10 0 0 9 15 13 7 13 3 16 9 10 13 0 2
24 1 0 0 9 15 13 9 7 9 1 9 16 15 0 13 12 9 9 1 10 9 1 9 2
22 15 13 0 16 9 1 11 4 4 13 16 15 13 10 9 1 11 1 9 7 9 2
48 7 16 10 0 9 3 4 13 9 1 10 10 11 2 3 4 15 3 13 1 15 15 13 1 9 2 15 15 13 1 9 2 15 15 13 0 9 7 15 15 13 0 9 1 9 1 9 2
13 3 13 15 0 3 3 14 13 9 1 0 9 2
7 11 7 9 2 10 9 2
24 10 9 4 3 13 1 11 2 7 15 13 15 3 1 14 13 0 9 1 9 13 1 15 2
31 9 13 0 1 0 9 2 1 9 3 10 9 4 13 2 0 9 2 1 10 10 2 7 0 13 0 1 9 1 15 2
13 15 13 3 0 1 11 7 11 2 9 13 9 2
16 1 14 13 10 9 13 11 10 10 9 1 11 7 11 12 2
10 15 13 3 3 10 0 15 4 13 2
30 9 1 2 11 8 2 2 2 11 8 2 2 2 8 8 2 7 2 9 2 4 4 0 13 1 9 10 0 9 2
19 15 4 1 7 1 13 1 10 9 15 13 2 9 2 1 10 0 9 2
20 9 1 11 13 3 3 0 2 9 13 2 9 13 0 2 9 13 3 1 2
4 9 13 0 2
13 15 13 3 3 3 0 15 15 13 1 11 11 2
13 1 7 1 11 10 13 16 9 13 0 1 0 2
9 7 2 3 4 15 13 3 0 2
22 11 4 10 0 9 13 1 0 9 2 15 13 9 7 15 13 0 1 14 13 0 2
11 15 13 0 15 13 15 3 1 10 9 2
14 7 9 4 13 1 0 9 1 11 2 11 7 11 2
21 3 13 15 3 9 1 15 10 15 13 10 0 1 2 7 3 15 4 13 3 2
36 3 13 15 14 4 13 1 10 9 1 9 15 13 1 9 3 15 13 1 2 15 15 13 2 0 2 7 3 10 9 13 15 1 10 9 2
5 3 13 9 1 2
21 0 13 4 15 13 16 9 13 1 12 9 2 10 0 2 0 9 7 1 9 2
25 0 9 13 15 15 13 2 11 9 2 3 1 11 2 3 16 15 13 10 9 1 0 9 2 2
28 15 13 1 9 0 2 13 14 13 0 0 7 2 0 2 2 7 15 4 13 0 7 0 14 13 1 9 2
15 9 1 0 9 13 0 9 1 10 12 9 11 7 11 2
16 15 13 1 9 9 15 13 1 9 2 1 9 1 9 3 2
7 13 11 9 1 0 9 2
17 10 9 4 4 13 1 1 9 10 2 7 4 13 0 0 9 2
28 11 13 1 14 13 9 1 10 9 2 7 4 13 14 13 1 9 3 2 7 3 13 10 0 9 15 3 2
12 9 1 9 13 15 15 13 2 0 2 9 2
13 15 4 13 1 1 9 1 9 15 13 1 9 2
19 15 13 15 16 15 13 16 15 4 13 0 0 9 15 4 13 1 9 2
8 10 0 9 1 15 13 11 2
28 15 4 13 0 1 9 3 2 7 1 0 9 13 15 2 0 2 9 2 0 1 9 1 0 7 0 9 2
8 10 9 13 15 0 1 1 2
9 15 13 9 16 15 13 1 9 2
23 9 2 7 3 9 2 13 2 10 0 9 1 0 9 1 10 0 9 2 2 11 2 2
7 9 3 13 2 0 2 2
19 15 4 3 13 1 10 9 1 9 1 10 9 2 15 4 13 15 0 2
13 3 4 15 13 15 1 15 15 13 10 0 9 2
26 4 15 13 1 9 1 10 9 1 11 2 7 13 15 14 13 1 3 11 2 11 7 11 11 13 2
22 4 15 13 1 10 0 9 1 10 9 2 7 13 15 14 13 3 9 7 9 13 2
25 13 15 14 13 1 10 9 1 10 9 2 7 13 15 1 10 9 15 13 3 15 3 3 13 2
12 10 0 9 3 13 2 15 13 3 1 2 2
6 15 13 15 3 1 2
9 6 2 15 15 4 13 9 1 2
16 15 13 9 1 10 9 1 10 9 2 11 9 7 10 9 2
21 9 9 1 10 9 13 1 13 15 3 1 9 10 0 9 13 1 15 1 9 2
20 15 4 13 1 15 2 7 3 0 1 16 9 13 1 10 9 15 13 1 2
9 0 9 13 15 3 10 0 9 2
15 9 4 3 13 1 9 1 15 9 13 15 0 1 15 2
27 15 13 3 1 16 16 15 13 1 1 10 0 9 13 15 1 0 9 2 15 13 9 2 9 7 9 2
13 9 13 1 14 13 10 9 1 9 1 0 9 2
11 15 4 3 13 1 9 15 13 10 9 2
9 0 9 13 0 0 0 1 9 2
8 15 13 3 0 9 1 9 2
20 15 4 13 10 0 9 0 2 3 16 15 4 0 13 1 16 15 13 1 2
9 1 9 4 10 9 4 13 0 2
16 15 15 13 3 7 7 1 10 9 2 13 1 9 1 9 2
15 2 13 10 9 1 10 9 2 7 3 1 9 12 2 2
10 3 13 15 0 16 9 13 10 9 2
21 16 15 15 0 13 10 9 13 9 15 13 2 9 2 2 4 9 13 0 0 2
31 16 15 13 9 7 13 10 9 2 4 15 13 16 15 13 10 9 1 11 2 16 9 15 13 1 0 9 3 13 3 2
10 1 10 0 9 13 3 15 10 9 2
20 3 4 10 9 0 13 2 1 0 9 2 3 16 9 13 14 13 15 0 2
7 3 13 3 10 0 9 2
4 9 13 0 2
16 7 13 15 9 15 4 13 1 10 9 2 7 15 13 9 2
21 3 9 1 11 4 2 13 2 9 1 10 15 0 9 2 7 9 4 13 0 2
7 9 13 10 0 9 3 2
12 15 13 14 13 1 0 2 0 9 1 9 2
19 3 4 15 3 13 14 13 9 1 14 13 1 9 7 13 9 1 15 2
25 7 2 16 9 1 11 4 13 1 1 10 9 1 15 9 13 15 3 3 0 16 9 13 9 2
16 3 4 9 13 1 9 1 14 13 15 1 16 9 13 0 2
14 9 13 0 2 7 15 1 9 13 0 1 14 13 2
11 3 13 15 16 10 9 13 2 0 2 2
27 3 13 15 9 10 2 15 13 16 9 10 13 0 9 2 16 9 13 3 15 13 7 16 9 13 0 2
14 15 13 10 9 1 10 9 2 16 9 3 13 15 2
20 15 4 0 9 13 9 2 9 7 9 2 2 13 15 10 9 7 9 2 2
11 2 13 15 0 14 13 1 10 9 2 2
14 10 0 9 13 15 16 15 4 13 9 1 0 9 2
19 15 4 13 9 10 0 2 7 4 15 13 10 9 4 0 9 13 0 2
40 16 15 13 9 1 9 9 7 9 4 15 0 13 3 16 9 9 13 9 1 10 0 9 15 4 13 1 10 9 2 16 11 11 13 9 1 10 0 9 2
6 3 4 15 0 13 2
12 0 9 7 9 1 14 13 15 13 10 9 2
6 10 10 9 13 9 2
41 16 15 13 9 1 12 9 2 16 9 9 4 13 1 9 10 1 9 2 16 9 9 4 13 10 0 9 2 13 9 0 1 16 3 9 4 13 0 1 9 2
2 9 5
10 9 13 3 0 2 16 15 13 9 2
23 3 4 15 3 13 10 9 1 3 15 4 13 9 1 14 13 15 1 14 13 1 9 2
43 15 13 15 15 4 13 1 9 7 9 2 7 11 2 15 4 13 1 1 0 9 0 2 13 16 15 14 13 9 1 9 13 15 15 3 4 7 13 7 13 1 9 2
29 15 13 9 15 13 15 1 9 2 15 4 13 1 9 1 0 9 7 15 4 1 10 9 13 0 15 9 13 2
28 3 4 15 3 13 16 11 13 14 13 1 10 0 9 2 13 0 7 13 11 10 9 15 4 13 0 1 2
21 3 4 15 15 13 1 9 3 10 9 13 16 9 3 13 15 15 13 0 1 2
23 1 9 4 15 3 3 13 15 16 3 3 11 11 4 13 1 9 2 15 13 15 0 2
26 10 0 9 13 16 0 9 1 11 11 4 4 13 1 0 1 11 11 16 15 4 4 13 1 9 2
2 9 5
11 9 1 9 2 3 9 2 13 3 0 2
15 1 9 1 9 1 9 1 9 13 15 10 9 1 9 2
5 13 9 1 11 2
8 15 13 3 1 0 1 15 2
20 9 1 1 9 9 1 9 9 2 10 9 1 9 7 9 7 9 1 9 2
24 9 4 3 13 1 9 9 2 7 16 15 4 13 15 1 14 13 9 13 3 15 10 9 2
2 3 2
17 9 13 0 2 15 13 0 2 7 15 13 15 3 1 1 9 2
12 3 2 9 9 2 13 2 0 1 9 2 2
7 13 15 1 2 13 0 2
4 13 1 9 2
8 13 1 9 2 13 1 9 2
11 9 13 12 16 15 13 15 1 1 9 2
17 3 13 15 0 14 13 1 9 1 0 2 13 10 9 10 9 2
6 9 4 13 1 9 2
15 1 10 9 9 2 9 7 9 13 3 9 0 0 0 2
10 4 15 13 15 1 7 13 0 3 2
2 6 2
4 13 1 9 2
15 12 9 11 11 0 13 15 15 1 10 0 9 1 9 2
7 9 13 15 12 2 12 2
2 3 2
6 3 4 15 13 0 2
9 13 9 3 2 13 11 7 11 2
8 13 1 16 15 13 3 0 2
9 3 13 15 1 9 15 13 1 2
5 13 10 0 9 2
4 3 0 9 2
5 9 13 0 12 2
2 0 2
4 0 11 3 2
4 3 0 9 2
15 13 1 9 1 9 2 7 13 12 1 14 13 1 9 2
21 0 2 15 13 3 10 9 1 9 2 7 15 13 3 10 0 1 9 1 15 2
20 6 2 13 1 9 2 9 3 1 9 7 9 2 1 12 10 9 2 2 2
8 3 13 15 9 7 13 9 2
11 4 3 13 10 0 1 9 1 9 3 2
17 7 2 9 13 0 12 2 15 13 0 9 16 15 13 9 3 2
7 3 4 15 3 13 0 2
18 6 2 15 13 15 1 1 14 13 10 9 1 3 15 3 13 9 2
4 13 1 9 2
7 7 2 15 13 14 13 2
7 13 15 0 14 13 9 2
13 13 15 15 13 3 0 16 15 13 14 13 15 2
20 15 13 3 3 10 9 1 9 2 3 13 15 1 10 9 7 13 1 9 2
6 15 13 15 13 0 2
34 3 13 15 3 3 14 13 15 10 1 14 13 1 10 9 16 15 10 13 15 15 4 13 2 3 15 4 13 7 3 15 4 13 2
5 15 13 10 9 2
23 7 2 15 13 3 10 9 2 7 15 13 10 9 15 2 0 3 2 13 1 11 2 5
13 0 13 2 15 13 3 9 1 14 13 15 0 2
4 3 13 9 2
64 13 1 15 2 13 15 1 15 13 15 3 3 7 13 15 0 1 12 2 12 9 16 15 13 1 9 2 13 15 15 13 1 11 2 3 11 2 7 13 16 2 3 1 9 13 15 14 13 11 2 2 16 15 13 10 9 11 7 10 10 2 0 9 2
22 9 1 14 13 15 2 13 1 15 15 4 13 2 1 3 14 13 1 9 4 13 2
29 7 16 15 2 13 2 3 0 2 0 9 2 2 13 10 9 15 4 13 1 14 13 2 15 2 3 0 0 2
25 15 4 3 13 14 13 9 9 9 2 7 3 4 15 13 2 3 4 15 13 14 13 15 0 2
21 9 13 16 15 3 13 14 13 15 0 2 16 15 13 0 14 13 1 0 9 2
28 1 1 9 4 15 13 1 10 0 9 2 3 13 15 0 9 1 11 16 15 13 0 14 13 1 0 9 2
44 15 4 3 13 3 16 3 16 15 4 13 1 10 0 9 1 14 13 1 15 13 15 3 0 1 10 9 9 3 1 14 13 15 2 16 15 2 3 2 4 13 15 3 2
32 15 13 3 0 3 15 13 1 2 3 15 4 13 14 13 9 2 3 15 3 4 13 14 13 15 10 16 15 13 10 9 2
17 15 15 0 1 15 13 1 13 16 15 3 13 15 15 13 3 2
31 13 15 3 15 15 4 4 0 13 1 10 0 9 1 10 9 2 7 13 1 1 14 3 4 13 10 9 0 0 9 2
8 7 15 4 15 13 1 15 2
16 2 6 2 2 13 15 3 2 13 3 10 0 9 2 2 2
2 9 2
3 11 11 5
17 1 10 12 9 0 9 4 15 4 13 1 10 9 0 1 9 2
6 12 1 14 13 0 2
41 16 15 13 0 13 0 1 10 9 0 9 0 1 9 10 2 9 1 11 2 7 10 9 9 2 15 15 1 10 9 13 9 1 16 15 13 14 13 1 9 2
7 1 0 9 13 15 9 2
37 15 13 1 1 9 0 9 2 1 9 1 9 1 15 15 3 13 9 1 14 13 1 16 9 3 4 13 9 1 14 13 15 0 1 10 9 2
25 15 13 9 15 4 13 15 1 15 1 9 1 9 2 7 15 13 3 3 3 1 1 10 0 2
12 15 13 3 3 9 15 4 13 1 1 9 2
15 1 9 1 9 13 0 0 0 9 1 1 11 0 9 2
16 9 15 4 13 1 14 13 0 9 1 14 13 14 13 9 2
3 13 9 2
3 13 9 2
13 13 14 13 9 1 9 15 0 13 3 0 1 2
14 13 14 13 1 9 1 10 9 7 13 9 1 9 2
44 1 15 13 15 3 12 9 2 14 13 16 15 13 10 0 7 0 9 2 1 10 0 9 2 12 9 2 10 0 9 7 10 11 0 1 9 15 13 1 14 13 9 10 2
24 15 13 10 9 1 14 13 15 10 2 7 15 1 15 2 1 16 15 0 13 15 1 15 2
32 1 9 1 15 4 15 0 13 0 9 1 0 9 15 1 9 13 10 0 9 1 10 10 0 9 0 2 7 15 13 0 2
3 7 15 2
34 15 13 14 13 1 10 10 9 3 2 16 11 2 9 2 9 2 9 10 7 15 1 10 0 9 10 13 15 1 15 1 0 9 2
14 15 13 14 13 9 1 9 15 0 13 3 0 1 2
18 15 13 14 13 1 0 9 15 15 4 13 1 1 9 15 3 13 2
15 15 13 14 13 1 9 10 7 13 15 1 9 1 9 2
22 10 9 15 0 13 4 13 10 12 9 1 9 10 16 9 10 0 13 15 10 9 2
6 13 15 13 3 3 2
9 15 13 3 1 10 0 1 15 2
24 15 13 10 9 15 0 13 0 1 1 2 15 1 9 13 13 9 1 15 2 9 1 15 2
12 7 1 9 13 0 10 0 9 1 15 10 2
51 10 1 10 0 9 1 9 13 0 1 9 15 4 13 14 13 15 1 1 9 1 14 13 1 15 10 2 15 2 7 10 10 0 2 16 15 3 13 9 1 10 0 9 15 0 4 4 13 1 0 2
20 0 13 1 15 3 2 3 16 15 13 3 0 0 14 13 15 1 11 11 2
43 15 13 3 0 10 9 14 13 9 1 16 15 10 13 1 7 4 13 1 10 0 9 2 0 9 2 0 2 1 10 0 9 15 4 13 14 13 15 1 1 14 13 2
21 15 13 3 1 15 3 0 14 13 0 1 11 11 2 7 3 13 10 9 3 2
33 9 1 10 15 13 14 13 7 13 1 3 0 10 9 13 2 7 15 13 3 1 10 9 3 16 15 13 14 4 13 1 9 2
8 3 16 15 3 4 13 0 2
9 3 16 15 3 13 14 13 9 2
66 7 16 15 13 10 9 2 7 10 10 2 13 1 2 9 13 0 2 0 7 10 1 10 0 9 15 13 1 16 10 9 13 0 9 15 13 10 0 9 1 14 13 15 15 4 13 1 10 0 2 3 15 4 13 15 2 7 15 15 4 13 1 14 13 15 2
2 6 2
19 15 13 3 10 9 7 10 9 15 15 13 2 15 13 15 2 2 1 2
12 3 4 15 3 3 4 13 10 9 1 9 2
16 2 15 4 13 15 1 16 15 13 10 9 1 9 10 3 2
28 15 4 3 3 13 11 1 9 2 7 13 3 1 10 9 1 9 1 10 0 9 15 13 12 9 1 11 2
21 9 15 0 4 13 1 10 9 9 2 7 1 9 13 15 0 0 1 9 2 2
5 15 13 1 9 2
33 15 13 1 9 15 13 9 10 3 16 15 3 13 9 2 7 15 13 1 0 9 15 13 0 9 3 16 15 3 13 11 11 2
24 15 13 3 3 10 0 9 1 0 9 1 9 15 4 13 1 15 2 0 2 1 1 1 2
18 3 13 15 14 13 9 16 15 3 13 3 9 1 9 13 15 1 2
6 11 13 0 0 9 2
3 3 12 5
27 15 13 0 9 16 0 9 15 13 3 9 1 9 10 1 0 9 2 7 15 13 1 3 14 13 1 2
45 10 0 9 13 1 10 9 0 1 15 1 3 2 15 13 3 16 15 13 0 1 9 1 14 3 13 15 15 13 2 7 10 9 15 13 3 7 3 2 16 15 13 10 9 2
8 3 13 15 15 3 0 0 2
2 0 2
7 3 13 10 9 1 15 2
20 15 4 13 10 12 9 1 9 15 13 9 1 1 14 4 13 1 10 9 2
17 1 9 2 3 13 15 3 12 9 2 12 9 16 15 13 15 2
30 0 13 13 15 9 3 15 13 7 13 9 3 16 15 13 15 1 9 2 7 3 1 2 1 14 13 0 0 1 2
11 3 13 15 1 1 10 9 1 12 9 2
27 15 13 15 3 13 14 13 1 10 9 16 15 4 13 15 0 1 9 7 13 16 15 13 10 0 9 2
18 4 15 13 10 9 15 13 1 14 13 15 0 1 9 1 12 9 2
27 15 4 13 15 0 1 9 2 9 7 9 1 12 9 1 2 7 15 13 3 15 15 13 15 1 3 2
5 15 13 0 0 2
47 3 13 15 15 10 2 16 15 13 9 14 13 11 9 1 14 13 9 1 14 13 1 9 2 13 15 3 3 0 14 13 1 1 10 0 1 11 7 13 9 1 1 9 1 9 10 2
22 0 16 15 1 11 4 13 15 3 2 7 15 13 1 9 9 1 14 13 9 10 2
2 9 2
7 15 13 10 9 1 15 2
12 3 13 3 15 7 11 11 7 9 5 11 2
26 15 13 15 1 1 10 9 1 11 2 3 9 2 7 13 0 1 9 1 14 13 10 9 1 15 2
21 11 7 11 13 0 9 2 7 13 1 9 0 1 14 13 1 1 10 0 9 2
7 9 13 1 9 7 9 2
26 15 13 3 3 0 16 15 13 2 7 15 13 0 16 15 13 15 1 14 13 15 1 11 1 9 2
21 15 4 3 13 1 11 1 10 9 3 2 1 14 13 10 1 3 9 1 3 2
41 15 13 9 1 9 3 1 9 7 13 15 15 13 11 7 11 2 7 0 13 15 3 7 13 1 10 0 9 7 13 16 15 4 13 15 1 14 13 1 15 2
5 15 13 15 3 2
8 15 13 0 7 15 13 15 2
6 0 9 7 0 9 2
4 7 0 9 2
7 15 13 15 13 0 3 2
11 1 9 1 11 13 15 3 9 1 9 2
19 15 13 1 0 9 1 9 1 11 1 11 1 14 13 10 1 10 9 2
24 15 13 3 0 3 2 7 15 4 13 1 10 9 15 4 13 14 13 1 15 10 1 9 2
6 10 9 13 1 11 2
15 15 13 15 3 2 7 13 16 15 13 0 2 9 2 2
9 3 13 10 10 9 15 4 13 2
16 4 3 4 13 15 2 7 13 3 15 15 4 13 10 9 2
7 1 15 15 4 13 15 2
8 15 13 14 13 15 1 9 2
7 0 13 15 9 1 15 2
38 1 9 13 15 3 1 11 2 7 3 15 4 13 0 9 1 9 1 12 12 9 2 7 15 13 0 0 1 0 9 7 9 2 0 9 2 2 2
13 3 13 3 10 9 1 10 10 9 15 4 13 2
10 1 9 1 10 9 3 1 10 9 2
25 16 15 0 13 15 15 13 1 9 3 1 9 2 3 4 15 1 9 13 16 9 10 4 13 2
34 7 16 15 3 13 1 9 15 13 9 0 2 7 16 15 3 13 2 7 4 2 13 14 13 9 1 11 1 9 1 12 9 9 2
11 3 13 10 9 1 15 7 3 0 9 2
12 15 13 3 3 15 13 10 10 9 1 15 2
28 3 13 15 16 15 13 10 0 9 1 14 13 1 10 9 1 11 2 7 13 14 13 15 1 10 0 9 2
11 1 10 9 13 15 1 9 1 11 11 2
27 3 4 15 13 1 10 9 1 11 2 16 15 13 1 2 13 1 9 2 7 13 1 10 9 1 11 2
25 3 1 9 13 10 9 2 11 11 2 15 0 1 16 9 1 11 3 4 13 1 9 10 3 2
30 15 13 10 15 0 0 2 7 1 15 15 3 4 13 10 9 1 10 9 2 3 13 15 1 15 15 13 3 0 2
4 13 15 11 2
21 1 3 9 2 13 14 13 9 1 14 13 10 10 0 9 15 13 16 9 13 2
10 13 3 15 1 9 1 10 1 9 2
7 13 15 15 15 4 13 2
8 15 4 13 10 9 1 9 2
55 1 15 15 3 13 11 2 7 3 13 14 13 9 1 14 13 2 3 13 15 15 13 9 3 7 13 1 15 3 0 15 13 1 15 16 15 13 1 9 1 14 13 9 2 7 15 13 1 16 15 13 1 15 3 2
22 0 16 15 15 13 14 13 9 13 1 1 1 15 2 3 16 15 4 13 10 9 2
25 15 10 4 3 13 15 10 9 7 10 9 15 13 0 10 9 7 10 9 2 9 13 0 2 2
5 9 4 13 0 2
14 10 9 2 7 3 0 2 3 13 15 15 1 9 2
23 15 4 13 16 15 3 13 10 0 9 15 15 13 9 1 2 7 10 0 2 0 9 2
20 15 13 15 0 10 9 15 13 1 1 11 1 14 13 11 7 9 1 9 2
23 15 13 0 16 15 3 4 13 3 0 1 2 7 0 16 10 9 13 10 9 1 9 2
7 3 13 15 7 9 10 2
8 15 13 3 3 0 1 15 2
6 13 1 11 2 3 2
11 3 13 10 9 1 15 1 9 11 9 2
18 15 13 3 12 9 1 9 2 13 3 3 2 15 13 0 3 2 2
22 15 13 0 0 9 7 9 16 9 4 13 1 9 7 9 13 14 13 15 1 3 2
15 3 13 15 9 1 11 1 10 1 10 0 9 15 13 2
11 15 13 16 15 13 1 11 1 1 1 2
22 15 7 15 13 14 13 15 1 11 11 1 14 13 0 9 1 14 13 15 10 9 2
18 15 13 1 14 13 9 2 7 3 4 15 13 9 1 9 7 9 2
3 7 9 2
20 0 13 11 1 9 1 14 13 15 14 2 13 2 16 15 13 1 1 9 2
16 15 13 0 9 1 9 10 16 11 4 13 1 10 0 9 2
19 1 15 4 15 13 1 9 2 15 13 0 0 0 9 1 11 7 11 2
5 13 1 0 9 2
22 11 13 3 0 1 1 16 15 13 10 0 15 13 2 7 15 13 3 10 0 0 2
21 15 13 9 1 9 1 0 9 2 7 13 1 11 1 14 13 15 14 13 9 2
11 3 13 10 9 14 13 1 10 10 9 2
19 15 13 9 1 15 3 1 14 13 1 12 0 9 11 4 13 1 11 2
2 0 2
2 0 2
11 15 13 0 14 13 0 9 1 9 10 2
4 6 2 6 2
13 9 13 1 9 12 7 1 12 9 13 15 11 2
17 15 15 13 3 13 15 3 2 7 15 13 3 10 0 9 9 2
13 15 13 1 15 15 4 13 1 10 0 9 1 2
22 15 4 13 1 9 10 2 13 0 9 1 15 7 13 9 1 15 10 1 10 9 2
9 15 13 1 1 10 15 3 0 2
3 13 15 2
6 13 3 1 9 3 2
13 15 13 0 2 7 15 13 3 9 1 10 9 2
14 3 13 15 0 9 1 9 2 15 13 0 3 0 2
20 15 13 0 2 7 15 13 1 9 9 1 15 9 1 12 0 7 12 0 2
8 15 13 10 1 10 12 0 2
7 15 13 10 9 1 9 2
10 15 13 15 3 1 10 9 1 9 2
18 15 4 13 0 2 13 1 9 1 11 7 13 9 1 9 7 9 2
8 15 4 13 10 9 1 9 2
13 15 4 13 1 10 9 15 4 13 1 1 9 2
7 15 4 13 10 2 9 2
4 10 0 9 2
4 3 13 15 2
12 3 13 10 9 1 15 10 1 9 2 3 2
9 15 4 3 13 1 10 9 1 2
5 3 13 15 1 2
3 6 11 2
2 11 5
29 1 10 0 9 1 10 9 15 3 13 3 0 1 1 9 1 11 2 3 13 15 15 3 10 9 0 1 9 2
88 15 13 0 9 9 15 13 1 9 9 2 7 0 1 15 10 2 2 9 2 9 15 13 1 9 7 0 9 1 11 2 0 9 1 9 1 0 11 1 10 9 2 15 13 15 13 9 16 15 4 13 10 7 10 9 2 7 13 9 1 9 2 9 2 9 7 10 9 2 7 13 15 4 13 15 2 3 3 1 0 9 2 7 3 3 1 9 2
26 15 4 4 13 1 0 1 10 9 7 4 0 13 1 1 1 15 15 13 1 10 9 2 9 2 2
12 10 0 0 9 13 10 9 15 13 15 11 2
13 11 13 0 9 7 0 10 9 15 15 0 13 2
27 15 13 0 9 3 1 15 13 9 15 4 13 2 7 9 1 10 9 13 16 15 13 9 1 9 10 2
30 15 4 13 1 14 13 1 10 9 16 11 13 1 9 1 15 2 3 13 15 1 0 1 9 7 13 1 1 11 2
8 15 13 3 15 11 13 1 2
8 15 13 1 9 10 1 9 2
19 9 10 13 9 2 7 15 13 0 1 16 15 15 13 1 11 13 0 2
4 11 13 0 2
15 15 4 0 13 1 16 15 0 13 0 9 1 10 9 2
29 1 14 4 13 15 0 1 10 9 10 1 9 2 3 13 15 10 9 1 9 16 15 13 1 9 14 13 1 2
13 15 13 0 3 2 7 15 1 11 13 14 13 2
23 15 13 9 1 9 1 11 15 4 0 13 1 9 15 13 1 11 0 12 9 1 9 2
34 3 2 16 15 3 13 0 14 13 15 2 7 15 3 13 3 10 0 9 1 0 9 13 1 3 16 15 4 13 15 9 1 9 2
6 15 13 15 0 3 2
13 15 13 0 9 1 9 16 15 13 0 1 9 2
10 10 0 9 13 0 14 13 1 9 2
14 7 15 4 0 13 16 15 3 13 1 15 1 3 2
36 1 10 0 9 4 15 3 13 1 9 1 14 13 1 9 1 11 7 3 4 15 3 13 3 0 1 9 2 7 3 0 1 1 9 2 2
10 10 10 9 13 14 13 15 1 9 2
2 13 2
13 13 10 9 15 13 1 9 2 3 1 11 11 2
9 10 0 9 13 7 9 7 9 2
23 15 13 3 12 9 7 10 0 0 9 2 7 15 13 15 3 10 9 13 1 0 9 2
10 15 13 0 1 10 0 2 0 9 2
4 3 13 15 2
8 10 9 1 0 9 1 9 2
8 15 13 3 15 13 3 0 2
5 16 15 3 13 2
7 15 3 13 3 1 9 2
3 13 0 2
7 13 0 1 10 0 9 2
3 15 13 2
12 7 9 13 16 15 1 10 9 4 13 9 2
5 15 13 3 3 2
5 11 13 3 3 2
16 15 13 3 12 9 15 4 13 1 14 13 9 1 10 9 2
5 15 13 11 1 2
14 15 4 15 3 3 13 3 1 14 13 9 7 9 2
24 3 13 15 14 13 10 9 1 0 9 1 11 2 11 2 11 7 11 11 5 0 11 3 2
21 15 13 10 9 1 11 1 9 7 13 0 1 10 9 1 3 15 4 13 15 2
13 3 4 3 11 13 9 1 9 1 9 1 11 5
17 7 1 0 9 1 9 2 3 4 15 0 13 15 14 13 9 2
18 11 13 1 0 9 9 1 9 7 9 1 16 15 1 9 13 15 2
5 7 15 13 0 2
21 0 13 15 3 1 10 9 2 3 13 15 0 0 0 9 1 9 1 10 9 2
36 3 13 15 10 10 9 7 9 7 9 13 14 13 9 1 10 9 2 0 16 15 13 3 0 9 15 13 2 13 10 9 7 13 0 9 2
10 3 13 15 0 9 1 9 2 9 2
3 3 11 2
10 15 4 13 15 12 9 1 10 9 2
12 15 13 14 13 10 7 10 0 1 15 3 2
10 3 10 9 13 1 9 7 10 10 2
4 9 1 9 2
2 9 2
10 15 13 0 1 0 9 1 10 9 2
2 6 2
2 9 2
6 13 3 1 1 0 2
9 13 1 9 1 14 13 15 0 2
3 9 12 2
11 2 11 2 4 3 13 10 9 1 15 2
10 15 13 15 1 10 9 7 13 9 2
8 15 13 0 1 15 2 11 2
3 9 12 2
5 11 11 11 12 5
4 9 9 9 5
25 6 3 2 15 13 0 15 13 1 0 9 1 0 0 9 7 9 2 7 15 13 1 10 9 2
11 3 4 9 10 13 3 0 9 2 2 2
20 16 9 13 0 3 13 15 3 0 7 13 1 10 0 9 15 15 13 1 2
4 6 2 3 2
20 10 0 9 13 3 0 0 7 0 16 15 13 1 1 16 15 13 1 9 2
11 6 2 6 6 13 7 13 1 9 2 2
13 7 3 13 15 0 10 9 16 15 13 1 3 2
8 6 6 6 13 15 15 3 2
11 15 13 2 13 7 13 1 9 2 2 2
34 1 0 9 1 9 2 13 15 15 1 9 7 13 0 1 1 9 7 13 1 10 0 9 2 16 15 13 9 2 10 0 9 2 2
20 7 16 15 13 9 10 13 0 2 3 4 15 3 13 10 0 9 2 9 2
27 16 15 13 9 13 15 9 1 16 15 3 13 0 1 9 1 10 9 2 15 15 0 13 12 0 2 2
32 3 13 15 0 0 1 10 9 15 13 15 3 2 7 15 13 0 3 1 14 13 15 1 16 15 13 15 13 9 1 9 2
17 15 13 3 15 16 10 9 13 3 3 0 1 9 1 10 9 2
25 15 4 13 16 15 13 7 13 15 1 16 15 13 1 14 13 9 1 9 1 14 13 1 9 2
10 7 9 1 9 13 15 3 14 13 2
35 2 6 6 2 15 4 13 1 1 1 10 9 2 15 4 3 3 13 2 2 13 9 2 7 13 15 1 3 1 9 1 9 1 9 2
10 15 13 0 0 9 1 9 10 9 2
21 0 9 13 15 3 16 9 13 3 1 9 2 7 15 13 1 10 9 15 13 2
6 2 9 2 9 2 2
34 6 2 15 13 3 10 9 1 9 16 15 13 1 1 15 1 14 13 1 16 15 13 1 9 2 15 13 3 10 2 0 2 9 2
13 15 13 3 1 15 15 13 16 15 13 14 13 2
4 2 8 8 2
3 8 8 2
14 8 8 8 8 8 8 8 8 8 2 8 8 8 2
12 8 8 8 2 8 8 8 8 2 2 3 2
2 1 2
8 0 9 1 0 9 7 9 2
44 1 15 13 15 0 1 10 9 15 13 2 13 7 13 2 2 7 10 9 15 0 13 3 2 9 2 9 9 2 9 9 2 9 9 2 9 9 2 9 9 2 9 13 2
9 0 9 1 15 13 0 13 0 2
2 9 2
4 10 0 9 5
9 10 9 3 4 15 3 0 13 2
37 1 10 0 3 13 15 15 1 10 9 2 7 1 14 4 13 9 11 11 11 11 9 1 11 1 10 9 4 15 13 15 1 15 10 12 9 2
8 7 15 13 3 13 15 13 2
31 15 13 3 16 0 9 15 4 13 9 1 14 13 0 0 0 1 10 2 16 15 13 9 9 1 14 13 10 10 9 2
45 15 13 1 9 1 9 1 14 13 10 9 2 7 13 10 0 1 10 0 9 1 11 11 15 13 1 10 9 1 10 0 9 7 2 13 15 2 7 10 9 1 10 0 9 2
7 0 9 14 13 1 1 5
14 7 15 13 3 0 9 9 1 3 15 4 13 1 2
10 10 3 0 13 3 3 3 2 3 2
29 0 1 15 13 0 10 9 1 10 0 9 1 12 15 13 15 2 7 15 13 10 9 1 14 13 3 9 1 2
33 10 13 3 10 9 1 9 15 13 2 10 0 9 7 14 4 4 13 1 1 0 9 10 9 9 16 15 13 1 1 9 9 2
35 0 13 3 9 1 16 15 13 1 1 10 9 2 3 3 0 1 9 2 7 15 4 3 13 10 0 0 0 9 1 3 15 13 1 2
79 1 10 10 9 3 13 15 16 15 0 3 4 13 15 1 1 10 9 7 13 16 15 4 13 16 10 9 3 0 7 0 13 16 15 4 13 1 9 2 1 14 13 16 15 13 1 9 16 9 10 13 9 1 14 4 13 15 0 2 7 1 10 0 7 0 9 1 10 0 9 2 7 1 16 9 13 1 9 2
6 3 2 15 13 0 2
8 10 9 4 0 9 3 13 2
17 15 13 16 12 9 1 15 13 10 10 0 9 1 15 15 13 2
44 15 13 3 9 1 16 9 13 2 7 16 3 0 1 15 13 1 10 9 2 7 4 4 13 1 10 10 9 1 15 15 4 13 1 0 7 1 2 15 13 15 0 1 2
23 11 11 9 13 1 9 1 11 11 9 7 10 0 9 15 13 9 9 1 10 0 9 2
26 15 13 10 9 10 9 15 13 1 2 15 13 3 2 0 2 16 15 3 13 10 9 2 13 9 2
9 7 9 13 16 9 3 13 9 2
5 15 13 3 9 2
19 15 13 16 15 4 13 15 7 13 15 2 13 7 0 9 7 0 9 2
25 7 4 13 9 1 15 2 1 14 0 4 13 16 15 3 13 2 0 2 2 16 15 13 15 2
12 16 10 9 3 13 0 3 3 15 15 13 2
5 15 13 10 9 2
25 7 15 13 10 9 15 4 13 7 10 9 15 4 13 3 1 15 15 1 0 7 3 13 15 2
9 15 4 1 9 3 13 9 9 2
5 15 13 3 0 2
20 7 15 13 16 9 13 1 9 7 9 9 2 7 15 13 16 15 13 1 2
14 15 16 15 13 1 16 10 9 3 13 10 0 9 2
7 4 9 10 13 0 3 2
4 0 2 6 2
10 7 3 7 0 4 15 3 13 9 2
24 3 15 15 13 15 9 2 7 3 0 15 15 13 15 7 13 15 1 15 15 13 1 9 2
18 7 9 4 13 3 12 2 7 15 13 0 0 0 1 10 0 9 2
12 10 9 13 3 7 0 15 15 13 1 9 2
28 15 15 13 1 9 2 15 15 13 16 15 13 15 2 15 15 13 16 15 4 13 15 15 13 15 3 13 2
20 15 15 13 3 7 13 15 0 2 0 1 16 15 13 10 10 9 7 9 2
5 15 13 3 9 2
4 15 13 9 2
3 11 9 5
3 6 11 2
12 15 13 3 14 13 0 1 10 0 9 10 2
12 6 2 6 2 15 13 9 15 4 13 2 2
7 11 4 13 10 0 9 2
45 15 13 3 0 1 15 3 14 13 1 1 15 2 7 15 4 13 0 3 7 3 2 1 11 7 1 11 1 9 1 9 2 1 9 2 9 2 9 2 9 7 9 1 9 2
25 7 15 4 3 13 0 9 3 1 3 2 7 3 4 15 13 0 9 3 1 10 0 9 10 2
10 3 3 13 15 15 13 1 11 11 2
14 15 13 9 1 10 9 2 7 13 0 1 10 9 2
40 15 13 3 0 1 9 2 11 13 16 15 4 13 1 15 12 9 0 1 14 13 1 9 2 7 15 13 10 9 4 13 1 10 9 3 2 7 9 13 2
6 7 15 1 9 10 2
15 15 13 3 10 0 0 9 10 9 11 13 1 1 9 2
10 15 4 13 1 1 9 2 1 9 2
20 15 13 9 13 15 2 15 13 12 2 7 3 13 15 1 1 14 13 15 2
10 15 13 15 3 0 2 0 1 9 2
8 7 15 4 13 15 13 0 2
14 9 13 0 2 1 1 1 16 9 0 4 13 0 2
6 7 15 13 10 9 2
16 13 15 15 4 13 16 9 13 1 3 1 9 2 0 3 2
32 11 4 0 4 13 1 9 7 13 9 2 15 4 4 4 13 7 13 1 10 9 2 7 15 4 4 13 10 3 0 9 2
5 15 4 13 15 2
28 15 13 14 13 15 0 9 2 11 2 7 15 13 3 3 0 14 13 9 1 16 15 13 10 10 9 10 2
22 9 13 3 3 9 2 7 15 13 15 0 1 14 13 1 1 10 9 9 1 9 2
18 10 1 9 15 13 9 2 13 3 0 0 2 1 14 13 15 0 2
14 9 7 9 4 3 13 10 0 9 1 10 9 10 2
14 2 6 2 7 15 4 0 13 10 9 1 10 9 2
11 15 13 15 15 0 13 15 1 10 9 2
25 14 13 0 1 14 13 10 0 9 1 14 13 0 7 0 1 10 9 10 2 13 15 13 0 2
7 0 15 0 13 9 2 2
24 10 9 4 15 3 13 1 10 9 2 3 16 15 13 15 15 4 13 16 9 13 1 9 2
16 9 13 0 1 10 9 2 9 1 9 1 0 2 0 9 2
17 15 4 4 13 1 14 13 1 9 2 7 1 10 0 13 9 2
5 1 0 9 11 5
2 3 2
20 15 4 4 13 16 10 7 10 9 4 13 1 10 9 1 10 9 1 11 2
6 15 13 3 0 0 2
23 11 13 3 10 15 15 13 2 7 0 1 2 7 15 13 15 15 4 13 9 2 11 2
6 0 1 15 2 11 2
10 11 13 15 0 1 14 13 15 3 2
11 2 7 1 15 2 3 13 0 9 3 2
8 13 15 1 7 13 9 2 2
2 9 2
4 7 0 9 5
15 1 9 4 15 13 9 2 13 15 2 7 13 15 0 2
5 15 13 15 0 2
19 15 4 3 13 9 15 15 13 4 0 13 1 10 0 9 7 9 0 2
7 15 13 15 10 9 0 2
21 3 13 15 1 16 15 13 7 13 16 15 1 9 13 0 1 7 9 7 9 2
18 10 9 15 13 15 2 13 16 15 13 1 9 1 10 9 9 3 2
19 3 13 15 14 13 1 10 0 9 0 15 10 0 11 13 3 1 11 2
4 3 0 0 2
23 1 15 4 15 13 10 9 15 4 13 16 15 13 0 1 9 1 14 4 13 7 13 2
18 16 15 13 1 11 2 4 15 13 15 3 16 10 0 9 4 13 2
9 15 4 3 13 0 2 13 15 2
8 7 3 13 15 14 13 0 2
13 15 16 15 4 13 1 15 16 15 13 1 9 2
23 13 16 15 13 9 2 13 1 10 0 9 2 7 2 1 14 13 15 0 1 2 13 2
24 3 2 15 13 0 0 2 7 15 13 3 15 15 4 13 10 0 9 2 7 15 3 13 2
23 15 13 3 10 0 9 2 7 10 9 1 9 13 15 1 15 10 12 9 1 10 0 2
18 15 13 3 9 1 15 15 4 13 1 15 16 15 13 15 0 1 2
21 7 16 15 4 13 1 10 12 0 9 1 10 0 2 13 15 14 13 1 9 2
8 4 15 13 10 9 2 3 2
6 10 0 2 0 9 2
27 10 0 9 4 3 13 10 0 9 2 10 0 9 1 3 0 2 10 9 1 9 7 10 9 1 9 2
7 7 15 13 15 0 1 2
9 7 15 4 13 10 0 0 9 2
41 9 13 3 10 3 0 2 3 16 10 0 9 16 15 13 16 15 13 15 1 10 0 9 1 9 2 0 4 13 3 3 0 16 15 3 0 13 1 9 2 5
25 3 2 3 1 0 9 1 9 2 13 15 13 0 1 0 9 2 3 10 9 1 9 1 11 2
17 15 13 3 10 1 14 13 0 7 0 9 16 15 4 13 15 2
3 0 1 2
32 10 0 9 2 11 1 9 1 0 9 1 9 2 15 15 13 1 15 10 1 9 2 13 3 10 9 15 4 13 1 15 2
9 13 10 0 9 1 7 1 9 2
6 1 14 13 9 1 5
12 11 13 1 10 9 3 15 4 13 1 9 2
8 7 15 13 15 1 14 13 2
8 7 15 13 3 0 10 9 2
2 9 2
5 15 13 3 0 2
3 3 0 2
5 3 0 14 13 2
5 3 0 14 13 2
3 3 0 2
14 3 13 15 3 10 9 15 10 9 13 9 1 9 2
5 1 0 9 3 2
3 15 12 2
3 1 9 2
3 7 9 2
13 0 2 3 13 3 3 11 11 1 9 7 9 2
13 15 13 3 1 10 9 1 14 13 10 0 9 2
6 7 13 10 0 9 2
15 15 13 9 13 3 0 14 13 1 10 9 1 10 9 2
9 16 9 13 3 0 1 10 9 2
14 15 13 3 0 14 13 1 9 2 1 10 10 9 2
25 15 13 3 3 9 3 4 13 3 0 9 1 9 1 10 9 2 15 15 7 9 13 1 9 2
9 7 3 13 15 9 1 10 9 2
3 10 9 2
5 3 13 15 15 2
5 1 14 13 9 2
6 1 14 13 1 15 2
3 13 15 2
2 9 2
4 11 11 11 5
4 11 8 8 2
3 1 9 2
13 11 11 11 2 11 11 2 11 11 2 11 11 2
5 2 3 1 9 2
8 11 11 7 11 11 11 2 2
2 9 2
5 11 11 11 9 2
50 11 11 2 9 2 9 2 2 11 11 11 2 9 2 9 2 2 11 11 2 9 2 9 2 2 11 11 11 2 9 2 9 2 2 11 11 2 9 2 9 2 2 11 11 2 9 2 9 2 2
10 2 3 13 15 1 1 10 0 9 2
11 2 15 13 9 1 10 0 9 7 9 2
17 13 15 1 0 0 9 2 16 15 13 0 14 13 1 1 9 2
38 2 15 13 15 1 9 9 2 11 11 2 2 2 11 11 2 2 2 11 15 1 2 2 11 11 2 7 2 11 11 11 11 2 2 11 11 2 2
16 2 15 13 15 10 1 9 1 1 2 7 15 13 0 9 2
19 2 15 13 10 0 1 10 9 1 15 2 14 13 2 13 2 7 13 2
6 2 14 13 0 9 2
9 15 13 3 3 10 0 15 13 2
9 2 15 13 10 9 1 10 9 2
23 2 15 13 10 0 9 15 13 1 9 1 11 1 14 13 1 9 2 9 7 0 9 2
15 2 3 4 15 13 14 13 1 9 2 10 0 9 11 2
30 2 15 1 9 13 0 9 1 11 1 9 2 7 10 9 13 10 9 7 15 13 15 3 1 15 15 13 9 3 2
5 9 13 1 9 2
8 2 3 4 15 13 1 9 2
23 2 15 13 1 16 15 13 1 1 9 1 0 9 1 9 15 10 13 10 0 9 1 2
7 2 15 13 10 0 9 2
19 2 15 13 10 9 1 2 11 11 11 11 11 11 2 1 11 11 11 2
4 15 13 15 2
7 2 15 13 10 0 9 2
9 2 15 13 9 1 9 1 11 2
15 10 9 1 0 9 7 0 9 13 10 9 1 15 10 2
6 2 15 13 10 9 2
13 2 15 3 1 11 13 10 9 14 13 0 1 2
19 11 11 2 1 11 11 7 11 11 2 13 15 0 15 4 13 15 1 2
11 3 4 1 3 9 10 11 11 4 13 2
13 2 15 13 10 0 0 9 15 4 13 9 1 2
17 2 0 0 2 11 13 9 2 2 10 3 0 9 1 11 11 2
6 15 13 9 1 9 2
4 15 13 3 2
7 2 15 13 1 10 9 2
9 2 15 4 13 0 7 0 1 2
28 3 3 0 9 2 7 1 10 9 3 9 2 2 2 2 2 9 11 13 1 0 9 1 9 2 9 2 2
9 2 13 15 9 14 13 1 9 2
5 2 15 13 0 2
6 13 3 1 11 11 2
8 2 15 1 9 13 0 9 2
4 2 0 11 2
14 9 13 15 1 15 1 14 13 3 0 10 9 13 2
10 3 4 15 3 13 10 12 10 9 2
30 2 16 9 4 4 13 1 9 1 10 2 9 2 7 9 4 13 9 1 9 1 11 15 0 13 15 1 14 13 2
6 2 15 13 10 9 2
7 2 10 9 13 10 9 2
6 15 13 0 1 9 2
6 2 15 13 9 9 2
9 2 2 11 11 2 2 1 9 2
14 15 13 15 1 14 13 10 9 9 15 9 3 13 2
8 2 3 4 15 13 9 9 2
9 2 1 14 13 1 9 1 9 2
10 2 3 4 10 9 1 10 9 13 2
16 2 15 13 3 10 0 9 1 11 16 9 13 10 0 3 2
6 2 13 9 7 9 5
4 2 0 9 5
4 2 0 9 5
5 2 4 13 9 5
9 9 13 0 9 16 11 13 9 2
27 2 15 13 3 0 1 16 9 3 4 13 1 9 2 13 11 11 11 2 9 1 9 1 11 0 9 5
25 15 13 1 16 11 9 13 11 9 1 9 1 9 1 11 9 2 16 9 4 13 1 1 9 2
18 11 9 13 1 9 7 1 9 7 9 1 10 9 1 11 0 9 2
21 1 9 13 9 9 15 13 9 1 0 9 1 9 2 0 9 2 9 7 9 2
28 11 13 16 9 13 10 9 14 13 2 7 13 16 9 1 9 4 13 2 16 9 7 9 4 13 1 9 2
18 2 15 4 3 13 10 9 1 9 1 9 0 1 9 2 13 15 5
18 11 11 11 11 2 9 7 0 1 11 1 11 1 11 2 13 0 2
26 2 15 4 13 0 0 9 2 7 9 4 13 9 15 15 4 13 0 9 14 13 1 2 13 15 2
14 11 11 2 9 1 9 1 11 9 2 13 9 9 2
21 15 13 16 15 4 13 9 1 9 2 16 15 4 13 16 9 4 13 1 11 2
21 9 11 4 1 0 9 13 1 0 9 1 11 2 7 16 9 4 13 9 3 2
25 11 13 1 9 0 1 11 9 2 7 13 1 9 1 9 16 15 7 9 1 9 1 11 13 2
21 2 9 4 13 15 1 9 1 0 9 2 7 13 9 1 9 2 9 7 9 2
26 16 15 4 13 10 9 1 9 1 12 9 2 4 15 3 13 10 9 3 1 1 11 2 13 15 2
24 11 1 9 13 15 13 0 16 9 13 9 13 15 1 9 2 16 9 0 4 13 1 9 2
20 2 15 4 0 13 1 14 13 10 0 9 2 7 10 0 9 2 13 15 2
20 11 11 11 2 9 1 11 9 2 13 15 4 13 9 1 9 1 0 9 2
18 2 16 9 13 15 1 9 15 3 13 9 1 2 13 9 0 9 2
22 15 13 9 1 9 7 9 2 7 15 13 3 15 13 0 14 13 9 2 13 11 2
9 15 13 3 0 1 9 1 11 2
14 2 16 15 13 9 1 9 2 13 0 13 10 9 2
17 15 13 3 10 9 15 13 9 1 14 13 1 9 2 13 9 2
29 11 13 11 13 0 9 1 11 9 2 7 13 3 9 1 1 11 2 16 4 15 13 15 15 13 0 7 0 2
11 2 13 1 14 4 13 1 9 1 11 5
2 9 2
5 2 4 13 9 5
4 4 13 9 5
3 4 13 5
3 13 11 2
4 9 3 9 5
7 2 4 13 0 0 2 5
8 2 3 15 15 4 13 2 5
9 2 15 13 0 0 2 13 9 2
4 3 13 15 2
11 9 13 1 1 11 11 16 15 4 13 2
18 9 13 0 1 9 2 7 15 13 3 16 9 15 13 15 13 9 2
24 13 15 10 0 9 1 0 0 9 1 11 16 12 0 9 13 10 0 9 1 11 0 9 2
32 11 13 9 16 12 0 9 1 11 11 11 2 11 2 1 11 4 13 10 10 9 1 10 9 15 13 15 11 11 1 11 2
13 9 1 11 13 3 1 1 16 15 13 10 9 2
11 9 13 1 9 2 7 12 0 13 15 2
5 10 9 4 13 2
14 2 10 12 13 15 1 10 9 2 10 0 10 9 2
25 15 4 3 13 9 2 7 15 4 13 1 15 7 13 1 9 9 2 13 9 11 11 1 11 2
19 2 15 13 12 0 9 2 7 15 13 3 1 1 16 15 13 10 9 2
12 15 4 3 13 1 10 0 1 2 13 11 2
14 15 13 16 15 3 13 10 9 1 11 11 1 11 2
28 2 15 13 1 0 9 7 15 13 3 0 14 13 15 16 15 13 0 14 13 1 9 1 11 2 13 9 2
13 9 4 4 13 1 0 9 7 1 11 7 9 2
11 9 4 3 13 10 9 1 9 1 11 2
23 11 4 13 1 15 2 7 13 14 13 1 9 1 2 11 11 2 2 15 15 4 13 2
11 15 4 13 15 14 4 0 13 1 13 2
24 1 14 4 13 1 12 9 1 11 2 13 15 0 1 14 13 9 1 9 1 14 13 9 2
4 15 13 11 2
6 15 13 9 1 11 2
9 15 13 0 16 15 13 1 9 2
34 11 13 16 15 4 13 1 11 1 10 9 9 2 7 9 1 12 9 15 13 1 9 1 0 9 2 13 0 3 0 1 10 0 2
17 15 13 0 1 1 11 11 2 1 10 9 15 13 0 1 9 2
19 15 13 1 15 12 9 1 9 7 9 2 7 15 13 3 14 13 15 2
2 9 5
17 7 15 13 3 15 9 13 1 16 15 13 1 9 0 10 9 2
20 15 13 3 10 9 1 0 9 2 7 9 15 13 1 11 13 15 3 1 2
7 3 13 15 15 15 13 2
12 2 15 13 14 4 13 16 15 13 1 3 2
9 1 10 13 12 9 0 1 9 2
7 15 13 15 13 0 9 2
6 0 13 15 1 15 2
8 15 13 0 2 1 1 9 2
15 15 13 9 1 9 2 3 16 15 3 13 9 1 9 2
11 15 13 16 15 13 15 1 9 7 13 2
9 10 12 13 2 13 15 3 2 2
7 15 13 10 12 15 13 2
11 15 13 1 12 2 12 9 2 13 15 2
6 15 13 14 13 0 2
22 9 13 10 9 15 15 13 2 13 1 10 9 7 13 1 1 9 1 10 0 9 2
15 3 13 9 9 2 7 13 0 1 9 1 14 13 9 2
10 15 13 15 4 13 9 15 13 1 2
10 15 13 9 1 2 0 7 0 2 2
20 2 15 13 1 15 9 1 12 9 7 9 2 7 15 13 3 14 13 15 2
8 15 13 0 15 3 13 9 2
7 7 15 4 13 15 0 2
17 7 15 13 0 7 0 16 10 10 4 13 1 11 2 13 15 2
9 2 15 13 10 0 9 1 9 2
14 15 7 10 9 4 3 13 9 7 9 2 13 15 2
12 15 13 0 1 2 1 9 1 10 12 9 2
24 3 13 15 16 10 0 9 2 15 13 1 1 9 1 9 0 10 9 9 2 4 13 9 2
19 2 11 11 2 13 10 0 0 9 2 1 12 9 2 10 3 0 0 2
5 7 2 15 13 2
27 10 9 9 1 16 11 13 9 1 10 9 9 3 7 13 16 15 13 10 9 1 9 2 13 9 0 2
13 9 13 9 1 3 2 7 3 13 15 10 9 2
22 11 13 10 0 9 7 1 11 7 11 2 7 15 13 3 10 9 1 15 1 9 2
17 15 4 13 11 7 13 16 9 4 4 13 2 7 3 13 9 2
22 15 13 1 9 11 11 13 15 1 1 10 0 7 0 9 11 11 11 11 1 11 2
9 15 13 14 13 1 0 1 9 2
10 2 15 13 1 10 9 1 10 9 2
27 15 13 0 0 1 9 1 2 7 13 15 16 15 13 1 0 1 9 10 2 13 9 11 11 1 11 2
6 11 13 3 1 9 2
23 1 9 2 3 13 9 14 13 10 9 3 15 9 4 13 0 2 2 2 13 15 11 2
10 0 1 9 13 9 1 11 10 9 2
15 15 13 3 9 1 11 2 7 13 0 1 9 1 9 2
21 15 13 0 1 9 1 9 2 7 0 9 13 15 10 9 1 10 9 1 11 2
6 3 1 13 11 9 2
11 2 15 13 16 15 3 4 13 1 11 5
25 15 13 1 9 2 7 13 16 15 13 1 1 11 11 9 2 0 9 2 2 13 9 1 11 2
16 9 11 11 1 11 11 11 13 3 1 9 1 15 4 13 2
11 2 9 15 4 13 1 2 13 3 0 2
3 7 0 2
14 15 4 13 1 1 0 9 2 7 3 13 10 0 2
17 10 0 0 14 13 1 2 13 9 1 0 0 9 2 13 11 2
13 15 13 3 1 16 11 11 4 13 15 1 11 2
30 11 13 1 9 3 1 12 16 15 13 1 9 1 9 7 13 1 10 9 1 9 2 15 15 13 15 14 13 0 2
11 3 4 15 13 1 2 0 0 0 2 2
11 11 13 9 4 13 9 1 9 0 9 2
7 2 15 4 4 4 13 2
14 9 4 13 15 0 0 7 13 1 9 2 13 15 2
14 2 15 15 4 13 2 4 13 7 13 15 12 9 2
12 15 13 15 1 10 0 7 0 7 0 9 2
11 15 13 0 9 1 10 9 1 10 9 2
17 15 4 3 13 0 9 1 15 1 9 1 9 2 13 15 1 2
16 11 11 4 3 4 13 1 9 2 1 10 10 9 1 12 2
12 15 13 9 1 10 9 15 13 1 3 1 2
20 11 13 3 15 15 13 2 7 15 4 13 0 7 13 0 0 16 15 13 2
10 3 1 12 4 15 13 1 15 0 2
12 11 4 3 13 1 11 7 13 1 0 9 2
18 11 11 1 11 11 11 13 3 0 1 16 15 13 9 1 0 9 2
4 2 0 0 2
15 16 3 15 4 4 13 2 4 15 3 13 15 1 15 2
16 15 13 3 15 15 13 0 1 14 13 9 10 2 13 15 2
20 16 11 11 11 4 13 0 9 1 9 2 13 15 1 12 9 1 11 11 2
14 2 15 13 9 13 16 15 13 10 9 15 4 13 2
25 15 4 3 4 13 1 10 9 3 2 7 15 13 0 0 15 13 14 13 9 1 15 1 11 2
7 15 13 0 2 13 15 2
8 9 10 4 13 9 1 9 2
9 2 15 4 13 9 1 9 3 2
8 15 13 14 13 9 1 9 2
17 7 3 4 15 3 13 15 1 9 7 13 9 3 2 13 15 2
2 9 2
11 13 7 13 9 1 12 2 7 13 9 5
5 0 1 11 9 5
3 1 9 5
4 12 9 0 5
9 9 1 11 13 9 13 3 0 2
3 0 9 2
11 0 13 11 12 9 15 4 13 1 9 2
14 12 1 15 13 10 12 0 9 13 1 7 1 9 2
21 11 13 11 1 14 13 0 1 9 1 9 1 9 1 11 11 11 10 0 9 2
21 1 9 9 1 11 9 4 10 0 9 1 11 0 9 1 9 1 9 0 13 2
23 0 9 13 10 9 1 9 13 3 0 2 7 1 10 3 0 9 4 4 13 1 9 2
21 15 13 1 16 9 13 1 10 9 16 11 13 1 13 0 1 9 1 9 1 2
7 2 15 13 10 0 9 2
15 10 9 1 9 13 10 1 9 15 4 13 0 9 1 2
36 1 10 10 12 9 1 9 4 9 13 10 2 7 15 4 0 9 13 1 10 0 9 15 13 1 9 2 13 9 1 11 2 11 11 11 2
21 1 9 13 15 3 7 0 11 11 7 11 11 15 13 15 0 1 9 1 9 2
7 15 13 9 13 3 0 2
14 9 11 11 13 16 10 9 13 10 9 9 7 9 2
35 2 15 13 10 9 1 14 13 9 1 10 0 9 2 7 15 4 3 13 1 9 1 16 15 4 13 0 9 1 10 9 2 13 11 2
23 1 9 9 13 11 3 9 1 14 4 13 10 0 0 9 1 10 12 0 9 1 9 2
11 2 15 13 1 16 9 13 0 1 9 2
10 3 13 15 15 4 13 0 7 0 2
23 7 0 4 15 3 3 13 1 10 9 1 9 2 13 11 9 11 11 11 2 1 11 2
12 11 13 3 9 1 1 12 9 9 1 9 2
30 10 0 9 13 15 1 1 12 7 12 9 9 2 16 9 1 9 7 9 1 9 13 1 9 12 1 12 9 9 2
11 0 13 11 12 9 15 4 13 1 9 2
14 12 1 15 4 10 12 0 9 13 1 7 1 9 2
7 13 1 0 9 1 9 5
6 2 9 13 0 9 5
7 2 15 4 13 3 0 5
3 13 9 5
6 2 13 10 0 9 5
9 0 0 9 13 0 9 1 9 2
8 15 13 0 9 0 0 1 2
2 9 2
9 9 11 11 1 9 1 9 11 2
21 9 1 11 11 4 13 9 1 0 9 2 7 3 13 0 9 1 3 0 9 2
9 15 13 16 15 4 13 9 9 2
23 2 10 0 9 13 0 1 16 3 0 0 9 15 13 2 3 0 13 15 10 10 9 2
19 0 9 13 1 9 1 0 9 1 1 1 9 16 15 13 9 7 9 2
20 15 13 0 9 16 15 13 1 1 10 10 3 1 11 2 13 9 11 11 2
13 15 4 1 1 12 9 13 1 9 7 0 9 2
26 7 4 3 0 13 1 9 1 0 9 1 9 2 16 15 13 15 13 9 1 9 1 10 0 9 2
11 2 15 13 10 9 1 14 13 1 11 2
30 1 9 15 13 15 2 1 1 11 7 11 2 13 15 3 16 15 13 0 0 1 15 1 14 13 9 2 1 9 2
29 16 15 3 4 13 1 9 2 3 4 13 1 15 1 10 0 9 2 13 15 10 7 0 9 1 14 13 15 2
14 11 13 9 4 13 0 7 1 9 1 9 7 9 2
6 2 15 13 0 9 2
17 15 4 13 1 10 10 9 2 0 15 15 13 9 1 10 10 2
14 15 13 0 0 2 7 15 13 3 9 10 0 9 2
9 15 13 0 10 0 9 1 9 2
9 15 13 0 9 9 2 13 15 2
10 2 9 13 9 13 0 16 15 13 2
17 2 15 15 3 1 9 13 2 13 16 15 3 13 9 1 9 2
12 15 13 3 3 16 9 3 13 15 15 13 2
9 15 13 9 13 0 16 15 13 2
18 7 3 16 9 3 13 15 2 13 15 3 10 0 9 1 10 9 2
21 9 13 1 10 0 9 11 11 2 11 2 13 16 11 13 0 1 9 1 9 2
23 2 15 13 10 0 9 15 13 0 0 1 14 13 9 1 14 13 9 7 13 1 9 2
27 16 15 3 4 13 10 0 9 1 9 4 13 1 9 10 2 13 0 9 1 11 1 11 2 11 11 2
12 2 13 15 0 9 4 13 10 0 9 10 2
3 2 6 2
12 1 15 15 13 9 13 15 3 3 3 0 2
9 7 1 9 11 13 15 0 0 2
12 9 13 0 0 7 13 0 0 16 15 13 2
17 16 15 13 0 0 4 15 13 10 0 9 1 9 2 13 15 2
24 9 1 11 2 11 11 2 13 9 1 9 13 0 3 1 16 9 1 11 13 0 0 0 2
12 2 1 14 13 13 9 9 1 0 0 9 2
6 9 10 13 0 9 2
18 1 10 9 13 10 9 0 16 15 13 16 15 4 13 0 7 0 2
10 9 4 13 1 14 13 9 1 9 2
23 11 2 15 3 13 9 1 11 11 2 13 15 13 0 14 13 0 0 9 1 10 9 2
43 2 15 13 16 15 1 9 1 10 9 4 13 9 2 7 3 4 15 13 3 0 2 13 11 7 13 1 10 1 16 11 13 10 0 9 2 11 1 11 2 1 9 2
15 11 13 16 11 1 11 4 13 14 13 0 9 7 9 2
16 2 4 15 13 10 9 1 3 0 9 1 11 4 4 13 2
12 2 15 13 0 1 1 16 9 4 13 1 2
30 7 16 15 13 0 1 15 2 3 13 15 10 9 1 16 15 1 11 13 0 9 1 1 0 9 16 15 13 0 2
15 15 13 3 14 13 0 0 1 14 13 16 15 13 3 2
15 3 0 4 15 3 13 7 13 12 12 0 9 1 9 2
24 2 3 16 3 15 13 0 9 1 9 2 13 15 0 2 13 11 11 2 9 1 11 11 2
17 2 15 13 3 0 0 9 1 9 2 7 15 13 0 0 10 2
34 15 13 3 9 1 15 1 9 16 9 4 13 15 2 1 9 1 4 15 13 0 1 11 7 0 9 1 9 3 16 15 4 13 2
27 15 13 3 0 1 0 9 2 7 15 13 15 13 0 16 9 13 10 0 9 16 15 3 13 1 9 2
10 16 3 13 15 9 15 3 13 0 2
11 15 13 16 9 13 10 0 9 1 9 2
25 2 9 1 11 11 13 12 1 12 9 2 7 15 13 15 10 16 3 15 13 0 1 14 13 2
20 1 14 13 10 9 15 13 7 13 15 0 0 1 9 13 15 0 1 9 2
10 9 1 9 13 0 7 0 7 0 2
19 15 13 10 9 9 3 15 13 0 16 15 13 7 13 15 15 4 13 2
9 3 13 15 0 3 0 1 9 2
34 15 4 13 9 1 9 1 7 1 9 1 14 13 15 15 13 1 15 2 7 0 1 0 0 9 13 9 0 1 9 2 13 11 2
16 15 13 15 14 13 9 1 9 7 9 13 0 1 9 9 2
22 2 16 9 13 15 15 13 2 4 9 13 0 0 7 13 10 0 9 2 13 11 2
13 3 12 9 1 9 1 11 11 4 13 1 9 2
10 7 2 13 11 2 15 13 3 15 2
13 2 10 1 10 0 7 0 9 13 15 9 1 2
14 0 10 9 1 10 0 9 1 10 0 9 13 3 2
17 10 9 13 15 3 0 0 1 9 2 1 9 9 1 11 11 2
8 11 13 3 3 3 11 11 2
17 0 9 13 3 1 11 2 11 7 11 2 7 3 13 15 15 2
6 0 7 0 1 9 5
9 11 11 11 13 0 16 9 13 5
2 9 2
11 11 11 11 13 0 1 10 0 9 11 2
10 3 13 2 11 2 7 0 7 0 2
44 3 16 15 13 0 9 0 4 13 1 15 10 0 9 7 9 2 13 2 11 2 15 1 1 10 0 9 2 16 15 13 9 16 15 13 9 2 7 9 13 1 0 9 2
10 1 13 15 0 10 10 9 7 9 2
6 7 3 2 10 9 2
4 15 13 12 2
16 12 9 4 13 16 9 13 9 2 3 12 9 1 11 9 2
20 10 9 1 9 1 11 13 10 9 0 2 13 1 11 2 11 11 11 2 2
9 10 9 13 15 10 9 1 9 2
6 0 11 13 1 9 2
13 0 13 15 0 16 15 4 13 10 0 0 9 2
13 9 1 2 11 2 13 3 9 1 10 0 9 2
27 9 13 1 9 2 7 3 4 15 13 2 10 10 9 0 1 9 1 9 1 7 1 9 3 13 0 2
11 0 13 9 15 15 13 1 9 1 9 2
21 7 15 13 16 9 9 4 13 14 13 10 0 9 1 10 0 0 9 1 9 2
16 9 1 0 0 9 13 1 9 7 10 0 15 13 1 9 2
7 3 13 9 0 7 0 2
20 9 2 3 2 16 15 3 13 1 15 10 9 7 12 2 7 0 0 9 2
11 1 1 1 12 13 15 0 9 1 11 2
15 3 1 9 13 15 14 13 10 9 15 1 9 4 13 2
30 1 2 11 2 13 15 9 15 13 15 1 1 11 2 9 15 13 15 1 11 2 7 0 1 1 10 9 1 11 2
8 15 4 3 13 14 13 9 2
29 7 10 0 2 0 9 1 0 0 0 9 7 9 2 0 1 10 0 9 1 9 2 4 13 10 0 10 9 2
34 1 9 13 15 9 1 2 3 13 1 2 15 2 2 2 0 1 1 11 9 1 10 0 2 9 16 15 13 14 13 7 13 15 2
3 2 9 2
20 2 13 11 1 11 2 12 9 16 10 0 9 3 4 13 1 9 1 11 2
31 7 3 13 3 0 9 7 10 9 2 1 12 9 16 15 2 7 9 2 15 9 13 0 3 1 2 0 13 1 11 2
28 3 1 9 9 13 15 10 0 9 0 9 14 13 1 10 9 15 3 0 13 14 13 15 1 10 0 9 2
12 1 9 13 2 11 2 10 9 1 0 9 2
8 7 9 13 0 7 0 0 2
10 0 13 9 10 0 0 2 0 9 2
19 9 13 1 9 13 1 9 13 1 9 1 10 0 7 1 10 0 9 2
19 0 1 10 9 9 1 9 1 0 9 2 13 9 1 9 7 0 9 2
12 9 13 1 12 9 2 7 13 3 0 0 2
12 11 11 11 13 14 13 9 1 10 0 9 2
8 1 7 1 13 15 2 3 2
9 15 13 10 0 2 0 1 15 2
15 10 3 0 9 13 9 1 11 11 9 1 2 11 2 2
24 11 13 3 0 16 9 13 2 7 13 15 15 13 1 10 3 0 0 0 7 0 0 9 2
21 9 4 13 9 1 10 9 1 14 13 10 9 16 9 13 9 2 7 9 9 2
9 9 13 16 15 3 13 0 3 2
4 9 13 0 2
9 1 9 11 13 15 10 0 9 2
34 0 1 1 10 0 9 2 13 15 3 10 0 9 1 11 2 11 11 11 2 7 0 11 2 11 11 2 2 15 11 13 3 1 2
10 0 0 13 15 0 14 13 1 9 2
16 2 11 2 4 0 13 2 1 0 9 1 0 2 0 9 2
17 3 0 13 15 0 16 15 3 4 13 1 9 7 9 1 9 2
10 2 8 2 8 8 8 8 8 8 2
5 12 9 1 11 5
7 11 11 2 9 1 11 2
7 11 11 2 9 7 9 2
6 11 11 2 9 11 2
9 11 11 2 9 1 11 7 9 2
12 15 13 11 11 1 9 15 3 4 13 1 2
10 2 8 2 8 8 8 8 8 8 2
18 15 4 3 13 11 11 7 13 15 15 13 1 9 15 4 13 1 2
25 11 13 0 1 14 13 1 9 16 15 13 2 7 1 11 13 10 0 1 11 9 0 1 15 2
39 11 2 7 11 15 15 13 1 11 2 13 1 9 1 15 10 1 9 2 1 9 2 9 2 9 1 9 1 9 1 11 7 9 0 9 1 10 0 2
6 15 13 1 15 10 2
6 7 15 13 3 3 2
14 1 11 12 9 9 13 10 9 0 9 1 10 0 2
20 10 9 13 1 1 14 13 15 2 15 13 1 1 10 9 2 9 7 9 2
18 3 13 15 9 1 15 2 13 15 7 13 1 9 16 15 4 13 2
4 7 9 13 2
16 13 3 0 0 1 16 15 13 10 9 2 0 9 0 9 5
3 11 11 5
46 16 11 11 13 1 9 1 9 9 2 13 15 0 12 9 2 7 10 9 1 0 9 15 13 9 1 9 2 11 2 15 13 3 0 2 2 7 2 3 4 15 13 9 2 2 2
26 3 13 9 1 11 9 2 9 15 13 1 9 10 7 9 11 2 11 2 11 15 13 1 9 10 2
10 13 15 0 1 3 0 9 0 13 2
5 3 13 11 9 2
36 9 15 3 4 13 1 1 1 9 1 11 7 11 2 13 0 15 13 0 0 14 13 1 9 1 9 10 2 9 2 9 7 9 1 9 2
19 2 15 4 3 3 13 15 3 1 9 2 7 15 4 3 3 15 13 2
4 11 11 13 2
14 15 13 1 1 15 15 13 1 2 9 13 1 15 2
6 0 2 0 7 0 2
31 2 13 3 0 0 1 16 15 13 10 9 2 0 9 0 9 2 2 13 11 11 1 10 9 1 11 1 9 7 9 2
11 1 11 13 9 3 3 15 13 14 13 2
6 15 4 0 9 13 2
14 2 15 13 10 3 0 0 9 16 9 3 13 9 2
22 7 16 10 1 15 1 7 1 7 13 9 7 9 2 13 9 11 11 2 11 2 2
55 15 13 1 9 1 15 15 13 13 9 0 9 2 1 9 2 1 9 9 7 1 9 1 9 2 16 15 0 4 13 1 9 1 10 9 13 1 1 11 11 0 9 2 7 0 9 1 9 2 7 1 9 7 9 2
24 2 9 15 3 13 0 0 2 1 9 10 9 9 2 13 0 0 9 1 15 10 1 11 2
8 3 13 15 15 2 13 15 2
20 2 15 15 13 0 9 3 1 9 2 4 0 13 0 7 3 13 0 9 2
15 15 15 13 1 14 13 7 13 0 9 2 13 0 0 2
35 15 13 10 0 9 15 4 13 1 10 0 16 9 4 13 0 0 7 13 16 15 13 0 9 2 13 9 11 11 1 11 9 2 11 2
30 16 11 11 2 11 2 13 10 9 1 10 12 9 2 4 11 11 2 11 2 3 0 13 14 13 15 1 1 11 2
26 15 4 13 1 12 9 2 0 10 1 15 10 7 9 11 11 2 7 10 1 15 10 1 11 11 2
34 11 11 2 11 2 4 13 0 0 2 1 10 9 1 9 1 15 7 9 2 9 9 2 0 9 2 11 7 11 11 15 13 9 2
38 9 11 11 2 11 2 13 3 0 0 2 1 9 1 0 9 13 1 11 2 9 7 9 1 9 15 13 1 9 9 4 13 1 11 1 12 9 2
13 2 13 15 15 13 1 16 11 13 10 0 9 2
5 2 15 13 15 2
16 15 13 3 0 14 13 15 1 0 9 1 16 15 13 0 2
15 15 13 1 3 9 1 15 10 13 7 3 15 4 13 2
22 1 9 13 15 10 9 1 11 13 10 0 0 9 1 9 1 9 15 13 1 9 2
13 15 13 0 9 1 0 9 2 13 9 11 11 2
13 11 13 15 13 0 9 1 3 0 9 4 13 2
36 15 13 3 3 10 9 1 14 13 16 9 3 13 1 9 2 7 13 16 15 13 14 13 15 0 0 1 15 10 16 15 13 1 10 9 2
8 15 4 1 10 13 0 9 2
13 2 15 4 0 13 10 9 1 11 1 0 9 2
23 3 4 15 13 9 14 13 15 0 1 16 15 13 1 14 13 1 15 15 4 13 0 2
12 9 13 1 7 1 3 0 2 3 1 9 2
13 10 9 1 11 13 1 14 13 1 0 9 9 2
24 2 10 9 1 9 11 2 2 13 11 11 2 11 2 2 7 13 1 9 1 9 11 9 2
17 2 11 2 2 13 11 11 2 11 2 1 10 9 1 9 11 2
39 2 10 9 2 9 2 9 2 9 2 10 9 2 10 9 2 8 8 8 8 8 8 2 2 13 9 1 11 11 2 11 2 1 10 9 1 9 11 2
19 9 11 11 2 11 2 13 12 9 1 10 9 1 15 10 0 1 9 2
18 2 15 13 7 13 1 15 16 11 13 15 1 1 9 1 9 9 2
14 3 9 1 9 4 13 13 15 3 3 13 15 1 2
3 0 2 2
11 2 9 1 15 15 13 1 9 4 13 2
4 15 13 15 2
12 2 15 4 3 0 13 10 0 9 1 9 2
10 0 9 13 3 0 1 1 10 9 2
23 15 4 3 3 13 1 10 9 16 9 13 0 0 1 14 4 13 2 13 9 11 11 2
14 2 13 15 10 9 0 0 1 14 13 0 1 0 2
12 2 15 13 3 1 16 15 13 14 13 9 2
9 0 13 1 1 14 13 0 0 2
20 7 15 13 0 16 15 13 0 0 2 16 1 7 1 9 13 16 9 13 2
18 15 4 3 13 16 9 7 9 13 0 0 0 10 9 1 10 9 2
15 9 11 13 9 1 11 13 3 10 10 1 11 7 11 2
27 2 15 13 3 10 0 9 2 3 16 11 4 0 0 13 1 14 13 1 9 7 3 13 0 0 0 2
9 13 15 1 15 9 13 1 9 2
8 15 13 15 15 3 1 11 2
6 2 0 9 1 11 2
11 11 11 13 3 0 16 15 3 13 9 2
59 13 0 9 1 9 1 3 2 2 13 9 11 11 11 2 11 2 1 10 9 1 15 10 7 9 11 11 1 9 2 16 11 11 2 11 2 13 1 9 1 15 10 1 9 1 11 11 2 1 0 9 2 9 1 9 7 0 9 2
26 2 9 13 15 1 9 7 9 2 2 13 11 11 11 2 11 2 1 9 1 15 10 7 10 9 2
15 12 9 1 11 1 11 4 13 9 1 14 13 0 9 2
44 2 9 1 14 13 13 0 2 7 9 15 13 0 1 0 9 13 0 0 0 1 14 13 9 1 15 15 13 0 0 2 13 9 11 11 1 11 1 11 7 11 2 11 2
12 15 13 9 1 14 13 13 10 9 1 9 2
19 2 10 9 13 1 16 15 13 15 14 13 1 0 1 0 0 0 9 2
34 9 13 16 9 3 4 13 3 16 15 13 16 15 13 1 9 2 7 16 9 3 13 1 9 16 15 13 1 15 15 13 1 9 2
18 15 13 0 7 0 0 9 1 10 9 1 9 16 15 13 0 9 2
20 0 4 11 11 7 9 11 11 13 9 1 14 13 9 1 12 9 1 11 2
18 1 9 13 15 14 4 13 9 1 9 1 9 7 9 1 10 9 2
24 2 9 10 13 1 16 11 1 15 10 13 1 1 14 13 9 1 15 15 4 13 1 10 2
12 7 10 10 13 3 11 7 11 2 13 11 2
25 9 13 9 0 4 13 15 16 15 13 1 9 2 3 13 15 1 10 9 1 15 15 13 0 2
30 1 0 9 13 15 1 0 9 0 9 7 3 3 0 9 1 9 15 15 0 13 1 10 9 2 1 9 1 9 2
15 11 13 9 13 1 10 10 9 1 10 9 1 0 9 2
6 15 13 3 3 0 2
18 2 7 15 13 3 3 9 7 10 9 15 13 0 1 9 7 9 2
5 15 13 1 15 2
24 0 9 13 1 9 0 0 1 3 15 13 1 11 16 9 7 10 9 13 3 2 13 11 2
3 7 0 2
9 10 9 7 15 13 1 14 13 2
25 7 15 13 3 1 11 1 9 2 7 3 4 15 13 1 11 16 15 13 15 2 13 11 11 2
6 2 11 13 10 9 2
13 3 13 15 1 9 1 9 15 13 0 7 0 2
10 15 13 10 0 10 1 11 7 11 2
20 2 13 15 1 9 1 14 13 10 10 9 1 15 10 2 10 10 1 11 2
17 2 15 13 3 1 9 1 15 10 2 7 15 13 3 11 0 2
13 15 13 0 9 2 10 9 16 15 13 0 9 2
13 15 13 10 3 0 0 9 16 9 3 13 9 2
14 7 16 10 1 15 1 7 1 7 13 9 7 9 2
13 15 13 15 3 1 10 9 16 10 9 4 13 2
16 2 13 15 0 1 16 10 1 15 15 13 1 4 4 13 2
20 2 15 13 3 9 1 9 7 15 13 3 1 15 15 13 0 1 14 13 2
14 2 0 9 1 11 13 3 16 15 4 13 14 13 2
18 15 4 3 3 13 15 3 1 9 2 7 15 4 3 3 15 13 2
25 16 15 13 16 15 1 10 4 13 1 9 1 15 7 9 2 13 15 16 15 13 0 1 9 2
10 2 10 9 7 15 13 1 14 13 2
23 7 15 13 3 1 11 1 9 2 7 3 4 15 13 1 11 16 15 13 15 2 6 2
15 2 15 13 3 0 1 11 7 15 13 3 15 13 11 2
18 13 15 9 1 9 7 13 15 0 1 14 13 1 9 1 0 9 2
14 15 13 3 0 1 1 9 7 15 13 10 0 9 2
9 2 13 15 15 15 3 13 1 2
27 2 15 13 16 15 13 15 15 3 13 1 1 10 9 3 2 7 13 0 1 14 13 1 9 1 10 2
6 3 13 15 0 9 2
11 4 13 16 15 1 9 13 9 1 11 2
10 15 13 3 3 1 9 1 0 9 2
14 1 9 4 15 13 10 1 9 2 7 3 3 0 2
18 2 7 15 4 13 1 9 1 10 9 7 1 11 11 7 11 11 2
22 2 6 2 15 13 3 12 1 10 9 2 15 3 13 1 11 7 13 1 1 10 2
11 15 13 1 10 9 1 11 1 0 9 2
19 13 15 13 0 0 14 13 9 1 10 10 9 16 15 13 9 1 9 2
15 2 13 15 1 9 1 14 13 10 10 9 1 15 10 2
11 2 15 13 3 3 0 7 0 1 15 2
15 11 13 10 0 9 14 13 1 1 15 10 13 0 1 2
16 2 13 15 0 1 16 10 1 15 15 13 1 4 4 13 2
27 2 6 2 15 13 14 13 0 1 9 1 15 15 13 7 15 13 3 3 0 1 16 15 4 4 13 2
15 1 11 13 15 9 1 9 15 3 3 13 1 9 1 2
8 15 13 10 0 9 1 15 2
17 2 15 13 1 9 1 15 15 13 2 16 15 13 1 9 3 2
11 15 13 3 1 9 1 9 7 0 9 2
11 15 13 3 3 0 1 15 15 13 1 2
18 15 13 3 3 1 9 2 7 15 4 3 3 13 1 1 10 9 2
10 15 13 15 3 1 9 1 9 10 2
8 15 13 3 0 9 1 9 2
18 2 15 4 13 1 11 11 1 9 2 1 9 1 9 11 5 11 2
15 2 15 13 3 9 7 15 13 10 9 1 15 13 15 2
11 15 13 3 10 9 15 4 13 0 9 2
6 4 3 13 10 0 2
22 15 4 3 3 13 10 0 9 15 13 2 15 13 3 0 1 9 10 1 10 9 2
10 2 13 15 15 15 3 4 13 1 2
10 2 15 13 3 1 9 1 15 10 2
14 0 13 1 9 1 9 7 9 10 7 10 0 9 2
7 15 13 3 11 1 9 2
16 2 13 15 0 1 16 10 1 15 15 13 1 4 4 13 2
13 2 6 2 7 15 13 3 1 15 15 13 0 2
14 7 15 4 3 13 0 0 16 15 4 13 9 3 2
19 13 1 9 1 9 1 11 9 11 2 11 2 11 2 11 11 2 3 2
9 11 2 11 7 11 13 1 15 2
11 11 13 16 9 13 2 8 8 8 2 2
18 2 15 13 10 0 9 2 7 15 13 15 7 13 3 2 13 11 2
13 2 1 11 13 10 0 3 1 15 2 13 11 2
12 2 15 4 13 10 9 15 13 1 10 9 2
18 7 15 13 1 0 9 2 7 4 13 0 1 9 1 14 4 13 2
10 3 2 15 4 13 15 2 13 11 2
23 10 0 9 13 14 13 15 1 1 9 11 11 1 14 13 3 15 4 13 1 9 1 2
10 11 13 9 11 11 2 7 9 11 2
7 2 13 15 13 15 0 2
12 11 2 15 4 3 13 15 0 2 13 11 2
11 15 13 3 15 15 4 13 1 9 10 2
28 2 9 1 10 9 1 12 9 4 13 0 7 0 2 13 11 2 15 13 16 15 4 13 3 1 10 9 2
17 2 1 9 1 10 10 9 13 15 0 9 1 11 2 13 11 2
17 11 4 13 1 2 13 11 2 7 13 16 9 1 4 13 0 2
28 2 15 13 1 11 0 9 0 0 7 0 0 1 3 1 14 13 3 1 9 15 4 13 0 2 13 11 2
31 11 13 16 11 4 13 10 9 16 15 2 0 1 9 2 9 2 0 9 7 10 9 4 4 13 9 0 1 0 9 2
17 2 15 13 3 10 9 0 7 0 9 2 15 13 11 0 9 2
19 11 11 4 13 1 9 1 11 9 1 11 1 9 16 15 4 13 9 2
16 11 11 7 9 11 7 11 4 13 3 1 15 2 1 11 2
22 11 11 13 10 0 9 1 11 0 9 1 0 14 4 13 0 9 1 10 0 9 2
20 11 13 9 11 2 11 2 11 11 2 11 2 11 2 11 2 11 7 11 2
20 1 9 13 15 3 1 14 13 10 0 9 11 2 15 3 4 0 13 3 2
16 11 11 4 13 0 1 10 9 1 14 4 13 11 10 9 2
22 10 12 9 11 13 14 13 1 1 9 13 11 7 11 2 12 0 0 0 0 9 2
22 11 4 13 11 11 1 9 1 11 12 9 2 15 15 13 15 12 1 11 11 12 2
14 3 13 15 3 11 15 3 4 4 4 13 1 11 2
20 1 11 13 11 9 1 16 10 0 9 4 13 1 9 1 14 13 10 9 2
16 2 8 8 8 2 2 12 0 9 2 13 15 0 1 9 2
22 1 9 1 11 13 11 11 3 16 15 4 13 9 11 11 1 14 13 15 1 9 2
9 3 13 15 0 16 11 13 9 2
26 11 13 9 7 9 11 11 2 15 15 13 10 9 3 0 9 2 3 1 9 1 11 11 1 9 2
11 2 11 4 13 10 0 9 2 13 11 2
18 11 13 1 16 15 13 10 0 9 1 11 2 1 0 9 1 9 2
21 2 9 4 13 10 10 9 1 15 2 7 15 7 11 13 1 15 2 13 11 2
11 1 11 9 1 11 13 15 1 11 9 2
12 15 4 13 16 11 3 0 4 13 1 9 2
12 1 9 9 1 11 2 13 15 3 1 11 2
19 10 0 0 9 4 13 9 1 10 10 0 9 2 1 11 1 12 9 2
11 11 11 13 1 0 12 0 1 11 11 2
22 1 12 9 1 9 0 1 2 13 15 1 16 3 10 9 4 13 1 10 0 9 5
11 11 13 0 9 1 9 1 14 13 9 2
14 14 13 10 0 9 4 15 13 2 13 9 11 11 2
18 9 11 11 1 11 13 10 0 0 0 9 2 1 11 11 11 9 2
11 11 13 3 3 11 11 1 9 1 11 2
25 1 9 12 9 2 13 11 1 12 9 2 12 1 11 2 1 12 1 11 11 2 1 11 9 2
17 9 13 1 0 9 2 7 3 3 13 11 11 3 1 9 9 2
23 11 11 11 13 16 11 9 4 13 16 9 1 11 2 11 0 0 9 2 4 13 1 2
12 11 13 12 9 1 11 12 9 0 1 9 2
8 9 4 3 3 13 1 11 2
21 7 9 12 9 2 15 4 13 14 13 1 9 2 4 3 13 15 1 7 1 2
18 9 11 11 11 13 3 11 11 1 9 1 9 11 2 12 9 2 2
16 1 12 9 1 9 0 2 13 11 1 12 9 1 10 9 2
31 9 4 13 11 1 9 1 9 2 1 0 14 4 13 1 10 0 9 2 7 13 11 13 12 0 9 1 12 1 11 2
29 3 4 9 3 13 10 9 1 11 7 11 2 16 15 13 11 13 0 3 2 7 1 11 16 11 13 0 3 2
12 0 13 11 11 1 12 0 9 1 11 11 2
27 9 1 11 13 3 16 10 0 9 13 1 1 14 13 0 9 2 7 3 13 0 9 1 11 0 9 2
15 11 13 3 16 11 11 13 9 11 2 15 13 12 9 2
6 15 13 11 12 9 2
15 3 1 11 12 2 13 11 3 1 10 0 9 1 12 2
12 11 13 3 11 11 1 9 1 11 12 9 2
21 11 11 4 3 13 15 12 9 2 7 13 3 1 14 13 0 1 10 0 9 2
12 15 13 1 1 11 2 11 2 11 7 11 2
24 1 0 4 11 13 1 1 0 9 1 9 2 7 3 3 13 15 1 1 14 13 1 11 2
15 9 13 3 10 9 1 12 9 1 12 9 1 9 0 2
17 1 11 13 12 9 1 9 0 2 7 11 9 13 0 3 3 2
30 11 13 16 9 1 11 11 9 3 13 0 1 14 13 9 2 16 15 13 16 15 15 13 11 3 3 4 0 13 2
34 12 9 1 9 4 13 1 1 11 2 7 3 16 15 3 13 12 9 1 12 9 1 11 1 11 2 13 11 16 11 4 13 9 2
27 3 9 11 11 13 11 9 2 1 12 9 2 7 13 16 11 11 3 3 4 13 0 1 7 13 9 2
29 15 15 13 9 11 2 12 9 2 2 11 2 12 2 2 11 2 12 2 7 11 2 12 2 13 3 3 0 2
19 7 3 1 15 13 11 2 11 7 0 10 9 16 11 13 1 12 9 2
5 11 2 11 2 2
20 2 15 13 11 11 2 15 13 9 10 2 13 11 11 1 11 9 1 11 2
8 15 4 13 1 11 1 12 2
10 1 11 13 10 9 3 0 1 0 2
7 2 15 4 13 3 0 2
5 15 13 1 9 2
16 15 13 10 0 9 1 15 15 4 13 1 15 2 13 11 2
33 9 11 11 11 13 16 9 9 13 16 11 11 13 9 2 7 13 3 3 2 1 10 0 9 1 12 1 11 1 12 1 11 2
5 11 2 11 2 2
17 9 1 11 9 1 11 13 3 16 11 13 16 11 4 13 9 2
12 9 13 7 13 1 9 2 13 7 13 15 2
10 1 9 13 9 2 11 8 11 2 2
22 7 11 7 11 13 3 11 11 1 9 2 1 16 15 13 9 1 10 0 9 11 2
10 3 11 13 11 9 2 1 12 9 2
8 3 13 9 16 11 13 11 2
8 11 13 3 16 11 13 9 2
12 11 12 9 13 0 1 11 11 2 13 11 2
6 15 13 11 12 9 2
8 15 13 3 3 12 1 12 2
11 11 13 3 16 11 11 13 11 12 9 2
14 1 9 13 9 16 15 4 13 11 11 2 12 2 2
23 15 13 15 10 9 1 12 0 9 2 3 12 1 10 0 9 12 15 13 1 14 13 2
11 11 13 1 3 12 9 2 1 11 9 2
13 11 9 13 3 16 11 4 13 10 9 1 11 2
13 9 13 16 11 4 13 1 12 9 1 9 12 2
21 1 9 13 12 0 15 4 13 14 13 1 11 2 7 12 15 3 3 13 0 2
20 11 13 3 16 11 11 13 11 12 9 2 9 11 12 9 7 9 11 12 2
12 11 9 13 3 16 11 13 11 2 12 2 2
17 11 13 3 16 11 13 11 2 12 2 2 7 11 2 12 2 2
13 9 11 13 3 16 11 0 13 11 2 12 2 2
6 10 10 13 3 11 2
13 11 13 3 16 11 13 12 9 2 1 11 12 2
13 3 12 9 1 9 1 11 4 3 3 13 1 2
20 3 13 15 0 0 2 7 11 13 1 12 9 1 11 12 9 2 1 11 2
8 11 4 13 9 10 0 9 2
11 3 12 9 9 4 3 13 1 1 11 2
13 1 11 9 4 11 11 13 11 7 9 12 9 2
22 9 13 0 16 11 11 13 3 1 14 13 10 12 9 1 11 2 8 11 11 8 2
7 11 7 11 13 10 10 2
12 10 0 9 1 11 9 1 11 13 1 9 2
12 9 13 1 16 15 13 15 1 9 7 13 2
19 3 12 9 13 11 7 11 1 11 1 12 9 1 9 0 2 1 11 2
13 11 13 1 12 9 1 11 12 1 10 0 9 2
10 0 12 9 9 4 13 1 1 11 2
15 11 13 0 3 1 10 0 9 2 3 0 1 9 11 2
28 16 11 11 13 1 9 2 4 15 3 13 1 10 9 15 13 1 12 2 1 9 2 11 11 13 0 2 2
27 16 12 9 1 9 4 13 1 1 11 2 9 1 9 11 11 2 13 11 7 11 1 12 1 12 9 2
27 11 13 15 13 3 0 14 13 10 9 1 11 2 16 11 7 11 3 4 13 11 1 0 9 1 9 2
17 1 10 9 1 9 0 1 11 13 11 1 0 12 9 1 9 2
10 11 13 3 12 9 1 9 3 0 2
9 9 1 11 13 1 3 12 9 2
20 11 11 13 0 1 11 11 1 9 0 9 2 1 10 0 2 0 9 9 2
13 7 0 13 0 0 9 1 11 2 11 7 11 2
14 11 13 0 9 1 10 9 2 1 0 12 1 12 2
10 11 13 12 2 7 9 11 12 9 2
9 1 10 9 13 9 12 0 9 2
18 1 10 0 9 11 13 11 3 1 1 12 9 1 9 1 11 12 2
11 12 9 1 9 4 3 13 1 1 11 2
12 1 11 13 15 9 1 0 0 9 1 1 2
21 1 10 4 3 0 9 1 9 13 1 10 0 0 9 11 2 15 13 0 0 2
14 0 1 10 0 0 9 1 1 3 13 12 9 0 2
16 15 13 16 11 4 13 10 0 9 1 14 13 9 1 11 2
11 11 11 13 1 1 14 13 9 1 11 2
35 9 11 13 0 16 15 13 16 9 13 0 9 1 14 2 13 1 0 9 2 16 15 13 0 1 14 4 4 13 1 2 0 9 2 2
30 15 4 13 1 10 0 9 1 9 1 11 2 15 3 1 10 0 9 3 13 0 1 14 13 9 1 11 0 9 2
14 11 13 3 16 11 11 4 13 11 7 9 12 9 2
10 9 13 0 0 2 1 10 0 9 2
30 1 11 2 11 7 11 4 9 3 13 2 7 9 13 15 13 3 0 14 13 1 9 1 15 15 4 13 10 9 2
19 3 11 9 13 16 11 13 11 2 7 9 13 3 16 9 4 13 11 2
9 3 11 13 11 13 11 7 11 2
19 15 4 13 16 0 1 10 0 9 4 13 1 0 9 9 12 0 9 2
13 9 11 13 3 11 1 0 9 1 9 11 11 2
5 9 13 12 9 2
14 11 11 13 1 1 14 13 11 0 0 9 1 11 2
20 15 13 16 11 13 1 11 11 9 2 15 15 13 16 15 13 1 9 12 2
19 11 2 11 2 11 7 11 13 16 11 11 13 11 2 7 9 12 9 2
25 9 11 9 13 3 16 11 11 13 3 1 14 13 11 2 1 16 12 9 1 9 4 13 1 2
5 9 13 12 9 2
14 9 13 3 1 1 9 11 1 12 1 11 12 9 2
10 1 11 4 12 9 1 9 13 1 2
5 9 13 12 9 2
16 11 13 16 11 3 13 1 9 11 2 1 12 1 12 9 2
7 11 13 3 12 9 1 2
20 1 11 13 15 0 0 9 2 12 2 12 2 16 12 9 9 4 13 1 2
9 11 13 3 12 9 1 1 9 2
19 9 11 10 9 13 3 16 11 11 13 3 1 14 13 11 11 12 9 2
15 11 13 16 11 11 13 12 0 9 2 1 12 1 11 2
11 11 13 12 1 11 2 1 12 1 11 2
17 1 12 9 1 9 0 1 11 13 15 0 9 1 11 7 11 2
21 15 4 13 1 0 12 9 9 2 7 15 13 3 0 12 9 1 10 0 9 2
21 1 11 13 11 3 1 12 1 12 9 2 1 16 12 9 1 9 4 13 1 5
23 11 13 9 12 16 11 4 13 9 1 11 9 2 15 15 13 9 1 1 9 1 12 2
21 3 4 0 9 3 4 13 1 0 9 7 0 9 1 10 12 9 1 0 9 2
22 15 13 3 3 0 14 13 16 11 4 13 10 9 1 11 2 10 10 9 1 11 2
5 11 9 1 11 2
4 3 13 15 2
13 16 11 13 11 9 1 11 2 13 9 1 9 2
13 2 15 13 0 2 13 9 11 11 1 11 11 2
15 15 13 11 0 4 13 10 0 9 2 16 15 4 13 2
12 2 3 13 15 9 1 14 13 10 0 9 2
17 15 13 3 15 4 13 15 11 4 13 3 2 13 15 1 8 2
25 11 13 11 11 1 9 1 11 2 12 9 2 2 11 11 2 12 2 7 11 11 2 12 2 2
9 0 12 0 9 1 10 0 9 2
45 10 9 13 11 11 1 9 1 11 2 12 2 2 11 2 12 2 2 11 2 12 2 2 11 11 2 12 2 2 11 11 2 12 2 2 11 2 12 2 7 11 2 12 2 2
33 1 9 13 11 16 11 4 13 12 1 12 9 1 11 2 15 13 10 9 1 10 10 9 1 10 0 9 2 16 9 13 15 2
7 0 12 0 9 1 11 2
7 11 11 11 13 1 11 2
32 10 0 9 9 15 13 14 13 15 1 11 9 1 11 13 1 9 16 11 13 10 0 9 1 9 1 10 0 0 9 11 2
23 11 11 13 10 1 11 0 9 0 2 7 4 13 0 9 1 0 9 1 9 1 9 2
14 1 9 1 9 13 15 1 9 1 9 9 1 11 2
19 2 0 1 9 15 4 13 1 1 9 2 13 15 0 1 16 15 13 2
26 15 4 13 1 9 1 9 2 3 16 15 13 0 1 14 4 13 9 1 10 0 9 2 13 11 2
20 1 0 9 13 15 3 0 0 9 1 14 13 2 1 10 1 11 7 11 2
10 1 11 13 3 9 1 1 10 9 2
12 15 13 3 1 14 13 9 1 9 0 9 2
18 16 15 13 1 9 16 9 0 13 2 13 15 9 1 14 4 13 2
24 1 10 9 13 9 1 0 9 2 1 10 9 11 7 1 11 2 9 1 9 9 11 11 2
20 9 4 13 16 11 4 13 9 0 2 7 1 10 0 9 1 9 13 9 2
28 1 9 13 9 1 11 2 11 11 2 11 2 11 2 11 2 11 11 7 1 9 1 11 11 7 11 11 2
7 11 13 11 2 13 11 2
9 9 4 1 9 13 1 0 0 2
10 9 11 11 13 1 11 9 1 11 2
4 9 3 3 2
16 15 4 13 1 9 1 9 7 9 15 3 13 1 1 9 2
14 9 1 9 15 3 13 1 2 7 9 4 13 3 2
18 1 9 15 3 13 0 0 2 13 11 11 1 12 1 12 1 11 2
4 13 15 0 2
20 3 1 9 13 15 1 9 7 11 2 7 15 4 13 9 1 11 11 11 2
14 9 1 11 13 11 9 1 12 1 12 2 1 11 2
25 15 13 10 9 9 13 4 13 1 9 2 7 3 0 13 15 1 1 16 11 13 9 1 9 2
5 9 13 12 9 2
29 11 13 3 16 11 11 4 13 1 11 2 12 2 2 11 2 12 2 2 11 2 12 2 7 11 2 12 2 2
14 15 13 9 15 1 9 4 13 1 0 9 1 9 2
18 10 9 13 16 11 11 13 1 12 9 1 10 9 1 9 11 11 2
22 1 11 2 16 12 9 1 9 3 4 13 1 2 13 11 1 1 12 9 1 12 2
28 11 9 13 3 16 11 11 4 13 0 9 1 9 2 3 16 11 3 13 12 0 9 1 12 1 11 11 2
59 9 11 13 11 4 13 13 11 2 12 9 2 2 9 11 11 9 11 2 12 2 2 11 11 2 12 2 2 11 9 11 2 12 2 2 11 2 12 2 2 11 2 15 13 9 1 11 11 2 2 12 2 7 11 11 2 12 2 2
33 1 11 2 16 9 13 1 10 10 9 1 10 0 10 9 2 16 9 13 15 2 13 11 9 16 11 4 13 12 1 12 9 2
12 0 13 9 16 11 11 4 13 11 12 9 2
11 3 13 9 1 12 9 2 1 15 11 2
30 11 4 13 1 9 1 11 2 7 9 4 1 9 1 9 13 0 1 1 14 13 14 13 1 1 10 0 0 9 2
10 3 1 11 13 9 9 12 0 9 2
13 0 13 15 12 9 1 10 12 9 7 11 11 2
19 1 9 15 3 13 3 0 2 13 11 11 1 12 1 11 12 1 11 2
20 11 12 9 13 1 10 0 0 0 9 11 11 2 11 11 2 11 7 11 2
18 1 11 13 3 11 11 1 12 9 1 12 9 1 11 11 1 11 2
16 12 9 1 9 4 3 13 1 2 7 11 13 1 12 9 2
19 11 13 3 11 11 1 9 1 11 11 2 10 9 15 13 1 0 0 2
16 1 9 13 15 3 1 16 11 11 13 10 0 0 9 11 2
13 1 9 13 11 12 9 2 1 12 9 1 11 2
10 11 13 11 11 1 9 1 11 11 2
5 9 13 12 9 2
18 1 11 11 13 9 9 16 15 13 0 9 2 12 9 1 12 9 2
20 11 11 2 9 1 11 1 0 9 2 13 11 13 9 2 1 12 0 9 2
22 2 9 13 16 10 9 15 4 13 1 9 1 9 0 13 1 1 9 2 13 11 2
18 10 0 9 13 0 0 2 0 7 0 0 1 1 0 10 0 9 2
19 15 13 15 0 1 9 14 13 16 0 9 0 13 1 1 9 7 3 2
31 15 4 3 13 16 9 7 9 1 11 4 13 0 9 1 10 0 9 2 9 15 3 3 13 15 1 14 13 1 9 2
33 2 15 4 3 13 1 1 1 16 9 3 4 13 1 14 13 9 15 3 4 13 14 13 1 1 9 1 0 9 2 13 11 2
14 9 12 2 0 9 2 13 9 1 10 0 9 11 2
28 0 13 9 1 11 11 2 15 9 13 14 13 1 1 11 2 7 11 11 2 15 13 1 10 0 0 9 2
8 0 13 10 12 9 12 9 2
27 0 9 1 11 2 16 12 9 1 9 4 13 1 2 13 1 11 16 9 3 13 12 9 1 12 9 2
6 11 13 1 12 9 2
13 12 9 1 9 4 13 1 1 11 2 13 11 2
17 0 13 11 1 12 9 1 10 0 9 2 1 12 9 1 11 2
18 11 13 12 9 2 7 16 3 11 13 14 13 9 4 9 0 13 2
23 7 3 4 3 10 9 1 9 13 2 7 15 13 3 3 12 9 1 9 15 4 13 2
6 11 13 11 1 12 2
16 15 13 1 9 0 9 3 9 1 0 9 1 9 1 11 2
16 1 11 13 9 3 0 2 16 9 13 14 13 9 1 9 2
26 1 0 9 4 9 4 13 1 1 1 12 9 1 9 2 13 11 2 7 12 9 2 1 11 11 2
19 1 11 13 9 1 11 0 9 1 11 7 11 2 12 9 1 12 9 2
20 9 13 3 16 11 0 13 11 2 7 11 1 9 1 11 2 12 9 2 2
14 3 11 11 11 10 9 13 16 11 13 11 12 9 2
17 9 12 13 9 1 12 9 2 15 1 3 13 12 1 12 9 2
27 9 13 9 11 7 11 2 10 0 0 0 9 11 2 11 7 11 11 2 7 10 0 0 0 9 11 2
31 15 13 3 0 1 12 9 1 9 15 4 13 1 2 7 11 11 11 4 13 10 0 9 1 11 11 1 9 11 11 2
13 3 3 4 12 9 1 10 0 9 13 1 11 2
15 9 12 13 9 1 12 9 2 1 15 10 0 9 11 2
24 16 11 3 13 14 13 9 12 9 2 13 9 10 1 14 13 9 1 11 0 9 0 0 2
8 11 13 0 9 1 1 9 2
19 0 13 12 9 16 11 11 13 0 0 1 14 13 9 2 12 9 11 2
23 1 9 1 15 15 13 0 1 9 1 9 1 15 2 13 12 9 11 2 12 9 11 2
23 1 11 4 15 0 3 13 14 13 10 9 1 10 0 0 9 11 1 9 2 0 9 2
7 15 13 9 12 0 9 2
5 11 13 12 9 2
12 10 0 9 13 14 13 1 1 11 7 11 2
29 3 13 15 3 0 0 9 15 4 13 1 2 7 1 11 13 11 11 1 0 9 1 12 9 2 1 11 11 2
8 1 11 13 11 1 12 9 2
12 15 4 1 9 13 16 11 4 13 10 9 2
13 1 11 4 11 11 13 1 10 9 1 14 13 2
6 7 2 15 15 13 2
20 1 9 2 3 13 10 9 1 10 1 10 0 9 2 9 15 13 0 9 2
8 10 0 9 13 0 1 9 2
14 15 13 16 9 13 10 0 9 1 10 9 1 9 2
24 1 15 15 13 16 9 13 0 2 13 12 9 1 9 7 12 9 1 9 1 10 0 9 2
21 11 4 13 10 0 9 1 11 11 11 1 11 11 1 14 13 15 15 13 9 2
22 3 13 15 0 2 1 9 2 1 12 9 2 7 0 2 1 9 2 1 12 9 2
22 16 9 13 0 1 13 15 15 13 9 2 4 9 1 10 0 9 13 0 7 0 2
13 1 11 13 11 11 15 14 13 10 9 7 13 2
25 9 13 1 11 2 15 13 10 0 0 9 2 7 13 1 11 2 10 9 9 1 10 9 13 2
21 1 15 15 3 13 0 1 14 13 1 7 11 7 11 2 13 11 10 0 9 2
5 11 11 1 9 2
9 15 13 1 11 0 11 1 9 2
7 9 11 11 13 9 10 2
10 15 13 14 13 1 11 9 11 11 2
12 15 13 3 15 15 13 1 3 2 14 13 2
15 10 0 9 4 13 9 0 9 2 1 9 11 7 11 2
17 10 9 13 1 0 9 1 9 2 3 16 11 13 11 1 12 2
20 11 13 16 1 12 9 4 13 1 10 9 16 9 4 13 1 1 0 9 2
13 9 4 1 10 13 1 11 7 11 2 0 9 2
25 11 13 3 1 16 10 9 4 13 1 16 10 9 13 10 9 1 11 1 1 10 9 1 11 2
22 9 1 0 9 2 7 0 1 11 2 0 2 13 1 14 13 10 0 9 1 9 2
6 7 15 13 3 9 2
17 11 11 11 11 12 9 1 11 11 11 13 7 0 7 0 0 2
2 9 2
14 15 13 12 9 15 13 0 14 13 1 1 1 9 2
23 11 2 12 9 2 2 11 11 2 12 2 2 11 11 2 12 2 7 11 2 12 2 2
21 11 11 4 1 9 13 11 2 11 7 11 11 1 14 13 10 9 1 14 13 2
18 11 11 13 0 10 0 0 9 2 7 11 13 14 13 15 1 12 2
15 3 13 10 0 9 16 15 13 10 0 0 9 1 11 2
14 0 9 1 11 13 16 9 13 0 1 9 1 0 2
15 15 13 0 1 11 14 13 15 1 12 1 9 12 9 2
15 11 13 11 9 1 11 1 9 11 11 7 9 11 11 2
13 0 1 9 13 9 11 11 2 15 13 1 11 2
18 9 13 1 0 9 1 10 10 2 7 16 0 9 3 13 14 13 2
7 15 13 3 1 11 11 2
19 3 13 15 1 10 12 9 0 11 11 2 15 4 13 1 9 1 11 2
10 10 0 9 13 1 9 12 0 9 2
8 1 15 13 10 0 9 11 2
18 11 4 13 10 9 12 9 2 4 15 13 10 9 1 14 13 9 2
20 11 13 11 1 12 2 7 9 13 0 1 9 15 11 13 1 12 7 12 2
12 1 9 4 15 13 0 0 1 9 1 9 2
14 11 9 1 0 9 13 11 10 9 1 3 12 9 5
9 10 9 13 3 1 10 0 9 2
32 11 2 11 2 11 13 10 9 1 11 1 12 2 11 11 4 13 1 9 1 11 2 16 11 11 4 13 1 7 13 11 2
22 15 13 3 1 9 1 14 13 11 11 11 2 3 1 11 11 10 0 9 1 11 2
15 9 11 7 11 4 2 15 15 4 13 2 3 13 3 2
7 0 13 1 9 1 9 5
4 9 13 0 5
25 9 10 4 3 13 15 15 13 2 1 11 11 2 10 9 15 13 10 9 9 13 1 1 9 2
20 9 13 1 0 9 2 16 9 1 16 15 13 11 16 15 13 11 13 0 2
9 3 3 0 2 4 3 15 13 2
19 7 9 13 10 0 14 13 3 13 2 13 9 2 1 10 9 1 11 2
22 16 15 13 9 1 11 8 11 2 11 11 7 11 13 15 0 14 13 3 15 13 2
16 7 15 1 9 15 13 0 0 9 2 15 15 13 1 9 2
11 15 13 3 9 1 9 1 9 11 11 2
7 13 9 1 9 1 11 2
10 15 13 1 0 9 1 12 15 13 2
30 10 0 9 4 13 1 1 10 0 9 2 16 12 9 0 1 10 12 9 2 7 11 11 2 13 15 15 13 9 2
20 15 13 0 14 13 9 1 14 13 0 9 2 3 0 15 13 10 0 9 2
22 3 4 15 13 0 1 3 9 13 2 7 3 10 0 9 4 13 15 15 13 9 2
13 9 11 11 13 9 16 15 3 13 1 1 9 2
35 9 11 11 1 11 1 11 11 11 13 11 13 12 9 9 1 9 2 16 9 9 11 11 3 13 12 9 9 1 14 13 2 1 11 2
28 7 2 15 11 10 13 10 0 1 14 13 2 15 13 14 13 1 16 9 13 16 9 1 9 13 12 9 2
10 10 9 13 16 15 3 4 13 9 2
6 0 1 9 1 11 2
23 11 11 4 13 15 1 1 9 7 9 2 7 11 11 11 4 13 1 15 9 7 9 2
31 15 13 1 14 13 1 3 16 15 13 0 15 15 13 9 2 1 0 15 13 10 11 11 1 11 11 9 1 1 12 2
3 0 9 5
15 10 0 9 1 9 15 13 1 10 0 9 9 1 9 5
3 0 9 2
20 9 13 10 0 9 1 14 13 9 10 1 10 0 1 0 9 1 0 9 2
14 11 11 1 11 2 1 9 2 7 11 11 1 11 2
29 11 13 10 0 2 0 0 9 15 13 0 1 9 7 1 2 7 13 3 0 1 9 1 10 9 9 1 9 2
23 16 15 13 9 1 9 1 9 13 15 11 2 10 0 9 1 10 1 11 2 0 9 2
28 11 13 1 9 3 1 9 1 10 9 3 16 15 4 13 16 15 0 13 9 7 3 4 13 14 13 9 2
39 1 10 9 1 0 0 9 13 3 11 15 1 14 13 10 0 0 9 10 9 2 7 3 4 9 13 1 10 9 15 13 10 0 9 1 0 0 9 2
7 7 3 3 15 4 13 2
27 2 11 0 2 13 10 9 3 10 9 1 9 13 9 0 9 1 14 13 0 1 0 0 9 1 9 2
32 9 13 10 9 2 7 0 13 15 0 15 13 15 1 10 1 10 0 9 1 11 11 0 9 2 11 11 11 8 11 2 2
38 1 3 1 10 9 13 9 16 9 4 13 1 10 0 9 7 0 9 10 0 2 7 3 13 14 13 9 7 13 1 1 0 11 2 11 8 11 2
27 9 4 1 10 9 13 9 1 0 9 2 13 15 10 9 1 9 7 13 15 9 1 10 9 0 9 2
30 16 2 11 0 2 1 9 1 15 4 13 1 1 15 1 9 1 10 0 9 13 3 7 0 10 0 7 0 9 2
41 1 10 0 9 1 0 9 7 0 0 9 2 13 15 10 9 1 9 15 0 15 15 13 13 15 1 14 13 16 15 15 13 1 1 9 13 9 1 0 9 2
35 9 13 3 10 0 9 1 14 13 9 10 1 10 0 1 0 9 1 0 9 2 7 13 3 1 14 13 1 1 9 1 9 7 9 2
20 0 13 11 11 2 15 13 0 0 11 11 2 10 0 9 1 9 1 11 2
22 3 4 15 3 13 9 0 9 16 15 13 1 14 13 10 9 1 10 9 1 9 2
33 15 16 11 13 10 1 0 0 9 1 9 1 9 0 9 2 13 2 11 0 2 10 0 9 1 10 9 1 9 0 0 9 2
36 9 9 1 0 9 13 9 1 10 0 9 7 10 0 9 1 9 0 0 9 1 10 9 1 9 7 9 13 1 3 9 10 0 1 0 2
18 16 9 13 10 3 0 0 0 9 3 2 13 3 10 9 1 0 2
30 0 13 15 16 15 13 3 0 1 10 9 1 9 9 16 15 3 1 9 13 0 14 13 1 9 1 10 0 9 2
12 2 11 0 2 13 10 9 15 3 4 13 2
33 3 16 15 4 13 1 10 0 9 2 13 15 3 0 7 0 16 16 15 3 13 15 1 2 13 15 0 9 4 13 10 9 2
42 9 9 13 1 3 9 1 14 4 13 10 9 15 13 3 0 7 0 0 16 15 1 9 1 0 9 3 13 15 13 1 1 14 13 0 7 13 1 10 0 9 2
7 11 13 11 9 1 11 5
2 9 5
4 1 1 9 5
2 13 2
3 11 11 5
9 11 13 11 0 7 0 0 9 2
9 11 13 11 0 7 0 0 9 2
15 3 13 10 0 11 2 9 1 0 9 2 9 7 9 2
12 7 10 12 9 0 9 15 13 9 1 9 2
9 11 2 13 10 0 9 1 11 2
30 15 13 15 14 13 1 3 2 7 16 15 13 1 12 9 4 15 13 1 15 9 7 13 1 10 9 1 12 9 2
11 15 13 1 2 7 13 10 10 10 3 2
34 9 1 9 13 1 0 0 9 7 10 0 9 2 7 13 10 0 9 1 11 0 9 2 15 4 13 1 1 9 1 10 0 9 2
25 11 9 4 13 0 0 7 9 4 13 1 14 13 10 0 2 0 9 1 10 0 0 1 9 2
40 2 1 9 13 15 10 9 2 7 16 15 13 9 4 15 13 9 3 2 13 12 9 0 11 11 11 2 15 13 1 9 9 16 15 13 9 1 0 9 2
7 3 4 15 13 3 0 2
27 1 14 4 13 1 4 15 2 10 0 9 9 7 0 9 2 13 0 9 2 7 3 13 1 0 9 2
14 15 13 1 10 16 10 0 7 0 9 13 9 10 2
25 11 4 13 10 0 9 1 0 9 2 13 13 10 0 9 11 7 10 0 9 2 11 11 2 2
20 9 13 1 0 9 1 14 13 12 9 9 1 11 2 7 13 10 0 0 2
44 10 9 1 1 10 0 9 13 15 9 1 10 0 9 2 15 1 10 0 7 0 9 13 15 3 0 16 15 13 3 1 14 13 1 9 7 9 2 3 1 14 13 1 2
2 6 2
36 1 16 9 0 9 4 13 1 13 15 1 10 9 2 3 1 10 9 9 7 0 0 10 15 4 13 1 14 13 10 9 1 9 0 9 2
45 15 13 1 16 15 13 1 2 3 16 15 13 1 1 9 1 0 9 7 0 9 2 7 3 2 3 1 11 11 11 2 13 15 1 9 10 1 0 9 16 0 9 13 9 2
25 9 1 13 1 9 12 2 1 16 12 9 13 0 1 10 0 9 15 13 0 0 1 15 10 2
42 9 13 0 7 0 2 7 16 11 9 13 14 13 9 2 0 3 1 2 13 15 1 9 1 9 7 3 13 15 2 1 10 9 2 10 9 1 10 0 10 9 2
25 11 4 13 10 0 9 1 0 9 2 13 13 10 0 9 11 7 10 0 9 2 11 11 2 2
20 9 13 1 0 9 1 14 13 12 9 9 1 11 2 7 13 10 0 0 2
37 9 13 10 0 9 1 11 0 2 0 7 0 2 15 13 15 1 1 10 0 9 3 9 13 0 2 9 13 1 2 7 9 9 13 0 0 2
41 2 11 13 10 0 9 9 2 0 1 15 13 0 1 10 9 15 10 0 9 3 4 13 15 9 1 2 13 11 11 2 12 2 15 13 1 1 9 1 9 2
13 7 3 3 3 13 11 10 0 9 14 13 9 2
24 2 9 13 3 1 0 9 2 1 14 13 1 2 1 14 13 2 13 7 13 2 13 11 2
24 10 0 9 13 3 0 1 9 2 7 9 13 0 7 1 9 3 0 1 10 0 9 9 2
11 10 0 2 0 9 13 3 1 10 9 2
33 1 9 1 0 7 0 9 2 13 0 9 0 0 0 2 7 10 0 13 0 16 15 13 10 0 9 15 11 7 11 13 1 2
5 9 3 13 0 2
5 12 9 0 11 2
14 11 13 10 1 0 9 1 11 15 13 9 1 9 2
12 15 13 1 7 1 12 9 13 15 1 9 2
17 9 13 10 0 2 0 9 3 9 13 3 1 9 15 13 1 2
38 9 13 1 10 1 10 0 9 2 9 2 2 7 4 0 13 1 10 9 2 7 10 9 0 9 2 15 15 13 9 16 15 4 13 9 1 1 2
49 9 13 1 9 2 7 1 0 0 9 13 0 9 15 13 1 9 1 9 7 4 13 15 1 0 9 2 9 2 9 7 0 9 9 1 1 9 2 9 2 2 0 9 1 0 2 0 9 2
12 1 13 10 9 3 0 16 15 3 13 9 2
26 9 13 0 2 9 2 16 15 13 9 2 10 0 9 15 13 1 10 0 9 7 13 1 0 9 2
27 10 0 9 11 11 2 3 1 11 9 2 13 3 10 1 10 0 9 15 3 13 10 0 9 1 9 2
23 11 2 15 13 9 1 9 1 9 2 13 11 9 1 11 7 10 0 9 14 13 1 2
32 1 0 2 0 7 0 9 13 11 0 1 0 2 0 9 15 13 9 2 9 7 9 2 9 2 9 1 9 2 7 9 2
27 15 13 3 10 0 9 1 0 2 0 9 2 7 13 3 0 1 9 2 3 9 13 0 7 0 9 2
41 0 11 13 10 0 9 1 9 2 16 10 0 9 13 9 15 13 1 0 9 1 0 9 2 1 1 9 10 0 2 0 9 11 2 15 13 1 1 7 1 2
24 3 13 15 2 9 2 2 0 2 0 9 15 3 13 9 2 7 10 0 0 9 1 9 2
15 16 15 13 11 11 13 15 14 13 9 16 15 13 9 2
15 9 2 9 2 13 10 9 9 1 11 2 7 4 13 2
30 11 11 13 3 1 11 7 13 10 0 9 1 9 15 3 13 0 9 2 0 9 13 16 9 13 9 1 9 2 2
18 16 9 2 9 7 0 9 4 13 3 13 15 3 1 9 1 9 2
52 9 13 15 3 10 9 7 13 3 1 1 8 9 1 0 9 1 9 2 3 11 13 9 12 2 7 15 4 13 1 16 11 3 13 15 0 16 9 13 14 13 9 2 7 15 13 3 2 11 11 2 2
6 9 13 1 11 11 2
2 11 2
4 2 0 0 5
3 9 3 5
2 9 5
11 3 1 9 9 13 11 11 3 10 9 2
13 10 0 9 11 11 11 13 1 11 11 0 9 2
4 9 2 11 5
9 11 11 11 13 1 9 11 11 2
4 9 2 11 5
8 10 0 9 11 11 11 13 2
19 2 15 13 0 0 0 16 10 15 13 2 7 10 9 13 1 10 0 2
11 15 13 0 0 14 13 9 1 10 0 2
17 15 13 3 10 9 2 7 0 13 15 0 0 16 12 9 13 2
29 15 13 0 13 3 9 7 9 15 13 1 9 2 7 16 10 10 1 15 13 13 15 0 10 9 15 13 0 2
20 2 15 13 1 10 9 10 10 9 14 13 9 1 7 15 13 15 0 1 2
14 15 13 3 0 14 13 3 15 4 4 13 1 15 2
24 1 2 0 16 15 13 7 3 2 10 9 13 1 10 0 2 11 11 13 3 11 0 2 2
19 11 11 13 0 7 13 7 13 10 9 1 1 10 0 9 1 12 9 2
6 15 13 15 0 9 2
25 11 4 0 13 1 9 7 13 1 9 1 9 1 11 11 11 2 7 9 13 3 1 14 13 2
11 9 13 1 1 10 0 9 1 10 9 2
5 15 13 1 12 2
30 2 15 4 13 15 2 7 15 13 16 15 15 3 13 15 2 13 15 0 2 2 13 11 11 1 9 10 9 9 2
17 1 9 1 12 4 12 9 13 1 9 1 9 1 10 0 9 2
9 11 13 1 11 11 11 1 11 2
9 15 13 10 0 9 9 1 9 2
4 2 11 2 5
2 9 5
6 0 9 1 0 9 2
5 9 2 11 11 5
45 2 9 7 9 1 11 2 15 13 10 7 10 9 2 15 2 13 10 0 11 11 10 0 9 1 11 1 2 16 9 13 0 1 1 10 0 9 2 7 9 13 9 1 9 2
40 11 11 4 13 9 1 11 9 1 10 9 2 7 15 13 1 7 1 0 9 1 9 16 15 13 11 2 7 2 15 13 3 1 1 16 9 4 13 0 2
27 15 13 0 1 10 9 2 7 4 13 0 9 1 2 11 11 11 11 2 2 7 13 0 9 1 15 2
35 0 0 9 9 14 13 2 7 3 10 0 9 1 0 2 0 9 2 7 9 2 13 0 9 1 0 9 7 0 9 1 10 10 9 2
25 11 9 13 3 0 1 10 9 10 9 2 7 15 13 1 15 7 9 1 10 0 9 1 9 2
48 9 11 11 13 3 10 9 16 15 13 11 0 0 9 2 16 11 11 7 11 11 13 10 0 9 1 9 1 9 1 9 7 12 9 1 14 13 9 2 3 16 9 13 15 10 0 9 2
49 11 11 1 9 13 0 0 1 9 10 9 2 3 0 10 0 9 2 16 10 9 2 15 3 3 13 14 13 9 1 2 13 1 15 1 14 13 0 9 1 2 1 0 0 9 1 14 13 2
43 15 13 0 0 9 1 9 2 7 16 15 13 1 15 15 13 2 4 15 13 1 15 16 15 13 0 0 1 9 1 9 2 7 13 1 10 9 7 13 10 0 9 2
31 15 4 13 0 9 1 1 9 2 7 0 16 9 4 13 1 14 13 1 9 2 13 11 7 9 10 0 9 15 13 2
32 9 14 13 15 13 10 9 15 0 1 2 7 1 10 9 9 1 0 9 2 13 15 14 13 3 1 0 9 7 0 9 2
10 7 15 13 0 9 3 0 15 13 2
12 9 7 11 11 2 15 13 10 9 2 15 2
6 9 11 11 13 0 5
6 2 13 10 0 9 5
5 9 1 11 1 5
4 0 7 0 5
5 13 10 0 9 5
14 11 13 1 10 9 1 10 9 1 11 1 11 9 2
16 1 9 12 4 11 13 9 1 9 1 11 11 9 1 11 2
36 2 9 11 9 13 10 0 9 2 7 1 10 9 7 1 0 11 1 11 2 13 9 11 11 1 10 9 1 9 1 11 0 9 10 9 2
7 2 11 13 10 0 9 2
14 15 4 1 15 13 9 7 1 9 7 1 14 13 2
20 15 13 3 10 0 9 7 9 2 7 13 9 1 10 0 9 7 1 9 2
24 15 13 1 9 0 1 10 9 2 9 2 9 7 9 2 7 13 3 1 15 2 13 11 2
25 9 11 13 1 10 9 10 0 9 1 11 7 11 2 7 4 13 1 9 1 9 1 11 1 2
15 15 13 3 11 11 1 9 1 9 7 13 14 13 9 2
20 2 15 13 10 9 1 14 13 15 10 7 4 13 9 1 14 13 7 13 2
11 9 13 15 1 14 13 1 10 0 9 2
8 15 13 0 1 10 0 9 2
23 11 1 9 13 1 10 0 9 7 13 10 9 2 13 11 1 10 9 1 11 9 12 2
15 0 9 13 15 3 1 1 11 7 13 9 1 1 11 2
6 2 9 13 10 9 2
6 10 9 13 10 9 2
14 10 9 13 16 15 13 0 7 4 13 1 1 9 2
17 15 13 3 3 15 2 7 9 1 15 15 13 13 0 1 9 2
8 15 13 14 13 9 1 9 2
14 0 1 10 9 13 15 9 1 9 2 13 11 3 2
16 11 13 1 1 11 2 13 9 1 11 7 13 9 1 11 2
37 12 9 0 13 15 1 11 0 9 1 14 13 9 2 7 1 10 9 1 9 7 12 9 1 0 9 2 4 15 13 1 9 1 11 1 12 2
9 15 4 13 1 0 9 1 12 2
14 15 4 3 13 0 1 11 2 7 13 1 0 9 2
19 2 1 11 11 9 4 0 9 13 10 1 10 0 9 2 7 0 9 2
18 15 13 10 0 9 1 14 13 15 2 15 13 0 1 10 0 9 2
37 0 13 15 10 0 9 2 0 7 0 7 13 7 13 15 1 10 0 0 2 0 9 1 11 2 13 9 7 9 11 11 11 1 10 0 9 2
20 1 16 9 11 9 13 0 1 9 2 4 15 13 1 1 9 1 9 11 2
6 3 13 10 1 9 2
23 2 9 11 11 13 10 1 10 0 9 1 16 15 13 9 14 13 3 16 15 13 0 2
6 11 4 13 0 2 2
20 2 13 3 10 0 9 16 10 9 7 9 9 11 11 13 3 1 10 9 2
8 8 8 8 8 2 8 2 2
7 2 9 11 11 13 0 2
9 10 9 1 0 9 4 13 1 2
10 0 1 9 2 15 10 0 13 2 2
6 2 13 15 0 0 2
9 9 1 10 0 9 0 9 2 2
6 2 13 11 11 11 2
11 10 0 9 2 10 0 7 0 9 2 5
11 2 4 4 13 16 9 11 11 13 0 2
16 10 1 10 0 7 0 0 9 15 4 13 9 1 14 13 2
4 0 0 2 2
8 2 8 8 8 8 8 8 2
6 8 8 8 8 8 2
11 8 8 8 8 2 8 8 8 8 2 2
18 2 0 1 10 10 13 15 9 1 11 0 9 7 10 0 1 11 2
8 13 1 9 2 11 11 2 2
5 9 13 1 9 5
3 0 9 5
3 0 0 5
8 0 7 0 0 2 13 9 2
18 1 9 4 15 13 1 12 9 1 9 15 13 9 1 14 13 9 2
5 9 2 11 11 5
26 15 4 13 1 1 12 9 1 9 15 13 9 1 14 13 9 1 9 2 13 9 11 4 13 1 2
25 2 15 13 0 9 3 1 15 13 1 1 0 9 1 14 4 13 9 7 3 3 13 0 9 2
25 15 13 0 2 0 7 1 0 9 0 7 0 0 2 13 9 1 11 2 11 11 2 1 9 2
11 0 9 13 1 10 0 9 1 12 9 2
17 10 9 15 4 13 2 13 9 2 16 9 1 9 13 0 9 2
23 9 13 10 0 11 13 15 3 13 9 2 13 1 16 15 13 9 1 14 13 0 9 2
36 1 11 13 15 3 15 15 4 13 1 14 4 13 1 0 9 2 3 4 15 3 13 10 0 9 7 13 9 15 3 13 9 1 14 13 2
20 0 1 15 15 3 13 9 2 13 3 3 0 7 1 0 9 2 13 9 2
6 2 15 13 0 0 2
25 15 14 13 9 13 10 1 10 0 9 1 9 7 1 10 10 7 1 10 1 9 2 13 11 2
25 15 13 3 10 9 16 15 15 4 13 1 14 13 9 1 9 2 0 13 0 1 1 9 3 2
4 2 11 2 5
7 3 4 15 13 0 9 5
4 0 1 9 5
5 13 15 1 9 2
4 3 3 11 5
6 9 1 9 13 3 2
18 9 1 0 9 1 11 1 11 13 0 1 15 7 10 9 1 10 2
19 4 15 13 3 1 9 2 13 10 0 9 1 3 14 13 9 1 9 2
5 9 2 11 11 5
13 0 9 13 15 13 10 1 10 0 0 15 13 2
35 3 13 3 10 0 9 9 1 11 16 15 4 13 3 0 15 13 2 13 7 13 2 1 1 1 16 10 0 9 0 1 13 12 9 2
14 9 13 1 0 9 2 7 1 3 0 13 15 0 2
19 10 0 9 1 9 15 4 13 9 2 13 2 0 9 1 0 9 2 2
15 1 9 13 15 3 12 9 9 1 9 7 9 1 11 2
11 15 13 3 12 9 3 0 1 1 11 2
19 9 15 13 0 9 1 12 2 4 15 13 1 10 9 2 13 1 0 2
16 0 9 7 0 1 10 0 9 2 1 9 2 13 15 3 2
15 9 15 13 1 9 13 1 16 15 3 4 13 0 9 2
8 3 4 15 4 13 9 3 2
28 16 15 4 13 1 14 13 0 16 7 15 7 9 13 0 1 3 1 2 13 15 1 0 14 13 0 9 2
13 1 10 0 13 15 0 14 13 1 1 9 0 2
29 13 15 15 1 9 0 1 9 2 13 15 3 14 13 15 1 2 3 15 0 13 9 13 1 9 3 1 9 2
11 9 0 13 3 10 9 2 1 0 9 2
19 15 13 3 0 9 16 15 13 10 11 12 7 10 11 11 0 0 9 2
15 16 15 13 10 9 1 0 9 1 11 13 0 0 0 2
13 10 9 13 15 1 9 11 8 11 2 1 11 2
17 1 0 9 13 15 9 2 16 15 1 9 0 13 3 0 1 2
34 1 9 13 2 3 2 16 10 0 9 13 0 1 15 15 1 0 9 13 9 2 7 16 15 3 3 13 10 9 1 10 0 9 2
16 1 9 13 10 9 10 7 0 7 0 9 11 8 11 11 2
10 13 15 10 9 1 14 13 1 11 2
14 4 0 9 0 13 9 2 7 4 15 3 13 9 2
3 13 9 2
11 13 1 12 9 2 13 3 1 1 9 5
2 0 5
3 10 9 5
3 0 9 5
3 0 9 5
13 3 10 9 13 0 9 16 12 0 13 14 13 2
8 10 1 15 13 1 1 9 2
3 0 9 2
29 9 15 13 0 9 1 12 9 12 9 13 3 10 0 9 1 9 2 7 13 3 0 1 9 1 12 9 9 2
4 9 2 11 5
13 2 15 13 0 0 1 16 15 13 1 1 9 2
20 15 13 10 9 1 16 9 13 0 1 14 13 1 1 9 2 13 11 11 2
28 3 1 11 11 11 4 15 13 10 9 1 8 11 11 2 11 1 9 1 11 0 9 2 11 2 1 11 2
16 1 9 4 15 13 12 0 9 1 14 13 1 12 0 9 2
8 5 10 9 13 9 1 9 2
10 5 10 9 13 12 9 1 12 9 2
13 9 13 1 9 7 13 12 9 9 1 10 9 2
21 10 9 13 1 1 12 2 12 9 7 13 10 9 1 14 13 1 9 1 9 2
11 1 3 13 10 9 1 12 2 12 9 2
19 5 10 0 9 2 15 13 1 9 2 13 12 9 1 12 9 1 9 2
11 15 13 3 10 0 0 9 0 1 9 2
17 10 12 9 15 13 1 1 9 13 12 9 1 9 1 12 9 2
12 1 9 13 15 10 9 2 9 2 1 12 2
18 2 15 13 1 15 1 11 10 9 1 14 13 1 9 2 13 11 2
18 9 1 10 9 13 14 13 3 0 9 2 9 3 2 13 1 9 2
19 0 3 13 15 3 15 15 13 9 15 13 13 0 9 1 12 9 9 2
11 15 13 1 9 10 9 1 12 1 9 2
10 1 12 9 4 15 13 1 12 9 2
10 3 13 9 10 9 1 12 1 9 2
16 9 15 13 0 9 1 12 9 13 3 10 0 9 1 9 2
15 2 15 13 15 3 16 15 13 0 9 1 14 13 9 2
12 9 4 13 1 1 10 0 9 16 15 13 2
12 15 13 15 0 3 1 10 9 2 13 11 2
12 15 13 3 1 3 9 13 16 9 13 1 2
27 2 15 13 16 9 4 13 1 3 0 9 9 13 14 13 2 7 13 3 15 1 9 3 2 13 11 2
7 9 13 7 9 7 9 2
17 15 13 10 9 1 12 9 7 4 13 7 13 1 7 1 9 2
14 1 9 1 10 12 9 4 15 13 7 13 1 0 2
14 3 13 15 15 16 3 10 1 15 13 1 1 9 2
9 2 1 15 13 15 3 0 0 2
31 0 13 15 4 13 1 0 1 9 1 14 3 13 2 7 15 13 0 9 15 13 16 9 13 0 1 9 2 13 11 2
21 2 15 4 3 3 13 16 9 13 14 13 0 16 15 13 14 13 2 13 11 2
12 7 15 13 16 9 13 0 16 15 13 9 2
12 2 15 13 0 9 1 14 13 1 0 9 2
14 9 13 0 1 9 2 15 13 0 9 10 0 9 2
14 14 13 1 0 9 13 0 1 10 9 2 13 11 2
17 15 4 3 13 16 9 1 9 13 15 1 9 1 10 12 9 2
22 2 15 13 10 9 1 16 15 4 13 2 3 16 15 4 13 0 9 7 0 9 2
17 15 13 16 9 0 13 15 16 9 13 15 1 9 2 13 11 2
10 9 13 3 16 9 13 0 1 9 2
25 2 15 13 3 16 0 9 13 0 2 16 15 13 0 14 13 1 9 7 10 9 2 13 11 2
18 1 1 1 16 9 3 13 2 3 13 15 0 1 9 1 12 9 2
12 9 4 13 1 16 15 13 3 0 15 13 2
18 3 13 15 15 15 4 13 9 1 9 15 13 0 9 1 9 10 2
10 15 13 3 12 9 0 1 1 9 2
12 10 10 13 3 9 0 2 7 3 3 0 2
6 0 14 13 9 3 5
3 13 3 5
5 2 3 13 3 5
4 13 14 13 5
5 4 13 1 9 5
6 0 9 1 12 9 5
6 2 9 1 9 0 5
22 9 1 11 4 13 12 9 2 7 13 1 14 13 0 0 2 13 11 9 11 11 2
9 1 11 13 11 11 1 0 9 2
21 10 9 1 11 13 1 12 9 7 13 9 1 12 9 2 1 9 11 11 11 2
6 9 2 11 11 11 5
20 10 0 12 9 4 11 11 2 12 2 13 9 1 10 0 9 11 1 9 2
13 2 15 13 1 1 9 1 9 1 10 10 9 2
18 9 13 14 13 10 0 0 0 1 10 9 7 3 13 15 1 3 2
8 3 4 15 13 0 0 9 2
23 3 3 1 11 13 9 0 1 9 15 9 3 0 13 9 1 14 13 1 2 13 15 2
17 1 11 13 12 12 0 9 9 1 14 13 9 1 9 1 9 2
9 12 9 13 1 14 13 1 9 2
7 13 10 0 9 1 11 2
23 11 11 2 12 2 1 11 4 13 9 1 11 1 12 7 4 13 0 1 11 1 12 2
15 7 15 7 11 13 9 4 13 14 13 1 0 9 1 2
10 2 15 13 3 14 13 1 1 9 2
14 0 9 13 1 9 1 14 13 1 15 9 15 13 2
9 11 13 3 1 9 2 13 11 2
38 1 9 1 9 13 15 7 9 1 1 10 3 0 9 15 15 4 13 0 7 0 3 15 15 13 2 1 9 2 9 7 0 9 1 9 1 9 2
12 9 13 12 9 7 13 0 1 1 12 9 2
10 2 15 13 15 14 13 3 1 11 2
15 15 13 3 0 9 1 16 15 13 0 15 2 13 15 2
31 9 1 10 0 9 4 13 12 2 12 9 1 9 1 12 2 7 13 1 14 13 0 0 2 13 11 9 2 11 11 2
25 1 10 9 15 13 1 10 9 2 13 11 7 10 9 16 11 4 13 0 16 15 0 4 13 2
10 2 9 13 14 13 2 7 9 13 2
12 7 9 1 11 4 13 1 1 0 9 3 2
19 15 13 1 14 13 10 9 16 9 1 11 13 14 13 15 2 13 11 2
10 2 7 3 4 9 13 13 3 0 2
15 2 6 2 15 13 1 12 2 12 9 1 2 13 15 2
28 3 4 15 13 0 1 0 9 2 7 15 13 3 0 1 1 9 16 15 13 10 0 9 3 2 13 11 2
11 4 15 13 9 1 9 1 9 7 9 2
9 7 4 15 4 13 1 0 9 2
7 13 15 9 1 10 9 2
18 0 9 4 13 0 9 9 7 9 1 16 9 4 13 7 9 13 2
14 0 9 4 13 1 9 1 16 9 4 13 1 9 2
9 2 3 13 15 9 4 13 0 2
32 2 1 1 1 9 13 15 2 1 9 15 4 13 2 3 16 16 15 13 9 1 10 9 2 13 15 3 0 14 13 9 2
7 15 4 3 13 10 9 2
16 13 15 1 10 9 7 9 2 13 15 3 0 14 13 9 2
21 3 4 3 9 3 13 14 13 16 15 4 13 9 1 1 10 0 13 4 13 2
22 10 0 9 13 14 13 2 7 15 13 3 1 14 13 0 2 0 9 2 13 11 2
16 11 9 4 1 9 1 15 13 9 1 11 1 12 7 12 2
22 2 1 9 1 10 0 9 13 15 16 11 4 13 1 9 1 9 7 11 0 9 2
15 11 4 3 13 1 1 9 1 9 2 13 11 1 9 2
26 0 9 13 3 12 9 9 1 0 9 7 9 1 9 1 9 1 9 9 1 12 2 1 11 11 2
20 10 0 12 9 4 13 1 9 9 1 10 9 1 14 13 0 9 1 9 2
40 9 11 4 2 1 1 1 9 1 1 1 12 9 2 3 13 14 13 9 1 9 1 10 9 1 11 8 11 2 3 0 1 11 2 13 9 11 1 9 2
21 9 13 9 1 0 1 12 9 1 9 2 1 9 1 10 9 1 9 1 9 2
30 2 3 2 1 15 1 9 2 4 9 13 0 13 1 9 9 13 2 13 11 11 2 0 1 9 9 2 1 11 2
23 0 11 11 15 13 1 11 13 9 1 14 13 13 15 2 3 16 15 3 13 15 0 2
11 2 15 13 0 0 9 9 2 13 11 2
20 0 11 11 11 1 11 11 11 4 13 9 1 9 1 12 7 13 9 0 2
18 15 13 16 9 1 9 1 9 4 13 1 12 9 1 9 1 12 2
20 2 15 13 10 9 1 16 0 9 13 9 1 9 1 11 3 1 1 9 2
13 10 0 9 13 3 3 10 0 9 2 13 15 2
27 1 9 9 4 15 13 12 9 1 10 9 2 7 9 4 1 9 1 10 0 9 13 0 1 1 12 2
10 1 12 9 3 13 15 1 9 12 2
39 2 15 13 0 14 13 3 9 7 9 4 13 15 0 2 15 13 3 1 9 1 11 2 7 15 13 10 9 1 16 15 13 9 9 3 2 13 11 2
21 1 9 13 15 1 10 10 12 9 0 9 1 11 11 1 11 11 3 1 11 2
23 9 15 1 12 13 1 12 12 9 2 13 3 9 1 12 12 9 7 1 12 12 9 2
12 2 15 13 0 1 9 1 9 3 4 13 2
16 10 9 13 15 1 9 0 1 1 9 7 1 10 0 9 2
23 1 10 9 13 15 0 1 10 0 2 0 9 15 15 13 10 9 1 11 2 13 11 2
6 9 13 0 0 9 5
6 9 1 11 0 9 5
3 2 9 5
26 9 11 10 13 0 1 14 13 10 0 9 2 15 4 13 1 9 1 0 9 1 9 9 7 9 2
10 15 13 9 11 11 2 9 1 9 2
30 11 11 4 9 13 1 9 1 12 9 1 14 4 4 13 0 1 14 4 13 1 12 0 9 15 9 4 4 13 2
27 16 11 3 13 10 10 9 2 13 11 1 14 13 15 15 0 13 1 9 1 9 1 9 10 1 11 2
29 9 4 13 1 9 1 9 2 7 13 0 1 14 4 13 9 1 9 9 2 13 15 7 13 9 0 1 9 2
9 9 4 13 1 9 2 11 2 2
26 16 9 13 2 13 11 16 15 3 13 10 9 2 7 4 13 9 1 2 9 1 9 7 9 2 2
11 9 13 0 1 9 9 1 12 9 9 2
16 9 13 3 3 9 1 11 9 2 15 13 9 1 10 9 2
17 9 13 3 0 16 15 13 1 16 11 13 0 2 7 13 3 2
22 1 9 4 11 4 13 16 15 13 1 15 10 1 2 10 9 1 11 0 9 2 2
22 15 4 13 9 7 13 15 0 0 16 11 13 0 1 9 7 9 1 9 1 11 2
17 1 10 9 1 1 11 13 9 12 9 15 4 13 1 9 0 2
26 10 9 1 12 9 2 3 12 9 2 2 10 9 7 10 0 9 1 10 0 9 11 2 11 2 2
11 11 13 15 3 2 13 9 1 2 9 2
22 15 4 13 10 0 9 16 15 13 1 9 1 9 2 15 4 13 0 0 1 9 2
29 2 15 4 13 1 10 9 9 13 15 13 0 2 15 15 13 0 1 7 13 9 1 2 13 10 9 1 11 2
27 0 9 4 13 1 16 15 4 13 10 0 9 1 9 1 9 9 2 1 16 15 4 13 14 13 15 2
16 9 1 11 13 3 0 1 11 7 13 0 0 1 9 11 2
31 9 13 10 0 9 1 0 9 2 15 13 10 9 9 2 9 2 7 13 1 9 1 11 9 2 15 13 0 10 9 2
9 11 4 3 13 1 14 13 9 2
5 0 9 1 9 5
10 13 1 12 7 10 0 9 3 0 5
6 13 3 1 12 9 5
4 13 15 1 5
5 2 13 3 0 5
9 1 13 9 0 1 9 7 9 2
5 1 13 9 0 2
22 2 15 4 13 9 7 13 15 13 15 15 3 13 14 13 3 2 13 10 0 9 2
20 15 4 13 15 1 1 9 1 11 11 1 14 13 15 10 9 1 10 9 2
12 7 15 13 3 0 1 2 7 13 3 9 2
8 2 3 3 13 15 0 3 2
19 7 15 13 3 16 15 13 9 1 10 9 7 9 1 12 2 13 15 2
9 0 0 4 13 1 15 9 9 2
27 0 1 9 13 9 0 1 0 2 7 15 13 0 0 14 13 15 1 15 15 13 3 1 14 13 9 2
21 10 3 0 13 15 1 3 9 12 2 12 7 10 0 9 16 9 1 9 13 2
33 2 15 13 15 4 13 3 0 9 2 7 15 13 16 15 4 13 0 1 2 13 11 11 2 12 2 7 11 11 2 12 2 2
11 10 12 4 13 15 9 1 9 12 1 2
20 1 9 12 13 15 14 13 1 1 9 15 4 13 15 3 0 9 1 9 2
18 2 15 4 13 3 3 0 2 7 15 4 13 15 0 2 13 11 2
12 15 13 1 9 1 9 7 9 11 11 11 2
22 15 13 9 1 12 9 0 1 9 2 7 13 15 13 9 14 13 9 0 1 9 2
7 2 15 4 13 0 9 2
15 15 13 0 1 0 9 7 9 9 1 9 2 13 15 2
10 2 7 10 9 13 15 3 1 9 2
18 2 3 13 9 1 12 7 12 9 2 7 9 13 0 2 13 9 2
6 2 13 15 0 15 2
13 2 6 2 16 15 13 1 1 9 3 2 3 2
4 15 13 0 2
11 0 9 12 13 15 15 1 1 10 9 2
27 2 6 15 3 2 3 13 9 2 13 15 3 0 15 13 2 7 13 14 13 1 9 1 10 0 9 2
17 15 1 15 13 9 15 1 1 14 13 15 9 15 4 13 1 2
16 2 13 14 13 9 2 9 2 9 7 9 1 2 13 9 2
11 1 9 4 9 10 13 1 11 11 11 2
9 9 9 12 13 1 1 9 10 2
12 2 15 13 3 0 3 10 9 2 13 15 2
7 2 7 9 4 15 13 2
17 2 16 15 3 4 13 3 3 0 4 15 3 13 15 10 9 2
6 10 0 9 1 12 5
5 2 4 13 9 5
4 9 13 0 5
4 11 0 9 5
3 11 9 5
3 11 9 5
5 11 9 1 9 5
4 9 1 11 5
7 11 11 0 9 1 9 5
5 9 1 11 9 5
3 11 9 5
3 11 9 5
4 9 1 11 5
10 0 9 4 13 15 1 9 15 13 2
14 10 9 7 9 13 3 16 12 9 4 13 1 9 2
24 1 9 1 9 1 11 11 2 11 11 11 2 3 4 15 13 15 1 16 9 13 0 9 2
25 2 1 9 4 9 3 13 9 1 10 9 2 3 4 9 13 1 7 15 13 1 1 0 9 2
14 15 13 3 16 9 4 13 9 1 9 2 13 15 2
34 15 13 12 9 9 4 13 9 1 2 7 1 16 15 13 10 0 15 13 16 15 3 13 9 1 9 7 1 16 9 13 10 0 2
19 2 16 9 13 15 1 3 13 15 0 7 0 1 16 9 13 10 0 2
13 9 13 1 9 9 7 15 9 13 2 13 11 2
11 1 9 2 13 15 10 0 9 1 9 2
15 10 0 10 9 4 13 13 16 9 1 9 13 15 0 2
7 2 9 13 10 0 9 2
12 15 13 1 9 3 0 1 16 15 13 9 2
8 9 4 1 9 13 0 9 2
11 7 13 15 2 3 4 15 13 10 9 2
10 15 4 13 9 1 9 2 13 15 2
20 9 4 3 3 13 1 9 2 7 3 1 9 7 15 4 0 13 0 0 2
20 2 10 9 13 9 1 14 13 9 1 14 13 16 15 3 4 13 1 9 2
10 9 1 14 13 10 9 4 13 0 2
14 3 13 12 9 1 9 15 4 13 15 1 1 12 2
27 7 0 9 2 0 9 7 0 9 13 11 9 1 9 10 2 15 13 1 16 9 9 1 3 4 13 2
7 1 12 9 9 4 13 2
13 15 4 13 15 14 13 10 0 9 1 9 3 2
10 15 13 3 12 9 16 11 13 9 2
20 11 9 13 16 10 9 1 9 13 1 10 0 2 9 2 1 10 0 9 2
11 0 9 1 9 13 1 10 9 1 11 2
11 16 9 13 9 13 15 9 1 9 3 2
10 7 9 13 3 9 1 9 1 9 2
29 2 15 13 0 9 11 4 13 10 10 0 9 2 7 3 13 15 9 3 4 13 1 15 1 10 9 1 9 2
23 7 1 9 13 15 0 16 15 13 15 10 9 15 4 13 16 9 13 9 1 9 3 2
16 3 4 15 0 13 10 0 0 9 1 9 1 2 13 11 2
14 0 9 13 11 10 0 9 1 9 1 9 1 9 2
11 11 13 1 10 9 3 3 0 1 9 2
16 3 1 9 1 9 13 11 11 9 1 14 13 9 1 9 2
16 11 13 3 11 7 9 1 14 13 9 1 9 1 9 12 2
24 15 13 9 10 1 9 10 9 2 7 9 13 3 16 15 13 11 4 13 9 3 1 9 2
18 11 9 13 16 15 13 14 13 1 10 9 15 4 13 1 0 9 2
37 15 13 0 10 9 15 4 13 9 1 10 9 2 7 13 1 16 10 9 13 9 1 9 7 10 9 1 10 2 0 2 0 9 1 0 9 2
17 9 13 1 16 0 4 13 9 1 11 9 1 0 9 7 9 2
17 9 7 9 4 13 1 9 1 16 9 4 13 1 9 1 9 2
9 2 3 13 15 14 13 10 9 2
12 3 13 15 9 1 9 11 11 7 3 15 2
9 15 13 10 9 15 13 10 9 2
14 16 15 13 0 9 3 4 15 13 1 9 1 9 2
19 7 15 4 3 13 1 16 9 13 10 0 0 9 1 9 2 13 11 2
11 11 13 14 4 13 0 1 10 9 10 2
24 0 1 9 15 9 13 2 4 3 3 13 13 3 16 15 4 13 1 1 12 9 1 9 2
19 0 15 13 1 9 15 0 4 13 1 9 11 13 0 9 13 1 9 2
16 1 11 2 13 15 0 12 0 15 13 13 0 12 9 9 2
9 0 0 13 9 1 1 12 9 2
15 9 13 1 16 11 13 9 1 11 9 1 9 1 9 2
15 2 1 11 4 13 10 9 15 13 1 10 0 0 9 2
22 16 15 13 1 9 1 9 9 3 4 15 13 16 15 13 9 7 9 2 13 11 2
23 15 13 1 9 0 16 11 2 1 12 9 1 11 2 13 1 9 15 13 9 1 9 2
22 15 13 9 1 11 11 1 14 13 1 15 15 13 13 10 2 0 9 2 1 9 2
17 1 12 9 9 1 13 15 1 9 7 13 9 1 14 13 9 2
20 11 13 3 9 1 14 13 1 16 15 3 13 10 0 9 1 9 1 9 2
14 7 12 9 1 16 15 4 13 9 2 3 13 9 2
8 2 15 13 0 1 9 9 2
12 9 1 9 1 11 13 16 9 4 13 0 2
8 3 13 15 10 9 15 13 2
8 9 1 9 13 3 0 3 2
19 7 15 4 3 3 13 1 10 9 16 0 0 9 13 9 2 13 11 2
8 9 11 11 13 9 1 9 2
9 11 4 1 9 13 9 1 9 2
21 15 13 1 10 1 14 4 13 9 9 1 14 13 1 10 9 1 11 1 11 2
31 15 13 1 9 1 9 16 9 13 10 9 7 12 10 9 7 13 15 1 9 1 9 1 11 2 15 13 11 0 9 2
15 1 9 4 0 12 9 13 2 1 10 0 9 11 11 2
27 0 0 1 9 4 1 10 13 1 14 4 13 1 9 1 1 3 1 12 9 9 1 10 0 9 11 2
16 1 9 1 9 3 4 11 13 1 9 1 9 1 11 1 2
17 2 3 13 15 3 3 10 9 2 7 10 9 15 13 10 9 2
12 15 13 1 16 15 4 13 9 1 10 9 2
18 15 13 0 16 9 13 16 15 0 13 9 1 10 9 2 13 11 2
14 11 11 13 10 0 9 11 7 11 1 9 1 9 2
12 15 4 13 0 9 1 9 1 10 0 9 2
13 9 13 14 4 13 1 12 9 9 1 0 9 2
23 1 11 4 15 13 15 1 9 2 16 9 1 10 0 9 4 13 3 0 1 0 9 2
15 0 9 11 11 1 11 7 11 13 1 1 9 1 9 2
18 11 13 0 1 11 16 15 13 16 9 1 9 13 1 9 1 9 2
11 9 13 1 9 1 11 2 0 11 2 2
20 1 12 4 11 11 0 13 1 14 4 13 1 9 1 10 9 0 1 11 2
23 2 9 15 13 3 1 13 16 9 3 4 13 1 1 3 15 13 14 13 10 0 9 2
24 15 4 13 9 7 3 13 15 10 9 2 7 0 4 15 3 13 15 0 3 2 13 11 2
26 9 0 1 12 1 12 9 15 4 13 14 13 1 12 9 2 4 13 1 9 1 12 1 12 9 2
10 9 13 0 7 0 1 3 0 9 2
20 1 9 13 15 0 16 11 9 13 1 9 1 15 10 1 12 9 1 9 2
17 11 11 13 7 13 9 7 9 2 15 13 1 1 9 1 11 2
5 9 13 12 0 2
12 9 1 9 13 1 9 1 1 12 9 9 2
16 9 13 3 16 9 4 13 0 12 9 9 1 9 1 12 2
16 1 10 0 9 1 9 1 11 9 13 15 1 10 1 9 2
13 2 15 13 10 0 0 9 1 9 1 11 2 2
24 9 11 11 2 11 2 13 16 15 13 0 1 1 15 15 13 1 2 9 1 9 9 2 2
14 15 13 16 15 13 0 14 13 1 3 9 13 3 2
17 1 16 3 15 13 3 3 4 11 3 13 1 10 0 0 9 2
11 1 10 4 9 13 1 14 13 9 10 2
14 2 15 13 9 1 0 9 7 10 0 9 1 9 2
15 15 4 13 9 9 1 14 13 15 0 9 2 13 11 2
26 10 0 9 1 9 11 13 1 9 1 16 15 13 1 7 1 1 9 0 9 1 11 11 1 9 2
16 1 9 1 9 13 9 13 16 9 13 1 1 10 0 9 2
15 3 1 13 0 1 9 9 1 9 1 10 0 0 9 2
35 0 13 3 9 9 16 11 7 11 9 13 9 1 10 0 9 1 11 11 11 2 15 15 13 1 9 1 12 9 1 11 9 7 9 2
15 2 15 13 15 13 0 9 15 4 13 1 10 10 9 2
19 15 13 1 0 9 2 7 4 13 0 0 9 7 4 13 1 0 9 2
6 15 13 10 0 9 2
5 9 13 10 9 2
7 3 4 11 9 13 1 2
10 15 4 13 15 0 3 2 13 11 2
28 1 9 1 9 12 13 9 1 9 1 10 0 9 11 11 14 13 0 2 1 0 9 0 9 9 1 9 2
30 16 11 11 11 11 4 13 0 0 9 13 15 10 9 15 13 1 15 12 9 1 9 2 9 7 10 9 1 9 2
19 1 9 4 11 13 0 0 2 7 9 1 9 13 1 1 12 9 9 2
14 1 9 4 11 13 7 13 1 0 0 9 7 9 2
11 2 1 9 13 15 9 1 10 9 9 2
10 1 9 13 15 3 9 15 13 3 2
9 11 13 3 1 15 2 13 11 2
20 1 9 12 4 11 13 1 9 1 9 1 9 1 9 0 1 2 9 2 2
23 9 12 13 15 0 1 11 16 11 3 13 1 9 11 9 1 14 13 9 1 10 9 2
9 11 13 3 14 13 9 1 9 2
12 11 13 14 13 10 3 0 9 1 10 9 5
18 10 9 4 13 1 10 9 0 1 16 15 13 10 10 9 1 9 2
8 2 1 9 4 15 13 0 2
11 15 13 10 0 9 14 13 15 1 11 2
8 3 4 11 13 10 0 9 2
12 15 13 3 3 15 4 13 1 10 10 9 2
10 15 13 0 1 10 9 2 13 11 2
7 2 11 4 13 10 9 5
2 9 5
3 0 9 5
5 9 1 12 9 5
6 2 9 13 3 0 5
15 9 1 12 2 12 9 9 13 1 9 1 10 0 9 2
8 9 13 0 1 11 1 11 2
15 0 1 9 0 4 13 9 7 9 1 9 1 10 9 2
2 9 2
8 9 2 11 11 11 5 11 5
22 16 15 13 10 12 2 12 9 1 9 4 10 0 9 3 1 11 1 11 13 10 2
2 9 2
8 9 2 11 11 11 5 11 5
20 9 11 11 1 11 11 13 15 13 0 14 13 1 0 11 1 11 1 11 2
11 2 11 13 0 0 1 1 10 9 9 2
11 15 13 0 9 1 11 2 11 7 11 2
22 15 13 10 9 0 9 1 15 15 13 1 11 2 13 11 11 1 11 11 1 11 2
19 15 13 3 1 16 15 13 10 9 1 2 0 2 7 2 0 2 9 2
16 10 0 13 3 10 0 9 1 11 7 11 2 16 11 13 2
10 9 1 0 0 9 13 0 1 9 2
16 10 0 9 1 11 13 16 12 9 9 13 10 9 0 13 2
7 4 13 0 9 1 9 5
12 2 15 13 3 9 1 10 9 9 1 11 2
13 9 13 16 9 13 9 7 0 9 2 13 11 2
10 15 13 16 11 4 13 0 0 1 2
7 2 11 4 13 10 9 2
12 15 13 3 0 1 9 2 13 15 1 11 2
17 11 13 3 16 15 13 0 9 1 9 1 9 1 9 1 9 2
20 15 4 3 13 10 0 0 9 2 7 4 13 9 1 9 1 9 7 9 2
22 2 15 13 15 15 13 0 9 2 13 11 7 13 1 10 9 1 12 9 1 11 2
14 10 9 16 15 4 13 1 11 4 15 13 0 0 2
33 3 16 15 13 0 9 1 9 1 9 2 13 3 9 1 9 2 11 11 11 2 16 9 4 13 1 10 0 0 9 1 11 2
12 15 13 3 9 15 13 16 11 13 1 9 2
17 13 15 16 15 13 9 1 11 2 3 13 15 3 13 10 0 2
26 15 13 3 16 15 13 0 9 7 16 9 4 13 9 1 0 9 2 11 13 10 0 9 1 15 2
7 10 0 9 13 9 3 2
17 13 15 16 15 13 9 1 11 2 3 13 15 3 13 10 0 2
6 15 13 3 10 9 2
21 15 13 3 16 15 13 0 9 7 16 9 4 13 9 1 0 9 2 13 11 2
13 2 15 13 0 1 16 0 7 0 13 1 9 2
9 7 1 11 13 9 2 13 11 2
17 1 9 1 9 1 9 13 15 0 12 9 1 9 0 1 11 2
15 9 13 1 3 1 12 9 9 2 7 12 9 1 9 2
21 3 1 9 13 3 12 9 1 11 9 1 9 2 1 10 9 1 12 9 9 2
20 1 12 9 3 13 11 16 15 1 9 1 9 13 9 1 9 1 10 9 2
14 0 13 15 12 9 1 9 1 12 9 9 1 9 2
17 2 10 9 9 4 13 16 9 3 13 3 0 0 15 15 13 2
9 3 13 15 3 1 10 0 9 2
13 0 9 13 16 15 13 2 7 15 13 0 0 2
11 10 9 1 9 13 0 0 1 9 9 2
17 13 15 9 1 9 2 3 13 15 3 9 2 13 11 11 11 2
14 10 0 9 1 11 3 3 13 10 9 1 3 11 2
12 12 9 9 13 1 1 9 1 11 1 11 2
7 9 13 1 12 9 9 2
13 3 13 15 0 1 9 2 7 15 13 0 9 2
16 2 15 13 9 1 12 9 9 1 9 2 7 15 13 3 2
13 1 10 9 3 3 2 13 9 11 11 1 11 2
16 1 10 0 9 1 11 13 15 0 1 0 9 1 0 9 2
9 2 15 13 10 10 9 1 11 2
8 12 2 12 9 13 1 9 2
20 15 13 0 9 2 7 15 13 0 1 9 2 13 9 11 11 1 11 12 2
13 0 1 11 7 11 13 15 0 0 9 1 9 2
13 1 11 13 15 12 9 1 9 2 1 11 12 2
15 0 1 15 13 0 9 2 3 16 10 0 9 13 0 2
26 1 11 13 15 9 7 9 1 10 1 11 2 11 2 11 2 11 2 11 2 11 2 11 7 11 2
19 1 11 13 9 1 12 9 7 0 9 1 12 9 1 11 3 1 9 2
10 2 15 13 1 15 9 13 0 0 2
5 15 13 3 0 2
23 3 16 9 13 0 15 2 4 15 3 13 3 16 15 3 13 3 0 9 2 13 11 2
16 15 13 16 9 1 10 9 9 3 13 0 1 9 10 9 2
4 9 11 11 5
4 9 1 9 5
3 9 9 5
4 1 1 9 5
4 10 10 9 5
4 0 7 0 5
17 11 11 13 10 9 15 7 4 13 1 7 13 2 13 11 11 2
3 9 9 2
8 11 11 13 1 11 0 9 2
7 9 2 11 11 2 11 5
9 11 11 13 0 1 9 1 11 2
20 15 13 3 10 11 11 2 11 11 7 11 11 15 13 9 1 11 0 9 2
21 7 16 15 13 0 9 7 3 0 9 2 4 0 9 9 2 11 11 2 13 2
14 11 11 11 13 1 1 10 1 12 9 1 10 9 2
10 1 9 13 15 0 1 10 0 9 2
25 3 1 9 13 15 10 0 9 2 9 2 11 2 2 15 15 13 3 1 9 7 9 1 9 2
18 16 15 13 10 0 9 3 1 11 11 2 13 15 10 9 1 15 2
21 12 9 7 1 12 9 0 9 0 2 13 11 7 9 11 1 9 0 0 9 2
47 1 1 1 16 15 1 0 9 4 13 9 7 9 3 2 13 11 1 14 13 10 0 0 9 7 9 1 11 9 2 10 0 0 2 0 7 0 9 15 9 0 13 3 4 13 1 2
5 3 13 15 1 2
20 9 9 4 13 1 11 1 12 1 11 2 11 11 2 11 11 7 11 11 2
23 15 13 12 9 1 1 9 1 10 0 9 2 15 9 9 13 10 9 1 2 11 11 2
9 15 13 1 9 2 9 7 9 2
2 3 2
25 1 10 0 9 1 10 0 9 2 13 9 1 10 0 9 2 10 9 2 15 15 13 1 9 2
31 10 9 2 3 0 2 11 9 2 2 4 4 13 1 3 0 7 0 16 15 13 0 1 9 7 1 1 9 1 9 2
38 1 9 1 9 9 4 9 13 9 1 9 1 11 2 11 11 11 11 2 7 11 11 2 11 11 11 8 11 2 2 1 9 7 9 1 0 9 2
18 3 13 9 1 10 0 9 1 10 0 7 0 2 1 3 0 9 2
18 11 13 3 1 1 15 7 0 13 15 1 10 9 7 9 1 9 2
23 9 1 2 11 11 2 13 1 1 16 9 11 4 13 10 9 1 10 0 9 11 11 2
15 15 13 1 15 10 9 7 13 9 13 1 9 1 9 2
9 1 10 9 1 13 11 0 1 2
28 2 8 8 2 2 13 15 2 7 15 13 1 1 16 15 13 1 1 9 1 9 1 9 0 7 0 9 2
9 10 9 4 13 2 9 13 9 2
12 16 11 13 10 9 2 13 15 3 1 9 2
23 15 13 3 9 1 9 9 1 9 7 9 2 7 15 13 0 10 0 9 1 10 0 2
25 0 9 2 0 9 7 9 13 10 9 1 9 2 16 9 4 13 1 10 9 1 10 0 9 2
17 15 1 11 2 11 2 1 9 1 11 11 13 9 1 10 0 2
25 11 11 2 11 11 2 11 11 7 1 7 1 11 11 13 1 10 9 1 0 9 1 0 9 2
34 0 1 9 2 11 7 11 2 1 10 0 9 11 11 2 16 10 11 13 1 11 2 13 11 11 2 11 11 8 11 2 1 12 2
27 0 13 10 0 9 1 9 9 1 9 1 10 0 9 15 13 9 9 2 1 1 9 11 9 1 12 2
41 16 10 9 13 0 1 0 9 2 0 9 7 9 1 9 2 13 11 11 10 0 9 1 10 0 7 0 9 2 1 0 9 1 0 9 1 9 1 10 0 2
15 11 11 13 3 9 9 2 7 4 13 0 1 9 9 2
14 13 1 10 0 9 1 11 11 7 0 11 1 9 2
9 15 4 3 13 10 9 1 9 2
15 3 1 9 2 4 9 0 13 1 10 9 7 10 9 2
25 16 10 0 9 11 11 13 11 9 2 11 8 11 2 1 12 2 4 9 3 13 1 10 9 2
28 16 10 0 7 0 9 0 13 1 1 9 0 1 9 2 9 7 9 1 9 2 4 9 3 13 9 9 2
33 9 9 4 1 3 0 13 1 10 10 9 15 13 1 10 9 2 10 9 1 14 13 1 10 10 9 7 13 15 10 10 9 2
17 9 13 15 3 0 0 0 2 7 1 10 0 0 7 0 9 2
19 9 13 2 1 10 10 9 2 1 1 9 15 13 15 1 3 7 3 2
22 16 10 9 13 10 9 1 9 2 13 10 9 0 1 1 9 2 1 9 7 9 2
10 10 4 13 1 9 1 10 0 9 2
21 15 13 0 7 13 1 1 9 2 16 9 7 0 13 1 1 9 1 0 9 2
26 9 4 3 13 3 1 9 2 7 13 1 1 15 15 3 13 3 2 1 9 2 7 15 13 0 2
50 9 9 13 3 1 9 2 1 16 9 2 0 9 7 0 9 13 15 2 16 15 13 9 2 9 7 9 1 0 0 0 9 2 9 2 9 2 11 11 11 2 16 0 9 13 1 9 1 9 2
23 9 13 10 9 2 16 3 10 0 9 13 0 2 1 10 9 15 13 0 7 0 0 2
23 16 10 0 0 9 4 13 0 1 9 2 9 7 0 9 2 3 13 9 10 0 9 2
17 1 9 2 11 2 11 11 8 11 2 2 13 11 11 1 9 2
15 10 9 13 0 1 11 11 2 15 13 10 0 1 9 2
16 10 9 4 13 14 13 1 9 10 2 1 10 9 0 9 2
21 15 13 3 10 9 1 10 9 2 3 3 1 9 2 7 3 1 0 10 9 2
16 15 13 10 0 0 2 7 0 9 15 13 0 9 1 9 2
14 10 9 1 15 13 10 9 11 1 2 10 9 2 2
6 15 13 1 1 15 2
21 15 13 10 0 7 0 1 9 10 2 15 13 10 9 1 10 0 7 0 9 2
10 10 1 9 1 11 11 9 13 3 2
27 10 0 7 0 9 13 1 9 1 9 2 16 11 13 10 0 7 0 9 15 13 10 9 1 0 9 2
11 3 4 15 13 16 11 9 13 11 11 2
25 15 13 16 15 4 13 10 9 9 1 14 13 3 0 1 9 9 15 13 1 1 9 1 9 2
9 7 11 7 11 13 1 9 3 2
15 7 3 0 9 4 13 10 9 13 1 0 9 11 11 2
37 16 15 1 12 13 10 9 1 2 11 11 11 2 7 13 15 1 0 9 7 0 9 2 13 15 0 3 1 10 0 9 2 1 10 0 9 2
18 1 9 4 11 1 0 0 9 13 1 10 9 1 1 10 0 9 2
38 1 9 1 9 13 15 0 1 7 1 1 9 1 10 0 9 2 7 13 3 0 1 9 16 9 1 10 13 0 1 10 0 9 1 10 0 9 2
35 15 13 10 0 1 9 15 13 16 15 13 3 0 1 9 2 15 15 13 1 9 1 10 9 15 0 4 13 0 1 9 1 10 0 2
17 15 13 3 0 11 9 11 11 2 15 3 13 1 9 1 9 2
20 1 9 1 10 9 1 9 2 13 15 16 9 4 13 10 0 9 1 11 2
21 15 4 13 1 10 0 9 2 11 11 2 2 15 3 13 9 9 1 0 9 2
27 1 10 9 4 15 3 13 1 15 7 13 15 0 2 7 1 0 4 9 3 13 10 2 0 9 2 2
29 11 13 0 9 1 9 1 9 2 7 15 13 1 9 2 11 11 2 1 12 16 15 1 9 13 10 0 9 2
24 1 9 13 15 10 9 15 13 9 9 2 16 9 2 9 7 9 13 1 1 10 0 9 2
30 10 2 9 9 2 2 0 1 9 1 10 0 9 7 9 2 0 0 1 0 9 1 11 11 1 0 9 1 15 2
12 1 9 4 15 13 2 13 7 13 1 15 2
6 11 13 9 11 11 2
4 9 1 9 5
4 9 1 9 5
3 0 9 5
5 0 2 1 9 5
2 9 5
3 0 9 5
2 9 5
4 13 1 9 5
24 4 10 0 0 9 0 13 3 0 16 15 13 14 13 1 9 0 16 10 1 15 0 13 2
24 1 9 13 15 9 0 1 9 0 1 9 2 7 1 10 0 9 4 15 13 1 1 9 2
27 15 4 13 9 1 0 9 1 11 7 11 2 0 1 16 15 3 13 0 1 12 9 14 13 15 1 2
7 9 7 9 13 0 0 2
32 16 15 10 13 9 7 4 13 10 9 1 10 0 0 9 2 13 15 0 1 10 9 1 3 0 15 13 14 13 0 9 2
19 3 13 15 15 1 14 13 10 10 9 2 3 1 14 13 3 15 13 2
38 15 13 3 0 14 13 9 2 7 15 13 15 1 10 9 15 13 15 0 0 14 13 1 16 15 4 13 1 0 9 7 13 14 13 10 0 9 2
6 10 9 1 15 13 2
10 2 15 13 15 13 3 11 3 13 2
33 15 13 10 9 2 7 3 9 13 16 15 4 13 0 14 13 1 0 9 2 3 16 15 3 13 10 9 1 10 0 9 2 2
9 15 13 1 14 13 9 1 9 2
2 0 2
16 10 10 9 4 15 13 1 14 13 15 15 13 0 0 0 2
15 15 4 3 3 13 10 9 1 14 13 15 10 1 9 2
18 15 13 0 3 14 13 15 3 1 9 7 13 14 13 1 1 9 2
30 0 9 13 1 1 14 13 9 1 11 1 9 2 7 3 13 15 15 15 3 13 10 9 1 9 15 13 1 9 2
24 9 13 1 3 9 3 10 0 15 4 13 1 7 1 16 15 3 4 13 9 15 13 1 2
23 16 9 1 10 9 13 1 9 13 15 0 9 15 13 1 14 13 9 1 9 7 9 2
15 9 1 10 9 3 13 1 9 2 7 13 1 0 9 2
20 2 15 13 3 10 9 1 14 4 13 10 10 0 0 9 1 1 9 2 2
23 15 4 13 16 9 13 9 0 2 7 10 9 13 15 3 1 16 0 9 13 0 9 2
35 15 4 3 13 1 10 9 15 10 4 13 13 1 2 9 2 9 7 9 2 2 7 15 4 1 9 13 10 0 9 1 1 0 9 2
39 0 13 15 15 15 13 1 10 9 3 1 9 13 0 1 2 1 9 1 9 7 9 0 1 9 2 7 9 13 16 9 1 10 9 0 4 13 9 2
23 1 0 9 13 9 0 0 2 7 0 9 13 15 0 1 14 13 10 0 7 0 9 2
9 7 1 10 9 13 9 1 9 2
12 15 4 13 0 0 1 16 9 3 13 9 2
4 15 2 0 2
8 7 4 9 13 10 0 9 2
5 6 2 0 3 2
15 0 9 4 3 13 0 1 14 13 15 1 10 0 9 2
21 0 1 9 13 15 3 0 5 9 7 9 2 7 1 10 9 13 9 10 9 2
7 15 13 0 0 10 9 2
37 7 9 1 9 2 15 13 15 15 13 0 5 9 9 2 10 9 1 4 13 10 9 2 7 15 13 14 13 9 2 0 16 15 3 13 0 2
7 0 14 13 0 1 15 2
7 6 3 2 7 1 9 2
28 9 4 3 13 0 1 9 2 1 1 1 16 15 10 9 13 0 9 2 9 15 15 13 4 13 15 0 2
17 16 9 13 0 1 9 2 13 15 0 14 13 10 9 1 9 2
26 9 7 9 13 3 1 9 2 15 13 3 9 1 14 13 1 0 9 2 1 9 13 0 0 9 2
12 3 13 15 15 10 0 7 0 9 4 13 2
4 15 13 9 2
11 9 13 16 15 13 1 9 1 0 9 2
20 15 13 3 0 9 16 4 9 13 1 9 2 4 15 13 12 9 3 0 2
5 15 13 15 15 2
16 6 2 9 13 3 3 0 15 15 13 2 15 13 3 0 2
8 9 13 10 9 1 10 9 2
12 15 13 3 3 0 0 1 15 15 13 0 2
19 7 15 13 0 7 0 9 16 10 0 9 1 9 1 9 0 13 1 2
21 15 13 10 2 7 13 16 9 4 13 0 9 2 7 10 9 13 3 14 13 2
26 9 13 9 10 2 7 13 16 3 0 9 4 13 0 1 14 13 10 10 9 1 9 1 0 9 2
16 3 13 15 10 0 9 7 13 14 13 9 1 9 1 9 2
35 9 1 10 1 11 0 9 13 15 1 1 9 2 15 13 1 12 2 16 11 11 7 15 13 14 13 10 10 9 1 10 2 7 13 2
3 2 9 2
10 15 13 3 1 10 9 1 11 11 2
9 15 13 3 1 14 13 9 2 2
15 0 13 15 1 9 1 0 9 1 11 2 11 7 0 2
18 15 13 3 9 2 16 15 15 3 4 13 9 7 9 2 13 0 2
17 7 3 13 9 2 10 0 9 14 13 9 2 9 7 9 1 2
18 3 13 9 15 1 16 15 2 0 1 0 0 2 4 13 15 9 2
27 7 16 15 13 16 15 4 13 0 2 7 16 9 13 15 2 13 15 14 13 9 1 1 10 0 9 2
39 1 9 1 14 13 0 9 7 13 0 2 3 16 15 4 13 9 1 14 13 1 9 15 13 1 2 13 15 9 1 9 1 14 13 9 1 14 13 2
34 1 14 4 13 15 0 1 9 7 9 1 10 0 9 2 13 15 0 1 9 10 2 9 13 3 10 0 1 15 15 13 15 1 2
19 7 9 1 0 9 1 9 2 3 1 1 2 13 16 9 13 1 9 2
28 15 13 3 0 10 9 1 16 10 9 4 13 1 9 7 13 9 1 1 9 1 16 9 4 4 13 15 2
30 1 9 4 9 9 3 13 0 2 7 15 13 3 9 1 10 9 15 13 16 15 4 13 12 7 12 9 1 9 2
25 7 4 0 10 0 0 9 13 3 0 16 15 13 14 13 1 9 0 16 10 1 15 0 13 2
35 15 13 16 0 9 3 13 14 13 9 1 9 2 7 15 13 10 10 9 15 13 16 15 13 0 1 9 2 7 3 13 9 1 9 2
29 15 13 15 15 13 15 13 0 3 1 14 13 9 2 7 13 3 0 1 14 13 16 15 3 4 13 10 9 2
4 10 0 9 5
25 9 2 9 7 9 13 1 9 1 11 2 9 11 11 7 9 11 11 13 9 2 9 7 9 2
15 1 12 9 4 13 2 7 11 9 13 9 13 9 9 2
15 2 15 15 13 1 1 2 4 13 1 11 2 13 11 2
14 0 12 9 1 9 13 15 10 9 1 9 1 11 2
5 11 2 9 12 2
9 9 4 13 1 9 3 1 9 2
14 1 9 1 9 4 9 11 11 13 10 9 0 9 2
22 15 13 9 7 9 2 1 15 7 9 11 11 2 7 1 9 15 4 13 1 9 2
15 9 1 11 13 1 1 9 1 14 13 9 9 1 9 2
27 10 9 4 13 1 10 9 1 9 2 7 13 0 1 9 1 9 1 11 11 1 9 2 3 1 9 2
10 15 13 3 10 9 2 13 15 15 2
22 15 13 0 14 13 2 7 9 4 13 0 2 16 9 13 14 13 9 15 4 13 2
11 0 16 9 13 9 1 4 13 1 9 2
13 1 9 1 9 13 0 9 1 1 10 0 9 2
12 15 13 0 1 0 7 0 0 14 13 1 2
11 0 13 0 9 16 15 13 0 1 9 2
24 1 9 13 9 11 16 9 1 16 15 4 13 0 13 0 2 16 9 7 9 13 3 0 2
10 9 7 9 11 11 13 14 13 1 2
8 15 13 1 9 11 7 13 2
5 2 15 13 3 2
5 11 2 9 12 2
25 2 9 1 16 15 13 9 2 13 16 10 9 4 13 15 1 15 2 13 11 11 2 12 2 2
8 1 9 1 9 13 10 9 2
17 2 0 9 7 0 9 2 2 13 9 1 10 9 1 11 9 2
19 2 10 9 14 13 1 2 2 13 11 11 7 11 11 0 1 10 9 2
25 11 13 1 10 9 16 2 15 13 0 1 1 15 7 9 0 9 2 2 7 16 15 13 9 2
22 9 13 3 16 2 10 0 9 1 10 0 9 1 9 1 11 9 13 3 0 2 2
10 15 13 1 12 9 16 9 13 0 2
11 1 12 9 3 13 15 9 1 0 9 2
21 11 11 13 16 10 1 9 15 13 1 1 9 4 13 1 9 15 13 1 1 2
22 1 9 13 15 1 10 9 16 0 9 1 11 1 9 12 2 12 3 13 1 9 2
5 15 13 3 0 2
11 11 13 15 1 7 13 9 1 9 11 2
17 2 15 13 16 10 9 4 13 7 13 1 0 3 2 13 11 2
22 9 12 13 11 11 1 11 9 1 11 2 1 14 4 13 9 7 13 9 1 11 2
22 16 11 4 13 1 11 1 14 13 9 1 9 1 11 2 13 9 1 9 1 11 2
17 11 7 9 4 13 9 2 15 13 10 0 9 7 4 13 9 2
7 9 1 11 4 0 13 2
8 3 13 9 1 10 0 9 2
5 15 13 15 0 2
14 15 13 0 1 0 9 1 10 0 0 9 7 9 2
14 9 11 13 3 14 13 10 0 2 16 15 4 13 2
19 15 13 0 14 13 9 7 3 4 13 10 3 0 3 1 10 0 9 2
12 15 15 0 13 1 11 2 13 9 15 1 2
13 1 11 13 9 7 9 1 9 1 11 1 12 2
10 9 13 1 9 1 14 13 10 9 2
10 11 9 13 16 0 9 4 13 1 2
8 0 9 13 10 9 1 15 2
13 10 0 1 9 15 13 1 9 2 13 1 11 2
9 1 10 0 9 13 15 1 9 2
12 12 9 13 15 2 7 15 13 15 1 9 2
10 9 13 2 7 1 12 4 9 13 2
8 9 4 13 9 2 1 9 2
11 11 11 13 1 10 1 10 9 1 11 2
6 3 13 10 9 9 2
10 15 13 1 0 9 1 3 12 9 2
4 15 13 0 2
16 9 4 13 16 15 3 13 2 4 13 1 10 0 0 9 2
5 15 13 1 9 2
10 16 15 13 2 13 15 0 9 1 2
13 10 13 0 9 2 0 1 9 2 9 7 9 2
11 1 9 12 13 15 10 9 1 11 11 2
18 15 13 9 7 9 11 11 2 15 4 13 1 11 1 11 1 11 2
9 15 13 10 9 15 4 13 1 2
9 9 13 9 11 1 9 1 11 2
20 1 0 9 13 9 2 11 11 2 2 10 9 15 4 13 15 14 13 0 2
23 1 10 9 1 1 11 13 11 10 9 1 11 0 9 2 0 11 11 11 1 9 12 2
10 0 1 9 15 4 13 2 13 9 2
18 11 9 4 13 1 9 15 4 13 1 2 0 0 7 0 9 2 2
18 11 13 16 9 13 2 8 8 8 8 8 2 2 9 9 7 9 2
17 1 10 12 9 15 13 7 13 0 2 13 11 11 7 11 11 2
36 2 15 13 16 9 13 9 1 9 1 11 0 9 16 15 13 9 1 15 15 4 13 2 7 15 13 10 9 9 7 9 2 13 11 11 2
12 15 13 11 7 13 3 0 15 4 13 9 2
14 15 13 3 10 9 7 13 14 13 2 0 0 2 2
5 1 13 15 0 2
11 2 15 4 3 13 9 2 2 13 15 2
9 9 13 1 9 1 9 1 12 2
23 16 11 9 13 0 2 7 13 1 0 9 7 9 2 13 15 9 0 1 14 13 15 2
23 15 13 0 1 14 13 2 7 1 9 1 9 13 11 14 13 1 9 1 9 1 11 2
18 2 3 13 9 16 15 13 14 13 10 10 0 15 4 13 1 15 2
13 10 9 9 13 2 13 15 9 1 9 10 9 2
6 7 15 13 0 9 2
4 15 13 15 2
20 9 1 10 9 1 11 13 1 1 9 2 16 11 11 7 11 11 4 13 2
15 0 9 9 13 2 13 7 13 1 9 2 4 15 13 2
8 9 2 9 7 9 4 13 2
11 12 9 4 4 13 7 10 9 13 1 2
19 9 2 10 0 0 7 0 9 1 9 2 4 13 1 2 7 15 0 2
9 3 11 13 9 1 14 13 15 2
15 9 1 9 4 13 1 11 11 2 10 0 9 1 9 2
23 15 4 13 1 1 10 9 1 11 7 13 9 1 9 2 7 9 2 15 15 4 13 2
22 9 11 7 9 11 13 1 10 0 9 1 9 15 13 9 1 14 13 1 9 9 2
14 10 0 9 11 11 11 13 1 11 1 14 13 9 2
9 1 9 4 12 9 13 13 1 2
7 15 13 0 9 1 9 2
11 1 9 13 10 9 1 0 9 1 11 2
14 11 9 2 11 2 13 1 0 9 7 13 0 9 2
22 2 9 13 15 3 3 16 15 13 9 2 1 16 15 13 11 1 12 2 13 11 2
16 1 12 13 11 10 9 1 0 9 13 1 0 9 1 11 2
6 11 11 13 1 15 2
8 1 12 0 9 13 1 11 2
26 2 0 15 4 13 1 14 13 0 2 13 0 7 13 3 9 1 14 13 15 1 9 2 13 11 2
18 1 9 13 15 16 9 13 10 0 0 9 1 0 9 9 1 11 2
17 4 15 3 13 1 15 9 15 15 7 9 11 11 13 1 1 2
12 15 13 1 14 13 9 2 7 13 15 13 2
19 1 1 9 13 11 3 0 14 13 16 10 1 9 13 9 7 9 10 2
20 11 11 7 11 11 13 1 15 9 11 11 11 7 10 0 9 11 11 11 2
12 9 13 14 13 1 9 2 7 4 13 1 2
18 15 13 9 10 7 13 16 9 4 13 9 7 16 9 4 13 1 2
12 9 4 13 1 10 9 2 7 4 3 13 2
11 9 13 9 1 9 1 9 7 13 1 2
3 15 13 2
9 9 4 13 14 13 9 1 9 2
19 15 13 0 7 4 13 16 9 3 13 2 15 13 3 14 13 15 0 2
14 15 13 0 1 9 11 2 16 15 13 1 1 9 2
15 10 1 9 13 10 9 1 1 9 7 1 1 9 10 2
13 0 13 9 11 1 14 13 0 9 1 1 9 2
28 0 9 13 1 2 15 13 1 1 9 7 9 7 13 9 2 15 13 7 13 9 1 9 16 15 13 1 2
12 0 4 9 4 13 1 0 7 0 0 9 2
15 1 9 13 9 2 11 1 11 0 0 11 11 9 2 2
14 11 13 12 9 0 16 15 13 15 2 0 1 11 2
24 9 1 9 13 16 15 7 11 11 4 13 0 9 1 9 7 9 2 1 9 1 10 9 2
17 2 15 13 9 10 2 15 2 0 1 15 2 13 15 1 9 2
8 15 13 1 12 9 3 1 2
19 15 13 1 9 3 0 15 13 9 2 0 9 4 13 1 9 1 9 2
14 9 7 9 16 15 13 0 9 1 9 13 3 3 2
7 1 11 13 0 9 9 2
17 9 11 13 9 9 13 14 13 9 7 9 2 1 9 1 9 2
18 16 9 13 1 1 9 7 13 1 14 4 13 2 13 15 3 9 2
24 1 10 9 13 9 15 2 7 15 13 0 14 13 15 1 9 16 9 7 9 13 1 9 2
19 9 1 14 13 15 13 3 0 2 16 9 13 1 10 9 9 1 15 2
26 9 9 13 16 10 12 9 4 13 1 14 13 9 2 16 10 10 13 0 1 9 1 14 13 9 2
22 9 13 1 15 2 16 15 13 9 1 9 10 2 10 9 15 13 16 15 4 13 2
6 15 4 13 15 0 2
20 11 11 7 11 11 4 13 10 0 9 1 10 9 2 16 9 13 1 9 2
20 9 13 3 1 16 9 1 9 13 0 1 8 9 1 14 13 15 1 9 2
15 1 10 9 1 9 7 9 7 9 1 0 9 13 15 2
8 15 13 15 2 15 13 15 2
8 10 9 13 9 1 14 13 2
11 1 9 13 9 1 1 9 1 11 11 2
20 2 15 13 1 9 1 16 0 9 13 15 2 1 9 4 15 13 1 9 2
25 16 15 13 3 1 1 15 2 13 15 1 14 13 14 13 9 0 2 14 13 9 2 13 11 2
17 15 13 16 15 3 13 14 13 0 2 15 13 15 15 3 3 2
22 2 15 4 13 1 14 13 9 16 15 13 1 11 2 15 13 9 10 2 13 11 2
12 15 13 1 1 16 15 4 13 10 0 9 2
13 2 15 4 3 13 3 0 9 1 10 9 1 2
16 1 9 4 11 1 9 13 9 2 7 4 15 7 15 13 2
7 15 4 13 0 1 9 2
21 7 15 4 13 0 1 9 2 13 15 13 1 9 2 1 9 1 3 10 9 2
23 9 13 3 16 15 13 15 14 13 1 2 3 1 0 9 2 16 15 13 7 9 13 2
18 9 11 13 0 9 1 9 2 7 1 0 9 13 15 1 9 10 2
8 2 13 15 3 2 13 11 2
12 15 13 1 9 2 10 9 1 10 0 9 2
16 9 13 0 2 9 13 15 0 1 9 2 16 15 4 13 2
8 15 13 15 1 9 1 9 2
11 7 9 4 13 7 13 1 9 1 9 2
10 10 0 9 4 0 13 1 1 11 2
16 11 13 3 10 9 1 14 13 10 0 9 2 7 4 13 2
26 15 13 9 1 12 0 9 2 13 15 3 1 9 7 13 15 1 2 3 16 9 13 1 9 9 2
13 1 10 0 2 0 9 7 9 4 15 13 9 2
11 2 15 13 3 1 15 0 9 0 9 2
13 15 13 15 2 7 1 9 1 9 13 15 13 2
20 15 13 0 14 13 1 9 1 9 2 1 14 13 9 1 15 15 13 15 2
19 3 0 15 13 1 9 2 3 0 13 9 1 14 4 13 2 13 11 2
16 2 15 4 13 16 15 3 4 4 13 1 16 9 13 15 2
11 2 10 9 4 15 13 1 2 13 11 2
11 9 11 13 0 1 10 10 9 1 9 2
12 2 15 13 3 3 14 13 1 15 10 9 2
20 10 12 9 13 1 10 0 9 2 16 15 4 13 0 9 1 10 0 9 2
22 3 0 1 9 9 4 10 12 9 13 1 9 2 9 4 13 2 15 13 9 1 2
9 9 2 1 0 9 2 4 13 2
8 10 10 9 13 1 14 13 2
21 11 11 7 10 0 9 13 1 1 14 13 2 16 15 13 14 13 1 9 10 2
11 9 13 15 1 12 9 2 1 10 9 2
11 9 13 1 16 9 3 4 13 1 9 2
11 9 7 10 0 4 13 1 10 10 9 2
13 15 13 9 2 9 11 11 11 13 1 10 9 2
9 15 13 15 1 2 10 9 3 2
18 16 11 11 13 1 7 13 1 9 2 13 15 15 13 1 1 9 2
11 2 15 13 3 15 15 13 2 13 15 2
8 9 11 13 1 9 1 9 2
9 1 3 10 9 13 15 15 0 2
25 15 13 1 3 15 13 3 9 1 9 2 1 10 9 15 13 16 15 4 13 0 1 0 9 2
21 1 9 13 15 1 9 0 9 2 3 13 15 3 10 12 9 9 13 1 9 2
26 1 9 7 1 10 0 9 11 11 11 9 1 9 13 15 3 10 0 9 9 4 13 15 1 9 2
23 11 11 13 16 15 1 9 3 4 13 1 2 16 15 3 13 14 13 9 15 4 13 2
7 7 12 9 13 15 1 2
9 15 13 1 10 9 7 4 13 2
12 2 15 13 9 1 14 13 1 2 13 15 2
6 2 4 15 13 9 2
9 2 15 15 13 3 2 13 11 2
24 12 1 12 9 1 11 4 13 2 7 9 13 1 1 9 2 15 4 13 1 10 0 9 2
8 9 13 1 0 9 10 9 2
26 9 1 9 2 9 11 11 11 2 13 1 10 12 9 1 9 2 3 9 1 11 11 7 11 11 2
19 15 4 13 1 14 13 9 1 9 16 9 13 15 2 7 13 1 9 2
13 10 0 1 9 9 4 13 2 13 11 1 9 2
26 15 13 3 3 9 4 13 1 14 13 2 16 11 1 9 13 12 9 1 9 1 14 13 1 9 2
11 10 0 9 13 3 1 9 1 0 9 2
19 2 15 13 0 9 1 14 13 1 15 15 13 1 11 2 13 11 11 2
9 15 13 3 9 15 3 4 13 2
18 3 1 11 11 13 15 1 1 14 13 1 10 0 9 1 12 9 2
9 15 13 0 2 1 14 13 15 2
18 2 15 4 13 15 0 2 13 11 2 1 14 13 16 15 13 0 2
13 15 13 10 12 9 15 13 1 15 1 10 9 2
20 15 15 13 1 4 13 2 10 10 4 13 0 1 12 9 1 14 13 9 2
16 2 11 13 15 3 10 9 1 14 13 1 1 2 13 15 2
12 11 13 1 9 1 9 15 13 3 0 1 2
17 2 11 11 13 10 3 0 9 2 15 3 13 15 2 13 15 2
11 11 13 0 1 11 1 10 9 7 9 2
14 1 12 13 11 9 1 16 9 1 11 4 13 1 2
5 9 13 1 9 2
8 15 4 13 12 9 1 9 2
10 9 11 11 4 13 10 9 1 11 2
5 13 15 1 3 2
10 15 13 9 1 10 0 9 1 11 2
13 11 13 16 15 13 0 7 13 15 1 1 9 2
8 9 13 9 16 9 13 15 2
23 2 15 2 9 2 15 13 0 0 9 1 11 2 15 13 3 0 15 13 0 10 9 2
15 10 9 13 11 11 11 9 7 13 16 15 3 4 13 2
12 10 9 1 9 1 11 13 1 9 1 11 2
15 9 15 13 1 2 13 1 10 9 1 10 9 1 9 2
4 10 12 13 2
5 11 13 9 0 2
25 15 4 13 1 1 0 9 1 9 1 11 7 13 3 1 9 1 10 16 15 13 1 7 13 2
16 15 13 3 3 0 16 15 4 4 13 15 15 13 1 11 2
17 15 13 3 1 16 9 3 4 4 13 2 16 15 4 13 1 2
2 9 5
12 15 4 13 15 15 4 13 11 10 0 9 5
12 11 13 1 1 10 9 1 9 7 0 9 2
5 3 13 15 1 2
10 15 13 9 2 0 13 15 9 12 2
6 1 13 15 0 9 2
11 9 13 1 15 0 9 7 13 0 1 2
16 1 10 0 9 13 15 15 1 9 2 1 9 1 1 9 2
4 15 13 0 2
12 3 13 15 1 16 10 9 4 13 1 15 2
9 11 11 11 13 12 9 7 0 2
13 0 9 4 15 13 1 16 15 13 10 0 9 2
35 15 4 13 9 1 9 2 1 15 10 2 13 9 2 13 15 1 9 2 13 1 16 15 3 13 14 13 16 9 13 1 9 1 9 2
16 9 2 15 0 13 3 0 2 13 0 7 0 1 1 9 2
19 9 2 15 13 14 13 15 0 1 7 13 1 15 2 13 3 3 1 2
12 3 13 15 11 7 9 15 4 13 1 15 2
5 11 13 3 0 2
8 15 13 3 11 13 15 1 2
6 15 4 4 13 15 2
24 3 4 3 9 1 11 13 15 1 9 15 4 13 1 3 16 9 13 0 7 0 1 9 2
17 9 10 13 9 1 15 15 13 2 15 15 13 9 15 3 13 2
4 15 13 15 2
20 2 15 13 0 15 4 4 13 16 15 13 0 0 1 1 15 2 13 11 2
18 1 9 13 10 0 10 9 1 14 13 1 1 9 15 13 0 1 2
13 9 7 9 13 9 1 14 13 16 15 13 9 2
11 11 13 15 15 13 1 14 13 9 1 2
12 0 12 0 13 1 9 2 7 13 3 1 2
10 9 13 10 9 0 16 11 13 15 2
9 9 13 1 9 2 0 1 9 2
8 11 4 13 9 0 1 15 2
7 9 13 1 9 1 11 2
15 15 13 10 0 1 9 2 7 15 13 0 1 14 13 2
15 16 15 4 13 15 10 2 4 15 13 15 3 2 9 2
2 11 5
19 15 13 9 1 16 9 13 1 1 9 7 13 15 1 1 10 0 9 2
12 7 15 13 10 9 1 0 1 9 1 9 2
11 15 13 1 10 0 9 1 9 1 9 2
13 1 15 15 13 1 14 13 2 13 10 0 9 2
13 15 13 9 1 15 2 7 13 15 1 1 9 2
5 9 13 1 11 2
17 9 13 15 1 9 2 3 11 0 1 9 4 13 1 10 9 2
17 15 13 15 3 0 15 13 2 7 13 10 12 9 0 9 10 2
6 10 12 9 13 11 2
11 10 1 10 0 4 13 16 15 13 1 2
11 1 9 13 15 0 1 1 9 1 11 2
9 10 9 1 12 9 1 10 9 2
10 9 1 0 9 1 11 7 0 9 2
5 9 13 1 9 2
7 12 9 15 13 0 9 2
12 9 13 1 16 9 13 1 0 9 1 9 2
14 10 9 1 12 0 9 2 15 13 1 9 1 9 2
3 0 9 2
8 7 15 13 3 15 15 13 2
5 9 13 0 9 2
13 0 4 15 13 1 10 0 9 2 7 13 0 2
7 15 13 3 1 0 9 2
18 16 15 13 12 9 4 15 3 13 13 1 0 0 9 1 9 10 2
7 1 10 9 13 15 9 2
18 15 13 10 0 9 15 4 13 2 15 4 13 15 1 15 1 15 2
2 9 5
13 9 13 9 2 7 13 1 9 0 9 1 9 2
21 16 15 13 1 9 13 15 0 1 10 10 9 10 2 7 15 13 0 1 9 2
15 11 13 15 0 9 4 13 15 1 9 16 15 13 1 2
15 1 10 13 15 0 1 2 7 13 14 13 1 15 0 2
6 9 13 3 10 9 2
13 13 10 0 9 16 15 13 3 15 0 13 1 2
6 15 13 9 1 9 2
8 15 13 0 9 1 11 9 2
15 11 13 10 0 9 1 9 2 0 9 7 10 0 9 2
21 15 4 3 13 1 9 2 7 15 13 3 3 0 14 13 1 16 15 13 9 2
11 15 13 3 3 0 9 16 9 13 1 2
14 11 13 0 0 2 15 13 0 9 2 15 4 13 2
18 1 12 9 13 9 1 11 1 16 11 4 4 13 1 10 10 9 2
28 7 15 13 3 2 1 9 1 11 9 2 16 15 13 1 1 15 16 3 15 13 0 15 15 4 13 1 2
6 15 13 10 0 9 2
13 9 13 3 1 15 9 2 11 9 13 0 0 2
16 0 3 0 13 9 14 13 9 2 7 9 13 15 3 3 2
14 10 9 13 15 9 15 13 11 1 9 2 1 9 2
9 7 15 7 9 4 13 1 9 2
18 1 9 13 15 10 9 3 0 16 9 13 15 1 1 9 10 9 2
5 11 13 0 3 2
14 1 9 1 9 13 15 16 15 13 15 1 1 9 2
7 15 13 10 9 1 9 2
16 3 13 15 1 9 1 9 2 9 1 9 2 16 9 13 2
9 9 13 1 14 13 10 0 9 2
6 9 13 3 1 15 2
7 15 13 3 9 7 9 2
16 11 13 3 10 9 1 14 13 15 15 0 13 1 9 10 2
8 7 15 13 3 0 1 9 2
5 7 15 13 9 2
14 1 0 1 0 9 1 11 9 13 11 11 11 9 2
12 15 13 15 13 9 0 2 3 16 9 13 2
7 9 4 3 3 0 13 2
25 2 10 9 13 9 16 15 3 13 15 15 4 13 2 7 16 15 3 13 15 1 14 13 15 2
12 15 13 3 3 15 7 10 10 2 13 15 2
7 1 9 13 15 12 9 2
14 1 10 3 0 9 13 15 0 1 7 9 7 9 2
18 10 0 9 13 16 9 1 9 13 1 9 2 7 10 9 13 9 2
20 16 15 13 1 9 2 13 9 7 14 13 0 9 7 13 10 9 1 9 2
9 11 4 3 13 16 15 4 13 2
12 15 13 11 1 9 9 1 14 13 0 9 2
17 10 9 13 11 15 16 15 3 13 9 1 16 15 4 13 15 2
14 9 13 3 0 3 0 9 15 13 1 9 1 9 2
10 2 15 4 0 13 16 15 13 0 2
16 15 4 3 13 0 1 14 13 1 9 15 3 13 15 0 2
7 7 15 13 3 11 3 2
10 15 1 9 1 2 15 13 15 3 2
9 3 4 15 3 13 15 1 9 2
14 15 4 13 16 15 4 13 2 7 15 13 15 3 2
11 15 13 3 1 10 9 16 15 13 11 2
8 9 13 3 3 1 10 9 2
23 9 11 11 11 2 15 13 9 1 10 10 3 12 9 1 9 2 13 1 10 15 13 2
10 9 13 9 1 9 1 9 1 9 2
6 11 13 9 1 9 2
17 1 10 9 13 15 0 14 13 1 9 9 2 16 15 4 13 2
13 0 13 15 0 2 10 9 1 16 15 13 0 2
23 0 1 13 15 3 16 15 4 13 16 15 13 3 0 15 13 1 2 3 0 9 13 2
5 7 15 13 15 2
27 2 10 9 13 0 1 10 2 7 15 13 3 9 1 14 13 16 11 13 0 1 1 10 2 13 11 2
13 9 2 15 1 9 4 13 9 2 13 11 0 2
12 15 13 0 0 16 15 4 13 1 11 9 2
15 10 0 9 13 10 9 2 10 9 15 13 9 1 9 2
29 2 3 15 13 9 2 13 15 15 0 1 16 15 4 13 9 0 1 15 16 15 13 9 1 0 2 13 15 2
5 13 11 1 15 2
7 13 16 15 13 1 15 2
9 15 13 3 0 15 4 13 15 2
2 9 5
18 11 13 10 9 15 13 10 9 1 12 9 1 1 9 3 1 9 2
5 15 4 13 9 2
18 11 13 11 9 1 10 9 15 13 10 0 9 1 9 1 11 9 2
22 2 16 11 3 13 15 1 11 9 2 13 15 15 0 1 16 9 4 13 1 15 2
17 15 13 0 1 14 13 16 15 4 13 15 3 0 2 13 11 2
8 3 13 3 11 7 9 15 2
8 1 1 11 13 15 0 1 2
15 9 13 1 9 1 10 0 9 2 7 15 13 0 9 2
11 1 9 13 9 9 10 0 9 1 9 2
7 15 13 0 0 9 0 2
29 2 9 13 0 9 7 9 13 1 15 15 4 4 13 1 0 2 7 13 3 9 2 13 11 12 9 0 9 2
19 15 13 15 15 13 9 1 9 1 7 9 7 9 16 15 13 12 9 2
8 9 13 11 3 0 15 13 2
17 13 15 1 1 1 9 16 9 13 2 13 14 13 9 1 9 2
16 9 13 12 9 2 15 4 3 13 15 1 3 9 13 1 2
17 9 4 13 15 16 16 15 13 15 2 13 9 1 14 13 15 2
17 9 13 15 4 4 13 1 10 10 9 2 1 14 4 13 15 2
8 9 13 15 1 10 0 9 2
7 2 15 4 3 13 15 2
8 15 13 0 1 14 13 11 2
11 7 15 4 13 1 9 16 15 13 15 2
4 3 13 9 2
11 13 15 10 10 15 13 9 7 13 9 2
15 1 0 9 13 11 9 1 11 16 15 13 15 1 9 2
6 15 13 9 1 9 2
17 9 13 10 0 9 2 15 13 14 13 15 0 1 15 1 15 2
9 15 4 3 13 15 1 1 15 2
2 11 5
22 2 1 1 15 15 4 13 1 1 10 9 4 15 3 13 10 9 1 9 1 11 2
27 16 15 4 4 13 10 9 1 15 15 3 4 4 13 1 14 13 1 9 4 15 3 1 9 13 1 2
27 1 1 1 3 12 9 3 13 9 16 9 15 3 13 1 9 3 4 13 1 12 9 16 15 4 13 2
33 1 3 12 9 3 13 15 10 9 15 13 1 16 15 3 4 13 9 15 3 13 1 9 1 16 3 9 4 13 9 1 9 2
14 15 4 13 0 1 9 1 11 1 0 1 12 9 2
26 15 4 3 13 16 15 4 13 9 13 1 10 9 2 7 14 13 16 15 3 4 13 15 13 0 2
9 3 11 11 2 11 1 9 2 2
7 11 13 3 9 13 15 2
14 10 9 13 15 9 1 10 0 9 1 9 1 9 2
21 9 4 13 2 0 1 9 1 9 2 7 13 0 9 1 1 9 3 1 9 2
16 1 13 12 0 9 15 4 13 1 9 1 16 15 4 13 2
9 1 14 13 15 15 13 1 9 2
20 9 13 12 7 12 9 0 2 7 4 13 15 10 16 9 13 1 1 11 2
18 9 13 1 9 3 3 0 15 13 9 1 2 7 13 15 13 0 2
12 1 9 13 9 0 0 9 2 7 9 13 2
14 1 10 0 13 15 1 9 2 13 0 7 13 0 2
12 15 13 1 9 1 9 2 13 9 1 9 2
19 11 7 9 13 1 9 1 9 2 15 13 0 1 1 14 13 1 9 2
21 16 11 10 0 9 13 1 10 9 1 2 13 15 1 9 2 1 9 7 9 2
24 15 13 0 1 16 15 4 13 14 13 1 9 1 9 9 7 16 9 4 13 3 0 9 2
7 9 13 0 7 0 1 2
5 9 13 3 15 2
10 2 15 4 13 1 1 13 15 10 2
10 15 4 13 10 9 14 13 1 9 2
4 15 13 9 2
8 1 9 1 11 13 9 0 2
16 10 9 13 16 15 0 13 9 1 9 7 9 1 11 9 2
20 2 15 13 9 1 16 9 13 1 9 7 0 9 1 0 9 2 13 9 2
10 15 13 16 9 3 13 3 15 13 2
9 10 9 13 11 1 9 1 9 2
5 15 13 12 9 2
5 9 13 1 9 2
16 2 9 13 15 13 16 15 4 13 0 2 13 11 1 9 2
7 15 13 3 3 0 0 2
25 13 3 16 9 0 9 4 13 15 2 16 11 4 13 9 1 14 13 9 1 14 13 9 10 2
14 0 1 9 13 9 1 11 16 15 3 4 13 0 2
19 9 13 1 9 2 13 15 1 2 7 13 15 4 13 9 1 10 9 2
8 11 13 15 3 1 1 9 2
24 2 16 15 4 13 15 10 4 15 13 15 3 2 9 2 13 11 2 7 13 14 13 15 2
23 1 10 9 13 11 9 1 9 2 13 15 1 2 7 13 15 1 1 9 7 1 9 2
9 11 13 1 7 13 9 1 9 2
8 9 13 16 3 13 15 3 2
5 15 4 13 9 2
11 7 15 13 15 16 9 15 13 13 9 2
7 7 10 9 13 3 1 2
9 9 13 15 2 13 2 13 15 2
14 16 15 0 13 11 1 9 2 13 15 3 15 13 2
4 9 13 3 2
13 2 15 13 1 16 15 3 13 15 2 13 9 2
7 7 3 13 15 3 0 2
4 9 13 0 2
5 15 4 13 0 2
6 2 13 11 1 15 2
7 13 16 15 13 1 15 2
9 15 13 3 0 15 4 13 15 2
6 3 13 9 1 9 2
21 16 15 13 0 2 0 9 1 15 15 13 9 2 13 11 9 13 15 1 9 2
10 16 9 4 13 9 2 13 15 0 2
5 3 13 15 0 2
13 13 2 13 0 9 1 9 7 13 9 0 9 2
16 10 9 13 9 1 0 9 1 15 16 15 13 1 1 9 2
10 3 13 15 16 15 13 1 1 9 2
7 16 9 13 0 1 9 2
23 16 15 4 13 10 9 1 14 13 10 0 9 2 13 1 9 2 7 13 15 1 9 2
13 3 13 9 15 0 1 9 1 16 9 13 15 2
18 2 9 13 10 0 9 2 15 13 14 13 15 0 1 15 1 15 2
9 15 4 3 13 15 1 1 15 2
18 7 15 13 3 3 3 0 9 7 10 0 9 13 15 2 13 11 2
12 11 9 13 3 0 1 14 13 15 15 13 2
15 9 11 11 11 13 15 1 10 0 9 1 9 1 9 2
10 10 0 9 15 13 0 1 14 13 2
13 15 13 9 1 9 2 7 13 3 1 11 11 2
21 10 9 13 9 16 11 9 13 0 2 7 4 13 16 15 13 1 9 1 9 2
9 15 13 3 16 9 13 10 9 2
14 2 15 13 9 16 15 4 13 15 15 0 4 13 2
21 15 13 0 1 16 15 4 13 3 0 1 15 2 7 0 1 16 9 4 13 2
21 7 15 13 15 3 2 7 13 3 15 0 0 1 15 1 15 15 13 1 9 2
7 0 13 11 0 1 11 2
10 11 11 11 1 9 13 10 0 9 2
14 15 13 1 10 0 1 1 9 2 7 1 1 11 2
9 10 0 9 13 15 1 1 11 2
18 3 13 9 0 13 7 13 1 9 2 16 9 13 1 9 1 9 2
8 11 13 15 1 0 7 0 2
25 15 11 3 13 2 13 16 9 3 13 16 15 13 1 15 15 1 2 16 15 4 13 9 1 2
7 1 9 13 15 1 9 2
11 9 2 11 2 1 11 11 13 11 9 2
9 15 13 1 15 1 7 1 3 2
37 2 15 13 3 0 15 13 16 15 13 15 2 16 15 4 13 9 1 9 7 15 2 7 15 13 10 1 15 15 13 3 15 0 13 15 1 2
12 15 13 0 0 1 14 13 15 2 13 11 2
10 15 13 0 16 9 13 9 1 9 2
6 9 13 3 0 9 2
21 2 1 10 9 15 13 13 15 0 16 11 4 13 15 15 4 13 2 13 11 2
6 9 13 0 7 0 2
10 1 0 7 0 9 13 11 0 0 2
5 15 13 1 9 2
12 3 1 11 13 15 1 11 2 11 2 11 2
3 9 9 2
12 0 4 9 1 10 0 13 1 9 1 9 2
12 11 13 9 7 13 3 1 0 9 1 9 2
6 1 13 15 1 9 2
7 3 13 9 1 9 0 2
6 15 4 4 13 15 2
7 7 15 13 15 15 13 2
10 9 13 1 10 0 1 9 1 9 2
15 9 13 3 9 1 9 1 9 16 15 13 1 1 11 2
23 11 7 9 13 9 1 14 13 2 13 9 2 13 9 2 13 9 2 13 15 1 9 2
4 13 1 9 2
10 2 15 13 3 3 0 14 13 9 2
23 10 10 13 1 0 9 15 4 13 1 9 2 15 4 13 1 16 9 3 13 0 9 2
12 15 13 3 3 0 14 13 1 2 13 11 2
6 15 13 15 1 11 2
16 1 11 9 13 9 11 11 1 12 0 9 14 13 9 1 2
8 7 9 13 15 0 1 10 2
10 10 1 9 13 15 1 10 0 9 2
6 9 13 9 1 9 2
5 0 9 7 9 2
25 2 15 13 1 10 10 9 15 13 1 9 2 13 9 1 11 2 7 13 10 0 9 1 15 2
14 9 10 13 0 2 9 1 10 0 2 7 9 13 2
14 1 0 9 13 9 0 1 16 15 3 13 1 9 2
11 11 4 13 1 9 9 1 9 0 9 2
12 1 9 1 10 12 13 9 0 2 9 0 2
9 15 13 2 7 13 0 13 0 2
2 0 2
2 0 2
14 9 11 13 0 1 3 15 13 3 0 1 1 9 2
8 2 13 3 9 2 13 9 2
17 9 13 3 3 0 1 15 2 13 15 2 7 13 15 13 0 2
5 15 13 0 3 2
5 9 2 13 9 2
20 15 13 15 3 1 16 10 0 9 4 13 1 15 10 16 15 13 12 9 2
10 11 13 12 9 0 16 9 13 1 2
21 9 13 0 7 0 1 2 7 11 13 15 13 3 10 9 1 14 13 1 9 2
8 15 13 3 0 2 3 0 2
35 15 13 3 0 1 15 15 4 13 9 16 15 13 3 15 13 1 2 0 1 16 9 4 13 15 2 7 15 13 15 3 1 10 9 2
11 9 13 15 13 10 9 1 9 1 15 2
13 1 12 1 9 13 15 2 0 2 0 9 2 2
32 15 13 16 15 13 0 16 9 13 0 2 3 4 15 13 3 15 15 13 2 16 15 13 1 7 13 15 1 10 0 9 2
15 2 4 15 3 13 0 9 7 9 2 4 15 13 0 2
9 7 15 13 3 3 0 7 0 2
12 15 13 1 9 16 15 4 4 13 0 9 2
15 15 13 9 1 16 15 3 13 0 10 9 2 13 11 2
4 15 13 9 2
13 11 9 13 10 10 9 1 9 1 11 7 9 2
23 15 13 9 3 4 13 10 9 2 7 16 9 13 0 3 1 14 13 9 1 15 10 2
18 7 9 13 16 9 2 11 9 2 3 13 10 9 1 9 1 9 2
10 15 13 16 10 9 13 1 12 9 2
18 9 13 15 13 0 9 16 9 13 0 1 9 1 0 9 1 9 2
11 15 13 9 13 0 1 9 1 9 9 2
15 0 9 1 9 13 9 9 7 13 9 13 1 0 9 2
19 11 7 9 13 3 15 13 0 16 9 13 10 10 9 1 9 1 15 2
37 2 15 13 3 0 1 15 15 4 13 9 16 15 13 3 15 13 1 2 0 1 16 9 4 13 15 2 7 15 13 15 3 1 10 0 9 2
9 7 15 13 9 15 13 9 9 2
9 16 9 0 13 2 13 15 15 2
15 1 10 9 4 9 1 11 7 9 13 10 0 10 9 2
15 7 15 13 10 0 9 15 4 13 3 9 13 15 1 2
25 10 1 15 13 9 1 15 15 13 4 13 15 2 13 15 1 1 9 1 9 10 2 7 13 2
17 15 13 15 2 1 9 1 14 13 9 7 1 15 10 7 9 2
11 9 13 0 0 16 9 13 15 0 0 2
6 9 1 9 15 13 2
21 16 15 13 16 15 13 2 13 0 2 13 1 9 1 3 2 13 0 14 13 2
14 16 15 13 14 13 15 0 9 1 10 9 1 9 2
12 15 13 1 10 0 9 1 16 9 4 13 2
6 15 13 1 10 9 2
24 9 15 9 13 1 1 14 13 9 2 13 10 10 15 4 13 1 9 1 9 1 10 9 2
17 16 0 13 9 1 7 9 7 9 2 13 9 0 0 1 9 2
15 9 13 16 9 9 13 1 9 1 11 0 9 1 9 2
6 9 13 9 1 0 2
6 3 13 3 9 9 2
26 3 16 0 13 16 12 0 9 1 10 0 13 3 1 10 9 15 13 0 0 9 7 13 15 3 2
12 1 9 4 10 9 13 1 2 10 9 2 2
8 0 9 13 9 1 9 9 2
20 15 13 1 16 9 13 0 1 0 9 2 16 15 13 15 1 0 7 0 2
8 10 9 13 10 9 1 9 2
12 9 13 0 16 11 9 13 9 1 0 9 2
11 9 13 9 14 13 9 1 9 1 9 2
4 3 13 9 2
6 3 13 3 9 9 2
6 9 9 13 0 9 2
23 9 1 9 1 10 9 15 13 0 0 2 15 13 1 9 2 0 9 2 9 1 9 2
12 10 9 13 15 1 1 11 1 10 9 9 2
4 15 13 9 2
5 13 1 0 9 2
27 13 1 10 9 16 9 13 15 13 0 0 1 15 2 7 13 14 13 1 11 11 7 10 0 9 3 2
18 1 12 9 2 3 0 1 16 9 1 9 13 3 1 12 0 9 2
8 1 9 9 2 0 9 12 2
5 2 13 1 9 2
8 13 0 0 1 10 7 10 2
3 0 9 2
8 13 16 15 13 0 1 15 2
13 13 16 15 4 13 10 0 9 7 13 0 2 2
13 1 9 13 9 9 1 9 7 13 15 1 9 2
8 7 9 13 3 0 0 9 2
15 16 9 13 3 15 13 9 2 13 9 16 15 13 9 2
20 16 9 13 0 7 13 0 9 1 9 2 13 9 15 13 9 1 10 9 2
6 15 4 3 13 15 2
8 15 13 0 1 14 13 11 2
2 9 5
35 2 15 13 3 0 2 7 13 10 9 1 9 15 13 9 14 13 14 13 15 2 3 16 9 13 16 9 13 3 1 15 9 1 9 2
9 3 0 4 10 9 9 13 15 2
21 13 3 9 3 3 0 9 1 15 2 15 3 13 10 9 2 7 15 13 9 2
17 11 4 13 9 1 9 2 7 13 16 9 4 13 15 15 13 2
15 11 4 13 1 9 1 9 2 7 0 4 3 13 15 2
6 9 13 1 9 0 2
7 3 4 15 13 1 9 2
20 10 9 1 9 12 13 9 1 9 1 9 2 15 13 1 10 9 1 9 2
7 15 13 15 15 4 13 2
11 1 0 9 13 9 16 15 13 10 9 2
11 15 4 13 15 1 14 13 15 1 15 2
10 15 13 1 14 13 15 1 1 9 2
21 2 15 13 0 0 2 7 13 10 9 1 9 15 15 3 4 13 1 0 9 2
29 1 14 4 13 1 10 9 1 0 9 13 15 3 1 9 2 15 13 3 15 13 3 9 13 2 13 11 9 2
6 15 13 10 0 9 2
10 9 13 9 3 15 4 13 1 9 2
12 9 13 15 4 13 0 2 7 0 7 0 2
5 1 10 0 9 2
12 7 15 13 3 3 0 9 4 13 1 9 2
10 9 13 1 9 1 16 15 4 13 2
7 13 16 15 4 13 0 2
28 7 1 16 15 13 10 9 1 15 15 4 13 2 13 15 16 9 4 13 14 13 9 1 11 16 15 13 2
17 2 15 13 0 1 15 2 2 13 9 2 7 13 15 10 9 2
7 2 13 0 1 9 2 2
22 3 13 9 1 2 1 14 13 15 15 13 0 2 14 13 2 13 1 9 1 9 2
24 15 13 11 2 7 3 1 1 2 16 9 13 0 2 4 9 13 9 1 10 9 1 9 2
7 3 13 15 9 13 0 2
8 1 1 9 13 9 1 11 2
13 15 13 15 9 2 3 1 1 9 4 15 13 2
16 1 15 15 13 1 14 13 1 9 1 9 2 13 15 1 2
16 15 13 12 9 7 4 13 15 1 14 13 15 1 9 10 2
4 3 13 9 2
5 11 13 1 9 2
10 1 15 15 13 1 1 9 13 9 2
18 2 15 4 13 1 1 10 9 2 15 4 13 15 2 13 10 9 2
14 15 13 9 1 15 16 9 10 7 15 13 3 0 2
7 9 13 1 9 1 9 2
9 11 13 1 10 9 15 15 13 2
13 2 15 13 1 10 0 9 1 16 9 4 13 2
6 15 13 1 10 9 2
10 9 15 13 1 9 13 9 1 9 2
9 15 13 14 13 15 2 13 9 2
8 7 9 13 3 1 14 13 2
9 1 1 11 9 13 15 1 9 2
10 15 13 2 7 4 11 13 1 9 2
8 13 15 16 11 3 13 3 2
12 11 13 12 9 16 15 0 4 13 1 9 2
16 1 9 13 15 7 9 0 9 2 7 15 13 3 0 1 2
10 11 13 3 0 9 3 7 13 9 2
9 9 11 11 1 11 11 13 9 2
13 15 13 3 10 9 1 9 15 4 13 0 9 2
6 2 15 13 1 9 2
9 1 3 4 15 13 10 9 1 2
10 1 3 2 13 11 1 10 0 9 2
33 10 0 9 13 1 9 10 1 9 15 13 15 0 0 2 7 11 13 9 1 16 15 4 13 7 13 9 3 1 3 1 9 2
6 15 13 14 13 0 2
5 11 11 13 9 2
2 13 2
6 11 13 0 1 9 2
5 3 13 15 0 2
7 15 13 3 1 9 9 2
8 7 15 13 1 9 1 9 2
19 15 13 1 10 1 1 9 16 9 15 13 1 9 1 9 10 13 0 2
11 9 13 3 1 0 9 1 9 1 9 2
16 1 9 13 9 2 15 13 0 0 9 2 0 3 1 9 2
18 2 15 13 16 15 13 0 9 1 15 2 1 9 2 9 7 9 2
12 15 13 15 3 16 11 4 13 9 1 15 2
13 15 13 3 16 15 13 3 0 3 2 13 11 2
16 9 13 9 4 13 1 1 9 16 0 9 3 13 0 9 2
14 2 10 9 4 3 13 3 3 3 16 9 13 0 2
20 4 15 13 15 4 15 13 10 9 1 10 9 2 1 14 13 1 0 9 2
9 7 15 13 3 16 15 13 0 2
5 9 12 13 15 2
10 11 13 3 3 9 14 13 15 0 2
7 9 13 9 1 9 10 2
11 11 11 13 0 0 1 10 0 0 9 2
19 15 15 4 13 2 4 13 15 0 2 4 13 9 1 14 13 15 10 2
6 10 0 9 13 9 2
8 3 13 15 1 1 11 9 2
5 9 13 11 12 2
16 3 13 11 14 13 3 2 3 13 15 15 1 15 15 13 2
9 9 10 9 13 15 0 1 9 2
16 0 13 9 1 9 2 7 9 13 3 0 10 12 0 9 2
14 1 9 2 12 9 0 2 13 3 9 1 11 9 2
10 9 13 10 10 2 7 9 10 10 2
17 2 13 15 10 9 7 9 15 13 3 0 2 13 9 7 9 2
20 3 13 15 3 3 2 2 13 15 1 10 1 10 0 9 15 13 1 9 2
14 11 11 4 13 0 2 0 9 2 14 13 9 1 2
6 7 15 13 15 3 2
17 2 0 9 13 15 1 15 1 9 0 16 15 13 0 1 9 2
6 11 13 10 10 9 2
7 15 13 10 3 0 9 2
8 15 13 15 1 9 1 15 2
7 15 13 0 1 15 3 2
12 15 4 13 16 15 4 13 1 15 15 13 2
7 11 4 0 13 1 15 2
6 3 4 9 13 3 2
12 7 13 9 3 16 15 4 4 13 1 9 2
14 11 11 2 9 1 9 1 11 2 13 3 1 9 2
11 10 1 15 15 3 13 2 13 0 9 2
16 15 13 11 15 10 0 1 11 4 13 1 11 1 9 10 2
13 4 15 3 13 9 7 9 2 4 15 13 0 5
4 9 11 11 5
7 15 1 15 4 13 9 2
7 15 13 0 14 13 15 2
20 9 7 9 13 9 1 14 13 9 16 15 13 16 10 9 4 13 1 9 2
27 7 9 7 9 1 9 7 9 13 3 3 9 1 16 15 4 0 14 13 9 1 11 9 2 13 11 2
31 2 7 15 13 0 16 15 3 13 1 11 9 1 9 1 15 16 15 3 13 9 1 2 7 16 15 0 9 13 0 2
22 1 9 4 15 0 1 0 9 2 7 10 9 7 9 15 13 15 1 10 10 9 2
17 9 4 1 9 13 10 9 1 9 1 3 11 3 13 1 9 2
26 15 4 3 4 13 1 9 1 9 1 9 2 1 14 4 13 1 9 9 1 14 13 1 9 10 2
5 4 9 4 13 2
25 9 13 3 0 14 13 9 2 7 10 0 13 10 9 1 14 13 1 1 9 15 13 0 1 2
17 15 4 9 13 16 9 15 11 13 9 1 4 13 1 10 9 2
40 2 9 9 13 1 2 1 0 9 1 9 7 10 0 9 15 13 16 9 13 16 15 4 13 2 13 9 15 4 13 1 16 15 4 13 1 9 10 9 2
22 10 9 13 1 9 1 9 7 9 2 3 3 9 1 3 9 7 9 13 15 3 2
16 9 13 3 9 1 9 2 9 2 9 7 1 10 9 9 2
19 9 13 14 13 9 2 7 13 15 16 15 13 0 1 0 1 11 9 2
5 4 15 13 0 2
19 2 15 13 15 2 7 0 9 4 13 0 0 9 16 15 13 1 9 2
26 16 15 4 13 1 10 9 1 14 13 0 2 4 11 9 13 9 1 14 13 15 15 4 13 15 2
6 4 10 9 13 3 2
12 9 13 1 1 9 1 16 11 9 13 0 2
24 11 13 3 12 9 2 13 0 9 7 13 3 1 9 1 0 9 2 16 9 13 1 11 2
14 13 15 15 15 13 16 9 4 13 9 1 11 9 2
8 15 13 0 15 4 13 0 2
4 9 1 11 5
25 2 6 2 15 13 9 4 13 9 16 15 13 3 16 10 0 13 9 1 11 16 9 13 0 2
13 15 13 3 0 16 10 9 1 11 9 13 3 2
34 9 4 13 15 1 16 15 13 0 9 1 10 9 1 16 15 13 0 9 1 11 16 9 13 1 2 3 4 15 13 1 1 15 2
6 10 0 9 1 9 2
17 0 13 1 0 9 1 9 15 13 11 9 2 15 13 0 9 2
14 9 13 11 9 2 15 3 13 9 1 9 7 9 2
15 9 13 16 10 12 9 13 3 1 10 9 15 13 15 2
15 15 13 16 9 9 13 0 1 1 9 1 9 1 11 2
6 9 13 9 1 0 2
11 10 9 13 9 1 9 3 9 13 1 2
17 9 13 3 1 1 9 2 7 13 14 13 1 0 9 1 9 2
9 2 15 13 0 9 1 9 9 2
15 9 13 9 1 14 13 1 1 9 2 1 9 1 9 2
21 1 10 9 13 9 10 0 0 9 1 14 13 9 2 13 9 1 9 1 11 2
11 2 15 4 15 13 16 9 4 13 1 2
20 2 9 1 0 9 15 13 3 1 10 0 9 2 4 13 1 9 1 9 2
16 16 3 10 9 4 4 13 9 2 4 9 4 13 1 9 2
8 2 15 13 15 1 11 9 2
11 2 16 9 0 0 4 13 1 1 9 2
32 15 13 0 0 16 15 3 4 13 10 9 15 13 9 1 2 7 15 13 0 16 15 4 13 15 3 0 1 1 1 15 2
15 15 13 15 4 13 9 1 14 13 15 15 4 13 1 2
5 15 13 11 9 2
17 0 1 9 13 15 10 12 15 13 9 1 15 15 13 3 1 2
12 2 15 13 0 15 4 13 0 2 13 9 2
15 15 13 16 11 9 2 10 0 9 2 13 10 0 9 2
23 2 15 13 3 15 16 15 13 2 7 10 0 12 9 15 13 13 15 15 0 7 0 2
14 15 13 0 2 13 0 7 13 1 10 0 1 9 2
10 15 13 15 13 9 15 13 1 9 2
18 2 13 15 0 1 14 13 9 1 12 9 16 15 13 0 1 9 2
27 2 15 13 1 10 9 1 14 13 3 9 13 15 2 7 13 15 4 13 1 9 10 16 15 13 0 2
11 15 13 0 1 9 16 15 13 1 9 2
29 2 15 13 15 12 9 1 9 2 3 13 15 7 13 15 16 15 3 13 14 13 1 15 15 13 0 1 9 2
13 2 13 15 15 1 14 13 10 9 1 1 9 2
25 2 6 2 16 9 1 15 13 0 7 0 2 7 1 9 13 15 3 0 3 2 3 13 2 2
27 2 11 13 0 15 4 13 14 13 1 16 9 13 1 9 1 9 2 7 13 15 4 13 1 0 9 2
6 13 15 3 0 9 2
10 2 6 2 13 1 9 13 15 15 2
11 15 13 0 16 9 13 1 9 1 9 2
21 9 1 9 7 9 4 1 0 9 13 0 2 7 4 1 10 0 9 13 0 2
20 9 13 0 1 15 2 7 13 3 16 9 4 13 10 0 9 1 9 10 2
7 7 9 10 13 0 3 2
27 7 3 1 9 1 15 15 0 13 1 9 15 13 1 1 9 1 9 2 13 15 0 1 11 7 9 2
22 2 15 13 10 0 9 15 4 13 2 15 4 13 15 1 15 1 15 2 13 9 2
25 2 15 13 9 1 15 16 9 10 7 15 13 3 0 7 0 2 3 4 15 0 4 13 1 2
12 15 13 3 15 15 13 1 15 2 13 11 2
7 9 13 15 0 0 9 2
13 15 13 0 0 1 16 10 10 13 15 1 15 2
10 16 15 13 14 13 9 1 14 13 2
7 3 15 4 13 9 9 2
14 2 0 1 15 13 0 7 0 1 3 15 13 15 2
13 4 10 1 15 13 2 4 9 10 13 0 0 2
17 15 13 0 0 1 16 15 4 13 0 14 13 15 15 13 1 2
17 2 7 16 15 13 1 9 15 3 13 15 0 2 3 13 1 2
21 9 1 0 9 13 15 1 1 9 15 13 1 9 1 0 9 16 15 13 15 2
15 15 13 3 0 14 13 10 9 3 0 1 15 3 0 2
2 3 2
21 1 9 13 9 9 7 0 0 1 16 9 10 3 4 4 13 15 15 10 13 2
23 11 13 1 10 9 1 12 9 10 10 9 1 9 2 7 13 9 1 9 1 0 9 2
32 0 13 15 1 11 12 2 7 13 1 1 14 13 2 11 9 2 2 10 9 1 9 1 9 15 13 1 9 7 0 9 2
12 9 1 9 13 15 1 9 1 14 13 1 2
19 9 1 9 13 15 0 0 1 2 7 11 13 14 13 15 13 9 10 2
8 2 15 13 10 9 15 13 2
15 15 13 14 13 15 0 2 3 16 10 9 4 13 10 2
79 9 4 0 1 9 1 11 11 11 2 11 9 2 11 9 2 11 9 2 0 9 11 11 11 1 11 9 2 0 9 11 11 1 11 9 2 0 9 11 11 1 11 9 2 9 11 11 1 11 9 2 11 9 11 11 11 2 11 9 9 7 9 11 11 11 2 0 9 2 9 11 11 1 11 1 11 7 9 2
12 2 16 9 13 2 13 15 3 0 14 13 5
6 2 4 9 0 13 2
5 0 9 7 9 5
3 13 9 5
9 2 15 13 11 1 14 13 9 2
7 2 15 13 1 12 9 5
10 2 15 13 12 9 16 9 4 13 5
9 2 13 15 3 9 1 0 9 2
5 2 15 13 9 5
4 9 13 0 5
2 11 2
3 13 9 5
5 15 13 9 1 5
5 15 13 15 1 5
6 15 13 15 9 1 5
3 12 9 5
21 1 9 4 9 7 9 13 1 11 1 14 13 0 9 0 9 1 9 1 9 2
2 9 2
23 11 9 11 11 2 9 11 11 7 0 9 11 11 1 9 9 1 11 1 9 0 9 2
4 9 2 11 5
45 1 9 13 3 9 1 11 9 2 9 2 2 11 11 2 0 9 11 11 7 9 11 11 1 10 0 9 1 11 1 14 13 1 9 0 1 9 1 11 7 1 9 0 9 2
36 15 4 13 1 14 13 16 0 9 13 10 9 1 0 9 15 4 13 1 11 1 0 9 11 11 7 0 9 11 11 1 9 2 13 11 2
2 12 2
11 11 11 2 11 2 13 0 9 1 9 2
11 2 9 13 0 1 9 1 9 1 9 2
7 15 13 1 10 0 9 2
12 4 15 0 13 2 7 4 15 13 1 9 2
5 9 11 11 13 2
28 2 15 13 9 15 3 4 13 1 9 2 7 15 13 9 15 3 7 0 13 1 1 9 2 1 0 9 2
30 7 9 7 9 4 13 1 9 1 9 15 3 13 1 0 9 2 7 3 15 4 13 0 14 13 9 1 11 11 2
14 3 15 4 13 2 4 15 4 4 13 1 1 1 2
14 16 9 13 1 9 1 9 2 13 15 0 1 15 2
12 15 13 1 9 1 10 0 9 2 13 11 2
2 12 2
13 11 11 2 11 2 13 1 9 1 9 7 11 2
12 2 15 13 1 10 0 9 1 9 7 11 2
21 4 9 13 16 0 9 4 13 16 15 4 13 0 9 1 9 10 12 9 13 2
3 11 13 2
17 2 15 13 0 0 9 1 16 15 4 13 9 1 9 1 11 2
17 15 13 0 9 1 9 15 13 0 2 9 1 9 2 7 9 2
22 2 16 15 4 13 1 0 9 7 9 2 15 4 15 13 2 13 11 11 11 11 2
16 2 15 13 3 2 7 15 13 7 9 7 9 2 13 11 2
2 12 2
15 11 11 2 11 2 13 1 9 1 9 2 9 7 11 2
12 2 15 13 1 9 1 9 2 9 7 9 2
13 13 9 15 13 0 1 9 1 9 2 13 11 2
14 2 0 13 15 15 13 10 0 9 1 9 7 1 2
30 7 15 4 13 15 16 15 13 0 1 0 9 15 13 1 9 2 1 10 9 2 16 15 13 0 3 2 13 11 2
5 9 11 11 13 2
17 2 15 13 0 9 2 16 9 4 13 1 10 10 9 1 12 2
7 15 13 0 9 7 9 2
17 2 3 0 13 11 1 9 1 14 4 13 10 9 2 13 11 5
17 2 15 4 13 0 1 15 1 14 4 13 9 2 13 11 11 2
2 12 2
13 11 11 2 11 2 13 9 1 11 9 1 9 2
14 2 15 13 11 0 9 1 14 13 9 2 13 11 2
29 2 15 4 13 1 10 9 1 11 1 3 15 4 13 0 7 0 13 9 1 14 4 13 10 9 9 1 9 2
19 1 9 9 4 15 13 10 9 2 15 4 4 13 1 1 9 1 9 2
18 15 13 0 9 15 15 4 13 10 0 9 1 2 13 9 11 11 2
18 2 15 4 0 13 16 9 4 13 0 9 2 13 11 11 11 11 2
20 2 10 9 13 3 9 1 15 15 13 2 7 4 13 9 0 0 7 13 2
14 15 13 9 16 10 0 9 4 13 0 1 11 9 2
11 15 4 3 13 9 2 13 9 11 11 2
7 2 16 15 13 1 9 2
16 4 15 13 1 16 9 9 13 15 13 0 2 13 11 11 2
11 2 15 4 13 10 0 9 2 13 11 2
2 12 2
10 11 11 2 11 2 13 1 11 9 2
12 2 3 0 9 1 11 13 15 2 13 11 2
14 2 15 13 12 9 0 2 7 12 9 1 10 9 2
12 15 13 3 10 9 1 11 2 13 9 11 2
14 2 11 13 10 9 1 9 15 13 0 1 1 11 2
12 4 15 3 13 10 9 1 11 2 13 11 2
25 2 15 4 0 9 13 9 1 15 15 13 1 2 15 4 3 13 10 0 1 10 9 15 13 2
18 15 13 9 1 12 9 2 7 15 13 0 1 9 2 13 11 11 2
2 12 2
9 11 11 2 11 2 13 1 9 2
29 2 15 13 15 1 9 1 9 1 9 7 11 15 13 1 16 15 13 12 9 7 12 9 15 16 15 13 9 2
22 2 10 0 9 13 9 1 13 9 1 9 2 7 15 13 9 1 9 1 10 9 2
26 15 13 10 9 15 4 13 1 9 2 16 15 4 13 9 1 9 1 11 0 2 13 9 11 11 2
17 2 13 15 10 0 9 1 9 1 14 13 1 9 2 13 11 2
21 2 0 13 15 3 15 2 15 13 9 1 9 7 13 1 10 0 9 1 9 2
8 15 13 10 9 15 4 13 2
16 15 4 3 13 16 9 13 3 0 1 10 9 2 13 11 2
10 2 15 13 12 9 16 9 4 13 2
19 13 15 0 16 15 1 10 9 4 4 13 1 9 1 9 1 10 9 2
21 2 15 4 4 13 9 0 2 7 15 13 10 9 1 10 10 9 2 13 11 2
2 12 2
11 11 11 2 11 2 13 9 1 0 9 5
16 2 11 13 1 1 10 9 16 15 13 9 15 13 0 9 2
13 15 4 13 14 13 0 1 16 15 4 13 15 2
6 11 4 3 13 3 2
11 10 0 9 4 13 9 0 7 13 9 2
16 13 15 10 9 16 15 13 3 9 1 15 1 10 0 9 2
5 9 11 11 13 2
14 2 15 13 12 9 1 0 9 2 12 1 10 9 2
9 15 13 1 10 0 9 0 9 2
20 15 13 0 1 15 14 13 9 7 9 1 2 7 15 13 0 16 15 13 2
15 15 15 13 10 9 13 16 15 13 0 7 16 15 13 2
20 16 15 1 9 13 1 9 2 7 13 1 9 7 13 0 9 2 13 11 2
12 2 10 0 9 1 10 0 9 13 0 9 2
26 1 9 13 15 16 10 9 15 13 1 9 2 13 16 15 13 0 9 1 15 2 13 9 11 11 2
16 2 4 9 13 15 1 3 15 13 1 9 1 9 1 9 2
39 2 4 13 0 9 1 14 13 15 2 7 15 13 10 0 7 0 9 15 15 13 1 1 14 13 1 2 7 15 13 3 1 9 16 15 13 0 9 2
18 15 13 1 14 13 1 11 7 9 1 13 9 2 13 9 11 11 2
2 12 2
11 11 11 11 2 11 2 13 9 1 11 2
15 2 13 15 0 1 16 15 13 0 9 1 11 7 9 2
4 9 11 13 2
17 2 6 2 15 13 0 1 15 3 15 4 13 1 9 1 9 2
16 15 4 3 13 16 15 4 13 1 14 13 0 1 16 9 2
11 2 15 4 13 9 7 9 2 13 9 2
18 13 3 9 10 0 9 1 16 15 3 13 0 3 9 2 13 11 2
15 2 10 9 13 16 15 4 13 1 9 1 14 13 0 2
27 1 0 9 7 9 13 15 1 9 1 9 2 7 3 15 4 13 16 15 13 1 0 9 2 13 11 2
18 2 4 15 13 0 14 13 9 7 9 1 10 0 9 2 13 11 2
11 2 15 13 3 0 14 13 15 7 13 2
23 10 9 13 14 13 10 9 15 13 2 15 4 13 7 15 4 13 1 3 2 13 9 2
2 12 2
6 0 9 11 11 13 2
16 2 15 13 16 7 9 0 9 7 9 4 13 9 1 9 2
16 2 15 4 13 10 9 2 13 11 13 2 1 9 1 9 2
18 9 15 4 13 1 9 0 9 3 13 1 9 2 3 1 0 9 2
11 9 4 13 1 10 0 15 13 1 9 5
7 2 9 4 13 1 11 2
19 10 0 9 4 13 1 3 16 15 4 13 10 9 1 10 9 13 9 2
11 9 1 9 13 16 15 13 9 1 9 2
8 15 4 3 3 13 1 9 2
19 0 9 4 3 13 2 7 9 4 4 13 1 9 1 15 2 13 9 2
17 2 9 4 1 10 9 13 1 1 9 1 9 7 9 7 9 2
14 2 15 13 0 0 1 9 2 15 15 13 0 9 2
25 15 4 13 10 9 1 11 2 15 13 3 7 13 10 9 1 9 2 9 7 9 2 13 11 2
2 12 2
7 9 11 11 13 10 9 2
17 2 16 15 4 4 13 15 0 2 13 15 0 9 1 9 9 2
8 2 9 15 13 15 1 11 5
2 9 5
4 0 1 15 5
4 13 1 9 5
3 11 9 5
4 13 1 9 5
2 0 5
4 13 1 9 5
2 11 5
2 9 5
3 13 9 5
4 10 0 9 5
5 2 9 0 9 5
6 2 15 13 9 10 5
2 9 5
8 1 1 11 13 10 0 9 2
6 9 4 13 1 9 2
19 10 9 13 11 11 2 12 2 13 1 9 1 9 2 12 9 1 9 2
7 9 1 9 0 9 12 2
14 9 4 3 13 15 2 1 15 15 13 10 9 13 2
25 9 13 9 1 9 1 11 11 11 1 11 9 2 7 13 10 9 13 1 9 1 9 0 9 2
5 9 13 11 11 2
11 15 13 15 1 10 9 7 9 1 9 2
7 15 13 1 14 13 1 2
12 1 0 9 13 15 3 12 9 1 1 9 2
13 3 1 16 11 13 1 9 2 13 9 15 13 2
7 10 9 0 2 9 9 2
26 11 11 13 1 1 11 1 10 9 2 15 13 1 9 1 9 1 14 13 10 9 15 13 12 9 2
19 9 11 13 1 7 13 0 1 9 2 16 15 3 4 13 7 13 9 2
9 13 15 15 15 4 13 1 11 2
5 15 13 1 9 5
9 11 13 10 9 1 10 0 9 2
9 1 0 9 13 15 9 7 9 2
7 9 13 9 7 9 9 2
11 15 4 13 1 11 11 7 13 1 9 2
12 11 9 13 14 13 9 2 7 13 10 9 2
13 1 0 9 13 15 0 1 9 1 11 0 9 2
8 1 10 9 4 15 13 9 2
18 1 1 0 9 1 10 9 13 9 1 10 9 2 9 10 0 9 2
5 1 10 9 1 2
9 1 9 13 11 1 9 1 9 2
11 15 7 9 11 11 11 13 1 10 9 2
7 15 13 10 9 15 13 2
30 11 13 16 11 13 0 2 7 13 16 15 3 4 13 1 1 15 7 13 10 9 2 1 9 1 14 13 1 9 2
12 7 11 13 3 15 2 7 9 13 3 9 2
11 11 13 1 15 9 7 13 9 1 9 2
11 15 13 0 0 2 7 15 13 0 1 2
36 11 7 11 4 13 1 1 10 9 2 15 4 13 15 16 15 13 1 9 7 13 1 3 0 9 15 13 2 7 16 15 13 0 1 15 2
19 1 9 4 9 13 1 10 9 16 11 3 13 0 3 1 14 13 1 2
13 15 13 0 3 3 0 1 14 13 1 10 9 2
15 11 13 15 1 1 10 9 1 11 2 13 9 1 15 2
6 10 0 9 13 1 2
8 11 13 3 10 9 1 15 2
16 15 13 1 11 2 16 11 13 9 1 14 13 10 10 9 2
18 7 11 13 3 1 1 11 2 0 13 15 3 1 3 2 13 15 2
13 11 13 15 4 13 1 2 7 11 13 15 3 2
14 15 4 13 15 0 2 3 16 3 15 4 13 1 2
13 11 13 9 1 9 10 2 15 15 13 1 9 2
6 15 4 13 9 3 2
25 2 0 2 15 13 1 2 7 15 13 1 3 1 12 2 12 9 7 13 1 15 2 13 11 2
20 4 15 13 2 13 15 1 16 15 4 13 10 9 15 13 14 13 1 9 2
11 2 16 3 2 13 15 1 2 13 15 2
5 0 1 1 11 2
7 9 11 13 0 1 9 2
21 15 13 10 9 1 16 15 4 13 1 9 1 9 2 7 13 15 0 1 15 2
5 13 9 1 9 5
7 13 15 0 0 1 9 2
3 0 9 2
22 9 11 11 4 13 9 1 0 9 15 13 10 9 1 9 15 13 9 1 9 10 2
2 9 2
18 16 9 1 10 9 13 9 1 16 15 3 13 0 9 2 13 0 2
2 0 2
16 3 10 9 1 0 9 1 9 1 9 2 13 1 0 9 2
5 13 10 0 9 2
14 9 4 3 13 1 14 13 10 9 9 0 0 0 2
19 3 4 9 1 9 1 1 9 1 9 0 13 13 0 9 14 13 1 2
35 9 1 2 4 15 13 9 1 1 9 16 15 13 15 1 9 2 2 4 13 0 1 9 1 9 2 1 1 3 3 0 1 0 9 2
32 3 4 9 11 11 13 1 10 9 15 4 13 1 10 0 0 9 1 9 1 10 3 0 9 10 9 13 1 1 10 9 2
46 11 13 9 2 11 11 2 2 7 13 16 15 13 14 13 9 10 9 7 10 9 1 14 13 0 0 1 15 1 9 1 15 15 13 1 1 14 13 1 9 1 9 10 1 9 2
15 9 13 9 1 0 9 16 10 9 4 13 1 1 9 2
39 2 15 14 13 3 2 2 2 13 10 10 9 2 7 2 9 1 16 15 13 15 2 13 1 9 15 1 9 4 13 1 0 7 0 0 9 1 9 2
19 9 13 0 2 15 13 3 14 13 9 1 9 16 15 13 15 1 9 2
33 16 9 13 9 1 9 10 2 13 0 7 0 9 1 0 9 2 7 9 13 3 10 10 9 1 9 9 13 1 1 9 10 2
23 3 4 9 15 13 9 1 9 13 1 10 9 1 9 7 9 2 3 16 9 13 1 2
24 9 13 1 0 9 9 1 14 13 1 1 9 1 9 7 13 9 1 9 1 9 7 9 2
11 16 9 10 9 13 1 9 2 13 3 2
21 7 1 0 9 1 11 1 9 4 15 13 15 13 14 13 10 9 1 0 9 2
16 7 3 13 15 3 14 13 1 16 15 13 10 9 1 9 2
14 10 9 4 13 1 11 9 2 7 3 13 1 9 2
13 13 15 9 7 9 2 13 15 1 15 1 9 2
3 10 0 5
16 9 11 11 2 12 2 13 15 4 13 9 1 9 1 9 2
3 1 12 2
12 9 11 1 0 9 1 9 1 11 1 11 2
5 9 15 13 12 2
8 11 11 7 11 11 1 9 2
3 1 12 2
4 16 15 13 2
19 11 2 3 2 1 9 1 11 1 9 11 11 1 9 1 11 1 12 2
2 0 2
13 11 11 1 9 1 15 15 13 3 0 0 1 2
9 11 11 2 11 11 7 9 11 2
18 15 13 0 9 12 7 9 4 3 13 0 10 10 3 1 11 11 2
23 15 13 12 9 2 9 1 11 2 7 10 1 10 0 1 9 15 4 13 1 10 9 2
14 1 9 1 9 13 15 1 9 2 15 13 0 9 2
8 2 4 15 13 0 1 11 2
8 15 4 13 10 9 1 11 2
6 0 11 11 13 9 2
25 15 13 0 7 0 2 15 13 9 15 13 9 1 2 13 9 1 9 1 11 7 9 1 11 2
9 3 10 9 1 16 9 13 1 2
19 15 13 3 14 13 15 0 9 2 7 13 11 13 0 9 7 0 9 2
9 15 13 10 0 9 15 13 15 2
7 9 11 4 13 1 9 2
13 12 12 9 4 13 2 3 10 9 13 1 9 2
17 9 13 0 2 15 13 3 9 1 0 9 2 15 13 9 12 2
13 15 13 1 9 15 13 1 2 15 13 1 9 2
12 1 9 1 12 9 13 15 0 9 1 9 2
13 1 1 11 13 15 10 0 9 16 9 0 13 2
22 15 13 3 15 13 2 9 15 13 16 15 12 9 0 4 13 10 9 11 4 13 2
8 11 11 4 13 0 1 9 2
13 10 9 13 15 9 11 1 1 9 2 11 2 2
22 1 9 13 9 9 1 9 1 11 2 16 9 7 10 12 9 13 1 9 1 11 2
12 2 15 4 13 1 2 7 3 4 9 13 2
15 3 10 9 4 15 13 1 9 1 14 13 1 15 3 2
22 11 11 13 1 1 10 0 9 16 15 13 7 13 0 1 9 10 1 11 1 11 2
29 1 10 12 9 13 15 0 1 0 2 15 13 3 3 0 1 9 1 15 15 10 9 13 9 1 9 11 11 2
13 10 0 0 9 1 12 4 13 1 9 11 11 2
19 9 4 13 1 9 2 7 0 3 1 13 11 9 2 9 11 11 11 2
12 10 9 1 12 13 11 11 2 9 1 11 2
25 16 15 13 1 9 2 13 15 3 10 0 9 1 10 0 9 13 15 1 1 9 16 9 13 2
11 9 13 3 14 13 9 10 3 1 9 2
23 15 13 3 1 15 15 1 9 15 3 13 14 13 9 1 2 7 15 13 15 0 0 2
12 0 1 2 11 2 13 9 1 10 0 9 2
16 9 13 1 0 9 1 9 2 9 2 9 2 9 7 9 2
20 2 3 13 15 9 1 15 15 13 16 10 0 9 13 1 14 4 13 9 2
5 2 15 13 15 2
13 2 15 13 1 0 9 16 9 4 13 1 15 2
20 7 15 13 15 3 0 0 2 15 13 15 10 9 1 14 4 13 3 0 2
18 10 9 4 15 13 1 0 9 2 7 15 13 0 0 1 10 9 2
16 2 13 15 10 14 13 16 15 13 1 10 9 15 4 13 2
16 2 9 13 3 1 9 15 13 1 2 7 1 15 15 13 2
14 1 14 13 15 0 15 15 3 4 13 2 7 13 2
22 3 1 1 10 10 9 2 2 11 2 11 2 2 4 3 10 9 13 1 0 9 2
24 2 15 13 3 0 2 7 13 0 9 1 14 13 11 2 15 13 10 0 9 1 0 9 2
8 9 13 1 10 9 1 9 2
11 2 15 4 13 16 15 3 13 1 9 2
9 2 15 13 3 1 9 1 9 2
14 9 13 9 1 10 9 15 13 1 1 14 13 0 2
18 1 15 13 15 14 13 1 10 9 3 0 0 16 15 4 13 0 2
12 15 13 3 14 13 2 7 15 4 15 13 2
5 2 15 13 15 2
4 2 10 9 2
15 10 1 10 0 1 11 13 3 1 14 4 13 12 9 2
18 15 13 15 16 1 10 0 9 2 4 15 13 7 13 1 10 0 2
8 10 9 15 13 0 10 9 2
23 3 13 15 3 3 7 4 13 16 10 10 9 4 4 13 1 16 15 13 1 0 9 2
27 2 11 2 11 2 4 13 1 12 12 9 1 9 1 12 2 7 13 10 0 0 9 1 9 10 9 2
13 15 13 12 9 2 11 7 13 11 9 1 11 2
17 15 13 3 10 9 1 11 2 16 15 4 13 1 0 0 9 2
3 1 10 2
11 7 9 15 13 15 4 13 10 0 9 2
12 2 15 13 10 9 15 13 9 14 13 3 2
13 14 13 15 15 3 4 13 0 4 15 3 13 2
17 15 4 13 9 15 7 13 2 7 15 13 14 13 15 1 9 2
11 2 15 13 3 0 1 14 13 0 9 2
5 2 6 2 6 2
3 2 6 2
6 2 6 2 10 9 2
10 15 13 16 15 4 13 0 3 0 2
17 16 15 3 13 15 15 13 1 15 9 1 14 13 10 0 9 2
14 2 16 10 9 13 15 0 2 4 15 3 13 9 2
7 2 6 2 15 13 3 2
2 3 2
15 7 10 9 13 15 3 16 2 3 13 15 0 0 2 2
7 2 13 9 15 1 15 2
10 2 15 13 1 9 15 4 13 15 2
16 3 13 15 1 1 15 2 10 15 15 3 3 13 1 15 2
4 2 15 3 2
4 2 10 9 2
6 7 15 4 13 15 2
18 9 1 9 7 1 14 13 10 9 1 14 13 10 9 2 13 0 2
13 7 16 15 3 13 1 9 2 2 0 15 13 2
6 2 7 13 15 0 2
18 11 11 4 13 1 15 9 2 13 15 1 9 2 7 13 1 9 2
16 15 13 9 1 9 11 11 2 13 9 1 0 9 7 13 2
4 2 6 3 2
9 15 4 13 15 10 1 0 0 2
12 2 4 15 14 13 13 10 9 1 0 9 2
7 2 9 1 9 2 6 2
8 15 4 3 13 9 1 15 2
16 15 13 11 11 15 1 9 13 15 0 0 14 13 0 9 2
19 15 13 9 2 9 1 9 2 2 7 13 9 2 0 2 0 9 2 2
16 2 15 13 11 0 2 7 15 13 1 10 9 10 0 9 2
21 15 13 10 9 2 7 13 0 0 0 16 15 13 14 13 15 10 1 1 9 2
11 2 13 15 2 0 2 0 9 2 9 2
9 2 6 2 15 13 3 3 15 2
15 7 15 4 13 10 9 16 3 3 10 9 4 4 13 2
22 3 13 15 3 16 15 15 13 2 0 2 0 2 9 2 13 7 13 2 11 2 2
8 2 4 3 15 0 0 13 2
9 2 6 2 15 13 3 0 9 2
13 15 13 1 10 9 1 1 15 15 13 10 9 2
15 1 9 1 9 13 15 9 1 10 9 15 13 1 9 2
15 15 13 10 9 1 9 2 11 2 13 1 9 11 11 2
5 2 15 13 9 2
6 10 0 2 0 9 2
24 15 13 10 9 2 13 11 2 15 1 9 4 13 14 13 9 15 13 3 1 9 13 1 2
14 11 11 11 13 3 16 2 11 2 11 2 13 0 2
8 9 1 9 13 0 3 0 2
10 11 13 3 12 9 16 9 13 15 2
10 15 13 0 1 9 2 9 1 9 2
24 1 0 9 13 9 9 0 9 1 9 2 7 9 1 9 2 11 2 7 2 11 11 2 2
12 15 13 9 1 9 2 11 7 10 0 9 2
14 3 1 12 4 15 1 11 13 1 2 11 11 2 2
18 15 13 9 16 15 13 1 10 0 9 1 0 9 1 9 1 12 2
17 2 1 9 13 15 0 0 0 2 7 13 3 1 9 1 9 2
17 15 13 10 9 15 13 0 0 9 2 7 13 3 10 0 9 2
16 1 10 9 13 15 0 2 13 0 9 7 13 3 1 12 2
13 1 10 9 4 10 9 4 13 1 1 10 9 2
13 9 13 11 11 2 15 13 10 0 9 1 11 2
35 11 11 11 4 13 1 11 0 9 2 4 13 9 11 11 2 13 9 1 11 2 7 13 15 1 16 0 9 4 4 13 15 1 9 2
7 2 15 13 15 1 15 2
11 2 16 15 4 13 15 15 13 9 1 2
17 7 16 15 14 13 10 0 1 10 2 13 14 13 10 0 3 2
14 11 11 13 12 9 7 4 13 15 1 1 14 13 2
7 15 13 1 1 9 12 2
7 15 13 9 15 13 15 2
19 9 1 11 4 13 15 10 0 9 2 7 15 13 1 9 1 11 9 2
10 10 9 13 15 1 9 1 12 9 2
6 15 13 3 9 13 2
10 13 15 15 15 4 13 9 1 9 2
4 13 15 9 2
7 6 2 15 13 3 15 2
23 16 15 1 0 9 13 11 11 1 11 1 11 9 1 11 2 4 15 4 13 1 9 2
15 15 13 0 9 1 11 2 7 13 0 0 1 14 13 2
13 15 4 13 10 10 9 2 3 13 9 1 10 2
14 12 9 1 13 15 1 1 11 11 1 11 1 9 2
8 9 13 1 12 9 12 9 2
11 1 10 9 4 15 13 10 9 1 11 2
14 15 13 10 9 0 1 10 10 9 1 9 7 9 2
12 9 15 3 4 13 1 0 13 1 0 9 2
13 2 15 4 13 3 0 9 2 15 13 1 9 2
21 15 13 0 0 1 15 14 13 10 9 2 14 13 15 15 0 4 13 1 1 2
7 1 11 4 15 13 0 2
19 1 10 9 13 15 1 9 2 15 15 4 13 16 15 13 9 1 9 2
14 9 13 3 3 0 2 7 15 13 0 0 1 15 2
11 10 13 15 1 10 9 2 15 13 9 2
20 15 13 3 3 3 1 9 1 10 9 2 7 15 13 10 0 9 1 9 2
5 2 1 15 3 2
19 2 15 4 13 1 1 10 9 15 10 9 1 11 7 11 4 13 1 2
17 15 14 13 3 1 2 13 0 1 2 13 10 0 7 0 9 2
16 1 0 9 13 15 1 10 0 7 0 9 15 13 1 9 2
11 2 7 3 13 15 3 3 9 1 9 2
25 2 15 13 15 15 4 13 1 9 16 9 13 1 0 1 15 2 3 13 9 1 9 7 9 2
7 15 13 15 13 0 0 2
10 11 1 11 13 12 0 9 1 11 2
11 15 13 1 9 2 7 13 14 13 9 2
11 1 12 13 15 1 9 1 2 11 2 2
23 1 12 9 4 15 13 12 9 2 7 10 9 9 1 15 1 11 9 1 11 11 11 2
19 0 2 1 10 0 9 2 4 13 3 0 0 9 2 0 1 0 9 2
12 15 13 3 7 7 1 9 10 2 0 7 2
29 3 0 4 15 13 15 1 1 12 9 1 10 2 11 2 2 10 9 15 4 13 15 1 10 9 1 0 9 2
13 2 16 10 0 9 13 0 2 13 3 3 9 2
10 15 13 3 3 10 9 1 0 15 2
13 16 10 0 9 13 3 0 4 13 0 1 0 2
25 3 13 15 3 3 2 7 15 13 3 3 16 15 13 9 1 0 15 4 13 1 1 15 3 2
14 16 15 13 0 1 1 9 2 13 15 1 10 9 2
13 15 13 10 9 2 16 9 4 13 15 1 9 2
33 10 0 13 10 0 9 15 13 16 15 13 1 0 9 2 7 15 13 0 1 16 15 13 10 0 9 2 3 0 2 3 0 2
10 2 3 0 9 4 15 13 1 11 2
17 2 15 4 13 9 1 12 0 9 2 7 1 12 7 12 9 2
7 2 3 4 15 13 9 2
8 13 3 11 9 1 10 9 2
26 2 1 14 4 13 12 7 12 9 1 9 1 12 2 13 15 0 10 9 7 9 15 4 13 1 2
13 15 13 3 15 15 4 13 1 1 7 1 9 2
23 3 4 15 13 1 11 11 11 2 15 13 10 9 15 13 3 0 9 1 14 13 1 2
35 7 1 10 9 4 15 13 0 1 14 13 1 10 15 1 14 13 10 2 9 1 13 2 2 7 3 10 0 9 1 10 0 0 9 2
19 15 13 0 9 13 1 9 16 15 13 1 3 1 11 2 11 7 11 2
8 7 15 13 15 3 2 3 2
23 3 13 15 1 9 0 9 3 1 1 11 2 7 4 13 0 1 1 11 1 12 9 2
12 2 15 13 1 1 16 15 13 9 1 11 2
16 2 15 4 13 9 1 10 9 1 9 1 9 1 0 9 2
13 16 15 3 13 2 4 15 13 0 14 13 9 2
11 15 13 10 3 0 9 1 15 3 1 2
7 15 15 13 2 15 13 2
22 16 15 13 1 9 1 9 2 4 15 13 1 1 11 1 10 0 9 1 9 10 2
24 15 4 13 0 9 2 15 4 13 9 2 9 7 9 2 7 1 1 0 9 13 9 11 2
7 15 13 10 9 14 13 2
8 2 13 15 0 2 13 15 2
9 2 15 13 3 0 2 13 11 2
7 2 6 2 15 13 15 2
11 11 13 0 2 13 9 2 13 7 13 2
7 15 13 1 9 1 11 2
23 15 13 15 15 1 9 4 13 1 15 16 2 9 13 0 2 7 11 13 15 0 2 2
19 9 15 13 9 10 1 2 13 10 11 11 1 14 13 1 10 0 9 2
10 2 11 13 10 0 9 15 13 1 2
16 15 13 10 9 1 9 2 7 10 0 9 1 15 1 15 2
22 0 9 1 9 13 15 10 0 9 10 9 4 13 1 15 10 2 13 15 1 9 2
22 1 9 13 15 16 11 13 0 0 1 9 2 10 9 7 9 15 13 14 13 9 2
16 16 15 13 1 7 13 2 13 15 10 0 0 9 1 15 2
7 13 9 16 15 13 1 2
12 13 1 10 9 7 9 15 13 1 9 10 2
12 7 15 13 11 16 15 4 13 15 10 0 2
18 3 13 15 3 1 10 9 2 13 15 7 15 10 10 0 9 9 2
4 7 13 0 2
8 1 10 9 10 3 0 9 2
7 2 13 15 0 3 0 2
7 2 6 2 13 15 15 2
7 15 4 3 15 13 1 2
10 11 13 1 10 0 9 10 1 9 2
5 4 15 13 0 2
7 6 2 15 13 0 0 2
23 2 15 4 3 13 15 3 16 15 13 9 1 9 3 1 2 7 15 13 14 13 15 2
12 15 13 3 3 0 0 1 9 7 9 10 2
8 10 12 13 1 9 1 12 2
16 15 13 9 1 10 0 9 2 11 2 2 16 11 13 9 2
13 15 13 1 15 2 7 10 9 13 15 1 15 2
18 1 12 0 9 2 13 15 1 11 11 1 14 13 10 9 1 9 2
10 1 10 9 9 13 15 9 1 11 2
4 15 13 11 2
19 2 15 13 15 4 13 2 15 4 3 13 9 7 13 15 0 1 9 2
16 12 9 1 13 15 3 2 0 1 9 7 13 15 1 9 2
14 15 13 10 0 9 1 15 2 7 0 0 1 15 2
14 15 13 0 0 16 15 13 14 13 1 10 0 9 2
6 9 1 13 1 11 2
21 1 9 1 11 13 15 1 1 9 2 15 13 0 2 9 1 15 13 14 13 2
22 15 4 13 12 9 16 15 13 1 9 16 11 13 1 1 9 12 12 9 1 9 2
3 15 13 2
11 2 15 13 1 10 9 1 14 13 9 2
5 15 13 3 0 2
15 16 15 13 1 11 4 15 1 7 1 13 9 1 9 2
14 10 0 15 13 16 15 13 1 2 13 14 13 9 2
15 2 15 13 0 0 2 11 2 13 9 7 13 10 9 2
14 2 7 13 15 9 14 13 15 15 4 13 15 1 2
12 0 9 12 13 15 9 1 10 9 1 11 2
7 12 9 12 9 1 9 2
20 7 16 11 11 13 1 9 1 2 11 2 11 2 2 13 9 0 10 9 2
11 2 0 13 15 3 9 7 9 1 15 2
22 15 13 0 0 1 2 15 13 10 9 0 9 2 7 13 3 0 1 9 1 15 2
14 15 4 10 9 13 2 15 4 3 13 14 13 9 2
18 15 13 10 0 9 2 16 15 13 1 10 10 9 7 3 4 13 2
5 2 15 13 0 2
4 2 0 9 2
7 11 13 0 7 4 13 2
4 9 10 13 2
17 15 13 1 10 9 15 13 1 15 15 0 4 13 1 10 9 2
11 15 4 13 15 2 7 15 4 13 15 2
8 15 13 1 10 3 0 9 2
16 15 13 3 0 14 13 1 2 1 14 4 13 0 1 9 2
21 16 15 13 0 9 1 15 3 2 3 13 15 16 15 13 14 13 9 1 15 2
20 15 13 3 0 14 13 13 2 7 15 13 0 14 13 15 14 13 0 0 2
39 2 15 13 15 15 13 4 13 1 1 9 3 1 15 3 3 2 13 11 11 16 15 13 9 1 9 1 2 11 2 11 2 1 11 1 12 9 3 2
11 2 11 11 4 13 15 1 10 0 9 2
23 15 4 13 15 9 7 9 2 7 15 13 15 4 13 3 1 9 2 13 10 0 9 2
15 1 1 9 13 9 2 15 10 9 13 12 9 7 9 2
10 11 13 15 1 2 13 15 1 9 2
11 3 13 15 2 11 2 1 10 0 9 2
36 2 9 10 13 15 3 1 1 15 15 13 2 16 16 9 0 13 0 7 9 13 2 4 15 13 0 9 16 3 10 9 3 4 13 15 2
9 2 4 15 13 0 0 1 9 2
3 2 6 2
6 15 4 13 0 0 2
6 2 4 15 13 0 2
5 2 6 2 1 2
17 15 13 0 16 15 13 0 2 16 15 13 9 1 10 0 9 2
14 1 10 0 4 15 3 13 14 13 3 0 1 9 2
11 7 10 9 13 9 2 3 1 11 11 2
7 2 15 13 3 1 9 2
4 10 0 9 5
26 16 12 1 9 1 9 0 9 2 11 2 13 1 11 1 14 13 2 13 15 3 3 1 9 9 2
10 1 1 13 9 7 13 1 0 9 2
2 9 2
3 11 11 2
11 11 11 2 12 2 13 10 0 11 11 2
24 15 13 0 1 10 9 1 11 1 9 2 7 13 0 1 9 1 16 15 4 13 0 9 2
9 3 1 9 1 11 11 1 11 2
5 0 9 1 9 2
8 10 9 4 13 1 9 11 2
6 13 0 1 9 9 2
3 0 9 2
10 1 11 4 9 13 2 1 9 9 2
8 15 13 11 11 7 11 11 2
5 13 0 1 9 2
5 11 11 1 11 2
3 0 9 2
21 10 1 9 15 13 1 11 1 12 9 3 13 1 3 12 9 7 0 9 9 2
13 15 13 0 14 13 10 9 0 16 10 0 13 2
4 1 1 9 2
15 11 11 7 10 10 9 13 1 1 10 0 9 1 11 2
8 10 0 13 1 11 1 9 2
5 1 10 9 9 2
18 1 11 13 15 9 14 13 10 10 9 1 9 1 9 2 11 2 2
16 15 13 3 0 14 13 9 7 9 2 7 13 15 0 9 2
3 9 13 2
15 10 0 9 1 11 2 1 9 7 9 2 13 12 9 2
10 3 0 11 13 0 1 10 0 9 2
19 9 11 11 7 11 11 13 13 1 12 9 1 11 11 1 9 1 11 2
10 15 13 0 9 1 0 7 0 9 2
19 1 9 13 10 0 9 1 10 0 9 2 15 4 13 1 10 0 9 2
3 15 13 2
25 2 8 2 8 8 8 8 8 8 8 2 8 8 8 8 8 8 8 8 8 8 8 8 2 2
10 1 15 13 12 12 9 7 13 1 2
9 3 3 13 10 0 0 9 9 2
23 15 13 10 0 9 1 14 13 16 15 1 9 13 10 0 9 1 14 4 13 1 9 2
7 3 13 9 1 1 15 2
10 10 0 9 1 9 7 9 4 13 2
26 15 13 0 9 11 11 11 2 9 0 9 2 15 13 1 12 0 7 12 0 9 2 13 1 11 2
8 0 9 13 1 11 1 9 2
24 1 9 13 15 11 1 11 1 12 9 1 11 2 7 11 11 11 1 11 11 11 1 11 2
9 15 13 9 3 3 9 13 15 2
11 15 13 1 11 1 10 0 9 1 15 2
33 1 9 12 13 9 1 10 9 1 11 2 11 11 2 16 9 1 11 13 10 9 14 13 9 1 10 10 0 9 1 1 9 2
26 2 8 8 8 8 8 8 2 8 8 8 8 8 8 2 8 8 8 8 8 8 8 8 2 2 2
5 15 13 3 9 2
22 15 13 3 9 2 10 0 9 11 4 13 1 9 7 9 2 16 9 13 1 11 2
29 15 13 3 9 1 9 1 1 2 10 0 11 2 0 11 11 2 2 1 9 1 11 2 11 2 11 7 11 2
16 7 15 13 3 16 15 4 13 0 14 13 1 9 1 11 2
11 11 2 9 12 13 1 1 14 13 9 2
13 15 13 11 11 2 9 15 13 9 1 10 9 2
3 9 11 2
30 9 15 1 10 9 1 12 9 4 13 1 10 11 11 16 2 4 15 13 9 10 2 3 4 15 13 10 9 2 2
8 11 13 9 0 9 1 11 2
10 15 13 10 12 9 15 4 13 9 2
10 15 4 13 1 9 0 9 1 9 2
14 15 13 9 16 11 7 11 13 10 9 1 10 9 2
13 11 11 13 9 11 11 7 11 11 2 1 3 2
15 9 13 1 9 2 7 15 13 3 0 9 16 11 13 2
16 11 13 9 1 3 12 9 2 1 10 0 0 9 1 11 2
5 15 13 10 9 2
3 1 13 2
4 12 9 0 2
8 11 11 13 1 10 0 9 2
12 1 9 1 15 13 10 10 9 2 11 11 2
6 15 13 0 0 1 2
6 15 13 9 1 9 2
20 15 13 16 15 13 0 14 13 10 0 9 2 7 16 15 3 4 13 0 2
15 10 0 9 13 3 15 13 14 13 9 1 10 10 9 2
9 2 15 13 3 15 13 3 0 2
24 15 13 3 10 10 9 3 1 1 2 7 15 4 13 3 0 1 15 15 13 2 13 11 2
26 3 2 16 11 9 2 11 11 2 13 1 10 0 9 2 13 15 3 1 10 0 9 1 11 9 2
10 15 13 11 11 7 13 1 11 11 2
16 15 13 1 15 0 9 13 1 16 9 10 13 1 0 9 2
19 2 13 15 15 11 9 13 2 16 15 13 16 10 9 4 13 1 9 2
3 2 6 2
20 1 11 13 9 12 9 2 7 15 13 15 3 15 14 13 9 1 12 9 2
15 15 13 3 1 15 13 0 16 9 10 4 13 10 9 2
13 10 0 1 15 13 3 9 1 9 2 13 11 2
4 1 1 9 2
25 11 11 2 9 15 1 15 15 13 15 13 3 3 0 1 11 2 13 9 16 11 13 1 9 2
9 15 13 9 7 13 11 2 9 2
9 3 0 1 13 11 11 1 11 2
19 15 13 9 3 1 9 1 11 11 2 13 15 9 7 13 15 1 9 2
15 1 1 9 13 2 11 8 8 8 2 2 16 9 13 2
7 9 1 9 13 15 3 2
26 15 13 0 1 0 9 1 2 11 2 2 7 15 13 3 0 9 2 15 13 9 1 3 0 9 2
11 1 9 1 11 13 15 9 7 0 9 2
18 10 9 13 0 9 2 1 9 7 9 13 1 1 10 9 1 15 2
12 1 10 12 13 15 2 11 11 2 11 2 2
21 10 0 9 1 11 1 9 2 13 0 1 10 9 2 15 13 3 2 11 2 2
11 3 1 13 11 11 7 13 1 11 9 2
13 9 13 16 9 7 9 4 13 1 1 9 10 2
24 15 4 3 3 13 1 15 16 10 0 9 13 16 15 2 13 9 1 9 1 10 9 2 2
6 9 13 0 1 9 2
14 15 13 1 3 15 13 9 11 4 13 15 10 9 2
14 16 15 13 10 0 9 13 9 1 14 13 15 9 2
16 10 0 9 13 3 15 13 15 13 14 13 11 2 11 11 2
7 11 13 3 0 15 13 2
14 15 13 0 1 15 2 7 13 3 9 10 1 9 2
6 3 13 15 0 9 2
12 10 0 9 13 15 15 4 13 9 1 11 2
16 2 15 13 9 15 13 1 2 11 2 13 2 8 0 2 2
23 7 3 4 15 13 0 14 13 1 9 1 9 7 4 13 1 10 0 9 2 13 11 2
22 10 10 9 13 16 9 13 9 4 13 1 1 9 1 9 1 15 11 13 1 9 2
19 2 1 15 15 4 13 1 9 1 9 7 3 1 9 2 13 15 15 2
10 9 13 15 13 0 16 15 13 3 2
10 2 13 9 3 1 1 2 13 9 2
8 2 6 2 15 13 3 0 2
12 15 13 16 15 4 13 9 2 3 1 1 2
14 15 13 1 15 11 13 1 16 11 4 13 1 11 2
7 2 13 3 15 0 9 2
10 2 15 13 0 15 4 13 1 15 2
31 16 15 13 0 1 9 1 11 2 3 13 15 15 13 0 14 13 3 0 9 15 13 7 3 0 9 15 4 13 3 2
16 7 15 13 0 15 15 13 1 14 13 2 13 15 1 11 2
15 2 7 13 15 9 13 10 10 9 1 9 1 1 11 2
5 2 15 13 15 2
29 15 13 2 10 9 3 1 11 13 0 2 7 15 13 0 16 15 13 9 1 11 1 11 2 7 15 13 15 2
11 11 1 11 13 0 15 15 4 13 1 2
12 2 13 9 1 11 1 10 2 0 2 9 2
9 11 13 1 1 9 10 10 9 2
9 2 6 2 15 13 3 0 0 2
17 15 13 16 15 13 10 10 9 1 0 2 7 9 13 10 10 2
13 15 13 1 10 0 9 1 9 1 10 0 9 2
27 15 13 3 9 1 16 15 13 0 1 11 1 9 2 15 13 3 12 9 1 11 16 3 9 13 0 2
16 7 15 13 3 0 9 16 10 9 13 9 13 1 1 0 2
21 11 4 3 13 12 5 9 2 16 9 11 3 4 13 9 9 1 10 0 9 2
21 1 12 9 2 0 9 12 2 13 9 0 3 16 12 5 9 4 13 1 0 2
27 9 13 16 15 4 13 9 1 3 0 10 0 9 1 10 9 4 13 2 7 3 0 10 9 4 13 2
19 10 9 4 13 10 9 3 2 7 10 0 9 13 3 1 12 9 9 2
15 1 9 4 15 4 13 10 9 1 10 1 9 1 11 2
8 15 13 15 1 10 0 9 2
24 1 9 15 13 15 2 13 15 2 11 11 11 2 11 11 11 11 11 2 11 11 11 2 2
13 15 13 1 1 15 15 13 1 10 0 0 9 2
23 2 11 2 13 9 1 11 16 15 0 13 2 1 1 9 2 1 9 1 12 5 9 2
3 2 0 2
12 15 4 13 10 0 9 1 10 9 1 9 2
16 0 9 2 0 9 7 0 9 2 0 9 2 0 0 9 2
19 1 9 2 16 15 13 1 9 1 9 10 2 13 15 16 15 13 0 2
19 15 13 3 10 9 16 15 13 0 0 9 2 1 11 11 7 11 11 2
13 2 15 1 10 9 13 15 15 13 1 1 11 2
6 2 6 2 0 9 2
17 16 15 0 13 2 3 13 1 12 9 1 9 1 11 1 11 2
10 15 4 3 1 7 1 13 10 9 2
22 1 10 9 2 16 3 0 1 9 10 13 0 2 13 3 9 1 11 0 3 1 2
24 15 13 10 1 9 15 13 1 14 13 9 0 11 2 7 3 3 9 7 9 1 9 10 2
13 15 14 13 0 9 3 1 13 16 15 13 9 2
11 2 13 15 0 9 1 0 2 9 2 2
8 2 6 2 6 2 3 3 2
9 15 13 1 14 13 9 0 9 2
25 15 4 13 0 16 15 13 0 1 10 0 9 2 7 15 13 3 1 9 10 1 10 0 9 2
15 10 9 13 3 1 15 15 13 2 7 15 13 0 9 2
17 9 13 3 2 7 15 13 10 9 1 9 15 4 13 1 9 2
11 10 9 9 13 2 13 0 9 1 9 2
4 9 13 1 2
17 9 11 10 9 2 11 8 8 2 2 13 3 3 0 1 9 2
27 7 3 16 10 9 1 9 13 7 9 7 9 9 1 14 13 9 2 13 0 1 9 1 9 0 0 2
18 12 9 1 9 1 0 9 4 9 13 2 3 16 9 4 13 9 2
23 1 15 13 15 10 9 1 10 9 7 9 1 1 12 9 2 15 3 4 13 0 9 2
2 9 2
10 2 15 4 13 10 9 2 10 9 2
2 9 2
11 2 4 15 3 13 10 9 1 10 9 2
2 9 2
3 2 6 2
2 9 2
11 2 4 15 3 13 10 9 1 12 9 2
2 9 2
3 2 6 2
2 9 2
11 2 4 15 3 13 10 9 1 12 9 2
2 9 2
13 2 6 2 15 4 3 13 10 9 1 12 9 2
9 15 13 15 11 13 14 13 1 2
12 9 13 9 2 3 0 3 12 9 4 13 2
15 1 9 13 15 3 1 9 1 9 15 13 0 1 15 2
7 9 13 1 9 1 9 2
22 1 9 13 15 1 9 1 15 15 13 2 7 3 0 15 13 7 3 0 15 13 2
24 1 10 9 0 9 2 16 10 9 13 10 10 16 9 13 2 13 10 12 9 1 10 10 2
12 2 6 2 13 15 3 13 1 1 15 2 2
9 15 13 1 1 11 11 1 11 2
13 2 13 15 1 1 9 1 10 0 9 2 11 2
9 2 15 4 3 13 11 7 11 2
12 15 13 12 9 9 7 15 13 12 9 9 2
9 15 4 3 13 9 1 9 3 2
27 0 13 15 0 16 15 13 1 11 2 7 16 15 13 0 2 16 15 13 0 9 7 9 1 0 9 2
10 7 15 13 3 9 15 13 9 1 2
25 15 13 3 3 15 13 1 9 7 15 13 3 0 0 1 9 15 4 13 1 15 1 3 15 2
16 7 16 15 4 13 2 3 13 15 3 1 11 1 10 9 2
35 15 13 3 15 13 9 15 13 1 10 9 2 7 16 15 13 3 1 15 1 14 2 15 13 2 13 9 1 14 13 1 10 0 9 2
14 2 13 15 0 10 9 16 15 13 0 9 1 9 2
15 2 15 13 1 14 13 9 1 11 2 3 10 10 9 2
22 15 13 15 15 13 0 1 2 16 0 9 4 4 13 1 0 9 7 0 9 0 2
18 2 7 15 4 4 13 1 16 11 7 11 4 13 1 10 0 9 2
19 2 15 13 3 3 1 14 13 10 9 1 9 7 13 16 11 13 10 2
8 7 15 7 9 13 10 9 2
7 15 13 3 14 13 11 2
26 15 13 10 9 1 16 16 15 4 13 12 9 1 12 9 1 11 2 3 4 3 9 13 3 0 2
6 7 2 15 13 15 2
3 11 13 2
9 7 1 10 9 13 15 0 0 2
28 2 0 9 4 13 1 16 11 9 4 13 10 9 2 16 0 9 13 0 1 0 9 1 14 13 0 9 2
4 13 15 15 2
34 2 15 13 3 9 1 10 9 2 7 15 13 16 16 0 10 0 9 4 13 1 2 4 15 13 10 9 1 10 9 2 3 10 2
16 9 13 3 1 2 7 3 1 9 13 11 1 12 2 12 2
34 15 13 12 9 0 9 2 7 4 3 9 13 15 15 13 1 1 12 9 2 13 15 15 1 10 9 12 9 16 9 13 1 9 2
20 11 11 13 9 1 9 2 1 11 9 2 13 9 7 13 1 1 0 9 2
8 11 13 1 10 3 0 9 2
4 9 13 1 2
9 15 13 1 10 0 9 1 9 2
5 1 9 13 9 2
20 15 13 0 1 9 2 7 0 1 15 4 0 16 9 11 11 9 3 13 2
3 11 9 2
4 3 13 11 2
7 1 13 10 9 1 9 2
7 15 13 0 3 10 3 2
9 15 13 0 9 1 10 9 1 2
7 10 1 15 13 1 9 2
14 15 13 16 11 13 0 1 11 1 10 9 9 3 2
7 3 4 15 13 3 0 2
12 10 9 1 9 13 0 1 9 1 9 10 2
11 2 11 12 2 2 13 15 1 9 10 2
7 15 13 1 9 1 9 2
3 9 13 2
11 0 4 2 11 12 2 7 9 13 3 2
16 9 1 13 15 1 1 11 2 1 0 9 1 9 7 9 2
12 1 9 13 11 3 0 15 11 11 13 0 2
17 9 4 13 1 10 0 9 2 7 4 13 1 0 9 1 11 2
31 1 0 9 1 9 4 12 12 9 13 3 1 9 1 14 13 9 2 4 13 0 1 9 7 13 12 1 9 0 9 2
32 1 9 1 1 9 13 15 11 11 2 15 13 9 1 9 11 2 11 8 11 11 11 2 1 11 2 11 7 9 1 11 2
27 15 13 16 9 11 2 11 11 11 11 2 4 13 1 1 11 2 7 4 13 9 1 11 11 1 9 2
9 15 4 0 3 13 1 11 11 2
11 15 13 3 9 1 11 13 0 1 9 2
26 2 11 13 7 0 9 2 9 2 9 7 11 2 7 3 13 15 3 1 14 13 0 0 1 11 2
9 15 13 2 9 13 0 1 11 2
16 11 13 0 1 9 1 11 2 11 2 11 2 11 7 11 2
33 16 15 13 1 15 3 1 11 2 4 15 13 9 1 15 2 7 9 10 13 16 15 13 15 15 13 0 11 1 11 1 15 2
21 15 13 1 16 9 3 13 12 9 9 1 11 2 1 9 1 12 12 1 12 2
16 9 1 11 9 13 3 1 1 0 9 2 7 15 13 9 2
24 3 9 10 2 11 11 2 10 1 9 1 11 2 4 13 1 10 0 9 1 10 0 9 2
13 2 15 13 15 15 13 1 14 13 11 1 11 2
18 15 13 16 0 9 4 13 0 3 0 2 7 13 9 13 3 0 2
20 16 10 9 4 13 9 0 9 1 0 9 2 4 15 13 0 2 13 15 2
16 9 9 12 1 11 7 11 13 0 0 1 15 9 1 9 2
33 3 13 3 10 0 1 9 3 1 9 2 7 3 16 15 0 13 0 1 14 13 11 2 11 7 11 2 13 9 3 0 1 2
10 1 0 9 13 9 11 11 1 9 2
13 15 13 1 9 2 7 1 9 13 0 10 10 2
30 11 13 0 0 1 9 2 16 0 13 15 13 0 9 1 9 1 12 9 3 2 7 16 15 3 3 13 9 0 2
8 15 4 3 9 13 1 15 2
13 1 9 4 11 10 0 13 1 1 12 2 12 2
15 11 11 13 0 1 16 11 3 4 13 14 13 1 9 2
22 16 9 10 13 1 9 2 13 15 9 0 9 1 9 7 13 15 1 15 1 9 2
22 10 9 1 9 13 1 9 1 11 7 13 15 0 0 1 10 9 9 13 1 9 2
18 3 1 2 1 10 1 10 0 9 1 9 2 13 10 9 1 9 2
2 9 2
3 11 11 2
15 15 13 9 10 16 15 13 1 1 9 3 1 1 9 2
36 2 8 8 8 8 8 8 8 2 8 8 8 8 8 8 8 2 8 8 8 8 8 8 2 8 8 8 8 8 8 8 8 8 8 2 2
8 9 13 12 2 12 1 11 2
10 9 13 3 12 9 10 1 12 9 2
16 1 9 13 15 11 9 7 9 11 11 15 13 9 1 9 2
13 3 1 4 9 13 1 2 10 10 2 11 11 2
17 15 4 13 1 10 0 9 15 13 1 9 16 15 13 1 9 2
5 2 15 13 0 2
23 16 15 13 12 2 12 1 9 2 4 15 13 15 10 9 1 14 13 1 10 0 9 2
8 15 13 15 3 1 14 13 2
10 3 1 13 15 9 11 11 1 0 2
10 2 13 15 0 1 16 15 13 11 2
3 2 0 2
10 15 13 3 1 9 3 1 10 9 2
6 7 9 4 13 0 2
15 2 3 15 4 13 1 14 13 11 1 11 1 12 9 2
5 2 6 2 11 2
4 8 8 8 2
6 11 11 1 0 9 5
14 3 0 15 13 15 13 0 14 13 1 15 1 9 2
2 9 2
13 0 9 13 3 9 1 9 2 0 3 1 9 2
16 3 13 9 11 11 10 9 1 10 2 11 15 13 2 9 2
17 2 15 13 0 1 16 15 13 15 13 3 0 1 10 10 9 2
11 3 13 15 10 0 0 9 2 13 9 2
2 9 2
14 9 1 9 4 13 0 1 0 9 1 9 1 9 2
4 3 13 10 2
4 11 11 9 2
2 8 2
14 15 13 3 1 9 1 9 1 14 13 9 1 9 2
2 9 2
16 11 11 1 10 0 9 11 13 9 7 9 1 10 0 9 2
2 9 2
21 1 9 11 1 11 13 9 9 0 1 14 13 9 9 1 1 0 0 0 9 2
7 2 3 0 2 3 0 2
18 9 13 14 13 0 0 7 13 10 9 1 9 2 13 9 11 11 2
21 2 16 15 13 9 2 13 15 16 15 13 0 1 1 9 2 13 11 11 11 2
15 9 7 10 0 9 13 10 0 2 0 9 1 1 15 2
24 9 1 9 1 9 1 11 13 0 10 3 12 9 9 1 9 2 16 15 13 1 10 9 2
34 9 4 11 13 1 15 16 15 4 13 9 1 11 11 11 1 9 2 11 15 13 2 1 11 12 1 3 12 12 9 12 9 0 2
13 2 15 13 10 0 0 9 1 15 2 13 11 2
21 2 7 15 13 0 1 14 13 1 1 10 9 2 7 13 15 0 0 1 9 2
25 11 11 2 15 3 4 13 0 1 11 12 0 9 2 13 10 0 0 0 9 1 10 0 9 2
18 2 15 13 16 15 13 15 1 2 3 16 15 13 15 2 13 15 2
18 2 7 15 13 0 1 16 15 13 15 13 3 0 1 10 10 9 2
19 3 13 15 10 0 0 9 2 13 9 2 15 13 12 1 9 1 9 2
12 10 9 1 9 13 9 0 1 1 9 9 2
43 9 15 1 9 13 9 2 4 13 10 9 15 13 1 10 0 10 9 1 9 1 0 2 7 15 13 10 0 7 0 9 16 15 0 4 13 3 0 9 7 0 9 2
8 7 3 0 9 7 0 9 2
7 2 3 0 2 3 0 2
26 9 13 14 13 0 0 7 13 9 2 13 10 9 1 9 2 3 0 2 13 9 11 11 1 11 2
24 1 10 0 0 9 1 1 11 13 12 9 1 14 13 0 0 9 7 9 1 9 9 1 2
30 3 9 1 2 11 15 13 2 1 0 9 1 9 2 7 10 12 9 1 10 0 9 2 11 11 11 2 1 11 2
11 2 15 13 3 1 9 2 15 13 9 2
7 15 4 3 13 10 0 2
26 15 13 1 1 0 2 0 9 7 1 1 10 9 2 16 15 13 1 14 13 10 0 7 13 9 2
19 15 4 13 1 14 13 1 15 9 1 9 2 13 11 2 15 13 1 2
10 2 7 10 0 9 13 3 3 0 2
16 15 4 3 13 0 14 13 1 15 7 13 9 9 0 0 2
22 15 13 0 16 15 15 13 15 1 15 13 0 2 3 13 15 3 13 15 1 9 2
10 15 4 3 3 13 1 9 7 9 2
42 11 11 11 2 15 13 9 1 2 11 15 13 2 7 4 13 1 12 9 7 12 9 1 9 2 13 16 15 13 0 9 15 13 16 15 10 13 14 13 1 9 2
8 2 10 0 9 13 1 9 2
12 3 13 15 0 9 2 3 9 2 3 9 2
26 1 9 4 3 0 9 7 9 13 0 0 2 7 9 4 13 15 0 0 7 0 9 2 13 15 2
25 11 11 2 15 13 9 1 11 9 7 9 7 0 9 2 13 3 9 4 13 0 0 1 9 2
15 2 15 13 12 9 15 4 13 1 10 9 2 13 15 2
15 2 0 13 15 9 1 15 15 4 13 1 15 7 3 2
14 15 13 10 9 1 10 9 3 3 9 13 3 0 2
16 3 13 15 0 9 1 2 7 15 13 0 9 2 13 15 2
20 1 10 0 9 13 15 1 10 16 2 8 8 8 8 8 8 8 8 2 2
11 7 10 9 10 0 9 2 15 11 13 2
12 15 13 1 9 9 13 14 13 9 1 9 2
27 1 9 7 9 13 3 10 0 2 9 2 2 9 2 9 2 9 2 9 7 9 2 1 10 0 9 2
25 3 1 9 13 2 9 2 2 9 2 9 2 9 2 9 9 7 9 2 10 9 1 0 9 2
9 3 13 9 2 7 9 13 15 2
24 2 3 13 11 11 2 9 13 0 2 7 15 13 0 14 13 10 1 15 2 13 11 11 2
14 16 9 13 13 1 14 13 10 0 9 1 10 9 2
12 3 13 9 15 1 1 10 0 9 1 9 2
12 2 9 13 1 0 9 2 13 11 11 11 2
18 2 3 13 15 9 1 9 7 9 1 9 1 11 11 7 11 11 2
15 9 13 0 2 3 4 9 13 15 7 9 13 0 0 2
5 9 13 0 9 2
11 2 7 9 13 3 3 2 13 11 11 2
11 2 9 13 1 0 1 1 9 1 9 2
11 3 13 15 0 7 0 1 9 7 9 2
26 7 9 15 13 1 10 9 1 10 9 3 2 13 3 14 13 1 10 0 13 1 9 2 13 15 2
12 7 9 13 3 10 0 9 1 9 1 0 2
27 2 15 13 10 9 1 9 1 9 3 2 1 9 2 9 7 0 9 2 13 9 1 11 2 11 11 2
23 2 7 16 9 13 9 2 13 15 1 16 15 13 2 0 13 0 2 15 13 1 9 2
22 7 13 15 3 0 3 15 4 13 2 7 3 13 15 15 0 7 0 3 1 15 2
21 15 13 3 3 15 13 10 0 2 13 11 2 15 13 9 13 0 1 10 9 2
21 2 15 13 1 16 15 13 1 10 10 9 2 7 4 13 10 10 0 0 9 2
15 9 13 15 3 3 2 7 15 13 0 9 2 13 11 2
18 9 1 2 11 15 13 2 2 11 11 2 13 1 9 1 11 11 2
26 15 13 0 1 9 2 9 2 9 7 0 9 1 9 15 10 9 13 1 1 9 1 9 1 9 2
18 3 13 15 9 15 13 3 0 1 10 0 9 1 9 1 3 0 2
8 3 1 9 2 9 7 9 2
13 7 3 0 9 1 9 7 9 7 9 1 9 2
7 12 9 13 1 10 9 2
30 1 9 1 14 13 1 11 1 14 13 9 7 13 1 9 7 9 16 15 13 9 2 4 11 3 3 13 0 9 2
23 2 9 2 4 15 13 1 15 15 3 2 2 13 15 0 1 9 2 13 15 7 13 2
5 2 0 1 9 2
10 11 11 11 13 3 3 0 1 9 2
22 3 13 15 16 15 13 10 9 7 10 9 2 7 13 1 1 7 0 9 7 9 2
14 11 4 13 1 10 12 9 1 2 11 15 13 2 2
25 2 15 4 13 1 9 1 9 2 15 15 4 13 7 10 9 15 4 13 16 15 13 3 9 2
9 9 4 13 1 9 7 13 9 2
15 7 15 13 0 9 1 9 2 3 16 15 4 13 0 2
10 9 13 15 3 10 9 1 1 9 2
21 2 15 4 3 13 1 9 1 9 1 14 13 15 0 7 0 2 13 11 11 2
20 2 15 13 7 9 7 15 16 15 13 15 2 15 15 3 13 9 1 9 2
7 15 13 0 0 1 9 2
17 3 13 9 1 0 9 1 9 2 7 9 7 9 13 10 10 2
13 1 9 13 12 9 0 11 11 1 9 7 9 2
17 10 9 1 0 7 0 9 2 0 0 1 9 2 13 1 15 2
22 10 0 9 4 3 3 13 11 13 1 9 16 15 13 1 11 11 11 10 9 9 2
24 7 10 0 9 15 13 1 11 1 12 1 14 13 1 10 0 9 2 13 3 10 10 9 2
20 0 1 15 4 15 2 1 0 11 11 9 2 13 1 2 11 15 13 2 2
27 2 15 4 13 15 12 9 9 2 13 15 1 10 0 9 15 13 14 4 13 9 1 16 9 13 1 2
13 2 9 13 0 2 7 3 4 15 13 1 9 2
11 15 13 2 7 15 13 3 0 1 9 2
18 7 12 9 9 13 3 3 0 13 1 9 1 10 0 9 1 11 2
6 15 13 0 12 9 2
16 9 13 10 0 0 9 1 9 7 0 7 0 9 1 9 2
35 2 15 13 10 9 1 16 15 4 13 0 1 9 2 13 11 2 15 4 13 16 15 13 12 9 0 7 13 10 10 9 3 3 0 2
11 16 15 13 9 13 15 14 13 15 3 2
17 2 10 0 13 16 15 0 3 13 3 0 1 9 2 13 15 2
13 2 7 9 13 3 0 1 16 15 3 13 0 2
22 15 15 4 13 10 0 9 4 13 0 1 1 9 2 16 15 3 13 12 9 0 2
25 15 13 0 14 13 15 15 13 0 2 15 13 16 9 13 15 7 13 2 15 13 15 2 2 2
23 7 3 16 15 13 10 3 10 11 13 1 15 10 0 0 9 2 13 15 0 1 9 2
28 2 9 13 10 12 9 1 9 1 9 16 15 4 13 1 3 0 9 1 16 15 13 0 1 2 13 15 2
16 2 7 15 13 15 0 0 16 15 13 1 10 9 1 9 2
20 15 13 3 3 3 15 13 9 1 14 13 1 10 9 16 15 4 13 0 2
8 11 11 13 3 0 1 9 2
18 2 1 9 13 15 16 15 1 9 3 4 13 10 9 2 13 15 2
37 2 7 15 13 15 13 0 14 13 3 10 1 10 9 13 10 10 9 2 16 9 7 9 13 3 1 10 9 7 10 9 15 13 10 0 9 2
12 15 13 10 9 1 16 15 13 15 15 13 2
16 15 4 13 12 9 2 9 2 9 2 9 7 9 1 9 5
3 11 11 2
2 0 2
14 11 4 13 10 10 9 1 9 7 13 0 9 1 2
2 0 2
10 9 4 3 13 1 9 1 12 9 2
6 2 10 0 0 9 2
3 1 9 2
12 9 15 1 3 4 13 1 9 1 1 11 2
8 15 13 10 9 1 11 11 2
29 3 4 9 1 9 7 9 11 11 13 1 10 9 2 1 9 1 0 0 9 1 9 2 11 10 0 9 2 2
6 2 15 4 13 9 2
27 3 13 15 9 2 9 2 9 2 9 7 9 2 13 11 16 15 13 3 1 9 13 1 9 11 11 2
23 3 4 15 13 1 0 9 2 9 7 9 15 4 13 1 1 3 12 9 1 12 9 2
26 15 13 0 9 1 9 1 9 2 9 15 13 9 1 10 9 7 9 15 13 1 14 4 13 11 2
25 1 9 1 12 0 2 12 1 9 15 13 1 9 7 10 9 1 10 0 9 7 10 9 1 2
31 1 9 13 15 3 9 1 10 12 9 0 9 15 13 1 9 1 0 9 7 9 2 9 10 13 14 13 9 10 2 2
29 0 13 1 9 7 9 11 11 13 1 9 1 9 1 10 9 0 16 15 13 2 1 10 9 1 13 10 9 2
37 2 15 4 13 1 9 1 9 1 0 9 2 7 15 13 1 10 3 0 9 1 10 10 9 16 15 13 9 1 14 13 15 1 10 0 9 2
14 7 15 13 9 1 9 1 10 10 9 2 13 11 2
16 2 3 4 15 13 14 13 10 10 9 3 0 1 9 10 2
15 2 15 13 0 14 13 9 1 15 15 13 0 1 15 2
8 9 13 0 9 7 0 9 2
14 15 13 14 13 15 1 9 7 9 2 9 7 9 2
14 15 13 0 14 13 15 1 12 0 9 2 13 15 2
17 2 13 15 3 3 0 15 13 0 16 15 4 13 10 10 9 2
9 2 1 0 9 13 15 3 15 2
13 15 13 10 0 9 2 7 15 13 10 0 9 2
7 15 4 3 13 9 3 2
19 1 9 1 14 13 9 1 15 4 15 3 13 14 13 1 10 0 9 2
15 9 13 14 13 10 0 2 15 10 4 13 15 3 1 2
20 2 9 1 9 10 13 0 0 2 13 15 0 1 9 1 9 14 13 15 2
20 2 15 13 0 9 10 15 13 9 1 9 7 13 15 4 13 15 1 15 2
18 1 10 9 4 15 13 15 1 15 1 12 9 1 14 13 15 1 2
18 15 4 13 1 16 15 13 1 0 2 16 15 4 13 0 1 10 2
10 2 13 10 9 0 0 2 13 15 2
9 2 6 2 15 13 3 0 0 2
6 10 9 13 10 9 2
12 7 9 13 0 16 15 13 16 15 13 9 2
10 15 13 1 1 10 0 2 0 9 2
13 15 13 3 16 15 13 12 7 0 16 15 13 2
5 9 13 3 0 2
9 15 13 10 9 16 15 13 15 2
15 7 3 13 9 14 13 2 7 14 13 0 2 13 11 2
18 9 10 13 10 0 9 1 11 7 13 1 12 7 10 0 9 3 2
21 1 9 1 9 1 9 10 4 15 3 13 9 2 10 1 12 9 2 1 9 2
14 15 13 1 10 9 16 11 13 10 9 1 10 9 2
17 3 1 10 9 13 9 16 15 13 10 9 15 13 10 10 9 2
10 0 9 4 9 13 1 11 1 11 2
15 11 9 2 9 11 11 2 4 13 10 10 9 1 9 2
37 15 4 3 13 1 10 9 2 1 10 10 0 9 2 10 9 15 4 13 9 10 0 9 1 10 9 16 11 7 10 9 13 1 15 1 9 2
11 1 9 1 9 4 9 2 9 2 13 2
19 3 4 11 11 13 10 9 2 9 11 11 2 1 11 2 11 7 11 2
36 15 13 1 15 10 0 9 13 1 15 15 13 15 1 9 2 7 9 4 3 13 1 9 16 10 12 13 1 9 7 13 1 0 7 0 2
9 1 9 4 15 13 9 1 9 2
24 15 13 0 14 13 1 9 1 10 9 1 0 9 2 7 15 13 3 11 11 0 0 1 2
9 2 15 13 0 0 2 0 9 2
8 7 15 13 3 1 10 9 2
22 15 4 3 13 1 15 14 13 10 0 9 1 12 16 10 9 1 11 13 1 9 2
23 3 13 15 1 16 9 4 13 3 0 1 9 10 16 10 9 3 4 13 1 0 9 2
19 3 16 9 1 9 7 10 15 4 13 1 9 2 3 4 0 13 3 2
15 2 15 13 0 0 1 16 15 4 13 7 13 15 1 2
9 9 13 3 15 10 1 9 10 2
2 11 5
18 9 11 11 2 12 2 1 9 2 9 7 9 1 16 9 4 13 2
2 9 2
5 2 15 13 3 2
7 11 7 10 0 9 11 2
4 0 1 9 2
10 2 15 13 3 3 10 9 14 13 2
10 3 16 15 13 1 15 2 13 11 2
7 15 13 0 14 13 0 2
2 9 2
10 9 1 10 0 9 1 10 0 9 2
2 9 2
9 9 4 13 1 11 11 1 12 2
3 0 9 2
12 2 4 15 13 10 10 0 0 9 10 9 2
4 9 7 9 2
13 11 7 9 11 11 15 4 13 0 9 1 11 2
4 9 7 9 2
11 11 7 9 11 13 1 9 1 9 11 2
7 11 13 3 1 1 11 2
4 9 1 9 2
12 12 0 9 7 12 0 2 0 13 9 11 2
10 15 13 0 9 2 9 13 1 9 2
44 7 9 2 9 13 0 1 11 2 15 13 1 1 9 15 13 1 9 2 1 0 9 7 10 0 9 1 9 12 2 7 15 13 1 9 1 10 0 11 1 9 1 11 2
18 1 9 13 11 11 2 9 2 9 2 9 2 9 7 9 1 11 2
10 15 13 9 1 9 1 10 0 9 2
13 0 2 0 9 13 15 1 1 10 0 0 9 2
8 10 0 9 13 1 1 9 2
6 2 15 13 0 0 2
14 9 13 1 9 1 9 2 7 11 13 1 1 9 2
6 2 0 2 0 9 2
4 0 7 0 2
13 7 3 0 9 7 9 15 13 1 1 10 9 2
5 15 13 3 0 2
8 15 4 13 0 7 0 3 2
10 16 9 13 10 9 7 9 4 13 2
21 16 11 13 1 9 7 9 0 1 0 9 7 1 11 2 4 15 0 13 9 2
13 10 9 13 10 0 9 1 0 9 1 11 9 2
11 15 13 3 7 13 2 13 1 10 9 2
10 11 13 3 1 15 10 9 1 9 2
12 15 4 13 1 9 7 13 1 10 0 9 2
13 9 12 2 1 9 9 2 13 11 12 0 9 2
4 15 13 11 2
13 1 9 13 15 1 9 2 9 2 9 2 9 2
34 3 2 12 9 0 2 13 10 0 9 15 2 2 2 15 4 13 2 9 9 2 16 9 13 1 0 9 2 0 9 2 0 9 2
8 15 13 10 9 9 1 9 2
8 9 13 3 0 0 1 9 2
16 15 13 0 0 1 9 3 2 7 3 13 15 15 15 13 2
13 9 13 7 13 2 7 3 4 15 7 15 13 2
13 1 10 0 9 4 9 10 11 13 12 1 9 2
11 2 10 0 9 13 10 10 9 1 9 2
14 3 13 15 1 9 10 14 13 9 1 9 1 9 2
8 2 15 13 0 0 1 9 2
15 1 10 9 13 15 3 0 0 9 1 9 1 10 9 2
4 0 1 15 2
9 10 0 9 13 14 13 1 9 2
16 3 4 15 13 1 2 3 4 15 13 0 2 3 13 15 2
6 15 13 3 3 0 2
16 2 4 15 13 1 1 10 9 2 7 15 4 13 11 0 2
15 3 4 15 13 11 2 11 2 6 2 3 0 1 11 2
6 15 13 0 3 1 2
8 9 1 13 15 1 0 9 2
9 11 13 7 13 1 9 7 9 2
10 15 13 15 13 7 13 3 10 9 2
4 3 1 9 2
19 2 15 13 0 0 1 9 2 7 15 4 13 1 14 13 15 1 9 2
6 3 13 15 0 9 2
7 2 13 15 0 14 13 2
5 2 6 2 1 2
12 15 4 13 1 15 0 9 16 15 4 13 2
26 1 7 1 13 15 3 0 16 15 13 10 9 9 2 7 15 4 3 13 10 9 1 9 1 15 2
13 2 13 15 0 1 16 9 10 9 13 14 13 2
3 2 6 2
10 7 15 4 3 4 13 9 1 9 2
10 15 4 3 13 9 1 9 7 9 2
6 15 4 13 1 9 2
5 15 13 0 0 2
6 11 13 9 1 9 2
7 2 15 13 3 9 15 2
10 15 4 13 7 13 2 13 7 13 2
7 7 1 12 13 11 3 2
3 1 9 2
17 15 13 12 9 1 9 2 11 9 2 7 2 11 0 9 2 2
13 12 0 9 2 0 9 1 11 2 0 11 11 2
11 7 3 3 2 1 9 2 13 15 15 2
36 11 11 2 15 4 13 9 1 12 9 2 13 10 9 9 1 9 7 11 13 1 10 9 16 15 13 2 0 14 13 9 1 11 11 2 2
6 15 13 0 1 11 2
11 2 15 4 3 4 13 3 15 15 13 2
8 3 4 15 13 9 1 11 2
7 15 13 15 0 0 1 2
4 2 3 15 2
10 2 15 13 3 15 15 13 1 10 2
24 16 3 9 13 2 7 9 4 13 1 1 15 15 0 13 1 1 2 3 13 15 0 9 2
5 2 3 13 9 2
8 2 15 13 15 3 0 1 2
13 7 15 13 3 15 15 13 10 0 9 1 9 2
38 9 7 9 1 14 13 1 3 2 13 1 0 9 2 13 0 9 2 16 15 13 3 15 13 2 16 15 4 13 1 10 9 2 13 0 1 15 2
15 15 13 1 10 9 16 15 3 13 9 1 14 13 3 2
8 7 15 4 15 13 15 1 2
4 15 13 0 2
10 7 15 13 3 14 13 0 1 9 2
10 2 7 15 13 3 3 0 1 9 2
3 2 6 2
9 2 7 15 13 10 0 0 9 2
10 7 15 13 0 9 14 13 0 1 2
8 2 3 4 15 13 9 10 2
10 2 3 0 2 0 7 0 1 15 2
18 7 15 13 3 0 1 14 13 9 7 13 13 16 15 13 3 0 2
8 15 13 3 15 13 15 13 2
9 2 4 15 13 1 11 11 3 2
7 2 6 2 15 13 15 2
8 15 13 10 0 7 0 9 2
24 15 13 15 13 0 0 1 10 9 16 15 13 3 7 3 2 3 16 15 13 0 0 9 2
9 2 3 4 15 13 9 12 9 2
9 3 13 15 1 2 13 15 11 2
3 2 6 2
6 15 4 3 13 15 2
15 11 11 2 10 0 9 2 13 1 1 9 16 15 13 2
11 7 15 4 3 13 3 0 14 13 9 2
10 11 11 13 7 0 9 7 9 1 2
22 11 11 2 12 2 13 1 9 11 2 7 13 12 9 16 11 13 1 10 0 9 2
12 2 15 13 1 9 15 0 9 13 1 9 2
7 15 13 15 0 7 0 2
3 2 6 2
16 15 4 13 1 7 0 7 0 9 2 15 2 1 0 9 2
13 3 13 15 10 0 1 10 15 13 0 7 0 2
13 15 13 1 9 1 0 9 2 0 9 2 0 2
7 1 1 10 9 13 9 2
8 2 10 10 9 4 15 13 2
7 15 13 9 2 13 15 2
14 15 13 3 3 9 13 1 9 1 10 9 1 11 2
2 6 2
9 12 1 12 9 13 15 10 9 2
15 15 13 1 0 9 2 7 3 3 0 16 15 13 0 2
14 2 7 15 13 10 9 1 9 15 13 0 1 9 2
16 11 13 14 13 3 1 9 2 13 1 9 2 9 2 9 2
5 16 15 13 0 2
10 2 15 13 14 13 1 9 1 9 2
12 13 9 15 13 1 9 2 16 15 13 1 2
38 3 13 15 16 15 4 13 10 0 9 2 3 3 16 15 4 13 3 0 9 2 7 3 16 15 4 13 15 1 7 13 1 15 15 3 4 13 2
24 15 13 0 0 9 1 9 2 7 15 13 3 3 0 14 13 1 15 1 14 13 9 10 2
11 15 13 3 16 15 3 13 10 0 1 2
7 9 13 15 9 1 9 2
18 1 12 4 15 13 2 7 15 4 13 16 15 4 13 9 7 9 2
6 9 13 3 10 9 2
7 2 15 13 14 13 9 2
5 15 13 1 9 2
6 9 13 0 1 9 2
10 2 15 4 13 0 3 1 1 9 2
5 15 4 13 1 2
15 11 13 1 9 2 13 14 13 1 9 7 9 13 1 2
32 10 0 9 1 12 2 1 10 0 9 15 15 13 3 10 9 1 9 2 13 0 1 10 0 9 1 10 0 9 1 11 2
24 9 4 13 1 9 2 9 2 9 7 9 2 7 1 9 13 10 9 15 0 1 10 9 2
22 11 13 1 1 9 2 9 15 15 13 15 2 13 1 9 7 13 15 1 1 9 2
40 15 13 9 1 10 9 2 12 9 2 10 0 9 0 1 9 2 12 9 2 10 9 2 9 7 10 0 9 1 9 15 4 13 1 10 9 1 1 9 2
20 15 13 9 1 10 9 1 12 2 1 9 7 10 0 2 1 9 7 9 2
22 3 4 0 1 11 9 7 4 13 7 13 1 2 7 1 10 9 1 9 13 9 2
4 12 0 9 2
3 12 11 2
16 1 9 4 10 9 13 1 9 1 11 2 0 1 1 9 2
8 9 13 0 2 0 7 0 2
5 2 0 9 2 2
5 2 0 11 2 2
7 2 10 9 1 1 2 2
5 2 9 9 2 2
7 2 0 2 0 11 2 2
6 2 9 13 0 2 2
5 2 0 11 2 2
10 2 7 3 13 10 3 0 9 10 2
17 15 13 3 11 13 11 2 1 10 9 15 1 9 7 9 13 2
11 15 13 9 2 9 7 13 9 1 9 2
9 1 9 13 10 0 2 0 9 2
16 1 10 9 1 1 0 9 4 15 13 10 0 9 1 9 2
10 11 2 11 2 11 2 11 7 11 2
9 9 4 13 12 9 1 12 9 2
8 1 10 9 4 11 13 9 2
23 15 4 13 9 2 15 4 13 9 2 13 1 9 7 9 2 13 9 2 9 7 9 2
48 9 1 9 2 16 15 4 13 9 2 16 15 4 13 1 9 2 16 15 13 9 2 16 15 4 13 10 12 0 9 1 9 2 6 2 10 15 2 4 11 13 7 13 1 1 10 9 2
10 2 4 15 13 16 15 4 13 9 2
3 2 6 2
12 15 4 13 15 1 14 13 9 3 10 9 2
6 9 12 9 1 9 2
15 2 4 10 10 3 13 15 15 4 13 1 15 1 9 2
3 2 6 2
6 6 2 15 13 15 2
23 7 16 11 11 1 10 0 13 13 14 13 9 1 10 15 2 4 15 4 4 13 1 2
23 1 15 13 10 9 15 4 13 1 9 16 15 13 1 15 7 15 3 13 9 1 9 2
19 15 4 4 4 13 0 9 1 9 2 7 15 13 9 15 13 15 10 2
10 11 4 13 1 9 1 11 1 9 2
12 15 13 2 13 9 13 1 9 7 13 1 2
15 9 12 2 3 10 0 9 0 2 13 9 1 1 11 2
5 15 13 1 9 2
17 15 13 1 16 15 13 10 9 15 13 7 13 1 9 1 9 2
4 15 13 15 2
11 11 4 13 0 1 1 9 7 13 1 2
7 2 15 13 0 3 0 2
15 15 13 9 7 13 0 0 9 14 13 1 10 10 9 2
18 7 10 10 10 2 15 13 1 9 14 13 2 15 13 3 10 9 2
6 15 13 3 0 9 2
14 15 13 10 1 14 4 13 1 1 9 1 10 9 2
8 15 3 13 15 13 0 9 2
15 15 3 13 16 15 3 13 1 15 15 13 0 1 15 2
8 15 13 15 15 13 1 11 2
7 15 15 10 13 4 13 2
10 1 12 9 4 15 13 3 1 11 2
9 1 0 1 9 4 15 13 0 2
7 1 12 9 13 15 9 2
10 11 13 9 7 13 15 1 1 9 2
12 2 15 13 0 0 1 15 14 13 10 9 2
4 15 13 15 2
7 15 4 13 1 12 9 2
11 1 9 4 15 13 0 0 1 0 9 2
10 7 1 9 13 11 7 11 10 9 2
6 10 15 13 1 15 2
7 15 13 10 3 0 9 2
17 10 9 15 11 13 1 2 1 12 2 13 9 2 0 9 2 2
6 15 4 13 1 15 2
8 11 13 1 15 1 1 9 2
8 2 0 13 3 1 10 9 2
12 15 13 0 2 15 13 0 1 3 15 13 2
8 16 15 13 1 7 13 9 2
15 15 13 3 0 9 15 13 0 14 13 16 15 13 15 2
8 15 4 3 13 3 1 9 2
8 13 16 15 13 9 1 15 2
15 15 13 9 1 1 9 7 1 1 9 1 9 7 9 2
15 2 15 13 3 2 7 13 3 2 3 0 1 9 10 2
14 15 4 13 15 3 10 9 13 1 10 9 2 3 2
15 2 16 15 13 1 10 0 9 3 2 10 9 13 1 2
15 2 16 15 13 15 0 16 15 13 3 9 10 13 15 2
5 3 15 13 15 2
5 3 0 15 13 2
11 15 4 13 7 0 7 0 1 9 10 2
8 15 4 15 13 1 0 9 2
7 11 4 13 15 15 3 2
18 2 15 13 10 10 9 14 13 10 9 1 1 14 13 15 1 15 2
4 10 10 9 2
20 15 4 13 0 7 0 1 15 10 2 13 15 1 7 13 3 0 15 13 2
19 15 13 0 13 15 4 13 3 0 0 9 3 16 15 13 15 10 9 2
14 15 13 3 10 9 0 9 2 1 14 13 10 0 2
22 10 9 13 11 10 12 9 1 9 2 1 9 2 1 9 7 1 12 9 1 9 2
18 15 4 13 1 9 7 13 9 2 7 9 12 13 15 0 1 9 2
6 15 13 0 1 9 2
5 13 9 1 9 2
4 13 1 9 2
7 13 14 13 10 0 9 2
10 2 1 0 9 4 15 13 0 9 2
10 3 13 15 1 3 7 13 14 13 2
4 15 13 9 2
4 0 7 0 2
22 7 0 13 15 15 15 3 13 15 2 7 3 13 15 10 7 10 14 13 0 1 2
20 16 15 4 13 15 2 3 13 15 1 2 13 1 15 2 7 3 13 15 2
6 15 13 10 0 9 2
11 10 9 13 10 9 1 9 7 1 9 2
19 15 13 3 7 13 7 13 1 10 9 2 7 9 13 0 1 12 9 2
5 2 15 13 9 2
8 2 15 4 3 13 15 3 2
6 3 13 15 9 2 2
11 10 9 4 13 15 14 13 0 1 10 2
11 3 13 15 1 11 10 0 9 13 1 2
9 15 13 1 10 9 3 1 9 2
6 13 15 0 1 11 2
8 15 4 3 13 3 0 9 2
15 7 3 10 9 4 13 10 9 15 13 9 1 14 13 2
28 15 4 13 11 9 2 10 9 15 13 9 1 14 13 1 11 10 12 9 15 3 4 13 15 1 10 9 2
3 15 9 2
16 10 0 9 15 4 4 13 16 10 0 9 13 1 11 0 2
10 2 6 2 15 13 3 3 1 15 2
10 15 13 3 16 15 13 1 10 0 2
8 15 13 1 15 1 0 9 2
8 15 13 9 3 1 9 10 2
15 15 13 15 1 9 2 1 9 2 1 9 2 1 9 2
7 9 1 9 2 1 9 2
6 2 15 13 3 0 2
18 16 15 13 10 9 0 1 10 2 4 15 4 13 3 0 1 15 2
15 7 15 13 3 3 15 4 4 13 3 0 15 15 13 2
8 3 1 9 13 9 10 9 2
5 15 13 10 9 2
6 2 11 8 8 2 2
22 2 16 15 13 15 2 3 16 15 13 9 2 13 15 9 9 13 1 10 9 1 2
4 15 13 9 2
6 15 13 0 7 0 2
16 15 13 10 0 9 14 13 10 10 9 4 13 1 10 9 2
5 15 13 1 9 2
13 1 13 11 1 9 15 4 13 1 9 1 9 2
11 9 7 9 1 11 13 15 1 10 9 2
8 10 9 0 13 15 3 3 2
32 7 1 3 14 13 15 1 2 4 15 3 0 3 13 16 15 3 13 1 9 1 9 16 11 13 1 10 0 9 1 11 2
5 2 15 13 0 2
9 15 13 1 9 3 1 15 10 2
9 15 13 10 9 1 10 0 9 2
10 7 15 13 3 7 13 15 0 0 2
6 15 4 3 13 1 2
9 2 4 15 13 15 0 0 9 2
14 2 15 4 1 10 9 13 15 9 1 14 13 9 2
7 15 13 0 9 13 0 2
16 1 10 9 1 9 2 16 15 13 7 13 7 13 0 0 2
28 7 3 10 9 2 3 9 12 1 9 2 13 11 1 15 9 2 0 9 7 9 7 13 15 1 1 9 2
11 3 13 15 0 9 7 3 13 15 3 2
14 3 13 15 2 3 13 15 2 3 13 15 10 9 2
7 1 3 4 15 13 3 2
9 2 15 13 10 0 9 14 13 2
12 2 15 13 10 9 15 13 14 13 1 9 2
3 2 6 2
13 1 10 0 13 3 13 15 14 13 1 1 9 2
7 13 1 10 9 1 9 2
5 10 9 15 13 2
19 15 13 0 1 15 2 7 15 13 0 9 1 14 13 0 1 7 1 2
11 11 13 15 4 13 15 0 14 13 0 2
27 2 7 15 13 0 2 7 10 0 15 13 2 13 14 13 1 10 9 2 10 9 2 3 15 13 0 2
18 16 15 3 13 9 7 9 13 1 9 1 15 2 13 15 1 15 2
11 15 13 1 9 1 9 1 9 1 9 2
6 2 3 13 15 0 2
6 7 15 13 3 0 2
8 11 11 4 3 13 14 13 5
2 11 2
11 3 13 10 0 9 10 13 1 10 0 2
6 2 15 13 0 0 2
20 16 10 0 9 13 0 0 2 13 10 9 1 2 0 1 1 9 2 0 2
8 3 13 15 9 1 9 10 2
15 2 9 13 15 16 15 13 7 16 15 13 1 7 13 2
9 9 13 16 15 0 13 1 9 2
23 16 15 3 4 13 9 1 9 2 13 15 15 1 9 2 11 2 1 11 7 13 9 2
12 3 13 15 3 0 14 13 9 15 15 13 2
10 15 4 13 16 15 13 10 0 9 2
7 15 13 10 0 15 13 2
3 2 6 2
7 15 4 3 13 1 15 2
7 13 3 15 13 10 0 2
7 3 13 10 0 9 1 2
11 2 15 4 13 0 9 7 0 10 9 2
13 3 11 1 9 2 1 0 9 7 3 10 9 2
7 13 3 14 13 1 9 2
22 15 13 0 0 0 9 1 11 2 15 13 0 0 1 15 15 13 0 1 1 11 2
11 9 7 9 13 10 0 9 3 1 11 2
5 10 9 9 13 2
8 2 2 11 2 1 11 11 2
5 3 13 15 3 2
15 2 13 10 9 1 9 1 0 11 1 3 10 9 3 2
8 15 13 0 9 15 13 9 2
16 9 13 10 0 10 1 15 7 15 13 3 1 10 10 9 2
5 15 13 10 9 2
28 2 15 13 0 2 7 13 15 12 9 15 3 4 13 0 2 3 13 15 10 0 9 15 13 11 1 11 2
6 3 13 15 3 3 2
9 10 9 13 15 1 14 13 1 2
11 2 15 13 1 1 11 1 10 9 3 2
9 7 13 3 9 1 14 13 11 2
8 3 13 15 9 1 14 13 2
8 13 15 1 9 16 15 13 2
16 2 15 13 15 2 7 6 2 15 13 0 9 16 15 13 2
11 13 15 1 16 15 3 13 3 0 9 2
16 15 13 14 13 9 2 7 15 13 0 1 10 9 15 13 2
7 15 13 15 1 1 9 2
16 2 13 15 13 0 1 9 15 13 9 1 14 13 10 9 2
18 16 15 3 13 0 2 13 15 9 1 14 13 7 13 3 1 9 2
11 10 9 4 15 13 2 16 15 13 9 2
13 2 3 4 15 13 0 1 9 7 13 10 9 2
5 3 0 13 15 2
4 2 15 13 2
19 1 9 13 15 0 0 2 7 15 13 3 9 16 15 3 13 3 0 2
13 13 14 13 1 0 9 7 9 12 9 1 9 2
6 15 13 15 9 1 2
6 2 0 10 0 9 2
6 13 0 0 7 0 2
12 15 15 13 15 1 1 0 2 4 15 13 2
9 7 15 13 16 15 13 15 0 2
8 15 13 15 1 15 1 9 2
5 2 10 0 9 2
12 10 12 9 13 15 1 16 15 13 14 13 2
13 2 16 15 13 3 2 13 15 9 7 9 10 2
6 15 13 1 12 9 2
19 3 13 15 1 15 11 10 2 16 15 13 10 1 9 2 9 7 9 2
15 10 0 11 9 10 4 13 7 9 10 1 11 11 11 2
8 15 13 10 0 15 13 3 2
10 2 15 13 0 0 1 14 13 9 2
20 9 10 13 3 10 0 3 2 7 15 13 3 1 9 16 15 13 1 9 2
11 15 13 15 10 0 12 9 16 9 13 2
22 2 16 9 13 10 9 9 2 13 15 15 1 7 13 1 15 15 4 13 1 9 2
11 13 0 1 14 13 1 2 11 11 2 5
6 9 13 9 1 11 2
7 9 13 15 15 4 13 2
4 13 1 9 2
8 9 11 11 7 9 11 11 2
2 11 2
21 3 10 9 1 9 13 3 0 1 1 2 11 11 2 9 1 11 11 1 9 2
4 2 11 2 2
19 9 11 11 0 9 13 1 9 1 10 0 11 11 1 2 11 11 2 2
20 10 9 1 11 11 1 9 1 11 11 4 13 10 0 9 1 9 1 0 2
32 16 2 11 11 9 2 3 13 1 1 9 1 11 11 1 11 0 9 2 13 3 9 1 3 15 13 14 13 0 0 0 2
15 10 9 4 15 3 13 1 10 0 0 1 14 13 9 2
4 9 13 1 5
21 10 9 4 13 10 9 0 1 11 2 3 1 11 7 10 0 11 1 11 9 2
21 9 13 15 1 9 1 1 9 2 7 13 1 10 0 15 4 4 13 9 9 2
26 15 15 4 13 1 2 4 3 13 7 13 1 1 9 2 16 10 9 13 15 0 12 9 1 9 2
20 15 13 1 15 0 9 2 7 10 9 15 13 15 11 9 1 9 1 9 2
10 2 10 0 12 9 10 9 13 0 2
13 15 13 3 9 1 10 11 11 7 10 0 13 2
12 7 15 13 3 3 9 4 13 1 10 9 2
10 0 13 9 3 9 7 9 13 3 2
16 15 13 1 11 7 1 11 1 10 9 2 13 9 11 11 2
3 0 9 5
29 9 11 11 13 16 15 4 13 14 13 9 16 10 0 9 13 1 10 9 2 3 13 1 11 0 9 7 9 2
19 2 15 13 0 1 10 0 0 9 9 1 10 9 7 10 0 0 13 2
16 13 1 13 9 10 0 9 2 10 9 15 13 1 10 9 2
19 7 13 15 0 0 1 15 2 13 15 10 9 15 13 0 1 3 9 2
15 15 13 10 9 1 9 9 1 9 2 1 14 4 13 2
25 15 13 3 10 9 1 9 1 9 2 10 3 0 9 1 9 2 9 1 9 2 7 3 0 2
16 15 13 0 9 15 4 13 1 10 9 2 13 11 1 11 2
3 2 0 5
21 9 2 15 4 13 12 0 9 1 9 1 10 0 9 2 4 3 0 13 9 2
11 2 13 1 0 9 7 13 10 0 9 2
20 0 0 2 15 13 15 1 10 9 15 4 13 0 9 7 0 9 1 9 2
22 15 13 0 0 1 16 15 4 13 10 10 9 2 13 10 0 0 11 11 1 11 2
15 11 13 3 1 9 7 9 2 7 13 10 9 1 9 2
17 2 15 13 0 0 1 9 14 13 15 10 2 7 0 7 0 2
19 15 13 3 15 13 0 16 15 13 0 9 7 13 15 1 10 10 9 2
14 15 13 3 3 9 2 13 15 1 9 2 7 13 2
25 2 16 15 4 13 10 9 10 9 15 10 13 0 2 4 15 13 1 16 15 13 3 0 1 2
16 7 1 9 4 15 4 4 13 1 16 15 4 13 15 10 2
17 15 13 0 1 9 16 15 4 13 1 1 10 9 1 0 9 2
6 1 10 9 1 9 5
14 11 4 13 0 1 14 13 1 9 1 9 1 11 2
28 15 4 3 13 1 15 10 0 0 1 9 7 13 0 9 1 0 2 16 10 0 4 4 13 0 1 9 2
13 11 4 13 1 11 2 15 3 4 13 10 9 2
21 15 13 10 1 10 0 15 4 13 15 14 13 1 1 9 1 9 10 0 9 2
20 2 2 11 11 2 13 10 9 15 13 9 1 14 13 16 15 13 0 15 2
19 1 9 13 15 15 1 10 9 2 7 3 13 10 0 9 1 1 15 2
8 15 13 0 10 0 9 3 2
26 9 11 13 16 15 13 9 15 13 1 9 10 0 9 16 15 13 15 9 1 2 11 11 9 2 2
11 2 15 13 10 0 1 14 13 10 9 2
24 15 13 15 0 15 15 13 15 4 13 1 1 2 7 15 13 9 1 14 13 15 1 3 2
32 15 13 9 1 14 13 3 1 15 2 7 10 0 9 2 7 16 0 13 14 13 3 1 15 4 15 0 13 2 13 11 2
6 2 13 9 10 9 5
28 2 9 15 13 16 15 13 1 11 1 9 2 13 15 16 10 0 3 13 3 1 9 15 3 13 15 1 2
21 15 4 13 3 0 14 13 3 2 1 16 15 13 0 1 14 13 15 1 9 2
15 1 10 9 13 15 14 13 9 10 9 2 13 11 0 2
21 1 1 11 13 15 1 11 0 1 10 9 9 2 7 3 15 13 7 13 9 2
21 2 15 4 13 14 13 15 1 3 10 0 0 2 7 3 4 15 4 13 1 2
36 15 13 3 3 16 15 1 9 3 13 9 1 10 9 2 15 13 10 10 15 13 1 15 2 7 15 4 3 3 13 10 9 15 13 15 2
15 16 15 13 10 9 2 13 15 0 1 9 2 13 11 2
18 2 13 15 0 1 15 14 13 1 2 11 11 9 2 9 1 11 2
21 2 14 13 1 10 10 9 13 10 0 0 9 2 16 15 4 13 9 14 13 2
19 7 15 4 13 0 2 3 15 13 13 4 15 10 9 0 1 15 3 2
5 3 13 15 9 5
12 15 13 0 1 9 11 11 7 9 11 11 2
6 3 4 15 3 13 2
8 13 14 13 9 1 11 11 2
14 1 0 9 1 11 13 10 10 10 12 9 7 9 2
5 10 0 9 13 2
10 7 15 13 1 9 1 9 1 9 2
5 3 3 1 9 2
19 9 11 11 13 9 1 14 13 11 0 9 3 15 13 9 1 10 0 2
28 3 0 2 1 10 10 9 1 9 2 13 9 11 11 9 1 14 13 2 11 2 2 11 11 7 11 11 2
4 1 0 9 5
17 7 4 15 3 3 13 15 3 2 3 4 15 3 13 3 0 2
38 2 15 13 1 9 1 9 1 9 1 9 2 7 3 13 15 1 9 14 13 1 9 2 13 11 11 2 13 1 10 12 9 1 9 11 7 11 2
9 9 1 11 9 1 11 13 0 2
25 2 15 13 1 15 15 13 10 12 15 13 16 15 13 1 14 13 2 13 9 11 11 7 13 2
26 1 9 13 15 7 9 1 11 9 1 11 9 1 12 9 2 1 9 1 9 13 15 3 3 0 2
20 11 11 13 2 1 10 0 10 9 2 0 9 0 15 15 13 15 1 9 2
24 2 15 13 1 9 2 7 15 13 9 2 13 11 2 15 3 13 10 1 9 9 1 9 2
14 7 15 13 15 13 0 0 14 13 14 13 9 3 2
5 15 13 3 9 5
6 15 13 11 11 3 2
28 15 13 3 0 0 9 1 15 7 15 7 11 11 16 15 4 13 1 1 9 2 1 9 9 7 0 9 2
14 3 13 15 15 3 13 10 9 9 14 13 9 3 2
30 2 15 13 10 9 9 15 4 13 1 2 1 14 13 9 0 9 2 13 11 2 7 13 1 9 15 13 9 9 2
15 2 16 15 13 0 9 13 15 3 0 2 13 15 0 2
11 1 11 13 15 3 0 14 13 1 9 2
11 2 3 12 1 12 15 13 3 13 9 2
19 10 0 9 13 0 0 1 10 3 0 9 2 1 9 2 13 11 11 2
4 7 13 1 2
8 1 9 1 10 10 0 9 2
7 7 1 10 0 9 1 2
8 2 3 13 15 0 1 9 2
23 16 15 13 3 0 1 1 10 9 7 9 7 3 2 13 10 0 0 11 11 1 11 2
3 13 3 2
10 15 13 10 9 0 1 9 1 9 5
15 2 15 4 13 1 9 16 9 3 13 0 1 12 9 5
16 3 4 0 9 13 1 1 0 9 2 13 9 11 1 11 2
9 13 14 13 10 0 9 1 9 2
16 11 11 1 11 13 10 0 1 14 13 9 7 10 0 9 2
24 7 0 0 0 9 13 3 9 1 9 2 16 9 3 13 16 15 4 4 13 1 10 9 2
2 9 2
7 11 11 5 11 5 11 5
5 2 15 13 0 2
13 16 11 13 9 1 15 2 4 15 4 0 13 2
22 15 13 3 3 9 1 10 9 14 13 9 1 0 9 2 13 11 11 2 12 2 2
12 15 13 3 1 9 7 10 0 9 1 11 2
20 12 9 0 11 13 3 1 1 9 1 11 2 16 10 0 9 13 1 9 2
6 2 9 10 4 13 2
14 15 13 1 9 2 7 15 1 9 1 9 13 1 2
8 10 0 9 13 15 1 9 2
14 7 15 13 1 15 9 2 9 7 9 1 9 10 2
17 9 10 13 15 0 1 9 2 16 15 4 13 16 15 13 9 2
7 3 13 15 15 1 9 2
21 7 15 13 0 9 0 0 1 16 11 4 13 15 7 13 1 15 2 13 11 2
9 10 11 13 10 0 9 10 9 2
13 1 10 0 9 2 13 11 7 9 0 1 3 2
12 2 15 4 3 13 3 0 7 3 7 3 2
13 7 10 9 13 15 9 10 16 15 4 13 9 2
7 11 13 9 2 13 9 2
9 1 9 13 11 9 1 11 11 2
11 15 4 3 13 1 1 0 1 12 9 2
24 11 13 15 1 11 1 11 2 15 1 9 1 9 1 11 7 11 13 9 1 10 0 9 2
13 2 16 11 4 13 1 9 2 13 15 9 10 2
14 1 12 9 1 0 11 2 13 15 3 1 1 12 2
20 15 13 0 2 7 3 0 3 1 10 9 1 1 12 9 9 2 13 15 2
18 1 11 7 11 13 0 9 1 9 12 9 2 10 0 9 1 11 2
15 2 0 13 15 0 14 13 0 9 7 13 1 10 9 2
8 3 0 9 2 3 0 9 2
18 1 11 9 2 4 9 13 16 15 13 0 0 14 13 3 0 9 2
16 7 3 13 15 10 0 9 1 9 2 1 9 1 11 11 2
12 10 0 1 10 9 4 4 13 2 13 11 2
12 2 1 9 13 15 9 0 9 1 0 9 2
13 15 4 13 16 1 12 12 9 2 13 12 9 2
11 15 13 16 10 0 9 13 10 0 9 2
34 2 10 0 9 13 3 7 0 0 9 2 1 16 9 0 3 4 13 10 0 9 7 9 14 13 0 9 1 0 9 2 13 11 2
7 2 11 13 3 10 9 2
13 9 4 3 3 13 3 1 14 4 13 10 9 2
24 9 13 3 9 3 2 7 1 10 0 9 13 9 3 0 1 12 9 1 9 2 13 9 2
25 2 16 10 0 9 13 1 14 4 13 15 1 9 10 2 3 13 10 0 0 9 9 1 9 2
24 15 4 13 1 9 16 9 3 13 0 1 12 9 2 16 9 13 1 9 9 2 13 15 2
11 10 10 9 13 16 15 13 0 1 9 2
17 12 9 1 9 13 1 9 2 7 0 9 13 0 0 9 1 2
5 11 13 3 0 2
21 15 13 1 16 1 10 12 9 1 11 3 2 3 13 9 1 9 15 13 1 2
19 2 9 4 3 4 13 1 0 1 10 0 9 2 7 15 13 10 10 2
8 3 4 0 0 9 13 9 2
23 10 0 9 13 3 1 9 1 9 2 7 15 13 9 9 1 9 1 9 7 9 9 2
7 2 9 13 3 9 9 2
19 10 0 9 13 0 9 7 9 2 7 3 13 15 0 9 2 13 11 2
13 2 1 7 1 4 15 3 13 16 15 13 9 2
17 3 0 15 4 13 2 4 9 1 11 13 0 2 13 15 1 2
17 9 1 11 13 10 0 9 1 10 0 9 2 7 10 0 9 2
20 2 15 13 1 7 1 0 1 15 16 15 13 2 7 15 13 15 13 0 2
11 15 4 3 13 14 13 15 2 13 11 2
5 7 0 13 15 2
13 11 13 1 1 0 11 1 14 13 3 9 13 2
15 15 13 3 10 0 9 1 1 2 3 11 3 13 9 2
16 2 15 4 13 15 4 4 13 9 10 9 1 9 1 9 2
22 4 15 13 2 13 15 3 16 15 13 1 10 0 9 2 7 16 15 13 1 9 2
7 15 13 15 2 13 11 2
21 2 10 9 13 15 3 1 9 10 1 11 1 1 2 3 15 4 13 12 9 2
7 9 3 1 13 3 0 2
10 3 10 9 13 1 16 15 4 13 2
17 15 13 3 1 12 9 2 7 10 9 13 15 1 1 0 9 2
15 12 9 7 10 9 4 13 7 13 16 15 13 3 1 2
16 2 0 13 15 3 0 15 13 0 1 16 15 0 13 9 2
9 15 13 1 9 2 9 7 9 2
7 15 13 0 1 0 9 2
15 1 0 9 13 11 3 1 9 1 9 10 1 1 11 2
19 2 15 13 3 1 16 15 13 1 15 9 2 7 1 15 15 4 13 2
7 1 15 15 13 9 10 2
6 16 15 13 9 10 2
11 3 13 15 15 16 15 4 13 1 9 2
14 10 9 4 13 1 11 9 2 7 3 13 1 9 2
13 13 15 9 7 9 2 13 15 1 15 1 9 2
9 3 4 11 2 12 2 13 1 5
6 13 9 1 10 9 2
3 13 9 2
13 9 11 11 13 11 9 1 3 14 13 10 9 2
12 0 9 1 9 4 13 10 9 1 9 10 2
23 11 4 13 10 0 9 1 9 16 15 13 12 9 2 7 13 0 1 14 13 1 9 2
19 2 15 4 13 1 14 13 10 9 2 13 9 11 11 1 11 1 11 2
30 9 1 10 0 9 11 11 4 13 9 1 1 16 15 13 7 9 7 10 0 9 1 14 13 15 13 10 0 9 2
15 0 9 1 0 9 1 9 4 13 10 9 1 9 10 2
34 11 0 9 13 14 4 13 10 0 9 3 1 9 7 10 12 9 1 9 7 9 2 1 14 4 13 1 7 1 1 9 0 9 2
39 2 16 15 13 16 10 9 13 1 9 1 14 13 10 10 9 13 15 7 1 9 9 7 9 2 7 13 3 9 9 1 1 9 2 13 11 1 11 2
3 13 3 5
19 11 13 3 9 1 14 13 9 1 9 2 7 9 13 14 13 9 9 2
23 3 13 10 0 9 1 11 1 14 13 1 9 1 14 13 10 0 9 1 14 13 9 2
10 15 13 3 1 14 13 15 1 9 2
22 2 11 13 10 9 3 2 3 1 10 0 2 1 1 1 16 15 3 13 12 9 2
8 7 15 4 13 0 1 9 2
13 15 13 14 3 13 15 3 0 1 1 10 9 2
34 15 13 15 1 9 15 4 13 15 1 2 7 3 15 4 13 1 9 2 7 15 4 13 14 13 15 2 13 11 9 2 11 11 2
15 1 16 10 9 1 9 13 9 1 11 13 9 14 13 2
8 3 13 11 9 14 13 1 2
14 9 13 0 1 16 15 3 13 12 9 3 14 13 2
5 2 15 13 0 5
7 2 15 13 10 0 9 2
6 15 13 0 0 9 2
10 1 10 9 4 15 13 0 1 15 2
36 15 13 0 1 9 14 13 16 15 4 13 2 7 15 13 3 15 15 13 0 1 15 2 13 11 11 1 10 9 1 10 0 9 11 11 2
33 15 13 16 9 4 3 13 15 1 14 13 10 9 2 7 16 15 13 10 10 9 4 15 13 3 1 14 13 10 13 1 15 2
15 2 15 13 10 0 9 2 7 9 13 15 3 0 9 2
8 15 4 13 3 9 1 9 2
20 3 4 15 3 13 1 2 3 16 15 13 16 9 10 13 0 2 13 11 2
22 11 9 13 10 0 0 0 9 2 3 16 15 13 10 9 14 13 9 1 14 13 2
13 7 3 9 13 1 14 13 1 10 9 7 9 2
5 4 3 13 15 5
15 9 13 3 9 0 1 16 11 4 13 1 14 13 15 2
28 2 15 13 10 9 14 13 15 3 1 3 2 7 15 4 7 9 7 0 9 13 0 1 2 13 11 11 2
22 11 9 13 10 0 0 0 9 2 3 16 15 13 10 9 14 13 9 1 14 13 2
13 7 3 9 13 1 14 13 1 10 9 7 9 2
35 9 1 10 0 9 1 10 0 9 2 11 11 2 13 16 10 9 1 11 9 13 1 9 1 14 13 10 10 9 13 1 10 0 9 2
29 15 13 3 1 10 9 1 10 0 9 15 13 16 10 9 15 13 7 9 7 9 4 13 14 13 1 0 0 2
6 4 3 13 1 11 5
20 10 1 11 0 9 13 14 4 13 1 11 11 1 11 3 1 9 1 9 2
26 15 4 13 15 14 13 0 16 10 9 4 4 13 9 1 9 1 11 9 2 13 1 10 11 11 2
25 11 9 11 2 15 13 9 2 4 13 16 15 13 9 4 13 10 7 0 9 1 14 13 15 2
17 1 9 4 3 9 13 1 11 2 1 9 15 4 13 1 11 2
19 9 4 13 1 10 0 9 2 7 4 0 13 1 9 1 0 0 9 2
22 10 9 1 0 2 9 7 9 4 13 14 13 1 1 9 1 14 13 11 7 9 2
24 2 16 15 4 13 1 9 13 15 1 9 2 7 1 3 4 15 13 0 1 9 1 9 2
12 15 4 3 13 16 15 4 13 1 15 3 2
24 15 15 13 3 0 13 16 10 0 9 3 10 9 13 15 9 13 2 13 11 9 2 11 2
21 11 13 12 0 9 2 11 2 12 2 2 11 2 12 2 7 11 2 12 2 2
23 2 0 9 4 13 1 1 15 16 0 9 10 4 4 13 1 11 0 9 2 13 9 2
3 0 9 5
17 1 12 13 0 9 10 0 9 2 15 3 13 1 9 11 11 2
7 9 13 3 1 10 0 2
13 9 13 1 10 12 9 0 9 15 3 13 9 2
17 15 13 3 14 13 2 7 15 4 3 13 1 10 10 9 9 2
14 15 13 3 3 14 13 10 0 9 2 13 11 11 2
12 1 0 9 13 9 1 9 16 9 4 13 2
10 9 13 16 15 13 1 9 10 0 2
7 9 13 0 9 1 11 2
4 13 10 9 5
12 11 11 1 9 2 0 9 7 9 15 13 2
2 9 2
11 0 9 1 9 13 11 9 1 0 9 2
13 3 13 15 7 9 11 11 11 3 1 11 11 2
2 11 2
14 1 9 1 11 11 1 12 2 13 15 9 1 9 2
16 11 13 9 2 13 9 1 9 7 4 13 1 11 11 11 2
3 0 9 2
7 1 9 1 11 11 11 2
12 15 13 15 15 4 13 1 10 0 12 9 2
11 15 13 1 1 11 11 11 1 9 9 2
54 2 15 13 0 14 13 1 9 1 14 4 13 1 15 2 13 15 2 4 13 1 15 2 13 15 2 4 13 1 15 2 1 16 15 4 13 9 10 1 10 9 2 7 3 13 15 10 0 9 2 13 11 11 2
7 2 7 3 13 15 3 2
6 2 2 13 15 1 2
3 2 6 2
10 3 15 13 1 11 11 2 13 15 2
38 15 13 3 2 1 9 1 11 11 11 1 11 11 7 13 1 14 13 1 9 2 7 15 13 0 9 15 4 13 15 1 1 10 0 2 0 9 2
12 15 13 15 15 4 13 1 10 0 12 9 2
7 15 13 3 15 4 13 2
30 7 16 11 13 10 0 9 7 13 1 11 1 12 2 13 15 3 16 15 4 13 1 0 9 1 9 1 9 10 2
15 15 13 3 16 10 0 9 10 13 1 9 1 14 13 2
12 11 13 1 11 11 1 14 13 0 1 9 2
12 15 13 3 1 1 11 11 11 1 9 9 2
13 2 3 13 15 0 14 13 1 11 2 13 11 2
11 2 15 13 14 13 1 1 10 0 9 2
9 7 15 13 10 9 14 13 3 2
18 15 13 15 13 1 1 9 2 1 15 15 0 13 14 13 1 1 2
7 15 13 3 0 1 11 2
21 15 13 3 3 0 14 13 1 3 2 7 15 13 15 1 1 0 9 0 9 2
27 15 4 13 1 10 9 16 15 13 12 2 7 15 13 0 14 4 13 10 0 9 2 10 9 2 3 2
17 1 11 4 15 13 1 10 0 9 10 2 2 11 11 11 2 2
21 15 13 1 9 2 11 2 15 13 1 9 1 0 9 7 15 13 1 1 9 2
12 15 4 13 15 1 15 15 13 2 9 2 2
5 15 4 13 9 2
4 13 15 3 2
28 7 3 4 9 15 13 11 11 7 13 9 10 1 0 11 2 1 10 9 13 10 9 1 9 9 7 9 2
21 3 1 11 11 4 15 13 10 10 12 9 1 9 2 10 9 2 9 7 9 2
28 9 2 11 11 2 13 11 1 10 2 0 7 0 9 1 9 7 9 15 13 10 9 1 9 1 9 2 2
33 15 4 13 7 13 2 1 9 2 1 9 2 1 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2
3 7 9 2
8 2 9 1 9 2 13 11 2
9 2 3 2 9 1 9 1 9 2
6 15 13 3 10 9 2
6 15 4 3 13 9 2
13 15 4 1 10 9 3 13 1 16 15 13 9 2
14 2 4 15 13 1 9 1 3 15 13 14 13 9 2
3 2 6 2
4 15 13 15 2
6 7 15 13 3 0 2
12 15 13 3 0 9 15 13 0 14 13 1 2
11 9 1 0 7 0 9 4 13 1 9 2
14 0 9 4 13 1 14 13 3 0 2 3 1 9 2
10 15 4 13 16 9 4 13 0 0 2
11 9 13 15 9 3 1 0 13 9 1 2
9 3 13 2 11 2 10 0 9 2
14 9 7 10 9 1 10 9 7 9 1 10 0 13 2
20 1 9 4 7 11 11 7 15 13 0 10 10 12 9 1 10 9 1 9 2
9 2 15 4 13 16 9 13 0 2
16 15 4 3 13 1 14 13 15 15 3 13 15 2 13 11 2
12 2 15 13 3 0 16 9 13 10 0 9 2
5 15 13 3 0 2
5 15 13 0 9 2
9 2 15 13 15 3 0 1 9 2
43 1 1 15 15 13 1 9 3 3 2 13 15 1 9 1 10 0 7 0 9 1 9 1 10 9 2 2 13 11 1 9 1 9 11 11 1 12 2 16 15 13 1 2
7 2 13 1 10 9 2 2
9 2 15 13 9 1 9 1 0 2
10 15 13 10 9 9 15 13 0 0 2
13 15 13 0 1 14 13 0 1 9 2 13 15 2
13 15 4 13 1 9 7 9 1 9 2 3 9 2
28 15 13 0 1 15 15 13 1 9 2 7 15 13 15 1 3 16 15 13 9 16 0 9 4 4 13 9 2
11 9 13 3 0 16 10 12 9 4 13 2
10 2 13 15 15 1 9 15 3 13 2
7 2 15 13 3 9 10 2
22 15 13 15 1 9 2 15 13 3 9 10 2 13 0 2 13 1 9 16 9 13 2
6 7 15 13 1 15 2
10 7 15 13 15 15 4 13 1 9 2
8 10 9 15 13 15 1 9 2
7 9 4 3 13 9 0 2
8 15 4 13 0 0 1 15 2
5 9 13 3 9 2
7 0 1 10 3 0 9 2
16 15 4 13 0 9 1 9 15 13 1 10 9 2 1 9 2
6 15 4 13 15 1 2
10 2 10 0 9 13 15 10 9 0 2
6 3 13 15 3 0 2
7 9 4 13 2 9 13 2
3 9 13 2
28 10 9 15 13 0 1 9 0 1 11 9 10 0 9 2 15 13 15 2 2 13 11 1 9 2 11 2 2
6 15 13 1 15 10 2
13 1 16 15 4 13 1 10 0 9 1 12 9 2
13 2 15 4 13 15 1 16 15 3 13 9 0 2
11 7 16 15 13 3 0 10 9 14 13 2
24 15 13 3 15 10 9 16 15 13 10 9 2 7 15 13 15 10 9 16 15 13 10 9 2
15 2 13 15 3 15 13 0 1 9 1 0 9 14 13 2
27 2 6 2 7 15 13 16 15 4 13 15 1 14 13 1 1 15 2 3 16 15 13 15 7 13 9 2
9 15 4 13 9 1 10 10 9 2
11 15 13 3 1 9 3 2 1 10 9 2
21 15 4 13 7 13 16 15 13 10 9 16 15 13 1 10 0 9 1 12 9 2
9 3 4 15 13 15 1 0 9 2
21 7 9 13 0 14 13 2 13 15 2 10 0 13 16 15 13 0 2 7 0 2
9 15 13 15 13 0 16 9 13 2
13 7 15 13 2 3 0 0 2 16 9 13 0 2
10 2 15 13 3 3 16 9 13 0 2
9 15 4 3 13 15 1 14 13 2
7 15 13 0 1 0 9 2
28 15 13 0 14 13 1 9 2 7 15 4 13 3 1 10 9 1 9 2 6 2 7 15 4 3 13 0 2
13 15 4 3 3 13 15 2 15 13 15 0 0 2
7 11 13 15 1 10 9 2
4 2 3 3 2
22 2 15 13 1 9 1 15 1 11 11 2 13 10 9 2 7 13 15 1 11 11 2
13 15 0 13 2 0 13 1 9 1 9 1 11 2
23 15 13 0 1 13 2 13 0 2 0 2 0 16 15 13 1 9 15 3 4 13 9 2
15 15 13 3 9 16 11 11 4 13 3 1 10 9 0 2
16 9 13 14 13 9 2 13 1 9 2 13 0 1 9 10 2
7 2 7 3 13 15 9 2
12 7 15 13 0 2 9 1 0 9 7 15 2
37 1 10 9 1 10 0 9 1 11 2 1 12 9 1 16 15 4 13 15 1 10 9 1 11 2 13 11 15 1 10 12 9 0 9 11 11 2
8 2 15 13 10 0 0 9 2
10 7 15 13 3 0 14 3 13 15 2
5 3 0 2 3 2
9 15 13 9 1 0 9 2 15 2
5 15 13 0 0 2
21 15 13 1 14 13 12 9 3 2 7 0 7 0 7 0 3 2 6 2 0 2
5 0 2 0 0 2
11 2 4 15 13 1 9 1 0 9 1 2
3 2 3 2
5 7 15 13 15 2
7 15 13 15 2 10 12 2
28 15 13 0 10 9 15 13 1 9 2 9 7 15 15 3 13 2 7 15 13 3 14 13 9 1 9 0 2
5 15 13 3 3 2
2 6 2
4 15 13 15 2
8 2 15 13 15 1 10 9 2
5 2 1 10 9 2
8 15 13 3 0 10 9 0 2
7 15 13 3 15 3 3 2
5 15 3 13 15 2
10 7 1 0 9 13 15 15 1 15 2
27 7 3 13 15 3 2 6 2 3 13 15 1 1 9 3 1 9 2 13 15 10 0 9 7 3 2 2
18 15 13 3 3 9 1 10 10 1 16 15 4 13 3 1 3 1 2
5 2 13 15 0 2
13 2 6 2 7 15 13 3 9 1 10 0 13 2
16 7 15 13 9 2 7 15 13 9 7 10 9 1 10 9 2
9 11 1 11 2 0 9 1 9 2
30 11 13 9 13 10 0 9 1 9 1 10 9 1 12 9 1 9 2 16 9 3 4 13 1 9 9 12 1 9 2
11 15 13 0 9 9 11 4 13 1 9 2
9 7 15 13 10 9 11 13 15 2
18 15 13 9 1 9 11 11 1 12 9 2 15 4 13 11 0 9 2
9 7 15 13 9 10 3 1 12 2
15 16 15 13 1 11 11 1 12 2 13 10 12 1 15 2
11 2 15 13 15 3 1 2 0 7 0 2
33 11 4 13 0 0 1 15 2 7 15 13 1 15 16 15 4 13 3 9 1 9 2 7 15 13 1 10 9 16 15 3 13 2
19 15 13 1 14 13 1 10 0 9 2 16 15 13 0 7 0 1 15 2
5 15 13 0 0 2
14 15 13 1 1 10 9 15 15 3 13 4 13 1 2
19 15 13 1 10 9 3 15 4 13 15 3 2 7 15 13 15 10 3 2
4 3 13 15 2
6 15 13 1 10 9 2
8 2 15 13 1 9 1 9 2
17 7 15 13 15 0 0 14 13 1 16 15 4 13 3 1 9 2
20 0 4 15 4 13 1 1 2 3 3 1 10 0 2 7 3 1 10 0 2
10 2 13 15 0 1 15 14 13 0 2
8 2 6 2 15 13 3 15 2
7 7 15 13 3 0 3 2
8 15 9 13 15 15 13 3 2
8 15 13 3 0 14 13 15 2
5 7 15 13 0 2
7 15 13 0 7 0 0 2
7 15 13 11 11 11 3 2
6 15 13 11 11 11 2
23 10 9 10 13 1 9 1 11 2 7 11 13 1 9 1 11 11 1 9 1 10 9 2
7 2 13 15 10 0 9 2
7 2 15 4 11 13 1 2
5 2 15 13 9 2
4 2 13 15 2
5 3 0 2 3 2
7 2 3 13 15 15 0 2
26 2 16 15 13 14 13 15 1 10 0 2 7 15 13 15 15 13 1 1 14 13 9 1 10 10 2
20 14 13 9 1 16 15 13 0 2 16 15 3 4 13 15 2 15 3 13 2
9 15 4 13 10 9 1 10 9 2
14 7 15 13 3 9 1 16 15 13 15 2 13 11 2
16 2 7 15 13 3 1 9 7 9 16 15 3 4 13 15 2
13 11 7 11 4 13 16 15 13 10 9 1 9 2
13 3 13 15 15 16 15 3 13 10 9 1 9 2
12 15 4 13 3 2 0 0 2 13 2 13 2
14 0 13 15 9 2 13 1 7 13 0 3 1 9 2
4 11 13 3 2
10 15 13 3 0 1 9 1 10 9 2
9 15 13 3 3 9 1 1 9 2
9 2 15 4 13 15 2 13 15 2
13 15 13 9 2 7 9 13 1 16 15 13 1 2
5 11 13 1 9 2
12 2 15 13 1 10 9 3 0 2 13 15 2
23 2 16 15 3 13 15 2 13 15 3 9 3 2 15 13 11 9 14 13 10 9 1 2
5 7 3 13 15 2
8 2 6 2 15 4 13 9 2
11 15 4 3 13 10 9 1 1 9 2 2
46 1 16 11 11 13 11 11 1 11 1 11 1 12 2 13 15 3 0 9 16 15 4 13 1 14 13 9 7 9 1 9 7 1 10 9 2 16 15 13 9 1 0 9 1 9 2
29 1 16 15 13 9 1 9 1 9 1 11 1 12 2 13 0 9 1 11 15 10 9 1 10 0 9 1 11 2
23 15 4 13 1 9 9 7 15 13 12 9 16 9 10 4 13 16 15 13 0 1 15 2
6 2 15 13 0 0 2
8 7 15 13 0 14 13 3 2
19 7 15 16 15 13 15 2 13 10 0 0 9 1 15 15 3 4 13 2
13 15 4 13 0 1 9 1 10 9 2 13 15 2
6 9 3 3 1 9 2
31 15 4 3 13 1 1 10 0 9 2 7 15 13 0 9 1 9 10 2 3 1 16 15 13 1 11 7 9 1 9 2
10 15 4 13 16 15 3 4 13 15 2
23 16 10 9 4 13 0 1 15 1 14 13 10 9 2 3 16 15 1 9 4 13 0 2
15 2 15 4 13 0 1 15 2 7 15 13 0 10 9 2
5 15 4 9 13 2
10 9 13 9 16 9 3 13 1 9 2
16 9 7 9 11 11 4 13 1 2 9 2 1 9 1 11 2
20 15 13 10 0 9 2 3 13 15 0 14 13 16 15 13 9 1 10 9 2
11 15 13 9 15 4 13 16 9 13 1 2
17 15 13 10 9 14 13 9 1 2 15 13 0 0 1 0 9 2
13 2 13 15 1 10 9 16 15 4 13 0 0 2
3 2 6 2
6 15 13 3 1 15 2
11 3 16 15 4 13 15 7 9 10 0 2
13 10 0 9 10 13 1 9 1 9 10 2 13 2
10 2 13 16 15 3 13 10 9 2 2
12 10 9 13 15 0 1 14 13 1 15 0 2
7 7 13 1 9 1 9 2
7 7 1 9 13 15 0 2
4 3 1 9 2
5 15 13 10 9 2
6 2 0 9 2 0 2
12 0 0 13 9 14 13 9 1 9 7 13 2
17 15 13 10 0 0 9 15 4 13 2 7 15 13 15 0 1 2
12 15 13 1 14 13 0 16 15 13 12 9 2
10 7 3 15 13 15 3 2 6 6 2
11 2 15 13 3 15 15 4 13 13 0 2
11 15 13 3 9 15 4 13 15 13 0 2
5 7 15 13 9 2
4 14 13 9 2
14 15 13 16 15 15 4 13 13 1 9 1 10 9 2
23 7 15 4 13 0 2 15 4 13 15 0 2 7 15 4 13 0 9 3 2 13 11 2
12 2 15 13 3 0 16 15 13 3 0 9 2
4 15 13 9 2
9 15 13 14 3 4 13 1 9 2
10 7 9 13 0 9 9 1 15 9 2
10 15 13 3 15 16 15 4 13 0 2
7 7 15 13 3 1 9 2
17 16 9 13 1 9 1 10 0 9 2 3 13 15 2 13 11 2
15 15 13 12 9 7 13 1 9 1 9 11 11 1 11 2
3 9 13 2
6 11 13 15 3 1 2
17 3 12 9 1 13 15 10 9 1 9 1 0 9 1 9 10 2
14 15 13 9 7 9 2 7 15 13 0 9 1 9 2
13 15 4 13 14 13 9 10 1 0 9 1 11 2
13 15 13 14 13 9 1 12 9 1 9 1 9 2
18 2 15 13 3 3 0 1 14 13 0 0 2 1 14 13 15 3 2
20 7 15 4 13 0 2 15 13 1 9 0 2 15 4 13 9 1 15 3 2
9 15 4 13 0 0 7 0 0 2
14 3 13 4 15 3 13 16 15 4 13 0 0 3 2
11 3 10 2 3 13 15 13 2 9 0 2
26 7 15 4 13 1 10 0 9 2 13 15 1 0 2 13 1 9 2 13 10 9 7 13 0 3 2
8 15 4 13 15 9 1 9 2
14 3 4 9 15 9 13 2 11 0 9 2 13 9 2
5 3 1 10 9 2
15 2 7 15 13 3 3 16 15 13 9 1 9 2 3 2
8 15 13 15 4 13 0 0 2
11 15 4 13 15 4 13 12 2 13 11 2
7 2 15 9 9 13 15 2
33 2 10 9 16 15 13 1 9 13 10 10 9 2 15 15 13 9 7 13 2 13 7 13 1 14 13 15 10 7 10 10 9 2
13 9 10 4 3 13 9 7 0 2 7 0 9 2
20 15 13 3 0 1 16 9 4 13 15 10 7 13 9 1 14 13 10 9 2
13 15 4 3 13 10 0 10 2 10 0 0 9 2
24 12 9 0 11 2 11 0 9 1 10 0 9 2 13 3 1 9 3 1 9 2 11 2 2
13 2 15 4 13 0 1 16 10 9 3 4 13 2
23 15 13 3 9 1 10 10 9 3 2 7 15 14 4 13 1 15 2 13 15 13 0 2
18 15 13 9 2 7 15 13 3 10 0 9 1 9 9 1 0 9 2
15 15 13 1 10 9 16 15 13 10 9 15 3 13 1 2
5 2 1 15 3 2
7 2 9 2 3 7 0 2
9 15 4 3 13 15 3 0 1 2
15 0 13 15 3 3 10 0 9 1 2 15 1 15 2 2
20 15 13 10 9 15 13 10 10 9 1 9 10 2 15 3 4 13 1 15 2
16 15 4 15 13 7 13 1 16 15 4 13 10 9 1 9 2
11 11 4 13 1 1 11 16 15 13 9 2
10 7 15 13 3 10 0 9 3 1 2
25 2 16 15 13 15 14 13 2 3 13 15 9 1 2 7 3 13 15 15 0 1 2 13 11 2
16 2 16 15 3 13 15 14 13 2 13 15 0 10 14 13 2
17 15 4 13 9 2 13 1 15 2 11 2 9 15 13 1 15 2
26 3 13 11 11 3 2 1 9 1 11 2 1 10 0 0 9 7 13 1 14 13 0 9 1 11 2
37 15 13 1 10 9 2 10 10 0 9 15 4 4 13 1 15 2 9 15 4 13 2 7 15 13 3 16 9 4 13 1 14 13 9 1 9 2
29 2 10 9 13 15 2 9 2 7 13 16 10 0 0 9 1 9 10 4 13 15 1 14 13 9 2 13 11 2
14 15 13 10 0 0 9 2 13 1 9 2 13 1 2
8 2 15 13 15 0 0 1 2
8 7 3 4 15 13 14 13 2
7 11 13 1 3 12 0 5
12 11 13 1 0 12 0 1 11 7 1 11 2
24 9 11 11 13 16 12 0 1 11 4 13 1 1 11 11 2 15 13 9 7 9 1 9 2
16 12 1 10 9 13 1 11 2 12 1 11 7 12 1 11 2
8 12 0 4 13 1 1 11 2
16 1 9 4 10 0 9 9 7 10 0 0 13 9 1 9 2
19 11 4 0 13 9 1 0 12 0 1 9 7 10 9 1 11 7 11 2
21 2 15 4 13 10 0 9 1 1 9 7 13 15 1 10 1 14 13 9 0 2
25 15 13 16 15 13 12 0 1 9 2 7 15 13 3 3 2 13 9 11 11 1 9 1 11 2
8 2 0 9 13 10 0 9 5
7 11 13 2 11 11 2 2
2 9 2
13 11 0 9 11 11 4 13 1 1 9 1 9 2
35 15 4 13 9 10 9 1 16 11 4 13 15 1 10 10 9 1 14 13 1 2 11 11 2 2 7 3 4 9 0 13 10 0 9 2
21 2 11 11 11 2 13 10 10 9 15 4 13 14 13 9 1 7 13 1 9 2
3 0 9 5
27 11 4 13 1 0 9 7 11 9 11 11 2 15 13 9 13 10 0 9 7 9 1 2 11 11 2 2
8 2 15 13 10 0 10 9 2
32 15 13 0 9 1 11 7 11 1 15 9 4 13 2 7 2 11 11 2 13 10 0 9 1 0 9 2 3 9 7 9 2
13 9 13 16 15 0 13 14 13 7 13 9 13 2
25 2 11 11 11 2 13 0 1 9 7 9 2 7 11 13 16 0 9 13 10 0 9 1 9 2
7 2 10 9 13 1 15 2
28 15 2 15 2 9 2 9 7 9 4 15 13 9 1 15 2 7 15 4 13 1 16 15 13 15 14 13 2
18 16 15 4 13 1 10 0 9 4 15 13 10 9 1 9 1 9 2
16 3 15 13 10 9 9 7 3 13 9 1 14 13 15 1 2
10 10 9 9 1 9 13 0 1 15 2
2 9 5
18 3 13 15 3 10 0 9 1 11 14 13 1 15 9 11 0 9 2
19 11 11 4 13 1 1 9 1 9 2 7 4 3 13 1 14 13 15 2
42 2 11 11 11 2 13 3 1 14 13 9 15 13 1 2 11 11 2 2 7 4 1 9 13 1 12 9 15 4 13 1 14 13 11 7 11 1 9 7 9 10 2
17 3 4 9 15 13 1 9 13 0 1 10 10 0 9 1 9 2
9 10 0 9 1 9 13 3 1 2
4 0 9 13 5
26 1 9 1 2 11 11 2 4 15 3 13 1 10 1 9 2 7 15 3 4 13 0 1 9 1 2
13 15 4 7 13 0 9 2 7 13 3 10 10 2
32 1 11 13 15 0 14 13 3 10 9 2 7 15 15 13 14 13 13 14 13 9 1 10 9 7 13 15 1 1 9 10 2
28 3 0 4 11 3 13 14 13 0 2 11 11 2 9 2 7 0 9 1 9 4 13 1 0 9 1 9 2
12 15 13 3 0 9 15 4 13 3 1 15 2
15 2 11 11 11 2 4 13 1 9 1 9 1 9 12 2
9 0 4 15 3 13 10 0 9 2
5 13 2 9 13 2
6 7 15 13 3 0 2
25 9 4 13 15 1 16 10 15 0 9 4 13 1 2 13 1 16 15 13 10 0 9 1 11 2
18 15 1 10 9 13 0 10 3 0 16 15 13 9 1 2 11 2 2
26 9 1 9 13 10 9 15 1 9 1 10 0 9 13 15 1 1 10 9 2 16 11 9 13 15 2
32 10 0 15 1 9 1 9 13 2 13 0 14 13 9 2 1 3 14 13 0 10 0 15 4 13 7 13 1 9 7 9 2
19 3 4 15 13 1 9 1 9 2 9 2 9 2 10 9 7 3 0 2
30 1 16 3 15 13 3 2 13 3 9 15 13 15 1 1 1 0 9 15 1 10 7 10 9 4 13 9 1 15 2
13 9 4 13 1 9 2 1 10 3 0 0 9 2
41 3 4 15 3 13 10 9 1 10 0 9 2 15 13 15 1 10 9 1 10 0 0 7 0 9 15 4 13 15 1 10 0 9 2 1 10 9 1 10 9 2
23 15 15 13 1 15 13 3 0 3 0 9 2 1 10 0 9 15 13 1 9 1 9 2
26 3 13 15 3 9 16 15 1 10 9 13 9 1 10 0 3 13 9 15 3 4 13 10 9 1 2
38 16 15 13 11 9 13 15 1 0 10 9 15 13 15 14 13 1 9 1 0 9 2 1 3 14 13 15 1 14 13 1 9 7 13 1 10 9 2
26 15 13 3 1 10 9 2 7 9 13 0 9 2 15 15 3 13 3 0 10 9 15 13 9 0 2
22 15 15 4 13 1 0 9 1 2 11 2 2 13 3 1 10 9 0 1 0 9 2
26 9 13 1 9 2 9 13 0 2 9 13 0 0 1 9 2 7 15 13 7 13 0 15 15 13 2
2 0 2
2 3 2
10 2 11 2 11 7 11 13 12 9 5
6 9 1 9 1 9 2
18 11 11 4 9 13 9 1 11 9 2 11 7 11 9 2 1 11 2
23 9 13 1 1 16 11 7 11 13 12 0 7 0 9 2 16 11 13 9 2 13 11 2
24 9 1 9 13 14 13 9 1 14 13 9 1 14 13 9 1 12 9 2 7 14 13 9 2
22 12 1 9 4 13 9 2 7 15 4 3 13 1 11 11 9 1 9 2 1 9 2
15 11 7 11 13 1 3 12 9 15 13 0 12 9 9 2
18 9 1 11 9 4 13 1 9 1 10 9 7 13 16 9 4 13 2
15 9 13 3 14 13 16 11 13 9 1 9 2 13 15 2
10 13 9 9 1 9 1 2 11 2 5
8 2 8 8 2 8 8 8 2
27 15 13 9 14 13 0 0 16 10 9 1 0 9 2 11 11 2 13 10 3 0 9 1 10 0 9 2
26 9 1 2 11 11 11 2 13 0 1 15 15 4 13 10 9 7 13 10 9 1 9 10 1 9 2
30 10 9 13 1 9 0 9 2 7 11 2 11 7 10 0 0 9 13 1 0 9 1 14 13 15 15 13 0 9 2
23 16 9 3 13 1 9 13 15 1 9 3 12 9 15 13 15 1 2 4 9 3 13 2
9 0 9 13 9 0 9 1 9 2
26 15 4 3 3 13 1 9 2 7 9 1 9 4 15 13 1 1 10 0 2 0 9 15 13 9 2
9 10 9 13 15 1 10 0 9 2
42 1 9 1 14 4 13 1 9 1 0 0 9 2 13 15 1 1 10 9 2 13 2 13 1 10 9 1 9 3 2 4 15 3 13 10 0 9 1 10 0 9 2
31 9 4 13 15 9 1 14 13 10 0 9 2 7 15 4 13 0 9 1 2 8 8 2 8 8 8 2 1 0 9 2
7 9 13 0 3 3 0 2
19 15 4 0 7 0 13 9 15 1 9 1 9 4 13 10 0 9 3 2
15 3 4 2 11 11 11 2 13 0 1 9 15 13 9 2
29 15 13 0 1 9 7 1 9 1 2 11 8 11 2 4 9 13 1 0 9 15 3 13 15 9 1 0 9 2
29 9 13 7 0 7 0 1 10 1 3 9 2 7 9 13 0 7 9 13 3 0 3 1 14 13 15 1 9 2
12 15 13 0 0 9 2 1 14 13 10 9 2
11 4 13 12 0 1 11 14 13 1 9 5
10 2 4 13 9 1 9 2 13 9 2
2 0 2
15 9 11 11 11 1 11 13 0 1 14 13 9 1 9 2
23 1 9 13 15 0 14 13 7 13 7 1 7 1 1 9 1 1 12 0 1 11 9 2
15 9 13 10 0 1 9 1 14 13 10 10 9 1 9 2
23 11 9 13 3 0 9 1 9 1 10 9 1 9 16 9 13 1 9 2 13 11 11 2
2 0 5
25 2 9 7 9 4 3 13 0 7 16 15 13 9 2 7 15 4 13 9 13 1 15 1 9 2
27 3 4 10 9 13 9 7 13 10 9 1 3 15 4 13 2 13 9 9 2 11 11 2 1 11 11 2
22 9 11 11 11 1 11 9 1 9 2 11 2 13 0 0 1 14 13 9 1 9 2
29 2 13 1 15 15 1 9 13 1 9 1 9 1 10 9 9 2 4 9 1 0 9 4 13 0 9 1 9 2
20 9 4 13 0 1 15 7 1 0 9 13 9 1 9 2 13 11 1 11 2
13 9 13 0 9 15 13 1 9 1 9 1 9 2
13 2 16 15 13 0 9 4 3 15 13 1 9 2
42 9 13 16 9 13 12 9 0 0 1 9 2 15 13 3 9 7 9 13 1 0 9 1 9 1 10 0 0 9 1 0 9 1 11 2 13 11 11 11 7 13 2
14 2 10 9 4 13 15 10 9 1 10 0 0 9 2
19 1 0 9 4 15 13 1 0 9 1 10 0 12 9 9 2 13 9 2
4 0 1 9 5
23 0 1 9 13 10 9 9 13 1 11 9 2 10 9 1 14 13 9 1 9 1 9 2
9 11 11 11 13 1 1 10 9 2
11 1 9 1 11 13 15 10 9 1 9 2
28 11 13 15 13 0 9 1 14 13 9 1 9 2 3 16 15 13 9 13 1 3 0 0 9 1 9 9 2
24 2 0 9 1 9 1 14 13 13 9 2 13 9 2 13 9 2 13 9 7 13 0 9 2
16 0 9 4 2 1 9 1 0 9 2 13 15 13 1 9 2
41 15 13 3 15 1 10 9 13 14 13 15 10 9 1 3 0 9 4 13 15 14 13 1 10 9 1 14 13 15 1 10 10 9 2 13 11 11 11 1 11 2
14 11 9 13 9 1 10 0 0 3 1 12 9 3 2
17 3 13 3 11 14 13 10 0 9 2 10 9 1 9 7 9 2
30 2 15 13 10 9 15 4 13 1 9 7 3 0 0 2 13 9 1 9 11 11 1 11 9 1 11 9 1 9 2
7 9 13 3 1 1 9 2
26 10 0 9 1 9 4 13 1 11 1 9 1 9 2 7 9 9 12 4 13 7 13 1 10 9 2
7 2 15 13 3 0 0 5
8 11 11 1 9 1 0 9 2
20 1 12 9 1 3 0 9 1 11 11 13 11 11 11 1 9 9 1 9 2
18 0 9 13 9 1 0 9 1 9 15 0 13 1 1 0 1 9 2
21 11 11 13 0 0 2 7 13 0 9 1 1 9 1 10 0 9 1 11 11 2
18 1 9 13 15 12 9 1 9 11 11 2 1 10 1 3 0 9 2
24 2 15 13 1 14 13 12 9 2 7 4 13 15 1 3 10 9 2 13 11 11 1 11 2
15 2 15 13 3 0 0 2 15 13 3 3 0 1 9 2
52 9 2 15 13 1 1 10 0 9 16 15 1 9 12 13 1 9 2 13 3 0 7 0 3 15 0 10 1 9 3 13 14 13 15 2 7 1 12 9 1 1 9 1 10 0 9 4 15 13 1 0 2
21 2 16 11 11 4 13 10 0 9 13 15 0 14 13 1 12 9 1 0 9 2
20 16 15 3 13 9 13 15 15 10 16 15 13 0 2 13 11 11 1 11 2
7 9 13 9 12 0 9 2
6 11 4 13 1 9 5
4 13 1 9 2
16 11 11 13 3 1 14 13 1 10 0 9 1 11 0 9 2
11 1 12 9 1 9 2 13 15 1 9 2
10 2 15 4 13 1 9 1 12 9 2
7 3 13 15 3 0 0 2
27 3 4 15 13 0 9 1 10 0 2 7 10 9 15 4 13 1 0 11 11 2 13 15 3 15 1 2
38 2 15 13 3 1 11 2 7 1 7 1 16 15 3 13 1 9 1 14 13 7 13 15 2 4 15 3 13 0 1 3 2 13 11 11 1 11 2
43 3 13 15 1 14 13 1 11 7 13 0 1 16 9 1 9 13 1 10 0 9 1 11 2 16 11 11 4 13 11 11 1 9 1 9 1 11 11 11 2 11 2 2
2 9 5
28 2 16 15 3 13 10 9 3 13 10 9 1 15 2 7 15 13 0 15 13 0 1 16 15 4 13 0 2
23 15 13 15 1 11 2 7 15 4 0 13 1 1 14 4 13 1 11 11 2 13 15 2
46 2 1 10 13 15 1 14 13 1 1 10 0 9 9 1 11 2 7 13 1 14 13 1 1 11 3 1 9 2 7 15 13 9 1 16 15 4 13 10 9 3 1 9 1 9 2
27 2 16 15 13 9 2 13 15 1 14 13 10 1 9 1 10 0 9 16 11 11 13 9 2 13 11 2
19 7 15 15 13 0 0 1 13 10 9 1 16 10 9 13 15 1 9 2
2 0 5
35 2 16 15 3 13 9 1 9 2 13 1 10 9 10 10 9 10 1 14 13 9 2 7 15 4 3 13 16 15 13 0 0 1 15 2
33 2 15 13 7 13 15 13 15 15 13 1 1 14 4 13 10 9 2 16 15 13 0 7 0 9 7 10 0 9 2 13 15 2
19 1 9 13 15 1 14 13 11 1 9 1 10 9 1 9 9 5 9 2
12 10 9 15 13 1 14 13 1 13 0 0 2
18 7 9 1 9 7 10 0 9 1 10 1 10 0 9 4 13 0 2
21 15 4 13 0 1 10 9 15 13 16 9 1 10 10 9 13 1 0 1 9 2
5 11 0 1 9 5
8 11 11 4 13 9 1 9 2
16 11 11 7 11 13 1 9 1 9 7 13 3 0 1 9 2
14 15 13 0 1 10 0 9 12 2 12 1 11 9 2
13 1 9 13 11 7 9 1 12 9 1 12 9 2
15 10 10 13 11 2 15 1 1 9 1 9 1 0 9 2
24 11 13 11 7 11 9 2 7 9 1 10 1 15 13 3 1 14 13 1 10 12 0 9 2
11 1 3 9 4 11 13 9 3 10 9 2
19 10 0 9 1 11 11 1 9 2 13 11 12 2 12 1 9 9 9 2
22 9 13 11 9 1 9 1 14 13 9 7 9 1 14 4 13 9 1 9 1 9 2
10 2 9 7 9 13 0 1 10 9 5
8 9 1 11 13 9 1 9 2
7 9 13 3 15 4 13 2
4 0 1 9 2
10 9 11 11 13 0 9 0 1 9 2
17 11 13 9 1 9 2 15 13 15 14 13 1 9 1 0 9 2
6 15 13 1 0 9 2
2 0 2
11 0 9 4 13 1 0 9 7 0 9 2
18 3 4 15 13 0 1 0 9 1 10 0 9 2 1 11 1 11 2
4 3 1 9 2
17 10 9 1 9 7 9 1 10 9 2 13 9 1 9 1 9 2
18 9 13 0 7 10 9 9 4 13 1 0 9 2 1 9 1 11 2
4 1 0 9 2
21 4 10 0 9 1 11 11 4 13 1 1 0 9 2 4 15 4 13 1 9 2
23 1 9 1 4 15 13 0 1 9 1 9 1 9 2 1 9 1 11 2 11 11 11 2
22 1 9 13 11 3 0 0 9 7 9 4 13 1 10 9 1 11 1 9 11 11 2
4 0 1 0 5
28 9 1 9 2 16 0 9 13 0 1 0 9 2 1 9 1 9 2 13 0 1 9 1 11 1 14 13 2
36 2 15 13 0 16 0 9 4 13 0 2 3 16 10 0 15 13 1 15 3 4 13 1 9 2 13 9 1 11 2 11 11 11 1 11 2
21 15 13 9 7 9 2 15 4 13 0 1 10 0 9 2 13 0 7 0 0 2
30 16 0 9 2 1 9 2 13 1 9 1 10 9 7 10 0 9 1 9 2 4 15 13 0 9 1 9 15 13 2
16 2 15 4 13 1 16 10 0 13 10 0 9 2 13 11 2
13 11 13 3 10 9 4 13 1 9 0 1 9 2
3 13 9 5
26 0 9 7 9 2 9 11 11 2 4 3 13 15 1 3 0 15 4 13 9 1 9 1 0 9 2
27 1 9 4 0 9 1 11 11 2 15 13 9 1 9 1 0 9 1 9 2 4 4 13 9 1 9 2
24 2 15 4 3 13 15 16 15 13 15 1 14 13 0 2 13 0 9 11 11 11 1 11 2
13 2 13 15 16 15 13 9 15 13 0 1 9 2
15 2 15 4 3 13 15 1 10 9 2 13 2 13 11 2
16 1 9 4 9 13 9 1 9 1 0 1 9 1 12 9 2
7 9 4 13 0 1 9 2
2 9 5
19 11 13 1 0 1 1 11 2 16 15 13 1 7 9 7 0 9 0 2
17 10 10 9 1 16 10 0 9 7 9 4 13 1 9 13 9 2
18 2 15 13 0 16 15 4 13 9 1 1 9 7 9 15 13 1 2
32 7 16 15 13 9 7 3 0 0 2 3 4 15 13 1 16 15 4 13 9 2 13 9 1 11 2 11 11 11 1 11 2
4 2 13 3 5
13 10 0 9 1 9 0 9 7 0 9 13 9 2
26 16 0 4 13 0 1 9 2 1 9 1 9 1 12 9 9 1 9 2 4 0 9 13 10 9 2
10 2 15 13 3 0 9 3 1 9 2
21 15 13 0 7 4 13 0 2 0 1 0 15 13 1 1 9 3 2 13 11 2
26 1 9 13 15 9 16 9 4 13 1 0 9 2 7 1 0 0 9 1 2 7 0 0 9 1 2
30 2 16 9 3 13 16 0 9 4 0 2 3 13 15 3 16 15 13 0 9 7 4 3 3 13 15 1 0 9 2
34 1 9 2 16 15 13 9 15 13 1 9 1 14 13 1 0 9 1 9 7 0 2 3 4 3 15 3 4 13 10 9 1 15 2
3 13 9 5
21 1 16 11 13 11 11 1 16 15 13 9 1 9 1 9 2 4 15 13 9 2
22 9 13 3 16 9 9 1 14 13 0 9 1 14 13 15 1 9 2 4 13 0 2
8 1 10 9 1 11 13 11 2
26 2 1 10 0 0 9 1 9 1 10 9 1 0 9 2 3 13 15 15 16 15 3 13 10 9 2
23 0 9 13 3 1 9 1 9 1 9 7 15 4 13 10 2 0 9 1 0 9 2 2
22 11 13 0 1 14 13 1 9 1 0 9 7 10 15 13 1 0 9 1 0 9 2
16 9 13 1 12 12 12 12 12 2 11 7 12 12 12 12 2
7 0 4 15 13 9 1 2
8 13 2 0 9 2 1 9 2
5 0 9 1 9 5
5 0 9 1 11 2
11 9 13 0 1 9 2 7 1 7 1 2
10 9 1 11 13 10 0 9 1 9 2
18 3 13 11 9 1 9 1 9 1 9 0 1 9 1 9 1 0 2
18 9 13 1 1 12 9 2 16 9 4 13 1 12 9 1 10 9 2
16 0 13 0 12 9 9 1 7 1 10 1 11 9 1 9 2
34 2 15 13 10 9 1 16 15 1 9 1 4 13 9 1 10 9 1 9 7 9 1 9 2 13 9 11 11 1 10 9 1 9 2
15 11 13 3 1 9 1 0 9 1 9 1 9 1 9 2
26 0 9 1 9 0 9 13 11 11 11 2 15 13 10 9 1 9 9 1 12 9 1 10 0 9 2
33 11 11 11 13 10 9 1 12 9 2 11 9 12 9 2 11 9 11 12 9 2 11 9 11 12 9 7 11 9 11 12 9 2
20 10 0 9 4 13 10 0 9 1 12 9 1 9 0 1 10 9 1 9 2
4 13 9 9 5
9 9 0 9 11 11 2 12 2 2
20 11 11 4 13 15 0 1 9 2 7 3 13 15 10 0 9 1 9 9 2
28 1 0 9 3 13 15 0 16 9 11 11 4 13 15 10 9 1 10 0 9 1 12 9 9 1 12 9 2
20 2 10 9 13 1 9 2 7 10 9 15 13 1 9 2 13 10 10 9 2
5 15 13 0 0 2
25 15 4 13 3 16 9 4 13 1 10 12 9 1 10 0 3 16 9 15 13 13 3 3 0 2
12 9 4 3 13 1 9 2 13 11 1 11 2
17 15 13 15 13 0 0 1 9 2 0 1 9 2 1 10 9 2
22 11 13 15 13 0 0 1 10 9 1 9 7 0 9 14 13 14 13 1 9 10 2
11 2 15 13 3 15 1 14 13 10 9 2
37 15 13 15 3 0 1 14 13 16 15 13 10 9 1 9 1 14 13 10 9 0 1 10 7 10 9 1 1 11 15 15 13 10 9 1 9 2
11 7 10 9 1 0 9 9 1 12 9 2
27 0 9 4 13 1 16 10 9 7 9 15 3 13 1 2 13 10 15 0 0 7 0 9 2 13 11 2
13 11 1 11 13 1 9 7 13 11 13 1 9 2
23 9 1 12 9 9 13 3 1 16 11 4 13 1 11 2 15 13 11 9 2 13 15 2
3 11 11 5
23 13 15 0 9 16 11 13 10 10 9 7 13 0 9 1 10 0 9 2 11 11 2 2
25 16 11 11 3 13 10 9 1 0 9 1 9 2 13 15 3 12 9 15 0 13 9 1 9 2
28 15 13 11 11 2 11 11 2 2 10 9 1 11 2 16 0 9 13 10 12 9 1 9 2 11 11 2 2
27 15 13 0 1 9 7 0 9 7 15 13 15 1 10 9 2 7 1 10 9 13 9 10 9 3 0 2
7 11 11 13 9 1 9 2
32 15 13 0 1 3 9 13 1 2 3 9 13 1 7 3 9 15 13 9 1 9 13 1 2 1 9 1 10 9 15 13 2
14 9 4 13 1 14 13 1 10 9 15 13 13 0 2
15 9 13 11 9 1 12 9 2 10 0 9 9 1 11 2
6 9 13 15 1 9 2
16 13 15 0 14 13 9 1 10 9 2 16 9 13 0 9 2
9 15 13 9 1 9 9 1 11 2
23 13 15 9 1 9 1 10 0 9 2 7 13 15 10 0 9 1 14 13 9 1 9 2
28 11 13 9 1 14 13 9 1 9 2 6 1 14 13 1 15 2 1 14 13 1 16 10 0 13 1 9 2
13 3 4 15 1 9 1 9 13 1 14 13 9 2
5 15 13 15 3 2
20 9 13 3 0 1 15 16 15 13 9 0 1 15 15 13 0 0 1 9 2
12 2 11 11 2 13 10 0 9 15 13 9 2
11 15 13 10 9 2 10 9 7 10 9 2
34 15 13 0 9 1 10 0 0 9 2 0 15 15 13 1 9 1 11 7 11 2 3 3 1 1 9 11 2 10 0 9 1 9 2
21 11 2 15 13 9 1 9 1 11 2 4 13 11 11 9 1 10 9 1 12 2
26 15 4 13 1 16 15 4 13 10 9 9 1 9 1 9 1 9 1 9 2 10 0 9 1 11 2
22 7 11 2 15 4 13 1 11 7 9 7 13 9 9 1 9 2 4 3 13 9 2
6 11 13 3 10 9 2
23 9 13 9 1 14 13 9 2 7 13 3 10 1 14 13 9 7 13 9 1 0 9 2
12 2 15 13 10 9 1 16 15 13 0 9 2
27 15 4 13 11 4 13 15 2 3 13 15 1 10 9 13 10 0 9 2 13 11 11 1 9 1 11 2
10 3 13 10 0 9 1 10 0 9 2
37 0 9 1 9 1 2 11 11 11 2 13 15 1 9 1 10 0 9 12 9 2 10 1 11 7 10 1 11 11 2 15 15 13 0 1 9 2
16 2 15 13 0 0 1 9 2 1 9 1 15 9 4 13 2
14 15 4 13 0 7 0 9 1 9 7 1 0 9 2
17 9 15 4 13 13 7 9 10 1 10 0 9 7 1 9 9 2
16 3 13 15 10 9 1 3 0 9 4 13 15 2 13 11 2
14 11 9 2 11 11 11 2 13 11 9 1 0 9 2
7 2 15 4 15 0 13 2
13 15 15 13 1 9 13 0 1 10 9 0 9 2
10 15 15 13 9 13 10 9 1 9 2
19 16 15 13 2 11 11 2 13 0 2 13 9 1 14 13 9 1 9 2
19 3 13 15 3 16 9 13 3 0 9 1 14 13 0 9 2 13 11 5
39 11 2 15 13 1 11 11 7 1 0 13 1 11 11 2 11 11 7 11 11 2 13 1 9 1 10 9 2 16 15 13 16 11 3 4 13 9 9 2
23 9 13 14 13 9 1 1 0 9 1 9 2 1 14 13 1 1 0 9 1 9 2 2
19 2 10 0 9 13 16 15 13 10 0 9 2 15 13 0 9 1 9 2
23 3 13 15 0 0 16 9 3 4 13 15 2 0 16 15 3 4 4 13 15 0 3 2
17 16 9 13 1 10 0 9 4 15 13 1 0 2 13 11 11 2
19 15 13 16 9 13 0 1 11 0 9 2 3 16 9 13 7 11 13 2
41 1 9 13 9 3 16 2 11 9 1 11 9 4 13 0 1 10 9 1 9 1 11 9 2 2 16 2 9 13 0 1 0 9 15 4 13 1 0 9 2 2
18 15 13 3 10 9 1 9 1 9 9 2 15 13 0 1 0 9 2
20 11 9 4 13 1 9 1 0 9 1 9 10 0 9 2 13 11 11 11 2
21 2 10 0 0 7 0 9 4 13 1 1 14 13 9 1 15 10 9 4 13 2
11 11 2 11 11 2 13 0 1 3 9 2
26 15 7 13 10 0 9 1 10 9 2 7 15 13 9 1 16 15 4 13 1 7 13 1 10 9 2
16 7 11 13 3 16 9 1 11 9 13 0 14 13 1 0 2
38 2 1 10 0 9 13 15 10 9 16 2 11 11 2 13 1 10 0 0 9 2 15 13 16 9 13 10 9 1 2 7 3 3 4 13 1 9 2
21 16 9 13 1 0 2 0 7 0 14 13 15 1 2 13 16 15 13 1 9 2
17 7 15 13 15 13 10 9 1 10 9 9 2 13 11 11 11 2
19 11 11 13 1 9 1 1 11 1 14 13 9 1 2 11 11 12 2 2
11 9 13 0 2 16 10 9 4 13 0 2
14 2 1 11 2 1 1 11 2 13 10 9 0 0 2
9 7 15 13 0 1 10 0 9 2
13 15 13 3 14 13 1 9 1 16 9 13 0 2
12 11 13 16 15 3 13 9 1 10 0 9 2
19 2 10 0 9 13 3 0 10 0 2 16 15 4 13 10 0 0 9 2
17 10 9 1 11 9 13 1 1 14 13 10 9 1 10 0 9 2
52 15 13 3 11 9 1 16 15 4 13 9 15 3 4 13 9 1 2 15 13 3 0 1 1 0 9 2 13 11 2 15 13 16 15 13 9 1 12 0 9 2 3 2 11 11 2 1 11 3 13 12 2
12 9 4 13 16 11 13 9 1 3 1 9 2
13 1 9 13 15 0 14 13 9 1 9 1 11 2
9 15 13 0 14 13 1 9 3 2
4 16 15 13 2
7 11 11 13 9 1 11 2
6 0 9 13 1 9 5
5 13 9 1 11 2
13 12 0 9 4 1 9 13 1 10 0 9 11 2
17 15 4 10 13 12 9 1 9 1 14 4 13 9 1 10 9 2
13 9 4 13 1 11 1 11 9 9 12 1 9 2
19 1 9 11 11 13 9 16 9 11 11 13 1 9 10 7 13 1 15 2
20 10 0 9 4 13 1 9 2 15 13 15 9 1 12 9 7 12 9 10 2
5 15 4 3 13 2
18 11 9 2 7 11 11 11 11 11 11 2 13 12 9 1 1 11 2
18 9 11 13 9 9 1 1 12 9 2 7 13 1 9 10 0 9 2
12 11 4 4 13 1 14 13 1 0 0 9 5
9 9 0 1 12 9 0 1 12 2
3 0 9 2
9 9 13 9 10 0 9 1 9 2
23 11 7 11 4 1 9 13 0 1 16 12 9 1 10 9 1 11 4 13 0 1 12 2
23 10 0 9 7 10 9 15 13 0 0 9 1 1 2 4 13 1 0 2 10 0 0 2
7 2 11 1 1 12 9 5
13 1 9 13 9 0 9 1 11 1 1 12 9 2
17 1 11 13 1 12 9 1 10 9 0 2 1 9 1 10 9 2
19 9 11 11 1 11 13 16 9 13 1 14 13 0 1 11 2 1 9 2
10 2 9 13 3 0 11 4 13 9 2
26 16 15 4 13 10 9 15 4 13 1 10 10 9 2 13 11 1 1 12 9 0 9 2 13 11 2
15 2 11 13 10 0 9 1 9 1 7 9 0 7 9 2
15 10 9 13 0 16 9 13 3 0 1 9 2 13 11 2
19 9 11 11 11 4 3 13 15 1 3 16 15 13 9 1 9 1 11 2
25 2 16 9 4 0 13 2 13 15 0 1 11 14 0 13 9 1 16 15 4 13 1 1 9 2
24 15 4 3 13 1 9 1 11 1 3 15 4 13 15 9 1 0 9 2 13 11 1 11 2
3 0 9 5
14 0 1 9 10 13 1 15 0 9 1 10 0 9 2
16 11 13 3 10 9 1 12 9 2 7 13 1 1 12 9 2
20 11 4 13 10 9 0 2 1 12 2 12 9 7 1 1 12 2 12 9 2
11 2 3 0 13 9 16 15 4 13 15 2
22 15 4 13 0 2 7 15 13 15 13 2 13 9 1 11 2 11 11 2 1 11 2
39 10 9 15 3 13 14 13 1 3 0 9 1 12 2 13 9 1 1 9 14 13 9 1 10 9 2 7 1 9 16 10 0 9 4 4 13 1 11 2
14 3 3 13 11 11 15 13 10 0 0 9 1 11 2
20 2 11 13 9 1 14 13 9 1 0 1 12 9 2 7 13 9 1 11 2
20 15 4 13 0 9 1 0 9 1 9 15 13 14 13 9 10 2 13 11 2
16 11 4 13 1 16 11 13 10 3 0 9 1 11 1 0 2
4 9 13 9 5
19 9 15 4 13 1 9 13 10 9 1 11 9 7 9 15 13 10 9 2
27 11 13 0 0 1 16 9 4 13 14 13 0 1 0 9 2 7 10 0 9 7 0 1 10 0 9 2
11 2 15 4 3 13 0 2 13 11 11 2
20 9 4 13 9 1 16 15 10 9 13 9 16 9 4 13 14 13 1 9 2
20 11 11 11 4 13 1 15 15 4 13 16 15 13 0 9 14 13 1 9 2
10 11 13 0 9 1 11 9 7 9 2
16 10 3 0 9 13 2 3 15 15 13 9 7 9 7 9 2
19 13 15 10 0 9 1 9 2 4 15 13 10 9 1 9 9 1 11 2
13 15 4 13 1 9 7 9 1 11 9 7 9 2
19 9 10 9 13 9 1 10 0 9 1 9 15 13 0 1 11 2 11 2
32 2 15 13 0 16 11 4 13 10 9 7 9 2 7 3 0 16 15 13 1 9 2 13 9 11 11 1 10 9 0 9 2
3 13 3 2
7 11 0 9 2 9 2 2
10 2 4 13 3 3 16 15 13 0 5
9 11 11 13 0 1 9 1 0 2
3 13 9 2
16 11 11 1 11 11 13 0 13 1 1 0 9 1 3 9 2
2 0 2
12 11 11 11 13 15 13 0 15 3 13 0 2
4 5 13 3 2
9 13 9 1 16 9 13 1 9 5
23 11 11 13 16 9 13 9 3 0 1 10 9 2 1 1 1 16 0 13 1 10 9 2
9 2 15 13 9 3 0 1 0 2
8 1 15 13 9 10 9 9 2
14 15 13 3 3 16 15 13 0 14 13 15 1 15 2
14 15 13 3 16 15 4 13 0 2 13 11 1 11 2
5 4 13 1 9 5
19 15 13 0 1 0 11 9 1 1 12 2 7 13 1 9 3 0 9 2
17 1 9 13 0 9 0 9 9 1 15 1 9 1 10 0 9 2
7 9 4 13 1 10 9 2
16 11 13 16 15 13 0 14 4 13 10 1 12 9 1 9 2
12 15 13 3 3 0 16 9 4 13 1 9 2
12 9 13 3 1 2 7 1 9 1 2 9 2
12 2 9 13 1 7 1 7 3 3 3 0 2
29 15 4 13 10 9 1 16 15 13 2 1 3 14 4 13 12 9 1 9 1 10 9 1 12 9 2 13 15 2
20 7 11 13 9 9 13 2 7 16 15 13 0 14 13 9 1 9 9 1 2
5 2 4 13 0 5
20 2 15 13 1 9 16 15 4 4 13 0 1 9 1 14 13 10 0 9 2
10 15 4 13 9 1 9 2 13 11 2
23 15 13 10 0 9 1 10 0 2 7 0 9 16 9 1 10 9 4 13 3 15 13 2
24 2 15 13 16 15 4 13 10 9 1 15 10 3 16 15 13 15 14 13 1 2 13 11 2
9 2 15 4 13 0 9 1 0 2
11 13 15 15 14 13 1 9 1 10 9 2
16 2 6 2 0 13 10 0 9 3 9 0 13 10 0 9 2
17 11 13 0 1 16 9 4 13 0 9 1 9 1 9 1 9 2
10 15 13 9 15 3 7 3 4 13 2
37 2 7 15 15 13 0 1 0 13 15 13 3 0 9 1 9 16 15 3 13 2 0 1 14 13 15 2 1 14 13 15 2 13 10 0 9 2
8 13 11 2 7 3 1 9 2
20 11 11 1 11 11 13 16 9 1 11 11 11 1 9 13 1 0 1 11 2
6 2 15 13 0 0 2
22 15 13 1 15 1 9 1 15 15 13 1 9 1 9 2 13 9 1 10 0 9 2
24 2 15 13 0 1 14 13 15 16 15 13 14 13 3 1 9 2 13 11 11 11 1 11 2
10 2 7 1 9 7 9 13 9 0 2
16 7 1 16 15 13 14 13 1 9 3 4 15 0 13 15 2
19 2 15 13 3 0 2 7 0 15 4 4 13 12 9 1 1 1 15 2
8 2 13 15 15 13 3 0 2
10 2 15 13 1 10 9 3 3 0 2
14 7 15 13 0 0 1 16 15 3 4 4 13 0 2
21 7 16 15 4 13 2 11 11 7 11 13 0 15 15 13 7 13 10 9 3 2
20 1 15 13 15 0 0 16 9 13 0 1 9 16 9 7 9 13 0 9 2
16 1 10 0 9 1 0 13 15 3 3 0 0 1 14 13 2
19 11 11 11 4 13 0 16 15 4 13 3 1 11 11 1 12 9 3 2
7 16 15 13 0 1 9 2
9 2 3 13 15 7 15 13 0 2
19 13 15 0 1 9 4 15 0 13 1 10 9 1 9 2 3 7 3 2
17 7 1 9 2 6 2 15 13 3 15 4 4 13 10 12 9 2
6 7 15 13 0 0 2
12 15 13 10 0 11 11 2 12 2 13 3 2
4 10 10 9 2
2 0 2
18 1 9 2 11 1 10 10 0 2 7 1 9 2 11 0 9 2 2
2 13 2
4 16 9 13 2
11 15 13 10 0 15 13 1 9 10 3 2
7 2 6 2 15 13 0 2
20 0 9 9 2 0 9 2 0 9 7 0 9 3 16 15 13 1 7 13 2
4 7 10 0 2
11 2 16 9 1 9 0 13 1 9 12 2
4 10 9 13 2
5 2 2 11 2 2
11 3 13 1 2 13 9 7 9 1 15 2
5 3 13 15 3 2
4 2 1 11 2
5 15 13 15 3 2
39 2 15 4 13 10 0 9 1 12 9 2 7 10 12 9 13 9 2 7 3 13 15 11 2 16 11 10 9 15 15 13 13 12 0 9 0 7 0 2
16 15 13 3 9 16 15 15 13 0 13 0 1 11 7 11 2
32 15 4 13 15 1 14 13 0 9 1 9 2 13 15 1 0 9 15 13 0 1 9 7 13 10 0 9 1 9 1 9 2
5 15 13 10 9 2
15 2 15 13 0 3 1 2 7 15 13 3 12 0 9 2
6 11 2 11 7 11 2
4 7 1 11 2
3 2 6 2
15 13 3 0 16 9 10 13 14 13 1 1 11 0 9 2
8 3 13 10 0 9 1 11 2
31 2 15 4 13 15 13 11 2 7 15 13 14 13 3 16 9 4 13 10 1 16 15 13 0 9 1 14 13 1 11 2
9 10 9 13 15 1 14 13 1 2
3 2 11 2
21 15 4 13 1 10 10 9 3 10 9 0 1 9 7 9 13 0 1 9 10 2
24 10 9 4 13 1 0 9 1 11 10 0 2 7 15 4 1 3 13 14 13 7 13 9 2
17 15 4 13 0 0 9 7 9 1 14 13 10 9 1 10 9 2
8 13 15 1 9 16 15 13 2
15 2 6 2 15 13 15 0 16 12 9 1 9 13 9 2
7 15 13 15 1 1 9 2
5 2 15 13 9 2
18 15 13 3 9 2 16 9 1 10 9 3 13 9 2 15 15 13 2
5 3 0 13 15 2
17 2 10 9 1 9 7 0 1 9 16 15 13 1 9 1 9 2
8 3 0 9 13 15 1 9 2
5 2 15 13 9 2
14 15 13 9 7 13 3 9 1 14 13 1 1 11 2
5 15 13 9 10 2
21 2 15 13 1 1 14 13 10 9 13 15 1 10 9 15 15 13 0 0 1 2
6 15 13 15 9 1 2
9 2 3 13 15 9 16 15 13 2
8 15 13 15 1 15 1 9 2
11 2 9 2 9 2 9 7 9 1 9 2
12 10 12 9 13 15 1 16 15 13 14 13 2
10 2 9 2 0 9 1 9 7 9 2
6 3 13 15 9 10 2
14 2 16 15 4 13 10 9 7 13 15 1 1 15 2
8 15 13 10 0 15 13 3 2
3 2 9 2
11 15 13 15 10 0 12 9 16 9 13 2
4 2 13 9 2
2 11 5
4 10 0 9 5
10 11 13 0 1 9 2 9 7 9 2
13 3 4 9 11 11 11 13 0 9 1 1 9 2
2 9 2
11 11 1 11 13 1 9 11 3 13 1 2
17 16 11 13 1 10 0 9 11 11 2 13 15 16 11 13 9 2
29 2 15 13 10 0 9 1 7 9 2 1 9 7 9 1 9 2 1 11 2 7 1 11 7 11 2 13 15 2
3 13 9 2
16 11 1 11 4 3 13 0 9 1 0 9 7 13 0 0 2
4 3 13 9 2
16 11 11 11 4 3 13 9 1 15 15 0 4 13 10 9 2
3 0 11 2
8 11 7 11 13 10 11 9 2
9 1 11 0 9 13 11 1 11 2
2 0 2
20 2 9 4 13 10 0 9 1 11 2 13 11 11 11 2 15 13 11 9 2
2 0 2
20 0 9 4 13 10 1 16 15 4 13 10 9 14 13 1 11 0 0 9 2
12 3 4 11 9 13 0 9 1 11 1 11 2
3 0 9 2
8 11 1 11 4 13 0 9 2
2 11 2
6 11 1 9 1 11 2
3 0 1 2
7 11 4 13 1 9 11 2
4 9 1 12 2
19 10 0 11 4 13 1 9 11 7 11 7 13 10 9 1 9 11 11 2
3 0 9 2
20 11 11 13 9 7 13 1 11 3 1 11 11 3 1 14 13 10 0 9 2
17 2 9 1 9 4 13 1 9 15 13 2 13 9 11 11 11 2
22 2 9 13 10 0 9 2 1 9 1 9 7 9 2 7 3 13 15 3 1 9 2
9 9 13 9 1 9 2 0 13 2
22 1 1 3 4 9 2 9 7 9 13 15 15 9 0 4 13 1 9 2 11 2 2
18 7 3 13 11 11 11 7 11 2 11 2 1 14 13 11 1 9 2
16 2 0 0 9 4 13 10 9 1 10 0 9 2 13 11 2
30 9 13 16 10 0 9 4 13 2 16 11 4 13 10 9 0 13 9 1 14 13 7 9 13 9 1 14 13 1 2
19 9 2 9 7 9 1 0 9 13 3 9 1 1 9 1 11 7 11 2
28 0 13 9 7 9 1 10 9 1 11 1 14 13 9 1 11 1 11 2 11 1 11 7 11 11 1 11 2
7 7 9 4 3 13 9 2
14 11 7 11 13 0 0 1 9 7 9 1 10 9 2
19 1 10 9 13 9 1 16 10 0 9 13 9 1 10 0 9 11 11 2
29 2 15 13 10 0 9 1 7 9 2 1 9 7 9 1 9 2 1 11 2 7 1 11 7 11 2 13 11 2
13 15 13 9 1 0 9 7 13 1 3 15 13 2
32 2 3 13 15 15 3 1 9 15 4 13 10 9 2 13 10 9 2 1 10 9 1 9 1 10 9 1 9 2 13 11 2
40 2 15 13 10 0 9 1 0 9 15 13 10 9 1 9 2 1 9 7 1 9 2 10 0 9 1 9 1 0 9 2 9 7 9 2 7 0 0 9 2
8 15 13 0 1 10 10 9 2
23 1 11 11 2 0 9 1 11 9 9 2 13 15 3 10 9 9 11 4 13 0 1 2
18 2 1 11 13 15 0 1 14 13 9 7 13 1 9 2 13 11 2
8 2 15 13 9 15 4 13 2
16 0 9 13 10 0 7 0 9 7 13 10 9 1 10 0 2
15 11 11 11 13 10 0 1 7 9 7 9 2 13 15 2
16 11 13 10 0 0 9 15 4 4 13 1 9 1 0 9 2
30 0 9 2 0 9 7 11 9 13 1 14 13 1 10 1 10 0 0 9 1 11 2 1 9 1 11 7 1 11 2
18 9 7 9 1 0 9 7 9 1 9 4 13 9 1 0 1 11 2
24 10 0 9 4 3 4 13 0 1 11 2 7 4 4 13 1 10 0 9 1 11 1 11 2
20 2 11 2 9 13 9 1 10 9 1 11 1 9 2 13 1 10 0 9 2
19 3 0 9 1 11 7 11 7 11 7 11 4 13 10 10 9 1 11 2
20 2 15 4 13 1 0 9 1 0 9 2 13 9 11 11 1 9 1 11 2
22 2 10 9 1 0 9 1 11 7 11 1 9 13 0 9 2 7 3 13 10 0 2
9 11 11 13 11 0 9 1 9 2
8 2 15 13 0 2 13 11 2
42 2 15 4 13 1 0 1 16 9 1 11 3 4 13 1 0 9 16 15 13 1 9 2 7 1 14 13 10 0 9 15 13 9 1 14 13 1 14 13 0 9 2
13 15 4 13 9 2 3 15 13 1 9 7 9 2
9 9 4 13 10 0 9 1 11 2
11 7 15 13 3 15 15 13 9 13 0 2
21 11 11 2 9 1 9 1 11 2 13 15 16 11 4 13 10 0 9 1 9 2
26 2 16 9 13 14 13 10 9 15 13 1 1 11 2 11 7 11 2 13 15 10 9 2 13 15 2
16 2 10 0 9 4 13 14 13 15 1 0 9 7 0 9 2
18 15 13 1 9 2 7 1 10 9 4 15 13 0 14 13 10 9 2
16 16 11 3 4 13 15 0 2 13 3 11 11 11 0 1 2
14 2 15 4 3 13 9 1 9 1 9 2 13 15 2
30 2 15 4 3 13 9 1 9 7 9 15 4 13 15 0 2 7 0 9 7 9 13 10 0 9 1 10 0 9 2
25 7 9 1 14 13 9 7 9 1 14 13 15 1 3 2 1 9 10 9 2 13 9 1 0 2
9 11 11 13 1 15 11 4 13 2
27 2 16 9 13 14 13 9 1 11 2 4 15 3 13 9 16 15 13 15 13 2 1 9 1 0 9 2
40 10 9 15 13 0 1 11 9 1 9 2 13 15 16 0 9 2 15 0 13 0 7 0 1 10 9 2 13 15 1 14 13 9 1 10 0 7 0 9 2
18 9 1 11 11 11 11 13 15 13 0 14 13 9 1 1 10 9 2
14 2 15 13 3 10 0 1 16 11 13 9 1 9 2
8 7 9 13 0 0 7 0 2
13 15 13 15 16 10 9 13 0 9 2 13 11 2
7 2 4 15 13 9 3 2
29 15 13 10 0 9 0 2 7 16 15 13 9 1 9 9 15 4 13 10 0 2 13 15 3 0 1 0 9 2
21 11 11 11 13 3 14 13 7 9 7 10 9 1 15 15 0 4 13 10 9 2
21 2 0 9 13 3 1 9 14 13 0 9 7 0 0 9 1 9 2 13 15 2
12 2 9 7 0 9 13 0 3 1 15 10 2
16 15 4 3 13 15 0 16 10 0 9 13 10 9 1 11 2
16 7 15 13 10 9 16 15 13 10 9 15 13 0 7 0 2
20 16 9 1 10 9 13 15 13 1 0 9 2 3 13 15 9 1 10 9 2
5 13 15 15 13 2
9 15 13 9 1 1 11 1 11 2
10 3 13 15 0 1 11 11 1 11 2
25 2 15 13 1 1 9 10 7 13 2 6 2 15 1 10 9 13 15 1 15 2 2 13 11 2
7 2 15 13 10 0 9 2
6 11 4 13 15 0 2
14 15 13 10 0 10 9 16 15 13 1 10 9 3 2
15 15 13 11 4 13 1 1 14 13 9 1 15 15 13 2
12 0 11 11 11 13 11 13 2 3 0 2 2
8 2 15 13 1 13 1 9 2
46 7 15 13 0 1 3 0 9 1 1 9 2 7 10 0 2 0 9 1 9 13 2 13 11 2 16 11 11 7 11 11 1 11 13 11 13 1 1 10 9 15 13 1 1 9 2
6 2 9 13 0 0 2
14 15 13 1 16 9 13 0 9 7 13 1 0 9 2
14 15 13 10 0 9 14 13 11 1 2 13 10 12 2
7 7 9 13 3 3 9 2
17 16 0 7 0 9 4 13 9 2 13 10 0 9 1 1 11 2
32 3 13 9 1 10 0 9 1 9 2 1 10 1 12 9 0 9 16 9 4 13 0 0 1 10 0 9 11 11 0 9 2
27 3 4 9 13 9 7 9 16 9 13 1 9 7 9 7 4 13 9 1 7 9 0 10 9 1 15 2
16 11 11 1 11 9 9 13 15 13 0 16 0 9 13 0 2
8 2 9 13 14 13 10 0 2
16 15 13 3 10 9 1 14 13 9 16 15 4 13 10 9 2
23 3 11 11 11 13 9 4 13 9 3 3 16 15 13 0 0 16 9 13 0 7 3 2
18 2 0 13 15 3 10 0 9 15 13 14 13 9 7 13 0 9 2
18 15 13 14 13 9 3 1 14 13 9 2 13 7 13 15 1 9 2
34 10 1 10 0 0 9 1 16 0 9 4 13 9 7 13 9 2 13 1 9 9 1 11 2 13 1 0 11 2 15 13 1 12 2
35 2 15 13 10 0 0 9 1 9 7 9 1 9 2 15 13 1 9 1 1 7 1 2 1 7 1 7 1 0 7 0 9 7 9 2
12 9 1 9 2 9 7 9 13 0 10 9 2
4 15 13 9 2
18 9 13 0 0 2 15 13 3 9 1 0 9 7 9 1 10 9 2
8 3 4 3 9 13 15 3 2
16 2 15 13 15 4 13 16 9 13 9 2 13 11 11 11 2
18 2 15 13 3 0 1 16 9 13 0 0 1 0 9 1 10 9 2
7 15 13 9 1 9 10 2
10 9 13 11 11 1 14 13 1 9 5
6 9 4 13 1 9 2
20 1 9 1 9 1 9 11 11 2 11 2 13 10 0 9 14 13 0 9 2
34 1 16 10 9 13 1 9 7 13 10 12 9 0 9 1 1 9 2 4 15 13 1 9 1 1 9 1 9 1 9 1 9 12 2
33 1 9 1 11 9 13 15 0 16 9 2 12 2 3 13 9 1 13 1 12 9 1 9 15 13 9 4 13 9 15 4 13 2
15 9 13 3 1 12 9 1 11 11 16 15 0 4 13 2
28 16 9 13 14 13 9 9 2 4 3 10 12 1 9 4 13 16 15 4 13 9 16 9 3 4 13 1 2
44 2 0 4 13 16 15 13 15 1 0 16 15 4 13 1 9 0 11 9 2 7 15 13 3 1 9 1 16 15 13 1 9 1 14 13 9 1 9 2 13 15 1 9 2
15 10 10 12 4 13 1 0 9 1 1 12 7 12 9 2
9 11 11 4 13 10 9 1 12 5
6 16 15 13 14 13 2
7 3 13 10 0 9 1 2
23 2 3 4 15 3 13 7 13 0 1 9 2 3 16 10 0 9 3 13 1 10 9 2
22 3 1 1 9 2 1 9 2 9 2 9 7 9 2 15 1 9 2 9 7 9 2
10 9 1 9 2 9 2 9 2 11 2
8 0 9 2 3 9 7 9 2
4 10 9 13 2
20 2 2 11 12 2 1 11 11 13 3 10 9 15 4 13 0 1 10 9 2
9 13 0 0 1 11 0 0 9 2
12 3 10 0 0 9 2 7 3 10 0 9 2
7 15 13 15 1 1 9 2
47 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 7 10 9 10 9 1 0 9 15 3 3 13 3 9 1 2
10 7 3 4 15 3 13 9 1 11 2
13 13 15 3 9 7 4 15 13 15 1 10 9 2
16 2 13 3 0 3 2 7 13 1 0 9 7 13 15 0 2
5 15 13 9 10 2
13 2 2 11 8 8 11 2 1 11 13 0 1 2
7 2 11 2 1 11 3 2
14 3 13 15 10 9 16 11 11 13 11 9 1 9 2
8 15 13 15 0 1 1 9 2
2 3 2
6 2 9 13 10 9 2
15 16 15 13 2 11 2 1 9 2 4 15 13 1 9 2
15 0 11 2 16 15 13 1 11 5 9 13 3 0 0 2
6 15 13 15 9 1 2
11 2 15 13 3 2 7 3 1 12 0 2
6 4 3 13 10 9 2
5 15 13 10 9 2
6 2 11 13 0 9 2
12 0 0 9 2 1 9 2 7 10 0 9 2
4 7 1 11 2
7 2 13 1 9 1 11 2
6 1 9 1 7 1 2
5 3 0 13 15 2
9 10 9 13 15 1 14 13 1 2
3 2 11 2
5 3 13 15 3 2
20 2 13 1 9 1 11 7 11 1 9 1 2 11 15 2 9 1 11 11 2
8 13 15 1 9 16 15 13 2
27 2 13 1 9 7 13 14 13 1 9 1 9 2 1 16 15 13 2 7 3 4 13 0 1 7 1 2
8 15 13 15 1 15 1 9 2
10 2 1 10 9 9 2 9 7 9 2
6 7 9 1 9 10 2
7 3 0 9 4 15 13 2
32 2 10 9 1 11 1 11 7 10 9 1 11 2 13 10 9 9 1 11 7 11 13 9 1 10 10 9 1 11 1 9 2
12 10 0 9 14 13 2 7 14 13 1 1 2
12 10 12 9 13 15 1 16 15 13 14 13 2
26 2 9 2 11 10 2 10 0 9 1 12 2 11 9 10 7 10 9 9 10 11 11 11 4 13 2
13 10 0 13 3 3 9 2 7 15 13 15 1 2
6 3 13 15 9 10 2
13 2 0 1 11 2 7 0 1 0 9 1 9 2
12 13 3 0 0 0 9 2 1 9 7 15 2
8 15 13 10 0 15 13 3 2
7 2 13 9 1 10 9 2
21 13 10 0 9 2 3 16 15 0 13 1 9 16 15 13 1 7 13 0 9 2
10 13 10 0 9 1 9 2 1 9 2
11 15 13 15 10 0 12 9 16 9 13 2
28 2 13 0 0 1 16 15 4 13 3 0 9 2 7 4 13 1 1 9 2 15 3 13 15 14 13 9 2
7 15 13 9 0 0 9 5
7 3 4 15 13 1 11 2
3 0 9 2
14 11 13 0 1 10 0 9 1 10 9 9 7 9 2
2 9 2
23 9 11 13 9 1 9 2 11 2 2 15 13 0 16 15 4 13 1 15 1 11 11 2
2 9 2
2 9 2
2 9 2
15 16 11 11 13 10 0 9 1 11 1 12 13 9 9 2
17 10 9 1 12 13 16 9 13 0 3 1 9 1 9 7 9 2
19 9 7 9 1 11 13 0 1 9 1 0 9 7 13 1 10 9 9 2
4 0 0 9 2
14 11 11 13 9 1 1 10 0 9 1 9 1 9 2
16 3 13 15 7 13 1 9 1 11 9 11 1 11 1 12 2
2 9 2
2 11 5
25 2 15 13 3 10 9 2 13 11 2 13 1 11 11 2 1 10 9 1 2 9 7 9 2 2
6 2 8 8 8 8 2
28 11 13 9 1 15 0 9 4 13 1 10 0 9 1 9 11 2 15 1 10 9 13 10 0 9 1 11 2
66 1 14 13 9 1 10 10 10 4 15 3 13 1 9 1 12 9 7 13 0 1 14 13 1 1 1 12 7 12 9 9 2 16 15 3 3 13 1 2 11 11 11 2 2 10 9 1 9 15 13 15 0 10 9 9 7 15 15 3 13 12 9 1 1 9 2
24 11 7 9 13 15 1 3 0 10 9 4 13 0 1 14 13 1 14 13 9 1 10 9 2
8 15 4 13 9 1 0 9 2
43 0 1 9 13 11 11 2 11 11 11 11 2 9 11 0 11 11 8 8 11 11 11 11 2 2 15 13 1 10 0 9 1 11 1 14 13 1 2 3 2 10 9 2
24 2 15 13 0 3 9 1 14 4 13 1 10 2 11 7 9 2 9 2 13 11 11 11 2
23 15 13 0 9 1 9 11 11 2 15 1 12 13 10 0 9 1 11 1 14 13 9 2
18 3 13 11 11 1 11 1 14 13 9 0 0 9 1 11 7 11 2
17 2 15 13 1 3 14 13 9 13 1 2 7 15 13 3 0 2
19 15 13 3 14 13 15 10 3 0 2 7 15 4 3 13 0 7 0 2
8 7 15 13 0 0 1 9 2
24 7 1 10 9 15 0 13 9 1 9 9 2 13 11 9 1 10 0 9 7 13 15 0 2
31 7 16 15 3 2 1 1 1 10 0 9 2 13 10 0 9 1 11 2 13 11 11 11 16 15 4 13 1 14 13 2
6 2 15 13 3 0 2
12 15 13 3 3 1 14 13 15 1 12 9 2
20 15 13 0 1 9 9 15 13 9 1 11 0 9 2 9 2 9 7 9 2
46 7 16 9 10 0 9 4 13 1 0 9 2 13 11 1 10 0 9 1 10 9 1 2 11 2 2 13 1 9 7 9 11 11 2 7 2 11 2 2 15 13 9 1 11 11 2
32 2 16 15 4 13 10 11 7 10 11 4 15 13 15 1 12 9 2 3 1 14 13 1 1 9 9 2 13 11 11 11 2
13 9 4 1 10 0 9 13 10 0 9 1 9 2
34 10 9 13 10 9 7 10 9 2 7 0 0 9 15 3 13 9 1 11 9 2 13 0 9 1 9 1 11 11 2 11 7 11 2
19 2 9 1 9 4 1 0 9 13 1 9 1 9 2 13 11 11 11 2
10 2 15 13 3 0 1 15 1 11 2
19 9 4 13 0 0 2 7 9 1 9 13 3 11 7 11 1 10 9 2
10 15 4 13 10 0 0 9 1 15 2
29 16 15 4 13 15 2 13 3 10 1 9 1 16 0 13 0 9 16 10 9 4 13 10 9 1 9 7 9 2
28 14 13 10 0 9 1 9 13 1 9 16 15 2 7 9 10 7 9 10 2 13 9 1 14 13 10 10 2
16 15 13 1 10 0 9 2 16 10 9 3 13 9 10 9 2
11 2 15 13 10 0 15 13 9 10 9 2
8 1 15 13 15 3 3 9 2
8 15 13 9 1 15 11 13 2
12 15 13 15 3 10 9 13 9 1 10 9 2
14 10 1 9 1 10 0 9 1 9 13 9 0 9 2
24 11 13 15 0 10 0 9 1 11 9 2 7 10 0 9 13 1 15 15 13 9 1 11 2
25 7 15 13 11 11 9 11 2 11 11 11 9 2 15 13 9 1 9 2 1 0 9 1 9 2
10 2 9 10 13 10 0 7 0 9 2
8 15 13 14 13 1 9 10 2
8 2 13 15 9 10 2 2 2
13 16 15 13 0 1 9 2 13 15 15 10 9 2
19 7 3 7 0 2 13 11 11 2 13 11 11 10 9 15 3 13 9 2
30 2 15 13 16 9 4 13 9 2 7 15 13 3 16 11 4 13 10 9 1 9 7 9 1 14 13 9 7 9 2
15 15 13 0 1 9 7 13 10 0 15 13 9 1 9 2
15 16 15 3 4 13 3 2 4 9 13 9 2 7 13 2
14 3 11 11 9 2 11 11 9 2 13 9 1 9 2
10 2 15 13 15 0 2 13 11 11 2
20 2 15 13 10 9 15 3 3 13 0 2 7 15 15 3 13 0 9 1 2
10 15 4 13 10 9 1 15 0 9 2
14 15 13 15 0 1 9 2 7 13 3 0 1 15 2
12 15 13 0 2 7 0 7 0 1 10 0 2
13 15 13 15 11 9 15 13 10 0 9 1 12 2
24 10 9 13 15 2 11 8 8 2 7 4 13 1 9 1 10 0 9 1 14 13 9 1 2
9 7 15 13 3 1 12 9 13 2
29 3 4 9 11 1 11 2 0 11 11 2 13 1 11 11 16 15 13 9 1 15 1 14 13 16 15 13 0 2
5 0 13 9 0 2
55 10 12 9 15 13 0 0 1 10 9 13 3 10 2 0 11 2 2 9 15 13 1 16 11 11 13 9 7 11 11 9 11 11 1 10 9 1 12 7 13 16 15 3 4 13 10 0 7 0 0 9 1 10 9 2
22 1 9 13 9 1 11 11 11 2 11 11 2 11 11 7 11 11 1 9 1 9 2
15 11 11 2 15 13 9 1 3 12 9 9 2 13 12 2
49 7 16 10 0 11 11 13 1 1 9 10 1 10 11 1 9 2 13 15 1 9 10 0 9 1 9 16 15 4 13 10 10 9 1 14 13 1 1 10 9 15 13 10 0 9 1 0 9 2
15 11 11 11 2 15 13 9 1 11 11 2 13 1 9 2
18 2 9 15 4 13 10 1 10 9 4 4 13 15 15 13 1 15 2
22 7 3 13 15 3 1 16 10 9 1 11 4 13 15 10 11 0 13 2 13 15 2
17 3 13 15 10 0 11 9 2 15 4 13 1 15 1 0 9 2
7 2 15 13 1 0 9 2
13 16 15 13 15 2 13 15 0 0 2 13 15 2
6 2 3 13 15 0 2
7 15 4 13 3 1 15 2
9 15 13 3 15 4 13 1 11 2
5 11 13 1 11 5
5 13 11 11 11 2
2 9 2
16 9 11 11 13 1 9 15 13 11 11 11 10 9 1 9 2
2 9 2
4 11 11 11 2
23 1 10 9 4 9 11 11 2 12 2 13 1 9 1 11 11 11 10 9 1 9 9 2
8 2 11 13 10 3 0 9 2
15 15 13 16 15 13 1 11 2 7 13 0 1 15 3 2
16 15 13 0 0 14 13 15 3 2 13 11 11 2 12 2 2
9 15 13 11 11 11 10 0 9 2
18 16 10 0 9 13 9 1 10 0 9 2 4 11 11 13 1 9 2
21 2 15 13 0 0 1 16 15 13 15 9 1 14 13 2 13 11 11 11 0 2
4 9 1 11 5
39 9 13 1 0 0 9 2 1 10 10 9 1 11 11 16 9 13 11 1 0 9 2 7 13 16 15 10 4 13 0 1 14 13 9 1 10 0 9 2
12 11 13 9 11 11 0 9 1 9 1 11 2
34 2 15 13 3 10 0 0 9 2 7 15 13 3 1 9 2 7 11 7 11 13 3 15 1 15 2 13 10 0 9 1 10 9 2
35 1 10 13 9 11 11 1 10 9 11 13 9 1 11 7 13 1 9 1 10 9 15 13 1 9 2 15 15 4 13 0 1 9 9 2
3 0 9 5
14 15 4 3 13 1 9 16 11 9 4 13 1 9 2
21 9 1 10 0 9 4 1 10 7 10 9 13 1 0 7 0 2 9 13 0 2
8 1 9 13 9 1 1 9 2
18 2 11 13 0 0 2 15 4 13 3 0 9 1 2 13 11 11 2
17 15 7 11 13 1 9 1 11 2 16 11 13 1 11 8 8 2
6 11 13 1 10 9 2
5 13 15 1 9 5
13 1 9 10 9 13 11 11 11 15 1 11 11 2
11 9 13 9 1 10 0 9 1 11 11 2
8 2 15 13 15 15 0 1 2
15 15 13 3 0 0 16 15 4 4 13 10 9 2 3 2
13 15 4 15 3 13 0 2 13 11 1 11 12 2
19 11 13 0 0 1 11 11 2 7 13 3 16 15 13 9 1 11 11 2
7 2 3 13 15 0 0 2
12 3 13 15 3 0 2 13 11 1 11 12 2
9 9 15 3 4 13 10 1 9 5
12 11 11 2 12 2 13 10 1 11 0 9 2
4 9 1 9 2
4 0 1 11 2
10 3 13 15 3 14 13 10 10 9 2
2 0 2
19 2 15 4 3 13 15 15 13 2 3 13 15 15 15 13 2 1 9 2
7 15 4 13 1 2 13 2
11 7 15 4 13 16 15 3 13 9 3 2
3 13 3 2
14 11 11 13 1 10 0 9 7 9 10 9 13 1 2
12 9 7 9 13 15 1 14 13 14 13 9 2
3 9 9 2
17 15 13 1 14 13 1 11 7 11 9 11 11 16 15 13 0 2
8 9 13 3 14 13 1 9 2
4 7 9 13 2
2 9 2
11 11 1 9 2 1 9 1 9 11 11 2
2 9 2
5 15 13 1 11 2
4 7 1 11 2
4 0 7 0 2
8 11 13 7 1 11 7 11 2
8 3 13 15 9 11 1 11 2
3 0 9 2
9 11 9 1 11 13 0 7 0 2
12 3 4 15 13 15 1 11 11 1 10 9 2
6 4 13 9 1 15 2
6 2 3 13 15 15 2
11 1 9 3 2 1 10 9 2 13 11 2
4 9 7 9 2
17 2 15 13 3 15 13 3 1 11 2 1 14 13 1 9 10 2
17 2 8 8 8 2 8 2 8 2 8 8 8 2 2 13 15 2
22 2 10 12 9 15 13 1 9 13 16 15 12 9 1 9 13 1 11 9 1 9 2
7 3 13 9 9 1 9 2
2 0 2
3 0 9 2
10 15 13 15 0 7 0 0 1 9 2
6 15 13 3 1 9 2
13 3 4 15 13 9 7 9 2 1 9 1 11 2
5 13 0 1 11 2
25 1 9 9 4 15 13 1 9 1 11 2 13 11 11 0 9 1 9 7 13 9 11 11 11 2
13 2 16 15 13 9 0 9 2 13 15 0 0 2
11 15 13 10 9 1 9 7 13 1 15 2
8 1 9 13 15 11 11 11 2
12 15 13 1 9 1 9 1 0 7 0 9 2
8 15 13 15 3 1 10 9 2
12 15 13 9 1 10 9 15 4 13 10 9 2
19 9 1 10 9 15 13 10 9 2 13 10 9 1 14 13 7 13 15 2
45 15 15 13 10 9 13 1 10 9 10 0 0 9 15 13 16 10 0 15 13 3 1 15 13 15 1 14 13 1 1 10 0 9 16 9 7 9 13 10 12 15 4 13 15 2
35 10 9 1 15 15 3 13 1 14 13 3 0 1 0 2 13 3 0 9 1 0 7 13 9 2 1 10 9 2 1 10 9 1 9 2
19 10 9 4 13 15 1 14 13 1 9 12 9 0 7 13 10 9 2 2
5 11 11 13 15 2
4 10 0 9 2
10 9 1 11 2 10 1 9 0 9 2
19 15 13 11 9 2 10 0 9 2 0 1 9 2 13 10 0 11 11 2
5 15 13 12 9 2
20 7 10 9 1 11 12 4 9 10 13 3 0 16 15 13 14 13 9 10 2
8 2 1 15 13 10 0 9 2
20 15 13 10 0 9 16 15 13 2 15 13 1 9 9 12 2 7 13 9 2
24 9 13 0 1 9 15 13 16 15 13 0 1 10 0 9 7 12 9 4 13 15 1 9 2
9 0 9 13 2 0 9 1 9 2
12 3 13 9 2 7 13 1 1 10 0 9 2
15 1 13 3 9 2 9 7 0 9 15 13 15 1 9 2
22 15 4 13 0 1 2 1 9 1 9 9 2 7 1 9 13 15 3 9 13 3 2
27 9 15 13 1 1 9 2 9 15 13 3 1 10 0 2 0 9 2 7 15 13 15 0 14 13 9 2
25 15 13 0 1 1 9 2 13 15 1 9 2 13 15 1 1 10 9 7 13 3 3 1 9 2
12 0 13 15 3 2 13 15 7 13 1 15 2
6 3 13 15 0 2 2
7 15 13 12 9 3 3 2
5 11 11 13 3 2
5 15 13 1 11 2
8 2 8 8 8 8 8 8 2
8 8 8 8 8 8 8 8 2
10 8 8 8 8 8 8 8 8 8 2
12 15 13 1 9 1 11 11 2 11 2 11 2
7 1 10 0 9 13 15 2
4 10 0 9 2
4 11 11 13 2
2 13 2
46 2 15 13 1 0 2 13 3 1 16 15 13 10 9 2 13 3 7 13 1 10 9 2 15 13 0 2 13 1 2 13 1 9 1 8 1 9 2 3 13 15 1 7 13 9 2
9 15 4 13 3 1 12 9 3 2
5 15 4 13 9 2
10 15 13 1 10 9 2 9 2 9 2
6 15 13 1 1 15 2
4 15 4 13 2
2 9 2
7 0 2 0 2 0 9 2
8 15 13 9 2 15 4 13 2
10 2 11 13 10 10 9 2 13 11 2
6 2 10 9 1 9 2
12 9 2 9 2 9 2 9 2 9 2 9 2
8 3 1 10 9 13 11 11 2
4 9 10 13 2
17 9 10 13 10 0 9 2 7 0 13 15 1 1 10 0 9 2
9 15 13 10 9 1 1 11 9 2
6 15 13 3 9 0 2
4 3 3 9 2
11 0 4 15 13 1 10 9 1 9 10 2
6 2 3 13 15 15 2
7 1 9 3 2 13 15 2
8 2 3 13 15 15 2 11 2
5 15 13 10 9 2
14 1 14 13 11 11 9 2 4 15 13 12 9 1 2
16 15 13 9 15 13 1 10 9 7 13 10 9 0 11 9 2
4 7 10 9 2
9 10 9 13 15 1 9 1 9 2
10 2 8 8 8 8 8 8 8 2 2
13 15 13 0 9 2 0 9 1 10 0 11 9 2
23 10 0 13 16 15 3 13 2 3 13 2 16 15 4 13 1 2 8 8 8 8 2 2
13 9 11 13 9 11 2 16 15 13 0 1 15 2
12 1 10 13 11 2 15 4 13 10 0 9 2
15 10 10 9 4 13 0 9 1 1 9 2 7 13 9 2
9 2 3 13 9 15 13 1 9 2
5 10 13 15 2 2
17 11 13 10 9 2 13 15 2 10 0 0 9 2 10 0 9 2
5 15 13 9 12 2
5 11 13 12 9 2
6 15 13 1 10 9 2
16 2 10 9 4 15 13 9 1 11 2 3 1 11 11 11 2
10 2 15 13 0 15 13 2 13 9 2
8 0 13 0 9 10 1 9 2
12 10 9 1 12 13 15 10 9 1 11 9 2
6 9 13 3 1 9 2
9 11 13 16 15 3 13 1 9 2
7 9 1 13 15 10 9 2
4 1 10 9 2
6 12 9 9 10 9 2
9 7 9 2 12 9 7 12 9 2
28 15 13 9 1 9 1 9 2 13 1 10 9 1 3 1 9 2 10 9 1 9 2 7 10 9 1 9 2
8 15 13 1 9 7 13 9 2
5 15 13 0 9 2
13 15 13 9 1 10 9 16 15 13 15 1 9 2
4 10 9 13 2
9 0 0 1 11 9 13 10 9 2
17 1 9 4 15 13 1 11 2 1 9 4 15 13 0 1 11 2
25 11 13 1 10 9 1 11 7 13 16 15 13 14 13 10 9 2 16 9 13 10 9 1 15 2
11 15 13 0 7 0 14 13 9 1 15 2
8 1 12 13 9 14 13 0 2
22 2 15 13 0 3 2 15 13 1 9 0 1 14 4 13 2 1 3 14 13 0 2
2 0 2
9 15 13 0 9 3 2 10 9 2
8 9 16 15 13 12 1 12 2
11 11 13 1 16 15 13 1 15 1 9 2
13 9 13 10 9 1 15 2 1 14 13 14 13 2
14 15 13 3 1 12 9 2 15 13 1 9 1 9 2
15 2 15 13 10 9 1 0 9 1 9 2 9 7 9 2
34 9 13 10 10 2 10 15 3 13 1 10 0 9 7 9 1 9 15 13 2 7 0 1 9 7 9 15 13 16 15 3 13 15 2
8 15 13 10 9 1 9 2 2
10 1 9 2 11 2 9 1 0 9 2
7 9 13 1 1 11 11 2
17 15 13 9 1 9 2 0 9 2 10 0 9 2 9 1 9 2
12 2 15 13 1 14 13 0 9 1 15 10 2
5 1 9 7 9 2
10 15 4 13 10 0 9 1 9 10 2
37 15 9 4 13 15 2 13 16 15 13 14 13 0 2 15 4 13 1 10 9 1 9 2 7 15 13 10 9 1 16 15 13 3 14 13 9 2
9 15 13 3 16 15 3 13 15 2
8 15 13 3 0 1 10 9 2
4 16 15 13 2
16 15 13 10 9 9 1 9 4 13 1 10 9 1 10 9 2
17 11 13 16 10 9 13 1 10 0 9 15 3 1 3 4 13 2
5 15 4 3 13 2
16 15 13 1 2 13 15 1 1 10 9 7 13 1 10 9 2
12 7 10 0 9 0 13 10 9 1 9 10 2
4 15 13 9 2
7 11 9 2 9 1 11 2
16 2 16 15 13 10 0 9 1 9 2 13 15 15 3 0 2
20 2 15 13 15 1 0 9 1 9 2 13 2 13 9 2 13 10 0 9 2
20 2 14 13 10 9 1 10 0 9 13 12 9 9 7 12 9 9 7 9 2
27 0 9 13 15 1 9 2 0 9 1 10 0 9 16 15 13 3 15 4 13 15 1 14 13 9 2 2
15 2 3 13 15 0 2 7 3 13 15 9 7 13 15 2
5 0 15 15 13 2
18 2 3 1 9 13 9 14 13 1 15 2 15 15 13 10 9 1 2
16 10 9 1 9 2 10 9 15 13 2 10 9 7 10 9 2
28 15 13 1 10 0 9 2 1 9 7 9 1 9 7 3 9 13 14 13 9 1 14 13 7 13 0 2 2
13 1 9 13 11 9 2 15 13 0 9 1 15 2
3 9 12 2
4 15 13 12 2
14 0 9 1 9 4 13 1 16 15 13 1 1 9 2
11 11 13 10 0 9 15 13 15 1 9 2
8 15 4 13 1 9 1 11 2
17 1 9 13 15 15 0 2 13 9 1 12 9 1 10 0 9 2
5 10 9 1 9 2
12 16 15 13 1 13 3 9 1 9 1 11 2
11 15 13 15 13 9 2 7 15 13 0 2
11 9 13 1 16 15 13 10 9 0 9 2
4 11 11 11 2
9 2 10 0 9 13 15 1 9 2
22 10 0 9 15 1 10 0 9 2 1 9 1 9 2 4 13 15 1 9 0 9 2
11 2 1 9 12 13 15 1 11 1 11 2
13 15 13 12 2 0 1 9 13 15 1 1 9 2
5 15 13 12 0 2
3 9 13 2
6 11 4 13 15 1 2
2 11 2
6 15 9 1 0 9 2
9 15 13 10 11 11 1 9 3 2
8 7 10 9 0 2 0 9 2
10 2 15 13 10 9 11 15 4 13 2
8 7 3 2 10 9 1 9 2
27 10 3 0 9 2 10 3 0 9 11 2 10 9 11 9 2 11 11 2 10 0 9 2 10 11 9 2
11 2 15 4 13 7 9 7 9 1 9 2
19 15 13 10 0 9 2 13 15 1 1 9 1 1 9 1 10 0 9 2
3 2 9 2
7 9 10 13 1 10 9 2
5 7 9 13 0 2
17 7 9 10 2 10 0 2 13 3 9 2 15 13 0 1 9 2
10 2 15 13 12 9 2 9 1 12 2
10 10 9 13 0 2 10 13 12 9 2
21 16 15 4 13 10 9 9 13 15 15 2 16 15 4 13 0 9 13 15 15 2
8 7 15 13 10 0 9 3 2
3 13 9 2
5 9 10 13 0 2
4 15 13 0 2
21 2 8 8 8 8 8 8 2 8 8 8 8 8 2 8 8 8 8 8 2 2
8 15 13 0 1 15 15 13 2
18 2 15 13 12 2 12 9 2 15 13 16 15 13 10 9 1 9 2
13 15 4 13 1 11 11 1 9 1 9 10 9 2
15 13 3 16 15 1 9 13 10 9 15 13 15 0 9 2
8 2 11 2 2 4 15 13 2
13 15 13 14 13 0 0 16 15 13 1 1 9 2
15 15 13 9 1 10 9 2 13 9 1 9 2 13 9 2
17 2 15 4 13 10 9 15 0 9 13 1 9 1 1 10 9 2
9 3 13 3 15 1 15 15 13 2
6 15 4 13 10 10 2
5 1 9 7 9 2
11 11 11 13 3 1 11 11 1 10 9 2
19 2 7 10 9 3 1 13 10 9 3 2 1 10 0 9 1 10 9 2
25 9 1 14 13 9 2 9 1 14 13 2 2 2 16 15 4 13 9 7 0 13 7 13 0 2
13 2 15 13 9 1 9 12 7 9 13 1 9 2
5 10 9 11 13 2
9 10 9 4 13 0 1 9 10 2
14 10 9 4 13 1 11 10 9 1 14 13 15 13 2
9 2 10 9 13 15 2 13 11 2
10 2 4 15 0 13 15 2 13 11 2
8 2 15 13 11 2 13 15 2
9 11 13 3 3 13 1 10 9 2
7 2 15 13 15 13 9 2
10 13 15 13 0 2 13 9 7 13 2
8 11 11 13 9 1 10 9 2
12 15 13 12 9 1 9 16 9 13 1 9 2
12 9 1 13 11 15 1 9 2 3 1 9 2
6 15 13 0 1 9 2
7 1 9 1 9 13 15 2
18 15 13 10 0 9 2 10 0 9 1 9 2 9 15 13 1 9 2
29 2 1 9 4 15 13 1 10 0 9 1 10 10 9 16 15 13 1 3 1 9 1 1 9 7 10 0 9 2
7 10 11 2 10 11 2 2
22 1 9 13 15 0 2 1 10 9 1 9 13 15 15 0 7 13 9 1 11 11 2
6 11 13 9 1 15 2
9 11 4 13 11 11 2 1 9 2
7 1 12 9 13 9 3 2
6 2 15 4 13 15 2
8 15 13 9 15 4 13 1 2
18 2 15 13 15 13 1 9 10 2 13 15 1 9 1 3 14 13 2
11 15 15 13 13 10 9 9 1 0 9 2
17 9 2 9 2 9 2 9 2 9 2 9 2 0 9 3 2 2
14 11 13 9 2 13 1 1 10 12 9 9 1 9 2
22 1 12 12 1 9 1 9 2 7 9 16 10 10 9 13 2 16 15 13 10 9 2
5 15 13 1 11 2
12 2 15 13 0 1 9 11 2 2 13 15 2
12 2 10 10 9 13 1 10 9 1 9 10 2
5 15 15 4 13 2
4 9 13 1 2
3 11 13 2
16 15 13 1 15 10 0 9 16 15 13 15 7 13 1 9 2
9 11 13 0 10 9 1 9 12 2
9 15 13 1 9 1 10 0 9 2
11 10 0 15 13 9 1 13 9 7 9 2
19 7 9 13 0 2 1 0 9 15 13 1 12 9 15 13 1 1 9 2
15 15 13 1 9 10 10 9 2 13 1 9 2 7 13 2
10 2 6 2 3 13 15 1 11 2 2
8 9 1 13 15 1 9 11 2
9 1 1 9 13 15 9 7 11 2
7 11 13 1 10 0 9 2
12 2 14 13 1 11 7 11 13 1 10 9 2
4 15 13 0 2
23 2 9 15 13 16 15 13 1 15 11 13 16 15 4 13 1 9 16 15 13 3 2 2
7 11 13 2 13 0 9 2
7 11 8 11 13 1 15 2
8 0 4 15 13 10 0 9 2
4 10 0 9 2
58 2 15 13 10 0 9 2 14 4 13 1 10 0 9 2 4 15 13 10 9 0 9 15 15 3 13 2 13 9 13 1 9 7 13 10 9 2 2 2 7 13 9 9 2 13 9 13 10 9 1 15 2 13 9 1 9 2 2
6 15 4 3 13 0 2
18 15 4 13 9 2 4 13 7 13 1 9 2 11 2 11 7 11 2
9 15 13 1 10 0 9 1 9 2
6 15 13 3 1 9 2
11 1 10 0 9 1 11 13 15 9 13 2
14 9 2 9 2 9 2 9 2 9 2 9 2 9 2
16 2 9 13 15 9 2 10 0 9 2 15 13 3 0 2 2
18 1 9 1 9 2 16 15 13 12 2 13 9 1 9 1 1 9 2
4 15 13 9 2
16 2 15 4 13 1 1 9 2 7 3 4 9 7 9 13 2
11 15 4 13 10 9 14 13 1 9 3 2
12 16 9 13 1 9 2 13 15 3 1 9 2
8 9 13 15 9 1 14 13 2
14 2 15 13 15 1 9 16 15 3 13 9 1 9 2
6 15 13 3 10 9 2
4 15 13 15 2
4 15 13 15 2
8 13 9 10 7 13 1 9 2
8 3 9 4 13 0 3 15 2
11 2 15 15 13 4 1 0 9 13 15 2
9 15 13 16 10 9 13 0 1 2
6 10 9 2 10 9 2
8 9 1 10 9 13 0 1 2
24 15 13 10 9 1 9 15 15 13 14 13 1 9 2 9 7 1 10 9 1 9 1 9 2
11 15 13 1 1 10 9 9 2 13 15 2
10 7 1 10 9 10 9 0 9 2 2
6 15 13 9 1 9 2
9 7 10 9 13 15 1 1 15 2
16 15 13 3 0 1 16 15 1 9 3 4 13 9 1 9 2
15 1 9 1 9 13 15 1 9 1 9 1 9 1 11 2
10 10 0 9 13 0 2 1 0 9 2
14 7 15 13 2 13 2 13 9 7 9 1 9 3 2
18 0 1 10 9 3 10 9 1 9 4 13 1 9 1 14 13 9 2
12 1 1 9 1 9 1 9 13 10 0 9 2
17 16 15 13 1 1 14 4 13 1 10 9 2 13 9 1 15 2
8 2 1 3 13 15 15 3 2
9 15 13 15 3 0 1 9 2 2
4 9 4 13 2
13 11 13 15 0 1 15 15 3 13 1 14 13 2
13 2 15 4 13 1 9 2 1 9 15 13 15 2
12 15 4 13 1 9 2 7 13 1 9 3 2
9 15 4 13 9 1 14 13 9 2
13 15 13 1 9 10 7 13 1 1 10 0 9 2
20 2 15 4 13 14 13 15 1 10 9 1 15 15 4 13 14 13 10 9 2
32 15 13 10 0 9 1 9 10 2 2 2 16 9 0 13 10 9 7 10 9 7 3 13 15 1 10 9 15 13 1 9 2
10 2 15 13 14 13 15 1 15 10 2
3 13 9 2
7 13 1 1 10 10 9 2
10 15 13 15 16 15 4 13 10 9 2
4 7 10 9 2
5 15 13 14 13 2
8 0 1 9 2 0 7 0 2
3 0 9 2
11 1 9 7 9 13 10 0 9 15 1 2
6 15 13 1 1 9 2
7 11 11 2 11 2 11 2
18 2 15 13 1 10 0 7 0 9 1 9 1 9 15 4 13 1 2
11 15 13 10 9 2 10 10 2 13 11 2
22 2 15 4 3 0 13 15 1 10 0 9 2 9 1 0 9 7 9 1 9 2 2
10 15 4 13 12 9 9 10 0 9 2
9 15 13 16 15 3 13 12 9 2
30 2 7 10 10 9 15 13 0 1 11 11 13 3 9 7 10 9 14 13 10 9 1 9 1 10 10 1 9 2 2
6 11 4 13 0 9 2
15 2 11 2 9 15 3 13 1 15 10 7 15 0 13 2
45 15 4 13 1 15 10 1 0 10 9 2 13 15 1 10 9 2 15 13 3 10 9 4 13 2 1 9 1 10 9 14 13 9 1 14 13 2 7 10 9 4 13 1 9 2
22 7 3 13 15 16 9 3 4 13 1 9 1 10 9 2 3 1 10 0 9 2 2
11 1 9 1 9 13 15 1 11 1 9 2
20 9 13 16 15 4 13 15 1 11 2 11 13 15 13 16 15 4 13 0 2
15 1 10 9 4 15 13 10 9 1 0 9 7 13 15 2
7 11 13 1 14 13 1 2
14 10 9 15 13 1 1 9 2 13 9 0 1 15 2
5 15 13 7 13 2
16 2 15 4 13 0 1 9 10 7 3 13 9 1 15 2 2
17 15 13 1 16 3 10 9 4 4 13 1 16 15 3 13 15 2
6 11 13 1 1 9 2
6 9 4 13 1 9 2
10 15 13 1 9 1 9 2 1 9 2
2 1 2
5 15 4 13 15 2
4 11 13 0 2
18 2 10 9 13 10 9 1 16 15 13 1 1 10 9 2 13 15 2
31 2 15 13 3 10 9 2 9 1 14 13 1 10 9 7 10 9 15 4 13 1 1 10 13 16 15 13 9 1 15 2
21 14 13 1 9 1 15 10 1 0 2 0 9 13 1 0 1 14 13 0 2 2
14 11 13 1 10 0 9 7 13 9 1 10 0 9 2
8 2 15 13 1 10 0 9 2
18 15 13 1 9 2 13 10 9 1 15 3 0 15 15 4 13 15 2
8 15 4 13 15 15 15 13 2
7 7 15 4 13 1 15 2
6 15 4 13 9 10 2
9 2 15 13 15 1 9 1 9 2
7 12 9 2 7 12 9 2
5 15 13 9 13 2
3 15 13 2
12 15 13 16 15 3 13 1 14 13 1 3 2
7 15 13 15 1 10 9 2
18 15 13 2 16 15 13 15 1 1 9 2 1 14 13 15 1 9 2
10 15 13 3 3 0 2 16 15 13 2
11 11 11 13 2 8 8 8 8 8 2 2
5 15 13 1 9 2
3 0 9 2
5 15 4 13 9 2
13 10 0 9 9 2 10 9 2 9 1 10 9 2
16 12 9 1 0 9 7 10 9 1 0 9 2 13 1 15 2
14 2 15 13 15 3 2 13 11 11 2 1 0 9 2
8 2 13 15 3 2 13 9 2
11 15 13 9 2 9 13 14 13 1 15 2
8 1 15 4 15 13 15 13 2
19 2 9 1 9 13 10 0 9 1 9 10 2 15 13 14 13 15 0 2
7 3 13 15 0 3 2 2
10 10 9 13 10 9 15 15 4 13 2
19 10 9 1 9 4 13 15 0 1 9 2 1 10 12 9 0 1 9 2
6 15 4 13 1 9 2
8 2 9 10 13 0 2 0 2
2 1 2
10 15 13 15 3 2 4 15 4 13 2
9 10 0 9 1 11 13 15 1 2
4 15 13 0 2
16 15 13 16 15 4 13 0 9 2 13 7 13 15 1 9 2
5 11 13 1 9 2
21 15 13 1 11 11 2 9 1 11 2 10 12 9 15 13 15 4 13 10 9 2
9 15 13 0 2 7 9 10 13 2
5 13 1 1 9 2
6 9 13 15 1 15 2
12 10 9 1 12 13 15 15 1 1 9 9 2
9 15 13 15 1 9 2 1 9 2
14 1 10 12 9 13 15 9 2 1 10 0 10 9 2
5 11 11 13 3 2
7 1 9 4 15 13 9 2
5 2 15 13 1 2
7 2 15 9 4 15 13 2
6 13 15 0 1 9 2
8 15 13 15 15 4 13 15 2
21 9 15 4 13 1 2 0 9 2 9 15 4 13 1 2 15 13 1 11 2 2
6 2 3 4 15 13 2
9 2 10 0 9 13 15 1 15 2
9 15 4 3 13 1 14 13 3 2
7 15 13 1 10 9 2 2
11 3 13 15 1 10 9 16 15 13 0 2
10 3 13 15 10 9 1 7 13 3 2
3 15 13 2
8 10 9 13 1 7 13 15 2
4 15 13 1 2
9 2 15 4 13 10 9 1 9 2
11 9 10 13 3 2 1 10 9 1 11 2
15 15 4 13 10 9 1 15 15 13 1 11 2 13 15 2
7 15 13 16 15 4 13 2
5 15 13 1 9 2
6 10 0 9 13 9 2
8 15 13 1 9 1 9 12 2
47 2 8 8 8 8 8 8 8 8 8 2 8 8 8 8 2 8 8 8 8 8 8 2 8 8 8 8 8 8 8 8 8 2 8 8 8 8 2 8 8 8 8 8 8 8 2 2
6 3 13 15 1 9 2
18 2 8 8 8 8 8 8 2 8 8 8 8 8 8 8 8 2 2
11 2 15 4 13 1 15 2 13 11 3 2
5 2 15 13 0 2
4 15 7 15 2
19 15 13 9 1 14 13 9 2 1 14 13 1 7 13 9 7 13 9 2
11 15 13 0 0 16 15 3 4 13 15 2
11 3 13 15 0 16 15 4 13 1 9 2
13 15 13 9 1 11 1 3 10 0 1 10 9 2
6 2 15 13 10 9 2
2 9 2
8 15 4 13 14 13 9 10 2
11 13 1 1 9 1 9 2 1 0 9 2
6 9 4 3 13 0 2
12 15 13 15 1 2 13 0 1 14 13 9 2
5 2 3 2 11 2
4 15 13 11 2
11 4 15 4 13 1 9 2 2 13 15 2
10 15 13 1 11 2 1 10 9 11 2
8 15 13 12 9 1 11 11 2
10 15 13 3 7 13 1 9 1 9 2
5 15 13 1 9 2
7 15 13 16 15 13 9 2
13 2 15 4 13 9 10 1 16 15 13 1 9 2
11 15 13 15 1 14 13 15 15 4 13 2
9 15 13 1 9 2 10 0 9 2
14 7 3 13 15 9 1 10 9 1 9 10 1 9 2
6 6 2 15 13 15 2
3 13 15 2
7 15 13 3 10 0 9 2
14 15 4 13 15 1 14 13 0 1 9 2 13 15 2
3 15 13 2
9 2 15 13 0 1 2 15 13 2
20 15 13 1 1 9 2 13 1 10 0 9 2 13 0 1 1 9 1 9 2
9 2 15 4 13 10 9 1 15 2
10 9 1 16 15 4 13 15 1 3 2
13 15 13 9 1 11 2 16 10 1 10 9 13 2
9 15 13 1 11 11 2 1 11 2
7 13 10 0 2 7 13 2
9 15 13 9 15 13 15 1 15 2
4 3 13 15 2
10 2 8 8 8 8 8 8 8 8 2
14 8 8 8 8 8 8 8 8 8 8 8 8 2 2
9 11 13 16 15 3 13 1 9 2
9 2 15 4 13 9 10 9 1 2
9 15 13 1 11 2 1 9 3 2
13 16 15 13 14 13 0 2 7 9 13 2 13 2
6 3 13 15 1 2 2
4 3 13 15 2
10 10 9 4 15 3 13 10 9 1 2
21 15 13 1 9 1 10 9 2 15 4 13 12 9 2 7 15 13 15 3 0 2
8 10 9 13 15 9 1 9 2
12 2 9 7 9 2 15 4 13 1 9 2 2
6 2 15 13 1 9 2
16 2 15 4 13 9 15 4 13 2 13 2 13 2 13 2 2
5 15 13 10 9 2
16 15 13 14 13 2 3 15 13 16 10 0 9 13 1 9 2
8 15 13 9 2 7 0 9 2
9 9 13 1 10 0 9 1 15 2
11 15 13 10 0 9 1 9 10 10 9 2
15 2 7 2 13 11 2 15 13 0 14 13 15 0 1 2
2 1 2
11 15 4 3 13 1 2 13 1 0 9 2
5 15 13 9 1 2
20 16 15 1 0 9 13 16 15 4 13 1 2 13 15 1 10 9 1 15 2
9 2 15 13 9 10 13 10 9 2
16 16 15 13 10 9 1 1 9 4 11 13 1 10 0 9 2
9 15 13 15 1 15 1 10 9 2
11 2 15 13 3 15 15 13 15 4 13 2
15 9 15 15 3 1 0 10 9 4 13 1 2 13 3 2
22 16 15 1 10 9 0 9 13 1 1 9 2 1 1 10 0 9 1 9 0 9 2
4 1 1 9 2
29 16 15 13 1 13 15 1 10 9 15 13 1 9 1 9 1 11 2 9 15 13 15 1 14 4 13 9 1 2
6 15 13 1 15 10 2
19 3 4 15 4 13 9 1 16 15 13 10 0 9 14 13 1 1 2 2
12 15 13 14 13 9 2 13 9 2 13 9 2
9 3 13 15 1 9 1 10 9 2
5 15 13 1 11 2
16 1 14 13 2 11 11 1 11 11 2 8 8 8 8 2 2
12 2 15 13 0 9 1 15 15 4 13 15 2
7 15 4 13 9 1 15 2
12 15 4 13 10 9 1 10 9 9 3 13 2
26 16 15 4 13 0 9 2 13 15 10 9 1 9 2 1 9 2 13 15 1 1 10 9 1 9 2
5 3 13 15 9 2
4 9 7 15 2
8 15 13 1 9 1 15 10 2
17 3 13 15 9 1 9 1 9 2 15 4 13 0 9 1 11 2
13 2 15 4 13 1 9 2 9 2 0 2 9 2
11 15 4 13 1 15 2 1 10 0 9 2
19 3 15 16 9 10 4 13 10 9 2 7 15 4 13 9 1 14 13 2
22 15 13 9 1 1 10 0 9 1 9 2 15 13 15 2 15 13 10 9 15 13 2
6 15 13 9 1 15 2
7 9 13 0 0 1 11 2
5 11 4 13 9 2
9 2 7 15 13 15 14 13 0 2
8 13 15 1 10 9 1 11 2
3 2 6 2
2 0 2
2 0 2
2 0 2
2 0 2
2 0 2
2 0 2
2 0 2
2 0 2
2 0 2
8 1 9 4 15 3 13 15 2
15 15 4 13 1 10 9 2 15 4 3 13 9 1 9 2
10 0 3 13 15 0 0 9 15 13 2
12 9 13 1 15 2 13 15 3 0 1 11 2
5 9 13 3 3 2
9 2 15 13 9 10 2 13 15 2
11 2 15 4 3 13 0 1 14 13 9 2
3 13 15 2
9 2 13 15 10 9 3 1 9 2
3 15 13 2
15 2 6 2 15 13 12 2 11 11 2 10 9 1 11 2
12 15 13 3 1 9 1 10 9 1 11 11 2
30 16 15 13 15 1 9 3 4 13 1 1 9 0 2 1 14 4 4 13 1 2 13 15 15 1 3 15 4 13 2
3 11 13 2
20 15 13 15 1 15 15 13 1 11 9 1 11 2 7 10 12 9 1 9 2
13 2 15 13 0 9 1 14 13 10 9 15 13 2
9 7 15 13 3 0 1 9 10 2
19 15 13 1 10 9 2 13 9 2 13 1 9 2 1 11 2 1 11 2
11 2 10 9 4 1 7 1 13 9 3 2
2 0 2
17 15 13 1 9 15 4 13 1 11 2 15 13 15 1 0 9 2
24 2 9 15 13 1 11 11 16 15 4 13 9 7 13 1 11 1 14 13 9 1 9 10 2
12 10 9 2 7 10 9 15 4 4 1 11 2
9 7 10 0 9 15 13 1 9 2
14 15 13 1 10 9 11 11 2 10 0 9 7 9 2
5 2 11 13 3 2
9 4 15 13 9 2 11 8 2 2
7 15 13 0 1 10 9 2
14 15 13 15 1 16 15 13 0 14 13 0 7 0 2
6 15 13 3 13 0 2
16 3 1 2 16 15 13 1 9 2 13 10 9 1 10 9 2
4 9 13 15 2
3 15 13 2
9 1 1 10 0 9 2 13 11 2
13 2 15 13 0 14 13 1 16 15 4 13 9 2
10 15 13 0 3 2 16 15 3 13 2
10 15 13 0 1 0 9 1 10 9 2
11 7 1 7 1 13 9 1 11 1 15 2
18 11 11 13 10 0 9 1 15 2 15 13 12 9 16 15 3 13 2
8 13 0 1 1 2 11 2 5
11 11 13 15 1 2 11 2 1 11 12 2
2 9 2
19 3 4 15 13 11 11 13 2 11 11 11 2 1 11 9 2 11 2 2
14 11 4 1 0 9 13 0 9 1 2 11 2 9 2
31 15 13 3 3 3 0 16 11 3 13 1 1 2 11 2 2 10 9 15 13 14 13 10 15 9 13 2 7 0 1 2
22 2 11 2 13 3 1 14 13 9 1 2 11 2 2 0 7 0 1 14 13 9 2
18 3 3 13 15 1 9 7 13 1 1 9 1 9 15 13 1 9 2
32 15 13 1 3 0 15 13 14 13 9 2 7 1 2 11 2 13 15 3 9 1 14 13 1 10 0 9 1 9 1 9 2
19 15 4 13 10 9 15 4 13 2 7 13 1 9 7 0 9 1 9 2
34 3 3 13 2 11 2 0 0 1 1 9 2 3 16 15 4 13 1 0 9 15 13 1 11 2 7 15 4 3 13 10 10 9 2
28 7 15 13 1 10 9 2 10 9 7 1 9 1 10 9 2 4 15 0 13 0 9 9 0 1 1 9 2
35 9 1 15 13 16 15 3 13 9 1 1 9 2 7 16 0 3 13 16 15 4 13 1 10 9 2 4 9 13 1 1 10 9 0 2
38 2 11 2 7 13 7 13 0 1 2 7 0 16 11 13 14 13 1 1 9 7 0 0 9 2 13 3 11 9 0 13 0 1 2 11 2 9 2
7 10 9 4 13 12 9 5
10 11 1 11 4 13 0 9 1 9 2
18 9 2 11 11 2 4 13 10 1 9 0 9 1 10 9 0 9 2
15 9 4 1 3 13 9 1 0 12 9 3 10 0 9 2
3 13 9 5
28 11 11 13 9 1 10 10 0 9 11 2 15 13 16 2 11 11 2 13 9 15 13 9 1 10 0 9 2
20 9 13 3 11 2 15 13 10 10 9 15 13 1 10 0 9 3 1 9 2
10 15 4 15 3 3 13 10 9 1 2
20 9 2 9 2 9 7 9 1 9 4 13 1 9 1 16 9 4 13 1 2
19 11 13 3 0 9 2 1 14 13 16 15 13 10 0 9 13 1 15 2
3 0 9 5
19 11 11 2 9 1 9 2 13 16 9 1 10 0 3 13 1 14 13 2
10 1 1 1 9 1 9 4 9 13 2
18 9 1 10 0 0 9 4 13 9 3 0 16 9 3 13 10 9 2
18 9 11 13 16 10 9 4 13 2 0 1 14 4 13 10 0 9 2
19 11 13 3 0 9 2 1 14 13 16 15 13 10 0 9 13 1 15 2
10 0 9 13 3 9 1 9 9 9 2
16 9 13 16 9 4 13 2 1 10 0 0 7 0 0 9 2
5 12 9 1 9 5
6 11 11 13 1 9 2
17 11 11 13 1 1 9 1 9 0 9 1 10 0 9 1 9 2
37 15 13 1 12 9 1 9 0 2 7 4 4 13 0 1 12 9 1 9 1 14 4 13 15 1 1 10 12 0 15 4 13 1 10 9 9 2
10 11 4 3 10 9 13 1 11 9 2
11 15 13 10 0 9 9 1 10 0 9 2
12 10 9 1 10 0 9 13 3 9 1 9 2
16 15 13 3 14 13 1 9 7 13 1 14 13 9 1 9 2
14 1 10 10 9 1 12 9 3 13 15 1 12 9 2
10 3 13 15 3 12 7 9 1 9 2
23 15 13 1 1 9 1 10 9 1 9 12 2 16 1 9 12 4 15 13 10 0 9 2
34 1 9 12 13 15 3 1 9 1 9 10 9 2 7 3 4 15 13 3 0 1 1 9 2 7 3 0 9 3 14 13 1 9 2
8 2 13 1 13 1 0 9 5
5 2 11 12 2 2
3 0 9 2
16 1 10 9 1 9 11 11 13 15 0 1 2 11 12 2 2
35 16 10 0 2 11 2 9 13 1 9 1 11 12 2 4 15 13 3 0 15 4 13 16 9 4 13 1 1 0 0 1 10 0 9 2
24 0 1 0 9 2 0 9 7 0 9 2 13 3 9 0 14 13 1 1 1 9 1 9 2
17 0 0 1 9 11 11 2 15 13 1 1 10 0 2 0 9 2
26 3 15 13 3 15 14 13 1 1 1 9 2 15 1 9 13 15 1 10 0 9 1 9 1 9 2
2 11 2
34 1 10 0 9 1 0 9 2 16 15 4 13 0 0 9 13 1 11 9 1 11 11 2 4 9 13 0 1 0 0 9 7 9 2
42 0 1 15 10 13 16 15 4 13 9 1 10 0 0 9 2 7 15 13 15 3 1 14 13 1 1 14 13 9 1 15 15 4 13 10 1 10 0 9 3 0 2
15 1 10 9 4 15 13 16 9 4 13 0 0 1 3 2
35 1 10 9 13 15 0 10 0 2 0 7 0 9 15 13 15 13 1 1 9 1 10 9 2 3 13 15 3 0 9 1 10 0 9 2
29 3 16 15 3 4 13 1 15 12 9 1 10 9 13 9 7 9 3 0 16 15 3 13 9 1 14 13 15 2
27 15 13 10 9 1 10 0 2 11 2 9 2 7 15 13 15 9 11 4 13 1 7 13 1 1 9 2
30 15 13 0 9 2 7 0 0 9 2 7 3 16 9 13 1 9 1 0 2 13 0 7 0 0 9 1 1 12 2
19 9 13 15 1 9 1 9 2 15 13 1 12 9 13 0 1 15 0 2
39 15 13 1 1 10 0 9 2 7 13 13 10 0 9 13 9 1 9 0 1 0 9 1 10 9 2 10 0 15 4 4 13 13 1 1 13 0 0 2
25 0 0 13 3 9 16 1 12 9 4 13 9 15 13 0 1 9 1 15 11 11 13 1 9 2
22 2 11 12 2 13 0 1 10 0 7 0 9 2 15 13 1 13 1 9 11 9 2
8 6 2 6 2 6 2 11 2
7 9 1 2 11 11 2 2
27 11 4 13 0 0 1 9 1 11 2 7 1 15 13 1 15 10 9 15 3 0 13 3 0 1 9 2
28 9 1 10 9 13 16 15 15 0 13 0 0 9 3 4 13 15 0 1 9 15 0 0 4 13 1 9 2
21 1 2 11 11 2 4 15 13 1 10 9 16 15 13 16 3 0 4 13 3 2
27 3 13 15 1 10 9 10 9 2 16 15 4 13 15 15 2 15 13 15 13 1 12 9 1 0 9 2
4 13 0 1 2
16 3 2 15 13 3 0 15 16 15 4 13 3 9 13 1 2
26 16 15 3 13 10 0 9 14 13 9 1 2 13 10 0 1 14 13 1 0 9 7 9 1 9 2
22 15 4 13 1 10 9 9 1 14 13 9 2 7 10 0 4 0 13 1 12 9 2
2 0 2
12 3 2 13 15 2 15 4 13 1 12 9 2
4 0 7 0 2
23 16 15 7 10 9 13 1 9 2 13 15 3 0 14 13 1 15 15 13 1 1 9 2
26 15 13 0 0 14 13 0 2 7 16 10 0 9 13 1 0 9 7 0 9 2 13 15 3 0 2
12 13 16 2 11 2 9 11 11 13 1 15 2
18 6 2 13 3 9 0 9 2 1 15 15 13 1 2 11 11 2 2
6 13 11 11 1 11 5
11 9 13 9 12 9 1 14 13 15 1 2
8 11 11 4 13 1 10 9 2
7 9 13 15 1 10 9 2
24 10 12 9 0 9 13 15 13 15 0 1 10 9 16 15 13 10 0 9 1 9 11 11 2
23 2 9 9 2 10 0 9 2 13 15 0 10 11 1 11 3 15 13 16 15 13 1 2
24 1 14 13 3 0 15 13 15 2 13 15 15 10 10 9 12 9 2 13 11 1 9 11 2
12 11 13 0 16 15 13 9 1 9 1 12 2
10 1 9 13 15 1 9 9 1 9 2
10 0 9 1 0 2 11 8 11 2 5
6 9 13 3 1 9 2
22 15 4 13 10 9 9 14 13 1 0 1 9 1 10 0 2 11 8 11 2 9 2
43 3 13 9 2 11 1 11 2 11 2 3 0 1 10 0 9 1 9 2 3 0 13 15 0 16 9 1 11 4 13 16 15 0 3 13 0 2 7 13 9 7 9 2
23 9 13 2 11 1 11 2 11 2 2 7 3 13 15 7 9 7 9 2 3 1 0 2
7 13 9 0 2 0 9 2
20 2 11 1 11 2 11 2 13 1 9 1 2 11 2 7 2 11 11 2 2
27 15 13 16 15 3 13 10 0 2 0 9 14 13 15 1 2 7 9 9 13 1 7 0 0 1 3 2
25 15 4 0 13 1 10 0 9 1 9 1 9 2 7 15 4 13 1 9 2 9 7 0 9 2
17 1 0 4 15 13 7 13 1 10 0 9 3 15 15 13 15 2
20 1 13 3 9 1 0 9 2 7 1 0 13 15 3 0 15 15 13 0 2
16 15 13 9 1 14 13 9 10 9 1 9 15 13 0 0 2
28 9 13 3 10 9 1 2 11 11 8 8 11 2 2 7 15 13 0 2 3 15 1 9 13 1 10 9 2
32 4 15 13 0 2 11 1 11 2 9 2 4 15 13 15 0 3 2 15 13 10 0 0 15 4 13 2 11 2 0 0 2
26 7 10 0 9 7 0 9 13 1 3 15 13 15 2 7 3 4 15 13 15 0 0 1 9 9 2
3 0 9 2
5 1 9 1 9 5
16 11 11 13 10 12 0 9 1 9 15 4 13 1 1 0 2
5 15 13 10 9 2
4 9 9 12 2
18 0 11 11 13 0 1 1 10 14 4 13 10 9 1 11 1 12 2
3 0 9 2
32 9 2 9 1 11 0 9 11 2 13 10 0 0 9 2 11 8 2 8 8 2 8 8 8 8 8 2 8 2 8 2 2
2 9 2
12 1 10 9 1 11 9 13 11 11 9 10 2
6 15 13 12 9 0 2
2 9 2
17 11 11 2 3 9 1 11 11 11 2 13 10 1 11 0 9 2
14 2 15 13 9 15 13 9 7 9 10 2 13 15 2
3 0 9 2
28 1 14 4 13 1 1 0 1 12 2 1 9 0 9 1 9 2 4 15 13 7 1 9 7 10 0 9 2
2 0 2
35 1 14 4 13 11 8 8 11 1 11 1 12 7 12 9 1 12 9 1 11 2 13 11 10 3 0 9 1 11 2 3 12 9 0 2
20 15 13 10 9 15 13 9 1 0 9 1 10 0 9 2 7 9 1 9 2
5 12 9 1 9 2
10 11 13 9 2 9 7 9 1 11 2
2 9 2
37 11 11 11 4 13 1 9 1 14 13 9 1 11 1 14 13 9 0 9 2 9 11 13 2 1 11 11 11 2 1 10 9 1 9 1 9 2
12 15 13 10 9 9 7 16 9 4 13 9 2
2 1 2
17 1 10 9 1 9 11 13 11 10 12 0 9 1 10 0 9 2
5 13 0 1 11 2
33 1 9 9 4 15 1 9 1 9 1 11 11 13 11 0 9 2 13 1 11 11 1 11 7 13 1 11 11 0 9 1 9 2
10 15 13 1 9 3 15 13 9 10 2
5 9 13 1 11 2
16 9 13 1 9 2 1 10 9 15 0 13 0 7 3 3 2
11 13 15 10 9 1 11 11 2 10 9 2
13 13 15 10 9 1 3 15 13 15 2 0 1 2
5 15 13 1 9 2
15 3 13 2 11 2 11 8 8 8 8 8 8 8 2 2
7 10 9 13 1 2 0 2
10 11 13 10 0 9 1 10 9 3 2
5 9 0 9 12 2
26 15 13 1 10 1 10 12 9 3 1 2 1 10 1 9 2 3 1 9 2 7 1 3 1 9 2
13 15 13 2 13 15 7 13 15 1 10 0 9 2
5 15 13 3 0 2
11 15 13 15 15 13 3 0 2 13 15 2
9 8 8 8 2 8 2 13 15 2
11 15 13 3 1 9 2 10 9 9 9 2
10 15 4 4 13 15 1 1 10 9 2
25 1 9 2 9 0 9 2 4 15 13 0 1 9 1 10 0 9 1 9 1 10 9 1 9 2
24 15 13 3 2 1 10 9 2 7 13 1 3 15 4 13 3 0 1 9 1 11 0 9 2
4 0 9 0 2
5 15 13 3 12 2
5 1 9 1 9 2
14 15 13 10 0 0 9 1 9 1 10 0 9 11 2
8 9 4 13 15 1 10 9 2
4 15 13 0 2
7 3 4 15 3 13 15 2
18 11 4 1 7 1 13 1 1 15 1 14 13 9 11 8 8 11 2
6 15 13 10 0 9 2
9 10 9 4 3 13 1 0 9 2
3 9 12 2
24 15 13 9 1 9 1 11 9 2 13 7 13 1 9 10 9 1 9 15 3 13 7 13 2
16 1 10 9 13 15 1 11 11 9 2 3 1 9 0 9 2
17 15 13 15 1 9 1 9 1 11 2 3 1 11 2 7 9 2
16 11 2 0 2 0 7 0 1 9 2 13 3 0 7 0 2
10 15 13 10 0 9 7 0 7 0 2
23 11 4 13 10 3 0 0 9 2 10 0 0 9 15 13 9 1 12 9 9 1 9 2
24 0 9 4 13 1 1 15 2 7 1 9 12 13 11 1 1 9 12 1 11 11 11 11 2
4 9 13 0 2
14 3 3 4 15 13 9 2 15 4 13 10 0 9 2
11 7 10 10 9 4 13 15 1 10 9 2
26 1 10 9 13 11 1 10 0 9 2 7 15 4 3 13 1 11 0 16 15 4 13 1 9 9 2
9 9 11 11 4 13 1 1 9 2
4 11 13 0 2
12 1 10 9 13 10 9 9 1 9 1 11 2
12 2 11 2 3 13 15 16 15 4 13 9 2
3 13 11 2
10 2 1 10 9 2 9 2 13 11 2
12 2 3 13 15 16 15 4 13 10 9 9 2
4 13 9 3 2
8 2 1 10 9 2 13 11 2
13 2 7 3 13 15 14 13 15 1 10 0 9 2
3 13 9 2
23 15 13 11 11 2 10 1 11 0 9 10 9 2 10 0 0 2 9 7 9 1 11 2
5 15 13 1 9 2
22 16 15 13 15 2 13 11 1 16 15 13 11 1 0 9 2 1 9 11 1 12 2
10 2 15 13 3 3 3 15 15 13 2
6 10 9 0 13 15 2
2 9 2
16 15 13 0 0 2 15 4 13 10 9 1 15 1 3 15 2
10 7 15 13 1 10 9 1 10 9 2
9 15 13 9 1 14 13 15 3 2
22 16 15 13 9 2 13 15 3 12 7 1 9 3 15 13 14 13 16 15 13 0 2
22 11 13 0 0 1 14 13 10 0 9 2 7 1 9 10 13 15 14 13 15 1 2
13 0 9 13 11 1 10 9 1 11 7 13 11 2
12 2 15 13 0 1 9 15 13 1 11 11 2
4 16 13 15 2
6 1 0 9 3 0 2
3 2 9 2
11 15 13 15 13 1 9 1 9 9 2 2
4 9 1 15 2
9 10 9 1 15 2 10 9 0 2
13 3 16 11 1 9 13 2 13 11 9 15 0 2
17 15 13 1 11 9 7 9 7 13 10 0 0 9 1 10 9 2
6 15 13 15 0 9 2
7 2 11 13 15 3 2 2
5 11 13 1 9 2
15 2 15 13 1 9 2 15 13 3 0 9 0 1 15 2
14 7 6 2 15 4 3 13 0 1 10 10 0 9 2
7 11 13 11 11 1 12 2
9 2 15 13 12 9 9 1 15 2
15 15 13 3 14 13 9 7 13 10 9 0 1 9 2 2
6 1 10 9 13 11 2
23 2 16 15 3 4 4 13 1 10 9 1 15 13 1 14 13 1 10 9 1 10 9 2
10 11 11 13 10 0 2 9 2 2 2
7 11 11 13 11 13 9 2
31 2 3 16 15 13 10 9 1 14 4 13 2 13 15 3 11 15 14 13 1 1 15 1 9 2 9 7 0 0 9 2
20 15 13 1 16 15 13 14 4 13 1 14 13 0 1 9 16 13 1 9 2
3 15 13 2
19 2 15 13 0 3 15 13 3 1 15 2 15 13 16 15 13 0 3 2
5 15 13 0 2 2
9 1 12 13 11 0 14 13 1 2
21 2 15 13 15 4 13 16 15 4 13 9 1 11 7 13 9 1 1 0 9 2
15 15 4 13 15 1 16 15 13 0 3 1 14 13 15 2
21 9 13 16 10 9 4 13 0 2 3 16 11 4 13 1 1 9 1 10 9 2
5 3 13 15 3 2
12 11 9 13 15 3 16 15 13 9 10 0 2
8 15 4 0 1 10 0 9 2
7 9 13 1 0 1 0 2
9 10 9 13 11 11 1 11 9 2
10 11 13 14 13 9 7 11 13 3 2
13 15 13 9 1 9 2 15 13 7 13 9 1 2
4 9 4 13 2
12 15 13 1 12 9 7 0 12 9 1 11 2
21 16 11 11 13 2 13 9 16 9 1 11 13 15 15 13 0 1 1 10 9 2
5 11 4 13 15 2
19 2 3 13 9 11 13 15 2 15 15 13 2 0 2 3 0 0 2 2
32 15 13 3 0 2 3 10 9 2 7 4 3 0 1 13 1 10 10 9 2 10 0 0 9 4 13 2 1 9 1 9 2
7 2 15 13 15 13 9 2
3 2 6 2
13 15 13 9 15 0 13 9 7 9 1 11 11 2
9 15 13 9 1 10 9 1 9 2
35 15 4 13 10 9 1 9 2 1 9 1 2 0 1 1 10 9 7 0 1 9 2 9 1 9 2 9 13 9 7 13 9 1 15 2
17 15 13 0 1 0 9 7 13 15 1 15 15 13 1 0 0 2
9 16 13 1 9 1 10 0 9 2
7 15 13 0 1 10 9 2
18 15 4 13 1 9 1 9 1 9 1 14 4 13 1 9 1 9 2
6 15 13 15 1 9 2
8 2 11 13 0 9 1 9 2
22 16 15 13 1 7 13 15 13 1 0 9 2 13 15 1 1 14 13 1 0 9 2
11 15 13 15 0 1 15 14 13 0 9 2
11 0 13 11 1 10 12 9 1 10 10 2
19 1 14 4 4 13 1 11 2 13 11 11 15 2 10 9 3 1 9 2
16 12 9 1 16 15 13 1 12 9 9 2 13 9 12 9 2
6 10 9 13 10 10 2
11 9 13 0 1 10 9 15 3 4 13 2
7 12 9 1 3 0 9 2
4 10 0 9 2
17 1 11 1 12 2 1 11 11 2 11 11 2 11 11 7 11 2
12 11 11 2 11 2 11 9 4 3 13 0 2
30 1 1 9 15 4 13 1 9 2 0 9 12 2 10 9 3 9 13 3 0 1 11 16 9 1 11 11 4 13 2
9 9 10 4 13 1 11 1 11 2
15 1 14 4 13 1 9 1 11 2 13 15 15 1 12 2
13 15 13 1 9 1 11 7 9 11 1 10 9 2
11 9 4 3 13 1 1 10 9 1 11 2
27 15 13 1 11 2 13 1 1 10 0 9 2 3 1 1 10 0 0 9 2 15 13 15 1 9 11 2
10 15 13 3 11 13 16 15 13 12 2
6 15 13 12 9 3 2
8 9 2 9 7 9 4 13 2
22 15 13 1 10 0 9 2 13 9 15 13 1 9 7 15 4 13 11 9 1 15 2
4 1 11 11 2
6 1 9 3 13 15 2
4 1 11 11 2
3 15 13 2
9 13 11 9 1 10 9 1 9 2
9 15 13 3 9 1 9 4 13 2
19 15 13 10 3 0 9 3 2 1 10 12 9 9 1 9 7 0 9 2
7 9 13 9 1 9 10 2
18 9 11 13 9 1 10 0 9 2 3 11 13 10 0 9 1 9 2
23 3 16 9 11 13 1 9 3 7 3 2 13 3 10 10 0 9 1 9 1 9 9 2
10 9 13 16 7 11 7 11 13 0 2
13 11 4 1 7 1 0 4 13 1 14 13 0 2
22 1 11 7 11 9 11 2 12 9 0 1 11 2 13 11 10 2 0 0 9 2 2
19 15 13 15 1 1 9 1 9 7 13 2 1 16 15 4 13 1 9 2
20 16 15 13 12 7 12 2 13 15 1 9 10 7 13 0 9 1 1 9 2
11 10 0 13 1 0 9 2 1 11 9 2
26 11 11 13 1 10 0 9 7 9 13 9 12 1 9 2 1 10 9 15 13 10 9 1 11 9 2
9 9 13 10 0 9 0 1 9 2
9 11 4 13 10 9 2 13 11 2
18 15 13 11 11 2 11 0 0 9 2 15 13 3 1 11 1 11 2
20 2 15 13 0 1 15 2 10 0 9 1 10 9 2 16 15 13 1 11 2
7 10 9 0 13 15 9 2
10 15 13 3 0 2 10 0 9 10 2
12 15 13 0 0 2 10 9 15 13 1 15 2
12 15 13 0 16 15 13 9 15 11 3 13 2
10 15 13 3 9 14 13 15 1 9 2
13 7 15 13 3 3 11 15 4 13 15 1 11 2
10 15 13 3 15 13 10 9 1 11 2
13 16 15 4 13 2 13 15 0 3 0 1 15 2
11 15 13 15 15 13 15 1 9 1 15 2
9 15 13 3 3 1 1 10 9 2
6 3 13 15 3 9 2
13 15 13 0 0 15 16 15 13 15 15 4 13 2
9 3 16 15 3 13 0 1 11 2
11 15 4 13 16 15 3 13 9 1 11 2
7 3 13 15 3 10 1 2
11 15 4 13 1 10 10 9 2 13 11 2
11 15 13 1 1 11 11 11 1 11 11 2
9 10 9 13 10 9 15 13 11 2
6 15 4 3 13 0 2
13 2 11 13 14 13 1 9 2 15 13 10 9 2
5 7 15 13 9 2
17 15 13 15 0 0 3 2 7 9 13 15 15 13 15 1 15 2
6 7 15 15 13 3 2
7 11 4 13 9 1 11 2
4 15 13 15 2
10 6 2 15 13 3 0 15 15 13 2
8 9 11 1 10 0 9 13 2
5 9 13 0 3 2
15 7 11 7 9 11 13 0 1 9 1 16 15 13 1 2
6 3 4 15 13 9 2
8 1 12 13 11 0 1 9 2
17 15 13 0 0 1 16 10 12 9 0 0 9 15 4 13 9 2
17 2 15 13 15 0 16 15 3 4 13 1 9 1 14 13 15 2
14 15 4 13 10 0 1 14 13 16 10 9 13 3 2
22 15 13 15 1 14 13 10 9 7 13 1 1 9 2 2 13 11 1 9 11 12 2
15 9 1 11 0 9 11 11 13 1 9 2 0 9 12 2
14 2 15 13 15 3 13 10 9 1 9 2 13 11 2
9 2 11 11 4 0 13 15 1 2
14 15 4 3 13 10 0 9 15 4 13 1 14 13 2
11 15 13 15 1 13 15 9 1 10 9 2
9 15 13 15 14 13 10 0 9 2
20 16 15 13 1 1 0 2 4 15 13 1 10 10 0 9 2 0 10 9 2
13 2 8 8 8 8 8 8 2 2 13 9 11 2
19 1 10 9 13 15 16 15 3 4 13 1 1 10 9 1 10 0 9 2
8 11 11 13 3 0 11 13 2
14 2 15 13 0 0 15 1 16 11 13 9 1 15 2
4 0 0 15 2
12 11 13 15 0 2 7 11 13 3 1 15 2
22 15 13 16 15 3 13 1 16 15 13 1 2 7 9 1 10 0 9 13 15 0 2
20 15 13 16 10 0 9 2 15 3 4 13 1 9 1 9 2 4 13 0 2
30 3 11 11 2 10 0 9 2 13 1 9 16 2 10 9 13 10 9 1 10 0 9 2 0 2 0 7 0 2 2
8 11 4 13 0 1 0 9 2
11 0 13 0 1 1 15 2 3 0 9 2
9 2 0 13 10 9 1 9 2 2
8 2 15 13 0 0 1 9 2
10 15 13 10 0 0 9 2 13 11 2
9 10 9 13 0 1 1 11 11 2
12 2 10 9 13 7 0 1 11 10 7 9 2
10 15 13 0 7 13 9 1 9 2 2
3 11 13 2
30 2 3 16 15 13 16 15 13 15 0 1 9 2 13 15 16 15 13 0 9 2 7 15 13 9 1 9 1 9 2
19 1 16 15 3 13 9 1 15 2 13 15 3 16 15 13 0 0 9 2
11 15 13 1 10 9 15 13 1 11 11 2
2 12 2
5 15 13 3 0 2
23 2 15 13 0 15 4 13 15 14 13 1 15 4 13 0 1 1 15 15 13 1 15 2
28 16 15 4 13 1 1 9 7 13 15 15 13 0 2 13 9 7 13 13 2 4 9 13 0 1 10 9 2
29 7 16 11 11 13 2 0 7 1 2 2 7 9 13 2 13 15 15 4 13 9 1 16 10 9 13 1 2 2
33 14 13 1 1 11 11 13 15 10 0 9 9 2 7 15 13 15 4 13 0 9 1 10 15 13 16 15 4 13 1 1 9 2
17 2 15 4 13 2 2 13 11 2 2 16 9 13 0 0 9 2
7 15 13 1 9 1 9 2
15 7 16 15 13 15 10 1 9 2 13 15 0 1 9 2
14 15 13 15 13 3 1 14 4 13 1 1 9 2 2
32 15 13 1 11 1 12 2 7 13 3 9 1 9 2 3 1 11 2 10 1 0 9 15 13 0 1 14 13 15 10 9 2
17 15 13 12 9 1 12 9 2 7 13 1 11 1 11 1 12 2
20 3 4 15 13 1 14 4 13 14 13 10 0 9 1 10 9 1 10 9 2
22 15 13 1 9 1 11 2 11 11 7 3 1 11 2 3 15 13 9 7 13 9 2
4 15 13 1 2
23 1 12 13 15 1 11 1 14 13 9 1 11 1 10 9 1 12 1 12 9 0 9 2
5 15 13 10 9 2
7 9 13 15 1 10 9 2
9 11 13 15 16 9 4 13 0 2
3 10 9 2
5 11 13 10 9 2
10 15 13 9 1 1 10 9 1 9 2
5 15 13 15 0 2
7 10 9 15 13 1 15 2
15 9 4 13 1 16 11 0 13 1 7 13 10 1 9 2
11 9 13 1 11 9 2 1 9 1 9 2
9 9 13 1 9 1 11 9 1 2
6 9 13 0 1 9 2
16 9 4 13 3 2 7 15 4 3 13 10 0 2 13 11 2
23 0 9 2 12 9 0 2 13 9 1 1 11 9 1 14 13 9 1 9 7 9 10 2
11 11 13 1 2 1 0 13 1 1 11 2
11 9 4 13 1 2 0 9 0 9 2 2
11 3 4 0 9 13 9 1 9 1 9 2
21 0 9 13 3 16 15 4 13 12 9 1 9 2 7 13 10 9 15 3 13 2
16 1 14 4 13 1 11 2 13 11 1 10 0 9 1 11 2
12 15 13 10 9 9 11 1 14 13 15 0 2
23 16 15 13 1 11 1 14 13 14 13 10 9 1 9 1 16 15 13 9 1 10 9 2
11 7 10 9 13 0 2 7 13 3 1 2
19 10 9 15 11 4 13 2 13 10 9 1 9 11 1 9 1 11 11 2
15 0 1 3 0 1 1 9 9 9 13 15 2 13 15 2
11 2 15 13 3 1 16 9 3 13 0 2
17 15 13 9 1 0 9 3 2 7 1 2 15 13 15 3 0 2
9 15 4 3 13 15 1 15 13 2
15 15 4 13 15 3 0 1 1 2 7 0 7 1 9 2
13 11 13 0 3 1 14 13 1 10 12 10 9 2
8 15 13 10 0 9 3 2 2
6 15 13 10 0 9 2
10 10 9 13 11 11 0 1 10 9 2
9 9 11 4 3 4 13 1 9 2
16 11 2 3 9 2 9 7 9 1 9 2 4 13 1 9 2
11 12 9 1 11 9 13 15 1 10 9 2
12 2 3 16 15 13 9 2 13 15 10 9 2
7 9 1 0 9 13 3 2
21 15 13 15 13 2 15 4 13 16 15 13 11 2 7 15 13 3 14 13 9 2
8 15 13 3 1 9 7 13 2
9 2 6 2 15 13 15 3 2 2
13 15 13 10 9 1 1 11 8 11 11 8 11 2
20 10 9 2 9 11 2 13 1 10 2 9 2 9 7 9 1 14 13 2 2
15 9 7 9 13 1 15 2 15 13 11 9 9 7 9 2
14 2 14 13 11 2 15 13 10 0 9 2 13 11 2
11 2 15 13 15 13 15 1 9 1 9 2
4 15 13 0 2
10 15 13 16 9 13 3 0 1 15 2
11 7 3 2 1 10 9 2 13 15 15 2
13 3 13 15 15 3 1 14 13 1 9 7 9 2
8 7 10 0 0 9 15 13 2
8 15 13 3 0 1 14 13 2
10 10 0 9 1 0 9 13 9 10 2
13 3 15 13 9 1 0 9 15 3 13 0 1 2
20 7 16 15 13 15 16 15 4 13 0 1 14 13 9 2 4 15 13 9 2
11 11 11 4 3 13 15 15 4 13 11 2
5 2 15 4 13 2
13 16 9 3 13 1 9 2 13 15 3 10 9 2
30 15 4 13 12 9 0 1 9 15 13 9 3 15 13 9 10 16 4 13 9 1 16 15 4 13 3 1 10 9 2
15 15 13 15 3 0 16 9 3 13 10 0 9 1 15 2
16 1 15 15 13 13 15 10 9 15 4 13 16 15 13 11 2
6 15 13 10 0 9 2
6 15 4 3 13 15 2
5 7 15 13 0 2
10 2 13 15 16 15 4 13 1 9 2
14 2 15 13 10 9 15 4 13 10 15 1 10 9 2
20 15 13 15 16 15 13 10 9 16 15 13 1 14 13 15 16 15 13 9 2
6 2 7 15 13 15 2
9 2 15 13 10 0 9 1 9 2
15 7 15 13 0 9 1 9 1 0 9 7 10 0 9 2
11 15 15 13 1 2 13 15 3 0 1 2
16 0 15 13 11 1 9 13 3 2 10 0 9 1 9 2 2
26 15 13 1 0 11 11 2 12 9 15 13 3 1 15 2 9 16 15 4 13 2 10 0 9 2 2
4 3 4 13 2
13 15 2 13 15 16 15 13 9 1 10 0 9 2
20 15 13 3 1 1 10 9 15 4 13 1 7 13 9 10 2 2 13 15 2
4 10 9 13 2
6 2 15 13 0 0 2
9 4 13 10 0 9 1 9 2 2
38 0 9 1 10 9 4 15 13 10 9 2 1 11 11 11 2 9 13 10 9 15 1 9 1 9 13 9 7 9 1 9 1 0 9 2 9 2 2
13 9 9 11 11 11 13 1 16 15 13 1 9 2
17 2 11 13 1 9 1 9 7 9 2 7 1 9 13 9 15 2
13 0 3 13 15 15 1 16 9 13 12 9 2 2
13 11 9 2 0 10 9 2 13 1 9 1 9 2
14 9 13 1 9 2 15 4 13 1 10 9 1 9 2
13 2 15 4 13 16 15 3 13 10 0 9 0 2
14 15 13 0 9 1 15 7 10 9 13 15 1 9 2
8 16 15 13 9 2 13 15 2
7 2 3 13 7 13 2 2
15 7 15 13 16 15 3 4 4 13 0 16 15 13 0 2
17 15 13 3 14 13 10 9 7 10 9 0 9 7 9 2 2 2
12 11 13 10 11 15 15 13 4 13 15 0 2
8 15 4 1 9 13 9 2 2
16 2 10 9 1 9 1 11 9 4 15 13 3 2 9 2 2
9 9 13 1 7 1 1 10 9 2
28 8 8 8 8 8 8 8 2 13 11 11 2 7 13 15 1 9 1 15 15 13 1 10 2 0 9 2 2
16 3 12 7 12 1 0 0 9 9 1 9 13 0 1 15 2
6 15 13 1 11 11 2
14 2 11 13 10 0 7 0 9 15 13 1 1 9 2
13 15 4 13 1 9 2 13 1 1 9 7 9 2
7 15 4 0 13 0 9 2
11 15 13 1 10 0 9 2 13 11 0 2
8 15 13 12 9 1 11 9 2
6 15 4 13 1 3 2
27 2 15 13 0 16 15 13 10 9 3 9 3 3 13 15 0 3 1 16 15 13 9 16 15 13 1 2
12 11 4 0 2 7 0 13 1 9 1 9 2
9 15 13 1 10 9 0 1 11 2
10 7 15 13 10 0 0 2 0 9 2
11 11 4 13 0 0 1 14 13 1 9 2
10 10 1 9 3 4 13 0 7 0 2
21 15 4 13 1 1 14 13 11 1 14 13 1 1 10 0 9 1 15 1 9 2
15 15 4 13 10 9 2 1 9 2 9 2 9 1 9 2
21 15 4 13 10 9 2 10 9 16 10 9 13 10 10 1 10 9 2 1 9 2
8 2 7 2 13 11 7 13 2
6 2 11 13 3 0 2
9 9 13 10 0 9 9 1 9 2
8 9 4 13 1 1 10 0 2
14 0 0 13 15 1 1 9 2 15 13 15 3 0 2
13 7 0 0 0 9 13 1 9 1 9 1 9 2
18 13 11 11 9 15 4 13 15 3 4 13 10 0 9 1 9 10 2
8 0 16 11 13 15 13 3 2
19 15 13 0 9 2 0 9 7 9 1 9 7 9 15 13 1 0 9 2
12 9 4 3 4 13 1 14 13 9 15 13 2
12 2 13 15 10 9 10 9 4 13 1 3 2
7 2 1 10 10 12 9 2
11 15 13 10 0 0 9 2 7 15 13 2
11 7 3 13 15 0 1 16 15 4 13 2
10 2 7 3 13 15 3 15 1 2 2
8 15 13 3 1 10 10 9 2
10 2 0 9 13 9 1 9 7 9 2
19 15 13 3 1 3 9 11 13 12 9 9 1 9 1 16 15 13 1 2
7 10 1 9 13 1 15 2
22 2 15 13 3 15 4 13 3 0 9 1 9 7 9 2 7 15 13 0 1 9 2
9 15 4 13 1 1 10 11 8 2
7 10 9 4 4 13 2 2
13 0 9 13 0 1 0 9 1 14 13 10 9 2
12 7 3 9 13 0 9 13 0 1 10 9 2
32 9 11 11 13 1 0 9 16 15 4 4 13 1 12 0 9 15 4 13 1 9 1 14 13 10 9 1 10 9 1 0 2
17 1 0 9 4 9 3 4 13 1 9 1 14 13 15 0 9 2
17 10 0 9 11 13 15 4 13 1 10 0 9 15 13 0 0 2
4 0 13 15 2
9 2 14 13 1 4 13 9 2 2
27 3 15 13 9 2 9 15 13 10 0 9 1 9 2 1 9 1 0 9 7 9 1 9 1 0 9 2
15 2 9 13 9 4 4 13 16 9 13 1 2 13 11 2
10 1 9 13 9 0 9 1 9 9 2
8 11 0 9 11 13 15 3 2
10 2 10 9 4 3 13 10 9 9 2
8 9 4 3 13 1 15 2 2
23 11 11 4 1 9 13 14 3 13 10 9 1 9 2 1 9 1 14 4 13 1 0 2
3 11 11 2
2 11 2
3 11 11 2
9 15 4 4 13 1 9 7 9 2
9 1 3 14 13 1 11 11 11 2
18 9 1 9 7 9 13 15 1 9 1 15 2 13 15 1 10 9 2
19 16 11 11 13 0 9 2 7 13 0 13 1 9 1 9 2 13 9 2
12 15 13 1 16 15 13 1 9 1 10 9 2
21 2 15 13 1 9 15 13 1 9 7 15 13 15 0 16 15 13 1 1 9 2
13 15 13 15 13 1 14 13 10 9 3 1 9 2
12 10 9 1 11 13 15 1 14 13 10 9 2
7 10 9 1 9 13 15 2
8 15 13 3 0 1 12 9 2
19 2 8 8 8 2 8 8 8 8 8 8 8 2 2 13 15 1 15 2
6 10 9 13 15 2 2
21 7 15 13 11 11 9 2 1 10 0 9 7 10 9 1 0 9 1 11 11 2
5 15 13 1 11 2
12 2 9 10 13 1 9 2 15 13 0 2 2
4 3 13 11 2
5 11 4 3 13 2
26 15 13 11 11 11 8 8 11 11 2 10 1 0 0 1 9 9 15 4 13 9 1 9 7 13 2
21 2 15 4 13 1 9 1 10 9 15 13 9 1 11 2 7 9 1 10 9 2
22 1 10 15 13 15 0 1 1 9 2 4 9 13 10 0 7 0 9 2 13 15 2
16 11 11 2 9 15 3 13 9 2 13 15 3 2 1 11 2
6 3 13 9 1 11 5
3 0 9 2
23 9 7 0 9 1 9 13 1 2 9 2 1 9 7 9 1 11 9 2 1 0 9 2
3 0 9 2
24 9 1 9 1 10 9 1 9 1 11 11 4 1 0 9 13 1 10 0 9 2 1 9 2
9 9 2 11 11 2 11 5 11 5
32 1 10 9 13 1 11 8 11 11 13 15 1 3 10 0 2 7 0 9 1 2 9 2 13 9 1 9 1 10 0 9 2
17 9 13 1 0 9 1 0 9 2 7 9 1 0 9 7 9 2
28 2 9 2 13 1 9 1 1 14 13 9 10 0 9 1 0 9 13 1 2 7 13 9 1 9 1 9 2
23 10 9 13 1 11 11 1 9 12 13 16 12 9 1 11 9 13 10 0 9 1 9 2
8 1 9 12 13 9 12 9 2
3 11 9 5
14 9 1 9 13 1 9 1 1 12 9 7 10 9 2
10 1 15 13 11 11 7 10 11 11 2
27 11 13 10 1 10 0 9 11 11 11 0 13 1 1 10 12 9 0 9 15 4 13 1 9 0 9 2
23 11 9 13 1 15 15 1 12 7 12 13 1 12 9 9 1 0 9 1 12 0 9 2
17 11 11 11 2 15 13 0 9 1 0 9 2 13 1 10 12 2
12 2 15 13 1 16 9 13 1 0 0 9 2
35 7 15 13 0 16 0 9 13 1 1 9 11 11 2 15 3 4 13 10 0 9 14 13 1 13 11 11 2 9 15 13 0 9 0 2
21 2 15 13 10 9 16 10 9 13 1 7 4 13 1 9 1 14 3 13 15 2
25 9 10 4 3 13 2 7 15 13 10 0 0 9 2 16 9 13 1 10 9 9 2 13 15 2
2 9 5
25 9 13 1 0 0 9 7 9 15 13 9 2 13 9 1 9 7 3 13 15 1 9 1 9 2
13 9 1 11 9 2 11 11 2 13 10 1 15 2
15 15 4 0 9 13 15 1 10 2 0 9 2 1 11 2
23 2 15 13 0 9 1 9 1 11 7 0 11 9 15 13 0 0 0 9 2 13 11 2
21 11 13 1 10 0 9 16 15 3 13 3 3 0 9 1 9 1 10 0 9 2
20 11 13 15 4 13 1 16 0 9 7 9 1 9 13 1 9 1 0 9 2
19 2 9 13 1 7 13 3 9 2 7 4 13 0 7 13 2 13 11 2
29 9 1 11 11 2 11 11 11 2 11 11 7 11 11 11 11 4 13 1 14 13 0 9 1 9 2 1 9 2
18 10 9 13 1 9 11 11 1 16 12 9 1 9 1 11 13 9 2
17 10 10 11 13 9 16 15 13 11 1 2 11 2 1 0 9 2
33 15 13 1 9 9 1 11 11 15 13 0 1 11 11 2 7 15 13 9 1 9 1 10 9 1 9 1 11 11 1 11 11 2
16 2 16 0 9 13 1 9 7 9 13 15 1 14 13 9 2
13 9 4 13 1 1 9 7 15 13 10 0 9 2
19 7 16 15 15 13 1 13 0 2 13 3 3 15 15 13 1 10 0 2
9 15 4 3 13 0 2 13 11 2
8 2 9 13 10 9 1 11 2
29 15 4 15 13 7 1 9 1 9 7 0 9 1 11 2 15 1 9 4 13 0 7 13 1 9 2 13 11 2
12 9 1 9 2 9 7 9 13 10 9 9 2
10 2 9 13 10 0 9 1 10 9 2
19 15 13 3 10 10 0 9 1 10 9 2 7 0 9 13 0 7 0 2
14 15 13 10 10 9 11 13 15 13 1 2 13 11 2
4 9 1 11 5
11 9 1 11 4 13 1 0 9 1 11 2
16 11 13 0 9 1 9 9 2 7 15 13 3 11 1 1 2
3 13 9 2
15 11 13 1 10 0 9 1 9 1 11 9 7 11 9 2
7 3 11 11 1 9 9 2
24 10 0 1 11 13 9 1 9 4 13 10 9 16 15 4 13 9 1 9 1 9 1 9 2
5 7 9 13 0 2
21 5 11 1 9 4 13 1 12 12 9 1 12 1 1 12 2 12 9 1 12 2
19 16 15 1 12 3 13 11 11 15 13 9 2 13 0 9 3 1 9 2
15 9 1 10 9 4 13 1 12 12 1 12 12 12 9 2
13 5 10 0 9 11 4 13 2 1 9 1 9 2
20 5 11 4 13 1 9 10 9 16 3 12 9 1 9 1 9 13 1 9 2
15 5 11 4 13 9 1 9 11 11 2 11 11 7 11 2
16 5 11 1 0 9 2 9 7 9 4 13 1 12 9 9 2
11 9 1 9 4 13 1 3 12 9 9 2
16 5 0 4 9 1 0 9 7 9 13 1 1 12 9 9 2
12 5 11 13 1 9 0 1 9 7 0 9 2
13 5 9 4 13 1 9 9 1 11 9 7 9 2
22 5 0 9 1 9 7 10 9 4 13 2 7 9 1 9 1 9 1 9 4 13 2
14 5 11 2 10 0 9 1 9 7 9 13 1 12 2
26 9 1 9 2 9 7 9 2 11 11 2 11 2 2 13 10 0 4 13 9 1 9 1 10 9 2
3 4 13 5
20 2 15 13 14 13 0 1 7 13 10 0 9 15 4 13 1 12 1 3 2
35 0 13 3 1 13 15 15 4 13 1 2 7 16 11 13 1 9 7 13 0 9 2 4 15 13 10 9 1 9 1 11 2 13 15 2
34 1 9 1 9 13 11 14 13 9 9 1 9 1 12 9 2 7 0 13 10 0 9 1 9 1 11 13 1 11 7 10 10 9 2
12 11 1 10 9 2 13 14 13 1 10 9 2
13 2 9 13 3 3 0 1 15 7 10 10 9 2
43 15 13 14 13 10 9 1 9 1 9 7 9 2 7 3 13 15 1 0 9 14 13 9 1 9 2 9 7 0 2 7 9 2 13 11 9 1 11 2 11 11 11 2
24 7 15 13 0 1 16 9 13 10 10 9 1 10 0 9 16 15 13 9 1 9 1 9 2
22 2 1 11 13 15 0 9 1 16 9 7 9 4 13 0 1 1 9 2 13 11 2
2 9 5
10 2 10 9 13 1 0 9 1 9 2
17 15 13 15 13 0 9 1 9 16 15 13 15 1 9 1 9 2
20 11 13 3 15 13 0 16 9 1 9 7 9 1 9 13 9 1 9 9 2
39 2 15 13 3 0 0 16 16 9 1 9 1 10 0 9 4 13 1 9 1 9 1 9 2 13 15 0 1 14 13 9 1 11 11 2 9 7 11 2
20 15 13 9 4 13 9 1 14 13 10 9 1 1 10 0 9 2 13 9 2
27 11 1 9 2 15 13 16 1 12 9 1 9 1 9 4 13 1 9 2 13 11 13 0 1 10 9 2
3 10 9 5
28 16 9 9 13 16 10 11 1 9 4 13 9 2 13 11 9 11 11 0 1 16 15 3 13 1 14 13 2
10 15 13 9 2 3 9 2 1 9 2
24 2 1 11 7 11 1 10 9 3 1 11 13 3 11 10 9 1 14 13 9 1 9 10 2
31 15 13 3 9 4 13 0 3 2 7 15 13 9 1 16 9 1 11 4 13 14 13 1 9 1 10 0 2 13 9 2
19 11 13 9 1 11 7 10 10 9 3 13 10 12 0 0 9 1 11 2
38 2 9 1 9 0 7 0 9 13 10 0 9 1 15 7 11 2 13 11 2 7 13 11 1 14 13 1 14 13 3 0 0 7 0 9 1 9 2
4 0 0 9 5
23 11 11 2 11 2 13 0 9 1 9 13 1 1 14 13 16 9 13 16 15 13 0 2
31 2 9 1 14 13 10 0 0 9 1 9 13 14 13 16 10 0 0 9 15 9 2 9 7 9 13 1 9 13 0 2
33 15 13 15 1 9 0 14 13 1 16 9 7 9 13 10 0 9 2 7 16 9 13 1 3 0 9 1 0 9 2 13 11 2
11 2 9 1 0 9 13 1 1 0 9 2
14 15 13 0 13 0 9 1 10 0 9 2 13 15 2
3 0 9 5
3 9 9 5
27 5 1 11 4 15 13 15 1 10 0 9 1 10 0 9 9 1 9 1 10 9 2 3 3 1 9 2
26 11 13 1 10 0 9 2 0 1 9 2 16 0 9 13 0 1 9 2 7 4 13 11 1 0 2
31 1 11 11 1 11 11 13 9 16 11 13 9 1 11 1 14 13 9 2 15 3 4 13 1 11 1 14 13 1 11 2
16 9 9 11 11 11 4 3 13 16 9 4 13 0 1 11 2
10 11 13 1 10 9 1 11 11 11 2
7 2 13 1 15 10 9 2
30 11 2 1 10 9 7 10 9 15 13 0 1 11 2 13 3 3 1 9 1 14 13 1 10 0 9 0 1 11 2
9 5 10 10 9 13 11 1 11 2
33 11 4 13 1 12 0 9 1 10 0 0 9 2 15 13 16 15 3 4 4 13 3 1 0 9 2 16 15 13 10 9 9 2
23 2 1 9 1 11 9 7 9 2 13 15 10 0 9 13 1 11 2 2 13 11 0 2
25 9 9 4 3 13 9 2 7 1 10 9 1 11 3 13 15 1 0 9 1 9 1 0 9 2
17 2 13 15 2 4 9 13 9 1 11 2 7 9 13 0 9 2
15 9 1 11 7 11 4 13 1 11 9 2 2 13 15 2
23 5 9 0 9 13 16 10 0 9 13 3 1 14 13 15 0 9 1 14 13 0 9 2
12 10 0 9 4 13 15 1 0 9 7 9 2
13 0 4 15 13 3 1 14 13 1 7 13 9 2
17 9 4 13 15 1 16 15 10 3 13 15 15 13 1 10 9 2
11 10 9 4 13 10 0 0 9 1 9 2
41 1 9 1 0 9 2 4 15 13 10 0 9 2 15 7 4 13 11 7 10 0 9 2 7 15 1 9 13 9 1 14 13 9 1 11 1 10 9 1 9 2
3 0 9 5
3 9 9 5
21 10 0 0 9 1 0 9 7 9 13 1 9 1 14 13 10 0 9 1 9 2
48 9 1 9 13 0 2 10 0 9 7 9 13 0 2 7 0 13 15 1 0 9 15 3 4 13 10 9 1 9 15 4 13 1 9 1 9 2 9 7 9 2 1 9 1 9 7 9 2
18 10 0 9 4 13 1 1 12 9 9 3 16 10 0 13 1 12 2
11 7 15 13 1 16 10 0 9 4 13 2
36 11 11 9 11 11 13 10 9 3 10 9 15 13 1 1 0 9 2 4 13 1 10 9 0 9 7 9 2 1 9 1 9 7 9 10 2
17 1 12 13 0 9 9 1 3 10 9 1 10 0 9 1 11 2
12 1 12 4 15 13 9 3 1 10 0 9 2
17 7 16 10 0 9 4 13 10 9 2 4 3 9 13 1 9 2
23 3 4 15 7 13 9 0 7 0 2 13 1 9 1 9 7 13 1 16 11 13 9 2
9 10 10 9 4 13 0 0 9 2
22 10 9 1 0 9 4 13 13 16 9 1 0 9 1 10 0 9 13 0 7 0 2
39 12 9 1 9 13 0 7 3 0 1 9 1 16 0 9 13 1 0 9 1 9 2 16 1 12 9 13 0 1 16 9 13 3 0 1 1 9 9 2
28 9 1 11 2 11 2 11 2 11 7 11 13 0 1 9 2 16 9 1 11 7 11 1 0 9 13 9 2
19 11 4 1 10 9 13 14 13 10 9 15 13 0 0 1 10 0 9 2
21 11 13 10 0 9 1 10 9 2 7 3 4 9 13 1 3 1 11 7 11 2
22 9 13 15 14 13 1 14 13 9 1 9 7 1 9 13 10 9 1 11 7 11 2
4 13 0 9 5
2 9 2
15 1 0 9 13 11 3 10 0 10 9 15 15 0 13 2
11 11 11 13 14 13 9 1 10 0 9 2
2 13 2
21 11 11 13 9 1 11 4 13 1 16 15 13 1 12 1 12 9 9 1 9 2
2 9 2
4 11 11 11 5
23 2 16 15 1 0 9 13 1 0 9 2 13 15 16 9 13 10 0 9 1 10 9 2
21 3 4 15 3 13 10 9 7 9 15 13 1 10 0 9 2 13 9 11 11 2
26 9 13 11 9 16 10 0 1 9 13 9 1 0 9 16 15 4 13 1 0 9 10 0 12 9 2
23 3 4 9 1 0 1 9 7 9 1 9 13 15 1 9 1 0 9 1 9 15 13 2
34 9 4 3 13 9 11 11 9 2 15 13 16 9 4 13 9 1 14 13 10 9 15 13 0 15 0 13 0 9 9 1 0 9 2
15 2 15 13 3 0 14 13 1 9 15 4 13 1 11 2
53 15 13 10 9 15 13 0 1 14 13 1 9 1 14 13 9 1 0 9 2 7 15 4 13 15 0 1 10 9 1 14 13 1 9 9 1 15 1 0 9 15 1 3 9 3 4 13 0 9 2 13 15 2
19 9 13 1 9 1 10 9 9 15 15 13 0 4 13 9 1 0 9 2
23 2 15 13 10 9 1 0 9 15 13 0 2 0 9 2 1 13 10 0 9 1 9 2
14 15 13 10 0 9 2 15 15 0 4 13 1 9 2
17 3 13 15 16 15 13 14 13 1 9 10 0 9 2 13 11 2
4 13 3 15 5
30 1 11 9 13 0 1 9 1 12 9 1 9 12 9 2 16 0 1 9 1 12 7 12 9 1 9 13 12 9 2
22 2 15 13 1 14 13 9 1 9 1 0 1 9 2 13 9 1 9 11 11 11 2
37 11 2 15 3 13 9 1 11 1 11 2 13 9 1 9 15 9 4 13 1 11 2 11 2 11 2 11 2 11 2 11 2 11 7 11 9 2
25 2 3 0 9 15 13 1 9 13 0 1 16 15 13 9 7 16 15 4 13 1 9 1 9 2
26 0 13 9 1 0 1 0 0 9 0 2 16 15 1 9 3 4 13 9 1 14 13 2 13 11 2
11 15 13 16 9 3 3 13 15 1 3 2
25 2 1 9 13 15 3 15 2 7 10 9 13 3 3 9 1 9 15 15 3 13 1 1 9 2
24 7 15 13 0 16 15 4 13 9 1 9 1 9 2 15 4 13 9 1 9 7 9 0 2
22 15 13 3 0 1 10 0 2 15 3 13 0 0 9 14 13 15 1 2 13 15 2
5 9 13 1 9 5
24 9 1 9 1 0 9 1 9 15 1 9 13 1 0 9 13 10 1 9 9 1 10 9 2
12 3 12 10 1 11 9 4 13 1 9 9 2
25 12 9 1 9 9 7 9 1 16 12 9 1 10 9 15 13 1 0 9 4 13 0 1 9 2
21 3 13 9 11 14 4 0 1 10 0 9 1 10 9 13 3 16 9 4 13 2
10 2 6 2 3 4 15 3 13 9 2
11 15 13 3 11 1 10 0 2 13 15 2
4 2 1 9 2
23 11 11 2 9 1 11 9 1 11 2 13 1 14 13 9 10 0 1 9 1 11 9 2
32 15 13 0 1 10 12 9 9 2 7 13 1 14 13 1 1 1 12 9 16 15 3 13 9 1 10 9 15 0 13 1 2
47 2 15 13 3 3 9 1 14 13 9 1 0 9 2 7 15 13 0 15 13 10 9 0 2 13 11 2 15 13 15 13 10 0 9 15 13 0 1 15 14 13 1 10 3 0 9 2
19 2 15 13 1 14 3 13 16 15 13 3 9 1 14 13 9 10 9 2
27 1 10 12 9 9 13 15 12 9 13 1 9 2 15 4 3 13 15 10 3 0 15 13 2 13 9 2
19 15 13 0 1 9 1 9 2 7 4 13 1 11 9 12 9 1 15 2
18 11 13 3 15 13 9 7 9 1 9 16 3 0 13 9 1 9 2
20 2 15 15 13 1 0 9 13 0 9 1 9 1 15 15 3 13 0 9 2
14 3 13 15 0 0 0 9 14 13 15 1 1 9 2
32 0 1 15 13 0 2 7 15 13 0 16 10 9 13 1 0 0 9 3 2 3 16 9 4 13 15 3 0 3 15 1 2
11 7 11 13 9 3 13 10 9 3 0 2
17 2 15 13 10 0 9 1 14 13 9 13 0 1 3 0 9 2
7 7 15 13 3 1 9 2
13 3 15 1 10 4 13 9 1 12 9 9 3 2
8 2 13 15 3 13 1 9 5
28 2 15 11 4 13 1 1 10 9 13 10 9 15 4 13 1 9 1 9 2 13 9 11 11 11 1 11 2
22 15 13 0 1 16 9 1 11 9 4 13 1 11 2 1 3 0 9 1 10 9 2
13 2 11 13 3 10 9 15 13 15 13 1 9 2
26 15 13 0 1 14 13 10 0 9 1 9 2 7 15 13 0 1 15 14 13 10 9 2 13 11 2
18 15 13 15 13 3 0 14 13 9 1 9 9 1 1 9 1 12 2
31 2 3 13 15 1 1 10 9 2 7 14 13 3 13 7 15 15 13 9 7 15 15 13 0 1 14 13 2 13 9 2
29 15 4 1 10 9 3 13 15 1 11 9 1 16 11 4 13 1 1 14 13 1 1 9 7 9 1 0 9 2
10 2 15 13 10 0 9 1 10 9 2
25 1 15 13 15 0 14 13 10 0 9 1 10 0 9 2 7 15 13 3 3 0 1 0 9 2
16 7 15 13 0 14 13 0 1 1 10 9 3 2 13 11 2
4 10 0 11 5
7 11 13 0 1 0 9 2
11 9 13 3 10 0 9 1 9 7 9 2
2 9 2
20 11 0 9 1 9 13 3 10 9 1 10 0 9 1 11 2 13 11 11 2
17 2 15 4 13 10 0 11 0 9 2 13 9 7 9 11 11 2
20 1 10 0 9 1 10 0 9 13 15 10 0 0 9 15 13 11 1 9 2
13 1 10 9 13 1 10 10 0 9 11 0 9 2
20 15 13 1 9 7 9 1 9 11 11 2 15 13 10 9 1 10 0 9 2
4 10 10 11 5
21 2 15 4 0 4 13 10 9 3 15 13 10 0 9 1 2 10 0 9 2 2
20 7 15 13 10 9 1 14 13 1 10 1 10 0 9 15 13 9 1 9 2
14 7 3 4 15 13 1 10 0 9 1 11 0 9 2
11 7 9 13 10 0 0 9 1 10 9 2
10 9 13 7 10 9 7 10 0 9 2
23 11 13 16 15 13 0 14 13 10 9 1 14 13 10 0 1 9 15 13 3 0 1 2
13 2 1 0 13 11 0 1 11 2 11 7 11 2
19 7 11 13 0 1 10 0 7 0 9 1 0 0 9 7 10 0 9 2
11 15 13 14 13 1 10 9 1 10 9 2
9 2 15 4 13 10 3 0 9 2
9 2 6 2 15 13 3 3 0 2
17 7 4 15 13 1 11 9 2 4 15 3 13 1 10 0 9 2
11 10 0 11 13 10 3 0 7 0 9 2
14 7 10 0 9 1 9 13 3 0 1 10 0 9 2
8 2 15 13 10 9 1 9 2
11 0 0 9 1 10 9 4 13 0 1 2
9 7 0 13 16 9 4 4 13 2
9 7 16 10 0 9 4 4 13 2
21 15 13 0 9 15 4 13 10 9 15 15 13 1 11 1 9 9 2 13 11 2
17 11 13 0 16 15 3 4 4 13 10 0 9 1 10 0 9 2
14 2 10 1 10 0 0 9 13 3 1 9 1 11 2
14 10 9 2 0 9 1 0 9 2 13 15 13 0 2
19 0 9 13 15 4 13 1 1 11 1 14 13 10 0 9 13 9 10 2
29 15 13 3 9 1 10 0 9 15 13 0 14 13 1 2 7 15 4 3 3 1 0 9 4 13 1 10 9 2
10 15 4 3 3 13 9 1 0 9 2
13 1 0 10 0 9 2 13 15 0 14 13 0 2
4 9 13 1 5
22 11 13 3 1 9 1 9 1 10 1 10 9 3 10 0 9 3 13 10 0 9 2
12 15 4 13 0 9 15 13 1 10 0 9 2
18 1 10 0 0 9 13 10 9 15 13 9 1 9 1 9 11 11 2
25 7 11 4 3 13 9 1 10 9 13 2 11 9 2 2 15 15 3 13 15 15 13 0 0 2
13 10 9 13 10 9 1 9 1 11 11 1 11 2
20 2 11 9 2 7 10 0 0 2 11 11 2 13 10 9 1 9 7 0 2
15 2 15 13 1 9 2 11 9 7 13 1 9 1 9 2
13 1 9 13 15 9 1 14 4 13 0 0 9 2
16 9 15 13 13 0 0 15 15 13 1 1 0 1 10 9 2
11 3 0 9 1 16 11 13 1 10 9 2
12 10 0 9 4 13 1 0 9 2 13 11 2
28 1 14 13 3 2 11 9 2 13 10 0 9 2 13 11 1 10 12 0 9 1 11 2 3 11 7 11 2
15 2 1 13 15 3 16 11 13 1 9 1 10 0 9 2
7 9 1 9 13 1 11 2
11 3 4 10 0 9 13 1 2 13 15 2
15 11 13 0 1 3 9 1 9 4 13 0 7 0 0 2
21 2 3 13 15 0 14 13 1 0 9 7 0 9 1 9 2 3 10 0 9 2
19 15 13 3 16 9 1 2 11 9 2 13 1 1 14 13 10 10 9 2
9 15 13 7 13 10 0 0 9 2
3 0 9 5
8 2 11 13 1 0 1 11 2
10 3 13 9 1 9 1 9 7 9 2
14 2 11 13 9 9 2 7 15 13 0 9 1 9 2
7 9 13 16 11 13 9 2
14 0 13 15 10 0 9 1 9 9 1 11 7 11 2
7 10 0 9 13 0 9 2
13 7 15 13 10 0 9 1 9 7 1 10 9 2
31 2 15 13 3 3 10 0 9 1 0 0 9 16 15 13 10 0 9 1 9 9 1 11 2 7 15 13 9 1 11 2
19 2 10 0 9 13 0 0 1 14 13 9 1 10 0 0 9 1 11 2
11 15 13 3 10 0 0 9 15 9 13 2
15 15 13 3 0 16 0 9 13 14 13 10 9 1 11 2
15 15 13 9 11 0 9 13 1 10 0 9 2 13 11 2
10 2 11 13 3 3 10 9 1 9 2
13 2 11 4 0 13 1 9 1 9 1 0 9 2
16 15 15 4 13 9 11 10 2 4 3 13 0 1 10 9 2
21 1 9 4 15 13 16 15 13 10 9 1 11 7 10 0 9 15 13 0 9 2
12 11 13 16 9 1 10 9 13 0 1 9 2
26 2 11 4 3 13 10 0 9 1 14 13 9 1 0 1 15 15 4 13 1 0 9 2 13 15 2
3 0 9 5
12 10 0 9 1 11 13 1 0 1 3 0 2
18 9 1 11 11 7 11 11 4 13 9 1 0 9 1 0 7 0 2
18 2 11 4 13 9 15 3 4 13 0 0 1 9 1 10 0 9 2
17 15 4 13 15 9 2 7 10 0 9 1 0 9 2 13 11 2
12 11 13 10 1 10 0 0 9 1 11 9 2
27 15 13 1 0 1 2 9 11 2 7 4 1 9 4 13 1 0 1 10 9 1 9 1 10 0 9 2
14 11 4 3 13 12 9 7 13 3 1 11 0 9 2
18 15 4 3 13 10 9 1 15 11 13 1 10 0 0 9 1 11 2
25 2 15 13 3 10 9 1 3 10 9 1 0 9 1 10 0 2 10 0 7 10 0 13 15 2
11 7 3 10 9 13 3 0 2 13 11 2
4 2 13 9 5
3 9 0 2
10 10 0 11 13 15 0 9 1 11 2
10 9 13 14 13 10 0 9 1 9 2
2 13 2
20 11 7 9 11 11 2 9 2 4 3 4 13 9 1 9 2 13 11 11 2
14 2 10 0 9 13 14 13 11 7 11 11 1 9 2
27 15 4 13 15 0 1 16 15 3 3 13 10 0 9 2 7 10 0 0 9 2 13 11 11 1 11 2
12 15 13 0 9 1 10 0 9 11 1 11 2
19 13 1 10 0 9 13 9 3 1 14 13 0 9 1 10 0 0 9 2
15 9 13 3 9 1 0 9 1 9 15 4 13 0 9 2
31 10 0 9 2 15 13 1 11 2 11 2 2 11 11 2 11 2 2 11 11 7 11 13 1 3 12 9 1 0 9 2
14 10 0 9 15 13 1 9 2 13 1 3 12 9 2
24 11 2 15 13 10 9 1 11 2 11 11 11 7 11 11 2 13 0 9 1 10 0 9 2
9 15 13 1 12 9 1 12 9 2
9 15 13 12 9 1 10 0 9 2
19 9 15 3 4 13 0 1 16 9 4 13 10 0 9 1 14 13 9 2
13 13 9 9 4 11 13 1 9 1 11 7 11 2
27 2 15 13 9 1 9 7 15 4 13 15 0 16 3 0 15 13 3 0 9 4 15 13 2 13 11 2
6 11 7 11 1 9 5
28 10 9 4 13 10 0 9 1 0 9 2 15 4 4 13 12 9 1 9 1 16 10 0 13 9 1 12 2
19 9 11 11 11 13 9 9 2 3 10 0 9 11 13 3 1 11 11 2
20 10 0 11 11 7 9 11 11 13 3 1 10 0 9 15 13 9 1 11 2
23 1 12 1 10 0 12 9 4 10 9 15 13 1 9 0 1 9 2 13 1 1 9 2
14 11 11 11 13 9 9 7 13 1 10 9 0 3 2
12 11 11 11 4 3 3 13 10 9 1 9 2
10 7 3 2 7 16 9 4 13 9 2
8 10 0 9 4 3 4 13 2
18 2 3 4 15 13 16 11 7 11 4 13 0 1 9 10 0 9 2
9 15 4 1 10 13 9 1 9 2
8 15 13 16 9 4 13 1 2
24 15 4 13 1 16 3 0 13 9 7 1 16 0 13 1 14 13 1 1 9 2 13 15 2
21 11 13 16 11 3 1 9 4 13 15 1 9 2 11 11 0 9 2 11 11 2
21 2 11 4 3 13 11 11 2 1 9 1 14 13 10 9 1 9 2 13 15 2
5 2 11 1 9 5
27 3 16 11 4 13 1 1 9 1 10 0 9 2 4 15 3 13 1 9 14 13 13 1 11 7 11 2
16 10 12 9 13 10 9 1 3 12 7 12 9 1 0 9 2
13 2 13 15 14 4 13 1 9 1 10 0 9 2
8 2 6 2 15 13 15 3 2
12 7 9 13 14 13 11 7 11 1 10 9 2
9 4 15 13 1 15 13 15 9 2
19 11 7 11 13 9 1 14 13 1 10 0 16 15 13 15 2 13 11 2
17 1 11 0 9 13 9 1 10 0 0 9 11 13 3 1 1 2
17 11 11 9 4 13 10 9 1 10 0 9 1 12 9 0 9 2
28 2 15 13 10 9 15 13 0 0 3 3 2 7 15 13 14 13 11 1 1 10 0 9 15 13 15 1 2
65 9 11 13 1 9 14 13 9 1 10 9 9 2 7 15 4 13 1 10 12 0 7 1 10 9 1 0 15 13 9 2 7 13 16 9 3 13 0 1 0 2 13 11 2 15 4 13 1 16 15 15 4 13 9 1 12 9 1 9 4 13 0 1 9 2
3 9 0 5
11 9 4 1 0 9 4 13 0 0 9 2
13 7 1 0 9 13 9 3 0 0 1 0 9 2
16 2 15 13 15 1 9 16 9 13 0 0 1 9 1 9 2
6 2 15 13 0 0 2
11 10 0 9 4 13 1 9 1 12 9 2
18 11 4 4 13 1 10 9 2 7 13 9 1 9 1 9 7 9 2
9 3 4 10 9 13 2 13 11 2
17 15 13 11 0 9 13 1 9 1 14 13 1 1 10 0 9 2
10 2 9 4 13 7 9 4 13 3 2
11 15 13 1 10 9 3 1 12 13 9 2
14 15 13 0 0 1 16 12 13 1 9 2 13 15 2
22 9 13 10 9 16 10 0 9 1 0 9 13 0 1 9 1 10 0 9 7 9 2
9 0 11 11 7 11 11 4 13 2
19 10 10 9 4 15 13 1 1 16 9 11 11 1 10 0 13 9 1 2
28 10 9 13 15 16 9 10 1 9 1 9 13 0 14 13 9 1 1 11 11 7 1 14 13 9 1 9 2
10 11 11 1 10 9 13 1 10 9 2
27 9 13 15 1 10 9 1 14 13 9 1 9 3 9 13 1 2 1 11 2 11 2 11 7 11 9 2
18 15 13 10 0 9 11 13 11 4 13 10 9 1 16 9 13 9 2
30 2 15 4 13 12 9 1 0 9 3 9 4 13 9 1 11 11 1 9 10 9 15 4 13 1 9 2 13 15 2
15 3 4 3 10 0 9 11 11 13 10 9 1 0 9 2
24 2 9 13 10 0 9 1 11 15 4 13 1 9 1 10 0 0 9 1 3 2 13 11 2
2 0 5
30 9 11 11 11 4 13 10 0 9 9 1 10 0 9 9 13 0 1 7 13 3 9 1 14 13 1 11 0 9 2
7 2 9 4 13 1 9 2
20 15 4 13 15 0 1 15 15 4 13 2 13 9 1 9 1 9 10 9 2
4 9 13 15 5
17 13 1 14 13 10 9 1 9 2 13 15 3 0 9 1 11 2
3 1 9 2
19 15 13 1 9 11 2 9 2 15 13 11 1 11 9 2 13 11 11 2
10 3 13 11 11 14 13 1 0 9 2
4 3 13 15 2
8 3 1 11 11 2 3 0 2
64 3 2 13 16 16 11 13 2 7 11 9 13 14 13 9 1 0 9 1 12 2 4 15 13 2 1 10 0 9 11 11 2 1 9 2 1 9 7 10 0 9 2 9 2 2 16 9 13 2 9 2 7 2 9 2 15 3 4 13 16 9 13 1 2
53 16 11 7 10 9 1 10 9 13 15 1 9 2 7 16 9 13 2 3 0 9 4 15 13 16 15 3 4 13 1 2 9 2 2 15 3 3 13 16 9 1 11 13 15 15 13 3 7 16 9 13 0 2
3 13 15 2
30 15 4 3 13 12 9 16 15 13 9 1 2 16 10 9 1 11 11 4 13 2 9 2 7 13 15 1 11 9 2
4 13 15 9 2
20 0 13 15 1 10 0 1 10 0 1 10 9 2 1 10 9 1 11 9 2
20 15 4 3 13 10 0 9 2 7 0 13 9 10 0 9 1 10 10 9 2
10 15 4 3 13 10 9 1 1 11 2
19 10 9 2 10 0 2 0 9 2 16 0 9 4 13 9 1 1 9 2
15 1 9 1 0 2 0 7 0 11 13 15 10 0 9 2
9 2 3 13 15 1 1 9 2 2
10 15 13 15 1 15 14 13 2 3 2
36 7 9 1 0 9 2 9 2 0 0 0 9 7 0 0 7 0 9 2 15 3 13 2 9 2 7 3 9 2 13 3 15 11 0 9 2
32 3 4 15 3 13 9 1 15 3 2 7 1 9 13 15 15 15 13 11 2 1 0 0 9 7 9 15 4 13 9 0 2
47 15 4 13 1 1 0 9 1 10 10 9 2 0 3 15 13 1 11 11 11 0 2 3 16 15 3 13 10 9 16 15 4 13 1 11 2 7 15 4 3 13 16 9 1 11 13 2
11 0 13 9 1 11 15 1 10 0 9 2
38 16 11 4 13 2 13 9 9 1 9 1 0 9 0 2 16 15 15 4 13 15 1 14 13 1 9 1 16 11 4 13 11 2 4 13 15 0 2
21 16 11 7 9 11 4 13 2 4 15 0 13 1 16 9 1 9 13 1 9 2
29 15 11 0 4 13 2 7 15 4 13 15 0 2 13 9 1 16 11 4 13 15 0 1 10 0 9 1 11 2
16 7 3 4 9 0 13 15 0 1 9 1 10 0 0 9 2
24 11 13 9 3 11 1 0 9 1 9 1 12 1 0 9 13 0 9 10 9 1 9 9 2
16 15 13 0 12 9 1 10 9 2 7 13 3 10 0 11 2
30 15 13 9 1 10 0 0 9 1 11 0 9 2 11 2 2 7 7 9 7 9 1 4 13 0 1 11 0 9 2
24 10 0 9 11 13 1 3 12 9 9 3 16 9 0 1 1 11 13 1 9 1 9 11 2
7 10 9 11 4 4 13 2
20 1 10 9 4 11 13 10 9 9 1 15 15 1 9 9 13 11 12 9 2
4 11 7 11 2
16 3 1 11 13 2 9 2 9 1 2 9 2 0 1 9 2
12 0 13 15 0 1 14 13 1 10 12 9 2
31 15 15 13 10 0 9 2 4 4 13 9 2 16 9 1 10 9 13 2 9 2 15 4 13 14 13 10 0 0 9 2
24 1 4 11 2 10 9 3 4 13 1 9 1 11 9 2 0 13 10 1 11 0 0 9 2
6 15 13 3 11 9 2
21 0 2 13 15 15 3 2 7 1 1 9 4 15 3 13 3 0 9 1 15 2
44 0 2 0 2 0 2 0 2 0 2 0 2 0 2 0 2 3 11 0 9 11 11 13 15 2 2 0 2 0 2 0 2 0 7 2 3 3 2 0 2 0 2 0 2
48 1 1 10 0 7 0 9 1 10 0 9 4 11 13 15 0 1 14 13 14 13 2 13 9 1 9 7 9 2 13 11 0 0 0 1 1 10 9 2 7 3 3 13 2 9 2 9 2
18 9 1 11 13 1 3 0 16 9 3 13 0 9 15 4 13 1 2
11 3 13 11 15 1 10 9 1 11 11 2
11 3 13 15 1 1 10 1 11 11 9 2
5 15 13 1 15 2
12 1 10 9 3 0 15 13 14 13 10 9 2
3 11 13 5
3 9 9 5
31 9 7 9 1 0 9 2 13 11 2 4 10 9 13 0 1 11 0 9 1 9 2 7 9 9 13 1 9 1 9 2
14 9 1 14 4 13 1 9 1 10 0 9 13 0 2
16 7 15 15 13 1 11 2 4 1 3 0 9 13 1 11 2
47 3 13 11 10 9 1 12 9 1 11 1 9 2 1 12 9 1 10 9 2 7 12 9 0 1 9 1 12 2 7 0 13 10 10 9 2 3 0 0 2 13 0 0 9 1 11 2
26 10 9 11 13 10 9 13 16 11 13 3 1 13 10 0 9 1 1 12 1 0 13 10 9 9 2
18 11 13 1 9 1 14 13 0 1 1 9 0 9 2 11 7 11 2
27 10 9 1 9 1 11 7 11 11 13 10 9 1 12 9 1 10 9 2 1 12 1 12 9 9 2 2
20 1 11 3 0 9 2 11 2 13 9 1 12 9 2 1 12 1 12 9 2
13 1 10 0 9 1 11 7 11 13 15 3 9 2
20 1 10 9 1 11 11 2 13 11 1 1 11 1 12 9 2 1 12 9 2
34 16 9 1 9 13 3 12 9 9 1 9 10 0 9 1 9 1 12 2 13 10 9 1 9 1 10 9 10 9 1 1 12 9 2
16 2 13 11 1 1 12 9 1 10 9 2 4 9 0 13 2
16 0 4 11 13 15 1 14 13 0 9 1 10 9 7 9 2
18 10 0 1 11 3 13 14 13 9 2 2 13 9 11 11 1 11 2
27 1 10 0 9 1 9 11 8 11 2 13 1 12 9 2 13 11 1 9 1 14 13 1 1 12 9 2
27 9 9 4 1 9 1 0 10 3 13 15 10 9 1 16 10 0 9 13 9 1 9 3 1 9 11 2
21 16 10 0 9 13 16 7 11 7 11 13 0 2 4 3 9 1 9 4 13 2
4 9 1 9 2
25 11 11 11 13 3 9 1 10 0 11 2 7 13 15 13 1 9 16 9 9 3 13 1 9 2
2 0 2
7 0 4 15 13 9 10 2
12 15 4 3 13 10 0 9 2 13 11 11 2
16 2 15 13 3 1 9 16 9 9 10 4 13 1 9 3 2
31 3 13 15 9 7 15 13 0 0 14 13 11 0 1 9 15 13 13 1 9 2 13 11 9 7 0 9 11 11 11 2
47 3 13 9 1 9 1 9 11 11 15 1 9 11 13 16 9 13 10 9 16 15 3 13 0 2 7 13 1 10 9 1 10 0 9 9 1 0 7 0 9 1 9 7 1 0 9 2
4 11 13 15 5
17 7 15 13 3 10 12 1 9 1 11 15 11 4 13 15 1 2
43 7 3 11 13 16 11 9 1 12 4 13 0 9 1 0 9 7 13 9 1 10 9 15 3 4 13 9 1 7 16 15 3 13 10 0 9 2 13 11 0 0 9 2
26 2 15 13 0 0 1 9 11 11 7 11 11 15 1 11 13 16 9 1 12 13 15 2 13 11 2
21 2 3 13 15 0 2 15 11 13 2 16 9 13 1 1 10 0 9 1 9 2
22 9 13 1 9 1 10 0 9 1 9 1 11 2 15 9 2 11 2 4 13 1 2
4 0 1 11 5
22 11 13 3 0 1 11 1 16 9 9 4 13 0 9 1 9 2 9 7 1 9 2
27 2 13 16 9 3 13 9 1 10 9 1 9 2 7 1 14 13 9 7 14 13 1 9 10 2 9 2
27 3 1 13 0 3 0 16 15 13 1 12 2 13 11 2 15 7 4 13 9 2 9 7 9 1 9 2
25 2 7 11 13 11 9 11 11 1 10 0 9 1 12 2 13 3 15 16 9 9 4 13 9 2
20 2 10 9 13 0 9 2 7 15 13 0 16 11 13 10 9 1 10 9 2
33 7 1 11 9 4 10 9 3 4 13 1 0 9 7 9 2 7 3 0 15 4 13 4 10 0 13 2 13 11 2 7 13 2
28 2 15 13 0 14 13 16 11 13 16 0 9 1 9 1 0 9 13 1 9 7 16 9 4 13 0 9 2
9 7 9 4 3 13 1 10 9 2
3 3 1 2
9 10 0 9 4 13 9 7 9 2
8 3 13 15 1 9 1 11 2
4 13 0 9 5
23 2 7 11 13 16 9 3 3 13 3 0 7 3 0 1 14 13 0 9 15 11 13 2
9 2 10 0 9 1 9 13 0 2
28 16 15 15 13 15 1 9 13 1 0 9 2 13 15 0 1 9 7 3 1 14 13 9 1 9 7 9 2
22 15 4 15 13 1 7 13 9 2 15 0 0 9 4 13 1 9 1 1 0 9 2
25 2 0 4 15 13 16 9 3 13 10 10 1 9 2 15 15 4 13 9 1 1 9 1 9 2
26 15 4 13 10 0 9 16 15 13 15 2 13 11 2 15 3 13 9 1 9 7 9 1 0 9 2
14 15 13 15 3 0 0 1 11 9 1 10 0 11 2
14 2 7 15 13 3 10 9 1 10 0 9 1 9 2
14 1 10 9 13 3 11 15 15 15 13 2 13 11 2
4 13 9 10 5
8 2 0 4 15 13 9 10 2
27 15 4 3 13 10 0 9 7 4 3 13 1 10 0 2 13 11 11 2 9 7 9 1 9 11 11 2
16 2 7 15 1 9 1 9 11 15 4 13 1 9 1 9 2
22 2 15 4 3 13 16 9 13 1 1 14 13 16 10 9 1 9 13 1 10 0 2
23 15 15 4 13 1 15 2 4 1 3 9 13 15 1 16 9 4 2 13 2 10 9 2
6 15 4 15 13 3 2
12 11 13 3 16 15 13 0 9 1 11 9 2
16 2 15 13 15 15 13 16 9 13 10 9 14 13 9 1 2
33 3 4 15 1 9 13 9 15 13 0 16 15 1 9 1 9 13 10 9 1 16 9 13 9 14 13 10 0 9 2 13 11 2
16 15 13 0 16 9 4 13 0 10 9 1 15 11 13 1 2
16 2 16 9 13 9 10 2 4 15 13 1 9 2 3 9 2
7 15 13 10 9 1 9 2
16 15 13 9 15 4 13 2 1 9 13 15 16 9 13 0 2
20 9 4 3 13 15 15 13 1 14 13 1 9 1 16 15 3 13 0 9 2
19 15 13 1 9 7 1 10 9 4 9 13 1 1 14 13 1 10 9 2
24 2 11 13 3 3 3 16 9 7 9 13 9 3 2 7 16 15 3 7 0 13 10 9 2
6 15 13 15 1 15 2
20 2 10 12 15 13 13 16 15 3 13 9 1 9 1 14 13 1 10 9 2
23 7 15 13 0 1 16 9 4 13 2 7 15 13 3 16 15 4 13 9 10 9 0 2
18 15 4 13 9 1 11 2 7 0 3 13 9 1 9 2 13 11 2
17 2 7 3 13 15 1 10 1 9 13 1 10 9 9 15 13 2
29 13 15 10 0 9 15 13 1 9 1 14 13 9 7 13 15 10 9 15 13 3 1 10 9 1 10 0 9 2
19 13 15 10 0 9 2 13 15 0 0 1 16 15 13 0 1 1 9 2
17 10 9 4 15 3 13 1 12 7 15 4 15 4 13 1 1 2
8 2 13 15 9 1 10 10 5
30 11 11 2 9 1 11 2 9 1 11 7 11 2 2 13 16 9 1 0 9 7 9 1 0 9 1 9 13 0 2
33 2 15 13 0 16 9 13 0 2 7 9 16 9 0 13 15 13 1 14 13 1 1 9 2 13 3 1 10 9 2 13 15 2
24 2 15 13 15 1 10 9 9 11 11 13 1 9 15 13 1 0 9 7 13 9 10 0 2
10 2 15 13 3 3 15 13 15 1 2
15 10 9 15 13 15 13 0 13 15 9 3 1 10 10 2
18 11 13 3 16 10 9 1 9 9 7 10 9 1 10 9 13 0 2
34 2 11 7 11 4 3 13 1 14 13 9 9 1 14 13 9 1 11 11 2 15 3 3 4 4 13 10 0 12 9 2 13 15 2
26 2 11 11 4 3 13 14 3 13 9 1 10 9 7 3 13 15 1 10 9 3 0 1 9 9 2
31 11 13 16 15 13 11 9 14 13 7 13 9 15 13 1 16 0 9 13 0 1 9 1 9 1 1 10 9 1 9 2
17 2 1 9 13 0 1 9 1 11 11 1 9 2 9 7 9 2
40 15 13 0 16 15 13 1 0 9 2 7 3 9 13 1 9 13 15 3 10 0 9 1 15 15 0 13 0 1 9 7 15 15 13 1 9 2 13 15 2
15 2 7 1 14 13 1 15 10 9 3 13 14 13 1 2
15 4 9 1 9 7 9 0 1 9 0 13 11 9 9 2
29 11 13 16 9 15 4 13 1 9 7 9 1 0 9 4 13 2 7 10 9 1 10 9 13 1 9 1 9 2
13 9 4 13 14 13 10 0 9 1 9 7 9 2
18 2 9 13 3 9 7 9 7 9 7 9 2 7 13 10 0 9 2
15 15 13 15 1 9 1 16 15 13 0 9 16 9 13 2
5 13 15 1 9 2
9 9 1 9 9 13 1 0 9 2
6 7 9 13 9 0 2
2 11 2
24 2 15 4 13 10 0 7 0 0 9 1 0 9 2 2 13 11 11 11 1 9 15 13 2
9 3 1 12 1 15 2 11 11 2
17 2 15 13 15 13 0 0 16 9 4 13 9 1 9 0 9 2
28 0 9 13 9 1 15 2 1 10 16 11 11 11 4 13 1 9 1 0 9 2 13 9 7 9 11 11 2
29 2 9 1 7 9 7 9 13 0 9 3 1 14 13 1 9 7 1 14 13 1 10 0 9 1 14 13 9 2
22 9 1 10 9 13 16 15 15 13 1 0 0 4 13 1 10 9 2 3 10 9 2
21 15 13 10 9 1 14 13 16 3 10 9 13 15 0 1 0 9 2 13 11 2
21 15 13 1 16 9 1 9 1 9 4 13 0 1 9 2 0 1 9 1 9 2
2 11 5
15 10 0 9 4 3 13 1 9 9 1 9 1 0 9 2
25 9 13 10 0 9 1 16 15 15 13 1 9 1 1 9 2 0 4 13 1 10 9 1 9 2
41 2 13 15 0 14 13 10 0 9 1 1 3 15 13 9 2 2 2 13 11 11 11 11 2 10 9 15 4 13 1 9 1 10 9 1 9 11 4 13 1 2
30 2 4 15 13 1 9 2 4 15 13 0 0 1 1 9 7 3 13 9 15 4 4 13 1 14 13 10 0 9 2
5 9 2 1 9 2
11 15 13 10 9 15 13 9 1 0 9 2
29 16 9 13 15 15 4 4 13 1 14 13 15 1 7 0 7 1 0 9 2 13 11 11 11 1 11 1 11 2
2 9 5
24 1 9 13 11 11 11 1 15 10 12 9 0 1 14 13 10 0 9 11 8 11 1 9 2
17 2 10 9 15 13 15 14 13 10 10 9 1 12 7 0 0 2
32 14 13 13 0 9 9 2 2 13 15 1 10 9 1 15 10 1 2 12 2 2 9 15 13 1 1 9 1 9 1 9 2
12 10 10 9 15 13 0 1 2 13 11 11 2
16 1 10 15 11 13 2 13 10 0 9 1 1 9 1 9 2
18 2 15 13 0 1 10 10 1 11 11 12 1 10 9 1 10 9 2
20 2 2 2 15 4 13 10 0 7 0 0 9 1 0 9 2 2 13 15 2
27 11 11 13 1 11 16 15 13 15 13 0 16 9 7 9 1 0 13 10 0 9 1 9 1 10 9 2
23 2 10 9 1 9 1 11 8 11 13 16 9 13 1 1 9 2 7 13 15 1 9 2
53 10 0 9 4 3 13 1 14 13 0 9 7 9 16 9 3 13 1 10 0 9 15 0 13 1 9 1 10 9 2 13 11 2 15 13 1 16 15 3 13 10 9 1 14 13 16 0 9 13 9 1 9 2
13 2 15 13 10 9 1 14 13 9 2 13 15 2
2 9 5
17 2 13 15 1 9 9 2 2 13 9 1 11 11 11 11 11 2
28 15 4 13 9 1 0 9 1 11 8 11 2 7 13 1 16 9 1 9 13 1 9 1 9 1 0 9 2
17 2 9 13 1 16 0 0 9 13 9 1 10 9 1 0 9 2
22 15 13 0 1 16 10 0 9 4 13 9 7 9 2 16 15 13 0 7 0 9 2
29 15 4 13 0 9 1 9 1 1 9 2 7 0 1 9 2 9 7 1 7 1 1 10 3 0 1 11 11 2
34 2 7 15 13 3 10 0 9 1 9 1 11 11 7 1 0 0 9 1 9 11 11 2 16 15 10 4 13 16 15 13 1 9 2
13 2 3 2 9 13 3 3 1 9 1 15 10 2
27 15 13 3 9 1 9 1 14 13 16 0 9 13 0 0 1 10 9 2 7 15 4 13 0 1 15 2
34 10 9 16 15 13 9 13 16 9 0 3 13 10 10 9 1 14 13 1 9 1 15 15 13 7 13 2 15 15 13 1 10 9 2
18 15 13 3 3 0 9 13 1 9 1 9 2 16 15 3 13 3 2
32 2 4 15 3 1 10 0 4 13 10 9 1 16 10 10 9 15 13 1 9 1 1 2 4 4 13 1 9 1 0 9 2
15 2 10 0 0 13 1 10 9 15 13 1 10 9 1 2
17 9 4 13 9 16 15 3 13 9 1 14 13 9 1 0 9 2
4 15 13 0 2
19 7 9 13 1 15 10 0 0 9 15 4 13 9 3 3 15 4 13 2
23 11 13 3 0 1 9 7 10 9 15 4 13 1 10 9 2 13 11 2 7 13 1 2
28 2 4 15 13 10 1 3 9 1 16 15 13 10 0 9 1 9 2 4 15 13 9 1 9 1 10 9 2
22 7 15 13 10 9 9 15 13 16 9 3 13 0 1 16 15 1 13 9 7 0 2
13 0 13 1 16 15 13 0 9 15 3 13 0 2
4 0 0 9 5
9 11 11 11 13 1 9 1 11 2
5 2 15 4 13 2
36 13 15 0 14 13 10 9 2 7 13 15 16 15 13 10 9 15 4 13 1 0 0 9 2 7 15 1 15 10 3 13 9 2 13 15 2
23 2 7 13 3 3 15 16 0 9 13 1 0 9 2 10 9 1 16 15 13 10 9 2
31 2 15 13 3 10 0 9 2 7 11 11 2 15 10 0 9 13 2 13 3 10 9 2 15 13 3 7 0 10 9 2
42 15 4 3 3 13 1 16 15 4 13 15 1 14 13 2 15 13 1 14 13 14 13 10 0 9 9 7 9 7 3 0 9 15 13 1 10 0 9 2 13 11 2
39 15 16 11 13 10 9 1 2 11 11 2 1 9 2 13 9 3 13 16 15 3 13 9 1 15 10 15 13 9 1 9 1 14 13 0 9 1 9 2
21 2 10 15 15 13 13 0 0 2 15 4 13 1 14 13 15 1 1 10 9 2
29 1 10 9 15 13 10 9 9 1 14 13 9 10 1 10 9 2 13 15 3 16 15 13 9 15 13 15 3 2
18 15 13 0 3 13 9 15 13 0 1 2 15 13 9 2 13 15 2
4 9 7 9 5
21 9 1 9 11 11 11 13 3 9 16 9 13 10 0 9 1 9 13 3 0 2
12 2 15 13 1 3 9 16 9 13 0 0 2
21 15 13 10 9 15 13 10 9 1 2 15 15 13 0 7 13 1 10 9 9 2
15 15 13 3 0 9 15 13 9 1 9 1 2 13 15 2
2 9 5
3 9 9 5
31 9 13 1 9 1 14 13 15 1 10 9 2 16 10 0 9 13 3 0 9 11 7 11 4 13 15 1 10 0 9 2
31 10 9 1 10 9 1 9 11 8 9 13 16 11 1 9 13 10 9 1 12 9 2 10 9 1 12 9 1 10 9 2
11 11 13 12 9 2 10 9 1 12 9 2
30 1 11 11 13 9 11 11 16 11 2 13 0 0 3 2 2 3 0 16 9 3 13 14 13 9 1 9 1 9 2
20 1 10 0 12 9 13 15 3 1 12 11 13 14 13 9 1 9 1 9 2
14 9 4 13 1 9 1 10 0 9 1 9 0 9 2
20 1 9 13 9 3 10 9 1 12 9 2 10 9 1 12 9 1 10 9 2
13 1 0 9 4 15 13 1 15 9 4 13 1 2
22 7 9 13 16 11 13 1 1 14 13 15 0 0 2 1 10 9 1 0 12 9 2
16 15 13 16 9 13 3 1 10 9 1 9 1 0 12 9 2
12 15 13 0 0 0 9 7 9 7 0 9 2
19 11 11 7 11 13 15 1 1 9 1 12 9 2 10 0 9 1 15 2
20 11 13 1 10 9 10 9 1 12 9 2 10 9 1 12 9 1 10 9 2
13 9 13 3 1 1 1 15 10 14 4 13 9 2
17 11 13 0 0 9 1 9 2 7 4 0 13 15 0 1 9 2
35 10 0 9 1 10 0 9 13 11 9 1 11 2 16 11 1 10 0 9 1 9 11 13 3 1 14 13 0 9 1 0 9 1 12 2
22 10 0 12 9 4 11 7 11 13 9 2 7 10 10 9 13 1 1 14 13 1 2
18 1 11 13 1 0 7 11 7 11 1 1 14 13 15 1 10 9 2
17 1 9 4 11 13 1 9 1 14 13 10 0 9 1 0 0 2
12 3 11 1 10 10 9 13 3 1 14 13 2
6 4 13 9 1 11 5
2 0 2
21 9 11 11 13 3 1 14 13 11 1 1 10 0 9 2 16 11 11 11 13 2
3 13 1 2
16 9 11 11 13 1 11 1 10 0 9 9 1 9 1 9 2
10 11 13 15 0 9 1 1 10 9 2
14 1 0 9 13 3 11 1 9 1 10 0 7 11 2
16 9 11 11 7 11 11 13 1 10 9 9 1 10 0 9 2
13 3 13 11 1 14 13 9 0 2 1 12 9 2
16 2 10 0 9 1 15 13 14 13 9 7 9 1 1 11 2
18 3 13 15 11 1 10 1 10 0 0 9 14 13 1 2 13 15 2
18 7 9 13 3 0 1 16 9 4 13 9 1 10 0 9 1 12 2
5 13 9 1 11 5
16 2 15 13 1 1 11 11 11 2 7 3 15 4 13 9 2
21 15 13 15 1 10 9 1 10 0 9 2 15 13 0 1 11 1 0 0 9 2
31 0 9 1 11 11 7 11 11 11 4 0 13 1 9 1 14 13 11 1 1 10 0 9 1 14 13 11 7 11 0 2
8 7 3 4 11 13 9 1 2
29 3 13 3 9 1 9 2 7 1 11 9 13 11 1 0 9 1 14 13 11 1 1 9 1 10 0 9 11 2
17 16 10 0 13 0 1 11 2 13 11 15 0 0 11 7 11 2
17 9 13 3 1 10 0 9 1 11 1 12 1 9 12 0 9 2
21 1 11 13 11 11 0 16 15 3 13 0 1 11 14 13 1 10 9 1 11 2
18 2 15 13 16 11 3 13 3 0 1 0 9 15 13 0 1 15 2
11 3 0 13 15 9 1 9 2 13 15 2
26 11 13 16 9 1 9 13 0 0 2 7 16 15 13 0 0 9 1 10 9 10 0 4 13 1 2
13 2 10 0 13 3 10 0 9 10 10 9 13 2
19 7 15 13 3 1 10 9 1 0 9 1 14 13 1 11 2 13 15 2
4 0 1 11 5
37 11 11 11 4 13 9 0 1 9 1 16 15 4 13 1 9 2 7 4 3 4 13 15 1 15 9 9 9 4 13 1 1 1 9 1 9 2
21 11 13 10 1 0 15 13 0 1 1 10 9 1 9 11 1 9 13 1 1 2
13 2 11 13 10 0 9 2 15 4 15 3 13 2
23 7 0 13 15 10 9 15 4 13 15 0 1 15 14 13 1 11 7 11 2 13 15 2
5 0 9 1 11 5
4 15 13 1 2
25 11 4 13 0 0 9 1 11 2 7 9 13 16 9 13 1 15 15 4 4 13 1 1 9 2
2 0 2
26 9 1 11 7 9 1 11 2 11 11 2 13 0 0 1 16 9 11 11 13 11 1 1 0 9 2
23 2 10 10 9 4 13 10 9 1 11 2 7 10 0 9 4 13 10 9 2 13 15 2
27 0 12 9 1 9 13 15 3 0 9 1 10 0 7 10 0 1 11 2 1 10 9 1 11 1 9 2
23 16 9 4 13 1 2 13 10 0 0 1 14 13 1 7 11 7 11 1 14 13 9 2
16 11 13 1 10 0 1 14 13 16 11 7 11 13 1 9 2
26 10 0 1 9 4 13 1 11 2 7 13 3 0 1 15 10 15 13 15 4 4 13 1 7 13 2
2 9 5
22 16 11 13 1 9 1 11 1 11 2 13 3 9 1 2 9 2 3 0 1 11 2
18 11 9 1 11 2 11 11 2 13 3 16 11 13 1 9 1 11 2
28 2 9 1 15 13 10 9 1 11 2 11 7 11 2 13 11 2 15 3 3 13 9 1 9 1 10 0 2
30 15 13 3 16 15 13 0 1 9 15 15 13 1 9 2 15 13 10 9 1 11 2 11 2 11 7 11 10 11 2
27 7 11 13 3 9 1 16 15 13 15 14 13 1 11 1 11 7 11 4 13 10 9 15 13 11 0 2
18 2 15 4 3 13 10 9 15 13 0 0 1 0 9 2 13 11 2
33 9 11 9 13 14 13 3 1 11 2 11 7 11 2 7 9 13 3 3 1 9 1 9 1 11 2 3 0 9 13 1 9 2
27 2 15 13 3 0 14 13 1 10 0 9 2 3 0 11 13 1 7 13 1 9 1 9 1 0 9 2
28 7 3 0 15 13 1 9 1 9 2 13 15 0 1 14 13 1 11 2 13 11 9 1 11 2 11 11 2
5 2 0 1 11 5
34 11 11 2 9 1 11 7 9 1 11 2 13 3 15 1 16 9 11 11 1 9 11 13 11 1 1 0 9 2 7 0 7 0 2
37 15 13 10 0 1 11 3 4 13 1 9 1 9 1 0 9 2 7 13 1 16 11 9 1 14 13 1 11 4 13 9 1 1 10 0 9 2
20 2 10 10 9 4 13 10 9 1 11 2 7 10 0 9 4 13 10 9 2
37 9 13 0 9 7 9 1 11 1 12 16 15 3 3 4 13 11 7 11 1 14 13 15 0 2 7 13 1 0 9 7 13 10 0 0 9 2
12 10 0 9 4 13 1 2 7 0 7 0 2
19 1 9 13 15 3 14 13 3 1 16 9 13 3 0 0 2 13 11 2
5 2 13 3 11 5
34 7 4 9 9 13 9 3 2 7 3 4 15 13 15 3 1 11 2 13 11 2 15 0 1 3 13 1 1 10 0 9 1 9 2
40 2 11 13 0 1 14 13 1 1 10 9 1 9 2 7 10 9 1 15 4 13 9 1 9 1 9 2 3 16 15 13 9 1 1 9 1 9 7 9 2
30 9 11 11 13 10 0 9 2 7 13 1 9 2 9 2 9 1 0 9 7 9 7 1 9 7 9 2 13 11 2
46 11 1 10 9 2 13 9 7 9 1 0 9 1 10 1 9 15 4 13 0 1 11 14 13 1 10 0 1 2 3 1 11 15 11 13 1 2 7 9 2 15 10 0 4 13 2
23 2 9 13 0 1 15 2 7 15 15 13 1 14 13 0 1 1 0 9 1 10 0 2
55 3 13 15 0 1 16 0 9 1 9 4 13 1 9 2 7 15 4 3 13 1 1 14 13 1 0 9 2 13 11 9 11 11 2 15 13 0 1 16 15 1 10 9 3 4 13 9 1 10 0 1 14 13 9 2
21 11 13 3 10 9 1 11 1 11 2 1 9 7 9 1 11 11 2 11 11 2
36 15 13 11 0 1 1 9 2 3 0 15 13 1 1 9 2 7 13 0 1 16 15 13 11 15 13 9 1 9 1 10 0 0 0 9 2
12 2 15 13 11 15 13 9 3 2 13 11 2
6 0 13 1 0 9 5
4 13 1 9 2
10 1 0 9 13 9 9 1 0 9 2
6 3 13 15 0 9 2
13 2 9 1 0 9 1 11 4 3 13 1 9 2
10 9 4 4 13 9 1 9 0 2 2
15 3 13 15 1 10 0 9 1 9 2 15 13 0 9 2
15 1 9 4 15 3 13 15 16 9 1 10 9 4 13 2
28 1 9 1 11 11 2 11 11 11 2 13 7 11 9 1 11 2 11 2 7 11 11 11 2 11 2 9 2
13 2 13 9 9 16 15 13 0 9 4 13 9 2
18 2 15 4 3 13 16 15 4 13 1 10 9 1 9 10 0 9 2
13 3 13 3 15 1 9 7 13 1 1 10 9 2
14 7 15 15 13 3 13 16 15 13 1 1 0 9 2
12 7 15 4 13 0 1 2 13 11 1 11 2
11 9 11 11 1 11 13 10 10 1 11 2
10 1 15 13 10 0 9 3 12 9 2
6 3 0 9 1 9 5
11 2 15 13 1 12 9 1 1 0 9 2
32 1 9 1 13 15 0 15 13 15 1 2 7 3 1 0 9 13 9 0 1 9 1 9 16 15 4 13 1 2 13 11 2
21 1 10 0 9 1 12 13 9 9 1 16 11 4 13 1 15 0 7 0 9 2
9 3 4 9 9 13 1 0 9 2
21 3 1 12 13 11 11 9 1 14 13 0 0 1 0 9 2 1 1 10 11 2
10 7 15 13 14 13 0 9 1 15 2
22 7 1 9 13 9 9 7 13 1 10 9 2 15 9 11 11 11 13 0 0 1 2
7 2 15 4 13 1 9 2
25 15 13 10 9 7 13 9 15 13 1 9 15 10 0 7 0 9 3 13 2 13 11 1 11 2
22 3 9 1 9 2 11 11 2 11 2 2 4 13 1 9 0 9 1 10 0 9 2
15 15 13 15 1 11 7 1 10 9 1 9 1 9 12 2
15 2 15 4 13 9 2 15 13 15 9 13 0 0 1 2
47 7 3 4 3 15 13 10 0 9 1 15 15 13 0 9 2 7 3 15 13 9 1 16 9 4 13 1 1 9 2 13 15 7 13 9 1 3 0 9 4 13 1 9 1 0 9 2
3 9 12 5
4 9 7 9 5
3 12 9 5
10 9 4 13 0 1 0 1 12 9 2
23 15 4 4 13 1 0 0 7 0 9 7 4 13 1 9 7 9 1 11 10 9 9 2
23 10 0 0 9 1 12 13 1 11 12 11 7 9 16 11 0 9 4 13 10 0 9 2
15 16 9 4 13 1 12 2 13 11 3 0 14 13 9 2
26 0 4 15 4 13 0 9 1 14 13 9 2 7 15 1 9 4 13 0 2 0 2 9 1 11 2
17 9 4 3 4 13 1 0 9 15 4 13 11 0 9 0 9 2
16 1 9 4 10 0 0 9 13 14 13 9 1 10 0 9 2
15 11 13 1 12 10 9 15 4 13 9 1 9 7 9 2
28 9 13 1 10 9 11 9 2 0 9 1 12 2 1 10 0 9 1 10 0 9 1 9 1 9 7 9 2
15 1 10 0 9 15 13 13 15 0 0 9 1 9 9 2
8 9 4 13 1 11 9 12 2
29 11 13 14 13 1 9 1 0 9 2 7 13 0 16 15 4 13 10 0 9 1 14 13 9 1 9 7 9 2
23 1 12 4 15 1 11 13 14 13 10 0 0 0 9 1 14 13 9 1 9 7 9 2
18 9 13 1 10 9 1 1 15 2 7 10 0 11 13 15 1 9 2
16 9 13 1 9 7 13 1 9 12 10 0 9 1 12 9 2
3 12 9 5
11 11 4 13 1 0 9 1 0 9 12 2
36 9 13 10 0 9 1 9 1 10 10 0 9 1 11 2 0 9 2 10 0 9 2 11 11 2 11 11 2 0 9 7 9 1 0 9 2
14 12 1 9 4 13 1 9 1 10 0 9 1 11 2
7 9 13 0 9 1 9 2
10 2 9 11 11 2 11 2 9 2 5
10 2 9 11 11 2 11 2 9 2 5
7 2 9 11 11 2 11 5
7 2 9 11 11 2 11 5
7 2 9 11 11 2 11 5
7 2 9 11 11 2 11 5
8 2 9 11 11 11 2 11 5
7 2 9 11 11 2 11 5
7 2 9 11 11 2 11 5
7 2 9 11 11 2 11 5
7 2 9 11 11 2 11 5
9 2 9 11 11 2 11 5 11 5
7 2 9 11 11 2 11 5
7 2 9 11 11 2 11 5
7 2 9 11 11 2 11 5
8 2 9 11 11 11 2 11 5
7 2 9 11 11 2 11 5
7 2 9 11 11 2 11 5
7 2 9 11 11 2 11 5
12 2 9 11 11 2 11 2 1 9 12 2 5
12 2 9 11 11 2 11 2 1 9 12 2 5
3 12 9 5
5 9 13 0 9 2
21 2 9 1 9 13 14 13 9 1 14 13 9 16 9 4 13 2 13 7 13 2
21 15 13 1 9 16 11 0 9 3 4 13 10 0 2 0 2 0 7 0 9 2
9 1 9 1 9 2 4 9 13 2
14 12 9 1 10 9 3 15 4 13 7 13 1 11 2
18 12 0 7 0 9 1 9 1 15 15 1 9 4 13 1 10 9 2
13 12 9 1 9 7 9 1 10 0 9 1 9 2
21 12 9 1 0 9 2 3 9 13 1 9 2 9 2 9 7 0 5 0 9 2
3 12 9 2
10 12 9 1 9 1 0 7 0 9 2
21 12 9 1 9 7 9 2 10 0 9 2 9 9 3 1 10 0 9 1 9 2
40 12 10 9 0 9 1 9 13 14 13 1 1 10 9 1 11 0 9 2 1 10 0 9 2 1 0 9 7 9 2 1 10 9 7 1 9 1 10 9 2
24 15 13 16 9 1 9 1 10 9 13 1 0 9 1 0 9 1 11 7 5 7 10 9 2
36 15 4 13 10 9 1 9 14 13 9 15 4 13 0 0 9 7 15 13 16 9 9 13 14 13 10 9 1 9 7 16 9 9 3 13 2
13 9 4 13 15 1 9 1 9 7 11 0 9 2
22 15 4 13 0 9 1 9 1 9 2 1 16 15 3 13 16 9 13 0 9 0 2
18 15 13 0 16 9 13 1 9 1 0 9 7 10 0 9 1 9 2
10 9 4 13 9 1 0 7 0 9 2
30 15 4 13 1 10 9 15 13 15 0 16 15 2 1 11 2 4 13 9 1 10 9 15 13 1 10 9 0 9 2
12 9 4 13 1 10 9 1 9 1 12 2 2
6 12 9 9 1 9 5
16 1 9 9 4 9 13 9 3 15 13 0 7 13 1 11 2
27 9 4 3 13 7 13 10 9 1 11 0 9 9 2 7 3 7 0 13 1 9 15 13 9 1 9 2
20 9 4 13 9 1 9 9 2 7 13 3 9 0 13 4 13 7 13 15 2
27 1 14 13 9 1 9 1 0 9 7 0 9 2 4 9 13 15 0 14 13 9 1 10 9 7 9 2
35 9 4 1 0 9 13 9 1 9 7 11 0 9 2 7 4 3 3 13 10 0 9 1 9 7 9 1 10 0 9 1 11 0 9 2
28 9 1 10 10 9 13 16 10 9 1 9 13 14 13 10 9 1 14 13 16 9 4 13 2 13 7 13 2
24 9 4 3 13 7 1 9 13 9 1 9 15 0 7 0 4 13 9 1 9 9 1 9 2
14 0 7 0 9 1 11 0 9 4 3 13 1 9 2
15 9 13 16 2 2 15 4 13 0 9 1 9 1 9 2
15 2 10 0 9 4 13 1 1 0 9 1 9 1 12 2
18 9 4 3 13 9 9 7 0 9 1 9 1 9 1 9 7 9 2
16 1 9 4 9 13 9 2 9 7 9 2 1 9 1 9 2
14 10 0 0 0 9 13 2 11 8 11 8 11 2 2
18 15 13 1 9 14 13 7 13 10 0 9 7 9 1 10 0 9 2
22 9 13 16 10 10 9 13 1 9 16 10 0 9 1 9 7 11 0 9 4 13 2
14 9 13 16 9 4 13 15 1 10 9 1 9 9 2
23 2 15 13 1 9 16 11 0 9 3 4 13 10 0 2 0 2 0 7 0 9 2 2
18 10 9 4 13 1 11 7 13 1 1 9 1 11 1 10 0 9 2
31 9 4 3 3 13 15 1 10 9 14 13 0 9 1 3 11 0 9 13 15 1 9 7 13 9 1 11 0 9 9 2
9 9 9 13 0 0 1 9 9 2
17 9 7 9 9 1 9 7 9 1 12 2 12 13 9 9 3 2
24 2 9 13 10 9 15 4 13 7 1 10 9 15 13 7 1 10 9 15 13 0 1 9 2
27 1 9 13 10 9 3 9 13 9 1 9 7 9 2 7 3 3 10 9 15 13 10 0 9 1 9 2
29 9 1 9 13 3 10 9 3 15 1 9 1 9 13 0 9 7 9 1 14 4 13 9 7 13 9 1 9 2
47 15 4 3 3 13 9 1 16 1 0 9 1 9 13 3 9 2 9 2 1 10 9 3 9 4 13 9 1 0 9 1 9 2 9 7 9 1 16 15 13 9 1 10 0 9 2 2
7 15 13 3 10 0 9 2
19 9 9 13 7 1 0 7 0 9 1 11 0 9 7 13 1 0 9 2
30 15 13 9 1 9 1 16 15 3 13 0 1 10 0 9 1 9 1 14 4 13 9 1 9 7 9 7 13 9 2
15 9 4 13 16 11 0 9 3 13 0 9 1 9 9 2
34 9 13 3 9 1 14 13 10 9 1 2 9 2 7 2 9 2 1 0 9 2 7 14 13 9 1 10 0 9 1 10 10 9 2
18 3 0 13 15 0 1 9 1 15 15 3 13 9 1 11 0 9 2
40 9 4 3 13 14 13 2 9 2 1 9 1 9 1 10 0 9 1 14 13 16 11 0 9 4 13 10 9 1 9 0 1 9 1 9 1 9 7 9 2
28 9 13 16 2 2 2 9 1 9 1 10 9 13 1 0 9 1 0 9 1 11 7 5 7 10 9 2 2
29 9 4 13 1 15 2 7 3 13 10 0 9 15 10 0 9 13 1 9 2 11 0 9 7 10 9 7 9 2
17 9 12 2 12 1 9 13 0 9 1 0 2 0 7 0 9 2
30 9 1 0 9 2 9 2 9 1 9 1 0 7 0 9 7 9 1 9 2 9 7 10 9 1 0 9 1 9 2
17 9 7 9 1 9 1 0 7 0 9 4 13 0 1 0 9 2
22 9 1 0 9 7 9 13 3 0 1 10 0 9 1 9 1 9 7 11 0 9 2
22 9 13 16 9 4 13 0 9 15 3 13 0 1 9 9 7 15 3 13 9 9 2
19 15 13 1 9 1 10 0 9 1 0 9 2 1 9 9 7 0 9 2
21 9 13 16 9 4 13 1 10 9 2 7 9 4 13 9 1 0 7 0 9 2
18 10 9 4 9 1 3 9 13 3 1 12 9 9 2 3 9 12 2
42 9 13 0 14 13 15 1 14 13 12 9 2 7 16 0 9 4 13 0 9 7 9 1 0 2 7 16 15 4 13 15 0 1 9 14 13 10 0 7 0 9 2
34 9 13 15 4 13 0 14 13 9 7 13 0 9 1 16 15 4 13 1 9 1 10 0 0 2 0 7 0 9 15 9 4 13 2
4 12 9 9 5
13 9 4 13 1 15 12 9 2 13 1 12 9 2
36 9 12 4 9 9 13 1 10 12 9 9 1 11 2 11 7 11 2 3 15 4 13 9 1 9 1 0 7 0 9 7 10 9 7 9 2
8 9 1 9 13 1 1 9 2
16 1 0 1 9 4 9 1 4 13 1 14 13 9 1 9 2
10 9 4 3 13 10 0 9 1 11 2
61 9 9 2 9 1 9 7 9 4 1 1 9 13 1 0 9 1 9 7 9 7 13 9 1 10 9 9 2 9 7 9 1 11 0 9 7 1 9 3 2 1 9 1 9 9 1 16 9 13 1 9 1 0 9 7 10 0 9 1 9 2
28 1 14 13 16 10 9 1 9 4 13 1 0 9 2 4 10 0 9 1 9 4 13 1 10 9 7 9 2
10 10 9 1 9 9 4 13 9 12 2
10 9 4 13 9 7 9 1 0 9 2
11 0 1 15 4 13 9 1 9 1 9 2
9 10 9 1 10 2 13 1 9 2
3 12 9 5
14 9 4 13 1 11 7 13 0 0 1 0 9 12 2
18 1 1 0 9 12 4 15 13 1 11 11 2 1 11 11 1 9 2
21 11 11 13 3 1 11 7 11 2 16 11 11 4 13 9 1 11 11 1 11 2
9 11 13 1 1 9 0 9 12 2
20 1 3 1 4 9 4 13 1 11 11 15 4 13 9 1 9 1 0 9 2
33 1 0 9 12 4 10 12 9 11 11 2 11 11 2 11 11 7 11 11 13 10 9 15 4 13 9 1 14 13 9 1 9 2
23 1 0 9 12 4 9 11 11 2 1 9 1 9 7 9 2 13 1 12 9 1 9 2
17 11 11 4 13 1 9 1 9 7 9 1 9 1 0 9 12 2
23 9 4 1 0 9 13 0 9 1 0 9 2 7 1 0 9 2 9 7 0 0 9 2
12 9 9 1 11 4 13 1 0 7 0 9 2
3 9 12 5
2 9 5
4 12 9 9 5
4 12 0 9 5
20 9 1 9 13 14 13 9 1 14 13 9 16 9 4 13 2 13 7 13 2
23 9 9 1 12 9 13 16 9 9 13 2 7 16 15 13 10 0 9 1 11 0 9 2
19 10 9 1 15 2 12 9 2 13 16 11 0 9 13 1 10 0 9 2
19 10 9 1 15 2 12 9 2 13 16 11 0 9 13 1 10 0 9 2
11 12 9 13 16 9 9 13 1 0 9 2
3 0 9 5
44 9 9 1 10 0 9 13 16 11 0 9 1 9 13 2 7 16 11 0 9 13 10 0 9 1 10 9 7 1 0 9 1 10 9 15 13 1 9 9 7 9 14 13 2
16 9 13 1 9 10 9 2 1 9 1 10 0 9 7 9 2
18 11 0 9 13 3 10 0 9 1 9 1 10 9 2 13 1 11 2
16 9 13 16 10 9 13 1 10 0 9 7 13 1 10 9 2
14 9 13 1 1 10 10 9 7 1 10 0 0 9 2
17 1 9 1 9 9 13 15 0 0 14 13 9 9 1 0 9 2
14 15 13 3 0 14 13 9 1 0 9 1 11 9 2
25 9 13 16 10 0 9 13 9 15 11 0 9 13 1 9 9 7 13 9 1 0 7 0 9 2
24 0 13 9 16 9 2 1 9 1 10 9 7 9 2 13 10 9 1 10 9 0 1 9 2
32 9 13 0 9 1 16 11 0 9 3 4 13 10 0 9 1 0 9 7 1 9 1 0 9 1 9 7 9 1 10 9 2
24 9 9 7 9 1 9 4 13 3 16 15 4 13 10 9 1 9 7 13 10 9 1 9 2
14 1 10 0 9 4 9 0 9 13 1 1 10 9 2
18 9 13 10 9 15 4 13 10 9 15 11 2 9 2 1 9 13 2
17 9 4 3 13 16 15 13 9 1 9 15 13 7 9 7 9 2
18 9 1 9 7 9 13 1 9 1 0 0 1 9 1 9 7 9 2
23 10 9 13 3 7 0 1 16 9 13 14 13 10 9 1 10 9 15 13 9 1 9 2
22 15 13 9 9 1 9 15 13 0 1 9 9 2 3 9 1 9 1 9 7 9 2
33 7 1 10 9 9 13 9 1 10 9 2 13 9 16 10 0 9 13 11 0 9 10 0 9 1 10 0 9 1 9 7 9 2
18 9 13 15 1 10 9 16 10 0 9 4 13 9 1 9 7 9 2
18 9 1 9 2 1 0 9 1 9 2 13 10 0 9 1 9 9 2
3 0 9 5
25 9 12 9 1 12 1 12 9 13 10 9 1 9 7 13 10 0 9 1 9 1 10 0 9 2
29 15 13 16 11 0 9 3 0 13 10 9 1 9 2 7 13 1 10 0 9 1 0 9 1 10 9 7 9 2
12 9 13 1 10 0 9 1 10 9 7 9 2
43 10 9 13 0 9 1 16 11 0 9 0 1 4 13 7 13 1 10 9 7 16 0 9 3 4 13 15 15 13 9 9 2 9 7 9 14 13 1 1 1 10 9 2
27 1 10 9 9 13 15 10 9 15 13 15 0 2 0 15 10 0 13 9 1 9 1 10 9 7 9 2
3 0 9 5
19 9 10 9 1 12 1 12 9 13 10 3 0 9 1 9 1 9 9 2
13 15 13 10 9 1 9 9 3 16 9 9 13 2
44 1 10 9 9 13 15 9 9 15 0 13 16 11 0 9 13 3 1 15 15 13 15 2 7 15 0 13 10 0 0 9 1 16 15 4 4 13 15 1 1 9 1 9 2
43 10 9 13 15 13 1 0 9 16 11 9 15 13 9 13 2 7 13 16 9 1 9 15 13 10 0 9 7 10 0 9 4 13 10 0 9 15 15 3 13 9 1 2
2 9 5
17 1 10 9 1 9 1 10 0 9 2 13 11 9 12 10 9 2
18 10 9 13 1 0 9 10 9 1 9 2 7 4 1 0 13 3 2
14 1 9 4 9 13 9 15 13 16 9 9 3 13 2
25 10 9 1 12 9 13 16 15 13 10 0 9 1 11 15 13 10 0 9 1 0 7 0 9 2
51 10 9 1 12 9 13 10 0 9 15 13 1 0 9 7 1 9 2 16 10 10 9 1 12 9 13 15 3 13 9 1 10 0 9 1 11 9 12 15 13 1 9 0 0 9 2 0 7 10 2 2
25 10 10 9 1 12 9 13 16 9 1 9 12 13 1 15 15 13 1 9 1 9 1 0 9 2
5 9 9 7 9 5
23 16 9 9 13 2 13 9 1 10 0 0 9 7 9 7 10 9 4 3 13 1 0 2
20 10 9 1 12 9 13 16 9 9 1 14 13 10 0 0 9 7 9 13 2
28 9 13 15 4 13 10 0 9 1 10 9 7 9 2 7 13 16 15 13 10 9 15 13 0 0 1 9 2
27 10 9 13 16 15 7 13 0 7 0 14 13 10 10 9 16 9 1 9 7 9 4 13 1 10 9 2
3 12 9 5
29 9 13 15 13 10 0 9 14 13 0 7 1 10 9 13 1 0 1 9 7 9 9 2 3 15 13 1 9 2
50 1 9 0 9 2 10 0 9 2 13 10 9 1 12 9 16 0 9 13 1 9 2 1 0 9 15 13 9 7 0 9 1 10 0 0 7 0 9 15 13 9 2 9 2 9 7 9 1 9 2
15 15 13 1 10 0 9 15 4 13 9 1 9 0 9 2
14 10 9 13 16 10 0 9 1 10 9 13 1 9 2
18 10 10 9 13 10 9 1 10 9 2 13 1 0 9 1 0 9 2
3 12 9 5
34 9 1 12 1 12 9 13 16 9 13 3 16 9 13 16 9 13 9 1 9 2 16 9 13 10 0 9 15 4 13 1 10 0 2
28 9 13 10 0 7 0 0 9 2 7 9 1 10 0 7 0 9 1 9 7 10 0 7 0 9 13 0 2
13 0 13 11 0 9 13 1 10 0 7 0 9 2
24 15 13 3 16 9 4 13 9 1 11 0 9 1 14 13 9 1 0 9 3 15 13 0 2
39 9 9 1 12 1 12 9 13 16 0 9 13 9 2 7 16 0 10 0 9 13 1 11 0 9 9 7 16 9 7 9 13 10 0 9 10 0 9 2
36 9 13 16 15 3 3 4 13 10 9 1 9 1 9 1 14 13 9 1 1 9 2 7 16 10 0 13 0 1 9 0 9 13 9 1 2
16 9 13 16 9 9 1 9 13 1 10 0 9 9 7 9 2
27 15 4 13 14 13 9 1 0 9 1 9 1 9 1 14 13 16 9 1 9 13 1 0 9 7 9 2
20 15 13 10 0 9 1 14 13 0 0 7 0 9 7 9 1 10 0 9 2
24 9 13 3 16 15 13 10 0 9 1 10 9 5 9 1 0 9 1 9 1 9 5 9 2
22 9 4 13 0 9 1 9 1 10 0 1 9 7 9 2 0 9 7 9 1 9 2
6 12 0 7 0 9 5
22 9 7 9 13 3 3 10 9 1 9 1 10 0 9 7 1 9 7 9 1 9 2
15 3 0 13 15 10 9 1 9 2 9 2 9 7 9 2
8 9 9 13 1 9 0 9 2
29 1 1 0 9 13 9 15 4 13 0 9 1 0 7 0 9 2 0 1 10 0 9 1 9 7 11 0 9 2
25 9 13 16 15 2 1 9 1 9 9 1 0 9 2 13 10 0 0 0 9 0 10 0 9 2
14 9 4 0 13 1 9 16 10 9 4 13 7 13 2
29 9 13 16 10 10 9 2 0 1 0 9 2 13 1 0 0 9 15 13 9 1 9 1 9 7 5 7 9 2
9 11 4 13 15 1 10 0 9 2
27 10 9 1 12 1 12 9 13 3 9 1 0 0 9 1 9 9 1 14 13 0 9 7 9 1 9 2
17 9 13 16 10 9 4 4 13 1 10 9 1 9 0 1 9 2
12 15 4 4 13 9 7 9 15 13 15 0 2
18 9 13 16 9 13 9 1 0 7 0 9 15 13 1 1 0 9 2
13 9 13 16 15 13 10 0 9 1 11 0 9 2
10 9 4 13 1 9 1 0 0 9 2
3 12 9 5
4 9 7 9 5
29 9 13 1 9 16 11 0 9 1 10 0 9 13 10 10 9 2 7 16 9 3 0 4 13 0 9 7 9 2
27 9 9 13 9 1 11 0 9 0 7 0 4 13 1 10 9 1 9 1 9 9 1 9 7 0 9 2
32 9 13 16 15 1 10 0 9 13 10 0 9 2 16 9 2 0 9 7 9 4 13 1 1 9 1 9 2 1 1 9 2
11 15 4 15 13 9 1 1 10 0 9 2
6 11 9 2 11 2 5
25 9 13 16 9 1 9 1 11 3 4 13 1 0 9 2 7 4 13 1 10 0 9 1 11 2
15 9 1 12 1 12 9 13 16 11 13 1 11 0 9 2
26 9 13 1 9 16 10 9 1 11 1 11 0 9 3 13 10 9 7 9 10 9 1 0 0 9 2
11 10 9 13 11 1 9 9 7 9 9 2
22 9 15 1 9 13 1 0 9 13 1 11 0 9 2 16 10 13 1 9 7 13 2
5 12 0 1 9 5
4 12 0 9 5
15 1 9 12 13 15 9 1 9 9 1 9 1 10 9 2
23 3 1 12 9 3 4 9 13 1 10 0 0 9 1 9 7 0 13 1 9 1 9 2
7 9 9 4 13 9 9 2
15 9 13 0 9 2 7 9 13 10 9 1 10 0 9 2
16 1 9 1 9 13 9 1 10 9 7 13 15 0 0 9 2
20 9 7 9 13 1 9 1 9 10 12 0 9 1 9 15 7 13 7 13 2
13 1 9 13 9 10 9 1 10 0 9 1 9 2
9 9 13 0 9 7 0 7 0 2
12 9 4 13 2 7 9 13 0 2 0 2 2
16 11 9 13 1 9 1 10 0 9 7 9 1 10 0 9 2
6 1 9 4 9 13 2
20 9 13 10 0 9 1 10 0 9 9 1 9 7 9 2 1 11 9 2 2
18 9 1 9 13 9 1 10 0 9 7 13 15 9 1 9 0 9 2
13 9 7 9 13 9 15 11 7 11 4 13 15 2
10 9 7 9 13 0 9 1 0 9 2
17 9 13 0 0 2 7 0 9 4 13 1 10 9 1 9 9 2
19 9 1 12 4 0 13 1 10 9 1 9 1 0 9 7 9 1 9 2
13 10 0 0 9 1 12 13 10 0 7 0 9 2
16 9 9 13 10 0 9 2 7 10 0 9 13 3 0 9 2
11 1 10 0 9 4 9 9 7 9 13 2
20 11 13 16 10 0 9 3 4 13 9 0 9 2 7 9 4 3 0 13 2
26 16 9 0 4 13 10 9 1 11 2 4 3 11 13 14 13 10 9 1 2 9 2 2 9 2 2
32 1 9 1 9 4 15 13 9 1 9 15 4 13 11 0 9 0 0 9 7 9 2 7 1 12 4 15 13 14 13 9 2
8 7 11 13 11 9 1 9 2
16 9 7 9 13 3 0 0 0 2 7 9 9 4 3 13 2
10 1 12 13 10 0 11 11 1 12 2
22 0 9 7 3 3 9 4 3 13 0 2 7 9 4 13 9 1 9 9 7 9 2
6 1 12 4 9 13 2
25 15 13 0 9 0 9 1 14 13 15 1 1 9 7 1 0 9 13 10 0 9 1 0 9 2
18 1 9 1 9 1 12 13 3 0 9 9 1 14 13 15 1 11 2
16 10 0 9 2 15 13 9 9 1 9 2 4 13 1 12 2
10 10 0 9 1 9 4 13 1 12 2
9 3 1 12 13 9 9 1 9 2
16 11 8 8 8 8 8 4 13 1 12 7 13 9 1 12 2
20 9 1 9 1 9 1 10 0 7 0 9 13 1 16 9 4 13 1 9 2
6 9 13 10 0 9 2
12 15 13 3 9 2 16 11 13 9 0 9 2
18 11 9 4 13 1 9 2 15 1 3 1 13 10 0 9 1 11 2
15 11 13 10 0 9 2 7 4 3 3 13 9 1 9 2
29 1 9 4 10 0 9 0 13 7 9 13 2 7 15 13 0 1 9 16 15 13 10 0 9 0 7 0 9 2
17 1 9 13 9 1 9 7 9 1 0 0 9 0 9 1 9 2
27 9 7 10 0 9 13 10 0 9 9 12 7 13 10 9 1 9 1 9 1 11 7 1 9 1 9 2
13 9 11 11 13 9 7 9 9 7 0 7 0 2
13 9 9 13 2 16 11 13 1 7 9 7 9 2
28 11 11 13 16 9 3 4 13 9 1 9 1 0 9 2 7 16 9 3 4 13 9 1 9 9 7 9 2
26 1 9 13 11 0 9 1 10 0 9 1 0 9 12 7 1 1 9 2 16 9 3 13 1 9 2
19 0 0 7 0 9 13 0 9 1 9 1 9 7 9 1 9 1 9 2
24 9 13 1 9 1 11 10 9 9 2 7 15 4 3 13 0 9 1 11 1 14 13 9 2
20 9 4 3 4 13 1 0 9 15 3 4 13 9 0 9 7 9 1 9 2
18 1 16 9 4 4 13 2 4 9 1 9 1 9 7 9 13 0 2
39 0 4 9 13 7 13 9 2 16 9 1 11 0 9 7 10 0 9 4 13 0 2 7 16 9 0 13 3 4 13 1 14 4 13 1 10 0 9 2
12 9 1 10 0 0 9 4 13 9 1 9 2
20 3 0 4 9 13 1 9 1 10 9 7 10 9 1 9 1 10 0 9 2
3 12 9 5
16 1 9 12 13 11 0 9 1 9 7 9 2 7 9 13 2
15 9 1 10 0 9 7 9 13 7 9 13 1 1 11 2
37 3 13 9 7 9 2 9 2 1 0 9 1 10 9 15 13 1 11 0 9 2 10 9 7 9 7 10 0 9 2 1 9 1 10 0 9 2
6 11 0 9 1 9 5
16 11 0 9 13 3 7 0 10 9 2 13 1 10 0 9 2
20 15 13 10 0 9 0 1 10 0 9 2 7 1 10 9 13 1 10 9 2
10 10 0 9 13 1 11 7 12 9 2
18 11 0 9 13 1 9 14 13 10 0 2 0 2 0 7 0 9 2
13 1 1 10 0 9 2 4 9 13 1 0 9 2
23 9 4 13 9 9 2 13 15 1 9 1 14 13 9 7 13 9 7 9 9 7 9 2
12 3 4 15 13 0 3 1 14 13 0 9 2
33 1 9 1 14 13 11 0 9 9 2 4 9 3 13 10 9 1 10 9 7 9 7 1 9 15 3 13 9 1 11 0 9 2
2 9 5
12 1 0 9 13 11 0 9 3 10 10 9 2
26 15 4 0 13 13 1 11 9 2 7 10 9 2 9 3 4 13 7 13 1 9 2 9 7 9 2
20 11 0 9 4 13 1 10 9 1 9 2 7 13 10 0 9 9 7 9 2
23 11 1 0 9 13 0 13 9 0 9 2 7 0 1 9 4 1 9 13 1 1 11 2
26 11 0 9 13 1 9 3 1 10 0 9 2 3 14 13 9 2 13 9 7 13 3 9 13 9 2
28 13 1 9 9 13 9 3 7 0 10 0 9 2 13 1 10 9 9 1 11 7 0 13 1 9 7 9 2
44 1 3 13 15 10 0 7 0 9 2 15 3 3 13 9 1 11 0 9 7 10 0 9 2 9 2 9 7 9 2 2 7 3 1 9 13 9 9 2 9 2 9 3 2
30 9 13 1 9 1 2 2 11 9 12 10 9 2 1 16 10 0 9 13 2 9 0 11 2 1 10 9 15 13 2
51 2 11 9 1 2 11 9 2 2 9 12 2 12 2 12 2 12 3 2 2 15 13 11 2 9 2 9 1 11 0 9 1 9 2 9 3 2 11 13 1 11 7 9 13 1 11 1 9 7 9 2
2 9 5
10 10 0 9 13 10 0 7 0 9 2
25 0 15 15 13 10 9 2 13 15 3 10 9 1 0 9 1 9 2 1 7 0 7 0 9 2
23 0 13 13 10 0 9 3 9 1 9 2 3 16 15 0 13 7 13 1 0 7 0 2
18 9 13 0 1 10 0 0 9 2 9 2 7 0 9 2 9 2 2
8 3 4 9 13 1 12 9 2
7 15 13 7 9 7 9 2
28 1 9 1 10 12 9 13 15 3 9 2 1 0 9 2 0 9 7 1 0 9 2 9 7 10 0 9 2
20 1 9 1 10 0 0 9 2 13 15 3 10 0 9 7 9 1 9 9 2
17 9 13 10 0 9 16 9 4 13 0 1 9 7 0 1 9 2
14 9 13 9 7 9 10 0 9 9 2 9 7 9 2
12 9 4 3 13 2 7 1 10 0 10 9 2
12 15 13 12 9 1 0 2 9 7 10 10 2
26 9 4 0 13 2 3 1 11 1 9 1 9 2 9 7 9 2 2 7 3 1 0 9 1 9 2
21 10 10 0 1 9 4 0 13 1 9 10 9 1 10 0 9 1 10 0 9 2
38 1 9 1 10 0 9 7 10 0 0 9 13 15 10 9 0 0 9 2 9 3 15 13 15 1 9 1 11 0 9 2 1 0 0 7 0 9 2
11 15 13 10 0 7 0 9 1 9 9 2
2 9 5
12 11 0 9 4 3 13 0 9 1 1 9 2
14 0 4 3 10 0 9 1 9 13 1 11 0 9 2
14 1 12 13 1 12 9 1 9 0 9 1 10 9 2
10 10 3 0 0 13 9 1 10 9 2
15 1 9 4 9 9 1 11 0 9 13 1 1 12 9 2
10 9 15 3 13 10 9 7 9 13 2
17 1 12 13 10 9 12 9 2 16 9 1 9 13 3 12 9 2
4 9 7 9 5
14 1 10 0 12 9 4 15 13 10 9 9 1 11 2
15 10 0 9 9 1 11 0 9 2 13 10 10 0 9 2
17 0 1 10 12 0 9 4 11 13 15 1 14 13 10 0 9 2
30 1 9 1 10 0 0 9 1 9 7 11 1 12 2 4 7 9 2 9 2 9 7 9 13 10 0 9 1 11 2
13 1 12 4 11 11 13 1 10 0 9 1 11 2
4 10 0 9 5
10 1 10 0 9 13 15 0 0 9 2
29 0 9 4 0 13 13 1 9 15 13 9 7 9 0 9 1 14 13 10 9 7 10 9 1 10 0 0 9 2
11 11 13 3 10 9 15 13 1 10 0 2
26 11 13 3 1 1 10 0 0 9 2 15 3 4 13 1 11 2 7 15 13 0 9 1 10 9 2
8 0 9 13 1 11 7 11 2
4 9 7 9 5
25 1 10 9 13 9 7 9 2 9 2 10 0 9 2 13 1 0 9 1 10 1 10 0 9 2
22 9 7 9 4 0 13 0 1 9 2 7 4 1 10 0 9 4 13 1 0 0 2
24 9 1 9 7 9 13 10 0 9 1 9 2 7 10 0 9 1 9 1 16 15 4 13 2
11 9 7 9 13 7 10 0 7 0 9 2
19 1 15 13 7 10 9 1 9 7 1 0 14 4 13 10 9 7 9 2
13 0 13 15 9 1 14 13 15 1 9 7 9 2
25 9 7 9 4 3 13 1 9 16 15 13 1 14 13 0 9 2 9 2 9 7 10 0 9 2
14 10 0 9 13 16 9 13 11 0 9 9 1 9 2
7 15 13 15 0 9 1 2
33 10 0 0 9 13 15 1 16 10 0 9 1 11 0 9 13 0 7 0 2 3 16 7 1 10 9 9 13 2 0 9 2 2
22 10 3 0 9 13 16 9 13 9 7 9 1 9 15 3 13 9 1 11 0 9 2
22 10 0 4 13 16 10 0 0 9 4 13 7 1 10 0 7 1 10 9 7 9 2
11 10 9 0 7 0 9 4 3 13 0 2
40 15 13 1 10 9 1 9 1 9 1 9 9 2 9 1 9 2 11 0 9 9 1 0 9 2 7 0 7 0 9 1 0 9 1 11 2 9 7 9 2
4 12 0 9 5
12 1 9 12 13 12 0 9 1 10 0 9 2
23 9 13 3 10 9 2 7 13 10 0 0 9 16 15 13 9 1 9 7 11 0 9 2
41 9 13 10 9 9 7 11 0 9 4 13 2 10 9 0 9 4 13 1 9 1 9 7 3 0 9 1 9 11 0 9 4 13 1 9 1 10 9 7 9 2
10 9 1 10 9 1 0 9 13 0 2
14 16 9 9 4 13 2 13 15 10 9 1 0 9 2
21 1 10 9 4 15 3 13 10 9 1 9 7 9 2 3 16 9 4 13 15 2
28 16 15 13 9 1 10 9 1 14 13 9 9 2 4 15 3 0 4 13 1 10 9 2 3 1 9 12 2
12 3 13 15 0 1 0 9 2 9 7 9 2
18 15 13 1 0 3 10 9 1 9 1 0 9 1 14 13 9 9 2
18 10 0 9 1 10 12 9 13 10 0 9 7 9 1 10 0 9 2
16 1 10 0 9 13 1 1 9 11 9 9 1 11 0 9 2
21 1 9 12 13 11 0 9 1 10 0 9 2 7 1 10 10 9 13 1 11 2
22 10 0 9 13 16 9 13 9 1 11 0 9 9 1 0 9 1 10 9 7 9 2
18 9 13 9 7 1 9 1 9 2 11 0 9 7 10 9 7 9 2
13 9 13 3 9 1 0 9 7 9 9 7 9 2
3 0 9 5
12 9 9 13 2 7 0 9 1 9 13 0 2
21 9 13 3 0 9 7 9 1 16 11 2 9 2 13 0 9 7 11 0 9 2
10 9 13 1 15 0 9 1 11 9 2
8 2 13 11 9 12 1 9 2
26 2 13 11 2 9 2 14 13 1 0 9 1 9 16 10 1 10 12 15 4 13 0 9 4 13 2
22 2 13 9 1 9 1 10 0 9 2 3 16 15 3 0 13 1 11 2 9 2 2
15 2 13 9 0 2 0 1 10 9 1 0 9 1 11 2
20 2 13 9 1 1 9 5 9 5 9 7 3 13 10 9 7 9 1 9 2
3 0 9 5
34 9 0 9 1 9 13 7 11 0 9 13 10 0 9 1 10 9 7 1 0 9 1 10 9 15 13 1 9 9 7 9 14 13 2
13 11 9 13 7 9 1 9 1 9 1 9 13 2
16 9 13 1 11 0 9 2 1 9 1 10 0 9 7 9 2
30 11 0 9 13 3 1 9 10 0 9 1 9 1 9 1 10 9 7 9 2 1 10 10 0 9 2 13 1 11 2
8 10 9 4 13 1 10 9 2
26 11 0 9 4 3 13 10 0 9 1 0 9 7 13 9 1 0 9 1 9 7 9 1 10 9 2
18 10 0 9 7 9 1 9 13 3 16 15 4 13 10 9 1 9 2
14 9 13 16 9 1 0 9 3 13 0 9 1 9 2
19 9 13 1 10 9 7 0 9 2 7 9 1 11 0 9 7 9 13 2
16 0 13 13 9 0 9 7 0 9 1 14 13 15 10 9 2
15 9 0 0 9 13 9 15 1 9 13 1 10 0 9 2
19 16 11 9 4 13 2 13 15 0 0 9 1 9 1 3 9 4 13 2
18 9 13 3 10 9 2 13 7 13 10 9 7 9 7 13 10 9 2
3 0 9 5
16 11 0 9 13 1 10 9 7 9 1 11 7 13 0 9 2
19 10 9 1 11 0 9 13 7 10 9 1 0 9 1 9 1 9 13 2
18 11 9 7 9 1 16 9 1 9 4 13 9 1 11 0 9 13 2
13 15 13 3 0 9 1 10 9 1 9 7 9 2
18 11 0 9 13 3 0 10 9 1 9 2 7 13 1 10 0 9 2
18 9 13 10 9 2 9 7 9 1 9 1 9 1 10 9 7 9 2
9 9 13 9 1 11 0 9 9 2
9 9 13 1 10 9 7 0 9 2
18 9 0 0 9 13 9 15 1 9 13 1 10 0 9 1 0 9 2
19 11 0 9 13 10 10 9 15 1 10 9 13 9 1 9 7 0 9 2
22 1 10 9 13 15 1 1 11 0 9 14 13 10 9 15 4 13 1 10 0 9 2
26 9 1 10 0 9 4 13 1 10 3 0 7 0 9 1 0 1 0 2 9 2 0 7 0 9 2
3 12 9 5
16 1 9 12 13 0 9 1 11 0 9 2 0 1 0 9 2
14 9 13 1 0 7 0 9 2 7 9 13 3 0 2
3 0 9 5
14 1 9 13 11 0 9 0 1 9 1 9 7 9 2
42 15 13 0 14 13 10 9 2 16 9 3 7 0 13 9 1 10 9 3 0 9 13 0 0 2 16 9 13 9 1 14 13 9 15 1 0 9 13 1 0 9 2
39 0 4 9 13 1 16 9 13 10 0 9 1 1 9 2 1 10 1 14 13 9 1 9 1 10 0 9 2 7 1 14 13 16 0 9 4 0 13 2
26 10 9 13 14 13 9 1 9 1 10 9 7 0 9 1 9 2 7 13 9 3 13 9 1 9 2
3 0 9 5
20 9 13 1 16 10 9 13 10 0 9 5 9 1 9 7 9 15 9 13 2
12 9 4 7 13 10 0 9 7 0 1 9 2
12 9 4 13 1 1 10 0 9 7 1 9 2
6 10 0 9 13 0 2
26 10 0 9 1 15 15 3 13 9 1 10 9 7 9 2 4 1 9 13 1 10 0 7 0 9 2
2 9 5
11 10 9 1 0 9 4 13 10 10 9 2
12 1 9 1 0 9 13 15 10 0 0 9 2
10 10 9 1 9 4 13 1 0 9 2
36 10 9 13 16 9 13 10 0 0 1 9 1 9 2 7 16 10 9 13 10 0 9 1 0 9 1 0 9 1 9 2 9 2 9 3 2
11 9 4 7 13 1 10 0 7 1 9 2
3 12 9 5
9 1 9 12 13 0 9 1 9 2
20 15 13 0 7 0 9 13 1 9 7 9 1 9 5 9 7 9 2 3 2
18 1 9 1 10 0 7 0 2 13 9 0 0 2 0 7 0 9 2
19 0 9 9 7 10 0 9 1 16 9 13 0 9 2 13 1 9 9 2
18 0 1 15 15 4 13 9 1 9 2 13 9 16 0 9 4 13 2
29 2 15 13 10 0 9 14 13 1 9 7 14 13 9 15 13 16 9 7 9 13 1 0 2 0 7 0 9 2
14 2 15 4 13 1 9 7 9 1 0 9 7 9 2
21 2 9 13 3 0 15 13 0 13 1 9 1 10 9 10 0 9 7 9 13 2
28 2 10 0 4 0 13 9 1 14 13 1 9 0 0 9 1 9 1 9 15 3 13 0 9 1 10 9 2
24 0 1 9 2 13 15 1 9 9 12 0 9 14 13 9 1 9 2 1 0 9 7 9 2
9 9 13 9 7 9 1 10 9 2
6 12 0 7 0 9 5
9 1 9 12 13 0 7 0 9 2
15 9 0 9 7 9 13 10 0 9 1 9 1 0 9 2
8 9 9 13 1 9 0 9 2
21 10 0 7 0 9 7 9 13 10 0 9 13 10 0 9 1 14 13 10 9 2
15 9 1 9 7 9 9 4 13 1 9 7 9 7 9 2
14 9 2 9 2 9 7 9 1 9 4 13 1 9 2
10 16 10 9 13 2 13 9 0 9 2
27 16 9 13 0 7 0 2 13 15 10 0 9 2 1 9 4 11 3 13 9 1 9 1 9 1 9 2
12 9 1 0 9 13 9 7 1 9 7 9 2
13 10 9 1 10 9 4 13 1 7 11 7 9 2
8 9 13 1 9 13 1 11 2
18 11 13 3 12 9 2 1 15 13 12 0 7 12 13 9 1 0 2
8 15 13 0 0 7 0 9 2
15 9 1 11 13 16 10 0 9 1 9 4 3 0 13 2
26 1 1 11 9 13 15 1 9 12 9 9 3 0 1 9 2 7 3 12 9 9 13 1 0 9 2
3 12 9 5
12 1 9 12 13 9 1 9 2 9 7 9 2
41 10 0 0 9 4 3 13 1 10 9 2 7 4 1 9 13 1 16 9 1 9 4 4 13 10 9 1 10 9 2 1 0 9 1 9 2 9 2 9 3 2
14 10 0 0 0 9 4 13 1 11 9 2 11 2 2
26 3 4 10 0 0 9 0 13 1 11 2 9 7 0 9 15 13 9 1 9 7 9 1 10 9 2
13 15 13 3 3 10 0 9 1 9 1 10 9 2
30 1 9 13 15 10 0 0 9 2 9 3 2 2 15 3 4 13 1 9 2 7 15 0 4 4 13 1 9 9 2
18 16 9 13 3 16 11 0 9 13 10 10 9 2 4 15 13 9 2
19 3 4 15 13 10 9 7 9 11 0 9 13 7 4 4 13 1 9 2
6 12 9 9 7 9 5
24 1 9 12 13 9 9 7 0 9 1 0 9 2 9 2 9 2 0 7 0 9 7 9 2
8 9 9 13 1 9 1 9 2
7 12 9 1 9 7 9 5
14 9 12 13 10 0 9 1 9 9 1 9 7 9 2
3 12 9 5
13 1 9 12 4 0 7 0 9 1 9 9 13 2
6 12 0 9 1 11 5
3 12 9 5
3 12 0 5
22 10 0 9 13 10 0 9 1 16 9 1 11 1 9 13 15 0 1 10 0 9 2
15 10 0 9 13 0 9 7 9 15 13 1 9 1 9 2
19 9 2 9 7 10 9 15 3 4 13 1 0 9 2 13 9 1 9 2
25 0 9 2 0 9 7 0 9 13 16 10 0 9 1 9 13 0 2 7 0 1 10 0 9 2
30 10 0 9 1 11 13 10 9 1 15 0 9 4 13 2 7 15 13 3 0 9 15 4 13 14 13 15 10 9 2
18 9 13 1 1 10 0 9 0 0 7 9 13 0 13 1 0 9 2
12 1 9 13 15 0 0 9 1 10 0 9 2
18 10 0 9 1 7 1 11 13 0 0 1 10 0 0 9 1 11 2
29 9 1 1 0 9 1 11 9 13 1 10 0 9 7 10 0 0 9 1 11 1 1 0 9 10 9 1 11 2
20 7 10 0 9 7 9 1 9 7 9 13 1 9 10 9 1 10 0 9 2
20 1 0 9 13 15 3 9 7 9 15 13 9 1 9 1 9 1 12 9 2
9 10 0 9 13 3 9 1 9 2
18 15 13 10 12 9 2 9 7 10 10 9 15 0 13 1 1 11 2
13 11 4 1 10 0 1 10 0 9 13 1 9 2
24 3 1 9 4 15 13 9 1 9 2 9 2 9 2 9 3 15 0 4 13 1 0 9 2
30 10 1 0 9 13 16 15 1 11 13 9 1 10 9 1 9 9 2 7 0 13 0 0 9 1 9 9 7 9 2
14 13 1 10 0 9 13 11 9 0 13 1 0 9 2
36 1 10 9 9 13 9 0 13 0 1 0 0 9 2 10 0 0 9 13 0 13 0 2 7 10 0 9 4 13 1 0 0 9 7 9 2
3 12 9 5
11 9 13 1 9 11 0 7 0 0 9 2
15 10 0 9 1 11 13 3 0 0 13 1 10 0 11 2
19 0 1 9 15 13 3 2 13 0 1 0 9 2 7 13 3 0 1 2
22 0 1 9 1 11 13 3 10 9 2 15 13 15 1 9 1 10 9 3 1 11 2
13 1 9 13 9 10 10 9 15 3 13 10 9 2
19 0 9 13 3 0 9 1 9 15 4 13 1 7 13 0 1 0 9 2
26 10 9 1 11 13 9 2 9 2 2 15 13 0 9 1 11 2 7 15 13 10 0 9 1 11 2
40 9 1 10 0 0 9 7 0 9 15 0 13 0 0 2 7 0 9 2 0 9 7 9 1 0 9 1 11 13 11 0 0 0 1 9 1 9 7 9 2
56 0 9 16 10 0 0 9 1 9 2 9 2 7 9 13 0 7 13 15 0 0 1 0 9 2 9 7 9 2 13 0 7 1 9 1 0 0 9 2 7 16 10 9 13 0 9 1 14 13 9 1 0 7 0 9 2
25 9 1 0 9 13 0 1 16 0 9 13 0 0 7 3 0 0 1 9 1 9 1 0 9 2
16 9 13 3 1 0 9 7 13 9 1 9 7 9 1 9 2
31 15 13 0 14 13 16 9 1 9 7 0 9 4 13 1 9 16 9 1 10 9 13 1 0 9 2 0 3 1 0 2
13 9 1 0 9 9 13 1 14 13 11 9 0 2
16 15 13 1 10 0 15 13 9 1 11 9 2 13 9 12 2
20 15 7 13 7 13 10 0 9 7 9 2 7 13 1 10 0 9 1 9 2
3 12 9 5
22 9 1 11 13 0 10 0 9 7 10 0 9 1 9 2 9 7 9 15 13 9 2
20 10 0 9 13 3 0 7 13 0 9 1 9 1 9 2 9 7 0 9 2
22 0 9 1 10 0 9 7 9 9 1 10 9 13 3 10 0 9 0 1 0 9 2
13 0 9 7 0 9 13 16 9 7 9 13 0 2
14 7 9 7 0 0 9 13 3 0 0 1 1 11 2
20 9 1 11 13 0 16 0 9 13 1 0 9 16 15 4 13 9 1 9 2
13 9 13 3 1 16 9 1 0 9 13 0 0 2
14 9 1 9 13 10 0 9 2 9 13 2 7 13 2
8 15 13 16 0 9 13 0 2
26 0 9 13 3 1 9 1 9 7 1 0 9 2 7 0 1 12 9 1 9 13 0 9 1 9 2
25 16 0 9 3 13 0 1 10 0 9 13 9 7 9 10 0 0 9 1 10 0 0 0 9 2
22 10 0 9 1 9 1 11 13 3 0 9 2 7 0 13 3 0 1 10 0 9 2
29 9 7 9 1 10 9 4 3 13 9 1 10 9 1 11 2 7 1 0 9 13 1 16 10 9 13 1 9 2
32 7 1 9 7 1 9 13 10 0 9 1 9 0 1 0 0 9 2 0 1 9 7 9 1 10 0 9 1 9 7 9 2
14 9 1 15 13 9 2 9 1 9 7 9 1 9 2
29 10 0 9 1 0 9 13 16 9 2 0 9 7 9 15 13 0 0 9 4 13 0 9 1 0 9 7 9 2
18 10 0 9 1 10 0 0 9 13 9 1 9 1 9 0 1 9 2
22 16 9 1 10 9 4 0 13 2 4 15 13 0 9 1 10 9 0 1 1 9 2
15 10 0 0 9 1 9 7 9 13 0 7 13 0 9 2
12 9 13 3 0 0 9 7 10 9 1 9 2
21 1 9 13 15 0 0 1 0 9 1 9 1 1 9 9 1 9 7 0 9 2
28 16 9 1 10 0 9 1 11 13 0 1 10 0 9 1 11 2 13 9 1 9 7 9 1 10 9 0 2
33 15 13 3 1 10 0 9 3 0 9 1 9 7 9 2 16 10 0 9 13 1 14 13 9 1 10 0 9 1 9 1 11 2
20 10 0 9 1 0 9 13 11 9 0 1 0 9 1 9 9 7 1 9 2
26 10 9 13 10 0 9 1 9 1 9 2 15 13 9 1 9 1 9 9 7 9 1 11 7 11 2
9 9 13 0 0 0 13 1 9 2
34 9 1 9 7 0 10 0 9 13 3 0 1 9 15 13 15 1 9 1 10 0 9 1 11 2 1 1 10 0 10 9 1 11 2
25 15 13 0 1 9 9 1 9 1 9 7 9 1 1 2 7 9 1 0 9 4 3 3 13 2
30 0 1 10 0 9 13 0 7 0 0 2 7 0 0 9 13 0 9 1 9 1 0 1 9 1 0 9 1 9 2
14 0 9 13 1 10 9 7 13 1 9 3 1 9 2
20 1 10 9 13 0 9 1 9 3 16 9 1 9 13 0 9 1 10 9 2
11 0 0 9 4 1 10 13 9 7 9 2
5 12 9 7 9 5
12 1 1 10 0 9 1 12 13 11 0 9 2
16 1 9 4 3 9 1 0 9 13 9 1 10 9 1 9 2
8 15 4 13 1 10 0 9 2
12 9 9 1 11 13 15 1 10 12 9 9 2
5 15 13 10 9 2
20 9 4 3 13 0 1 0 9 15 3 4 13 9 1 9 1 10 0 9 2
16 11 4 0 13 13 10 0 9 1 15 15 4 13 15 3 2
12 9 4 4 13 1 9 1 0 7 0 9 2
38 16 10 0 1 9 0 4 13 1 9 2 7 13 0 9 1 9 2 4 11 1 9 1 10 0 12 9 13 1 10 9 1 9 2 9 7 9 2
15 1 11 13 9 1 0 9 2 7 1 0 9 1 9 2
22 16 11 0 13 10 9 1 9 7 9 2 13 15 3 3 0 1 10 9 3 3 2
26 16 9 13 1 11 1 12 7 1 1 3 12 2 13 15 9 1 10 0 9 15 13 9 1 9 2
16 9 4 0 13 2 7 0 9 4 0 13 1 9 1 11 2
13 1 1 12 13 9 1 9 2 3 7 0 9 2
10 1 10 0 9 13 9 1 0 9 2
10 10 0 9 13 1 9 12 2 12 2
34 9 1 11 9 1 9 13 1 11 9 7 9 1 11 2 9 0 9 1 11 7 9 1 10 0 9 1 9 1 9 1 0 9 2
20 1 9 1 9 13 15 3 11 7 11 2 3 11 15 13 10 9 1 11 2
26 1 9 1 9 1 9 1 9 13 11 9 1 9 2 16 7 11 2 11 7 0 10 9 13 0 2
24 10 9 9 4 13 1 14 13 9 2 7 1 12 4 1 9 1 11 13 1 9 7 9 2
14 1 12 13 10 9 9 10 0 9 1 10 0 9 2
15 10 0 9 1 11 4 13 9 1 10 9 1 1 9 2
26 1 9 4 9 1 0 9 9 3 13 1 0 9 1 9 2 16 1 11 4 9 13 3 7 0 2
15 3 10 9 15 13 0 1 14 13 1 9 4 4 13 2
17 15 13 0 9 1 9 2 7 0 1 10 0 9 4 0 13 2
28 9 1 9 2 9 7 9 13 3 0 1 9 1 9 7 9 2 7 0 4 13 7 13 1 3 10 9 2
16 0 1 0 9 1 9 13 9 15 13 15 1 9 7 1 2
17 9 13 1 0 9 1 9 2 16 0 9 7 9 13 1 9 2
21 9 13 0 1 9 1 9 7 9 1 9 1 9 1 10 0 9 1 10 9 2
11 15 13 0 1 9 1 9 1 10 9 2
13 9 1 0 9 13 3 0 14 13 1 10 9 2
21 9 4 13 1 10 9 7 0 9 2 15 13 15 0 1 9 14 13 0 9 2
36 9 1 9 13 0 1 10 9 15 13 10 0 0 9 2 3 1 11 9 7 0 1 10 0 9 11 2 11 2 11 2 11 7 1 11 2
13 15 13 3 0 9 7 0 9 1 9 1 11 2
16 10 0 9 1 11 13 0 1 10 0 9 1 9 7 9 2
29 0 13 0 0 9 2 9 2 9 2 9 2 9 2 1 0 7 0 9 2 7 1 10 9 13 10 9 9 2
16 1 9 7 9 13 15 9 1 9 1 9 7 0 0 9 2
25 15 4 4 13 10 9 9 1 9 1 0 9 7 9 2 7 15 13 9 1 9 1 10 9 2
45 16 0 1 9 1 11 13 1 9 2 13 15 9 1 14 13 16 15 13 9 1 9 1 9 2 7 0 9 2 9 2 9 3 2 2 9 1 0 9 7 9 1 0 9 2
9 15 13 3 0 9 1 0 9 2
20 9 1 9 4 13 0 2 7 7 9 9 7 9 13 0 1 9 1 9 2
5 12 9 1 11 5
16 15 13 12 9 1 10 0 9 1 11 2 7 15 13 1 2
24 1 9 13 15 9 1 0 9 1 1 1 9 2 1 10 1 11 2 1 11 7 1 11 2
3 12 11 5
11 11 13 11 0 9 2 7 13 1 11 2
16 11 13 9 1 11 2 7 9 7 0 9 13 10 9 3 2
14 9 13 1 1 9 1 9 1 9 1 10 12 9 2
19 1 12 13 11 11 11 11 11 9 1 11 1 10 0 9 11 11 11 2
27 1 16 9 12 4 13 1 12 2 13 15 3 3 1 11 12 0 1 11 9 13 9 1 9 1 11 2
8 1 9 13 9 9 1 11 2
23 0 9 1 10 0 9 1 11 2 11 12 7 11 2 13 1 3 12 12 9 1 9 2
32 10 0 12 12 9 4 15 13 1 10 0 9 1 9 1 9 2 9 7 9 2 7 3 1 10 0 9 1 10 0 9 2
17 15 13 1 9 3 12 9 1 11 2 3 3 12 13 0 9 2
16 10 0 9 9 1 0 9 4 3 13 9 1 9 13 9 2
11 15 13 3 10 0 9 1 9 7 9 2
15 11 1 11 2 11 2 13 0 3 12 9 1 0 9 2
32 10 0 9 1 11 1 10 9 13 10 0 1 9 1 0 9 1 9 2 7 15 4 13 1 9 16 9 13 3 12 9 2
13 11 13 1 9 1 10 0 9 1 0 0 9 2
39 1 10 0 9 4 15 13 9 15 4 13 0 9 1 9 2 0 4 13 9 1 9 1 11 1 9 1 9 1 11 11 7 10 0 9 1 9 11 2
3 12 11 5
11 11 13 9 0 0 9 2 0 1 11 2
14 1 11 9 1 12 4 15 3 4 13 9 1 9 2
16 11 4 13 16 11 4 13 9 1 0 7 0 9 1 11 2
18 1 9 13 3 12 9 1 9 7 9 1 9 1 1 9 12 9 2
14 11 11 11 13 9 7 13 10 0 1 9 1 9 2
15 9 13 10 0 9 1 9 7 13 9 2 9 7 9 2
10 1 9 12 9 13 1 11 9 1 2
17 1 9 1 9 13 1 12 9 1 9 2 10 0 13 1 9 2
27 9 13 0 1 9 0 1 9 15 15 4 13 9 1 9 7 9 9 1 0 0 9 1 9 1 9 2
3 12 11 5
18 11 2 15 13 1 11 2 13 1 9 10 12 0 0 9 1 11 2
16 1 9 13 15 9 1 10 9 1 9 1 9 3 1 9 2
21 11 13 3 12 9 2 0 0 1 1 3 12 9 3 2 16 9 13 3 12 2
18 9 13 1 11 7 11 7 13 12 9 9 1 10 0 9 11 11 2
23 10 0 9 2 11 11 2 13 10 9 9 1 9 1 0 9 1 9 1 10 0 9 2
17 1 12 13 11 10 9 2 7 1 0 9 4 9 13 1 9 2
15 9 1 11 4 10 0 12 9 4 13 1 12 0 9 2
31 1 9 12 13 12 9 1 9 1 11 1 9 1 11 1 11 2 7 1 9 12 4 12 9 13 1 10 9 1 9 2
3 12 11 5
18 11 13 1 11 2 7 13 1 12 10 0 9 1 0 9 1 11 2
15 11 11 13 1 9 12 9 1 11 1 12 9 0 9 2
23 1 10 0 13 3 12 9 7 9 1 11 2 7 9 13 9 2 9 7 10 0 9 2
22 9 12 5 12 4 11 13 0 2 7 15 13 0 10 9 11 11 13 1 9 9 2
9 9 1 9 1 9 4 4 13 2
24 9 7 9 1 11 13 0 0 9 2 7 9 4 13 1 16 9 4 13 0 0 1 9 2
19 9 4 0 13 9 1 16 15 4 13 1 1 0 9 7 9 1 9 2
24 9 1 11 4 13 0 1 9 2 7 15 4 13 10 3 0 9 1 11 11 1 9 9 2
3 12 11 5
30 11 11 11 11 11 2 11 2 4 13 9 1 11 1 11 11 1 12 2 16 9 4 13 1 9 11 11 11 11 2
10 11 11 13 9 10 0 9 1 9 2
22 3 1 12 13 9 14 13 9 0 0 2 7 0 1 12 13 11 11 0 9 3 2
18 9 1 11 13 1 9 0 0 1 11 15 13 1 11 1 10 9 2
14 15 13 15 1 10 9 1 12 7 12 9 1 11 2
18 11 11 4 13 1 9 1 9 1 10 0 9 1 1 11 2 11 2
29 16 15 13 9 1 9 1 10 9 2 13 9 1 14 4 13 1 12 7 12 9 9 1 9 1 12 9 1 2
19 16 11 3 4 13 2 4 9 13 1 1 9 1 9 3 0 1 0 2
13 12 9 1 9 1 11 2 1 0 9 1 9 5
5 12 11 7 9 5
24 11 13 9 1 11 1 10 0 9 2 11 2 2 13 9 9 12 9 12 7 12 9 12 2
7 11 9 4 13 1 11 2
6 0 13 9 1 11 2
2 11 5
2 11 5
2 11 5
4 11 7 9 5
2 11 5
2 11 5
3 11 11 5
22 9 1 10 9 13 16 9 13 10 9 15 13 1 10 9 15 3 13 0 1 9 2
22 1 9 4 11 13 9 1 16 10 9 1 11 11 4 13 1 9 1 9 1 11 2
34 10 9 13 9 1 16 9 13 9 1 9 1 9 2 13 9 1 11 1 12 9 12 9 12 7 9 13 1 9 9 12 9 12 2
11 3 13 9 1 11 1 0 9 1 9 2
35 11 13 10 0 9 1 9 1 11 1 11 1 9 2 11 9 2 11 11 2 11 2 11 9 1 0 9 7 11 1 11 1 0 9 2
20 0 10 9 13 1 10 9 10 0 9 1 9 15 13 9 1 9 1 11 2
65 15 13 0 11 15 13 9 1 11 7 13 9 1 9 2 11 2 9 7 9 15 13 10 9 1 9 1 9 7 9 2 11 7 9 15 13 9 9 1 9 7 9 1 0 9 2 13 0 0 9 2 7 11 15 13 9 1 9 1 9 7 9 1 11 2
12 11 13 9 1 10 0 9 0 9 1 11 2
20 10 0 0 9 2 0 0 9 7 0 9 13 1 9 9 9 12 10 9 2
12 1 9 7 9 13 9 1 0 9 7 9 2
3 12 9 5
3 12 9 5
18 1 12 4 9 1 10 0 9 1 11 13 1 11 2 11 7 9 2
22 11 9 2 11 2 13 9 1 9 2 16 11 1 9 2 11 2 3 4 13 9 2
13 9 13 16 11 13 9 15 1 9 13 0 9 2
42 1 14 13 10 0 9 7 9 7 0 13 10 0 9 1 9 1 11 13 11 1 9 9 9 12 2 12 2 12 2 11 9 1 11 1 1 14 13 9 0 9 2
19 15 4 13 1 1 9 12 2 16 11 13 9 7 9 1 11 7 11 2
26 1 9 1 0 9 1 11 13 0 9 13 10 9 3 9 1 0 9 15 13 9 1 9 7 9 2
15 15 13 0 11 2 11 2 11 2 11 7 11 1 11 2
42 1 9 13 10 0 9 9 9 1 9 1 10 0 9 2 13 1 1 10 9 2 2 0 9 2 9 2 9 1 9 1 9 13 1 9 7 9 1 9 1 9 2
15 9 4 13 9 1 14 13 9 1 0 9 1 10 9 2
12 9 9 1 10 9 1 9 1 11 13 3 2
5 12 11 1 9 5
29 11 1 9 13 9 1 10 9 1 11 2 1 0 9 7 9 2 3 9 7 9 1 9 1 9 13 1 9 2
34 11 1 9 13 1 9 9 1 14 13 0 9 7 9 1 0 9 7 9 1 9 1 9 1 9 1 0 9 7 9 2 11 2 2
43 11 1 9 13 3 9 1 9 2 3 14 13 9 1 0 0 9 1 9 2 7 13 9 2 14 13 9 1 0 9 15 9 13 7 14 13 9 1 9 13 1 9 2
6 9 13 0 9 1 2
16 9 1 9 2 3 9 7 9 1 9 1 9 13 1 9 2
8 9 1 9 1 9 7 9 2
13 9 1 9 7 0 10 9 13 1 9 1 11 2
4 12 11 9 5
27 11 9 7 9 13 0 0 1 9 1 0 9 2 9 1 9 2 9 1 0 9 7 9 1 0 9 2
9 11 13 7 13 9 1 10 9 2
15 0 4 15 13 9 15 13 9 2 7 11 13 3 9 2
14 1 9 1 0 0 9 4 15 13 11 15 13 9 2
10 11 13 3 9 1 9 1 0 9 2
3 12 11 5
8 11 13 9 1 9 0 9 2
17 11 13 0 9 1 10 10 0 9 1 9 15 13 9 1 11 2
19 9 1 9 7 9 1 9 1 10 9 9 13 0 9 4 13 1 11 2
4 12 11 11 5
14 11 11 13 10 0 0 7 0 9 1 9 1 11 2
21 9 13 9 1 0 7 0 9 2 9 1 9 7 0 9 1 0 7 0 9 2
16 10 0 9 1 9 13 3 14 13 0 9 1 9 7 9 2
3 12 11 5
12 9 1 9 7 9 1 11 13 1 11 9 2
30 11 13 9 1 9 1 9 1 11 9 7 1 9 2 1 9 1 9 13 1 9 9 12 9 12 1 9 1 9 2
15 0 13 9 11 1 9 1 9 1 9 1 9 1 9 2
3 12 11 5
44 11 13 9 1 16 9 15 13 1 9 13 9 15 4 13 1 14 13 9 1 10 0 9 1 10 9 9 12 9 12 9 12 12 1 11 1 11 11 9 12 13 1 11 2
22 15 13 10 9 1 9 1 11 2 7 9 1 11 13 9 1 9 1 9 1 9 2
3 12 11 5
35 9 1 9 1 9 15 13 1 9 12 9 12 9 12 1 9 2 9 2 7 9 2 13 1 11 2 1 9 1 9 1 9 7 9 2
18 9 15 13 9 1 9 2 13 0 9 1 9 1 9 2 9 3 2
4 12 0 9 5
5 12 11 1 11 5
17 11 13 9 0 9 1 11 7 4 13 10 0 9 9 1 9 2
17 10 9 9 15 1 9 4 13 1 0 9 2 4 13 1 9 2
20 15 13 10 9 1 10 9 2 7 13 3 9 2 3 9 1 10 0 9 2
33 11 13 9 1 10 0 0 9 1 11 1 9 1 10 0 9 2 3 9 1 9 7 9 1 9 15 13 0 1 9 7 11 2
25 11 13 10 0 9 1 10 0 9 1 0 9 1 11 2 1 9 2 12 0 9 1 9 2 2
17 1 9 13 11 9 2 7 9 13 9 16 11 13 9 1 9 2
30 1 9 9 9 12 2 12 2 12 2 13 11 1 1 14 13 10 10 9 1 9 2 3 15 13 1 9 1 9 2
26 9 4 13 12 9 12 2 7 13 3 10 0 9 1 12 0 9 10 9 2 12 9 7 12 9 2
17 1 9 1 10 9 15 13 2 13 9 1 9 2 9 7 9 2
18 1 9 1 9 13 15 10 9 16 9 1 9 7 9 13 0 3 2
10 1 9 13 9 1 3 9 7 9 2
23 1 9 13 9 9 15 13 9 7 9 7 0 13 9 9 1 9 1 7 1 1 11 2
12 9 13 1 9 0 1 10 9 7 10 9 2
18 11 13 0 9 1 9 7 9 2 0 1 9 14 13 7 13 9 2
5 12 11 1 11 5
21 11 1 11 13 10 0 9 1 9 1 9 1 11 13 1 9 9 12 9 12 2
23 11 13 9 2 9 2 2 15 13 9 1 9 1 10 10 0 9 15 13 1 9 9 2
18 1 9 1 0 9 7 9 1 9 7 9 13 9 0 9 1 9 2
9 15 13 1 0 9 1 9 9 2
20 11 1 11 13 9 1 10 0 7 0 9 16 15 13 9 1 10 0 9 2
16 1 10 9 13 9 1 9 1 9 15 4 13 9 1 9 2
19 11 4 0 13 1 16 11 0 9 13 7 13 0 0 1 9 1 9 2
25 1 10 9 4 9 13 14 13 9 7 9 1 9 1 10 1 9 7 9 1 11 1 10 9 2
6 9 1 9 1 11 5
15 12 11 11 11 7 11 11 4 3 13 1 9 7 9 2
31 10 9 9 15 13 1 9 1 9 4 1 11 13 11 11 11 2 11 2 2 15 13 10 0 0 9 13 11 7 9 2
32 15 13 1 10 9 1 9 2 9 2 9 7 9 7 10 9 0 9 1 9 1 9 7 9 7 0 9 1 9 7 9 2
33 10 0 9 11 2 12 9 2 13 1 1 9 3 7 0 0 9 2 7 4 13 0 9 2 9 1 9 1 9 7 9 2 2
18 15 13 3 0 9 1 16 11 4 13 9 1 14 13 9 1 11 2
24 10 0 0 9 1 11 1 10 0 9 1 10 0 9 4 4 13 1 10 0 9 1 11 2
4 12 11 11 5
7 12 11 11 9 7 9 5
26 11 11 13 10 12 9 0 9 15 13 1 1 11 2 12 9 1 1 11 7 12 9 1 1 11 2
11 9 13 3 12 9 1 7 9 7 11 2
20 15 13 15 12 9 1 1 9 1 9 1 5 7 5 7 1 5 7 5 2
19 9 13 1 12 9 2 10 0 11 7 11 2 1 10 0 2 0 9 2
24 1 12 13 11 11 10 9 1 11 11 2 13 9 12 9 12 9 12 1 11 11 9 12 2
32 10 0 9 13 3 10 10 1 11 11 7 11 2 1 9 1 10 0 9 15 4 13 1 9 1 9 12 9 12 9 12 2
24 11 13 3 1 11 11 2 3 16 0 9 4 13 1 11 11 1 9 1 9 15 9 13 2
34 16 11 11 13 10 9 1 9 2 13 16 9 15 11 13 0 1 2 3 13 1 9 1 11 11 16 15 3 4 13 9 1 9 2
5 12 9 7 9 5
6 12 9 1 11 11 5
18 11 11 4 13 1 0 9 2 7 9 13 0 1 0 9 1 11 2
21 10 0 9 11 2 12 9 2 1 11 13 3 0 7 13 10 0 9 1 12 2
14 3 13 15 9 7 1 9 7 0 10 9 1 9 2
22 9 13 1 9 1 0 7 0 9 1 10 0 9 1 11 15 13 1 5 7 5 2
12 9 13 1 10 9 15 0 13 0 9 1 2
16 9 13 1 10 0 9 2 7 13 1 1 12 9 1 11 2
29 0 1 0 9 3 1 9 4 11 11 13 1 3 0 9 16 10 0 9 1 9 13 0 0 1 10 0 9 2
27 9 13 3 0 1 0 9 2 13 13 9 0 9 2 1 9 1 9 2 0 9 7 0 9 1 9 2
9 0 9 1 9 13 0 1 9 2
13 9 9 7 9 1 10 9 13 16 9 13 0 2
13 9 7 9 13 0 1 9 1 0 7 0 9 2
21 13 1 11 4 11 11 13 0 9 2 7 1 9 13 9 15 13 10 0 9 2
10 9 13 1 0 9 2 9 7 9 2
10 15 13 3 9 7 9 1 11 11 2
5 0 9 13 0 2
5 9 13 3 0 2
4 9 13 3 2
9 15 13 10 0 0 9 1 9 2
12 9 13 3 1 10 0 0 1 9 7 9 2
12 9 13 0 16 9 13 1 1 11 11 3 2
13 9 13 12 0 9 7 13 15 3 0 1 11 2
13 9 4 3 13 9 7 9 1 0 9 1 9 2
4 9 13 3 2
15 11 1 11 13 10 12 9 15 3 13 1 1 0 9 2
21 10 13 1 10 9 1 9 15 15 13 4 13 0 1 9 1 12 7 12 9 2
4 9 13 0 2
18 11 9 13 10 0 9 1 0 9 2 7 10 9 9 13 1 9 2
17 15 4 13 7 13 10 0 9 1 0 9 1 9 1 11 11 2
13 0 11 11 13 15 3 0 9 1 9 7 9 2
16 1 9 13 15 0 9 1 9 7 9 15 4 4 0 13 2
6 9 4 3 4 13 2
16 1 0 4 15 13 10 0 9 1 9 2 9 7 0 9 2
18 9 1 0 9 4 3 13 1 9 1 10 9 15 13 1 11 9 2
23 15 4 13 0 9 0 1 0 9 2 7 0 16 15 4 4 13 9 1 0 9 0 2
6 0 9 13 0 9 2
12 9 7 9 1 9 13 10 0 9 1 9 2
11 15 13 0 9 2 3 15 13 0 9 2
6 12 9 1 0 9 5
30 10 0 0 9 1 9 1 11 11 13 15 1 9 2 7 15 13 9 1 14 13 1 16 11 11 13 0 1 9 2
19 9 4 2 9 2 13 1 12 1 9 7 9 1 9 1 9 1 9 2
20 9 13 10 9 1 10 0 9 2 7 9 13 0 9 1 11 11 1 9 2
11 15 13 3 0 9 1 9 7 10 9 2
23 1 15 13 9 1 10 9 16 10 0 0 9 13 0 1 10 9 3 1 12 2 12 2
14 0 1 9 13 9 1 9 2 3 7 0 1 9 2
11 0 9 13 16 10 9 13 9 1 9 2
17 15 13 9 1 10 0 9 7 0 9 1 9 2 1 10 9 2
9 10 0 0 9 4 13 1 12 2
11 1 15 13 15 3 9 7 0 9 3 2
17 1 9 1 9 12 2 12 4 15 13 0 0 9 1 11 11 2
34 1 10 9 4 9 1 11 11 13 1 11 2 7 9 1 10 0 9 1 9 1 0 1 9 1 11 13 16 9 4 13 1 3 2
22 1 9 13 3 11 11 10 12 9 1 11 15 0 1 13 1 10 0 0 9 9 2
10 1 9 4 15 13 10 0 0 9 2
12 15 4 13 1 12 7 13 3 10 0 9 2
20 1 9 1 10 9 4 9 3 13 9 1 7 0 13 10 0 9 7 9 2
5 12 9 1 9 5
14 9 1 11 11 1 9 13 1 0 0 7 0 9 2
13 15 13 15 1 0 9 7 1 12 1 9 11 2
17 10 0 9 1 11 11 13 1 0 9 2 7 13 3 1 11 2
13 1 9 13 15 0 12 9 15 13 1 11 11 2
15 9 1 9 13 1 9 1 9 2 7 3 13 3 9 2
4 9 13 0 2
23 9 13 1 1 9 7 13 3 3 2 3 1 9 2 7 13 1 9 1 10 0 9 2
8 9 1 11 11 13 3 0 2
15 1 12 13 10 9 15 10 0 9 4 13 1 9 1 2
26 15 13 0 7 13 1 11 15 13 15 1 11 10 10 7 0 9 1 14 13 1 9 7 0 9 2
6 9 13 10 0 9 2
16 9 1 9 4 13 0 2 7 13 0 7 1 9 7 9 2
19 15 13 9 1 10 0 9 7 9 1 11 2 13 1 10 0 0 9 2
10 15 13 3 0 9 1 9 1 9 2
16 9 1 11 11 13 3 1 10 0 0 1 10 0 5 9 2
8 1 9 13 15 10 0 9 2
27 1 0 9 0 9 4 9 13 3 0 16 15 4 13 0 14 13 15 1 14 13 16 9 4 4 13 2
25 15 13 10 0 9 1 9 7 10 0 2 7 15 4 3 13 1 1 10 9 1 9 7 9 2
16 3 4 3 0 9 13 15 1 9 1 9 16 9 13 15 2
6 12 9 1 11 11 5
4 12 0 9 5
17 1 11 9 9 12 13 0 9 7 9 7 0 9 1 11 11 2
14 10 9 13 1 11 11 3 1 10 9 15 4 13 2
24 15 13 0 1 11 9 3 2 9 12 0 9 10 9 2 2 7 4 3 13 1 0 9 2
28 12 10 0 9 1 11 13 1 10 9 0 9 1 9 2 11 11 2 2 13 11 9 1 11 12 9 12 2
28 16 9 13 10 9 1 9 1 12 2 13 10 9 2 9 2 9 7 9 9 2 13 3 11 9 9 12 2
12 10 9 13 3 16 15 4 13 9 1 9 2
7 11 11 13 10 10 9 2
22 1 9 1 9 13 10 0 9 2 15 13 15 1 9 13 1 9 9 12 9 12 2
29 1 1 15 13 9 12 9 12 9 12 1 11 0 9 9 1 14 13 10 0 9 1 1 12 0 9 1 9 2
29 1 9 13 1 9 9 12 9 12 4 10 9 13 1 14 13 10 12 9 9 2 3 10 0 9 13 1 9 2
30 12 1 9 1 11 4 10 9 13 1 10 0 12 9 9 2 9 1 11 7 11 12 9 12 7 12 9 12 2 2
29 1 11 4 9 13 1 1 11 0 9 9 1 11 9 1 11 7 11 1 12 2 11 11 12 9 12 0 2 2
6 12 9 9 1 9 5
32 9 1 9 1 11 12 1 0 12 9 3 2 11 11 2 12 2 2 4 1 10 0 11 9 13 1 10 9 1 12 9 2
31 9 13 16 9 1 11 11 2 12 2 1 11 7 11 11 2 12 2 1 11 4 13 1 0 9 7 1 3 0 9 2
13 1 9 13 15 16 0 4 13 12 9 1 9 2
10 1 15 4 15 13 12 9 1 9 2
12 9 1 9 1 12 9 4 3 13 1 9 2
22 0 13 9 7 13 12 9 1 15 1 14 13 16 15 4 13 9 1 1 11 9 2
3 0 9 5
37 9 4 3 13 16 3 13 9 1 16 2 9 2 4 4 13 0 9 1 10 9 7 1 10 10 9 16 15 4 4 13 1 1 9 1 9 2
42 3 4 0 1 10 12 9 13 1 0 0 2 0 7 1 0 9 2 7 9 13 3 3 3 1 9 1 16 2 9 2 0 9 1 9 3 4 13 1 0 9 2
4 0 14 13 5
35 2 15 4 13 0 14 13 9 1 9 2 13 9 2 9 11 11 11 1 11 2 7 15 13 3 10 0 9 14 13 15 0 1 3 2
12 15 13 15 13 0 1 9 3 14 13 9 2
4 13 1 9 5
27 1 1 0 9 1 10 9 2 13 15 3 14 13 10 9 7 13 10 9 1 0 3 1 9 7 0 2
28 0 13 3 16 9 1 15 13 3 0 7 0 2 1 10 9 1 16 11 13 1 1 11 1 9 1 9 2
32 1 15 13 15 16 15 0 9 4 13 1 7 3 9 13 15 2 13 15 15 10 9 1 16 15 4 13 15 10 10 9 2
14 15 13 0 10 9 1 16 10 9 4 13 11 11 2
3 0 9 5
31 9 13 1 9 16 0 1 9 1 10 0 12 9 16 9 13 9 2 4 13 10 0 9 1 16 11 3 0 13 15 2
22 10 0 9 13 10 0 9 1 15 2 7 9 13 1 9 16 9 13 1 1 9 2
3 13 9 5
11 0 13 1 9 7 13 15 1 12 9 2
9 3 13 15 1 11 12 1 9 2
24 1 11 12 13 15 1 9 7 13 10 9 1 9 7 9 3 16 9 3 4 13 1 9 2
19 3 13 15 1 1 10 10 9 2 13 15 1 9 7 13 14 13 9 2
12 9 15 4 13 1 2 9 2 13 15 0 2
11 15 13 1 9 7 13 1 1 11 12 2
20 16 15 13 15 1 14 4 13 13 9 1 1 15 2 13 3 9 15 1 2
5 13 9 1 9 5
14 1 9 1 9 13 15 11 7 13 15 1 1 9 2
17 3 13 15 11 15 13 15 1 9 1 9 1 9 7 1 15 2
5 13 1 14 13 5
9 9 13 15 0 16 15 13 0 2
20 15 13 0 1 16 15 13 1 14 13 2 7 16 9 13 16 15 4 13 2
20 15 13 15 0 0 16 10 9 13 10 9 1 10 3 0 9 1 0 9 2
21 15 4 13 1 7 1 2 7 4 1 9 13 15 1 14 13 10 12 1 9 2
15 3 13 10 9 1 10 9 7 9 16 15 4 13 9 2
3 0 9 5
40 10 0 9 2 7 9 1 14 13 9 2 4 13 1 0 1 9 7 9 1 9 0 9 12 16 0 13 9 2 13 15 1 10 9 7 13 1 11 12 2
15 3 9 10 3 13 9 9 1 16 9 4 13 1 9 2
3 0 9 5
14 9 4 3 13 16 10 9 4 13 1 3 0 9 2
6 11 11 13 0 9 2
29 1 10 9 7 9 1 10 12 0 3 16 9 4 13 2 4 0 13 1 10 3 0 7 1 9 3 0 9 2
26 1 14 13 15 1 1 9 13 9 9 1 10 0 9 3 0 13 9 1 2 0 9 1 15 2 2
29 9 13 3 16 11 2 15 13 9 1 11 2 4 4 13 10 3 0 7 0 9 7 9 16 3 15 4 13 2
4 13 10 9 5
19 16 15 13 9 13 9 1 16 0 4 13 0 1 9 1 12 0 9 2
10 9 4 13 1 10 0 7 0 9 2
5 15 13 10 9 2
3 0 9 5
16 11 4 3 13 15 1 14 13 9 0 9 1 9 1 9 2
13 9 4 1 9 13 1 1 11 1 14 13 9 2
18 13 15 9 4 11 3 13 1 9 2 7 3 4 11 13 11 1 2
7 7 11 4 13 1 11 2
29 9 13 0 1 9 1 10 9 1 15 15 13 1 12 9 3 2 16 11 13 1 1 9 1 0 9 1 11 2
10 10 9 4 9 13 3 0 0 0 2
18 10 10 1 14 13 1 1 9 7 1 1 10 0 9 1 0 9 2
3 11 13 5
7 9 1 11 13 3 9 2
16 11 11 13 15 10 1 16 15 13 10 9 1 9 1 9 2
11 15 15 4 13 2 7 0 0 1 9 2
21 11 11 11 4 13 1 1 9 1 9 1 9 2 7 9 15 0 3 13 9 2
14 11 11 11 4 13 3 1 9 7 13 3 1 3 2
4 0 1 9 2
8 7 11 4 4 13 0 1 2
24 9 13 0 2 16 11 11 13 9 1 10 9 2 7 3 0 16 11 11 13 3 1 9 2
28 7 14 13 9 0 1 11 11 13 3 9 2 7 10 9 4 3 10 9 15 13 9 13 15 14 13 1 2
17 3 13 15 15 10 9 1 2 16 11 11 13 10 9 1 9 2
15 3 15 13 3 0 1 9 15 15 13 0 14 13 1 2
8 14 13 10 9 13 3 9 2
3 0 3 5
15 3 3 13 15 9 16 3 0 9 13 9 14 13 1 2
17 10 9 13 12 2 12 2 3 4 11 11 0 13 1 0 9 2
22 12 9 0 13 11 11 0 1 9 1 16 9 11 11 11 13 10 9 1 1 9 2
11 1 10 9 13 9 11 11 11 3 0 2
14 11 0 9 13 3 1 9 2 9 15 3 4 13 2
12 11 11 4 13 9 1 9 1 10 9 9 2
4 4 13 3 5
21 2 15 13 3 14 13 9 2 15 13 3 0 10 7 9 2 13 9 11 11 2
11 16 1 9 13 0 9 9 1 9 9 2
8 10 9 13 3 3 0 0 2
25 11 13 15 15 13 10 9 3 2 7 11 4 13 1 10 9 7 13 0 7 0 9 1 9 2
11 7 15 13 0 0 1 1 15 11 13 2
2 9 5
8 11 4 13 1 9 1 9 2
6 15 4 13 9 9 2
21 12 1 10 12 0 9 13 1 9 1 9 15 3 13 0 1 9 1 0 9 2
29 3 4 15 3 13 15 1 10 3 0 9 1 9 2 1 10 9 15 3 13 10 0 9 1 14 13 9 12 2
21 1 10 0 9 1 0 9 2 7 9 1 10 0 9 2 4 11 13 1 9 2
4 9 1 11 5
17 11 4 13 10 9 1 9 9 2 15 15 1 9 4 13 1 2
7 10 9 13 9 1 9 2
15 12 9 1 12 9 13 9 1 1 10 0 9 1 9 2
14 2 9 15 4 13 3 1 9 13 0 0 1 15 2
48 10 9 15 4 13 1 3 4 13 0 7 13 10 9 2 0 4 10 9 13 15 2 7 3 13 15 0 16 15 4 13 0 0 9 2 13 10 0 9 11 11 1 9 0 9 1 11 2
5 13 15 1 9 5
24 10 9 15 3 4 13 3 0 16 11 13 9 2 13 16 9 13 15 1 9 1 0 9 2
8 0 9 9 1 11 13 0 2
16 3 1 1 9 13 11 14 13 15 10 9 1 9 1 11 2
16 12 9 2 15 0 11 11 2 13 1 7 3 4 9 13 2
3 11 10 5
11 9 13 15 0 1 3 10 9 1 11 2
21 3 13 15 11 15 13 11 7 1 10 9 13 15 10 9 9 15 4 13 1 2
17 2 9 1 11 13 3 10 0 9 15 4 13 3 0 10 9 2
10 15 13 0 0 7 13 3 0 3 2
13 7 15 13 9 15 4 13 1 2 13 11 11 2
6 9 1 9 1 9 5
22 2 14 13 9 1 9 1 10 9 15 3 4 13 2 4 3 13 1 9 1 11 2
9 2 15 4 4 13 9 1 15 2
16 15 13 3 1 1 9 10 1 9 1 16 15 4 13 9 2
4 0 1 9 5
18 2 15 13 0 1 15 15 4 13 2 13 9 1 10 9 1 11 2
19 15 13 1 0 9 2 0 1 9 7 1 10 9 15 13 13 3 0 2
4 13 15 0 5
18 2 3 4 3 9 13 9 1 14 13 15 1 9 16 9 13 9 2
11 15 13 10 10 9 7 0 9 1 9 2
7 0 4 15 3 13 15 2
26 15 4 3 13 1 0 1 9 16 15 4 13 9 1 1 9 2 13 9 15 3 4 13 12 9 2
5 13 9 7 13 5
17 2 15 4 13 16 9 4 4 13 3 1 9 16 9 4 13 2
8 1 3 12 9 4 9 13 2
11 3 13 3 10 12 0 3 2 13 9 2
15 15 13 16 9 1 9 13 0 1 15 15 0 4 13 2
5 1 10 0 9 5
9 9 13 14 13 1 10 0 9 2
22 1 11 9 2 15 13 9 9 2 13 9 10 0 9 15 0 13 0 1 9 10 2
13 2 13 15 1 16 9 13 1 9 1 9 10 2
16 15 13 9 11 11 2 15 13 10 12 9 0 9 1 11 2
28 1 9 1 9 7 9 9 4 15 13 9 1 1 9 1 9 1 16 9 1 9 1 11 7 11 4 13 2
3 0 9 5
11 9 1 11 7 11 13 0 1 0 9 2
18 7 1 16 11 13 0 2 7 13 10 12 0 9 2 13 9 1 2
19 1 10 0 9 13 9 15 1 12 2 12 2 16 11 13 14 13 9 2
11 2 15 4 13 16 15 13 0 14 13 2
10 9 4 13 3 0 9 3 1 9 2
19 4 15 13 0 0 2 4 15 4 13 10 9 2 13 9 11 11 11 2
3 9 13 5
16 11 4 3 13 9 1 11 1 12 9 2 7 13 9 0 2
25 15 13 3 0 1 16 11 13 0 16 10 9 13 1 0 9 2 7 15 13 9 1 10 9 2
3 1 9 5
16 7 16 11 9 13 1 9 1 9 1 0 9 2 13 9 2
22 15 13 15 9 1 0 9 2 1 1 1 16 9 3 13 9 1 14 13 9 10 2
4 13 3 0 5
9 11 13 10 9 1 0 0 9 2
25 7 11 11 7 11 11 13 9 1 9 2 7 13 1 9 9 16 15 4 13 0 1 11 1 2
5 13 15 1 9 5
17 11 11 4 0 13 11 1 9 2 7 13 15 3 1 9 9 2
11 10 0 0 0 9 4 9 13 9 9 2
21 2 15 13 9 15 4 13 1 9 10 15 3 13 0 1 15 14 13 9 9 2
41 15 13 14 13 10 9 1 9 1 14 4 13 1 10 9 3 0 0 11 13 2 15 13 14 13 0 0 1 9 7 15 13 14 13 0 1 10 0 9 9 2
26 15 13 12 9 0 2 7 4 13 1 16 15 4 13 10 0 9 1 9 1 10 9 1 9 10 2
16 7 9 13 15 3 0 2 13 10 0 0 11 11 1 11 2
24 2 7 3 13 15 1 10 9 1 11 1 9 9 2 1 3 14 13 15 3 3 2 11 2
15 2 15 13 1 0 9 16 15 13 9 1 11 1 9 2
29 15 13 3 9 2 7 3 13 15 0 1 16 15 4 13 9 1 14 13 1 1 9 9 16 15 13 15 3 2
6 7 15 13 15 3 2
22 15 4 13 1 9 0 9 10 2 7 13 10 0 9 1 14 13 10 10 3 3 2
20 15 4 13 15 10 0 9 10 9 2 16 15 13 1 0 3 1 10 9 2
20 13 1 16 3 1 12 9 4 15 13 10 0 9 2 7 15 13 15 0 2
12 15 13 0 9 1 9 10 2 9 1 9 2
43 1 12 9 3 13 11 11 10 9 1 9 11 11 7 0 9 11 11 2 16 15 13 1 10 9 9 15 13 16 15 13 1 14 4 13 1 9 1 11 1 9 9 2
20 15 13 3 10 9 1 11 7 11 2 7 11 9 4 13 1 1 11 9 2
11 7 15 13 1 16 9 13 11 11 9 2
17 3 16 9 1 9 13 14 13 9 1 0 3 16 11 4 13 2
26 2 15 13 3 16 15 13 1 11 2 7 15 13 3 16 11 1 1 9 13 1 15 1 0 9 2
28 15 4 13 10 0 9 1 11 2 7 15 13 0 3 0 0 1 9 15 4 13 1 7 9 10 1 9 2
19 15 13 0 7 0 14 13 0 1 14 13 1 9 10 15 15 10 13 2
17 3 3 13 15 15 0 2 0 2 2 7 15 13 10 0 9 2
16 11 13 3 3 15 15 4 13 1 16 9 9 3 13 0 2
15 2 3 15 13 1 9 2 3 15 13 15 10 0 9 2
27 7 1 9 13 15 1 14 13 1 9 2 7 3 3 4 15 13 1 0 9 15 0 13 14 13 0 2
5 13 14 13 0 2
19 3 1 11 4 15 13 1 14 13 1 9 1 14 13 0 3 1 9 2
34 3 13 15 15 1 10 0 9 1 3 14 4 4 13 15 10 9 1 10 0 0 9 2 7 13 9 1 14 13 1 0 0 9 2
27 7 15 13 16 9 13 1 0 9 3 1 9 2 15 4 3 13 9 1 15 7 13 15 10 0 9 2
4 13 1 11 5
6 2 3 13 9 3 2
19 2 3 13 3 15 16 15 13 1 1 9 11 2 7 15 13 3 3 2
17 15 13 0 10 0 9 1 14 13 0 1 11 1 10 9 1 2
29 15 13 9 1 11 2 7 15 13 3 16 15 13 0 1 9 7 1 9 1 10 0 0 1 0 12 9 3 2
31 15 4 13 1 11 9 3 12 9 10 9 9 16 15 13 3 2 15 4 13 12 9 1 11 2 7 15 13 3 0 2
5 15 13 3 0 2
23 15 13 3 14 13 10 0 9 1 9 1 10 0 9 10 9 1 11 9 13 1 15 2
26 15 13 3 1 9 2 7 13 16 10 0 13 1 2 13 11 2 7 13 1 1 9 1 0 9 2
9 2 0 3 4 15 13 1 9 2
10 15 13 14 13 2 0 3 1 9 2
20 7 3 1 10 9 2 15 13 3 16 15 13 0 9 3 2 13 15 0 2
4 9 1 9 2
8 2 3 13 10 9 1 9 2
9 2 3 13 15 1 9 1 9 2
21 15 13 10 0 9 1 14 13 11 1 0 9 1 9 2 7 15 4 15 13 2
32 15 13 0 16 15 4 13 10 9 9 1 9 7 3 13 9 2 7 15 13 15 3 0 10 1 9 15 13 2 13 15 2
19 15 13 16 9 1 11 13 14 13 0 0 3 16 11 3 13 7 13 2
23 7 15 4 3 13 15 1 15 11 13 15 2 15 4 3 13 1 14 13 0 3 3 2
8 2 15 13 10 9 1 9 2
13 2 15 13 3 10 9 2 1 14 13 15 3 2
36 7 9 4 0 13 10 9 16 15 13 14 13 10 9 15 7 11 11 4 13 1 2 7 16 15 13 14 13 10 9 0 0 15 9 13 2
25 16 9 13 14 13 1 10 9 1 3 2 13 15 16 9 4 13 1 11 9 1 10 0 9 2
19 16 11 4 13 15 1 0 0 9 4 3 11 11 11 13 10 0 9 2
23 15 13 3 0 9 1 10 9 2 7 11 13 10 0 10 9 9 1 15 11 3 13 2
22 7 15 13 0 3 1 14 13 16 15 0 3 13 0 16 10 9 13 10 12 0 2
13 3 10 0 9 4 13 1 10 0 1 11 3 2
4 15 3 13 2
15 11 11 13 16 15 0 3 4 13 10 9 1 10 9 2
2 9 5
26 2 15 13 14 13 15 1 0 9 3 2 7 15 13 0 0 16 15 3 13 9 1 10 0 9 2
18 15 13 14 13 9 1 10 9 1 9 2 7 15 13 0 0 9 2
30 13 1 16 15 4 13 9 16 15 13 12 9 2 13 11 2 7 13 1 10 9 1 11 2 11 2 11 7 11 2
34 2 15 4 13 1 1 14 13 1 3 12 9 1 11 2 7 3 13 15 0 0 9 1 14 13 1 0 9 3 1 11 10 9 2
25 7 15 13 3 10 9 2 15 4 3 13 1 15 14 13 3 16 15 13 1 9 1 9 3 2
12 2 10 9 4 15 13 1 9 2 13 15 2
23 2 15 13 12 9 15 13 1 2 7 15 13 16 15 13 1 0 9 1 11 1 11 2
16 15 13 9 2 7 4 13 0 1 10 0 12 2 12 9 2
14 10 9 13 15 1 12 9 2 7 15 13 15 0 2
8 15 13 10 9 9 1 9 2
5 13 14 13 9 5
26 12 9 1 11 13 14 3 13 9 10 1 11 9 16 3 11 9 13 15 1 14 13 9 1 9 2
11 2 1 10 0 9 13 9 12 9 0 2
14 1 9 4 15 13 10 1 10 0 0 9 1 9 2
27 16 15 4 13 10 9 15 13 0 16 15 13 0 0 1 9 2 13 9 1 10 0 9 1 11 9 2
19 15 13 9 9 16 10 9 15 13 9 1 0 9 4 13 1 0 9 2
13 1 9 15 13 0 1 11 2 13 15 12 9 2
24 15 13 3 3 3 14 13 15 1 16 12 9 4 13 15 1 1 9 1 9 2 13 9 2
40 2 15 13 3 0 1 10 9 2 16 16 15 4 13 1 9 2 4 15 13 15 0 1 14 13 13 14 13 9 10 1 9 2 13 9 1 9 1 9 2
6 9 13 1 1 9 5
9 10 0 9 4 3 13 1 9 2
19 15 13 10 0 9 1 0 0 9 1 9 2 13 9 11 11 1 11 2
14 1 9 13 11 11 10 9 1 12 1 9 1 9 2
24 9 4 3 13 1 1 9 2 15 13 10 9 15 13 1 9 10 9 1 10 0 1 9 2
12 10 9 13 16 9 13 16 9 13 12 9 2
7 10 9 4 15 3 13 2
29 2 15 4 13 15 13 3 14 4 13 9 1 9 7 1 9 7 3 1 9 2 13 15 15 13 11 1 11 2
23 9 13 0 9 1 9 2 7 11 11 13 3 16 9 4 13 1 14 13 9 1 9 2
14 0 4 15 13 1 14 13 0 9 1 1 10 9 2
16 9 15 4 13 1 9 2 4 0 13 7 1 9 7 10 2
24 10 9 1 9 13 12 1 9 1 9 1 0 2 16 12 1 15 4 13 9 1 0 9 2
11 9 11 11 13 16 9 13 1 9 1 2
9 15 13 3 16 15 3 13 0 2
11 7 15 4 13 1 14 13 1 1 15 2
21 2 1 9 13 15 9 1 16 15 4 13 1 1 9 7 14 13 9 1 9 2
15 1 10 9 13 10 9 1 7 1 10 13 15 1 9 2
26 15 13 10 9 15 13 9 2 7 15 4 13 3 1 15 7 13 1 1 10 9 2 13 11 11 2
8 11 11 13 2 9 9 2 5
38 1 0 9 1 12 9 1 10 0 9 4 11 11 1 11 13 1 2 11 11 2 7 13 0 10 0 9 16 10 0 9 1 11 4 13 0 9 2
8 9 13 15 1 10 0 9 2
30 7 3 0 1 11 2 15 1 0 13 11 11 2 4 13 9 1 10 9 1 9 1 15 2 10 0 11 1 11 2
28 11 11 7 11 11 1 11 11 1 11 13 1 10 0 9 2 11 8 8 2 15 0 1 9 1 0 9 2
8 10 0 9 1 10 0 9 2
33 10 0 12 0 9 4 0 13 16 11 11 11 11 11 13 0 9 16 15 1 9 1 2 11 9 2 2 13 9 1 0 9 2
19 9 4 3 13 1 16 11 9 13 9 0 9 1 2 11 7 11 2 2
59 3 10 9 1 11 11 11 13 1 1 9 1 16 9 4 13 2 7 15 4 13 11 11 11 10 9 16 15 1 10 9 4 13 1 15 10 10 9 15 13 1 1 14 13 10 0 9 2 16 9 13 0 7 16 15 13 0 15 2
20 15 13 1 0 2 11 9 2 15 13 0 9 1 9 1 9 2 7 9 2
12 7 15 13 3 10 9 1 10 9 1 9 2
15 11 11 13 10 9 2 3 9 11 11 7 9 11 11 2
17 10 0 9 1 9 11 11 15 1 10 9 4 13 10 0 9 2
31 3 9 2 7 2 9 2 15 9 10 13 2 11 11 11 2 4 13 9 1 10 0 9 15 4 13 1 1 9 9 2
21 7 1 9 1 9 0 9 2 13 15 3 14 13 11 1 9 1 9 7 9 2
19 3 13 0 1 12 9 15 2 7 1 15 13 7 9 7 0 0 9 2
6 9 11 11 13 0 2
7 2 3 4 15 13 9 2
27 0 0 16 15 13 3 15 4 13 2 1 12 4 13 1 9 1 9 7 0 4 13 1 9 10 3 2
43 15 13 10 0 9 14 13 10 9 2 0 9 2 1 15 1 9 3 2 4 13 1 1 9 7 9 2 7 3 13 15 0 14 13 2 13 10 0 2 7 0 11 2
7 9 2 7 9 1 9 5
9 1 12 13 11 11 1 11 11 2
16 1 9 13 9 3 3 0 1 9 1 10 0 9 1 3 2
10 9 13 0 9 7 10 0 9 9 2
15 9 13 1 11 11 2 15 13 9 1 1 12 9 9 2
13 1 11 9 1 9 11 9 1 11 13 9 0 2
9 3 0 7 9 13 15 15 13 2
14 9 13 1 2 7 9 13 1 9 7 0 7 0 2
19 3 0 16 9 10 13 9 1 14 13 9 1 15 9 13 2 7 3 2
7 9 13 0 1 9 9 2
10 9 1 15 13 16 9 13 1 9 2
28 16 15 13 1 9 7 16 11 11 13 0 1 14 13 1 1 15 1 10 9 2 4 9 13 1 12 9 2
23 2 13 15 0 1 1 10 9 15 4 13 2 13 15 12 9 0 2 2 13 15 15 2
5 2 6 2 6 2
14 15 4 3 13 16 15 3 13 9 2 13 11 15 2
16 15 13 15 0 1 2 7 9 1 10 9 13 3 1 9 2
8 15 4 13 0 1 10 9 2
16 2 4 15 13 10 9 1 9 2 4 15 13 1 10 9 2
22 7 9 13 3 0 2 7 1 10 9 2 15 13 9 16 15 13 15 2 13 11 2
13 2 15 13 9 1 14 13 12 9 7 10 9 2
10 2 1 10 9 13 15 10 9 0 2
14 15 13 9 2 13 11 2 13 1 9 7 13 1 2
16 2 15 15 4 13 1 15 1 3 2 13 3 0 1 9 2
10 1 15 13 15 9 1 9 15 13 2
20 16 15 13 9 1 10 9 15 13 10 9 2 4 15 13 1 9 0 0 2
17 2 15 4 3 13 0 14 4 13 9 1 7 15 7 10 9 2
5 2 15 13 0 2
15 1 3 15 4 13 2 3 4 15 3 13 3 1 15 2
17 16 0 1 10 10 1 9 4 13 15 0 9 2 13 3 0 2
11 7 1 15 10 7 1 9 2 13 11 2
10 15 4 13 1 10 0 9 1 9 2
17 1 9 13 10 10 10 9 15 4 13 1 11 7 13 15 0 2
17 2 0 13 0 1 2 7 4 1 9 4 13 1 10 0 9 2
12 1 9 13 15 10 9 15 4 13 0 9 2
9 3 15 4 1 10 9 13 0 2
5 16 15 13 0 2
8 0 15 13 15 2 13 11 2
17 0 1 9 1 9 4 13 15 1 10 9 1 11 11 10 9 2
13 11 11 13 3 10 9 15 4 13 11 11 0 2
11 9 4 15 3 13 15 9 13 1 9 2
19 2 15 4 13 10 9 2 7 4 3 13 10 0 2 13 9 11 11 2
10 3 4 15 3 13 15 15 1 9 2
11 1 10 9 4 10 9 3 13 1 9 2
24 3 13 11 11 10 9 0 14 13 15 1 2 16 15 13 16 15 4 13 12 9 1 9 2
14 2 15 13 3 0 2 13 15 7 13 15 0 1 2
12 4 15 13 2 4 11 13 0 1 12 9 2
5 0 7 0 11 5
14 2 15 4 3 3 13 0 14 13 1 10 0 9 2
36 3 4 3 9 13 15 1 14 13 9 9 10 2 3 14 13 15 1 1 9 7 13 15 1 16 11 11 13 9 7 13 14 13 9 3 2
10 15 13 11 0 9 11 11 1 11 2
36 1 3 4 9 4 13 1 2 10 9 2 1 10 0 9 2 3 13 15 16 9 13 1 1 14 13 15 1 15 15 4 13 10 0 9 2
36 10 0 11 7 11 9 4 1 9 13 15 1 1 9 9 2 7 13 3 0 1 9 9 1 11 16 9 4 13 15 9 7 10 9 9 2
18 1 14 4 13 10 9 9 7 13 15 3 1 10 9 9 1 11 2
12 2 0 9 13 0 2 7 1 15 7 9 2
40 15 13 0 1 9 15 13 1 10 9 2 7 15 13 3 10 9 15 4 13 3 1 9 15 3 4 13 9 2 1 16 15 13 1 0 1 9 9 1 2
12 15 13 3 1 9 2 13 10 0 0 11 2
5 2 3 0 3 2
25 15 13 9 9 1 14 13 0 9 7 13 9 1 16 9 13 14 13 9 1 15 15 4 13 2
29 11 9 1 14 13 1 11 0 9 7 9 15 13 9 1 14 4 13 10 9 2 13 15 0 7 0 1 1 2
22 7 15 11 0 1 15 13 3 2 13 0 9 1 9 1 9 7 9 2 3 9 2
13 2 15 4 13 3 9 7 0 9 1 15 3 2
24 0 9 2 0 9 2 0 9 2 0 1 9 7 0 0 9 4 3 4 13 9 3 0 2
24 1 0 9 13 15 3 9 2 7 15 3 4 13 9 7 13 0 3 1 14 13 0 0 2
37 15 13 3 9 0 2 7 4 13 0 1 2 13 9 11 2 15 3 13 16 15 3 13 0 0 1 16 15 13 10 12 1 9 15 13 9 2
3 13 9 5
26 3 13 15 16 16 10 0 9 4 13 15 2 4 3 7 15 1 9 7 9 1 9 4 13 15 2
8 2 15 4 13 9 1 15 2
23 15 13 15 3 10 10 15 13 1 1 9 1 15 7 3 0 4 13 9 2 4 13 2
35 3 13 15 3 16 9 1 9 3 13 9 1 10 0 9 1 0 9 1 9 7 9 2 16 15 4 4 13 1 9 1 9 7 9 2
32 1 9 16 15 4 13 1 9 7 9 2 13 7 9 7 9 1 15 0 3 16 15 13 1 9 1 15 2 13 11 11 2
5 11 0 1 9 5
17 2 15 13 0 1 3 10 9 4 13 15 9 1 9 1 9 2
18 1 9 4 15 3 13 0 3 0 0 1 9 2 13 9 11 11 2
27 2 15 13 16 15 4 13 0 14 13 9 1 9 1 10 9 2 7 13 9 13 15 2 13 15 1 2
11 9 11 4 13 0 1 9 1 9 9 2
11 2 15 13 3 0 1 1 9 1 9 2
36 15 13 0 0 9 1 9 1 9 2 3 4 15 3 13 1 1 10 9 3 2 13 11 2 15 1 10 9 13 16 11 11 3 4 13 2
35 2 7 11 13 15 0 0 9 1 2 0 13 15 0 0 2 7 15 4 13 10 9 13 15 0 3 16 15 4 13 3 0 15 13 2
26 1 9 9 1 9 2 16 15 13 12 2 12 1 11 2 13 11 7 0 7 0 7 13 12 9 2
10 15 13 10 1 15 15 13 1 15 2
20 13 15 3 9 1 2 9 2 10 2 4 15 13 0 0 2 13 11 11 2
5 9 13 1 11 5
27 1 12 9 4 15 13 10 0 9 1 9 1 11 2 7 3 0 13 9 1 11 7 11 1 1 3 2
21 7 3 2 0 1 9 13 9 0 1 15 15 13 0 1 1 10 0 12 9 2
11 7 15 13 3 1 14 13 12 2 12 2
19 9 1 11 13 3 3 1 1 14 13 15 0 9 1 9 1 11 9 2
28 7 15 13 0 1 10 0 9 2 7 1 12 9 1 9 13 15 1 1 16 9 7 0 9 4 13 9 2
17 1 1 3 13 3 11 1 1 10 9 15 9 1 9 4 13 2
13 2 15 15 13 10 0 12 9 13 0 1 15 2
16 0 0 2 2 13 10 0 0 9 2 11 11 2 1 9 2
6 2 9 13 0 3 2
21 14 13 12 2 12 1 10 9 13 0 0 2 7 9 1 9 13 0 1 0 2
13 3 0 13 15 3 15 4 13 2 13 15 1 2
5 0 9 1 9 5
25 9 13 1 0 0 1 11 9 2 7 1 10 0 9 13 9 1 0 9 1 11 11 1 9 2
31 1 10 9 13 15 3 0 1 7 13 16 9 4 13 1 9 2 7 9 1 10 9 1 11 10 0 13 14 13 9 2
17 9 1 15 13 16 15 3 4 13 0 1 9 1 10 10 9 2
24 3 12 0 9 4 13 2 7 1 10 10 9 4 15 13 0 1 14 13 10 9 1 9 2
14 2 15 13 3 14 13 15 15 15 4 13 1 9 2
22 15 13 3 9 1 9 2 10 0 9 13 3 2 9 13 3 0 7 9 13 3 2
29 0 13 15 3 9 1 9 0 3 2 7 10 9 15 13 3 13 9 3 0 2 13 11 11 2 9 0 9 2
18 1 1 1 0 9 10 0 9 13 15 0 7 13 1 10 0 9 2
12 15 13 0 1 9 7 13 0 14 13 15 2
17 4 0 1 11 9 13 10 9 1 9 4 3 9 13 0 1 2
34 1 9 13 15 0 9 13 1 9 2 11 4 13 1 14 13 9 3 2 7 4 3 13 1 10 0 9 16 15 13 15 9 9 2
3 9 13 5
23 1 9 13 9 11 9 1 10 9 2 0 15 15 13 1 11 11 11 1 11 11 11 2
4 10 9 13 2
22 11 4 13 9 0 2 15 13 0 1 9 2 7 15 13 0 0 9 1 0 9 2
17 9 13 2 7 15 13 0 7 0 16 11 1 9 4 13 9 2
10 1 10 0 9 13 15 9 1 9 2
23 1 10 0 9 13 11 11 11 0 0 3 1 0 9 2 7 13 0 1 9 11 11 2
23 11 4 3 13 1 10 9 1 0 1 3 14 13 2 7 13 1 3 11 1 1 9 2
16 12 9 0 13 15 10 10 9 2 11 11 2 15 13 1 2
28 1 10 0 9 1 11 7 11 11 11 13 9 1 9 1 11 2 15 13 15 0 16 15 13 1 12 9 2
10 3 1 13 15 15 14 13 1 9 2
9 0 1 1 9 0 9 1 9 2
11 12 9 1 9 4 15 13 1 11 9 2
24 1 10 9 4 15 13 9 2 1 14 13 9 1 11 9 16 15 13 1 1 14 13 9 2
19 2 15 13 12 2 12 2 13 15 14 13 1 1 9 16 9 4 13 2
5 7 1 1 9 5
16 2 2 11 2 13 15 1 1 9 7 13 1 10 0 9 2
11 3 13 4 11 13 12 0 9 1 9 2
14 2 15 15 13 1 1 9 1 9 13 0 1 9 2
25 11 11 11 13 0 0 2 11 11 11 13 16 15 0 13 0 2 7 11 11 13 10 0 9 2
28 7 1 13 13 9 3 0 1 9 2 7 15 4 13 0 0 4 15 13 0 9 1 9 11 2 13 11 2
14 10 9 4 11 13 15 0 9 2 1 9 1 11 5
14 2 15 13 0 14 13 1 10 9 2 13 11 0 2
11 1 11 4 3 3 13 15 1 11 11 2
10 15 13 15 10 0 0 0 1 9 2
5 9 7 0 9 5
2 11 2
20 9 13 10 0 9 1 9 1 9 11 11 7 11 11 2 11 2 11 11 2
24 15 13 15 1 10 9 2 13 15 1 9 1 12 9 3 2 7 13 0 1 9 1 11 2
13 2 15 4 13 1 1 10 9 1 9 1 12 2
17 1 10 4 15 13 10 0 9 1 11 11 7 11 11 1 12 2
13 10 9 1 9 13 15 0 3 15 13 1 11 2
14 7 10 3 0 9 13 3 9 1 11 11 1 12 2
17 2 11 13 1 9 2 2 13 9 11 11 2 13 11 11 11 2
27 3 13 15 10 0 9 15 4 13 1 0 1 9 2 0 0 3 1 11 11 2 7 9 1 11 11 2
11 1 0 9 13 15 10 0 9 1 9 2
18 10 9 4 15 7 9 13 1 11 1 10 9 2 13 15 7 13 2
3 1 11 5
20 9 11 11 2 0 1 11 1 11 2 13 3 9 1 12 1 10 0 9 2
13 15 13 14 13 1 9 1 11 1 9 1 9 2
10 3 15 13 9 1 9 2 13 15 2
22 16 15 13 3 0 1 9 2 13 15 0 0 16 15 13 14 13 15 1 10 9 2
7 15 13 0 9 1 12 2
9 11 13 16 15 13 10 0 9 2
22 1 16 15 4 13 1 9 2 13 15 9 1 0 9 2 9 7 9 1 11 11 2
9 2 11 11 13 1 10 10 9 2
12 7 15 13 3 1 1 14 13 3 1 15 2
8 15 4 0 13 2 13 11 2
5 2 11 11 2 5
20 3 13 15 0 9 1 9 10 2 3 16 10 10 4 4 0 13 1 9 2
17 15 13 1 1 11 11 2 15 13 9 2 11 11 2 1 11 2
16 3 4 15 13 9 10 9 10 9 2 3 13 11 10 9 2
14 7 15 4 0 13 1 9 1 14 13 1 0 9 2
15 3 13 11 11 1 1 9 1 11 11 9 1 11 9 2
8 2 11 11 13 10 0 9 2
9 1 12 9 3 13 15 10 9 2
24 10 9 0 13 15 9 2 7 15 13 1 10 9 1 11 11 7 11 11 11 1 11 11 2
7 15 13 10 0 0 9 2
10 9 13 15 3 0 7 0 10 9 2
17 10 0 13 3 0 0 1 9 1 10 9 15 13 1 1 1 2
24 1 16 9 13 1 7 9 4 13 1 2 13 15 0 0 3 1 9 16 15 13 9 13 2
14 1 9 13 3 10 9 1 15 7 13 3 1 15 2
16 15 13 10 0 0 9 1 7 0 7 0 2 13 11 11 2
2 0 5
27 3 16 15 13 9 7 9 2 4 0 11 11 11 13 0 1 10 0 9 15 11 4 13 10 0 9 2
14 15 13 0 16 9 7 9 4 13 3 0 14 13 2
15 2 15 13 3 16 9 13 0 1 9 15 3 13 9 2
19 7 15 4 13 0 1 10 9 1 9 15 3 13 15 1 9 14 13 2
21 6 2 15 13 3 1 7 1 13 9 2 1 11 11 2 15 13 10 0 9 2
15 15 13 10 1 15 1 10 9 14 13 2 13 11 11 2
10 2 7 15 13 3 1 9 1 11 2
7 2 6 2 15 13 15 2
7 15 13 15 0 2 15 2
2 9 5
14 11 11 13 3 0 9 1 9 1 9 1 9 9 2
11 2 15 13 3 10 0 9 1 9 3 2
12 15 13 3 0 0 2 15 15 13 0 0 2
6 7 0 0 1 15 2
9 15 13 9 1 11 3 1 9 2
8 1 0 9 13 15 3 15 2
22 3 13 15 3 0 9 10 12 9 9 1 1 2 11 11 2 2 13 11 11 11 2
6 9 1 11 1 9 5
3 13 9 5
4 9 0 9 5
13 11 9 4 13 9 1 9 1 14 13 1 9 2
14 11 11 11 2 9 1 11 9 2 3 0 1 9 2
7 11 13 0 0 9 12 2
17 9 2 0 2 3 0 2 4 0 1 1 3 4 13 1 9 2
6 9 2 11 11 11 5
9 13 0 10 9 1 11 9 9 5
25 2 15 4 13 9 1 16 15 4 13 1 9 2 13 11 11 11 2 9 1 11 9 1 11 2
23 0 0 4 13 7 13 1 9 1 14 13 2 1 9 1 10 0 9 1 9 0 9 2
21 9 1 11 11 7 11 4 3 13 10 9 1 9 1 3 9 1 11 4 13 2
28 15 9 4 13 13 16 15 3 4 13 1 16 0 9 1 11 9 1 11 7 1 11 9 1 11 4 13 2
13 3 4 15 13 10 9 7 9 16 9 4 13 2
3 13 3 2
7 2 4 13 15 10 9 5
3 13 3 2
5 13 9 1 11 5
3 13 3 2
4 9 1 9 5
20 2 9 13 14 13 16 9 13 2 13 0 9 11 11 1 11 11 7 11 2
8 9 1 9 13 1 10 9 2
10 11 13 10 12 9 1 9 1 9 2
12 3 9 1 10 0 2 0 9 13 9 3 2
8 2 15 13 3 0 1 9 2
26 10 9 9 13 9 1 14 13 14 4 13 1 9 2 7 13 15 3 13 1 15 14 13 10 9 2
21 0 9 4 3 13 0 9 2 0 1 15 15 13 1 9 10 2 13 9 11 2
31 16 3 9 13 9 1 9 9 2 4 10 12 9 13 2 7 4 3 13 1 12 9 1 11 9 7 12 1 11 9 2
9 13 0 10 9 1 11 9 9 5
8 9 13 9 13 9 1 9 5
5 11 2 11 2 2
31 9 4 13 1 9 16 15 13 10 9 1 9 1 9 13 9 11 1 11 1 16 15 4 13 9 1 9 9 1 9 2
13 2 15 13 3 14 13 1 1 3 0 9 3 2
36 15 15 4 13 13 16 15 3 13 10 0 9 2 7 16 9 0 13 12 2 12 9 0 2 13 9 11 11 1 11 9 1 11 1 11 2
18 9 4 3 13 9 15 4 13 2 7 4 13 15 12 2 12 9 2
25 15 4 3 13 16 15 13 9 15 4 13 2 7 11 13 16 9 3 13 0 0 1 10 9 2
15 2 15 13 3 3 0 14 13 10 9 15 13 1 9 2
24 15 4 1 10 13 1 3 15 15 13 2 13 14 13 1 15 10 9 1 9 2 13 15 2
12 9 13 1 0 9 7 9 1 9 1 9 2
27 2 15 4 3 13 1 10 9 1 10 9 2 7 15 4 4 13 1 10 9 9 1 9 2 13 9 2
22 0 9 1 9 4 10 9 13 1 9 1 16 15 4 13 9 1 9 1 11 9 2
34 2 15 13 0 16 15 13 15 15 13 0 14 13 0 1 2 7 3 4 9 13 16 15 13 10 9 1 10 12 9 2 13 11 2
4 2 11 2 5
5 9 13 1 9 5
6 9 2 9 7 9 5
2 9 5
5 0 9 1 9 5
20 0 10 9 1 9 1 11 2 7 11 7 11 13 1 9 15 4 13 9 2
10 3 13 9 1 1 9 0 1 9 2
8 9 4 15 13 9 1 9 2
9 9 2 11 2 11 2 11 2 5
22 9 7 9 4 13 1 9 1 11 10 0 9 2 7 10 9 13 9 1 0 1 2
13 9 13 0 9 1 11 7 1 2 7 1 11 2
22 1 11 7 11 10 9 13 15 3 1 1 7 1 9 2 1 0 9 0 9 9 2
23 1 10 0 4 15 13 1 9 2 7 1 9 13 15 10 9 7 9 2 7 3 9 2
4 3 0 9 2
7 3 13 9 16 15 13 5
28 15 13 15 0 9 0 1 1 11 7 11 1 9 9 2 1 9 1 1 0 7 0 9 1 9 0 1 2
14 3 3 13 15 0 9 2 15 13 1 9 1 9 2
11 9 4 1 10 0 13 15 1 12 9 2
17 10 9 13 9 9 1 9 1 7 4 3 13 11 7 9 1 2
23 9 13 3 1 9 2 3 1 9 1 9 2 13 0 9 11 11 1 11 9 1 11 2
9 0 9 1 9 13 9 1 9 2
17 1 9 1 10 9 9 9 4 15 13 1 12 7 12 9 9 2
23 9 13 15 0 9 16 9 4 13 14 13 1 9 2 7 15 4 3 13 9 1 11 2
14 2 1 9 13 15 9 7 0 9 2 13 9 11 2
13 3 13 15 9 1 10 0 9 1 3 0 9 2
16 9 7 9 1 12 9 4 9 13 9 0 1 9 1 11 2
21 1 9 13 15 9 9 13 0 9 7 0 0 9 1 0 9 1 11 7 11 2
17 2 9 13 9 1 11 7 1 0 0 9 1 9 2 13 9 2
27 1 1 9 4 15 3 13 10 10 9 1 1 1 2 7 1 11 4 15 13 0 9 1 0 9 9 2
4 9 7 9 5
2 9 5
8 9 13 9 1 9 1 11 2
17 9 13 10 9 2 0 0 2 1 9 1 10 0 9 1 11 2
8 9 2 11 11 5 11 11 5
20 9 4 13 14 13 9 1 9 1 11 0 9 1 9 2 16 12 9 13 2
3 13 3 2
5 12 13 1 9 5
21 9 1 16 9 13 2 13 16 9 13 16 15 15 13 9 2 3 13 1 9 2
38 2 9 1 9 13 14 13 16 9 4 13 1 1 9 7 1 1 9 2 3 16 15 13 10 0 9 2 9 2 1 11 2 13 9 1 10 9 2
3 13 3 2
5 2 13 0 9 5
21 2 9 15 15 13 13 9 13 0 0 1 9 2 13 9 11 11 1 11 9 2
14 1 15 11 13 1 4 9 4 13 10 9 1 12 2
24 2 15 4 15 3 13 2 7 15 15 4 13 13 16 9 13 1 15 15 13 0 1 9 2
13 7 9 13 3 0 0 2 13 11 11 1 11 2
21 15 4 3 13 15 1 9 1 1 9 2 7 13 16 15 13 9 0 1 9 2
7 1 9 4 15 3 13 2
3 13 3 2
6 2 13 9 1 9 5
3 13 9 5
17 9 11 11 13 1 9 0 9 11 11 0 0 9 1 0 11 2
13 9 11 11 13 1 11 11 0 0 9 1 11 2
8 9 2 11 11 11 5 11 5
16 9 4 13 10 0 7 0 0 0 9 1 9 1 0 9 2
15 2 9 1 11 11 11 11 11 13 10 9 1 11 11 2
40 9 13 3 3 10 0 9 1 10 0 9 7 9 2 7 3 10 9 1 10 9 15 13 15 1 10 0 9 1 11 2 13 0 9 1 9 2 11 11 2
21 11 13 16 9 13 10 9 1 10 0 9 1 0 9 1 10 0 9 1 11 2
21 0 0 9 7 10 0 9 1 9 2 9 7 9 4 13 10 9 1 0 9 2
29 2 9 1 11 4 13 1 1 10 0 9 1 11 1 11 2 11 11 7 9 11 11 11 2 11 2 1 11 2
23 11 11 13 14 13 10 0 9 1 9 1 9 1 9 2 9 7 9 2 13 11 11 2
28 9 1 9 1 11 4 13 1 9 1 11 1 11 2 7 9 1 11 13 1 9 1 10 0 9 1 11 2
16 10 0 9 1 11 2 11 11 7 11 1 11 13 0 9 2
18 10 9 7 9 1 9 13 9 1 0 9 2 7 9 13 0 9 2
7 9 13 1 9 12 0 2
9 9 2 7 3 9 1 11 11 5
5 11 2 11 2 2
22 1 10 0 9 1 9 13 9 1 11 11 9 1 10 9 1 12 9 1 12 9 2
15 1 15 12 9 1 9 13 16 12 13 7 12 13 0 2
22 3 16 0 3 13 0 9 1 9 1 0 1 9 2 13 15 3 9 15 13 9 2
34 3 16 0 13 1 10 9 2 13 15 3 0 9 1 16 10 0 0 9 13 10 0 9 1 9 2 0 0 1 3 15 4 13 2
23 9 13 3 0 1 12 9 7 3 13 15 0 15 13 1 16 9 1 9 4 4 13 2
14 1 12 9 1 9 13 15 0 0 0 9 15 13 2
9 1 9 11 13 9 10 3 0 2
22 9 7 9 1 0 9 9 1 13 16 9 3 13 15 0 1 14 13 10 9 0 2
14 3 13 9 1 11 1 11 9 1 10 0 9 3 2
9 9 13 3 0 0 1 12 9 2
23 9 13 0 1 1 9 1 10 1 9 2 11 2 16 9 3 13 10 9 1 12 9 2
4 2 11 2 5
7 13 9 2 13 1 9 5
10 12 9 13 1 11 1 14 13 9 2
13 1 9 13 12 1 15 1 1 2 13 11 11 2
4 11 11 11 5
5 9 2 11 11 5
28 2 15 13 1 9 1 10 9 7 13 1 10 0 12 2 2 13 11 11 11 1 10 9 1 11 11 9 2
16 11 11 11 7 11 11 11 7 11 11 11 13 1 1 9 2
18 10 0 9 13 1 11 1 9 9 1 14 13 1 10 9 1 11 2
15 7 9 13 3 12 1 15 9 7 13 1 9 1 9 2
18 2 11 13 12 9 1 16 11 4 13 1 9 1 11 2 13 11 2
4 11 13 11 5
3 0 9 5
4 9 3 3 5
3 4 13 5
26 2 13 11 1 1 11 1 0 9 7 0 9 2 13 15 0 2 13 9 1 11 2 11 11 11 2
27 15 13 1 16 0 9 1 9 13 0 7 0 1 10 9 9 15 15 4 13 1 1 16 11 11 13 2
18 11 13 16 9 13 16 9 15 13 1 11 4 4 13 1 0 9 2
17 1 9 1 11 7 11 13 15 10 9 1 0 9 1 0 9 2
6 2 15 13 0 0 2
21 15 1 11 4 3 1 10 10 9 0 9 13 9 1 10 9 1 9 1 9 2
32 15 13 3 2 3 15 13 15 1 11 7 11 2 16 15 4 13 9 15 13 3 2 7 16 0 9 4 13 2 13 11 2
17 9 4 3 4 13 1 0 9 1 9 11 11 7 9 11 11 2
11 2 15 1 11 13 9 1 15 1 9 2
7 15 4 3 3 13 9 2
16 1 9 13 15 1 9 7 13 16 15 3 0 4 13 0 2
37 15 13 1 16 9 9 15 13 0 9 9 1 0 9 9 2 3 13 1 9 1 14 4 13 1 10 9 15 4 13 1 0 0 9 1 9 2
23 2 16 11 13 9 1 11 2 13 9 1 11 7 13 9 9 3 13 3 15 10 9 2
14 15 4 3 13 1 9 7 15 4 3 13 1 9 2
16 15 4 13 7 0 9 7 9 1 10 0 9 2 13 11 2
27 15 13 16 3 0 1 10 0 9 1 0 9 10 0 9 4 13 1 9 7 13 0 9 1 0 9 2
23 2 11 13 10 1 10 9 15 4 13 15 2 7 15 4 3 0 13 1 3 0 9 2
17 7 16 11 13 1 0 9 4 0 9 1 9 1 11 13 15 2
10 2 3 4 3 9 13 1 9 9 2
21 2 3 0 15 3 4 13 10 0 9 1 9 1 11 2 13 15 3 3 9 2
29 3 13 15 16 9 13 14 13 1 9 11 13 1 1 1 10 9 7 13 1 9 10 9 1 9 2 13 11 2
5 2 3 0 0 5
2 0 5
19 9 15 4 13 1 9 1 11 11 1 11 13 3 0 0 2 1 9 2
18 9 1 11 11 1 11 16 11 11 4 13 0 1 10 9 1 9 2
7 9 2 11 2 11 11 5
14 9 4 1 9 13 1 12 0 9 2 13 11 11 2
3 13 3 2
4 9 1 11 5
45 9 1 9 4 13 10 0 9 1 9 2 16 9 1 9 13 16 15 3 13 15 1 16 15 13 1 9 1 10 0 7 10 9 2 16 15 13 1 15 10 1 9 1 9 2
3 13 3 2
2 9 2
5 2 11 4 13 5
23 0 1 9 2 9 11 11 2 4 3 13 1 1 0 9 2 7 13 16 0 13 0 2
9 2 15 13 3 3 0 0 0 2
12 15 13 3 3 10 0 2 13 11 1 9 2
18 9 13 3 1 10 0 9 2 7 13 14 13 0 1 9 1 9 2
15 1 0 4 9 13 1 1 9 1 9 1 9 10 9 2
5 9 13 1 9 5
3 13 9 5
3 12 13 5
2 13 5
6 9 13 9 1 9 2
2 9 5
5 9 2 11 11 5
20 9 13 16 10 9 13 1 10 12 0 1 9 15 13 1 9 1 11 9 2
25 2 15 4 13 16 10 9 1 10 9 4 13 7 13 2 13 9 11 11 1 11 9 1 11 2
25 9 13 0 1 9 1 9 2 7 15 13 9 11 11 1 11 9 15 13 15 1 9 1 9 2
22 15 13 16 9 4 13 1 16 15 4 13 9 1 9 1 10 9 1 9 1 11 2
19 2 15 4 13 9 1 9 15 4 13 1 9 2 13 11 11 1 11 2
9 15 13 16 9 4 13 7 13 2
11 2 15 4 3 13 9 1 9 1 9 2
16 3 13 15 3 10 9 9 15 4 13 1 9 7 10 9 2
10 15 13 3 0 1 9 2 13 11 2
16 11 13 16 12 9 3 0 4 13 1 12 9 1 1 9 2
26 9 13 10 9 1 11 9 2 16 10 9 1 9 4 13 2 0 1 9 1 10 9 1 12 9 2
24 9 0 1 9 9 4 13 1 10 9 9 1 9 7 9 1 9 1 9 0 1 1 9 2
36 3 0 4 15 13 12 9 1 11 9 7 12 1 11 11 7 12 10 1 9 11 2 11 2 11 2 11 2 11 2 11 2 11 7 11 2
24 1 0 12 9 13 15 3 1 9 2 7 11 13 9 4 13 1 1 10 0 9 3 0 2
21 0 1 9 1 9 15 13 0 1 11 2 4 10 1 10 0 0 13 1 9 2
20 2 15 13 0 1 10 15 15 4 13 9 2 9 7 0 9 2 13 11 2
2 11 2
5 0 9 1 9 5
5 11 2 11 2 2
23 10 0 9 15 13 0 9 1 9 1 10 9 1 11 9 2 4 13 1 9 1 9 2
7 15 4 0 13 1 9 2
15 10 0 9 13 0 1 9 1 0 2 1 11 11 9 2
11 9 1 9 13 0 1 9 12 9 9 2
17 15 4 4 13 12 1 10 0 1 9 2 15 13 1 9 9 2
6 9 13 1 1 9 2
16 9 4 3 13 2 13 9 11 11 1 11 11 9 1 11 2
33 0 1 9 12 4 10 12 0 9 13 1 1 9 2 7 1 10 9 0 13 9 2 15 13 0 9 1 0 9 2 13 1 2
18 2 15 4 13 0 1 9 1 9 2 7 9 4 1 13 1 0 2
14 9 13 0 9 2 7 9 13 1 9 2 13 9 2
17 2 1 3 15 13 13 15 12 9 2 7 15 4 0 13 0 2
10 15 13 0 7 13 1 15 0 9 2
37 15 13 1 1 16 9 13 9 1 9 1 10 0 9 15 13 0 1 1 9 2 7 1 9 7 1 9 2 13 10 9 1 11 16 9 13 2
5 9 13 1 0 2
26 2 15 13 0 16 15 13 0 2 7 15 13 9 1 16 15 13 10 9 2 13 9 11 1 11 2
21 9 15 4 13 1 9 2 4 13 9 1 9 7 4 1 10 4 13 1 9 2
4 2 11 2 5
9 9 13 12 9 9 1 11 9 5
5 11 2 11 2 2
24 9 1 10 9 1 9 1 11 1 11 4 1 11 9 13 1 9 1 12 9 1 0 9 2
30 9 4 13 1 14 4 13 12 9 9 1 9 1 11 7 1 9 1 11 1 12 9 1 3 11 7 11 8 11 2
30 9 15 4 13 1 12 9 13 0 0 0 9 15 13 16 9 4 13 1 11 7 11 1 10 9 16 15 4 13 2
35 1 9 13 9 16 0 9 13 0 1 10 0 9 1 0 9 15 4 13 0 7 1 9 1 0 9 16 15 13 14 13 15 15 13 2
19 9 13 0 7 16 10 9 13 2 4 15 1 0 9 13 1 0 9 2
11 15 13 11 15 4 13 9 1 11 9 2
5 9 13 0 0 2
11 15 4 3 13 10 9 1 12 9 9 2
12 11 13 10 9 1 16 9 3 4 13 9 2
18 3 13 15 16 10 9 13 9 1 0 9 2 15 9 3 13 1 2
4 2 11 2 2
5 9 13 11 11 5
6 11 11 2 11 2 2
29 11 11 13 0 7 13 0 1 9 1 9 9 1 9 1 11 11 9 2 7 10 9 3 1 9 13 1 15 2
15 11 13 1 10 0 9 2 7 15 13 15 0 1 9 2
28 15 13 0 7 13 0 9 2 3 1 16 10 9 1 10 0 9 13 16 9 4 3 13 16 9 4 13 2
36 1 16 15 13 1 9 3 13 3 11 10 9 2 7 13 1 10 0 1 14 13 10 9 2 7 9 13 1 1 10 0 9 3 1 9 2
34 9 13 1 15 2 7 3 13 15 10 9 1 11 2 15 13 10 9 9 1 14 13 1 1 9 1 3 0 9 1 10 9 9 2
17 2 15 13 0 0 0 1 9 10 2 7 3 4 15 13 0 2
53 16 15 13 1 9 1 9 7 13 16 15 13 3 0 1 10 3 0 2 13 15 0 1 1 14 13 10 0 9 1 9 1 9 2 7 1 10 10 9 13 15 1 9 2 13 11 11 1 10 9 1 9 2
4 2 11 2 5
5 10 9 1 11 5
3 0 9 5
3 0 9 5
4 13 10 9 5
18 11 11 11 13 3 9 1 10 0 0 9 1 9 1 9 1 11 2
12 7 15 13 0 0 1 3 9 4 13 15 2
21 11 11 11 4 13 12 1 10 1 15 12 0 0 0 0 9 1 9 1 9 2
10 7 10 0 9 13 15 3 9 1 2
12 11 13 0 0 1 9 10 0 9 13 1 2
4 9 2 11 5
7 2 15 4 13 10 9 2
10 15 13 12 0 1 10 9 1 11 2
6 12 9 7 12 10 2
14 1 11 13 15 15 1 11 1 9 15 13 3 1 2
19 7 10 1 10 13 15 3 1 9 2 3 3 0 2 13 9 1 11 2
17 3 13 15 3 1 9 1 10 9 15 1 11 11 13 12 9 2
15 3 13 15 3 1 12 10 1 11 9 7 9 1 9 2
11 9 1 10 12 9 13 1 3 12 9 2
9 11 11 13 15 15 13 1 9 2
5 7 3 13 9 2
8 2 15 13 3 0 1 9 2
14 15 13 0 9 1 9 2 13 11 1 9 1 11 2
12 15 13 16 15 13 10 0 0 9 1 9 2
28 16 15 3 13 1 1 11 13 15 15 16 9 1 9 13 0 0 1 1 10 9 1 10 0 9 1 9 2
14 3 13 15 15 1 14 13 9 1 14 13 1 9 2
32 2 1 10 0 3 13 15 1 9 0 1 9 1 9 1 11 2 7 15 13 15 13 0 14 13 3 15 13 15 1 11 2
23 1 10 0 13 15 9 1 10 9 7 15 13 1 1 10 0 9 1 9 2 13 11 2
27 2 15 13 1 9 1 10 9 7 13 1 10 0 12 2 2 13 11 11 11 1 10 9 1 11 11 2
16 0 12 13 10 12 9 9 2 9 2 9 2 9 7 9 2
8 2 6 2 15 13 3 12 2
10 9 13 15 3 9 1 2 13 11 2
27 10 12 15 3 1 11 13 1 1 9 13 11 11 11 7 11 11 11 7 11 11 11 2 15 13 9 2
11 1 9 13 10 12 9 9 1 1 11 2
36 2 1 9 16 9 13 13 15 10 9 1 9 15 13 1 9 7 13 3 0 15 13 1 14 13 16 15 3 4 13 1 9 9 1 9 2
21 0 13 15 3 0 9 15 13 3 16 15 13 3 0 14 13 1 9 1 15 2
10 15 13 10 9 3 0 13 10 9 2
13 15 4 13 10 9 14 13 15 1 2 13 11 2
20 11 13 10 12 9 1 11 15 3 13 1 10 0 9 1 9 1 0 9 2
5 11 13 1 9 5
13 11 11 11 13 1 1 9 1 9 1 11 9 2
8 3 13 11 1 10 0 9 2
9 11 11 11 9 13 9 1 11 2
5 9 13 11 11 2
4 9 2 11 5
9 2 15 13 9 1 0 7 9 2
11 15 4 15 13 15 15 13 1 14 13 2
6 15 13 10 0 9 2
8 11 13 9 1 3 10 9 2
10 15 13 3 3 9 15 13 10 9 2
19 11 4 3 13 0 0 7 0 16 15 13 7 13 7 15 13 0 9 2
12 15 4 13 0 1 15 1 9 2 13 11 2
7 13 9 0 3 9 12 5
10 10 9 13 3 0 1 15 1 11 2
9 12 2 13 14 13 9 3 9 2
11 12 2 13 10 0 9 1 9 1 9 2
9 12 2 13 10 9 1 0 9 2
10 12 2 4 3 13 9 11 1 9 2
15 10 2 9 2 2 11 11 4 13 16 10 9 13 0 2
17 11 9 2 12 1 10 9 2 4 13 0 0 1 11 3 0 2
22 1 9 13 15 1 15 11 4 13 1 1 12 9 7 13 9 1 9 2 1 9 2
17 9 1 11 2 11 11 11 2 13 3 9 1 11 13 3 0 2
18 2 15 13 1 1 10 9 15 13 1 7 15 13 1 0 1 15 2
10 15 13 0 1 1 11 2 13 11 2
4 11 13 0 2
16 2 15 13 0 0 9 7 13 0 9 7 0 9 1 9 2
9 15 4 3 13 10 1 0 3 2
12 11 13 9 3 0 1 9 2 1 12 9 2
17 12 2 1 12 0 2 9 4 13 1 1 1 0 9 1 9 2
3 9 9 2
21 11 2 11 2 12 2 2 11 2 11 2 12 2 2 11 2 11 2 12 2 2
4 2 11 2 5
6 11 1 9 1 11 5
5 11 2 11 2 2
8 11 11 13 14 13 1 9 2
13 9 13 3 12 9 1 9 1 9 9 1 11 2
9 11 11 13 10 0 9 1 9 2
22 11 13 1 9 1 9 2 7 13 15 1 11 11 1 10 9 1 12 9 1 9 2
11 1 12 9 13 15 0 9 1 1 9 2
7 11 13 3 1 12 9 2
23 9 13 0 1 0 9 2 7 1 12 9 1 0 9 13 15 3 0 15 13 1 9 2
20 12 9 13 1 1 9 11 11 1 11 2 15 3 13 3 12 9 1 11 2
13 11 11 13 1 9 1 9 1 12 9 1 9 2
8 15 13 12 9 1 11 11 2
10 11 11 11 13 0 3 1 0 9 2
8 9 13 9 12 1 11 9 2
16 11 11 4 13 15 1 12 9 1 12 9 7 3 12 9 2
4 2 11 2 5
8 9 13 12 9 9 1 11 5
5 11 2 11 2 2
21 1 12 9 9 13 1 9 1 14 13 0 1 9 1 0 9 1 11 1 11 2
26 3 0 0 13 9 1 11 2 16 1 9 1 9 9 13 14 3 13 3 9 2 1 11 9 11 2
42 11 4 13 9 1 14 13 1 12 9 9 2 12 9 9 2 1 14 13 9 1 9 7 9 1 10 0 9 1 11 2 15 10 0 9 4 4 13 1 0 9 2
8 2 9 13 0 0 1 9 2
26 15 13 3 0 1 14 13 1 9 2 7 9 1 9 13 16 15 13 0 2 13 11 11 1 11 2
16 15 13 15 3 13 0 14 13 16 10 9 13 10 0 9 2
12 3 11 13 16 9 1 11 3 13 0 0 2
43 2 9 7 10 9 13 9 7 13 9 1 11 2 7 9 13 0 1 9 1 9 1 14 13 1 9 15 1 0 9 4 13 0 0 2 13 11 11 1 11 1 11 2
4 2 11 2 5
4 9 1 9 5
11 11 5 11 2 11 2 11 11 11 2 2
23 11 7 10 0 9 13 9 1 10 0 9 11 2 11 7 11 1 9 1 9 1 11 2
22 9 4 1 9 13 9 9 2 7 10 0 13 1 16 9 4 13 1 0 1 9 2
20 3 12 9 7 11 13 9 1 10 0 9 1 9 1 10 0 9 1 11 2
19 9 13 7 10 0 9 7 0 0 9 2 15 13 10 0 0 1 9 2
25 9 13 1 10 0 9 1 0 9 1 9 7 10 2 0 9 7 9 1 10 0 0 9 2 2
21 3 10 0 9 11 7 11 13 15 9 1 9 2 13 11 9 11 11 1 11 2
19 7 15 13 10 9 1 11 1 16 10 0 9 13 1 2 13 15 1 2
35 2 9 1 10 0 0 9 7 9 13 0 9 7 4 3 13 9 1 10 0 9 1 10 9 2 13 9 7 9 11 11 2 11 2 2
4 2 11 2 5
7 11 11 13 1 1 9 5
5 11 2 11 2 2
9 9 13 9 1 9 11 11 9 2
14 11 13 1 10 9 3 15 13 9 1 10 0 9 2
15 1 0 9 13 0 11 9 1 10 0 9 2 13 11 2
31 7 16 11 13 11 0 9 2 4 10 0 9 13 0 9 1 15 2 0 9 3 3 1 9 4 13 15 1 9 10 2
25 0 13 11 0 9 2 7 1 9 1 9 13 9 0 1 0 9 7 9 2 13 10 0 9 2
36 9 11 11 11 13 9 10 1 10 9 1 10 10 9 2 16 9 11 11 3 13 10 0 9 0 1 10 9 1 10 0 9 1 11 9 2
10 10 9 11 11 4 13 15 1 9 2
31 9 2 15 3 13 9 1 10 0 2 0 9 2 4 13 16 11 9 14 13 1 13 2 10 9 1 10 0 9 2 2
15 1 10 9 1 9 11 8 11 9 9 2 13 11 9 2
16 2 15 13 1 11 16 15 13 12 16 10 9 13 10 9 2
8 15 4 13 3 1 12 9 2
32 9 10 13 10 9 1 10 0 9 9 7 10 0 9 2 13 9 1 9 2 15 13 12 9 1 9 1 16 15 4 13 2
4 2 11 2 5
10 9 13 1 9 1 9 1 11 11 5
5 11 2 11 2 2
18 9 13 3 1 9 1 3 10 9 4 13 7 13 1 9 11 11 2
11 9 4 0 13 10 10 9 2 1 9 2
13 9 13 1 12 9 1 10 0 9 1 11 9 2
18 12 9 4 13 7 12 13 16 9 2 10 9 2 13 10 10 9 2
5 9 13 9 3 2
27 10 9 2 15 13 1 9 1 9 2 4 13 7 13 1 10 9 1 9 16 15 13 10 9 1 9 2
12 0 4 10 9 13 1 10 9 12 9 1 2
11 15 4 13 1 10 10 9 2 1 9 2
24 9 13 9 16 9 0 4 13 1 9 15 4 13 15 10 2 7 9 10 4 3 3 13 2
26 9 13 3 3 9 1 9 2 7 15 4 3 4 13 10 9 1 9 11 11 11 2 15 4 13 2
4 2 11 2 5
7 13 9 1 0 0 9 5
24 11 11 11 13 1 1 12 7 13 1 0 9 1 9 1 12 9 9 1 9 1 9 9 2
17 9 1 11 11 11 13 10 9 1 10 0 9 2 1 12 9 2
13 10 9 13 3 1 9 1 9 1 11 1 9 2
4 9 2 11 5
21 9 13 9 1 11 1 11 0 1 9 2 16 15 13 9 1 10 9 1 9 2
25 9 1 11 9 13 10 9 1 10 0 9 2 0 1 11 11 1 11 1 12 2 1 12 9 2
7 2 15 13 10 0 9 2
11 15 13 9 1 9 7 1 9 7 9 2
14 10 9 13 0 0 2 13 9 11 11 11 1 9 2
31 11 11 13 1 9 12 3 1 9 2 7 13 0 1 0 9 7 13 0 12 0 9 1 9 11 11 1 11 1 9 2
12 0 11 11 4 13 1 9 1 9 1 12 2
16 15 13 0 1 9 7 13 9 1 11 11 1 11 1 11 2
15 0 0 13 9 9 1 9 1 16 15 13 10 0 9 2
20 11 11 13 9 1 9 1 11 10 9 7 13 1 9 2 1 10 1 9 2
19 12 13 3 10 0 9 1 9 11 11 4 13 0 1 9 1 0 11 2
10 1 9 9 13 15 0 0 1 12 2
9 1 9 4 15 13 1 1 12 2
4 2 11 2 5
5 11 2 11 12 2
19 11 11 11 11 1 9 1 12 9 9 1 9 1 9 1 11 1 9 2
7 9 2 11 11 5 11 5
2 9 2
17 11 13 9 9 1 11 9 1 16 0 9 4 13 1 0 9 2
6 2 9 11 11 11 5
5 2 9 11 11 5
5 2 9 11 11 5
18 10 0 9 13 1 9 2 7 15 13 0 1 14 13 10 0 9 2
17 10 9 15 1 9 1 10 0 13 14 13 9 2 4 13 15 2
13 2 15 13 3 1 0 9 2 1 9 11 11 2
6 11 11 2 11 2 2
10 15 4 3 13 9 7 9 10 9 2
13 15 4 13 9 1 11 9 7 16 11 4 13 2
39 10 9 4 0 13 1 1 16 11 9 10 4 13 10 9 2 7 3 0 16 11 1 9 1 9 4 13 15 13 10 9 15 13 1 9 7 9 9 2
38 15 15 15 4 13 0 14 4 13 1 9 7 9 2 13 16 15 15 13 1 11 2 13 0 2 16 15 13 0 0 9 1 3 10 9 4 13 2
6 1 11 13 15 0 2
19 2 11 4 3 13 10 0 9 1 0 9 7 13 10 0 0 9 2 2
4 2 15 13 2
7 2 10 0 0 9 2 2
24 1 15 15 13 1 15 11 10 9 3 4 13 2 13 15 0 1 16 15 3 0 4 13 2
7 10 9 13 3 0 0 2
21 13 15 16 11 0 0 9 1 10 9 13 0 2 7 13 15 3 9 1 9 2
4 9 11 11 2
26 16 9 11 4 13 1 2 7 15 15 13 1 11 2 13 11 9 16 11 4 13 10 0 0 9 2
28 15 13 10 9 15 11 4 13 1 11 1 0 9 0 2 7 15 13 11 9 16 11 0 13 10 10 9 2
8 15 4 11 3 0 3 13 2
29 7 15 13 0 16 15 4 13 10 9 1 10 0 9 1 11 7 3 1 10 0 9 1 10 0 9 1 9 2
6 11 11 2 11 2 2
10 15 13 3 0 0 14 13 0 1 2
66 15 13 3 0 16 15 4 13 9 2 7 1 10 9 2 15 13 10 1 10 3 0 9 1 10 0 2 4 15 13 2 9 9 7 3 0 9 1 10 0 9 1 0 9 2 13 15 3 1 10 9 3 1 0 0 16 15 13 9 1 14 13 10 10 9 2
33 16 15 13 2 0 13 1 2 14 13 9 1 11 1 14 4 13 15 1 9 2 13 15 10 0 7 1 10 9 10 0 9 2
33 3 13 15 9 3 3 16 15 3 3 1 9 4 13 16 15 4 13 15 2 7 15 13 16 15 13 0 1 16 15 4 13 2
10 7 3 13 10 9 1 9 7 9 2
74 13 15 10 9 1 10 9 15 13 1 11 7 9 1 9 1 16 11 3 4 13 10 0 9 2 7 13 15 16 15 4 13 11 10 9 16 15 16 15 13 10 3 0 9 1 10 9 2 10 3 0 9 1 9 7 10 0 9 2 1 0 4 13 1 1 2 4 15 13 2 14 13 9 2
4 9 11 11 2
34 15 4 13 11 9 1 1 9 2 7 4 3 13 1 16 15 13 10 9 1 9 1 11 2 7 10 9 4 4 13 10 9 1 2
20 1 10 9 4 11 2 0 1 9 1 9 2 13 1 10 9 1 10 9 2
19 15 4 13 9 7 1 7 1 10 9 1 7 10 9 1 9 1 11 2
23 15 9 11 13 16 15 13 9 1 10 9 7 10 9 2 13 3 10 0 0 0 9 2
14 15 13 0 1 16 0 9 9 13 10 9 1 9 2
38 9 13 16 15 3 13 10 0 9 1 14 13 0 9 1 9 1 10 9 2 3 0 13 1 10 9 16 15 1 9 13 1 10 9 1 0 9 2
19 15 13 16 9 4 13 10 0 9 1 14 13 15 15 13 9 1 9 2
4 3 13 9 2
25 4 15 13 9 1 10 9 16 15 13 10 3 0 9 1 9 1 15 9 11 3 13 1 1 2
7 11 11 11 2 11 2 2
25 11 13 3 0 0 1 16 9 3 13 0 9 1 14 13 1 9 15 4 13 1 0 0 9 2
14 15 13 10 0 9 1 9 1 15 9 0 4 13 2
29 15 13 0 10 9 15 4 13 16 15 13 0 1 3 0 9 16 15 4 4 13 0 2 0 9 2 1 9 2
7 15 13 15 13 3 0 2
16 7 16 9 3 13 11 0 9 2 13 15 0 0 1 15 2
25 1 0 9 2 1 11 7 11 2 4 15 13 0 0 16 10 0 9 4 13 0 1 1 9 2
30 15 4 4 13 1 16 15 14 13 3 1 0 0 9 4 13 0 3 1 14 4 13 1 10 0 9 1 10 9 2
8 13 9 0 1 10 10 9 2
4 9 11 11 2
29 9 1 9 1 0 9 7 10 9 1 15 1 10 9 15 13 2 15 13 15 1 9 11 1 9 1 9 9 2
23 15 13 9 16 3 9 11 10 9 13 15 7 3 1 9 13 1 15 1 10 0 9 2
9 15 4 3 13 1 0 9 3 2
25 15 13 16 15 4 13 0 1 10 9 15 4 4 13 1 0 1 9 1 10 0 9 7 9 2
28 15 4 13 16 15 13 9 1 15 14 13 10 0 2 0 9 7 15 14 13 1 10 0 9 0 1 9 2
13 15 13 1 10 9 16 15 4 13 1 10 9 2
24 15 13 3 0 1 9 2 7 9 13 9 15 13 0 1 10 9 15 1 9 13 1 9 2
20 13 15 1 10 9 15 13 9 2 3 9 2 4 9 13 1 10 10 9 2
22 3 4 15 13 15 16 15 1 9 7 1 9 13 0 9 16 15 13 9 1 15 2
6 11 11 2 11 2 2
9 10 9 13 3 1 9 7 9 2
52 16 0 3 4 13 1 1 2 4 15 0 9 13 1 11 10 9 1 11 11 2 3 15 13 16 15 13 7 0 7 0 0 14 13 9 1 11 15 3 13 2 7 15 4 13 10 9 1 9 1 11 2
31 1 10 9 9 13 15 1 9 16 15 13 1 10 9 2 7 16 15 4 13 1 0 9 1 14 13 0 9 1 11 2
36 15 4 0 13 0 0 0 9 15 4 13 0 0 9 2 7 15 4 10 13 15 1 0 16 15 4 13 3 0 7 14 13 7 14 13 2
12 13 15 0 3 16 9 13 9 1 10 9 2
25 4 11 13 1 9 1 9 15 13 9 1 9 2 1 14 13 1 16 15 4 13 1 10 9 2
4 9 11 11 2
20 15 4 13 15 10 9 15 4 13 1 9 2 1 12 1 0 9 1 9 2
31 15 4 3 13 9 1 14 13 1 9 1 1 10 9 2 7 15 13 3 10 9 1 14 13 16 15 13 15 1 9 2
34 7 15 13 15 13 0 16 15 13 0 9 1 10 9 2 7 3 0 16 15 13 0 0 9 1 15 15 3 4 13 1 10 9 2
6 15 13 15 13 0 2
20 15 13 3 16 9 1 10 0 9 4 13 0 7 0 0 16 15 4 13 2
33 16 15 13 9 1 9 1 0 9 2 13 15 10 9 16 15 4 13 0 14 13 10 0 9 1 16 10 0 9 13 1 9 2
18 15 4 13 16 15 13 0 0 9 1 9 1 3 0 15 4 13 2
36 10 9 4 1 9 13 16 15 13 9 1 14 13 10 10 9 1 9 2 7 15 13 0 9 15 13 1 1 14 13 9 15 4 13 9 2
19 15 13 11 9 2 11 2 15 15 13 1 9 1 9 2 7 3 11 2
6 11 11 2 11 2 2
6 15 13 9 1 9 2
21 15 15 15 13 1 2 13 0 0 9 1 11 10 9 1 11 9 10 0 9 2
35 3 13 15 3 1 16 9 13 9 1 0 9 2 15 3 4 13 0 2 7 15 13 3 0 1 16 10 0 9 3 13 9 1 9 2
38 4 15 3 13 0 14 13 1 9 1 14 13 9 1 0 1 9 1 10 3 0 9 2 1 3 14 13 15 1 10 0 9 16 15 4 13 0 2
4 9 11 11 2
10 15 13 0 16 1 9 13 15 9 2
41 15 13 9 1 16 15 13 0 1 10 9 2 3 0 15 15 4 13 1 14 13 0 9 2 7 16 9 1 10 9 15 13 2 13 1 9 1 14 13 15 2
9 3 13 13 15 9 1 9 1 2
17 15 13 16 15 13 0 1 10 0 9 14 13 1 10 0 9 2
26 15 13 3 1 10 9 16 15 14 13 0 9 3 4 13 1 14 13 15 14 13 1 9 0 9 2
28 15 4 13 15 16 11 2 15 3 13 10 1 15 15 13 1 0 9 2 13 9 1 10 10 1 9 9 2
2 9 2
7 15 13 9 2 11 11 2
6 11 11 2 11 2 2
9 1 10 9 13 11 10 0 9 2
15 10 1 9 1 9 13 16 9 0 9 4 13 1 12 2
32 9 9 1 14 13 9 1 9 1 11 13 0 10 9 16 15 0 13 9 1 11 1 9 2 3 15 1 4 13 1 9 2
16 1 3 1 9 15 13 9 13 1 9 2 13 9 10 10 2
20 1 11 13 1 10 9 9 13 1 9 9 2 16 9 13 1 11 13 9 2
7 4 9 13 9 1 15 2
4 9 11 11 2
24 15 4 1 10 0 13 15 10 9 16 11 4 13 10 1 3 9 1 9 16 15 13 9 2
16 3 1 0 10 9 3 13 15 1 1 11 10 9 1 9 2
25 15 4 11 13 0 0 1 1 0 9 2 7 15 4 3 13 1 10 0 13 1 9 1 15 2
24 15 4 3 1 0 9 13 11 9 16 15 13 9 1 9 2 7 11 9 1 15 1 9 2
24 15 13 16 15 15 4 13 1 10 9 2 4 13 0 7 4 13 1 11 9 1 0 3 2
53 3 16 15 13 0 1 16 15 13 9 0 2 7 16 15 13 9 15 13 1 9 1 10 9 2 13 15 16 11 4 13 10 10 9 16 15 13 10 9 15 13 14 13 1 0 9 1 9 1 10 10 9 2
26 16 15 3 13 15 2 4 15 1 9 13 3 10 10 16 11 13 9 2 9 2 9 7 0 9 2
2 9 2
6 11 11 2 1 9 2
2 9 2
8 15 13 3 0 1 10 9 2
7 11 11 11 2 11 2 2
12 15 13 0 1 16 9 11 3 4 13 3 2
16 1 0 9 4 11 13 9 1 9 1 9 1 9 1 11 2
44 1 0 1 15 13 15 10 0 9 16 15 1 11 1 10 9 7 9 4 13 9 2 1 3 14 13 9 7 1 0 9 7 1 9 1 10 9 15 13 0 9 1 9 2
6 15 13 10 0 9 2
6 15 13 0 0 9 2
25 1 0 9 4 15 13 16 9 4 13 10 9 1 9 1 10 9 15 9 13 1 9 1 10 2
15 15 13 0 9 16 0 9 4 13 0 9 1 10 9 2
27 1 10 9 13 9 11 11 10 9 15 13 1 9 1 10 9 2 9 13 2 11 4 13 1 1 11 2
19 15 4 13 9 10 0 9 1 14 13 11 2 9 13 2 9 1 9 2
18 13 15 10 0 9 1 11 1 10 9 1 14 13 11 9 1 0 2
2 9 2
13 9 13 9 11 1 14 13 15 1 10 0 9 2
14 15 13 10 9 15 13 3 0 9 15 13 1 9 2
9 15 13 12 9 15 13 15 1 2
4 11 11 11 2
5 15 4 13 15 2
4 9 11 11 2
29 15 13 9 11 9 1 16 15 1 11 4 13 1 9 9 1 0 9 2 1 9 2 9 7 3 3 1 9 2
15 15 13 0 1 16 15 13 10 0 9 15 3 13 1 2
29 15 15 13 1 9 2 13 3 16 15 4 13 9 1 9 1 11 2 7 1 10 9 4 15 13 9 1 9 2
24 9 13 1 10 9 16 16 15 4 13 9 1 9 1 11 2 4 15 13 1 10 0 9 2
12 3 4 15 13 9 15 13 10 0 0 9 2
20 15 13 1 11 9 10 0 9 15 15 4 13 2 0 1 9 1 10 9 2
43 16 15 13 9 1 11 9 7 0 9 0 1 11 2 13 15 10 9 1 14 4 13 15 1 15 11 4 13 1 10 9 2 7 3 3 16 15 13 9 9 1 15 2
16 11 4 3 2 15 9 11 13 1 2 0 3 13 10 9 2
7 11 11 11 2 11 2 2
26 15 13 3 3 10 9 1 9 2 15 13 0 15 4 13 0 10 0 9 1 9 16 15 13 15 2
17 15 13 0 1 16 0 9 1 11 4 13 1 0 9 10 9 2
5 15 13 0 9 2
9 7 15 13 3 10 9 1 3 2
15 15 13 3 10 0 9 2 15 13 3 1 9 1 9 2
27 15 4 13 9 1 3 12 9 2 7 15 9 13 2 13 16 15 4 13 14 13 15 1 12 9 1 2
10 15 13 0 9 2 7 15 13 9 2
35 16 11 4 13 15 1 9 2 16 15 4 13 1 0 9 2 7 16 15 4 13 1 9 2 13 15 0 1 14 13 10 0 9 3 2
22 13 9 14 13 16 11 13 10 0 9 1 11 1 10 0 9 15 4 13 1 9 2
4 9 11 11 2
32 13 15 3 4 13 16 11 13 9 1 3 10 10 9 15 15 0 4 13 9 1 0 7 1 11 16 15 13 9 1 9 2
10 15 4 15 3 13 1 11 1 9 2
15 15 13 10 9 1 1 10 9 15 4 13 1 9 9 2
30 10 0 9 1 15 13 16 15 3 4 13 15 1 9 1 9 16 15 13 10 9 1 9 15 13 10 0 0 9 2
21 9 4 2 1 9 1 11 9 2 13 1 3 14 13 1 9 1 10 0 9 2
14 15 13 15 13 16 15 13 9 1 11 1 14 13 2
41 16 10 9 13 1 9 2 16 15 13 15 15 13 9 1 9 2 16 15 13 10 9 15 13 0 1 15 2 16 15 13 3 0 9 13 2 3 13 15 0 2
34 15 9 11 3 13 1 2 13 9 1 1 9 7 1 16 10 0 9 13 1 9 2 7 2 9 13 2 0 10 0 9 4 13 2
23 15 13 3 10 0 9 2 9 13 2 1 9 1 10 0 9 9 11 13 15 13 1 2
2 9 2
11 7 15 2 9 2 13 10 9 1 9 2
7 15 13 3 1 10 9 2
7 1 9 11 11 1 9 2
27 2 15 13 0 0 16 10 0 9 13 0 9 2 9 2 9 7 10 0 9 1 14 13 10 0 9 2
43 13 15 0 16 9 3 13 0 1 15 2 7 3 13 15 3 10 9 1 11 7 9 2 15 13 1 9 10 0 9 2 2 3 15 4 13 1 11 0 9 12 2 2
6 11 11 2 11 2 2
13 15 13 1 9 2 15 15 0 3 13 0 1 2
28 15 4 13 16 16 9 13 1 0 9 16 15 13 1 9 1 9 1 9 2 3 13 15 12 0 0 9 2
14 1 10 9 13 15 0 1 9 2 3 0 0 9 2
6 7 15 13 0 9 2
32 2 1 1 1 10 0 9 1 0 9 1 9 4 15 1 9 12 2 12 13 1 12 13 3 12 12 9 1 0 9 2 2
24 15 4 0 13 1 0 9 15 4 13 2 7 16 15 3 13 1 9 2 15 9 3 13 2
7 15 13 15 13 1 9 2
13 2 9 13 2 2 7 15 13 0 9 1 9 2
33 4 15 1 0 9 13 1 2 9 13 3 2 16 15 13 10 0 9 2 7 16 15 1 9 13 1 1 10 9 15 13 0 2
4 9 11 11 2
20 15 13 1 1 16 11 13 14 13 9 1 9 1 9 2 7 3 1 9 2
10 15 13 1 1 16 15 13 10 9 2
25 15 15 13 9 1 9 10 0 9 2 13 15 10 9 13 1 16 15 4 13 10 9 1 9 2
34 7 15 13 15 3 10 9 1 2 15 13 0 0 1 3 3 0 9 15 4 13 2 7 15 13 0 1 16 15 13 10 0 9 2
36 16 15 13 2 15 13 16 15 4 4 13 0 16 15 13 15 15 13 0 2 3 0 9 2 15 3 3 13 0 0 9 2 7 3 9 2
24 7 1 10 15 9 4 13 0 1 9 1 12 2 4 0 9 1 10 9 13 0 7 0 2
14 7 15 4 13 15 15 4 13 1 10 9 1 9 2
25 15 13 1 10 9 10 0 9 12 16 15 1 9 4 13 16 0 9 1 12 4 13 12 12 2
5 2 9 13 2 2
10 2 4 15 4 13 10 9 2 9 2
21 2 3 4 9 13 2 15 13 0 7 13 16 15 4 13 12 12 9 1 12 2
15 1 15 13 12 12 0 0 9 2 7 12 12 0 9 2
6 11 11 2 11 2 2
15 15 13 3 1 9 2 15 15 0 3 3 13 0 1 2
22 15 4 3 13 16 15 13 16 9 1 10 9 13 1 10 0 9 15 15 13 1 2
16 1 11 13 15 10 0 9 1 11 1 0 12 9 0 9 2
15 1 9 15 13 12 9 2 13 15 12 9 15 13 9 2
15 1 9 15 13 12 9 2 13 15 12 9 15 13 9 2
12 15 13 3 1 1 10 0 0 9 1 11 2
6 13 9 15 13 0 2
22 7 16 15 3 13 15 2 15 4 15 13 1 16 15 0 4 13 10 9 1 15 2
4 9 11 11 2
27 15 13 16 11 10 9 2 1 10 0 9 2 3 13 0 1 10 0 13 1 10 9 15 13 1 9 2
30 16 15 4 13 11 11 2 4 15 3 13 16 15 4 13 10 9 15 4 13 0 2 16 15 13 9 15 13 9 2
37 7 15 13 3 9 0 9 15 13 11 9 10 9 2 15 13 3 9 1 16 15 4 13 10 9 1 9 1 11 1 9 1 1 9 1 11 2
12 7 15 13 15 16 15 13 10 0 9 1 2
6 11 11 2 11 2 2
14 15 4 13 16 15 13 10 0 0 1 9 1 9 2
5 15 13 0 9 2
12 2 9 4 1 9 13 1 0 9 1 9 2
25 1 9 13 9 16 9 3 13 9 0 16 15 1 10 13 0 7 0 10 0 9 1 0 9 2
7 15 4 9 3 0 13 2
31 15 4 3 0 13 16 15 13 3 0 9 1 9 1 9 7 9 2 7 4 3 13 9 1 9 1 12 9 1 9 2
11 3 4 9 13 9 1 9 1 9 2 2
4 9 11 11 2
11 9 9 4 1 10 9 13 1 0 9 2
14 15 13 1 0 1 16 0 9 13 1 9 0 0 2
31 15 4 0 13 1 16 15 13 0 0 2 7 16 15 7 4 13 1 10 0 0 9 1 9 2 7 16 9 4 13 2
8 9 1 9 13 3 0 9 2
28 1 10 4 15 7 13 3 9 1 3 12 9 9 4 13 1 2 7 3 15 4 13 10 0 9 1 9 2
18 1 1 1 9 9 13 15 1 10 0 9 1 9 1 10 0 9 2
20 1 12 4 3 10 9 1 9 13 1 10 12 9 1 9 1 10 0 9 2
20 10 9 13 16 9 1 9 4 13 1 9 1 9 1 9 1 9 7 9 2
15 10 10 9 4 13 0 9 1 11 7 4 13 10 9 2
15 15 4 1 9 1 9 13 1 12 10 0 9 1 11 2
10 10 9 1 9 7 10 9 1 9 2
13 10 9 13 0 7 4 13 10 0 9 1 9 2
25 15 4 3 3 3 13 16 3 9 1 9 1 9 7 10 0 9 1 9 4 13 1 10 9 2
28 15 13 3 10 0 9 1 3 0 16 15 4 13 1 9 1 14 13 15 1 1 11 3 0 1 0 0 2
6 11 11 2 11 2 2
22 3 4 15 13 16 15 13 0 1 16 9 13 16 15 13 16 9 3 13 9 0 2
23 16 15 13 9 1 14 13 10 9 1 9 1 9 1 9 1 9 2 13 15 9 1 2
66 16 9 3 13 16 15 13 1 14 13 10 9 1 9 7 1 9 1 9 2 13 15 16 9 3 3 4 13 1 15 15 3 4 13 2 3 10 9 16 15 13 0 9 2 10 9 1 9 2 3 15 4 4 13 0 3 14 13 1 1 15 15 13 1 9 2
23 4 9 13 15 1 16 9 16 15 13 0 9 13 2 7 16 9 3 3 4 4 13 2
4 9 11 11 2
17 15 13 0 16 15 1 11 13 1 9 1 10 9 1 0 9 2
41 15 4 0 13 9 1 2 7 15 13 16 15 4 13 0 0 2 16 10 9 4 13 1 10 9 3 1 9 2 3 16 11 4 13 9 7 13 10 9 3 2
44 15 4 3 0 13 1 9 2 7 15 13 1 10 10 9 0 3 1 14 13 16 15 3 4 13 16 15 4 13 2 0 7 0 16 9 1 11 4 13 1 10 0 9 2
35 13 15 0 2 13 15 3 10 9 14 4 13 15 3 1 9 2 7 1 10 9 4 15 3 4 13 0 9 1 10 9 1 3 0 2
24 16 15 13 1 10 0 9 2 3 4 10 0 9 4 13 1 1 11 3 0 1 0 0 2
16 15 4 13 0 16 3 9 9 4 13 1 9 1 10 9 2
6 11 11 2 11 2 2
6 15 13 3 1 9 2
42 15 13 15 13 0 16 9 13 16 15 1 9 13 1 9 9 2 16 15 3 3 13 15 15 9 13 1 2 7 16 15 4 13 10 9 1 10 9 1 0 9 2
17 16 15 13 1 9 1 9 7 1 9 2 13 0 1 1 9 2
8 3 0 15 13 2 3 0 2
31 10 9 13 15 0 14 13 1 9 1 0 9 16 15 1 9 13 9 0 0 2 7 15 13 0 10 9 9 13 1 2
38 16 15 4 13 9 2 4 15 3 13 1 12 9 2 10 9 1 16 15 3 4 13 0 1 12 9 1 9 1 9 7 9 2 7 13 10 0 2
28 1 9 13 15 0 15 0 13 0 1 9 1 10 12 9 2 15 4 3 13 1 9 0 1 1 12 9 2
4 9 11 11 2
37 16 9 4 13 2 13 15 1 10 9 16 15 4 13 9 14 13 10 0 9 1 2 3 16 9 13 15 0 0 7 0 16 15 13 1 9 2
12 16 15 13 2 4 0 12 9 3 13 9 2
34 15 4 3 1 0 13 16 15 13 12 9 13 0 3 15 13 1 9 2 7 15 4 1 10 9 3 13 16 15 4 13 9 3 2
13 16 9 3 4 13 2 13 12 9 3 0 0 2
14 3 13 15 3 0 10 9 7 13 15 3 1 0 2
6 11 11 2 11 2 2
16 2 9 4 13 16 11 13 1 9 1 10 9 1 9 9 2
17 9 1 9 13 3 0 16 10 9 1 12 9 13 0 1 9 2
28 1 11 4 15 3 13 14 13 9 3 16 9 13 16 15 13 2 7 3 13 15 3 14 13 1 0 9 2
26 10 9 4 11 13 1 9 1 9 15 13 0 1 15 15 13 1 10 9 2 1 14 13 9 2 2
4 9 11 11 2
21 15 13 0 0 9 1 16 9 13 14 13 0 9 1 10 9 1 10 0 9 2
22 9 13 16 10 0 4 13 9 1 9 9 2 7 4 3 13 1 0 9 7 9 2
12 10 9 4 3 13 1 14 13 15 0 9 2
28 0 1 9 1 9 15 13 0 9 2 7 3 9 1 9 13 0 2 4 15 13 0 14 13 9 1 9 2
33 0 4 1 10 9 4 13 0 0 0 9 1 9 1 16 15 1 9 13 9 7 3 4 13 0 1 10 0 9 1 9 9 2
19 1 7 1 9 12 4 15 1 9 13 0 9 1 9 1 9 1 9 2
13 0 4 9 1 9 13 1 9 7 9 1 9 2
18 10 0 9 13 16 9 1 10 9 1 9 13 3 1 9 1 9 2
6 9 4 13 1 9 2
27 16 0 9 7 9 1 9 13 10 9 1 10 9 15 4 13 1 9 2 4 10 0 9 13 1 9 2
25 16 9 13 7 13 1 0 9 1 10 0 9 2 7 13 1 0 2 13 10 9 1 0 9 2
34 9 1 16 15 4 13 0 7 0 9 1 9 13 0 16 15 13 0 16 9 1 0 9 13 9 1 10 1 9 0 0 0 9 2
22 9 13 14 13 9 1 14 13 7 13 10 9 1 16 15 13 10 9 1 10 9 2
47 1 9 1 14 13 9 1 9 1 0 9 1 9 13 3 3 10 0 9 9 1 9 15 4 13 3 1 9 1 10 0 9 0 1 9 2 7 1 14 13 15 7 13 0 0 0 2
6 9 13 15 1 0 2
14 1 9 1 9 1 12 4 15 3 13 9 1 9 2
23 9 13 14 13 11 9 1 14 13 9 1 10 0 9 1 12 12 9 1 9 1 9 2
20 9 13 1 16 9 4 13 1 12 12 9 2 15 15 4 13 1 1 11 2
16 9 1 9 13 16 0 9 1 9 1 9 1 9 13 0 2
14 15 4 3 13 9 1 10 0 9 1 9 1 9 2
34 0 13 1 16 15 4 13 0 14 13 1 9 1 14 13 9 9 1 14 13 9 1 10 9 1 14 13 1 15 7 13 0 9 2
10 15 4 3 4 13 0 9 1 9 2
18 15 13 9 1 14 13 1 1 11 1 10 0 9 1 9 1 9 2
6 11 11 2 11 2 2
27 3 4 15 13 16 15 13 0 1 16 9 3 13 16 15 4 13 1 10 9 1 9 1 9 1 9 2
21 15 13 0 1 16 15 3 4 4 13 1 9 1 9 2 0 13 10 0 9 2
4 15 13 0 2
39 16 9 13 16 2 0 13 1 2 16 9 9 3 13 0 3 2 7 16 15 4 2 13 2 14 13 9 2 13 3 0 3 0 15 15 4 13 1 2
22 15 13 3 3 0 3 0 15 9 13 1 9 2 1 10 9 3 3 15 13 15 2
23 3 13 9 0 1 16 15 4 13 1 9 1 9 9 2 3 3 9 13 1 12 9 2
30 4 9 13 16 15 4 13 1 15 9 13 2 3 14 13 9 2 7 16 15 13 9 1 9 1 9 15 3 13 2
4 9 11 11 2
91 16 15 13 15 3 0 1 14 13 16 2 0 13 1 2 16 9 3 13 0 3 2 13 15 10 9 1 1 10 9 1 11 11 10 0 9 2 1 3 10 9 9 3 2 3 15 13 1 10 2 9 2 1 9 2 7 3 15 13 16 1 9 4 9 7 0 1 12 0 9 13 9 7 9 0 3 12 9 9 2 7 16 12 9 9 1 15 13 0 9 2
13 3 15 13 0 16 10 9 13 3 1 0 9 2
11 3 13 15 16 15 13 9 1 0 9 2
17 1 10 9 13 15 3 16 15 13 3 16 15 13 14 13 9 2
11 15 3 1 13 16 15 4 13 0 9 2
12 15 15 13 2 13 10 9 15 4 13 1 2
42 9 13 1 10 9 15 11 11 13 1 2 16 2 9 13 9 1 14 13 1 11 1 9 1 0 9 1 9 15 4 13 11 0 1 9 1 9 15 13 1 2 2
6 15 4 4 13 1 2
6 11 11 2 11 2 2
22 3 4 15 3 13 16 15 4 3 13 0 1 16 15 0 13 10 9 15 13 3 2
55 10 9 15 13 1 11 2 13 0 0 0 1 1 10 9 15 13 1 15 2 7 3 13 15 3 16 10 9 0 9 13 9 1 14 13 1 15 10 0 9 2 7 15 13 3 0 1 16 10 1 15 13 1 11 2
16 15 4 13 3 10 9 16 3 13 15 9 15 13 10 9 2
38 7 1 12 9 4 15 3 13 10 10 9 0 2 7 10 9 4 13 9 1 10 7 10 9 2 1 16 11 3 4 4 4 13 9 1 10 9 2
18 3 4 15 3 13 0 9 2 1 14 4 13 10 9 1 10 9 2
60 16 9 13 16 15 4 13 10 9 1 9 1 9 1 9 2 7 16 15 13 0 1 15 9 13 2 16 15 4 13 0 1 9 1 10 9 2 4 15 3 13 9 1 10 9 3 15 0 13 15 2 15 4 13 0 9 1 11 9 2
4 9 11 11 2
47 15 13 0 1 9 11 11 1 16 15 4 13 1 16 15 13 9 1 11 3 16 15 13 9 2 15 13 16 15 13 0 2 7 16 0 9 4 13 15 9 1 9 1 9 1 9 2
6 3 13 15 3 9 2
44 15 13 3 3 7 9 7 0 1 9 4 13 1 9 5 9 16 15 4 13 9 1 0 9 1 9 2 3 16 15 3 13 0 1 3 12 9 16 15 13 10 0 9 2
21 0 15 9 15 13 1 9 2 4 13 1 1 2 4 15 3 13 3 7 3 2
32 7 15 13 0 2 15 15 13 2 16 15 13 14 13 1 15 9 13 1 10 9 1 9 2 15 15 13 1 10 10 9 2
2 9 2
16 11 13 9 9 1 11 9 1 16 0 4 13 1 0 9 2
14 2 9 11 11 11 2 9 11 11 2 9 11 11 5
18 10 0 9 13 1 9 2 7 15 13 0 1 14 13 10 0 9 2
17 10 9 15 1 9 1 10 0 13 14 13 9 2 4 13 15 2
12 2 15 13 1 0 9 2 1 9 11 11 2
6 11 11 2 11 2 2
21 15 4 13 10 9 13 15 4 13 10 0 9 2 16 15 13 1 9 1 9 2
11 7 15 4 13 9 1 10 10 0 9 2
18 1 9 13 15 0 16 11 13 14 13 1 11 9 1 9 1 9 2
24 9 13 14 13 1 9 1 9 1 9 1 9 2 7 3 4 15 13 0 0 3 1 9 2
18 15 4 13 1 9 1 9 1 9 15 11 4 13 1 14 4 13 2
10 11 9 13 0 1 9 1 11 9 2
22 11 4 13 9 1 11 1 14 13 12 9 2 7 3 1 14 13 9 1 10 9 2
49 15 4 13 16 11 3 3 13 15 1 0 14 13 1 10 9 1 0 2 1 7 1 16 15 4 13 10 10 9 1 1 15 2 1 9 1 14 13 14 13 9 1 11 2 15 13 0 0 2
5 9 11 11 11 2
11 16 15 13 9 2 13 11 9 10 10 2
27 15 13 15 13 0 0 14 13 1 9 1 0 0 9 16 15 3 13 1 9 15 4 13 1 0 9 2
22 9 13 0 16 15 13 0 0 2 7 15 13 15 16 15 3 13 9 1 14 13 2
13 16 15 13 11 9 2 13 11 0 1 10 9 2
29 15 13 2 3 0 15 13 2 10 9 15 4 13 14 13 0 1 1 3 12 2 15 13 9 1 9 1 11 2
33 7 9 1 9 7 1 0 4 13 1 1 10 9 1 9 1 9 2 7 3 1 9 15 4 13 10 1 15 15 13 1 9 2
31 10 9 13 0 2 16 15 4 13 15 9 15 13 0 1 9 1 9 1 11 2 7 0 9 4 13 0 1 10 9 2
23 7 15 13 0 14 13 16 9 3 4 13 1 9 1 2 7 13 10 9 1 0 9 2
29 3 13 15 0 16 15 13 3 16 10 0 9 3 13 1 16 9 1 0 0 9 16 15 13 9 2 13 1 2
17 3 13 11 0 0 7 4 3 13 1 7 13 9 1 10 9 2
26 7 15 13 3 1 16 15 3 4 13 14 13 1 10 0 9 2 7 3 13 1 10 0 0 9 2
6 11 11 2 11 2 2
9 9 13 3 2 0 0 9 2 2
39 9 13 16 11 3 13 3 0 0 9 1 11 2 7 16 15 4 13 1 10 0 9 2 15 15 13 4 13 2 4 15 13 14 13 0 9 1 11 2
7 9 1 10 9 13 3 2
18 15 15 13 9 3 2 13 16 11 13 0 1 14 13 1 11 9 2
7 11 13 3 1 10 9 2
28 2 15 13 14 4 13 10 9 1 10 9 15 13 1 9 1 10 9 2 7 4 13 11 9 1 9 2 2
50 15 13 16 15 13 7 13 16 15 4 13 10 0 9 1 9 1 10 9 2 3 16 15 4 13 1 1 10 9 7 13 1 9 9 2 7 1 14 13 9 1 9 7 13 0 0 9 1 11 2
5 9 11 11 11 2
3 1 0 2
33 15 13 15 13 0 0 16 15 3 13 1 10 0 9 15 4 13 1 0 9 2 16 15 4 13 1 0 9 15 13 0 0 2
20 15 4 1 10 0 9 7 10 0 9 13 11 7 11 9 9 1 10 9 2
28 11 11 13 3 3 0 1 1 9 12 16 11 3 4 13 11 14 13 9 1 15 15 4 13 10 0 9 2
8 15 13 15 13 10 0 9 2
44 3 13 15 3 3 9 7 11 15 13 16 9 4 13 1 11 1 9 2 15 15 4 13 2 7 15 4 13 9 1 12 9 1 15 15 10 12 0 9 1 11 4 13 2
11 1 11 9 1 10 9 13 15 10 9 2
12 15 13 0 0 1 14 13 15 1 11 9 2
2 9 2
7 15 13 9 2 11 11 2
6 11 11 2 11 2 2
58 11 4 3 13 14 13 1 1 10 9 16 15 13 9 1 9 1 9 2 7 15 13 16 10 9 15 4 13 2 13 1 0 9 7 3 0 9 2 7 15 13 1 1 16 15 3 13 1 14 13 0 9 1 0 0 0 9 2
19 15 13 1 14 13 1 9 1 9 1 9 1 11 15 13 14 13 9 2
24 3 13 15 3 16 15 13 0 1 9 1 9 1 0 0 9 1 15 11 4 13 1 1 2
45 7 15 11 0 3 13 2 13 16 16 15 13 7 1 10 0 9 7 1 0 9 2 13 15 0 0 1 10 9 15 15 13 1 10 3 0 9 2 0 1 1 0 0 9 2
66 10 9 1 9 13 16 15 4 13 15 14 13 9 15 11 4 13 2 3 16 15 4 13 1 9 1 14 13 0 9 1 11 1 9 1 14 13 9 2 7 1 10 9 13 1 0 1 10 0 0 9 2 0 16 11 13 1 1 15 1 9 7 9 1 11 2
5 9 11 11 11 2
48 1 10 0 13 15 3 0 1 9 2 16 16 15 13 9 15 13 0 0 2 1 14 13 9 2 15 4 13 14 13 10 0 0 9 2 3 4 15 1 15 10 13 1 10 0 0 9 2
37 15 13 3 1 16 16 15 13 15 1 1 10 9 2 3 4 15 1 10 9 13 0 1 10 9 15 15 4 13 1 14 13 1 0 0 9 2
15 15 13 16 15 13 0 0 9 15 3 13 1 0 9 2
32 16 15 13 9 1 10 0 2 3 0 0 9 2 13 15 16 9 1 14 13 1 0 0 9 15 13 0 2 4 13 0 2
8 7 15 13 10 9 1 15 2
51 15 13 2 1 0 2 16 15 16 15 4 13 3 0 15 11 11 3 13 9 1 2 13 0 1 15 9 9 13 1 9 1 9 2 16 11 3 4 13 11 14 13 9 1 15 15 4 13 0 9 2
2 9 2
7 11 11 11 2 1 9 2
7 11 11 11 2 11 2 2
19 9 13 0 1 16 15 13 0 1 0 9 2 16 15 13 10 0 9 2
26 1 11 1 1 9 13 15 16 9 13 3 2 7 16 15 13 0 9 1 9 1 9 1 0 9 2
30 9 13 3 16 9 1 10 9 15 13 0 2 7 15 15 3 4 13 10 1 3 0 1 2 13 16 15 13 0 2
7 15 13 3 10 0 9 2
11 15 13 9 1 14 13 10 9 1 9 2
40 13 15 11 9 16 15 3 4 13 9 1 0 9 1 14 13 1 10 0 0 9 1 0 9 2 15 15 3 13 0 9 1 2 7 15 3 0 13 0 2
9 13 15 15 15 0 13 11 9 2
13 14 13 9 1 9 1 9 1 14 13 15 0 2
5 9 11 11 11 2
44 6 2 15 13 3 11 9 2 7 15 13 1 10 0 9 15 15 13 2 16 10 9 2 0 2 1 14 13 1 9 1 0 9 2 13 16 15 13 0 3 9 1 15 2
38 15 13 0 0 1 7 4 3 13 9 1 11 1 9 1 16 10 9 3 13 3 1 9 2 3 3 13 3 2 7 9 13 14 13 15 0 0 2
31 7 15 13 0 9 15 0 13 1 15 2 7 15 13 16 15 13 0 14 13 9 1 2 3 16 10 9 4 13 0 2
37 15 13 15 16 9 7 9 4 13 15 9 1 14 13 16 13 15 13 2 7 0 1 14 4 13 9 1 9 1 9 2 15 11 11 11 13 2
6 15 13 3 11 9 2
2 9 2
6 11 11 2 1 9 2
6 11 11 2 11 2 2
40 15 4 0 13 9 14 13 16 15 1 10 9 13 15 3 1 9 15 13 0 1 11 9 1 9 1 9 2 7 15 4 3 13 14 13 0 9 1 15 2
8 3 13 15 1 10 0 9 2
18 15 13 0 16 16 15 13 9 2 13 11 9 1 11 3 0 1 2
21 3 2 1 16 15 4 13 9 2 13 15 1 9 0 1 10 9 15 11 13 2
32 16 15 13 1 9 1 2 13 15 10 0 9 1 14 13 16 15 1 12 4 13 3 0 9 1 15 15 4 13 1 9 2
26 3 13 9 3 15 3 1 9 4 13 1 9 15 13 16 15 4 13 10 9 15 4 13 1 11 2
7 7 3 13 9 1 11 2
25 10 0 9 10 1 14 13 0 9 13 15 11 4 13 1 1 16 15 0 4 13 14 13 9 2
30 16 15 13 9 2 3 4 15 13 1 0 9 1 10 0 0 9 2 7 15 13 3 0 1 10 9 15 13 1 2
5 7 10 9 13 2
15 10 9 13 15 9 4 13 14 13 1 14 13 11 9 2
5 9 11 11 11 2
11 15 13 0 0 1 11 0 9 1 9 2
28 15 4 13 16 10 9 3 2 15 0 13 0 1 10 9 2 4 13 0 3 2 1 14 13 9 1 9 2
31 15 13 0 0 15 11 11 13 2 16 15 13 3 0 1 11 14 13 9 1 11 16 15 13 0 9 0 1 0 9 2
30 3 1 10 9 4 15 13 9 1 2 15 13 15 13 2 1 12 9 1 9 1 9 9 1 14 13 9 1 11 2
33 4 15 1 9 13 10 12 0 9 1 11 2 4 10 9 2 1 15 15 13 2 13 1 12 2 7 15 4 13 15 3 0 2
10 3 13 15 3 3 15 13 0 9 2
65 16 15 13 14 13 9 2 4 3 11 3 13 1 1 11 10 9 9 1 9 15 13 15 2 3 0 15 13 2 3 3 2 7 15 13 0 1 2 9 13 2 0 9 2 13 2 9 2 3 15 4 13 7 9 7 10 9 1 9 1 14 13 15 1 2
2 9 2
7 7 3 4 9 13 9 2
5 9 11 11 11 2
7 15 13 15 10 9 1 2
2 9 2
6 11 11 2 1 9 2
6 11 11 2 11 2 2
49 15 13 1 3 0 0 16 9 13 1 15 15 13 1 1 10 9 2 7 15 13 3 0 15 13 1 16 15 3 0 3 1 3 4 13 15 1 16 9 1 11 4 13 1 14 13 10 10 2
7 10 9 13 1 12 9 2
13 16 9 13 1 0 9 2 10 9 13 15 3 2
25 9 1 10 9 13 3 3 16 15 13 0 1 1 9 9 1 14 13 15 10 0 9 1 11 2
9 10 0 9 15 4 13 2 13 2
56 3 13 15 3 0 1 10 9 15 1 11 11 13 2 3 16 15 1 9 13 0 1 9 1 0 9 1 9 2 9 2 15 4 13 1 10 9 16 15 13 0 9 1 9 2 1 3 14 13 9 3 0 1 10 9 2
17 13 15 0 3 16 9 13 14 13 1 10 0 9 1 10 9 2
5 9 11 11 11 2
47 16 15 13 9 2 13 15 3 0 1 15 14 13 10 0 9 1 15 2 16 15 3 13 0 9 1 15 1 10 9 15 13 1 9 2 7 15 4 3 1 10 0 9 13 10 9 2
45 7 15 13 1 16 11 13 1 10 9 2 11 11 13 15 2 1 15 15 3 13 2 1 9 1 10 0 0 9 2 7 15 13 15 15 11 11 11 13 1 1 11 1 9 2
26 15 13 15 13 0 9 2 7 15 13 16 15 4 4 13 16 15 13 15 13 1 10 0 0 9 2
44 6 2 15 13 3 0 1 10 9 15 11 11 7 10 4 13 1 16 15 13 9 1 9 2 15 15 1 0 9 13 0 1 2 15 0 3 4 4 13 1 0 0 9 2
22 7 15 13 3 16 15 13 9 1 9 1 10 9 1 16 15 10 13 9 1 15 2
42 15 4 1 9 3 13 1 9 9 0 15 13 16 15 13 9 1 16 10 0 9 1 15 13 10 9 1 10 9 2 7 10 9 13 15 1 0 3 1 9 3 2
2 9 2
13 3 13 15 0 1 10 9 2 1 11 11 11 2
7 11 11 11 2 11 2 2
17 15 13 3 10 9 1 9 2 0 1 10 9 1 11 1 9 2
6 1 0 9 13 15 2
8 2 9 13 11 1 11 2 2
13 7 1 1 9 13 15 1 9 11 11 1 11 2
24 2 0 1 12 13 11 9 1 16 15 13 14 13 1 9 0 15 10 0 9 13 1 2 2
12 9 13 10 9 1 9 9 15 13 1 11 2
35 1 12 13 15 12 12 2 7 3 1 16 11 13 1 2 13 15 1 12 12 12 2 7 1 12 13 15 3 1 1 9 1 12 12 2
9 9 13 3 0 1 1 10 9 2
22 4 11 13 0 7 13 9 1 16 15 3 13 1 12 12 9 10 9 1 9 1 2
40 10 9 4 15 13 1 0 9 1 10 0 9 16 15 3 13 9 1 9 1 10 9 15 3 4 13 1 11 2 7 10 0 9 15 13 1 10 0 9 2
15 4 11 0 13 12 12 1 9 1 9 1 9 7 10 2
5 9 11 11 11 2
4 15 13 0 2
41 9 13 15 0 0 1 16 15 4 13 1 9 7 9 1 10 9 9 2 7 10 9 13 1 9 3 0 9 3 1 11 2 1 10 0 9 0 1 11 9 2
14 15 13 16 10 9 13 14 13 9 7 9 1 9 2
19 0 4 10 9 4 13 10 9 1 0 9 1 14 13 1 11 1 9 2
17 15 13 15 0 1 2 7 15 13 15 1 10 9 1 14 13 2
19 7 15 16 15 13 0 9 1 11 2 13 3 16 10 15 3 13 9 2
35 15 13 1 9 1 10 0 9 2 7 3 13 15 3 16 14 13 1 10 9 3 1 0 13 0 1 9 2 16 15 13 10 9 0 2
33 0 1 1 10 9 3 15 4 13 0 0 9 1 0 9 3 2 3 13 15 0 7 13 0 3 16 15 13 9 1 10 9 2
17 16 10 9 13 10 0 0 9 7 9 2 4 3 15 13 1 2
17 15 13 16 15 4 13 10 9 15 13 0 7 3 0 0 0 2
7 11 11 11 2 11 2 2
8 11 11 1 10 0 11 13 2
25 2 15 13 10 9 1 16 11 13 10 0 9 0 2 7 16 15 3 13 0 15 13 1 11 2
24 15 13 3 0 9 14 13 9 1 11 2 7 3 13 9 1 16 15 4 13 1 9 2 2
16 10 3 0 13 3 9 3 2 16 15 4 13 1 10 9 2
29 9 1 9 13 3 3 16 15 3 4 13 1 10 9 2 7 16 9 13 0 0 1 15 15 4 13 11 9 2
23 3 13 15 1 1 16 11 3 4 13 10 9 1 14 13 9 9 1 10 0 0 9 2
38 7 16 9 13 1 16 3 10 4 13 0 9 2 3 13 3 15 1 9 2 3 0 15 13 2 1 10 9 15 3 3 13 1 12 12 1 9 2
32 3 0 4 10 0 9 1 9 1 9 1 10 10 10 15 13 2 13 16 11 13 1 10 0 0 15 13 9 7 3 9 2
5 9 11 11 11 2
23 13 15 3 13 16 15 15 4 13 0 9 2 0 3 13 9 1 11 1 10 10 9 2
36 15 13 10 9 1 9 1 15 2 7 15 13 15 15 13 10 9 2 15 13 9 2 3 0 9 2 3 16 3 10 9 4 13 0 3 2
38 15 13 0 14 13 1 0 9 3 2 16 15 13 9 7 9 1 1 9 15 13 3 0 15 4 13 9 1 11 2 7 3 3 0 15 4 13 2
9 15 13 3 3 0 15 13 9 2
10 3 13 15 0 14 13 1 0 9 2
22 15 13 16 10 9 7 9 15 3 13 2 13 0 2 7 15 13 0 9 1 11 2
47 15 13 0 1 9 11 1 12 9 2 7 15 13 16 9 3 13 0 0 1 0 9 2 7 15 13 3 0 1 14 13 1 10 9 7 13 10 9 15 13 1 1 14 13 1 9 2
8 15 13 15 0 3 1 3 2
6 11 11 2 11 2 2
18 11 13 0 1 16 15 4 13 10 0 9 1 9 1 9 7 9 2
19 7 1 10 9 13 15 0 1 10 9 15 4 13 1 11 9 7 9 2
71 7 16 15 13 9 1 15 2 4 15 3 13 9 1 9 1 9 1 7 9 1 9 2 7 9 1 9 1 10 0 9 1 9 2 16 15 13 0 7 0 0 9 2 7 3 15 4 13 16 9 4 13 12 9 1 9 16 15 4 13 10 9 7 4 4 13 9 1 10 9 2
38 1 9 4 15 0 3 13 10 9 7 9 15 13 0 0 1 10 0 9 7 10 9 2 7 15 13 16 11 13 16 1 9 13 3 9 3 0 2
5 15 4 13 9 2
16 13 15 0 3 14 13 10 0 9 1 11 1 10 10 9 2
5 7 9 9 12 2
14 15 13 16 10 9 13 0 1 1 9 1 0 9 2
11 15 4 11 13 1 1 14 13 10 9 2
5 9 11 11 11 2
45 1 10 0 4 15 13 16 15 13 0 1 16 11 13 16 15 1 9 13 0 1 10 9 15 13 1 10 9 7 9 2 7 15 13 16 15 13 10 0 9 1 15 1 11 2
35 3 13 15 0 1 9 11 1 2 15 15 3 3 4 13 10 9 9 2 16 15 13 0 1 10 3 0 9 15 15 13 1 0 9 2
14 15 13 3 16 9 3 13 3 0 15 15 4 13 2
33 15 13 0 9 1 0 9 1 9 1 1 10 9 15 13 1 9 7 9 2 15 4 3 0 13 3 1 10 9 7 10 9 2
22 7 15 13 15 3 1 2 15 13 0 1 3 10 12 9 2 7 13 14 13 9 2
18 16 15 13 0 9 2 13 15 0 1 9 11 1 16 15 13 0 2
19 15 4 11 0 13 2 7 1 11 7 1 9 15 3 13 1 1 11 2
33 9 13 15 1 9 2 15 4 13 7 1 9 1 10 9 2 9 1 9 2 7 10 9 15 4 13 1 0 9 1 3 9 2
2 9 2
7 15 13 0 1 10 9 2
6 11 11 2 11 2 2
35 16 15 13 9 0 9 2 4 15 13 16 15 13 9 13 10 0 9 3 1 9 2 3 16 3 15 4 13 9 1 10 10 0 9 2
31 15 4 13 9 9 1 9 1 10 9 15 13 1 11 9 2 3 15 13 9 1 9 7 1 0 9 7 1 0 9 2
20 3 13 15 3 0 1 16 15 3 13 14 13 15 16 15 13 9 7 9 2
7 7 15 4 3 13 9 2
6 10 9 4 11 13 2
5 9 11 11 11 2
30 13 15 1 10 0 13 16 15 13 11 9 2 16 15 13 9 7 9 1 16 15 13 14 13 9 1 15 1 9 2
9 15 13 15 3 15 14 13 1 2
39 16 15 13 9 15 13 1 9 1 10 9 7 3 1 9 2 13 11 0 1 16 15 4 13 9 2 7 16 15 4 13 0 9 1 9 1 10 9 2
13 7 1 10 9 1 9 13 15 0 1 12 9 2
11 10 12 13 9 2 7 10 10 13 9 2
31 1 7 1 12 4 9 13 2 3 16 9 1 0 9 1 12 12 9 3 4 13 1 9 2 13 0 9 15 4 13 2
39 9 4 3 1 9 1 9 1 0 9 13 1 0 9 1 9 1 16 9 1 0 9 4 4 13 10 9 1 14 13 1 15 7 13 1 0 0 9 2
22 10 0 9 4 13 14 13 9 2 3 16 9 1 9 3 13 0 1 9 1 9 2
12 3 4 9 1 9 13 15 15 13 1 12 2
18 15 13 0 9 3 1 9 9 1 16 0 9 13 1 9 0 0 2
21 3 4 15 3 13 1 9 1 10 0 0 9 1 9 2 7 10 9 1 9 2
58 10 9 15 10 9 13 2 3 0 15 13 2 13 3 16 15 3 13 9 1 0 0 9 2 3 15 15 13 1 9 7 13 3 1 9 7 9 2 16 15 13 15 1 10 9 2 3 2 4 15 13 2 9 0 1 0 9 2
32 15 13 1 10 9 11 3 4 13 7 13 1 11 2 7 3 1 9 1 9 15 13 0 1 10 10 2 1 9 1 9 2
6 11 11 2 11 2 2
16 3 0 15 13 2 13 9 9 16 15 4 13 1 10 9 2
31 7 10 9 13 15 9 1 16 15 13 3 15 15 13 2 15 13 7 13 2 7 15 13 3 3 10 0 1 1 15 2
6 7 10 9 13 3 2
16 4 15 1 10 12 9 13 0 2 0 2 0 9 1 9 2
5 9 11 11 11 2
38 3 0 15 13 10 10 9 2 13 15 3 3 13 1 2 7 15 13 3 13 1 9 1 10 9 15 13 0 1 9 2 7 3 1 9 7 9 2
6 15 13 10 0 9 2
11 3 13 3 10 9 1 11 11 9 3 2
37 6 2 15 4 13 9 1 0 9 1 10 9 15 15 3 4 13 1 1 2 3 3 1 10 2 7 15 13 10 12 15 3 0 13 1 9 2
28 15 13 3 16 15 3 13 1 9 1 11 15 15 13 13 0 1 10 10 9 2 1 9 1 9 1 9 2
2 9 2
7 15 13 9 2 11 11 2
6 11 11 2 11 2 2
15 1 0 7 1 0 9 13 3 9 1 0 9 0 0 2
21 3 1 4 10 0 9 13 16 9 1 11 13 3 3 1 2 3 3 1 9 2
26 7 15 13 16 16 0 9 13 16 9 0 13 1 9 1 9 2 3 13 15 10 9 1 0 9 2
7 7 10 9 1 9 13 2
41 16 15 13 14 13 9 2 16 15 13 14 13 9 2 7 16 15 13 14 13 10 9 1 9 2 4 15 13 3 1 16 9 1 9 1 9 7 9 4 13 2
32 1 11 13 15 10 0 9 16 15 4 13 2 3 16 15 4 13 10 0 0 9 1 9 1 9 1 9 7 9 7 9 2
6 7 10 9 13 3 2
23 16 15 13 15 2 4 15 13 3 1 9 1 15 15 13 11 9 2 7 3 13 15 2
8 15 4 13 10 9 1 9 2
5 9 11 11 11 2
32 13 15 3 13 16 11 13 9 1 16 0 13 4 15 3 13 16 0 9 13 0 0 1 9 1 10 9 2 3 10 0 2
33 7 15 13 10 9 0 9 1 9 15 15 13 3 3 14 13 1 2 7 13 1 14 13 2 7 15 4 13 1 10 9 10 2
22 16 15 13 9 1 9 1 9 7 9 2 4 3 11 13 9 1 14 13 10 9 2
9 15 4 1 4 13 1 10 9 2
17 16 15 13 9 2 13 15 0 9 2 15 15 3 4 13 1 2
6 11 11 2 11 2 2
16 3 4 15 13 9 16 15 4 13 1 14 13 10 9 9 2
23 11 4 9 1 9 13 1 16 11 4 13 1 10 9 1 9 2 9 2 9 7 9 2
8 15 4 10 0 9 13 1 2
37 7 3 13 9 1 10 9 1 11 11 10 9 16 15 15 11 13 1 3 2 7 15 4 13 1 9 2 13 12 9 2 9 7 9 5 9 2
7 15 13 11 1 1 9 2
5 9 11 11 11 2
13 6 2 15 13 1 10 12 9 2 9 7 9 2
30 7 15 4 3 13 16 15 1 15 13 1 0 9 2 15 15 3 9 11 13 1 16 11 4 13 11 13 1 1 2
27 1 9 1 9 7 9 2 15 15 4 13 1 1 1 9 1 11 11 2 13 15 3 1 9 7 9 2
23 16 15 13 14 13 1 15 11 3 4 13 1 2 7 15 15 10 1 0 9 4 13 2
2 9 2
8 3 13 15 0 1 10 9 2
2 9 2
8 15 13 9 2 11 11 11 2
7 11 11 11 2 11 2 2
17 15 13 15 9 9 1 16 15 13 9 1 11 15 13 10 0 2
72 1 10 9 4 15 3 13 9 16 15 3 13 0 1 16 15 3 1 15 10 13 9 13 1 9 1 9 15 4 13 10 0 1 10 9 9 1 10 9 2 7 16 15 13 9 15 4 13 1 9 2 15 13 10 0 2 7 15 1 10 0 9 7 9 13 10 9 1 14 13 1 2
35 16 15 3 4 13 1 11 1 9 16 10 9 13 9 4 13 2 13 15 15 15 13 16 15 13 10 9 1 14 13 1 1 10 9 2
16 7 15 13 3 9 1 10 9 13 1 9 2 7 9 9 2
5 9 11 11 11 2
14 15 4 1 9 13 15 0 1 9 11 9 1 15 2
40 15 13 0 16 4 10 15 2 3 15 15 13 1 0 9 2 13 1 9 1 10 9 2 3 13 15 10 3 3 3 0 2 7 0 9 7 9 1 15 2
38 16 10 9 9 13 1 9 1 9 2 4 15 15 13 1 9 1 15 2 4 13 1 9 1 9 7 9 1 0 9 2 0 1 9 1 10 9 2
36 15 4 15 3 13 0 14 13 10 0 9 1 1 9 2 15 4 13 3 7 3 3 10 9 13 2 3 0 15 13 15 1 15 2 3 2
2 9 2
6 11 11 2 1 9 2
6 11 11 2 11 2 2
49 15 13 15 10 13 9 1 14 13 9 1 15 15 4 13 3 2 7 15 15 4 13 0 2 7 15 4 3 13 14 13 1 10 0 0 9 1 9 1 15 15 4 13 1 9 11 1 9 2
39 10 9 13 16 15 3 13 0 14 13 1 15 15 4 13 1 9 1 9 2 16 11 4 13 9 1 15 1 10 9 1 9 7 1 10 9 1 9 2
31 9 13 16 3 11 3 13 0 1 14 13 1 1 11 9 15 13 1 0 9 1 15 15 13 1 0 9 1 11 9 2
27 11 13 1 0 0 7 0 1 11 9 1 10 9 0 1 9 2 7 3 1 15 11 4 13 1 9 2
36 13 3 3 15 9 1 14 13 9 15 13 1 0 9 2 7 15 4 13 10 9 1 10 9 15 13 1 10 3 0 7 0 7 0 9 2
5 9 11 11 11 2
28 15 13 1 3 0 0 1 10 0 9 16 15 4 13 1 9 16 15 13 1 0 9 1 11 9 1 9 2
11 15 4 3 3 13 15 3 1 10 9 2
20 15 4 3 13 10 9 9 1 9 7 1 0 2 0 7 10 9 1 9 2
33 15 4 9 0 13 1 7 13 14 13 9 1 2 7 1 10 9 2 3 15 13 9 2 13 15 3 10 9 1 15 1 9 2
13 3 13 3 11 10 0 9 1 14 13 10 9 2
22 15 13 1 0 3 1 9 15 3 4 13 10 9 2 7 15 15 4 13 9 1 2
22 7 15 4 3 2 15 15 4 13 0 2 13 10 9 3 0 10 9 15 4 13 2
49 16 15 4 13 10 0 9 1 11 9 2 13 15 3 0 0 9 1 2 15 4 15 13 4 13 10 10 1 2 7 15 13 3 16 11 4 13 0 1 15 1 10 9 16 15 4 13 1 2
2 9 2
8 15 13 3 0 1 10 9 2
6 11 11 2 11 2 2
7 15 13 10 9 1 9 2
26 15 13 16 11 2 11 11 2 1 9 13 1 9 1 14 13 0 9 1 14 13 9 1 1 9 2
15 1 9 13 10 0 9 16 11 13 0 9 1 10 9 2
18 15 13 16 10 9 1 9 4 13 10 9 1 1 9 3 1 9 2
45 1 9 13 15 10 9 16 10 9 1 9 2 0 7 9 2 4 13 1 9 2 7 16 15 13 9 2 13 15 3 11 15 4 13 1 0 9 2 7 15 13 10 0 9 2
21 13 9 15 13 0 7 0 16 11 4 13 9 9 1 14 4 13 10 9 0 2
4 9 11 11 2
45 16 15 13 9 1 9 1 9 2 0 7 9 1 10 2 13 15 3 15 13 10 9 14 13 1 7 13 9 1 15 2 15 4 15 13 1 10 9 15 13 0 1 10 9 2
28 16 15 13 9 2 4 15 13 10 0 9 1 11 1 16 9 1 10 13 10 9 9 10 4 13 1 15 2
24 15 13 10 10 9 1 15 15 3 13 1 11 2 16 15 13 0 9 15 13 9 1 9 2
28 1 11 13 15 3 16 15 13 9 10 15 1 9 4 13 1 14 13 10 9 15 13 0 1 14 13 9 2
32 3 4 3 3 15 15 4 13 10 9 2 9 2 4 13 0 9 1 14 13 10 9 15 4 13 1 10 9 11 4 13 2
48 1 9 15 11 4 13 2 15 3 13 1 11 1 9 2 13 15 16 15 13 10 9 15 15 3 4 13 1 9 2 7 16 9 7 9 1 9 7 9 13 10 9 15 9 10 4 13 2
33 15 13 3 0 16 15 13 1 10 9 15 10 0 4 13 2 7 15 13 15 10 9 1 1 10 9 16 15 13 1 10 9 2
6 11 11 2 11 2 2
46 15 13 0 15 9 13 2 16 9 13 10 0 7 1 10 9 0 9 1 11 2 7 1 9 1 12 9 2 1 10 9 9 3 2 13 12 0 9 0 2 7 15 4 13 9 2
11 15 13 11 11 2 11 11 7 11 11 2
26 7 15 15 13 1 9 1 10 0 9 1 9 2 13 16 15 0 13 10 0 9 1 9 1 11 2
27 4 15 4 13 10 9 7 13 0 0 9 2 4 3 15 1 9 1 7 1 4 13 9 0 1 11 2
36 15 13 0 9 1 9 1 9 16 9 13 0 1 9 2 7 15 4 13 0 14 13 9 7 1 11 7 11 7 1 0 9 1 10 9 2
15 4 9 13 10 9 2 3 16 9 4 13 1 1 9 2
4 9 11 11 2
31 1 10 9 1 10 9 13 15 3 1 9 1 14 4 13 16 15 13 9 15 4 13 9 1 16 0 9 4 13 0 2
22 15 13 0 9 15 13 1 16 10 9 13 0 7 3 2 15 13 1 9 1 10 2
32 15 4 3 13 16 1 11 9 4 15 13 9 1 11 1 9 2 7 3 4 3 11 4 13 3 10 9 15 11 3 13 2
32 7 10 9 2 7 15 15 15 3 13 1 11 2 13 16 15 13 14 13 10 9 15 1 9 13 2 1 10 9 15 13 2
45 15 4 13 1 16 15 4 13 0 1 9 1 11 9 7 10 9 15 13 2 15 15 13 15 4 13 1 11 9 2 7 15 15 13 10 10 0 9 16 15 4 13 1 9 2
12 1 15 4 3 11 1 10 9 13 10 9 2
6 11 11 2 11 2 2
7 15 13 10 9 1 9 2
26 9 13 0 9 1 9 16 9 11 11 7 10 3 3 4 13 0 9 1 9 7 9 11 11 11 2
20 1 15 13 11 16 11 3 13 9 1 9 16 15 13 9 11 1 0 9 2
28 9 13 9 15 4 13 0 9 1 9 7 10 9 2 7 1 0 9 13 9 3 3 0 9 1 9 10 2
25 11 9 13 3 3 0 1 9 1 15 11 13 16 15 13 10 0 9 1 9 1 12 2 12 2
20 9 1 15 13 3 14 13 9 1 9 7 3 13 1 9 1 9 1 9 2
14 11 9 1 11 13 0 16 9 13 0 9 1 0 2
25 7 10 9 1 9 11 13 16 15 13 16 9 13 1 9 1 9 9 7 11 9 1 0 9 2
4 9 11 11 2
26 11 9 1 0 9 1 10 9 13 10 9 1 10 9 1 11 11 1 10 9 15 4 13 1 11 2
9 15 13 9 1 11 9 1 15 2
20 11 9 4 13 1 10 0 9 1 11 11 9 7 9 1 9 1 11 9 2
42 1 16 9 4 13 0 2 4 11 13 9 1 11 11 11 2 15 13 16 15 4 13 3 0 2 7 11 4 13 9 1 11 11 2 15 13 15 4 13 3 0 2
62 11 9 13 1 10 9 1 10 9 15 10 0 4 13 11 11 11 1 9 2 7 10 9 15 13 1 14 13 10 9 1 9 1 9 2 7 1 1 15 4 15 13 1 1 10 9 15 13 14 13 9 1 0 0 9 1 9 1 10 12 9 2
6 11 11 2 11 2 2
14 15 4 3 13 15 0 0 1 9 7 0 1 9 2
53 3 13 15 0 13 1 11 2 15 13 0 16 9 15 11 4 13 2 13 1 9 1 9 7 3 3 1 9 1 7 9 7 9 2 16 15 1 10 9 1 14 13 0 9 1 9 0 13 0 9 1 9 2
25 15 13 3 10 9 16 15 13 9 2 7 3 4 15 3 4 13 1 0 9 1 10 0 9 2
50 7 10 9 13 3 16 3 9 4 13 15 1 10 9 16 15 13 10 9 1 11 2 15 1 10 9 4 13 1 11 1 14 13 15 1 14 13 1 0 9 1 9 1 11 11 7 10 0 9 2
4 9 11 11 2
36 1 9 1 11 9 1 0 9 13 15 3 10 0 9 1 10 9 15 11 4 13 9 1 2 7 1 10 9 15 11 11 4 13 9 1 2
10 15 4 3 13 9 1 9 1 9 2
25 1 10 9 2 15 3 13 0 2 7 1 10 9 0 0 2 13 3 11 1 10 9 1 9 2
11 15 13 3 1 9 16 11 13 10 9 2
14 15 4 13 16 11 3 13 10 0 0 9 1 11 2
17 15 4 13 10 9 1 9 1 9 1 10 9 15 11 4 13 2
2 9 2
9 10 9 4 4 13 1 11 11 2
27 9 13 0 1 16 15 13 0 1 9 2 7 1 11 9 4 11 13 16 9 11 3 4 13 10 9 2
6 2 10 9 4 13 2
6 11 11 2 11 2 2
7 15 13 10 9 1 9 2
14 11 4 13 16 15 4 13 10 0 9 1 10 9 2
15 15 4 13 10 0 9 0 9 2 1 13 15 0 9 2
18 11 13 16 10 0 9 3 4 13 15 1 10 0 9 7 10 0 2
28 15 13 3 9 1 10 9 2 7 10 9 4 13 15 1 10 0 7 0 9 2 7 15 13 3 9 9 2
42 16 10 0 9 1 9 13 15 14 13 14 13 15 1 10 0 9 2 4 15 13 2 13 2 13 2 13 2 0 1 9 2 16 15 13 1 9 2 13 7 13 2
9 15 4 13 1 9 3 1 11 2
10 13 9 15 1 10 0 9 1 11 2
21 7 10 9 4 9 7 11 13 14 13 1 14 13 10 9 1 9 1 10 9 2
5 9 11 11 11 2
25 13 15 0 13 16 15 13 0 16 1 11 13 0 9 2 15 3 13 1 9 15 15 4 13 2
15 3 13 15 0 3 10 9 1 15 9 11 3 13 1 2
29 9 15 13 1 10 10 9 2 13 9 1 9 9 2 7 9 4 13 1 1 1 9 1 15 15 4 13 15 2
6 15 4 13 11 9 2
31 15 4 3 13 9 1 10 9 7 9 2 7 15 15 0 13 10 9 15 11 13 2 13 0 0 9 1 9 1 15 2
31 7 15 15 3 4 13 15 2 7 15 4 13 1 10 9 15 11 13 1 2 13 0 10 0 9 10 9 1 14 13 2
6 11 11 2 11 2 2
5 15 13 10 9 2
17 15 4 0 13 1 10 9 2 7 15 13 15 1 9 14 13 2
8 15 13 9 1 0 0 9 2
4 10 9 13 2
38 15 13 1 9 9 1 0 9 2 1 4 15 13 16 15 4 13 9 1 0 9 16 9 3 4 13 11 7 13 10 9 15 15 3 4 13 1 2
7 13 15 0 9 1 9 2
12 7 4 15 13 10 9 15 13 1 1 9 2
5 9 11 11 11 2
18 1 10 9 13 10 9 3 3 10 9 1 9 1 9 2 1 9 2
32 16 9 13 16 9 4 13 9 1 10 0 9 2 7 15 13 1 1 0 9 7 9 2 4 15 13 9 1 9 1 15 2
12 15 13 0 1 9 2 9 7 9 14 13 2
24 7 10 0 9 2 7 15 13 0 7 10 2 4 0 3 13 10 9 1 9 1 0 9 2
4 16 15 13 2
17 9 15 0 13 11 9 1 0 9 2 13 9 1 9 1 15 2
28 7 16 15 3 13 15 2 7 3 4 13 1 0 9 2 13 15 3 9 9 14 13 1 7 13 10 9 2
7 7 15 4 0 4 13 2
2 9 2
16 10 0 9 13 3 3 2 7 15 13 1 1 10 0 9 2
4 9 1 11 5
4 9 11 11 2
21 1 16 9 11 13 14 13 1 2 4 11 1 10 0 9 1 11 13 15 9 2
16 9 1 9 13 10 0 9 1 9 1 10 0 9 7 9 2
11 15 13 0 9 1 9 1 9 7 9 2
16 9 13 10 9 1 11 9 7 13 1 9 1 9 1 11 2
24 15 4 13 10 9 1 9 1 14 13 9 1 9 15 4 13 1 0 7 0 9 1 9 2
5 11 13 9 9 2
9 15 13 10 9 1 9 7 9 2
5 15 13 0 9 2
20 15 13 10 0 9 2 10 0 9 2 7 15 13 1 10 0 9 1 9 2
11 15 13 15 2 7 15 13 15 1 9 2
43 1 9 1 14 13 2 2 10 0 9 2 10 9 15 13 0 1 10 0 9 2 10 9 16 3 0 9 13 0 2 0 9 2 0 9 2 0 9 7 0 0 9 5
8 15 13 9 1 10 0 9 2
6 15 13 9 1 11 2
7 9 9 4 3 13 15 2
16 15 4 13 1 10 9 1 0 9 2 0 9 7 0 9 2
28 9 1 15 15 13 10 0 9 2 13 16 15 13 9 1 9 1 15 7 9 1 10 10 9 7 1 9 2
12 10 9 13 15 1 15 1 1 10 0 9 2
22 1 10 10 9 13 10 0 0 9 14 13 9 1 9 15 3 13 10 9 1 9 2
6 11 4 13 1 15 2
13 10 0 9 1 10 9 13 9 2 9 7 9 2
9 10 0 9 13 3 14 13 9 2
10 1 9 2 9 2 9 7 0 9 2
4 15 13 9 2
4 15 13 9 2
4 15 4 13 2
40 10 7 10 1 15 4 13 9 2 7 9 2 1 14 13 9 1 15 7 10 2 7 4 13 16 10 9 15 3 13 1 9 1 15 2 4 9 13 1 2
13 15 4 13 9 1 14 13 15 2 13 7 13 2
9 15 4 13 0 9 15 13 9 2
6 0 9 13 0 9 2
6 0 9 13 0 9 2
4 15 13 11 2
9 15 4 13 1 14 13 7 13 2
11 4 15 13 2 4 9 13 10 0 9 2
9 0 9 13 3 0 1 0 9 2
13 0 9 13 14 13 9 1 15 7 10 0 9 2
12 0 9 13 14 13 1 9 9 1 0 9 2
7 9 13 10 0 1 15 2
17 0 9 13 14 13 16 10 9 4 13 15 0 3 0 1 9 2
26 0 9 13 14 13 10 0 9 1 9 1 9 2 3 16 15 4 13 7 0 9 7 0 9 0 2
11 9 9 2 9 7 9 13 11 0 9 2
7 15 4 13 9 1 9 2
7 15 4 13 15 14 13 2
7 15 4 13 0 14 13 2
15 10 9 13 14 13 15 15 1 9 13 0 2 1 9 2
13 0 4 11 13 10 0 9 2 0 9 1 9 2
13 3 1 9 13 15 3 0 9 1 9 7 9 2
9 15 13 0 9 1 9 1 9 2
11 15 4 13 3 0 9 1 10 0 9 2
16 3 4 15 13 0 9 1 10 9 1 9 2 3 1 9 2
14 3 4 15 13 10 9 15 13 15 15 15 4 13 2
21 3 4 15 13 10 9 16 0 13 7 13 2 7 16 15 13 9 1 10 0 2
17 3 4 15 13 9 7 9 15 13 15 0 14 13 9 7 9 2
9 1 10 0 9 13 15 0 9 2
14 9 9 13 0 0 1 15 15 13 9 1 0 9 2
13 15 4 4 13 16 9 9 13 0 1 10 9 2
15 15 13 1 10 0 9 1 0 9 3 1 10 0 9 2
9 15 4 13 0 9 1 14 13 2
5 9 9 4 13 2
14 7 9 1 0 9 4 3 3 13 1 0 0 9 2
13 15 4 13 9 1 0 9 7 0 9 1 9 2
49 15 4 13 0 7 13 16 15 4 13 9 10 1 10 0 9 2 0 1 14 13 1 9 1 9 15 13 0 9 2 9 1 9 2 9 1 9 7 9 2 9 1 9 7 9 1 0 9 2
15 9 4 13 10 0 9 7 13 15 0 1 9 7 9 2
10 9 9 4 13 16 15 0 13 15 2
9 7 9 4 1 9 13 1 9 2
9 9 7 9 4 13 10 0 9 2
10 3 13 9 3 0 7 9 3 0 2
9 3 4 15 13 10 9 7 9 2
26 9 4 13 14 13 10 9 1 0 15 13 14 13 0 9 2 7 15 3 4 13 10 10 9 0 2
11 11 4 13 1 9 1 9 1 0 9 2
16 9 13 1 0 9 1 9 7 9 1 7 0 7 0 9 2
12 15 13 16 0 9 4 13 10 9 1 9 2
18 9 7 9 1 10 9 1 9 4 13 9 1 9 7 10 0 9 2
9 3 13 0 2 0 9 1 9 2
7 0 7 0 9 4 13 2
9 9 7 9 13 0 0 1 15 2
7 9 4 13 10 0 9 2
17 15 4 13 9 1 9 7 13 9 9 1 14 13 15 10 9 2
65 15 4 13 10 0 9 9 1 0 9 0 2 2 10 0 9 15 13 0 9 1 0 9 2 7 15 13 10 0 9 2 10 0 9 15 13 9 9 2 7 16 15 13 9 1 9 7 9 2 10 0 7 0 9 2 0 9 1 9 2 9 7 9 10 5
9 15 4 13 0 1 9 1 9 2
11 11 4 3 13 15 1 10 0 0 9 2
9 9 4 13 11 9 1 10 9 2
8 9 4 13 1 9 1 9 2
16 15 15 13 1 9 2 13 15 15 13 1 1 9 7 9 2
7 3 13 9 10 0 9 2
14 9 13 0 9 2 0 9 2 0 9 7 0 9 2
16 9 4 13 1 0 9 2 9 7 1 16 0 13 14 13 2
18 9 4 13 9 1 14 13 9 3 16 9 7 9 1 9 13 0 2
8 15 13 15 0 0 9 1 2
8 11 4 13 10 9 1 9 2
26 9 4 13 1 10 0 9 1 9 1 9 7 9 7 4 1 9 1 15 13 1 0 9 7 9 2
20 1 9 1 0 9 4 9 11 3 13 0 9 1 10 9 2 7 9 13 2
10 10 9 13 1 0 9 1 10 9 2
10 1 10 0 9 13 0 9 1 9 2
7 1 9 9 13 15 0 2
26 9 4 13 9 1 14 13 1 16 11 1 9 4 13 10 1 10 9 1 14 13 9 1 0 9 2
14 9 1 9 1 11 4 13 1 9 1 10 0 9 2
18 11 4 13 0 0 9 7 0 9 13 1 14 13 3 0 0 9 2
21 9 4 13 9 1 10 0 9 1 9 7 9 1 14 13 9 9 1 9 11 2
19 9 13 10 9 1 10 0 9 9 16 9 13 3 1 14 13 1 9 2
11 11 4 13 9 1 10 9 1 10 9 2
26 15 13 1 1 9 1 11 9 2 15 4 13 1 14 13 9 7 13 10 0 9 1 9 1 9 2
25 9 7 0 9 4 13 9 0 1 2 7 4 13 1 9 1 9 7 9 1 0 1 0 9 2
9 1 14 13 9 4 0 9 13 2
5 3 4 15 13 2
13 0 9 4 13 15 2 7 15 4 3 13 15 2
25 9 4 13 7 13 0 9 1 0 9 1 9 2 0 0 7 1 9 1 10 0 7 10 9 2
19 15 13 1 0 9 1 10 9 15 13 15 0 9 7 0 9 1 9 2
18 10 0 13 9 1 9 2 0 7 0 9 13 3 10 9 14 13 2
25 13 15 0 1 0 9 15 3 13 2 3 13 15 9 1 9 2 3 13 15 9 7 13 9 2
6 15 13 15 10 1 2
13 9 13 9 2 7 9 13 15 0 1 0 9 2
21 15 0 9 13 2 4 15 13 3 0 16 9 7 13 7 13 1 10 0 9 2
3 0 9 2
18 10 9 1 15 2 7 10 9 1 9 15 13 3 16 15 13 15 2
4 9 13 9 2
18 9 13 3 1 9 1 14 13 9 1 9 2 9 2 9 7 9 2
8 1 0 9 13 15 0 9 2
7 15 4 15 13 1 1 2
7 0 9 13 3 0 9 2
11 0 0 9 13 10 0 9 1 0 9 2
4 9 4 13 2
14 10 0 9 1 9 4 13 2 0 9 7 0 9 2
17 9 15 4 13 1 9 14 13 9 1 9 2 13 9 1 9 2
10 9 4 13 1 1 11 1 0 9 2
8 10 0 9 13 10 0 9 2
14 0 9 1 9 9 13 16 9 3 13 10 0 9 2
11 9 13 10 9 7 1 9 7 0 9 2
23 9 4 13 1 9 1 10 0 9 1 14 13 10 9 15 13 15 0 9 7 0 9 2
19 4 15 13 0 1 9 1 9 7 9 2 13 11 0 9 7 0 9 2
8 0 9 7 9 4 3 13 2
11 3 4 11 13 16 11 13 10 0 9 2
22 9 4 3 13 9 1 10 0 9 1 9 0 9 1 9 7 9 1 9 1 11 2
11 15 13 1 0 9 1 0 7 0 9 2
18 1 10 0 9 4 15 13 0 9 1 14 13 10 0 7 0 9 2
14 15 13 0 9 2 0 0 9 7 0 9 1 9 2
10 15 13 9 2 9 2 9 7 9 2
19 1 12 9 4 9 13 1 1 10 0 9 9 1 10 0 9 0 9 2
12 10 0 9 13 15 0 14 13 7 13 11 2
16 9 4 13 1 14 13 11 10 9 1 11 9 1 9 12 2
16 15 4 13 9 1 9 2 9 7 0 9 1 9 7 9 2
14 9 4 13 11 9 1 9 7 9 2 1 1 11 2
7 11 9 13 3 11 9 2
15 9 4 13 10 9 15 0 13 0 9 1 10 0 11 2
13 15 13 3 10 9 1 9 7 9 1 10 9 2
8 10 0 9 13 1 0 9 2
7 10 0 9 13 1 11 2
17 15 4 4 13 1 16 10 0 9 13 10 0 0 9 2 9 2
7 15 13 0 9 1 11 2
30 9 13 9 1 9 1 9 1 9 1 11 1 12 2 7 4 13 0 1 10 9 15 4 13 1 9 7 10 9 2
21 15 4 13 11 10 0 9 1 9 7 9 1 9 1 11 1 10 9 1 9 2
10 15 13 10 0 7 0 9 1 9 2
19 15 13 14 13 1 14 13 0 1 9 1 10 0 9 9 1 11 11 2
9 9 4 13 10 9 13 11 9 2
15 11 4 13 10 0 9 1 11 1 9 7 9 1 11 2
17 15 4 13 10 9 1 10 0 9 1 9 7 10 0 0 9 2
12 15 4 13 0 1 10 0 0 9 1 11 2
7 10 0 9 13 11 0 2
10 11 13 10 9 1 11 7 11 9 2
22 15 4 13 10 0 7 0 9 1 11 2 0 1 9 1 0 9 7 9 1 9 2
16 9 1 11 13 1 9 7 9 2 15 13 3 9 1 9 2
10 1 9 13 9 1 9 9 1 9 2
5 15 13 10 9 2
19 9 4 13 9 2 9 13 2 15 13 0 9 1 14 13 15 1 9 2
7 9 4 13 10 0 9 2
11 15 13 10 0 9 1 0 9 7 9 2
11 9 4 13 10 9 1 0 9 1 9 2
12 9 13 1 9 2 7 9 13 1 0 9 2
8 15 13 7 4 13 10 9 2
23 1 9 13 12 9 1 9 9 1 9 15 0 9 13 1 2 15 13 12 9 10 9 2
7 15 4 15 13 15 1 2
15 15 4 13 1 1 14 13 9 1 10 9 1 0 9 2
28 9 4 13 9 1 16 11 13 7 13 3 1 10 0 9 15 13 1 11 2 11 2 11 11 7 0 9 2
12 15 13 16 9 7 0 4 13 1 7 13 2
19 15 13 10 9 2 10 9 1 15 2 10 9 15 15 4 13 9 1 2
8 3 15 4 13 15 1 9 2
25 15 13 10 0 9 1 14 13 9 2 13 9 7 13 9 2 0 7 0 2 15 13 0 9 2
12 10 9 4 13 0 1 0 9 7 0 9 2
14 15 4 13 9 1 10 9 2 9 2 9 7 9 2
11 15 4 13 9 1 9 9 7 9 9 2
16 15 4 3 13 9 1 9 2 9 7 15 15 0 13 9 2
16 9 7 9 1 9 13 10 0 1 10 9 1 9 7 9 2
10 9 4 13 0 7 13 9 1 11 2
17 9 7 9 13 10 0 9 1 10 9 1 14 13 9 7 9 2
17 9 2 9 2 9 2 9 2 9 7 9 2 0 7 0 9 2
9 9 4 13 7 13 10 9 0 2
5 9 13 9 9 2
10 15 13 1 10 9 1 9 7 9 2
5 11 13 9 9 2
4 9 1 11 5
5 9 11 11 11 2
21 1 9 9 4 9 15 1 3 13 10 9 1 11 2 13 16 15 13 10 9 2
19 10 9 1 9 1 11 2 11 11 7 11 4 1 10 9 13 15 9 2
19 11 13 1 9 1 0 9 1 9 7 10 9 15 4 13 1 14 13 2
10 9 9 4 13 1 9 1 0 9 2
16 11 13 10 9 1 9 7 9 9 7 10 0 7 0 9 2
34 11 4 13 10 9 13 1 2 2 9 1 9 7 9 2 0 9 2 9 1 9 2 9 1 9 2 9 2 9 7 9 1 0 5
9 1 10 0 9 13 15 0 9 2
7 0 13 3 16 15 13 2
7 9 1 11 13 15 10 2
18 15 13 10 9 1 0 9 1 10 0 9 2 9 2 9 7 9 2
13 9 9 13 14 13 9 7 9 2 9 7 9 2
7 7 15 4 3 4 13 2
11 1 9 1 9 4 15 13 9 7 9 2
11 1 9 1 9 4 15 13 9 7 9 2
16 1 9 1 9 7 9 1 9 4 15 13 0 9 7 9 2
22 11 13 14 13 10 9 1 10 9 9 2 1 9 2 9 2 0 9 7 0 9 2
7 9 13 10 9 1 11 2
17 11 13 15 1 0 16 10 9 2 9 7 9 4 13 7 13 2
10 11 9 4 13 1 11 1 0 9 2
12 11 4 13 10 9 1 11 1 10 0 9 2
8 10 0 9 13 9 1 15 2
17 11 13 14 13 9 15 13 0 9 1 10 0 9 1 0 9 2
9 15 13 3 0 1 9 7 9 2
18 7 3 1 1 10 0 9 13 15 0 1 9 2 9 7 0 9 2
5 11 13 0 9 2
12 4 15 13 15 2 13 15 9 1 0 9 2
12 1 0 9 4 11 13 1 10 0 0 9 2
13 9 4 13 1 9 1 7 10 0 9 7 9 2
7 11 4 13 9 7 9 2
18 2 15 4 13 10 0 9 1 15 15 13 0 2 0 7 13 9 2
13 2 15 4 13 10 9 7 13 9 1 0 9 2
11 2 15 4 13 9 7 13 9 1 11 2
13 2 15 4 13 0 9 1 0 1 9 7 9 2
13 2 15 4 13 1 9 2 13 9 7 13 0 2
14 2 15 4 13 0 0 9 1 9 1 9 7 9 2
9 11 4 13 9 7 10 0 9 2
10 2 15 4 13 2 10 0 11 2 2
11 2 15 4 13 9 7 9 0 1 9 2
16 2 15 4 13 9 1 9 1 14 13 1 0 9 7 9 2
11 2 15 4 13 0 9 1 10 0 9 2
25 2 15 4 13 1 9 1 10 0 9 1 9 7 9 2 7 1 9 9 1 3 14 13 9 2
12 11 4 13 9 1 11 7 1 10 0 9 2
7 15 4 13 10 0 11 2
18 11 13 1 9 16 11 9 1 11 13 1 9 7 10 9 1 11 2
14 15 13 0 9 1 14 13 9 1 9 1 10 9 2
11 0 9 7 9 4 4 0 13 1 9 2
10 9 1 11 4 4 13 1 0 9 2
16 11 4 13 0 1 14 13 9 9 2 1 1 9 1 9 2
15 16 9 0 9 4 13 0 2 4 9 1 10 0 13 2
19 11 13 16 11 4 13 1 9 1 10 0 9 1 9 2 9 7 9 2
15 9 4 13 7 3 13 1 12 9 1 3 9 1 12 2
6 9 4 13 0 9 2
15 11 4 13 9 7 13 16 9 13 1 9 1 0 9 2
16 3 1 11 4 9 1 10 0 7 10 0 13 10 0 9 2
17 11 4 13 1 10 9 1 0 9 1 14 13 9 1 1 9 2
17 9 4 13 7 9 2 9 7 9 1 9 1 0 9 1 9 2
12 15 13 3 0 0 14 13 9 1 0 9 2
10 1 9 13 9 1 9 9 7 9 2
13 11 4 13 9 1 16 9 13 9 1 10 9 2
14 9 9 1 0 14 13 10 9 1 9 9 4 13 2
4 9 13 0 2
7 10 9 4 13 0 9 2
7 11 4 13 1 0 9 2
9 7 0 7 0 9 4 13 0 2
17 10 0 9 1 9 4 4 13 1 12 0 9 1 10 0 9 2
10 11 4 13 9 7 1 10 13 9 2
20 11 4 13 1 11 1 0 14 13 9 1 1 15 15 13 9 1 0 9 2
21 9 9 4 4 13 2 7 11 4 13 10 0 9 16 15 13 9 13 1 9 2
8 9 7 9 4 13 0 9 2
11 10 0 4 13 1 1 14 13 0 9 2
25 15 13 11 9 16 11 4 13 10 9 15 13 1 9 0 16 15 13 0 9 2 9 7 9 2
6 11 13 0 1 9 2
22 9 9 7 9 2 10 9 7 9 2 13 3 10 0 9 11 13 1 9 1 9 2
10 11 4 3 13 9 1 9 7 9 2
11 9 4 13 9 2 9 2 9 7 9 2
12 15 4 13 9 1 9 2 9 7 0 9 2
17 11 4 13 1 10 0 9 7 16 15 13 9 2 9 7 9 2
17 15 4 13 0 9 1 14 13 9 9 1 9 2 9 7 9 2
3 9 13 2
15 9 4 13 1 10 0 9 1 14 13 0 7 0 9 2
11 9 7 9 4 13 0 9 7 9 13 2
5 11 4 13 9 2
11 9 1 9 4 13 7 9 0 9 13 2
13 11 4 3 13 0 9 1 0 0 9 1 12 2
10 10 0 9 1 9 4 13 1 9 2
11 15 4 4 13 9 1 9 9 7 9 2
16 11 13 1 9 10 0 9 1 9 2 0 1 9 7 9 2
6 11 4 13 1 9 2
24 10 0 9 7 10 0 9 1 9 4 13 1 3 14 13 0 9 15 13 9 1 0 9 2
13 9 1 9 2 9 7 9 1 9 4 4 13 2
8 15 4 4 13 1 0 9 2
9 9 1 0 0 7 0 4 13 2
7 10 0 9 13 10 9 2
8 9 1 0 9 4 3 13 2
15 11 4 13 9 9 1 9 16 0 9 7 9 4 13 2
25 11 4 13 9 1 9 1 0 7 0 9 2 3 16 15 4 13 10 9 15 13 0 1 0 2
7 11 4 13 9 1 9 2
8 10 0 9 13 0 1 9 2
9 9 1 9 14 13 1 1 11 5
4 9 1 9 2
8 10 9 13 1 9 1 9 2
17 9 1 9 13 1 9 2 7 9 13 0 9 9 14 13 1 2
6 9 2 11 5 11 5
5 2 5 11 2 5
9 9 1 9 14 13 1 1 11 5
25 12 9 1 16 10 0 9 13 1 11 2 13 0 9 14 13 1 1 10 0 7 0 0 9 2
17 9 0 9 13 0 9 11 11 11 11 1 14 13 1 1 9 2
15 15 13 9 1 10 0 9 2 1 9 1 0 0 9 2
22 11 13 10 0 1 10 9 15 4 13 9 1 9 2 7 1 9 13 9 1 9 2
23 7 9 1 9 7 9 13 0 2 7 0 13 0 1 15 15 4 13 1 9 0 9 2
18 2 10 0 9 13 14 13 1 12 9 7 10 0 9 1 0 9 2
30 15 13 1 12 9 2 7 15 13 0 1 9 7 10 0 14 13 15 2 13 9 11 11 1 11 1 11 1 11 2
26 1 1 10 0 7 0 9 4 9 13 1 12 9 1 10 0 9 15 4 13 10 9 1 0 9 2
31 2 15 13 0 9 7 10 9 9 7 9 2 13 11 11 1 11 16 15 13 9 15 4 13 1 1 1 1 9 11 2
21 2 15 13 3 9 1 14 13 15 2 3 16 15 3 13 3 0 2 13 15 2
19 0 0 4 13 16 9 4 13 1 1 10 9 1 14 13 11 1 9 2
19 16 9 15 4 13 1 9 2 4 13 1 9 2 13 15 1 0 9 2
23 2 15 13 3 10 9 16 9 3 4 13 0 2 7 16 15 3 4 13 10 0 9 2
9 9 15 13 3 2 13 3 0 2
16 9 13 16 15 4 13 15 1 1 9 7 3 2 13 11 2
27 10 0 9 13 11 1 9 1 11 11 11 2 3 9 1 1 12 9 1 10 13 9 1 10 0 9 2
12 9 13 10 9 1 11 7 10 9 10 9 2
20 16 11 11 13 9 7 11 1 9 2 4 15 13 9 7 9 1 0 9 2
11 0 13 3 0 1 9 1 10 0 9 2
13 2 15 13 16 15 13 0 1 9 10 0 9 2
21 7 15 13 10 0 9 2 10 0 9 13 15 15 4 13 1 9 1 1 9 2
13 15 13 16 15 4 13 9 7 9 2 13 11 2
14 10 0 9 11 2 9 2 4 13 13 10 0 9 2
26 11 13 0 1 0 9 1 9 11 11 9 2 7 13 3 10 0 7 0 0 9 13 1 10 9 2
19 2 1 9 4 11 13 1 12 7 12 9 1 9 7 13 3 3 9 2
25 7 15 13 1 14 13 10 0 0 9 1 9 7 4 0 13 10 0 9 1 9 2 13 11 2
20 3 11 0 0 9 7 11 1 9 4 13 14 13 10 0 9 2 1 11 2
23 9 15 4 13 1 14 13 9 1 11 2 4 4 13 1 0 9 1 11 9 1 9 2
18 1 15 15 4 13 1 1 0 9 2 13 10 0 9 11 11 11 2
33 2 15 4 13 0 2 7 15 13 10 0 9 1 15 2 13 11 1 9 1 10 9 1 11 7 10 9 13 1 10 0 9 2
8 9 1 0 9 13 1 9 5
5 2 11 11 2 5
23 15 13 9 0 9 11 2 15 9 13 1 9 2 15 1 9 13 1 0 9 1 11 2
15 11 13 16 15 4 4 13 9 7 13 9 1 0 9 2
15 10 0 13 1 9 1 9 0 7 0 1 10 9 9 2
10 1 10 13 11 10 1 9 1 15 2
27 0 9 3 13 15 14 13 9 1 9 2 15 4 13 10 9 1 10 12 9 7 10 9 1 10 0 2
15 9 4 4 13 1 1 10 0 9 1 12 2 1 11 2
19 7 16 10 0 9 4 13 2 13 9 11 11 1 1 14 13 1 9 2
14 0 15 13 9 13 1 11 9 1 14 13 15 1 2
24 10 0 0 9 4 13 7 13 12 9 0 2 0 9 12 1 10 2 9 2 1 11 11 2
6 15 4 13 1 9 2
5 0 9 1 9 2
16 11 13 3 1 9 0 9 2 0 15 15 13 1 0 9 2
7 11 9 13 12 0 13 5
3 0 9 2
8 11 9 11 11 4 0 13 2
33 9 13 9 10 0 0 9 1 14 13 15 1 12 0 2 0 15 9 1 10 9 13 9 1 3 12 9 7 0 9 1 13 2
4 9 2 11 5
4 2 8 2 5
7 11 9 13 12 0 13 5
27 10 0 9 13 9 9 7 9 2 7 13 3 1 14 13 9 1 9 1 9 1 9 2 7 10 9 2
23 0 9 2 0 9 7 10 0 9 1 14 13 9 0 1 0 9 1 10 9 1 12 2
16 15 13 1 9 15 13 1 9 16 10 0 9 13 9 9 2
42 9 13 16 9 13 0 3 1 16 11 2 11 0 9 2 11 2 7 11 0 9 13 9 1 16 11 13 10 10 9 1 12 9 9 1 9 9 4 13 1 9 2
35 9 1 14 13 12 0 0 12 9 1 14 13 10 10 9 16 15 4 13 1 2 1 12 9 1 9 1 9 2 13 1 15 15 13 2
27 7 15 13 3 16 11 1 9 13 1 0 9 1 14 13 1 0 9 15 4 13 1 3 12 9 3 2
33 1 9 1 9 9 13 10 0 9 3 1 14 13 12 9 1 9 1 9 2 3 0 1 9 1 12 9 15 4 13 1 9 2
14 3 3 10 9 13 9 1 14 13 9 2 13 9 2
8 9 13 15 3 0 1 1 2
19 11 13 1 9 2 7 3 9 13 0 1 14 13 1 12 9 1 9 2
22 9 4 13 1 1 1 12 9 10 9 2 13 15 1 9 15 4 13 1 9 9 2
13 10 0 9 13 1 9 1 15 15 11 4 13 2
24 7 9 13 0 1 9 15 1 12 9 3 4 13 1 14 13 10 0 9 1 12 9 9 2
10 3 13 11 1 12 9 9 10 9 2
19 9 1 11 2 11 7 11 4 10 0 9 13 10 0 9 7 9 9 2
17 1 10 9 13 10 0 9 1 14 13 9 1 9 1 12 9 2
27 1 9 4 11 3 1 0 9 4 13 1 0 9 2 15 15 4 13 10 10 12 9 0 1 1 9 2
22 9 4 3 3 13 1 15 9 7 11 0 9 13 1 10 0 9 1 10 10 9 2
32 0 9 1 1 12 4 13 16 0 9 15 3 4 13 1 1 9 1 9 1 14 13 11 2 4 4 13 1 3 0 9 2
5 3 13 11 9 5
7 7 9 9 13 1 9 5
3 13 9 2
17 9 11 11 4 13 1 14 4 13 10 0 9 1 0 1 9 2
17 11 11 13 1 9 2 7 11 13 15 13 3 0 14 13 9 2
8 9 2 11 11 11 2 11 5
5 2 11 11 2 5
8 2 15 13 0 7 0 0 2
25 15 13 1 10 9 15 10 9 4 13 2 13 11 9 11 11 1 11 11 1 9 9 1 11 2
9 1 9 13 11 10 0 0 9 2
12 9 1 11 13 12 9 1 10 12 0 9 2
24 3 11 2 12 2 12 2 7 11 2 9 2 4 13 14 13 9 1 11 10 12 0 9 2
20 2 15 13 0 9 15 4 4 13 7 15 4 13 15 9 7 9 1 9 2
20 1 9 7 9 13 15 1 9 1 9 2 3 4 15 1 9 13 1 9 2
18 15 4 15 4 13 1 7 3 13 15 9 1 0 9 2 13 11 2
30 2 1 10 0 13 15 3 0 1 14 13 15 2 7 3 3 0 13 15 0 3 2 7 15 13 14 13 0 9 2
36 1 10 0 3 4 11 11 7 11 11 11 13 1 9 2 7 3 13 15 1 7 10 12 13 0 1 15 2 13 9 11 11 1 11 11 2
19 11 11 13 3 12 9 1 9 7 13 3 1 1 9 1 9 1 9 2
20 1 11 13 10 0 9 10 9 2 7 4 0 13 1 9 0 1 9 9 2
14 1 9 13 11 1 9 12 9 1 1 1 0 9 2
2 9 2
13 3 13 9 1 11 11 0 9 1 11 1 9 2
20 11 11 4 3 13 1 14 13 3 1 9 2 7 4 3 13 12 0 9 2
8 9 2 11 11 11 2 11 5
28 2 16 15 4 13 10 12 0 0 9 2 3 13 15 15 4 13 12 9 0 16 15 13 3 2 13 11 2
18 1 3 10 0 9 3 13 11 11 0 9 1 9 16 15 13 9 2
9 1 9 9 13 9 3 9 12 2
19 3 12 9 13 1 1 11 7 11 15 13 3 9 12 7 12 1 9 2
27 7 1 1 1 16 9 13 1 0 9 7 16 9 13 1 9 2 13 9 1 16 15 13 9 1 9 2
31 2 15 4 3 13 16 15 4 13 15 1 10 9 15 13 3 1 9 2 16 13 15 15 13 1 14 13 9 1 15 2
17 7 15 13 15 13 3 0 14 13 9 1 9 2 13 11 11 2
23 2 15 13 15 4 4 13 12 9 0 1 9 1 16 15 4 13 9 1 14 13 9 2
34 11 2 11 7 11 13 3 0 1 16 15 13 15 13 3 0 9 1 9 16 15 4 13 10 9 1 10 1 15 2 13 9 11 2
5 0 9 1 11 5
5 2 5 11 2 5
4 9 1 11 5
20 11 11 2 12 2 13 15 10 0 9 1 9 1 9 9 1 10 0 9 2
4 6 2 11 2
9 11 11 4 0 13 9 1 9 2
4 9 2 11 5
13 9 2 15 4 13 1 11 2 13 1 10 9 2
19 0 13 11 12 9 1 9 2 7 15 13 1 12 9 9 1 11 11 2
16 1 12 9 7 12 9 1 9 4 15 0 13 1 10 9 2
8 1 9 13 15 9 1 11 2
10 2 15 13 9 1 14 13 1 9 2
16 9 4 13 0 9 1 15 16 15 4 13 3 2 13 11 2
26 11 7 11 13 9 1 12 9 3 14 13 2 7 11 13 0 1 9 1 9 12 2 12 7 12 2
5 3 13 11 9 5
3 1 9 2
16 1 9 4 11 13 1 15 10 0 9 15 13 1 9 11 2
5 9 2 11 11 5
5 2 11 11 2 5
22 15 13 0 9 16 11 7 9 11 2 12 2 13 9 1 11 11 11 11 1 11 2
42 16 15 13 9 1 0 12 9 1 9 1 9 2 13 15 0 15 13 9 1 16 9 7 9 9 2 15 10 9 1 9 13 9 11 2 13 0 0 2 13 11 2
10 15 15 4 13 1 10 9 0 9 2
28 10 9 1 10 0 9 13 3 1 11 16 11 13 9 1 7 13 15 1 9 2 1 9 1 0 1 9 2
16 1 0 9 13 15 9 1 9 2 15 4 13 1 1 0 2
2 9 2
12 9 13 1 10 12 9 9 1 9 7 9 2
6 9 13 9 11 9 2
7 9 13 1 9 1 9 2
5 9 2 11 11 5
12 3 1 9 1 9 0 9 13 9 1 9 2
15 1 9 13 11 3 0 1 1 9 16 9 4 13 1 2
20 16 15 13 1 16 9 4 4 13 2 4 15 13 1 10 0 9 1 9 2
34 2 15 13 10 9 15 13 1 14 13 9 2 7 15 4 13 0 9 1 15 2 13 11 11 11 15 13 9 1 11 1 11 11 2
11 15 13 11 4 13 9 1 0 9 1 2
17 2 15 13 0 14 13 7 9 7 9 9 1 9 2 13 11 2
5 9 13 0 9 5
5 2 11 11 2 5
18 0 9 3 0 1 9 4 13 3 0 9 1 9 2 11 12 2 2
20 10 9 13 15 3 13 2 7 13 15 2 3 0 16 15 3 13 0 2 2
7 3 13 9 3 0 0 2
3 13 3 2
8 2 11 2 9 1 0 9 5
21 10 0 9 2 11 11 2 2 15 13 0 9 2 13 9 9 1 10 0 9 2
21 15 4 3 13 9 1 10 9 7 1 9 7 9 2 7 9 1 9 1 9 2
21 15 13 2 11 12 2 9 0 0 9 2 7 1 10 9 4 15 13 0 0 2
3 13 3 2
10 3 13 2 11 11 8 11 2 9 5
30 11 11 4 13 1 0 1 11 12 7 11 12 2 3 15 4 13 15 1 9 9 1 0 11 11 11 7 11 11 2
14 11 7 11 9 4 13 16 9 13 1 0 1 11 2
24 3 15 13 1 10 0 9 4 15 3 13 1 0 7 0 9 1 9 9 1 10 0 9 2
10 13 15 1 10 9 15 13 1 9 2
6 13 10 9 1 11 2
7 0 9 1 9 1 11 5
2 0 2
13 9 11 11 13 15 13 0 1 10 9 1 11 2
4 9 2 11 5
5 2 5 11 2 5
7 0 9 1 9 1 11 5
18 9 1 10 0 9 1 11 13 0 1 16 10 9 13 0 7 0 2
7 9 11 11 13 9 0 2
18 1 9 12 9 1 9 11 1 1 11 13 15 1 9 1 9 9 2
12 15 13 9 1 0 9 7 13 9 1 9 2
7 9 13 1 9 7 9 2
15 9 1 9 13 0 0 7 0 0 9 13 0 1 9 2
16 9 4 3 13 9 1 2 9 2 7 2 9 2 1 9 2
14 15 13 1 9 15 0 9 3 13 1 9 1 11 2
13 10 10 9 13 1 11 1 11 1 10 9 3 2
32 1 9 1 11 4 15 3 13 2 11 2 2 9 1 10 0 9 15 13 9 3 1 10 0 9 1 11 1 12 9 3 2
13 9 15 13 2 13 1 14 4 4 13 1 9 2
18 11 13 1 10 9 16 15 13 2 0 2 16 15 13 9 1 9 2
11 2 9 13 0 7 13 3 1 1 11 2
22 15 13 10 9 15 13 1 9 1 11 2 15 13 9 7 9 0 0 2 13 9 2
10 3 9 11 11 13 9 1 10 0 2
24 2 10 9 1 0 9 13 10 0 7 0 9 15 15 3 4 13 1 9 1 2 13 15 2
16 9 1 9 13 15 13 0 9 1 9 1 9 15 13 1 2
10 2 15 13 0 16 0 9 13 15 2
26 1 1 1 10 0 9 15 13 2 4 15 3 4 13 14 13 9 2 13 10 1 9 1 9 11 2
22 1 10 9 1 9 2 11 11 2 13 10 0 9 9 15 1 1 9 9 1 9 2
20 9 7 9 4 4 13 0 9 2 7 9 13 15 10 2 3 0 9 2 2
17 1 9 1 9 4 15 3 4 4 13 2 9 2 2 1 11 2
4 9 1 11 2
7 2 13 3 9 1 9 5
8 11 4 13 12 9 1 9 5
4 13 1 9 2
12 12 9 13 9 1 9 1 11 2 1 11 2
5 9 2 11 11 5
5 2 11 11 2 5
33 15 13 11 15 1 9 4 13 16 15 13 12 9 1 0 9 9 7 11 13 9 1 9 2 16 11 9 2 11 2 4 13 2
7 12 9 13 9 1 9 2
31 11 11 2 9 1 11 11 2 11 2 2 13 15 1 16 15 13 0 9 1 9 16 15 13 0 9 9 12 1 9 2
28 2 1 10 9 13 15 11 10 9 14 13 11 2 7 15 4 3 13 1 16 15 13 9 0 2 13 11 2
6 1 11 13 15 9 2
10 12 13 9 0 9 1 9 1 9 2
19 9 13 3 9 1 1 11 10 9 0 2 3 12 2 3 4 9 13 2
12 11 13 14 13 1 1 0 7 13 3 1 2
15 3 13 7 9 7 11 9 16 15 13 9 0 1 9 2
19 12 13 11 9 1 16 15 13 9 1 9 1 9 2 7 13 11 0 2
10 11 13 3 9 1 9 13 1 9 2
16 2 15 13 3 0 9 15 13 1 9 1 9 2 10 9 2
23 1 0 13 15 1 9 7 3 13 15 1 14 13 11 2 16 15 13 9 2 13 9 2
12 0 11 11 2 12 2 13 1 9 1 9 5
3 0 9 2
13 9 1 9 4 11 11 13 1 10 9 1 11 2
10 15 13 3 0 15 15 13 1 9 2
8 15 13 10 0 9 1 9 2
4 9 2 11 5
5 2 11 11 2 5
19 9 1 9 4 11 13 1 15 15 0 13 0 9 1 9 11 1 11 2
31 3 13 0 11 11 11 2 12 2 2 13 1 0 9 1 11 9 2 1 15 15 13 1 10 0 9 16 11 4 13 2
19 15 13 16 10 1 9 4 4 13 11 7 13 15 1 1 9 1 9 2
10 1 9 13 10 9 15 13 15 1 2
14 9 4 4 13 9 3 9 16 9 13 9 1 11 2
8 0 9 13 1 1 0 9 2
19 2 15 13 3 1 9 1 9 1 9 2 9 15 13 7 9 15 13 2
15 15 13 1 9 2 7 16 15 13 1 13 9 3 1 2
12 3 13 11 11 11 1 9 10 1 9 11 2
4 9 2 11 5
26 9 11 2 15 13 1 11 1 10 0 9 2 13 10 9 7 13 10 0 9 1 10 0 7 0 2
10 3 13 0 9 16 9 4 0 13 2
12 2 0 9 13 1 11 1 9 3 1 9 2
10 10 0 0 9 13 0 0 1 9 2
14 15 13 1 11 3 2 13 11 11 1 10 0 9 2
17 10 0 9 13 14 13 9 2 7 15 13 9 1 9 7 9 2
22 9 11 11 13 9 4 13 1 9 1 10 9 1 14 13 1 9 2 13 11 11 2
14 9 13 15 0 1 16 9 13 0 15 4 13 9 2
9 9 4 4 13 11 1 9 11 2
18 11 11 2 9 1 11 9 1 9 2 13 15 13 0 14 13 9 2
14 2 15 13 0 7 3 0 1 15 14 13 1 9 2
15 3 13 15 1 1 0 9 2 13 11 1 1 11 11 2
15 3 13 0 7 0 9 0 1 14 13 11 1 1 9 2
2 0 2
17 3 13 10 0 9 9 1 9 1 9 11 3 11 11 4 13 2
4 9 2 11 5
14 2 10 9 4 13 15 15 13 1 14 4 13 11 2
23 9 13 1 15 1 1 7 15 13 0 0 0 2 13 9 1 9 1 11 2 11 11 2
17 9 11 13 3 0 1 9 3 12 9 4 13 0 9 1 9 2
33 9 11 7 11 11 13 1 9 1 1 11 7 13 10 12 9 1 11 11 11 2 15 13 3 12 9 1 9 1 10 0 11 2
12 11 11 4 13 7 13 2 16 9 4 13 2
18 15 13 14 4 4 13 1 9 15 13 15 0 1 0 9 1 11 2
4 11 1 11 5
5 2 5 11 2 5
26 11 11 11 13 9 1 11 11 11 16 9 13 11 11 12 2 12 1 10 9 1 10 0 9 9 2
2 13 2
19 11 11 11 13 1 10 1 11 11 11 0 9 16 9 13 1 11 9 2
4 9 2 11 5
13 15 13 9 15 13 9 1 10 9 1 0 9 2
18 11 11 13 0 1 9 16 11 13 9 1 9 12 1 12 1 9 2
15 11 11 2 11 11 7 11 11 13 10 10 9 1 11 2
13 9 13 12 9 7 13 10 0 9 1 11 9 2
16 0 13 1 16 3 11 11 13 10 12 9 1 11 1 11 2
8 9 13 11 0 11 1 11 2
12 9 13 11 10 9 1 11 11 11 1 11 2
15 2 15 13 14 13 15 2 13 9 11 11 0 1 9 2
16 11 0 9 11 11 13 10 9 1 9 7 9 12 1 9 2
10 15 1 14 13 10 0 9 11 11 2
13 11 13 1 10 0 1 9 1 11 1 10 9 2
8 11 13 11 13 9 1 9 5
9 2 15 13 3 11 1 14 13 5
4 13 1 9 2
17 3 13 0 11 11 1 9 15 4 13 2 16 9 1 11 13 2
7 9 2 11 11 2 11 5
5 2 11 11 2 5
3 2 0 2
2 0 2
2 0 2
24 13 15 1 10 9 16 11 13 10 9 0 2 2 2 13 9 11 11 1 10 9 9 9 2
22 2 15 13 1 9 1 11 2 7 15 13 0 9 1 15 2 13 11 1 11 11 2
33 16 11 2 15 13 10 9 1 9 1 9 1 11 10 9 2 13 1 9 1 9 1 11 9 2 13 9 0 1 0 1 9 2
9 9 11 11 13 9 1 0 9 2
27 2 16 15 13 0 4 15 0 13 9 1 10 9 1 9 2 7 15 4 13 0 3 0 9 1 10 2
18 4 15 13 10 9 16 15 13 10 9 15 4 13 1 11 9 3 2
12 2 15 13 10 9 2 7 15 13 0 0 2
10 7 15 4 3 13 1 15 0 9 2
9 15 13 0 2 15 4 13 15 2
14 7 10 0 13 1 9 2 11 10 9 2 11 11 2
2 13 2
23 9 1 11 11 2 11 11 2 13 0 1 11 9 9 1 9 1 11 7 11 1 11 2
7 9 2 11 11 2 11 5
35 11 13 15 13 1 1 11 14 13 1 16 11 13 0 9 1 14 13 9 1 9 2 7 13 3 1 9 1 16 9 4 13 10 9 2
32 2 13 15 9 1 10 1 11 0 9 2 3 4 15 13 9 1 15 2 3 1 9 2 7 0 16 15 13 15 1 9 2
38 16 15 13 1 10 9 15 15 13 2 4 15 3 13 15 9 16 15 4 13 1 2 7 13 10 10 13 10 10 9 2 13 15 2 7 13 1 2
18 2 9 13 0 9 2 7 15 4 13 3 15 9 9 15 4 13 2
5 15 13 10 9 2
19 7 0 13 13 15 1 15 15 13 1 2 7 4 13 1 1 0 9 2
15 7 15 13 0 0 1 10 9 15 13 1 3 0 0 2
27 1 0 9 1 11 11 1 16 11 13 14 13 1 11 11 11 10 9 1 9 2 13 9 10 9 0 2
8 2 6 2 15 13 15 3 2
16 15 13 15 3 0 2 7 13 16 15 13 10 9 1 9 2
9 3 4 15 13 2 13 11 11 2
7 1 11 0 9 13 11 2
16 2 11 11 4 13 16 15 13 15 15 13 1 2 13 11 2
12 11 13 9 1 11 2 7 3 0 11 9 2
31 2 15 13 3 7 0 16 7 11 7 11 13 0 9 1 15 2 7 15 13 1 10 9 15 15 4 4 13 7 13 2
5 15 13 0 0 2
4 13 9 3 2
23 3 11 11 11 11 2 15 3 4 13 9 1 10 9 3 2 13 0 0 1 9 9 2
7 2 15 13 15 13 0 2
12 15 9 13 10 9 7 13 0 9 1 9 2
8 11 11 13 10 9 15 13 2
15 15 13 3 1 10 9 2 13 15 1 11 9 9 9 2
12 3 9 1 11 7 9 9 13 1 9 9 2
35 2 15 4 4 13 10 9 9 15 4 13 1 9 7 15 13 9 15 13 0 1 9 1 15 15 13 2 13 9 11 11 1 11 9 2
6 2 15 13 0 0 2
21 15 13 0 9 1 10 9 2 13 11 11 2 0 9 1 11 2 1 11 12 2
7 3 13 9 15 13 0 2
5 2 15 13 9 5
5 2 15 13 0 2
23 10 0 9 2 3 2 13 1 14 4 13 11 11 2 12 2 1 9 1 11 1 11 2
6 9 2 11 11 11 5
5 2 11 11 2 5
7 3 13 0 9 11 11 2
19 10 9 4 1 0 9 13 9 1 9 2 7 13 16 15 4 13 9 2
8 15 4 3 13 1 10 9 2
31 2 15 13 16 15 13 1 7 13 10 0 9 0 9 2 13 1 9 7 3 13 1 9 1 10 0 13 2 13 11 2
10 9 1 9 13 1 11 9 9 9 2
8 9 4 0 13 1 0 9 2
14 2 15 13 10 0 9 1 14 13 0 1 10 9 2
25 15 13 15 13 3 0 1 9 9 16 15 3 13 10 9 1 14 13 15 10 9 2 13 11 2
17 9 7 9 4 13 16 3 10 9 4 4 13 1 16 9 13 2
25 9 13 16 9 1 9 2 7 16 9 1 9 3 13 3 0 1 10 0 9 2 13 9 9 2
16 15 13 3 16 9 4 13 10 9 15 3 13 0 1 11 2
9 0 13 1 1 10 0 9 9 2
16 10 0 9 4 13 16 15 13 1 1 9 0 1 9 12 2
9 15 4 3 13 16 9 13 9 2
31 9 11 11 13 16 15 13 0 16 10 0 9 4 13 9 2 16 9 13 12 9 0 2 16 10 0 9 13 12 9 2
14 9 13 10 9 1 10 9 9 12 7 9 9 12 2
12 15 4 3 4 13 1 1 11 9 9 12 2
41 1 9 13 15 0 0 16 15 13 9 1 14 13 1 1 9 2 13 10 9 2 4 13 2 13 9 2 13 1 1 9 7 13 15 1 9 3 1 10 9 2
12 9 13 10 9 1 16 15 13 9 1 9 2
7 0 13 15 13 1 9 2
12 9 13 16 9 1 9 3 13 15 1 9 2
24 0 13 15 1 14 13 15 10 9 1 9 2 7 10 9 2 3 16 15 3 13 0 3 2
13 10 9 13 10 0 9 2 3 13 15 0 9 2
6 15 13 0 1 0 2
5 13 9 13 0 5
4 13 1 9 2
9 1 9 13 3 9 1 0 9 2
10 9 4 13 1 9 1 11 11 11 2
4 9 2 11 5
5 2 11 11 2 5
18 11 9 13 1 9 10 9 3 9 11 11 15 13 1 10 10 9 2
15 9 4 13 1 10 9 16 15 13 1 1 9 0 9 2
21 1 9 1 9 13 11 16 9 11 11 13 1 9 1 11 0 12 9 0 9 2
17 15 13 9 15 13 11 11 1 9 1 12 0 9 15 13 15 2
12 9 4 3 13 3 0 15 13 9 1 9 2
8 11 0 9 13 1 0 9 5
15 11 13 9 10 0 9 1 10 0 9 1 10 0 9 2
2 9 2
12 1 0 9 1 11 13 11 11 10 0 9 2
7 3 13 15 10 0 9 2
4 9 2 11 5
24 9 15 4 13 9 13 1 10 0 9 9 2 7 13 9 1 11 11 1 9 1 10 9 2
25 1 9 13 10 2 0 0 9 2 1 9 1 9 15 13 9 1 9 1 9 2 9 7 9 2
35 2 10 0 9 11 11 13 0 0 1 10 0 9 7 13 0 0 9 2 13 15 1 9 2 3 9 13 1 9 16 15 13 0 11 2
13 15 13 3 0 9 10 0 9 4 13 1 9 2
15 1 10 4 15 4 13 16 9 9 13 1 11 11 9 2
23 10 0 9 13 11 2 15 0 13 1 12 9 2 1 10 9 11 11 2 0 9 2 2
21 11 13 0 9 2 7 9 13 0 9 1 10 0 9 2 9 7 9 0 9 2
25 1 1 1 10 9 9 3 13 0 15 13 10 0 1 11 11 2 15 3 3 13 10 0 9 2
41 1 9 13 15 3 16 11 13 10 0 9 1 0 9 3 16 15 13 12 9 2 7 16 15 1 9 3 13 12 9 10 9 7 0 13 9 1 9 1 9 2
23 2 10 0 9 11 11 13 15 1 9 2 9 1 9 1 0 9 2 13 15 1 9 2
6 0 9 13 1 11 5
4 9 7 9 5
16 2 0 1 11 4 13 1 9 7 9 1 9 1 1 9 2
11 15 13 3 3 10 0 9 2 13 11 2
2 9 5
23 2 15 13 16 9 1 0 9 13 0 1 9 1 0 9 2 7 16 15 13 10 9 2
19 15 4 13 0 14 4 13 1 15 1 10 9 1 10 0 2 13 11 2
3 13 9 5
5 11 13 12 9 5
5 2 11 11 2 5
17 2 1 9 1 10 0 0 9 2 3 13 1 11 1 9 2 2
25 10 0 9 1 11 1 11 13 10 1 9 1 9 15 13 1 1 0 9 1 0 9 1 9 2
2 9 2
20 9 11 11 1 11 4 13 9 1 14 13 10 9 15 4 13 1 1 9 2
11 3 13 15 1 9 1 10 9 1 11 2
6 9 2 11 11 11 5
3 1 9 2
21 10 0 9 9 4 13 3 1 9 1 10 0 9 1 11 1 9 1 0 9 2
6 9 2 11 11 11 5
3 0 9 2
19 9 11 11 7 9 11 11 1 11 13 1 9 1 9 1 11 1 11 2
6 9 2 11 11 11 5
20 3 9 1 9 1 9 7 11 13 9 14 13 1 1 0 9 1 0 9 2
22 1 3 4 15 13 1 9 1 9 2 9 2 9 7 10 9 0 9 1 12 9 2
18 10 1 15 15 13 14 13 10 9 1 9 1 9 13 11 1 11 2
25 0 9 1 9 13 15 1 9 10 2 10 9 1 10 0 9 11 2 1 9 1 10 0 9 2
6 1 10 13 0 1 2
25 0 9 13 1 9 10 2 1 9 1 16 15 4 13 0 1 9 1 9 15 13 9 1 11 2
15 2 15 4 13 0 14 13 3 9 4 13 1 10 9 2
33 15 4 13 0 9 2 13 11 11 2 15 1 0 9 4 13 1 14 13 7 13 10 0 9 2 15 3 4 13 0 1 11 2
20 1 0 9 1 9 13 15 14 13 1 9 7 9 1 9 1 10 0 9 2
11 0 1 9 13 9 1 14 4 13 1 2
22 9 11 11 13 16 7 9 7 11 4 13 1 9 1 10 0 9 9 1 11 13 2
30 2 10 0 9 15 13 13 16 15 13 1 9 1 11 7 13 16 15 13 12 9 1 9 7 13 2 11 11 2 2
16 3 13 15 16 15 13 0 2 3 1 11 9 2 13 15 2
26 9 11 11 11 13 15 4 13 0 9 1 14 13 10 10 9 15 4 13 1 7 1 9 7 9 2
15 0 1 9 13 1 9 15 4 13 9 13 7 13 9 2
17 10 4 13 3 0 0 9 1 9 1 0 9 2 9 7 9 2
17 1 9 13 10 0 9 9 15 4 13 1 10 0 9 1 9 2
22 11 13 16 9 1 9 3 13 10 9 1 10 10 0 9 15 13 1 9 1 9 2
23 1 9 13 10 9 1 0 9 15 13 0 9 1 9 16 10 0 9 1 11 13 0 2
22 2 10 0 15 13 16 15 13 3 1 9 1 1 11 0 9 13 9 9 11 11 2
8 3 1 13 11 9 11 11 2
22 15 13 0 9 16 15 15 3 4 13 9 13 9 1 14 13 10 9 2 13 15 2
11 11 13 0 9 1 9 1 10 0 9 2
16 2 15 4 13 0 1 10 0 9 2 3 15 13 1 15 2
25 0 9 1 9 13 1 9 16 9 13 0 2 7 15 4 13 1 1 10 0 9 2 13 15 2
14 9 13 15 13 0 14 13 10 0 9 1 1 11 2
28 2 15 13 10 0 9 2 7 15 13 3 0 16 15 4 13 0 1 14 13 15 1 11 9 2 13 15 2
20 11 9 4 13 1 1 12 9 1 9 2 9 2 9 7 0 9 1 9 2
14 12 9 2 10 9 7 9 4 13 10 9 1 11 2
43 9 13 1 0 0 9 1 11 11 2 11 9 11 11 7 11 9 11 11 2 1 9 1 11 2 11 11 2 9 1 10 0 9 1 11 7 0 9 1 11 7 11 2
22 11 4 3 13 9 1 11 0 9 1 11 2 9 7 0 0 9 1 1 1 9 2
24 15 13 9 1 11 15 4 13 9 1 14 13 9 7 13 1 16 15 4 13 1 10 9 2
9 10 9 4 3 13 1 9 10 2
16 2 15 4 13 9 1 9 1 11 7 9 7 9 1 11 2
25 1 9 4 9 1 0 9 13 9 1 9 1 11 2 13 9 11 11 1 11 9 1 11 11 2
4 0 1 1 5
12 9 1 11 9 13 12 9 0 1 1 9 2
8 10 0 9 1 11 13 0 2
20 2 4 15 13 1 11 4 15 13 0 1 9 2 13 11 11 2 12 2 2
22 15 13 1 11 11 1 11 2 15 13 10 9 1 11 16 9 4 13 14 13 0 2
17 10 9 13 1 11 11 1 9 1 11 4 13 14 13 12 9 2
18 10 9 1 11 9 1 11 1 4 3 13 1 14 13 12 9 0 2
23 2 15 13 0 9 2 7 15 4 13 15 13 9 2 13 11 11 2 12 2 1 11 2
3 0 9 5
18 11 11 13 15 1 9 1 14 13 11 15 13 3 1 9 1 11 2
33 9 1 3 0 10 9 4 13 14 13 1 9 7 9 1 11 4 13 10 0 12 9 2 13 0 9 1 11 9 2 11 2 2
23 0 9 13 10 9 9 10 0 4 13 14 13 2 7 13 10 9 1 9 1 10 9 2
8 2 15 13 0 9 1 11 2
28 10 0 9 1 9 13 0 1 1 12 9 3 2 13 9 11 11 1 11 9 1 9 7 9 2 11 2 2
3 9 13 5
11 11 13 10 9 1 1 7 1 1 9 2
9 15 13 1 15 12 9 1 11 2
18 1 0 9 15 13 15 1 9 9 2 13 9 1 9 7 9 0 2
7 2 15 13 1 10 9 2
32 10 9 1 9 4 13 10 0 9 2 7 1 1 1 15 13 10 0 9 9 1 9 1 9 2 13 9 11 11 1 11 2
17 15 13 1 0 9 7 9 0 1 9 1 10 0 9 1 9 2
19 2 16 15 13 1 13 11 10 0 0 9 2 7 15 4 13 10 9 2
23 3 13 15 0 0 9 3 2 15 13 16 15 3 13 10 9 9 1 9 2 13 11 2
5 13 0 1 1 5
10 9 1 9 13 0 0 1 1 1 2
19 1 9 13 10 9 1 9 1 12 9 1 9 2 13 11 9 1 12 2
8 1 1 13 9 1 12 9 2
9 9 1 11 13 3 10 0 9 2
10 9 13 0 1 9 16 9 13 0 2
17 9 15 13 1 9 2 13 11 11 2 11 2 11 7 11 11 2
19 15 13 3 10 9 16 9 13 0 2 13 9 1 11 9 9 1 12 2
14 2 15 13 3 9 13 1 9 2 13 9 11 11 2
9 2 7 15 13 15 3 0 9 2
18 0 9 13 3 0 9 0 0 14 4 13 2 13 11 11 1 11 2
3 0 9 5
11 9 1 9 1 11 13 0 1 1 9 2
22 0 11 2 11 7 9 11 13 15 1 9 2 7 13 10 12 9 1 0 0 0 2
28 10 9 1 0 9 13 11 2 11 7 11 2 16 3 12 9 13 9 1 1 0 9 2 13 9 1 11 2
25 10 1 9 13 16 9 1 9 13 0 2 7 1 12 9 1 10 0 1 9 13 1 12 9 2
8 2 11 13 11 0 0 9 2
36 15 13 0 14 13 16 1 1 1 10 9 1 9 10 0 4 13 2 3 4 9 1 9 7 9 13 2 13 9 11 11 1 11 1 11 2
7 11 1 14 4 13 1 2
6 2 15 13 1 13 5
3 0 9 5
3 13 9 5
6 13 9 1 0 9 5
5 2 11 11 2 5
21 16 11 11 11 2 12 2 13 1 14 4 13 0 2 13 0 0 1 1 9 2
7 15 4 3 4 13 9 2
3 1 9 2
22 10 0 11 11 11 4 13 16 15 13 1 7 13 15 1 9 16 9 4 13 9 2
4 9 2 11 5
22 15 13 9 1 10 9 1 16 15 4 13 1 1 9 7 1 1 9 1 9 9 2
12 2 15 13 16 15 3 13 10 0 1 15 2
8 15 13 16 15 13 1 13 2
25 3 3 3 3 0 1 9 2 7 10 9 9 2 13 10 1 11 9 11 11 11 1 11 11 2
9 2 15 13 0 1 9 1 11 2
9 13 15 9 1 15 16 15 13 2
11 2 6 2 15 13 3 15 2 13 15 2
16 15 13 1 12 0 2 0 7 9 1 9 1 9 1 9 2
21 3 12 1 15 13 1 1 9 2 16 9 13 9 1 9 1 10 9 1 9 2
30 15 13 1 16 11 13 10 9 1 3 15 13 15 3 4 13 1 9 1 9 7 9 1 11 16 9 1 9 13 2
14 11 13 15 13 0 7 13 16 11 4 13 15 9 2
13 16 11 13 1 1 9 13 15 9 1 10 9 2
13 1 9 13 9 11 11 16 15 13 10 0 9 2
26 11 11 11 13 16 11 13 16 15 4 13 15 16 15 13 15 1 9 1 9 3 16 9 4 13 2
22 2 15 13 16 15 13 14 13 10 0 9 1 14 13 10 9 15 13 2 10 0 2
20 15 13 0 0 16 15 3 4 13 10 9 1 3 15 13 2 13 11 11 2
8 2 15 4 13 1 10 9 2
14 2 6 2 15 13 15 0 0 1 16 15 3 13 2
12 15 13 10 10 9 9 13 1 10 0 9 2
21 1 9 13 11 9 11 11 11 1 14 4 13 12 9 1 3 15 3 13 9 2
19 2 1 9 4 11 13 16 15 4 13 15 15 4 13 7 13 1 9 2
10 15 13 15 0 1 2 13 11 11 2
19 15 13 16 11 4 13 15 1 9 9 1 14 13 1 9 1 11 9 2
33 16 11 0 1 9 1 9 1 0 13 1 9 2 13 15 16 15 13 10 9 1 11 11 7 11 11 9 15 13 15 0 0 2
10 1 9 13 11 10 9 2 0 2 2
28 2 15 13 0 0 1 16 15 13 14 13 1 9 2 7 15 13 0 9 15 13 9 9 2 13 11 11 2
14 2 4 15 13 15 1 3 15 13 14 13 10 9 2
13 2 6 2 15 13 0 0 1 15 2 13 9 2
14 9 13 10 9 1 9 1 11 1 9 1 0 0 2
17 2 0 13 15 16 15 4 13 0 9 1 15 2 13 11 11 2
16 1 9 15 13 0 9 4 15 13 1 12 9 1 11 9 2
11 15 13 1 9 0 1 9 1 10 9 2
22 1 7 1 1 9 4 15 0 13 9 1 9 1 9 15 0 4 13 0 1 15 2
2 9 2
5 9 15 13 11 5
3 13 0 5
2 9 5
4 13 1 9 5
4 11 13 3 5
11 10 0 9 4 13 14 13 0 9 1 2
4 9 7 9 2
9 15 4 3 13 10 0 9 3 2
11 10 9 4 9 11 13 1 12 9 9 2
10 9 10 13 9 1 10 9 1 9 2
5 15 13 15 3 2
12 11 4 13 1 14 4 13 0 9 1 9 2
18 14 13 1 9 15 13 1 10 0 7 0 9 2 13 10 0 9 2
15 11 4 13 16 15 13 2 3 16 15 13 15 15 13 2
13 3 13 15 16 9 1 11 4 13 9 1 11 2
13 15 13 0 9 1 0 0 9 1 0 0 9 2
16 7 15 13 16 9 4 13 3 2 7 13 9 1 0 9 2
14 15 13 3 9 1 16 0 9 13 10 9 1 11 2
9 9 1 9 4 13 1 0 9 2
20 0 9 2 1 9 1 10 9 9 2 4 13 9 1 9 1 9 1 11 2
15 0 9 15 13 1 0 0 9 2 4 13 1 10 9 2
16 15 13 0 14 13 1 9 9 1 10 0 0 9 1 9 2
8 1 11 13 0 9 10 9 2
15 15 4 13 2 3 1 9 10 2 1 10 9 1 9 2
25 1 9 1 10 0 9 13 10 10 9 3 2 15 13 15 1 1 9 2 7 13 9 1 9 2
5 10 13 0 9 2
12 7 10 0 9 1 11 13 10 9 1 9 2
11 11 13 3 9 1 9 9 1 0 9 2
17 1 9 1 11 1 0 12 9 3 2 13 9 1 1 0 9 2
9 0 1 9 4 13 0 1 15 2
14 15 13 0 9 1 16 0 9 13 1 1 0 9 2
17 9 13 14 13 10 0 0 1 10 0 10 15 13 0 1 9 2
10 10 0 4 15 13 0 14 13 1 2
15 10 10 4 13 1 2 7 13 1 1 10 10 7 0 2
8 8 8 8 2 13 9 15 2
7 9 13 1 10 0 9 2
10 15 13 0 1 0 1 9 7 9 2
13 15 13 15 3 13 10 12 9 2 15 15 13 2
22 10 12 9 13 9 1 0 7 0 2 7 15 13 1 9 1 9 2 9 7 9 2
8 9 13 1 7 9 7 9 2
10 9 13 0 2 7 13 9 1 9 2
8 3 10 9 2 3 0 9 2
10 3 10 0 9 13 1 9 1 9 2
10 9 1 0 9 13 3 2 9 1 2
11 10 9 4 3 4 13 1 10 0 9 2
15 3 1 0 9 4 15 13 9 2 9 7 9 1 11 2
10 10 10 9 4 4 13 2 0 0 2
12 11 13 2 1 9 2 14 13 0 10 9 2
6 15 13 1 0 9 2
5 0 4 15 13 2
16 9 4 13 15 2 16 15 0 13 1 9 1 14 13 9 2
11 7 0 4 9 4 13 3 0 15 13 2
25 1 10 9 15 9 11 3 4 4 13 16 15 13 10 0 9 2 16 9 13 0 10 0 9 2
19 15 13 0 9 1 14 13 1 10 9 1 9 2 1 9 7 1 9 2
8 10 9 16 9 13 0 9 2
17 11 4 4 13 9 1 14 13 10 10 9 15 10 13 0 1 2
3 0 3 2
18 7 16 15 13 15 10 9 2 13 15 0 0 9 1 10 10 9 2
13 15 13 1 10 0 9 15 4 13 10 0 9 2
16 1 10 9 15 15 4 13 1 9 2 7 1 10 0 9 2
10 16 15 13 9 2 4 15 0 13 2
20 7 15 4 4 13 2 7 15 4 4 13 3 0 15 13 1 10 0 9 2
16 15 4 13 15 1 1 9 2 7 15 4 13 15 15 13 2
9 3 3 4 15 13 15 1 9 2
17 15 13 0 0 9 1 16 0 9 13 1 9 1 10 0 9 2
7 0 9 13 0 1 9 2
22 7 16 15 13 10 9 15 4 13 1 9 2 7 16 15 10 4 13 0 7 0 2
13 15 4 1 10 13 10 0 7 0 9 1 11 2
13 9 4 13 10 9 3 3 9 13 0 15 1 2
23 15 13 15 13 1 14 13 0 1 11 2 1 10 16 0 13 16 15 3 4 13 0 2
14 13 4 15 2 4 11 4 13 1 14 13 0 9 2
19 11 2 11 0 0 9 2 4 3 4 13 1 0 9 1 9 7 9 2
33 15 4 13 0 1 15 15 4 13 1 15 15 13 3 2 7 1 15 15 4 13 1 10 0 9 2 15 15 13 3 1 1 2
25 15 13 0 1 10 9 16 10 0 0 9 15 13 10 9 1 10 0 9 2 13 3 11 11 2
15 15 13 15 13 15 1 16 9 1 11 3 13 3 0 2
14 16 15 13 0 15 13 10 0 9 9 10 13 1 2
17 16 15 0 7 0 13 0 1 9 14 13 0 9 1 9 10 2
15 9 2 9 7 9 4 13 14 13 1 1 0 9 10 2
14 16 15 13 1 9 2 4 15 13 15 1 9 9 2
8 7 15 4 13 15 1 9 2
9 11 9 13 11 13 9 1 9 5
4 13 11 11 5
6 2 4 3 13 9 5
5 2 11 11 2 5
29 1 10 9 1 9 11 13 9 11 9 10 9 1 10 9 7 10 0 9 1 16 9 4 13 1 9 1 9 2
2 9 2
19 9 11 11 13 3 9 2 7 13 3 9 11 9 13 1 9 1 9 2
6 9 2 11 11 11 5
4 9 2 11 5
31 1 9 13 9 1 10 0 9 11 16 9 4 13 1 9 1 15 15 13 2 7 3 1 9 1 9 15 4 13 1 2
14 11 4 1 9 13 1 9 1 1 10 9 11 11 2
26 2 7 9 13 0 16 9 13 1 9 15 3 13 10 9 1 2 0 9 2 2 13 15 1 9 2
2 9 2
4 9 1 15 2
36 9 13 3 1 10 9 15 13 1 14 13 0 1 9 16 9 13 2 7 13 1 11 11 7 11 11 1 10 9 1 1 10 9 11 11 2
17 2 15 13 0 14 13 16 9 3 13 1 9 16 9 4 13 2
12 11 11 13 16 9 13 1 15 11 13 0 2
15 11 11 7 11 11 13 0 16 11 13 15 1 11 11 2
16 3 13 15 15 13 16 9 13 1 9 9 2 13 15 0 2
29 9 11 11 11 13 16 15 4 13 0 1 10 9 14 13 9 1 9 1 10 9 9 11 4 13 9 1 9 2
23 2 15 13 0 3 10 2 0 2 9 1 10 9 2 7 13 15 1 15 1 0 9 2
20 15 10 13 3 0 0 9 1 10 9 7 10 9 2 13 11 1 11 11 2
24 15 13 3 11 11 1 9 2 7 13 16 9 3 4 13 9 1 14 13 10 9 1 11 2
16 2 15 13 16 0 9 13 15 7 0 7 9 4 13 3 2
17 7 15 4 13 11 11 1 9 3 2 15 13 0 15 13 9 2
20 0 9 13 10 9 1 15 1 10 9 2 7 1 0 1 9 2 13 11 2
15 2 11 13 3 10 0 2 0 9 2 15 13 0 9 2
14 3 13 15 10 9 3 1 0 9 7 10 9 0 2
10 16 15 13 0 7 0 2 13 15 2
25 9 13 16 11 13 9 1 9 1 11 2 7 13 16 9 3 13 15 1 15 15 13 1 11 2
22 2 3 13 15 10 0 9 3 1 11 2 7 3 10 9 1 14 13 9 1 11 2
16 3 10 9 1 9 1 11 7 10 9 2 13 15 1 9 2
15 11 11 13 9 4 13 9 1 9 11 7 9 1 9 2
20 2 9 4 13 1 15 16 15 3 13 9 2 7 11 15 13 9 1 11 2
17 7 16 11 13 10 9 4 10 0 9 2 13 11 2 13 0 2
11 15 13 10 0 7 0 9 2 13 9 2
17 15 13 3 1 15 15 13 10 2 15 2 1 2 15 2 9 2
12 2 15 13 3 9 15 15 13 1 10 9 2
29 15 0 9 13 0 0 9 3 9 2 0 2 9 2 9 2 9 7 3 0 4 13 9 1 9 2 13 15 2
7 3 13 15 9 0 9 5
3 0 9 5
4 0 0 9 5
2 9 5
3 0 9 5
3 9 0 5
4 0 1 9 5
4 11 1 9 5
5 0 1 9 10 5
3 9 11 5
5 11 2 11 2 5
12 1 0 9 2 1 0 9 2 13 10 9 2
10 15 13 1 9 7 9 1 9 10 2
4 9 7 9 2
24 9 11 11 2 12 2 1 11 13 0 1 14 13 0 1 9 1 14 13 0 9 1 11 2
10 15 13 9 7 9 1 9 1 11 2
6 9 2 11 11 11 2
3 0 9 2
16 9 11 1 11 11 13 0 9 1 9 7 9 1 9 11 2
6 9 2 11 11 11 2
2 9 2
26 9 11 13 0 9 2 3 9 4 13 1 9 7 13 0 9 1 3 9 7 9 13 1 1 11 2
6 9 2 11 11 11 2
2 11 2
12 9 1 11 13 10 0 9 1 0 7 0 2
11 1 1 9 13 0 7 0 9 7 13 2
6 9 2 11 11 11 2
4 9 1 11 2
18 9 13 1 9 11 1 11 2 3 10 1 12 9 0 9 4 13 2
13 9 13 1 9 7 9 1 9 15 13 1 9 2
6 9 2 11 11 11 2
3 9 11 2
15 11 11 2 12 2 1 9 1 9 15 4 13 1 12 2
16 15 13 9 1 1 11 1 14 13 2 13 9 7 0 9 2
6 9 2 11 11 11 2
3 9 9 2
13 11 11 11 2 12 2 13 9 11 11 1 11 2
18 15 13 16 0 0 9 13 14 13 1 11 1 9 1 14 13 1 2
6 9 2 11 11 11 2
14 9 13 11 11 2 12 2 1 9 1 10 0 9 2
18 9 9 2 9 7 9 13 9 1 15 1 14 13 10 0 1 9 2
18 15 13 3 0 16 11 9 11 11 10 9 13 0 0 9 1 11 2
31 1 11 2 1 9 7 9 2 13 10 9 1 11 2 11 0 7 0 9 1 0 9 2 3 0 9 11 13 10 9 2
38 2 15 13 0 0 1 9 2 1 3 0 9 7 0 9 15 15 13 3 2 13 11 11 16 15 13 15 1 9 7 13 9 1 10 9 1 9 2
9 15 13 0 1 0 7 0 9 2
8 15 13 9 1 10 0 9 2
11 2 3 13 15 14 13 2 13 15 0 2
6 3 1 13 15 1 2
10 0 9 0 13 15 0 9 7 9 2
13 9 9 13 11 1 7 9 2 9 7 1 9 2
17 15 4 13 2 13 1 9 2 13 7 13 1 0 7 0 9 2
24 9 13 10 1 9 1 2 11 0 0 9 2 2 10 9 15 13 1 11 1 11 1 12 2
48 10 1 11 0 9 13 10 9 15 1 10 13 0 16 2 15 0 9 13 9 0 1 14 13 10 0 0 9 2 15 1 9 1 10 9 7 9 4 13 15 1 10 0 9 1 9 2 2
26 9 13 0 9 1 0 9 2 7 3 0 13 0 9 1 9 2 1 11 1 11 7 11 1 11 2
19 11 9 13 11 11 2 11 2 15 13 1 11 11 2 1 9 1 9 2
13 3 13 15 9 1 9 7 0 9 0 1 9 2
21 1 9 4 9 7 9 13 1 11 0 2 11 7 9 2 1 0 11 11 11 2
21 1 0 9 3 13 0 1 11 0 13 9 1 14 13 9 2 9 9 7 9 2
21 13 15 1 0 9 2 13 15 3 9 2 9 7 0 9 2 16 15 13 0 2
10 1 9 13 9 0 0 0 7 0 2
18 1 11 4 15 13 9 1 9 1 9 2 1 14 13 9 3 0 2
10 3 4 15 13 1 1 10 0 9 2
14 1 9 13 10 9 0 10 10 11 1 10 0 9 2
17 3 4 15 13 1 9 7 13 0 9 15 13 3 9 13 1 2
25 3 13 15 1 1 9 1 9 3 9 13 1 9 2 7 4 13 3 9 13 1 10 0 9 2
10 9 1 11 13 1 10 0 9 11 2
23 3 13 9 1 10 0 9 3 9 13 2 3 16 9 13 0 0 0 7 0 1 9 2
13 9 13 1 9 1 11 7 11 2 10 0 11 2
21 9 13 3 0 1 9 1 9 2 3 9 1 9 2 9 7 9 13 1 9 2
26 1 9 13 10 9 1 0 9 7 1 0 2 0 9 1 1 9 1 10 1 9 0 9 2 11 2
19 10 1 12 9 0 9 13 1 9 10 0 9 1 0 9 7 0 9 2
12 0 9 7 9 13 1 0 9 9 0 9 2
24 9 3 13 0 16 10 0 9 4 13 1 9 0 9 7 0 0 9 1 11 11 1 12 2
16 1 11 7 11 2 7 3 0 1 0 9 1 11 7 11 2
18 10 9 1 1 12 9 0 9 1 0 9 13 12 9 1 0 9 2
15 9 1 9 13 9 9 1 9 2 0 9 7 0 9 2
10 9 1 11 13 0 1 3 9 13 2
22 15 13 1 0 9 1 12 9 1 9 2 7 13 7 9 2 9 2 9 7 9 2
18 0 9 13 15 3 0 14 13 1 1 9 2 7 9 13 12 9 2
13 9 13 3 0 1 1 9 2 7 9 13 9 2
39 15 13 15 10 9 1 9 1 11 7 11 2 3 1 10 9 1 9 7 9 1 10 12 15 13 0 3 2 11 2 12 2 7 11 11 2 12 2 2
12 9 13 1 12 9 7 13 12 9 12 9 2
9 16 15 13 0 9 13 10 9 2
15 2 15 13 10 9 3 0 15 13 2 13 9 11 11 2
14 15 13 3 9 15 13 2 7 16 15 13 0 9 2
6 7 9 13 3 3 2
11 1 1 11 13 15 1 1 10 0 9 2
10 3 4 10 0 0 9 13 10 9 2
39 7 16 9 11 11 2 12 2 13 10 0 9 1 9 2 7 16 2 11 2 0 13 1 9 1 9 7 9 1 14 13 1 9 2 13 7 13 9 2
17 0 13 9 1 10 9 13 1 15 15 4 13 1 1 9 1 2
16 9 13 1 1 0 9 2 0 9 7 0 9 1 0 9 2
13 3 4 15 3 13 15 1 0 9 3 0 9 2
7 2 15 13 3 3 9 2
7 15 13 9 1 10 9 2
9 0 15 13 0 2 13 15 0 2
9 1 9 13 11 15 1 0 9 2
11 15 1 0 1 10 0 1 9 7 9 2
13 9 7 9 4 3 13 10 0 9 1 0 9 2
17 10 1 9 0 9 13 1 9 11 11 2 0 0 1 1 9 2
24 3 13 15 9 0 9 1 9 2 7 1 9 9 12 1 9 1 9 13 15 3 15 13 2
18 11 11 11 2 12 2 13 1 9 2 1 0 9 7 9 1 9 2
9 15 13 15 15 13 7 13 9 2
12 11 13 10 9 1 11 2 7 13 1 3 2
14 2 15 4 13 1 16 0 9 13 14 13 1 11 2
22 15 13 0 1 9 10 2 7 15 4 13 1 16 3 3 0 13 3 2 13 11 2
2 3 2
20 11 13 10 9 1 12 9 15 13 1 1 11 2 3 3 1 11 7 11 2
8 9 13 10 0 9 1 11 2
18 1 9 1 12 9 13 3 2 1 15 1 12 1 7 1 9 11 2
2 9 2
21 0 11 11 13 0 1 11 1 11 9 1 11 12 9 1 9 2 9 7 9 2
5 0 9 1 9 2
13 13 15 10 10 9 1 9 2 13 15 1 11 2
10 9 1 11 13 10 7 10 0 9 2
17 9 13 2 7 13 1 1 12 9 2 12 9 9 9 1 11 2
13 4 15 13 9 2 13 11 11 1 11 1 11 2
2 3 2
12 10 0 9 1 15 15 13 9 7 0 9 2
29 15 4 13 0 1 16 15 4 13 12 9 1 10 9 2 0 9 2 9 7 9 2 7 15 13 3 0 0 2
2 13 2
18 0 9 1 9 1 11 2 1 0 9 2 1 0 9 1 0 9 2
6 15 13 1 11 11 2
