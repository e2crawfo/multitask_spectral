605 11
20 13 3 15 16 16 0 13 15 9 3 10 9 7 9 3 3 13 1 9 9
3 6 13 15
13 13 7 3 13 16 15 15 13 9 13 15 9 9
14 3 1 9 15 13 16 3 13 12 9 0 7 0 13
13 10 13 15 13 7 10 13 1 15 13 15 3 13
12 13 3 15 0 3 9 15 10 1 9 0 13
7 6 13 15 16 13 9 15
9 13 9 15 3 1 9 3 1 9
8 13 3 9 15 16 13 9 13
12 16 3 9 10 1 15 9 13 10 9 3 3
11 7 15 15 13 13 13 1 9 15 9 12
10 13 7 3 9 15 10 1 9 16 13
13 3 13 9 0 9 0 13 7 9 0 9 0 13
19 15 3 15 13 9 15 7 13 0 13 15 9 0 15 13 9 15 1 9
6 7 13 9 13 15 13
4 15 13 13 15
6 3 1 11 0 9 13
5 7 13 7 13 15
9 9 13 15 3 13 7 13 9 15
5 7 13 1 15 11
9 13 7 3 3 15 9 9 0 13
10 7 13 1 9 13 7 13 1 15 9
10 15 13 3 0 13 13 15 9 7 13
5 7 13 13 1 15
7 3 3 13 13 0 7 0
8 3 3 7 9 13 7 9 13
8 7 11 13 15 7 13 0 13
12 7 13 11 3 13 1 15 12 0 13 7 13
5 13 16 9 3 13
5 3 13 1 9 15
5 3 3 13 15 15
20 15 3 15 13 15 1 9 9 13 3 15 15 1 9 9 15 15 1 9 13
13 10 13 15 15 13 7 10 15 13 13 10 13 15
17 0 13 7 0 13 0 0 13 7 0 13 7 0 13 7 0 13
1 9
8 15 3 9 7 9 1 11 13
9 13 10 9 9 13 7 13 7 13
16 3 16 1 11 13 9 10 13 1 15 3 15 13 1 0 9
7 3 13 3 10 1 0 9
4 3 13 15 13
3 15 15 13
2 15 13
4 3 13 0 9
3 7 15 13
23 7 13 12 12 0 9 10 13 15 13 1 9 11 7 13 15 1 9 9 3 13 15 9
13 7 3 13 15 1 3 15 9 16 13 10 9 3
8 13 3 1 10 9 7 13 15
2 15 13
16 7 13 1 9 1 9 15 13 1 10 0 9 7 13 15 0
15 0 3 9 15 13 1 9 13 0 9 7 9 1 11 13
4 13 7 3 13
12 13 11 9 1 9 7 13 9 9 1 9 9
10 15 13 9 15 10 0 1 15 3 13
9 7 3 13 10 9 15 13 1 15
4 15 15 7 15
16 15 0 9 10 0 16 1 9 3 9 10 0 13 7 13 15
13 7 3 9 13 13 7 13 1 0 9 7 3 13
11 7 11 13 13 9 15 13 15 7 13 15
7 7 13 3 1 11 1 9
7 15 13 13 9 3 12 9
6 7 15 9 13 1 15
6 7 13 11 13 1 15
15 7 13 9 16 13 1 15 0 9 7 3 13 1 0 9
5 7 15 13 1 15
9 7 13 1 10 9 10 13 13 9
28 7 11 13 1 9 15 1 9 7 3 9 1 11 13 1 15 7 1 11 7 1 9 7 1 11 7 3 11
17 7 11 10 11 7 11 9 11 7 13 15 9 11 15 13 9 9
12 7 16 9 1 15 13 3 13 13 10 9 0
5 7 13 1 15 9
9 7 15 10 9 1 9 1 9 13
24 7 15 13 1 9 0 7 13 9 13 7 13 7 13 12 12 7 12 12 7 12 12 7 13
27 7 0 13 3 10 1 0 13 15 16 13 0 9 3 1 9 13 15 7 3 13 9 1 15 7 0 13
6 16 15 13 9 13 13
15 0 3 9 9 13 3 9 3 9 3 9 9 1 0 9
3 13 0 9
8 7 13 10 9 7 13 9 0
30 3 15 3 9 1 9 13 7 9 0 13 13 7 13 1 15 0 9 7 10 1 9 9 13 7 9 3 13 15 13
3 15 9 15
10 13 3 3 3 12 12 7 13 1 9
3 7 15 13
12 7 3 11 13 1 15 15 10 1 15 9 13
5 9 9 15 13 15
5 7 13 13 1 15
7 7 3 13 10 9 7 13
8 7 3 13 9 15 3 1 15
10 3 3 13 1 9 3 13 16 13 3
12 13 3 11 13 16 15 15 9 13 11 0 13
4 7 13 15 16
10 7 3 13 0 9 9 13 13 9 15
60 7 13 15 10 9 15 0 9 0 13 13 13 9 7 9 7 15 9 16 3 13 9 3 13 13 9 10 0 7 1 9 16 13 3 13 7 0 13 0 15 13 1 13 9 9 7 9 7 9 7 9 3 3 13 15 10 9 7 10 9
6 13 9 15 7 9 15
10 7 10 13 1 9 0 13 10 13 9
8 10 15 0 3 13 7 13 9
4 7 13 1 15
7 7 13 15 16 9 3 13
3 7 13 15
6 7 13 9 9 12 9
10 7 13 15 13 3 1 9 13 1 9
12 9 13 3 13 7 9 13 3 13 7 3 13
15 7 13 1 11 7 13 1 15 0 7 13 15 16 15 13
11 7 13 11 7 9 15 1 9 11 10 11
3 15 13 11
8 15 3 13 9 15 13 13 15
16 7 9 15 13 13 0 3 9 0 3 9 1 9 3 13 13
2 0 13
7 7 3 13 13 1 9 9
15 7 3 3 15 13 13 15 7 13 7 13 9 15 7 13
6 7 13 1 9 13 13
4 15 0 10 13
8 7 11 13 15 1 9 13 15
4 7 13 1 11
12 7 15 15 15 13 3 15 13 7 10 13 15
26 7 15 15 13 12 0 0 10 13 1 15 0 13 15 3 16 13 9 1 9 15 7 13 13 1 9
7 7 16 9 13 13 3 13
6 7 13 11 13 1 15
8 3 13 1 15 9 16 13 15
5 7 15 13 1 15
6 13 9 15 7 9 15
5 13 3 13 9 0
5 13 1 15 11 13
19 13 7 3 1 9 13 1 11 7 13 13 15 11 7 13 7 13 0 13
6 7 11 13 3 1 15
7 7 15 13 15 13 1 15
5 9 11 11 13 15
9 7 15 13 9 15 13 13 1 11
20 7 16 1 13 11 1 11 7 11 1 9 0 13 12 9 15 7 13 1 15
16 7 13 10 9 1 11 7 13 1 15 9 15 7 13 1 15
13 7 13 9 3 13 9 13 16 3 13 15 1 15
5 7 13 13 1 15
6 9 6 9 15 13 13
5 7 13 3 1 11
6 7 13 1 15 3 13
6 7 13 11 13 1 15
12 3 0 13 7 0 0 15 13 15 7 3 13
10 13 7 13 10 9 7 13 10 9 0
10 9 13 16 0 13 7 3 9 15 15
1 9
3 7 0 3
10 15 13 9 11 7 9 11 7 9 11
3 0 0 9
7 7 15 3 3 13 15 13
3 13 1 9
3 7 15 13
4 9 10 9 13
4 15 13 0 13
9 7 13 12 9 15 13 7 1 15
1 13
9 7 15 13 9 1 15 7 13 15
9 7 15 13 10 9 0 13 1 15
12 15 13 9 10 0 7 1 12 9 0 0 13
2 15 13
1 13
9 7 1 0 3 10 13 13 1 11
24 7 3 1 9 9 13 10 0 9 1 10 0 7 9 7 15 10 9 13 11 13 15 1 11
9 7 11 3 9 3 13 16 13 11
9 15 3 13 16 13 15 13 9 9
3 0 9 9
8 13 7 3 9 0 7 13 15
8 0 13 7 15 15 3 13 13
3 6 11 13
35 7 3 1 9 13 16 13 9 15 13 0 9 13 11 1 11 0 9 15 13 3 15 13 9 9 13 13 3 1 11 7 13 10 9 11
9 15 13 15 10 9 1 9 10 9
1 13
12 7 15 13 16 13 7 13 13 1 15 3 13
6 7 9 10 13 0 13
1 6
6 13 3 1 15 10 9
18 15 13 11 10 13 1 9 9 7 13 13 13 1 15 7 13 15 0
8 7 13 3 10 9 1 15 13
16 0 13 0 7 9 0 13 7 13 15 9 9 9 11 9 15
5 13 15 1 9 15
12 13 9 15 9 7 13 9 15 1 9 9 15
17 13 11 9 15 13 9 3 13 1 9 15 11 7 9 15 1 9
9 13 3 9 15 10 3 13 13 15
11 7 11 9 15 13 9 0 7 13 7 13
11 13 3 16 0 13 3 13 9 1 13 15
12 9 1 9 9 7 1 9 9 1 9 0 9
48 7 16 13 9 9 15 1 9 11 13 15 1 11 13 1 9 3 13 13 1 9 9 16 15 0 13 9 0 9 13 7 16 13 1 15 9 3 13 13 1 9 9 9 9 7 12 0 9
14 6 0 13 1 9 7 9 0 1 11 7 1 9 13
12 7 13 10 9 15 9 15 1 11 1 9 9
4 7 13 1 15
4 9 13 1 9
12 13 3 15 16 13 9 1 9 0 13 9 11
4 3 13 1 15
15 13 9 1 9 15 7 13 9 15 7 13 9 1 9 15
5 7 13 1 15 9
5 7 13 15 11 13
18 7 13 15 11 1 9 9 1 11 7 9 13 1 15 9 13 1 15
8 0 9 13 9 0 1 9 15
30 7 1 9 13 15 16 0 9 13 1 9 11 1 11 16 13 9 1 9 12 7 9 12 16 13 9 0 1 15 9
1 13
14 15 9 0 16 1 9 7 9 13 10 0 9 7 13
5 15 13 11 9 9
7 16 3 13 13 13 1 11
8 13 1 15 16 9 0 13 9
1 13
7 7 9 9 13 1 13 15
5 15 13 1 9 15
16 7 1 0 13 7 13 9 9 11 13 1 9 7 13 1 15
5 7 15 13 1 15
14 3 13 10 0 9 10 9 7 0 13 7 10 9 13
15 3 0 13 15 13 11 16 0 13 15 7 15 1 15 13
5 13 3 11 1 15
52 7 16 13 9 13 9 15 7 13 1 15 12 15 3 9 13 11 15 7 13 11 7 11 9 15 11 7 11 11 7 11 11 7 11 11 10 11 7 11 10 13 11 11 11 7 11 11 15 7 13 13 15
13 13 1 0 9 7 13 16 6 9 15 0 1 9
5 3 13 10 13 15
12 7 16 9 13 10 9 13 15 15 15 9 13
4 13 7 13 15
23 7 3 13 13 1 9 15 9 13 15 13 9 10 1 9 15 0 1 9 15 9 3 13
14 0 13 9 13 9 15 13 7 13 7 13 9 1 9
10 7 15 13 1 11 13 15 3 13 16
7 7 13 1 0 13 7 13
27 16 3 1 13 9 10 9 3 6 13 13 9 9 0 9 15 7 15 0 9 7 9 10 9 0 1 15
5 7 13 15 9 15
19 1 7 3 0 9 13 0 1 9 7 9 7 9 0 7 0 0 13 9
11 6 10 1 9 0 7 9 13 1 9 13
9 7 10 0 1 9 9 0 15 13
8 13 9 9 13 7 13 7 13
5 11 13 15 15 13
5 3 15 13 1 15
6 7 15 9 13 9 15
4 9 15 13 15
4 0 3 13 13
7 7 0 1 9 13 10 13
15 13 3 1 15 9 7 9 15 7 3 13 13 15 1 9
5 3 3 3 13 13
12 15 13 0 16 7 9 13 7 9 7 13 15
5 13 3 15 11 13
26 13 3 13 10 13 7 13 1 11 7 13 13 10 9 1 15 9 13 13 7 13 1 9 11 7 13
5 13 3 15 13 15
4 15 10 13 15
14 3 15 13 13 15 9 1 10 9 9 13 1 15 16
7 3 13 16 3 13 7 13
11 7 13 15 13 9 9 7 13 15 10 0
13 11 15 9 13 7 15 13 0 1 15 15 13 0
4 13 15 15 13
9 7 13 13 15 13 15 9 9 12
33 7 15 3 13 15 13 16 9 3 13 0 13 16 13 9 9 0 13 7 13 1 0 13 7 9 7 9 7 13 7 0 9 13
18 13 3 1 0 9 3 9 12 13 11 7 11 7 11 13 1 9 13
7 7 9 13 1 10 9 13
10 7 13 9 15 16 13 15 7 3 13
15 7 15 3 13 0 9 7 13 13 1 15 16 3 13 15
5 7 13 1 15 11
5 3 13 15 9 13
2 13 15
5 13 3 1 15 11
5 3 15 1 9 13
10 7 13 10 1 15 0 7 13 1 15
10 7 15 11 15 1 9 13 1 9 13
10 7 13 1 16 9 15 13 13 1 9
9 7 6 9 15 13 13 15 7 13
4 0 13 7 13
13 3 15 15 13 15 0 13 7 15 13 15 15 13
8 9 15 13 9 0 7 13 0
8 9 9 13 12 7 13 13 0
8 9 13 3 13 7 3 9 13
30 7 15 9 13 13 1 0 9 1 9 15 3 13 3 13 13 3 0 1 12 12 13 10 1 12 12 12 13 1 15
13 7 13 9 7 9 13 16 0 0 13 7 13 15
13 3 13 15 9 13 1 9 9 9 1 12 13 0
13 7 13 0 13 9 15 13 9 7 9 15 3 13
5 7 13 15 10 9
10 7 13 13 1 9 7 13 9 7 9
12 9 15 3 1 15 13 7 15 10 15 15 13
9 15 13 16 9 15 13 9 1 15
9 13 15 9 7 13 3 13 12 12
4 7 15 15 13
12 13 3 10 15 3 10 9 0 13 7 13 15
7 7 0 15 13 9 13 11
21 3 16 12 9 1 9 13 1 15 7 12 9 1 9 13 15 13 13 15 13 15
5 7 3 13 1 15
5 7 15 13 9 13
4 7 10 12 3
4 13 3 1 9
6 7 13 9 7 13 15
9 7 15 1 9 3 3 13 15 0
4 7 15 13 15
3 13 3 9
18 9 13 15 16 3 13 3 10 0 9 9 0 9 7 3 3 0 9
5 7 11 13 15 13
3 10 9 13
5 3 12 15 9 13
3 7 15 13
18 7 15 3 9 0 13 7 13 10 9 0 1 15 7 3 13 10 13
8 13 3 11 13 15 13 1 15
7 7 15 9 13 13 9 9
11 7 13 15 13 13 16 1 0 9 13 13
13 13 3 12 9 15 13 15 12 9 7 13 1 15
4 7 13 0 13
9 1 9 15 13 15 0 9 7 0
18 7 3 9 15 0 15 3 13 15 13 1 15 13 3 7 13 1 15
4 3 13 10 9
5 9 13 10 9 15
5 9 15 9 9 13
9 13 15 3 15 12 9 7 13 15
9 3 15 15 13 1 15 9 0 13
6 13 3 10 9 10 9
10 13 7 13 9 0 7 13 10 9 0
8 13 3 16 1 15 0 9 13
3 13 3 13
5 7 0 13 0 3
11 7 16 13 0 3 11 13 1 9 16 13
7 7 0 11 13 1 9 9
5 1 15 3 0 13
6 7 0 13 15 13 13
7 3 13 9 9 3 12 12
11 7 9 3 13 7 3 13 3 1 15 11
20 3 16 13 9 16 11 13 3 7 9 15 13 1 9 7 13 1 11 13 11
6 15 13 16 13 9 9
4 6 6 13 15
16 15 15 13 15 9 1 15 13 7 10 13 1 15 3 13 3
5 3 13 1 15 3
5 15 13 10 9 9
4 6 6 13 15
7 3 0 13 10 9 15 13
7 7 13 15 15 15 3 13
4 9 9 0 13
8 13 7 3 3 9 9 10 9
6 3 13 10 9 13 15
6 15 3 13 16 0 13
21 16 15 13 9 15 13 13 1 10 9 1 7 9 13 7 15 3 1 15 15 13
6 13 11 7 13 1 15
13 3 3 1 9 13 10 9 16 0 13 1 9 11
10 11 16 13 3 0 9 13 15 0 13
13 13 15 7 3 13 7 3 13 15 15 3 13 13
3 0 13 11
4 3 3 13 15
5 13 7 13 1 15
6 13 11 7 13 1 15
6 3 15 13 7 9 15
7 3 15 13 15 3 13 13
6 9 16 3 13 1 15
6 0 15 13 0 13 15
9 10 3 9 3 13 1 9 1 9
7 16 9 11 13 9 11 13
12 3 3 3 1 15 15 3 13 7 15 15 13
7 16 9 13 3 3 13 15
4 6 6 13 15
2 13 11
6 3 13 10 9 1 15
12 9 15 13 0 3 7 9 15 16 0 13 13
12 3 9 7 10 13 15 3 16 15 9 13 13
12 9 13 11 9 13 7 13 15 9 7 13 15
9 3 3 13 15 7 10 9 3 13
9 15 15 13 1 0 16 13 15 9
15 7 3 3 13 3 13 7 15 13 15 10 9 15 3 13
13 13 3 0 9 10 9 15 13 0 7 13 1 15
2 13 15
19 13 7 3 16 9 0 3 13 7 16 15 9 13 7 9 15 13 0 13
8 3 15 13 9 16 13 1 15
5 3 3 15 0 13
19 0 9 13 7 10 9 9 15 13 7 10 0 9 13 1 9 7 13 0
4 15 13 10 9
9 3 0 9 13 15 3 13 0 9
3 15 0 13
3 13 15 11
9 13 3 9 10 9 16 13 1 15
33 16 0 13 9 1 15 9 9 13 7 3 13 13 13 10 13 15 9 13 7 13 1 10 9 15 13 16 13 16 13 9 9 13
19 13 3 3 11 15 13 9 9 7 13 9 15 9 15 15 9 11 0 13
5 13 1 15 10 9
5 3 13 10 9 15
11 13 3 11 13 15 3 12 9 13 1 9
3 13 9 15
15 6 9 15 13 16 15 13 11 9 9 10 1 10 9 13
2 7 13
11 3 11 3 13 1 15 15 13 1 10 9
6 13 3 10 9 3 13
5 13 15 7 13 13
16 13 3 12 10 9 15 11 11 10 11 15 13 15 1 13 15
23 0 9 9 3 15 13 1 9 13 16 13 11 1 11 13 9 9 7 13 13 15 7 13
7 3 10 9 13 1 15 3
4 6 6 13 15
6 7 3 13 1 0 9
5 3 9 13 0 9
7 3 0 9 9 1 15 13
19 13 15 9 7 13 15 9 16 3 13 9 7 13 9 7 13 7 13 15
10 3 3 13 16 13 9 7 16 13 9
3 9 7 9
4 15 13 15 13
11 3 13 1 15 3 10 9 13 1 15 13
5 13 3 1 15 11
7 9 3 0 9 1 15 13
3 7 3 13
7 1 9 9 15 9 0 13
8 15 13 10 9 7 9 7 9
5 15 13 15 13 9
5 3 15 1 9 13
10 7 15 13 15 16 15 13 7 15 13
12 7 10 9 15 13 13 15 7 10 13 15 9
11 16 13 15 3 15 13 16 15 13 1 9
9 15 9 1 15 13 9 0 13 15
14 1 0 13 13 9 15 16 9 0 13 7 13 15 9
8 3 9 3 13 15 13 15 9
6 16 15 13 3 15 13
3 13 15 3
14 7 3 13 1 10 13 15 7 15 1 15 3 13 15
13 7 1 9 16 1 9 15 13 7 3 3 13 15
9 3 13 1 10 9 15 1 15 3
9 9 16 13 9 13 16 13 9 15
17 1 0 9 1 9 15 13 7 3 13 15 16 15 13 9 1 15
2 3 13
23 13 15 9 16 9 15 13 15 3 13 15 9 15 9 16 15 15 13 15 13 15 9 0
4 15 1 15 13
5 15 13 15 9 15
15 7 15 9 15 13 15 13 15 16 13 12 3 15 12 13
19 7 11 13 9 7 10 9 7 9 9 13 7 0 1 9 7 9 7 9
5 3 3 15 3 13
18 7 11 11 13 9 13 15 7 13 10 0 9 9 7 13 15 9 0
15 10 3 9 13 0 10 9 7 13 1 11 1 9 10 9
13 7 10 0 9 13 11 1 9 15 7 1 9 15
3 13 15 11
7 13 15 10 9 10 0 9
5 13 7 13 1 15
2 13 11
6 7 3 9 15 13 3
11 7 0 13 3 13 3 1 9 7 13 15
3 0 9 9
2 13 15
6 7 11 9 3 13 15
7 16 0 13 3 13 9 9
15 7 16 13 9 0 13 10 9 16 3 13 13 13 9 0
11 7 9 13 9 1 9 13 1 15 15 9
6 13 3 16 9 0 13
19 16 3 15 3 13 15 0 13 3 3 15 13 15 7 15 13 1 15 9
14 3 9 9 9 1 11 11 0 13 15 9 9 7 9
10 7 16 15 9 11 3 13 0 13 15
22 9 13 3 9 13 13 15 9 15 1 9 0 16 9 15 13 0 7 0 9 9 15
11 7 3 3 13 13 7 13 15 9 7 9
9 3 3 3 13 7 13 7 13 9
4 15 15 13 3
10 16 13 9 9 11 3 9 9 9 13
4 13 1 9 9
5 3 13 1 9 15
20 16 16 13 1 9 15 9 11 7 13 1 9 15 16 9 15 13 1 0 13
5 7 3 13 1 13
3 3 3 13
6 13 13 10 15 3 13
2 3 13
2 13 3
8 7 0 16 13 15 1 9 13
8 1 9 13 3 9 7 9 9
22 3 13 15 0 9 7 13 9 9 15 1 13 15 13 9 9 15 0 7 13 7 13
4 9 15 3 13
4 13 10 13 15
10 16 13 13 1 15 1 15 9 9 13
8 3 13 1 9 7 13 9 9
5 7 16 0 13 13
3 15 9 9
8 13 3 9 9 7 13 9 9
5 15 9 13 7 13
2 13 15
16 13 3 9 9 9 7 9 7 9 7 9 7 9 1 9 0
3 3 13 13
7 7 9 9 13 15 15 9
12 15 13 11 7 15 11 7 15 11 7 15 11
9 13 9 10 0 7 9 10 0 13
4 16 15 0 13
7 15 7 3 13 15 3 13
7 15 7 3 0 7 15 0
5 13 15 1 10 9
14 15 3 3 3 1 9 15 9 16 0 13 13 7 13
30 7 10 9 0 13 3 15 7 9 9 1 9 3 13 7 16 13 13 13 7 1 9 15 3 13 7 9 9 3 13
8 15 3 13 15 9 16 9 13
3 9 13 13
10 7 9 13 3 13 1 9 1 0 13
22 16 3 15 13 15 10 13 9 1 9 9 13 3 9 15 0 13 13 1 9 13 13
6 3 9 15 9 15 13
6 1 9 3 11 13 13
10 0 7 3 13 1 9 16 9 15 13
4 13 15 15 13
7 3 13 3 15 9 9 13
7 9 13 3 9 7 9 15
6 13 15 13 3 15 11
10 7 16 0 13 9 1 13 7 13 13
1 13
16 15 3 13 7 13 3 9 15 0 13 7 13 3 13 9 9
19 16 13 9 16 3 13 9 3 13 10 9 7 1 10 9 13 1 10 9
25 7 16 13 9 7 13 15 9 7 15 9 7 13 15 9 16 9 13 7 9 3 13 3 9 13
2 3 13
4 7 16 9 13
11 13 3 1 9 1 9 7 3 9 1 9
6 10 0 9 15 0 13
10 16 9 15 13 1 12 7 0 12 7
28 7 9 9 13 15 13 7 10 9 15 1 15 0 3 13 7 0 15 15 13 7 3 15 7 9 9 1 15
7 3 3 10 13 1 11 13
13 13 3 15 13 1 16 13 15 9 15 1 9 15
15 16 1 9 1 9 13 1 11 15 15 9 16 0 3 13
1 0
7 3 1 9 9 1 0 9
21 3 3 9 15 0 0 13 13 13 1 9 9 3 13 16 9 15 13 0 1 9
11 3 13 15 15 9 13 1 15 16 9 13
2 13 13
6 13 15 3 1 9 0
11 7 3 13 1 0 9 9 13 13 1 11
54 7 0 1 15 0 9 9 13 16 3 13 13 1 15 0 7 1 9 10 13 0 15 1 0 9 15 13 7 13 1 15 13 16 13 1 13 3 15 1 15 9 16 1 0 9 10 1 15 9 1 0 13 1 15
8 3 0 9 9 1 15 10 6
24 7 1 0 9 7 9 9 13 15 1 0 9 3 16 13 7 16 9 13 15 13 9 1 15
6 7 13 15 13 1 11
14 9 15 15 13 13 1 9 15 13 7 13 1 15 9
22 7 13 9 15 16 1 0 9 10 0 9 1 9 10 0 9 13 13 16 1 11 13
23 3 9 15 13 1 9 9 13 15 3 13 1 9 15 1 9 9 9 9 1 9 11 11
36 13 3 10 0 9 9 1 10 13 13 1 15 7 13 3 15 13 1 15 7 13 13 16 10 13 9 11 7 15 1 11 13 7 13 1 15
14 13 3 3 7 13 16 13 1 10 9 0 13 1 9
12 3 9 11 13 15 13 0 16 12 1 15 13
10 1 11 3 13 3 1 9 13 1 15
15 1 9 9 0 7 0 7 1 9 7 9 1 9 7 9
8 15 7 3 9 9 9 1 9
3 3 15 13
16 7 3 13 15 1 11 3 9 13 9 9 15 7 1 15 13
8 1 15 13 15 0 13 10 9
23 3 1 9 13 7 1 9 0 13 1 0 9 13 15 13 9 15 7 9 9 1 10 0
12 3 3 3 16 0 9 7 15 9 7 1 9
11 7 1 11 15 13 9 15 7 9 1 15
10 15 3 13 9 3 1 9 7 1 9
35 1 9 0 9 13 9 1 9 9 15 1 9 11 7 1 9 9 1 15 7 1 15 7 15 9 1 15 13 15 1 9 9 9 1 15
16 3 10 3 9 13 0 13 7 0 7 9 9 0 7 9 13
7 3 6 13 15 0 15 9
16 7 3 9 13 15 0 13 16 15 13 16 3 9 9 13 15
10 7 13 0 16 0 11 13 15 9 9
12 7 1 15 3 15 13 1 9 13 13 3 15
2 3 15
5 15 13 7 3 13
26 7 16 13 13 3 13 9 16 9 13 7 13 16 15 1 15 15 13 1 15 13 7 13 15 1 15
3 15 15 13
3 7 13 3
30 3 13 16 3 13 3 0 3 13 13 15 7 15 13 15 0 3 3 13 15 16 3 9 9 9 9 9 9 9 9
6 0 13 13 3 1 9
6 0 3 3 13 15 9
5 13 15 10 0 15
29 13 16 3 3 13 1 10 13 15 1 9 11 1 0 9 15 13 0 16 15 13 10 13 15 7 13 13 9 11
9 7 3 15 13 16 3 13 7 13
13 7 16 13 11 1 11 1 9 15 13 16 13 13
15 13 16 0 13 1 11 13 13 3 15 0 3 11 9 9
16 15 15 13 9 3 13 15 1 9 11 11 13 13 1 15 13
11 3 0 3 3 1 11 13 13 11 13 13
12 3 3 15 16 13 0 1 9 10 9 13 13
7 13 15 16 3 13 1 15
17 7 0 13 13 1 0 3 7 3 3 1 16 15 13 0 1 15
5 0 3 13 12 9
8 7 15 9 1 11 9 9 13
11 7 13 15 9 13 16 9 13 15 9 13
11 15 13 1 15 1 9 16 3 9 0 13
13 7 16 15 3 13 7 13 13 16 1 15 3 13
6 16 13 9 9 3 13
3 9 3 13
18 3 3 3 0 15 13 13 9 13 7 13 15 13 16 1 15 9 13
6 1 9 13 13 1 11
50 7 9 0 13 1 9 1 10 0 9 15 13 15 7 13 15 0 9 13 15 11 9 13 13 7 13 7 13 1 0 1 11 11 16 13 1 9 10 13 9 9 9 15 1 9 1 15 1 11 11
16 6 3 3 13 9 7 0 7 13 9 10 0 7 0 9 13
30 7 10 0 1 15 13 0 3 13 7 13 1 9 10 13 1 15 15 7 9 1 11 11 7 9 1 15 9 9 6
13 15 13 0 13 3 15 13 1 15 9 16 13 15
19 15 9 0 1 9 15 3 13 7 15 0 13 1 9 9 16 13 9 13
9 13 3 3 9 7 3 9 1 9
10 3 3 9 13 13 15 9 3 9 15
30 13 3 13 9 15 9 7 13 9 9 7 0 9 1 9 9 9 1 15 13 9 9 15 13 15 9 10 0 0 13
7 15 3 7 1 9 7 9
15 7 16 13 1 9 0 15 9 9 13 7 15 13 3 13
37 0 3 13 1 15 15 3 1 11 11 15 1 9 13 3 9 13 13 15 0 9 7 15 0 13 9 9 13 1 9 9 13 7 9 13 3 9
13 3 3 13 15 16 13 15 3 13 7 15 0 13
26 9 0 1 9 11 9 11 11 1 11 1 9 9 1 9 13 9 1 9 10 15 1 9 13 13 0
10 7 16 15 3 13 3 0 15 9 13
19 13 0 15 13 15 1 9 1 11 7 0 9 15 15 9 13 1 9 9
20 15 7 13 15 7 13 7 13 7 13 1 15 0 13 7 9 9 13 1 15
12 3 7 1 11 7 12 9 7 12 9 15 13
19 7 15 13 9 9 9 15 13 9 9 1 0 16 13 1 15 15 9 13
40 3 15 15 13 13 1 9 7 9 9 15 3 13 13 15 3 13 1 9 9 15 7 3 13 9 1 15 15 9 1 9 7 9 13 7 13 13 1 9 9
8 1 15 13 9 9 1 9 9
18 7 9 9 13 1 9 15 1 15 3 13 13 1 12 9 7 13 13
13 15 9 3 13 9 15 1 9 16 3 13 1 9
8 1 9 13 1 10 3 9 13
12 13 10 1 11 9 7 11 7 10 0 15 9
31 3 3 15 13 9 13 16 13 1 15 9 9 9 13 3 3 9 9 7 3 13 3 9 9 15 3 13 1 15 15 13
8 0 3 13 16 1 0 13 13
10 13 3 15 9 13 15 1 9 11 11
22 0 7 3 15 13 1 9 9 16 15 10 13 10 13 1 9 9 3 13 1 10 13
5 3 13 9 7 9
3 13 10 0
3 9 3 13
7 9 9 15 11 11 1 15
48 1 15 3 13 3 1 15 16 15 0 13 10 9 9 15 7 13 15 9 9 15 7 9 9 1 9 16 13 9 9 15 11 11 1 15 7 15 1 15 1 9 9 15 7 9 15 11 11
12 7 9 13 9 15 1 9 9 7 1 9 11
8 3 13 15 1 15 16 13 15
4 1 11 0 13
20 0 10 9 7 15 9 0 16 11 11 13 1 10 9 0 13 15 0 13 15
20 1 15 13 13 15 9 7 9 9 13 1 11 3 13 9 9 1 9 7 9
3 0 10 9
11 9 13 12 9 9 9 3 13 7 15 9
13 7 10 0 3 13 9 13 7 13 15 0 1 9
8 13 1 15 0 7 1 9 3
6 7 0 13 16 13 13
14 13 3 9 9 13 9 3 13 7 0 10 9 9 15
5 15 3 3 3 13
7 1 9 16 3 13 15 13
3 1 11 0
26 9 13 0 9 15 1 15 13 1 9 7 9 1 11 11 10 0 9 13 1 9 0 15 13 1 15
7 13 9 9 13 3 9 13
6 16 13 3 15 13 15
23 7 0 9 9 13 13 9 0 13 9 0 15 13 15 7 13 1 9 15 15 13 9 9
31 3 1 0 13 15 13 1 9 7 13 13 0 13 9 15 13 1 9 0 3 13 15 7 3 3 3 1 9 9 13 0
20 13 1 9 9 7 9 11 11 15 13 13 0 7 0 1 9 15 7 9 15
3 9 13 9
3 11 1 11
5 3 3 13 15 9
24 13 3 0 0 0 13 3 10 1 9 15 13 13 15 9 15 13 13 15 3 13 13 1 9
8 7 15 15 0 13 15 9 13
7 6 9 15 15 13 1 9
