700 11
5 13 2 16 13 2
11 14 13 2 3 14 13 2 3 15 13 2
6 15 9 14 13 0 2
22 14 13 2 9 9 2 9 7 9 13 2 3 13 15 2 16 0 9 13 1 9 2
5 14 4 15 13 2
7 14 3 3 13 1 15 2
5 7 14 13 3 2
19 1 3 0 9 9 13 9 1 9 2 0 1 0 0 9 7 9 9 2
20 14 13 15 0 9 2 14 13 9 1 9 2 9 14 1 9 0 14 13 2
7 0 9 13 0 7 13 2
13 16 9 13 13 9 9 2 7 0 1 9 13 2
8 14 14 13 13 1 15 9 2
12 3 9 13 1 13 9 1 0 2 9 9 2
12 1 9 13 9 12 8 2 13 9 1 9 2
7 9 0 9 13 1 9 2
7 3 13 1 0 0 9 2
11 1 9 13 13 15 1 0 9 0 9 2
9 13 3 1 9 0 9 1 9 2
6 2 7 3 13 13 2
8 2 9 13 1 9 0 9 2
4 2 9 13 2
8 13 9 2 13 15 1 9 2
10 1 0 9 13 1 15 0 9 9 2
5 9 13 0 9 2
5 13 15 1 13 2
3 9 13 2
6 1 9 9 13 9 2
3 13 15 2
11 3 1 0 3 9 9 13 0 0 9 2
7 1 9 0 13 3 13 2
9 13 15 1 15 9 1 0 9 2
7 9 13 14 1 9 9 2
13 1 9 13 0 9 9 13 15 3 1 9 9 2
5 9 9 13 9 2
13 3 0 9 9 0 9 9 14 13 15 14 9 2
7 9 3 14 13 13 9 2
26 9 9 2 13 3 3 1 9 2 1 0 1 0 0 9 13 1 0 2 8 2 9 1 9 9 2
9 1 9 0 9 13 9 0 9 2
7 9 13 15 0 9 9 2
8 9 4 13 1 9 0 9 2
8 1 9 13 15 13 12 9 2
9 9 13 13 0 9 9 9 9 2
10 13 3 9 13 9 0 0 1 9 2
16 1 0 9 9 0 13 13 0 9 2 0 13 13 15 9 2
19 9 0 0 9 1 9 0 4 9 0 9 9 1 0 8 2 9 9 2
5 13 15 12 9 2
17 16 9 4 13 1 9 0 9 2 13 15 0 9 1 9 9 2
5 9 9 0 13 2
4 9 13 15 2
16 0 9 9 13 2 16 9 9 13 0 2 7 14 13 0 2
10 9 13 0 9 1 9 8 2 9 2
9 1 9 0 8 2 13 15 9 2
10 1 9 1 9 9 13 13 9 9 2
7 13 4 1 15 1 9 2
23 0 9 13 3 13 1 9 9 7 9 2 0 13 1 9 9 13 3 1 9 0 9 2
9 1 9 2 9 15 9 13 0 2
12 9 14 12 9 1 13 9 13 15 1 15 2
38 3 9 9 2 13 9 2 13 1 9 2 13 1 0 9 9 9 1 9 2 13 1 9 2 13 15 3 1 9 7 9 13 9 13 13 1 9 2
12 9 13 0 9 7 13 3 0 2 0 9 2
6 13 15 9 2 9 2
6 1 9 13 15 9 2
6 9 15 1 9 13 2
23 2 13 4 15 13 13 15 1 13 1 9 2 7 13 1 9 2 16 13 9 1 15 2
8 9 9 9 1 9 13 0 2
17 9 9 9 14 13 1 9 2 16 1 9 9 13 0 1 9 2
12 14 9 9 14 13 2 13 15 1 9 0 2
12 14 9 9 13 2 16 9 9 13 15 3 2
9 1 13 9 3 13 9 9 9 2
16 9 14 13 2 0 1 9 13 1 9 13 9 0 1 9 2
10 14 1 9 13 15 2 16 13 9 2
4 13 15 9 2
4 13 1 9 2
13 14 1 0 9 0 9 13 9 0 1 9 9 2
20 13 15 2 16 0 9 13 1 9 0 9 9 9 2 0 3 13 1 9 2
17 13 15 9 9 1 0 9 1 9 0 2 0 13 0 9 0 2
7 9 9 9 13 1 0 2
7 14 13 9 1 13 9 2
4 9 13 9 2
10 2 1 0 0 9 9 13 1 9 2
7 15 9 1 9 14 13 2
17 2 14 9 13 2 14 13 4 13 9 2 13 9 14 2 2 2
11 13 3 1 9 2 16 13 0 13 9 2
4 9 13 15 2
10 9 2 13 1 9 2 4 14 13 2
9 1 0 9 0 9 13 12 8 2
8 9 9 9 13 3 1 9 2
13 3 9 13 9 2 9 2 9 13 1 0 9 2
16 2 13 9 1 9 7 13 2 16 13 3 13 1 9 9 2
2 13 2
7 9 13 9 1 9 9 2
18 9 7 13 2 13 9 7 13 9 2 0 1 0 9 13 1 9 2
8 1 0 9 9 13 0 9 2
10 9 13 1 9 2 16 4 13 9 2
10 1 9 1 9 12 9 13 0 9 2
9 0 9 13 1 0 9 9 9 2
6 7 9 14 15 13 2
12 1 9 9 0 4 13 12 9 8 0 9 2
10 9 3 13 12 9 7 9 0 13 2
20 1 0 12 9 2 1 14 9 9 13 9 1 13 7 9 0 9 0 9 2
15 9 9 13 2 16 1 0 9 9 13 1 0 9 9 2
14 9 13 13 2 14 0 9 13 9 1 9 13 0 2
12 14 3 1 9 1 9 13 9 1 13 9 2
15 9 14 13 13 9 1 9 13 9 1 9 0 1 9 2
9 9 4 13 13 1 15 14 3 2
22 13 13 1 12 0 9 1 0 9 2 7 9 9 13 2 16 9 3 4 15 13 2
10 0 9 13 9 1 9 7 13 9 2
9 13 15 0 9 1 15 13 9 2
11 13 4 13 2 3 13 9 9 1 9 2
8 9 0 9 13 1 0 9 2
8 1 9 13 15 14 9 9 2
7 3 13 15 13 1 9 2
8 9 1 9 9 9 13 0 2
7 9 4 13 1 0 9 2
6 0 9 0 13 0 2
18 14 0 9 13 0 9 1 9 0 9 1 9 13 15 0 9 9 2
8 9 1 9 13 9 12 9 2
5 9 13 1 9 2
16 1 9 9 2 14 13 15 9 2 0 13 1 9 1 9 2
22 9 0 7 9 9 1 9 3 13 1 9 1 9 0 9 2 9 7 9 0 9 2
16 0 9 3 14 13 9 9 2 1 9 13 1 9 9 9 2
12 3 1 9 9 1 9 13 13 1 13 9 2
13 9 13 1 9 1 0 9 2 15 9 13 0 2
11 9 13 9 1 9 1 12 9 1 9 2
4 14 13 15 2
12 3 13 2 16 9 1 9 9 0 13 0 2
8 9 9 13 13 9 9 0 2
13 1 0 9 13 12 9 2 0 13 1 0 9 2
6 14 13 15 9 0 2
12 1 0 9 4 4 1 9 0 1 0 9 2
5 14 13 0 9 2
17 9 1 9 14 13 2 9 13 13 1 0 9 9 1 9 0 2
9 9 13 2 16 9 13 1 9 2
8 1 9 13 4 3 0 9 2
19 13 3 0 1 9 9 2 16 1 13 9 13 1 9 9 13 9 9 2
10 9 13 15 1 9 13 3 1 9 2
10 9 13 9 7 9 13 1 9 9 2
9 1 0 9 0 9 13 3 3 2
10 14 14 4 13 0 9 7 0 9 2
23 13 15 9 2 13 1 9 9 13 3 13 9 7 13 15 3 2 13 13 9 13 9 2
8 7 14 0 3 9 13 9 2
7 13 14 14 0 9 9 2
12 1 9 14 13 9 3 0 1 0 9 9 2
7 14 13 2 9 14 13 2
6 2 13 4 9 2 2
3 9 13 2
16 1 9 9 7 9 0 13 14 0 9 9 1 9 9 0 2
18 14 14 1 0 9 9 0 4 13 7 7 9 2 7 14 9 0 2
11 1 14 12 9 9 9 9 13 0 9 2
17 9 13 1 9 1 9 2 1 0 13 1 9 1 9 1 9 2
12 3 13 12 9 2 7 9 14 13 13 9 2
13 13 1 9 1 13 0 9 9 7 13 1 9 2
6 14 13 15 1 9 2
4 9 4 13 2
8 13 15 13 1 0 9 0 2
22 13 1 13 2 16 1 9 0 13 15 9 1 13 9 0 1 9 9 0 7 0 2
4 13 15 12 2
5 0 13 3 0 2
12 13 4 2 16 13 0 2 16 13 1 9 2
8 1 9 1 3 14 13 9 2
14 9 9 9 13 9 1 9 2 13 9 7 13 9 2
8 3 13 13 9 9 2 2 2
3 9 13 2
7 0 9 9 13 0 9 2
8 13 14 1 9 3 0 9 2
26 16 9 13 15 1 0 9 1 9 1 9 9 2 9 9 13 15 1 9 2 0 13 1 9 0 2
13 0 9 4 13 1 9 2 7 9 13 1 9 2
10 1 0 9 1 9 13 12 8 9 2
5 13 1 15 9 2
7 13 4 13 1 0 9 2
8 9 0 3 13 1 0 9 2
5 9 0 4 13 2
10 9 0 1 9 13 9 9 9 0 2
18 1 0 9 13 15 0 0 9 7 14 9 0 9 13 0 9 9 2
24 1 9 13 2 16 9 1 9 1 0 9 4 13 1 9 7 3 13 0 9 13 3 3 2
6 9 13 1 0 9 2
4 14 13 15 2
4 2 13 15 2
6 16 0 9 13 0 2
7 2 7 15 9 9 13 2
4 2 14 13 2
4 2 0 13 2
8 9 13 1 3 0 0 9 2
7 7 13 15 1 9 3 2
3 2 13 2
5 13 15 9 13 2
5 2 13 2 2 2
3 13 9 2
5 2 13 15 3 2
4 9 14 13 2
3 13 9 2
8 3 13 9 13 15 0 9 2
5 3 13 15 3 2
8 9 13 15 9 1 9 9 2
15 1 12 9 9 13 15 1 13 0 9 1 3 13 9 2
11 13 2 16 13 1 9 12 9 9 0 2
11 14 3 3 13 15 9 14 0 2 0 2
11 4 13 3 0 7 0 9 1 9 9 2
16 1 3 14 13 0 9 2 7 1 9 13 1 0 9 9 2
16 14 14 13 9 2 16 13 15 1 9 1 9 7 15 9 2
13 0 9 1 9 9 13 13 1 9 9 9 9 2
12 9 13 0 9 2 0 4 13 1 0 9 2
8 3 3 9 13 1 9 9 2
7 1 0 9 13 14 9 2
9 9 4 13 1 9 9 9 0 2
6 3 4 13 9 0 2
13 9 8 2 9 9 13 1 9 9 0 1 9 2
8 1 9 13 13 1 9 0 2
6 9 1 9 14 13 2
5 14 13 1 9 2
5 9 13 3 3 2
4 9 13 15 2
22 9 13 1 9 2 13 15 7 13 9 2 9 13 2 16 15 9 13 15 0 9 2
7 13 2 16 3 4 3 2
6 9 14 13 15 9 2
4 13 15 13 2
4 13 15 13 2
4 2 14 13 2
7 9 9 13 7 13 15 2
4 3 14 13 2
3 14 13 2
7 9 13 1 9 1 9 2
9 9 9 14 13 2 9 14 13 2
6 2 13 15 1 9 2
10 13 9 7 13 2 16 0 3 13 2
4 9 13 15 2
10 2 9 13 9 7 13 15 13 9 2
4 2 14 13 2
9 2 9 13 15 13 0 7 0 2
5 2 3 9 13 2
10 1 9 9 0 9 3 13 0 9 2
15 9 9 2 1 9 0 9 1 9 2 3 13 1 15 2
8 9 9 13 9 1 13 9 2
7 9 7 9 13 1 9 2
7 9 13 15 1 0 9 2
6 14 13 3 1 15 2
15 13 1 0 9 1 0 0 9 2 1 0 13 3 15 2
22 14 13 0 9 2 1 0 1 9 14 13 0 9 2 16 9 3 3 13 15 13 2
10 7 14 13 0 1 15 0 9 2 2
20 16 13 1 9 2 9 13 1 9 9 7 13 15 1 9 1 0 9 9 2
11 13 15 15 9 0 2 16 3 13 0 2
11 9 13 14 1 9 7 13 1 15 13 2
10 14 13 2 1 9 13 0 9 9 2
26 15 13 1 0 9 2 0 1 0 9 13 0 9 2 16 13 14 15 13 0 9 1 3 0 9 2
8 9 9 13 9 2 9 13 2
18 9 9 13 1 9 1 0 9 0 7 13 1 0 9 1 0 9 2
11 7 14 2 3 7 3 13 14 0 9 2
16 1 0 9 0 9 0 13 1 0 9 2 7 3 15 13 2
19 0 0 9 13 4 13 1 9 2 7 9 14 13 15 1 9 0 9 2
7 1 9 0 13 15 9 2
10 3 1 9 0 9 9 13 1 9 2
13 9 0 13 1 13 0 9 2 16 0 4 9 2
10 3 1 9 1 9 13 0 9 9 2
4 13 2 9 2
10 13 0 9 9 2 13 4 0 9 2
8 9 13 1 9 9 1 9 2
5 14 13 9 9 2
8 1 9 13 15 1 9 0 2
7 1 9 9 13 0 9 2
6 3 14 13 0 9 2
9 1 13 9 13 15 9 1 9 2
10 1 3 0 9 9 9 13 9 0 2
8 9 1 9 13 14 12 9 2
10 13 2 14 3 13 14 4 9 13 2
11 9 0 2 16 13 2 13 15 1 9 2
5 7 3 9 13 2
9 7 9 1 9 14 13 1 9 2
7 13 15 3 7 13 3 2
4 7 13 9 2
8 3 13 9 7 13 15 9 2
5 7 13 1 9 2
5 7 9 9 13 2
5 9 9 4 13 2
6 13 3 2 9 9 2
18 1 9 1 13 15 9 13 15 9 9 9 1 9 9 0 9 9 2
16 2 13 15 2 16 0 9 1 9 1 0 9 13 15 13 2
15 14 9 14 13 1 9 1 9 2 7 14 1 15 13 2
7 9 13 13 1 9 9 2
5 2 13 9 9 2
9 1 15 13 9 9 9 9 9 2
17 2 1 0 14 9 9 9 13 1 0 9 9 1 9 0 13 2
14 13 14 4 14 2 16 0 9 4 13 1 9 9 2
4 13 1 9 2
8 2 9 9 2 13 9 9 2
17 2 13 14 4 13 2 9 9 2 16 0 9 4 13 9 0 2
15 2 1 9 9 13 9 9 2 0 3 4 13 1 9 2
6 2 13 4 9 0 2
3 13 3 2
6 2 9 4 14 13 2
6 13 1 15 14 13 2
9 2 15 14 3 13 13 1 9 2
8 13 1 15 7 13 15 3 2
11 14 3 13 4 1 9 9 9 2 2 2
8 2 14 13 9 2 2 2 2
6 1 9 13 0 9 2
12 3 15 13 4 2 16 0 9 13 3 0 2
10 3 14 9 9 0 14 13 1 9 2
6 2 7 13 9 9 2
9 7 14 13 1 15 1 0 9 2
7 1 9 9 13 15 9 2
11 2 3 15 13 4 1 0 9 2 9 2
9 14 1 0 9 13 14 4 3 2
5 13 13 0 9 2
7 2 14 13 1 0 9 2
21 1 9 0 2 13 3 1 15 9 7 0 9 13 15 13 2 7 13 0 9 2
12 3 2 1 9 9 2 13 4 14 13 9 2
13 14 13 4 9 1 15 9 2 16 13 13 0 2
21 0 0 9 14 15 13 2 7 15 2 0 9 1 9 2 13 4 15 14 9 2
5 2 7 9 13 2
12 13 4 0 9 2 16 14 13 9 1 9 2
4 3 15 13 2
6 13 1 9 9 9 2
24 16 9 13 15 0 1 0 9 1 9 1 9 7 9 0 2 9 0 13 15 0 0 9 2
5 2 9 14 13 2
6 2 9 0 14 13 2
22 9 0 13 9 9 9 9 2 7 9 13 9 9 0 2 0 1 9 9 9 9 2
14 1 9 1 9 0 9 0 9 13 15 1 9 9 2
11 13 4 1 9 0 9 7 3 13 9 2
7 13 9 14 13 9 0 2
18 0 1 15 15 1 9 13 2 7 9 9 1 0 9 13 15 0 2
9 16 3 13 2 3 14 4 13 2
20 9 1 9 0 13 13 1 0 9 1 9 2 9 7 0 9 13 0 9 2
14 1 9 13 9 1 9 0 1 9 0 9 1 9 2
7 13 8 2 12 9 9 2
12 1 0 9 0 9 13 14 12 8 9 9 2
8 9 13 15 1 9 9 0 2
15 13 14 9 1 13 9 0 1 9 2 9 7 9 0 2
9 13 9 9 13 14 12 9 9 2
12 9 9 0 1 9 13 0 9 1 9 9 2
15 9 13 1 9 13 9 2 7 9 14 13 14 0 9 2
8 3 1 9 9 9 9 13 2
20 9 9 9 13 13 1 9 0 0 9 2 0 9 0 14 1 9 14 13 2
7 9 3 13 9 0 9 2
10 4 13 9 9 7 13 1 0 9 2
9 13 15 9 9 7 9 1 15 2
5 13 15 1 9 2
8 12 9 9 13 1 9 9 2
5 7 9 15 13 2
9 12 9 13 13 0 9 0 9 2
10 0 9 1 9 9 13 1 0 9 2
6 9 15 13 0 9 2
18 9 0 14 13 9 1 9 2 4 13 9 0 7 9 13 1 9 2
13 14 13 15 13 9 1 0 9 1 9 0 9 2
8 14 14 13 15 1 9 3 2
6 1 9 13 12 8 2
11 13 15 0 9 0 7 14 13 0 9 2
10 0 13 14 9 13 13 0 9 9 2
8 12 9 1 14 13 9 0 2
18 9 1 9 9 9 13 13 0 9 9 2 0 13 0 2 0 9 2
13 7 9 2 13 9 2 13 9 7 13 0 9 2
10 1 0 9 0 9 13 13 0 9 2
25 9 9 9 2 13 1 9 9 1 9 2 13 1 9 9 1 9 9 0 2 13 13 15 9 2
12 14 13 14 7 0 9 2 7 0 9 9 2
7 13 7 0 9 7 9 2
7 1 0 9 14 14 13 2
10 9 9 9 3 13 15 1 9 9 2
15 13 15 2 16 1 9 9 9 9 0 13 0 9 0 2
4 9 13 9 2
12 13 1 0 9 9 9 7 13 9 1 9 2
19 9 13 15 2 3 13 15 2 14 1 9 13 15 9 1 9 0 9 2
3 14 13 2
8 14 9 0 9 13 1 9 2
3 13 15 2
8 3 13 2 16 4 13 9 2
10 8 2 9 9 13 15 0 9 13 2
3 13 9 2
14 9 13 15 1 9 2 0 13 0 1 9 9 9 2
5 9 0 14 13 2
8 9 0 13 13 1 9 9 2
9 13 15 14 9 2 13 0 9 2
12 1 9 13 15 13 3 1 9 9 1 9 2
16 3 1 9 1 9 13 15 1 9 9 9 2 1 0 13 2
4 7 9 13 2
9 3 13 9 2 1 0 15 13 2
3 3 13 2
7 9 13 15 3 1 9 2
21 1 9 9 9 13 15 13 0 9 2 16 13 2 9 14 3 15 13 1 9 2
5 14 9 13 13 2
3 9 13 2
14 13 15 0 9 13 4 1 9 7 13 4 1 9 2
12 1 9 2 0 9 14 13 14 9 1 9 2
10 2 9 1 9 13 9 1 9 9 2
21 0 9 0 9 2 13 9 9 0 1 9 0 2 16 15 13 4 1 9 9 2
13 1 3 0 9 9 14 0 9 13 4 1 9 2
13 9 13 2 16 13 15 9 7 13 15 1 9 2
10 13 0 9 1 9 0 14 0 9 2
8 1 0 9 9 3 13 9 2
5 13 4 15 9 2
5 14 15 15 13 2
3 14 13 2
4 9 13 9 2
5 13 4 0 9 2
13 13 15 3 2 16 9 13 15 0 1 0 9 2
10 13 1 15 0 9 2 13 1 9 2
9 13 1 15 1 0 9 0 9 2
6 13 4 3 15 9 2
8 9 0 4 13 1 0 9 2
6 9 0 9 13 0 2
6 9 13 15 1 9 2
6 13 1 13 9 9 2
4 13 9 13 2
4 14 13 9 2
3 13 3 2
8 13 1 13 9 9 9 0 2
15 9 9 1 13 9 13 4 13 1 9 13 9 0 9 2
9 2 9 1 9 13 1 13 9 2
6 9 15 13 1 9 2
4 9 13 0 2
7 13 2 16 9 4 13 2
22 1 9 9 13 2 16 9 13 9 1 9 9 1 9 9 1 13 7 13 9 0 2
15 2 13 9 2 9 9 2 9 13 3 13 9 0 9 2
25 1 0 9 13 2 16 9 9 13 0 7 0 9 2 13 0 9 0 9 7 3 13 15 9 2
10 13 1 13 1 9 1 13 9 0 2
3 3 13 2
9 13 9 0 13 9 1 9 9 2
7 13 13 9 9 1 9 2
6 2 13 4 13 9 2
8 2 13 14 4 13 9 0 2
4 2 13 3 2
6 2 3 13 1 9 2
4 2 3 13 2
6 9 13 15 1 9 2
4 9 13 0 2
6 2 9 0 4 13 2
2 13 2
6 2 13 2 9 9 2
3 2 13 2
12 9 13 0 9 1 9 1 9 9 9 0 2
4 14 13 9 2
10 13 2 16 13 9 13 0 9 9 2
2 13 2
6 13 1 13 9 9 2
18 3 13 13 1 9 13 1 9 2 0 13 9 13 1 9 9 9 2
7 2 0 9 9 0 13 2
9 2 13 2 16 9 0 4 13 2
7 13 1 13 1 9 0 2
4 9 13 0 2
10 9 1 9 9 13 1 13 0 9 2
6 9 13 15 1 9 2
6 13 1 13 9 9 2
3 13 9 2
6 2 13 2 9 9 2
4 14 13 9 2
7 14 13 9 1 9 9 2
3 13 3 2
2 13 2
3 13 9 2
3 14 13 2
10 14 9 1 9 14 13 14 13 9 2
5 13 1 15 9 2
6 9 13 15 1 9 2
6 13 1 13 9 9 2
5 2 9 13 9 2
5 0 9 13 9 2
19 1 0 9 4 13 3 1 15 2 7 3 13 1 13 1 9 9 9 2
6 13 1 13 9 9 2
5 14 13 0 9 2
4 13 1 9 2
13 13 2 16 4 13 9 0 7 3 13 15 13 2
7 2 13 3 2 9 9 2
9 1 9 9 13 9 1 13 9 2
22 13 14 9 1 9 9 9 2 0 1 9 0 9 13 2 16 13 9 1 13 9 2
2 13 2
12 13 3 2 9 1 9 13 1 13 0 9 2
4 13 1 9 2
6 9 13 15 1 9 2
7 3 15 13 1 0 9 2
6 13 9 9 9 0 2
7 9 14 13 9 9 0 2
13 9 15 14 13 2 9 14 4 13 1 13 9 2
3 2 13 2
8 2 13 1 13 12 9 8 2
13 2 14 4 9 13 1 9 9 2 3 1 9 2
11 3 13 9 0 7 9 13 0 0 9 2
13 13 7 9 2 13 12 9 7 14 3 13 3 2
15 7 9 14 13 0 9 2 9 13 1 0 9 9 13 2
15 1 9 9 0 13 3 1 9 2 0 13 1 13 9 2
13 1 0 9 13 15 3 9 0 9 0 2 0 2
15 14 0 9 9 13 9 2 13 9 0 2 0 0 9 2
22 1 9 9 13 1 9 1 9 9 0 2 8 2 9 9 2 13 13 0 9 0 2
11 13 15 9 9 9 1 9 1 9 0 2
4 2 0 13 2
7 9 13 1 9 9 0 2
7 2 14 13 2 3 13 2
27 12 8 2 8 13 9 0 9 2 12 8 2 8 13 4 1 9 2 7 0 12 8 2 8 13 9 2
22 13 2 16 9 9 13 1 0 8 2 0 9 9 0 2 13 1 0 8 2 9 2
5 9 0 13 3 2
9 9 1 9 13 1 9 13 9 2
22 1 9 9 2 3 13 15 0 9 0 2 1 0 9 13 13 1 9 0 12 9 2
7 13 9 9 7 13 13 2
7 13 1 9 9 2 13 2
10 9 1 9 13 3 1 9 2 13 2
5 13 15 13 9 2
18 13 9 2 13 1 9 9 2 13 0 9 9 7 13 15 1 9 2
22 1 9 8 2 13 15 1 9 9 9 13 1 9 0 7 0 2 13 0 9 0 2
5 13 15 1 9 2
5 7 3 13 9 2
7 7 3 4 13 2 2 2
6 0 15 13 9 9 2
3 7 4 2
10 2 16 15 2 9 2 0 9 13 2
7 7 9 3 13 1 9 2
5 7 13 1 9 2
9 1 0 0 9 0 9 13 0 2
4 9 15 13 2
13 13 15 14 2 16 9 13 13 1 9 9 0 2
18 12 0 9 1 9 9 1 9 1 9 0 13 1 0 1 0 9 2
7 14 3 3 13 15 9 2
8 3 13 15 9 14 1 9 2
11 0 9 13 3 9 0 7 9 0 9 2
10 13 15 3 12 9 0 7 9 0 2
22 1 9 0 0 9 13 15 1 0 9 7 3 2 13 9 1 9 2 13 13 9 2
22 9 13 1 9 0 9 3 0 9 9 7 13 2 16 15 9 13 15 13 0 9 2
8 0 9 13 15 1 9 9 2
23 13 9 2 13 1 15 0 9 7 13 1 9 9 9 2 1 9 14 9 13 1 9 2
8 3 3 13 3 1 15 9 2
15 13 15 0 9 1 0 9 1 9 7 13 15 15 3 2
13 9 13 9 7 13 13 2 16 9 13 3 0 2
6 9 13 15 13 9 2
6 7 9 3 15 13 2
6 7 14 3 13 9 2
10 13 1 9 2 13 0 9 7 9 2
10 13 14 12 9 2 3 15 15 13 2
13 14 13 13 2 16 9 1 9 1 15 14 13 2
12 13 15 2 16 15 9 13 9 1 0 9 2
6 13 4 14 1 9 2
7 0 9 13 15 1 9 2
9 9 13 15 3 1 0 1 9 2
12 13 15 15 3 2 16 13 15 1 9 0 2
15 13 9 0 1 13 9 7 9 9 1 13 9 9 0 2
25 12 9 13 0 9 9 0 2 0 7 13 13 2 16 4 15 3 3 15 13 1 9 12 9 2
14 13 15 13 9 7 13 9 1 9 0 9 0 9 2
17 2 13 1 0 2 13 9 2 13 1 9 7 9 2 7 9 2
10 0 1 9 9 13 15 15 1 9 2
5 2 13 1 9 2
9 2 14 13 15 3 1 0 9 2
3 13 9 2
10 9 13 1 9 2 1 9 13 9 2
10 13 4 1 9 7 13 4 15 9 2
11 13 4 1 15 7 1 9 13 4 9 2
4 14 3 13 2
2 13 2
8 9 13 1 0 0 2 2 2
6 13 15 15 2 2 2
5 3 13 1 14 2
2 13 2
2 13 2
4 3 9 13 2
21 13 4 15 14 3 1 9 9 2 13 4 15 1 9 7 3 13 4 1 9 2
5 13 15 7 13 2
5 13 1 0 9 2
4 13 0 9 2
12 9 1 9 0 9 13 13 15 1 0 9 2
5 13 2 9 13 2
6 13 15 1 9 0 2
9 9 13 1 9 7 13 1 9 2
8 1 9 13 0 9 0 9 2
4 9 13 9 2
7 9 13 15 1 0 9 2
6 9 15 13 1 9 2
3 13 9 2
8 9 13 15 3 1 9 9 2
12 1 9 9 1 9 13 15 9 1 0 9 2
7 1 9 13 15 1 9 2
9 9 13 0 9 1 0 9 9 2
10 1 9 1 9 13 9 9 1 9 2
8 4 13 1 9 1 0 9 2
9 9 13 15 1 9 8 2 9 2
7 2 1 9 3 9 13 2
16 3 2 1 9 2 4 3 2 13 13 0 9 7 0 9 2
19 1 13 9 1 9 1 9 2 1 9 9 0 13 0 9 1 9 9 2
15 1 9 0 9 2 9 13 0 9 0 0 9 1 9 2
13 2 13 9 2 16 4 9 3 14 1 0 9 2
15 13 14 4 3 0 2 16 9 9 13 13 1 0 9 2
6 9 13 9 15 3 2
7 2 13 15 3 0 9 2
17 9 13 14 0 2 13 9 9 7 13 2 16 13 9 1 9 2
23 1 9 9 13 3 0 9 2 9 9 7 9 13 1 9 13 15 3 0 7 3 0 2
4 9 3 13 2
19 13 9 9 2 9 7 9 13 15 1 9 2 9 7 9 13 1 9 2
11 14 1 9 0 9 2 1 9 13 9 2
6 2 13 0 14 3 2
6 0 9 3 13 4 2
10 2 14 9 14 13 15 1 9 9 2
5 9 13 1 9 2
4 15 9 13 2
5 2 7 13 9 2
6 9 9 13 12 9 2
14 1 9 13 15 9 7 13 15 1 0 1 0 9 2
8 7 14 12 13 1 0 9 2
18 0 9 13 9 0 9 9 2 0 9 9 9 7 0 9 9 9 2
11 0 9 9 0 9 13 1 9 0 9 2
9 15 9 13 9 9 7 9 9 2
6 13 1 9 12 9 2
11 13 13 3 9 2 1 0 13 9 0 2
7 9 0 13 13 0 9 2
18 7 9 13 15 2 16 13 0 9 2 1 9 9 13 14 9 9 2
19 0 9 13 9 7 9 9 0 4 13 1 9 9 9 1 9 0 9 2
12 12 13 9 2 0 9 0 13 12 9 9 2
3 9 13 2
16 12 9 2 0 3 13 1 9 13 2 13 9 1 9 9 2
14 0 13 9 9 0 1 9 1 9 0 13 15 3 2
12 13 13 9 2 13 7 14 1 13 1 9 2
10 1 13 9 9 9 13 9 13 9 2
10 9 1 12 9 13 9 1 12 9 2
12 1 0 0 9 9 13 3 9 1 9 0 2
14 0 1 9 0 13 12 9 0 2 7 14 12 8 2
10 0 1 0 9 0 13 1 9 9 2
19 9 13 1 9 2 16 9 13 9 2 0 0 4 13 1 9 0 9 2
10 3 1 0 9 13 9 0 1 9 2
11 1 9 13 1 9 8 2 1 9 9 2
9 1 9 0 13 9 14 0 9 2
16 1 15 9 9 13 4 14 9 1 9 2 13 9 1 9 2
10 1 9 13 4 2 1 9 3 13 2
6 9 13 9 1 9 2
4 9 15 13 2
9 2 13 2 9 2 13 0 9 2
4 2 13 15 2
10 9 13 0 2 7 13 9 1 9 2
15 9 9 2 1 9 2 13 2 13 15 9 2 13 9 2
4 9 13 9 2
9 2 14 13 1 0 9 2 9 2
5 3 3 13 4 2
8 2 13 2 9 13 9 9 2
17 9 13 9 0 2 1 0 13 14 9 1 9 2 9 7 9 2
20 3 14 13 1 15 13 2 16 15 9 13 14 1 9 9 2 1 9 9 2
7 9 9 13 0 0 9 2
16 13 9 12 9 0 7 0 9 0 2 3 13 15 12 9 2
30 1 0 8 2 13 9 1 9 9 0 1 9 9 7 9 7 9 0 2 7 14 9 1 9 9 1 9 9 0 2
20 1 0 9 2 3 13 0 9 2 1 15 9 13 3 12 9 9 7 9 2
22 15 9 1 12 9 13 0 2 13 12 9 1 9 0 2 4 13 9 0 7 0 2
7 9 0 13 9 0 9 2
10 9 13 4 3 1 9 9 7 9 2
10 14 12 1 15 13 1 8 2 0 2
14 1 9 13 12 9 2 13 1 9 0 1 0 9 2
17 2 16 14 13 9 1 13 15 1 9 2 7 15 3 14 13 2
15 14 13 13 9 9 7 9 2 16 3 13 1 0 9 2
10 2 0 9 13 15 3 13 1 9 2
9 2 3 13 9 0 9 1 9 2
16 2 1 9 9 9 9 13 2 16 14 13 9 1 9 13 2
16 9 2 0 13 4 1 9 9 1 9 2 13 9 1 9 2
13 1 9 14 13 9 2 7 13 13 1 9 0 2
6 3 15 0 9 13 2
5 13 9 1 9 2
6 1 0 9 15 13 2
15 13 1 9 7 13 15 0 13 2 7 13 15 0 13 2
5 0 9 13 0 2
6 9 9 4 3 13 2
7 9 3 13 1 0 9 2
17 13 9 0 2 0 9 2 13 9 1 9 2 0 15 13 9 2
8 1 0 9 13 15 9 0 2
4 13 2 2 2
7 15 9 13 1 0 9 2
10 9 0 9 4 13 1 0 9 9 2
8 9 13 7 13 15 1 9 2
11 9 9 13 0 2 9 9 0 4 13 2
11 13 0 13 1 0 9 1 9 9 9 2
9 0 9 13 9 0 9 7 9 2
6 0 9 13 1 9 2
21 3 8 2 8 2 0 2 12 2 1 13 9 0 2 1 9 9 9 13 9 2
6 13 4 7 9 0 2
8 3 15 13 7 13 0 9 2
12 13 4 7 2 16 14 13 9 0 1 9 2
10 14 9 13 15 9 1 9 12 9 2
12 3 13 9 8 2 2 0 13 0 1 9 2
7 9 9 1 9 14 13 2
11 1 9 0 2 0 9 13 15 0 9 2
6 1 9 9 13 0 2
5 0 9 3 13 2
5 9 13 1 9 2
7 7 9 13 15 1 9 2
12 16 9 13 9 1 13 9 2 9 14 13 2
10 1 9 9 9 13 9 9 1 9 2
7 9 13 15 1 12 9 2
6 9 13 15 1 9 2
19 1 9 9 1 9 9 13 9 0 1 12 9 2 9 0 7 0 9 2
10 1 0 0 9 4 14 9 9 0 2
8 3 13 15 9 0 1 9 2
17 9 14 13 1 9 2 16 13 4 0 9 1 9 9 1 9 2
7 13 15 1 9 1 9 2
17 1 0 9 0 9 1 9 7 9 13 13 9 1 9 1 9 2
6 13 15 14 1 9 2
6 9 13 0 9 9 2
19 1 0 9 7 13 9 9 9 9 13 15 1 0 9 2 16 13 9 2
18 16 1 13 9 9 13 13 9 2 4 3 13 1 9 7 13 9 2
15 9 9 2 13 1 9 2 13 1 9 0 12 0 9 2
13 13 2 16 13 3 3 13 1 13 0 0 9 2
12 1 0 9 9 13 1 9 9 13 0 9 2
10 15 9 3 13 14 15 14 1 9 2
14 13 2 13 2 13 2 3 13 14 13 9 0 9 2
19 1 9 2 13 0 9 7 9 0 9 2 13 4 1 9 13 3 9 2
9 13 13 9 9 2 7 14 9 2
10 0 9 13 1 9 1 12 9 9 2
18 13 3 13 2 16 9 13 15 9 0 9 2 15 0 9 7 9 2
10 3 1 0 9 13 9 1 9 9 2
4 13 3 0 2
7 7 13 15 3 1 13 2
5 13 12 1 9 2
9 7 14 13 3 0 2 1 9 2
12 7 9 2 1 0 9 2 13 3 3 3 2
5 3 13 4 15 2
