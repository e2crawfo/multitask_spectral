1684 17
14 15 1 11 11 2 11 11 7 11 14 0 9 13 2
26 10 9 1 9 1 11 9 13 2 15 14 11 1 9 13 7 0 13 1 9 14 9 13 4 4 2
14 11 1 9 11 1 11 7 11 1 1 1 0 13 2
26 15 11 1 12 9 1 7 11 1 12 9 1 2 9 2 13 1 12 3 0 9 7 9 9 13 2
7 15 9 14 12 9 13 2
14 15 0 9 7 0 9 1 12 10 14 0 9 13 2
14 15 11 9 13 2 15 10 0 13 7 0 14 13 2
17 9 13 16 10 9 1 11 1 11 1 13 1 1 9 13 4 2
11 9 1 11 7 11 1 9 1 9 13 2
18 0 9 11 1 13 2 15 11 9 1 0 9 13 4 14 0 13 2
11 9 1 9 1 11 9 1 0 9 13 2
13 0 9 1 11 2 11 7 11 1 9 0 13 2
6 15 10 9 14 13 2
12 15 9 11 11 2 11 11 7 11 11 13 2
9 10 9 1 0 9 13 4 4 2
19 9 13 16 15 10 9 13 2 15 9 13 11 1 11 1 9 13 4 2
19 11 1 9 16 11 9 1 9 2 3 9 9 2 14 15 13 4 4 2
6 11 11 13 4 9 2
22 11 9 1 0 9 2 11 2 1 9 11 11 1 9 1 9 0 13 4 4 4 2
8 12 9 1 9 13 4 4 2
16 0 13 1 9 1 11 11 1 0 9 1 9 13 4 4 2
8 9 1 9 11 11 13 4 2
23 9 3 9 0 13 9 1 9 7 9 1 12 9 1 9 1 1 11 1 13 4 4 2
14 9 1 9 9 1 9 1 9 1 9 1 13 4 2
9 3 12 9 0 9 13 4 4 2
19 12 9 1 9 1 9 11 1 9 13 1 9 14 11 9 1 13 4 2
8 15 11 1 9 9 13 4 2
31 11 1 10 9 1 11 11 1 9 9 7 9 1 1 13 4 4 10 9 1 1 11 1 11 9 1 9 13 4 4 2
22 10 9 11 11 1 9 1 9 13 4 2 10 9 11 9 1 9 1 9 13 4 2
16 10 9 9 9 11 1 9 13 7 15 9 9 1 13 4 2
14 11 9 1 9 13 14 11 1 9 0 13 4 4 2
16 11 9 1 0 9 1 0 11 9 11 11 1 13 4 4 2
15 10 0 9 1 11 7 11 1 9 1 9 13 4 4 2
22 11 11 1 0 10 0 9 1 9 13 1 1 15 0 9 1 9 1 9 13 4 2
10 9 11 1 1 1 10 9 0 13 2
37 12 9 1 1 11 11 1 15 15 9 11 1 15 0 13 9 1 15 1 0 13 4 15 9 1 13 9 9 1 1 9 11 1 11 11 13 2
15 10 9 9 11 1 9 1 9 15 2 15 9 1 13 2
21 13 4 16 15 9 1 9 11 1 15 9 11 1 9 13 4 2 15 13 4 2
10 10 9 1 9 1 9 9 13 4 2
9 15 1 9 2 9 13 4 4 2
35 12 0 9 14 0 13 16 11 9 1 9 1 12 9 1 9 1 9 1 9 1 9 13 4 15 0 9 13 7 11 11 1 9 13 2
14 9 15 9 1 13 4 7 9 11 1 9 13 4 2
12 11 0 0 11 9 1 9 10 14 0 13 2
17 10 9 1 9 1 13 4 9 1 9 1 9 15 13 4 4 2
21 9 1 9 11 9 1 9 1 9 13 4 15 11 11 1 9 1 13 4 4 2
9 15 9 1 12 9 13 4 4 2
7 10 9 10 9 13 4 2
19 11 9 1 11 11 2 11 7 11 1 9 9 1 0 9 13 4 4 2
16 10 9 1 9 11 1 9 1 0 9 1 1 13 4 4 2
34 9 1 9 9 12 1 1 9 12 9 1 13 4 4 7 9 9 12 1 1 9 12 9 1 9 9 1 9 2 9 13 4 4 2
14 9 1 9 12 9 1 1 9 1 12 1 13 4 2
13 11 9 1 9 9 7 9 1 1 13 4 4 2
16 9 1 9 9 1 11 9 1 1 9 1 9 13 4 4 2
12 9 1 12 9 0 9 1 9 13 4 4 2
20 9 1 9 1 13 4 4 7 9 1 1 9 1 9 1 9 13 4 4 2
16 9 7 0 9 1 9 1 9 11 1 9 1 13 4 4 2
19 0 9 15 9 1 0 13 15 13 9 2 15 9 9 1 13 4 4 2
15 13 4 4 16 9 1 9 1 11 9 0 9 1 13 2
14 9 1 1 15 1 13 9 1 9 9 13 4 4 2
7 9 15 9 0 13 4 2
14 11 1 11 1 11 11 1 1 11 11 11 0 13 2
10 10 9 11 11 1 12 9 1 13 2
11 11 11 1 9 9 11 1 9 13 4 2
25 11 11 1 9 11 1 9 13 4 2 15 1 9 11 1 15 9 13 16 9 1 9 13 4 2
12 10 0 9 1 9 1 9 3 0 13 4 2
9 9 11 1 9 1 9 0 13 2
9 10 9 12 9 9 1 0 13 2
12 11 11 9 9 11 1 1 14 13 4 4 2
8 11 9 11 1 0 9 13 2
28 0 9 1 9 1 13 4 9 1 9 15 12 9 13 2 1 9 11 9 1 9 11 1 1 0 13 4 2
20 11 9 1 9 9 1 1 0 13 7 15 12 9 0 7 12 9 0 13 2
28 0 9 15 13 16 10 9 1 1 0 11 9 15 14 11 1 11 9 1 9 1 13 4 4 2 13 4 2
7 10 9 1 12 9 13 2
11 10 9 0 2 0 2 9 1 0 13 2
33 0 9 11 11 1 9 11 1 9 1 9 1 0 9 0 13 4 7 15 10 9 1 13 4 9 2 9 1 1 9 13 4 2
13 11 10 9 1 9 13 7 9 1 14 13 4 2
12 15 9 1 9 3 9 1 1 0 13 4 2
14 9 11 1 9 0 9 1 1 1 9 1 0 13 2
10 15 9 1 9 1 9 13 4 4 2
10 11 1 1 0 10 9 12 0 13 2
14 3 1 12 9 1 12 9 0 9 1 13 4 4 2
10 9 1 9 1 0 9 13 4 4 2
16 9 1 0 9 1 11 11 11 2 9 11 1 0 13 4 2
23 9 1 9 10 9 1 13 4 4 10 0 9 1 1 9 13 4 4 7 9 13 4 2
9 10 9 1 1 11 11 0 13 2
18 0 9 1 1 0 9 9 1 9 1 1 9 1 9 13 4 4 2
11 11 9 11 1 9 9 1 3 0 13 2
17 11 1 0 0 9 9 1 9 11 1 9 3 0 13 4 4 2
11 9 1 11 9 1 11 1 9 0 13 2
14 11 9 1 1 12 11 9 11 1 11 9 1 13 2
13 9 9 1 10 9 15 1 9 13 13 4 4 2
4 15 13 15 2
13 11 1 0 9 1 12 9 13 2 11 7 11 2
15 11 9 1 1 1 14 10 0 0 9 1 13 4 4 2
10 10 0 9 1 11 13 4 4 4 2
8 11 1 9 1 9 13 4 2
13 9 2 9 9 2 9 9 7 9 9 13 4 2
29 11 11 11 1 0 9 11 1 9 9 1 13 1 9 13 4 4 7 15 11 1 15 9 1 9 1 14 13 2
14 11 11 9 1 9 1 9 13 13 1 9 13 4 2
42 11 0 0 9 11 11 11 1 13 16 16 11 1 0 11 11 11 1 15 9 1 9 1 13 1 9 13 4 16 11 15 0 9 13 1 1 1 9 13 4 4 2
32 7 11 11 1 15 1 15 9 1 13 13 4 15 1 0 9 1 1 11 1 15 9 1 13 1 0 9 0 14 13 4 2
28 11 11 11 1 11 11 11 1 11 0 0 9 1 11 1 15 9 1 13 1 1 1 9 2 9 13 4 2
66 7 15 15 9 14 13 4 4 16 9 2 9 14 0 9 1 13 4 7 11 1 14 0 9 1 9 13 1 1 1 0 11 11 11 11 1 11 1 13 4 16 11 1 11 11 1 0 9 1 0 9 1 9 15 13 4 15 15 1 15 13 1 0 9 13 2
12 10 9 1 11 1 9 9 14 0 13 4 2
14 9 9 1 9 9 11 11 11 11 1 0 9 13 2
11 11 11 11 11 11 0 9 1 9 13 2
22 11 1 11 11 1 9 9 1 9 13 4 1 3 13 4 1 11 0 0 9 13 2
28 12 0 9 1 11 1 11 1 9 9 13 9 9 1 12 9 9 1 9 13 4 7 12 9 0 13 4 2
35 11 1 0 13 1 12 0 11 9 9 1 9 1 9 13 1 1 0 9 9 11 11 11 11 1 12 0 9 1 11 1 1 0 13 2
27 9 13 4 4 4 16 15 11 1 12 9 13 7 10 3 15 11 11 11 1 12 9 9 13 4 4 2
19 0 9 1 1 2 9 9 1 9 1 9 11 1 0 11 11 11 13 2
26 9 1 13 16 11 11 1 11 11 1 11 1 12 9 1 9 9 1 1 11 1 13 1 9 13 2
34 9 13 16 11 2 11 7 0 0 9 1 11 2 11 9 9 1 9 2 9 1 11 3 1 11 1 1 12 0 9 13 4 4 2
15 11 9 1 11 9 7 11 1 1 10 0 0 9 13 2
29 11 1 11 11 11 1 1 0 11 7 11 11 11 11 7 15 0 0 11 11 11 1 14 0 9 2 9 13 2
13 11 11 2 11 1 1 11 1 11 1 9 13 2
16 11 11 9 1 9 1 13 1 3 15 15 0 11 9 13 2
17 16 2 11 11 9 1 9 9 1 1 14 0 9 13 4 4 2
24 15 0 9 1 1 11 11 1 11 1 9 11 11 1 13 4 1 9 9 1 14 0 13 2
22 11 11 1 0 9 1 13 9 1 12 9 1 13 1 1 9 0 13 4 4 4 2
60 11 11 11 11 1 9 7 11 2 11 1 11 11 11 11 1 11 1 9 1 13 16 11 11 11 11 11 2 11 2 1 9 9 1 1 9 1 13 9 1 0 13 1 9 13 4 4 7 15 1 14 12 12 9 9 13 1 9 13 2
23 11 1 13 16 9 1 0 13 1 9 15 12 9 1 9 1 1 0 13 1 0 13 2
41 15 13 16 9 9 1 12 12 9 1 1 14 9 13 4 1 1 10 9 9 2 9 1 0 13 13 4 4 7 10 9 1 1 9 1 9 3 13 4 4 2
29 11 1 13 16 9 9 1 9 7 9 1 1 0 9 1 14 9 1 13 1 1 1 10 9 9 14 13 4 2
33 11 1 13 16 15 9 13 16 11 7 9 9 1 9 1 14 9 1 9 7 9 2 9 1 9 1 12 12 9 9 13 4 2
35 11 1 12 9 1 0 9 9 11 1 10 9 9 1 0 13 4 4 15 0 9 1 9 1 9 1 9 1 9 1 9 1 9 13 2
18 11 1 9 9 1 0 13 1 10 0 9 1 9 11 11 11 13 2
10 11 11 11 11 1 11 1 9 13 2
42 11 1 13 13 2 15 11 1 10 9 1 9 1 0 13 4 4 15 0 9 1 9 1 9 1 9 1 9 1 0 7 0 9 1 9 13 1 9 13 4 4 2
25 11 1 13 1 9 15 15 13 15 15 12 9 1 11 1 12 9 11 11 1 9 2 9 13 2
47 15 11 1 11 1 9 2 9 1 15 9 13 16 11 11 11 1 9 9 14 15 14 12 9 9 1 9 13 4 4 2 15 15 11 1 9 1 1 12 11 11 1 9 2 9 13 2
16 15 11 1 13 16 11 10 9 9 1 0 0 13 4 4 2
16 11 1 11 1 9 1 10 9 1 0 13 1 9 13 4 2
13 15 11 11 11 1 1 13 10 9 1 9 13 2
15 11 1 13 16 11 11 3 14 11 11 11 13 4 4 2
12 15 1 1 10 9 9 1 9 2 9 13 2
22 0 13 16 11 1 11 1 11 0 11 11 11 1 9 13 1 1 0 13 4 4 2
14 11 7 11 1 15 11 1 10 9 1 10 9 13 2
25 11 1 13 16 10 9 9 1 15 9 1 15 9 1 9 9 11 11 11 1 0 13 4 4 2
11 11 1 15 0 9 13 1 9 13 4 2
19 11 1 11 1 9 13 4 13 4 16 11 1 9 0 9 1 3 13 2
16 11 1 9 1 1 9 9 1 11 1 10 9 0 13 4 2
24 0 3 9 1 11 1 0 10 9 1 0 9 13 7 11 1 9 1 1 9 1 9 13 2
11 15 11 1 1 1 11 11 11 0 13 2
18 7 11 1 2 9 2 1 1 9 15 0 9 1 9 13 4 4 2
23 11 1 11 1 9 1 13 4 13 4 16 0 9 1 11 11 1 13 15 9 14 13 2
20 13 4 4 4 16 9 1 9 1 13 9 7 9 1 1 9 13 4 4 2
16 9 9 1 9 13 7 14 11 1 9 1 9 1 3 13 2
19 12 9 0 9 1 12 2 12 9 13 1 9 1 13 9 13 4 4 2
11 9 1 9 1 1 0 9 0 13 4 2
28 7 15 10 9 1 14 9 9 11 1 11 1 9 1 9 13 16 11 1 9 11 1 9 1 9 14 13 2
26 11 9 11 11 11 1 3 11 11 1 13 16 11 1 9 1 3 14 0 9 1 9 13 4 4 2
20 3 11 11 15 9 1 13 4 7 15 10 9 1 3 14 9 1 9 13 2
18 10 9 11 1 9 11 11 1 13 16 11 11 7 11 1 1 13 2
11 13 4 9 7 9 1 15 15 0 13 2
30 7 9 15 9 1 3 0 0 9 1 13 15 15 13 0 13 16 3 9 1 1 12 11 9 1 9 1 15 13 2
12 3 2 9 11 1 1 11 7 11 0 13 2
17 7 2 10 14 10 12 9 1 11 11 1 13 1 0 13 4 2
24 15 10 11 11 13 2 15 9 11 1 3 13 4 7 15 0 13 1 14 15 9 14 13 2
29 16 0 3 11 11 1 13 1 0 13 11 15 10 9 1 9 1 9 1 0 13 1 1 11 0 13 4 4 2
13 9 1 9 13 11 11 9 1 1 0 14 13 2
5 15 11 1 13 2
7 15 15 9 1 9 13 2
14 11 11 11 1 9 9 9 1 11 11 1 9 13 2
11 7 2 15 11 11 1 9 13 4 4 2
15 3 11 7 11 11 1 9 1 11 11 9 13 4 4 2
17 11 1 9 13 11 1 10 9 1 9 1 11 1 9 9 13 2
23 11 1 11 1 9 1 13 1 9 13 1 9 13 7 2 11 9 3 15 9 13 4 2
27 11 11 1 13 11 1 9 1 9 10 9 1 13 4 4 4 15 15 11 1 15 0 9 1 13 4 2
18 11 1 15 13 2 11 1 1 11 1 13 4 15 9 1 1 13 2
30 11 1 11 1 11 13 4 11 1 11 1 9 11 11 11 1 9 9 13 16 2 9 2 9 7 9 1 13 13 2
26 11 1 11 1 9 9 1 9 13 4 9 13 4 16 15 1 1 11 11 1 9 1 9 13 4 2
14 11 11 1 11 11 1 15 9 9 1 1 9 13 2
9 15 1 11 9 1 9 0 13 2
10 3 11 1 11 11 1 9 13 4 2
13 16 2 10 9 1 12 9 1 11 0 0 13 2
13 9 1 9 1 11 11 1 11 11 1 13 4 2
16 11 15 9 11 1 1 11 11 1 9 1 9 1 0 13 2
18 9 1 1 11 12 9 1 13 1 9 9 1 1 11 1 14 13 2
20 11 1 11 0 0 0 9 1 11 9 13 0 0 9 1 12 9 13 4 2
20 11 11 2 11 1 10 9 0 11 11 2 11 11 1 9 1 9 1 13 2
23 11 0 12 0 9 1 9 1 13 16 10 9 1 12 9 13 4 7 12 0 13 4 2
8 9 1 12 9 14 0 13 2
35 0 9 1 13 16 11 1 11 11 11 1 11 1 9 1 9 9 1 0 9 1 1 9 1 9 13 4 7 15 1 1 9 13 4 2
14 0 9 1 14 11 9 13 10 9 1 9 13 4 2
11 7 9 1 9 1 1 1 15 14 13 2
24 0 9 1 1 1 13 4 16 10 9 1 11 11 11 1 1 1 3 1 9 0 13 4 2
21 11 11 2 11 1 11 11 1 0 0 11 1 9 13 4 11 9 10 9 13 2
20 0 13 16 11 1 11 1 11 11 11 11 1 1 0 9 1 9 13 4 2
17 10 9 1 11 14 13 4 7 15 9 1 12 9 13 4 4 2
12 11 1 9 1 12 12 9 1 9 0 13 2
20 0 9 9 1 11 1 12 0 9 1 11 11 1 1 9 9 0 13 4 2
39 9 9 11 11 11 1 11 1 13 16 0 9 9 1 9 1 11 11 1 0 13 4 1 9 1 1 9 9 1 9 1 12 9 11 0 13 4 4 2
24 15 13 16 0 0 9 11 11 11 1 11 11 1 11 1 9 1 0 13 1 9 13 4 2
20 11 1 11 11 1 9 9 11 11 1 1 11 1 0 13 11 13 4 4 2
14 11 1 11 1 11 1 0 9 0 13 1 9 13 2
32 9 9 1 13 16 11 1 11 7 11 1 1 0 9 9 1 9 0 13 1 3 9 1 9 1 1 9 9 0 13 4 2
15 0 9 1 11 11 1 10 9 1 3 14 9 0 13 2
21 11 11 15 2 11 11 11 2 13 1 9 1 10 9 1 0 13 4 4 4 2
30 9 1 0 9 1 0 13 4 9 1 13 7 9 1 9 9 1 9 13 1 1 9 1 1 14 10 9 13 4 2
15 15 9 15 2 11 11 11 2 1 9 13 4 4 4 2
19 0 0 9 9 1 2 9 9 2 1 9 1 0 0 13 1 9 13 2
24 9 1 9 13 16 10 14 10 0 9 15 1 15 9 0 13 0 13 9 9 1 13 4 2
26 10 0 9 1 15 0 9 1 15 9 1 1 15 9 0 13 1 1 11 11 11 13 1 9 13 2
16 11 11 11 1 1 12 9 9 1 1 9 13 1 9 13 2
23 7 9 9 1 13 15 0 9 2 9 1 10 0 9 13 16 10 9 0 14 13 4 2
22 9 9 14 10 9 1 9 13 1 1 15 1 9 1 10 9 1 9 13 4 4 2
35 16 11 9 1 1 0 11 11 2 11 1 14 9 9 1 9 13 4 1 9 13 2 7 9 1 9 1 10 9 15 1 9 1 13 2
21 10 9 1 14 11 11 11 13 1 1 9 7 0 9 1 9 13 1 9 13 2
19 7 15 0 9 9 1 10 9 1 0 9 1 9 0 13 1 9 13 2
38 15 13 4 1 9 2 9 2 9 2 9 2 9 2 9 2 9 7 9 2 9 2 9 7 9 1 0 9 1 11 11 11 13 4 0 13 4 2
23 10 9 1 1 14 10 9 1 13 11 11 11 1 15 14 12 9 9 0 13 4 4 2
12 15 1 12 9 9 9 1 13 4 4 4 2
10 9 1 13 9 0 9 1 13 4 2
28 11 11 11 1 9 13 1 9 1 9 13 16 9 1 9 1 13 4 9 1 9 1 0 9 0 13 4 2
9 10 9 13 15 9 1 13 4 2
12 9 15 9 1 12 9 9 1 13 4 4 2
33 15 14 12 12 9 9 14 0 13 4 4 7 9 11 1 10 9 1 9 0 13 1 1 10 14 10 12 12 9 10 9 13 2
16 10 9 1 10 9 1 9 9 1 1 0 13 1 9 13 2
27 11 11 11 11 1 11 1 13 16 11 2 11 1 9 1 9 13 1 9 1 9 1 9 13 4 4 2
42 11 1 15 11 11 9 1 11 11 11 2 11 2 1 12 9 1 1 9 1 13 16 11 2 11 1 9 1 9 13 1 9 12 0 9 1 9 1 13 4 4 2
20 16 9 1 9 13 4 7 9 13 4 2 16 3 10 9 1 9 13 4 2
36 11 2 11 1 9 1 0 9 1 1 1 11 11 1 13 16 9 13 1 9 1 11 2 11 1 9 1 9 13 1 9 1 9 13 4 2
15 15 13 16 9 1 0 9 1 9 9 1 9 14 13 2
45 9 1 9 1 9 13 4 11 11 1 13 16 9 9 9 1 9 0 13 1 1 3 11 11 7 11 11 1 0 0 9 7 15 0 9 1 9 1 9 1 9 1 13 4 2
42 11 1 13 16 11 3 10 9 1 9 13 4 4 16 11 1 11 11 11 1 11 0 9 7 9 1 1 15 9 1 9 14 13 4 1 15 9 1 0 13 4 2
13 9 15 0 13 4 1 0 9 1 0 13 4 2
26 15 13 16 9 9 1 9 1 9 1 9 1 9 1 9 9 7 9 9 1 9 1 13 4 13 2
33 11 1 1 9 0 13 1 9 1 1 1 11 11 1 13 16 15 0 13 16 11 1 9 1 15 14 3 9 13 4 4 4 2
29 15 13 16 11 11 1 1 0 9 0 13 13 4 7 15 1 0 9 9 1 1 0 9 1 9 13 4 4 2
23 11 11 1 1 11 1 11 1 13 16 15 11 1 0 9 1 13 4 1 1 1 13 2
32 9 1 1 0 11 11 1 0 11 11 11 1 13 16 11 11 2 11 1 11 1 0 9 1 9 1 15 15 9 14 13 2
41 15 13 16 9 1 1 9 1 9 13 4 4 7 15 9 1 9 13 1 13 4 2 7 9 1 9 1 9 14 13 4 1 1 1 15 1 9 14 13 4 2
26 11 1 9 11 11 1 11 1 9 1 1 13 16 11 11 1 0 9 1 13 4 1 1 1 13 2
27 15 13 16 15 1 1 15 9 14 13 4 4 16 11 7 15 9 0 9 1 13 1 9 1 0 13 2
22 15 13 16 9 1 13 4 0 13 7 9 9 1 15 9 1 9 14 13 13 4 2
15 9 1 3 13 4 9 1 9 1 15 14 0 14 13 2
26 11 1 9 1 11 1 13 4 16 15 0 9 1 3 15 0 0 9 1 0 13 1 9 1 13 2
11 16 10 9 1 9 9 1 9 13 4 2
30 11 1 13 16 11 9 3 2 3 0 9 1 13 1 9 1 13 1 9 13 4 2 7 9 1 15 0 13 4 2
25 11 10 9 1 13 1 1 0 9 1 15 13 13 4 2 7 9 9 1 1 1 15 13 4 2
19 15 1 11 1 11 11 7 11 11 1 15 13 9 1 13 1 9 13 2
37 0 3 11 11 1 9 11 11 11 1 9 1 9 13 4 9 11 11 11 1 13 16 9 1 9 0 13 4 16 10 9 9 1 9 13 4 2
17 11 1 13 16 11 1 14 15 1 1 15 9 0 14 13 4 2
41 15 13 16 10 0 13 16 10 9 1 9 1 13 7 15 9 13 1 13 15 11 11 9 1 1 13 7 13 4 16 10 9 9 1 1 9 1 0 14 13 2
35 16 9 1 1 0 9 1 1 12 1 10 9 0 13 2 7 0 9 1 1 1 9 1 13 9 1 1 15 1 14 0 14 13 4 2
13 15 15 9 13 0 13 16 15 9 1 9 13 2
23 11 7 9 1 11 2 11 7 11 11 1 10 9 1 14 9 1 9 0 13 4 4 2
15 11 1 9 1 1 13 1 1 9 13 12 13 4 4 2
22 9 1 12 9 11 2 11 7 11 1 9 15 14 9 1 0 9 1 13 4 4 2
28 11 2 11 7 11 1 9 1 9 2 9 1 9 13 4 4 3 11 7 11 1 15 15 9 14 13 4 2
19 9 1 9 1 9 10 9 1 13 4 1 1 9 1 0 13 4 4 2
13 11 1 12 12 1 10 9 9 1 0 13 4 2
12 9 1 12 1 1 12 9 9 1 0 13 2
15 0 9 1 13 16 10 9 1 9 1 9 13 4 4 2
26 11 1 9 11 11 1 9 1 13 16 11 1 9 1 12 9 1 11 1 11 11 11 0 13 4 2
17 10 9 1 11 11 1 12 9 1 11 9 1 0 13 4 4 2
21 11 1 13 16 9 1 9 7 15 9 1 13 1 9 1 1 0 13 4 4 2
15 11 1 9 2 9 0 9 1 9 1 9 1 1 13 2
12 9 14 1 9 7 9 9 0 2 0 13 2
17 0 9 1 9 1 1 10 9 1 9 9 1 0 13 4 4 2
26 9 9 1 0 9 1 9 9 1 9 1 9 1 1 10 9 1 9 9 1 9 1 0 13 4 2
14 0 0 9 1 9 1 1 1 9 9 13 4 4 2
12 9 1 1 11 7 11 1 9 14 0 13 2
18 11 1 11 9 1 9 1 12 9 1 12 1 10 9 0 13 4 2
21 11 11 11 1 11 11 11 1 0 9 9 11 11 1 9 1 9 1 13 4 2
36 9 1 9 9 1 13 4 16 15 9 9 1 9 2 9 1 9 9 1 9 1 1 11 11 1 11 9 1 13 9 9 1 9 13 4 2
23 9 1 15 14 13 4 16 15 9 1 10 9 1 9 1 1 15 9 1 9 13 4 2
20 9 1 9 9 1 11 11 11 1 11 9 1 13 9 1 9 14 13 4 2
20 11 1 11 11 1 9 1 15 9 1 9 1 3 14 9 1 9 13 4 2
29 15 9 13 16 15 1 15 0 9 1 13 4 9 9 1 9 1 9 11 11 1 0 9 9 1 1 13 4 2
13 11 1 15 0 9 1 9 9 1 9 13 4 2
34 7 9 9 1 11 1 9 7 0 9 1 9 14 13 1 9 1 0 13 4 7 0 9 1 1 15 9 1 0 13 4 4 4 2
43 9 1 13 15 9 1 11 1 13 4 16 15 15 11 1 0 13 15 10 0 9 1 15 9 9 13 2 7 15 1 14 15 9 14 13 16 15 3 0 13 4 4 2
34 15 15 14 9 13 16 9 9 1 9 2 9 1 9 9 1 9 1 1 11 11 1 11 9 1 13 9 2 9 1 9 14 13 2
14 11 11 11 11 11 1 14 15 9 0 13 4 4 2
36 9 1 13 13 16 9 15 9 1 9 13 1 9 1 1 9 1 1 13 4 4 2 15 11 9 13 1 9 13 9 1 1 13 4 4 2
13 15 13 16 9 1 1 9 1 9 10 0 13 2
19 11 1 13 16 9 1 0 7 0 9 13 1 9 13 3 13 4 4 2
11 9 7 11 12 14 9 1 12 9 13 2
20 10 9 13 16 9 9 1 9 2 9 7 9 1 9 1 9 13 4 4 2
15 15 13 16 10 9 1 9 9 1 1 9 0 13 4 2
22 0 0 9 1 9 15 15 9 13 4 4 2 7 10 9 9 1 9 14 13 4 2
25 9 9 11 11 11 1 11 1 0 9 1 9 13 4 13 16 15 9 3 1 0 13 4 4 2
22 15 13 16 11 1 9 9 1 13 4 9 10 9 13 4 2 7 9 1 13 4 2
46 3 2 11 1 11 11 1 13 4 11 11 11 1 11 9 7 11 11 1 11 11 11 11 1 9 9 11 11 11 1 9 1 10 14 10 12 9 0 13 1 9 1 3 9 13 2
8 10 9 1 15 9 14 13 2
12 15 9 7 9 1 9 1 9 9 14 13 2
20 15 13 16 9 1 9 13 1 1 11 15 14 13 13 4 2 15 13 4 2
45 0 13 16 9 1 9 1 0 9 1 9 13 4 9 9 11 1 11 1 9 1 13 4 16 0 2 9 1 9 1 0 13 1 1 15 14 10 14 10 12 9 0 13 4 2
23 7 10 9 1 9 13 1 11 1 11 11 11 1 11 1 9 1 3 9 13 4 4 2
28 11 1 9 1 10 14 10 12 9 13 1 9 11 1 0 13 1 1 1 13 1 15 10 9 1 13 4 2
15 0 11 1 13 16 0 9 1 10 9 14 13 4 4 2
7 15 15 15 9 14 13 2
26 11 11 11 11 1 11 11 11 11 11 11 11 11 11 11 1 0 9 1 13 10 0 13 4 4 2
14 9 1 1 9 1 1 1 10 9 9 1 9 13 2
26 9 9 9 9 9 11 11 1 13 16 10 9 1 9 7 9 1 1 9 13 4 4 15 13 4 2
11 9 1 13 16 15 9 1 9 13 4 2
15 0 9 1 9 1 1 10 9 1 9 13 0 14 13 2
49 9 1 9 1 9 9 2 9 7 9 1 9 1 13 9 2 9 1 9 2 0 9 2 13 9 1 9 2 9 9 1 9 13 1 0 9 7 9 1 1 9 10 15 1 9 13 14 4 2
31 9 1 13 16 15 9 1 10 3 9 13 1 9 1 1 11 9 1 10 9 1 9 13 9 1 9 1 14 13 4 2
25 9 9 9 9 1 9 1 13 16 11 11 9 7 9 1 9 7 15 1 9 1 13 0 13 2
10 11 11 11 11 1 9 14 15 13 2
23 9 1 13 16 9 1 0 9 1 9 11 11 11 1 9 9 9 7 9 9 1 13 2
14 9 1 13 16 15 15 9 0 0 9 1 1 13 2
24 11 11 1 13 16 10 9 1 0 13 4 1 3 10 9 1 12 9 9 9 0 13 4 2
35 10 9 1 1 11 11 11 11 1 1 10 9 13 7 15 9 1 12 2 12 9 1 1 9 1 1 13 1 9 1 15 0 9 13 2
30 9 1 13 16 10 9 1 9 1 1 9 15 15 9 1 9 2 9 7 9 1 9 9 13 1 1 0 13 4 2
19 11 11 11 1 9 11 11 1 9 1 9 14 15 9 1 9 14 13 2
12 11 9 1 10 9 1 9 11 1 9 13 2
29 9 1 0 9 11 11 1 9 1 9 1 0 9 1 9 0 9 9 1 13 16 15 0 9 1 13 4 4 2
22 9 9 1 14 11 11 7 11 1 9 9 9 1 9 1 1 0 9 2 9 13 2
15 10 12 14 9 1 9 7 9 9 1 1 3 9 13 2
20 9 1 9 1 11 1 0 9 1 1 9 1 11 11 11 1 11 13 4 2
26 11 11 9 1 0 9 1 9 9 1 0 13 4 4 7 0 9 1 9 1 9 13 4 4 4 2
36 11 11 1 9 11 11 1 9 1 9 11 11 7 9 9 1 9 11 11 11 11 1 9 1 13 1 3 9 9 1 9 0 13 4 4 2
43 9 9 1 11 11 1 11 11 1 11 1 9 1 0 13 4 1 12 9 9 9 1 0 13 7 13 16 9 1 0 13 1 3 11 11 1 9 1 9 13 4 4 2
14 11 11 1 1 14 9 1 9 11 11 1 13 4 2
24 7 2 9 9 9 11 11 1 9 1 9 9 1 13 4 1 9 1 9 1 9 13 4 2
9 15 15 9 9 15 1 9 13 2
13 9 11 11 1 12 9 1 9 1 13 4 4 2
21 7 2 9 1 0 9 1 15 9 13 4 13 16 15 0 9 1 13 4 4 2
16 15 9 13 16 9 1 13 4 1 15 1 9 13 4 4 2
18 9 1 9 1 9 13 4 7 15 1 9 1 15 9 1 9 13 2
16 12 9 13 9 1 1 9 1 15 9 1 13 1 9 13 2
25 9 1 1 9 1 9 1 15 9 1 1 1 13 15 15 13 2 15 13 14 4 16 0 13 2
17 15 1 9 1 13 2 9 14 13 4 4 16 15 9 0 13 2
7 7 9 1 15 9 13 2
19 11 11 1 14 11 1 9 1 9 0 13 9 1 13 1 9 13 4 2
38 9 1 1 0 9 11 1 11 1 11 11 1 13 9 1 13 9 1 9 13 7 13 16 9 1 9 1 1 9 1 12 9 1 9 1 13 4 2
29 15 13 16 15 15 10 9 1 9 1 13 4 9 7 11 1 13 4 15 1 1 1 9 2 9 13 13 4 2
21 15 9 13 16 9 9 1 9 1 0 14 13 4 7 15 0 9 0 13 4 2
29 15 9 13 4 9 9 1 9 11 11 11 1 13 16 0 9 1 13 4 1 3 9 15 9 1 14 13 4 2
31 11 1 0 9 7 11 1 0 11 11 11 11 1 11 1 13 16 15 9 9 11 11 11 1 15 13 15 15 13 4 2
30 11 1 11 11 1 9 9 13 4 1 0 13 4 11 1 13 16 15 15 1 11 1 1 1 15 9 14 13 4 2
9 15 15 9 1 9 1 9 13 2
29 0 13 16 11 1 9 9 2 9 2 9 2 0 9 9 7 0 9 1 10 9 1 0 13 1 9 13 4 2
28 9 1 13 13 16 11 1 9 1 9 13 4 9 1 10 0 9 1 1 10 9 9 9 1 12 9 13 2
17 9 11 1 0 9 1 9 1 3 10 9 1 1 13 4 4 2
17 7 10 9 1 9 1 12 12 9 1 15 9 13 1 9 13 2
32 11 11 11 11 1 9 11 11 1 13 16 9 1 0 9 11 1 11 1 9 1 14 11 0 15 9 1 0 13 4 4 2
19 10 9 15 15 9 2 9 1 11 1 9 1 12 9 9 13 4 13 2
20 15 13 16 10 9 1 9 13 4 9 1 9 11 1 9 1 12 13 4 2
18 10 9 1 9 1 9 1 12 11 2 11 11 11 2 9 13 4 2
13 15 1 14 10 9 1 10 14 10 12 9 13 2
13 10 9 1 9 1 14 9 1 12 11 9 13 2
54 0 9 1 0 9 1 9 12 9 14 9 13 1 3 11 11 11 2 11 2 1 10 9 12 12 9 9 1 9 1 13 4 9 1 9 12 9 14 9 7 9 1 9 12 9 14 9 13 4 1 9 13 4 2
39 11 9 11 11 1 15 9 1 13 16 16 0 9 1 9 0 9 1 0 13 4 2 16 9 11 2 11 1 1 15 9 9 14 12 12 12 9 13 2
39 9 15 9 1 9 2 9 13 4 11 1 13 16 9 9 9 1 1 15 3 0 9 13 4 4 7 3 14 9 1 13 1 1 10 13 1 9 13 2
29 12 9 1 9 1 15 13 16 9 9 1 0 9 1 13 1 1 0 9 1 14 1 9 10 9 13 4 4 2
18 15 1 14 11 11 1 9 1 14 10 9 1 0 13 4 4 4 2
31 0 13 16 0 9 9 1 9 7 9 1 9 1 9 1 1 14 9 9 1 1 12 12 9 1 9 14 0 13 4 2
16 15 1 1 9 9 15 9 1 10 9 1 9 13 4 4 2
38 15 13 16 16 0 9 1 0 9 1 9 0 9 1 14 13 4 16 0 9 9 1 1 9 9 1 9 1 9 1 12 12 9 1 9 13 4 2
19 0 11 9 1 10 9 1 9 1 12 12 9 1 9 13 4 4 4 2
38 0 13 16 9 9 1 9 1 9 1 9 1 9 2 9 13 1 1 11 11 11 11 11 11 11 0 9 11 11 11 11 1 1 9 13 4 4 2
15 15 1 14 11 11 1 9 1 14 9 9 13 4 4 2
28 10 9 1 9 1 9 1 9 13 1 9 1 1 11 11 11 11 1 0 9 1 0 9 1 9 13 4 2
31 11 2 11 1 0 9 7 11 7 0 0 9 1 9 1 9 1 9 13 1 1 9 1 9 9 1 9 13 4 4 2
17 15 1 9 0 9 1 13 9 9 1 14 3 9 13 4 4 2
21 0 9 1 1 9 1 0 9 1 13 9 1 15 10 9 1 9 13 4 4 2
15 0 9 1 1 9 1 15 1 9 13 4 1 9 13 2
39 9 1 1 0 9 1 9 11 11 11 1 12 9 1 13 9 1 0 9 1 10 9 1 9 13 15 0 9 1 9 1 9 13 1 9 13 4 4 2
14 12 9 1 10 9 1 11 11 11 1 0 13 4 2
36 9 1 1 9 13 4 16 9 1 12 9 11 2 11 2 11 2 11 2 11 7 11 7 0 0 11 1 9 1 9 9 1 13 4 4 2
18 10 9 1 9 9 1 13 4 4 7 15 9 1 9 13 4 4 2
19 0 3 11 1 9 1 9 10 13 1 1 15 13 1 9 14 0 13 2
14 15 14 10 9 13 4 4 15 9 1 13 4 4 2
44 0 9 1 9 1 9 1 1 13 1 12 9 1 13 13 16 15 14 15 9 1 9 13 14 4 4 7 9 1 10 9 1 12 9 3 15 15 9 1 9 13 4 4 2
19 11 1 12 9 9 9 13 4 4 7 15 12 9 14 9 13 4 4 2
27 11 11 1 9 9 1 9 1 13 0 11 1 9 9 11 11 1 9 13 1 9 1 0 9 13 4 2
23 11 1 1 11 1 11 11 13 4 4 7 11 1 15 9 1 0 9 1 11 13 4 2
10 12 0 11 1 9 0 13 4 4 2
31 15 1 11 1 0 9 13 4 2 15 10 9 11 2 11 1 12 9 1 13 1 9 1 9 1 9 1 9 13 4 2
22 11 9 9 9 9 1 0 9 1 11 1 9 1 13 9 1 9 2 9 13 4 2
16 11 11 9 11 1 9 1 0 9 1 0 13 13 4 4 2
12 7 9 1 15 9 1 3 15 9 13 4 2
23 15 3 9 9 1 9 13 4 2 15 9 1 9 13 4 1 1 15 11 11 13 4 2
32 9 11 11 1 13 16 11 1 9 1 0 9 1 9 1 12 0 9 13 4 7 15 9 1 0 9 1 11 13 4 4 2
31 11 1 0 9 1 11 10 9 1 9 1 13 4 4 2 15 9 1 13 1 9 1 9 1 9 1 0 9 13 4 2
18 11 9 9 1 9 9 1 0 9 1 10 9 1 14 9 13 4 2
23 0 9 11 11 7 11 11 11 1 10 9 15 0 0 9 1 0 13 9 1 0 13 2
12 16 15 9 13 4 16 11 3 0 13 4 2
24 9 9 11 11 7 11 11 14 11 1 9 2 9 13 7 9 1 9 13 15 13 4 4 2
42 11 11 11 11 2 11 2 1 11 11 11 11 2 11 2 1 9 9 11 11 1 11 1 9 1 0 13 4 7 0 12 9 1 15 9 13 1 0 9 13 4 2
43 15 1 11 11 11 11 11 11 11 11 11 1 9 1 13 12 9 7 0 9 1 9 1 11 2 11 11 11 2 9 1 9 13 1 0 9 1 9 13 1 9 13 2
10 11 11 10 9 1 9 1 9 13 2
28 11 11 11 1 9 1 12 0 9 1 11 1 0 9 1 9 1 0 13 4 12 0 9 1 0 13 4 2
18 9 1 9 1 11 1 1 11 11 11 7 11 11 11 1 9 13 2
51 9 1 9 11 11 11 1 13 16 9 1 1 9 11 11 1 12 12 12 12 12 12 9 1 9 0 13 4 1 1 1 11 9 1 9 0 13 1 1 1 12 9 1 9 1 9 1 9 13 4 2
18 15 1 14 15 11 1 9 7 9 1 9 1 14 13 4 4 4 2
39 0 13 16 9 1 11 11 11 11 11 11 11 11 11 1 9 11 2 11 2 11 2 11 7 11 2 11 1 11 9 1 13 9 1 9 13 4 4 2
14 9 1 9 11 2 11 1 9 1 15 9 14 13 2
15 0 12 9 1 11 1 0 9 1 9 11 11 0 13 2
28 15 9 1 11 2 11 1 11 9 1 9 13 1 1 9 12 12 9 1 13 12 12 9 13 4 4 4 2
36 10 9 11 11 11 1 11 1 0 9 7 9 1 0 11 2 11 11 9 11 11 11 7 12 9 1 12 12 9 1 9 1 9 13 4 2
35 0 9 11 2 11 1 12 0 0 9 1 9 1 11 9 1 1 9 13 4 7 3 1 15 0 9 1 9 1 9 1 9 13 4 2
50 9 1 9 11 1 13 16 9 1 9 1 1 10 9 3 13 16 11 11 11 11 11 11 11 1 0 11 9 1 9 1 1 10 9 14 11 11 11 7 11 1 13 9 1 9 1 14 13 4 2
27 15 13 16 9 1 10 9 1 9 14 13 1 15 15 1 9 13 4 2 15 3 0 7 0 0 13 2
25 9 1 0 9 1 1 9 13 1 12 12 9 1 12 12 1 9 15 14 9 1 13 4 4 2
14 15 9 14 13 4 4 7 9 9 1 14 9 13 2
14 16 10 0 9 15 9 2 9 1 9 14 13 4 2
26 15 1 14 10 9 1 1 11 11 11 11 15 1 10 9 1 15 0 9 9 14 0 13 4 4 2
22 9 7 9 1 15 9 7 9 9 1 13 1 9 1 14 9 14 13 4 4 4 2
17 11 11 11 1 9 1 1 12 12 9 0 9 9 1 0 13 2
13 15 9 1 9 13 1 1 9 14 1 9 13 2
16 9 11 11 15 3 0 9 0 9 1 0 13 4 13 4 2
15 0 9 1 9 1 1 14 9 1 9 9 13 13 4 2
26 11 11 1 9 9 11 11 11 1 9 1 13 15 9 1 0 0 9 1 0 9 9 13 4 4 2
15 10 9 1 12 12 9 9 7 9 1 9 13 4 4 2
11 9 13 4 1 10 0 9 15 1 13 2
14 7 15 0 9 1 9 1 9 14 0 13 4 4 2
30 0 9 1 9 1 9 13 7 11 11 11 1 0 9 9 11 11 1 1 15 10 14 9 13 0 13 4 4 4 2
6 7 9 13 14 15 2
29 15 1 1 11 11 11 11 1 9 9 1 1 15 9 1 10 9 1 9 1 13 15 9 9 0 14 13 4 2
12 9 9 1 1 9 1 9 9 13 14 13 2
31 11 11 1 9 9 1 9 9 1 9 1 13 11 1 12 9 1 9 13 1 3 15 0 9 0 13 1 9 13 4 2
21 7 0 9 7 9 9 9 1 15 9 0 9 1 1 0 13 1 9 13 4 2
47 11 11 11 11 1 1 9 1 1 11 11 11 2 11 2 7 11 11 11 11 11 2 11 2 1 9 1 13 16 15 9 13 4 1 9 1 9 1 1 11 1 15 9 0 13 4 2
21 15 13 16 9 13 4 1 9 1 0 7 0 9 1 1 1 9 13 4 4 2
19 16 15 9 13 16 9 0 9 11 9 1 1 15 1 1 9 13 4 2
30 11 9 1 9 9 9 11 11 1 0 11 11 1 10 9 1 1 11 9 1 11 1 9 1 13 1 9 13 4 2
33 11 1 9 1 9 1 9 2 11 2 11 2 1 9 1 1 12 9 1 1 11 1 11 1 1 13 1 9 1 9 13 4 2
31 0 9 11 11 11 1 13 16 11 9 1 1 13 4 4 2 7 10 3 16 15 9 13 4 4 16 15 0 13 4 2
25 10 3 9 1 9 1 13 4 0 9 1 9 1 0 13 1 1 11 11 1 1 9 13 4 2
17 11 11 1 1 9 1 9 15 11 1 9 1 14 13 4 4 2
26 11 1 0 11 11 11 1 0 9 1 12 9 1 1 0 9 1 9 13 1 9 9 1 13 4 2
16 0 9 1 0 9 1 1 0 9 1 9 13 1 9 13 2
22 15 9 13 1 15 0 13 16 15 0 2 0 13 4 7 15 9 1 0 13 4 2
16 15 9 9 10 9 1 9 2 9 13 1 9 13 4 4 2
26 13 4 4 16 11 11 1 9 9 1 0 9 1 9 11 11 11 2 11 0 11 11 11 13 4 2
7 11 11 1 11 13 4 2
17 0 14 9 9 9 1 10 9 1 10 0 9 1 15 13 4 2
10 15 11 1 1 0 9 9 13 4 2
11 11 1 15 9 13 15 15 15 3 13 2
17 11 1 9 1 1 15 9 2 9 7 9 1 0 9 13 4 2
9 15 1 15 9 7 9 13 4 2
40 11 1 9 11 11 1 1 11 14 12 9 1 9 1 0 2 0 13 4 2 7 9 9 1 15 9 9 13 1 1 9 1 9 2 9 13 1 9 13 2
13 3 1 11 1 9 11 11 1 10 9 13 4 2
9 11 1 13 11 11 9 9 13 2
14 15 9 1 11 1 9 13 15 9 1 0 13 4 2
8 11 11 11 1 9 1 13 2
17 3 1 15 1 15 8 13 11 1 12 0 9 1 0 13 4 2
15 11 11 1 1 15 14 11 0 11 1 0 14 13 4 2
24 11 1 9 1 9 13 16 9 9 1 9 13 1 9 1 1 15 1 15 9 14 13 4 2
21 15 1 9 9 10 9 1 9 2 9 13 0 9 1 13 1 9 13 4 4 2
25 11 1 9 1 0 9 11 11 2 11 11 7 11 11 1 12 9 1 9 13 1 9 13 4 2
25 10 3 9 11 1 9 9 11 11 11 1 9 13 16 11 11 1 9 9 1 12 9 13 4 2
12 16 15 15 9 1 9 13 1 9 13 4 2
11 15 13 16 10 9 1 9 15 13 4 2
13 10 9 1 9 1 0 9 1 13 4 4 4 2
10 9 1 9 1 9 1 14 9 13 2
34 11 11 11 2 11 2 9 9 1 10 13 12 9 13 1 11 9 1 9 1 9 1 11 1 9 14 1 12 9 9 1 13 4 2
24 0 12 9 1 11 9 9 1 0 13 1 9 13 4 9 1 9 2 9 9 2 9 13 2
20 11 11 11 1 9 1 9 1 9 1 0 9 1 1 9 9 7 9 13 2
12 15 1 15 9 14 13 7 9 14 0 13 2
31 11 2 11 7 11 1 9 9 1 9 1 13 16 9 1 11 1 9 13 15 11 9 9 1 0 13 1 9 13 4 2
30 11 9 11 11 11 1 13 16 9 1 15 9 1 9 1 9 14 1 0 9 7 9 9 9 9 1 9 13 4 2
39 11 1 1 2 9 1 13 4 16 10 9 1 0 13 1 1 9 9 1 9 0 13 4 16 15 12 12 11 9 7 15 12 12 9 0 13 4 4 2
15 15 15 14 13 16 9 1 9 9 1 10 9 0 13 2
32 11 1 3 13 16 9 1 0 9 7 9 2 3 1 9 3 11 2 11 2 11 2 11 7 11 1 14 9 2 9 13 2
30 11 1 9 11 11 11 1 13 16 11 2 11 2 11 11 2 11 2 11 7 11 1 14 9 13 7 9 13 4 2
19 16 2 3 1 9 0 13 1 1 10 9 9 1 3 14 12 9 13 2
23 11 1 9 13 4 11 1 12 0 9 1 1 10 0 9 1 9 15 0 9 0 13 2
13 3 0 9 13 2 10 0 9 1 0 9 9 2
20 3 9 9 1 10 0 0 9 1 10 9 1 9 10 9 1 13 4 4 2
39 15 1 11 1 13 0 9 2 11 1 0 9 7 11 11 1 9 13 4 9 1 9 14 9 14 13 2 15 9 1 1 9 1 13 4 1 9 13 2
20 3 9 1 10 9 1 9 11 1 0 0 9 1 1 10 0 3 13 4 2
28 0 9 1 11 11 11 1 9 1 1 11 1 9 1 13 1 13 4 7 3 9 9 1 14 13 4 4 2
13 12 9 1 11 11 1 11 1 11 9 13 4 2
24 15 11 1 11 11 9 1 13 7 9 1 11 1 11 9 1 9 1 9 13 9 13 4 2
10 11 10 9 9 1 9 1 9 13 2
18 15 11 15 13 1 9 1 14 13 2 7 10 9 9 13 4 4 2
8 15 0 11 9 1 9 13 2
15 11 1 9 1 9 1 1 9 1 9 9 13 4 4 2
18 15 14 13 4 4 4 16 11 11 1 9 1 13 1 0 13 4 2
21 15 1 11 9 7 11 1 0 9 1 9 14 9 1 1 2 9 13 4 4 2
41 16 2 9 1 11 9 11 11 2 11 11 11 2 9 1 0 9 7 11 0 12 9 1 9 1 1 9 7 9 9 1 9 1 14 12 9 9 13 4 4 2
45 13 1 9 9 1 9 9 1 9 0 13 4 13 4 4 16 9 9 0 2 0 7 0 9 1 1 9 2 9 7 9 1 0 9 1 12 0 9 1 1 3 13 13 4 2
21 9 9 1 13 13 16 0 9 1 10 0 9 1 9 9 14 15 0 9 13 2
18 11 11 11 11 1 9 1 0 13 2 7 11 11 11 9 9 13 2
19 10 0 13 2 11 11 1 10 9 1 11 9 2 9 1 9 13 4 2
23 15 14 13 4 4 4 16 3 11 10 9 1 0 14 13 2 16 11 1 9 13 4 2
19 16 9 9 11 11 1 13 13 16 15 11 1 11 1 0 9 13 4 2
6 15 9 13 4 4 2
37 11 1 0 9 11 1 0 9 2 9 1 9 2 9 7 9 9 1 9 13 15 0 2 0 2 9 9 7 9 1 9 1 0 9 13 4 2
32 11 1 11 11 11 2 11 2 7 0 9 1 1 9 9 13 4 9 1 9 7 11 9 11 11 9 1 0 9 1 13 2
40 15 11 1 11 9 1 9 11 11 1 11 11 1 1 9 11 13 4 16 11 11 11 2 11 2 1 9 11 11 1 11 1 0 9 11 11 1 9 13 2
27 11 1 11 1 11 1 13 16 11 11 1 9 1 9 11 2 11 2 7 11 2 11 1 1 9 13 2
6 15 9 11 1 13 2
14 15 13 16 15 11 11 1 11 1 9 1 13 4 2
11 15 15 9 11 1 9 13 4 4 4 2
16 11 1 1 1 11 1 13 16 15 11 1 9 1 1 13 2
63 15 0 9 14 13 4 16 11 11 11 11 1 11 1 11 11 1 0 11 11 11 11 1 9 1 9 9 9 1 0 13 1 9 1 9 1 0 13 4 2 7 9 12 9 1 12 9 3 11 14 9 1 10 9 9 1 9 1 13 9 13 13 2
9 15 9 1 1 0 13 4 4 2
34 9 1 9 1 9 13 4 11 1 13 16 15 9 9 1 10 9 9 1 0 13 1 9 0 13 4 2 15 15 1 13 4 4 2
21 15 0 11 11 11 1 9 13 16 15 13 16 9 1 9 1 0 9 13 4 2
19 3 15 9 9 1 0 13 1 9 0 13 4 7 15 0 13 4 4 2
40 7 15 15 1 11 11 9 1 9 1 9 9 1 9 1 9 0 13 15 1 13 4 15 3 9 1 9 13 4 9 1 9 1 1 10 9 13 4 4 2
18 11 1 13 16 9 9 1 1 0 9 1 9 1 13 1 9 13 2
10 11 1 14 10 9 9 1 13 4 2
15 11 1 11 9 1 14 9 1 9 9 1 9 13 4 2
15 15 9 1 10 9 1 0 9 1 9 1 13 4 4 2
20 15 1 9 1 1 11 11 11 11 11 11 1 11 11 1 9 1 9 13 2
9 15 9 1 9 1 9 13 4 2
13 15 1 9 9 1 9 1 0 13 1 9 13 2
25 11 1 15 13 15 9 13 16 15 1 11 9 15 13 4 9 7 0 9 1 9 13 13 4 2
14 15 0 9 1 3 13 10 9 1 0 13 4 4 2
20 11 11 11 11 11 11 0 13 1 3 9 9 1 9 13 1 13 4 4 2
28 11 11 11 11 1 10 9 1 9 1 9 2 9 1 1 11 11 1 9 1 0 9 9 1 9 13 4 2
22 11 7 9 1 9 1 0 13 16 10 9 1 0 13 1 15 10 9 13 4 4 2
29 11 11 11 11 9 11 11 11 1 13 13 16 10 9 1 0 13 1 1 15 10 14 10 12 9 1 9 13 2
23 10 3 10 9 1 13 9 1 1 9 2 9 13 4 7 15 9 2 9 0 13 4 2
22 9 11 1 9 1 0 13 16 15 10 9 1 11 11 1 0 13 4 0 14 13 2
17 16 11 11 1 11 11 1 9 1 15 0 13 4 1 9 13 2
20 11 1 10 9 1 14 13 15 0 13 1 9 2 9 1 13 9 13 4 2
9 10 9 1 14 9 13 4 4 2
14 10 9 1 9 9 1 9 1 14 0 13 4 4 2
24 9 1 0 9 1 11 1 9 13 4 1 3 9 15 15 9 2 9 0 13 1 13 4 2
26 11 1 9 13 16 9 0 13 1 3 10 9 1 1 9 13 1 9 1 9 9 1 0 13 4 2
17 9 15 1 10 9 1 9 1 0 9 9 1 9 13 4 4 2
23 15 1 9 10 9 1 9 2 9 1 13 11 11 1 1 14 9 2 9 13 4 4 2
33 11 11 1 0 9 11 11 1 9 9 7 15 9 1 13 9 1 9 1 11 1 0 9 1 9 1 11 1 9 1 9 13 2
19 11 11 11 11 1 9 1 13 10 9 9 1 11 2 11 1 9 13 2
12 9 1 0 9 1 9 14 9 13 13 4 2
10 10 9 1 11 1 9 14 13 4 2
19 9 1 0 13 1 1 11 1 1 11 11 1 0 9 1 9 13 4 2
16 9 3 14 11 11 9 13 16 0 9 0 9 1 13 4 2
15 7 0 9 9 1 1 15 0 9 1 9 14 13 4 2
23 9 1 9 13 4 11 1 0 9 11 11 11 1 13 16 15 9 1 9 9 1 13 2
11 11 11 1 9 0 9 9 1 9 13 2
19 9 11 11 1 13 16 11 11 11 11 7 11 1 9 1 13 4 4 2
19 0 9 11 11 1 13 16 11 11 1 9 9 13 15 9 1 9 13 2
24 9 1 0 9 11 11 11 1 13 16 11 11 1 9 1 0 11 9 1 9 0 9 13 2
31 11 1 11 9 11 11 1 13 16 10 9 11 1 9 1 13 4 2 15 15 14 13 4 4 7 11 11 15 14 13 2
15 11 9 11 11 11 1 0 9 1 1 9 1 0 13 2
16 15 13 13 16 11 9 1 15 9 1 10 9 1 13 4 2
33 9 1 11 1 0 9 7 9 9 1 9 11 11 2 9 11 11 11 2 11 11 11 2 9 11 11 7 11 11 14 0 13 2
12 9 1 9 9 1 0 9 11 11 1 13 2
32 0 11 9 1 3 1 9 13 4 11 11 11 2 11 2 1 11 1 9 9 1 0 9 1 0 13 4 1 9 13 4 2
23 11 7 9 9 1 9 9 1 0 9 11 1 9 1 0 9 1 14 12 9 1 13 2
27 9 9 0 9 1 1 9 1 1 11 1 1 9 2 11 9 1 1 9 9 7 9 9 1 9 13 2
34 11 1 12 9 1 1 11 9 1 1 9 13 4 11 9 11 11 1 11 1 13 16 9 9 1 13 13 16 9 9 0 13 4 2
28 16 11 11 1 1 9 13 13 4 16 15 14 15 0 9 1 9 9 1 9 1 13 9 1 9 13 4 2
33 14 9 2 9 11 1 11 1 11 1 9 9 1 10 9 1 9 1 13 1 11 1 9 1 1 1 15 9 0 13 1 13 2
19 9 1 0 9 1 14 13 16 11 1 0 9 9 1 1 0 13 4 2
30 15 13 13 16 9 9 1 11 1 0 2 0 13 1 1 11 1 11 1 9 1 9 1 12 9 0 13 4 4 2
25 11 1 13 16 10 9 1 11 1 15 9 0 13 4 7 9 9 1 9 9 1 0 13 4 2
19 15 13 16 12 9 9 9 13 1 11 1 11 1 0 9 0 13 4 2
31 11 1 3 3 9 13 1 0 13 4 4 16 11 1 11 1 11 1 1 9 9 1 9 9 1 9 0 14 13 1 2
16 10 9 1 9 1 9 9 1 1 14 10 0 9 13 4 2
16 9 9 9 1 10 9 13 1 13 4 9 1 14 9 13 2
27 9 9 1 13 13 16 11 11 11 7 11 11 2 11 11 2 11 9 1 10 9 1 3 13 4 4 2
11 7 0 9 9 9 14 13 1 9 13 2
25 3 9 9 1 11 11 11 2 11 11 2 11 11 2 11 11 2 11 11 7 11 11 0 13 2
23 11 11 11 2 11 2 7 11 11 2 11 2 9 1 1 0 9 1 0 13 4 4 2
10 15 1 0 9 0 13 4 4 4 2
29 15 11 1 11 2 11 2 11 7 11 9 1 0 9 1 13 16 9 1 0 9 1 9 3 14 9 13 4 2
19 0 11 11 1 11 1 11 9 1 11 9 1 9 1 15 9 13 4 2
18 3 12 0 9 1 13 16 15 14 9 9 9 1 14 13 4 4 2
13 0 9 9 1 14 15 9 1 9 14 13 4 2
6 11 9 1 9 13 2
22 9 1 0 0 9 11 11 11 11 2 11 2 1 9 1 12 9 1 13 4 4 2
38 11 1 12 9 3 11 0 11 2 11 11 1 9 1 9 9 1 11 11 11 1 11 1 9 1 13 4 13 16 15 15 14 9 1 0 14 13 2
37 11 1 9 1 9 13 1 0 9 11 1 13 16 11 11 16 11 11 1 9 1 1 9 13 1 1 0 13 16 15 9 13 1 1 0 13 2
32 9 1 9 1 9 1 11 11 1 13 16 9 1 0 9 0 13 1 9 9 1 9 13 1 1 15 9 0 13 4 4 2
20 11 1 13 16 9 1 9 1 9 1 9 1 9 1 15 9 13 4 4 2
9 15 10 9 1 9 1 9 13 2
22 15 13 16 9 1 9 1 12 14 12 0 9 1 1 9 9 1 9 13 4 4 2
13 15 9 1 10 9 1 1 15 9 13 4 4 2
12 16 11 1 10 9 1 9 1 9 14 13 2
15 11 11 1 13 16 11 7 11 1 9 9 9 13 4 2
26 11 1 9 1 1 11 1 1 9 9 11 11 11 7 0 9 1 11 8 8 11 11 14 3 13 2
16 11 11 1 10 9 1 11 1 9 1 0 9 9 13 4 2
14 11 1 11 1 3 10 9 12 9 13 1 9 13 2
18 11 1 11 9 1 11 11 9 1 9 1 1 1 0 9 13 4 2
17 9 1 12 9 1 13 1 9 13 7 12 9 0 13 4 4 2
20 7 11 9 1 14 0 9 1 1 1 9 7 9 9 0 9 1 0 13 2
24 0 9 1 1 11 9 9 1 11 9 1 11 11 9 1 9 1 1 1 0 9 13 4 2
17 9 1 12 9 1 13 1 9 13 7 12 9 0 13 4 4 2
22 15 1 10 0 9 1 9 1 1 1 12 2 9 1 9 3 14 0 13 4 4 2
13 9 1 11 1 9 1 9 9 9 13 4 4 2
19 11 9 1 14 0 9 1 1 1 9 7 9 9 0 9 1 0 13 2
34 0 9 1 9 1 13 16 11 9 7 11 9 1 1 12 1 1 12 9 9 1 9 13 4 1 1 1 9 9 0 13 4 4 2
13 9 1 12 12 9 9 1 9 1 13 4 4 2
19 0 9 1 11 11 7 0 11 11 1 14 0 2 0 9 13 4 4 2
18 9 1 9 9 1 15 1 9 1 12 9 10 9 0 13 4 4 2
9 0 9 9 1 9 12 9 13 2
20 9 9 1 9 13 4 16 9 12 9 3 14 0 9 1 9 13 4 4 2
23 9 9 1 11 11 1 11 11 1 1 9 1 9 1 1 9 1 9 13 4 4 4 2
16 10 9 1 10 12 9 9 13 4 7 12 9 9 13 4 2
20 0 9 1 11 11 1 10 12 9 9 13 4 7 15 1 12 9 13 4 2
11 9 1 12 9 10 9 0 13 4 4 2
21 11 1 12 9 1 1 1 12 9 9 13 4 4 15 9 1 12 9 10 13 2
9 16 12 9 9 1 9 1 13 2
9 7 11 9 1 1 13 4 4 2
17 15 12 1 1 12 9 9 13 4 15 9 1 12 9 10 13 2
21 0 11 11 1 12 1 1 1 12 9 9 13 4 15 9 1 12 9 10 13 2
21 10 9 1 12 1 1 12 9 9 0 13 4 4 15 9 1 12 9 10 13 2
19 9 9 1 1 9 1 12 1 1 12 9 9 1 9 1 13 4 4 2
16 9 1 0 9 1 1 0 11 1 9 14 10 9 0 13 2
14 9 1 9 1 0 9 9 1 1 3 0 13 4 2
17 7 12 9 1 9 13 7 12 9 1 9 1 14 0 9 13 2
11 9 1 1 9 1 12 9 10 9 13 2
13 11 11 1 10 9 1 1 9 9 3 14 13 2
19 10 3 9 9 1 3 11 11 1 10 9 1 9 1 9 0 13 4 2
23 7 9 9 1 13 13 16 9 1 12 9 3 0 9 1 9 13 1 9 13 4 4 2
13 0 12 9 1 1 15 1 1 9 0 13 4 2
39 0 9 13 1 9 7 12 12 9 1 15 9 1 0 9 13 1 1 11 11 11 11 2 11 2 1 9 1 11 1 0 9 9 11 1 0 13 4 2
13 10 9 3 0 9 9 13 1 11 1 9 13 2
25 9 1 12 9 1 1 11 1 15 9 13 4 7 15 14 12 14 9 1 12 12 9 13 4 2
12 11 1 10 9 1 0 9 9 1 9 13 2
23 9 9 1 13 13 16 10 9 14 11 11 1 13 4 4 15 11 9 1 9 13 4 2
31 11 11 11 11 11 1 11 1 9 1 13 16 15 11 9 9 9 1 9 9 0 13 1 1 1 9 13 1 13 4 2
34 15 13 4 1 16 11 9 9 12 9 13 1 3 12 12 1 9 1 9 10 9 0 13 11 1 13 2 9 10 9 1 9 13 2
11 9 1 15 15 1 1 9 13 4 4 2
43 15 3 2 3 13 4 1 1 10 9 1 13 4 16 15 13 1 1 15 11 11 11 1 1 13 7 14 11 1 13 1 11 9 1 0 9 13 1 9 1 9 13 2
18 16 15 9 9 9 0 13 1 1 10 9 1 15 9 14 13 4 2
23 11 11 11 1 13 16 11 1 9 1 11 9 9 1 0 13 1 1 1 15 9 13 2
13 15 9 2 9 1 9 7 11 1 9 0 13 2
29 9 1 13 16 0 9 13 1 9 1 1 14 9 0 14 13 1 9 1 9 13 1 1 3 0 9 13 4 2
14 11 9 1 11 11 11 1 9 9 1 9 13 4 2
11 13 4 4 16 9 1 9 13 4 4 2
29 15 9 13 4 13 4 4 16 9 9 1 9 7 0 9 1 9 12 1 12 13 4 1 1 10 9 13 4 2
28 0 9 9 11 11 1 13 4 16 9 1 9 9 1 11 11 1 9 1 9 9 11 11 1 9 13 4 2
44 11 1 9 11 11 1 9 1 11 0 11 11 11 11 11 11 11 11 11 11 2 11 2 1 0 12 9 1 11 1 13 16 11 1 11 11 1 9 1 3 9 13 4 2
15 9 9 1 10 9 13 15 1 15 15 9 0 13 4 2
42 11 11 1 11 9 1 9 9 1 9 13 4 11 1 13 16 2 16 9 15 10 9 1 0 9 1 9 13 4 7 10 9 1 9 13 4 16 15 15 0 9 13
17 15 3 13 16 15 10 9 1 10 0 9 1 15 9 13 4 2
24 15 15 14 13 16 10 9 1 15 11 11 1 9 1 0 2 0 9 9 1 9 13 4 2
21 11 11 1 9 9 14 13 1 9 15 13 16 9 1 9 1 9 1 9 13 4
21 9 1 3 13 4 16 10 9 1 11 1 9 9 11 11 1 14 15 9 13 2
20 9 1 9 1 9 11 11 1 11 1 9 2 9 1 11 13 1 9 13 2
13 9 1 1 15 11 11 11 1 9 1 14 13 2
26 14 12 9 1 11 1 0 9 11 11 11 1 11 1 9 1 13 9 1 11 1 9 13 4 4 2
15 3 9 1 9 9 1 11 1 9 13 1 0 13 4 2
19 15 9 1 11 1 13 16 15 11 1 0 11 11 1 9 1 9 13 2
13 11 11 1 9 13 15 9 12 9 1 0 13 2
20 10 3 15 11 11 1 9 1 14 13 7 11 7 11 1 15 9 1 13 2
9 9 1 14 12 9 15 1 13 2
17 15 13 16 11 1 11 11 11 1 9 1 15 9 0 13 4 2
14 15 0 9 13 15 9 1 9 3 13 1 9 13 2
14 15 13 16 15 9 11 11 11 1 9 1 14 13 2
23 15 13 16 11 1 9 13 1 1 15 9 1 9 1 9 1 9 1 9 14 13 4 2
16 11 1 13 16 15 15 9 1 9 9 9 1 13 4 4 2
15 3 10 9 1 1 9 1 15 9 1 15 9 14 13 2
6 15 12 0 9 13 2
29 11 1 9 14 1 11 1 13 4 9 1 1 1 11 1 13 16 15 11 11 7 11 1 9 1 9 14 13 2
7 15 11 1 0 9 13 2
15 11 1 0 9 1 1 1 15 13 16 15 0 9 13 2
23 15 13 16 10 9 1 9 0 13 7 9 2 9 1 13 1 3 15 9 13 9 13 2
15 15 13 16 15 9 14 13 2 16 0 9 1 9 13 2
23 11 1 11 11 1 9 11 11 1 9 9 11 11 1 13 4 9 1 0 13 4 4 2
17 1 11 2 11 1 3 9 1 10 9 1 9 1 0 13 4 2
15 15 9 13 16 15 10 0 0 9 1 14 10 9 13 2
26 9 1 10 9 1 14 0 9 13 16 11 11 1 15 0 9 1 11 9 11 11 1 9 13 4 2
13 11 11 1 13 16 10 9 1 15 9 14 13 2
21 11 9 1 9 13 4 9 9 1 15 9 1 11 9 1 15 9 14 13 4 2
23 11 11 1 9 1 0 9 9 1 9 13 4 15 13 16 9 9 11 1 9 9 13 2
12 11 1 9 1 1 15 11 13 1 9 13 2
21 10 9 13 4 1 16 15 11 11 11 14 13 2 15 13 16 15 0 9 13 2
9 15 2 11 1 15 9 14 13 2
27 11 11 11 9 11 11 11 1 13 16 11 9 9 1 9 1 9 11 1 11 9 1 9 1 14 13 2
12 15 13 16 10 9 9 1 11 9 14 13 2
18 11 1 9 1 9 1 11 1 13 16 0 9 11 1 14 0 13 2
14 11 1 9 11 1 9 1 13 1 1 13 4 4 2
27 15 9 13 4 13 16 15 9 1 1 7 3 1 15 14 9 1 11 11 1 9 11 1 9 14 13 2
25 11 1 13 16 10 9 15 9 9 1 11 9 1 1 15 14 9 1 0 9 1 9 14 13 2
13 15 9 1 10 9 1 0 9 1 9 13 4 2
26 11 1 13 16 16 9 1 15 9 1 9 13 4 16 11 11 11 2 11 2 1 15 9 11 13 2
23 15 9 13 4 13 16 11 1 9 0 13 4 4 15 9 1 12 1 10 9 14 13 2
10 15 13 16 11 11 1 9 13 4 2
14 11 1 12 9 1 9 1 11 1 9 13 4 4 2
27 15 13 16 11 7 11 1 1 9 7 9 1 1 9 1 11 0 13 4 7 15 0 9 11 1 13 2
21 11 1 13 16 9 1 9 13 4 4 16 10 9 1 1 11 7 11 0 13 2
36 9 9 11 7 11 1 9 1 9 1 12 0 9 1 9 13 11 1 1 13 4 4 7 15 15 12 0 9 1 9 1 9 13 4 4 2
16 15 1 11 11 1 9 1 9 1 9 10 0 13 4 4 2
23 9 11 11 3 1 11 11 1 9 13 0 9 1 0 13 1 9 1 9 13 4 4 2
14 9 1 11 1 0 9 1 0 13 1 9 0 13 2
10 15 0 3 11 9 1 9 13 4 2
32 13 4 4 16 0 0 9 1 10 9 1 9 12 12 9 13 7 15 11 1 0 9 11 11 11 11 1 9 1 9 13 2
21 10 9 9 1 0 9 9 11 11 1 0 9 11 11 1 0 12 9 1 13 2
30 15 13 16 10 9 1 12 0 9 1 0 2 0 9 1 9 13 4 4 2 15 15 0 13 1 9 13 4 4 2
15 15 13 16 15 1 12 9 1 9 12 9 1 1 13 2
15 11 1 9 1 10 9 1 11 1 11 1 13 4 4 2
11 15 9 12 9 13 7 9 12 9 13 2
16 9 11 1 13 16 15 10 9 1 15 9 1 1 13 4 2
22 15 9 13 16 9 1 9 1 1 10 0 9 1 9 13 11 1 1 13 4 4 2
19 15 13 4 16 9 9 9 1 1 1 9 13 7 9 1 3 0 13 2
14 15 13 16 15 1 1 9 1 9 0 13 4 4 2
15 0 9 1 9 1 9 11 1 11 11 11 11 1 13 2
16 10 9 1 9 9 1 9 9 1 9 1 13 1 9 13 2
40 11 11 1 0 9 1 1 9 1 13 4 1 9 1 9 9 1 9 1 9 14 13 2 7 9 1 9 9 7 9 9 1 0 9 1 9 13 4 4 2
21 11 11 1 0 9 1 9 1 1 1 9 1 9 9 1 9 1 0 9 13 2
14 9 1 9 11 11 1 15 9 1 0 13 4 4 2
32 7 11 11 1 13 13 16 0 12 9 1 11 11 1 9 1 1 9 1 9 1 9 1 9 10 9 1 3 13 4 4 2
22 10 3 11 11 1 9 1 9 1 1 12 12 12 9 1 9 9 1 0 13 4 2
17 15 1 0 9 1 1 9 1 9 9 13 1 15 9 14 13 2
24 11 11 1 10 9 1 1 0 9 1 0 9 9 2 11 2 1 15 9 1 9 14 13 2
15 0 9 9 1 9 1 14 9 1 9 0 13 4 4 2
16 0 9 9 1 9 1 1 9 1 14 0 13 1 9 13 2
22 10 9 13 16 11 11 10 9 1 9 1 15 14 9 1 13 1 1 0 14 13 2
29 16 2 9 1 11 11 1 9 9 7 9 9 1 9 9 1 12 1 12 9 1 9 1 0 9 13 4 4 2
44 11 11 1 9 9 7 9 9 1 13 4 0 9 1 1 15 1 9 13 1 1 9 1 0 9 1 10 9 1 9 13 4 2 15 1 1 9 1 9 1 9 13 4 2
22 9 9 2 11 11 2 1 9 1 0 9 9 11 11 1 12 9 9 0 13 4 2
13 15 1 11 11 1 12 12 9 1 9 13 4 2
19 9 1 15 9 1 0 9 9 1 13 4 15 9 1 10 0 9 13 2
33 11 11 1 9 7 9 11 11 11 1 11 1 13 16 11 11 1 11 11 1 9 13 1 1 11 2 11 1 15 9 13 4 2
17 11 7 11 11 1 10 0 0 9 1 1 9 1 9 13 4 2
19 15 13 16 11 11 1 12 0 9 1 15 11 11 1 14 12 9 13 2
24 16 2 0 9 9 1 1 0 9 9 15 0 9 9 1 0 12 9 1 9 13 4 4 2
33 11 9 1 11 1 9 1 1 9 1 11 9 1 9 11 11 1 13 4 16 9 7 11 1 9 1 9 1 13 15 9 13 2
26 15 13 16 15 11 1 1 1 9 1 9 1 9 14 13 2 16 15 1 3 13 13 1 9 13 2
12 15 13 16 15 9 12 0 9 1 9 13 2
22 11 1 11 1 9 1 9 13 4 11 11 1 15 0 9 1 7 12 0 9 13 2
15 11 1 13 16 9 1 9 7 9 1 1 9 13 4 2
19 16 0 9 1 9 1 9 14 13 1 15 9 15 9 13 1 9 13 2
23 15 1 1 13 4 9 1 13 4 15 13 2 2 15 14 10 14 9 0 13 0 13 2
9 15 9 13 4 7 15 9 15 13
25 0 7 0 9 13 1 1 15 9 9 1 14 9 13 4 13 16 9 1 9 1 9 13 4 2
24 3 11 11 1 11 1 11 1 1 9 1 9 13 4 11 1 9 1 0 13 1 9 13 2
39 11 11 1 9 1 13 16 3 0 9 2 0 9 7 9 1 11 1 15 13 4 0 13 16 9 1 10 14 9 13 15 0 15 12 9 1 9 13 2
22 15 13 16 10 9 11 1 9 1 9 13 4 4 15 3 14 15 9 1 9 13 2
15 15 9 13 16 11 9 1 13 9 1 0 14 13 4 2
9 15 15 9 1 9 1 9 13 2
30 11 11 11 1 15 9 9 7 11 9 11 11 1 9 1 13 4 13 16 15 9 1 15 1 1 15 9 14 13 2
13 11 1 13 16 9 1 9 2 9 13 4 4 2
43 0 11 9 1 11 1 11 9 1 9 9 9 2 9 2 1 9 11 11 1 11 11 9 1 1 1 10 9 13 1 1 9 2 9 7 0 9 1 9 13 4 4 2
35 0 9 11 11 1 9 1 9 13 4 9 11 11 11 1 9 1 11 1 9 2 9 2 9 9 7 11 11 11 13 1 9 13 4 2
13 0 9 1 9 1 1 11 1 9 13 4 4 2
42 9 9 1 13 16 9 1 11 9 1 11 7 0 9 1 0 13 1 1 1 10 9 13 1 1 9 1 9 2 9 2 9 9 7 11 11 11 13 1 9 13 2
25 0 9 1 9 1 13 16 11 1 9 7 9 9 1 0 13 10 9 1 9 1 9 13 4 2
17 15 9 1 9 13 1 1 9 1 11 1 9 13 1 9 13 2
20 0 11 11 7 11 1 0 9 11 11 1 0 9 1 0 13 4 4 4 2
18 11 9 1 15 1 0 11 0 13 4 1 3 15 0 13 4 4 2
29 0 13 16 11 11 1 12 9 9 1 9 1 11 1 11 1 12 9 1 11 11 1 9 1 9 13 4 4 2
15 15 1 11 1 11 1 11 11 1 1 0 13 4 4 2
16 3 1 11 1 0 0 9 1 15 0 9 1 13 4 4 2
29 11 11 1 11 11 11 1 1 11 9 11 11 1 9 1 1 11 9 11 1 1 9 0 13 1 9 13 4 2
25 11 1 13 16 11 1 9 11 1 15 9 1 13 16 11 15 9 1 9 13 1 1 0 13 2
16 15 13 16 11 11 11 14 15 9 1 9 1 1 0 13 2
35 11 1 13 16 15 11 11 11 0 13 1 9 1 11 9 1 9 1 1 0 13 1 3 11 11 1 14 15 9 9 0 13 4 4 2
22 9 1 0 9 1 0 9 1 9 13 4 11 11 1 12 0 9 1 9 13 4 2
9 10 9 13 9 9 11 11 1 2
23 11 1 11 1 1 9 13 16 9 1 3 10 9 13 1 9 2 9 1 0 9 13 2
15 10 9 1 10 9 1 11 1 9 1 0 13 0 13 2
12 15 13 16 3 14 15 2 9 2 1 13 2
21 9 1 9 1 1 1 15 13 16 10 9 10 13 4 16 9 1 9 13 4 2
13 9 1 15 9 9 0 13 1 10 9 14 13 2
18 11 1 15 0 9 1 9 1 1 11 1 11 1 1 0 13 4 2
17 9 11 11 14 10 9 13 15 11 1 11 11 1 9 13 4 2
11 7 10 9 1 15 9 0 13 4 4 2
32 15 9 1 9 1 9 13 4 15 13 16 15 15 9 2 9 11 11 7 15 3 13 1 9 1 9 1 14 15 14 13 2
22 9 1 11 11 1 13 16 15 0 9 13 16 11 0 9 1 1 9 1 9 13 2
14 11 11 1 9 1 9 11 1 12 0 9 9 13 2
30 15 13 16 15 11 1 1 1 10 14 13 7 11 1 0 9 13 7 15 9 13 1 1 15 9 9 1 14 13 2
29 11 11 11 2 11 2 1 11 2 11 9 9 13 1 1 11 9 11 11 7 15 9 11 11 1 9 13 4 2
28 9 9 1 1 11 1 1 0 11 9 1 13 1 1 9 1 11 9 11 11 1 14 9 13 4 4 4 2
42 11 9 2 9 9 2 11 11 1 1 1 12 0 9 9 1 13 4 16 9 1 9 11 11 1 11 1 0 9 9 1 13 1 1 11 7 11 1 9 13 4 2
18 2 11 11 2 1 1 9 1 11 1 14 9 13 4 1 9 13 2
32 0 9 1 1 11 1 13 1 0 9 7 15 1 12 12 0 9 1 13 1 1 10 0 9 9 1 14 0 13 4 4 2
39 9 2 9 2 9 11 11 2 11 7 11 1 15 9 9 1 9 1 11 1 9 1 9 14 13 1 1 11 1 11 11 11 7 11 1 9 13 4 2
16 9 11 11 11 1 13 16 15 9 1 0 9 1 9 13 2
7 2 9 15 15 14 13 4
31 11 0 9 1 9 11 11 11 1 13 16 0 9 1 1 1 12 9 1 9 13 1 15 9 1 9 1 9 13 4 2
18 16 11 14 9 1 0 13 7 9 1 9 13 16 15 14 9 13 2
15 15 13 16 11 9 1 15 1 14 9 1 9 14 13 2
36 16 11 9 1 0 14 13 4 16 15 0 13 4 16 11 9 1 9 1 0 13 4 4 7 14 12 14 9 1 9 1 9 13 4 4 2
41 11 1 9 13 16 9 1 11 11 1 10 9 1 9 1 1 1 12 9 13 4 15 1 11 11 7 15 12 9 9 1 9 13 4 7 15 1 9 13 4 2
14 15 9 1 11 11 1 12 9 13 1 14 9 13 2
17 0 13 16 12 9 1 11 11 2 11 1 9 13 4 4 4 2
53 11 11 2 11 11 2 11 11 7 11 11 1 9 13 1 9 1 9 1 9 13 4 11 1 13 16 2 15 0 14 9 1 9 13 16 9 1 10 9 9 1 11 11 1 9 1 0 9 1 0 14 13 2
26 11 1 11 11 11 11 1 9 1 0 9 11 11 11 11 2 11 2 1 0 9 1 0 13 4 2
29 9 9 1 11 9 9 1 11 11 1 9 0 13 1 3 0 9 14 15 0 9 10 9 1 9 13 4 4 2
20 9 11 11 1 1 14 12 9 1 9 1 15 0 9 1 10 9 13 4 2
15 0 9 1 9 13 4 15 11 9 1 9 1 13 4 2
22 9 1 0 9 1 0 9 7 9 9 1 9 14 0 9 1 1 0 9 1 13 2
51 11 9 9 0 11 9 1 0 11 9 1 0 0 9 1 11 1 11 9 7 9 1 0 9 11 11 11 1 11 1 9 13 4 1 9 13 2 15 11 1 11 11 7 11 1 11 11 1 9 13 2
41 9 1 1 11 1 9 12 9 14 9 1 15 9 13 4 16 9 9 11 11 11 10 9 1 9 1 12 12 9 1 10 9 1 9 1 9 13 4 4 4 2
55 9 11 2 11 1 1 13 4 11 9 1 11 1 11 1 11 11 2 9 11 11 11 2 11 11 11 2 11 11 11 2 11 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 7 11 11 11 13 2
19 9 1 3 13 4 9 1 11 11 11 7 11 11 11 1 9 0 13 2
20 11 1 9 13 1 9 1 1 0 9 11 11 11 0 13 9 1 13 4 2
20 11 11 1 11 11 11 1 9 1 15 9 1 0 14 13 4 1 9 13 2
48 11 11 11 11 11 1 9 7 11 1 9 1 9 11 11 11 1 11 11 11 1 0 9 13 4 1 9 13 4 13 16 10 9 1 9 13 4 4 2 15 1 11 1 9 14 14 13 2
18 9 1 11 1 11 11 11 11 11 2 11 1 9 1 0 13 4 2
19 15 1 9 1 10 0 9 1 12 9 9 1 9 1 9 13 4 4 2
9 15 10 10 9 14 13 4 4 2
25 10 9 1 0 9 12 9 1 10 13 2 15 10 9 1 14 10 9 1 0 9 14 0 13 2
14 16 9 1 10 9 1 9 1 15 13 4 9 13 2
26 9 1 10 9 1 9 1 1 11 11 11 11 11 1 13 16 15 12 10 0 9 13 4 4 4 2
12 15 13 16 0 9 0 13 9 1 9 13 2
11 15 9 1 15 9 14 0 2 0 13 2
11 10 9 1 0 9 12 9 1 10 13 2
20 10 9 1 10 9 1 1 13 1 9 1 14 10 9 1 9 14 0 13 2
26 15 13 16 10 9 9 1 12 12 9 1 9 13 2 7 3 14 15 0 9 1 0 13 4 4 2
26 15 1 0 9 12 9 1 13 4 4 2 7 9 1 9 13 16 15 1 14 15 0 13 4 4 2
11 9 1 10 9 1 11 11 1 0 13 2
35 9 1 9 13 4 15 13 16 15 9 1 9 1 9 1 0 9 0 13 7 15 10 9 1 9 1 13 4 14 0 9 13 4 4 2
22 15 13 16 15 15 15 14 13 16 10 9 1 0 13 1 9 7 9 0 13 4 2
27 15 13 16 9 1 9 1 1 16 9 9 1 1 9 14 13 4 16 15 10 14 9 1 9 9 13 2
23 0 9 9 9 0 13 1 1 15 9 9 1 11 11 2 2 11 2 1 9 14 13 2
30 11 11 11 11 11 2 11 2 1 11 1 15 14 10 0 9 1 9 13 4 2 15 0 9 9 1 10 9 13 2
30 9 1 9 1 0 2 0 13 1 1 2 0 0 9 2 1 9 1 0 7 0 2 0 0 2 9 0 13 4 2
39 9 1 9 1 13 4 4 16 10 13 10 9 9 9 1 3 13 2 10 9 13 2 15 9 7 9 0 13 7 9 1 9 1 0 13 1 9 13 2
40 12 0 0 9 1 3 9 1 1 2 0 9 2 1 9 0 13 9 13 4 4 2 3 9 1 15 9 15 0 13 1 9 13 9 1 9 13 4 4 2
25 0 9 1 15 9 0 13 14 10 9 1 9 1 13 1 1 0 9 7 9 0 13 4 4 2
40 9 9 1 9 9 2 1 9 0 13 4 9 1 15 14 13 4 16 0 9 0 7 0 9 1 15 14 0 9 15 9 1 14 15 9 9 14 13 4 2
30 9 1 13 4 4 16 0 9 2 9 9 7 0 9 13 4 9 1 9 1 9 1 9 7 9 1 9 13 4 2
40 11 11 9 7 0 11 11 11 11 1 11 1 13 16 15 11 1 9 1 9 1 3 14 12 9 1 1 11 2 11 9 7 9 9 1 9 1 9 13 2
29 11 1 13 16 11 11 1 10 9 13 1 9 1 15 12 9 1 1 11 11 11 7 11 9 11 11 1 13 2
21 11 0 11 11 11 1 1 0 9 1 9 13 1 3 9 1 9 13 4 4 2
26 11 11 11 11 1 9 1 14 11 1 13 9 1 15 13 16 15 15 1 9 9 0 13 4 4 2
27 0 13 16 11 1 15 9 1 13 4 16 11 11 1 10 9 13 1 9 1 9 7 9 1 9 13 2
23 15 1 11 1 13 16 11 11 9 1 0 9 1 9 9 9 13 1 9 13 4 4 2
15 15 13 16 15 1 1 9 9 1 9 13 4 4 4 2
31 14 12 12 9 1 15 12 9 11 1 9 1 1 9 13 15 9 1 9 1 11 9 11 1 9 1 9 13 4 4 2
13 9 9 9 11 11 11 1 11 1 10 9 13 2
20 11 1 9 11 11 11 1 11 11 1 1 9 1 9 1 0 13 4 4 2
41 9 1 9 1 1 11 1 11 11 9 11 11 1 12 12 9 1 9 11 11 11 11 1 9 1 9 1 1 11 1 13 1 9 2 9 1 9 13 4 4 2
19 11 11 1 9 1 11 14 11 9 13 1 1 11 1 3 13 4 4 2
24 11 2 11 2 1 11 11 1 13 4 11 14 11 10 9 11 1 9 1 1 9 13 4 2
26 7 9 9 1 15 14 11 13 7 14 11 14 11 1 10 9 13 15 9 13 1 9 13 4 4 2
19 15 13 4 4 16 11 1 0 13 1 1 12 12 9 1 9 13 4 2
25 0 9 11 11 1 11 1 9 13 7 11 9 1 0 11 11 11 1 1 9 13 1 9 13 2
10 11 9 1 9 1 9 13 4 4 2
23 9 9 1 1 9 1 13 4 9 1 13 2 7 11 15 1 9 13 1 1 14 13 2
6 0 9 3 9 13 2
24 10 9 9 1 12 12 9 13 1 15 9 13 16 12 12 12 12 9 1 9 0 13 4 2
23 10 9 9 1 9 13 1 9 1 13 4 11 9 1 11 11 11 1 1 13 1 13 2
14 9 1 15 9 13 7 9 1 1 15 13 4 4 2
22 11 1 13 16 15 11 1 10 9 13 4 11 9 0 9 1 9 1 13 4 4 2
28 11 1 11 11 1 11 9 11 11 1 0 9 13 1 9 13 1 9 1 9 1 15 11 1 9 13 4 2
22 9 1 11 11 1 9 11 11 1 11 11 1 10 9 15 11 1 9 1 13 4 2
30 15 13 16 0 9 13 1 9 13 1 11 11 1 9 1 9 1 15 12 9 1 1 15 9 13 1 1 13 4 2
14 9 1 11 1 11 1 9 1 0 9 0 13 4 2
31 11 11 1 13 16 9 1 9 2 9 9 7 0 0 9 1 13 4 13 4 16 9 11 11 1 11 1 9 13 4 2
12 15 13 16 9 10 9 1 15 0 9 13 2
10 11 13 4 16 11 15 15 9 13 2
11 15 10 9 1 11 1 0 13 4 4 2
19 11 9 13 1 3 9 11 11 15 0 9 1 9 11 11 1 9 13 2
17 15 0 10 9 1 14 11 11 1 9 1 13 1 9 1 13 2
13 11 1 0 2 0 9 15 10 9 1 0 13 2
20 15 11 2 11 7 0 11 11 15 9 1 9 13 1 9 13 4 4 4 2
31 11 9 1 1 11 1 10 9 1 0 9 10 0 9 13 13 16 15 9 7 0 9 1 9 1 9 1 1 0 13 2
25 15 10 9 13 15 11 1 0 9 13 4 7 0 12 9 1 12 1 10 9 1 9 13 4 2
24 0 9 15 13 16 11 9 13 1 3 14 10 9 1 9 1 9 9 1 9 13 14 4 2
30 11 1 10 9 1 11 1 9 9 1 14 13 13 4 4 4 15 9 1 9 1 9 13 10 0 0 13 4 4 2
13 15 10 9 1 9 1 9 1 9 13 4 4 2
17 0 9 14 9 1 9 1 9 0 13 1 9 3 13 4 4 2
15 9 1 1 9 1 9 9 1 10 13 4 1 9 13 2
25 10 9 13 16 11 11 1 9 1 1 11 9 7 0 2 0 9 1 1 10 9 13 4 4 2
19 11 11 11 11 14 9 1 9 13 1 3 9 13 1 9 13 13 4 2
27 9 2 9 1 9 1 11 11 1 9 13 4 1 11 9 11 11 11 1 15 10 9 1 9 14 13 2
16 13 15 16 12 0 11 11 11 13 11 1 9 1 13 4 2
23 11 15 0 13 16 9 2 9 1 0 13 1 11 11 1 9 1 11 1 9 14 13 2
18 15 15 15 1 11 11 2 11 11 1 9 13 14 0 13 4 4 2
23 15 0 9 1 11 0 9 1 1 9 2 9 1 2 9 2 9 13 1 13 4 4 2
22 11 10 9 11 1 11 11 11 11 11 13 7 11 1 15 10 9 9 13 4 4 2
17 15 1 14 11 11 1 9 11 9 13 14 3 0 13 4 4 2
29 9 2 9 1 15 9 1 11 10 9 0 13 4 4 16 15 11 1 3 14 9 1 13 1 9 13 4 4 2
11 11 11 1 10 9 15 1 14 13 4 2
16 2 11 11 2 1 15 13 2 0 3 9 11 1 14 13 4
24 11 1 13 1 3 15 15 15 9 13 16 15 13 16 15 13 16 15 1 9 1 9 13 2
27 15 11 1 9 1 9 13 9 1 9 13 4 7 10 9 1 11 9 1 1 0 9 0 13 4 4 2
23 11 11 11 11 1 9 13 1 1 11 9 1 1 11 1 9 13 10 0 13 4 4 2
8 10 9 1 14 9 13 4 2
12 11 1 9 13 7 11 13 11 1 13 4 2
21 11 13 4 2 2 15 9 9 15 14 13 4 16 15 1 9 1 9 14 13 2
16 3 2 15 11 1 9 13 7 9 15 11 1 0 9 13 2
24 11 13 4 2 2 10 9 15 11 1 0 13 4 4 10 9 14 15 1 9 2 9 13 4
15 11 1 15 13 16 15 11 1 14 15 15 9 13 4 2
23 15 15 13 16 9 2 9 1 9 13 9 1 9 13 16 0 9 2 9 0 9 13 2
22 15 15 9 1 0 13 7 15 9 1 14 15 9 2 9 1 9 0 13 4 4 2
29 0 9 1 3 2 3 13 11 11 11 1 9 11 11 11 11 1 9 1 11 11 1 0 9 13 1 13 4 2
30 7 10 9 1 9 11 1 13 1 15 9 11 11 1 0 13 4 15 9 7 0 15 9 1 13 1 9 13 4 2
12 11 9 1 0 9 1 9 1 14 0 13 2
16 11 11 1 9 1 1 11 9 1 11 1 9 13 4 4 2
46 9 11 11 11 7 9 11 11 11 1 9 1 11 1 11 1 9 11 11 1 9 13 16 9 1 9 11 9 1 1 11 1 13 4 7 11 1 9 1 9 11 9 1 13 4 2
31 9 1 11 9 1 9 13 16 11 1 0 9 13 4 7 11 1 9 1 1 9 7 0 9 1 1 13 1 1 13 2
38 9 1 11 9 1 9 1 13 16 15 9 9 1 10 9 1 9 13 16 16 11 1 9 11 9 1 13 4 4 16 11 9 1 9 14 14 13 2
22 11 9 1 9 11 11 1 13 16 15 10 9 1 9 9 11 11 11 1 9 13 2
14 11 1 15 1 13 9 1 11 9 1 9 13 4 2
27 9 1 9 15 9 1 9 1 14 0 9 13 4 13 16 15 10 9 1 0 7 0 9 14 13 4 2
23 11 1 11 11 1 9 1 11 11 9 1 10 0 9 1 9 13 4 0 13 4 4 2
15 11 11 11 11 1 11 1 12 9 1 9 13 4 4 2
14 15 1 1 15 11 11 1 14 9 1 13 4 4 2
33 0 13 16 11 11 11 1 9 1 0 9 1 9 1 9 1 11 11 11 1 11 7 11 11 14 11 11 1 0 13 4 4 2
13 11 11 7 11 11 11 1 9 1 9 13 4 2
13 12 9 1 9 1 1 11 11 1 9 13 4 2
13 0 13 4 9 1 1 11 9 1 9 13 4 2
21 0 9 1 1 0 9 1 11 1 12 0 9 1 1 11 1 15 9 0 13 2
24 11 11 11 7 11 11 11 11 11 1 13 10 9 1 9 14 9 9 7 9 13 1 13 2
9 7 11 9 1 15 9 14 13 2
28 1 15 11 11 11 11 11 11 11 1 9 1 12 9 1 9 9 1 9 13 7 10 9 1 15 9 13 2
17 15 10 9 14 0 14 13 7 3 15 9 13 1 9 14 13 2
19 9 1 9 11 11 1 9 9 9 13 11 11 11 1 9 13 1 13 2
16 15 9 1 1 14 9 10 9 1 0 9 1 9 0 13 2
21 9 1 9 1 1 9 1 9 9 1 9 13 15 1 9 1 15 0 13 4 2
26 0 9 1 9 9 11 11 1 1 14 9 9 13 1 11 11 11 1 1 12 9 1 0 13 4 2
8 15 12 9 7 12 9 13 2
9 15 9 12 9 0 13 4 4 2
19 0 13 1 1 0 9 11 11 2 11 2 11 7 11 11 14 0 13 2
44 11 9 0 13 4 1 9 1 0 0 9 13 4 11 11 11 1 11 1 13 16 9 1 9 2 9 1 9 1 16 15 1 9 0 13 16 15 10 9 1 1 9 13 2
17 11 1 0 13 4 1 9 1 11 11 11 1 12 9 0 13 2
20 11 1 13 16 15 10 0 9 1 9 1 13 4 9 0 13 1 9 13 2
22 11 11 1 9 7 11 2 9 9 1 11 11 1 9 1 9 1 14 10 9 13 2
25 11 1 12 9 9 1 11 1 13 16 11 1 9 15 9 1 1 9 1 13 1 1 0 13 2
19 15 13 16 9 9 1 1 9 1 9 2 9 1 15 1 0 9 13 2
47 3 11 1 9 9 11 11 11 2 11 1 9 9 11 11 11 7 11 2 11 2 1 9 9 11 11 1 12 0 9 9 1 13 16 11 11 1 11 13 4 1 0 9 13 4 4 2
40 11 1 9 1 9 2 9 13 7 11 9 1 9 1 9 13 4 1 1 1 10 9 1 13 16 16 11 1 1 0 9 13 16 11 0 9 15 14 13 2
36 0 9 1 11 7 11 2 11 2 9 1 13 1 3 11 11 7 11 1 13 16 11 11 11 1 0 11 11 11 1 9 1 9 13 4 2
19 15 15 14 10 9 1 11 11 11 1 9 1 9 13 1 1 13 4 2
12 11 11 1 10 9 9 1 9 1 14 13 2
27 9 1 9 9 1 11 7 9 2 3 1 9 1 9 1 15 9 1 13 9 2 9 1 8 13 4 2
11 15 9 1 9 9 1 9 13 4 4 2
34 9 1 0 9 1 1 0 9 15 13 4 4 9 1 0 9 1 9 13 10 13 4 4 7 15 15 9 1 15 9 13 4 4 2
41 11 1 11 11 8 13 12 9 2 9 1 1 11 2 11 2 11 1 12 9 1 15 9 1 0 13 16 0 9 15 13 14 9 1 9 0 13 4 4 4 2
7 9 1 1 0 14 13 2
29 10 9 1 3 13 0 9 1 13 16 3 13 2 9 13 7 16 9 14 13 16 9 1 9 1 9 13 4 2
4 9 10 13 2
11 15 0 13 16 9 1 9 13 4 4 2
9 0 9 1 9 0 13 4 4 2
11 9 9 9 7 10 14 9 15 9 13 2
13 9 1 1 0 9 1 14 10 9 1 9 13 2
24 0 9 1 14 10 0 9 1 13 4 1 9 13 7 10 9 1 9 0 9 14 13 4 2
31 11 2 11 2 11 2 11 2 11 2 11 7 11 11 1 0 9 11 2 9 9 2 11 11 11 1 11 1 13 4 2
21 10 9 1 11 11 1 9 9 2 11 11 2 11 1 11 11 1 13 4 4 2
8 15 9 9 11 7 11 13 2
13 9 1 9 1 1 11 11 1 11 1 9 13 2
10 11 11 1 15 11 11 11 11 13 2
19 9 1 1 15 0 9 1 3 0 9 13 7 15 11 1 9 13 4 2
22 9 13 4 16 10 9 1 1 11 7 11 1 9 9 1 9 13 9 13 4 4 2
19 15 3 13 16 9 15 9 1 1 13 4 14 9 1 1 13 4 4 2
8 7 2 3 1 9 14 13 2
17 9 1 15 13 1 12 2 12 9 1 1 14 9 13 4 4 2
6 9 13 4 4 4 2
8 15 9 1 9 13 4 4 2
16 11 11 11 11 11 1 9 1 3 9 13 1 9 13 4 2
24 7 2 9 1 1 3 0 9 15 13 16 9 1 13 4 9 1 9 1 15 0 13 4 2
32 11 11 1 13 1 1 11 11 11 11 11 2 11 2 9 1 12 11 11 11 2 11 2 11 2 11 2 9 13 4 4 2
21 11 11 11 1 12 0 9 1 13 13 16 0 9 11 11 1 9 13 4 4 2
13 16 15 15 0 9 1 15 9 14 13 4 4 2
41 11 1 11 1 11 11 11 2 11 11 11 11 11 1 9 13 4 11 11 1 13 16 9 9 1 11 11 1 9 13 1 3 15 9 7 9 13 0 13 4 2
13 15 1 14 9 9 1 14 9 1 9 13 4 2
14 15 1 9 2 9 7 9 1 9 1 9 13 4 2
13 15 3 13 16 9 3 9 2 9 7 9 13 2
11 15 9 1 9 13 16 15 3 9 13 2
21 7 15 15 1 10 14 0 9 13 16 9 1 13 9 1 9 1 15 0 13 4
33 15 13 16 11 1 11 11 13 1 9 1 1 11 11 11 12 12 9 9 1 13 4 4 7 12 9 1 14 0 13 4 4 2
25 15 3 13 16 2 3 9 10 9 1 13 16 10 9 11 1 9 13 15 15 15 0 13 4 2
18 15 1 15 0 13 1 14 9 13 16 10 9 1 9 14 13 4 2
34 2 11 11 11 11 11 2 11 2 1 9 11 11 11 1 13 16 11 2 11 2 11 7 11 1 11 11 11 2 11 11 13 4 2
24 9 9 11 11 11 1 13 4 9 7 9 1 1 9 1 9 1 13 1 9 13 4 4 2
19 3 0 3 9 9 11 11 1 9 14 9 1 9 1 9 13 4 4 2
11 15 14 9 1 9 2 9 13 14 4 2
21 16 2 11 1 9 1 1 15 1 9 9 1 13 9 1 15 15 9 14 13 2
41 9 11 11 11 2 11 2 1 12 9 2 11 1 12 9 7 11 11 2 11 2 1 12 9 1 1 9 1 13 9 1 13 1 15 9 1 9 13 4 4 2
31 16 9 1 15 9 1 1 10 9 13 4 15 0 9 14 13 1 1 9 1 15 11 11 1 0 9 13 1 13 4 2
33 9 1 9 1 13 4 16 15 13 16 0 9 7 9 1 10 9 1 9 1 0 13 4 2 15 15 11 11 11 13 4 4 2
49 9 1 0 9 14 0 13 1 13 4 4 16 15 9 13 4 4 16 9 7 9 2 15 1 9 1 9 13 4 2 15 9 7 9 13 1 3 11 11 11 1 0 13 7 15 1 1 13 2
48 16 15 9 7 9 13 1 3 9 1 15 9 13 4 15 14 9 9 15 1 9 13 7 16 9 7 9 9 1 1 14 11 11 11 1 13 16 15 1 9 1 9 1 9 9 9 13 2
42 9 1 13 13 16 0 9 9 11 11 1 11 11 11 1 13 9 13 1 10 9 13 4 4 15 15 13 1 14 13 7 10 9 1 10 9 1 9 13 4 4 2
16 15 1 9 1 1 14 12 14 9 1 9 1 9 13 4 2
13 15 9 13 4 16 9 1 10 9 1 13 4 2
18 0 3 9 9 11 11 1 9 14 9 1 9 1 9 13 4 4 2
33 11 1 9 7 9 1 14 12 9 1 9 1 12 9 11 1 13 4 15 11 1 9 13 4 4 16 15 0 11 1 1 13 2
25 11 1 9 13 16 15 9 1 9 1 9 1 11 11 11 11 11 7 0 9 1 9 13 4 2
24 9 1 3 14 11 1 1 1 11 1 1 1 15 9 13 4 2 15 15 1 9 13 4 2
20 9 9 1 0 11 11 11 11 1 9 1 0 11 11 2 11 2 13 4 2
52 0 0 9 1 1 12 9 1 1 11 11 2 11 2 1 0 13 1 3 0 9 13 1 9 11 11 11 1 9 1 1 10 9 1 9 13 4 16 11 11 2 11 2 1 9 9 1 0 13 4 4 2
23 15 0 14 13 1 15 9 1 9 13 4 16 15 9 1 14 0 11 11 13 4 4 2
11 7 15 11 1 15 9 0 13 4 4 2
41 11 11 2 11 2 1 9 11 11 1 9 1 13 16 9 1 15 0 13 4 16 11 1 15 9 0 13 4 4 7 9 1 10 0 9 1 0 13 4 4 2
18 11 1 11 11 1 13 15 9 1 15 9 0 13 1 9 13 4 2
27 9 1 11 11 1 11 1 13 13 16 9 1 15 9 9 13 4 4 7 10 9 1 0 13 4 4 2
14 9 1 1 9 1 15 1 9 11 1 14 13 4 2
33 0 13 16 11 1 9 1 0 13 1 3 11 11 11 11 1 9 13 4 4 7 15 1 9 1 11 1 9 9 9 14 13 2
13 11 1 1 9 1 12 9 14 0 13 4 4 2
17 9 1 11 7 11 1 1 15 9 1 9 1 9 1 9 13 2
23 11 1 13 16 11 7 0 9 1 9 1 9 9 1 9 9 1 1 15 14 0 13 2
20 11 9 9 1 9 1 1 9 7 0 0 9 1 9 9 1 9 0 13 2
27 0 9 1 0 13 4 16 11 1 9 1 14 11 11 2 11 2 11 2 11 7 11 1 9 13 4 2
9 10 9 1 0 9 9 9 13 2
20 9 3 14 11 7 11 1 9 9 9 1 1 14 10 9 1 9 9 13 2
36 9 1 1 9 1 11 1 1 14 10 9 1 13 4 16 15 10 9 1 9 9 9 1 13 15 1 0 0 9 0 12 9 1 0 13 2
17 9 1 15 10 9 1 9 1 9 1 9 13 1 9 13 4 2
17 9 1 13 16 9 1 3 10 9 11 11 1 9 9 1 13 2
22 3 11 11 1 9 11 11 0 9 1 9 1 13 9 1 9 9 1 13 4 4 2
30 13 4 4 4 16 9 9 9 11 0 9 11 11 1 9 13 4 4 7 15 15 10 9 1 9 14 13 4 4 2
17 9 1 9 1 13 16 11 11 1 12 12 0 0 9 0 13 2
19 15 1 12 12 9 1 9 13 4 4 4 7 15 9 0 13 4 4 2
12 11 1 0 0 9 1 12 12 9 0 13 2
21 11 1 0 9 11 1 9 1 9 9 1 9 11 1 9 1 12 9 1 13 2
37 0 11 1 1 14 9 1 9 9 2 11 7 11 1 14 10 9 1 0 9 13 7 9 1 11 9 1 9 1 9 1 13 9 1 9 13 2
21 11 11 11 11 1 12 9 1 10 9 1 9 13 2 7 9 15 0 14 13 2
28 9 1 9 1 3 10 9 13 7 3 11 1 9 1 9 13 16 9 9 9 1 0 9 1 1 0 13 2
19 15 1 12 9 1 9 1 9 0 13 4 7 10 9 1 9 13 4 2
26 9 1 11 1 11 11 11 1 9 13 4 13 16 10 9 1 11 11 11 1 9 0 13 4 4 2
52 9 1 11 1 9 2 11 7 0 0 9 9 1 3 0 13 2 9 1 12 1 12 12 1 9 13 2 9 1 0 9 1 0 13 2 0 9 1 0 9 13 4 7 11 9 1 0 13 1 9 13 2
24 9 1 9 9 13 14 11 1 11 11 1 9 1 9 1 13 9 13 4 10 9 1 13 2
17 15 9 1 0 9 13 4 9 9 1 9 1 9 1 1 13 2
15 11 1 11 11 11 1 9 9 1 0 13 1 9 13 2
24 10 3 9 9 7 9 1 1 10 9 9 2 9 13 2 15 9 1 9 1 9 0 13 2
15 9 1 11 1 9 13 1 9 13 7 9 1 9 13 2
18 11 1 13 16 10 9 1 9 13 15 1 11 11 0 13 4 4 2
24 9 1 15 9 1 9 1 1 13 13 15 15 9 1 9 13 2 15 12 9 0 13 4 2
12 15 12 9 1 0 13 1 9 1 0 13 2
19 9 1 9 1 9 13 4 4 2 15 1 12 1 9 13 4 4 4 2
9 15 13 16 12 9 14 0 13 2
11 10 9 1 12 11 1 12 9 13 4 2
12 9 1 9 1 9 1 12 0 9 13 4 2
23 11 1 10 9 1 9 13 16 11 1 11 9 1 3 9 7 15 9 1 9 13 4 2
19 15 13 16 15 9 7 9 1 1 0 9 2 9 13 1 9 13 4 2
13 15 13 16 10 9 0 13 15 15 1 9 13 2
20 9 1 0 9 1 9 1 9 1 15 9 1 9 9 1 0 13 1 13 2
10 0 9 11 1 9 1 0 14 13 2
15 15 13 13 16 9 9 1 9 13 1 9 13 4 4 2
20 9 1 11 1 9 11 11 1 13 16 11 1 11 9 1 9 13 4 4 2
28 9 1 11 11 1 9 0 13 16 11 11 1 9 13 1 9 13 4 2 15 9 1 15 9 1 13 4 2
13 15 13 16 0 9 15 13 16 9 9 15 13 2
15 15 1 11 1 13 16 9 1 10 9 1 9 13 4 2
17 9 1 9 1 1 12 9 3 10 9 1 9 1 9 0 13 2
10 15 1 11 1 3 9 1 9 13 2
26 15 0 9 15 13 16 11 9 1 0 9 1 1 0 13 4 4 2 15 9 12 9 1 1 13 2
28 9 1 9 1 13 1 9 1 0 0 13 4 9 1 15 10 9 3 1 12 2 12 14 10 9 13 4 2
39 11 11 11 11 1 2 11 11 2 9 1 9 1 13 1 3 0 12 9 1 10 9 1 9 1 13 1 1 11 15 9 1 9 13 1 9 1 13 2
32 15 10 9 0 9 1 9 0 14 13 4 15 9 1 9 2 10 9 1 13 1 9 13 15 9 1 0 9 13 4 4 2
28 9 1 9 9 13 1 1 11 11 11 11 1 0 11 11 1 10 9 1 0 9 9 1 11 9 13 4 2
12 10 9 0 9 1 9 9 1 13 4 4 2
22 15 1 14 10 9 10 9 1 1 11 1 9 1 9 1 14 13 4 4 4 4 2
29 7 9 1 9 13 16 9 11 1 9 10 11 11 11 11 1 1 15 1 10 12 12 9 9 9 1 9 13 2
18 0 9 11 1 13 1 3 14 0 9 1 9 2 9 0 14 13 2
24 11 11 11 11 9 11 11 11 1 1 11 11 11 1 1 15 10 9 1 10 9 13 4 2
26 9 11 2 11 1 0 9 1 12 12 7 0 9 1 12 12 9 1 10 9 1 9 1 13 4 2
27 9 1 9 9 13 16 9 11 1 10 9 1 1 0 12 9 9 1 14 12 9 9 14 13 4 4 2
26 15 11 11 11 1 1 0 12 9 1 10 12 12 9 1 13 1 1 12 12 9 9 13 4 4 2
11 15 1 10 12 12 12 9 1 9 13 2
20 0 0 9 1 12 12 12 1 9 1 1 12 12 9 9 13 1 9 13 2
23 7 11 11 11 1 13 1 3 15 10 12 12 12 9 9 13 12 12 9 9 13 4 2
10 16 9 1 3 1 10 9 13 4 2
12 7 9 1 15 1 1 9 9 0 14 13 2
19 15 1 11 1 9 10 12 9 1 13 14 13 15 9 9 3 10 13 2
26 15 11 11 2 11 11 2 11 2 11 11 2 11 2 11 2 11 2 11 2 11 7 11 11 13 2
25 7 0 0 9 1 1 0 12 12 9 13 1 1 15 1 0 9 15 9 14 14 13 4 4 2
14 9 1 0 9 1 3 10 9 1 9 0 14 13 2
31 9 1 12 0 9 1 0 9 13 11 11 11 2 11 2 1 1 13 1 1 9 9 9 1 9 1 9 13 4 4 2
18 10 9 1 2 9 9 2 1 9 1 1 9 9 0 13 4 4 2
30 11 11 11 11 1 9 1 1 9 9 1 9 0 9 13 1 9 13 7 9 1 9 1 9 1 3 1 9 13 2
25 9 11 11 11 1 9 1 0 9 1 12 9 1 13 4 9 9 1 9 1 9 13 4 4 2
13 9 11 11 7 9 11 11 11 9 1 9 13 2
18 9 1 12 9 1 0 9 13 1 9 1 1 1 9 0 13 4 2
27 11 11 2 11 1 0 11 11 11 11 1 12 0 9 1 0 9 13 11 1 1 13 1 9 13 4 2
24 10 9 1 9 1 1 11 1 11 11 1 9 11 11 11 1 9 1 9 9 0 13 4 2
10 9 1 10 9 15 9 13 4 4 2
18 9 1 13 4 16 10 9 0 9 1 9 1 1 1 10 3 13 2
18 15 11 1 1 13 4 1 0 11 1 9 1 13 9 0 13 4 2
31 0 9 11 1 10 13 4 9 1 1 13 9 1 9 1 13 4 16 15 11 11 1 9 1 9 1 9 9 0 13 2
16 11 11 11 11 11 1 11 9 1 9 9 9 1 0 13 2
15 15 1 14 12 0 9 1 11 7 11 1 9 13 4 2
30 7 9 11 1 0 11 11 11 1 9 1 1 11 1 9 9 1 1 10 9 13 16 11 11 1 0 9 13 4 2
29 11 12 12 1 9 1 1 9 1 3 0 9 13 7 11 1 9 15 1 13 9 2 9 1 9 13 4 4 2
18 0 9 11 1 11 11 1 9 1 11 1 13 16 15 1 1 13 2
14 11 1 10 9 1 10 15 0 0 9 1 9 13 2
15 10 9 13 4 16 11 1 1 1 15 9 1 9 13 2
35 15 11 1 0 9 9 1 13 0 13 7 9 1 13 13 16 0 9 1 16 0 9 9 13 4 4 16 0 9 1 15 9 14 13 2
17 0 9 11 1 0 9 1 12 9 1 10 1 9 0 13 4 2
22 11 1 13 16 11 1 0 0 9 9 9 2 9 9 7 9 9 1 9 13 4 2
10 15 1 0 0 9 1 9 13 4 2
23 10 9 1 13 13 16 11 11 1 13 9 1 9 13 4 4 15 11 15 9 13 4 2
10 7 11 10 9 13 1 0 14 13 2
13 15 1 14 15 11 11 1 9 1 0 9 13 2
18 16 10 9 1 13 13 16 10 9 1 13 0 13 1 9 14 13 2
22 11 1 9 2 9 2 11 2 9 1 11 1 9 13 9 1 9 1 9 13 4 2
17 15 9 1 1 13 16 14 15 1 9 1 15 14 0 13 4 2
11 11 13 9 13 7 9 13 14 13 4 2
19 11 1 11 11 11 1 0 12 9 1 13 1 10 9 11 1 9 13 2
22 11 9 1 9 9 1 12 9 13 2 15 9 9 1 9 1 1 9 0 13 4 2
8 11 1 15 0 9 9 13 2
16 15 15 11 11 11 0 11 11 11 1 9 1 15 9 13 2
19 15 11 1 11 11 11 11 11 2 11 2 1 9 2 9 0 13 4 2
13 11 1 9 7 0 9 1 11 1 0 13 4 2
11 13 1 1 11 1 12 9 13 4 4 2
29 15 9 1 15 9 1 13 7 13 4 4 7 15 1 11 1 9 1 15 9 7 0 9 1 9 13 4 4 2
30 16 15 15 15 9 14 0 9 1 14 13 4 2 7 9 1 9 13 4 16 3 14 15 11 1 14 9 13 4 2
9 9 1 9 1 11 9 13 4 2
12 15 9 1 15 9 13 9 1 13 4 4 2
15 9 1 9 1 11 1 9 1 9 1 9 8 13 4 2
14 15 0 9 1 13 4 4 7 15 9 13 4 4 2
11 15 9 1 9 1 15 9 13 4 4 2
21 12 9 0 7 12 9 9 1 11 9 1 9 1 12 9 1 0 13 4 4 2
13 9 1 9 9 1 11 1 13 1 9 14 13 2
18 9 1 13 16 11 9 1 0 10 9 13 2 15 13 14 4 4 2
14 16 15 0 9 11 1 9 9 1 0 13 4 4 2
8 11 11 11 1 11 1 13 2
14 11 1 9 1 11 0 11 11 1 15 15 9 13 2
16 15 1 11 1 11 1 11 7 11 11 1 15 9 1 13 2
27 11 1 11 1 9 13 16 15 9 1 13 1 9 1 0 0 9 1 9 2 9 13 14 9 14 13 2
43 11 1 11 11 11 11 11 1 1 1 0 11 1 13 4 16 11 9 9 9 1 0 9 1 0 13 7 12 9 1 13 13 1 9 1 11 1 9 1 9 13 4 2
28 11 1 11 9 1 1 11 1 11 11 11 11 7 11 1 11 11 11 1 10 9 1 9 2 9 13 4 2
27 9 2 9 1 11 1 9 13 4 16 11 10 9 1 0 9 1 9 2 9 1 1 14 15 9 13 2
26 11 1 13 16 11 3 14 14 10 9 13 4 4 4 16 9 9 1 10 9 1 13 9 13 4 2
18 11 1 13 16 15 13 4 16 11 1 15 9 1 0 13 4 4 2
20 11 1 13 16 11 11 11 1 13 1 11 1 10 9 11 1 13 13 4 2
10 10 9 1 1 10 9 9 13 4 2
20 15 1 11 11 1 9 13 4 16 11 0 9 1 1 0 9 0 13 4 2
17 15 1 14 11 0 9 1 0 9 2 9 1 1 14 9 13 2
28 11 1 11 1 10 9 1 9 13 4 15 13 4 16 0 9 1 9 1 11 14 15 9 1 9 14 13 2
43 9 2 9 2 9 7 9 1 12 0 9 1 0 0 9 11 11 11 9 11 9 9 1 9 11 11 1 11 7 11 9 1 0 9 1 9 1 1 9 1 13 4 2
11 15 12 9 1 9 1 1 9 13 4 2
17 9 1 9 1 1 11 7 15 9 1 9 1 9 1 13 4 2
24 11 11 1 11 1 9 11 11 1 9 1 15 9 13 7 9 13 11 11 13 1 9 13 2
15 11 11 1 3 15 9 9 2 9 2 11 11 1 13 2
19 11 1 11 9 1 9 11 11 1 3 9 13 11 11 13 1 9 13 2
11 10 14 9 1 10 9 11 11 13 4 2
27 10 3 9 13 1 11 9 1 9 9 1 0 9 1 9 11 11 14 15 9 1 1 11 11 13 4 2
20 11 1 1 9 14 12 12 9 9 1 12 9 1 11 1 9 1 13 4 2
12 11 1 9 1 9 13 9 9 3 13 4 2
19 11 1 9 13 9 1 1 13 4 11 11 1 9 2 9 1 9 13 2
27 9 1 13 14 11 1 9 11 7 11 1 3 13 9 13 4 2 7 11 1 9 9 1 9 13 4 2
20 9 1 9 1 14 9 13 2 15 11 0 13 9 1 9 1 1 13 4 2
13 9 9 11 11 7 11 11 1 3 15 13 4 2
20 11 11 1 9 1 12 9 1 9 7 9 1 12 9 1 0 9 0 13 2
32 11 1 9 11 11 1 9 1 11 1 11 11 2 11 2 11 2 11 7 11 1 1 9 0 13 9 9 13 4 4 4 2
23 15 9 13 1 9 1 15 12 0 9 1 9 13 2 15 9 1 1 15 9 13 4 2
21 9 1 11 9 9 1 1 11 11 7 15 9 11 1 9 1 9 1 13 4 2
11 15 1 10 12 12 9 1 9 0 13 2
24 11 11 11 2 11 2 9 11 11 1 9 1 13 13 4 9 0 13 9 14 13 4 4 2
29 15 9 1 11 1 13 16 15 11 1 11 11 1 0 9 1 15 15 13 1 1 3 14 11 11 1 9 13 2
42 11 11 1 12 0 9 11 11 7 15 0 9 11 11 1 9 1 13 16 11 1 11 11 1 15 11 11 0 9 1 0 9 1 13 4 1 1 15 11 11 13 2
34 15 13 16 11 11 1 0 9 1 0 9 13 4 4 4 2 15 1 1 15 15 15 13 4 7 11 1 9 1 13 1 0 13 2
19 0 11 11 1 0 13 4 12 0 9 1 9 1 11 1 9 13 4 2
8 10 9 11 1 9 1 13 2
21 9 9 1 13 16 11 11 1 9 1 0 13 4 0 9 1 15 10 9 13 2
22 9 9 1 13 16 0 13 4 9 1 0 11 1 0 9 1 9 13 4 4 4 2
31 9 1 13 16 9 1 12 9 1 9 13 4 2 15 1 12 1 11 1 11 11 1 0 11 9 1 9 13 4 4 2
16 0 0 9 1 12 1 12 9 1 9 1 0 13 4 4 2
12 15 11 11 1 0 11 1 0 13 4 4 2
26 11 1 0 0 9 7 9 9 1 9 1 1 11 1 0 9 1 0 9 3 0 9 14 0 13 2
22 9 1 0 9 1 9 13 1 1 9 1 9 13 4 7 9 9 1 9 13 4 2
39 0 9 1 1 11 1 0 9 7 15 1 0 9 11 1 13 4 4 9 1 1 1 9 1 11 1 11 9 2 11 7 15 13 9 1 0 9 13 2
10 10 3 9 1 9 9 1 9 13 2
12 10 9 1 11 1 12 9 14 0 13 4 2
17 0 9 1 11 7 11 9 1 12 0 9 1 12 9 13 4 2
16 11 11 9 1 11 1 9 2 9 1 1 9 1 13 4 2
15 9 1 9 1 12 9 9 9 7 12 11 0 13 4 2
26 12 0 9 1 11 9 11 9 1 11 9 1 0 13 4 12 9 1 9 1 11 9 0 13 4 2
12 9 1 9 1 13 1 3 9 13 4 4 2
22 12 0 9 1 11 1 11 1 9 1 1 9 1 11 11 1 12 0 9 13 4 2
13 10 9 1 9 1 12 9 9 14 0 13 4 2
43 0 11 11 7 11 1 11 9 11 11 11 1 11 1 15 9 7 11 1 9 11 11 1 9 9 1 0 13 1 9 13 1 9 1 12 0 9 1 1 9 13 4 2
19 11 10 9 0 9 1 0 0 9 0 13 1 3 1 0 13 4 4 2
33 11 1 11 1 9 1 9 2 9 9 11 11 11 1 1 9 13 4 2 15 1 15 12 9 1 0 9 1 13 4 4 4 2
25 15 1 2 9 1 11 1 9 11 11 11 7 11 11 1 11 1 9 13 1 9 0 13 4 2
32 11 1 9 1 15 9 0 14 13 1 1 1 9 13 1 14 9 0 13 4 2 7 9 1 9 9 13 1 9 13 4 2
11 15 13 16 9 15 1 3 1 9 13 2
20 15 1 2 11 11 11 1 11 1 11 11 1 0 9 9 0 13 4 4 2
23 11 1 9 11 1 11 11 1 9 7 11 1 0 0 9 1 1 9 9 13 4 4 2
23 0 9 1 13 16 10 9 12 9 0 9 9 1 9 1 13 1 1 13 4 4 4 2
53 11 11 2 11 1 12 9 1 13 16 0 9 1 9 1 9 11 11 7 11 11 1 0 9 9 11 11 11 1 9 1 11 11 11 11 11 2 11 2 11 2 1 12 0 9 1 9 2 9 13 4 4 2
19 11 2 11 1 9 1 9 0 9 11 11 11 7 11 11 13 4 4 2
20 11 1 11 2 11 1 9 1 1 9 9 1 1 1 9 2 9 13 4 2
22 15 1 15 1 12 9 1 1 10 14 10 12 9 1 9 2 9 0 13 4 4 2
10 0 9 14 10 9 1 12 9 13 2
33 11 1 12 0 9 1 11 11 1 9 1 11 11 1 9 1 9 13 16 12 9 1 1 1 10 9 3 3 0 13 4 4 2
23 0 13 16 9 7 11 2 11 1 1 1 9 9 9 1 9 11 1 0 13 4 4 2
22 10 9 1 9 1 0 9 11 2 11 1 9 9 1 9 13 1 9 0 13 13 2
35 9 9 11 11 11 1 9 9 11 11 1 11 7 11 9 9 1 9 1 9 1 9 1 1 0 0 0 9 1 9 13 1 13 4 2
25 0 9 1 11 1 10 9 13 4 13 16 12 9 1 9 9 1 14 11 1 9 13 4 4 2
36 0 13 16 9 9 1 9 1 9 1 9 1 1 9 2 9 9 1 9 0 13 1 3 0 9 9 9 1 9 1 9 0 13 4 4 2
25 10 9 1 0 9 1 11 11 2 11 11 7 11 9 1 9 7 11 11 1 9 9 0 13 2
35 10 9 11 11 11 11 1 9 1 9 1 9 1 9 1 0 9 1 1 0 9 1 1 1 7 9 13 1 15 9 13 1 9 13 2
22 12 9 9 1 9 1 1 10 9 11 7 11 1 9 1 12 9 1 12 9 13 2
21 9 1 12 9 11 11 11 1 1 12 0 9 0 13 12 9 9 1 9 13 2
51 11 1 9 1 9 13 14 11 1 11 1 13 16 9 9 9 1 9 13 7 15 0 9 1 9 1 1 3 9 13 1 0 13 2 16 16 9 14 1 11 1 15 9 1 0 9 1 13 4 4 2
26 11 11 11 11 11 7 0 11 9 11 11 1 15 13 16 0 0 9 1 9 9 9 1 9 13 2
43 11 11 9 9 1 11 11 9 11 11 1 11 1 9 13 1 9 1 1 1 11 1 13 16 15 9 10 9 1 1 14 13 2 7 15 3 15 9 11 1 13 4 2
44 9 1 9 1 1 0 9 9 1 9 2 9 13 1 11 1 9 1 1 1 0 9 1 13 16 15 11 14 13 2 15 0 9 0 9 1 10 9 1 0 13 4 4 2
24 11 11 11 1 9 9 1 11 1 0 9 1 1 11 2 11 1 9 1 9 13 4 4 2
16 11 11 1 9 2 11 2 1 0 9 1 1 13 4 4 2
22 9 1 13 4 4 16 14 15 9 7 9 1 9 1 9 1 9 13 4 4 4 2
23 9 1 9 9 1 9 13 7 0 9 13 1 9 1 11 1 10 9 1 9 13 4 2
22 0 9 1 1 11 11 11 1 9 2 11 11 11 11 11 11 2 1 13 4 4 2
25 0 9 1 1 11 11 1 9 2 11 11 11 11 2 11 11 11 11 11 2 1 13 4 4 2
15 9 1 9 1 1 10 9 15 9 1 0 14 13 4 2
21 9 1 9 9 1 1 1 11 2 11 11 1 13 1 12 0 9 1 13 4 2
34 11 11 11 2 11 1 9 1 9 9 1 9 9 1 0 9 13 4 1 9 0 9 1 9 1 9 1 9 1 1 1 3 13 2
45 11 11 1 9 9 7 9 11 11 1 2 11 11 2 1 13 16 9 1 12 9 9 13 4 1 15 13 9 1 9 13 1 9 13 2 15 11 11 11 11 1 0 9 13 2
33 11 2 11 0 13 4 11 11 11 11 1 10 9 2 9 9 1 9 9 1 0 9 1 12 1 13 12 9 13 1 9 13 2
29 15 1 14 11 11 1 9 9 1 9 9 12 1 13 12 9 13 7 9 1 12 9 9 13 1 14 9 13 2
34 0 9 1 9 1 9 1 0 13 4 4 9 1 9 13 1 1 11 1 0 9 1 9 1 0 9 1 0 9 0 13 4 4 2
19 10 9 1 13 1 9 1 9 1 0 9 1 0 9 13 1 9 13 2
21 3 14 0 9 1 9 1 9 1 14 9 9 0 9 1 1 1 3 10 13 2
22 10 9 1 13 1 9 1 0 9 1 9 1 9 1 9 1 9 13 1 9 13 2
19 0 13 16 0 10 9 1 9 1 9 1 3 9 1 9 13 4 4 2
35 9 1 0 9 1 9 1 11 1 13 16 10 9 1 9 1 11 11 11 11 1 0 9 1 9 1 10 9 1 9 1 9 13 4 2
38 11 9 1 9 1 14 9 13 16 0 9 9 1 1 0 9 9 12 9 13 1 9 13 7 13 1 9 1 15 13 12 9 1 13 1 9 13 2
22 9 1 9 1 9 1 9 9 1 9 14 13 4 4 2 7 9 1 1 14 13 2
31 9 1 9 13 4 11 11 1 9 9 11 11 11 1 1 0 7 0 9 1 9 1 13 4 15 1 0 9 0 13 2
22 11 1 13 16 16 0 9 1 12 12 1 1 10 9 12 12 9 1 9 13 4 2
32 10 12 12 12 12 12 9 1 9 9 1 11 11 11 1 9 13 4 4 4 7 0 7 0 9 1 1 10 0 14 13 2
21 11 11 1 9 11 11 1 13 16 0 9 1 9 1 15 9 14 13 4 4 2
30 9 1 9 10 10 9 1 0 13 1 11 11 1 9 13 15 9 9 1 13 4 0 9 1 9 1 1 14 13 2
20 11 2 11 11 11 1 9 1 14 12 1 13 12 12 9 13 4 4 4 2
14 11 11 11 1 0 9 1 1 12 12 9 13 4 2
14 15 10 9 11 11 1 0 9 1 1 13 4 4 2
22 11 2 11 7 11 9 1 0 9 9 1 9 1 1 12 2 8 12 9 13 4 2
27 11 11 11 1 9 1 9 1 1 0 9 9 1 11 11 1 12 9 1 9 0 13 1 9 13 4 2
47 9 11 11 11 7 9 11 11 11 1 9 1 11 11 11 11 11 7 9 1 9 1 9 1 1 11 11 11 7 9 9 1 0 9 13 1 3 13 16 9 10 9 1 0 14 13 2
32 9 1 13 16 9 1 9 9 1 1 10 2 15 9 0 9 1 0 13 4 2 2 9 9 12 9 1 9 0 13 13 2
18 9 1 13 16 9 9 1 9 13 1 3 11 11 1 9 13 4 2
32 11 11 1 0 9 11 11 11 1 9 1 13 16 9 9 1 9 0 13 1 3 9 10 14 9 13 15 11 11 9 13 2
18 11 9 9 1 9 1 1 9 9 1 0 7 0 9 0 13 4 2
32 0 13 16 11 11 2 11 1 9 9 9 9 9 1 0 9 9 1 13 4 4 16 9 9 1 1 10 9 13 4 4 2
21 0 9 1 9 2 15 9 1 9 14 13 4 2 15 1 9 13 4 4 4 2
11 9 9 1 0 9 0 13 4 4 4 2
11 15 9 1 1 14 10 9 13 4 4 2
26 11 1 9 9 1 1 13 4 4 12 9 9 1 9 0 13 4 1 9 9 1 9 13 4 4 2
25 9 7 9 1 9 1 13 9 1 9 1 1 11 1 11 13 4 10 9 11 13 4 4 4 2
42 10 9 1 11 11 1 9 1 13 16 11 11 1 15 9 1 1 0 9 2 9 9 2 9 2 9 9 2 9 7 9 9 1 9 1 12 0 0 9 13 4 2
15 11 11 11 2 11 2 15 9 9 1 9 13 4 4 2
23 9 1 13 16 9 1 9 7 9 9 1 12 9 1 9 1 13 9 13 4 4 4 2
18 9 1 11 11 1 11 1 11 1 9 11 1 1 0 13 4 4 2
13 15 1 10 9 1 9 9 1 11 13 4 4 2
18 15 11 1 11 1 13 4 9 1 1 10 9 1 9 13 4 4 2
19 7 11 1 12 1 12 9 9 1 9 1 9 1 0 13 1 9 13 2
28 9 1 13 16 11 11 1 9 7 9 2 9 9 1 9 1 9 1 9 13 4 7 15 0 11 13 4 2
25 9 1 1 9 1 1 9 1 9 1 13 16 0 9 1 1 9 1 13 9 9 1 13 4 2
26 11 1 13 13 16 9 1 0 13 1 12 9 1 1 14 0 9 1 1 12 9 9 1 13 4 2
8 9 1 15 9 9 1 13 2
11 15 1 9 1 0 13 1 1 13 4 2
15 15 9 13 4 4 10 3 12 10 9 9 1 13 4 2
11 15 13 16 10 9 9 9 1 13 4 2
22 0 9 11 11 11 1 12 9 1 9 1 9 1 9 1 0 0 9 1 0 13 2
25 0 9 9 1 1 12 9 9 1 0 0 9 1 13 1 9 13 1 10 9 1 0 13 4 2
40 0 9 1 9 9 11 11 1 13 16 0 9 1 11 11 14 11 11 2 11 11 14 11 2 9 11 14 11 7 11 11 11 11 9 1 13 0 13 4 2
25 15 13 16 10 9 11 0 11 11 11 1 1 11 11 1 0 0 9 1 13 1 9 1 13 2
26 9 9 1 9 1 10 9 1 0 13 15 13 4 16 10 9 0 9 1 9 13 1 9 1 13 2
21 9 1 1 11 11 1 1 11 11 11 1 3 1 9 7 9 1 9 0 13 2
40 9 1 9 1 9 13 4 0 9 11 11 11 2 11 0 0 9 11 1 9 11 11 1 0 9 1 13 4 9 1 9 9 9 1 11 1 9 13 4 2
10 9 1 1 11 7 15 9 0 13 2
21 11 9 1 13 13 16 15 9 9 1 3 11 1 9 1 9 13 1 9 13 2
10 15 9 1 13 14 0 13 4 4 2
23 9 0 9 1 9 11 11 11 1 13 13 16 9 1 1 11 7 15 9 1 9 13 2
23 0 13 16 11 11 11 2 11 0 11 11 11 2 11 11 1 9 11 11 1 9 13 2
26 10 0 9 1 12 9 1 0 14 12 9 1 2 11 11 11 2 9 1 9 1 9 13 4 4 2
14 9 0 9 1 13 7 15 0 9 14 13 4 4 2
21 0 11 1 9 1 15 11 11 1 9 1 12 9 1 9 13 1 9 13 4 2
51 9 1 9 9 1 9 9 11 11 11 11 1 15 9 1 9 1 13 4 16 2 11 11 11 2 0 9 1 9 11 11 1 9 0 13 7 9 13 1 9 13 14 10 0 9 1 9 13 4 4 2
22 11 9 12 12 9 11 11 1 9 1 1 12 0 9 1 9 13 1 9 0 13 2
14 7 2 9 1 9 9 1 1 14 12 12 9 13 2
13 9 1 9 15 11 2 11 13 15 11 3 13 2
6 15 1 11 14 13 2
8 9 1 9 1 0 9 13 2
21 15 1 14 12 9 1 10 9 1 9 1 9 1 9 1 9 1 9 13 4 2
7 11 7 15 9 0 13 2
17 15 13 13 16 15 0 9 1 1 1 9 1 15 9 14 13 2
14 11 1 9 1 9 13 16 9 11 1 9 13 4 2
10 15 1 15 0 9 1 0 14 13 2
17 10 9 1 9 13 1 3 12 0 9 1 14 9 13 4 4 2
31 9 9 1 0 9 1 9 11 11 11 1 13 13 16 11 7 15 9 1 9 1 15 9 14 13 2 16 0 9 13 2
31 11 11 11 1 0 9 11 11 1 11 1 13 16 15 9 9 9 1 11 1 9 11 11 1 9 1 9 1 9 13 2
42 9 9 1 11 9 9 1 13 1 3 9 1 9 1 11 1 13 16 15 10 14 0 9 13 16 12 9 1 10 9 1 0 13 4 7 15 9 1 13 4 4 2
27 15 9 13 16 9 1 1 13 4 9 0 9 1 0 13 7 15 9 1 0 9 0 7 9 1 13 2
29 11 1 13 16 10 9 7 12 9 9 1 0 0 9 1 9 1 15 9 13 1 9 1 15 0 7 0 13 2
29 15 13 16 15 15 1 1 0 9 0 13 4 7 9 1 1 13 4 16 10 9 0 9 1 0 7 0 13 2
31 9 9 1 11 1 0 2 0 9 1 13 9 1 11 2 11 2 11 11 1 12 0 9 9 1 12 9 1 13 4 2
19 9 1 11 1 9 2 9 1 9 1 0 12 9 1 14 0 13 4 2
12 9 11 11 1 9 11 11 13 4 4 4 2
33 9 9 1 1 2 11 9 1 11 9 1 9 7 9 1 0 9 1 1 9 1 11 2 11 2 11 1 9 11 11 13 4 2
23 11 11 1 9 1 11 9 1 11 1 12 9 11 11 11 7 11 11 11 1 0 13 2
19 9 9 1 11 9 1 11 9 9 1 11 1 12 9 1 9 0 13 2
12 11 11 9 1 9 1 12 9 1 13 4 2
18 11 9 1 9 1 13 4 11 9 1 9 1 12 9 0 13 4 2
35 9 9 11 11 1 9 11 11 1 11 11 11 1 9 0 13 11 9 1 11 11 11 2 11 2 1 11 1 0 13 1 9 13 4 2
28 15 1 14 11 1 9 1 1 9 13 1 11 1 15 0 9 9 1 1 0 9 1 13 1 9 13 4 2
45 11 1 9 11 11 1 11 1 11 11 1 9 0 13 11 1 11 1 11 11 11 1 9 13 1 1 11 1 0 13 1 9 13 7 13 16 11 1 9 1 13 4 4 4 2
38 11 1 9 13 16 15 11 1 9 11 11 11 11 1 11 1 9 1 15 9 1 13 13 4 2 15 15 13 4 16 9 9 1 15 9 13 4 2
16 11 11 7 0 11 1 11 9 9 1 0 9 0 13 4 2
18 0 13 16 11 11 1 13 0 9 1 1 0 13 9 1 9 13 2
13 9 1 9 1 9 11 11 1 12 0 13 4 2
17 15 9 11 1 12 9 0 9 7 12 9 0 9 1 0 13 2
10 9 11 9 12 13 12 9 1 13 2
26 9 9 1 0 9 13 1 9 1 9 10 0 0 0 9 1 9 1 9 13 1 9 13 4 4 2
24 11 11 11 11 1 9 9 1 1 9 1 13 16 15 9 9 1 9 2 9 13 4 4 2
10 10 9 1 14 9 2 9 0 13 2
46 11 1 9 1 9 1 15 9 1 9 13 4 1 9 13 4 11 11 1 13 16 9 1 10 9 13 4 4 2 7 9 1 0 9 13 1 1 1 15 0 9 1 9 13 4 2
34 15 1 11 9 11 11 11 1 1 11 1 11 11 1 9 13 4 11 9 11 11 1 13 16 15 10 9 9 1 9 13 13 4 2
6 15 15 9 13 4 2
8 15 15 9 14 13 4 4 2
28 13 4 4 4 16 11 1 9 1 9 9 1 10 0 9 1 9 1 9 1 13 11 11 1 9 13 4 2
14 15 11 11 1 13 16 9 9 9 1 1 13 4 2
37 9 9 9 13 1 0 9 1 9 1 9 1 9 13 4 4 2 7 15 13 13 16 15 0 0 0 9 1 9 1 9 1 9 13 4 4 2
30 0 9 1 0 9 1 9 1 9 1 1 11 1 11 1 11 1 2 12 0 9 7 9 2 0 13 1 13 4 2
32 9 9 7 0 9 1 15 0 9 1 9 1 1 11 1 9 13 4 1 3 11 10 9 1 9 13 1 0 13 4 4 2
28 12 9 15 2 15 1 15 13 4 9 1 15 9 1 9 1 9 1 13 1 9 13 1 0 13 4 4 2
14 12 9 1 1 12 0 0 0 9 11 1 0 13 2
32 10 9 1 12 9 1 0 0 9 7 0 9 1 9 1 9 1 13 1 9 13 1 0 13 4 12 0 9 2 0 13 2
44 9 1 11 1 9 9 11 11 1 1 9 13 1 0 9 9 11 11 11 1 13 16 12 9 1 15 0 9 1 0 13 4 9 1 9 1 0 9 1 9 2 9 13 2
31 12 9 1 1 9 1 9 13 4 11 1 13 16 11 1 0 11 11 1 1 11 1 11 11 11 1 9 1 9 13 2
18 11 1 0 9 13 7 15 14 9 1 9 1 9 1 9 14 13 2
36 9 2 9 1 1 11 1 0 13 16 15 15 11 1 13 9 1 11 1 0 11 1 9 1 9 9 1 15 9 1 9 1 0 14 13 2
7 9 1 9 13 4 4 2
20 9 1 13 4 4 16 12 9 9 7 9 1 9 13 1 0 13 4 4 2
33 9 1 9 1 9 1 11 1 11 11 1 10 9 1 0 9 0 13 1 13 2 15 9 1 12 9 1 1 9 13 4 4 2
18 12 9 1 0 9 1 9 13 1 1 3 9 1 9 1 9 13 2
20 0 9 1 13 1 1 14 12 9 9 1 9 13 7 9 13 1 0 13 2
22 0 9 11 1 12 0 0 9 1 9 13 1 9 1 12 9 1 0 13 4 4 2
8 9 1 11 1 10 9 13 2
26 11 1 9 9 11 11 1 13 16 9 1 9 1 0 10 12 9 1 0 13 9 13 4 4 4 2
19 11 1 13 16 10 9 1 0 9 7 9 1 1 15 9 0 13 4 2
14 15 13 16 9 1 9 9 1 9 1 9 13 4 2
26 11 1 9 12 9 1 9 13 4 2 7 11 1 9 1 0 12 9 1 9 1 9 13 4 4 2
11 9 1 9 12 1 12 9 1 1 13 2
13 9 1 10 9 11 9 1 11 9 1 1 13 2
13 10 9 15 9 2 9 1 9 0 13 4 4 2
8 0 13 16 9 9 13 4 2
39 11 1 11 11 1 13 1 0 9 1 9 1 1 0 9 1 9 1 13 4 11 2 11 11 7 11 11 1 13 9 1 9 13 1 9 13 4 4 2
36 11 9 1 12 9 1 9 0 9 1 0 13 1 0 0 9 9 11 11 11 1 13 16 0 9 1 9 1 1 9 9 1 0 9 13 2
23 0 9 1 9 1 1 11 1 13 9 9 1 0 9 1 9 1 9 13 4 4 4 2
10 15 9 7 9 9 1 1 9 13 2
35 9 1 11 11 1 9 1 13 4 16 11 11 1 0 0 9 1 9 1 10 9 1 0 9 1 9 1 1 0 9 1 9 13 4 2
32 9 1 13 16 10 14 9 1 9 1 11 9 1 13 11 9 1 1 13 1 9 9 2 9 7 0 9 1 9 13 4 2
11 10 9 1 9 1 10 9 13 4 4 2
19 15 1 0 9 1 11 1 0 9 1 10 0 9 13 1 14 9 13 2
22 9 1 13 16 9 1 9 1 9 13 1 3 10 9 9 9 13 11 13 4 4 2
12 0 9 1 12 9 9 9 1 9 13 4 2
18 15 1 10 9 0 7 0 11 2 11 7 11 9 1 0 9 13 2
19 9 9 11 11 11 1 13 16 3 0 9 1 11 1 9 0 13 4 2
36 11 11 11 11 2 11 2 1 12 9 1 9 13 1 9 1 9 1 9 11 11 2 9 9 2 9 7 12 0 9 1 0 13 4 4 2
29 10 9 1 9 11 1 12 9 1 11 11 11 2 11 2 1 0 13 1 1 0 9 1 9 13 1 9 13 2
22 9 1 1 11 1 11 11 11 1 11 11 0 11 1 9 1 12 9 1 0 13 2
18 3 1 15 0 9 2 9 2 11 11 11 1 9 1 0 13 4 2
15 9 1 10 15 1 11 11 1 0 9 1 13 4 4 2
54 11 11 1 9 1 1 11 1 9 1 1 9 9 11 11 11 2 9 1 9 11 11 11 2 9 11 11 2 9 11 11 2 9 9 11 11 7 11 11 2 9 9 11 11 7 9 11 11 11 1 0 13 4 2
26 11 11 1 9 9 1 9 1 13 4 9 1 0 9 9 13 4 1 3 9 1 0 13 4 4 2
29 9 1 1 15 1 11 11 11 1 1 11 11 11 1 11 11 2 11 2 11 7 11 1 1 0 13 4 4 2
26 11 11 1 9 1 11 11 1 11 9 1 9 1 1 9 1 0 9 1 15 9 1 13 4 4 2
22 9 1 1 10 9 1 1 11 9 1 9 1 1 1 15 9 1 9 14 13 4 2
19 15 1 9 1 11 11 1 9 1 1 0 9 13 1 9 13 4 4 2
11 15 1 9 1 11 11 11 1 9 13 2
19 9 1 11 1 9 9 1 1 9 13 7 10 0 9 13 1 9 13 2
17 15 1 10 9 1 9 1 9 13 4 10 9 0 13 4 4 2
22 9 1 9 1 1 9 11 11 11 1 14 9 9 1 1 9 13 1 1 13 4 2
27 9 0 13 1 1 9 1 9 13 1 9 13 4 9 1 0 13 7 3 14 9 13 1 9 13 4 2
14 11 1 11 1 9 1 0 13 10 9 1 9 13 2
14 15 1 11 11 1 0 11 11 11 0 13 4 4 2
22 11 9 1 9 9 7 15 9 0 11 11 11 1 9 13 11 11 11 1 9 13 2
9 11 15 1 0 9 13 4 4 2
8 11 10 9 11 11 11 13 2
26 11 11 1 0 2 0 13 4 9 9 11 11 11 1 9 1 11 9 1 9 9 11 11 9 13 2
38 10 9 11 1 9 9 1 11 1 9 13 4 9 9 9 11 11 11 1 11 11 1 9 1 9 2 9 9 1 0 9 13 1 1 13 4 4 2
24 11 1 9 2 9 2 9 2 9 7 9 9 1 11 11 1 9 1 9 0 13 4 4 2
16 7 11 11 1 9 9 9 9 9 1 0 9 13 4 4 2
24 11 11 11 1 9 9 2 11 2 11 2 11 11 11 1 11 9 1 9 0 13 4 4 2
26 0 9 1 13 16 11 11 11 11 11 11 11 2 11 2 1 14 0 9 2 9 13 1 9 13 2
22 11 1 11 9 1 9 9 11 11 1 9 9 1 9 2 9 2 0 13 4 4 2
30 11 1 0 9 11 11 2 11 11 2 11 11 11 7 11 11 11 1 9 9 9 2 9 2 9 1 0 13 4 2
15 15 9 1 13 4 0 9 1 9 1 1 1 0 13 2
26 9 9 1 0 9 1 1 0 7 0 11 1 9 11 9 1 9 9 9 1 9 1 13 4 4 2
14 7 0 12 0 9 1 15 1 10 9 14 13 4 2
32 16 9 1 9 13 4 16 0 0 9 1 10 9 1 0 13 1 14 15 9 1 9 1 10 9 1 9 13 4 4 4 2
15 0 9 1 9 11 11 1 11 1 12 9 1 9 13 2
26 15 13 16 11 0 9 1 13 1 12 1 12 1 9 1 11 9 1 9 1 15 9 14 13 4 2
24 7 15 10 9 13 1 1 12 0 9 11 7 11 1 9 1 15 1 9 14 13 4 4 2
15 10 9 1 9 1 1 1 3 15 9 14 13 4 4 2
12 12 1 9 1 11 9 0 0 0 9 13 2
13 10 9 11 1 9 1 12 0 9 1 13 4 2
12 3 11 9 1 12 9 11 11 1 13 4 2
10 15 0 9 13 15 9 0 13 4 2
18 10 9 11 7 11 11 9 1 9 1 14 9 2 9 13 4 4 2
25 7 11 11 1 10 9 14 12 13 7 15 11 11 1 12 9 1 9 1 11 9 1 13 4 2
26 11 9 11 11 1 13 16 15 1 9 1 10 9 1 1 10 9 1 9 1 9 0 13 4 4 2
9 15 9 1 12 9 0 13 4 2
34 15 13 4 11 11 11 1 11 11 9 1 0 9 1 13 9 1 1 0 11 11 11 11 11 1 15 12 9 1 15 0 13 4 2
25 15 11 1 0 9 11 11 11 7 11 11 1 9 1 9 11 9 11 11 1 9 1 13 4 2
35 15 13 13 16 11 11 1 0 9 1 9 14 12 9 1 9 1 13 7 10 12 9 1 9 1 1 11 11 1 15 9 0 13 4 2
15 15 13 16 15 14 0 9 1 10 9 15 13 14 13 2
40 11 1 11 7 11 1 9 0 9 11 11 1 14 13 2 15 11 11 1 9 1 11 11 1 0 9 2 9 1 11 1 9 1 13 1 0 9 13 4 2
5 11 15 14 13 2
9 7 15 9 13 1 0 14 13 2
33 11 7 11 1 1 11 1 11 1 1 9 9 9 1 9 1 9 1 1 11 11 1 9 12 9 1 9 1 15 13 4 4 2
19 11 9 9 11 2 11 11 1 1 9 9 1 9 1 9 2 9 13 2
24 9 1 13 13 16 12 9 1 9 9 9 9 9 13 1 9 7 9 1 9 1 9 13 2
21 0 13 16 11 7 11 1 11 1 1 9 9 9 1 12 9 0 13 4 4 2
14 9 9 1 9 1 1 0 9 1 9 13 4 4 2
13 7 0 9 1 9 2 9 1 9 13 4 4 2
26 9 1 9 1 9 9 1 0 9 1 1 11 1 11 11 1 11 11 1 1 12 0 0 9 13 2
18 10 9 11 11 1 9 12 9 9 13 0 9 9 12 9 11 13 2
18 9 1 10 9 11 11 2 11 2 11 2 11 7 11 9 1 13 2
24 9 1 10 9 11 1 11 11 11 1 9 12 9 13 4 0 9 9 12 9 11 11 13 2
16 11 1 11 11 11 11 1 11 1 11 11 11 1 9 13 2
28 11 1 11 1 11 9 13 1 1 9 13 7 9 13 16 0 9 1 0 13 1 1 13 4 9 0 13 2
28 11 1 13 16 9 1 9 9 1 9 1 9 1 0 13 4 16 15 15 2 15 1 0 9 13 13 4 2
13 9 9 1 9 1 14 12 9 1 9 0 13 2
12 11 1 11 11 11 1 14 11 1 9 13 2
22 11 1 11 1 9 0 13 7 0 9 1 1 11 1 11 1 9 1 14 9 13 2
31 9 9 9 9 9 11 11 1 9 7 9 1 9 1 9 1 11 11 2 11 2 9 11 11 1 11 1 9 13 4 2
23 11 11 11 1 11 9 1 11 1 12 9 7 9 1 9 1 12 0 9 1 9 13 2
11 11 1 9 14 9 2 9 0 13 4 2
15 9 9 7 9 1 1 15 13 11 9 9 1 0 13 2
25 11 2 11 1 0 11 11 11 11 1 13 4 16 9 1 9 0 13 15 1 3 0 9 13 2
21 10 9 9 1 11 11 11 11 1 13 4 4 4 2 15 3 11 1 9 13 2
15 15 9 13 16 10 9 1 3 13 9 1 9 0 13 2
26 11 11 11 11 11 11 11 1 11 1 9 1 0 9 2 9 1 13 16 15 0 9 13 13 4 2
12 7 15 1 0 9 1 15 9 14 13 4 2
14 1 15 2 9 12 9 9 1 9 9 14 13 4 2
9 15 9 1 9 1 9 0 13 2
26 11 1 10 9 1 14 10 9 13 16 2 9 9 2 9 1 11 11 11 1 13 13 4 4 4 2
25 15 13 16 2 9 9 2 9 9 1 11 1 9 13 7 9 9 9 1 15 9 13 4 4 2
28 11 1 13 13 16 9 1 9 0 13 15 1 0 9 13 7 15 1 15 0 7 0 0 9 1 9 13 2
10 0 11 11 1 15 0 9 14 13 2
27 15 13 13 16 11 1 10 9 1 1 10 9 0 13 7 11 1 0 13 1 1 15 14 0 9 13 2
21 11 10 9 1 14 10 0 13 16 9 9 1 11 1 3 10 13 13 4 4 2
9 7 9 1 11 1 0 9 13 2
13 9 9 1 11 1 12 9 1 9 0 13 4 2
17 15 1 9 1 12 1 12 9 11 1 11 1 1 13 4 4 2
30 11 1 9 13 1 3 11 1 13 1 9 1 1 1 9 13 4 1 11 1 13 16 11 1 9 15 13 4 4 2
10 9 1 9 15 14 9 13 4 4 2
8 0 9 14 9 13 4 4 2
10 15 2 11 1 15 15 9 14 13 2
24 11 11 11 1 1 1 9 13 4 1 15 13 16 15 15 1 1 15 9 14 13 4 4 2
25 15 15 9 1 1 1 9 13 4 1 11 1 13 16 15 1 1 15 14 0 14 13 4 4 2
16 16 2 0 9 11 1 9 9 1 12 9 0 13 4 4 2
21 9 1 9 1 13 9 9 7 11 11 12 9 3 0 2 8 9 13 4 4 2
20 9 9 1 13 13 16 10 9 9 9 1 1 9 1 9 12 12 9 13 2
30 7 11 11 1 1 10 9 9 1 9 12 12 9 13 1 9 13 2 15 0 9 1 1 1 14 12 9 10 13 2
19 7 9 1 13 13 16 10 9 9 1 9 0 9 1 1 1 10 13 2
17 9 9 7 11 11 1 9 9 1 1 0 9 1 0 13 4 2
35 9 9 7 9 1 3 0 9 11 11 11 11 11 11 11 16 11 1 13 13 16 10 9 9 1 9 10 13 1 9 13 4 4 4 2
22 9 9 9 13 4 16 10 9 9 1 1 9 1 9 0 9 1 1 1 10 13 2
13 9 1 1 10 9 9 9 14 12 12 9 13 2
13 15 0 9 1 9 1 14 12 12 9 10 13 2
11 0 9 9 1 9 12 12 9 13 4 2
29 11 11 9 9 1 10 9 1 9 14 13 4 7 15 1 10 9 9 9 1 14 12 9 1 9 13 4 4 2
16 10 9 11 7 11 1 10 9 1 9 9 9 1 13 4 2
11 0 9 12 12 9 9 1 9 13 4 2
19 11 1 13 13 16 10 9 1 9 1 9 9 1 9 1 14 13 4 2
21 15 13 13 16 15 1 10 9 0 9 1 13 4 15 0 9 1 0 13 4 2
30 12 9 1 10 9 1 13 4 11 11 11 1 9 1 9 1 0 13 1 1 9 1 0 9 1 9 0 13 4 2
22 9 1 9 1 10 9 0 13 4 4 7 15 9 1 9 1 1 13 4 4 4 2
27 3 0 9 1 9 1 9 1 1 0 9 7 9 1 11 11 11 11 1 14 9 1 9 13 4 4 2
11 0 9 1 0 13 4 1 0 9 13 2
38 9 9 9 9 9 11 11 1 13 16 11 11 11 11 1 9 1 12 9 9 1 0 13 4 4 4 7 15 9 1 0 9 1 0 13 4 4 2
15 9 1 15 9 1 9 13 4 15 0 13 4 4 4 2
12 11 11 1 13 16 15 15 9 1 1 13 2
20 11 1 13 16 10 9 9 1 15 9 1 8 13 1 0 9 13 4 4 2
22 9 9 9 9 9 1 1 9 1 9 1 11 11 11 11 1 14 9 13 4 4 2
30 11 11 1 13 16 0 9 1 1 15 9 7 9 1 9 13 1 9 1 15 9 7 9 1 0 14 13 4 4 2
12 11 1 13 16 11 11 1 14 10 9 13 2
20 15 1 9 9 7 9 1 9 1 1 9 13 1 9 1 0 13 4 4 2
17 16 10 9 1 9 1 9 9 1 0 13 4 16 15 14 13 2
10 16 15 9 7 9 1 9 14 13 2
22 15 15 14 0 13 4 7 15 9 2 9 7 15 0 9 3 10 9 1 13 4 2
11 15 9 1 9 14 9 7 9 14 13 2
23 11 11 1 13 16 15 9 7 9 2 9 1 9 13 1 1 1 0 9 1 9 13 2
19 9 1 9 1 9 1 0 13 4 9 9 1 9 1 9 13 4 4 2
32 9 1 9 1 0 9 13 4 16 2 9 1 9 1 1 0 9 14 9 1 11 1 1 9 1 1 13 1 9 13 4 2
44 9 1 1 15 9 1 0 9 9 1 0 9 1 13 4 0 9 1 0 9 1 13 4 4 4 2 14 10 9 9 1 0 9 1 9 15 0 0 9 1 10 14 13 2
28 11 1 0 9 2 9 2 11 11 13 4 16 9 1 10 9 1 1 9 1 13 1 9 13 4 4 4 2
25 10 9 9 1 11 11 11 2 11 2 7 11 11 1 9 9 1 14 9 9 1 0 13 4 2
27 9 1 9 9 11 11 11 13 4 16 9 1 9 1 10 9 9 1 0 9 1 0 13 4 4 4 2
10 9 1 11 9 1 12 9 9 13 2
14 11 1 11 7 11 9 9 14 9 1 1 0 13 2
11 15 9 13 1 3 9 1 0 9 13 2
23 9 1 9 1 1 9 14 1 12 9 1 9 9 0 13 1 1 0 13 4 4 4 2
11 9 9 1 0 9 0 0 9 1 13 2
25 0 9 9 11 11 1 13 0 11 11 1 9 9 1 9 13 14 9 1 9 9 13 4 4 2
23 0 9 1 1 9 1 0 9 13 4 4 16 15 9 1 1 0 9 1 1 0 13 2
22 11 2 11 7 11 1 13 1 11 2 11 7 11 1 9 7 9 9 14 13 4 2
37 9 1 12 9 9 0 13 1 3 11 1 9 12 13 12 9 1 0 9 1 1 9 2 9 1 1 11 9 1 9 9 1 9 13 4 4 2
22 15 0 9 1 9 1 1 9 12 9 1 14 9 1 0 9 13 9 13 4 4 2
34 0 9 11 11 11 11 1 9 9 1 1 9 9 13 9 1 9 11 11 1 13 4 9 9 1 13 15 3 1 9 1 13 4 2
29 10 9 1 1 11 14 1 9 1 9 9 1 13 11 11 13 4 7 11 14 1 9 1 9 9 1 13 4 2
14 15 1 9 11 11 1 10 9 1 0 9 0 13 2
20 9 9 1 3 9 9 9 1 0 9 11 1 11 9 1 15 9 1 13 2
16 3 9 1 11 11 11 1 9 9 1 9 1 0 13 4 2
19 7 0 9 1 1 9 1 9 9 1 10 9 14 0 9 1 9 13 2
29 0 3 11 9 7 11 11 11 1 9 1 11 9 1 9 11 11 1 9 1 9 1 9 1 9 15 9 13 2
14 0 9 1 14 1 11 1 9 13 15 9 13 4 2
8 9 1 9 1 1 13 9 2
26 3 10 9 1 9 1 13 4 16 10 9 1 9 1 15 9 1 9 1 1 9 0 13 4 4 2
39 9 1 10 9 1 10 14 9 1 11 1 9 1 0 9 1 13 12 9 1 9 13 16 12 9 1 15 9 1 13 4 7 15 9 1 14 13 4 2
23 16 11 1 13 16 15 3 9 1 14 13 2 16 9 1 9 1 1 9 1 13 4 2
9 10 9 11 1 9 12 9 13 2
5 0 13 9 11 2
30 11 9 1 12 2 12 9 1 9 1 9 15 0 13 16 9 11 0 13 7 9 1 15 13 1 1 9 14 13 2
18 9 14 1 14 12 12 1 10 9 9 11 1 9 1 1 13 4 2
13 15 14 9 14 10 9 1 0 9 13 4 4 2
13 11 1 0 9 1 9 1 9 13 1 9 13 2
25 16 9 1 11 1 11 1 10 9 1 13 9 1 1 10 9 1 11 9 1 9 14 9 13 2
18 3 1 11 9 1 9 1 1 11 9 1 9 1 9 0 13 4 2
17 10 9 1 11 9 1 0 13 9 1 10 9 1 13 4 4 2
12 11 9 1 1 9 1 0 9 9 13 4 2
54 16 11 9 1 9 9 2 9 9 2 11 11 1 13 16 10 9 1 9 2 9 7 9 1 12 9 3 13 9 1 9 13 1 9 1 1 11 11 1 9 2 9 1 1 9 9 10 14 10 13 1 9 13 2
21 11 9 1 14 11 11 1 9 2 9 1 9 13 1 1 0 13 4 4 4 2
17 9 1 13 13 16 11 1 9 15 1 9 1 9 14 0 13 2
15 9 1 1 13 10 9 15 10 9 1 0 14 13 4 2
28 0 9 11 1 11 11 11 2 11 2 1 9 11 11 2 11 11 7 11 11 1 9 1 10 9 13 4 2
11 10 9 15 1 12 1 9 1 0 13 2
30 9 1 1 11 11 1 11 9 11 2 11 1 9 1 0 14 9 13 4 2 15 10 9 0 9 9 1 9 13 2
23 11 1 9 1 3 0 9 9 1 9 14 13 4 2 15 9 14 12 9 13 4 4 2
16 15 1 0 9 1 9 1 9 2 9 1 9 2 13 4 2
21 10 9 1 10 9 9 1 1 9 13 1 1 9 0 13 1 9 13 4 4 2
10 15 9 14 12 12 9 13 4 4 2
19 10 9 1 11 11 7 0 10 9 1 0 9 1 9 1 9 13 4 2
22 10 9 9 1 9 1 1 7 0 9 1 13 7 15 1 10 9 1 9 13 4 2
5 10 9 0 13 2
25 15 0 13 4 16 10 9 1 15 9 9 1 13 7 15 0 13 1 1 9 1 9 0 13 2
11 15 9 1 9 1 9 14 13 4 4 2
15 9 1 10 9 1 10 0 9 1 9 14 9 13 4 2
24 11 13 4 16 10 9 1 9 1 9 2 9 7 0 9 1 0 9 7 9 14 13 4 2
9 15 9 12 12 9 13 4 4 2
6 9 1 9 0 13 2
23 9 13 16 10 9 1 10 3 0 9 0 13 1 1 9 13 1 9 13 4 4 4 2
34 10 9 1 9 2 9 1 9 0 13 1 1 9 1 10 9 14 9 13 4 2 15 10 3 0 13 9 1 9 1 9 13 4 2
35 11 1 13 9 1 1 1 15 13 16 15 1 9 1 1 1 12 9 1 9 13 4 2 15 10 3 1 0 9 9 9 1 9 13 2
31 11 1 1 9 9 13 1 9 13 4 11 1 13 16 16 0 9 1 9 13 4 16 10 14 10 9 0 13 4 4 2
18 11 11 1 9 11 1 9 9 0 9 1 13 9 9 1 13 4 2
17 15 9 9 1 1 9 1 9 0 9 2 9 2 1 13 4 2
8 12 9 1 9 1 9 13 2
10 9 1 11 9 3 0 13 4 4 2
24 11 1 11 7 11 9 1 12 9 7 15 1 12 9 0 9 9 13 11 1 9 13 4 2
6 9 0 9 1 13 2
21 11 11 11 11 1 9 11 11 1 1 0 9 12 12 9 1 9 1 9 13 2
8 15 12 12 9 1 9 13 2
19 9 11 11 1 13 16 9 9 1 11 11 1 9 9 0 13 4 4 2
32 10 9 1 0 9 11 11 2 9 9 11 11 2 11 11 2 11 11 2 11 11 2 11 11 7 9 11 11 14 0 13 2
11 10 9 11 1 12 9 0 9 0 13 2
18 11 7 11 9 11 11 14 1 9 9 9 1 1 9 13 4 4 2
35 12 9 1 0 9 1 9 11 11 14 1 0 9 13 7 12 1 11 1 9 11 14 1 9 1 1 11 9 1 1 15 9 13 4 2
12 9 12 9 1 9 1 9 14 0 13 4 2
17 11 1 11 11 11 11 7 9 9 11 11 10 9 1 0 13 2
21 9 13 16 9 1 11 11 11 11 1 9 14 1 9 1 9 9 0 13 4 2
9 9 13 1 9 12 1 9 13 2
15 15 1 15 0 9 1 3 9 1 9 1 9 13 4 2
29 11 1 9 13 9 11 14 1 9 1 0 13 7 11 1 9 1 9 7 0 0 9 1 9 14 1 9 13 2
18 9 1 13 16 11 1 9 12 9 1 14 12 9 11 1 0 13 2
20 10 9 9 1 1 11 11 1 0 11 9 1 9 1 9 14 13 4 4 2
26 3 11 1 9 1 13 16 9 1 9 1 1 9 1 0 9 1 11 1 9 1 0 13 4 4 2
19 0 9 1 9 13 4 4 4 7 10 9 1 3 9 13 4 4 4 2
28 11 1 10 0 9 1 1 0 13 1 1 1 12 9 9 14 13 4 7 9 1 0 9 1 9 0 13 2
19 0 9 1 1 12 9 1 9 1 13 4 9 1 9 0 13 4 4 2
24 3 11 1 0 9 1 1 11 1 11 0 9 9 1 9 1 3 13 1 9 14 13 4 2
23 11 7 11 9 9 1 9 1 9 1 13 4 0 9 1 3 13 1 9 14 13 4 2
16 15 1 12 12 9 1 11 1 0 9 9 1 9 13 4 2
20 9 1 9 1 9 1 13 0 0 11 11 1 13 1 1 9 1 9 13 2
15 11 1 3 0 9 14 9 12 1 12 9 1 13 4 2
10 15 9 1 9 1 9 10 13 4 2
15 11 1 9 1 1 1 10 9 1 14 9 14 13 4 2
12 15 1 11 1 0 9 1 9 1 9 13 2
20 9 9 1 13 13 16 0 12 9 1 9 0 13 7 9 1 9 0 13 2
20 11 9 12 9 1 11 9 1 10 9 1 9 1 0 9 13 4 13 4 2
30 3 2 3 9 13 7 11 1 13 9 1 9 1 9 7 9 1 9 13 16 13 9 0 2 0 9 1 13 4 2
8 15 9 14 9 1 13 4 2
18 16 0 9 7 9 1 1 9 13 7 0 9 1 15 0 13 4 2
16 9 1 1 15 15 9 1 9 1 13 15 9 1 3 13 2
28 9 1 9 1 1 11 1 13 7 9 13 15 0 9 14 13 2 7 9 1 1 10 9 3 9 13 4 2
14 9 1 13 1 1 10 9 1 9 1 9 13 4 2
20 9 1 9 14 9 1 10 9 1 9 13 4 15 3 10 9 13 4 4 2
17 11 1 12 9 0 9 11 1 13 12 9 1 10 13 4 4 2
32 9 15 11 9 1 13 4 9 15 2 15 9 13 9 1 13 15 15 11 1 9 13 13 1 1 10 9 1 9 13 4 2
14 9 1 9 1 13 4 15 15 9 7 9 3 13 2
14 9 1 9 11 1 9 1 1 12 12 9 10 13 2
10 11 9 1 9 12 1 12 9 13 2
8 9 1 9 1 0 9 13 2
18 9 9 1 11 7 11 1 9 1 1 14 0 13 1 13 4 4 2
17 11 1 11 0 11 1 9 7 9 1 1 9 13 4 4 4 2
20 11 11 9 1 1 0 9 1 9 13 4 11 1 14 9 13 4 4 4 2
21 9 9 11 11 1 13 16 9 7 0 9 1 1 9 1 0 9 13 4 4 2
23 11 11 11 11 1 10 0 0 9 1 9 13 4 4 4 7 9 1 9 13 4 4 2
24 9 1 9 9 11 11 1 13 16 10 9 7 9 9 9 1 9 13 1 9 13 4 4 2
28 11 1 11 11 1 11 11 11 1 11 1 13 9 1 9 13 4 13 16 0 9 1 9 13 4 4 4 2
14 11 1 11 11 11 11 1 9 9 0 13 4 4 2
15 11 1 9 9 11 11 1 13 16 9 1 9 0 13 2
14 7 9 1 1 1 9 9 1 0 13 4 4 4 2
18 9 1 1 9 0 13 1 3 9 1 0 9 1 9 1 13 4 2
26 11 9 1 11 1 9 11 1 9 1 1 9 9 13 11 14 1 9 1 9 9 1 13 4 4 2
18 9 11 1 0 9 1 13 4 9 9 1 9 1 9 1 13 4 2
15 15 1 9 1 1 9 11 11 1 9 0 13 4 4 2
18 9 0 13 1 9 1 14 12 12 9 1 9 11 11 1 9 13 2
19 10 9 1 9 1 11 11 11 1 0 9 9 13 9 1 0 13 4 2
7 9 9 1 9 0 13 2
15 11 11 1 11 11 12 9 1 1 11 11 1 9 13 2
14 15 13 13 16 9 0 13 1 15 9 14 14 13 2
15 16 15 0 9 14 13 16 9 1 9 14 13 14 4 2
16 11 1 11 12 9 1 1 11 11 1 11 9 1 1 13 2
24 15 13 13 16 9 0 13 1 15 9 14 14 13 16 10 9 9 1 9 1 13 4 4 2
19 11 1 11 1 15 9 11 1 1 11 9 1 11 11 1 9 13 4 2
22 10 9 11 11 11 1 11 11 1 12 9 1 1 11 11 1 9 1 9 13 4 2
32 10 9 1 13 13 16 15 9 9 1 9 14 13 4 2 15 15 13 1 15 9 14 13 16 9 15 1 9 13 13 4 2
12 15 13 16 15 0 9 13 1 9 13 4 2
22 11 1 9 13 16 11 14 1 11 1 9 1 9 1 3 9 13 1 9 13 4 2
12 0 9 7 9 1 1 9 9 1 13 4 2
10 11 1 0 9 14 12 9 13 4 2
11 10 9 1 0 9 13 1 14 9 13 2
21 11 9 1 0 9 7 9 1 9 1 9 1 1 0 9 0 2 0 13 4 2
8 9 15 9 1 14 13 4 2
18 11 1 9 1 14 9 13 1 9 9 13 4 15 9 1 13 4 2
10 15 1 9 12 9 1 1 13 4 2
13 9 7 9 1 11 1 1 9 9 0 13 4 2
12 11 1 9 1 9 1 3 9 13 4 4 2
14 0 9 9 11 9 1 12 9 1 9 13 4 4 2
28 11 7 9 11 11 1 11 2 11 7 11 2 11 11 11 1 0 9 1 1 10 9 9 0 13 4 4 2
29 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 11 2 11 2 11 7 11 1 9 9 1 13 4 2
14 9 1 1 11 2 11 2 11 11 0 13 4 4 2
11 9 11 11 1 1 14 13 4 4 4 2
14 11 1 9 1 12 9 1 10 0 9 13 4 4 2
20 11 1 9 1 10 0 9 7 9 9 1 13 9 9 9 1 13 4 4 2
27 11 11 1 9 1 0 9 7 9 1 9 1 1 14 12 12 9 1 11 1 0 11 11 1 9 13 2
25 11 11 1 0 9 0 2 0 9 1 9 1 1 9 1 11 7 0 9 1 9 2 9 13 2
17 11 1 9 1 14 0 9 1 9 1 1 9 2 9 13 4 2
7 10 3 12 12 9 13 2
9 9 1 9 12 12 9 13 4 2
18 11 11 1 9 1 9 1 0 9 1 14 0 0 9 1 9 13 2
18 9 1 12 9 1 9 1 9 1 0 9 14 11 11 1 13 4 2
35 15 9 13 4 4 16 16 0 9 9 11 11 1 11 1 9 1 1 0 13 4 16 11 11 1 0 16 0 9 11 0 14 13 4 2
16 0 13 16 15 1 10 9 1 12 9 14 13 4 4 4 2
35 0 11 11 1 11 1 9 1 9 1 0 13 9 1 13 4 9 1 1 9 1 0 9 1 0 13 1 9 11 11 1 13 4 4 2
10 15 1 14 0 9 14 13 4 4 2
20 10 3 11 11 1 1 1 12 9 13 1 9 14 9 1 1 13 4 4 2
13 15 9 1 11 11 11 11 1 9 1 9 13 2
15 9 1 9 1 1 14 9 7 9 1 9 11 1 13 2
26 11 9 9 1 0 9 9 1 10 9 1 13 4 1 13 16 10 9 1 15 15 14 14 13 4 2
15 11 9 1 14 10 9 1 15 9 0 13 4 4 4 2
55 9 1 9 9 1 9 1 0 13 1 9 1 13 4 9 9 1 11 1 9 13 4 16 15 11 2 11 2 7 11 1 11 7 11 1 10 9 13 1 13 2 15 14 11 1 1 9 1 13 0 0 9 13 4 2
22 9 9 1 9 13 16 3 9 2 9 0 9 1 9 13 1 13 9 14 13 4 2
15 9 9 1 11 9 1 14 10 9 13 1 9 14 13 2
19 9 1 9 1 15 10 9 1 12 1 1 12 9 9 0 13 4 4 2
12 15 3 11 1 12 9 9 13 4 4 4 2
16 11 9 1 12 9 1 1 9 1 9 9 3 13 4 4 2
9 15 10 9 13 4 0 14 13 2
19 9 13 1 3 16 0 9 10 9 11 1 3 12 9 9 0 13 4 2
19 16 11 1 15 14 10 9 13 1 14 9 1 9 0 14 13 4 4 2
19 11 1 1 15 11 1 9 13 4 15 9 1 9 9 13 1 9 13 2
32 15 15 11 9 1 10 9 13 1 15 9 14 13 2 7 11 7 11 2 11 1 9 1 1 15 9 13 1 0 14 13 2
23 15 9 10 9 1 9 13 1 12 12 9 1 0 0 9 1 1 1 13 4 4 4 2
27 9 1 13 16 15 11 11 11 11 1 10 9 1 9 14 13 16 9 1 9 12 9 1 13 4 4 2
36 9 1 9 11 11 1 13 16 0 9 1 9 1 13 11 11 1 9 13 4 4 4 7 16 9 9 15 13 1 9 13 16 9 13 4 2
20 11 2 11 1 0 9 1 1 11 1 0 9 1 1 11 11 11 9 13 2
29 11 9 1 0 9 1 1 11 11 1 9 11 11 1 1 0 9 1 9 11 11 1 13 11 1 1 0 13 2
12 10 3 11 2 11 11 1 0 9 13 4 2
14 12 9 1 13 1 11 9 11 11 1 9 13 4 2
25 9 9 13 1 3 11 1 11 11 0 11 11 11 1 11 1 0 11 11 1 0 9 9 13 2
14 0 9 1 1 9 1 1 0 9 1 9 0 13 2
21 9 9 1 0 11 11 1 9 1 13 0 9 9 1 1 11 13 4 4 4 2
7 0 9 1 10 13 9 2
26 9 11 1 13 16 11 11 1 1 11 1 9 15 11 13 15 9 1 7 11 1 9 9 13 4 2
28 11 11 1 11 11 2 11 11 2 1 0 9 1 1 15 9 1 9 1 11 2 11 7 11 13 4 4 2
22 10 9 2 11 11 2 9 1 11 11 1 11 13 4 4 15 9 2 9 13 4 2
7 15 1 15 11 13 4 2
21 0 9 1 1 10 9 14 12 12 9 1 11 11 1 0 9 1 9 13 4 2
11 16 10 9 0 9 1 1 10 10 13 2
12 0 9 12 12 9 1 11 1 9 13 4 2
19 10 3 11 1 11 11 1 12 9 1 11 1 9 9 1 9 13 4 2
16 15 1 14 9 1 1 13 1 9 1 9 12 13 4 4 2
21 9 14 1 9 1 0 0 9 13 11 1 9 1 12 9 1 0 13 4 4 2
17 11 1 0 9 7 9 11 11 1 9 1 12 9 1 9 13 2
16 11 1 12 9 1 9 1 9 0 13 1 9 0 13 4 2
15 9 14 1 0 9 1 15 14 12 12 9 1 9 13 2
21 11 11 1 9 9 11 1 15 9 11 11 1 9 1 10 9 1 9 13 4 2
15 15 9 2 9 2 9 2 9 15 1 9 1 9 13 2
18 11 1 12 9 1 9 13 9 1 0 9 1 9 13 4 4 4 2
20 12 9 7 0 9 1 9 1 1 11 1 9 1 12 9 1 9 13 4 2
9 15 1 10 9 1 9 13 4 2
15 11 11 11 1 9 12 9 1 9 1 0 13 4 4 2
13 11 11 11 1 9 1 10 9 1 0 9 13 2
13 3 12 9 10 0 9 1 13 9 13 4 4 2
11 10 9 1 9 7 0 0 9 0 13 2
16 11 1 9 7 9 15 9 0 13 1 1 15 13 4 4 2
15 11 1 0 11 11 11 14 15 12 9 9 13 4 4 2
18 9 1 9 11 11 11 1 13 16 11 15 9 13 15 13 4 4 2
8 15 10 9 1 0 9 13 2
20 15 0 11 9 1 1 15 15 9 1 9 1 9 1 9 13 15 13 4 2
15 11 1 15 9 13 4 7 15 9 9 1 0 13 4 2
17 10 9 11 15 9 1 1 15 13 7 11 1 1 9 0 13 2
20 11 2 11 1 11 1 0 0 9 11 11 11 10 9 1 9 13 13 4 2
15 11 11 11 1 9 0 13 1 10 9 12 9 0 13 2
14 9 1 9 11 9 9 1 9 1 11 11 13 4 2
20 3 1 15 9 1 12 9 1 9 13 2 15 9 1 11 9 1 0 13 2
30 10 9 1 11 1 10 9 1 12 9 9 1 9 1 0 9 13 4 2 15 12 9 1 1 9 13 4 4 4 2
8 15 14 10 9 9 1 13 2
12 9 11 1 10 9 10 9 1 9 13 4 2
19 12 9 1 1 11 0 13 4 16 15 0 13 1 1 11 1 9 13 2
9 11 7 11 1 10 9 0 13 2
