80 11
13 0 2 0 0 9 9 9 1 2 15 13 4 2
13 0 9 14 14 2 11 9 14 9 9 0 13 2
20 3 2 15 9 2 11 9 11 9 9 13 4 14 13 4 14 9 11 13 2
25 10 9 2 0 11 9 9 11 14 2 0 9 14 14 11 11 2 11 9 0 9 14 13 4 2
18 15 9 9 9 13 4 14 2 9 9 13 13 4 14 9 11 13 2
17 11 9 0 11 11 9 11 9 0 9 9 0 14 15 9 13 2
5 15 13 14 2 2
10 9 9 13 14 2 3 9 14 13 2
10 9 9 0 9 2 9 9 13 4 2
18 9 9 3 13 0 9 1 13 4 0 9 9 9 14 13 4 4 2
18 3 2 10 9 2 11 2 11 9 9 14 9 9 13 4 15 9 2
25 11 9 9 14 9 9 14 9 10 9 13 9 9 13 4 14 2 3 13 4 14 9 11 13 2
11 11 13 11 9 11 9 11 9 13 4 2
18 11 9 14 2 3 9 13 1 11 9 14 11 0 9 3 13 4 2
4 9 14 12 2
30 11 9 0 12 9 9 13 11 11 14 2 0 12 9 9 13 9 14 2 0 12 9 9 13 11 11 14 9 13 2
12 11 11 12 9 13 9 9 0 9 14 11 2
22 9 9 9 0 9 14 14 2 9 14 2 9 14 0 9 14 14 10 9 13 4 2
14 9 0 11 1 0 0 9 14 9 13 14 9 9 2
43 10 9 2 15 0 9 14 2 9 14 13 9 1 13 0 9 11 3 9 13 9 9 13 4 4 14 13 2 11 9 9 0 11 9 13 13 14 11 15 9 13 4 2
24 11 9 9 0 9 13 9 9 1 11 9 0 9 9 13 14 9 13 0 9 13 4 4 2
12 11 11 7 11 9 11 9 9 11 9 13 2
49 9 11 9 0 9 9 11 11 2 11 9 9 11 11 2 11 11 2 11 11 9 0 9 9 9 11 11 2 11 9 9 11 11 2 11 9 9 11 11 2 11 11 2 11 11 9 13 4 2
18 11 11 11 9 14 2 11 11 11 9 14 15 9 1 9 13 4 2
10 9 1 9 13 2 0 9 13 4 2
14 9 11 0 11 9 1 13 2 9 9 9 3 13 2
11 9 9 13 11 9 10 9 14 13 4 2
8 9 9 9 11 9 13 4 2
4 9 13 4 2
8 3 11 9 14 9 3 13 2
16 3 2 11 9 2 9 9 3 15 13 11 9 9 9 13 2
18 3 2 11 9 0 9 13 11 9 0 9 12 11 9 1 9 13 2
25 11 11 11 9 11 11 2 11 9 11 9 11 11 9 9 10 9 13 14 10 9 13 4 4 2
10 11 9 11 11 9 0 9 13 4 2
19 12 9 9 14 9 11 9 0 3 13 14 11 14 11 9 11 11 13 2
31 11 11 9 11 9 1 0 15 2 11 11 9 12 9 9 14 9 3 13 1 2 0 9 14 3 13 14 9 13 4 2
13 12 9 9 3 11 9 0 9 11 11 9 13 2
11 12 9 0 0 9 9 3 9 3 13 2
24 3 12 9 14 0 9 9 13 1 2 3 0 0 9 7 9 3 13 1 14 9 13 4 2
14 9 3 0 9 13 0 9 13 14 10 9 3 13 2
14 11 7 11 1 11 14 11 14 3 9 13 4 4 2
14 15 1 2 11 9 0 9 0 9 14 3 13 4 2
10 9 11 0 9 13 9 13 4 4 2
21 15 1 11 9 1 9 7 9 9 1 9 13 14 2 15 13 1 14 13 4 2
12 12 9 14 3 11 13 1 14 3 13 4 2
15 12 9 14 1 9 1 11 9 0 9 3 13 1 13 2
18 3 9 9 2 13 0 11 9 2 9 13 1 14 12 9 14 13 2
19 11 2 11 9 14 9 0 9 1 0 9 9 9 13 14 9 13 4 2
14 12 9 9 14 9 9 3 9 9 14 9 1 4 2
16 9 9 9 13 9 14 3 12 9 14 3 0 9 13 4 2
20 11 9 1 13 9 9 9 9 14 9 9 13 14 11 9 14 9 3 13 2
13 3 11 9 9 11 1 14 9 0 9 13 13 2
19 9 2 11 9 9 2 9 9 2 11 9 9 3 13 14 9 13 4 2
13 3 11 9 9 9 0 9 9 13 11 11 13 2
14 3 9 9 0 9 11 13 14 13 14 11 11 13 2
31 0 9 0 11 11 9 13 11 9 9 14 11 9 7 11 9 9 2 11 2 9 9 9 13 4 14 11 9 13 4 2
8 15 0 9 14 11 13 4 2
13 12 9 14 0 9 9 0 11 11 9 13 4 2
18 11 9 15 0 9 13 11 1 3 13 11 9 3 13 13 11 11 2
24 11 1 9 13 4 9 1 11 9 11 11 3 13 4 14 9 13 4 11 9 9 11 11 2
11 15 9 9 13 3 13 14 14 15 13 2
19 11 9 9 13 11 7 11 0 9 9 0 9 9 0 14 15 3 13 2
6 11 1 9 13 4 2
14 0 9 2 11 2 3 13 9 13 4 4 14 13 2
10 3 3 15 9 13 14 15 9 13 2
8 11 0 9 9 13 11 13 2
33 0 11 11 2 11 9 13 14 9 7 11 11 2 11 11 9 13 14 9 15 12 14 14 0 2 9 9 13 9 9 13 13 2
12 3 15 2 11 2 11 2 9 9 3 13 2
13 15 11 9 14 9 14 0 9 14 13 9 13 2
19 9 2 9 2 9 2 9 2 9 2 11 14 9 1 14 0 9 11 2
11 15 1 9 14 11 9 13 4 13 11 2
9 3 14 11 0 9 14 3 13 2
8 3 13 9 13 14 9 13 2
4 3 3 13 2
4 9 1 13 2
10 9 9 0 9 13 3 13 13 15 2
22 11 11 9 9 9 9 1 0 0 9 11 9 9 1 3 13 4 4 14 15 13 2
11 0 0 9 1 12 12 12 11 13 4 2
13 3 3 10 9 9 2 9 13 13 4 13 15 2
15 11 11 9 9 0 14 11 9 11 11 9 10 13 4 2
