271 11
15 13 1 15 10 0 9 1 10 11 2 13 3 1 11 2
3 10 11 0
20 2 11 2 13 10 9 1 9 0 2 9 9 2 7 10 9 1 10 9 2
32 10 9 13 10 9 1 10 9 0 1 10 0 9 0 1 11 2 13 1 10 9 0 15 13 3 10 9 1 9 7 9 2
18 1 13 10 9 0 1 10 9 2 11 13 3 3 3 1 10 9 2
23 10 9 1 11 13 13 11 1 10 9 0 2 1 13 10 9 1 13 9 0 1 0 2
18 10 9 1 10 9 3 13 10 9 0 2 10 9 1 10 9 0 2
9 9 1 10 9 1 10 11 13 9
26 10 9 3 1 10 0 11 1 11 13 10 9 1 10 9 1 10 9 0 1 10 9 1 10 9 2
29 10 11 1 10 11 13 10 9 1 10 3 12 9 0 2 15 3 13 9 0 1 9 2 1 10 9 1 11 2
32 16 10 9 3 13 9 2 7 13 13 1 15 2 10 9 13 13 3 3 10 3 0 2 15 3 13 9 1 10 9 0 2
24 10 9 13 0 16 13 2 3 2 10 9 1 10 9 2 1 10 9 2 1 10 9 0 2
26 13 10 9 0 1 0 9 2 15 13 13 0 7 0 2 1 10 10 9 13 0 13 15 13 13 2
18 9 1 10 11 2 11 2 2 1 12 2 13 16 12 9 1 9 2
14 1 10 9 2 12 9 13 9 7 12 9 2 9 2
19 10 9 13 1 12 7 12 9 1 9 7 10 9 2 1 12 7 12 2
6 11 13 12 1 13 9
3 1 10 11
15 10 11 2 11 2 13 3 12 9 1 13 9 1 9 2
21 13 13 10 9 1 10 9 11 2 11 2 7 10 9 11 2 1 10 9 11 2
26 15 12 13 13 3 10 9 11 2 12 2 13 13 9 12 1 11 3 9 1 10 9 1 10 11 2
10 15 13 13 1 12 9 1 10 11 2
9 12 1 15 13 10 9 2 11 2
4 9 13 10 9
35 1 10 9 2 10 9 1 10 9 1 10 9 11 13 1 13 10 9 1 10 9 13 1 10 9 13 1 10 10 9 1 10 9 0 2
21 10 9 1 10 9 0 13 13 10 9 1 10 9 0 1 10 9 1 9 0 2
15 1 10 9 1 10 10 9 0 2 10 9 13 3 0 2
11 15 13 3 9 1 9 1 10 9 13 2
35 10 9 3 0 1 10 9 1 10 9 1 11 13 1 16 15 13 9 1 9 1 9 15 13 13 1 10 9 1 9 0 1 10 9 2
22 1 10 10 9 2 13 10 9 0 1 0 9 13 10 9 2 15 13 10 9 0 2
21 11 13 16 3 10 9 1 9 9 13 9 12 2 3 10 9 13 1 9 12 2
10 11 13 10 9 1 13 1 10 9 2
34 10 9 13 4 13 1 10 9 1 10 9 2 2 3 13 16 13 10 9 7 3 13 3 2 13 9 15 15 13 1 13 10 9 2
20 3 1 10 9 2 10 9 13 7 13 13 13 7 3 13 13 15 13 2 2
35 10 9 3 13 0 1 10 9 2 16 1 13 15 9 0 1 13 7 13 9 2 15 3 13 10 9 1 9 3 13 1 10 9 0 2
7 11 2 12 2 9 12 2
26 10 9 2 13 1 9 7 9 2 13 10 9 1 9 0 1 10 9 1 10 9 1 10 9 12 2
15 15 3 13 13 1 10 9 2 13 13 10 9 1 9 2
7 9 2 12 11 2 3 2
14 9 2 1 10 9 12 2 1 10 9 1 10 0 9
4 9 2 13 15
3 9 1 9
24 1 9 1 10 11 1 9 2 1 11 2 10 9 13 16 9 3 3 13 15 13 1 9 2
24 2 10 9 13 13 1 10 9 15 15 13 1 10 9 2 1 10 9 7 1 10 9 0 2
4 9 13 0 2
7 15 3 15 13 1 9 2
10 1 15 9 7 9 13 9 0 2 2
11 11 2 15 10 9 13 3 2 1 9 2
13 9 7 9 13 9 15 13 10 2 9 11 2 2
20 9 1 10 9 1 9 7 9 13 9 0 1 15 13 1 10 0 1 10 11
28 10 9 1 9 1 10 11 13 13 3 10 9 1 9 7 10 9 1 9 3 9 1 15 13 1 10 9 2
18 13 15 15 13 10 9 1 10 11 2 13 3 1 10 0 9 0 2
15 11 13 13 10 13 9 2 11 2 2 1 10 9 0 2
17 3 1 10 11 2 11 13 10 9 1 10 9 1 2 11 2 2
25 11 13 13 1 10 9 1 10 9 2 11 2 2 15 13 10 9 11 1 10 9 1 12 9 2
15 7 10 9 1 9 12 9 13 16 10 9 3 13 0 2
24 13 0 9 3 10 9 1 10 9 2 11 2 2 15 13 10 9 13 1 11 1 12 9 2
24 11 13 9 3 9 0 2 13 13 1 11 1 12 9 2 7 10 9 3 13 1 10 9 2
25 1 10 9 0 2 11 7 11 13 1 9 13 1 10 9 1 10 11 1 10 9 1 10 9 2
18 11 13 10 9 1 10 9 1 9 2 15 13 10 9 1 9 0 2
17 13 15 2 1 15 2 1 10 2 9 1 9 1 10 9 2 2
17 3 2 1 10 9 0 1 0 9 2 15 13 1 13 10 9 2
41 1 15 2 3 2 13 0 16 10 10 11 13 3 10 2 9 2 1 10 9 2 15 13 0 2 7 16 13 1 2 13 15 2 1 10 10 9 0 1 9 2
7 9 1 10 11 13 1 9
10 10 9 11 3 13 10 9 1 11 2
11 3 2 13 13 9 1 9 1 10 9 2
20 10 9 2 1 9 1 9 1 10 10 9 2 13 13 10 9 1 10 9 2
9 9 13 1 10 9 1 10 9 2
20 1 15 2 15 13 1 10 9 1 9 0 1 9 0 2 1 9 1 12 2
21 2 3 1 10 9 2 10 11 0 13 1 13 10 9 1 10 9 1 10 11 2
32 10 11 1 10 11 13 1 13 1 10 9 7 1 13 15 1 13 10 9 1 15 2 3 2 13 10 9 2 2 13 11 2
17 10 9 1 10 0 9 0 13 1 9 0 2 13 1 10 11 2
10 3 13 9 1 10 9 1 10 9 2
9 10 9 13 13 3 1 10 9 2
18 10 11 13 11 2 11 2 2 11 7 11 2 11 2 2 1 15 2
14 13 10 9 1 15 10 9 13 1 9 7 1 15 2
30 1 9 15 10 10 9 13 2 1 10 9 1 10 9 1 10 9 0 2 10 9 3 3 13 10 0 9 1 11 2
23 10 9 0 13 1 10 9 0 2 1 15 11 13 1 10 9 2 16 0 1 9 0 2
20 13 15 10 12 9 7 10 9 15 13 2 13 9 7 3 2 3 2 9 2
28 13 15 2 3 2 10 9 0 15 13 1 10 9 1 12 2 3 10 9 0 2 1 10 9 1 10 11 2
10 3 13 10 9 1 10 9 1 13 2
15 11 2 11 2 11 7 3 10 11 13 9 1 10 9 2
10 10 9 13 16 10 9 13 13 13 2
19 15 13 13 13 1 10 9 1 9 1 9 1 13 1 10 9 1 13 2
24 10 9 13 9 1 10 11 2 11 2 1 10 11 1 13 10 9 1 10 9 1 10 9 2
17 1 10 9 2 10 9 1 11 3 13 13 10 9 1 10 9 2
3 9 7 9
13 10 9 13 13 10 11 1 13 9 2 13 11 2
21 2 10 11 13 13 1 12 9 2 7 12 1 10 9 13 10 15 1 10 11 2
12 13 13 9 2 3 1 10 9 2 2 13 2
23 1 10 9 0 2 3 13 13 1 11 1 13 9 0 2 7 13 9 0 1 10 9 2
27 2 1 10 9 1 9 1 10 9 2 13 13 10 9 1 10 9 0 1 10 9 0 16 15 13 11 2
15 3 2 1 10 9 0 1 10 0 12 9 2 2 13 2
1 9
19 13 13 16 3 13 1 12 9 1 13 10 9 2 13 1 10 9 0 2
8 2 12 9 1 9 13 9 2
33 15 13 13 10 9 0 2 1 15 15 13 10 9 11 2 11 2 1 10 9 2 2 1 10 9 1 10 11 2 1 12 9 2
9 7 15 13 13 1 12 9 2 2
17 15 13 10 9 1 10 9 1 10 9 1 10 2 9 0 2 2
20 2 10 9 13 16 13 9 12 2 7 12 9 3 10 9 13 3 0 2 2
10 13 10 9 2 11 13 10 9 13 2
5 10 9 15 13 2
11 15 13 1 10 9 1 10 9 2 9 2
5 9 11 13 1 9
35 10 9 11 2 1 10 11 2 13 9 9 1 10 9 2 9 2 1 10 9 1 10 0 9 1 10 11 1 11 2 9 1 10 11 2
31 10 9 15 13 11 3 3 13 9 1 9 7 13 13 3 1 10 9 1 10 9 1 12 9 1 10 9 1 10 9 2
53 11 7 11 13 10 11 10 9 1 10 11 2 11 2 7 1 10 11 2 11 2 13 3 10 9 1 2 11 2 1 10 11 2 9 0 0 2 13 1 10 11 2 2 15 13 9 0 1 9 1 10 11 2
17 1 15 2 10 9 1 10 9 3 13 13 10 9 1 10 11 2
22 3 13 9 2 3 13 11 2 16 10 9 13 1 11 13 13 2 9 1 9 2 2
10 10 9 0 3 13 10 9 1 9 2
22 10 9 1 9 13 13 1 10 9 11 7 11 2 1 10 11 2 3 1 10 11 2
13 13 1 9 1 10 11 2 13 13 1 12 9 2
18 10 0 1 15 2 1 10 9 1 12 9 2 13 9 1 12 9 2
5 11 13 10 12 9
19 11 2 12 2 9 2 2 13 3 1 10 9 1 11 1 10 9 0 2
6 15 13 13 1 9 2
20 13 4 13 1 10 9 2 3 10 9 11 2 12 2 13 1 10 10 9 2
13 11 13 13 1 12 13 7 3 13 9 1 9 2
6 9 13 9 1 10 9
23 9 1 10 9 1 10 11 13 10 9 1 10 9 0 1 11 2 10 0 1 10 9 2
16 10 9 13 1 3 12 9 1 11 2 10 9 1 10 9 2
17 10 9 13 1 12 9 1 10 9 1 10 9 11 7 10 9 2
8 2 3 13 9 1 13 15 2
19 10 9 1 10 9 1 9 13 0 2 2 13 11 2 9 1 10 11 2
8 10 9 1 10 9 13 0 2
26 7 2 13 11 2 9 1 10 11 2 2 13 3 1 10 9 1 9 16 13 1 9 3 13 2 2
9 9 11 13 16 13 9 1 10 11
28 10 11 13 1 13 10 9 0 1 10 0 9 2 9 1 10 11 2 1 9 1 10 0 9 1 10 11 2
35 10 9 11 2 13 1 10 9 1 10 9 1 10 9 1 12 1 12 1 11 3 2 13 2 16 13 13 9 7 9 1 10 9 2 2
19 11 3 13 9 16 10 9 11 13 10 10 9 2 13 1 12 1 9 2
20 2 16 15 13 2 13 16 13 0 2 1 10 9 3 13 3 2 2 13 2
4 13 15 13 11
34 13 1 10 9 12 1 9 1 12 2 1 11 2 11 13 10 9 0 1 10 9 2 1 12 2 3 13 9 0 1 10 9 0 2
24 1 12 2 1 13 10 9 0 7 0 1 10 9 2 11 13 10 11 2 13 1 0 9 2
6 11 13 9 1 10 11
3 2 9 2
11 2 11 2 2 9 1 9 2 11 2 12
9 9 13 12 9 1 9 1 10 11
16 10 11 2 11 2 13 9 12 9 1 10 11 2 1 11 2
11 15 3 13 9 1 9 13 1 10 9 2
15 10 9 1 9 15 13 10 9 13 13 1 9 12 12 2
24 1 11 2 9 1 10 9 2 3 13 13 12 9 1 10 10 9 1 10 9 1 10 9 2
6 11 13 9 1 10 11
37 10 11 13 13 10 9 1 9 1 10 11 2 9 0 1 9 1 10 9 1 10 9 1 10 9 2 1 11 2 9 1 10 9 1 10 11 2
17 10 9 13 13 1 10 9 1 10 9 0 2 1 10 0 9 2
10 10 9 0 13 13 1 10 9 12 2
15 11 13 10 9 1 13 1 10 9 2 13 13 10 9 2
16 2 3 15 13 13 9 0 1 10 9 16 10 9 13 2 2
19 10 9 11 2 9 13 1 13 13 9 0 1 10 9 2 3 13 13 2
7 2 13 10 9 3 0 2
17 3 2 10 9 13 13 10 9 3 1 9 7 3 1 9 2 2
10 1 10 9 2 11 13 13 10 9 2
11 2 11 13 10 9 1 13 15 13 2 2
53 13 1 10 9 1 10 9 1 12 2 9 0 1 10 9 9 1 9 7 9 0 7 13 1 13 1 10 9 13 1 10 9 11 1 10 11 2 10 9 13 9 1 9 2 1 9 1 10 0 9 1 9 2
5 9 2 9 12 2
18 10 9 13 10 9 1 9 1 10 9 1 10 11 2 1 10 11 2
18 13 10 9 0 2 1 11 7 11 2 9 15 1 10 9 15 13 2
15 16 15 13 2 15 13 13 1 9 3 13 1 10 11 2
43 9 1 10 11 1 10 11 2 13 1 10 11 2 13 9 1 10 9 2 9 1 9 2 13 1 10 9 1 10 11 3 1 9 7 9 0 1 16 10 0 13 13 2
28 1 10 9 2 13 0 10 9 1 10 9 0 1 10 11 1 16 15 13 10 9 0 1 15 1 10 11 2
9 2 13 13 10 9 1 12 9 2
9 13 3 0 16 1 3 12 9 2
14 13 4 13 2 3 2 1 13 10 9 1 12 9 2
11 13 10 9 0 2 2 13 11 2 12 2
32 10 9 15 13 1 10 9 1 11 13 10 9 11 2 15 13 13 1 10 11 2 16 10 9 1 10 11 13 10 10 9 2
26 1 10 9 2 11 2 10 0 9 1 10 9 1 10 9 2 13 3 10 0 9 1 10 9 0 2
28 1 10 9 2 10 3 9 13 1 10 11 2 1 9 1 10 9 15 2 1 10 9 2 13 1 10 11 2
25 3 2 10 9 13 10 9 1 9 12 12 0 1 10 11 2 15 13 1 10 9 1 10 11 2
27 10 9 1 10 9 13 3 1 10 9 1 10 9 7 1 10 9 2 0 1 10 9 1 10 9 0 2
26 1 10 11 2 10 9 13 1 9 12 9 1 12 1 9 12 9 1 12 2 7 10 12 9 2 2
27 1 10 9 2 10 9 13 1 12 9 2 13 10 9 1 9 12 9 1 12 1 9 12 9 1 12 2
1 9
39 10 9 11 2 11 2 13 3 9 1 10 9 1 10 9 0 1 9 1 9 1 12 2 13 16 10 9 13 10 9 0 1 9 12 9 1 10 9 2
28 16 13 1 3 12 9 1 10 9 2 10 9 13 13 16 13 1 10 11 2 3 10 11 13 1 10 9 2
15 10 9 1 10 9 13 1 10 9 2 9 1 11 2 2
9 10 10 9 13 3 1 10 9 2
10 10 9 7 11 3 13 1 10 9 2
17 1 13 10 9 2 1 10 12 9 1 9 10 9 13 10 9 2
12 10 11 1 11 13 1 12 9 1 9 0 2
1 9
38 0 1 9 2 10 9 1 10 11 1 10 11 13 13 3 1 10 9 1 10 9 2 1 3 12 9 3 2 7 13 10 9 1 9 1 10 9 2
24 10 9 10 13 10 9 1 9 1 10 11 2 15 13 3 3 10 9 16 10 11 1 11 2
28 1 15 3 1 10 9 7 9 1 11 11 13 10 9 0 2 1 9 1 10 9 1 11 2 11 7 11 2
25 3 13 13 9 0 1 10 9 2 13 11 2 7 13 3 10 9 1 13 10 0 9 1 9 2
22 1 11 2 12 2 9 1 10 11 2 2 3 15 13 13 3 12 9 1 9 2 2
22 1 15 2 9 3 13 13 16 13 13 10 9 1 9 1 10 9 1 10 9 0 2
7 9 0 3 13 10 9 9
3 9 1 9
23 10 9 13 13 13 1 10 11 1 9 1 12 2 16 10 9 13 4 13 12 9 3 2
27 13 1 10 11 2 11 2 2 10 9 0 13 13 1 15 1 10 9 2 11 2 11 7 11 2 3 2
20 7 2 3 1 10 9 2 10 9 1 10 9 0 13 10 9 1 9 13 2
27 10 9 1 10 9 9 7 10 9 1 9 1 9 13 2 13 9 1 10 9 12 2 13 9 3 0 2
18 2 13 1 10 9 2 2 13 1 10 11 11 2 9 1 10 11 2
18 15 13 2 3 2 16 3 10 2 9 9 13 9 1 0 9 2 2
7 9 13 13 13 1 10 11
24 11 13 12 9 13 2 13 7 1 9 13 2 1 10 9 1 10 9 11 2 9 0 2 2
17 11 7 11 13 13 4 13 1 9 2 15 15 13 13 1 9 2
10 9 13 13 1 9 1 9 1 10 11
30 9 1 10 11 7 11 1 10 11 13 13 1 9 3 1 10 9 1 10 11 2 11 2 9 0 1 10 11 2 2
6 10 9 13 9 0 2
9 1 10 9 2 13 11 2 12 2
19 10 9 13 13 1 10 9 11 2 12 2 13 1 12 9 1 10 11 2
18 10 9 13 0 1 10 11 1 10 11 2 13 1 10 11 1 12 2
9 9 13 11 7 13 1 9 1 11
38 10 9 0 0 1 9 13 10 9 1 10 11 2 10 9 0 13 1 11 2 11 2 7 15 13 1 10 9 1 10 9 1 11 2 11 7 11 2
39 10 9 13 1 10 9 11 13 1 10 9 1 13 3 1 10 9 1 10 9 10 0 9 1 11 1 12 1 12 2 12 1 12 1 10 0 9 2 2
13 10 9 1 10 9 13 11 2 15 13 12 9 2
22 1 10 9 1 10 9 2 13 1 10 9 10 11 7 10 11 2 0 9 1 9 2
28 10 0 9 1 10 9 13 10 9 11 2 13 1 13 9 1 9 1 9 2 15 13 13 1 12 12 11 2
19 9 1 10 9 11 2 15 13 9 7 13 13 1 10 9 1 10 9 2
22 2 10 11 13 3 12 9 1 9 7 10 9 0 2 2 13 10 9 1 10 11 2
18 1 11 2 10 9 13 10 0 9 1 10 9 1 9 1 10 9 2
17 11 15 13 10 9 15 10 9 13 13 1 10 9 13 10 9 2
15 13 1 10 9 2 13 13 0 9 7 13 1 10 9 2
11 9 0 15 13 1 10 10 9 1 9 2
6 3 13 9 3 0 2
14 11 10 9 3 13 9 15 13 1 13 1 10 9 2
20 10 9 13 0 7 10 11 13 13 3 10 9 0 3 9 1 10 0 9 2
20 10 9 7 10 9 13 1 13 10 9 0 2 3 2 13 3 1 9 0 2
2 9 0
21 13 1 9 1 10 11 10 9 1 9 1 13 10 9 1 9 1 10 0 9 2
17 15 13 13 1 11 2 3 9 1 10 13 9 1 10 9 0 2
2 9 0
34 13 0 9 2 1 10 0 2 10 9 1 10 9 1 10 9 2 11 2 1 10 9 15 13 1 10 9 1 9 1 10 9 0 2
15 13 0 2 13 0 1 10 9 7 13 3 1 10 9 2
6 11 1 10 9 1 11
33 1 2 11 2 2 11 2 1 11 2 11 13 10 9 1 15 10 2 10 0 9 2 0 0 2 15 13 1 13 1 10 9 2
9 13 3 10 0 9 1 10 9 2
25 11 13 10 0 11 1 13 10 10 9 2 10 1 10 9 15 13 1 10 0 0 10 0 9 2
13 2 11 2 13 10 9 1 10 9 1 10 9 2
21 11 2 11 2 13 10 9 1 10 9 1 9 9 1 9 2 11 7 11 2 2
41 11 3 13 1 9 1 10 9 2 13 1 10 9 1 11 2 7 3 13 1 10 9 1 10 9 2 15 13 1 15 13 2 11 13 0 1 2 11 2 2 2
31 16 10 9 13 10 11 2 13 13 10 10 9 3 1 10 9 3 1 10 9 2 2 13 15 16 10 0 13 10 0 2
21 13 2 1 10 9 3 0 1 10 9 2 10 11 13 9 3 0 16 10 11 2
6 13 1 12 1 12 2
19 3 13 2 1 9 1 10 11 2 16 10 11 3 13 13 1 10 9 2
13 7 3 1 10 11 3 10 11 13 10 9 0 2
18 10 9 13 1 10 9 2 11 2 15 15 13 0 1 10 12 9 2
13 1 10 9 13 3 9 2 9 7 9 1 9 2
5 10 9 13 0 2
13 15 13 2 13 1 9 1 10 9 0 2 11 2
37 1 13 16 10 10 9 13 2 3 2 10 10 9 11 2 3 1 10 9 1 10 11 2 12 1 12 2 1 10 9 1 10 9 1 10 11 2
21 3 10 9 13 1 10 9 1 11 2 10 9 11 15 13 1 13 10 10 9 2
12 2 13 1 3 2 6 2 3 1 11 2 2
7 3 11 13 1 10 9 2
16 1 10 12 9 1 10 0 9 2 3 12 13 1 10 9 2
10 1 10 12 0 9 2 12 13 9 2
8 10 15 13 10 9 1 11 2
17 9 0 1 10 15 13 13 2 9 7 10 3 0 9 1 9 2
22 10 11 3 13 7 10 9 1 10 9 3 13 3 13 10 0 9 1 10 9 0 2
5 10 9 2 11 2
5 10 9 2 12 9
43 1 10 9 0 1 10 9 15 13 10 12 0 9 1 10 9 0 2 10 9 2 9 7 9 1 10 11 11 7 10 9 1 10 11 7 9 1 10 9 1 9 11 2
15 11 13 16 10 9 1 10 9 13 13 3 1 10 9 2
11 2 9 13 3 2 7 9 13 10 11 2
11 2 9 13 3 2 7 9 13 10 11 2
4 9 1 9 2
28 2 10 9 13 3 0 16 13 16 13 1 13 10 10 9 0 1 12 9 2 2 13 11 2 1 10 11 2
10 13 9 15 13 9 1 9 1 9 2
18 10 9 13 10 9 1 10 11 2 1 12 9 1 9 1 11 2 2
24 11 3 13 13 9 1 9 2 16 3 3 13 13 7 13 13 1 9 1 9 1 10 9 2
23 7 15 13 16 13 15 13 2 3 10 0 2 1 9 15 13 10 9 1 10 9 0 2
19 11 2 10 9 13 16 10 9 13 9 1 9 2 1 9 7 1 9 2
19 11 1 10 9 1 10 9 2 15 13 3 10 9 1 9 7 1 9 2
10 15 13 3 13 1 13 10 9 0 2
21 10 9 13 10 9 15 13 1 10 0 10 9 1 9 2 13 15 10 9 0 2
6 9 0 13 11 1 11
12 11 13 10 0 9 1 10 11 1 10 9 0
34 10 9 11 2 9 1 0 9 1 10 9 2 13 13 1 10 0 9 1 10 11 1 11 2 15 13 10 12 0 9 1 10 9 2
32 11 2 9 12 1 10 9 0 2 13 1 10 9 0 1 10 9 11 1 12 2 12 7 12 2 1 12 1 10 9 0 2
18 1 10 0 9 1 10 9 2 11 13 13 1 10 9 1 10 11 2
