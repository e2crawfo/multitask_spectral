150 17
10 15 14 13 1 10 9 15 3 3 2
48 2 3 13 15 3 10 9 9 7 13 1 10 9 15 2 7 13 15 10 9 0 14 13 15 3 2 9 0 9 14 13 1 12 9 1 9 7 12 1 9 2 7 3 12 9 1 9 2
99 2 13 10 9 16 13 3 0 1 11 11 2 10 9 9 1 9 9 2 9 7 9 1 9 10 9 14 13 1 1 9 12 8 1 9 10 11 2 12 2 8 12 1 12 2 1 9 1 10 9 9 7 9 2 9 1 9 10 9 7 1 9 10 9 2 2 12 2 8 8 12 1 12 2 2 7 1 10 9 9 2 9 7 9 2 11 9 9 2 2 12 2 8 8 12 1 12 2 2
32 1 9 10 14 13 9 1 9 10 11 1 11 8 11 1 10 9 1 11 3 16 14 13 15 0 1 9 9 10 9 0 2
26 13 9 1 9 1 15 7 1 10 9 9 1 9 7 13 9 13 15 10 9 14 0 1 11 15 2
9 10 11 13 0 1 14 9 3 2
28 2 13 9 11 0 1 11 7 1 9 10 11 1 9 14 9 1 9 1 9 10 7 1 9 1 11 11 2
30 2 11 13 14 11 14 9 3 16 14 13 1 9 14 13 9 1 1 9 11 7 14 13 15 9 1 15 14 9 2
15 9 10 9 1 9 10 11 11 14 11 9 10 9 0 2
4 3 1 9 2
13 13 9 9 1 10 9 2 7 13 9 0 1 2
19 13 11 10 9 1 9 10 9 16 13 1 11 7 1 11 9 10 9 2
23 1 10 9 14 13 1 9 13 9 1 9 10 11 11 7 9 9 1 9 1 8 9 2
18 2 14 13 15 9 7 9 9 7 10 9 1 9 1 2 14 9 2
32 2 11 2 10 9 0 15 2 2 13 10 11 2 2 16 13 9 1 1 10 9 2 7 16 13 15 9 1 10 9 1 2
41 13 1 10 9 11 9 0 14 0 14 13 9 2 15 7 10 9 0 14 13 10 9 2 10 9 2 9 10 9 2 7 10 9 0 1 10 9 9 10 9 2
13 13 0 1 9 14 13 9 1 9 1 9 10 2
20 13 3 1 12 9 0 9 7 9 9 1 9 1 9 2 1 9 1 9 2
26 13 10 9 1 1 9 9 14 13 1 9 1 9 9 9 10 9 14 13 10 9 1 9 3 1 2
16 11 14 11 11 0 7 9 11 14 13 9 0 11 14 0 2
26 12 2 14 13 9 10 9 0 14 13 9 10 11 2 9 11 2 1 9 1 1 2 9 0 2 2
10 10 9 10 14 13 1 9 0 9 2
16 1 9 10 9 0 1 9 9 14 13 10 9 0 9 3 2
15 7 9 9 7 9 1 9 0 10 9 9 9 1 12 2
21 13 10 9 9 9 1 10 11 9 14 9 1 9 0 10 16 14 13 9 1 2
17 13 0 14 13 9 1 12 9 10 1 3 2 13 12 1 11 2
6 13 10 9 1 9 2
15 13 9 11 1 9 1 9 13 9 0 0 14 13 1 2
37 13 15 10 9 7 10 9 15 7 13 1 9 1 16 9 0 2 1 9 1 9 1 13 0 10 9 15 14 9 1 9 1 9 7 1 9 2
29 13 9 1 3 2 7 15 9 2 16 1 9 10 9 13 0 1 10 9 2 7 13 1 1 9 1 9 15 2
13 13 10 9 0 7 13 10 9 0 1 10 9 2
11 1 9 14 13 9 15 2 1 10 9 2
18 14 13 1 9 15 2 14 13 1 9 15 2 14 13 1 9 15 2
9 13 13 14 0 14 13 10 9 2
22 13 10 11 10 9 1 9 9 2 9 7 9 16 13 15 10 9 14 9 1 9 2
11 13 9 1 1 9 3 1 10 9 10 2
8 9 1 9 14 13 9 9 2
41 13 11 14 11 1 11 11 9 10 9 10 1 2 13 9 15 1 9 14 13 1 9 9 1 9 11 11 7 14 13 3 1 9 9 10 9 10 2 11 11 2
23 13 1 1 10 9 10 14 13 15 9 14 13 14 0 1 10 9 14 9 1 10 9 2
37 13 0 12 9 1 9 14 9 1 12 9 12 1 2 2 9 10 11 2 2 10 9 2 9 10 11 0 2 9 11 2 9 9 2 8 11 2
10 2 13 15 10 15 2 2 13 15 2
9 13 10 9 10 14 13 1 9 2
19 1 9 14 13 9 1 9 15 1 13 15 10 9 0 14 13 9 1 2
16 13 9 9 1 1 9 1 2 1 9 3 7 1 9 9 2
75 13 9 1 10 9 1 10 9 2 11 11 2 1 11 11 11 1 9 10 11 2 1 10 9 13 3 1 2 14 0 1 9 9 9 2 9 9 7 9 1 11 11 10 9 1 10 9 0 2 9 1 9 10 11 2 9 14 13 1 9 1 9 14 13 1 9 1 16 10 2 11 9 11 2 2
90 8 1 10 9 2 9 2 9 7 9 14 13 1 9 7 14 13 1 9 1 7 14 13 1 9 9 1 9 10 9 1 9 1 9 2 13 15 7 15 2 1 10 9 10 7 1 9 2 0 2 1 1 7 1 9 1 9 2 1 10 9 10 9 14 13 15 7 15 1 9 14 13 1 9 1 9 10 9 10 7 14 13 0 7 0 1 10 9 10 2
8 14 8 8 7 14 8 15 2
22 13 10 12 9 1 9 9 9 3 1 15 2 16 14 13 15 3 1 9 9 1 2
13 13 11 14 0 16 13 9 0 1 9 1 3 2
27 2 13 15 14 13 9 9 9 1 10 9 1 12 9 14 13 3 2 7 13 15 14 13 10 9 0 2
11 9 11 12 2 12 9 11 12 2 12 2
11 13 9 1 9 10 11 14 13 3 3 2
26 13 11 11 2 10 12 9 10 1 10 9 7 10 12 9 10 3 2 1 9 1 9 10 11 11 2
137 12 13 9 10 9 13 1 9 1 9 10 9 10 1 9 10 9 1 9 9 1 10 9 13 1 10 9 8 7 1 10 9 14 13 1 7 14 13 1 15 1 7 2 1 10 9 10 1 9 2 13 15 1 9 1 9 9 10 9 14 13 10 9 8 1 9 10 9 8 1 9 2 1 14 13 10 9 10 15 2 7 3 10 9 2 9 0 2 9 2 7 9 10 2 1 14 13 9 1 1 9 1 15 15 14 9 1 9 2 14 13 10 9 10 14 0 1 9 13 0 10 9 0 1 9 8 7 15 1 9 9 0 1 9 3 1 2
16 13 15 1 9 10 9 14 9 1 10 9 1 9 1 12 2
47 13 15 0 1 9 0 2 7 14 0 1 15 13 9 1 9 3 1 9 10 11 7 9 14 9 1 9 10 9 0 1 9 1 11 2 13 9 0 3 0 3 7 3 14 13 1 2
33 16 2 1 15 10 14 9 13 14 11 9 1 9 9 9 10 9 2 13 15 10 14 13 10 9 9 7 9 0 1 9 0 2
19 2 13 10 9 10 1 1 9 1 9 9 14 13 0 1 10 9 0 2
60 8 16 9 15 2 3 2 14 13 10 9 1 9 0 2 13 15 2 3 0 16 14 13 1 10 9 7 1 9 14 13 1 9 1 1 9 1 1 9 0 2 1 9 10 9 0 14 13 10 9 14 13 1 9 1 9 1 10 9 2
7 13 15 13 1 9 9 2
18 13 10 9 1 9 0 1 9 10 9 12 1 9 11 11 3 3 2
34 13 9 0 3 1 10 9 1 9 14 9 1 9 1 9 0 2 16 10 9 0 2 13 9 0 15 15 1 9 1 9 1 9 2
17 9 14 13 9 0 1 10 9 2 13 9 3 1 10 9 0 2
23 13 15 15 11 8 11 2 0 10 11 11 11 2 10 9 11 8 11 7 11 8 11 2
28 14 0 13 9 1 11 0 1 9 1 9 14 9 1 9 7 1 9 0 14 9 1 10 9 14 13 15 2
24 13 9 9 7 9 1 9 1 9 9 9 9 7 9 9 10 0 7 14 13 14 0 1 2
34 14 13 11 9 10 9 9 0 2 14 13 15 9 7 9 3 7 3 2 7 13 15 0 2 9 2 14 13 10 9 1 10 9 2
7 0 1 9 2 13 9 2
34 1 9 15 14 13 0 1 9 10 12 9 13 14 11 7 14 11 2 11 14 11 2 11 11 2 11 14 11 11 7 11 14 11 2
10 13 10 9 16 13 1 9 0 1 2
16 1 9 2 14 0 10 9 14 13 1 9 1 7 10 9 2
41 8 9 2 9 14 9 1 9 1 9 9 1 8 2 13 9 3 0 1 9 9 2 8 2 2 13 9 1 9 9 9 0 8 7 1 9 8 1 11 9 2
66 8 1 10 9 0 2 13 15 1 10 9 7 13 10 9 1 7 10 9 1 2 7 13 15 0 1 10 9 7 1 10 9 2 7 0 7 0 1 10 9 2 14 13 0 1 9 9 10 9 10 7 14 13 1 9 1 9 1 9 15 1 9 10 9 10 2
18 14 13 1 16 9 9 1 9 14 13 15 1 9 9 1 9 11 2
15 2 14 13 15 1 15 16 9 7 9 1 9 1 9 2
16 9 9 14 13 1 7 15 0 7 15 1 9 1 9 9 2
17 13 10 9 1 12 2 7 13 11 7 11 1 9 1 3 0 2
5 13 15 1 9 2
30 13 15 9 7 9 1 9 16 13 15 0 14 9 1 9 15 2 13 2 13 0 10 9 15 16 13 3 1 15 2
44 13 10 9 10 1 9 1 10 9 1 1 9 0 0 9 13 0 14 0 1 13 10 9 0 7 9 9 1 9 10 9 15 11 7 13 10 9 1 10 9 0 15 11 2
10 13 15 9 16 14 13 15 1 9 2
6 13 1 15 13 3 2
22 1 15 2 13 10 9 9 1 12 9 1 2 9 1 9 2 9 2 9 7 9 2
7 2 9 1 2 14 11 2
21 13 9 0 1 9 10 3 2 10 9 0 1 11 10 9 16 1 9 9 9 2
151 8 13 10 9 10 9 9 7 10 9 2 16 1 1 2 1 9 14 13 1 14 9 1 9 8 7 16 0 1 1 10 9 10 14 13 10 9 9 7 10 9 1 14 13 10 9 9 10 1 9 1 9 14 13 1 9 14 13 1 9 2 14 13 9 9 1 9 7 1 9 14 9 1 9 10 9 9 7 10 9 10 1 9 1 2 10 9 7 10 9 13 9 1 10 9 1 9 14 0 2 13 10 9 2 1 9 2 14 9 16 13 10 9 9 14 13 10 9 7 10 9 8 1 9 1 10 9 7 1 10 9 14 13 1 15 1 9 8 9 1 10 9 1 9 1 9 1 10 9 10 2
32 13 0 9 9 9 3 14 13 10 9 1 9 9 10 9 11 2 1 9 1 9 10 9 0 10 2 13 12 9 9 1 2
23 16 16 14 13 1 9 3 13 9 1 2 7 13 15 15 13 15 2 0 1 9 9 2
21 14 13 15 1 15 13 1 9 1 9 10 9 7 10 9 1 9 7 1 9 2
14 13 10 9 2 10 9 7 10 9 1 9 1 9 2
9 2 13 3 10 9 13 0 1 2
33 13 1 11 8 1 11 11 14 13 9 9 9 10 9 10 1 10 9 10 12 9 16 15 1 9 1 9 10 9 9 14 9 2
9 11 9 1 2 2 13 2 2 2
18 16 13 10 9 1 7 13 15 9 0 16 14 13 15 10 9 3 2
26 13 10 9 1 10 9 14 13 10 9 0 1 9 1 12 9 1 9 2 1 9 1 10 9 10 2
20 13 0 1 9 16 1 9 3 13 9 10 9 0 1 10 9 1 10 9 2
16 1 10 9 2 13 0 10 9 10 14 9 1 9 9 9 2
41 15 15 10 2 9 2 2 10 9 0 13 0 16 13 10 9 3 2 9 0 9 16 14 13 9 9 2 7 9 9 2 9 10 9 2 16 10 9 1 9 2
20 13 15 1 9 1 11 14 0 1 9 0 7 13 15 15 10 12 9 1 2
16 8 2 13 10 9 1 14 13 11 11 14 0 1 9 10 2
5 13 10 9 15 2
28 1 9 12 9 14 9 1 9 1 10 9 10 2 14 13 10 9 12 9 1 9 10 9 14 13 9 1 2
59 2 11 14 14 13 1 10 9 14 9 1 11 2 16 13 15 1 9 1 11 1 9 14 9 2 7 13 10 9 1 10 9 14 13 15 9 1 9 11 7 14 13 9 1 15 1 10 9 14 9 1 9 11 16 13 11 11 11 2
26 14 13 10 9 9 0 1 10 9 2 16 13 0 1 10 9 14 9 14 13 9 1 9 1 9 2
80 8 10 9 14 13 1 9 8 13 15 1 9 10 11 1 9 3 0 16 13 9 15 1 10 9 7 16 13 10 9 1 8 3 1 9 7 9 14 13 10 9 10 1 9 10 9 14 13 1 9 10 9 10 1 9 13 10 9 8 1 9 1 9 15 16 13 15 1 9 1 9 9 14 13 1 15 1 9 8 2
8 9 11 1 9 1 12 9 2
23 13 10 9 14 9 9 3 3 10 9 1 14 13 10 9 8 1 9 1 10 9 0 2
23 1 9 9 1 9 10 14 13 1 9 1 9 0 10 9 2 13 9 0 0 1 11 2
8 13 1 3 1 9 10 9 2
37 13 9 15 15 1 10 9 14 13 11 1 9 1 9 11 9 3 1 10 9 15 16 10 9 1 9 2 10 9 9 14 13 1 11 15 2 2
23 2 14 13 9 16 13 9 1 9 0 9 14 9 1 10 9 2 2 13 10 9 11 2
3 11 11 2
36 16 13 10 9 1 14 13 10 9 2 14 13 15 3 1 9 1 10 9 1 9 10 9 9 7 14 13 10 9 1 1 9 3 1 9 2
17 9 2 1 9 0 0 13 10 9 1 9 9 7 9 1 8 2
5 13 0 10 9 2
8 14 13 15 10 9 1 11 2
44 16 13 15 1 1 13 9 1 2 13 9 1 14 13 15 1 9 11 2 11 2 1 11 2 16 13 1 9 15 14 13 15 14 1 9 7 1 9 10 9 14 13 15 2
7 14 13 9 16 13 15 2
26 1 9 2 13 9 1 14 13 16 14 0 1 10 9 2 7 9 10 14 13 1 9 1 9 10 2
45 13 10 9 1 9 0 2 12 1 11 9 9 2 12 1 11 11 2 12 1 9 9 7 9 2 1 10 9 9 2 2 12 1 9 9 7 9 9 7 12 1 9 10 11 2
23 13 9 14 9 14 13 9 9 1 9 14 9 1 9 9 1 10 9 1 10 9 9 2
66 1 9 10 9 1 9 1 2 14 13 1 9 1 9 14 13 9 3 1 10 9 16 1 1 16 12 9 0 2 7 13 1 9 11 15 2 14 13 9 10 1 9 1 9 1 2 7 14 13 10 9 7 10 9 9 1 10 9 3 2 7 1 1 9 1 2
14 1 9 13 10 9 0 0 1 10 9 10 14 0 2
6 13 15 9 10 9 2
21 13 15 3 1 9 0 16 14 13 1 9 9 7 9 1 9 1 1 10 9 2
13 2 1 9 1 9 10 9 9 2 2 14 13 2
35 13 9 1 1 9 3 12 2 13 9 1 9 3 1 9 11 7 2 16 14 13 2 9 0 11 14 11 3 1 9 1 10 9 0 2
6 13 11 3 1 9 2
10 1 9 14 12 14 13 15 1 9 2
7 2 13 9 0 3 1 2
7 9 0 0 14 13 1 2
89 8 14 13 10 9 9 1 9 1 10 9 1 9 14 13 1 9 8 16 13 7 1 14 13 9 9 1 1 9 1 9 0 14 13 1 10 9 14 9 1 9 1 10 9 7 9 1 9 9 13 14 13 10 9 0 14 9 1 10 9 16 16 13 9 1 9 10 9 8 14 13 10 9 10 10 9 1 9 0 10 9 7 14 14 13 1 10 9 2
7 13 9 0 1 10 9 2
24 1 9 11 13 15 1 9 1 9 10 11 2 1 9 11 2 1 9 11 7 1 9 11 2
75 13 11 2 12 2 14 13 10 9 10 9 14 9 1 9 1 2 9 2 2 7 3 0 7 14 13 1 10 9 9 14 13 9 1 10 9 7 1 9 9 1 2 13 15 0 2 16 15 2 9 14 9 1 9 1 10 9 1 9 10 9 14 13 1 9 1 9 10 9 1 9 13 3 2 2
19 2 13 15 1 9 10 9 2 7 13 10 9 1 1 7 13 9 1 2
22 2 16 13 15 10 9 3 13 9 1 2 13 15 1 9 1 9 2 14 13 9 2
9 14 13 9 7 14 13 9 15 2
12 13 15 10 9 7 10 9 14 13 10 9 2
12 13 9 1 9 14 13 9 0 1 9 1 2
36 13 9 0 1 9 8 9 9 7 9 16 14 13 10 9 3 10 9 1 15 1 12 9 10 2 9 0 14 9 7 9 14 13 1 3 2
26 11 1 10 9 14 13 9 9 1 9 1 9 0 2 16 3 2 13 0 7 9 15 9 10 9 2
29 14 13 15 16 3 7 9 1 9 2 7 9 9 9 9 0 2 16 14 13 15 9 0 14 13 1 9 3 2
23 2 13 15 10 9 3 3 1 10 9 7 14 13 15 10 9 1 9 2 9 7 9 2
83 10 9 2 0 2 7 10 9 2 0 2 2 13 15 9 10 9 10 9 2 10 9 7 10 9 2 13 15 10 9 7 10 9 9 10 9 2 13 10 9 2 14 13 0 1 9 2 1 9 14 9 1 10 9 1 15 14 9 2 13 10 9 2 14 13 0 1 9 7 14 13 3 1 10 9 2 10 9 7 15 1 9 2
15 13 9 3 1 10 9 14 13 1 10 9 0 1 9 2
7 13 9 0 15 1 9 2
3 9 9 2
14 16 3 7 3 13 15 1 9 14 14 13 14 9 2
22 1 9 13 10 9 7 10 9 0 2 13 9 14 13 1 10 9 16 10 9 0 2
