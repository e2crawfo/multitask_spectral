4798 11
9 0 9 1 1 9 0 13 13 2
5 9 2 9 9 0
15 9 13 16 0 13 0 9 1 1 9 0 14 13 13 2
16 1 9 0 2 0 1 12 9 9 1 9 9 9 9 13 2
34 7 9 3 10 9 14 3 13 13 7 3 1 9 9 2 9 7 9 16 15 1 9 9 15 13 2 0 1 9 10 9 13 13 2
15 3 9 13 16 10 9 1 9 9 9 1 9 13 13 2
33 1 0 9 1 9 0 16 9 3 3 0 1 9 0 9 13 2 7 9 9 14 13 16 1 9 15 1 12 9 0 13 13 2
16 1 1 10 9 2 9 0 10 9 2 9 15 14 0 13 2
24 16 10 9 0 9 13 13 2 9 15 13 1 9 9 7 9 0 9 0 1 9 9 13 2
13 9 10 9 1 9 0 9 9 1 9 13 13 2
5 9 2 9 0 9
16 9 0 9 13 1 9 9 9 7 0 9 9 9 9 13 2
37 1 9 9 0 9 1 9 2 9 9 13 2 9 0 9 13 13 9 0 1 9 0 0 1 9 9 7 9 10 9 1 9 9 2 0 13 2
38 10 9 13 2 10 12 9 9 9 9 16 9 9 0 1 12 9 9 9 1 9 13 7 1 9 9 13 0 1 9 0 14 3 9 9 9 13 2
11 9 0 1 9 4 1 9 9 9 13 2
5 9 2 9 0 9
19 9 1 9 9 1 9 0 1 9 2 0 1 9 0 1 9 0 13 2
29 1 9 9 1 9 2 9 12 1 9 9 13 2 9 0 0 1 9 0 9 9 1 9 9 9 0 9 13 2
48 9 1 9 7 9 9 9 0 1 9 9 9 0 7 9 1 10 9 13 16 9 3 0 9 9 9 16 1 9 1 9 9 9 9 13 2 1 9 9 0 1 9 10 9 16 9 13 2
23 1 9 9 2 9 1 9 0 9 9 3 1 9 9 1 9 9 9 0 9 13 13 2
3 9 9 9
8 9 9 9 9 9 0 13 2
29 1 10 7 4 9 0 10 9 14 9 13 7 1 15 9 13 2 4 9 15 14 0 9 0 7 9 0 13 2
14 9 9 13 16 9 9 14 1 9 7 9 9 13 2
17 9 0 15 2 9 1 9 0 2 0 7 9 1 10 9 13 2
22 9 9 2 9 2 9 2 9 7 9 1 9 1 9 9 1 9 9 1 9 13 2
16 1 0 9 9 15 1 9 9 0 0 1 9 9 15 13 2
13 9 15 9 9 13 7 9 9 9 1 15 3 2
13 9 1 9 12 1 9 15 1 9 9 9 13 2
15 1 9 1 9 1 9 9 0 1 9 9 9 0 13 2
31 9 9 1 10 9 3 1 9 0 1 9 15 1 9 13 7 1 9 1 15 1 9 2 0 9 9 9 2 9 13 2
11 1 9 1 9 9 9 9 0 9 13 2
31 3 10 9 1 9 10 9 0 15 13 16 1 9 9 2 9 0 1 9 7 9 9 15 2 16 1 9 9 9 13 2
28 9 0 9 1 9 9 0 14 1 9 13 16 1 15 9 0 2 9 0 7 9 0 1 9 0 9 13 2
21 9 9 1 9 9 9 7 9 16 13 7 1 9 0 2 9 9 2 9 13 2
20 9 0 1 9 9 9 7 9 0 9 1 9 9 9 0 7 0 9 13 2
35 9 1 9 15 9 7 9 9 14 1 9 9 0 7 0 9 9 15 9 13 7 9 14 1 9 13 16 3 1 9 9 15 0 13 2
26 9 0 7 1 10 9 0 9 2 1 9 0 9 9 13 7 9 0 1 9 9 15 14 9 13 2
45 1 9 9 15 9 13 9 13 2 9 7 9 13 9 13 2 9 9 1 9 13 7 3 2 9 1 9 9 7 9 13 13 2 7 9 1 9 0 1 9 7 0 9 13 2
28 16 9 9 0 0 9 0 13 2 9 9 15 2 9 7 9 9 7 9 15 9 1 9 1 9 15 13 2
31 9 9 0 7 1 10 9 0 2 1 9 7 9 9 0 9 0 9 15 14 9 13 7 9 0 1 9 10 9 13 2
25 9 7 9 9 16 1 9 9 13 2 9 0 15 14 13 7 1 9 0 15 1 12 9 13 2
20 9 3 13 1 9 9 15 9 13 7 9 14 13 16 3 0 9 15 13 2
27 3 15 1 0 9 13 16 0 13 13 16 1 9 2 9 7 9 9 9 0 7 1 9 9 0 13 2
16 9 3 9 13 13 16 9 9 0 1 9 9 7 9 13 2
45 7 3 0 13 16 9 15 14 1 9 0 9 13 7 1 10 9 1 1 9 15 9 0 14 9 13 2 1 9 0 7 0 1 9 13 1 9 0 2 0 7 0 1 9 2
33 9 3 1 1 15 13 16 1 3 13 9 0 15 14 9 1 9 13 7 3 3 9 7 9 16 1 9 10 9 9 13 13 2
35 9 3 9 13 9 9 9 15 13 2 1 9 9 13 7 3 7 13 9 15 14 1 9 0 9 13 2 1 9 9 1 9 0 13 2
23 3 16 9 9 16 13 9 9 0 1 9 2 9 7 9 15 13 2 1 9 9 13 2
20 7 1 9 9 7 9 4 13 9 12 1 9 0 9 0 1 9 9 13 2
18 9 0 9 7 9 0 15 2 3 1 9 3 0 15 3 0 13 2
15 9 1 1 15 13 16 9 14 13 16 3 9 13 13 2
13 1 10 9 2 3 1 1 9 1 9 0 13 2
11 15 1 1 9 0 1 9 0 9 13 2
14 9 0 1 9 9 2 9 9 0 1 9 15 13 2
26 15 3 13 13 1 9 9 1 9 0 1 9 9 15 2 9 13 16 1 9 9 9 9 9 13 2
5 9 0 9 9 9
6 9 1 9 13 13 2
6 9 9 1 9 13 2
10 9 2 9 2 9 2 3 15 13 2
5 9 2 9 13 2
6 9 1 9 9 13 2
11 9 2 9 9 13 2 9 15 3 13 2
20 9 1 9 9 14 1 9 13 2 9 0 13 2 9 14 1 9 0 13 2
21 1 9 7 9 7 9 1 9 13 2 1 9 0 9 13 7 1 9 13 13 2
3 3 13 2
8 9 2 3 3 0 15 13 2
7 9 15 3 13 2 6 2
15 9 2 2 9 14 13 2 13 3 15 13 9 2 13 2
10 9 1 9 0 13 7 3 9 13 2
34 9 2 3 3 15 13 2 1 9 9 13 2 9 9 13 1 9 2 7 1 13 9 7 9 13 7 9 13 3 15 13 2 6 2
5 1 9 9 13 2
19 9 2 0 7 1 9 7 9 14 9 13 2 2 9 0 16 9 13 2
6 9 13 7 9 13 2
12 9 2 6 2 6 2 9 15 13 13 9 2
7 3 3 13 13 0 13 2
2 6 2
12 2 9 13 2 13 9 15 4 12 9 13 2
18 2 7 0 9 13 2 9 9 14 1 9 13 2 7 1 15 13 2
23 1 9 2 9 16 9 9 13 7 1 9 1 9 13 13 7 3 9 14 13 2 13 2
12 2 9 9 1 9 9 1 9 7 9 13 2
16 1 9 15 1 9 9 15 14 1 13 7 1 15 9 13 2
6 9 1 9 13 13 2
16 9 9 7 9 0 2 0 9 2 9 1 9 0 9 13 2
4 9 9 13 2
6 9 1 1 9 13 2
9 9 2 9 15 4 12 9 13 2
10 9 2 3 9 13 2 1 9 13 2
7 2 9 9 14 13 2 2
3 3 13 2
12 9 2 3 9 2 2 3 9 15 9 13 2
8 9 2 3 2 9 9 13 2
13 9 16 3 1 9 13 2 0 13 1 9 15 2
5 9 2 9 13 2
3 9 13 2
10 6 2 2 9 1 13 2 9 13 2
16 9 16 1 9 9 9 13 2 15 14 1 10 9 9 13 2
5 9 2 9 2 2
14 9 3 13 7 9 0 2 7 0 15 2 0 13 2
5 9 1 9 13 2
11 9 9 15 14 9 13 7 3 0 13 2
9 9 2 9 2 12 9 9 13 2
16 9 1 9 9 1 9 7 9 14 1 9 0 13 2 13 2
18 9 1 9 7 1 9 9 13 2 9 13 9 9 15 14 0 13 2
9 9 0 13 7 1 3 0 13 2
36 9 2 3 13 9 15 13 2 3 9 0 13 2 15 9 15 13 1 15 13 2 9 14 1 9 15 0 13 2 13 2 9 9 9 15 2
8 10 3 13 13 1 9 15 2
8 9 2 2 13 2 1 9 2
8 9 14 1 9 1 9 13 2
9 9 2 9 16 3 13 10 9 2
2 3 2
6 7 1 9 9 3 2
7 9 1 1 9 9 13 2
9 9 2 1 9 13 9 15 13 2
7 2 9 16 0 13 2 2
2 13 2
18 9 1 9 9 9 1 9 9 7 9 3 0 7 9 15 2 13 2
8 3 1 9 13 7 9 13 2
9 9 12 9 9 15 14 9 13 2
11 1 10 9 13 7 9 14 1 9 13 2
16 2 1 9 9 0 9 2 1 9 9 1 9 9 13 2 2
4 9 9 13 2
7 12 9 15 14 0 13 2
21 1 1 9 9 13 1 2 9 2 9 2 9 2 7 9 15 9 9 0 13 2
8 9 14 13 7 9 9 13 2
6 15 14 1 9 13 2
7 9 2 9 9 3 13 2
28 9 9 2 2 1 9 7 1 9 9 13 2 9 15 2 9 7 2 9 9 9 9 1 9 14 9 13 2
8 9 0 13 7 3 9 13 2
13 9 2 2 1 9 7 3 13 2 9 13 2 2
3 3 0 2
9 9 9 9 9 14 1 9 13 2
14 1 9 15 2 9 9 9 2 7 9 9 0 13 2
12 9 9 13 7 9 9 15 13 7 9 13 2
9 9 1 9 7 9 9 14 13 2
7 9 2 13 15 9 13 2
6 9 2 15 9 13 2
4 9 13 9 2
13 9 9 1 9 9 16 1 15 9 9 13 13 2
12 0 9 1 9 1 1 9 7 9 9 13 2
13 2 9 0 9 2 9 2 15 13 9 2 13 2
6 0 2 15 13 6 2
28 9 2 16 9 9 0 13 13 2 7 1 9 9 13 2 9 9 13 13 2 2 9 9 1 9 13 2 2
4 9 2 13 2
22 9 9 0 13 7 9 9 9 15 13 7 1 9 9 7 9 9 9 1 9 13 2
10 9 1 1 9 9 2 1 9 13 2
3 9 13 2
4 9 3 13 2
25 9 16 9 9 14 0 13 7 13 2 2 9 9 1 9 13 2 9 9 14 1 1 9 13 2
23 9 9 9 14 0 13 7 13 2 2 9 9 1 9 13 2 9 9 9 14 0 13 2
16 9 12 14 0 13 7 13 2 2 9 9 1 9 13 2 2
8 9 9 14 9 13 7 13 2
17 9 1 9 1 1 9 7 9 9 16 1 15 13 2 13 13 2
8 12 1 9 9 15 14 13 2
11 9 9 13 7 9 13 1 9 9 13 2
5 9 2 9 9 2
5 9 9 0 13 2
14 16 15 13 1 9 9 13 4 9 0 14 0 13 2
12 9 13 3 9 13 16 7 9 13 0 13 2
13 15 13 16 9 9 14 1 9 0 3 13 7 2
18 9 9 2 0 9 9 1 9 9 13 13 7 1 9 9 9 13 2
9 9 2 1 9 2 2 9 13 2
6 9 2 9 9 13 2
13 2 7 9 14 1 15 13 2 9 2 0 13 2
9 9 2 2 1 9 2 0 13 2
7 9 9 14 1 9 13 2
7 9 9 14 1 9 13 2
10 9 15 9 14 13 7 3 9 13 2
11 9 9 9 9 2 9 14 1 15 13 2
10 9 9 15 14 1 9 3 13 13 2
6 9 1 9 0 13 2
7 9 9 14 13 1 9 2
9 9 9 9 14 1 9 0 13 2
12 9 9 9 9 0 1 9 1 9 15 13 2
8 9 9 14 1 9 9 13 2
8 12 12 9 9 1 9 13 2
9 9 0 13 9 13 2 3 13 2
11 9 9 1 15 13 7 9 15 0 13 2
6 9 9 1 9 13 2
15 7 9 9 9 14 0 13 2 7 1 1 15 9 13 2
4 9 3 13 2
4 9 2 9 2
22 2 9 3 1 9 0 13 7 9 15 14 13 2 7 1 9 9 1 9 13 2 2
11 9 9 9 15 14 13 7 1 9 13 2
5 13 2 0 9 2
9 9 1 15 9 13 16 2 13 2
6 9 9 2 9 9 2
6 9 1 9 0 13 2
8 9 14 3 13 7 0 13 2
18 9 9 1 9 13 2 7 3 9 15 9 14 1 9 13 7 13 2
2 13 2
3 9 9 2
9 9 9 1 9 7 9 13 13 2
10 9 9 14 13 7 3 1 15 13 2
11 9 14 1 9 9 13 2 1 9 13 2
9 15 0 1 9 9 16 9 13 2
9 9 1 9 0 1 9 9 13 2
4 9 9 2 2
5 1 15 9 13 2
11 1 9 9 13 16 1 9 9 0 13 2
22 9 15 14 0 1 9 13 7 15 15 16 15 7 9 1 9 0 15 14 9 13 2
15 9 1 10 9 0 13 16 4 1 15 9 9 0 13 2
18 9 0 9 15 14 9 13 16 9 14 1 3 1 1 9 15 13 2
20 9 9 13 3 15 14 3 13 16 1 9 13 7 3 1 9 0 0 13 2
21 7 15 15 16 13 12 9 7 9 7 9 9 16 12 9 7 1 9 15 7 2
19 9 1 9 9 13 2 2 9 9 1 9 13 2 9 15 14 9 13 2
23 1 9 9 13 16 1 9 1 9 9 9 0 13 2 1 9 16 1 9 1 9 13 2
11 9 1 9 9 13 2 15 14 9 13 2
6 9 15 9 13 13 2
14 1 12 9 2 1 9 0 2 9 9 14 0 13 2
7 9 9 15 14 0 13 2
6 9 3 9 1 9 2
11 2 9 1 9 0 15 14 9 13 2 2
20 9 3 9 1 9 13 2 1 10 9 9 14 9 13 16 3 0 9 13 2
6 2 9 9 13 2 2
17 9 1 2 9 9 1 9 13 2 1 1 9 9 2 9 13 2
18 9 13 7 0 1 9 16 13 9 13 2 9 9 14 1 9 13 2
4 9 2 9 2
4 9 9 13 2
12 9 1 9 9 9 2 9 13 2 9 13 2
24 9 1 0 9 9 1 9 13 13 7 1 9 0 13 2 16 9 13 10 9 14 0 13 2
20 9 1 9 9 13 7 0 2 3 7 3 0 9 0 9 13 2 9 13 2
10 9 9 15 3 1 9 16 9 13 2
5 9 1 15 13 2
7 9 0 13 7 9 13 2
5 13 9 2 15 2
5 3 1 9 13 2
6 9 9 1 9 13 2
2 13 2
7 9 2 9 9 2 9 2
4 9 2 13 2
10 9 2 9 13 1 10 9 9 13 2
14 9 3 9 13 7 3 0 9 13 7 0 9 15 2
4 9 2 3 2
2 6 2
6 16 13 2 9 13 2
5 1 9 9 13 2
17 7 1 9 9 1 9 1 9 7 3 9 13 9 1 15 13 2
5 13 13 2 3 2
4 9 9 13 2
5 9 2 9 9 2
9 9 15 14 9 13 7 9 13 2
7 9 2 13 2 9 13 2
9 9 3 9 13 7 0 9 13 2
6 9 2 9 13 9 2
35 1 9 15 2 2 3 15 15 14 0 7 0 13 7 0 1 9 9 13 16 2 16 13 13 3 15 7 4 9 2 9 13 2 9 2
18 15 1 9 16 3 13 1 15 9 9 13 2 12 1 12 9 13 2
6 9 1 9 15 13 2
7 9 2 0 3 13 9 2
6 12 9 0 9 13 2
9 9 2 1 9 9 2 9 13 2
14 9 1 9 9 2 9 9 1 9 15 1 9 13 2
7 9 9 14 1 9 13 2
13 9 15 1 15 2 15 3 2 1 9 3 13 2
11 9 7 9 15 9 1 1 15 9 13 2
13 1 9 9 13 7 3 9 15 1 15 0 13 2
18 9 10 9 15 0 9 9 13 16 3 10 9 9 1 9 9 13 2
9 9 2 2 16 13 2 2 6 2
5 9 15 3 13 2
3 9 13 2
9 9 16 1 9 0 13 13 13 2
4 9 3 13 2
15 9 2 2 0 7 1 9 9 3 3 2 4 9 13 2
9 9 13 2 9 9 16 9 13 2
2 9 2
14 7 1 9 7 9 15 14 13 2 1 15 9 13 2
8 9 0 3 9 15 14 13 2
19 2 1 9 1 9 9 2 7 15 14 1 9 9 9 13 7 9 13 2
17 15 1 9 9 13 2 9 15 14 1 9 9 13 7 9 13 2
4 9 3 13 2
27 9 16 1 9 15 2 3 2 9 13 7 15 14 0 13 2 3 9 9 9 14 1 9 1 9 13 2
3 9 13 2
7 9 14 1 9 15 13 2
12 15 14 3 0 13 2 9 9 1 9 13 2
7 9 14 13 7 3 13 2
6 9 1 9 3 13 2
6 9 15 14 0 13 2
9 9 13 7 3 9 1 9 13 2
13 9 9 14 13 7 1 9 9 9 13 7 13 2
7 9 2 2 9 2 13 2
5 3 1 9 13 2
14 1 9 9 13 2 16 3 9 15 1 9 9 13 2
14 7 9 9 3 1 9 0 15 1 9 2 9 13 2
19 9 16 9 13 2 9 1 9 13 1 9 1 9 2 9 1 9 13 2
18 9 9 13 16 2 3 13 2 2 3 9 14 1 9 0 13 2 2
17 9 9 9 0 13 7 9 14 13 16 1 9 9 3 3 13 2
19 9 0 1 9 13 2 9 13 7 3 1 9 13 7 15 14 9 13 2
6 9 9 9 9 13 2
18 9 3 13 7 3 7 1 9 15 13 15 14 9 13 7 9 13 2
10 9 3 1 9 9 9 14 9 13 2
50 9 0 13 2 1 9 15 16 9 13 7 3 1 1 15 13 7 0 13 2 7 2 9 1 9 15 13 13 2 7 1 9 7 1 9 2 1 9 2 13 3 9 15 14 9 13 7 9 13 2
10 9 9 1 1 9 15 1 9 13 2
15 9 1 9 9 0 13 13 7 15 14 1 9 15 13 2
4 9 9 13 2
4 9 9 13 2
9 9 9 14 1 9 0 13 13 2
7 9 9 3 13 7 13 2
11 9 1 9 0 13 7 9 9 9 13 2
11 9 9 14 13 7 13 7 1 9 13 2
20 9 9 9 14 1 9 1 9 9 13 2 9 9 14 1 9 1 9 13 2
8 9 1 9 7 1 9 13 2
13 9 2 2 1 9 2 16 9 13 2 9 13 2
7 9 2 3 15 0 13 2
8 9 2 3 15 16 0 13 2
17 9 2 2 1 0 9 2 0 13 2 7 9 13 2 9 13 2
7 9 9 14 1 9 13 2
22 9 1 9 9 9 9 1 9 13 2 9 1 9 13 13 16 9 14 1 9 13 2
19 9 1 9 7 9 14 0 7 0 0 13 2 7 9 14 1 15 13 2
14 9 2 2 1 9 2 9 9 2 9 13 3 9 2
10 9 2 10 9 14 9 13 2 9 2
26 9 1 9 7 1 9 9 14 9 13 2 9 1 9 13 7 13 16 10 9 9 2 1 9 13 2
27 9 3 12 12 2 1 9 2 15 9 14 9 13 16 0 7 0 13 2 7 9 1 9 13 1 9 2
6 9 2 6 2 9 2
8 9 9 9 9 1 9 13 2
7 13 1 9 9 14 13 2
5 9 16 3 13 2
7 9 2 3 9 9 13 2
14 15 15 13 2 3 9 0 13 16 1 9 0 13 2
16 9 2 2 1 9 2 3 2 3 2 13 9 16 13 13 2
22 2 7 15 1 9 0 13 2 9 9 13 13 1 9 2 1 9 2 9 1 9 2
10 9 1 9 15 9 13 7 0 13 2
3 9 13 2
21 9 2 9 9 2 9 9 9 13 2 9 9 0 16 13 1 2 0 9 13 2
10 9 2 9 9 2 9 9 9 13 2
6 13 15 15 9 13 2
11 7 15 15 14 3 3 13 1 9 9 2
15 9 9 1 9 9 2 7 9 2 9 2 1 9 9 2
12 9 9 1 12 9 7 9 1 9 0 13 2
13 9 14 1 9 2 7 9 9 14 1 9 13 2
9 9 1 9 9 13 9 14 13 2
26 9 2 2 1 9 9 9 2 9 9 2 15 9 15 0 13 9 2 1 9 9 13 9 0 13 2
9 9 1 9 13 13 7 0 13 2
21 9 16 3 9 13 2 9 15 1 0 9 2 1 3 2 9 14 0 15 13 2
14 9 2 13 9 2 13 9 15 3 13 2 9 15 2
6 3 13 9 13 9 2
18 9 2 2 1 9 7 1 9 9 13 2 6 2 3 9 13 6 2
15 2 1 9 2 6 2 16 13 13 2 9 1 9 13 2
26 9 9 15 14 1 9 2 16 9 9 13 2 9 13 2 9 1 9 13 7 9 0 15 0 13 2
11 9 1 9 9 0 9 1 9 9 13 2
10 9 0 9 9 13 7 1 9 13 2
16 9 1 9 15 9 13 7 1 9 0 13 7 1 9 13 2
12 9 9 9 7 9 3 2 1 15 9 13 2
6 9 9 1 9 13 2
15 9 1 9 2 9 13 2 13 13 7 9 15 9 13 2
12 3 9 3 0 13 7 9 15 1 9 13 2
21 9 0 13 2 9 15 1 9 9 16 1 9 13 13 2 1 1 9 9 13 2
7 9 2 3 15 13 9 2
3 3 13 2
6 9 1 9 15 13 2
8 9 1 9 9 14 1 13 2
13 2 9 14 13 2 9 2 9 2 3 13 9 2
18 9 0 9 13 7 10 9 9 15 1 9 13 7 15 14 9 13 2
7 9 2 1 9 9 13 2
6 9 0 13 7 13 2
6 9 3 1 15 13 2
10 9 2 2 0 1 9 2 3 13 2
9 9 9 9 13 7 3 1 9 2
6 9 2 3 3 9 2
6 9 3 9 13 13 2
6 9 1 1 9 13 2
18 9 15 1 9 9 13 7 0 9 13 16 1 9 1 9 9 13 2
15 9 1 9 13 7 9 0 2 7 9 15 2 0 13 2
17 9 9 9 14 13 7 9 0 9 9 2 15 14 0 9 13 2
10 9 2 3 13 3 13 2 9 13 2
9 2 9 2 13 3 13 2 9 2
8 2 9 2 3 9 9 13 2
15 9 1 9 13 7 1 9 1 15 9 13 16 9 13 2
10 9 9 2 9 13 2 3 13 9 2
7 9 9 13 7 9 13 2
14 9 0 9 13 1 9 9 2 9 1 9 9 13 2
7 2 16 13 9 13 2 2
27 9 2 3 9 13 7 9 13 9 14 13 2 9 9 9 9 14 1 13 7 3 9 13 2 9 13 2
24 9 1 9 9 15 14 1 9 15 13 7 9 9 14 16 3 9 15 14 13 2 1 13 2
7 9 2 3 15 13 3 2
9 2 9 2 9 9 13 1 9 2
5 13 3 13 9 2
4 9 9 13 2
15 9 2 9 13 2 9 13 9 1 15 13 13 2 9 2
14 16 1 9 9 16 13 9 13 2 13 16 0 13 2
4 9 13 9 2
8 9 2 3 3 13 3 13 2
8 9 9 9 2 9 14 13 2
6 9 9 14 0 13 2
6 9 1 9 0 13 2
6 9 15 0 9 13 2
8 9 9 0 1 9 13 13 2
10 9 2 3 2 13 9 2 3 13 2
12 9 2 3 2 9 2 13 2 1 15 13 2
17 1 9 9 9 13 2 16 7 9 0 13 9 2 9 2 13 2
14 9 9 14 2 16 0 9 9 0 15 13 2 13 2
10 9 2 2 1 9 2 9 0 13 2
4 9 0 13 2
14 13 9 2 9 0 13 7 9 1 9 15 0 13 2
5 9 2 3 9 2
15 9 1 9 9 9 13 7 9 9 14 16 0 13 13 2
6 9 2 6 2 6 2
8 2 3 1 15 2 12 13 2
9 9 9 9 14 13 7 0 13 2
10 9 9 9 14 13 7 1 9 13 2
31 10 9 1 9 9 9 13 13 7 3 9 7 9 16 1 15 9 13 13 2 1 9 9 2 1 9 1 9 9 13 2
9 9 1 9 9 2 9 7 9 2
28 3 13 16 3 9 9 13 7 3 13 16 10 9 13 13 2 3 9 13 7 10 9 14 13 1 9 13 2
20 9 13 16 1 9 1 9 9 0 9 9 9 9 1 9 9 0 9 13 2
13 7 3 3 10 9 3 3 1 9 15 16 13 2
57 3 9 1 9 15 14 9 0 1 15 0 13 13 7 12 2 12 9 9 0 16 13 13 16 1 9 9 13 7 10 9 0 9 13 13 16 9 0 9 9 16 10 9 14 9 9 13 7 15 16 13 7 9 1 9 13 2
18 9 1 3 9 9 13 7 15 3 9 14 9 13 16 1 9 13 2
28 16 9 9 13 2 9 3 0 1 9 13 2 16 9 16 1 9 0 13 9 13 2 15 16 1 9 0 2
18 10 9 16 9 15 14 3 13 2 1 9 7 9 9 0 0 13 2
21 7 16 0 9 13 7 9 14 9 13 2 13 16 3 2 1 10 9 16 13 2
11 15 1 9 9 9 1 9 0 0 13 2
24 3 2 16 0 9 13 2 3 9 13 7 13 9 13 2 1 9 9 9 7 9 9 2 2
19 1 15 2 9 16 1 9 13 2 1 12 9 9 0 9 13 1 9 2
18 0 1 15 7 1 10 9 1 9 9 16 3 1 9 1 9 13 2
44 9 9 7 9 13 2 9 7 9 0 1 9 13 16 15 15 15 9 9 9 0 13 16 0 1 9 16 13 2 13 9 3 0 13 2 3 9 9 9 1 9 9 13 2
69 1 15 1 9 9 13 7 9 0 13 16 1 12 9 0 13 7 15 7 10 9 15 13 1 9 0 15 2 9 7 9 2 16 9 9 9 13 2 15 15 9 13 16 16 15 0 9 13 1 15 13 7 13 16 9 3 0 13 16 3 9 13 16 10 9 13 1 12 2
53 1 10 9 2 1 9 9 7 9 9 9 13 7 1 10 9 13 16 9 2 9 7 9 2 14 1 10 9 9 13 2 2 15 13 3 9 14 9 13 7 16 1 15 9 13 2 13 1 10 9 9 13 2
31 2 1 0 2 16 13 1 3 1 10 9 9 13 2 3 9 13 16 4 13 13 7 9 13 3 1 9 15 9 13 2
38 3 13 13 16 1 9 13 16 9 1 10 9 1 15 15 13 2 7 9 9 15 1 9 2 1 9 7 15 9 9 3 0 9 0 7 0 13 2
16 1 9 7 9 10 10 9 12 9 0 1 9 9 9 13 2
54 16 0 10 9 13 2 12 9 1 12 9 9 3 13 16 9 7 9 0 9 15 3 9 9 3 9 0 10 12 13 2 9 0 7 9 0 7 9 0 2 16 15 15 15 14 1 9 13 16 3 9 3 13 2
20 10 9 12 1 0 9 13 16 9 13 13 2 16 3 15 1 9 0 13 2
37 13 1 9 10 9 3 13 2 7 3 1 9 1 9 7 9 9 2 16 9 9 7 9 9 16 9 15 3 16 0 1 15 13 2 0 13 2
53 13 16 1 10 9 13 1 10 9 16 1 9 0 13 2 16 0 9 13 7 13 16 9 9 3 9 0 7 9 0 13 2 7 9 9 15 1 9 9 9 13 2 13 13 10 9 3 9 1 9 9 13 2
67 15 9 0 14 1 10 9 9 13 16 16 0 9 13 7 13 1 9 2 1 10 9 16 9 13 7 13 10 9 14 9 13 2 1 9 15 9 13 1 9 2 1 9 2 9 7 9 0 2 9 0 2 7 9 2 16 15 15 1 12 9 13 2 9 0 9 2
17 16 13 9 0 9 14 9 13 2 13 16 9 0 9 9 13 2
23 16 13 9 0 9 9 14 9 13 2 13 16 15 1 9 0 3 9 9 9 15 13 2
19 15 3 9 13 16 10 9 3 9 9 15 13 7 3 9 9 0 15 2
8 15 9 13 16 15 9 13 2
28 3 9 0 9 1 9 2 9 0 9 1 9 9 1 9 2 9 0 9 1 1 9 0 9 7 9 7 2
17 15 9 13 16 15 9 0 13 13 16 10 9 0 9 15 13 2
40 1 9 7 16 3 9 0 14 9 13 2 13 16 3 9 0 9 13 2 10 9 14 15 9 13 16 13 16 15 3 15 14 1 9 7 9 9 13 2 2
10 9 15 15 13 16 15 0 9 13 2
33 15 1 12 9 0 9 13 13 9 9 13 0 9 16 1 10 9 13 9 13 2 7 13 1 0 7 0 0 0 14 9 13 2
41 1 12 9 0 13 3 3 10 9 3 9 16 10 9 4 1 13 16 15 14 1 9 9 13 7 13 15 13 2 16 9 7 9 7 9 13 2 3 3 13 2
7 3 9 9 7 9 13 2
46 1 12 9 0 2 9 1 15 13 16 13 10 9 1 9 9 9 7 9 9 1 9 7 9 7 9 15 0 12 10 9 1 9 13 2 16 3 15 13 2 3 3 15 4 13 2
11 3 9 0 9 16 9 1 0 9 13 2
5 3 3 15 13 2
4 9 16 13 2
4 9 7 9 2
12 15 16 13 9 9 13 2 3 13 9 13 2
2 3 2
14 3 1 9 15 7 9 7 9 15 1 9 9 13 2
26 15 14 3 1 9 13 16 3 9 10 9 10 9 13 7 9 9 15 15 9 13 7 3 9 3 2
12 9 7 9 2 9 3 15 14 13 13 3 2
10 3 9 14 16 13 2 13 1 9 2
29 9 9 1 9 16 9 13 0 0 13 2 9 16 9 13 9 13 7 13 2 1 9 0 15 13 1 10 9 2
12 15 13 1 12 9 0 1 15 9 13 13 2
17 7 15 9 13 16 15 1 9 0 13 7 9 13 3 0 13 2
19 16 15 16 9 14 1 9 13 7 7 9 7 3 2 9 7 9 14 2
46 1 3 16 9 9 13 7 9 13 2 1 15 15 0 13 1 9 7 15 9 7 9 15 7 9 16 1 9 9 12 10 9 1 15 9 13 7 12 10 9 14 16 1 15 13 2
15 1 3 2 1 12 9 0 9 16 0 13 7 7 0 2
17 16 9 0 14 9 13 2 16 1 9 9 0 9 16 9 13 2
12 16 9 9 0 7 0 16 13 7 9 9 2
33 15 1 9 9 7 9 12 9 0 2 4 13 2 9 16 13 0 13 7 1 1 9 0 3 13 1 9 7 9 15 9 13 2
17 1 15 2 9 0 15 14 9 13 1 9 1 9 9 7 9 2
8 7 9 14 3 1 15 13 2
27 13 15 16 9 13 2 3 9 13 9 9 14 9 1 9 13 16 0 13 2 9 13 9 9 15 13 2
27 15 16 10 9 16 1 9 2 9 7 7 1 1 9 7 10 9 0 13 2 3 9 1 15 9 13 2
17 9 13 1 9 9 1 10 9 9 13 7 13 9 0 9 13 2
8 9 0 7 9 3 9 13 2
84 3 2 16 1 9 0 13 2 1 3 9 9 9 0 13 7 1 3 9 13 13 2 7 16 9 0 10 9 0 14 1 9 13 2 9 16 13 3 1 9 9 9 1 9 13 7 13 2 10 9 1 9 9 13 2 10 9 1 9 9 16 9 15 1 15 15 13 2 9 13 16 3 1 9 9 15 9 13 7 1 9 13 13 2
26 15 13 13 15 14 1 9 0 0 13 2 1 9 16 9 1 15 9 13 7 16 13 9 0 13 2
20 10 9 13 16 9 13 2 9 15 1 9 0 9 0 13 2 16 9 13 2
11 16 1 9 9 9 0 14 1 9 13 2
33 16 13 1 9 9 9 13 16 3 3 13 16 9 7 9 9 0 13 7 15 7 3 13 1 9 13 16 12 10 9 16 13 2
19 16 13 9 14 9 13 2 9 13 1 10 9 9 9 15 1 9 13 2
14 9 2 15 15 14 9 13 3 16 9 9 13 13 2
16 16 15 9 13 16 15 13 13 16 9 1 9 13 7 3 2
17 9 16 3 1 9 9 1 15 13 15 13 16 15 3 9 13 2
12 13 9 15 15 13 16 9 13 9 9 13 2
8 16 13 16 15 0 9 13 2
23 9 2 9 7 9 2 7 9 15 9 0 13 16 3 3 7 1 9 0 1 9 13 2
21 7 15 13 0 9 13 16 9 9 2 13 9 13 16 1 3 3 9 13 13 2
58 16 9 9 13 9 16 1 9 15 13 7 9 13 7 9 4 15 14 9 13 7 9 10 9 15 14 13 2 3 3 9 9 14 13 2 16 9 14 13 2 9 14 16 13 7 9 9 14 16 13 2 9 1 9 9 0 13 2
19 3 15 13 1 9 0 15 9 7 9 12 9 0 1 9 14 9 13 2
20 3 15 16 9 0 16 9 16 15 14 13 2 9 13 7 16 15 13 3 2
10 9 13 1 9 2 9 15 13 2 2
43 10 9 15 13 1 9 15 7 9 9 7 9 9 9 9 9 9 13 2 7 16 9 0 13 2 1 9 9 0 15 2 16 12 9 0 1 9 13 2 15 13 15 2
14 15 13 0 9 12 13 7 3 9 13 1 9 9 2
8 15 13 13 9 9 15 13 2
15 9 15 13 10 9 13 2 7 13 2 15 16 9 9 2
23 3 16 9 9 9 7 9 9 0 13 2 3 9 1 15 7 13 13 16 4 3 13 2
16 9 16 3 9 4 13 2 9 16 9 9 7 9 4 13 2
49 1 15 7 13 2 12 9 13 9 9 15 9 13 2 1 15 7 13 13 9 15 9 10 0 13 2 12 9 13 16 9 9 16 9 9 9 3 1 9 9 0 13 2 9 9 0 9 15 2
7 3 13 3 10 9 13 2
19 15 1 9 9 0 7 0 13 16 9 4 13 2 1 15 7 15 13 2
13 9 15 9 13 16 9 14 13 7 13 9 15 2
11 3 2 3 7 3 2 9 9 0 13 2
8 9 9 1 10 9 0 13 2
7 9 9 13 16 9 13 2
12 3 9 1 9 1 9 15 15 0 9 13 2
27 7 9 16 1 9 9 7 9 0 13 15 13 16 9 9 13 9 14 13 7 9 14 15 15 9 13 2
18 3 9 9 0 13 1 9 9 2 7 15 1 9 15 15 0 13 2
15 0 9 15 15 13 16 9 9 1 1 9 15 3 13 2
28 3 1 10 9 16 15 13 2 15 15 7 9 13 15 9 9 9 14 3 9 15 13 13 16 9 9 13 2
30 3 9 9 9 13 7 13 16 15 9 0 9 0 15 15 14 13 13 16 1 9 15 13 9 7 9 1 9 13 2
10 7 3 9 15 14 13 7 0 13 2
18 13 10 12 16 16 13 0 13 2 7 15 9 15 14 0 0 13 2
5 15 13 9 13 2
19 9 13 16 9 15 9 13 9 0 13 7 3 9 13 7 9 0 13 2
17 3 9 9 16 9 13 9 9 14 13 13 7 1 15 9 13 2
17 15 10 9 13 16 15 1 9 0 0 13 9 13 7 9 13 2
17 3 16 10 9 9 13 10 9 0 15 13 1 10 9 7 9 2
23 3 15 4 9 14 13 16 9 13 7 16 1 12 9 9 0 9 13 2 3 9 13 2
21 3 1 1 9 15 10 9 13 2 15 9 0 13 2 9 7 9 0 9 13 2
14 3 16 0 7 0 13 7 3 7 9 14 0 13 2
21 7 13 13 1 1 9 16 9 13 9 9 0 13 2 0 9 13 7 9 13 2
6 3 1 15 9 13 2
8 9 0 15 10 9 0 13 2
14 16 1 9 16 13 0 9 0 3 13 2 9 13 2
21 10 9 16 16 9 15 15 14 1 9 9 9 9 13 2 1 10 9 9 13 2
22 16 15 1 9 3 9 7 9 9 13 2 15 15 14 4 9 13 1 10 9 9 2
7 9 13 15 9 0 13 2
34 9 13 9 0 13 7 16 9 9 14 9 13 2 4 1 10 9 7 9 7 1 10 9 9 13 16 9 15 15 14 4 9 13 2
21 12 9 15 15 15 14 13 0 1 9 2 1 15 7 9 15 14 1 15 13 2
23 12 9 16 13 2 9 15 15 4 13 2 1 3 15 4 1 10 9 15 9 0 13 2
10 1 9 9 9 1 9 3 9 13 2
14 16 3 15 7 15 13 9 16 1 10 9 9 13 2
19 15 16 13 16 9 0 9 1 10 9 9 13 7 9 9 16 10 9 2
39 9 9 2 9 0 9 0 9 2 16 3 9 9 9 13 2 3 9 13 2 9 0 9 0 2 9 9 7 9 9 12 9 9 16 3 3 9 13 2
25 1 9 15 2 9 2 15 9 7 10 9 16 9 9 0 14 9 13 2 3 4 9 15 13 2
29 12 1 9 10 9 13 16 15 13 2 9 15 9 13 2 9 15 9 1 9 7 9 1 9 7 9 15 13 2
14 9 16 9 9 9 13 7 9 0 1 15 0 13 2
20 1 0 9 0 13 2 7 15 9 1 9 9 7 9 9 1 9 0 13 2
32 9 13 16 9 13 16 10 9 7 9 9 13 1 9 10 9 0 0 2 7 9 16 13 15 13 16 9 9 9 9 13 2
18 0 1 15 7 1 10 9 7 9 9 0 9 3 3 16 0 13 2
18 10 10 9 1 9 9 13 7 3 16 1 9 7 9 1 9 13 2
13 1 1 9 16 1 10 9 13 1 15 9 13 2
14 10 9 3 1 10 9 16 9 9 13 15 9 13 2
26 3 12 1 9 1 9 0 9 12 9 9 0 13 7 12 1 15 1 12 1 9 15 12 9 13 2
38 1 12 9 15 1 15 9 13 2 3 7 3 9 1 15 9 13 7 9 9 1 10 9 1 9 0 13 2 16 3 1 9 15 15 14 0 13 2
44 9 0 13 15 9 9 15 14 9 13 7 9 13 16 9 7 9 15 14 1 9 9 9 0 9 13 13 7 15 1 9 13 13 7 16 9 1 9 13 1 9 9 13 2
15 9 9 9 13 7 13 15 13 15 14 1 9 9 13 2
17 7 9 16 0 13 7 9 1 9 13 7 15 1 15 9 13 2
42 9 15 1 9 10 9 14 13 7 9 13 7 13 16 9 15 1 10 9 13 7 3 13 7 15 14 0 13 2 9 16 12 9 1 9 0 13 2 13 1 9 2
6 1 10 9 3 13 2
24 7 3 12 1 9 16 9 9 0 13 13 15 13 16 15 9 0 14 1 9 10 9 13 2
9 10 9 16 9 1 9 9 13 2
29 1 10 9 16 0 0 13 2 9 9 15 1 9 1 15 13 2 9 7 9 16 9 0 1 9 9 15 13 2
12 16 3 9 13 9 15 1 9 15 0 13 2
17 0 9 0 13 2 3 1 9 9 7 15 9 0 1 9 13 2
22 9 13 16 9 13 7 13 9 0 13 2 7 15 9 1 9 9 7 9 9 13 2
15 9 13 1 9 9 13 2 7 15 9 10 9 14 13 2
11 1 10 9 15 9 15 1 9 9 13 2
24 9 9 9 1 9 0 9 1 9 9 9 13 7 7 9 9 7 9 9 9 9 7 2 2
21 9 9 2 9 9 2 1 10 9 12 9 13 1 9 9 13 7 13 1 9 2
11 9 16 15 10 9 14 13 9 0 13 2
26 1 12 9 16 0 7 0 3 13 2 9 16 1 9 1 9 15 2 0 13 2 13 7 9 13 2
40 3 1 15 7 9 14 0 13 2 13 13 16 9 15 1 9 10 9 2 16 13 7 9 9 1 1 10 9 1 9 2 3 9 2 9 7 9 3 13 2
14 16 15 10 9 14 1 9 12 9 0 1 9 13 2
8 16 0 13 15 3 0 13 2
7 9 15 3 9 16 13 2
16 1 15 3 0 13 16 9 13 7 9 13 7 9 16 13 2
29 16 9 1 15 9 0 13 2 3 9 13 16 10 9 14 9 13 2 1 15 7 9 13 2 16 9 9 13 2
16 3 9 1 10 9 12 9 9 0 16 13 2 9 13 13 2
9 9 9 9 16 1 15 0 13 2
28 15 13 9 15 3 0 13 7 9 1 15 7 9 15 1 12 9 0 0 1 9 12 9 1 15 0 13 2
42 12 1 9 0 15 2 16 3 9 16 13 1 9 9 9 2 1 15 7 0 13 1 9 9 2 15 13 16 1 9 0 16 9 1 15 9 0 13 2 9 13 2
24 1 9 9 2 15 9 15 1 12 9 16 3 4 9 9 13 2 0 7 0 7 0 13 2
34 1 9 15 7 9 7 9 13 7 7 9 13 7 7 10 9 14 16 13 9 13 2 13 1 9 15 1 9 1 9 0 9 13 2
8 16 9 12 9 9 0 13 2
7 3 15 0 9 9 13 2
52 12 1 9 16 15 13 1 9 1 9 2 3 15 1 15 9 13 2 7 15 1 9 9 0 9 13 2 15 13 16 1 10 9 16 13 13 10 9 9 13 2 3 13 13 13 3 13 3 9 15 13 2
4 9 13 2 2
5 9 2 15 13 2
26 10 10 9 1 9 2 9 9 7 9 9 13 2 12 9 16 3 13 2 13 3 0 13 16 13 2
30 16 12 9 9 1 0 9 9 13 7 13 1 9 9 9 9 16 9 13 13 7 1 10 9 13 2 13 7 13 2
6 16 1 9 9 13 2
15 0 9 16 1 15 9 13 2 3 13 10 9 13 13 2
38 9 9 9 13 15 0 13 1 10 9 1 15 9 13 2 3 9 0 7 0 7 0 13 2 10 9 1 12 9 13 2 10 9 1 9 15 13 2
21 7 9 9 9 3 13 15 0 13 1 9 0 9 15 13 2 7 9 9 9 2
18 12 1 9 0 9 15 9 9 13 2 1 9 15 9 3 0 13 2
29 15 1 9 9 9 2 12 9 9 13 13 16 9 9 1 15 13 13 7 16 9 13 2 7 1 9 9 0 2
46 3 9 16 15 13 1 1 15 9 0 13 16 1 9 9 0 13 2 12 9 1 9 15 9 0 16 13 9 1 15 15 0 13 2 0 13 7 12 9 9 14 13 1 9 9 2
7 7 1 9 9 0 13 2
38 3 0 13 1 0 9 16 1 9 9 13 7 3 9 13 16 9 9 13 16 0 13 7 3 9 9 14 0 13 7 3 12 9 13 7 9 13 2
8 15 1 9 9 3 9 13 2
23 1 1 15 1 9 15 12 9 9 13 7 9 14 9 13 7 13 10 9 1 9 13 2
13 1 1 10 9 16 13 16 9 9 15 15 13 2
19 3 1 9 9 9 7 9 9 9 15 13 2 7 9 14 15 15 13 2
28 9 15 15 13 16 1 10 9 12 9 3 0 7 0 1 9 13 7 15 7 9 0 13 1 10 9 13 2
5 3 1 15 13 2
16 0 9 16 9 4 1 3 13 2 16 15 13 10 9 13 2
16 1 10 9 13 13 3 9 13 2 13 3 10 9 9 13 2
52 13 3 10 9 13 16 15 13 2 16 9 3 1 9 10 9 13 16 9 16 13 9 13 2 1 9 10 9 13 9 2 13 3 9 13 2 3 9 13 16 1 15 9 9 1 9 9 13 2 3 3 2
31 3 10 9 0 7 10 9 14 16 13 0 13 2 12 9 1 9 1 9 0 7 0 2 3 1 9 10 9 14 13 2
15 3 1 12 9 9 1 10 9 2 10 9 9 9 13 2
31 3 9 9 13 0 13 2 7 16 3 1 9 9 13 7 12 9 0 2 3 12 9 1 9 10 9 7 9 9 13 2
9 15 10 12 9 9 14 16 13 2
19 15 12 9 1 9 9 14 10 9 13 7 9 15 14 1 9 9 13 2
19 12 9 16 13 1 1 9 9 0 13 16 1 9 9 0 9 9 13 2
7 1 1 9 3 9 13 2
22 12 9 0 16 1 10 9 13 7 3 9 13 13 13 2 9 7 9 10 9 13 2
7 10 9 9 3 0 13 2
63 9 16 0 1 9 9 13 13 7 9 1 15 9 13 13 2 1 9 1 10 9 13 13 7 1 9 15 15 3 9 13 13 2 3 9 15 9 7 9 16 1 15 1 9 9 13 7 1 15 1 9 12 9 16 13 7 15 1 9 9 9 13 2
7 12 9 9 9 3 13 2
22 12 9 9 0 13 2 16 1 9 9 0 16 9 9 14 1 12 9 0 0 13 2
23 15 15 15 9 13 1 0 9 0 16 9 14 13 2 3 13 7 13 7 9 14 13 2
16 7 1 9 0 12 9 13 16 3 9 9 9 7 9 13 2
10 13 13 16 15 3 1 10 9 13 2
27 16 1 9 13 7 3 2 9 14 3 13 7 9 14 3 7 15 14 9 13 7 1 12 9 0 13 2
13 7 15 7 10 9 9 9 7 9 1 9 13 2
15 10 9 14 16 15 13 15 12 9 13 2 9 7 9 2
40 1 9 1 9 9 3 3 9 13 2 9 16 9 13 1 12 9 2 12 9 15 3 2 9 13 2 15 14 1 12 9 13 2 2 16 9 14 0 13 2
19 13 13 9 1 9 0 13 7 10 10 9 14 9 9 13 16 9 13 2
27 7 1 9 0 9 14 13 2 16 3 4 13 9 10 9 10 9 15 9 12 12 9 1 15 0 13 2
26 1 9 13 13 16 9 16 1 10 9 1 9 9 13 1 9 16 3 1 9 13 2 3 0 13 2
16 1 15 3 9 13 16 10 9 4 1 9 0 3 0 13 2
35 15 16 13 9 1 1 9 13 2 15 9 7 0 7 7 0 13 2 9 13 2 13 2 9 0 2 7 15 9 0 7 1 10 9 2
5 15 3 0 13 2
14 9 16 3 9 3 0 7 3 0 7 3 0 13 2
11 15 10 9 14 1 9 13 2 3 9 2
9 9 9 10 9 1 9 9 13 2
16 10 9 3 9 13 7 15 1 9 13 3 7 3 9 13 2
13 12 9 1 9 9 16 1 9 9 0 9 13 2
32 15 1 12 9 13 10 9 16 4 9 13 7 1 12 9 13 2 1 12 9 13 9 9 14 13 3 2 9 9 0 13 2
23 1 10 9 2 9 13 16 4 15 14 1 9 3 13 7 13 15 9 0 14 9 13 2
7 4 1 9 0 9 13 2
22 16 15 9 0 13 2 15 9 1 9 9 13 2 7 1 9 9 10 9 9 13 2
16 3 1 9 13 16 9 9 0 0 15 13 16 9 0 13 2
41 1 9 0 2 15 13 1 10 9 0 13 7 0 13 2 7 13 13 10 9 9 2 9 9 0 14 1 3 13 7 16 9 15 14 1 9 9 13 7 3 2
14 9 13 9 15 16 9 10 9 14 1 9 9 13 2
18 9 15 0 13 3 9 15 9 0 7 0 13 7 15 3 0 13 2
31 10 9 16 1 9 15 0 13 7 10 9 12 9 0 1 15 0 13 2 9 12 9 0 13 2 9 2 9 7 2 2
62 15 3 1 15 13 12 9 9 16 9 7 9 7 1 10 9 13 1 3 9 1 12 1 9 0 9 13 2 7 16 13 1 9 0 15 2 15 15 0 1 10 9 13 2 1 9 2 16 15 10 9 14 13 13 1 9 7 1 15 13 9 2
7 7 9 14 13 9 13 2
15 1 10 9 2 15 9 13 16 3 9 9 9 9 13 2
29 15 9 13 1 10 12 2 12 9 12 9 12 9 14 9 13 16 9 0 15 3 0 13 2 7 0 9 13 2
28 3 1 9 15 1 9 0 15 2 9 16 9 13 7 9 15 13 2 0 9 13 2 1 9 9 0 13 2
20 15 15 14 1 9 16 13 0 13 7 1 9 7 9 16 9 1 9 13 2
12 9 9 2 3 1 1 9 9 9 9 13 2
20 15 9 0 15 13 16 1 9 9 9 9 13 2 16 9 0 15 9 13 2
21 0 9 13 16 9 13 7 9 13 16 1 10 9 3 9 13 7 3 0 13 2
21 1 10 9 9 16 4 13 15 13 16 9 0 0 0 13 13 1 9 9 13 2
31 3 13 16 15 0 9 1 15 14 1 9 0 1 9 7 9 7 2 0 12 9 0 13 13 7 1 10 9 9 13 2
24 15 13 9 9 3 13 2 16 3 1 0 9 9 13 2 1 10 9 16 1 9 0 13 2
40 15 16 1 9 9 9 7 2 7 9 13 13 16 10 9 4 1 10 9 10 9 16 13 13 2 16 9 9 3 13 7 16 1 10 9 15 9 13 13 2
26 15 12 9 13 7 4 15 9 1 9 15 13 16 9 9 13 2 16 1 10 9 9 14 9 13 2
15 9 9 9 0 1 0 9 9 13 2 3 9 0 13 2
19 1 10 9 9 14 1 13 7 9 15 15 14 1 9 9 0 9 13 2
20 3 10 9 16 1 15 9 13 2 3 1 9 15 9 13 7 3 9 13 2
20 3 9 1 9 15 9 0 13 7 16 10 9 1 9 9 13 7 7 0 2
20 9 0 9 16 1 9 0 13 7 9 15 15 13 16 13 7 0 15 13 2
36 15 9 13 1 10 9 7 10 9 12 10 9 0 13 7 0 16 13 7 12 10 9 0 16 13 16 15 15 1 9 13 7 0 16 13 2
38 1 9 15 9 15 0 13 2 16 13 9 0 15 15 14 13 2 7 9 9 0 13 7 15 14 16 1 0 9 9 13 2 7 1 12 9 0 2
19 15 4 9 13 16 16 15 0 15 13 7 7 10 9 1 9 15 13 2
13 10 9 9 13 16 15 16 9 13 9 15 13 2
50 3 9 13 9 13 1 10 9 16 3 1 15 9 13 2 16 16 9 13 2 10 9 1 9 13 2 9 0 9 0 2 9 9 2 16 3 3 2 15 1 3 9 7 9 9 13 2 9 13 2
6 9 9 1 9 13 2
14 9 0 15 1 15 9 13 7 13 10 9 14 13 2
19 3 1 15 9 13 2 13 10 9 9 9 13 2 13 9 14 9 13 2
13 16 1 10 9 0 9 14 1 9 9 15 13 2
28 9 9 16 3 9 13 2 1 9 9 9 0 2 1 9 0 13 7 9 13 7 13 15 1 9 9 13 2
13 9 9 1 9 9 7 9 9 15 15 9 13 2
36 10 9 9 13 7 13 3 14 9 13 2 10 9 3 9 9 2 9 7 9 3 9 14 0 9 7 9 13 7 15 9 13 9 0 13 2
33 15 13 1 15 9 13 7 13 16 10 9 14 13 0 13 2 7 15 0 13 7 10 9 16 0 13 2 13 3 0 2 13 2
14 9 9 2 9 9 2 16 3 9 0 13 16 13 2
24 1 9 9 10 9 3 0 13 7 9 15 14 13 7 3 13 16 9 15 9 15 16 13 2
7 9 9 16 3 9 13 2
20 9 9 0 1 9 2 9 0 1 1 9 9 0 1 9 1 9 13 13 2
36 9 2 12 2 9 13 16 9 9 0 1 12 12 9 13 2 7 9 0 9 3 0 14 1 1 9 9 2 9 9 12 9 2 9 13 2
40 0 9 1 1 9 1 9 0 1 9 13 13 2 9 16 3 9 0 1 1 15 16 16 9 3 10 3 16 9 13 1 9 13 7 3 2 9 13 13 2
22 0 1 3 9 9 9 9 9 0 0 13 1 9 9 9 12 9 0 0 13 13 2
22 9 0 15 13 16 0 13 9 3 9 13 16 9 0 14 3 0 1 9 9 13 2
33 9 9 9 0 9 2 9 13 16 9 3 0 1 9 0 14 9 13 16 9 0 1 9 2 9 7 9 16 0 0 13 13 2
19 9 0 16 1 9 12 1 9 9 13 2 10 9 9 14 9 13 13 2
29 9 2 9 7 9 2 12 2 9 13 16 9 9 0 9 0 2 9 7 9 13 16 1 9 0 16 0 13 2
43 1 15 3 2 9 9 1 15 9 13 16 9 9 0 14 4 1 9 3 9 9 1 9 3 7 0 9 0 13 2 9 2 12 2 9 2 12 2 9 2 12 2 2
26 10 9 1 9 1 9 9 9 3 9 0 2 0 2 0 7 3 1 9 9 0 7 9 0 13 2
38 9 0 9 0 1 1 9 9 0 15 13 16 15 0 9 13 1 9 7 0 1 9 9 13 1 1 9 2 9 2 12 2 9 9 2 12 2 2
20 10 9 1 9 9 9 9 7 9 9 9 13 2 9 7 15 2 12 2 2
18 10 9 0 1 10 9 0 0 2 9 0 1 9 0 1 9 13 2
22 9 9 0 9 0 13 1 9 1 9 7 9 0 0 2 3 9 9 7 9 9 2
24 9 16 9 0 9 0 13 1 9 16 0 9 9 13 2 9 0 13 7 0 7 0 13 2
15 1 9 9 9 3 0 1 9 9 0 2 0 4 13 2
18 9 0 1 1 9 0 9 9 9 13 16 9 1 9 15 9 13 2
47 9 0 1 9 9 3 0 9 9 9 7 9 13 7 3 0 10 9 9 0 2 0 1 9 0 7 0 2 9 0 2 9 9 2 9 7 9 0 13 2 9 2 9 2 12 2 2
36 1 9 9 9 9 2 12 2 2 2 9 7 9 3 1 1 9 0 3 13 16 3 9 9 0 0 13 7 3 12 9 9 9 9 13 2
11 3 9 13 0 1 15 3 1 9 13 2
32 9 0 1 3 9 13 1 9 2 9 2 9 9 7 9 2 3 9 0 7 9 0 16 3 9 1 15 0 1 15 13 2
27 2 9 0 1 1 9 9 0 2 9 7 9 0 14 16 9 9 9 7 9 9 13 2 0 13 13 2
30 1 9 0 2 10 9 9 12 9 9 0 14 0 13 13 16 9 13 1 2 0 2 2 0 2 7 2 0 2 2
16 9 2 0 2 0 9 0 7 0 9 1 9 14 9 13 2
38 9 9 2 0 2 9 9 9 0 13 2 1 9 7 9 9 1 9 9 0 7 9 9 0 9 13 2 9 2 12 2 12 2 9 2 12 2 2
23 10 9 0 1 9 1 1 9 0 1 9 16 9 13 13 2 9 2 12 2 12 2 2
37 1 10 9 2 9 0 1 9 0 13 2 1 10 9 16 3 0 9 0 9 1 9 9 0 13 2 9 7 9 2 12 2 9 2 12 2 2
32 7 9 0 13 2 9 9 2 12 2 7 1 1 9 9 1 9 9 0 1 9 9 0 13 2 9 2 9 2 12 2 2
16 1 10 9 2 9 0 9 9 0 2 9 0 2 9 13 2
29 9 2 12 2 9 13 16 9 2 0 2 1 9 12 9 7 9 0 9 12 9 1 9 9 0 14 9 13 2
24 9 2 0 2 1 9 0 9 9 9 3 7 3 0 13 7 1 10 9 0 16 9 13 2
21 10 9 0 9 9 0 9 13 7 1 9 9 0 9 7 9 0 9 9 13 2
24 9 2 0 2 16 9 13 16 1 9 13 3 9 1 9 13 7 7 9 16 3 0 13 2
26 15 0 1 9 16 9 9 13 9 13 7 1 9 0 16 9 9 7 9 0 14 13 2 9 13 2
16 10 9 3 0 1 9 2 0 2 0 13 7 9 0 13 2
36 1 1 9 9 2 15 9 0 14 1 9 9 9 0 7 1 9 9 16 1 1 9 0 7 9 7 9 9 0 7 0 13 2 9 13 2
35 9 0 1 9 1 9 9 1 9 9 9 9 7 9 9 9 12 9 13 13 2 3 9 9 9 1 9 9 0 1 9 9 9 13 2
19 9 9 9 1 0 9 10 9 1 9 9 2 1 9 9 0 13 13 2
19 9 0 9 9 9 3 0 13 2 9 9 12 12 12 1 12 12 9 2
16 1 1 9 9 9 9 10 9 0 13 16 9 15 0 13 2
14 9 0 9 9 9 7 9 3 7 0 9 9 13 2
27 1 9 10 9 4 1 9 2 9 2 1 9 9 9 9 7 2 9 2 1 9 9 9 9 9 13 2
11 0 9 0 9 1 9 9 9 13 13 2
20 1 9 12 3 9 9 9 12 2 12 9 9 1 9 9 9 9 9 13 2
28 12 9 1 0 10 9 13 1 2 2 9 0 2 1 9 9 9 7 9 9 1 9 9 9 1 9 12 2
36 9 9 1 9 0 1 12 12 9 13 2 1 9 7 2 9 2 9 0 2 1 9 12 7 12 12 1 12 2 12 12 9 14 9 13 2
26 3 7 10 12 9 3 9 13 2 9 9 9 1 9 14 16 1 9 9 10 9 13 2 9 13 2
15 10 9 1 9 0 1 9 9 0 1 9 0 9 13 2
25 10 9 0 9 0 9 0 7 9 0 0 13 16 9 9 1 1 9 9 0 15 14 9 13 2
13 9 0 1 9 13 16 1 9 12 9 13 13 2
44 9 9 0 9 9 13 16 9 0 1 9 2 7 9 0 0 1 9 2 7 9 16 1 9 0 1 9 13 0 1 9 0 9 0 9 13 2 9 0 9 2 12 2 2
39 1 9 12 2 12 9 9 1 9 9 9 9 0 9 1 9 0 9 2 9 7 9 15 1 9 9 9 7 9 9 9 9 13 2 9 2 12 2 2
13 9 0 14 9 1 9 12 7 12 9 13 13 2
12 3 0 1 12 9 1 9 9 0 9 13 2
18 9 0 9 0 2 9 9 1 9 13 16 0 1 9 1 9 13 2
26 9 0 0 1 10 9 9 9 9 1 9 3 7 0 9 9 9 1 9 7 9 9 1 15 13 2
42 1 9 12 9 0 9 13 16 9 9 9 3 9 14 0 13 7 1 9 9 0 13 2 7 0 1 9 1 15 9 13 16 1 9 9 9 0 1 15 9 13 2
15 9 0 9 13 16 9 9 0 14 0 9 0 9 13 2
37 10 9 3 1 9 12 1 9 9 1 9 9 9 9 13 7 3 1 9 9 1 9 9 12 2 9 2 12 2 7 1 9 9 12 9 13 2
25 7 1 9 9 9 9 16 9 9 13 2 0 13 16 9 0 14 0 9 9 13 16 0 13 2
16 9 9 1 9 0 9 13 16 1 9 9 9 0 13 13 2
38 9 2 12 2 9 13 16 1 9 9 1 9 0 1 9 0 1 9 0 2 9 9 13 3 9 4 9 9 7 9 14 1 9 3 9 9 13 2
10 10 9 3 1 12 9 0 9 13 2
17 1 9 9 12 2 0 9 0 13 16 1 9 9 9 9 13 2
20 15 0 15 13 16 9 1 9 2 3 1 1 9 1 9 9 9 0 13 2
27 0 9 9 13 16 9 9 7 9 15 14 9 13 2 3 16 0 1 9 7 1 9 0 0 13 13 2
40 16 1 9 1 9 0 1 9 1 9 0 2 9 9 0 7 0 2 16 9 9 0 2 1 9 7 9 15 9 13 16 9 14 9 0 9 15 9 13 2
17 9 0 16 1 9 1 9 0 2 9 0 14 1 9 9 13 2
42 9 9 9 9 1 9 7 9 9 0 10 9 16 1 9 16 1 9 2 9 2 9 13 7 7 2 1 1 0 2 1 9 0 16 1 9 0 9 13 0 13 2
70 12 2 9 12 2 12 2 9 2 1 9 9 2 0 12 2 0 13 16 9 0 1 9 9 0 13 7 16 3 9 4 0 9 0 13 2 9 2 10 9 9 0 1 9 7 9 9 16 10 9 14 9 13 2 9 2 10 9 9 1 9 0 9 16 1 9 0 0 13 2
26 12 2 9 7 9 0 1 9 0 1 9 9 0 13 7 0 13 0 9 7 9 7 9 0 13 2
22 12 2 9 9 0 16 1 9 9 13 13 4 1 9 9 7 9 1 9 0 13 2
31 12 2 10 9 9 4 9 13 16 9 7 9 9 0 1 9 0 1 9 13 7 9 0 1 10 9 0 7 0 13 2
31 12 2 1 9 0 9 0 9 12 7 12 4 9 2 9 7 9 9 0 0 14 16 3 1 9 9 13 2 0 13 2
16 10 9 3 0 13 2 7 9 0 16 1 10 9 9 13 2
18 9 0 16 1 9 0 9 13 4 9 0 14 1 10 9 9 13 2
42 12 2 1 9 4 9 14 13 16 1 9 16 9 3 7 3 0 13 2 9 7 9 9 0 9 13 2 3 15 7 10 9 1 9 9 12 1 10 9 0 13 2
9 10 9 0 9 0 1 9 13 2
35 12 2 1 9 0 4 1 9 9 7 9 7 9 9 0 9 13 2 7 9 0 9 0 14 4 1 9 9 1 9 0 0 9 13 2
22 7 1 9 7 9 0 15 4 1 9 0 9 7 0 9 9 9 10 9 9 13 2
33 12 2 1 9 16 9 0 2 3 9 2 9 2 9 7 9 0 9 2 16 9 0 1 12 9 13 2 1 9 9 0 13 2
15 9 9 12 2 12 1 9 9 9 9 1 15 0 13 2
47 10 9 9 13 16 9 0 1 9 2 9 2 9 7 9 2 7 9 0 16 1 9 9 9 13 2 1 1 9 0 9 7 9 13 2 9 9 9 9 10 9 9 0 14 0 13 2
19 9 9 0 1 9 0 1 9 2 4 1 9 0 1 9 0 9 13 2
24 1 9 7 1 9 0 0 9 9 13 2 7 10 9 9 13 13 2 9 9 0 0 13 2
11 9 9 0 4 1 9 15 9 9 13 2
30 1 1 9 9 0 1 9 7 9 2 4 1 15 9 13 16 3 1 10 9 9 1 9 2 1 9 15 9 13 2
35 12 2 9 0 2 0 16 9 12 2 12 15 14 0 13 2 13 9 0 1 9 9 13 2 7 9 0 1 9 0 14 13 9 13 2
29 12 2 9 0 1 9 9 0 1 9 0 4 3 9 13 16 3 9 9 1 9 2 1 9 15 2 4 13 2
20 9 9 4 15 14 1 9 0 13 16 9 0 1 9 9 7 9 0 13 2
57 12 2 10 9 0 7 9 1 15 3 1 9 7 9 9 1 9 0 7 9 1 9 9 13 2 1 10 9 2 9 0 4 1 1 9 9 7 9 1 15 1 9 9 9 15 7 9 9 0 1 9 0 1 9 15 13 2
29 12 2 1 1 9 0 7 0 2 9 0 4 0 9 0 9 7 9 0 7 9 0 1 1 9 0 15 13 2
34 12 2 9 9 2 9 2 1 9 1 15 7 3 9 9 1 9 0 9 9 9 13 2 4 9 0 1 9 1 9 0 0 13 2
24 12 2 9 9 0 14 1 9 7 9 0 1 9 13 7 10 9 0 9 0 0 15 13 2
23 9 1 10 9 1 15 9 0 13 16 3 1 9 1 9 0 2 1 10 9 0 13 2
28 1 9 7 9 9 9 0 0 13 16 1 9 9 0 2 16 9 9 0 0 1 9 9 13 2 9 13 2
13 1 9 1 9 15 2 0 1 1 15 9 13 2
26 10 9 12 9 13 7 15 1 9 15 0 13 7 3 9 0 12 9 0 13 16 13 1 9 9 2
11 9 1 9 9 9 0 1 9 0 13 2
11 3 3 0 0 13 7 12 9 0 13 2
26 1 1 9 9 15 7 9 0 7 3 9 10 9 9 0 13 7 1 9 12 9 1 15 9 13 2
29 1 9 0 9 3 0 13 2 3 12 9 3 9 9 1 9 9 0 15 3 0 13 7 15 12 0 0 13 2
11 15 1 10 9 9 14 13 3 9 0 2
14 1 9 0 16 9 15 13 2 3 0 10 9 13 2
13 15 14 13 7 4 9 13 2 1 1 3 13 2
5 3 9 0 13 2
20 9 14 16 9 13 2 3 15 15 2 15 13 13 7 1 1 9 9 13 2
25 9 9 15 7 9 3 9 13 16 1 10 9 3 0 13 1 9 16 9 1 9 15 9 13 2
45 3 9 9 13 16 9 0 13 7 15 1 9 9 16 13 9 13 7 9 9 13 13 7 12 9 13 7 1 9 16 9 13 13 7 13 7 13 7 1 12 9 0 9 13 2
13 15 1 9 10 9 7 9 10 9 3 0 13 2
5 15 9 9 13 2
29 9 3 0 9 0 15 15 13 7 3 9 15 9 14 1 15 0 13 16 0 13 13 9 15 15 14 0 13 2
11 9 9 1 10 9 9 12 9 0 13 2
8 13 2 16 9 13 0 13 2
7 9 9 7 10 9 13 2
24 1 9 15 2 9 16 3 13 3 0 9 13 1 9 16 4 9 1 9 9 1 9 13 2
40 15 9 14 9 13 7 15 15 16 1 9 0 13 16 9 1 9 9 13 2 7 3 9 0 4 9 0 13 2 3 13 1 10 9 13 13 7 7 3 2
40 9 16 1 9 0 13 7 9 13 9 3 9 0 13 10 9 9 15 13 2 16 15 0 9 15 13 16 1 9 9 16 9 13 7 16 13 7 16 13 2
33 10 9 15 9 13 15 9 14 1 9 13 7 12 9 0 0 13 13 7 3 1 9 15 13 16 9 3 9 9 14 9 13 2
16 3 15 4 3 10 9 14 9 13 1 1 10 3 9 13 2
15 1 9 15 2 1 10 10 9 0 7 0 7 0 13 2
20 3 1 9 0 15 12 9 0 13 1 9 16 12 9 1 9 9 13 13 2
17 15 3 0 13 7 1 12 9 1 10 9 12 9 15 9 13 2
15 10 12 9 2 12 9 12 9 14 1 15 15 9 13 2
34 1 10 9 3 10 9 13 2 7 3 9 3 9 15 14 0 13 7 9 13 16 9 0 13 7 9 9 13 16 9 1 9 13 2
8 9 13 7 15 16 9 13 2
29 10 9 16 1 1 9 1 9 0 13 2 15 15 0 13 7 10 9 9 2 16 9 0 13 2 3 9 13 2
8 9 15 1 9 9 0 13 2
17 1 9 0 9 0 9 13 2 7 3 15 9 0 9 9 13 2
42 15 15 14 1 2 9 9 2 9 13 7 9 13 2 7 1 9 9 1 10 7 3 9 13 10 9 14 13 2 13 2 16 1 10 9 2 9 9 2 9 13 2
30 16 9 0 13 13 7 2 9 9 2 12 3 1 15 9 13 7 9 0 1 15 9 13 2 13 3 9 13 13 2
44 7 9 9 12 9 9 13 2 12 15 7 9 16 4 9 13 7 3 9 0 9 13 7 1 12 9 9 13 2 12 9 0 14 13 7 12 9 1 9 0 15 3 13 2
23 3 9 9 3 9 9 13 7 9 3 0 16 13 7 3 10 9 9 13 1 15 13 2
26 15 1 9 15 7 1 9 0 15 3 15 13 7 16 9 15 14 16 13 2 12 0 1 9 13 2
23 7 9 9 2 13 12 0 9 13 1 9 0 15 7 9 13 13 2 1 15 9 13 2
4 9 13 13 2
5 6 2 9 13 2
17 9 16 13 9 13 16 3 9 13 9 3 13 2 3 9 9 2
16 15 3 15 9 13 0 13 2 16 9 9 3 0 0 13 2
31 3 16 9 13 3 9 13 7 3 1 12 9 2 3 0 13 2 3 12 2 12 9 0 2 15 9 9 9 14 13 2
26 3 12 9 13 16 15 15 15 12 9 0 1 15 13 2 15 9 7 9 13 7 9 7 7 9 2
11 3 10 9 9 9 13 16 3 9 13 2
19 1 1 15 12 9 0 13 2 16 15 9 15 9 0 9 9 14 13 2
25 9 0 15 13 16 9 3 0 1 9 16 1 9 0 13 0 13 2 16 1 9 9 0 13 2
48 9 0 13 16 10 9 15 14 9 13 2 3 1 2 9 9 2 13 16 9 9 2 1 15 7 9 13 2 12 9 0 7 0 13 2 7 7 9 9 16 0 13 2 9 14 9 13 2
18 13 13 16 0 13 10 9 13 7 10 9 0 14 1 9 9 13 2
8 16 9 13 10 9 14 13 2
4 3 0 13 2
18 10 9 16 9 13 2 9 7 9 7 9 2 9 15 16 9 13 2
17 10 9 1 2 9 9 2 13 7 9 13 1 10 9 3 13 2
29 3 9 9 16 0 13 2 3 9 0 13 7 3 12 9 0 7 0 16 13 2 0 15 9 16 1 9 13 2
28 15 15 15 0 13 7 0 15 16 15 9 13 2 15 9 0 13 7 9 0 1 15 0 2 0 2 13 2
7 9 13 16 3 0 13 2
29 7 10 9 0 15 2 16 3 1 15 13 9 7 13 1 9 0 2 9 9 0 9 14 1 1 10 9 13 2
67 15 15 15 1 9 13 7 13 16 0 9 3 9 0 13 7 0 13 7 3 9 9 13 2 7 7 9 1 9 13 3 0 13 2 0 13 2 7 9 1 10 9 0 13 2 3 9 0 13 2 3 3 0 7 0 13 7 0 2 0 9 16 15 1 9 13 2
45 3 16 13 1 9 2 9 9 0 14 1 9 0 9 13 2 9 9 0 3 1 15 0 7 0 13 13 2 9 3 0 13 2 16 1 9 7 16 1 9 7 3 1 9 2
20 1 9 0 9 13 2 3 3 1 9 9 9 13 16 9 1 15 9 13 2
12 3 15 0 13 7 7 1 0 10 9 13 2
15 1 10 9 15 9 10 9 14 1 9 10 9 9 13 2
24 16 1 9 12 7 0 10 9 14 1 9 9 12 7 0 10 9 9 13 2 9 0 13 2
89 9 13 12 2 12 9 10 9 16 13 2 12 9 1 15 9 13 16 10 9 1 9 2 9 9 2 2 16 15 15 13 13 2 9 13 7 13 16 10 9 3 1 15 0 7 0 13 7 16 3 9 2 9 9 2 13 7 9 15 2 10 9 1 9 3 13 16 15 12 9 1 9 15 13 16 12 1 9 14 9 13 7 3 12 9 0 14 13 2
16 15 3 9 0 13 7 3 10 9 14 13 7 13 9 13 2
7 9 13 12 9 0 13 2
34 12 9 0 16 10 9 14 0 13 15 13 16 3 9 13 16 10 9 3 16 9 0 7 0 16 9 13 12 9 0 13 2 13 2
6 15 1 9 0 13 2
6 15 9 15 14 13 2
5 12 9 0 13 2
18 12 9 2 3 1 9 9 2 15 15 1 10 9 15 15 0 13 2
33 3 12 9 9 9 13 2 2 9 2 15 16 10 9 1 9 7 9 15 13 7 3 4 9 13 2 3 13 9 0 13 2 2
13 15 12 9 13 1 9 13 16 10 9 0 13 2
9 16 3 9 9 15 15 9 13 2
33 1 9 3 0 16 1 9 13 2 7 15 9 13 3 0 13 2 15 13 16 9 2 3 15 15 14 1 2 6 2 9 13 2
71 15 9 13 16 16 10 0 13 7 0 13 7 3 15 15 14 1 9 9 7 9 9 13 2 16 15 13 12 9 0 13 13 2 4 15 10 9 14 13 13 2 7 3 9 0 9 15 1 3 1 10 9 0 13 2 7 16 9 7 9 1 15 9 13 2 15 10 9 14 13 2
17 9 1 10 9 9 13 16 15 9 16 1 9 9 13 0 13 2
16 9 15 9 13 16 9 4 3 9 13 2 7 3 13 13 2
21 10 9 13 13 16 9 15 9 9 13 7 12 9 4 13 16 15 9 9 13 2
10 16 9 0 13 13 13 2 15 13 2
5 1 9 9 13 2
23 1 9 0 9 13 1 9 9 16 1 9 12 10 9 0 2 1 9 9 3 9 13 2
6 1 10 9 15 13 2
12 15 1 10 9 3 9 14 0 10 9 13 2
4 16 3 13 2
69 3 1 15 7 9 14 1 15 9 13 16 9 13 2 15 3 9 13 2 1 9 15 7 9 3 9 13 13 16 3 13 2 7 15 13 13 13 2 7 15 3 9 13 2 16 12 9 9 16 9 0 13 2 0 13 7 1 15 0 13 7 3 0 13 9 14 9 13 2
15 12 9 15 13 16 10 9 14 13 7 1 15 9 13 2
6 15 3 9 0 13 2
30 16 15 9 13 1 9 2 1 10 9 1 15 12 9 0 1 9 13 16 1 12 9 7 7 12 9 1 9 13 2
27 3 12 9 13 16 15 1 12 9 9 13 7 3 13 9 2 9 0 13 2 12 9 0 1 15 13 2
4 3 9 13 2
6 9 15 9 3 13 2
29 3 15 4 15 14 13 2 12 9 9 9 1 9 13 2 16 15 10 9 14 13 2 16 9 15 0 13 13 2
61 9 13 16 7 15 3 3 1 15 7 9 7 9 3 9 15 9 13 7 1 9 13 2 13 9 14 9 13 2 4 12 9 0 1 9 13 7 12 16 1 9 2 16 15 12 9 13 2 1 9 15 2 16 9 13 16 4 9 15 13 2
6 10 9 14 13 13 2
16 9 0 15 13 16 9 14 13 0 10 9 2 16 0 13 2
44 10 9 0 1 0 9 15 0 12 9 3 9 13 13 2 16 15 16 9 14 13 16 9 9 13 2 13 16 9 2 15 0 15 13 3 2 9 1 10 9 9 13 13 2
33 10 9 0 15 13 16 15 12 9 0 13 16 9 9 9 13 7 1 12 9 0 2 16 12 10 9 0 7 12 10 9 0 2
4 15 9 13 2
34 9 13 16 10 9 3 13 2 3 10 9 12 9 0 13 2 12 9 3 0 2 16 9 0 13 7 15 9 13 13 1 9 0 2
27 3 9 9 16 13 9 13 16 12 9 1 10 12 9 13 2 16 3 0 7 0 13 7 3 0 13 2
11 1 9 9 13 7 13 4 3 9 13 2
11 0 9 9 1 0 9 9 3 0 13 2
7 1 9 15 1 9 13 2
11 7 9 16 13 1 9 13 7 0 13 2
33 7 3 9 16 9 0 3 9 9 13 7 3 12 9 13 2 9 16 3 1 9 15 9 16 0 13 2 12 9 0 1 9 2
23 1 9 0 12 9 3 0 13 2 9 9 7 9 2 16 15 9 9 7 9 9 13 2
13 7 1 9 0 9 13 9 13 10 9 9 13 2
7 10 9 9 14 0 13 2
8 16 9 0 9 13 2 3 2
15 1 9 2 9 15 1 10 9 3 0 1 9 0 13 2
24 9 9 0 9 0 15 3 12 9 9 0 10 9 13 7 1 1 9 0 16 9 0 13 2
23 3 10 9 13 7 3 10 9 9 3 0 13 16 12 9 9 0 13 7 9 1 9 2
18 3 16 13 9 13 16 15 1 12 9 9 13 13 2 3 0 13 2
13 7 3 10 9 14 13 2 0 1 9 9 0 2
8 3 13 9 0 13 2 3 2
24 16 1 9 0 12 9 9 13 7 3 15 7 12 9 1 15 13 7 7 1 15 0 13 2
24 16 1 15 13 2 3 15 9 3 1 9 13 2 7 16 1 15 13 2 9 9 0 13 2
56 3 9 0 14 13 1 7 3 1 12 9 0 9 13 2 16 12 9 9 15 14 9 13 7 12 9 10 9 13 7 3 9 0 9 15 1 0 10 9 13 7 12 9 0 13 7 9 1 9 9 10 9 1 9 13 2
12 3 3 9 14 9 0 13 2 10 9 13 2
13 3 0 13 1 12 9 12 1 15 3 0 13 2
7 3 1 9 0 10 9 2
17 12 9 3 9 9 1 9 13 7 9 9 0 13 2 7 3 2
16 1 9 0 16 13 15 13 16 3 9 14 0 7 9 13 2
19 1 10 9 12 9 0 13 2 7 3 0 0 13 2 3 12 9 13 2
25 10 9 2 9 9 0 2 1 3 9 0 13 7 0 13 7 13 9 13 15 0 13 7 0 2
33 1 9 0 15 9 14 13 16 0 7 0 13 7 9 14 13 16 0 7 0 13 2 7 3 3 2 15 12 9 0 15 13 2
8 9 13 16 13 3 9 13 2
6 1 1 9 9 13 2
29 9 14 15 1 9 9 13 16 9 9 0 9 13 3 2 1 9 0 15 15 2 12 9 0 7 9 9 0 2
25 3 13 16 3 1 10 9 15 15 13 3 7 12 9 0 13 7 3 9 4 1 15 9 13 2
6 3 1 9 9 13 2
16 12 9 9 13 2 12 1 9 9 15 9 13 1 9 9 2
56 9 0 9 13 16 1 9 0 9 13 7 0 1 9 3 10 7 9 1 12 9 3 13 16 0 13 3 4 9 15 13 2 12 9 12 2 0 14 1 9 15 13 2 7 3 9 3 1 9 13 16 9 9 14 13 2
18 0 9 14 9 13 2 16 9 0 16 13 2 7 0 9 9 13 2
9 9 0 13 7 9 0 16 13 2
41 15 1 9 0 15 9 14 9 13 16 0 13 1 9 0 12 9 9 16 9 13 2 7 3 13 9 13 16 3 9 13 16 9 15 3 0 13 7 9 13 2
8 9 9 3 1 9 0 13 2
7 3 2 15 12 9 13 2
47 9 0 15 13 16 15 12 9 1 9 13 1 9 2 9 12 2 16 9 9 13 7 9 12 9 14 9 13 16 9 9 13 7 3 3 9 13 7 15 10 9 15 14 1 9 13 2
11 3 9 1 9 13 7 12 9 0 13 2
12 15 1 15 9 13 16 13 1 10 9 13 2
21 0 15 7 10 9 16 9 9 0 3 9 13 13 2 7 1 10 9 0 13 2
18 15 3 9 13 16 9 15 14 3 9 13 2 16 9 15 0 13 2
17 7 16 9 13 2 0 9 13 2 16 9 1 15 9 0 13 2
38 13 1 12 10 9 9 13 16 0 9 13 2 16 15 15 3 9 1 9 0 9 13 7 9 3 4 10 9 0 15 14 1 1 9 0 15 13 2
37 13 16 9 3 1 9 9 9 1 9 2 0 1 9 9 13 13 2 15 9 13 1 9 10 9 0 9 1 9 13 2 15 10 9 9 13 2
18 3 2 1 9 15 13 16 9 1 3 12 9 1 9 15 9 13 2
37 13 9 10 9 3 9 13 2 12 9 13 16 1 9 4 9 13 7 9 13 7 1 9 9 9 13 7 9 0 13 7 1 9 9 9 13 2
22 16 15 13 12 9 16 9 1 9 15 13 13 2 16 1 3 15 14 13 2 13 2
11 3 15 1 9 9 15 15 14 0 13 2
18 9 13 16 9 13 0 13 2 7 3 0 1 9 13 7 9 0 2
6 1 9 15 16 13 2
17 1 9 9 10 9 3 0 13 16 9 10 9 0 15 9 13 2
32 15 3 13 3 1 9 0 15 15 9 13 2 16 9 0 13 13 2 7 15 9 13 2 16 9 4 1 10 9 9 13 2
12 13 3 9 13 16 9 15 15 4 9 13 2
18 9 0 12 9 1 9 9 9 13 7 3 16 13 9 15 14 13 2
17 3 16 13 9 14 9 13 2 9 0 13 2 9 15 15 15 2
17 9 1 15 9 13 2 7 15 0 13 16 3 1 0 9 13 2
3 9 13 2
23 3 2 16 9 15 13 2 1 9 0 9 1 9 9 9 1 12 2 12 9 9 13 2
17 9 12 9 3 0 7 0 7 0 2 3 9 13 1 0 9 2
18 3 15 0 13 2 13 9 13 1 9 16 9 1 15 0 15 13 2
9 3 13 16 3 2 3 0 13 2
12 15 9 13 16 0 13 9 13 7 7 13 2
52 9 16 1 9 15 0 13 15 13 16 1 9 0 13 12 9 0 16 1 9 13 2 9 13 7 1 9 12 9 1 9 15 13 7 1 15 9 13 2 1 9 9 7 2 1 10 9 1 15 9 13 2
12 12 3 9 3 9 13 2 3 9 9 9 2
31 9 9 1 9 15 16 9 15 13 7 10 9 16 1 15 13 7 9 16 9 1 15 13 2 3 1 10 9 0 13 2
9 9 9 13 9 15 4 0 13 2
7 10 9 1 3 9 13 2
17 15 12 1 0 9 15 9 9 13 2 16 1 9 13 13 15 2
15 9 9 1 9 9 3 0 13 7 9 16 1 15 13 2
28 1 9 3 3 0 13 7 1 9 9 16 13 2 9 13 1 9 0 9 13 16 12 1 15 9 9 13 2
24 1 9 9 1 15 0 13 7 1 9 0 16 9 9 1 15 9 13 7 3 1 15 13 2
26 3 1 10 9 9 9 15 14 13 9 2 16 9 15 15 14 13 2 16 3 1 9 15 9 13 2
25 1 9 15 7 9 15 3 10 9 13 2 9 16 15 9 9 14 13 2 9 15 3 0 13 2
32 7 10 9 16 15 1 9 13 2 4 9 15 3 0 7 0 13 7 3 9 15 15 0 7 0 7 12 9 0 1 9 2
15 13 16 10 9 0 9 13 7 3 15 14 3 9 13 2
7 9 9 15 3 9 13 2
29 3 1 15 7 12 9 1 12 9 1 15 9 13 2 9 14 0 13 7 12 9 0 14 3 1 9 0 13 2
11 1 9 9 9 9 12 9 9 3 13 2
13 7 9 13 3 10 9 2 3 9 0 16 13 2
10 3 9 15 14 13 1 1 9 15 2
10 10 0 9 14 3 1 9 15 13 2
10 16 3 1 9 13 9 15 14 13 2
16 16 3 9 9 0 0 9 13 7 9 1 15 9 13 13 2
2 13 2
31 3 15 10 9 14 13 7 9 13 1 10 9 9 16 0 1 13 2 9 9 13 7 3 16 9 2 9 3 1 13 2
29 3 9 16 15 4 13 1 9 12 9 13 16 9 13 7 9 16 15 13 1 9 12 2 12 9 13 16 13 2
21 7 0 13 16 9 0 2 10 9 9 9 13 2 7 0 3 13 13 3 13 2
14 15 7 4 13 16 0 13 13 7 0 13 7 13 2
10 7 3 9 9 9 10 9 9 13 2
15 9 16 9 13 0 13 2 7 9 12 9 0 9 13 2
8 10 9 1 1 9 0 13 2
17 1 9 15 9 0 13 16 9 0 1 9 0 1 15 0 13 2
15 10 9 9 1 15 1 9 0 13 7 15 15 9 13 2
6 7 1 3 9 13 2
20 3 2 10 9 9 14 9 0 1 15 15 0 13 2 16 9 9 13 3 2
15 15 13 12 9 13 7 13 7 10 9 13 7 9 13 2
16 3 9 0 1 9 9 13 16 13 9 1 10 9 4 13 2
14 15 1 10 9 3 3 1 9 13 2 1 9 13 2
9 1 10 9 12 9 1 9 13 2
9 1 9 16 1 3 13 13 13 2
31 15 1 9 9 13 7 3 9 1 15 13 3 10 9 14 13 2 0 13 1 9 16 13 9 14 9 13 2 9 13 2
11 15 0 13 12 9 1 9 9 9 13 2
11 1 9 15 7 10 9 9 9 9 13 2
38 3 15 16 1 9 3 9 13 2 3 4 9 13 16 9 0 13 7 3 15 13 1 12 9 13 7 1 12 9 12 9 0 13 7 9 0 13 2
43 9 16 16 0 13 2 13 9 13 1 12 9 7 1 12 9 9 7 9 0 7 13 12 9 0 1 9 13 7 15 1 9 9 9 13 16 15 15 1 3 0 13 2
25 9 9 0 13 7 15 16 1 9 9 9 0 13 2 7 3 1 10 9 16 1 9 9 13 2
22 3 1 9 0 9 9 16 10 9 10 9 14 3 1 9 13 2 13 2 9 13 2
10 7 9 13 2 1 3 9 7 9 2
9 3 3 12 2 12 9 9 13 2
29 9 0 16 1 9 2 1 9 0 2 1 9 9 7 1 9 13 2 1 9 13 7 3 3 3 1 9 13 2
16 3 12 1 0 9 16 15 1 3 13 2 10 9 0 13 2
7 1 9 0 3 0 13 2
11 3 9 1 9 1 9 9 14 9 13 2
6 0 13 2 9 13 2
19 9 0 3 0 13 2 3 0 7 9 15 3 0 13 7 1 9 13 2
18 3 0 7 0 13 7 9 9 3 0 13 7 9 9 16 10 9 2
12 15 15 3 0 13 2 1 0 9 14 13 2
5 9 0 0 13 2
5 3 3 9 13 2
7 3 15 7 9 13 13 2
12 12 9 13 9 7 9 13 7 12 14 13 2
6 9 9 3 0 13 2
22 1 10 9 7 9 13 7 9 13 7 0 13 7 1 9 13 2 9 0 0 13 2
11 9 9 13 16 10 9 0 7 0 13 2
24 10 9 7 12 9 0 0 9 13 16 9 7 9 16 13 9 0 13 7 9 9 9 13 2
22 15 14 16 13 16 1 12 9 9 2 1 0 9 2 10 10 9 9 1 9 13 2
19 13 16 4 1 1 9 9 13 2 13 10 9 0 9 0 14 13 13 2
14 9 9 13 10 9 0 14 2 9 15 9 0 13 2
7 10 9 9 0 9 13 2
49 10 9 16 1 12 9 0 13 2 0 13 4 3 9 1 15 13 2 3 9 16 3 2 1 10 9 16 15 9 13 2 9 10 9 12 9 13 2 9 16 9 7 9 13 1 9 15 13 2
40 9 16 1 9 1 15 9 13 13 2 12 9 0 7 10 9 9 9 14 13 2 9 9 13 2 1 9 7 3 10 9 13 7 9 0 3 3 0 7 2
32 9 16 9 13 7 10 10 9 13 1 9 16 12 9 13 13 16 13 2 9 2 9 9 14 13 2 9 9 14 0 13 2
6 3 3 3 0 13 2
23 3 15 9 13 16 9 9 3 9 13 7 9 14 0 13 7 1 9 7 9 9 13 2
5 10 9 0 13 2
9 9 9 9 9 0 7 0 13 2
15 3 9 2 9 15 16 10 9 4 9 14 13 2 13 2
25 3 9 16 1 9 9 13 2 9 13 1 9 0 2 9 0 7 0 7 0 7 12 9 9 2
26 15 7 10 9 9 13 7 3 9 13 7 9 9 13 7 12 9 16 13 2 3 13 9 16 3 2
31 7 9 9 1 9 16 9 0 13 2 1 9 16 1 9 9 7 12 0 1 9 9 1 9 9 13 2 13 3 13 2
11 9 1 9 15 13 2 13 9 3 13 2
16 10 12 9 9 13 7 10 9 16 1 9 9 13 9 13 2
14 16 3 9 13 9 3 13 7 3 9 13 16 13 2
9 9 9 14 15 15 9 13 13 2
3 0 13 2
6 15 15 9 13 13 2
4 9 0 13 2
9 16 0 9 1 9 10 9 13 2
19 3 9 1 9 2 9 12 9 2 13 3 7 0 9 9 0 9 13 2
18 15 4 13 16 9 13 9 0 12 10 9 0 2 9 0 7 0 2
30 9 13 16 15 9 1 9 3 0 13 7 15 9 1 9 1 0 9 15 16 13 7 0 1 12 9 9 0 13 2
12 1 9 15 7 1 9 15 10 9 13 13 2
12 3 3 16 0 13 7 15 13 1 15 13 2
21 1 9 2 1 9 0 2 9 12 9 2 2 3 15 9 9 0 7 0 13 2
14 3 9 1 15 13 7 3 13 10 9 14 9 13 2
20 3 15 9 13 16 1 0 9 0 2 9 15 9 2 9 13 1 0 9 2
14 9 13 10 0 9 1 9 9 9 7 9 9 13 2
11 3 15 9 9 15 16 15 15 0 13 2
37 9 16 3 9 13 2 9 1 15 13 16 3 9 0 1 9 9 9 13 16 16 9 9 15 0 13 2 15 9 15 14 0 13 2 0 13 2
22 16 9 9 15 0 13 2 15 1 1 9 3 9 14 13 16 13 2 9 9 13 2
39 7 15 1 9 13 16 15 15 7 15 9 1 15 15 9 13 2 16 16 1 9 9 10 12 9 1 15 13 2 0 9 9 13 7 3 9 9 13 2
13 7 10 9 13 2 1 9 0 15 7 9 13 2
13 3 9 0 13 7 3 13 13 16 1 15 13 2
16 10 1 15 9 1 9 0 7 0 13 16 9 13 1 9 2
35 1 15 7 15 3 9 14 0 13 7 3 13 1 10 9 0 7 0 7 13 9 10 9 9 13 7 1 10 9 10 12 9 9 2 2
26 1 9 15 2 9 16 1 9 9 7 9 9 13 2 3 9 0 13 16 10 12 9 1 15 13 2
45 9 10 12 9 16 1 0 12 9 9 0 2 12 9 9 0 13 7 3 16 3 10 12 9 1 15 9 13 7 15 9 1 9 7 9 0 13 2 0 9 14 15 13 13 2
29 3 9 0 3 13 16 16 15 1 15 13 2 9 0 13 7 0 13 7 3 1 9 15 1 15 9 9 13 2
8 3 9 0 3 15 9 13 2
22 1 9 15 7 1 0 9 9 2 7 0 9 15 4 12 10 9 14 1 15 13 2
23 16 1 9 4 12 10 9 14 13 7 15 14 1 9 0 9 13 1 1 9 0 13 2
12 9 0 16 15 9 9 13 7 9 13 13 2
26 15 7 10 12 9 1 15 13 2 3 0 13 7 15 14 15 13 16 9 0 2 10 9 3 13 2
34 3 12 9 13 16 1 15 9 7 9 13 7 9 13 2 3 9 13 16 1 15 9 15 14 13 7 3 16 3 1 15 9 13 2
21 9 3 0 13 16 16 13 13 15 13 16 1 3 2 15 9 0 14 9 13 2
2 6 2
23 16 9 1 10 9 0 9 13 7 9 10 9 9 13 16 9 13 9 0 14 0 13 2
11 13 15 1 9 0 9 13 16 0 13 2
14 9 16 9 7 9 1 15 9 13 16 9 0 13 2
25 13 9 9 7 1 15 13 16 9 15 0 13 2 3 1 0 9 7 9 7 9 7 9 2 2
12 15 9 13 7 9 1 9 7 9 0 13 2
28 16 1 10 9 2 9 7 9 1 15 9 13 3 0 13 2 16 15 13 7 13 2 9 10 3 9 13 2
10 1 10 9 0 13 16 9 0 13 2
12 3 1 10 9 13 16 15 9 4 0 13 2
54 9 1 9 1 9 9 13 2 0 9 15 13 16 0 9 9 0 13 2 9 9 13 7 7 16 1 9 3 9 13 2 0 9 15 13 16 10 9 14 1 12 9 1 9 9 2 9 15 13 2 15 16 3 2
14 16 1 9 0 13 12 9 9 13 7 3 9 13 2
6 16 3 9 0 13 2
8 3 9 13 10 9 0 13 2
13 3 0 10 9 3 0 13 7 3 9 0 13 2
58 15 9 13 9 7 9 16 1 9 9 13 2 1 9 3 1 12 9 9 0 15 7 15 1 15 9 13 7 9 0 13 1 9 9 13 7 3 9 15 14 9 13 7 3 10 9 16 3 9 13 16 12 9 0 3 9 13 2
11 3 15 0 13 2 16 9 13 7 9 2
11 15 7 12 10 9 0 0 14 9 13 2
22 3 15 7 13 2 15 1 9 0 13 1 9 15 7 4 1 9 0 16 13 3 2
7 15 1 9 15 9 13 2
20 9 16 13 1 15 9 13 2 4 0 13 2 3 1 15 7 3 0 13 2
6 1 10 9 9 13 2
18 1 9 0 9 9 7 9 13 16 1 9 3 0 1 15 0 13 2
11 16 13 2 16 15 0 13 4 0 13 2
44 3 3 1 15 0 13 7 9 1 9 3 1 15 0 13 16 3 10 12 9 4 1 15 0 13 7 0 13 1 9 9 7 3 0 13 16 10 12 9 0 1 9 13 2
40 3 9 9 1 9 2 7 3 9 13 16 4 1 1 15 9 13 7 9 9 15 0 13 7 10 9 1 15 13 13 1 12 9 0 9 13 7 0 13 2
10 3 15 16 9 12 9 9 13 7 2
7 1 3 1 9 9 9 2
12 3 1 9 9 0 13 7 9 0 7 0 2
10 1 9 0 9 9 0 13 7 9 2
42 9 16 9 9 13 7 9 0 15 2 0 10 9 13 16 12 9 10 9 14 13 2 16 10 9 16 4 10 9 14 13 2 3 9 0 13 2 3 9 15 13 2
14 4 9 13 13 1 9 9 16 9 9 15 9 13 2
15 9 16 3 16 13 12 9 0 9 13 2 0 15 13 2
12 16 9 13 9 3 0 13 7 9 3 0 2
3 0 13 2
17 1 1 9 15 2 15 9 0 14 9 13 7 9 0 14 9 2
17 15 7 9 1 15 12 9 0 9 9 3 0 13 7 3 9 2
19 3 9 4 9 13 16 9 14 13 0 7 0 9 9 14 1 9 0 2
5 15 3 9 13 2
20 15 13 16 9 1 15 13 16 15 12 9 9 0 14 1 12 9 0 13 2
22 9 13 10 9 12 12 9 13 7 12 12 1 12 9 1 15 9 9 3 9 13 2
14 7 10 9 1 12 9 13 13 7 15 16 0 9 2
11 1 9 15 1 3 9 1 9 0 13 2
14 15 9 13 3 9 1 9 9 9 9 14 13 13 2
56 10 2 9 12 9 2 9 16 1 15 13 2 1 9 12 9 15 12 2 12 9 9 13 7 12 9 0 12 9 4 10 9 9 9 12 1 9 15 13 3 7 9 12 2 12 13 1 9 15 1 3 12 9 13 13 2
20 1 9 7 15 9 13 7 16 10 12 9 2 12 9 13 3 9 0 13 2
12 1 15 2 9 12 9 0 13 9 13 13 2
18 9 13 16 13 13 9 10 9 15 12 9 9 13 1 12 9 15 2
38 3 9 1 12 9 0 0 2 1 9 3 0 9 2 1 1 9 2 12 2 12 9 9 13 2 7 12 9 12 9 14 13 1 12 9 9 13 2
19 15 16 9 1 9 2 9 1 9 7 12 9 9 13 16 1 9 13 2
13 1 9 15 2 9 1 9 0 1 9 9 13 2
19 16 9 3 0 13 7 15 9 9 15 15 14 13 2 7 1 9 3 2
15 15 12 1 9 13 16 9 13 7 1 9 16 9 13 2
39 9 3 9 0 13 7 10 9 9 9 9 1 9 0 7 9 7 9 0 9 9 13 7 15 7 3 1 9 1 9 0 13 1 1 9 7 9 9 2
31 7 15 9 15 1 9 0 15 13 16 1 3 1 9 9 0 2 10 9 9 1 10 9 13 16 0 1 9 9 13 2
20 9 13 1 10 9 1 9 1 9 9 9 9 13 7 10 9 0 0 13 2
8 3 9 3 9 9 15 13 2
9 1 10 9 2 9 9 0 13 2
23 16 9 16 3 15 9 0 13 2 3 1 9 13 10 9 0 13 2 16 9 0 13 2
5 16 3 9 13 2
5 15 15 9 13 2
12 13 2 9 9 3 0 13 7 9 0 13 2
8 9 12 9 1 9 9 13 2
27 16 15 7 10 9 3 4 1 9 13 16 9 1 15 13 2 9 15 0 13 2 15 3 13 9 13 2
32 15 0 13 16 10 9 9 12 9 0 13 7 0 13 1 9 7 9 9 13 2 7 9 1 9 12 9 3 2 3 13 2
12 1 10 9 2 4 9 1 9 15 3 13 2
15 0 1 10 9 13 16 9 0 13 16 9 9 0 13 2
36 16 10 9 13 2 3 1 9 16 0 9 0 13 2 3 15 4 3 9 0 13 2 1 9 7 3 15 0 13 7 1 12 9 9 13 2
7 3 2 9 15 15 13 2
7 16 15 9 0 15 13 2
17 16 1 1 9 0 3 3 9 13 7 3 9 7 9 14 13 2
17 16 15 1 9 9 13 2 16 13 12 9 1 10 9 9 13 2
10 4 10 9 0 13 7 10 9 13 2
50 9 16 1 10 9 13 2 15 13 16 10 9 12 10 9 15 2 3 2 10 9 1 9 0 1 0 1 15 15 9 13 2 1 0 1 0 3 0 2 7 1 0 1 3 3 10 9 14 13 2
25 1 9 3 15 2 3 1 9 1 9 9 9 13 2 16 3 10 9 15 14 16 1 9 13 2
15 1 9 0 13 16 9 13 10 9 4 3 9 0 13 2
43 10 9 3 3 13 2 9 14 9 13 2 3 3 9 13 1 9 7 1 10 9 13 15 1 15 9 13 2 7 1 10 9 2 16 9 13 2 16 0 13 1 15 2
22 1 9 0 3 13 1 9 7 1 9 0 3 0 13 7 3 1 15 15 9 13 2
12 3 1 9 7 9 15 3 9 13 0 13 2
10 9 1 15 15 7 9 0 0 13 2
11 15 1 10 9 0 1 9 3 0 13 2
22 1 9 9 2 3 15 16 9 0 13 2 0 0 13 2 16 10 9 0 14 13 2
13 3 1 10 9 16 9 0 13 13 2 9 13 2
6 15 1 9 0 13 2
50 1 12 9 0 13 16 3 3 9 13 16 9 16 1 9 12 9 9 13 2 0 13 0 13 7 0 13 3 9 0 13 2 7 9 16 0 13 2 9 0 13 2 16 9 2 9 0 9 13 2
11 0 13 10 9 1 9 12 9 9 13 2
15 10 9 7 15 3 2 9 12 9 3 13 2 0 13 2
23 7 16 9 0 16 9 13 12 9 13 7 12 9 0 12 9 0 2 3 9 9 13 2
21 1 9 2 1 9 9 0 13 13 16 3 3 9 2 9 12 9 2 9 13 2
44 15 9 13 1 9 15 13 16 12 9 0 1 9 0 1 9 0 13 7 9 13 16 15 13 7 9 16 9 1 9 15 13 3 1 9 9 2 9 12 9 2 14 13 2
13 9 3 2 9 0 2 9 9 2 9 2 9 2
23 15 15 9 13 2 1 15 0 7 1 15 0 13 7 15 7 9 13 4 9 15 13 2
13 1 9 7 15 13 9 0 4 9 14 9 13 2
16 9 0 1 9 15 13 16 1 9 0 9 1 9 9 13 2
13 16 1 9 9 9 9 7 9 9 15 14 13 2
25 3 10 9 16 13 0 13 1 9 9 0 13 7 0 13 9 16 15 13 13 2 15 13 13 2
21 3 9 16 3 10 9 14 13 2 10 9 14 13 16 15 3 1 15 0 13 2
24 7 15 0 13 16 15 14 4 13 2 1 15 7 9 9 2 9 1 9 13 7 4 13 2
9 1 9 15 3 1 9 9 13 2
20 1 15 7 9 9 13 7 1 9 9 15 9 7 9 2 9 7 3 13 2
4 3 9 13 2
11 0 15 0 13 7 10 9 14 0 13 2
10 15 9 0 13 16 9 14 0 13 2
18 3 1 9 0 2 9 12 9 2 2 9 12 1 9 13 1 9 2
4 3 0 13 2
26 16 1 1 10 9 9 7 0 2 3 0 13 7 13 12 9 0 0 13 7 12 9 0 0 13 2
4 7 0 13 2
13 15 13 16 9 14 0 13 2 16 10 9 0 2
13 1 10 9 16 10 9 13 2 9 13 0 13 2
11 16 1 12 9 9 0 0 9 0 13 2
24 7 15 13 16 16 0 10 9 14 16 1 9 13 2 13 13 2 3 13 1 15 9 13 2
5 15 9 0 13 2
7 3 10 9 4 9 13 2
7 9 0 3 10 9 13 2
8 3 15 15 13 7 7 13 2
17 9 16 13 15 13 16 1 9 1 1 9 0 4 9 9 13 2
16 0 13 3 1 0 9 10 12 9 2 9 0 16 13 13 2
9 1 10 9 2 0 9 15 13 2
34 0 9 16 0 13 3 9 13 2 15 13 16 15 1 0 9 16 4 3 9 13 2 12 1 9 10 9 13 16 1 15 9 13 2
11 3 9 1 3 9 1 1 15 9 13 2
14 15 4 1 9 9 13 16 9 13 0 9 9 13 2
33 0 15 7 0 1 10 9 16 4 1 15 9 13 2 1 9 9 1 9 9 16 1 9 0 13 2 9 0 7 0 9 13 2
19 3 9 16 9 9 13 2 10 9 1 9 13 16 15 15 9 14 13 2
15 9 15 13 16 15 3 9 9 13 16 10 9 14 13 2
11 9 1 10 9 13 16 0 13 7 0 2
14 1 15 15 9 13 16 0 13 9 0 10 9 13 2
27 15 3 13 16 1 9 12 9 0 7 9 7 7 12 9 0 13 9 13 16 1 9 15 3 9 13 2
18 3 3 13 9 13 16 1 9 0 13 7 7 1 9 15 0 13 2
7 1 10 9 3 9 13 2
10 1 2 9 12 9 2 3 9 13 2
20 3 9 13 16 1 9 2 1 9 0 13 7 3 1 9 9 4 9 13 2
10 3 9 0 7 0 13 1 9 9 2
5 9 9 0 7 0
29 0 13 16 1 9 0 0 9 9 0 7 3 0 13 2 2 1 12 9 0 2 13 1 9 2 9 9 2 2
58 7 9 0 9 15 13 16 1 9 13 1 9 9 10 9 3 1 9 9 7 9 15 0 13 7 1 9 7 9 9 0 13 13 2 1 9 16 9 3 1 9 9 9 13 7 9 16 3 9 1 9 9 9 7 9 9 13 2
53 1 0 10 9 2 3 3 4 13 1 0 9 0 2 9 9 2 9 12 2 1 9 9 9 13 16 1 15 2 3 9 9 1 9 7 9 0 9 2 9 16 9 9 7 9 13 2 9 1 12 9 13 2
27 7 9 1 15 9 13 16 3 9 1 9 0 7 0 3 9 9 1 9 9 9 0 3 9 9 13 2
53 7 1 15 7 9 9 1 10 9 9 1 9 10 9 13 2 7 3 9 3 0 13 2 7 1 10 9 12 1 12 9 7 10 12 9 1 9 9 0 9 9 0 13 2 15 16 1 9 9 0 9 9 2
39 9 16 9 13 9 15 14 1 15 0 13 2 9 9 1 9 2 9 2 1 9 13 2 16 10 9 3 1 9 7 9 0 1 10 9 3 9 13 2
24 1 9 0 0 13 16 9 9 2 12 9 13 7 7 9 9 1 9 2 0 2 1 13 2
34 1 9 2 0 1 9 7 1 9 13 7 7 9 15 1 9 0 7 0 0 13 2 1 2 1 9 2 13 1 2 9 9 2 2
64 3 1 15 1 9 2 9 0 1 10 9 0 3 9 14 1 9 10 0 16 0 13 7 3 1 9 9 0 13 2 1 9 9 0 1 9 9 0 16 1 9 0 3 1 9 3 1 9 13 13 1 9 9 9 0 3 9 7 9 9 7 9 9 2
50 9 0 14 4 16 1 9 16 1 9 7 9 13 13 2 7 3 0 7 0 13 2 7 1 15 1 9 9 9 13 2 9 13 7 16 1 9 16 1 9 13 13 2 3 0 9 9 9 9 2
42 1 0 9 9 9 1 9 0 9 9 15 2 0 9 3 0 9 13 2 3 2 9 9 9 0 10 9 16 9 7 9 15 10 9 14 0 9 9 9 13 13 2
46 0 2 9 9 1 9 16 1 9 9 9 13 13 16 16 9 14 1 15 13 16 9 9 1 9 9 0 13 13 2 15 15 13 16 4 1 9 7 9 9 15 1 15 9 13 2
22 0 2 1 10 9 1 1 15 9 9 13 1 9 2 9 7 9 9 0 10 9 2
46 0 2 1 15 0 2 9 9 9 9 1 9 1 9 9 9 0 13 16 9 0 0 2 0 14 16 13 9 0 13 2 1 9 12 9 2 7 0 2 12 9 9 2 9 13 2
21 16 0 13 16 9 10 9 9 9 0 9 0 0 7 7 12 9 0 0 13 2
30 1 9 2 9 2 3 9 10 9 0 1 9 13 16 2 9 2 9 0 9 7 1 9 9 9 2 12 9 13 2
95 0 9 16 9 9 0 9 2 9 12 9 2 13 2 9 3 0 13 2 16 3 9 14 9 0 7 0 13 7 9 13 16 16 9 9 9 9 7 9 14 13 16 10 2 9 2 0 14 13 7 2 9 2 1 15 13 16 9 0 9 15 14 13 7 7 9 13 16 2 9 0 2 14 16 4 1 10 9 13 4 1 9 7 9 0 9 13 7 7 15 14 9 13 2 2
13 0 9 16 1 10 9 13 2 2 9 2 13 2
24 10 9 9 0 13 7 9 0 2 0 10 9 0 16 10 9 15 14 3 1 9 3 13 2
12 1 9 15 13 16 10 9 12 9 0 13 2
10 9 9 0 9 16 0 7 0 13 2
8 9 0 1 9 10 9 1 7
38 1 10 9 15 16 1 9 0 9 9 13 7 10 9 14 13 2 7 10 9 10 9 13 16 0 9 1 9 1 7 9 2 3 1 15 9 13 2
18 1 10 9 12 9 0 1 9 12 9 1 9 1 9 0 9 13 2
30 9 9 0 16 15 9 9 14 1 15 13 2 13 7 15 1 9 0 9 0 14 16 4 9 13 1 15 9 13 2
51 1 10 9 3 12 1 9 16 3 1 9 0 7 0 1 15 9 13 7 3 0 10 9 1 9 13 16 1 9 15 13 13 1 1 2 9 2 9 1 9 14 9 13 1 9 10 9 0 9 13 2
27 10 10 9 1 9 0 9 13 2 1 9 16 1 9 15 9 13 13 1 9 16 1 9 15 9 13 2
10 3 4 12 9 0 16 1 9 13 2
41 7 9 1 9 0 9 10 9 7 9 0 1 10 9 3 13 16 1 9 9 16 13 2 9 9 16 13 2 9 15 16 13 2 1 9 0 9 16 9 13 2
17 0 9 9 0 2 9 0 7 0 2 1 1 9 0 7 0 2
31 9 9 0 1 9 0 16 9 15 14 0 13 2 7 9 10 9 1 9 9 7 9 15 2 3 0 7 0 13 2 2
8 9 9 3 0 1 10 9 0
52 1 9 7 9 9 7 7 9 0 2 3 3 1 9 1 13 2 12 9 16 1 9 12 1 9 0 1 9 10 0 2 9 14 1 9 9 9 0 13 2 9 15 9 13 16 9 0 2 9 13 2 2
67 9 0 2 1 10 9 4 13 16 16 9 1 10 9 15 9 9 14 9 13 7 1 9 9 0 13 13 2 3 0 1 9 2 2 3 1 3 9 9 1 9 16 4 9 0 13 0 4 13 2 7 1 3 10 9 9 9 1 9 0 15 13 13 2 4 13 2
93 1 0 10 9 14 16 4 9 13 16 3 9 10 9 1 9 9 15 14 9 13 2 7 3 9 15 14 1 1 9 0 10 9 16 1 9 9 13 2 0 13 7 1 9 2 3 16 10 9 13 2 10 9 1 15 9 13 7 1 0 2 9 1 9 7 9 9 7 9 13 2 3 15 7 1 12 9 0 1 9 13 7 1 9 9 13 16 9 15 9 0 13 2
10 1 9 7 9 10 9 0 13 13 2
49 1 9 0 9 9 9 12 9 9 9 9 9 9 9 9 1 9 9 9 9 9 13 7 1 9 10 9 16 12 9 15 1 9 9 0 1 9 13 13 2 1 12 9 1 9 9 9 13 2
52 1 9 9 9 9 9 9 9 9 7 12 1 9 10 9 2 1 9 9 9 9 0 13 2 3 9 16 1 12 12 9 0 3 3 1 9 0 9 0 1 9 13 9 9 0 9 9 14 0 13 13 2
21 9 9 9 9 9 14 12 1 9 3 0 7 0 1 9 9 7 9 9 13 2
29 9 9 9 9 7 9 1 9 1 9 9 12 9 9 0 13 2 9 1 10 9 1 9 9 12 0 9 13 2
25 15 13 2 10 9 4 1 9 12 9 0 1 9 9 9 0 7 1 9 0 1 9 0 13 2
64 1 9 9 9 9 9 1 9 1 9 12 9 10 9 13 2 3 12 9 1 9 9 13 1 9 7 9 9 9 9 10 9 13 7 1 9 9 0 9 9 9 1 10 9 0 13 7 15 1 9 13 16 9 9 2 9 9 15 14 16 1 9 13 2
42 9 9 9 16 0 13 16 1 9 9 9 9 10 9 1 10 9 1 9 9 9 13 7 9 15 1 10 9 13 16 1 9 9 7 9 7 9 15 9 9 13 2
53 9 9 10 9 9 9 1 9 1 9 9 1 10 9 2 13 2 9 9 12 0 1 9 9 13 16 9 1 15 0 13 2 15 1 3 4 9 13 2 1 9 7 10 9 9 9 14 1 9 0 9 13 2
49 1 10 9 13 13 13 2 1 9 9 7 9 9 9 7 9 0 1 9 0 7 0 2 1 9 9 9 9 9 2 9 0 1 9 9 1 9 9 0 7 0 1 9 9 9 9 9 13 2
18 9 7 9 0 10 9 2 0 9 9 9 9 0 7 9 9 13 2
36 1 9 9 10 9 0 2 9 10 9 1 9 9 9 0 9 1 15 0 13 7 9 7 9 9 9 9 9 3 1 10 9 0 4 13 2
53 1 9 9 9 9 12 9 9 9 9 9 1 9 0 1 9 1 9 13 7 9 0 9 9 0 9 1 9 9 0 9 9 0 0 1 9 9 0 7 9 9 9 9 9 0 1 9 0 7 1 9 13 2
53 9 9 7 9 1 9 9 9 1 9 9 9 7 9 1 9 9 9 9 1 9 0 7 9 9 1 9 0 10 9 9 13 16 9 15 9 14 0 13 7 9 1 9 9 12 7 12 9 0 9 13 13 2
22 0 9 9 1 9 9 9 9 9 0 9 7 9 9 9 3 3 9 9 9 13 2
26 1 9 12 9 9 1 9 9 9 1 12 9 1 9 12 9 9 0 9 1 9 9 9 9 13 2
24 9 9 1 9 9 1 9 9 9 1 9 9 9 13 2 9 9 1 9 0 0 4 13 2
28 15 9 13 2 16 1 9 1 9 1 10 9 9 7 9 1 9 9 13 9 0 1 1 15 9 4 13 2
30 1 1 9 9 9 9 9 9 9 9 2 9 9 9 0 1 9 1 9 9 9 9 0 1 9 9 2 9 13 2
56 1 10 9 13 13 13 2 1 9 9 0 15 1 9 1 1 9 7 7 9 9 0 9 9 9 9 1 9 9 16 9 7 9 16 10 9 14 1 9 9 1 9 9 3 9 13 2 9 0 14 1 9 15 0 13 2
31 9 9 9 9 1 3 9 9 9 9 7 7 9 0 15 13 13 7 3 9 9 1 9 9 9 7 9 15 13 13 2
31 16 15 0 9 9 1 10 9 13 2 3 1 9 9 7 9 9 13 16 9 9 0 1 10 9 1 9 9 0 13 2
75 0 1 9 13 16 3 3 9 9 0 9 0 1 9 0 9 9 1 12 1 9 9 3 9 0 16 1 9 9 1 9 0 9 13 2 1 9 0 0 13 13 7 16 0 13 1 9 0 7 0 1 10 9 9 0 1 9 9 16 1 9 9 13 1 9 13 7 3 1 9 16 9 0 13 2
34 7 9 9 9 1 9 9 1 9 7 9 0 7 1 1 9 0 9 13 16 1 9 10 9 2 3 9 9 13 15 14 9 13 2
68 9 1 9 7 9 0 15 15 13 16 1 1 10 9 0 16 1 9 0 0 1 9 9 1 9 9 0 9 13 13 2 1 9 9 0 13 13 7 3 1 9 9 9 9 13 7 9 7 9 10 9 0 14 1 9 0 0 13 7 1 9 0 9 10 9 0 13 2
26 9 9 1 10 9 2 15 14 1 15 13 16 1 9 9 1 9 15 9 0 0 14 3 9 13 2
17 0 13 9 9 7 9 0 1 9 0 1 9 9 0 4 13 2
16 9 9 9 0 7 9 9 9 3 3 1 9 9 9 13 2
63 1 9 9 9 1 10 9 1 9 1 9 7 9 0 9 0 1 9 9 13 2 1 9 7 9 0 1 9 7 9 15 9 13 2 3 0 9 16 1 9 15 13 13 7 9 16 9 15 1 9 9 13 2 7 15 9 9 13 0 7 0 13 2
36 9 9 9 13 2 9 0 9 9 0 9 1 9 9 9 16 10 9 15 9 1 9 9 13 2 9 9 9 7 9 1 9 0 9 13 2
52 9 1 9 1 15 16 3 1 9 9 0 15 9 9 0 1 9 1 9 4 13 2 9 13 2 16 3 1 9 9 0 13 2 7 0 13 1 9 10 9 1 9 9 2 9 9 0 3 0 9 13 2
47 9 9 1 9 15 16 9 9 0 9 9 7 9 1 9 13 2 13 2 9 7 9 9 3 15 14 1 1 9 0 9 13 7 9 7 9 10 9 1 1 9 9 0 0 14 13 2
45 9 9 9 0 9 7 9 14 0 7 9 1 9 9 13 7 13 2 9 0 9 9 9 1 9 2 9 9 1 9 12 9 13 7 15 1 9 9 9 0 10 9 4 13 2
24 9 16 1 9 1 9 0 12 9 1 10 9 1 9 7 9 0 1 3 10 9 9 13 2
52 9 9 1 9 0 0 9 9 9 13 7 13 2 9 0 9 1 10 9 7 9 1 1 9 1 9 7 9 1 9 9 9 13 7 9 0 16 13 1 9 9 0 9 2 9 0 7 9 9 13 13 2
41 9 9 16 1 10 9 13 2 0 13 1 9 9 16 9 0 14 1 9 0 9 4 13 2 3 7 9 9 9 1 9 7 9 0 15 9 0 7 0 13 2
38 12 9 9 9 9 9 1 9 2 9 1 9 9 9 0 7 0 1 9 7 9 9 0 1 9 2 9 0 2 9 7 9 1 9 12 9 13 2
37 1 9 9 9 1 9 2 10 9 16 3 1 9 9 1 9 0 9 9 7 9 9 13 2 0 13 1 9 9 0 12 9 1 9 0 13 2
33 9 2 10 9 14 1 9 1 9 0 16 1 9 3 9 15 7 7 9 0 9 1 9 0 1 9 1 9 13 2 9 13 2
12 12 9 0 9 0 1 9 9 9 13 13 2
23 9 0 9 0 16 9 0 9 9 1 9 9 1 1 9 9 9 9 2 0 15 13 2
32 1 9 0 1 9 16 9 0 16 3 9 1 9 9 0 9 13 13 2 3 1 9 0 9 9 15 1 10 9 0 13 2
48 10 9 0 16 9 9 0 2 0 9 1 9 15 13 7 16 9 0 15 2 1 9 0 1 9 9 13 13 2 1 0 9 0 7 3 1 9 0 9 9 9 9 9 9 14 9 13 2
9 9 9 1 9 9 9 13 13 2
10 9 9 9 0 1 9 9 14 13 2
7 1 9 13 7 13 13 2
69 9 7 9 9 0 9 1 9 0 7 9 7 9 0 15 1 9 0 9 2 0 9 9 13 16 9 0 9 2 9 9 9 1 9 0 1 9 13 16 9 1 9 9 14 3 1 9 12 9 13 13 7 1 10 9 2 9 9 9 16 9 9 9 16 13 14 9 13 2
49 9 0 9 9 1 9 1 9 9 9 9 0 9 9 13 13 2 12 1 9 9 1 9 0 9 13 16 12 9 0 13 16 9 9 9 1 9 1 9 0 14 1 9 9 9 0 4 13 2
38 10 9 3 1 15 7 9 13 7 13 13 3 10 9 14 1 9 15 1 9 13 16 1 9 15 1 9 0 1 9 9 0 1 9 9 9 13 2
72 16 12 9 7 9 9 0 7 0 1 1 15 13 16 1 9 10 9 9 0 7 0 2 1 15 9 9 13 3 0 9 13 2 7 3 1 9 9 9 0 9 3 0 13 16 1 9 10 9 9 2 9 7 1 9 1 9 9 9 13 16 1 9 0 9 1 10 9 9 9 13 2
28 9 3 9 0 9 0 1 9 1 9 0 12 9 0 1 9 9 9 9 1 10 9 9 9 7 9 13 2
67 15 9 0 9 9 13 16 3 9 0 1 15 1 9 0 2 0 7 0 13 7 3 4 13 16 1 9 13 16 9 10 9 16 0 1 9 10 9 7 9 0 0 13 16 1 9 1 9 1 9 0 0 2 9 9 0 7 0 7 3 0 14 1 9 13 13 2
15 9 16 9 0 13 7 7 1 10 0 13 16 9 13 2
42 0 16 13 16 16 9 1 9 1 9 1 9 0 9 1 9 13 2 4 10 9 1 15 0 13 16 10 9 1 9 7 9 9 7 9 9 7 9 0 9 13 2
6 9 1 10 9 13 2
59 1 10 9 9 9 13 13 2 1 9 9 9 7 10 9 9 16 1 9 9 0 9 0 15 14 9 13 2 9 9 9 1 9 2 9 1 9 0 2 9 7 9 2 2 1 9 9 9 1 9 0 9 3 9 1 9 0 13 2
39 9 9 9 9 0 1 12 9 0 2 0 13 16 9 0 2 9 9 1 10 9 9 13 13 9 9 0 1 9 0 1 9 9 1 9 9 4 13 2
74 9 16 1 9 12 9 0 1 9 9 0 7 9 9 16 1 9 9 9 13 13 13 2 9 1 10 9 13 16 9 0 1 9 16 0 1 9 15 14 9 7 9 9 0 0 9 13 1 9 9 1 9 1 9 9 0 9 1 9 13 2 16 10 9 16 1 9 9 9 0 9 16 13 2
38 1 10 9 12 1 9 0 0 7 3 9 9 9 16 12 1 9 0 9 13 1 9 16 10 9 1 9 7 7 9 16 1 9 9 13 9 13 2
39 9 10 9 15 13 16 15 15 0 13 1 9 9 16 1 9 9 7 9 1 9 1 9 0 13 9 0 13 2 7 9 10 9 9 1 10 9 13 2
26 9 9 0 15 13 16 15 3 1 9 0 9 13 7 13 16 9 9 9 14 1 9 0 4 13 2
25 15 9 16 1 9 9 13 1 9 9 0 1 10 9 9 13 16 3 0 7 9 16 9 13 2
35 9 9 10 9 0 14 1 9 12 1 9 0 9 13 16 13 13 2 4 9 14 1 9 13 2 7 3 4 15 14 1 3 9 13 2
34 12 9 1 9 9 9 9 1 9 0 15 2 9 7 9 9 2 13 13 2 0 9 13 16 9 9 9 0 1 9 9 0 13 2
33 9 9 0 1 3 9 13 13 16 9 7 9 0 1 9 1 9 0 9 7 9 9 9 0 1 9 12 9 0 9 13 13 2
27 9 1 9 0 7 0 1 9 9 0 2 3 15 14 1 9 7 9 9 0 9 0 0 13 2 3 2
39 9 1 15 13 16 10 9 0 9 9 7 9 13 7 3 15 1 9 9 0 9 9 1 9 13 2 1 15 9 9 7 9 9 9 9 0 13 13 2
40 9 2 10 0 7 0 13 2 1 1 9 7 9 4 9 0 14 16 1 10 9 13 7 1 10 9 0 13 16 15 3 1 1 12 9 9 0 9 13 2
18 9 16 1 9 9 9 9 0 1 9 9 1 9 0 9 0 13 2
25 9 16 9 9 1 9 9 10 9 14 1 0 9 15 12 0 13 7 1 9 0 15 0 13 2
25 15 1 1 15 13 16 1 9 0 9 15 2 1 9 0 9 13 7 15 14 1 15 0 13 2
23 3 9 16 9 9 1 9 1 9 0 0 9 13 13 2 1 10 9 16 9 13 13 2
28 9 13 2 9 16 9 13 1 9 9 0 9 1 9 9 0 9 13 9 0 13 2 9 15 14 9 13 2
32 9 16 16 1 9 0 0 9 9 13 7 1 9 9 9 9 0 7 0 1 9 13 10 9 14 13 2 3 1 9 0 2
12 1 10 9 3 10 12 9 9 1 9 13 2
48 1 9 13 4 1 9 9 9 9 14 1 9 15 9 15 13 7 1 9 0 1 10 9 9 0 13 16 9 9 0 1 0 9 0 15 0 13 10 9 7 9 14 1 3 9 15 13 2
116 9 9 9 0 15 14 1 9 1 9 2 12 9 9 0 1 9 2 9 13 16 9 1 15 14 1 1 13 2 9 0 9 1 9 9 9 9 2 9 7 9 9 0 9 1 9 9 9 1 9 9 0 1 9 1 12 9 0 1 9 9 7 9 0 1 9 7 9 15 1 9 13 13 13 16 0 9 9 0 9 1 9 0 7 0 1 9 9 0 1 9 9 1 13 7 3 3 1 9 9 9 1 9 2 9 0 9 7 9 9 0 9 9 13 13 2
86 1 9 9 9 2 9 0 7 0 1 9 7 9 9 0 9 15 13 16 9 1 9 0 1 9 9 0 9 0 1 9 0 14 0 1 9 2 9 2 9 9 0 2 9 1 9 9 9 15 7 0 9 9 0 1 9 0 7 9 9 9 13 7 1 9 0 0 9 9 9 7 7 9 7 9 0 15 3 9 9 9 9 7 9 0 2
23 9 9 9 9 7 9 9 9 9 16 9 9 0 9 7 9 0 9 14 9 9 13 2
85 9 7 9 1 9 0 9 0 1 9 9 2 9 7 9 9 0 1 10 9 9 7 9 9 7 9 0 7 0 1 9 0 7 3 9 0 0 1 9 9 0 9 15 9 15 13 16 9 0 1 9 0 9 9 0 1 9 7 9 9 1 9 2 16 3 13 1 9 9 0 1 9 12 9 9 9 0 9 14 0 13 2 9 13 2
35 0 10 9 2 9 9 9 0 12 9 13 16 1 15 9 1 9 2 9 9 7 9 9 0 7 9 9 9 0 7 0 9 13 13 2
38 1 10 9 16 9 9 0 2 9 0 9 2 9 9 2 9 9 7 9 9 0 9 7 9 1 9 9 15 9 13 2 12 9 1 9 0 13 2
21 9 9 16 1 9 0 9 0 1 9 9 1 9 7 1 9 9 9 0 13 2
36 9 16 9 13 1 9 10 9 0 13 16 9 1 9 9 0 1 1 9 0 7 9 15 7 9 9 13 7 1 9 9 9 15 13 13 2
44 9 9 9 0 16 0 7 1 12 9 0 1 9 9 0 0 16 0 13 9 12 0 9 9 1 9 9 0 2 9 2 9 7 9 9 7 9 3 1 9 9 13 13 2
41 9 9 1 9 2 9 0 7 9 9 0 2 13 13 2 9 9 9 0 1 9 9 9 0 7 9 0 9 0 1 9 15 2 9 14 1 9 0 0 13 2
47 9 15 13 16 9 9 1 10 9 7 9 9 13 13 2 0 9 7 9 0 7 0 9 0 1 9 9 7 9 9 15 7 0 1 15 9 7 9 16 1 9 0 9 13 2 13 2
8 1 10 9 9 0 0 13 2
34 9 9 0 1 9 0 4 0 7 0 13 7 1 9 9 7 9 9 0 1 9 9 2 9 14 1 9 9 1 9 15 9 13 2
16 9 10 9 1 9 9 0 7 7 9 0 7 0 9 13 2
35 16 10 9 1 1 9 9 0 0 9 13 13 16 9 9 0 15 13 13 9 0 9 0 9 9 1 9 9 0 1 9 9 15 13 2
50 3 9 0 1 9 9 9 9 1 9 1 9 9 10 9 1 9 9 1 9 0 1 9 1 9 9 0 2 9 4 13 7 9 0 1 9 9 9 10 9 1 9 1 9 1 9 9 9 13 2
36 4 9 13 1 9 9 2 0 1 9 0 9 0 15 14 1 9 13 7 1 3 9 1 9 9 9 16 1 10 9 0 9 13 2 13 2
20 9 1 9 15 13 16 9 0 1 9 0 3 13 9 10 9 14 0 13 2
44 1 10 9 9 0 1 9 2 1 9 0 9 1 9 0 9 0 13 7 3 1 9 16 1 9 15 9 7 9 0 9 13 2 0 15 7 4 15 14 1 12 9 13 2
30 3 9 0 0 13 1 9 9 1 9 9 0 2 9 14 1 1 9 9 0 13 7 15 14 1 9 15 0 13 2
52 9 9 9 0 10 9 14 9 13 16 9 0 1 9 0 7 0 1 9 0 2 9 0 7 0 1 9 9 0 9 13 7 9 0 7 0 1 9 9 0 1 1 9 9 7 9 0 1 9 0 13 2
23 9 9 9 13 1 9 9 9 16 1 15 9 0 9 9 15 14 1 9 0 9 13 2
8 9 9 9 9 9 0 13 2
49 16 10 9 0 7 0 9 1 9 0 9 7 3 3 1 0 9 0 1 9 9 9 13 2 7 9 0 15 1 9 9 15 1 0 9 9 0 9 7 9 0 1 9 9 1 9 13 13 2
9 9 0 9 1 10 9 0 13 2
28 9 1 9 9 15 3 1 9 9 9 1 9 1 15 13 13 7 15 1 3 1 9 9 1 9 9 13 2
13 1 10 9 9 9 9 9 15 14 1 9 13 2
79 10 9 16 0 13 7 1 9 1 15 7 15 1 9 12 9 1 9 9 9 9 1 9 9 9 0 9 13 7 1 9 15 9 9 9 9 0 1 0 9 0 1 9 7 9 0 13 9 15 14 1 1 9 0 9 7 9 0 9 9 9 9 9 9 9 7 9 15 1 9 0 1 9 7 9 3 9 13 2
70 1 10 9 9 13 1 9 16 9 1 3 9 1 9 0 13 9 1 9 0 7 9 9 15 13 7 3 1 9 15 3 1 10 9 0 9 7 9 0 7 0 9 9 1 9 13 13 16 3 0 10 9 7 9 14 1 1 13 7 9 9 14 0 1 9 7 9 13 13 2
18 10 9 3 1 9 9 7 9 0 13 13 7 10 9 16 3 13 2
61 15 9 13 9 16 1 10 9 3 0 13 7 9 13 2 12 9 7 9 9 13 2 13 1 1 9 0 9 9 9 15 14 9 13 7 3 1 9 0 1 9 0 9 9 0 1 9 9 9 7 9 0 1 15 1 1 9 9 9 13 2
27 9 13 9 7 9 1 9 9 9 13 16 10 9 7 10 9 9 9 12 12 9 9 9 3 9 13 2
39 15 1 9 13 2 3 12 9 3 1 9 9 1 9 9 1 9 0 9 13 7 1 9 15 7 9 7 9 15 0 1 9 0 7 9 9 9 13 2
32 9 15 9 13 16 9 7 9 7 9 1 3 9 7 9 0 13 2 3 10 9 7 10 9 2 3 10 9 7 9 0 2
16 4 9 14 1 9 9 7 9 9 13 3 9 9 7 9 2
23 4 9 13 16 9 9 7 9 1 9 15 13 16 9 9 7 15 1 10 9 9 13 2
26 15 4 15 14 0 1 15 13 16 9 13 15 13 7 7 9 15 13 2 16 9 9 7 7 9 2
10 15 12 1 9 0 0 9 16 13 2
43 10 9 7 0 13 3 9 0 1 12 9 0 12 9 7 9 16 3 0 1 0 9 13 14 9 13 2 1 9 7 1 9 15 3 9 3 1 9 9 0 0 13 2
25 16 10 9 9 0 9 0 7 1 10 9 9 7 9 1 9 1 9 9 7 9 7 9 13 2
12 1 9 9 9 15 14 1 10 9 9 13 2
34 9 0 9 9 13 16 9 9 9 1 9 7 7 9 13 7 9 9 9 1 9 9 13 7 4 13 16 10 9 9 9 0 13 2
13 9 13 13 0 9 9 1 9 9 0 0 13 2
18 10 9 9 0 9 14 9 13 7 9 9 9 7 9 14 9 13 2
62 9 0 15 13 16 16 9 3 9 13 1 9 9 1 15 9 13 7 7 16 9 7 9 1 10 9 9 13 9 13 2 7 9 0 9 7 9 0 9 1 12 9 10 9 14 1 9 15 1 9 13 16 9 0 0 13 9 10 9 13 13 2
13 15 15 13 7 13 7 3 9 7 9 9 13 2
9 9 3 9 0 1 9 9 13 2
15 1 9 1 12 12 9 7 0 15 1 0 9 9 13 2
24 1 1 9 0 0 10 9 7 9 9 9 7 9 9 7 7 10 9 7 10 9 9 13 2
6 9 9 7 9 9 2
62 9 9 16 9 1 9 9 9 9 9 14 1 9 9 9 1 10 9 9 13 13 2 9 9 9 9 0 2 13 2 9 9 0 9 9 13 16 1 9 9 0 1 9 0 9 9 0 3 1 15 13 7 15 1 9 9 9 9 1 9 13 2
38 9 9 1 13 7 13 1 9 13 2 9 15 13 16 9 15 14 9 13 7 1 9 9 13 2 9 10 9 13 16 1 9 12 9 9 15 13 2
23 15 13 2 15 9 13 16 1 1 9 9 13 1 9 7 9 0 1 1 9 9 13 2
30 15 13 1 9 0 13 2 16 3 9 10 9 14 16 13 2 1 9 7 15 13 1 9 7 13 7 13 9 13 2
71 9 1 9 2 9 7 9 9 9 1 9 1 9 9 9 0 9 1 9 9 0 14 0 13 7 9 13 2 15 9 13 2 7 9 14 1 9 9 13 16 1 9 0 15 1 9 9 2 9 2 9 1 9 12 9 0 7 9 9 9 0 9 13 7 1 10 9 0 16 13 2
28 9 9 13 2 3 1 9 12 9 9 1 9 0 9 7 9 9 0 13 16 10 9 1 9 15 0 13 2
49 1 3 9 16 9 1 9 9 9 14 13 9 13 9 0 14 1 9 0 1 9 13 7 1 3 7 9 9 1 9 9 0 7 9 9 1 9 9 9 13 1 10 9 1 9 9 0 13 2
43 9 9 9 9 0 1 9 1 9 1 0 9 10 9 1 9 9 0 9 1 9 9 9 9 3 1 9 9 9 7 9 0 9 13 2 3 9 9 9 3 0 13 2
7 0 9 15 9 9 13 2
25 0 1 12 9 13 16 10 9 0 0 2 1 9 9 13 13 7 15 14 16 1 15 15 13 2
28 9 15 14 16 13 9 2 3 13 16 1 9 9 16 10 9 14 13 7 10 0 0 14 1 9 0 13 2
37 1 9 12 9 1 3 9 15 14 1 9 13 2 10 9 12 9 2 9 7 9 7 9 2 9 10 9 14 13 7 3 1 9 9 9 13 2
19 9 16 16 13 2 13 2 15 15 1 9 13 16 3 1 9 9 13 2
6 16 13 2 9 9 2
29 1 10 9 7 9 7 3 9 0 16 9 13 1 9 15 13 7 13 13 2 9 15 3 9 9 13 7 13 2
10 15 3 14 1 9 15 13 10 0 2
19 15 15 12 9 9 1 9 13 2 12 9 13 6 13 3 3 13 2 2
23 3 7 7 13 9 15 13 2 13 1 9 0 9 13 7 13 2 6 15 7 7 7 2
12 16 13 12 9 7 12 9 4 9 13 3 2
32 3 12 9 13 2 12 9 7 12 9 16 3 13 13 1 9 15 2 7 1 3 16 9 15 1 9 10 9 13 2 13 2
5 13 2 9 9 2
8 13 2 15 0 13 9 13 2
23 1 9 15 9 13 2 3 1 9 13 2 9 9 15 9 15 13 2 9 13 10 9 2
33 0 9 0 1 15 13 2 9 15 15 7 9 15 14 0 9 13 7 13 2 2 0 12 7 9 1 9 9 0 12 9 13 2
7 15 9 13 2 15 13 2
5 9 13 9 9 2
5 15 4 9 13 2
33 10 3 9 2 1 9 15 2 12 9 0 9 13 7 13 2 9 12 9 13 1 9 2 12 9 1 15 13 2 12 9 13 2
8 13 10 9 12 0 13 13 2
8 3 15 10 9 12 0 13 2
8 0 12 9 0 16 3 15 2
20 3 2 9 9 15 16 16 0 9 0 13 2 1 9 0 3 12 0 13 2
12 10 9 15 12 9 13 2 10 9 0 13 2
13 9 13 1 0 2 12 9 9 13 16 9 13 2
4 6 9 2 2
3 9 13 2
9 10 9 1 9 15 9 15 13 2
15 1 15 15 9 1 13 2 13 16 12 9 0 9 13 2
15 12 9 0 13 2 0 9 0 13 9 14 13 1 9 2
22 12 9 0 1 10 9 13 2 7 13 1 9 15 16 9 0 7 0 15 9 13 2
5 9 15 9 13 2
6 13 2 9 9 9 2
7 15 3 9 15 9 13 2
8 9 15 0 2 9 15 0 2
11 3 9 13 1 10 9 9 1 9 13 2
7 9 9 1 9 9 13 2
30 9 9 0 9 9 0 9 3 9 13 2 9 9 9 9 1 9 3 1 1 9 0 9 0 12 9 9 13 13 2
35 9 9 13 2 1 9 3 3 12 12 7 12 12 9 9 1 9 9 13 16 10 9 1 9 3 1 12 12 7 12 12 9 13 13 2
36 15 13 2 1 9 7 9 15 9 9 0 3 9 9 2 9 0 7 9 9 13 2 7 1 9 9 1 9 9 3 3 0 1 9 13 2
46 15 1 9 9 9 9 1 9 14 9 9 9 10 9 0 9 13 7 13 2 9 9 1 9 1 9 12 1 1 9 12 0 12 9 9 13 16 0 1 9 0 9 15 13 13 2
26 9 13 2 9 13 1 9 3 9 9 9 1 9 1 1 12 12 9 1 9 13 16 3 3 13 2
40 15 9 9 9 0 1 3 1 9 14 3 12 12 9 0 9 9 0 9 13 7 13 2 0 9 0 0 1 9 0 1 9 1 12 12 9 1 9 13 2
29 15 16 13 2 1 9 9 9 9 16 12 9 9 13 2 16 1 9 9 2 9 7 9 7 9 9 13 13 2
57 9 9 0 9 9 0 9 13 2 1 9 9 1 9 9 9 9 9 9 0 1 9 9 9 9 9 13 7 1 9 10 9 9 9 0 9 9 13 7 1 9 9 1 9 9 9 7 7 1 9 9 9 0 9 9 13 2
31 15 13 2 1 9 9 9 9 9 9 2 9 1 9 9 1 9 9 1 9 9 9 1 9 9 9 1 9 9 13 2
42 9 9 9 9 9 9 1 9 0 1 9 0 9 0 1 9 9 9 13 1 9 9 0 9 9 1 9 7 9 9 9 9 9 0 9 9 9 9 9 4 13 2
35 1 9 9 0 9 9 9 9 9 9 1 9 0 1 9 0 9 13 2 0 1 9 1 9 9 13 7 10 9 9 0 14 9 13 2
47 9 9 9 1 9 1 10 9 16 16 10 9 9 0 9 9 4 13 7 3 13 2 1 9 0 4 1 9 9 16 9 4 13 9 13 7 9 2 9 9 1 9 7 9 9 13 2
34 9 9 1 9 9 9 0 9 9 13 2 1 9 0 4 9 9 13 7 10 9 7 9 13 4 9 9 1 9 9 1 9 13 2
18 1 9 9 3 9 3 13 2 3 1 9 7 9 9 1 9 13 2
60 9 9 9 1 9 1 10 9 16 16 9 9 9 9 1 9 12 9 9 0 9 9 4 13 7 3 13 2 15 1 9 0 1 9 0 13 9 0 9 7 9 9 9 9 0 1 9 0 9 13 7 9 10 9 9 14 0 4 13 2
59 9 9 1 9 9 10 9 1 1 15 16 9 9 13 1 9 9 9 9 9 9 1 9 12 0 9 13 2 13 2 10 9 7 9 0 13 7 9 13 7 10 9 7 9 13 9 9 0 1 9 0 7 10 9 9 9 9 13 2
37 9 9 9 1 9 1 10 9 16 16 1 9 0 13 9 7 9 9 9 14 9 13 7 3 13 2 9 9 0 13 7 9 9 16 9 13 2
63 9 9 9 1 9 9 9 9 1 1 15 16 12 9 16 1 9 9 9 9 13 13 2 13 2 15 9 13 16 9 1 9 0 13 7 9 7 9 13 7 9 16 1 9 9 9 9 13 2 9 7 9 7 9 16 0 13 7 9 0 9 13 2
66 9 9 9 1 9 1 10 9 16 3 9 9 9 9 0 1 9 9 13 13 2 13 2 10 9 1 9 9 16 0 9 7 9 13 2 9 9 1 12 9 7 1 12 9 0 13 7 12 9 1 3 1 12 9 14 15 16 1 12 9 4 9 1 9 13 2
40 9 0 1 9 0 1 12 9 9 0 13 2 9 9 15 16 0 13 7 9 9 7 9 0 16 0 13 2 7 1 10 9 1 9 0 4 9 0 13 2
45 9 9 9 1 9 1 10 9 16 16 9 0 1 0 9 1 9 9 9 9 4 13 7 3 2 13 2 1 15 9 0 13 7 15 0 13 16 9 1 9 3 0 9 13 2
34 10 9 1 9 9 9 13 2 3 1 10 9 9 0 16 1 9 0 13 16 9 9 9 0 7 9 12 0 9 1 9 15 13 2
43 9 9 9 1 10 9 16 1 9 9 9 0 9 9 9 0 1 12 9 13 1 9 0 10 9 0 9 9 9 2 9 2 3 1 9 9 9 12 7 9 9 13 2
14 9 9 7 9 15 1 10 9 12 1 12 0 13 2
19 3 1 9 9 9 2 9 2 9 1 9 1 9 1 9 9 9 13 2
6 9 9 9 15 13 2
24 1 9 15 1 9 9 2 9 2 9 13 7 9 13 16 0 9 9 9 2 9 2 13 2
15 9 9 16 9 13 7 9 9 0 9 9 14 9 13 2
25 7 15 7 15 0 9 9 9 2 9 2 13 7 1 9 16 3 0 13 7 1 15 9 13 2
25 10 0 9 1 3 9 9 9 9 2 9 2 1 9 12 7 1 3 1 9 7 9 9 13 2
12 9 15 14 1 9 7 9 1 9 9 13 2
14 7 13 1 9 16 9 0 13 10 9 14 9 13 2
17 16 9 13 10 9 9 9 2 9 2 9 13 16 9 4 13 2
32 9 2 9 7 9 9 16 7 10 9 9 7 9 14 9 7 9 13 2 9 7 9 7 9 7 9 14 1 9 9 13 2
17 9 9 1 9 9 2 9 2 13 7 9 13 16 9 9 13 2
31 9 9 2 9 2 1 9 1 0 9 9 7 9 13 2 15 1 9 9 13 16 9 14 16 9 0 13 13 9 13 2
29 3 9 9 2 9 2 9 13 16 16 9 15 9 1 9 9 13 2 9 9 0 9 7 9 1 15 9 13 2
25 3 9 7 9 1 10 9 13 7 13 16 9 9 3 9 0 13 7 9 14 1 9 0 13 2
24 3 16 9 13 1 10 9 9 9 2 9 2 1 9 7 9 7 9 7 9 9 0 13 2
20 1 15 9 2 9 2 1 9 9 2 9 2 9 14 9 13 7 9 13 2
54 9 9 13 13 16 1 9 9 1 0 1 12 12 9 9 2 9 2 14 9 13 16 9 9 9 9 1 9 1 10 9 7 9 9 16 9 9 2 9 2 9 9 9 7 9 9 13 1 10 9 9 13 13 2
18 1 3 9 0 0 9 9 2 9 2 9 10 9 15 14 9 13 2
20 9 9 16 1 9 9 1 9 9 9 0 13 13 2 1 9 9 9 13 2
20 1 9 8 9 2 9 2 16 1 1 15 13 13 13 2 9 15 3 13 2
4 13 2 9 2
8 13 2 9 9 15 3 13 2
4 13 2 9 2
7 9 13 2 9 7 9 2
26 16 9 8 9 2 9 2 9 14 1 9 9 9 13 2 9 9 2 9 2 13 2 6 1 15 2
13 16 12 9 16 13 13 9 10 15 14 9 13 2
9 10 9 9 9 7 9 9 13 2
54 1 9 16 3 9 9 1 9 7 9 9 13 7 0 13 16 9 0 9 13 9 15 14 9 9 13 2 9 9 1 9 9 15 7 7 12 9 3 9 0 15 2 9 9 2 10 9 0 7 0 14 9 13 2
28 9 16 9 0 9 7 9 1 9 15 9 13 13 2 9 9 16 1 9 9 9 2 9 0 9 13 13 2
14 3 9 16 1 9 9 2 9 2 1 9 13 13 2
6 9 0 10 9 13 2
13 1 9 9 7 9 9 9 10 12 9 0 13 2
11 9 1 9 9 2 9 2 9 13 13 2
10 9 1 10 9 9 14 0 13 13 2
24 10 9 1 9 10 9 2 1 9 15 13 7 13 2 3 1 10 9 9 1 9 13 13 2
5 9 10 9 13 2
9 3 1 10 9 9 0 13 13 2
3 1 13 2
6 9 15 7 15 13 2
11 1 10 9 12 9 0 7 9 9 13 2
11 7 9 9 16 9 7 9 13 9 13 2
60 9 10 9 16 13 9 9 9 2 9 2 14 9 9 1 9 13 16 1 9 9 9 9 2 9 2 9 7 9 9 3 9 13 7 9 13 2 16 3 9 9 2 9 2 13 7 1 9 13 2 16 9 13 1 9 13 15 9 13 2
14 1 1 9 9 2 9 2 16 9 9 14 9 13 2
14 9 0 9 16 16 9 9 9 13 7 7 9 9 2
30 9 1 9 16 9 9 13 7 9 15 1 9 2 9 13 16 9 9 16 9 9 9 9 13 14 1 9 9 13 2
23 9 9 14 1 9 1 9 13 2 9 13 2 9 7 9 9 15 9 2 9 2 13 2
5 1 9 9 13 2
12 9 1 9 9 13 16 3 7 3 4 13 2
23 10 9 9 15 13 7 15 7 10 12 9 9 7 9 2 1 10 9 9 15 0 13 2
16 1 9 9 9 13 16 9 13 7 10 7 2 8 8 8 2
24 9 1 9 14 16 1 9 9 0 13 13 1 9 13 2 7 15 7 9 9 9 4 13 2
16 9 9 2 9 2 10 9 0 1 9 14 12 12 9 13 2
22 13 9 9 15 0 9 16 1 9 15 13 7 9 9 9 13 2 9 12 9 13 2
21 1 3 1 1 9 1 9 15 9 13 13 16 9 9 15 14 9 9 13 2 2
12 15 9 13 16 1 9 9 1 15 9 13 2
9 7 1 9 9 1 15 9 13 2
9 10 9 16 9 3 9 4 13 2
18 9 16 0 1 9 7 9 9 7 9 9 13 9 14 9 13 13 2
8 9 1 9 9 9 0 13 2
12 15 16 1 9 3 9 13 2 3 16 13 2
15 10 9 1 9 9 13 7 1 9 15 7 9 15 13 2
57 3 1 9 0 1 10 9 16 9 9 9 0 13 13 2 9 9 2 9 2 13 2 15 9 13 16 15 9 9 9 14 1 9 9 15 9 8 9 8 9 1 9 12 9 7 1 1 15 9 16 15 15 1 9 13 13 2
14 9 16 1 9 13 7 9 15 9 12 12 9 13 2
11 9 13 2 15 6 9 1 15 9 13 2
46 0 13 9 9 2 9 2 3 9 7 1 9 13 16 12 9 9 7 9 0 13 2 7 9 1 9 9 7 9 15 13 16 1 9 9 9 9 1 9 9 7 9 9 9 13 2
49 1 9 1 9 0 16 9 13 9 9 12 9 13 7 9 7 3 9 0 0 13 2 9 16 0 9 13 2 13 9 9 7 9 9 14 1 9 9 13 16 3 9 7 9 1 1 9 13 2
42 9 9 1 9 9 9 9 7 9 16 1 3 3 1 9 9 2 9 2 0 9 9 13 1 9 9 0 13 2 16 9 9 2 9 2 10 9 14 1 15 13 2
36 9 0 9 13 16 9 9 2 9 2 1 9 12 10 9 2 9 0 3 13 13 9 15 14 1 1 9 9 7 7 9 9 9 13 13 2
13 9 9 9 2 9 2 0 1 1 9 9 13 2
6 9 14 1 9 13 2
13 1 9 13 16 9 1 9 15 9 0 13 13 2
8 1 9 13 2 12 9 13 2
13 7 15 7 9 7 9 1 1 9 0 9 13 2
32 0 15 7 9 1 9 9 9 2 9 2 9 13 2 10 9 9 9 2 9 2 2 9 9 9 7 9 14 1 9 13 2
14 7 15 7 10 9 14 1 9 9 2 9 2 13 2
32 16 1 15 1 10 12 9 9 13 2 9 0 9 4 13 7 9 9 2 9 2 9 14 1 9 9 2 8 8 2 13 2
27 9 13 2 16 1 9 9 13 15 16 1 15 13 1 9 15 1 9 15 7 1 1 9 15 9 13 2
7 9 0 15 14 9 13 2
36 12 9 9 9 9 13 7 3 9 1 9 0 7 9 9 13 7 1 9 16 9 9 4 9 1 9 9 13 7 10 9 1 9 9 13 2
48 12 9 1 9 9 16 1 9 12 1 9 9 1 9 9 13 2 9 9 1 13 7 13 1 9 2 9 15 1 10 9 14 9 0 13 7 9 3 0 15 1 9 14 1 9 9 13 2
52 10 9 16 1 15 9 9 9 9 9 7 9 0 7 9 9 9 9 9 9 16 9 13 2 9 9 15 1 9 1 0 1 9 9 13 7 9 13 16 1 10 9 2 15 1 9 9 0 16 9 13 2
33 9 9 9 9 16 1 10 9 9 13 2 13 2 9 16 15 1 9 1 9 9 0 15 0 13 2 3 0 7 0 0 13 2
50 16 9 9 9 2 9 0 13 7 3 16 1 12 9 3 2 9 1 9 9 9 7 9 1 9 1 15 9 13 13 16 3 13 1 15 9 13 7 3 12 9 1 9 0 1 10 9 9 13 2
32 9 9 2 13 2 9 9 1 9 9 9 2 12 9 0 7 0 13 7 1 15 2 3 9 1 9 7 9 1 9 13 2
45 9 9 2 13 2 0 9 13 7 13 1 10 9 2 1 9 0 9 9 9 9 13 16 1 9 15 2 9 7 9 9 13 7 1 15 2 3 9 0 7 7 0 9 13 2
35 15 1 9 9 1 9 9 10 9 0 2 13 2 3 9 16 1 10 9 7 9 13 9 13 2 9 0 7 9 9 0 1 9 13 2
33 9 9 2 9 13 2 15 1 9 9 9 9 9 16 15 14 9 9 7 9 12 9 13 2 13 10 9 0 7 0 14 13 2
58 9 9 9 9 16 16 1 10 9 9 13 2 10 9 0 14 0 13 7 13 2 9 16 1 10 9 1 1 9 9 0 13 2 0 0 13 7 9 9 1 9 9 0 7 9 9 15 1 9 9 0 15 2 0 7 0 13 2
34 9 9 13 2 16 15 3 1 10 9 13 9 0 1 9 14 9 13 7 9 13 16 9 1 3 1 9 9 3 0 16 9 13 2
55 15 1 9 1 10 9 16 9 9 10 9 1 9 7 9 0 15 3 9 1 9 0 13 2 9 9 13 16 9 1 9 1 9 0 7 9 0 9 0 1 9 0 13 7 9 7 9 15 14 9 9 9 15 13 2
26 9 2 1 0 9 1 9 9 2 9 15 9 9 9 9 0 9 3 1 9 9 0 14 0 13 2
32 9 9 9 16 3 1 9 0 9 13 7 1 9 9 0 13 2 1 0 9 9 9 9 1 9 9 9 0 1 15 13 2
30 1 1 9 9 1 9 9 16 1 9 9 0 9 13 9 9 10 9 1 12 1 12 9 9 1 12 9 9 13 2
20 3 1 0 9 9 9 0 9 2 12 9 0 0 1 9 1 9 9 13 2
42 9 9 0 9 0 9 10 9 14 9 0 9 2 9 0 9 9 9 2 9 12 9 2 9 0 9 9 2 9 9 9 9 2 9 9 7 9 9 9 9 13 2
20 9 9 9 9 9 13 2 9 10 9 0 0 12 12 9 9 1 9 13 2
19 15 16 13 2 1 9 12 9 0 1 9 9 3 12 9 15 0 13 2
29 15 9 9 10 9 14 12 9 9 13 7 13 2 10 9 9 12 12 7 12 9 9 14 1 9 9 9 13 2
27 1 9 0 9 12 9 0 7 9 1 9 9 2 9 2 9 2 9 2 9 2 9 7 9 9 13 2
18 9 9 9 9 1 9 9 0 0 1 12 12 7 12 9 9 13 2
15 9 9 10 9 1 9 9 0 9 9 7 9 9 13 2
32 7 1 9 9 9 9 9 9 9 9 12 9 9 1 9 9 9 9 1 9 9 9 13 13 16 9 0 2 0 16 13 2
29 9 7 9 1 9 9 3 1 9 0 9 7 9 9 0 2 9 1 12 9 9 7 9 1 9 9 0 13 2
37 1 9 9 0 9 9 0 9 2 9 9 7 9 16 12 9 1 9 0 9 13 2 10 12 1 9 9 1 9 0 1 9 9 7 9 13 2
28 10 9 1 9 0 9 12 7 3 1 9 9 0 9 12 7 9 9 9 0 1 9 9 9 9 9 13 2
20 9 1 9 9 9 1 1 9 9 2 9 0 9 14 16 1 15 13 13 2
17 9 7 9 0 7 0 1 9 9 7 1 9 9 3 9 13 2
39 9 7 9 9 0 1 9 12 9 0 13 16 9 10 9 1 9 0 1 9 9 12 9 1 15 1 0 9 9 9 0 1 0 1 9 0 0 13 2
9 9 16 9 1 9 9 9 13 2
26 9 16 1 9 0 1 10 9 9 0 7 9 1 9 1 9 13 2 3 1 9 9 0 9 13 2
36 9 9 0 16 1 12 9 9 7 1 0 9 9 4 13 9 1 9 7 9 0 7 9 9 9 0 16 1 9 9 9 9 0 4 13 2
22 9 9 0 1 0 9 0 9 9 1 9 2 1 9 9 7 9 9 9 13 13 2
22 1 10 9 9 12 9 1 9 9 9 2 9 9 7 9 0 0 9 9 9 13 2
22 1 9 9 9 10 9 16 9 9 0 1 9 9 9 1 9 1 9 1 4 13 2
41 10 9 1 9 12 9 9 1 9 9 1 9 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 7 9 1 0 9 9 9 1 9 13 13 2
30 9 9 16 1 9 9 0 1 10 9 9 13 2 9 9 1 9 9 9 15 1 12 9 9 7 9 0 9 13 2
22 15 1 10 9 1 1 9 0 9 9 1 9 0 2 0 7 0 9 14 9 13 2
44 1 10 9 12 1 9 9 9 2 1 9 1 9 0 1 9 9 9 0 7 0 0 2 9 9 13 16 9 0 1 9 9 0 0 15 2 3 1 9 9 9 0 13 2
18 0 9 9 0 0 1 9 9 9 0 1 9 9 9 9 0 13 2
50 1 10 9 9 0 9 1 9 9 0 1 9 9 2 9 2 9 2 9 7 9 0 9 0 7 0 2 9 2 9 0 2 9 2 9 2 9 7 9 9 7 9 9 0 7 0 0 9 13 2
25 10 9 1 9 9 0 9 0 1 9 9 1 9 7 9 0 9 9 0 9 7 9 9 13 2
6 9 1 9 9 1 9
29 9 9 9 9 1 9 9 9 9 9 0 9 1 9 2 9 7 9 9 9 9 1 9 14 1 1 13 13 2
31 1 9 0 16 9 0 1 9 0 9 9 9 1 9 1 9 1 13 13 2 3 9 1 9 9 1 10 9 9 13 2
46 1 9 9 9 16 1 9 9 0 9 0 9 1 9 0 13 2 9 1 9 9 2 9 9 2 9 9 2 9 9 2 9 9 7 0 9 0 1 9 0 1 9 13 13 13 2
38 9 9 9 9 9 9 1 1 9 0 1 1 9 1 9 9 0 1 10 9 0 13 2 10 0 9 13 16 9 3 9 1 12 9 9 0 13 2
28 15 13 2 9 10 9 9 7 9 1 9 1 9 1 0 1 10 9 0 2 0 7 9 9 9 9 13 2
21 1 9 0 9 1 9 0 1 9 9 1 9 0 15 14 1 9 9 9 13 2
30 7 9 0 9 16 16 1 9 0 13 2 9 1 9 0 15 14 1 9 9 9 2 9 7 9 0 0 9 13 2
12 9 9 9 0 9 1 9 3 1 9 13 2
10 9 0 1 9 0 1 9 13 13 2
37 9 0 1 9 9 9 9 0 16 1 9 12 9 3 0 9 9 9 9 9 13 2 3 1 9 9 0 1 9 9 1 9 9 9 9 13 2
41 1 9 9 0 9 9 0 2 9 9 0 0 2 9 0 9 0 9 7 9 2 9 0 0 2 9 2 9 7 9 0 1 9 9 13 16 1 9 13 13 2
38 10 9 16 1 9 9 15 0 9 12 9 9 13 2 0 9 1 9 12 1 9 0 7 1 9 9 1 9 9 13 16 1 9 12 16 9 13 2
28 10 9 3 1 9 12 7 3 1 12 9 12 0 1 9 9 9 9 9 1 9 9 13 16 3 9 13 2
18 0 9 0 1 9 9 0 2 9 0 1 9 7 9 9 0 13 2
35 1 0 9 0 2 9 12 9 12 0 13 16 1 9 9 0 1 9 9 9 13 7 4 1 15 1 9 0 9 9 1 9 9 13 2
34 3 1 9 9 0 9 7 9 9 0 16 1 12 9 9 13 9 9 2 9 7 9 0 7 9 9 16 1 9 7 9 9 13 2
27 9 0 9 9 1 0 9 15 1 9 9 9 9 1 9 9 9 1 9 12 1 12 9 14 9 13 2
15 9 9 9 0 14 1 9 12 1 12 1 9 13 13 2
26 1 10 9 9 1 9 9 0 7 9 1 9 9 0 1 9 9 1 9 9 0 10 9 9 13 2
30 1 9 9 16 9 1 9 9 0 7 9 9 9 9 7 9 16 1 9 13 1 9 9 0 1 9 9 0 13 2
25 9 9 9 0 14 3 9 9 9 1 1 9 9 9 7 9 7 9 1 1 9 0 4 13 2
11 9 0 7 9 16 3 9 9 4 13 2
23 9 0 1 9 9 1 9 9 0 9 0 1 9 9 2 9 2 9 7 9 0 13 2
16 9 9 9 10 12 9 9 0 14 1 9 0 1 9 13 2
13 9 9 9 9 9 1 9 0 1 10 9 13 2
42 9 0 9 9 16 1 0 9 9 9 9 1 9 9 9 9 13 13 1 12 9 7 12 9 2 1 9 12 9 0 9 0 14 1 9 0 9 9 1 9 13 2
34 9 9 16 1 9 7 9 1 9 0 0 13 1 12 9 1 9 2 12 1 12 2 7 9 12 1 12 1 9 9 9 0 13 2
51 9 9 15 1 9 0 1 9 1 9 2 9 7 9 9 13 16 1 12 9 12 1 12 7 12 9 1 9 7 9 9 13 7 9 14 1 9 12 1 12 9 13 7 3 1 9 0 9 9 13 2
26 9 0 9 9 14 1 10 9 2 9 9 2 9 9 2 9 9 2 9 9 7 9 9 9 13 2
48 10 9 1 9 1 9 9 13 16 1 9 3 1 9 9 2 9 9 15 1 9 0 9 13 13 7 1 9 0 12 9 1 12 9 1 12 9 1 9 0 0 1 9 0 9 13 13 2
33 9 9 9 1 10 12 9 0 2 12 9 7 0 9 13 13 16 1 9 0 7 12 9 9 13 7 1 9 0 9 9 13 2
27 1 9 0 9 2 9 7 9 1 9 0 7 0 13 7 9 0 7 9 3 9 0 14 1 9 13 2
38 9 0 1 0 9 9 9 9 9 16 1 9 9 0 13 2 9 9 1 9 1 9 0 9 7 9 9 1 9 1 9 9 1 9 9 9 13 2
21 1 9 0 9 9 9 7 1 9 9 9 0 9 0 1 9 0 9 9 13 2
15 1 9 0 2 9 9 0 13 7 9 1 9 0 13 2
13 9 9 0 7 9 3 9 0 14 1 9 13 2
24 9 9 3 1 0 9 9 2 3 0 13 7 9 0 9 1 0 9 10 9 9 13 13 2
15 1 9 9 1 9 12 9 9 9 1 12 9 9 13 2
19 9 0 12 9 9 16 9 9 9 9 0 1 9 14 1 9 15 13 2
39 9 9 1 0 9 9 2 9 9 1 12 9 13 16 12 9 0 1 9 0 9 10 9 1 10 9 1 9 13 7 1 9 12 1 3 0 13 13 2
11 0 9 0 9 9 1 9 9 13 13 2
24 10 9 12 9 9 2 12 2 12 9 9 7 12 9 9 13 7 1 12 9 13 13 13 2
26 10 9 0 9 0 2 9 0 2 0 9 9 7 9 0 13 7 9 0 15 9 12 9 14 13 2
22 1 10 9 9 0 9 9 7 9 9 0 16 9 13 13 7 9 15 12 9 13 2
34 9 0 10 9 0 1 9 13 13 7 1 15 9 0 1 9 7 9 9 16 1 9 13 13 7 1 10 9 9 7 0 0 13 2
15 9 10 9 0 13 9 15 14 1 9 9 9 9 13 2
21 1 9 9 9 0 9 9 9 2 9 9 9 9 9 9 3 1 9 9 13 2
53 1 9 9 0 9 9 9 2 9 10 9 9 9 9 9 9 9 2 9 9 12 7 12 7 12 9 9 9 13 7 9 10 9 9 9 1 9 9 10 9 1 9 9 0 15 1 9 1 9 9 13 13 2
26 9 0 9 0 9 1 9 9 14 1 9 1 9 13 7 0 13 3 10 9 14 1 9 9 13 2
47 1 9 10 9 9 9 12 9 13 16 9 0 15 9 9 9 0 13 7 9 0 15 9 9 9 14 9 13 16 1 9 16 1 10 9 9 13 2 3 0 13 7 9 0 9 13 2
23 15 0 13 10 9 3 1 9 9 9 13 7 15 14 1 9 0 1 10 9 9 13 2
13 9 0 9 13 9 0 9 0 9 9 9 13 2
34 1 9 9 2 9 9 1 9 9 0 1 12 9 2 1 9 0 9 13 7 9 9 9 10 9 13 16 9 9 14 1 1 13 2
48 10 9 3 1 9 9 12 9 9 0 9 2 3 7 3 1 9 0 15 2 9 13 16 10 9 3 1 9 1 9 2 9 0 1 9 0 15 14 1 0 1 9 9 9 1 9 13 2
20 9 0 0 13 9 9 12 9 14 1 9 1 9 0 1 9 15 9 13 2
13 10 9 12 0 2 12 9 1 9 9 0 13 2
37 15 9 9 9 9 0 0 10 9 14 1 9 9 13 7 3 9 1 15 13 7 9 0 1 9 9 9 9 14 3 1 9 9 9 9 13 2
22 10 9 12 9 3 1 9 9 2 9 0 15 14 13 7 9 1 9 15 0 13 2
17 9 0 13 1 9 10 9 2 9 9 7 9 14 16 9 13 2
34 0 1 9 9 1 9 1 9 9 13 7 9 1 9 14 3 3 13 16 3 9 13 9 15 13 1 9 7 9 14 0 9 13 2
65 9 13 2 9 7 9 0 15 1 3 9 13 9 14 1 9 9 9 9 7 1 9 9 13 7 3 16 15 1 9 0 9 13 16 1 9 9 13 2 10 9 16 9 13 4 1 15 1 9 9 1 9 9 13 2 1 10 3 2 1 15 9 4 13 2
41 15 9 9 0 9 14 16 0 13 7 9 13 2 1 9 9 13 3 13 16 9 0 0 1 9 9 9 13 7 9 16 15 14 1 15 9 13 9 0 13 2
71 15 0 9 0 9 9 9 9 14 9 0 9 1 15 9 13 7 13 2 9 7 9 9 9 1 9 9 7 9 0 1 9 9 13 2 7 15 1 3 1 9 0 1 9 9 9 9 13 7 16 9 13 9 4 9 13 3 1 9 1 9 7 9 15 1 9 9 1 4 13 2
40 9 9 9 9 9 9 13 2 9 9 0 13 1 10 3 1 10 9 16 13 9 7 7 9 9 7 7 9 9 14 9 13 2 1 9 9 3 9 13 2
47 9 9 9 9 9 1 9 10 9 16 12 9 9 9 0 9 1 9 9 0 13 7 9 1 9 0 9 13 13 2 1 9 10 9 7 9 0 9 1 9 1 9 9 0 9 13 2
84 15 1 9 10 9 16 1 15 7 1 9 9 9 9 0 13 7 9 0 15 1 9 9 9 13 2 9 13 2 15 9 13 3 12 9 9 13 16 9 13 9 9 0 14 1 9 9 9 7 9 9 0 14 1 9 1 9 0 13 1 15 9 7 9 0 1 9 0 1 9 9 13 7 9 9 1 9 9 9 7 9 1 13 2
38 9 9 16 1 9 9 9 0 7 1 1 9 1 9 1 9 9 9 0 1 9 9 13 7 9 13 2 15 9 0 9 9 14 9 9 9 13 2
24 9 9 9 9 9 13 2 9 9 7 9 0 13 9 13 16 3 12 9 1 9 0 13 2
41 15 4 3 0 13 7 9 9 14 1 9 9 0 13 1 9 1 9 0 9 9 2 9 15 14 9 13 7 9 0 13 1 9 15 2 10 9 14 9 13 2
28 9 13 2 15 16 9 9 0 13 9 9 9 14 13 7 9 14 0 13 2 7 13 3 10 9 14 13 2
56 9 9 9 9 9 1 9 1 9 9 9 13 2 15 1 10 9 16 9 9 1 0 9 1 9 15 2 0 9 13 1 0 9 1 15 13 16 9 0 14 9 7 9 14 0 13 2 13 16 10 9 13 9 9 13 2
38 9 9 9 9 9 9 13 2 15 0 13 16 9 9 13 7 3 3 1 9 9 1 13 2 3 3 15 9 14 13 7 3 12 9 16 0 13 2
34 9 1 9 9 9 7 9 9 0 13 2 1 9 0 1 9 9 9 0 4 13 7 9 0 1 9 0 2 0 9 9 4 13 2
9 9 1 9 9 0 9 3 13 2
22 9 9 9 0 9 9 9 1 9 9 16 1 9 9 0 9 13 13 2 0 13 2
22 1 9 9 9 9 2 9 9 9 13 13 12 9 1 9 9 9 15 14 9 13 2
31 9 0 9 16 1 15 9 0 3 0 9 13 2 1 9 9 13 7 1 9 0 9 1 9 0 9 9 3 13 13 2
22 12 12 9 10 9 1 9 9 13 7 9 1 12 9 9 1 9 0 1 13 13 2
19 9 9 9 9 0 13 2 9 0 9 13 16 1 15 9 0 9 13 2
21 15 13 2 9 0 1 9 1 9 3 1 9 9 13 7 3 9 0 15 13 2
39 10 9 1 9 9 12 9 0 1 9 9 0 1 9 9 0 9 1 9 13 2 7 1 9 9 9 1 9 12 9 1 9 2 1 9 9 9 13 2
11 12 9 0 1 9 9 15 14 0 13 2
10 12 9 0 1 9 9 9 9 13 2
41 1 9 9 0 9 2 12 9 0 1 1 9 9 9 9 1 9 9 9 9 9 2 9 9 3 1 12 9 9 1 9 9 0 1 9 2 15 14 0 13 2
25 9 0 9 13 2 9 0 1 10 9 9 13 1 0 9 1 13 9 9 9 1 15 9 13 2
13 9 9 2 10 9 0 14 3 1 9 9 13 2
25 9 9 9 9 2 9 9 12 9 9 14 1 12 1 9 9 9 0 10 9 9 7 9 13 2
25 9 9 9 1 9 9 9 13 2 10 9 1 9 9 1 12 9 0 1 10 9 1 9 13 2
29 1 9 9 1 10 9 12 9 2 12 9 7 12 9 0 7 1 9 9 0 0 9 9 0 1 10 9 13 2
5 12 9 0 13 2
17 12 9 1 9 9 9 1 9 9 0 13 1 10 9 9 13 2
30 9 3 1 9 12 9 1 9 12 9 1 9 12 9 9 2 1 9 9 13 7 9 9 16 1 9 15 0 13 2
46 10 9 1 9 0 0 9 13 7 3 1 9 9 7 9 0 13 2 7 9 7 9 3 9 0 13 16 9 9 0 9 0 13 16 9 14 9 7 3 9 9 15 14 0 13 2
5 3 9 4 13 2
7 9 0 1 9 9 13 2
24 9 9 9 9 1 9 9 13 13 1 9 9 1 9 15 2 15 14 1 9 1 9 13 2
27 9 9 9 0 9 9 9 9 0 14 1 12 9 0 13 7 1 3 9 9 0 13 12 9 9 13 2
19 9 16 9 0 9 13 15 9 13 16 9 13 9 9 15 14 0 13 2
45 9 9 9 9 1 9 10 9 1 10 9 13 16 9 9 1 9 15 14 1 9 12 1 12 1 9 12 9 1 9 9 13 7 12 9 3 12 9 1 10 9 14 9 13 2
24 9 10 9 1 10 9 0 1 12 9 9 0 13 2 7 1 0 9 9 9 3 0 13 2
13 9 13 16 9 1 10 9 13 16 9 9 13 2
27 15 9 13 16 9 0 1 9 9 9 1 9 13 2 7 3 0 13 16 9 7 9 10 9 3 13 2
39 1 3 7 9 0 1 9 1 9 9 0 0 13 2 10 9 1 9 13 16 9 9 0 13 1 9 9 0 9 13 7 1 10 9 1 9 9 13 2
14 10 9 3 1 9 9 7 9 1 9 9 13 13 2
27 9 1 9 1 10 9 9 0 14 1 9 13 7 1 9 9 2 9 9 13 7 1 9 9 9 13 2
16 1 9 12 16 9 1 9 2 9 9 13 2 1 9 13 2
20 7 9 9 9 7 9 9 0 7 9 9 9 1 0 9 14 0 13 13 2
10 9 3 9 13 16 9 16 9 13 2
20 9 9 9 9 9 9 0 13 2 12 9 9 1 9 9 9 9 13 13 2
24 3 0 1 15 1 9 13 13 13 7 15 1 12 9 9 0 13 2 9 9 7 9 9 2
21 1 12 9 9 0 2 12 9 1 9 7 9 1 9 0 10 9 9 13 13 2
25 12 7 12 9 1 12 9 0 0 13 7 9 0 7 1 9 9 12 9 9 0 14 4 13 2
30 9 9 13 16 9 9 9 14 1 1 12 9 0 1 9 9 2 9 2 9 7 9 9 13 7 3 9 0 13 2
19 15 13 3 9 9 1 9 7 9 1 9 9 0 10 9 9 9 13 2
29 9 13 2 9 0 3 0 13 3 7 15 14 1 13 1 9 9 9 1 10 9 9 1 1 9 0 9 13 2
35 3 9 9 9 0 0 13 2 15 9 12 9 0 1 1 12 9 0 1 9 9 7 9 14 9 13 16 3 9 9 0 14 0 13 2
22 9 0 16 1 9 0 9 9 13 13 2 9 9 1 9 9 9 1 9 9 13 2
19 10 9 16 9 2 12 9 13 2 1 9 9 9 1 9 13 13 13 2
14 9 10 9 0 9 0 12 2 12 12 9 13 13 2
11 7 9 0 1 9 7 9 1 9 13 2
17 9 0 9 10 9 2 9 1 9 9 9 1 9 9 9 13 2
36 7 9 13 1 10 9 12 9 0 0 1 9 12 2 12 12 9 9 13 7 1 9 10 12 9 1 0 9 9 9 1 15 0 4 13 2
20 9 1 9 9 9 13 16 0 1 12 9 3 1 10 9 1 9 13 13 2
21 9 0 16 1 9 9 16 0 1 9 9 13 9 12 1 9 3 9 0 13 2
49 9 7 9 1 9 0 0 9 9 1 9 7 9 9 3 13 13 7 9 1 9 9 0 10 9 9 16 1 9 0 9 1 9 0 3 1 9 2 12 9 0 9 13 2 0 7 0 13 2
33 1 9 9 0 9 2 9 9 9 9 13 9 0 14 16 12 9 0 1 9 9 1 9 1 9 9 13 13 13 14 1 13 2
35 12 1 9 16 1 9 0 13 9 9 1 10 9 13 16 1 9 12 1 9 9 9 1 9 9 1 9 9 9 7 1 9 0 13 2
38 1 0 9 9 2 9 9 9 13 16 1 9 9 0 1 9 9 1 3 9 16 1 9 12 1 12 1 9 0 1 9 9 9 1 9 0 13 2
40 10 9 16 1 9 0 7 0 9 9 16 1 9 15 9 13 13 1 9 0 16 1 9 9 7 1 9 9 0 9 9 9 9 13 13 13 2 9 13 2
50 9 0 9 0 13 16 9 1 9 9 1 9 7 9 0 13 16 3 1 9 9 9 0 13 7 12 1 9 16 9 9 1 3 13 13 10 13 16 1 9 9 1 9 9 1 9 1 9 13 2
16 1 9 9 0 1 9 12 9 1 9 12 9 0 13 13 2
39 0 9 9 3 1 15 7 9 9 14 1 9 1 9 0 9 13 2 12 9 0 1 9 7 9 9 9 7 9 9 16 9 15 1 9 13 0 13 2
28 16 10 9 1 9 9 9 9 0 7 0 13 2 2 7 1 9 9 9 9 1 9 0 9 15 0 13 2
36 9 1 9 9 9 15 14 3 9 0 9 13 7 9 13 16 1 9 0 1 9 9 13 2 16 15 1 9 16 3 1 9 13 0 13 2
25 9 0 9 15 13 16 9 9 13 9 14 1 9 9 9 13 16 9 1 9 9 0 9 13 2
21 1 10 9 1 10 9 9 0 4 13 16 9 0 14 1 9 9 0 9 13 2
38 9 9 7 9 9 9 0 9 7 9 2 16 9 14 3 3 9 16 1 1 9 0 13 2 1 1 9 15 0 13 2 1 9 9 9 0 13 2
84 7 10 9 16 9 15 9 0 14 1 9 1 13 7 16 9 16 1 9 1 9 0 13 13 9 15 14 1 9 9 13 2 7 1 9 0 7 9 0 9 9 0 13 2 9 1 9 9 9 7 9 9 2 1 1 15 9 9 1 10 9 0 13 2 9 1 9 0 9 13 7 0 1 9 0 1 9 9 13 7 3 9 13 2
41 3 9 0 0 7 0 2 1 9 9 13 7 10 9 16 1 9 0 2 7 0 2 7 0 2 7 9 0 13 9 9 13 7 3 9 1 9 10 9 13 2
44 16 7 9 9 14 1 9 1 9 9 13 2 9 9 0 9 9 13 16 15 14 9 0 13 7 0 13 2 16 3 1 15 9 9 0 9 15 14 3 1 9 13 13 2
30 9 1 9 9 15 1 9 13 7 16 9 0 9 7 9 15 14 1 9 10 9 13 2 9 13 16 9 14 13 2
7 9 9 0 9 0 13 2
28 9 1 15 13 16 9 15 15 2 3 1 15 16 0 9 9 15 1 9 13 2 1 3 9 1 4 13 2
9 16 7 1 9 0 9 15 13 2
24 1 9 9 15 1 9 9 1 9 13 16 1 3 9 9 1 9 0 1 9 0 13 13 2
37 9 0 14 16 1 9 9 9 13 1 1 9 0 16 1 9 13 7 1 1 9 0 13 13 13 2 7 9 1 15 13 7 1 9 9 13 2
6 9 9 0 9 13 2
39 1 9 7 9 0 9 0 9 9 0 14 1 9 0 9 7 9 9 9 14 1 15 9 13 13 2 0 1 9 7 3 9 1 10 9 0 0 13 2
24 9 9 0 1 12 1 12 9 9 9 13 7 0 9 0 9 9 7 9 1 9 9 13 2
26 1 9 0 16 9 9 9 9 13 2 1 9 9 7 9 1 1 9 0 9 9 12 0 9 13 2
32 9 9 2 10 9 14 12 9 7 9 9 12 9 9 13 2 1 9 7 9 0 0 9 9 1 9 0 2 12 9 13 2
12 10 9 1 1 9 9 9 16 9 0 13 2
26 9 9 9 12 1 9 10 9 13 2 9 0 9 9 0 1 1 9 0 2 9 0 7 0 13 2
38 9 7 9 4 1 9 0 1 1 9 9 9 0 9 13 7 13 16 9 1 9 0 2 3 3 0 1 10 9 13 16 1 12 9 3 9 13 2
11 9 0 1 9 9 9 2 10 9 13 2
22 9 16 1 9 0 1 9 9 9 9 9 1 9 9 9 9 13 2 10 9 13 2
36 9 9 9 9 1 9 9 0 9 1 9 13 2 12 9 9 0 1 9 9 2 2 3 1 9 1 9 9 9 0 9 0 9 0 13 2
33 9 9 1 12 9 0 9 9 16 1 15 9 9 9 9 13 2 0 1 15 13 16 9 15 3 1 9 2 10 9 0 13 2
26 1 9 1 9 9 0 2 9 0 1 9 1 9 1 9 0 1 9 9 1 9 0 0 9 13 2
24 9 9 9 9 9 0 0 13 16 1 9 15 9 9 0 1 9 9 9 9 0 9 13 2
22 1 0 9 9 1 9 9 2 9 9 9 0 0 14 1 9 10 9 9 9 13 2
22 9 9 9 9 9 9 13 2 9 0 14 1 9 9 9 9 1 9 9 13 13 2
38 9 0 16 9 0 15 1 9 9 0 9 13 2 9 0 9 10 9 0 1 9 4 13 7 9 0 1 9 7 9 0 1 9 14 9 4 13 2
39 9 9 9 0 9 1 9 10 9 13 2 9 10 9 9 1 9 9 9 1 9 9 9 13 1 15 7 9 1 9 9 0 1 9 9 7 9 13 2
26 9 0 9 1 9 13 10 9 9 1 1 9 0 1 9 13 2 15 14 3 1 9 1 9 13 2
32 9 0 9 0 9 1 9 9 9 0 9 10 9 13 16 9 0 0 1 9 14 1 9 9 0 1 1 9 0 9 13 2
24 9 9 9 1 9 9 0 9 9 9 16 9 1 9 0 10 9 1 10 9 14 9 13 2
17 9 9 9 1 9 9 15 14 1 12 9 12 12 0 9 13 2
26 1 10 9 12 9 9 9 7 12 9 9 9 9 9 0 16 0 1 9 9 9 13 2 9 13 2
33 9 9 0 7 9 16 1 12 1 9 9 9 9 13 13 2 9 9 1 9 9 9 1 9 12 2 12 12 9 1 9 13 2
48 1 9 9 9 2 1 10 9 9 16 0 9 9 0 13 7 1 1 15 9 1 9 9 9 2 9 9 1 9 12 9 0 9 13 2 12 1 12 12 9 9 9 1 9 13 13 13 2
32 10 9 9 16 1 9 9 0 1 12 1 0 7 0 9 9 9 1 9 13 2 1 9 0 1 9 1 9 13 13 13 2
40 9 0 1 9 9 0 9 0 2 9 9 0 13 7 1 9 9 9 9 9 2 9 0 1 9 0 9 7 9 9 0 2 9 9 7 9 9 0 13 2
28 9 9 16 1 9 13 9 0 1 9 9 9 1 9 0 9 13 2 9 9 9 2 9 7 9 9 13 2
54 1 9 15 7 0 1 9 9 9 0 7 9 9 0 14 9 0 13 2 7 9 13 9 0 1 9 0 1 1 9 9 13 7 1 9 16 9 9 15 14 1 9 13 13 2 4 9 9 9 0 14 9 13 2
52 1 9 9 10 9 16 1 10 9 0 1 9 9 0 1 9 9 13 13 2 0 9 9 0 13 16 1 9 1 9 9 7 9 9 13 7 3 1 9 9 9 9 1 9 0 7 9 1 15 9 13 2
30 9 9 0 9 9 13 2 0 9 9 0 1 10 9 1 9 9 2 9 1 9 12 2 12 9 9 9 13 13 2
15 10 9 9 2 0 9 9 9 0 9 0 1 9 13 2
61 9 9 9 9 2 9 9 1 9 1 10 9 13 2 1 9 0 9 9 2 9 9 1 9 9 12 9 9 13 1 9 16 0 9 9 1 9 12 1 9 9 0 9 1 9 12 2 12 2 12 9 0 1 9 0 1 9 0 0 13 2
24 9 9 9 3 1 9 9 0 9 9 13 2 7 1 9 9 9 10 9 16 9 13 13 2
16 1 15 7 9 9 9 9 9 9 0 1 10 9 13 13 2
13 9 9 7 9 1 9 9 1 9 9 9 13 2
38 9 9 9 9 9 9 9 9 1 9 13 2 1 9 7 0 1 9 1 9 0 9 9 13 2 7 1 9 9 7 9 1 9 9 9 0 13 2
33 1 9 9 2 12 0 1 9 9 1 9 9 9 2 12 0 1 9 9 0 7 9 7 12 0 0 1 9 9 0 9 13 2
24 1 9 9 0 1 9 9 9 0 2 9 7 9 1 9 9 0 0 7 9 0 9 13 2
23 1 9 9 0 2 9 12 9 1 9 9 9 0 1 9 1 9 0 0 0 9 13 2
19 1 9 0 3 4 1 9 9 12 0 1 9 1 9 9 9 9 13 2
42 9 9 1 9 9 9 0 0 1 9 1 9 1 9 9 13 16 1 9 10 9 9 1 9 0 9 13 7 1 9 1 9 2 9 9 1 9 0 9 13 13 2
17 9 9 7 9 1 9 9 16 1 9 9 9 0 9 13 13 2
24 9 9 9 1 12 12 9 1 9 9 7 9 0 9 9 9 1 9 0 0 9 4 13 2
37 1 9 9 9 1 9 2 9 9 9 7 9 9 9 9 2 1 9 0 9 9 14 1 9 7 9 9 1 9 12 2 12 12 9 9 13 2
16 1 10 9 3 12 9 9 0 1 9 0 0 9 4 13 2
20 9 1 10 9 1 9 9 15 1 9 9 9 1 9 1 9 0 4 13 2
37 9 9 9 13 2 10 9 13 1 15 9 0 1 9 9 9 2 9 0 2 9 0 7 0 2 9 7 3 9 9 7 9 9 0 9 13 2
21 1 10 9 2 9 0 0 3 9 2 9 7 9 0 1 9 7 9 0 13 2
20 9 13 2 9 9 13 1 9 1 9 0 1 9 15 1 9 0 9 13 2
7 0 9 9 9 9 13 2
21 9 0 9 9 9 16 0 9 9 13 2 13 16 1 9 0 9 9 9 13 2
20 9 9 9 12 0 2 3 1 9 9 0 1 9 9 9 9 1 9 13 2
21 15 13 16 0 1 9 9 13 1 9 9 13 7 3 9 9 1 9 13 13 2
30 9 1 9 12 2 16 0 9 3 1 9 0 0 2 0 9 13 7 1 10 3 2 12 9 0 9 9 13 13 2
26 15 16 12 9 16 9 9 13 13 2 12 9 3 1 9 12 9 9 9 9 9 14 1 9 13 2
35 1 10 9 4 1 9 9 9 9 9 1 9 2 9 1 9 1 9 2 9 0 1 12 9 7 9 7 9 1 9 12 9 9 13 2
19 1 9 13 16 9 0 12 1 0 9 9 9 9 9 1 9 0 13 2
49 16 9 0 9 1 9 9 1 9 0 3 3 0 13 2 7 1 9 3 0 10 9 16 9 9 9 9 7 3 9 1 9 0 13 2 9 9 7 9 9 14 16 1 10 9 1 9 13 2
22 3 0 13 13 16 3 9 1 9 9 16 9 0 1 0 9 9 9 9 0 13 2
8 0 13 16 0 9 9 13 2
10 16 10 9 7 9 14 3 9 13 2
6 16 0 9 0 13 2
4 3 0 13 2
13 9 15 1 9 9 0 0 1 10 9 0 13 2
17 9 9 9 9 7 9 9 0 1 9 0 9 7 9 0 13 2
32 16 1 9 1 9 9 13 3 9 12 9 1 9 9 13 16 16 3 1 9 0 9 9 13 3 1 1 9 15 9 13 2
2 9 2
11 16 1 15 0 13 2 9 9 15 13 2
17 15 9 9 14 1 9 15 0 13 2 3 9 1 15 9 13 2
14 9 9 9 13 2 3 15 7 9 9 1 15 13 2
14 15 15 4 9 1 9 14 13 7 9 14 9 13 2
14 16 1 0 9 1 9 9 13 2 3 9 9 13 2
12 0 9 9 9 2 9 9 0 1 9 13 2
8 9 2 0 9 9 9 13 2
14 15 9 13 16 0 9 12 9 3 0 2 9 13 2
17 1 9 9 2 9 1 9 13 7 9 0 1 9 0 9 13 2
20 1 10 9 1 9 9 9 0 13 7 3 9 0 7 0 1 9 9 13 2
25 9 9 9 1 9 9 2 10 9 9 9 13 7 0 1 9 9 0 0 1 9 9 9 13 2
46 1 9 4 1 1 10 9 2 1 9 0 0 1 9 7 9 9 13 7 3 9 1 9 0 1 9 9 7 7 9 1 9 0 1 9 9 9 13 16 0 9 0 1 9 13 2
25 1 9 9 2 9 0 4 1 9 9 1 9 9 16 9 9 9 3 0 9 13 2 9 13 2
13 1 9 9 0 2 9 9 1 9 0 9 13 2
32 9 9 13 16 9 0 9 14 1 9 0 7 0 9 13 7 9 7 9 9 14 1 9 9 13 16 9 3 9 0 13 2
18 1 9 9 16 9 1 9 7 9 15 1 9 0 2 0 7 0 2
32 1 9 0 9 9 9 9 14 9 13 16 9 0 1 9 15 9 0 14 13 2 9 2 9 7 9 7 1 15 9 13 2
40 9 16 9 9 13 0 9 0 13 16 1 9 0 1 9 9 13 7 9 0 15 1 9 9 1 9 9 2 9 7 9 9 9 7 9 9 9 9 13 2
29 9 1 9 16 1 15 9 1 9 9 0 2 9 0 1 9 7 9 9 9 9 0 0 9 13 2 9 13 2
31 16 10 9 7 9 3 9 9 7 9 9 0 13 2 9 16 1 9 9 9 13 2 16 9 1 9 0 1 9 13 2
14 9 1 9 1 0 9 9 10 9 14 4 9 13 2
22 9 7 9 0 15 14 1 9 0 9 13 7 1 9 0 1 9 0 15 9 13 2
13 1 10 9 16 13 1 9 0 7 0 9 13 2
28 1 9 9 9 0 15 7 9 15 14 0 1 9 0 9 13 7 1 9 0 9 13 2 3 9 7 9 2
8 3 7 1 9 0 9 13 2
7 1 9 0 9 9 13 2
11 1 9 9 0 9 1 9 9 9 13 2
11 9 0 9 2 1 9 9 0 9 13 2
15 1 9 9 16 0 9 0 9 7 9 13 2 9 13 2
14 9 15 14 0 9 13 7 15 14 1 9 0 13 2
14 1 9 9 0 1 12 9 9 13 7 9 0 13 2
17 10 9 9 1 9 0 7 9 15 14 1 9 0 9 9 13 2
9 9 0 14 1 9 0 9 13 2
25 9 0 12 9 13 16 9 13 1 2 9 2 9 2 9 2 9 0 7 9 2 9 7 9 2
41 9 0 1 9 9 0 9 1 9 0 13 1 2 2 9 9 2 9 2 9 2 1 9 9 9 9 1 9 1 9 10 9 9 9 1 9 0 1 9 13 2
16 1 9 9 9 9 0 2 0 1 9 1 9 9 0 13 2
27 9 9 2 9 2 9 2 9 9 1 9 9 2 9 0 9 2 9 0 1 1 9 0 9 9 13 2
19 9 1 9 9 2 9 0 1 9 0 0 1 9 1 9 0 9 13 2
34 9 9 7 9 0 2 0 2 0 2 1 9 9 9 16 9 0 9 13 1 9 0 1 9 1 9 16 9 0 13 2 9 13 2
13 16 1 9 1 9 0 9 0 10 9 9 13 2
25 9 9 0 0 13 16 1 9 0 9 7 9 9 2 3 9 1 9 0 3 9 14 9 13 2
19 9 9 9 9 9 3 0 13 7 16 4 10 9 1 9 9 9 13 2
12 9 0 9 1 12 9 0 7 0 9 13 2
13 9 0 0 9 9 2 9 2 9 7 9 13 2
60 7 13 9 1 9 9 2 9 2 9 2 9 7 9 9 2 9 0 2 9 2 9 2 9 2 9 0 2 9 2 9 2 9 2 9 2 9 9 2 9 2 9 2 9 0 2 9 9 7 3 15 14 9 9 0 9 1 9 13 2
6 9 9 0 0 13 2
12 9 0 9 0 9 13 16 0 9 0 13 2
31 9 9 3 9 1 9 1 9 1 9 0 1 9 9 13 2 7 4 1 12 1 12 9 9 0 1 9 9 9 13 2
18 16 1 9 9 0 9 10 9 1 9 0 9 1 9 9 9 13 2
37 9 0 9 2 9 0 13 16 3 7 1 15 9 0 13 7 1 9 7 9 0 1 9 9 2 9 9 7 9 9 1 15 0 9 0 13 2
12 10 9 7 9 7 9 13 9 14 9 13 2
24 9 16 0 13 9 0 0 13 13 16 3 9 14 1 9 0 9 9 15 2 0 9 13 2
37 1 10 9 9 16 0 13 3 9 9 0 7 0 3 9 2 9 2 9 7 9 2 9 0 7 0 1 9 13 7 9 0 9 14 0 13 2
12 10 9 0 13 9 14 1 9 0 0 13 2
12 9 0 7 9 0 2 1 9 10 9 13 2
23 3 9 0 10 9 1 9 0 13 15 14 0 9 2 9 2 0 9 7 3 9 13 2
21 7 9 15 13 0 1 9 2 9 13 7 1 9 2 9 7 0 9 9 13 2
21 9 0 0 13 2 9 0 13 13 7 1 10 9 10 9 0 9 14 0 13 2
41 1 9 0 0 2 12 9 0 1 9 0 9 2 10 9 14 1 13 7 0 1 12 9 9 9 14 0 13 7 9 0 2 0 7 0 9 9 0 14 13 2
27 1 1 9 2 9 0 2 9 14 1 15 1 9 7 9 13 16 9 0 10 9 1 1 15 9 13 2
25 3 7 9 9 1 9 12 1 9 9 9 9 16 1 12 9 9 9 13 13 2 1 1 13 2
30 9 0 0 2 9 1 9 7 9 0 14 1 9 9 13 7 1 9 9 0 15 14 0 13 7 1 1 13 13 2
39 3 2 16 9 16 1 9 9 9 13 2 3 7 9 9 0 2 9 14 9 13 7 10 9 1 9 13 16 9 0 7 0 16 1 10 9 0 13 2
27 1 9 9 2 10 9 7 9 1 9 9 13 1 10 9 9 0 2 9 9 9 14 1 9 9 13 2
25 9 0 7 0 10 12 16 9 7 9 1 1 15 1 9 9 13 16 9 1 9 15 9 13 2
16 1 9 9 2 9 0 9 3 9 14 1 1 9 4 13 2
23 10 9 9 14 0 9 9 2 9 7 9 13 7 9 7 9 9 14 1 9 9 13 2
21 9 0 9 1 1 9 1 10 9 0 2 9 0 2 9 7 9 0 9 13 2
26 9 1 1 9 0 13 2 16 3 9 9 1 9 15 13 16 12 9 7 12 9 14 0 9 13 2
14 1 9 7 9 7 9 0 1 1 10 9 0 13 2
21 3 16 9 0 1 9 0 0 13 2 3 9 9 13 16 9 9 14 9 13 2
32 7 10 9 1 9 0 1 9 0 7 0 9 13 7 7 1 9 9 9 9 0 9 9 13 16 1 15 9 7 9 13 2
28 9 2 0 9 0 13 16 9 0 1 1 9 1 9 0 7 1 1 9 0 1 9 1 9 0 9 13 2
15 16 9 1 9 9 0 1 9 2 0 9 7 9 13 2
55 1 9 9 2 0 9 3 12 1 9 16 1 9 0 1 9 9 0 9 9 13 2 0 1 9 9 0 0 1 9 9 13 13 7 10 9 9 9 9 0 14 13 13 16 3 10 9 3 1 9 10 9 9 13 2
16 9 15 13 16 3 9 0 1 1 9 9 10 15 0 13 2
17 3 1 9 0 1 13 16 9 15 2 9 9 9 9 9 13 2
15 9 10 9 1 9 9 1 9 9 2 9 15 14 13 2
46 15 3 9 9 9 7 9 9 9 9 7 9 15 1 9 12 9 0 9 13 16 1 9 10 9 7 1 9 0 2 9 7 1 9 9 9 1 10 9 1 1 13 7 0 13 2
15 1 0 9 9 3 9 13 13 16 9 0 1 9 13 2
73 16 15 9 9 9 14 1 9 1 9 13 13 2 9 10 9 4 13 16 3 9 13 2 9 9 9 0 14 9 13 4 2 3 0 1 9 9 9 7 0 15 13 2 7 4 1 1 9 9 0 1 9 9 2 9 2 9 2 9 9 2 9 2 9 7 9 0 10 9 16 0 13 2
24 9 9 0 7 0 2 15 1 9 9 9 9 7 7 9 16 1 1 15 13 2 9 13 2
41 1 9 1 9 0 2 12 9 0 0 13 12 9 14 9 9 7 9 9 13 7 9 0 15 14 0 1 0 9 9 7 9 0 0 1 12 9 0 9 13 2
14 0 13 16 10 9 9 0 0 14 1 9 4 13 2
20 3 9 1 10 9 16 16 15 3 0 13 7 6 2 1 9 9 9 13 2
49 1 9 2 9 9 0 1 9 3 1 9 12 9 9 13 2 16 1 10 9 16 9 9 7 9 1 9 0 7 0 9 13 2 9 0 1 10 9 15 14 9 13 7 1 9 9 16 13 2
37 7 0 1 9 0 16 1 9 9 13 7 16 15 7 12 9 0 13 7 9 7 9 1 15 9 13 7 9 1 1 9 15 9 10 9 13 2
23 3 9 16 9 15 14 9 13 2 9 15 1 9 1 9 9 0 7 0 15 9 13 2
27 9 9 9 1 9 15 1 10 9 13 13 16 9 9 0 0 1 9 2 9 0 1 1 9 9 13 2
44 16 9 1 9 2 1 9 9 7 0 13 7 3 1 10 9 1 1 9 9 13 1 9 7 9 1 9 1 9 9 13 7 1 9 15 13 16 9 0 1 9 15 13 2
13 10 12 9 3 9 15 14 1 10 9 9 13 2
19 1 9 0 9 0 0 9 15 14 9 13 7 1 9 9 9 9 13 2
23 1 1 9 7 9 0 2 15 1 9 1 9 9 15 1 9 0 7 9 0 9 13 2
16 10 9 9 14 1 9 13 7 15 14 9 9 1 9 13 2
19 16 1 9 1 9 1 10 9 16 9 4 9 14 9 13 2 9 13 2
24 16 2 9 7 9 1 9 9 7 9 9 7 9 9 9 1 1 10 9 9 3 0 13 2
45 9 9 1 9 9 1 9 0 9 13 2 3 1 15 7 9 9 1 9 9 13 7 9 9 9 14 9 13 2 9 14 1 9 9 1 9 13 16 4 1 9 7 9 13 2
11 9 1 9 9 9 9 7 9 9 13 2
21 1 10 9 0 9 7 9 9 9 7 9 0 14 9 13 7 1 9 9 13 2
34 9 0 7 10 9 9 1 10 9 1 9 9 7 9 9 13 7 3 1 9 9 7 9 12 9 1 9 13 16 3 1 9 13 2
40 9 1 9 9 7 9 9 9 1 9 7 9 9 14 9 13 16 1 9 0 9 7 9 9 13 7 9 7 9 1 9 9 9 9 15 9 14 9 13 2
15 3 1 9 9 4 9 9 0 7 9 1 9 9 13 2
34 1 10 9 9 1 9 9 9 1 9 9 9 13 7 9 1 9 9 9 15 14 9 13 7 1 15 1 9 9 9 15 9 13 2
45 10 9 1 10 9 12 9 0 13 7 10 9 7 9 9 1 12 9 0 0 3 1 15 9 13 13 2 1 1 16 4 10 9 14 9 13 16 9 9 9 14 1 9 13 2
20 3 1 10 9 2 9 9 3 9 13 7 9 10 9 14 1 9 9 13 2
11 10 9 0 4 1 9 1 9 9 13 2
31 1 9 10 9 9 14 1 9 9 13 7 9 9 7 9 0 15 14 9 13 7 9 1 9 7 9 1 9 15 13 2
11 9 1 9 9 1 9 7 9 0 13 2
29 1 9 9 9 2 15 4 9 14 1 9 9 13 7 15 14 9 13 1 9 9 9 15 14 13 7 9 13 2
15 9 9 14 1 9 9 9 1 9 0 9 3 9 13 2
23 3 1 15 1 9 13 16 1 1 9 9 9 1 9 9 1 9 13 7 3 9 13 2
25 3 9 9 9 3 9 12 1 9 0 9 13 16 1 9 0 3 13 9 9 9 7 9 13 2
33 1 9 12 9 0 13 13 7 9 9 9 16 3 1 9 9 13 13 3 13 7 7 15 7 9 9 0 1 9 9 9 13 2
43 3 9 9 9 1 9 9 9 9 14 12 9 9 13 7 9 16 0 13 16 10 3 9 9 9 1 9 9 0 1 9 9 9 13 16 1 10 9 9 9 13 13 2
20 10 9 1 9 9 7 9 9 9 13 7 3 1 12 9 0 9 9 13 2
29 1 9 0 10 9 2 9 3 9 0 2 9 9 2 9 2 9 0 2 9 9 7 9 7 9 1 9 13 2
27 9 1 9 9 1 9 9 1 10 9 0 13 16 16 9 0 13 16 1 12 1 12 9 9 13 13 2
20 16 0 13 9 3 9 13 13 7 3 9 12 9 9 0 9 9 15 13 2
29 16 1 9 9 13 1 9 9 9 1 9 1 9 1 9 9 13 16 1 9 9 10 9 9 3 0 9 13 2
8 3 9 1 9 9 9 13 2
33 9 9 9 3 9 14 16 9 0 9 14 1 9 13 7 3 9 1 9 0 1 12 9 7 7 0 1 12 9 14 0 13 2
34 9 9 13 9 16 9 0 13 7 7 1 9 9 9 0 9 0 2 9 0 13 2 1 9 9 0 1 9 1 9 9 9 13 2
21 7 13 13 16 9 0 9 0 3 9 7 9 0 1 9 9 9 14 9 13 2
15 9 1 9 2 9 9 7 9 9 16 1 9 9 13 2
8 9 1 9 9 3 4 13 2
17 10 9 4 1 9 9 1 9 1 9 9 13 1 9 9 13 2
19 9 9 1 9 0 9 0 12 9 7 1 12 9 12 9 12 9 13 2
11 1 10 9 9 9 9 7 9 9 13 2
31 7 9 0 1 9 0 3 9 9 1 9 9 9 2 9 9 2 0 9 9 7 9 9 7 0 9 9 9 9 13 2
15 9 0 1 1 9 0 9 1 9 1 9 9 9 13 2
21 1 10 9 9 13 9 1 9 13 13 7 1 9 9 2 9 9 14 0 13 2
11 9 9 10 9 1 9 9 0 9 13 2
30 1 9 0 9 16 9 9 7 9 0 9 16 9 3 9 13 7 7 9 9 9 7 9 9 13 2 9 9 13 2
25 9 9 13 7 9 9 9 9 13 7 1 9 0 9 9 1 9 9 9 9 9 7 9 13 2
35 7 0 9 0 13 7 7 9 9 9 14 0 13 7 3 9 0 13 7 16 9 16 13 9 13 2 9 9 9 9 15 14 0 13 2
8 9 16 12 9 9 9 13 2
19 9 9 9 14 0 13 7 1 9 9 16 9 0 13 2 1 9 13 2
13 9 9 14 0 13 7 9 9 9 1 9 13 2
11 7 1 9 9 0 7 9 9 0 13 2
12 9 9 1 9 9 1 9 9 3 3 13 2
40 9 0 9 13 16 9 9 0 2 9 9 7 9 9 13 7 1 9 9 7 9 9 9 13 7 1 9 1 9 2 9 2 9 2 9 7 2 9 13 2
19 1 9 9 0 2 9 2 9 0 7 0 2 9 9 7 2 0 13 2
9 9 0 13 7 0 9 9 13 2
7 7 9 9 9 0 13 2
7 9 1 9 9 9 13 2
8 9 9 1 9 9 13 13 2
7 1 9 1 3 13 13 2
14 9 9 1 9 9 9 9 9 9 9 14 13 13 2
12 9 0 9 9 9 1 9 0 9 13 13 2
13 9 9 9 9 9 14 1 9 9 9 13 13 2
15 10 9 16 9 9 1 9 9 1 9 0 9 13 13 2
14 0 1 9 7 9 1 15 9 1 9 0 13 13 2
16 15 0 9 13 7 0 9 1 9 9 1 9 0 13 13 2
13 9 15 1 9 0 9 0 1 9 9 13 13 2
15 0 9 0 15 1 1 9 9 1 9 0 9 13 13 2
13 9 1 9 9 9 1 9 1 9 10 9 13 2
15 16 9 9 15 14 1 9 9 1 9 0 9 13 13 2
13 3 1 9 0 9 10 9 0 1 9 13 13 2
6 9 9 9 9 13 2
40 9 9 9 9 9 2 9 2 9 7 9 0 9 9 9 9 2 3 1 9 0 7 0 1 9 9 9 2 9 9 2 1 9 0 9 1 9 9 13 2
18 9 9 9 1 9 12 1 9 0 7 0 1 9 9 1 9 13 2
30 9 15 9 9 9 9 9 9 9 9 2 1 9 0 7 1 9 9 7 9 9 7 9 15 9 9 7 9 13 2
25 7 16 1 9 9 9 9 9 9 2 9 9 0 9 9 13 7 1 9 9 0 15 9 13 2
68 9 1 9 9 9 0 7 0 1 15 9 13 1 1 9 1 9 0 0 7 0 9 0 13 7 1 9 1 9 0 2 1 9 9 0 16 9 13 1 3 7 15 16 1 9 12 1 9 0 7 0 2 16 1 9 9 7 9 7 16 1 9 9 7 9 9 13 2
43 15 1 1 9 7 9 0 1 9 7 9 0 1 9 9 9 2 0 9 9 1 9 0 9 13 7 1 9 7 9 7 9 0 7 0 1 9 9 9 0 9 13 2
28 9 9 0 15 1 9 9 9 0 0 2 12 9 9 1 9 7 9 7 9 9 7 9 9 0 13 13 2
64 9 9 9 2 1 3 7 10 9 9 7 9 1 9 9 0 14 0 1 9 7 9 9 9 13 7 13 1 10 0 9 9 9 12 1 9 9 0 7 0 2 9 1 9 13 7 1 9 0 0 7 0 2 15 16 1 9 0 9 9 1 9 13 2
47 9 12 9 9 0 15 9 0 1 12 9 9 13 16 3 1 9 9 7 9 0 1 9 9 9 9 3 9 9 2 9 9 9 2 9 9 9 2 9 9 9 9 9 7 2 13 2
31 7 9 12 9 1 9 7 9 3 9 9 2 9 9 7 9 9 7 9 0 1 15 9 0 7 0 14 1 9 13 2
26 3 15 9 1 9 9 9 0 9 9 9 0 7 0 9 9 0 9 9 0 15 9 9 13 13 2
57 9 9 0 9 10 9 0 14 1 9 9 9 7 9 2 1 0 9 0 9 7 9 9 9 7 9 0 15 9 9 9 9 9 9 9 9 13 2 1 10 9 1 9 9 0 2 9 9 7 1 9 9 7 9 9 13 2
31 9 9 0 9 9 2 1 9 9 0 15 1 10 9 2 1 9 1 9 1 12 9 0 0 2 1 9 15 9 13 2
62 9 10 9 16 1 9 9 9 0 0 9 13 1 10 9 13 2 9 9 2 9 9 2 9 9 2 9 9 2 9 9 2 9 9 2 9 9 2 9 9 9 2 9 9 9 2 9 9 2 9 9 9 2 9 9 2 9 9 7 9 9 2
25 1 10 9 9 9 1 9 9 0 1 9 9 9 9 1 9 1 13 7 3 1 9 9 13 2
9 9 12 9 0 2 0 9 13 2
17 10 9 2 0 9 1 9 9 9 13 16 1 9 9 9 13 2
19 0 9 9 1 9 9 9 13 16 1 9 9 9 1 9 12 9 13 2
15 10 9 0 1 9 1 9 0 9 1 9 0 0 13 2
12 0 9 2 1 9 1 9 9 9 9 13 2
28 9 9 9 9 3 1 9 9 0 9 9 9 13 2 1 9 0 12 12 9 0 1 9 1 9 9 13 2
50 9 16 1 9 9 1 9 15 9 13 13 2 1 9 1 10 9 1 12 12 9 9 9 13 1 9 7 9 0 1 9 9 12 12 7 12 9 0 2 1 12 12 9 1 9 9 9 13 13 2
17 15 9 9 1 10 9 14 12 12 7 12 9 9 1 9 13 2
25 9 9 16 13 2 1 9 9 0 9 12 12 7 12 9 0 1 12 12 9 9 1 9 13 2
32 1 9 15 2 1 9 9 9 0 1 9 10 9 1 12 12 9 9 9 13 16 1 1 9 9 0 12 9 9 13 13 2
26 9 9 13 2 16 1 9 10 9 7 1 9 9 0 1 12 12 9 1 9 0 9 9 13 13 2
41 9 9 1 9 0 0 9 9 9 13 7 13 2 1 9 9 0 12 9 9 1 10 9 9 13 16 1 9 9 0 12 9 7 12 12 9 15 9 13 13 2
22 9 9 13 2 16 12 12 9 1 9 9 1 9 9 0 7 9 9 9 13 13 2
42 9 9 9 9 0 9 0 1 9 0 1 9 10 9 14 1 9 12 9 9 9 13 7 13 2 16 1 10 9 12 12 9 9 0 16 1 9 9 0 0 13 2
16 9 9 9 9 0 1 9 9 0 14 12 9 9 9 13 2
28 15 16 9 13 16 1 9 0 12 12 9 1 9 9 9 7 9 0 7 9 0 0 1 9 9 9 13 2
58 9 9 1 9 15 16 9 9 1 9 9 0 1 9 0 1 9 15 9 13 13 2 15 1 9 0 1 9 9 13 3 9 0 13 0 1 9 12 13 7 1 9 0 9 9 1 9 0 1 9 9 7 9 1 9 13 13 2
35 15 1 9 9 9 1 9 12 9 7 13 2 1 9 12 3 9 1 9 9 7 9 9 9 13 7 10 9 9 13 9 9 4 13 2
9 9 9 12 12 9 9 9 13 2
23 9 9 0 9 9 13 9 0 9 1 9 9 1 9 9 1 0 1 12 12 9 13 2
30 1 9 9 10 9 1 9 1 9 9 2 9 1 12 9 9 12 2 9 9 0 7 0 1 10 9 9 13 13 2
61 1 9 9 13 13 9 0 0 1 10 9 1 12 12 7 12 12 9 1 0 1 12 12 9 1 9 12 13 7 9 9 7 9 9 9 0 9 0 7 0 9 1 12 12 9 1 9 12 1 0 1 12 12 9 1 9 12 9 13 13 2
50 1 9 9 7 9 9 0 7 0 16 1 9 9 9 7 9 1 12 12 9 9 0 7 12 12 9 9 0 1 9 12 1 12 12 9 9 0 7 12 12 9 9 0 1 9 12 9 13 13 2
45 1 9 10 9 2 9 9 0 2 1 9 9 0 1 9 9 12 9 1 9 9 1 9 16 1 9 12 9 9 13 13 2 13 13 9 15 1 9 0 9 0 9 0 13 2
25 7 1 9 1 9 0 2 1 0 9 9 9 0 9 0 0 1 9 1 9 7 3 9 13 2
37 1 9 10 9 9 9 0 1 9 9 9 0 10 9 13 2 1 9 0 9 9 9 9 9 13 9 0 0 16 2 1 9 10 9 0 13 2
13 9 13 15 15 16 13 13 9 7 9 13 13 2
36 3 9 1 9 1 9 9 9 0 1 9 9 9 7 9 9 2 9 13 7 3 9 9 7 9 9 0 2 13 13 7 13 7 13 13 2
14 9 9 13 2 9 15 0 1 9 9 7 9 13 2
19 13 6 9 2 3 9 7 1 3 13 13 9 7 9 3 1 9 13 2
23 1 9 1 1 12 9 0 3 9 13 2 3 1 0 9 1 10 9 3 9 0 13 2
9 10 9 1 9 7 9 15 13 2
16 10 9 1 9 9 1 9 15 1 9 0 7 0 9 13 2
10 10 9 13 16 15 4 15 9 13 2
23 9 1 9 3 9 13 3 7 9 15 9 9 7 9 9 1 9 0 7 9 0 13 2
8 10 9 1 9 9 9 13 2
28 16 9 15 13 9 7 1 9 1 1 1 9 0 13 7 9 9 9 13 1 9 7 9 3 9 13 2 2
26 9 9 9 13 2 9 1 9 9 9 13 9 1 15 9 13 7 9 9 16 15 13 7 9 13 2
14 13 3 9 1 9 3 9 1 15 15 0 13 13 2
13 9 9 13 7 9 13 14 3 13 7 7 13 2
11 15 16 13 1 13 7 13 15 13 13 2
25 9 14 15 15 9 13 1 9 2 13 2 3 16 1 10 9 16 1 9 13 1 9 9 13 2
18 15 7 13 7 13 13 2 10 10 9 9 13 7 1 9 12 9 2
45 1 9 9 9 16 1 9 9 0 0 13 13 13 13 1 9 7 9 0 9 13 3 9 14 0 13 2 9 9 13 7 9 14 1 13 7 13 7 9 1 1 9 9 13 2
54 3 9 1 9 9 13 9 9 7 9 16 1 9 9 9 9 7 9 9 9 15 9 13 7 13 2 1 9 12 7 9 9 1 9 9 0 7 1 9 9 9 0 1 9 12 9 2 3 9 9 9 9 13 2
68 9 9 9 3 1 9 1 9 9 13 2 9 9 0 15 14 9 13 7 1 1 9 0 9 9 9 13 7 9 16 13 1 0 9 10 9 1 15 1 9 13 13 15 1 15 4 10 9 0 9 13 7 16 9 13 0 13 1 0 10 9 9 13 3 0 4 13 2
60 9 1 9 0 7 0 7 1 9 1 1 9 1 9 9 9 16 3 1 9 12 9 0 1 9 9 0 13 13 9 9 0 7 9 0 13 16 15 1 9 9 9 9 1 9 9 9 1 9 9 7 9 0 7 0 0 13 7 13 2
57 9 1 9 3 9 9 1 9 9 1 9 10 9 0 1 9 0 9 9 9 13 16 1 15 9 13 7 9 0 15 13 16 10 9 7 9 3 7 3 1 9 9 7 1 9 1 9 13 16 1 9 0 9 9 13 13 2
36 0 13 16 9 0 9 9 1 9 9 1 9 9 7 9 9 3 1 9 9 16 3 0 9 9 14 1 9 9 9 9 13 2 4 13 2
22 9 9 4 1 10 0 9 9 0 7 0 13 16 1 9 0 9 3 9 9 13 2
21 9 0 0 1 9 0 13 7 10 14 3 9 0 9 7 9 15 1 4 13 2
8 10 9 1 3 9 4 13 2
20 9 7 9 9 9 0 7 9 9 9 9 9 9 13 16 1 1 9 13 2
23 9 0 1 9 1 9 9 7 9 0 1 12 9 0 2 9 7 9 0 14 9 13 2
8 9 10 9 2 3 0 13 2
32 9 1 9 12 9 9 9 9 12 2 9 0 9 7 9 9 12 7 9 0 9 12 10 9 14 3 2 0 7 0 13 2
51 4 1 9 7 9 0 16 1 10 12 9 1 9 0 7 1 9 0 1 9 9 0 9 13 13 16 9 13 7 9 13 16 9 0 9 9 3 0 9 13 2 7 3 9 7 9 0 0 13 13 2
18 9 0 9 9 9 9 2 0 0 1 9 9 9 0 1 9 13 2
27 9 0 2 9 9 7 9 0 9 13 16 9 3 9 1 9 9 0 1 12 9 9 7 9 9 13 2
15 9 12 9 9 9 7 9 12 9 9 9 9 0 13 2
25 1 9 9 9 10 12 9 7 12 9 0 1 9 14 13 13 2 9 15 14 1 9 9 13 2
55 3 9 16 9 10 9 14 1 9 1 9 9 9 7 9 13 16 1 12 9 0 1 9 13 13 1 9 1 9 0 7 1 9 1 9 0 7 9 2 9 0 1 9 0 14 3 1 9 9 7 9 15 9 13 2
29 9 0 9 0 7 9 7 9 9 9 1 9 1 9 9 0 2 0 2 9 9 9 0 1 10 9 13 13 2
51 10 9 13 16 1 9 9 0 1 9 9 1 9 9 9 0 14 13 9 13 2 1 9 7 9 9 0 7 0 9 15 3 1 0 9 9 13 16 9 0 0 1 9 2 1 15 0 7 0 13 2
26 1 9 0 2 3 12 9 0 1 9 1 9 0 9 7 1 9 9 7 9 1 9 0 9 13 2
21 9 0 2 3 1 1 9 7 9 13 1 1 9 0 1 9 0 9 0 13 2
16 9 0 0 16 1 9 9 9 13 2 10 9 14 9 13 2
39 7 9 0 9 0 2 0 1 9 7 9 0 7 0 7 9 0 2 0 16 9 2 9 2 9 7 9 9 9 9 9 7 9 0 1 9 9 13 2
23 10 9 7 9 9 9 3 13 16 9 0 2 9 13 2 3 9 7 9 7 9 0 2
23 1 9 9 2 1 9 0 2 4 1 12 9 0 7 0 1 1 9 7 9 0 13 2
18 9 7 9 0 4 1 1 9 7 9 1 9 0 1 9 0 13 2
27 10 9 16 9 1 9 0 2 1 9 9 0 7 0 2 9 13 2 3 13 9 0 1 1 13 13 2
26 9 9 9 9 2 1 9 9 7 9 9 7 9 15 1 9 0 9 7 9 0 15 14 9 13 2
41 9 0 7 9 0 9 16 9 0 7 0 1 9 9 13 7 1 9 7 9 9 1 9 7 9 1 9 7 9 15 13 2 9 0 1 10 9 1 9 13 2
28 7 1 9 9 7 9 1 9 0 7 0 13 2 10 9 2 9 7 9 0 7 0 14 0 7 0 13 2
5 9 9 14 13 2
43 9 9 1 9 9 0 15 13 13 2 9 9 9 9 0 9 9 9 9 1 9 0 3 9 0 1 1 9 16 1 1 9 0 7 9 9 9 0 9 13 9 13 2
50 15 1 9 3 1 9 9 13 2 3 9 0 7 9 9 0 9 0 1 9 9 1 9 9 13 7 1 1 9 0 7 9 0 7 9 9 0 9 0 1 9 9 9 7 9 7 9 9 13 2
36 9 9 9 9 13 2 15 1 9 9 7 15 9 9 7 9 1 9 0 7 15 9 7 9 9 7 9 9 13 16 16 9 9 14 13 2
61 15 13 2 9 13 16 9 0 13 1 9 1 9 12 9 0 2 9 1 9 9 7 9 9 14 1 9 9 13 1 9 7 9 12 9 0 1 12 9 1 9 0 0 2 0 2 0 7 0 1 9 9 0 7 9 0 9 0 9 13 2
45 9 9 9 13 2 15 1 10 9 9 9 13 16 9 12 16 0 9 9 0 14 13 1 13 9 9 9 0 14 16 9 9 1 10 9 0 13 2 1 3 9 0 9 13 2
14 9 9 9 1 9 9 12 9 9 9 9 13 13 2
40 1 9 3 9 9 9 9 9 9 7 9 9 9 9 9 9 12 9 1 9 0 9 9 9 9 9 14 13 7 9 9 1 9 12 9 15 9 0 13 2
49 9 12 9 10 9 1 9 9 9 9 9 9 13 13 7 3 9 1 9 9 16 9 1 9 0 1 9 12 9 10 9 9 0 13 2 1 9 1 15 7 9 0 1 10 12 9 9 13 2
15 1 9 1 12 12 9 7 0 15 1 9 0 9 13 2
26 0 9 0 9 7 9 9 9 9 0 2 9 7 9 1 9 9 9 0 9 9 1 9 0 13 2
17 1 10 9 0 2 12 9 2 9 7 9 9 9 9 9 13 2
51 10 9 1 9 3 9 9 1 9 9 7 9 9 1 9 0 9 9 7 9 9 9 9 7 9 9 9 0 1 9 0 0 0 13 7 12 9 1 9 0 9 2 9 2 9 7 9 9 9 13 2
15 9 0 9 9 1 9 9 9 2 1 9 9 9 13 2
32 1 9 10 9 16 1 9 9 9 13 7 9 9 9 15 12 9 13 9 12 9 9 9 1 9 9 9 9 7 9 13 2
15 9 9 1 10 9 9 13 1 9 9 3 1 9 13 2
30 9 9 0 9 9 7 9 7 9 7 9 13 2 9 9 0 1 9 9 1 9 0 1 9 9 9 9 9 13 2
23 9 9 13 2 10 9 0 0 16 0 9 9 7 9 13 1 9 9 9 3 13 13 2
24 15 13 2 9 2 1 9 7 9 9 9 10 9 3 9 15 14 1 9 9 1 9 13 2
18 9 0 13 2 9 9 0 7 9 0 1 9 10 9 0 13 13 2
32 1 9 15 2 1 9 1 9 9 9 9 2 9 0 9 1 9 0 9 13 2 16 9 9 0 9 1 10 9 0 13 2
34 9 0 13 2 3 1 9 9 9 7 9 9 0 9 2 9 9 7 9 15 1 9 9 9 0 2 9 7 9 0 9 9 13 2
18 12 9 1 9 9 2 12 9 0 14 1 9 0 1 9 9 13 2
21 1 9 10 9 16 9 15 1 9 3 7 3 9 13 2 12 9 9 9 13 2
16 15 9 9 9 0 0 1 9 9 0 9 9 9 13 13 2
27 9 9 12 12 7 12 12 9 9 1 9 0 13 16 10 9 1 0 1 12 12 9 9 0 9 13 2
20 9 7 9 9 0 9 1 12 9 0 1 9 9 9 0 7 0 9 13 2
35 9 9 9 0 7 0 9 0 13 2 10 9 16 1 9 9 9 9 13 1 9 9 2 9 0 7 9 9 0 3 0 2 9 13 2
42 9 9 9 13 2 1 9 0 7 9 9 0 9 3 1 9 0 9 9 13 16 10 9 1 9 1 9 9 9 2 9 9 10 9 14 16 1 9 0 9 13 2
34 1 9 9 0 9 1 9 9 9 2 9 0 0 7 9 0 9 13 7 0 9 15 9 9 9 1 9 0 7 9 9 9 13 2
11 9 9 1 9 9 9 1 9 0 13 2
45 1 10 9 16 1 9 9 9 9 7 9 1 9 1 9 9 13 2 9 1 9 9 9 16 9 15 9 2 9 7 9 9 9 13 2 1 10 9 9 7 9 0 9 13 2
42 9 9 1 9 1 9 7 1 9 1 10 9 16 9 10 9 13 1 9 7 9 9 10 9 13 2 13 2 9 0 1 9 0 7 0 0 9 7 9 13 13 2
12 16 9 0 16 4 0 1 9 0 3 13 2
24 15 13 2 1 1 9 0 1 9 3 2 9 0 16 4 1 9 9 7 9 0 9 13 2
28 9 9 1 9 1 10 9 16 9 9 9 9 15 13 2 13 2 9 0 9 9 9 2 9 7 9 13 2
23 9 9 1 9 10 9 2 1 9 9 0 9 1 9 7 10 9 15 1 9 9 13 2
8 9 9 1 9 1 9 13 2
29 9 9 9 9 0 9 9 16 1 12 1 9 9 9 9 1 9 0 2 1 9 9 1 0 9 2 9 13 2
29 10 9 16 1 9 0 1 12 1 9 9 0 1 9 9 1 9 13 13 2 9 13 9 15 1 9 9 13 2
32 9 16 1 10 9 9 13 2 13 10 9 1 9 9 16 1 10 9 1 9 1 13 13 2 9 0 14 1 15 9 13 2
45 1 13 7 9 16 1 0 9 1 9 10 9 1 9 13 2 9 0 9 9 9 2 9 9 9 0 10 9 1 9 9 2 7 9 0 9 0 2 1 9 7 9 9 13 2
12 9 1 9 0 1 9 0 1 9 1 13 2
30 12 9 1 9 0 7 0 9 0 0 0 1 9 0 3 1 9 1 9 0 1 9 9 0 9 1 9 1 13 2
37 10 9 1 9 12 9 0 1 9 1 9 9 9 9 13 16 0 9 10 9 1 9 9 2 0 7 1 9 0 9 3 0 1 9 9 13 2
18 1 10 9 9 9 9 7 9 1 1 12 9 1 9 0 9 13 2
23 9 0 1 10 9 0 9 0 0 9 1 9 12 9 13 16 9 9 9 9 0 13 2
40 1 9 9 0 9 9 0 9 2 9 0 10 9 0 14 9 0 1 9 9 2 9 2 9 2 9 7 2 1 9 0 1 9 9 1 12 9 9 13 2
37 10 9 16 0 9 0 0 2 0 2 0 2 0 2 0 7 15 16 0 9 13 7 1 1 12 9 7 1 9 12 9 1 9 9 9 13 2
22 9 0 9 13 16 9 9 0 0 1 9 7 9 13 16 0 1 9 15 13 13 2
30 10 9 9 1 9 12 0 1 9 9 7 9 9 0 9 9 13 7 1 9 9 0 1 9 9 9 9 4 13 2
6 9 9 9 9 13 2
27 9 9 9 0 9 9 9 9 0 0 7 12 9 0 1 9 0 9 9 12 9 9 0 9 9 13 2
36 1 9 9 9 9 2 9 9 7 9 15 0 9 12 1 9 0 9 12 9 9 0 0 9 0 9 14 1 9 9 1 15 9 13 13 2
21 9 10 9 1 9 0 12 9 9 7 12 9 0 9 1 9 9 12 9 13 2
20 0 9 0 1 9 9 16 1 9 0 1 9 15 9 13 13 2 9 13 2
22 9 16 1 0 9 2 0 9 2 0 9 9 2 0 9 7 0 9 9 13 13 2
53 9 9 9 9 9 9 3 3 1 9 12 1 9 9 2 9 7 9 9 9 0 13 13 7 12 1 0 9 0 1 10 9 1 9 13 16 4 15 14 1 9 9 0 7 9 12 9 1 12 9 9 13 2
19 12 7 0 9 0 9 9 9 1 10 9 2 3 1 9 9 9 13 2
23 1 9 9 9 9 2 12 9 9 9 9 7 9 1 9 0 7 0 10 9 9 13 2
30 9 9 9 1 9 9 9 9 0 0 9 1 9 12 7 0 9 13 16 1 9 12 9 0 9 9 9 4 13 2
37 1 9 9 9 2 12 9 1 9 9 0 9 0 1 9 9 9 2 1 9 9 9 9 13 16 1 9 12 9 9 10 9 1 9 1 13 2
49 9 9 0 9 16 9 9 1 15 13 7 9 0 1 10 9 16 1 15 9 0 13 13 7 9 9 7 9 7 9 9 9 1 9 7 9 7 10 9 0 14 4 1 9 0 9 9 13 2
40 9 0 2 9 9 9 9 9 7 9 9 10 9 1 9 0 9 1 9 9 9 0 0 2 9 1 9 9 7 1 9 7 9 1 9 9 9 13 13 2
21 1 10 9 16 16 9 0 9 9 7 9 1 9 13 13 2 9 9 4 13 2
42 7 9 10 9 9 9 7 9 0 13 1 9 9 16 1 3 9 7 9 0 2 0 9 1 10 9 9 9 0 13 13 7 16 10 9 9 0 15 14 9 13 2
45 7 1 9 0 9 7 9 1 9 7 9 9 9 0 1 9 0 13 16 9 3 9 1 9 7 9 1 9 7 9 0 1 13 7 9 1 15 9 9 7 9 1 9 13 2
18 1 1 9 0 16 9 9 2 9 2 1 9 0 7 0 9 13 2
24 1 0 9 9 13 7 15 13 9 9 2 9 2 3 10 9 14 0 13 7 1 9 13 2
51 3 16 9 13 9 9 13 9 0 9 9 2 9 2 14 1 1 13 1 16 2 9 7 9 15 1 9 9 2 9 2 9 9 13 7 16 15 9 9 2 9 2 7 9 15 1 9 9 0 13 2
19 1 10 9 1 9 7 9 9 7 9 9 9 2 9 2 14 9 13 2
29 16 9 9 1 9 9 2 9 2 14 13 13 2 1 3 7 9 9 13 2 9 9 2 9 2 1 15 13 2
13 1 9 9 9 9 14 1 9 15 13 7 13 2
15 9 13 13 1 1 9 9 3 9 1 1 9 13 13 2
14 9 9 2 9 2 13 2 10 9 1 15 13 9 2
20 9 0 16 3 9 9 9 2 7 9 9 14 9 13 2 9 9 9 13 2
33 9 1 9 16 9 7 9 2 9 2 7 9 7 9 1 9 13 1 1 9 9 9 13 2 1 9 9 2 9 2 9 13 2
12 9 9 2 9 2 2 9 16 1 9 13 2
31 9 9 9 9 2 9 2 16 3 9 9 14 1 9 13 2 9 13 16 9 9 0 1 15 7 9 7 9 15 13 2
20 3 7 9 2 1 9 7 9 9 9 1 1 9 9 2 9 2 9 13 2
38 9 9 2 9 2 1 15 13 2 6 9 16 1 15 15 9 13 2 1 9 15 9 13 2 3 1 9 15 7 9 16 9 15 14 13 9 13 2
15 10 9 16 15 7 9 15 2 9 2 15 14 9 13 2
25 9 9 7 9 16 1 9 9 2 9 2 1 10 9 1 9 9 1 9 13 13 3 0 13 2
30 10 9 0 9 3 9 13 16 9 9 2 9 2 1 9 13 2 9 9 9 0 13 7 3 9 15 9 13 13 2
35 3 7 3 1 9 9 7 9 1 9 2 1 10 9 12 1 12 9 12 9 10 9 12 1 9 9 2 9 2 9 1 9 13 13 2
21 9 7 9 15 13 1 9 0 7 9 0 9 9 2 9 2 14 1 9 13 2
25 3 1 9 13 16 9 9 2 9 2 14 3 9 9 9 2 9 2 16 1 9 0 0 13 2
25 3 1 9 9 9 9 2 9 2 9 1 9 13 13 2 3 9 1 9 2 9 2 3 13 2
15 9 9 0 16 0 1 9 9 13 15 14 1 9 13 2
24 10 9 7 9 1 9 0 0 9 9 2 9 2 1 9 7 9 9 14 3 0 13 13 2
41 9 9 2 9 2 0 13 3 1 15 1 9 16 9 13 1 9 9 1 9 7 9 9 1 9 9 2 9 2 13 2 3 9 13 7 9 15 14 0 13 2
14 3 7 9 9 2 9 2 1 9 12 9 9 13 2
29 9 9 13 16 15 9 0 13 7 9 9 7 9 2 9 9 2 9 2 13 2 1 9 9 1 15 9 13 2
29 3 7 9 2 9 2 1 9 9 9 7 9 9 9 9 13 7 13 2 9 15 14 1 9 1 15 9 13 2
29 10 9 1 9 13 16 0 1 9 9 9 2 9 2 3 15 16 1 9 9 7 9 9 13 13 9 9 13 2
13 9 9 9 2 9 2 1 9 9 9 9 13 2
6 9 0 7 0 13 2
13 9 9 2 9 2 9 9 7 9 15 14 13 2
8 13 2 12 12 9 9 13 2
13 9 9 2 9 2 13 2 9 15 1 9 15 2
3 9 13 2
9 9 13 2 13 1 10 9 13 2
24 9 9 2 9 2 13 2 3 1 15 7 1 9 13 9 15 14 13 7 10 9 14 13 2
19 9 9 9 2 9 2 1 9 2 3 9 9 15 9 2 9 2 13 2
11 0 13 16 9 1 9 15 9 0 13 2
16 9 16 3 13 1 10 9 1 9 9 7 9 15 9 13 2
30 12 9 16 9 9 2 9 2 3 1 9 9 13 13 2 9 13 16 9 9 9 14 1 9 9 2 9 2 13 2
17 10 9 2 1 9 9 2 9 2 12 9 13 7 12 9 0 2
25 9 2 9 2 1 9 15 0 9 9 13 13 2 7 9 14 9 9 9 7 8 8 13 13 2
15 9 9 2 9 2 13 2 9 9 14 1 3 9 13 2
39 9 9 10 9 14 16 13 16 13 9 9 2 9 2 14 1 12 9 0 9 13 16 9 0 1 9 9 14 0 13 7 9 15 14 3 9 13 13 2
31 10 9 0 9 13 1 9 9 0 9 2 9 2 2 9 9 9 9 16 1 10 9 9 9 9 9 2 9 2 13 2
22 1 9 9 16 9 1 9 9 15 1 9 13 2 1 9 9 2 9 2 9 13 2
28 1 9 9 2 9 2 13 2 16 9 9 15 1 9 7 9 7 9 15 7 9 9 15 1 15 13 13 2
13 9 9 2 9 2 13 2 1 15 3 9 13 2
16 9 13 2 15 14 13 2 9 15 13 7 1 15 9 13 2
13 9 9 2 9 2 13 2 10 9 9 15 13 2
20 7 15 16 9 15 14 13 2 15 14 9 7 9 13 7 1 15 9 13 2
18 10 9 9 0 7 0 12 9 9 7 9 2 7 9 7 9 13 2
20 7 7 9 0 1 9 9 2 16 9 0 0 3 9 9 9 14 9 13 2
13 1 9 0 15 14 9 13 7 1 15 9 13 2
18 10 9 9 2 9 9 9 13 7 9 9 9 9 9 2 9 15 2
24 9 9 9 13 16 1 9 9 9 2 9 2 9 15 1 9 2 0 7 9 15 0 13 2
20 1 9 9 16 9 0 7 0 1 1 9 2 9 2 7 9 15 9 13 2
35 9 0 2 1 9 9 16 9 0 9 9 1 9 13 13 2 9 9 2 9 13 2 9 9 14 0 0 13 7 9 15 14 3 13 2
20 7 9 2 9 9 14 1 9 13 2 1 9 0 7 0 15 9 0 13 2
14 9 16 1 9 9 1 9 9 13 7 13 2 13 2
33 7 3 16 9 9 9 13 13 1 9 9 9 13 7 13 2 6 8 9 10 9 16 1 15 9 13 3 1 9 9 15 13 2
11 9 10 9 13 16 3 9 9 13 13 2
18 9 9 14 1 9 9 13 16 9 9 9 9 2 9 2 14 13 2
16 9 9 15 14 13 7 9 7 9 13 7 1 15 9 13 2
15 10 9 9 9 7 9 9 2 9 2 1 10 9 13 2
10 0 13 9 1 9 9 7 9 13 2
42 15 1 9 1 9 9 1 9 2 3 1 15 7 9 9 14 9 13 7 9 13 2 1 9 1 9 13 2 1 1 9 7 9 7 9 7 9 1 15 0 13 2
8 9 15 1 9 9 13 13 2
14 9 16 9 1 9 9 13 7 9 1 15 0 13 2
18 9 9 9 1 9 9 9 2 9 2 9 0 7 0 14 9 13 2
26 9 9 2 9 2 9 9 14 1 9 9 9 13 2 9 15 1 10 9 16 13 2 1 9 13 2
19 1 9 15 7 9 13 9 1 9 15 13 9 7 9 15 14 9 13 2
27 16 9 9 13 16 9 15 13 2 15 14 1 9 13 2 9 15 14 9 13 7 9 15 14 0 13 2
41 9 9 9 0 13 16 10 9 9 13 2 15 14 13 7 1 9 13 2 9 7 9 9 14 9 13 2 9 3 0 1 15 0 13 2 7 1 15 9 13 2
9 9 9 9 9 9 9 9 13 2
15 1 9 9 2 9 1 9 9 1 9 9 9 9 13 2
15 9 9 13 10 9 14 0 13 7 9 15 14 9 13 2
8 9 1 9 1 9 9 13 2
12 9 13 2 15 3 9 14 9 7 9 13 2
9 7 9 15 14 1 9 9 13 2
19 10 9 3 1 9 9 16 9 13 13 2 3 3 0 7 1 9 0 2
45 3 7 9 9 9 1 9 9 1 9 9 9 7 9 9 13 7 1 9 9 1 9 9 9 9 9 13 2 7 1 9 15 9 9 13 2 9 3 9 13 9 9 14 13 2
18 7 9 14 16 9 13 1 9 15 9 13 2 9 15 14 9 13 2
15 1 9 9 9 9 9 12 9 7 12 9 14 9 13 2
21 9 15 3 9 14 9 7 9 13 7 10 9 14 1 9 7 9 13 2 13 2
21 1 9 9 13 16 9 1 9 1 9 9 2 9 2 3 1 9 15 9 13 2
14 9 14 0 13 7 9 15 14 1 9 1 9 13 2
16 7 7 9 9 0 1 9 7 9 14 1 1 9 9 13 2
26 0 1 12 9 1 9 2 9 7 9 9 0 9 1 9 9 9 15 1 9 0 9 14 9 13 2
45 1 9 1 9 1 15 7 9 7 9 0 3 10 9 0 13 1 9 9 7 9 7 9 7 9 13 2 9 9 0 7 9 3 9 1 0 9 9 7 9 9 9 13 13 2
46 9 9 9 13 2 9 7 9 15 0 1 9 9 7 9 0 9 0 2 9 2 13 7 13 16 3 9 16 9 0 2 9 2 9 13 1 9 0 12 9 1 9 0 0 13 2
35 9 2 0 9 9 1 9 3 9 14 9 0 7 9 0 7 9 0 9 9 1 9 9 7 9 7 9 9 7 9 0 9 13 13 2
52 9 7 9 16 1 9 9 9 7 1 9 9 13 13 2 9 9 7 9 15 14 0 13 13 7 10 9 0 0 13 7 0 2 9 0 13 7 3 9 0 7 9 0 7 9 0 14 4 0 9 13 2
39 10 9 0 13 2 9 1 9 0 9 0 1 9 7 9 0 9 0 1 9 7 9 9 7 9 7 9 0 13 7 9 16 9 10 12 9 0 13 2
36 9 9 9 13 2 9 9 9 1 9 9 16 9 14 0 13 7 10 12 9 0 15 14 0 13 9 1 1 9 9 9 7 9 0 13 2
51 9 13 2 15 16 3 9 9 9 7 9 7 9 14 13 4 0 1 15 1 9 13 7 3 3 9 7 0 2 9 7 9 14 1 3 16 9 9 7 9 0 7 0 9 13 1 0 7 9 13 2
40 9 1 9 0 9 7 9 9 0 7 0 9 9 9 9 9 9 1 9 9 0 9 13 16 0 9 7 9 13 16 1 9 9 9 7 9 9 13 13 2
28 9 9 1 9 0 1 15 7 12 9 0 1 0 9 9 13 2 10 9 0 14 9 9 7 9 13 13 2
86 10 12 9 14 10 9 9 13 13 2 9 16 3 9 14 0 13 7 3 0 9 14 7 15 14 9 1 9 9 1 9 0 7 9 1 9 9 9 0 0 13 7 13 2 7 9 0 16 8 1 9 9 7 9 9 1 9 13 7 3 7 3 1 9 1 0 9 13 7 10 9 0 14 9 1 0 7 9 9 9 7 0 9 9 13 2
34 9 1 0 9 1 9 0 7 0 12 9 9 13 7 13 16 10 9 0 7 9 0 10 1 0 9 1 3 9 7 9 0 13 2
48 0 9 9 0 13 16 1 9 9 0 0 13 7 9 7 9 1 15 1 9 7 9 0 13 7 1 1 9 9 9 7 9 13 9 9 0 16 1 9 9 0 9 0 7 0 13 13 2
31 1 9 9 10 9 2 15 0 1 15 9 0 7 0 13 2 9 9 1 1 9 0 7 9 0 7 9 9 0 13 2
45 1 9 10 9 9 13 13 2 9 0 9 3 9 0 9 7 9 9 9 13 7 1 9 9 1 9 0 7 9 9 0 9 13 7 3 0 9 0 13 7 1 9 9 13 2
59 9 3 9 1 9 16 15 14 9 7 9 0 9 9 13 0 13 2 13 9 15 14 1 9 16 3 3 9 1 9 7 9 7 9 13 2 3 1 9 15 9 0 1 9 1 9 13 7 9 15 1 15 7 15 12 13 0 13 2
43 1 10 9 13 13 2 9 0 7 9 0 16 9 9 9 7 9 1 9 0 13 2 16 15 9 0 9 13 1 9 1 9 13 16 13 9 9 0 15 13 7 3 2
30 9 13 2 9 9 9 1 9 7 9 7 9 7 9 3 1 9 0 9 9 9 1 9 0 7 9 1 9 13 2
35 9 9 13 13 2 9 7 9 4 3 0 9 13 16 1 9 0 9 9 0 13 2 9 7 0 7 9 7 9 0 9 9 0 13 2
49 9 1 9 10 9 16 3 15 9 1 9 7 9 1 9 9 9 13 9 13 16 1 10 9 3 4 9 7 9 7 9 9 3 0 7 0 7 0 1 9 13 16 15 4 1 15 9 13 2
41 9 16 1 9 7 1 9 0 1 9 13 7 15 9 7 9 9 1 15 9 13 2 3 0 7 0 1 9 0 7 0 13 16 9 0 14 1 9 13 13 2
32 9 13 13 2 9 7 9 7 9 9 0 9 3 13 16 9 0 14 1 9 13 7 3 9 15 16 9 1 9 15 13 2
16 0 9 16 16 9 13 16 9 13 16 1 9 9 9 13 2
27 16 3 1 9 1 9 0 7 0 9 13 7 16 0 1 9 9 0 9 0 9 0 13 1 9 9 2
58 9 9 9 1 9 13 2 9 0 7 0 9 0 13 7 0 7 13 16 9 7 9 15 1 9 0 9 1 9 9 9 7 9 9 1 1 15 13 3 1 1 15 2 7 9 9 0 14 1 9 13 16 8 8 8 8 8 2
38 1 9 10 9 12 0 9 9 13 13 16 9 9 10 9 14 9 7 9 9 13 7 9 9 14 1 9 9 9 13 7 9 14 0 7 0 13 2
42 1 0 9 0 9 9 9 2 9 9 3 0 13 2 1 9 7 9 1 9 12 9 1 9 0 9 0 12 1 9 9 0 12 9 9 13 7 1 9 0 13 2
50 1 9 0 9 9 9 16 9 9 1 9 9 0 9 9 0 13 3 1 9 9 9 9 7 9 16 10 12 1 9 9 9 9 0 13 1 9 0 7 0 9 13 7 9 1 9 0 9 13 2
20 9 9 1 9 0 1 9 9 9 1 9 12 9 1 9 0 0 13 13 2
13 7 9 9 1 12 9 9 1 9 0 0 13 2
23 0 9 14 1 10 9 9 9 1 12 9 9 13 16 1 9 12 7 0 9 13 13 2
25 9 1 9 10 9 3 12 9 0 0 12 9 0 1 9 9 0 12 14 9 9 9 13 13 2
30 1 9 9 9 9 7 9 9 9 1 9 9 10 9 2 9 0 9 1 9 0 1 9 9 9 9 9 9 13 2
55 9 9 2 9 9 9 0 1 9 9 9 9 13 2 1 9 9 0 9 1 9 7 9 15 1 9 1 10 9 2 9 9 1 9 0 9 9 9 7 1 9 0 9 9 2 1 9 0 9 9 9 9 9 13 2
63 15 13 2 9 1 10 9 1 9 0 9 13 7 1 15 1 9 1 9 9 2 1 12 9 0 16 10 9 9 13 0 9 9 9 7 9 7 9 0 0 13 13 16 9 13 1 9 10 9 0 9 4 3 9 9 1 9 9 0 0 9 13 2
27 9 9 9 9 9 9 1 9 9 9 1 9 1 9 9 9 9 9 9 9 0 9 1 9 9 13 2
25 10 9 1 9 12 1 12 9 9 0 1 9 9 0 13 7 1 15 9 12 9 9 4 13 2
36 9 9 9 9 9 9 16 1 9 9 13 13 2 1 9 1 9 9 9 9 1 9 0 9 10 9 1 9 1 9 0 9 1 9 13 2
12 10 9 1 12 9 9 7 9 0 4 13 2
21 9 9 9 9 12 9 9 9 9 1 9 9 9 1 9 9 1 9 9 13 2
21 9 0 9 9 0 1 9 0 1 9 0 9 9 9 0 1 9 9 9 13 2
21 1 9 0 9 10 9 9 0 9 0 1 9 9 9 1 9 1 9 1 13 2
33 3 1 15 2 9 12 7 12 0 9 9 1 9 9 9 13 16 1 9 10 9 12 9 9 9 9 15 14 1 9 4 13 2
57 9 9 9 9 9 9 0 9 13 16 9 9 14 1 9 13 2 15 1 9 13 16 9 9 9 9 9 1 9 9 4 13 16 9 9 10 9 1 9 9 7 9 15 1 9 9 9 9 9 12 9 14 1 9 4 13 2
29 1 9 9 9 0 9 9 12 9 1 9 9 9 9 12 9 1 9 9 7 1 9 12 9 0 9 4 13 2
10 9 9 9 12 9 9 14 9 13 2
34 9 0 9 9 0 1 9 9 2 9 9 9 12 9 9 3 1 9 9 14 9 13 7 9 9 14 1 9 10 9 1 9 13 2
17 9 9 0 1 10 9 1 9 0 0 9 7 9 0 9 13 2
38 9 9 15 1 9 0 1 9 0 1 9 13 7 15 14 1 9 1 0 9 3 0 1 9 9 1 9 9 9 16 12 9 9 13 2 0 13 2
20 9 9 16 9 9 1 9 0 9 13 2 0 9 0 1 9 1 9 13 2
34 0 9 9 15 13 16 12 12 7 12 12 9 9 9 0 1 9 1 9 13 16 1 9 1 9 3 1 15 12 9 0 13 13 2
29 9 9 0 9 9 9 13 16 9 9 9 1 9 7 9 9 0 9 2 1 9 9 9 9 9 1 9 13 2
22 1 10 9 2 9 0 1 0 9 1 9 9 9 9 9 0 1 9 9 13 13 2
29 9 9 9 9 13 2 12 9 0 0 1 9 9 2 12 1 9 9 1 9 0 9 1 9 9 9 13 13 2
19 9 1 15 9 13 16 16 9 9 13 2 9 0 0 0 9 4 13 2
59 9 0 9 2 12 1 9 9 9 1 9 0 9 0 13 7 1 10 9 2 10 9 0 0 0 1 9 10 9 0 0 13 13 7 9 15 13 16 3 1 9 1 9 9 9 13 7 9 9 9 9 1 9 9 9 14 0 13 2
19 10 9 1 9 0 1 9 9 0 1 9 9 9 0 9 2 12 13 2
26 9 1 9 0 9 13 1 12 9 9 7 9 9 9 3 9 13 13 7 1 9 10 12 9 13 2
32 9 9 9 13 13 16 9 9 1 10 12 9 1 9 0 7 9 0 1 9 0 13 7 1 12 9 9 7 9 0 13 2
10 3 9 9 1 15 13 7 9 13 2
22 10 9 1 9 9 0 12 9 9 7 9 1 9 9 1 9 1 9 10 9 13 2
23 12 1 9 9 9 1 9 9 9 0 9 7 9 14 9 13 7 1 10 9 9 13 2
13 12 9 0 0 9 0 10 9 14 9 13 13 2
33 9 9 9 14 9 13 13 16 1 9 15 4 9 0 14 9 13 7 1 1 15 1 9 0 9 7 9 0 16 1 9 13 2
24 10 9 9 1 9 0 0 13 7 3 1 9 0 9 1 9 4 10 9 14 1 9 13 2
40 9 16 1 10 9 9 13 2 13 1 12 9 9 9 9 1 9 9 9 7 9 0 16 9 13 7 3 9 9 0 14 16 1 9 1 9 9 9 13 2
18 9 9 9 9 2 9 0 1 9 0 1 9 0 1 9 9 13 2
36 9 9 1 10 13 7 13 9 13 2 16 9 0 9 0 1 9 1 9 9 9 9 9 9 0 13 2 9 12 9 1 9 0 4 13 2
26 9 9 13 2 9 0 4 1 12 9 9 7 3 1 9 9 1 10 9 2 1 9 15 9 13 2
21 0 1 9 9 9 9 1 9 16 1 9 9 9 9 9 13 2 0 9 13 2
18 9 0 9 9 9 9 9 9 1 9 9 7 9 7 9 15 13 2
41 9 9 9 9 9 9 9 9 13 2 1 9 9 9 0 0 9 16 3 9 9 1 9 0 0 15 14 9 13 13 2 4 10 9 14 1 9 0 9 13 2
38 9 10 9 1 12 9 10 9 9 0 13 13 7 10 9 1 15 7 0 9 7 9 9 9 9 13 2 1 9 10 9 13 9 0 14 9 13 2
33 0 1 12 12 9 1 9 0 9 9 9 1 9 0 13 7 9 9 9 0 15 7 9 9 2 9 2 1 9 9 9 13 2
21 1 9 9 9 1 9 2 9 12 9 1 12 9 0 9 1 10 9 9 13 2
12 0 9 0 9 0 0 1 12 12 9 13 2
23 9 9 1 1 9 9 9 9 1 1 0 9 9 1 9 9 1 9 9 9 9 13 2
42 9 9 9 9 13 2 9 9 9 12 9 3 1 9 1 9 9 9 9 13 7 3 9 0 1 1 9 7 9 7 9 9 0 1 9 10 9 1 9 13 13 2
22 1 9 9 0 9 2 1 9 0 9 9 9 9 9 2 12 9 0 3 9 13 2
21 9 9 9 13 2 12 9 9 9 0 7 0 7 9 9 0 10 9 9 13 2
41 1 9 9 2 10 12 9 1 9 9 15 14 1 9 9 13 16 9 9 0 0 7 12 9 9 0 1 9 9 9 1 12 9 1 9 1 9 0 9 13 2
11 1 9 0 9 9 9 0 9 0 13 2
17 9 9 9 0 9 10 9 1 9 9 9 10 9 14 13 13 2
38 9 9 16 1 3 9 12 9 14 1 9 9 13 13 2 9 13 2 1 9 13 9 0 1 9 15 9 13 16 9 9 9 1 9 9 9 13 2
26 9 10 9 16 1 9 9 0 13 2 13 2 16 13 9 15 14 1 9 13 3 10 9 14 13 2
24 0 9 10 9 9 9 9 13 16 9 9 9 9 12 14 1 9 12 1 9 9 9 13 2
43 3 1 9 9 0 3 2 9 15 1 1 9 9 3 9 1 9 9 9 16 9 3 1 15 1 12 9 10 9 9 13 13 7 3 12 9 15 14 9 13 2 13 2
69 12 1 9 1 10 9 1 9 15 13 16 3 1 9 9 0 9 9 9 0 9 1 9 1 9 9 9 15 14 1 10 9 9 13 7 9 9 12 9 10 9 13 1 10 9 1 12 9 0 7 9 9 9 7 9 9 9 9 1 15 1 3 9 1 9 0 0 13 2
28 9 9 16 1 0 10 9 7 9 9 9 9 9 1 1 9 9 9 12 9 10 9 9 0 14 9 13 2
38 9 9 1 10 9 13 13 2 1 12 1 0 9 9 9 0 2 12 9 9 9 9 9 9 1 9 9 1 9 9 9 0 7 1 9 9 13 2
53 1 9 10 9 1 9 9 9 9 9 9 2 9 0 1 9 9 1 9 9 0 7 0 9 13 16 9 15 1 9 9 9 0 9 1 15 0 13 7 9 7 9 9 9 9 9 3 1 10 9 0 13 2
60 15 0 13 9 9 1 9 9 0 9 0 9 15 1 9 9 9 9 13 7 13 1 10 9 7 9 0 15 7 1 9 9 9 13 2 7 1 10 9 9 0 9 13 1 10 9 9 9 1 9 9 7 9 9 9 15 9 13 13 2
65 9 0 9 3 9 9 0 16 1 9 0 0 2 3 1 9 12 9 9 2 9 0 7 9 0 1 9 7 9 9 7 9 0 9 9 0 13 4 1 9 9 9 1 9 9 2 3 1 9 9 13 16 9 7 9 0 7 0 1 9 1 9 13 13 2
11 0 9 7 9 1 9 9 10 9 13 2
26 1 9 7 0 12 9 1 9 0 9 0 9 13 13 2 9 3 9 1 9 0 3 9 4 13 2
64 16 9 9 13 16 13 3 1 9 9 7 9 0 1 15 13 13 7 3 10 9 0 0 13 16 1 10 9 3 3 9 13 13 16 9 9 9 1 0 9 9 9 15 1 9 9 13 16 4 1 12 9 0 7 0 1 1 15 9 7 9 9 13 2
29 1 10 9 9 12 9 1 9 0 16 1 9 9 9 9 9 9 1 9 9 0 13 2 1 3 9 0 13 2
55 1 9 7 0 1 12 9 1 9 9 0 9 13 7 9 9 4 1 1 9 0 9 9 12 9 0 14 16 9 15 1 9 0 13 13 0 13 2 3 1 9 9 15 1 9 2 15 14 1 9 0 15 1 13 2
75 9 9 16 1 9 1 9 13 13 2 1 9 12 0 9 9 9 9 9 16 9 9 9 9 13 2 1 9 9 9 13 16 9 7 9 0 1 9 13 2 1 9 7 9 0 9 9 9 3 1 9 10 9 9 13 2 13 13 9 9 1 9 1 9 10 9 16 0 13 2 1 9 3 13 2
59 9 9 9 9 9 3 1 9 9 1 10 9 1 9 15 13 2 9 9 1 10 9 0 13 7 9 10 9 14 1 9 0 13 2 16 16 9 1 9 9 10 9 9 13 2 1 9 1 9 15 1 9 0 9 1 9 9 13 2
19 9 12 0 9 9 7 9 1 9 7 9 7 9 0 1 9 9 13 2
78 9 9 9 10 9 9 0 1 9 10 9 1 9 13 2 7 9 0 7 0 9 9 7 9 9 9 1 9 10 9 13 7 16 9 9 9 9 13 2 1 0 9 1 9 7 9 0 2 9 9 13 2 7 9 9 16 1 9 10 9 9 13 2 1 9 9 0 9 1 9 10 9 9 9 1 9 13 2
31 9 9 9 1 9 13 2 1 9 9 9 0 10 9 9 0 13 2 7 1 9 2 16 9 13 2 1 9 9 13 2
11 1 9 12 9 0 1 10 9 9 13 2
46 9 7 9 12 7 12 9 12 9 1 12 7 12 9 12 7 12 7 12 9 12 1 9 0 9 9 0 1 9 9 0 9 0 9 13 7 9 9 0 1 10 9 9 13 13 2
16 9 0 9 0 9 9 9 2 9 1 3 1 9 9 13 2
19 1 10 9 1 9 12 9 1 9 9 7 12 9 1 9 9 9 13 2
37 9 1 9 0 9 1 9 9 9 12 9 16 1 9 9 0 0 2 0 2 0 2 0 1 9 9 0 0 1 10 9 0 13 2 9 13 2
23 10 9 1 9 12 9 1 12 9 9 0 13 16 12 9 15 9 7 12 9 9 13 2
22 9 9 12 9 1 12 9 2 1 9 9 2 0 1 12 9 1 9 9 0 13 2
27 1 10 9 1 9 3 12 9 0 1 12 9 1 9 1 12 9 1 9 7 9 0 1 9 4 13 2
17 9 9 12 9 1 9 9 9 1 9 1 9 9 9 4 13 2
7 12 9 1 9 0 13 2
33 12 9 0 9 9 1 9 12 9 0 2 16 3 1 9 9 12 9 9 0 9 0 9 1 9 2 0 13 2 3 13 13 2
52 9 9 9 9 9 9 9 9 9 1 9 1 12 1 9 9 9 9 13 2 9 9 0 2 12 0 7 12 9 0 16 9 15 0 13 9 9 1 9 9 1 9 15 1 9 12 9 9 0 0 13 2
34 16 3 1 15 9 13 13 16 9 1 10 9 0 13 2 7 9 0 9 7 9 1 9 0 9 9 9 14 1 9 0 13 13 2
34 10 9 0 16 9 9 13 9 13 16 9 0 9 0 9 0 3 9 7 7 9 9 0 9 0 1 9 9 0 9 7 9 13 2
33 9 0 9 3 9 13 16 1 9 12 1 3 3 12 9 1 9 9 16 1 9 0 9 13 13 2 9 15 14 1 9 13 2
10 9 9 2 9 0 9 0 14 13 2
31 9 0 9 9 13 2 1 3 9 0 12 9 1 9 9 1 9 9 0 1 9 0 1 9 9 15 14 1 9 13 2
53 1 9 9 9 9 9 9 10 9 3 0 16 3 1 9 0 0 13 7 1 9 16 1 9 0 13 2 1 9 1 9 9 15 9 13 2 9 12 9 0 1 9 0 13 7 12 9 14 1 9 9 13 2
50 1 1 10 9 12 9 1 9 0 9 0 9 1 9 0 0 13 7 12 9 1 12 9 9 9 0 1 9 0 9 13 1 9 7 1 9 12 3 1 12 2 12 9 9 1 9 0 9 13 2
26 9 9 1 9 0 7 0 9 9 13 9 9 0 1 9 0 9 1 9 9 9 9 9 13 13 2
26 9 0 7 0 9 9 13 13 12 9 1 9 12 1 12 1 9 9 9 9 15 14 1 9 13 2
42 1 9 1 15 7 1 9 1 9 9 2 9 0 1 9 0 9 13 7 12 9 9 9 1 9 9 0 9 13 2 9 9 9 1 9 9 0 0 3 9 13 2
36 1 9 7 9 9 1 9 0 1 9 9 13 2 0 13 9 9 9 1 9 0 7 0 9 2 3 1 9 0 9 9 9 0 9 13 2
8 0 9 9 1 9 0 13 2
17 9 0 7 9 9 13 0 9 9 0 1 9 9 14 0 13 2
17 9 10 9 1 12 9 9 0 13 16 1 9 9 0 13 13 2
35 9 9 9 2 9 9 12 9 12 9 14 1 9 9 12 9 9 2 1 9 9 2 9 9 0 2 9 7 9 2 1 9 9 13 2
23 9 9 2 1 9 9 13 2 10 0 9 9 13 16 9 9 1 3 1 15 13 13 2
22 9 9 9 13 16 9 9 10 9 2 1 9 9 0 9 0 1 9 9 9 13 2
36 9 9 12 0 2 9 10 9 2 1 12 9 9 0 13 16 13 13 3 9 1 1 9 1 10 9 9 1 9 1 9 9 0 13 13 2
15 9 13 16 9 10 9 2 15 14 0 9 9 4 13 2
31 9 9 0 9 1 10 9 1 9 1 9 0 10 9 9 0 14 1 9 16 1 9 9 7 9 9 13 2 9 13 2
12 9 0 0 1 12 9 9 0 9 13 13 2
8 12 9 9 9 14 9 13 2
28 12 9 1 0 12 2 12 7 12 2 12 9 9 1 9 9 0 9 2 9 9 9 9 9 14 9 13 2
17 9 9 9 9 9 9 10 9 14 9 9 1 9 9 9 13 2
9 10 9 9 0 7 0 13 13 2
20 9 9 9 9 13 2 9 9 9 12 9 0 1 1 9 0 9 9 13 2
30 9 9 9 9 9 0 9 1 9 0 9 9 9 13 2 10 9 3 1 9 0 13 7 1 9 9 9 9 13 2
28 15 13 2 9 3 10 9 0 14 1 9 1 9 0 9 13 7 15 14 1 9 1 1 9 0 3 13 2
20 9 9 13 2 9 12 9 0 1 9 1 9 9 1 9 9 1 9 13 2
13 9 9 3 9 0 14 1 1 10 9 0 13 2
18 9 13 9 0 16 1 3 1 9 9 9 13 2 15 9 0 13 2
26 9 0 9 9 1 9 13 2 0 9 1 15 7 1 9 9 9 1 9 9 9 13 9 9 13 2
14 7 9 0 1 10 9 0 2 1 3 0 13 13 2
37 9 9 9 9 9 9 9 7 9 1 9 9 9 0 9 16 1 3 12 9 0 9 1 9 13 2 0 13 16 10 9 9 2 0 4 13 2
61 9 9 13 16 9 1 9 9 2 9 12 9 0 1 9 1 9 9 0 0 13 3 7 1 9 1 9 9 2 3 12 9 0 1 9 0 13 1 9 7 1 9 9 0 12 9 0 1 9 9 13 7 9 9 9 16 1 9 9 13 2
36 9 9 9 9 9 9 9 9 9 1 9 2 13 2 9 16 1 9 0 9 13 2 1 0 9 16 9 13 2 12 12 9 9 9 13 2
30 9 9 16 16 9 9 9 9 7 9 9 9 9 13 2 13 2 9 0 13 16 9 0 2 1 9 9 0 13 2
30 1 9 9 9 2 9 9 1 9 9 16 1 0 9 1 9 0 1 9 12 9 13 2 0 9 1 9 0 13 2
46 1 10 9 13 13 16 1 12 9 0 2 0 1 9 1 9 9 9 1 0 9 9 9 7 7 1 9 9 9 9 13 7 9 9 9 9 1 9 9 9 0 1 9 9 13 2
20 9 12 9 9 9 1 9 2 9 9 1 9 0 14 1 9 0 9 13 2
34 9 1 9 1 9 1 9 7 7 9 1 13 16 9 9 2 0 9 0 9 9 13 7 1 9 9 1 1 9 0 9 9 13 2
24 1 9 9 10 9 2 9 9 9 0 1 9 1 9 9 9 1 9 9 9 16 9 13 2
35 1 10 9 0 13 16 1 9 9 16 10 9 12 9 9 9 13 2 3 1 12 9 9 0 13 16 9 0 1 9 1 9 0 13 2
16 9 9 16 9 1 0 9 9 9 9 7 9 0 9 13 2
31 0 9 9 1 9 9 15 1 9 0 13 7 9 9 1 9 9 1 10 9 0 9 1 0 9 9 7 9 9 13 2
22 9 1 15 9 9 13 1 9 9 1 9 0 2 10 9 1 9 9 0 9 13 2
22 1 12 9 9 1 9 2 9 0 9 9 9 1 9 9 0 7 9 9 9 13 2
18 9 9 0 1 9 2 9 2 9 7 9 0 9 9 16 9 13 2
32 3 1 9 9 9 1 9 0 2 9 12 9 1 9 2 9 0 0 13 16 9 7 9 9 1 9 9 9 15 9 13 2
30 1 9 9 9 2 10 9 14 9 0 9 9 1 12 9 9 2 12 9 0 7 12 9 1 9 9 9 13 13 2
39 1 9 9 9 1 9 9 9 13 13 16 9 12 9 12 0 0 0 13 13 16 3 9 0 7 0 13 2 9 16 1 9 0 7 0 1 9 13 2
22 9 2 9 2 9 7 9 2 12 9 13 16 9 1 15 1 0 9 9 0 13 2
33 1 10 9 1 10 12 9 1 9 9 2 12 9 3 9 1 9 9 0 13 2 10 9 1 9 1 10 12 9 12 9 13 2
36 1 9 10 9 2 9 0 9 9 1 9 9 13 1 9 7 9 1 9 0 9 0 0 1 9 1 9 9 9 9 1 9 0 9 13 2
43 9 2 9 1 9 7 9 9 2 9 9 7 9 3 9 2 9 9 9 1 9 2 9 9 7 9 9 1 9 9 13 16 1 9 1 9 9 1 9 13 13 13 2
25 9 0 9 9 9 7 9 0 9 9 9 9 1 15 7 9 12 9 0 0 0 14 9 13 2
26 1 0 9 9 9 9 9 9 9 2 9 0 9 1 9 0 9 7 9 9 0 0 9 9 13 2
33 1 10 9 1 1 0 9 9 10 12 9 1 15 2 9 9 0 1 1 9 9 0 9 1 15 1 9 9 0 0 9 13 2
33 1 9 0 9 0 9 9 16 7 1 9 0 9 9 0 0 9 0 1 9 9 13 9 9 1 9 9 14 1 9 9 13 2
42 9 13 2 0 9 10 9 1 9 9 9 1 9 1 9 0 9 9 7 9 9 9 4 13 16 1 9 0 1 9 12 1 0 9 1 9 0 0 9 13 13 2
43 10 9 0 13 2 1 9 0 9 9 0 9 9 0 9 9 14 9 13 7 1 9 0 9 9 15 1 9 3 9 1 9 9 0 1 9 0 1 9 0 4 13 2
33 9 9 1 9 9 1 9 9 9 2 9 0 9 14 3 1 9 9 1 9 7 1 9 9 9 1 9 12 2 9 4 13 2
35 1 9 9 9 1 9 2 9 9 9 9 9 9 13 2 9 10 9 0 1 9 0 1 9 9 1 9 7 9 0 9 15 4 13 2
39 10 9 1 9 1 9 9 9 9 9 9 0 9 7 9 9 0 9 9 13 2 9 12 2 12 2 12 7 12 9 1 9 0 1 9 9 4 13 2
47 1 9 10 9 2 9 7 9 1 9 9 0 7 0 12 9 0 9 9 9 1 9 9 9 12 1 9 9 4 13 7 9 9 0 1 9 15 9 0 9 1 12 9 9 12 13 2
30 1 9 10 9 2 9 0 9 9 13 1 9 12 9 9 9 0 7 1 9 0 2 1 1 9 9 9 9 13 2
40 9 10 9 16 1 9 9 7 9 13 13 0 1 12 12 9 7 9 0 15 12 2 12 9 9 0 12 2 12 9 9 7 12 2 12 9 9 4 13 2
21 9 9 10 9 9 1 9 0 9 12 9 0 12 9 7 9 12 12 9 13 2
17 9 9 1 9 9 0 1 9 2 1 9 9 9 9 4 13 2
29 9 9 0 9 16 1 9 9 0 1 12 9 9 9 1 9 9 9 9 13 2 1 0 9 0 9 9 13 2
34 9 9 9 9 9 9 13 16 9 2 3 12 2 12 9 9 9 0 13 16 1 1 9 3 1 15 2 12 9 9 0 13 13 2
36 9 0 13 2 9 9 7 9 9 1 9 9 9 1 9 0 16 1 9 1 3 9 9 9 9 13 2 1 9 0 9 9 0 9 13 2
24 9 0 9 1 9 0 0 9 0 0 2 9 2 9 7 9 9 0 1 9 0 9 13 2
38 0 9 9 13 16 9 1 9 12 2 12 9 9 7 9 1 12 2 12 9 9 3 1 9 1 9 0 7 0 9 9 1 9 9 0 9 13 2
30 9 1 12 2 12 9 9 2 9 0 1 12 2 12 9 9 7 9 1 12 2 12 9 9 1 9 0 9 13 2
14 9 0 16 0 1 12 9 13 2 9 0 14 13 2
9 9 7 9 9 9 14 9 13 2
23 9 0 16 1 1 9 1 15 0 13 0 1 15 1 9 9 9 1 9 0 9 13 2
41 9 9 0 9 1 9 2 9 1 9 12 1 12 0 0 14 1 9 12 9 1 9 9 13 7 3 1 10 9 12 0 10 9 9 15 14 1 9 13 13 2
15 12 9 9 9 7 9 15 0 1 9 0 7 0 13 2
23 9 9 9 13 16 9 7 9 9 16 0 7 0 13 9 12 9 0 1 9 0 13 2
13 16 1 9 0 12 2 12 9 9 9 0 13 2
15 9 12 9 9 13 16 9 0 9 9 7 9 0 13 2
27 1 9 9 9 9 2 1 10 9 1 12 9 0 10 9 1 9 9 9 9 9 1 10 9 9 13 2
21 1 1 9 9 9 7 9 9 10 9 1 9 12 1 12 12 9 0 9 13 2
45 1 10 12 9 2 12 9 9 13 16 9 9 1 9 9 7 9 1 9 4 1 15 9 13 2 7 9 0 1 15 1 9 9 9 9 9 2 9 7 9 1 9 9 13 2
34 12 9 9 9 9 13 2 9 4 1 9 7 9 0 9 13 2 0 9 3 9 13 16 9 13 9 13 16 9 9 1 9 13 2
28 10 9 0 13 16 1 9 9 7 9 0 1 9 9 9 1 9 2 9 1 9 7 15 15 9 13 13 2
26 12 1 9 16 1 12 1 9 0 9 9 9 9 13 2 13 2 10 9 15 1 9 9 9 13 2
19 3 1 9 9 9 13 7 15 13 10 9 9 0 14 1 9 9 13 2
23 12 9 0 9 0 13 13 16 13 9 9 14 1 9 12 9 1 9 0 0 9 13 2
27 9 1 10 9 0 13 13 16 1 9 0 9 13 7 3 9 13 7 9 0 16 13 15 14 0 13 2
11 10 9 3 1 9 0 9 9 13 13 2
23 9 9 1 9 3 9 13 9 9 7 9 0 7 9 10 9 14 1 9 0 9 13 2
22 10 9 3 9 9 9 1 9 0 1 9 15 13 9 15 14 1 9 0 9 13 2
25 9 0 9 9 0 9 1 10 9 3 0 13 7 9 9 10 9 9 0 1 15 12 9 13 2
22 9 9 9 0 9 9 3 1 9 9 1 9 9 9 2 13 9 9 9 9 13 2
43 1 9 9 1 9 2 9 9 1 9 1 9 9 9 9 9 9 2 1 9 9 9 15 13 2 1 9 9 1 9 9 2 9 9 0 14 1 9 0 9 13 13 2
26 1 9 9 9 9 13 16 1 1 9 9 9 0 2 9 9 9 9 9 9 9 16 9 13 13 2
30 10 9 3 1 10 9 13 16 9 9 9 3 1 9 9 1 9 9 9 13 9 9 14 1 9 9 9 9 13 2
29 12 9 0 9 9 13 2 9 0 0 9 9 9 3 1 12 9 0 1 9 9 15 1 9 0 9 4 13 2
55 10 9 14 9 9 9 9 1 9 9 2 9 7 9 2 9 9 1 9 0 15 1 9 9 9 9 9 9 1 9 9 9 16 1 15 13 13 2 9 0 9 9 9 9 1 3 9 9 4 13 2 9 13 13 2
10 9 7 9 0 9 1 9 9 13 2
13 9 9 15 14 1 9 9 9 13 7 0 13 2
12 1 9 16 15 15 14 3 13 7 9 13 2
24 7 9 0 13 16 1 9 7 9 9 9 14 1 1 15 0 13 7 15 14 1 9 13 2
29 3 1 9 9 13 7 1 15 9 13 7 9 13 16 9 9 1 15 13 2 16 1 3 9 1 9 15 13 2
12 3 1 15 3 9 13 7 3 9 0 13 2
32 9 9 13 7 1 9 15 13 2 7 9 1 9 15 0 13 2 7 16 3 1 15 0 13 9 1 9 14 9 9 13 2
23 9 9 14 1 15 13 7 15 15 1 9 9 1 1 15 9 1 9 13 7 9 13 2
16 3 1 9 1 9 13 7 9 13 16 9 14 1 9 13 2
8 9 16 10 13 1 9 13 2
57 9 9 13 2 3 2 16 9 0 14 1 9 13 7 1 9 9 0 9 13 7 1 10 9 15 14 9 9 7 9 9 13 2 1 9 7 4 10 9 0 7 0 14 3 9 9 16 1 9 3 13 2 1 15 3 13 2
27 7 9 16 7 13 16 4 9 9 14 9 13 2 3 13 2 9 1 10 9 1 15 3 9 13 13 2
35 13 10 9 13 1 15 9 13 2 16 3 9 9 7 9 9 1 1 9 9 7 9 13 7 3 15 16 1 9 9 1 9 13 13 2
18 1 9 15 0 13 2 16 15 1 9 10 9 1 10 9 13 13 2
21 1 10 9 13 2 16 9 15 9 15 14 1 9 13 7 1 15 9 13 13 2
9 13 16 9 0 15 14 13 13 2
16 15 9 9 7 9 13 16 3 1 9 13 7 3 9 13 2
23 9 15 13 16 3 9 13 7 0 13 2 7 9 7 9 15 1 9 13 7 0 13 2
54 1 9 13 16 13 16 1 15 9 1 10 9 9 0 16 9 1 9 9 0 13 9 0 13 2 7 9 10 9 16 9 1 1 9 9 13 7 9 15 14 0 13 2 3 1 9 0 1 9 9 9 9 13 2
11 9 0 1 9 0 1 9 9 0 13 2
17 9 13 1 9 7 9 1 9 0 1 9 7 9 9 9 13 2
18 7 1 1 9 0 9 9 7 9 9 2 0 1 9 0 0 13 2
51 1 9 9 9 1 9 2 9 9 0 9 13 2 9 1 9 0 7 9 1 9 0 1 9 13 13 2 7 10 0 9 13 16 9 13 9 7 9 0 1 9 0 1 9 0 0 1 9 0 13 2
27 9 10 9 1 9 9 9 9 1 12 9 7 12 9 1 9 13 13 2 1 12 9 0 9 13 13 2
28 9 1 10 9 1 9 9 9 1 9 12 1 12 2 0 1 9 0 13 7 1 9 9 1 9 9 13 2
37 10 9 1 13 9 0 12 9 0 1 9 0 1 9 9 9 0 7 10 9 0 9 13 7 9 9 7 9 0 1 9 0 1 15 0 13 2
36 9 0 1 9 1 9 0 2 12 9 0 1 9 9 1 9 0 7 12 2 12 9 0 1 9 9 9 7 9 0 1 9 0 9 13 2
11 9 1 9 9 0 9 1 9 0 13 2
40 9 0 1 9 7 9 0 3 1 0 9 0 13 1 9 10 9 16 9 0 0 9 13 0 13 2 9 9 9 9 7 9 0 9 16 1 15 0 13 2
28 9 9 1 9 15 13 13 2 9 9 9 9 9 9 9 1 9 0 1 9 12 1 12 0 9 4 13 2
39 9 9 9 9 2 12 9 13 16 3 1 9 0 7 0 9 9 13 2 3 7 9 0 1 9 10 9 3 1 9 0 2 3 9 0 1 9 13 2
26 9 1 9 9 9 13 2 9 0 16 0 1 9 9 7 9 13 2 1 9 9 9 0 0 13 2
42 1 9 9 9 1 9 2 9 1 9 9 9 9 9 13 9 16 0 9 9 7 9 1 9 9 9 7 9 13 2 12 9 0 1 15 1 9 9 0 9 13 2
33 10 1 9 13 16 1 9 9 9 9 9 0 1 9 0 16 9 9 9 15 0 1 12 9 13 2 1 12 9 16 0 13 2
20 9 9 9 9 7 9 9 9 9 9 9 1 9 9 10 9 14 0 13 2
22 9 9 7 9 9 0 9 1 9 9 14 16 9 1 15 9 13 13 2 0 13 2
13 9 10 9 0 9 9 9 7 0 9 9 13 2
28 10 9 1 9 9 9 1 12 9 13 16 3 9 9 0 3 9 9 2 9 9 0 2 7 9 9 13 2
17 9 13 9 12 9 1 9 0 1 9 1 3 9 0 9 13 2
43 9 1 9 9 13 3 1 0 9 2 9 9 7 9 15 14 9 13 7 9 9 14 16 0 9 9 7 9 13 7 1 9 0 9 1 9 13 2 1 9 9 13 2
27 9 9 13 9 0 9 9 9 1 12 9 0 13 7 9 9 0 0 1 1 9 9 0 14 9 13 2
34 9 16 1 9 9 1 9 9 9 13 9 13 16 9 3 9 9 14 16 9 0 1 9 9 9 13 1 9 0 9 1 1 13 2
18 12 1 9 13 2 15 9 13 16 9 9 1 10 9 1 1 13 2
7 15 9 3 0 9 13 2
35 1 10 9 0 13 16 3 9 0 13 9 0 3 9 14 16 9 9 2 9 2 9 7 9 9 9 9 13 2 1 9 1 9 13 2
40 10 9 9 0 1 9 9 1 9 9 9 14 1 9 9 13 16 16 1 9 7 7 1 9 9 13 7 9 1 9 9 0 7 10 9 0 1 9 13 2
44 3 1 15 7 9 9 12 9 1 9 9 9 13 16 9 15 12 9 9 9 9 1 9 3 0 3 9 7 9 13 2 9 9 9 1 9 9 9 15 12 9 9 13 2
19 3 1 9 12 9 9 1 9 3 12 0 9 9 9 0 9 13 13 2
39 16 9 9 1 10 9 12 9 9 13 16 1 0 9 0 13 1 15 9 13 7 9 3 13 16 9 3 1 9 12 9 1 9 1 10 9 9 13 2
10 1 9 0 10 9 1 9 0 13 2
15 9 9 1 3 9 7 9 9 1 0 9 15 9 13 2
40 1 9 9 0 9 9 1 9 12 15 13 16 9 15 9 1 15 9 13 2 10 9 1 9 7 9 13 2 4 12 9 0 16 9 9 9 14 9 13 2
10 9 9 15 0 13 7 9 15 0 2
33 10 9 1 9 9 2 13 3 1 9 7 9 1 9 13 2 16 7 0 2 9 9 7 9 7 9 7 9 9 7 9 13 2
16 9 9 9 2 9 2 1 9 9 0 7 1 9 0 13 2
8 9 15 14 1 10 9 13 2
10 3 9 13 2 9 2 9 2 9 2
5 15 9 9 13 2
14 3 9 1 9 15 13 7 13 2 15 9 0 13 2
16 16 10 9 14 1 15 13 1 9 0 9 9 0 1 13 2
11 3 16 9 3 9 15 14 9 15 13 2
10 15 9 13 4 9 15 14 9 13 2
17 12 1 9 0 1 9 9 1 9 1 9 10 9 14 9 13 2
15 9 16 9 0 1 9 9 13 13 2 12 9 9 13 2
21 0 13 13 16 9 9 9 9 13 7 3 9 12 12 9 9 1 9 9 13 2
11 1 10 9 12 12 9 14 9 9 13 2
11 15 9 12 9 3 10 9 14 9 13 2
30 0 13 13 16 1 9 1 9 12 9 2 9 12 9 9 1 9 13 7 1 10 15 9 3 4 12 9 9 13 2
5 16 13 16 2 2
11 9 0 9 12 1 9 9 0 13 13 2
21 10 9 14 9 9 9 1 9 9 9 15 9 2 1 9 12 3 1 9 13 2
19 9 9 9 1 9 9 9 13 2 7 3 1 10 9 9 9 13 13 2
26 1 9 7 1 9 13 13 2 10 9 12 9 13 7 1 10 9 9 0 7 9 0 13 13 13 2
9 9 13 2 12 13 2 12 13 2
17 9 9 9 15 13 1 9 13 7 3 9 15 13 7 9 13 2
6 10 9 16 9 13 2
18 9 15 13 1 9 13 7 15 15 1 9 9 9 7 9 0 13 2
9 9 9 9 13 16 9 9 13 2
11 15 13 7 9 9 15 1 12 9 13 2
4 7 15 13 2
15 9 9 7 9 7 9 9 12 9 1 9 15 3 13 2
4 0 9 13 2
15 9 9 10 9 1 9 9 13 7 1 9 0 0 13 2
7 9 7 9 15 0 13 2
18 3 9 1 10 9 9 9 14 13 13 16 10 9 0 7 0 13 2
24 9 13 2 15 12 9 9 0 7 0 13 7 4 3 12 9 2 0 7 0 7 0 13 2
23 15 16 4 3 9 9 9 9 13 2 9 13 2 9 13 7 10 9 7 10 9 13 2
11 0 13 16 9 15 0 7 0 9 13 2
11 15 4 9 13 3 15 0 7 0 13 2
10 9 9 13 2 9 16 1 9 13 2
5 9 1 9 13 2
12 9 15 1 9 1 9 2 0 7 0 13 2
7 9 15 13 3 15 13 2
12 9 15 13 1 9 13 7 1 0 9 13 2
4 1 9 13 2
5 9 3 9 13 2
16 9 9 13 16 3 9 1 9 1 9 2 1 9 13 13 2
27 9 9 13 16 9 7 9 12 9 1 9 9 9 9 13 13 7 1 1 9 2 0 7 0 9 13 2
17 9 9 9 9 15 14 13 7 13 2 9 15 13 9 14 13 2
9 9 15 13 9 9 14 9 13 2
15 9 15 13 9 9 14 1 9 13 2 13 1 9 13 2
6 9 1 15 9 13 2
3 9 13 2
3 9 13 2
3 9 13 2
30 15 0 9 9 9 1 9 13 7 15 13 9 15 13 16 9 9 14 1 7 13 7 12 9 0 15 1 9 13 2
18 9 0 16 9 0 1 9 9 13 13 2 9 2 0 7 0 13 2
4 15 9 13 2
11 9 13 7 3 0 10 15 14 0 13 2
26 4 15 1 7 1 9 13 16 9 9 9 15 14 13 16 1 9 1 9 13 15 1 15 9 13 2
19 15 9 13 3 10 9 0 1 9 15 9 13 7 9 1 9 9 13 2
12 9 9 16 9 9 0 14 13 3 0 13 2
28 9 9 9 13 7 9 1 1 9 9 2 9 0 1 9 9 9 13 7 13 2 10 9 12 9 9 13 2
8 16 9 9 15 13 2 13 2
7 1 10 9 3 9 13 2
13 16 10 9 0 13 3 9 13 1 15 9 13 2
11 9 13 2 9 13 1 9 0 9 13 2
15 9 15 13 16 1 9 0 9 9 13 9 3 9 13 2
20 9 13 2 9 0 7 0 13 7 15 9 13 2 16 9 13 1 15 13 2
16 9 9 10 9 9 7 9 14 1 9 13 7 0 9 13 2
13 9 7 9 1 0 9 9 15 13 7 0 13 2
12 9 3 9 0 16 9 9 13 9 9 13 2
16 9 9 9 7 9 15 14 13 7 1 12 9 1 9 13 2
4 9 9 13 2
7 9 15 3 9 14 13 2
3 9 13 2
6 9 1 9 9 13 2
12 3 0 13 7 1 1 9 9 15 14 13 2
12 9 15 13 1 9 13 7 9 9 14 13 2
19 9 9 9 14 1 9 9 13 7 13 16 15 9 0 7 1 9 13 2
7 3 9 9 9 9 13 2
17 15 1 1 9 13 13 7 9 9 15 14 0 1 9 13 13 2
11 9 1 9 15 13 7 9 3 0 13 2
10 9 9 1 3 9 0 9 14 13 2
9 3 9 0 1 9 9 9 13 2
16 9 9 15 14 0 13 7 1 9 0 9 9 1 9 13 2
8 9 9 3 1 9 0 13 2
3 9 13 2
10 9 0 7 0 1 9 9 9 13 2
22 9 9 1 9 7 9 15 0 13 1 1 9 9 13 7 1 9 0 1 9 13 2
9 9 1 9 9 13 7 9 13 2
9 15 15 14 9 13 7 3 13 2
15 9 9 1 9 9 9 13 7 9 13 7 1 9 13 2
11 10 9 9 13 16 10 9 9 0 13 2
15 10 9 12 9 9 1 9 7 9 7 9 1 9 13 2
16 9 9 3 1 9 9 13 7 9 9 15 14 3 9 13 2
11 9 3 0 9 14 1 9 9 3 13 2
18 9 7 9 1 9 9 9 13 16 10 9 13 1 9 9 9 13 2
8 12 9 9 13 7 9 13 2
9 9 3 0 1 10 9 9 13 2
14 9 7 9 1 0 9 0 1 9 0 9 0 13 2
23 15 1 9 9 0 9 1 9 9 14 1 9 15 13 16 9 0 14 1 1 15 13 2
9 9 3 1 9 9 9 9 13 2
13 3 9 0 9 13 7 13 2 15 15 14 13 2
17 9 9 9 14 9 13 7 13 10 9 1 9 7 9 15 13 2
13 9 9 13 2 15 15 14 13 2 9 15 13 2
12 9 1 9 15 9 9 14 13 7 9 13 2
11 3 9 2 3 9 1 1 10 9 13 2
17 9 1 1 9 7 9 9 9 13 7 1 9 1 9 9 13 2
5 9 9 15 13 2
11 7 3 9 9 13 1 9 9 9 13 2
9 10 3 9 14 9 13 0 13 2
5 15 1 9 13 2
6 3 9 9 9 13 2
4 3 0 13 2
8 15 9 9 14 9 13 13 2
12 0 13 7 1 9 1 9 7 9 9 13 2
12 9 9 9 1 9 13 2 9 9 9 13 2
3 0 13 2
20 15 7 9 9 1 9 9 9 13 9 9 3 3 9 13 7 1 9 13 2
8 9 9 13 7 13 3 13 2
6 3 10 9 9 13 2
5 9 9 0 13 2
11 15 14 9 13 7 13 2 15 9 13 2
12 9 13 2 3 15 9 13 7 9 14 13 2
11 9 9 13 2 15 13 16 1 15 13 2
12 9 13 2 16 13 13 2 3 3 9 13 2
10 9 9 13 2 15 3 9 9 13 2
16 9 13 2 3 2 15 9 9 13 7 9 9 14 16 13 2
20 3 15 13 13 2 15 10 9 13 16 9 0 15 14 9 1 9 0 13 2
16 9 9 13 2 15 16 3 1 9 7 9 15 9 0 13 2
11 3 2 15 10 9 13 7 15 14 13 2
16 9 0 9 0 13 7 13 2 15 10 15 14 1 9 13 2
6 15 16 9 9 13 2
6 9 9 13 2 9 2
4 13 9 13 2
15 7 9 9 0 13 16 10 10 9 14 1 15 9 13 2
10 15 13 9 12 1 10 9 9 13 2
6 9 13 2 3 9 2
18 9 9 0 1 9 0 13 7 9 15 14 1 9 9 9 9 13 2
13 9 9 1 9 13 2 9 9 1 15 9 13 2
7 0 13 1 15 9 13 2
10 9 9 13 2 15 1 9 15 13 2
10 9 13 2 15 16 9 13 9 13 2
13 13 16 7 15 10 9 13 15 1 15 9 13 2
12 9 9 9 0 15 14 1 1 9 0 13 2
14 0 9 9 1 9 13 2 9 9 1 15 9 13 2
19 12 9 1 9 15 1 9 15 13 2 9 13 15 15 14 1 15 13 2
19 9 2 9 9 9 9 13 7 13 2 3 3 15 14 1 9 0 13 2
7 9 9 15 14 0 13 2
10 9 9 13 2 1 15 9 13 13 2
12 15 3 12 9 9 13 13 16 1 9 13 2
20 9 9 13 2 9 16 15 9 13 3 9 1 3 9 13 16 9 0 13 2
9 9 16 15 9 13 9 9 13 2
11 15 13 1 9 3 9 0 1 9 13 2
26 9 3 9 13 7 13 2 10 9 3 3 9 1 3 9 13 16 0 13 0 1 9 13 7 3 2
14 1 9 9 1 7 13 2 1 9 2 9 7 9 2
8 1 9 15 9 13 0 13 2
15 16 9 13 9 14 1 9 0 13 7 9 1 9 13 2
13 9 9 1 9 0 13 7 9 13 2 13 13 2
5 13 1 9 13 2
4 9 3 13 2
15 9 1 9 7 9 13 9 13 2 15 1 15 9 13 2
32 9 9 9 0 7 0 15 14 9 13 16 9 9 14 0 13 7 3 9 9 15 1 9 0 1 9 13 7 12 9 13 2
5 9 9 0 13 2
8 9 14 1 9 13 7 13 2
7 3 9 13 1 3 13 2
14 9 1 9 13 16 9 9 9 9 9 14 9 13 2
11 3 9 9 15 13 2 9 13 15 13 2
7 9 9 15 14 0 13 2
8 3 9 9 13 2 3 9 2
11 10 9 0 7 0 1 9 9 9 13 2
9 9 1 9 1 9 9 9 13 2
8 1 9 7 9 16 9 13 2
15 3 9 13 16 1 9 0 1 10 9 1 10 9 13 2
9 9 9 0 15 14 1 3 13 2
12 16 9 0 13 2 9 0 14 3 13 2 2
16 9 12 9 16 3 1 7 0 13 13 2 1 15 9 13 2
22 9 1 0 13 2 15 12 9 13 7 13 9 13 16 3 12 9 16 1 9 13 2
7 0 1 9 13 2 3 2
7 9 1 9 13 2 3 2
4 10 15 13 2
9 9 9 2 3 9 13 9 13 2
17 9 2 15 15 15 16 9 15 0 1 9 13 13 9 13 2 2
7 13 3 9 9 15 13 2
13 3 9 13 2 3 16 9 1 9 15 9 13 2
3 9 13 2
11 1 9 15 13 9 9 7 9 15 13 2
10 9 16 15 13 9 1 13 15 13 2
9 9 9 1 15 9 9 15 13 2
8 10 9 3 9 0 1 9 2
10 12 9 9 13 7 9 9 15 13 2
10 1 9 15 14 9 1 15 9 13 2
10 3 1 15 9 1 15 9 15 13 2
9 9 13 0 2 1 10 9 9 2
5 9 2 3 9 2
7 16 9 1 9 15 13 2
8 1 9 10 9 15 0 13 2
13 16 15 10 9 9 1 1 9 7 9 15 13 2
10 16 0 3 9 1 9 13 10 9 2
11 9 16 9 1 15 2 7 9 15 13 2
30 9 1 9 0 7 0 7 9 0 0 0 9 1 15 7 9 15 2 9 9 1 9 9 12 9 9 9 14 13 2
32 9 9 9 2 9 9 7 9 0 9 9 1 9 12 9 0 0 9 13 7 1 9 9 9 9 2 9 0 15 9 13 2
33 9 9 1 9 13 16 1 9 1 9 9 2 9 0 9 9 1 1 9 7 9 1 9 9 12 9 14 1 9 15 4 13 2
36 9 9 13 2 9 7 9 1 9 9 9 0 2 1 9 9 12 9 9 13 16 13 1 10 9 9 0 9 1 9 7 9 0 9 13 2
33 15 1 1 9 0 9 9 9 0 13 2 9 0 1 9 0 13 7 9 9 0 16 1 12 9 9 9 15 14 9 4 13 2
29 9 9 9 9 9 16 13 2 9 1 9 9 0 3 9 9 0 13 7 9 15 14 1 9 0 15 9 13 2
31 9 9 0 9 0 1 12 7 0 9 9 0 9 0 9 9 13 2 9 9 9 13 7 1 12 2 12 9 13 13 2
46 9 9 9 9 9 1 9 13 2 1 9 9 9 0 9 12 16 1 12 9 9 9 13 13 2 9 9 1 1 9 0 1 12 2 12 9 1 12 2 12 9 9 0 13 13 2
23 9 1 9 0 1 9 15 13 2 9 9 0 7 0 9 1 1 9 12 9 13 13 2
32 15 9 9 9 0 14 12 2 12 9 9 13 7 13 2 9 0 9 9 0 1 9 12 7 12 12 2 12 9 13 13 2
25 9 9 0 9 0 1 1 9 9 13 2 9 9 9 12 7 9 1 12 2 12 9 13 13 2
27 15 9 13 2 16 9 0 3 13 13 7 9 1 9 9 0 13 10 9 9 1 1 12 9 4 13 2
26 9 9 1 9 12 7 12 12 2 12 9 13 13 16 1 9 12 7 12 1 12 2 12 9 13 2
8 6 9 9 7 9 3 13 2
72 9 7 9 0 9 9 16 1 9 9 9 7 9 1 9 9 13 13 2 16 9 1 1 12 9 1 9 9 9 0 9 0 9 3 1 9 9 9 10 9 9 13 7 1 9 10 9 1 9 7 9 9 0 2 9 9 9 0 7 9 7 9 1 1 9 9 9 14 9 13 13 2
69 1 9 7 1 9 9 0 9 9 9 0 9 3 1 9 9 7 9 9 0 10 9 0 13 7 0 13 13 15 1 9 9 9 9 10 9 9 9 9 1 9 9 9 9 13 2 9 9 9 7 1 10 9 1 9 9 0 1 12 9 3 9 9 9 1 10 9 13 2
34 1 9 9 3 9 9 0 0 13 7 3 9 9 9 9 10 3 0 16 4 1 9 9 1 9 16 9 9 14 0 13 0 13 2
37 9 9 9 9 7 9 9 1 10 9 9 7 9 9 7 9 9 9 9 9 1 9 15 9 9 10 9 9 0 1 9 9 14 3 0 13 2
16 1 9 0 9 9 1 9 9 0 1 9 9 9 13 13 2
22 7 1 0 9 10 9 3 1 9 9 7 9 1 9 9 7 9 0 9 13 13 2
39 9 9 0 9 16 16 3 3 1 9 7 9 9 0 10 9 9 13 2 1 0 9 9 15 3 1 9 9 0 1 9 7 9 9 9 9 9 13 2
13 9 9 9 1 9 9 15 9 9 14 0 13 2
43 1 9 1 9 0 9 0 9 7 7 1 9 9 10 9 9 10 9 9 10 9 3 9 13 16 16 9 9 1 9 9 16 3 7 16 3 9 0 1 9 9 13 2
34 16 1 9 15 9 9 7 0 0 7 9 9 0 0 13 1 9 4 1 9 0 10 9 9 7 9 0 7 7 0 14 9 13 2
29 16 9 9 9 9 9 1 9 1 9 9 9 1 9 9 2 3 1 9 9 7 9 0 1 9 9 9 13 2
31 9 9 0 13 7 1 9 9 16 3 9 0 1 9 1 9 9 4 13 7 3 1 9 9 1 1 9 0 4 13 2
29 0 9 10 9 9 9 9 9 7 9 1 9 0 9 7 1 1 9 9 7 9 10 9 0 1 9 0 13 2
15 9 0 7 0 9 0 9 4 1 10 9 0 9 13 2
26 9 12 12 9 0 9 13 16 4 1 9 7 1 9 9 7 9 9 0 7 0 1 15 9 13 2
35 9 0 9 9 0 9 1 9 9 9 9 14 1 10 9 9 13 1 9 10 9 1 9 1 9 0 7 9 7 9 9 9 4 13 2
5 9 0 0 13 2
74 9 9 1 9 0 15 2 9 7 9 0 2 13 13 2 9 9 13 16 1 9 3 1 9 0 7 0 3 1 9 13 7 9 1 15 15 13 16 9 1 9 1 9 12 9 7 9 1 9 15 0 13 7 1 9 9 1 3 7 9 9 1 9 10 9 0 15 14 1 9 0 3 13 2
16 7 10 9 1 9 9 9 9 0 9 1 0 0 0 13 2
35 1 12 9 0 1 9 15 2 10 9 1 1 9 0 0 9 0 16 13 16 1 9 9 1 9 9 3 9 0 14 1 1 4 13 2
43 9 1 10 9 9 13 16 3 1 9 9 7 9 9 1 12 9 0 13 13 7 9 3 0 13 1 15 10 9 13 7 9 15 9 1 9 9 0 7 9 0 13 2
55 10 9 1 9 9 1 9 0 9 13 1 9 9 0 12 9 2 1 15 7 9 14 1 9 13 2 3 1 1 9 7 9 9 9 2 9 9 15 14 9 13 7 1 9 9 7 9 0 14 16 1 9 9 13 2
43 1 9 7 9 9 9 0 14 1 9 9 9 16 9 1 9 0 13 2 1 9 13 1 3 16 9 0 1 9 9 10 9 7 9 14 1 9 13 13 9 0 13 2
39 3 3 0 13 16 9 0 1 9 9 1 9 0 13 7 9 13 16 1 9 9 9 9 12 9 1 9 1 9 9 9 7 9 0 1 15 9 13 2
14 16 0 13 16 1 9 9 13 7 9 13 9 13 2
43 1 10 9 10 9 16 1 9 1 9 13 9 0 9 1 9 9 9 9 14 1 12 9 7 9 14 1 9 0 13 2 3 0 7 0 1 1 9 9 0 9 13 2
42 9 1 9 0 9 9 9 9 9 9 14 1 9 1 9 0 9 13 7 13 13 2 9 9 0 9 0 1 9 9 9 9 0 1 9 0 9 0 9 13 13 2
28 9 9 9 0 13 2 9 9 9 2 9 0 9 2 9 9 1 9 0 9 9 2 9 9 2 9 13 2
39 9 9 9 13 16 9 0 9 0 1 9 0 0 13 7 1 10 9 1 9 0 16 9 13 16 10 9 9 12 9 1 9 9 1 9 14 3 13 2
7 15 13 2 9 9 13 2
6 9 1 9 9 13 2
9 9 1 9 9 15 4 3 9 2
43 9 0 13 16 2 1 9 13 15 9 13 1 10 9 2 9 9 14 16 3 1 1 9 9 9 13 2 0 13 2 9 16 9 9 14 1 1 9 0 9 13 13 2
23 1 9 9 9 2 9 9 1 9 0 0 13 16 10 9 0 14 1 9 9 9 13 2
26 15 13 2 1 9 16 15 0 13 7 10 9 14 13 2 1 15 9 4 13 1 9 9 9 13 2
16 9 3 0 13 9 9 13 7 13 10 9 0 14 0 13 2
25 1 9 9 9 15 1 9 0 7 9 0 13 16 9 9 0 1 9 12 9 1 9 0 13 2
23 1 9 9 9 1 9 0 2 10 9 9 13 1 9 9 9 1 9 0 9 9 13 2
21 9 13 3 16 9 0 9 9 0 0 13 2 3 10 9 9 9 0 4 13 2
35 1 10 9 9 9 9 9 16 9 0 13 2 9 9 9 9 9 0 1 9 9 15 1 9 0 9 2 9 9 0 9 14 9 13 2
45 10 9 9 13 16 2 9 9 1 9 9 9 15 1 9 7 9 13 16 1 15 0 13 7 13 2 10 10 12 9 3 7 1 9 0 9 0 13 13 9 1 9 9 13 2
31 1 10 9 9 9 9 9 16 13 16 2 9 9 9 9 0 9 9 9 0 7 9 1 9 0 9 1 9 13 13 2
27 9 9 9 9 9 9 1 9 9 13 2 16 9 9 9 9 0 13 7 9 0 1 9 9 13 13 2
42 1 9 9 2 9 9 1 9 0 2 9 13 1 9 2 7 9 9 9 1 10 9 16 9 0 0 1 9 9 13 3 9 1 9 7 9 1 1 9 9 13 2
66 9 9 9 0 13 2 9 9 9 9 13 16 9 9 9 4 1 9 1 10 9 0 3 13 7 1 3 7 15 1 9 1 1 9 9 9 16 9 1 15 9 13 1 0 9 9 9 9 13 1 9 13 16 10 9 9 9 1 9 9 1 9 0 0 13 2
41 9 9 16 1 10 9 9 13 16 2 9 9 9 2 9 0 9 9 9 1 9 0 1 9 9 2 9 2 9 9 1 9 0 1 9 9 1 10 9 13 2
62 9 9 1 9 15 2 9 9 1 9 9 2 13 13 2 1 9 0 2 7 3 1 9 12 9 1 9 2 15 3 1 9 0 1 9 7 9 13 1 9 7 9 0 13 1 9 15 1 9 7 9 2 7 1 9 7 9 1 9 7 9 2
20 15 1 0 9 9 0 7 0 9 13 16 4 9 15 14 1 1 0 13 2
20 1 9 15 2 10 15 16 1 9 9 7 9 9 0 4 1 9 9 13 2
28 9 9 0 7 0 7 0 1 10 9 2 9 7 9 0 14 1 15 1 9 13 7 15 14 1 9 13 2
32 1 9 16 9 1 9 7 9 7 9 13 2 4 9 13 16 16 9 9 0 7 9 9 13 7 7 9 1 9 13 13 2
19 16 9 0 13 13 7 7 9 10 9 1 9 9 7 9 9 9 13 2
35 9 2 9 9 0 7 0 13 16 9 14 1 9 3 13 7 1 1 15 2 0 9 9 7 9 14 13 7 3 9 0 1 15 14 2
13 15 15 1 9 7 9 9 0 9 16 9 13 2
30 0 13 9 0 16 16 1 9 9 0 9 9 13 2 9 9 0 15 7 9 7 9 9 0 14 9 9 13 13 2
25 9 9 3 1 9 0 7 0 0 13 16 0 9 7 0 9 15 2 3 0 13 7 3 0 2
22 10 9 16 3 9 15 14 1 1 9 0 2 7 7 9 9 2 0 7 0 13 2
29 10 9 1 9 0 9 15 3 13 16 9 0 7 9 0 0 10 9 14 9 9 9 13 16 9 0 9 13 2
25 1 10 9 16 10 9 7 9 0 0 9 9 15 13 2 9 7 9 16 9 15 14 9 13 2
24 9 15 9 7 9 0 13 16 3 3 1 9 13 7 3 9 15 14 1 9 10 9 13 2
18 9 16 9 0 15 7 9 0 9 9 13 2 1 15 3 0 13 2
58 1 10 9 7 9 9 14 1 9 0 16 1 9 9 0 7 0 15 9 13 2 1 9 13 7 1 9 1 9 0 0 7 9 16 1 15 9 13 7 9 13 2 9 7 9 0 7 0 15 15 14 9 9 7 3 9 13 2
17 9 15 1 10 9 0 1 10 9 7 9 7 9 3 0 13 2
14 10 9 13 16 13 7 4 1 9 9 0 0 13 2
64 1 9 1 9 0 9 0 9 1 9 9 9 1 1 9 9 0 16 9 9 0 1 9 9 7 9 0 9 1 9 10 9 2 4 9 9 1 9 7 9 0 1 10 9 14 13 16 1 9 0 9 15 14 1 9 0 0 13 7 1 15 9 13 2
16 10 9 16 1 9 0 7 7 1 9 0 0 9 0 13 2
43 16 1 10 9 2 9 1 9 1 9 1 9 9 9 0 1 1 9 13 2 1 9 16 3 1 9 13 2 15 13 16 4 0 0 13 9 2 9 0 13 7 0 2
23 16 1 10 9 13 16 9 0 13 2 3 3 9 9 13 2 9 1 15 14 9 13 2
18 16 3 13 3 9 0 15 14 1 1 10 9 0 7 0 9 13 2
33 16 15 9 0 7 3 0 1 9 0 9 3 9 9 1 10 9 13 16 9 1 1 9 13 7 1 10 9 9 9 14 13 2
27 7 7 1 15 7 9 0 15 3 9 0 15 14 13 7 1 9 10 9 9 3 1 10 9 0 13 2
3 9 13 2
17 16 3 2 3 9 7 3 9 3 13 7 1 10 9 9 13 2
49 16 9 15 13 13 16 9 0 0 2 9 1 9 0 15 9 13 7 9 9 15 2 3 13 3 15 7 3 1 15 9 7 9 0 15 1 9 9 13 7 1 9 0 7 0 0 9 13 2
49 9 13 10 9 7 9 9 1 15 9 13 7 1 15 13 16 3 13 1 9 9 0 2 1 9 0 9 7 9 13 16 15 1 15 3 1 9 15 1 9 2 9 7 3 9 9 9 13 2
22 7 1 3 9 0 7 0 13 9 9 7 9 9 7 9 9 7 9 14 1 13 2
24 3 3 9 0 7 9 9 13 13 7 1 9 9 0 0 9 13 9 0 15 14 9 13 2
20 9 0 16 9 9 2 3 1 15 9 13 2 3 3 0 1 10 9 13 2
33 3 1 9 9 9 2 9 1 9 7 9 0 1 9 13 16 1 9 0 2 3 9 9 9 7 9 9 9 7 9 4 13 2
23 9 7 9 0 16 3 13 3 3 0 1 9 9 2 10 9 16 1 9 9 9 13 2
32 1 9 9 2 0 13 9 13 16 9 2 9 7 9 7 9 15 14 9 13 7 15 14 1 9 7 9 7 9 9 13 2
4 16 9 13 2
57 9 9 9 9 1 9 1 9 2 16 9 13 3 13 2 1 9 9 13 13 2 12 1 9 9 9 1 1 9 15 2 1 9 13 13 2 1 9 9 12 9 9 9 13 16 3 13 7 1 9 0 9 13 16 3 13 2
47 9 10 9 15 13 16 9 9 1 9 3 1 10 9 9 9 9 14 13 7 1 15 9 13 16 9 9 1 9 9 0 13 2 9 16 0 13 7 10 9 0 9 14 1 9 13 2
37 7 9 13 10 9 9 16 9 13 1 9 9 9 1 9 9 13 3 9 13 7 3 3 1 12 7 12 9 13 13 16 15 3 9 9 13 2
69 16 10 9 14 1 1 9 9 7 9 10 9 7 9 15 9 13 7 1 9 7 9 7 9 9 9 9 9 16 9 13 2 3 4 13 9 15 13 13 16 9 1 9 9 0 13 7 3 13 3 13 7 3 9 9 3 0 7 9 0 1 9 7 9 0 1 9 13 2
43 9 0 9 0 1 9 0 9 9 12 7 0 9 12 7 9 2 1 9 1 10 9 2 9 13 16 9 16 13 16 3 13 7 7 13 16 3 13 7 3 16 13 2
39 9 13 9 1 10 9 9 13 7 1 15 13 16 3 9 9 1 9 0 16 9 0 1 9 1 15 1 9 9 9 12 9 13 3 13 16 3 13 2
63 16 9 9 9 14 13 7 13 16 15 1 9 12 9 7 12 9 0 9 9 13 7 9 1 9 9 13 13 7 16 9 1 9 3 1 9 9 0 1 9 15 7 1 9 15 9 7 9 1 9 9 13 13 16 1 9 9 9 0 1 9 13 2
33 1 9 0 9 9 12 7 12 2 16 1 9 12 9 3 1 9 9 2 9 9 1 9 1 9 13 2 9 0 15 3 13 2
19 16 13 16 9 14 0 13 7 1 9 15 3 9 9 14 13 0 13 2
29 7 9 9 13 2 9 0 15 9 12 9 7 9 0 13 2 16 0 9 9 0 9 10 9 0 7 0 13 2
16 1 9 0 4 9 1 9 13 16 1 9 0 9 9 13 2
12 9 3 13 2 9 15 1 9 0 3 13 2
16 15 1 10 9 3 1 9 13 9 9 7 7 9 0 13 2
19 7 9 13 2 10 9 9 1 15 2 9 9 7 9 9 9 9 13 2
44 10 9 2 16 12 1 12 9 9 9 1 10 9 13 2 3 1 9 2 7 1 10 9 9 7 0 13 7 16 4 13 16 9 9 16 9 9 9 14 13 13 3 13 2
49 16 1 9 3 1 9 9 0 1 15 9 7 1 9 1 9 2 1 10 9 2 9 0 9 2 9 9 2 9 2 9 0 13 16 1 10 9 7 0 3 1 9 2 9 9 0 9 13 2
16 16 12 9 1 10 9 9 15 14 1 9 10 9 9 13 2
38 16 4 13 9 13 1 1 3 13 7 0 1 9 13 7 1 9 9 16 13 3 13 2 1 1 9 7 9 7 9 9 9 13 7 1 9 13 2
53 16 15 9 1 9 9 13 16 13 1 9 13 3 13 7 1 10 9 9 13 7 15 15 9 7 9 7 9 7 9 14 9 13 7 3 3 1 12 7 12 9 4 1 9 9 9 9 13 16 3 4 13 2
16 16 1 10 0 9 9 9 15 14 2 9 0 13 7 13 2
17 16 9 1 15 13 0 9 9 7 0 9 9 9 3 0 13 2
35 16 15 9 9 14 1 10 9 0 7 0 7 0 13 16 13 1 9 0 9 13 16 9 9 7 9 0 13 7 1 10 9 9 13 2
112 13 16 1 9 0 9 1 9 7 9 9 9 1 9 0 7 13 13 16 15 1 9 9 9 0 13 7 15 9 16 1 9 0 7 0 15 1 9 2 9 2 9 9 0 2 16 1 1 9 2 9 1 9 2 1 9 2 16 13 16 3 13 7 7 13 16 3 13 7 3 13 16 1 12 9 9 9 2 9 1 9 15 16 9 9 9 13 1 9 9 9 13 13 7 1 9 15 2 16 1 9 9 0 7 0 2 9 7 9 13 13 2
28 3 1 9 0 9 9 9 7 9 9 0 2 3 12 9 12 9 0 7 0 15 13 7 1 7 0 13 2
36 1 9 12 2 12 2 12 9 0 1 9 1 9 9 13 2 3 9 9 9 7 9 9 0 1 9 9 1 9 0 2 3 0 9 13 2
82 7 9 9 1 9 13 2 9 1 9 1 9 9 15 0 13 7 1 3 9 9 0 13 7 3 16 1 9 1 9 9 10 9 9 7 9 7 9 0 15 1 9 0 9 15 7 9 15 14 9 13 7 1 9 15 7 9 0 1 9 9 9 9 13 2 16 0 13 1 9 10 9 1 9 1 12 9 9 0 0 13 2
48 9 1 9 0 13 2 1 15 10 14 9 13 16 13 9 0 0 9 13 2 1 9 7 9 9 0 3 9 16 0 13 7 9 0 0 3 9 0 16 0 13 2 9 1 9 9 13 2
16 16 13 9 9 0 14 16 1 9 13 9 13 16 3 13 2
22 7 9 2 1 9 13 2 3 1 9 10 9 16 9 15 1 9 0 13 13 13 2
14 3 9 1 9 0 9 0 1 9 9 0 13 13 2
18 16 3 9 9 1 9 9 15 4 13 16 9 0 3 9 14 13 2
23 3 9 9 16 1 9 9 0 15 15 7 7 9 9 9 15 1 9 9 9 9 13 2
42 1 9 10 9 9 9 1 9 9 7 9 7 9 9 0 13 2 1 9 0 2 9 9 13 1 9 1 9 2 9 13 7 7 1 9 0 9 1 15 0 13 2
45 4 9 0 14 1 9 7 1 10 9 1 9 9 13 7 3 9 15 13 2 3 4 1 9 0 1 15 9 9 13 2 3 9 9 7 7 9 9 14 1 9 9 4 13 2
10 9 1 9 10 9 7 9 0 13 2
34 10 9 9 7 9 1 9 9 1 9 7 9 9 14 1 9 13 0 13 7 9 1 10 10 9 9 7 9 15 14 9 13 13 2
50 13 16 9 9 2 16 9 9 1 9 3 1 9 2 3 7 15 9 9 9 9 7 9 9 9 0 14 1 9 7 1 1 16 9 13 7 9 9 7 9 7 9 9 0 14 16 9 13 13 2
31 1 9 0 9 16 1 9 9 7 9 7 1 1 9 9 2 1 9 2 9 2 9 9 0 2 9 13 16 3 13 2
47 3 3 3 1 12 7 12 9 15 9 10 9 0 13 7 3 13 9 3 7 3 15 14 16 9 9 0 7 9 1 9 9 7 9 1 9 9 1 9 13 2 1 9 9 9 13 2
63 0 13 16 9 9 9 0 7 9 9 2 3 7 3 1 9 9 9 13 2 7 9 9 1 9 10 9 1 9 1 9 7 9 9 0 15 0 13 13 7 9 9 7 9 7 9 14 1 9 7 9 9 7 9 7 9 9 9 13 7 13 13 2
36 16 1 10 9 0 7 0 9 16 9 7 9 9 15 15 14 1 9 9 9 1 9 13 2 9 9 9 1 9 7 9 7 9 0 13 2
46 1 9 12 9 3 1 9 9 0 10 9 9 1 9 1 9 9 9 1 9 9 9 2 3 9 12 9 14 1 15 13 7 1 1 9 9 7 9 0 9 13 7 1 9 13 2
20 1 9 9 16 16 9 9 1 9 9 7 9 9 13 10 9 1 9 13 2
31 9 12 9 1 9 9 0 16 16 1 9 9 0 9 0 9 13 2 9 9 7 9 0 9 1 9 0 9 9 13 2
60 9 9 9 9 0 9 9 1 9 9 9 1 9 9 1 9 9 9 13 2 9 0 9 9 13 16 9 9 1 9 9 9 9 9 1 12 9 14 9 13 7 15 1 9 0 9 9 0 9 1 1 9 9 1 9 10 9 9 13 2
31 9 9 0 1 13 7 13 1 9 9 0 13 2 15 0 13 10 9 7 9 0 9 13 2 10 9 3 0 9 13 2
18 9 9 1 9 0 9 9 9 9 9 9 7 9 9 0 4 13 2
8 9 9 0 1 12 9 13 2
28 9 0 9 0 0 9 1 9 9 2 9 1 9 7 9 0 9 13 7 10 9 14 1 9 0 4 13 2
39 9 9 1 9 9 9 7 9 9 1 9 9 0 9 9 9 9 13 2 9 0 9 1 9 9 7 9 1 9 0 9 0 7 0 1 15 9 13 2
50 9 9 9 14 0 1 12 9 9 10 9 13 7 13 2 9 0 9 9 9 7 9 1 9 15 9 9 9 9 13 13 16 1 9 9 0 2 0 7 9 0 10 9 1 9 9 0 15 13 2
45 9 1 9 1 15 16 4 1 3 9 9 9 1 10 9 13 13 2 13 2 15 9 9 9 9 4 1 9 0 1 9 0 7 0 15 9 13 7 1 9 9 9 15 13 2
37 9 9 1 9 1 9 9 0 9 0 1 9 9 0 13 2 9 0 9 7 9 1 1 9 9 9 9 7 9 0 9 14 9 1 9 13 2
49 9 1 9 1 15 16 1 9 9 0 1 9 9 0 3 12 9 9 9 1 9 9 13 7 9 1 9 9 13 2 13 2 10 9 9 2 9 7 9 9 0 3 9 0 9 0 9 13 2
32 9 2 9 2 9 7 9 0 14 9 9 12 9 0 13 7 13 2 10 9 1 9 0 1 9 7 9 0 9 9 13 2
24 9 9 3 9 9 13 16 9 9 3 0 9 9 9 14 0 13 16 9 9 0 0 13 2
37 9 9 9 1 9 13 2 9 15 15 13 16 9 1 9 0 1 9 9 16 9 9 2 9 2 9 7 9 9 13 12 1 0 9 13 13 2
52 9 9 1 1 9 9 13 2 10 9 16 15 1 9 0 13 15 13 16 1 10 9 1 9 9 9 1 9 9 13 7 1 9 1 9 16 16 9 7 9 0 13 2 1 9 9 0 1 9 9 13 2
28 15 9 13 2 1 9 0 13 3 0 9 9 1 9 14 9 13 7 3 3 1 9 9 9 1 9 13 2
41 9 9 13 2 9 1 9 9 1 9 0 1 9 9 7 9 9 0 13 16 10 9 7 9 0 16 1 9 9 0 7 9 9 9 9 4 13 2 9 13 2
23 9 9 13 2 4 1 9 0 1 9 10 9 9 13 7 9 7 9 0 16 9 13 2
39 9 9 16 13 2 4 1 9 0 9 13 7 9 0 0 13 7 15 9 1 10 9 9 13 16 1 9 9 9 13 16 9 9 7 9 1 9 13 2
3 9 13 2
38 9 9 1 9 0 9 9 16 1 9 13 2 1 9 15 9 16 9 13 7 9 14 16 9 9 13 9 13 9 13 16 13 15 9 9 0 13 2
48 9 16 9 9 0 14 0 13 9 9 9 14 0 13 3 7 16 0 13 2 13 9 9 13 16 13 3 4 13 7 3 4 13 7 16 9 1 1 9 9 13 9 15 0 13 3 0 2
34 9 9 13 2 16 15 1 9 0 13 9 0 9 1 9 15 13 7 3 15 1 9 2 1 9 0 16 9 1 9 13 9 13 2
31 8 8 3 1 9 13 13 9 15 12 9 13 2 9 9 1 9 9 7 9 9 10 9 16 1 9 7 9 9 13 2
18 3 10 9 9 14 16 9 7 9 13 16 9 1 15 9 13 13 2
34 1 9 0 15 1 9 13 13 2 8 8 8 8 8 8 8 8 8 9 8 8 8 8 8 8 8 8 8 8 8 8 8 8 2
22 1 12 9 9 15 2 9 0 9 9 13 16 9 1 9 7 9 9 9 0 13 2
21 9 16 16 9 9 15 14 1 9 13 1 9 9 15 0 13 16 10 9 13 2
29 9 7 9 7 10 9 9 15 14 1 9 9 13 13 2 3 1 9 2 9 7 9 9 9 10 9 14 13 2
8 9 9 0 9 14 9 13 2
12 1 9 9 12 9 0 1 9 9 9 13 2
24 10 12 9 3 1 9 9 13 7 9 9 2 9 7 9 1 9 1 9 10 9 14 13 2
31 9 9 9 0 7 0 2 9 1 9 9 9 2 9 1 9 9 1 10 9 9 13 16 3 9 15 1 9 9 13 2
38 1 9 9 2 9 9 14 9 9 9 13 7 1 1 9 13 7 9 15 10 9 0 13 16 15 9 9 14 0 13 7 9 14 1 9 13 13 2
15 9 9 13 9 9 14 0 13 7 1 9 1 9 13 2
27 9 16 9 13 9 9 14 1 9 1 9 13 2 16 9 3 9 7 9 1 1 9 14 1 9 13 2
46 9 9 16 9 8 9 1 9 9 2 9 2 7 9 15 1 9 13 2 16 9 9 14 0 13 2 1 9 13 7 0 9 13 2 1 9 9 16 9 13 2 9 10 9 13 2
17 9 13 9 13 9 7 9 14 1 10 9 9 7 9 9 13 2
29 9 16 1 9 9 9 9 0 13 2 1 0 9 2 1 9 0 13 16 9 9 7 9 1 9 15 14 13 2
23 10 9 9 2 1 9 9 9 9 13 2 16 3 13 16 9 9 7 9 9 9 13 2
17 0 13 9 9 7 9 9 15 3 9 7 9 1 9 9 13 2
18 10 9 16 1 9 9 12 9 0 1 9 7 9 0 7 0 13 2
23 16 9 7 9 7 9 16 1 9 9 15 7 1 1 7 1 9 0 13 2 0 13 2
36 9 9 9 2 9 2 1 9 9 9 10 9 13 2 8 8 8 8 8 8 2 8 8 8 8 8 8 8 8 8 8 8 8 8 8 2
27 10 9 0 2 9 1 9 9 1 1 7 1 9 1 9 9 1 9 9 3 9 13 1 9 9 0 2
20 10 9 0 1 3 13 16 9 9 1 1 9 0 3 9 9 13 1 9 2
17 7 10 9 3 7 3 9 9 7 9 7 9 9 14 9 13 2
17 0 13 16 9 0 1 9 7 9 9 9 7 9 14 0 13 2
23 9 9 1 9 9 12 2 16 3 3 1 9 9 9 2 9 2 1 9 9 9 13 2
15 9 9 2 9 2 14 1 9 0 9 9 9 0 13 2
9 9 0 2 9 1 9 9 13 2
27 9 16 1 1 9 9 0 7 0 13 2 3 9 2 3 1 9 9 1 9 12 0 9 0 13 13 2
46 1 10 9 16 1 9 12 9 1 3 2 12 9 0 1 1 9 9 13 2 0 2 9 7 9 9 2 0 2 9 9 9 2 9 2 7 9 7 9 7 9 7 9 8 9 2
15 9 13 9 14 1 9 12 9 0 7 9 0 0 13 2
27 1 15 7 1 9 7 9 7 9 9 3 0 13 2 9 1 10 9 0 13 16 9 3 9 0 13 2
26 1 15 9 3 9 9 7 9 1 15 13 16 1 9 9 0 14 1 15 13 7 9 1 9 13 2
13 9 0 9 2 1 9 0 13 16 3 9 13 2
16 7 9 15 3 9 7 9 7 9 0 15 14 0 13 13 2
18 3 9 9 13 16 9 7 9 9 1 9 9 1 9 0 9 13 2
10 1 9 3 0 9 7 9 9 13 2
11 1 9 9 13 16 15 1 9 9 13 2
18 9 1 9 9 13 16 1 9 9 13 16 9 7 9 15 9 13 2
28 9 14 9 13 7 1 9 9 7 9 1 15 0 9 9 13 7 13 10 9 14 9 13 7 1 9 13 2
9 10 9 9 14 1 9 9 13 2
15 1 12 9 2 9 9 7 9 14 1 9 15 9 13 2
23 0 9 15 1 9 15 13 16 10 9 7 9 15 14 3 7 3 1 9 9 9 13 2
11 13 2 9 0 13 16 9 15 0 13 2
16 15 1 9 10 9 13 9 13 16 9 4 1 15 9 13 2
34 9 9 1 9 15 13 16 9 9 7 9 15 14 9 13 7 9 1 9 1 15 9 13 2 9 9 9 7 9 9 15 13 13 2
17 1 9 9 2 9 13 9 1 9 9 7 9 9 14 9 13 2
5 9 9 9 13 2
15 1 9 1 9 9 9 9 16 3 9 13 13 9 13 2
7 16 1 9 9 9 13 2
6 9 1 9 9 13 2
21 9 1 9 0 7 9 9 2 1 9 0 2 9 9 0 9 7 9 13 13 2
16 0 7 0 1 9 9 13 16 3 1 9 9 15 13 13 2
20 1 15 1 9 9 15 1 9 7 9 1 9 13 13 3 9 7 9 13 2
10 9 9 9 16 3 9 9 15 13 2
14 9 12 7 12 7 12 9 1 9 9 9 9 13 2
13 3 9 13 1 10 9 9 0 1 9 9 13 2
20 1 9 9 16 9 3 13 16 3 9 0 14 1 9 9 9 9 9 13 2
7 1 9 9 9 9 13 2
11 9 9 2 9 2 7 9 1 9 13 2
9 15 14 16 1 9 9 9 13 2
8 9 9 1 9 9 0 13 2
13 9 9 2 9 2 13 13 2 10 3 9 13 2
34 1 9 9 9 1 9 9 9 1 9 2 9 0 9 1 9 1 9 9 1 9 0 0 9 13 16 1 9 10 9 9 9 13 2
41 9 12 9 9 1 9 9 9 9 13 16 9 0 9 1 9 16 1 10 9 9 13 2 9 15 14 1 12 12 9 0 13 16 1 9 9 9 9 9 13 2
65 1 9 9 9 9 2 0 4 12 12 9 1 9 9 13 7 3 12 9 0 13 16 9 15 14 1 9 9 9 9 13 2 9 16 1 9 9 9 9 1 9 9 9 13 3 1 12 9 9 3 9 1 15 1 15 4 13 2 9 16 3 9 15 13 2
40 1 9 9 9 2 9 0 9 9 12 9 9 13 16 1 9 7 9 0 10 9 9 13 7 9 9 9 14 0 13 1 1 9 9 7 9 0 9 13 2
35 1 9 1 0 9 9 9 9 2 12 9 1 9 0 1 9 0 9 9 13 16 9 0 9 13 16 1 1 9 9 9 9 9 13 2
33 1 10 9 0 9 9 1 9 13 16 1 0 9 0 1 9 7 9 1 9 13 16 1 0 9 9 1 1 9 9 13 13 2
23 1 9 9 9 9 9 9 2 9 7 9 9 7 9 16 1 9 7 9 9 0 13 2
32 9 12 9 1 9 9 13 2 1 9 12 9 12 9 1 9 1 1 10 9 1 9 13 16 9 15 14 1 9 9 13 2
34 0 9 2 9 9 7 9 1 9 9 0 13 16 9 15 4 9 9 0 13 16 1 9 9 1 9 15 1 10 9 9 0 13 2
35 1 10 9 9 16 1 9 9 9 9 9 1 9 10 9 2 1 9 10 9 1 9 12 12 9 1 9 2 9 0 1 9 0 13 2
18 1 9 9 9 9 9 2 1 9 9 9 9 1 9 16 0 13 2
30 0 1 9 0 9 1 9 9 9 9 9 2 9 15 14 0 9 13 7 9 9 7 9 9 1 9 9 9 13 2
28 9 9 0 9 9 13 2 9 9 9 9 1 9 9 0 13 7 9 9 9 3 9 1 10 9 4 13 2
35 9 9 9 9 1 9 1 9 0 1 9 9 9 9 1 9 0 13 2 9 9 9 13 16 1 15 7 9 9 0 9 0 9 13 2
31 15 13 2 1 9 0 1 10 9 0 9 7 12 9 1 12 9 9 1 9 12 9 1 12 0 9 9 1 9 13 2
28 9 1 9 1 9 9 12 0 0 9 12 9 0 0 9 0 0 1 9 1 9 9 0 7 9 9 13 2
54 9 0 9 7 9 9 9 9 9 2 9 7 9 3 9 13 2 9 0 4 1 1 9 9 9 0 0 9 0 7 1 9 0 7 1 9 0 1 9 9 13 13 7 7 9 0 14 1 1 1 9 9 13 2
29 9 16 4 1 9 0 7 9 1 9 1 9 9 0 7 1 9 9 0 7 9 1 9 0 0 1 9 13 2
41 1 1 9 10 9 0 2 3 9 9 1 9 1 9 9 0 12 9 7 1 9 9 12 13 16 9 9 9 9 2 9 1 9 7 9 9 1 15 0 13 2
46 1 9 9 0 9 2 0 9 9 9 9 0 9 12 2 12 9 7 1 9 9 9 12 2 12 9 7 1 9 9 9 9 0 7 10 9 0 1 9 9 9 1 0 4 13 2
11 9 0 4 9 1 9 9 9 13 13 2
42 9 0 9 7 9 9 1 9 9 9 0 3 9 12 0 0 9 12 7 1 1 9 0 9 9 2 9 7 9 13 7 9 9 9 10 9 1 10 9 9 13 2
53 9 9 1 9 12 0 1 9 0 9 13 2 9 0 9 9 1 9 9 9 7 9 9 9 0 9 9 1 9 0 2 9 0 1 9 9 9 7 9 15 1 9 0 1 9 7 9 7 9 9 13 13 2
11 7 15 9 15 13 1 9 15 9 13 2
29 9 9 2 9 9 9 0 9 9 16 3 1 9 0 1 0 9 9 9 9 13 2 1 9 9 9 9 13 2
39 7 1 9 9 3 2 13 2 15 10 9 1 9 9 9 9 13 7 16 9 9 9 2 9 15 13 16 3 1 9 13 7 1 3 9 9 14 13 2
70 15 16 9 12 0 1 9 0 9 9 13 7 3 1 9 9 9 9 13 7 1 9 0 9 9 2 9 2 7 9 0 9 13 7 1 9 9 9 9 13 2 13 2 15 3 1 9 9 9 16 1 9 9 13 16 16 9 15 7 7 9 15 14 1 15 9 9 9 13 2
32 15 1 9 15 16 3 9 9 9 13 7 1 9 0 0 13 2 9 13 2 15 9 15 14 1 3 2 0 9 9 13 2
49 9 9 1 9 1 9 9 9 9 9 9 9 2 9 2 2 9 9 0 9 14 3 0 9 13 7 13 2 9 2 9 0 9 2 9 1 9 1 9 9 15 7 9 9 1 1 9 13 2
64 1 10 9 2 9 9 9 2 9 7 9 9 0 9 9 7 9 0 1 9 2 9 9 13 16 9 9 3 0 2 9 0 15 14 1 13 7 3 9 1 9 9 0 1 9 9 7 9 7 9 9 7 9 1 9 9 1 10 9 1 9 0 13 2
10 9 9 9 9 9 9 0 9 13 2
34 9 9 9 9 12 7 12 0 9 2 1 9 9 0 9 9 2 1 9 0 9 16 9 9 9 9 0 13 13 2 1 9 13 2
45 9 0 9 9 9 9 9 9 2 1 9 10 9 13 2 9 2 9 2 0 9 9 9 9 1 12 7 0 9 9 0 9 7 9 12 12 1 9 9 2 1 9 1 13 2
38 2 9 2 9 0 9 7 9 13 7 9 15 16 1 9 9 1 9 0 13 2 9 9 13 16 2 9 2 15 14 1 9 13 7 1 9 13 2
23 1 9 9 9 9 9 12 1 9 0 9 2 9 3 12 9 1 9 9 9 9 13 2
37 9 9 2 9 9 7 9 9 9 9 3 1 9 9 9 1 9 1 9 1 9 9 1 15 13 1 3 9 9 9 9 2 9 9 0 13 2
56 9 9 1 10 9 9 13 2 15 10 9 14 1 9 9 16 13 2 9 13 2 16 13 9 1 9 13 16 1 9 9 3 3 9 0 7 9 0 7 12 9 9 13 16 1 9 3 10 9 2 9 7 9 9 13 2
7 7 7 9 12 9 13 2
8 7 3 9 15 9 0 13 2
15 3 9 16 9 13 7 0 13 2 9 15 9 0 13 2
36 9 9 9 9 1 15 13 2 3 1 10 9 16 15 1 1 10 9 13 2 1 9 0 1 1 9 9 7 9 7 9 9 3 9 13 2
32 9 9 9 13 2 15 13 15 1 1 9 3 9 13 2 7 9 9 1 12 9 0 1 0 9 9 12 9 0 14 13 2
36 15 9 13 2 15 13 16 1 10 9 9 1 9 9 4 9 9 9 7 7 10 9 14 16 1 9 0 2 7 0 7 7 0 13 13 2
29 16 15 7 3 1 1 15 9 13 16 13 15 0 13 7 15 0 13 2 9 13 15 14 3 1 9 3 13 2
45 9 9 2 9 9 9 12 1 0 9 9 9 13 2 16 0 9 15 1 9 2 9 2 14 9 16 12 0 13 2 13 16 10 9 16 12 9 3 1 9 1 9 1 13 2
29 1 9 9 9 9 9 16 9 9 0 9 1 9 9 9 13 2 15 0 9 4 13 16 10 9 14 9 13 2
36 9 0 9 1 9 9 7 9 0 9 1 9 9 1 9 9 2 9 2 9 7 9 0 7 0 9 0 7 9 9 1 9 9 0 13 2
30 9 9 10 9 12 9 1 9 0 1 9 9 0 9 2 9 9 7 9 0 9 0 9 1 9 9 1 13 13 2
52 1 9 9 9 1 9 10 9 2 9 1 9 9 7 9 15 1 9 0 9 2 1 9 2 1 9 9 7 9 9 7 9 1 9 9 2 9 2 9 2 9 2 9 7 9 1 9 9 3 9 13 2
33 1 0 9 10 9 9 9 9 1 9 0 9 0 9 7 9 9 9 9 0 9 1 9 9 9 0 9 1 9 9 15 13 2
38 1 9 9 9 2 1 9 9 1 9 9 7 9 0 9 16 1 12 9 9 13 13 2 1 9 9 0 1 9 9 0 7 0 1 9 0 13 2
45 1 9 9 9 2 15 0 9 1 9 1 9 9 9 13 16 0 1 12 9 1 10 9 1 9 2 1 15 9 13 13 16 1 10 9 12 9 9 15 14 1 9 9 13 2
11 9 13 9 0 1 9 12 9 0 13 2
13 9 9 1 9 9 9 9 1 9 1 9 13 2
21 9 1 9 9 1 9 9 9 9 1 0 9 9 3 1 9 9 1 9 13 2
27 1 10 9 16 1 9 9 0 9 9 1 9 13 2 0 1 12 9 0 1 9 0 1 9 1 13 2
25 10 9 1 9 9 9 7 9 0 2 9 9 9 2 9 9 0 9 0 9 7 9 9 13 2
19 9 9 1 9 9 9 9 1 9 12 9 1 9 9 0 9 9 13 2
21 10 9 1 9 9 9 0 9 9 7 9 0 7 9 0 9 1 9 0 13 2
26 9 9 9 9 9 9 1 9 9 9 2 12 9 0 9 0 1 9 14 1 9 7 9 1 13 2
26 15 1 9 9 0 13 2 10 9 0 13 9 13 16 9 0 9 15 13 16 9 7 9 9 13 2
48 12 9 0 2 1 9 0 7 1 9 7 9 7 9 0 2 1 9 9 9 7 9 9 13 13 7 15 9 0 13 16 1 10 9 9 13 2 16 13 2 8 8 8 8 8 8 8 2
44 15 4 1 9 9 7 9 13 2 3 3 1 0 9 9 9 2 1 9 15 2 1 9 15 2 1 9 7 1 9 15 16 4 1 15 9 13 2 3 4 15 14 13 2
29 9 0 9 0 7 0 10 9 14 1 9 9 13 7 1 9 13 16 4 10 9 0 9 14 1 9 9 13 2
12 12 9 0 1 9 9 0 1 9 9 13 2
33 9 10 9 2 1 1 9 3 1 9 15 2 7 1 1 9 0 0 9 3 1 9 15 1 9 13 7 10 9 9 14 13 2
100 1 9 9 0 7 0 10 9 9 16 9 15 15 14 1 9 0 7 0 9 7 9 13 16 15 14 1 9 7 1 9 9 0 9 13 2 10 9 0 9 9 14 1 12 9 0 0 1 9 9 9 16 1 9 9 13 13 2 15 16 9 14 1 9 9 15 13 7 1 9 12 9 10 9 0 7 10 9 0 14 13 7 1 15 9 13 7 15 14 9 13 2 16 9 1 9 9 0 13 2
20 3 10 9 14 1 9 15 9 9 13 7 15 15 14 13 7 3 0 13 2
58 3 1 12 9 16 10 9 1 9 0 7 0 9 3 0 0 13 13 3 0 2 0 2 0 2 0 2 1 9 0 16 0 2 0 2 0 2 0 7 1 9 0 2 16 9 9 1 10 9 13 1 9 7 1 9 0 13 2
36 9 10 9 14 13 7 1 15 1 9 13 2 1 15 7 9 9 9 14 16 1 10 9 1 9 13 7 1 10 9 16 9 13 9 13 2
43 3 16 9 1 9 9 13 7 1 10 9 16 9 13 2 13 9 9 15 1 10 9 13 7 15 9 15 13 16 1 9 9 9 15 2 1 9 15 1 10 9 13 2
26 1 9 2 1 9 1 9 9 2 9 16 1 9 13 7 10 9 1 9 7 9 10 9 9 13 2
31 1 10 9 2 9 0 10 9 16 1 9 4 9 14 1 9 0 7 0 15 9 13 7 3 13 2 3 9 0 13 2
12 9 15 14 1 9 13 7 1 9 9 13 2
12 9 3 9 0 1 10 9 9 7 9 13 2
12 1 9 9 13 16 15 1 15 3 9 13 2
37 10 9 9 0 16 9 9 7 3 0 7 0 13 10 3 10 9 14 1 9 7 9 9 13 16 9 9 1 10 9 3 1 9 13 7 13 2
51 0 15 13 16 10 9 2 9 9 1 9 7 9 14 9 13 2 1 15 7 9 7 9 15 9 0 13 2 7 12 9 9 9 16 3 0 13 1 15 1 9 3 3 13 2 1 15 1 9 13 2
15 9 10 3 15 14 0 7 0 13 16 9 9 15 13 2
38 1 9 9 7 9 13 13 16 1 1 9 1 9 9 7 9 0 13 7 15 10 9 13 7 9 15 7 9 9 1 9 7 9 1 15 9 13 2
71 16 7 9 13 7 1 1 9 13 2 10 9 13 1 10 9 13 2 9 16 13 2 9 9 1 10 9 13 16 0 13 2 9 9 13 2 7 9 13 3 2 9 15 10 9 13 7 4 10 9 13 2 15 15 1 13 7 10 9 0 7 0 7 0 14 1 10 9 9 13 2
9 0 13 16 9 16 1 9 13 2
60 9 13 16 3 9 2 9 1 8 9 9 3 0 7 0 15 15 9 13 7 13 16 10 9 14 1 15 13 2 4 3 15 1 15 9 13 2 9 16 0 13 7 15 14 1 9 15 15 13 7 3 9 0 15 14 1 9 9 13 2
34 9 7 9 15 9 9 2 16 9 9 9 2 9 9 3 12 9 3 9 7 9 2 10 9 0 14 1 9 7 9 15 9 13 2
13 9 0 1 10 9 9 9 7 9 15 14 13 2
41 9 0 0 2 9 0 0 2 9 7 9 0 2 0 1 9 7 9 16 0 13 1 12 9 1 9 3 13 2 9 0 0 7 0 14 1 10 9 9 13 2
29 1 10 9 9 2 1 9 7 9 15 2 9 9 9 14 1 9 13 7 0 9 13 2 15 9 0 9 13 2
18 1 9 15 15 2 1 10 9 9 1 9 8 9 1 9 9 13 2
28 3 10 9 9 9 13 2 16 1 9 9 7 9 9 1 9 9 7 1 9 12 0 16 9 9 13 13 2
41 0 9 0 12 9 0 1 15 9 13 2 16 15 3 9 1 9 0 10 9 14 3 0 9 13 2 7 3 9 9 0 13 16 9 1 9 0 9 9 13 2
46 15 3 1 9 9 7 1 15 16 1 9 7 9 2 3 9 13 13 16 1 1 9 9 9 0 9 13 7 9 15 9 13 16 9 0 13 10 0 9 14 1 10 9 0 13 2
20 3 1 9 0 1 1 9 0 7 1 9 0 1 1 9 10 9 9 13 2
45 15 16 15 1 10 9 9 13 2 1 9 12 1 9 0 9 9 9 9 9 9 9 13 16 9 1 10 9 13 7 15 1 9 15 16 9 13 7 0 7 0 13 9 13 2
35 3 15 9 1 10 9 13 16 1 9 10 9 13 2 0 9 10 9 0 7 0 1 15 9 13 16 15 3 15 1 15 14 9 13 2
12 10 9 2 0 2 0 2 0 7 0 13 2
11 0 13 2 1 9 1 15 9 9 13 2
17 0 13 2 9 15 1 9 2 1 9 9 7 9 7 9 13 2
8 0 13 2 0 7 0 13 2
37 0 13 2 1 10 9 0 0 9 3 1 9 2 1 9 9 2 10 9 2 0 1 9 7 9 13 7 9 15 14 15 0 13 2 0 13 2
21 9 9 7 9 9 13 2 9 2 0 2 9 2 0 2 9 2 9 1 9 2
16 0 13 7 3 9 0 1 9 2 15 14 0 7 0 13 2
13 0 13 2 9 15 14 1 9 7 9 9 13 2
10 1 9 2 9 7 9 9 15 13 2
19 0 13 16 9 9 2 7 9 9 2 16 9 13 2 9 7 9 13 2
19 3 0 13 2 3 9 15 14 1 9 0 13 2 3 1 9 9 13 2
4 3 0 13 2
30 16 9 15 14 1 9 16 15 0 13 2 9 13 16 1 9 9 9 13 1 9 7 9 9 15 14 1 9 13 2
11 3 0 7 0 7 0 7 9 9 13 2
28 1 0 9 10 9 2 1 9 9 1 3 9 1 12 7 12 0 2 10 9 14 1 9 10 9 13 13 2
57 15 15 1 10 9 14 3 0 13 2 0 9 7 9 15 10 3 13 16 1 9 9 15 14 1 9 9 13 13 7 9 10 9 16 1 15 3 9 9 13 2 9 15 13 7 0 13 16 10 9 1 15 0 1 4 13 2
41 3 3 1 15 7 9 9 9 13 7 9 9 7 9 1 9 3 13 2 1 10 9 16 0 10 9 16 13 9 14 1 9 9 13 2 13 7 1 9 13 2
25 16 15 13 16 16 9 0 1 9 9 13 2 9 14 1 9 13 16 9 9 14 1 15 13 2
31 0 13 16 1 10 9 16 9 9 1 10 9 13 13 2 3 9 9 2 7 9 9 7 10 9 16 1 15 9 13 2
24 9 15 1 10 9 13 16 9 16 15 1 9 15 0 13 2 1 10 9 9 1 9 13 2
76 3 9 10 9 1 9 9 1 15 13 16 16 9 8 9 1 12 9 13 2 3 0 13 16 9 15 14 13 7 1 9 15 1 3 13 7 10 9 16 15 1 9 13 13 2 15 14 1 9 15 9 13 2 13 2 10 9 9 13 2 9 15 14 13 2 7 9 10 9 14 1 9 9 13 13 2
28 1 12 9 0 1 9 9 9 13 2 9 9 9 9 1 9 13 2 7 10 9 9 13 7 9 9 13 2
48 12 9 13 1 9 9 13 16 9 9 10 9 1 9 15 9 13 2 9 0 13 7 13 1 9 1 9 9 9 13 7 9 15 14 0 13 2 3 16 13 1 9 10 9 2 9 13 2
53 3 1 9 2 3 9 1 9 2 1 1 9 7 7 9 2 9 0 1 9 13 2 3 12 9 12 9 1 9 9 9 9 9 9 16 12 1 9 9 13 1 9 9 13 16 15 9 13 2 7 9 13 2
7 9 9 13 7 9 13 2
21 15 9 0 13 16 9 15 14 0 13 13 2 16 3 0 13 1 15 9 13 2
22 3 9 1 9 13 7 9 15 15 14 0 13 7 1 9 13 16 9 15 14 13 2
14 9 16 1 9 0 2 10 9 7 9 14 9 13 2
16 9 15 9 13 16 9 0 15 14 1 9 7 9 9 13 2
17 16 1 9 0 13 2 1 7 1 9 15 13 2 9 1 13 2
29 1 9 2 9 1 9 9 9 0 2 3 1 9 16 9 9 1 15 15 13 9 13 16 9 1 15 9 13 2
12 12 9 0 0 9 13 7 9 15 14 13 2
19 9 16 9 14 13 13 2 9 13 2 15 9 0 0 1 9 9 13 2
28 10 9 0 1 15 16 16 9 13 2 13 9 9 13 2 16 1 9 9 13 7 9 13 2 6 9 9 2
6 1 15 9 13 13 2
49 9 7 9 15 9 10 9 14 13 2 16 1 15 9 13 7 9 13 16 1 9 15 9 13 2 0 13 1 9 13 7 13 2 9 15 14 13 2 15 16 13 7 0 13 9 15 14 13 2
21 3 1 9 9 13 13 2 9 13 16 15 3 16 15 14 1 10 9 0 13 2
14 9 1 9 0 15 9 13 16 1 15 0 9 13 2
43 1 9 0 0 2 16 7 9 9 14 1 10 9 7 9 9 13 2 13 2 8 8 8 2 3 2 9 9 7 9 13 2 16 9 13 2 15 2 9 10 9 13 2
4 15 0 13 2
25 1 9 9 10 9 7 13 9 13 2 1 9 7 9 13 2 1 9 0 0 13 7 9 13 2
52 12 1 9 9 9 15 3 13 16 15 0 9 13 2 3 9 13 2 3 9 13 2 3 9 15 14 1 9 9 13 2 3 1 9 9 13 2 3 1 15 3 13 2 3 1 15 0 13 2 0 13 2
12 10 9 15 13 16 9 9 14 0 15 13 2
19 15 9 16 9 0 9 7 1 9 9 7 9 7 9 2 9 0 13 2
8 1 9 9 2 0 0 13 2
18 1 9 9 9 2 1 9 9 9 9 2 0 7 0 7 0 13 2
18 9 0 15 16 1 9 15 13 2 0 2 9 0 15 0 7 0 2
11 3 1 9 2 15 14 0 7 0 13 2
48 1 9 1 9 9 0 16 3 4 13 9 9 3 0 13 1 15 15 9 7 9 13 2 9 1 13 2 1 15 7 9 15 14 9 13 2 16 10 9 0 13 9 9 15 14 9 13 2
7 10 9 0 9 9 13 2
18 15 14 16 1 10 9 2 1 10 9 2 1 10 9 0 9 13 2
32 9 15 10 13 16 9 13 9 0 4 1 9 7 1 9 0 13 2 3 2 1 9 0 7 0 16 13 0 7 0 13 2
17 9 9 0 7 0 13 2 7 9 7 9 7 9 15 0 13 2
17 15 1 9 2 1 9 2 1 9 0 7 1 9 3 0 13 2
12 10 9 1 9 0 2 1 9 3 0 13 2
35 9 15 1 9 2 9 0 13 2 1 9 9 2 3 0 13 2 0 16 13 2 10 9 9 7 9 7 9 16 13 2 3 9 13 2
18 9 7 9 15 15 14 1 9 15 15 1 9 0 13 2 0 13 2
5 1 15 9 13 2
21 16 9 15 14 0 13 2 1 9 15 9 13 13 2 7 9 1 9 0 13 2
29 9 13 1 9 15 1 9 9 13 7 1 9 9 13 2 15 15 16 1 3 9 9 13 7 1 9 9 13 2
31 9 14 1 9 9 13 2 1 9 9 13 2 1 9 9 9 14 13 2 1 9 15 9 13 7 1 15 9 9 13 2
27 9 15 12 9 13 2 9 15 1 9 13 16 1 9 9 0 13 13 9 9 15 9 9 7 9 13 2
21 13 16 3 12 9 1 9 16 1 9 9 3 9 0 9 15 14 0 13 13 2
16 8 9 9 13 16 3 12 9 1 9 9 15 9 0 13 2
7 9 9 0 7 0 13 2
28 10 9 16 9 0 14 1 9 7 9 0 9 13 7 9 13 2 10 9 1 0 1 9 9 1 9 13 2
6 9 9 1 15 13 2
36 1 9 15 2 9 15 14 9 13 15 10 9 13 16 9 0 10 9 9 9 9 9 9 13 7 1 9 1 1 15 2 10 14 3 13 2
17 9 15 10 3 9 13 16 9 15 1 9 1 9 9 9 13 2
12 9 9 14 1 9 0 7 9 0 9 13 2
48 9 9 7 9 9 7 9 13 2 13 9 9 13 16 1 15 15 7 16 1 15 2 15 15 16 0 9 13 2 9 15 12 9 0 1 9 12 9 9 13 7 12 9 1 9 0 13 2
19 9 0 1 9 14 1 9 7 9 7 9 7 9 7 9 7 9 13 2
10 1 9 0 9 7 9 7 9 13 2
32 3 1 9 9 2 1 9 9 7 9 9 7 1 9 9 9 16 10 9 16 13 1 10 9 0 12 9 1 9 9 13 2
5 15 16 9 13 2
22 13 2 8 8 8 8 2 16 9 0 9 13 16 10 15 1 15 9 13 13 2 2
15 9 15 9 13 16 1 9 9 3 15 14 13 9 13 2
20 15 3 9 1 9 13 16 13 10 9 0 0 14 16 0 13 2 9 13 2
7 3 1 9 2 0 13 2
6 1 9 15 0 13 2
10 1 9 15 2 9 10 0 9 13 2
27 1 9 15 2 1 10 9 16 3 9 9 13 2 9 9 0 9 1 1 9 0 7 9 9 0 13 2
6 15 9 0 9 13 2
11 9 0 9 15 13 2 0 7 0 13 2
65 9 16 9 9 9 1 9 14 13 10 9 0 2 10 9 9 2 10 9 9 1 9 1 1 9 2 10 9 0 2 10 9 1 9 0 9 10 3 9 0 7 0 7 0 1 9 10 9 9 13 16 0 13 7 9 13 16 15 3 13 15 14 9 13 2
24 15 9 7 9 9 7 9 13 2 13 9 9 13 2 16 1 15 15 2 7 16 1 15 2
16 15 15 16 0 9 13 2 9 9 16 1 10 9 9 13 2
27 1 10 9 16 9 4 9 13 2 15 10 9 16 3 7 3 1 10 9 9 13 7 9 13 9 13 2
51 10 15 9 7 10 15 9 1 9 13 2 12 9 16 1 15 13 2 16 9 0 1 15 7 9 1 9 15 13 7 1 15 9 13 7 1 1 15 3 0 13 2 7 0 13 1 9 15 9 13 2
21 16 9 13 1 10 9 1 9 15 13 2 9 16 9 13 2 7 15 0 13 2
30 3 7 3 9 13 2 9 1 15 9 9 1 15 13 2 12 9 1 9 15 15 9 13 16 1 15 10 9 13 2
20 9 13 2 16 13 1 15 9 13 2 9 0 13 7 9 1 9 0 13 2
11 1 10 9 0 15 15 13 16 0 13 2
5 3 9 9 13 2
18 9 1 15 9 13 2 7 15 13 2 9 9 9 13 2 15 13 2
5 15 16 0 13 2
15 16 1 9 9 9 13 2 3 9 13 9 3 13 13 2
22 15 9 14 9 13 7 13 2 3 13 2 13 2 3 2 13 2 3 0 4 13 2
32 1 3 9 9 13 16 13 15 4 1 9 9 13 2 9 13 16 1 3 9 2 9 3 9 13 16 9 4 1 9 13 2
14 9 14 12 9 13 2 10 1 9 0 9 9 13 2
33 15 1 9 2 9 13 16 9 15 0 13 2 7 9 16 13 16 15 9 0 13 2 1 15 9 13 7 1 1 15 0 13 2
21 9 16 13 16 9 13 2 7 9 15 14 9 13 7 1 9 13 2 3 9 2
32 9 0 9 12 1 9 9 16 13 2 16 9 16 15 14 1 9 13 2 9 1 9 15 13 7 1 9 9 9 16 13 2
19 0 3 1 9 9 2 9 9 1 9 13 2 7 9 15 14 9 13 2
36 15 9 13 16 1 9 15 9 7 9 0 7 9 0 1 9 0 3 13 2 7 9 1 9 16 1 9 15 9 9 13 2 3 0 13 2
83 10 9 0 2 10 9 0 2 10 9 0 7 1 9 2 9 13 16 9 9 14 16 0 12 9 13 1 12 9 1 9 13 7 9 7 9 14 3 13 7 9 14 9 13 2 16 15 9 0 13 2 9 1 15 9 9 1 9 9 9 14 1 9 13 13 2 7 15 1 1 9 13 7 1 1 9 13 7 9 7 9 13 2
9 15 2 9 1 9 10 9 13 2
2 9 2
13 1 15 9 13 16 15 14 1 9 9 9 13 2
34 15 13 16 9 15 0 1 9 9 13 2 15 14 1 10 9 0 7 0 0 13 7 1 10 9 0 2 15 14 1 10 9 13 2
2 9 2
44 9 9 9 14 1 9 9 15 13 2 9 1 9 9 7 9 1 9 10 9 14 9 15 13 2 15 14 1 9 0 9 9 15 9 13 7 9 14 9 10 9 9 13 2
26 15 0 13 15 9 16 1 9 0 7 1 10 9 0 1 9 9 13 2 1 9 3 15 9 13 2
36 10 9 16 16 0 13 16 3 1 9 15 9 13 16 9 13 2 3 15 1 15 9 13 2 1 15 7 9 0 14 1 15 15 9 13 2
9 3 3 10 9 2 9 0 13 2
35 3 1 9 0 9 16 1 9 9 13 2 9 1 9 0 7 0 9 7 9 1 9 7 9 0 9 9 16 3 1 10 9 9 13 2
19 9 2 12 9 0 1 9 12 9 9 13 7 12 9 1 9 0 13 2
39 15 1 9 15 3 13 2 9 0 13 2 9 0 1 9 0 7 0 7 0 9 7 12 9 1 9 7 12 9 1 9 9 10 9 7 10 9 13 2
25 3 1 9 16 1 9 9 1 9 13 2 15 1 9 7 9 9 13 2 10 9 3 0 13 2
18 15 13 1 9 9 13 16 9 15 14 0 7 1 9 9 9 13 2
17 7 3 1 10 12 9 0 9 0 0 7 9 0 9 9 13 2
5 16 9 0 13 2
21 9 0 2 9 0 13 16 1 9 9 0 1 9 13 13 2 7 0 16 13 2
48 1 15 7 9 1 9 1 9 13 2 7 3 9 0 13 2 1 9 9 2 1 9 9 9 13 7 9 0 9 1 9 2 1 9 2 1 9 7 1 9 0 0 7 9 1 9 13 2
9 1 9 0 2 9 0 0 13 2
16 9 1 3 13 13 7 10 9 14 1 9 9 15 13 13 2
39 3 1 9 15 1 9 0 7 0 15 16 12 9 1 9 7 1 9 15 15 0 1 9 13 2 7 10 9 9 7 10 9 0 9 0 14 9 13 2
28 3 9 1 10 9 13 2 3 9 0 1 9 13 2 7 1 15 15 0 16 13 7 9 0 9 16 13 2
24 9 0 0 13 2 1 9 0 2 3 0 1 9 2 1 9 9 0 2 3 0 1 9 2
10 0 13 16 10 9 0 1 9 13 2
51 3 16 9 15 2 9 0 7 0 13 2 13 1 9 9 9 14 1 9 15 15 9 13 7 9 9 13 2 7 3 13 9 13 2 13 3 15 16 1 3 13 2 3 1 0 12 9 3 0 13 2
12 0 13 16 10 9 1 15 0 9 9 13 2
65 10 9 16 9 15 0 13 16 12 7 12 9 3 1 15 3 9 1 9 9 13 16 16 0 13 2 1 10 9 0 3 7 0 2 7 0 16 9 0 15 13 9 13 13 2 7 9 7 9 9 7 9 10 9 15 14 9 13 7 0 13 7 1 13 2
52 1 9 2 9 13 2 7 9 13 2 9 13 2 7 9 13 2 9 0 13 2 7 1 1 9 9 7 9 9 13 2 9 9 7 9 13 2 7 1 9 9 13 2 3 9 2 3 16 10 9 13 2
28 10 9 16 15 9 13 2 9 15 13 2 15 1 9 10 9 0 0 9 13 2 1 9 15 9 9 13 2
31 3 1 9 0 7 1 15 9 2 10 9 16 1 9 9 7 9 9 13 2 9 9 13 2 9 15 2 9 9 13 2
40 15 0 13 16 1 9 7 9 15 9 13 2 7 15 9 0 9 13 7 13 16 10 9 9 2 9 9 9 7 9 9 2 1 3 9 7 9 9 13 2
48 16 9 9 13 2 4 13 16 1 10 9 2 9 9 3 3 9 13 2 15 16 9 0 7 0 14 13 2 9 7 9 7 9 0 0 7 1 1 9 7 0 1 9 9 9 0 13 2
10 9 9 13 2 7 9 9 3 13 2
18 9 0 1 9 13 2 7 10 9 0 9 1 9 9 0 13 13 2
56 9 1 0 15 16 12 9 0 0 13 2 15 14 1 9 0 7 0 9 13 7 1 9 9 7 9 9 9 13 2 10 9 9 0 13 1 15 9 13 7 15 14 9 13 2 3 13 2 10 9 13 2 0 15 13 2
15 1 9 9 13 2 7 9 1 1 9 7 9 7 9 2
20 9 1 9 0 13 7 15 9 13 2 7 9 1 9 0 1 3 9 13 2
7 3 0 1 9 13 2 2
10 15 16 9 0 13 2 13 9 13 2
19 15 1 15 9 7 15 9 12 9 0 9 9 13 16 0 1 9 13 2
40 3 9 16 0 13 2 16 9 9 16 9 15 15 14 13 2 15 14 13 2 0 13 2 15 14 13 2 0 13 2 1 10 9 13 2 9 0 14 13 2
5 15 16 9 13 2
43 16 12 9 0 13 7 1 9 9 13 3 10 9 9 16 0 9 9 1 9 13 7 13 2 15 16 13 9 14 1 9 9 13 2 9 13 9 0 1 15 9 13 2
33 16 9 0 1 9 13 2 0 1 9 9 9 13 2 3 9 15 13 13 2 3 9 15 1 9 9 13 2 3 9 9 13 2
26 6 2 9 0 13 16 1 9 9 7 9 7 9 15 15 2 10 3 14 16 9 15 13 2 13 2
12 10 9 2 9 13 2 10 9 2 9 13 2
37 9 14 1 9 7 1 9 13 2 10 9 13 2 9 0 13 2 10 9 13 2 9 0 0 13 2 10 9 13 2 9 13 2 9 16 15 2
33 0 13 16 1 9 16 1 9 15 7 9 15 9 13 13 7 1 9 15 12 9 0 7 9 9 13 2 9 0 13 9 13 2
37 3 2 15 9 14 3 1 9 0 7 3 1 9 0 13 2 15 9 14 1 9 13 7 9 15 1 9 9 1 9 2 9 0 14 9 13 2
22 9 15 9 0 13 13 2 1 9 0 13 2 1 9 0 13 2 9 9 13 13 2
20 1 10 9 0 2 9 0 1 9 2 9 2 9 7 9 9 0 13 13 2
14 9 12 9 9 1 15 9 13 13 7 1 15 13 2
14 1 9 9 0 3 9 13 2 1 10 9 0 13 2
8 9 1 9 1 10 9 13 2
5 3 10 9 13 2
12 15 1 10 9 9 1 10 9 14 9 13 2
30 3 16 13 10 9 14 1 12 9 9 13 2 15 9 13 9 2 7 9 12 9 0 13 7 9 0 1 15 13 2
28 9 15 1 1 9 13 16 15 15 1 1 9 13 7 15 1 9 1 15 9 13 2 9 0 2 9 13 2
20 9 1 9 7 9 7 9 0 7 0 13 2 13 9 15 1 9 9 13 2
6 9 0 2 9 13 2
26 9 13 16 9 2 9 0 13 2 0 1 3 1 9 9 13 2 15 15 16 1 15 15 9 13 2
24 1 1 9 9 2 10 9 16 1 1 15 9 7 9 0 13 2 1 9 16 0 9 13 2
46 1 9 9 13 2 1 9 9 9 13 2 1 9 9 13 2 1 9 0 9 13 2 1 9 0 9 13 2 15 9 9 0 13 7 9 1 9 7 9 15 15 9 14 9 13 2
25 1 9 9 15 7 9 0 9 0 9 1 1 9 1 9 9 1 9 9 0 1 9 9 13 2
9 15 1 12 1 9 0 9 13 2
29 12 9 3 1 9 1 9 0 1 12 9 9 13 16 3 1 9 9 2 9 1 9 15 1 9 0 9 13 2
27 3 13 9 15 14 9 13 7 16 1 9 1 15 16 15 9 9 14 13 13 1 9 0 9 0 13 2
70 9 0 2 1 9 9 1 15 2 9 1 9 7 9 9 16 15 0 13 3 0 13 2 7 1 9 1 9 9 1 1 1 9 7 9 15 1 9 0 16 1 10 9 9 13 2 9 9 13 0 9 13 7 4 1 9 10 9 9 13 16 1 9 0 1 9 15 9 13 2
24 1 10 9 15 13 1 1 9 9 9 0 1 9 9 0 1 9 9 13 7 9 9 13 2
56 1 10 9 9 13 16 1 9 1 9 9 2 15 14 9 13 2 16 1 9 0 13 1 9 9 16 10 9 1 15 9 13 1 9 9 9 9 15 9 7 9 9 1 9 14 13 16 9 1 9 0 1 15 9 13 2
35 0 9 0 0 0 9 0 9 16 0 1 12 9 1 9 15 13 2 1 9 0 9 9 15 14 1 9 0 1 9 1 9 0 13 2
53 0 1 9 0 9 1 9 1 9 9 1 9 1 9 1 9 0 9 9 0 9 9 2 1 1 9 9 9 1 9 0 7 9 15 1 9 0 9 13 16 3 12 9 3 1 9 10 9 1 15 9 13 2
45 1 10 9 1 9 13 2 1 9 1 9 9 9 0 1 9 2 9 0 9 9 16 1 9 1 9 0 1 9 9 0 14 4 13 2 0 1 9 0 15 14 1 9 13 2
34 15 1 9 13 16 12 9 0 9 9 13 2 9 0 0 9 9 9 3 1 12 9 0 1 9 9 15 1 9 0 9 4 13 2
53 10 9 14 9 9 9 9 1 9 9 2 9 7 9 9 9 1 9 0 15 1 9 9 9 9 9 9 1 9 9 9 16 1 15 13 13 9 0 9 9 9 9 1 3 9 9 4 13 2 9 13 13 2
6 9 1 9 9 13 2
29 9 3 9 7 9 9 2 9 9 1 9 9 9 9 9 13 16 4 1 9 12 9 1 9 0 14 9 13 2
25 1 9 9 9 2 9 9 1 9 9 9 9 13 1 9 9 9 15 1 9 9 0 15 13 2
23 12 9 0 1 9 0 1 9 9 13 7 12 12 9 1 9 10 9 9 14 9 13 2
21 9 16 9 15 0 13 13 1 9 1 9 9 9 15 1 9 0 0 13 13 2
27 9 9 13 16 0 9 0 9 1 15 13 13 7 1 9 9 0 9 3 1 9 1 9 9 13 13 2
22 9 9 0 9 16 9 9 9 9 0 9 13 13 2 9 0 9 3 9 13 13 2
17 9 9 3 1 9 9 7 1 9 9 9 13 16 0 9 13 2
28 9 16 1 9 9 1 9 9 9 9 1 9 13 2 9 13 16 0 1 9 0 1 9 1 9 13 13 2
23 9 9 9 13 2 9 1 9 9 0 9 13 13 2 16 10 9 1 9 9 9 13 2
9 9 1 9 9 9 1 9 13 2
30 9 9 9 9 9 9 9 2 1 9 0 1 9 0 7 9 0 9 0 13 7 9 0 12 9 1 9 13 13 2
13 9 0 9 9 13 9 0 1 9 9 9 13 2
18 1 9 9 0 1 9 10 9 16 1 12 9 9 9 0 13 13 2
29 10 9 1 9 12 2 12 9 9 1 9 9 0 9 9 9 1 9 0 2 9 9 1 9 9 14 9 13 2
23 10 9 1 9 0 1 9 0 9 1 9 9 9 2 9 2 9 9 7 9 9 13 2
18 9 9 9 9 2 9 10 9 14 9 9 2 9 10 9 9 13 2
35 9 0 9 1 9 0 10 9 12 9 9 13 16 9 15 14 9 7 9 0 0 13 7 1 10 9 9 9 9 1 9 14 0 13 2
40 1 9 9 9 2 0 9 0 1 10 9 1 9 9 0 9 9 9 9 13 2 7 9 10 9 3 9 9 13 7 13 16 10 9 9 0 1 9 13 2
35 9 9 9 9 13 2 10 9 1 9 0 9 1 9 7 9 9 1 9 9 9 15 4 13 16 9 9 1 9 0 7 0 4 13 2
24 10 9 7 9 16 1 9 0 13 13 2 1 9 9 9 9 0 2 1 9 9 9 13 2
23 12 9 9 0 9 1 9 9 9 12 9 9 9 9 1 9 9 9 0 14 9 13 2
25 9 9 2 9 0 1 9 12 12 9 13 7 9 9 9 9 9 1 1 10 9 9 9 13 2
28 9 9 9 9 9 9 9 9 0 13 2 9 9 9 1 9 9 1 9 12 9 9 1 9 0 9 13 2
22 1 10 9 2 9 9 1 9 9 9 9 2 9 12 9 0 12 9 14 9 13 2
11 9 10 9 1 9 9 9 0 9 13 2
36 10 9 1 9 1 9 9 2 1 0 9 9 2 9 9 2 9 7 9 9 14 16 1 9 9 9 0 13 2 1 9 9 9 4 13 2
18 9 9 0 1 9 9 9 12 9 9 14 12 12 9 9 13 13 2
22 9 1 9 0 1 12 12 0 12 1 12 0 0 9 9 14 1 1 9 9 13 2
10 9 10 9 9 9 9 14 9 13 2
16 12 9 0 1 9 9 1 9 9 1 9 3 9 9 13 2
60 1 9 9 9 1 9 2 9 9 9 12 0 0 16 3 9 15 14 1 9 9 9 9 9 13 2 9 13 2 9 13 16 9 0 15 1 9 9 1 9 9 3 9 1 9 9 9 3 1 9 9 1 15 2 1 9 0 0 13 2
23 15 1 10 9 13 16 13 1 12 9 9 1 9 2 0 1 12 9 9 1 9 13 2
27 15 13 2 1 9 9 1 9 12 2 1 9 0 1 0 9 10 9 9 13 7 9 15 14 0 13 2
45 1 9 10 9 2 9 9 1 9 10 9 1 9 2 1 9 0 1 9 9 7 9 0 1 9 0 0 13 13 2 7 1 9 13 16 10 9 1 1 9 9 16 0 13 2
17 9 13 2 9 3 9 2 9 9 7 9 1 10 9 0 13 2
30 15 13 2 10 9 1 9 9 0 1 9 0 13 13 7 16 1 9 9 13 2 12 9 0 0 1 9 0 13 2
20 10 9 9 13 16 9 12 9 9 0 9 1 9 2 1 9 0 9 13 2
14 9 0 9 9 14 9 7 1 3 13 7 3 13 2
28 10 9 13 2 1 9 13 9 0 14 1 9 1 9 0 1 9 9 0 3 9 7 9 1 9 9 13 2
28 9 0 9 1 9 9 9 1 9 1 1 9 1 9 0 9 0 9 0 9 9 9 14 1 15 15 13 2
17 10 9 9 9 1 9 1 9 12 1 12 1 9 9 9 13 2
13 9 9 0 10 9 12 1 12 1 9 9 13 2
14 9 9 1 0 9 9 9 9 16 1 9 0 13 2
24 1 9 0 9 0 9 9 0 9 0 1 9 9 2 12 9 9 7 9 1 15 9 13 2
10 1 10 9 9 0 1 9 9 13 2
28 9 0 1 9 1 9 9 0 1 9 9 2 9 2 9 7 9 0 13 7 1 9 10 9 14 9 13 2
34 1 9 0 9 0 1 9 9 2 9 9 12 9 9 14 0 9 9 0 13 7 9 0 0 1 12 9 0 1 9 9 9 13 2
21 1 10 9 9 9 0 9 9 7 0 9 9 10 9 14 16 1 15 9 13 2
21 9 2 9 7 9 1 9 12 9 0 9 9 1 9 9 0 1 9 9 13 2
10 10 9 9 3 1 9 0 4 13 2
6 9 9 3 9 13 2
15 9 0 7 0 2 9 0 0 9 9 9 14 9 13 2
12 1 10 9 4 1 9 9 9 0 9 13 2
22 9 9 9 7 9 9 9 2 12 9 14 9 13 16 1 1 9 9 0 9 13 2
18 10 9 0 7 0 0 16 9 9 13 13 2 9 1 9 13 13 2
36 9 16 10 12 9 3 0 9 13 2 9 9 15 1 9 0 9 13 7 1 9 0 9 9 14 9 13 7 10 9 9 1 1 9 13 2
12 10 9 1 9 12 9 7 9 9 0 13 2
32 9 0 9 13 7 1 1 15 9 7 3 1 15 9 7 9 0 9 9 7 1 9 16 9 7 9 0 9 9 9 13 2
22 9 16 12 9 9 13 2 10 9 0 9 1 9 13 16 9 9 9 9 15 13 2
24 10 9 0 13 9 0 9 9 14 9 13 16 1 9 9 10 9 1 9 9 0 9 13 2
28 1 9 9 2 1 9 9 1 9 9 2 16 9 16 1 9 9 0 13 2 9 9 9 0 9 9 13 2
10 16 9 0 0 9 0 1 9 13 2
42 9 1 9 9 13 16 1 0 9 9 0 13 2 7 9 1 9 9 1 15 9 13 16 1 9 9 9 0 13 2 7 9 10 9 15 1 9 0 3 13 13 2
12 1 9 0 13 13 16 9 0 9 0 13 2
22 3 3 15 10 9 13 16 1 9 9 0 9 3 0 0 13 7 3 9 0 13 2
18 15 15 9 13 7 15 9 13 2 16 1 9 9 1 9 0 13 2
18 3 1 9 9 15 15 13 7 10 9 0 1 10 9 1 1 13 2
11 15 2 16 9 15 13 7 7 9 15 2
10 16 9 15 13 7 7 9 0 15 2
17 9 10 9 9 1 9 15 7 9 10 9 9 1 9 15 13 2
9 9 15 15 9 0 9 9 13 2
2 9 2
7 3 9 9 13 3 13 2
9 9 9 9 9 9 12 9 13 2
27 1 9 0 9 9 0 2 9 9 13 1 9 9 9 1 9 0 1 9 0 7 9 0 0 0 13 2
18 9 9 9 13 16 9 9 10 9 1 9 0 1 12 9 9 13 2
30 1 1 10 9 2 9 9 9 7 9 1 9 14 1 9 12 1 12 1 9 3 9 9 7 9 9 9 9 13 2
31 10 9 1 13 10 9 9 9 9 0 13 2 9 9 7 9 0 1 9 0 0 2 9 0 7 9 0 0 0 13 2
20 10 9 9 13 2 9 9 12 9 0 0 9 9 16 9 9 7 9 13 2
17 9 13 2 1 10 9 9 7 9 0 1 10 9 3 0 13 2
20 9 9 13 16 9 9 1 10 9 9 0 1 9 9 7 9 0 9 13 2
28 9 0 9 9 9 13 9 7 9 0 0 1 9 9 9 13 7 10 9 9 9 7 9 1 1 9 13 2
24 1 9 9 12 1 9 9 12 9 9 9 0 2 9 9 9 9 9 0 9 9 0 13 2
16 1 10 9 12 9 9 15 14 1 15 7 9 15 9 13 2
34 15 13 9 13 1 9 10 9 2 9 3 1 9 1 9 9 0 7 9 9 13 2 1 9 13 16 3 0 13 13 7 13 13 2
10 9 9 1 9 3 2 9 9 13 2
4 13 9 13 2
11 6 2 1 9 15 7 9 9 0 13 2
19 3 16 13 9 2 3 1 9 7 9 7 15 13 2 3 9 13 13 2
6 9 9 3 9 13 2
4 1 15 13 2
4 3 9 13 2
7 9 9 9 9 9 13 2
8 9 9 13 1 9 15 13 2
8 9 3 1 9 9 4 13 2
25 9 12 7 0 9 9 9 0 9 9 9 9 9 1 9 12 9 1 9 7 9 9 9 13 2
23 1 10 9 9 9 7 9 9 2 9 9 2 9 9 7 9 9 9 15 14 9 13 2
46 9 9 16 1 1 9 9 0 9 7 9 9 2 9 15 0 13 13 9 9 9 1 9 9 13 7 0 13 9 15 14 1 12 9 9 13 7 9 9 15 14 1 12 9 13 2
32 1 9 12 9 0 9 9 9 0 9 1 9 9 13 16 9 10 9 9 14 1 1 9 9 9 9 9 9 1 9 13 2
27 1 9 12 9 9 9 12 9 9 13 16 9 9 9 14 1 9 13 16 0 9 10 9 1 9 13 2
21 16 9 9 9 7 9 9 1 9 1 9 15 1 9 9 1 9 0 9 13 2
17 9 0 9 9 9 0 9 9 2 9 9 9 9 9 9 13 2
42 1 9 10 9 9 9 9 7 9 9 1 9 1 9 12 7 12 9 1 9 0 7 0 9 9 9 13 7 9 9 1 9 0 9 9 9 9 14 1 9 13 2
28 9 9 9 9 16 1 9 9 0 9 9 0 9 9 13 2 9 9 9 3 1 9 1 9 1 9 13 2
43 9 9 16 1 1 9 0 9 0 9 9 7 9 9 9 2 9 15 0 13 13 3 0 13 1 12 9 1 9 9 9 13 16 12 9 13 7 1 9 1 3 13 2
15 0 9 9 9 1 9 9 9 1 9 12 1 9 13 2
34 9 9 9 3 1 10 9 1 9 7 9 9 9 15 14 1 1 9 15 9 13 13 2 1 9 13 2 7 9 9 1 9 13 2
37 12 9 0 0 16 0 9 3 1 0 9 9 9 9 0 1 9 9 14 1 9 9 13 2 3 1 9 13 0 9 14 1 10 9 9 13 2
49 1 0 9 9 9 9 2 9 9 9 1 9 0 9 1 9 12 0 2 9 1 12 1 9 0 9 13 7 1 9 10 9 9 13 16 16 9 7 9 9 1 9 15 9 13 13 7 6 2
44 1 9 16 1 10 9 0 9 13 2 1 10 9 9 13 13 16 9 1 9 0 2 9 0 1 9 9 13 7 9 1 15 14 1 9 9 0 7 1 9 0 13 13 2
43 9 9 1 9 9 15 9 13 13 16 9 0 16 1 9 1 9 9 0 9 7 1 9 15 16 9 9 0 13 13 2 13 7 1 15 10 9 1 9 0 0 13 2
37 1 9 9 0 2 9 15 15 14 16 1 9 7 9 15 13 7 9 7 9 16 9 9 15 14 9 13 2 1 9 0 1 9 9 1 13 2
12 9 1 1 9 9 0 7 3 9 9 13 2
45 15 3 9 9 13 16 15 13 9 9 13 7 15 1 15 9 0 13 2 3 2 7 9 0 1 10 9 7 1 10 9 2 1 9 7 9 9 7 1 9 15 0 0 13 2
17 9 9 7 9 3 1 15 1 9 2 0 13 2 9 0 13 2
50 12 9 1 9 9 13 13 1 9 9 13 13 7 15 15 14 9 0 13 2 3 7 7 13 1 9 13 16 13 15 14 13 2 16 9 13 13 7 1 9 15 13 9 15 14 9 15 15 13 2
8 3 10 9 13 7 13 2 2
10 3 9 3 13 7 9 15 13 2 2
5 15 3 0 13 2
30 3 1 15 16 9 13 2 12 0 13 2 12 0 0 1 9 15 15 13 2 9 1 9 7 9 9 2 0 0 2
5 9 15 14 13 2
22 9 13 16 9 0 1 15 13 2 13 1 15 13 2 9 15 1 10 9 13 13 2
11 9 9 2 9 13 2 9 13 0 13 2
52 10 9 0 1 15 9 1 9 9 2 1 9 2 1 9 2 1 9 9 13 9 14 1 9 9 13 2 7 9 13 2 9 0 13 2 9 9 13 16 9 7 9 1 9 2 1 9 9 15 9 13 2
13 9 0 2 9 1 9 7 9 1 9 9 13 2
50 3 9 7 9 1 15 9 0 13 2 7 10 9 16 9 14 3 13 16 1 1 10 9 9 9 13 2 9 0 7 0 7 9 1 9 9 1 9 9 13 2 15 1 10 9 13 16 9 13 2
14 9 0 1 9 10 9 1 9 13 16 10 9 13 2
10 9 0 2 9 0 7 0 9 13 2
42 9 13 16 10 9 16 1 9 9 13 2 0 13 2 0 13 2 9 15 0 13 2 9 15 0 13 2 15 15 0 13 2 9 15 0 13 2 16 10 9 13 2
10 9 9 0 2 12 0 1 9 13 2
44 9 0 13 16 9 0 7 9 0 0 1 1 15 9 0 13 2 9 2 9 2 9 2 9 2 9 2 9 2 9 1 9 7 9 1 9 7 9 9 1 15 0 13 2
11 9 9 7 9 16 12 1 9 9 13 2
6 9 13 3 9 13 2
24 10 9 2 9 9 7 9 9 7 9 9 16 13 2 9 10 14 13 2 13 10 9 13 2
13 12 0 1 9 2 9 0 7 0 7 0 13 2
58 9 13 16 10 9 1 9 0 2 9 10 9 0 7 9 13 2 1 9 0 2 9 15 0 1 9 0 13 16 10 9 13 2 1 10 9 13 2 1 9 0 2 1 9 0 7 0 16 13 2 3 9 7 9 9 0 13 2
7 9 9 10 9 3 13 2
13 9 9 7 9 7 9 7 9 10 9 0 13 2
26 10 9 16 13 10 9 0 7 10 9 0 14 3 1 9 1 10 9 1 9 9 13 2 3 13 2
34 15 9 13 1 15 7 9 1 10 9 16 9 13 9 9 9 0 13 7 9 0 1 10 9 1 9 1 9 10 9 1 9 13 2
25 1 15 9 9 13 7 9 15 7 9 14 1 9 9 0 7 9 9 13 7 0 16 9 13 2
11 9 13 3 13 2 9 1 10 9 13 2
42 15 3 9 4 13 16 15 10 9 1 9 0 9 13 7 15 1 9 9 0 1 9 13 2 10 3 13 16 3 9 9 15 14 16 13 7 9 15 14 16 13 2
79 3 15 3 16 15 15 14 1 9 0 9 13 2 3 9 13 2 7 16 1 10 9 16 1 10 9 13 2 1 10 9 16 1 9 0 13 2 9 13 2 10 9 13 16 10 9 3 1 9 13 1 10 9 9 13 7 10 9 3 9 9 13 7 9 15 14 13 2 10 9 13 13 13 16 9 13 3 13 2
10 6 2 9 13 2 9 9 14 13 2
7 3 9 13 3 13 2 2
18 9 16 13 2 3 12 9 9 0 14 1 9 15 15 3 13 2 2
13 9 14 16 13 2 3 9 1 15 9 13 2 2
13 9 3 13 3 13 2 3 16 3 13 3 13 2
103 10 9 16 1 9 13 7 9 9 0 13 2 4 16 3 0 13 2 16 15 1 15 14 0 13 13 2 15 14 0 13 13 2 9 0 13 2 16 1 15 9 13 2 1 15 9 13 2 9 9 4 13 2 16 15 9 2 9 7 9 7 9 1 9 13 2 1 9 10 9 9 4 9 13 2 9 0 13 7 1 9 13 2 4 9 1 9 9 0 14 9 13 7 12 9 0 13 16 4 1 9 13 2
3 9 15 2
11 9 12 9 0 13 2 12 9 0 13 2
28 12 9 9 16 9 9 0 13 2 0 13 2 7 1 9 9 2 9 4 9 0 13 2 10 9 3 13 2
67 10 9 1 15 13 16 10 9 16 9 13 7 9 0 13 13 2 9 0 13 7 3 9 0 2 9 0 2 9 0 2 9 0 2 1 9 7 1 9 10 9 1 9 1 9 13 7 3 13 2 16 10 9 4 1 9 7 1 9 1 9 9 15 15 9 13 2
24 9 2 0 13 2 9 2 9 13 2 7 9 16 0 13 2 4 9 13 7 1 9 13 2
6 3 10 9 1 13 2
17 10 9 16 13 4 1 9 13 2 10 9 1 9 1 3 13 2
13 9 2 9 0 13 7 4 3 0 7 0 13 2
19 1 9 7 1 9 0 9 2 9 1 9 4 9 13 7 9 9 13 2
50 1 9 0 7 0 9 2 1 9 0 2 1 9 2 1 9 9 7 9 9 2 3 1 9 0 2 4 9 0 7 0 7 0 2 3 9 0 2 9 0 2 9 0 7 9 0 14 9 13 2
6 9 2 10 9 13 2
30 1 9 10 9 3 13 7 9 14 1 9 13 2 10 9 9 2 12 9 0 7 9 1 9 13 7 0 16 13 2
38 10 9 2 0 16 13 2 16 10 12 9 2 12 9 12 9 2 16 9 1 9 9 13 2 4 13 16 1 9 0 2 9 7 9 9 13 13 2
10 3 2 12 9 1 10 9 0 13 2
28 15 9 15 13 16 9 0 1 10 9 9 13 2 7 7 9 16 1 9 9 0 0 13 2 3 9 13 2
31 12 9 1 10 9 0 13 2 12 15 16 9 16 9 1 9 15 0 13 13 2 1 9 13 7 3 1 15 9 13 2
80 0 15 7 10 9 14 1 7 13 2 10 9 13 16 12 1 9 0 7 0 7 0 9 13 2 7 1 9 9 13 2 7 1 9 9 13 2 7 1 9 9 9 13 2 7 1 9 9 7 9 9 13 2 1 9 9 7 9 9 9 13 2 16 10 9 13 2 9 3 9 13 2 4 1 15 9 9 9 13 2
26 0 1 15 2 9 0 13 16 4 1 10 10 9 9 13 7 15 15 14 1 9 7 9 9 13 2
8 9 0 2 9 1 9 13 2
26 9 7 9 7 9 9 13 16 9 7 9 7 9 1 9 13 7 9 9 15 15 14 1 9 13 2
7 9 2 9 15 9 13 2
15 16 13 9 1 9 13 2 4 9 7 9 1 9 13 2
20 10 9 1 9 2 15 13 16 15 1 9 9 1 15 1 9 0 9 13 2
18 16 9 2 9 7 9 1 9 9 9 13 2 9 0 9 4 13 2
7 15 2 10 9 0 13 2
26 1 9 9 13 2 1 9 9 0 13 2 1 9 9 9 7 9 1 9 14 1 9 0 9 13 2
25 3 1 9 0 1 9 9 13 16 1 15 1 10 12 9 9 13 2 7 1 10 0 9 13 2
67 15 13 1 9 9 13 2 7 1 9 7 9 9 0 13 2 15 16 3 2 1 9 7 9 9 0 13 1 9 7 9 9 13 7 1 9 9 9 0 14 13 2 3 15 7 0 13 0 16 13 7 9 12 15 2 9 9 13 2 9 9 7 9 7 9 13 2
47 1 9 9 2 12 1 9 9 7 9 9 0 9 0 13 2 12 1 9 9 9 1 9 9 9 0 9 13 2 12 1 9 9 9 0 0 13 2 12 1 9 9 9 0 0 13 2
52 3 10 9 0 13 2 9 16 13 2 0 15 15 13 16 15 1 15 9 9 13 2 7 16 12 9 1 12 9 9 0 13 2 12 9 1 12 9 0 9 0 13 2 3 0 2 15 13 0 16 13 2
23 10 9 16 1 9 1 9 9 13 2 15 0 10 9 13 16 1 9 7 9 9 13 2
21 10 9 16 1 9 7 9 9 13 2 0 10 9 13 16 1 9 9 0 13 2
12 3 9 1 9 13 2 7 10 9 0 13 2
76 0 13 10 9 16 1 9 0 9 13 2 1 10 9 16 1 9 0 9 13 2 13 16 15 1 9 9 7 9 13 2 7 10 9 16 1 9 9 0 13 2 1 10 9 16 1 9 0 9 13 2 7 1 9 9 0 13 2 13 15 1 9 7 9 7 1 9 9 9 13 2 9 14 9 13 2
26 15 1 9 13 7 7 0 13 3 13 2 7 9 13 7 0 13 2 4 15 14 9 7 0 13 2
48 16 7 9 14 16 9 7 9 1 9 10 9 13 15 1 9 0 0 13 2 15 16 3 12 9 0 1 12 9 9 13 7 0 1 9 0 9 13 2 3 9 0 13 2 9 4 13 2
53 9 16 1 15 9 13 2 12 9 0 7 12 9 0 13 2 13 1 7 12 9 0 14 9 13 2 9 0 9 0 7 0 14 9 13 2 1 3 3 12 9 9 13 2 12 9 2 16 12 9 12 9 2
18 16 10 12 9 12 9 3 9 13 2 10 9 3 7 3 4 13 2
65 3 10 9 16 13 15 10 9 14 1 9 9 13 7 1 15 9 9 14 0 9 15 15 13 2 9 13 16 1 9 0 7 1 9 15 9 13 13 2 7 15 15 13 16 12 9 0 0 1 9 9 13 13 16 4 9 9 7 9 15 9 14 3 13 2
4 3 9 13 2
11 1 15 7 9 9 7 9 0 14 13 2
42 15 0 13 9 0 13 2 7 1 9 0 13 7 4 15 14 16 9 9 7 9 7 9 7 9 0 13 2 3 9 13 2 0 13 9 13 7 9 16 13 13 2
6 3 2 4 9 13 2
5 3 4 0 13 2
17 1 15 7 16 15 1 9 9 13 2 9 9 1 9 4 13 2
46 15 16 1 9 15 15 13 2 1 9 9 15 15 13 2 1 9 9 15 15 13 2 1 9 9 13 2 1 9 9 9 13 2 10 9 10 9 0 1 9 10 9 9 4 13 2
22 16 16 1 9 13 2 1 15 7 0 13 9 15 14 9 13 2 15 15 0 13 2
4 3 9 13 2
15 1 15 7 16 9 13 7 9 14 13 2 9 4 13 2
39 4 9 13 2 16 9 14 13 2 16 9 7 9 14 13 2 16 4 1 1 9 15 14 16 9 9 7 9 15 13 2 15 14 9 13 7 9 13 2
21 10 9 7 9 0 2 1 9 0 9 13 13 2 15 10 9 13 16 0 13 2
34 3 3 1 9 0 15 2 10 9 16 15 9 13 16 15 0 1 9 9 13 2 15 1 9 7 9 9 13 15 14 0 9 13 2
37 16 15 14 0 1 15 16 3 9 13 2 9 13 2 9 12 9 3 3 0 13 2 7 0 16 13 2 13 1 7 9 13 7 0 15 13 2
41 0 15 13 16 15 1 15 9 0 9 13 13 7 9 13 2 7 3 16 16 13 7 9 1 10 9 2 9 16 1 10 9 9 13 2 16 1 15 9 13 2
16 9 1 10 9 9 13 2 0 15 13 16 1 9 9 13 2
32 10 12 9 4 0 13 2 3 10 9 0 0 9 7 9 13 2 3 9 0 0 9 7 9 1 9 7 9 9 9 13 2
46 16 12 9 10 9 14 13 13 2 10 9 9 13 9 13 16 1 10 9 16 1 9 7 0 13 2 9 15 15 14 1 9 9 7 9 16 9 1 15 1 9 13 2 3 13 2
37 3 12 9 2 9 13 1 15 7 12 9 7 12 9 2 15 15 9 13 7 0 9 13 2 7 9 0 1 15 16 9 13 2 15 3 13 2
15 15 9 9 13 2 1 10 12 9 0 13 9 9 13 2
39 3 12 9 1 10 12 9 9 13 2 1 10 9 1 9 9 13 7 1 10 9 9 9 13 2 3 1 9 0 16 9 13 7 13 9 0 14 13 2
25 15 1 9 9 2 1 9 9 2 1 9 9 2 1 9 9 2 13 0 9 13 7 9 13 2
10 15 0 13 1 9 0 9 9 13 2
91 16 10 9 9 0 7 0 1 9 0 9 9 13 2 3 0 13 2 16 9 7 9 7 9 1 9 0 13 2 4 9 9 0 13 2 7 1 15 0 15 13 16 13 1 9 0 9 13 2 9 9 2 9 9 2 9 9 2 9 9 0 9 14 9 13 7 1 9 13 2 10 9 9 13 16 1 9 9 7 9 7 9 9 9 4 9 13 2 16 9 2
80 3 7 9 7 9 0 9 0 9 1 9 9 13 2 15 1 1 9 15 13 7 9 0 14 16 9 13 7 1 9 0 13 9 13 2 15 10 9 13 16 9 0 9 3 1 15 2 9 15 14 1 9 7 1 9 13 7 9 0 14 13 2 15 13 2 15 16 9 15 14 9 13 7 13 3 9 0 9 13 2
25 16 9 13 1 9 9 1 9 9 2 9 1 9 13 2 0 13 16 9 1 9 15 3 13 2
14 9 1 9 15 2 16 9 9 0 1 9 3 0 2
9 3 15 15 1 15 14 16 13 2
101 3 15 16 1 9 7 9 9 0 13 16 1 10 9 13 7 13 7 9 0 3 13 2 3 16 13 15 15 14 1 9 9 9 9 13 7 3 4 9 0 13 7 9 0 13 7 9 9 7 9 7 9 13 2 10 9 16 9 9 7 9 9 13 16 0 1 12 9 1 10 9 9 13 7 12 9 9 1 10 12 9 13 2 3 10 9 16 1 15 9 1 10 9 9 13 2 13 9 9 13 2
7 10 9 9 15 13 2 2
8 10 9 2 16 10 9 0 2
45 16 3 16 15 9 9 9 9 14 9 13 2 13 13 7 9 15 14 9 13 2 9 13 9 0 1 9 9 13 7 0 16 9 9 7 9 7 9 9 9 14 1 9 13 2
80 12 9 16 9 13 16 9 10 9 13 2 7 1 0 9 2 16 15 3 1 9 2 9 13 16 1 9 9 1 9 9 1 9 9 9 13 2 15 9 9 14 13 7 9 9 14 9 13 2 9 9 1 10 9 16 13 2 7 3 9 1 9 0 2 1 9 0 7 1 9 0 13 2 0 1 10 9 0 13 2
17 9 9 16 12 9 1 9 13 9 14 9 13 7 1 9 13 2
21 16 9 1 9 10 9 13 2 10 9 2 3 9 7 9 14 1 9 9 13 2
34 15 16 9 1 9 13 2 3 9 1 9 16 13 2 7 1 1 9 9 13 16 3 1 9 4 9 13 7 1 15 9 9 13 2
37 3 9 1 9 13 2 7 1 1 9 9 13 16 9 9 1 9 0 2 9 9 7 9 9 9 7 9 0 7 9 1 0 7 9 14 13 2
35 0 13 16 15 0 13 2 15 9 10 9 13 16 9 14 0 13 7 0 1 9 13 2 3 2 15 0 13 2 15 0 7 9 13 2
31 9 0 9 3 1 15 1 10 9 9 9 9 9 7 9 14 0 13 2 7 9 15 0 13 16 3 13 9 7 9 2
24 6 2 15 9 2 15 9 7 9 7 9 14 0 13 2 9 0 4 9 15 14 9 13 2
21 9 1 9 13 7 1 9 13 2 9 4 13 16 15 1 9 10 9 9 13 2
33 9 9 13 2 15 14 16 13 2 15 16 16 13 2 15 0 1 10 9 7 9 13 2 10 9 13 2 3 1 15 9 13 2
21 10 9 0 7 0 16 9 9 9 14 1 9 0 13 2 15 13 3 9 13 2
49 9 1 10 9 2 10 9 14 1 9 13 13 2 3 1 15 9 13 2 7 13 16 9 1 15 0 13 2 15 16 13 2 12 0 13 2 0 16 9 15 13 2 16 1 9 15 0 13 2
42 13 1 7 7 10 9 0 1 9 0 13 7 10 9 1 9 9 1 9 9 13 2 9 15 0 13 1 9 9 0 13 2 7 4 13 10 9 0 14 0 13 2
11 9 15 9 1 9 15 13 2 9 0 2
2 9 2
9 13 9 0 7 0 14 9 13 2
11 9 0 1 9 10 9 0 9 0 13 2
29 0 13 1 9 0 2 12 9 1 9 1 12 9 2 12 9 16 1 12 9 0 0 13 7 1 9 0 13 2
41 9 13 10 9 16 10 9 1 9 0 13 2 12 9 13 2 10 9 16 10 9 0 0 13 2 9 0 13 2 3 2 15 9 7 9 0 7 9 0 13 2
9 9 1 9 0 1 10 9 13 2
56 9 10 9 14 9 13 2 10 9 14 1 10 9 9 3 9 2 3 9 2 3 9 0 2 10 9 16 9 9 13 13 16 13 1 9 9 0 13 10 9 14 1 9 7 9 7 9 7 9 9 16 13 2 9 13 2
5 9 1 9 13 2
16 10 12 9 16 1 1 9 9 13 2 9 0 14 9 13 2
28 16 9 1 15 15 14 0 13 7 9 0 1 7 0 13 2 16 9 15 14 1 10 9 0 7 0 13 2
44 13 2 9 15 16 9 7 9 1 9 9 3 9 13 2 12 9 13 2 7 10 9 16 10 9 0 1 9 2 9 15 14 1 1 0 3 9 13 2 12 9 0 13 2
49 15 1 9 9 2 10 9 16 1 1 9 9 13 16 9 9 16 13 1 7 7 9 7 9 13 13 2 9 7 9 7 9 7 9 7 9 15 9 13 2 15 4 1 15 9 13 7 13 2
35 16 9 1 9 13 7 9 13 2 15 13 16 9 0 9 14 9 13 13 7 9 0 9 14 2 1 15 9 13 13 2 9 15 13 2
30 10 9 16 1 9 0 9 9 13 2 15 13 3 9 14 13 13 2 16 3 13 13 2 4 9 13 2 9 13 2
96 15 12 9 13 2 7 9 9 0 2 3 1 9 9 13 2 9 0 4 9 15 14 0 13 2 4 3 1 1 10 9 16 1 9 0 13 2 1 9 0 13 2 1 9 9 0 13 2 1 9 0 1 10 9 0 13 2 9 7 9 15 14 0 13 2 10 9 1 1 9 16 16 3 13 2 7 1 9 9 7 1 9 9 3 9 13 9 7 9 4 9 15 14 0 13 2
23 13 9 7 9 7 9 13 2 7 9 15 14 0 13 2 15 9 15 1 9 0 13 2
8 3 9 9 9 15 0 13 2
13 9 15 2 9 1 9 9 13 2 9 9 13 2
63 15 10 9 16 9 13 16 3 3 9 1 10 9 0 7 0 7 0 7 0 7 0 7 0 7 0 7 0 13 2 15 16 9 13 2 1 10 9 0 13 2 1 9 13 16 13 2 1 9 13 16 13 2 4 13 16 15 9 13 2 9 13 2
87 3 9 9 9 1 10 9 2 12 9 3 0 7 0 13 2 13 9 14 1 9 10 9 0 7 0 13 2 13 9 14 1 9 0 13 2 13 9 14 1 9 0 13 2 13 9 14 1 9 0 16 1 9 0 13 1 9 9 2 1 9 9 2 1 9 9 0 13 2 13 1 9 9 13 7 9 9 13 2 13 9 0 1 9 0 13 2
15 15 16 9 13 15 1 9 9 7 9 13 2 15 13 2
35 15 16 1 10 9 13 2 3 2 9 9 13 2 9 13 7 13 9 14 13 7 0 16 13 7 1 9 9 9 15 15 14 9 13 2
16 9 9 9 13 16 9 13 2 4 3 9 1 15 9 13 2
20 15 9 16 1 9 0 9 9 13 2 1 9 7 9 0 10 9 9 13 2
26 13 10 9 16 13 10 9 14 9 13 2 10 9 13 16 15 1 9 0 13 7 9 13 16 13 2
10 3 3 9 9 9 0 7 0 13 2
30 1 9 12 9 9 16 9 0 1 9 13 7 9 3 12 9 13 16 1 15 7 9 7 9 7 9 15 0 13 2
21 16 10 9 0 7 0 7 0 7 0 0 13 16 9 13 7 13 16 3 13 2
43 16 9 9 1 9 9 7 9 15 1 15 2 3 1 9 9 0 9 15 16 9 9 9 13 2 3 9 1 1 9 7 9 0 0 16 15 16 10 9 14 13 13 2
95 3 3 15 13 9 9 9 9 2 9 0 1 9 0 7 9 0 0 7 0 13 7 3 3 15 7 3 9 0 0 7 9 16 1 9 7 9 1 1 9 9 2 3 9 9 4 9 13 2 3 9 14 9 13 7 15 16 1 9 1 1 9 9 9 9 9 1 9 13 2 3 3 9 9 9 9 10 9 7 9 7 9 7 9 14 13 7 3 1 9 9 9 9 13 2
4 9 0 13 2
66 9 15 13 16 9 9 3 1 1 9 9 9 13 7 1 1 15 1 9 9 7 9 9 0 16 13 7 9 10 9 7 9 14 3 12 9 12 9 1 15 7 3 13 7 1 10 9 1 9 15 9 0 2 1 9 9 9 9 13 7 9 1 9 15 13 2
29 3 9 9 0 7 9 0 9 0 9 12 16 13 9 10 9 14 1 9 0 9 0 13 7 1 9 9 13 2
25 9 15 9 13 16 13 1 9 9 13 2 16 9 1 9 9 0 0 0 7 0 9 13 13 2
44 9 16 3 7 7 3 13 7 13 16 9 0 7 0 1 9 0 7 0 13 2 7 9 9 0 1 9 0 7 0 13 7 9 9 0 1 0 0 1 9 0 4 13 2
40 9 13 9 7 9 0 1 1 9 9 1 9 9 7 9 7 9 7 9 7 9 7 7 9 16 9 7 9 13 13 7 10 15 9 9 12 9 0 13 2
17 3 9 0 9 1 9 15 13 16 9 14 1 10 9 0 13 2
21 0 13 16 9 9 0 1 10 9 16 1 9 12 9 9 9 13 16 3 13 2
42 1 9 0 0 13 2 7 4 1 9 7 1 10 9 16 13 6 1 9 1 9 15 12 9 9 13 16 9 0 13 2 9 0 1 9 7 9 0 1 9 13 2
23 9 9 9 9 1 9 14 1 9 0 15 13 13 7 13 10 9 14 9 15 9 13 2
31 9 9 7 9 0 9 14 1 9 9 9 1 9 7 9 0 13 13 7 13 10 9 7 9 14 1 9 15 9 13 2
30 3 10 9 16 9 9 13 16 3 13 2 1 12 9 0 13 2 7 10 9 10 9 13 16 1 9 9 13 13 2
24 13 16 16 9 7 9 7 7 10 9 9 0 13 13 2 15 3 1 1 9 9 9 13 2
18 1 10 9 9 9 13 15 1 12 9 0 2 0 7 0 9 13 2
21 9 12 1 10 12 9 9 9 15 13 7 3 1 10 12 13 0 7 0 13 2
11 15 0 13 16 9 9 15 9 0 13 2
12 10 9 16 9 1 9 7 9 0 0 13 2
19 3 16 3 1 9 7 9 0 13 2 7 9 0 16 1 15 9 13 2
42 12 16 13 12 9 9 7 9 14 0 13 7 1 9 9 0 9 7 9 7 9 7 9 9 0 2 12 9 1 12 9 2 1 9 9 0 1 9 0 13 13 2
13 16 1 9 9 15 14 9 13 2 13 3 13 2
8 9 0 14 1 3 9 13 2
11 9 0 12 12 9 1 9 9 9 13 2
10 9 9 0 1 9 0 0 13 13 2
14 9 9 0 4 1 9 1 9 0 7 0 9 13 2
12 9 9 1 9 9 0 7 0 9 0 13 2
18 9 9 1 9 0 9 7 9 3 9 0 9 0 7 0 13 13 2
9 9 9 1 9 9 9 9 13 2
12 9 9 1 9 3 1 9 0 0 4 13 2
12 9 13 9 0 9 0 9 7 9 9 13 2
18 9 9 9 1 9 0 7 9 9 15 1 9 0 1 9 9 13 2
19 9 1 9 12 9 12 0 0 16 9 10 9 0 1 15 13 9 13 2
21 9 9 9 1 1 9 9 1 9 9 9 9 9 9 0 1 9 14 9 13 2
15 9 9 0 3 9 0 2 9 0 14 3 0 13 13 2
6 9 0 9 9 13 2
24 9 9 9 9 9 7 9 0 7 9 9 9 9 1 9 9 9 9 9 9 9 9 13 2
27 9 9 1 10 9 9 0 9 9 9 14 1 9 9 0 7 9 1 9 9 0 1 9 9 9 13 2
35 1 9 9 9 1 9 9 9 9 9 9 9 9 9 2 9 9 9 9 0 9 2 9 7 9 9 7 9 9 9 9 16 9 13 2
27 9 9 9 9 9 9 9 1 12 9 0 9 13 16 0 9 12 9 9 1 9 0 9 9 4 13 2
30 1 9 9 9 2 15 1 9 13 16 9 9 13 1 9 9 2 9 9 1 9 14 1 12 12 9 9 9 13 2
23 9 0 13 15 1 9 9 9 0 13 7 1 12 9 0 9 0 1 10 9 0 13 2
61 9 9 9 9 9 1 9 1 9 9 9 9 0 9 2 9 9 14 9 0 7 3 0 13 7 9 13 2 9 0 4 1 9 9 0 7 9 0 15 2 1 9 12 9 0 2 0 2 0 7 0 2 9 0 15 14 9 7 9 13 2
88 1 9 9 9 0 9 9 1 9 1 9 0 9 0 9 1 9 9 2 9 7 9 9 0 7 0 1 9 2 9 1 9 7 9 9 0 2 0 7 0 9 0 14 0 13 7 9 13 2 10 9 1 9 1 9 9 1 9 9 0 9 2 9 9 0 9 9 14 1 9 9 0 9 0 7 0 1 10 9 0 7 9 10 9 2 0 13 2
56 15 2 9 9 0 14 9 7 9 9 0 9 13 7 1 9 1 9 0 9 13 2 9 0 2 9 9 7 9 9 2 9 7 9 13 16 1 15 9 1 9 9 7 9 0 9 9 2 9 0 7 0 13 7 13 2
67 9 9 9 2 1 9 1 9 0 9 0 1 9 9 13 2 1 9 0 10 9 2 9 1 9 9 13 13 7 3 16 4 1 9 1 9 0 2 0 7 0 1 9 1 9 9 7 9 0 1 9 9 1 9 9 9 1 9 9 0 9 9 13 7 9 13 2
74 9 9 16 1 9 9 9 7 9 0 9 0 9 2 9 1 9 14 9 9 0 7 9 9 9 13 7 13 2 9 9 0 7 1 9 0 9 9 1 9 9 9 7 9 1 9 1 9 0 7 0 2 4 1 9 0 9 7 9 3 9 0 2 0 0 2 0 2 0 7 0 13 13 2
35 9 9 16 1 9 9 9 0 9 0 9 2 9 0 9 14 0 1 9 0 1 9 9 13 7 1 9 9 0 9 0 9 9 13 2
36 15 1 9 1 9 9 9 9 0 9 1 9 1 9 0 9 13 2 9 7 9 9 9 0 9 1 9 9 1 9 9 9 9 0 13 2
27 9 9 16 9 1 9 9 7 9 0 9 0 14 0 13 7 1 9 0 7 0 9 1 9 9 13 2
23 9 9 3 9 13 2 9 10 9 1 9 9 9 9 9 9 9 12 9 9 4 13 2
63 9 9 9 9 9 9 1 9 1 9 9 0 9 1 9 10 9 9 13 2 9 9 9 9 3 1 12 9 0 7 0 1 10 9 13 16 3 1 9 9 9 2 1 9 9 10 9 9 15 14 1 9 9 9 13 7 1 9 9 0 9 13 2
61 9 9 9 1 9 1 9 1 0 9 9 9 9 9 13 2 1 9 15 9 0 9 0 9 9 13 16 1 9 9 0 13 10 9 14 1 9 9 13 7 9 0 9 9 9 1 10 9 7 9 7 9 0 9 9 9 14 0 13 13 2
21 9 9 9 1 9 0 1 9 9 1 9 12 9 9 13 2 9 9 9 13 2
34 9 9 9 9 9 9 9 9 9 1 9 9 1 9 9 13 1 9 9 9 9 9 9 9 14 1 9 0 9 7 9 9 13 2
30 1 10 9 16 9 9 9 1 9 0 9 9 13 2 9 9 9 7 9 9 0 1 9 9 0 0 9 13 13 2
53 9 9 9 1 9 15 13 13 2 1 9 9 9 0 7 9 9 0 1 9 7 9 1 9 2 3 9 9 0 7 0 9 0 13 16 9 15 2 9 9 0 7 0 10 2 9 7 9 9 9 13 13 2
38 9 9 9 9 0 0 1 9 1 9 9 9 0 2 9 9 9 9 2 9 9 9 0 2 9 9 9 9 2 9 0 9 7 10 9 0 13 2
14 9 9 10 9 2 9 9 14 1 9 0 9 13 2
16 12 9 9 9 9 3 13 2 9 9 9 9 3 0 13 2
25 9 9 13 2 3 1 1 9 1 9 16 1 9 15 1 9 9 13 2 9 0 9 4 13 2
24 15 0 13 2 9 9 3 1 9 9 0 1 9 9 9 2 1 9 9 9 9 0 13 2
42 9 9 13 2 9 9 1 9 9 9 15 1 9 9 9 9 1 9 0 9 13 7 0 13 9 9 1 9 1 9 9 16 1 3 9 13 9 13 2 9 13 2
52 15 9 0 14 1 12 9 9 13 7 13 2 3 9 16 1 15 9 13 9 13 7 3 1 15 7 1 9 13 2 9 13 13 9 1 9 0 16 16 1 1 15 9 13 2 1 9 0 2 9 13 2
34 9 9 9 9 13 2 10 9 9 13 9 9 1 0 9 0 9 9 2 9 9 14 1 9 13 7 9 15 14 1 9 9 13 2
44 15 1 9 1 10 9 16 16 9 9 1 9 7 7 9 9 9 9 9 9 13 2 13 2 9 9 13 7 15 13 9 9 13 7 10 9 9 1 9 9 9 9 13 2
45 9 1 9 9 9 9 9 9 7 9 9 13 2 1 10 9 1 9 9 9 9 9 13 7 10 12 9 13 16 1 10 9 9 1 9 0 9 0 13 7 9 7 9 13 2
5 9 9 0 13 2
37 9 9 1 9 9 13 2 9 9 9 9 9 9 9 1 9 9 0 0 1 9 9 9 9 9 13 7 3 1 9 9 0 9 14 9 13 2
56 1 10 9 16 9 9 9 13 2 13 13 2 1 1 9 10 9 3 0 1 9 0 7 1 1 9 0 1 9 0 2 1 9 9 9 2 9 9 9 1 9 0 9 9 2 3 1 9 3 1 9 9 9 0 13 2
32 1 9 9 9 13 2 3 2 1 9 0 2 3 1 9 0 2 3 9 9 9 13 13 7 9 9 9 9 14 9 13 2
23 9 9 9 9 9 0 9 9 1 9 9 9 9 7 9 9 9 0 9 7 9 13 2
43 9 9 1 10 9 1 9 1 9 0 9 9 1 9 9 9 9 9 0 9 13 2 9 9 0 1 10 9 1 12 9 3 0 1 12 9 0 1 9 0 9 13 2
48 9 1 9 1 9 9 9 0 1 12 9 0 13 2 9 0 1 10 9 1 7 0 13 7 10 9 13 1 9 0 7 0 9 7 1 9 1 9 2 9 7 9 9 0 9 13 13 2
27 9 9 9 0 1 9 1 9 10 9 1 9 9 9 9 9 13 16 1 9 2 9 1 9 9 13 2
33 9 9 9 9 9 0 7 9 0 14 0 9 13 7 13 2 10 9 1 9 9 9 16 9 0 13 7 9 0 14 13 13 2
15 9 9 9 0 1 9 1 9 9 0 10 9 9 13 2
57 9 9 16 1 10 9 1 9 10 9 16 1 9 9 9 9 1 9 9 0 10 9 1 9 0 9 9 13 13 13 2 9 3 9 7 9 0 9 0 1 9 0 16 1 0 9 9 0 13 1 9 9 9 9 4 13 2
42 9 9 9 0 1 9 9 0 7 9 1 9 9 10 9 9 13 7 13 2 10 9 3 9 0 1 9 0 7 1 9 1 9 0 0 1 9 9 9 0 13 2
4 3 0 13 2
9 9 0 9 0 9 3 0 13 2
30 9 1 9 16 9 9 9 14 13 2 3 13 16 1 9 2 9 7 9 13 7 9 15 14 1 3 9 0 13 2
51 1 9 9 1 9 7 9 16 1 9 9 9 13 2 3 13 16 9 9 9 7 9 1 9 9 1 9 9 0 7 9 9 14 13 3 7 1 3 10 9 9 9 7 9 2 15 14 9 4 13 2
33 1 9 0 2 15 9 7 9 1 1 9 9 14 1 9 9 7 9 1 9 1 13 16 15 3 9 9 7 9 3 9 13 2
35 3 9 7 9 1 9 10 9 0 9 2 1 9 13 7 10 9 9 1 10 9 2 1 9 0 9 9 2 3 1 9 9 4 13 2
50 9 9 13 9 16 1 0 9 16 1 9 9 3 2 9 13 2 3 1 9 0 7 0 1 9 10 9 9 1 9 7 0 9 9 9 0 1 15 2 9 13 7 1 9 9 15 9 13 2 2
67 9 0 15 16 9 9 1 10 12 9 4 3 1 9 10 12 9 1 9 7 9 0 15 0 13 13 7 1 10 9 0 13 13 16 3 10 12 9 1 0 9 7 9 3 2 0 1 9 1 9 7 9 7 9 0 9 14 1 9 15 9 0 15 13 9 13 2
40 9 0 10 9 15 13 16 9 0 9 9 2 16 9 16 1 9 7 9 13 2 7 3 9 9 0 13 16 1 3 12 1 9 7 9 16 9 9 13 2
78 0 9 9 1 9 10 9 0 7 0 15 13 16 3 1 10 3 2 9 1 9 0 0 9 13 7 9 13 16 1 12 9 0 13 9 0 0 0 9 14 1 12 9 0 7 0 2 9 13 7 9 13 16 9 1 15 0 13 7 7 1 15 13 7 10 9 9 1 15 13 2 3 9 9 9 9 13 2
49 10 9 0 7 0 1 9 0 9 7 9 1 10 9 9 0 9 9 0 1 9 0 0 9 13 7 3 1 9 9 2 9 2 9 7 3 9 10 12 1 12 9 0 13 16 13 13 13 2
68 16 9 0 9 15 1 9 0 7 9 9 7 9 7 9 7 9 0 7 9 7 9 0 0 14 13 16 9 0 13 7 3 0 13 2 1 3 9 9 9 13 13 7 4 1 9 3 9 0 9 1 9 14 1 9 0 7 0 15 9 7 1 9 9 7 9 13 2
14 1 9 3 0 1 12 9 1 9 9 9 13 13 2
57 7 3 9 9 9 9 14 16 1 15 9 0 9 9 9 14 1 15 9 13 14 9 13 13 2 16 1 3 9 16 9 9 1 15 13 7 1 9 15 9 13 7 3 9 9 14 13 1 9 9 7 9 9 9 4 13 2
66 16 1 9 0 9 1 9 9 9 12 9 7 3 9 0 7 9 9 9 13 13 16 3 9 7 9 3 9 13 2 1 3 9 1 9 1 9 13 2 1 9 10 9 3 9 9 1 9 9 13 7 9 9 3 9 0 9 16 9 0 7 0 15 14 13 2
28 1 9 7 9 9 9 3 0 7 9 9 0 13 4 1 9 9 9 13 16 9 0 9 1 9 9 13 2
28 12 1 9 13 9 9 9 1 9 1 9 0 9 0 9 1 9 14 0 7 0 1 9 9 0 13 13 2
16 9 1 9 0 3 1 0 9 9 9 1 9 7 9 13 2
45 16 9 7 7 10 9 0 9 1 9 15 1 12 9 9 13 2 9 9 9 1 9 9 1 9 9 13 13 7 15 9 0 15 1 9 9 9 0 15 14 1 9 4 13 2
28 9 3 1 9 9 13 7 10 9 16 13 9 9 15 4 13 7 0 13 16 1 9 9 1 9 9 13 2
20 1 10 9 9 1 9 9 1 9 7 3 9 0 9 1 9 9 0 13 2
19 12 3 9 0 7 9 9 1 9 3 1 9 0 9 9 14 0 13 2
32 1 9 1 10 9 4 3 1 9 9 3 9 9 0 9 13 16 9 9 9 7 9 9 9 9 1 9 9 1 9 13 2
50 16 9 9 13 16 9 0 1 12 9 0 2 9 9 7 9 14 13 7 9 7 9 9 15 14 1 9 1 9 13 1 15 9 13 7 10 9 15 9 0 9 7 9 9 14 1 9 4 13 2
34 16 9 9 13 16 12 9 0 1 9 9 7 9 9 13 7 0 1 9 13 15 14 1 9 0 7 9 0 9 13 16 9 13 2
35 9 7 9 9 9 1 9 0 15 1 9 2 9 2 9 7 9 2 2 13 13 2 9 1 12 9 0 1 9 0 15 9 0 13 2
38 3 1 9 9 9 1 9 1 9 2 9 0 0 9 0 13 7 7 3 16 9 0 0 13 4 1 9 0 9 0 14 1 3 1 15 9 13 2
36 9 0 1 0 9 0 1 9 16 9 1 9 9 0 9 15 13 2 3 9 0 13 16 9 9 1 0 9 1 9 9 15 1 9 13 2
26 9 1 9 9 0 16 1 9 1 1 9 1 9 9 9 0 13 2 9 0 14 1 9 13 13 2
34 15 7 9 9 1 9 15 1 3 9 13 13 2 9 9 7 0 1 9 7 9 0 13 16 9 1 10 9 1 9 0 9 13 2
41 7 3 1 9 13 15 1 9 9 9 1 9 0 9 0 16 3 1 9 9 9 1 9 9 0 3 1 9 0 1 9 9 9 13 2 1 9 15 9 13 2
49 10 9 1 9 7 9 9 0 15 7 9 9 1 10 9 0 12 9 0 13 7 15 15 16 9 13 2 9 0 15 9 14 1 9 9 0 3 13 7 1 9 12 9 0 0 9 13 13 2
40 16 15 9 9 9 1 9 9 7 9 13 7 10 9 16 9 13 0 13 9 0 14 1 9 0 7 9 9 15 3 13 7 1 9 12 9 0 9 13 2
33 1 9 0 2 9 3 9 1 15 13 2 9 9 12 9 1 9 12 9 0 3 9 10 9 0 1 9 12 9 7 9 13 2
29 7 9 0 1 10 9 0 13 16 9 0 1 9 0 7 0 1 9 9 10 9 0 1 9 14 1 9 13 2
68 9 1 9 9 0 13 13 1 9 12 9 0 16 1 9 1 9 0 9 0 13 2 9 13 7 10 9 7 9 0 15 13 16 13 1 12 9 9 9 9 14 9 13 7 1 9 0 2 1 9 12 9 0 0 9 9 0 1 9 14 1 9 9 9 1 9 13 2
25 3 9 9 1 9 9 0 15 13 16 9 13 2 1 9 9 13 2 9 0 1 9 0 13 2
20 3 10 9 1 9 9 1 9 9 0 15 13 7 1 1 9 15 9 13 2
49 1 10 9 2 10 9 4 0 13 15 9 9 13 16 15 14 1 9 0 1 9 0 9 13 2 3 15 7 15 0 13 10 9 9 9 12 9 0 14 1 9 13 7 9 0 14 9 13 2
55 1 9 9 0 9 1 9 0 12 9 9 9 9 0 1 9 0 7 0 1 9 1 9 9 7 1 1 12 9 9 0 0 1 9 2 9 13 9 15 14 1 9 9 9 1 9 0 9 9 1 15 9 0 13 2
105 1 9 9 9 9 9 9 0 9 16 9 3 9 9 2 9 9 2 9 9 2 9 7 2 14 0 13 2 9 9 1 9 9 9 15 1 9 0 9 9 0 9 1 9 9 9 1 9 15 16 9 0 9 1 9 9 0 1 9 15 1 9 7 9 9 15 9 13 13 2 9 9 7 9 9 0 13 2 7 3 1 9 9 9 9 9 1 9 9 13 13 2 9 13 9 1 9 9 9 1 9 0 9 13 2
42 1 9 9 9 9 9 9 9 9 9 0 7 9 9 0 9 13 9 0 1 9 9 1 9 10 9 9 9 9 9 9 0 0 9 9 14 1 9 9 9 13 2
22 7 9 9 9 1 1 9 0 9 0 16 1 15 13 16 15 1 9 9 9 13 2
50 1 9 0 1 9 9 9 0 1 9 9 9 9 9 1 9 9 1 9 1 10 9 13 16 1 9 0 9 9 9 1 9 9 0 7 9 16 9 0 13 13 1 9 1 9 0 9 9 13 2
50 1 9 9 0 16 9 13 13 1 9 9 9 2 9 9 2 9 9 9 2 9 0 9 9 2 9 9 9 1 1 1 9 2 9 9 9 9 9 9 1 9 7 0 9 0 0 9 13 13 2
14 9 9 9 9 1 9 0 9 0 1 9 9 13 2
47 12 1 9 0 1 9 9 0 0 1 9 15 13 2 9 9 1 9 0 1 9 1 10 9 7 9 1 9 1 9 9 9 9 9 1 9 3 3 0 9 7 9 15 3 0 13 2
52 9 0 16 1 9 0 1 0 9 9 9 1 9 9 7 9 15 9 13 13 9 13 13 7 9 0 1 1 9 9 9 9 1 9 0 7 0 1 9 9 0 9 1 9 0 9 1 9 0 13 13 2
54 16 9 0 9 9 1 9 7 9 9 7 9 1 15 16 9 0 0 4 15 14 1 9 13 7 1 9 9 9 13 2 9 3 9 9 9 7 1 9 9 9 0 9 14 1 9 3 0 9 0 9 13 13 2
36 1 10 9 0 9 13 16 10 9 9 9 9 1 9 0 9 14 0 9 0 1 9 10 9 13 7 9 1 9 3 9 3 0 9 13 2
50 16 9 0 7 0 2 1 9 0 15 0 9 1 9 0 0 1 9 0 9 13 2 7 15 1 9 9 9 1 9 9 13 2 15 16 2 1 9 9 0 2 9 2 10 9 9 9 0 13 2
7 9 1 9 7 9 13 2
36 9 2 1 10 9 2 12 1 9 9 9 1 9 14 2 3 9 9 0 9 1 9 9 9 1 9 13 16 1 9 0 9 1 9 13 2
27 10 9 0 15 13 16 3 9 14 1 9 3 9 13 7 9 9 1 9 14 1 9 12 9 13 13 2
8 9 9 9 0 1 3 13 2
36 7 3 13 16 1 9 1 9 4 9 9 15 14 1 9 9 1 9 15 0 13 7 15 10 9 13 16 1 9 1 9 9 0 9 13 2
48 1 9 10 9 0 16 2 9 1 9 9 1 9 2 0 9 9 9 9 7 9 9 9 13 16 1 9 15 2 1 9 10 9 2 4 9 9 9 14 1 9 0 1 9 9 9 13 2
23 7 16 4 9 13 16 10 9 2 9 9 0 9 1 9 0 9 15 14 1 9 13 2
29 7 3 16 9 15 13 13 16 9 0 7 0 1 9 7 9 7 9 2 9 15 14 1 10 9 0 13 2 2
54 9 9 1 9 1 0 9 1 9 9 9 0 9 13 7 13 13 2 1 9 7 9 9 0 0 9 0 9 14 9 9 9 0 4 13 2 9 7 9 0 1 1 9 9 9 0 9 2 16 9 1 9 13 2
25 9 7 9 0 9 9 15 14 1 9 9 9 9 13 16 4 9 9 15 14 1 9 9 13 2
43 9 3 9 0 1 9 9 13 2 1 9 1 12 12 9 7 0 9 9 9 1 9 9 9 13 1 9 9 0 1 9 9 1 9 9 12 9 1 9 9 9 13 2
49 9 9 9 9 9 1 9 1 9 2 9 1 0 9 9 9 15 2 9 9 14 0 13 2 1 9 1 9 9 9 0 9 1 9 9 9 0 1 9 1 9 9 9 9 9 1 9 13 2
17 9 10 9 9 9 9 12 9 0 0 0 1 9 0 0 13 2
36 15 1 10 9 1 9 1 9 13 2 16 9 9 1 9 9 0 1 9 9 1 9 12 9 12 2 10 9 3 1 10 9 9 1 13 2
23 15 1 9 1 9 12 1 9 0 9 1 9 9 1 0 9 9 1 9 9 9 13 2
16 1 9 9 10 9 0 9 0 1 9 10 9 14 9 13 2
31 9 1 12 9 12 0 3 0 9 13 16 1 9 9 9 10 9 16 3 1 9 9 13 9 1 9 15 9 1 13 2
24 15 9 9 13 1 9 9 0 4 9 14 3 1 9 0 9 7 9 15 1 9 9 13 2
23 9 0 9 0 0 1 9 9 13 7 10 9 14 1 9 1 9 9 9 1 9 13 2
32 1 9 9 0 9 9 12 9 0 1 9 12 9 13 16 12 1 15 3 1 9 9 0 13 7 0 3 0 9 13 13 2
29 1 9 9 10 9 9 0 4 1 9 9 12 9 0 1 9 9 9 9 1 13 7 10 9 9 9 0 13 2
19 1 9 9 1 3 9 13 9 1 9 3 9 0 7 9 9 14 13 2
24 9 0 1 10 9 13 9 0 1 9 9 9 1 9 0 3 9 2 9 7 9 9 13 2
27 9 0 13 9 9 1 9 10 9 1 9 9 0 16 9 0 13 2 9 0 1 9 10 9 13 13 2
16 1 9 9 10 9 9 9 9 0 1 9 9 9 13 13 2
27 9 9 9 9 9 7 9 0 9 9 1 9 9 13 16 9 9 1 9 3 1 9 0 0 4 13 2
66 9 16 1 9 9 9 9 1 9 9 9 9 9 13 1 1 9 7 9 9 1 9 13 2 0 9 1 1 10 12 9 1 9 14 9 0 9 1 9 9 9 1 9 13 7 1 15 1 9 12 9 9 9 13 16 4 1 9 7 9 0 1 15 9 13 2
31 9 13 2 1 9 9 0 15 9 7 9 0 13 1 9 9 0 16 1 9 9 0 13 9 7 9 15 14 9 13 2
46 15 1 1 10 9 1 1 9 9 0 9 1 9 9 13 2 1 9 0 15 1 9 9 7 9 0 9 13 13 7 15 9 7 9 10 9 1 9 10 9 9 1 10 9 13 2
62 9 9 7 9 0 1 9 9 9 0 7 9 0 13 2 9 15 13 16 1 9 3 9 9 9 7 9 7 9 7 9 9 0 0 13 7 9 1 9 16 9 7 9 1 15 3 9 7 9 9 7 9 10 12 9 0 13 1 3 0 13 2
65 15 1 1 9 9 9 9 13 2 9 9 7 9 0 1 1 9 0 7 0 9 13 13 7 15 9 9 0 13 16 9 14 1 1 9 1 9 13 7 3 15 1 9 9 7 9 9 1 15 1 9 0 0 13 7 9 15 14 16 3 1 9 9 13 2
35 9 13 2 9 16 1 9 0 9 13 7 9 13 9 13 16 0 9 14 16 1 9 0 9 15 9 4 13 2 9 9 9 0 13 2
68 9 9 1 1 9 9 9 9 1 9 0 7 9 1 9 9 13 2 9 9 9 9 9 1 12 12 9 1 12 12 9 2 9 0 7 0 9 2 9 9 1 0 9 9 2 9 9 9 1 9 9 7 9 7 9 9 15 1 9 0 1 3 1 9 9 9 13 2
14 15 9 13 2 3 9 2 9 0 3 3 9 13 2
31 10 9 16 9 0 1 9 7 7 9 0 1 9 1 1 12 9 7 7 9 2 9 9 1 9 0 7 0 15 13 2
21 9 13 2 9 13 1 9 0 9 9 0 9 0 0 1 9 7 9 9 13 2
16 1 9 12 9 0 16 12 9 0 9 7 9 9 13 13 2
33 15 9 13 1 9 10 9 16 9 0 1 9 7 9 9 0 2 0 7 0 1 9 13 2 9 9 0 15 14 0 4 13 2
48 9 9 7 9 0 16 9 9 1 9 0 0 7 0 7 0 9 14 0 9 7 9 13 2 1 9 9 9 0 1 9 0 1 9 9 9 13 16 3 15 14 1 3 9 9 4 13 2
14 9 13 2 15 9 13 16 1 9 1 15 3 13 2
14 9 13 7 13 7 13 2 6 8 9 15 16 13 2
10 9 9 9 3 9 9 14 9 13 2
4 3 6 9 2
13 9 15 14 16 9 13 2 16 3 9 4 13 2
40 8 8 16 1 9 1 9 9 13 2 7 1 9 7 9 7 9 7 9 15 9 13 2 1 9 13 2 15 9 1 9 13 7 9 14 16 3 9 13 2
9 9 9 2 9 9 9 13 13 2
7 9 0 7 0 13 13 2
6 9 9 9 13 13 2
19 9 1 9 0 2 7 9 0 2 9 7 9 9 9 9 9 15 13 2
19 3 2 10 3 9 9 13 9 9 7 9 7 9 0 14 1 9 13 2
13 9 1 9 9 7 9 1 10 9 9 13 13 2
10 13 9 1 9 0 9 9 0 13 2
38 3 16 9 0 9 0 13 2 9 9 13 2 7 9 1 9 9 1 9 13 16 9 10 12 9 15 13 3 9 9 9 8 9 9 7 9 9 2
25 9 10 3 0 7 9 7 0 13 16 3 9 16 9 9 9 9 13 16 13 1 9 9 13 2
20 9 1 9 13 2 6 9 2 3 9 1 9 16 1 15 13 1 15 13 2
14 9 3 4 13 16 7 15 14 1 9 9 9 13 2
18 7 13 16 15 14 9 13 16 12 9 7 12 9 1 9 15 13 2
9 3 4 9 14 1 9 0 13 2
18 9 1 9 9 13 13 16 15 9 13 16 3 1 15 9 9 13 2
17 1 9 9 16 15 14 1 9 15 9 7 9 15 9 1 13 2
28 15 9 9 0 7 9 0 13 2 16 9 0 9 7 9 15 14 1 9 0 16 9 0 13 2 9 13 2
20 1 9 7 10 9 3 16 9 9 13 9 13 2 9 1 9 15 9 13 2
33 9 16 9 15 3 9 9 2 9 9 13 1 9 9 9 9 13 2 7 1 9 9 9 9 1 9 7 9 9 9 0 13 2
18 7 3 16 1 9 9 0 13 9 15 14 9 1 9 1 9 13 2
32 3 10 9 9 2 9 0 1 9 9 9 0 13 2 16 3 0 13 0 9 7 9 9 0 16 1 9 7 9 4 13 2
8 9 3 1 9 15 9 13 2
7 9 9 9 9 9 13 2
15 15 1 9 15 7 9 15 3 9 14 1 9 13 13 2
11 9 9 13 9 14 1 9 9 9 13 2
5 9 0 13 13 2
4 9 0 13 2
35 9 9 13 16 1 9 16 9 3 0 13 7 9 9 9 1 10 9 0 1 10 9 7 9 0 9 13 1 9 1 9 9 9 13 2
9 9 13 2 9 14 9 9 13 2
20 9 1 0 15 7 1 9 9 1 9 13 1 9 13 7 1 9 9 13 2
18 13 2 13 16 1 9 9 7 9 9 16 1 9 10 9 13 13 2
8 15 16 16 1 9 9 13 2
24 15 0 13 16 3 1 9 15 2 3 3 1 0 9 9 2 3 9 9 7 9 0 13 2
14 3 1 15 15 9 0 13 16 9 1 15 9 13 2
12 9 15 9 14 1 9 9 15 15 9 13 2
12 9 13 1 10 9 9 15 1 9 9 13 2
15 9 7 9 9 9 1 9 9 3 1 9 9 9 13 2
22 16 9 1 9 1 9 0 1 9 13 13 2 8 8 9 16 1 9 10 9 13 2
33 9 1 9 8 9 9 13 2 16 15 1 9 13 7 9 14 9 13 7 9 9 13 2 15 13 7 1 15 9 9 9 13 2
21 16 9 13 2 9 14 9 13 7 9 13 1 9 9 9 7 9 7 9 9 2
34 9 9 9 0 3 1 9 1 9 9 9 9 9 1 9 9 9 9 9 13 7 9 9 0 9 9 9 1 9 9 10 9 13 2
56 1 10 9 13 13 13 2 9 15 1 15 13 16 1 9 9 10 9 7 9 10 9 0 1 9 7 9 7 3 9 16 1 3 10 9 13 2 0 13 7 1 9 7 9 0 7 9 9 0 9 9 1 3 9 13 2
47 3 1 9 16 1 9 9 9 9 13 2 9 0 1 9 9 9 0 1 9 1 9 1 9 1 9 3 9 1 9 13 2 7 9 9 2 9 9 1 9 0 14 1 9 0 13 2
25 3 9 1 9 0 13 7 1 9 9 9 1 9 9 16 9 15 16 0 9 0 13 2 13 2
17 9 0 3 1 9 1 9 9 9 16 9 0 1 15 9 13 2
44 15 9 16 1 9 9 9 1 9 9 9 0 7 0 13 13 13 2 1 9 9 9 0 1 13 7 9 0 9 9 0 1 9 9 7 9 9 1 9 1 9 9 13 2
44 9 13 2 3 9 9 14 16 1 9 7 9 9 9 9 0 1 15 15 9 13 1 9 13 7 9 0 0 3 9 0 2 9 0 2 9 9 7 2 14 3 0 13 2
10 9 1 9 0 9 9 9 9 13 2
39 1 9 9 0 9 7 9 9 0 7 9 9 12 1 9 9 9 9 9 9 1 9 10 9 1 9 9 1 9 0 1 9 9 9 1 9 1 13 2
35 1 9 9 0 9 9 0 9 2 1 10 9 12 9 1 9 9 9 9 1 9 0 9 2 9 7 9 9 1 9 9 9 9 13 2
38 10 9 9 9 9 0 9 9 2 9 2 9 2 9 7 9 3 9 9 2 9 9 9 2 9 9 9 2 9 9 9 7 9 9 9 9 13 2
17 0 9 10 9 9 9 9 13 16 1 9 9 9 9 13 13 2
22 9 9 9 9 7 9 0 9 9 9 9 1 10 9 1 9 0 1 10 9 13 2
10 9 9 9 1 9 1 9 1 13 2
17 9 9 9 1 0 9 9 9 1 9 9 1 1 9 9 13 2
27 10 9 1 9 9 9 9 13 1 9 12 9 1 9 9 9 9 9 7 9 9 9 9 9 13 13 2
19 9 9 9 9 9 14 9 0 9 13 16 9 15 3 0 7 0 13 2
22 9 10 9 0 0 13 16 15 1 9 15 1 9 9 0 1 9 0 9 9 13 2
18 9 9 9 1 9 9 9 16 3 1 9 9 1 9 13 13 13 2
41 9 9 9 9 1 9 9 1 9 9 1 9 0 9 9 15 1 9 2 9 9 15 14 9 9 13 7 13 2 10 9 9 14 0 13 7 9 14 0 13 2
17 10 9 1 9 9 9 13 2 0 9 10 9 1 9 15 13 2
45 9 3 1 9 9 1 0 9 9 9 9 13 7 1 1 9 0 16 9 0 9 1 9 9 13 2 13 2 10 9 1 10 9 16 9 9 1 9 9 9 9 13 2 13 2
30 1 9 10 9 2 9 9 0 9 9 13 16 9 13 1 9 9 9 7 9 1 9 7 9 9 7 9 1 9 2
9 9 9 9 9 1 9 9 13 2
31 9 9 9 9 9 9 1 9 9 9 9 9 9 7 9 0 7 9 9 9 9 9 9 9 2 1 10 9 9 13 2
34 1 10 9 9 1 9 9 2 9 9 2 9 9 2 9 9 2 9 9 2 9 9 2 9 9 7 9 9 1 9 13 13 13 2
53 9 0 1 10 9 16 1 9 9 9 0 9 2 9 9 7 9 0 7 9 0 9 2 9 7 9 9 1 9 13 13 2 9 1 9 7 9 0 15 14 1 9 9 9 1 9 9 9 7 9 9 13 2
41 9 9 8 9 9 9 9 9 1 9 9 7 9 9 0 2 1 9 9 0 13 2 10 9 1 9 9 9 7 9 9 0 1 9 0 1 9 0 0 13 2
15 15 1 9 7 9 9 9 9 9 0 9 7 9 13 2
33 9 9 16 9 9 0 14 9 9 9 13 7 13 2 9 0 9 9 2 9 7 9 9 0 14 1 9 1 9 15 9 13 2
28 15 9 13 2 9 9 0 1 10 9 9 0 13 16 9 9 9 1 0 9 10 9 1 9 0 0 13 2
38 1 9 9 9 9 9 9 2 9 0 1 9 2 9 7 9 9 0 2 9 9 0 9 2 9 7 9 9 7 9 9 9 1 10 9 9 13 2
9 9 0 0 9 9 14 9 13 2
19 9 9 9 9 0 2 0 1 9 2 9 0 9 9 9 14 9 13 2
50 1 9 9 0 9 9 9 9 2 10 9 0 9 0 9 9 14 1 9 12 9 9 1 9 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 7 9 1 9 15 13 2
18 16 1 10 9 9 9 9 9 7 9 9 9 1 9 9 9 13 2
20 12 7 0 9 9 9 7 9 9 1 12 1 12 9 1 9 1 9 13 2
34 1 10 9 1 9 1 1 9 2 0 1 9 2 2 9 0 2 9 2 9 9 2 0 9 9 9 1 9 9 10 9 9 13 2
39 9 2 0 1 9 2 3 1 15 9 0 9 9 0 9 9 9 14 1 9 15 13 7 1 9 9 9 9 0 9 1 9 9 9 1 9 1 13 2
30 12 9 9 9 9 0 9 13 2 10 9 1 9 0 12 12 12 9 1 9 15 14 1 9 9 9 9 13 13 2
48 9 9 1 9 9 9 9 9 0 9 9 1 9 13 2 10 9 1 9 9 0 7 0 1 9 9 2 9 7 9 2 9 2 9 2 9 0 9 2 9 0 7 9 0 9 13 13 2
20 15 16 13 2 9 9 0 3 12 9 0 9 0 9 0 9 14 9 13 2
34 15 13 2 1 9 9 12 12 9 1 9 9 2 12 12 12 9 1 9 9 0 7 9 1 9 0 2 0 7 0 9 13 13 2
23 9 13 2 9 3 9 0 1 9 9 9 12 9 7 1 9 9 12 9 9 13 13 2
24 10 9 1 9 0 10 9 2 0 9 1 9 9 13 16 9 3 9 16 1 15 4 13 2
18 1 10 9 2 9 9 9 0 0 7 0 1 12 9 0 15 13 2
27 1 9 9 16 1 9 9 13 7 1 15 9 13 2 9 0 9 0 13 16 3 1 9 0 9 13 2
56 9 16 1 10 9 9 1 9 1 9 13 1 15 9 15 1 10 9 13 3 13 2 9 0 1 9 9 16 3 1 12 9 9 9 13 13 7 1 9 0 15 1 9 9 9 9 9 13 13 7 1 15 7 9 13 2
25 1 15 1 15 1 9 15 13 9 0 16 1 9 4 9 15 14 1 9 9 9 13 9 13 2
43 9 0 16 9 9 9 15 1 0 9 9 7 9 9 13 13 7 9 15 16 0 13 1 9 0 1 15 9 13 7 1 10 9 13 16 1 9 9 9 9 9 13 2
12 10 9 3 1 9 0 1 9 9 13 13 2
19 1 9 9 9 9 0 9 1 9 1 12 9 0 15 0 9 0 13 2
10 9 0 3 1 9 0 16 0 13 2
38 3 1 9 2 7 3 3 1 9 7 1 9 15 2 1 9 9 0 1 9 16 1 9 9 13 13 2 9 14 9 0 2 0 7 3 0 13 2
90 7 9 16 1 9 0 9 1 9 1 9 0 9 13 9 13 16 1 3 9 15 1 9 0 9 0 9 13 2 9 16 1 9 7 9 9 13 2 1 9 1 12 1 9 15 13 7 3 1 9 15 1 9 7 9 2 7 1 1 15 9 0 13 2 1 9 15 9 13 2 7 9 15 9 0 0 3 9 9 7 9 7 9 14 1 15 9 13 13 2
36 9 10 9 15 13 16 1 9 9 0 7 9 9 0 9 16 1 9 15 9 13 2 9 9 9 9 3 0 7 9 1 15 3 0 13 2
18 0 9 16 1 9 1 9 9 7 9 9 13 1 9 15 9 13 2
10 1 9 9 2 9 10 9 0 13 2
32 0 1 12 9 3 1 9 15 1 9 13 16 1 9 9 9 9 9 13 7 15 1 15 1 9 12 9 14 1 1 13 2
56 0 13 16 15 10 9 13 1 9 13 2 7 9 16 1 12 12 9 1 9 1 9 9 0 1 9 13 1 9 15 13 13 16 1 10 9 15 14 16 13 1 9 13 2 1 15 9 9 15 1 9 0 13 0 13 2
16 10 9 3 0 13 2 16 9 9 1 10 9 0 13 13 2
28 0 9 16 1 9 9 1 9 13 2 9 0 13 2 7 10 9 1 9 9 16 1 9 0 9 13 13 2
14 9 16 1 10 9 9 13 1 9 0 9 13 13 2
46 9 1 9 9 2 1 0 1 9 9 2 16 13 9 13 16 9 9 1 9 0 0 7 9 1 9 0 1 1 9 9 13 2 1 9 15 1 10 9 9 1 9 9 15 13 2
22 1 10 9 2 9 0 2 0 1 9 9 2 9 13 16 10 9 14 9 0 13 2
45 9 9 10 12 9 14 16 9 1 9 9 9 15 13 13 7 0 9 7 9 1 9 9 13 1 9 9 13 7 10 9 14 16 1 9 7 9 9 9 9 13 1 15 13 2
22 1 10 9 2 1 10 9 9 16 16 1 9 10 9 9 7 9 13 2 0 13 2
64 1 10 9 2 9 16 1 9 15 1 9 7 9 0 13 7 9 9 0 13 7 1 9 15 3 9 0 0 13 16 9 3 9 1 9 12 9 0 1 15 0 13 2 1 9 9 1 9 9 0 7 0 0 13 16 10 9 1 9 9 1 9 13 2
33 1 9 0 10 9 0 16 1 9 9 7 9 1 9 13 13 15 13 16 3 3 1 9 0 3 9 9 14 1 9 9 13 2
42 3 9 16 1 9 9 0 2 0 7 0 9 9 9 2 9 0 2 13 13 13 2 7 9 3 0 9 1 9 0 9 13 13 2 0 1 10 9 0 3 13 2
31 9 9 3 9 13 13 16 12 9 0 1 9 16 9 13 13 7 9 10 9 14 16 1 9 9 0 9 15 0 13 2
45 1 3 9 9 1 9 9 1 13 7 15 1 9 15 14 2 16 1 3 3 9 0 15 7 9 1 9 0 9 9 0 7 9 9 9 9 13 2 1 9 15 9 13 13 2
18 1 9 7 15 1 9 9 9 1 3 9 3 9 1 9 9 13 2
41 3 13 16 9 9 9 2 1 9 9 0 7 9 9 0 1 9 12 9 0 1 13 7 9 7 9 2 1 1 9 0 9 2 1 9 7 9 10 9 13 2
26 4 13 16 9 9 0 1 3 9 14 13 7 9 15 14 1 9 9 16 1 15 9 13 9 13 2
23 3 1 10 9 9 9 9 9 13 2 16 9 0 15 9 1 9 9 0 0 15 13 2
26 3 9 9 1 0 0 9 0 13 7 9 9 0 9 2 16 1 9 3 0 7 3 0 15 0 2
6 10 9 12 9 13 2
16 7 9 10 9 9 7 9 7 9 10 9 14 1 15 13 2
50 16 9 10 9 9 0 9 1 9 0 0 13 3 1 10 9 13 16 15 1 9 9 15 7 1 9 9 7 9 15 2 9 0 7 9 1 9 7 9 7 9 0 7 0 0 1 10 9 13 2
62 3 1 9 9 9 0 9 2 0 9 16 13 15 13 16 9 7 9 0 0 16 9 13 7 13 0 13 2 9 9 14 13 7 1 9 7 9 9 0 15 9 13 7 1 9 7 9 10 9 7 9 1 15 13 2 9 0 1 9 15 13 2
23 9 16 9 13 7 9 16 13 2 7 9 7 9 9 9 7 9 0 1 15 0 13 2
10 9 9 3 9 7 9 14 13 13 2
11 10 9 1 9 0 2 9 9 9 13 2
11 9 0 7 0 1 9 9 9 9 13 2
24 9 9 9 0 14 16 15 7 9 9 9 9 13 7 9 0 1 9 9 0 9 13 13 2
29 12 9 0 7 0 10 9 2 9 9 9 9 9 0 0 9 9 13 7 9 14 1 9 0 15 1 9 13 2
17 9 1 9 9 9 9 13 7 1 9 1 9 9 0 13 13 2
56 12 4 9 15 9 2 9 0 9 9 2 7 9 0 9 15 13 16 1 9 0 7 0 15 10 9 0 14 0 13 7 1 9 13 7 9 0 1 9 7 1 15 9 9 7 9 0 7 0 1 9 0 1 9 13 2
22 3 9 7 9 9 7 9 0 16 9 0 13 1 9 9 15 1 10 9 0 13 2
17 10 0 7 9 15 1 9 9 2 1 9 9 1 9 13 13 2
23 10 9 1 9 9 8 0 13 7 9 9 9 9 9 15 14 1 9 9 1 9 13 2
41 0 13 16 0 9 3 1 10 9 2 9 9 16 9 9 9 9 9 9 7 9 9 1 15 14 1 9 13 1 9 9 9 2 1 9 9 7 9 9 13 2
29 12 9 1 9 10 9 2 1 9 1 10 9 16 3 1 15 2 1 9 12 9 9 9 13 13 16 13 13 2
30 9 9 9 9 9 13 2 3 1 9 12 9 9 9 1 9 12 12 9 2 9 1 9 9 9 9 9 9 13 2
29 9 9 9 13 2 9 9 2 9 7 9 10 9 1 9 0 9 1 9 9 9 9 9 9 2 0 13 13 2
37 15 13 2 3 1 9 9 12 0 9 0 9 2 9 0 2 9 7 9 1 9 12 12 9 9 9 0 13 16 10 15 1 10 9 9 13 2
39 9 0 13 2 1 9 9 9 9 9 2 10 9 1 10 9 9 4 13 7 12 0 9 10 9 0 12 12 9 9 9 0 0 9 1 9 4 13 2
60 9 9 9 9 2 9 9 9 0 1 9 14 1 9 9 12 12 7 12 9 9 13 7 13 2 3 9 9 2 9 2 9 7 9 9 9 9 1 9 9 9 13 16 1 10 9 10 9 9 0 9 9 1 9 9 9 9 4 13 2
19 9 12 12 7 12 9 1 9 1 9 0 9 9 1 10 9 9 13 2
22 9 9 9 9 9 0 9 9 13 2 9 1 9 9 2 9 7 9 9 0 13 2
18 15 13 2 9 9 1 9 9 2 3 0 1 9 0 9 13 13 2
23 15 13 2 9 9 9 9 9 16 1 9 9 9 0 9 3 1 9 0 9 0 13 2
29 1 10 9 9 9 9 7 9 0 7 0 9 9 16 12 9 0 7 0 10 9 14 1 9 9 0 13 13 2
20 9 9 16 1 9 9 1 10 9 13 1 9 9 1 9 0 0 4 13 2
22 9 9 9 13 2 9 9 9 1 9 12 12 9 1 9 0 9 10 9 9 13 2
23 9 9 13 2 10 9 9 9 1 9 1 9 9 9 2 1 1 9 12 9 9 13 2
40 15 13 2 9 13 16 3 0 1 12 12 9 9 9 9 9 7 9 1 9 9 13 16 1 9 1 9 2 1 1 9 0 12 1 12 9 9 4 13 2
52 9 7 9 1 9 7 9 7 7 9 0 0 13 16 9 15 9 9 7 7 9 9 13 7 7 1 9 1 9 9 7 9 1 9 1 9 7 9 9 7 9 1 9 9 1 9 9 7 9 9 13 2
18 9 4 13 16 1 3 9 7 9 9 7 9 1 15 9 0 13 2
24 9 0 2 9 9 7 9 1 9 9 9 7 9 2 9 3 0 1 9 9 1 9 13 2
12 16 9 10 12 9 7 9 9 9 0 13 2
43 10 9 1 9 0 9 13 7 1 9 7 9 2 9 9 7 9 7 9 14 9 13 7 1 9 9 7 9 7 9 0 7 0 2 9 9 0 0 7 0 15 13 2
31 1 3 9 16 3 9 9 7 9 0 13 13 2 9 1 9 9 7 9 9 9 7 9 7 9 9 1 9 15 13 2
20 9 1 9 9 0 7 9 9 0 1 9 7 9 7 1 9 0 9 13 2
39 9 9 9 1 3 9 9 13 16 9 0 9 7 9 9 1 9 15 13 7 7 1 9 0 9 9 1 15 1 9 2 15 14 9 13 2 9 13 2
16 9 7 9 12 9 13 16 9 1 9 9 1 9 14 13 2
37 7 9 16 1 9 0 9 7 9 13 2 9 1 9 16 0 7 0 1 9 13 2 9 9 13 16 9 1 15 0 7 0 9 14 13 13 2
41 15 16 1 9 9 0 9 1 9 9 9 0 2 9 9 13 7 3 10 9 1 15 1 9 9 9 9 13 2 12 9 0 13 16 1 9 10 9 0 13 2
63 4 9 0 1 9 7 9 0 1 9 9 9 1 9 9 0 1 9 9 9 7 9 9 9 2 9 13 7 1 9 7 9 9 1 9 0 1 9 9 9 7 9 9 13 7 1 9 9 0 1 9 0 9 0 2 9 9 1 9 14 9 13 2
28 9 0 9 9 1 0 9 1 0 9 9 9 9 9 16 1 9 9 9 13 2 1 12 9 9 9 13 2
32 9 9 1 9 0 7 9 9 1 9 0 2 12 9 9 15 1 0 9 9 13 16 1 9 0 9 7 9 9 9 13 2
27 9 1 0 9 15 1 1 9 1 9 12 1 12 0 13 7 3 9 1 9 14 1 10 9 0 13 2
54 15 1 0 9 15 1 1 9 1 9 0 9 13 7 1 9 7 9 0 14 1 9 12 1 12 1 9 15 1 9 13 13 2 1 9 10 9 1 9 12 1 12 9 13 7 1 9 9 3 1 9 0 13 2
18 1 10 9 9 9 0 1 9 9 13 7 9 9 1 9 0 13 2
41 9 9 9 0 9 15 16 1 9 0 10 9 1 0 9 15 1 9 12 1 12 1 9 1 9 9 13 7 3 9 0 15 14 1 9 12 1 12 9 13 2
26 15 1 0 9 15 1 9 9 9 0 13 7 1 9 12 1 12 1 10 9 1 9 9 0 13 2
17 9 9 10 9 1 9 0 13 7 9 9 0 1 9 0 13 2
16 1 0 9 2 9 9 1 9 0 1 12 9 9 9 13 2
23 9 9 10 9 9 1 10 9 1 9 0 10 9 1 9 1 9 1 9 9 9 13 2
43 9 9 16 1 9 9 0 7 0 15 14 1 9 0 10 9 13 13 2 1 9 0 1 9 1 9 9 0 15 1 9 12 1 12 0 13 7 1 9 9 9 13 2
36 9 1 9 1 9 0 0 13 13 2 9 9 9 2 9 7 9 14 1 9 1 9 12 1 12 2 12 1 12 7 12 1 12 9 13 2
22 1 10 9 9 0 1 9 9 9 13 7 9 9 7 9 3 1 9 9 9 13 2
34 1 9 0 2 9 9 9 0 0 3 1 9 1 9 1 9 7 9 1 9 0 1 9 9 0 0 13 7 1 9 1 9 13 2
21 9 9 1 9 0 10 9 16 9 12 1 9 9 9 0 13 1 9 0 13 2
15 9 9 1 10 9 12 9 9 7 12 9 9 13 13 2
29 9 9 2 9 9 12 7 0 0 9 9 9 0 9 9 7 12 9 0 9 9 9 1 10 9 14 9 13 2
40 1 9 0 9 9 9 9 1 9 9 12 9 7 9 12 9 2 12 9 0 15 14 1 9 7 9 1 1 9 9 9 9 7 9 9 9 0 4 13 2
43 9 0 0 1 9 9 9 9 15 13 16 9 0 9 9 13 10 9 12 1 12 9 9 9 16 9 9 7 9 9 1 9 9 1 9 9 9 9 0 9 4 13 2
45 1 9 0 2 9 9 9 9 9 1 9 9 9 0 9 0 7 9 15 1 9 9 13 2 15 9 0 1 9 7 9 9 9 0 13 7 1 9 9 9 1 9 9 13 2
46 9 7 9 9 1 9 9 0 9 0 13 16 0 9 9 9 9 9 9 13 7 9 9 1 9 9 9 9 0 4 13 7 1 9 9 1 9 9 9 0 9 0 9 13 13 2
35 15 1 9 13 16 9 9 9 9 0 9 9 9 13 16 9 9 9 13 7 9 9 16 1 9 9 1 9 0 15 9 0 13 13 2
31 1 9 10 9 9 9 9 9 9 0 1 9 9 9 13 16 9 0 3 1 9 9 1 9 0 9 9 9 9 13 2
23 9 9 9 0 9 16 1 9 9 1 9 9 0 9 0 9 1 9 9 0 9 13 2
26 9 9 9 9 0 16 1 9 9 9 15 2 9 13 16 1 9 9 9 1 9 9 0 9 13 2
37 1 10 9 2 9 9 2 12 9 9 9 9 0 1 9 15 16 9 15 1 9 0 9 13 13 16 9 9 3 1 9 9 9 9 13 13 2
15 1 9 9 0 9 9 16 1 9 9 7 9 9 13 2
26 9 9 10 9 1 9 9 9 1 9 1 9 9 12 9 9 7 12 9 9 9 1 9 9 13 2
20 9 9 9 7 9 16 1 9 9 9 3 1 9 9 1 9 0 13 13 2
18 9 9 13 13 15 1 9 16 13 1 9 9 9 0 1 9 13 2
56 9 9 1 10 9 9 0 13 16 15 16 1 1 13 2 3 1 9 16 10 9 1 9 9 7 9 0 0 1 9 0 1 9 13 2 9 9 1 15 13 16 9 9 9 12 0 9 1 12 9 0 15 0 4 13 2
16 0 9 15 16 9 9 1 9 9 7 9 1 9 15 13 2
75 1 9 9 0 2 1 9 0 2 9 1 9 9 9 2 9 9 7 0 9 9 0 9 9 16 9 14 1 9 0 1 9 13 1 1 9 12 9 9 7 12 9 9 1 9 9 9 9 9 9 13 7 9 16 1 15 9 13 13 2 7 1 10 9 2 10 12 9 9 0 14 9 13 13 2
46 1 9 0 2 9 2 9 9 9 9 7 9 9 2 9 9 9 9 14 1 9 9 9 9 9 9 9 0 9 13 1 9 7 10 12 1 9 9 9 1 9 9 9 9 13 2
20 3 9 9 1 1 9 9 0 1 12 9 0 9 0 9 16 1 9 13 2
37 9 9 9 1 9 9 9 16 12 3 0 13 2 1 9 1 9 9 9 13 2 1 9 7 9 9 7 9 9 9 9 9 9 9 9 13 2
64 1 10 9 2 9 9 9 12 9 0 9 0 9 7 9 9 9 9 7 9 9 16 9 9 0 14 1 9 13 7 1 9 0 1 9 9 13 16 1 0 9 0 1 9 9 15 2 9 0 0 13 7 1 9 10 9 1 3 9 0 9 13 13 2
35 10 12 9 2 1 9 9 9 1 9 0 9 13 7 3 0 13 16 16 9 15 1 1 9 9 0 10 9 9 9 4 13 7 3 2
25 1 10 9 13 13 2 9 9 9 9 9 1 9 1 9 9 0 9 1 9 9 9 9 13 2
25 9 9 9 12 9 13 16 1 9 0 9 2 12 9 1 9 15 2 12 9 7 12 9 13 2
18 9 9 1 12 9 0 13 13 2 9 9 1 9 1 9 9 13 2
46 1 10 9 13 13 13 2 0 9 3 1 9 9 1 1 9 7 9 9 1 15 1 9 9 9 16 1 9 9 1 9 0 13 2 15 3 1 9 9 3 10 9 14 9 13 2
46 15 1 9 3 1 9 9 13 2 9 9 9 7 9 0 0 0 13 2 10 9 1 9 0 7 9 0 1 9 9 7 1 1 15 9 9 9 2 1 9 1 9 9 0 13 2
35 9 1 9 9 10 9 9 13 2 1 9 3 1 9 2 12 1 9 0 2 9 1 15 9 13 7 13 2 13 1 15 3 13 13 2
9 13 2 9 7 0 7 9 13 2
16 9 15 15 13 16 9 16 9 1 10 9 9 13 14 13 2
8 15 13 2 13 2 9 13 2
4 9 9 13 2
22 9 13 2 9 13 2 13 16 9 13 13 2 9 9 13 2 3 9 9 13 13 2
7 16 16 13 2 3 9 2
48 9 9 1 9 1 15 16 9 9 2 9 7 9 9 14 9 13 7 15 14 1 9 7 0 7 9 0 13 2 9 13 2 1 9 1 3 9 0 1 1 9 9 0 2 9 0 13 2
53 9 16 9 0 14 0 10 9 9 0 0 7 1 9 9 0 13 7 9 13 2 16 16 9 12 9 1 9 16 1 10 9 2 1 9 7 9 13 1 9 9 0 7 9 0 9 1 15 1 9 9 13 2
19 15 13 2 3 2 9 7 9 0 15 1 9 9 9 9 3 9 13 2
20 15 13 9 9 14 1 9 7 1 9 9 16 1 9 15 9 13 2 13 2
20 15 13 9 7 9 9 14 1 9 9 0 2 1 9 7 9 7 9 13 2
22 15 13 9 7 9 9 13 2 16 1 9 9 9 9 13 7 1 9 12 0 13 2
3 9 13 2
16 9 9 9 13 13 16 9 1 9 0 1 9 0 9 13 2
35 10 9 13 13 2 1 9 9 0 9 2 9 9 16 1 9 9 9 13 1 9 10 9 13 2 1 9 0 9 1 9 0 9 13 2
39 1 9 9 9 0 1 9 16 1 9 9 15 1 9 9 13 9 1 9 9 0 14 16 9 13 13 7 10 9 9 9 9 9 0 1 9 0 13 2
27 9 9 1 9 1 9 1 9 9 0 13 2 16 9 9 1 9 13 1 15 4 9 9 9 14 13 2
34 15 9 1 9 14 9 9 0 9 13 7 9 13 2 9 0 4 1 9 9 0 2 9 9 13 13 7 1 9 9 0 9 13 2
64 15 1 9 15 16 1 9 9 9 0 9 2 9 7 9 9 0 14 0 13 2 9 13 2 9 9 9 1 9 1 9 0 9 2 0 13 9 1 9 13 1 9 0 0 2 9 15 14 1 9 16 9 9 0 7 9 0 14 0 13 2 9 13 2
38 12 9 0 1 9 9 9 9 13 16 15 1 15 9 13 2 12 9 9 9 9 1 9 3 12 9 1 9 0 7 1 9 12 9 9 9 13 2
25 1 9 9 9 9 9 10 9 9 1 12 9 7 1 9 0 1 9 12 9 0 0 13 13 2
44 12 9 0 1 9 9 9 16 13 9 15 0 13 2 13 2 0 9 9 9 0 9 9 1 9 12 0 1 12 9 0 13 16 9 1 9 9 12 9 1 9 0 13 2
37 15 13 2 1 9 9 1 9 0 1 3 16 12 9 1 9 9 9 9 9 13 2 3 12 9 9 9 9 9 0 1 12 9 9 9 13 2
22 1 9 9 9 9 9 9 2 9 1 9 2 1 10 9 9 1 9 0 9 13 2
19 10 9 9 9 7 9 9 0 9 7 9 9 9 1 9 9 13 13 2
17 9 9 15 0 13 9 9 1 9 9 3 3 12 9 9 13 2
12 16 9 9 9 7 9 9 12 9 9 13 2
39 1 10 9 9 10 9 9 12 9 1 1 12 9 0 12 9 2 9 0 9 9 12 12 9 2 9 9 12 12 9 7 9 9 12 12 9 9 13 2
30 9 9 9 7 9 0 13 9 9 1 9 9 9 9 9 9 0 9 7 9 1 9 7 9 9 10 9 13 13 2
31 12 9 1 9 13 1 9 9 0 3 0 9 1 9 9 9 13 16 15 9 9 9 13 7 3 9 7 9 9 13 2
27 9 1 9 13 2 15 3 13 2 15 9 9 13 7 3 10 9 13 15 13 16 9 9 12 9 13 2
25 12 9 0 0 16 9 9 7 9 9 7 9 2 7 9 1 15 0 13 7 0 9 9 13 2
27 7 12 9 0 16 13 16 1 9 13 2 7 3 9 0 1 15 9 13 7 1 1 15 3 0 13 2
11 15 3 1 9 0 0 13 2 7 15 2
4 3 9 13 2
9 9 9 1 9 0 9 9 13 2
15 9 13 9 2 9 7 9 14 3 13 9 0 13 13 2
102 0 7 0 13 7 0 1 15 0 7 0 7 0 13 7 10 9 14 15 9 3 1 15 7 15 14 3 13 1 9 1 9 9 13 3 0 7 0 13 7 16 9 9 13 7 9 9 13 1 9 9 0 9 4 13 16 1 9 7 9 15 13 7 15 3 9 9 14 13 7 1 9 9 7 9 9 7 9 9 9 13 16 9 0 13 7 9 0 2 7 1 10 9 10 9 2 9 0 15 14 13 2
31 16 9 9 12 7 12 9 3 1 9 9 1 9 9 1 9 13 2 1 1 9 1 9 9 1 12 9 0 9 13 2
32 9 9 9 0 9 9 1 9 9 13 7 9 13 1 9 7 9 9 7 1 9 3 16 3 9 7 9 15 13 9 13 2
44 9 9 13 2 1 15 7 9 9 9 0 13 7 9 12 9 2 9 9 14 13 16 1 9 9 2 1 9 13 1 9 0 16 0 15 13 7 1 9 9 0 14 13 2
31 7 9 15 2 16 0 7 0 13 2 9 1 9 9 0 13 2 9 1 9 0 9 13 16 1 9 9 9 13 13 2
45 9 1 9 15 9 13 2 16 9 13 9 9 9 9 16 1 9 13 13 1 9 1 15 9 9 0 15 9 15 14 0 13 7 10 9 9 13 16 9 1 9 0 15 13 2
9 9 3 12 9 0 1 9 13 2
12 15 1 1 9 13 7 9 9 9 15 13 2
27 9 9 1 9 10 9 13 2 3 1 15 7 9 9 15 14 9 13 2 9 1 9 7 9 0 13 2
20 9 1 15 0 13 15 14 13 2 7 9 0 15 14 1 9 9 15 13 2
16 10 9 2 9 15 14 1 9 13 2 7 1 9 9 13 2
17 3 9 1 9 9 13 2 7 9 0 2 9 9 14 9 13 2
15 3 1 15 7 9 1 9 9 13 12 9 9 0 13 2
8 9 9 9 9 9 9 13 2
8 9 9 13 9 15 15 13 2
5 15 3 9 13 2
16 3 9 1 9 10 9 9 13 16 13 2 13 2 9 13 2
10 13 2 16 9 13 1 9 15 13 2
21 1 10 9 9 9 2 9 0 13 2 7 1 10 9 13 9 9 14 0 13 2
26 9 9 13 16 9 9 7 3 9 4 1 9 9 9 13 7 0 13 16 9 1 9 9 9 13 2
16 7 15 16 0 13 16 9 9 0 13 7 9 9 0 13 2
8 7 9 13 2 7 9 13 2
35 16 9 1 9 9 7 9 0 1 9 9 14 9 13 7 1 9 7 9 9 9 1 13 7 0 13 1 9 10 9 0 3 9 13 2
26 10 9 14 15 1 9 13 2 9 15 0 13 7 0 1 9 9 2 7 9 9 9 16 13 13 2
23 9 9 16 1 9 0 9 9 13 1 9 13 7 12 9 0 9 13 7 9 15 13 2
4 15 9 13 2
38 1 9 15 9 13 7 13 2 9 9 9 2 9 9 13 2 15 16 13 9 13 4 9 14 13 2 7 16 13 0 13 3 1 9 4 9 13 2
45 9 15 16 1 9 0 9 13 7 3 9 15 13 9 13 2 9 1 9 13 2 9 14 13 2 16 2 1 9 0 0 1 9 0 13 1 10 9 9 13 2 7 3 13 2
8 0 9 0 1 10 9 13 2
42 12 9 0 16 3 0 16 13 2 16 9 15 14 1 9 13 2 3 1 9 9 2 7 9 0 2 9 1 9 15 13 2 9 9 9 2 15 16 9 14 13 2
19 7 9 15 3 1 9 15 13 2 9 14 13 7 9 1 9 9 13 2
15 9 0 16 16 15 14 1 15 9 13 2 12 9 13 2
17 9 13 7 15 14 1 9 13 16 10 9 14 9 1 9 13 2
27 7 1 10 9 16 9 9 13 16 15 9 13 16 1 9 12 9 0 1 9 13 13 16 10 9 13 2
8 7 13 2 8 8 8 8 2
41 9 1 0 9 16 9 1 9 9 13 2 1 0 9 15 13 13 2 1 9 9 9 2 3 9 0 9 13 3 9 9 1 1 9 0 7 9 0 0 13 2
28 12 9 0 13 0 9 9 13 16 9 13 13 3 9 15 2 1 9 15 2 3 9 13 16 1 9 13 2
26 0 13 9 2 9 0 9 9 9 2 9 9 14 2 1 9 1 9 0 15 13 1 10 9 0 2
7 3 7 0 13 9 13 2
42 9 13 9 13 16 16 9 13 7 9 13 2 9 0 15 16 13 2 7 10 9 0 1 9 9 16 9 13 1 10 9 9 9 0 13 2 3 10 9 9 9 2
31 1 3 1 10 9 9 7 9 1 15 0 13 13 2 9 9 0 15 1 10 9 13 2 9 9 0 1 10 9 13 2
3 15 13 2
15 10 9 16 9 9 15 14 0 13 2 9 15 3 13 2
6 9 9 2 9 12 2
9 0 9 1 9 15 15 16 13 2
21 8 16 12 9 7 9 1 9 13 3 9 9 9 12 9 0 1 9 13 13 7
63 12 12 9 13 1 10 9 15 15 9 0 14 1 9 9 9 9 0 7 12 9 0 15 15 9 13 7 9 13 2 12 9 1 9 15 1 9 13 16 13 2 7 9 0 2 9 7 9 1 9 9 7 9 9 13 7 9 9 9 9 9 13 2
63 9 9 16 9 9 9 9 13 16 3 1 9 9 9 9 13 16 9 9 15 14 1 9 9 2 9 13 7 15 1 9 9 9 9 13 16 9 9 12 9 9 7 12 9 9 13 12 9 3 15 16 9 7 9 15 0 13 9 0 0 13 13 2
36 9 9 9 9 9 9 14 13 16 15 14 3 1 9 13 7 3 13 7 9 1 9 13 1 1 9 7 9 9 13 7 9 14 0 13 2
54 15 13 0 13 9 9 13 2 7 0 9 9 15 13 7 9 1 9 9 13 7 9 1 15 16 9 9 9 13 13 16 1 12 12 9 9 13 2 7 9 16 10 12 12 9 14 1 9 13 9 9 9 13 2
21 3 9 1 15 0 16 9 9 2 12 9 13 1 1 9 9 9 9 9 13 2
22 15 14 16 13 2 16 10 9 2 0 9 1 9 9 13 16 9 15 1 9 13 2
35 15 9 13 16 12 7 3 12 9 0 9 9 7 9 1 9 9 13 13 13 16 9 9 0 13 2 7 9 15 1 10 9 9 13 2
35 3 9 9 13 16 15 9 9 13 16 1 9 7 16 1 9 9 2 16 1 8 8 7 16 1 9 2 16 1 9 7 16 1 9 2
5 9 1 15 0 2
76 15 0 13 16 10 9 12 12 9 9 9 9 13 13 7 12 9 15 14 9 13 2 10 9 9 9 9 9 2 10 9 14 2 3 1 12 12 9 2 7 1 12 12 9 9 13 7 1 9 9 0 15 13 7 3 1 10 9 2 9 3 0 13 16 13 2 10 3 13 13 2 10 3 13 13 2
25 9 13 10 9 0 9 15 16 1 9 9 9 7 9 3 0 13 16 9 15 14 9 9 13 2
11 10 9 3 9 15 3 0 7 0 13 2
24 1 9 9 7 9 0 9 9 2 9 0 9 9 2 3 1 9 0 0 9 0 4 13 2
21 10 9 1 9 9 1 9 0 9 1 9 9 0 7 9 0 0 1 9 13 2
12 9 16 0 9 9 1 15 1 9 4 13 2
30 1 9 9 9 0 4 9 9 0 3 2 7 9 7 9 9 0 1 9 7 9 1 9 0 14 1 9 9 13 2
20 1 10 9 9 9 3 9 9 1 9 9 7 15 14 9 13 0 4 13 2
17 9 9 9 0 13 9 0 9 1 9 9 9 9 12 9 13 2
7 9 16 9 14 9 13 2
17 9 0 9 13 16 9 2 9 2 9 7 9 9 14 9 13 2
23 9 9 9 9 1 12 9 2 10 9 14 16 9 9 13 1 9 7 9 9 13 13 2
19 9 9 9 13 2 9 16 9 13 9 9 14 9 13 2 1 9 13 2
22 9 9 9 1 9 9 16 13 2 9 1 9 1 9 9 3 9 7 9 9 13 2
30 9 13 2 3 1 15 13 9 0 3 9 9 14 9 13 7 9 3 9 13 2 7 9 0 15 14 9 13 13 2
19 9 16 9 1 9 9 7 9 9 13 2 0 1 9 9 14 9 13 2
21 10 9 3 1 1 9 9 7 9 7 7 10 12 1 0 9 9 0 9 13 2
18 9 0 1 9 9 9 0 9 1 9 9 0 7 7 9 9 13 2
27 9 0 13 16 9 9 1 9 9 15 1 9 9 0 2 9 1 9 0 1 9 9 9 14 9 13 2
47 9 9 2 9 9 9 13 2 9 9 9 0 14 9 13 7 16 9 9 9 9 7 9 9 14 1 9 13 10 9 9 1 9 13 7 9 1 0 7 0 9 9 9 15 9 13 2
44 9 9 9 9 9 1 9 0 16 9 9 9 7 9 9 14 1 9 13 13 2 0 13 16 10 9 3 1 9 9 1 9 15 1 12 7 12 9 9 0 14 9 13 2
22 9 1 9 13 16 1 9 9 1 9 9 9 0 7 9 15 1 9 9 0 13 2
27 1 9 0 9 9 9 0 9 2 9 9 9 9 1 1 9 9 1 9 12 9 9 1 9 0 13 2
64 1 9 9 9 2 1 10 9 16 1 9 2 1 1 9 9 7 9 9 9 9 13 2 12 9 1 9 16 9 9 9 1 9 7 9 13 2 1 9 9 0 2 9 15 14 1 9 0 9 9 7 9 1 9 9 9 7 0 9 9 15 9 13 2
28 1 9 9 16 9 9 9 1 9 1 9 9 9 1 9 0 0 2 16 9 9 0 13 13 2 9 13 2
22 1 10 9 16 1 9 9 9 1 9 9 9 9 13 2 9 12 12 9 9 13 2
30 9 0 1 9 9 0 0 1 9 1 9 9 9 9 0 0 1 9 2 9 2 9 7 9 1 9 0 9 13 2
31 9 9 1 9 9 7 9 15 2 1 9 9 9 9 9 1 9 2 1 9 9 10 9 1 9 1 9 7 9 13 2
28 9 9 0 1 15 13 16 1 9 9 9 9 2 9 3 1 9 9 9 9 13 7 16 1 15 0 13 2
37 1 9 1 9 9 0 2 1 9 9 9 9 1 9 2 4 9 0 14 9 13 7 1 9 15 1 9 9 0 1 9 9 0 16 9 13 2
22 1 9 2 9 9 9 13 16 9 9 9 9 1 9 9 7 9 16 9 0 13 2
17 1 9 9 0 9 2 12 9 0 9 9 9 1 9 9 13 2
19 9 10 9 9 13 9 1 9 0 7 9 0 0 14 1 9 9 13 2
23 1 9 1 10 9 2 9 9 1 9 0 1 9 13 13 13 16 1 15 1 9 13 2
18 1 10 9 1 9 0 0 1 9 7 9 0 0 9 9 13 13 2
35 10 9 0 0 9 13 16 1 0 9 9 13 0 1 9 0 14 3 9 9 1 9 0 9 13 7 1 9 15 1 9 0 0 13 2
11 0 1 12 9 9 1 9 9 9 13 2
32 0 1 12 9 1 9 12 9 9 1 9 9 9 13 7 12 9 1 9 10 12 9 2 1 9 9 0 9 9 9 13 2
59 9 9 9 9 9 0 9 1 9 0 9 9 0 1 9 0 1 9 12 7 0 16 9 9 0 1 9 15 1 9 9 9 9 13 2 13 2 1 1 9 1 9 9 7 0 1 12 9 1 9 9 9 3 1 9 9 13 13 2
25 9 0 9 13 9 9 16 9 9 15 14 13 2 13 0 9 9 9 1 9 1 9 9 13 2
21 1 9 9 1 9 2 10 9 0 1 9 13 7 1 9 9 0 9 9 13 2
24 9 9 13 2 9 9 0 1 12 9 0 1 9 9 9 15 3 1 9 1 10 9 13 2
28 15 16 13 2 16 9 9 10 9 0 13 2 7 3 3 0 13 16 15 14 1 9 9 9 9 9 13 2
30 10 9 13 2 9 1 9 9 0 3 13 1 10 9 9 13 7 9 1 9 9 0 3 4 1 9 9 9 13 2
47 9 9 1 9 0 1 9 9 9 9 1 9 1 15 16 9 9 0 9 9 9 9 1 0 9 1 9 1 9 9 9 13 2 13 2 10 9 2 9 7 9 0 1 0 9 13 2
27 1 0 10 9 2 9 1 9 9 0 9 3 9 9 2 1 10 9 1 9 2 9 1 9 13 13 2
25 9 0 9 10 9 2 9 9 9 9 13 16 1 9 9 1 9 9 1 9 9 2 9 13 2
21 10 9 13 2 9 0 2 1 9 9 0 0 2 3 1 0 9 9 0 13 2
21 9 0 16 3 1 9 9 9 0 13 3 1 12 9 9 1 9 9 9 13 2
18 7 9 9 2 10 9 14 1 9 0 13 7 9 1 9 0 13 2
35 1 9 9 2 1 1 9 3 9 13 13 16 9 9 9 1 9 1 1 9 0 2 1 12 9 9 0 2 12 9 0 0 9 13 2
55 1 9 10 9 2 9 0 15 2 9 0 0 0 7 0 13 16 1 9 9 9 9 9 1 9 12 2 9 1 13 7 9 1 9 0 2 1 9 9 0 1 9 2 9 0 2 7 9 9 7 9 2 9 13 2
34 9 0 9 13 2 9 14 16 0 9 1 9 12 9 13 13 7 1 3 1 15 1 9 9 0 9 13 13 2 9 0 9 13 2
86 1 9 9 9 1 9 2 9 9 9 9 1 9 9 9 9 13 2 9 0 1 9 12 1 9 12 12 9 9 2 10 12 2 12 9 12 9 1 1 15 13 16 10 12 9 12 9 1 0 9 1 9 13 16 0 9 15 1 9 12 13 7 1 9 12 7 12 9 0 1 0 9 1 9 13 7 9 0 1 9 9 1 9 3 13 2
24 10 9 13 16 9 12 16 1 9 12 2 12 12 9 9 13 2 3 9 1 9 9 13 2
13 9 13 2 9 10 9 1 12 1 12 9 13 2
19 9 0 12 9 0 0 1 9 14 1 9 9 1 9 9 0 9 13 2
10 9 0 1 9 9 9 9 9 13 2
33 9 9 1 9 9 16 1 9 9 1 9 3 9 13 0 2 1 9 0 13 7 1 9 1 9 9 0 9 13 7 9 13 2
25 9 0 1 0 9 1 9 9 12 0 9 13 7 1 10 9 9 1 10 9 9 0 9 13 2
20 9 1 3 0 9 9 1 9 13 16 13 1 9 9 0 9 7 9 13 2
34 9 0 9 0 13 16 1 10 9 9 0 13 7 9 9 0 13 1 9 15 1 9 0 9 9 13 16 9 0 14 1 9 13 2
24 10 9 0 0 1 9 12 9 9 0 13 7 0 12 2 12 9 9 7 12 9 9 13 2
24 9 9 9 0 9 16 1 9 0 1 9 9 0 1 9 9 1 13 13 2 9 9 13 2
39 1 9 9 1 9 9 12 0 16 1 9 12 9 1 9 12 7 0 9 9 9 9 14 1 9 13 2 3 1 9 9 9 9 0 14 1 9 13 2
17 9 1 9 12 1 9 0 9 1 12 9 9 0 9 9 13 2
31 9 15 16 9 9 13 1 9 9 9 9 13 7 9 0 9 9 16 1 9 12 13 16 1 0 9 0 9 9 13 2
28 9 1 9 1 9 15 16 1 0 9 9 0 9 14 1 9 0 9 16 9 9 13 1 9 9 9 13 2
18 9 9 1 9 12 3 1 9 9 15 9 1 9 9 9 9 13 2
23 9 16 1 9 12 9 3 9 9 13 1 9 12 1 12 9 9 9 14 1 9 13 2
24 1 9 9 16 9 15 1 9 9 1 9 13 2 9 16 0 13 1 9 9 9 0 13 2
59 1 9 9 9 1 9 9 9 13 10 9 3 1 9 9 13 2 7 9 0 9 9 9 2 10 9 14 1 12 9 16 1 9 9 0 13 13 2 9 13 7 13 16 12 2 12 1 12 9 9 10 9 0 1 9 9 9 13 2
26 9 9 9 0 10 9 9 1 9 9 0 13 13 16 9 9 1 10 9 13 9 0 1 9 13 2
29 15 13 2 9 9 0 1 10 12 9 3 3 1 9 9 13 16 12 7 12 9 3 1 1 9 0 13 13 2
31 9 9 0 9 9 7 9 9 0 0 9 13 13 13 2 7 1 3 9 9 9 9 14 3 1 1 9 9 13 13 2
8 6 9 2 15 3 0 13 2
7 9 0 7 9 0 13 2
18 1 9 0 9 13 7 9 0 14 13 16 1 10 9 1 15 13 2
20 1 9 7 9 1 9 9 0 9 13 7 3 13 16 1 1 9 1 13 2
11 1 10 10 9 9 9 7 9 1 13 2
10 3 15 15 14 1 9 9 9 13 2
24 3 9 16 1 13 7 1 10 9 13 2 7 9 15 9 0 9 9 9 14 1 9 13 2
18 10 9 0 1 9 16 1 9 9 7 9 9 13 9 3 0 13 2
23 9 13 16 15 14 1 9 15 13 2 16 9 10 9 0 9 14 1 9 0 15 13 2
26 6 9 0 9 2 16 10 9 0 14 16 9 0 7 0 13 7 9 9 15 13 2 0 4 13 2
7 6 9 2 15 3 13 2
16 9 0 15 3 9 9 13 7 15 14 1 9 9 0 13 2
26 9 15 1 15 1 9 7 9 9 13 7 10 9 15 14 1 13 16 13 2 9 15 3 0 13 2
36 3 1 0 9 9 9 0 15 14 16 3 9 0 9 13 13 2 7 9 0 15 14 2 6 9 15 1 0 9 13 16 1 15 9 13 2
12 7 15 7 9 15 14 3 1 9 4 13 2
28 1 0 9 7 9 4 13 2 7 1 15 9 3 9 1 9 0 7 0 2 0 9 15 9 15 4 13 2
13 9 15 2 10 9 9 13 2 1 15 9 13 2
16 16 15 16 15 9 9 15 15 14 1 9 15 1 4 13 2
34 1 1 9 0 1 9 9 1 9 9 9 2 9 9 9 10 9 1 1 9 9 0 0 7 9 0 1 9 9 9 9 9 13 2
59 1 9 9 0 9 2 1 1 9 0 1 9 9 9 9 9 0 1 9 7 9 0 12 1 9 9 16 9 9 9 0 7 9 9 0 1 10 9 13 2 9 0 1 1 9 9 0 7 9 9 0 1 9 9 10 9 13 13 2
81 1 1 10 9 2 10 9 3 0 13 16 9 0 7 0 9 1 0 9 1 12 9 0 1 12 9 1 9 9 7 9 0 9 13 16 1 9 9 7 9 1 10 9 3 0 16 1 0 7 0 9 0 1 9 13 2 9 13 7 1 9 10 9 7 9 9 13 16 3 9 1 9 9 0 7 0 15 14 9 13 2
45 10 9 0 13 2 9 0 16 1 9 9 0 7 0 1 9 9 9 13 2 3 9 9 14 9 13 2 7 10 9 16 1 9 9 0 0 13 2 13 13 1 9 9 13 2
34 9 9 0 9 9 16 3 9 9 13 7 9 3 1 9 9 9 7 3 1 9 9 13 13 9 9 9 12 9 9 15 14 13 2
82 1 9 9 13 7 13 9 9 0 13 16 9 15 0 13 2 7 16 9 13 7 13 9 9 13 2 9 15 14 9 15 14 1 9 0 13 7 1 9 9 15 13 2 15 3 9 1 9 9 9 13 7 15 1 10 9 16 9 15 14 1 9 0 13 2 9 13 7 9 9 13 16 1 10 9 1 12 9 0 9 13 2
32 9 9 15 3 9 14 1 0 9 13 7 9 9 1 9 9 0 9 9 7 9 9 15 14 9 0 0 1 9 0 13 2
22 3 9 13 16 9 1 9 12 0 15 0 13 7 13 2 9 15 14 9 12 13 2
25 9 9 3 0 9 13 7 9 9 14 16 9 15 0 13 7 9 15 14 0 13 13 2 13 2
17 10 9 13 2 15 1 15 9 13 16 9 15 14 9 12 13 2
7 15 3 9 15 14 13 2
43 10 9 1 9 15 9 13 7 13 2 9 9 15 9 12 14 9 13 7 9 0 9 14 9 13 7 15 3 9 15 3 9 9 9 13 7 3 9 15 3 9 13 2
27 10 9 16 9 9 13 13 3 0 13 7 1 9 9 13 2 9 15 14 16 12 0 1 15 0 13 2
39 9 9 9 15 14 16 13 7 10 9 9 15 14 16 9 15 14 1 10 9 9 1 10 9 9 13 13 13 2 0 7 9 14 1 10 9 9 13 2
36 10 9 13 7 1 0 15 16 15 16 13 1 9 13 2 13 2 1 10 9 9 9 9 13 7 1 9 9 15 3 9 1 1 15 13 2
14 0 15 2 1 15 9 13 7 1 9 9 9 13 2
12 15 16 9 15 14 13 7 10 9 1 8 2
24 1 9 15 16 1 1 15 13 16 9 15 14 0 13 2 15 3 9 9 15 14 13 13 2
39 1 15 7 12 9 12 1 9 1 9 15 0 13 7 3 9 0 15 14 1 9 15 9 13 7 9 13 2 15 1 3 9 2 9 9 15 3 13 2
28 7 15 10 12 9 9 2 1 9 15 0 13 7 3 15 1 9 9 15 0 13 16 9 0 7 0 14 2
54 9 9 0 13 2 15 1 9 9 15 3 0 13 7 1 9 9 16 1 9 13 2 9 14 7 12 9 9 14 1 9 9 9 9 13 7 9 14 9 13 7 9 9 14 9 9 13 7 9 13 7 9 13 2
77 7 3 16 1 9 9 9 1 13 2 1 9 0 0 9 13 7 9 12 9 9 16 1 10 9 13 2 9 9 14 3 13 7 16 10 9 9 9 0 10 9 13 7 15 3 13 15 14 1 15 0 13 7 16 15 14 1 10 9 0 13 2 3 16 3 9 0 1 15 0 13 7 15 14 3 13 2
5 9 9 0 13 2
36 9 9 9 9 9 9 9 9 13 2 9 0 9 9 1 9 9 0 1 9 12 1 9 12 9 1 9 3 12 9 14 1 9 4 13 2
21 1 9 9 9 2 9 13 2 9 15 9 9 0 1 12 9 1 9 14 13 2
31 9 4 1 9 9 9 13 16 16 12 9 14 1 9 9 9 13 7 15 7 12 9 0 14 1 9 9 0 0 13 2
18 9 9 9 1 9 9 12 9 0 1 9 0 9 9 0 9 13 2
15 1 9 9 2 1 9 10 9 12 12 9 9 4 13 2
27 9 13 2 1 12 9 10 9 12 0 4 9 7 9 14 1 9 9 3 1 1 9 0 9 0 13 2
20 9 9 1 9 12 9 2 12 1 9 9 9 1 10 9 9 1 9 13 2
8 9 9 9 0 9 9 13 2
27 9 0 9 9 9 2 9 9 1 9 1 9 0 1 9 2 9 9 9 9 9 0 9 14 9 13 2
22 1 9 9 2 16 9 9 9 9 2 15 1 9 9 2 1 9 1 9 0 13 2
36 9 0 9 9 9 2 3 1 9 9 9 9 0 10 9 1 9 9 1 9 9 0 7 9 1 9 2 15 14 1 9 1 9 9 13 2
29 9 1 9 1 9 0 9 13 2 9 9 0 1 12 9 14 16 1 9 9 7 9 15 9 13 2 9 13 2
27 1 1 10 9 2 9 13 16 9 9 9 10 9 0 7 0 9 0 10 9 7 9 15 14 9 13 2
31 1 0 9 0 9 9 0 9 13 13 16 9 0 9 0 0 1 9 9 3 9 0 0 2 9 7 15 1 9 13 2
44 15 1 9 13 16 9 0 0 13 13 16 9 9 9 9 9 0 14 9 13 2 9 9 0 14 9 13 2 9 9 14 0 13 7 3 1 1 15 1 9 9 0 13 2
29 9 0 16 1 9 16 3 9 13 13 0 13 16 9 9 1 9 9 9 13 7 9 9 1 9 9 0 13 2
14 9 0 13 9 9 0 1 9 0 0 9 0 13 2
20 0 9 0 9 0 9 13 7 1 9 1 9 0 2 9 7 9 0 13 2
35 9 9 3 12 9 9 14 1 9 1 15 9 9 13 7 13 16 9 10 9 9 2 9 9 9 0 9 0 14 1 9 0 9 13 2
29 9 3 14 15 1 9 0 9 2 9 13 7 9 0 7 9 0 14 9 13 9 7 9 16 9 9 9 13 2
15 7 15 2 9 12 0 9 0 0 9 9 1 9 13 2
34 15 10 9 14 12 9 3 1 9 7 9 9 13 7 13 16 15 12 9 1 9 9 1 13 7 3 3 15 14 13 1 9 13 2
13 9 9 2 9 3 1 7 1 10 9 9 13 2
14 12 7 12 12 9 9 13 7 12 12 9 0 13 2
51 16 10 9 2 15 16 1 9 9 9 9 13 13 2 15 3 9 16 1 9 1 9 0 2 9 1 9 0 9 13 2 1 10 9 12 1 9 0 13 7 13 2 9 9 2 9 9 3 14 13 2
19 7 15 16 9 9 13 15 0 13 0 13 13 2 9 1 9 15 13 2
60 9 0 2 9 0 16 1 9 13 13 2 7 15 9 13 0 16 12 1 0 9 14 1 9 9 9 7 9 9 1 9 15 13 13 3 9 1 15 13 2 0 13 16 13 9 9 15 1 3 13 16 15 9 9 0 13 7 9 13 2
20 7 16 1 9 15 9 13 2 13 2 9 9 2 7 9 3 14 3 13 2
16 9 0 9 0 0 13 2 9 2 10 9 9 9 3 13 2
19 7 15 16 3 1 9 7 9 9 1 9 9 0 13 13 13 2 6 2
11 12 9 13 16 15 16 1 15 9 13 2
14 7 15 13 2 9 9 0 15 13 9 0 13 13 2
11 0 9 12 13 2 15 9 9 14 13 2
6 1 9 13 2 6 2
9 13 2 9 9 9 14 16 13 2
4 13 2 6 2
10 10 12 13 1 9 7 9 0 13 2
40 16 9 1 9 1 9 9 9 9 13 2 13 2 9 0 2 9 13 16 12 12 9 9 0 1 9 13 16 9 9 13 7 9 9 1 9 9 9 13 2
60 15 16 9 0 9 9 9 13 9 9 1 10 9 2 1 9 0 9 9 9 9 9 13 16 1 9 15 9 7 9 9 13 2 9 12 9 2 12 9 2 2 1 3 12 9 9 13 16 1 9 9 10 9 2 0 1 9 15 13 2
27 3 16 9 9 3 13 2 3 10 9 0 2 9 15 13 12 9 13 2 7 1 9 0 9 9 13 2
64 3 9 16 9 9 2 1 9 0 9 9 13 16 15 9 1 10 9 7 9 13 0 13 7 3 9 9 2 9 9 9 9 9 9 9 9 2 9 13 13 16 10 9 9 9 9 9 15 13 15 1 10 9 7 10 3 13 0 13 1 15 9 13 2
54 9 16 2 3 16 9 9 9 0 7 9 9 16 1 9 15 1 9 13 2 13 1 10 9 0 9 13 2 1 9 15 7 9 15 13 9 1 9 9 1 9 2 9 9 13 1 10 9 2 1 9 15 3 2
59 9 1 10 9 13 16 15 12 9 13 1 9 9 15 16 9 0 13 7 9 0 13 2 7 9 3 13 7 9 3 13 7 9 9 15 13 2 7 9 12 9 9 9 1 9 1 9 13 7 15 12 9 1 10 9 7 9 13 2
47 10 9 9 9 7 9 12 9 0 13 1 9 12 9 0 1 9 2 7 9 12 9 0 13 12 9 0 1 9 9 2 7 1 3 16 9 1 9 9 13 13 9 1 9 9 13 2
11 15 13 2 3 1 9 9 1 9 13 2
14 12 9 9 14 13 1 9 15 1 9 9 0 13 2
31 0 9 1 9 9 9 15 2 7 0 9 1 9 0 15 2 7 12 12 9 9 9 0 16 1 15 9 13 16 13 2
26 15 3 13 16 9 9 9 3 0 16 15 9 15 14 16 1 9 7 7 1 9 13 13 0 13 2
46 15 9 14 0 13 7 9 15 14 13 16 15 14 1 9 15 1 9 13 2 7 9 16 1 0 15 12 9 9 9 9 2 0 9 15 14 9 13 7 1 10 9 0 9 13 2
38 15 3 1 9 9 13 2 7 1 9 9 9 15 14 1 9 15 1 15 7 15 9 13 9 3 1 9 9 0 1 9 13 2 7 3 9 13 2
2 3 2
40 9 15 13 16 9 9 9 15 9 3 2 16 3 1 9 2 1 9 9 9 9 2 9 9 9 2 1 9 1 9 9 13 7 1 9 1 9 13 13 2
151 15 1 9 9 2 1 9 13 2 15 2 1 3 13 16 9 13 7 9 9 13 2 10 12 12 9 2 15 2 1 9 9 12 9 3 9 2 9 1 9 13 7 1 3 13 7 9 9 12 9 13 13 9 9 9 2 9 2 16 1 9 9 3 9 7 9 13 7 9 13 7 7 9 9 13 7 7 9 7 9 13 7 9 7 9 7 9 2 3 0 9 13 12 9 0 1 9 0 2 0 2 16 12 9 9 1 9 15 13 2 7 9 16 1 10 9 7 9 1 9 15 9 9 14 9 13 0 13 7 9 16 0 7 0 1 9 9 13 2 3 9 7 9 14 1 13 1 9 9 13 2
33 1 9 15 7 10 9 16 1 9 0 9 3 13 7 0 1 9 9 16 9 12 9 0 13 13 9 15 3 7 0 16 13 2
55 1 1 15 2 16 9 16 9 3 13 2 9 0 1 10 9 9 9 16 1 3 15 13 9 1 9 9 13 16 1 9 9 10 9 0 2 9 1 9 15 7 15 13 7 9 1 9 15 7 15 13 9 9 13 2
18 3 13 2 15 3 13 16 9 15 14 1 9 13 7 9 15 14 2
31 1 9 15 7 1 9 9 9 9 9 2 10 9 9 13 2 7 0 13 3 1 9 9 14 3 16 3 13 0 13 2
49 15 16 13 9 9 15 13 7 15 13 9 15 13 16 9 1 9 9 13 9 15 15 13 2 12 9 3 16 9 1 9 9 7 9 1 9 13 2 13 1 9 0 9 1 9 7 9 13 2
71 9 0 3 0 7 0 13 1 9 9 7 9 0 0 1 12 9 2 0 7 0 7 0 15 14 1 9 9 13 2 7 1 15 1 1 9 9 9 7 9 7 1 1 9 0 9 1 9 13 7 3 1 9 12 9 9 2 9 1 9 9 13 2 9 9 2 1 9 9 13 2
11 9 0 9 13 7 13 2 9 2 9 2
35 9 9 1 9 1 9 13 7 13 2 3 2 9 10 9 13 7 15 9 9 9 13 2 7 13 3 10 9 9 15 1 3 9 13 2
9 9 15 13 2 7 9 15 13 2
27 1 9 7 9 4 13 1 1 15 2 15 3 13 16 9 13 16 9 1 9 9 13 16 10 9 13 2
66 0 1 15 2 9 9 15 2 1 9 12 0 2 9 13 13 1 9 9 12 9 3 7 9 7 9 9 9 12 9 3 7 9 7 9 9 7 9 12 9 3 9 13 10 9 14 16 15 13 1 9 10 9 12 9 0 15 13 16 9 9 7 9 0 13 2
87 1 1 15 15 2 16 9 13 9 13 2 3 13 16 9 9 9 9 9 9 12 0 0 14 13 16 12 7 12 9 15 14 1 9 13 7 12 7 12 9 3 16 10 9 16 15 3 12 12 0 13 12 0 2 12 0 12 9 3 1 9 0 0 2 1 9 9 13 7 1 9 7 9 13 7 10 9 12 9 9 1 10 9 0 13 13 2
26 15 13 9 15 14 13 2 7 15 1 0 9 3 0 9 1 9 9 13 16 13 9 13 7 3 2
40 9 15 15 16 9 0 13 9 13 15 16 13 2 7 15 7 13 9 13 7 13 15 10 9 16 15 1 9 9 1 10 9 13 9 13 1 9 10 9 2
5 15 9 9 13 2
24 13 16 3 9 9 15 0 13 2 16 15 1 9 0 0 9 13 2 7 9 1 9 13 2
47 0 13 16 12 9 9 13 2 15 3 1 10 9 0 9 13 16 10 9 12 9 1 9 9 13 2 7 0 1 15 9 13 16 10 9 0 13 7 0 2 7 10 9 9 9 13 2
72 9 9 0 13 16 3 0 13 1 9 9 9 7 9 9 7 9 9 7 0 1 15 9 9 3 9 2 7 3 9 15 14 3 9 16 3 0 13 1 9 0 16 9 1 9 13 13 13 9 13 7 3 9 7 9 9 0 13 16 9 3 9 10 9 14 9 13 2 3 2 3 2
12 3 7 9 13 13 0 13 9 3 13 13 2
31 1 1 15 2 10 9 2 10 9 9 2 10 9 2 10 9 0 9 9 13 7 9 13 7 1 9 0 13 13 13 2
26 9 9 13 9 9 9 9 9 14 2 12 9 0 0 1 9 15 13 16 9 9 9 15 9 13 2
7 15 9 9 9 0 13 2
25 10 9 3 12 9 1 15 1 9 13 13 7 9 15 16 0 13 7 4 0 15 1 9 13 2
41 9 2 16 9 9 13 3 9 9 14 13 2 7 16 9 9 9 9 7 9 14 13 7 3 12 9 3 13 3 9 14 0 13 7 9 13 9 3 9 13 2
42 12 9 9 1 9 9 9 9 9 13 2 9 1 0 9 13 7 9 13 2 7 9 0 13 2 9 9 13 7 3 13 2 9 9 3 15 7 9 15 14 13 2
38 9 1 9 9 13 2 9 2 10 9 7 3 9 15 14 15 0 13 1 9 13 2 7 9 13 16 9 13 10 9 14 1 15 13 3 0 13 2
10 1 10 9 10 9 14 15 9 13 2
14 3 2 15 12 2 12 9 16 3 13 9 0 13 2
24 15 4 13 2 7 15 4 13 2 3 4 1 9 10 0 9 9 16 9 13 9 13 13 2
19 9 16 0 13 2 9 16 3 1 10 9 0 9 2 3 9 0 13 2
8 15 9 14 13 7 4 13 2
69 10 9 0 1 10 9 12 0 7 1 10 9 0 0 3 15 13 16 1 9 9 9 9 1 9 0 0 13 9 1 10 9 7 9 1 15 16 13 2 16 12 12 12 9 0 9 9 9 0 2 0 13 7 2 10 9 1 9 0 13 2 9 16 9 0 1 9 13 2
109 9 3 14 2 1 10 9 0 2 7 10 9 0 1 10 9 2 3 15 13 13 16 1 9 0 0 13 9 14 1 9 9 13 9 15 13 16 9 10 9 1 12 12 7 12 12 13 1 9 16 0 13 1 9 9 9 9 2 15 14 3 13 2 7 1 15 15 10 12 7 12 12 9 14 12 12 9 13 7 1 9 15 12 12 12 13 1 9 7 9 13 7 12 9 16 12 12 12 13 9 9 13 16 9 15 14 0 13 2
36 10 9 9 15 13 2 7 10 9 9 15 13 2 7 15 9 7 1 9 9 15 9 2 9 9 0 13 2 3 1 9 9 9 0 13 2
44 9 1 15 13 7 1 9 9 9 9 0 7 0 2 1 1 10 9 16 3 13 2 10 9 0 9 16 3 9 0 9 13 7 2 3 13 1 9 9 9 1 9 13 2
81 9 1 9 0 1 9 9 13 16 8 9 9 9 13 2 9 0 7 0 0 1 9 13 16 1 0 12 9 9 9 9 9 3 3 0 13 16 12 9 13 9 0 9 0 9 13 7 16 9 0 13 7 9 0 2 3 3 10 9 7 9 9 16 9 7 9 7 2 13 2 9 14 13 7 9 13 7 3 9 13 2
27 7 9 9 13 16 1 9 9 13 7 13 13 9 9 9 0 4 13 3 16 9 9 7 9 13 13 2
70 9 15 9 1 10 9 13 16 16 9 3 13 7 1 9 13 7 9 7 9 0 9 9 7 9 7 9 1 3 13 15 16 9 7 9 13 0 13 2 7 16 9 9 13 13 2 15 9 0 13 2 9 9 9 2 16 7 9 13 1 9 2 1 13 10 9 16 9 13 2
103 1 9 13 16 1 9 9 0 16 0 1 9 1 9 9 13 7 9 1 9 15 9 13 13 1 9 9 12 9 9 9 0 13 1 9 2 9 9 0 9 16 16 9 9 9 2 16 9 9 9 9 13 7 9 15 1 9 13 9 7 9 7 0 7 0 7 15 9 9 1 15 9 13 7 1 9 4 13 16 15 9 0 16 13 1 10 9 2 9 16 2 9 2 2 15 16 13 1 9 12 9 0 2
7 9 15 1 9 9 13 2
71 7 16 9 9 13 7 9 13 3 13 16 9 9 9 0 13 7 9 1 9 9 13 1 10 9 13 16 1 9 9 9 9 2 1 9 9 9 2 9 9 9 1 12 9 0 9 13 16 12 9 1 9 9 0 12 3 1 9 16 9 9 9 9 9 9 9 1 9 9 13 2
32 1 10 9 1 10 9 1 3 1 9 9 2 10 9 9 0 13 16 2 1 9 9 9 13 2 9 9 9 0 4 13 2
96 15 1 9 10 9 2 1 9 9 9 1 9 9 7 9 16 12 9 0 9 13 1 9 0 13 2 9 9 2 9 9 2 9 13 15 1 9 13 16 9 9 9 14 1 9 13 7 9 13 16 9 9 1 9 9 13 2 7 10 9 14 1 15 9 13 16 9 12 12 9 1 9 9 0 15 9 1 9 9 2 9 9 1 15 0 13 7 1 10 9 3 0 1 9 13 2
17 13 9 13 1 9 9 16 15 14 1 15 13 1 9 7 9 2
81 7 9 1 9 2 3 15 1 10 9 1 3 9 1 15 9 13 13 7 9 0 16 15 13 13 10 9 1 10 9 7 9 0 15 13 7 9 16 15 13 13 1 15 9 9 15 14 13 2 7 9 14 16 1 9 9 13 13 15 1 9 15 13 2 7 10 9 3 1 9 15 1 2 3 1 9 9 9 15 13 2
62 1 9 15 13 16 15 9 9 15 13 7 10 9 14 1 10 9 13 16 1 10 9 9 1 9 9 1 0 15 7 1 15 9 13 1 15 13 2 9 2 15 9 9 15 14 1 10 9 9 15 1 9 13 7 1 10 9 1 15 0 13 2
18 15 3 1 9 3 9 13 16 9 15 1 9 1 9 12 9 13 2
104 2 9 9 12 2 7 1 9 9 9 16 13 16 9 1 9 13 2 7 1 15 3 0 2 4 1 12 9 16 0 13 7 15 15 16 10 9 9 9 14 1 9 13 2 0 13 2 7 10 9 14 1 9 9 9 9 9 9 9 7 9 7 9 9 9 9 3 13 2 9 9 9 12 2 7 9 9 9 9 16 1 9 9 9 1 15 15 13 7 3 0 9 15 9 0 0 9 13 16 9 0 9 13 2
44 7 3 10 9 13 16 9 9 9 12 12 9 13 7 9 10 15 3 12 12 9 9 13 2 7 1 10 12 9 0 2 3 9 9 9 13 16 15 14 12 9 9 13 2
11 2 9 3 15 0 13 2 9 12 2 2
31 13 1 9 15 15 9 13 2 16 7 12 12 9 16 3 16 12 12 9 16 13 12 9 0 3 9 1 9 15 13 2
33 10 9 12 9 0 13 16 2 6 15 9 0 13 16 12 12 9 0 13 13 7 9 9 14 13 7 1 9 9 9 9 13 2
6 9 1 10 0 13 2
85 16 9 15 14 1 9 7 9 9 9 13 7 1 12 9 15 14 1 9 9 9 13 3 3 1 9 0 9 7 9 9 15 13 7 13 16 9 15 9 13 1 9 9 15 16 16 9 1 9 13 1 9 0 13 7 9 15 13 16 1 0 13 1 10 9 9 15 1 9 16 3 9 9 13 7 10 9 14 9 9 9 1 15 13 2
18 1 9 16 9 9 9 13 12 9 1 9 15 7 9 4 0 13 2
126 9 15 2 1 9 9 2 1 9 9 9 9 13 16 16 3 1 9 9 13 7 7 3 1 9 2 7 3 9 15 2 9 7 9 13 7 3 13 2 10 9 3 9 9 9 13 16 9 12 7 12 9 9 13 2 0 1 9 9 16 12 12 9 9 1 12 13 2 1 1 9 9 9 9 0 13 7 9 16 9 15 1 9 0 16 15 14 1 9 13 0 13 2 7 1 9 2 16 9 12 12 9 1 12 13 9 9 13 7 9 13 16 16 9 13 16 12 9 9 1 1 10 9 9 13 2
103 7 3 1 9 12 16 13 9 7 9 15 1 9 9 0 13 7 9 14 3 13 7 6 1 9 13 16 0 13 7 9 0 13 2 3 15 7 9 13 16 9 9 9 9 13 2 9 9 9 7 9 13 16 10 9 9 14 1 9 15 16 13 2 3 3 10 9 9 16 1 10 12 9 9 1 9 9 0 7 0 2 3 9 9 7 9 15 1 9 15 16 9 7 9 7 9 9 13 3 0 13 13 2
16 3 3 9 2 16 9 9 0 13 13 1 9 16 9 13 2
52 1 10 9 16 9 0 13 1 9 7 9 7 9 7 3 9 7 9 9 9 9 2 7 12 12 9 1 9 9 0 16 15 9 9 15 13 9 16 9 13 13 7 3 12 12 9 1 9 16 9 13 2
40 3 9 15 3 1 12 9 9 13 16 9 10 9 13 10 9 9 1 9 13 7 9 13 3 9 1 15 13 7 7 13 12 9 1 9 9 0 7 0 2
14 10 9 1 12 9 9 0 9 0 14 9 9 13 2
15 12 12 9 3 2 1 9 9 9 9 9 13 13 2 2
53 9 9 13 2 1 15 7 9 1 12 12 9 9 7 9 7 9 9 2 9 13 7 3 2 15 15 14 1 9 12 9 9 2 1 12 9 2 9 9 0 1 9 9 2 7 9 0 0 1 9 9 13 2
48 15 9 14 1 9 9 13 7 9 9 14 1 9 15 15 9 13 16 12 7 0 9 13 7 16 1 10 9 12 0 7 9 16 13 13 7 15 13 16 9 1 9 0 3 9 0 13 2
31 1 9 16 3 12 9 7 0 1 9 9 13 7 3 15 10 9 13 16 15 15 9 13 7 9 14 3 15 4 13 2
17 1 1 10 9 2 15 9 15 14 13 9 16 9 9 0 13 2
37 9 13 2 15 12 9 9 9 7 9 1 9 7 9 0 13 2 7 3 1 9 9 0 14 13 16 2 8 8 8 8 7 8 8 8 8 2
79 15 9 13 16 10 9 16 9 0 4 13 16 9 9 1 15 9 13 2 7 16 1 10 9 9 9 0 13 13 3 9 0 9 1 9 10 9 0 16 13 0 13 12 9 0 14 9 13 16 2 3 15 1 9 0 2 9 1 9 16 9 15 1 9 13 7 1 9 0 13 1 12 9 9 0 0 9 13 2
16 16 2 10 9 0 1 9 13 16 13 2 9 14 0 13 2
12 9 0 0 1 0 9 9 13 3 9 15 2
34 7 16 9 9 14 1 10 9 0 13 9 13 2 15 9 14 0 13 15 9 9 14 1 9 9 0 13 2 9 9 9 12 2 2
25 12 9 0 3 4 9 15 14 0 9 9 13 16 1 9 12 9 9 0 8 0 3 13 13 2
30 9 13 16 12 9 3 2 15 15 1 9 9 9 9 16 9 0 10 9 13 1 9 13 2 9 9 9 12 2 2
59 9 0 9 13 16 1 9 0 13 0 9 9 9 14 1 9 9 7 9 9 13 7 15 9 13 7 16 10 9 9 13 7 0 13 13 10 9 9 3 3 0 1 9 9 9 9 13 7 16 13 3 15 1 9 0 13 0 13 2
15 0 9 9 7 9 9 0 1 9 9 2 9 9 13 2
23 2 9 9 2 9 12 2 7 15 9 13 16 9 12 7 0 12 9 1 1 15 13 2
93 10 9 16 15 1 1 9 9 9 13 3 1 9 7 0 13 3 15 7 2 9 3 9 16 9 0 16 1 9 13 7 7 1 9 13 7 7 1 9 13 7 7 1 9 13 2 1 3 13 1 0 9 10 9 7 9 15 16 9 9 15 14 13 7 13 9 14 9 13 7 0 9 0 1 9 0 9 9 13 16 1 9 10 9 7 9 9 15 9 14 9 13 2
99 9 0 1 15 13 16 12 9 0 1 9 9 9 9 1 9 1 9 9 0 9 2 7 0 9 1 9 9 9 13 16 9 9 7 9 9 9 2 9 3 9 9 14 16 1 9 9 2 9 1 9 9 13 2 3 9 13 16 15 9 9 14 1 12 9 9 13 7 1 9 9 15 14 16 1 9 13 16 1 9 13 7 0 9 16 2 9 0 15 9 9 9 3 9 14 1 9 13 2
87 2 9 9 9 12 2 9 9 9 9 16 16 9 9 10 9 1 9 15 13 2 0 0 1 15 13 16 9 9 9 9 9 9 9 0 1 9 9 0 16 1 9 9 9 13 2 9 2 1 9 9 9 0 2 1 10 9 16 15 1 9 9 7 9 13 2 1 9 1 9 10 9 16 3 9 9 13 2 9 13 16 9 14 3 9 13 2
19 9 1 9 0 7 0 7 9 0 0 0 9 1 15 7 9 15 13 2
21 9 9 1 9 9 12 9 9 9 14 13 2 9 2 12 12 12 12 12 12 2
74 2 9 9 9 12 2 7 15 1 9 9 13 16 12 7 0 9 3 16 15 7 9 9 1 9 13 2 9 9 9 13 15 14 1 1 9 9 13 16 9 0 13 7 13 2 9 15 9 0 13 7 12 9 3 1 15 1 9 9 9 9 9 7 9 14 9 13 16 9 9 9 13 13 2
20 9 9 13 16 13 2 9 16 9 14 1 9 9 0 3 1 9 9 13 2
85 6 9 12 9 16 1 9 9 7 9 9 0 9 7 9 7 9 7 9 3 9 13 2 7 15 1 9 0 7 9 1 15 1 9 15 15 9 9 0 7 9 9 0 0 7 0 13 1 9 9 7 1 9 9 0 7 9 3 0 9 13 15 1 9 9 16 9 9 9 9 0 9 1 15 0 13 2 9 9 1 15 9 0 13 2
17 9 3 0 1 15 9 13 2 16 1 9 15 10 9 0 13 2
16 9 7 9 9 15 0 9 2 9 1 15 7 9 9 13 2
17 0 7 0 7 0 7 3 15 9 2 3 9 1 15 9 13 2
18 3 9 0 7 0 13 1 9 9 2 9 1 9 9 9 0 13 2
17 0 3 9 15 9 1 9 7 9 2 9 16 1 9 0 13 2
14 15 0 1 9 9 9 2 15 0 14 9 9 13 2
20 3 1 9 10 9 13 15 14 2 16 15 14 13 1 10 9 7 0 13 2
18 9 1 9 13 10 9 9 2 16 9 9 0 1 10 9 0 13 2
30 9 9 3 1 9 1 9 9 7 9 0 7 9 0 9 13 16 9 1 9 9 0 7 9 9 9 7 9 13 2
76 9 9 9 9 9 7 9 0 0 7 9 0 14 1 9 9 0 1 9 9 0 1 9 9 0 1 9 9 13 7 13 2 10 9 7 9 13 16 0 1 9 9 9 2 9 9 7 9 0 7 0 13 2 9 0 14 1 9 13 7 1 9 9 9 0 1 1 15 3 1 1 9 7 9 13 2
58 9 9 0 14 1 0 9 9 7 9 9 7 9 0 7 9 1 9 0 13 7 13 2 9 7 9 9 16 13 1 9 9 0 7 0 7 16 13 1 9 9 7 9 0 9 3 7 9 0 7 0 13 2 4 3 13 13 2
122 9 1 9 0 1 9 15 1 9 1 9 9 9 0 7 9 0 1 9 9 0 9 13 2 9 7 9 9 0 1 9 15 3 9 13 16 9 0 1 9 9 0 1 9 0 9 13 7 1 9 9 0 7 0 2 9 1 9 0 9 7 9 1 9 0 16 9 0 1 9 9 0 13 4 1 9 9 9 7 9 7 9 7 9 9 1 0 9 9 9 0 13 7 15 10 9 0 13 16 9 0 10 9 9 9 9 1 9 13 7 9 15 1 9 0 9 0 9 3 9 13 2
53 9 9 9 13 2 3 9 1 9 9 0 7 9 9 9 7 9 13 7 1 9 10 9 9 0 16 9 1 15 14 1 9 9 13 7 1 9 9 2 9 0 14 0 13 1 9 9 0 9 0 4 13 2
59 1 9 0 1 10 9 9 13 2 15 3 9 9 9 7 9 9 13 9 9 7 9 13 16 1 9 9 7 9 9 7 0 9 9 7 9 15 0 13 7 1 1 15 9 7 9 2 9 9 7 9 1 1 9 14 1 9 13 2
16 9 15 0 7 0 7 1 9 1 9 0 7 9 0 13 2
21 3 3 9 7 3 9 3 0 1 12 9 9 0 2 9 0 7 9 0 13 2
24 4 9 0 7 0 0 1 9 7 9 9 2 9 7 9 9 9 14 16 9 9 9 13 2
20 7 3 1 9 7 9 1 9 13 16 1 9 10 9 9 7 9 13 13 2
56 9 9 9 13 16 3 9 9 0 1 9 9 13 7 13 2 1 3 9 13 16 1 9 9 0 1 9 2 9 2 9 7 9 4 9 9 3 0 9 7 9 7 9 9 2 9 7 9 7 9 0 7 0 16 13 2
16 1 15 13 16 9 14 3 1 15 15 1 9 9 9 13 2
46 9 1 0 9 0 2 1 9 9 7 9 9 7 9 9 7 9 9 16 9 13 7 13 2 15 16 2 3 1 9 16 13 7 9 7 9 9 14 1 1 9 9 7 9 13 2
17 8 8 10 9 9 9 16 9 15 14 9 13 13 9 13 13 2
22 0 13 16 15 1 0 9 7 9 3 0 13 1 9 7 9 1 9 7 9 13 2
28 16 15 9 13 7 15 13 13 9 15 14 1 9 0 7 0 0 13 2 9 13 2 16 15 15 0 13 2
7 15 13 2 6 0 13 2
9 13 2 3 8 8 9 3 13 2
6 9 1 9 9 13 2
7 9 13 2 15 9 13 2
17 9 3 9 13 16 13 3 1 15 15 9 14 1 3 9 13 2
19 7 9 9 7 9 1 9 8 9 2 9 2 0 13 1 9 9 13 2
19 9 8 8 9 9 13 16 12 9 0 9 9 9 3 13 7 9 13 2
9 9 8 9 9 9 14 9 13 2
14 13 2 10 9 9 15 9 13 7 15 16 9 13 2
20 1 9 7 9 15 1 9 16 9 1 9 1 9 13 13 9 7 9 13 2
23 9 1 9 2 10 9 9 8 9 13 2 16 16 2 9 9 14 9 7 9 0 13 2
17 16 2 1 9 9 9 2 9 2 9 1 10 9 0 0 13 2
19 8 8 9 1 9 0 9 16 1 9 15 9 13 7 1 9 9 13 2
38 9 16 1 9 1 9 9 7 9 0 13 2 9 8 9 14 9 9 13 7 9 14 9 9 2 9 1 9 9 16 13 7 13 2 6 9 9 2
9 15 9 9 7 9 0 14 13 2
5 15 9 9 13 2
10 16 13 9 3 1 15 9 9 13 2
20 15 16 9 13 7 13 2 10 9 9 15 14 1 9 13 7 1 9 13 2
8 13 2 1 9 16 15 13 2
13 9 1 15 13 2 15 0 7 0 10 9 13 2
3 3 13 2
30 9 1 9 0 16 9 13 16 1 9 9 9 7 9 15 9 15 1 1 9 9 13 16 13 9 1 9 9 13 2
28 9 9 0 9 7 9 16 12 9 0 13 2 12 9 9 9 14 9 13 7 1 9 9 0 9 9 13 2
17 12 9 0 16 4 13 16 9 0 15 9 9 7 9 9 13 2
6 1 9 9 9 13 2
13 1 9 16 9 9 2 10 9 0 0 0 13 2
15 9 16 1 9 13 16 9 9 0 1 9 9 13 13 2
8 9 0 9 7 3 9 13 2
31 9 9 9 2 9 2 1 9 7 7 0 1 9 9 2 9 2 7 9 16 9 14 3 13 2 9 0 9 9 13 2
18 9 1 9 9 9 13 16 9 13 7 9 14 1 9 9 9 13 2
11 9 9 14 1 9 1 9 9 0 13 2
15 9 1 1 15 13 7 13 10 9 9 9 9 0 13 2
11 9 9 1 9 13 7 9 14 9 13 2
14 9 1 9 13 16 9 14 1 9 9 9 13 13 2
9 9 10 9 14 1 9 0 13 2
35 9 8 9 1 9 9 1 13 7 9 13 16 1 9 9 2 9 7 9 9 13 7 15 1 9 9 2 9 2 9 7 9 0 13 2
20 7 13 9 14 9 1 9 13 16 3 9 13 2 9 0 1 9 15 13 2
17 9 13 2 10 9 10 9 13 16 10 9 1 15 0 13 13 2
31 2 9 9 9 12 2 9 9 9 2 9 2 16 1 1 9 13 13 2 9 15 14 1 9 1 9 15 9 0 13 2
5 9 13 2 9 2
2 9 2
4 9 0 13 2
8 9 16 1 9 9 9 13 2
11 9 13 2 15 13 10 9 1 9 13 2
3 0 13 2
7 10 9 1 10 9 13 2
7 9 7 9 16 9 13 2
19 16 9 7 9 13 13 9 9 14 1 9 9 13 2 9 0 9 13 2
60 9 1 9 9 14 1 9 13 7 15 1 9 9 2 9 0 7 0 7 0 16 9 9 0 14 0 13 2 1 9 9 16 3 1 9 7 9 15 9 13 2 9 0 9 9 3 9 0 1 9 16 1 9 1 13 1 9 0 13 2
16 9 9 13 2 9 9 9 1 9 14 15 15 1 9 13 2
8 1 9 12 0 1 9 13 2
16 9 13 2 9 2 9 7 9 7 9 14 1 1 15 13 2
16 1 9 9 13 16 10 9 1 1 15 13 9 0 0 13 2
7 10 9 9 9 9 13 2
11 10 9 1 9 16 9 1 9 13 13 2
12 3 1 10 9 13 2 9 15 3 13 13 2
10 0 9 13 7 9 15 14 3 13 2
22 1 9 15 13 16 3 1 15 15 9 14 9 13 15 16 0 7 0 9 9 13 2
14 15 16 9 7 9 14 9 13 15 9 9 15 13 2
12 15 1 1 15 16 9 9 13 7 9 0 2
14 9 0 9 0 1 9 9 7 9 9 1 9 13 2
7 3 0 9 9 9 13 2
12 1 9 9 9 2 9 2 1 9 9 13 2
36 9 2 3 1 9 9 9 2 9 2 9 13 7 1 9 9 13 16 1 9 13 7 3 16 9 9 14 1 9 13 2 1 9 9 13 2
25 1 9 9 9 7 9 9 16 1 9 9 13 7 13 2 15 13 16 15 9 9 7 9 13 2
34 9 1 9 9 7 9 9 7 9 7 15 15 7 9 9 7 9 9 14 9 13 7 1 9 13 16 1 9 13 7 9 13 13 2
26 9 15 3 10 9 14 13 16 1 9 9 3 15 7 9 16 1 9 13 2 9 9 1 9 13 2
27 9 2 9 1 9 9 1 9 14 0 13 7 13 2 10 9 1 9 9 0 7 0 7 0 9 13 2
20 1 10 9 16 9 2 9 7 9 7 9 13 2 9 1 9 9 9 13 2
20 16 10 9 2 9 15 9 13 2 0 13 15 3 1 9 15 1 9 13 2
18 9 3 1 9 9 2 3 9 1 9 1 9 1 9 9 0 13 2
11 1 9 0 9 7 9 16 1 15 13 2
11 1 9 1 9 1 9 12 0 9 13 2
21 9 9 9 9 2 9 2 3 16 9 13 2 9 1 9 9 7 9 9 13 2
26 9 3 1 9 9 9 2 9 2 1 9 13 2 13 1 9 2 9 2 9 0 1 9 13 13 2
11 9 13 2 15 15 0 13 7 0 13 2
14 9 13 2 9 2 9 2 0 9 15 13 16 13 2
24 8 9 13 2 9 9 0 1 15 13 16 9 4 1 1 9 9 15 15 14 1 9 13 2
17 9 1 8 9 13 2 3 3 9 9 15 2 9 2 15 13 2
20 8 9 13 2 7 1 3 7 9 8 9 9 2 9 2 14 13 15 13 2
8 9 9 0 9 3 0 13 2
28 15 1 9 9 13 9 7 9 9 9 9 2 9 2 14 9 13 2 16 16 13 9 9 3 9 3 13 2
14 0 15 7 13 9 9 9 2 9 2 14 0 13 2
31 9 1 1 9 9 2 9 2 3 9 7 9 9 1 10 9 16 15 14 9 9 0 9 9 13 9 0 7 0 13 2
19 9 13 1 0 9 15 2 9 7 9 9 9 2 9 2 1 9 13 2
6 15 9 9 0 13 2
27 9 13 15 14 15 9 7 9 13 2 3 0 7 0 13 7 15 14 16 15 3 13 9 7 9 13 2
13 0 1 15 7 9 9 1 9 7 9 9 13 2
8 15 3 13 1 9 9 13 2
25 9 9 0 9 9 1 9 9 0 0 10 9 9 13 2 1 9 0 9 9 2 9 0 13 2
44 9 9 9 9 1 9 0 13 9 3 9 9 15 14 1 9 9 0 9 0 9 9 13 7 1 10 9 9 13 16 4 9 9 9 14 1 0 9 9 0 2 9 13 2
54 15 9 13 2 9 1 9 1 9 15 2 9 1 9 0 13 2 4 9 15 14 9 1 9 7 9 13 16 3 15 1 15 1 9 7 9 1 9 9 7 9 0 1 9 0 7 9 0 0 2 9 0 13 2
21 9 9 13 2 9 15 1 9 0 7 9 0 0 7 0 9 7 9 9 13 2
47 9 9 0 9 13 2 4 1 9 1 9 15 9 13 7 1 9 9 15 15 7 9 0 16 1 9 0 13 2 9 7 9 9 14 9 7 9 0 14 1 9 7 9 9 9 13 2
71 15 13 2 10 9 13 16 1 9 1 10 9 4 9 0 7 0 15 15 14 9 13 7 9 9 9 14 1 9 9 0 7 9 9 0 1 9 9 15 9 13 7 1 7 15 9 0 2 0 7 0 15 14 1 9 0 0 13 2 1 9 1 9 0 9 15 1 0 4 13 2
35 9 1 9 9 16 1 12 9 3 9 13 1 0 9 7 1 9 9 9 9 0 9 1 9 9 0 1 9 10 9 1 9 13 13 2
31 10 9 16 0 1 12 9 9 0 1 9 1 9 9 9 13 1 0 9 9 1 9 9 1 9 9 1 9 13 13 2
36 1 9 9 0 2 9 0 3 1 9 9 1 9 0 2 9 0 2 7 1 9 9 15 7 9 15 9 1 9 14 1 9 9 13 13 2
31 1 9 9 0 9 9 0 9 2 1 9 0 1 10 9 9 0 0 16 1 9 9 0 7 0 13 1 9 1 13 2
34 10 9 0 16 0 1 12 9 3 1 9 13 2 1 9 12 2 12 9 7 1 9 9 1 9 0 9 0 9 1 9 9 13 2
37 0 1 9 10 9 2 9 0 0 1 9 0 9 9 2 1 1 9 9 7 0 9 9 1 9 9 9 0 1 9 0 1 9 1 4 13 2
37 10 9 0 16 9 15 1 0 1 12 9 13 2 0 1 9 0 3 1 9 0 7 9 9 9 0 14 1 9 0 1 9 9 9 9 13 2
17 9 0 1 9 12 0 1 9 1 9 9 9 9 1 9 13 2
31 12 9 0 0 1 9 9 9 0 12 9 2 9 2 0 9 9 1 9 0 9 9 2 1 9 9 9 12 9 13 2
19 2 9 2 3 1 9 9 0 9 9 0 9 0 9 9 13 13 13 2
31 9 9 9 2 12 1 0 9 0 13 16 9 9 1 9 9 10 9 2 9 9 1 9 1 9 9 9 14 9 13 2
26 1 9 9 0 9 2 9 2 1 9 16 1 9 9 10 9 9 13 1 9 9 9 9 13 13 2
47 9 9 9 9 13 16 1 9 9 7 1 9 9 1 9 0 13 7 2 10 9 1 3 1 9 0 1 9 9 9 2 9 9 2 9 9 2 9 9 2 9 9 9 0 13 13 2
19 10 9 16 2 1 12 9 9 9 1 9 9 1 9 9 13 13 13 2
23 3 1 9 9 9 2 9 9 1 9 9 9 2 9 2 9 7 9 9 0 0 13 2
15 3 1 9 0 0 1 12 9 1 10 9 9 13 13 2
50 16 2 9 9 7 9 9 9 7 9 9 7 9 9 1 10 9 1 9 9 9 9 0 1 9 9 7 9 9 0 9 7 9 1 9 9 9 13 7 10 1 9 0 9 9 9 1 9 13 2
18 0 9 9 0 9 0 9 9 1 12 1 12 9 9 3 0 13 2
57 9 9 9 10 9 2 1 9 9 9 9 9 13 16 9 9 15 14 3 1 9 1 9 0 9 9 13 7 12 9 0 1 9 2 9 2 2 2 9 2 2 2 9 2 2 9 16 0 15 13 7 9 9 9 13 13 2
7 12 9 9 1 9 9 9
32 9 9 9 0 1 9 0 9 9 0 1 9 9 0 9 7 9 9 9 7 9 1 9 9 2 9 1 9 9 9 13 2
53 10 9 1 9 0 9 1 9 0 13 7 9 15 0 9 9 9 2 9 2 1 9 9 1 9 9 2 9 9 1 9 9 9 7 9 9 1 9 9 9 9 9 9 1 9 9 1 9 9 2 4 13 2
7 9 1 9 9 9 13 2
11 9 9 1 9 1 9 9 1 9 13 2
45 1 10 9 9 0 3 9 9 1 1 9 9 0 1 9 2 9 9 9 1 9 9 7 9 9 7 9 9 9 1 1 9 9 0 1 9 7 9 15 1 9 9 4 13 2
42 1 10 9 9 9 9 2 9 9 9 2 9 9 9 2 9 9 9 2 9 9 2 9 9 7 9 9 1 9 9 13 16 1 1 9 0 9 1 9 4 13 2
11 9 9 1 9 1 12 9 9 4 13 2
8 9 9 0 7 0 9 13 2
20 9 0 15 1 9 0 2 9 9 0 14 3 7 3 1 9 0 13 13 2
16 9 3 1 9 9 1 9 9 0 1 9 9 9 9 13 2
26 9 9 0 9 1 9 9 13 2 9 0 12 12 7 12 9 0 7 0 1 9 10 9 9 13 2
25 9 9 13 2 12 12 7 12 9 1 9 0 1 9 7 9 9 0 13 7 9 9 0 13 2
42 9 2 9 0 7 0 0 7 9 10 9 14 1 9 0 2 12 12 7 12 9 9 9 13 7 13 2 1 10 9 12 12 7 12 9 9 0 1 9 0 13 2
25 15 13 2 1 9 12 2 9 9 0 7 0 0 1 0 7 0 12 12 7 12 9 13 13 2
28 9 0 9 1 9 9 12 9 9 13 7 0 1 9 0 2 9 9 0 2 9 7 0 9 1 9 13 2
28 9 7 9 0 9 0 9 9 9 9 7 9 13 16 3 1 9 9 0 1 9 9 7 9 9 13 13 2
25 9 9 1 9 0 9 9 9 13 2 9 9 1 9 0 9 3 1 10 9 1 9 1 13 2
33 9 9 9 1 13 7 9 1 9 1 9 13 2 1 9 10 9 2 12 9 9 7 12 9 9 0 1 1 10 9 9 13 2
23 15 9 9 7 9 9 14 12 12 9 7 9 9 7 9 14 9 12 12 9 9 13 2
43 9 1 9 1 15 16 9 9 0 9 9 0 13 7 3 1 9 9 16 13 0 13 2 13 2 1 9 1 10 9 9 4 3 9 13 7 12 9 3 13 0 13 2
21 15 13 2 1 9 1 9 9 0 1 9 9 0 7 9 9 9 0 13 13 2
32 9 9 0 9 9 13 2 1 9 9 1 0 9 9 2 12 12 7 12 12 9 1 9 0 0 7 9 10 9 9 13 2
39 9 9 13 2 1 10 9 16 1 9 9 9 0 9 13 12 12 7 12 9 1 9 0 0 9 13 7 12 12 9 1 9 16 9 7 9 13 13 2
20 15 13 2 1 1 15 1 9 9 0 12 9 0 16 1 10 9 13 13 2
29 9 13 2 9 0 10 9 1 3 1 9 10 9 1 9 9 9 1 12 9 1 9 1 12 9 0 13 13 2
29 15 9 9 9 1 9 0 10 9 14 12 9 1 10 9 13 7 15 14 3 0 1 9 1 0 9 9 13 2
18 1 9 9 12 12 9 9 7 12 12 7 12 12 9 9 9 13 2
34 9 9 9 9 13 2 1 9 9 9 9 2 15 3 9 12 9 9 9 2 9 14 0 13 16 4 12 9 1 15 14 9 13 2
35 9 9 9 2 16 1 9 9 9 9 9 13 2 13 2 9 12 0 9 9 1 9 9 0 3 1 9 9 7 1 9 16 0 13 2
19 15 13 2 15 1 9 7 9 9 9 9 10 9 15 14 1 9 13 2
30 9 13 2 1 9 9 1 9 9 9 9 1 9 9 2 9 0 1 9 12 9 9 9 1 9 14 0 9 13 2
35 15 1 9 15 16 9 0 9 9 10 9 1 9 13 2 13 2 9 0 15 9 9 3 7 9 0 16 1 9 12 1 9 4 13 2
14 15 9 9 9 9 14 0 1 12 12 9 9 13 2
26 9 9 1 12 0 9 9 9 2 12 1 9 0 7 0 9 2 3 1 9 9 0 1 9 13 2
34 9 9 0 9 2 13 2 1 9 10 9 1 9 12 1 9 9 0 2 3 9 0 1 9 7 9 10 9 1 9 13 13 13 2
34 9 9 13 2 9 9 3 0 1 9 10 9 2 1 9 0 1 9 9 13 7 1 9 0 1 9 9 9 9 3 9 13 13 2
34 1 9 15 2 9 1 10 9 1 9 0 13 13 7 9 9 0 15 2 3 1 9 12 0 0 1 9 9 9 9 9 13 13 2
24 9 9 0 9 13 16 9 0 10 9 1 9 3 1 9 7 1 9 0 1 9 9 13 2
26 9 10 9 1 9 0 7 1 9 0 13 7 1 9 0 1 12 12 9 2 3 10 9 9 13 2
22 0 9 9 9 0 9 16 1 9 9 13 13 3 1 12 9 1 9 15 9 13 2
40 9 9 0 9 9 9 10 9 14 9 9 9 1 9 9 0 7 0 1 9 2 9 7 9 9 7 7 9 1 0 9 0 1 9 9 9 0 9 13 2
26 9 9 9 9 0 9 14 1 9 9 3 9 2 9 2 9 2 9 7 9 2 3 0 9 13 2
76 15 13 2 1 9 7 9 12 2 12 9 9 9 9 14 1 9 13 3 12 9 9 9 9 1 9 15 9 13 7 1 12 12 9 9 16 1 9 9 13 9 1 9 12 12 9 1 9 2 9 9 9 0 10 9 14 1 9 13 7 1 12 12 9 9 9 0 9 12 12 9 9 9 9 13 2
16 1 10 9 12 9 1 9 2 9 7 9 10 9 9 13 2
30 9 0 2 9 2 9 0 9 9 9 2 9 9 9 2 9 0 7 9 7 9 1 9 1 9 1 10 9 13 2
21 1 9 9 9 1 9 0 7 9 0 9 2 9 0 7 9 16 1 9 13 2
8 9 16 1 9 0 0 13 2
40 9 2 1 9 9 0 1 9 2 9 12 12 9 9 9 0 9 0 12 9 9 13 7 9 9 9 0 13 7 9 9 1 9 9 2 9 9 0 13 2
14 9 7 9 0 9 9 0 2 10 9 0 15 13 2
78 16 9 1 9 9 9 0 9 9 13 16 13 2 16 9 1 9 1 9 9 0 9 16 1 9 12 9 0 0 9 15 9 7 9 1 9 9 7 1 9 13 2 9 13 2 16 13 2 0 1 9 7 9 4 13 16 1 9 9 0 7 9 1 9 2 9 7 9 2 1 9 9 13 2 1 9 13 2
20 9 1 9 1 9 1 9 9 2 1 9 9 9 15 1 9 0 9 13 2
16 9 9 1 1 12 9 0 2 1 9 9 0 9 9 13 2
4 9 2 9 2
34 9 9 1 9 9 9 1 9 9 9 0 1 9 13 16 0 1 9 0 9 13 7 9 10 9 1 9 0 14 16 1 9 13 2
52 9 9 9 9 9 13 2 3 9 9 9 9 14 1 9 9 15 9 4 13 16 1 9 15 1 9 16 9 9 13 9 13 13 9 0 1 9 9 14 1 9 9 9 16 9 7 9 9 13 9 13 2
36 1 10 9 13 13 2 9 0 1 9 9 13 16 9 0 4 13 3 7 9 9 9 13 1 9 9 9 9 13 16 1 9 9 13 13 2
41 9 16 9 9 9 7 9 9 9 1 9 13 16 9 1 12 9 9 9 1 9 7 9 13 16 1 10 12 9 9 9 9 9 9 10 12 9 14 13 13 2
45 9 9 13 2 16 9 13 9 0 9 7 9 14 9 13 15 14 1 12 9 0 16 1 9 1 10 9 1 9 13 0 4 13 7 16 9 1 10 9 1 9 0 0 13 2
23 9 1 9 16 1 9 1 9 15 9 13 13 9 0 13 16 1 9 0 9 13 13 2
41 16 1 9 0 9 9 7 9 1 9 0 15 3 1 9 9 13 13 7 9 0 1 9 0 1 9 0 16 15 16 9 0 13 1 9 9 9 13 13 13 2
10 12 9 0 1 9 9 9 1 13 2
36 1 9 0 9 9 9 9 9 7 9 16 1 9 9 13 2 9 9 12 9 1 9 9 15 1 9 1 9 15 1 9 10 9 1 13 2
31 1 0 9 10 9 2 9 9 0 7 0 0 13 7 9 9 7 9 9 1 10 12 9 13 9 9 14 9 9 13 2
12 1 9 0 2 9 9 1 9 0 9 13 2
33 1 9 0 9 0 14 3 12 1 12 0 13 7 1 9 0 1 1 9 0 15 12 1 12 0 13 7 1 9 9 9 13 2
42 1 9 0 2 9 9 1 9 0 9 0 15 14 3 12 1 12 9 13 7 1 9 0 1 1 9 9 0 12 1 12 9 14 0 13 7 1 9 9 1 13 2
24 1 0 9 10 9 9 9 7 9 9 9 9 0 7 0 9 15 1 9 1 9 15 13 2
9 12 9 1 9 9 1 9 13 2
31 9 9 9 1 9 0 1 9 16 1 9 0 9 1 9 0 7 9 0 0 13 2 9 12 9 9 7 12 9 13 2
45 1 10 9 16 1 9 9 0 13 7 9 9 1 9 13 2 9 9 1 9 16 1 9 0 13 13 2 1 1 9 9 1 9 1 9 0 0 13 7 1 9 9 9 13 2
13 16 9 9 0 9 0 1 9 9 9 0 13 2
30 1 1 9 9 0 9 0 9 1 9 2 9 9 9 0 9 9 0 9 9 1 9 0 1 9 0 14 9 13 2
37 1 10 9 16 9 3 1 9 12 9 1 12 9 1 9 9 9 9 0 0 13 2 9 0 9 0 9 15 1 9 12 9 1 9 0 13 2
32 1 9 9 9 1 9 2 12 9 9 9 9 16 13 9 15 9 13 2 1 10 9 13 2 9 1 12 9 9 4 13 2
48 0 9 1 9 9 9 1 9 7 9 0 9 1 13 7 13 1 9 9 9 13 16 15 0 1 9 9 1 9 15 13 7 9 16 1 15 13 13 7 0 10 9 1 9 15 0 13 2
22 15 0 9 13 16 9 1 9 9 12 9 0 9 0 7 0 1 3 9 9 13 2
16 9 1 9 9 7 9 0 1 9 1 9 9 9 9 13 2
4 9 2 9 2
19 9 12 1 0 9 9 16 0 1 9 13 2 1 12 9 3 0 13 2
23 9 0 13 2 9 9 9 9 9 16 1 9 9 9 9 13 2 9 10 9 13 13 2
27 10 9 16 9 9 15 12 2 12 9 13 1 9 12 9 3 1 9 0 1 12 12 9 9 13 13 2
16 15 0 9 15 14 9 1 9 7 9 9 0 9 13 13 2
24 9 9 3 3 9 9 9 13 7 9 0 16 9 13 7 1 9 9 0 9 0 16 13 2
46 0 3 13 16 9 16 0 13 2 9 9 9 7 9 7 9 9 0 14 9 9 0 13 2 9 13 16 1 9 1 10 9 9 13 2 15 1 9 9 10 9 9 15 3 13 2
50 9 9 1 9 9 16 9 7 9 15 14 4 1 0 9 9 9 13 2 13 2 2 0 1 9 9 2 9 9 13 2 9 9 7 9 7 2 7 9 16 9 9 7 9 1 9 0 9 13 2
17 9 9 9 0 16 9 9 9 13 16 1 9 9 0 0 13 2
34 16 10 9 9 0 1 9 13 7 9 0 1 9 15 13 2 3 0 0 13 9 13 16 9 1 9 9 9 7 9 9 9 13 2
66 9 1 9 16 1 10 9 1 9 9 7 9 9 13 13 9 9 9 0 1 9 9 9 0 7 9 0 7 1 0 9 9 13 13 7 1 9 9 9 15 9 9 9 9 0 7 12 9 0 7 3 9 0 9 13 16 9 0 1 9 14 9 7 0 13 2
31 9 16 1 3 1 9 13 13 15 16 2 9 9 1 3 9 1 15 9 13 16 10 9 1 12 9 7 9 9 13 2
33 9 9 1 9 15 12 9 0 9 7 9 14 9 12 9 13 16 1 9 0 1 9 7 9 2 9 7 9 0 14 1 13 2
94 9 3 1 9 1 9 10 12 9 16 12 9 9 14 9 15 13 7 9 14 3 0 9 0 13 7 9 0 16 9 14 1 9 7 9 9 0 13 13 13 2 9 16 15 14 0 9 13 2 9 0 1 9 13 7 1 9 2 0 9 13 7 0 13 16 1 9 9 13 9 16 1 10 9 13 7 15 14 1 9 9 1 9 9 13 2 0 1 10 9 0 9 13 2
16 1 9 0 9 0 1 9 15 15 14 16 0 9 0 13 2
27 1 10 9 2 0 1 9 9 1 1 9 7 9 2 12 9 0 1 12 9 9 9 7 9 0 13 2
73 1 9 0 2 12 9 9 7 9 1 9 7 9 15 9 1 9 9 15 13 7 1 9 1 10 9 1 9 9 0 9 9 9 13 7 3 16 4 9 15 14 1 15 9 13 2 9 13 16 1 12 9 2 1 9 1 9 15 7 9 9 9 0 1 9 15 2 9 15 14 9 13 2
12 1 10 9 2 9 9 0 0 9 0 13 2
32 9 3 9 13 1 9 16 1 15 13 2 1 9 0 9 13 7 9 15 14 1 9 7 9 7 9 9 9 9 3 13 2
24 3 9 0 7 9 0 15 1 1 9 9 9 0 13 13 2 3 1 10 9 0 9 13 2
64 9 7 9 9 0 16 9 13 3 1 9 0 9 0 9 2 9 0 1 15 13 9 13 16 1 12 9 0 9 13 7 9 9 7 9 15 1 9 7 9 14 1 9 9 13 7 1 9 0 2 9 15 14 1 9 0 0 1 9 7 9 0 13 2
24 9 0 10 9 2 0 9 9 0 1 9 9 9 2 7 0 9 10 9 2 1 9 13 2
50 2 9 2 1 9 0 9 2 9 9 9 13 16 1 15 13 2 0 1 9 16 12 9 0 14 1 9 1 1 9 0 9 1 9 13 3 3 13 9 9 15 14 1 9 9 7 9 9 13 2
48 9 7 9 10 9 0 0 1 9 7 9 0 1 9 9 1 9 9 0 13 2 3 9 0 0 7 0 9 10 9 7 9 13 16 3 9 15 1 9 0 1 9 7 9 0 4 13 2
33 9 16 9 9 2 9 1 1 9 9 7 9 10 9 13 7 13 1 9 9 7 9 15 9 0 9 0 7 3 0 9 13 2
33 16 9 3 13 7 13 16 1 9 7 9 10 9 0 13 2 7 9 9 9 3 9 7 9 9 1 9 9 14 0 13 13 2
63 1 10 9 9 0 1 0 9 15 1 9 0 9 9 10 9 7 9 14 1 9 9 9 13 16 1 0 9 9 12 3 9 1 9 7 9 16 1 9 0 2 9 7 9 9 13 0 1 15 13 16 9 9 1 9 0 9 3 7 3 9 13 2
39 9 9 1 10 12 9 0 1 9 2 9 7 9 0 7 0 13 16 1 9 9 7 9 0 9 7 9 15 1 9 9 1 9 9 9 9 13 13 2
43 12 1 9 0 7 9 0 1 9 9 15 13 16 15 14 1 9 7 9 9 7 9 0 9 13 7 3 1 9 7 9 0 7 0 0 9 0 14 1 9 9 13 2
37 9 0 13 16 9 12 9 7 9 0 1 9 10 9 13 7 15 9 9 0 13 16 9 9 1 9 15 13 7 9 15 1 9 0 15 15 2
32 9 7 9 0 15 1 9 9 0 10 9 14 1 9 13 16 3 12 9 1 9 0 15 1 9 9 0 7 0 9 13 2
123 9 0 10 9 14 4 1 1 9 9 9 13 16 9 9 14 3 1 9 7 9 9 0 2 0 7 0 15 13 7 0 13 1 9 0 7 0 15 1 9 9 9 0 7 0 1 9 9 0 13 2 3 16 9 0 0 9 1 0 9 0 15 16 9 9 0 9 13 2 3 0 1 10 9 1 9 7 9 9 7 9 15 1 9 9 9 9 9 9 13 13 2 16 15 16 9 14 9 12 9 7 9 13 7 16 9 16 9 3 9 9 7 9 9 14 1 9 0 1 9 0 13 2
54 1 9 9 10 9 3 9 0 9 13 16 0 13 9 1 9 0 1 9 9 1 9 9 15 0 13 2 15 16 3 9 0 7 1 9 9 9 0 2 7 9 16 1 9 9 9 15 14 1 9 9 13 13 2
45 0 13 16 10 9 1 9 7 9 9 9 7 9 13 16 3 1 9 0 7 0 7 1 9 9 9 13 7 9 0 3 1 9 7 9 15 9 7 9 0 14 9 13 13 2
39 9 9 9 0 9 0 9 1 9 1 9 13 7 13 13 16 1 0 9 0 3 12 9 9 7 9 1 9 1 9 7 9 9 13 7 13 13 13 2
49 9 0 9 1 9 15 9 7 9 16 1 15 9 13 1 3 0 9 9 7 9 14 1 9 9 13 13 7 10 9 7 9 9 3 1 9 9 7 1 9 1 9 7 9 9 15 13 13 2
28 16 1 9 13 16 9 9 9 0 9 1 9 9 2 9 7 9 0 1 9 7 9 9 9 1 9 13 2
21 3 16 9 9 0 1 9 0 9 1 9 13 13 2 9 0 9 0 0 13 2
24 9 9 1 9 12 9 9 9 9 13 13 2 9 0 12 12 9 9 9 0 14 9 13 2
50 10 9 13 13 2 1 9 9 15 2 9 9 9 9 0 1 9 9 9 1 9 10 9 13 2 9 0 0 1 9 7 9 2 9 7 9 7 9 13 2 7 10 9 9 9 9 9 0 13 2
45 15 16 9 0 1 9 9 1 9 9 0 9 9 13 2 9 13 2 3 1 12 9 0 1 9 2 12 9 1 9 0 13 16 12 9 1 9 1 12 9 0 1 9 13 2
65 10 9 0 1 9 1 15 16 12 9 0 0 7 0 1 9 0 13 2 13 2 9 16 1 9 9 9 0 13 0 1 9 0 1 9 9 13 1 9 0 2 9 9 16 9 13 3 9 13 9 14 1 9 1 9 15 13 7 1 9 9 16 9 13 2
14 15 9 13 2 9 0 9 1 9 0 9 13 2 2
5 9 3 4 13 2
58 9 9 1 9 2 9 9 0 3 4 13 2 2 13 2 9 9 1 9 7 9 0 1 9 13 16 9 9 0 1 9 0 2 9 9 7 9 0 14 1 9 9 13 7 9 9 7 9 1 9 9 7 9 0 14 0 13 2
32 9 1 9 7 9 9 1 9 7 9 9 0 9 2 9 13 7 9 9 0 7 9 7 9 0 9 9 14 1 9 13 2
84 3 1 9 0 9 16 1 9 9 15 9 13 2 9 7 9 0 7 3 0 15 14 1 10 9 0 1 9 0 1 9 7 9 9 13 7 1 9 9 9 9 7 9 0 10 9 9 0 9 9 1 9 13 16 9 9 7 9 9 0 1 9 1 10 9 10 9 1 9 13 16 9 9 9 7 9 0 14 1 9 9 0 13 2
70 0 9 10 9 2 9 7 9 9 0 7 7 0 9 2 3 9 9 0 13 16 1 9 9 1 9 7 9 7 9 1 9 9 0 9 13 7 1 9 9 9 0 2 9 1 9 7 9 0 7 7 2 9 9 0 0 7 0 9 9 9 9 0 7 9 9 15 9 13 2
82 1 9 2 9 0 0 16 1 9 15 16 9 0 9 14 1 9 9 1 9 7 9 13 2 1 9 9 7 9 9 2 3 1 9 1 10 9 13 16 3 1 9 1 9 9 9 13 7 15 7 1 9 0 7 0 2 0 2 0 7 0 1 9 9 13 16 9 9 9 1 9 7 9 1 9 9 14 1 9 0 13 2
52 9 0 9 0 1 9 0 7 3 1 9 0 2 9 7 9 9 0 14 9 13 7 3 9 9 7 9 1 9 9 0 7 9 14 1 9 0 7 9 7 9 9 0 14 1 9 9 7 9 9 13 2
34 16 2 4 9 0 2 9 9 7 9 14 9 13 7 1 0 9 9 1 15 2 9 14 1 9 10 9 7 9 9 0 0 13 2
73 1 10 9 9 13 9 2 9 7 9 0 2 9 9 0 15 14 3 1 9 9 7 0 13 7 9 0 1 9 0 14 16 9 13 2 12 9 0 0 9 14 1 9 9 1 9 7 7 9 1 9 13 7 16 2 9 7 9 0 14 0 9 13 2 1 9 9 7 9 0 15 13 2
65 7 1 10 9 2 3 9 0 9 1 9 0 9 2 1 9 9 0 9 9 13 7 9 15 1 9 14 1 9 7 9 9 13 7 1 9 1 9 9 7 9 1 9 9 0 2 9 9 9 0 7 9 0 1 9 9 9 14 1 9 0 10 9 13 2
27 4 10 9 14 1 9 0 13 7 0 13 16 15 9 0 1 9 9 15 7 9 1 9 15 9 13 2
51 9 7 9 14 0 13 7 1 9 9 0 2 9 14 9 13 7 9 0 14 1 9 9 7 9 15 13 7 10 9 1 9 15 7 1 9 9 15 2 1 9 9 9 9 7 9 9 9 9 13 2
9 9 16 9 9 15 14 13 13 2
39 9 0 1 9 9 1 9 9 0 15 1 9 9 13 7 1 9 1 9 9 13 2 1 9 12 1 9 15 9 1 9 0 13 7 1 15 9 13 2
21 9 15 1 15 7 1 15 9 13 13 12 9 1 9 15 14 1 9 15 13 2
86 15 12 9 9 0 13 1 15 7 1 9 9 12 9 15 0 9 0 13 7 15 1 15 7 1 15 9 13 13 1 9 9 15 1 12 1 9 9 9 9 13 7 9 15 14 16 0 1 12 12 9 9 13 1 10 9 1 9 13 7 9 0 9 9 12 12 9 1 9 9 9 1 15 13 16 1 10 9 1 9 9 9 15 0 13 2
37 15 9 13 2 12 9 3 1 10 9 16 1 9 10 9 1 9 0 9 13 16 3 9 13 16 9 1 3 9 1 9 9 0 9 13 13 2
14 10 9 9 13 2 1 9 9 15 9 15 0 13 2
35 9 1 9 9 15 9 13 7 16 15 16 0 13 9 13 9 15 13 7 1 9 0 9 14 9 13 7 9 9 14 15 15 9 13 2
65 1 10 9 1 9 9 16 1 9 9 13 13 13 7 1 9 9 2 9 7 9 15 9 12 12 9 14 9 13 7 3 13 9 9 14 0 13 16 9 13 16 9 9 14 1 9 0 13 13 1 9 0 9 13 7 1 9 9 0 9 9 9 15 13 2
28 7 9 9 1 9 0 1 15 13 16 9 0 9 15 1 9 1 9 7 9 9 2 9 14 9 13 13 2
24 15 1 9 10 9 0 13 7 1 9 9 9 9 15 1 15 13 16 9 15 9 13 13 2
31 7 9 9 1 9 9 9 7 9 0 7 9 9 3 1 15 13 15 1 10 9 7 9 0 9 14 1 15 9 13 2
43 1 9 10 9 9 9 2 9 10 9 0 14 1 9 9 7 9 0 7 9 1 9 12 9 16 1 9 9 13 1 9 1 9 9 13 7 1 15 9 1 9 13 2
41 7 15 1 15 1 9 9 9 1 9 9 13 16 1 3 9 7 3 1 9 9 1 9 0 13 2 7 9 9 9 9 14 1 9 7 9 1 9 9 13 2
38 9 9 1 9 9 9 7 0 1 9 9 9 13 2 16 9 10 9 1 9 9 12 12 9 9 9 0 7 9 9 2 9 0 14 9 13 13 2
46 9 3 1 9 9 7 9 0 9 9 13 16 9 1 9 9 12 16 12 9 3 1 9 9 1 9 16 15 14 9 10 9 9 13 9 13 7 1 9 9 16 9 9 13 13 2
41 1 9 10 9 2 9 1 9 10 9 0 0 7 9 9 16 9 14 1 9 13 3 9 15 14 9 13 13 7 1 9 9 9 9 14 1 9 1 9 13 2
6 9 2 9 0 9 2
29 9 9 0 9 9 9 9 13 2 1 1 9 9 0 1 12 9 0 2 3 12 9 13 7 12 9 0 13 2
29 1 9 9 9 1 9 2 9 10 9 13 2 1 9 9 9 9 1 9 9 12 9 13 7 12 9 0 13 2
31 10 9 13 2 1 9 9 9 0 1 9 9 16 1 9 9 7 9 9 0 13 2 12 9 1 9 12 9 13 13 2
8 9 9 1 9 1 9 13 2
6 9 2 9 0 9 2
26 3 1 9 1 9 9 9 1 9 2 3 12 1 9 9 9 9 9 9 10 9 7 9 9 13 2
66 1 9 9 0 9 1 9 1 9 0 9 2 1 9 9 0 16 1 12 9 9 7 9 9 9 9 7 9 9 1 9 1 9 9 1 9 9 9 13 2 12 9 13 13 7 9 0 1 9 0 13 16 12 1 15 1 9 9 9 1 9 9 0 13 13 2
48 1 1 10 9 2 9 0 9 3 1 1 9 10 9 9 13 7 9 0 16 10 9 1 9 9 1 9 13 2 1 1 9 9 9 0 1 9 13 16 9 9 7 9 15 14 9 13 2
41 9 7 9 0 1 9 15 13 13 2 7 9 9 0 14 16 2 16 1 10 9 1 1 9 9 9 13 13 2 1 9 0 7 1 9 12 9 0 9 13 2
27 1 10 9 9 1 9 9 0 9 0 7 0 14 1 1 9 9 9 0 7 0 1 15 1 9 13 2
19 1 10 9 0 2 1 3 9 1 9 9 13 16 3 9 0 9 13 2
51 9 16 9 9 3 1 15 14 3 0 13 1 9 9 16 1 10 9 13 13 9 13 7 1 3 16 3 9 15 1 9 9 15 9 13 7 1 9 9 0 0 16 9 1 10 9 1 15 9 13 2
75 16 9 9 0 15 9 9 14 2 16 3 13 13 2 1 13 2 4 13 16 9 9 16 9 9 15 14 13 7 9 15 14 0 13 12 9 3 1 9 15 2 3 1 9 16 15 1 15 13 13 7 13 13 2 1 9 9 0 7 0 2 1 9 9 7 9 0 0 16 9 9 13 9 13 2
42 16 9 9 0 9 1 9 3 3 9 13 13 2 9 0 9 13 13 16 9 2 0 1 15 16 9 9 7 9 0 0 15 13 2 9 9 10 9 0 0 13 2
65 1 9 9 7 9 0 16 1 9 0 9 9 9 1 9 12 1 9 0 13 2 9 9 9 9 9 7 9 9 9 1 9 0 15 1 9 9 1 9 7 9 9 13 16 9 0 9 1 12 9 1 9 16 9 1 9 9 15 13 13 2 0 13 13 2
35 3 9 3 1 9 9 1 9 0 7 9 0 2 16 3 9 13 13 2 9 0 1 9 13 16 9 9 1 9 7 9 14 0 13 2
31 13 16 1 10 9 9 0 7 9 9 9 13 7 9 4 1 9 7 9 15 9 7 9 9 1 9 15 14 9 13 2
62 13 16 9 0 9 0 0 2 9 2 16 1 9 9 2 15 16 3 9 3 1 9 9 9 13 7 9 9 7 9 15 1 9 9 7 9 16 13 13 7 0 13 2 1 9 10 9 1 9 9 0 15 9 0 9 9 9 9 14 9 13 2
52 16 9 9 16 9 9 9 12 9 14 16 1 9 10 9 0 13 13 1 9 13 2 16 9 9 1 9 9 3 1 9 1 10 9 16 1 15 9 13 2 7 9 9 1 9 0 7 0 9 9 13 2
66 16 1 9 0 2 9 0 9 9 16 9 16 9 0 15 1 9 7 9 13 2 1 9 13 0 13 16 15 2 9 12 9 3 1 9 1 9 9 9 1 9 10 9 9 0 13 13 13 7 12 9 0 12 7 0 1 9 9 15 14 1 9 9 13 13 2
29 9 0 9 13 13 16 9 9 2 1 9 15 1 9 9 15 1 9 9 0 1 9 0 9 9 13 13 13 2
35 16 1 10 9 9 13 13 13 16 9 9 0 0 1 9 0 9 13 7 9 9 15 14 12 1 9 0 1 9 9 1 9 9 13 2
47 9 0 9 2 8 8 8 8 8 9 9 2 16 1 9 9 9 0 13 13 2 16 9 9 1 10 9 1 9 9 9 9 9 0 1 9 13 16 3 1 9 1 9 9 0 13 2
21 16 9 1 10 9 9 13 15 1 9 9 0 7 9 0 9 9 14 9 13 2
72 9 1 10 9 16 1 9 9 9 3 9 13 9 0 15 13 16 9 1 15 13 16 9 9 0 9 14 16 1 9 9 9 0 13 9 13 12 2 10 9 3 2 1 9 9 9 9 9 1 10 9 16 9 9 9 13 2 1 9 0 7 1 9 0 1 9 9 0 0 3 13 2
18 9 9 1 10 9 1 9 1 9 2 9 1 9 9 0 9 13 2
18 9 9 0 9 0 13 2 7 9 9 9 0 3 0 9 0 13 2
17 9 0 9 12 9 3 1 9 1 9 0 1 9 9 9 13 2
44 1 9 0 9 0 7 1 9 0 0 9 16 3 9 16 13 9 14 9 13 16 1 15 13 0 9 1 9 12 9 9 13 13 7 7 3 9 0 1 15 9 13 13 2
59 9 1 9 9 9 1 9 9 0 9 0 3 1 9 9 13 7 1 9 16 9 13 13 2 7 9 0 9 10 9 14 1 9 0 9 7 9 13 7 1 9 9 7 9 9 14 1 9 0 7 0 15 1 9 3 0 13 13 2
75 9 16 16 1 9 7 16 1 9 2 9 9 9 7 9 7 9 0 13 12 2 9 1 9 1 9 9 16 13 13 13 7 13 16 15 7 9 7 9 9 9 9 1 9 9 9 1 9 9 13 16 9 0 14 9 13 7 9 9 15 9 13 16 9 9 9 13 7 1 9 0 9 9 13 2
10 9 9 12 9 1 9 1 9 13 2
9 9 9 14 16 1 10 9 13 2
58 9 9 1 9 9 7 3 9 9 10 9 2 0 1 9 0 15 1 9 9 9 7 9 0 10 9 2 1 10 9 16 0 9 13 16 1 9 9 9 9 9 1 9 9 9 2 9 0 1 9 9 9 1 9 9 13 13 2
12 3 1 9 1 9 9 16 9 9 13 13 2
24 9 16 1 9 9 1 9 9 13 3 1 9 9 13 16 1 9 0 1 10 9 13 13 2
44 1 9 16 9 9 1 9 9 0 13 10 9 1 9 16 9 13 2 7 16 0 13 16 9 1 9 16 13 13 7 3 1 10 9 1 9 9 1 9 0 9 13 13 2
33 1 10 9 2 16 1 9 0 9 9 1 9 15 13 2 9 1 9 15 1 9 1 9 0 7 1 9 9 0 16 0 13 2
41 9 0 15 13 16 15 9 0 13 13 2 7 15 16 7 9 15 1 9 1 9 15 1 9 7 9 0 9 13 7 3 9 13 16 3 1 15 9 4 13 2
51 9 0 1 9 16 3 0 13 13 9 15 1 9 9 0 13 16 1 9 15 12 1 9 0 9 2 9 2 9 7 9 9 9 1 9 13 7 3 0 13 16 9 3 9 1 10 9 16 13 13 2
17 9 9 1 9 15 1 9 8 8 8 9 9 9 9 13 13 2
19 15 9 13 16 9 10 9 14 1 9 7 9 9 9 9 9 13 13 2
10 3 7 9 9 14 1 9 13 13 2
17 9 0 1 9 9 9 9 15 1 9 9 9 2 9 2 13 2
37 1 10 9 3 9 0 1 9 9 13 2 7 9 15 1 9 9 9 0 1 9 1 1 9 9 16 9 9 9 9 9 13 2 9 13 13 2
17 9 0 10 12 9 2 1 9 15 9 0 15 2 9 13 13 2
36 9 9 3 1 15 0 9 1 9 0 9 13 13 16 12 1 15 9 13 16 15 9 9 9 2 1 9 9 9 9 2 1 9 13 13 2
28 7 9 9 0 1 15 13 16 15 9 16 1 3 1 9 9 13 13 1 9 9 15 1 9 9 13 13 2
41 1 9 9 1 3 9 0 0 9 13 7 0 9 0 15 9 13 16 9 9 9 9 1 9 12 9 1 10 9 9 13 13 7 1 9 9 15 0 13 13 2
14 16 9 0 1 9 9 0 0 9 9 9 9 13 2
16 12 2 9 1 9 9 1 8 9 1 10 9 9 13 13 2
63 1 9 9 9 9 9 2 9 0 9 9 0 2 9 9 1 8 9 1 3 9 9 9 0 9 2 9 9 13 16 1 9 15 9 0 1 9 9 13 1 9 0 16 2 1 3 16 1 9 9 7 0 15 13 2 1 9 0 0 0 13 13 2
50 9 1 8 9 9 13 16 3 1 9 9 9 9 0 9 3 10 9 14 9 13 13 2 7 3 1 10 9 1 9 0 13 7 9 0 14 1 9 9 16 1 9 12 9 0 13 9 13 13 2
31 12 2 9 1 12 9 1 9 9 2 1 9 12 9 13 13 16 1 12 9 12 9 0 1 12 9 0 4 9 13 2
25 9 9 13 9 13 16 10 9 12 9 16 9 15 0 13 13 7 1 9 9 0 0 9 13 2
24 1 15 9 7 8 9 1 10 9 9 0 13 13 7 3 1 15 16 9 9 9 3 13 2
19 7 1 3 9 9 9 0 1 9 9 9 9 1 9 0 9 13 13 2
25 0 9 9 1 9 0 1 9 0 9 0 9 9 9 7 1 9 9 0 1 9 9 9 13 2
43 1 10 9 9 9 9 7 7 9 0 9 9 9 2 9 2 9 2 9 7 9 0 0 9 12 7 12 9 9 2 7 9 15 1 9 9 9 7 9 9 4 13 2
49 1 9 9 0 9 9 0 9 2 1 9 9 9 9 9 0 9 0 1 9 0 0 0 16 1 9 9 1 9 9 0 3 1 9 7 9 0 3 12 9 0 0 9 13 1 9 13 13 2
28 10 9 16 1 9 7 9 1 9 0 7 1 9 0 9 13 0 9 12 2 12 1 12 2 12 9 13 2
29 1 12 9 15 9 9 13 16 9 9 12 9 7 9 12 9 9 0 2 9 2 9 2 9 7 9 2 13 2
39 9 0 0 1 9 9 0 0 1 9 12 7 12 9 9 2 9 9 0 9 9 1 9 9 0 7 9 0 0 1 9 9 1 0 9 10 9 13 2
37 0 13 9 1 9 9 9 2 1 9 9 9 2 1 9 9 2 9 9 2 1 9 16 9 9 7 9 0 9 13 16 1 10 9 9 13 2
36 16 9 0 9 0 9 9 7 9 1 9 0 7 9 1 0 9 13 16 1 9 9 0 7 1 12 9 1 12 9 1 10 9 0 13 2
4 9 2 9 2
25 9 9 0 1 9 9 16 1 9 9 13 2 1 9 9 9 1 9 9 1 9 15 9 13 2
68 9 9 9 10 9 9 9 1 12 9 0 1 12 9 0 9 1 9 9 9 1 9 9 9 2 9 0 9 9 2 1 9 15 9 13 7 13 2 9 13 9 7 9 15 1 10 9 9 14 9 13 13 16 1 9 9 0 13 13 16 10 9 9 9 0 15 13 2
35 15 16 1 1 9 9 9 9 1 9 1 9 0 9 9 13 13 2 1 9 3 9 13 7 1 1 16 9 9 1 15 9 9 13 2
50 9 9 9 3 1 9 0 1 9 0 1 9 0 9 2 9 9 1 9 9 14 3 9 13 7 13 2 9 15 15 13 16 9 0 1 9 9 13 2 9 1 9 9 1 9 9 9 13 13 2
18 15 13 2 10 9 9 13 9 1 9 13 16 9 15 14 0 13 2
15 9 9 13 2 3 0 13 15 1 9 9 9 9 13 2
29 3 1 9 9 2 1 9 15 7 9 9 9 2 3 9 9 9 0 9 13 16 12 9 1 9 13 13 13 2
51 12 9 3 9 9 9 9 1 9 9 9 1 9 9 9 13 7 9 1 15 3 9 13 7 12 9 3 1 15 9 1 9 1 9 9 2 9 9 2 1 15 9 13 7 1 9 12 0 9 13 2
39 9 16 9 1 9 0 9 9 9 7 9 9 12 10 9 3 1 9 9 9 9 9 13 2 3 1 9 10 9 9 0 13 7 1 10 9 9 13 2
45 9 1 9 7 9 9 3 3 13 16 9 15 3 1 9 9 9 9 13 13 7 15 0 13 15 13 16 12 9 16 1 9 9 0 9 9 9 13 1 9 9 1 9 13 2
25 9 9 16 1 9 9 1 9 9 9 13 13 2 1 9 9 9 9 9 9 14 1 9 13 2
23 9 9 7 9 0 9 9 0 9 9 2 12 2 12 2 7 1 9 0 9 0 13 2
19 9 9 3 12 9 9 9 9 13 7 1 12 1 0 9 9 9 13 2
41 9 15 1 12 9 0 9 7 3 16 0 13 9 0 7 9 0 13 2 16 1 9 9 9 0 16 0 13 7 3 9 9 15 1 9 1 10 9 13 13 2
24 9 9 9 0 9 0 0 9 7 9 9 9 13 7 9 0 15 3 1 9 9 13 13 2
34 15 1 9 9 7 16 9 13 7 9 0 7 0 16 1 9 9 1 9 9 15 13 2 1 0 9 0 9 9 1 9 13 13 2
49 9 3 1 9 9 0 1 9 15 13 2 10 9 14 1 9 0 7 0 7 0 16 9 15 1 15 9 0 13 13 2 7 3 3 13 16 3 9 9 9 13 16 4 15 14 1 9 13 2
13 9 13 16 1 1 9 9 1 9 9 0 13 2
21 6 9 15 16 4 9 15 14 16 1 15 9 13 7 1 9 10 9 9 13 2
28 1 3 9 0 1 9 1 9 9 13 2 9 13 7 9 0 13 7 9 9 9 9 14 1 9 9 13 2
47 3 0 13 9 7 9 14 16 1 10 9 2 1 9 0 15 13 16 3 7 3 2 3 3 7 3 3 1 9 9 0 1 0 7 9 13 16 1 1 9 0 1 9 9 9 13 2
20 3 7 3 10 9 0 7 0 16 9 0 14 1 9 0 0 13 9 13 2
30 3 9 1 9 9 16 9 9 9 13 1 9 13 2 7 3 10 9 14 13 16 9 0 9 14 1 9 0 13 2
21 6 9 9 9 2 15 3 0 9 9 15 13 2 7 3 3 1 9 9 13 2
42 16 7 1 15 9 0 13 7 3 1 9 15 13 2 10 9 1 9 1 15 13 2 15 13 7 9 0 1 9 9 15 7 1 9 15 14 1 15 1 9 13 2
20 7 3 0 13 1 10 9 9 0 7 0 9 9 1 9 0 15 0 13 2
13 3 0 13 1 10 9 9 9 9 3 13 13 2
18 3 13 16 13 1 0 9 9 16 3 3 7 0 13 2 9 13 2
30 3 13 16 13 1 10 9 9 2 1 9 9 0 2 9 13 16 3 1 15 13 2 9 13 16 3 9 9 13 2
25 3 13 16 13 3 10 9 13 16 1 9 0 1 9 0 2 0 9 1 9 9 0 13 13 2
6 9 2 9 0 9 2
27 1 9 9 1 9 0 9 9 9 9 1 9 7 9 0 1 9 9 7 9 9 9 7 0 13 13 2
30 10 9 1 9 9 9 12 12 9 9 9 12 12 9 9 13 13 7 9 1 15 9 9 9 9 9 1 9 13 2
32 10 9 0 16 1 12 9 9 0 7 0 9 13 13 12 9 9 7 9 12 9 9 13 7 0 9 9 9 9 13 13 2
28 9 10 9 0 0 16 1 9 9 0 0 7 0 13 13 13 2 9 1 10 9 0 0 9 0 9 13 2
42 9 1 10 9 15 13 16 1 9 9 13 2 1 9 1 9 9 9 16 10 9 9 1 15 1 9 1 9 15 9 13 2 3 9 0 9 16 1 1 4 13 2
15 10 9 0 0 9 0 1 1 9 9 1 9 9 13 2
18 12 9 9 1 10 9 1 10 9 0 7 0 0 9 13 4 13 2
19 0 9 1 9 1 9 0 16 1 9 12 12 9 9 13 9 4 13 2
6 9 2 9 0 9 2
21 9 1 9 7 9 0 1 9 9 9 16 9 9 0 7 9 13 2 9 13 2
19 9 7 9 9 13 16 9 0 1 9 9 9 1 9 1 9 0 13 2
13 9 9 9 9 0 1 9 0 1 9 9 13 2
15 3 1 9 9 2 9 9 14 0 1 9 0 0 13 2
53 9 0 1 9 9 7 9 0 16 9 0 1 9 0 1 15 0 13 2 1 9 9 9 9 13 7 9 9 1 10 9 9 0 13 2 10 9 16 1 9 9 9 2 9 0 7 3 9 0 1 9 13 2
40 9 9 9 9 14 1 10 9 7 1 9 1 9 2 9 2 9 2 9 2 9 2 9 2 9 0 2 9 2 9 7 7 9 9 7 1 9 9 13 2
14 1 9 9 0 1 10 9 9 7 9 0 9 13 2
38 9 1 13 9 0 9 1 12 9 0 1 15 9 0 9 13 7 9 0 1 9 9 0 7 9 0 13 7 9 0 1 9 9 0 16 0 13 2
19 1 9 0 2 15 1 9 0 9 9 9 1 9 9 1 9 0 13 2
56 9 9 9 9 9 7 9 0 1 9 9 9 13 2 9 9 9 14 12 9 3 7 1 9 9 9 9 1 9 0 13 16 3 1 15 10 9 1 9 16 12 12 9 3 1 9 9 1 9 13 13 2 9 13 13 2
6 9 2 9 0 9 2
16 9 13 16 9 9 0 1 9 9 9 1 9 0 9 13 2
39 9 9 2 9 9 1 9 9 2 1 9 9 1 9 1 9 9 9 16 1 1 9 9 13 7 13 2 9 9 0 1 9 9 9 1 9 0 13 2
36 9 1 9 9 9 9 7 0 9 9 9 0 1 9 7 9 9 9 9 16 9 1 9 13 2 9 0 1 9 9 1 1 9 9 13 2
44 9 9 13 2 3 10 9 1 9 0 0 13 7 1 9 16 3 9 9 0 1 9 9 0 2 9 2 9 9 1 9 7 9 1 15 9 13 2 9 9 9 0 13 2
37 9 1 9 9 9 13 16 9 14 1 9 0 9 9 0 9 13 7 1 10 9 16 9 9 1 9 15 13 2 9 0 1 9 14 9 13 2
7 9 1 9 9 9 13 2
4 9 2 9 2
39 12 9 0 9 9 13 2 16 9 9 9 9 16 1 9 9 7 9 0 0 13 2 3 1 9 0 9 13 2 7 9 13 9 0 15 9 13 13 2
41 9 9 9 1 10 9 13 2 9 1 9 15 1 9 0 7 0 2 9 13 16 9 15 1 9 9 9 1 9 9 9 1 9 2 3 1 9 9 13 13 2
35 9 9 9 9 1 9 2 9 9 1 9 9 13 2 1 3 16 0 1 9 9 13 2 9 0 13 7 15 16 9 13 2 9 13 2
27 15 13 16 9 3 9 4 13 7 4 10 9 3 1 9 10 9 13 2 3 7 9 9 0 4 13 2
20 12 9 1 9 9 9 9 9 1 9 9 12 9 0 10 9 14 9 13 2
16 10 9 3 1 12 9 0 13 9 9 9 9 0 9 13 2
22 10 9 1 9 0 1 9 12 1 12 1 9 9 9 0 13 7 1 9 0 13 2
32 9 10 9 9 1 9 9 9 9 14 1 9 15 0 13 7 1 9 0 1 9 9 7 9 13 7 10 9 14 9 13 2
4 9 2 9 2
28 12 9 9 0 9 9 9 9 9 9 13 2 1 12 1 9 9 9 0 1 9 12 9 0 9 13 13 2
30 9 9 9 9 9 1 13 7 13 1 9 13 2 3 9 9 9 1 12 0 10 9 1 10 9 9 9 13 13 2
31 10 0 7 9 13 2 3 9 0 16 13 9 1 9 10 9 1 9 9 1 12 2 12 1 12 2 12 9 9 13 2
35 1 9 10 9 9 0 2 10 9 1 9 1 9 12 9 1 9 9 12 12 7 12 9 9 1 9 1 9 12 2 12 9 9 13 2
31 9 9 13 2 12 9 9 1 9 9 9 13 16 15 0 9 0 1 9 9 1 10 9 13 16 1 9 9 9 13 2
29 9 9 0 12 9 0 9 2 9 2 9 7 9 13 16 12 9 3 1 9 9 1 0 9 1 9 13 13 2
17 9 0 9 13 9 0 9 14 1 1 9 9 7 9 9 13 2
29 1 9 10 9 2 9 0 0 12 9 0 1 9 9 13 16 9 9 1 9 0 9 13 7 15 14 0 13 2
14 10 9 9 9 9 9 1 1 9 7 9 9 13 2
49 9 9 1 9 0 9 0 9 13 9 16 9 15 0 1 9 0 13 2 0 1 9 7 9 0 0 13 7 9 16 1 9 9 0 9 1 9 7 9 9 13 2 0 1 10 9 0 13 2
23 9 10 9 0 13 9 14 1 9 9 9 13 16 1 9 0 1 9 7 9 13 13 2
33 10 9 13 1 9 3 0 16 9 1 9 13 2 9 0 9 14 9 7 0 13 7 9 14 1 1 9 7 9 0 9 13 2
6 9 0 9 2 9 2
25 9 13 2 4 1 9 0 9 1 9 9 1 9 9 9 0 3 1 9 9 0 0 9 13 2
31 9 9 1 9 9 7 9 15 1 9 12 9 9 0 2 1 9 9 9 9 10 9 0 1 9 9 9 0 0 13 2
25 9 9 0 1 15 13 16 9 9 9 1 9 9 16 9 0 0 13 2 1 9 0 9 13 2
27 1 1 9 16 9 9 1 9 15 0 1 12 2 12 9 1 9 13 12 9 0 0 9 0 0 13 2
22 9 9 13 2 9 9 16 9 9 0 9 13 16 9 9 9 0 0 14 9 13 2
11 10 9 13 9 9 0 1 9 0 13 2
20 9 0 1 9 9 1 9 16 1 9 9 9 13 13 1 9 0 9 13 2
24 10 9 9 1 9 9 7 9 0 14 1 9 9 13 7 15 14 1 9 0 9 9 13 2
10 10 9 9 9 0 9 0 9 13 2
17 12 9 0 1 10 9 1 9 9 9 12 0 12 0 9 13 2
22 1 9 0 3 9 0 9 1 1 13 7 9 9 7 9 0 0 9 16 9 13 2
25 10 12 9 3 1 9 9 9 9 1 9 9 10 0 2 9 0 9 14 16 1 15 9 13 2
21 15 3 1 12 9 9 13 16 9 9 9 13 7 9 16 1 9 9 9 13 2
17 1 9 9 0 9 3 1 9 9 0 9 1 9 0 9 13 2
22 10 9 16 1 9 9 0 0 13 2 7 3 0 13 7 9 7 9 1 9 13 2
24 1 9 1 10 9 9 16 9 13 0 9 4 13 7 4 9 0 9 14 1 15 9 13 2
14 9 0 9 9 9 1 9 9 0 14 9 13 13 2
27 9 9 9 1 9 1 13 1 9 16 0 9 9 7 9 13 2 9 9 0 1 9 0 1 15 13 2
22 1 10 9 2 9 1 9 12 9 7 12 9 9 13 16 9 9 15 14 9 13 2
24 1 9 0 1 9 2 9 9 1 9 9 13 7 9 9 9 1 9 15 1 9 9 13 2
22 9 15 13 16 9 16 1 9 9 9 0 13 2 9 9 0 1 9 15 0 13 2
27 9 9 13 16 1 1 9 9 0 3 9 0 1 9 12 9 0 9 7 9 15 1 9 9 0 13 2
19 9 0 9 13 13 16 0 9 10 9 1 9 9 9 0 14 9 13 2
23 16 4 9 13 16 12 9 0 9 9 0 1 9 0 3 9 9 9 1 9 15 13 2
47 9 13 9 9 1 9 9 9 13 2 16 1 9 9 9 9 9 1 9 9 7 9 7 9 13 2 9 9 0 9 13 2 9 9 0 13 7 9 9 0 16 1 9 9 4 13 2
71 9 2 9 9 9 16 9 0 15 14 3 1 9 9 0 0 7 9 9 9 7 9 7 9 9 7 9 9 9 7 9 9 9 7 16 9 9 9 13 2 3 1 1 9 9 9 0 7 9 0 1 9 0 7 0 1 9 0 13 7 1 9 9 9 7 9 7 9 9 13 2
80 9 16 1 10 9 2 9 0 9 1 9 9 0 7 9 9 9 9 9 0 9 0 9 2 9 0 1 9 9 9 13 7 1 9 9 0 7 9 9 9 10 9 1 9 13 1 9 9 15 9 7 9 9 0 1 9 9 0 13 16 1 9 9 7 9 0 9 9 9 9 7 15 1 9 7 9 0 9 13 2
65 1 9 9 0 15 1 15 7 0 1 12 9 1 9 0 9 13 2 3 9 13 1 12 1 10 9 2 9 0 0 7 9 0 9 9 9 9 1 9 9 7 9 9 16 1 12 9 13 9 0 9 7 9 9 14 1 10 9 0 9 13 2 9 13 2
28 16 3 7 9 0 13 2 9 0 9 9 9 1 9 12 9 0 7 0 0 1 9 9 0 7 0 13 2
117 1 9 9 10 9 0 1 10 9 16 9 1 9 0 1 9 9 9 9 9 16 1 9 7 9 0 9 7 9 7 0 1 9 9 9 7 9 9 1 9 1 9 13 2 9 13 1 9 9 10 9 7 3 1 9 0 1 15 1 9 1 9 9 9 3 9 7 9 13 16 9 9 9 9 9 7 9 9 0 15 14 16 3 0 1 9 0 7 0 9 9 13 1 9 13 16 1 10 9 9 10 9 7 9 9 9 9 1 9 12 1 9 0 9 9 13 2
153 9 9 9 9 16 15 1 9 0 1 9 7 9 9 9 9 1 9 9 7 9 7 9 7 9 9 0 13 2 16 1 10 9 13 16 10 9 14 1 9 13 2 7 9 0 7 9 0 15 9 1 9 10 9 13 2 1 3 1 9 9 7 9 0 9 2 9 9 9 1 9 9 9 1 10 9 0 2 9 1 9 0 2 1 9 9 7 9 0 9 9 9 2 9 0 7 9 9 9 9 9 9 9 0 9 9 7 9 0 9 9 9 9 16 1 10 0 9 9 15 1 9 9 9 9 0 13 2 9 1 9 14 1 9 0 1 9 9 13 7 1 9 9 0 16 9 0 15 14 13 9 13 2
39 3 1 9 1 9 0 7 9 0 1 9 9 9 1 1 9 0 9 9 9 9 9 9 0 1 9 1 9 12 9 9 0 1 9 9 9 9 13 2
57 9 9 9 2 9 0 0 13 16 9 0 9 15 14 1 9 9 9 13 7 1 9 4 13 15 1 9 0 7 0 1 9 9 9 9 1 9 2 3 9 0 14 9 13 7 1 9 15 9 9 14 1 9 9 15 13 2
28 9 10 9 3 1 9 9 15 9 13 7 15 14 0 9 15 13 7 10 9 3 9 1 9 9 15 13 2
35 9 1 9 9 9 9 13 13 7 1 9 9 15 3 9 9 9 12 9 16 9 9 9 2 9 9 7 9 14 1 9 9 13 13 2
30 13 16 1 9 12 9 0 2 0 7 0 9 13 13 7 6 2 1 10 9 10 9 3 0 1 12 9 0 13 2
42 9 9 9 0 13 7 1 10 9 9 15 1 10 9 0 13 7 1 10 9 9 9 13 13 16 3 1 9 0 13 2 16 9 9 7 9 9 3 9 13 13 2
38 7 1 9 1 9 9 9 9 13 13 16 15 1 9 9 9 9 0 13 2 16 0 13 16 1 9 9 0 2 9 9 9 1 9 15 9 13 2
19 9 9 2 9 9 7 9 13 16 1 9 9 1 9 1 9 9 13 2
44 0 13 1 10 9 3 1 9 7 9 2 12 9 9 7 9 0 0 9 13 7 1 9 0 7 0 7 0 9 0 13 7 9 1 9 9 0 1 9 0 9 13 13 2
14 10 9 3 0 13 16 4 1 15 0 9 9 13 2
25 1 10 9 3 13 13 16 1 9 10 9 2 9 0 7 0 9 1 3 9 1 9 9 13 2
41 1 10 9 1 9 0 13 16 12 9 7 9 1 9 1 9 13 7 12 9 0 7 0 1 9 13 16 9 15 1 9 9 9 0 2 1 10 9 0 13 2
55 3 9 9 9 1 10 9 2 9 0 9 9 9 1 9 9 9 13 7 9 9 9 10 9 14 9 13 16 9 1 9 2 9 7 9 0 1 9 0 9 10 9 13 7 9 0 9 13 16 1 9 9 4 13 2
54 9 9 0 12 9 1 12 9 2 9 12 9 1 12 9 2 9 12 9 2 9 0 12 9 2 9 9 12 9 2 9 9 0 12 9 2 9 9 7 9 12 9 2 9 9 12 9 2 7 9 12 9 13 2
20 9 1 9 9 1 9 1 9 9 9 7 9 9 9 9 7 9 0 13 2
25 1 9 9 9 1 9 13 16 15 3 1 15 1 9 9 0 9 13 16 0 1 15 0 13 2
15 1 9 9 2 9 12 9 7 3 9 12 9 0 13 2
29 3 1 9 10 9 9 13 2 12 2 1 9 0 9 13 13 7 1 9 9 9 15 1 15 0 10 9 13 2
26 1 9 12 9 0 9 13 12 9 9 9 9 9 9 0 7 0 13 2 0 1 9 12 9 13 2
22 0 13 9 3 9 9 7 9 14 1 15 0 13 13 16 1 9 0 1 9 13 2
9 1 10 9 9 9 3 0 13 2
46 7 9 9 1 10 9 9 13 13 7 0 1 9 13 16 9 16 1 9 10 9 9 13 7 1 9 15 2 9 15 14 9 13 13 7 9 15 14 3 9 9 3 0 9 13 2
50 9 0 16 1 10 12 9 0 13 15 13 16 9 9 9 9 13 16 1 9 1 9 9 13 2 1 9 7 9 9 9 9 13 16 1 9 2 9 0 2 9 7 1 9 0 1 9 0 13 2
24 12 1 9 9 9 15 13 16 1 9 9 9 2 9 7 9 0 14 1 15 9 13 13 2
17 7 1 9 9 9 9 1 1 9 7 9 9 2 12 9 13 2
133 15 1 9 9 13 13 16 1 9 0 0 13 7 1 9 0 0 3 9 9 2 9 0 13 13 2 9 9 1 9 9 13 2 9 9 15 1 10 9 15 16 9 9 9 14 3 7 3 13 7 9 9 16 1 9 9 9 9 9 14 3 13 2 1 10 9 9 9 9 9 9 9 0 1 9 9 1 9 13 2 1 10 9 15 9 9 0 15 13 16 1 9 1 9 13 7 9 9 9 16 0 13 2 16 1 9 13 16 9 9 9 0 13 2 9 15 14 1 9 0 16 9 9 13 4 13 16 1 9 9 9 13 2
42 12 2 1 9 1 9 9 13 13 2 9 10 9 9 7 9 13 7 9 15 9 2 16 1 9 9 0 2 0 9 13 7 9 0 14 1 9 9 16 0 13 2
18 1 10 9 1 9 9 2 1 1 15 16 15 9 13 9 0 13 2
36 3 13 16 9 10 9 13 2 16 0 13 16 15 3 9 0 13 2 7 3 1 9 9 9 13 2 16 9 3 1 9 0 1 9 13 2
13 9 9 1 9 9 9 13 7 1 15 13 13 2
16 9 9 9 12 9 13 1 9 7 9 9 9 12 9 13 2
17 1 9 9 3 9 1 9 13 2 7 1 9 9 9 0 13 2
9 1 10 9 9 9 0 9 13 2
27 1 9 9 9 9 1 9 13 2 1 9 7 1 9 3 1 9 2 9 1 9 9 9 9 13 13 2
11 1 10 9 16 9 1 9 9 9 13 2
15 7 1 9 0 2 9 9 1 9 0 9 13 8 8 2
20 12 2 3 7 3 9 13 1 9 3 1 9 10 9 1 9 9 13 13 2
18 16 3 9 9 0 15 13 7 10 9 1 9 9 0 9 0 13 2
32 12 2 1 9 1 9 12 9 0 2 9 0 1 10 9 0 13 2 16 3 1 9 0 4 1 15 12 9 0 9 13 2
94 12 2 16 1 10 9 0 9 16 1 3 9 13 3 9 13 13 2 7 1 9 1 15 16 12 9 1 9 9 0 7 0 16 9 9 9 9 7 9 9 9 0 9 0 13 2 9 9 1 9 0 10 9 9 0 13 7 1 9 9 4 13 3 9 0 3 1 9 9 3 9 14 1 9 15 1 9 13 7 1 9 0 3 9 13 13 1 10 12 9 0 9 13 2
43 9 10 9 1 9 9 15 1 9 2 0 9 0 1 9 1 9 3 1 9 9 14 1 9 13 7 1 1 15 0 9 13 13 7 13 1 9 0 10 9 9 13 2
22 7 1 9 9 9 0 1 9 13 7 9 9 0 1 9 15 9 9 9 13 13 2
50 13 3 9 1 9 0 1 9 15 9 1 9 2 9 2 9 7 9 9 2 9 0 7 0 1 15 3 0 13 7 1 9 9 9 9 9 9 9 0 9 9 1 9 1 9 0 9 9 13 2
14 1 15 7 9 14 0 3 12 9 1 9 13 13 2
37 0 13 3 9 0 1 3 13 13 3 9 9 1 9 15 9 9 1 3 9 9 13 7 0 13 16 9 12 9 0 16 1 15 9 13 13 2
27 1 9 1 9 0 3 9 7 9 0 7 0 13 13 1 12 9 0 16 9 9 9 7 9 9 13 2
17 16 10 12 9 1 3 1 9 13 7 9 0 15 16 0 13 2
16 7 3 16 4 1 9 9 7 9 3 1 9 9 9 13 2
25 9 9 9 1 9 9 9 16 1 9 0 9 13 13 7 15 16 1 10 12 9 0 9 13 2
17 16 9 0 16 1 9 7 9 9 1 9 9 9 3 9 13 2
12 1 10 9 16 10 9 9 9 9 15 13 2
54 9 9 9 13 16 1 9 10 9 9 0 9 13 16 9 7 9 1 3 9 9 13 7 9 9 1 9 1 9 12 9 0 0 4 13 2 3 7 1 1 10 9 0 1 10 9 2 4 12 9 0 9 13 2
48 3 1 9 9 9 9 1 9 0 7 0 13 7 0 9 7 9 13 16 9 0 3 1 9 0 10 9 0 14 9 13 7 10 9 0 9 9 9 1 9 9 9 0 9 1 9 13 2
15 1 3 10 9 0 9 9 9 7 9 1 9 9 13 2
15 1 9 9 4 9 1 9 9 10 9 1 15 0 13 2
32 16 9 15 1 9 9 14 1 9 13 13 7 16 10 9 9 13 2 9 10 9 0 13 2 9 10 9 1 10 9 13 2
15 1 9 15 16 9 9 3 0 1 9 7 9 0 13 2
69 0 13 9 7 9 9 1 9 0 13 16 9 0 2 9 2 9 0 2 9 7 9 1 9 0 1 9 7 9 9 0 7 9 10 9 13 16 3 4 9 10 9 14 16 1 15 0 13 2 3 7 9 7 9 0 9 9 9 13 7 9 15 1 9 9 9 9 13 2
36 16 9 9 2 9 2 9 7 9 16 1 9 13 2 4 1 9 9 9 13 2 7 9 13 16 9 3 9 16 1 9 13 3 0 13 2
26 3 1 9 13 16 9 9 9 3 9 9 9 9 14 1 9 13 7 9 9 0 14 0 13 13 2
29 16 1 9 0 3 1 9 0 9 0 1 9 0 1 9 13 2 0 13 1 9 9 9 10 9 16 9 13 2
75 1 9 9 9 9 7 0 9 0 13 16 1 9 9 15 1 9 0 1 9 9 13 7 1 9 9 16 1 9 9 1 9 0 13 4 9 3 9 9 2 9 9 9 7 9 14 9 13 16 9 0 13 2 1 15 7 9 10 12 9 1 9 9 1 9 9 9 9 1 9 0 9 13 13 2
38 16 9 15 1 9 9 7 9 0 13 13 7 3 15 0 13 7 15 1 9 16 1 9 9 13 2 9 13 1 9 7 15 1 15 0 9 13 2
13 3 10 0 9 2 1 1 10 9 9 13 13 2
29 16 9 13 1 9 16 1 1 9 1 15 9 13 2 9 0 9 13 7 1 9 10 9 12 9 0 9 13 2
27 16 0 9 13 15 1 9 0 1 0 9 1 9 0 0 4 13 7 4 1 1 15 9 0 13 13 2
39 9 0 16 0 9 13 9 12 9 13 16 1 9 15 1 15 9 7 9 9 13 16 3 15 1 9 13 13 7 7 15 7 0 9 15 1 9 13 2
25 3 4 1 10 9 9 0 13 2 16 1 9 0 15 1 15 0 13 7 1 9 1 9 13 2
9 1 10 9 12 9 0 9 13 2
20 1 9 1 9 1 9 9 2 9 1 9 13 13 16 3 9 9 9 13 2
15 1 9 9 9 9 12 16 9 9 1 9 9 0 13 2
10 7 1 9 16 9 9 9 0 13 2
8 16 1 9 9 0 9 13 2
15 1 9 9 0 1 9 0 1 9 9 9 13 13 13 2
12 16 15 14 9 9 13 2 15 9 9 13 2
12 1 9 9 9 0 16 1 10 9 0 13 2
41 1 9 1 12 9 1 9 9 9 1 9 0 16 12 9 9 2 0 1 9 9 13 7 0 9 9 16 9 15 9 9 13 2 9 12 7 12 2 12 2 2
25 1 9 9 9 1 9 9 9 9 13 13 7 1 9 0 9 10 9 1 9 9 9 0 13 2
9 3 9 0 1 9 9 9 13 2
11 16 1 9 10 12 9 1 15 0 13 2
24 9 9 9 13 7 16 1 15 9 9 7 9 14 0 9 13 13 2 9 9 1 1 13 2
30 16 9 9 0 1 9 9 2 9 12 2 9 12 2 12 2 9 13 13 16 9 1 9 9 9 1 1 9 13 2
29 16 9 1 9 9 1 9 2 9 12 2 2 9 9 2 9 12 2 7 1 9 9 2 9 12 2 13 13 2
10 9 9 9 1 9 9 9 13 13 2
9 1 9 10 9 1 9 9 13 2
15 16 1 9 9 0 1 9 7 0 9 15 3 9 13 2
26 1 9 9 2 9 9 9 2 9 12 2 13 13 16 1 15 1 9 15 14 1 9 9 9 13 2
23 1 9 9 1 9 3 13 13 16 15 1 9 12 0 9 9 13 7 1 9 9 13 2
5 3 1 9 13 2
17 3 1 9 1 9 1 9 9 9 13 2 9 2 9 12 2 2
33 1 9 9 16 3 9 2 9 15 9 13 13 7 1 12 0 1 9 1 1 9 7 9 9 1 9 9 9 9 9 9 13 2
74 1 9 9 2 9 15 9 9 9 13 7 1 9 15 1 9 16 9 13 13 2 9 12 2 7 1 9 1 9 9 9 9 1 9 9 1 9 7 0 9 15 9 13 13 2 9 9 2 9 12 2 9 9 13 16 3 1 9 13 7 1 9 12 0 1 9 9 9 15 1 9 15 13 2
10 9 9 9 15 14 12 0 13 13 2
18 9 0 9 10 9 13 16 9 9 7 9 9 2 12 9 0 13 2
33 1 9 15 1 9 7 9 9 9 9 9 0 13 7 1 9 1 9 9 9 1 9 7 9 15 3 1 0 9 9 13 13 2
40 3 1 10 9 13 16 9 9 1 9 0 1 9 13 7 9 9 1 9 3 13 7 1 1 15 9 9 13 7 0 13 16 10 12 9 1 15 0 13 2
9 9 9 9 0 1 9 9 13 2
11 7 9 9 1 9 0 1 9 9 13 2
24 0 15 7 9 9 9 9 14 0 13 16 9 9 9 7 9 9 14 1 15 9 0 13 2
16 9 9 9 1 9 9 9 1 9 1 1 9 9 9 13 2
14 9 9 1 9 9 13 13 16 9 9 14 9 13 2
26 10 9 9 1 9 9 1 9 9 0 13 2 3 1 1 9 9 9 1 9 9 9 7 9 13 2
27 7 15 1 0 9 9 16 9 13 13 7 13 2 3 9 1 9 7 9 7 9 7 9 15 9 13 2
17 1 9 10 9 9 9 9 15 14 1 9 9 0 9 13 13 2
14 1 10 9 15 9 13 16 4 1 1 15 9 13 2
26 1 9 9 1 9 9 9 9 9 9 1 9 9 9 13 16 1 9 9 2 9 7 9 9 13 2
36 7 3 12 9 1 9 9 1 15 9 13 13 2 1 9 7 9 9 15 0 13 2 0 13 16 15 9 0 2 0 13 7 1 9 13 2
12 1 15 9 9 15 1 9 9 0 0 13 2
17 9 9 1 9 13 2 1 10 9 2 9 9 1 9 0 13 2
28 1 9 9 15 1 9 9 13 16 15 1 9 1 9 13 16 1 9 9 13 7 1 9 1 9 4 13 2
14 16 0 13 0 13 7 4 1 10 9 16 9 13 2
41 1 9 9 9 12 9 1 9 9 9 13 7 1 9 15 9 1 9 9 0 1 9 9 13 7 9 16 1 10 12 9 9 13 0 1 9 1 9 15 13 2
27 1 9 1 9 13 13 16 13 9 13 16 1 9 1 9 13 7 3 1 9 7 9 15 9 9 13 2
17 1 10 9 0 13 16 9 1 9 13 7 9 14 1 9 13 2
24 7 9 13 16 15 0 13 7 3 0 13 16 1 3 1 9 13 7 3 13 7 13 13 2
9 16 4 1 9 9 0 0 13 2
10 7 1 9 0 4 1 15 9 13 2
11 16 10 9 1 9 9 0 9 9 13 2
37 15 1 9 1 9 0 13 9 0 7 0 1 9 13 2 7 1 15 9 0 13 16 9 9 1 15 13 7 1 10 9 9 1 15 0 13 2
18 1 9 1 1 12 9 1 9 9 9 7 0 9 9 9 13 13 2
23 9 9 1 9 13 2 1 9 7 9 9 2 9 9 14 1 9 9 1 9 13 13 2
16 7 10 9 3 0 7 0 9 13 7 4 1 15 9 13 2
49 1 1 9 9 2 9 9 13 16 1 9 13 7 1 9 0 9 9 13 2 7 9 9 9 1 9 9 15 0 13 7 9 10 9 16 9 2 9 2 9 9 7 9 9 1 15 9 13 2
10 16 9 0 1 9 9 3 9 13 2
42 1 9 9 9 9 1 9 9 2 9 12 2 7 9 9 2 9 9 9 12 2 12 2 9 1 10 12 9 1 9 13 7 10 9 1 9 10 12 9 13 13 2
19 1 9 9 9 9 16 3 2 1 1 9 7 9 15 9 0 16 3 2
11 9 1 15 13 16 10 9 12 13 2 2
16 1 9 7 1 9 2 9 9 2 9 9 2 9 13 13 2
31 0 15 7 9 9 9 0 13 7 9 9 7 9 1 9 1 15 9 9 15 1 9 7 9 15 1 9 9 0 13 2
19 9 9 16 1 10 9 9 13 13 7 4 1 1 10 9 16 9 13 2
29 1 9 0 9 9 2 16 9 1 9 15 1 9 7 0 9 15 2 9 9 9 2 9 9 12 2 13 13 2
21 9 9 1 9 9 15 14 1 9 12 9 16 1 9 9 0 13 2 13 13 2
12 16 4 15 14 1 3 9 9 0 9 13 2
7 16 9 9 0 15 13 2
22 1 9 9 10 9 1 9 9 0 9 15 0 13 7 9 1 10 9 9 9 13 2
15 1 9 1 9 0 2 9 9 1 9 9 1 9 13 2
25 7 1 9 9 15 0 13 2 16 1 9 0 13 13 16 1 9 9 0 1 9 12 9 13 2
10 7 13 16 1 3 1 9 9 13 2
15 10 9 0 9 13 7 9 9 2 10 9 14 9 13 2
16 9 9 9 1 9 16 0 13 7 0 13 7 4 9 13 2
32 9 9 1 9 1 9 9 1 9 7 9 15 1 9 14 1 9 0 13 13 7 1 3 9 1 9 10 9 9 13 13 2
11 16 4 15 14 1 9 9 0 9 13 2
39 9 9 1 12 9 1 9 9 9 2 9 9 7 9 9 13 13 16 15 1 9 13 7 16 1 9 15 9 13 2 16 9 15 1 9 1 9 13 2
21 9 9 1 9 9 12 9 9 9 14 13 9 2 12 12 12 12 12 12 13 2
14 1 9 1 9 9 2 9 9 0 1 9 9 13 2
22 15 0 1 9 13 2 3 1 9 9 0 13 7 1 9 9 0 2 15 0 13 2
10 3 9 9 1 9 15 9 13 13 2
17 15 1 9 15 14 9 13 7 9 9 10 9 14 9 9 13 2
11 16 9 9 15 1 9 9 0 0 13 2
7 16 10 9 0 9 13 2
15 9 9 1 9 2 9 9 7 9 13 16 1 9 13 2
32 15 16 1 9 15 9 13 7 1 9 0 13 16 1 1 1 9 9 13 7 3 0 13 7 16 4 1 9 0 0 13 2
8 9 1 9 0 3 0 13 2
16 15 9 13 7 1 9 9 9 9 3 13 7 9 0 13 2
21 9 9 15 14 9 9 9 13 13 7 13 13 16 1 9 9 1 9 13 13 2
12 9 9 9 9 13 16 15 1 9 9 13 2
29 1 10 9 4 13 9 15 1 9 9 0 0 13 2 1 3 9 0 1 1 9 1 9 9 10 9 0 13 2
19 7 9 9 1 9 1 9 9 13 13 16 9 0 9 15 0 9 13 2
31 9 16 1 9 1 9 1 9 9 9 13 13 16 15 1 9 9 13 2 7 1 1 9 10 9 1 9 9 13 13 2
21 16 1 9 1 9 9 9 0 9 13 16 3 0 13 16 1 10 9 9 13 2
61 1 0 9 9 9 16 1 15 1 12 9 9 13 13 2 1 1 9 1 9 7 0 9 15 9 13 2 7 12 9 0 13 1 10 9 0 7 0 13 7 9 1 9 0 0 13 16 1 1 10 9 9 13 2 16 9 0 9 0 13 2
40 1 9 1 9 0 4 13 16 9 9 1 9 0 0 13 2 12 2 9 0 16 1 9 13 7 1 1 10 9 1 10 9 9 1 15 1 9 13 13 2
26 12 2 9 9 16 1 9 0 7 9 0 0 1 9 13 16 4 9 10 9 1 9 9 13 13 2
35 1 9 9 10 9 0 13 16 9 9 9 0 9 13 16 0 1 9 14 9 13 13 7 3 15 13 16 13 10 9 14 3 9 13 2
12 3 9 9 0 9 0 9 9 1 9 13 2
6 1 9 9 9 13 2
17 9 15 9 9 9 13 2 3 7 1 15 9 13 9 9 13 2
18 9 10 9 1 15 9 9 13 2 9 10 9 1 15 9 0 13 2
18 3 9 0 16 1 15 3 9 13 2 10 9 16 9 13 9 13 2
17 9 13 0 1 9 15 7 9 9 2 13 1 9 9 9 13 2
17 16 9 9 0 0 13 2 10 9 9 1 9 15 9 9 13 2
18 1 10 9 9 13 10 9 16 3 2 1 9 9 15 9 9 13 2
18 1 10 3 9 9 16 13 0 2 3 3 9 9 9 9 0 13 2
11 9 13 1 9 2 16 3 9 9 13 2
9 1 9 0 0 1 15 9 13 2
49 16 9 9 9 9 3 13 10 9 14 1 9 13 2 0 13 9 1 9 1 9 15 1 1 10 9 0 9 13 16 9 7 9 16 1 9 1 9 13 9 7 9 15 1 9 9 9 13 2
32 9 0 1 10 9 0 16 1 9 0 15 9 7 9 9 14 0 9 15 9 13 13 2 0 9 7 9 15 14 9 13 2
39 1 9 9 0 2 9 2 15 1 9 16 0 9 0 0 7 0 9 0 7 9 0 13 2 1 9 7 9 3 13 1 15 7 3 9 1 15 13 2
15 1 15 9 9 1 9 7 9 15 1 9 9 9 13 2
24 9 9 9 0 14 9 1 9 0 13 16 9 15 14 9 13 7 15 16 9 14 9 13 2
42 3 13 2 8 8 8 2 8 8 8 2 12 2 1 1 9 0 7 0 13 7 1 1 9 0 7 0 13 2 1 9 9 9 13 7 1 9 3 9 16 13 2
11 1 9 10 9 9 7 9 0 13 13 2
30 15 9 1 9 9 9 2 9 2 13 7 15 9 1 9 9 9 2 9 2 13 16 15 15 13 9 1 9 13 2
13 16 9 0 9 9 14 1 1 3 9 9 13 2
32 9 16 13 2 3 7 1 9 0 1 1 10 9 9 13 9 13 1 9 9 7 13 2 8 8 8 2 15 7 9 15 2
13 3 13 2 8 8 8 2 8 8 8 8 8 2
17 16 9 1 9 9 13 2 9 1 9 9 9 1 15 0 13 2
17 9 16 1 10 9 1 9 13 2 8 8 8 8 8 8 13 2
29 7 9 9 0 7 0 9 14 3 9 13 16 1 1 9 0 7 0 13 7 1 1 9 1 9 7 9 13 2
20 1 9 10 9 7 13 13 16 9 13 7 9 2 16 9 13 7 7 9 2
13 9 10 9 0 1 9 8 8 8 8 9 13 2
9 6 2 1 9 9 0 7 0 2
24 9 16 1 10 9 9 15 9 7 9 14 13 7 1 10 9 9 15 1 9 15 0 13 2
9 3 3 9 0 7 3 9 0 2
13 10 9 7 10 9 13 3 15 1 9 9 13 2
32 7 10 9 9 1 9 16 13 2 3 1 9 9 10 9 9 13 2 7 13 2 8 8 8 8 8 8 8 8 8 8 2
18 12 2 6 9 9 1 9 7 9 15 1 1 9 0 14 9 13 2
23 7 1 1 9 9 16 9 10 3 7 3 13 1 9 9 0 9 9 1 15 9 13 2
17 12 2 1 1 9 16 10 9 7 3 9 13 9 4 0 13 2
53 12 2 9 15 14 1 9 1 9 7 9 7 9 1 9 9 13 7 1 15 3 1 9 9 0 13 16 9 7 1 1 9 15 9 13 16 15 12 9 13 2 7 9 0 15 13 7 7 3 15 9 13 2
55 0 9 13 7 9 7 9 1 15 0 13 7 1 9 0 7 7 9 9 1 15 1 13 2 3 7 9 13 7 0 13 16 9 0 1 9 7 9 15 1 15 9 13 15 16 1 9 7 9 15 15 14 0 13 2
23 1 9 9 0 9 9 1 9 16 4 0 13 7 1 10 9 9 0 9 15 9 13 2
20 1 9 9 12 9 0 1 1 15 9 13 13 13 7 1 1 15 13 13 2
12 9 0 1 9 9 0 13 2 8 0 8 2
26 12 2 1 1 9 0 7 0 13 7 1 3 9 9 1 1 9 13 2 8 8 8 8 8 8 2
44 12 2 9 7 9 1 1 15 15 14 1 9 9 0 1 13 2 10 9 16 1 1 9 0 7 0 13 13 1 9 9 0 1 1 9 1 9 9 9 13 7 9 13 2
52 1 3 9 7 9 1 9 9 13 7 9 9 9 9 7 9 15 13 2 9 14 0 13 2 9 9 14 0 13 2 9 9 0 14 9 13 7 3 10 9 7 9 14 1 9 13 16 9 9 13 13 2
39 0 13 1 9 1 12 9 0 0 12 9 13 16 1 9 9 9 0 1 9 9 7 9 9 13 2 3 9 0 16 1 9 9 12 1 9 0 13 2
29 10 9 7 9 9 9 13 2 9 9 0 7 0 13 2 9 9 9 9 7 3 9 14 1 9 9 0 13 2
19 1 15 9 9 1 3 9 13 1 9 9 14 9 13 7 0 9 13 2
17 3 3 1 9 9 3 0 7 3 0 7 3 0 7 3 0 2
4 9 2 9 2
25 9 9 0 9 13 9 9 2 3 2 9 12 9 1 9 3 12 12 9 1 9 14 9 13 2
31 1 9 12 9 0 2 9 9 9 9 0 9 1 10 9 0 9 9 13 7 9 9 9 9 9 0 1 9 13 13 2
25 1 9 9 9 12 0 1 9 9 2 9 9 7 9 1 9 1 9 9 1 9 0 4 13 2
20 1 9 10 9 1 9 9 9 7 9 0 2 9 9 9 1 9 4 13 2
24 9 9 9 9 9 9 0 0 0 1 9 1 9 9 13 2 15 1 9 0 10 9 13 2
27 9 9 9 0 9 0 16 9 9 0 9 13 2 0 9 9 15 14 1 9 9 9 0 9 0 13 2
34 1 10 9 9 9 9 9 0 1 9 9 1 9 1 1 0 9 9 9 13 7 13 2 9 9 0 13 1 9 0 0 0 13 2
22 15 1 9 13 2 16 9 0 0 14 9 13 9 13 1 9 0 9 1 0 13 2
30 9 0 13 2 9 9 0 9 9 13 16 9 9 1 9 12 1 9 9 0 9 1 9 9 7 9 9 13 13 2
31 9 9 0 9 0 16 13 2 1 9 1 9 0 9 1 9 1 9 0 2 9 7 9 9 3 0 1 15 4 13 2
40 9 9 0 9 0 9 13 2 15 13 9 9 0 1 9 0 13 7 1 9 16 9 0 9 1 9 15 13 13 1 9 9 1 9 9 1 9 9 13 2
26 9 9 9 1 9 9 1 9 9 13 2 3 12 12 9 9 1 9 12 12 9 9 9 9 13 2
38 9 9 13 2 9 1 9 12 1 12 9 0 9 1 9 9 9 0 0 2 0 7 0 13 16 9 0 9 1 10 9 0 9 1 9 0 13 2
26 15 13 2 9 15 1 9 12 12 9 9 7 9 9 0 9 2 9 0 9 9 1 9 14 13 2
35 9 13 2 3 12 12 9 9 1 9 12 12 9 9 9 1 9 1 9 13 16 12 12 9 15 1 9 0 7 9 9 0 0 13 2
25 15 0 13 2 16 3 12 12 9 9 2 12 12 9 9 7 12 12 9 9 1 9 9 13 2
43 9 9 9 9 9 0 3 9 2 9 9 7 9 2 9 9 7 9 7 7 9 9 0 1 9 9 1 9 0 14 1 9 9 9 9 1 9 9 9 0 9 13 2
28 9 9 9 0 9 9 0 1 9 1 9 9 7 9 9 0 1 9 7 9 0 1 10 9 14 9 13 2
35 1 10 9 13 13 2 9 0 1 9 9 2 9 0 7 9 0 9 16 12 9 1 12 9 9 1 9 0 0 7 0 9 13 13 2
28 10 9 1 9 1 9 9 9 9 9 13 16 9 0 0 1 9 9 0 12 2 12 12 9 9 13 13 2
31 9 9 9 0 14 1 0 1 1 9 0 0 13 7 9 1 9 7 9 2 9 9 7 9 16 3 0 9 13 13 2
41 1 10 9 16 1 9 9 9 0 1 9 9 9 9 13 7 9 13 13 16 9 9 1 9 0 1 9 0 0 7 9 9 3 1 9 9 0 0 13 13 2
47 10 9 13 2 9 9 9 9 13 13 2 16 9 0 12 12 9 9 0 1 9 13 7 1 3 16 9 9 12 9 9 0 0 12 12 9 1 9 1 9 0 1 9 9 0 13 2
42 9 9 0 9 0 9 9 13 2 1 9 9 0 16 9 9 1 9 9 9 1 9 9 13 13 16 9 9 10 9 9 1 9 1 9 0 9 0 0 9 13 2
17 9 9 9 9 9 13 2 9 9 0 1 9 1 9 0 13 2
40 9 9 9 1 9 10 9 13 2 9 0 2 9 1 9 0 7 0 2 9 9 2 9 0 7 9 9 0 1 9 7 9 0 9 9 0 1 9 13 2
27 15 13 2 9 0 0 9 4 1 9 0 9 13 7 9 0 2 9 7 9 0 9 1 9 9 13 2
24 9 9 9 13 2 9 0 1 9 9 1 9 0 0 9 13 16 4 1 10 9 9 13 2
