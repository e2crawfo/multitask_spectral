8800 17
3 10 9 0
10 10 11 13 10 9 1 10 9 0 2
28 13 12 1 10 3 0 9 1 10 11 2 13 1 11 2 15 13 1 13 10 9 0 7 10 9 1 3 2
67 13 3 10 9 1 10 9 1 2 10 9 1 10 9 2 2 1 0 9 1 10 9 1 10 9 0 2 13 1 11 2 11 2 11 7 9 7 11 2 7 10 9 0 1 10 9 1 10 9 2 15 1 15 13 10 9 2 9 2 1 15 12 7 1 15 12 2
56 3 13 1 13 2 1 10 9 15 13 2 10 10 2 9 0 2 2 9 1 9 1 10 15 13 13 1 10 9 0 3 1 9 1 10 9 1 9 2 1 10 9 2 13 15 1 10 11 7 13 15 1 10 11 2 2
60 7 3 2 1 10 12 9 15 10 11 3 13 1 10 9 1 10 9 13 1 10 9 2 13 13 15 10 9 1 10 9 3 0 2 15 10 9 2 3 1 9 1 10 9 2 13 13 3 1 10 9 2 1 13 10 9 1 10 11 2
33 7 10 9 2 3 13 3 1 10 9 2 2 13 10 9 2 15 13 16 10 9 1 10 9 13 2 13 15 1 9 0 2 2
18 7 3 2 16 15 3 13 2 1 10 10 9 2 1 10 9 0 2
56 2 13 15 1 9 3 2 16 2 16 10 9 13 1 4 13 2 15 3 13 3 2 16 2 1 10 9 2 2 10 9 0 13 10 9 2 10 15 3 13 3 15 13 13 1 10 11 2 2 13 13 9 1 10 9 2
24 15 13 4 1 13 10 9 2 3 16 2 1 10 9 2 10 9 1 10 11 13 3 13 2
18 15 3 3 13 2 3 15 1 11 2 7 15 13 4 1 13 9 2
5 10 9 1 12 9
6 2 9 2 1 10 9
48 10 0 9 0 1 2 9 2 1 9 2 10 9 0 11 2 13 10 9 1 10 9 13 15 13 9 1 11 2 11 2 10 9 0 13 2 11 2 15 13 13 10 9 1 2 9 2 2
17 1 10 9 2 10 9 13 16 10 9 13 7 13 10 9 0 2
24 2 13 1 13 10 9 1 10 0 9 2 13 11 2 9 1 9 1 10 11 1 10 11 2
45 10 11 13 13 1 10 11 1 3 12 9 7 13 15 1 10 9 7 1 10 9 15 15 13 13 3 1 10 9 2 13 4 13 1 10 9 1 12 9 0 2 12 9 2 2
21 11 13 3 13 1 10 9 1 3 13 13 1 10 9 3 1 13 1 10 9 2
29 11 2 15 13 10 9 1 11 1 10 9 1 9 1 11 2 3 3 13 1 10 9 15 10 9 0 15 13 2
22 2 3 13 1 13 16 2 1 13 10 9 2 15 13 1 13 3 10 9 2 13 2
11 2 10 9 9 13 10 9 1 13 2 2
23 11 13 3 16 2 1 10 0 0 2 10 11 13 10 10 9 12 9 3 1 10 9 2
1 11
15 3 1 10 11 2 10 9 13 1 10 9 0 3 13 2
42 10 9 0 2 1 10 9 2 9 0 1 2 9 2 7 1 9 2 13 9 0 1 10 10 9 2 3 1 9 2 10 3 11 2 11 2 11 2 11 7 11 2
44 10 12 0 9 13 15 1 13 10 9 1 11 1 10 9 7 10 0 2 10 0 1 9 1 10 9 0 2 13 13 1 10 9 1 11 2 11 2 2 15 13 0 9 2
25 10 2 9 9 2 0 2 1 9 1 10 11 2 13 15 1 13 10 9 1 10 9 1 9 2
8 15 2 3 13 2 3 13 2
5 12 9 1 12 9
32 10 9 2 1 13 1 9 1 10 9 1 0 2 13 1 10 11 2 13 13 1 12 9 1 9 2 9 0 1 10 11 2
11 1 3 3 10 11 13 13 1 10 9 2
58 2 10 9 13 3 3 13 2 16 13 3 0 16 16 13 3 10 9 1 9 1 10 9 2 2 13 10 9 11 2 1 10 9 1 10 11 2 13 16 2 1 10 9 0 2 2 16 10 9 13 13 2 15 13 1 13 2 2
40 1 15 3 12 9 1 10 9 0 1 10 11 2 11 2 2 10 9 1 9 3 13 1 10 9 1 10 9 1 9 1 10 9 3 13 3 13 1 13 2
11 10 0 9 13 1 10 11 3 13 9 2
29 12 9 2 13 12 9 2 13 3 1 13 1 10 9 13 1 13 9 13 0 1 9 7 9 1 9 13 3 2
36 10 9 2 1 15 10 11 13 9 2 13 1 10 9 13 16 10 9 1 9 13 1 10 11 13 12 9 1 10 0 9 1 12 1 9 2
40 10 9 2 13 1 10 9 1 13 10 9 1 9 2 1 13 10 9 1 10 9 0 1 1 10 9 12 1 9 2 2 13 1 10 11 10 9 2 11 2
29 1 15 2 13 10 0 2 2 13 13 10 9 2 10 9 13 13 7 2 1 15 2 10 9 15 13 13 2 2
27 7 15 13 10 9 16 10 9 13 1 13 10 9 1 10 11 13 1 13 9 1 10 9 0 1 9 2
25 10 9 1 10 9 3 13 2 3 2 13 3 1 10 9 0 1 10 9 1 15 3 12 9 2
18 3 0 13 10 9 2 11 2 15 13 10 9 1 2 10 9 2 2
27 16 13 10 9 2 15 13 10 9 1 9 1 10 9 15 13 10 9 2 15 1 15 13 10 9 2 2
34 1 16 3 13 9 2 9 13 1 10 9 16 15 13 1 10 9 1 10 9 1 10 9 2 1 10 9 15 13 1 2 9 2 2
48 3 2 1 10 11 2 15 3 13 13 2 10 9 1 10 0 9 1 10 9 0 13 1 10 9 1 11 1 13 10 9 1 10 11 0 2 3 2 10 9 13 1 10 9 1 10 11 2
40 1 10 9 1 9 1 10 9 2 11 13 1 3 12 12 9 16 2 10 11 13 1 10 9 0 7 16 10 9 13 4 13 1 10 9 1 10 9 2 2
27 3 13 1 10 9 1 10 9 2 10 9 0 13 16 2 13 10 9 1 15 10 11 13 10 9 2 2
19 10 9 0 13 1 9 0 7 9 1 9 0 1 10 9 0 7 0 2
5 10 9 1 10 9
50 9 0 2 2 11 2 13 15 1 10 9 1 11 2 9 1 11 2 13 10 9 1 11 15 2 13 12 9 2 13 13 10 10 9 0 1 15 13 1 10 11 1 10 9 2 9 1 10 9 2
76 13 10 9 1 10 9 1 11 2 1 10 9 13 2 10 9 1 10 9 2 11 2 13 16 10 9 0 15 13 1 10 9 1 11 2 2 7 3 15 13 1 10 9 1 10 11 15 13 2 1 9 0 2 10 9 13 1 10 9 1 10 9 1 10 9 15 15 13 1 10 9 1 10 11 2 2
17 1 10 9 1 10 11 2 10 9 1 9 13 3 1 10 9 2
25 2 15 3 13 0 1 13 1 10 9 0 2 7 13 16 15 13 10 9 0 1 10 9 0 2
21 7 16 12 1 10 10 9 13 10 9 1 10 9 0 2 15 3 15 13 2 2
3 9 2 11
3 9 2 11
12 10 0 9 1 11 2 15 3 3 13 13 2
14 11 13 11 2 10 9 2 1 15 13 10 9 0 2
1 11
24 1 10 0 9 15 13 10 9 1 10 11 2 10 9 11 13 10 9 15 3 13 10 9 2
19 0 2 0 2 13 2 13 10 11 10 11 7 3 10 9 13 13 15 2
17 11 2 13 1 10 0 9 1 10 11 2 10 9 1 9 0 2
20 1 10 10 9 3 13 10 9 2 16 10 9 1 10 9 3 13 0 9 2
33 13 3 15 13 10 9 7 3 13 1 10 9 10 0 9 1 9 2 7 13 16 13 1 9 7 3 1 9 2 3 13 3 2
31 1 13 10 9 0 1 10 9 0 2 13 3 1 10 9 10 10 9 2 10 13 1 10 9 11 2 1 15 15 13 2
13 10 9 15 10 9 9 13 2 3 13 15 2 2
4 13 15 2 2
35 2 13 15 13 2 3 2 16 15 13 1 10 9 0 2 3 13 1 10 9 11 2 15 13 2 3 2 13 10 9 1 10 9 11 2
73 9 0 2 15 10 15 13 13 2 3 0 2 13 3 16 2 1 10 9 13 1 10 9 9 15 2 1 9 2 15 3 13 13 10 9 1 10 9 2 11 2 2 10 9 1 10 9 11 3 15 15 13 1 10 10 9 1 9 7 2 3 2 2 10 13 9 1 10 9 1 10 9 2
26 10 11 13 3 1 13 10 11 1 10 9 0 2 12 2 2 13 1 10 9 1 10 11 1 9 2
37 10 9 13 1 13 13 1 10 9 1 11 2 3 16 10 11 13 3 3 2 12 2 7 10 9 0 3 13 13 15 1 10 9 1 10 9 2
40 7 10 9 0 7 0 1 11 2 3 3 3 13 13 9 1 9 2 13 2 3 3 2 1 10 9 1 11 2 13 10 9 1 13 10 9 1 10 9 2
25 10 11 13 10 10 9 0 2 1 11 7 11 3 13 7 13 1 10 9 1 11 1 10 9 2
28 3 2 10 11 13 1 12 9 2 1 10 9 11 2 1 3 2 1 13 10 9 7 10 9 11 3 0 2
27 3 3 13 3 10 12 9 2 11 2 11 7 11 2 2 13 11 10 9 1 2 9 2 1 10 9 2
55 1 15 2 7 3 16 10 9 13 3 3 13 1 10 3 13 7 0 9 2 10 11 13 3 0 1 10 9 2 13 10 0 9 1 10 9 1 10 9 0 1 10 9 2 13 1 10 9 7 10 9 1 10 11 2
11 10 2 9 2 15 11 13 13 3 0 2
52 7 13 15 3 16 10 11 7 10 9 2 13 2 1 9 1 10 9 13 2 10 9 7 10 9 1 10 9 3 9 1 9 0 1 10 0 0 2 3 3 13 1 9 1 12 2 1 0 1 10 0 2
11 10 9 0 13 3 1 10 9 3 0 2
39 7 9 1 10 9 13 2 3 2 10 9 0 1 10 11 2 15 13 3 1 13 10 9 3 9 7 3 3 10 9 1 10 10 9 1 10 9 0 2
6 9 7 9 1 10 9
29 3 1 9 7 9 3 13 2 1 10 9 1 10 13 9 2 10 9 1 10 9 7 1 10 9 1 10 9 2
50 13 10 9 0 7 0 1 10 11 2 1 10 0 9 2 7 3 10 9 13 13 9 1 10 10 9 2 15 15 13 3 1 13 10 10 9 1 10 9 2 1 15 15 13 7 1 10 0 9 2
45 12 10 11 13 13 1 10 9 0 9 10 0 9 7 2 1 10 10 9 2 13 10 2 0 2 2 2 11 2 7 2 11 2 2 1 13 10 10 9 7 3 10 10 9 2
43 9 1 9 0 2 11 12 2 2 11 2 2 2 1 9 9 2 11 12 2 2 11 2 2 2 1 9 0 2 11 12 2 1 9 0 2 11 12 2 2 9 2 2
1 11
4 11 2 12 2
35 3 1 10 0 9 1 10 11 2 13 1 11 7 11 2 11 13 13 15 3 10 2 0 9 2 1 10 2 0 9 2 2 11 2 2
59 10 11 2 15 13 10 9 1 12 2 13 13 0 1 13 10 10 9 1 9 2 7 13 11 7 11 1 13 10 10 9 0 1 15 13 13 10 9 0 1 15 13 1 10 9 1 11 1 13 10 9 7 15 13 10 12 12 9 2
39 10 2 9 2 13 0 10 0 9 1 10 0 9 1 9 2 3 12 1 15 10 9 2 2 15 13 13 10 9 13 2 3 1 10 9 15 13 0 2
33 3 2 10 9 1 11 2 9 1 10 9 0 1 12 2 13 9 1 10 11 1 13 11 1 13 10 0 9 1 11 7 11 2
9 15 1 10 12 9 13 10 9 2
6 3 2 15 13 9 2
11 10 9 16 10 9 1 9 13 3 0 2
37 11 16 10 9 13 3 0 2 10 11 13 10 9 1 10 9 3 1 10 10 9 7 13 3 10 9 1 9 16 10 9 2 1 9 1 11 2
37 11 7 11 16 10 9 13 3 0 2 7 7 0 7 0 16 1 10 0 9 1 10 9 7 10 11 13 3 0 7 13 1 9 1 9 0 2
21 1 10 9 2 15 13 15 1 12 9 0 2 3 7 3 1 10 9 1 11 2
38 3 2 10 11 13 10 9 2 1 9 1 11 2 1 10 9 1 10 9 13 1 11 2 7 13 10 9 15 3 15 13 1 10 9 1 10 9 2
36 3 2 10 11 13 9 1 10 9 2 13 10 9 1 9 7 13 10 9 3 1 10 0 9 13 1 11 2 1 13 9 1 11 1 11 2
20 1 10 9 1 9 2 10 9 13 1 9 0 10 9 15 13 1 10 9 2
43 1 10 9 1 10 9 1 9 13 2 13 13 3 0 9 10 9 1 10 9 0 3 1 10 9 0 2 7 10 0 9 7 10 9 1 10 9 1 10 9 7 9 2
1 11
1 11
10 11 13 0 9 1 10 11 1 10 11
59 10 11 2 11 2 2 9 1 10 9 1 12 1 9 2 13 10 0 9 1 10 11 1 10 11 2 9 1 15 11 13 1 12 2 1 2 3 2 13 10 10 9 0 1 15 1 10 11 2 3 1 10 9 1 10 9 1 12 2
35 10 9 15 13 10 0 9 1 10 11 7 1 10 11 7 15 3 13 10 9 1 10 9 1 11 2 10 0 0 9 0 1 10 9 2
48 10 9 13 12 1 10 12 9 0 13 1 11 3 7 3 2 1 10 11 2 1 10 11 2 3 15 13 10 9 1 12 9 1 0 2 10 9 1 10 15 13 12 9 15 13 1 11 2
31 3 2 1 10 9 0 1 10 11 7 1 10 10 9 1 10 9 2 10 9 13 1 10 0 12 9 1 10 0 11 2
29 1 15 13 2 1 10 12 9 2 11 2 1 3 2 1 10 9 1 11 2 11 13 13 1 10 9 1 9 2
18 3 10 0 9 3 11 13 2 3 9 2 10 9 1 10 10 9 2
41 7 13 15 16 10 10 9 1 12 9 2 1 13 1 10 11 1 11 2 13 13 10 9 3 1 10 10 0 9 1 10 11 2 1 12 1 12 1 9 13 2
20 11 13 3 9 1 13 16 10 9 1 9 1 10 9 13 3 1 10 9 2
12 2 16 13 13 2 15 13 3 0 16 15 2
18 15 13 2 10 9 11 13 2 16 13 13 2 6 2 2 2 13 2
4 7 16 13 2
11 2 15 13 3 1 3 16 10 9 11 2
4 13 13 2 2
5 7 13 10 9 2
8 2 10 9 13 13 3 0 2
15 13 15 3 15 13 13 1 10 11 16 10 9 13 2 2
4 9 0 13 6
4 1 10 10 9
4 11 2 1 11
12 3 1 10 11 10 9 13 13 1 9 0 2
39 10 9 1 10 9 1 10 9 1 13 15 3 13 1 10 9 2 13 9 0 2 15 13 10 9 1 13 10 9 2 1 10 9 1 10 9 0 2 2
44 10 11 2 10 9 13 13 1 13 2 13 13 1 10 9 1 9 2 9 2 9 3 7 9 1 15 10 9 1 10 9 11 1 2 10 0 7 13 2 13 13 3 9 2
47 13 4 1 13 10 9 1 9 1 10 11 2 10 9 2 1 10 9 1 10 0 9 2 13 10 9 0 1 11 2 10 9 13 3 2 15 10 10 9 15 10 9 13 1 10 9 2
12 13 2 1 10 9 2 10 10 9 1 9 2
10 9 1 11 2 11 3 2 13 2 9
37 11 3 13 10 0 9 15 13 9 1 9 1 10 9 1 11 2 15 13 16 2 1 15 15 13 0 2 10 9 3 13 10 9 1 10 11 2
31 3 2 13 1 13 1 10 9 2 3 1 10 9 2 10 9 1 16 10 9 12 13 12 9 2 0 2 1 10 9 2
45 13 15 16 10 9 1 11 3 13 10 9 0 2 7 3 2 0 2 2 3 2 10 9 10 9 13 16 13 10 9 2 13 1 2 11 2 2 1 15 13 10 9 1 9 2
45 10 9 2 3 13 1 10 9 15 15 13 1 10 11 1 10 9 2 13 15 16 11 13 10 9 1 10 11 2 11 13 2 0 7 3 2 2 13 2 1 10 9 1 11 2
24 3 2 3 1 10 2 9 2 2 0 1 0 2 9 2 2 3 10 9 0 3 15 13 2
15 1 12 3 13 1 10 9 10 9 1 10 2 0 2 2
49 10 0 9 1 10 11 13 13 13 15 15 2 13 10 9 2 13 10 9 1 10 9 2 10 9 0 1 10 11 2 11 2 2 15 3 13 10 16 10 9 1 10 9 3 13 1 10 9 2
56 1 9 0 7 1 9 2 10 9 1 11 3 15 13 1 13 10 11 2 10 9 13 2 3 2 13 1 10 11 2 11 2 2 1 10 0 9 0 1 10 11 2 15 3 13 1 15 9 1 10 0 9 1 10 11 2
44 3 2 1 12 9 2 3 10 11 13 3 13 2 1 10 9 15 13 2 1 10 9 2 1 9 0 2 10 11 2 7 15 15 13 10 9 1 10 0 2 10 11 2 2
38 11 15 2 1 10 9 2 13 3 13 2 3 1 10 9 1 10 9 2 3 15 13 10 11 7 10 11 2 2 3 1 10 11 13 1 10 11 2
19 10 9 13 1 10 9 1 12 2 1 10 9 1 11 2 1 10 11 2
40 10 9 13 1 9 1 10 9 1 10 9 1 9 2 3 10 9 0 1 0 1 10 0 9 0 13 1 10 9 1 11 2 1 10 10 9 2 10 11 2
21 10 9 1 10 9 13 1 10 9 15 10 9 13 3 10 2 9 1 11 2 2
53 1 10 9 2 10 11 2 11 2 13 1 10 9 1 10 9 0 2 10 9 0 11 13 1 4 13 2 7 10 9 2 13 1 13 1 11 1 10 9 1 10 9 1 12 2 13 3 13 9 1 10 11 2
5 10 9 1 10 9
34 10 0 13 16 2 3 3 2 11 13 15 16 10 9 0 13 4 1 10 10 9 7 4 1 10 11 2 10 9 1 10 0 9 2
31 2 13 1 10 9 1 9 2 2 13 13 10 9 11 0 2 13 1 9 2 7 12 9 2 7 13 15 1 10 11 2
12 12 1 10 0 2 11 2 13 1 10 9 2
10 2 13 10 10 9 2 13 13 2 2
13 3 3 2 10 9 13 15 10 9 1 10 9 2
25 1 10 9 15 15 13 2 13 10 0 9 2 3 12 9 2 7 10 12 9 13 1 10 9 2
34 1 1 10 9 0 11 2 13 1 10 11 2 10 9 7 9 13 16 13 1 1 10 12 9 1 3 1 2 3 2 13 10 9 2
28 13 1 10 9 1 11 1 10 9 2 10 0 9 13 13 1 9 1 10 12 9 0 1 13 9 3 3 2
56 1 10 12 9 1 10 9 2 10 9 1 9 1 10 9 13 13 3 7 1 12 9 10 9 13 1 10 9 2 0 1 13 9 1 10 9 1 1 10 9 15 13 10 9 1 9 1 10 9 11 2 1 10 9 0 2
21 10 9 1 10 9 3 13 10 0 9 1 10 9 1 10 9 3 10 9 13 2
52 10 9 13 10 3 13 9 1 10 9 2 3 9 2 9 0 2 9 0 7 1 9 3 1 10 9 1 9 10 9 1 10 11 3 13 10 9 7 9 1 9 1 10 9 1 9 15 13 1 10 9 2
20 3 1 10 9 0 1 10 9 2 10 2 9 0 2 13 3 1 12 9 2
18 10 11 13 13 10 11 1 12 9 1 9 2 12 9 1 9 2 2
32 10 11 13 10 2 9 2 7 10 2 9 2 15 13 13 10 9 1 9 2 3 10 15 13 1 10 9 1 10 10 9 2
44 10 9 0 1 10 9 3 13 13 0 7 10 9 13 1 10 9 1 10 9 3 3 12 9 1 10 11 1 13 10 11 1 10 9 13 1 9 7 9 1 10 9 0 2
17 10 11 13 10 3 0 9 1 2 9 2 1 9 1 10 11 2
3 11 13 9
21 10 11 2 10 0 0 9 0 1 9 2 13 13 10 9 1 10 10 9 0 2
25 10 9 13 13 3 0 10 9 1 10 9 2 15 13 1 13 10 0 9 1 10 10 0 9 2
14 10 9 13 2 3 10 9 2 1 12 7 12 9 2
46 1 10 0 9 1 10 0 9 2 10 9 1 9 0 1 10 11 13 10 9 1 12 9 1 0 9 1 10 9 0 2 1 10 9 1 12 9 1 9 2 12 9 1 9 2 2
4 9 1 10 11
43 10 9 13 1 10 9 1 10 11 13 16 10 9 1 9 0 2 13 1 10 11 2 1 9 1 9 1 10 0 12 9 1 13 13 0 1 10 9 1 9 1 11 2
18 10 3 9 3 13 4 13 1 9 0 3 1 10 9 1 10 0 2
21 10 9 1 10 9 13 15 1 9 13 1 10 9 1 13 10 9 7 13 9 2
75 10 9 0 2 1 10 9 1 15 13 9 1 10 9 1 2 10 9 2 1 10 9 2 13 1 10 9 16 3 13 10 0 7 1 10 9 1 10 9 2 11 2 7 1 10 9 0 2 11 2 7 16 13 1 10 0 9 10 9 0 2 1 16 15 13 13 10 9 1 10 0 2 1 2 2
35 13 15 3 1 10 9 16 3 13 1 10 9 0 7 1 10 0 7 1 10 0 7 16 13 10 9 1 10 10 9 2 9 7 9 2
10 2 2 9 2 11 2 1 10 11 2
3 10 9 0
8 3 13 10 9 2 13 15 2
14 3 13 11 13 15 15 13 1 10 9 1 10 11 2
12 3 13 2 7 2 3 3 13 9 0 2 2
16 3 3 15 15 13 1 16 10 0 0 13 13 10 10 9 2
21 10 9 13 2 3 0 2 10 9 3 13 7 15 13 1 13 15 1 0 9 2
21 3 3 13 1 10 9 0 1 13 1 10 9 1 9 0 1 10 2 9 2 2
26 13 1 15 13 1 10 9 1 10 11 1 11 2 1 13 10 2 9 2 15 3 13 9 1 9 2
3 13 9 2
12 13 9 2 3 3 13 10 9 1 10 9 2
6 1 10 9 13 12 2
2 11 13
18 10 9 1 11 1 10 11 13 1 13 10 9 1 10 9 0 0 2
14 13 10 9 0 2 10 0 9 0 2 1 10 9 2
14 10 9 2 3 0 2 13 1 13 3 3 13 9 2
19 3 2 13 1 13 15 10 9 1 10 9 1 10 0 9 1 10 9 2
13 10 9 11 13 12 9 2 13 1 10 12 9 2
6 11 13 9 1 10 9
4 9 2 0 2
43 10 11 13 3 2 3 0 2 13 1 10 9 1 9 1 10 9 1 10 9 0 15 2 1 13 15 2 13 13 10 9 1 10 9 1 11 1 3 12 9 1 12 2
32 10 9 13 13 1 13 3 10 9 1 10 9 2 9 0 1 10 9 1 10 9 2 2 15 3 13 13 1 9 13 3 2
27 1 10 9 2 10 9 13 15 2 3 1 9 1 10 9 0 7 12 1 9 1 10 0 9 0 2 2
20 1 11 2 10 9 13 1 9 1 9 1 9 2 1 9 1 10 10 9 2
13 3 2 13 13 15 10 9 13 3 3 15 13 2
21 2 3 2 10 9 13 1 13 10 9 0 2 2 13 10 10 0 1 10 11 2
14 10 9 1 9 13 15 1 9 0 2 1 10 9 2
14 1 10 9 1 10 9 2 13 10 9 1 10 9 2
25 2 10 0 9 1 10 9 13 13 10 9 7 13 1 10 9 0 10 9 7 9 1 13 13 2
11 10 9 13 1 15 2 2 13 10 11 2
36 1 10 11 2 10 9 13 10 9 3 2 1 10 9 1 9 0 2 3 9 1 10 9 1 11 7 11 1 10 11 13 3 13 10 9 2
14 10 9 13 13 3 1 9 2 2 1 9 3 2 2
39 1 10 9 10 0 9 13 10 9 1 3 15 13 13 1 10 9 1 10 9 0 3 10 9 13 2 16 15 3 13 9 13 1 10 9 1 10 11 2
7 7 3 13 15 0 9 2
16 10 9 1 9 0 15 13 13 1 11 7 10 10 9 0 2
18 13 0 13 1 10 9 0 1 10 11 2 10 9 0 0 7 11 2
20 10 9 13 16 10 9 0 13 13 10 9 0 1 10 9 2 1 10 9 2
6 15 13 3 10 9 2
44 0 1 10 9 13 10 9 1 0 9 2 3 1 9 3 1 9 2 7 1 11 2 1 10 9 15 2 1 10 0 9 1 10 10 9 7 1 10 9 2 13 1 13 2
29 15 1 10 9 13 10 9 2 13 15 12 9 1 9 1 9 7 10 9 1 12 12 1 12 12 9 1 9 2
24 1 10 13 9 1 10 9 2 11 13 16 2 10 9 3 13 13 1 9 2 7 1 9 2
27 13 15 16 10 11 7 10 11 13 13 1 10 11 7 10 11 7 10 11 1 10 11 2 7 13 9 2
8 3 15 13 10 10 9 2 2
26 1 10 9 1 10 11 2 10 9 11 3 13 9 1 9 13 7 13 10 0 9 3 10 3 0 2
19 2 13 16 10 11 3 13 1 15 13 1 10 11 2 3 13 1 15 2
16 10 9 1 9 13 13 0 9 7 15 3 13 13 10 9 2
16 15 13 10 9 1 9 7 3 13 13 15 13 3 0 2 2
6 9 2 3 13 0 2
16 13 13 1 11 2 7 3 13 13 15 1 13 7 1 13 2
21 3 13 10 9 1 10 9 2 7 13 9 2 16 13 16 15 13 15 1 13 2
11 9 2 3 13 10 10 9 1 10 9 2
4 2 3 13 2
4 3 0 2 2
15 1 10 9 2 3 13 10 9 1 13 1 9 2 9 2
50 13 1 10 9 15 1 9 13 10 0 9 1 11 2 13 3 12 9 1 10 3 13 9 1 10 11 2 15 15 13 13 1 10 9 10 9 1 10 11 13 1 10 9 15 15 13 1 10 9 2
63 13 16 10 9 1 13 10 9 13 1 10 9 1 10 9 2 11 2 3 9 1 11 7 11 2 15 1 10 9 13 2 3 9 1 10 9 2 2 10 9 1 9 0 15 13 10 10 9 2 2 2 10 0 9 13 1 13 10 9 1 10 9 2
72 2 10 9 1 10 9 13 0 2 10 0 9 13 1 9 7 9 2 1 10 11 1 10 9 1 10 9 2 3 1 9 7 9 2 15 1 3 3 15 13 3 1 13 1 10 9 1 10 9 1 11 2 13 15 10 11 2 15 13 13 10 9 3 7 13 9 1 13 9 2 2 2
30 13 1 13 9 10 9 1 10 11 1 13 10 9 0 1 13 10 9 1 10 11 2 1 10 9 1 10 9 9 2
18 10 10 9 3 13 16 10 9 3 13 9 7 13 13 1 10 9 2
27 3 10 9 0 13 2 1 12 2 10 9 1 10 11 2 3 3 13 1 10 11 2 13 10 0 9 2
28 3 10 0 7 0 9 1 10 9 2 3 13 10 11 1 10 9 0 2 1 10 9 15 13 10 10 9 2
51 10 9 1 10 9 2 1 10 9 1 10 11 13 1 10 9 0 1 10 9 0 2 3 10 0 9 1 9 1 10 9 2 3 10 9 1 10 9 1 10 9 1 10 10 9 15 13 10 9 0 2
34 3 2 15 1 10 9 13 1 10 11 2 13 16 10 11 13 4 2 13 2 1 10 9 7 16 13 0 9 1 10 9 1 12 2
33 3 1 10 12 9 2 13 10 0 9 1 10 0 9 0 1 10 9 0 1 10 9 1 10 9 2 3 2 3 2 10 11 2
11 10 9 3 13 1 10 9 13 1 11 2
27 2 13 3 0 16 10 11 13 13 1 10 9 1 10 11 2 2 13 1 10 11 10 9 1 10 9 2
32 1 10 9 1 10 9 2 13 15 3 10 9 1 10 11 15 2 1 10 0 9 1 10 9 0 2 13 1 13 12 9 2
20 13 15 3 12 12 9 2 1 10 9 1 9 1 13 15 1 10 12 9 2
12 2 10 9 15 13 1 10 9 1 10 9 2
13 13 10 0 9 1 10 0 2 2 13 10 0 2
4 11 13 1 11
14 11 13 10 0 9 15 13 13 3 1 10 12 9 2
24 3 2 1 10 9 1 9 3 0 2 13 10 9 1 9 1 0 9 13 1 9 1 9 2
37 7 13 3 13 1 9 3 15 1 10 9 0 11 15 13 10 9 0 7 0 7 3 10 9 0 1 10 1 10 10 12 9 1 9 1 9 2
20 1 9 2 13 3 10 9 1 10 11 13 13 1 10 9 1 9 3 0 2
39 1 9 1 12 2 13 15 10 9 1 10 11 1 10 9 15 13 10 9 0 1 10 9 1 9 0 2 1 13 13 9 1 10 9 1 10 9 0 2
24 1 10 10 9 2 13 1 13 10 9 0 15 13 13 3 3 10 9 1 10 9 1 9 2
36 15 13 13 10 9 1 13 2 7 10 9 1 16 10 9 13 13 1 10 9 1 9 0 15 13 3 1 13 3 13 10 10 2 9 2 2
33 3 2 10 9 13 15 1 16 10 9 13 1 13 1 10 9 1 11 1 10 9 1 9 1 10 9 1 10 9 1 10 9 2
24 1 9 0 13 1 10 2 11 2 2 10 9 13 4 13 1 10 0 9 1 10 9 11 2
34 16 11 13 13 2 1 9 13 2 10 10 9 2 1 12 9 2 13 1 13 15 2 3 1 10 9 1 9 0 1 10 9 0 2
36 3 1 10 9 1 9 2 11 13 1 13 10 9 0 1 10 0 9 1 10 9 2 13 1 10 9 1 13 9 0 1 15 15 13 0 2
21 10 9 13 0 9 11 7 10 10 9 13 4 13 3 10 9 1 10 0 9 2
18 10 9 7 9 2 13 2 3 10 9 0 1 10 11 2 1 11 2
13 1 15 13 11 2 10 9 1 10 9 1 10 11
28 11 2 9 2 7 11 2 9 1 10 11 2 13 15 1 10 9 1 10 11 1 9 13 1 10 9 1 9
17 11 3 13 13 10 9 0 16 13 13 11 2 13 10 9 0 2
12 10 9 13 10 9 7 13 15 1 10 11 2
10 10 0 9 1 10 9 13 1 4 13
24 1 10 10 9 13 15 9 15 13 1 10 9 0 11 2 3 15 13 1 15 13 13 13 2
46 10 11 13 3 10 9 1 13 9 1 10 9 1 11 2 9 2 2 11 2 9 2 7 11 2 9 2 2 15 13 1 10 11 2 1 10 9 1 10 0 13 10 9 1 9 2
28 3 11 13 13 2 1 10 9 1 10 9 13 1 9 0 13 1 10 11 7 11 2 3 15 13 10 9 2
24 16 11 13 0 2 15 13 10 9 7 3 10 9 3 13 3 0 1 10 9 1 10 11 2
11 15 13 10 9 15 3 3 13 1 9 2
31 3 2 1 10 9 13 1 10 9 1 10 11 2 10 9 2 13 1 10 9 2 3 13 10 9 15 13 13 10 9 2
15 1 10 9 2 3 13 13 1 10 9 1 2 13 2 2
3 9 7 9
15 11 3 13 15 13 10 9 2 7 3 13 9 1 13 2
4 2 3 13 2
13 3 2 10 9 1 10 9 13 13 1 10 9 2
21 3 13 11 2 1 10 11 2 15 13 10 9 1 9 0 1 10 9 1 11 2
28 2 13 16 9 0 7 0 13 1 10 9 15 13 1 9 1 10 9 1 10 9 1 10 9 1 10 9 2
30 10 9 2 10 9 2 10 9 2 10 2 9 2 1 10 11 15 13 13 15 13 10 9 1 10 2 9 2 2 2
115 10 9 13 13 12 2 2 11 2 2 9 1 10 9 0 13 10 9 1 10 9 0 2 2 2 11 2 2 11 3 9 1 9 7 9 1 10 9 0 7 0 1 10 9 2 2 2 11 2 2 11 3 9 1 9 7 9 2 9 0 1 10 9 1 9 0 2 2 2 11 2 2 11 3 9 13 1 9 0 2 1 10 9 1 9 1 9 2 7 2 11 2 2 11 3 9 1 9 1 10 9 0 2 13 10 9 1 10 9 1 9 1 9 2 2
6 11 2 9 2 13 2
28 2 1 10 0 9 10 9 13 13 1 10 2 9 2 1 10 11 2 1 9 0 7 15 13 9 1 11 2
40 10 9 1 10 11 13 12 9 1 9 1 11 7 1 10 9 0 1 10 11 2 1 10 9 1 9 7 9 1 10 9 2 1 10 9 0 1 10 9 2
12 3 2 13 13 9 1 9 0 1 10 9 2
14 13 15 13 1 10 9 0 2 16 13 10 9 3 2
38 7 13 15 10 9 2 3 13 10 9 2 13 9 2 3 16 13 9 13 1 13 15 7 13 9 1 12 2 9 2 15 13 9 0 1 11 2 2
16 10 0 9 13 13 1 10 9 1 10 9 13 1 10 11 2
22 1 10 0 9 10 9 13 15 0 2 2 13 15 3 0 9 7 9 2 2 13 11
18 1 10 11 2 10 12 9 1 10 9 13 10 9 0 1 10 9 2
12 13 0 1 9 2 9 1 9 0 1 9 2
25 10 9 13 9 1 9 1 9 1 13 9 1 9 1 10 9 13 1 10 9 1 10 11 13 2
15 13 10 9 0 1 13 13 10 9 2 7 13 15 3 2
12 9 2 11 2 11 2 7 11 2 11 2 2
24 11 2 11 2 11 2 11 2 11 2 11 2 11 2 12 2 2 11 7 11 2 12 2 2
13 13 10 9 3 13 10 0 9 0 1 10 9 2
22 1 10 9 13 15 1 10 9 1 9 15 3 13 7 15 13 10 9 1 9 0 2
15 3 15 13 0 3 13 13 10 9 1 10 2 11 2 2
21 13 13 16 3 15 15 13 2 3 15 15 13 13 3 13 1 10 0 9 0 2
48 13 1 10 9 14 9 0 2 3 13 1 9 1 3 13 10 9 1 10 10 9 2 1 10 9 3 13 2 15 3 13 12 1 10 9 15 13 1 10 9 12 1 10 10 9 10 9 2
12 10 9 13 1 10 9 13 1 10 9 3 2
14 13 10 9 1 10 9 15 15 13 2 2 11 2 2
17 1 15 15 13 3 13 0 1 10 9 2 10 9 13 9 0 2
9 3 10 10 9 13 9 7 15 2
21 3 2 3 2 13 10 9 0 1 10 9 15 15 13 9 13 3 10 9 0 2
21 3 13 0 13 16 13 10 9 1 13 9 1 10 9 2 0 2 1 10 9 2
49 13 1 10 9 15 13 10 9 2 13 1 10 2 9 2 0 2 0 7 1 0 9 2 10 9 13 1 9 1 9 2 13 10 9 2 13 10 9 1 9 2 13 10 9 2 13 10 9 2
11 10 10 9 13 1 10 3 0 15 13 2
9 9 0 0 3 3 1 9 1 12
16 10 9 0 0 3 13 13 15 10 9 2 3 13 10 11 2
40 12 9 1 10 3 0 9 1 13 1 10 9 1 10 11 7 10 11 2 1 10 9 1 10 0 9 2 13 13 0 9 7 13 1 10 9 1 10 9 2
27 1 10 11 13 15 13 1 10 9 13 1 10 9 2 15 13 13 15 9 1 10 3 9 1 10 9 2
14 3 13 10 9 2 1 10 0 9 0 1 10 9 2
9 1 11 2 10 9 3 13 0 2
20 1 12 7 12 2 10 9 1 10 9 1 9 13 1 12 9 1 12 9 2
24 13 15 13 16 10 9 1 10 9 0 15 2 1 13 9 2 13 13 1 9 1 12 9 2
29 2 11 2 2 9 15 13 13 1 10 0 9 2 13 13 1 10 9 11 7 11 7 1 10 9 11 7 11 2
22 13 1 10 11 2 10 9 13 13 10 2 9 0 7 0 1 10 9 1 11 2 2
30 1 10 9 1 11 7 10 9 11 2 13 3 10 9 13 1 10 9 15 13 10 9 1 10 9 1 10 9 11 2
23 1 10 9 2 10 9 13 0 2 7 1 10 9 10 0 9 1 10 9 13 3 0 2
14 3 16 10 9 13 1 13 10 9 1 10 12 9 2
65 10 9 0 1 10 9 1 10 9 11 2 11 2 13 10 9 1 10 9 0 13 1 10 11 1 13 10 9 1 10 9 2 1 10 9 1 13 10 9 1 10 12 9 13 1 10 9 0 3 0 1 10 9 2 12 3 9 0 7 10 0 3 9 0 2
26 11 13 3 10 9 1 10 9 0 11 2 11 7 10 9 1 10 11 11 2 10 9 1 10 9 2
16 10 9 13 13 1 10 9 2 15 3 13 13 1 10 9 2
46 15 1 15 13 1 10 9 1 10 0 9 2 3 2 3 11 7 10 11 13 3 10 9 2 9 2 2 16 15 1 10 2 9 2 15 1 10 9 13 1 13 15 10 9 0 2
44 11 13 10 0 15 13 1 13 0 7 13 2 13 1 10 10 9 9 1 9 0 2 0 1 10 9 1 10 9 0 2 1 10 0 9 0 1 10 2 9 2 1 11 2
51 16 15 13 3 3 13 1 2 11 2 2 10 9 1 10 10 9 1 9 7 1 10 11 2 15 3 13 1 10 9 2 3 13 0 16 1 10 0 0 9 13 1 10 0 9 10 9 13 1 11 2
54 10 9 0 13 2 11 2 2 10 0 2 9 2 13 1 10 0 9 1 9 7 15 3 13 13 1 10 9 1 10 9 13 0 1 9 1 9 0 2 15 3 15 13 1 13 1 10 2 0 2 11 7 11 2
16 1 9 2 10 9 13 10 0 9 1 10 9 1 10 9 2
11 3 2 13 15 10 9 1 9 7 9 2
29 11 2 1 10 10 9 1 10 9 2 13 15 10 9 7 11 13 13 1 11 1 15 15 13 3 10 9 13 2
62 7 11 13 15 16 15 13 1 13 2 3 3 15 13 13 9 10 3 3 13 10 10 9 2 1 15 15 11 2 2 16 15 1 10 9 13 1 10 9 2 2 15 13 16 3 13 13 10 12 9 1 11 7 15 16 13 10 9 1 15 12 2
38 7 13 3 1 10 9 1 11 16 13 13 3 2 7 15 3 2 3 9 7 9 3 3 13 10 9 2 10 9 7 10 9 0 2 0 7 0 2
36 3 2 13 10 9 16 9 7 9 2 1 10 0 9 1 10 9 2 3 3 13 3 1 10 0 9 2 10 9 0 1 9 3 1 9 2
9 2 7 15 13 1 13 10 9 2
59 10 9 13 3 9 15 13 10 9 1 10 9 0 1 10 9 1 10 9 2 10 9 1 10 9 1 10 11 2 7 13 1 10 9 1 9 1 10 9 1 10 9 2 13 2 3 2 10 9 1 10 9 0 1 10 0 9 11 2
55 1 10 9 3 13 2 13 15 13 1 10 11 16 13 10 9 1 10 11 2 13 10 9 1 13 10 9 1 10 9 7 10 9 0 2 13 1 0 10 9 1 10 11 7 13 9 1 9 1 9 0 1 10 9 2
63 7 3 13 3 0 16 10 9 11 15 2 3 9 2 13 10 9 1 10 9 15 15 13 2 13 9 1 13 10 9 1 10 15 13 1 13 1 10 9 2 1 13 10 9 1 13 10 9 3 0 16 11 13 9 1 13 15 1 2 10 9 11 2
25 2 7 2 16 10 9 11 13 13 9 1 10 9 2 13 16 2 3 2 13 1 10 10 9 2
33 10 9 13 4 13 1 10 9 1 10 9 2 11 2 15 3 13 1 10 9 1 9 2 3 1 10 9 1 10 2 9 2 2
17 2 10 11 3 3 13 10 9 2 16 13 1 13 10 10 9 2
29 7 2 3 3 3 13 0 16 13 4 13 10 0 9 2 1 15 3 15 13 13 1 10 9 11 1 11 2 2
50 11 13 2 3 2 16 11 13 12 1 10 9 15 13 1 4 13 1 10 9 2 13 15 4 13 10 9 1 10 9 1 9 2 1 10 0 9 1 12 1 10 9 1 10 11 2 1 10 11 2
32 1 10 9 2 10 9 13 4 13 1 9 1 12 7 2 16 10 9 13 1 11 2 15 13 2 10 0 9 2 1 9 2
27 2 1 12 3 13 13 10 9 1 10 0 11 2 11 2 7 3 3 13 0 15 1 10 11 1 12 2
32 7 2 13 3 0 13 10 9 1 9 0 15 13 13 10 9 1 10 9 2 15 13 13 1 9 0 1 10 9 0 2 2
20 11 2 7 13 3 9 3 2 13 12 12 2 1 10 9 2 10 11 2 2
32 13 10 9 3 13 1 10 9 1 10 9 15 13 10 10 9 2 7 13 1 10 0 2 16 13 10 9 16 13 1 15 2
18 13 0 16 13 1 13 10 9 1 10 9 13 3 1 10 9 0 2
14 9 2 7 15 13 10 10 9 1 10 9 0 0 2
14 15 3 13 16 13 1 10 9 1 9 1 10 9 2
34 10 11 13 3 13 13 10 9 1 10 9 1 3 12 9 0 1 10 11 2 7 13 13 13 10 9 1 13 12 13 1 10 11 2
51 1 10 9 1 11 2 10 9 3 13 13 2 10 9 0 1 10 11 13 16 15 13 10 9 1 12 9 1 9 11 2 1 10 9 1 12 9 2 1 13 13 1 11 2 1 10 9 1 10 11 2
48 10 11 2 0 1 10 9 1 10 11 7 1 11 2 3 15 13 13 2 1 10 9 1 10 9 2 1 13 1 10 10 9 10 9 1 12 9 2 1 10 9 13 1 12 9 1 9 2
42 1 10 11 2 11 2 9 1 10 9 1 11 2 0 1 10 9 0 2 13 10 9 1 10 9 1 12 9 0 2 1 13 10 9 1 11 15 13 1 10 11 2
27 1 15 2 15 13 13 4 1 10 9 7 4 1 9 2 3 1 10 9 1 10 9 13 1 10 11 2
6 2 11 2 1 10 11
6 11 3 3 1 10 9
43 10 11 13 9 1 10 10 9 10 11 2 1 12 2 13 1 13 2 1 12 2 10 9 1 10 11 1 10 11 2 11 2 2 15 15 13 1 10 0 1 12 9 2
3 11 1 11
9 11 1 10 9 1 10 2 9 2
18 10 11 13 9 7 9 2 7 2 3 13 0 1 13 2 10 11 2
19 10 9 13 13 3 2 1 11 2 1 10 9 1 10 11 2 11 2 2
47 11 13 2 1 10 11 2 10 9 1 10 9 15 13 2 10 9 3 0 1 10 9 2 2 1 13 13 1 10 2 9 2 1 10 9 2 13 1 10 2 9 1 10 10 9 2 2
31 10 9 1 9 0 13 15 1 10 9 1 10 9 3 3 1 9 2 3 1 9 1 10 9 1 10 9 1 10 9 2
74 3 2 11 2 15 13 10 9 2 0 2 2 1 10 9 15 13 1 10 9 7 13 1 10 9 2 0 2 0 2 1 10 9 7 1 10 9 2 13 3 10 9 0 2 7 13 0 1 10 9 2 2 1 10 9 0 7 0 2 1 10 9 0 2 10 9 1 10 9 7 1 10 9 2
17 1 10 9 1 9 13 2 10 0 9 1 0 9 13 10 9 2
32 2 11 2 2 13 10 9 1 9 1 10 9 2 15 13 1 15 0 2 0 7 0 2 0 7 0 2 9 1 10 9 2
16 11 2 9 15 13 10 10 9 1 10 9 1 10 9 0 2
54 3 13 9 1 9 2 7 1 10 10 9 2 15 3 13 1 3 1 13 10 9 1 10 9 1 12 1 10 9 3 0 2 7 0 2 0 1 10 9 2 10 2 9 2 2 7 10 9 3 2 9 0 2 2
64 11 13 10 9 13 1 9 3 0 2 15 13 10 9 1 15 9 1 10 3 0 9 1 10 9 2 10 9 1 10 9 1 9 1 10 9 0 2 10 9 1 10 9 2 2 3 13 3 1 13 3 0 10 9 0 2 3 0 2 15 3 15 13 2
42 10 9 13 13 1 9 2 9 0 2 2 1 9 1 9 2 13 15 1 15 12 12 9 0 2 0 2 7 1 16 10 9 15 13 1 10 9 0 1 10 9 2
15 13 10 9 1 10 9 2 1 10 9 7 1 10 9 2
33 1 12 2 10 9 1 10 11 13 16 10 9 13 9 0 1 10 12 9 1 9 7 13 13 10 9 1 9 2 13 1 12 2
51 1 10 9 1 9 1 9 2 10 11 13 3 13 1 12 9 1 9 10 9 1 10 9 1 9 2 13 15 1 12 9 2 1 10 12 9 15 15 13 1 9 2 7 13 12 0 13 1 10 9 2
36 11 13 3 16 10 9 1 12 2 12 13 13 1 10 9 0 1 13 13 1 15 2 3 2 1 10 9 1 10 9 2 9 1 10 0 2
22 10 11 13 1 13 0 9 1 10 9 0 7 10 9 1 9 13 13 1 0 9 2
26 16 10 11 3 13 13 10 0 9 2 13 3 13 16 10 11 13 12 1 10 0 9 1 10 9 2
6 11 3 13 1 10 9
39 1 10 9 1 13 10 11 2 10 11 13 3 13 13 1 10 9 1 10 9 1 10 10 12 9 0 2 11 7 11 2 15 15 13 1 13 10 11 2
57 10 9 2 15 13 10 9 0 1 10 9 1 11 2 13 3 1 10 9 1 11 2 3 12 9 3 1 10 10 9 13 4 13 1 10 9 1 10 9 0 1 10 9 0 2 13 3 3 13 1 10 9 1 10 9 9 2
34 1 10 9 1 11 7 11 2 10 9 0 1 10 11 13 1 10 10 9 10 9 2 1 9 1 10 0 11 2 15 15 13 13 2
10 15 13 10 9 2 15 13 10 9 2
5 15 3 13 13 2
7 15 13 10 2 9 2 2
26 13 10 9 2 10 9 2 15 9 2 7 10 9 2 1 13 12 9 11 1 11 2 1 10 9 2
79 3 13 15 2 7 3 15 13 3 1 13 16 1 10 9 3 13 3 15 2 13 10 0 9 2 7 2 3 1 10 9 3 13 13 7 10 9 7 10 9 2 13 1 10 0 9 1 13 10 9 10 15 13 1 10 9 1 10 9 0 2 13 15 3 10 9 2 13 3 15 2 1 15 3 13 1 4 13 2
5 10 9 1 11 2
3 10 9 2
16 10 9 13 2 11 2 2 7 13 13 1 10 11 1 12 2
26 3 1 2 11 2 2 1 2 11 2 2 1 2 11 2 2 1 2 11 2 2 1 2 11 2 2
13 3 1 2 11 2 2 7 3 3 1 10 9 2
21 2 11 2 13 3 3 0 7 0 3 10 9 3 13 0 7 13 1 10 9 2
11 10 9 1 10 9 13 10 9 1 9 2
44 10 9 13 0 2 0 7 0 3 1 10 9 1 11 2 16 10 0 13 9 15 15 13 3 1 10 9 0 1 3 3 13 13 7 3 15 15 13 0 1 3 13 13 2
45 11 1 10 9 13 9 1 10 2 11 2 2 7 13 9 1 10 11 1 13 10 9 1 2 11 2 2 13 1 4 13 15 15 1 0 15 13 1 9 1 13 3 12 9 2
32 13 16 13 16 2 10 9 13 10 9 1 0 15 13 1 10 9 1 10 9 15 15 13 13 9 0 0 1 10 9 2 2
77 10 9 3 13 2 7 10 9 13 15 9 0 2 7 0 1 10 10 9 2 10 9 3 1 9 13 15 2 10 0 2 10 9 2 10 9 2 10 9 1 10 0 2 13 10 9 0 15 3 13 3 13 7 13 2 7 11 15 13 9 2 10 9 13 2 10 9 7 10 9 2 7 3 13 10 9 2
6 11 13 1 10 9 2
18 3 1 10 9 2 13 1 12 9 1 9 2 13 12 9 1 9 2
12 13 15 1 10 9 15 3 13 9 1 15 2
17 3 15 13 9 1 10 9 1 10 9 3 10 9 13 13 9 2
15 10 9 3 13 1 10 9 13 2 11 2 2 1 11 2
10 3 9 3 3 3 11 13 10 9 2
50 3 1 10 9 3 1 10 9 7 10 11 2 11 2 3 15 13 10 9 0 0 1 10 0 9 1 10 9 13 1 10 9 1 10 9 7 15 13 10 9 1 10 9 0 1 10 9 1 9 2
19 13 15 13 10 9 1 10 11 1 13 1 10 9 10 9 0 7 0 2
25 3 13 10 9 1 13 10 9 3 0 3 15 1 10 0 9 1 10 9 1 15 3 13 9 2
25 7 1 10 9 0 2 1 15 10 9 13 0 2 7 15 10 9 13 2 13 10 9 1 9 2
50 2 10 9 1 10 11 2 10 9 2 13 3 13 1 10 11 2 1 11 2 10 9 0 13 2 11 2 2 7 2 13 1 10 9 3 0 7 1 10 9 3 0 1 10 9 2 2 11 2 2
85 16 1 10 0 9 1 10 9 1 12 10 9 1 10 9 1 10 12 2 0 9 2 13 3 13 2 1 10 0 9 1 10 10 9 2 9 13 1 15 0 12 1 15 10 11 13 10 11 1 10 9 1 12 1 9 1 12 2 1 11 2 10 2 9 2 13 13 9 1 10 3 0 2 9 2 1 10 9 1 10 11 7 1 11 2
35 10 0 9 1 10 0 9 2 0 2 13 1 10 9 1 10 11 2 1 10 10 12 0 9 1 11 2 13 13 3 10 2 9 2 2
30 9 2 2 7 3 2 3 3 1 10 9 13 1 13 1 10 9 2 7 1 10 9 0 2 10 9 1 10 9 2
23 9 2 2 3 13 7 13 9 1 10 9 0 15 13 16 13 1 10 9 1 10 9 2
23 7 2 13 9 2 13 3 13 1 16 10 11 13 13 7 2 3 2 13 13 9 0 2
14 13 15 2 3 13 7 10 0 7 10 0 2 13 2
42 9 13 2 10 9 11 2 9 2 9 0 7 0 9 1 10 11 1 10 11 1 9 1 12 1 11 2 13 10 9 1 15 15 13 10 2 11 2 1 10 11 2
18 1 9 1 10 9 1 9 1 10 9 0 2 13 10 9 7 9 2
18 3 1 10 9 1 10 9 2 13 16 10 9 13 4 1 13 9 2
13 1 3 3 13 0 1 0 9 1 10 10 9 2
12 11 2 1 3 9 13 10 0 11 1 9 2
37 3 13 3 10 9 1 10 9 1 13 0 9 0 7 1 9 2 11 13 16 2 1 15 13 10 9 2 2 13 1 13 16 13 3 7 3 2
15 10 9 3 13 3 3 9 10 9 0 2 7 10 9 2
24 1 10 9 2 13 16 10 2 9 7 10 9 1 10 9 2 13 10 0 9 1 10 9 2
32 1 10 10 9 2 10 10 9 3 13 10 9 1 16 10 9 1 10 11 13 1 10 9 0 1 10 9 1 10 9 0 2
23 3 2 10 0 9 0 2 3 1 10 9 2 13 3 1 13 13 1 10 9 1 9 2
42 1 10 9 2 13 16 10 2 9 13 0 1 13 10 9 1 10 9 1 9 2 1 9 1 10 9 1 9 13 2 2 13 3 13 10 9 1 1 13 10 9 2
24 1 10 11 2 3 13 10 9 1 10 9 7 10 9 2 13 10 9 1 10 9 1 9 2
32 11 13 10 9 1 10 11 1 13 10 9 1 9 1 11 2 15 3 13 1 13 2 7 13 10 9 1 10 9 1 9 2
6 10 9 0 0 2 0
23 11 13 15 3 13 1 10 9 15 13 4 15 13 3 1 10 11 2 7 13 10 9 2
26 3 13 1 15 2 1 10 9 1 10 9 15 13 10 9 1 9 13 2 9 0 1 10 10 9 2
17 2 1 9 2 11 2 3 13 1 10 10 9 15 13 13 2 2
11 13 10 0 9 2 13 3 15 13 2 2
5 2 11 2 2 11
21 12 9 1 13 10 9 1 11 1 10 9 11 2 10 9 15 15 13 10 9 2
34 12 1 10 3 0 9 1 10 0 9 2 11 13 10 9 1 9 7 10 9 1 13 7 15 13 1 10 9 15 13 9 1 11 2
43 13 1 10 9 1 10 0 11 2 1 15 15 13 10 0 9 0 2 3 13 13 3 2 11 13 13 15 1 10 9 15 15 13 10 9 1 13 7 15 13 13 15 2
26 13 1 10 9 1 13 0 7 0 1 10 9 2 10 9 13 9 2 13 9 2 13 1 10 9 2
72 1 10 9 1 15 11 13 10 9 7 10 9 1 13 10 9 2 1 15 15 13 13 3 2 1 15 13 2 1 9 0 2 10 9 2 11 2 2 1 10 0 9 15 15 13 10 9 2 1 10 9 7 9 1 10 9 0 13 1 11 2 2 10 0 9 15 13 1 10 9 0 2
7 13 15 3 1 10 9 2
10 11 2 9 2 13 1 10 9 0 2
35 7 11 13 10 10 9 1 15 1 10 15 15 13 1 10 9 1 11 2 13 1 12 9 1 10 9 1 10 9 2 13 13 3 12 2
7 13 1 10 2 9 2 2
2 13 2
7 2 10 9 13 9 2 2
9 13 10 9 3 0 1 10 9 2
58 1 9 1 10 2 15 13 10 9 1 13 1 1 10 9 15 1 10 9 3 0 1 10 9 1 9 2 13 15 1 13 2 3 2 10 9 1 13 9 1 9 1 10 9 2 1 10 9 7 3 10 9 1 10 9 1 9 2
29 1 10 10 9 2 11 13 12 9 0 9 2 11 7 11 2 15 13 1 15 15 13 13 10 9 0 1 11 2
36 2 3 10 11 13 0 1 13 3 16 13 0 13 1 10 9 0 2 2 10 9 13 1 16 2 15 13 9 1 13 10 0 9 0 2 2
16 11 13 10 10 9 1 10 9 1 10 9 1 10 9 13 2
24 2 10 10 9 2 13 7 0 2 1 13 4 1 13 10 11 2 3 15 13 13 0 2 2
27 7 13 1 10 2 9 7 1 10 9 2 1 10 11 3 10 9 0 1 13 9 1 10 10 0 9 2
66 11 13 1 10 9 1 9 1 10 9 1 2 11 2 2 10 9 15 13 1 10 9 1 10 9 1 11 2 9 1 12 2 2 1 15 13 13 10 9 1 10 9 3 0 2 1 9 0 7 0 2 7 3 0 2 1 10 9 1 10 12 9 1 10 11 2
46 2 10 0 9 1 10 9 13 13 3 10 9 0 1 10 10 9 0 1 13 2 1 10 9 0 1 10 10 9 2 9 1 9 2 9 0 7 9 1 0 2 2 13 10 9 2
16 2 3 10 0 11 3 13 1 4 13 3 12 1 10 11 2
26 7 13 13 15 3 3 16 10 10 9 2 7 2 13 13 7 13 2 10 10 9 13 3 13 2 2
15 9 0 1 10 9 11 1 11 2 12 0 7 12 13 2
12 13 10 9 1 10 9 1 10 10 9 11 2
1 9
19 11 7 11 13 15 1 11 2 13 16 10 11 13 13 1 9 7 9 2
14 9 1 10 9 13 3 7 11 13 1 9 1 10 9
10 9 3 13 10 9 1 13 1 10 9
9 11 13 10 0 9 1 10 9 2
15 13 9 1 13 15 9 1 13 1 9 2 7 13 0 2
34 1 10 0 9 3 13 13 15 7 13 2 11 2 2 1 10 11 2 1 11 2 7 2 11 2 2 1 10 11 2 1 10 11 2
3 7 13 2
21 10 9 13 15 3 1 10 9 15 13 2 1 11 2 1 10 9 1 10 9 2
17 1 10 9 1 15 13 13 10 9 1 9 1 10 9 3 0 2
8 9 1 10 11 1 11 13 9
5 10 9 1 10 9
16 10 9 1 10 11 1 11 3 13 13 10 9 1 10 9 2
9 9 1 9 2 13 13 10 9 2
23 3 2 3 2 15 13 1 10 9 15 10 9 13 13 10 9 7 15 10 9 3 13 2
9 3 2 13 16 13 13 10 9 2
5 11 13 13 9 0
33 10 11 13 1 10 9 1 10 11 16 13 13 10 9 0 13 1 10 9 1 9 2 13 9 0 0 7 0 13 1 10 11 2
52 10 9 13 16 10 9 3 2 10 9 2 12 9 3 0 16 10 9 2 3 13 0 1 10 9 7 13 13 10 9 1 10 9 0 2 15 10 9 1 10 11 13 1 13 2 16 10 9 3 13 13 2
9 10 11 7 10 11 13 10 11 2
30 10 9 1 9 13 13 1 10 11 7 1 10 11 3 1 10 9 1 9 13 13 16 10 9 13 9 1 10 9 2
43 10 11 2 10 0 9 1 10 11 15 13 10 9 2 13 3 13 10 9 1 10 11 13 1 10 9 1 16 10 9 13 2 1 10 9 2 1 10 9 7 9 0 2
37 7 10 9 1 10 11 1 10 9 0 2 13 1 9 1 10 12 9 2 13 10 9 3 1 13 10 9 0 1 10 0 1 10 9 1 9 2
22 11 2 9 0 7 9 13 2 13 10 9 7 13 11 2 9 1 9 2 7 11 2
19 11 3 15 13 3 1 9 2 3 13 13 1 15 15 15 13 1 13 2
12 13 15 1 10 9 2 15 13 1 0 9 2
21 2 13 10 9 3 2 2 13 15 0 2 7 3 15 13 1 13 1 10 9 2
17 3 3 11 15 13 1 10 9 2 15 13 1 16 13 3 9 2
10 10 9 2 1 9 13 2 13 15 2
16 7 3 11 13 10 0 9 1 10 9 3 1 10 9 13 2
8 2 15 13 15 13 13 2 2
8 11 2 12 1 9 1 12 2
29 13 9 9 7 11 13 10 9 3 1 10 9 1 10 11 2 13 1 10 11 7 10 9 0 9 1 10 11 2
34 9 1 10 11 13 15 1 9 0 2 13 9 1 10 9 2 15 15 13 13 2 3 10 9 1 9 2 3 12 9 1 9 2 2
23 10 9 13 9 3 10 9 1 10 9 0 1 11 7 10 9 1 10 11 2 1 10 2
23 1 10 9 11 2 13 15 1 10 9 2 0 1 10 9 0 7 0 1 10 9 2 2
36 1 9 13 1 10 0 9 1 10 9 2 10 11 13 2 1 10 9 0 1 10 9 13 2 12 9 2 3 15 12 16 1 10 9 0 2
24 10 0 1 10 9 2 3 15 1 10 9 2 13 16 2 10 9 13 3 1 10 9 2 2
14 1 15 10 9 13 13 10 11 2 1 10 9 0 2
16 2 16 11 3 13 1 10 9 2 10 9 13 1 11 2 2
13 9 1 10 11 15 13 1 10 9 1 10 9 2
16 10 9 3 1 13 1 10 11 15 13 10 9 1 10 11 2
9 9 0 1 10 11 3 13 9 0
7 11 13 1 10 11 1 9
63 10 11 2 11 2 13 3 2 1 13 2 3 2 0 2 10 9 0 13 1 10 9 11 2 1 10 9 1 10 9 1 10 9 0 1 11 1 10 9 0 11 2 13 16 13 13 10 10 9 1 13 10 9 1 10 11 0 1 10 9 1 9 2
48 10 9 1 13 9 2 13 1 10 9 1 9 1 10 9 1 10 9 1 9 1 10 9 1 9 1 10 9 0 1 11 2 13 1 4 13 1 9 15 13 9 1 10 0 9 1 9 2
44 3 12 9 1 9 1 9 2 1 9 7 1 9 0 2 13 13 1 10 9 1 12 1 12 1 9 1 10 9 1 9 1 10 11 2 11 2 2 1 10 11 2 11 2
16 15 13 13 16 10 9 13 10 9 1 13 10 9 1 9 2
18 13 3 10 9 0 1 10 9 15 13 13 2 13 15 13 1 9 2
7 1 10 9 2 10 9 2
25 3 2 1 10 11 3 13 0 9 1 10 9 1 10 9 16 13 9 1 10 0 9 1 11 2
30 16 10 9 0 2 3 2 13 1 10 9 1 12 1 12 9 2 13 10 15 1 10 9 7 10 9 13 10 9 2
31 13 15 10 9 7 3 13 13 10 9 1 10 9 1 10 11 7 13 10 9 0 1 15 10 11 13 9 1 10 11 2
33 3 2 10 11 2 11 2 13 3 10 11 1 10 3 9 1 10 9 1 10 9 11 2 1 10 9 1 10 9 1 15 13 2
47 10 9 1 11 13 10 9 1 12 9 1 13 2 13 10 11 1 10 10 0 9 13 10 9 2 15 2 16 13 0 1 10 11 2 15 13 13 10 9 1 10 12 7 12 12 9 2
8 1 12 7 12 9 2 3 2
3 11 13 11
30 10 11 13 1 10 11 2 11 2 10 9 11 2 2 9 2 1 9 0 2 7 11 2 2 9 2 1 9 0 2
29 7 10 0 0 9 1 11 13 1 11 2 1 10 9 0 2 1 3 0 1 10 11 7 3 9 1 10 11 2
33 1 10 9 0 1 10 9 1 10 9 2 11 2 13 7 13 10 0 9 15 15 13 1 13 10 9 1 11 1 12 2 11 2
27 11 13 1 10 9 1 10 9 2 13 1 9 3 13 1 9 1 10 9 0 2 13 3 9 7 9 2
7 7 13 3 15 15 13 2
23 1 10 9 13 9 2 13 9 0 2 1 16 12 9 13 1 10 9 1 10 9 0 2
10 10 11 13 15 2 13 15 1 11 2
7 7 11 13 1 13 15 2
49 10 9 0 1 10 11 2 11 2 13 13 2 1 10 9 13 2 13 0 1 13 10 9 0 1 13 12 9 0 2 12 9 7 12 9 2 1 13 1 13 1 10 0 9 2 1 10 11 2
38 11 13 16 10 9 0 13 15 13 2 1 9 2 1 16 10 11 13 10 10 2 9 2 1 9 7 9 2 3 1 10 9 1 10 12 9 0 2
23 10 9 0 13 9 1 10 9 1 12 9 2 10 9 7 9 0 1 13 10 9 0 2
4 10 9 1 9
49 3 1 10 9 13 12 9 2 10 9 0 1 2 3 2 13 10 9 1 9 1 10 9 7 2 1 0 9 2 10 9 1 13 10 10 9 1 9 0 1 10 12 9 1 10 9 0 0 2
34 10 9 13 13 13 3 10 9 1 10 9 1 13 10 10 9 2 2 3 13 1 10 9 7 10 2 0 9 2 2 2 13 11 2
4 9 11 1 11
6 11 1 9 1 10 9
34 10 9 11 2 11 13 1 10 9 1 10 0 11 1 11 2 9 0 1 10 2 9 2 1 9 2 1 10 9 1 10 0 9 2
48 10 9 1 9 1 10 0 2 11 2 11 2 1 11 2 13 1 10 9 1 10 11 10 9 9 1 9 1 13 10 9 1 10 9 2 15 15 13 1 0 9 1 10 9 1 10 9 2
12 10 9 13 3 13 1 10 11 2 1 11 2
9 3 2 10 9 10 0 13 15 2
16 11 13 15 2 13 15 7 13 15 2 1 9 1 10 9 2
20 10 11 2 1 10 11 13 10 9 15 15 13 13 1 10 9 1 10 11 2
10 1 11 2 10 9 3 13 3 13 2
20 1 10 10 9 1 11 2 3 2 11 2 13 10 9 7 13 1 10 11 2
30 15 13 0 16 2 1 10 9 2 10 9 13 10 9 0 7 0 15 2 1 10 9 2 1 10 11 13 4 13 2
9 9 0 13 9 1 9 1 10 9
53 10 9 0 1 10 11 7 1 10 11 13 3 1 10 11 9 0 13 10 9 0 1 12 9 1 9 1 10 9 7 10 9 1 9 1 10 9 1 9 1 10 9 13 1 10 9 2 13 10 9 0 11 2
32 10 12 9 13 13 9 1 10 9 0 1 10 0 9 1 15 12 2 1 12 1 9 1 11 2 7 13 15 10 9 0 2
45 10 9 13 0 9 1 9 2 12 1 10 12 9 1 9 0 2 10 9 2 12 9 13 1 10 9 1 10 9 1 10 9 7 10 9 3 2 11 2 2 9 1 10 9 2
16 10 9 7 10 9 0 1 10 9 13 3 13 1 10 9 2
21 10 9 2 13 11 2 13 13 1 10 9 2 7 13 1 9 1 9 1 9 2
35 10 9 13 13 3 13 1 9 7 13 1 10 9 1 9 7 13 1 9 1 9 1 10 9 2 13 10 9 13 1 10 11 7 11 2
30 1 10 9 1 9 13 1 10 9 13 4 13 2 11 13 16 3 13 13 10 2 9 1 10 9 1 10 9 2 2
35 1 10 11 13 13 10 9 1 10 9 2 16 1 9 1 9 3 13 2 16 3 13 4 13 10 0 9 1 9 0 13 1 10 9 2
11 10 9 13 0 7 13 1 10 12 9 2
70 10 9 9 11 2 3 2 1 3 15 13 1 10 9 1 13 10 12 9 2 3 1 13 16 13 2 0 9 0 2 1 10 9 1 10 9 1 10 9 2 15 3 15 13 2 1 10 9 1 9 0 2 15 3 13 15 1 15 15 10 9 1 9 7 10 9 0 13 2 2
8 9 15 15 13 10 9 0 2
31 2 13 16 13 0 15 12 9 1 13 15 3 13 1 15 15 12 13 13 16 10 15 3 13 9 7 3 13 15 2 2
44 10 9 1 10 9 13 4 1 4 13 13 2 3 2 0 1 2 13 9 0 2 2 16 3 2 1 10 9 3 10 9 13 4 13 1 10 9 3 10 9 15 13 2 2
44 11 2 13 13 1 10 9 1 12 9 2 1 13 1 10 9 1 10 0 9 2 9 1 9 1 10 9 0 1 12 2 12 2 9 1 10 9 1 11 2 0 9 2 2
12 1 10 11 13 13 2 3 2 3 12 9 2
7 10 9 13 10 0 9 2
8 15 13 13 3 3 10 9 2
26 10 9 1 9 0 1 12 9 2 13 1 0 2 13 13 1 9 1 12 1 9 2 3 1 12 2
27 16 10 9 1 9 1 0 13 10 9 1 9 0 2 0 13 16 15 13 1 10 9 1 10 10 9 2
9 3 0 3 13 13 10 9 0 2
7 2 11 2 2 1 11 2
15 15 13 2 1 15 2 10 0 9 0 1 10 0 9 2
9 11 2 3 3 11 2 13 1 9
5 9 1 10 0 9
10 2 12 9 0 15 13 9 0 2 2
32 3 15 13 10 11 2 14 11 2 15 1 3 12 9 1 9 1 10 9 13 1 9 1 10 0 9 7 10 9 1 9 2
16 1 10 9 2 3 2 13 3 2 11 2 2 10 9 0 2
1 9
53 2 11 2 2 10 9 1 9 1 9 1 11 2 13 1 12 1 11 2 11 7 11 2 1 10 9 1 9 1 10 9 2 11 2 2 1 11 2 13 4 13 1 12 1 9 1 10 9 11 1 10 11 2
45 2 11 2 13 10 9 1 10 9 2 9 1 11 2 15 13 1 10 9 13 1 10 9 7 15 13 4 13 2 1 10 9 2 1 10 11 2 11 2 12 2 2 1 11 2
77 10 9 13 3 13 2 13 1 10 2 11 2 13 11 7 11 2 9 2 12 7 12 9 2 3 2 13 1 12 1 12 9 1 9 2 11 2 9 2 12 9 2 13 1 12 9 2 11 2 9 2 12 9 2 13 1 12 9 2 7 11 2 12 9 2 0 9 1 10 9 11 2 13 1 12 9 2
19 3 13 9 2 3 15 13 1 10 9 1 9 2 3 1 10 9 0 2
19 1 10 9 1 10 11 2 10 9 13 0 1 10 9 0 3 13 13 2
12 7 3 10 0 9 1 10 11 15 13 13 2
18 13 15 3 1 3 13 4 13 2 13 1 10 9 13 1 10 11 2
23 10 0 9 2 1 3 13 9 2 13 1 3 13 10 9 7 13 15 3 15 15 13 2
18 3 2 13 16 13 9 1 9 1 9 2 3 1 9 0 1 10 2
5 0 9 1 10 11
29 10 9 13 1 10 9 1 9 2 15 1 10 9 3 13 3 13 2 13 1 13 9 2 15 3 3 13 13 2
15 15 10 9 13 13 3 13 13 3 0 15 13 1 13 2
14 13 13 10 9 7 13 10 9 1 9 1 10 9 2
16 16 3 15 13 3 13 16 13 9 1 13 1 10 9 0 2
9 15 3 3 15 13 3 15 13 2
7 11 13 9 0 1 10 11
3 11 1 11
43 10 2 11 2 15 11 13 1 10 11 13 15 1 10 9 0 1 9 7 9 1 9 3 13 9 2 10 11 2 10 0 9 2 1 11 2 7 10 9 0 1 9 2
8 10 9 2 15 2 13 3 2
25 10 9 0 11 13 15 1 10 9 0 7 13 3 1 10 9 15 15 0 13 2 10 9 11 2
44 13 15 3 2 13 15 10 9 7 13 10 9 0 1 10 9 1 10 9 2 7 13 1 13 10 9 0 1 10 9 13 1 10 10 9 3 1 10 9 13 1 10 9 2
14 2 13 0 2 10 9 13 15 1 10 9 7 13 2
16 7 2 1 15 15 13 1 10 0 9 2 10 11 13 13 2
19 3 2 3 13 13 2 10 2 11 2 7 10 11 3 13 13 9 2 2
8 11 13 3 1 10 10 9 2
12 1 10 9 1 13 13 1 10 10 9 0 2
15 2 13 16 13 1 10 11 13 16 15 13 3 10 11 2
16 13 15 1 13 2 7 13 13 10 9 2 2 13 10 9 2
15 10 9 1 10 9 13 2 13 1 10 9 1 10 9 2
9 2 10 11 13 9 1 13 0 2
25 13 3 2 13 3 16 13 10 10 9 2 16 13 1 10 10 9 7 10 9 15 13 11 2 2
38 1 10 9 2 13 13 10 9 1 11 2 15 2 1 10 10 9 2 15 13 1 10 10 9 3 13 13 1 2 9 7 9 1 10 0 9 2 2
21 7 10 15 13 10 9 0 2 11 2 10 9 1 10 9 0 1 10 0 9 2
10 10 9 13 3 1 9 1 10 9 2
15 3 2 16 10 9 13 1 13 1 15 2 1 10 9 2
19 11 2 12 1 10 9 0 1 15 13 10 9 1 10 9 13 10 9 2
10 3 3 13 9 3 1 3 10 9 2
6 7 15 13 3 0 2
35 7 1 10 10 9 1 15 10 9 13 10 9 0 1 10 9 0 2 13 4 13 10 9 1 10 9 2 15 3 16 3 13 9 0 2
29 16 13 1 12 1 10 9 1 10 9 0 1 10 11 2 3 3 2 3 0 2 7 13 9 0 15 15 13 2
50 1 9 1 11 2 1 10 11 2 9 1 10 11 13 2 1 15 3 1 3 2 10 9 2 3 13 1 10 9 1 11 2 15 13 12 9 1 9 0 2 1 9 1 10 9 1 10 12 9 2
26 1 10 9 1 10 9 13 13 12 9 2 1 15 10 9 1 10 9 2 15 13 2 3 2 13 2
20 10 11 13 3 10 9 0 3 11 2 13 1 10 9 1 9 2 3 13 2
41 9 0 1 9 2 12 9 3 11 7 12 1 11 2 13 13 2 1 10 9 1 9 2 1 10 9 1 11 2 1 9 1 10 9 1 10 11 1 10 11 2
15 10 9 2 0 1 10 9 2 13 13 1 10 9 0 2
30 11 2 1 9 1 9 2 15 13 1 10 11 2 2 10 13 11 13 10 10 0 9 1 10 9 7 3 1 9 2
29 1 13 2 10 9 11 13 1 10 9 1 12 9 7 13 1 11 1 3 9 1 13 10 0 9 1 10 9 2
1 13
5 9 1 10 9 2
27 1 10 9 2 11 13 13 10 9 1 10 9 3 13 1 9 1 10 9 2 1 9 1 9 1 9 2
46 1 11 10 9 13 10 9 1 10 9 2 15 10 9 13 13 2 1 11 3 13 9 3 1 9 1 9 2 7 1 9 10 15 13 3 3 3 1 11 13 10 9 1 12 9 2
43 13 9 0 7 3 1 2 9 2 2 16 10 9 3 13 1 10 9 13 10 10 9 7 10 9 1 10 15 15 13 13 2 1 10 9 3 2 3 3 13 10 15 2
8 10 9 13 13 3 10 9 2
33 1 15 15 13 9 1 10 12 9 1 9 1 9 7 9 2 10 0 9 13 1 15 3 2 1 9 1 13 3 1 10 11 2
46 1 10 9 2 10 9 3 13 9 3 13 13 2 10 9 15 13 1 4 3 13 1 13 1 10 9 13 1 10 9 2 1 10 9 13 1 10 9 1 10 9 1 10 9 13 2
51 13 15 1 9 3 0 2 3 13 0 13 3 10 9 1 10 9 1 9 2 2 13 16 13 10 9 1 9 1 10 9 1 9 1 10 9 2 1 13 1 0 9 2 2 15 13 13 10 10 9 2
42 1 15 2 10 9 13 13 1 9 0 1 10 0 2 13 15 1 10 9 15 13 2 13 2 10 9 7 13 15 2 3 2 2 1 0 9 2 1 1 10 9 2
55 10 9 2 15 13 13 10 9 1 10 11 7 1 11 1 10 9 0 1 10 9 2 13 1 13 13 3 9 1 0 9 2 7 10 9 2 13 3 1 10 0 9 0 2 13 13 15 1 10 9 0 1 10 11 2
34 9 1 11 13 1 10 11 16 2 1 13 10 9 2 11 13 13 10 9 0 1 9 1 10 9 0 7 1 10 9 3 1 9 2
25 11 3 13 2 11 2 2 3 2 1 10 9 1 10 9 0 11 2 13 10 9 1 9 0 2
23 1 10 9 2 10 9 0 13 10 9 1 11 2 10 9 0 15 13 1 2 11 2 2
7 10 9 13 1 10 11 2
6 2 11 2 15 13 2
3 10 9 2
26 13 1 10 9 1 9 0 1 15 13 10 2 11 2 2 10 15 13 1 10 9 1 9 2 11 2
24 1 11 2 10 0 9 15 13 1 10 9 13 3 10 9 2 0 7 13 3 10 9 0 2
45 13 1 2 11 2 2 7 3 13 2 11 2 2 13 1 10 9 10 2 1 10 9 1 9 1 9 7 9 2 2 2 11 2 7 3 2 1 9 1 11 2 2 11 2 2
8 11 13 13 9 1 10 9 0
56 10 9 1 10 9 1 10 9 7 9 1 10 2 11 2 2 10 0 7 0 9 1 10 11 13 1 10 9 1 2 10 9 0 1 10 9 2 2 13 3 9 1 13 9 1 10 11 7 13 10 9 1 10 10 9 2
13 10 9 1 10 13 9 13 15 0 1 10 9 2
13 1 11 2 3 10 9 13 2 10 9 13 0 2
19 1 10 11 2 3 1 9 13 2 13 10 9 1 10 9 1 10 9 2
12 13 15 10 9 1 10 11 1 10 0 9 2
20 7 10 9 3 0 1 10 9 13 1 10 0 9 10 9 1 9 1 9 2
4 13 10 11 2
29 3 15 13 16 10 9 1 13 10 9 15 13 13 3 0 2 13 1 13 10 10 9 1 9 1 12 7 12 2
30 2 2 2 10 10 9 1 10 9 13 13 0 2 12 9 1 10 10 0 13 1 10 9 1 10 11 1 10 9 2
22 1 12 9 13 15 1 10 9 1 10 9 1 10 11 2 3 10 9 13 10 9 2
12 3 13 13 2 7 15 3 15 13 1 13 2
24 3 13 10 9 1 10 9 2 7 3 10 9 7 10 9 2 15 13 1 13 10 10 9 2
10 13 1 13 10 9 1 9 3 0 2
11 15 13 13 3 1 10 9 1 10 9 2
14 15 13 13 1 11 2 9 1 11 2 1 15 13 2
45 1 10 9 3 0 1 13 2 1 10 9 1 11 2 13 15 15 1 15 15 13 1 10 9 1 11 2 3 1 9 1 10 9 2 3 3 10 9 13 13 1 10 11 2 2
27 13 15 1 10 10 9 2 1 10 9 2 1 10 9 2 3 1 10 2 9 2 2 1 10 10 9 2
8 7 1 10 9 1 10 9 2
16 10 9 0 2 2 11 2 2 9 13 1 10 9 1 12 2
12 7 10 9 1 10 9 13 1 10 0 9 2
4 11 13 3 2
6 13 0 1 10 9 2
2 1 11
8 9 11 2 11 2 11 7 11
13 9 1 10 11 13 3 1 10 0 9 1 9 0
3 10 9 0
26 10 9 1 10 9 0 7 1 10 9 0 13 3 13 15 1 10 0 9 1 9 0 1 10 9 2
40 10 9 0 7 0 3 13 10 10 9 1 10 0 9 2 7 10 9 0 1 10 11 13 1 13 0 9 1 10 0 9 0 13 1 15 2 0 9 2 2
54 10 9 13 1 10 9 13 10 11 2 7 13 13 1 10 10 13 2 9 0 2 2 15 2 1 10 9 1 10 9 1 10 9 0 2 13 13 1 10 9 13 1 10 11 1 10 9 0 1 10 2 9 2 2
47 11 13 13 3 9 1 10 10 0 9 10 10 9 11 2 15 13 1 10 9 13 2 7 11 2 10 9 1 12 9 2 13 9 2 15 1 10 9 13 13 1 10 9 1 10 11 2
27 11 2 11 2 11 2 11 2 11 2 11 2 11 7 11 13 10 9 2 15 13 13 1 10 9 11 2
27 10 9 1 10 0 9 13 10 12 12 9 7 10 0 9 13 13 10 9 1 10 11 1 10 9 0 2
33 10 11 2 10 10 9 1 10 9 1 11 2 13 3 1 10 9 1 10 9 1 10 9 1 10 9 11 1 10 10 9 11 2
19 1 9 1 10 9 0 2 11 13 15 1 0 9 0 7 1 9 0 2
30 11 2 15 13 1 10 9 1 9 2 13 12 9 1 9 2 13 12 9 2 7 13 13 9 1 10 10 9 11 2
44 10 9 1 10 11 2 11 2 13 3 1 10 10 9 10 0 9 2 11 2 9 2 2 11 2 9 2 2 11 2 11 2 11 2 11 2 11 2 11 2 11 7 11 2
41 13 3 9 13 15 1 10 9 1 10 9 2 10 11 13 2 1 10 0 9 2 1 10 9 1 13 10 12 12 9 2 9 3 0 1 15 1 10 9 13 2
27 1 10 10 9 2 10 9 13 2 1 15 2 10 10 9 1 10 15 15 13 1 10 9 1 10 9 2
63 1 11 2 10 9 13 2 16 13 10 9 1 10 9 15 13 10 9 1 0 9 1 10 9 2 2 1 13 9 10 0 9 1 10 9 15 13 10 9 7 1 10 0 9 1 10 10 9 1 10 9 0 2 3 13 3 9 7 9 1 10 9 2
1 9
22 1 10 9 0 2 10 9 0 15 13 1 10 9 13 10 9 3 0 16 10 9 2
48 2 1 10 0 9 2 10 9 0 13 3 3 13 2 3 2 1 10 9 2 13 1 9 1 10 9 2 13 10 9 2 13 9 1 10 9 2 2 13 10 9 0 1 10 11 2 11 2
29 2 1 10 9 0 2 10 9 3 13 7 10 9 13 2 3 2 13 9 0 2 3 10 9 7 10 9 2 2
40 1 11 1 10 9 1 10 0 0 13 10 9 11 2 0 1 10 2 11 2 7 15 1 10 0 9 13 9 1 0 9 3 10 9 11 7 10 9 11 2
30 10 11 13 15 1 11 2 0 13 1 10 0 12 2 11 2 2 13 3 10 9 15 3 13 10 9 7 10 9 2
10 3 3 13 11 2 9 1 10 11 2
24 7 10 0 9 13 16 10 9 1 10 9 1 10 10 9 13 10 2 9 2 7 10 9 2
58 1 12 9 7 3 13 1 10 10 0 2 15 3 13 3 12 9 1 9 3 13 10 10 0 9 1 9 0 2 1 11 2 13 10 2 9 9 2 11 2 10 9 15 13 10 9 1 13 2 0 2 1 9 1 10 0 9 2
18 2 3 1 13 2 13 10 9 1 10 9 7 13 3 1 15 2 2
6 2 10 11 2 2 12
29 9 13 1 10 9 1 10 9 1 10 9 1 9 2 1 10 9 7 10 9 13 1 10 9 0 1 9 3 2
40 10 9 15 11 13 1 10 9 15 13 10 11 1 10 11 7 15 13 1 10 9 1 10 11 3 13 9 11 2 7 10 9 1 10 9 1 10 12 9 2
52 13 10 9 0 1 10 9 1 10 12 9 1 9 13 1 10 2 9 2 15 10 9 13 1 12 9 3 15 13 1 10 11 7 15 13 1 10 9 0 13 10 10 2 9 2 1 10 9 7 10 9 2
9 2 10 9 1 10 11 2 2 12
42 10 9 13 13 1 10 9 1 15 13 3 12 9 2 1 10 9 1 11 2 1 10 11 2 3 13 3 12 9 1 9 2 1 10 9 1 12 1 12 1 9 2
52 12 9 3 3 2 10 9 1 10 9 13 10 9 1 10 10 12 9 2 13 3 2 9 0 2 2 13 1 4 13 2 3 16 10 10 9 2 13 1 10 9 11 1 9 1 9 2 13 10 11 12 2
35 13 10 9 0 2 13 7 13 2 1 10 9 11 2 2 11 2 2 1 11 2 1 9 1 9 1 10 11 2 1 9 13 1 9 2
20 2 13 10 9 2 11 2 15 15 13 3 16 13 16 13 10 10 0 9 2
9 13 16 13 0 13 10 9 0 2
38 10 0 9 1 10 9 2 13 1 13 1 13 1 10 9 2 15 13 1 13 7 15 13 1 13 2 7 10 9 13 9 2 13 9 1 13 2 2
10 9 7 9 1 10 9 1 10 9 2
7 13 1 11 13 12 9 2
14 13 1 9 2 13 10 9 3 2 7 15 1 9 2
45 16 13 2 13 16 1 15 2 3 1 10 10 9 2 3 13 10 9 2 13 7 13 1 10 9 7 13 2 3 13 3 2 3 13 13 9 7 0 9 1 13 10 10 9 2
26 9 2 9 0 1 10 9 1 9 1 10 2 11 2 2 15 15 13 1 10 11 2 1 10 11 2
3 11 2 3
29 9 2 9 1 9 1 10 9 0 1 10 11 2 11 2 1 13 1 10 11 2 1 15 3 2 1 10 11 2
3 9 2 3
15 3 10 9 13 13 1 10 9 2 3 13 10 9 11 2
6 9 3 0 7 0 2
33 16 3 13 2 3 13 10 9 0 2 3 10 2 9 2 2 3 15 13 1 10 9 10 9 0 15 13 1 10 9 1 9 2
5 10 9 13 15 2
50 10 9 13 16 10 11 2 1 9 7 1 15 2 3 7 3 2 1 10 9 15 13 2 13 13 10 9 1 13 10 9 15 13 10 9 1 9 2 10 9 0 1 15 13 10 9 1 10 9 2
17 16 10 11 13 10 9 1 9 2 1 9 7 3 1 9 0 2
19 15 13 3 0 2 15 13 3 3 0 7 0 16 10 9 1 10 11 2
10 13 3 1 10 9 1 9 1 9 2
19 10 11 3 13 12 9 1 10 9 2 7 3 13 0 13 16 13 13 2
15 10 11 13 10 10 12 9 2 7 15 13 16 13 13 2
79 1 15 2 10 0 9 1 10 11 13 13 15 10 9 2 13 2 11 2 2 11 1 9 2 1 10 9 1 10 9 0 0 1 10 9 0 1 10 9 7 10 9 2 1 10 0 9 1 10 9 1 10 11 2 11 2 7 1 15 15 13 1 10 10 9 1 9 0 1 9 1 10 9 0 1 10 9 0 2
23 1 15 2 10 9 13 16 3 13 0 13 1 10 9 10 9 1 10 9 1 10 9 2
14 10 9 1 11 13 10 9 1 9 13 1 10 9 2
54 10 0 9 13 1 10 9 1 10 9 13 1 10 9 2 1 10 9 1 9 2 1 10 9 0 7 1 10 9 1 9 15 13 1 4 13 1 10 9 0 2 0 9 2 1 10 9 7 9 1 10 0 9 2
20 10 9 2 1 13 3 3 2 13 4 13 1 1 10 9 1 10 0 9 2
32 10 0 9 1 10 9 13 1 10 9 1 10 9 3 0 2 15 9 13 1 12 7 3 13 13 13 3 1 13 12 9 2
21 3 12 9 13 15 13 2 1 9 1 10 9 2 1 13 3 9 2 3 9 2
42 2 7 3 2 3 2 2 3 13 16 3 13 1 13 2 13 3 1 13 9 13 1 13 3 10 9 2 2 13 10 9 1 10 11 2 15 13 1 13 10 11 2
16 1 10 9 1 10 11 2 2 10 9 3 13 1 13 2 2
30 3 1 10 11 2 10 9 1 10 11 1 10 11 13 13 0 9 1 9 1 10 9 13 1 13 9 1 10 11 2
35 1 10 10 9 1 9 2 10 9 13 1 4 13 16 10 9 3 13 13 3 2 2 1 12 1 12 9 2 2 1 10 2 11 2 2
9 9 13 1 9 1 10 9 1 11
5 9 13 3 1 11
14 10 9 3 13 9 2 1 1 15 15 15 10 13 2
37 7 2 10 0 9 1 10 9 15 13 10 11 1 10 11 1 10 11 2 1 10 9 0 1 11 2 13 13 10 9 1 10 9 1 10 9 2
44 13 1 11 2 10 9 13 13 10 9 0 1 10 9 1 3 1 10 9 2 3 2 1 12 9 2 13 4 1 4 4 10 10 9 7 1 4 10 9 1 10 10 9 2
25 3 2 1 10 9 1 9 1 15 13 10 2 9 2 2 10 9 3 13 9 3 1 10 9 2
6 2 13 13 15 3 2
32 13 13 13 10 9 1 13 10 9 1 10 11 7 13 1 9 1 10 9 0 2 2 13 2 13 16 13 10 9 9 12 2
26 10 9 2 1 10 9 2 13 13 15 1 10 9 1 9 1 11 1 10 10 9 1 2 9 2 2
12 10 9 0 7 1 10 10 9 13 15 0 2
15 2 15 13 1 10 10 9 10 9 2 2 13 10 0 2
10 10 9 1 11 13 4 1 4 13 2
12 1 3 2 10 9 13 1 9 7 1 9 2
36 9 7 9 13 3 3 2 16 3 13 13 12 9 2 7 9 13 9 1 9 15 10 9 2 1 9 1 9 7 9 1 9 3 13 13 2
9 9 2 9 1 10 9 1 12 9
4 11 1 9 0
34 10 9 11 13 1 10 9 2 1 10 0 9 13 1 11 2 1 11 2 10 0 9 0 1 10 9 2 13 10 9 1 12 9 2
20 10 0 0 13 13 1 10 10 9 1 12 1 9 1 12 2 1 12 9 2
26 10 9 13 10 10 9 1 12 9 2 13 3 1 12 9 0 7 10 0 9 13 1 10 0 9 2
16 1 13 13 10 10 9 1 12 9 2 12 9 7 12 9 2
48 10 11 3 13 2 10 11 2 7 3 13 1 13 2 1 10 11 1 10 9 3 2 1 10 9 2 1 10 11 2 1 0 9 3 1 10 9 1 10 9 1 10 9 1 12 9 2 2
39 7 1 10 9 1 11 13 3 1 13 10 9 1 10 9 11 2 13 1 10 9 1 10 0 11 1 11 7 13 1 10 9 0 1 10 10 9 0 2
29 3 16 2 3 2 10 0 9 1 10 9 2 10 11 2 13 10 11 3 2 10 9 0 2 2 1 13 11 2
43 7 10 9 13 3 16 13 1 10 9 1 10 9 2 3 12 12 9 1 10 9 1 10 12 9 2 0 1 10 9 1 11 7 2 13 2 1 10 0 9 0 2 2
14 1 13 9 2 10 11 13 1 13 9 1 10 11 2
29 7 1 13 15 1 10 11 2 3 13 9 2 3 2 1 10 9 2 15 3 3 13 10 9 3 1 10 11 2
9 13 16 13 1 13 10 11 11 2
72 1 10 9 3 0 2 7 3 13 1 10 10 9 2 13 9 1 11 7 1 11 2 3 2 9 15 2 1 11 7 11 2 13 10 9 1 9 0 0 1 2 1 10 9 12 2 13 9 3 1 10 9 0 7 0 1 10 9 0 1 10 9 2 3 1 10 9 1 10 9 0 2
30 13 10 9 1 10 9 1 13 10 9 0 1 10 10 9 2 15 13 1 13 10 0 1 9 1 9 1 10 9 2
26 10 9 0 2 1 10 10 9 0 2 13 15 9 2 7 2 16 13 2 10 10 9 1 10 9 2
44 13 15 1 15 10 2 9 2 2 16 10 9 2 15 15 13 3 1 1 10 9 12 2 13 13 3 1 2 9 2 2 7 13 1 10 9 1 11 3 2 9 0 2 2
58 1 15 2 13 16 13 0 10 9 2 2 2 7 2 3 3 1 10 0 9 2 15 13 13 13 1 10 10 9 2 3 3 13 2 1 9 7 0 9 7 1 9 3 0 16 15 13 1 10 9 13 7 9 0 13 7 13 2
152 1 11 2 15 13 9 1 10 9 0 1 9 0 1 10 10 2 1 0 9 2 9 1 10 3 0 9 0 7 9 1 10 0 7 0 9 0 7 0 1 10 9 2 11 2 10 10 9 2 13 1 10 13 9 1 9 2 1 16 13 10 9 1 10 9 3 10 9 1 10 9 1 10 9 2 9 13 13 9 1 10 10 0 9 2 13 3 13 2 3 10 9 2 3 1 9 0 2 13 3 3 9 2 3 10 9 1 9 13 7 13 1 13 0 9 1 9 1 13 9 0 1 10 9 7 1 10 9 2 3 10 9 0 2 10 9 7 10 9 13 10 9 1 10 9 2 1 10 9 2 2 2
34 13 15 3 16 13 13 0 7 0 10 9 0 1 10 11 7 13 15 13 16 10 9 9 3 13 3 1 12 2 3 1 10 9 2
19 7 15 3 13 10 9 1 10 9 2 10 9 1 10 9 13 10 11 2
12 10 11 7 10 11 13 12 9 0 3 0 2
14 10 10 9 3 9 2 7 3 3 9 2 13 13 2
21 10 15 3 15 13 1 10 11 2 3 10 9 13 1 10 0 9 1 10 9 2
40 1 15 2 13 10 9 13 10 11 1 3 13 13 10 9 0 1 10 11 2 7 3 13 9 0 0 1 15 13 2 16 13 0 13 10 9 1 9 0 2
25 10 9 1 11 13 1 10 13 9 2 1 9 1 10 9 1 9 1 10 9 9 2 10 11 2
36 1 10 9 1 9 1 10 9 2 10 9 0 13 1 9 10 9 1 10 10 9 1 10 9 2 15 13 1 13 1 10 9 1 10 9 2
23 1 10 9 1 15 13 0 10 9 1 10 9 2 0 9 1 15 13 13 1 9 0 2
28 1 12 1 9 0 2 10 9 1 11 13 9 1 9 2 1 10 9 1 10 9 1 10 9 1 10 11 2
22 10 0 9 1 10 3 12 9 13 13 3 9 13 1 15 1 10 9 1 10 9 2
3 9 13 9
38 10 9 0 13 2 3 2 10 12 9 15 13 12 9 1 10 9 1 3 12 9 1 10 11 2 1 13 13 10 9 2 1 10 9 2 1 11 2
28 3 13 13 10 9 1 10 9 1 10 9 0 1 11 2 1 11 2 10 9 13 0 1 9 2 13 13 2
7 10 9 13 1 13 3 2
9 0 9 13 3 13 1 10 9 2
30 10 12 9 13 13 2 3 2 1 15 3 0 2 10 12 9 15 13 2 12 1 15 13 2 1 10 9 1 11 2
20 10 9 2 10 9 7 10 9 2 13 15 1 3 12 9 1 9 1 11 2
24 1 10 9 1 12 9 3 1 10 9 2 10 9 15 13 15 1 10 9 1 11 7 11 2
31 10 9 13 13 9 1 10 9 1 15 13 13 13 15 1 10 9 13 13 10 9 2 16 10 9 15 13 1 0 9 2
30 10 9 13 1 13 12 9 1 10 9 1 10 9 1 10 9 15 15 13 12 12 9 2 13 13 3 12 0 9 2
48 10 12 9 2 10 0 9 1 9 1 10 9 1 10 11 1 12 9 2 7 10 9 1 12 2 13 15 2 13 12 9 2 1 10 9 1 11 2 13 1 9 7 9 1 10 9 13 2
20 1 10 9 2 2 3 13 13 10 9 1 16 10 9 15 13 1 11 2 2
4 13 1 9 0
4 11 13 11 2
45 10 9 0 11 2 12 2 13 13 1 11 2 1 10 10 9 2 2 11 2 2 13 1 10 9 13 2 13 3 2 1 10 9 0 2 10 9 1 10 9 2 10 9 11 2
26 10 9 13 13 1 10 9 1 13 1 12 1 9 2 7 3 3 13 13 10 9 1 11 1 11 2
6 9 0 13 1 11 2
30 9 13 1 11 2 11 7 11 13 13 3 2 1 10 11 1 11 2 1 10 9 1 10 9 1 9 0 2 11 2
18 10 9 13 1 10 9 1 10 9 13 1 10 10 9 2 1 11 2
17 11 13 9 1 10 9 0 1 9 2 1 9 1 9 7 9 2
17 9 13 1 10 2 9 2 9 13 1 10 9 1 10 9 1 9
8 11 7 12 9 13 1 10 11
20 12 9 1 9 7 10 9 1 10 11 13 3 13 1 10 9 1 10 11 2
10 9 0 13 10 9 13 1 10 9 2
14 10 0 1 10 9 0 13 3 13 10 9 1 9 2
14 10 13 9 1 10 2 9 2 3 13 10 10 9 2
26 10 9 11 13 1 10 9 1 10 9 1 10 9 2 1 12 2 1 10 0 9 0 0 2 11 2
36 3 1 11 2 9 1 10 10 9 2 10 10 9 13 1 10 9 1 15 11 13 0 1 13 10 9 1 10 2 9 2 1 10 9 0 2
10 10 11 13 10 0 13 1 10 9 2
48 1 9 1 12 2 10 2 12 11 2 2 11 2 9 1 10 11 2 11 2 9 2 7 11 2 9 0 2 13 13 1 13 15 1 13 10 10 9 3 1 10 10 9 0 13 4 13 2
13 1 10 9 2 13 12 9 15 13 3 1 11 2
17 3 2 10 9 13 15 1 10 0 9 1 9 1 10 10 9 2
38 3 2 10 9 13 13 1 10 9 0 2 10 9 15 11 13 1 13 1 10 10 9 1 10 9 2 15 13 1 10 9 13 1 10 9 2 11 2
15 2 3 13 15 1 10 9 1 15 2 2 13 10 9 2
16 3 2 1 9 1 10 9 2 10 9 13 13 1 10 11 2
29 10 9 13 13 1 13 15 1 10 9 1 10 9 1 9 1 10 10 9 2 3 16 13 1 4 13 10 9 2
27 2 16 13 13 15 2 13 16 15 13 1 15 2 16 3 15 10 13 3 13 10 9 7 13 10 9 2
20 3 13 13 16 13 9 15 13 1 3 13 3 12 9 2 2 2 13 11 2
3 9 1 11
3 11 13 13
20 10 9 11 2 0 9 1 10 9 1 11 2 13 1 4 13 1 10 9 2
25 10 9 13 13 12 9 2 1 16 13 4 13 10 9 1 10 9 15 3 13 1 10 9 0 2
17 3 3 3 13 2 7 13 10 9 2 3 10 9 0 1 9 2
10 2 13 13 2 7 3 13 13 15 2
6 13 3 1 15 2 2
28 10 11 13 10 9 1 11 3 9 0 2 7 15 13 10 0 9 3 13 1 10 9 7 9 1 10 9 2
19 7 10 0 3 13 10 9 2 7 10 9 13 10 9 1 9 1 9 2
48 2 3 15 13 2 1 10 0 9 2 13 0 10 9 2 2 13 10 9 1 10 9 2 13 10 12 9 1 10 0 1 12 12 9 1 9 2 7 2 1 9 2 1 12 9 1 9 2
26 13 15 2 3 2 1 10 2 9 0 1 15 13 2 7 13 15 10 9 1 10 9 1 12 9 2
25 1 10 9 2 15 3 13 1 10 9 3 11 13 1 10 9 2 13 13 9 1 15 15 13 2
9 2 16 13 1 3 2 15 3 2
26 15 13 10 9 13 1 10 9 1 9 2 15 13 2 3 2 10 9 1 10 9 13 1 10 9 2
28 13 9 3 11 16 2 2 1 15 15 13 0 7 0 2 2 10 9 13 13 1 13 2 10 9 0 2 2
11 7 2 3 13 3 9 1 9 1 9 2
25 16 13 1 3 2 15 3 2 16 13 3 2 13 15 3 15 2 12 2 15 3 10 9 13 2
9 13 0 9 1 9 2 2 13 2
5 11 13 1 9 2
14 2 7 16 10 9 13 10 9 2 3 13 0 2 2
5 11 13 3 3 2
34 1 13 1 9 2 10 9 13 1 10 9 16 2 1 9 1 10 9 1 10 9 0 1 12 2 15 13 4 13 9 1 10 9 2
6 3 13 1 10 9 2
20 2 13 15 16 3 3 2 1 10 9 0 2 10 9 13 9 1 10 9 2
12 16 10 9 13 1 11 1 9 1 9 2 2
3 7 13 2
8 2 3 13 1 9 1 9 2
11 10 9 1 10 9 13 13 1 10 9 2
29 13 3 13 10 9 1 10 11 1 13 13 10 9 2 7 3 15 13 13 10 11 1 10 9 1 10 9 2 2
5 9 0 1 10 11
35 10 12 0 9 0 13 3 1 10 9 1 13 9 0 1 10 9 1 12 12 9 1 9 2 1 12 9 1 9 2 1 12 7 12 2
32 12 0 1 10 9 13 13 3 1 9 1 10 9 1 10 11 2 9 7 9 0 2 13 10 9 0 1 10 9 1 9 2
59 10 9 2 13 1 10 9 1 10 11 2 11 2 9 2 2 7 1 10 11 2 11 2 9 2 2 1 10 9 1 9 0 2 13 15 1 13 10 9 1 10 9 1 9 2 13 16 10 11 13 13 1 10 0 9 1 10 11 2
35 1 10 9 2 10 9 0 13 12 9 1 10 11 2 11 2 10 9 7 12 1 12 2 9 15 1 10 9 1 12 9 13 1 11 2
5 11 13 1 11 2
41 10 11 13 3 1 9 1 10 9 0 13 10 9 1 9 7 11 13 9 1 10 9 0 1 10 0 9 1 15 13 13 10 9 1 9 7 9 1 10 9 2
46 10 9 3 13 3 2 3 2 16 15 13 13 7 13 1 10 9 1 11 2 7 13 3 16 13 10 9 2 0 2 7 2 13 13 10 9 3 2 2 1 15 2 13 9 2 2
15 15 13 16 10 10 9 13 13 1 10 11 10 9 13 2
29 13 16 13 2 13 9 0 1 10 9 1 10 11 2 2 3 1 15 13 1 10 9 13 1 10 9 1 9 2
19 2 10 11 13 1 13 10 0 9 1 10 9 1 13 9 2 2 13 2
21 11 2 1 13 4 13 2 13 16 13 1 11 13 12 9 2 1 9 1 12 2
45 1 10 9 1 11 2 13 10 0 9 2 13 3 3 0 1 10 11 13 15 15 13 1 10 11 1 10 9 0 2 16 15 13 1 10 0 10 9 15 13 1 10 9 0 2
36 3 1 11 2 10 9 13 15 3 1 11 2 1 10 9 1 10 11 7 1 10 0 9 1 11 2 13 9 12 2 12 1 10 11 2 2
41 1 12 1 9 2 10 11 2 15 3 13 13 1 12 9 2 13 1 11 2 11 2 11 2 11 2 11 2 11 2 13 1 11 7 2 3 2 13 1 11 2
31 1 10 0 9 1 10 9 2 13 15 2 1 10 9 7 9 0 2 10 11 2 11 2 11 2 11 2 11 7 11 2
46 1 10 9 13 1 9 2 13 15 15 1 9 12 2 1 10 11 2 3 10 9 13 10 9 11 2 15 13 10 9 9 12 2 9 12 2 1 11 2 1 10 9 1 10 11 2
37 10 9 11 13 1 10 9 1 11 7 13 10 9 1 10 11 13 10 10 9 13 3 13 7 0 1 10 9 2 1 9 1 12 1 10 11 2
29 1 10 9 13 13 3 0 9 0 10 9 2 9 7 9 0 13 13 10 9 1 9 1 9 1 9 7 9 2
35 1 10 10 9 13 15 3 10 9 1 10 0 9 0 1 10 2 11 2 2 10 9 1 9 1 10 9 1 10 11 7 1 10 11 2
43 10 9 1 10 9 1 10 9 11 13 10 9 2 1 10 9 1 9 1 9 1 10 10 9 1 1 10 9 1 10 9 1 9 15 1 10 9 13 13 9 1 9 2
66 1 10 9 1 10 9 10 9 13 1 13 3 13 3 9 1 12 9 1 9 0 1 10 0 9 1 10 9 7 12 9 1 9 1 9 1 10 9 1 0 9 1 9 2 3 13 1 9 0 2 15 3 1 10 10 0 9 1 9 15 13 13 1 10 9 2
27 10 11 13 10 13 9 0 3 10 0 9 1 16 15 15 13 16 10 9 1 10 9 0 3 13 13 2
9 9 1 10 11 13 1 10 11 0
3 10 9 0
23 10 9 0 2 15 3 13 1 13 15 1 9 1 10 11 0 2 13 13 15 10 9 2
16 13 10 9 1 10 9 13 7 13 2 7 3 15 13 3 2
21 13 10 9 1 16 3 13 1 13 10 9 0 7 13 10 0 9 1 10 9 2
9 1 10 9 0 2 10 9 13 2
47 11 2 1 10 11 2 13 3 3 13 4 13 15 2 7 16 3 13 1 13 3 2 13 10 9 1 10 11 2 16 10 9 13 1 10 11 13 13 1 3 13 10 9 1 9 0 2
32 3 11 13 0 1 15 13 16 10 9 13 3 13 13 2 7 3 13 2 3 13 10 9 1 10 9 7 9 1 10 9 2
34 13 1 10 9 7 10 9 1 10 9 3 0 2 15 3 13 9 1 9 13 10 9 7 15 13 13 15 1 9 1 0 7 9 2
35 11 2 1 10 11 2 11 2 2 13 16 10 0 9 15 13 1 13 10 9 1 11 1 9 1 11 2 1 15 13 10 9 1 9 2
21 1 9 2 3 13 9 2 10 9 13 15 1 13 15 15 13 3 1 10 9 2
22 10 9 1 11 3 13 11 2 10 9 1 11 3 13 10 2 10 2 9 3 3 2
32 1 10 9 1 9 15 10 11 13 4 1 13 2 13 13 16 10 9 3 13 10 0 9 16 3 15 13 13 10 0 9 2
31 1 3 13 12 1 10 9 1 10 9 2 3 13 13 1 10 9 1 10 11 2 10 9 2 3 2 3 13 13 15 2
27 10 9 0 13 15 13 2 7 10 9 13 3 0 16 10 9 13 3 16 4 13 10 9 1 10 9 2
51 13 15 16 10 0 9 1 9 13 3 3 3 10 11 2 1 13 1 10 11 10 10 2 9 2 1 9 2 10 9 1 16 10 9 0 13 10 9 2 15 13 1 10 9 10 0 9 1 10 9 2
10 10 9 13 15 3 1 11 1 11 2
22 10 9 13 15 2 11 3 13 2 1 9 13 1 10 11 7 13 10 9 1 13 2
12 2 10 11 13 3 10 9 2 2 2 13 2
12 10 12 9 0 13 7 11 13 3 13 15 2
10 9 1 11 0 1 10 9 1 10 9
33 10 0 9 0 1 11 2 15 13 1 13 9 3 1 10 9 1 10 0 11 2 3 11 2 2 13 0 1 9 1 10 9 2
37 13 15 10 9 13 1 10 9 2 11 2 13 1 13 1 10 9 10 0 9 1 10 0 9 1 9 7 9 1 16 15 13 10 0 9 0 2
40 1 10 11 13 13 1 10 9 2 10 9 13 13 2 1 10 0 9 1 9 2 10 9 15 3 15 13 13 7 13 1 10 9 0 13 1 9 7 9 2
21 3 13 4 13 15 1 10 9 15 13 13 10 9 2 13 1 10 9 1 9 2
19 13 10 9 1 10 1 10 9 7 1 10 0 9 3 13 1 9 0 2
18 3 7 3 2 13 1 10 11 10 0 1 2 11 2 1 10 11 2
18 11 2 1 10 11 2 13 2 11 2 2 10 0 9 1 10 11 2
7 9 0 1 10 9 1 11
34 2 11 2 13 10 9 15 13 1 10 9 0 15 10 11 2 11 2 13 2 1 12 7 12 1 9 2 1 10 11 2 1 11 2
38 3 1 9 1 10 9 0 0 1 9 7 9 2 13 13 10 9 1 10 9 0 1 10 9 1 10 11 2 11 2 3 1 10 9 1 10 11 2
42 10 9 13 15 1 12 0 9 2 10 9 1 10 9 0 1 9 2 10 9 0 1 10 11 7 10 9 1 10 9 1 10 11 2 9 1 9 2 9 0 2 2
10 10 9 0 2 11 2 13 10 9 2
14 9 2 15 13 10 9 1 13 1 9 7 1 9 2
32 9 2 1 10 9 13 15 13 10 9 1 10 9 2 13 15 10 9 2 7 3 12 9 2 13 15 10 9 1 10 9 2
16 1 10 9 2 3 15 15 15 13 13 10 9 1 10 9 2
30 1 10 9 13 1 10 9 2 13 15 9 1 9 7 12 9 13 4 13 1 12 9 1 9 2 1 9 1 9 2
7 13 10 9 1 10 9 2
9 3 1 12 3 10 9 13 9 2
25 11 2 1 9 1 11 2 3 11 2 13 10 0 9 1 11 1 13 10 9 2 2 11 2 2
8 10 9 1 10 9 13 11 2
24 10 9 1 10 9 11 2 10 2 9 2 13 10 9 1 10 9 1 13 13 10 0 9 2
20 3 15 1 9 1 11 2 11 2 1 3 12 9 2 1 15 10 9 11 2
42 13 1 10 9 2 11 13 3 1 11 2 13 2 3 10 9 2 10 9 1 11 2 2 11 2 2 7 13 9 1 10 0 9 13 1 10 9 3 0 2 11 2
39 16 15 3 1 3 13 2 13 1 10 9 0 2 3 1 3 3 10 9 13 10 10 2 9 2 2 13 15 2 1 10 9 2 10 9 1 10 9 2
7 13 10 0 2 11 2 2
30 10 9 13 10 9 7 11 1 1 10 9 1 10 0 0 9 13 7 13 15 1 9 1 10 9 1 10 10 9 2
17 3 15 13 10 9 1 10 2 9 2 13 3 12 9 1 0 2
50 13 0 10 9 1 2 11 2 2 11 2 2 10 9 15 13 10 0 0 7 10 9 1 9 1 10 9 12 2 15 13 1 15 10 10 9 7 13 1 10 9 10 9 1 9 2 10 0 2 2
22 2 11 2 13 13 1 12 1 0 1 2 11 2 2 10 0 3 7 10 0 3 2
34 13 12 9 3 1 2 11 2 2 2 11 2 13 10 9 0 1 15 13 3 1 9 0 2 1 10 9 7 1 10 9 1 9 2
52 7 10 9 0 13 3 1 15 3 1 10 9 12 1 9 2 10 9 2 1 10 9 1 10 11 2 1 10 11 2 7 13 1 10 10 9 7 1 10 10 9 1 10 9 2 9 12 2 1 10 11 2
59 10 10 9 2 1 10 9 1 10 9 2 13 1 10 9 7 3 1 10 10 9 10 9 1 9 7 9 0 2 9 12 2 2 10 9 11 2 9 12 2 2 11 2 9 12 2 2 11 2 9 12 2 7 11 2 9 12 2 2
20 3 3 2 1 10 0 9 1 10 11 2 10 9 13 0 2 13 10 9 2
31 1 10 9 2 9 7 9 13 15 2 1 10 10 9 1 9 2 10 9 2 10 9 2 9 1 9 2 9 7 9 2
16 9 2 13 15 1 3 0 1 2 11 2 10 10 0 9 2
26 9 2 13 16 10 0 13 16 2 11 2 13 10 0 9 10 2 1 10 9 2 2 13 3 15 2
23 10 9 13 3 3 10 9 2 13 13 1 10 15 2 3 13 3 12 7 12 9 0 2
16 3 15 13 10 9 0 1 15 1 10 10 9 2 1 9 2
6 16 13 10 9 0 2
19 3 2 3 2 13 10 9 3 1 10 9 2 13 1 12 1 10 9 2
7 9 1 9 13 1 10 11
47 10 9 1 11 1 10 11 13 1 10 13 9 2 1 9 2 7 1 10 9 1 9 15 13 1 4 13 1 10 11 1 10 9 1 9 1 10 9 2 10 9 1 10 9 1 11 2
35 1 10 9 13 13 2 1 10 2 12 0 1 9 13 1 15 12 7 15 12 9 2 15 13 13 2 1 10 11 2 1 13 10 9 2
4 11 13 3 0
9 10 11 13 13 3 0 10 11 2
42 1 15 2 3 1 10 9 3 13 1 3 2 13 10 9 1 10 9 1 10 10 9 2 1 13 13 10 9 1 10 9 2 2 13 2 3 10 9 3 1 9 2
46 1 9 1 10 2 9 2 9 2 15 13 3 10 9 1 10 11 2 10 9 13 3 13 9 1 16 10 11 2 15 13 1 10 9 13 1 9 2 13 13 3 1 10 9 0 2
28 3 2 10 9 1 10 9 2 13 1 3 2 13 1 10 9 1 10 9 0 2 3 13 1 10 0 9 2
8 10 9 3 13 10 10 9 2
47 7 2 1 10 0 9 1 10 9 1 10 9 2 13 15 1 13 3 3 1 10 2 11 2 2 9 1 9 1 10 9 0 3 3 13 2 7 1 10 3 0 7 0 2 11 2 2
32 10 9 1 11 3 15 13 2 3 16 1 10 9 13 0 1 10 9 0 2 15 3 15 13 1 10 9 15 15 10 13 2
30 1 9 15 3 15 13 1 13 2 1 9 15 13 3 0 2 15 2 1 2 13 3 10 0 9 16 10 9 0 2
7 1 9 2 10 0 9 0
10 2 13 15 3 1 10 2 11 2 2
35 13 12 9 1 10 9 1 11 2 7 3 13 2 15 13 1 10 11 2 3 13 11 1 13 2 11 2 3 1 10 9 1 10 11 2
10 11 13 15 16 13 13 1 10 9 2
14 1 10 9 0 13 1 15 2 7 13 16 13 13 2
23 3 2 10 9 1 10 9 13 3 13 2 13 1 10 11 7 3 3 13 1 10 11 2
6 10 9 13 3 0 2
9 7 10 9 1 10 9 13 0 2
16 10 10 9 13 15 1 13 3 10 10 9 1 10 1 11 2
39 3 13 16 13 10 0 9 15 13 1 10 9 2 15 3 13 3 13 7 0 2 7 15 13 2 3 2 16 13 13 10 9 0 1 10 2 11 2 2
34 13 1 13 1 11 16 13 3 0 1 10 11 2 3 10 9 3 13 3 2 3 3 2 10 9 0 1 10 9 1 9 1 11 2
5 13 1 10 11 2
5 7 13 3 0 2
18 7 13 13 16 10 9 0 1 10 10 0 9 13 13 0 7 0 2
38 10 9 0 2 1 15 10 9 2 13 13 3 13 2 2 13 11 15 3 13 16 2 11 2 13 10 10 0 9 1 10 11 1 9 1 10 9 2
5 10 9 1 10 9
4 10 9 1 11
37 3 2 1 0 9 1 2 9 2 2 13 1 13 12 1 10 0 9 1 10 9 15 13 13 10 0 9 1 10 9 1 10 9 3 15 13 2
54 13 15 1 10 9 1 10 11 2 10 3 0 9 1 10 9 1 10 9 1 9 1 9 0 7 10 11 2 15 1 12 9 13 12 9 1 10 9 1 9 1 9 1 10 11 1 10 9 15 15 13 10 9 2
16 9 0 1 11 2 10 11 13 1 10 11 2 1 10 9 2
4 1 10 9 2
27 1 10 9 1 10 11 2 13 1 10 11 1 10 11 2 13 13 15 10 9 2 11 2 2 1 11 2
35 10 9 13 11 2 9 2 2 11 2 9 2 2 11 2 9 2 2 11 2 9 2 2 11 2 9 2 7 11 2 9 1 9 2 2
4 1 10 9 2
24 10 9 7 10 10 9 2 11 2 13 10 9 1 12 3 10 9 1 15 15 13 9 0 2
26 2 1 13 10 9 0 1 10 12 9 2 3 1 15 12 3 10 11 15 13 3 2 2 13 11 2
26 2 16 10 9 1 10 12 9 2 9 7 12 12 2 13 0 2 13 10 9 3 1 10 0 2 2
21 11 3 15 13 3 1 10 9 0 15 2 3 2 13 13 2 10 9 7 9 2
13 2 10 9 13 0 1 15 7 3 15 13 3 2
6 13 3 1 15 13 2
23 3 16 13 13 1 9 0 1 15 15 13 1 11 2 7 2 3 13 0 2 9 2 2
13 1 9 2 10 10 9 13 0 1 10 9 0 2
17 2 10 3 0 13 13 15 1 10 9 2 1 0 10 9 11 2
30 10 2 0 2 11 3 13 16 13 15 12 7 10 9 7 10 9 13 9 7 9 7 3 13 10 9 1 12 2 2
24 1 10 11 2 10 9 1 10 9 12 1 15 12 13 10 9 0 1 10 9 1 10 9 2
25 1 13 10 9 1 9 0 2 10 0 11 13 10 9 1 9 7 10 9 1 9 7 1 9 2
23 12 1 10 9 1 10 0 11 13 3 13 10 0 9 1 10 9 1 11 7 1 11 2
35 1 10 9 2 15 13 10 10 1 10 12 9 2 1 10 9 1 9 2 15 13 13 1 16 10 9 1 10 12 9 3 13 10 9 2
39 10 10 9 15 13 1 10 10 2 9 1 9 2 2 3 15 13 10 11 2 16 13 16 10 9 13 10 1 13 1 10 9 11 16 1 15 1 11 2
19 3 2 10 0 2 9 2 13 9 15 3 13 1 10 9 12 1 11 2
22 10 11 2 1 10 9 2 1 15 13 1 12 1 12 13 15 3 1 10 0 9 2
28 13 2 1 15 12 2 15 15 13 10 9 3 0 7 2 1 15 2 13 15 15 13 10 0 9 1 9 2
13 3 10 9 1 10 11 13 13 2 15 13 15 2
10 3 15 13 10 9 1 10 10 9 2
14 10 9 3 0 16 3 13 0 13 3 1 10 9 2
13 3 2 11 13 16 13 13 0 13 3 3 3 2
17 2 13 16 13 0 13 3 3 1 10 9 2 2 13 10 9 2
21 2 13 16 13 13 0 13 15 10 1 10 9 1 10 9 7 1 10 10 9 2
11 13 16 13 3 0 13 1 1 10 11 2
27 10 0 9 13 13 16 13 10 9 3 1 15 15 13 10 11 7 16 13 1 10 15 1 10 15 2 2
53 1 11 2 10 9 13 10 9 1 10 9 3 13 1 10 9 2 9 10 1 13 10 9 7 13 10 9 1 10 0 9 2 15 3 13 10 9 1 13 1 10 0 9 1 10 9 1 10 0 9 1 9 2
45 10 9 13 3 13 1 11 7 11 2 10 1 12 9 2 1 12 1 10 11 2 15 13 13 2 12 2 2 1 10 9 2 1 10 11 2 1 10 11 2 7 1 10 11 2
39 3 3 2 13 10 0 11 2 15 13 13 3 10 11 2 1 12 2 7 10 11 2 9 1 12 9 1 10 11 1 10 11 2 2 10 1 12 9 2
32 10 9 0 1 10 0 13 3 15 10 9 1 10 9 2 16 10 0 7 10 0 1 10 9 0 13 13 3 1 12 9 2
36 9 0 1 10 11 2 15 2 3 1 2 1 10 9 13 2 13 13 10 11 2 13 1 13 10 9 0 2 3 13 10 2 9 0 2 2
24 12 9 1 12 9 13 3 15 1 10 9 15 13 10 9 1 10 9 0 1 10 9 0 2
31 3 2 10 9 13 1 10 9 1 10 11 2 15 13 13 1 11 1 12 7 13 1 13 10 0 9 1 10 9 0 2
69 1 10 0 9 2 10 11 13 13 10 9 2 12 2 1 11 1 10 11 2 3 10 9 0 2 12 2 1 10 11 1 10 11 7 1 10 11 1 10 11 2 13 13 1 12 10 9 13 1 10 0 9 2 15 13 12 9 1 15 13 2 12 9 7 3 12 9 3 2
40 10 9 13 3 13 2 13 3 1 9 0 1 9 0 2 7 10 0 9 1 10 11 13 15 0 2 13 10 9 1 9 2 3 13 2 1 10 9 0 2
17 10 9 13 15 1 10 9 1 10 9 1 9 1 9 1 10 9
31 9 2 13 10 10 9 1 9 1 11 2 13 15 1 10 9 1 10 11 13 10 9 1 11 1 10 9 1 10 9 2
14 7 3 13 10 9 1 10 9 2 3 12 0 9 2
19 13 12 9 2 3 2 13 3 1 10 9 2 9 1 15 15 13 3 2
36 13 16 1 10 10 9 2 15 13 3 12 7 12 9 2 13 3 10 9 2 1 13 13 1 10 9 15 13 3 3 0 16 10 1 15 2
12 10 9 1 9 7 9 13 3 1 0 9 2
13 9 2 10 10 9 13 15 15 13 1 9 12 2
6 13 15 3 15 13 2
11 11 2 11 12 2 1 10 9 0 1 11
4 9 1 10 9
46 1 10 9 1 15 10 11 13 13 10 9 1 10 9 2 13 12 12 9 0 1 10 11 2 1 10 9 1 11 7 1 10 11 2 13 1 13 1 10 9 1 10 9 3 13 2
21 13 1 10 11 2 13 15 3 1 10 9 1 10 9 13 7 1 10 9 13 2
37 10 11 13 10 0 9 0 1 10 11 2 13 12 9 1 10 9 1 10 9 0 1 12 9 1 10 0 9 0 2 7 12 9 1 10 11 2
40 1 9 1 10 11 1 12 12 9 1 9 7 13 10 0 1 12 12 9 2 10 11 13 1 12 12 9 0 2 1 10 9 2 1 12 12 9 1 9 2
74 3 13 1 13 2 16 1 10 9 13 1 10 9 12 1 9 1 9 1 10 9 0 11 2 9 11 2 1 11 2 10 9 1 10 9 1 11 2 11 2 3 15 13 3 10 9 1 10 11 2 7 3 15 12 0 13 1 10 9 15 13 10 9 0 11 7 10 9 11 2 0 9 11 2
95 15 13 16 10 9 2 13 1 0 9 1 10 2 9 2 0 2 13 4 13 1 13 1 10 0 9 13 1 11 7 10 11 7 2 13 10 9 1 10 9 2 11 13 10 9 0 1 11 7 11 13 10 9 1 10 9 0 1 16 15 13 10 0 9 1 10 0 0 1 10 9 0 1 10 10 0 9 2 2 13 15 3 9 0 16 11 13 1 4 13 2 10 2 9 2
60 1 15 13 10 0 9 1 10 2 0 9 2 2 1 9 12 2 12 9 2 11 13 1 12 9 1 0 1 10 2 9 2 1 11 2 1 11 12 2 7 13 13 3 1 10 0 9 1 10 9 1 9 2 13 0 9 1 10 9 2
14 2 10 9 13 3 13 7 13 13 1 10 9 2 2
20 11 3 13 1 10 2 9 2 10 0 9 2 7 13 10 9 1 10 9 2
7 2 13 16 13 3 3 2
24 10 9 13 15 2 3 3 7 3 1 10 9 2 15 15 13 1 13 10 9 1 10 9 2
13 10 9 13 3 2 7 10 9 3 13 13 2 2
39 1 11 2 10 9 0 13 10 9 1 10 0 2 3 13 1 10 10 11 9 12 0 16 10 0 9 2 1 9 2 15 15 13 1 10 2 9 2 2
41 10 9 0 13 1 3 15 13 1 10 9 1 10 9 2 15 13 11 3 13 2 3 16 13 1 11 10 9 0 15 13 13 10 2 9 2 1 10 10 9 2
5 13 0 2 3 2
13 3 1 15 2 1 10 11 13 15 3 1 11 2
8 7 13 15 10 15 1 3 2
18 16 1 10 0 9 0 10 9 3 13 1 12 2 7 1 12 9 2
4 1 13 11 2
24 2 13 16 10 11 13 1 10 9 1 15 15 13 1 10 9 2 1 10 9 1 11 2 2
29 9 2 15 13 10 9 15 3 13 1 10 9 2 7 1 10 11 2 1 10 9 0 13 1 15 2 11 2 2
24 9 2 13 15 3 13 16 10 9 1 9 0 13 13 10 9 0 7 1 9 15 13 13 2
12 10 9 1 9 0 13 13 3 1 12 9 2
26 3 13 10 9 2 0 2 1 0 9 2 13 1 10 10 9 15 10 9 13 13 1 12 1 12 2
91 13 15 0 13 10 9 1 9 0 1 10 11 2 11 2 7 1 10 11 2 1 10 9 0 1 10 9 1 9 0 7 2 3 16 15 2 16 10 9 13 3 2 1 10 9 2 16 13 13 1 16 10 0 9 13 9 1 9 7 1 9 1 10 11 7 1 10 11 2 16 13 13 16 10 9 0 7 0 15 13 1 15 13 1 10 11 7 1 10 11 2
18 7 10 9 13 4 4 1 10 9 0 7 3 3 4 1 10 11 2
6 2 13 1 10 9 2
4 9 1 10 9
5 10 9 1 9 0
18 12 9 2 10 9 1 11 7 15 0 2 13 15 1 13 1 9 2
33 10 0 13 1 13 16 13 13 1 10 9 1 10 9 1 9 7 16 13 13 9 1 13 10 9 1 9 0 1 10 9 13 2
2 3 2
32 16 10 9 1 9 1 11 13 15 16 3 12 9 1 10 9 1 9 0 13 9 2 1 15 13 2 1 12 7 12 9 2
26 1 16 15 13 10 9 3 2 13 9 15 13 1 4 2 13 2 2 15 13 1 10 9 1 9 2
12 1 15 2 1 11 10 9 13 10 9 3 2
23 2 1 10 9 2 3 13 3 10 9 2 3 13 16 13 10 9 15 13 13 10 9 2
12 3 2 1 15 3 3 13 2 13 1 13 2
17 3 3 3 15 13 13 10 9 7 10 9 0 2 2 13 11 2
26 10 9 13 16 3 13 13 1 13 15 1 10 9 2 7 13 1 10 9 16 10 9 3 13 2 2
13 3 3 15 13 16 10 9 1 10 9 15 13 2
39 3 3 2 10 11 13 1 13 1 10 10 9 2 1 10 9 1 10 9 1 10 11 2 3 11 13 2 7 3 3 1 10 9 3 10 9 15 13 2
22 3 16 2 3 2 10 9 2 1 10 9 2 13 9 2 10 9 13 7 13 9 2
22 11 13 13 10 15 15 13 1 10 9 7 15 13 1 13 10 9 3 1 10 9 2
5 10 9 1 10 9
23 10 9 3 13 10 9 2 13 13 10 10 9 1 9 2 15 13 1 15 10 0 9 2
7 10 9 3 13 2 13 2
80 11 7 11 13 10 0 9 0 2 10 9 1 11 2 9 13 1 13 10 9 0 15 1 10 9 13 3 3 16 0 2 13 10 9 1 9 1 10 15 15 13 1 10 10 9 3 0 1 10 9 1 10 0 9 2 7 10 9 1 11 2 16 13 3 15 13 13 10 9 1 10 9 2 13 3 10 10 9 0 2
90 10 9 0 1 13 12 9 0 2 3 7 3 13 1 11 2 10 9 7 10 9 1 13 2 1 15 2 3 2 10 9 1 11 13 0 2 2 13 16 2 3 16 10 9 2 10 9 13 10 9 1 9 2 10 9 1 10 9 1 10 9 1 10 9 7 2 1 15 2 10 10 9 0 2 3 3 3 13 1 10 9 2 13 10 9 7 13 10 9 2
29 13 15 12 1 10 0 9 1 10 9 1 10 9 2 10 9 13 2 3 3 2 13 3 10 0 9 0 2 2
9 3 3 1 13 3 11 15 13 2
5 9 3 1 10 11
65 10 9 11 2 10 9 11 2 10 9 11 2 10 9 11 7 10 9 11 13 10 0 1 13 10 9 1 10 0 9 1 10 11 1 9 2 9 15 13 1 4 13 1 11 2 11 2 7 15 13 13 1 12 9 1 9 2 3 12 12 9 2 1 9 2
36 11 2 9 12 1 10 2 9 2 0 2 13 10 9 1 13 10 9 11 2 12 7 12 2 2 13 1 15 13 1 10 9 1 10 9 2
28 10 9 13 12 9 1 10 9 2 1 12 1 10 9 2 15 4 1 13 10 0 9 1 12 9 10 9 2
22 11 13 13 1 10 0 9 10 9 11 2 15 13 10 9 11 2 12 7 12 2 2
45 11 2 15 1 10 0 9 13 13 10 9 2 3 1 13 13 9 1 10 10 9 1 10 9 11 2 13 1 13 10 10 0 9 2 13 10 9 1 10 10 9 1 9 0 2
37 11 2 15 13 10 9 11 2 12 2 12 7 12 2 2 13 13 1 10 0 9 10 9 1 10 9 1 11 2 11 2 7 11 2 11 2 2
37 3 11 3 13 9 1 13 10 9 11 2 12 2 12 7 12 2 2 13 3 1 10 9 11 2 15 13 10 10 9 11 2 12 7 12 2 2
32 3 2 10 0 0 11 13 10 9 3 0 1 10 0 9 2 13 10 9 11 2 0 1 9 3 0 2 1 12 7 12 2
23 1 10 0 9 2 11 13 10 9 1 10 9 1 11 2 11 2 7 11 2 11 2 2
8 2 11 2 1 9 13 1 11
23 15 13 15 12 9 16 10 9 1 10 11 2 13 11 2 10 9 15 13 1 10 9 2
25 2 10 9 13 10 9 1 10 9 2 1 10 9 15 10 9 13 13 1 10 9 3 13 2 2
45 11 2 9 1 10 2 11 2 2 10 9 0 1 10 9 1 11 7 13 1 11 2 13 1 10 2 11 2 16 13 1 13 10 2 11 2 1 10 9 1 11 7 10 9 2
4 13 9 1 11
37 10 9 1 10 9 0 11 2 9 1 2 11 2 2 13 1 10 9 1 10 11 2 13 3 13 2 13 3 10 11 2 1 10 9 1 11 2
38 10 9 1 10 9 0 13 12 1 10 12 9 13 1 9 2 1 10 9 1 11 2 9 1 10 9 1 10 9 0 3 15 13 16 11 13 13 2
22 10 9 1 2 11 2 2 9 0 1 10 11 2 13 1 10 0 11 15 3 13 2
53 10 10 9 13 13 1 9 2 1 10 9 1 9 2 1 10 9 13 1 10 9 11 2 15 13 10 9 1 10 9 2 10 10 9 1 10 9 1 10 9 7 10 9 0 2 1 9 1 9 1 10 9 2
45 1 10 9 15 13 1 10 9 1 9 1 10 9 2 1 10 9 1 9 0 2 10 9 13 1 11 13 16 2 10 9 1 11 2 13 11 2 15 13 1 9 1 9 2 2
8 13 1 12 1 9 1 12 2
7 9 2 6 2 1 15 2
36 15 13 13 16 2 1 10 9 1 15 13 13 10 9 1 10 9 1 10 9 2 13 3 13 16 10 9 0 13 1 10 11 13 13 0 2
10 15 13 10 0 9 7 9 3 0 2
21 10 9 1 16 10 9 1 9 3 13 2 3 2 3 0 3 13 13 10 9 2
36 9 2 13 13 16 3 15 13 1 10 9 1 12 9 7 16 10 9 1 10 9 13 13 2 1 10 9 2 1 13 1 12 9 7 3 2
71 10 10 9 13 10 9 9 2 13 1 10 9 1 9 2 13 3 1 10 9 9 1 9 7 1 9 2 7 10 9 0 2 15 1 10 9 1 10 0 2 13 2 3 2 1 10 9 1 9 1 9 1 10 9 1 9 7 1 10 9 1 9 2 9 2 9 7 9 1 9 2
53 10 9 1 11 2 10 9 1 9 1 0 9 2 13 2 1 10 9 2 1 12 2 9 2 2 3 3 16 15 12 15 13 0 9 1 10 9 1 10 11 2 10 9 0 13 1 10 9 1 12 9 2 2
49 10 9 1 10 11 1 12 9 2 9 1 9 1 0 9 2 0 1 10 9 1 10 9 13 1 10 9 0 0 2 3 13 1 4 13 1 10 9 1 9 7 3 13 13 12 2 9 2 2
40 1 10 11 2 11 2 2 11 13 12 9 1 9 7 13 12 9 1 9 2 1 10 0 12 9 1 12 2 15 13 1 10 9 0 1 12 9 1 9 2
29 10 9 1 9 1 10 9 1 10 9 13 2 13 15 1 12 9 2 1 12 9 1 10 12 0 9 1 12 2
42 1 9 13 15 10 9 1 12 9 1 10 9 7 10 9 1 12 9 1 10 9 2 15 13 10 9 1 12 9 1 10 9 0 0 2 1 10 10 9 1 12 2
39 10 9 1 10 11 2 11 2 13 12 9 1 9 1 9 1 10 9 2 1 0 9 1 12 2 3 10 9 1 10 11 13 12 9 1 10 10 9 2
25 2 10 9 13 13 3 0 1 10 9 2 3 1 9 3 3 2 2 13 10 9 1 10 9 2
21 2 13 1 15 13 2 1 9 1 13 10 9 1 10 9 7 1 10 9 2 2
20 10 9 0 1 10 9 0 1 9 0 2 11 2 9 1 10 11 2 13 2
10 2 13 16 13 9 1 11 13 2 2
22 7 13 1 9 15 3 13 13 9 15 3 13 13 3 10 9 15 11 13 1 13 2
27 10 9 0 1 2 11 2 13 15 1 10 9 0 2 9 3 10 9 13 4 13 3 16 1 10 9 2
48 0 16 3 13 10 0 9 3 1 9 2 7 3 1 10 9 13 10 9 1 10 0 2 7 10 9 13 1 11 3 1 11 13 3 3 9 0 2 3 13 3 1 10 9 1 10 9 2
50 3 0 16 15 2 10 9 13 1 11 3 13 10 0 9 2 7 13 3 10 9 1 2 11 2 2 1 10 9 13 1 10 10 9 7 1 10 10 0 2 7 1 10 9 1 13 1 9 0 2
46 0 1 10 9 1 11 13 9 7 9 2 7 10 9 15 13 13 9 1 10 9 1 10 9 13 2 16 15 13 1 10 9 3 9 2 7 2 16 15 13 2 10 9 3 0 2
16 13 2 1 15 2 9 0 7 0 2 1 13 10 9 0 2
29 1 3 13 10 9 1 10 9 0 2 10 9 1 9 7 1 9 2 7 3 1 10 9 1 13 7 1 9 2
27 10 9 13 13 13 2 3 2 10 12 9 15 13 10 9 0 1 11 7 11 2 9 2 9 7 9 2
22 2 11 13 13 11 1 10 10 9 2 3 13 10 9 7 10 9 2 2 13 11 2
22 3 3 13 9 1 9 2 16 2 10 10 0 9 13 13 2 13 10 9 0 2 2
15 1 10 10 9 2 10 10 9 3 13 13 1 10 9 2
18 2 15 13 10 9 0 7 10 10 9 13 13 15 2 13 15 2 2
22 10 9 13 16 11 13 11 1 10 11 2 15 1 12 2 15 3 13 2 0 2 2
14 2 3 13 15 1 15 15 13 10 9 1 13 0 2
7 3 13 9 1 9 2 2
9 3 3 2 3 2 13 10 9 2
7 2 1 10 9 0 2 2
18 3 1 10 2 9 1 10 9 2 7 1 10 9 1 10 9 0 2
46 2 1 10 9 2 10 9 0 13 13 1 10 11 2 13 10 9 1 10 11 2 15 13 3 12 9 1 9 2 2 13 11 2 15 2 3 2 13 10 2 9 2 1 10 9 2
44 2 10 11 13 10 0 9 3 11 13 10 9 0 2 3 10 9 0 2 15 2 1 12 2 16 3 13 10 9 1 10 9 1 11 2 13 3 13 1 9 1 10 11 2
8 2 10 9 0 1 13 13 2
9 11 13 15 1 10 9 1 11 2
10 11 2 1 10 11 2 13 10 15 2
11 10 9 13 7 10 9 1 10 9 13 2
3 9 2 12
28 2 10 9 15 13 1 10 9 13 0 2 0 2 13 3 2 10 9 13 2 2 13 10 9 1 10 9 2
9 2 10 10 9 13 13 9 0 2
20 1 15 13 2 10 9 13 13 1 9 1 9 7 3 1 9 2 2 13 2
28 1 13 2 10 9 13 10 9 1 10 9 2 2 1 13 10 9 7 2 16 0 2 13 1 10 9 2 2
35 10 9 13 9 1 10 9 1 10 9 1 9 0 1 10 9 1 11 7 1 10 9 1 10 11 2 9 9 1 10 9 1 9 3 2
6 9 0 13 9 0 2
24 11 7 15 1 10 10 9 13 3 10 9 11 3 2 9 0 2 1 10 9 1 10 11 2
24 3 0 2 10 9 1 10 2 9 2 13 1 16 13 2 13 3 2 10 9 1 10 9 2
8 3 2 10 9 13 3 0 2
38 3 3 10 9 13 3 13 15 2 3 10 9 15 13 1 9 2 3 10 9 3 13 3 13 1 9 2 1 15 15 10 9 1 9 13 13 13 2
9 10 9 13 1 11 13 3 0 2
20 1 10 9 15 15 13 13 10 9 2 3 10 9 1 10 9 1 10 9 2
12 9 12 2 13 1 10 9 10 2 3 0 2
20 9 12 2 13 10 9 2 9 7 9 2 13 3 1 10 0 9 1 9 2
11 9 12 2 13 1 10 9 2 13 12 2
41 9 12 2 13 10 9 1 10 9 10 1 10 10 9 2 7 1 15 1 10 9 13 1 12 1 12 2 0 2 0 2 3 2 2 13 10 0 9 1 9 2
22 9 12 2 13 1 10 0 9 7 13 13 12 7 15 9 1 9 13 9 3 13 2
5 16 3 2 6 2
3 2 13 2
18 16 3 2 13 10 9 12 1 12 13 15 13 3 13 10 9 0 2
20 13 2 3 2 13 10 0 9 1 15 1 10 9 1 9 1 10 10 9 2
16 7 2 1 13 1 12 1 12 2 13 13 1 12 1 12 2
5 7 13 9 0 2
11 13 9 1 9 1 9 1 10 10 9 2
14 1 13 10 9 2 10 9 1 10 11 13 12 9 2
22 10 9 1 11 2 1 10 2 9 2 1 11 2 13 13 10 12 9 1 10 0 2
7 9 1 12 9 13 1 9
5 11 13 9 1 11
22 10 9 1 10 0 11 13 4 1 13 1 10 9 0 10 9 1 10 9 1 11 2
44 10 11 0 13 2 1 10 9 1 9 2 10 9 1 9 1 9 1 10 9 1 10 9 7 13 10 9 1 9 1 10 9 1 10 12 9 3 1 10 9 13 1 12 2
43 10 9 13 1 10 9 0 13 1 9 10 9 1 10 11 1 10 9 1 9 0 2 13 15 10 0 9 1 9 2 7 13 15 9 1 13 10 9 1 10 10 9 2
50 11 13 1 9 0 1 13 16 10 11 1 10 9 2 3 2 1 10 10 9 0 2 2 13 13 10 2 9 3 13 1 10 9 0 2 2 1 10 9 1 10 11 7 2 1 15 2 3 13 2
27 10 9 0 13 2 3 2 10 9 9 1 13 10 9 15 13 10 9 2 10 9 0 1 10 9 2 2
16 10 9 1 10 11 13 7 13 3 10 9 1 10 9 0 2
25 2 10 9 2 1 13 10 9 2 13 10 9 0 3 1 10 9 0 2 2 13 10 9 11 2
21 1 10 11 2 11 13 1 13 10 9 1 10 9 1 9 1 10 10 9 0 2
26 2 15 13 7 13 1 11 1 1 10 12 9 7 1 15 13 1 10 9 10 9 1 10 9 2 2
39 3 2 10 9 0 13 2 9 1 9 13 2 7 13 1 13 10 9 1 10 9 1 10 9 2 1 15 13 10 9 1 9 1 10 9 1 10 9 2
7 9 0 1 9 1 10 9
6 11 13 9 1 10 11
30 10 9 2 11 2 13 3 2 16 13 13 1 10 9 10 9 1 10 9 0 15 10 10 9 13 1 10 0 9 2
49 10 9 2 13 1 10 9 1 9 2 13 1 10 9 1 10 9 15 10 9 1 10 11 2 11 2 15 13 1 13 13 10 10 9 1 9 1 10 9 1 13 10 9 1 9 1 10 11 2
48 11 2 15 15 13 1 10 0 9 2 13 16 10 10 9 2 13 1 13 9 2 7 16 10 10 9 13 13 3 2 1 15 3 13 10 9 1 2 13 10 9 1 16 3 13 9 2 2
25 10 9 1 15 13 13 9 1 9 3 0 16 10 0 13 9 3 0 2 1 12 1 12 9 2
52 3 2 10 9 2 9 1 10 11 2 13 16 2 3 13 9 0 2 0 7 0 15 15 13 13 16 10 9 1 10 9 13 0 1 10 10 9 2 1 15 15 10 9 0 13 4 13 1 10 9 2 2
26 10 0 9 0 1 10 9 13 2 1 11 2 2 10 13 9 13 1 10 9 7 1 10 9 2 2
30 2 10 9 13 10 0 9 1 9 1 10 9 2 13 1 0 9 1 10 9 15 13 1 10 9 0 2 2 13 2
6 9 0 13 3 1 11
50 10 9 0 2 11 2 7 10 9 1 10 9 0 2 11 2 13 3 1 11 2 9 1 9 1 10 11 0 7 10 9 1 11 2 13 3 1 10 9 0 11 10 9 1 10 9 1 10 11 2
25 10 9 1 10 0 9 11 2 11 1 10 9 0 1 12 2 12 7 12 2 13 15 1 0 2
10 7 10 9 1 15 13 13 3 0 2
17 9 2 9 2 9 13 10 9 1 10 9 13 1 9 1 11 2
9 10 0 13 1 10 9 7 3 2
12 10 9 1 10 9 2 3 2 13 10 9 2
14 7 3 1 10 9 3 13 10 9 0 1 10 11 2
7 10 0 9 1 10 9 2
12 7 1 10 9 13 3 10 9 1 0 9 2
4 13 13 13 2
10 7 15 13 2 3 2 13 10 9 2
61 16 2 9 13 2 10 9 1 9 3 11 2 11 2 11 2 11 2 11 2 11 2 11 7 11 3 15 13 15 2 13 10 9 1 3 2 1 10 9 2 1 13 1 10 11 13 10 9 1 10 9 1 15 10 9 13 13 1 10 9 2
49 16 9 0 3 13 1 10 9 2 15 2 1 9 3 2 11 2 2 2 11 2 2 2 11 2 7 2 11 2 2 13 1 10 11 12 9 0 1 10 9 1 10 9 0 1 10 9 12 2
3 9 1 11
1 11
3 11 13 9
50 10 9 1 10 11 2 11 2 2 11 2 13 3 1 10 9 1 10 9 11 1 10 9 1 16 1 1 10 9 1 9 13 13 1 11 10 9 1 9 15 13 1 15 13 10 11 2 11 2 2
34 15 9 2 12 9 2 13 11 2 15 9 2 12 9 2 11 1 10 9 2 13 1 10 9 1 10 9 1 9 9 2 12 9 2
21 10 9 1 9 3 0 13 3 2 3 1 13 2 1 10 0 9 1 10 9 2
23 1 10 9 0 0 2 10 9 13 3 0 16 10 9 13 10 9 7 13 1 10 9 2
29 10 9 3 15 13 7 2 1 10 9 15 10 9 1 10 10 9 15 13 2 13 1 15 2 13 10 10 9 2
44 10 0 9 1 10 11 2 13 1 11 2 9 1 10 9 11 2 7 10 11 0 13 3 10 9 1 9 0 2 1 15 15 13 1 13 10 0 9 1 10 0 9 0 2
33 10 11 2 1 10 9 11 2 2 15 13 10 11 2 13 3 3 12 9 1 10 9 1 9 15 15 13 1 10 0 9 12 2
46 1 10 9 13 4 13 2 3 2 12 9 1 9 1 10 11 2 15 1 10 11 7 1 10 11 2 10 0 9 0 9 2 7 15 1 10 9 11 2 13 1 10 9 0 11 2
57 1 9 2 10 10 9 13 1 9 1 10 10 9 1 13 10 0 9 2 16 13 0 16 10 9 0 1 12 1 10 9 13 1 10 9 1 9 15 13 3 12 9 1 10 9 1 10 11 2 15 13 1 12 9 1 9 2
20 1 10 3 0 2 9 1 9 2 1 10 9 15 1 10 11 13 10 9 2
10 13 15 15 13 10 9 1 10 9 2
27 13 15 15 13 10 9 2 7 3 10 9 7 9 7 9 2 10 9 1 9 2 10 9 1 10 9 2
42 10 9 15 13 1 11 2 11 2 11 7 11 2 1 10 2 13 2 3 2 10 9 0 1 10 11 2 10 9 1 13 3 9 3 0 1 10 9 1 10 9 2
27 10 9 1 9 2 13 3 1 10 9 2 11 2 2 13 4 13 1 9 2 1 11 2 1 10 11 2
15 13 3 9 9 0 2 3 13 7 3 0 13 10 9 2
27 13 16 10 9 1 10 9 2 1 10 9 1 10 10 9 2 13 1 15 10 9 0 1 9 1 9 2
38 16 10 10 13 9 11 13 9 1 10 9 1 10 1 10 0 9 1 10 9 0 13 10 9 2 3 0 2 1 10 9 1 10 10 9 1 9 2
24 3 3 7 3 3 2 3 15 13 2 13 2 15 3 2 1 10 9 1 15 15 3 13 2
30 3 2 15 2 7 10 9 1 9 15 15 13 1 10 11 2 1 10 13 9 2 2 13 15 13 1 10 10 11 2
45 10 9 13 1 11 2 9 0 7 9 2 2 11 2 9 2 2 11 2 9 2 7 11 2 9 2 13 1 10 9 2 1 10 9 0 1 10 9 2 1 10 11 1 11 2
52 10 2 0 2 9 2 13 1 12 9 2 1 10 1 10 9 3 13 1 10 9 2 0 2 13 1 10 9 11 7 1 10 9 1 11 2 1 10 11 2 11 11 2 9 12 2 2 1 10 9 7 9
4 1 10 11 2
27 10 9 1 9 13 1 10 11 13 3 1 10 9 1 11 1 9 1 10 9 0 7 0 1 10 11 2
43 10 9 0 13 1 2 11 2 13 10 9 1 10 9 2 15 13 1 10 11 7 13 1 1 10 11 2 3 1 13 10 9 1 10 9 1 10 9 7 1 10 9 2
50 10 9 1 10 9 13 1 2 9 0 2 9 1 9 2 2 2 2 0 9 2 0 9 2 2 2 2 10 9 2 3 9 2 11 3 0 2 2 7 2 13 2 13 2 13 11 1 13 2 2
14 1 10 9 2 11 2 9 1 10 11 2 3 13 2
34 2 3 13 13 16 10 9 0 13 13 2 16 10 9 13 1 13 2 16 10 9 0 2 10 9 7 10 9 13 1 13 15 2 2
42 2 13 13 1 13 10 10 9 10 3 0 0 2 1 10 9 3 13 0 9 2 2 13 11 2 10 9 0 1 10 9 12 2 1 10 11 2 13 1 10 11 2
19 2 3 13 3 9 1 13 9 0 7 3 13 3 3 1 15 13 2 2
15 13 10 0 0 13 13 10 9 1 9 1 9 1 9 2
20 1 3 16 11 13 13 3 0 1 10 0 1 10 9 1 10 12 9 0 2
20 7 2 1 16 13 13 2 10 9 13 16 10 11 3 13 1 10 9 11 2
25 11 13 16 15 13 1 13 1 10 9 11 2 1 10 11 2 0 7 3 16 13 1 15 13 2
33 1 10 9 1 10 9 1 10 9 1 9 1 15 2 3 10 11 3 15 13 1 13 10 2 9 2 1 10 9 1 10 9 2
56 13 9 3 10 12 9 2 1 15 3 15 13 9 0 2 13 1 9 1 10 9 7 9 13 1 10 9 1 10 11 1 11 2 10 9 3 13 7 13 1 15 13 11 2 9 15 1 10 10 9 3 13 1 9 2 2
39 10 9 13 10 9 1 12 1 10 9 2 15 13 3 10 9 2 1 10 15 10 9 13 13 10 9 1 9 3 3 1 15 13 4 13 1 10 9 2
40 1 13 16 10 9 13 4 13 2 10 12 9 13 3 1 10 9 11 2 1 9 0 2 10 9 1 10 9 13 11 2 7 13 10 9 15 13 1 11 2
26 1 10 9 1 10 11 1 10 11 2 9 1 15 3 13 13 10 9 2 3 13 13 10 9 0 2
21 1 13 3 3 13 10 10 9 3 0 1 10 9 0 2 10 9 13 1 13 2
41 3 2 3 2 10 9 0 2 1 10 9 2 3 13 13 3 10 9 0 2 0 2 2 7 3 10 0 0 1 13 0 9 0 7 1 13 9 0 7 0 2
36 13 15 16 10 9 0 3 13 0 1 9 0 1 0 9 2 10 3 10 9 2 10 9 2 10 9 1 10 9 2 1 10 9 0 2 3
51 10 9 0 1 10 9 0 13 13 10 9 1 2 1 10 9 2 10 9 0 0 13 9 0 0 7 0 1 10 12 9 1 10 9 2 3 10 9 0 13 3 3 13 1 10 0 9 1 10 9 2
24 15 13 13 2 3 2 16 10 9 0 1 10 9 0 13 3 0 16 15 1 10 9 0 2
26 10 9 1 10 11 1 11 7 1 10 11 13 10 9 1 10 9 1 11 1 16 13 9 1 11 2
9 10 9 0 13 4 13 1 9 2
36 11 2 9 1 10 9 1 11 1 10 9 1 10 9 2 13 13 1 9 0 16 10 9 3 13 1 9 1 10 9 1 9 1 13 9 2
52 10 9 13 2 3 2 10 2 0 9 2 1 10 9 1 10 11 1 10 9 0 2 13 1 10 11 2 7 2 15 13 13 10 9 1 9 1 10 9 1 10 9 13 1 10 9 1 9 0 0 2 2
44 13 3 16 13 13 10 9 2 3 3 13 1 10 9 2 15 13 10 9 1 15 13 13 13 10 9 1 9 0 1 9 15 2 3 13 4 13 1 10 0 9 0 2 2
45 11 13 2 1 10 15 2 10 2 0 9 1 9 0 0 2 3 13 4 13 10 9 1 15 10 9 7 10 9 13 9 13 1 9 2 1 10 9 1 10 10 9 0 2 2
52 10 9 1 9 1 10 9 1 0 3 3 13 13 2 1 9 1 10 11 2 1 10 0 9 0 15 13 3 1 2 0 9 2 10 11 13 1 10 9 1 10 9 0 1 9 7 3 13 1 9 0 2
44 13 10 9 0 0 2 0 2 0 2 13 7 1 0 9 0 2 13 10 9 7 10 9 15 3 13 1 10 9 1 9 0 7 0 15 10 9 3 13 2 13 7 13 2
5 9 13 1 12 9
31 10 9 15 13 1 10 9 1 10 9 13 1 10 9 1 11 2 11 7 11 2 13 13 3 13 1 10 9 1 3 2
51 10 9 1 10 9 0 2 1 10 0 9 1 10 9 1 10 11 1 0 9 2 3 11 7 11 2 3 3 13 9 7 13 1 9 2 3 13 10 9 1 10 11 2 3 11 15 13 1 0 9 2
37 3 2 10 9 1 10 11 2 11 7 11 2 3 13 1 11 2 13 1 13 1 3 10 9 1 10 11 2 3 11 3 13 1 10 9 0 2
7 10 0 9 13 1 9 2
30 1 10 0 9 2 1 10 11 13 13 10 15 1 15 1 3 13 10 9 2 10 11 3 13 10 9 1 10 9 2
24 7 10 9 0 1 10 11 11 13 1 13 15 1 10 9 7 1 10 9 1 10 10 9 2
53 3 3 1 3 3 13 1 13 9 1 10 11 2 7 3 13 16 2 1 3 3 12 9 1 9 2 13 10 10 11 1 13 10 9 1 10 9 1 11 2 1 13 15 10 9 1 10 0 9 1 10 9 2
1 11
6 9 0 13 15 1 9
44 3 12 9 1 9 0 13 15 3 1 10 11 2 13 1 10 9 0 11 10 9 1 10 9 0 7 1 10 9 1 9 7 10 9 1 10 9 1 9 2 9 7 9 2
17 1 10 9 2 13 1 10 9 7 10 2 9 2 1 10 9 2
37 1 10 9 2 10 9 0 3 13 10 9 13 2 13 1 10 12 7 15 12 9 1 9 2 3 1 10 9 1 10 11 15 13 10 0 9 2
26 1 10 9 1 10 9 0 2 10 9 13 15 1 12 9 1 9 2 3 13 3 13 9 7 9 2
29 1 15 15 13 1 10 9 1 9 2 10 11 13 10 9 1 10 9 1 15 13 10 9 1 10 10 9 0 2
14 10 9 0 0 2 0 2 0 7 0 13 0 9 2
15 11 2 1 10 9 2 9 1 9 2 10 11 13 0 2
32 11 2 10 11 13 3 7 13 16 3 13 1 9 10 2 12 3 0 9 1 9 1 10 9 2 3 15 13 1 10 9 2
9 15 13 16 10 9 3 13 13 2
42 13 1 13 16 13 3 16 10 9 13 16 10 9 13 13 1 10 15 2 7 13 3 16 15 13 1 10 9 1 9 2 12 9 16 13 10 9 13 1 15 13 2
16 13 4 10 9 2 4 9 2 9 2 9 2 4 9 2 3
19 9 2 12 9 2 11 2 11 2 11 2 11 2 11 2 11 7 11 2
10 9 0 2 12 12 9 2 2 11 2
29 3 1 10 9 1 11 2 1 10 9 11 2 3 10 11 13 1 4 13 3 9 2 7 9 2 1 10 11 2
13 10 9 1 9 1 10 9 0 13 3 10 11 2
34 13 3 2 1 9 1 10 11 2 10 0 11 2 13 1 10 9 1 11 2 13 3 2 1 9 0 2 1 10 9 1 10 11 2
9 1 3 16 13 3 13 3 11 2
70 9 3 3 3 15 13 15 1 10 3 0 9 1 9 7 9 1 10 9 2 10 11 13 3 1 12 9 1 0 9 1 10 9 1 10 9 2 13 10 3 13 9 1 9 2 10 11 2 10 9 0 13 13 1 10 11 7 1 10 11 2 3 1 11 2 2 7 10 11 2
59 13 12 9 1 10 9 0 1 10 9 1 10 9 0 1 10 11 2 13 3 1 10 9 1 9 0 7 1 9 1 16 2 3 1 10 9 0 15 13 1 4 13 1 10 9 2 10 9 13 13 1 10 9 15 10 10 9 13 2
34 3 3 13 10 9 0 2 10 9 13 10 9 1 10 11 2 7 10 9 1 9 13 10 9 0 1 10 11 2 16 10 9 13 2
8 2 9 1 10 11 1 10 11
7 9 1 10 11 1 10 11
10 9 1 10 11 1 10 11 2 11 2
14 10 0 9 13 10 9 3 9 0 1 10 12 9 2
56 13 2 3 2 10 9 1 10 11 2 1 10 9 0 7 0 2 10 9 0 1 10 9 0 7 2 3 2 10 9 1 10 11 1 10 9 1 9 1 10 11 1 10 9 0 7 10 9 0 7 0 1 10 9 0 2
21 1 10 9 2 13 11 2 11 2 11 2 11 2 11 2 11 2 11 7 11 2
34 3 2 10 0 9 13 13 1 10 9 3 0 1 10 9 1 15 15 13 11 2 1 10 9 1 10 10 9 7 1 10 10 9 2
27 1 13 1 10 9 0 2 15 13 10 11 2 2 13 1 10 9 9 3 11 2 11 2 11 7 11 2
22 11 2 11 7 11 13 1 9 0 2 7 10 9 11 13 10 9 1 10 9 0 2
36 1 10 9 0 1 10 0 9 10 0 13 3 13 10 10 9 2 3 1 10 9 0 1 11 7 11 7 10 0 9 15 11 13 1 11 2
18 10 9 2 13 2 3 10 9 9 16 11 13 1 13 15 1 11 2
21 10 11 13 1 13 1 10 9 2 3 11 13 1 10 9 10 9 13 1 11 2
20 3 2 3 13 16 10 9 13 13 1 10 9 0 2 13 10 9 1 9 2
27 13 1 13 1 13 11 2 10 9 11 13 13 1 10 9 0 7 13 10 0 9 1 10 9 1 11 2
17 10 9 0 13 2 3 10 0 9 0 13 3 1 10 9 0 2
7 3 10 9 1 10 9 2
56 10 9 1 12 9 1 9 2 3 12 9 1 9 1 10 9 0 2 13 1 10 9 0 1 10 9 1 12 2 9 2 0 2 13 0 1 10 9 15 10 9 1 11 2 1 10 11 2 11 2 2 13 1 10 9 2
84 13 1 9 3 13 1 9 13 1 10 9 0 1 10 9 12 7 10 2 9 0 2 13 1 9 1 10 9 0 1 10 3 0 9 1 11 2 10 9 13 13 10 9 1 10 9 0 2 1 10 9 15 13 13 10 9 0 7 2 1 9 1 10 9 0 2 13 0 9 2 15 1 10 9 7 1 10 9 2 1 10 10 9 2
76 1 15 2 0 1 15 13 1 10 10 9 2 10 9 2 1 10 1 3 13 2 9 11 2 2 13 13 10 9 1 10 0 9 2 3 0 2 13 1 10 9 7 1 15 13 1 10 9 16 10 11 13 10 10 9 2 3 0 7 2 3 2 13 1 10 9 0 2 15 15 10 9 13 1 9 2
50 13 2 3 2 10 9 13 1 10 9 0 11 2 15 13 2 0 2 10 9 1 11 2 2 16 15 13 15 2 10 9 13 1 15 2 13 10 10 9 2 2 11 13 10 10 9 1 10 9 2
22 2 16 15 13 10 9 1 13 10 9 2 13 16 13 13 10 0 9 2 2 13 2
13 9 1 9 13 2 1 9 1 9 2 10 9 2
35 13 1 10 9 11 1 10 9 1 12 2 10 9 13 13 0 2 1 10 9 2 10 9 1 10 9 1 10 9 2 13 15 1 9 2
45 13 10 9 12 9 1 13 9 2 11 2 9 2 2 11 2 9 2 2 11 2 9 2 2 11 1 10 9 2 9 2 2 11 2 9 2 7 11 1 10 9 2 9 2 2
28 3 7 9 2 1 10 9 2 10 9 0 1 13 2 1 9 2 10 9 7 9 1 10 9 0 3 0 2
7 1 10 9 1 10 11 2
9 15 15 13 9 13 13 3 3 2
52 1 10 12 9 2 13 4 13 2 11 2 2 9 1 10 9 1 11 2 2 9 1 9 0 3 9 1 11 2 11 2 11 7 11 13 2 13 2 1 9 13 1 9 0 1 10 11 2 11 7 11 2
14 10 9 0 13 1 11 7 10 9 7 9 1 11 2
18 1 15 13 15 2 1 9 2 10 9 2 9 11 2 11 7 11 2
23 10 9 13 9 1 10 10 9 7 1 10 9 0 2 12 7 12 2 3 1 10 9 2
15 10 11 13 10 9 0 1 10 0 9 1 10 9 0 2
12 10 9 3 13 3 1 10 9 1 10 9 2
27 11 2 1 10 9 2 13 10 9 1 10 11 2 13 10 0 9 15 10 9 0 13 1 10 10 9 2
31 7 10 9 1 11 13 16 13 3 1 13 1 9 1 11 15 2 1 9 1 11 7 11 2 13 10 9 1 10 9 2
15 11 13 3 12 9 10 13 1 10 9 1 10 9 0 2
34 10 9 1 11 13 10 12 9 3 7 3 1 12 9 1 10 9 10 11 13 1 10 9 1 10 9 2 1 9 1 10 9 11 2
52 1 10 10 9 1 10 2 9 2 2 9 1 3 12 9 1 10 11 1 11 2 12 1 10 11 2 2 3 10 11 1 11 13 4 13 10 9 0 13 1 11 7 13 13 1 10 13 11 2 1 12 2
18 9 3 1 3 12 9 1 10 11 2 3 1 12 2 1 10 11 2
48 3 2 1 10 9 1 10 0 11 2 13 1 10 9 1 10 9 1 10 9 7 10 9 15 15 13 1 10 9 2 13 15 10 9 0 1 10 9 1 0 9 13 13 1 10 9 11 2
32 13 15 1 10 11 1 11 2 13 1 10 11 7 13 1 10 9 11 2 13 1 10 9 0 2 11 2 1 10 9 0 2
28 10 9 1 11 1 13 10 9 1 2 11 2 2 13 1 9 2 1 10 9 0 1 9 0 1 10 9 2
20 1 10 9 2 13 3 10 9 1 9 0 13 1 11 2 10 0 9 0 2
11 13 13 10 9 1 9 13 1 9 0 2
19 3 2 13 10 9 1 13 1 13 1 10 9 15 13 1 10 9 0 2
19 13 10 9 1 9 0 7 10 9 15 15 13 13 10 9 13 1 11 2
14 12 9 0 1 10 10 9 13 2 3 13 12 9 2
14 13 15 1 10 9 1 9 11 2 15 13 1 11 2
28 13 9 7 15 13 10 9 1 10 9 13 13 1 10 9 0 7 0 1 10 9 2 16 3 1 15 9 2
70 3 10 9 13 1 13 1 10 9 1 10 11 7 10 9 1 10 9 1 11 13 9 0 1 10 9 1 9 13 2 13 15 15 10 0 9 0 2 0 7 2 9 2 2 13 2 15 15 13 1 10 9 13 2 3 16 15 13 1 10 9 7 1 10 9 13 1 10 9 2
52 10 9 13 15 3 1 15 7 2 3 15 13 10 9 7 13 13 15 1 1 10 9 0 2 13 1 13 15 10 9 13 2 10 10 9 0 2 15 15 13 10 9 1 10 11 7 1 10 9 3 0 2
40 13 15 10 9 1 11 2 3 13 10 9 1 10 9 1 13 9 7 1 13 2 1 10 9 2 10 9 1 9 0 1 10 9 2 1 10 9 1 9 2
18 7 10 9 13 15 3 2 13 10 9 1 13 1 10 9 1 15 2
24 13 15 3 2 1 10 9 1 10 9 2 13 3 1 10 11 1 10 9 15 13 1 11 2
44 13 1 10 9 1 11 7 1 10 11 2 1 10 9 1 11 2 3 10 9 1 10 9 13 9 1 9 13 2 13 10 0 9 1 10 11 1 11 2 3 15 13 9 2
17 10 9 15 15 13 13 15 1 10 11 1 10 9 1 10 9 2
34 10 10 9 0 1 10 9 1 11 2 3 2 1 10 9 15 15 13 1 10 9 2 1 15 13 9 2 1 16 15 3 15 13 2
22 3 2 10 0 9 1 9 1 10 9 2 1 10 9 7 1 10 9 1 10 9 2
53 10 9 0 1 10 0 9 1 10 9 2 3 10 9 1 10 9 15 13 13 1 9 10 9 13 1 10 9 1 10 9 7 3 15 13 13 1 10 10 9 2 15 3 3 15 13 1 10 9 13 7 0 2
10 3 2 3 13 13 15 7 13 15 2
19 3 2 10 9 13 13 10 10 9 1 10 9 0 7 13 1 10 9 2
17 2 7 10 9 13 15 1 3 13 0 2 2 2 13 15 3 2
4 3 10 9 0
41 1 10 9 1 13 9 1 15 10 9 13 13 1 10 0 9 2 13 16 3 13 3 10 9 15 3 13 13 1 10 9 0 2 9 1 9 0 7 9 0 2
26 10 9 13 3 0 16 3 10 10 9 13 13 7 13 2 3 2 1 10 9 1 10 9 1 9 2
16 13 15 1 10 0 9 1 10 9 1 2 10 13 9 2 2
35 1 10 9 1 10 0 2 13 12 9 1 15 13 1 10 9 7 3 13 10 0 9 15 3 15 13 1 10 9 1 10 10 9 0 2
31 13 3 0 1 3 10 9 2 7 3 15 13 10 9 1 10 9 13 13 1 10 9 1 9 1 10 0 9 3 0 2
11 13 10 9 2 10 9 3 13 13 0 2
16 3 3 2 1 15 15 13 13 3 13 2 13 3 12 9 2
31 3 3 16 10 9 3 1 10 10 9 15 1 10 9 13 13 10 9 1 10 10 9 3 15 13 9 1 10 10 9 2
23 1 10 9 2 10 10 9 13 1 10 9 1 10 9 2 3 13 13 12 1 12 9 2
28 16 13 4 13 9 3 1 10 10 9 7 16 13 10 9 15 13 1 13 10 9 1 9 1 10 9 0 2
5 9 0 3 1 9
25 10 9 0 11 13 12 1 10 9 13 1 10 11 1 10 9 2 11 2 2 15 13 1 11 2
32 3 13 10 9 1 10 9 1 10 9 0 7 10 9 13 1 10 9 1 10 9 2 10 9 0 7 10 9 1 10 9 2
15 10 0 9 2 13 1 9 2 13 12 9 1 0 9 2
39 1 11 2 10 11 13 10 11 2 9 15 13 13 1 10 9 1 13 1 10 9 0 2 12 9 7 10 9 2 2 3 10 9 13 13 10 9 0 2
26 1 10 10 9 2 10 11 13 3 1 10 0 11 2 3 1 0 9 2 1 12 9 1 10 9 2
16 10 11 3 13 0 9 2 16 13 1 10 11 1 10 11 2
24 3 2 11 2 11 2 11 7 11 2 10 9 2 13 10 9 13 7 13 1 10 9 13 2
13 10 9 13 13 7 0 2 10 9 0 7 0 2
11 13 10 9 1 13 2 13 13 7 0 2
19 1 10 9 13 9 1 9 2 10 9 0 1 9 7 10 9 1 9 2
27 1 1 10 9 0 1 9 2 10 9 13 15 10 9 15 13 7 13 2 2 10 9 2 1 15 2 2
5 12 9 1 10 9
60 1 11 2 10 9 1 10 9 13 0 9 1 10 9 1 15 0 13 2 1 9 1 10 11 2 15 13 1 10 0 9 2 7 1 10 11 2 15 2 1 13 2 13 1 10 0 9 1 10 11 7 1 10 11 7 3 13 10 9 2
51 11 7 11 13 3 10 0 9 2 15 1 12 9 2 12 9 13 7 12 13 2 13 1 10 11 2 3 1 12 9 2 1 10 11 2 1 12 2 10 10 9 2 2 7 1 10 11 2 1 12 2
28 10 0 9 13 1 15 9 2 1 10 9 1 10 11 1 10 11 2 12 2 2 1 10 9 13 1 11 2
38 1 10 9 2 10 11 13 13 1 10 9 1 10 11 2 12 2 2 13 10 0 9 1 10 9 2 3 10 11 13 7 13 10 11 2 12 2 2
31 1 10 9 1 10 11 2 10 11 3 13 1 10 9 1 9 2 15 13 10 9 1 11 1 15 13 1 10 0 9 2
10 11 3 13 9 1 10 9 1 10 9
8 11 7 11 13 3 1 10 9
78 10 9 1 16 10 9 1 2 11 2 13 10 9 13 13 13 15 2 3 2 1 10 9 1 10 2 11 2 15 13 3 1 2 9 2 2 1 10 9 2 15 13 1 13 1 15 2 2 7 15 1 10 9 1 9 1 9 1 10 9 13 2 2 9 11 2 10 10 9 13 10 10 9 1 10 9 2 2
12 13 15 2 3 2 16 13 15 13 10 9 2
16 7 3 2 11 7 11 13 2 3 2 10 9 1 10 9 2
41 1 10 9 1 11 7 1 11 2 13 3 10 9 1 10 9 1 11 2 11 7 11 13 10 0 13 1 10 2 9 2 2 9 1 11 2 13 15 1 11 2
17 7 1 13 10 9 2 2 13 10 9 15 3 15 13 13 2 2
11 11 2 1 10 9 13 1 2 9 2 2
6 0 2 10 9 13 2
8 3 1 15 3 10 11 13 2
15 3 13 10 9 1 9 1 10 0 9 0 1 10 9 2
12 13 15 13 13 10 9 1 10 9 3 13 2
45 7 13 13 10 9 0 1 10 9 2 1 13 3 13 1 10 9 15 2 3 2 1 10 11 15 13 9 2 2 3 3 1 9 3 13 10 9 13 9 2 3 2 1 11 2
49 13 1 10 9 7 1 10 9 1 10 9 1 10 0 9 1 10 9 0 2 1 10 9 9 1 9 7 9 2 13 9 1 11 13 3 13 9 1 15 15 3 3 13 9 1 13 10 9 2
25 10 9 1 10 2 11 2 13 3 0 7 0 1 13 0 7 2 3 2 13 10 9 0 0 2
42 16 13 1 10 12 9 10 9 3 0 1 10 9 2 10 9 1 10 11 13 10 9 15 13 1 10 9 1 10 9 0 3 1 1 10 9 1 9 1 10 9 2
53 1 10 0 9 1 10 12 0 9 2 13 15 1 2 10 9 0 1 10 9 1 13 3 10 9 0 1 10 9 1 13 0 9 7 0 9 2 1 10 9 1 10 9 0 1 10 11 7 1 10 11 2 2
46 1 12 9 1 9 1 10 11 2 12 1 15 1 10 9 1 11 2 13 13 15 3 10 9 0 1 9 0 1 10 11 2 11 2 2 13 1 12 1 13 10 9 1 10 9 2
35 10 9 1 10 9 13 16 10 11 2 1 10 9 1 11 2 13 13 1 12 1 12 9 1 10 9 1 10 9 1 9 1 10 11 2
42 7 10 9 13 1 10 9 10 9 1 10 9 0 2 16 10 11 0 1 13 1 10 0 9 13 10 9 1 10 9 1 10 9 15 13 3 12 9 1 10 9 2
8 9 1 9 13 12 9 1 12
5 11 13 9 1 9
57 10 9 1 9 1 9 0 7 1 10 9 1 10 0 9 2 10 9 1 9 3 0 1 10 9 3 1 15 7 1 10 9 1 10 10 9 3 10 9 1 9 1 9 1 9 7 1 9 13 10 12 0 9 1 10 11 2
3 9 1 9
2 9 0
6 10 11 13 1 0 2
40 3 12 9 1 13 13 10 11 1 9 2 13 1 10 11 2 13 1 10 9 1 10 2 9 2 12 9 15 13 1 10 9 1 10 9 2 11 7 11 2
27 10 11 13 10 10 0 11 1 15 13 10 11 2 1 12 2 1 10 9 1 10 9 13 1 10 11 2
35 1 10 9 1 10 9 2 9 1 10 11 13 9 7 9 1 10 9 1 9 2 3 13 11 2 9 1 10 11 2 7 11 2 9 2
49 11 2 9 1 10 11 2 1 10 9 1 10 2 11 2 2 13 16 3 13 2 1 15 15 1 15 15 13 2 9 0 1 15 13 7 13 16 10 11 1 11 13 10 9 3 0 1 11 2
33 10 9 2 1 9 0 2 1 3 12 9 1 0 2 13 13 3 11 2 9 1 10 9 2 3 13 13 10 9 1 9 0 2
47 10 9 13 1 10 9 13 10 9 3 13 1 10 9 1 11 2 7 3 3 2 1 10 9 1 10 9 11 7 11 2 13 1 9 1 10 11 2 15 13 1 10 2 9 0 2 2
37 1 10 10 9 1 15 13 13 10 9 2 10 9 2 1 9 1 10 11 2 13 3 13 9 0 15 13 3 1 13 9 1 9 7 9 0 2
44 1 10 9 11 2 1 9 1 10 11 2 10 9 0 2 13 13 10 9 0 1 10 0 2 11 2 7 13 10 9 0 1 11 1 10 9 1 10 9 1 10 9 2 2
17 10 9 13 3 13 10 9 7 13 10 10 9 1 9 7 9 2
34 3 2 3 10 9 0 11 2 11 7 11 13 1 10 9 2 2 10 10 9 13 11 2 3 13 11 2 2 2 13 10 9 3 2
6 7 11 13 10 9 2
13 2 13 10 9 0 15 3 3 13 13 3 2 2
21 10 0 9 13 10 2 9 2 11 15 13 0 9 1 10 9 1 10 11 0 2
68 13 1 10 9 1 12 1 12 9 0 2 10 0 1 15 1 11 2 1 11 2 11 2 0 11 2 13 13 1 13 0 10 9 3 1 13 13 11 2 9 1 9 9 2 2 12 1 10 9 1 0 9 10 9 1 10 9 13 2 9 2 9 2 12 2 12 2 2
37 2 3 13 13 0 9 3 2 7 3 13 1 13 10 9 3 13 15 3 0 2 2 13 10 9 1 10 9 1 12 2 12 2 12 7 12 2
24 10 9 13 15 2 7 3 13 15 1 13 1 10 9 0 15 13 1 10 9 1 10 9 2
20 10 9 13 15 0 1 10 9 0 7 13 9 1 10 9 13 1 10 9 2
40 11 2 1 10 11 2 13 16 2 1 2 9 2 2 10 9 13 7 10 9 1 10 9 0 13 10 9 3 13 1 10 9 1 10 9 0 1 10 9 2
22 10 9 13 1 10 9 1 12 7 10 9 13 1 10 9 1 10 0 9 1 9 2
29 10 9 1 9 1 11 13 3 10 9 1 10 11 2 15 13 1 13 13 1 12 9 1 9 0 1 10 9 2
24 10 11 13 10 9 13 7 10 9 13 13 15 1 13 10 9 0 1 10 9 1 9 13 2
51 10 11 2 11 2 13 1 12 15 1 0 9 1 9 1 9 0 2 13 10 11 2 11 2 2 15 13 10 9 1 10 9 13 10 2 9 2 2 3 3 1 10 9 2 1 10 9 1 10 11 2
27 10 9 15 13 13 3 0 16 10 9 1 10 9 1 10 11 13 13 0 1 10 9 0 1 10 9 2
37 3 1 10 9 3 15 13 10 9 1 10 9 1 10 2 3 2 2 0 1 10 9 15 13 10 9 13 1 10 9 1 10 9 1 10 9 2
22 7 3 3 1 10 9 3 13 10 9 1 10 15 13 13 10 9 1 10 12 9 2
14 1 10 12 9 1 10 9 2 10 9 13 10 15 2
47 16 15 2 3 2 1 10 0 9 1 10 9 13 0 1 10 3 0 1 10 12 9 13 2 15 13 2 3 1 9 2 10 9 1 10 9 13 1 10 9 1 10 11 7 10 11 2
49 2 16 15 13 1 13 2 10 9 13 13 1 12 7 12 9 2 2 13 11 2 9 1 10 9 1 10 11 1 10 11 2 15 13 1 15 2 9 0 2 1 10 2 3 2 1 10 11 2
10 12 9 2 10 9 2 10 9 1 9
6 10 9 1 15 15 13
9 13 15 1 11 2 11 7 11 2
6 12 9 2 10 9 2
24 13 15 1 10 9 15 10 0 13 2 2 11 2 2 2 15 10 0 13 7 10 0 13 2
33 13 15 1 10 9 0 2 13 1 10 9 13 2 10 9 11 2 7 1 10 9 3 10 0 2 10 9 1 11 2 15 13 2
11 1 10 9 2 13 15 10 9 1 9 2
39 10 0 9 1 9 2 15 15 10 11 13 3 1 10 9 2 1 10 11 2 7 1 10 15 15 13 2 3 3 16 2 0 9 2 13 1 10 9 2
13 9 2 0 2 1 0 9 7 0 9 1 9 2
22 9 2 3 12 11 2 13 2 1 10 9 3 13 2 1 9 1 10 12 0 9 2
21 2 13 10 0 9 15 15 13 0 1 13 10 9 1 9 1 10 9 0 0 2
12 11 13 3 0 1 10 9 7 1 10 9 2
16 11 13 1 10 9 1 9 1 10 9 1 10 9 0 13 2
10 10 11 13 1 13 15 1 10 9 2
8 1 11 2 3 13 13 15 2
7 11 2 9 0 1 10 11
3 2 11 2
44 2 3 16 13 10 9 0 2 3 1 10 9 15 13 1 10 9 0 1 10 0 12 9 7 2 1 0 9 2 16 10 11 13 3 3 13 1 10 9 16 1 10 9 2
26 1 11 3 13 9 13 10 9 16 15 13 1 10 9 1 10 10 9 1 13 2 10 9 0 2 2
40 3 13 2 3 2 10 9 1 10 9 1 9 1 13 16 2 3 13 13 10 0 9 1 10 9 0 1 13 7 1 10 9 0 1 9 1 10 9 2 2
30 11 13 16 10 9 1 11 2 13 1 0 9 1 10 9 2 3 13 10 9 1 2 10 9 0 1 10 11 2 2
38 1 10 2 11 2 2 9 0 1 10 9 2 10 9 13 13 15 2 13 1 10 10 9 1 10 15 13 13 2 10 9 1 9 1 10 11 2 2
80 1 9 1 10 11 2 12 1 10 9 1 10 2 11 2 13 9 1 10 9 1 9 1 10 9 13 1 12 1 9 0 2 13 1 10 9 1 10 9 15 13 13 1 10 11 10 9 0 1 11 2 10 9 1 10 9 2 11 2 7 11 2 0 1 10 11 2 7 15 13 13 1 9 2 16 13 3 1 9 2
52 10 10 9 13 16 15 13 1 10 9 13 13 1 13 16 13 10 9 1 9 1 10 9 1 11 2 15 13 13 13 1 10 9 2 3 10 2 9 13 1 10 9 13 13 1 9 13 1 10 9 2 2
3 9 1 11
37 1 9 1 11 2 10 11 2 11 2 13 15 13 1 10 9 1 9 1 10 9 0 2 0 10 9 1 0 9 2 3 1 9 1 9 0 2
32 1 13 2 10 11 13 9 10 9 1 10 9 1 10 9 2 9 3 1 9 7 9 1 10 9 0 2 3 1 10 9 2
47 10 9 1 11 13 1 10 9 1 9 3 13 3 9 1 9 2 10 9 2 13 1 9 2 3 13 4 13 1 9 2 1 3 12 9 2 15 13 9 1 10 9 0 1 15 13 2
19 7 1 9 1 9 1 10 9 7 10 9 1 10 9 13 10 9 0 2
41 3 2 13 3 10 11 2 1 10 2 9 2 13 1 10 9 1 10 9 0 13 15 10 9 2 13 9 7 9 0 15 13 13 1 9 7 3 1 10 9 2
17 13 15 1 10 9 7 2 3 2 10 10 9 13 13 1 9 2
3 11 13 9
24 3 2 11 13 1 10 9 10 9 1 11 7 11 7 3 9 1 9 2 9 7 9 0 2
43 10 0 9 13 3 1 11 13 1 10 9 0 3 10 9 13 13 1 10 9 7 3 13 1 10 9 1 13 1 12 9 2 13 10 9 0 1 10 9 2 11 2 2
18 10 9 13 1 10 9 2 7 10 9 13 1 13 7 13 13 3 2
50 11 13 13 10 9 1 10 11 2 7 3 13 4 1 13 1 10 11 2 13 16 10 11 2 3 13 3 10 9 2 7 16 13 10 9 7 1 15 16 10 9 2 13 1 13 10 9 0 2 2
61 10 11 13 16 13 1 10 9 0 7 16 13 10 9 13 1 13 10 9 1 10 9 2 13 3 0 1 0 2 16 16 13 13 1 10 9 1 10 9 0 9 13 3 13 3 10 9 0 2 1 10 9 1 10 9 1 10 11 2 11 2
35 10 9 3 13 1 10 9 2 9 2 1 10 9 2 11 2 2 13 1 10 11 1 11 7 10 11 2 3 1 10 11 2 11 2 2
34 7 10 9 13 0 1 12 1 9 7 13 0 16 2 1 10 10 9 1 9 1 10 9 2 0 9 1 10 9 13 1 13 15 2
17 2 15 13 0 2 13 10 0 9 2 15 3 13 16 13 2 2
15 11 2 12 9 2 13 1 10 9 1 10 9 2 3 2
26 1 10 9 2 13 1 10 9 1 10 9 1 10 2 11 2 2 15 13 1 10 9 1 10 9 2
5 7 3 15 13 2
9 2 13 10 9 7 10 9 0 2
7 13 13 1 13 11 2 2
11 10 0 9 13 1 10 0 9 1 11 2
17 2 10 9 13 15 15 13 10 9 13 3 0 16 10 9 2 2
25 10 9 13 2 3 1 10 9 1 11 2 1 10 9 1 10 0 9 1 11 2 2 11 2 2
60 11 13 16 11 3 13 9 1 13 10 10 9 1 1 10 0 9 2 15 13 13 2 3 13 10 9 1 10 9 13 1 10 9 2 7 1 1 15 13 10 0 9 1 10 9 2 10 9 2 10 9 1 10 9 2 3 2 10 9 2
24 10 9 2 13 1 12 2 13 10 9 1 10 0 9 2 1 15 10 9 13 13 10 9 2
48 9 2 0 9 2 2 9 2 2 9 0 2 11 2 2 9 2 2 9 0 2 2 9 2 2 13 15 1 10 9 15 2 1 10 9 7 10 9 2 13 13 1 10 0 9 1 9 2
4 11 7 11 13
48 10 11 13 13 1 13 1 10 11 13 1 9 13 10 9 0 15 13 10 12 9 2 1 10 9 0 1 9 1 9 2 16 10 9 0 3 13 10 10 9 0 1 10 9 1 12 9 2
58 10 9 1 11 2 11 2 13 13 10 9 1 11 2 7 13 16 10 11 13 1 13 13 10 9 1 10 12 9 2 1 15 1 10 9 1 9 2 9 2 9 7 9 0 1 10 9 1 10 9 2 9 0 2 9 7 9 2
28 10 9 1 10 9 1 10 9 0 0 13 13 1 11 1 10 0 9 2 3 1 10 9 1 10 9 0 2
5 11 13 9 1 9
23 1 11 1 12 1 9 2 11 13 1 11 2 3 12 9 2 13 15 3 1 10 11 2
33 1 10 9 1 10 13 9 13 13 1 10 9 0 1 10 0 9 1 10 11 2 1 10 11 2 1 13 13 10 9 1 9 2
17 9 0 13 16 10 0 13 13 10 9 1 10 9 1 10 9 2
26 1 10 9 2 11 13 9 7 16 13 13 9 2 13 3 10 10 9 1 10 9 3 1 10 9 2
22 0 2 13 10 9 9 2 11 2 2 13 13 0 7 16 13 10 9 1 10 9 2
27 10 9 3 13 13 1 10 9 1 10 11 15 15 13 1 9 0 1 10 11 2 11 7 1 10 11 2
17 10 9 1 10 9 13 1 10 10 9 1 10 11 2 11 2 2
34 3 1 10 11 2 10 11 13 13 0 10 9 13 1 10 11 7 13 10 9 1 10 9 1 10 9 1 10 9 1 10 10 11 2
21 10 9 13 16 10 11 13 12 9 2 12 0 2 0 2 7 15 0 2 13 2
29 10 0 9 13 4 13 1 10 11 2 1 10 11 2 1 12 9 7 13 15 1 13 13 1 10 9 1 11 2
40 13 1 9 1 9 2 11 13 10 9 13 1 10 9 1 9 2 15 3 13 1 10 9 1 10 0 13 3 12 9 2 1 10 9 0 1 15 13 0 2
30 12 9 3 3 2 10 11 13 10 9 7 13 10 9 1 10 9 1 10 9 1 10 11 2 1 15 13 13 3 2
6 9 1 10 9 0 9
38 10 11 13 2 1 12 2 10 9 0 9 1 12 12 9 1 9 2 12 12 9 1 9 2 2 15 13 10 9 1 12 9 1 10 9 1 12 2
47 10 9 2 11 2 13 3 16 2 1 10 9 13 2 10 9 0 13 10 9 0 1 12 12 9 1 9 2 3 12 12 9 1 9 2 2 13 10 9 1 12 9 1 10 9 0 2
25 10 9 13 10 9 1 12 9 2 15 13 1 12 12 9 1 9 2 12 12 9 1 9 2 2
31 10 0 9 0 1 10 9 0 13 4 13 1 12 2 1 10 9 1 12 12 9 1 9 2 12 12 9 1 9 2 2
4 9 1 10 11
20 10 11 13 10 9 1 10 9 0 1 10 9 1 9 1 10 9 0 11 2
53 10 0 9 2 10 9 0 9 11 2 13 1 10 0 9 10 0 9 1 10 9 2 15 13 10 9 1 9 1 10 9 1 10 12 9 1 9 2 3 12 9 1 9 2 7 10 9 1 10 9 1 9 2
24 10 11 13 3 13 10 9 1 10 0 9 1 10 9 0 13 1 10 9 0 0 2 11 2
42 13 15 3 10 9 2 1 10 9 2 1 10 0 9 1 10 9 1 9 1 10 9 0 11 2 10 9 0 13 1 3 12 9 1 9 2 3 12 12 9 2 2
8 3 10 9 1 9 13 3 2
6 7 2 3 2 13 2
23 13 10 9 1 10 11 11 1 15 13 10 9 1 10 9 1 9 13 1 10 0 11 2
42 2 3 2 7 13 15 1 10 9 3 0 2 13 0 16 15 13 10 0 9 1 10 9 0 1 10 9 2 13 15 10 9 1 10 9 7 10 9 1 10 9 2
33 3 2 7 13 15 1 10 9 3 0 2 13 1 13 16 13 13 10 9 0 1 10 11 1 10 9 1 10 9 9 0 2 2
55 16 10 9 2 11 2 15 13 1 9 7 9 2 1 11 7 1 10 11 2 1 10 9 1 10 9 7 1 10 9 1 10 11 2 3 10 11 15 13 13 1 9 1 13 10 9 1 9 1 10 0 9 1 9 2
59 1 10 9 2 10 9 15 15 13 1 13 3 10 9 1 9 0 3 10 9 1 9 7 10 9 0 1 15 15 13 2 9 2 2 13 13 10 9 0 1 10 0 11 2 3 1 10 9 13 13 1 10 9 1 11 1 10 11 2
38 10 9 0 13 1 10 11 2 1 10 9 2 1 11 2 1 10 11 2 1 10 9 1 10 11 2 11 2 11 2 11 2 11 2 11 7 11 2
26 13 1 10 11 2 1 10 9 2 10 12 0 9 7 13 10 12 9 7 11 3 13 1 10 9 2
20 3 2 3 2 3 1 0 9 9 3 10 9 7 10 9 13 1 10 9 2
42 11 13 1 11 2 11 2 2 15 3 13 10 9 0 1 12 9 2 11 2 11 2 12 9 2 2 11 2 11 2 12 9 2 7 11 2 11 2 12 9 2 2
36 3 13 10 11 0 2 9 2 2 13 10 11 2 11 2 11 2 11 2 11 2 11 2 11 7 11 2 1 10 9 0 1 13 10 9 2
29 10 9 0 0 2 1 10 9 2 13 1 10 9 1 10 0 9 1 11 2 1 10 11 2 1 9 7 9 2
18 10 9 0 13 1 10 0 9 2 7 1 10 9 13 0 10 11 2
35 11 13 1 11 2 11 2 12 9 2 2 11 2 0 2 12 9 2 2 11 2 11 2 12 9 2 7 11 2 11 2 12 9 2 2
23 10 0 9 1 10 9 0 13 10 9 1 10 9 0 2 13 1 12 9 2 1 11 2
36 2 13 16 13 13 10 9 1 10 9 1 10 9 11 2 2 13 1 10 9 1 9 1 10 9 11 2 9 1 10 9 2 13 10 11 2
17 2 13 16 13 4 1 13 10 9 1 9 1 10 0 9 2 2
21 1 10 9 2 11 13 2 2 9 1 10 1 10 0 9 7 10 0 9 2 2
42 3 3 1 10 9 1 10 11 15 10 11 13 4 13 1 12 9 1 10 9 2 1 12 9 1 9 15 2 15 13 13 1 10 9 11 2 11 2 11 7 11 2
18 10 0 2 10 3 0 1 10 9 2 13 13 3 1 10 9 13 2
64 16 15 13 3 13 13 2 13 15 10 9 1 12 9 1 9 1 10 11 2 10 11 7 10 11 2 7 10 9 1 12 0 9 13 1 13 3 10 10 9 1 9 2 10 11 2 11 2 7 10 11 2 11 2 2 15 1 10 9 1 10 9 0 2
40 10 9 1 10 12 9 13 3 1 15 13 3 10 9 0 1 10 9 13 1 13 10 9 1 9 2 13 10 9 13 3 9 1 10 0 9 1 10 9 2
55 7 10 9 1 10 9 1 11 15 13 1 10 9 0 2 1 10 9 1 13 9 3 10 10 9 15 13 13 10 9 3 2 3 13 1 3 0 2 3 16 10 9 13 10 0 9 1 10 9 1 10 9 1 9 2
53 1 10 9 13 2 10 11 11 2 15 13 3 3 1 10 9 0 1 9 2 13 10 9 0 1 10 9 0 3 13 1 10 11 2 3 10 11 15 13 2 1 10 9 0 2 1 10 9 1 10 9 0 2
53 1 10 9 1 10 9 2 11 2 10 9 2 15 13 13 3 1 10 9 13 1 10 11 7 1 10 11 2 13 1 10 9 2 13 10 9 1 9 1 10 0 9 7 13 16 10 9 13 0 1 9 2 2
12 10 9 11 13 1 10 9 2 1 10 11 2
5 10 9 13 3 2
5 9 2 12 1 9
10 9 0 1 10 9 2 1 10 11 2
9 13 1 10 9 12 1 10 9 2
41 3 13 10 9 2 9 0 2 9 1 10 9 2 0 2 9 2 9 2 9 1 9 2 9 2 3 2 2 1 15 10 9 13 3 0 7 10 9 3 0 2
28 3 1 15 3 1 10 9 2 0 7 0 2 13 10 9 0 2 7 3 12 2 1 10 9 7 10 9 2
23 15 10 2 1 10 9 0 1 12 2 3 13 1 10 9 3 10 9 2 3 10 9 2
29 10 9 0 3 13 3 16 10 9 1 10 9 1 10 9 2 1 9 3 13 1 10 9 0 7 1 10 9 2
38 13 0 16 10 9 0 13 3 9 1 13 12 3 13 9 1 10 9 0 2 3 1 10 9 15 13 1 4 1 13 1 10 9 1 10 9 0 2
67 1 10 10 9 1 9 1 11 3 13 13 12 3 9 1 13 2 3 13 10 0 9 1 10 9 1 9 1 11 2 3 10 1 10 9 0 2 1 10 9 0 1 10 0 11 2 15 3 13 10 9 1 13 1 13 15 3 0 1 10 9 1 9 1 10 9 2
22 7 13 13 1 13 16 10 9 1 9 13 13 3 1 13 10 0 9 1 9 0 2
46 16 10 9 1 10 11 13 4 13 1 10 9 1 10 9 1 10 9 2 3 10 9 1 10 0 9 1 11 15 15 13 0 2 13 13 13 10 9 0 1 10 9 1 10 11 2
26 13 15 16 1 15 15 13 1 13 9 1 9 7 1 3 13 3 7 10 9 1 9 7 10 9 2
28 1 10 9 2 13 16 10 0 9 1 9 1 10 11 2 2 11 2 2 11 2 12 2 13 10 0 9 2
82 16 2 1 1 15 15 13 2 2 10 11 13 13 10 9 0 1 10 15 13 13 1 10 9 1 13 10 9 0 1 10 9 7 1 10 9 7 10 9 15 15 13 1 9 1 10 9 2 16 13 9 0 0 2 1 3 13 13 1 10 9 13 7 1 15 13 9 13 1 15 13 2 2 9 2 2 3 13 13 10 9 2
29 10 0 9 1 10 11 1 10 9 13 13 12 9 2 1 10 9 1 10 11 2 13 13 1 10 9 3 0 2
16 2 1 10 9 10 9 13 4 13 3 9 1 9 0 2 2
31 15 13 10 9 0 15 3 13 4 13 1 15 2 13 15 13 10 9 1 10 9 1 10 9 1 10 11 7 1 15 2
90 1 10 9 1 9 7 9 1 10 9 2 13 9 1 10 9 2 10 9 1 10 11 13 10 9 13 1 10 9 1 10 9 1 13 1 13 9 0 2 13 3 13 2 1 7 1 10 9 1 10 9 1 10 11 2 2 15 15 13 1 2 9 2 2 2 7 13 13 10 9 0 1 10 9 1 10 9 3 0 1 10 9 15 13 10 9 1 10 9 2
5 9 1 9 1 11
3 9 1 11
26 10 9 0 1 9 1 10 11 13 10 11 1 10 9 1 11 2 11 7 1 10 11 1 10 11 2
72 13 1 10 11 2 10 9 1 10 9 1 10 11 2 1 10 11 2 1 10 9 1 10 11 2 2 1 10 11 7 10 9 0 1 10 11 13 0 1 13 16 10 9 13 13 1 10 11 2 11 2 13 1 10 0 9 9 2 13 3 15 3 15 13 10 9 1 2 9 0 2 2
47 3 2 10 10 9 0 13 13 2 1 10 0 9 1 10 11 2 9 2 1 13 10 9 1 16 13 13 10 9 1 13 1 10 11 7 1 10 9 1 9 1 10 11 2 11 2 2
15 9 1 10 11 13 13 9 1 9 1 10 9 1 10 9
2 11 0
20 11 13 10 0 9 1 10 9 1 9 1 9 0 15 10 11 13 1 13 2
65 1 15 13 1 10 11 2 7 13 1 10 9 1 10 9 1 10 9 0 2 10 9 0 13 3 10 10 9 1 10 9 2 9 13 1 2 10 9 7 10 9 1 9 7 9 1 10 9 1 10 9 2 7 1 10 2 9 1 10 9 7 10 9 2 2
31 3 3 15 13 13 1 10 9 1 13 12 9 7 10 9 1 9 2 3 13 13 1 10 9 1 16 10 9 13 13 2
26 13 15 2 1 7 1 9 2 1 13 4 2 7 3 4 2 1 10 10 9 13 1 10 9 13 2
17 13 10 9 2 7 10 9 2 2 1 9 15 10 9 13 13 2
4 7 3 13 2
50 3 2 13 15 16 2 1 9 0 2 10 9 1 10 9 2 3 10 9 0 2 15 15 13 13 1 10 3 0 2 13 1 4 13 2 7 13 1 10 0 9 2 1 16 10 0 13 13 3 2
8 13 10 9 2 7 3 13 2
42 10 9 13 13 1 10 9 0 1 10 11 2 11 2 7 1 10 11 2 11 2 2 7 13 15 1 10 9 1 9 1 10 9 1 9 1 10 9 0 1 11 2
1 11
3 9 13 0
10 11 2 11 7 11 7 11 2 11 2
26 3 2 1 11 2 13 15 10 9 1 10 9 1 10 9 1 10 11 2 1 13 9 12 1 9 2
63 10 9 1 9 15 13 10 12 0 3 1 9 2 7 15 13 10 11 1 13 10 9 15 15 13 2 1 11 2 12 9 1 10 2 11 2 2 3 10 11 13 13 1 10 11 13 15 0 9 1 15 13 10 9 1 10 2 11 2 1 10 9 2
9 3 2 1 10 9 15 13 0 2
47 3 3 1 10 9 0 15 13 13 10 9 1 10 9 15 13 11 1 10 0 11 2 10 9 13 10 10 9 1 11 1 10 0 2 13 10 9 1 9 3 0 2 3 15 1 11 2
59 3 3 0 16 10 9 13 1 10 9 0 13 13 16 10 9 0 3 13 2 3 16 1 9 7 9 1 15 13 15 3 15 13 1 13 1 10 9 1 15 15 13 1 9 0 7 1 15 10 9 15 13 1 9 0 1 15 10 2
19 10 9 13 4 1 4 13 3 2 3 1 9 15 13 7 13 9 0 2
31 13 9 1 15 10 9 1 10 0 9 0 1 9 1 12 2 10 0 9 1 10 9 1 10 9 1 9 1 10 9 2
30 13 1 10 9 0 2 1 0 9 0 2 10 11 13 3 13 2 13 10 10 9 1 10 0 0 1 10 9 0 2
53 1 3 2 13 3 13 7 13 7 2 3 3 13 2 13 10 9 1 9 1 9 7 9 13 1 9 1 10 9 0 7 0 2 13 3 1 10 9 13 1 10 0 9 7 10 2 9 2 2 13 10 11 2
24 3 2 2 11 2 7 2 9 2 13 1 9 1 10 9 2 7 2 9 2 13 1 9 2
9 10 2 9 2 13 15 1 9 2
8 10 10 9 13 1 13 15 2
4 9 1 10 11
6 9 13 9 1 10 9
68 10 9 3 1 10 9 0 13 1 13 10 9 1 10 10 9 2 1 10 0 9 15 15 13 1 10 9 1 10 9 2 13 15 10 9 0 1 10 9 15 13 10 9 1 10 9 0 1 10 9 2 7 13 13 3 2 1 16 10 9 15 13 13 13 10 9 0 2
24 3 10 9 13 1 10 9 1 10 9 1 10 11 2 13 3 2 0 2 10 12 9 13 2
25 16 1 13 10 9 1 2 9 2 2 10 9 3 3 13 3 0 2 1 10 9 13 3 3 2
15 1 10 11 11 13 1 9 1 9 2 13 10 0 9 2
13 11 13 1 12 1 9 1 11 7 12 1 11 2
29 1 10 11 2 11 2 11 2 13 1 10 9 2 13 1 10 9 1 12 1 11 2 11 2 7 12 1 11 2
35 1 10 11 2 11 13 10 10 9 11 1 0 1 10 9 1 13 10 9 0 2 1 12 1 9 2 13 10 0 2 11 2 1 12 2
36 1 13 10 9 2 10 9 1 10 11 13 3 13 1 11 2 11 2 15 13 10 9 1 12 1 9 1 11 16 12 1 11 2 15 1 11
5 11 13 2 13 2
30 10 9 11 2 11 2 13 3 10 9 1 11 13 1 11 1 10 0 9 2 13 3 1 10 9 1 10 0 9 2
19 10 9 0 13 10 0 9 1 10 0 9 1 10 9 2 13 12 9 2
17 2 3 13 1 13 9 1 10 9 7 1 10 9 15 13 3 2
28 1 9 1 10 9 2 10 9 13 1 13 9 7 13 1 10 0 9 2 3 1 10 9 2 2 13 11 2
22 13 2 3 2 1 10 0 9 2 10 9 13 3 1 13 10 9 1 10 0 9 2
27 10 9 13 1 10 9 11 2 11 2 15 13 10 9 1 9 1 9 2 13 3 10 9 1 10 9 2
3 9 3 13
9 0 9 1 11 2 3 13 3 2
50 11 2 10 9 0 15 13 3 2 1 10 9 13 2 13 13 10 0 9 1 10 9 0 1 10 9 0 11 2 3 13 3 13 10 9 1 0 9 2 13 10 9 2 11 2 1 10 9 13 2
21 11 2 9 1 10 11 7 9 1 10 11 2 11 2 2 13 13 10 9 0 2
44 10 9 1 10 11 13 0 2 13 13 1 3 12 9 1 9 2 1 9 1 12 2 7 10 9 1 10 9 1 10 0 12 9 13 13 3 10 9 15 13 10 10 9 2
52 10 9 3 13 3 0 1 10 10 9 1 9 2 15 15 13 3 1 9 1 10 9 1 10 9 7 1 10 9 1 10 9 1 9 1 10 9 1 12 9 1 9 1 10 11 2 13 1 9 7 9 2
33 3 1 10 9 1 12 2 10 9 1 10 11 13 2 1 9 2 3 12 9 1 9 1 10 9 0 1 10 9 1 10 9 2
25 13 15 16 10 9 13 13 1 10 10 3 9 1 9 2 15 3 13 0 13 1 10 9 0 2
39 1 2 11 2 2 10 9 13 13 10 9 3 3 0 2 10 0 9 0 2 7 13 2 1 15 2 3 2 10 9 13 9 2 9 2 9 1 9 2
2 13 2
48 7 15 3 15 13 1 10 9 13 16 2 1 10 9 1 9 0 2 7 1 10 9 1 9 2 0 2 1 9 0 2 13 9 10 9 13 1 9 2 9 2 9 7 9 2 9 13 2
8 10 9 13 2 9 1 9 2
55 3 2 1 10 0 9 2 11 2 9 7 9 1 11 1 10 9 1 10 9 2 13 1 10 9 15 10 9 15 13 13 1 11 2 13 1 13 1 10 9 1 10 9 2 1 10 2 9 2 1 15 11 13 11 2
17 7 2 1 10 9 2 11 13 16 2 1 15 2 13 10 9 2
68 3 2 13 1 13 15 1 10 9 10 9 1 10 9 2 1 10 9 7 1 10 9 2 1 10 9 2 1 10 0 7 1 10 9 2 1 10 9 15 15 13 2 9 15 13 15 9 2 13 2 3 2 7 2 3 2 10 9 15 13 10 9 1 9 1 10 9 2
43 3 2 10 9 1 15 11 2 11 2 13 1 10 9 1 9 13 7 13 10 9 7 10 9 1 11 2 3 10 9 1 15 15 15 13 13 1 10 9 1 10 9 2
44 1 10 9 13 1 10 9 0 1 13 10 9 1 10 9 1 10 9 9 2 10 11 13 10 10 9 1 10 9 0 1 9 1 9 1 10 9 1 10 9 1 10 9 2
78 3 13 3 11 9 1 9 2 9 1 15 10 9 13 1 10 0 2 7 11 2 1 10 10 9 2 11 2 2 1 15 13 15 1 10 10 9 1 10 9 2 13 16 11 13 10 9 1 11 1 12 2 13 1 15 13 9 1 9 1 12 2 9 1 15 9 1 10 11 2 1 9 2 13 10 10 9 2
33 13 3 1 10 9 10 9 1 10 9 1 10 9 12 1 9 1 12 9 2 15 13 13 13 15 15 13 1 13 3 12 9 2
60 3 2 13 15 10 11 2 13 1 10 9 1 10 9 13 1 10 9 1 10 9 7 1 15 13 10 9 11 2 11 2 10 9 11 7 10 9 11 2 1 15 13 10 9 1 13 1 10 0 9 15 15 13 1 10 9 1 10 11 2
14 13 15 10 9 1 9 1 11 2 15 10 11 13 2
2 9 0
20 13 10 9 1 10 0 9 0 2 10 11 13 10 9 1 3 1 9 13 2
25 1 10 9 2 3 3 10 9 15 13 1 13 1 15 13 1 0 9 2 3 9 1 9 0 2
9 10 9 11 13 1 10 12 9 2
34 1 10 9 2 9 1 0 9 1 10 9 11 2 15 13 1 10 0 9 2 1 10 9 1 10 9 1 11 2 12 12 9 2 2
34 13 15 16 11 2 3 1 11 2 13 1 10 0 9 2 7 10 0 9 1 10 9 13 0 7 1 10 9 0 13 15 10 9 2
49 10 9 11 2 9 1 10 11 2 1 15 13 11 1 12 2 12 2 12 2 12 9 3 1 13 13 1 10 10 9 10 10 0 9 1 9 2 13 10 0 9 7 13 10 9 0 1 11 2
36 1 11 2 12 12 9 2 2 1 10 11 7 3 1 9 2 10 9 13 10 9 11 2 15 13 1 10 9 10 9 11 1 12 2 12 2
19 11 1 10 0 9 0 2 13 1 10 9 1 10 3 0 9 0 9 2
30 9 7 9 1 15 10 9 0 2 10 9 0 0 2 10 9 7 10 9 0 7 10 9 0 15 13 1 0 9 2
24 3 1 11 2 11 2 11 2 11 7 11 2 13 10 9 1 10 11 15 13 1 10 11 2
3 9 0 2
4 9 11 11 2
8 9 2 12 2 1 10 9 2
6 11 13 9 3 0 2
35 10 9 7 9 0 11 2 12 9 2 9 2 13 9 12 2 2 13 3 10 9 1 10 0 9 1 9 0 1 10 9 1 10 11 2
51 1 9 1 9 13 3 1 10 9 1 10 9 2 10 9 0 11 2 12 9 2 11 13 16 2 1 2 9 1 9 2 2 13 16 2 10 0 9 1 9 0 2 0 2 9 2 13 1 10 11 2
13 2 1 13 10 9 1 10 9 0 2 2 13 2
41 10 9 13 13 1 13 2 11 2 2 10 9 13 1 11 2 1 11 2 7 13 13 2 11 2 2 15 13 1 9 10 9 2 10 9 1 15 15 13 0 2
33 1 9 13 13 10 9 1 10 9 1 2 11 2 2 10 9 1 13 1 10 9 11 1 9 1 10 2 9 2 0 1 11 2
3 10 0 11
49 10 11 13 1 13 16 13 10 9 3 0 1 10 11 2 11 2 2 1 15 13 1 10 9 1 9 10 10 0 9 1 9 2 13 10 10 9 1 10 11 1 10 0 9 1 12 2 12 2
60 1 9 1 10 9 3 11 2 9 0 1 10 9 1 10 11 2 15 13 10 10 9 1 13 10 9 1 10 9 1 10 11 2 13 3 1 13 13 15 1 10 9 1 10 9 2 16 10 9 3 13 13 1 1 10 9 1 10 9 2
38 1 9 1 10 11 2 11 13 13 10 10 9 2 1 13 0 10 9 3 13 1 10 11 2 15 15 13 4 13 1 10 10 11 1 10 13 9 2
27 11 13 10 10 9 0 1 10 9 2 13 16 10 9 1 9 1 10 11 1 9 15 13 13 12 9 2
45 2 15 13 0 13 0 2 2 13 11 2 13 13 16 13 13 10 9 3 2 3 13 9 13 2 1 0 9 1 10 11 2 13 1 13 3 15 9 1 9 0 1 10 9 2
28 1 11 2 1 1 10 9 12 2 10 11 13 3 12 9 1 10 10 9 1 9 1 10 9 1 10 11 2
47 10 9 1 10 9 1 10 11 1 9 0 1 10 9 13 2 1 10 0 9 2 1 10 9 1 10 9 1 9 1 10 11 0 2 15 13 3 1 10 9 10 10 0 9 1 9 2
18 2 3 15 13 13 16 13 2 2 2 13 11 2 1 13 10 9 2
47 3 1 9 0 1 10 9 1 10 10 9 7 10 0 9 1 1 15 2 13 10 0 9 2 3 11 13 3 10 9 3 13 13 7 13 10 9 1 10 10 9 1 10 9 1 11 2
94 10 9 3 1 10 9 1 10 9 15 2 1 3 12 9 2 13 10 11 0 7 10 9 1 10 11 2 13 13 10 9 3 15 13 2 10 9 1 13 9 1 10 9 11 2 13 1 9 1 9 1 10 9 1 10 9 1 10 9 1 10 9 2 1 15 15 13 13 10 0 9 1 16 13 13 10 13 9 0 15 13 10 9 7 9 1 10 9 1 10 10 9 2 2
26 11 13 3 10 2 9 2 0 1 10 11 2 15 15 13 3 1 10 9 1 10 11 2 11 2 2
29 10 9 0 13 10 3 0 1 10 0 9 1 9 1 9 2 13 1 12 9 1 9 10 10 9 1 9 11 2
25 10 11 13 3 13 10 10 12 9 1 10 0 9 1 10 9 0 2 10 9 15 13 10 9 2
97 3 1 10 0 7 0 9 1 10 11 2 13 12 9 2 7 1 10 0 9 13 1 10 9 13 1 10 9 0 2 3 1 10 9 1 11 2 11 13 10 3 0 1 10 12 9 15 13 1 9 2 13 11 7 11 2 2 10 11 13 1 11 16 10 10 9 13 1 13 2 13 10 9 1 16 15 13 13 1 9 1 9 1 10 11 7 10 11 2 10 12 9 13 1 10 11 2
31 11 13 15 13 12 1 15 3 13 1 10 0 9 2 10 9 13 3 1 10 10 11 2 9 0 1 10 2 11 2 2
16 2 10 11 13 9 2 15 13 10 9 3 13 1 10 9 2
17 13 0 3 13 16 15 13 10 9 1 9 2 3 15 1 9 2
15 10 9 13 1 13 9 2 7 3 13 15 1 13 2 2
42 3 2 11 2 9 1 10 11 2 13 3 16 2 1 10 9 1 15 13 1 10 0 11 2 11 2 11 13 13 2 16 3 3 15 13 3 10 9 1 10 9 2
34 1 2 13 9 16 13 9 0 7 0 1 10 9 2 2 10 9 13 3 10 9 7 3 3 15 13 16 13 9 1 13 10 9 2
12 3 3 15 13 3 7 3 13 10 9 0 2
12 13 2 9 13 2 1 9 1 10 9 2 2
19 10 9 1 10 11 13 3 16 13 0 13 10 9 13 10 9 1 11 2
18 2 13 13 1 12 9 2 7 16 3 13 0 9 13 10 9 2 2
6 9 13 15 1 10 11
28 10 9 7 10 9 15 15 13 1 13 9 1 10 11 2 13 10 9 1 12 9 2 13 13 1 10 11 2
21 3 2 2 10 9 3 13 13 16 3 13 1 4 13 10 9 2 2 13 11 2
50 1 10 12 12 9 15 10 11 13 3 13 13 1 10 9 1 9 1 10 9 2 2 15 13 2 3 2 3 7 1 15 13 13 2 3 16 1 10 9 1 9 3 0 3 15 13 3 12 9 2
78 13 10 9 1 15 13 1 10 11 1 10 0 9 1 10 9 2 1 9 1 9 1 10 0 0 7 10 9 0 1 10 9 2 10 9 13 3 2 1 15 2 10 9 2 11 2 10 0 1 10 11 2 11 2 7 3 9 1 10 11 7 1 10 11 2 10 0 9 13 13 1 10 11 1 10 0 9 2
38 1 10 3 0 9 1 10 9 0 1 10 9 1 10 9 2 15 13 2 0 2 7 2 0 2 2 11 13 10 9 1 10 0 9 1 10 11 2
42 2 1 10 0 9 2 15 3 10 11 13 1 9 0 2 2 2 13 10 9 2 13 1 10 0 9 1 10 9 1 11 2 15 15 13 1 10 10 9 1 11 2
10 9 1 10 11 2 9 13 2 9 0
32 10 11 2 11 2 2 10 9 0 15 13 10 9 7 10 9 2 13 4 1 13 10 9 2 1 10 9 0 1 10 9 2
32 15 15 13 13 10 9 11 2 1 10 9 13 2 1 15 15 13 13 2 10 3 0 9 1 10 9 0 1 10 11 2 2
75 13 1 10 11 2 10 9 0 2 11 2 13 10 9 2 12 9 0 1 10 9 7 1 10 9 1 10 9 2 2 13 2 2 1 10 9 0 2 13 4 10 9 1 10 9 7 4 10 10 9 1 10 9 1 9 7 1 10 9 1 13 10 10 9 13 2 1 10 9 0 1 10 9 2 2
31 10 9 13 16 13 13 10 9 1 10 11 1 13 10 9 1 9 1 0 2 13 10 9 1 13 10 9 1 10 9 2
19 3 3 1 10 11 3 13 13 2 1 3 2 10 9 1 9 1 9 2
49 1 10 9 1 15 2 3 1 9 1 10 11 2 3 1 9 1 10 9 13 3 12 9 2 13 0 1 10 9 16 10 9 1 9 0 15 13 1 12 9 2 1 10 9 0 13 1 12 2
28 10 9 13 4 13 1 10 9 2 3 1 10 11 2 1 15 10 9 0 1 9 13 1 12 1 12 12 2
10 3 1 11 7 1 10 11 13 9 2
54 15 15 13 2 3 2 13 16 1 10 9 10 9 1 9 1 10 9 1 9 1 11 3 13 10 12 9 7 10 9 1 10 9 1 9 1 12 1 9 13 13 10 9 15 13 1 10 9 3 0 1 10 9 2
13 2 10 9 13 16 10 9 0 13 1 10 9 2
19 3 10 9 13 13 3 2 13 10 12 9 2 3 13 15 1 10 0 2
64 3 16 3 15 13 13 10 9 15 3 13 13 3 10 9 15 13 2 2 13 11 2 13 16 10 11 3 13 15 16 13 1 10 9 1 10 9 7 13 16 10 9 3 13 1 13 3 10 9 2 3 13 10 9 1 10 11 2 1 15 10 11 13 2
21 10 9 1 9 1 9 0 9 13 13 1 10 11 1 11 7 11 1 9 13 2
10 10 11 3 13 10 9 1 10 9 2
27 1 10 9 2 10 11 3 13 1 13 0 9 1 9 1 9 0 2 7 13 13 9 0 2 1 11 2
37 15 16 2 13 4 13 11 2 11 2 2 1 15 3 13 10 9 13 1 13 9 15 13 4 1 13 1 9 1 10 11 2 2 13 10 9 2
17 1 10 9 1 10 9 0 15 13 2 0 2 13 10 9 13 2
16 15 1 10 11 2 3 2 15 13 10 9 1 10 10 9 2
7 11 13 10 0 1 13 2
20 3 2 13 15 10 9 11 7 10 9 11 2 9 1 10 9 2 0 2 2
13 10 11 13 0 7 13 10 9 3 1 10 9 2
19 3 1 10 9 1 12 9 0 1 11 2 3 13 3 7 13 1 11 2
32 10 3 0 9 1 10 11 2 1 10 11 2 1 10 9 2 13 3 7 2 1 10 9 2 11 13 1 3 1 10 9 2
21 16 10 0 9 1 10 9 13 13 1 10 0 9 0 2 10 0 13 3 3 2
9 10 9 13 10 9 1 10 9 2
21 7 10 0 9 1 10 9 1 10 9 1 10 9 13 13 10 9 1 10 9 2
21 1 10 9 1 10 9 2 1 10 9 0 1 10 11 2 11 13 10 9 0 2
17 15 13 3 10 0 0 9 1 12 2 15 10 0 9 13 13 2
17 10 9 1 9 13 1 10 9 10 9 2 15 1 0 9 3 2
12 10 2 9 2 13 10 0 9 1 10 9 2
19 13 13 1 10 9 0 2 13 1 10 9 2 1 9 1 9 1 9 2
31 3 10 9 0 3 13 13 10 9 1 10 9 1 12 1 12 9 1 9 7 13 1 10 9 0 1 12 9 1 9 2
18 1 10 9 1 10 9 13 15 12 9 7 13 13 12 9 1 9 2
45 3 1 10 9 13 10 0 9 0 15 13 10 9 7 15 13 1 10 9 2 3 16 13 13 10 9 1 9 13 2 0 7 0 1 10 9 1 12 9 2 15 13 10 9 2
14 10 9 1 10 9 2 9 7 9 3 13 13 15 2
12 10 9 13 13 7 13 1 9 0 7 0 2
6 11 2 10 0 9 0
2 3 0
51 2 13 16 13 0 2 2 13 10 0 1 10 9 11 2 10 0 9 0 1 10 11 1 10 9 1 10 9 2 3 12 1 10 13 9 1 10 2 9 2 0 2 16 13 1 10 9 1 10 9 2
23 0 16 10 10 9 2 10 11 2 10 11 13 9 0 7 0 2 3 0 7 3 0 2
35 10 9 1 2 9 0 1 9 1 10 10 9 2 2 1 10 9 1 11 2 13 1 10 9 1 9 10 9 7 10 9 1 10 9 2
47 9 7 9 13 1 3 13 7 13 2 7 13 0 16 10 9 11 2 2 11 2 2 13 13 1 10 0 9 1 10 11 2 13 1 10 9 1 9 15 13 7 13 1 10 10 11 2
4 9 1 10 9
27 10 9 1 10 11 13 3 1 10 9 2 13 10 11 2 1 13 1 10 11 1 10 11 2 1 11 2
43 10 9 1 9 13 13 3 10 9 1 9 1 10 9 2 1 10 9 1 9 0 2 0 13 7 9 1 9 0 2 10 9 1 10 9 2 11 2 7 2 11 2 2
39 10 10 9 13 13 1 10 9 1 10 9 11 2 13 9 1 10 2 11 2 2 2 10 9 13 3 10 0 1 10 9 1 10 9 2 11 7 11 2
10 9 1 10 11 7 11 13 9 1 9
6 1 10 9 1 9 0
26 13 3 13 10 9 1 9 0 15 13 13 10 9 1 10 9 0 7 15 1 10 9 1 9 0 2
34 13 1 10 9 11 2 10 9 2 13 1 9 1 10 9 1 10 11 7 1 10 11 2 13 12 9 1 13 10 9 7 13 9 2
21 3 2 13 2 2 3 13 10 11 15 13 3 2 2 7 10 2 9 0 2 2
19 2 10 9 0 3 13 9 1 10 9 9 1 13 7 13 10 0 2 2
2 0 9
12 1 10 0 9 2 13 3 4 13 10 9 2
54 13 15 16 2 3 13 9 1 10 9 7 9 1 10 9 9 0 7 1 10 9 1 10 9 0 0 2 1 3 13 1 9 1 9 2 3 13 7 13 1 10 9 0 1 9 2 1 0 9 1 10 11 2 2
43 13 15 3 10 9 1 10 9 2 13 9 1 9 7 9 0 1 10 11 7 9 1 15 13 2 3 1 10 9 0 2 13 10 9 13 3 0 7 13 9 0 2 2
34 3 1 10 9 2 13 10 9 11 2 9 1 10 11 2 7 10 9 11 2 9 1 10 11 2 15 13 10 9 1 10 9 0 2
41 1 10 9 7 9 1 10 0 2 10 3 12 9 2 9 2 0 1 9 0 0 7 0 2 9 7 9 2 13 13 1 10 2 9 0 2 2 7 9 0 2
28 10 9 13 13 1 9 1 10 9 7 9 1 10 2 9 1 9 2 2 13 3 1 9 1 10 9 0 2
27 3 1 10 9 2 10 9 13 15 1 2 9 0 2 2 1 9 0 2 1 13 9 1 10 9 0 2
47 2 11 2 13 10 9 1 0 9 1 10 0 9 1 10 11 2 2 11 2 1 15 10 0 9 1 10 11 13 13 10 9 1 15 10 1 15 13 10 10 2 0 9 7 9 2 2
38 10 9 1 11 2 11 2 13 3 10 9 0 1 11 2 13 13 3 1 11 2 3 13 10 10 9 11 2 7 3 1 11 3 13 1 4 13 2
44 11 2 1 15 10 9 1 9 13 1 2 9 2 2 13 9 1 10 11 1 10 11 7 3 13 1 4 13 1 9 1 13 13 10 9 0 1 13 10 10 9 1 9 2
3 10 9 0
22 10 9 11 2 1 15 13 10 9 0 2 13 1 13 0 10 9 1 3 0 9 2
30 3 13 13 1 16 10 9 11 13 1 10 10 9 1 10 9 1 10 9 0 12 1 10 0 9 1 10 10 9 2
13 13 16 13 10 9 2 7 1 9 0 7 0 2
58 10 9 2 0 7 0 2 13 10 9 1 0 9 2 7 3 13 9 1 10 9 0 1 11 1 10 15 3 0 9 2 11 2 1 10 11 2 9 2 2 11 2 1 10 11 2 9 2 7 11 2 1 10 11 2 9 2 2
35 1 9 2 11 3 3 13 9 1 13 11 2 1 10 11 2 0 1 10 9 7 0 0 2 2 7 11 2 1 10 11 2 0 2 2
12 10 9 1 15 0 13 13 9 1 10 9 2
16 3 2 13 1 10 9 1 9 3 13 11 2 1 10 11 2
17 15 13 15 3 1 10 9 1 11 13 13 10 9 1 0 9 2
29 9 0 1 15 13 0 1 10 9 1 9 15 15 13 1 11 7 13 7 13 10 9 1 10 9 0 7 0 2
48 11 2 15 15 13 2 3 13 2 1 15 13 9 1 10 9 1 10 10 2 0 9 2 2 13 10 9 1 10 2 13 3 12 9 2 1 10 11 2 9 0 15 10 9 11 13 3 2
3 13 11 2
43 2 3 13 10 9 13 1 13 2 11 13 15 2 1 10 9 0 0 2 1 10 9 1 11 2 2 13 0 13 10 11 0 2 2 7 13 16 10 9 13 10 9 2
17 13 10 9 3 13 7 13 10 9 15 13 0 13 1 9 2 2
4 9 2 6 2
19 13 15 1 13 7 13 0 9 16 13 1 13 10 9 1 10 10 9 2
14 9 2 10 9 13 1 9 7 13 1 10 10 9 2
12 10 9 1 0 9 13 15 1 10 10 9 2
8 13 10 9 1 10 10 9 2
11 9 2 10 2 9 2 13 3 1 11 2
16 9 2 13 3 13 16 11 13 15 3 1 10 9 1 9 2
19 7 16 13 3 10 10 9 2 15 1 3 15 9 13 10 9 3 15 2
10 16 13 13 2 13 12 9 7 12 2
12 10 9 1 3 13 0 7 3 13 10 0 2
32 10 9 2 1 10 0 12 9 2 9 7 9 13 9 1 9 1 10 9 7 1 10 9 0 2 9 3 13 1 9 0 2
31 1 9 2 3 2 11 13 10 9 1 9 2 15 13 13 0 7 1 10 9 13 1 9 2 1 13 3 13 10 9 2
11 11 13 12 9 1 9 1 2 11 2 2
10 10 9 1 10 11 1 10 9 11 2
21 15 15 13 11 13 10 9 1 3 12 9 2 3 12 5 16 1 10 9 0 2
22 1 10 10 9 13 12 9 0 10 9 1 9 13 2 1 10 9 1 9 15 13 2
33 2 10 0 9 13 3 10 9 2 2 13 11 2 12 1 10 0 1 10 9 1 10 9 1 11 2 9 1 10 9 1 11 2
18 3 2 10 11 13 1 10 10 9 2 13 1 9 10 9 0 0 2
19 13 2 3 2 10 9 1 10 9 0 1 13 1 10 9 9 1 9 2
42 10 11 0 13 16 13 1 9 10 1 13 1 9 10 9 1 9 2 13 15 0 2 1 10 0 1 10 9 1 10 9 0 2 1 15 15 13 1 13 9 0 2
21 9 13 1 10 11 2 11 2 11 2 11 7 11 13 3 1 13 1 10 11 2
39 7 10 9 1 9 13 13 1 10 9 1 10 9 1 16 3 13 13 3 1 13 9 7 16 10 11 3 13 10 9 0 2 13 15 10 10 0 9 2
40 1 10 9 1 10 11 7 1 10 9 15 3 3 15 13 2 11 13 3 13 13 3 3 9 1 10 9 15 13 1 10 9 2 13 10 9 1 10 11 2
21 9 15 2 3 2 13 1 13 13 1 9 1 10 9 15 15 13 1 10 11 2
54 2 1 10 0 11 3 10 9 13 13 2 3 10 9 1 10 9 0 1 10 9 7 15 1 10 9 1 9 2 13 1 10 0 9 2 7 15 13 13 2 3 13 10 9 1 9 1 10 11 7 10 9 2 2
70 10 9 1 10 11 1 10 11 2 11 2 11 2 1 10 9 2 13 16 10 9 1 10 9 15 13 10 9 1 10 11 2 15 13 13 2 1 10 0 2 1 10 9 2 13 13 9 1 10 11 2 11 2 16 10 9 13 1 10 10 9 2 3 1 10 9 1 10 11 2
4 9 2 0 2
26 2 2 11 2 2 13 1 10 9 1 11 2 11 2 7 13 1 10 9 1 11 2 13 1 13 2
15 13 11 7 11 1 10 11 2 3 1 10 9 1 9 2
37 11 13 10 0 2 7 13 16 11 2 10 9 1 9 2 13 1 13 1 10 10 9 2 11 2 2 9 2 1 13 16 10 10 9 0 13 2
48 11 13 16 2 1 10 10 9 0 2 15 2 13 3 13 3 13 9 1 13 2 7 2 0 9 1 9 7 9 7 15 2 2 15 13 10 9 1 10 9 15 15 13 13 3 2 9 2
20 2 11 2 2 1 11 2 1 11 2 3 13 1 4 13 1 10 9 0 2
23 11 13 10 9 1 10 10 9 15 15 13 1 13 1 10 0 9 1 0 1 10 11 2
7 1 3 3 13 13 13 2
38 3 13 13 10 9 15 13 11 1 13 9 1 10 9 1 10 0 10 9 2 3 15 3 3 13 1 13 3 1 2 11 2 7 1 2 11 2 2
25 10 9 1 9 2 13 7 0 2 13 3 3 13 10 9 2 3 1 15 1 0 9 1 9 2
18 7 10 9 13 1 13 1 10 9 0 9 13 1 12 9 0 0 2
2 9 0
28 2 10 9 1 10 9 13 13 15 1 9 0 2 2 13 11 2 9 1 10 0 9 1 9 1 10 11 2
6 7 15 13 15 2 2
13 11 13 10 10 9 1 10 11 2 1 10 11 2
22 0 9 1 10 9 1 10 11 1 10 9 1 10 11 7 1 10 11 1 10 11 2
44 10 9 13 13 13 15 1 10 9 1 10 9 0 1 10 9 1 9 2 13 1 10 9 1 10 0 9 1 9 2 7 13 10 9 1 10 10 9 0 1 10 9 0 2
60 16 3 13 2 3 2 10 0 9 1 10 9 1 10 9 1 9 1 10 9 2 10 9 0 13 1 13 15 15 3 13 1 10 9 1 11 2 11 7 11 2 10 9 0 1 10 9 0 2 1 15 10 9 13 3 10 9 13 0 2
3 9 1 11
5 10 9 13 10 9
79 9 1 10 12 9 15 13 3 9 1 10 9 1 10 11 2 9 1 10 11 2 0 1 10 11 7 1 10 9 9 1 10 9 2 10 11 2 13 15 2 1 10 9 2 1 10 9 2 1 13 10 9 3 13 13 10 9 0 15 13 10 10 9 15 3 13 4 1 13 1 13 0 10 9 13 1 10 9 2
54 1 10 9 1 9 2 13 3 1 10 9 2 13 15 2 3 2 10 9 2 1 10 0 2 3 12 9 0 13 1 10 9 1 10 11 2 2 1 10 10 2 10 9 0 2 11 2 11 2 11 2 11 2 3
37 9 15 13 1 10 10 9 9 1 9 7 9 1 9 0 1 9 1 9 1 9 2 9 1 9 1 9 1 9 1 13 3 12 9 1 9 2
38 13 1 9 1 11 2 10 9 1 15 2 3 1 10 9 2 7 1 10 9 0 2 2 10 0 9 13 10 1 10 9 0 3 1 10 10 9 2
15 10 9 3 3 13 9 1 9 1 9 1 9 1 9 2
30 11 2 2 11 2 2 13 10 0 9 0 1 9 2 9 13 1 10 11 2 15 13 1 10 0 9 1 10 11 2
22 10 9 1 10 11 13 10 9 2 3 13 10 12 0 1 10 9 1 10 12 9 2
19 10 11 2 1 12 9 1 10 12 0 9 2 13 10 9 0 1 9 2
24 3 2 13 1 13 15 10 11 2 9 1 9 2 1 10 11 2 1 10 9 12 1 9 2
1 11
21 11 2 2 0 2 2 13 10 9 1 10 11 2 15 3 15 13 1 10 11 2
19 1 10 0 9 1 10 12 9 2 11 2 1 10 11 2 13 10 9 2
10 10 11 2 1 11 2 13 1 9 2
20 1 10 11 2 3 13 10 11 2 13 1 9 7 10 9 13 1 10 11 2
1 9
3 10 0 9
46 13 1 10 9 11 2 1 10 0 9 1 9 1 10 9 2 3 10 9 7 10 9 15 13 1 10 9 1 9 2 13 13 1 10 9 2 3 0 13 10 9 0 1 10 9 2
21 7 11 13 13 1 10 9 1 10 2 9 1 15 13 2 1 10 9 3 0 2
38 10 10 9 13 13 15 1 10 11 2 3 11 13 10 9 1 12 1 10 12 9 1 10 2 3 0 7 3 0 9 1 10 9 2 2 10 9 2
28 13 3 12 9 2 12 1 13 1 11 2 10 0 9 1 10 11 2 7 12 1 13 1 11 2 1 11 2
42 11 3 13 10 9 0 7 2 1 15 13 10 0 1 12 1 10 9 1 11 2 15 1 11 2 9 1 11 2 15 13 16 3 10 9 13 0 1 10 0 11 2
39 1 15 2 1 15 13 10 9 1 11 2 13 16 13 3 3 16 10 11 2 15 3 13 1 15 1 11 10 9 1 13 13 1 10 11 2 9 2 2
5 11 13 1 10 9
20 10 11 13 13 1 1 10 9 1 10 9 12 12 9 1 9 1 9 0 2
32 7 2 1 10 9 13 1 10 9 2 1 10 9 1 0 9 11 2 1 12 2 10 9 1 12 13 1 10 9 7 9 2
28 10 13 2 9 0 2 2 11 2 7 10 9 1 0 9 11 13 9 1 10 9 0 1 9 1 9 0 2
7 11 13 9 1 10 9 0
59 10 11 13 3 16 10 10 9 2 11 2 3 13 10 9 1 9 15 15 13 13 1 10 9 1 9 1 11 2 13 13 10 11 1 9 0 13 10 9 1 9 1 10 9 0 2 1 9 1 13 13 1 10 9 1 10 9 0 2
68 2 10 9 1 10 11 13 16 10 11 13 13 10 9 2 13 3 1 13 9 3 9 2 9 1 15 13 10 9 1 10 9 2 2 13 1 10 11 10 9 1 10 9 1 10 11 1 11 2 11 2 13 16 13 13 1 10 11 7 1 10 11 10 9 1 9 0 2
16 7 2 10 9 13 1 10 9 15 13 13 2 2 13 11 2
33 2 10 11 13 13 1 15 15 15 3 13 2 15 3 13 1 13 10 9 1 10 11 2 13 15 10 9 1 10 9 0 2 2
31 2 10 9 13 10 9 1 10 9 1 13 2 3 2 7 13 15 0 1 15 13 2 10 9 2 10 9 1 10 10 2
15 3 13 10 0 9 15 3 13 1 10 10 9 1 9 2
22 1 10 9 2 13 15 15 13 13 10 9 1 10 9 7 1 13 1 10 0 0 2
18 10 9 13 1 10 9 0 7 0 2 1 15 2 10 10 9 2 2
35 13 1 10 10 9 7 1 9 13 1 9 0 2 11 13 16 10 0 9 1 10 9 3 13 10 0 9 1 13 1 12 1 12 9 2
12 3 3 2 10 9 0 13 13 13 10 9 2
30 3 2 16 15 13 1 9 1 10 9 7 16 10 0 9 1 13 13 9 15 13 1 13 2 10 9 13 10 9 2
3 15 13 2
20 15 3 2 16 13 0 1 13 1 10 9 1 10 9 1 10 9 7 3 2
39 9 1 9 0 7 1 10 0 2 9 2 1 9 7 9 0 13 1 10 9 12 9 3 15 3 0 1 13 9 1 0 13 1 10 9 1 10 9 2
19 7 15 16 13 10 9 2 0 2 1 10 2 9 0 2 1 10 9 2
31 10 3 0 13 10 11 2 7 11 2 1 10 2 9 1 10 9 2 11 2 3 1 9 0 1 9 0 1 10 11 2
10 10 15 13 10 11 2 9 0 0 2
21 10 2 9 2 1 11 7 1 11 13 3 3 1 10 11 2 7 3 13 13 2
30 15 1 10 9 13 3 3 3 1 10 0 9 0 7 1 10 12 9 1 10 0 9 13 15 3 3 1 10 9 2
21 10 11 13 2 10 9 13 1 13 9 0 2 7 13 15 9 1 10 9 0 2
19 10 9 15 13 1 13 0 2 1 12 9 15 13 3 1 13 3 13 2
21 10 11 13 10 9 1 10 0 9 1 11 2 7 1 10 9 1 10 9 13 2
44 11 13 10 9 1 10 9 2 3 3 3 1 10 9 11 13 1 10 9 1 10 9 2 13 1 11 13 1 10 9 1 10 9 1 10 9 11 2 13 10 9 1 11 2
29 11 13 3 1 10 9 2 13 11 0 1 10 9 1 10 9 2 9 15 13 10 9 0 1 10 2 9 2 2
20 11 13 1 11 1 13 9 1 10 9 1 10 11 0 1 10 9 2 11 2
33 10 9 1 10 11 1 10 11 13 10 9 1 13 16 2 2 1 12 2 3 13 10 9 13 2 1 10 9 2 1 11 2 2
37 1 11 2 2 3 10 9 0 1 10 11 7 1 11 13 13 0 9 1 10 0 9 7 13 2 9 1 11 16 10 9 7 9 13 13 2 2
30 10 9 1 10 9 0 13 9 1 10 9 0 1 13 16 2 1 10 9 0 3 13 13 10 9 1 10 9 2 2
7 2 13 2 13 9 1 11
37 11 2 12 1 10 12 9 2 13 2 1 10 0 9 1 10 11 2 15 13 3 10 9 13 1 12 2 13 3 10 9 1 10 9 0 11 2
27 10 0 9 1 11 1 11 13 12 9 2 13 10 9 0 1 12 7 13 10 9 1 9 1 10 11 2
16 3 3 10 9 1 10 9 13 2 1 10 11 2 9 9 2
8 10 9 1 10 11 13 13 2
7 3 3 13 10 9 0 2
14 3 1 11 2 12 1 10 9 1 10 9 1 11 2
14 7 2 1 11 2 3 15 13 10 9 1 10 9 2
25 13 16 15 3 13 10 9 13 1 10 10 9 1 10 11 7 13 3 0 1 13 9 0 13 2
18 10 9 1 12 12 9 1 10 11 1 10 11 13 3 13 1 11 2
23 10 9 13 16 3 15 13 13 10 9 1 10 9 2 7 3 13 13 15 1 12 9 2
36 13 0 2 3 2 1 15 13 16 2 16 10 11 13 10 9 1 10 9 2 10 9 0 13 1 13 10 9 2 16 15 3 13 4 13 2
33 10 9 0 1 9 7 10 0 9 1 9 1 10 9 13 3 1 10 9 1 10 11 2 1 10 9 1 12 2 3 13 13 2
23 11 13 16 15 13 1 10 9 1 10 9 1 10 11 2 1 15 13 10 9 1 9 2
50 10 0 9 13 10 9 2 0 2 2 13 15 1 10 9 2 9 2 0 13 10 10 9 0 2 1 10 9 2 11 13 1 13 10 9 0 2 2 1 10 9 2 1 0 1 9 1 0 9 2
33 7 2 1 9 1 10 9 2 13 15 1 10 9 0 0 15 13 10 9 13 1 13 10 9 1 10 9 2 1 12 9 10 2
24 10 9 2 3 13 1 10 9 1 9 1 9 2 3 13 13 3 1 10 9 1 10 9 2
43 11 13 15 3 13 1 10 9 7 13 15 3 13 1 10 9 1 10 9 2 2 15 13 1 3 0 9 2 2 13 2 2 15 13 10 9 1 10 10 9 0 2 2
19 2 12 1 10 9 15 3 15 13 13 10 9 1 10 9 1 10 9 2
41 7 10 9 15 13 4 13 3 13 13 9 2 2 13 10 9 2 15 13 10 9 1 10 10 9 1 15 13 16 2 3 13 0 9 7 0 9 16 13 2 2
2 11 13
24 11 2 15 13 3 1 10 9 2 13 0 1 15 13 10 9 15 3 13 10 9 1 11 2
14 10 9 13 10 9 1 2 0 9 2 1 10 11 2
34 2 13 9 1 9 2 2 2 3 15 13 10 9 3 3 15 13 2 2 2 13 15 1 10 9 2 2 2 16 13 3 10 9 2
10 2 7 10 9 13 1 4 13 2 2
27 3 11 13 2 10 9 13 1 10 9 2 15 13 10 15 13 7 15 15 13 13 3 1 13 1 11 2
8 1 15 2 11 13 0 9 2
45 12 7 15 13 10 10 9 2 3 13 10 9 0 1 15 2 10 0 9 13 16 2 1 10 0 2 15 13 10 13 9 1 11 7 2 1 10 0 2 10 9 13 3 0 2
36 15 13 3 1 15 15 15 13 2 9 1 11 2 2 1 15 15 15 13 13 16 2 13 10 10 9 2 2 7 13 16 15 13 1 13 2
3 15 13 2
4 9 0 13 13
4 13 15 10 11
5 11 2 1 11 2
17 10 0 9 0 13 1 13 1 10 9 11 3 13 1 10 11 2
20 1 11 2 15 13 13 10 9 2 13 10 0 9 15 3 15 13 4 13 2
14 13 9 1 10 9 1 11 3 11 13 11 1 9 0
6 10 9 1 13 10 9
10 11 13 1 13 10 11 1 10 9 2
11 13 16 16 3 13 1 9 2 13 13 2
7 10 11 13 1 10 9 2
9 10 9 0 13 10 9 1 13 2
11 10 9 1 10 9 13 13 7 13 15 2
5 10 9 13 15 2
11 11 13 1 11 16 10 9 13 10 9 2
10 7 10 9 13 13 1 9 1 9 2
27 10 11 13 3 10 9 13 1 10 0 11 1 13 10 9 1 11 2 15 13 13 10 9 1 12 9 2
31 10 9 13 1 10 9 0 13 4 1 10 9 1 10 9 1 9 7 4 1 10 12 9 0 2 11 2 11 7 11 2
61 13 16 10 9 13 3 3 13 2 1 13 9 1 9 7 1 10 0 9 0 2 10 9 13 1 10 9 1 10 11 7 1 10 9 13 1 10 9 0 2 9 1 10 9 0 0 2 13 1 9 10 9 7 9 1 10 11 2 11 2 2
6 11 13 9 1 10 11
35 10 11 13 1 13 9 1 10 9 1 10 9 0 1 10 11 2 13 3 13 1 10 10 9 0 16 13 11 1 10 9 1 10 9 2
19 10 9 1 10 9 0 13 3 16 10 11 13 1 13 10 9 0 9 2
22 10 9 2 11 13 3 2 16 10 11 13 13 10 9 13 1 10 11 2 11 2 2
25 9 10 0 1 10 9 1 10 9 0 2 1 16 10 9 1 10 11 2 11 13 1 10 9 2
6 11 13 9 1 10 11
49 1 10 9 1 10 9 2 15 11 13 3 0 1 10 9 2 10 9 13 3 13 2 2 15 9 2 13 2 2 2 2 2 7 13 9 0 7 0 1 9 2 9 2 9 15 13 9 0 2
48 10 2 9 2 0 13 13 10 9 1 10 9 1 10 9 2 7 12 7 10 15 13 13 1 9 7 9 1 9 7 9 2 16 10 10 9 7 9 13 2 3 2 10 9 7 10 9 2
23 3 2 10 9 13 1 10 9 1 10 9 0 1 10 9 0 2 7 13 15 1 15 2
68 10 9 13 3 13 3 9 2 3 3 3 9 2 0 2 2 16 0 7 3 2 0 7 3 2 10 9 13 10 10 9 2 10 10 9 2 10 10 9 0 7 0 2 9 2 9 2 9 2 9 2 13 2 7 10 10 9 0 7 0 2 9 2 9 2 3 2 2
46 7 10 10 9 2 7 10 9 15 13 2 13 13 1 9 3 0 7 0 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 2 9 1 9 2
72 3 2 13 1 10 9 10 9 0 1 10 9 2 2 0 10 9 2 2 1 3 13 1 10 0 1 10 2 9 2 7 1 10 2 9 1 9 2 2 7 10 9 0 2 2 1 15 13 2 2 2 1 3 13 2 2 2 15 13 2 2 2 9 1 9 2 2 2 0 9 2 2
81 10 9 2 7 2 9 2 2 3 15 13 10 9 2 2 2 11 2 13 7 13 1 10 9 0 2 0 2 0 2 0 1 15 1 10 2 9 2 7 1 10 2 9 2 2 15 3 13 3 1 10 9 1 10 9 2 7 1 10 10 9 2 13 0 10 10 2 9 0 2 7 13 10 9 1 10 10 2 9 2 2
19 10 9 0 1 10 9 7 10 9 3 13 13 9 0 1 10 0 9 2
16 3 13 10 9 2 9 1 10 0 9 0 1 10 12 9 2
31 9 0 13 3 10 9 0 0 2 13 1 13 13 10 9 1 16 10 9 3 13 3 1 13 10 9 1 10 9 0 2
42 7 10 9 0 7 10 9 13 16 13 10 9 0 1 10 12 9 2 3 10 11 7 10 11 13 13 10 9 0 1 10 9 2 16 1 10 9 13 3 10 9 2
24 10 9 13 9 1 10 9 1 10 0 9 1 10 11 2 11 2 9 13 1 10 9 11 2
23 1 10 11 2 10 0 9 1 10 9 1 1 10 9 13 3 4 13 10 9 3 0 2
78 15 16 2 2 1 10 9 2 7 13 3 1 16 11 7 11 13 7 13 2 0 9 2 10 10 9 1 9 7 9 2 13 10 9 13 15 1 10 9 13 10 9 0 1 10 10 9 1 10 9 2 1 11 7 1 0 9 2 3 16 13 10 9 1 10 9 0 1 10 9 0 7 1 9 10 9 2 2
3 3 1 11
5 0 13 15 1 11
27 10 0 9 1 10 9 0 2 11 2 13 13 15 3 1 11 1 13 10 9 15 15 13 1 10 9 2
56 13 3 15 10 9 1 10 9 11 7 1 10 9 1 10 11 2 11 2 3 13 10 9 15 13 13 2 1 10 9 0 1 11 2 10 9 0 7 10 9 0 15 13 13 2 1 9 2 10 9 1 9 0 1 11 2
24 10 9 13 1 10 9 1 10 9 1 9 1 10 11 3 10 9 0 13 3 10 0 9 2
9 10 11 3 13 1 10 9 0 2
13 10 9 0 1 10 2 9 2 13 1 12 9 2
45 1 10 9 1 10 9 13 13 12 9 1 9 1 11 1 12 9 2 1 10 9 0 13 1 12 9 2 1 12 13 1 10 0 9 1 10 10 9 2 13 1 12 1 9 2
55 10 9 1 10 9 1 9 1 10 11 13 13 1 10 9 1 9 1 11 2 9 1 11 2 1 9 13 1 10 9 1 9 1 10 11 2 1 10 10 9 1 10 9 0 2 1 15 9 3 0 13 1 9 0 2
17 9 1 10 9 0 13 3 13 1 13 9 1 13 10 10 9 2
54 1 10 9 1 9 13 1 10 9 2 11 2 11 2 2 13 15 16 1 12 2 9 1 10 9 1 10 11 2 1 9 1 12 2 10 9 2 13 3 13 1 10 9 2 9 2 9 7 9 2 1 10 9 2
53 7 10 9 3 13 1 10 9 1 10 11 2 1 9 1 12 2 16 10 9 9 1 10 9 1 10 9 3 13 13 1 9 0 2 3 10 9 13 2 7 13 13 2 1 10 9 7 9 1 10 9 2 2
106 7 1 10 9 1 10 9 2 7 3 1 10 9 0 1 2 11 2 2 10 9 1 11 15 11 13 3 3 1 10 9 1 10 9 1 10 11 2 13 15 3 10 9 1 10 1 10 10 9 15 15 13 13 2 3 10 1 10 9 2 11 2 2 15 13 2 11 2 2 2 16 15 1 10 9 15 15 13 2 2 11 2 2 13 3 1 9 1 0 9 1 10 9 0 13 1 9 2 13 13 3 2 1 9 0 2
1 11
11 11 2 11 2 9 2 12 1 9 2 9
56 1 10 9 1 3 12 12 9 7 3 10 9 15 13 13 3 3 1 10 9 12 7 3 10 9 0 0 13 1 10 9 0 1 10 9 2 10 9 1 3 13 1 10 9 1 9 13 16 2 10 9 13 3 0 2 2
37 10 12 0 7 12 13 13 9 0 1 10 9 0 0 2 15 13 1 9 1 9 10 9 1 10 9 1 11 2 11 7 11 2 1 9 0 2
24 1 10 9 0 1 12 2 13 12 0 2 7 1 10 0 1 12 10 9 13 1 12 0 2
6 13 1 10 2 11 2
23 1 10 11 2 10 9 1 10 11 13 3 0 3 1 13 10 9 1 9 15 15 13 2
24 13 9 1 15 2 1 10 9 1 1 10 9 2 3 10 9 13 10 0 9 1 15 13 2
17 10 9 13 15 13 1 13 9 1 13 10 9 15 15 13 13 2
54 9 15 2 1 10 9 13 3 1 10 9 1 10 11 7 1 10 11 2 3 15 13 1 10 9 1 10 9 2 7 1 10 13 9 1 9 7 1 10 9 15 13 10 9 1 10 9 16 10 9 2 10 9 2
33 10 9 15 15 13 1 13 2 1 10 10 0 9 2 1 9 3 15 13 3 13 1 10 9 15 1 10 9 13 10 12 9 2
55 7 1 10 3 13 9 1 9 2 3 11 2 1 9 1 11 2 13 16 2 3 13 9 1 9 3 0 2 7 13 1 10 9 1 10 9 1 10 9 1 10 11 1 13 3 13 3 13 3 0 16 1 10 9 2
28 3 10 2 11 2 2 10 9 1 10 11 2 1 9 13 3 1 10 9 1 10 9 2 13 13 1 15 2
69 1 10 0 7 0 9 0 7 10 13 9 1 10 9 1 10 0 7 0 9 2 13 10 10 0 9 2 7 1 10 9 1 9 1 9 2 10 10 9 13 4 1 2 13 2 10 0 9 1 9 0 2 0 7 0 2 13 3 10 9 1 10 9 0 1 10 9 13 2
27 13 0 13 3 1 10 9 1 9 0 7 13 10 9 0 1 15 15 13 13 10 9 1 3 0 9 2
37 13 9 1 9 2 1 10 9 2 9 0 2 9 1 9 1 10 9 7 1 10 11 2 9 1 10 9 1 9 3 0 1 10 11 2 3 3
14 10 9 0 7 3 0 15 10 9 0 13 13 3 2
36 7 15 15 13 3 0 1 15 13 16 10 10 9 13 1 10 9 11 13 13 1 10 9 1 10 0 9 2 3 10 10 10 9 7 9 2
35 13 13 3 1 10 0 9 1 10 9 2 15 3 0 15 13 2 3 2 1 13 9 1 2 9 2 7 15 13 1 13 10 0 9 2
28 7 10 0 9 1 10 11 13 16 10 0 9 0 13 13 10 9 1 13 10 9 15 13 7 13 1 9 2
67 1 3 2 10 9 3 15 1 11 7 1 10 11 13 3 0 1 13 3 7 10 9 2 0 7 3 2 1 10 11 7 3 2 13 10 9 1 9 3 0 16 2 1 15 13 13 2 3 3 13 4 10 9 15 15 13 13 3 3 4 9 1 9 1 3 13 2
6 9 1 11 3 13 9
54 3 3 1 9 1 9 3 10 11 13 10 9 1 10 0 9 1 10 9 1 10 9 2 15 13 3 12 9 2 10 9 1 9 0 2 15 1 12 2 9 2 0 13 10 9 1 10 12 0 9 1 10 11 2
12 3 1 10 11 7 1 10 11 3 15 13 2
36 10 11 13 1 13 1 10 9 1 10 11 2 1 13 10 9 2 13 13 2 3 2 10 9 1 10 1 3 13 1 10 9 1 10 11 2
30 15 1 10 9 1 10 9 0 2 10 11 2 1 10 9 15 10 11 13 10 2 10 11 2 13 11 1 9 2 2
37 11 2 9 2 13 10 9 1 10 12 9 7 13 16 2 10 9 0 13 13 1 10 11 2 2 1 15 10 9 13 4 13 2 1 13 9 2
17 3 16 10 11 3 13 3 10 11 13 10 9 1 10 12 9 2
41 9 13 13 13 10 11 1 10 9 1 10 11 2 15 3 13 13 10 9 0 2 1 10 10 9 7 1 10 10 9 2 7 1 9 3 10 9 3 13 13 2
40 3 2 1 10 9 1 10 9 1 10 0 9 1 10 9 2 10 9 13 1 10 9 3 0 15 13 10 0 9 1 10 9 1 10 9 1 10 0 9 2
60 10 9 15 13 3 1 10 9 1 9 13 2 3 2 10 9 1 9 1 10 11 13 10 0 9 1 10 9 9 2 9 7 2 3 2 10 9 1 10 11 13 13 3 10 9 1 9 7 0 0 3 1 10 12 9 2 7 12 9 2
26 10 0 9 13 1 12 1 9 2 3 10 9 0 0 13 1 10 9 1 12 9 2 1 10 10 9
48 11 2 9 0 2 13 2 1 10 9 13 1 10 9 2 16 12 9 0 3 13 9 0 1 10 9 0 1 10 11 7 13 1 10 9 0 1 10 9 0 15 13 10 0 9 0 0 2
1 11
2 9 13
33 3 1 0 9 1 10 9 2 11 2 3 10 2 9 12 2 1 10 9 2 11 2 11 2 2 13 10 9 1 10 10 9 2
54 1 10 10 9 2 11 2 15 13 3 9 1 10 9 1 10 11 0 7 15 3 15 13 3 3 9 1 10 11 2 2 13 10 11 2 1 9 0 7 2 3 13 1 10 9 1 13 10 9 1 10 9 2 2
28 1 1 10 9 1 10 13 9 2 10 11 13 4 1 13 10 9 1 10 9 2 1 1 10 9 1 9 2
35 10 9 13 1 9 1 9 0 7 0 1 13 10 9 0 1 10 12 9 15 13 13 1 10 9 2 16 10 11 13 13 9 1 9 2
70 10 11 13 13 1 10 9 1 10 9 12 2 1 10 9 1 10 9 1 9 1 9 13 1 10 0 11 2 0 11 2 2 10 11 7 10 9 0 11 2 13 1 10 9 10 11 4 10 9 1 10 9 7 4 1 10 9 1 9 1 13 10 9 1 9 0 1 9 13 2
6 0 9 1 10 9 0
34 10 9 1 9 0 13 4 1 4 3 13 1 10 9 1 9 1 10 9 7 1 10 9 3 0 2 3 1 10 9 12 1 12 2
26 10 9 1 10 9 13 13 10 9 0 1 9 1 9 13 1 10 9 1 9 0 2 3 10 11 2
9 7 3 13 0 1 10 9 0 2
5 9 0 1 10 11
39 1 10 11 1 10 0 9 2 10 2 9 2 0 1 12 9 1 9 2 2 10 9 0 13 2 3 2 13 1 10 0 9 3 3 12 9 1 9 2
12 10 9 15 2 3 2 3 13 10 11 13 2
54 2 13 3 16 10 9 1 10 9 13 1 4 13 1 10 9 0 7 0 2 7 3 10 9 3 15 13 1 10 9 1 10 9 15 13 10 11 7 15 13 10 9 0 1 10 9 1 10 9 2 2 13 11 2
40 1 10 10 9 2 11 13 13 16 10 9 13 1 15 10 9 13 1 10 9 1 10 0 9 2 12 9 2 2 13 16 10 0 11 13 13 10 11 3 2
17 2 10 11 13 13 10 9 2 7 10 9 13 0 2 2 13 2
3 9 2 11
3 9 2 11
65 1 10 9 1 10 9 1 10 11 1 10 9 1 10 9 15 13 11 2 0 9 1 9 13 1 10 9 7 10 10 9 2 15 2 13 9 0 1 10 0 7 0 9 15 13 13 1 9 7 1 9 2 1 9 7 1 9 2 1 9 7 1 9 2 2
5 1 0 9 0 2
3 9 2 11
82 1 10 9 1 10 11 2 10 9 13 13 10 9 1 10 9 1 9 1 9 2 10 9 11 2 1 12 9 2 1 12 9 2 10 11 2 10 13 9 1 12 9 2 1 13 2 1 12 9 2 7 10 13 9 0 11 2 3 10 1 12 9 7 10 11 2 10 3 0 2 9 2 1 10 9 2 15 13 12 12 9 2
51 1 10 9 2 13 15 3 10 9 1 9 1 10 0 11 2 10 13 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 7 11 2 10 0 13 10 2 11 2 1 10 9 2
47 1 9 0 2 13 15 10 11 2 10 0 9 1 12 9 2 1 9 1 12 9 2 13 1 10 9 1 9 2 1 12 9 2 7 10 11 2 10 9 1 9 1 9 1 9 9 2
54 1 10 9 2 10 9 3 13 15 2 13 10 0 9 13 1 10 11 2 1 12 9 2 15 15 13 13 1 9 0 1 0 9 2 1 10 0 7 0 9 11 7 1 10 13 11 2 9 1 9 0 7 0 2
44 1 9 2 13 10 9 0 7 0 1 9 1 9 7 0 2 3 9 2 1 10 0 9 15 13 10 9 1 10 9 2 1 10 9 2 10 11 2 7 11 2 11 2 2
34 1 10 9 1 12 3 12 12 9 0 13 1 10 11 2 13 0 9 2 1 13 1 10 9 7 9 1 10 9 1 10 9 11 2
24 13 15 16 3 12 12 9 13 13 10 10 9 7 9 7 15 13 1 9 0 1 10 9 2
69 3 1 9 0 13 2 1 9 15 13 13 1 10 0 9 2 3 1 10 9 0 2 10 9 15 13 1 3 2 9 7 9 1 9 0 3 3 13 9 2 9 2 9 2 9 0 2 9 13 2 9 13 2 9 7 9 13 1 9 1 15 15 13 13 9 1 9 0 2
72 10 9 1 9 9 0 1 11 13 15 1 10 9 7 9 1 9 0 1 9 13 15 9 2 1 9 1 9 1 9 1 9 0 2 1 9 1 9 2 1 2 9 1 9 2 7 1 2 9 2 1 9 1 10 9 11 2 11 2 11 7 2 1 10 9 2 9 1 9 1 9 2
30 15 1 10 13 2 9 1 9 2 13 13 1 10 11 2 1 10 11 2 11 2 7 1 10 9 11 2 11 2 2
27 10 9 1 10 9 15 1 10 9 1 3 13 1 10 9 13 10 9 7 2 3 2 10 9 1 9 2
53 1 10 9 13 3 13 12 1 15 2 15 15 13 0 1 10 9 0 7 1 10 9 0 7 15 15 15 13 3 1 10 0 7 15 13 13 3 1 0 1 10 9 0 2 15 15 13 13 1 10 10 9 2
56 9 3 1 10 9 2 11 2 9 1 10 11 2 13 9 0 1 10 9 1 10 9 2 10 9 0 1 10 9 2 10 9 0 2 10 9 1 10 0 9 1 10 9 3 0 7 10 9 0 1 10 9 1 10 9 2
17 1 10 9 1 11 1 10 9 0 1 10 9 1 10 9 0 2
24 2 13 1 11 3 13 1 10 10 9 2 16 10 9 1 10 11 13 13 3 1 15 2 2
12 13 13 10 9 0 1 10 9 15 13 13 2
30 3 13 9 2 3 2 16 10 10 9 15 13 1 10 9 1 9 7 9 2 13 16 15 13 0 1 10 9 9 2
8 15 3 13 4 13 1 9 2
13 1 10 9 13 2 13 1 0 9 10 9 0 2
23 13 10 9 13 7 10 9 15 13 3 13 10 9 1 10 0 9 15 13 1 10 9 2
28 13 2 1 10 9 2 16 10 9 13 13 3 2 16 10 9 1 10 11 13 15 1 10 9 1 10 9 2
13 7 10 9 13 1 13 16 13 13 10 10 0 2
28 1 10 9 1 10 9 1 10 9 2 13 9 1 15 13 7 13 13 7 13 2 16 13 13 10 9 0 2
31 1 10 9 2 13 10 9 1 10 9 13 0 1 10 9 2 1 13 10 9 3 2 1 13 9 1 10 9 1 9 2
11 7 13 16 10 9 13 1 13 1 12 2
22 3 2 12 1 10 10 9 13 10 9 1 11 7 11 2 7 3 10 9 1 11 2
36 10 9 0 1 10 0 13 3 1 10 2 9 1 9 2 1 10 9 0 1 10 9 2 1 13 15 1 10 9 0 1 10 9 1 9 2
42 1 13 10 11 1 10 9 0 1 10 9 2 11 2 13 1 10 9 1 10 9 2 13 16 10 11 13 2 13 10 9 1 0 7 3 0 9 1 9 0 2 2
5 11 1 9 1 9
25 10 11 7 10 11 13 10 9 1 9 1 13 1 11 2 10 11 2 15 13 9 0 1 11 2
41 10 9 13 13 1 10 9 1 10 9 7 2 1 10 0 9 2 10 11 13 12 5 1 10 9 7 10 11 12 5 2 13 10 9 4 1 13 10 9 0 2
18 13 13 10 9 1 12 5 1 10 9 0 2 3 1 12 9 0 2
4 13 13 12 9
18 10 9 13 1 13 9 1 10 9 0 7 1 10 9 1 10 9 2
31 7 2 16 15 13 16 10 9 1 9 1 11 13 3 0 16 10 1 10 11 2 15 3 13 15 16 13 13 16 3 2
8 3 1 10 0 9 1 9 2
1 0
3 11 2 11
5 10 9 13 15 2
16 10 9 1 10 9 2 7 10 9 1 10 9 15 15 13 2
30 10 9 0 1 10 9 1 10 11 13 12 1 10 9 15 10 9 0 1 9 0 3 13 4 1 13 1 9 13 2
15 13 3 2 12 9 1 0 9 0 2 1 9 3 9 2
36 16 10 9 13 0 2 3 1 10 9 1 10 9 13 1 10 9 3 1 10 9 15 15 13 2 2 1 10 9 10 9 3 13 9 0 2
16 16 11 7 11 13 2 3 2 10 9 0 1 13 7 13 2
29 16 13 13 0 2 1 0 9 2 16 13 0 2 1 13 0 9 2 16 13 13 7 13 15 1 13 9 0 2
8 3 12 9 1 10 11 1 9
9 2 9 1 9 2 3 13 9 2
48 2 10 9 13 1 15 2 15 13 10 9 2 13 15 1 15 2 2 13 11 2 9 1 9 1 11 2 3 15 13 1 13 1 10 9 13 1 10 11 2 11 2 2 3 2 1 11 2
7 2 11 2 13 10 0 9
5 10 9 13 1 11
4 11 2 1 11
13 13 10 2 11 2 1 12 2 13 15 1 12 2
30 10 9 13 13 10 9 1 10 9 2 7 10 0 13 13 15 0 2 1 3 1 12 9 2 1 10 9 1 11 2
6 7 3 13 10 9 2
29 10 9 13 3 3 13 16 10 11 15 13 3 1 11 2 7 16 15 13 1 10 9 2 7 3 10 9 13 2
31 10 9 0 1 10 9 1 9 13 10 9 1 16 10 11 13 13 1 10 9 1 9 2 10 9 15 13 0 9 0 2
16 13 10 9 1 10 9 1 10 11 13 10 9 1 10 9 2
23 10 9 1 11 1 13 10 9 1 9 13 1 11 1 12 13 1 10 10 9 1 11 2
18 11 2 10 9 0 13 10 0 9 2 13 3 3 0 1 10 9 2
28 13 0 16 1 10 9 10 9 0 15 13 13 1 13 10 9 1 10 9 2 9 1 9 3 0 1 11 2
10 7 10 9 1 11 3 13 3 0 2
8 10 9 1 10 9 13 15 2
13 10 9 1 10 9 13 1 10 9 13 13 0 2
9 12 1 10 12 9 13 1 9 2
34 10 11 0 13 16 10 9 13 13 3 1 10 9 1 10 9 2 3 1 10 0 9 1 10 9 2 7 2 3 2 13 3 13 2
18 1 10 9 1 9 2 13 15 10 0 9 1 10 9 1 10 9 2
30 10 11 13 13 1 13 7 13 10 9 1 16 10 9 13 4 10 9 1 10 9 7 1 10 9 7 4 10 11 2
32 13 15 15 13 3 13 1 10 9 2 13 15 2 3 15 13 2 16 10 9 1 10 11 13 10 9 0 1 10 9 0 2
34 1 1 11 10 9 13 3 1 9 2 13 1 10 9 13 1 9 1 10 0 9 2 10 11 13 1 10 0 9 1 10 9 0 2
43 3 0 2 16 16 13 0 9 0 2 10 11 3 3 13 4 7 4 10 9 1 10 10 11 13 1 10 9 3 0 2 7 3 0 1 15 15 3 13 3 1 13 2
10 10 9 2 3 2 13 13 1 9 2
6 10 9 13 10 9 2
12 10 9 1 10 9 7 1 10 10 0 9 2
34 1 15 13 10 9 13 1 9 1 10 9 1 10 9 3 0 1 10 9 0 2 11 13 10 9 1 9 1 10 11 2 11 2 2
47 2 15 13 15 1 10 9 1 10 9 2 2 13 11 2 15 13 10 9 0 1 11 1 10 9 1 10 11 1 10 11 7 10 0 9 2 15 3 13 13 3 10 10 9 1 11 2
36 13 1 13 1 10 9 11 1 10 11 1 12 2 11 2 1 12 9 2 13 1 1 10 9 1 10 9 13 10 0 0 9 1 10 11 2
7 2 13 9 10 9 10 2
38 3 13 1 13 0 7 0 2 7 13 16 10 9 3 13 16 13 1 10 9 2 2 13 10 9 1 10 9 0 2 1 15 13 10 10 0 9 2
4 9 1 10 11
6 9 1 9 0 1 9
23 10 9 13 1 13 15 2 9 1 10 9 2 2 7 10 9 1 10 9 1 9 3 2
27 3 12 9 1 10 9 0 13 13 1 9 2 13 10 9 1 10 11 2 11 2 2 3 13 1 11 2
40 10 9 1 10 2 11 2 1 11 2 11 2 13 13 1 9 1 12 9 1 9 7 12 9 1 9 1 13 13 10 9 1 10 11 2 13 3 10 11 2
32 10 9 13 13 1 12 9 2 13 1 10 9 1 15 13 3 1 10 9 7 1 13 13 2 10 9 1 15 13 13 2 2
39 10 9 13 13 1 2 1 9 13 1 9 1 12 2 13 13 10 9 1 10 9 1 10 11 2 9 11 7 10 9 11 2 9 15 10 11 13 0 2
52 3 1 10 9 2 11 13 13 2 9 3 2 1 10 9 2 1 9 0 1 13 0 0 2 2 1 15 15 13 13 1 10 9 13 2 0 16 2 1 10 9 1 9 1 10 9 2 15 13 9 2 2
34 1 9 2 10 9 13 3 13 13 9 1 13 2 2 7 3 3 1 13 2 2 3 13 2 13 10 9 7 9 1 15 13 2 2
68 10 9 13 2 3 2 16 10 9 1 11 2 13 0 7 3 0 7 0 1 13 3 10 9 1 10 9 1 10 2 3 10 9 1 10 10 0 9 2 1 10 9 7 1 10 9 1 15 13 3 9 2 9 7 9 1 10 9 1 10 9 0 3 15 15 13 2 2
23 1 9 1 10 11 2 11 13 16 15 13 1 13 2 0 9 1 9 15 3 13 2 2
3 7 13 2
16 2 16 3 13 1 4 7 4 15 15 13 2 3 13 2 2
9 9 1 0 1 10 2 9 0 2
21 10 9 13 3 16 10 9 1 10 9 1 10 9 0 2 13 15 1 13 2 2
37 13 1 10 11 1 10 11 2 15 13 1 10 9 1 11 2 11 13 16 2 10 9 1 9 13 13 15 3 7 10 9 13 1 10 9 2 2
51 13 10 9 1 10 9 1 2 13 10 9 0 0 7 0 1 10 9 0 7 0 2 7 3 13 1 10 9 2 13 13 1 10 10 9 1 10 9 2 9 7 1 10 0 9 1 10 9 0 2 2
25 1 13 10 9 0 2 11 13 16 10 9 0 1 10 9 0 13 13 9 0 2 13 7 13 2
14 1 15 2 13 2 2 13 10 9 1 9 0 2 2
4 11 13 11 3
53 10 9 1 10 9 0 13 3 10 9 2 16 15 1 10 9 15 13 9 1 10 9 3 1 10 9 1 10 9 1 9 13 3 13 1 10 9 1 10 10 9 3 13 1 9 10 9 15 13 1 10 9 2
29 13 3 1 10 11 2 1 9 2 13 1 10 9 1 10 11 1 10 9 1 10 11 7 13 12 2 9 2 2
17 13 3 10 9 0 0 2 1 9 0 7 9 0 1 9 0 2
16 7 9 2 16 13 2 3 13 2 2 15 13 1 10 9 2
13 3 15 13 3 3 2 9 1 9 2 1 11 2
8 15 13 10 0 9 15 13 2
56 1 10 9 2 0 7 0 9 1 12 9 2 1 9 0 13 15 10 9 1 2 11 2 1 11 2 11 2 2 2 11 2 1 11 2 11 2 2 2 11 2 1 11 2 11 2 7 2 11 2 1 11 2 11 2 2
29 10 9 2 9 1 9 0 9 13 3 10 9 1 10 9 0 11 2 1 10 10 10 11 13 13 12 9 10 2
41 10 12 9 1 11 13 0 1 10 9 2 13 2 10 0 9 1 12 1 10 9 0 3 0 2 3 0 2 13 3 0 9 1 10 9 2 2 1 13 11 2
29 3 11 15 13 13 1 10 9 0 1 2 11 2 1 11 2 9 13 1 10 9 11 2 13 1 10 0 9 2
57 2 1 10 9 1 12 7 12 2 10 9 0 1 11 13 10 9 0 7 9 1 9 0 2 1 10 9 1 10 9 1 9 15 13 10 9 1 10 9 1 9 0 7 1 9 3 1 10 9 1 10 9 0 1 10 9 2
62 3 2 10 9 13 1 0 9 1 9 2 3 1 10 9 1 9 1 9 15 10 9 3 13 2 1 13 13 1 10 9 1 9 7 10 9 13 1 13 2 1 10 9 2 10 0 9 0 1 15 13 13 10 9 1 10 9 2 2 13 11 2
64 10 9 0 1 10 9 2 9 2 2 10 0 9 1 9 1 10 0 9 2 10 9 1 9 7 9 1 10 9 0 7 0 2 10 9 0 7 10 9 7 9 0 1 10 9 0 1 11 2 9 13 10 12 9 1 9 2 13 10 9 15 11 13 2
79 10 9 2 15 13 13 10 9 1 10 9 1 11 12 9 1 10 9 0 0 1 10 11 2 13 3 12 9 2 13 10 2 0 9 2 1 10 9 0 2 10 11 2 7 10 11 2 11 2 13 16 2 1 11 13 15 3 7 13 15 3 2 2 1 10 9 1 10 9 1 10 11 7 10 9 1 10 9 2
5 3 3 15 13 2
21 3 13 16 10 9 13 3 13 1 10 9 11 3 15 13 16 13 1 9 0 2
32 15 15 13 2 13 11 2 15 13 10 9 0 1 10 9 13 3 12 9 2 13 16 3 13 9 13 10 9 1 10 9 2
23 2 3 0 10 9 13 1 10 10 9 2 3 0 10 9 13 13 2 2 13 10 9 2
18 15 16 10 10 9 13 3 10 9 1 9 1 10 9 1 10 9 2
37 3 10 9 13 1 10 9 1 10 9 13 2 9 0 12 2 13 3 0 1 12 3 1 10 10 7 10 9 1 9 1 10 12 9 13 0 2
21 2 10 9 15 13 10 9 1 10 9 13 3 13 0 1 13 10 9 1 9 2
18 1 15 2 13 15 3 13 2 1 10 9 3 0 2 2 13 11 2
6 2 10 9 13 3 2
42 10 9 2 11 2 2 13 1 12 1 9 0 2 1 10 9 15 13 1 13 13 1 10 9 2 11 2 7 15 13 1 9 13 1 10 11 13 15 10 0 9 2
60 2 10 12 9 15 13 10 9 3 2 11 7 11 2 13 2 1 10 9 1 10 9 15 13 3 2 16 10 9 1 13 1 15 12 1 10 9 15 13 1 10 9 15 15 13 2 15 11 2 9 0 2 10 11 2 9 1 9 0 2
9 2 15 13 9 2 9 7 9 2
28 1 9 1 12 13 13 12 2 12 2 9 2 1 15 15 13 13 3 1 15 13 1 10 9 1 10 9 2
66 1 10 9 2 3 13 2 3 9 2 1 10 11 2 1 10 13 9 2 10 10 9 1 2 9 2 2 2 9 15 13 15 1 13 2 2 2 0 2 2 7 10 9 1 10 2 9 2 3 9 1 13 1 15 13 1 9 2 9 2 1 10 0 2 0 2
51 1 9 1 9 1 10 9 2 1 10 9 11 2 13 13 1 10 11 10 9 3 1 9 1 10 11 2 10 9 13 13 13 15 1 10 0 9 7 10 3 0 2 13 1 10 2 9 2 1 11 2
36 3 1 15 2 3 1 10 9 1 11 2 13 4 13 3 1 9 10 9 3 13 1 10 11 2 1 15 15 13 15 1 10 11 7 11 2
44 3 1 15 2 10 11 13 13 10 9 1 10 11 2 1 10 9 11 2 1 10 0 9 1 10 11 13 11 2 10 0 9 1 10 11 2 7 9 1 10 12 0 9 2
69 1 9 1 9 2 9 1 9 2 13 13 12 0 9 1 10 11 15 13 13 10 9 3 13 1 2 11 2 2 3 12 9 0 1 10 9 2 10 9 13 11 1 10 9 13 1 10 11 2 7 3 12 1 9 2 7 3 12 9 1 10 11 1 2 11 2 1 11 2
54 10 9 1 10 2 9 2 2 15 13 12 9 2 10 15 1 2 9 2 7 13 1 12 9 2 1 10 0 7 10 0 2 2 13 1 10 9 11 2 0 1 10 9 0 1 10 9 11 2 0 1 10 11 2
38 3 10 9 1 10 9 0 2 15 15 13 13 1 12 9 2 10 9 2 10 0 9 7 10 2 9 2 2 13 3 1 13 1 15 13 4 13 2
30 2 13 1 9 1 10 9 2 1 15 10 11 2 7 3 13 3 9 13 1 15 1 15 2 13 1 10 11 11 2
34 10 11 13 16 10 9 7 10 9 1 9 13 13 10 0 9 2 9 7 9 2 1 10 9 2 1 15 13 1 10 9 1 9 2
11 10 9 13 3 0 2 16 13 1 15 2
36 16 13 13 2 9 0 2 1 10 11 13 15 1 13 12 1 9 2 10 15 16 2 3 2 1 10 11 2 11 2 11 2 11 7 11 2
29 3 16 13 13 2 3 1 9 0 2 1 11 2 11 2 11 2 11 7 11 2 10 9 1 9 13 1 12 2
45 10 11 9 1 10 11 13 3 1 11 7 13 4 1 13 2 1 10 9 7 1 10 9 2 1 10 9 1 11 1 11 1 3 12 9 1 9 15 3 13 13 1 10 11 2
59 1 10 10 9 1 11 2 10 9 0 9 13 12 9 9 2 12 9 7 12 9 2 15 13 1 9 1 9 1 11 2 1 10 9 13 1 10 9 1 10 9 1 9 2 11 2 15 13 10 9 1 10 11 1 11 2 11 2 2
8 11 13 15 1 10 2 11 2
37 10 9 1 10 9 13 13 9 1 10 11 1 10 9 2 11 2 2 15 3 13 1 0 9 16 2 11 13 12 9 1 9 1 10 11 2 2
54 3 1 10 9 0 13 1 10 9 1 11 2 10 13 9 13 2 3 0 7 0 2 16 2 10 9 3 13 9 1 10 9 2 2 7 13 10 9 1 10 9 1 10 9 0 1 10 9 1 9 1 10 9 2
78 1 9 13 2 16 15 13 3 12 12 9 1 9 0 2 1 9 2 1 10 10 9 1 9 2 13 15 3 12 12 2 10 9 15 15 13 1 10 9 2 12 12 9 1 11 1 9 2 0 2 1 3 12 12 9 1 9 3 1 2 0 2 2 2 1 10 0 9 13 13 3 1 10 9 1 10 0 2
13 10 9 1 10 10 9 13 1 3 13 3 3 2
22 13 3 16 10 9 2 15 3 12 12 2 15 13 1 10 9 1 3 12 12 9 2
22 10 9 3 13 13 15 15 13 1 10 9 1 10 9 13 3 1 0 9 1 9 2
34 13 10 9 3 1 2 11 2 2 1 11 2 15 3 13 1 9 1 9 2 10 9 1 9 13 1 10 9 1 12 12 9 2 2
19 10 9 1 9 1 10 11 2 11 7 11 3 13 3 12 9 1 9 2
16 10 0 9 0 15 13 10 9 13 10 11 1 2 11 2 2
32 10 9 1 9 1 10 11 3 3 13 9 1 9 2 7 3 3 13 1 10 9 1 10 9 2 16 3 15 13 1 9 2
19 9 2 1 10 9 1 15 13 2 13 1 13 1 13 13 10 9 0 2
4 9 2 13 2
8 9 2 3 13 10 10 9 2
24 13 10 9 0 3 10 9 2 7 2 16 3 15 13 2 15 3 3 13 1 15 10 9 2
10 11 0 13 13 1 13 9 1 10 11
8 9 13 1 10 11 1 10 11
15 10 11 1 10 11 13 13 1 13 10 9 1 10 11 2
12 1 10 9 2 3 10 9 0 1 10 9 2
19 7 10 9 13 3 4 13 10 9 13 1 10 9 1 15 10 9 13 2
14 9 0 13 15 3 7 13 10 9 1 10 0 9 2
13 13 0 9 2 0 9 2 0 9 2 0 9 2
6 3 2 10 0 9 2
17 13 13 1 13 1 15 2 7 13 13 10 9 1 12 1 9 2
69 1 10 9 1 9 0 1 10 9 1 10 9 0 2 2 11 2 2 9 11 2 12 2 2 11 2 2 9 11 2 12 2 7 2 11 2 2 9 11 2 12 2 1 13 13 10 9 1 10 11 2 15 13 1 13 10 11 2 2 11 13 15 3 1 11 1 10 9 2
8 13 1 12 2 1 10 11 2
53 3 1 13 11 7 11 1 10 11 2 13 15 2 1 12 2 1 10 9 2 11 2 2 2 13 13 2 1 11 2 11 2 11 7 11 2 12 1 10 9 15 3 13 13 1 16 11 3 13 1 10 9 2
28 13 1 10 11 2 10 9 13 13 13 10 9 2 1 10 9 15 3 13 7 13 2 10 9 2 3 2 2
22 15 13 2 1 11 2 10 9 10 1 3 15 13 2 3 0 2 1 10 9 13 2
60 3 3 1 13 4 13 16 2 1 10 9 1 10 9 1 3 2 10 11 13 12 9 2 10 11 2 1 12 9 2 10 11 2 1 12 9 7 10 11 2 1 12 9 2 2 10 9 1 10 9 0 1 10 11 1 13 1 10 9 2
9 2 13 3 1 13 1 10 9 2
9 3 13 1 10 9 2 13 11 2
31 7 10 11 2 1 12 9 2 7 3 9 1 10 11 2 13 16 10 9 2 13 3 10 9 15 3 13 1 13 2 2
25 1 10 9 1 10 9 2 11 2 13 15 1 13 16 2 3 15 13 1 9 1 10 9 0 2
11 13 9 0 15 3 13 1 10 9 2 2
28 7 1 10 0 1 10 11 2 11 2 10 9 13 2 13 3 9 2 3 3 13 1 10 9 1 9 2 2
22 10 9 13 1 15 1 10 9 0 1 10 9 1 10 9 3 1 10 9 1 11 2
18 2 13 9 15 3 13 1 10 9 1 9 16 3 13 9 0 2 2
25 3 2 13 3 13 10 9 1 15 13 13 7 3 13 2 1 15 2 1 13 9 16 13 13 2
21 2 13 16 3 16 10 9 3 13 10 9 2 2 13 2 1 9 2 10 9 2
16 11 2 3 13 1 13 10 11 2 1 12 2 13 10 9 2
17 3 16 15 2 13 13 1 10 9 1 13 1 13 10 9 3 2
8 3 13 1 9 1 10 9 2
12 9 2 13 9 1 15 2 16 13 1 11 2
10 13 15 1 10 9 0 2 3 13 2
5 11 2 13 2 9
51 10 9 0 11 13 1 10 9 2 1 9 0 2 1 10 9 1 11 2 1 11 2 1 10 9 1 0 9 13 7 0 2 10 9 3 0 1 10 0 1 10 9 2 10 9 2 13 2 11 2 2
31 2 13 10 9 13 3 1 15 2 13 10 9 1 10 2 11 2 2 15 13 13 1 10 11 2 10 3 0 9 0 2
45 16 10 2 9 2 13 10 9 1 9 7 1 9 1 9 2 1 15 10 9 2 1 13 3 10 9 1 10 9 2 13 2 3 1 15 2 10 9 1 10 9 1 10 10 2
33 3 10 9 1 10 9 13 1 10 9 2 13 9 1 9 15 13 10 9 1 10 9 0 1 10 9 1 10 9 1 10 11 2
49 2 7 10 9 1 10 9 2 2 13 2 10 0 9 1 10 9 1 15 15 13 10 9 1 10 9 15 3 13 10 9 1 10 9 0 2 1 10 9 2 1 10 9 0 7 1 10 9 2
12 10 9 1 10 2 9 2 13 3 12 9 2
21 13 16 2 1 10 0 9 2 10 9 1 9 0 13 1 10 9 0 7 0 2
35 10 9 1 10 9 13 1 13 1 10 0 9 1 10 11 2 2 10 9 13 1 10 11 2 2 16 10 9 13 0 1 10 9 3 2
29 10 9 1 10 11 2 3 1 13 10 9 15 10 0 11 13 1 10 9 2 3 13 10 9 1 10 9 0 2
35 10 9 1 10 11 13 1 10 9 1 10 9 1 10 9 2 1 10 9 2 16 10 0 9 13 1 10 11 3 13 3 10 9 0 2
42 7 10 9 1 10 11 2 13 10 0 9 16 10 9 0 1 10 9 13 10 9 0 7 16 10 9 0 15 13 2 3 2 3 2 10 9 15 13 1 10 9 2
20 10 9 1 9 13 13 2 3 2 10 9 0 1 10 11 1 10 0 9 2
46 1 1 10 9 2 10 9 1 9 1 10 11 2 13 16 10 10 9 0 13 13 15 3 0 2 2 13 11 2 13 10 9 1 10 9 0 15 13 1 10 9 0 1 10 9 2
22 1 15 2 10 11 13 1 13 10 2 0 9 2 1 10 9 0 2 13 10 9 2
50 10 9 1 10 11 1 10 9 13 3 10 9 0 1 10 9 1 10 9 13 1 10 9 2 3 10 1 10 9 0 2 15 13 10 15 13 3 13 9 1 9 2 2 3 12 9 1 10 9 2
31 10 9 13 13 2 3 2 10 9 1 9 2 10 9 1 9 2 9 2 7 10 9 1 9 15 13 10 9 3 0 2
23 11 2 9 1 11 1 10 11 2 11 2 2 13 10 0 9 1 10 9 0 1 9 2
34 13 1 10 11 2 10 9 13 1 10 9 12 1 12 9 0 1 11 0 2 12 1 10 11 2 12 1 10 11 7 15 1 11 2
23 2 1 3 12 9 1 10 9 2 3 1 12 1 12 9 15 13 13 10 9 0 2 2
14 9 15 13 10 11 1 13 10 9 1 12 9 0 2
35 12 1 10 9 0 2 1 9 1 9 1 12 7 12 2 13 12 12 9 2 13 12 9 2 12 1 10 9 7 12 1 10 11 2 2
13 1 10 9 2 13 3 1 12 9 1 10 9 2
23 10 9 13 3 2 16 10 9 0 3 13 9 1 9 0 1 12 1 10 9 1 11 2
11 2 1 12 2 13 10 9 1 9 13 2
14 1 10 9 0 13 15 9 1 9 0 1 12 2 2
26 10 0 9 0 2 15 13 13 1 10 11 1 12 7 12 2 13 12 9 7 13 3 12 12 9 2
20 10 11 13 10 9 1 10 11 2 15 13 2 3 1 10 9 1 10 11 2
4 13 3 0 2
50 10 9 7 9 13 1 10 9 1 10 9 1 10 9 2 13 2 12 2 10 9 1 10 9 9 2 1 10 9 1 10 11 1 1 11 2 1 10 9 2 1 15 3 13 10 9 1 10 9 2
5 12 9 3 13 2
6 10 9 3 13 13 2
30 1 10 9 2 10 9 13 1 10 9 0 1 10 9 13 13 1 9 2 15 13 10 0 9 3 1 10 10 9 2
24 15 13 1 3 13 13 3 10 2 9 2 1 10 9 2 16 15 13 12 1 1 10 9 2
16 7 3 13 1 15 13 1 10 9 2 15 15 13 15 12 2
11 3 2 10 9 1 9 13 15 10 9 2
9 3 13 10 0 16 3 13 9 2
10 16 10 9 2 10 9 2 15 13 2
2 0 2
18 7 2 1 3 15 13 9 2 16 15 13 2 10 9 13 3 0 2
13 13 3 0 16 10 9 15 15 13 15 13 11 2
7 11 2 13 3 1 13 2
6 13 15 16 10 9 2
28 1 10 0 9 2 10 10 9 13 15 1 10 9 15 13 1 10 0 9 2 1 9 2 0 9 2 9 2
35 1 10 9 3 13 1 10 9 1 10 9 2 15 3 3 15 13 13 1 16 10 0 3 3 13 3 10 0 2 13 3 10 9 0 2
43 3 2 3 1 10 9 2 3 13 1 4 1 10 9 7 4 1 10 9 1 10 11 7 1 10 9 1 11 2 3 13 9 13 2 3 2 3 13 3 1 13 11 2
11 9 2 3 13 3 13 10 9 1 11 2
13 10 9 13 9 2 3 2 1 9 7 9 0 2
38 3 2 3 2 1 9 1 10 11 2 11 2 9 2 13 1 9 1 11 2 1 10 0 9 2 1 10 9 1 10 9 13 1 11 1 10 9 2
57 13 9 1 10 9 1 10 9 15 13 10 9 1 10 11 13 10 11 1 10 9 1 10 9 1 9 2 11 2 13 10 9 1 10 11 2 13 13 3 2 16 2 13 2 2 10 9 1 10 3 15 13 1 10 11 2 2
31 3 16 11 2 1 10 9 1 11 2 3 13 2 0 9 2 7 2 0 2 2 13 1 15 4 4 2 13 3 2 2
41 3 2 11 13 15 1 10 9 13 1 10 11 2 1 10 9 1 10 9 1 11 2 1 15 13 16 10 0 9 2 1 11 3 13 2 9 1 10 11 2 2
3 2 1 11
2 11 2
28 3 2 1 10 9 2 3 2 1 10 9 7 1 10 9 2 9 2 1 10 9 2 9 2 1 10 9 2
2 11 2
9 9 12 7 12 2 1 10 9 2
51 10 11 13 13 1 13 10 10 9 0 1 11 2 1 13 10 9 7 10 9 0 0 2 1 10 9 1 13 1 10 9 1 16 10 9 15 13 1 10 9 1 9 1 9 2 13 3 10 9 11 2
39 9 1 10 11 0 13 16 10 11 13 1 10 9 1 10 9 1 10 9 0 1 10 9 1 9 1 10 11 2 3 1 10 9 1 10 9 1 9 2
41 10 9 13 16 10 0 13 16 10 9 13 10 0 9 1 10 9 13 1 10 9 1 10 9 2 13 1 10 9 1 10 9 1 11 2 13 15 1 10 9 2
55 10 9 13 2 16 10 9 0 1 10 11 3 15 13 13 2 16 10 11 0 13 0 1 2 2 3 1 10 11 2 2 13 9 1 16 11 13 10 10 9 1 9 1 9 0 2 13 1 13 3 1 10 9 0 2
4 9 13 7 13
36 10 9 1 12 9 10 9 13 13 1 10 9 13 13 1 10 9 1 10 12 9 7 13 1 10 11 1 11 2 11 2 13 3 9 0 2
43 11 13 1 10 9 2 9 2 1 10 9 1 11 2 1 12 9 1 10 9 0 1 11 2 1 10 11 2 3 13 13 1 10 9 7 15 13 10 9 1 10 9 2
24 10 9 1 10 9 13 10 9 15 15 13 1 10 9 0 2 1 9 1 9 7 13 3 2
14 7 10 9 13 1 9 1 13 2 2 13 0 2 2
22 13 1 9 1 11 1 10 9 1 10 9 13 1 9 2 13 3 13 1 12 9 2
37 3 2 13 15 13 3 10 9 0 15 1 3 13 9 2 9 2 9 7 10 9 1 0 9 2 13 9 1 10 0 15 13 3 1 10 9 2
47 7 10 9 13 1 13 2 3 2 15 1 10 9 3 0 1 10 9 0 0 7 10 9 0 2 15 3 10 1 11 2 15 15 13 13 13 1 10 9 7 10 9 1 10 9 0 2
3 9 1 9
82 10 9 0 1 3 2 1 15 13 12 9 2 7 10 9 0 15 15 15 13 13 1 16 9 0 13 13 10 9 1 10 11 2 10 0 11 2 1 12 9 2 7 15 1 10 11 2 10 9 11 2 1 12 2 13 3 1 13 10 9 1 3 12 9 2 11 2 7 1 10 9 1 9 1 10 11 2 11 2 10 9 2
37 1 13 10 9 1 10 9 0 1 10 9 2 10 9 13 2 16 15 13 1 10 0 9 1 13 2 10 9 1 9 1 9 15 13 10 9 2
27 10 9 3 13 12 1 10 9 1 10 9 7 13 15 1 9 1 10 9 1 10 9 13 1 10 9 2
48 16 10 9 13 3 0 1 10 10 9 13 13 1 10 11 2 3 1 10 9 3 0 2 10 9 13 1 13 2 9 2 1 10 9 1 2 1 3 2 13 10 2 9 2 1 10 9 2
36 10 9 1 9 2 13 10 9 0 1 15 1 12 2 9 2 1 10 9 1 10 9 1 10 11 2 2 13 10 9 3 13 1 10 11 2
34 1 10 9 2 2 10 9 1 10 11 3 13 13 9 1 9 1 10 9 2 2 7 2 13 10 9 1 10 9 15 13 9 2 2
29 7 13 3 16 10 9 1 10 11 1 9 2 13 1 11 2 2 13 10 9 0 1 10 9 1 10 11 2 2
38 10 9 13 10 10 9 0 1 11 3 13 2 10 0 2 7 13 3 13 10 9 1 10 9 0 2 16 2 10 9 13 1 13 10 10 9 2 2
42 13 3 16 10 10 9 1 11 13 1 10 9 0 1 10 9 0 2 3 10 11 13 1 10 9 2 15 13 4 13 1 10 11 2 15 13 13 1 10 9 0 2
5 9 1 11 1 11
2 13 13
36 10 9 1 10 9 7 10 9 1 10 9 1 11 1 10 9 1 10 9 13 10 9 1 10 9 1 12 9 2 1 13 3 2 1 11 2
33 13 1 10 11 2 1 9 1 10 11 2 10 9 13 1 10 9 1 9 1 10 9 0 1 9 1 11 7 1 10 0 9 2
4 11 13 9 0
50 10 11 13 13 1 10 9 1 10 11 10 9 15 13 1 12 9 10 9 0 2 13 1 16 2 1 12 2 10 9 2 1 13 12 9 1 10 9 1 10 9 0 2 13 1 13 1 12 9 2
30 10 9 2 3 13 1 10 11 0 2 13 1 13 13 10 12 9 0 2 11 2 11 2 11 2 11 7 11 2 2
45 10 0 0 1 10 9 1 9 1 9 2 11 2 13 16 10 11 2 11 2 2 10 9 1 9 1 13 10 9 0 1 10 9 1 12 9 2 13 0 1 13 13 1 9 2
11 7 15 2 1 0 9 2 13 1 9 2
44 1 10 9 0 1 10 9 0 2 11 2 13 15 1 10 11 13 2 1 10 9 1 12 9 2 1 10 2 9 13 1 9 2 7 10 9 3 13 10 9 1 10 11 2
33 2 10 9 3 15 13 1 10 9 2 2 13 3 11 2 13 15 1 10 9 0 13 1 10 11 1 10 11 2 11 7 11 2
10 2 10 10 9 0 13 12 9 0 2
8 15 13 13 10 10 9 2 2
5 9 0 1 10 11
37 10 9 1 0 9 13 3 2 1 10 9 2 1 10 9 1 10 11 2 1 11 2 1 10 9 1 9 13 1 10 9 0 1 10 9 11 2
20 0 1 10 9 0 1 10 9 1 10 9 2 11 13 0 1 0 1 9 2
39 10 2 9 11 2 2 10 9 1 10 9 1 11 1 10 9 15 3 13 10 9 1 10 11 2 3 13 2 3 2 10 9 0 15 10 9 0 13 2
40 3 15 13 10 9 1 10 2 0 9 0 2 2 3 0 2 12 1 10 9 1 10 10 9 2 16 3 13 13 1 12 13 1 10 9 0 1 9 0 2
25 10 9 2 1 10 9 1 10 9 7 10 9 13 1 10 9 0 2 13 15 9 1 10 9 2
28 10 0 9 13 13 1 10 9 1 10 0 9 0 2 1 10 11 13 1 10 9 1 10 9 1 10 9 2
3 10 0 9
18 10 9 0 11 13 2 1 10 9 2 12 1 10 10 3 13 9 2
29 15 16 10 9 11 2 1 9 3 9 3 13 10 9 2 13 10 9 13 10 9 1 10 9 1 10 9 0 2
10 13 12 9 1 10 9 1 10 9 2
13 13 15 3 9 7 9 0 2 3 15 13 3 2
8 13 1 13 15 1 10 9 2
8 13 15 10 9 1 10 9 2
3 13 15 2
5 13 4 13 9 2
5 11 13 10 9 2
4 13 10 9 2
3 13 9 2
13 13 1 10 9 7 1 10 9 7 13 15 3 2
21 3 3 13 16 13 10 9 16 10 9 13 1 10 9 1 10 9 15 3 13 2
4 3 2 13 2
38 11 13 13 10 2 9 1 10 9 2 7 13 1 10 10 9 2 11 2 16 1 10 9 1 11 1 11 2 10 9 13 1 10 9 1 10 9 2
6 13 10 2 9 2 2
10 10 9 2 15 2 13 1 10 9 2
19 12 9 7 9 1 9 1 13 2 13 7 13 10 9 13 1 10 11 2
45 3 1 10 9 2 1 10 9 0 1 11 2 10 9 13 15 1 10 9 7 13 15 1 13 2 11 2 2 2 11 2 2 2 11 2 2 3 13 0 10 9 1 10 11 2
22 9 7 9 1 10 11 13 2 13 1 10 9 7 9 13 15 13 9 10 9 13 2
20 13 15 10 9 11 7 10 9 15 11 13 1 10 9 1 10 2 11 2 2
29 11 2 9 1 10 9 15 13 13 1 11 2 13 13 1 13 10 9 13 3 1 10 9 0 13 1 10 11 2
12 9 0 2 7 15 13 13 10 9 1 9 2
10 2 13 1 10 10 9 1 11 2 2
31 3 2 1 10 9 1 9 7 9 2 13 15 2 11 2 2 10 9 13 7 13 1 10 0 1 10 12 9 1 9 2
11 2 13 7 13 15 1 10 9 1 9 2
8 2 2 2 12 12 3 13 2
3 2 13 2
3 2 13 2
7 13 10 10 9 2 2 2
22 1 10 9 1 10 0 9 2 10 0 9 13 1 9 13 7 13 13 1 10 9 2
4 9 1 13 9
47 10 9 0 0 11 13 1 10 9 1 10 11 1 13 3 9 1 10 11 1 10 9 1 13 10 9 1 10 9 0 1 11 2 13 1 10 11 7 13 0 1 10 9 0 7 0 2
31 10 12 9 3 1 9 1 10 9 2 1 12 9 15 2 13 4 1 12 7 12 7 4 3 1 10 9 1 10 11 2
10 12 1 15 13 1 10 9 3 13 2
9 2 3 3 13 10 10 9 9 2
12 13 1 15 9 1 9 13 2 2 13 11 2
40 3 10 9 1 9 1 11 7 10 11 13 2 10 9 13 1 13 10 9 1 10 11 2 3 9 0 13 3 3 12 9 1 9 0 1 10 9 1 9 2
22 1 10 9 1 10 9 1 10 11 2 11 2 1 10 9 0 2 13 13 10 9 2
29 1 10 9 0 1 10 9 1 10 11 2 1 10 9 1 11 2 11 2 13 12 9 0 7 15 12 13 13 2
23 11 3 13 1 11 3 1 13 10 9 1 10 11 1 15 13 13 3 1 10 9 11 2
35 10 9 0 1 10 11 2 15 3 13 1 13 10 0 9 1 9 0 1 11 2 13 1 15 10 9 3 0 1 13 1 10 9 0 2
32 12 9 3 1 10 0 9 1 11 1 10 11 2 13 10 9 1 13 1 13 10 9 1 10 9 1 10 11 1 10 9 2
78 10 9 1 10 9 1 2 9 0 2 1 10 9 1 10 11 3 13 3 1 10 9 15 10 9 0 13 1 10 9 1 10 11 1 11 7 1 11 2 11 3 13 13 10 9 1 10 9 15 13 13 1 10 11 9 3 1 15 13 10 9 1 11 2 2 7 10 0 13 16 10 11 0 13 10 9 0 2
14 3 1 15 13 3 11 13 3 3 13 1 10 10 9
41 1 10 0 9 15 13 1 10 11 15 15 13 1 13 10 11 1 10 9 1 10 0 9 0 7 15 15 13 16 13 13 2 3 3 2 10 9 2 11 13 2
15 2 15 15 13 13 10 9 1 10 9 13 10 9 2 2
28 15 13 10 13 9 1 10 9 0 2 11 2 1 10 9 1 10 11 2 3 10 9 1 9 1 10 11 2
32 7 2 13 2 2 10 9 7 10 9 1 10 9 3 13 4 13 1 10 9 1 15 13 2 7 1 15 1 10 9 2 2
17 1 10 13 9 0 2 1 11 13 10 9 1 9 3 3 13 2
40 1 10 2 9 2 13 1 10 9 15 13 16 13 7 3 13 2 10 9 1 9 13 1 13 1 10 9 1 10 9 7 13 1 15 2 1 9 1 9 2
22 2 13 15 0 2 2 13 9 1 10 9 2 2 13 1 10 9 1 10 9 2 2
6 2 11 2 13 1 11
19 15 3 13 1 10 9 1 11 2 11 2 13 3 1 13 1 10 11 2
33 2 11 2 2 3 15 15 13 2 13 12 9 7 13 1 10 9 2 1 10 9 1 10 9 2 1 9 1 10 13 9 0 2
45 1 12 9 3 2 11 2 13 15 9 1 10 9 15 13 1 10 9 1 9 7 1 9 2 1 10 9 1 10 11 7 11 2 7 1 10 9 0 1 15 15 13 1 15 2
7 11 13 1 11 2 12 2
4 11 13 10 9
25 11 13 10 9 1 10 9 1 3 1 10 11 7 10 11 1 15 13 12 9 1 10 9 0 2
35 11 13 1 13 10 9 0 2 1 15 13 2 1 10 0 9 7 1 10 9 1 9 2 10 9 15 13 10 9 1 10 9 1 11 2
20 1 10 9 13 2 10 9 13 1 13 1 10 9 2 1 10 9 1 9 2
9 7 13 2 7 3 2 13 15 2
17 10 11 13 12 1 10 9 1 9 1 0 9 1 10 10 9 2
12 13 3 16 10 9 13 2 1 10 10 9 2
5 2 3 13 2 2
13 10 2 9 2 1 10 9 3 13 1 9 0 2
21 15 13 1 10 9 2 13 1 10 9 0 7 13 1 10 9 15 13 3 9 2
8 10 0 13 2 13 15 2 2
8 10 9 13 3 13 1 15 2
4 9 12 2 9
31 10 11 2 3 2 13 13 10 9 1 10 2 9 0 1 10 0 9 1 9 7 9 2 1 10 9 15 1 15 13 2
23 15 3 2 3 13 13 9 0 2 13 15 1 10 9 1 10 2 9 0 1 9 2 2
30 1 10 9 1 10 9 0 2 10 9 13 13 9 1 10 9 1 10 9 0 2 0 2 0 7 1 9 1 9 2
23 3 15 13 10 9 1 10 9 0 2 16 2 15 15 13 2 13 13 10 10 0 9 2
2 12 9
49 1 15 13 1 10 9 2 13 10 9 13 1 9 0 7 0 2 13 1 12 9 1 10 9 2 11 13 12 7 12 9 7 13 1 10 9 2 16 10 10 9 13 10 9 1 9 1 9 2
38 13 15 16 2 1 10 9 2 11 15 13 1 9 2 16 3 13 10 9 7 13 10 9 1 10 9 2 1 3 13 1 10 0 9 1 10 9 2
46 7 3 10 9 13 15 2 13 10 9 1 10 9 0 2 3 0 16 15 2 10 9 1 9 0 7 0 3 9 1 9 15 13 13 1 10 9 2 1 9 9 7 1 10 9 2
51 10 9 1 15 13 1 10 9 7 3 13 1 10 9 1 10 9 2 1 15 13 1 9 10 9 13 7 0 1 11 2 15 3 13 13 12 7 15 9 2 13 2 2 3 15 3 2 7 3 13 2
16 1 12 9 2 11 13 1 4 13 3 1 9 1 10 9 2
13 1 10 9 1 10 10 9 0 2 10 9 0 2
17 13 10 9 0 13 13 1 10 9 12 9 1 12 9 1 13 2
5 7 13 13 15 2
49 13 3 0 16 15 13 1 10 0 9 2 1 10 9 3 2 13 10 9 2 10 9 13 1 10 9 1 10 11 10 9 1 9 2 7 13 16 1 15 13 2 1 15 7 1 9 0 2 2
24 11 3 13 1 9 1 12 9 2 3 12 9 2 2 1 10 10 9 0 1 13 12 9 2
37 10 9 9 13 13 1 10 9 1 9 1 11 7 1 10 9 1 10 9 0 2 15 13 10 9 1 10 9 1 10 9 1 10 9 0 11 2
14 10 9 1 9 1 10 9 1 3 12 9 1 9 2
31 1 11 2 13 15 10 9 1 12 9 2 1 10 9 11 1 13 1 12 9 2 1 10 9 15 13 11 1 10 9 2
44 1 10 9 0 2 11 13 10 9 7 2 1 10 9 1 10 9 2 10 9 13 1 10 9 0 2 1 10 9 11 1 13 12 9 1 10 9 1 10 9 1 10 9 2
10 10 9 1 10 10 9 13 10 9 2
25 1 11 2 3 2 13 10 9 7 10 9 11 13 12 9 0 2 1 10 9 0 1 12 9 2
11 11 3 13 1 10 9 9 1 12 9 2
40 11 13 10 9 1 10 0 1 10 9 1 10 9 1 9 1 10 9 7 13 16 10 0 9 2 13 2 1 10 0 2 10 9 0 1 10 9 0 2 2
42 1 10 0 9 15 13 1 10 0 9 15 15 13 1 10 9 1 10 9 2 11 3 13 9 1 13 1 10 9 1 10 0 9 13 2 3 2 13 1 10 9 2
15 2 10 9 3 0 13 3 1 10 9 1 13 10 9 2
37 3 13 1 11 2 3 13 11 11 2 9 2 15 13 1 10 0 9 2 2 13 3 1 13 3 1 10 11 0 2 3 1 10 9 1 13 2
18 3 2 13 15 13 1 13 10 10 10 0 9 16 10 9 3 13 2
4 11 13 4 13
31 11 2 1 12 9 2 13 10 11 1 10 10 9 1 10 11 1 10 0 9 1 10 11 2 11 2 13 1 10 9 2
18 11 2 1 10 11 2 13 10 0 9 1 10 9 2 1 12 9 2
19 10 11 13 10 10 0 9 1 10 9 7 13 1 0 9 1 10 11 2
18 1 10 11 2 3 3 13 10 9 1 10 9 7 13 1 12 9 2
3 11 13 11
26 10 11 13 13 1 12 12 11 1 10 9 1 11 2 15 13 12 9 1 9 7 13 13 1 11 2
30 1 10 9 13 1 10 9 2 15 13 10 9 1 9 7 13 13 1 12 2 10 9 13 13 3 12 9 1 9 2
32 16 10 11 2 15 3 13 10 9 1 9 1 10 9 2 13 1 10 9 1 10 9 2 15 13 10 9 1 12 12 9 2
25 11 13 1 11 10 10 0 9 1 10 9 2 15 13 13 1 10 11 3 10 0 1 10 9 2
8 3 12 9 13 1 9 0 2
39 10 9 13 1 10 9 1 10 9 2 13 1 10 9 1 10 9 2 13 1 10 9 7 2 1 12 9 0 2 13 10 12 9 9 2 11 7 11 2
19 3 2 1 10 9 1 11 13 1 9 0 3 1 0 9 1 10 9 2
29 3 1 10 9 2 15 13 12 9 2 11 7 11 13 1 13 10 9 1 10 0 9 2 15 1 12 9 0 2
18 10 12 9 13 1 13 1 10 9 2 3 15 1 0 9 1 9 2
2 11 9
16 2 11 2 13 3 10 9 1 10 9 0 1 10 9 11 2
37 0 2 0 2 0 7 0 2 13 1 2 11 2 13 2 1 9 2 10 9 2 10 9 1 15 15 2 1 15 2 13 15 1 10 10 9 2
16 10 9 0 1 10 9 2 10 9 2 13 1 12 12 9 2
27 1 10 9 1 11 2 11 2 2 10 9 1 2 11 2 13 1 10 9 3 2 1 10 9 1 11 2
18 10 9 2 13 1 12 2 13 12 9 1 10 9 3 1 13 13 2
8 9 0 1 10 9 1 10 11
24 12 9 1 9 1 10 9 1 10 11 13 4 3 13 2 13 10 9 1 10 11 1 11 2
26 12 1 10 9 13 13 1 10 9 1 9 2 1 16 10 9 0 1 9 15 13 13 1 10 9 2
28 10 9 13 4 13 1 10 9 1 9 7 9 13 7 13 4 4 13 3 1 10 9 1 10 9 1 9 2
39 10 9 1 10 11 13 1 10 11 16 2 10 9 13 13 3 1 9 2 2 13 3 10 9 1 9 1 10 9 13 1 10 9 2 15 13 1 9 2
37 13 3 3 13 10 9 1 10 9 1 10 11 7 10 11 2 1 15 13 0 10 9 1 10 9 0 1 10 1 0 9 2 13 1 10 11 2
10 10 0 9 13 13 1 9 1 9 2
25 11 13 13 16 15 13 3 1 10 9 1 11 2 7 3 10 9 0 13 15 10 9 13 13 2
16 10 12 9 0 1 9 1 10 0 9 1 9 3 13 0 2
25 10 9 11 13 10 0 1 13 1 9 2 13 1 10 0 9 1 10 9 9 0 1 10 9 2
16 13 15 12 2 15 3 15 13 2 7 3 3 13 10 9 2
12 10 9 2 3 0 2 13 3 10 0 9 2
45 1 10 0 13 1 12 9 1 10 10 9 0 2 12 2 1 12 2 7 3 1 10 0 9 2 10 9 3 13 12 2 15 13 3 3 16 9 2 1 12 2 7 3 13 2
9 13 0 12 1 13 1 10 9 2
16 15 13 1 9 13 11 2 11 2 2 1 10 9 1 9 2
29 13 10 9 12 7 13 1 10 9 11 2 9 2 7 1 10 9 11 2 10 9 0 2 9 2 2 1 9 2
10 1 9 2 3 2 15 13 1 9 2
38 1 10 0 9 13 1 10 9 1 10 12 9 1 13 1 10 9 7 13 10 0 0 9 1 10 9 11 15 1 10 9 0 2 1 9 1 9 2
7 13 10 9 11 1 9 2
14 13 10 0 9 1 13 13 10 0 9 0 1 12 2
7 1 3 13 9 10 11 2
18 10 11 2 11 2 9 2 3 3 13 1 10 9 13 1 10 11 2
25 0 10 13 1 13 16 10 9 13 13 1 9 2 1 13 13 3 2 2 1 3 13 9 2 2
17 10 9 13 13 2 3 13 2 1 10 9 1 10 9 2 11 2
1 11
5 13 1 10 10 9
15 12 9 1 10 9 13 1 10 9 13 1 10 9 3 2
4 9 0 1 11
45 10 11 2 11 2 13 1 10 9 1 10 9 10 9 1 10 11 2 3 1 10 9 1 11 1 11 2 13 9 1 10 9 1 11 2 13 10 11 3 1 9 0 1 11 2
27 11 13 9 0 1 10 11 1 12 7 13 13 1 11 1 10 9 1 10 10 9 0 1 10 9 0 2
17 10 9 13 13 1 11 2 9 1 10 9 9 7 10 0 9 2
40 10 9 2 11 2 13 13 1 10 9 0 1 11 2 3 1 10 10 9 0 2 2 13 9 2 1 10 9 1 11 2 13 13 12 9 2 1 12 9 2
70 3 2 3 2 10 11 2 13 1 10 9 13 1 3 0 1 10 15 15 13 13 1 10 9 1 9 1 10 9 0 2 13 10 0 9 0 1 9 1 9 1 9 2 13 13 9 1 10 9 0 1 15 13 13 10 10 9 2 1 10 9 1 10 9 1 10 2 11 2 2
4 11 13 9 0
15 11 2 7 10 9 0 3 13 9 0 1 10 0 9 2
5 11 2 1 9 2
45 7 3 13 3 9 2 16 10 9 15 13 1 10 7 1 15 9 3 1 10 9 2 13 1 4 13 10 9 1 9 1 10 9 13 10 9 15 15 13 16 13 4 13 3 2
12 7 10 9 1 9 13 13 13 3 12 9 2
27 13 1 13 0 10 9 13 15 1 10 9 1 15 13 1 9 1 12 9 1 12 1 10 9 1 9 2
20 3 13 13 3 2 1 9 0 7 1 9 2 1 10 9 3 13 13 9 2
16 10 9 0 3 15 13 1 10 9 1 11 2 11 7 11 2
33 2 15 13 1 3 13 9 1 9 2 13 1 13 15 13 10 9 7 1 13 3 1 10 10 9 2 3 13 10 9 13 2 2
7 13 1 10 9 13 10 9
60 2 15 2 1 11 2 3 13 16 13 13 9 1 11 2 15 3 13 10 10 9 2 16 10 9 13 15 15 13 2 2 13 1 10 11 11 2 2 16 13 10 9 0 7 3 13 9 2 3 3 10 9 2 15 13 10 9 0 2 2
30 3 1 10 9 0 3 10 9 2 1 9 12 1 10 9 0 3 0 1 11 2 13 10 9 1 10 12 9 0 2
35 11 13 3 3 10 11 1 11 2 10 0 9 1 11 2 1 10 11 1 12 2 13 0 2 2 7 3 13 15 13 13 3 12 9 2
49 2 10 9 1 11 13 0 7 3 0 1 15 2 2 13 2 13 9 1 9 1 9 15 2 1 10 0 12 9 2 1 9 7 9 1 10 9 1 11 2 13 9 1 10 9 1 9 0 2
48 3 1 9 1 10 11 2 10 9 13 13 1 12 1 12 9 2 13 3 1 13 10 9 2 13 1 11 2 2 10 9 7 10 9 13 1 10 9 1 10 11 2 3 13 9 12 9 2
12 10 0 13 10 0 15 3 13 1 10 11 2
18 3 2 13 15 3 13 10 9 1 10 11 2 15 13 12 1 12 2
11 10 10 9 2 13 11 2 13 13 3 2
5 11 2 11 13 3
31 10 11 13 3 10 9 1 10 11 2 11 1 3 2 1 10 9 1 10 11 2 13 3 9 1 10 9 1 10 11 2
38 10 9 1 10 9 2 1 10 0 9 1 10 9 0 7 13 1 13 9 1 10 9 1 10 9 1 10 9 11 2 13 0 1 10 9 1 11 2
23 10 9 13 1 10 9 7 10 9 2 10 0 13 1 10 11 2 1 13 10 9 0 2
2 9 0
11 2 13 9 7 9 2 10 9 0 2 2
28 3 1 9 1 10 10 2 10 9 1 10 10 9 0 13 10 9 0 15 13 10 9 7 10 9 3 13 2
70 10 0 9 2 13 3 10 9 0 7 10 9 0 7 0 1 11 2 13 15 10 9 1 10 9 3 10 9 1 10 9 0 13 10 9 0 1 10 15 13 0 2 7 3 15 9 1 10 9 0 2 7 15 15 13 0 2 3 0 1 10 9 15 13 9 0 1 9 0 2
49 13 15 1 10 9 3 0 2 16 2 1 10 9 0 15 0 2 10 9 13 13 10 9 1 13 10 0 7 0 9 1 9 2 9 0 7 9 0 2 3 16 15 13 16 13 0 7 0 2
26 10 9 0 13 3 1 9 0 7 2 0 7 3 2 9 0 15 13 1 10 9 1 9 1 15 2
12 2 10 9 1 15 2 3 9 1 10 9 2
35 1 10 9 1 10 11 1 15 10 9 1 10 9 7 9 13 10 9 1 9 1 10 9 0 2 13 10 9 1 10 9 13 1 9 2
13 3 10 9 11 2 11 13 15 1 13 10 9 2
27 7 16 10 9 13 13 10 9 1 10 9 1 10 9 2 10 9 13 0 2 3 1 9 3 1 9 2
22 10 9 0 3 13 13 13 11 7 13 10 9 1 10 11 7 1 10 10 0 9 2
20 3 3 13 4 1 13 10 9 1 10 9 1 10 9 13 10 9 13 15 2
30 3 13 3 13 16 10 10 9 13 1 10 9 1 9 9 13 16 10 9 13 13 1 10 11 1 9 2 3 9 2
46 10 0 9 1 12 9 13 3 1 9 1 11 7 1 10 11 2 3 1 10 9 1 10 9 1 10 9 2 13 13 1 10 11 1 10 9 7 13 10 9 13 1 10 9 0 2
27 13 15 1 10 0 1 12 9 2 15 13 13 10 9 7 10 9 1 10 9 13 1 10 9 1 9 2
38 10 9 13 3 3 1 10 9 1 10 9 1 9 1 10 9 1 9 1 9 2 3 13 2 7 13 1 13 10 9 1 9 0 13 1 10 11 2
32 10 9 1 10 9 13 2 1 9 2 1 10 9 7 1 9 1 15 10 0 13 1 10 9 13 10 11 1 10 10 9 2
14 3 13 13 10 9 1 10 9 1 9 7 9 13 2
6 9 1 11 13 1 11
39 10 12 9 1 10 9 1 10 9 1 10 11 1 11 2 13 1 10 9 1 3 2 13 13 3 12 9 3 1 10 11 2 1 10 9 2 1 11 2
26 10 10 9 13 13 1 10 12 9 13 1 11 1 10 9 12 1 9 7 10 9 1 10 0 9 2
25 10 11 13 16 10 9 15 13 1 10 9 11 2 9 15 15 13 1 13 13 10 9 3 13 2
17 13 3 1 11 2 10 9 2 1 12 7 12 9 2 13 13 2
19 1 10 12 9 2 3 13 1 9 1 9 2 13 13 3 12 12 9 2
9 10 9 1 15 13 13 3 13 2
5 9 1 9 1 11
23 1 9 1 10 9 13 2 3 12 9 1 9 2 13 4 13 1 10 9 2 9 2 2
18 1 10 2 9 2 1 10 11 2 13 10 12 9 1 9 1 12 2
46 2 10 9 13 3 13 1 10 9 1 10 9 1 9 2 1 10 9 1 10 9 1 10 9 13 1 9 1 9 7 1 10 9 1 10 0 9 1 9 2 2 13 10 10 9 2
1 11
5 3 13 10 9 2
40 10 9 0 11 2 11 2 9 2 7 11 2 11 2 0 2 13 3 10 9 1 9 1 10 11 2 13 13 10 9 13 1 13 10 9 1 10 12 9 2
28 10 9 13 1 10 9 1 10 9 15 13 1 10 9 1 10 9 7 15 3 13 3 10 9 1 10 9 2
23 10 9 13 13 13 3 10 10 9 15 2 13 15 2 13 13 1 10 9 1 10 9 2
33 2 13 1 9 1 10 0 9 1 10 9 2 3 13 10 9 0 2 2 13 11 7 11 1 10 9 1 9 0 15 13 3 2
20 1 10 11 2 10 11 13 16 11 13 9 1 1 10 9 1 10 0 9 2
27 3 2 16 13 13 3 13 10 9 1 10 9 2 10 11 13 4 1 13 10 10 0 9 1 11 0 2
20 10 0 9 1 3 13 1 10 9 15 13 10 11 1 10 11 2 12 2 2
16 3 13 11 2 11 2 12 2 7 11 2 11 2 12 2 2
11 10 9 1 10 9 1 9 2 10 9 2
6 11 2 2 11 2 2
15 15 13 2 3 10 9 1 10 9 1 10 9 1 9 2
5 13 10 9 1 9
9 11 13 9 1 9 1 10 0 9
33 10 11 13 13 10 9 1 9 13 1 13 1 13 10 9 1 10 9 15 1 10 0 9 13 10 9 1 10 9 9 7 9 2
39 15 15 13 13 10 9 2 11 2 15 13 10 9 1 3 1 13 15 1 10 9 1 10 9 1 11 2 10 9 3 13 2 7 3 3 13 9 13 2
12 2 11 2 2 1 3 1 10 11 2 1 11
3 11 13 9
16 2 11 2 13 10 9 13 1 11 15 13 11 1 10 0 2
28 10 9 1 10 2 9 2 1 15 15 13 10 9 1 13 10 9 15 3 13 13 2 7 9 7 13 9 2
5 10 9 3 0 2
21 9 13 9 1 13 10 9 1 10 9 1 9 0 3 15 1 10 11 2 1 11
8 13 9 1 10 9 1 10 11
46 10 11 2 1 10 11 2 13 13 3 10 9 1 10 11 1 3 13 10 10 10 9 1 9 0 1 10 9 1 9 0 15 2 13 12 9 7 0 2 15 13 1 9 1 9 2
33 13 10 9 1 10 9 13 1 10 9 13 1 10 11 2 15 13 10 9 1 10 9 7 13 10 10 9 1 10 9 1 11 2
27 10 9 1 10 11 13 2 3 2 4 1 13 10 9 0 1 10 9 1 10 9 13 1 10 9 0 2
9 3 13 13 10 9 1 10 11 2
40 1 10 9 2 1 9 2 1 10 9 1 10 11 2 1 11 2 3 3 13 13 10 9 1 10 9 1 9 1 10 9 2 13 1 13 1 10 10 9 2
12 9 15 15 13 1 13 10 9 1 10 9 2
19 9 3 2 13 2 3 2 0 2 16 10 9 13 3 1 10 9 13 2
16 13 1 10 9 1 11 2 1 10 11 2 7 13 1 11 2
13 1 10 9 13 0 7 13 15 1 9 1 9 2
7 13 15 1 12 1 9 2
17 1 13 10 9 15 13 10 10 9 1 9 2 10 9 1 15 2
20 13 1 10 9 1 10 9 2 13 1 10 9 1 13 3 3 2 1 13 2
19 1 10 9 2 13 15 13 2 1 10 9 2 1 10 9 1 10 9 2
48 10 9 13 1 4 13 1 10 11 7 10 11 2 11 2 3 13 3 13 2 9 0 1 16 10 9 13 10 10 9 2 7 13 10 9 0 2 3 3 10 9 15 13 0 1 10 9 2
20 7 10 11 2 11 2 13 2 13 10 9 1 10 9 1 10 9 1 9 2
27 10 9 1 10 9 1 10 2 9 2 13 13 7 0 2 15 13 10 0 9 1 10 9 1 10 11 2
21 3 10 9 13 1 10 11 13 1 10 11 2 1 10 11 2 9 1 15 13 2
18 3 16 10 9 13 10 9 1 10 11 1 10 9 1 10 10 9 2
22 13 3 2 13 13 1 10 9 9 2 1 9 0 7 1 9 13 1 10 9 2 2
13 1 10 10 9 2 13 3 12 9 1 10 11 2
11 12 1 15 13 1 15 7 13 15 3 2
17 13 11 2 10 9 1 9 0 1 11 15 15 13 1 10 9 2
10 13 15 10 9 1 9 7 13 15 2
21 2 13 1 11 2 13 1 10 10 9 11 7 13 13 16 15 15 13 13 2 2
12 1 10 9 0 2 10 9 2 13 1 11 2
19 13 15 1 10 11 1 13 15 1 15 15 13 2 7 10 9 13 0 2
18 13 0 9 1 10 9 1 10 9 13 13 15 1 10 9 1 9 2
24 1 10 9 0 2 13 15 10 9 1 10 9 2 13 15 13 10 9 7 13 1 10 9 2
36 13 1 10 9 0 13 15 12 9 1 2 9 2 2 9 0 2 1 1 10 9 2 1 10 10 9 0 2 10 3 0 7 1 9 0 2
30 13 1 10 11 2 13 13 12 9 1 10 9 1 9 2 13 12 9 1 9 1 10 9 1 9 7 1 9 0 2
37 2 9 1 10 9 2 2 9 1 10 9 1 10 9 15 15 13 9 1 10 0 9 0 1 10 9 1 10 9 2 13 10 0 9 1 11 2
18 11 2 13 10 9 1 10 11 2 2 13 10 10 9 7 13 9 2
3 15 13 2
4 1 3 2 2
12 2 13 16 10 9 13 10 9 1 9 2 2
28 10 9 1 10 9 15 13 1 10 9 1 10 11 2 11 2 1 10 9 1 10 11 13 10 9 1 9 2
10 3 2 3 3 13 4 13 1 9 2
35 15 16 11 2 9 7 3 9 1 10 11 2 13 13 10 9 3 13 1 11 16 13 13 10 9 1 9 1 10 9 1 10 9 0 2
14 15 11 3 13 2 13 15 1 13 10 9 1 9 2
28 15 13 3 2 10 9 1 10 9 2 13 1 11 10 9 1 13 10 9 1 10 9 15 13 1 10 11 2
14 10 9 13 13 1 13 7 13 2 3 2 12 9 2
41 3 13 9 1 9 1 10 9 1 10 9 2 10 9 1 13 13 1 12 9 1 10 9 0 13 2 13 9 2 7 13 4 13 10 3 0 9 1 10 9 2
10 11 13 11 3 2 9 1 10 11 2
37 11 2 0 9 1 10 9 0 1 10 11 7 11 2 13 3 1 11 16 2 11 13 9 1 13 1 13 10 9 1 10 11 1 10 11 2 2
19 1 10 9 1 10 9 1 10 9 0 2 10 9 3 3 13 3 0 2
20 3 12 9 1 10 9 13 9 7 3 3 12 9 13 9 0 1 10 0 2
23 12 1 10 9 0 1 10 9 13 13 16 10 9 3 13 1 10 9 1 10 9 0 2
50 1 3 13 13 2 2 3 13 3 1 10 9 0 2 13 9 1 10 9 15 10 9 13 2 2 3 13 10 9 0 1 10 9 2 15 13 3 9 7 9 1 15 3 13 3 13 13 15 2 2
70 11 2 13 1 10 9 1 10 9 2 13 3 3 1 15 13 16 10 2 9 3 13 10 9 0 1 10 9 2 7 2 13 10 9 15 10 9 13 13 1 10 9 0 1 3 13 15 1 10 10 9 2 13 3 16 10 9 7 15 1 10 11 2 1 10 9 13 15 2 2
41 10 9 13 13 3 1 10 9 2 13 13 1 10 9 1 9 1 13 1 10 9 1 10 9 15 13 1 10 9 1 10 11 2 1 12 1 12 1 9 0 2
22 1 3 2 13 13 9 1 10 9 13 10 9 7 13 9 1 10 9 1 9 0 2
46 1 10 9 13 2 13 12 10 9 3 2 15 13 9 15 13 1 10 9 2 10 9 7 10 9 0 1 1 10 9 0 2 9 7 10 9 1 11 1 10 11 7 1 10 9 2
18 15 13 15 1 10 9 1 10 9 0 13 1 10 11 2 11 2 2
32 10 9 13 12 1 10 3 0 9 1 10 9 1 10 9 2 13 13 10 9 1 10 2 9 13 2 1 10 9 0 9 2
7 10 9 13 4 13 9 2
31 3 2 13 11 1 9 2 2 10 9 13 16 13 13 2 9 1 9 1 9 0 2 1 10 0 2 0 7 0 9 2
40 10 9 13 1 10 9 0 1 10 11 13 1 10 11 2 1 15 2 3 2 15 13 10 9 1 10 9 1 10 11 7 15 13 1 10 11 2 11 2 2
41 10 9 13 16 2 10 9 1 9 7 0 9 15 13 1 9 15 13 4 13 1 9 1 13 13 9 0 2 13 1 15 1 10 9 4 13 1 13 13 2 2
15 9 2 13 0 16 10 9 3 13 13 16 13 9 0 2
27 7 13 1 13 16 2 1 10 9 2 13 0 13 10 9 1 13 1 9 7 1 13 9 1 9 0 2
19 7 13 16 10 9 15 10 9 13 2 3 10 9 1 10 11 15 13 2
2 9 0
9 9 2 13 1 13 1 10 11 2
3 2 11 2
2 11 13
40 10 9 11 2 11 2 13 3 10 0 9 1 10 11 2 13 1 11 7 10 11 2 1 10 9 1 12 9 7 13 1 10 0 9 1 10 9 0 0 2
3 11 13 9
27 10 11 2 11 2 13 13 1 9 1 12 3 12 9 1 9 1 9 1 9 13 1 0 7 0 9 2
30 10 9 0 1 10 9 0 1 10 11 13 1 12 9 1 9 2 0 1 10 11 2 1 10 11 7 1 10 11 2
35 10 9 13 13 1 12 7 13 10 9 1 9 0 2 9 1 9 1 9 1 10 11 2 3 10 9 1 9 1 10 9 1 0 9 2
29 3 2 1 1 10 9 1 12 10 11 13 13 12 9 1 10 11 2 1 10 9 0 1 9 13 1 10 9 2
4 9 1 10 11
7 9 2 13 3 7 13 2
30 10 9 2 1 10 9 15 13 2 13 10 9 0 1 10 9 1 9 7 10 2 9 2 3 13 13 1 10 9 2
61 10 9 13 2 1 0 9 2 10 9 0 2 15 13 3 10 9 1 2 9 0 2 7 10 9 1 13 2 9 2 1 10 9 1 10 9 2 13 2 3 2 16 15 13 1 9 1 10 9 1 9 3 0 2 1 9 7 1 9 13 2
17 13 0 16 15 13 1 10 9 3 13 10 9 7 10 10 9 2
26 10 9 0 1 3 15 13 13 10 9 13 1 10 9 1 9 11 2 1 10 13 9 12 1 9 2
44 10 9 13 13 1 12 1 10 3 13 9 1 10 11 2 11 2 9 1 9 1 10 11 1 10 11 0 2 11 2 1 10 11 1 10 11 2 7 11 2 1 10 11 2
26 15 15 13 2 3 2 3 13 16 15 13 13 9 3 1 10 9 15 13 4 4 13 13 3 9 2
30 3 13 10 9 2 10 9 3 13 10 9 1 13 3 13 1 13 15 1 15 15 13 3 13 13 1 10 10 9 2
16 1 15 2 3 3 2 13 1 13 15 1 13 1 10 9 2
9 3 13 13 13 9 1 10 9 2
40 15 15 3 13 13 16 15 13 13 1 13 2 1 0 9 2 16 10 9 3 1 10 9 1 10 9 13 3 3 2 7 1 9 0 2 10 9 1 9 2
24 13 10 11 7 10 0 9 0 2 10 9 1 10 9 13 4 4 3 13 3 15 1 0 2
51 9 15 2 13 3 10 9 3 13 1 13 10 9 1 10 11 1 10 9 1 10 9 0 2 3 13 4 13 1 10 9 2 10 9 0 1 10 9 0 3 13 10 9 1 10 0 9 1 10 9 2
18 3 2 10 9 2 3 13 1 10 9 1 10 9 2 13 10 9 2
33 1 10 0 1 10 9 2 10 9 13 1 13 15 7 10 9 13 13 3 12 9 1 9 1 10 9 1 10 9 1 10 9 2
13 13 2 7 10 15 13 3 13 1 10 9 0 2
17 13 15 1 9 1 9 7 1 9 7 9 2 9 1 9 2 3
10 10 9 3 13 13 3 1 10 9 2
40 13 10 9 1 10 9 1 10 9 1 9 7 9 1 9 0 2 10 9 3 15 13 1 10 9 0 2 3 13 2 3 2 3 1 12 1 9 1 12 2
26 3 2 13 16 15 1 9 1 9 13 3 1 10 0 9 7 16 10 9 1 9 0 13 0 9 2
12 13 13 1 15 2 3 3 13 13 1 11 2
11 10 9 0 13 3 1 10 13 9 0 2
23 12 1 9 2 10 9 13 3 1 10 9 1 16 15 13 1 10 11 1 10 9 12 2
1 9
4 11 13 1 11
56 10 9 0 1 10 11 13 3 10 11 2 15 13 1 11 2 1 15 13 1 10 9 10 11 2 1 12 2 12 1 10 9 2 2 1 10 0 7 0 9 1 10 9 2 1 15 13 3 11 2 11 2 11 7 11 2
29 10 11 13 10 0 9 1 13 1 9 10 12 9 0 15 13 2 3 2 10 9 1 10 9 1 10 9 11 2
53 1 10 0 0 1 10 9 2 15 13 10 9 2 10 9 1 9 1 10 9 0 13 13 15 3 1 10 0 9 1 12 2 13 15 2 1 10 9 2 1 10 9 3 0 15 13 0 9 1 10 9 0 2
24 2 16 15 13 9 1 10 9 2 10 10 9 13 1 10 9 0 2 2 13 10 10 9 2
40 1 3 13 0 16 10 11 13 3 3 10 10 9 2 10 9 1 10 10 9 13 13 3 0 16 1 10 9 13 2 1 10 9 1 10 9 0 2 13 2
43 13 3 9 0 10 11 2 1 10 9 13 3 0 2 10 10 0 1 10 11 13 16 10 11 13 4 1 13 10 2 9 0 2 2 16 3 13 3 10 0 9 0 2
34 10 9 13 13 16 10 11 13 1 13 3 12 2 9 0 2 1 10 11 15 13 10 9 0 1 15 12 1 10 10 0 9 13 2
99 10 9 1 11 7 10 9 0 15 13 10 11 1 11 2 13 1 9 10 2 9 2 0 2 9 1 10 9 2 15 13 1 4 10 11 7 1 4 3 2 13 2 1 10 10 9 0 2 13 2 3 2 10 0 9 15 10 9 0 13 1 13 3 1 10 9 1 10 11 2 11 13 10 0 9 1 10 0 9 0 1 10 11 2 3 1 10 9 1 10 2 9 2 15 13 1 10 9 2
4 2 9 0 2
1 11
5 11 13 15 1 11
75 10 9 1 10 11 13 3 13 10 9 1 10 9 1 10 0 9 0 0 11 1 10 10 9 1 11 2 10 9 1 10 9 0 1 10 11 1 10 9 1 11 2 2 1 15 13 16 10 9 0 13 1 4 13 2 10 9 2 1 10 9 15 15 13 13 3 12 9 7 0 1 10 9 0 2
37 10 11 13 10 9 13 1 10 0 9 2 15 2 13 1 10 9 1 9 2 13 1 10 9 0 15 15 13 13 7 3 13 10 9 1 9 2
47 13 1 10 9 1 10 9 2 1 10 9 13 13 1 10 9 1 3 12 12 9 1 10 9 2 13 13 15 1 10 9 1 10 9 2 1 13 3 1 10 10 9 7 9 1 0 2
55 1 10 9 1 0 9 2 3 10 9 1 10 11 2 10 9 1 9 7 10 9 1 9 1 10 11 2 10 9 1 10 9 2 1 13 11 2 13 13 10 9 3 13 2 2 13 10 9 15 13 0 7 0 2 2
42 3 1 11 2 2 10 9 1 10 9 13 16 10 9 13 1 13 9 1 9 0 2 7 10 0 0 2 3 13 13 1 10 9 1 10 9 1 11 2 11 2 2
33 10 9 1 10 11 13 1 13 13 1 10 11 2 11 2 1 12 2 13 10 9 13 1 10 9 1 10 11 13 10 10 9 2
22 3 13 2 13 2 1 10 9 2 10 0 9 1 10 11 2 1 11 7 11 2 2
29 10 9 1 9 0 2 3 13 2 9 2 2 13 2 3 0 2 1 13 10 9 0 1 10 9 1 10 0 2
39 10 9 3 13 2 1 9 9 2 13 13 3 12 1 10 3 0 9 2 0 1 9 2 2 16 13 10 9 1 10 9 1 10 9 1 10 9 0 2
31 13 15 16 10 9 15 13 3 2 1 10 9 2 10 9 1 10 9 13 1 13 15 1 9 13 1 13 1 10 9 2
20 1 3 16 2 3 10 9 13 0 2 10 9 3 13 13 7 13 10 9 2
20 10 9 13 16 1 9 1 10 9 1 9 13 13 1 9 1 10 9 9 2
55 1 10 0 3 13 2 15 13 1 10 9 0 1 10 9 1 10 9 2 10 9 13 1 13 10 9 1 10 9 9 0 2 3 2 13 1 10 10 9 0 1 9 2 1 10 10 9 2 2 3 2 1 10 9 2
35 1 10 9 13 10 9 1 13 10 9 0 2 13 3 13 13 10 9 1 10 9 0 2 13 1 2 9 1 11 2 1 10 9 9 2
45 10 11 13 2 10 9 2 1 10 9 1 9 0 13 1 10 11 2 16 3 15 13 2 9 0 2 1 10 12 9 1 10 9 11 2 11 2 13 1 12 1 9 1 11 2
34 10 9 13 13 3 1 11 1 10 9 0 1 10 11 2 11 2 3 1 15 13 13 1 10 9 1 10 9 11 7 10 9 11 2
6 10 9 0 1 10 11
43 10 9 0 13 4 1 13 10 9 1 10 11 2 7 1 10 9 3 13 16 1 12 2 7 10 9 13 13 10 9 1 10 2 9 2 2 3 10 9 2 11 2 2
29 10 9 13 13 15 3 1 10 9 1 10 9 0 2 10 9 0 1 10 9 1 12 15 13 3 1 9 0 2
8 13 9 1 10 11 1 10 11
47 10 9 2 13 2 12 9 1 10 9 3 0 1 10 9 11 0 2 10 9 1 10 9 3 0 1 10 11 2 2 15 3 13 10 9 1 10 9 7 15 13 3 1 10 10 9 2
18 1 13 2 13 15 1 10 9 1 10 9 1 10 9 2 10 11 2
24 3 12 9 3 2 12 1 10 9 3 15 13 1 0 9 2 13 10 0 13 13 10 9 2
37 10 9 1 10 9 1 9 15 3 13 4 13 1 10 11 13 1 10 9 1 10 9 2 1 10 9 15 15 13 1 10 10 9 1 10 11 2
23 2 1 10 10 9 2 13 3 13 13 9 13 1 10 9 2 7 3 1 10 9 11 2
16 13 15 1 9 0 15 13 13 0 1 10 9 1 10 11 2
32 3 2 3 13 1 13 1 9 1 10 11 2 1 10 9 1 9 15 13 4 1 13 1 9 0 2 3 13 10 9 0 2
16 7 0 16 13 13 10 9 3 1 13 10 9 0 0 2 2
4 9 1 10 11
29 2 11 2 13 10 9 1 10 9 15 13 13 1 10 0 9 12 7 12 1 9 1 10 11 2 1 10 11 2
44 13 3 1 11 7 11 2 10 9 13 1 10 2 0 9 2 1 10 9 1 11 2 15 13 1 10 9 10 9 1 9 1 10 9 0 13 1 11 1 10 9 1 11 2
38 1 11 2 9 1 10 11 2 9 15 13 10 9 2 10 9 13 3 12 1 10 10 9 0 13 10 0 9 0 1 10 9 1 10 9 7 9 2
27 10 9 2 13 3 1 9 0 1 9 0 2 13 15 3 1 10 9 0 7 13 1 1 10 10 9 2
51 1 10 9 13 13 15 9 1 9 7 9 2 9 0 7 0 2 2 9 1 9 0 2 9 2 9 2 9 2 9 1 10 9 1 11 7 1 11 1 9 7 9 7 10 9 1 9 1 10 11 2
30 13 15 3 10 9 1 10 2 9 2 1 10 11 1 10 9 1 10 9 2 3 1 10 9 0 1 10 9 0 2
19 3 12 9 1 9 13 2 1 10 11 2 13 10 9 1 10 9 13 2
54 10 9 0 13 10 9 1 10 9 0 9 2 15 13 1 10 9 13 9 1 2 9 1 9 2 0 2 1 10 9 13 1 10 9 1 9 13 1 11 2 11 1 10 9 2 2 9 1 10 9 1 9 0 2
11 3 13 13 9 1 10 9 1 10 9 2
36 1 10 11 2 10 9 0 13 1 10 9 1 9 1 9 10 9 1 11 7 11 2 13 3 1 12 9 7 12 9 1 9 1 11 2 2
27 1 10 9 1 10 9 1 10 9 0 1 10 9 0 2 13 13 0 7 0 9 1 9 1 10 9 2
29 10 9 7 10 9 0 13 4 1 13 3 9 13 1 10 9 2 1 3 13 10 9 0 1 10 9 1 11 2
16 10 9 3 13 1 13 11 2 12 9 1 9 1 10 9 2
3 10 9 2
16 15 13 1 13 1 10 9 2 1 10 9 2 1 10 9 2
9 15 3 13 3 13 1 10 9 2
4 10 10 9 2
4 9 13 1 11
33 10 0 9 1 10 9 0 1 9 3 13 9 1 10 9 1 10 9 2 16 10 12 0 13 10 10 9 7 13 10 9 0 2
53 10 11 13 3 10 11 1 12 7 13 3 12 9 2 10 11 13 13 1 10 9 1 10 11 1 12 7 13 1 12 7 10 11 13 1 10 10 9 10 11 1 12 2 13 12 9 2 7 1 15 12 9 2
5 11 13 1 10 11
3 11 1 9
7 11 1 9 13 1 10 11
31 11 2 9 2 13 16 1 10 0 9 10 9 1 10 9 1 10 11 13 13 1 13 1 10 9 15 3 13 1 11 2
38 1 13 0 9 7 10 9 1 10 9 0 1 10 9 0 7 1 13 3 10 9 1 10 9 1 10 9 1 0 9 2 11 3 15 13 1 9 2
46 2 13 13 3 0 1 10 11 3 1 11 2 2 13 3 2 1 10 11 2 10 9 1 10 11 2 1 10 9 15 13 1 9 12 9 1 10 9 1 10 9 1 10 12 9 2
1 9
36 13 15 10 9 2 1 9 2 1 0 7 13 9 1 9 7 9 13 1 10 9 0 1 10 9 0 2 13 1 10 0 1 10 9 0 2
45 10 10 9 0 2 10 9 1 9 1 10 9 7 10 9 1 9 13 9 1 9 0 1 0 9 13 2 7 9 1 10 9 13 0 10 9 1 10 9 3 13 1 10 0 2
9 3 2 10 0 3 13 1 15 2
18 1 13 10 9 11 2 13 9 13 13 3 2 13 9 2 13 3 2
46 10 10 9 11 2 1 0 9 2 13 1 15 13 2 13 15 1 10 9 2 13 10 9 1 15 15 13 1 10 9 2 7 13 10 9 0 13 10 9 2 13 15 1 10 9 2
14 13 2 3 2 10 9 1 10 0 2 0 7 13 2
12 9 3 13 1 10 9 11 2 7 3 13 2
47 2 11 2 13 10 0 1 13 13 7 10 9 1 10 9 1 10 9 3 0 0 1 10 9 13 1 4 13 1 10 9 13 1 2 7 3 1 2 10 9 3 2 3 2 3 0 2
6 2 7 10 9 1 11
16 3 3 15 13 13 2 1 10 9 2 1 10 2 11 2 2
117 16 2 3 1 10 9 1 12 2 13 13 1 9 7 9 2 1 10 9 0 1 11 2 10 9 1 10 9 1 10 9 12 3 0 7 2 3 2 1 12 2 1 11 2 11 13 2 7 13 10 13 9 2 1 15 13 1 1 10 9 1 10 0 10 9 3 0 2 13 10 9 1 10 0 0 3 13 1 10 9 1 10 9 2 1 0 9 1 9 0 7 1 10 0 9 13 9 13 1 9 1 9 3 0 7 0 1 15 13 1 10 9 1 10 9 0 2
9 10 9 0 13 3 1 10 11 2
18 1 10 9 1 10 9 13 10 9 15 13 3 3 12 9 13 9 2
42 1 13 10 10 9 2 10 9 13 3 10 9 1 10 9 1 10 11 7 10 11 2 11 2 1 13 3 10 9 2 15 13 1 10 11 3 12 12 9 1 9 2
55 10 9 0 13 3 1 10 9 1 10 9 1 10 9 2 13 1 9 0 10 9 1 10 11 13 13 1 13 10 9 1 9 1 10 9 1 11 2 7 10 9 1 10 1 13 10 9 15 13 13 1 10 9 0 2
5 10 0 7 10 0
9 10 0 9 3 13 1 10 0 2
15 10 11 2 11 7 10 11 2 11 2 1 10 0 9 2
13 10 11 2 11 7 10 11 2 11 1 10 9 2
5 10 11 2 11 2
31 7 2 15 1 3 3 1 15 2 10 11 2 11 15 2 3 3 2 13 10 9 1 10 9 7 10 9 15 15 13 2
18 10 9 15 13 10 9 7 13 1 10 9 13 13 1 10 0 9 2
20 10 9 3 2 10 13 2 0 7 0 9 0 2 13 9 1 10 9 0 2
18 10 9 0 2 10 9 13 7 0 2 10 9 0 2 0 1 13 2
6 13 15 13 3 3 2
23 3 2 1 10 9 2 11 13 10 0 9 1 12 9 0 1 9 2 13 10 0 9 2
6 15 13 16 15 13 2
5 10 9 1 11 2
5 10 9 1 11 2
5 10 9 1 11 2
20 10 11 13 10 9 13 1 10 9 1 10 12 0 1 10 9 1 10 0 2
16 10 9 0 1 10 9 1 10 9 2 10 9 15 15 13 2
16 10 9 0 2 15 1 10 9 13 13 7 13 1 10 9 2
4 9 12 2 9
28 3 2 3 1 9 1 10 11 2 1 10 11 13 15 10 9 2 13 1 13 15 1 10 11 1 10 11 2
27 1 10 11 2 10 9 13 1 10 11 7 10 11 13 1 13 9 2 13 15 1 10 11 1 10 11 2
43 1 10 2 10 9 1 10 9 2 2 1 11 2 10 9 1 10 9 11 2 10 9 1 11 2 3 9 1 10 2 0 11 2 13 13 2 1 13 2 1 10 9 2
42 11 13 10 0 9 7 10 9 0 13 16 10 10 9 13 2 1 10 9 2 0 2 3 10 9 15 2 13 10 9 2 1 11 13 1 13 10 9 0 2 11 2
32 10 9 1 10 13 1 13 1 9 7 3 2 1 10 0 9 0 2 10 9 1 11 13 10 9 1 9 13 10 10 9 2
25 3 12 12 9 13 3 10 9 1 11 2 10 9 1 10 9 1 9 0 7 10 9 1 9 2
19 13 10 9 2 13 12 9 7 13 13 1 1 10 9 1 10 10 9 2
29 3 2 13 10 9 1 10 9 1 11 1 10 11 7 10 9 3 13 0 9 1 10 15 11 13 1 15 13 2
44 13 15 10 9 1 10 9 1 10 9 1 10 9 2 11 2 11 2 11 2 2 7 10 9 1 10 9 2 11 2 13 3 9 1 10 9 7 10 9 12 1 10 11 2
30 12 1 10 9 0 1 10 9 13 16 11 2 9 2 15 13 1 10 9 1 10 9 10 9 3 0 1 10 9 2
29 3 0 1 15 13 13 1 13 0 9 1 10 9 1 10 10 9 7 1 13 13 1 10 0 9 1 9 0 2
12 1 15 2 13 15 10 9 3 11 13 9 2
65 10 10 9 7 9 1 9 11 13 1 10 9 0 7 2 3 3 2 10 9 1 10 9 2 11 2 0 1 10 2 9 2 1 10 9 1 10 11 2 2 13 1 10 9 2 0 1 3 13 1 10 9 1 10 9 2 13 10 0 11 1 11 7 11 2
1 11
4 9 1 10 11
36 11 13 10 9 1 10 10 9 2 13 1 10 9 9 7 2 1 12 9 1 10 9 2 13 10 2 9 2 0 15 3 13 1 10 9 2
25 13 13 3 12 9 1 10 9 1 10 9 1 10 11 1 9 2 15 13 10 11 1 10 11 2
31 1 10 9 2 10 11 13 1 10 9 3 12 2 1 11 2 12 2 2 7 13 10 9 1 10 0 9 1 10 9 2
40 10 9 13 10 9 1 13 2 13 10 9 1 10 9 1 11 2 3 13 0 7 13 10 9 1 15 13 9 2 1 9 0 1 10 9 1 10 9 2 2
66 1 9 1 10 11 2 11 2 9 1 10 9 1 9 1 10 9 2 10 9 1 9 1 10 9 7 10 11 2 13 13 10 9 2 15 2 1 10 9 2 13 10 9 13 3 1 10 9 1 10 9 2 1 10 9 3 10 15 15 13 1 10 9 1 9 2
33 3 1 3 10 11 13 1 9 10 9 1 10 9 1 10 9 1 9 1 13 1 9 2 3 3 10 9 13 0 1 15 13 2
47 11 2 13 12 9 1 10 9 1 9 0 13 1 10 11 2 13 16 10 9 1 10 11 3 13 9 1 10 9 1 10 9 1 10 9 1 10 9 2 13 10 9 1 11 7 11 2
11 9 2 1 0 2 13 16 15 13 13 2
7 9 2 6 2 3 13 2
19 3 13 13 10 9 1 9 1 10 11 15 13 9 15 3 13 4 13 2
22 16 10 9 13 13 2 15 3 15 13 13 2 10 9 13 13 3 9 2 0 9 2
22 10 9 13 1 10 9 1 10 9 0 2 1 10 9 1 10 9 7 1 10 9 2
28 10 9 13 10 0 9 0 7 3 10 9 1 10 9 7 1 10 9 7 1 10 9 1 10 9 1 9 2
11 10 9 13 16 13 13 1 10 9 0 2
27 10 9 1 10 9 13 13 16 15 2 1 1 10 9 1 12 2 15 13 1 10 12 9 1 10 9 2
11 1 9 2 13 16 15 13 16 13 3 0
4 9 2 3 2
43 1 13 15 10 9 2 13 10 0 9 0 0 1 10 9 1 12 9 7 10 9 0 1 10 11 2 1 10 9 1 9 2 10 9 15 13 10 9 1 10 12 9 2
64 3 2 11 2 15 13 13 10 10 0 9 1 10 9 0 2 7 11 2 1 10 9 13 7 10 9 1 10 11 2 13 15 1 10 9 1 9 0 2 13 3 3 0 9 0 2 15 0 1 10 9 1 10 9 1 10 11 7 10 11 2 1 12 2
44 10 9 3 0 2 15 3 13 3 12 9 1 9 1 9 15 13 13 2 13 4 1 13 9 7 13 10 9 1 10 10 9 13 2 1 10 9 1 9 7 9 3 13 2
38 10 9 1 10 9 1 9 2 3 9 1 9 2 13 9 1 9 2 13 13 10 9 1 10 9 2 13 1 12 12 9 2 1 10 11 1 12 2
55 11 2 11 3 15 13 13 10 10 9 1 11 15 2 1 9 1 10 2 1 9 1 10 9 15 13 1 10 9 1 10 9 1 10 9 1 10 11 2 1 9 1 10 2 0 2 1 10 11 2 13 15 1 11 2
27 10 9 0 13 1 10 9 0 7 2 1 10 9 2 3 13 10 9 2 13 10 10 9 1 0 9 2
8 10 0 0 11 13 1 13 2
44 11 2 10 9 0 13 10 9 1 13 10 2 9 2 1 15 2 12 2 1 10 10 9 2 3 10 9 13 13 13 1 10 9 0 11 2 11 2 16 1 10 9 0 2
26 10 9 13 16 11 15 13 13 2 1 10 9 1 10 9 2 3 12 1 10 0 9 1 10 11 2
32 16 2 1 15 13 2 10 11 13 1 12 9 2 11 13 9 1 9 7 3 13 13 15 1 9 1 13 9 1 10 9 2
21 15 13 10 9 1 10 10 0 9 13 1 10 9 13 9 1 10 10 0 9 2
24 10 9 0 7 0 1 15 10 9 13 1 13 13 9 1 10 9 13 1 10 10 0 9 2
18 15 13 2 13 0 1 10 9 13 1 13 10 9 7 13 1 9 2
28 2 9 3 0 1 10 9 1 10 9 2 16 10 0 13 9 2 7 10 0 9 3 3 15 15 3 13 2
13 10 9 13 13 3 9 1 10 9 1 10 9 2
17 3 16 15 13 3 10 9 0 7 3 0 2 1 9 0 0 2
32 10 9 15 13 1 10 9 13 3 0 13 3 4 13 3 10 0 9 1 10 9 0 2 15 1 15 13 1 13 1 13 2
24 3 13 16 13 9 2 9 7 9 2 13 13 15 13 3 2 10 10 9 1 10 9 2 2
64 1 3 2 3 2 10 0 9 13 1 10 9 1 10 11 7 2 16 13 13 1 10 2 9 1 10 9 3 2 2 10 9 0 3 13 1 13 16 2 16 15 13 2 2 3 13 16 13 12 9 10 16 10 9 15 3 13 0 1 13 10 9 2 2
61 1 10 9 1 10 9 2 11 13 16 3 10 0 9 3 13 10 2 9 1 0 9 7 9 2 1 10 9 0 1 15 1 10 9 2 3 16 10 11 13 1 10 9 1 10 9 2 1 10 9 3 7 1 10 9 1 10 9 0 2 2
22 1 11 2 1 10 11 2 13 0 10 9 2 11 2 2 1 9 1 9 1 11 2
31 10 9 11 13 12 9 1 9 7 10 11 13 10 9 1 10 9 0 2 1 10 11 2 10 9 0 1 10 9 2 2
13 9 1 13 12 9 0 7 12 0 1 9 11 2
39 3 15 13 16 11 7 10 10 9 3 13 1 10 9 1 10 9 16 15 13 1 10 9 1 10 9 2 1 10 2 9 2 7 1 10 9 1 9 2
42 1 10 0 9 2 10 9 13 1 10 9 1 9 2 2 11 2 2 15 13 15 1 13 1 10 9 1 15 15 13 16 1 10 2 9 2 7 10 9 1 11 2
20 11 13 1 9 10 9 7 10 9 2 7 13 10 10 9 3 1 10 9 2
43 1 15 13 9 3 2 11 2 2 2 11 2 7 10 2 11 2 2 13 13 15 3 13 0 16 10 11 7 10 11 13 13 10 9 1 10 9 1 2 0 9 2 2
65 2 11 2 13 2 3 2 10 9 3 0 1 10 9 2 1 10 10 13 9 1 9 15 13 10 11 3 2 1 9 7 9 2 1 13 1 10 9 3 1 10 9 13 7 1 10 9 15 11 13 1 10 9 0 2 2 9 2 2 15 13 1 15 13 2
10 2 13 1 10 11 13 10 9 2 2
37 9 13 3 1 10 9 1 10 9 2 16 10 0 2 9 2 1 11 1 10 9 13 1 10 11 2 3 13 10 9 1 10 9 1 10 11 2
20 10 9 13 15 2 11 2 7 2 16 15 2 0 2 2 13 1 10 15 2
24 9 3 1 10 0 9 1 11 2 15 3 13 1 11 1 15 13 1 10 0 1 10 11 2
27 10 9 13 1 10 0 9 2 1 9 1 10 0 2 7 13 3 0 1 10 9 2 12 9 1 11 2
34 3 2 10 9 13 3 12 9 1 10 0 9 1 10 11 2 1 9 1 11 7 9 1 11 2 1 10 9 0 2 1 12 9 2
25 9 1 10 9 1 10 11 2 1 12 9 1 9 2 15 13 12 1 10 9 0 1 10 11 2
4 9 13 9 0
8 9 0 1 10 9 1 10 11
17 1 10 11 2 10 12 9 1 9 0 0 1 10 9 13 0 2
17 1 10 11 13 3 3 9 10 9 0 1 10 11 2 1 11 2
8 9 2 2 9 2 1 10 11
3 9 1 9
42 12 9 0 13 3 13 13 15 10 9 1 10 11 1 10 2 9 2 1 10 11 1 9 2 15 1 3 7 3 13 1 10 9 1 11 2 1 10 11 1 11 2
26 3 1 13 13 10 9 0 3 1 10 9 1 10 12 9 13 2 10 9 3 13 13 3 3 3 2
41 1 9 3 10 9 1 10 11 2 10 9 1 10 11 7 10 9 1 10 11 2 0 9 1 10 9 2 2 1 10 11 3 3 13 16 13 13 10 9 0 2
28 10 9 1 10 11 13 10 9 0 1 13 10 9 3 15 13 10 9 15 13 3 10 9 1 9 7 9 2
44 13 2 3 3 2 1 15 13 1 9 7 13 1 9 1 10 9 1 9 7 10 0 9 7 9 1 9 0 2 7 3 1 10 0 9 1 9 15 1 15 13 13 0 2
30 10 9 1 10 11 7 1 10 11 2 1 10 10 0 9 2 13 1 9 10 9 1 10 9 1 15 2 9 2 2
22 13 9 1 13 10 9 7 1 15 13 1 10 9 0 7 0 2 3 13 10 9 2
51 3 16 2 13 11 2 2 2 10 9 13 10 9 1 10 9 3 3 13 2 16 15 13 13 3 3 13 1 15 16 3 10 3 0 1 1 10 9 13 3 13 13 3 9 16 15 15 3 13 2 2
4 1 13 4 2
2 2 9
49 1 12 2 13 12 9 1 15 10 9 2 13 1 0 9 7 9 0 15 13 1 10 9 1 15 13 1 9 0 15 13 1 10 9 1 9 2 3 10 11 1 11 2 13 2 11 2 2 2
35 1 10 9 2 10 9 1 10 9 2 13 3 0 2 2 16 2 3 15 13 13 0 9 2 15 13 1 15 13 1 10 9 1 9 2
40 10 12 0 9 1 10 9 13 10 13 2 9 1 9 0 2 2 3 10 11 2 7 15 1 9 0 2 1 15 15 3 13 13 10 11 2 1 10 11 2
73 1 10 9 0 2 1 15 10 9 13 10 10 9 2 7 3 2 1 10 9 1 11 2 3 13 13 9 0 2 2 10 9 1 9 0 2 13 1 10 9 12 7 13 1 10 9 1 10 9 1 12 2 13 10 9 13 1 10 9 2 13 1 10 2 9 2 1 10 9 1 10 9 2
28 13 2 3 2 1 11 2 15 13 12 9 1 10 9 1 10 9 2 13 10 9 1 10 11 1 10 11 2
25 10 0 1 11 2 12 9 13 1 9 2 13 1 10 11 3 12 12 9 7 13 1 13 9 2
12 1 11 1 10 11 2 11 13 3 10 9 2
29 1 11 7 10 10 9 1 9 2 11 3 13 10 0 9 7 2 3 2 13 3 1 13 10 9 1 13 9 2
20 10 9 0 13 3 10 9 2 13 1 10 9 1 10 9 7 13 10 9 2
36 11 13 12 9 1 10 11 1 10 9 13 2 3 3 1 12 0 9 1 10 9 2 1 11 2 3 0 2 1 10 9 15 13 3 11 2
24 13 10 9 0 2 15 15 13 1 10 9 1 10 9 7 10 9 3 0 1 10 0 0 2
20 13 3 7 10 11 13 1 13 10 11 1 12 9 1 11 7 12 1 11 2
7 13 3 1 10 9 0 2
22 10 9 13 16 3 13 10 10 2 9 1 9 2 3 10 9 13 1 13 10 11 2
27 3 16 2 3 2 13 1 10 9 16 13 10 11 2 13 3 16 3 11 13 13 10 10 9 3 0 2
31 13 0 16 10 9 13 13 2 7 3 13 2 10 9 1 9 1 13 10 9 1 13 16 10 11 13 10 9 1 11 2
21 2 1 10 9 13 3 0 13 12 9 1 10 9 2 2 13 10 9 0 11 2
51 1 9 0 1 10 9 2 7 2 1 10 9 1 13 10 9 0 2 2 10 9 1 10 11 2 13 13 1 9 10 9 1 9 2 2 13 2 10 9 15 10 9 3 13 1 13 2 1 10 9 2
27 1 10 9 1 10 9 1 10 9 2 1 13 1 10 11 10 0 1 10 11 2 2 13 3 0 2 2
76 11 2 9 1 10 11 2 13 15 1 13 2 1 10 9 2 16 2 2 1 12 9 1 0 9 1 10 0 9 2 2 13 1 9 1 12 2 2 10 9 13 10 9 13 2 7 16 2 10 9 13 2 1 10 11 2 1 10 10 9 2 2 10 0 9 7 9 1 10 9 13 2 1 10 9 2
5 7 3 3 13 2
11 7 10 9 1 10 9 3 13 3 0 2
15 10 9 9 13 2 3 2 10 0 9 2 13 0 9 2
28 1 15 1 10 9 1 10 9 13 1 9 1 10 9 1 9 1 9 2 10 9 13 3 0 2 1 9 2
20 3 15 13 2 3 2 16 1 1 10 9 1 10 9 15 13 9 1 9 2
33 10 9 11 13 1 9 2 13 15 1 10 12 9 2 3 12 9 2 3 10 11 13 12 9 1 15 13 15 1 10 12 9 2
17 1 9 2 1 10 11 13 15 12 9 1 9 2 3 12 9 2
17 10 11 13 1 12 9 1 9 2 3 12 9 16 1 10 9 2
18 3 3 1 13 2 10 11 3 13 1 13 1 10 9 1 10 11 2
49 10 0 1 10 9 0 13 1 13 11 7 2 3 2 1 10 9 13 1 10 9 1 15 13 13 1 10 9 1 9 0 0 2 7 3 13 10 9 3 1 10 11 1 10 9 1 0 9 2
17 10 0 9 1 10 9 1 3 13 11 2 11 2 11 7 11 2
34 10 9 1 10 0 9 1 10 9 1 9 1 10 9 1 0 9 0 13 2 3 2 15 10 11 13 1 10 9 1 10 9 0 2
48 13 1 10 9 0 1 12 2 10 9 0 13 1 10 9 0 1 10 9 1 10 11 13 3 1 10 0 9 7 13 13 1 10 0 11 2 2 10 9 0 13 3 13 1 10 9 0 2
37 7 10 9 1 10 11 13 9 1 10 9 2 1 10 9 1 10 2 9 2 3 13 2 9 2 1 13 10 0 9 1 9 1 13 10 9 2
56 16 13 13 10 9 0 1 10 9 3 1 9 0 2 15 3 13 13 3 2 2 10 0 15 15 13 13 4 1 13 10 9 13 1 10 2 9 0 1 12 9 1 10 9 1 10 9 1 10 9 0 2 2 11 2 2
54 3 1 10 9 13 1 10 9 12 1 10 9 12 2 10 9 13 13 3 10 2 9 7 9 0 13 1 10 9 2 2 1 13 1 10 9 1 9 2 15 13 16 13 10 9 2 1 9 0 7 1 9 2 2
9 10 9 1 12 9 3 13 0 2
34 15 13 3 1 10 9 0 1 10 9 1 10 11 2 15 10 9 13 1 10 11 2 3 1 10 9 15 13 4 13 1 10 11 2
7 10 9 3 3 13 0 2
18 13 15 10 9 1 11 7 11 2 9 1 9 1 11 0 1 11 2
41 1 10 9 2 1 10 10 9 13 15 1 10 9 1 10 9 13 2 1 10 9 1 9 2 10 10 9 15 13 13 10 9 2 12 1 11 2 12 1 11 2
10 2 9 1 10 9 1 13 13 2 2
31 9 2 0 9 1 10 9 1 10 9 13 15 1 10 9 7 1 10 9 1 10 9 1 10 9 15 10 9 15 13 2
5 13 15 10 9 2
19 1 15 13 15 3 10 9 7 13 15 13 3 2 7 1 10 10 9 2
20 10 9 1 10 11 13 10 9 1 10 9 2 13 3 1 10 9 1 9 2
15 10 10 9 1 10 9 13 3 13 1 10 9 1 9 2
53 10 9 13 13 15 1 10 9 1 15 13 10 9 7 13 2 3 10 9 1 10 11 15 2 1 12 7 12 2 13 13 10 9 1 9 1 12 9 2 1 10 9 1 12 9 1 10 11 2 11 7 11 2
74 1 13 10 9 2 15 3 1 10 12 9 1 10 11 2 11 2 13 12 9 1 9 2 2 10 11 13 10 9 1 10 9 1 10 9 1 9 2 10 9 13 13 1 10 9 1 9 0 2 7 2 1 10 9 2 13 0 2 13 10 9 1 10 9 7 1 10 9 1 2 9 2 2 2
44 13 10 11 16 2 13 10 9 0 1 3 10 9 1 13 10 9 7 10 9 0 1 10 9 1 9 0 2 1 10 9 1 13 10 9 15 13 10 9 1 0 9 2 2
52 1 10 9 13 15 10 13 9 0 1 10 9 2 10 2 9 2 1 10 9 1 9 2 10 2 3 13 2 9 7 10 9 1 9 1 9 2 13 2 3 0 2 2 3 9 0 1 10 9 1 9 2
32 3 2 10 11 13 13 3 1 11 2 1 15 15 13 13 1 10 9 7 13 10 9 1 10 11 1 16 13 13 10 9 2
68 2 10 9 9 13 15 16 15 15 15 13 1 13 13 0 7 16 10 9 13 9 1 13 13 2 7 13 15 16 13 13 1 16 15 13 1 10 9 0 2 2 13 15 11 2 10 9 1 13 10 9 1 10 9 1 1 10 9 0 1 10 9 3 13 10 9 0 2
46 10 9 2 3 2 1 10 9 1 10 15 13 1 10 11 10 9 2 11 2 2 13 1 10 11 16 2 10 9 0 3 13 13 10 9 1 10 9 1 10 9 2 11 2 2 2
5 9 1 11 13 11
37 10 11 1 10 11 13 3 11 7 13 10 11 2 15 13 10 9 1 10 9 11 2 11 3 1 13 13 10 9 1 13 11 1 9 1 9 2
47 10 9 0 13 2 0 2 10 9 1 11 2 7 13 16 3 13 13 1 10 9 10 9 1 10 9 15 15 13 13 2 1 15 10 9 1 10 11 3 13 4 15 13 1 10 9 2
41 1 15 2 13 10 2 9 1 9 2 1 10 9 7 13 10 10 9 1 10 9 1 11 2 1 13 10 9 1 2 10 9 0 15 3 15 13 3 13 2 2
21 3 13 1 13 16 11 15 13 1 10 9 2 3 1 10 0 9 1 2 11 2
43 10 9 0 1 9 1 9 13 12 9 1 9 2 3 10 9 1 10 9 13 12 12 9 1 9 0 2 12 9 13 1 9 1 9 7 3 12 9 1 9 0 2 2
41 3 2 1 9 1 10 9 11 13 1 10 9 2 11 2 2 13 13 12 9 1 9 1 2 11 2 1 15 10 9 2 13 12 9 1 9 15 3 15 13 2
24 10 11 13 16 2 1 10 9 2 3 13 0 13 10 12 9 1 9 13 1 10 13 9 2
39 1 10 9 1 10 9 2 11 2 2 15 15 15 13 1 10 9 1 10 9 13 10 9 7 10 9 1 16 10 11 13 1 13 9 1 10 9 2 2
11 3 3 2 1 10 11 13 2 11 2 2
36 7 10 9 1 10 9 3 0 1 10 9 13 1 10 0 9 1 10 9 13 1 13 1 10 0 9 1 15 10 9 13 13 1 10 9 2
24 1 10 9 2 10 9 1 10 9 13 1 13 12 9 15 3 13 13 2 9 7 0 9 2
36 10 9 13 1 10 9 1 10 9 13 3 13 10 9 1 10 9 1 13 15 3 1 10 9 1 10 9 1 13 1 10 9 1 10 9 2
23 13 3 16 10 9 2 11 2 13 1 10 0 9 1 9 1 10 9 3 13 1 11 2
69 10 0 9 15 13 1 10 9 0 13 10 9 15 13 13 10 9 0 2 11 13 9 0 2 1 13 10 9 2 11 2 1 13 10 9 2 3 2 16 2 1 15 2 13 10 9 1 9 2 10 9 0 13 10 0 9 1 15 15 13 13 10 9 1 9 2 2 13 2
19 2 11 13 3 2 13 11 1 13 1 4 2 13 1 10 9 0 2 2
59 1 10 9 0 13 1 10 11 2 10 0 9 1 10 9 0 1 13 10 9 1 10 9 13 1 10 9 0 2 2 11 13 13 15 1 10 9 2 15 15 13 13 10 9 2 7 13 13 1 10 9 11 2 15 13 3 1 11 2
3 9 7 9
21 10 11 13 1 10 9 13 10 0 9 1 9 1 10 9 1 10 11 1 12 2
29 1 10 9 0 13 13 3 10 9 1 12 9 2 0 1 12 9 1 10 9 13 3 2 1 10 11 1 12 2
28 7 3 10 9 0 13 13 1 9 2 10 9 1 11 13 10 9 0 2 1 10 0 12 9 1 12 9 2
29 10 9 0 1 11 13 13 9 7 13 10 9 3 10 9 13 13 1 15 2 7 3 13 16 15 13 13 2 2
20 9 1 9 2 10 9 1 9 0 13 13 10 9 0 1 10 9 15 13 2
15 16 3 15 13 9 1 15 2 13 15 15 3 13 13 2
17 1 10 9 0 1 9 1 10 11 2 1 11 2 13 12 9 2
24 1 15 13 2 9 13 10 2 9 2 7 2 15 2 13 1 10 9 2 10 2 9 2 2
10 11 1 10 9 1 10 11 1 10 11
50 11 2 11 2 11 2 11 7 11 2 10 0 15 3 13 9 1 10 11 2 13 10 9 13 7 3 13 1 10 11 1 13 10 9 1 10 11 1 10 9 7 9 0 1 10 9 1 10 9 2
26 10 11 13 3 13 13 1 10 9 1 11 2 11 2 11 7 11 2 11 2 11 2 11 7 11 2
25 3 1 10 9 1 11 7 1 10 9 2 10 11 13 3 13 10 9 1 10 9 1 10 9 2
18 3 10 0 9 3 13 13 10 9 0 1 9 1 9 1 10 11 2
31 1 10 2 9 2 1 10 9 13 15 3 15 13 13 1 10 9 1 9 0 7 0 1 9 2 9 2 9 7 9 2
22 10 9 13 1 13 10 9 7 13 3 1 12 7 12 9 2 12 1 12 9 2 2
38 10 9 1 10 9 1 10 9 2 13 1 9 7 1 10 11 2 13 1 12 7 12 9 2 12 1 12 2 2 9 1 15 10 9 13 12 9 2
17 10 0 9 13 13 1 10 9 0 1 10 9 7 13 1 9 2
35 15 1 10 9 13 15 3 1 10 9 0 1 12 9 1 9 7 1 10 9 15 13 13 1 1 10 12 12 9 2 12 12 9 2 2
35 7 11 2 9 1 11 2 9 7 9 1 12 1 10 9 2 10 11 2 2 3 13 10 9 1 16 10 11 0 13 9 1 10 9 2
22 11 13 3 16 10 9 3 13 13 1 10 9 1 10 10 9 15 13 1 10 11 2
23 1 10 9 10 11 13 9 1 10 9 0 1 15 1 10 9 0 2 13 13 10 9 2
16 1 15 15 13 1 10 11 0 2 13 15 12 9 1 11 2
23 1 10 0 2 1 12 9 2 13 13 12 9 1 9 2 1 10 9 0 1 12 9 2
23 1 10 0 2 1 12 9 2 13 13 12 9 1 9 2 1 10 9 0 1 12 9 2
41 7 1 10 0 2 1 12 9 2 13 13 12 9 1 9 2 1 10 9 0 1 12 9 2 15 13 1 13 10 9 1 10 9 1 10 9 0 1 0 9 2
10 2 15 13 0 1 15 3 13 2 2
24 11 2 1 10 9 1 10 11 2 1 10 9 1 10 9 1 10 11 2 2 11 2 2 12
32 2 10 11 13 2 3 1 10 9 1 9 2 13 10 9 1 10 10 9 2 7 1 10 0 9 2 13 9 7 9 2 2
7 10 9 13 3 10 9 2
14 3 13 13 15 2 3 13 13 1 15 13 1 15 2
17 13 15 2 1 3 7 3 2 15 15 13 7 15 15 13 3 2
34 10 9 1 13 1 9 13 13 1 10 9 1 10 11 7 1 10 10 9 1 10 9 2 15 13 10 0 9 1 10 9 0 0 2
38 2 3 10 9 3 13 3 2 13 0 13 10 9 2 2 13 12 1 10 9 1 10 9 1 9 0 15 13 1 10 9 1 10 9 1 10 11 2
28 10 9 1 12 9 13 1 13 10 9 0 0 1 10 9 0 13 15 1 10 9 13 1 10 9 1 11 2
40 2 13 13 1 9 0 9 10 9 0 1 10 9 2 1 10 9 3 15 13 2 16 3 3 13 9 0 1 10 9 2 2 13 11 2 15 13 3 9 2
37 10 9 1 10 9 2 15 13 13 1 10 9 1 10 11 2 13 1 9 1 10 9 1 13 1 10 11 0 1 10 9 1 10 9 7 9 2
32 3 1 10 0 9 12 2 10 9 0 13 13 15 1 10 9 11 1 13 2 3 2 10 9 1 10 9 1 10 9 0 2
10 3 2 10 9 13 15 1 10 9 2
43 3 3 1 15 15 15 13 3 1 10 9 3 0 1 10 11 2 7 3 1 10 9 15 10 9 1 11 13 1 13 7 2 3 2 1 15 15 10 9 13 1 13 2
32 1 10 9 13 3 1 10 11 2 10 11 13 1 11 12 1 10 12 9 1 15 13 2 13 10 11 3 1 10 9 0 2
19 1 12 1 9 2 13 15 16 13 3 1 10 2 9 2 0 1 11 2
14 3 13 0 3 2 7 10 9 3 13 3 13 9 2
27 10 9 1 10 11 2 10 0 15 13 1 15 12 15 3 13 2 13 3 13 7 13 13 1 10 9 2
30 10 9 13 1 10 9 1 10 0 9 11 2 11 13 1 13 10 9 1 3 7 13 2 3 2 13 10 10 9 2
33 10 9 0 1 10 9 2 9 1 10 9 0 2 13 13 1 10 9 1 10 0 9 2 9 15 13 1 10 9 11 7 11 2
14 1 10 10 9 2 13 10 9 13 1 9 1 9 2
27 10 9 1 10 9 0 13 13 1 10 9 1 10 9 2 13 1 9 2 13 0 9 1 10 9 13 2
32 3 1 11 2 10 0 9 2 1 10 9 2 10 9 0 13 1 13 9 1 10 9 3 10 9 15 13 1 13 10 9 2
32 13 15 13 2 3 1 10 9 15 13 3 1 10 9 13 13 2 13 10 9 8 1 10 9 1 2 3 2 13 10 9 2
19 1 12 2 10 9 13 13 7 2 12 9 3 2 15 13 1 10 15 2
20 3 2 10 9 0 1 10 0 9 0 13 3 1 13 10 9 1 10 11 2
35 10 9 2 7 3 10 11 2 13 13 16 10 9 0 13 3 1 10 9 10 10 9 0 16 10 9 0 2 1 10 9 2 10 9 2
50 16 10 11 13 13 10 12 9 2 13 3 1 10 9 1 11 13 10 9 1 10 9 0 2 13 3 16 10 9 2 9 2 2 13 1 10 11 2 13 13 1 10 11 2 15 13 2 9 2 2
25 9 2 3 10 9 1 10 9 13 1 10 9 2 13 1 13 1 10 9 7 13 1 10 9 2
18 13 15 10 9 1 13 1 10 9 7 13 15 2 1 9 1 9 2
13 9 2 15 10 10 9 1 10 9 1 10 9 2
27 9 2 10 11 13 15 1 10 9 2 3 9 2 7 3 13 9 1 10 10 9 7 1 10 10 9 2
27 3 2 1 10 9 2 10 11 13 10 11 2 13 3 10 11 15 2 3 2 13 13 10 11 1 13 2
6 9 2 1 10 9 2
1 11
7 3 13 10 9 1 10 9
36 2 10 9 1 13 10 9 2 7 1 13 10 10 9 2 7 1 13 15 2 13 4 13 7 13 3 9 1 10 9 0 1 10 9 2 2
35 15 13 12 1 10 9 0 1 10 9 1 10 11 1 10 9 2 15 13 13 13 10 9 2 0 2 1 13 10 9 1 10 9 0 2
36 3 10 9 3 13 13 15 3 16 11 7 11 13 1 10 9 1 10 9 2 16 1 10 9 10 9 1 11 13 3 13 1 10 9 12 2
47 15 16 2 3 1 10 9 2 1 10 0 13 13 10 9 15 13 15 1 9 1 10 9 13 2 3 2 3 12 9 3 12 2 2 13 15 1 10 9 10 9 1 9 7 10 0 2
5 3 3 13 3 2
62 10 9 1 10 9 1 10 9 1 9 1 10 9 0 3 13 13 1 10 9 1 10 9 0 2 1 12 1 9 1 12 2 15 13 13 9 1 10 9 15 13 1 10 9 10 11 2 11 2 7 10 11 2 11 2 1 10 11 2 11 2 2
8 3 10 9 1 9 1 10 9
3 9 13 11
13 13 1 9 0 2 10 11 7 10 11 13 3 2
31 10 9 13 1 10 9 1 10 9 13 1 13 9 0 7 3 13 10 9 15 13 1 11 1 13 10 9 1 10 9 2
1 11
12 12 11 2 10 9 1 10 11 13 1 11 2
7 12 11 2 10 9 1 11
37 0 9 1 10 9 0 0 2 1 15 12 9 1 9 15 13 1 13 2 13 2 13 9 7 1 13 9 0 2 10 11 13 10 9 13 9 2
15 7 1 15 13 3 0 1 2 9 2 2 9 0 2 2
45 13 12 9 2 9 1 10 9 7 9 1 9 0 13 3 12 0 7 13 10 9 2 3 10 9 0 13 2 11 2 13 2 1 9 2 10 13 9 1 10 9 1 9 0 2
34 13 15 15 15 13 3 2 1 10 9 2 13 3 1 9 3 13 1 10 9 2 1 10 15 10 9 13 4 13 1 9 3 0 2
25 13 2 13 15 1 10 11 2 3 15 13 11 2 1 11 1 13 16 13 3 0 1 10 9 2
32 13 2 1 10 9 15 15 10 13 2 10 9 1 9 2 0 1 15 1 10 9 1 10 11 2 3 3 0 1 10 9 2
24 7 2 3 13 10 9 1 9 1 10 9 2 3 13 1 13 7 1 13 3 1 10 11 2
31 9 7 9 2 10 11 3 13 9 1 10 9 7 1 10 9 2 10 0 9 13 1 16 2 1 9 2 13 15 9 2
35 13 7 13 7 10 9 1 9 13 15 1 0 9 2 10 10 9 2 10 10 9 2 10 10 9 2 10 10 9 13 15 1 10 15 2
12 3 13 3 13 2 3 3 3 13 15 13 2
25 11 13 10 0 1 13 3 10 9 2 1 10 0 9 2 1 10 10 9 0 1 11 2 11 2
22 1 10 9 2 11 13 10 10 9 13 9 7 13 3 2 1 10 9 2 13 9 2
16 10 9 1 10 11 11 13 10 0 1 13 15 2 9 3 2
29 3 13 1 10 11 7 1 11 2 11 13 13 10 9 1 10 10 9 1 15 13 1 10 10 9 10 9 3 2
7 10 9 13 1 13 10 9
48 10 9 0 1 10 11 2 11 2 2 13 1 10 0 9 1 10 9 0 2 11 2 2 13 16 10 9 13 3 1 13 7 16 10 9 1 9 0 13 12 1 10 9 0 1 10 9 2
20 10 9 1 10 11 13 4 13 1 10 9 0 15 13 9 1 11 1 9 2
44 10 11 13 1 10 9 10 9 1 12 9 15 13 1 10 9 10 0 9 1 9 0 2 10 9 1 9 7 9 2 10 9 1 9 7 10 9 1 9 1 10 9 0 2
33 10 0 9 1 10 11 2 13 1 12 2 13 16 10 9 1 10 9 13 1 13 7 3 13 13 16 10 9 13 10 9 0 2
10 3 2 13 10 9 2 3 13 9 2
20 10 11 13 10 9 1 9 15 13 13 1 12 1 10 11 7 1 10 11 2
34 7 10 11 13 4 1 13 10 9 0 1 10 0 9 2 15 15 13 9 1 9 2 1 10 9 1 3 12 9 1 10 10 9 2
25 10 9 0 13 15 1 10 9 1 9 2 16 13 13 1 13 10 9 1 9 1 10 0 9 2
10 3 2 10 11 13 10 9 15 13 2
26 13 10 9 1 10 9 13 1 10 11 7 1 11 2 11 7 11 2 3 10 9 13 1 10 9 2
16 10 9 1 10 11 1 10 11 13 10 9 1 9 1 9 2
23 10 9 0 13 1 10 9 1 3 12 9 1 10 11 2 3 1 10 11 2 1 11 2
2 9 3
26 13 10 9 0 2 10 9 13 3 9 1 9 1 10 9 1 10 9 13 9 2 13 9 7 9 2
13 3 1 15 15 13 1 10 2 9 1 9 2 2
29 1 10 9 2 10 11 13 1 12 9 1 10 9 2 13 3 10 9 1 10 9 1 10 9 3 13 13 0 2
13 2 15 13 1 13 9 7 15 13 13 1 13 2
21 7 2 13 2 13 16 10 9 3 13 1 4 13 1 10 9 0 1 10 9 2
23 13 1 4 13 1 10 0 16 15 13 12 7 12 9 3 16 10 9 1 10 9 2 2
16 1 11 2 10 9 0 1 11 13 3 10 0 1 12 9 2
15 2 3 2 16 13 13 10 9 1 10 9 1 10 11 2
75 3 16 13 9 1 10 9 1 9 0 2 11 7 11 2 15 2 1 15 13 10 9 1 10 9 2 13 1 16 15 3 13 13 10 0 2 7 2 0 2 16 10 9 1 10 9 13 10 9 1 10 9 1 10 9 1 9 0 2 15 13 10 9 0 1 10 9 1 10 0 1 0 9 2 2
2 9 13
15 10 9 9 1 10 11 13 1 13 9 1 10 9 0 2
33 9 13 16 10 9 13 13 10 10 9 1 10 0 9 1 10 0 9 1 10 9 0 7 0 2 3 13 13 1 10 0 9 2
7 10 9 11 13 12 9 2
39 10 9 0 1 11 7 11 13 3 13 10 9 1 10 9 1 10 9 2 15 15 13 2 13 2 1 10 9 1 10 9 7 1 10 9 1 10 9 2
88 3 2 16 1 10 2 9 2 1 10 2 9 2 10 9 1 10 11 13 13 2 3 2 10 9 1 11 2 3 10 0 9 0 0 1 10 9 2 11 2 3 13 0 9 2 13 1 0 9 1 10 11 1 10 11 2 2 13 0 12 9 2 10 10 16 11 2 1 12 9 1 10 11 2 15 3 13 10 0 0 9 1 10 11 1 10 9 2
41 10 9 1 10 11 13 0 16 13 1 10 9 1 16 10 0 13 1 0 2 1 10 9 15 13 13 15 1 10 9 1 9 0 15 13 1 13 10 0 2 2
15 10 9 1 9 1 10 9 13 10 9 2 1 0 9 2
42 1 10 11 2 10 9 2 1 9 0 1 9 2 1 10 11 2 1 10 9 1 15 10 9 11 13 10 9 0 2 3 13 3 16 10 0 12 9 1 10 9 2
23 3 2 10 13 7 13 2 9 0 0 3 0 2 2 10 11 2 13 16 3 15 13 2
53 10 11 2 15 13 10 9 0 1 10 9 1 10 9 1 9 2 7 10 9 3 3 0 1 10 9 0 1 10 9 2 3 13 3 16 10 9 1 12 9 1 9 0 1 10 9 13 1 10 9 3 13 2
7 10 9 1 15 2 13 2
42 15 13 13 2 3 16 13 1 13 2 13 10 9 0 1 10 12 9 1 10 11 2 15 13 13 15 1 10 11 1 10 11 1 12 2 3 3 3 10 9 2 2
32 3 1 2 1 10 9 2 13 10 9 2 13 1 10 9 1 11 7 11 2 15 3 13 10 10 9 1 10 9 1 11 2
28 10 0 9 2 10 11 13 13 1 10 11 2 1 10 9 3 7 0 1 10 12 9 1 11 1 10 11 2
15 15 2 1 10 9 15 13 2 3 3 13 9 7 9 2
149 1 10 9 0 1 15 13 13 13 10 9 7 10 9 3 0 1 10 10 9 0 7 0 2 10 9 11 2 3 13 1 10 9 0 2 7 3 3 13 1 11 7 1 10 11 2 13 15 2 1 10 2 1 10 9 1 10 9 0 2 1 10 12 9 2 1 13 10 9 15 2 1 10 9 2 13 1 10 9 1 10 11 7 1 10 0 9 1 15 13 1 1 10 0 9 1 10 9 1 10 9 7 1 10 9 0 1 10 10 9 2 9 1 10 9 0 1 10 9 1 9 1 10 9 7 1 10 9 15 12 9 13 1 13 1 9 0 2 13 1 10 9 0 15 13 1 10 0 2
188 10 12 9 2 11 7 10 11 2 13 15 7 13 15 1 10 9 0 2 1 10 9 2 1 10 9 1 10 9 0 2 1 10 9 0 1 10 9 0 2 1 2 11 2 7 10 9 1 9 0 7 0 2 1 1 10 2 11 2 1 11 2 1 10 2 11 2 1 11 2 1 10 2 11 2 1 11 7 1 10 2 11 2 1 11 2 13 1 10 9 1 10 9 15 13 10 2 11 2 1 11 2 15 1 10 0 2 1 10 9 0 1 10 9 0 2 10 0 9 1 11 2 11 2 2 2 3 11 13 3 9 1 10 11 2 0 2 2 3 13 7 1 10 9 2 2 1 10 9 0 7 1 10 9 11 2 13 1 10 9 1 10 9 15 15 13 1 10 9 0 2 1 13 10 0 9 1 9 2 1 11 15 13 10 9 1 15 2
8 9 1 9 13 9 1 12 9
4 13 1 10 9
26 10 11 1 11 13 10 9 0 1 10 9 1 10 9 1 9 2 1 15 13 13 9 9 1 9 2
49 1 15 15 15 13 2 10 9 1 9 1 10 9 13 1 10 9 1 9 2 1 10 2 11 2 7 1 10 9 2 11 2 2 1 9 0 2 13 1 9 0 1 10 9 2 3 1 11 2
25 3 2 11 13 16 13 10 2 9 1 11 2 1 10 0 9 1 9 1 10 9 1 10 9 2
25 2 13 10 9 15 3 13 1 12 9 7 13 10 9 1 15 13 2 13 16 13 15 3 13 2
22 10 9 13 16 10 9 13 3 15 15 13 7 13 10 9 1 13 13 10 9 2 2
58 1 10 9 1 12 9 10 9 11 2 1 10 11 2 13 10 10 0 9 1 10 2 11 2 2 3 13 1 10 11 2 2 13 1 3 12 9 10 9 11 2 11 2 7 10 9 11 2 11 2 2 3 2 0 7 0 13 2
29 10 9 13 3 13 1 11 2 9 1 10 9 1 10 11 2 15 13 10 9 1 10 9 7 3 3 15 13 2
6 10 9 3 13 10 9
28 1 10 11 2 10 9 0 13 0 3 1 10 9 2 15 15 13 13 10 9 1 10 9 1 10 9 11 2
25 10 11 13 15 3 13 2 7 15 13 1 10 9 7 2 1 15 10 2 3 13 1 10 9 2
23 3 3 1 10 9 1 10 9 1 11 2 13 10 11 2 3 1 10 0 11 1 11 2
6 3 1 9 2 11 2
12 7 1 10 11 13 0 13 10 9 1 9 2
22 10 9 1 12 1 9 13 4 13 2 3 2 3 10 9 1 10 9 1 10 9 2
45 1 10 9 1 10 9 2 3 2 10 9 0 13 10 9 1 10 9 13 1 9 1 9 2 15 2 1 13 15 2 13 10 11 3 1 10 9 12 1 10 9 1 10 9 2
42 2 1 10 0 9 2 9 13 2 2 13 2 13 10 9 2 13 10 9 1 10 9 7 13 3 2 16 3 13 9 2 2 13 1 10 11 10 9 1 10 11 2
48 2 3 3 13 10 9 1 10 9 1 10 9 2 3 13 15 13 7 1 10 9 2 16 10 11 13 1 10 0 11 2 13 10 9 1 10 11 2 7 10 11 7 10 11 13 10 9 2
66 10 9 13 15 2 13 0 9 1 13 2 3 3 9 2 7 3 13 4 1 13 10 11 0 2 2 2 13 10 9 2 13 15 13 1 10 9 1 10 9 1 10 9 15 13 3 10 9 1 10 9 0 2 16 3 13 13 0 1 11 3 1 10 11 2 2
62 10 9 0 13 10 11 2 1 9 1 11 2 1 10 10 11 2 15 13 16 10 9 1 10 9 0 13 10 9 1 9 7 9 2 13 15 1 13 10 10 9 2 13 16 15 15 13 1 10 11 13 10 9 0 1 10 9 0 7 10 11 2
35 7 2 1 10 9 1 9 2 3 13 13 1 10 10 9 1 9 2 11 2 2 11 13 3 13 13 1 2 3 0 2 10 9 0 2
7 10 0 1 10 10 9 2
12 11 2 1 12 9 1 10 0 1 10 11 2
30 12 1 10 12 9 13 0 2 12 1 10 12 9 3 13 9 7 3 12 1 10 12 0 13 13 10 9 1 9 2
14 15 13 10 9 3 0 1 10 11 1 10 9 0 2
51 9 2 3 1 15 13 1 10 9 1 10 9 2 13 10 9 15 10 9 7 10 9 0 13 1 10 11 7 15 13 1 13 1 10 9 1 10 9 1 9 2 3 1 15 13 1 10 9 1 9 2
21 3 13 16 10 0 9 2 13 1 10 9 3 0 2 13 1 13 10 9 0 2
15 9 2 13 16 13 10 9 3 0 2 15 15 13 13 2
19 7 13 15 15 9 2 3 10 9 1 10 9 7 10 9 1 10 9 2
25 11 13 2 1 10 9 2 10 9 1 10 11 7 11 3 13 1 10 9 1 10 13 9 12 2
47 13 1 10 9 1 10 9 15 13 1 10 9 7 3 13 10 10 9 1 9 2 13 0 9 10 9 1 15 13 9 1 13 10 10 9 2 3 3 10 2 9 0 2 2 1 9 2
12 7 3 10 9 1 13 10 9 1 10 9 2
16 13 10 10 9 1 13 1 13 1 10 9 13 1 10 9 2
44 1 10 9 1 11 2 3 3 13 3 12 9 1 13 1 9 2 11 13 1 10 2 9 7 9 0 1 10 9 0 2 1 2 13 16 3 15 13 13 10 9 3 2 2
19 2 3 13 9 7 13 9 13 0 16 15 3 13 3 10 9 13 0 2
13 3 13 1 13 16 3 15 13 13 15 3 2 2
25 10 9 2 1 10 0 9 2 2 13 16 13 10 9 1 13 15 13 10 9 0 2 2 13 2
1 11
4 9 1 9 0
33 1 9 1 10 9 2 10 9 0 1 10 11 1 11 2 11 2 13 3 10 9 1 11 1 9 1 10 9 1 10 9 0 2
38 1 10 9 2 12 9 13 2 2 10 9 13 10 9 1 10 9 1 15 12 1 10 9 2 13 3 13 10 9 3 1 13 2 10 9 0 2 2
7 9 1 10 11 13 1 11
6 1 10 9 1 10 11
49 1 10 9 1 10 11 2 3 1 9 1 10 9 13 1 12 2 10 9 1 10 9 1 10 9 0 1 10 11 13 1 13 15 1 3 2 1 11 2 1 13 13 3 10 9 1 9 0 2
8 7 15 13 1 10 9 0 2
3 2 0 2
12 1 10 9 3 13 10 9 0 1 10 9 2
32 15 13 13 13 9 2 13 9 13 1 13 1 10 9 1 9 2 13 13 1 10 9 9 1 9 13 2 13 13 1 11 2
13 2 1 10 9 2 0 2 3 1 13 10 11 2
9 2 13 2 3 2 10 9 0 0
51 10 9 13 1 11 13 15 1 16 10 9 2 1 13 9 2 2 13 13 3 10 10 9 2 2 13 16 2 10 9 13 1 15 13 1 10 9 16 10 9 3 13 15 1 13 1 10 9 13 2 2
16 2 16 3 15 13 10 9 2 10 9 13 13 10 9 2 2
50 1 10 9 1 10 9 1 10 9 0 0 2 10 9 0 13 0 1 13 16 2 10 9 13 13 2 2 1 10 2 9 1 10 9 1 10 9 2 2 3 16 2 10 9 3 13 7 13 2 2
19 1 10 10 9 2 15 13 15 1 10 9 1 15 10 9 0 13 13 2
19 2 3 1 10 9 1 10 9 2 13 0 16 10 11 15 13 13 2 2
4 9 1 10 11
4 11 13 1 11
36 10 11 13 13 1 1 10 9 1 9 12 0 9 1 10 9 1 10 9 0 1 9 2 1 2 13 10 9 2 1 10 9 1 9 0 2
45 10 9 11 2 3 13 2 13 3 13 1 10 9 1 11 1 10 11 1 10 11 2 7 13 1 10 9 1 9 0 7 1 10 9 1 10 9 1 9 1 10 9 1 9 2
20 10 9 1 10 9 13 13 1 10 9 1 11 1 10 9 7 1 10 9 2
26 10 9 1 10 9 1 10 11 13 16 2 10 0 9 1 10 9 1 9 13 3 13 7 13 2 2
17 2 13 0 13 10 9 1 10 9 7 13 10 9 2 2 13 2
22 10 9 3 13 13 3 10 9 2 15 13 9 1 10 9 1 10 9 0 1 9 2
31 3 1 10 9 2 12 9 1 10 9 2 13 1 10 9 11 10 9 1 9 2 9 0 7 3 12 9 1 10 11 2
33 10 9 13 3 12 9 1 13 10 9 1 10 9 1 9 2 3 1 13 10 9 11 7 2 3 2 13 10 9 13 1 11 2
42 10 9 1 10 0 2 3 1 13 10 9 1 10 9 1 10 11 2 3 13 13 1 10 9 1 10 9 11 7 3 13 1 1 10 9 1 10 11 1 10 11 2
42 1 13 10 9 1 10 9 2 13 13 1 10 9 1 10 11 1 10 11 2 13 1 10 10 9 1 0 2 3 0 1 10 0 9 1 10 9 1 10 9 13 2
23 2 15 13 10 9 2 2 13 10 9 1 10 11 2 3 1 13 10 9 1 10 9 2
23 10 0 9 1 10 9 13 13 1 10 9 11 7 1 10 9 11 2 15 1 12 9 2
34 15 2 9 1 10 9 1 9 1 12 7 0 1 10 2 9 2 0 2 13 15 3 3 10 0 9 1 10 9 1 10 11 0 2
32 16 3 13 12 9 1 9 2 10 9 13 16 10 10 9 1 9 13 0 2 3 1 15 13 10 9 13 1 10 0 9 2
16 10 9 13 0 1 11 7 0 1 10 11 2 11 7 11 2
27 10 10 2 9 2 1 10 9 1 10 0 9 1 10 11 2 13 1 10 9 1 12 9 1 10 9 2
14 10 9 1 12 9 2 1 10 9 1 12 1 9 2
31 3 0 13 1 10 11 2 10 0 9 1 10 9 0 13 15 13 11 1 10 0 9 1 10 9 0 1 10 9 0 2
9 3 13 10 0 9 1 10 9 2
28 11 2 10 9 1 11 2 1 10 9 2 13 10 0 9 1 9 2 13 10 12 9 1 9 1 10 9 2
16 3 2 13 3 2 13 12 2 9 2 1 10 12 9 0 2
38 13 15 10 9 1 0 9 2 1 15 13 12 2 9 2 2 15 15 13 13 10 9 1 10 9 1 10 12 9 1 10 12 0 9 1 10 9 2
16 10 9 2 15 13 10 0 9 1 10 9 0 2 13 0 2
18 2 16 13 3 3 2 3 2 2 10 9 1 10 9 13 0 2 2
14 9 2 3 13 9 0 2 3 13 1 10 9 0 2
11 13 16 3 13 9 1 10 9 1 3 2
13 10 9 1 10 9 13 10 9 1 10 9 0 2
8 2 9 2 2 13 10 9 2
21 13 13 1 10 15 16 13 13 15 1 10 9 2 3 1 15 2 7 1 15 2
14 10 9 13 1 15 7 3 15 3 13 13 9 10 2
8 13 10 0 9 15 2 9 2
5 15 13 1 13 2
21 15 15 13 1 15 13 10 9 1 10 15 13 7 15 10 15 13 2 7 3 2
13 16 10 9 13 9 3 13 16 15 13 10 9 2
17 7 16 10 9 13 1 9 2 3 13 16 13 13 10 0 9 2
27 11 13 1 10 11 13 1 10 9 7 16 13 13 10 9 3 2 13 10 9 1 9 13 1 10 9 2
19 3 2 10 9 1 10 9 1 10 11 2 13 13 1 9 1 10 9 2
47 7 2 13 11 2 10 11 13 10 9 1 13 10 9 0 15 13 1 10 11 13 10 9 0 7 12 9 1 9 2 1 13 10 9 1 10 11 2 1 10 9 1 9 1 10 11 2
40 11 2 1 12 9 2 9 1 0 7 0 9 0 2 12 2 1 10 9 2 13 1 10 9 13 10 9 7 13 13 1 10 10 9 3 1 10 0 9 2
60 10 10 9 2 13 1 10 9 0 11 7 11 2 3 15 13 2 7 10 9 13 3 15 1 10 10 9 2 1 10 9 1 11 1 10 9 0 2 1 9 3 1 13 2 7 1 10 0 1 10 9 1 10 9 2 11 2 3 9 2
33 13 10 9 1 9 2 1 11 2 15 13 10 9 2 0 2 16 13 10 9 1 10 9 13 1 12 9 2 2 1 13 11 2
3 7 13 2
28 2 3 13 1 10 11 3 13 3 9 1 9 13 2 13 10 9 0 1 10 9 7 13 3 15 1 13 2
28 3 10 12 9 13 10 9 1 12 7 12 9 7 13 13 2 1 15 2 3 10 11 13 13 3 9 2 2
34 11 13 3 10 9 1 10 9 1 10 9 15 13 1 10 9 1 10 9 3 15 13 3 1 10 0 2 1 13 1 4 3 13 2
15 2 3 1 10 9 13 13 1 10 9 1 10 9 2 2
4 11 1 10 11
10 2 13 0 13 10 11 1 10 9 2
50 9 2 1 12 1 12 2 7 9 1 10 11 2 1 10 9 1 10 9 1 12 2 11 13 2 3 2 10 9 1 10 11 1 10 11 2 10 0 0 9 0 1 11 2 1 13 1 10 9 2
49 9 0 2 3 3 15 13 10 9 1 10 0 9 2 13 1 10 9 1 10 9 7 1 10 9 2 1 10 11 0 7 10 11 0 2 11 13 16 10 9 1 9 0 13 1 11 13 0 2
50 13 0 10 0 9 0 1 10 11 2 3 3 1 10 9 1 10 11 2 13 1 12 2 7 2 1 15 13 2 10 9 1 10 11 13 1 16 15 15 13 1 10 0 9 1 9 7 1 9 2
7 2 3 3 13 13 3 2
15 13 10 9 13 1 9 2 10 9 13 2 10 9 13 2
15 1 10 9 2 3 13 10 9 2 13 1 10 9 2 2
5 3 0 7 0 2
13 10 0 9 13 1 10 9 2 1 10 9 0 2
28 13 10 0 9 7 13 2 10 11 1 10 9 1 10 9 12 2 13 2 10 0 9 1 11 7 11 2 2
49 13 10 9 1 10 9 0 2 11 15 2 3 2 2 3 13 13 10 9 1 11 7 11 7 2 3 2 13 10 9 3 0 1 10 9 13 1 10 9 0 7 1 10 9 0 7 0 2 2
3 9 2 11
3 9 2 11
1 9
5 12 7 0 9 2
38 1 10 9 7 9 1 9 11 3 1 10 9 3 11 13 10 10 9 2 3 1 13 4 13 1 10 10 0 9 1 10 9 13 1 10 9 11 2
42 11 13 10 9 1 10 9 2 15 3 13 1 10 9 2 1 10 9 3 1 2 11 2 2 3 13 0 9 1 2 11 2 2 2 11 2 2 2 11 2 2 2
23 7 10 9 13 1 13 1 10 9 0 2 1 10 9 1 10 9 1 10 9 1 9 2
24 10 11 13 3 10 9 1 10 12 9 1 15 13 3 1 10 12 9 1 10 9 1 9 2
26 3 1 9 0 2 10 11 13 1 9 0 1 1 10 12 9 2 1 1 10 9 0 13 1 13 2
19 15 1 10 9 0 1 3 13 13 10 9 0 1 10 9 1 10 9 2
28 1 10 9 13 10 9 1 10 9 1 9 0 2 15 1 9 13 3 12 9 2 13 10 9 1 9 0 2
39 1 10 9 1 9 2 1 15 13 1 10 12 9 2 3 12 9 16 1 10 9 0 2 10 9 11 13 9 1 10 9 1 10 12 9 1 10 9 2
4 9 2 9 0
37 11 13 1 13 9 0 1 10 9 3 13 13 10 10 9 0 1 10 9 1 9 13 1 13 10 9 1 10 9 7 13 15 10 9 3 0 2
10 11 3 2 1 10 0 7 13 9 0
38 10 9 13 13 0 7 10 10 0 9 7 10 9 13 3 13 13 10 10 12 9 7 2 3 3 2 9 1 9 13 1 13 15 3 15 13 12 2
26 10 9 11 13 3 3 12 0 2 9 2 1 12 9 1 10 9 2 1 9 1 10 10 0 9 2
4 9 1 10 11
41 10 9 1 10 9 1 9 12 1 10 11 13 1 10 9 1 10 9 7 1 10 9 1 10 9 9 2 15 13 1 13 10 9 1 10 9 1 10 9 0 2
15 3 13 13 12 9 1 10 9 11 2 1 10 9 0 2
51 3 2 10 11 13 1 13 9 1 9 7 13 10 9 1 10 9 1 10 11 2 3 1 10 2 9 2 1 10 9 2 15 3 13 2 7 13 10 9 16 10 10 2 7 1 10 9 15 3 13 2
36 10 9 13 3 7 15 2 1 12 9 2 13 12 9 1 9 1 10 0 2 10 11 2 15 3 13 1 10 11 7 3 13 1 10 11 2
29 10 11 2 10 9 2 13 13 3 1 10 11 7 13 3 10 9 1 10 10 9 13 1 13 15 10 0 9 2
29 10 11 13 1 13 10 9 1 10 11 2 3 2 10 9 0 7 1 9 2 7 3 13 10 11 1 10 11 2
37 10 11 13 1 13 7 13 1 15 15 13 1 13 3 13 9 1 10 11 2 1 10 9 15 3 13 13 1 10 9 1 10 9 1 10 9 2
21 10 11 2 1 11 1 9 2 2 13 2 10 9 1 9 1 10 9 1 11 2
22 10 11 13 13 1 10 9 1 10 11 7 13 10 10 9 1 9 13 1 10 11 2
38 13 3 10 9 3 10 9 1 9 7 9 13 1 13 3 13 7 2 1 10 9 1 10 0 9 1 9 2 10 9 1 10 9 13 15 13 0 2
18 1 1 11 2 12 9 1 9 2 15 13 13 0 9 1 10 9 2
5 6 2 6 7 6
25 10 0 9 1 9 1 9 1 9 2 9 7 9 13 10 9 13 1 10 9 1 10 9 0 2
49 10 9 13 3 13 1 10 9 1 10 9 11 12 1 3 13 12 9 13 2 13 13 1 10 9 2 13 15 0 7 0 2 13 13 0 2 1 10 9 1 9 1 10 9 1 10 0 9 2
13 1 10 11 2 1 10 9 2 13 15 10 11 2
1 9
39 1 10 11 13 13 2 3 1 10 9 1 10 9 1 10 11 2 10 9 0 2 11 2 2 1 9 1 11 2 11 2 11 2 11 2 11 7 11 2
4 1 10 9 2
1 11
5 11 13 9 1 9
58 10 9 0 1 10 11 2 10 9 0 1 11 10 9 15 13 1 9 1 10 13 9 2 13 1 10 11 1 11 10 9 1 10 9 13 3 1 10 9 7 15 13 1 10 9 1 10 9 1 12 9 1 10 9 13 1 9 2
5 9 0 13 10 9
78 1 10 9 1 3 1 10 11 2 15 13 9 1 10 0 9 1 9 1 9 1 9 2 10 11 13 1 3 4 10 9 0 1 9 7 1 4 13 10 9 0 2 13 2 3 2 10 9 1 9 1 1 10 9 1 12 9 1 9 2 1 12 9 2 1 9 1 9 1 9 1 9 1 10 9 1 11 2
13 11 2 10 9 1 10 9 7 10 9 3 13 2
10 13 2 1 0 9 2 3 3 13 2
16 1 12 1 9 1 12 3 13 13 1 10 9 9 10 9 2
26 15 3 13 13 1 0 9 2 3 1 9 0 1 9 1 12 2 7 3 13 2 1 3 2 9 2
20 10 9 2 1 9 0 2 3 0 2 13 13 1 10 9 9 1 10 9 2
31 3 3 0 2 10 9 3 3 13 13 13 1 10 9 2 15 3 13 1 13 0 13 3 10 9 13 1 10 0 9 2
5 9 2 7 3 2
113 1 11 2 11 13 3 16 10 9 0 1 9 1 10 11 13 10 9 1 10 9 11 2 11 2 7 3 3 10 9 1 10 11 2 1 10 9 15 3 13 1 11 7 10 9 15 15 3 13 13 12 9 1 10 11 2 10 9 11 2 11 7 10 0 9 1 10 11 1 11 7 1 3 1 11 7 11 2 11 2 2 7 3 10 9 1 10 11 2 11 2 11 2 13 10 9 13 3 13 2 3 10 9 1 10 11 7 10 0 9 1 11 2
22 15 13 1 10 11 2 1 10 9 0 1 11 2 1 15 13 1 9 1 10 9 2
25 3 3 11 13 13 3 10 9 2 1 10 0 9 1 16 10 9 13 1 10 9 3 7 3 2
18 2 3 1 10 9 1 10 9 0 1 10 9 2 3 13 9 2 2
31 7 13 10 9 1 13 2 1 10 10 9 2 1 10 0 9 1 10 9 2 10 0 9 3 0 1 13 10 0 9 2
20 7 13 2 1 10 9 0 2 10 9 0 1 11 2 13 1 3 12 9 2
4 3 10 0 2
4 11 1 10 11
10 2 3 13 15 13 1 11 13 2 2
36 1 13 1 9 2 13 13 16 10 9 0 1 13 1 10 11 13 10 0 9 2 1 15 12 13 2 1 9 7 9 2 10 9 1 9 2
26 3 0 2 1 10 0 0 9 2 15 3 13 13 1 15 12 2 13 10 9 1 12 9 1 9 2
41 10 11 2 10 11 2 10 11 2 10 11 2 10 11 2 10 11 2 10 11 7 10 11 13 15 1 10 15 3 13 7 2 13 15 2 0 9 13 1 13 2
66 16 1 15 13 15 13 1 4 13 2 9 7 9 1 10 11 2 9 1 10 11 7 1 10 11 2 9 1 10 9 2 11 7 11 2 2 9 1 10 9 2 11 7 11 2 2 0 1 10 9 1 9 2 3 15 1 11 2 2 2 10 9 13 13 9 2
40 3 13 1 9 1 10 11 2 9 7 9 1 9 13 10 9 1 10 9 2 1 11 2 1 11 2 10 9 1 10 11 13 3 1 9 13 1 10 9 2
20 13 2 16 2 13 10 9 1 9 2 7 13 15 1 10 2 0 9 2 2
30 3 13 1 13 10 9 1 10 9 1 10 11 2 2 15 3 13 10 1 10 9 2 2 13 1 10 9 7 9 2
12 3 15 13 1 13 3 3 3 13 3 0 2
15 10 9 3 13 1 13 1 10 11 7 1 10 10 9 2
14 2 3 13 2 13 2 2 13 10 0 1 10 9 2
8 13 10 9 13 2 9 0 2
24 7 3 2 10 9 13 2 1 10 9 13 1 10 2 11 0 1 10 9 1 10 9 2 2
24 7 10 0 1 10 9 13 15 13 12 9 2 1 11 2 3 13 1 10 0 9 1 11 2
16 9 13 9 0 1 12 1 12 9 1 10 11 7 13 1 9
10 11 1 10 9 1 10 9 1 10 9
37 11 2 9 7 0 9 2 13 13 4 13 1 10 9 1 11 1 10 9 0 7 1 9 1 10 11 2 1 13 10 9 1 3 1 10 11 2
17 2 3 13 1 10 9 2 7 13 13 1 10 9 2 2 13 2
8 3 2 10 9 3 13 15 2
7 11 13 1 2 9 2 2
8 13 2 9 2 1 10 9 2
15 3 13 10 0 9 15 15 13 13 2 15 1 10 9 2
15 7 1 15 15 2 1 13 12 9 1 3 2 15 13 2
6 2 13 2 9 9 2
4 13 13 3 2
30 3 13 10 9 3 0 2 7 15 13 3 2 1 13 13 10 9 2 2 2 13 15 1 10 9 15 15 13 13 2
13 3 2 10 0 9 2 10 0 9 13 15 3 2
37 7 13 1 10 9 1 13 2 3 2 0 2 16 10 9 1 10 9 13 10 9 1 12 9 2 9 7 9 2 13 3 2 1 13 12 9 2
10 15 13 16 3 15 13 10 10 9 2
19 7 3 13 16 13 1 10 9 3 15 13 1 10 10 9 10 0 9 2
5 3 13 10 9 2
26 3 13 10 0 9 1 9 1 13 3 2 7 1 9 0 2 10 9 1 10 9 7 1 10 9 2
28 1 0 15 13 2 13 15 10 9 0 1 15 13 0 1 10 2 9 1 10 11 2 1 15 15 13 9 2
2 11 2
24 9 1 9 1 11 13 10 9 1 10 9 1 10 9 0 9 15 13 1 10 9 1 11 2
9 15 13 3 10 2 9 0 2 2
13 7 15 15 13 3 1 10 9 13 2 0 2 2
101 1 10 9 2 7 3 1 11 2 12 9 2 10 9 1 10 2 9 2 1 10 2 9 2 2 10 9 1 13 2 9 2 1 2 9 2 2 7 3 10 9 1 13 10 9 1 10 9 2 10 0 2 9 1 9 2 1 10 15 13 3 0 13 16 10 9 13 13 2 7 10 9 1 9 2 1 10 15 13 3 0 13 16 10 2 9 2 2 3 2 0 2 2 13 13 0 2 1 9 2 2
6 13 15 3 1 9 2
3 7 9 2
33 7 13 13 1 9 2 7 13 13 2 3 2 1 10 9 1 9 13 1 10 9 1 10 9 2 15 13 10 9 1 10 9 2
37 9 0 2 7 3 9 2 1 10 10 9 13 1 10 9 13 13 1 10 9 0 1 12 9 2 3 13 1 10 11 2 0 11 2 1 9 2
24 10 10 9 13 3 3 9 1 12 9 1 12 9 0 2 15 15 13 13 1 10 10 9 2
1 11
4 9 1 10 9
38 0 0 1 10 11 7 1 10 11 13 3 13 13 10 9 1 10 12 9 1 10 0 9 0 15 13 12 0 1 9 1 10 9 13 1 10 11 2
33 10 9 7 9 0 2 11 2 13 13 15 3 1 10 11 1 13 13 10 9 2 13 1 10 11 10 9 1 11 2 9 0 2
27 13 9 1 11 2 12 2 7 3 13 13 10 10 0 9 2 16 3 3 15 13 13 3 1 10 0 2
21 11 13 16 3 13 10 9 3 1 9 7 13 11 1 13 10 11 3 10 9 2
16 10 9 0 1 15 12 13 3 0 16 10 9 1 10 9 2
10 11 2 10 0 2 11 2 10 0 2
29 11 13 1 11 2 11 2 2 1 12 2 7 13 15 1 10 11 2 1 3 13 10 9 1 10 9 0 0 2
29 13 0 1 11 2 1 12 1 12 2 3 13 12 9 7 2 1 12 2 13 1 10 9 3 9 1 10 11 2
16 1 10 9 2 1 10 9 1 10 9 2 13 1 13 0 2
19 10 0 9 13 15 10 9 1 12 9 1 10 9 2 1 12 1 11 2
1 11
30 10 9 0 1 10 11 2 11 2 3 15 13 3 3 10 2 9 1 10 9 2 1 10 9 1 10 10 9 11 2
9 7 15 13 1 16 13 10 9 2
19 16 1 10 9 10 9 15 13 10 0 9 2 3 13 3 0 16 11 2
12 11 2 12 9 2 13 1 10 11 1 12 2
22 3 13 0 1 10 11 2 9 0 2 9 1 10 11 7 9 1 11 1 10 11 2
10 13 3 9 7 2 9 2 1 11 2
27 1 10 11 2 13 13 10 9 2 13 10 9 1 10 2 0 9 0 1 1 10 9 1 10 9 2 2
19 10 9 1 10 11 13 15 1 10 11 1 11 1 13 10 9 1 11 2
17 1 10 9 3 13 2 3 2 10 9 0 1 10 2 9 2 2
35 10 9 1 9 0 2 10 9 1 10 9 2 9 1 15 3 11 13 0 1 0 2 13 9 1 10 0 15 15 13 1 10 0 9 2
44 10 12 9 1 10 11 1 3 12 1 10 11 2 1 10 9 0 2 13 3 10 9 1 10 9 0 1 10 9 1 11 7 3 13 1 15 10 9 0 1 10 10 9 2
16 1 10 0 9 2 10 9 1 10 9 13 1 13 10 15 2
17 11 13 15 2 1 15 2 1 13 1 10 9 13 11 1 11 2
35 1 10 9 1 11 2 10 0 9 1 10 11 13 13 9 0 1 10 9 2 13 16 10 10 9 15 13 3 0 1 10 9 1 9 2
17 16 3 0 2 10 9 1 10 11 3 13 13 10 10 9 0 2
16 3 10 9 11 2 10 9 2 13 2 3 2 10 9 0 2
56 10 9 7 9 1 10 9 1 9 1 9 1 11 7 11 13 1 10 9 1 10 11 11 2 10 9 1 10 9 11 11 2 15 13 2 1 1 10 9 1 12 2 13 10 9 1 12 12 9 1 10 9 1 10 11 2
16 10 9 11 13 1 10 9 1 10 11 9 2 1 15 13 2
62 13 10 9 0 1 12 12 9 0 3 1 10 9 1 11 2 11 2 2 11 2 11 2 2 11 2 11 2 2 11 2 11 2 2 11 7 11 2 11 2 7 11 2 11 2 1 10 11 2 10 9 0 1 10 12 9 1 9 1 10 11 2
32 13 3 12 9 1 9 1 15 12 9 0 13 1 10 11 13 10 9 1 9 1 10 9 1 10 9 7 9 11 7 11 2
54 10 9 1 10 2 9 0 2 2 9 2 9 2 2 1 10 9 7 1 10 2 9 1 10 9 0 2 2 3 10 10 2 9 2 1 10 9 1 10 2 9 2 7 1 10 2 9 2 13 15 1 10 9 2
34 2 11 2 13 3 10 9 1 10 9 1 15 11 13 1 11 2 1 10 9 12 2 3 13 10 9 2 10 9 1 11 7 11 2
34 3 2 11 13 15 1 9 1 9 2 1 10 9 2 12 2 1 11 2 1 10 9 0 2 7 3 1 10 10 9 2 1 11 2
36 1 12 2 1 10 11 2 13 10 11 2 1 12 2 1 10 11 2 11 2 13 15 3 1 9 2 1 10 11 7 1 12 13 10 11 2
35 3 1 10 9 1 10 9 2 13 10 9 1 10 11 2 1 11 2 7 13 10 9 1 9 7 10 11 2 1 12 2 1 10 11 2
23 1 10 0 9 1 9 1 12 9 2 1 10 9 1 9 2 7 11 7 11 13 0 2
45 2 13 3 13 9 16 2 1 13 1 10 9 2 11 2 7 1 10 10 9 2 1 16 13 9 0 1 10 9 1 9 3 13 2 3 13 1 13 10 9 2 2 13 11 2
20 2 10 9 11 13 3 1 13 10 9 2 2 13 2 1 10 9 2 11 2
35 1 10 11 13 2 10 11 13 1 10 11 10 9 1 10 0 9 2 3 15 13 16 10 9 1 10 9 2 1 9 2 13 1 12 2
27 10 9 3 0 1 10 9 1 10 2 9 1 9 2 2 1 12 9 2 1 10 0 9 1 12 9 2
23 15 13 2 10 11 13 16 10 12 9 1 13 13 2 7 3 13 10 9 1 10 9 2
23 11 2 9 2 3 13 2 3 13 2 1 10 9 13 1 10 9 0 1 10 9 11 2
11 7 1 15 13 10 9 0 1 10 9 2
15 13 15 10 9 13 1 10 11 1 10 9 1 10 9 2
54 11 13 2 3 1 15 2 16 10 9 3 10 11 13 13 10 9 13 2 0 2 2 3 2 1 10 9 11 2 10 2 9 2 13 10 0 13 1 10 9 13 2 7 3 1 10 9 1 10 9 1 10 9 2
48 1 10 9 3 15 1 10 9 2 1 15 10 9 1 9 13 4 7 4 1 9 13 3 2 10 9 0 13 2 1 10 9 1 11 2 13 1 16 10 9 15 13 3 1 10 9 0 2
31 3 2 10 9 13 10 9 1 11 13 10 0 9 15 13 1 15 10 9 1 11 13 13 1 13 10 9 1 12 9 2
37 1 10 9 1 10 9 0 1 10 9 1 10 9 2 12 9 1 10 9 13 16 13 0 1 12 9 2 16 12 9 13 9 0 1 12 9 2
99 13 10 9 2 10 11 13 16 2 2 16 13 10 9 16 1 10 9 2 9 0 2 1 9 2 9 7 9 2 0 7 3 0 2 15 13 10 9 1 9 1 15 10 9 0 13 0 1 12 9 1 10 9 1 9 2 13 3 0 10 9 1 10 0 1 10 9 13 10 9 9 0 2 9 1 10 12 7 15 12 9 2 12 9 1 10 9 2 7 12 9 13 9 0 1 12 9 2 2
4 9 1 10 9
19 1 10 9 2 1 9 1 10 9 2 1 11 2 10 9 13 3 0 2
18 1 10 9 2 1 10 10 9 2 1 11 2 10 9 13 3 0 2
24 16 10 10 0 9 2 2 11 2 2 3 13 10 9 1 10 9 2 2 11 2 13 15 2
18 7 2 3 1 15 13 1 10 9 2 12 13 15 12 9 1 9 2
1 11
1 11
34 9 1 10 9 1 12 9 7 9 1 10 9 1 10 11 2 11 13 12 1 10 9 1 10 9 1 10 0 9 0 1 10 11 2
25 1 13 1 9 1 12 7 13 1 9 1 12 2 13 12 9 2 10 9 13 10 9 1 9 2
1 11
9 9 1 9 7 9 1 10 9 0
5 11 13 13 1 11
14 10 11 13 13 10 9 3 1 10 9 0 1 11 2
41 10 9 13 13 3 2 3 1 10 9 1 10 9 1 10 9 15 15 13 1 10 9 1 9 1 10 9 2 13 15 1 10 9 0 3 13 13 3 12 9 2
28 15 13 12 1 10 12 9 15 10 9 13 1 9 1 10 9 15 13 3 13 13 3 10 9 1 10 9 2
23 3 2 13 3 1 10 9 10 9 13 1 10 9 1 10 9 1 10 9 1 10 9 2
20 13 15 16 10 10 9 13 3 13 1 10 0 9 16 10 9 3 13 13 2
4 9 13 1 9
27 10 11 13 1 13 10 9 1 11 2 1 12 9 2 10 9 13 13 2 3 3 2 1 11 2 11 2
55 11 2 10 2 0 2 1 10 11 0 2 15 13 9 1 10 0 9 7 13 3 9 2 13 10 9 1 9 9 1 10 0 9 0 2 15 13 2 1 9 1 9 2 10 9 11 7 11 2 9 1 10 9 11 2
36 10 2 9 2 0 3 13 9 1 9 2 2 3 9 1 10 9 0 13 1 9 0 2 2 16 2 10 9 13 0 2 7 13 9 2 2
5 2 13 10 9 2
38 1 10 12 9 2 11 2 2 11 2 2 2 11 2 1 10 2 9 2 1 10 11 7 1 10 11 2 3 13 13 7 13 1 9 1 10 9 2
28 3 13 10 9 1 10 9 1 10 11 7 1 10 9 1 10 11 7 3 13 2 10 9 1 10 9 2 2
53 3 2 1 12 9 15 13 15 3 2 13 15 3 10 9 1 10 2 9 2 1 10 11 2 11 2 2 2 3 12 9 1 9 15 13 3 13 7 15 13 15 1 10 15 2 2 7 13 3 10 10 9 2
34 2 10 10 9 13 3 13 1 10 11 2 10 9 1 9 1 15 13 9 2 1 15 9 1 10 2 9 2 7 1 10 9 2 2
7 9 13 11 16 13 0 13
8 3 10 9 13 15 3 13 2
54 7 3 0 3 3 15 13 3 1 10 9 3 2 3 1 13 10 9 2 1 13 1 9 2 2 2 7 3 13 3 10 10 9 2 13 15 2 3 13 3 3 2 2 2 7 13 15 1 10 9 1 10 9 2
8 3 13 13 9 7 13 9 2
16 3 13 10 9 1 10 9 15 13 3 1 10 9 1 11 2
10 13 10 9 9 2 3 6 2 2 2
11 10 9 1 10 9 1 9 13 10 9 2
6 3 13 1 15 13 2
21 7 3 15 13 10 0 9 1 10 9 15 13 16 10 9 0 13 10 9 13 2
8 7 3 13 3 13 15 13 2
11 1 9 2 3 15 13 13 3 7 3 2
6 3 13 0 10 0 2
28 1 10 9 10 9 13 15 2 10 9 7 10 0 0 2 10 11 2 11 2 7 10 11 2 9 7 9 2
18 9 2 9 1 9 2 9 0 7 10 9 13 15 11 13 1 13 2
3 13 15 2
2 9 13
20 3 1 12 9 1 13 10 9 10 9 13 15 3 2 3 1 9 7 9 2
26 10 0 13 13 1 10 9 1 10 9 1 10 9 3 13 10 9 2 7 10 9 2 1 9 0 2
28 13 12 1 10 0 9 1 10 9 15 10 9 1 11 13 1 10 13 9 0 2 7 10 0 9 1 9 2
6 9 1 10 11 1 9
4 10 9 1 11
33 13 1 10 9 0 2 13 1 10 13 9 12 1 9 2 1 11 2 10 9 11 2 12 1 10 0 9 0 1 10 9 0 2
20 10 9 1 10 10 9 3 3 13 13 2 3 1 10 9 0 2 11 2 2
25 10 0 9 13 13 15 1 10 9 1 11 2 1 12 12 9 2 3 1 11 13 3 12 9 2
20 1 10 9 1 12 1 9 1 12 1 9 10 9 13 13 1 12 9 0 2
49 3 2 10 0 9 15 13 9 1 10 9 1 10 11 2 1 10 9 1 11 7 11 2 13 1 13 15 1 10 9 1 3 2 1 13 4 13 13 1 10 9 2 1 9 1 10 9 0 2
36 3 2 13 1 10 11 2 1 10 9 1 10 10 0 9 0 1 10 11 2 11 13 1 13 10 9 1 10 9 1 10 11 1 9 0 2
18 15 13 2 13 15 13 13 1 10 0 12 9 2 15 11 13 0 2
29 11 13 1 10 9 0 2 11 2 16 13 1 10 9 2 9 0 7 9 2 16 2 13 10 9 1 10 9 2
37 10 9 13 16 2 1 11 2 10 9 13 3 1 10 9 1 10 9 1 10 11 1 10 11 2 3 1 11 13 0 1 10 9 1 10 11 2
28 2 15 13 16 13 13 15 1 10 11 2 7 1 10 9 0 13 15 2 3 15 13 2 2 13 15 11 2
18 2 10 11 13 3 10 10 9 7 2 1 10 9 2 13 15 2 2
6 9 1 10 11 1 11
5 10 9 1 10 9
17 1 10 9 13 10 9 2 1 10 9 13 10 9 7 10 9 2
31 10 12 9 1 10 11 1 10 11 13 15 1 10 9 7 9 2 13 3 3 1 9 2 16 10 9 15 13 1 9 2
9 15 13 10 0 2 15 7 15 2
6 11 2 13 1 3 2
6 11 2 13 1 3 2
1 11
8 13 1 13 15 1 10 9 0
31 12 2 10 9 13 10 9 0 2 0 2 1 15 10 9 13 9 7 3 13 13 3 1 10 10 9 7 9 2 2 2
6 2 15 13 10 11 2
8 15 2 1 11 2 15 3 2
5 3 10 9 13 2
9 2 13 12 9 3 1 10 9 2
20 15 13 1 10 9 2 3 3 15 1 0 13 1 10 9 2 7 13 15 2
47 13 7 13 16 13 10 9 1 9 2 15 3 13 9 2 7 3 13 2 11 2 3 13 3 2 13 15 10 9 1 10 9 2 3 13 16 13 2 16 13 0 2 16 13 10 9 2
21 3 13 13 2 11 2 2 7 15 15 13 3 13 7 10 9 13 1 13 2 2
16 12 9 3 2 13 11 2 1 10 9 1 10 9 1 11 2
16 2 15 3 13 9 7 15 3 13 2 2 7 3 13 2 2
20 16 15 13 1 10 9 1 11 1 10 9 1 15 2 13 15 15 13 13 2
13 10 10 9 13 15 2 13 13 15 1 10 9 2
9 3 15 13 2 3 13 0 2 2
28 3 15 13 15 13 10 0 9 1 10 9 3 0 1 10 9 2 11 13 15 16 13 16 13 12 9 0 2
8 2 12 1 15 13 10 9 2
29 13 10 9 3 0 1 9 1 13 1 10 9 0 7 15 13 13 10 9 1 13 9 1 10 9 0 0 2 2
47 3 3 13 1 13 2 3 2 16 10 0 9 1 10 9 13 0 1 10 11 2 10 9 3 0 1 10 9 2 3 10 9 1 10 9 13 3 0 16 1 10 10 9 1 10 9 2
22 2 3 2 2 13 11 2 2 10 9 13 1 13 1 9 3 0 3 10 9 2 2
16 10 9 1 9 1 10 0 9 0 2 3 2 13 3 0 2
46 1 10 9 2 15 13 10 9 1 9 1 9 0 2 3 12 9 1 9 2 2 7 1 12 1 12 9 1 9 10 10 9 13 1 10 9 0 2 1 3 12 12 9 1 9 2
6 0 9 3 1 10 11
5 11 13 10 9 11
22 10 9 13 10 9 0 1 10 9 1 10 11 2 15 13 10 9 1 10 9 0 2
25 1 10 9 0 2 10 9 13 0 2 13 16 10 9 1 10 9 11 2 10 9 0 1 9 2
7 2 7 0 1 10 11 2
44 1 10 11 2 15 13 13 1 10 0 9 1 10 11 2 1 15 13 13 1 10 9 1 10 9 1 10 9 2 13 12 1 10 12 9 1 9 13 1 10 9 1 11 2
27 10 9 1 10 11 13 3 3 16 16 11 13 1 15 1 10 9 1 10 10 9 13 9 1 15 13 2
33 10 9 1 9 3 13 2 13 10 11 2 13 1 13 10 9 1 10 9 1 10 9 1 10 0 9 12 2 9 1 10 9 2
32 3 1 10 0 9 1 9 2 13 13 12 9 2 10 11 13 13 10 9 0 1 10 11 1 13 1 13 10 9 1 11 2
33 7 3 1 10 0 9 0 2 1 9 1 9 2 9 7 9 1 9 2 10 9 0 1 10 9 13 16 3 13 13 1 3 2
31 10 9 1 3 2 13 1 11 2 10 15 15 13 10 9 1 9 0 2 13 1 15 2 16 10 10 11 13 13 0 2
39 13 10 9 0 1 10 9 0 1 10 9 2 11 2 9 0 2 13 10 9 1 10 0 7 10 0 2 10 9 7 10 9 2 10 0 7 10 0 2
6 3 2 13 9 0 2
7 1 15 2 13 9 0 2
56 13 10 9 10 9 1 9 1 10 9 2 13 16 2 10 9 2 1 10 9 1 9 15 13 3 12 9 1 9 2 10 9 1 10 9 1 10 9 7 9 1 10 9 16 10 9 1 10 10 9 2 1 10 10 9 2
9 13 10 9 13 10 9 1 9 2
43 13 10 9 1 10 9 0 1 10 9 13 13 10 9 0 7 13 1 10 9 7 3 13 2 1 15 13 13 10 9 1 10 9 2 13 10 9 13 15 10 0 9 2
3 10 9 13
24 3 10 9 2 13 3 1 9 15 13 9 1 10 10 9 2 3 1 9 13 13 10 9 2
27 3 13 13 10 10 9 13 1 10 9 3 0 7 13 1 10 9 16 13 13 10 9 1 15 13 9 2
35 1 10 9 2 13 15 1 10 9 1 9 1 9 1 9 7 1 9 1 9 0 3 13 1 10 9 2 13 11 1 12 1 9 2 2
50 13 1 10 11 3 1 10 9 1 10 11 2 10 9 3 13 10 9 1 13 11 2 3 1 10 9 1 10 11 2 7 11 2 3 9 1 10 11 2 10 9 15 13 10 12 11 0 3 13 2
57 13 10 9 0 2 10 9 0 11 2 9 1 10 9 2 3 13 9 1 13 16 10 11 13 10 9 1 9 1 10 2 9 7 9 2 13 1 10 9 1 10 9 1 10 9 1 10 11 7 1 10 9 1 10 10 9 2
35 10 11 13 3 7 10 11 2 3 1 10 10 9 1 10 9 1 10 11 2 11 2 13 3 10 9 1 13 1 13 10 9 1 11 2
43 2 3 1 13 10 9 1 10 9 11 13 1 10 9 0 1 10 9 0 7 13 16 13 3 10 9 15 10 10 11 3 13 2 2 13 11 1 10 11 13 12 9 2
28 3 2 3 2 10 11 13 10 9 1 9 13 1 10 9 1 13 3 10 9 1 10 9 1 10 10 11 2
6 11 13 9 1 10 11
26 2 13 1 10 11 13 10 9 0 1 10 9 2 13 12 9 3 3 13 3 10 9 1 10 11 2
31 13 1 10 0 9 13 10 9 2 7 2 13 15 1 10 9 2 13 13 1 13 10 9 3 10 9 2 2 13 11 2
8 11 2 1 10 11 2 1 11
10 10 12 9 1 10 0 9 1 10 11
39 10 9 1 10 9 1 10 9 1 10 2 3 13 2 0 9 0 1 10 11 2 11 2 13 9 0 1 10 9 1 3 1 10 11 2 1 10 11 2
8 1 10 11 13 13 10 9 2
32 3 12 12 9 13 1 10 11 2 2 9 2 3 13 1 10 11 2 3 13 3 3 12 12 9 2 9 0 1 10 9 2
20 10 9 1 10 9 1 10 9 13 1 10 9 1 11 10 9 1 0 9 2
11 2 1 3 2 10 9 13 0 1 9 2
9 10 9 13 10 9 2 2 13 2
11 10 9 13 2 3 2 10 10 0 9 2
18 2 7 13 10 9 1 10 0 9 3 2 2 13 2 1 0 9 2
28 13 9 1 15 2 16 10 9 13 15 3 10 9 1 3 12 9 2 13 3 2 10 10 9 1 10 9 2
26 2 1 10 9 1 10 9 2 13 1 10 9 10 9 7 10 9 1 13 2 16 13 3 13 2 2
31 3 13 13 9 1 10 10 9 2 11 13 3 10 9 2 13 3 10 9 2 13 10 9 7 3 13 13 10 10 9 2
34 3 2 13 1 13 10 9 1 10 10 9 2 15 2 1 12 1 10 9 0 1 11 2 13 13 15 10 9 2 13 15 10 9 2
25 2 15 13 3 1 15 16 2 3 13 1 9 3 13 16 3 13 15 2 13 15 7 13 0 2
7 1 15 13 2 2 13 2
9 10 9 1 11 3 13 3 0 2
15 10 9 0 1 10 9 1 10 0 9 1 10 11 13 2
23 10 9 13 3 13 9 1 10 9 1 10 9 1 10 9 2 10 11 7 10 10 9 2
25 2 10 0 9 1 10 11 13 4 13 1 10 9 1 10 9 2 2 13 11 2 10 9 0 2
8 9 1 10 9 1 10 11 2
33 10 9 15 13 10 9 1 10 9 1 11 2 11 2 1 13 10 9 7 10 9 0 13 3 1 0 9 2 1 13 10 9 2
17 11 13 16 10 9 0 13 10 0 9 1 9 13 1 10 9 2
52 1 10 9 13 1 10 10 0 1 10 9 1 10 9 0 2 1 11 2 13 9 1 10 9 1 10 9 1 10 9 1 10 9 1 10 9 2 10 9 1 9 1 10 9 1 9 7 10 9 1 9 2
19 9 15 2 3 1 11 2 10 11 7 10 11 1 10 11 13 13 13 2
5 9 1 10 11 2
34 10 11 13 15 1 13 10 9 1 10 9 1 13 1 10 11 7 9 0 2 13 10 9 1 10 9 1 9 13 1 12 12 9 2
36 10 9 2 1 12 9 7 12 9 3 2 13 15 1 10 9 1 10 9 1 10 9 0 1 10 9 2 13 3 1 10 11 7 10 11 2
27 10 9 2 11 2 13 10 9 0 1 10 9 0 1 10 9 2 13 10 9 1 10 9 1 9 0 2
27 1 9 2 10 9 1 9 1 12 9 13 13 1 10 9 0 1 13 10 9 1 10 9 0 7 0 2
71 1 10 9 1 10 10 9 0 1 10 9 0 2 10 11 2 11 2 13 10 9 1 0 9 0 3 2 3 2 1 10 9 7 9 2 1 9 0 2 1 10 9 0 2 1 10 9 0 2 9 2 9 7 9 2 7 2 3 2 3 2 1 10 9 0 2 1 10 9 13 2
38 3 11 3 2 1 0 9 13 1 12 1 9 1 12 2 13 10 9 1 15 11 2 1 10 9 0 1 13 2 10 9 0 1 0 7 13 2 2
18 10 9 13 1 13 1 10 9 10 9 15 2 3 2 3 3 13 2
28 3 2 3 1 10 9 0 2 10 11 13 10 0 1 10 9 0 1 10 9 7 10 9 13 1 12 0 2
6 1 11 13 9 0 2
14 1 10 9 13 1 10 9 10 9 1 9 1 11 2
14 12 9 3 3 10 11 13 10 9 1 10 9 0 2
28 1 10 11 2 11 2 11 2 1 10 2 13 2 1 10 9 2 1 10 9 13 1 10 9 2 11 2 2
12 10 9 1 9 11 13 10 9 2 11 2 2
9 11 13 10 9 1 10 9 11 2
12 1 10 9 2 1 10 11 2 1 10 11 2
14 1 10 9 13 1 10 9 13 10 11 7 10 11 2
31 10 9 2 1 9 1 9 15 3 13 3 11 2 13 10 10 9 1 10 9 3 9 2 12 9 2 7 10 0 9 2
27 9 1 9 2 7 1 12 9 1 10 9 7 1 12 1 10 9 0 2 10 11 2 10 1 10 9 2
27 13 3 10 9 1 10 11 1 10 0 2 9 2 2 3 15 1 11 7 11 2 15 3 13 10 9 2
28 9 0 2 10 9 1 10 0 11 2 13 1 10 9 2 13 3 3 9 1 9 2 13 3 1 4 13 2
55 3 1 10 11 2 1 10 9 13 3 2 13 13 1 10 11 1 10 9 1 12 9 1 9 1 11 2 2 1 3 13 10 9 15 15 13 1 10 9 13 1 10 9 2 10 9 11 13 1 10 9 1 10 9 2
32 13 15 16 1 9 2 3 10 9 1 10 9 13 10 9 1 10 9 7 10 9 3 13 10 9 1 10 9 1 10 9 2
1 9
5 10 9 1 10 9
25 3 13 1 9 1 15 3 15 13 2 16 10 9 2 0 7 0 2 15 13 1 10 0 9 2
43 10 9 3 0 2 3 0 7 0 16 10 9 13 3 13 1 9 0 1 10 11 2 10 10 9 15 13 10 10 9 2 12 9 3 13 1 10 9 1 9 1 11 2
3 11 2 11
7 11 13 11 1 13 9 2
31 10 11 13 13 3 10 9 1 9 1 10 0 9 2 1 13 10 9 1 9 7 13 10 9 1 9 13 1 10 9 2
55 10 9 13 3 13 1 10 9 1 10 11 2 1 10 10 3 0 9 1 10 9 1 10 9 0 2 1 15 15 13 10 9 1 10 9 1 13 10 9 1 10 11 1 10 9 1 13 2 3 2 10 9 0 0 2
35 10 9 13 16 10 11 13 12 9 1 12 2 1 12 9 10 9 2 3 10 9 13 1 12 9 1 12 1 12 9 1 10 0 9 2
43 10 11 13 16 1 10 12 0 9 10 9 9 13 10 0 9 2 7 13 10 9 1 10 9 0 7 0 9 1 10 9 2 16 10 9 1 9 3 13 1 4 13 2
28 1 15 15 15 13 2 10 9 1 10 0 9 1 10 9 13 3 13 2 16 10 9 3 3 13 4 13 2
31 3 15 2 10 9 1 10 11 13 4 1 13 15 7 1 4 15 1 10 9 13 1 10 9 1 10 9 1 10 11 2
41 13 10 9 1 10 9 1 10 11 1 10 11 7 1 10 11 2 15 13 4 1 13 10 10 9 1 13 10 9 3 13 0 10 10 9 1 9 1 10 9 2
26 1 11 2 9 0 1 10 11 2 10 9 1 11 1 10 11 13 2 10 9 1 10 9 0 2 2
35 13 2 10 9 13 10 9 1 16 2 3 13 13 10 9 1 13 1 10 9 1 10 9 15 3 13 13 3 10 9 1 10 9 2 2
38 10 9 1 10 9 1 11 13 2 3 2 13 3 13 13 10 9 1 10 9 7 2 3 2 13 2 15 13 10 9 1 10 9 1 10 9 2 2
49 1 10 9 1 10 11 2 13 10 11 2 10 9 1 10 9 1 10 11 13 9 1 10 10 9 2 16 15 13 3 13 1 10 11 2 10 9 0 2 1 10 0 11 2 15 3 15 13 2
27 2 13 12 9 1 9 1 10 9 2 10 0 7 15 0 2 2 13 11 2 9 1 9 1 10 11 2
12 2 3 2 13 0 3 1 10 9 0 2 2
60 13 1 10 9 3 13 1 10 9 2 10 9 11 2 13 1 10 9 1 10 11 2 13 2 1 10 9 1 12 1 12 2 3 13 10 9 1 10 9 1 10 9 3 13 10 9 1 9 1 10 9 2 13 1 10 9 7 10 9 2
42 1 9 1 10 11 7 1 15 11 2 10 12 9 0 13 1 10 9 2 2 15 13 10 9 13 1 10 11 2 13 0 1 10 9 10 9 1 9 1 10 11 2
40 3 2 1 10 12 9 13 15 10 9 2 10 9 0 2 10 9 2 10 0 2 10 9 7 10 9 3 15 1 10 9 7 15 1 10 9 2 1 10 2
23 12 1 11 2 10 11 13 1 9 1 10 9 2 13 13 1 10 9 0 1 10 11 2
38 12 1 11 2 10 11 13 1 10 9 1 10 11 2 1 10 9 1 10 9 0 1 12 9 7 10 9 1 10 0 9 1 10 9 1 12 9 2
1 11
22 11 13 9 1 10 9 2 15 1 15 13 13 1 3 12 9 7 13 10 9 0 2
11 13 10 0 9 1 10 9 2 11 2 2
1 11
16 11 1 10 11 2 1 10 9 1 10 9 0 1 10 9 2
9 9 0 1 10 11 13 13 12 9
9 11 3 13 7 13 9 1 10 9
34 12 9 1 10 9 0 1 10 9 1 10 11 2 13 0 10 9 1 10 11 2 10 9 0 1 10 11 13 1 13 10 10 9 2
19 10 9 13 3 0 1 10 9 15 3 1 10 11 15 13 3 1 15 2
23 13 3 1 3 13 15 13 1 13 10 9 2 15 15 13 7 15 15 13 13 1 13 2
14 10 9 13 3 1 10 9 1 15 13 1 10 9 2
9 1 10 9 10 9 13 10 9 2
43 10 9 15 13 1 15 13 11 2 9 1 10 9 0 7 1 10 0 9 0 7 0 2 1 11 2 9 1 10 9 0 7 9 1 16 10 9 13 1 13 1 11 2
23 7 15 3 13 16 10 9 1 1 11 7 10 9 0 13 3 3 3 0 7 3 0 2
26 10 11 13 16 1 13 10 9 1 12 9 1 9 0 2 13 0 10 9 1 12 9 1 12 9 2
37 10 9 2 13 13 10 0 0 9 1 9 0 7 0 1 10 9 1 10 9 1 13 13 3 1 10 9 1 10 9 0 2 2 13 10 9 2
17 10 0 9 2 1 12 12 9 2 13 3 13 1 10 10 9 2
5 9 13 1 10 11
34 10 11 13 3 11 1 13 1 10 0 9 10 9 1 10 11 1 15 13 9 1 13 10 9 1 11 2 1 10 9 1 10 9 2
68 2 1 16 13 3 13 1 10 9 0 2 10 9 0 13 16 10 9 0 13 10 9 1 11 1 16 13 10 9 7 1 16 15 13 1 9 0 2 13 10 10 9 2 2 13 10 11 2 9 15 13 1 10 9 1 10 9 1 10 11 2 1 10 9 13 1 11 2
62 10 9 11 13 13 1 10 10 9 11 2 0 11 2 1 10 0 1 12 2 12 2 2 12 2 15 13 16 10 9 12 1 10 9 13 13 1 10 2 9 1 10 9 13 2 2 11 2 1 12 9 1 10 10 9 13 1 10 9 1 9 2
28 11 2 9 12 1 10 2 9 2 2 13 13 1 10 9 11 2 0 11 2 1 10 0 1 12 2 12 2
24 0 13 3 10 9 1 10 9 1 10 9 1 11 2 1 10 9 13 2 10 13 1 9 2
36 11 2 9 1 10 9 0 2 13 13 1 11 1 12 2 12 2 7 11 2 9 1 9 9 2 13 13 1 11 1 12 2 12 7 12 2
39 3 15 13 15 13 3 3 10 9 1 10 9 3 13 4 13 2 11 13 16 13 2 13 13 1 10 9 2 13 3 10 9 3 10 9 15 13 2 2
19 2 16 15 13 13 2 13 4 13 3 3 13 1 10 9 2 2 13 2
10 2 10 9 3 13 16 15 13 9 2
7 3 15 13 13 3 9 2
44 13 15 16 10 9 13 13 1 10 9 2 15 13 13 10 9 1 10 9 1 15 13 2 2 13 10 9 2 13 16 13 3 13 10 9 13 16 10 9 13 9 1 15 2
10 2 11 2 13 9 1 9 1 10 11
7 11 7 11 13 1 10 9
43 1 10 9 0 7 1 10 9 2 10 9 0 2 0 7 0 1 10 11 1 11 3 13 13 3 1 10 11 7 1 10 11 2 12 1 10 12 9 15 13 1 11 2
29 15 13 10 9 1 15 13 10 9 1 9 2 11 2 2 15 13 1 10 10 9 1 9 10 9 1 10 9 2
42 1 10 9 1 10 9 2 13 15 9 1 10 11 2 7 13 10 9 3 1 10 2 9 2 1 10 9 2 15 13 11 3 3 10 9 2 13 10 10 9 0 2
16 15 3 2 10 9 15 13 1 10 2 9 2 13 3 13 2
2 10 9
34 3 9 1 10 0 2 10 0 9 3 15 13 1 10 9 0 7 13 3 13 1 10 0 9 0 2 15 3 13 9 1 0 9 2
26 10 9 7 10 9 1 9 0 13 2 1 0 2 10 9 1 9 1 10 9 0 2 15 15 13 2
20 12 9 1 10 9 1 11 2 10 9 13 13 15 10 9 0 1 10 9 2
7 9 0 13 9 1 9 2
50 10 9 13 2 11 2 13 3 10 9 1 10 9 1 10 11 9 7 1 10 10 9 2 15 13 1 10 11 2 7 13 13 15 16 3 13 13 10 9 1 10 11 2 13 3 1 11 10 11 2
45 10 9 13 16 10 9 3 13 7 15 15 13 3 1 9 13 1 10 9 0 1 13 16 10 9 13 1 10 9 10 9 11 2 12 9 2 7 10 10 9 11 2 12 9 2
14 10 12 9 13 13 12 9 1 10 11 1 10 11 2
26 1 13 10 11 2 10 9 11 13 10 9 2 11 2 1 13 10 11 1 10 9 0 1 10 9 2
28 10 9 15 13 9 1 10 11 1 2 10 9 1 9 2 15 10 9 2 11 2 13 1 2 3 0 2 2
81 10 9 13 1 12 2 9 1 15 10 11 1 10 11 2 3 1 10 11 2 13 1 10 9 11 2 13 1 10 11 10 9 1 15 15 13 1 13 10 9 0 1 9 1 1 10 9 1 12 12 9 7 1 13 1 12 9 10 9 1 10 9 0 1 10 9 2 3 9 1 10 9 1 10 9 0 1 11 7 11 2
5 9 1 9 1 11
29 10 11 13 3 10 10 9 1 10 9 1 10 11 7 1 10 11 2 1 10 9 2 1 10 11 1 10 9 2
32 10 9 13 1 10 9 1 11 2 9 2 2 11 2 9 2 2 11 2 9 2 2 11 2 9 2 7 11 2 9 2 2
35 10 9 13 13 2 1 10 9 1 10 9 11 2 10 9 11 1 11 2 3 10 2 11 2 7 10 9 2 11 2 2 10 1 11 2
8 1 11 13 15 3 10 11 2
30 1 10 9 1 10 11 13 2 1 10 9 2 10 11 1 10 11 2 15 13 13 1 11 2 11 2 11 7 11 2
10 10 9 13 13 1 10 9 1 11 2
6 1 10 9 1 10 9
60 3 2 10 0 9 1 13 1 10 9 1 9 0 9 2 1 9 7 9 1 11 2 12 1 10 3 0 9 0 2 13 1 10 9 11 7 11 2 7 10 9 1 10 9 1 11 2 11 2 1 10 9 1 11 2 15 13 9 0 2
18 10 9 0 13 1 10 9 0 7 3 0 1 10 9 1 10 11 2
25 7 3 1 10 9 2 10 3 12 9 15 15 13 1 10 11 13 1 10 0 9 13 1 11 2
21 1 10 0 9 2 10 0 9 0 13 1 10 9 13 13 10 9 1 10 9 2
27 10 9 0 2 7 0 9 1 9 13 2 13 1 13 10 0 7 0 9 0 2 3 1 10 0 9 2
33 3 1 11 2 1 10 0 9 1 10 9 2 7 1 12 9 1 10 9 1 11 15 2 1 9 2 13 10 0 9 1 9 2
16 1 13 2 11 13 3 10 9 7 10 9 15 15 13 13 2
5 10 9 15 13 2
6 10 9 15 15 13 2
19 10 11 13 10 9 1 10 9 2 16 13 13 1 10 11 2 1 12 2
38 10 11 2 1 12 9 1 11 2 13 1 10 9 7 13 3 12 9 2 10 15 13 3 2 7 12 9 2 15 15 13 10 0 9 1 10 11 2
45 1 10 9 2 10 9 1 11 13 13 15 1 13 13 2 1 10 9 2 10 0 9 0 1 10 9 1 9 2 12 9 0 2 1 12 2 9 1 15 15 13 1 10 11 2
20 10 9 1 10 11 13 15 1 9 9 1 12 9 1 10 9 1 10 9 2
43 10 9 0 1 9 13 1 12 9 2 9 15 15 13 1 10 9 0 1 9 0 13 1 10 11 2 1 9 2 15 13 1 10 11 10 9 0 1 12 9 1 9 2
31 10 9 1 9 2 15 13 1 12 9 1 9 2 13 1 10 9 10 9 9 1 12 9 1 9 2 13 1 10 11 2
50 10 9 0 1 10 9 1 10 11 13 13 2 1 9 2 3 7 1 9 2 15 13 10 9 1 9 1 9 2 9 0 7 9 2 13 1 10 9 1 9 2 2 1 13 1 9 1 10 11 2
29 10 9 13 12 9 2 2 13 10 9 13 1 10 9 2 10 9 7 10 9 1 10 9 13 1 10 9 2 2
2 9 0
7 9 1 10 11 13 9 0
34 11 2 9 0 2 13 10 9 1 10 9 1 10 9 1 10 11 1 16 13 10 10 9 1 9 1 10 9 0 2 3 1 9 2
18 10 11 0 13 3 1 10 9 2 13 13 1 10 11 2 11 2 2
33 10 9 1 10 11 7 10 11 13 3 13 1 10 9 13 1 10 2 11 2 2 1 11 2 1 10 0 0 11 7 13 9 2
36 10 11 13 10 9 1 10 9 11 16 10 9 0 1 10 9 1 9 13 1 12 9 7 13 0 1 12 1 9 1 10 9 1 10 9 2
13 10 11 13 13 1 12 9 1 10 9 1 9 2
16 10 9 1 10 9 13 1 13 9 1 10 9 12 1 9 2
2 11 13
40 10 0 9 1 9 1 10 11 2 11 2 13 13 1 10 11 1 10 9 0 1 9 2 1 10 9 1 10 9 0 1 10 9 1 12 9 1 10 9 2
51 1 10 9 2 10 11 2 9 2 2 1 11 2 13 13 10 9 0 1 12 9 1 10 9 2 1 12 9 1 10 11 2 0 2 2 1 10 9 0 11 2 7 12 9 1 10 11 2 0 2 2
29 11 2 10 9 1 12 9 2 15 13 3 10 9 1 12 7 12 2 13 1 10 9 1 10 9 1 12 9 2
4 9 1 10 11
7 13 9 1 10 2 11 2
4 11 7 11 3
25 11 2 9 0 9 1 9 2 13 3 10 12 9 15 13 13 10 9 1 10 11 1 10 11 2
8 10 9 11 7 11 13 3 2
47 10 11 2 0 2 1 10 11 2 1 10 11 2 13 10 9 15 10 9 13 1 10 9 0 2 1 12 9 2 13 15 10 11 2 1 12 2 10 11 7 10 11 2 10 1 12 2
18 1 10 9 0 2 1 9 10 2 10 9 13 7 13 15 13 0 2
19 13 1 10 9 2 13 13 7 13 10 9 15 15 13 9 13 12 9 2
14 3 13 13 12 2 1 10 0 15 13 1 10 9 2
21 13 1 10 10 9 1 9 2 13 3 13 1 10 9 1 10 10 9 1 9 2
21 3 15 15 13 2 16 3 15 13 16 13 13 15 1 2 10 9 1 10 9 2
21 3 13 0 1 2 1 10 9 1 12 9 2 13 13 13 15 13 1 10 11 2
10 7 13 16 10 10 9 13 10 9 2
3 11 2 11
30 13 15 16 10 9 1 10 11 7 13 10 0 9 2 7 13 15 10 9 0 2 7 13 13 3 1 10 9 0 2
7 11 13 13 10 0 9 2
22 11 13 10 10 0 9 1 10 0 9 2 1 10 9 1 10 10 9 1 10 11 2
47 0 2 1 10 9 1 12 9 1 9 13 2 1 10 9 1 9 0 2 10 10 9 11 13 12 9 1 10 0 9 12 2 1 10 9 1 10 11 3 13 3 9 1 10 9 0 2
56 10 9 1 9 13 3 1 9 2 1 10 9 1 11 7 11 2 11 13 13 2 1 13 1 10 9 1 9 0 1 10 9 1 10 9 1 10 9 1 10 12 2 11 2 9 3 0 1 10 9 2 1 11 2 11 2
22 10 9 13 1 9 1 10 12 9 2 13 15 3 1 10 12 9 7 13 0 9 2
25 12 9 0 13 10 9 0 1 10 9 1 9 2 3 13 1 9 1 10 9 0 2 13 9 2
22 10 9 11 1 10 11 13 12 9 2 3 10 11 2 1 11 2 13 15 12 9 2
26 10 11 2 1 10 9 2 13 1 10 12 9 2 3 12 9 2 1 11 2 15 13 1 9 0 2
41 11 2 1 9 1 10 9 13 15 1 9 2 1 10 9 11 1 13 15 1 10 12 9 2 3 12 9 1 10 9 7 3 1 10 9 0 1 10 12 9 2
26 2 1 10 10 9 10 9 13 3 0 2 2 13 10 2 9 2 2 15 13 13 10 9 3 0 2
23 9 13 16 10 9 1 10 11 13 13 1 10 9 1 11 7 11 0 1 10 9 9 2
26 1 10 10 9 1 9 0 2 15 15 13 0 9 2 3 1 10 10 9 1 9 2 13 10 0 2
36 10 3 3 12 9 1 9 15 13 1 10 9 1 10 9 13 13 1 10 9 1 9 1 12 9 1 9 2 3 2 10 9 1 12 9 2
28 1 10 9 3 13 0 10 9 1 10 9 13 10 15 3 13 10 0 9 1 9 2 1 10 9 1 9 2
20 10 2 9 1 10 9 2 13 2 1 11 2 10 9 3 0 1 10 9 2
25 1 10 9 13 15 2 3 2 0 13 1 10 9 1 10 9 2 1 9 1 13 15 3 0 2
20 12 1 10 9 13 10 0 9 1 10 0 9 15 13 10 9 1 10 9 2
39 10 9 13 1 12 7 13 1 16 10 9 9 13 1 10 10 12 9 1 10 10 9 1 9 0 7 12 9 1 10 9 13 16 13 1 9 13 1 9
7 11 13 2 12 2 10 11
2 0 3
35 10 9 2 1 12 2 1 10 11 1 10 11 13 0 2 3 3 13 0 16 15 15 15 13 3 1 10 11 15 13 1 13 1 9 2
29 15 13 2 15 13 10 9 0 2 3 3 1 10 9 13 1 10 10 9 13 13 9 1 9 2 0 7 9 2
13 10 9 1 10 9 13 15 1 10 9 2 0 2
5 9 13 1 10 9
14 11 2 15 3 0 1 10 9 7 11 13 1 9 0
49 15 13 0 13 1 10 11 2 1 9 1 9 7 9 2 9 2 9 0 2 9 2 9 2 9 2 9 7 9 0 2 3 13 9 0 10 9 1 11 2 2 10 3 0 1 10 9 2 2
27 10 12 9 13 13 1 10 9 2 7 3 1 9 1 10 9 0 2 3 10 3 0 1 10 0 9 2
70 1 15 15 13 9 1 10 9 2 0 13 1 0 3 0 13 1 0 2 2 10 9 13 16 10 9 1 10 9 1 10 9 13 3 13 2 16 2 10 9 1 9 1 10 9 13 3 2 13 1 10 9 1 10 9 13 10 9 1 11 3 0 1 15 1 10 9 0 2 2
13 3 2 10 9 13 10 12 9 13 1 10 9 2
53 10 9 0 9 1 10 9 13 15 1 10 9 1 9 1 12 9 1 9 2 15 13 3 12 9 16 15 13 1 10 9 0 1 10 9 1 12 2 7 15 15 13 3 1 10 9 1 10 9 0 1 11 2
28 3 9 1 10 9 13 13 15 1 10 9 0 7 2 1 10 9 2 3 12 9 13 4 13 1 10 9 2
29 10 9 0 0 1 9 0 2 1 10 9 2 13 15 1 12 9 1 9 3 1 10 9 0 3 3 13 9 2
1 11
5 9 13 9 1 9
36 10 9 13 2 3 1 10 9 2 12 9 1 9 1 10 9 1 0 9 1 11 2 13 10 9 1 12 9 2 15 3 13 10 9 0 2
10 9 2 9 1 10 9 2 9 3 2
13 9 0 0 2 13 3 2 1 10 9 1 10 9
31 1 12 7 12 1 9 13 1 11 2 10 9 11 2 11 12 1 10 11 2 9 1 9 2 1 15 11 13 3 9 2
26 10 11 13 1 12 1 3 12 9 7 3 13 1 1 10 12 9 7 0 2 1 9 1 12 9 2
15 13 10 9 1 9 3 0 1 10 9 7 12 1 10 0
22 2 7 10 10 9 13 3 0 3 10 10 9 15 13 10 9 1 10 9 15 13 2
30 10 9 3 13 1 9 13 10 11 2 10 11 7 2 3 10 11 2 3 10 0 9 13 1 11 2 11 7 11 2
52 9 15 13 1 16 10 11 13 3 0 1 10 9 0 13 1 10 9 2 3 3 10 9 1 9 1 10 11 13 10 9 0 1 15 15 13 12 1 10 9 0 1 0 9 1 10 9 1 10 10 9 2
68 10 9 2 3 2 15 3 13 1 13 1 10 9 10 9 11 2 13 15 2 9 2 2 13 15 16 11 13 2 1 0 9 2 10 9 1 10 11 1 10 9 0 2 2 13 15 1 11 1 15 13 16 10 9 15 10 9 13 1 10 9 13 0 1 13 10 9 2
16 10 9 13 15 2 13 15 2 3 2 16 15 15 13 0 2
8 2 15 13 3 9 1 15 2
17 15 3 13 10 9 13 10 9 1 9 2 15 13 3 10 9 2
21 13 1 10 9 1 10 10 9 2 11 13 13 10 9 2 1 9 1 10 9 2
10 2 10 9 3 3 13 3 0 2 2
39 2 6 9 2 13 15 10 9 2 16 15 13 3 9 1 15 7 15 3 3 13 1 9 3 1 10 10 9 2 2 13 2 0 2 10 9 1 9 2
38 1 10 9 0 2 10 2 9 2 1 10 11 1 10 9 1 10 9 13 13 1 10 9 13 1 10 9 2 1 9 0 1 10 11 7 10 11 2
26 2 13 10 9 1 13 13 10 9 7 2 3 2 10 10 9 1 16 10 9 13 13 3 3 13 2
40 3 2 10 9 13 1 13 16 10 9 13 16 4 13 3 2 3 13 1 13 16 10 9 13 16 15 13 2 7 1 13 10 9 0 2 2 13 10 9 2
42 11 13 16 2 3 1 10 9 0 2 10 9 7 10 9 1 10 9 1 10 9 13 13 2 1 9 1 10 11 2 1 1 10 9 1 10 9 7 9 1 12 2
65 2 10 9 1 10 11 7 1 10 11 2 1 10 9 1 10 11 2 3 13 4 1 13 10 9 1 13 0 9 1 9 1 10 9 2 2 13 10 9 2 15 13 16 1 13 9 3 13 4 13 10 9 1 10 9 1 9 1 10 9 1 11 7 11 2
27 2 10 0 9 1 3 13 10 9 1 9 13 1 16 2 3 2 15 13 10 9 2 2 13 10 9 2
4 11 13 1 13
6 10 0 9 1 10 11
18 10 11 13 3 1 11 10 10 0 9 1 10 9 0 2 1 12 2
28 3 13 1 10 9 1 10 11 2 11 13 1 13 10 0 9 1 10 9 2 7 2 3 2 1 10 0 2
16 3 0 13 10 11 2 15 13 1 13 10 9 1 10 9 2
18 7 2 1 10 9 1 12 9 2 10 9 1 11 13 10 10 9 2
6 9 0 1 10 9 0
8 11 13 9 1 9 1 10 11
44 10 9 13 1 10 9 13 1 10 10 9 16 15 13 1 10 9 1 10 9 3 13 4 13 1 10 9 1 9 1 10 11 10 9 0 1 10 9 13 1 9 1 9 2
46 11 13 0 1 10 9 1 10 9 1 10 9 15 1 15 15 13 13 3 10 9 1 1 15 13 4 3 13 7 2 1 10 11 13 2 13 3 13 1 13 10 9 1 10 11 2
31 1 10 9 1 3 2 10 9 1 10 9 0 3 13 10 9 1 10 9 3 13 13 10 9 1 10 9 15 15 13 2
40 13 3 16 2 15 13 3 1 13 2 7 2 1 15 2 13 1 10 9 1 3 13 9 13 1 9 3 16 13 13 2 0 9 15 13 4 1 13 2 2
26 7 13 10 9 1 16 10 0 9 13 3 10 9 1 9 2 13 10 9 1 10 9 1 12 9 2
7 1 11 10 9 13 0 2
33 16 10 11 13 10 9 1 16 13 10 9 1 9 13 1 13 3 16 10 9 1 10 0 9 0 13 13 1 10 0 9 0 2
21 3 2 11 13 16 10 9 13 1 10 9 0 13 0 1 10 9 1 10 0 2
51 1 13 10 9 2 13 16 3 13 3 10 9 1 10 9 13 1 2 10 9 3 2 1 10 9 0 2 9 15 15 13 13 16 10 9 1 12 5 1 10 9 13 1 11 13 2 1 15 2 9 2
26 1 10 15 2 13 11 2 10 11 13 1 15 0 2 13 2 7 13 1 13 0 10 9 0 2 2
10 10 9 13 2 3 2 13 3 12 2
38 10 11 13 1 15 13 3 10 9 0 2 1 10 9 0 2 3 16 1 10 9 1 11 3 13 10 9 0 1 10 9 0 15 13 3 1 13 2
4 3 3 13 2
7 3 13 3 1 10 9 2
2 3 2
24 10 13 9 2 1 10 9 1 10 9 2 13 15 1 10 9 1 10 11 7 1 10 9 2
20 9 3 9 3 16 10 11 2 10 9 0 3 0 7 13 1 10 10 9 2
19 3 10 11 1 10 11 13 13 1 13 2 10 0 9 1 9 1 9 2
18 3 1 10 9 1 2 1 10 0 9 2 13 1 10 9 15 0 2
35 10 9 0 13 10 11 1 10 10 9 1 13 9 0 2 3 10 11 2 15 13 10 9 1 12 9 2 7 10 11 2 1 0 9 2
50 10 9 13 2 10 11 13 10 9 1 10 9 3 1 10 2 11 2 2 13 10 9 0 9 2 13 13 16 10 11 13 9 11 1 10 9 1 11 2 1 10 9 1 10 11 2 1 10 9 2
5 11 13 10 9 2
22 1 10 11 7 1 10 11 13 13 10 9 1 13 2 7 1 3 13 2 9 0 2
29 15 15 13 1 13 2 1 10 9 1 12 2 10 9 1 9 0 1 9 0 2 11 2 1 10 9 0 2 2
36 11 2 10 0 2 13 10 9 1 16 10 2 9 13 2 7 16 2 10 2 9 2 0 13 15 15 13 13 9 2 9 7 9 0 2 2
36 3 0 1 10 9 9 2 9 13 10 9 0 11 2 15 13 10 9 1 10 9 0 2 3 10 9 13 12 9 3 16 10 9 1 9 2
52 10 3 9 1 10 11 13 16 15 13 1 13 1 10 9 1 16 2 10 9 13 13 1 10 9 1 10 9 2 2 7 13 16 2 10 9 1 13 0 2 3 13 13 0 1 9 1 10 10 9 2 2
45 1 9 1 10 9 1 10 10 9 7 1 13 1 10 9 10 9 2 13 2 2 10 9 1 10 9 13 4 13 2 1 2 3 2 13 1 10 0 9 1 10 9 1 11 2
43 11 13 16 10 9 1 10 9 0 13 13 0 3 13 1 10 9 0 2 7 3 13 4 13 10 10 9 1 9 15 15 13 2 2 10 9 0 7 10 9 0 2 2
56 3 2 10 11 13 15 13 1 13 9 1 9 1 9 1 9 1 15 13 1 10 9 1 10 9 1 12 9 1 10 9 2 12 9 2 1 10 9 3 0 7 1 10 0 9 15 13 10 0 9 1 15 1 10 9 2
4 7 3 13 2
19 13 12 9 3 13 3 7 15 2 1 13 0 2 13 1 13 1 9 2
32 3 2 13 3 1 10 0 9 1 10 9 1 10 11 2 1 10 9 1 2 1 10 9 2 3 15 13 13 3 12 9 2
16 2 2 2 3 1 10 9 2 15 10 9 1 10 0 9 2
18 3 15 13 1 13 10 11 3 10 13 9 15 13 10 9 1 9 2
12 13 10 13 9 1 13 10 9 1 10 9 2
52 10 0 1 10 9 1 9 1 10 9 2 1 10 11 2 3 13 2 3 2 1 10 11 2 12 9 0 2 12 9 2 12 9 1 9 7 12 9 1 10 2 3 10 2 9 15 3 13 10 0 9 2
34 3 2 16 13 10 9 2 1 9 7 1 9 2 3 2 2 3 13 13 13 3 16 2 1 10 9 2 15 13 10 2 9 2 2
67 13 1 10 9 1 10 9 0 2 10 9 0 2 3 1 10 10 9 2 11 2 13 10 11 1 10 9 1 13 10 9 1 11 1 10 10 9 15 13 10 9 7 15 15 13 1 10 9 1 10 11 13 1 10 11 2 15 3 13 1 10 9 1 10 9 0 2
32 11 2 9 2 13 16 2 3 2 10 9 1 10 9 2 13 4 13 1 10 0 9 1 10 11 2 1 13 1 9 2 2
44 10 9 1 12 9 2 11 2 15 15 13 1 13 9 1 10 9 0 13 1 10 9 1 10 10 9 1 11 2 15 13 3 1 9 0 1 9 2 13 15 1 10 9 2
32 10 9 1 9 1 10 11 13 0 1 15 1 11 2 13 9 15 13 10 9 0 13 1 10 9 3 9 1 10 9 13 2
8 10 11 13 2 3 2 10 9
51 10 9 1 9 7 1 10 9 1 9 3 0 1 9 2 13 1 13 10 9 1 10 9 0 2 13 1 13 10 9 1 10 10 9 1 9 1 10 9 2 13 10 9 13 1 10 11 2 11 2 2
31 1 1 10 9 12 2 10 9 1 10 9 13 1 10 9 13 3 0 7 2 1 9 1 15 2 13 0 13 15 3 2
39 10 0 9 1 10 9 13 2 3 2 3 10 9 0 7 10 0 9 1 10 9 13 15 1 10 9 0 0 7 13 15 1 10 9 7 1 10 9 2
27 3 3 3 15 13 10 0 9 1 10 9 0 7 10 0 9 1 10 9 1 10 9 13 1 10 9 2
65 3 3 13 10 9 7 10 9 3 0 3 10 9 13 1 13 10 9 3 3 2 13 15 3 1 1 10 9 0 2 13 10 9 1 9 1 9 0 1 10 9 3 0 2 1 10 9 1 10 9 2 15 13 9 1 10 9 1 10 9 1 9 13 9 2
4 10 9 3 0
10 9 1 10 11 13 1 10 9 1 11
15 11 13 15 1 11 2 15 1 10 9 2 3 0 2 2
13 11 7 11 13 9 0 1 10 9 1 10 9 2
15 13 3 3 10 9 1 10 11 13 15 6 13 1 13 2
15 0 13 16 11 13 1 10 9 10 9 0 2 1 9 2
15 0 13 10 9 1 10 9 1 11 7 10 9 1 11 2
39 10 9 1 10 9 0 2 11 2 1 10 9 0 2 11 2 13 16 3 13 2 10 9 0 2 1 13 10 9 1 11 3 9 1 10 9 3 13 2
35 10 10 11 13 2 0 2 10 9 1 11 7 10 9 0 1 15 15 13 3 10 9 0 3 13 15 3 0 1 13 13 10 10 9 2
90 1 10 9 13 1 13 10 9 1 10 9 2 10 0 9 13 15 1 10 10 12 9 1 10 9 1 10 9 0 2 10 9 15 13 3 10 9 2 2 1 15 13 10 2 9 1 9 2 1 10 9 15 13 13 1 10 0 9 1 10 11 7 10 2 0 9 0 9 2 15 13 10 9 1 10 9 1 10 15 13 1 10 0 9 7 15 15 13 3 2
60 13 1 10 9 1 10 9 2 1 10 9 13 1 10 9 11 2 11 13 16 2 10 9 0 3 13 3 10 9 1 9 7 1 9 2 1 13 1 2 9 0 2 2 7 13 13 3 3 10 9 0 2 15 13 10 9 7 10 9 2
20 7 3 13 1 13 1 10 9 1 2 10 0 9 3 13 0 1 9 2 2
25 15 13 15 1 10 0 9 0 1 10 11 13 3 1 10 11 0 2 11 2 1 10 9 0 2
19 9 0 13 16 9 1 10 9 1 10 0 9 3 13 1 13 11 0 2
7 9 1 11 1 9 1 9
43 10 11 1 11 13 10 9 10 9 1 12 9 2 0 2 13 2 0 1 10 9 1 11 2 13 1 13 4 7 4 13 10 9 1 12 9 2 0 1 10 10 9 2
31 10 13 9 13 13 1 10 9 2 3 1 10 9 13 13 10 9 1 10 9 0 3 15 13 1 10 11 1 13 9 2
34 10 9 2 1 10 9 13 2 13 1 10 9 1 10 9 2 1 10 9 0 2 1 10 9 0 2 10 9 3 13 1 10 9 2
30 1 10 9 1 15 13 1 9 2 10 9 13 15 1 15 2 13 15 10 9 2 13 15 7 13 15 1 10 9 2
11 3 13 15 10 9 7 13 13 10 9 2
33 10 9 13 9 7 2 10 9 3 3 2 13 10 9 1 10 9 2 1 12 9 2 15 13 1 10 9 7 13 10 13 9 2
1 11
6 9 13 9 1 10 11
14 1 10 11 2 1 11 2 13 13 10 9 1 9 2
41 1 10 9 0 13 13 10 9 1 9 1 9 7 9 1 0 0 2 10 0 1 15 13 9 1 10 9 1 9 13 7 13 1 9 1 10 9 1 10 9 2
27 1 13 10 9 2 10 9 1 10 9 1 9 0 13 3 13 1 10 9 7 10 9 1 10 11 0 2
2 0 9
4 9 2 9 0
18 9 0 7 9 0 13 10 9 0 1 10 0 9 1 10 9 0 2
21 15 1 10 10 9 0 7 1 10 9 1 10 9 1 10 9 1 9 1 9 2
2 0 9
16 3 12 9 15 13 3 2 3 10 9 0 13 1 10 11 2
28 1 10 9 0 13 1 13 9 1 10 9 2 10 9 13 1 11 13 1 13 15 1 10 9 0 7 13 2
15 1 10 9 15 13 10 9 1 9 13 10 9 3 0 2
17 10 9 11 13 1 10 12 9 2 3 12 9 1 10 9 0 2
24 10 9 13 3 10 9 1 10 9 1 10 9 1 2 11 2 2 13 0 9 1 10 9 2
16 13 2 3 2 0 16 3 3 10 12 9 13 13 3 13 2
52 3 2 13 10 9 0 2 2 10 9 0 13 1 10 9 0 1 10 9 1 9 0 2 1 10 9 1 0 9 2 1 10 9 1 9 15 13 10 9 0 7 2 1 10 9 2 13 3 10 10 9 2
86 3 2 3 2 15 3 13 10 9 1 10 9 2 13 10 9 1 10 9 1 11 2 9 2 3 2 10 9 1 11 2 2 15 2 3 2 13 1 16 10 11 13 1 13 9 1 13 2 1 10 10 9 0 1 9 2 10 9 1 10 10 9 7 13 10 10 9 2 9 2 9 7 9 2 15 3 3 3 13 13 1 13 1 10 9 2
90 10 9 1 13 9 1 10 9 1 10 11 13 13 1 10 9 0 1 10 9 9 2 9 1 10 9 1 10 9 0 2 1 10 9 1 10 9 1 10 0 2 15 13 1 13 0 9 1 10 9 13 1 10 0 1 13 1 13 0 1 10 9 13 15 13 10 9 2 3 0 2 15 13 10 9 0 2 11 7 11 2 7 13 10 9 0 1 10 9 2
51 3 2 10 9 1 10 9 1 10 9 7 10 9 1 9 0 13 9 0 1 10 10 9 1 10 9 1 13 2 13 3 1 13 10 9 0 1 10 9 7 2 3 2 1 10 9 0 1 10 9 2
26 1 10 9 1 10 9 2 9 1 10 9 2 15 13 10 9 2 13 7 13 13 15 15 15 13 2
24 3 11 13 3 13 3 0 1 10 9 2 13 10 9 3 0 1 10 9 15 15 13 13 2
22 7 10 9 13 16 3 1 11 3 10 9 0 13 10 0 9 7 9 1 10 9 2
11 3 13 1 10 9 10 9 3 13 13 2
11 13 3 13 9 0 1 10 9 0 13 2
22 10 0 1 10 9 13 10 0 1 12 9 2 9 1 10 11 1 11 7 9 3 2
21 13 1 10 9 0 2 7 10 10 9 13 3 10 9 2 10 9 2 10 9 2
7 2 15 13 1 10 9 2
20 3 1 10 9 1 9 2 13 16 13 10 10 9 1 15 2 2 13 11 2
18 3 3 13 15 1 10 9 1 9 7 3 13 15 13 2 9 2 2
11 13 1 13 2 13 9 2 13 10 9 2
10 10 2 9 2 0 15 13 13 9 2
50 1 10 0 9 2 10 9 3 13 13 2 9 1 10 9 2 16 2 3 12 9 1 9 0 15 13 2 10 9 3 13 2 2 13 11 2 15 13 13 10 9 1 10 9 12 2 0 15 13 2
31 3 2 1 10 9 1 10 9 2 11 7 11 2 3 1 9 1 10 9 2 13 1 13 9 1 10 9 11 7 11 2
39 3 2 11 13 12 1 10 9 0 1 10 9 1 10 9 2 15 15 13 13 12 1 10 0 0 1 10 9 0 15 10 10 9 13 1 10 9 0 2
6 13 10 9 3 13 2
36 11 13 15 3 2 3 13 2 1 10 9 1 15 13 0 10 11 1 10 11 2 11 2 7 13 10 9 1 2 3 13 10 10 9 2 2
38 13 13 13 9 1 10 9 3 1 10 11 2 11 13 16 2 10 9 13 16 4 13 1 10 11 15 13 10 9 1 10 9 7 13 10 9 2 2
13 1 15 13 9 1 10 9 2 13 1 10 9 2
12 2 15 13 10 9 1 9 3 13 15 2 2
47 11 13 10 11 1 13 10 9 2 0 7 0 2 1 10 9 2 2 13 9 1 9 1 9 10 15 13 13 1 10 11 1 10 9 1 9 0 1 10 9 1 10 0 9 0 2 2
27 11 3 13 13 10 2 9 2 1 10 9 7 13 13 10 9 0 1 10 11 0 2 1 9 1 9 2
4 9 1 10 9
31 10 9 1 10 9 1 9 1 13 1 10 9 13 10 9 2 1 10 13 9 2 1 10 11 2 11 2 1 10 11 2
33 12 1 10 9 13 1 10 11 13 10 9 1 10 9 1 10 11 1 10 9 1 9 7 1 10 9 1 10 9 0 7 0 2
54 12 9 15 2 1 15 13 1 10 9 0 2 2 3 13 1 0 2 7 13 13 10 9 1 12 15 13 10 9 1 10 9 2 13 15 3 0 9 7 9 1 10 9 1 10 9 1 10 9 0 1 10 9 2
42 10 2 9 1 9 1 10 9 1 10 9 1 10 9 2 1 13 1 10 9 13 15 1 10 9 1 10 11 2 15 13 10 9 0 2 2 13 1 9 0 2 2
21 13 2 1 15 2 16 2 10 9 1 9 1 9 13 1 4 13 1 9 2 2
56 10 9 1 10 9 0 13 16 10 9 3 0 9 13 9 0 1 10 9 1 10 9 9 1 10 9 2 16 10 9 1 9 0 1 10 9 13 10 9 1 10 9 7 16 10 9 13 13 1 10 9 1 9 1 9 2
29 10 2 9 1 10 9 2 13 9 0 1 10 9 1 10 9 7 13 11 1 13 1 10 9 7 1 13 11 2
47 7 10 9 1 10 9 1 10 10 9 1 9 7 2 3 2 10 0 9 1 10 9 0 2 13 1 16 10 9 13 3 15 15 13 13 2 3 13 13 11 1 10 9 1 10 11 2
5 11 13 1 10 9
2 1 9
6 11 2 10 9 1 11
23 10 11 13 10 0 9 1 10 11 2 3 1 15 1 15 15 13 13 2 10 9 2 2
28 13 10 9 13 11 2 13 1 15 2 7 15 3 13 13 10 9 1 10 9 1 10 9 1 10 9 0 2
5 2 10 9 0 2
37 10 9 1 11 2 11 2 13 1 10 9 1 10 11 1 12 1 9 1 10 9 1 9 13 3 0 1 15 15 13 1 10 9 1 10 9 2
15 13 2 3 2 10 9 15 3 13 13 1 10 10 9 2
32 13 16 13 1 10 9 0 1 15 13 1 9 3 0 1 9 2 3 13 10 9 1 9 13 1 2 9 2 2 1 12 2
26 3 2 16 10 9 13 2 7 13 2 0 2 16 13 9 3 0 15 3 13 13 2 7 3 2 2
35 3 2 13 15 10 0 9 1 9 1 10 10 9 1 9 0 2 3 0 2 1 13 3 1 10 9 1 10 9 7 1 10 0 9 2
14 13 15 10 10 9 15 13 1 3 0 3 0 9 2
28 7 2 16 10 9 13 13 10 9 2 13 10 9 2 13 0 16 10 9 13 1 10 9 2 15 3 13 2
103 3 2 13 1 10 0 9 1 10 10 9 2 15 3 13 2 13 16 13 2 3 2 10 9 0 2 1 9 0 2 0 2 3 2 2 1 10 9 1 10 3 0 2 3 1 10 9 0 2 9 1 9 1 9 1 10 11 2 10 9 0 3 13 3 9 1 15 2 1 10 11 1 10 11 2 2 7 1 10 9 1 10 9 1 10 9 0 1 10 9 0 1 10 10 9 3 9 0 2 0 7 0 2
53 1 10 9 2 13 13 10 9 1 13 10 9 7 13 13 10 9 1 10 0 9 7 1 10 0 9 7 2 3 2 1 13 10 9 1 10 10 9 1 10 9 0 1 10 9 2 13 15 1 10 9 0 2
24 1 10 9 2 11 2 2 3 1 10 11 2 13 1 13 1 10 9 1 15 1 13 15 2
65 13 1 15 13 10 9 0 1 10 0 9 2 13 7 1 0 2 1 10 9 1 10 9 1 10 11 2 13 12 9 2 2 2 1 9 3 13 7 3 13 3 11 2 15 3 13 1 10 9 2 7 1 10 15 15 13 10 9 0 2 0 7 0 0 2
61 13 15 16 13 3 10 0 9 1 0 9 2 10 0 2 1 10 9 0 1 10 0 11 13 9 0 1 10 11 2 15 3 13 1 10 9 0 2 1 10 9 15 13 13 3 1 10 9 1 10 9 1 10 12 9 16 10 15 3 13 2
12 10 9 1 9 1 9 13 3 15 13 13 2
19 13 15 2 3 2 3 13 0 1 10 9 10 9 1 9 1 10 11 2
22 3 2 10 9 0 13 13 3 0 1 15 15 15 13 1 10 11 16 10 9 0 2
21 1 10 9 2 3 10 9 0 13 1 13 10 9 1 10 9 2 1 9 0 2
42 1 10 9 2 13 13 10 9 1 10 0 2 3 1 15 3 2 13 2 10 0 9 1 10 9 1 9 2 2 1 3 1 10 9 10 9 13 1 13 10 9 2
45 0 1 10 10 2 9 2 1 11 2 13 10 9 2 7 3 13 10 9 1 15 1 12 9 2 1 12 13 12 9 2 3 13 15 1 15 12 2 13 9 1 9 7 9 2
28 10 0 1 10 9 3 13 13 1 10 0 9 0 2 15 10 9 13 3 15 13 13 1 10 9 1 9 2
52 1 13 10 9 11 2 10 9 3 1 10 0 9 13 1 15 2 0 9 2 0 1 9 0 2 2 3 13 10 9 1 10 9 15 2 3 1 13 1 10 9 2 13 1 13 3 16 3 1 10 9 2
45 1 9 0 2 10 9 13 3 13 9 1 10 2 0 9 2 15 1 15 15 13 7 15 1 10 9 1 10 9 13 2 3 3 9 13 1 9 16 3 9 1 9 0 2 2
35 10 9 1 13 1 10 9 1 10 11 13 15 15 13 9 1 10 9 1 9 2 1 10 9 1 10 11 7 1 10 9 1 9 0 2
44 1 10 0 2 10 9 1 10 9 1 10 9 13 10 9 1 10 9 15 13 1 16 2 1 10 9 2 13 11 2 3 12 0 1 10 9 13 13 13 1 13 0 9 2
19 9 2 13 2 3 2 2 9 1 9 1 9 7 9 1 10 9 2 2
25 15 15 10 11 13 13 2 10 9 1 9 1 10 9 1 0 9 2 1 15 13 10 9 2 2
6 10 9 13 13 4 13
1 11
2 12 9
1 0
2 9 2
9 1 3 9 13 13 9 1 11 2
5 13 10 9 13 2
10 9 2 13 10 9 2 10 9 3 2
9 3 13 3 0 1 10 10 9 2
19 13 16 10 9 0 15 13 16 3 13 13 2 7 13 2 7 13 13 2
22 7 3 13 9 2 1 15 13 2 1 10 9 0 1 10 9 0 2 13 15 3 2
41 13 16 10 9 15 10 9 13 16 13 1 10 9 2 1 10 9 7 10 10 9 1 10 9 13 15 1 13 1 10 9 7 3 1 13 7 3 13 10 9 2
14 9 2 3 16 13 13 2 3 15 13 1 10 9 2
9 3 3 2 10 9 0 13 0 2
42 1 13 0 2 11 7 10 10 9 13 3 0 9 1 10 9 2 3 1 10 10 0 9 0 1 10 9 2 16 3 3 1 10 9 15 13 13 15 0 7 13 2
48 10 0 2 7 3 2 13 2 2 9 13 13 1 10 9 1 10 9 2 11 2 11 2 11 2 7 10 9 0 0 13 3 3 0 9 1 10 0 9 0 1 10 11 2 13 1 9 2
51 1 13 16 13 10 9 0 1 10 10 0 9 1 2 9 1 10 9 2 1 10 11 2 1 10 9 1 10 11 13 1 11 2 11 2 11 13 16 15 10 7 10 10 9 1 10 11 13 13 3 2
54 1 10 9 2 10 3 0 13 15 1 16 13 13 10 9 0 1 10 11 2 16 3 13 13 3 2 7 3 16 3 13 1 10 9 2 7 3 13 10 0 9 16 9 0 13 13 1 10 9 1 0 9 0 2
26 2 13 13 10 9 1 1 10 9 1 10 11 2 2 13 11 1 10 9 1 11 2 1 10 11 2
4 7 13 3 2
14 2 16 13 3 2 10 9 13 3 10 9 0 2 2
9 7 1 15 13 15 2 13 3 2
8 2 15 3 15 13 1 3 2
29 13 1 1 10 11 2 1 10 11 7 1 10 9 1 10 11 2 1 15 13 2 7 13 9 7 9 0 2 2
2 11 2
51 1 10 9 2 10 0 9 1 10 10 9 13 10 9 1 0 9 2 10 9 1 9 1 9 1 9 7 9 2 10 9 1 10 9 1 9 15 13 13 0 9 1 10 9 1 9 0 7 0 0 2
14 11 13 16 11 13 0 1 13 9 7 1 13 9 2
24 2 12 9 2 10 11 2 10 11 7 10 10 9 13 1 9 7 13 1 10 9 1 11 2
19 10 11 13 13 16 15 13 10 9 3 2 1 9 2 13 13 10 9 2
12 1 10 9 2 10 10 9 3 13 1 13 2
10 13 10 9 7 13 15 10 0 9 2
21 10 10 9 13 7 13 3 1 10 10 0 9 2 2 13 10 9 2 2 2 2
21 10 10 9 13 1 10 9 1 13 3 1 13 16 10 9 15 13 11 7 11 2
14 16 3 13 12 9 1 9 2 13 7 13 1 9 2
22 2 13 10 0 9 0 7 13 0 1 13 10 9 1 10 9 1 10 3 13 9 2
13 13 10 9 0 13 1 10 11 2 3 9 2 2
14 13 0 1 10 0 9 1 10 9 2 1 10 11 2
13 13 12 9 2 13 13 3 13 2 1 10 0 2
13 3 2 13 15 9 1 9 1 10 3 0 9 2
21 7 13 16 13 3 1 13 1 10 0 9 2 1 10 9 0 7 1 0 9 2
43 1 10 0 9 2 1 10 9 1 10 9 1 10 9 0 13 1 10 9 2 10 9 1 10 0 9 13 3 9 0 2 15 13 1 12 9 10 9 13 1 10 9 2
35 1 10 9 1 11 2 11 2 11 7 11 10 9 13 10 9 1 9 0 7 3 1 9 1 13 16 10 9 3 13 9 1 10 9 2
42 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 7 11 13 10 0 13 1 11 2
16 13 3 2 1 15 13 1 10 9 2 11 2 11 7 11 2
63 10 9 13 13 1 10 9 0 1 11 2 10 9 1 9 2 13 1 10 9 1 10 9 0 1 10 9 2 1 10 0 9 1 9 1 13 1 9 2 9 7 9 2 13 1 10 9 2 1 10 9 7 1 10 9 1 9 1 12 0 9 0 2
50 2 3 13 9 16 13 10 9 1 15 7 16 13 13 2 2 13 12 1 10 9 1 10 9 2 10 9 11 2 9 1 10 2 11 2 7 10 9 15 3 13 10 9 1 10 9 1 10 11 2
26 11 13 3 1 10 9 0 2 9 1 10 9 2 7 13 0 13 1 9 3 0 1 10 10 9 2
26 10 9 13 0 7 10 11 2 16 1 10 0 9 1 9 10 0 13 3 13 15 2 13 10 9 2
80 1 10 13 9 2 10 11 13 1 10 11 2 1 9 0 2 10 9 1 9 1 10 9 1 9 2 7 3 1 9 2 11 2 1 10 11 2 13 1 10 9 10 9 1 10 9 2 9 15 10 9 13 1 2 9 0 2 2 13 16 10 9 13 1 10 9 1 10 9 7 3 13 1 4 13 2 15 3 13 2
46 3 2 10 11 13 1 13 1 10 9 2 1 10 9 1 11 2 15 13 15 13 1 10 9 1 10 2 9 1 10 9 15 13 7 13 1 10 11 7 1 10 9 1 11 2 2
59 11 13 16 10 11 13 10 9 1 10 9 1 11 1 0 9 1 9 0 7 2 13 3 12 1 10 0 9 0 1 10 9 2 1 10 9 1 15 13 1 12 1 10 0 9 0 1 10 9 2 2 13 1 10 9 0 7 0 2
42 10 9 0 1 10 11 13 15 3 1 10 9 0 1 10 11 1 13 10 2 9 2 1 10 9 7 1 10 11 15 13 1 10 9 0 1 10 9 1 10 9 2
24 10 9 1 10 9 1 10 11 2 10 9 0 2 13 12 1 10 9 1 9 1 10 9 2
34 10 9 1 10 9 2 1 11 7 11 2 1 9 1 9 0 0 3 15 13 3 1 9 1 10 9 1 10 9 0 1 10 11 2
4 2 7 11 3
11 10 11 2 11 13 3 15 1 10 9 2
37 15 13 13 3 1 10 9 1 10 9 1 10 11 2 3 1 10 11 13 12 9 1 10 11 1 3 13 1 10 9 0 1 10 2 0 2 2
20 13 0 16 10 9 13 10 13 15 2 16 9 7 9 13 7 9 13 9 2
11 1 10 9 2 10 11 13 1 10 9 2
39 10 9 1 10 9 13 3 3 13 2 1 12 9 1 9 1 13 1 10 9 1 12 9 7 1 13 0 13 1 10 2 9 2 1 13 15 15 13 2
2 9 12
9 13 10 0 9 2 1 12 9 2
19 3 11 7 11 13 10 12 0 9 2 7 10 11 3 13 1 10 9 2
27 10 11 2 11 1 3 3 13 1 13 9 2 7 13 13 10 11 2 11 1 12 1 9 15 15 13 2
27 16 10 11 13 3 10 11 7 10 11 13 10 11 2 13 11 7 11 3 1 15 9 1 10 11 13 2
2 9 12
85 10 9 0 1 10 9 2 13 1 10 11 2 13 10 9 1 10 9 0 1 9 1 10 9 2 1 12 9 0 2 9 1 10 9 0 2 9 0 1 10 9 1 10 9 7 9 1 10 9 1 9 13 2 9 1 9 1 9 13 10 9 9 7 0 7 9 1 10 9 1 10 9 2 1 13 16 15 15 13 9 7 9 1 9 2
14 2 10 9 9 13 4 13 13 10 9 1 10 9 2
13 3 13 10 9 7 10 9 15 13 10 9 2 2
12 10 0 9 13 15 13 10 9 0 7 0 2
18 10 11 3 13 2 1 10 9 2 1 12 9 9 7 12 9 9 2
15 2 10 9 13 4 13 9 1 10 10 9 13 9 2 2
3 9 7 9
6 11 13 1 10 9 2
38 15 3 13 10 9 13 10 9 1 10 11 2 0 1 13 16 10 9 1 10 9 1 9 1 11 13 1 10 0 1 10 9 2 13 10 9 11 2
11 10 9 1 11 13 16 10 9 3 13 2
47 1 10 9 12 1 9 10 9 1 10 9 13 16 3 13 10 9 1 11 1 10 9 1 13 10 9 1 10 9 7 13 15 0 1 10 9 0 2 3 1 15 13 1 10 9 0 2
18 1 3 2 15 13 2 1 10 9 1 11 2 10 9 1 10 9 2
31 13 15 10 9 7 1 15 13 16 11 13 13 10 9 1 10 10 9 2 1 13 1 10 0 9 1 10 2 11 2 2
32 13 10 9 2 13 15 1 10 9 0 1 3 2 16 11 2 13 16 10 9 3 13 1 10 9 1 9 1 10 9 2 2
15 1 13 1 10 9 2 13 10 9 2 2 10 9 2 2
12 13 3 10 9 1 10 11 2 13 1 9 2
21 11 2 13 15 1 10 9 7 13 1 9 2 13 10 2 11 2 1 10 9 2
15 7 3 13 10 15 15 13 13 3 10 11 7 15 13 2
15 9 2 1 9 1 9 2 9 1 9 2 9 1 9 2
7 9 2 13 10 9 10 2
34 9 2 13 10 9 1 13 9 1 10 15 13 13 2 7 13 16 13 13 2 16 3 10 9 3 13 3 1 10 9 1 10 9 2
12 10 11 13 13 10 9 0 1 10 10 9 2
17 3 13 10 9 1 10 9 1 11 2 13 10 9 1 9 0 2
24 3 15 13 10 9 0 2 13 10 9 1 10 11 2 11 2 2 16 3 13 1 10 9 2
17 3 3 10 11 3 13 7 13 10 9 3 13 13 10 9 0 2
14 1 15 2 16 15 13 13 2 13 15 1 10 11 2
33 3 10 9 13 2 10 9 0 13 1 15 9 9 1 10 2 9 3 2 1 10 9 13 1 10 9 1 10 9 0 1 11 2
41 10 9 0 2 1 10 9 0 2 10 9 0 9 13 9 0 7 1 10 9 1 13 13 1 10 9 2 13 3 1 10 9 1 10 9 2 7 13 10 9 2
35 3 2 10 9 0 7 13 13 3 13 9 1 10 9 2 7 3 1 9 0 2 0 7 0 2 13 1 9 0 7 13 1 10 9 2
36 3 2 10 2 9 1 10 9 13 1 12 2 3 13 10 9 1 10 9 7 1 10 0 9 13 1 4 13 15 3 13 13 10 9 0 2
13 2 13 1 9 1 9 2 9 1 10 9 0 2
14 13 10 9 1 10 9 1 10 10 9 1 10 9 2
55 13 3 12 9 2 7 15 13 12 2 2 13 3 2 1 10 9 1 10 2 11 2 2 11 2 9 1 12 1 10 12 9 1 0 1 11 2 15 13 3 12 9 13 1 13 4 13 2 13 7 13 1 10 9 2
42 12 1 10 9 1 10 11 2 3 15 13 13 12 9 11 2 9 1 10 11 2 13 13 10 9 1 10 9 0 1 10 9 0 2 1 15 13 13 1 9 0 2
27 3 2 1 10 9 0 1 9 7 2 1 10 15 2 1 10 9 1 10 9 3 1 10 0 9 0 2
34 10 11 13 15 13 1 10 0 9 2 13 10 9 7 13 10 9 0 2 1 10 9 1 15 13 1 10 9 1 15 14 7 9 2
13 11 3 13 10 9 0 2 7 13 10 9 0 2
21 2 10 9 0 2 1 10 11 2 13 13 10 9 2 13 15 1 10 9 0 2
19 7 10 9 1 10 10 9 3 15 13 1 10 9 1 10 9 0 0 2
10 3 13 10 9 0 2 1 9 2 2
27 10 9 13 10 9 1 13 15 15 13 7 3 13 16 13 0 13 15 1 10 9 16 13 10 0 2 2
5 10 9 1 10 9
39 11 2 1 12 2 13 3 13 13 2 2 13 13 2 3 2 16 10 9 13 9 1 9 2 9 13 3 1 10 9 1 10 11 1 10 9 1 11 2
11 1 16 13 13 3 0 3 3 13 9 2
58 10 9 1 12 9 13 10 0 1 13 1 10 9 0 16 2 3 1 9 2 13 13 9 1 10 11 2 1 12 7 12 1 10 9 13 2 9 15 13 9 1 10 9 1 12 9 1 10 11 1 11 7 10 9 1 10 11 2
32 10 9 2 13 15 2 13 1 9 1 10 9 13 2 3 3 1 10 9 1 10 11 7 13 1 10 9 1 9 3 13 2
68 1 9 1 10 0 9 1 10 9 2 10 11 2 11 13 12 1 10 2 9 2 2 9 2 1 11 2 15 13 3 1 10 9 1 10 11 2 11 2 7 13 0 16 10 9 13 0 9 2 13 2 3 2 16 10 9 2 7 3 3 1 12 9 2 13 3 0 2
30 2 1 10 9 13 10 9 2 1 9 1 10 2 0 1 15 2 2 11 1 10 12 9 1 10 2 11 2 2 2
61 2 2 10 9 1 10 11 7 1 10 11 3 3 13 13 10 9 0 1 10 9 1 10 9 1 10 10 2 14 2 9 2 11 2 2 15 13 4 4 3 9 0 1 10 9 1 9 0 7 4 13 3 2 2 2 11 2 2 9 2 2
37 3 1 10 0 0 1 10 9 2 10 9 2 11 2 2 13 1 11 2 15 3 13 1 10 11 2 13 15 3 0 2 3 13 10 9 0 2
24 13 3 1 13 16 15 13 1 12 1 10 3 0 9 0 1 10 0 9 2 1 9 0 2
42 10 9 1 10 9 2 13 1 10 9 3 9 0 1 10 11 2 13 13 10 9 1 10 10 9 2 0 2 0 7 0 2 7 3 13 15 1 10 0 9 0 2
43 13 2 1 9 1 9 7 9 2 9 1 9 2 13 1 10 9 1 10 9 1 10 9 0 7 1 10 9 1 9 7 9 2 11 13 13 3 15 1 13 10 9 2
45 10 11 2 11 2 13 1 13 10 9 1 12 9 1 9 2 2 1 13 13 9 1 10 9 13 1 10 9 1 10 9 1 9 0 2 2 13 1 10 11 10 9 2 11 2
18 3 1 10 9 2 10 11 13 10 11 2 10 9 11 7 10 11 2
20 10 9 13 13 1 9 2 16 10 9 3 13 1 10 9 12 2 12 2 2
34 10 9 0 1 10 9 13 13 1 12 9 1 9 2 1 15 12 9 13 1 10 9 1 10 11 1 11 7 10 0 1 10 9 2
51 1 11 13 13 12 9 2 2 10 9 0 1 9 13 1 10 9 1 10 12 9 1 9 2 2 13 2 1 10 2 1 10 9 2 9 2 9 2 9 7 1 10 9 1 10 0 9 0 1 9 2
6 11 13 10 9 1 11
11 2 3 13 10 9 3 1 10 9 0 2
23 13 1 10 9 1 9 1 9 0 2 10 9 1 10 9 0 0 13 10 9 1 9 2
39 11 2 12 9 2 9 1 12 2 3 13 3 1 10 9 1 10 9 0 0 2 3 13 10 9 2 10 9 2 10 9 1 9 2 3 10 9 0 2
44 9 0 1 10 11 1 9 0 1 10 11 2 13 11 1 13 9 13 1 9 1 9 1 10 9 7 13 10 9 0 1 10 9 15 13 10 0 9 1 9 1 0 9 2
3 9 1 12
3 10 9 0
28 10 9 13 1 10 9 1 10 11 13 13 3 10 9 1 15 13 13 2 1 10 10 9 1 9 7 9 2
29 13 1 10 9 1 13 1 10 11 2 1 11 2 1 10 11 2 3 10 9 1 10 12 9 15 13 13 3 2
29 9 0 13 15 15 13 2 1 11 2 10 11 7 10 11 2 7 15 13 1 10 9 1 10 9 2 1 12 2
29 11 2 9 1 10 11 2 13 12 9 1 13 10 11 2 1 10 9 1 15 2 9 2 11 13 3 12 9 2
15 0 1 10 9 2 10 0 11 13 1 13 9 1 15 2
18 3 2 13 4 1 13 1 9 1 10 9 1 9 13 1 10 9 2
27 11 13 13 1 13 13 11 1 10 9 2 3 1 15 15 13 13 1 13 10 9 15 3 13 10 9 2
14 11 3 13 10 9 2 7 10 15 13 10 10 9 2
31 10 11 2 0 1 10 9 13 2 13 3 13 1 10 9 2 3 13 10 0 9 1 10 11 2 13 1 10 0 11 2
11 10 9 3 0 1 13 9 1 10 11 2
26 10 11 13 10 9 0 1 13 2 9 2 1 10 9 1 10 11 1 10 9 1 13 7 13 9 2
33 13 10 9 1 10 11 15 13 0 9 15 13 4 13 1 10 9 3 1 10 9 0 2 1 15 13 13 2 0 11 0 2 2
1 11
14 10 9 3 13 1 13 9 1 9 0 1 10 11 2
25 11 13 10 9 1 9 9 2 0 2 1 15 13 16 10 9 13 1 10 9 9 1 10 11 2
29 10 11 13 15 3 3 3 1 10 11 1 10 0 9 2 7 13 1 4 13 1 10 9 13 3 1 10 11 2
19 3 2 13 3 9 1 11 1 10 11 2 15 13 13 1 10 10 9 2
1 9
28 1 10 9 1 10 10 9 0 2 10 9 1 10 0 1 10 11 3 13 3 16 10 9 1 10 9 0 2
50 3 3 10 9 0 1 11 13 16 2 10 9 13 10 9 2 3 1 10 9 0 2 1 13 1 10 9 10 0 1 10 9 0 2 1 10 0 9 1 10 10 9 7 1 13 10 9 0 2 2
9 3 15 3 13 10 9 10 11 2
28 1 11 2 10 9 1 10 0 13 13 1 10 9 2 15 10 9 1 10 11 2 3 0 2 13 7 13 2
24 1 10 11 2 13 10 9 0 3 10 9 13 2 3 2 10 10 9 1 10 9 1 11 2
5 2 11 2 1 11
6 13 10 9 1 10 9
21 16 10 9 1 9 3 13 1 15 2 11 13 13 10 0 9 1 13 10 9 2
44 3 10 2 9 0 2 1 10 10 9 13 2 3 3 2 0 9 13 2 1 0 9 2 10 9 1 9 1 10 9 15 13 2 3 10 10 9 1 10 9 13 0 9 2
36 1 10 9 1 10 9 13 1 0 9 0 0 1 10 9 1 10 9 2 1 10 9 1 10 9 15 13 1 13 1 10 9 1 10 0 2
8 10 9 13 3 1 10 9 2
20 3 10 0 15 13 1 13 1 10 11 2 1 13 1 9 1 11 2 11 2
42 3 1 13 13 1 9 1 9 1 10 0 9 1 10 9 2 15 13 1 13 1 9 0 3 0 2 9 7 9 2 0 2 2 2 10 9 13 3 0 9 0 2
14 1 9 2 11 7 11 13 15 1 10 9 1 9 2
25 1 10 9 2 11 2 11 2 1 9 2 2 11 7 11 2 1 9 2 13 3 1 10 0 2
4 11 1 9 0
32 3 13 9 7 9 1 10 9 1 10 11 2 10 11 2 3 1 3 3 13 9 1 10 9 0 2 13 10 9 7 9 2
34 10 9 13 13 15 15 13 16 13 1 10 9 15 3 13 1 10 9 7 1 10 9 1 10 9 2 10 9 7 9 1 10 9 2
48 13 3 2 7 16 10 9 1 10 9 0 1 9 2 10 9 15 13 13 9 2 13 13 1 9 2 15 13 16 10 11 13 2 1 13 2 1 12 1 9 2 3 2 1 10 0 9 2
50 3 1 10 2 9 2 2 13 15 3 13 16 1 10 11 15 13 1 9 1 9 2 16 13 13 1 10 9 10 9 3 2 1 10 9 2 15 13 10 9 1 10 9 1 9 1 10 9 0 2
26 3 1 10 9 1 10 9 15 13 10 9 1 10 9 3 0 13 1 9 0 1 9 1 10 9 2
34 1 13 10 9 1 2 11 11 2 7 1 11 2 11 2 2 13 10 9 1 11 2 11 7 11 2 1 9 1 10 9 1 11 2
37 10 9 1 11 7 11 13 10 0 9 7 9 1 10 9 1 11 2 13 15 3 1 10 9 1 10 9 1 10 9 0 0 1 10 9 0 2
59 1 3 15 13 13 1 10 9 1 9 1 10 9 1 10 11 2 1 10 9 1 10 15 15 13 1 10 9 1 10 9 0 1 10 11 2 10 9 1 11 13 10 0 9 1 10 9 1 9 1 2 9 2 1 10 9 0 13 2
51 1 10 0 9 1 10 9 2 1 10 9 13 2 12 13 13 1 10 9 1 9 7 12 13 7 12 13 13 1 10 11 2 13 11 1 10 9 1 9 1 10 9 1 11 2 9 1 10 11 2 2
11 12 15 13 3 13 1 10 9 1 9 2
31 9 1 10 11 2 3 0 2 13 9 1 12 9 0 7 12 13 1 9 2 1 10 9 12 1 9 2 1 10 11 2
8 10 9 13 13 1 10 9 2
33 11 13 16 10 2 0 9 1 9 0 1 10 9 1 9 13 13 16 10 11 3 13 3 1 9 0 2 3 1 10 9 2 2
11 9 2 3 13 3 10 9 1 10 9 2
39 13 10 10 9 2 10 9 15 13 9 1 9 0 2 10 9 13 1 10 9 0 2 15 1 10 0 2 7 1 10 9 0 2 3 15 13 1 11 2
6 3 2 3 13 9 2
10 1 9 3 13 10 9 1 10 9 2
46 10 9 0 2 1 9 1 9 2 7 16 10 9 1 10 9 0 13 13 1 9 2 10 9 3 15 13 3 1 10 9 0 2 0 2 11 2 15 13 1 10 9 1 10 11 2
6 9 1 9 13 10 9
68 1 10 9 0 15 10 11 13 4 1 13 1 10 9 1 10 0 9 1 9 1 9 1 9 2 10 9 1 3 1 10 9 0 0 13 1 13 15 3 13 1 10 9 1 9 2 1 10 0 9 1 9 1 10 0 9 1 13 0 1 10 9 1 10 9 1 3 2
8 9 0 1 10 9 1 10 11
5 15 13 1 10 9
9 13 9 1 10 9 1 10 11 2
37 10 9 13 1 10 9 0 13 1 4 13 7 10 9 1 10 9 13 16 13 9 1 9 1 10 15 13 1 10 9 1 10 2 9 0 2 2
30 9 3 15 1 10 11 2 11 7 11 13 1 9 3 0 10 9 15 10 9 13 13 1 10 9 13 1 10 9 2
79 1 10 11 2 10 9 13 1 12 3 13 3 1 13 10 9 1 12 12 9 13 1 10 0 9 2 15 1 1 10 9 1 10 9 1 10 0 9 1 12 13 13 16 2 15 13 1 10 0 9 10 0 9 1 10 9 1 10 9 1 10 9 2 7 1 0 1 10 9 1 10 9 7 1 10 9 9 2 2
31 3 2 7 15 13 13 10 9 0 1 10 10 9 2 11 13 16 10 9 1 10 0 9 13 13 1 11 10 9 0 2
37 1 10 9 0 0 2 1 15 11 13 10 9 1 10 9 2 13 1 3 0 16 10 9 0 13 1 13 1 13 3 1 10 9 1 10 9 2
33 15 13 13 15 1 0 9 16 10 9 13 1 11 2 3 13 10 9 12 9 7 12 9 13 13 1 10 9 1 2 9 2 2
23 1 10 9 2 10 9 1 10 9 13 15 1 10 9 1 10 9 1 13 1 15 13 2
31 3 1 10 9 1 10 9 3 11 13 13 1 13 10 9 2 13 3 10 9 1 10 9 3 13 1 10 0 9 0 2
35 11 2 9 0 1 10 11 2 13 10 9 1 10 9 0 2 2 15 13 10 9 1 10 10 9 7 1 10 9 13 1 10 9 2 2
28 2 15 13 16 10 9 1 11 13 3 0 3 2 1 12 9 2 10 9 13 3 1 15 13 9 0 2 2
64 11 2 10 9 7 9 0 2 13 10 9 0 15 10 10 9 13 1 13 2 3 1 10 9 1 10 9 2 1 10 9 0 13 1 13 9 7 9 2 10 9 15 13 10 9 0 2 10 9 13 7 13 1 9 0 2 1 16 10 9 13 10 9 2
1 11
13 2 13 10 9 1 3 13 15 13 3 10 9 2
4 1 2 11 2
20 2 13 10 9 15 13 3 3 13 1 10 11 1 9 13 3 1 10 11 2
34 13 1 13 12 9 3 0 1 9 1 10 9 0 2 1 10 9 1 9 1 10 9 1 10 9 7 1 10 9 1 13 1 15 2
12 2 2 2 7 10 9 0 13 3 10 15 2
19 13 13 15 9 3 0 3 1 10 9 0 7 15 3 13 1 10 9 2
16 10 0 1 15 13 13 15 1 10 9 0 7 0 0 2 2
15 11 13 1 11 2 1 11 2 1 15 9 12 1 9 2
22 3 1 10 9 1 11 2 1 13 10 9 1 10 9 2 1 10 9 1 10 9 2
29 7 13 10 9 1 9 1 9 7 9 1 10 9 2 1 10 0 9 1 10 9 1 10 9 1 10 9 0 2
43 16 13 9 1 9 15 13 13 3 3 1 10 0 9 1 9 0 15 13 1 10 0 9 1 10 9 13 7 10 0 9 1 10 9 2 15 13 3 15 13 1 11 2
44 11 13 3 10 9 1 10 9 0 2 1 10 9 0 0 2 10 11 2 7 10 9 3 0 9 2 10 11 2 13 3 10 11 0 2 11 2 13 9 1 9 1 12 2
91 2 13 0 13 16 13 11 15 13 11 2 7 3 2 7 13 0 16 11 13 9 0 7 0 2 16 15 13 1 10 9 1 10 9 0 2 2 13 11 2 13 10 11 2 1 10 11 2 10 11 2 1 10 11 2 10 11 2 1 10 11 2 10 11 2 1 10 11 2 10 11 2 1 10 11 2 7 10 11 2 1 10 11 2 10 2 0 1 9 2 2
6 9 2 1 10 0 2
34 10 9 0 7 10 9 1 10 9 3 0 13 1 10 9 2 7 11 13 15 15 13 0 9 1 9 13 1 9 2 3 12 9 2
43 1 10 0 9 1 10 9 13 10 11 13 10 9 1 9 1 12 9 2 1 10 9 7 13 12 2 3 2 12 9 1 10 9 2 15 13 1 10 9 1 10 9 2
32 3 3 1 15 2 3 2 3 10 11 15 13 3 13 2 16 13 1 13 13 10 9 1 9 2 16 2 15 3 15 13 2
11 10 9 13 13 1 10 15 2 1 15 2
12 1 15 13 9 0 2 16 13 10 9 13 2
22 3 13 0 1 10 9 1 10 9 0 2 15 1 10 9 13 1 10 9 1 9 2
20 13 13 3 10 9 15 13 1 10 9 2 15 13 0 1 10 9 1 9 2
22 3 2 13 10 9 7 16 15 13 16 13 10 9 0 1 15 2 13 1 9 2 2
7 13 13 15 13 4 13 2
30 2 3 13 16 10 9 3 2 3 0 1 10 9 2 7 3 10 11 2 1 9 2 16 13 0 1 10 9 2 2
8 1 10 10 9 2 11 13 2
12 2 3 13 9 2 3 13 13 10 9 2 2
7 7 13 16 13 13 3 2
27 15 13 1 15 0 7 15 0 9 1 10 9 13 2 3 2 10 9 1 9 2 10 9 1 10 11 2
41 3 10 0 9 1 9 13 1 16 10 9 1 10 9 1 11 3 15 13 13 2 15 2 3 2 13 10 9 1 2 13 2 10 9 1 10 9 1 0 9 2
91 3 2 1 10 10 0 11 2 11 3 9 2 1 10 9 11 2 11 13 1 10 9 7 1 11 1 3 13 13 1 10 11 2 11 13 13 1 13 1 10 9 7 1 9 10 0 9 2 13 3 3 3 16 10 10 9 0 15 2 0 7 0 2 13 10 10 9 1 15 13 1 10 2 9 2 0 1 15 11 7 11 13 13 3 2 1 1 10 9 2 2
56 3 11 13 13 1 10 11 7 15 13 13 2 1 10 2 11 7 11 2 10 9 1 11 13 15 7 2 1 10 10 9 2 13 1 13 15 1 10 9 1 10 9 15 2 3 2 13 13 13 1 10 9 1 10 9 2
42 11 13 10 9 2 7 13 0 16 11 13 1 13 10 9 1 2 9 2 1 10 9 2 1 9 1 10 9 2 16 13 10 9 15 15 13 10 9 1 10 9 2
11 13 16 13 10 9 1 1 10 0 9 2
28 1 10 9 1 10 11 2 10 12 9 13 13 1 10 9 11 2 10 9 0 7 3 15 0 1 10 9 2
22 10 10 0 13 11 2 9 2 2 11 7 11 2 13 2 7 11 2 3 9 2 2
39 9 2 13 15 0 2 1 10 9 0 2 1 9 0 3 10 10 2 16 2 1 10 0 2 10 9 7 10 9 13 10 9 0 1 15 1 10 9 2
16 9 2 15 13 13 10 9 10 9 3 0 2 1 10 0 2
18 13 3 1 10 9 10 0 9 1 10 9 1 10 11 2 11 2 2
21 1 10 11 2 1 11 2 10 9 1 11 13 10 0 9 1 9 1 10 11 2
80 10 9 0 13 13 1 10 9 1 10 9 2 13 2 10 9 1 9 2 2 2 13 10 9 3 9 1 10 9 7 1 9 1 9 15 13 9 1 10 10 9 2 2 1 10 9 15 13 2 1 10 9 2 2 13 1 10 9 1 9 7 9 15 15 13 1 10 9 1 9 7 9 15 15 13 1 0 9 2 2
17 3 2 10 9 13 13 9 13 1 15 15 15 13 13 1 9 2
37 10 9 0 1 10 9 2 11 2 2 13 1 10 11 7 15 10 11 13 2 13 3 13 1 10 9 0 1 13 10 9 0 7 1 13 15 2
64 13 10 9 3 1 10 9 1 10 9 1 11 13 10 9 3 0 2 16 13 10 9 0 2 16 13 10 9 15 13 2 1 10 2 1 10 9 0 1 10 9 13 1 10 11 1 10 9 0 2 16 13 13 1 10 9 3 0 1 10 9 0 0 2
15 11 13 15 1 10 9 1 10 9 1 10 9 1 9 2
36 1 10 9 2 13 9 1 10 10 9 7 9 2 13 9 1 9 7 13 13 2 3 1 10 9 0 0 2 10 9 1 10 9 0 0 2
24 10 9 1 9 1 11 2 1 10 10 11 2 7 11 2 9 1 10 11 2 13 10 9 2
2 9 0
5 11 13 1 10 11
21 11 2 9 13 13 1 13 1 10 11 1 10 9 1 10 9 1 10 9 0 2
20 10 9 13 9 0 1 10 11 2 7 13 3 13 1 10 9 0 1 11 2
26 12 3 13 16 15 13 3 13 10 9 2 1 10 9 1 10 0 9 1 10 9 7 1 10 11 2
37 11 2 15 3 3 13 1 13 9 10 2 13 9 1 10 9 0 2 3 1 13 7 1 10 11 2 1 15 10 9 3 13 9 1 10 11 2
8 2 3 10 9 13 13 0 2
14 3 15 13 13 10 9 3 1 10 9 1 10 9 2
13 3 13 16 10 9 0 13 16 15 13 15 2 2
15 10 9 13 10 9 1 15 15 13 1 10 9 1 9 2
25 3 15 13 13 1 10 9 16 11 13 10 9 7 12 9 3 13 16 15 13 1 10 13 9 2
47 11 13 10 9 1 10 9 1 10 9 7 9 2 13 11 2 10 9 13 15 13 2 1 12 1 9 2 13 1 10 11 2 7 1 15 1 11 13 13 10 0 0 1 0 9 0 2
87 10 10 9 13 16 10 2 9 0 7 10 9 1 9 1 15 0 2 15 13 2 0 2 1 10 9 15 13 13 1 10 11 2 1 10 10 9 1 11 1 12 2 2 13 1 9 0 9 1 9 2 9 7 9 7 1 15 13 1 10 9 2 1 13 1 13 10 9 1 9 0 7 1 13 7 13 10 9 1 9 2 9 7 1 9 2 2
50 2 1 3 12 9 2 10 9 1 10 11 13 10 9 0 9 2 13 0 13 9 1 16 2 1 10 0 9 15 11 13 2 10 9 1 10 9 1 10 9 15 13 1 10 13 9 1 10 9 2
27 1 9 2 13 1 9 0 10 9 0 1 10 0 9 1 10 11 2 2 13 2 1 13 2 10 9 2
32 10 11 13 13 1 10 9 1 10 11 10 9 15 3 13 1 10 9 1 11 2 1 9 1 10 9 0 15 13 1 11 2
84 10 9 13 4 13 1 0 9 2 3 1 10 9 2 9 2 1 10 9 0 13 13 10 9 1 10 11 2 11 2 2 1 11 2 10 9 2 1 10 9 1 10 9 2 15 13 1 10 9 1 9 1 10 9 1 10 9 0 2 7 15 13 10 9 0 1 10 9 1 11 1 10 11 2 13 1 10 11 2 13 11 9 2 2
41 2 13 9 0 1 10 10 9 2 2 13 1 10 11 10 0 9 0 2 9 11 2 12 9 2 13 3 2 1 10 9 0 1 10 9 2 1 13 10 9 2
37 2 1 10 9 2 15 13 1 13 13 10 9 1 10 11 1 9 3 10 11 2 16 15 13 10 9 1 9 1 10 9 1 10 10 9 2 2
1 11
25 1 10 0 9 1 15 13 1 11 10 9 13 10 9 1 10 11 2 1 10 12 2 9 2 2
20 10 9 3 0 1 9 2 1 10 9 0 1 15 13 13 10 10 9 0 2
38 13 1 13 1 10 10 9 7 13 13 1 10 9 1 10 10 7 13 10 9 0 3 13 10 2 9 2 1 10 9 13 1 13 10 0 9 0 2
21 13 3 10 9 7 10 9 1 10 9 13 1 13 15 1 10 9 1 10 9 2
10 1 12 9 13 10 9 1 10 11 2
16 1 10 10 9 0 13 12 9 0 7 12 9 13 1 9 2
16 10 9 1 9 15 13 2 13 2 1 10 9 1 10 11 2
25 9 3 1 9 13 0 1 11 7 10 9 0 0 7 0 13 13 1 12 1 15 7 13 0 2
26 15 13 1 10 9 1 16 13 10 1 10 9 0 1 10 11 7 3 1 10 9 0 1 10 9 2
38 10 9 1 9 7 9 1 10 10 9 3 13 15 2 3 2 7 3 13 13 1 10 0 9 1 16 13 13 1 10 9 1 10 9 1 10 11 2
19 10 9 3 13 10 9 0 1 10 0 2 1 10 9 10 9 1 9 2
30 11 13 10 9 1 0 1 10 9 2 7 10 9 1 10 9 13 10 9 1 10 9 1 9 0 1 10 9 0 2
6 3 2 1 9 13 2
30 13 15 15 13 3 1 10 9 1 9 0 7 9 7 9 2 9 2 7 1 10 0 9 1 9 0 1 10 9 2
55 10 9 1 11 15 13 1 10 9 0 15 2 10 9 2 13 13 1 10 9 2 2 11 2 2 1 10 9 11 2 1 15 15 13 16 10 9 1 9 1 10 9 13 15 3 10 9 1 9 7 9 1 10 9 2
28 15 12 13 10 9 16 10 9 13 10 9 0 1 10 9 1 9 1 12 9 2 7 15 13 0 1 15 2
6 9 1 10 11 1 11
3 12 9 0
36 11 13 3 2 1 10 9 11 2 10 0 9 1 10 11 2 15 1 10 9 15 13 1 10 9 1 10 11 2 1 10 11 2 1 11 2
14 11 2 1 10 9 2 13 10 9 1 10 9 11 2
38 15 13 10 0 9 1 13 10 0 9 1 10 10 9 15 13 9 1 10 9 1 10 11 2 15 13 1 10 9 1 12 9 2 12 1 15 0 2
67 3 2 1 3 13 4 13 1 12 2 13 9 10 9 0 11 2 10 11 2 2 10 9 0 1 11 2 9 2 7 11 2 9 2 2 15 13 13 1 10 0 9 1 10 10 9 2 12 2 1 10 9 1 2 9 2 1 9 1 10 9 0 11 2 11 2 2
21 2 11 2 13 10 9 1 11 2 11 2 9 2 2 11 7 11 2 9 2 2
5 11 2 1 0 2
20 2 9 2 2 10 9 1 10 9 13 15 1 13 10 9 1 10 9 0 2
20 1 10 9 2 15 10 9 15 13 13 10 9 1 13 10 9 1 10 9 2
7 7 13 16 13 10 0 2
8 10 15 15 13 1 10 9 2
35 13 16 10 9 1 10 9 7 1 10 9 13 15 1 13 10 9 1 10 15 10 9 13 13 2 7 3 3 1 13 1 15 0 9 2
15 13 0 16 13 10 9 2 7 3 15 13 13 10 9 2
6 15 3 13 10 9 2
15 10 0 2 1 15 2 13 16 10 9 13 0 1 9 2
3 10 0 9
10 11 2 13 10 0 9 1 10 11 2
43 3 0 1 10 9 1 10 9 1 10 11 1 13 10 9 1 10 2 9 1 9 0 2 13 1 10 11 2 10 11 3 13 13 0 9 1 10 9 1 10 10 9 2
47 7 2 1 10 9 1 9 15 3 15 13 1 13 1 10 9 1 10 11 2 10 9 1 10 11 7 10 9 0 2 11 2 3 13 10 2 9 2 1 10 9 1 13 1 10 11 2
21 3 13 2 16 2 10 9 2 0 2 3 2 1 3 13 10 9 1 10 9 2
36 1 10 9 2 3 2 13 9 1 9 2 3 10 15 13 1 10 2 11 2 2 10 9 2 9 1 11 2 13 1 9 1 10 11 2 2
20 2 0 9 2 9 0 2 9 3 0 1 10 9 7 15 13 1 9 0 2
11 9 2 9 1 10 9 1 9 0 0 2
18 0 9 2 9 0 2 9 15 13 9 0 1 10 9 1 10 9 2
22 9 2 9 1 9 2 9 1 10 9 0 1 13 10 9 7 10 9 2 3 2 2
16 0 9 2 9 0 2 9 15 13 1 9 1 10 0 9 2
18 9 2 9 1 9 0 0 2 9 1 10 9 0 1 13 3 2 2
22 0 9 2 9 0 2 9 15 13 7 3 13 3 0 2 7 15 13 1 9 0 2
8 9 2 9 1 10 9 2 2
17 10 9 15 13 9 13 2 10 9 2 3 0 2 1 9 2 2
59 1 10 9 1 10 9 13 1 10 9 1 9 2 1 10 9 7 1 10 9 2 2 13 15 2 3 2 12 1 10 9 3 0 2 2 10 9 1 10 9 1 10 9 2 9 10 9 13 1 13 11 15 3 13 1 10 9 0 2
65 10 9 1 10 9 2 1 10 15 13 13 10 9 1 9 0 2 10 9 1 10 9 2 3 13 7 3 1 9 7 9 2 7 10 9 1 10 9 2 3 12 12 9 1 10 9 13 2 13 15 1 10 9 3 0 1 10 9 0 1 9 1 9 0 2
54 7 10 9 1 12 1 12 1 10 11 2 1 15 13 9 10 9 0 1 10 9 0 2 13 13 10 9 2 1 15 1 10 9 1 13 10 9 13 9 0 2 1 16 10 9 13 9 10 1 13 10 9 0 2
45 10 9 13 3 10 9 0 1 10 15 15 13 13 10 9 1 9 2 16 13 13 10 9 0 16 13 10 9 1 9 0 3 13 10 10 9 16 13 10 9 15 15 13 9 2
25 13 1 10 9 1 10 11 2 13 1 10 9 2 10 9 13 13 10 9 0 1 13 10 9 2
35 0 13 10 9 7 0 10 9 1 10 9 2 15 10 13 9 13 1 13 2 13 10 9 2 15 13 1 10 9 7 13 13 10 9 2
24 1 1 15 15 13 1 10 9 1 10 9 11 2 10 9 13 2 1 9 2 15 3 13 2
42 15 13 2 13 2 15 13 1 10 9 1 10 9 2 7 10 9 13 3 1 13 1 10 9 10 9 1 10 9 2 2 1 13 15 2 2 1 10 9 2 3 2
17 2 3 13 10 9 15 13 13 10 9 3 1 10 9 0 2 2
23 3 3 3 11 2 9 0 2 13 10 0 9 1 10 9 0 15 2 3 2 13 0 2
13 1 11 2 10 9 13 1 4 13 1 12 9 2
30 3 2 10 0 9 1 9 1 10 9 0 1 9 0 0 1 10 9 0 2 1 0 1 10 11 7 1 10 11 2
15 3 1 10 9 3 2 1 10 9 2 10 9 13 0 2
24 7 2 3 2 3 3 10 9 1 10 9 3 13 13 10 9 3 1 9 1 10 9 0 2
5 9 1 9 1 11
29 10 9 13 3 1 9 1 10 9 1 9 0 11 2 1 11 2 3 13 1 13 9 1 10 9 7 9 13 2
7 11 13 13 15 1 10 9
6 2 11 2 1 9 13
44 10 11 13 4 1 13 15 1 10 9 2 1 12 12 9 2 1 10 9 1 10 9 2 11 2 2 1 11 7 11 2 1 9 1 11 2 13 1 10 11 2 11 2 2
47 13 3 1 10 9 1 10 9 0 1 10 11 2 1 9 1 12 2 3 13 1 9 1 12 2 1 10 11 2 13 11 1 9 2 10 9 3 13 4 13 1 9 2 9 1 12 2
26 11 2 9 0 1 10 11 0 2 13 7 13 16 10 9 1 10 9 0 13 3 0 16 13 3 2
29 1 10 9 1 10 9 0 2 10 9 13 1 10 9 1 9 2 13 9 13 2 1 13 10 9 1 0 9 2
16 2 3 2 10 11 13 10 0 9 15 13 1 13 9 2 2
33 3 10 9 2 1 9 2 10 9 0 3 13 1 10 9 0 12 9 13 2 9 2 0 1 10 9 1 15 9 2 2 13 2
10 1 15 2 3 13 10 9 1 9 2
16 10 9 13 16 15 13 1 9 13 1 10 9 1 9 0 2
14 7 2 2 1 10 9 16 10 11 2 2 13 11 2
27 3 2 11 13 3 10 0 9 1 9 1 10 9 7 13 15 1 13 9 2 1 13 10 9 2 11 2
35 2 3 2 10 9 13 3 3 13 0 7 10 9 1 10 13 9 1 9 1 10 9 13 13 9 1 9 0 2 2 13 10 13 9 2
21 11 13 15 1 13 13 1 10 9 7 13 10 9 1 9 2 16 13 1 9 2
5 9 1 10 9 3
6 11 13 9 1 10 11
50 10 9 1 10 11 2 11 2 13 3 10 9 1 13 10 9 1 9 1 10 9 1 10 11 1 12 1 16 13 10 10 9 1 10 9 1 10 9 2 7 11 2 1 9 2 13 1 10 9 2
30 2 1 10 9 7 9 1 9 1 10 9 11 3 13 3 15 1 13 2 16 13 15 1 15 15 13 2 2 13 2
38 10 9 0 3 13 2 13 2 1 10 9 0 2 1 9 1 9 2 1 10 9 1 9 1 9 1 9 2 1 9 1 9 13 13 1 10 9 2
20 10 2 9 2 13 2 3 2 13 1 13 10 2 9 9 2 1 9 0 2
49 3 2 1 10 11 2 10 0 1 10 0 9 0 1 10 9 1 10 9 0 2 10 2 9 1 11 2 2 3 1 10 9 1 10 9 0 2 13 13 10 9 0 2 11 2 7 10 11 2
23 10 9 1 10 9 1 10 9 13 2 3 2 13 1 9 1 2 9 7 1 9 2 2
40 10 9 1 2 11 2 13 10 9 1 9 0 11 2 15 2 1 12 2 13 10 9 1 10 9 7 1 10 9 3 2 0 2 0 2 0 7 13 2 2
13 11 13 16 2 3 2 10 9 13 13 1 9 2
9 2 10 9 13 0 2 10 0 2
19 15 13 3 0 2 10 3 0 2 10 3 0 2 10 3 1 9 2 2
12 10 9 1 9 2 1 10 9 13 10 9 2
27 11 7 11 13 10 9 1 2 9 1 9 2 2 1 1 15 13 7 13 15 15 13 1 10 9 3 2
30 10 9 2 1 10 9 1 10 2 9 1 9 2 2 13 13 13 15 13 13 7 3 13 10 9 1 10 9 0 2
27 10 9 3 2 9 1 13 1 15 1 10 9 2 13 13 15 16 15 13 3 7 13 2 13 15 2 2
27 12 1 11 2 9 0 1 9 1 10 9 1 11 2 9 1 10 11 2 13 4 13 1 13 1 11 2
23 10 11 2 10 11 2 10 11 7 10 11 13 10 9 1 10 9 12 1 9 1 11 2
11 12 1 11 2 2 13 15 9 0 2 2
11 3 12 12 0 13 10 10 9 1 11 2
24 13 10 9 1 3 12 9 1 10 11 7 10 9 1 10 9 13 1 10 10 9 1 9 2
9 2 10 9 13 1 10 9 2 2
20 1 10 12 9 2 10 9 11 13 1 10 9 2 13 10 9 1 10 9 2
17 10 0 13 1 10 9 2 13 9 0 7 13 2 6 11 2 2
2 9 13
48 10 9 1 10 11 2 9 11 2 13 13 1 10 9 1 10 9 1 10 11 2 11 2 2 13 4 13 2 1 10 13 9 2 10 9 1 10 9 11 2 1 10 9 1 10 9 0 2
27 3 2 10 9 11 13 13 10 9 1 10 11 2 7 2 1 10 0 9 2 13 13 10 9 3 0 2
25 13 0 16 10 9 0 0 13 3 0 13 9 0 2 3 3 15 1 9 0 2 0 7 0 2
39 10 9 13 1 9 3 15 13 13 1 10 9 10 9 15 13 1 13 10 10 9 7 9 1 10 9 1 9 15 1 10 9 7 1 10 9 13 9 2
46 7 3 13 1 9 3 15 13 10 9 1 10 9 1 10 9 1 10 9 2 13 13 16 15 13 1 9 1 13 9 0 2 0 7 0 2 1 15 10 9 0 13 0 9 0 2
43 10 9 13 3 16 3 13 9 1 15 13 10 9 0 1 10 9 2 16 13 10 9 1 10 9 1 10 9 15 13 16 15 13 3 1 10 9 3 0 1 10 9 2
32 2 3 1 12 2 10 9 13 0 7 2 3 2 13 1 13 9 0 1 10 9 1 15 10 9 3 13 3 3 0 2 2
33 7 13 16 2 1 3 1 10 9 2 10 11 2 15 13 10 9 0 1 13 12 9 2 13 1 13 3 15 2 10 9 0 2
11 10 9 1 10 9 0 13 1 10 9 2
51 10 2 11 2 2 15 13 1 4 13 12 9 1 9 2 13 1 13 10 10 9 2 13 10 9 2 11 2 1 13 15 10 9 0 2 15 2 1 11 13 2 13 10 9 1 9 1 10 0 9 2
47 7 2 1 9 2 13 15 1 10 9 1 2 11 2 10 9 1 0 11 2 1 10 9 1 10 9 1 9 2 11 2 7 10 9 2 1 11 2 1 10 9 15 13 1 10 9 2
28 11 13 12 12 9 7 13 1 9 13 1 10 2 11 2 2 13 2 1 10 10 9 2 1 11 7 11 2
11 15 13 16 10 9 13 3 1 10 9 2
6 11 2 3 3 13 2
21 13 13 10 9 0 1 10 9 1 10 9 0 2 10 9 0 7 10 9 0 2
32 16 13 1 11 2 10 0 9 1 9 15 3 13 1 9 3 13 1 10 9 0 7 1 10 9 0 2 7 1 10 9 2
20 13 9 3 13 15 2 1 15 2 3 13 13 13 10 9 1 10 10 9 2
30 3 2 1 10 11 2 15 1 3 13 3 3 13 2 10 9 13 13 15 1 9 7 13 1 10 9 1 10 9 2
12 3 2 15 13 13 15 1 10 9 0 0 2
17 11 2 13 1 3 13 13 1 16 15 13 3 1 10 9 0 2
18 16 10 9 1 9 1 11 13 13 3 2 10 9 13 1 13 15 2
15 10 9 13 10 9 2 10 9 13 1 13 9 3 0 2
27 15 1 10 9 13 4 13 1 10 9 0 1 9 2 3 3 1 11 3 1 10 11 7 1 10 9 2
9 13 10 9 0 1 9 7 9 2
45 1 10 9 13 2 11 13 16 16 11 3 13 10 9 1 10 9 0 13 13 13 1 10 9 2 16 10 9 13 1 13 13 10 10 9 1 13 7 10 9 1 15 13 13 2
45 10 9 13 10 9 1 10 9 3 15 1 12 2 9 1 15 12 12 9 15 13 1 9 1 10 11 2 3 15 1 10 10 9 3 15 13 1 13 1 10 9 1 10 11 2
43 10 9 13 13 10 9 1 10 9 15 13 2 3 10 9 0 1 10 9 3 10 9 1 10 9 1 11 15 15 13 13 3 12 9 2 13 9 13 1 10 9 0 2
23 7 13 0 10 9 1 10 10 9 1 9 2 13 15 3 10 9 0 13 1 10 9 2
62 3 13 9 2 3 16 10 9 13 2 1 10 9 1 0 9 0 2 9 2 7 9 2 9 13 13 12 9 1 10 9 1 9 2 1 11 2 7 10 9 1 11 2 1 9 2 7 16 10 9 15 13 1 13 11 2 13 1 11 7 11 2
71 3 2 10 9 3 3 13 3 1 10 11 2 1 13 16 10 9 13 13 1 1 10 9 1 10 9 2 1 10 9 0 2 1 10 9 1 10 9 11 2 13 2 2 13 1 13 3 9 1 10 9 2 10 9 3 1 10 9 15 13 10 9 1 9 1 9 1 9 0 2 2
43 7 11 2 10 9 1 10 9 2 0 2 0 1 10 9 0 2 13 0 1 15 13 1 10 9 16 2 2 1 10 0 9 1 9 2 10 11 13 13 10 9 13 2
23 15 1 10 9 13 1 10 9 3 13 2 3 2 9 1 10 9 0 15 3 15 13 2
56 3 2 3 10 0 9 13 16 16 13 10 9 2 10 11 13 10 9 1 9 1 10 9 1 10 9 2 10 9 3 13 3 13 16 2 13 4 13 1 12 1 9 1 10 0 9 9 15 13 3 10 9 0 2 0 2
37 3 2 3 13 3 10 11 1 13 15 2 7 10 9 0 1 10 9 1 10 9 13 16 2 1 3 2 2 10 11 13 13 10 9 0 2 2
28 10 9 13 16 13 0 10 9 1 10 10 9 1 10 2 9 2 7 10 2 9 2 1 10 11 13 13 2
24 2 16 15 13 10 9 2 3 13 10 9 13 15 10 9 1 13 10 11 2 2 13 11 2
38 2 13 10 9 0 1 10 9 15 13 7 3 16 3 15 13 13 10 9 9 1 9 1 10 9 0 2 13 16 13 13 1 10 9 2 2 13 2
58 1 10 10 9 1 9 1 10 9 1 10 9 2 13 1 10 9 7 3 1 10 9 2 10 9 1 9 2 10 9 1 15 10 9 15 13 7 15 10 9 13 1 13 16 10 9 13 13 2 13 3 13 10 9 1 10 9 2
17 10 9 13 3 16 11 13 1 10 10 9 15 13 13 1 9 2
6 2 15 13 3 0 2
10 10 10 9 13 3 0 2 2 13 2
45 1 10 9 1 10 9 2 10 10 0 9 1 9 1 10 11 2 11 13 9 10 1 13 3 12 9 1 10 2 9 2 2 7 3 13 3 15 15 10 9 0 13 1 11 2
43 2 10 3 0 13 13 16 13 0 1 13 9 1 10 2 9 2 2 2 13 15 2 13 15 1 10 9 1 10 11 1 11 2 0 11 2 7 11 2 0 11 2 2
26 7 10 9 3 13 13 3 1 10 9 0 2 1 10 9 1 11 7 11 1 10 9 1 9 0 2
27 10 9 0 13 10 3 0 11 7 10 9 11 1 12 2 12 2 13 10 9 7 10 9 1 12 9 2
45 2 13 13 1 10 0 9 16 13 13 15 7 16 3 13 13 16 10 9 13 3 2 2 13 11 2 15 3 13 16 15 12 13 1 13 3 12 9 3 1 10 9 15 13 2
28 11 3 13 13 0 1 10 9 1 12 2 10 0 9 1 15 10 9 13 13 3 1 10 9 1 10 9 2
1 9
13 1 11 2 10 9 13 10 9 7 3 13 13 2
34 2 3 13 1 10 9 2 13 16 3 13 10 9 2 16 10 9 13 10 9 1 10 9 2 7 1 10 10 9 13 10 9 2 2
15 3 2 13 2 2 13 16 3 15 13 1 12 9 2 2
18 1 10 9 0 2 11 7 11 13 1 10 9 2 13 1 10 9 2
19 2 1 10 9 2 10 9 13 16 3 13 10 9 2 2 13 10 9 2
9 7 10 9 3 13 1 4 13 2
32 13 15 10 9 1 9 3 0 7 11 13 1 13 10 9 2 13 13 4 13 7 16 10 0 9 1 10 9 13 4 13 2
13 10 9 13 7 13 1 10 9 1 10 12 9 2
26 15 15 13 13 3 3 1 10 9 10 10 9 13 15 7 1 10 9 9 3 13 2 2 13 11 2
9 2 15 13 1 13 9 1 9 2
22 15 13 1 13 1 15 2 1 10 9 2 1 10 9 2 1 10 15 2 2 13 2
22 3 2 11 13 13 10 9 15 13 10 9 3 13 12 9 2 1 13 13 10 9 2
34 13 1 10 11 2 11 13 3 13 2 13 10 9 3 13 10 9 1 10 9 0 1 10 0 1 10 9 0 1 10 10 9 2 2
16 10 11 3 15 13 9 7 10 10 9 3 3 15 13 3 2
9 13 13 2 1 13 9 1 9 2
23 1 10 2 9 1 9 2 0 2 13 3 12 12 2 0 2 1 10 9 1 10 9 2
11 1 3 2 13 13 12 9 1 9 13 2
6 1 13 13 10 9 2
5 1 15 13 13 2
15 1 3 13 13 1 10 9 1 15 13 1 10 9 13 2
13 1 10 9 1 10 9 2 13 10 9 1 9 2
16 10 9 13 9 1 13 1 12 9 1 10 0 9 1 9 2
16 1 10 0 9 2 10 0 9 1 10 11 13 2 13 2 2
12 3 13 10 3 13 2 9 1 9 2 0 2
8 9 13 2 9 2 1 10 11
5 9 0 1 10 11
6 2 11 13 10 9 2
14 7 1 3 13 11 2 3 13 15 13 9 9 2 2
49 1 9 0 1 10 9 2 13 10 9 1 10 0 9 1 10 9 2 10 9 2 1 9 13 2 13 1 10 10 9 10 9 1 10 12 9 0 1 10 9 13 3 1 10 9 2 1 11 2
51 3 1 13 10 0 9 7 10 0 9 1 10 9 2 10 9 13 15 1 10 9 1 10 0 9 12 1 9 2 9 2 1 10 12 9 1 10 9 2 1 10 9 1 9 1 10 11 2 10 11 2
12 2 9 11 2 13 9 3 7 1 10 9 0
4 0 9 1 11
13 10 0 9 13 15 1 3 12 9 1 10 11 2
35 10 2 9 11 2 2 1 10 11 2 13 1 4 9 1 10 9 1 9 0 7 1 4 9 1 9 1 15 13 1 10 9 1 9 2
32 10 9 13 3 13 4 13 10 9 15 15 13 13 1 9 2 2 3 13 2 1 10 9 2 7 13 13 16 15 13 9 2
95 10 9 1 10 11 11 13 13 13 9 1 10 9 0 1 10 9 2 1 15 13 10 9 1 10 10 9 2 1 2 13 13 1 10 9 1 10 9 2 2 3 13 13 10 9 1 10 9 1 15 15 13 1 10 11 2 10 0 9 0 2 2 3 1 10 9 1 10 11 15 2 1 10 9 0 1 10 11 2 15 13 13 13 1 13 10 9 2 1 10 9 1 9 2 2
44 10 2 9 1 9 2 1 15 13 10 11 13 10 9 1 10 9 1 10 9 1 10 11 2 7 3 3 10 9 0 1 10 9 1 9 1 10 9 0 13 1 10 11 2
4 13 1 13 9
9 13 1 11 7 11 2 15 13 2
11 2 15 13 10 9 13 9 7 9 2 2
19 2 10 9 7 9 1 10 9 13 15 1 10 9 3 13 10 9 2 2
22 13 16 15 13 1 9 0 2 16 10 9 2 9 2 3 15 13 1 15 13 9 2
24 13 10 12 0 9 2 3 2 2 7 13 9 0 1 10 9 1 10 9 7 1 10 9 2
26 3 15 13 15 11 2 11 2 10 9 13 1 10 9 7 15 13 10 9 1 11 1 10 0 9 2
18 7 11 2 15 13 3 0 9 7 10 13 9 13 1 10 0 9 2
20 13 11 2 11 2 11 2 11 2 15 13 10 9 1 10 10 9 7 9 2
15 10 9 2 7 0 7 0 2 10 9 1 9 13 13 2
16 13 0 16 10 9 13 13 1 10 9 0 2 7 15 13 2
6 10 9 13 1 11 2
6 7 10 2 9 2 2
11 3 2 13 0 1 13 15 15 7 3 2
13 3 2 13 10 9 1 9 15 13 13 1 10 11
22 10 9 1 10 9 1 9 0 13 2 3 0 2 3 1 10 9 1 10 3 0 2
16 1 10 11 13 10 9 1 13 9 1 9 0 1 9 0 2
30 10 9 3 2 15 13 10 9 1 15 13 13 9 2 1 15 3 13 10 9 0 1 9 1 9 1 10 9 2 2
20 3 2 1 13 13 10 9 0 1 9 15 13 13 1 11 7 1 10 9 2
27 10 11 3 3 13 10 9 0 1 10 9 2 15 13 13 1 10 9 1 9 7 9 1 9 1 11 2
23 3 2 12 1 10 9 13 1 10 9 13 15 1 10 13 10 9 1 13 1 10 9 2
8 7 3 3 3 15 13 13 2
16 3 2 10 11 13 16 13 13 12 9 1 10 9 1 9 2
21 12 1 10 9 11 2 11 7 15 1 10 11 1 9 1 10 11 2 11 2 2
47 10 11 13 15 3 1 10 9 1 9 1 9 2 9 2 9 0 7 9 2 13 3 13 1 10 9 10 9 2 3 2 9 2 1 9 7 9 1 9 2 9 0 7 9 1 9 2
33 10 9 13 9 10 9 2 15 13 1 10 9 1 9 0 7 0 1 9 7 9 0 2 3 0 1 10 9 0 7 10 9 2
21 1 13 1 10 3 0 2 10 11 13 10 9 1 9 0 0 1 10 9 0 2
7 0 9 1 9 1 10 11
6 11 2 1 9 1 9
17 10 11 13 10 0 9 1 9 15 13 1 10 9 1 10 9 2
37 10 9 1 9 1 10 9 2 10 9 1 9 2 10 9 1 9 7 1 9 1 9 13 15 1 10 9 1 10 9 2 13 1 12 9 0 2
22 10 0 2 9 2 2 13 1 10 9 0 1 2 9 2 2 11 2 13 10 9 2
14 10 9 1 10 9 13 3 10 0 9 1 10 9 2
85 10 11 13 1 13 1 10 9 3 12 9 0 2 10 0 16 10 9 13 10 9 1 10 9 2 2 1 13 10 9 1 10 0 9 1 10 0 7 3 13 9 1 11 2 10 9 3 13 1 13 16 13 13 15 1 10 9 1 13 9 1 10 9 7 15 2 1 15 2 13 13 1 15 3 1 10 10 9 1 9 2 1 10 11 2
33 1 11 2 10 9 1 10 10 9 13 13 15 1 10 12 12 7 12 12 9 2 9 15 15 13 2 0 2 1 10 9 0 2
42 11 2 3 1 10 11 2 11 7 10 10 9 0 7 0 2 13 10 9 1 10 9 2 13 10 9 0 1 10 11 7 11 2 7 3 1 9 13 1 10 11 2
8 9 0 0 1 9 1 10 9
9 10 2 9 1 15 2 1 12 9
32 10 9 0 13 3 0 1 10 0 11 2 15 13 3 3 7 15 13 10 0 11 1 12 2 1 10 9 15 13 12 9 2
56 3 1 15 10 9 13 10 9 1 15 15 3 13 13 10 9 1 10 10 9 2 3 1 11 15 13 9 0 1 0 2 15 13 10 9 1 9 2 3 10 9 13 13 1 13 3 1 10 9 15 10 9 1 15 13 2
61 1 10 9 2 1 10 9 1 10 10 15 13 7 13 0 9 1 10 9 2 7 15 13 10 15 15 3 15 13 1 10 13 9 0 2 2 13 13 13 2 13 7 13 2 10 9 1 10 9 0 2 10 9 0 7 10 9 1 10 9 2
50 1 10 9 0 7 0 1 10 15 13 10 9 0 2 16 10 9 1 10 9 3 13 1 10 9 3 15 15 13 2 2 13 10 11 2 11 2 1 13 15 1 13 1 13 10 9 1 10 9 2
11 7 15 13 10 9 1 10 9 3 13 2
9 15 13 10 9 1 10 9 13 2
10 15 13 10 9 1 10 9 0 0 2
23 15 13 3 10 11 1 10 9 1 10 9 1 9 15 3 13 1 9 1 9 1 9 2
22 1 3 13 10 9 13 1 9 1 9 1 9 15 13 3 13 7 13 1 10 9 2
26 1 15 13 10 9 1 10 9 13 1 10 9 1 10 9 7 9 15 13 9 1 10 9 1 9 2
27 15 13 4 13 1 10 9 1 10 10 9 7 9 2 13 1 10 9 1 9 3 13 1 9 1 9 2
34 7 10 9 1 9 1 10 9 0 2 13 1 10 9 2 1 10 9 1 9 2 1 10 9 0 7 0 13 0 1 10 9 0 2
6 7 10 9 3 13 2
26 3 2 1 10 9 1 3 2 10 9 13 2 1 10 9 1 10 11 2 13 15 13 13 7 13 2
16 2 7 10 9 13 15 3 13 2 2 13 10 9 2 11 2
21 2 10 9 13 15 16 15 13 2 7 3 2 9 3 2 13 15 2 2 13 2
43 10 9 13 4 1 10 11 1 10 11 7 4 3 1 10 9 2 15 13 16 10 9 3 13 13 1 10 9 1 10 9 2 16 13 13 2 13 4 13 9 1 9 2
50 3 1 9 2 3 10 11 13 3 10 9 1 10 9 2 11 2 9 1 10 11 2 13 12 1 10 9 1 13 15 1 10 9 1 10 9 7 1 13 1 10 9 0 10 9 1 10 10 9 2
5 11 2 1 10 11
15 9 2 1 10 9 2 10 0 9 13 16 13 1 9 2
10 3 2 3 13 15 3 7 1 15 2
17 10 9 1 10 9 1 10 9 13 1 13 9 0 2 1 15 2
6 13 15 1 10 9 2
1 11
11 10 11 13 2 11 2 2 1 10 11 2
20 11 10 11 1 10 11 13 3 1 10 9 2 1 10 11 2 2 11 2 2
32 9 0 7 1 10 11 2 11 2 13 15 13 1 13 10 9 0 15 1 10 9 13 12 0 1 10 9 1 9 1 11 2
68 10 9 0 1 10 11 2 11 2 13 3 16 10 11 1 11 13 13 10 9 1 10 11 2 11 2 1 10 9 1 16 15 13 3 1 10 11 2 10 9 0 15 13 10 9 1 12 1 10 10 9 0 2 0 1 10 11 2 13 13 10 0 1 10 9 1 11 2
3 11 13 2
17 1 9 7 15 0 1 10 9 0 13 1 11 7 3 1 11 2
7 13 10 9 1 9 0 2
5 10 9 13 0 2
44 13 1 13 15 3 1 10 9 1 9 1 10 9 2 10 9 11 2 11 2 13 3 10 0 9 1 10 0 9 1 9 1 10 11 15 3 15 13 1 11 2 11 2 2
38 3 2 10 9 1 10 2 9 2 3 13 3 13 2 1 10 9 11 2 11 2 1 13 13 9 1 10 9 2 3 2 1 10 0 9 1 9 2
25 15 15 10 9 13 13 15 2 1 10 0 9 1 9 3 0 2 1 13 10 10 9 1 9 2
26 11 13 1 13 15 3 0 7 13 13 1 10 2 9 2 2 13 1 10 9 1 9 1 10 9 2
13 3 3 2 13 10 9 1 11 13 10 10 9 2
28 2 10 9 13 15 3 16 2 13 2 10 9 1 9 1 10 9 2 2 13 15 2 1 13 10 9 0 2
24 2 16 10 9 1 11 13 10 9 0 16 10 1 11 2 13 16 13 3 13 3 0 2 2
7 11 1 0 2 3 7 3
59 1 10 9 1 10 11 1 10 11 13 3 1 10 0 9 2 3 1 10 11 13 13 3 10 9 1 10 9 1 9 1 9 0 2 2 10 9 1 10 9 7 10 2 9 2 13 1 10 10 9 13 3 1 10 9 1 10 9 2
29 10 9 13 3 2 3 1 10 9 1 13 1 10 9 0 15 13 10 9 1 10 11 1 10 9 1 10 11 2
44 3 2 10 11 13 15 13 1 10 9 1 9 15 10 11 13 13 2 13 13 15 1 9 1 9 0 1 13 10 9 1 10 9 15 10 9 13 1 13 10 9 1 11 2
38 3 1 10 9 15 13 10 9 0 7 13 1 4 15 1 10 9 7 1 4 1 10 9 1 12 1 10 12 9 2 10 9 1 10 9 3 13 2
13 3 3 13 10 9 1 2 6 2 1 10 9 2
14 13 10 9 15 15 15 13 1 10 9 7 3 13 2
21 13 1 9 1 15 13 10 9 13 7 13 15 1 10 9 15 3 13 1 13 2
4 13 9 13 2
12 3 2 3 3 2 3 15 13 1 10 9 2
48 3 13 1 10 0 9 2 1 15 12 1 15 13 1 9 0 2 1 10 9 0 1 9 0 2 0 9 1 15 10 9 1 10 9 15 13 1 10 9 1 9 2 1 9 1 9 2 2
15 10 0 9 13 13 3 10 9 7 13 10 9 1 9 2
11 13 15 0 2 1 10 9 7 1 9 2
14 3 1 10 9 2 13 15 2 3 2 1 0 9 2
21 13 10 9 1 10 11 2 15 13 10 9 1 13 1 10 9 15 13 1 15 2
13 2 10 9 13 1 13 10 9 1 10 10 9 2
23 3 13 9 1 15 13 1 3 7 15 1 13 16 10 9 1 10 9 3 15 13 2 2
11 9 0 3 10 9 2 11 2 13 13 2
5 2 3 13 15 2
14 3 3 3 10 9 3 15 13 1 10 10 9 2 2
17 10 11 2 10 11 7 10 11 13 1 10 11 1 10 13 9 2
41 10 11 13 3 1 10 9 1 11 2 3 13 1 10 10 0 9 12 1 10 9 3 0 1 10 0 9 2 10 9 1 10 9 3 13 1 10 2 9 2 2
62 3 1 10 9 1 9 2 10 11 1 11 7 10 11 1 11 13 15 3 0 1 9 2 13 1 10 10 9 3 0 1 9 2 3 10 11 1 11 13 15 3 0 2 13 9 2 10 1 10 9 11 2 9 1 10 9 2 15 13 3 9 2
44 11 2 11 2 2 1 9 2 11 2 11 2 2 1 9 2 11 7 11 2 11 2 2 3 2 1 9 7 9 2 13 15 1 10 9 3 0 2 1 10 9 1 11 2
18 10 9 1 10 9 2 9 13 13 2 3 13 15 1 0 7 13 2
19 13 16 10 9 13 10 9 7 16 10 9 13 1 10 9 7 10 9 2
15 10 9 13 1 10 9 0 10 13 9 1 10 9 0 2
5 9 3 3 0 2
20 13 1 16 10 0 1 10 12 1 10 12 9 3 13 15 10 9 13 13 2
14 15 2 13 3 9 2 13 16 3 13 0 1 15 2
4 10 9 1 11
17 10 0 11 13 13 9 2 9 7 9 1 10 9 2 9 2 2
42 12 9 1 10 9 0 1 10 11 2 1 10 13 7 3 13 9 0 2 2 1 15 13 12 3 0 9 2 2 9 1 9 2 9 1 9 0 0 3 13 2 2
5 9 7 9 0 2
24 13 7 13 3 1 10 11 1 12 1 11 1 10 7 15 9 2 1 0 7 0 9 2 2
11 13 16 13 12 1 11 7 15 1 11 2
4 10 9 0 2
21 6 2 3 13 3 12 9 1 9 7 9 0 1 9 2 7 10 9 1 13 2
38 15 13 3 0 7 10 9 1 16 13 13 1 10 9 15 2 1 15 13 10 9 2 13 16 3 13 12 2 7 12 9 15 13 13 1 10 9 2
10 12 9 1 10 7 12 9 1 10 2
8 13 10 9 1 10 9 11 2
21 2 10 9 13 1 10 9 2 13 13 3 12 9 2 7 3 13 1 12 2 2
3 7 13 2
15 2 7 13 3 3 7 13 1 13 16 13 12 9 2 2
20 10 9 13 16 2 1 9 3 15 2 2 10 9 13 10 13 1 12 2 2
33 3 13 9 1 10 2 16 13 9 2 7 1 10 9 2 10 0 9 0 2 0 1 10 9 0 2 1 13 13 1 9 0 2
32 10 11 7 10 11 13 3 0 2 16 2 3 9 2 15 13 10 9 1 9 1 10 9 7 13 10 9 0 1 10 9 2
21 13 3 0 2 15 1 10 10 9 7 9 7 15 1 10 10 9 7 0 9 2
14 3 1 10 10 9 0 2 13 15 1 10 0 9 2
22 7 13 3 15 13 16 2 13 10 9 10 0 9 1 10 9 2 2 13 10 9 2
19 10 11 13 13 9 2 16 10 11 3 13 9 1 10 9 1 10 9 2
59 10 9 0 1 9 3 15 1 10 9 1 10 11 2 1 10 11 7 1 0 10 9 13 1 10 9 0 7 9 13 3 0 1 10 9 1 0 9 2 3 1 9 3 13 7 10 9 3 13 13 3 1 10 0 12 7 12 9 2
23 16 10 9 13 1 9 2 13 1 13 3 10 9 15 1 9 13 1 10 11 1 11 2
25 10 9 1 13 1 10 9 13 3 4 13 1 10 9 1 9 15 3 13 10 9 1 10 11 2
32 3 12 9 13 12 9 1 10 11 2 11 2 13 0 15 13 1 10 9 1 9 2 12 9 2 7 1 10 9 2 12 2
43 1 10 9 2 10 9 3 3 13 10 9 0 16 13 10 9 3 2 10 9 1 10 0 2 2 1 13 13 4 13 1 10 9 1 10 9 2 11 2 1 10 11 2
10 10 9 13 4 13 1 13 10 9 2
12 12 1 15 13 1 13 10 9 1 9 0 2
15 1 10 9 3 10 9 13 13 2 10 10 9 3 13 2
14 7 13 1 15 15 2 16 3 3 13 10 10 9 2
27 10 10 9 13 1 13 16 10 9 1 9 0 3 15 13 13 2 16 10 10 9 15 13 1 15 13 2
3 2 3 2
21 3 2 13 3 10 9 1 10 9 15 3 13 9 1 10 13 9 1 10 9 2
22 7 3 2 3 2 13 10 9 1 9 1 10 9 1 9 1 13 9 1 10 9 2
18 7 3 2 13 10 9 0 1 10 9 15 10 9 13 1 4 13 2
10 9 1 10 9 1 12 9 1 10 9
4 11 13 1 11
54 3 1 10 9 1 9 0 2 10 9 1 9 1 10 11 13 3 10 10 9 1 9 2 13 10 9 1 10 9 1 12 2 1 11 2 1 10 9 1 12 9 13 1 11 1 12 9 1 10 9 1 10 9 2
28 1 10 9 2 10 11 13 15 1 10 0 9 1 10 2 11 2 2 3 10 11 13 10 11 1 10 9 2
48 2 10 11 13 10 9 0 1 10 9 1 10 9 1 10 9 2 7 3 13 0 16 10 9 15 13 1 10 11 3 7 3 13 10 9 1 10 9 2 2 13 11 2 0 1 10 11 2
26 2 3 10 9 13 3 13 2 15 13 13 1 10 11 2 7 3 13 15 15 13 16 13 9 2 2
31 3 2 13 0 10 10 9 1 9 1 13 10 9 1 10 11 2 13 11 2 9 0 1 10 2 9 2 1 10 11 2
29 7 10 9 1 9 2 13 10 11 2 13 1 13 9 1 10 9 2 13 16 3 13 10 9 1 10 10 9 2
53 10 0 9 13 10 9 2 13 10 9 1 2 9 0 2 7 13 13 2 10 9 1 10 9 1 9 7 1 10 9 2 1 10 9 2 16 15 13 2 13 3 1 10 9 2 13 1 10 9 15 15 13 2
40 13 1 10 9 1 2 11 2 2 0 2 7 2 11 2 2 9 2 7 1 11 2 10 2 11 2 13 10 9 13 1 0 9 0 2 3 1 9 0 2
56 1 10 11 2 10 9 2 13 1 10 0 12 9 1 9 1 3 12 9 1 9 2 13 3 13 1 10 11 7 1 10 11 2 2 3 13 4 13 10 9 2 10 9 13 4 13 1 10 9 1 10 2 11 2 2 2
56 10 9 13 1 10 2 11 2 3 13 0 1 10 9 13 13 1 10 11 3 2 9 1 9 0 1 10 9 1 10 9 2 2 13 15 1 2 0 10 9 1 9 3 13 0 7 15 13 9 0 7 9 3 0 2 2
27 10 9 1 10 11 1 11 13 10 9 1 10 9 7 10 9 1 10 9 1 10 10 9 1 10 11 2
28 10 9 13 13 1 10 9 0 7 2 1 10 9 2 3 10 9 1 10 9 0 13 1 10 9 13 13 2
24 13 10 9 1 9 3 10 9 1 10 9 0 7 11 13 0 1 9 3 0 1 9 13 2
36 13 15 13 1 10 9 7 13 0 3 13 9 0 2 3 0 1 10 9 2 1 13 10 9 1 15 13 10 9 1 10 9 12 1 9 2
30 1 10 9 7 1 10 9 2 1 1 10 9 2 15 13 2 1 10 10 9 2 10 9 0 1 10 9 1 12 2
3 7 3 2
7 13 10 9 2 10 11 2
18 16 13 12 9 0 1 10 11 7 2 3 2 10 11 13 10 11 2
8 3 13 10 9 13 12 9 2
9 1 10 9 13 3 0 10 9 2
76 16 2 13 10 9 2 13 10 0 9 1 10 9 2 2 10 9 0 1 10 9 2 10 9 1 9 0 1 10 10 9 2 10 10 9 0 7 10 9 16 10 9 1 10 9 3 13 10 1 10 9 1 9 1 10 9 0 7 0 2 13 10 9 0 1 10 9 1 10 9 15 15 13 9 2 2
19 15 2 13 2 2 1 10 0 9 1 9 2 1 9 7 1 9 2 2
65 10 2 9 0 2 15 10 9 13 13 1 10 9 13 1 15 13 3 0 1 10 2 9 1 9 7 1 13 9 0 2 3 10 0 2 7 15 13 2 1 15 2 3 0 1 10 0 9 1 9 1 10 9 2 1 10 3 0 9 1 0 7 0 9 2
31 10 0 9 15 15 13 1 10 9 15 13 13 10 9 1 9 1 11 13 15 1 9 1 9 1 9 13 1 10 9 2
40 1 9 0 2 3 13 2 1 9 0 1 13 7 0 2 10 9 3 0 13 1 13 1 9 0 2 3 15 13 1 9 1 9 0 7 1 10 0 9 2
25 16 1 10 11 13 9 0 7 0 3 0 1 13 10 9 2 1 10 0 9 0 15 3 13 2
38 1 10 0 9 0 1 11 2 10 11 2 10 9 0 13 2 1 9 0 2 13 10 9 15 13 10 9 7 15 1 10 9 13 13 15 3 9 2
35 10 9 1 10 11 3 13 3 1 10 10 9 2 13 15 3 2 16 3 13 10 9 1 10 11 0 1 13 9 2 3 10 11 2 2
19 1 10 0 1 10 9 13 11 2 15 13 13 13 3 1 10 0 9 2
32 10 2 9 2 13 3 2 1 9 2 1 10 9 13 1 10 11 2 15 13 10 9 1 10 9 1 10 9 1 10 11 2
16 3 1 10 0 9 2 10 9 13 13 1 13 9 1 10 9
9 11 13 2 12 2 10 11 1 11
5 10 2 9 2 13
19 10 9 2 10 11 3 3 13 13 13 3 12 9 1 10 9 1 11 2
20 13 15 3 2 13 10 11 3 13 7 13 3 10 2 9 2 1 10 9 2
13 7 2 1 10 9 2 3 15 13 1 10 9 2
3 11 3 13
27 10 9 1 12 9 0 7 12 1 10 9 1 10 11 13 3 12 1 10 9 0 1 10 9 9 0 2
16 13 1 10 11 2 11 2 2 10 9 13 13 1 10 11 2
26 1 10 9 1 10 10 9 0 2 13 1 0 1 10 9 7 13 13 1 13 16 13 9 1 11 2
41 15 13 4 10 10 9 1 10 9 2 4 2 3 2 7 4 15 1 10 9 0 2 2 13 11 2 13 16 10 0 9 1 9 13 1 10 0 9 1 9 2
27 2 13 10 0 9 15 13 10 10 9 2 1 15 15 15 13 4 7 4 16 10 9 13 13 1 3 2
17 9 3 13 10 0 9 1 15 13 2 16 3 15 13 13 2 2
27 11 13 16 10 9 1 11 3 13 9 7 9 2 9 3 2 0 2 2 2 15 2 7 2 3 2 2
29 11 3 15 15 13 1 10 9 7 13 15 1 10 0 2 9 2 2 15 1 9 1 9 0 13 2 13 2 2
53 1 10 9 1 10 11 13 0 13 11 3 3 1 15 13 3 7 2 1 10 9 1 10 9 2 10 2 3 0 1 10 2 2 2 13 10 9 1 13 15 15 1 10 15 3 2 0 2 7 2 0 2 2
17 7 11 13 1 10 2 11 2 15 13 1 10 9 2 0 2 2
6 2 13 10 9 0 2
12 13 10 10 9 2 10 9 1 13 9 0 2
24 1 13 10 0 9 7 2 3 1 15 15 15 13 2 13 3 2 2 15 15 3 2 2 2
5 13 10 9 0 2
5 13 1 9 0 2
4 9 1 13 2
10 13 9 15 1 10 9 3 13 13 2
12 10 10 9 15 13 1 10 9 13 0 2 2
15 10 9 11 13 3 1 10 0 9 7 1 3 10 0 2
17 3 2 13 1 13 12 0 9 0 1 11 2 13 3 1 11 2
56 10 13 9 13 16 10 9 1 10 0 9 1 10 9 2 1 1 10 9 1 12 13 13 10 9 1 3 12 2 11 2 11 7 11 2 2 13 13 10 9 1 9 2 1 12 9 1 12 1 12 9 2 2 1 12 2
27 1 9 2 10 9 0 13 3 12 9 1 10 9 1 10 9 0 2 2 15 3 13 1 10 11 2 2
27 1 10 9 2 2 10 0 9 0 7 13 0 0 7 9 0 15 13 10 9 1 10 0 9 0 2 2
29 12 9 2 10 11 13 9 1 10 11 7 10 11 2 10 11 1 10 11 7 10 11 7 13 9 1 10 11 2
14 9 0 2 3 13 13 2 10 9 1 9 13 13 2
25 9 2 13 0 9 1 10 9 1 13 9 2 13 3 3 10 10 9 2 1 13 1 10 9 2
45 1 9 13 1 10 2 11 2 2 10 11 13 15 2 1 10 9 3 3 0 16 13 1 12 2 12 2 9 1 15 13 10 9 15 13 1 10 9 1 10 9 1 9 2 2
31 3 2 13 2 2 11 13 1 10 9 1 10 9 1 10 9 1 9 2 13 10 9 0 7 10 9 0 13 0 2 2
7 11 2 0 9 1 9 2
13 13 9 15 3 2 3 13 13 10 0 9 0 2
8 3 2 3 0 2 3 13 2
10 11 2 0 1 13 7 1 13 9 2
8 9 3 0 2 7 3 0 2
3 3 13 2
12 12 1 10 9 3 0 1 10 11 2 0 2
4 7 10 9 2
10 3 2 10 9 3 0 1 10 11 2
26 2 7 10 9 13 3 0 1 10 10 9 16 15 13 1 13 13 3 1 3 15 13 1 10 9 2
6 2 7 3 13 3 2
7 10 10 9 3 13 3 2
23 15 10 9 13 13 10 9 1 9 1 10 9 0 15 13 10 9 7 9 0 1 9 2
22 15 13 13 10 9 1 1 10 9 1 13 16 10 9 1 10 11 13 10 0 9 2
25 1 13 10 0 9 1 10 9 15 13 1 10 9 0 2 10 11 13 10 9 0 13 1 11 2
3 11 13 11
31 10 11 13 1 10 2 11 2 2 1 11 2 13 3 1 12 9 13 1 10 9 1 10 9 1 10 11 2 10 11 2
20 10 11 13 1 12 12 9 3 0 2 15 3 13 13 1 12 1 10 9 2
32 13 3 11 13 10 12 9 0 15 13 10 9 2 7 3 13 16 10 11 13 1 10 9 2 13 15 1 10 2 9 2 2
27 3 2 1 10 9 10 9 1 10 9 13 0 1 15 1 9 3 10 9 2 9 2 9 7 10 9 2
21 3 12 9 2 10 9 1 10 9 3 13 9 2 1 10 9 7 1 10 9 2
34 13 3 9 0 15 13 16 10 9 13 10 0 9 2 3 2 16 13 10 2 9 2 13 12 1 10 9 1 9 1 10 9 0 2
20 10 9 1 10 9 0 13 3 0 2 16 13 16 4 13 1 10 9 0 2
39 9 2 13 3 10 9 1 10 0 2 9 2 2 15 13 1 13 9 2 7 2 1 13 10 11 1 13 10 9 2 10 9 13 13 1 10 10 9 2
6 13 15 13 1 13 2
23 10 0 9 1 10 9 13 9 0 2 3 9 13 1 9 0 2 9 2 9 7 13 2
13 7 3 13 1 13 15 1 10 9 1 10 11 2
21 15 13 10 9 2 13 10 9 1 2 9 2 7 1 10 9 2 3 15 9 2
13 11 2 3 3 13 3 2 3 15 13 13 13 2
27 13 0 2 13 15 3 1 10 9 7 13 16 2 1 15 1 9 2 13 3 3 0 13 10 9 0 2
23 13 12 9 2 10 15 0 2 7 13 10 9 15 3 13 1 10 9 1 10 0 9 2
11 3 13 9 1 13 10 9 1 9 0 2
13 11 2 13 0 2 3 3 15 1 13 10 9 2
17 13 9 1 15 13 13 10 9 15 13 10 9 1 10 10 9 2
34 10 0 2 9 2 1 12 9 13 4 13 1 9 15 13 0 9 1 9 2 3 10 9 1 9 1 9 7 1 10 9 1 9 2
47 10 9 1 10 11 7 10 11 2 15 13 10 9 1 10 9 1 10 11 2 9 7 11 13 1 9 13 1 10 10 9 2 13 4 3 13 1 10 9 2 3 10 11 7 10 11 2
22 11 3 13 9 1 0 9 1 10 0 9 1 16 3 15 15 13 1 10 10 9 2
45 13 1 10 9 1 2 13 2 1 10 9 3 3 0 2 15 1 10 9 1 10 9 2 11 13 13 1 10 9 3 2 0 9 2 2 7 0 9 1 10 9 1 10 9 2
24 3 13 10 9 1 10 10 9 2 11 2 7 10 9 1 10 9 13 3 13 1 10 9 2
23 1 10 0 9 2 13 15 1 10 9 1 9 1 10 9 15 13 1 10 9 10 9 2
49 3 10 9 0 13 13 10 9 1 9 1 9 1 13 1 9 7 3 9 2 13 3 0 10 9 1 9 1 9 0 1 9 0 1 13 3 9 15 10 9 3 13 1 10 9 7 10 9 2
7 13 9 1 9 1 10 11
31 13 13 10 9 1 10 9 1 10 9 15 2 9 2 13 13 1 10 9 2 1 10 9 1 10 11 2 1 10 11 2
35 2 10 9 13 0 2 13 3 3 2 7 10 9 13 0 2 15 13 0 10 9 1 10 9 2 2 13 10 9 1 10 11 2 11 2
21 3 1 15 13 11 7 10 10 9 2 10 9 2 3 2 13 13 1 10 11 2
40 2 10 9 11 2 15 13 1 11 1 10 11 2 13 15 16 3 13 9 13 10 9 3 13 1 10 9 2 2 13 3 1 10 11 10 0 9 2 11 2
45 2 12 1 10 9 16 15 13 15 3 13 13 16 13 1 10 11 9 3 13 1 10 9 1 12 12 9 2 2 13 12 1 10 10 9 1 10 11 0 15 3 13 10 9 2
50 11 2 15 13 3 9 0 1 10 9 1 10 9 1 11 2 13 16 3 15 13 1 13 13 13 1 10 9 2 7 13 16 10 9 15 13 1 16 2 10 9 13 9 15 13 1 4 13 2 2
43 10 9 1 3 1 10 11 13 15 3 1 10 10 9 3 13 1 10 9 1 9 2 15 13 10 9 1 10 9 1 9 2 15 15 13 13 3 15 13 1 10 9 2
51 1 10 9 1 13 10 9 2 10 11 13 1 0 1 10 9 10 9 0 1 9 1 9 1 1 10 9 1 12 9 1 9 2 1 10 9 1 11 2 11 1 12 9 7 1 10 9 1 12 9 2
16 1 10 9 13 1 10 9 2 3 13 13 12 9 1 9 2
18 10 9 11 13 2 1 10 9 13 2 9 0 13 1 12 12 9 2
67 10 9 13 13 1 10 9 1 9 0 1 10 10 13 11 2 3 13 1 10 11 2 1 10 9 1 12 12 9 2 2 1 9 1 3 13 1 10 10 9 9 0 1 9 0 1 9 1 9 2 3 0 1 9 0 0 2 2 13 10 9 1 10 9 3 13 2
12 3 0 2 10 11 13 9 1 12 12 9 2
50 10 9 1 9 13 1 12 9 1 9 2 10 9 0 13 13 1 12 9 1 9 2 1 12 12 9 13 1 12 2 2 3 10 9 0 13 12 12 9 2 3 12 9 16 1 10 9 0 2 2
11 9 0 1 10 9 1 10 9 13 0 9
7 10 0 9 1 10 9 9
19 13 0 9 0 7 13 13 13 1 10 9 1 10 9 1 10 9 11 2
4 10 10 9 2
23 3 15 13 13 3 3 15 13 4 4 3 13 1 3 13 1 10 9 13 1 10 9 2
22 7 13 0 16 10 9 15 15 13 13 10 1 15 13 13 10 9 15 13 10 9 2
27 13 15 1 12 1 10 9 0 13 1 10 11 2 1 10 9 1 10 9 1 9 1 9 1 10 9 2
40 11 13 15 1 13 16 10 9 3 13 4 13 7 10 10 9 2 11 2 13 10 9 1 10 9 13 13 7 13 13 1 11 2 13 10 9 13 1 15 2
24 10 9 0 13 1 13 12 9 1 10 11 7 12 9 1 10 11 2 1 13 10 9 13 2
28 1 10 0 2 13 15 10 9 11 2 9 1 11 7 15 15 13 1 10 9 13 2 1 9 1 10 9 2
18 10 9 1 10 11 13 1 10 0 11 2 1 9 1 0 9 0 2
21 2 10 9 15 13 10 9 1 10 9 7 3 10 9 2 2 13 11 2 9 2
40 1 10 9 0 2 15 0 13 1 10 9 2 10 11 13 9 0 7 9 2 9 0 7 10 9 1 9 2 13 3 1 10 0 9 1 10 10 9 0 2
32 7 10 9 1 10 10 9 13 2 10 9 0 0 2 10 9 7 10 9 0 13 2 1 9 0 2 10 9 1 10 9 2
29 3 2 10 9 1 9 1 9 13 13 3 10 9 0 3 0 2 16 13 2 3 2 0 9 2 13 9 2 2
57 10 2 9 2 1 10 9 11 2 0 0 7 0 9 1 10 9 2 1 10 9 11 2 12 9 2 3 13 10 9 1 10 9 0 9 2 3 1 10 9 1 15 10 9 13 3 2 1 10 9 2 1 10 9 1 11 2
24 10 9 7 9 1 10 9 2 15 13 13 15 1 10 9 0 2 3 13 13 1 10 11 2
50 1 10 9 1 10 9 1 10 9 2 10 9 1 9 1 10 11 13 3 1 10 11 2 13 1 10 11 2 10 9 0 1 13 12 0 9 1 9 1 11 7 13 1 10 9 12 9 1 9 2
35 10 9 1 10 11 13 16 10 9 13 13 1 10 9 1 10 9 1 10 9 0 2 10 9 15 1 10 9 2 3 13 10 9 2 2
30 10 9 1 10 9 13 1 10 9 1 9 0 0 1 10 9 1 10 9 1 10 0 9 1 10 9 1 10 9 2
44 3 2 10 9 1 10 9 1 9 2 13 1 10 11 2 13 16 10 9 1 9 1 9 1 10 11 13 3 0 2 1 15 13 13 1 12 9 1 12 1 12 1 12 2
24 1 12 9 2 10 9 13 13 12 12 9 1 9 2 12 9 1 9 2 2 13 10 9 2
56 13 16 10 9 15 13 3 1 10 9 0 1 10 9 7 3 13 10 9 1 10 9 1 10 9 2 9 13 2 1 13 13 15 1 15 13 1 10 9 3 2 15 13 10 12 12 9 1 9 2 12 9 1 9 2 2
24 10 9 0 13 15 1 10 9 0 1 2 9 0 2 2 1 15 15 13 9 1 9 13 2
22 1 12 1 3 2 13 12 9 1 15 15 13 10 9 1 9 0 1 12 12 9 2
25 10 9 13 10 9 13 1 12 12 9 2 13 10 9 1 10 9 1 12 2 1 12 12 9 2
4 0 13 9 0
51 10 11 2 11 2 11 2 2 13 1 11 2 1 10 11 2 13 3 10 9 13 13 12 9 1 2 10 9 2 1 10 11 7 13 10 9 1 9 1 10 9 2 1 10 9 1 10 9 0 2 2
42 1 10 9 13 1 9 0 2 10 11 2 13 10 9 1 10 0 9 2 13 1 9 0 7 0 2 7 2 13 1 9 10 9 13 1 12 1 9 1 12 2 2
35 10 11 13 10 10 2 9 0 2 1 10 9 1 10 11 2 11 2 11 2 7 13 10 2 9 0 1 10 9 0 1 10 9 2 2
61 13 10 0 1 10 0 9 1 9 1 12 9 1 9 1 12 9 15 10 11 13 1 10 9 1 9 2 11 13 0 1 10 9 1 10 9 15 13 2 1 10 9 2 3 13 1 10 9 0 2 7 3 1 10 0 9 1 15 15 13 2
58 10 9 2 15 13 10 9 1 11 2 13 1 13 10 9 1 12 9 2 13 9 7 13 10 9 1 10 9 2 3 10 9 13 13 2 16 2 1 10 9 2 13 1 13 15 1 0 9 1 9 7 10 9 15 13 1 9 2
21 13 3 1 13 1 10 9 1 10 10 9 1 9 2 13 15 3 13 1 9 2
28 1 10 9 2 10 9 13 0 1 13 2 13 1 10 9 13 9 7 13 10 9 1 13 3 10 10 9 2
16 13 12 9 1 9 1 10 9 2 1 10 9 1 10 9 2
26 1 10 9 1 9 10 2 9 1 2 9 2 2 2 1 10 9 1 10 9 2 13 1 0 9 2
1 11
5 3 12 9 1 11
38 10 9 1 9 7 10 9 1 10 0 12 9 1 10 11 2 1 9 1 11 2 13 3 13 1 10 9 1 15 13 9 1 10 9 1 10 11 2
16 10 11 2 15 2 13 3 3 7 1 15 9 1 10 9 2
15 15 13 0 13 2 13 13 2 13 10 9 1 10 11 2
11 13 10 9 2 13 13 3 15 13 3 2
6 15 3 3 13 0 2
8 15 13 1 10 0 9 0 2
14 9 1 10 11 13 2 9 0 1 10 9 2 1 9
6 9 1 13 1 10 11
15 13 10 9 1 10 9 1 9 13 10 9 1 10 11 2
67 10 9 13 3 2 15 13 9 1 10 9 13 1 10 2 9 0 1 10 9 2 7 15 13 10 9 3 0 1 10 9 1 0 2 13 10 9 1 10 9 1 9 1 9 1 10 11 7 10 9 1 10 9 1 2 9 2 7 1 10 9 0 1 0 7 0 2
11 10 9 13 3 10 9 13 7 3 13 2
56 10 11 13 13 13 1 10 9 2 11 2 10 9 1 10 9 1 13 10 9 2 3 0 2 3 0 1 12 9 2 2 1 10 9 1 10 9 1 10 9 7 13 15 1 13 4 13 2 15 9 3 2 1 10 9 2
63 2 10 9 1 10 9 2 12 2 1 10 9 1 15 3 10 11 13 13 13 3 0 16 10 0 9 13 9 15 13 0 1 13 1 10 0 9 1 9 2 3 13 10 9 1 9 0 7 9 1 9 1 10 11 2 2 13 11 2 1 10 11 2
30 2 3 10 9 15 13 2 2 13 3 2 2 10 9 13 10 9 1 13 13 1 10 9 1 9 2 1 10 9 2
16 10 9 13 2 1 11 2 1 10 9 1 13 1 10 9 2
59 10 11 2 15 3 15 13 13 1 15 13 2 1 13 9 1 9 2 2 13 16 10 9 1 10 9 1 9 0 1 10 9 13 3 3 0 1 10 0 7 0 9 15 13 2 3 0 2 16 10 9 0 3 13 3 1 10 9 2
1 11
5 10 9 1 10 9
18 13 12 9 1 10 11 16 10 10 9 0 13 2 10 9 0 2 2
22 13 12 9 2 13 3 13 10 9 15 15 13 3 0 9 1 10 11 1 10 0 2
13 2 3 13 13 1 10 9 2 2 2 13 11 2
16 13 2 3 2 12 1 10 9 3 13 1 10 9 1 12 2
19 1 10 9 1 12 9 2 13 10 11 1 13 13 10 11 1 10 11 2
6 13 9 1 10 9 2
14 1 9 2 13 1 10 9 13 9 2 13 3 9 2
43 9 1 16 13 1 9 1 10 11 2 1 10 9 1 2 9 13 2 1 10 9 1 10 9 1 11 2 2 3 15 15 13 1 10 9 1 10 9 1 10 13 11 2
26 13 3 13 10 9 1 10 9 1 10 9 0 3 13 1 10 9 1 10 9 2 11 7 11 11 2
31 10 9 1 10 9 1 10 11 13 3 9 0 10 11 2 15 3 13 13 2 9 2 15 13 13 10 9 1 10 9 2
28 3 13 2 3 2 10 9 1 13 10 9 1 10 9 1 12 9 2 15 1 15 1 3 12 9 1 9 2
16 10 9 13 3 13 1 10 9 11 1 10 9 1 9 0 2
38 15 13 13 13 9 2 3 1 15 13 13 10 9 1 9 1 9 0 2 1 10 9 13 2 1 10 9 1 12 12 9 2 13 3 1 10 9 2
43 2 13 0 16 15 15 13 2 2 13 10 9 1 10 9 2 1 10 9 15 3 1 10 9 13 9 1 10 11 2 1 10 11 2 7 15 15 13 4 1 13 3 2
32 13 1 10 2 9 2 13 1 10 9 1 9 7 13 1 9 13 1 10 0 9 1 15 12 1 10 9 15 13 1 13 2
23 10 2 1 9 2 13 1 10 9 7 1 10 9 1 10 12 9 1 10 2 9 2 2
42 0 13 10 9 1 10 2 9 2 15 13 13 1 12 9 7 1 10 2 9 2 13 3 1 10 9 7 3 1 10 9 1 10 9 2 3 13 9 1 10 9 2
44 3 2 3 2 10 9 7 9 13 9 1 10 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 7 11 2
54 1 10 9 2 1 10 9 3 0 2 13 9 1 10 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 7 11 2
9 10 9 1 9 2 2 9 2 2
15 9 2 10 9 13 15 7 3 13 2 3 2 10 9 2
27 3 2 15 15 15 13 2 1 13 10 9 7 10 10 9 2 13 16 10 9 1 10 11 13 3 0 2
40 10 9 1 9 3 13 13 2 1 3 2 15 3 2 16 1 10 9 13 10 9 15 13 10 9 1 10 9 2 10 9 1 11 2 1 10 9 0 0 2
7 13 13 10 9 1 9 2
24 9 2 7 3 10 11 13 1 13 10 9 1 7 1 9 2 1 10 0 9 1 10 9 2
12 9 0 1 9 1 10 9 11 13 9 7 9
4 11 1 10 9
33 13 13 7 13 1 10 9 0 9 2 10 9 11 13 3 13 7 15 3 13 10 9 15 13 10 9 1 10 11 2 10 9 2
13 1 10 9 2 1 10 9 3 10 9 13 13 2
10 1 10 9 2 10 9 1 11 13 2
17 1 13 10 9 11 2 2 3 13 1 10 9 1 10 9 2 2
31 10 11 1 10 11 2 10 10 9 1 9 13 1 10 11 2 13 15 3 1 10 11 13 1 10 9 1 10 13 9 2
14 9 2 10 11 2 11 2 3 13 13 10 9 3 2
26 2 13 1 12 9 1 15 13 1 13 9 0 15 13 10 9 0 1 10 9 2 2 13 10 9 2
49 11 2 10 9 0 2 13 13 1 13 10 9 0 1 10 9 7 13 2 13 2 10 10 9 7 13 1 9 1 10 9 2 7 2 3 3 1 13 2 1 15 3 11 13 13 10 9 2 2
16 11 2 9 2 13 2 3 0 2 10 9 13 1 10 9 2
30 2 10 9 3 15 13 1 13 1 0 9 1 10 9 1 10 9 1 10 0 9 2 9 7 13 2 2 13 11 2
6 11 13 9 1 10 11
38 10 11 13 13 3 2 1 9 1 10 9 2 10 3 9 2 1 10 13 9 2 1 10 9 11 2 11 2 1 10 0 9 1 10 2 11 2 2
30 10 9 0 13 3 1 13 10 9 1 10 9 2 15 13 4 13 1 9 1 10 9 1 9 13 1 13 10 9 2
38 1 10 9 1 10 11 2 10 9 13 13 1 10 11 7 10 11 13 10 9 3 1 13 2 2 3 13 15 13 16 10 9 3 15 13 9 2 2
15 10 9 1 10 9 13 3 13 1 10 9 1 10 9 2
36 16 15 3 13 1 13 15 2 10 11 13 13 10 9 3 10 11 13 1 13 10 9 15 13 10 9 1 13 1 11 7 3 1 10 11 2
8 11 1 10 11 7 1 10 11
10 10 2 9 2 2 1 10 9 0 2
22 10 0 9 2 0 1 10 9 2 10 9 0 7 0 2 13 1 9 12 9 13 2
14 13 3 2 13 15 15 15 13 10 9 3 3 0 2
21 1 10 9 15 15 13 2 10 9 0 2 1 10 9 2 10 9 1 10 9 2
6 11 7 11 1 9 2
1 11
2 1 11
8 1 11 2 11 2 11 7 11
34 2 3 13 10 9 0 2 3 2 13 10 9 2 2 13 1 10 11 10 9 0 1 10 11 1 13 10 9 1 10 2 0 2 2
30 2 11 2 11 7 11 13 10 9 15 13 2 2 13 2 1 3 13 16 11 3 13 13 15 2 16 13 13 15 2
2 1 11
27 10 9 1 10 0 1 10 11 2 2 10 9 0 1 10 9 2 2 3 13 13 10 0 9 1 9 2
31 11 13 10 9 1 10 9 2 11 2 1 11 2 7 1 10 9 1 11 2 10 9 1 10 9 1 11 2 1 11 2
5 9 0 1 9 0
4 10 9 1 11
32 10 9 1 10 9 0 1 9 1 10 9 0 1 9 0 2 1 9 1 10 9 0 2 13 1 4 13 1 10 9 0 2
23 3 2 1 10 11 2 13 15 3 10 9 13 1 12 9 1 9 1 13 7 9 0 2
21 1 11 2 9 1 10 11 2 10 9 13 13 10 9 1 9 1 10 0 9 2
9 1 11 2 3 11 13 13 10 9
3 2 11 2
23 10 12 9 15 13 1 9 2 13 11 2 13 10 0 9 2 13 9 0 1 10 9 2
19 10 9 1 10 9 13 1 10 9 2 13 9 3 13 11 13 10 9 2
46 13 13 10 2 9 1 10 11 2 2 10 9 13 16 13 1 10 2 9 0 2 2 1 10 9 2 7 13 16 15 2 13 13 13 1 10 9 0 7 13 1 10 9 0 2 2
14 1 3 1 13 10 9 1 10 0 9 13 10 9 2
34 10 9 1 10 9 1 10 9 2 13 11 2 2 13 0 1 10 9 7 1 10 9 2 7 2 0 9 2 1 13 1 10 9 2
42 2 13 0 13 9 3 0 2 1 13 13 2 16 9 3 0 15 2 3 2 3 13 0 2 2 13 2 13 2 10 9 2 1 15 10 9 13 13 1 10 11 2
11 3 13 16 10 0 2 13 13 3 2 2
41 1 11 2 10 9 3 13 10 9 1 10 9 1 9 1 10 11 2 1 10 9 0 15 13 1 10 9 1 12 9 2 1 10 11 1 13 1 10 12 9 2
10 1 11 2 10 9 0 13 12 9 2
53 12 10 9 15 15 13 2 1 9 2 1 10 0 9 1 10 9 1 10 9 13 10 9 2 11 2 13 1 10 9 7 1 10 9 1 10 9 2 7 11 2 10 9 13 9 1 10 9 0 1 10 9 2
59 9 0 2 0 13 7 9 1 10 9 1 9 1 10 11 2 11 13 1 10 9 10 9 1 10 9 0 7 1 10 11 2 15 13 1 13 1 15 15 13 1 10 9 1 10 9 1 10 9 2 3 11 3 13 13 10 10 9 2
19 7 2 13 3 3 10 9 0 2 3 13 10 9 13 16 11 13 13 2
29 1 10 9 1 10 9 2 1 0 9 0 7 1 12 9 0 2 10 9 1 10 11 3 13 1 10 12 9 2
15 3 2 1 12 1 9 13 10 10 9 1 12 0 9 2
31 7 2 1 10 9 1 10 9 2 13 13 1 13 7 13 2 1 13 7 1 13 10 2 9 2 7 10 2 9 2 2
1 9
18 13 1 10 11 2 1 11 2 1 10 9 2 10 11 7 10 11 2
23 0 1 10 9 1 1 10 0 9 12 2 1 9 1 9 2 1 10 9 1 10 9 2
18 10 2 11 2 3 13 10 0 1 9 1 10 0 9 0 7 0 2
48 9 0 1 15 13 10 11 1 10 9 15 13 13 2 10 9 7 9 1 10 9 1 10 9 2 2 1 16 10 15 2 13 1 9 1 10 9 0 1 9 7 9 1 10 9 0 2 2
35 1 3 2 10 9 3 13 13 1 10 9 2 1 13 1 10 0 9 1 2 9 2 3 13 7 10 15 3 13 13 1 9 3 13 2
7 9 2 11 13 1 10 11
34 10 9 0 9 2 11 2 13 3 16 10 9 0 9 11 13 13 12 9 1 9 2 3 12 9 1 9 2 1 10 9 0 11 2
24 10 9 13 9 1 10 9 9 2 7 3 15 1 10 9 13 1 10 9 13 10 9 13 2
35 10 11 3 13 13 10 10 9 1 10 9 1 10 9 1 10 9 1 10 11 2 10 0 9 13 10 9 3 0 1 10 9 0 11 2
8 9 2 11 3 0 1 10 11
56 11 2 1 11 2 9 1 10 11 2 11 2 1 0 2 13 3 10 9 3 0 1 10 9 1 10 12 9 1 9 1 10 11 2 0 1 10 11 7 9 0 7 2 11 2 11 1 9 2 9 15 10 9 15 13 2
30 11 13 10 0 9 1 9 2 13 10 10 0 9 1 10 9 1 10 11 1 10 11 2 9 11 2 2 13 1 9
19 1 10 9 1 12 9 2 11 2 2 11 2 11 2 13 15 1 9 2
13 13 15 1 10 9 3 10 0 2 7 13 13 2
4 1 10 9 2
69 1 10 9 1 9 13 1 10 9 3 2 11 2 2 2 1 15 2 3 13 13 12 2 2 2 10 9 1 10 9 0 1 10 9 1 10 11 1 13 2 10 9 1 9 1 10 2 9 1 10 0 9 2 2 3 13 1 11 2 1 10 9 11 2 7 10 15 2 2
4 7 10 9 2
34 10 0 9 2 3 2 13 13 10 9 1 13 1 11 2 1 12 12 9 1 10 2 9 1 10 9 1 10 9 2 2 1 12 2
24 1 10 9 13 10 0 9 1 9 7 10 9 1 10 9 15 13 1 13 1 10 10 9 2
6 2 13 9 11 2 2
9 16 13 15 10 9 1 10 9 2
8 2 6 2 15 3 13 15 2
22 15 3 13 1 13 2 2 15 2 1 10 9 3 15 13 2 13 13 10 0 9 2
14 13 15 13 16 10 9 13 1 10 10 9 2 9 2
6 13 15 1 10 9 2
28 15 13 9 0 2 16 10 9 13 15 15 3 15 13 1 10 10 9 2 1 10 10 9 1 13 10 9 2
33 13 2 1 10 10 9 1 13 2 16 10 9 1 9 2 15 15 13 1 13 9 3 0 2 12 1 10 0 9 1 10 9 2
35 3 13 9 10 3 10 9 13 3 1 10 9 2 0 1 13 1 4 13 2 13 2 1 10 9 1 13 1 4 13 1 10 10 9 2
24 15 15 13 1 10 10 9 2 1 3 9 2 1 7 1 9 2 3 13 9 1 10 9 2
27 7 15 15 3 13 1 10 9 2 3 13 2 1 15 15 13 1 13 2 16 13 1 15 15 15 13 2
20 3 13 9 10 15 13 10 9 0 2 15 15 15 13 16 15 13 7 13 2
16 13 0 2 13 15 9 2 13 1 9 10 9 1 10 10 2
47 3 3 3 2 13 15 9 2 9 1 15 10 2 9 2 13 4 13 1 10 9 1 9 2 3 13 10 9 1 10 9 7 10 9 0 2 3 13 3 3 10 9 1 10 9 0 2
19 1 10 10 9 2 11 13 10 9 3 0 2 12 0 9 1 10 10 2
15 3 15 13 13 16 10 9 13 10 10 9 1 10 15 2
18 13 15 10 10 9 1 9 2 7 15 1 15 10 9 13 1 9 2
12 13 10 9 0 1 10 9 0 15 15 13 2
26 10 9 3 13 1 10 9 16 13 9 1 10 10 2 7 1 10 10 9 2 7 1 10 10 9 2
30 15 13 15 13 10 2 9 1 10 9 2 2 7 3 15 13 1 10 10 0 9 2 15 13 13 1 10 10 9 2
23 3 13 9 10 1 15 10 9 2 10 9 2 10 9 2 10 9 7 10 9 13 13 2
21 7 2 3 2 10 10 9 13 0 1 15 13 10 9 2 10 9 2 10 9 2
10 16 11 13 9 0 2 0 7 0 2
12 13 10 0 1 9 2 15 1 9 1 9 2
14 3 2 13 10 0 2 15 15 13 2 15 15 13 2
22 1 10 9 2 13 3 0 3 13 9 13 2 2 0 2 2 1 9 7 9 0 2
4 15 13 15 2
38 13 10 9 1 10 9 0 2 7 13 15 1 9 2 1 9 0 2 1 10 9 15 3 13 13 15 15 15 13 2 3 15 13 2 15 15 13 2
55 1 10 9 2 10 11 13 10 10 0 9 2 11 2 7 10 9 11 2 9 15 13 13 10 9 1 10 11 1 10 9 2 13 1 10 9 1 2 9 2 2 13 1 10 9 7 1 10 9 1 2 9 2 2 2
52 1 10 9 1 10 11 2 11 2 2 10 11 13 4 1 13 11 2 11 2 2 13 1 10 10 11 2 7 11 2 11 2 2 13 1 9 2 15 13 9 0 1 9 1 9 13 1 11 1 10 9 2
38 1 10 9 2 3 13 3 12 9 1 10 1 15 9 2 3 3 12 1 12 12 9 13 10 9 1 9 1 9 2 9 1 9 2 9 7 9 2
49 10 10 9 2 3 2 1 10 9 1 10 11 2 13 10 9 1 10 11 1 13 10 9 3 0 1 10 9 1 10 9 1 2 9 2 13 1 11 2 13 1 11 11 2 9 0 1 11 2
64 1 15 15 10 11 13 2 10 9 15 13 13 10 9 0 1 10 9 1 13 15 1 10 9 1 10 11 1 10 9 0 13 3 1 13 1 10 9 1 10 0 9 1 10 9 1 10 9 2 7 15 3 1 10 9 1 13 2 9 0 1 9 2 2
19 3 2 1 10 0 9 10 11 13 13 10 9 1 9 1 9 7 9 2
37 13 10 9 1 10 9 0 1 10 9 1 9 2 15 13 1 3 12 9 1 12 1 15 0 12 2 15 13 3 0 9 1 9 1 10 9 2
64 3 10 9 1 10 9 0 13 10 9 1 10 11 1 13 2 3 1 10 13 9 1 2 9 2 11 2 10 9 1 9 0 2 3 10 1 10 9 1 10 11 2 1 10 11 7 1 10 11 2 15 9 12 1 10 0 9 2 3 2 1 10 11 2
48 13 3 10 9 1 13 1 10 9 0 1 10 9 1 11 2 1 10 9 1 10 0 9 1 10 9 2 2 1 15 15 10 9 13 13 12 9 1 9 2 1 10 9 13 1 10 9 2
9 11 13 13 10 9 1 2 9 2
46 10 11 2 11 2 13 13 1 10 10 9 2 1 10 0 9 2 13 1 12 1 9 2 1 16 13 10 9 1 2 9 2 2 1 13 10 9 1 9 1 10 9 1 10 9 2
33 1 10 10 9 2 10 9 11 2 2 13 0 9 1 10 11 2 2 1 15 15 13 10 10 9 2 1 9 2 1 10 9 2
5 11 2 1 10 11
8 9 2 9 7 9 1 9 2
19 2 3 3 3 13 13 16 10 9 1 10 9 13 4 13 1 9 0 2
27 10 9 3 10 9 15 13 13 0 7 15 1 15 13 13 16 10 9 0 3 13 0 2 2 13 11 2
44 2 7 15 15 15 13 13 16 2 3 13 2 3 2 10 9 15 13 1 10 9 7 15 3 13 13 1 10 9 0 15 10 9 3 15 13 2 13 0 13 15 10 9 2
9 7 3 15 13 3 1 9 0 2
12 13 0 9 15 13 13 10 9 1 9 2 2
13 10 9 13 16 3 13 9 15 13 10 10 9 2
36 2 10 9 15 15 13 3 13 2 15 13 10 10 9 1 9 0 2 13 10 9 1 0 9 2 15 3 13 13 10 9 2 2 13 11 2
43 2 13 3 9 15 13 10 9 1 9 2 3 10 0 2 7 13 3 9 1 2 9 2 9 2 15 10 9 13 1 13 10 9 2 3 13 9 1 10 9 1 9 2
25 7 13 0 13 10 9 13 1 10 9 1 10 9 0 2 15 13 10 9 1 9 0 2 2 2
12 10 9 13 1 4 13 3 1 11 7 11 2
11 10 0 9 13 16 10 9 1 10 9 2
57 3 2 13 15 10 9 1 10 9 1 10 9 7 1 10 10 9 2 13 1 10 9 13 2 13 7 3 2 3 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 7 9 2 3 11 2 11 2 11 2
34 1 10 0 12 9 2 10 9 13 13 9 1 9 1 9 2 3 1 9 0 2 2 9 0 1 9 7 9 2 16 13 3 9 0
25 2 10 9 12 2 9 1 12 2 13 3 2 9 11 2 2 13 10 0 9 13 1 10 9 2
11 15 12 2 9 1 12 2 13 11 2 2
33 10 9 13 15 1 10 2 9 2 2 9 1 11 7 11 2 15 13 10 9 1 9 0 3 10 9 0 1 10 9 13 13 2
67 1 9 2 13 15 9 2 15 10 9 1 10 9 13 3 13 2 13 7 13 2 1 10 9 7 3 1 11 7 11 2 11 2 11 2 11 2 11 2 11 2 11 2 10 9 2 0 2 1 11 2 9 1 9 0 1 11 2 11 2 11 2 11 2 11 2 3
53 13 15 13 0 13 1 10 9 3 13 7 0 2 11 7 11 13 13 10 9 1 10 9 1 15 10 2 11 7 11 7 13 1 16 10 9 13 1 10 9 0 1 12 1 15 2 1 10 9 1 10 0 2
38 3 13 7 13 10 0 9 1 10 9 2 1 15 12 1 15 12 2 13 1 12 7 12 2 2 1 10 0 9 1 11 2 11 2 11 7 11 2
39 11 7 11 13 9 1 15 10 9 1 9 7 9 7 1 10 11 7 10 9 0 13 3 0 2 11 2 11 2 11 2 9 0 1 11 7 11 2 2
45 11 2 13 10 9 1 15 15 13 10 10 9 1 10 9 7 9 1 10 2 9 2 2 1 9 1 11 7 9 1 11 2 11 2 11 7 11 2 7 10 13 9 1 11 2
49 7 2 3 2 11 2 15 13 10 9 1 10 10 2 9 2 2 13 10 9 3 0 2 3 12 9 13 1 9 13 2 3 10 9 7 10 9 13 0 2 7 10 9 0 15 13 3 0 2
33 10 9 13 15 1 10 0 9 7 10 9 1 10 9 13 12 1 10 9 1 13 2 1 13 1 10 11 10 10 9 2 11 2
25 10 0 13 16 2 11 13 10 9 15 13 13 1 10 9 7 15 13 10 9 1 10 9 13 2
17 13 10 9 0 2 1 9 9 2 0 7 0 1 13 9 2 2
38 1 10 9 1 9 13 1 11 2 11 13 16 10 9 0 1 11 13 13 9 1 10 9 1 10 0 9 2 1 10 9 1 15 13 10 10 9 2
25 10 9 2 10 9 2 0 15 13 1 10 9 13 10 9 0 1 10 9 1 9 7 1 9 2
43 10 9 1 10 9 2 1 10 9 2 1 10 9 1 10 9 0 2 13 10 10 9 1 10 9 2 1 10 9 1 13 10 9 0 15 13 1 10 9 10 9 0 2
43 0 1 10 9 1 9 0 1 11 2 11 13 10 2 11 2 1 11 1 10 0 9 0 2 10 9 2 1 10 10 9 0 2 13 3 10 9 1 9 0 7 0 2
43 1 10 9 1 11 2 11 2 11 2 10 9 3 13 3 13 1 0 9 2 3 1 0 9 1 10 9 0 7 13 2 0 7 0 2 0 1 10 0 9 1 9 2
52 10 9 1 10 10 0 9 13 4 13 2 3 1 10 11 2 1 11 2 9 3 13 4 13 2 1 9 1 10 9 1 9 2 10 9 0 2 10 9 13 10 9 1 10 9 1 10 9 1 10 9 2
49 13 15 2 1 10 9 11 2 15 13 10 9 2 1 10 9 0 2 0 1 13 2 1 10 9 0 2 10 9 13 1 10 0 9 1 9 13 1 9 1 10 11 2 11 2 11 7 11 2
30 1 10 9 1 9 2 10 9 1 10 10 9 2 1 10 9 1 10 9 0 2 13 13 1 13 9 2 13 11 2
38 16 10 9 1 10 9 2 3 9 2 13 13 3 0 1 10 11 2 1 10 9 13 13 10 9 13 13 10 0 9 1 10 9 1 10 0 9 2
36 7 3 3 10 9 0 3 13 1 10 9 1 13 10 9 0 2 1 15 2 13 16 15 15 13 13 1 13 10 9 1 10 9 1 9 2
24 16 10 11 13 1 10 9 1 10 9 13 3 0 16 15 13 9 1 12 0 9 1 9 2
20 7 13 16 13 13 3 0 1 10 0 2 7 15 13 10 10 9 1 9 2
2 9 13
15 10 9 1 9 1 11 3 13 15 2 7 3 10 9 2
31 11 13 10 9 7 10 9 1 10 9 2 10 9 11 13 1 9 7 10 9 11 7 11 13 10 9 2 7 3 3 2
31 10 10 9 0 13 15 1 10 9 1 10 9 1 10 9 1 9 1 10 9 2 15 3 13 1 10 9 1 10 9 2
19 11 13 12 1 10 9 15 15 13 0 7 3 15 13 3 10 9 13 2
10 3 3 1 9 2 13 10 9 0 2
3 9 1 9
3 11 1 11
65 10 9 2 11 2 13 3 3 1 11 2 3 13 1 10 11 2 1 11 2 11 2 2 1 13 9 1 10 9 0 1 10 11 1 10 9 1 10 11 15 15 13 1 12 1 9 1 11 2 3 13 13 10 9 13 10 9 1 10 9 1 9 1 11 2
26 1 10 9 9 2 10 9 13 3 12 9 1 1 10 11 2 11 7 11 2 13 3 1 12 9 2
27 3 15 13 16 10 9 1 10 9 0 7 13 1 10 9 0 13 13 10 9 1 10 9 1 10 9 2
34 10 9 3 13 3 10 9 1 10 9 1 0 1 10 9 0 13 9 2 9 2 2 3 3 13 1 10 9 1 0 9 1 9 2
24 10 9 13 13 16 10 9 13 3 1 9 13 1 10 11 2 15 13 10 9 1 15 12 2
9 9 1 10 11 13 1 12 1 9
5 11 3 13 9 13
24 10 11 2 11 2 13 1 13 15 1 10 9 1 10 9 1 9 2 7 3 3 13 9 2
31 10 9 13 3 2 1 10 9 1 10 9 2 7 1 0 9 2 16 15 13 10 9 3 13 1 10 11 7 10 11 2
27 16 3 15 13 10 9 1 0 9 2 13 0 16 10 11 13 10 9 0 1 10 12 9 1 10 11 2
32 2 10 9 13 2 3 2 16 10 9 3 13 4 13 1 10 9 1 9 0 2 2 13 11 2 9 1 11 1 10 11 2
23 3 2 10 9 1 11 3 13 1 12 9 1 13 10 9 0 1 15 15 13 0 13 2
13 7 10 9 1 10 11 1 10 9 13 3 0 2
19 11 13 9 1 10 0 9 1 9 2 3 1 10 9 1 10 9 0 2
48 16 10 9 1 10 11 13 13 3 12 9 1 10 9 13 2 13 15 10 9 15 13 1 9 10 9 0 1 10 10 9 2 15 13 1 12 12 9 1 9 2 3 12 9 1 9 2 2
26 11 13 16 10 9 13 13 0 9 1 10 11 1 10 9 7 10 9 1 10 9 0 1 10 9 2
19 10 9 13 2 1 10 0 9 1 10 9 2 1 10 9 1 10 9 2
22 2 10 9 3 13 4 13 1 10 9 0 2 2 13 10 9 1 10 11 2 11 2
15 2 10 9 1 10 9 7 1 10 3 9 3 13 0 2
8 10 3 9 13 13 9 2 2
26 10 9 13 1 10 9 1 2 3 2 10 11 2 13 10 9 15 13 13 3 10 9 1 10 9 2
28 1 11 7 1 10 11 10 9 3 13 0 2 7 1 10 10 9 1 10 11 3 13 2 16 1 9 0 2
16 10 9 0 13 13 10 9 1 2 9 2 0 0 7 0 2
28 13 15 2 3 2 10 0 9 1 10 9 1 12 1 9 1 10 9 2 7 9 2 7 9 1 10 11 2
16 7 3 1 9 2 1 2 9 0 2 1 13 10 3 0 2
8 3 10 11 13 13 10 9 2
7 7 15 13 13 10 9 2
22 9 7 9 2 1 10 9 2 11 2 2 1 10 9 2 1 10 11 2 1 11 2
10 1 11 2 13 13 10 11 2 11 2
40 2 11 2 15 13 9 1 10 11 7 1 10 11 2 13 1 10 11 1 10 9 1 13 1 10 9 1 10 10 12 0 9 2 0 9 1 10 11 2 2
57 11 13 1 11 2 15 13 13 1 10 9 11 2 10 9 1 10 10 9 1 10 11 7 2 3 1 10 9 1 10 9 2 13 1 15 1 10 9 1 10 9 2 13 1 9 1 10 9 7 1 10 9 1 10 11 2 2
38 2 13 16 10 11 13 10 9 2 13 0 9 2 7 13 3 16 10 11 2 1 15 15 13 1 10 9 2 13 3 0 1 10 9 16 10 11 2
21 10 9 1 10 11 13 3 0 16 10 9 13 15 3 3 3 1 10 9 2 2
31 10 9 13 1 10 9 1 11 2 11 2 7 13 2 1 10 2 9 1 11 2 11 2 11 2 11 2 11 7 11 2
9 9 1 10 9 1 9 1 11 2
10 1 10 9 1 10 11 2 1 11 2
9 0 1 10 9 1 12 1 9 2
2 9 0
4 11 2 1 11
28 13 13 1 12 1 9 1 10 9 1 9 0 2 3 10 9 1 10 10 9 13 13 1 10 9 1 11 2
23 1 9 1 10 0 9 2 15 1 10 9 1 10 9 0 13 13 13 1 10 10 9 2
3 11 13 3
24 3 12 9 13 1 9 1 3 1 10 0 9 1 10 11 2 15 15 13 1 12 1 9 2
104 1 10 9 13 9 9 3 2 11 2 2 1 10 9 11 2 11 2 2 2 11 2 2 1 11 2 13 10 0 9 2 9 2 0 2 2 11 2 2 1 11 2 11 2 2 2 11 2 2 1 10 9 11 2 2 11 2 2 1 11 2 11 2 2 2 11 2 2 1 10 9 11 2 2 11 2 2 1 10 9 11 2 2 11 2 2 1 10 9 11 2 7 2 11 2 2 1 10 9 11 2 1 10 2
55 1 10 11 7 10 11 2 10 9 1 10 9 13 13 1 10 9 11 2 11 2 2 11 2 11 2 2 11 2 11 2 2 11 2 11 2 2 11 2 11 2 2 1 10 9 0 7 1 10 9 1 10 9 0 2
38 10 9 13 3 10 9 1 10 9 0 0 2 9 1 9 1 10 9 11 2 10 9 1 10 9 0 11 7 10 0 9 0 1 10 9 1 11 2
38 1 13 10 11 1 10 9 1 13 2 3 1 10 9 1 10 9 1 10 9 2 13 4 13 10 9 1 9 1 10 9 0 7 12 9 1 9 2
23 3 13 13 15 13 10 9 0 2 7 15 13 10 9 1 10 9 0 0 1 10 9 2
46 1 10 9 15 13 9 10 9 1 15 10 9 1 10 9 13 13 2 10 9 11 2 13 16 10 9 3 3 13 13 2 7 16 2 10 9 13 13 10 9 0 1 10 11 2 2
18 9 2 13 13 13 10 9 1 10 9 0 2 3 10 11 13 13 2
23 9 2 1 3 2 10 9 1 10 11 1 10 9 13 4 13 1 13 10 0 9 0 2
23 10 9 1 15 13 13 13 1 10 9 10 9 15 3 13 1 10 9 1 10 0 9 2
12 3 13 9 1 13 2 3 2 10 10 9 2
22 13 10 9 0 7 0 2 9 1 9 0 7 9 0 1 13 9 2 9 2 9 2
50 1 10 9 0 2 13 1 10 11 7 3 2 13 2 13 15 1 13 9 1 10 9 1 10 9 7 9 2 10 9 15 13 13 7 15 15 13 1 13 13 10 0 0 1 10 9 1 0 9 2
45 3 1 13 13 12 0 9 7 10 10 9 1 9 0 2 13 16 10 9 3 0 15 13 13 2 13 2 1 10 9 1 11 2 13 10 9 2 13 15 0 7 0 1 13 2
50 13 3 3 1 15 2 1 10 9 1 10 9 1 11 1 10 9 1 10 9 1 10 9 1 10 9 12 2 1 10 9 1 13 9 1 13 3 2 1 9 7 9 1 13 10 9 1 10 11 2
45 1 10 9 1 11 2 13 3 1 13 10 9 1 11 2 1 10 9 15 13 13 10 9 2 3 13 3 7 3 2 7 15 13 1 13 7 1 13 1 13 10 9 13 15 2
9 12 1 10 0 9 13 10 9 2
20 15 13 15 13 16 10 15 13 9 1 10 9 7 10 9 2 1 10 9 2
25 13 16 15 15 13 13 0 7 0 2 3 1 15 13 13 2 7 16 10 10 9 13 3 13 2
20 1 10 9 2 13 9 1 10 0 2 1 15 13 13 10 9 1 10 9 2
21 3 2 3 2 10 9 0 7 0 3 15 13 1 10 9 0 2 1 10 9 2
8 1 12 2 13 1 9 0 2
21 13 9 2 13 1 13 9 2 13 0 1 13 7 1 13 9 0 1 10 15 2
1 11
4 10 9 1 9
37 10 9 1 10 9 1 9 1 9 2 15 13 13 3 12 9 1 9 2 13 12 1 10 9 1 13 1 10 0 9 1 9 0 1 10 9 2
44 3 1 10 9 2 15 13 3 9 0 2 10 9 0 13 13 10 9 1 9 1 15 1 10 9 2 1 12 0 9 1 9 2 9 1 9 2 2 9 2 13 7 9 2
28 1 10 9 1 10 9 7 1 10 9 0 1 10 9 3 15 13 9 2 10 9 0 13 3 13 10 9 2
30 3 2 13 10 9 3 13 15 13 10 9 1 0 9 0 1 10 0 9 1 9 3 9 1 9 7 9 1 9 2
75 13 15 3 16 2 1 9 1 12 2 3 10 11 13 10 0 9 3 0 1 3 2 13 10 9 11 2 13 1 10 11 2 1 10 9 1 11 2 12 9 1 9 1 11 2 2 1 15 13 13 12 12 9 1 9 2 3 13 15 13 1 10 9 1 12 9 13 9 1 10 9 1 9 0 2
48 10 11 2 15 13 1 9 10 0 9 1 9 0 0 0 1 9 2 13 13 10 9 1 10 9 3 10 9 1 2 9 2 13 3 13 2 16 15 13 10 9 0 1 9 1 10 9 2
46 16 10 0 9 1 10 9 15 13 13 1 10 9 1 10 9 13 2 1 10 9 0 10 9 13 16 15 13 4 3 13 2 13 2 3 2 10 9 1 15 13 9 0 1 9 2
38 3 2 15 15 13 13 3 10 0 9 1 10 9 13 13 2 1 10 9 1 10 9 2 9 15 13 1 13 3 0 10 9 1 10 0 9 0 2
13 10 9 13 3 10 9 1 11 1 10 0 11 2
35 13 15 1 10 11 2 11 13 10 9 1 9 1 10 9 2 2 13 3 10 9 1 9 1 2 13 9 3 13 3 4 1 13 2 2
31 3 1 10 9 1 10 9 13 15 16 15 13 0 1 2 13 15 15 13 1 10 9 7 3 13 16 13 1 9 2 2
44 1 10 9 1 9 1 2 9 2 2 10 9 1 9 1 9 2 10 9 1 9 0 2 10 9 1 9 7 10 9 3 2 10 11 13 10 0 9 1 2 13 10 9 2
80 13 10 9 13 3 9 1 11 1 15 13 10 9 2 1 15 10 2 3 1 10 9 10 1 10 9 13 1 13 11 2 10 13 9 1 9 2 11 2 1 10 9 0 2 7 10 9 7 9 0 1 11 2 10 9 1 11 2 13 3 9 1 13 10 9 15 13 1 10 9 1 10 0 9 1 10 9 2 11 2
58 10 9 13 15 2 3 2 1 10 9 1 10 9 7 13 16 10 9 0 2 0 1 10 9 0 3 1 10 9 1 10 9 2 13 1 13 10 9 0 15 3 15 13 2 3 15 13 2 3 15 13 1 10 9 0 7 0 2
26 7 10 9 15 13 13 1 10 9 1 10 9 1 9 1 10 15 13 9 1 10 9 1 10 9 2
12 2 13 10 9 1 9 7 9 1 10 11 2
58 11 13 10 11 1 13 9 0 1 10 11 2 10 9 13 1 10 11 1 12 2 1 10 9 1 10 11 2 7 1 13 10 9 1 9 1 10 9 13 1 10 9 0 2 16 15 13 10 10 9 1 10 9 0 1 10 9 2
26 1 15 2 10 11 0 13 1 3 10 9 1 10 9 1 10 9 1 10 9 1 10 12 9 0 2
24 2 10 9 0 13 10 0 9 1 13 10 9 1 10 11 7 10 11 2 2 13 9 11 2
23 7 10 9 1 10 9 0 13 13 1 10 0 1 10 11 3 12 9 1 2 9 2 2
44 15 16 10 9 1 10 9 0 13 10 9 0 1 10 11 2 15 13 1 10 9 13 13 10 10 9 1 9 1 10 11 2 11 2 2 15 13 13 1 10 9 1 9 2
26 10 9 1 10 9 13 13 10 9 13 10 9 13 2 7 13 1 10 9 1 9 1 10 12 9 2
48 10 9 1 10 11 2 15 13 3 12 0 2 13 1 12 2 3 10 9 1 10 0 11 13 10 9 1 10 9 2 15 2 1 10 0 9 2 13 13 9 7 15 13 3 1 10 9 2
23 1 10 11 2 10 9 0 1 13 10 9 1 10 9 1 9 13 11 2 11 7 11 2
21 7 10 9 13 3 13 1 10 2 9 2 0 2 13 1 11 2 11 7 11 2
17 1 11 2 12 12 9 2 2 10 9 13 11 2 11 7 11 2
22 1 3 2 13 10 0 9 1 10 9 9 11 1 10 2 9 2 0 1 10 11 2
18 1 10 9 0 1 10 9 0 2 3 12 13 3 7 15 13 13 2
29 10 9 0 11 13 1 10 9 11 1 12 2 12 2 12 2 7 11 13 13 1 10 9 11 1 12 2 12 2
9 3 2 10 9 3 15 13 3 2
44 1 13 16 10 2 9 2 13 1 10 9 2 10 9 13 3 13 10 0 11 2 3 13 11 2 10 9 1 11 2 7 3 3 13 10 9 1 10 9 7 10 9 0 2
33 1 10 9 15 10 9 13 3 1 13 1 10 9 2 10 9 1 10 9 0 13 2 1 9 2 10 9 1 15 3 15 13 2
15 1 13 3 10 9 3 13 2 3 2 1 10 0 11 2
25 10 0 9 13 3 3 0 1 13 7 2 13 10 9 2 16 13 10 1 10 9 3 3 3 2
4 11 13 13 9
44 10 9 11 2 9 1 10 9 2 13 15 3 1 10 9 1 10 9 13 3 0 7 1 15 2 7 1 10 13 9 2 13 1 10 11 10 9 1 10 9 1 10 9 2
16 10 11 13 13 10 9 1 10 9 15 3 13 13 1 11 2
37 10 9 13 3 2 1 10 9 2 1 10 9 7 13 13 10 10 9 1 10 9 1 10 9 1 10 9 2 13 3 10 9 1 10 0 9 2
39 3 12 9 13 13 3 1 10 9 0 1 11 2 1 10 9 1 0 9 7 10 9 2 3 3 1 9 1 10 7 15 13 13 1 10 9 3 0 2
62 10 0 9 1 15 13 9 13 1 10 9 1 11 2 1 10 9 0 1 10 0 9 0 2 3 3 12 9 13 1 10 9 1 13 1 10 9 1 10 9 1 10 10 9 2 11 2 3 1 10 0 12 9 13 1 12 7 12 9 1 9 2
9 13 1 10 11 2 11 13 0 2
19 2 3 13 10 11 1 13 10 9 7 3 13 15 1 13 1 15 2 2
13 7 2 1 9 2 13 1 10 10 9 2 11 2
28 10 9 1 11 13 15 1 10 9 1 10 11 2 1 12 1 9 1 12 2 15 13 10 9 1 10 11 2
15 9 15 13 13 1 10 9 2 1 9 1 10 9 12 2
19 11 2 1 10 9 2 13 13 9 1 16 10 9 13 0 7 13 15 2
20 2 13 0 13 16 10 9 1 10 9 1 10 11 13 13 13 10 9 2 2
32 7 13 10 9 1 15 13 2 10 9 1 10 11 7 10 10 9 2 1 3 9 1 10 11 13 1 10 9 1 10 9 2
4 2 11 2 2
9 9 0 2 3 10 9 15 13 2
7 7 11 13 1 13 9 2
17 2 13 10 9 15 13 1 13 1 10 9 2 2 13 10 9 2
12 13 15 16 10 9 15 13 3 1 10 9 2
4 2 9 2 2
5 13 15 10 9 2
4 13 1 15 2
51 11 2 11 2 7 11 2 11 2 13 10 9 2 15 0 2 15 0 2 15 13 1 11 16 11 2 9 2 13 16 13 13 1 10 11 9 15 15 13 10 9 1 15 11 13 10 9 1 9 0 2
35 1 10 9 2 10 9 13 1 10 0 9 2 11 2 11 2 2 10 9 2 10 10 9 2 11 2 11 2 2 7 10 9 2 11 2
4 10 9 1 11
32 1 10 9 2 10 11 13 10 11 13 3 15 13 13 1 15 2 9 0 2 13 10 9 0 2 10 9 0 2 10 9 2
8 7 15 13 3 1 10 9 2
47 10 9 1 0 9 13 3 1 10 9 1 9 1 10 9 1 9 2 3 0 7 0 13 2 7 13 1 10 9 1 10 9 1 2 9 2 2 9 2 1 10 11 7 1 15 11 2
32 1 10 12 9 2 10 2 9 1 10 11 2 13 10 9 7 13 15 1 10 9 1 2 13 15 10 9 1 10 9 2 2
16 1 10 2 0 2 2 10 11 13 0 1 13 12 0 9 2
37 13 0 10 0 9 1 9 1 10 9 1 13 10 0 9 0 1 12 9 1 10 9 1 10 11 15 15 13 13 12 9 1 10 9 0 0 2
23 10 9 7 10 9 13 3 1 12 7 12 9 1 15 12 7 12 13 1 10 9 0 2
6 11 13 9 1 10 11
3 13 10 9
23 10 9 13 4 13 10 9 1 9 1 9 1 10 9 1 9 7 9 1 10 9 0 2
31 10 9 13 13 3 10 9 7 10 9 1 10 9 1 9 2 1 16 10 9 13 13 1 9 1 10 9 1 9 0 2
24 13 10 9 3 3 1 10 9 1 10 10 0 11 2 3 10 9 13 3 2 7 13 9 2
14 3 13 0 13 10 9 0 7 10 9 13 0 9 2
7 3 1 11 2 15 13 2
29 9 2 9 1 10 9 1 9 2 9 15 13 0 1 15 13 7 10 9 3 15 3 13 9 1 10 10 9 2
2 9 0
8 12 13 1 10 11 1 10 11
30 10 9 13 2 1 10 9 1 3 2 15 3 16 12 9 1 10 11 2 1 11 2 1 10 9 1 10 9 0 2
19 10 9 0 2 15 13 9 1 10 9 2 13 13 9 1 9 1 9 2
67 1 12 1 10 9 2 10 9 13 12 9 2 10 9 1 12 9 2 10 9 1 12 7 12 9 1 9 1 12 2 7 12 9 2 15 13 1 12 9 2 10 9 1 12 7 12 9 1 12 2 2 3 1 10 10 9 2 13 4 3 13 10 0 9 1 9 2
20 12 5 1 10 9 13 13 1 9 0 7 0 1 10 11 1 11 7 11 2
15 10 10 9 13 1 9 1 9 3 11 2 11 7 11 2
54 10 2 11 2 2 9 2 11 7 11 2 13 10 9 1 10 9 1 10 11 2 3 13 1 12 9 2 12 9 2 1 10 2 9 1 10 9 2 2 11 2 11 2 11 2 11 7 11 2 3 13 13 2 2
21 1 13 1 10 9 1 10 9 0 1 10 9 1 10 11 2 10 9 15 13 2
28 13 0 13 9 1 9 0 2 3 10 9 2 13 3 1 9 0 2 13 13 1 13 9 1 10 10 9 2
12 3 13 10 9 13 1 10 9 1 10 9 2
21 2 15 13 10 9 0 1 13 9 2 2 13 1 10 11 11 2 1 10 11 2
35 2 1 10 9 2 10 9 1 10 9 13 13 15 1 13 10 9 1 10 9 1 10 9 1 10 9 2 13 10 9 1 10 9 2 2
25 10 11 13 3 16 10 9 1 10 11 7 10 11 1 10 9 1 10 9 0 3 13 3 13 2
17 10 9 1 10 9 9 1 10 11 13 13 12 1 10 0 9 2
43 10 11 13 4 1 13 10 9 0 1 10 9 1 9 2 16 0 1 12 9 2 7 2 3 2 10 11 13 13 2 3 2 10 10 9 1 10 9 0 1 10 11 2
27 3 2 10 9 1 10 11 13 13 2 1 12 9 0 2 1 10 11 2 1 10 11 7 1 10 11 2
53 10 9 13 3 2 9 2 1 10 9 1 9 0 1 10 9 2 15 13 13 3 2 2 1 13 13 1 10 9 1 10 9 1 10 9 13 1 13 10 9 1 9 0 2 1 13 10 0 9 1 10 9 2
13 11 13 10 9 1 9 1 11 1 12 1 12 2
27 3 2 1 10 9 2 13 1 10 9 1 11 2 13 1 13 10 9 0 2 3 1 10 9 1 9 2
14 13 13 1 10 9 3 3 0 2 10 0 9 11 2
18 10 9 13 15 10 9 2 13 4 13 9 1 10 11 1 10 11 2
6 1 12 13 1 11 2
24 13 15 1 10 10 9 11 2 3 15 10 9 9 15 3 13 13 1 10 9 1 10 9 2
15 11 13 15 1 10 0 9 1 10 9 1 10 9 13 2
23 1 10 9 0 2 11 13 1 10 10 9 0 3 1 13 1 11 2 1 13 1 11 2
20 12 1 10 9 13 1 10 9 13 10 9 1 9 0 1 10 9 1 11 2
48 1 10 9 0 13 2 3 2 15 13 10 9 1 2 9 2 1 10 9 1 11 1 10 11 1 11 1 10 9 1 13 10 0 9 13 1 10 0 9 1 9 2 0 2 1 10 11 2
63 1 13 13 1 10 11 1 11 10 3 0 9 1 9 1 9 1 11 2 10 11 0 3 13 1 10 9 1 10 9 0 2 15 13 10 0 9 1 3 13 13 10 9 2 3 10 9 1 10 9 2 11 2 13 1 10 11 7 3 13 1 11 2
2 9 13
45 3 2 3 12 9 3 1 10 9 3 1 10 0 9 1 9 1 10 9 2 15 13 10 0 9 1 9 1 10 9 7 10 9 2 13 13 13 1 13 10 9 1 10 9 2
26 10 9 13 1 10 9 2 13 1 10 9 1 10 9 1 10 9 1 10 9 3 13 13 0 9 2
35 7 3 10 9 0 13 1 9 1 9 0 2 13 10 9 7 13 9 1 10 9 1 10 10 9 1 9 2 13 10 9 1 10 11 2
31 10 9 1 10 9 13 16 2 1 10 9 1 10 9 2 10 9 13 1 13 3 1 10 9 2 13 9 1 10 9 2
43 12 1 10 9 3 13 9 1 10 11 2 13 16 10 9 0 13 3 13 2 16 10 9 13 13 7 16 10 9 1 10 9 13 4 4 13 1 10 9 1 10 9 2
38 2 3 13 2 9 2 1 10 9 2 2 13 10 9 2 15 13 16 10 9 1 10 9 1 10 9 1 10 9 1 10 9 13 4 4 3 13 2
29 7 13 3 10 11 1 3 13 13 1 10 0 9 1 10 11 2 1 13 16 10 9 15 13 1 10 0 11 2
43 10 9 13 10 0 9 3 1 10 9 1 10 9 2 10 9 15 13 2 3 2 1 13 9 1 10 9 1 10 9 13 10 0 3 13 1 16 2 3 13 9 2 2
87 1 10 0 1 10 9 2 10 9 15 13 13 1 10 9 15 13 1 13 1 15 13 1 11 2 13 1 10 0 9 1 9 2 13 2 9 2 7 15 13 16 15 13 1 10 9 2 1 10 9 0 1 12 2 12 2 0 9 7 0 9 2 13 10 10 9 1 9 0 2 9 13 2 2 2 1 15 15 13 10 9 1 10 9 1 13 2
37 1 0 1 10 9 2 13 13 10 9 1 2 10 9 13 3 1 11 2 3 13 1 10 9 1 10 9 1 10 9 2 1 9 1 9 2 2
7 1 9 2 15 13 13 2
49 3 2 3 13 11 2 9 1 10 11 2 2 3 3 13 13 10 9 1 10 9 1 13 1 10 9 2 3 3 15 13 15 13 9 1 9 2 10 9 0 1 10 9 3 3 13 13 2 2
24 3 2 1 10 9 13 3 13 10 9 1 10 9 1 9 1 9 2 16 13 13 15 2 2
47 11 3 13 9 1 16 15 13 1 2 10 9 13 1 10 9 0 1 10 9 1 13 10 9 2 3 13 1 10 9 2 1 13 2 1 13 13 3 16 13 10 9 1 13 9 2 2
5 11 13 0 9 0
9 12 9 1 10 9 1 10 9 0
33 12 1 10 9 1 11 1 10 9 1 10 11 1 10 11 2 11 2 13 13 10 9 0 2 13 10 9 15 10 11 3 13 2
23 13 15 1 10 9 1 10 9 1 12 9 1 10 9 1 10 9 0 1 10 9 0 2
7 0 9 1 9 1 10 11
4 11 13 13 9
37 10 11 2 10 0 9 0 0 1 9 1 10 11 2 13 13 13 1 13 10 9 1 9 1 13 10 10 9 1 12 12 9 1 10 9 12 2
42 10 9 13 3 13 1 10 11 2 15 13 9 1 10 11 7 1 10 11 7 13 1 12 12 9 1 9 13 1 12 9 1 9 2 1 9 0 1 12 12 9 2
8 13 1 10 9 1 9 13 2
17 1 12 9 2 13 15 1 15 1 15 2 13 15 3 10 9 2
3 10 9 2
6 7 3 13 10 9 2
24 1 10 9 1 15 13 1 10 9 0 1 10 11 13 2 1 10 9 0 2 10 9 9 2
11 13 15 7 10 9 13 1 13 1 9 2
12 13 3 10 2 11 2 2 1 10 10 9 2
17 13 15 10 9 1 10 9 2 7 3 3 13 15 15 0 13 2
13 15 10 13 15 3 2 7 13 15 1 13 3 2
82 3 0 1 10 10 9 1 9 2 1 0 9 1 10 9 0 2 10 9 1 10 11 13 12 9 3 1 10 9 13 1 10 11 7 10 11 1 10 9 0 1 10 9 1 10 9 0 1 12 2 7 12 9 3 1 10 9 1 10 10 2 11 2 2 10 0 9 2 2 10 9 15 13 1 10 11 10 0 9 1 13 2
51 11 13 10 9 15 13 10 9 2 15 13 10 9 1 10 9 0 1 10 9 2 1 10 0 9 1 9 2 1 12 2 1 10 9 15 13 3 12 12 9 1 9 7 13 12 9 1 9 1 9 2
27 1 10 10 9 1 9 1 9 0 2 3 13 10 9 1 10 11 2 10 9 0 13 1 13 10 9 2
64 13 10 9 1 10 9 1 10 9 1 10 9 1 10 9 0 1 11 2 1 10 11 2 2 1 10 11 1 10 9 1 10 0 9 1 9 11 2 7 1 10 11 1 13 10 9 1 0 9 1 10 9 1 10 2 9 2 13 9 7 9 1 9 2
39 1 10 11 2 13 10 2 9 2 11 1 10 9 7 9 1 9 1 9 0 2 9 1 9 7 1 9 2 3 1 10 9 0 7 1 9 1 9 2
27 13 3 10 0 9 13 1 10 9 0 9 11 1 13 9 0 1 10 9 0 15 10 9 13 1 13 2
52 1 9 1 11 2 1 10 11 2 10 10 9 1 9 7 9 0 13 0 7 2 1 10 11 1 10 9 2 10 0 9 1 10 0 9 0 1 9 2 1 12 12 9 2 2 13 10 9 1 10 9 2
30 10 11 13 1 13 10 9 1 10 0 9 2 10 11 2 1 10 9 1 9 1 10 0 9 1 2 9 2 0 2
37 10 0 9 13 1 9 2 9 0 7 9 1 10 9 1 10 10 9 0 1 10 9 1 10 9 2 9 2 9 0 2 9 7 9 1 9 2
58 2 13 10 9 9 1 13 10 9 1 10 11 1 10 9 1 10 2 9 2 2 2 13 1 10 9 2 11 2 11 2 9 2 15 13 13 16 2 10 9 1 10 9 1 10 2 9 2 13 10 9 1 10 0 12 9 2 2
45 9 0 1 10 9 13 10 9 1 10 9 0 7 1 10 9 3 15 15 2 3 2 13 13 10 0 9 2 13 15 3 10 9 7 10 9 0 7 2 3 2 10 9 0 2
14 10 11 13 3 3 10 9 1 9 0 1 12 9 2
35 10 9 13 1 10 11 13 1 10 9 2 7 10 9 2 0 2 13 13 3 2 15 13 3 12 9 1 10 9 13 13 1 10 9 2
27 1 10 9 3 3 13 13 2 10 11 13 1 12 9 7 1 10 9 0 1 12 9 1 10 9 11 2
21 10 9 1 10 9 3 13 3 13 16 13 10 9 13 10 9 0 1 12 9 2
32 3 2 10 9 1 10 9 1 11 13 10 9 1 10 9 13 7 13 0 9 1 10 0 9 2 15 13 10 9 1 11 2
18 10 9 0 13 1 13 10 9 1 10 9 1 11 1 10 9 9 2
24 10 11 13 10 9 1 10 9 2 7 10 9 1 10 11 13 3 1 13 15 1 10 9 2
35 7 10 9 0 3 13 0 9 7 13 13 10 9 2 16 3 13 13 1 10 9 1 3 13 13 9 2 15 13 10 9 1 10 9 2
53 2 1 10 9 2 13 3 15 1 13 2 2 13 11 2 15 13 10 10 2 9 0 2 1 16 2 10 9 1 9 1 10 9 0 7 10 9 0 2 13 1 13 10 2 9 2 1 10 11 1 10 11 2
7 11 13 1 10 10 9 2
13 2 13 1 13 10 9 1 10 0 9 7 9 2
29 1 11 2 3 2 10 0 9 7 10 9 13 10 10 9 2 7 2 3 2 3 13 10 9 0 2 2 13 2
39 1 13 10 9 13 1 9 1 9 1 10 11 2 11 13 2 10 9 1 9 0 2 2 15 13 15 1 13 1 9 13 1 10 0 9 1 10 9 2
38 1 10 9 0 2 10 9 13 0 7 1 9 2 1 11 7 10 11 2 1 10 9 0 10 9 13 3 1 10 9 10 0 9 3 1 10 9 2
14 9 0 2 10 9 1 15 2 10 9 3 1 9 2
25 11 2 15 13 10 9 13 10 0 9 0 7 3 15 13 10 9 1 10 10 1 10 9 0 2
28 2 1 10 9 13 1 10 9 13 16 3 13 3 15 2 2 13 15 10 9 15 13 10 9 1 9 0 2
22 10 9 0 11 13 15 0 1 10 9 1 10 11 2 15 13 2 9 7 9 2 2
38 10 9 13 3 16 10 2 10 11 13 2 3 2 1 13 13 3 10 9 15 13 10 9 0 0 15 13 10 9 1 9 1 9 1 10 9 2 2
22 15 16 10 9 1 10 11 1 10 9 13 13 1 10 9 0 1 10 9 2 11 2
50 2 3 13 10 9 1 10 9 2 11 2 13 3 10 9 2 7 10 9 1 9 9 7 1 10 11 2 7 3 10 9 0 1 10 9 0 1 10 9 0 1 10 9 2 2 13 10 9 0 2
26 1 11 2 3 15 13 1 10 9 1 9 2 7 3 1 10 9 3 10 11 13 1 13 10 9 2
25 2 3 10 9 1 10 9 7 1 10 9 3 13 1 10 9 3 10 11 13 10 9 0 2 2
2 11 2
2 11 2
10 9 1 9 1 10 9 1 10 9 2
12 9 2 7 9 2 1 10 9 1 10 9 2
54 10 9 1 0 9 2 1 15 10 9 0 13 9 1 10 9 1 9 0 2 13 10 9 1 10 9 1 9 1 10 9 1 10 11 2 13 10 9 3 9 1 9 2 1 10 9 15 13 3 1 11 15 13 2
45 1 10 0 9 2 11 13 10 9 9 1 0 9 2 3 10 9 1 13 10 9 1 10 9 15 13 2 3 1 10 9 15 13 13 10 9 15 10 9 1 10 9 3 13 2
11 3 13 15 15 13 10 9 2 11 2 2
1 9
31 3 15 2 13 3 13 10 9 0 0 15 13 4 13 1 10 11 2 9 1 10 11 2 13 9 1 10 9 1 9 2
52 11 2 9 1 10 11 2 11 2 1 10 9 1 10 9 2 13 1 10 9 9 0 1 10 9 1 10 9 2 13 7 1 10 9 13 1 9 15 13 13 1 11 7 1 10 2 9 1 10 9 2 2
2 9 0
34 10 9 1 10 9 1 10 11 1 10 11 2 3 13 3 7 9 2 13 13 10 9 1 10 0 9 1 11 1 10 10 0 9 2
36 10 9 15 15 13 1 10 12 9 3 13 1 10 9 15 13 2 7 13 1 13 2 15 15 13 2 13 9 2 7 15 13 13 1 3 2
30 1 9 2 7 1 10 9 1 10 9 0 2 0 7 0 1 10 9 1 10 9 2 3 2 7 1 10 0 3 2
18 13 15 15 3 13 2 3 1 10 0 9 1 9 13 1 10 9 2
28 9 2 10 9 13 10 9 1 9 1 15 13 7 13 1 10 11 2 3 10 9 15 13 4 13 7 13 2
20 16 13 10 9 2 10 11 13 13 10 9 2 15 13 13 3 10 10 9 2
26 13 0 16 15 13 10 9 13 16 13 0 1 10 11 7 1 10 9 13 10 9 16 3 13 15 2
70 10 9 1 9 1 10 11 9 7 9 2 11 2 10 9 2 7 11 2 10 9 2 13 15 3 0 1 10 2 11 2 15 13 15 13 7 13 10 9 1 10 9 2 3 1 10 9 0 2 11 2 13 10 9 1 10 9 0 2 15 15 13 1 10 9 1 9 7 9 2
6 11 2 12 2 12 9
1 11
2 1 11
8 1 11 2 11 2 11 2 11
31 10 9 13 16 10 9 13 3 9 1 13 0 9 1 9 7 13 10 11 1 13 10 10 9 1 10 9 1 10 9 2
23 2 10 11 3 15 13 13 1 10 0 9 0 1 10 9 1 9 2 2 13 10 9 2
33 10 9 1 10 11 2 11 2 1 15 13 10 10 9 1 10 9 13 16 15 13 13 16 10 9 1 9 15 13 1 0 9 2
26 2 10 9 3 13 10 9 3 13 0 13 1 13 10 9 7 15 3 13 0 13 2 2 13 11 2
23 2 10 11 13 1 10 9 7 3 13 9 1 16 13 13 1 9 15 3 3 0 2 2
3 10 9 13
33 0 1 10 0 9 1 10 9 15 13 1 13 9 1 9 1 13 10 10 9 2 3 3 13 0 0 1 2 13 2 13 2 2
39 3 3 7 1 10 9 0 2 10 9 13 1 13 16 10 9 1 10 9 13 4 13 1 16 13 13 10 9 1 10 2 3 9 0 2 1 15 13 2
62 10 9 1 9 2 1 10 10 0 9 2 1 15 3 1 10 10 9 2 13 3 10 9 1 13 13 1 10 9 2 1 15 15 13 16 13 3 13 1 10 11 10 0 9 1 9 15 13 10 9 1 10 9 1 9 2 1 9 7 1 9 2
17 11 7 11 13 1 9 2 13 9 2 9 2 13 7 10 9 2
19 10 0 13 10 9 1 10 9 13 16 3 15 13 7 16 3 13 13 2
40 3 3 12 0 9 2 13 9 7 9 1 10 9 1 10 9 2 13 10 11 2 3 13 1 10 11 2 3 13 10 0 1 10 9 2 13 1 10 11 2
23 10 9 1 10 9 3 13 4 13 7 10 9 9 13 13 2 1 9 2 1 10 9 2
9 2 13 16 10 9 13 3 0 2
30 1 10 9 2 10 0 9 13 4 10 10 9 0 7 4 10 10 9 2 2 13 1 10 11 11 2 1 10 11 2
5 12 9 1 9 2
3 11 9 0
25 11 2 10 11 0 1 12 9 2 13 13 7 13 3 1 13 13 3 12 9 1 9 1 9 2
40 13 15 13 1 10 9 0 2 9 1 9 7 0 1 9 2 7 2 3 1 13 16 10 10 2 9 2 15 13 0 9 3 7 9 2 13 1 13 9 2
43 13 16 2 15 3 16 10 0 13 15 13 4 13 2 2 11 13 16 13 13 10 9 0 1 9 1 9 2 9 1 10 9 7 1 10 9 0 1 9 1 10 9 2
32 2 13 13 10 9 1 10 9 7 3 10 2 9 2 0 3 10 0 2 15 13 10 9 9 1 9 7 1 9 0 2 2
32 9 15 13 10 9 1 13 9 1 13 3 1 3 13 13 3 2 2 15 3 13 0 1 15 2 3 3 1 10 11 2 2
27 0 1 13 15 13 10 0 9 2 2 16 13 10 9 0 2 2 2 11 13 1 10 9 1 10 9 2
35 0 13 16 13 10 9 15 13 10 9 1 10 9 7 15 13 13 9 3 13 1 10 9 2 2 9 7 10 9 13 1 10 9 2 2
22 11 13 16 10 9 13 4 13 1 10 9 13 15 13 10 11 7 2 9 0 2 2
15 7 3 13 1 10 9 2 1 10 9 1 10 9 2 2
60 10 9 0 1 12 9 1 9 0 1 9 11 2 12 9 1 9 2 12 9 2 10 9 1 9 0 11 2 10 9 0 11 2 10 9 1 9 2 10 9 1 9 11 7 10 9 1 12 9 2 13 10 9 13 1 10 9 1 9 2
18 10 9 2 3 1 13 1 10 11 1 11 2 13 13 1 10 11 2
46 1 13 1 11 2 13 1 11 7 1 11 2 13 10 10 9 1 9 0 1 9 1 9 0 2 15 13 1 4 13 1 11 2 3 13 1 13 9 1 10 9 3 13 3 0 2
42 1 10 11 13 13 2 10 11 13 1 13 10 9 1 10 9 1 10 9 3 1 10 10 9 0 15 2 16 3 13 10 9 3 0 1 10 9 3 2 11 2 2
24 3 2 1 10 10 9 1 9 15 15 13 2 13 10 9 0 1 10 9 1 10 9 0 2
38 10 9 13 15 2 1 13 3 10 9 0 2 3 10 9 13 10 9 13 2 1 15 10 9 1 11 2 11 7 11 13 13 10 2 9 2 0 2
18 2 11 2 13 9 1 10 10 9 2 15 13 2 1 10 9 0 2
57 10 9 1 10 9 3 0 1 10 9 1 11 1 11 13 13 10 9 2 0 2 1 10 10 9 2 3 10 9 1 10 11 1 10 9 1 9 7 2 9 2 3 13 4 13 10 9 1 10 9 1 10 10 9 3 0 2
43 13 10 9 3 13 1 9 1 9 2 15 2 3 2 15 13 0 2 13 15 3 1 10 9 0 2 15 13 1 10 10 0 9 10 9 2 15 15 13 1 10 9 2
66 10 9 13 0 7 0 2 13 1 9 0 1 10 9 3 0 1 11 2 11 2 0 1 9 1 9 7 9 1 9 0 2 15 1 10 9 0 1 10 0 9 3 13 3 16 10 9 2 7 15 13 10 10 9 0 7 0 9 2 1 10 9 1 10 9 2
7 3 12 9 1 9 7 9
21 10 11 13 3 12 9 1 10 9 0 1 9 2 13 3 10 9 1 10 11 2
26 2 13 15 1 0 2 13 1 10 10 9 2 2 13 11 2 2 10 9 1 9 1 10 10 9 2
18 3 15 3 15 13 1 10 9 1 10 9 0 2 2 1 10 11 2
21 2 13 13 16 15 13 13 10 9 1 10 9 15 13 3 1 10 9 0 2 2
43 12 0 9 13 15 15 13 10 0 1 9 2 13 2 7 0 2 1 10 10 9 1 10 9 2 1 10 9 2 1 10 2 0 2 2 1 10 9 2 1 10 9 2
18 1 10 9 2 11 13 13 10 9 1 15 13 1 4 13 10 11 2
56 2 13 1 10 9 1 15 13 10 9 2 10 9 7 10 9 1 10 9 7 1 0 9 1 10 9 1 10 9 1 10 9 15 1 10 10 0 9 3 15 13 1 15 15 13 10 9 0 15 10 9 13 13 13 2 2
34 11 2 15 13 1 13 10 9 1 10 9 2 13 3 10 10 9 1 16 10 11 13 2 10 0 9 1 10 9 1 10 11 2 2
3 2 13 2
42 2 13 13 9 1 10 9 7 1 10 9 1 10 10 9 2 1 10 10 9 7 1 10 10 9 0 1 9 0 15 15 13 1 13 7 1 13 13 1 13 2 2
4 10 9 1 9
63 10 9 1 13 1 10 9 0 1 10 9 0 1 10 11 10 9 13 1 10 9 2 16 3 1 10 9 15 15 13 3 1 10 11 2 13 3 12 9 7 10 0 9 13 1 3 3 13 1 0 9 2 13 1 10 11 7 1 11 10 9 13 2
31 15 13 1 10 9 2 1 12 2 1 13 10 3 3 13 11 2 7 11 2 3 13 3 13 2 13 13 3 12 9 2
47 12 2 1 10 9 0 2 11 2 3 9 13 1 10 11 2 2 10 9 1 10 11 13 12 9 2 13 10 0 9 1 10 11 2 7 13 2 3 2 10 0 9 2 1 10 11 2
10 11 2 11 7 11 13 1 10 9 2
15 10 0 9 13 13 10 9 1 10 0 9 1 10 9 2
54 3 2 10 9 13 13 1 10 9 1 10 9 1 10 9 13 1 10 9 1 10 9 1 9 1 10 9 3 15 13 13 10 9 2 10 9 3 0 2 2 7 13 10 9 1 10 9 1 10 9 1 9 0 2
20 1 10 9 12 1 9 2 10 9 13 1 10 2 9 2 1 10 9 0 2
28 12 9 3 11 13 15 1 10 9 1 10 9 0 1 13 1 10 9 1 9 2 9 2 9 7 9 2 2
26 1 10 9 0 2 10 9 13 4 13 2 13 4 13 10 9 1 3 12 9 1 9 1 10 9 2
46 1 10 9 2 13 13 10 9 1 9 0 1 12 9 1 9 0 2 10 9 2 10 9 1 9 7 10 9 0 1 10 9 1 10 9 0 1 12 9 2 9 2 12 9 2 2
6 2 9 2 1 10 9
32 2 13 10 9 3 13 2 3 0 7 3 13 2 2 13 1 10 11 11 2 15 13 0 1 15 15 15 13 1 10 9 2
44 1 10 9 3 1 10 9 2 15 13 2 1 10 9 2 10 9 1 10 11 7 10 9 0 1 0 9 2 3 10 9 1 9 2 0 7 0 2 10 9 7 10 9 2
24 10 9 15 13 13 1 9 2 7 15 11 3 13 9 1 13 1 2 9 1 9 0 2 2
19 2 15 13 10 9 1 9 2 3 0 7 0 1 10 9 2 2 13 2
21 10 11 13 13 16 13 9 1 9 1 11 7 11 2 15 15 3 13 7 13 2
36 2 10 10 9 3 13 0 2 3 13 0 1 10 10 9 13 15 2 13 13 3 13 0 7 1 9 10 9 3 10 9 13 2 2 13 2
15 10 9 13 2 1 10 10 9 2 16 10 9 13 0 2
2 9 2
30 2 3 2 10 9 0 2 3 0 2 15 2 13 1 10 9 15 3 3 13 2 2 13 15 1 10 9 1 9 2
54 10 9 1 10 9 0 2 3 13 1 9 0 2 15 13 3 10 9 1 10 0 2 3 2 11 2 7 2 11 2 2 13 3 0 2 16 10 9 2 16 3 15 13 1 10 9 0 3 0 2 13 3 0 2
21 10 9 1 10 2 9 2 7 10 2 9 2 13 10 9 0 15 3 15 13 2
12 2 13 13 1 10 9 1 10 9 7 13 2
19 7 15 13 1 10 9 13 15 1 10 9 1 13 1 10 9 1 9 2
11 7 3 3 13 9 15 13 10 9 0 2
5 3 15 1 9 2
11 2 2 9 12 2 13 13 10 9 0 2
9 3 2 13 10 9 2 3 0 2
14 2 15 13 13 10 9 0 2 7 10 9 15 13 2
16 15 13 10 15 1 10 9 0 2 7 10 10 9 15 13 2
20 15 13 10 10 9 2 13 15 2 0 1 13 10 9 2 2 9 12 2 2
16 7 2 3 2 10 9 13 13 7 13 10 9 1 10 9 2
21 2 2 3 10 9 13 13 2 3 13 3 3 1 10 9 16 10 9 13 0 2
13 1 10 9 15 13 9 1 9 2 2 13 15 2
8 7 15 13 1 10 9 13 2
19 10 9 13 1 10 9 1 10 9 2 1 15 13 10 9 1 10 9 2
18 7 10 9 13 9 7 3 9 2 2 13 15 2 2 9 12 2 2
27 10 9 2 3 2 13 3 13 1 10 11 2 15 9 13 10 10 0 0 2 1 10 9 1 12 9 2
31 10 2 9 11 2 2 1 15 13 12 9 0 7 10 9 2 13 12 1 10 9 1 9 2 13 10 9 1 10 9 2
23 10 11 13 3 10 0 9 1 10 9 15 13 10 9 7 15 13 10 9 1 10 11 2
26 10 9 1 10 9 3 13 15 7 10 11 13 16 10 9 1 11 13 1 9 1 9 1 10 11 2
39 10 9 13 3 13 13 1 10 9 13 10 9 1 10 11 2 7 10 11 2 11 2 13 1 13 10 9 3 13 13 15 1 9 1 13 1 10 9 2
5 9 2 13 2 9
42 12 9 0 2 10 11 2 11 2 11 2 7 10 11 2 11 2 2 13 10 9 1 9 1 9 1 9 0 15 13 1 10 9 1 10 9 9 13 2 11 2 2
31 10 9 13 2 1 10 10 9 2 10 9 1 10 0 9 1 9 0 1 10 9 2 1 13 1 10 0 9 1 9 2
32 10 11 13 15 2 3 2 13 15 1 10 9 1 10 9 0 7 13 9 0 1 9 7 9 1 10 9 1 10 12 9 2
16 3 10 2 9 1 10 9 2 3 1 10 9 7 9 2 2
83 2 2 2 1 12 2 1 10 11 2 10 9 0 13 10 9 13 2 11 2 1 15 13 1 10 9 1 10 2 9 13 1 10 9 2 1 10 9 7 1 10 9 2 2 2 10 2 9 7 9 0 2 2 15 13 1 13 10 9 0 2 0 2 0 2 2 0 16 13 1 10 0 9 1 9 2 13 1 9 7 9 2 2
23 7 13 16 2 3 15 13 13 1 10 9 1 10 9 0 1 10 9 1 10 9 2 2
38 1 3 1 3 2 10 9 13 4 1 13 10 9 2 13 3 1 10 9 0 13 1 10 9 1 9 2 1 15 10 9 13 10 9 1 10 9 2
28 3 2 10 9 1 10 9 1 9 13 1 10 9 13 16 3 13 1 0 10 9 0 2 15 1 10 11 2
38 13 12 10 0 9 0 2 10 9 1 9 13 1 10 9 1 9 2 10 9 1 10 9 1 11 13 9 7 9 2 7 3 10 9 1 10 11 2
35 10 9 1 10 9 0 2 11 2 13 3 2 9 1 10 9 1 9 2 2 13 16 10 9 13 2 1 12 9 2 7 3 1 9 2
59 1 10 9 1 3 2 1 11 2 11 13 13 13 10 9 0 1 13 10 9 1 10 9 1 10 11 1 10 9 0 1 10 11 7 1 10 9 1 9 2 7 11 3 13 3 2 3 3 13 9 1 9 1 10 12 12 9 0 2
49 10 9 1 10 11 13 3 10 9 1 10 9 2 13 1 12 1 9 2 1 16 12 12 9 13 13 1 11 2 16 13 3 16 11 13 10 10 9 1 10 2 9 0 2 1 10 12 9 2
14 11 13 16 10 9 13 9 1 9 7 3 1 9 2
9 10 9 1 10 9 1 11 13 11
40 10 9 1 11 2 15 13 10 9 11 2 13 12 9 2 10 9 1 10 10 9 7 10 9 1 10 10 9 1 12 9 1 10 9 11 2 9 1 11 2
19 3 1 10 9 2 11 2 3 3 13 10 15 2 2 13 10 10 9 2
4 11 1 10 9
33 11 9 13 3 13 10 9 0 2 13 10 9 0 2 10 0 9 2 12 5 2 1 10 9 13 10 11 13 1 10 9 11 2
8 13 9 2 3 2 10 9 2
21 3 3 16 1 10 9 1 10 9 2 10 9 1 10 11 13 2 3 2 13 2
13 7 11 7 10 9 3 13 10 9 1 15 13 2
13 15 15 13 9 2 7 3 3 13 15 13 13 2
16 15 1 10 9 1 10 0 9 13 1 10 9 1 10 11 2
6 2 11 2 13 1 11
17 1 10 0 9 12 2 2 11 2 13 4 13 1 10 9 0 2
14 10 9 13 3 1 10 9 13 1 10 11 1 11 2
21 1 15 2 10 9 1 10 9 0 11 1 10 9 1 10 12 9 13 4 13 2
4 11 13 0 9
23 2 11 2 13 10 9 1 10 0 9 0 15 13 9 2 1 10 9 2 1 10 11 2
14 1 10 9 1 11 2 10 9 13 9 0 1 11 2
11 10 9 1 10 0 0 13 13 1 11 2
22 10 9 15 13 1 10 12 9 1 10 9 2 13 1 9 2 9 2 9 7 9 2
21 2 13 10 9 1 10 11 2 2 13 10 9 11 2 13 9 1 10 9 2 2
15 1 11 2 11 7 11 2 10 9 13 13 3 1 11 2
23 10 9 2 15 13 4 15 13 3 1 10 9 2 13 10 12 9 1 9 1 10 9 2
17 1 10 9 1 10 9 1 10 9 2 13 10 9 13 10 9 2
10 9 1 10 9 0 3 13 10 9 2
16 10 9 11 2 1 10 11 2 13 13 1 11 1 9 12 2
13 10 9 1 9 1 10 9 0 13 1 9 12 2
14 10 9 13 13 3 9 1 10 9 1 10 9 0 2
21 9 1 10 9 1 10 9 1 10 11 13 13 1 10 9 1 10 9 7 9 2
31 1 10 9 2 10 0 9 2 11 2 13 10 9 1 9 0 1 13 10 9 1 10 9 1 13 10 11 1 9 0 2
28 10 9 1 9 1 10 11 2 11 2 13 3 16 10 9 2 11 3 13 13 10 9 16 3 13 9 10 2
14 10 9 0 1 10 9 13 1 10 11 9 12 9 2
28 16 3 13 9 1 9 7 9 1 10 9 1 9 2 10 9 13 13 1 10 9 1 9 1 9 1 9 2
38 3 2 1 10 9 1 10 9 1 13 1 10 9 0 2 10 9 13 1 10 9 10 9 1 10 9 2 13 1 9 12 9 10 9 1 10 11 2
25 10 9 13 10 9 1 9 1 10 9 0 7 10 0 9 13 1 3 13 9 1 10 0 9 2
35 13 15 15 13 2 13 2 2 3 2 15 13 1 10 9 0 1 12 9 2 11 2 10 9 7 9 1 9 0 7 0 1 9 0 2
4 11 2 3 2
7 3 3 13 15 13 3 2
14 15 13 10 9 16 13 15 13 10 9 1 10 11 2
9 15 3 3 13 16 3 13 3 2
15 11 2 7 15 10 9 13 1 10 9 1 10 9 0 2
5 11 2 10 9 2
16 3 12 9 13 13 10 10 0 2 3 10 9 13 3 12 2
18 10 9 13 13 10 9 1 10 9 1 10 9 7 13 10 10 0 2
15 16 15 13 10 9 2 13 9 0 7 13 10 9 0 2
19 10 11 7 10 11 13 13 1 9 1 10 9 7 1 10 10 10 9 2
24 10 9 1 10 9 15 13 9 1 10 9 13 3 13 4 13 3 1 10 9 1 10 9 2
23 10 9 1 10 11 2 11 2 12 2 13 16 13 13 9 9 1 10 9 1 9 3 2
28 11 13 3 16 10 9 13 13 2 9 0 1 13 13 1 10 9 7 9 1 10 9 2 0 1 10 9 2
24 2 10 11 13 13 1 10 9 1 10 11 7 1 10 11 2 1 10 11 2 2 13 11 2
25 11 2 9 1 10 9 2 13 16 10 11 2 15 13 1 10 11 1 9 7 13 3 3 2 2
21 10 11 2 10 9 12 9 2 1 9 12 2 13 10 9 3 0 1 10 11 2
9 10 0 1 9 13 9 12 12 2
40 10 9 1 10 9 1 9 15 13 13 3 1 10 9 1 10 11 2 1 10 0 9 12 13 13 1 10 11 2 15 3 13 9 1 9 1 10 9 0 2
22 2 1 10 9 2 3 13 10 9 2 13 16 4 13 10 9 2 1 3 13 13 2
15 3 3 3 13 10 9 1 13 10 9 2 2 13 9 2
5 11 11 2 9 2
5 11 13 1 10 11
31 10 9 1 10 11 13 10 0 2 11 2 2 1 15 11 13 10 9 1 9 0 15 13 1 10 9 1 13 10 9 2
23 1 10 0 9 2 11 2 12 2 10 2 11 2 2 10 9 13 10 9 1 12 9 2
16 11 3 13 1 10 9 10 9 1 13 1 10 9 1 9 2
11 15 12 13 9 1 12 1 9 1 12 2
5 10 9 1 10 11
43 13 3 3 1 15 15 15 13 10 9 1 10 0 9 1 10 11 3 12 9 3 1 10 9 15 2 1 10 9 1 10 9 2 13 10 9 11 1 10 0 9 0 2
41 1 10 9 2 10 12 9 3 13 1 13 10 9 1 11 2 10 11 2 10 11 7 10 11 2 13 13 10 10 9 1 9 1 9 2 3 2 1 12 9 2
28 11 13 13 10 9 11 1 10 10 9 7 2 1 15 2 13 10 10 9 0 2 13 10 9 1 9 0 2
29 10 11 13 12 1 10 9 15 13 1 10 9 13 1 10 0 11 2 1 12 1 9 1 0 1 9 1 11 2
24 9 1 9 0 1 0 1 10 11 2 11 7 11 13 13 1 11 2 1 10 11 1 11 2
7 10 9 13 10 9 0 2
29 12 1 10 0 13 11 2 15 13 3 12 9 2 1 12 9 15 13 1 13 10 2 9 2 1 0 1 0 2
20 3 9 2 15 13 13 10 9 0 1 10 9 0 2 15 13 1 9 0 2
17 11 13 1 10 3 0 9 1 10 9 1 10 9 1 10 9 2
9 10 9 13 9 10 1 10 9 2
36 9 1 9 7 9 2 3 11 2 11 2 11 7 11 2 13 10 10 7 0 9 16 11 7 15 15 15 13 13 1 9 1 13 3 9 2
8 3 15 13 10 9 1 15 2
4 9 2 11 2
18 13 16 3 13 13 9 0 7 9 1 9 1 10 9 13 1 11 2
15 13 16 10 9 1 9 2 3 2 13 10 9 1 11 2
4 13 10 9 2
9 1 10 9 2 10 9 3 13 2
12 11 3 15 13 1 10 9 1 9 7 9 2
20 10 10 9 0 13 16 11 13 1 13 3 2 3 15 13 1 12 9 0 2
30 7 10 11 7 10 9 13 9 0 1 13 10 9 1 10 9 1 10 9 1 11 2 15 13 10 9 13 1 9 2
17 10 9 1 10 9 13 10 9 13 13 10 9 2 1 10 9 2
15 1 10 9 2 10 9 1 10 9 13 13 1 10 9 2
14 2 10 0 9 1 10 9 1 10 11 3 13 0 2
20 13 10 9 2 2 13 10 9 11 2 12 2 0 9 1 10 9 1 9 2
10 2 13 11 1 10 12 9 1 9 2
14 10 9 1 10 9 13 13 9 3 2 2 13 11 2
23 1 13 10 9 1 12 9 1 9 2 10 11 3 13 3 16 10 10 9 13 3 3 2
17 10 9 1 10 9 13 9 1 10 9 1 10 9 7 10 9 2
8 2 3 13 13 9 1 9 2
31 7 13 9 15 13 4 13 1 10 9 1 13 10 9 2 2 13 11 2 9 1 10 11 2 15 13 10 9 1 9 2
7 9 13 3 10 9 1 9
19 10 9 15 13 10 9 0 1 9 3 13 13 0 9 1 10 9 12 2
24 10 0 9 1 10 11 2 11 2 13 9 1 12 5 1 10 9 13 1 10 9 1 0 2
31 11 2 15 13 10 9 1 10 0 9 1 10 9 2 11 2 2 1 10 11 2 13 10 9 1 10 9 1 10 9 2
23 1 15 2 10 9 1 10 9 1 10 9 7 1 10 12 0 9 1 9 3 13 9 2
2 9 0
2 0 9
29 11 2 10 9 2 15 13 9 1 10 9 1 10 12 9 1 9 1 10 9 0 2 13 12 9 1 0 9 2
14 13 13 9 13 2 13 9 2 9 2 9 7 9 2
19 1 9 1 9 1 10 9 1 10 9 2 9 1 10 9 1 10 9 2
5 1 12 1 9 2
12 9 1 10 9 2 1 9 12 1 9 12 2
36 10 9 1 10 9 1 10 9 0 7 1 10 9 1 9 7 9 13 10 0 9 1 13 10 9 3 13 1 10 2 9 1 10 9 2 2
71 3 15 13 3 1 10 9 1 10 9 3 13 13 9 0 1 10 9 0 2 3 1 15 13 13 10 0 9 0 1 10 9 7 9 1 10 0 2 7 3 3 1 10 9 1 10 9 13 13 7 13 10 9 1 10 9 0 15 10 9 0 13 13 1 15 13 0 1 10 9 2
23 10 9 13 15 1 10 9 1 13 7 13 10 9 1 9 2 9 7 9 1 10 0 2
28 15 13 16 13 15 16 10 9 13 0 1 9 15 10 0 9 13 2 3 13 10 9 0 1 13 15 13 2
23 7 2 3 2 10 15 15 10 9 13 3 13 1 4 13 1 9 15 13 10 9 0 2
31 3 10 0 9 1 15 13 10 9 13 10 9 13 1 9 1 9 7 2 3 2 10 9 0 13 13 10 9 1 9 2
32 13 3 3 0 16 13 0 13 3 1 10 9 1 10 9 0 1 13 13 1 9 1 15 15 13 13 0 1 10 9 13 2
28 1 10 0 9 1 3 13 1 13 10 9 1 10 11 2 1 12 9 2 10 9 13 10 9 1 10 9 2
20 3 2 10 9 13 15 13 3 1 10 9 1 10 9 3 11 2 11 2 2
1 9
22 12 9 0 2 1 3 12 9 10 2 13 13 1 9 0 1 10 9 1 10 9 2
12 15 13 13 1 9 1 12 9 1 12 9 2
16 10 9 2 0 1 10 9 2 13 13 3 1 9 1 9 2
10 9 13 16 10 9 13 13 0 0 2
1 11
33 10 9 1 9 1 10 9 11 2 1 9 1 12 2 13 9 1 10 9 1 9 12 9 2 1 10 9 1 11 2 11 2 2
16 10 9 13 4 13 1 9 2 9 2 9 1 9 7 9 2
26 10 9 13 15 16 10 9 1 10 13 1 10 11 2 7 0 16 15 9 13 2 1 9 12 9 2
4 9 1 10 11
26 9 7 9 1 9 13 13 1 0 9 1 11 1 10 9 1 10 9 1 3 2 1 10 9 0 2
12 9 1 9 13 1 3 12 9 1 10 11 2
15 13 1 10 9 13 7 10 0 13 10 9 15 13 9 2
38 1 13 10 0 9 2 10 9 1 10 11 13 1 10 9 16 13 16 3 13 1 9 10 0 9 15 13 10 10 9 1 15 13 2 3 16 3 2
23 16 10 9 13 1 10 9 0 2 10 9 13 13 16 10 9 13 9 0 2 13 15 2
29 3 10 9 1 13 10 9 13 9 3 1 10 9 15 13 10 9 2 10 9 1 11 13 13 10 9 1 9 2
24 3 13 15 10 9 13 7 3 13 15 10 9 2 1 9 13 2 1 10 9 0 7 0 2
20 10 9 13 10 11 2 15 13 9 1 9 0 2 1 16 10 9 13 9 2
15 10 9 13 13 1 9 7 9 2 15 13 13 15 0 2
3 13 10 9
24 10 9 0 13 16 10 9 3 13 3 2 13 13 9 0 1 9 1 9 1 15 13 2 2
2 1 9
14 1 11 2 1 10 11 2 1 10 9 7 10 9 2
14 2 13 16 13 3 7 13 3 2 16 9 13 2 2
17 9 1 10 11 0 15 13 1 9 7 9 1 11 2 11 2 2
4 13 10 0 11
6 13 9 7 10 9 2
6 9 1 10 9 12 2
35 10 9 0 1 9 13 10 9 1 10 9 1 11 2 13 9 1 15 1 10 9 2 2 9 1 9 1 10 11 7 9 1 10 9 2
13 10 9 0 2 15 13 1 10 11 2 3 13 2
5 9 1 15 12 2
11 11 13 10 9 1 10 11 1 10 9 0
14 11 13 1 10 9 1 11 2 16 15 13 13 3 3
21 3 3 2 10 9 15 3 13 1 10 9 2 13 1 10 9 1 10 9 0 2
15 15 15 13 2 13 9 1 9 1 10 9 1 10 11 2
12 11 13 1 10 9 1 10 9 1 10 9 2
5 2 15 13 3 2
13 15 15 13 1 10 11 13 10 0 2 2 13 2
15 11 13 10 9 1 10 9 2 3 13 13 1 10 9 2
11 11 13 16 10 11 3 13 10 10 9 2
15 11 13 9 1 10 9 1 12 9 2 11 2 1 11 2
53 10 0 9 0 1 10 11 1 12 9 13 9 3 2 3 10 9 11 13 1 10 9 10 9 3 13 11 2 15 13 13 12 9 1 12 9 1 10 9 1 13 0 9 0 7 0 1 10 9 1 10 9 2
12 10 9 0 1 10 9 13 11 2 11 2 2
24 15 13 13 1 10 11 7 1 10 11 2 1 15 1 10 0 9 0 1 9 0 7 0 2
31 10 9 13 3 1 10 9 0 1 11 2 1 10 11 2 9 0 1 10 9 2 1 10 9 0 2 9 1 11 2 2
12 10 9 0 1 10 9 13 1 9 12 9 2
13 10 0 9 1 10 9 13 1 13 10 9 13 2
39 1 10 11 2 3 10 9 1 10 9 1 10 9 13 1 9 1 0 7 0 9 3 2 3 13 1 13 16 10 9 13 9 1 10 9 1 10 9 2
13 10 9 1 9 13 1 10 9 13 13 1 9 2
31 2 10 9 1 9 0 13 10 9 13 9 2 2 13 10 9 1 11 1 10 11 2 11 2 9 1 9 1 10 11 2
33 2 3 13 1 9 1 9 2 7 15 13 10 9 0 2 2 13 3 10 9 2 1 9 1 10 9 1 9 2 1 10 11 2
24 11 13 10 9 0 1 12 2 1 10 11 2 9 1 15 13 10 0 9 1 10 9 0 2
8 9 13 1 9 7 9 13 13
40 10 11 2 12 9 1 9 1 11 2 13 3 1 10 9 10 9 0 11 2 12 2 13 1 13 1 10 9 10 9 11 2 12 2 1 10 9 1 9 2
13 10 9 11 2 12 2 13 16 11 13 10 9 2
33 11 13 13 1 11 1 13 15 13 1 10 9 13 2 9 1 15 13 10 9 1 10 11 1 10 9 11 2 3 10 9 13 2
31 2 10 9 1 10 9 13 9 1 10 9 7 2 3 2 1 10 9 1 9 15 11 13 13 1 11 2 2 13 11 2
27 11 13 16 13 13 10 9 1 10 0 9 2 15 13 3 1 10 9 15 9 1 15 13 1 10 9 2
7 2 13 10 9 0 0 2
14 10 0 9 1 10 9 3 13 0 3 1 10 9 2
13 13 3 2 3 13 13 10 9 13 2 2 13 2
10 15 13 13 9 7 9 1 10 9 2
19 1 10 9 2 13 10 0 9 13 3 3 1 9 1 9 1 13 13 2
23 10 9 13 13 1 13 10 9 15 13 3 1 13 1 9 13 1 10 9 1 10 9 2
6 13 9 1 0 9 0
33 9 0 7 0 1 9 13 1 10 9 1 9 0 15 3 13 1 10 9 1 10 9 2 13 10 9 1 10 11 2 11 2 2
9 2 13 10 9 1 10 0 9 2
19 13 15 3 13 10 9 0 1 10 9 1 10 9 2 2 13 10 9 2
31 10 9 0 1 10 9 13 10 9 1 10 0 9 1 10 9 3 1 10 9 0 2 15 13 13 1 10 9 15 13 2
10 11 3 13 3 10 9 1 10 9 2
18 2 10 9 1 10 11 13 0 2 2 13 3 3 1 13 1 11 2
6 10 9 0 3 13 2
22 7 13 9 1 13 16 2 1 10 12 9 2 3 13 10 10 9 1 13 10 9 2
23 10 0 9 13 13 10 9 1 10 9 0 1 10 9 1 9 1 10 9 1 10 10 2
24 15 13 13 10 9 1 9 15 13 13 9 1 13 15 1 10 9 15 13 1 15 1 15 2
52 3 2 10 9 1 10 11 1 10 11 13 10 9 7 10 9 1 13 10 9 2 15 2 1 15 15 13 1 10 11 11 2 13 1 10 11 2 7 10 9 2 0 2 15 13 1 10 9 0 7 13 2
18 10 0 9 1 10 9 1 0 9 13 1 10 9 1 10 9 0 2
38 1 10 9 2 13 13 3 10 10 9 0 7 0 13 1 10 9 1 10 9 1 10 9 2 1 9 0 2 9 7 9 13 1 10 10 9 9 2
10 9 1 13 2 13 2 1 10 9 12
25 11 2 9 1 10 11 2 11 2 2 13 16 10 9 1 13 13 1 10 9 1 9 1 12 2
17 2 1 12 13 10 0 9 1 9 2 7 3 0 2 2 13 2
14 1 15 2 3 10 9 1 9 0 13 0 7 0 2
6 11 13 1 13 1 9
16 10 11 13 1 13 9 1 10 9 1 10 9 2 11 2 2
17 3 2 1 10 9 0 13 1 9 7 13 1 9 1 9 0 2
20 10 9 13 16 10 9 13 1 11 2 9 0 13 1 9 1 10 9 13 2
24 2 11 2 2 10 9 1 10 11 2 13 10 9 1 9 12 9 3 2 9 1 9 2 2
19 10 9 2 11 2 7 2 11 2 7 10 9 2 11 2 13 10 9 2
13 11 7 11 13 1 10 9 1 10 9 1 9 2
11 15 13 16 10 9 13 10 9 1 9 2
20 11 3 13 1 11 1 10 12 9 1 9 2 7 13 13 1 10 12 9 2
10 10 9 13 15 10 9 0 7 0 2
67 3 13 15 2 7 13 10 11 2 13 1 10 9 0 2 10 10 9 3 10 11 1 11 1 15 13 13 0 2 13 10 9 1 10 0 7 13 15 2 3 2 1 10 9 0 2 0 2 15 13 13 10 9 2 10 0 9 2 3 15 13 1 10 0 9 13 2
23 10 9 2 11 2 2 13 1 10 11 3 2 11 2 2 13 13 1 10 9 1 11 2
45 10 9 2 13 1 10 9 9 2 13 3 13 4 13 1 10 10 9 1 10 11 2 11 2 2 11 2 2 1 15 2 2 15 11 13 1 10 10 9 1 9 0 3 0 2
5 11 13 9 1 9
28 11 13 12 9 0 1 10 9 1 10 9 1 11 1 10 9 3 1 10 9 1 10 0 9 1 9 0 2
26 2 3 13 10 9 1 10 9 2 13 1 10 11 16 13 10 9 1 10 9 2 2 13 10 9 2
21 1 10 10 9 2 10 9 3 13 13 1 9 3 10 9 0 3 13 10 9 2
1 11
35 1 9 1 10 9 2 11 13 10 9 1 10 9 1 10 9 1 11 2 15 13 10 9 0 1 13 13 10 9 1 9 1 10 11 2
32 11 13 16 10 9 1 9 1 10 11 7 1 10 9 1 9 1 10 9 1 11 3 13 2 0 2 2 7 3 13 9 2
26 10 9 13 1 9 1 10 9 1 11 2 9 1 10 9 2 1 10 9 1 9 0 1 10 11 2
9 11 13 10 9 1 12 1 9 2
11 11 1 10 9 11 13 1 13 9 12 2
20 10 9 3 13 16 10 9 1 9 1 10 11 7 1 10 9 13 10 9 2
18 10 9 1 10 9 2 11 2 13 16 10 9 0 13 4 13 3 2
12 10 9 15 13 13 1 15 13 12 9 2 2
42 3 15 13 9 3 2 3 10 9 1 11 2 11 2 13 13 10 9 1 10 9 10 9 0 15 2 3 2 3 13 1 10 9 1 11 7 13 11 1 10 9 2
47 1 9 1 13 9 2 11 13 11 7 2 1 10 9 0 2 13 15 16 2 3 10 9 1 10 9 13 13 1 10 11 2 15 13 1 3 2 7 1 10 9 1 9 1 10 9 2
10 10 9 1 9 1 10 9 13 0 2
41 10 9 13 3 9 10 9 1 9 2 10 9 1 9 2 10 9 7 10 9 15 13 10 9 3 11 13 13 10 9 1 10 9 2 13 10 9 1 10 9 2
16 13 15 1 10 0 9 1 10 9 1 10 9 0 1 11 2
4 2 11 2 2
43 13 1 10 9 2 11 2 2 10 9 1 10 11 2 10 10 15 13 11 1 10 9 2 2 10 9 13 10 12 9 1 11 1 10 10 9 1 10 0 1 10 9 2
16 1 10 0 9 1 2 11 2 13 0 9 0 1 9 0 2
10 1 11 2 15 13 3 1 10 9 2
39 1 10 10 9 2 15 13 13 1 9 2 9 7 3 10 9 0 2 13 9 1 9 2 9 0 2 2 9 2 9 2 9 2 9 2 9 7 9 2
30 1 10 9 2 13 9 1 9 15 13 2 3 2 10 9 1 10 9 7 10 9 0 2 1 9 0 1 10 11 2
26 1 10 9 1 10 9 2 10 9 13 13 9 0 2 3 9 7 10 9 2 15 13 1 10 9 2
22 1 15 2 15 13 13 13 10 9 0 1 13 10 9 0 1 10 9 1 10 9 2
24 1 13 1 10 9 13 1 10 9 13 2 11 13 13 10 9 1 10 0 9 2 11 2 2
17 10 9 13 16 2 1 9 1 9 2 10 9 13 16 4 13 2
17 1 15 2 2 3 10 0 9 13 13 10 9 1 10 9 2 2
18 1 15 2 9 7 9 3 13 16 13 9 1 11 13 10 0 9 2
34 2 10 9 1 10 11 13 9 1 13 10 9 1 9 7 9 2 7 3 1 10 9 15 13 10 0 1 9 12 2 2 13 11 2
1 9
20 1 13 3 1 10 9 1 11 2 11 7 11 3 13 3 9 1 10 9 2
15 13 10 12 9 11 7 11 7 15 13 1 11 2 11 2
30 1 15 13 0 13 10 9 3 10 9 1 9 9 1 9 7 1 10 9 2 1 10 9 1 10 9 1 10 9 2
18 3 13 0 13 10 10 9 1 10 9 1 15 13 10 9 1 9 2
31 1 10 9 13 0 13 9 1 9 0 7 0 1 10 9 1 10 9 7 13 0 9 1 10 9 7 9 1 10 9 2
4 11 13 0 2
4 13 9 0 2
10 13 9 2 9 0 15 13 9 0 2
18 10 9 13 13 1 10 9 0 2 15 13 1 15 10 0 0 9 2
19 13 13 1 10 11 2 13 1 10 11 2 1 9 12 9 1 12 9 2
24 3 13 10 9 11 2 1 10 9 0 2 11 2 2 13 10 0 9 2 7 15 3 0 2
19 2 11 2 2 9 1 9 1 10 9 1 10 11 2 13 12 12 9 2
22 10 12 9 1 10 11 13 3 13 2 1 0 9 13 1 10 9 3 3 16 0 2
13 15 3 10 9 13 1 10 9 13 1 10 9 2
18 10 9 0 2 0 2 13 16 10 9 3 13 13 3 3 13 13 2
8 3 13 10 9 1 10 9 2
28 2 10 11 13 10 0 9 0 2 2 13 10 9 1 10 9 2 11 2 1 10 9 1 10 2 11 2 2
6 11 2 13 2 10 9
18 9 0 13 9 1 9 2 9 13 16 2 9 13 1 10 9 2 2
24 10 9 3 13 10 2 9 1 12 9 2 1 0 9 1 10 9 1 10 0 7 0 9 2
9 11 2 11 2 9 1 10 11 2
9 11 2 11 2 9 1 10 11 2
31 1 10 9 13 2 10 11 13 12 9 2 15 13 10 9 1 12 11 2 9 12 2 1 10 12 9 1 10 9 13 2
41 2 10 9 13 13 16 10 11 13 10 9 1 9 1 10 10 9 2 2 13 11 2 9 1 10 11 1 10 11 2 10 1 10 12 9 13 1 13 10 9 2
3 9 1 9
12 10 15 3 15 13 13 1 10 9 1 11 2
16 1 10 0 9 1 9 0 2 11 13 3 1 10 0 9 2
25 13 10 0 9 2 7 10 0 9 13 15 15 3 13 10 9 2 7 13 0 2 13 9 0 2
28 16 11 2 1 10 9 2 11 2 2 13 16 10 9 1 11 13 3 10 9 2 10 9 13 3 10 9 2
14 2 10 9 13 11 2 13 10 9 1 10 0 9 2
28 10 9 13 10 9 0 0 1 10 9 2 13 16 10 9 11 2 9 2 3 13 13 2 1 9 1 12 2
37 2 10 9 1 10 9 3 13 1 10 0 9 0 2 15 13 10 9 1 9 2 9 7 9 2 15 1 10 9 1 9 2 2 13 10 9 2
27 10 9 13 9 1 9 0 2 3 13 10 9 2 1 13 7 13 9 3 1 9 0 1 10 9 0 2
17 11 2 15 13 10 9 15 10 9 1 10 9 13 1 10 9 2
14 9 2 3 13 10 9 1 10 9 1 13 10 9 2
25 3 10 9 1 9 15 13 1 10 9 7 1 10 9 13 2 10 9 1 9 0 13 13 3 2
32 13 13 2 1 10 0 2 10 9 0 13 1 10 9 2 7 13 16 9 0 13 13 3 3 16 15 2 3 16 10 9 2
26 9 2 10 9 0 1 10 11 13 10 9 0 1 12 1 10 9 3 1 10 0 9 1 10 9 2
5 11 2 15 13 2
2 9 0
2 9 2
7 2 15 13 10 9 0 2
23 10 9 0 13 9 1 11 2 10 9 13 12 9 9 1 11 2 3 13 10 10 9 2
13 1 3 13 9 1 10 9 2 3 13 1 13 2
21 13 1 9 2 10 9 13 3 10 10 10 9 1 15 13 12 5 1 10 9 2
3 9 0 2
23 1 3 1 10 9 2 10 11 13 1 11 2 1 13 15 3 13 2 13 9 1 9 2
12 7 2 16 13 3 13 13 15 2 0 2 2
49 1 10 0 9 2 12 2 15 13 2 11 2 2 2 11 2 2 2 11 2 2 2 11 2 2 2 11 2 2 2 11 2 2 7 2 11 2 2 2 7 15 13 3 15 15 13 3 13 2
27 3 2 12 13 3 10 0 9 1 11 2 16 15 13 1 9 2 1 10 9 0 2 1 10 12 9 2
32 10 9 13 16 2 3 2 3 13 10 0 9 2 3 15 1 10 9 0 2 0 2 13 1 13 10 0 9 1 10 9 2
28 10 9 0 2 13 2 2 15 13 3 13 10 9 2 13 3 9 0 10 0 2 10 9 3 13 1 9 2
16 1 10 9 1 10 11 2 16 15 13 10 9 1 10 9 2
2 9 0
23 12 9 1 10 9 0 13 0 1 10 9 13 2 1 9 13 1 10 9 0 1 11 2
2 9 0
35 3 12 5 1 10 9 1 10 9 13 16 10 10 9 13 10 9 1 10 9 1 10 9 2 3 12 5 13 16 10 9 13 10 9 2
5 11 15 10 9 2
26 11 2 3 13 10 9 0 2 13 10 9 1 16 15 13 13 13 1 10 9 1 9 0 7 0 2
53 10 9 13 0 9 1 10 9 1 10 9 7 13 15 1 10 11 2 1 10 11 2 1 11 2 3 10 9 13 1 9 12 2 9 12 12 2 1 10 9 7 9 12 2 9 12 12 2 1 9 1 9 2
32 11 7 10 12 9 13 1 9 1 10 9 1 10 11 1 11 2 11 2 1 10 9 11 2 0 1 10 9 1 10 11 2
18 10 9 2 13 1 10 9 2 13 9 12 12 2 9 12 9 2 2
45 10 9 13 0 1 10 10 9 2 3 13 10 9 0 7 10 9 1 10 9 15 13 10 9 1 10 9 7 10 9 1 9 1 10 9 2 7 3 10 9 1 9 0 0 2
71 1 10 9 13 2 15 3 13 3 9 0 2 7 10 9 3 13 1 10 9 1 10 0 12 9 2 15 13 13 10 9 0 1 10 10 0 1 9 0 2 13 15 1 10 9 1 9 0 2 11 2 2 1 10 9 1 10 9 2 11 7 9 2 7 1 10 9 2 11 2 2
7 10 9 1 9 13 3 2
8 13 10 9 0 1 10 11 2
7 7 15 13 13 0 9 2
8 3 2 10 9 13 10 9 2
29 13 16 10 9 1 10 10 9 0 10 9 3 13 4 13 1 9 13 1 10 9 0 7 10 9 1 10 11 2
7 13 3 2 3 13 9 2
14 13 10 9 1 10 9 7 1 10 9 1 10 9 2
3 15 10 2
25 10 9 13 1 10 10 0 9 2 9 7 9 11 2 10 9 1 13 10 9 0 1 10 9 2
33 1 10 9 2 15 15 13 13 10 9 7 10 9 1 10 9 13 3 3 2 13 10 9 2 10 9 2 10 9 7 10 9 2
28 13 10 9 3 0 2 15 13 10 9 1 10 9 0 7 1 10 9 13 1 10 9 1 10 2 9 2 2
17 1 15 13 2 11 2 15 13 13 10 9 2 13 10 0 9 2
30 1 10 9 13 10 9 11 2 1 10 11 2 7 10 9 11 2 1 10 11 2 10 2 9 2 13 1 10 9 2
31 1 12 9 2 10 9 13 16 13 10 9 1 9 1 9 7 13 1 13 10 9 3 10 9 13 1 10 9 13 13 2
17 11 13 9 12 9 1 13 2 11 2 1 10 9 1 10 11 2
58 10 2 9 11 2 3 13 1 10 11 2 1 10 9 1 9 1 10 9 2 11 2 1 9 12 9 1 9 0 2 10 9 1 10 9 1 2 9 2 9 0 7 9 2 1 3 12 9 13 1 10 9 15 13 10 9 3 2
33 10 9 2 13 9 2 13 13 13 2 9 0 2 2 1 10 9 1 10 9 1 10 9 1 10 9 11 7 1 10 9 11 2
5 11 7 11 13 3
16 10 9 1 10 11 13 1 10 9 2 1 10 9 1 9 2
7 10 9 13 13 3 0 2
21 3 1 10 9 2 10 9 13 1 10 11 2 3 13 13 1 10 9 1 9 2
26 13 1 13 10 9 1 9 1 9 2 11 2 1 10 9 11 2 13 9 1 10 9 7 13 11 2
27 13 3 13 1 10 9 7 9 1 13 10 9 1 10 9 2 3 1 10 0 9 1 10 9 1 10 11
5 11 13 10 11 2
22 1 12 10 9 2 2 11 2 13 13 1 13 10 12 9 1 9 1 10 9 0 2
21 16 1 10 9 3 3 13 10 9 2 3 10 9 3 13 10 9 1 10 9 2
10 11 13 15 13 1 10 9 3 0 2
16 15 13 3 0 0 2 16 10 9 13 13 1 13 1 15 2
27 10 9 2 11 2 2 9 11 2 2 1 11 2 13 10 10 9 1 10 9 7 10 9 1 10 9 2
2 11 12
17 10 9 1 10 9 13 10 9 0 1 13 12 9 1 9 0 2
16 10 9 13 1 10 0 9 12 2 1 10 9 1 10 9 2
7 10 9 13 1 11 12 2
2 11 12
22 3 12 12 9 13 9 0 1 10 11 2 11 2 1 10 9 13 2 1 10 11 2
23 1 10 9 0 1 10 9 2 11 2 10 9 1 10 9 13 13 10 9 1 10 9 2
1 11
14 15 13 16 10 9 1 10 9 13 13 0 9 0 2
21 3 1 13 3 9 0 1 10 2 11 2 2 11 13 10 9 1 9 1 9 2
5 11 13 9 1 9
22 9 1 10 11 13 3 1 11 2 11 2 10 9 13 1 9 0 1 10 11 0 2
16 1 15 2 9 1 9 1 9 1 9 13 13 1 10 9 2
30 10 11 7 9 1 10 11 13 16 9 1 9 13 9 1 12 7 12 9 0 16 15 13 1 10 11 1 10 11 2
9 9 7 9 13 10 9 1 10 11
30 1 13 13 10 9 1 10 9 1 9 7 1 10 9 1 10 11 2 10 9 1 10 11 7 10 11 13 10 9 2
15 3 2 10 9 7 10 9 13 13 3 1 13 10 9 2
11 15 13 13 10 2 9 2 1 10 9 2
20 3 3 13 9 3 0 2 3 15 1 10 11 2 10 9 13 13 1 13 2
7 11 13 10 9 1 10 9
19 10 9 13 4 13 3 3 9 2 7 3 10 9 1 9 0 1 10 9
5 1 10 9 1 9
16 3 11 13 1 13 3 1 10 9 2 13 9 1 10 9 2
23 3 13 16 2 3 1 10 9 3 0 1 10 9 2 11 13 1 9 13 1 10 9 2
30 10 9 0 2 0 2 0 1 10 9 2 3 13 1 2 11 2 2 9 11 2 13 3 13 10 9 1 10 9 2
19 3 9 2 11 13 10 9 1 3 13 15 2 7 13 0 13 1 15 2
22 3 10 9 1 10 9 13 13 3 10 9 0 2 13 1 10 11 13 10 0 9 2
2 9 13
31 10 11 13 1 10 11 10 9 1 12 12 9 1 9 2 1 10 9 1 12 12 9 1 9 1 10 9 1 10 9 2
29 1 10 9 2 10 9 1 10 9 13 0 1 15 13 1 10 9 0 2 12 5 1 12 5 1 10 9 2 2
16 11 3 13 13 16 10 11 2 11 2 13 1 13 10 9 2
17 11 13 10 9 1 9 1 12 5 1 9 2 3 1 10 11 2
19 2 10 10 11 13 16 1 9 15 15 13 7 10 9 13 2 2 13 2
48 1 10 9 0 2 10 9 12 1 10 9 12 2 10 9 13 13 1 12 9 1 10 9 0 2 3 12 9 0 1 10 11 7 1 9 1 10 11 13 1 13 10 9 1 10 10 9 2
21 10 9 13 1 10 9 1 10 9 2 13 1 10 9 1 10 9 1 10 9 2
19 10 9 13 1 10 11 7 1 10 11 10 9 1 9 0 1 10 9 2
10 9 1 11 13 15 9 1 10 0 9
15 3 12 9 1 9 13 13 10 9 1 11 1 3 3 2
12 10 9 1 10 11 13 13 12 9 1 9 2
18 10 9 0 1 10 9 1 9 13 3 13 4 13 1 10 0 9 2
15 10 12 9 1 10 11 13 9 0 15 13 10 9 0 2
20 1 10 9 1 10 11 13 12 9 11 2 1 10 11 7 12 9 1 9 2
17 1 10 0 2 13 0 10 11 2 10 11 2 10 11 7 10 11
12 10 9 13 13 12 9 1 15 1 10 9 2
13 16 3 13 9 2 10 9 1 9 13 13 0 2
15 1 10 9 12 2 10 11 3 13 10 9 1 10 11 2
21 12 9 3 1 10 9 2 10 9 0 3 3 13 13 1 10 9 1 10 9 2
29 1 10 9 1 10 9 2 10 9 11 13 10 9 0 1 9 12 9 1 13 15 13 9 15 13 1 10 9 2
24 3 10 9 13 10 11 1 12 10 9 13 13 1 10 11 2 7 10 9 13 9 1 15 2
25 10 9 13 16 10 9 2 11 2 15 3 13 10 11 1 12 2 13 10 0 1 13 10 9 2
24 10 9 1 11 1 12 1 10 11 2 13 10 9 2 13 10 9 1 10 9 2 1 11 2
22 3 2 10 9 13 0 9 1 9 2 9 2 9 1 9 2 9 7 9 1 9 2
21 10 0 13 15 13 1 11 2 3 1 9 7 9 2 3 13 13 9 1 9 2
5 10 9 13 0 2
12 11 13 7 13 3 15 13 13 1 10 9 2
17 0 13 1 10 9 2 13 16 13 0 2 13 15 13 3 2 2
11 10 9 13 2 3 2 13 1 10 9 2
55 1 10 9 1 9 2 10 9 1 10 11 3 13 3 0 1 10 9 2 10 9 1 15 13 9 0 1 13 11 3 13 9 2 10 0 15 13 9 0 1 10 9 2 10 9 1 13 9 1 10 9 1 10 9 2
37 1 10 9 1 10 9 2 10 9 0 2 11 2 13 10 9 1 12 9 2 1 15 12 9 13 16 10 9 13 13 10 0 9 1 10 9 2
39 1 9 1 10 11 2 10 9 1 10 9 3 10 9 2 10 11 0 7 10 9 1 11 7 11 2 1 10 11 2 13 3 9 12 9 1 9 0 2
30 10 2 9 1 9 2 2 9 1 10 9 3 10 12 9 1 16 10 9 13 1 9 2 13 9 0 1 10 9 2
9 10 9 13 12 1 10 9 0 2
18 1 10 9 1 10 11 2 13 15 1 10 10 9 2 13 10 9 2
22 10 9 13 13 1 9 7 13 1 9 13 1 10 9 1 11 2 9 1 10 11 2
37 1 10 11 2 1 10 9 13 1 10 9 10 11 13 10 9 1 9 12 12 3 12 9 1 9 1 9 1 9 1 11 2 3 1 13 13 2
2 9 0
16 1 15 2 13 16 15 13 10 9 0 1 13 9 1 9 2
29 10 9 13 13 1 10 9 1 13 10 9 1 10 9 1 0 9 1 10 9 0 2 1 10 9 1 13 9 2
24 3 3 15 13 10 9 1 10 9 2 13 16 10 9 13 1 9 0 10 9 1 10 9 2
25 10 9 1 10 9 13 1 13 3 1 10 9 0 2 15 3 13 13 1 10 0 9 1 9 2
30 13 10 9 1 10 9 0 1 10 9 15 13 1 10 9 7 13 9 1 16 3 13 9 1 10 9 2 13 11 2
5 13 9 1 10 9
29 13 13 3 1 10 9 11 2 1 11 2 9 9 1 11 2 2 10 9 1 10 11 1 10 9 11 2 12 2
23 11 13 1 9 0 1 10 9 2 9 1 10 9 0 1 9 1 9 1 10 9 2 2
6 9 13 9 0 1 11
29 10 9 11 2 13 1 10 9 1 13 13 9 3 10 9 11 2 13 10 9 1 9 1 10 9 2 11 2 2
24 1 10 9 2 11 2 2 10 9 13 9 1 15 11 13 13 9 0 1 10 9 2 11 2
22 10 9 13 9 1 12 5 1 10 9 1 10 9 1 15 15 13 1 13 10 9 2
16 3 2 13 9 1 9 7 9 1 9 1 15 13 13 3 2
13 10 9 1 10 9 13 13 10 9 1 10 9 2
20 13 0 13 9 0 2 1 10 15 13 13 9 1 9 1 10 2 11 2 2
11 10 9 2 3 2 3 13 9 7 9 2
9 10 9 13 2 13 10 9 2 2
35 10 9 13 16 10 9 0 1 10 9 13 10 9 0 1 10 0 9 2 16 15 3 13 10 9 1 13 15 7 3 13 9 1 15 2
13 10 9 13 1 10 0 9 1 10 7 1 15 2
17 15 2 9 2 9 7 0 9 2 13 10 0 9 1 15 10 2
11 13 10 9 13 10 9 0 1 10 9 2
16 3 2 10 9 13 1 10 9 0 13 1 9 0 7 0 2
24 3 13 15 0 2 1 9 0 2 0 7 0 2 13 10 9 1 9 1 10 9 1 9 2
29 10 9 13 15 2 1 10 9 1 10 9 0 2 1 9 1 9 1 10 9 2 1 10 9 7 1 10 9 2
17 10 9 3 3 13 12 9 1 9 1 9 13 1 9 1 12 2
11 7 2 1 10 9 2 13 13 12 9 2
48 3 13 10 9 2 16 10 0 9 0 1 9 13 15 3 3 3 1 10 9 1 9 13 2 1 15 2 13 1 13 10 9 1 10 9 2 16 15 9 13 2 0 13 10 9 1 9 2
29 13 13 10 9 0 2 3 10 9 1 10 9 2 7 2 3 2 13 10 9 1 9 3 13 3 10 9 0 2
21 13 3 13 16 10 9 13 2 3 13 2 13 1 10 9 10 9 15 15 13 2
30 1 10 9 0 3 1 9 12 7 10 9 13 16 3 13 9 1 3 2 10 0 9 13 3 13 1 10 13 9 2
32 10 9 1 11 3 13 9 1 12 1 10 3 13 9 0 1 11 2 10 11 2 15 13 1 12 1 10 11 1 10 11 2
32 10 9 2 1 13 0 9 15 3 15 2 13 2 1 10 11 2 3 11 2 13 1 11 13 10 9 3 0 1 10 9 2
22 1 10 11 2 11 13 1 0 2 1 12 5 2 1 10 9 1 9 2 1 10 9
12 11 13 10 0 1 10 11 2 1 12 5 2
8 13 0 10 9 0 7 0 2
12 10 9 1 13 13 13 10 9 1 10 9 2
28 1 12 9 10 9 3 3 13 10 9 1 10 9 2 11 2 1 10 10 11 2 7 11 2 1 10 11 2
8 13 10 9 15 13 10 11 2
10 13 10 0 9 0 15 13 1 11 2
20 10 9 3 15 13 9 2 7 2 3 2 15 13 16 13 13 10 9 0 2
17 1 10 0 9 2 9 0 13 1 10 9 1 9 1 10 9 2
12 10 9 3 13 10 9 2 3 3 13 11 2
14 10 9 13 10 9 0 2 10 9 13 10 9 0 2
15 3 3 2 11 13 13 10 9 0 2 13 12 9 0 2
26 1 10 9 11 7 1 10 9 11 2 10 9 11 13 15 3 1 10 9 0 7 13 13 3 3 2
12 15 15 13 9 1 10 11 2 1 10 11 2
17 10 9 0 13 1 10 11 16 3 13 9 7 9 1 10 11 2
8 10 11 0 3 13 10 9 2
10 10 9 13 13 1 9 1 10 9 2
19 10 9 1 10 11 13 1 10 9 1 3 7 3 13 3 1 10 9 2
10 10 11 13 1 10 9 1 9 13 2
23 10 11 3 3 13 10 9 0 1 10 9 2 7 13 16 3 12 9 13 13 10 9 2
31 1 9 0 2 13 10 9 1 9 1 9 15 2 1 13 10 9 1 9 2 13 1 10 0 9 9 0 1 10 0 2
45 13 16 15 13 2 1 10 11 2 1 10 9 1 9 0 0 2 15 13 13 2 1 10 0 9 2 10 9 0 1 10 9 7 13 1 10 9 0 1 13 1 10 9 0 2
21 2 10 10 9 13 0 1 15 1 11 16 1 10 11 15 13 15 1 9 2 2
19 10 9 13 16 3 1 13 1 10 11 13 10 9 3 13 2 10 11 2
19 3 13 2 1 10 11 2 10 12 9 1 10 9 1 9 1 10 9 2
33 2 16 13 16 13 10 9 0 2 15 13 13 10 9 0 2 2 13 11 1 12 9 1 9 1 11 2 3 2 1 10 9 2
30 11 13 16 10 11 13 13 10 9 7 9 1 10 10 9 1 9 1 10 9 1 10 9 1 10 9 0 7 0 2
12 10 9 1 10 9 13 13 0 1 10 11 2
36 10 9 13 1 10 0 11 2 1 10 9 1 10 9 2 13 1 10 11 2 9 11 2 11 2 11 7 13 2 3 2 1 10 9 11 2
28 10 9 1 11 3 13 1 13 0 9 1 10 9 1 10 9 1 10 9 11 2 1 10 9 1 10 9 2
28 3 13 16 13 0 2 13 3 0 10 9 13 12 11 16 11 13 9 1 9 13 1 10 9 1 9 13 2
2 13 2
30 3 13 10 9 2 11 13 1 13 11 12 9 1 16 10 9 13 1 10 9 1 10 9 2 13 10 9 1 9 2
7 10 9 1 11 13 0 2
12 10 9 1 10 11 13 1 10 9 1 12 2
8 3 13 16 13 13 10 9 2
12 13 15 13 1 10 9 1 13 15 10 9 2
3 9 13 9
33 10 0 1 10 9 1 11 1 10 9 1 10 11 2 9 1 9 2 13 9 1 10 9 1 9 2 9 7 9 7 13 9 2
25 10 9 13 12 5 1 9 1 11 2 11 7 11 7 12 5 3 12 5 1 9 1 10 9 2
6 10 9 13 12 5 2
46 10 11 1 10 11 7 1 10 11 2 9 1 9 2 15 13 3 1 9 1 10 11 2 9 1 10 9 1 10 11 2 3 1 10 9 1 10 9 1 10 9 2 1 10 9 2
12 10 9 13 12 5 7 10 9 13 12 5 2
15 10 9 2 1 9 2 13 3 12 9 7 12 12 9 2
6 11 13 9 9 2 11
20 9 1 10 9 13 9 0 1 10 11 1 3 13 9 1 9 2 1 11 2
38 10 9 1 10 11 2 11 2 12 2 13 13 10 9 1 10 11 1 13 10 9 12 9 0 15 15 13 13 13 1 9 1 9 0 1 10 9 2
33 15 13 10 9 0 1 3 13 3 10 9 1 13 10 9 1 10 9 1 9 7 1 3 13 10 9 13 1 10 9 1 15 2
7 10 9 13 0 9 0 2
32 11 2 15 13 1 10 11 7 1 10 10 9 0 15 13 11 1 13 1 10 11 2 13 13 15 13 1 9 1 10 9 2
18 10 9 13 3 0 16 3 7 12 1 10 0 9 13 0 1 11 2
22 10 9 15 13 1 3 2 13 2 10 9 2 1 10 9 1 10 9 1 10 11 2
16 13 16 10 9 0 13 15 13 1 10 9 1 9 1 9 2
36 3 13 10 9 1 10 9 0 7 2 1 10 9 1 9 2 13 10 9 15 13 13 10 9 0 1 10 9 10 9 0 7 10 9 0 2
27 1 13 10 9 1 10 9 2 11 13 10 9 1 9 13 1 10 9 0 1 10 9 2 11 2 1 11
26 1 13 10 9 2 10 9 1 10 9 13 10 9 1 10 9 1 10 9 1 10 9 1 10 9 2
19 3 13 2 2 10 9 13 1 9 0 13 1 4 13 1 10 9 2 2
14 3 12 12 9 13 1 10 9 2 1 10 9 11 2
7 10 9 11 3 13 3 2
15 13 1 10 9 1 9 2 11 2 13 3 1 10 9 2
9 1 11 2 11 2 13 13 2 2
27 10 9 11 13 3 16 10 9 11 2 11 2 9 1 10 9 13 9 1 10 9 11 2 13 13 2 2
15 2 15 13 13 1 10 11 2 2 13 11 2 1 9 2
15 11 13 1 10 11 1 12 9 7 13 13 1 10 9 2
11 10 9 1 10 9 13 13 3 3 0 2
7 9 13 10 0 2 9 2
26 13 1 10 9 0 13 1 9 1 10 9 13 1 13 9 2 9 7 9 3 0 7 1 0 9 2
25 7 13 0 9 1 13 1 9 10 2 1 9 7 9 1 10 9 2 13 10 9 1 10 9 2
47 10 9 11 2 9 1 10 9 0 15 15 13 1 12 9 2 13 10 9 1 13 10 9 1 10 9 13 1 10 9 11 3 9 1 10 9 15 2 1 12 2 13 1 9 12 9 2
43 10 9 1 10 9 11 2 9 11 2 13 16 10 9 1 10 9 13 15 1 10 2 9 2 1 10 9 15 4 4 0 1 10 11 2 13 1 10 9 1 10 11 2
26 10 9 13 0 1 10 9 1 9 0 13 1 10 9 11 7 13 1 13 3 15 13 3 3 13 2
20 1 3 2 10 11 13 1 1 12 9 2 1 10 9 13 1 10 9 0 2
12 1 10 9 2 10 0 9 3 13 9 10 2
11 15 13 10 9 1 10 9 1 12 9 2
25 10 9 1 10 9 1 10 11 2 11 2 2 11 2 13 10 9 1 11 1 10 2 11 2 2
5 11 11 2 9 2
20 11 2 9 1 10 0 2 13 16 10 9 13 1 10 11 13 1 10 9 2
14 2 15 3 3 13 13 1 10 9 0 2 2 13 2
16 10 9 1 11 3 13 3 9 12 9 1 13 10 10 9 2
18 13 10 9 11 2 10 0 9 1 9 1 9 2 1 10 10 11 2
19 13 10 0 2 10 10 9 1 10 9 3 15 13 1 10 9 1 11 2
22 10 9 13 10 9 0 2 11 2 15 3 13 10 9 2 13 10 9 1 9 0 2
15 1 15 2 10 9 0 3 15 13 1 13 10 10 9 2
13 1 10 9 2 12 1 15 3 13 13 10 11 2
9 15 13 10 10 9 1 10 9 2
12 10 9 1 12 3 13 13 0 1 10 11 2
20 10 9 2 15 1 10 9 12 13 10 9 0 2 13 1 13 1 10 0 2
10 3 2 3 13 13 1 10 12 0 2
25 1 12 2 1 10 9 1 11 2 10 9 13 1 0 9 2 9 15 13 0 9 1 10 9 2
9 11 13 1 10 11 1 12 1 12
26 10 11 13 1 12 1 12 1 10 11 2 1 11 2 3 1 10 9 1 10 9 11 2 1 11 2
16 1 10 11 2 13 10 0 9 1 10 9 1 13 10 9 2
17 11 2 9 1 10 9 1 11 2 13 10 9 1 10 12 9 2
32 11 2 13 9 1 10 9 1 10 9 2 13 10 9 1 10 12 9 2 1 9 1 9 1 10 9 11 2 1 10 11 2
20 1 15 13 10 9 2 1 10 11 10 0 9 13 1 11 2 1 12 9 2
17 3 3 2 10 9 11 13 16 10 9 0 13 1 10 0 9 2
12 13 10 9 1 10 9 13 10 9 3 0 2
3 9 2 9
2 9 0
27 10 9 11 13 2 3 10 9 0 2 10 9 1 13 10 9 1 10 9 1 10 9 1 15 3 13 2
19 13 3 13 1 10 9 1 10 9 16 13 10 10 9 7 13 10 9 2
30 3 2 10 9 1 10 9 1 13 9 0 1 10 9 11 2 3 10 9 13 1 10 9 1 3 2 13 1 9 2
31 16 3 13 1 10 11 1 3 2 13 3 0 2 1 10 9 1 0 9 0 2 15 10 9 13 10 9 7 15 13 2
19 11 3 13 9 1 13 10 9 2 11 2 9 1 10 11 2 1 12 2
44 10 9 13 10 2 9 0 2 1 10 0 9 1 10 9 2 12 9 0 1 10 9 1 10 11 1 10 9 1 10 11 1 10 2 9 0 2 13 1 10 9 1 11 2
24 10 9 1 11 13 16 15 3 13 13 3 1 9 7 9 2 1 11 3 13 2 3 13 2
26 10 9 13 10 9 1 16 10 11 13 10 9 1 10 9 15 13 16 10 9 13 13 1 10 11 2
8 11 2 3 13 9 1 9 2
6 3 13 13 9 0 2
27 3 13 13 9 1 10 9 0 7 2 1 10 9 0 2 10 11 13 13 10 9 1 9 1 10 9 2
7 13 1 10 9 1 9 2
34 11 2 7 1 10 9 1 15 10 0 9 13 13 2 16 10 9 13 13 1 10 9 2 3 13 0 10 9 0 2 10 9 0 2
6 9 0 13 13 13 9
48 10 9 1 9 2 11 2 2 1 10 9 1 10 9 11 2 11 2 2 13 13 13 1 10 9 1 10 9 1 10 9 1 9 0 1 10 11 2 11 2 13 1 15 3 9 1 9 2
51 1 10 10 9 13 3 1 10 11 2 15 13 13 13 10 2 9 1 9 2 1 10 9 1 10 9 1 15 11 13 16 10 11 2 16 13 10 9 0 2 13 13 2 10 9 1 10 9 0 2 2
42 9 0 2 9 1 10 9 7 12 1 10 9 1 10 11 1 10 9 1 11 2 11 13 3 10 9 9 1 10 9 2 10 9 1 10 9 7 1 10 9 0 2
16 11 2 15 13 10 9 0 1 9 1 10 9 1 10 9 2
1 9
27 1 13 15 13 1 10 9 7 1 10 9 1 10 9 1 10 9 1 10 11 2 11 13 3 9 3 2
29 1 10 9 11 2 13 1 11 10 9 1 10 9 1 10 9 2 3 3 13 13 13 9 1 9 2 0 9 2
6 9 13 9 1 10 11
29 10 9 9 2 0 0 9 1 9 1 10 9 2 13 9 1 10 9 1 10 12 9 11 2 10 13 1 11 2
20 10 9 13 10 9 3 1 9 1 10 9 1 9 7 1 9 1 10 9 2
6 3 2 10 9 13 2
15 11 2 1 15 3 13 9 15 3 13 1 10 10 9 2
8 11 2 3 2 7 1 3 2
21 10 9 1 10 11 13 10 9 1 10 0 9 3 15 2 13 1 10 9 2 2
14 1 3 2 10 9 1 11 13 3 4 13 10 9 2
13 2 10 9 3 15 13 2 2 13 1 9 11 2
35 10 9 15 13 3 1 16 2 16 13 10 9 2 13 15 13 9 1 11 7 13 10 9 1 9 1 10 9 1 10 9 1 10 11 2
16 10 9 1 11 1 15 13 9 3 13 10 9 15 15 13 2
19 2 15 3 13 13 10 9 11 2 2 13 11 2 11 2 2 1 11 2
21 11 13 10 9 1 13 1 10 9 11 2 15 15 13 1 9 1 3 13 11 2
18 2 1 15 13 13 9 1 10 9 2 13 9 7 9 2 2 13 2
22 1 13 10 9 0 1 11 2 13 10 9 0 11 2 11 2 2 9 1 10 9 2
23 2 15 13 3 7 13 9 12 9 2 12 5 1 10 9 1 10 9 2 2 2 13 2
7 13 11 2 1 10 11 2
1 9
29 1 10 10 9 2 10 0 9 1 15 13 2 12 5 2 13 16 11 13 9 1 9 1 10 9 1 10 9 2
22 13 10 0 9 2 3 2 15 13 0 1 10 9 1 13 16 11 3 13 13 9 2
5 13 3 12 5 2
14 1 15 12 5 2 13 9 7 3 1 13 10 9 2
18 11 13 16 13 10 9 1 10 9 1 13 1 10 9 0 2 11 2
14 1 11 2 11 3 15 13 15 1 9 1 10 9 2
21 2 13 13 16 10 9 1 11 7 15 1 10 11 13 9 1 10 0 9 0 2
17 3 2 13 13 9 1 10 9 1 10 9 0 2 2 13 11 2
1 11
5 7 15 13 13 2
7 11 2 7 13 10 9 2
16 15 13 10 9 1 12 9 2 13 16 10 9 13 15 13 2
17 13 10 9 1 13 2 7 13 16 15 15 13 1 13 10 9 2
13 13 16 10 9 2 11 2 13 13 1 0 9 2
22 10 9 1 11 2 15 13 9 0 2 13 9 7 13 13 1 9 7 9 1 9 2
5 1 13 1 11 2
34 10 9 1 10 9 13 1 10 9 15 11 13 1 9 1 12 1 10 2 11 2 1 10 9 11 2 1 10 9 13 1 10 11 2
13 2 10 9 1 10 9 15 13 7 13 10 9 2
17 13 10 9 7 13 1 13 10 9 1 10 9 2 2 13 11 2
12 1 10 9 1 9 13 9 0 1 12 9 2
20 1 10 9 1 10 9 2 4 3 13 15 9 1 9 13 11 2 11 2 2
4 9 1 13 0
16 11 3 3 3 10 9 13 13 10 9 1 10 9 3 0 2
27 10 9 13 0 2 9 1 9 2 9 1 9 7 9 1 9 2 9 0 2 9 0 1 10 10 9 2
22 13 10 9 1 3 13 3 15 2 13 3 1 13 1 10 9 7 13 13 10 9 2
3 3 3 2
21 16 13 10 9 1 9 1 10 9 3 10 9 1 9 2 13 15 13 10 9 2
13 3 3 13 16 3 13 16 10 9 3 15 13 2
5 1 10 9 1 9
6 13 10 9 1 9 2
3 13 0 2
3 13 9 2
3 13 9 2
7 7 3 13 10 9 10 2
10 2 15 3 13 9 2 13 0 2 2
2 6 2
3 7 9 2
2 9 2
3 11 9 2
16 10 9 0 13 10 9 9 2 10 9 1 9 7 12 9 2
2 6 2
5 13 10 9 2 2
3 13 9 2
7 7 10 9 1 10 9 2
5 11 2 11 7 11
4 7 10 9 2
7 2 11 13 10 9 2 2
7 2 9 0 3 11 2 2
11 7 9 1 9 1 9 13 9 1 0 2
6 2 15 13 13 2 2
4 2 6 2 2
6 2 15 13 13 2 2
8 2 6 2 15 13 13 2 2
9 2 6 13 16 15 13 13 2 2
3 13 0 2
5 13 0 7 13 2
5 3 1 10 9 2
11 13 1 10 9 10 12 9 1 10 11 2
12 0 13 10 11 15 13 13 1 10 10 9 2
2 0 2
2 13 2
6 9 1 10 9 3 2
6 13 9 1 10 9 2
9 10 11 1 10 11 13 10 9 2
12 15 13 10 0 9 1 10 11 2 10 9 2
10 3 10 11 7 10 11 3 13 9 2
16 3 1 10 11 2 1 11 2 11 2 10 9 13 10 9 2
6 9 2 13 10 9 2
5 13 9 1 9 2
10 7 3 11 2 9 2 9 7 9 2
12 7 15 13 16 13 10 9 7 13 10 9 2
8 9 1 10 9 2 11 2 2
3 9 0 2
8 10 9 1 9 13 3 0 2
10 3 3 1 10 9 13 1 10 9 2
29 1 10 11 15 3 13 1 12 9 1 9 0 2 9 2 9 2 9 2 9 2 9 2 9 2 9 7 9 2
10 7 13 9 15 3 13 1 10 9 2
2 6 2
7 9 13 13 10 9 10 2
6 12 9 13 1 9 2
23 10 9 1 9 11 2 1 10 9 2 9 2 13 9 1 9 1 9 7 13 9 0 2
6 9 2 1 9 12 2
17 1 10 9 2 10 0 13 10 11 2 13 9 1 10 9 2 2
19 7 13 12 3 0 2 3 1 15 2 10 9 13 3 1 9 1 9 2
9 2 13 10 9 3 0 7 0 2
14 10 9 13 1 9 1 9 2 16 15 13 3 3 2
14 3 1 11 2 15 13 13 10 9 2 2 13 9 2
2 10 9
24 1 11 2 10 12 9 3 0 1 10 9 13 9 1 10 9 1 10 0 9 1 10 11 2
20 10 9 0 2 1 15 10 1 10 11 2 13 13 1 9 13 1 10 9 2
28 1 15 13 13 10 9 1 10 9 10 9 1 9 3 13 10 9 2 15 13 16 13 9 1 10 3 9 2
60 1 11 2 1 10 11 2 1 10 9 3 0 2 13 9 1 10 9 2 13 10 9 1 9 2 11 2 2 13 1 12 9 0 2 9 1 10 9 9 0 2 9 1 9 2 9 0 2 9 1 9 2 9 1 9 7 9 1 9 2
22 10 9 2 13 2 10 9 7 13 13 1 9 15 13 9 0 2 3 9 7 9 2
37 13 0 16 13 10 9 1 16 10 10 9 2 15 13 9 0 15 13 10 9 1 9 7 9 1 9 1 10 9 2 13 10 9 1 10 9 2
9 3 13 13 13 10 9 1 11 2
13 15 13 10 9 1 9 1 13 10 9 1 9 2
9 11 13 1 10 9 1 10 9 2
15 11 13 10 9 1 10 11 0 7 10 9 1 10 9 2
38 2 10 11 3 13 10 9 15 13 9 1 10 11 2 2 13 10 9 0 2 13 13 10 9 1 2 9 0 2 13 1 10 10 9 1 10 11 2
52 2 15 3 13 13 16 10 9 3 0 3 10 1 10 11 13 13 9 3 13 13 1 3 2 2 13 2 13 15 1 10 9 1 10 0 9 1 10 11 2 15 13 1 10 9 1 10 9 1 10 11 2
83 12 2 10 0 2 13 15 15 10 11 13 7 13 3 9 0 10 9 1 10 9 0 13 7 0 7 3 1 9 0 1 9 2 13 0 1 10 9 10 9 7 9 0 13 10 9 2 7 10 9 1 10 9 1 9 1 9 7 1 9 2 1 9 0 7 9 1 10 9 0 2 13 10 9 1 9 1 10 9 1 9 13 2
45 10 15 2 0 7 0 2 13 1 13 10 9 0 1 10 9 2 1 10 9 0 2 1 10 9 13 1 10 10 9 0 1 9 1 10 9 1 9 2 13 15 9 7 9 2
30 10 9 3 13 0 3 1 10 11 1 0 9 1 9 1 9 0 1 13 10 9 1 10 9 0 1 10 9 11 2
25 10 9 1 9 13 1 10 9 1 10 9 0 13 1 12 5 1 10 9 0 1 12 5 3 2
52 10 9 13 1 10 0 9 1 2 11 2 2 1 9 13 1 11 7 3 1 9 1 9 2 13 10 9 1 11 2 15 1 12 13 10 9 0 2 0 7 0 1 13 10 9 1 10 9 2 11 2 2
14 10 0 2 12 9 2 2 0 7 0 11 13 13 2
37 10 9 15 1 13 13 1 2 11 2 2 11 2 3 3 13 3 13 1 10 9 1 10 9 16 2 1 10 9 2 11 3 13 1 10 9 2
1 9
30 1 10 9 2 10 0 7 0 9 15 13 2 13 9 7 9 10 9 0 13 3 3 16 10 9 1 10 9 0 2
27 3 15 12 13 13 2 2 11 2 2 2 11 2 2 2 11 2 2 2 13 10 9 1 10 10 9 2
24 7 9 1 9 1 10 9 2 15 3 13 10 9 1 13 1 10 2 9 2 1 10 9 2
23 1 12 1 15 2 2 11 2 7 2 11 2 2 10 1 9 1 11 2 13 10 9 2
5 11 13 2 11 2
21 10 9 15 11 13 1 9 1 12 7 9 1 12 13 0 9 1 10 9 1 12
18 10 9 11 2 12 2 13 15 13 1 13 10 9 1 10 9 0 2
30 9 15 13 2 13 1 13 2 11 2 2 9 1 11 15 10 9 13 1 0 9 1 9 1 12 7 9 1 12 2
25 10 9 13 13 10 2 9 2 1 9 1 12 2 1 10 9 2 1 10 9 1 2 11 2 2
4 15 1 10 9
15 1 10 9 1 10 10 10 9 1 9 13 10 10 9 2
6 13 15 1 10 9 2
23 10 0 9 1 10 9 1 10 9 1 10 11 1 10 11 13 10 9 0 1 10 9 2
38 13 10 9 15 13 10 9 15 13 1 13 7 2 3 2 13 2 13 9 1 10 9 7 13 2 3 2 10 9 2 15 13 9 2 9 7 9 2
35 13 16 9 3 9 2 9 7 9 2 13 10 9 1 10 9 1 10 9 2 13 3 16 3 2 13 10 9 1 10 9 1 10 9 2
32 11 2 11 2 11 7 10 10 2 9 2 2 9 0 1 10 9 2 13 16 10 9 1 10 9 0 13 1 10 9 0 2
16 10 0 9 13 10 9 0 1 10 9 2 15 13 10 9 2
14 1 10 9 0 1 9 2 10 9 13 10 12 9 2
19 15 13 13 1 11 2 9 3 13 13 10 9 2 1 9 1 12 9 2
29 3 1 10 10 9 2 3 10 9 13 3 10 9 2 10 9 0 2 10 9 2 10 9 7 9 0 7 0 2
17 10 9 1 11 2 1 13 13 13 1 10 11 2 13 10 9 2
15 10 9 2 3 3 13 7 0 2 13 1 13 1 9 2
8 10 11 13 10 9 3 0 2
8 13 1 15 12 7 15 12 2
9 10 9 11 13 13 10 0 9 2
32 3 13 3 15 15 13 1 13 3 10 9 1 9 0 2 3 13 10 9 1 10 11 7 13 10 9 1 10 9 0 0 2
13 7 10 9 13 1 10 9 1 9 1 10 9 2
33 3 1 10 0 9 0 2 10 9 1 10 9 0 1 10 9 1 10 10 9 1 10 9 0 13 9 0 0 1 10 9 0 2
47 13 0 13 2 3 2 1 10 9 0 1 10 9 1 9 0 2 15 10 9 0 1 11 7 11 1 10 9 1 10 9 0 0 1 10 9 1 10 9 13 3 1 10 9 1 9 2
19 11 13 1 10 9 1 9 1 11 2 11 2 2 7 3 13 13 9 2
7 2 3 13 1 10 9 2
10 13 16 3 13 9 0 2 2 13 2
7 1 12 15 3 13 13 2
13 2 10 11 13 13 10 10 9 7 13 10 9 2
7 13 13 7 3 13 13 2
13 7 13 3 13 10 9 1 10 9 2 2 13 2
13 11 13 16 13 10 9 0 1 11 1 12 9 2
6 3 13 13 9 0 2
17 13 16 13 13 3 9 1 10 10 9 0 13 1 3 12 9 2
27 10 9 11 13 3 10 2 9 2 1 10 9 2 3 1 11 2 2 1 10 9 0 1 13 9 2 2
19 3 2 13 10 9 16 13 10 9 2 1 13 15 1 10 9 3 13 2
7 9 1 10 9 2 3 2
18 3 2 3 2 7 3 3 3 15 13 1 10 0 9 1 10 9 2
24 1 9 2 10 9 1 9 3 0 13 1 10 9 1 10 11 2 1 10 11 2 1 9 2
45 1 3 13 10 9 1 10 9 0 13 10 9 2 16 15 3 13 4 13 1 10 9 1 10 9 15 13 3 12 9 1 9 2 3 3 16 10 9 0 1 10 10 9 0 2
11 10 9 11 3 13 13 10 9 1 11 2
18 1 15 2 10 9 1 10 9 13 10 2 9 0 2 1 10 9 2
14 2 13 1 9 13 10 9 1 10 11 2 2 13 2
21 11 2 3 2 13 16 10 9 13 13 10 9 7 2 13 10 9 2 1 11 2
11 10 9 13 13 10 0 9 1 15 13 2
22 10 9 1 9 1 10 11 2 11 2 13 16 10 9 13 13 10 9 1 10 11 2
13 2 15 15 15 13 13 10 9 1 10 9 0 2
5 10 9 13 0 2
12 10 11 13 1 13 10 9 1 9 7 9 2
17 16 15 3 13 10 9 2 13 4 13 9 0 2 2 13 11 2
24 2 10 9 0 13 15 13 13 1 13 9 0 1 10 9 7 9 0 2 2 13 10 9 2
14 10 9 13 10 9 1 10 9 13 1 9 1 9 2
18 7 13 10 9 1 9 2 3 15 15 13 11 1 10 9 1 12 2
18 10 11 3 13 10 9 3 10 9 13 1 9 10 9 1 10 9 2
24 3 3 10 9 13 1 9 7 3 10 9 3 13 9 1 9 2 10 9 13 13 3 9 2
17 10 11 13 3 10 9 7 10 9 0 3 0 2 3 10 9 2
16 10 9 0 1 9 3 13 2 13 2 10 9 1 10 9 2
20 1 10 9 1 10 9 0 2 13 0 13 15 7 13 10 9 1 10 9 2
21 10 9 2 10 9 1 9 13 11 2 13 10 9 1 9 12 12 7 13 13 2
10 10 9 13 13 1 11 1 10 9 2
15 10 9 1 10 9 1 10 9 13 13 1 10 9 0 2
27 2 13 9 2 1 10 9 13 9 0 2 3 13 10 9 10 2 2 13 11 2 12 2 9 1 9 2
20 11 13 1 10 9 11 2 11 2 3 1 10 0 9 1 9 1 10 9 2
16 13 1 12 9 3 2 11 13 16 3 13 10 9 3 0 2
10 2 1 12 9 16 10 9 13 0 2
13 1 10 9 2 13 10 9 3 0 2 2 13 2
20 10 9 1 10 11 13 16 10 9 1 9 13 1 9 12 9 1 10 11 2
20 1 12 2 3 2 10 9 1 10 0 9 1 10 11 1 10 11 13 13 2
10 2 13 13 10 9 1 9 1 12 2
17 10 9 13 13 15 1 0 9 7 10 9 0 2 2 13 11 2
23 1 10 11 13 13 10 11 2 11 2 2 1 9 1 10 11 2 11 2 11 7 11 2
7 10 11 13 1 9 0 2
7 7 13 0 10 9 11 2
33 13 3 2 13 10 9 0 7 15 2 16 13 1 10 10 9 0 2 10 11 2 13 13 10 9 0 15 10 9 13 7 13 2
35 11 2 12 2 9 1 9 1 10 9 1 11 2 11 2 2 13 9 1 10 9 1 11 1 10 11 7 9 1 10 11 2 11 2 2
18 13 9 1 10 9 7 1 11 1 10 9 1 11 2 9 11 2 2
24 3 1 15 11 13 1 10 9 2 15 13 13 3 3 0 16 10 9 3 13 13 1 15 2
18 7 13 10 9 16 15 13 10 9 1 10 2 10 9 1 10 9 2
37 13 10 9 1 10 9 7 9 1 10 9 1 10 9 12 7 13 10 9 1 16 15 3 15 13 13 3 13 10 9 1 16 13 15 1 9 2
13 2 1 10 9 2 13 3 10 11 2 2 13 2
36 3 1 11 2 10 9 1 9 1 10 9 13 12 9 1 13 7 10 9 3 13 1 13 15 13 15 1 10 9 0 1 10 11 2 11 2
23 1 15 2 10 9 0 1 10 9 13 4 13 1 10 9 1 10 11 11 2 11 2 2
26 1 11 2 10 9 1 9 13 2 10 9 1 9 2 1 10 9 10 0 9 0 1 10 9 0 2
18 2 13 10 9 0 1 13 10 9 15 13 13 10 11 1 10 11 2
25 10 9 0 1 13 10 9 2 10 9 7 15 13 10 9 1 9 1 10 9 2 2 13 11 2
4 13 9 0 2
19 16 15 13 15 2 13 1 13 1 9 0 7 13 10 9 1 10 9 2
13 13 3 1 10 11 2 9 2 7 13 10 9 2
3 1 10 9
9 2 3 13 3 10 15 1 2 11
21 10 9 13 1 10 9 7 15 13 1 15 15 3 13 13 10 9 1 10 9 2
3 15 13 2
18 13 13 16 13 10 9 7 13 1 10 9 1 10 11 7 13 2 2
92 10 11 13 10 9 1 10 11 2 3 1 9 7 1 9 2 7 9 1 10 10 9 13 10 11 2 15 13 13 15 13 2 1 11 1 11 2 13 16 2 1 10 9 1 11 1 15 13 2 10 11 13 13 10 11 2 1 10 9 12 2 15 3 15 13 1 9 0 1 10 9 2 1 10 0 9 2 0 1 10 9 1 10 9 7 1 10 9 1 10 9 2
16 10 11 3 13 1 10 10 9 16 15 13 13 1 10 11 2
40 7 3 13 1 15 16 3 13 10 0 9 1 15 3 11 2 10 0 2 9 2 2 15 1 15 9 13 10 9 1 10 10 9 7 9 1 10 9 0 2
27 3 11 13 13 1 10 10 9 0 2 13 11 2 15 13 16 10 11 13 10 9 1 9 7 1 9 2
4 9 13 9 0
12 10 11 7 11 13 9 1 10 9 0 3 2
14 10 11 13 10 9 1 11 7 11 2 1 10 9 2
16 10 11 13 1 9 10 9 1 11 7 11 2 1 10 9 2
7 9 9 13 12 1 10 11
36 9 1 10 11 13 1 10 9 0 10 9 1 12 9 2 13 1 13 1 13 11 2 9 9 13 1 10 9 3 3 1 10 9 1 12 2
13 10 9 13 9 1 13 10 12 9 0 1 9 2
24 10 9 11 13 1 10 9 1 12 9 2 3 9 1 10 9 9 1 10 9 1 10 9 2
6 11 13 9 1 12 9
14 11 2 12 2 13 13 1 12 9 1 9 1 11 2
23 15 13 7 13 12 9 1 10 9 1 15 13 10 9 1 10 9 1 15 15 13 0 2
12 10 9 13 1 9 2 9 7 9 1 9 2
19 13 10 0 9 1 10 11 15 10 9 13 10 9 11 3 10 9 0 2
19 10 9 1 9 13 1 10 11 13 13 1 10 9 1 10 11 2 11 2
11 1 10 9 2 3 13 9 1 10 11 2
31 3 2 10 9 0 13 1 13 10 9 1 10 9 1 10 9 11 2 1 11 12 7 12 2 7 3 13 1 10 9 2
1 9
17 3 13 3 11 10 0 9 1 10 9 15 13 13 9 1 9 2
21 3 0 3 9 2 10 9 11 13 10 9 1 10 9 1 9 13 1 10 11 2
10 10 11 13 10 9 1 10 9 0 2
23 10 9 1 10 9 13 3 13 1 15 1 9 3 2 1 12 9 2 1 10 9 2 2
43 10 9 13 10 9 1 10 9 0 2 9 1 9 13 2 13 1 10 9 1 10 0 9 2 2 13 10 9 1 10 9 1 9 0 2 2 7 9 1 0 9 0 2
34 10 9 13 1 10 9 13 1 9 0 10 9 1 10 9 0 2 16 10 9 13 10 2 9 0 1 10 9 2 13 10 9 2 2
10 10 11 13 13 10 9 0 1 12 2
24 1 9 0 2 10 9 13 9 1 12 9 1 9 1 9 1 9 1 9 0 1 9 0 2
21 10 9 0 13 10 9 1 10 9 1 0 9 13 2 9 0 7 13 9 0 2
26 3 2 10 9 3 13 3 1 10 9 0 1 11 2 11 1 15 13 1 10 11 2 11 7 11 2
30 10 9 2 3 2 13 10 9 0 7 0 1 10 10 9 1 9 0 0 1 10 9 1 10 9 1 10 9 0 2
27 1 10 11 2 13 0 10 9 1 11 7 11 13 13 1 9 16 15 13 13 9 10 1 3 12 9 2
18 2 3 13 16 13 12 9 1 9 1 9 7 9 2 2 13 11 2
28 10 11 13 13 10 9 1 10 9 1 9 7 9 1 10 0 9 2 7 10 9 1 10 9 13 10 9 2
21 1 10 9 2 10 11 13 10 9 2 7 3 3 13 3 13 1 13 10 9 2
21 10 9 0 13 16 13 15 15 15 13 1 10 9 1 10 9 1 10 0 9 2
34 10 9 13 1 13 1 10 9 1 12 9 1 9 1 10 10 9 1 10 9 13 7 13 1 9 12 9 10 16 10 13 1 12 2
13 10 9 1 10 9 3 13 4 13 1 10 11 2
29 10 9 11 13 16 2 13 3 12 9 2 1 10 9 1 10 11 1 10 9 1 10 11 1 9 1 10 9 2
25 10 9 13 1 10 9 13 10 9 1 10 2 9 2 7 3 1 10 9 1 10 0 12 9 2
24 11 13 16 1 3 10 9 13 13 16 2 13 3 10 9 0 7 0 15 13 13 13 2 2
9 2 7 15 13 13 2 2 13 2
29 10 9 13 16 13 1 10 9 1 10 11 2 11 2 16 13 3 10 9 13 1 15 1 13 16 3 13 9 2
1 9
10 13 1 9 0 1 11 2 11 2 2
1 11
1 3
30 1 10 9 2 13 1 11 7 13 10 9 2 11 2 1 9 1 11 2 9 1 10 11 1 10 9 1 10 9 2
15 1 10 9 13 1 11 1 13 1 10 9 2 11 2 2
32 1 11 2 10 9 1 10 9 1 10 9 13 1 9 12 9 2 9 12 9 2 7 10 9 1 9 2 1 9 12 9 2
45 1 10 9 1 10 9 2 10 9 1 10 9 13 13 1 10 9 1 10 11 2 9 15 13 1 10 9 0 1 10 9 2 1 10 9 1 12 12 9 2 15 13 4 13 2
7 9 13 9 13 7 13 13
5 9 3 13 15 13
23 10 9 1 10 11 13 13 1 10 9 1 10 9 2 3 10 9 13 13 1 10 9 2
26 15 1 10 9 11 2 3 13 13 10 9 2 2 12 2 13 1 10 9 13 16 10 9 13 13 2
2 11 12
21 10 11 13 16 13 13 12 9 1 9 2 1 12 9 2 10 9 1 10 9 2
21 10 9 1 0 9 13 11 2 1 12 9 2 11 2 12 2 7 11 2 12 2
2 11 12
17 10 11 1 10 11 13 10 9 1 10 9 11 2 9 1 11 2
11 10 9 13 13 1 10 9 1 10 9 2
17 10 9 11 7 10 9 1 10 9 2 11 2 13 3 10 9 2
23 13 1 12 2 10 9 1 2 11 2 1 0 0 1 10 9 3 13 12 9 3 3 2
21 1 15 13 9 3 13 2 3 10 9 11 2 10 9 0 11 7 10 9 11 2
11 11 13 10 0 1 13 9 1 10 9 2
25 1 12 2 13 2 11 2 2 0 9 1 10 9 1 15 13 9 1 10 9 0 1 10 9 2
25 1 13 10 9 2 13 4 13 9 1 10 9 7 0 9 2 1 9 1 13 10 9 1 9 2
20 10 9 13 10 9 1 10 9 0 2 15 13 1 10 9 0 1 10 9 2
16 9 7 9 13 9 1 10 9 7 13 10 9 1 10 9 2
19 3 1 10 9 1 10 9 2 13 15 10 9 1 12 9 2 3 13 2
12 2 13 10 9 0 7 0 2 2 13 11 2
8 1 10 9 2 9 13 13 2
22 13 15 13 9 2 9 9 7 9 2 2 9 0 2 15 13 3 2 7 9 13 2
34 10 9 2 13 1 10 9 11 7 11 1 10 9 1 9 1 10 9 1 9 11 2 13 10 9 1 9 1 9 7 9 13 0 2
18 2 10 9 1 9 13 16 13 0 2 3 16 0 2 2 13 11 2
1 9
9 11 13 10 9 1 10 0 9 2
6 13 1 10 9 11 2
9 3 2 15 13 1 10 9 0 2
6 13 1 9 1 9 2
9 11 2 3 2 13 1 10 11 2
15 10 11 13 4 13 10 0 1 10 0 1 13 1 11 2
8 11 13 12 9 1 9 1 12
21 10 11 1 11 13 1 10 0 12 9 1 10 9 12 9 1 9 1 10 9 2
44 10 9 1 10 9 2 11 2 13 16 2 1 10 9 1 10 9 1 10 9 2 10 9 1 10 9 1 10 9 1 10 9 2 9 7 9 13 13 10 9 1 10 9 2
29 11 13 13 10 9 1 10 9 1 10 11 13 1 10 9 1 13 16 10 9 1 10 9 13 7 3 9 0 2
28 1 10 9 2 10 9 13 13 1 13 10 9 1 10 9 15 13 13 0 13 1 10 9 1 9 7 9 2
35 11 13 13 3 1 10 9 10 9 1 10 9 12 1 10 9 2 15 13 16 9 13 13 3 12 5 1 10 9 1 9 1 10 9 2
13 10 9 7 9 13 16 13 12 5 1 10 9 2
5 9 13 9 1 9
22 10 9 11 13 10 9 11 1 13 12 1 10 12 9 1 10 9 15 13 1 9 2
12 10 9 1 9 13 10 9 1 9 7 9 2
21 13 10 0 9 15 10 9 13 10 9 1 10 9 1 10 9 1 10 9 0 2
6 9 0 13 1 10 11
22 10 9 1 10 11 13 4 13 3 3 1 10 11 2 9 1 9 1 9 1 9 2
10 10 9 13 13 1 10 9 1 9 2
10 10 9 13 1 10 9 11 7 11 2
16 13 13 3 10 0 9 1 10 9 7 3 13 4 13 9 2
9 10 11 7 10 11 13 13 9 2
12 10 11 13 13 9 1 13 3 13 10 9 2
1 13
10 1 9 1 10 9 7 1 10 0 9
33 12 1 10 10 9 1 10 9 0 1 15 13 10 9 13 10 0 9 1 9 0 7 0 1 10 9 0 7 1 10 9 0 2
35 13 0 1 16 15 13 3 1 13 1 10 9 1 10 9 0 1 10 10 2 3 1 10 9 1 10 9 13 1 10 9 0 1 10 11
23 16 13 10 9 3 3 13 1 13 15 1 10 9 0 2 9 15 15 13 3 16 15 2
14 10 9 13 13 13 16 9 13 10 9 1 10 9 2
1 9
19 16 13 1 9 2 13 0 9 10 9 3 13 15 13 10 9 1 10 11
12 13 10 9 1 10 11 15 13 13 10 9 2
12 9 1 10 11 13 1 10 9 13 10 9 2
23 10 11 13 9 1 10 9 0 15 13 10 9 1 10 9 3 1 10 9 1 10 9 2
18 12 1 9 2 11 13 1 13 10 9 1 10 11 1 11 7 11 2
12 15 13 13 1 11 2 13 9 1 10 9 2
13 10 9 13 1 12 5 1 10 0 13 1 13 2
8 11 13 3 10 9 12 1 9
25 10 0 9 1 10 11 3 1 11 7 3 1 10 11 2 13 10 9 12 1 9 1 10 9 2
58 10 9 0 2 15 13 1 11 2 11 2 1 10 9 2 2 11 2 11 2 9 12 2 7 11 2 9 12 2 2 13 10 9 1 10 0 9 1 9 1 10 9 2 13 1 10 9 2 0 7 0 9 0 7 9 0 7 0
23 13 1 10 12 9 1 10 9 0 2 10 9 1 10 9 1 9 13 3 10 9 0 2
17 3 0 1 10 9 1 11 2 11 7 11 1 10 9 1 12 2
12 13 10 9 7 13 10 9 2 0 7 0 2
8 10 9 13 3 9 1 9 2
1 9
20 1 9 1 10 9 1 10 9 1 10 9 11 2 11 13 3 10 0 9 2
13 11 13 10 9 1 9 1 9 1 10 9 1 11
34 13 1 10 9 1 9 1 10 9 2 11 2 11 13 10 9 1 9 1 10 9 13 2 11 2 7 15 13 1 10 9 1 9 2
25 0 1 10 9 3 0 1 9 1 10 9 0 2 11 13 10 9 3 0 1 10 9 0 0 2
10 10 9 1 9 3 9 3 13 0 2
19 15 13 16 13 1 10 11 1 9 1 9 2 1 10 9 1 10 9 2
14 1 12 9 1 10 9 2 9 13 9 1 10 9 2
9 13 3 12 9 0 1 10 9 2
10 3 1 9 2 13 9 1 10 9 2
16 1 15 2 10 9 3 13 9 1 13 10 9 1 10 9 2
16 2 15 13 9 1 13 13 2 16 10 9 13 13 0 3 2
21 13 15 2 1 10 9 1 9 1 10 9 2 13 10 0 9 2 2 13 11 2
21 10 9 1 10 9 1 10 11 13 1 9 12 2 1 9 0 2 1 10 11 2
22 1 10 9 11 10 9 1 10 10 9 13 1 9 12 1 9 1 12 9 1 9 2
17 10 11 13 9 0 1 9 12 16 10 9 13 13 10 9 12 2
13 1 10 9 10 9 13 10 9 0 1 15 12 2
5 9 1 11 13 9
41 10 9 0 13 10 9 1 10 11 1 10 9 0 2 1 9 2 12 9 0 7 3 12 9 1 10 9 2 10 9 1 10 9 1 10 9 1 12 1 15 2
14 10 9 13 13 1 10 9 1 10 0 1 10 11 2
5 9 13 13 0 9
18 10 9 1 10 9 0 13 3 16 10 9 13 13 0 9 7 9 2
18 7 9 1 9 1 10 9 13 3 0 2 13 10 9 11 1 11 2
36 9 0 2 1 10 9 1 15 13 1 10 9 3 13 13 9 1 9 0 1 15 3 13 2 1 9 0 2 1 10 9 1 9 1 12 2
83 9 0 2 10 9 1 10 11 2 1 15 13 10 9 12 2 12 2 12 7 12 1 10 9 9 12 2 1 12 2 13 4 1 9 7 4 1 11 1 10 9 12 1 10 9 9 12 2 1 12 1 9 1 12 2 7 1 9 1 10 9 1 10 9 2 16 15 13 3 1 10 0 9 0 1 10 9 0 1 15 1 9 2
90 9 0 2 10 9 1 10 9 0 1 9 13 1 9 1 10 11 2 1 10 9 2 13 4 3 1 10 9 13 1 10 9 12 2 9 0 2 1 10 9 9 12 2 1 12 2 1 10 9 1 10 9 9 12 2 1 12 2 1 10 9 1 9 1 12 2 7 4 1 9 2 1 10 9 1 9 1 10 9 1 9 1 10 9 12 1 9 1 12 2
8 9 13 13 9 0 1 10 11
31 10 9 1 10 11 13 13 10 9 0 1 10 9 2 9 1 9 1 10 9 2 2 15 13 1 10 9 12 1 9 2
9 3 10 9 2 10 9 13 13 2
28 10 9 13 3 13 9 2 9 1 9 2 13 13 1 9 1 9 2 15 13 1 12 1 12 9 1 9 2
6 9 13 13 13 1 9
30 10 9 1 11 2 12 9 1 9 1 11 2 13 12 9 13 1 13 10 9 0 11 2 12 2 1 10 0 9 2
16 11 2 12 2 11 2 12 2 7 11 2 12 2 13 0 2
12 1 10 9 11 2 11 13 13 1 10 9 2
6 10 12 9 13 13 2
9 11 2 12 2 9 1 10 11 2
16 2 15 13 10 9 15 15 3 13 2 10 9 0 2 0 2
16 1 10 9 3 2 1 10 9 1 9 2 15 15 13 3 2
20 15 15 15 13 1 9 13 10 9 1 10 9 7 13 10 9 1 11 2 2
6 11 2 12 2 9 2
11 2 13 10 9 0 7 13 9 3 0 2
11 13 10 10 9 1 15 7 1 10 11 2
19 13 3 0 1 16 13 10 9 1 10 9 1 10 11 2 11 2 2 2
10 11 13 9 1 13 11 1 12 1 12
25 10 11 13 3 10 9 1 10 0 11 2 1 13 11 1 12 1 12 2 1 11 2 11 2 2
15 10 9 11 13 10 9 1 11 1 10 12 9 1 9 2
23 10 9 11 13 12 9 3 7 13 10 9 1 10 9 1 10 12 9 1 10 0 9 2
34 10 9 0 13 15 1 15 13 10 9 13 2 12 7 12 9 2 1 16 10 9 15 13 3 1 10 9 2 13 9 13 1 9 2
19 13 10 9 2 10 9 1 9 13 0 2 3 9 3 13 1 10 9 2
36 3 13 9 1 10 9 13 13 3 1 10 9 13 2 3 2 10 9 0 15 13 10 11 7 2 3 2 10 9 0 1 12 1 9 12 2
8 7 1 10 9 1 10 9 2
17 15 13 16 2 15 13 3 2 10 9 1 10 9 13 1 9 2
10 9 11 13 7 13 10 9 1 10 9
39 10 9 7 9 0 1 9 11 7 10 12 9 13 10 9 1 3 1 10 9 1 11 2 3 1 13 13 10 9 1 10 9 1 10 9 11 1 11 2
23 10 12 9 13 9 1 10 11 2 11 2 2 9 0 15 13 1 10 9 1 10 9 2
25 15 15 13 3 7 1 10 9 1 10 9 1 9 1 10 9 1 9 9 1 9 1 10 9 2
6 11 13 9 1 10 9
21 10 9 11 13 3 16 10 9 0 10 0 1 12 13 9 1 9 1 10 9 2
21 10 9 13 1 10 9 1 10 9 2 11 2 13 1 10 9 13 1 10 11 2
23 10 9 13 1 10 9 1 13 2 13 7 13 10 9 1 9 1 10 9 1 10 9 2
26 11 13 16 10 9 1 10 9 13 10 9 1 12 9 2 15 3 13 13 1 10 9 1 10 9 2
22 1 11 2 10 9 1 10 9 13 1 10 9 1 10 9 13 10 9 1 10 9 2
21 10 9 1 10 11 2 9 11 2 13 16 13 2 9 13 1 13 15 3 2 2
17 10 9 2 3 2 3 13 15 1 13 10 9 1 10 9 0 2
19 10 9 11 13 10 9 15 3 13 10 9 1 13 10 9 7 9 11 2
35 2 15 13 10 0 9 2 7 13 10 0 9 2 2 13 11 2 15 13 10 9 1 11 2 9 1 9 0 2 7 1 10 9 11 2
7 11 2 3 2 7 13 2
10 11 2 10 9 13 13 13 10 9 2
3 0 1 13
26 11 2 9 1 10 11 2 13 3 13 4 13 1 10 9 1 10 9 1 10 9 1 13 10 9 2
7 10 9 0 13 13 3 2
8 10 9 11 13 9 1 9 2
2 9 0
27 10 9 1 10 11 13 16 10 9 11 2 9 1 10 9 2 13 9 1 10 9 7 9 1 10 9 2
17 1 9 1 10 9 1 10 9 2 15 13 16 3 13 10 9 2
32 15 3 3 13 10 9 7 10 9 1 10 15 13 13 11 3 13 9 1 2 9 0 13 2 1 15 15 13 1 10 9 2
28 10 0 9 0 13 13 10 9 1 10 9 1 3 12 12 9 1 10 11 13 1 12 1 10 9 1 11 2
28 1 10 9 2 11 13 10 9 1 9 1 9 0 1 10 9 7 13 10 0 9 1 15 13 1 10 9 2
8 9 0 13 13 9 1 10 9
32 9 1 0 9 1 9 0 7 0 13 15 13 2 1 13 10 9 2 1 13 10 9 1 10 9 2 13 10 9 7 9 2
25 15 2 3 2 13 13 1 9 10 10 9 0 7 0 15 13 13 10 9 0 7 1 0 9 2
7 10 9 13 0 2 13 2
12 10 9 0 15 13 1 10 9 13 0 9 2
8 15 3 15 13 1 10 15 2
39 7 15 1 15 13 9 1 3 13 10 9 1 10 9 1 10 9 7 1 13 13 1 10 9 2 7 1 13 1 10 9 1 9 1 10 9 1 9 2
10 3 7 1 10 12 9 13 10 9 2
14 15 1 9 13 0 2 7 13 1 11 7 13 3 2
24 15 1 15 12 3 13 0 2 7 13 1 10 9 3 13 1 10 9 7 3 13 13 9 2
9 3 9 1 13 2 16 13 0 2
10 13 10 11 1 11 15 13 10 9 2
16 1 9 1 11 7 11 7 9 3 1 10 9 1 10 11 2
25 1 9 13 1 10 9 13 1 11 2 11 13 10 9 1 10 2 9 2 1 10 9 1 11 2
16 10 9 2 13 3 1 10 9 0 2 13 10 9 1 9 2
24 10 9 0 13 13 2 13 3 10 9 13 1 2 11 2 1 11 7 2 11 2 1 11 2
10 10 11 13 3 1 10 9 1 11 2
14 3 10 9 0 13 1 10 9 1 10 2 11 2 2
14 3 2 13 0 10 9 1 10 10 9 1 10 9 2
12 1 10 9 13 10 9 2 11 2 1 11 2
22 10 0 2 11 2 13 2 11 2 1 10 9 11 7 2 11 2 1 10 9 11 2
11 10 10 9 13 1 10 2 9 2 13 2
80 2 11 2 1 11 2 2 11 2 1 11 2 2 11 2 2 1 11 2 2 11 2 1 11 2 2 11 2 1 11 2 2 11 2 1 11 2 2 11 2 1 11 2 2 11 2 1 11 2 2 11 2 1 11 2 2 11 2 1 11 2 2 11 2 1 11 2 2 11 2 1 11 7 10 9 0 2 11 2 2
6 11 13 9 13 1 9
16 10 9 15 10 9 3 13 3 13 10 9 2 7 10 9 2
8 10 9 0 13 10 0 9 2
27 10 9 1 10 0 9 13 10 9 11 1 10 9 0 2 1 10 9 1 12 9 2 1 10 0 9 2
16 15 0 13 13 1 10 9 1 16 3 15 13 1 10 9 2
35 1 10 9 2 3 1 10 9 2 9 1 10 9 1 10 0 9 1 11 2 11 2 11 2 11 7 9 2 13 10 9 1 10 9 2
38 3 9 1 10 9 1 10 9 2 10 9 0 13 10 9 1 10 11 2 10 9 1 9 0 15 13 13 3 1 10 9 1 9 3 13 1 9 2
27 2 13 13 12 9 1 10 9 2 13 3 9 1 9 1 9 7 15 13 9 1 9 2 2 13 9 2
27 1 9 2 10 9 13 1 10 9 1 15 13 1 12 9 0 15 3 13 1 10 9 2 11 7 11 2
31 10 9 13 1 10 9 10 9 3 0 2 15 13 1 15 15 13 1 10 9 0 10 9 0 2 3 13 1 10 9 2
6 10 9 13 3 0 2
28 10 9 13 10 9 1 9 7 1 9 11 1 10 9 1 10 9 13 7 13 10 9 1 9 1 10 9 2
28 1 10 9 13 2 10 9 1 10 11 13 2 9 2 10 9 1 10 9 7 13 2 9 2 10 9 0 2
18 10 9 13 13 10 9 1 10 9 7 13 10 9 1 10 9 0 2
15 10 9 1 10 9 1 10 9 13 1 9 12 1 9 2
9 15 1 15 13 0 2 9 12 2
9 1 9 2 9 13 2 0 2 2
16 10 9 1 10 9 1 10 11 13 13 1 10 9 1 11 2
14 3 1 10 9 1 10 9 2 7 1 10 9 0 2
10 9 2 9 2 9 1 9 7 9 2
27 10 12 9 3 13 1 4 13 2 7 13 10 9 2 13 1 9 1 10 9 13 0 2 7 3 13 2
26 1 10 9 2 1 11 2 12 9 1 10 9 1 10 11 2 2 11 13 10 9 1 11 7 11 2
18 13 16 11 13 0 3 7 16 11 13 0 7 16 3 13 1 13 2
20 1 10 9 2 13 12 9 1 10 9 1 10 9 2 3 11 13 1 13 2
17 3 15 13 2 1 10 9 2 9 1 10 9 13 13 10 9 2
11 13 10 9 1 10 2 9 1 10 9 2
27 10 9 13 2 3 2 10 9 1 13 9 3 13 1 10 9 1 13 2 7 3 3 13 15 15 13 2
18 3 10 9 1 10 9 1 15 13 13 1 10 9 1 9 1 9 2
41 10 9 3 13 1 10 2 9 1 10 0 9 2 2 15 13 13 3 1 10 9 0 2 7 3 10 10 9 1 15 10 9 13 10 9 13 1 10 10 9 2
23 16 10 9 13 10 9 7 9 1 10 9 1 10 9 7 16 2 3 2 13 1 15 2
15 16 3 13 15 2 1 3 13 13 10 9 1 10 9 2
16 11 13 1 10 9 1 11 7 11 2 9 2 1 10 9 2
8 13 12 9 0 7 12 0 2
27 15 13 16 10 9 11 7 11 2 1 10 11 2 13 13 10 9 0 2 1 9 1 12 1 10 11 2
38 9 1 11 2 11 13 12 9 3 10 9 2 10 9 7 12 9 13 1 11 2 0 1 11 2 1 10 11 2 1 13 3 9 1 10 9 11 2
33 11 2 15 13 13 9 1 11 2 1 10 11 2 3 13 1 12 9 2 13 9 1 15 13 9 7 9 1 13 1 10 11 2
31 1 11 2 9 1 10 11 1 10 11 2 11 2 2 10 9 15 13 1 9 1 10 9 1 13 9 0 1 10 11 2
27 3 1 11 2 10 9 13 0 10 9 1 10 9 1 10 9 16 10 11 13 10 9 0 1 9 0 2
20 1 10 9 1 3 2 1 10 9 2 9 2 13 2 10 9 1 10 11 2
21 10 9 13 10 9 1 16 10 10 9 13 0 1 13 10 9 0 1 10 9 2
8 3 2 13 13 3 12 9 2
16 15 1 0 9 13 1 10 11 2 11 2 7 1 10 11 2
4 9 13 12 9
12 10 11 2 11 2 13 3 12 9 1 9 2
18 12 1 10 9 11 2 12 1 10 11 7 10 11 2 1 10 11 2
20 13 13 10 11 2 10 11 7 10 11 2 15 3 13 4 1 13 1 9 2
27 2 10 9 1 10 9 1 9 0 13 10 9 1 15 13 1 10 15 2 3 10 9 13 12 9 3 2
20 15 13 10 9 1 9 1 9 12 5 0 1 10 15 2 2 13 10 9 2
24 10 9 1 10 9 1 9 1 10 9 3 13 0 9 1 10 9 2 9 2 7 10 9 2
22 10 9 1 9 1 9 11 2 12 2 13 1 12 9 2 13 10 9 1 10 9 2
11 2 15 13 9 1 10 9 1 10 9 2
3 13 13 2
4 13 9 2 2
14 10 9 13 10 9 1 10 9 1 9 1 10 9 2
16 2 13 13 1 10 9 2 1 10 9 7 10 9 10 2 2
23 10 9 11 2 13 1 9 13 16 10 9 0 13 13 0 13 1 10 9 1 10 9 2
30 2 16 10 9 13 10 0 9 1 10 9 1 10 9 1 10 9 1 9 0 1 9 13 9 1 15 2 2 13 2
15 15 16 15 13 15 13 10 9 1 10 9 0 2 13 2
27 10 9 1 10 11 2 11 1 10 11 2 13 13 10 0 9 1 15 13 13 1 10 11 1 10 11 2
14 10 9 13 0 2 7 13 10 0 9 1 9 12 2
20 15 13 1 9 0 2 13 13 10 11 2 11 2 3 9 1 10 11 2 2
21 10 9 13 1 9 1 9 3 2 1 9 12 2 7 9 13 2 9 12 2 2
11 2 11 2 13 9 13 1 10 9 1 9
5 1 10 9 1 9
27 13 15 1 9 1 10 12 9 15 11 13 1 10 11 2 1 12 9 1 11 2 11 2 11 7 11 2
31 3 13 9 1 9 2 3 13 9 0 9 2 3 13 9 0 2 3 13 9 1 10 9 0 2 3 13 13 1 9 2
17 2 13 3 13 1 10 9 9 0 1 12 5 2 2 13 11 2
29 10 9 15 13 13 13 10 9 1 10 9 1 9 2 3 2 2 15 3 13 1 3 12 5 1 10 9 13 2
10 10 9 13 13 1 12 5 2 13 11
37 10 9 10 2 1 10 9 2 10 0 0 15 13 1 10 9 1 10 0 9 1 10 9 2 13 1 10 10 9 1 9 15 13 1 10 9 2
37 1 10 9 1 10 9 1 2 11 2 2 13 10 9 1 12 1 10 0 9 0 0 2 3 13 15 0 1 13 10 9 13 3 1 10 11 2
1 9
20 10 9 1 9 1 10 11 13 13 9 1 10 9 1 0 9 1 9 0 2
20 13 13 9 1 9 1 10 9 1 10 9 11 3 0 1 12 1 12 9 2
38 10 9 13 10 9 1 10 9 12 9 13 7 9 12 9 1 9 1 10 9 2 13 1 10 0 9 2 7 9 12 9 15 10 9 13 1 13 2
47 11 13 16 1 10 9 12 9 10 9 13 1 13 9 12 9 1 9 1 9 0 2 7 9 12 9 1 9 1 9 1 9 7 10 9 12 9 1 9 1 9 1 9 1 10 9 2
4 11 13 10 9
15 10 9 1 9 1 10 11 13 12 5 1 12 7 12 2
18 10 9 1 10 9 13 13 1 10 9 1 10 9 1 10 9 0 2
20 1 12 1 12 2 10 9 1 9 0 13 1 12 9 1 12 9 1 9 2
17 0 9 2 3 13 13 1 10 9 1 10 9 1 13 10 9 2
17 10 9 1 10 9 2 3 3 2 3 13 10 9 1 10 9 2
6 11 13 9 1 9 2
8 11 13 9 11 1 15 1 11
35 10 9 11 13 3 1 10 9 1 10 9 0 1 10 9 12 1 12 7 10 0 9 1 10 9 11 1 10 9 1 10 9 1 11 2
27 10 9 13 1 10 9 1 10 9 1 10 9 1 9 2 9 7 9 7 9 1 10 9 1 10 9 2
25 10 9 1 10 11 2 11 2 13 16 10 9 13 13 12 5 1 9 1 10 9 1 10 11 2
43 1 10 9 1 10 11 2 11 2 10 9 13 16 10 9 1 9 7 9 13 10 9 10 10 9 0 1 12 2 9 1 15 13 13 10 0 9 1 9 1 9 0 2
10 10 9 13 1 9 12 9 1 12 2
25 1 10 0 11 2 9 1 10 11 2 9 1 10 9 1 10 11 2 2 9 7 9 13 13 2
16 2 13 1 9 15 13 10 9 7 13 10 9 2 3 11 2
17 11 13 13 2 7 1 10 9 15 3 13 2 2 13 10 9 2
40 10 0 2 1 10 9 1 10 9 2 13 1 10 9 1 10 11 2 9 3 0 16 10 10 11 13 3 9 0 2 15 15 13 9 2 1 10 0 11 2
41 3 7 3 1 15 2 13 10 9 1 10 11 2 15 13 1 10 9 1 10 9 2 7 13 10 9 0 2 7 13 1 10 9 1 0 1 10 9 1 9 2
10 3 2 10 0 13 13 10 0 9 2
6 7 13 13 3 15 2
76 13 13 10 9 15 15 13 1 10 9 15 13 10 0 9 1 10 9 1 10 9 2 3 10 9 1 11 13 10 9 2 1 12 2 12 2 3 12 9 13 10 9 2 15 2 1 10 9 2 3 13 7 9 0 1 10 9 2 7 9 0 1 10 9 2 10 9 13 1 11 2 10 0 9 0 2
9 10 9 13 13 1 9 7 9 2
4 13 0 9 2
18 9 1 9 3 3 13 0 2 1 3 10 9 2 9 2 9 2 2
29 1 9 1 10 9 2 13 15 16 10 9 15 10 11 13 1 10 9 3 13 1 10 9 2 7 1 10 9 2
65 10 9 13 2 3 2 1 10 9 1 16 10 9 0 1 10 11 15 13 1 15 15 13 1 12 9 2 1 10 9 0 15 15 13 9 7 1 10 9 0 15 13 2 0 1 9 0 2 10 9 1 13 1 10 9 1 9 1 10 9 1 10 0 9 2
15 10 9 0 3 13 13 1 11 10 9 1 13 10 9 2
24 3 3 15 13 16 13 10 0 9 1 10 9 2 15 13 3 13 7 3 13 1 10 9 2
34 16 15 13 2 3 2 10 10 9 1 10 9 2 3 3 3 10 9 13 1 10 9 1 10 9 2 7 1 10 9 1 10 9 2
19 16 3 13 1 10 9 1 10 9 0 2 3 13 13 1 3 1 9 2
7 2 10 9 13 13 3 2
11 7 3 13 15 1 13 1 10 9 2 2
23 10 9 13 13 10 9 1 10 9 2 13 10 9 1 10 9 0 1 9 7 13 9 2
9 9 1 10 9 13 0 2 13 9
18 9 1 10 9 7 9 1 10 9 13 0 7 3 0 2 1 11 2
23 10 9 7 9 0 13 1 10 9 1 10 0 9 1 10 9 1 10 9 2 11 2 2
22 1 10 9 1 3 2 13 3 12 9 13 1 10 9 1 11 2 10 0 1 11 2
18 10 9 1 10 9 1 3 1 11 7 11 7 11 13 13 1 11 2
5 2 13 1 15 2
13 7 3 13 13 16 10 9 13 0 10 9 2 2
16 2 13 13 16 15 15 13 2 7 16 15 13 1 10 9 2
16 7 3 13 9 3 10 2 16 10 9 3 13 0 7 0 2
5 13 3 10 9 2
12 3 15 13 13 10 9 3 15 13 10 9 2
28 16 15 13 13 15 2 13 13 3 10 9 2 3 15 1 10 9 1 10 9 2 3 13 13 10 9 2 2
12 2 15 13 13 2 2 13 11 1 10 9 2
16 2 13 16 13 3 1 10 9 0 1 13 1 10 9 2 2
19 10 9 13 10 10 9 0 1 10 9 1 13 10 9 1 10 0 9 2
52 3 1 10 9 2 0 9 1 10 9 0 3 13 13 10 9 0 2 9 1 10 9 7 1 10 9 2 13 1 10 9 0 2 13 1 10 9 10 9 1 9 0 7 0 1 15 15 10 9 13 13 2
30 9 0 2 9 1 9 1 10 9 2 9 1 9 7 9 3 13 10 9 1 10 9 0 1 10 9 1 10 9 2
40 10 9 1 9 7 1 9 15 3 13 1 12 9 13 1 13 10 9 2 10 9 2 10 9 0 1 10 0 9 1 10 9 0 1 10 10 9 1 9 2
26 11 2 12 2 9 2 13 9 1 10 11 2 11 2 7 9 1 10 11 1 10 11 2 11 2 2
24 11 13 1 11 2 3 2 1 10 9 15 13 13 2 15 13 1 10 9 3 0 1 11 2
29 11 13 11 1 15 13 3 1 9 7 2 3 2 13 10 9 13 1 10 10 9 15 15 13 13 1 10 9 2
25 11 2 11 2 13 3 3 1 10 9 1 11 7 3 13 10 0 9 1 9 2 13 13 1 11
18 10 9 13 12 9 2 1 10 9 1 12 9 2 7 13 9 12 2
14 10 0 9 1 10 9 13 9 12 7 12 1 9 2
2 3 13
7 11 13 0 0 1 11 2
17 10 12 9 1 9 13 1 11 7 13 1 10 9 1 12 9 2
11 11 2 12 9 2 13 9 1 12 9 2
21 10 9 2 9 7 13 1 13 9 2 13 15 2 3 2 1 13 1 9 13 2
34 3 13 13 16 10 9 13 0 2 7 3 16 13 10 0 9 0 2 9 2 1 13 10 0 3 3 1 13 15 15 13 10 9 2
26 10 9 0 2 0 7 0 3 13 1 15 13 2 16 10 9 1 10 9 0 3 13 1 9 0 2
22 16 10 9 0 13 3 0 15 13 2 7 13 16 3 13 1 13 3 0 1 9 2
27 11 2 12 2 9 1 9 0 1 10 11 2 11 2 2 13 0 1 10 11 1 10 11 2 11 2 2
45 12 9 13 9 3 1 10 9 2 1 10 9 2 9 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 7 11 2
14 1 10 9 0 13 0 11 2 11 2 11 7 11 2
7 10 9 0 13 1 11 2
23 1 10 9 13 13 9 1 10 9 1 10 9 1 9 1 9 1 11 2 1 10 11 2
8 13 10 9 1 9 1 10 11
19 9 1 10 9 1 10 9 7 9 1 10 11 13 10 9 0 2 9 13
8 10 9 0 13 3 13 3 2
10 10 11 2 11 2 13 9 12 9 2
15 13 10 0 9 1 0 1 9 0 2 9 12 9 2 2
22 10 9 13 1 10 9 1 9 2 1 10 11 2 1 9 1 9 1 9 1 9 2
40 10 9 11 13 1 9 1 10 10 9 7 9 1 10 9 2 7 13 1 9 1 12 5 2 13 10 9 1 10 11 3 0 1 10 9 1 10 9 0 2
30 13 10 9 1 10 15 13 1 12 2 1 10 11 2 3 2 13 2 12 5 1 9 1 10 9 0 1 9 0 2
27 10 9 13 1 10 9 1 13 10 9 1 13 10 9 0 1 10 9 2 7 13 10 9 1 0 9 2
5 10 9 13 13 2
22 10 9 0 1 10 11 13 13 1 9 12 1 10 9 1 9 1 10 0 9 12 2
20 10 9 11 0 13 1 12 9 2 1 9 1 9 1 12 5 1 10 9 2
2 13 11
42 13 10 9 11 3 10 9 1 9 1 12 7 12 9 3 13 13 10 9 1 9 13 1 10 15 1 11 1 10 9 2 1 10 9 1 10 9 7 1 10 9 2
18 11 13 10 9 1 9 2 15 13 1 9 7 9 1 10 9 13 2
20 10 9 13 10 3 0 9 1 10 0 9 11 2 1 10 11 2 1 11 2
2 13 3
27 11 2 9 1 10 9 0 1 11 2 13 13 1 10 11 10 0 9 15 13 13 15 13 1 10 11 2
21 13 15 1 10 11 10 9 1 9 11 7 9 11 1 10 0 9 13 1 11 2
21 13 10 9 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 7 11 2
9 3 13 0 11 2 11 7 11 2
20 10 9 13 13 13 10 9 1 2 9 1 9 2 1 10 9 1 10 9 2
21 10 9 1 9 1 9 2 1 10 9 2 13 1 10 9 1 11 7 10 11 2
25 1 10 9 2 10 9 1 11 2 11 2 13 16 13 1 13 1 10 9 1 16 13 10 9 2
21 3 2 15 13 1 10 9 7 15 13 0 1 13 15 2 3 1 10 9 2 2
38 1 10 9 1 3 2 1 10 9 1 10 11 2 9 1 10 9 2 11 13 16 2 3 13 13 7 13 9 10 9 1 9 2 13 1 10 11 2
18 11 10 11 13 15 13 1 10 9 1 10 10 9 2 1 9 0 2
20 11 3 13 10 9 16 13 10 9 10 10 2 15 13 10 9 1 10 11 2
10 13 10 9 7 13 10 9 1 11 2
17 13 13 9 13 1 9 2 9 2 9 2 10 10 9 1 9 2
19 2 3 13 13 9 2 9 13 2 9 1 9 7 3 13 13 10 9 2
12 13 16 10 2 9 2 13 10 0 9 2 2
6 10 9 13 12 9 2
24 11 13 9 0 2 13 1 10 9 1 10 9 2 7 13 13 1 10 9 1 10 10 9 2
22 1 10 11 2 3 10 9 1 9 13 0 1 10 9 2 13 3 9 7 9 13 2
18 15 13 13 3 1 10 9 0 7 0 1 10 9 1 13 10 9 2
7 9 13 10 9 1 10 9
17 9 9 13 9 12 1 9 12 1 10 0 1 12 9 13 1 11
30 1 10 9 13 2 10 9 1 9 0 13 13 1 10 9 2 10 9 0 13 9 0 1 10 9 0 1 10 9 2
17 9 12 0 2 10 0 11 13 10 9 1 9 12 1 12 9 2
29 12 9 3 2 10 11 2 13 10 9 1 9 12 1 10 9 1 9 1 10 12 9 0 15 13 13 1 9 2
20 1 10 11 1 11 2 10 10 9 13 3 12 9 2 10 9 1 10 9 2
9 10 9 13 13 10 9 0 12 2
18 10 9 1 10 11 13 1 10 11 2 12 2 1 10 9 1 9 2
7 11 13 1 10 9 1 11
14 11 13 1 10 9 1 3 1 11 2 13 1 11 2
15 10 9 13 10 9 15 15 13 1 3 13 1 10 11 2
29 2 3 13 9 2 9 2 9 0 7 9 0 3 1 12 9 2 2 13 10 9 11 2 15 13 3 1 11 2
16 10 9 2 13 15 2 13 9 13 7 3 13 13 1 9 2
13 15 13 16 10 9 1 10 9 3 13 10 9 2
13 11 13 16 10 9 15 13 3 3 1 15 13 2
14 1 15 2 10 3 12 9 0 13 13 1 0 9 2
6 9 0 13 1 12 9
19 10 9 1 10 9 11 2 11 7 11 13 0 12 9 2 1 9 0 2
25 13 0 13 10 12 9 1 10 9 1 10 9 0 1 12 9 2 13 15 10 9 1 10 9 2
13 15 13 1 10 9 1 12 5 1 10 9 0 2
2 9 13
15 10 9 11 13 10 11 1 10 9 11 2 13 1 11 2
43 10 9 1 9 1 10 11 15 13 1 10 9 1 10 11 2 9 0 1 11 2 7 1 10 11 2 11 1 10 11 2 13 10 9 1 10 11 2 9 0 0 0 2
9 10 9 7 10 9 0 13 9 2
16 3 2 10 9 11 2 0 1 10 9 2 13 1 10 11 2
3 9 2 9
2 9 13
20 10 9 0 13 10 9 1 10 9 3 0 7 13 16 10 1 10 9 13 2
42 16 3 3 13 4 3 13 2 10 9 1 10 9 1 10 9 11 13 15 3 3 3 13 2 13 9 1 16 10 9 13 1 13 1 9 1 10 0 9 1 13 2
42 10 0 9 15 13 1 11 3 13 16 10 11 13 10 9 1 9 13 1 10 11 1 11 7 16 2 1 10 9 2 10 9 1 11 13 1 10 9 1 10 11 2
5 13 10 9 0 2
51 3 10 9 13 1 10 9 13 3 10 9 1 10 11 15 13 13 10 0 9 11 1 9 1 9 1 10 9 2 3 3 13 9 13 9 1 16 10 9 13 3 13 10 9 1 11 2 1 10 9 2
7 9 13 0 9 1 10 9
44 9 1 10 11 1 10 11 1 10 9 1 9 1 10 9 13 16 10 11 13 10 9 1 1 12 5 1 10 9 1 10 9 15 13 4 13 1 13 10 9 1 10 9 2
15 10 9 13 15 1 10 9 1 10 9 0 1 10 9 2
10 10 9 13 10 11 7 3 13 9 2
10 9 1 11 13 2 13 2 1 10 11
27 10 11 2 11 2 13 13 10 0 9 1 10 10 9 2 10 9 1 10 9 1 10 9 2 10 11 2
45 10 9 2 13 1 12 9 1 10 11 1 10 11 1 13 10 10 10 9 1 9 2 13 13 10 0 9 1 9 1 9 2 13 1 9 1 9 13 1 10 9 1 10 9 2
22 10 9 3 13 1 10 11 13 9 0 7 9 1 9 2 13 3 11 2 11 2 2
31 1 15 13 10 9 1 10 9 1 10 11 2 10 11 13 13 1 10 9 2 13 9 7 9 1 10 9 1 10 9 2
1 9
31 10 9 11 13 9 2 9 2 9 2 9 2 7 13 1 9 1 10 9 1 12 1 12 7 1 12 1 12 1 9 2
15 13 1 10 9 11 2 1 11 2 1 12 9 1 11 2
19 11 13 13 10 9 1 10 11 1 13 10 9 1 10 11 7 13 11 2
19 10 9 13 16 10 11 13 10 9 2 1 13 10 9 1 9 0 2 2
36 11 2 15 13 0 7 15 13 9 1 10 11 2 13 16 10 9 1 10 9 2 1 10 9 13 16 10 9 13 3 0 1 10 9 2 2
31 1 10 9 13 1 10 11 2 10 9 1 10 9 13 16 2 10 9 1 11 13 1 10 9 0 2 1 10 10 9 2
18 7 10 9 1 10 9 1 0 7 0 1 10 9 9 3 15 13 2
15 1 10 9 2 15 13 3 10 9 13 10 9 0 2 2
4 2 13 9 2
19 10 9 0 13 4 13 1 12 9 0 16 10 9 13 0 2 2 13 2
9 10 9 13 4 13 1 9 0 2
9 3 13 9 0 1 10 9 0 2
4 11 2 9 2
3 11 1 9
32 10 9 0 2 11 2 13 10 9 1 11 2 11 2 2 10 0 9 1 10 9 15 13 10 9 1 9 11 2 11 2 2
21 13 1 10 9 0 1 11 2 10 0 13 3 1 10 9 11 2 11 7 11 2
6 10 9 13 1 11 2
34 1 11 2 13 13 10 9 10 9 1 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 7 11 2
20 10 9 13 4 13 3 1 10 9 0 2 13 3 10 9 0 1 9 0 2
17 15 13 12 9 3 3 16 11 13 10 9 12 9 3 2 3 2
21 1 10 9 2 10 9 1 11 13 13 3 12 9 1 3 2 16 13 12 9 2
23 10 9 13 13 1 10 9 1 9 2 7 10 9 13 1 13 1 10 2 0 9 2 2
12 15 13 1 10 9 1 10 9 9 7 9 2
33 10 9 9 13 13 1 10 9 7 2 3 2 3 13 13 1 10 9 2 10 10 9 1 10 9 13 1 10 9 1 10 9 2
24 10 9 1 10 9 13 0 1 10 9 1 10 0 3 13 9 1 10 9 2 7 3 9 2
18 15 1 10 9 13 0 9 3 2 15 13 9 1 10 9 3 9 2
22 10 9 13 3 13 10 9 1 9 7 13 1 10 9 1 10 9 2 1 10 11 2
12 3 13 10 9 0 2 0 2 0 7 0 2
15 10 9 3 13 10 9 1 9 2 13 10 9 1 9 2
87 13 1 10 9 2 10 9 13 1 10 9 1 10 9 2 10 9 13 1 10 9 1 10 9 2 1 10 9 1 10 9 2 11 13 10 9 1 10 11 2 1 10 11 3 0 7 3 0 2 13 1 10 9 2 1 10 9 2 1 10 9 2 1 10 9 2 1 10 9 2 1 10 9 13 1 10 0 9 1 10 9 0 1 0 9 0 2
26 6 2 9 11 2 13 15 1 10 9 1 3 9 2 13 15 10 9 1 10 9 7 1 10 9 2
40 3 2 1 10 9 3 15 13 10 9 2 15 15 13 9 1 10 10 9 2 10 0 9 13 1 10 9 1 10 9 2 1 15 13 10 9 7 10 9 2
20 15 13 16 3 10 9 13 9 7 15 13 3 2 1 10 9 1 10 9 2
2 11 12
11 10 11 13 9 12 10 11 2 1 11 2
24 10 9 13 1 10 9 1 15 13 11 2 9 1 10 9 2 11 2 2 10 9 3 0 2
5 10 9 13 13 2
1 11
9 10 11 13 13 3 2 1 11 2
36 10 9 1 10 9 2 9 11 2 11 2 2 13 16 10 9 13 13 10 9 1 9 0 2 1 10 9 1 10 9 7 9 1 10 9 2
27 10 9 13 1 9 12 9 2 0 1 9 12 9 2 1 9 12 9 1 10 9 0 2 15 13 13 2
25 10 0 9 1 10 9 1 9 13 10 9 1 9 0 2 1 9 1 10 9 2 1 12 9 2
39 10 9 1 12 9 0 1 10 11 1 10 9 1 10 9 1 9 1 11 2 11 2 13 1 13 3 1 11 1 10 9 1 13 1 13 10 9 0 2
22 12 9 1 12 9 1 10 9 1 10 11 3 13 3 1 10 11 1 10 10 9 2
38 10 9 1 10 11 1 10 9 2 11 2 13 16 13 13 1 12 9 1 10 13 9 13 1 11 10 9 13 1 10 9 0 13 1 10 10 9 2
35 10 9 13 13 9 13 1 12 9 1 11 3 9 12 9 2 9 15 13 1 10 11 2 11 2 7 11 2 11 2 13 1 10 9 2
6 11 0 15 13 1 9
23 11 2 1 10 9 11 7 11 2 9 7 9 1 10 11 2 13 10 9 1 10 11 2
39 1 10 0 9 2 10 9 13 12 1 10 9 2 0 1 10 9 1 9 1 10 9 2 1 13 10 11 1 10 9 0 2 1 10 11 2 1 12 2
42 11 2 9 1 10 11 2 13 10 9 0 7 10 3 12 9 1 9 1 13 10 9 1 10 9 1 10 0 2 3 1 10 9 0 1 10 11 1 10 0 9 2
6 13 13 1 10 0 2
20 1 10 9 2 11 3 13 10 9 0 15 15 13 1 10 9 1 10 9 2
15 13 10 11 3 1 10 9 1 9 1 9 1 10 9 2
23 2 16 13 0 13 2 10 11 3 13 10 9 0 2 2 13 11 2 9 1 10 11 2
27 13 16 10 0 9 15 2 3 1 10 11 2 13 9 0 2 15 13 1 13 0 9 13 1 10 9 2
18 1 10 9 1 10 0 9 2 11 13 10 9 1 10 9 0 11 2
12 1 12 9 2 13 2 11 2 2 1 11 2
18 10 9 11 13 1 10 11 1 9 1 10 9 11 7 1 10 11 2
4 11 13 1 9
37 1 10 9 2 9 12 2 10 11 2 11 2 13 10 9 0 1 9 1 10 11 2 1 10 11 2 9 0 2 2 1 10 11 1 10 11 2
14 10 9 13 13 3 9 1 9 7 9 1 10 11 2
3 11 13 9
4 9 1 10 9
37 9 1 10 9 1 11 1 10 0 9 11 13 15 1 10 9 1 10 9 1 10 9 15 13 9 1 10 11 1 11 7 1 10 11 1 11 2
36 11 13 1 12 5 1 12 5 1 10 9 2 12 9 0 1 9 2 7 1 12 5 1 12 5 1 10 9 1 10 11 2 12 9 2 2
35 12 1 9 1 12 2 10 11 2 1 10 11 2 13 1 10 9 3 3 1 13 1 10 9 0 1 11 2 13 10 9 1 12 9 2
7 9 1 0 1 12 2 12
22 12 1 9 1 12 2 10 9 0 11 2 1 10 11 13 1 10 9 0 1 11 2
15 1 10 12 9 7 9 15 13 1 10 9 2 12 13 2
17 9 15 10 9 1 10 9 1 10 11 1 10 9 1 10 9 2
18 9 0 3 3 15 13 1 9 1 9 2 1 13 1 9 7 9 2
6 9 13 9 0 1 11
32 10 2 11 2 13 10 9 0 1 10 9 1 10 11 1 3 2 1 10 9 1 10 9 7 10 9 1 10 9 1 9 2
23 1 10 9 1 9 12 2 10 9 13 15 13 1 10 9 1 10 9 1 9 1 9 2
17 15 15 13 9 2 13 13 1 10 9 13 1 10 9 1 9 2
31 10 9 13 13 1 10 11 1 12 9 7 13 12 9 1 9 1 10 9 1 10 9 2 1 9 0 2 9 7 9 2
10 11 13 10 9 1 10 0 9 1 11
11 9 13 9 1 0 1 10 2 11 2 2
30 1 10 9 0 1 10 9 2 10 9 11 13 13 9 2 1 9 0 2 1 10 9 15 13 10 13 2 11 2 2
1 9
8 9 1 9 1 10 9 13 3
16 13 9 1 9 0 10 9 1 10 9 1 10 9 2 9 2
7 11 2 11 7 11 13 2
3 13 11 2
5 15 15 13 0 2
6 2 0 2 7 0 2
20 10 9 13 13 2 3 2 9 1 9 0 2 9 1 9 7 9 1 9 2
24 9 1 10 11 2 1 9 1 9 2 13 16 10 9 13 1 13 10 0 9 1 10 9 2
14 9 0 3 11 7 11 13 9 1 13 1 10 11 2
21 15 13 2 3 2 16 10 9 0 1 11 7 10 9 15 13 1 9 1 9 2
33 1 10 9 2 10 11 13 9 0 1 10 9 1 10 11 1 10 0 9 1 10 11 2 10 9 0 0 2 13 1 12 2 2
2 0 9
42 13 12 10 9 1 10 9 15 13 10 9 1 9 1 10 9 2 10 9 3 13 4 13 2 10 9 1 9 0 13 4 13 7 11 13 1 10 9 1 10 9 2
2 9 0
25 9 0 13 1 13 9 10 9 2 13 1 10 9 2 13 16 10 9 1 10 9 13 10 9 2
20 10 9 13 1 10 9 1 0 9 13 11 2 11 2 11 2 11 7 11 2
15 1 0 9 2 13 11 2 11 2 11 2 11 7 11 2
15 1 10 9 2 13 11 2 11 2 11 2 11 7 11 2
26 10 11 13 13 1 10 2 11 2 7 1 10 9 2 11 2 2 7 13 10 9 1 10 9 11 2
27 10 9 13 9 1 10 9 2 0 9 1 9 2 0 9 1 9 2 0 9 1 9 0 2 1 15 2
2 10 9
4 9 1 10 9
3 1 10 9
13 10 11 13 10 9 0 2 7 13 10 9 1 13
3 1 10 9
10 11 7 11 13 3 7 13 11 7 11
4 9 1 10 9
3 1 10 9
14 10 11 3 15 13 1 10 9 1 10 9 1 10 9
29 11 2 9 0 1 10 11 2 13 16 10 9 3 13 10 9 2 7 16 10 9 1 9 3 13 13 1 9 2
20 15 13 16 10 9 0 1 10 9 3 13 13 15 12 5 13 1 10 11 2
14 10 9 2 3 2 13 13 10 9 0 1 10 9 2
8 11 7 11 13 13 1 10 11
13 0 9 1 9 1 10 12 0 9 1 10 9 2
28 11 7 11 13 1 10 11 2 1 10 11 2 1 9 3 13 1 10 9 0 10 9 11 7 10 9 11 2
19 10 0 9 1 13 13 11 2 15 13 10 3 9 11 1 12 7 12 2
4 11 13 0 2
20 11 2 1 12 9 7 9 12 1 10 9 2 13 10 0 9 1 10 9 2
24 2 13 9 13 1 10 9 2 3 2 2 16 3 13 13 0 1 13 11 2 2 13 11 2
3 13 1 13
43 11 2 16 10 9 15 13 1 10 9 1 13 10 10 9 1 10 9 13 3 1 10 11 2 13 13 16 2 3 3 13 1 10 9 2 13 9 0 2 3 7 3 2
22 16 13 10 9 3 10 9 1 15 13 2 13 13 3 16 10 10 9 13 13 0 2
7 13 0 13 3 10 15 2
7 13 3 1 11 10 9 11
22 10 12 9 1 10 9 1 10 9 1 9 13 9 1 9 12 9 1 10 0 9 2
7 13 13 3 12 12 9 2
19 10 11 13 1 10 11 2 9 0 1 11 2 7 13 13 1 10 9 2
5 9 0 13 10 11
23 10 11 1 10 11 13 3 16 1 9 2 9 12 2 10 11 2 11 2 13 9 12 2
14 10 9 13 1 12 5 2 0 1 10 11 1 9 2
28 10 9 15 13 10 9 2 11 2 9 3 2 3 13 13 2 16 10 9 13 13 1 10 11 1 9 12 2
7 9 1 11 13 13 9 12
31 13 13 1 10 0 9 12 2 1 10 9 1 10 9 2 1 10 9 2 10 9 2 11 2 2 13 1 10 9 11 2
27 9 1 10 9 1 10 11 2 15 13 13 10 0 9 1 9 1 12 2 11 13 10 9 1 10 9 2
32 3 1 9 2 1 10 9 1 10 9 2 13 15 10 9 1 10 9 11 2 1 10 0 9 1 10 0 9 2 7 11 2
15 10 9 13 10 9 1 10 9 15 13 0 9 1 9 2
13 9 1 10 9 13 13 1 10 9 1 9 2 2
13 2 9 1 9 1 9 0 1 10 12 0 9 0
13 11 15 13 1 9 2 1 10 9 1 10 11 2
42 10 9 11 2 12 1 10 9 1 10 9 0 1 10 9 2 13 13 15 1 10 9 0 1 10 0 9 1 13 10 9 1 2 10 9 2 15 13 1 10 9 2
21 2 3 13 16 13 9 2 13 13 15 13 1 10 10 9 7 9 2 2 13 2
30 11 2 12 2 13 16 13 10 2 9 2 15 3 13 9 1 10 9 2 3 15 13 1 10 9 2 1 9 13 2
25 2 13 9 7 2 3 13 10 9 1 9 1 10 9 2 13 13 10 9 2 2 13 10 9 2
3 9 1 11
19 2 3 13 16 15 13 13 10 9 2 7 13 15 15 13 1 15 2 2
15 11 2 9 0 1 10 11 2 3 1 10 2 11 2 2
17 11 7 10 9 15 15 13 13 1 10 9 1 10 9 1 3 2
24 15 13 1 10 9 1 3 12 9 7 13 1 13 1 10 9 11 1 10 9 1 10 9 2
20 1 9 1 10 9 2 15 13 10 9 16 11 13 10 9 9 15 3 13 2
8 15 13 1 13 9 1 9 2
18 1 10 9 2 10 9 13 1 9 13 1 12 9 2 1 9 0 2
11 1 10 9 3 13 9 13 1 12 9 2
5 15 13 9 0 2
18 10 9 0 13 1 9 0 13 2 9 11 2 1 9 1 12 9 2
11 10 9 0 13 0 1 10 0 9 11 2
5 9 13 9 1 12
49 10 11 2 11 2 13 4 1 13 1 10 9 10 9 1 9 1 10 9 1 10 12 9 0 13 1 10 9 1 12 9 1 10 9 12 1 10 11 2 1 10 11 2 9 0 1 11 2 2
27 10 9 13 3 10 9 1 9 1 10 11 13 10 9 1 13 1 10 9 2 1 12 1 9 1 12 2
24 3 2 3 3 2 1 10 9 0 2 10 11 13 1 10 9 1 10 9 16 3 13 9 2
21 13 0 10 9 1 10 11 2 11 2 2 11 2 11 2 7 11 2 11 2 2
16 1 10 9 0 2 11 7 11 13 13 3 9 1 10 9 2
25 10 11 13 3 1 11 2 1 10 9 2 1 10 9 1 10 11 2 9 2 2 10 9 0 2
23 10 11 1 11 2 11 2 13 9 2 1 10 9 2 1 10 11 2 1 10 9 11 2
17 1 11 2 10 9 13 13 9 1 9 2 9 1 9 7 9 2
28 1 11 2 13 3 10 9 1 10 9 1 10 11 2 9 2 1 10 9 1 9 1 10 9 1 10 9 2
22 1 9 0 2 9 1 10 11 7 1 10 11 13 9 1 9 7 1 9 1 9 2
27 10 9 13 4 13 1 10 9 11 2 15 13 10 9 1 9 1 9 15 3 13 13 3 10 9 0 2
11 1 9 2 12 9 3 13 13 10 9 2
29 2 13 13 12 9 1 10 12 9 7 13 10 9 2 2 13 10 9 1 9 11 2 12 2 12 1 10 9 2
29 3 2 3 10 0 9 7 9 2 13 2 10 9 1 15 13 2 0 10 9 1 15 1 13 13 1 10 9 2
48 3 2 10 9 3 13 13 13 1 10 9 9 15 3 13 16 15 13 10 9 1 10 9 2 13 7 13 9 7 9 0 2 13 9 0 2 13 10 9 0 2 13 9 7 10 10 9 2
6 9 13 13 9 7 9
27 1 13 10 9 1 10 9 1 11 1 10 9 1 10 11 2 12 9 0 13 3 10 9 1 10 11 2
20 11 7 11 2 9 7 9 2 13 13 1 10 0 9 1 9 15 13 13 2
33 3 1 15 10 9 2 10 11 2 15 13 9 1 10 11 7 9 1 11 2 15 13 10 9 1 10 9 7 10 9 1 9 2
6 9 13 13 13 1 11
37 2 15 13 13 2 2 13 10 9 11 2 12 2 1 10 9 1 10 11 1 11 2 3 13 3 10 9 2 11 2 1 10 9 11 2 12 2
8 11 3 13 16 3 13 13 2
3 3 13 2
18 11 13 16 10 9 1 10 9 13 2 13 3 2 10 9 1 11 2
34 1 12 9 13 2 7 10 0 1 9 2 10 9 13 3 2 1 10 0 9 2 16 11 13 13 15 1 10 9 0 1 10 9 2
20 2 11 2 2 15 10 11 13 3 1 10 11 2 13 10 0 9 1 11 2
20 10 10 9 13 2 1 12 2 10 9 1 9 1 10 9 2 2 11 2 2
7 11 1 15 13 1 10 11
21 10 9 0 2 12 2 15 13 1 11 2 1 10 9 1 10 11 1 12 9 2
18 1 12 2 11 13 10 11 2 10 0 9 1 10 9 1 10 9 2
6 9 13 1 13 10 9
21 11 2 12 2 1 10 11 2 1 10 0 9 2 13 9 1 9 2 1 11 2
9 11 15 13 1 10 9 1 9 2
15 3 12 5 1 10 9 1 10 9 13 13 1 9 0 2
38 2 10 9 1 10 9 13 16 2 3 1 12 9 2 10 9 13 13 12 9 2 10 9 7 10 9 2 2 13 10 9 11 2 12 2 11 2 2
28 7 10 11 15 13 16 9 1 10 11 2 3 9 2 13 3 2 15 13 10 9 1 10 9 7 13 13 2
2 6 2
5 9 1 10 9 2
8 7 13 15 15 3 3 13 2
8 10 11 1 10 2 9 2 2
8 10 11 10 9 13 10 9 2
4 15 13 13 2
8 13 13 3 9 1 10 9 2
2 6 2
31 1 10 9 1 10 9 11 2 10 9 13 9 1 1 12 5 1 10 9 2 13 9 0 7 9 1 10 9 1 9 2
27 10 9 11 13 13 1 10 9 2 1 10 9 2 10 9 1 10 0 9 13 1 9 0 1 10 11 2
9 10 11 13 3 13 9 1 9 2
28 10 9 11 3 13 9 2 1 10 2 1 10 11 1 11 2 10 11 2 10 11 2 10 11 7 10 11 2
37 9 1 10 11 2 1 10 0 12 9 11 13 10 9 1 11 2 10 9 2 1 10 2 11 2 2 10 9 1 10 9 1 9 2 11 2 2
13 13 1 10 9 2 11 13 1 13 1 10 11 2
24 2 13 0 2 15 13 12 9 0 16 15 13 2 2 13 1 11 1 13 10 9 1 9 2
22 13 10 9 2 10 9 1 10 9 2 7 13 1 10 11 13 10 9 1 10 9 2
9 11 13 10 9 7 15 13 2 11
12 9 13 10 9 1 9 2 1 10 9 0 2
11 10 9 11 13 10 11 1 9 1 9 2
4 7 13 3 2
24 1 10 9 7 10 9 13 1 12 9 7 0 2 13 10 9 1 9 12 9 1 10 9 2
40 1 10 9 1 10 9 1 15 13 10 9 1 10 9 1 10 11 2 13 1 12 9 1 9 2 13 1 9 2 7 13 12 1 10 9 1 9 7 11 2
14 15 13 13 10 9 7 10 9 13 1 10 10 9 2
7 10 9 13 15 13 13 2
13 1 13 10 9 1 10 9 2 11 3 13 9 2
24 1 11 2 10 9 1 13 13 0 1 9 1 9 2 9 2 9 2 9 1 9 7 9 2
29 1 10 9 1 10 9 2 11 13 13 1 10 9 0 7 1 10 9 15 13 1 10 9 1 13 10 9 0 2
29 10 9 1 10 9 1 10 11 13 13 9 1 10 12 9 1 10 9 1 10 9 1 10 9 11 7 10 0 2
29 1 10 11 2 10 9 13 1 10 9 1 9 7 16 15 13 10 9 2 1 10 0 9 1 10 9 1 9 2
11 15 3 13 13 10 9 11 2 11 2 2
30 1 10 9 1 10 9 0 1 10 9 2 13 15 10 9 1 9 1 10 9 2 9 3 13 1 10 9 1 9 2
40 7 10 9 1 10 9 0 2 9 13 1 9 1 9 0 15 13 10 9 1 10 9 2 7 10 9 1 10 9 13 13 1 9 1 10 9 1 10 9 2
18 11 13 16 3 13 10 9 1 9 7 16 10 9 13 13 1 9 2
26 3 2 13 3 13 2 16 9 13 15 2 2 7 16 2 1 3 10 9 13 13 1 10 9 2 2
30 1 15 15 10 9 13 2 10 9 0 3 13 13 1 13 9 1 10 9 1 9 1 10 9 0 15 13 10 9 2
23 2 3 13 13 9 15 13 10 9 1 10 9 2 2 13 11 2 1 13 1 10 9 2
34 13 1 10 9 1 10 11 1 10 9 2 10 9 13 13 0 1 3 13 2 1 3 2 9 0 0 1 10 9 1 10 9 0 2
21 15 13 16 10 11 1 11 13 13 16 3 13 9 0 1 10 9 1 10 9 2
1 9
38 1 15 15 13 13 1 10 0 9 0 2 11 13 3 13 9 1 10 13 2 9 0 1 9 2 1 10 9 0 9 15 13 13 9 1 10 9 2
31 10 9 13 15 1 13 16 13 13 1 9 1 9 1 10 9 11 1 10 9 1 10 0 9 1 9 1 10 9 0 2
11 10 9 2 1 10 11 2 13 3 0 2
18 10 9 13 12 9 2 10 11 2 12 2 10 11 13 0 1 12 2
12 10 9 1 9 1 10 12 9 13 10 9 2
6 10 9 11 13 0 2
18 13 13 1 10 9 13 1 11 1 11 2 0 9 1 10 11 9 2
15 3 10 11 2 13 10 9 1 10 9 2 13 1 3 2
20 15 13 16 10 9 1 10 9 13 10 9 15 13 10 11 1 10 9 0 2
22 1 15 2 3 1 12 2 13 1 13 10 9 0 1 10 9 2 13 10 9 0 2
22 3 15 13 10 0 9 0 0 1 10 9 1 10 11 2 9 15 13 10 11 2 2
31 3 2 3 13 13 9 3 1 9 12 9 1 10 0 12 9 1 10 11 7 15 9 12 9 1 10 11 2 13 11 2
39 1 10 0 12 9 2 3 1 10 11 2 10 11 13 9 12 9 1 10 9 1 0 9 7 9 1 0 9 2 13 11 1 9 1 10 9 0 11 2
8 2 13 9 1 10 9 12 2
48 12 1 10 9 1 15 13 10 9 1 10 9 0 2 1 12 2 10 9 0 13 1 10 9 0 13 12 5 1 10 9 1 9 13 1 10 11 7 13 10 0 1 12 5 1 10 9 2
34 10 9 13 1 9 1 10 9 0 2 1 15 10 9 13 13 10 0 9 0 13 2 7 10 9 13 13 1 13 15 1 10 9 2
26 1 10 9 0 1 0 9 1 9 2 11 13 2 3 2 13 10 9 1 9 1 10 9 1 9 2
33 15 13 1 10 9 2 15 13 10 9 1 10 9 1 9 0 0 2 16 10 9 13 13 3 10 9 1 9 1 10 10 9 2
5 9 13 10 0 9
4 9 13 9 0
6 10 9 13 1 9 2
31 10 9 13 1 10 9 13 1 10 9 1 12 5 1 10 9 1 10 9 13 1 12 5 1 10 9 1 10 0 9 2
38 11 2 9 1 10 11 2 13 10 9 13 1 9 0 2 7 16 10 9 1 9 13 10 9 0 1 10 9 0 1 9 1 10 9 1 12 9 2
23 10 9 1 9 2 1 10 9 0 0 2 13 10 9 1 10 9 9 2 9 0 2 2
17 3 13 10 11 16 3 13 1 15 15 3 13 2 10 9 2 2
21 10 9 1 10 9 9 2 9 0 2 13 9 1 10 9 7 9 1 10 9 2
23 10 11 13 10 9 13 7 13 1 10 0 7 3 0 9 1 9 1 9 1 9 0 2
30 2 10 9 3 13 9 1 10 10 9 7 13 13 3 3 1 10 11 2 2 13 11 2 12 2 9 1 10 11 2
14 10 9 13 4 13 1 10 9 1 10 2 11 2 2
16 10 9 2 16 13 13 2 13 13 3 13 3 1 10 9 2
17 1 10 9 1 10 9 2 10 9 1 10 9 13 10 9 0 2
12 1 10 9 2 13 10 9 1 10 9 0 2
31 10 9 13 10 9 1 9 1 10 9 1 10 9 1 10 9 2 15 3 13 10 9 1 9 1 10 9 1 10 11 2
24 10 9 1 9 1 10 11 13 3 16 10 9 3 13 15 13 1 16 13 13 1 10 9 2
12 11 13 10 0 9 1 10 2 1 12 9 2
8 11 13 1 13 2 1 12 2
9 11 13 1 10 9 2 1 12 2
24 3 2 11 3 13 10 0 9 1 9 2 12 2 2 1 12 1 11 7 3 12 1 11 2
9 10 9 13 0 2 7 3 13 2
16 13 16 15 13 3 1 9 7 1 9 16 10 9 13 9 2
28 3 3 15 13 10 9 1 10 9 2 13 10 9 2 7 10 9 2 15 13 10 9 1 16 3 13 9 2
15 15 13 10 9 2 16 13 1 13 16 10 9 13 13 2
10 9 13 1 12 11 12 9 1 12 11
9 9 1 10 9 2 13 1 0 2
2 9 0
14 1 13 1 10 11 2 13 10 9 0 1 9 0 2
12 3 13 1 10 9 0 7 10 9 1 9 2
21 3 1 10 9 0 1 10 9 0 2 13 0 13 10 9 1 13 13 1 10 9
9 13 10 9 1 13 10 9 0 2
26 10 9 13 10 9 1 10 9 7 10 9 2 3 0 2 1 10 9 1 10 9 7 1 10 9 2
33 1 10 9 2 16 10 9 1 10 9 1 10 0 13 13 1 12 9 2 15 1 10 9 7 1 10 9 13 4 13 3 3 2
11 13 3 15 15 13 1 10 9 1 9 2
20 3 2 13 10 9 1 10 9 0 1 12 9 7 3 13 13 10 9 13 2
9 9 1 10 9 1 9 3 13 3
34 10 9 1 10 9 2 11 2 13 16 10 9 1 9 1 10 9 1 9 1 9 2 0 1 10 9 1 10 9 2 13 3 13 2
29 1 10 9 1 11 1 10 11 2 11 2 10 9 1 9 13 3 1 10 0 9 1 9 2 7 13 0 3 2
28 11 13 16 10 9 3 13 1 9 10 9 1 10 9 13 15 13 7 13 1 10 9 1 13 10 9 11 2
13 2 3 3 15 13 16 10 9 13 13 7 3 2
5 13 1 9 2 2
35 10 9 2 3 2 3 13 1 10 9 1 10 2 9 1 9 2 1 9 0 2 7 13 13 1 10 12 9 15 13 10 9 1 11 2
20 7 10 9 2 3 2 13 10 15 3 1 10 9 1 10 9 1 10 9 2
51 12 9 1 10 9 1 11 2 1 10 9 9 3 1 10 9 13 10 0 9 2 11 13 10 2 0 1 10 9 0 7 0 1 10 9 7 9 2 7 1 10 2 0 7 0 9 1 10 9 2 2
7 9 13 9 2 13 2 2
15 10 9 7 9 11 3 13 9 1 10 0 1 10 9 2
16 1 15 2 10 9 13 2 9 13 2 13 1 9 0 2 2
14 10 9 13 13 3 3 1 10 9 1 10 9 0 2
19 10 9 1 10 11 13 16 10 9 13 12 5 1 10 0 9 1 9 2
20 10 9 13 10 9 1 10 9 0 13 1 10 11 2 1 9 1 10 11 2
23 10 9 1 9 15 13 3 9 1 9 7 1 9 13 9 1 12 5 1 10 9 0 2
5 13 1 10 9 2
3 13 15 2
5 9 13 10 9 2
5 3 1 10 9 2
13 10 9 3 13 13 1 13 9 15 13 10 9 2
19 1 10 11 2 9 0 2 3 15 13 11 1 12 9 10 9 2 3 2
7 0 9 13 9 2 13 9
12 9 1 10 11 13 16 10 9 13 0 9 3
35 10 9 2 9 2 13 3 0 1 13 9 3 16 15 3 13 2 1 9 1 10 0 9 1 10 9 1 10 11 2 2 11 2 2 2
11 10 9 13 4 13 3 1 9 1 9 2
20 15 13 9 13 3 0 1 10 9 2 9 3 10 9 13 1 10 9 2 2
12 10 9 3 13 10 9 1 13 1 10 9 2
26 1 13 10 0 9 0 2 11 13 10 9 1 10 9 11 2 15 13 13 1 10 9 1 10 9 2
22 10 9 0 2 1 10 0 9 2 13 10 9 1 10 11 7 13 13 1 10 9 2
8 9 1 9 1 15 7 11 2
16 1 10 9 2 13 10 9 0 2 1 15 12 5 1 9 2
33 11 2 1 9 1 10 9 2 3 13 16 2 1 9 2 3 15 13 13 3 2 7 1 9 10 9 13 0 1 10 9 2 2
16 3 15 13 16 1 9 10 2 9 2 1 9 13 4 13 2
4 9 2 3 2
12 7 2 1 9 2 10 9 13 10 9 3 2
9 1 9 2 13 15 10 10 9 2
5 9 13 9 1 9
6 9 7 9 13 1 13
21 10 11 13 1 13 10 9 1 9 1 9 1 13 3 15 13 13 10 0 9 2
29 2 13 13 10 9 2 10 9 11 2 1 10 11 2 1 13 10 9 1 10 10 9 1 9 2 2 13 11 2
53 3 15 2 7 3 2 3 1 10 0 9 1 9 2 2 10 9 11 13 0 9 1 13 10 9 1 10 11 2 12 9 1 9 2 9 1 12 5 13 2 10 9 1 9 2 9 2 1 9 2 9 2 2
12 1 10 9 2 10 0 9 1 10 9 0 2
26 3 15 2 3 10 9 1 13 9 2 2 10 11 13 10 9 1 10 9 1 10 11 15 15 13 2
18 15 1 10 9 1 10 9 1 10 9 13 3 9 10 9 1 9 2
23 3 2 13 12 9 15 13 1 2 2 2 10 9 1 11 13 13 10 9 1 12 9 2
8 10 11 3 13 13 10 9 2
26 10 9 2 13 1 10 9 11 2 12 2 13 9 1 10 9 1 10 9 13 2 1 0 10 9 2
16 10 11 13 12 9 1 10 9 0 13 10 9 1 10 9 2
22 1 13 1 9 2 10 9 1 9 13 13 3 16 13 10 9 1 9 2 13 11 2
6 10 9 13 9 0 2
15 1 11 2 1 10 9 2 10 9 13 3 0 7 0 2
16 15 13 16 3 13 9 1 10 9 1 10 9 1 10 9 2
5 13 10 9 1 9
21 9 13 0 9 1 13 9 1 9 1 10 9 1 0 9 2 13 3 10 0 9
15 1 10 9 1 10 9 1 9 3 13 13 3 10 9 2
19 13 10 9 13 10 9 7 13 10 9 1 9 1 10 9 9 1 9 2
29 10 11 13 1 10 11 12 9 1 9 9 1 13 2 15 13 13 10 9 0 1 10 9 1 10 9 7 9 2
5 9 1 11 13 13
26 10 11 1 10 11 13 3 9 1 10 9 1 10 9 0 1 11 1 10 9 1 13 0 9 0 2
39 1 11 2 10 11 2 11 2 10 9 0 1 10 11 2 13 10 9 0 1 10 9 1 10 9 1 3 13 16 10 9 1 11 13 10 9 1 9 2
20 10 9 13 16 13 3 12 9 1 11 1 10 9 0 1 13 9 1 9 2
13 2 10 9 15 13 4 13 13 2 2 13 9 2
21 3 10 12 9 13 1 10 11 13 12 9 1 9 0 2 0 2 0 7 0 2
14 10 9 0 13 9 12 12 2 0 1 9 12 12 2
20 10 9 0 13 10 0 9 1 10 11 2 9 12 12 2 9 12 12 2 2
11 13 13 1 10 11 7 13 1 10 11 2
15 11 2 10 9 3 13 10 9 1 10 9 1 10 9 2
23 11 2 3 13 13 13 3 1 10 9 1 10 9 16 3 15 13 13 9 1 10 9 2
13 9 13 13 12 5 3 2 1 10 9 1 11 2
43 10 9 0 1 10 9 0 13 13 1 12 5 16 10 11 13 10 9 1 10 9 0 1 10 9 1 10 9 7 10 9 1 10 9 1 9 1 10 11 2 11 2 2
15 3 10 9 13 1 10 9 1 10 9 15 13 10 9 2
29 10 9 1 9 1 10 9 1 10 9 1 9 1 10 9 13 13 1 13 1 9 12 9 10 11 2 11 2 2
36 10 9 13 16 13 1 12 5 1 12 5 10 0 1 10 9 1 10 9 15 13 13 9 1 10 11 1 13 10 9 1 9 1 10 11 2
21 10 9 13 13 3 9 12 9 1 10 11 2 3 1 9 15 13 1 10 9 2
6 10 9 1 10 9 11
23 10 9 13 2 1 10 9 2 10 9 3 0 1 10 0 9 1 10 9 1 10 9 2
64 13 3 10 9 1 10 9 1 10 9 13 1 13 1 9 1 10 9 2 1 10 0 9 0 1 10 9 0 0 10 9 15 13 9 1 9 7 9 2 9 1 11 1 11 2 13 1 10 10 9 0 2 9 2 9 0 2 9 7 9 1 10 0 2
12 10 9 0 0 13 3 1 9 0 3 11 2
2 9 13
32 11 2 9 1 10 11 2 13 16 10 9 13 3 3 10 9 2 11 2 2 15 13 1 13 7 13 9 1 10 9 2 2
15 13 16 15 13 1 12 9 2 3 10 9 13 1 11 2
25 10 9 13 13 10 0 9 1 10 9 1 10 9 7 2 1 10 12 9 2 3 13 13 9 2
6 2 13 3 13 2 2
23 3 2 10 9 13 13 13 10 9 0 1 10 9 2 3 10 9 0 13 1 12 9 2
11 13 1 10 9 1 10 9 2 11 13 2
9 2 13 0 2 7 13 15 2 2
42 1 13 13 1 9 16 2 1 10 0 7 0 7 10 0 2 2 13 1 10 0 7 0 2 11 13 16 10 9 0 2 1 10 0 9 2 13 13 1 10 9 2
26 11 13 1 10 11 1 9 1 10 9 2 3 13 3 1 10 11 2 3 13 1 9 1 10 9 2
4 13 0 1 11
25 2 11 2 2 1 12 2 13 10 9 2 1 10 9 13 2 10 9 13 10 9 3 16 0 2
10 3 3 1 15 3 2 11 2 13 2
26 10 9 1 11 1 10 9 1 10 9 0 0 13 10 9 3 0 2 10 9 1 9 1 13 0 2
17 3 1 15 10 11 1 2 11 2 13 1 10 9 1 10 9 2
23 10 9 1 11 13 3 2 1 11 15 13 1 13 9 1 10 9 1 10 9 1 9 2
22 7 1 10 9 13 10 9 0 15 13 10 9 0 1 10 0 9 1 10 9 12 2
34 1 11 7 11 2 3 13 1 9 0 0 10 9 11 2 0 2 11 2 2 11 2 0 2 11 2 7 11 2 0 2 11 2 2
25 3 2 10 9 1 10 11 1 10 11 13 10 9 1 10 9 1 10 0 9 1 10 0 9 2
29 10 9 13 12 9 1 11 2 0 2 9 2 7 12 1 11 2 0 2 11 2 1 10 0 9 2 11 2 2
9 10 9 13 13 1 10 10 9 2
8 3 13 13 12 9 1 11 2
2 13 3
13 10 11 13 9 0 16 15 13 1 10 0 9 2
21 10 9 13 12 5 1 9 12 9 7 10 9 2 12 5 2 1 9 12 9 2
27 10 11 3 13 0 9 2 13 9 1 9 1 15 13 13 10 9 1 10 0 9 1 9 1 10 11 2
2 10 9
32 10 9 11 2 1 10 9 1 11 2 13 16 2 1 9 2 13 13 10 9 2 3 1 9 1 10 11 7 1 10 11 2
20 13 16 2 1 10 0 9 1 9 2 10 9 0 1 9 13 1 12 5 2
17 1 13 10 9 2 10 9 13 10 9 1 9 1 3 12 9 2
10 13 13 10 9 1 12 9 7 9 2
26 1 11 2 13 12 9 0 2 11 7 11 2 7 12 9 2 11 7 11 2 10 1 10 11 2 2
23 10 9 13 13 1 11 3 2 10 9 1 9 1 10 9 2 2 3 10 0 9 13 2
11 11 13 3 10 9 1 10 9 1 11 2
6 2 3 13 15 13 2
17 13 0 2 2 13 15 15 11 13 1 1 10 9 1 10 9 2
5 13 3 13 10 9
69 10 9 0 1 12 1 9 1 12 1 10 11 2 11 2 13 16 2 10 9 1 9 1 9 1 10 9 9 2 9 1 9 7 9 2 1 10 9 2 13 13 1 13 1 9 0 2 3 13 7 13 1 10 9 7 9 1 9 0 1 9 2 1 9 1 10 9 2 2
31 10 9 13 3 16 12 5 1 10 9 13 16 4 13 7 13 13 9 1 9 7 9 1 10 10 9 0 1 10 9 2
13 10 9 1 9 1 9 7 9 13 9 3 0 2
3 9 7 9
68 10 11 1 10 11 13 16 2 3 10 9 13 9 1 9 1 9 2 9 7 1 9 13 1 2 9 2 7 2 9 1 9 2 7 13 1 10 9 13 1 3 12 9 2 13 0 10 9 1 10 13 9 1 10 9 1 9 1 10 11 2 11 2 9 11 12 2 2
3 11 2 9
72 10 9 1 10 11 13 4 13 1 9 2 16 2 16 1 9 1 12 11 2 1 0 9 3 1 10 9 2 13 1 9 1 9 7 9 1 10 9 7 1 15 13 2 1 9 1 10 9 2 7 16 1 9 1 12 11 3 13 4 13 1 9 2 11 2 9 0 11 9 12 2 2
23 1 15 2 15 13 10 9 1 10 9 13 10 9 1 10 9 0 2 3 11 7 11 2
3 1 10 0
34 3 13 1 10 0 1 10 11 2 15 13 13 1 9 1 11 2 10 9 0 13 10 9 1 10 9 1 10 9 1 10 0 9 2
8 2 11 2 9 1 10 11 2
21 2 15 13 16 13 1 12 9 7 13 1 15 10 2 1 10 9 13 13 2 2
9 2 11 2 9 1 10 9 0 2
13 2 9 2 3 13 10 9 1 10 9 1 9 2
11 10 9 1 10 9 1 3 13 13 3 2
23 1 11 2 9 7 9 1 10 11 1 9 2 1 10 9 2 15 13 7 13 9 2 2
24 3 2 10 0 9 1 9 13 13 1 9 15 13 10 9 15 10 9 13 1 15 15 13 2
39 1 13 1 10 9 2 11 13 10 9 1 9 0 2 9 0 2 15 13 7 13 1 10 9 0 1 10 9 1 11 2 9 11 2 11 7 9 2 2
9 13 3 10 9 3 10 9 13 2
4 9 1 10 11
17 9 11 13 9 2 1 10 11 2 2 16 9 3 13 9 2 2
14 15 3 13 2 7 13 0 13 10 9 1 10 11 2
16 3 13 10 9 13 15 3 3 7 3 3 10 11 13 13 2
17 13 0 10 9 0 1 10 9 2 1 9 0 7 1 9 3 2
5 9 1 10 9 0
14 3 1 15 13 2 1 16 13 0 13 1 10 9 2
18 3 2 10 9 13 0 2 11 13 13 1 10 11 0 7 10 11 2
19 10 9 13 12 9 1 9 2 9 12 12 2 7 9 12 12 1 9 2
18 13 15 1 12 2 13 10 9 1 10 9 7 15 13 9 12 12 2
11 2 11 2 3 13 13 1 10 9 12 2
16 11 3 13 10 9 0 1 12 9 2 11 2 11 7 11 2
13 1 10 11 2 10 9 13 1 10 11 1 11 2
18 10 11 2 1 11 2 9 1 10 11 2 3 13 9 1 10 9 2
32 1 10 11 2 10 9 1 10 11 2 11 2 3 13 13 10 9 1 11 2 7 15 3 13 16 13 3 10 2 11 2 2
14 10 9 1 9 13 10 9 3 0 2 1 10 9 2
11 10 9 2 15 13 16 13 1 12 9 2
24 1 10 9 1 9 2 12 5 1 10 9 1 10 9 1 9 13 13 13 1 9 7 9 2
33 1 10 9 1 9 1 10 9 0 0 2 10 0 3 13 1 12 5 2 1 12 5 1 10 11 2 9 15 3 13 10 9 2
6 9 1 11 13 12 9
33 12 9 13 1 10 9 13 1 10 9 1 3 1 10 9 12 1 10 9 11 2 15 13 11 1 11 2 1 10 9 1 11 2
8 12 9 7 10 11 15 13 2
6 15 13 1 9 0 2
16 10 9 1 10 9 7 10 9 1 10 11 13 1 10 9 2
13 10 9 3 3 13 15 13 10 9 1 10 9 2
6 11 13 9 1 13 9
19 9 1 10 11 3 13 16 10 9 13 13 16 2 13 9 13 7 13 2
36 10 9 1 11 1 10 11 2 11 2 13 16 10 11 13 13 9 1 10 9 2 3 3 2 1 9 12 2 9 1 15 13 10 9 0 2
21 3 2 1 10 9 0 2 1 9 1 10 11 2 10 9 13 13 1 9 12 2
25 1 11 2 10 11 13 13 9 3 10 9 13 1 10 9 13 2 2 3 13 1 10 9 2 2
28 10 9 2 3 2 13 3 9 1 10 9 0 2 15 15 10 3 13 2 3 13 2 16 10 9 7 9 2
29 1 15 2 13 10 2 9 2 1 10 9 7 3 1 10 9 1 10 9 0 2 13 0 13 9 0 16 0 2
21 10 2 9 2 3 13 1 10 9 2 13 15 2 3 2 10 9 2 10 9 2
13 7 2 1 10 9 2 13 9 0 1 10 9 2
78 10 9 1 10 9 2 1 10 9 13 1 10 9 0 7 0 2 10 15 11 3 13 2 1 9 1 10 9 12 2 3 13 16 10 9 0 15 13 1 10 9 1 10 9 1 13 1 10 9 0 1 10 9 0 7 1 15 2 13 15 2 13 15 1 9 0 1 10 9 2 1 15 15 13 10 9 0 2
34 1 10 9 2 10 11 3 13 9 1 13 10 9 1 10 9 1 10 11 3 13 13 3 9 3 0 2 11 2 11 7 11 2 2
28 2 1 10 0 9 2 15 13 10 9 2 7 1 13 9 7 1 13 10 9 1 10 11 2 2 13 11 2
26 2 10 9 1 10 9 2 3 2 13 13 3 1 10 9 2 3 13 10 11 2 2 13 10 9 2
8 2 13 13 1 10 9 2 2
31 10 9 1 9 2 1 13 13 3 2 13 1 4 13 1 10 9 1 10 9 0 2 15 3 13 10 9 0 0 0 2
54 1 3 12 9 2 10 11 13 15 1 10 9 1 9 0 0 1 10 9 1 9 0 7 1 10 9 0 2 15 13 13 3 3 1 10 9 0 1 10 9 0 1 10 9 0 0 2 3 1 10 9 1 11 2
7 11 13 11 3 1 10 9
19 10 0 9 1 10 11 1 9 1 10 9 12 13 3 1 10 12 9 2
27 10 11 15 13 1 0 9 1 10 9 0 2 13 13 10 9 1 10 9 1 10 11 2 1 10 11 2
15 10 9 13 10 9 0 1 10 9 1 10 9 1 10 11
30 10 9 2 11 2 13 1 9 1 10 9 1 10 9 1 9 2 1 9 1 10 0 9 1 9 13 1 10 9 11
14 1 10 9 2 13 10 9 1 10 9 1 10 9 2
12 7 2 1 10 9 12 2 10 9 13 9 2
8 11 13 13 10 9 1 9 2
14 10 9 13 10 9 2 15 10 9 13 1 10 9 2
6 12 9 13 9 1 9
34 10 9 1 9 1 10 11 13 13 13 1 10 9 1 12 9 2 11 2 11 2 0 1 10 11 1 10 11 2 2 11 7 11 2
32 10 12 0 13 13 1 10 9 1 9 2 3 13 3 9 1 10 9 7 3 9 1 10 0 9 1 9 1 9 2 10 11
13 7 13 3 1 9 7 9 1 13 1 10 9 2
1 9
17 1 15 3 13 3 0 1 10 9 2 10 9 13 1 10 9 2
27 10 9 13 1 10 9 2 13 1 10 12 9 2 3 13 10 0 1 10 9 2 7 15 13 13 3 2
10 10 11 13 13 1 9 1 9 0 2
11 10 9 1 15 11 13 13 1 12 9 2
14 10 9 1 15 13 13 0 7 10 9 13 3 13 2
17 10 9 13 1 10 9 1 11 2 10 1 10 0 9 1 11 2
17 1 10 9 2 10 9 13 13 1 9 1 9 1 9 1 9 2
13 15 13 10 9 15 13 2 3 3 13 1 9 2
38 7 11 2 13 15 1 10 9 0 7 10 9 2 13 10 9 0 1 10 10 9 2 15 3 1 10 9 13 10 9 1 9 7 9 2 1 9 2
42 0 2 0 2 1 10 9 3 2 2 1 10 9 1 10 9 1 9 0 2 16 13 10 12 9 2 2 3 13 10 9 0 1 13 1 11 2 10 9 1 9 2
15 7 0 2 7 3 3 0 13 10 2 11 2 1 11 2
6 13 10 9 3 0 2
22 13 3 1 13 10 0 1 11 2 7 10 9 1 10 9 0 3 13 3 1 13 2
23 9 3 13 1 10 9 11 2 13 10 9 1 12 9 2 0 7 1 9 1 10 9 2
14 7 13 3 1 10 9 2 9 7 9 1 10 9 2
16 13 10 9 0 2 1 10 9 0 1 10 9 0 1 9 2
7 9 1 9 0 13 9 13
14 10 9 13 3 1 10 9 0 1 10 9 1 9 2
20 10 9 1 9 0 1 10 11 13 12 9 0 1 10 9 1 10 0 9 2
31 1 12 2 10 9 1 10 9 11 1 10 11 13 10 9 13 1 11 2 9 15 13 1 10 9 0 7 1 10 11 2
13 3 1 11 15 15 13 0 11 13 10 0 11 2
20 13 9 7 9 2 15 13 3 1 10 9 0 1 10 9 0 2 12 2 2
43 3 1 10 9 1 9 1 12 2 13 10 9 2 10 9 2 13 9 0 0 1 15 1 9 0 2 13 10 9 0 7 10 9 0 7 13 1 10 9 9 1 9 2
12 10 9 13 13 1 10 9 1 10 9 13 2
3 13 9 2
27 10 9 1 10 11 13 13 1 10 9 0 3 10 9 0 2 1 9 13 1 10 9 2 13 10 9 2
1 13
8 9 1 9 15 13 1 10 9
17 1 9 1 9 12 2 9 13 9 0 2 9 1 9 7 10 9
17 10 9 1 9 3 13 12 5 1 10 9 15 13 1 10 11 2
17 10 9 2 3 2 13 10 0 9 1 10 9 7 13 10 9 2
12 13 9 0 2 9 0 1 9 7 10 9 2
17 13 9 1 9 12 2 9 12 12 2 1 9 2 1 9 0 2
18 13 9 3 0 2 3 10 9 2 1 9 12 2 9 12 2 3 2
13 13 15 2 9 3 2 13 1 10 9 13 2 2
24 11 2 12 2 2 1 12 9 1 11 2 10 9 13 12 9 2 9 1 9 7 12 9 2
35 10 9 2 1 9 0 2 13 9 2 13 1 9 12 2 9 12 12 2 2 12 9 2 1 9 12 2 9 12 12 2 2 12 9 2
21 10 9 1 9 2 1 9 2 9 2 9 7 9 0 2 13 12 5 3 0 2
15 1 10 9 2 10 9 13 1 9 12 2 9 12 2 2
40 1 10 9 3 0 2 11 13 10 9 1 10 15 13 3 10 10 9 2 9 0 13 1 10 9 1 10 9 0 7 13 1 10 9 13 1 10 9 0 2
38 10 9 1 10 0 9 13 10 9 15 10 9 13 1 11 1 10 9 12 2 13 1 9 1 9 2 1 9 13 1 9 1 9 2 3 13 13 2
21 10 9 1 11 15 13 2 3 2 1 10 9 1 10 9 0 11 1 10 9 2
18 15 13 12 9 1 10 9 1 10 11 2 1 10 9 1 10 9 2
15 13 10 3 0 9 3 13 1 10 9 0 1 10 9 2
9 2 11 13 0 9 1 10 9 2
28 13 10 9 1 15 13 9 1 10 9 2 2 13 11 2 15 10 12 1 10 0 9 15 10 11 3 13 2
18 2 1 10 9 3 11 2 10 9 13 3 0 1 10 10 9 2 2
27 11 2 12 2 9 1 10 0 9 2 13 3 1 10 9 7 13 1 4 13 1 10 9 1 10 9 2
14 11 2 12 2 9 1 9 2 13 13 1 10 9 2
38 10 9 11 2 12 2 13 16 13 1 10 9 1 9 1 10 9 2 1 10 0 9 2 7 13 10 9 13 1 10 9 1 10 9 1 10 9 2
23 1 10 9 1 10 9 2 10 9 13 1 12 9 1 12 9 0 2 1 10 10 9 2
25 2 13 10 9 0 1 0 15 13 10 9 1 10 9 1 9 7 1 10 9 2 2 13 11 2
9 11 13 16 10 9 13 13 3 2
19 1 10 9 11 2 9 1 10 11 13 9 13 1 10 9 7 13 9 2
21 1 10 0 12 9 1 10 9 13 13 1 10 11 12 9 9 1 12 1 9 2
13 10 9 13 10 15 13 1 9 1 10 9 13 2
31 10 9 1 10 11 2 11 2 13 16 10 9 1 9 7 9 1 10 9 13 10 9 1 10 9 1 9 13 7 13 2
22 3 1 9 3 1 9 2 10 9 13 3 12 12 9 2 1 10 11 1 10 9 2
31 13 10 9 1 10 9 2 13 1 10 9 1 10 9 7 13 12 9 3 1 10 9 1 11 2 9 1 10 11 2 2
54 1 13 10 0 9 1 10 11 1 13 13 2 1 12 2 1 10 9 0 1 9 1 9 0 1 10 9 1 9 0 2 10 11 2 13 1 12 2 3 13 3 2 16 3 3 13 10 9 1 9 7 1 9 2
11 9 0 13 12 5 1 10 0 9 1 11
36 10 9 1 10 9 0 1 10 9 1 11 1 10 0 9 1 9 13 1 12 5 1 9 0 2 1 9 1 10 11 1 9 1 10 11 2
32 1 15 13 1 10 9 13 12 5 2 13 10 9 1 9 2 12 5 2 2 9 2 12 5 2 7 9 2 12 5 2 2
8 1 12 13 9 1 12 5 2
23 1 10 0 9 1 10 9 13 10 9 1 9 2 12 5 2 7 9 2 12 5 2 2
33 3 10 0 9 2 1 10 9 0 2 13 1 10 9 2 2 12 2 2 9 0 2 12 5 2 7 9 2 2 12 5 2 2
15 10 9 9 2 3 2 13 13 10 0 9 1 10 9 2
15 3 10 11 13 13 10 9 0 7 13 10 9 1 9 2
17 10 11 3 13 9 1 10 9 7 10 9 1 12 9 1 9 2
22 10 9 2 15 13 1 10 9 1 10 9 2 13 9 7 9 1 13 9 3 0 2
17 13 10 9 1 10 0 9 2 10 9 3 13 1 10 0 9 2
22 10 9 13 10 9 7 13 10 9 1 12 1 12 9 1 16 10 9 13 9 0 2
27 7 13 2 1 10 9 10 1 10 9 1 10 9 2 16 1 13 9 10 9 13 0 2 3 9 13 2
17 13 10 9 1 10 9 2 11 13 10 9 1 15 13 15 9 2
27 7 1 10 0 9 2 10 9 0 13 9 1 9 2 9 7 3 10 9 1 13 9 1 10 0 9 2
9 7 15 13 10 9 1 9 13 2
18 7 13 10 9 13 10 10 9 13 1 10 9 1 9 1 10 9 2
4 9 1 10 11
16 10 11 1 11 13 9 0 1 9 12 9 1 10 0 9 2
10 15 13 1 12 5 1 10 9 0 2
4 9 1 10 11
27 10 9 0 1 10 11 1 10 0 9 13 1 9 12 9 2 1 10 9 1 12 5 1 10 9 0 2
21 13 9 3 1 10 0 9 1 11 1 10 9 10 0 9 0 1 11 7 11 2
19 1 10 11 2 11 13 9 12 1 9 1 0 13 9 7 9 1 11 2
13 1 10 9 2 10 11 13 10 9 1 10 11 2
22 16 10 9 13 12 1 12 1 10 0 9 3 13 3 16 10 0 9 1 10 9 2
12 3 16 10 11 13 1 0 9 7 0 9 2
37 3 16 10 0 13 1 9 3 13 1 11 2 15 13 13 3 3 2 1 10 9 1 11 1 10 0 7 10 9 1 11 1 10 9 1 11 2
16 3 2 1 10 0 9 1 10 12 0 9 0 11 7 11 2
27 10 9 2 1 10 9 1 11 2 3 13 3 1 10 9 2 1 11 1 10 0 7 11 1 10 9 2
31 7 13 9 1 11 13 10 9 1 9 1 10 9 1 11 7 13 1 9 3 1 10 9 2 16 10 9 13 10 9 2
39 1 10 9 2 3 10 9 13 9 1 9 1 10 9 0 2 10 9 1 0 9 13 9 2 9 2 9 7 9 0 1 13 16 10 9 15 13 3 2
4 9 13 13 2
13 13 13 10 9 3 10 9 0 1 10 10 9 2
11 9 1 10 9 3 13 15 1 10 9 2
9 7 13 13 10 9 1 10 9 2
20 1 10 9 11 2 10 2 11 2 13 10 9 1 10 11 2 12 9 2 2
9 13 9 1 9 0 2 3 9 2
12 13 10 9 1 9 1 11 7 2 11 2 2
12 1 9 1 9 1 9 7 1 10 9 12 2
25 13 1 9 0 7 13 2 10 12 9 13 9 1 13 3 10 9 1 10 9 0 1 10 11 2
10 13 9 1 9 1 15 12 1 12 2
6 9 2 9 12 12 2
37 13 15 10 9 1 11 2 12 9 1 9 1 11 2 12 1 10 12 9 13 1 10 9 2 9 1 9 2 2 9 0 1 10 9 1 9 2
12 1 11 2 10 9 7 15 0 11 13 0 2
30 1 10 9 1 9 2 10 0 9 1 12 9 13 13 1 10 9 7 10 9 11 13 1 13 10 9 1 10 9 2
25 13 16 10 9 1 9 13 12 1 10 0 9 2 13 15 2 1 10 9 1 10 9 1 11 2
12 13 2 3 2 10 2 9 2 1 10 9 2
13 11 3 13 13 1 10 9 1 16 15 13 9 2
11 13 15 2 1 9 0 2 1 10 9 2
8 10 9 13 3 0 2 0 2
21 10 11 1 11 13 2 1 10 9 13 2 10 9 9 1 9 11 1 9 12 2
32 1 10 9 1 11 2 10 11 13 1 9 12 2 16 13 1 10 9 1 10 9 2 13 10 9 1 9 1 9 12 2 2
5 3 13 9 0 2
11 10 11 2 1 3 0 2 13 9 0 2
17 10 9 1 11 3 13 10 0 1 13 1 9 10 9 1 9 2
8 10 9 11 13 10 9 0 2
27 11 3 13 1 9 0 7 11 13 10 9 1 10 9 1 9 1 9 0 2 3 15 1 10 9 11 2
21 3 10 9 13 10 9 13 1 10 9 1 9 2 10 0 9 1 9 1 12 2
22 11 2 9 1 11 2 13 1 10 9 3 7 3 3 13 3 4 13 1 10 9 2
36 10 11 2 10 11 7 10 11 13 9 0 15 13 13 10 9 13 1 9 0 1 9 7 13 10 9 0 1 13 13 7 13 1 10 9 2
36 3 2 10 11 13 10 9 0 1 9 1 13 9 1 10 9 2 13 10 0 9 1 9 7 10 11 13 10 0 9 1 10 9 1 11 2
2 11 12
18 10 11 1 11 13 3 9 12 9 2 3 1 9 13 1 10 11 2
32 1 10 9 2 9 12 9 13 13 1 10 9 1 9 1 10 9 7 1 10 9 1 10 12 9 1 9 13 1 10 9 2
2 11 12
9 11 13 1 12 9 10 10 11 2
22 10 9 1 11 2 11 2 13 16 12 1 10 9 13 13 10 9 13 1 10 9 2
19 1 15 2 10 9 0 13 13 1 10 0 9 10 9 1 10 9 11 2
6 9 1 10 9 13 9
24 9 1 10 9 1 10 11 2 13 1 10 9 1 10 9 2 13 1 13 9 1 10 9 0
21 10 9 2 9 7 9 13 1 10 9 0 1 10 9 3 13 3 12 9 0 2
13 15 13 1 13 10 9 1 10 9 1 10 9 2
22 10 12 9 1 10 0 13 3 13 1 10 9 0 2 15 13 9 0 1 10 9 2
22 13 1 10 9 0 2 11 2 10 9 1 9 13 15 13 10 13 9 1 10 9 2
7 15 13 1 10 9 0 2
28 2 3 1 15 7 15 3 10 9 13 13 10 9 1 10 9 7 3 3 13 13 3 2 2 13 10 9 2
15 7 13 16 15 13 1 10 9 10 9 0 1 9 13 2
7 6 2 13 1 10 9 2
11 6 2 9 1 10 9 0 1 10 11 2
4 13 3 15 2
20 1 9 1 9 2 3 2 15 15 13 1 9 13 13 10 9 1 10 9 2
3 6 11 2
9 11 13 9 0 1 10 11 7 11
24 10 11 13 3 3 10 9 13 1 10 11 7 11 1 10 9 12 1 9 7 12 1 9 2
27 10 11 2 9 1 9 1 9 1 9 1 1 12 9 2 13 12 5 1 11 7 12 5 1 10 11 2
27 10 9 13 9 1 9 1 12 9 0 1 11 7 12 9 0 1 10 11 2 1 9 1 10 9 0 2
22 10 9 1 10 11 13 1 11 1 10 9 1 3 2 1 10 9 13 1 10 9 2
12 13 13 1 10 9 1 9 2 9 7 9 2
22 11 13 16 13 13 9 1 10 2 9 0 2 1 10 9 1 2 13 2 10 9 2
10 2 7 13 13 9 1 9 0 2 2
16 9 1 10 9 1 9 1 9 0 2 9 0 2 9 7 9
17 9 0 7 0 1 9 2 3 1 10 15 13 9 1 9 7 9
45 10 9 1 13 13 13 0 2 13 15 15 9 1 2 13 2 12 5 2 3 2 13 15 10 10 9 0 2 13 1 12 5 2 7 3 15 13 1 10 9 0 10 9 0 2
26 1 10 0 9 1 10 9 1 12 5 2 10 9 13 1 12 5 2 1 10 9 1 12 5 3 2
22 3 2 10 9 1 9 12 9 2 13 1 10 0 9 1 10 9 1 9 12 9 2
13 1 10 0 9 2 1 9 12 9 7 3 3 2
5 13 10 9 3 2
26 10 9 1 10 9 0 3 13 10 9 2 3 13 1 13 9 1 16 10 9 13 7 13 10 9 2
40 10 9 13 1 10 9 1 9 1 10 9 11 2 11 2 1 10 9 11 2 11 2 2 9 0 15 13 9 0 1 10 9 2 10 9 11 2 11 2 2
15 12 9 3 2 12 9 0 13 13 10 9 1 10 11 2
36 10 9 1 10 9 13 13 3 1 10 9 11 2 1 10 9 11 2 9 2 7 1 9 1 10 11 11 7 11 2 9 15 13 10 9 2
23 10 9 1 10 9 7 10 9 1 10 0 9 1 10 9 1 11 13 13 9 12 12 2
12 13 13 3 10 0 0 1 10 9 1 9 2
15 10 9 1 10 9 0 13 15 13 10 9 1 10 9 2
30 3 2 1 15 13 1 10 9 0 1 10 9 0 2 11 7 10 9 1 10 9 13 10 9 1 13 10 9 0 2
16 13 13 12 9 1 10 9 7 1 10 12 9 13 1 11 2
21 10 9 13 3 10 10 9 7 9 1 10 11 1 10 11 3 9 1 9 0 2
24 10 9 2 1 10 12 0 9 2 13 9 1 9 0 1 10 9 11 13 13 15 1 9 2
31 13 1 10 9 2 1 10 9 2 13 0 2 0 7 0 2 13 10 9 13 1 10 9 1 10 9 0 1 10 9 2
14 1 10 9 2 10 10 9 13 13 13 1 10 9 2
2 9 13
28 0 9 1 10 11 1 10 9 12 2 10 0 9 11 7 10 0 9 11 13 13 3 1 9 1 9 0 2
19 13 1 10 9 1 10 11 7 13 1 10 10 9 15 13 13 10 9 2
19 12 9 11 13 1 11 16 13 13 10 9 11 2 9 1 10 9 11 2
23 11 13 16 3 13 9 1 13 9 7 13 1 11 16 15 13 1 10 9 1 10 9 2
15 1 15 2 10 9 13 13 10 9 15 13 10 12 9 2
16 2 3 10 9 0 2 3 13 1 10 9 1 10 11 2 2
1 9
24 1 11 2 10 9 1 10 11 3 3 13 13 2 1 15 13 16 10 9 13 9 7 9 2
7 13 16 10 9 2 13 2
8 15 10 0 9 16 3 13 2
9 2 3 15 3 0 13 10 0 2
12 1 13 1 13 2 13 13 10 9 10 9 2
12 13 10 9 7 15 13 10 9 1 10 0 2
3 2 9 2
11 2 3 13 10 9 2 1 3 13 13 2
5 1 10 9 1 9
10 0 9 2 10 11 3 13 10 11 2
17 3 2 13 10 0 15 15 13 9 1 13 1 10 9 1 12 2
10 16 3 13 10 9 0 2 10 11 2
9 15 13 10 12 9 1 10 11 2
6 7 3 13 10 9 2
7 2 10 11 13 0 2 2
10 7 10 9 13 15 13 1 10 11 2
9 15 13 3 12 9 1 10 9 2
8 13 12 1 10 9 1 10 11
2 6 2
11 0 9 2 10 11 13 10 9 1 9 2
5 9 1 10 9 2
8 1 10 9 0 1 9 12 2
3 0 2 2
13 1 15 13 1 10 9 2 1 15 13 10 9 2
5 0 13 9 12 2
4 7 13 3 2
11 3 10 9 13 10 9 7 8 13 3 2
7 3 15 13 13 10 11 2
12 13 9 12 1 15 13 10 9 1 10 9 2
5 10 11 3 13 2
6 16 13 15 15 13 2
10 13 16 10 0 15 13 1 10 9 2
40 10 9 13 10 0 9 1 10 9 1 11 2 1 10 2 9 2 15 13 10 9 1 10 9 1 10 9 2 15 13 9 2 13 10 9 0 1 10 9 2
32 10 9 1 11 13 1 10 9 1 10 9 1 10 9 15 2 13 16 13 15 1 10 9 2 13 13 10 0 9 1 9 2
8 2 13 1 10 9 1 9 2
6 13 10 9 1 9 2
26 13 1 9 7 9 2 2 13 12 1 10 9 1 10 9 2 10 9 2 1 10 9 2 9 2 2
8 13 10 0 9 1 9 3 2
52 10 9 1 2 11 2 13 13 1 10 9 1 2 13 2 1 10 2 11 2 2 10 1 10 9 3 0 1 10 9 0 7 1 0 9 1 10 9 15 13 10 9 1 12 1 10 3 0 1 10 9 2
3 9 13 9
33 10 9 1 9 0 1 10 11 2 11 2 13 3 1 10 11 1 10 11 16 10 9 3 13 9 12 9 1 10 9 1 9 2
8 13 13 13 10 9 12 9 2
9 10 9 3 13 13 12 12 9 2
30 10 9 0 13 13 1 9 0 2 11 2 11 2 2 1 10 9 1 9 1 9 7 1 10 9 1 10 9 0 2
27 10 9 1 0 9 7 10 9 1 9 2 1 9 0 2 13 9 2 9 7 9 2 2 13 10 9 2
9 11 13 1 13 7 15 13 1 9
11 9 3 13 1 10 9 2 7 13 1 9
31 10 9 11 2 10 9 11 7 10 9 11 13 3 1 10 9 1 10 9 11 2 1 11 2 1 10 11 2 11 2 2
20 1 10 9 2 9 15 13 1 10 9 0 1 15 1 11 7 11 13 9 2
14 16 3 13 10 9 2 10 9 13 15 1 10 9 2
31 1 10 10 9 2 10 9 13 16 10 9 13 0 2 2 7 3 13 13 15 3 2 16 13 13 9 1 10 9 2 2
11 13 3 13 0 16 10 9 13 9 0 2
35 1 10 9 1 10 11 2 11 2 12 2 10 9 0 13 13 1 13 10 9 7 9 1 9 1 9 1 9 2 9 0 7 9 0 2
12 1 10 9 2 10 11 13 9 1 10 9 2
17 10 9 13 9 0 1 10 11 7 13 10 9 13 1 10 9 2
13 10 9 13 0 2 1 9 2 7 1 10 9 2
4 11 13 9 3
20 9 13 10 9 0 1 10 9 1 13 2 15 15 13 1 10 0 9 7 9
9 11 13 3 13 1 10 9 0 2
13 7 10 9 13 13 16 10 9 3 13 0 9 2
21 10 9 13 10 0 9 1 9 0 7 15 13 10 9 7 10 9 1 10 9 2
27 7 16 1 10 9 0 1 10 9 10 9 7 10 9 13 10 9 1 15 15 13 1 9 3 3 0 2
41 13 10 9 1 10 11 2 9 13 12 9 3 1 10 9 11 2 12 2 9 1 12 1 10 3 0 9 0 1 10 9 2 10 11 2 13 1 12 9 2 2
2 9 0
32 12 9 0 7 12 9 15 13 1 10 0 9 1 9 1 10 11 1 13 9 1 10 9 0 1 10 12 9 1 10 11 2
3 9 1 9
28 10 9 0 13 16 10 9 3 0 1 9 1 10 11 13 2 9 2 9 2 9 2 9 2 9 7 9 2
30 1 11 2 11 2 13 1 10 9 0 7 9 1 9 0 2 1 9 2 13 2 0 1 10 9 1 10 9 2 2
11 3 13 1 10 11 11 2 9 1 11 2
21 11 13 9 10 9 0 2 1 10 9 2 1 9 0 7 1 9 15 13 9 2
30 10 9 1 10 9 13 1 13 1 10 9 1 9 1 10 9 1 10 9 2 11 2 15 13 1 9 1 10 11 2
42 13 1 10 9 1 10 9 1 9 2 11 2 7 10 9 1 10 9 1 10 9 2 11 2 11 2 2 7 1 10 9 2 11 2 11 2 7 11 2 11 2 2
11 11 13 9 1 10 9 1 9 7 9 2
11 11 13 13 1 13 3 10 9 13 9 2
3 9 1 11
6 9 13 1 9 12 12
8 9 1 10 9 11 2 11 2
6 9 2 9 12 12 2
16 12 5 1 9 1 10 11 2 11 2 9 0 1 10 11 2
9 9 1 10 9 2 9 12 12 2
3 1 10 9
20 10 11 2 13 1 11 2 13 13 10 9 0 1 9 1 9 1 10 9 2
18 3 13 1 10 11 2 10 9 15 13 3 3 0 1 10 10 9 2
20 1 10 9 2 10 9 13 1 9 1 9 1 9 1 9 2 1 12 2 2
26 1 10 9 2 10 9 2 11 2 13 13 1 9 1 10 10 9 1 12 9 7 15 13 1 11 2
10 7 11 13 11 7 15 13 15 13 2
3 13 10 9
24 10 11 2 9 11 2 13 1 10 9 0 7 15 13 1 13 1 13 1 11 1 12 9 2
4 9 1 10 9
20 9 11 2 1 10 11 2 13 16 10 9 13 9 1 10 9 1 10 9 2
21 10 9 0 1 9 1 9 13 10 9 10 9 3 0 16 13 13 1 12 9 2
3 13 9 2
10 13 16 3 13 10 0 9 1 13 2
5 13 16 13 3 2
15 15 13 10 0 9 2 7 13 16 13 13 10 0 9 2
3 13 15 2
14 13 13 10 9 2 13 7 15 13 12 5 1 15 2
11 13 13 12 1 10 0 9 1 10 9 2
5 15 13 10 9 2
12 7 3 15 15 13 3 2 9 1 9 2 2
2 6 2
11 13 10 9 1 13 3 1 15 13 3 2
11 7 10 9 15 13 13 1 15 13 0 2
13 15 13 1 10 9 3 0 2 3 0 1 11 2
10 15 3 13 13 16 3 3 15 13 2
11 15 15 13 1 10 9 7 13 1 13 2
13 13 1 13 3 7 13 13 10 9 0 1 15 2
25 3 15 13 1 10 9 3 15 15 15 13 2 15 3 13 16 13 10 10 9 0 3 1 3 2
5 13 10 9 3 2
13 15 13 13 15 13 3 2 13 13 1 10 9 2
28 13 16 13 13 3 7 13 1 10 9 16 15 3 13 13 13 3 2 16 13 10 10 10 9 3 1 3 2
13 3 10 9 13 0 1 10 9 0 1 10 11 2
11 3 1 11 2 13 9 3 11 7 11 2
11 3 15 13 9 2 13 9 1 13 0 2
11 11 15 13 13 2 15 13 3 13 15 2
9 11 2 13 2 2 15 13 11 2
6 2 15 13 13 2 2
45 2 3 13 1 10 11 1 9 2 13 10 9 0 1 10 9 2 16 1 15 3 13 9 1 9 7 15 13 13 0 9 2 9 2 9 7 9 1 9 1 9 1 9 2 2
37 2 13 1 10 9 10 9 0 7 10 9 1 9 2 7 13 15 1 10 9 1 10 9 1 10 9 2 15 13 16 13 4 13 1 9 2 2
35 3 2 1 10 9 15 13 10 9 12 2 11 13 10 12 9 2 13 1 10 9 2 1 13 1 10 12 12 9 1 9 1 10 9 2
9 9 3 2 13 13 10 9 11 2
44 1 10 9 1 9 1 11 7 11 2 9 3 2 10 9 13 10 9 1 16 3 13 0 1 13 9 1 10 9 1 11 2 13 1 10 9 3 1 13 13 1 10 9 2
12 2 10 9 1 10 11 13 10 9 13 2 2
12 1 10 9 0 1 10 9 1 9 2 11 2
16 13 0 7 13 1 10 9 1 10 11 1 12 9 1 9 2
27 7 13 10 9 1 10 10 9 1 10 9 2 13 3 1 9 13 1 10 9 1 10 9 7 10 9 2
27 3 1 10 11 2 11 13 15 1 10 9 15 13 1 9 1 10 9 1 9 1 10 11 7 10 11 2
18 13 13 1 9 1 12 2 10 9 3 1 10 9 1 10 12 9 2
18 13 1 10 9 2 11 2 2 9 1 10 11 2 13 1 10 9 2
7 10 9 13 13 1 9 2
34 2 13 15 1 10 9 15 13 1 9 1 9 7 13 2 1 10 9 1 10 9 2 13 15 13 10 9 2 2 13 11 1 11 2
38 2 15 3 13 13 9 1 10 9 0 2 2 13 10 9 1 10 11 2 15 13 0 10 11 13 10 9 1 11 1 10 9 15 3 13 10 11 2
27 10 9 1 10 11 2 11 2 2 9 1 10 9 1 10 9 2 13 10 10 9 0 1 10 9 0 2
16 1 10 11 2 3 12 12 9 13 3 10 9 1 10 9 2
8 9 1 9 13 16 13 13 9
30 10 9 1 10 9 11 2 10 2 11 2 2 13 1 10 9 10 9 1 11 2 12 2 13 1 10 9 1 9 2
21 9 1 2 11 2 2 11 13 13 1 10 9 2 1 10 11 2 9 0 2 2
13 10 9 13 13 13 10 9 12 12 1 10 9 2
28 1 10 9 1 11 2 11 2 10 9 13 16 15 13 0 2 1 13 3 10 9 1 10 9 1 10 9 2
10 11 13 16 10 9 3 13 12 9 2
18 1 10 9 2 1 12 2 11 13 1 10 9 7 13 10 9 9 2
17 1 2 11 2 2 11 13 10 0 9 0 7 15 13 1 9 2
36 2 15 13 10 13 7 0 9 2 1 15 13 15 10 11 2 15 3 1 11 2 11 2 11 2 2 11 2 7 15 13 2 13 0 2 2
42 10 9 2 13 10 9 2 13 10 9 1 9 15 13 1 10 9 10 9 1 9 2 15 13 10 9 1 9 15 13 1 10 9 2 3 13 1 10 11 7 11 2
23 13 10 15 16 9 2 9 7 9 2 9 1 9 0 16 10 9 7 0 16 10 9 2
26 10 9 0 13 1 9 12 9 1 9 12 9 2 9 1 9 3 1 10 9 0 3 1 10 9 2
24 10 9 0 2 13 10 9 0 2 13 1 9 12 9 1 12 2 1 9 12 9 1 12 2
31 10 9 0 1 9 13 10 9 1 12 5 1 10 9 1 9 13 13 1 12 9 1 12 1 12 9 1 10 9 13 2
35 10 11 2 15 13 10 9 2 13 10 9 13 1 12 5 1 12 1 12 5 1 12 2 9 1 10 9 1 12 5 1 10 10 9 2
38 1 10 9 1 10 9 2 11 13 16 10 9 13 1 10 9 1 10 9 2 13 1 13 3 12 5 1 10 9 2 1 10 9 1 10 9 11 2
2 9 13
44 10 11 2 0 2 13 12 1 10 12 9 13 1 13 1 9 1 9 12 9 1 13 10 9 1 9 1 10 9 1 10 11 2 1 11 2 13 1 10 9 1 10 9 2
2 9 13
21 10 11 13 9 1 10 9 1 11 13 16 10 9 1 9 1 9 13 10 11 2
30 10 9 13 12 9 1 9 1 10 10 1 10 12 9 3 0 1 10 11 9 0 2 9 2 9 2 9 7 9 2
46 10 0 9 1 10 9 13 10 9 2 1 12 2 1 10 11 2 1 10 10 9 7 1 10 9 2 15 13 10 9 0 1 10 9 2 9 2 9 2 9 7 9 1 10 11 2
21 1 10 9 15 15 13 2 9 2 2 12 5 3 13 9 13 1 10 9 0 2
17 13 3 0 16 15 15 15 13 9 7 1 9 2 12 5 2 2
26 13 1 16 13 1 10 9 1 10 9 1 10 9 1 9 2 12 5 13 3 7 12 5 13 3 2
35 13 1 16 11 13 10 0 9 2 10 9 13 13 10 9 2 13 15 13 2 1 2 3 1 10 9 0 2 13 15 13 1 10 9 2
27 13 1 10 9 2 11 2 2 11 13 13 1 10 9 1 15 13 9 1 10 9 1 9 1 10 9 2
7 9 13 1 12 9 1 9
24 10 11 13 10 9 1 12 1 10 9 15 13 10 0 9 11 2 13 10 0 9 1 3 2
37 10 0 9 13 13 10 9 1 2 9 1 10 9 2 3 15 13 1 10 9 1 10 9 11 2 9 2 2 3 1 10 9 0 1 12 9 2
7 9 13 9 0 1 9 0
30 15 3 3 13 10 9 7 13 13 10 9 1 10 9 0 13 13 1 10 9 1 9 0 13 1 10 9 1 11 2
33 3 13 1 9 0 2 10 9 13 13 1 10 9 7 13 10 9 1 13 0 7 13 9 0 16 13 1 15 1 9 1 9 2
34 10 9 1 10 9 2 1 11 2 13 13 10 9 0 7 10 9 1 9 1 10 9 13 2 9 13 1 9 1 9 7 9 2 2
18 12 1 10 9 13 10 9 1 10 9 15 13 1 9 1 13 9 2
13 3 2 10 9 1 9 3 13 13 1 10 9 2
22 10 9 3 13 1 10 9 13 2 13 7 13 10 9 7 10 9 1 10 9 0 2
23 7 15 3 13 9 1 10 9 1 10 9 1 9 0 1 10 9 2 13 10 9 0 2
18 10 9 3 13 1 10 9 1 10 11 7 3 13 13 1 10 9 2
34 15 13 13 2 3 2 0 9 1 9 7 12 9 1 9 2 7 3 13 9 0 1 10 9 2 13 16 13 9 1 1 12 9 2
39 10 9 15 13 3 12 9 1 9 12 1 13 10 9 1 9 0 13 1 13 10 9 1 9 1 10 9 13 1 10 9 7 13 10 9 1 9 0 2
42 10 9 3 13 9 2 13 1 10 0 9 1 10 9 11 2 15 13 10 0 9 2 1 10 11 2 1 10 9 1 10 0 9 13 1 10 9 7 1 10 9 2
9 11 13 2 10 9 1 10 9 2
27 3 13 15 15 10 9 13 3 9 0 1 10 9 2 3 15 13 2 0 2 2 13 1 10 10 9 2
15 1 10 9 2 10 9 13 9 1 13 10 9 10 9 2
15 11 13 16 10 9 0 13 3 10 9 1 10 0 9 2
21 2 13 10 9 1 3 13 15 2 2 13 11 2 9 1 9 1 10 9 11 2
26 10 9 13 16 13 10 9 1 10 9 2 1 11 2 15 3 13 13 16 10 9 13 0 7 0 2
16 3 2 13 1 13 16 10 10 9 13 2 0 2 2 2 2
11 13 16 15 2 13 2 3 3 10 11 2
14 7 15 13 1 13 3 13 1 13 10 9 1 9 2
20 1 10 9 2 10 9 3 0 13 13 10 9 0 7 10 9 1 10 9 2
8 15 13 13 9 1 13 15 2
17 10 9 11 2 11 2 3 3 13 13 1 10 9 1 10 9 2
22 9 1 10 9 2 11 13 10 9 13 10 9 1 11 2 1 12 1 9 1 12 2
30 10 9 1 11 2 11 2 11 2 2 7 10 9 13 1 10 11 1 10 9 2 11 2 3 3 13 13 10 9 2
6 11 13 4 13 1 11
25 11 13 16 13 2 10 9 2 13 1 9 2 1 11 2 9 1 12 13 16 13 3 15 1 12
24 10 9 11 13 13 10 9 0 11 9 1 10 11 1 10 0 9 2 9 2 1 10 11 2
23 10 9 11 13 3 16 10 9 0 13 13 3 10 9 1 10 9 15 15 13 3 0 2
16 10 9 1 9 1 10 9 11 3 13 9 1 10 9 0 2
54 10 9 1 9 2 3 15 1 10 0 9 2 13 12 9 1 9 1 9 2 1 9 1 9 1 9 0 7 0 2 2 9 2 9 2 9 2 9 2 13 1 10 9 2 2 9 0 2 9 1 9 0 3 2
13 10 9 1 10 1 10 11 13 13 3 1 11 2
15 2 13 16 15 3 13 10 11 3 1 13 13 3 2 2
11 11 2 13 2 1 10 11 10 9 0 2
34 10 9 13 13 1 10 0 9 10 9 1 9 1 10 0 9 15 13 13 3 2 1 10 0 2 2 1 10 10 9 7 9 2 2
5 11 13 9 1 11
7 2 9 2 13 9 7 9
22 1 3 10 9 1 9 1 10 11 13 9 0 1 10 9 0 11 2 2 9 2 2
25 10 9 13 9 1 10 9 2 11 2 1 10 11 2 15 13 10 9 0 1 9 1 10 9 2
14 10 0 1 10 9 11 7 11 13 1 9 10 9 2
13 2 13 16 10 11 13 0 1 15 15 13 13 2
27 10 9 13 13 10 9 3 0 1 10 9 16 13 4 13 1 10 9 2 2 13 11 2 1 10 11 2
26 1 10 9 11 2 1 10 11 2 2 3 10 9 0 13 13 10 9 1 10 9 1 10 9 2 2
25 1 11 2 10 9 1 10 11 13 9 1 10 9 13 2 1 10 9 13 2 1 10 9 11 2
6 9 13 12 5 1 11
30 10 11 2 11 2 1 11 13 10 0 9 1 9 1 9 1 12 5 2 1 15 12 5 13 1 0 9 1 9 2
18 1 9 1 10 9 0 2 3 10 11 13 1 12 5 2 13 9 2
27 10 9 13 1 10 11 2 11 2 7 13 10 9 1 10 9 1 9 1 12 1 12 9 0 1 11 2
29 10 11 2 1 9 1 9 1 12 1 12 9 2 13 1 12 5 2 1 15 12 5 1 10 10 9 1 9 2
30 13 2 3 2 10 9 3 3 0 1 10 9 1 10 9 7 3 0 2 0 7 0 2 1 10 9 1 10 9 2
23 13 10 9 1 9 7 9 15 15 11 7 11 13 2 7 15 10 9 3 13 1 9 2
10 11 2 12 2 13 0 1 10 11 2
8 10 9 1 10 9 13 0 2
20 2 11 2 13 10 0 1 10 11 2 9 13 1 11 1 10 9 1 12 2
48 11 2 9 2 2 11 2 0 2 2 11 2 9 2 7 11 2 9 2 13 1 10 9 1 10 9 2 10 9 1 11 2 9 1 9 7 10 9 1 10 9 13 0 7 0 1 11 2
20 1 10 9 15 10 9 13 13 2 11 2 2 2 11 2 7 2 11 2 2
4 11 2 9 2
9 13 16 10 10 9 3 13 13 2
15 13 10 9 0 1 10 9 0 2 0 2 13 7 0 2
24 15 3 13 16 2 1 10 9 2 15 13 10 9 1 10 0 2 0 7 0 9 1 15 2
18 1 10 9 1 10 9 1 10 9 2 3 13 10 9 1 10 9 2
11 10 9 13 9 2 9 2 9 7 9 2
8 10 10 12 9 3 13 13 2
14 10 9 13 16 13 15 13 0 10 9 1 10 9 2
13 13 15 13 3 1 11 2 11 2 11 7 11 2
24 1 10 9 1 11 2 13 1 12 10 9 1 9 13 1 10 11 1 10 9 1 10 9 2
7 9 13 1 9 1 10 11
46 10 9 1 10 9 1 10 0 12 9 13 1 16 10 9 0 11 13 0 9 1 9 1 9 2 9 7 9 0 1 9 1 10 9 13 1 10 11 2 1 10 9 1 10 11 2
40 10 9 11 13 1 10 9 1 12 12 9 2 7 10 11 2 9 1 9 1 10 9 7 9 1 11 1 10 11 1 11 2 1 10 9 1 13 10 9 2
15 1 10 9 2 11 13 10 9 1 10 9 1 10 11 2
10 15 13 16 10 9 13 2 0 2 2
8 11 13 10 9 1 0 9 2
17 1 10 9 2 10 9 1 10 9 0 13 16 15 13 10 9 2
8 11 13 9 1 10 9 1 11
23 10 9 7 9 11 13 1 10 9 12 1 9 2 1 10 9 2 10 0 9 1 11 2
17 10 11 13 13 1 10 9 11 2 12 2 1 10 9 1 11 2
16 10 9 1 10 9 1 9 13 13 1 10 11 1 10 9 2
2 10 9
28 12 2 9 13 13 1 10 0 9 2 9 1 9 2 1 16 10 9 1 10 9 1 11 13 10 9 0 2
16 1 10 12 9 2 12 13 9 1 10 11 2 11 7 9 2
21 16 15 13 13 13 2 3 9 2 12 5 2 1 10 9 0 13 13 1 11 2
23 11 2 9 2 9 0 1 9 0 1 10 11 7 9 0 1 9 0 2 9 11 2 2
3 9 0 2
11 11 2 13 13 1 10 9 1 10 11 2
12 13 0 7 9 1 10 11 2 9 11 2 2
40 3 1 10 0 2 9 2 2 10 0 9 15 11 13 2 11 2 7 2 11 2 13 3 1 10 9 1 10 9 2 1 10 9 0 2 1 10 9 0 2
16 1 9 2 13 1 0 10 9 1 10 10 9 1 15 13 2
16 1 2 11 2 2 10 9 7 10 9 13 1 10 9 0 2
31 1 10 11 2 1 12 2 10 9 1 9 2 11 2 11 2 2 13 13 3 9 1 10 9 0 2 11 2 11 2 2
22 15 13 1 10 9 1 10 9 2 1 10 9 1 11 2 15 13 1 10 11 2 2
37 10 9 1 10 11 13 9 1 12 9 2 13 12 9 7 12 9 1 9 2 13 13 10 9 13 1 10 9 2 1 9 7 9 1 9 0 2
33 15 13 10 9 0 13 1 10 9 3 12 9 1 9 1 12 9 2 13 10 9 11 7 10 9 1 10 9 11 1 10 9 2
16 10 9 3 13 10 9 1 13 10 9 1 3 12 12 9 2
20 13 1 10 9 2 10 9 11 15 13 0 1 10 9 0 1 13 10 9 2
34 2 3 13 10 9 0 1 13 1 10 9 0 2 1 11 2 2 15 13 9 1 13 0 2 2 13 10 9 1 9 1 10 11 2
25 10 9 13 1 11 13 10 10 9 15 13 10 0 2 11 2 1 10 9 0 2 13 1 11 2
25 1 10 9 1 10 9 1 3 2 15 1 10 9 1 10 2 11 2 13 15 13 1 10 9 2
14 11 13 16 13 13 1 13 10 9 0 1 10 9 2
22 10 9 1 10 11 2 11 2 13 10 9 1 10 9 1 10 0 7 11 1 9 2
31 2 16 15 13 0 2 10 11 13 1 10 9 10 9 2 7 1 11 15 13 1 9 1 10 9 7 13 10 9 2 2
1 13
8 9 13 9 1 9 1 10 9
35 10 11 13 2 1 10 0 9 2 10 9 1 10 9 1 10 9 2 11 2 1 13 10 9 0 15 13 1 10 9 1 10 9 0 2
30 10 11 2 11 2 2 15 13 1 10 9 2 9 7 9 1 10 9 0 1 9 0 2 13 13 1 10 9 11 2
21 11 7 11 3 13 2 1 10 9 2 15 10 9 13 7 15 13 13 10 9 2
42 3 2 3 10 9 1 15 10 9 13 13 3 1 10 9 13 13 10 9 1 10 0 9 2 13 9 3 11 2 11 2 2 11 2 11 2 7 11 2 11 2 2
13 9 1 10 9 0 3 13 0 9 1 10 9 2
32 11 7 11 13 13 16 10 9 1 10 9 13 0 1 13 10 9 1 10 9 2 1 15 10 9 3 13 10 9 0 0 2
21 1 13 10 9 1 9 2 10 9 13 3 10 9 1 13 10 9 1 10 9 2
23 10 9 1 10 9 13 10 9 1 10 9 0 1 10 9 1 12 9 0 1 0 9 2
17 10 9 13 10 9 0 1 9 12 9 1 10 9 1 10 9 2
20 10 9 2 1 13 9 12 9 2 13 13 1 10 9 1 10 9 1 12 2
13 10 15 3 13 1 10 9 1 9 1 10 9 2
30 1 10 9 1 9 11 2 10 9 13 4 13 1 10 9 13 10 9 1 10 9 2 1 10 9 1 10 9 0 2
26 7 13 15 13 10 9 1 13 1 9 1 10 9 1 16 10 9 13 13 3 13 7 13 10 9 2
3 13 10 9
33 11 2 1 10 11 2 13 10 2 9 2 1 10 9 1 10 9 1 3 2 2 15 13 13 13 10 9 1 10 9 0 2 2
2 10 9
24 9 1 11 2 2 13 3 1 10 9 10 9 1 9 3 13 1 10 9 1 10 9 2 2
20 10 11 13 9 12 9 1 10 9 2 3 1 10 9 1 10 11 2 11 2
22 1 10 0 9 2 1 10 9 12 1 9 2 13 13 3 12 9 1 9 1 11 2
29 11 13 16 10 9 13 1 10 9 13 10 9 1 12 9 1 9 2 9 12 9 2 1 9 1 10 9 0 2
38 1 15 2 10 9 13 16 10 9 13 10 9 1 9 1 12 9 1 9 2 9 12 9 2 7 13 10 9 1 12 9 1 10 9 1 10 9 2
19 1 10 9 2 13 15 16 10 9 1 10 9 13 10 12 9 1 9 2
15 10 9 13 13 1 10 9 1 10 9 1 10 9 12 2
23 10 9 1 10 11 13 15 1 10 9 1 9 1 10 9 1 10 9 0 1 10 9 2
28 10 9 2 13 1 10 0 9 2 13 10 9 1 10 11 1 0 9 2 1 12 5 1 10 9 1 9 2
28 10 9 1 10 9 1 10 9 0 0 13 13 1 10 9 1 10 10 9 15 13 10 9 1 10 9 11 2
7 9 13 10 9 11 7 11
43 10 9 1 10 9 11 2 1 10 11 1 10 11 2 7 11 2 9 0 1 10 11 2 3 9 1 10 11 1 10 9 1 10 11 13 9 1 9 1 10 9 0 2
21 15 13 10 9 1 10 12 9 1 10 9 1 10 9 7 1 10 9 0 0 2
12 11 2 3 13 13 1 10 9 1 10 11 2
13 11 2 13 13 1 9 2 13 16 13 13 0 2
15 13 1 10 10 9 7 13 13 1 10 11 1 10 9 2
7 9 1 9 13 9 1 11
21 9 1 2 11 2 13 1 10 11 1 13 1 10 9 10 9 1 2 11 2 2
23 10 0 9 0 1 10 11 13 3 1 11 10 9 11 2 9 1 10 0 2 11 2 2
7 9 13 13 12 5 1 9
44 10 9 1 9 1 10 11 2 11 2 13 12 9 1 9 2 15 13 10 9 1 12 5 1 9 1 10 9 3 0 2 3 13 13 12 9 2 3 1 9 1 10 9 2
15 10 9 0 1 9 1 10 9 1 9 13 1 12 9 2
25 1 10 10 9 1 10 9 13 2 3 10 9 13 12 9 1 9 2 10 9 13 1 12 5 2
17 10 9 0 1 10 9 13 1 12 9 2 1 9 1 10 11 2
11 2 16 3 13 15 2 10 9 13 3 2
16 10 9 1 10 9 13 13 1 10 9 0 2 2 13 11 2
23 3 1 9 3 0 2 1 12 1 12 9 2 10 9 13 13 1 13 10 9 1 11 2
23 10 11 2 3 2 13 10 9 1 10 9 15 13 10 9 1 10 9 1 10 9 0 2
24 10 11 13 12 9 13 1 10 9 1 9 2 9 2 9 2 9 2 9 2 9 7 9 2
8 1 9 2 13 10 9 0 2
7 2 13 0 1 10 9 2
2 13 2
8 13 10 9 1 15 13 2 2
12 13 1 13 10 9 1 11 7 11 2 13 2
10 2 3 13 13 1 15 15 13 2 2
6 7 13 13 15 13 2
18 1 10 9 1 10 9 7 1 10 9 2 10 9 0 13 13 0 2
18 7 3 15 13 2 1 10 9 2 2 16 3 13 9 1 13 2 2
16 3 11 13 1 10 9 9 1 10 9 13 1 10 9 13 2
26 10 9 2 1 9 2 13 10 9 11 1 10 11 2 15 1 3 12 9 0 15 13 1 10 9 2
16 10 11 13 1 10 9 1 10 11 2 13 3 13 10 9 2
7 3 2 3 13 10 9 2
17 10 9 1 10 9 0 13 13 1 10 12 9 1 10 0 9 2
11 11 13 1 10 9 7 13 1 10 9 2
12 11 13 3 10 9 1 13 1 10 9 0 2
24 9 13 10 0 9 1 10 9 1 10 9 7 10 9 1 10 9 1 9 13 13 13 1 2
9 2 9 2 13 10 9 1 10 9
17 9 2 9 1 12 9 2 13 1 9 1 9 2 1 10 11 2
8 3 2 0 9 2 1 10 9
19 2 11 2 13 10 9 1 9 15 13 4 13 1 9 1 10 9 0 2
53 10 0 1 10 9 13 10 9 1 9 1 9 2 0 2 0 2 0 2 0 2 0 2 7 13 9 13 1 10 9 0 1 10 9 15 13 10 0 9 1 10 9 1 10 9 12 2 3 13 1 10 9 2
12 10 9 1 10 9 13 16 10 9 13 0 2
14 10 9 1 10 11 2 11 2 3 13 1 9 3 2
10 15 13 12 5 1 9 1 9 0 2
14 10 9 1 10 9 13 1 9 1 10 0 9 12 2
17 11 2 10 9 13 1 10 9 2 1 10 9 2 1 10 9 2
17 15 13 13 10 9 1 9 2 3 15 13 1 10 9 1 9 2
7 11 2 3 13 10 9 2
7 9 13 2 9 2 1 9
1 11
24 10 9 11 13 13 10 9 1 10 9 15 13 13 1 10 9 1 10 0 2 13 10 9 2
19 10 9 2 11 2 13 1 10 9 1 10 9 3 7 11 3 13 13 2
8 9 1 10 11 13 13 9 0
20 10 9 9 1 10 11 13 13 1 9 10 9 1 10 9 1 10 9 11 2
14 10 9 1 9 13 9 1 9 2 13 1 10 9 2
21 1 11 2 9 1 9 2 10 9 1 9 13 13 1 10 9 13 1 9 13 2
25 9 1 9 1 9 13 10 9 1 10 12 13 9 2 13 10 9 1 10 9 15 15 10 13 2
26 1 9 2 11 13 1 10 11 1 9 1 10 11 1 11 2 1 13 10 0 9 1 10 9 11 2
10 10 9 13 3 10 0 9 1 9 2
17 1 15 12 2 10 9 1 2 11 2 13 10 0 9 1 9 2
27 2 13 0 15 1 3 2 2 13 13 10 9 0 2 15 13 1 10 9 3 9 1 10 0 9 12 2
39 2 9 0 2 1 10 9 2 10 9 7 10 9 1 9 13 13 3 9 1 2 11 2 1 11 2 9 1 10 11 2 1 10 9 0 1 10 9 2
28 9 3 0 15 3 13 10 9 13 13 9 0 2 9 0 13 7 9 0 1 10 9 2 9 7 9 2 2
15 9 13 13 16 10 9 13 13 10 9 1 10 10 9 2
22 10 9 15 13 1 13 9 13 13 9 1 10 9 7 1 10 9 7 10 0 9 2
5 9 13 13 9 0
19 9 1 10 11 2 15 13 9 0 1 9 0 2 13 4 13 1 10 11
29 3 9 13 1 10 9 0 7 2 3 2 13 1 9 1 11 2 13 3 9 0 10 9 7 9 1 9 0 2
31 10 11 2 9 0 1 10 11 2 13 1 10 9 11 10 9 1 10 9 1 9 1 9 13 9 13 1 13 9 0 2
7 10 9 13 9 12 12 2
23 10 9 1 9 13 0 2 7 3 10 9 15 13 1 13 10 2 9 0 1 9 2 2
52 1 12 1 10 9 3 0 1 10 9 2 10 9 13 1 10 2 9 2 0 1 9 1 9 2 10 9 11 2 13 13 10 9 1 9 0 1 10 9 2 1 11 2 9 1 10 9 0 1 10 9 2
14 10 9 13 13 10 9 1 9 1 9 1 13 9 2
37 15 13 4 13 1 9 13 1 10 9 1 9 0 13 10 9 0 1 10 9 7 1 10 9 0 7 10 9 15 13 13 10 9 1 10 9 2
47 1 11 2 9 13 1 9 2 10 9 13 4 13 1 12 9 2 9 0 1 9 2 0 2 0 2 0 3 2 2 9 0 7 9 1 10 9 1 9 2 9 2 9 2 9 2 2
1 11
30 13 10 9 1 9 2 13 16 2 13 0 9 1 16 9 13 10 9 1 10 9 15 10 9 1 10 11 13 2 2
1 11
34 10 9 0 13 16 10 9 1 10 9 13 10 9 1 9 1 12 9 1 13 10 9 15 13 9 1 13 1 9 1 9 7 3 2
5 11 13 10 0 9
35 10 11 13 10 0 9 1 10 9 1 10 11 2 1 3 12 9 2 2 1 9 2 9 2 1 13 10 11 12 9 1 12 1 12 2
23 3 10 9 11 13 10 9 1 9 1 10 11 2 10 1 10 3 13 9 1 10 9 2
9 15 13 12 9 7 13 12 9 2
12 10 11 13 3 12 9 7 3 13 12 9 2
23 1 10 11 2 10 9 1 10 9 13 11 2 1 12 9 2 13 1 11 2 1 12 2
5 1 10 9 1 9
17 3 2 3 2 10 9 1 10 9 0 13 10 9 1 10 11 2
30 3 2 3 2 3 13 10 9 0 7 10 9 0 10 15 13 10 9 0 1 10 9 0 2 7 3 10 9 0 2
12 7 2 3 2 10 9 3 13 1 10 9 2
30 13 1 12 2 10 9 11 2 9 2 13 10 9 0 0 15 13 9 1 10 9 13 9 1 10 9 1 0 9 2
33 11 13 12 9 1 9 0 7 2 3 1 11 2 13 13 9 1 9 7 2 3 2 13 15 1 10 9 1 10 9 1 9 2
15 13 10 9 2 11 15 13 13 1 10 9 1 10 0 2
22 16 3 13 3 9 3 0 2 10 0 13 13 10 9 1 10 9 2 10 9 11 2
28 10 9 1 10 9 1 9 13 1 10 13 9 2 11 2 2 11 2 2 0 9 1 12 9 1 10 9 2
30 10 9 3 13 16 1 10 9 1 9 10 9 13 1 10 9 10 9 1 10 9 1 10 9 0 1 10 9 0 2
16 16 10 0 13 9 2 10 9 13 16 10 9 3 13 13 2
5 11 13 0 9 0
27 10 11 13 3 10 11 1 11 1 12 1 12 1 11 7 13 10 12 9 1 13 10 9 1 10 11 2
20 10 9 13 15 12 0 13 1 10 11 7 10 9 1 10 11 1 10 11 2
18 1 11 2 3 13 0 13 15 3 1 10 9 1 9 1 0 9 2
13 13 9 1 9 1 9 15 13 10 9 1 9 2
10 1 12 9 7 15 13 13 0 9 2
21 1 10 9 2 11 13 9 1 9 1 13 10 9 7 13 10 10 9 1 13 2
25 1 10 9 1 10 9 13 10 9 1 10 9 2 9 2 9 0 2 9 2 9 0 7 9 2
9 2 13 9 15 13 10 9 0 2
22 13 10 10 9 15 13 16 10 9 0 15 13 1 13 9 2 2 13 11 2 12 2
17 2 13 0 13 10 9 1 10 9 13 2 2 13 11 2 12 2
26 11 13 16 3 1 10 9 1 9 13 10 9 1 2 0 9 2 2 16 3 13 1 10 10 9 2
15 2 10 9 13 0 16 10 9 3 13 10 9 1 15 2
18 15 13 10 9 7 13 10 9 1 9 13 2 2 13 11 2 12 2
14 1 11 2 10 9 13 1 2 9 2 1 9 0 2
34 2 15 3 13 10 9 1 10 9 2 7 13 9 3 9 0 7 0 3 1 9 3 10 9 1 10 11 1 10 9 2 2 13 2
42 1 10 9 0 2 10 11 13 12 2 9 2 2 1 9 12 9 1 9 2 1 16 10 9 1 10 9 13 10 9 1 10 9 3 1 13 10 9 1 10 9 2
9 10 9 13 13 3 1 13 9 2
23 10 9 11 13 3 2 1 11 2 10 10 9 1 10 0 9 0 3 9 1 10 11 2
19 10 9 1 10 11 2 11 2 13 16 10 9 0 13 13 9 1 11 2
24 2 13 3 1 11 16 10 11 3 13 10 9 1 13 10 9 16 15 13 1 10 9 2 2
15 2 10 9 13 10 9 0 1 9 2 1 13 3 13 2
26 10 9 13 13 1 9 1 9 2 9 2 1 10 9 1 9 7 1 10 9 1 9 13 1 9 2
7 11 4 15 3 13 1 9
23 10 9 1 10 11 13 10 2 11 2 2 9 13 1 9 1 10 9 0 2 11 2 2
12 13 12 9 2 12 5 2 1 12 12 9 2
8 11 13 10 0 9 1 10 11
11 10 9 13 3 10 9 1 10 9 0 2
26 1 10 9 2 11 3 13 1 12 5 1 10 9 1 9 1 9 2 12 9 3 1 10 0 9 2
19 1 1 12 9 1 10 9 1 10 9 2 11 3 13 1 15 12 5 2
19 11 13 1 10 0 9 7 13 10 0 9 1 11 2 11 2 11 2 2
35 1 10 9 11 13 1 10 0 9 2 15 0 13 2 11 2 13 1 12 5 2 12 9 0 1 10 9 1 10 9 1 10 10 9 2
23 11 13 16 2 3 13 13 15 2 1 10 0 9 0 13 1 10 9 1 10 9 11 2
31 2 15 13 0 1 10 9 11 2 0 1 10 9 2 0 1 12 9 1 9 2 15 3 13 9 10 1 10 9 2 2
20 1 11 2 2 15 13 16 13 10 9 2 1 10 9 0 2 13 13 2 2
15 10 9 13 16 13 1 10 11 1 16 10 9 13 0 2
16 10 9 13 13 2 1 0 9 2 10 9 1 11 1 12 2
39 10 9 13 16 2 13 9 2 10 9 1 12 3 3 13 13 3 16 3 13 0 10 9 1 10 9 13 1 10 11 2 13 1 9 12 9 1 9 2
3 9 1 12
28 10 11 13 16 11 7 11 2 13 1 10 11 1 10 9 1 9 0 2 13 4 13 1 10 11 1 11 2
25 9 13 1 10 11 2 1 12 9 2 13 9 1 12 5 1 9 1 11 1 10 11 2 11 2
3 9 1 12
23 10 9 0 11 2 0 2 7 11 2 0 2 13 16 10 11 0 13 9 1 10 9 2
19 10 9 13 1 10 9 0 3 1 10 2 11 2 2 13 1 10 11 2
23 13 7 13 0 1 9 0 1 11 2 3 15 1 10 9 2 15 1 10 11 7 9 2
26 10 9 1 10 0 1 11 2 11 2 2 1 11 2 11 2 7 1 10 11 3 13 1 10 9 2
18 1 10 9 2 10 9 13 10 9 1 13 3 10 9 1 10 9 2
48 10 9 13 1 10 9 3 1 10 9 2 9 1 11 2 1 13 1 10 11 2 1 10 0 2 9 1 10 9 2 2 10 9 1 10 0 9 1 10 0 2 13 9 1 10 9 2 2
29 1 10 9 1 10 9 15 13 1 10 10 9 2 10 9 12 2 10 2 11 2 2 13 3 1 10 0 9 2
22 15 13 10 9 0 2 1 9 0 1 9 0 7 0 9 2 0 1 13 13 13 2
12 10 2 11 2 7 10 11 13 3 3 13 2
34 10 2 11 2 13 9 7 9 13 1 9 7 13 3 1 10 9 2 3 10 11 2 3 13 2 13 3 0 7 2 3 2 0 2
24 10 9 11 13 1 9 7 9 0 3 1 10 9 1 11 1 13 10 9 1 10 9 0 2
25 15 13 10 0 9 15 10 9 13 2 1 15 10 9 0 7 10 9 1 9 13 3 12 9 2
13 3 2 13 1 15 13 16 13 0 9 1 9 2
20 3 3 1 15 3 1 10 10 9 3 13 10 9 0 7 0 1 10 9 2
36 3 10 9 13 1 9 1 10 9 0 13 1 9 2 10 9 13 1 10 9 3 10 15 2 13 10 9 15 13 10 0 1 10 0 9 2
9 13 0 16 15 13 13 10 0 2
28 10 0 2 3 2 13 16 1 10 9 10 10 9 13 1 9 7 13 13 10 9 1 10 9 1 10 9 2
15 11 2 10 11 13 9 1 9 3 0 1 10 0 9 2
9 10 9 2 3 2 15 13 13 2
26 11 2 3 13 13 16 15 15 13 2 13 3 16 1 12 9 10 9 1 10 11 13 1 10 11 2
40 3 13 16 10 9 13 3 0 2 1 10 9 1 9 1 9 1 9 2 1 15 13 13 10 9 0 2 15 13 1 12 5 1 12 5 1 10 9 0 2
32 7 16 15 13 1 9 7 11 13 3 2 12 9 7 9 1 9 2 10 9 3 13 10 9 1 10 9 1 11 7 11 2
1 9
24 13 1 12 1 10 11 3 10 9 13 11 2 11 7 11 2 10 9 11 13 1 10 9 2
27 2 15 13 1 13 16 13 1 10 9 1 9 2 2 13 10 9 11 2 0 1 10 9 1 10 9 2
17 1 12 9 1 9 1 10 9 2 12 13 15 0 1 10 9 2
1 9
34 2 13 13 2 2 13 10 9 1 10 9 2 11 2 9 0 1 10 9 1 11 2 11 2 2 11 2 11 7 11 2 11 2 2
57 1 13 10 9 1 3 9 1 10 12 0 1 10 9 9 2 9 2 9 2 9 2 13 7 3 12 9 2 10 9 13 16 16 10 9 15 13 1 13 10 9 1 10 9 2 10 9 13 1 9 10 9 1 10 9 0 2
13 2 10 9 13 3 3 13 2 2 13 9 11 2
33 10 9 1 13 10 9 1 10 9 1 10 9 0 13 13 1 9 1 10 9 1 10 9 1 10 9 2 12 2 12 7 12 2
20 13 1 9 10 9 1 10 9 13 0 13 1 10 9 13 1 15 1 11 2
30 3 3 1 10 9 1 10 1 10 9 3 9 3 10 11 2 10 11 7 10 11 13 3 3 3 16 3 13 13 2
45 1 10 9 1 15 13 10 9 13 2 15 13 10 9 13 10 9 13 13 2 1 9 1 11 2 10 2 9 2 1 10 9 1 9 2 11 2 11 2 11 2 11 2 11 2
24 9 2 10 9 0 13 13 2 3 2 10 9 13 1 10 9 1 10 9 1 13 0 9 2
34 9 2 10 0 9 1 13 10 9 13 11 2 12 2 10 9 13 13 1 10 9 1 3 2 1 13 1 10 9 0 2 11 13 2
21 1 10 9 13 13 10 9 1 13 16 10 9 13 1 10 9 13 1 10 9 2
1 9
17 1 11 2 10 9 1 10 11 3 3 13 10 9 1 9 11 2
21 10 9 15 13 13 10 9 7 2 1 10 9 2 10 9 13 13 1 10 9 2
6 9 13 9 1 9 0
27 10 9 1 9 0 1 10 11 1 10 9 13 13 10 9 1 9 0 1 9 1 10 9 1 10 11 2
22 10 9 13 13 10 9 3 0 1 9 1 10 9 0 1 10 0 9 1 10 9 2
20 10 0 9 1 10 9 13 3 7 13 1 10 9 12 1 11 2 11 2 2
8 9 13 1 10 9 9 1 9
52 10 0 9 13 1 10 9 1 9 1 12 9 0 1 11 13 13 1 10 11 10 11 2 1 10 9 1 9 1 9 0 2 9 0 15 13 9 0 2 9 1 10 9 0 7 9 0 1 10 9 2 2
25 10 9 13 13 1 9 13 1 10 11 9 1 9 1 9 1 10 11 1 10 9 1 10 9 2
6 9 1 10 9 12 2
28 10 9 7 9 0 11 13 1 10 11 16 13 1 10 9 10 9 1 10 9 2 1 10 11 1 10 11 2
15 3 13 1 10 11 2 15 3 15 13 1 13 9 0 2
10 3 13 1 10 9 11 2 1 11 2
9 3 15 13 9 7 9 1 9 2
18 10 9 11 13 16 15 13 13 1 9 7 13 13 10 9 1 9 2
11 2 10 9 2 10 15 9 1 13 2 2
22 10 9 13 1 10 11 7 13 3 12 9 1 10 9 1 10 9 2 1 10 11 2
15 1 10 9 2 12 9 13 13 7 13 13 1 10 11 2
4 15 13 3 2
83 3 2 13 15 10 9 3 0 2 3 3 13 1 10 9 0 1 10 9 13 2 10 9 13 13 15 15 13 1 10 9 1 2 9 0 7 0 2 2 13 10 9 2 0 2 7 10 9 0 1 15 13 15 10 9 13 1 10 9 7 1 10 2 9 2 2 10 9 0 2 13 2 2 10 9 0 7 3 2 10 9 0 2
46 10 9 2 3 0 2 13 1 10 9 13 1 10 9 14 12 1 10 11 2 11 2 2 13 1 10 11 2 15 13 10 2 9 2 7 13 13 10 13 9 1 10 2 9 2 2
26 15 13 0 9 1 13 10 9 0 7 10 9 0 1 10 9 0 1 10 11 2 13 10 9 0 2
62 3 9 1 10 9 11 2 15 1 12 9 1 10 9 1 10 9 13 10 9 1 10 9 7 13 1 9 1 11 2 9 1 11 2 2 13 16 10 9 1 11 13 1 13 10 9 1 10 9 2 15 13 9 1 10 9 11 13 10 10 9 2
27 10 9 1 13 0 9 3 1 10 9 3 13 2 3 2 16 13 0 7 0 13 10 9 1 10 9 2
18 15 13 1 0 9 1 9 0 2 15 13 3 1 13 0 1 13 2
57 3 2 16 10 9 13 1 10 9 1 16 13 1 10 0 13 2 13 7 13 1 10 9 13 1 10 9 10 9 15 13 10 9 2 13 15 3 3 0 13 15 13 1 10 9 1 10 9 1 10 9 13 1 10 10 11 2
9 1 15 2 3 13 9 1 9 2
16 13 2 13 0 2 10 10 9 1 10 9 1 10 0 9 2
19 7 2 3 1 13 3 10 9 1 10 9 2 11 13 4 1 13 3 2
19 10 0 11 2 11 2 7 11 2 11 2 13 2 7 10 9 15 13 2
16 13 0 13 10 9 1 15 2 13 2 13 3 10 0 9 2
23 2 13 1 9 7 13 13 13 9 1 9 7 15 15 13 3 7 1 9 1 9 2 2
16 10 9 1 11 13 1 3 10 9 1 10 9 1 10 11 2
7 13 15 1 10 9 0 2
9 11 3 13 1 10 9 1 11 2
11 13 1 15 10 0 9 1 9 1 9 2
7 3 2 3 13 4 13 2
6 10 9 13 1 9 2
9 7 10 9 3 0 3 13 13 2
7 3 13 13 15 1 9 2
18 3 15 13 1 10 9 1 10 9 15 13 3 2 1 13 10 9 2
6 15 13 3 10 9 2
21 10 9 13 16 10 9 15 13 4 13 1 10 9 3 13 4 13 1 9 0 2
20 3 12 9 13 1 10 9 1 10 9 0 1 10 11 2 3 10 9 13 2
26 9 1 10 9 0 13 13 10 9 1 10 9 13 9 1 9 1 10 9 1 10 9 1 9 0 2
36 1 11 2 12 9 0 2 9 0 2 13 13 3 3 1 10 9 0 2 11 2 2 15 13 10 9 1 11 7 11 1 13 13 10 9 2
8 10 9 3 13 1 4 13 2
24 16 13 15 13 1 10 9 2 3 13 13 10 15 1 10 10 9 2 3 13 3 1 11 2
18 13 1 9 2 1 0 9 2 13 13 10 9 1 11 1 10 11 2
6 9 13 9 1 10 11
30 10 9 11 7 11 13 3 2 1 9 13 1 10 11 2 11 2 2 16 13 9 1 10 9 1 10 11 7 11 2
33 10 11 7 10 11 13 13 1 11 2 0 1 10 9 0 2 1 13 10 9 0 1 10 9 1 10 11 1 10 9 2 11 2
29 1 10 9 2 1 9 7 9 2 3 10 9 0 1 9 13 12 9 2 10 9 1 10 9 13 13 1 9 2
27 1 10 9 3 0 2 3 10 9 3 13 1 12 9 1 9 2 10 9 13 9 2 15 13 10 9 2
14 1 10 10 0 9 2 11 13 9 12 9 1 9 2
14 1 15 13 10 9 11 2 9 7 9 0 1 11 2
38 10 9 1 10 9 1 10 11 2 11 2 13 16 10 9 1 9 13 13 16 11 3 13 13 1 10 9 13 1 16 15 13 10 0 9 1 9 2
23 3 10 9 1 9 1 9 0 2 1 10 9 1 10 11 2 13 13 12 9 1 9 2
30 13 15 10 12 9 2 13 15 1 12 9 1 9 2 3 12 5 1 10 12 9 1 9 0 9 13 1 10 9 2
38 3 1 10 9 1 12 1 12 1 10 0 9 1 10 12 9 2 9 1 10 11 2 10 9 0 11 13 10 9 0 1 10 9 0 1 10 9 2
8 15 13 1 9 10 12 9 2
10 2 10 9 1 10 11 13 10 9 2
14 15 13 1 1 1 10 9 7 15 13 2 2 13 2
2 9 12
15 10 9 7 9 0 11 13 13 1 11 10 9 2 11 2
20 15 13 10 0 1 10 9 1 9 0 1 10 9 1 10 9 1 10 11 2
2 9 12
13 10 11 1 10 11 13 13 10 9 0 1 9 2
14 15 13 13 10 9 15 13 1 11 1 10 9 11 2
15 9 13 10 9 1 9 0 15 13 10 9 0 1 9 2
21 3 13 16 10 9 10 13 10 9 1 9 15 13 9 7 1 9 15 13 9 2
9 1 15 13 1 9 2 13 0 2
17 1 15 13 2 13 3 13 10 0 9 13 1 13 10 9 3 2
21 13 3 15 15 13 13 1 10 9 1 15 13 9 1 15 13 10 9 2 3 2
16 7 1 10 9 1 10 9 1 10 9 2 15 13 10 9 2
18 16 15 13 10 9 0 2 3 13 9 13 10 9 1 10 10 9 2
22 1 10 9 13 2 13 13 9 1 10 11 10 9 1 9 1 9 13 1 10 11 2
23 13 1 10 11 2 10 9 1 9 0 2 1 9 7 9 2 13 15 1 10 0 9 2
9 15 3 13 4 13 1 10 11 2
11 15 13 3 1 13 9 0 1 9 12 2
14 1 15 12 2 3 13 13 10 12 9 1 10 11 2
16 10 9 1 13 10 9 1 10 9 13 13 10 9 1 9 2
15 11 13 3 1 9 2 7 3 13 10 0 1 10 9 2
10 3 0 2 13 13 1 10 11 0 2
12 13 3 0 9 7 13 3 13 1 10 9 2
18 10 9 13 1 15 13 2 16 15 1 10 9 13 13 9 1 13 2
16 10 9 13 3 10 0 9 2 9 15 13 0 1 10 11 2
24 10 9 13 16 15 13 10 9 15 13 9 1 13 10 9 1 13 10 9 1 10 0 9 2
14 1 15 2 13 2 13 10 9 1 9 1 10 0 2
29 1 15 15 13 13 10 9 0 1 10 9 1 10 11 2 10 9 1 11 3 13 4 13 1 9 7 9 0 2
44 1 12 9 2 3 2 10 9 1 10 9 2 15 3 3 13 13 1 13 10 11 7 13 10 9 2 3 2 10 9 1 10 2 9 0 2 1 10 9 3 15 13 9 2
13 10 0 9 13 1 10 9 1 11 2 1 12 2
9 3 1 15 2 13 1 10 9 2
7 10 9 13 13 3 0 2
29 10 9 2 11 2 13 1 10 11 1 9 2 1 11 2 16 11 3 13 9 1 13 10 9 0 1 10 11 2
15 1 10 0 9 2 1 10 9 2 11 2 2 11 13 2
13 2 13 16 3 13 10 9 1 13 3 3 3 2
18 1 10 11 2 13 13 1 10 9 7 1 10 9 1 10 9 2 2
29 13 13 16 7 10 9 2 7 10 10 9 1 15 2 13 1 10 9 13 1 11 10 9 15 15 13 3 15 2
28 10 9 1 10 10 9 13 2 3 2 1 10 9 2 10 1 10 9 1 9 1 10 11 7 1 10 11 2
25 3 13 10 0 9 2 7 13 3 13 10 0 2 16 11 7 10 9 15 13 1 10 10 9 2
8 10 0 13 12 9 1 15 2
30 13 3 13 16 11 13 1 9 0 1 10 9 11 2 13 10 9 1 9 1 10 9 15 15 13 7 15 15 13 2
29 1 15 2 10 9 3 13 13 1 10 9 0 1 10 9 2 11 2 15 3 13 10 9 1 9 1 10 9 2
19 11 13 1 10 9 9 0 2 10 15 15 13 1 13 10 11 1 3 2
35 3 13 13 2 3 2 15 13 10 9 15 11 13 3 13 1 10 9 2 1 10 9 1 16 13 9 1 10 9 1 13 10 9 0 2
21 10 9 11 2 15 13 9 1 10 11 2 3 13 1 13 10 9 9 1 11 2
20 7 13 9 1 10 9 1 10 9 2 3 10 9 11 2 15 13 10 9 2
16 1 10 9 3 3 0 2 1 10 9 11 15 13 0 9 2
8 1 10 10 9 15 13 3 2
38 3 13 13 1 10 9 1 9 2 3 2 13 11 7 11 1 10 9 1 10 9 2 7 15 13 16 10 9 1 11 13 2 1 10 0 2 0 2
13 6 2 11 7 11 13 3 10 9 1 10 9 2
6 3 13 10 0 9 2
15 10 11 13 1 13 10 12 9 1 13 10 0 9 0 2
38 3 11 2 10 0 9 13 1 2 2 9 1 10 9 2 2 2 9 1 10 9 2 2 2 9 1 10 9 2 7 2 9 1 10 9 0 2 2
13 1 13 10 9 2 10 10 11 13 9 1 11 2
17 2 15 13 1 13 1 10 9 0 1 15 1 10 9 11 2 2
4 0 2 13 2
15 2 3 2 1 10 9 13 2 1 10 9 0 13 2 2
8 13 9 1 9 1 10 9 0
26 13 1 10 9 1 10 9 1 10 12 9 10 9 11 2 9 1 10 11 1 9 7 9 1 12 2
18 10 9 13 13 9 1 10 11 2 11 2 2 3 11 13 1 12 2
17 1 10 9 13 3 1 11 2 10 11 13 13 1 10 12 9 2
48 10 11 13 10 0 9 1 10 9 1 9 1 10 9 2 9 7 9 0 2 15 1 10 11 2 13 1 16 10 9 1 10 11 1 10 9 1 10 9 13 9 12 9 1 10 9 13 2
49 10 9 13 12 9 1 10 11 2 2 10 9 1 10 9 1 9 7 9 13 3 0 16 10 1 10 10 9 1 10 11 2 9 3 13 2 7 13 10 9 0 1 10 9 1 9 0 2 2
29 13 1 9 10 11 2 10 11 13 3 10 9 13 3 11 2 9 0 15 13 10 9 1 9 0 1 10 11 2
45 10 11 2 15 3 13 13 1 10 11 3 13 1 9 1 12 7 12 2 13 10 9 1 12 9 1 16 10 9 0 13 1 10 9 1 10 15 10 11 13 9 1 10 9 2
22 3 1 15 2 10 11 13 13 9 0 1 1 12 5 1 10 9 1 10 9 0 2
27 9 1 10 9 0 11 2 2 13 3 0 2 2 2 11 13 10 9 0 3 0 3 1 12 7 12 2
11 10 0 9 1 10 9 13 10 9 11 2
13 15 13 1 10 9 0 1 10 9 1 10 11 2
16 1 10 9 7 10 9 2 10 9 3 3 13 1 10 9 2
7 11 2 9 1 10 11 2
17 2 10 11 1 9 13 10 9 16 10 9 1 10 11 1 9 2
11 15 13 10 9 7 13 10 9 1 15 2
8 7 10 9 13 1 13 9 2
17 10 0 13 16 10 11 3 13 0 7 3 15 13 3 10 11 2
20 16 15 3 13 3 13 13 9 1 15 1 15 13 1 10 9 7 13 2 2
8 9 11 2 9 1 10 11 2
8 2 3 13 10 9 2 9 2
18 10 9 13 10 9 0 7 13 13 1 10 9 1 15 15 15 13 2
19 10 9 1 10 9 13 13 1 10 9 13 10 9 1 10 10 9 0 2
5 13 10 9 2 2
10 10 9 1 10 11 3 13 10 9 2
21 13 3 0 2 13 1 9 2 9 7 9 3 1 10 9 2 13 2 2 3 2
23 10 10 9 1 10 9 2 1 11 2 13 1 2 9 0 1 11 2 11 2 11 2 2
6 13 2 9 0 2 2
31 10 9 13 10 9 1 13 1 10 9 10 9 1 9 10 9 13 10 2 9 2 7 3 1 9 1 10 2 9 2 2
14 2 1 3 10 9 1 9 1 15 2 2 13 11 2
29 2 10 0 2 10 9 2 13 16 13 3 10 9 1 9 2 3 10 0 2 10 9 2 1 13 10 9 2 2
1 13
6 9 13 13 1 12 9
32 10 9 15 10 11 13 13 1 10 9 1 12 9 13 12 9 2 10 11 2 10 11 2 1 10 9 11 2 7 10 11 2
26 3 13 0 13 9 1 10 9 2 1 11 2 12 2 9 0 1 10 9 11 2 15 13 10 11 2
10 9 1 10 9 12 13 12 9 1 11
21 9 1 9 13 1 10 9 2 13 1 9 2 13 4 1 9 1 3 9 12 12
48 10 9 1 13 2 1 9 0 2 13 1 10 9 1 10 11 1 10 9 12 2 13 1 9 1 10 0 9 1 11 1 9 12 12 2 9 0 1 12 9 0 12 9 2 3 10 9 2
16 10 9 13 1 10 9 11 2 1 10 11 2 9 0 2 2
21 11 2 9 1 10 11 2 11 2 0 2 13 13 1 9 1 11 1 10 9 2
13 15 13 10 9 1 10 9 13 1 12 1 9 2
12 13 13 3 9 1 11 2 15 13 10 9 2
34 10 9 2 15 13 13 9 3 1 10 9 2 13 13 10 9 11 2 9 11 2 9 11 7 9 1 10 11 2 3 1 10 11 2
18 1 10 9 2 10 10 9 13 10 9 1 10 9 1 10 9 0 2
13 3 13 13 10 11 2 9 1 9 1 10 11 2
17 15 13 13 1 10 9 1 3 12 9 7 1 13 13 15 12 2
28 10 11 13 3 1 10 9 2 9 1 10 11 2 1 10 11 2 13 9 7 13 1 10 0 9 1 9 2
2 9 13
1 11
38 11 10 9 0 13 1 10 10 0 9 2 15 13 10 1 10 9 0 1 9 2 1 10 9 0 1 9 2 1 10 9 7 9 1 9 7 9 2
17 13 10 9 1 10 9 15 13 10 9 1 10 9 1 10 9 2
9 13 10 9 0 1 15 2 9 2
43 13 16 1 10 0 9 1 10 9 15 13 10 9 1 9 16 13 15 13 10 9 2 10 9 1 10 9 2 10 9 1 10 9 13 1 10 0 9 1 10 9 0 2
16 13 15 15 13 1 10 9 15 13 13 7 13 9 1 9 2
25 3 2 10 9 0 13 3 1 10 9 1 10 0 9 16 13 10 9 2 2 3 2 10 9 2
5 3 15 13 3 2
13 11 2 13 2 3 13 3 0 9 1 10 9 2
15 2 15 13 13 10 9 1 10 9 2 2 13 2 13 2
6 10 9 13 0 13 2
12 11 2 9 1 9 2 9 1 9 7 9 2
9 10 9 2 9 7 9 0 3 2
4 9 13 10 9
7 9 7 9 3 15 13 2
19 15 13 10 9 15 13 1 10 9 1 10 9 1 10 9 0 1 9 2
19 3 10 9 11 2 11 2 13 10 10 9 1 10 9 0 1 10 9 2
11 11 13 13 1 10 9 11 2 11 2 2
19 2 1 10 9 1 3 2 2 13 1 15 2 13 10 9 1 10 11 2
7 1 9 15 3 13 0 2
18 1 10 9 2 10 9 11 2 13 9 2 13 15 1 10 9 0 2
21 1 10 9 2 10 9 13 1 11 2 11 2 7 10 9 11 13 1 10 9 2
12 11 13 16 2 11 2 13 10 0 9 10 2
34 11 13 9 1 11 2 13 1 12 2 2 15 13 1 3 12 9 10 11 2 9 1 9 1 9 3 9 7 9 1 10 9 0 2
23 10 9 13 15 13 10 9 1 10 9 1 11 7 2 3 2 13 9 12 1 10 9 2
27 3 1 13 3 2 10 9 13 10 9 1 9 7 10 9 1 10 9 1 9 7 15 13 1 10 9 2
23 2 15 13 16 13 1 15 13 15 7 1 3 13 13 7 13 10 9 2 2 13 11 2
18 7 2 3 10 9 13 13 10 9 2 12 10 9 1 10 9 13 2
5 11 3 13 1 9
4 3 1 10 11
14 11 13 10 0 9 0 1 13 10 9 1 10 9 2
14 13 10 2 11 2 2 1 10 9 11 2 1 12 2
9 15 13 0 1 10 10 10 9 2
9 11 15 13 11 7 13 12 9 2
17 3 9 2 13 1 13 7 3 13 13 1 9 2 3 10 9 2
37 1 11 2 16 3 13 13 10 9 0 15 13 1 10 9 1 9 1 10 9 7 9 10 9 1 10 0 9 2 1 15 13 10 9 1 9 2
8 2 3 3 13 1 13 0 2
14 10 9 13 0 7 10 9 13 15 2 2 13 11 2
28 1 15 2 10 0 9 13 0 1 10 9 2 3 10 11 15 13 1 10 9 1 9 13 1 4 3 13 2
26 15 3 13 4 13 16 10 9 7 9 1 9 3 13 4 13 1 10 9 0 1 15 1 10 9 2
1 3
31 10 11 3 3 13 10 13 9 1 10 9 1 10 9 1 13 13 9 1 10 9 1 9 1 9 0 1 10 9 11 2
8 10 11 3 13 13 10 9 2
2 1 9
24 16 10 11 13 9 1 10 9 0 1 10 9 1 11 2 10 0 13 0 1 9 1 9 2
30 7 10 2 11 2 2 12 2 7 3 10 2 11 2 1 9 7 9 2 12 2 13 1 10 9 3 0 2 0 2
20 13 2 11 13 11 1 15 15 15 13 1 0 2 1 0 7 2 0 2 2
24 10 9 7 9 0 1 10 9 0 0 15 13 2 1 11 2 9 7 9 0 1 10 9 2
3 2 9 2
41 10 9 13 10 9 1 9 0 1 3 1 10 9 0 1 10 9 2 9 1 10 11 2 11 2 2 9 7 9 1 9 1 10 11 2 11 2 1 9 0 2
16 2 1 12 9 2 10 9 13 15 13 9 3 1 9 0 2
9 16 13 0 2 10 9 13 13 2
14 1 15 2 15 3 13 13 1 13 10 10 9 2 2
11 15 13 10 9 0 1 10 9 7 9 2
8 1 9 2 13 9 1 10 9
19 10 9 11 13 10 9 1 9 3 12 1 10 9 1 10 10 0 9 2
18 2 13 16 3 13 13 15 15 13 2 7 13 1 9 2 2 13 2
19 11 2 15 15 13 1 10 9 15 13 13 1 10 9 7 1 10 9 2
22 1 10 9 11 2 10 9 0 1 10 9 15 13 1 9 15 13 1 9 1 9 2
12 10 9 13 16 10 9 1 10 9 13 0 2
11 2 10 9 13 0 7 13 13 9 2 2
17 10 9 13 13 15 15 13 1 10 9 1 10 9 12 1 9 2
7 11 13 9 1 9 1 9
23 9 13 13 1 1 12 9 7 13 1 10 10 9 2 11 13 9 0 13 9 1 10 9
19 10 11 13 3 10 0 9 1 9 1 10 11 1 13 9 1 10 9 2
15 10 9 13 4 13 1 12 9 7 13 1 10 10 9 2
32 13 10 0 9 0 1 9 13 1 10 11 1 10 9 1 10 9 2 10 1 10 9 1 13 9 15 13 10 9 0 13 2
34 10 9 1 10 9 13 10 9 1 12 1 10 9 13 1 11 2 10 0 15 13 2 1 10 10 9 2 13 11 1 10 10 9 2
22 16 13 10 9 1 10 11 2 11 15 13 10 0 9 13 1 10 9 1 10 9 2
34 1 9 1 10 9 1 10 9 7 1 9 1 10 9 1 10 0 12 9 1 9 2 10 9 13 13 3 1 9 0 1 12 9 2
24 16 10 9 13 1 10 0 12 9 1 9 2 10 9 13 13 1 10 9 2 1 12 9 2
19 1 10 12 9 2 1 10 9 1 9 13 13 1 10 9 1 10 11 2
25 13 3 0 10 9 2 10 9 1 10 9 7 2 3 2 1 10 11 2 11 2 13 10 9 2
8 13 10 9 1 9 1 9 0
19 10 9 1 9 0 1 9 13 9 1 12 5 13 1 10 9 1 9 2
13 13 13 12 9 1 9 1 12 1 10 9 0 2
16 1 10 10 9 1 10 9 13 10 9 13 3 0 12 5 2
8 10 9 13 13 1 10 11 2
10 1 9 13 13 12 9 0 1 9 2
14 13 1 10 9 0 2 10 0 13 9 1 12 5 2
23 3 2 16 10 9 1 9 13 13 1 10 10 9 1 12 2 13 15 9 1 12 5 2
14 1 10 0 9 1 12 13 13 12 9 1 10 9 2
27 1 10 9 2 9 12 9 13 13 1 10 9 12 9 3 1 9 7 9 1 12 9 7 9 1 9 2
34 1 15 2 13 10 9 7 9 1 10 9 1 10 11 2 9 12 9 2 2 11 2 9 12 9 2 7 11 2 9 12 9 2 2
32 11 13 3 16 10 9 13 10 9 1 9 1 9 1 10 9 7 16 9 12 9 13 4 13 3 1 9 1 10 0 9 2
43 1 13 16 10 9 13 10 9 7 10 9 1 10 9 0 2 10 9 13 1 13 9 1 15 9 2 15 15 13 1 10 9 1 10 10 9 2 1 3 10 9 11 2
19 1 10 9 15 13 1 10 9 1 10 9 2 10 9 13 1 10 9 2
10 9 0 13 13 1 10 9 1 9 2
8 9 13 13 9 1 9 1 9
31 10 11 13 3 16 13 13 10 9 1 10 9 11 15 13 10 9 1 9 1 9 1 9 1 15 13 0 1 10 9 2
16 10 9 13 13 1 10 2 11 2 1 10 9 12 1 9 2
31 1 10 9 0 1 10 10 0 9 2 15 13 16 10 9 3 13 13 2 9 1 9 0 2 1 9 1 10 9 2 2
8 10 9 13 3 7 13 0 2
48 3 13 1 10 9 1 9 2 9 1 9 7 9 15 13 1 3 13 10 9 1 10 9 1 10 9 1 9 2 3 1 13 9 7 9 0 2 1 13 10 9 3 0 1 10 9 3 2
27 10 9 1 10 9 13 9 2 13 13 15 1 10 9 0 2 10 9 7 9 1 10 0 1 10 9 2
23 10 0 13 2 1 0 9 2 10 9 7 10 9 2 3 16 15 13 9 1 9 0 2
19 3 13 13 15 2 3 2 13 15 10 10 9 2 3 13 3 12 9 2
25 3 13 1 9 9 13 7 0 15 13 1 10 9 3 9 1 9 7 1 15 3 9 1 9 2
32 10 0 13 3 2 3 2 16 12 9 13 15 1 13 10 9 1 3 12 5 1 10 9 13 1 10 9 7 1 10 9 2
45 13 13 2 16 10 0 3 13 3 1 10 13 9 1 9 1 10 12 9 2 15 13 3 1 10 9 1 10 0 9 0 2 3 3 15 13 3 0 7 15 13 1 15 3 2
15 10 11 13 3 10 9 0 7 13 10 9 1 10 11 2
11 16 15 13 2 13 15 1 9 3 0 2
34 3 2 16 15 13 13 10 9 2 3 2 13 13 9 2 7 15 2 7 13 15 13 13 1 10 9 7 10 9 15 13 4 13 2
21 10 9 1 10 9 3 13 4 13 1 10 9 2 13 10 9 1 9 7 9 2
5 11 13 9 12 9
42 10 9 1 10 9 0 0 7 13 11 2 12 2 13 13 9 12 9 1 10 9 1 11 3 9 1 10 9 1 10 9 15 13 1 12 9 0 1 9 1 12 2
32 10 9 1 9 1 12 1 10 9 13 12 9 1 9 0 1 11 15 13 1 12 9 2 12 13 7 9 12 9 1 9 2
21 10 9 2 10 9 1 10 9 0 2 10 0 9 0 7 10 3 0 13 3 2
12 15 13 13 1 10 9 15 13 1 10 11 2
6 2 13 2 13 2 2
22 10 3 0 13 15 2 7 3 10 9 15 13 2 1 2 13 0 2 10 0 0 2
5 13 10 0 9 2
12 10 0 11 13 13 2 3 2 13 10 9 2
30 3 10 9 1 10 9 13 11 2 10 9 13 13 1 9 0 7 9 2 13 15 2 1 13 10 9 1 10 9 2
26 10 9 13 16 13 13 9 0 1 10 9 1 13 13 10 9 7 16 10 11 13 3 13 10 9 2
26 1 13 10 9 1 10 9 2 10 11 13 9 7 9 15 13 1 10 9 15 1 10 0 9 0 2
15 15 13 1 12 9 2 10 0 2 10 9 7 10 9 2
23 1 10 9 1 15 2 10 9 13 0 7 13 10 9 1 10 9 1 9 0 7 0 2
24 1 10 9 1 9 1 9 1 12 2 3 2 10 9 13 1 13 12 5 1 0 12 5 2
9 10 9 13 1 10 9 2 9 2
11 1 10 0 2 10 9 13 10 9 0 2
17 10 9 13 13 10 9 1 10 9 7 13 13 15 1 10 9 2
27 1 10 9 1 12 9 2 1 9 2 9 2 9 7 9 2 15 13 13 1 10 9 2 13 9 3 2
2 13 13
16 10 11 13 10 9 1 10 12 9 1 10 9 1 10 11 2
11 10 12 9 1 10 9 13 1 10 9 2
4 9 1 10 9
20 11 2 9 0 1 10 11 2 13 1 10 11 1 9 1 9 1 10 9 2
7 3 13 15 13 1 11 2
6 2 10 9 13 0 2
10 16 3 13 15 2 13 13 10 9 2
21 10 10 9 3 13 9 2 2 13 10 9 1 11 1 10 9 1 11 2 11 2
19 10 9 13 3 10 9 1 9 1 10 9 2 1 10 9 1 10 11 2
14 13 0 9 1 10 9 2 7 9 0 9 7 9 2
9 15 13 15 1 10 9 1 10 9
22 11 2 9 7 9 1 9 2 12 2 2 13 10 0 9 0 1 9 1 10 11 2
8 1 12 2 13 9 1 9 0
20 11 2 9 15 13 1 10 9 12 1 15 12 7 13 10 9 0 1 9 2
9 11 3 13 13 16 3 13 11 2
43 10 9 13 10 9 7 10 9 2 1 10 0 9 2 13 12 9 2 12 9 7 13 12 13 1 10 9 12 1 10 9 2 15 13 13 1 2 9 1 10 9 2 2
30 3 1 10 9 2 10 9 1 10 9 2 11 2 13 16 10 9 1 10 11 2 11 2 13 10 9 1 10 9 2
5 11 13 12 9 0
12 9 0 13 1 9 10 12 9 0 1 9 2
19 2 11 2 2 11 2 7 2 11 2 2 11 2 13 13 1 10 11 2
18 2 11 2 13 13 1 9 15 13 1 10 0 9 1 10 0 9 2
10 10 15 1 10 9 13 13 9 12 2
17 13 3 10 10 9 2 15 13 3 9 1 9 1 9 1 9 2
22 10 0 9 1 10 9 2 12 9 2 3 13 13 1 10 9 1 9 1 10 9 2
16 10 0 13 13 1 9 2 9 7 9 1 9 1 10 11 2
28 10 9 2 15 13 3 12 9 1 9 2 13 16 13 1 10 9 1 9 2 3 3 0 2 1 10 9 2
25 13 1 15 10 9 1 11 2 1 9 3 2 3 1 10 11 2 1 10 9 0 1 10 11 2
30 15 13 10 9 2 15 13 13 3 3 2 15 13 10 9 1 12 1 10 9 3 0 7 0 1 10 9 2 11 2
23 15 13 15 13 7 15 13 10 9 1 15 13 1 13 10 9 1 10 9 1 10 9 2
17 11 13 10 9 1 13 10 9 1 10 0 15 3 13 13 9 2
9 7 9 13 9 2 15 13 9 2
19 3 2 1 10 9 1 11 2 13 10 9 1 9 1 9 1 10 11 2
34 7 3 1 10 2 9 2 0 0 2 10 9 11 13 10 9 1 10 9 1 10 11 1 10 9 1 10 9 1 3 12 12 9 2
24 2 3 13 1 10 9 2 7 3 13 13 1 10 9 2 2 13 11 1 10 9 1 11 2
12 3 2 10 9 3 15 13 1 10 0 9 2
21 2 10 10 9 13 13 1 12 9 2 2 13 11 2 9 1 11 1 10 11 2
18 11 13 16 13 3 1 13 10 9 0 1 10 9 1 10 0 9 2
9 11 13 10 2 9 0 2 1 11
24 10 9 11 13 13 10 2 9 1 9 2 3 2 1 10 9 2 1 10 11 2 1 11 2
14 2 13 15 3 13 1 10 9 2 13 10 9 0 2
10 2 13 13 10 9 1 10 9 2 2
10 15 13 0 10 9 1 10 9 11 2
17 10 9 13 3 10 9 1 9 1 0 1 12 9 15 13 9 2
18 2 15 2 1 3 0 16 13 2 13 13 1 10 9 1 10 9 2
13 0 1 10 9 2 13 16 13 10 9 0 2 2
10 10 9 13 12 5 1 9 1 12 2
2 10 9
33 10 9 1 10 9 0 2 13 1 10 2 11 2 2 13 16 13 10 9 1 9 0 7 0 16 1 10 9 1 9 7 9 2
25 1 10 9 1 11 2 10 9 1 10 11 13 15 1 13 10 9 0 2 10 9 2 10 9 2
18 1 10 9 2 13 15 1 10 9 1 15 15 13 1 10 9 12 2
29 3 1 10 9 2 1 10 9 3 15 13 1 13 10 9 15 13 10 9 0 2 3 2 11 2 13 10 9 2
17 10 9 13 1 10 9 1 15 10 9 1 9 13 13 0 3 2
16 11 3 13 1 10 9 3 13 2 9 2 9 3 3 2 2
13 7 3 1 15 2 11 2 13 1 12 9 13 2
28 2 13 1 9 7 0 2 2 13 11 2 1 9 1 9 1 9 1 9 2 1 10 9 13 1 10 9 2
10 11 2 10 9 1 9 13 10 9 2
16 11 2 13 7 15 13 13 3 2 1 10 9 1 15 13 2
15 1 15 2 10 9 13 3 13 3 16 13 10 10 9 2
8 13 12 9 3 1 10 9 2
26 10 9 15 9 0 7 0 3 13 13 10 9 1 10 9 1 10 9 0 13 9 1 10 9 0 2
16 10 11 13 1 12 1 10 3 0 9 0 13 1 10 9 2
31 10 9 1 16 10 9 0 13 1 13 2 3 2 9 1 9 13 3 13 10 9 1 10 9 1 10 9 1 10 9 2
1 11
16 1 10 11 2 13 12 9 15 13 13 10 9 1 10 9 2
7 10 9 13 13 1 9 2
32 10 9 1 10 9 1 11 2 9 2 9 12 2 1 10 11 2 13 16 2 10 9 13 10 0 9 7 10 0 9 2 2
19 3 2 10 9 13 10 9 0 7 13 13 10 9 15 13 1 10 9 2
45 13 15 1 10 9 1 9 13 2 0 1 13 15 1 10 9 1 10 9 0 1 10 9 1 15 10 9 0 15 13 1 16 3 13 0 2 7 1 16 10 9 13 1 13 2
34 15 13 13 10 0 9 1 13 3 10 9 0 7 2 3 2 13 13 10 9 1 9 0 2 15 1 3 13 10 9 1 9 3 2
6 11 13 13 9 1 9
10 10 11 3 13 3 9 1 10 11 2
25 10 9 13 3 11 1 13 16 15 2 13 1 10 9 2 1 10 9 1 10 0 9 1 9 2
32 3 1 13 2 11 13 10 0 9 1 10 11 2 11 2 2 13 9 15 13 13 2 13 2 1 10 0 9 15 13 13 2
17 3 13 9 0 1 10 9 0 1 10 9 7 15 1 10 9 2
30 15 13 3 1 10 9 2 9 0 2 2 3 2 10 0 13 1 10 11 1 10 0 9 7 9 1 9 7 9 2
16 9 13 9 3 0 7 1 10 9 0 2 1 3 12 9 2
29 3 10 9 13 9 0 1 15 1 10 9 2 7 13 13 15 1 9 2 1 10 9 0 2 1 10 1 9 2
37 1 10 9 13 9 10 10 11 2 10 9 13 1 9 9 2 12 5 2 15 13 3 1 10 9 7 3 1 9 1 10 9 0 1 10 9 2
15 15 13 10 9 3 0 7 13 0 1 13 10 9 0 2
32 15 1 12 2 13 9 0 2 0 7 0 2 15 15 13 10 9 0 13 3 10 9 1 10 9 0 1 9 0 7 9 2
23 3 1 10 9 1 10 9 3 0 2 13 10 11 2 12 5 9 2 12 5 11 2 2
24 15 13 10 0 9 2 9 12 2 13 10 9 0 3 2 0 2 7 1 9 7 9 0 2
33 10 9 13 1 10 0 9 1 10 9 1 10 9 7 10 9 0 1 10 11 2 3 12 9 13 1 10 9 1 10 9 0 2
5 11 13 9 1 9
30 10 9 11 2 12 9 2 12 9 7 12 9 2 2 13 3 16 2 3 1 10 9 2 10 0 9 13 10 9 2
37 2 3 13 9 13 3 1 13 9 1 10 9 2 2 13 10 9 2 15 2 1 10 9 2 3 13 3 9 2 13 13 3 9 1 10 9 2
57 10 9 1 10 11 13 10 11 1 10 9 1 9 1 10 9 7 13 16 10 11 13 9 1 13 1 10 11 2 9 12 9 13 1 3 1 12 2 9 12 9 1 9 7 10 9 12 9 13 3 9 0 2 3 1 10 11
31 3 2 10 11 2 15 13 10 9 0 0 2 3 13 16 10 11 13 9 12 9 1 9 0 2 13 15 1 9 0 2
30 13 15 15 15 13 1 2 9 2 1 10 9 1 9 12 2 3 2 13 15 13 1 10 9 1 9 12 7 3 2
15 16 10 9 13 13 2 10 9 1 9 13 10 0 9 2
11 10 9 1 10 2 9 2 3 13 0 2
51 10 9 13 10 9 0 2 1 15 10 9 1 9 13 1 10 9 1 10 9 0 2 10 9 0 15 13 10 11 2 10 0 9 0 1 10 9 1 10 11 7 3 10 0 7 0 9 1 0 9 2
29 1 10 11 2 10 11 2 1 3 1 10 9 1 10 9 2 13 12 5 1 10 9 1 10 9 1 12 5 2
9 11 13 16 10 9 13 9 1 9
33 10 11 2 11 0 2 13 10 9 1 10 9 1 10 9 1 10 9 1 10 9 1 10 9 1 10 9 1 11 2 11 2 2
28 1 10 0 9 12 2 11 2 12 2 13 13 1 10 9 1 10 9 3 12 9 13 15 13 1 10 9 2
8 15 12 13 1 9 12 12 2
26 2 15 13 10 9 1 15 13 2 1 15 15 1 15 13 2 2 13 2 1 0 9 1 10 9 2
14 13 2 3 2 13 10 9 2 1 9 1 10 9 2
27 11 2 1 10 9 2 13 10 0 1 10 9 15 15 13 9 7 9 1 13 1 10 9 2 3 3 2
3 3 13 9
14 9 1 11 2 11 3 13 3 10 9 2 9 2 2
37 15 15 13 3 13 16 13 9 1 10 9 1 13 15 1 10 9 2 1 10 9 1 11 15 13 13 10 9 1 10 11 3 1 10 0 9 2
3 9 1 9
33 9 1 10 11 3 13 10 9 1 13 10 0 9 0 1 13 9 1 10 9 1 2 13 2 10 9 0 1 10 0 9 11 2
11 2 15 13 3 1 10 9 13 0 2 2
4 9 0 13 13
26 3 13 10 9 0 1 13 10 9 1 2 9 2 2 3 10 9 3 13 7 15 13 1 10 9 2
46 15 13 10 0 9 1 10 0 9 1 9 2 1 15 13 10 9 11 2 11 1 10 11 2 2 11 2 2 11 1 10 11 2 2 7 11 2 9 1 10 11 1 10 11 2 2
9 9 13 10 2 9 2 1 10 9
23 10 0 9 1 10 9 7 9 13 1 10 9 1 9 7 9 1 9 15 13 10 9 2
26 10 10 9 13 1 9 1 12 9 12 1 9 1 10 9 9 7 15 1 9 1 10 9 1 9 2
17 1 10 9 2 15 13 1 10 11 2 13 12 9 1 12 9 2
5 10 11 13 13 2
4 13 12 9 2
17 10 10 9 13 13 12 11 2 10 11 2 12 11 7 10 11 2
8 2 13 0 1 10 0 9 2
17 15 13 0 2 13 10 9 9 1 10 9 2 13 10 9 0 2
7 7 10 9 13 9 2 2
15 2 11 2 1 10 9 1 11 3 10 9 1 10 9 2
9 2 13 9 0 2 3 13 9 2
12 10 11 3 13 9 0 1 13 10 9 0 2
8 1 15 13 3 9 1 9 2
19 11 13 13 3 1 10 9 2 1 13 13 3 2 1 10 0 9 2 2
35 9 1 10 11 13 16 10 9 13 9 1 9 2 9 1 9 2 0 9 1 9 2 3 1 11 7 1 10 9 7 3 1 9 0 2
24 2 13 9 1 9 7 9 15 3 13 13 10 9 2 2 13 11 2 9 0 1 10 11 2
28 10 9 2 1 9 1 9 2 12 9 1 9 1 11 2 2 13 15 13 1 10 11 2 3 13 12 9 2
43 3 10 0 9 13 10 9 1 10 9 2 9 1 9 0 13 13 1 10 9 2 10 9 13 3 2 11 15 13 10 9 1 11 7 3 11 2 13 13 2 13 9 2
17 1 10 9 1 10 9 2 10 9 15 13 1 9 0 2 0 2
18 10 3 0 9 1 9 2 9 7 9 13 2 3 1 10 9 0 2
9 9 0 2 9 7 9 13 13 2
8 10 9 13 10 9 3 0 2
27 10 0 13 1 10 9 1 10 9 7 9 9 1 13 9 0 1 10 9 13 1 13 9 0 1 9 2
7 11 13 9 1 10 9 0
21 9 1 10 9 1 10 9 13 1 10 9 2 9 13 9 12 12 1 9 1 9
28 10 9 15 13 1 10 9 1 10 9 0 2 1 3 2 13 9 1 10 9 1 12 9 1 9 1 9 2
18 10 9 13 1 9 12 12 1 9 2 1 9 1 10 9 1 9 2
39 10 9 13 13 1 10 9 1 3 1 10 9 1 10 9 0 2 9 11 2 11 2 2 15 13 10 9 3 13 1 9 9 0 1 10 10 9 0 2
24 11 15 13 2 13 2 1 10 9 7 1 10 9 1 13 10 9 1 10 9 1 10 9 2
31 1 10 9 2 10 9 1 10 9 1 10 9 1 10 9 1 9 13 1 10 9 1 10 9 2 9 11 2 11 2 2
27 11 3 13 13 10 9 1 10 9 1 12 12 9 1 10 9 1 10 9 1 9 1 9 1 10 9 2
19 10 0 9 13 1 10 9 1 9 1 10 9 2 15 15 13 9 12 2
23 1 10 9 2 15 3 13 15 13 1 10 9 1 10 9 3 1 10 9 1 10 9 2
19 10 9 1 10 9 2 11 2 13 16 10 9 1 10 9 13 10 9 2
28 0 1 10 9 1 10 9 2 13 13 0 2 3 13 7 3 13 2 1 0 2 15 15 13 10 9 0 2
38 10 9 1 11 7 11 13 16 10 9 7 10 9 1 9 0 9 13 10 0 9 1 10 9 7 13 9 15 10 9 1 10 9 3 13 1 13 2
29 11 2 12 2 9 1 11 1 10 11 1 11 2 13 0 1 10 9 1 9 1 11 1 10 11 2 11 2 2
13 13 9 0 1 11 1 10 11 2 9 11 2 2
5 11 13 0 1 9
44 10 9 1 15 10 9 1 10 11 2 11 2 13 1 10 0 9 12 1 9 1 11 2 10 9 0 2 13 4 13 1 10 9 2 13 3 10 9 1 11 2 11 2 2
15 10 9 13 4 13 1 9 7 13 10 9 1 10 9 2
9 10 9 13 10 13 9 1 9 2
7 11 13 10 9 12 1 11
2 1 11
11 13 3 3 1 11 10 9 1 9 9 2
12 10 0 9 13 10 11 2 1 10 9 11 2
28 10 9 15 13 1 10 0 9 1 9 7 9 13 1 10 11 2 15 13 1 10 11 2 1 10 9 12 2
3 3 15 13
40 9 13 1 11 13 3 2 1 9 1 9 2 16 11 2 11 2 13 13 1 13 9 1 11 16 10 9 13 16 13 3 13 10 9 1 9 1 10 9 2
2 9 0
38 3 2 10 9 1 10 11 13 10 9 1 10 9 1 10 9 1 10 9 1 10 9 0 1 16 10 11 13 15 11 13 13 1 10 9 1 11 2
4 9 7 11 12
8 12 9 13 10 12 9 1 11
18 10 0 9 1 10 9 2 11 2 13 11 13 1 10 2 9 2 2
4 2 11 2 2
26 10 0 9 1 11 2 3 1 10 11 2 13 4 13 1 10 9 11 2 1 11 2 1 10 11 2
12 3 10 9 0 13 1 3 12 9 1 9 2
18 1 10 9 2 10 9 1 10 9 13 10 9 1 12 9 1 9 2
10 10 9 1 10 9 13 3 13 9 2
24 10 9 1 10 9 13 12 9 1 9 1 10 9 0 7 3 12 9 1 9 1 9 0 2
28 10 12 0 9 13 2 1 10 9 2 10 10 9 1 13 3 13 10 11 1 10 11 2 15 13 9 13 2
19 13 2 11 2 2 1 2 11 2 2 10 9 13 3 0 16 15 2 2
50 1 10 9 13 1 16 10 9 3 13 1 3 16 10 9 13 10 9 2 10 9 13 10 9 2 0 2 1 10 9 0 2 3 15 2 1 9 2 10 2 10 9 13 10 9 1 11 1 11 2
37 10 11 13 1 13 16 10 0 9 1 10 9 2 11 2 2 1 10 9 1 10 0 9 1 10 9 2 10 11 2 13 10 9 1 10 9 2
11 7 16 3 11 13 1 10 9 1 13 2
21 11 2 10 9 13 2 13 3 13 1 0 9 7 1 10 9 1 13 10 0 2
17 13 10 9 3 16 9 2 7 13 13 3 13 13 10 9 0 2
27 10 9 1 10 9 2 7 2 1 9 2 1 10 9 2 13 3 16 10 9 1 10 9 1 10 9 2
21 10 9 3 15 13 1 16 10 9 13 10 9 1 10 9 7 1 10 9 11 2
26 10 9 13 1 10 0 9 1 12 9 2 10 9 13 9 7 10 9 13 1 2 0 2 13 3 2
16 10 9 13 1 10 9 2 16 13 1 10 9 1 10 9 2
8 11 13 10 9 1 10 11 2
14 10 9 13 9 1 12 9 2 0 1 10 12 9 2
24 15 3 13 4 13 1 10 9 1 10 9 7 13 9 1 12 9 1 10 9 1 10 9 2
38 10 9 13 13 10 9 1 10 9 1 10 9 13 7 13 10 9 15 15 13 1 10 9 7 13 2 1 10 9 2 10 9 1 10 9 1 9 2
27 9 13 13 13 1 10 9 9 1 11 2 12 2 0 9 2 11 2 11 2 2 9 12 2 9 11 2
19 1 9 0 2 13 2 12 2 12 1 9 7 9 2 1 9 10 9 2
16 1 10 9 13 1 10 9 13 10 9 11 7 10 9 11 2
24 1 10 9 3 0 13 15 1 10 9 11 2 15 1 10 9 13 9 13 7 10 9 0 2
13 9 13 3 1 10 11 2 1 10 9 1 11 2
30 10 9 15 13 10 9 1 9 0 1 10 9 13 10 9 11 2 15 13 3 10 9 1 13 10 9 1 10 9 2
16 10 9 1 10 9 13 3 3 1 10 9 0 1 10 9 2
11 10 9 1 10 9 13 3 1 10 11 2
23 2 1 10 9 0 2 3 13 13 10 9 13 0 2 2 13 10 9 11 2 11 2 2
34 10 11 13 10 0 9 0 2 7 13 1 10 12 9 1 10 9 3 13 1 10 9 11 1 11 2 3 15 13 13 1 10 9 2
8 3 2 11 13 10 12 9 2
17 1 10 12 9 2 10 11 13 1 13 1 9 7 13 10 9 2
13 10 11 3 13 13 13 7 13 9 1 10 9 2
32 10 9 1 10 9 13 11 7 10 9 1 10 9 13 11 2 13 1 10 9 1 10 11 2 0 2 1 9 1 10 9 2
30 10 9 13 4 13 1 10 9 0 0 11 2 15 13 9 1 10 9 0 1 12 1 10 9 1 10 9 0 0 2
20 11 7 11 2 13 2 13 13 11 12 9 3 2 7 15 3 13 1 9 2
10 10 9 13 13 7 13 1 10 11 2
24 9 1 10 11 2 3 2 13 9 1 10 9 1 9 0 2 1 10 9 1 9 12 12 2
26 10 9 1 11 2 11 2 2 1 10 11 2 3 13 10 9 1 10 9 0 1 13 9 7 9 2
16 9 0 13 1 10 9 1 13 9 1 9 1 9 1 9 2
52 13 15 13 2 1 10 9 2 7 1 2 0 9 2 2 16 10 9 1 10 0 9 1 9 3 13 2 1 9 2 10 9 15 13 10 9 0 1 10 10 9 0 1 10 9 1 10 9 1 9 0 2
21 3 2 1 10 0 9 2 10 9 13 13 2 16 13 10 9 16 13 10 9 2
23 1 10 0 9 2 10 9 13 1 10 9 15 13 10 9 16 13 10 9 1 10 0 2
23 10 9 1 10 9 1 9 13 10 9 1 10 9 1 10 9 1 9 0 1 10 9 2
66 15 13 4 13 1 16 15 13 16 10 0 9 1 10 9 13 1 9 0 1 10 9 1 10 9 3 13 0 16 10 9 13 1 10 9 1 10 9 1 10 9 1 10 0 9 15 13 1 9 1 9 1 10 9 2 1 2 3 3 2 13 10 9 1 11 2
16 11 2 1 10 9 1 2 11 2 2 3 13 10 9 0 2
14 11 2 10 9 13 12 9 1 10 9 1 10 9 2
11 3 1 13 1 11 2 3 13 10 9 2
30 16 10 9 13 1 9 2 1 9 2 13 16 13 13 10 9 2 13 10 9 2 15 13 1 13 1 10 9 3 2
34 13 3 2 1 10 9 1 9 0 2 13 12 1 10 9 7 3 13 15 15 12 2 13 3 10 9 2 15 13 10 1 10 9 2
25 2 15 13 0 2 16 13 13 10 9 7 3 13 3 9 0 3 15 3 1 9 2 2 13 2
29 10 9 0 1 10 9 13 4 13 3 2 13 10 9 2 16 3 13 10 11 15 13 13 9 0 1 10 11 2
9 9 13 0 2 9 2 1 10 9
14 13 1 9 2 10 9 13 0 9 1 9 1 10 9
26 10 9 0 13 1 13 10 0 2 9 2 1 13 10 9 1 9 3 1 10 9 1 10 9 0 2
24 13 15 1 10 9 1 13 2 15 13 1 13 1 10 9 3 11 2 11 2 11 7 11 2
20 3 3 13 1 10 11 2 10 9 13 13 9 7 13 10 3 0 9 9 2
34 13 1 9 2 10 9 13 9 7 13 1 13 9 0 1 9 0 1 10 9 2 3 9 1 9 2 9 1 9 7 9 1 9 2
30 10 9 2 3 3 13 1 10 9 1 10 11 2 13 16 10 9 0 1 10 9 2 11 2 13 13 1 10 9 2
13 1 9 0 2 11 13 13 7 13 1 10 9 2
22 10 9 13 3 10 9 1 10 9 0 1 10 9 1 10 11 2 0 1 10 9 2
1 11
23 10 9 11 2 11 2 13 1 12 5 1 12 5 2 13 12 9 0 1 10 0 9 2
9 3 13 13 0 9 1 10 9 2
1 11
12 11 2 11 2 13 12 9 2 13 12 5 2
12 10 9 3 13 13 10 9 1 10 0 9 2
31 10 9 1 9 1 10 9 11 13 1 12 9 0 2 1 15 7 1 15 2 1 1 10 11 2 15 13 1 12 9 2
13 10 9 1 10 9 13 1 10 9 11 7 11 2
30 15 15 13 13 7 13 3 1 13 1 3 15 13 1 10 9 15 15 13 13 7 10 9 15 13 1 10 9 0 2
20 1 10 9 15 15 13 2 3 13 1 10 9 2 1 10 9 1 10 9 2
12 7 1 10 10 9 15 15 13 1 13 9 2
27 7 3 13 1 10 9 0 2 13 13 10 9 2 13 9 1 15 7 13 9 1 3 13 9 1 9 2
74 9 13 10 9 1 10 9 1 9 1 9 0 0 1 10 9 0 7 0 2 1 10 9 0 2 1 10 9 0 9 12 2 1 12 1 9 1 12 2 16 2 1 10 9 1 9 1 10 9 1 11 2 11 2 13 13 2 1 9 0 7 1 0 9 2 10 9 1 10 11 1 10 9 2
16 9 13 0 10 9 1 10 9 1 9 0 1 10 9 0 2
16 10 9 1 10 9 15 13 1 10 9 1 10 9 1 3 2
18 1 10 11 7 1 10 11 2 13 15 1 10 9 11 10 0 11 2
24 7 13 3 0 13 3 12 9 0 1 10 9 2 10 1 10 9 2 13 1 11 7 11 2
32 1 10 9 3 0 1 10 9 2 2 11 2 2 10 0 2 10 9 13 13 10 9 1 10 9 1 9 7 1 10 9 2
7 10 9 0 13 10 9 2
20 10 9 13 16 10 9 1 10 11 13 10 9 3 0 1 10 2 11 2 2
18 10 9 1 11 7 11 13 13 1 10 9 1 15 1 11 7 11 2
23 10 9 1 10 9 13 13 15 9 1 10 13 1 10 9 1 11 2 3 2 11 2 2
20 1 15 2 13 13 10 12 9 3 10 9 1 10 9 2 1 13 10 9 2
21 1 10 9 2 13 13 10 9 13 12 9 1 9 1 9 2 9 12 9 2 2
13 1 12 13 12 9 1 9 2 9 12 9 2 2
14 7 1 10 9 0 1 10 9 3 1 12 1 9 2
2 12 9
15 1 11 2 2 3 13 0 10 9 13 1 10 9 2 2
35 1 12 9 2 10 0 9 1 10 9 7 9 0 15 13 13 1 10 9 1 9 1 10 9 1 11 2 16 15 13 13 1 9 0 2
22 10 9 1 10 11 13 13 3 1 10 9 11 15 13 9 1 10 9 1 10 11 2
22 11 13 12 1 10 3 0 9 1 11 2 15 13 10 9 1 10 9 1 10 9 2
19 3 2 3 15 13 13 1 10 9 13 7 3 0 15 10 9 13 13 2
21 3 2 16 13 13 10 9 2 15 3 13 2 3 7 3 2 3 3 15 13 2
10 11 2 12 2 13 0 1 10 11 2
8 10 9 1 10 9 13 0 2
6 11 15 13 9 1 12
22 10 9 0 2 11 2 13 16 13 10 9 1 10 9 1 12 16 13 13 1 12 2
13 3 1 12 9 2 11 3 13 4 13 1 12 2
13 2 13 12 9 7 13 1 15 13 2 2 13 2
7 9 13 12 9 1 10 11
19 12 9 13 12 9 1 11 3 2 1 10 9 0 1 9 2 11 2 2
20 3 13 13 9 1 10 9 16 13 4 13 16 10 9 13 9 1 10 9 2
21 10 9 13 1 10 9 1 10 9 2 15 13 3 13 1 10 2 9 2 0 2
9 13 15 1 10 9 1 10 9 2
17 10 9 0 2 7 3 1 10 9 1 9 0 2 13 10 9 2
11 13 15 1 9 1 13 10 0 9 9 2
17 3 10 9 1 9 1 10 9 13 3 1 15 15 13 10 9 2
29 10 11 13 13 1 10 9 13 2 1 10 9 1 10 9 1 10 9 1 9 1 10 9 11 2 9 0 2 2
17 13 1 10 9 11 2 10 9 13 10 9 2 15 13 13 3 2
5 12 9 13 10 11
23 10 11 13 1 10 0 9 12 9 2 15 13 10 9 1 13 10 9 1 11 7 11 2
20 10 9 1 9 13 1 10 9 7 9 1 9 2 3 10 9 13 12 9 2
20 10 11 13 10 9 1 10 9 1 9 1 10 11 2 9 1 10 11 2 2
8 9 1 9 1 11 3 13 11
20 10 9 1 10 11 13 3 2 1 11 2 1 10 9 1 9 1 10 11 2
11 11 13 1 12 3 9 0 1 10 9 2
12 11 7 11 3 13 1 10 9 1 10 9 2
13 13 3 10 9 1 9 1 9 0 7 9 0 2
26 10 9 13 3 9 1 10 9 7 1 10 9 1 9 2 1 13 1 0 9 10 9 1 10 9 2
17 10 9 1 10 9 13 13 1 10 9 1 13 10 9 1 9 2
32 10 9 1 10 11 13 13 1 16 10 10 9 0 13 10 0 9 1 9 0 1 9 0 2 13 2 3 2 1 9 2 2
15 15 13 2 3 2 16 10 9 0 0 13 13 1 12 2
24 10 9 13 0 1 10 9 2 9 2 1 10 0 1 9 12 9 1 9 0 1 10 9 2
26 1 10 0 9 2 13 10 9 1 9 12 9 1 10 9 1 10 9 2 1 10 9 1 10 11 2
29 11 13 16 10 9 3 13 1 9 0 1 9 2 7 3 1 9 1 2 9 2 2 9 13 3 9 9 2 2
32 15 13 2 3 2 16 10 9 0 13 7 10 9 1 9 1 9 0 1 10 9 13 1 9 12 9 1 10 9 1 12 2
18 1 13 13 10 9 0 2 11 13 3 16 13 13 10 9 1 11 2
24 2 13 3 13 1 10 9 2 7 10 9 11 13 9 3 0 1 13 10 9 2 2 13 2
6 9 13 9 1 10 11
55 10 9 1 10 9 13 2 3 1 9 1 10 9 1 9 2 16 10 9 1 10 9 11 7 1 10 9 13 11 1 9 0 1 9 1 10 9 1 9 2 13 9 0 1 15 15 10 9 1 10 9 13 13 2 2
45 1 10 9 2 2 10 9 0 1 13 10 9 0 1 9 1 10 9 13 9 1 10 11 7 1 10 11 2 1 10 9 1 13 10 9 1 9 13 7 9 1 10 11 2 2
4 9 13 13 9
19 9 1 10 11 13 13 1 10 0 9 0 1 3 13 1 13 1 10 11
32 0 1 10 0 9 1 10 9 11 2 10 9 1 10 11 3 13 10 9 1 10 9 1 3 13 1 10 11 1 10 9 2
21 10 9 13 0 13 10 0 9 1 11 13 1 10 9 1 10 9 7 9 0 2
17 11 13 16 15 12 13 9 1 9 0 1 9 1 10 9 0 2
24 10 9 1 11 13 1 10 9 1 10 9 3 1 10 9 7 1 11 13 1 10 9 0 2
9 10 9 13 16 13 13 10 15 2
15 2 10 15 13 4 13 2 7 13 13 16 13 0 2 2
19 10 9 13 10 9 0 7 10 9 0 7 10 0 9 13 11 7 11 2
28 11 15 13 3 1 10 9 7 13 15 1 10 9 1 10 1 10 9 2 3 2 11 2 7 2 11 2 2
12 3 13 9 10 2 11 2 7 2 11 2 2
12 10 9 1 10 11 13 16 13 13 10 15 2
9 10 0 9 13 13 3 1 9 2
18 1 15 15 13 1 9 0 2 11 13 13 9 0 2 1 12 9 2
31 10 9 13 3 9 1 10 9 2 3 0 2 1 10 9 0 0 7 15 13 1 15 15 13 1 3 0 1 10 9 2
15 15 13 1 13 15 3 2 1 16 15 13 1 9 10 2
14 3 2 13 1 3 16 15 13 13 10 9 1 11 2
18 10 11 13 16 10 9 3 13 13 10 9 2 7 13 9 1 9 2
20 11 2 9 1 10 9 2 13 16 10 9 13 1 9 1 10 9 1 9 2
6 11 13 9 1 10 11
23 3 1 10 0 9 10 11 15 13 10 11 13 1 9 7 13 9 1 9 1 10 9 2
61 10 9 13 1 10 9 11 2 9 0 1 10 9 7 9 1 10 9 2 15 13 13 1 13 10 9 1 10 9 7 1 10 9 13 1 12 9 2 10 9 0 7 10 9 0 1 10 11 12 3 13 12 9 1 10 9 2 15 13 13 2
19 1 15 2 10 9 1 10 11 1 9 1 9 13 0 2 1 10 9 2
10 10 9 13 10 9 0 1 10 11 2
27 13 10 9 0 16 13 13 10 9 2 13 1 2 9 0 2 1 13 2 3 2 3 9 1 9 0 2
15 15 13 1 10 11 10 10 9 1 10 9 1 10 9 2
29 3 2 10 0 9 1 10 9 13 2 2 2 13 10 9 0 1 13 13 3 9 1 9 13 1 9 0 2 2
21 2 13 10 9 0 0 7 15 13 13 1 10 9 0 3 0 2 2 1 11 2
53 10 9 1 10 9 1 11 1 10 11 13 9 3 1 10 12 9 1 11 2 13 1 10 9 13 2 7 13 1 10 12 9 1 11 2 13 1 10 0 9 12 2 3 13 10 9 1 10 9 1 10 11 2
47 0 13 1 10 11 2 1 12 9 2 11 13 16 13 13 1 13 1 10 9 1 10 9 1 10 9 2 9 16 15 13 1 11 1 13 1 10 9 1 15 13 10 9 0 1 12 2
19 1 10 0 9 2 13 10 9 1 15 13 10 9 1 11 1 10 11 2
23 15 3 13 1 10 9 1 9 13 10 9 11 2 15 3 3 13 13 10 9 1 11 2
17 15 13 10 9 1 15 3 13 1 10 9 3 7 13 10 9 2
15 11 13 0 1 10 9 7 2 1 10 9 2 13 9 2
11 10 0 9 13 1 10 11 2 9 2 2
24 10 9 13 3 11 13 13 13 1 10 9 11 1 10 9 1 3 1 9 15 13 13 9 2
6 15 3 13 2 3 2
4 3 9 9 2
7 3 10 9 1 10 11 2
5 3 9 7 9 2
3 2 6 2
9 3 13 0 10 11 13 15 13 2
16 13 0 15 13 10 9 1 11 2 16 10 9 13 13 0 3
12 10 11 2 3 2 3 13 13 1 10 9 2
8 2 9 2 2 3 13 3 2
20 15 13 1 11 2 13 10 9 1 10 9 1 9 11 2 3 2 1 9 2
22 1 10 9 0 2 10 9 13 10 9 2 3 13 1 9 0 15 13 1 10 9 2
18 1 10 9 11 2 15 13 10 9 1 10 9 13 1 10 9 0 2
49 7 2 1 11 2 10 0 9 7 9 15 15 13 13 9 1 10 0 9 15 10 9 1 10 9 1 10 11 13 1 10 9 1 10 9 1 13 10 9 1 10 9 7 10 9 1 10 9 2
4 15 12 5 2
14 1 12 2 10 9 1 9 0 13 9 1 12 5 2
14 9 1 10 11 13 9 1 9 12 9 1 10 11 2
24 3 2 10 9 1 9 1 10 9 2 15 13 1 12 5 2 3 13 10 9 1 12 5 2
36 13 10 9 2 1 15 2 1 10 9 11 2 11 2 2 1 10 9 11 2 11 2 11 2 2 1 10 9 11 2 9 1 10 11 2 2
29 10 9 1 10 9 0 1 10 9 3 13 1 10 0 9 0 2 10 11 2 7 1 10 11 2 9 1 9 2
21 10 9 13 10 9 2 1 9 13 2 1 12 9 1 9 7 12 9 1 9 2
15 1 12 2 15 13 12 9 1 9 7 12 9 1 9 2
40 1 10 9 1 10 9 11 13 13 12 9 7 10 9 1 12 9 2 13 13 10 9 1 9 7 3 13 1 13 9 12 12 1 10 9 1 12 12 9 2
12 9 1 10 9 13 1 10 9 1 10 9 2
12 2 13 1 9 1 12 9 7 3 13 9 2
14 1 10 0 12 9 2 10 9 1 9 13 12 5 2
11 3 2 13 1 12 5 7 12 5 2 2
19 10 9 13 1 12 12 9 1 9 0 2 13 0 9 1 10 10 9 2
20 10 9 1 10 9 13 12 5 2 1 12 2 3 1 9 0 7 1 9 2
7 11 13 9 1 10 11 2
4 13 2 1 13
15 13 9 0 2 0 7 0 1 15 13 9 1 10 11 2
14 3 2 16 10 9 1 10 9 3 13 4 13 3 2
29 1 9 0 2 10 9 13 1 10 9 1 10 9 3 0 7 0 2 1 0 9 1 13 10 9 7 10 9 2
25 13 15 13 1 10 0 9 0 7 13 1 10 9 1 10 9 7 9 2 9 0 1 10 9 2
5 11 13 9 1 9
17 13 9 12 13 10 9 1 15 15 10 9 0 13 15 13 1 13
14 1 10 9 0 2 10 9 1 9 13 1 10 9 2
37 10 9 13 1 10 9 16 2 3 2 13 13 1 9 2 13 13 10 9 1 10 9 0 7 13 4 1 13 1 10 10 9 1 9 1 9 2
13 16 15 13 13 1 10 9 2 3 10 9 13 2
24 7 2 1 16 10 9 13 4 3 13 2 13 0 16 15 13 16 10 9 13 3 13 15 2
8 2 1 13 2 13 10 9 2
6 1 10 9 15 13 2
9 10 9 3 1 10 9 15 13 2
9 13 16 13 3 2 2 13 11 2
19 13 10 9 1 10 9 15 13 10 2 0 2 2 3 10 9 1 11 2
21 1 10 9 1 10 9 2 3 2 10 0 9 1 10 9 13 13 1 10 9 2
9 10 9 1 11 13 1 9 13 2
52 12 1 10 0 1 10 9 1 10 9 1 10 11 2 15 3 13 15 13 2 13 10 9 11 2 13 1 10 9 0 10 2 9 2 3 0 1 10 9 2 2 15 13 3 12 9 2 3 10 3 0 2
12 2 15 3 2 13 9 1 9 2 2 13 2
19 10 9 1 10 9 0 11 7 11 7 10 9 1 10 11 3 13 13 2
30 2 10 11 7 10 11 13 10 2 9 2 0 2 13 12 1 10 9 0 1 10 11 2 15 3 3 13 15 13 2
26 13 3 1 10 9 1 10 9 2 9 11 2 10 9 0 2 0 9 2 3 0 2 2 13 11 2
22 10 9 0 13 15 3 0 1 9 0 2 16 10 9 13 1 15 10 9 3 13 2
41 13 10 9 1 15 11 13 0 3 1 13 0 2 11 2 10 9 2 13 0 3 1 13 0 2 7 11 2 10 0 9 1 9 2 3 13 7 0 7 0 2
24 1 10 9 2 3 1 10 9 2 11 13 1 10 9 1 10 11 2 11 2 7 15 13 2
41 2 15 13 1 16 3 15 13 10 9 2 3 15 13 10 9 7 16 3 13 12 9 1 9 1 10 9 7 3 10 12 9 2 3 13 2 2 13 10 9 2
12 15 13 13 10 0 9 1 10 9 1 11 2
38 3 1 10 9 3 2 13 1 10 11 2 11 2 2 11 13 1 10 9 2 12 9 3 1 13 15 13 1 15 3 13 7 0 9 1 10 9 2
4 13 9 0 2
48 1 3 0 2 10 9 2 11 2 2 11 2 13 10 9 1 10 10 0 9 2 13 1 11 2 15 3 13 10 9 1 11 2 9 1 11 2 1 10 9 2 11 2 2 13 1 12 2
8 11 13 16 3 13 9 1 11
20 9 1 10 11 2 11 2 13 13 1 9 1 10 9 1 10 9 1 10 11
18 10 9 1 10 11 2 11 2 13 13 9 1 10 9 1 10 11 2
38 3 1 10 9 2 11 13 16 13 1 9 1 16 10 9 0 13 10 9 1 10 9 1 9 13 1 10 9 1 9 1 10 9 11 2 13 9 2
24 7 2 1 10 11 2 10 9 1 9 1 10 11 2 11 2 13 16 10 9 3 13 13 2
21 1 11 2 10 9 0 13 16 10 9 1 10 9 13 3 9 10 9 7 9 2
13 9 2 9 1 10 9 13 1 10 9 1 9 2
22 16 10 9 1 10 9 3 13 9 0 1 10 9 11 2 10 9 0 13 10 9 2
34 13 0 16 2 3 2 10 9 13 3 0 16 1 10 11 7 13 13 2 1 10 9 11 2 10 10 9 1 13 10 9 1 9 2
8 16 13 13 2 13 10 9 2
18 3 2 15 13 16 10 9 13 10 9 15 3 13 0 1 10 11 2
14 11 3 13 0 10 9 1 11 1 10 0 12 9 2
25 13 3 1 9 9 15 15 13 1 12 1 10 9 2 11 2 2 3 13 10 9 1 10 9 2
4 13 10 9 2
22 2 10 9 3 13 13 1 13 10 9 1 10 9 1 9 3 13 9 1 9 2 2
34 3 2 1 10 9 15 2 3 2 13 10 9 1 10 9 1 9 0 7 2 3 2 1 9 0 2 13 1 10 9 1 10 11 2
22 10 9 0 13 15 1 10 9 1 9 2 1 10 9 1 12 9 1 10 10 9 2
25 10 9 0 1 10 9 1 11 13 1 10 9 1 9 12 9 2 1 9 12 1 10 9 2 2
20 1 10 9 2 10 9 13 9 1 10 9 3 1 10 9 1 10 0 9 2
30 13 0 13 16 10 9 13 10 9 1 13 9 0 1 10 9 2 15 3 13 13 1 10 9 1 10 2 9 2 2
30 13 10 9 0 1 10 9 0 2 13 1 15 10 9 3 3 0 2 1 9 1 9 1 9 7 10 9 1 9 2
6 13 10 9 3 9 2
33 11 2 10 9 1 9 0 1 10 9 1 10 9 1 10 9 2 12 1 9 2 1 10 9 12 1 10 9 13 1 12 12 2
34 16 10 9 13 1 10 9 12 1 9 2 13 13 10 9 0 1 1 10 9 12 12 9 2 1 3 12 12 9 2 13 10 9 2
7 10 9 13 10 0 9 2
8 11 13 9 1 13 1 10 9
32 1 10 9 11 2 12 1 10 9 0 1 10 9 1 9 1 10 11 2 13 0 13 10 9 1 10 11 1 10 9 11 2
13 10 9 2 13 2 2 13 13 1 10 9 2 2
25 1 10 9 1 10 11 1 10 9 1 10 11 2 10 9 13 16 10 9 13 2 9 13 2 2
38 3 1 10 11 2 10 9 1 10 11 2 10 11 13 12 9 13 1 10 9 2 1 10 11 2 9 2 10 11 2 9 2 7 10 11 2 9 2
18 2 16 13 10 12 9 2 13 1 12 5 1 9 1 10 9 13 2
14 13 16 2 13 10 0 2 13 9 2 2 13 11 2
30 11 13 16 10 9 13 16 4 13 1 2 9 2 2 9 1 10 10 9 2 2 15 3 13 9 1 10 9 13 2
30 2 15 13 16 13 10 9 1 13 10 9 13 1 10 9 7 3 13 13 16 10 10 9 1 10 9 13 9 2 2
17 11 13 3 1 11 7 3 13 13 1 10 9 0 1 10 9 2
9 15 3 13 2 3 2 12 9 2
27 1 10 9 0 2 3 13 0 11 7 11 2 11 2 7 10 9 1 2 9 2 2 11 2 11 2 2
18 15 13 4 13 1 13 9 1 0 2 9 1 10 9 7 9 0 2
17 10 9 11 2 15 13 10 0 1 10 9 2 15 13 1 13 2
9 9 13 3 1 10 9 1 10 9
1 11
35 10 9 11 13 10 9 0 1 10 9 2 1 12 9 2 2 9 11 2 11 2 7 11 2 11 2 2 3 2 1 10 10 9 11 2
28 12 9 1 10 9 7 10 9 13 16 13 1 11 2 16 10 9 2 11 7 11 2 13 9 0 1 9 2
22 2 13 1 10 11 16 15 13 10 11 2 2 13 10 9 2 11 2 1 10 11 2
22 10 9 13 1 11 1 2 11 2 13 15 2 11 2 2 1 9 0 13 1 11 2
23 10 9 2 1 11 2 15 13 1 9 1 10 9 2 10 0 9 7 10 9 1 9 2
32 2 13 10 9 15 13 1 9 7 15 13 16 13 1 10 9 10 9 0 1 10 9 2 10 9 1 9 0 7 0 2 2
23 0 7 0 1 10 9 1 10 11 2 11 13 12 1 10 9 3 0 1 10 9 0 2
34 3 2 1 13 10 9 13 1 11 2 15 3 13 13 3 9 1 10 11 2 15 13 1 13 15 1 10 9 2 3 13 1 11 2
15 9 1 10 9 1 11 2 11 13 10 9 1 10 9 2
20 1 2 11 2 15 13 2 11 2 2 10 9 13 10 9 1 2 0 2 2
20 10 9 1 11 15 10 11 13 3 13 15 2 11 2 2 1 9 1 11 2
25 2 13 15 1 10 3 0 7 0 9 1 10 9 2 15 13 1 10 0 9 2 2 15 13 2
44 10 9 1 11 13 10 0 9 2 7 13 0 2 13 1 10 0 9 16 10 9 7 10 9 13 9 0 7 16 10 9 1 10 9 13 13 9 1 10 9 1 10 9 2
28 11 13 1 9 7 13 10 9 1 10 9 1 10 9 1 9 0 0 1 13 2 1 10 9 1 10 9 2
53 11 13 10 9 1 9 13 7 9 0 7 13 10 9 1 13 2 9 2 2 10 9 0 1 13 9 1 13 2 3 15 10 13 1 10 9 1 10 11 2 9 1 10 11 2 2 9 1 9 1 10 11 2
6 15 13 11 7 3 13
13 10 9 11 13 3 15 16 15 13 1 10 9 2
26 11 13 10 9 2 11 10 9 2 16 2 3 1 10 9 2 15 13 9 1 10 9 1 10 10 2
23 3 2 11 13 10 9 2 11 13 10 2 9 2 1 10 9 7 13 15 9 7 9 2
20 3 13 1 11 10 9 1 10 9 2 1 16 15 15 13 3 1 10 9 2
29 10 9 0 13 15 1 2 11 2 2 12 2 2 15 13 2 0 2 7 11 13 16 15 15 13 10 9 0 2
17 11 13 10 9 2 0 7 0 2 11 13 3 0 7 3 13 2
21 11 13 0 1 13 2 11 13 0 7 2 3 2 13 9 1 10 9 2 13 3
15 11 13 0 3 2 11 13 2 0 2 2 1 9 0 2
17 10 9 1 10 11 3 9 3 13 13 1 15 1 9 3 9 2
27 15 12 13 0 3 1 10 9 3 0 2 0 7 0 2 3 1 15 3 2 0 2 2 0 7 0 2
22 1 10 9 1 10 9 2 10 9 13 13 1 10 9 2 1 0 9 7 1 9 2
15 10 9 13 1 10 9 11 2 9 1 10 9 1 11 2
17 10 9 2 13 16 13 1 9 12 12 2 13 15 10 9 13 2
8 10 9 13 2 7 15 13 2
11 2 6 2 2 13 10 9 1 10 9 2
20 13 1 12 9 2 10 9 13 12 9 15 13 13 10 10 9 1 10 9 2
12 13 3 0 7 13 3 9 1 13 9 0 2
36 10 9 13 0 7 0 7 10 10 9 13 13 1 9 2 9 7 9 2 13 1 10 0 9 2 9 2 2 2 9 2 7 2 9 2 2
20 1 9 1 11 2 10 11 13 10 9 1 10 11 7 10 9 1 10 9 2
24 10 0 13 13 1 10 9 1 10 11 7 1 10 9 10 9 3 1 10 9 1 10 11 2
15 10 3 0 2 3 2 13 10 9 15 10 9 13 13 2
15 1 15 13 1 10 9 1 10 9 1 10 15 13 13 2
36 13 3 16 2 3 10 9 0 15 13 1 10 9 1 9 1 10 9 0 0 15 13 10 11 2 13 12 9 2 13 10 9 1 10 11 2
62 3 2 16 10 9 3 13 0 7 13 3 10 9 1 10 9 0 2 15 13 3 13 1 10 9 0 7 0 1 10 9 1 9 1 3 13 10 9 2 15 3 13 13 1 16 13 7 3 13 10 9 7 16 13 10 9 1 10 9 7 9 2
31 16 13 1 10 11 10 9 1 9 1 10 9 11 2 10 0 9 13 10 9 1 10 9 1 10 9 15 13 10 11 2
40 1 10 9 1 10 9 1 11 2 11 2 10 9 15 13 1 10 9 0 2 16 10 9 13 13 1 10 9 1 10 9 1 10 11 1 10 11 2 11 2
11 15 3 13 10 9 0 13 1 10 9 2
5 10 9 1 10 9
2 3 13
25 3 13 2 10 9 1 10 9 13 10 9 0 7 15 1 10 9 2 10 9 1 10 9 0 2
26 9 13 1 10 9 12 7 12 3 1 10 9 11 2 11 2 11 2 11 2 11 2 11 7 11 2
14 13 2 9 13 1 9 13 1 9 1 10 10 9 2
9 11 2 10 9 9 13 10 9 2
23 3 10 9 15 13 13 2 13 10 9 1 13 9 0 7 10 9 3 13 13 9 0 2
14 7 10 9 1 10 9 13 10 9 1 9 2 3 2
7 11 2 6 1 10 9 2
5 9 0 7 9 0
72 10 9 13 1 10 11 2 1 12 2 1 15 10 9 13 11 13 13 10 9 1 10 9 9 2 9 0 13 10 10 9 7 1 10 10 9 0 2 3 13 13 1 10 9 0 2 0 1 10 11 1 12 2 3 1 10 9 0 1 9 2 13 10 9 1 10 9 1 10 9 0 2
41 3 2 10 9 1 10 9 13 16 10 9 0 1 9 13 3 13 1 10 9 1 9 0 2 9 11 2 1 2 11 2 2 9 11 2 12 2 9 12 2 2
4 3 13 0 2
13 3 12 13 0 13 13 1 10 11 1 10 9 2
25 10 9 11 2 11 2 13 9 1 9 0 1 10 9 2 15 13 1 9 7 9 1 12 9 2
57 10 10 9 15 13 1 10 9 1 10 9 0 13 1 10 9 1 9 0 2 10 9 0 1 10 9 1 9 1 12 7 12 9 13 1 10 9 13 9 12 9 1 10 10 0 9 7 13 10 9 1 13 10 9 12 9 2
42 10 9 13 13 0 10 9 1 10 9 2 10 11 13 9 1 9 1 9 13 9 7 9 15 13 13 1 10 9 0 2 13 10 0 9 1 10 2 9 2 0 2
12 11 13 9 2 9 7 9 1 10 9 11 2
18 11 13 9 12 12 1 13 9 1 10 9 7 13 10 9 1 11 2
3 2 6 2
8 3 13 1 11 1 9 10 2
8 13 3 1 9 2 2 13 2
17 15 13 1 10 9 1 12 9 1 11 13 1 13 9 1 11 2
15 2 13 0 10 9 13 15 1 13 10 9 2 2 13 2
12 10 9 13 15 1 10 9 7 3 15 13 2
25 10 9 2 2 16 10 11 13 10 9 1 3 13 13 10 11 1 10 0 9 2 9 2 2 2
13 10 11 2 3 13 1 9 2 2 1 10 9 2
15 2 15 13 10 9 1 10 9 2 13 13 10 9 2 2
29 10 9 1 10 9 2 15 13 1 10 9 1 10 9 2 13 9 1 9 1 10 9 1 10 9 1 12 9 2
15 13 1 13 10 9 13 7 10 9 13 15 1 10 9 2
25 13 13 1 13 10 9 2 3 2 13 13 2 9 2 2 9 1 9 1 9 2 1 10 9 2
31 1 10 9 2 13 10 9 1 10 9 0 1 10 0 9 1 9 7 13 10 9 0 1 10 9 13 13 10 9 0 2
30 2 13 0 13 3 16 10 9 1 10 9 1 10 9 1 10 9 13 13 1 12 5 1 10 9 1 10 9 0 2
14 10 0 13 3 0 16 13 9 12 9 2 2 13 2
25 11 13 3 16 10 9 1 9 13 1 10 9 1 10 9 15 15 13 1 10 10 9 1 9 2
33 9 2 13 1 10 0 9 12 2 1 10 11 2 11 2 12 2 2 9 1 10 9 1 10 9 1 9 1 10 9 1 11 2
16 10 9 13 4 13 1 10 0 9 12 2 1 10 9 12 2
25 9 1 9 2 10 11 13 12 9 1 10 9 2 11 2 2 15 13 1 12 1 12 1 9 2
6 9 1 10 9 12 2
13 10 9 3 13 10 9 1 10 9 0 1 9 2
7 9 13 10 9 13 1 11
18 10 12 11 1 2 11 2 13 10 9 1 10 9 1 10 9 1 12
5 11 13 10 9 2
10 2 11 13 3 13 1 10 9 2 2
18 10 9 1 12 2 9 11 2 13 3 10 0 9 13 1 10 9 2
32 10 9 13 10 9 0 1 10 9 1 10 9 1 12 2 3 3 1 10 9 1 10 9 0 2 1 12 1 9 1 12 2
31 15 13 10 9 1 15 11 13 1 13 10 9 1 10 9 1 13 15 10 9 0 1 10 9 15 13 1 11 7 9 2
25 1 10 9 2 10 9 13 15 1 10 0 9 3 2 1 13 1 10 0 9 2 2 11 2 2
12 3 1 10 9 11 13 1 10 9 0 11 2
28 10 9 3 13 0 1 10 9 7 1 10 9 1 10 9 3 1 10 12 9 1 15 13 13 1 10 9 2
18 7 3 3 1 15 3 3 15 13 13 2 13 9 1 10 0 9 2
61 1 13 10 9 1 9 2 13 15 13 10 10 9 1 9 2 9 0 7 11 10 11 1 10 11 13 10 9 1 13 1 10 9 0 9 1 10 9 7 1 10 9 1 10 9 2 15 2 13 2 13 4 13 3 3 10 11 7 10 9 2
64 7 10 9 13 3 10 9 1 10 2 9 2 2 10 9 0 2 10 0 9 2 13 10 0 9 1 9 7 9 1 10 9 0 2 0 1 13 13 1 9 3 0 1 9 7 9 7 2 3 13 10 9 2 13 3 16 2 3 15 13 13 3 2 2
36 11 9 10 13 9 3 11 13 10 9 1 9 1 9 1 10 11 15 13 10 9 0 3 15 13 2 13 15 10 9 0 1 13 10 9 2
14 2 15 13 9 1 10 11 15 13 9 1 10 9 2
21 16 11 2 10 9 2 9 7 9 13 15 13 3 13 16 13 13 10 9 0 2
6 3 15 15 13 15 2
9 7 2 15 3 2 2 13 11 2
46 1 10 9 2 3 1 13 1 10 9 1 11 2 11 2 2 3 13 13 10 9 1 10 9 1 3 2 11 13 16 13 13 10 9 1 10 9 11 2 11 2 1 10 9 0 2
12 11 2 3 15 13 10 9 1 15 13 13 2
4 11 2 3 2
16 9 13 15 2 13 15 13 0 2 3 13 10 9 1 9 2
7 10 0 9 3 13 13 2
3 10 9 12
25 2 9 0 1 9 1 11 2 12 9 1 11 2 13 13 3 1 10 11 2 11 2 1 11 2
9 10 9 13 10 9 1 10 9 2
9 10 9 1 11 13 12 9 13 2
6 11 13 12 9 0 2
8 9 0 1 10 11 13 1 9
20 10 9 0 1 11 13 1 9 3 2 1 9 1 10 9 13 1 10 11 2
21 10 9 13 1 9 0 1 10 11 1 10 11 2 15 13 10 9 1 12 5 2
11 1 11 2 10 9 13 13 1 13 3 2
6 15 13 9 1 11 2
6 11 13 10 3 0 2
15 13 2 13 12 9 7 13 1 10 9 1 10 0 9 2
16 2 15 13 3 1 15 2 6 2 2 2 13 11 1 11 2
13 10 9 13 13 9 1 10 9 1 9 12 12 2
11 10 9 1 9 12 12 13 9 1 9 2
17 16 10 9 1 10 9 13 0 2 13 0 13 9 1 9 0 2
11 1 10 9 0 10 9 13 1 9 12 2
26 16 3 13 15 13 1 10 9 0 2 13 9 2 3 10 11 2 9 12 2 15 13 9 1 9 2
34 1 11 2 9 1 9 1 10 11 2 10 9 2 13 1 10 9 1 12 9 2 13 1 10 9 0 1 10 9 13 1 10 9 2
19 10 9 1 9 1 10 11 13 13 1 10 9 15 13 3 1 10 9 2
28 11 2 10 9 13 12 9 13 1 9 0 1 9 1 9 7 12 9 1 9 2 15 13 9 0 7 9 2
19 1 9 1 9 1 10 9 1 10 9 7 9 1 10 9 1 10 9 2
12 9 1 10 9 2 1 9 12 1 9 12 2
5 1 12 1 9 2
6 9 13 12 9 1 9
39 10 0 9 1 9 1 10 11 13 1 10 0 9 1 9 12 9 1 9 2 9 2 7 13 1 12 5 1 12 5 3 0 16 10 1 10 9 0 2
12 10 11 11 7 11 13 10 9 12 7 12 2
19 13 9 1 12 9 1 9 2 9 2 2 15 13 13 9 1 10 9 2
7 11 15 13 9 1 10 11
28 10 9 7 9 1 9 2 11 2 13 13 1 10 0 9 9 1 10 11 1 10 9 1 11 2 11 2 2
12 13 10 10 0 9 1 10 9 1 10 9 2
18 3 11 13 0 1 10 9 3 9 2 10 9 11 13 7 13 6 2
17 13 1 13 1 10 9 2 11 13 1 13 4 13 3 1 10 9
3 9 2 9
1 9
23 3 1 10 11 2 10 9 13 10 9 15 15 13 1 9 1 9 7 1 9 1 9 2
60 10 9 1 9 7 10 9 1 10 9 0 13 1 9 9 1 10 11 1 10 9 1 10 9 12 2 3 2 1 10 9 3 13 2 10 9 13 4 13 1 10 9 13 1 10 9 11 2 1 13 7 13 10 9 1 10 0 9 0 2
13 3 13 3 9 1 10 9 1 10 11 1 3 2
54 10 0 9 1 12 9 13 10 9 1 10 11 13 4 13 3 0 7 1 9 15 13 2 13 7 13 1 10 9 1 10 10 10 9 2 7 13 3 15 12 1 10 9 1 10 9 1 10 9 13 1 10 9 2
24 3 1 10 11 2 3 2 10 9 1 10 11 0 13 16 13 12 9 1 10 0 12 9 2
23 13 1 9 1 10 9 7 1 10 9 2 10 9 13 9 1 12 9 1 13 10 9 2
10 10 9 13 13 10 9 1 10 9 2
25 1 10 9 1 10 9 2 11 2 10 9 13 4 13 3 1 10 9 1 9 7 9 1 9 2
5 9 13 1 9 13
28 1 10 9 12 1 9 1 12 2 9 0 3 13 10 9 0 1 10 11 2 13 1 11 2 1 10 11 2
31 10 11 2 3 1 10 0 9 1 10 9 2 11 2 13 1 9 1 10 11 7 10 9 1 10 9 2 11 7 11 2
20 10 0 2 9 0 2 2 15 3 13 3 10 11 2 13 15 1 10 9 2
4 7 10 11 2
25 1 10 11 2 1 11 2 13 15 1 11 2 9 1 10 9 1 10 9 0 1 10 9 0 2
17 11 2 1 10 9 2 13 13 3 2 7 13 15 1 10 9 2
13 10 11 2 3 2 13 3 3 0 16 10 11 2
10 11 13 13 3 10 9 1 9 0 2
5 3 13 10 0 2
10 7 15 13 1 11 7 13 10 9 2
21 3 13 13 1 10 0 9 1 10 9 0 1 10 9 1 9 7 9 1 9 2
22 3 13 13 1 10 9 1 10 9 1 13 10 9 1 10 9 0 1 10 9 0 2
11 7 13 0 9 1 10 9 1 10 9 2
38 10 9 3 13 13 1 10 9 13 1 10 11 2 15 13 13 0 1 13 9 13 1 9 7 13 9 0 1 9 15 13 9 1 9 1 10 9 2
32 9 13 1 9 15 13 9 1 10 9 1 12 7 12 13 16 12 9 13 4 13 1 9 1 9 13 1 10 9 1 9 2
3 1 10 9
41 3 9 13 1 10 11 2 10 9 1 10 9 1 10 9 1 10 2 11 2 1 9 12 9 13 16 4 13 10 9 2 1 12 9 0 2 13 7 1 9 2
13 13 1 12 9 7 9 10 9 0 1 10 9 2
2 9 0
13 10 11 13 9 12 9 1 9 1 10 9 0 2
27 1 10 9 11 2 10 9 13 10 9 1 9 15 15 13 3 9 1 10 9 0 2 1 10 11 2 2
21 1 10 9 2 15 13 13 10 9 2 1 10 9 1 9 2 1 13 12 9 2
6 9 13 1 12 5 0
23 10 9 1 9 13 1 10 9 2 1 10 9 2 9 0 1 12 5 2 1 10 11 2
20 10 9 0 2 1 9 1 0 1 9 2 13 13 1 10 9 1 10 11 2
21 3 2 10 9 13 9 1 12 5 2 1 10 15 10 9 1 9 13 12 5 2
6 9 1 10 11 13 13
22 10 9 15 15 13 3 1 10 11 2 1 11 2 13 13 1 10 9 1 10 9 2
28 2 3 13 0 1 13 13 1 10 9 2 2 13 11 2 12 2 15 13 10 9 1 10 9 11 2 12 2
11 15 13 10 9 1 10 11 1 10 9 2
3 9 13 9
48 10 9 11 2 13 1 10 9 1 10 11 2 11 2 1 13 10 9 1 9 1 10 9 2 13 3 16 2 16 13 2 13 13 9 1 10 9 1 13 9 7 13 9 0 1 10 9 2
24 1 10 9 1 3 2 10 9 13 13 10 9 1 10 9 1 13 16 13 7 3 10 9 2
20 1 10 9 11 2 2 11 2 13 3 12 1 10 0 9 1 10 9 0 2
19 13 9 1 10 11 2 9 1 10 11 2 9 0 1 9 1 10 11 2
22 13 10 9 0 1 10 9 1 10 9 1 10 9 2 10 2 11 2 2 11 2 12
4 9 3 13 9
15 9 13 10 9 0 3 1 15 13 10 9 0 1 9 2
13 10 10 9 1 10 9 13 0 2 9 7 9 2
22 10 9 13 10 0 9 0 13 13 1 10 9 0 1 9 7 9 1 9 1 9 2
13 2 10 9 1 10 9 13 10 9 1 10 9 2
8 15 13 13 2 2 13 11 2
17 1 15 2 10 9 13 1 10 9 1 9 0 1 9 1 9 2
19 13 16 10 9 13 13 2 1 9 1 9 0 1 9 1 9 0 2 2
19 10 9 1 10 9 13 4 13 3 1 10 9 1 10 9 1 10 11 2
21 7 15 2 1 10 11 2 1 13 2 9 2 2 1 2 10 9 1 3 2 2
4 9 1 10 9
19 11 13 1 10 9 7 1 10 9 13 16 3 13 15 1 10 10 9 2
13 7 16 2 3 2 3 13 1 10 9 1 11 2
18 10 9 3 13 1 15 1 11 2 1 10 9 1 10 9 1 11 2
24 2 3 13 10 9 0 2 7 15 13 15 1 13 10 9 1 9 1 10 9 2 2 13 2
13 1 15 2 10 9 13 13 2 1 15 15 13 2
15 11 3 13 13 16 10 9 1 10 9 13 13 10 9 2
8 9 13 9 1 9 1 10 9
23 10 11 3 13 3 10 9 13 2 11 2 1 9 1 9 13 1 10 11 2 1 11 2
26 1 9 7 9 2 9 1 15 10 2 9 2 13 13 1 10 9 2 10 9 13 10 9 1 9 2
16 3 2 13 1 10 9 1 10 9 1 10 9 1 12 9 2
22 10 9 3 15 13 1 9 0 1 13 1 10 0 9 0 0 1 9 7 9 0 2
31 7 13 10 9 0 1 9 13 1 9 1 9 0 2 9 1 11 7 9 1 9 1 12 9 15 13 3 9 12 9 2
8 2 9 2 13 9 1 10 11
34 9 1 9 1 11 2 11 2 13 16 13 9 0 1 13 9 1 10 9 15 13 9 0 1 10 9 2 16 10 9 15 13 13 2
11 11 13 10 9 0 1 10 11 7 11 2
32 10 9 13 16 13 13 3 10 9 0 2 1 15 11 2 1 10 11 2 11 2 1 10 11 2 7 11 2 1 10 11 2
30 10 9 13 1 10 2 9 2 2 9 7 9 1 10 0 11 2 9 1 10 11 2 10 9 13 1 10 0 9 2
13 11 13 13 10 11 1 10 9 7 1 10 9 2
5 3 2 3 13 2
11 1 15 2 13 11 2 9 1 10 9 2
14 11 13 10 9 1 13 9 1 10 9 1 10 9 2
28 1 13 10 9 1 10 10 9 2 15 13 10 10 9 1 12 9 0 2 1 10 9 1 11 7 1 11 2
11 15 1 15 13 0 2 0 2 1 9 2
22 1 10 9 2 1 10 9 2 1 10 9 13 10 9 1 13 2 3 1 3 13 2
47 11 2 9 1 10 9 2 3 13 15 10 10 9 15 13 2 7 13 12 9 1 10 9 1 10 10 12 9 1 2 3 2 13 10 9 0 7 10 9 0 1 10 9 1 10 9 2
15 1 10 9 1 10 9 13 13 12 9 1 9 7 9 2
14 10 9 1 9 13 1 13 12 9 0 1 10 11 2
14 7 10 9 1 9 13 1 13 12 12 9 1 9 2
43 10 9 13 13 1 11 2 0 1 10 9 1 10 9 1 10 0 9 1 10 11 2 11 2 2 1 10 0 9 1 10 11 7 1 10 9 11 1 10 9 0 11 2
30 1 10 9 2 11 13 10 12 0 9 1 10 9 1 11 2 15 13 1 4 13 1 9 0 13 1 10 9 11 2
14 15 13 10 9 1 10 0 2 13 1 13 10 9 2
16 3 13 3 2 7 13 16 3 13 13 10 0 9 1 11 2
9 10 9 13 3 13 10 9 0 2
15 2 3 2 13 3 10 9 7 15 15 12 9 1 9 2
23 7 15 15 13 13 3 1 9 1 10 9 2 15 13 9 2 9 7 9 3 13 13 2
7 3 13 0 2 2 13 2
10 3 2 1 10 9 1 10 9 0 2
14 10 9 13 9 0 2 7 3 13 13 1 10 9 2
2 11 12
23 10 11 2 9 13 1 10 9 1 11 2 13 13 10 9 1 10 9 1 9 1 9 2
15 9 1 12 1 12 9 13 13 1 13 9 1 9 0 2
2 11 12
32 10 11 1 10 11 13 16 11 13 1 10 12 9 0 15 13 12 5 1 9 0 1 10 0 9 1 9 2 13 1 12 2
13 1 10 9 2 10 9 13 13 3 12 12 9 2
6 11 13 9 1 10 11
13 11 13 16 9 1 9 0 13 10 11 1 13 9
15 10 11 13 9 1 10 11 1 10 9 0 1 10 11 2
23 10 9 13 10 9 15 13 1 10 9 1 10 11 16 13 9 1 10 9 0 1 11 2
7 10 9 13 3 1 11 2
33 2 16 10 9 1 10 9 13 13 1 10 9 1 10 9 2 10 9 13 1 12 5 1 12 5 1 10 9 2 2 13 11 2
18 10 9 1 10 9 2 1 15 2 13 12 5 1 10 9 1 9 2
12 10 9 3 13 10 9 0 13 1 10 9 2
15 9 0 2 9 12 12 2 1 10 9 2 9 12 12 2
22 3 1 10 0 2 10 9 0 13 1 10 11 15 13 9 9 12 2 1 10 11 2
7 9 13 9 0 1 10 9
11 11 13 10 9 3 13 1 10 9 0 2
44 3 2 10 9 1 10 9 13 1 10 9 15 1 10 9 1 10 9 2 7 11 13 3 1 10 9 0 1 10 11 1 10 9 7 1 10 9 1 2 0 2 3 9 2
19 10 9 1 11 13 1 13 1 10 9 15 3 13 0 1 10 9 0 2
32 1 10 9 7 9 1 10 9 2 10 9 13 3 1 10 0 2 3 16 13 1 10 10 9 0 2 10 10 9 1 9 2
6 13 10 9 1 10 9
16 9 1 9 15 13 2 3 2 10 9 7 10 9 1 10 11
29 10 9 2 1 10 9 13 1 10 9 1 10 9 2 11 2 7 10 9 1 10 11 2 1 10 9 2 11 2
28 13 13 9 0 1 10 9 7 1 10 9 13 1 10 9 1 10 9 2 1 10 9 7 1 10 9 0 2
10 9 0 1 10 9 0 13 12 5 2
25 10 9 0 1 10 9 1 9 3 0 1 10 9 1 11 13 1 9 12 5 2 1 10 11 2
15 10 9 13 3 0 16 10 13 1 9 2 12 5 2 2
11 10 0 9 13 1 10 9 1 10 11 2
13 11 1 11 13 9 1 12 1 10 9 1 10 11
30 10 11 13 3 1 11 11 2 10 2 11 2 2 9 1 12 1 10 9 1 10 11 2 9 0 15 13 9 2 2
29 2 11 2 13 13 1 10 9 1 10 11 2 1 10 9 2 3 13 13 12 9 1 9 1 11 2 11 2 2
21 11 1 11 2 15 3 13 13 1 10 11 1 12 9 1 9 2 1 10 11 2
19 10 9 1 11 1 10 9 1 10 9 13 13 1 10 0 1 10 9 2
27 9 13 1 10 9 1 10 9 1 10 9 13 2 1 10 9 0 2 1 10 9 1 10 9 13 9 2
34 3 16 15 2 10 9 1 10 9 13 16 2 1 10 9 0 2 3 15 13 13 3 10 9 1 10 9 13 9 1 10 9 0 2
27 1 9 1 11 2 9 1 10 9 2 10 9 1 10 11 2 11 2 13 10 9 1 11 1 10 9 2
12 2 10 9 1 10 9 13 0 2 2 13 2
17 13 1 10 9 1 10 9 2 11 13 10 9 7 13 10 9 2
8 11 13 10 9 1 10 9 2
14 13 1 10 9 1 9 2 13 10 9 1 10 9 2
22 10 11 3 13 1 13 9 1 9 0 1 10 11 2 11 7 11 2 1 12 9 2
25 10 0 9 1 9 2 13 1 11 2 13 1 10 9 1 9 7 10 9 1 9 1 0 9 2
7 2 13 10 9 0 2 2
24 1 11 2 10 0 9 7 9 13 12 5 1 10 9 2 15 13 1 9 12 9 1 12 2
13 2 1 10 0 9 13 15 12 5 2 2 13 2
6 11 2 13 16 3 2
14 10 10 9 13 13 1 10 9 0 1 10 9 0 2
44 2 11 2 2 12 1 10 9 0 1 10 9 2 13 10 10 9 1 10 9 1 13 7 13 10 9 1 10 9 15 13 10 9 1 10 9 1 10 9 1 10 9 0 2
7 10 9 1 9 13 0 2
17 12 1 10 9 15 10 9 3 13 13 13 10 9 1 10 9 2
6 11 13 1 10 9 2
15 11 13 10 9 1 9 7 9 1 13 10 9 1 9 2
12 3 15 13 16 10 9 0 13 1 10 11 2
20 10 9 13 10 9 0 2 15 3 15 13 13 1 10 9 1 9 1 11 2
49 9 0 7 0 3 10 9 0 1 10 9 1 9 13 1 9 0 1 10 9 0 1 10 11 2 1 10 9 1 16 13 10 9 1 10 9 2 3 3 16 10 9 15 13 1 13 10 9 2
37 3 13 1 11 2 9 1 10 9 3 13 2 7 1 11 10 9 2 1 10 9 0 1 10 9 2 9 13 2 13 10 0 9 1 10 9 2
25 10 9 13 13 10 9 1 10 9 2 13 1 10 11 7 1 10 9 7 13 1 10 9 11 2
13 11 2 12 2 13 13 1 9 0 1 10 11 2
17 2 10 9 13 1 13 15 13 1 2 9 9 2 1 10 9 2
22 9 13 16 3 10 9 13 10 9 15 13 10 9 1 3 12 9 2 2 13 11 2
10 10 9 13 4 13 1 9 1 9 2
18 13 2 13 2 1 10 9 1 10 9 2 3 1 10 9 1 9 2
10 10 9 1 10 9 3 3 13 13 2
60 11 13 12 9 1 10 9 2 10 9 1 10 11 7 10 9 1 10 10 9 0 2 1 9 1 12 3 1 12 9 2 2 10 9 1 2 10 9 0 2 2 1 12 1 12 9 2 7 10 9 1 10 9 1 10 9 1 10 11 2
26 10 9 11 13 1 0 9 1 10 9 1 3 1 9 1 10 9 0 7 1 9 0 1 10 11 2
9 11 13 9 1 9 7 11 13 9
11 9 0 13 2 9 2 1 9 1 10 9
11 11 7 11 13 0 9 0 1 10 9 2
14 10 9 7 9 11 13 1 10 9 10 9 1 13 2
27 3 10 9 1 10 9 7 10 9 1 10 9 3 13 13 12 9 1 9 1 10 11 2 11 7 11 2
2 9 0
24 10 9 1 10 9 11 7 11 2 9 0 1 11 2 13 1 10 9 12 1 9 1 12 2
35 10 9 11 2 1 10 9 1 12 9 2 2 3 1 13 1 10 9 2 13 1 10 9 2 13 1 10 9 2 13 10 9 7 13 2
19 10 11 2 9 0 1 3 12 9 1 9 2 13 10 9 3 1 11 2
46 10 9 2 0 1 10 9 1 12 2 3 13 10 9 1 10 9 1 10 9 1 10 11 2 9 1 12 2 2 1 10 11 2 9 1 12 2 7 1 11 2 9 1 12 2 2
11 10 9 0 1 10 9 3 13 13 9 2
27 11 13 16 3 10 9 7 9 0 11 13 9 1 13 1 10 9 1 11 2 1 10 9 2 1 11 2
15 2 10 9 1 9 13 13 13 10 9 2 2 13 11 2
9 10 9 13 10 9 1 10 9 2
12 2 10 9 1 9 0 13 0 2 2 13 2
5 2 1 11 3 2
14 10 9 1 3 13 3 13 1 9 1 10 9 12 2
11 16 13 13 0 16 13 16 13 0 2 2
19 1 15 13 3 0 13 10 9 0 1 10 9 15 13 1 10 9 0 2
14 3 2 13 15 15 13 13 1 10 9 1 15 13 2
12 15 13 3 13 10 9 2 15 13 3 13 2
15 10 9 2 10 9 3 10 9 13 13 2 3 13 0 2
2 15 13
7 0 9 1 3 12 9 2
11 13 10 9 2 15 13 15 1 15 1 9
18 0 16 10 9 13 16 13 10 10 9 1 13 10 9 1 10 9 2
15 10 9 2 13 7 13 13 2 2 10 0 1 10 9 2
35 10 2 9 2 0 15 13 10 9 3 7 13 10 9 3 7 15 13 13 10 9 2 13 15 13 3 10 9 13 1 10 9 9 0 2
20 13 16 3 15 13 10 0 9 0 1 10 9 15 13 15 13 1 13 13 2
26 7 10 9 3 13 15 13 1 10 9 7 10 9 1 15 13 0 1 13 10 9 1 10 10 9 2
31 10 9 1 9 0 13 15 13 1 10 9 1 9 7 10 9 0 1 10 0 9 1 10 9 13 13 7 13 1 3 2
11 10 9 13 10 9 2 3 10 9 0 2
28 10 9 1 10 9 13 1 10 9 1 10 10 9 1 10 9 7 3 1 10 9 0 15 13 1 10 9 2
33 1 9 2 13 11 7 11 2 1 10 11 2 1 13 1 13 10 9 13 1 10 9 1 9 0 13 1 10 9 1 12 9 2
25 1 9 2 13 10 11 1 10 9 1 12 9 1 10 9 1 9 13 13 1 9 13 10 9 2
23 1 10 9 1 3 2 10 9 13 13 1 9 1 9 1 10 11 2 15 13 1 9 2
22 1 10 9 2 15 13 10 9 1 10 9 13 13 1 12 1 10 9 1 12 9 2
17 10 9 13 13 1 10 9 1 10 9 1 11 2 9 0 2 2
17 1 9 1 9 7 9 2 10 9 1 10 11 13 10 12 9 2
4 3 13 9 2
16 3 1 10 9 2 10 9 13 10 9 3 1 10 9 0 2
15 1 12 2 12 9 1 10 11 13 13 1 10 9 1 11
18 11 2 3 15 13 13 10 9 15 13 9 0 3 15 1 10 9 2
28 10 9 3 13 13 13 10 9 0 1 10 9 13 1 10 9 1 13 7 1 13 1 10 9 1 10 9 2
13 10 9 3 0 7 0 13 15 1 11 7 11 2
32 10 10 9 13 1 9 0 2 13 10 9 1 13 12 1 10 0 9 1 10 10 9 2 15 13 10 1 10 9 1 9 2
19 11 2 10 9 13 13 1 10 9 15 10 9 13 13 1 10 9 0 2
15 13 13 9 0 2 13 0 9 2 7 16 3 13 9 2
26 15 13 1 10 9 15 10 9 13 1 13 10 10 9 1 10 9 2 1 10 9 7 1 10 9 2
14 3 13 16 10 9 13 0 1 10 0 9 15 13 2
14 10 10 12 9 3 13 10 9 12 12 9 1 9 2
7 9 2 9 12 1 9 2
7 1 10 9 2 9 12 2
23 3 3 13 16 10 11 13 10 9 1 10 9 1 15 7 13 1 10 9 1 10 9 2
16 15 13 10 9 1 10 11 2 0 1 10 9 1 10 9 2
46 3 13 10 9 2 7 0 10 9 1 15 10 9 0 13 1 10 9 10 9 1 9 0 2 13 10 9 2 13 9 1 10 9 15 15 13 1 9 2 7 9 1 13 10 9 2
8 11 13 10 0 9 1 10 11
26 10 9 13 10 9 3 1 9 1 11 2 13 1 10 9 1 10 11 2 12 1 12 2 2 3 2
16 2 10 9 13 3 1 10 11 16 15 13 1 10 3 0 2
13 3 2 15 13 9 1 10 9 1 13 9 2 2
13 0 2 1 10 9 0 7 9 1 10 9 0 2
10 0 2 1 10 9 7 9 1 9 2
32 1 15 13 1 9 0 13 10 9 1 9 13 11 2 12 9 2 9 7 9 1 10 11 7 11 2 9 1 10 9 11 2
26 10 12 9 13 9 1 10 9 1 10 0 9 13 1 10 11 1 10 9 1 10 9 2 1 9 2
17 10 9 1 11 13 13 1 10 9 1 10 9 2 1 10 11 2
17 10 9 13 13 9 12 9 2 1 9 12 9 2 1 13 15 2
26 13 2 10 9 13 3 13 10 11 2 1 9 7 9 2 1 10 11 2 16 10 9 3 13 13 2
26 10 0 9 1 11 13 1 10 9 7 9 1 10 9 7 13 9 1 10 9 0 1 10 9 12 2
16 10 9 13 11 2 11 2 11 2 11 7 10 12 0 9 2
6 10 9 13 10 9 2
4 3 15 13 2
15 13 10 9 13 1 9 2 9 1 9 0 7 10 9 2
10 1 10 9 2 13 9 0 7 0 2
17 1 10 9 0 2 3 2 13 15 3 1 3 15 7 15 13 2
4 13 13 3 2
8 3 15 13 3 3 11 13 2
8 10 9 3 13 9 1 9 2
13 3 15 13 10 9 3 13 13 1 10 9 13 2
23 10 9 13 10 9 1 12 9 15 13 13 1 10 9 1 10 9 1 10 11 1 11 2
14 1 10 9 1 10 9 2 11 2 15 12 13 13 2
15 10 9 11 2 11 2 13 13 1 13 1 11 10 9 2
20 11 3 13 1 11 16 13 0 2 7 13 1 13 10 9 1 10 11 0 2
12 11 13 1 10 9 1 11 2 1 10 9 2
10 10 9 1 11 13 13 1 10 9 2
7 10 9 13 1 10 9 2
12 11 13 13 3 1 9 1 10 9 1 11 2
23 10 9 13 1 9 2 1 11 2 3 1 13 1 9 1 10 11 7 13 9 1 9 2
6 10 12 9 13 13 2
8 11 2 6 2 13 1 12 2
13 11 2 15 10 9 13 13 1 15 1 9 0 2
3 11 13 9
3 2 9 2
2 13 2
25 3 2 3 13 16 3 15 13 10 9 0 2 7 13 1 13 13 0 13 15 3 10 0 9 2
15 1 10 9 0 2 13 3 1 13 10 9 2 9 2 2
12 7 2 1 10 9 0 2 13 11 7 11 2
21 10 9 1 9 2 13 1 10 0 9 0 2 13 15 7 15 9 1 10 9 2
26 7 10 0 9 1 10 9 1 9 1 9 1 9 13 13 10 0 9 15 11 13 1 10 9 13 2
13 10 9 1 10 9 2 11 2 3 13 9 13 2
17 11 13 13 15 1 10 11 2 7 10 11 2 11 2 3 13 2
32 10 9 13 2 3 2 9 0 1 10 11 2 11 2 7 3 13 1 11 16 15 13 1 13 11 1 10 9 1 10 9 2
35 10 9 13 9 1 10 9 2 11 2 2 13 1 10 11 2 11 2 2 1 10 11 2 1 10 11 2 11 2 2 9 1 10 9 2
24 13 1 10 9 12 9 0 13 10 9 1 10 9 7 10 0 1 9 13 1 9 1 9 2
12 10 9 1 10 9 1 10 9 3 13 13 2
31 10 9 0 1 10 11 3 13 10 9 1 10 9 1 10 9 1 10 11 1 13 10 9 1 9 0 1 10 9 0 2
62 1 10 9 1 16 10 9 1 10 9 0 3 13 1 10 9 1 9 1 10 11 3 1 10 9 0 1 10 11 7 10 11 2 11 13 16 15 13 13 10 9 1 9 13 3 13 10 9 1 10 11 2 7 10 9 0 7 0 1 10 11 2
6 9 1 10 9 13 9
12 9 7 0 13 3 10 9 12 1 10 11 2
11 13 9 2 15 13 10 9 1 9 0 2
10 13 10 9 1 9 1 9 3 0 2
16 10 9 0 13 13 3 10 9 1 9 1 10 9 7 9 2
6 9 1 11 13 9 0
19 10 9 0 0 13 0 1 13 10 9 0 1 10 9 0 1 10 11 2
23 1 15 13 1 13 10 9 2 10 11 13 1 10 10 9 0 10 9 1 10 9 0 2
12 15 3 13 10 9 1 9 0 1 10 11 2
26 15 13 10 9 1 10 11 1 11 2 11 2 2 10 1 10 3 0 9 1 9 0 1 10 11 2
29 2 10 9 3 3 13 3 9 2 16 10 9 13 1 13 2 2 13 1 10 11 10 9 11 2 1 10 11 2
20 10 0 13 16 1 10 9 3 15 13 10 2 9 2 1 10 9 1 11 2
42 10 9 0 2 11 2 13 9 1 10 2 9 2 3 13 3 1 10 9 7 13 1 11 3 10 0 9 2 0 1 10 9 1 9 2 1 10 9 1 10 9 2
21 15 2 3 7 3 2 13 1 10 9 1 16 15 13 10 9 1 2 9 2 2
22 10 9 11 2 15 3 13 9 1 10 9 2 15 13 1 15 13 3 0 1 13 2
6 2 13 10 9 0 2
11 3 13 4 13 1 10 9 1 9 2 2
20 10 9 2 3 2 2 11 2 13 2 13 16 13 2 3 16 9 3 9 2
26 10 9 11 13 10 2 9 2 0 2 1 13 10 9 1 10 9 1 13 15 3 9 1 10 9 2
27 10 9 2 13 9 0 7 0 9 1 9 16 10 9 0 2 2 13 10 9 1 10 0 9 2 11 2
29 9 1 10 11 1 11 2 11 2 13 10 9 1 10 0 9 1 10 9 1 10 11 2 2 2 11 2 2 2
32 1 15 2 10 11 13 13 10 9 1 11 2 11 2 11 2 11 7 11 2 11 2 11 7 11 2 11 2 11 7 11 2
9 10 9 13 13 0 1 15 9 2
31 10 9 11 7 9 11 13 3 1 10 9 7 10 9 11 2 10 9 11 7 10 9 11 13 13 1 10 9 1 12 2
28 13 2 11 2 12 2 3 13 12 1 10 9 1 10 11 1 10 9 1 10 9 1 10 9 1 10 9 2
21 10 9 13 1 10 9 1 12 9 7 2 1 9 2 13 1 10 9 1 0 2
10 11 13 10 0 9 3 1 10 11 2
5 2 13 3 13 2
18 10 9 13 13 0 7 15 13 13 3 13 13 10 9 2 2 13 2
12 1 10 9 2 10 9 13 13 1 10 11 2
13 2 3 13 13 3 3 7 13 10 9 3 2 2
19 16 10 9 11 13 1 10 9 2 11 13 3 10 10 9 1 10 9 2
17 3 1 10 9 1 11 2 15 12 13 0 13 10 2 11 2 2
2 13 2
81 9 0 2 1 10 9 13 7 13 1 9 2 1 15 13 9 1 9 1 9 1 9 1 9 7 1 9 15 13 10 9 13 1 10 9 1 10 9 13 2 10 9 1 10 9 2 1 9 1 9 2 13 13 1 10 9 1 10 9 1 10 9 7 2 3 2 1 9 2 13 10 9 12 1 10 9 9 12 1 12 2
35 9 0 2 10 11 2 11 2 3 13 4 13 1 10 9 13 1 10 9 0 2 1 9 0 2 1 9 2 1 9 0 7 1 9 2
9 13 15 1 10 11 3 1 10 9
11 9 3 13 0 1 10 9 1 9 7 9
5 1 10 2 11 2
24 10 9 15 15 13 3 15 13 13 1 10 9 13 1 9 13 0 1 15 1 10 9 0 2
26 1 10 10 0 9 2 13 3 10 10 9 15 1 10 0 9 15 13 9 0 2 13 7 15 13 2
12 13 13 10 10 9 1 13 1 13 10 9 2
34 1 13 10 9 2 10 12 0 9 3 0 1 15 13 1 9 1 10 11 13 13 1 0 0 9 0 7 13 3 12 9 1 9 2
18 15 7 10 9 2 9 1 0 9 2 3 3 0 2 13 10 9 2
17 10 10 9 13 13 1 10 11 2 9 1 9 12 2 1 9 2
21 10 9 13 1 10 2 0 9 2 1 10 9 1 13 3 2 9 3 15 2 2
16 7 15 13 1 10 9 1 10 9 11 2 16 3 15 13 2
4 3 13 0 2
25 10 9 13 1 10 11 2 13 1 10 9 1 12 1 10 9 13 1 10 9 11 2 10 9 2
19 11 2 12 2 12 1 10 9 1 10 9 2 13 10 9 1 10 9 2
50 3 2 10 9 13 9 2 13 9 2 13 9 2 13 10 9 2 10 0 9 1 10 11 2 15 13 9 0 2 15 2 13 4 2 16 4 1 13 1 10 9 2 15 15 3 3 13 9 0 2
37 13 9 2 9 7 13 2 1 10 9 0 1 9 12 1 9 2 7 13 3 1 10 9 15 2 3 13 11 2 13 2 0 1 13 13 2 2
3 15 3 2
3 15 13 2
11 10 0 9 1 9 11 2 12 2 13 2
21 13 9 1 10 11 2 11 13 0 10 10 9 0 2 15 2 13 1 13 2 2
8 2 13 0 3 2 2 13 2
28 10 9 0 13 10 9 0 1 10 9 1 10 9 2 13 10 0 2 9 2 2 9 13 1 0 1 9 2
29 1 13 10 9 1 10 9 1 9 13 2 10 9 13 1 10 9 1 10 9 7 6 2 13 13 10 9 0 2
34 3 2 13 9 1 9 1 10 9 0 1 10 0 9 2 1 0 1 10 0 9 2 3 15 13 10 9 1 9 1 10 9 0 2
27 10 9 1 10 9 0 13 10 9 1 10 9 1 9 3 0 2 9 15 13 0 9 1 10 9 0 2
22 1 10 9 1 10 11 2 10 9 0 1 9 13 13 1 12 9 1 9 1 9 2
13 1 10 9 13 2 10 9 13 12 9 1 9 2
7 9 1 10 11 13 1 11
23 10 9 1 10 11 1 10 11 2 11 2 12 2 13 1 10 9 1 9 3 1 11 2
37 15 13 0 10 11 12 1 0 9 1 10 11 2 1 10 11 2 9 0 2 2 3 2 3 2 13 10 9 1 10 9 7 13 1 10 9 2
22 3 2 10 11 7 10 11 2 3 2 13 9 3 0 12 5 7 12 5 2 3 2
27 10 9 13 16 10 9 1 12 13 1 12 5 1 12 5 10 9 0 1 10 9 1 10 11 1 12 2
7 9 1 10 9 13 9 0
26 10 9 1 10 9 2 11 2 13 10 9 1 10 11 3 1 13 15 1 10 9 0 1 10 9 2
45 2 13 3 9 0 2 1 10 9 0 2 0 7 0 1 15 10 9 0 1 10 9 2 2 2 13 13 3 10 9 15 10 9 13 2 2 13 2 1 9 13 1 10 9 2
8 11 13 1 9 1 9 1 11
12 10 9 1 11 13 13 10 0 9 1 9 2
40 10 9 1 10 9 1 10 9 1 9 1 11 13 1 9 0 1 10 11 2 11 2 11 2 11 2 11 2 11 2 11 7 11 2 1 10 9 11 2 2
13 10 9 0 13 1 12 1 13 10 9 1 11 2
11 2 13 10 9 15 3 13 1 15 13 2
27 13 1 10 9 1 10 9 7 3 13 15 1 10 9 0 2 2 13 11 2 12 2 9 1 10 11 2
28 1 10 9 1 9 1 10 11 2 11 2 2 3 13 0 9 2 3 13 4 13 10 9 15 13 13 2 2
36 15 13 10 0 9 1 9 1 9 1 10 9 1 11 1 10 9 3 10 0 9 1 9 1 10 9 1 10 9 1 10 9 1 10 9 2
23 1 10 9 2 3 9 1 10 9 1 9 13 13 1 10 9 1 2 9 2 7 9 2
20 10 0 13 1 10 9 1 9 13 1 10 9 1 10 9 0 1 10 9 2
30 10 9 13 1 4 13 16 9 15 13 1 10 9 1 11 13 13 16 10 9 13 7 13 10 9 13 1 10 9 2
20 10 9 13 13 7 3 13 10 9 7 13 10 9 3 1 12 9 1 9 2
74 1 10 9 2 9 1 10 9 15 13 3 12 2 7 12 9 0 2 10 11 2 15 3 13 13 0 7 13 11 7 11 1 10 9 2 7 10 11 2 15 13 10 16 10 9 1 10 9 1 9 1 10 11 2 1 10 9 1 9 1 10 9 1 10 9 2 11 2 2 11 2 3 13 2
7 9 13 1 10 10 9 2
35 10 0 11 13 10 9 7 13 12 9 0 1 10 9 1 10 2 9 2 11 7 13 9 1 10 9 1 9 2 11 7 1 10 11 2
12 1 10 9 2 10 11 13 10 9 3 0 2
19 2 16 15 13 12 5 1 10 12 9 2 13 16 15 13 13 10 9 2
9 13 13 15 13 1 10 9 2 2
6 11 13 3 10 11 2
29 10 9 3 15 13 1 9 15 13 1 12 5 1 12 5 1 10 9 1 15 13 2 13 2 9 0 7 9 2
18 3 1 10 9 1 12 9 7 12 9 3 10 9 13 10 0 9 2
21 13 12 5 1 0 7 0 2 12 5 1 0 7 0 7 12 5 1 9 0 2
1 9
37 10 0 9 1 11 1 9 0 13 1 10 9 1 15 15 13 10 9 1 10 9 7 13 1 9 1 0 9 2 3 10 9 1 10 9 11 2
2 9 13
20 10 11 0 9 0 1 9 0 13 13 13 9 12 12 1 10 9 1 9 2
22 10 9 2 15 13 9 12 9 1 12 2 13 13 1 9 10 12 9 1 10 11 2
7 10 9 13 13 10 9 2
19 10 9 2 3 2 3 13 15 13 13 3 1 10 9 1 10 0 9 2
19 15 16 10 9 1 9 3 13 3 10 9 1 9 12 9 1 10 9 2
13 13 3 13 10 9 1 12 9 1 10 12 0 2
9 1 3 2 10 9 13 3 13 2
10 10 9 13 3 0 1 10 0 9 2
22 11 2 9 1 10 11 1 10 11 2 13 1 9 10 9 1 12 5 7 12 5 2
20 10 9 13 13 7 13 10 11 1 10 0 9 2 1 10 9 12 7 12 2
19 10 10 9 11 13 9 1 10 10 9 1 13 10 10 9 1 10 9 2
25 10 9 11 13 13 1 9 1 10 11 1 10 9 1 10 9 13 1 10 9 15 13 10 9 2
16 1 10 9 2 13 11 2 10 9 13 13 0 1 10 9 2
23 10 0 9 13 13 1 10 9 1 9 1 10 11 2 15 13 3 1 12 9 1 9 2
21 3 13 13 1 10 10 9 10 12 9 1 10 11 2 10 9 0 1 10 9 2
19 2 15 13 1 10 9 9 1 10 9 2 2 13 10 9 11 2 12 2
2 10 9
32 1 10 9 1 9 1 9 1 9 0 2 9 11 13 13 1 10 9 16 10 9 1 10 9 13 4 15 13 1 10 9 2
27 9 13 1 13 9 1 9 1 15 7 12 9 1 10 2 1 10 9 2 15 13 9 0 1 9 9 2
3 2 0 2
3 2 0 2
20 3 15 13 1 10 9 15 13 16 10 9 3 13 10 9 3 13 16 15 2
36 7 2 9 1 10 9 2 13 10 9 15 13 10 9 3 13 16 10 9 2 13 1 13 10 9 2 15 3 1 10 9 1 10 9 2 2
35 13 16 10 11 2 10 15 15 13 10 0 11 2 13 10 9 1 2 9 2 2 3 9 15 13 10 9 1 9 0 3 1 10 9 2
10 2 11 2 13 10 9 1 13 9 2
16 1 9 2 13 9 1 9 1 9 2 9 2 9 7 9 2
8 13 9 12 2 1 10 11 2
3 9 12 2
19 2 11 2 13 10 9 1 9 2 13 1 9 15 13 13 9 1 9 2
9 13 4 13 1 10 11 1 9 2
8 13 1 9 12 1 9 12 2
11 2 11 2 13 10 9 1 9 1 9 2
16 13 1 9 1 9 7 9 2 15 13 10 9 1 10 9 2
11 13 9 12 1 10 11 2 9 12 2 2
32 15 13 2 3 2 16 10 9 9 13 1 10 9 13 10 9 15 10 9 13 13 1 10 9 15 13 10 9 1 10 9 2
21 11 2 1 10 9 0 11 2 13 2 16 3 13 0 10 9 9 1 10 9 2
19 7 13 16 10 9 9 13 1 10 9 13 10 9 0 1 10 9 0 2
31 1 10 9 1 10 9 2 10 9 0 13 13 1 13 10 9 1 10 11 2 9 0 1 10 11 2 3 1 10 11 2
24 10 9 0 1 10 11 2 11 2 13 3 1 11 16 10 9 1 10 9 1 9 13 13 2
25 11 13 16 10 11 13 13 16 3 3 13 10 9 1 11 13 10 9 12 12 13 1 10 9 2
8 11 2 10 9 13 15 13 2
8 11 2 1 15 13 10 9 2
7 2 11 13 1 13 2 2
9 13 3 15 13 3 15 2 9 2
5 16 13 3 13 2
6 2 13 15 1 13 2
9 9 13 9 1 12 9 1 10 9
36 10 9 1 10 11 2 11 2 2 1 10 11 2 13 3 2 13 13 2 1 10 9 1 9 1 10 9 1 9 2 10 9 1 12 9 2
21 1 9 1 10 9 2 10 9 13 10 9 1 10 0 9 1 12 5 1 12 2
20 10 11 2 11 2 13 1 10 9 1 9 1 12 9 15 13 9 1 9 2
45 1 10 9 1 10 11 2 11 2 10 9 1 10 9 3 13 13 1 10 9 2 13 1 10 9 0 1 10 9 3 10 0 9 1 10 9 1 9 1 10 9 1 10 9 2
29 1 15 2 10 9 1 9 1 10 9 1 10 0 9 13 4 13 1 10 9 0 3 10 9 7 15 1 9 2
7 10 9 3 3 13 0 2
23 1 10 9 11 2 12 2 2 13 9 15 15 13 2 1 10 9 1 13 10 9 2 2
31 3 2 10 9 1 10 0 7 11 15 13 10 9 1 10 9 1 10 9 1 10 9 15 13 1 13 9 1 10 9 2
9 11 3 13 10 9 1 10 9 2
21 1 13 9 2 13 13 1 10 11 10 9 1 13 1 10 9 15 13 13 3 2
9 13 10 9 1 9 1 10 9 2
8 13 13 9 1 10 9 0 2
23 16 10 11 3 13 10 9 13 2 15 13 13 1 10 9 1 9 10 9 15 13 13 2
23 3 13 13 12 9 1 9 0 2 1 13 10 9 1 10 9 1 10 9 1 10 9 2
8 11 13 11 7 11 13 15 12
5 1 10 9 1 9
36 10 11 13 3 10 11 2 3 1 10 9 0 2 1 12 1 12 2 1 10 9 3 0 7 0 1 10 0 9 9 1 10 11 1 12 2
36 13 1 10 9 1 9 2 10 9 11 2 9 1 10 11 2 13 1 9 10 9 0 11 2 10 9 1 10 9 13 13 1 10 0 9 2
27 1 10 9 0 1 10 9 11 2 10 9 1 9 13 1 12 9 2 13 9 1 12 9 1 10 9 2
27 1 10 9 0 1 9 2 10 9 1 9 0 1 9 13 1 12 9 2 1 12 9 1 10 9 0 2
7 0 9 13 9 1 10 9
18 13 10 9 1 9 0 7 13 3 0 13 9 1 10 9 1 10 9
17 10 9 1 10 9 1 10 9 13 13 1 10 0 7 0 9 2
47 9 0 2 9 1 9 7 10 9 13 13 1 10 9 3 1 15 15 13 1 13 9 3 13 1 10 9 7 0 1 10 9 1 10 9 1 10 9 1 0 9 1 10 9 1 9 2
36 2 10 9 13 16 10 9 13 15 0 13 3 10 9 13 10 9 3 7 1 10 9 7 9 2 2 13 10 9 1 9 0 11 2 12 2
21 2 10 9 1 10 9 13 10 12 9 1 10 9 1 10 10 9 2 2 13 2
19 1 10 11 2 9 7 10 9 13 1 13 9 1 0 9 1 10 9 2
14 1 10 11 2 10 9 3 13 1 10 9 1 15 2
19 10 9 15 13 13 13 10 9 3 0 1 10 9 1 15 13 1 15 2
45 10 9 15 13 2 13 9 1 9 7 9 1 15 10 9 3 13 7 0 2 9 2 0 2 7 0 2 13 2 2 7 13 1 9 0 0 3 0 3 2 3 15 13 13 2
5 15 15 13 3 2
12 1 15 12 2 11 2 11 7 11 13 3 2
25 11 2 15 13 1 10 11 1 10 9 2 3 13 9 0 1 10 0 9 2 1 10 9 12 2
29 10 9 3 13 13 0 2 13 13 3 10 11 16 10 9 0 3 2 3 13 15 2 10 9 13 1 10 9 2
3 13 15 2
24 1 10 9 1 12 9 2 10 9 0 1 10 11 13 16 12 1 15 13 9 1 9 0 2
21 13 10 9 15 2 1 10 9 2 13 13 2 10 9 0 13 1 10 11 2 2
47 13 1 10 9 11 2 11 2 2 11 2 1 9 2 11 2 2 11 2 11 2 2 11 2 11 2 2 11 2 11 2 2 11 2 11 2 2 11 2 11 2 7 11 2 11 2 2
15 1 15 2 13 3 0 10 9 0 1 3 1 10 9 2
11 11 13 13 10 9 1 10 9 1 9 2
16 2 3 13 9 1 10 9 1 15 15 7 10 11 13 2 2
28 1 10 0 9 2 13 13 1 10 9 10 9 1 10 9 15 3 13 1 10 9 15 13 1 13 10 9 2
9 3 12 9 13 13 1 10 9 2
13 1 10 9 2 12 13 9 7 0 1 10 9 2
29 1 10 9 13 10 2 9 1 10 9 2 2 11 2 10 9 11 7 10 9 11 2 9 1 10 9 0 11 2
22 10 9 1 10 9 13 16 11 13 13 1 9 10 9 1 10 9 0 1 10 9 2
16 15 13 13 10 9 1 11 1 13 16 15 13 1 10 9 2
21 10 9 0 1 10 2 11 2 2 1 11 2 13 12 1 10 9 1 10 9 2
25 1 10 9 2 10 9 13 9 2 9 2 9 2 9 2 9 2 11 2 7 2 0 2 9 2
16 12 1 9 2 13 1 9 10 9 1 10 11 7 9 11 2
13 12 1 9 2 11 13 10 9 1 10 9 11 2
37 10 9 13 1 10 2 9 2 1 10 9 12 13 13 3 3 9 1 10 9 1 15 10 9 13 13 1 10 9 1 9 15 13 10 9 0 2
20 10 11 13 3 12 9 1 10 9 1 10 10 9 3 9 0 1 10 9 2
22 2 10 9 13 10 9 0 2 2 2 2 13 10 9 0 1 10 9 1 10 9 2
33 10 9 13 13 10 9 0 1 13 10 9 3 2 1 10 9 2 1 9 15 10 9 0 3 13 3 3 10 9 1 10 9 2
18 1 10 11 2 10 9 13 13 3 1 10 9 7 3 1 10 9 2
14 10 9 13 13 2 2 13 11 1 10 11 1 12 2
2 9 13
15 10 9 13 16 10 11 3 13 10 11 0 1 10 11 2
32 7 13 16 10 11 13 9 12 9 1 13 1 10 9 2 1 10 11 2 1 10 9 1 10 11 2 9 1 10 11 2 2
3 1 10 9
24 11 2 1 10 11 2 13 16 10 9 12 9 13 9 1 2 9 1 9 2 1 10 11 2
22 2 7 10 11 1 10 11 3 13 13 10 9 7 13 9 1 10 9 2 2 13 2
23 10 9 0 1 10 9 1 9 13 10 11 2 11 2 2 10 9 0 13 1 10 11 2
28 2 13 10 9 1 13 2 13 1 9 7 3 13 15 2 2 13 3 11 2 9 1 10 11 1 10 11 2
11 11 2 11 7 11 13 9 1 10 11 2
18 13 1 9 1 10 11 10 9 1 3 1 2 11 2 1 10 11 2
48 13 1 10 9 13 2 10 0 9 1 9 1 10 9 0 7 1 10 0 9 1 10 9 13 1 10 9 1 16 10 11 13 13 1 10 0 9 1 10 9 1 10 0 9 1 10 9 2
19 10 9 13 1 10 9 1 10 11 1 9 7 9 3 13 13 1 9 2
23 10 9 13 16 10 9 13 1 10 9 15 10 9 13 1 10 0 9 1 12 3 13 2
25 10 9 1 10 0 7 0 9 13 1 10 9 16 15 13 13 0 1 10 9 1 10 9 0 2
15 10 9 1 10 9 1 10 9 13 10 0 1 12 9 2
14 13 3 2 11 13 10 9 0 2 7 3 13 15 2
18 3 13 2 9 2 16 2 13 1 10 9 0 2 15 3 13 9 2
6 9 13 0 1 10 9
15 3 13 0 13 16 10 9 0 13 10 9 1 10 0 9
1 11
13 10 9 12 13 10 9 1 9 1 10 9 0 2
14 3 12 9 13 4 13 1 10 10 9 0 1 9 2
35 12 10 9 1 10 9 13 1 10 9 1 10 9 2 9 1 10 9 0 2 9 0 1 9 1 9 1 0 7 0 9 0 7 0 2
11 9 13 1 9 13 1 10 9 1 10 9
29 11 2 12 2 13 1 10 0 9 13 1 10 9 1 9 1 10 9 1 15 13 2 15 13 1 10 9 11 2
15 10 9 13 1 10 9 2 1 10 11 2 9 0 2 2
13 10 10 12 9 15 13 1 10 9 13 15 13 2
7 9 13 7 13 9 7 9
28 10 9 1 10 9 1 10 9 12 1 10 9 11 1 10 9 11 1 10 9 1 3 13 9 1 10 9 2
27 10 9 13 10 9 1 10 9 11 2 15 13 1 10 11 13 1 11 2 12 2 15 13 1 10 9 2
27 10 0 9 13 1 12 9 15 3 13 1 13 12 9 1 10 9 0 1 10 9 13 3 13 1 11 2
24 2 11 2 16 13 12 1 10 0 9 1 10 11 2 3 3 13 1 10 9 13 1 9 2
39 10 9 1 9 1 10 9 1 10 9 1 11 2 2 2 13 0 1 10 9 16 2 1 10 9 1 9 2 10 9 13 7 13 10 9 1 11 2 2
17 10 9 0 2 3 11 2 2 13 1 10 9 13 1 9 2 2
8 9 13 15 1 10 9 0 2
49 10 9 3 0 1 11 2 15 1 2 13 12 1 10 0 9 1 10 11 2 13 3 10 0 9 0 1 10 9 2 13 1 10 9 1 10 9 1 9 15 3 13 10 9 11 1 10 9 2
31 10 9 11 13 10 0 9 0 2 1 9 1 10 11 7 3 10 9 2 3 3 9 2 13 10 9 1 9 1 11 2
17 11 2 3 15 13 1 9 2 3 15 13 3 1 10 9 0 2
22 3 15 13 1 10 9 2 13 15 1 9 15 13 15 15 13 13 10 9 1 11 2
24 11 2 9 3 10 11 2 15 13 1 9 13 1 15 1 10 11 2 13 3 10 9 0 2
5 2 9 2 9 2
8 15 10 9 13 1 10 9 2
7 2 9 2 9 2 9 2
6 9 1 15 3 13 2
22 10 9 13 1 10 11 2 11 2 15 13 9 0 1 12 9 1 9 1 10 11 2
23 1 10 9 1 9 2 10 9 9 13 1 12 9 1 10 9 7 10 9 2 12 9 2
11 10 9 1 11 13 12 9 1 10 9 2
2 1 9
23 10 9 3 13 9 13 1 10 11 7 1 10 9 1 10 9 1 9 13 1 9 0 2
2 9 13
18 10 9 11 7 10 9 13 13 1 13 9 1 9 13 1 9 13 2
39 3 2 10 9 0 9 11 7 11 2 9 1 10 9 1 10 11 7 11 2 3 2 15 13 1 10 9 0 0 11 2 11 2 7 11 2 9 2 2
7 9 1 10 11 13 12 0
23 3 12 9 13 7 12 15 13 1 10 0 9 0 1 9 1 9 0 1 11 2 11 2
12 9 1 10 9 11 13 9 1 10 9 11 2
5 13 10 9 1 9
22 1 10 9 1 10 9 1 10 9 2 13 13 0 1 10 9 0 1 10 0 9 2
25 9 2 13 10 9 7 9 1 0 9 1 10 9 1 9 7 9 13 1 10 9 7 9 0 2
12 1 13 13 10 9 1 11 2 11 13 13 2
12 2 13 10 9 2 7 3 13 10 10 9 2
8 3 3 13 10 11 1 15 2
10 15 13 10 10 9 2 2 15 13 2
15 1 11 2 13 13 10 9 1 10 9 0 1 10 9 2
17 2 13 10 9 1 10 11 7 15 13 3 13 10 9 3 2 2
41 10 9 13 1 11 13 10 9 1 13 10 9 1 10 11 15 13 13 10 9 1 10 9 1 10 9 1 10 0 9 12 2 3 13 10 11 13 1 10 9 2
21 10 9 1 11 3 13 13 16 10 9 0 13 16 10 9 1 10 9 13 13 2
28 15 13 10 9 3 13 1 10 9 1 10 9 2 3 2 15 13 9 1 9 0 1 10 9 1 9 0 2
30 1 10 9 1 3 2 10 9 1 12 9 13 13 13 1 10 9 1 10 9 1 11 2 12 9 1 9 1 11 2
25 10 11 13 3 12 9 1 9 1 11 7 12 9 1 10 9 11 2 1 11 2 1 10 11 2
2 0 9
23 10 0 9 15 15 13 9 1 9 0 1 10 9 13 1 10 9 1 10 9 1 12 2
1 11
32 13 16 10 11 2 11 2 2 13 1 10 9 1 10 9 13 2 13 13 10 9 2 11 2 3 9 1 9 1 10 11 2
1 11
16 13 9 13 1 11 2 9 1 11 7 11 1 10 9 11 2
27 10 9 13 16 10 9 1 10 11 13 3 13 1 10 9 1 10 9 1 10 9 16 13 13 1 3 2
26 3 1 10 9 13 1 10 9 1 13 10 0 9 2 10 9 1 10 0 9 15 13 10 9 13 2
8 10 9 11 13 1 10 9 2
26 10 0 9 13 13 1 10 11 2 15 1 9 1 12 13 10 0 9 1 9 13 1 9 1 9 2
47 10 11 13 3 12 9 2 9 12 9 2 1 10 9 13 1 10 9 1 10 11 2 13 3 10 0 9 1 10 9 1 10 9 0 1 11 7 10 0 1 10 11 2 13 1 12 2
7 9 13 9 1 10 10 9
23 10 9 11 2 9 1 10 11 2 13 1 12 1 10 9 15 13 10 9 1 10 9 2
25 10 9 1 10 9 2 13 1 12 9 2 1 11 2 1 10 9 11 2 13 3 10 9 11 2
1 9
22 3 1 13 10 9 1 9 1 10 9 11 1 11 2 10 0 9 11 13 15 12 2
