5396 17
8 3 2 13 9 9 12 13 2
30 7 2 2 9 0 9 0 7 0 13 13 7 9 0 7 0 12 9 13 9 0 13 9 13 9 2 13 4 11 2
12 11 10 13 4 12 9 2 9 13 0 9 2
8 15 7 14 7 13 4 13 2
19 11 2 11 2 11 2 11 2 11 7 0 11 9 0 13 4 9 10 2
24 11 9 4 11 9 9 13 4 7 2 10 9 11 13 4 2 13 13 4 10 9 9 10 2
17 15 9 0 4 11 2 7 9 13 9 0 13 2 12 9 13 2
9 7 2 15 9 13 9 13 4 2
16 9 13 13 4 2 9 13 4 2 7 15 13 4 9 9 2
3 10 13 2
7 11 12 9 9 9 13 2
12 0 9 2 7 2 9 13 4 3 13 4 2
5 2 9 0 13 2
19 11 9 9 9 13 4 7 2 9 13 9 9 13 2 9 13 13 4 2
19 2 9 10 14 4 9 9 13 2 9 0 13 9 10 7 0 9 7 2
10 11 3 13 11 9 10 13 4 13 2
14 13 9 12 0 13 4 11 9 2 7 10 0 13 2
17 7 2 12 9 11 11 9 9 13 4 2 9 0 9 13 9 2
7 2 13 4 11 9 2 2
9 12 9 10 13 13 9 13 4 2
10 9 13 13 2 7 9 13 9 13 2
9 2 9 14 13 9 12 9 13 2
18 11 11 7 11 11 13 2 7 9 13 13 0 9 2 7 11 9 2
15 10 14 4 13 2 7 12 9 13 4 10 10 13 4 2
16 9 9 10 13 4 2 3 13 4 2 7 11 13 13 4 2
4 9 9 13 2
9 3 0 13 9 9 13 13 4 2
10 12 9 0 3 13 2 9 9 9 2
11 9 0 13 9 13 7 3 9 13 4 2
6 3 9 13 13 4 2
14 11 9 7 2 11 11 0 9 10 9 13 4 13 2
14 0 13 9 13 2 7 13 9 13 3 0 13 4 2
18 12 9 9 0 13 4 7 2 11 9 12 9 13 3 9 13 3 2
20 11 9 9 14 4 9 0 10 9 9 13 2 9 9 2 10 9 0 13 2
14 9 9 11 11 13 4 2 7 11 11 13 4 9 2
12 15 9 9 0 9 9 13 2 9 9 13 2
16 9 2 13 4 13 2 13 4 9 0 2 13 7 0 13 2
17 9 9 9 9 2 7 2 13 13 4 7 0 9 13 13 4 2
26 9 2 9 7 9 0 0 9 0 13 9 13 13 9 10 3 15 13 14 4 9 7 9 0 10 2
5 3 13 13 10 2
10 11 11 9 0 14 4 9 10 13 2
8 11 9 12 13 4 9 9 2
14 9 10 12 9 3 11 11 9 9 13 4 9 10 2
7 12 9 14 4 3 13 2
15 14 4 9 9 3 13 2 7 0 10 9 0 13 4 2
13 9 9 0 9 13 4 2 3 2 9 7 9 2
24 11 9 2 7 2 9 0 13 4 2 7 11 9 2 9 9 0 12 13 4 2 12 2 2
5 2 13 4 2 2
25 9 13 9 10 11 2 12 2 9 13 4 9 9 13 9 2 7 9 11 2 9 2 13 4 2
8 7 2 3 9 10 13 4 2
22 9 12 0 9 13 9 13 4 11 2 9 0 9 13 2 7 9 13 4 12 9 2
14 9 0 9 13 4 9 7 10 13 4 9 13 9 2
5 2 9 13 4 2
10 13 13 9 3 9 9 0 13 4 2
9 9 9 9 13 9 9 13 4 2
15 14 4 9 9 3 13 2 7 3 13 9 13 13 4 2
6 11 9 13 9 13 2
4 13 9 9 2
13 7 2 3 2 12 9 13 9 9 9 13 2 2
6 9 13 2 13 4 2
12 11 11 0 7 11 11 11 7 9 13 4 2
7 9 9 9 7 13 4 2
10 14 4 13 2 7 9 3 13 4 2
8 10 9 0 13 4 13 9 2
14 2 9 13 4 15 14 13 3 11 11 7 11 2 2
6 11 13 4 9 13 2
7 7 10 13 3 13 3 2
12 3 2 11 9 0 12 2 9 13 4 9 2
18 9 10 13 3 11 9 12 9 13 13 4 9 9 9 13 13 4 2
10 13 4 9 9 10 13 7 13 9 2
15 3 2 11 13 7 11 13 4 2 3 9 13 4 9 2
19 10 9 2 9 9 7 9 0 9 3 13 2 3 13 4 9 9 10 2
10 11 9 9 12 13 13 4 9 11 2
5 9 13 13 9 2
11 3 9 0 7 12 9 13 7 13 4 2
7 2 9 9 9 12 13 2
5 2 9 13 4 2
8 11 11 13 9 9 13 4 2
16 2 11 3 9 0 13 2 3 13 7 9 3 3 13 4 2
13 15 7 3 13 13 4 2 3 13 4 9 2 2
16 15 9 3 9 13 2 10 3 13 3 2 15 9 13 13 2
10 0 0 12 9 13 2 9 13 0 2
11 11 12 9 0 0 13 4 9 7 9 2
16 9 9 9 10 13 4 12 9 2 3 10 9 13 13 4 2
13 11 9 13 4 2 11 11 0 9 13 3 13 2
17 9 12 2 10 7 10 13 2 3 13 4 14 9 7 14 9 2
16 11 3 13 4 3 2 7 9 0 13 10 9 12 13 4 2
7 7 9 13 4 15 9 2
11 10 9 0 13 4 3 11 7 11 13 2
6 14 9 13 9 13 2
13 11 9 9 9 0 13 2 7 9 13 0 3 2
11 2 9 12 9 10 13 4 9 13 9 2
10 7 3 13 4 2 7 10 13 9 2
28 7 2 11 9 13 4 2 11 9 13 4 9 9 12 9 13 4 13 2 7 3 14 4 9 9 13 13 2
10 14 13 13 9 9 13 9 13 4 2
17 9 13 2 9 9 13 9 13 2 7 9 13 13 9 13 2 2
8 11 9 9 7 13 4 9 2
7 9 11 12 9 13 4 2
5 9 9 13 13 2
15 9 12 13 11 9 13 4 9 9 9 9 9 13 4 2
13 9 13 9 10 9 13 4 2 9 2 13 4 2
8 11 9 9 9 13 4 9 2
13 11 9 13 4 11 2 2 9 13 2 4 13 2
13 11 13 13 4 9 2 7 11 11 13 13 4 2
16 9 3 13 4 13 2 7 9 9 13 4 9 2 12 2 2
6 11 9 13 13 4 2
18 9 0 13 9 9 2 9 0 9 2 13 4 2 9 13 4 9 2
5 9 13 4 10 2
6 9 10 9 9 13 2
22 9 13 9 11 9 0 9 0 13 4 7 3 13 4 11 10 9 7 9 9 9 2
11 9 12 13 4 9 0 13 2 0 13 2
7 9 10 13 4 9 9 2
7 11 14 4 9 13 11 2
10 11 9 13 4 2 9 0 9 13 2
5 11 9 13 10 2
8 9 0 13 9 13 13 4 2
6 9 13 2 7 9 2
13 10 9 2 0 9 10 2 13 9 9 13 4 2
17 11 9 10 13 4 12 9 13 2 7 10 7 3 0 13 13 2
20 9 11 2 11 2 11 2 11 2 11 7 11 9 9 13 4 2 12 5 2
18 9 9 3 13 4 2 3 9 14 13 7 3 9 0 13 4 2 2
14 3 13 4 9 10 9 11 11 0 7 11 11 0 2
15 6 2 9 9 13 2 7 9 13 10 9 13 9 13 2
28 9 2 9 0 13 10 0 10 13 4 9 0 13 2 7 0 2 7 2 9 0 13 7 0 13 9 4 2
17 9 9 13 13 9 0 9 9 0 2 0 9 13 4 3 13 2
16 12 12 9 3 13 4 9 2 7 12 9 9 13 4 11 2
11 2 0 9 13 9 13 9 0 13 2 2
9 2 11 13 4 9 11 10 2 2
9 9 12 13 7 9 12 13 4 2
10 9 9 13 14 2 7 12 13 4 2
13 9 0 0 10 13 4 2 7 2 9 9 0 2
5 11 13 9 13 2
10 9 13 2 13 13 4 11 13 4 2
7 10 12 13 9 13 4 2
11 3 2 11 9 3 13 4 13 4 11 2
11 9 9 0 9 7 9 9 12 13 4 2
11 11 13 4 9 2 11 9 7 11 9 2
9 2 9 13 2 9 4 15 13 2
20 13 2 9 10 13 13 2 12 9 2 0 9 2 9 0 0 12 13 4 2
9 11 9 3 13 4 9 13 9 2
3 6 13 2
16 9 0 12 13 7 9 0 13 9 12 9 12 13 13 4 2
21 10 9 2 2 9 13 10 13 4 9 13 9 13 2 7 12 9 0 13 4 2
11 9 9 2 0 2 13 4 2 11 9 2
8 11 7 11 13 3 0 13 2
10 11 8 11 0 13 4 9 0 9 2
17 11 2 7 2 10 9 13 13 4 2 9 14 4 15 13 11 2
13 9 2 3 2 9 13 9 13 7 9 13 4 2
20 10 9 0 13 4 2 9 9 3 13 13 3 11 14 4 13 9 0 13 2
10 2 11 9 9 9 9 13 13 2 2
15 3 2 13 2 9 13 7 13 13 4 2 13 10 9 2
8 9 13 4 9 9 9 13 2
7 9 12 13 4 11 13 2
17 2 12 9 0 13 4 11 2 7 10 13 4 9 0 13 4 2
22 11 11 0 8 12 9 10 7 12 9 10 13 4 11 2 12 9 12 9 9 13 2
13 9 13 13 9 9 9 15 9 3 3 13 4 2
11 11 11 9 3 13 4 2 0 13 11 2
21 9 11 9 13 11 9 13 4 2 13 9 9 13 3 13 12 9 9 13 4 2
9 3 13 4 12 9 0 13 9 2
16 9 0 13 10 2 13 9 9 9 0 13 2 9 7 11 2
13 2 9 9 9 13 9 12 13 14 4 13 2 2
7 7 9 0 13 4 13 2
25 11 11 11 9 2 7 2 12 13 4 9 9 10 2 13 4 9 10 9 12 9 9 9 13 2
4 2 13 3 2
8 2 9 10 9 11 13 2 2
9 3 13 3 2 9 13 4 3 2
9 2 9 13 9 13 10 9 13 2
5 13 9 13 13 2
17 9 13 3 12 9 2 11 11 9 14 4 3 11 9 9 13 2
13 11 7 11 9 9 9 13 13 4 11 7 11 2
22 9 13 4 9 12 2 9 10 9 0 13 4 2 3 9 9 13 12 9 13 4 2
18 12 12 9 9 9 9 13 4 2 7 11 9 9 0 12 13 4 2
9 9 13 9 14 4 13 9 13 2
12 9 2 9 7 9 0 13 9 10 9 0 2
5 13 4 9 9 2
13 0 9 13 4 9 2 7 10 9 13 4 2 2
20 2 14 13 9 10 9 13 13 2 7 15 7 9 13 4 11 2 3 2 2
6 2 9 13 13 9 2
15 11 13 4 11 11 9 0 2 9 2 9 7 9 2 2
9 9 10 13 4 2 9 13 4 2
8 7 2 15 9 12 13 4 2
20 9 0 12 9 10 3 13 4 2 2 9 0 2 0 9 13 4 9 7 2
15 11 11 9 3 13 4 12 9 10 2 7 0 13 13 2
14 9 11 12 9 13 2 7 9 0 13 4 10 12 2
10 3 13 9 9 0 9 13 13 4 2
16 9 12 13 4 11 2 7 3 11 13 4 2 9 9 13 2
12 9 0 13 9 12 9 7 10 9 13 4 2
21 3 13 9 2 12 2 9 0 9 0 13 2 7 9 13 13 2 9 2 9 2
14 9 2 7 2 3 0 13 4 9 11 9 10 13 2
31 11 9 12 9 9 13 4 9 9 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 7 11 9 2 3 2
5 11 9 13 4 2
17 11 7 11 13 4 9 9 13 11 13 9 3 13 14 13 3 2
5 9 13 9 13 2
5 10 10 13 4 2
21 14 13 9 2 10 9 3 9 13 4 7 2 3 13 13 7 4 13 13 4 2
6 2 13 4 11 2 2
13 12 9 3 3 13 4 7 10 9 0 13 4 2
17 3 9 12 9 13 4 11 2 12 2 12 2 12 7 12 2 2
10 2 9 9 13 4 15 9 9 13 2
8 9 11 13 4 2 9 12 2
10 9 9 2 11 7 11 13 4 9 2
20 9 10 9 13 10 13 4 9 10 2 7 9 2 12 9 13 9 13 4 2
10 3 2 9 13 2 9 0 13 4 2
16 9 12 14 13 9 11 13 9 13 2 7 9 10 13 4 2
8 3 13 7 2 9 3 13 2
16 15 12 9 9 13 3 9 3 0 13 4 7 2 13 4 2
6 2 9 12 13 4 2
3 13 4 2
11 7 9 10 9 13 4 10 9 13 9 2
6 9 10 13 4 9 2
11 2 11 2 2 13 3 13 4 9 9 2
10 9 11 13 4 7 10 3 13 4 2
5 3 13 9 13 2
16 12 9 13 11 11 11 0 2 7 9 9 9 13 4 9 2
6 10 2 10 3 13 2
9 7 9 9 3 13 13 13 4 2
14 11 11 9 9 7 3 9 9 0 7 3 13 4 2
5 9 9 7 13 2
6 9 9 13 4 9 2
7 10 10 13 3 2 13 2
17 2 9 13 4 12 9 13 4 11 9 7 12 14 4 3 13 2
9 2 9 14 4 3 13 2 2 2
11 11 9 2 11 2 9 0 2 13 4 2
22 3 9 0 12 9 13 2 9 9 0 9 13 4 3 2 9 0 13 11 9 9 2
7 14 13 9 13 4 0 2
12 0 13 4 2 9 13 13 13 4 13 4 2
9 9 13 4 9 2 9 2 9 2
10 15 2 9 13 2 9 0 13 4 2
12 11 0 9 13 4 11 2 0 9 11 13 2
25 11 7 11 9 13 4 9 13 2 0 13 4 11 9 0 12 12 9 7 3 13 4 9 9 2
17 10 2 11 9 10 13 4 9 2 0 12 2 13 13 4 11 2
20 9 3 13 4 2 7 3 13 4 2 14 13 3 2 7 9 12 0 13 2
11 3 13 4 9 12 9 13 7 3 13 2
23 0 9 9 9 12 13 4 7 3 13 4 9 13 9 2 3 13 4 3 13 4 9 2
12 9 10 9 13 7 9 3 13 4 9 0 2
10 10 10 13 3 10 9 10 13 4 2
13 7 2 9 12 9 13 4 2 12 13 4 9 2
7 13 13 12 9 3 13 2
3 9 13 2
31 9 9 13 4 11 2 9 0 13 4 9 0 2 13 9 13 13 7 13 9 13 13 2 9 7 9 9 13 4 11 2
11 9 9 0 10 9 2 9 2 13 4 2
7 3 2 11 13 4 11 2
8 11 13 4 12 7 11 12 2
10 9 0 13 4 11 2 11 7 11 2
10 9 9 0 13 4 3 11 7 11 2
13 7 2 14 2 15 9 13 3 9 0 13 4 2
11 12 7 12 9 9 9 12 13 4 9 2
4 9 13 4 2
6 2 11 3 13 4 2
13 9 11 13 4 10 12 9 14 4 9 12 13 2
16 9 14 4 13 3 13 4 9 2 7 0 13 4 13 4 2
11 9 10 9 9 13 4 7 3 13 4 2
12 0 13 12 9 15 13 2 7 3 13 4 2
11 9 9 12 9 13 7 12 12 13 4 2
10 9 9 0 7 9 0 13 4 9 2
11 9 13 2 11 9 2 7 11 13 9 2
10 9 13 9 13 2 9 13 4 2 2
7 9 13 2 3 13 13 2
16 9 13 4 2 7 12 9 9 13 13 4 2 3 13 13 2
12 9 13 4 7 2 9 9 2 9 0 13 2
10 9 9 12 9 9 9 13 4 11 2
12 9 9 10 0 13 9 13 13 4 10 9 2
14 12 9 9 13 4 3 9 0 13 7 0 9 13 2
22 3 2 9 2 9 3 13 2 9 2 15 9 2 9 9 2 9 9 2 13 4 2
15 0 13 15 9 0 10 0 13 4 7 9 0 13 13 2
10 12 13 4 9 2 9 11 9 9 2
9 7 14 4 9 11 3 3 13 2
6 9 9 13 9 13 2
4 9 0 13 2
11 9 13 2 12 9 9 13 9 0 13 2
10 7 2 0 10 14 4 15 9 13 2
8 9 10 9 9 3 13 4 2
20 9 10 11 2 11 2 11 8 9 11 2 11 2 11 7 11 9 13 4 2
8 9 13 4 3 13 4 11 2
8 12 9 9 13 13 11 3 2
18 10 9 9 2 10 14 4 13 2 7 9 10 13 9 13 9 13 2
13 9 9 10 13 13 4 13 2 9 9 13 3 2
10 3 2 13 9 9 0 13 4 11 2
8 9 9 9 8 0 13 4 2
14 2 11 10 9 13 4 2 7 3 15 9 13 2 2
15 9 10 13 3 7 13 4 10 9 13 4 11 9 3 2
7 7 3 13 7 13 4 2
7 15 0 13 11 14 13 2
7 0 13 4 3 9 9 2
18 11 9 9 2 2 14 11 2 14 11 9 3 13 14 13 10 3 2
22 12 7 12 9 9 14 13 0 2 7 0 13 12 9 9 0 9 13 9 10 9 2
16 2 11 7 11 3 9 13 10 13 2 3 9 0 14 13 2
14 9 13 2 9 10 9 9 9 7 9 13 13 4 2
9 7 12 9 0 10 13 11 9 2
14 3 12 9 13 2 7 3 10 13 4 10 12 9 2
8 3 2 12 9 10 13 4 2
12 10 13 9 13 10 9 12 9 13 13 4 2
10 3 3 13 4 15 9 9 13 9 2
16 9 12 9 9 13 13 4 2 7 12 9 13 4 11 9 2
15 9 13 4 3 2 9 9 9 9 13 4 9 9 9 2
14 9 10 0 13 9 9 7 9 0 12 9 13 9 2
9 9 10 9 0 13 3 2 3 2
20 9 13 4 15 9 0 2 7 15 9 13 13 4 9 11 2 9 13 2 2
6 11 10 9 13 13 2
18 11 12 9 9 13 4 2 7 9 12 2 12 9 9 13 9 13 2
11 0 9 0 7 0 14 4 3 13 13 2
12 10 0 9 12 13 4 2 10 13 13 4 2
14 11 9 12 9 2 11 7 11 11 9 2 13 4 2
15 11 9 9 11 2 11 9 9 9 13 4 2 12 2 2
7 2 9 13 9 13 2 2
5 7 9 13 4 2
8 12 9 13 9 10 13 4 2
20 11 2 9 9 13 9 9 13 3 13 4 9 10 2 9 13 7 3 13 2
8 4 13 10 9 13 9 13 2
5 9 13 4 3 2
7 14 4 13 0 7 9 2
5 9 13 4 3 2
15 13 4 15 9 2 13 15 9 2 13 7 9 9 13 2
8 2 3 7 13 13 9 10 2
23 11 2 9 0 2 3 13 14 4 13 13 4 11 2 7 11 14 13 15 9 9 13 2
12 9 13 0 9 10 2 9 14 13 9 0 2
11 12 9 2 9 9 7 0 13 4 0 2
8 13 9 12 11 2 9 13 2
13 9 14 13 0 9 2 7 9 3 13 4 9 2
16 12 9 11 13 12 9 7 9 13 4 3 11 9 13 4 2
7 0 9 13 9 13 3 2
20 9 0 13 13 4 2 7 9 13 13 4 3 13 9 2 9 0 10 13 2
13 11 9 13 4 2 0 0 9 13 4 11 11 2
24 0 9 9 13 13 2 7 3 13 9 13 2 9 13 13 2 3 13 3 2 9 13 2 2
9 7 11 13 4 3 9 13 4 2
4 3 13 9 2
4 10 9 13 2
6 7 11 13 13 4 2
11 9 10 9 13 7 3 9 13 13 9 2
8 11 9 14 4 13 9 9 2
5 2 13 3 2 2
9 11 9 13 4 9 9 13 4 2
9 0 13 2 13 7 9 13 4 2
8 14 4 3 10 3 9 13 2
8 11 12 9 13 9 13 3 2
7 10 13 9 0 0 12 2
4 13 15 13 2
3 9 13 2
14 11 11 9 0 9 0 13 9 13 9 13 13 4 2
11 9 13 4 7 9 14 4 13 2 7 2
12 9 13 13 13 4 2 13 4 9 9 13 2
4 13 4 9 2
8 11 9 9 13 4 11 11 2
5 9 12 13 4 2
11 9 0 13 7 9 13 9 2 9 13 2
14 10 10 12 9 9 12 7 9 9 7 9 12 13 2
14 11 9 13 9 13 9 12 9 9 9 14 4 13 2
7 13 4 9 13 4 11 2
14 3 2 10 13 7 9 12 12 9 9 13 9 9 2
11 13 4 2 7 13 9 13 13 0 13 2
21 11 3 13 2 11 10 9 0 9 13 7 3 13 13 4 9 0 12 13 4 2
5 9 0 13 3 2
11 9 12 9 13 9 13 4 12 9 9 2
10 3 2 9 0 0 13 4 9 9 2
8 11 10 13 7 0 9 13 2
8 2 2 14 2 2 13 4 2
14 11 11 11 9 9 13 4 3 9 9 12 12 9 2
17 9 2 9 2 9 7 9 2 7 9 13 4 9 9 13 2 2
12 3 0 13 4 2 3 13 15 9 13 9 2
18 11 9 0 13 4 2 3 9 3 9 2 7 9 10 13 4 11 2
27 9 11 8 3 10 13 14 4 7 2 11 9 10 13 4 9 2 7 9 9 12 9 13 4 11 9 2
8 12 9 13 4 9 9 13 2
12 3 9 0 13 4 2 9 0 13 4 3 2
18 3 14 4 13 2 3 14 13 9 13 4 13 9 2 11 11 9 2
13 2 11 9 9 13 9 0 14 4 9 13 9 2
8 3 10 9 10 7 13 4 2
14 3 12 10 13 4 11 7 10 7 13 13 4 3 2
15 11 9 9 9 13 4 11 9 13 9 7 13 4 11 2
9 11 2 3 2 12 9 13 4 2
18 3 3 13 4 2 9 10 13 13 4 2 7 9 0 3 0 13 2
11 2 12 12 9 9 0 9 13 4 3 2
7 9 9 13 2 9 13 2
5 11 9 13 4 2
7 9 14 4 0 13 9 2
22 9 13 9 9 0 13 9 13 7 13 3 2 9 12 7 12 5 0 13 9 13 2
25 11 8 11 13 4 2 2 11 2 9 9 12 9 13 9 12 9 13 13 7 13 7 4 2 2
15 11 11 15 9 10 13 3 13 4 2 7 10 13 4 2
11 2 9 7 9 13 9 9 12 13 2 2
3 3 13 2
5 0 13 4 12 2
7 9 0 9 10 13 4 2
16 11 2 9 13 9 13 2 9 10 9 0 13 13 4 3 2
5 3 13 4 9 2
7 2 13 9 9 12 2 2
7 2 9 9 12 13 4 2
5 9 9 13 4 2
9 9 13 9 2 10 9 13 9 2
18 11 2 7 2 12 9 9 9 9 13 4 9 9 13 4 13 4 2
7 13 2 12 13 4 11 2
7 9 2 9 2 9 13 2
21 2 9 9 0 13 0 13 12 9 13 9 13 2 7 9 3 0 13 10 2 2
6 3 9 9 13 4 2
17 9 13 13 9 9 9 2 7 11 2 11 7 11 9 13 4 2
11 13 9 9 13 7 9 9 9 13 13 2
13 9 9 2 9 0 13 2 9 9 13 13 4 2
10 3 2 12 9 13 4 0 13 9 2
8 9 7 9 13 13 0 13 2
13 9 13 7 13 4 2 3 9 7 9 13 4 2
8 2 14 4 15 3 3 13 2
19 7 3 11 9 13 10 13 4 7 13 3 2 9 3 13 4 9 13 2
7 11 9 13 4 10 9 2
8 9 9 7 9 9 9 13 2
11 9 3 0 9 7 14 3 9 13 4 2
12 9 9 0 13 13 13 4 9 10 9 0 2
16 3 2 9 2 9 7 9 9 9 9 13 4 0 0 13 2
12 3 2 3 12 9 13 4 9 0 13 4 2
10 9 11 13 4 13 9 13 11 9 2
19 2 9 13 4 9 9 7 11 9 9 7 9 13 4 9 13 13 4 2
9 11 7 11 9 9 13 4 11 2
6 2 11 8 0 13 2
9 9 13 9 12 9 13 13 4 2
8 9 12 9 9 13 9 13 2
17 13 9 9 13 2 9 14 4 9 10 9 13 9 9 13 13 2
8 9 7 14 4 3 0 13 2
30 10 13 2 11 12 9 9 13 4 13 12 9 0 9 13 2 12 12 9 2 2 7 11 9 9 13 9 13 4 2
9 11 9 11 8 11 8 0 13 2
8 10 9 13 13 4 11 9 2
6 3 14 4 15 13 2
6 2 9 9 13 4 2
17 7 2 3 9 12 0 13 4 7 2 3 13 4 9 3 9 2
19 12 9 0 2 9 2 15 9 7 9 10 9 13 13 9 13 13 4 2
12 3 2 2 9 0 2 13 0 13 13 4 2
7 10 13 9 13 4 9 2
10 12 9 2 9 0 9 13 13 4 2
6 2 9 13 9 13 2
5 9 10 13 4 2
22 9 3 13 4 3 11 9 13 2 7 9 9 13 13 4 11 9 2 9 0 9 2
15 11 3 7 3 13 4 9 10 9 2 9 13 4 9 2
10 0 10 2 11 9 9 13 9 13 2
7 7 9 2 14 13 9 2
17 12 9 11 9 0 12 13 4 2 7 9 11 7 11 13 4 2
6 12 9 13 12 9 2
11 11 9 0 9 3 13 4 13 4 11 2
21 11 9 13 12 9 10 9 13 4 3 13 4 10 12 9 13 12 9 9 9 2
10 11 11 0 11 13 4 13 12 9 2
11 9 10 13 2 7 2 14 4 15 13 2
16 11 9 10 9 9 12 9 9 13 4 11 9 13 4 9 2
11 10 13 9 10 13 4 9 0 2 7 2
9 9 10 3 0 13 4 10 9 2
10 11 2 7 2 9 0 12 13 4 2
14 9 13 9 11 9 13 4 2 11 11 9 0 13 2
17 12 2 11 13 4 9 9 13 3 9 9 9 9 0 12 13 2
8 11 9 15 14 13 13 4 2
15 3 2 9 9 10 13 4 13 4 2 11 7 11 9 2
13 3 13 4 9 2 9 13 7 11 11 9 13 2
7 7 11 3 13 10 13 2
17 2 9 12 13 9 13 4 2 9 9 10 0 13 13 4 2 2
12 9 13 4 9 0 3 13 4 9 0 11 2
15 3 13 4 3 2 15 9 9 2 9 7 10 9 13 2
13 11 14 4 9 13 2 7 3 9 0 13 4 2
17 9 3 13 13 4 3 11 11 9 9 9 11 12 9 9 9 2
14 0 9 9 9 9 13 9 2 13 13 13 13 13 2
10 11 13 9 7 9 9 9 13 4 2
13 3 13 4 9 2 9 9 13 4 7 9 13 2
12 9 12 9 3 13 4 2 11 2 11 2 2
11 9 10 12 9 3 9 13 4 9 9 2
14 12 2 11 9 12 2 11 4 9 13 13 4 11 2
9 11 2 9 0 2 13 11 9 2
11 9 9 0 13 4 7 9 12 9 13 2
7 14 13 9 0 9 9 2
16 3 2 7 2 10 9 9 13 4 9 9 7 3 13 4 2
16 7 9 13 13 2 7 2 13 4 9 2 13 4 15 9 2
5 12 9 13 4 2
11 15 0 2 9 12 13 4 9 0 13 2
10 9 15 7 2 7 2 14 4 13 2
13 9 13 9 9 2 9 2 13 4 9 13 11 2
14 9 10 2 11 7 0 9 13 4 9 9 9 10 2
7 2 0 13 9 13 4 2
21 9 9 12 13 9 12 9 9 13 9 2 10 9 13 7 10 10 9 13 4 2
23 3 13 4 2 9 0 2 13 4 2 11 11 11 11 9 0 9 9 13 14 4 2 2
11 10 9 12 9 9 13 9 13 13 4 2
13 11 11 2 12 9 0 9 2 13 4 11 9 2
10 11 2 11 9 12 9 13 4 9 2
15 11 9 9 14 4 3 13 2 7 9 9 9 10 13 2
19 9 9 0 9 0 0 9 12 13 4 2 7 10 9 0 9 13 4 2
6 2 11 9 13 4 2
12 9 9 3 0 13 7 2 9 13 13 4 2
15 9 2 3 13 4 9 7 0 9 2 9 13 3 13 2
6 3 11 13 13 4 2
7 9 10 13 4 0 9 2
13 14 4 3 13 13 2 7 0 13 4 9 13 2
13 11 9 9 13 4 9 0 2 9 9 0 2 2
21 9 13 13 4 2 7 11 9 0 9 9 12 9 13 4 2 0 3 13 13 2
19 11 11 9 9 13 4 12 11 9 13 4 3 9 12 9 13 4 9 2
9 11 9 0 2 11 12 9 13 2
7 11 9 11 9 13 4 2
19 11 2 9 2 13 4 9 13 4 2 13 4 2 7 14 4 3 3 2
16 7 2 12 9 3 13 4 9 2 12 9 9 0 13 4 2
11 9 2 7 2 9 13 9 14 4 13 2
19 3 9 10 3 13 4 11 9 0 2 12 9 2 2 7 14 4 13 2
9 15 9 14 13 9 2 0 3 2
9 14 4 9 13 7 13 10 13 2
6 9 9 13 4 0 2
18 9 13 4 9 3 13 2 12 9 3 13 4 2 7 3 13 4 2
16 9 9 9 0 2 9 9 7 9 13 9 0 13 10 9 2
5 10 13 4 15 2
12 9 0 7 9 9 7 13 13 0 9 13 2
11 10 2 9 9 13 4 9 10 13 4 2
9 10 2 13 9 13 9 13 4 2
20 9 2 9 2 9 9 2 9 2 9 2 9 2 9 2 13 4 9 9 2
21 9 13 3 2 9 12 9 11 0 13 9 10 13 9 13 9 12 13 13 4 2
15 3 14 4 13 11 2 7 9 0 10 9 13 9 13 2
22 11 12 9 13 4 9 12 9 2 7 3 13 4 7 2 12 9 13 4 9 13 2
18 3 12 9 12 13 4 2 11 13 9 9 0 7 0 13 13 4 2
8 9 2 7 2 0 9 13 2
13 12 9 13 9 2 3 12 9 0 9 13 4 2
17 0 9 9 13 4 2 13 9 9 10 13 4 11 0 9 13 2
14 9 2 9 0 10 13 2 13 9 13 3 9 10 2
8 11 9 7 14 4 9 13 2
6 13 4 9 13 4 2
14 0 10 9 10 0 9 13 7 15 9 9 13 13 2
19 9 10 0 9 13 9 13 4 7 9 9 12 9 2 0 3 2 13 2
24 13 9 13 4 2 7 9 9 3 13 4 2 9 0 13 13 4 7 2 9 9 13 4 2
12 15 13 4 15 13 7 14 4 0 9 13 2
12 2 9 9 13 2 7 10 10 0 13 2 2
4 9 11 13 2
13 6 2 15 9 10 13 9 13 2 3 0 13 2
12 9 7 13 4 9 7 14 4 9 0 13 2
7 2 3 9 0 13 2 2
35 3 13 4 11 0 13 4 9 2 11 9 13 4 9 0 12 14 4 13 7 2 7 9 10 3 13 4 3 3 13 4 9 9 0 2
7 13 12 9 13 4 11 2
10 0 13 0 9 9 0 13 9 13 2
10 9 10 9 13 4 10 9 0 13 2
4 10 13 4 2
15 9 11 11 0 13 4 2 7 9 11 11 0 13 4 2
19 13 4 9 9 12 13 4 9 9 9 11 9 2 7 12 9 13 4 2
12 9 11 9 13 4 7 13 4 9 13 0 2
11 2 13 9 13 9 14 4 9 13 2 2
8 11 11 9 0 13 4 3 2
19 11 9 9 0 13 2 9 9 0 7 13 9 2 7 9 9 13 4 2
14 2 3 3 13 4 13 7 0 13 13 7 13 4 2
4 13 13 13 2
11 9 0 13 9 2 9 13 13 9 13 2
5 11 13 4 9 2
7 9 9 13 4 9 10 2
4 10 13 4 2
10 13 4 9 14 4 9 0 13 7 2
17 11 2 11 2 11 2 11 2 11 2 3 9 13 13 4 11 2
14 11 11 9 9 13 4 9 9 9 2 11 7 11 2
12 9 13 9 0 9 13 13 13 4 11 9 2
7 11 9 7 13 13 4 2
4 15 9 13 2
17 9 13 2 9 9 13 9 7 2 13 9 14 4 9 13 13 2
7 3 14 4 10 15 13 2
35 2 9 13 9 11 11 13 9 13 4 2 7 9 0 9 0 13 4 2 7 9 14 4 9 13 2 9 9 7 9 13 9 13 2 2
13 11 9 11 13 9 13 12 12 9 9 13 9 2
3 13 13 2
13 11 11 0 13 4 12 2 7 11 11 0 12 2
6 9 10 13 9 9 2
27 9 12 9 9 13 4 2 12 9 13 9 2 7 9 10 12 9 10 9 12 9 13 9 13 4 11 2
10 3 9 3 13 9 0 9 9 13 2
12 9 12 9 13 2 7 11 9 9 13 4 2
6 9 13 9 13 9 2
28 3 13 4 14 4 9 0 13 11 9 2 0 9 13 4 2 7 11 9 9 9 9 9 7 9 13 4 2
8 11 9 10 9 13 4 3 2
7 2 9 13 2 9 9 2
17 9 0 3 13 2 9 0 14 4 3 13 9 9 0 9 12 2
18 11 9 3 13 4 11 0 9 2 7 9 9 13 9 7 9 13 2
7 9 9 7 11 13 9 2
9 9 0 13 2 12 9 13 4 2
10 11 11 14 4 3 13 11 11 9 2
11 9 9 13 4 7 9 9 9 13 4 2
18 12 9 9 9 13 7 3 13 9 13 4 2 0 2 11 11 9 2
8 9 10 9 0 13 4 9 2
7 10 11 9 13 13 4 2
11 9 13 4 9 2 9 0 9 13 9 2
18 11 13 4 9 10 3 9 2 7 11 13 4 12 2 12 9 10 2
14 13 3 9 13 14 4 10 9 0 3 0 13 4 2
3 13 4 2
11 9 10 0 7 9 12 9 9 13 4 2
12 11 9 9 13 4 2 9 9 0 9 13 2
12 7 2 3 15 14 13 15 13 4 11 9 2
12 7 9 13 4 11 11 9 0 12 9 9 2
8 2 6 2 13 7 3 13 2
16 11 9 13 9 13 2 15 9 2 13 13 4 11 9 0 2
10 9 9 9 9 9 9 13 4 3 2
17 11 7 11 2 12 7 12 13 2 0 9 13 2 9 0 13 2
4 0 9 13 2
7 11 9 13 4 11 9 2
18 3 2 7 2 11 3 13 2 7 10 9 14 4 9 13 9 13 2
9 3 13 4 9 13 4 9 12 2
8 9 9 10 13 4 9 2 2
11 11 13 4 9 9 13 4 2 12 9 2
9 2 0 2 13 4 10 10 9 2
12 0 9 9 13 4 7 9 9 9 13 4 2
5 11 11 3 13 2
14 7 9 13 4 3 2 9 0 0 15 13 4 13 2
9 11 9 12 9 0 10 13 4 2
9 9 13 3 7 9 10 13 4 2
8 9 9 13 4 11 11 9 2
14 11 10 9 12 13 4 9 2 11 9 9 13 4 2
12 11 2 7 2 12 13 4 7 12 9 13 2
4 7 0 13 2
9 11 7 11 14 4 3 9 13 2
9 3 13 4 12 9 11 9 9 2
6 12 9 0 13 4 2
9 14 13 9 0 9 10 9 13 2
9 3 13 4 9 9 13 9 7 2
12 2 10 13 15 9 0 2 7 3 13 0 2
16 13 2 11 11 9 13 7 10 9 13 13 4 11 7 11 2
16 2 9 0 9 0 13 4 2 7 9 7 3 0 13 15 2
3 11 13 2
14 10 13 7 2 9 10 9 13 4 9 13 14 13 2
5 10 9 13 4 2
9 2 11 2 10 13 4 0 10 2
3 10 13 2
9 11 9 0 7 9 0 13 4 2
24 11 13 14 13 0 2 7 11 9 9 0 13 13 4 2 7 3 13 13 4 10 9 13 2
11 2 9 0 7 0 12 13 13 4 2 2
18 0 9 9 7 0 9 13 4 2 7 10 13 4 13 14 13 9 2
9 9 9 13 9 0 13 10 9 2
9 12 9 13 4 3 9 9 13 2
8 14 13 15 13 4 9 9 2
4 3 3 13 2
17 12 9 11 11 0 13 4 2 7 9 9 11 11 0 13 4 2
8 9 10 10 9 7 13 4 2
13 11 9 13 4 2 7 2 9 13 4 11 11 2
8 3 9 9 13 9 13 4 2
9 10 10 13 4 9 13 13 4 2
8 2 13 9 9 13 4 9 2
8 2 11 9 12 9 13 4 2
15 3 13 7 13 9 13 2 0 13 4 2 7 15 9 2
8 12 7 11 9 13 13 4 2
8 9 13 3 13 4 9 0 2
10 11 13 9 7 9 9 9 13 13 2
10 9 9 13 4 2 9 9 9 13 2
7 9 13 9 2 9 13 2
12 2 9 9 9 9 12 9 10 13 4 2 2
5 12 9 13 4 2
19 9 3 0 13 4 2 13 4 9 0 13 4 2 7 9 0 13 4 2
9 9 12 9 13 4 9 13 13 2
3 10 13 2
10 7 2 9 13 9 13 0 13 4 2
6 15 9 2 13 13 2
22 11 12 9 0 13 7 9 0 13 11 9 11 9 0 7 11 11 9 13 9 13 2
8 9 0 9 13 2 0 13 2
10 9 9 13 4 2 7 3 13 4 2
6 11 11 13 13 4 2
13 0 12 9 2 7 2 9 13 4 12 9 9 2
12 3 2 9 7 9 13 9 0 9 13 4 2
8 12 2 9 13 9 7 9 2
14 3 0 13 4 9 9 9 10 13 7 9 9 13 2
25 12 13 4 11 9 9 12 9 13 7 2 11 2 9 9 0 0 13 9 13 9 13 9 13 2
9 13 4 9 12 13 4 11 9 2
8 9 9 9 13 9 13 4 2
11 9 10 14 4 9 12 13 4 9 13 2
19 9 7 11 9 13 4 9 9 9 11 11 7 11 11 9 13 3 9 2
7 2 14 13 2 14 2 2
14 9 3 13 4 2 9 14 4 9 9 13 9 13 2
5 9 3 13 4 2
7 3 13 4 9 11 9 2
15 11 9 9 9 13 9 13 3 9 13 9 0 13 9 2
25 3 7 2 11 3 13 13 4 7 3 2 12 9 12 9 2 9 9 13 4 13 4 9 9 2
17 7 14 4 15 9 13 2 7 10 15 9 13 7 13 9 13 2
6 13 9 7 0 13 2
12 9 10 2 3 0 13 4 15 9 13 2 2
7 9 13 9 0 13 4 2
15 2 9 9 9 0 12 13 9 13 13 13 0 13 4 2
6 13 4 10 13 4 2
9 9 0 0 0 13 7 13 13 2
8 3 11 12 9 0 13 13 2
8 15 9 10 9 13 4 10 2
8 9 7 9 10 13 4 9 2
13 10 13 4 9 0 13 9 9 13 13 9 9 2
9 11 13 4 14 13 9 13 13 2
8 7 2 9 13 11 13 4 2
6 11 14 13 9 0 2
8 9 0 13 9 9 13 4 2
10 11 13 9 14 4 13 11 13 9 2
5 2 13 13 4 2
8 9 9 13 9 0 13 11 2
9 9 0 13 9 0 13 2 7 2
14 9 0 13 4 9 2 7 9 14 4 0 9 13 2
13 13 3 3 2 3 2 13 4 9 9 10 13 2
6 13 2 3 13 2 2
6 3 3 13 10 13 2
7 3 13 4 12 9 13 2
9 12 9 10 0 13 9 9 7 2
18 9 13 9 2 9 0 0 9 13 9 13 2 3 9 9 12 13 2
16 9 9 2 11 9 13 9 13 2 13 9 12 9 13 4 2
5 11 9 0 13 2
7 3 2 9 10 13 4 2
6 2 10 13 4 2 2
5 13 4 9 13 2
6 9 12 12 13 4 2
10 3 2 11 12 9 9 0 13 4 2
14 0 13 4 11 11 2 11 11 7 11 11 13 4 2
14 9 12 13 4 2 7 3 9 13 10 9 0 12 2
5 3 9 13 4 2
10 9 9 13 2 9 0 13 4 3 2
10 11 13 11 2 0 2 13 13 11 2
6 13 13 11 9 0 2
4 9 13 10 2
7 7 3 2 9 13 4 2
12 11 13 13 4 2 11 7 9 9 13 13 2
7 9 9 13 9 13 9 2
10 10 13 2 9 2 12 9 13 4 2
10 11 13 4 0 9 9 10 13 4 2
15 9 13 4 3 13 4 3 7 9 9 0 13 4 2 2
20 13 4 9 11 9 13 9 13 13 13 4 2 7 2 3 2 14 4 13 2
20 7 2 11 7 11 9 13 4 2 9 9 10 9 9 12 13 9 9 13 2
8 9 0 9 13 9 13 9 2
7 9 0 13 4 0 9 2
21 11 9 13 10 9 13 7 2 11 9 0 9 13 10 9 7 12 9 13 4 2
10 11 9 0 12 13 4 11 11 9 2
9 9 9 13 4 9 3 7 3 2
19 3 9 13 3 2 9 10 7 9 10 13 4 11 7 11 9 9 10 2
4 9 13 4 2
12 9 9 10 9 13 9 13 4 9 0 9 2
5 11 9 13 4 2
9 14 4 2 3 2 9 12 13 2
12 3 2 9 0 12 13 7 9 13 4 3 2
4 9 9 13 2
15 11 9 13 9 2 9 2 13 4 9 12 9 9 13 2
7 9 10 12 9 13 4 2
11 13 9 0 7 2 7 10 9 0 13 2
6 11 14 4 9 13 2
5 11 13 4 3 2
6 3 9 9 13 0 2
7 9 9 13 9 13 13 2
11 6 2 9 13 9 14 4 9 0 13 2
10 11 7 2 9 10 9 13 13 4 2
6 11 9 13 9 10 2
15 9 0 13 2 13 4 9 9 3 13 4 11 11 9 2
27 14 12 14 12 9 11 7 11 13 0 2 7 3 9 13 9 10 9 13 2 9 9 13 2 12 9 2
9 13 7 15 15 9 13 4 9 2
10 2 13 9 9 13 13 9 13 2 2
13 11 12 9 13 11 2 7 12 9 3 13 4 2
18 12 9 0 9 2 11 11 7 10 9 9 13 9 13 4 2 3 2
4 3 10 13 2
17 13 9 9 0 13 9 13 7 9 3 13 4 2 9 8 3 2
19 9 2 9 9 0 12 13 4 2 9 9 9 9 13 7 9 13 13 2
12 7 2 9 9 13 4 9 13 10 9 13 2
13 11 9 13 4 2 2 9 13 13 4 9 2 2
16 2 9 7 2 14 13 3 0 2 0 13 11 10 9 2 2
28 9 10 9 7 9 13 4 9 10 9 9 9 13 2 9 7 9 9 13 2 9 9 7 9 9 13 2 2
28 2 3 9 14 4 9 13 2 9 11 9 9 0 13 4 2 7 12 9 0 13 4 9 2 2 13 4 2
11 2 15 9 10 9 13 7 13 4 2 2
9 0 9 13 9 13 4 3 9 2
15 9 10 13 2 9 12 13 4 2 7 9 9 13 10 2
8 9 9 11 12 9 13 13 2
5 3 13 4 9 2
5 9 13 2 14 2
11 11 11 0 10 12 9 9 13 4 3 2
6 9 13 4 9 13 2
8 9 9 12 13 4 9 11 2
6 3 13 4 9 0 2
5 3 14 4 13 2
6 9 9 13 9 2 2
14 9 12 13 9 13 3 9 0 9 13 4 9 9 2
18 10 12 9 9 0 13 9 13 2 7 15 14 4 13 9 13 4 2
23 11 14 4 9 0 13 11 2 11 2 3 11 9 4 7 2 10 3 13 9 13 4 2
11 9 12 13 4 2 7 9 13 4 12 2
20 3 2 9 13 10 9 0 11 9 13 13 4 7 10 10 9 0 13 4 2
8 10 9 2 11 11 13 4 2
11 0 9 7 12 11 9 13 4 13 4 2
7 3 13 4 12 9 7 2
15 9 9 0 0 13 9 2 7 9 13 2 9 13 4 2
4 9 0 13 2
6 9 9 13 9 13 2
11 11 9 13 4 2 12 9 13 13 4 2
11 2 9 9 13 4 7 10 9 0 13 2
5 9 10 9 13 2
13 9 2 9 2 9 7 9 2 13 13 4 9 2
8 11 13 2 11 11 13 4 2
17 2 15 13 4 14 13 15 3 0 7 14 13 0 9 2 7 2
6 2 9 3 13 4 2
10 11 11 0 13 12 2 9 0 12 2
5 2 2 13 4 2
7 13 10 9 13 4 13 2
9 9 11 13 9 7 12 9 13 2
6 2 11 9 9 13 2
20 9 10 9 13 7 9 13 9 2 9 13 13 13 7 14 13 11 9 10 2
8 12 9 13 4 9 0 12 2
5 9 9 13 4 2
5 12 9 13 4 2
11 9 9 9 13 4 11 2 10 9 13 2
12 7 2 12 9 9 10 9 0 13 4 2 2
19 3 7 3 13 4 11 9 2 7 13 9 10 12 9 13 2 12 2 2
15 3 13 4 12 12 9 2 11 7 11 2 11 13 4 2
10 12 9 0 9 0 13 4 9 9 2
11 7 2 9 9 9 7 13 4 9 10 2
9 11 11 0 7 13 13 4 9 2
7 10 7 9 13 4 9 2
6 10 10 9 13 9 2
5 3 13 4 9 2
7 10 9 13 4 3 9 2
10 9 9 13 9 9 13 4 11 9 2
12 11 9 13 13 4 2 9 14 4 9 13 2
14 2 14 4 12 9 9 13 9 13 2 13 7 2 2
6 11 13 4 9 9 2
11 12 9 9 11 9 9 0 9 0 13 2
9 9 13 4 10 2 3 9 13 2
10 9 10 12 9 9 7 9 13 4 2
4 13 13 4 2
14 11 9 13 4 7 10 9 9 0 7 9 0 13 2
13 11 9 9 3 0 13 2 7 9 9 13 4 2
22 3 2 11 9 9 13 4 11 11 9 11 9 9 9 12 13 13 4 9 12 9 2
7 14 4 9 12 9 13 2
10 11 12 9 13 4 12 9 13 9 2
9 11 9 9 7 9 13 4 3 2
8 11 9 13 13 13 13 4 2
14 9 3 13 4 2 9 12 2 9 13 13 9 13 2
11 9 13 4 9 0 10 9 9 13 4 2
17 9 13 3 13 9 2 7 2 2 0 2 13 4 13 4 11 2
10 10 11 12 9 13 9 9 13 4 2
19 9 9 10 0 13 2 9 0 14 13 2 9 0 9 13 13 4 9 2
7 10 0 13 13 13 9 2
7 9 13 10 13 2 8 2
9 9 13 2 11 12 9 0 13 2
18 3 2 11 9 2 2 11 9 9 9 13 2 9 7 14 13 2 2
6 3 13 4 9 13 2
7 11 3 13 4 11 9 2
14 9 13 4 2 9 13 13 2 7 9 13 9 13 2
5 6 2 9 13 2
20 2 13 4 9 13 3 2 3 9 13 7 10 13 13 4 2 2 13 11 2
6 2 13 4 11 2 2
4 15 13 4 2
16 11 12 9 13 9 13 2 11 13 4 2 7 12 9 0 2
10 9 10 13 4 9 9 3 13 4 2
17 2 3 9 12 13 9 13 2 15 13 2 7 14 13 10 2 2
6 0 13 7 2 6 2
24 3 2 9 3 13 4 13 4 2 0 4 2 13 13 4 2 9 12 13 7 9 13 4 2
12 9 2 7 2 11 13 4 9 0 2 12 2
12 2 9 10 9 9 9 7 9 0 13 13 2
7 3 2 3 13 9 9 2
7 3 13 4 9 11 9 2
17 15 9 7 0 7 13 4 2 3 2 9 7 9 12 15 9 2
12 0 13 4 9 9 13 2 9 2 13 4 2
18 11 2 11 9 2 9 13 4 9 2 7 9 9 9 0 13 4 2
7 12 9 9 13 13 4 2
7 2 14 13 10 13 4 2
16 15 13 2 15 9 0 13 3 9 13 4 2 12 9 13 2
14 3 2 9 2 15 9 13 4 7 10 9 13 4 2
5 2 3 13 4 2
6 3 9 2 0 13 2
13 9 0 13 4 11 9 2 9 9 13 9 13 2
10 2 9 0 13 13 9 13 4 2 2
7 2 3 3 13 4 2 2
16 12 9 2 9 9 13 4 9 13 9 2 11 9 13 4 2
8 2 11 2 15 15 13 4 2
15 11 14 4 0 13 10 9 2 7 10 9 13 13 4 2
11 12 7 3 11 2 11 2 13 4 9 2
6 9 13 3 13 4 2
11 9 9 13 13 4 2 7 13 13 4 2
21 9 10 13 4 9 9 13 4 2 7 12 9 13 4 11 2 9 0 2 3 2
20 9 13 2 2 9 11 9 13 9 13 2 13 13 9 7 13 9 13 2 2
19 11 9 2 0 9 11 3 13 4 9 9 9 13 13 2 9 13 2 2
19 9 9 9 3 13 4 9 0 7 2 0 2 2 9 9 9 2 9 2
10 2 11 2 0 9 13 2 13 2 2
17 13 4 2 9 0 12 9 13 13 2 9 0 7 9 0 2 2
5 9 9 13 4 2
6 14 4 3 10 13 2
16 11 2 15 10 13 14 4 13 13 4 9 2 9 13 4 2
5 3 11 9 13 2
8 9 9 10 14 13 9 3 2
21 7 2 11 9 3 13 13 4 2 7 11 7 11 9 0 13 13 4 9 10 2
7 9 13 4 9 9 0 2
9 14 13 9 2 9 3 0 13 2
5 2 13 9 13 2
12 3 2 9 0 9 9 0 7 0 13 4 2
12 13 4 12 9 12 2 12 9 9 13 4 2
9 11 9 9 13 4 9 12 9 2
15 9 13 13 4 9 2 3 9 9 13 7 11 13 13 2
11 9 0 12 13 4 9 2 9 13 13 2
9 9 10 13 13 4 3 7 2 2
7 2 15 13 4 3 9 2
4 0 13 4 2
5 12 9 13 4 2
9 9 9 13 7 9 0 13 15 2
7 12 9 13 7 12 9 2
9 10 9 9 9 13 13 13 4 2
9 11 11 0 13 4 9 9 0 2
10 11 9 9 13 4 11 2 9 9 2
11 11 9 13 4 7 12 13 4 12 9 2
11 11 9 13 9 9 0 13 4 13 9 2
5 15 3 13 13 2
26 9 10 0 9 9 13 4 2 7 11 2 11 7 11 13 4 9 9 9 10 0 9 12 13 4 2
9 9 0 13 14 13 10 9 13 2
6 2 10 14 13 9 2
7 2 14 2 14 13 0 2
4 7 13 13 2
7 11 9 10 9 13 4 2
8 11 7 13 13 4 11 9 2
20 9 0 13 4 2 9 2 9 7 2 9 2 9 13 2 14 4 9 13 2
11 12 9 9 13 4 3 11 2 11 2 2
19 11 9 14 4 13 2 11 2 11 2 11 7 11 10 9 12 13 4 2
15 11 9 13 4 2 2 14 13 9 9 9 13 4 2 2
16 3 2 9 9 13 2 9 13 7 9 13 4 2 9 13 2
10 14 4 13 11 9 13 4 7 14 2
18 9 10 9 13 4 11 11 9 11 9 9 9 13 4 9 9 9 2
22 9 13 2 14 13 9 12 9 3 0 13 4 12 9 3 11 13 9 13 14 4 2
14 7 9 10 0 13 9 13 2 9 3 13 7 4 2
9 2 9 9 13 13 4 2 14 2
4 15 13 4 2
5 9 13 4 11 2
6 7 9 0 13 4 2
6 12 9 0 13 4 2
9 3 9 0 9 0 10 13 4 2
7 11 9 13 12 9 13 2
11 11 9 13 13 4 12 9 13 4 9 2
12 9 9 3 7 13 2 0 0 13 4 15 2
20 3 11 13 13 9 13 2 7 13 9 13 2 13 9 9 0 13 9 13 2
4 14 13 0 2
12 9 12 11 12 9 13 4 11 2 11 2 2
12 11 9 0 12 9 13 4 11 2 9 13 2
23 9 10 3 13 4 12 3 11 13 7 10 3 11 13 2 15 9 2 3 13 9 13 2
13 15 8 9 10 13 4 2 7 3 9 0 13 2
6 3 14 13 13 9 2
9 12 0 2 7 2 0 13 4 2
5 10 13 9 10 2
18 9 12 13 13 13 2 7 13 13 4 2 11 11 9 13 9 13 2
11 14 13 9 12 9 13 11 8 9 0 2
35 9 12 2 12 9 13 4 9 9 0 13 9 2 7 9 12 0 12 9 13 13 4 2 11 2 11 11 2 11 2 11 7 11 2 2
14 14 13 15 10 13 2 7 2 9 10 9 13 4 2
6 11 13 4 11 9 2
17 11 9 11 8 11 2 11 9 11 8 11 2 9 9 13 4 2
19 9 9 13 3 2 9 9 9 9 13 13 4 2 0 13 13 9 13 2
5 14 4 9 13 2
7 2 9 9 8 0 13 2
6 11 9 0 13 4 2
10 9 13 14 4 13 13 4 9 10 2
12 9 13 13 4 10 9 9 10 9 13 4 2
8 7 2 9 12 10 13 4 2
8 11 3 13 9 13 4 9 2
17 2 9 10 2 9 0 9 9 0 9 7 2 13 4 9 0 2
16 11 9 13 4 9 10 9 13 4 9 10 13 13 2 3 2
13 0 13 2 7 2 0 13 2 15 14 4 13 2
7 9 9 13 4 2 3 2
27 11 0 13 9 11 13 4 9 13 4 9 13 2 7 3 9 9 13 4 2 8 10 9 12 13 4 2
9 2 3 13 9 9 13 4 2 2
7 10 2 12 13 9 13 2
7 14 4 12 10 3 13 2
8 11 9 0 12 9 13 4 2
6 11 7 9 0 13 2
6 9 9 9 13 4 2
16 2 11 15 9 13 4 9 2 9 12 11 13 4 3 2 2
8 11 2 9 12 9 13 4 2
14 2 9 13 4 13 4 9 2 7 0 3 13 13 2
10 11 3 14 4 13 9 0 9 0 2
13 14 4 0 13 2 0 9 10 13 4 2 3 2
7 7 10 13 13 10 9 2
25 11 9 0 13 2 7 9 0 10 13 4 2 11 11 9 0 12 8 3 10 13 13 4 3 2
10 7 9 0 10 9 0 10 13 4 2
9 12 9 13 7 3 0 9 13 2
5 12 9 13 4 2
6 2 3 2 15 13 2
14 2 11 13 13 3 13 4 9 0 13 4 11 9 2
11 9 9 13 2 0 10 13 4 9 0 2
10 2 11 11 9 3 0 13 4 2 2
12 2 9 13 9 13 4 7 13 13 4 2 2
6 3 2 11 9 13 2
10 9 0 9 9 7 9 13 13 4 2
14 10 11 10 9 13 4 9 2 9 9 10 9 13 2
10 0 13 9 2 11 7 9 10 13 2
16 9 13 4 3 9 0 7 0 14 4 3 9 9 13 7 2
11 7 9 10 10 9 7 9 9 13 4 2
28 15 9 10 2 9 0 13 9 0 13 2 10 13 9 9 2 9 9 2 9 9 7 9 9 0 9 13 2
7 9 0 12 9 13 4 2
8 2 7 9 9 10 13 3 2
8 14 13 10 9 13 4 9 2
11 11 7 9 2 9 9 2 13 4 13 2
7 9 3 0 13 13 4 2
6 9 0 10 13 9 2
16 11 11 11 9 7 11 11 11 11 9 0 11 13 4 3 2
5 9 13 3 11 2
11 13 2 12 2 7 11 7 11 13 4 2
7 2 9 14 13 0 2 2
6 9 9 13 4 3 2
14 11 11 7 11 9 9 9 13 4 2 7 2 11 2
5 10 9 13 10 2
9 9 10 13 4 3 13 4 9 2
5 2 13 2 9 2
5 13 3 13 4 2
16 9 0 9 0 9 12 13 4 9 9 12 9 0 9 13 2
20 11 7 11 9 13 13 13 9 9 9 7 11 14 4 15 9 13 13 4 2
6 9 14 13 13 13 2
8 3 2 10 9 13 13 4 2
10 11 11 9 9 2 9 12 13 4 2
10 2 13 2 13 2 9 0 2 2 2
8 0 2 9 0 13 4 0 2
8 9 13 13 4 2 9 13 2
5 9 13 9 13 2
21 9 9 2 11 9 2 11 9 2 11 11 9 7 11 7 11 11 9 13 4 2
7 13 9 9 13 13 4 2
6 3 13 4 9 3 2
7 9 2 7 2 9 13 2
10 11 9 7 11 11 9 9 13 4 2
7 11 11 11 13 4 9 2
7 9 7 3 13 4 2 2
11 12 12 9 12 9 13 4 12 11 9 2
9 9 10 13 4 9 13 4 9 2
6 9 7 3 13 4 2
8 13 7 9 13 13 4 11 2
9 3 13 9 13 4 13 4 9 2
7 11 11 9 0 13 4 2
14 3 13 4 9 0 13 3 13 4 3 12 9 13 2
8 12 9 10 9 13 4 11 2
9 9 10 13 13 4 9 9 13 2
5 2 9 0 13 2
6 9 13 12 9 13 2
21 13 9 10 11 13 4 2 3 0 2 13 0 7 9 0 13 4 9 13 4 2
7 9 0 14 4 3 13 2
16 7 3 13 4 9 7 13 4 9 13 13 4 9 13 4 2
15 7 2 9 10 2 10 9 9 9 13 13 4 9 13 2
16 7 2 12 9 3 13 3 13 4 11 7 9 13 13 4 2
8 9 0 13 4 9 11 9 2
8 3 0 13 2 9 7 9 2
7 2 0 9 9 14 13 2
7 11 9 13 4 13 13 2
16 9 13 11 7 11 13 0 0 2 7 11 13 14 13 0 2
12 12 9 13 13 7 15 14 4 0 0 13 2
8 11 9 11 9 9 0 13 2
16 7 2 14 4 10 13 7 3 9 9 3 13 9 13 9 2
10 9 13 9 2 10 9 13 4 3 2
8 11 9 9 0 13 4 9 2
16 9 10 9 7 9 9 13 4 2 7 9 7 9 13 13 2
21 11 13 13 2 9 0 2 14 13 13 9 2 0 9 9 13 4 9 13 4 2
10 14 4 2 7 2 9 0 13 9 2
13 11 11 0 9 13 4 3 9 0 0 9 13 2
17 11 11 9 9 12 13 4 9 13 4 2 9 7 9 2 13 2
14 11 11 9 9 13 7 9 0 9 13 13 4 11 2
31 2 9 13 11 2 9 9 9 9 9 9 2 2 7 2 9 13 11 2 7 2 11 2 12 2 2 9 10 9 2 2
13 7 3 10 7 3 7 3 13 4 9 0 10 2
14 11 11 11 13 4 13 9 2 0 0 9 13 3 2
7 9 0 7 0 13 4 2
17 9 3 13 4 13 7 2 9 3 13 2 12 9 9 13 4 2
9 9 10 13 0 13 7 15 14 2
17 11 9 9 13 9 9 9 13 2 9 13 4 10 9 0 13 2
10 9 10 13 2 10 9 13 9 13 2
8 9 13 9 10 10 9 12 2
8 7 2 9 0 11 13 4 2
8 2 11 13 7 13 4 2 2
14 9 10 13 9 13 9 9 0 13 13 4 9 9 2
10 11 7 11 9 10 12 9 13 4 2
14 3 9 3 13 4 2 7 9 7 9 0 13 4 2
8 9 13 13 11 11 8 11 2
4 13 3 13 2
16 9 13 9 2 3 13 4 9 2 0 2 13 4 13 4 2
9 14 13 10 9 11 11 11 9 2
7 9 9 13 9 7 13 2
22 9 9 13 4 9 9 10 2 7 9 13 4 9 2 9 2 3 13 4 10 9 2
13 2 12 2 12 9 12 13 9 13 4 11 9 2
8 0 9 3 13 9 13 9 2
4 10 13 4 2
8 2 9 10 0 13 4 3 2
9 11 7 11 13 7 9 13 4 2
19 7 2 2 12 9 13 9 0 8 9 0 13 9 0 9 2 11 9 2
20 11 11 11 9 12 9 9 0 13 4 2 7 12 9 9 0 7 13 4 2
15 14 13 13 11 3 13 2 10 9 0 13 3 3 13 2
13 9 9 2 7 9 13 9 11 13 4 9 9 2
10 3 7 0 13 4 12 12 9 9 2
11 12 9 9 2 9 2 11 9 12 13 2
15 11 2 7 2 9 12 9 13 3 2 3 3 13 4 2
8 3 2 11 12 9 12 13 2
9 3 12 9 13 4 9 13 9 2
5 14 13 9 7 2
9 9 13 9 2 10 9 12 13 2
10 2 9 9 12 9 9 12 13 2 2
13 9 13 9 2 9 7 2 11 11 10 13 9 2
7 7 2 9 9 13 4 2
15 3 14 4 9 12 13 9 13 2 7 9 13 9 13 2
10 10 2 3 9 10 9 10 13 4 2
19 9 9 13 4 11 9 2 7 12 9 0 9 13 4 11 9 0 13 2
4 13 13 4 2
20 0 9 3 0 13 4 2 7 9 3 3 13 7 2 13 9 10 13 3 2
8 9 0 9 13 11 13 4 2
4 9 13 13 2
12 9 9 9 12 9 9 13 4 11 9 9 2
10 2 9 9 0 13 4 9 4 2 2
8 9 12 14 4 9 13 13 2
11 3 2 11 10 9 12 9 13 13 4 2
7 9 0 13 9 13 13 2
10 2 9 10 3 7 13 4 2 11 2
13 9 0 9 9 9 13 4 2 11 13 13 4 2
9 2 11 9 9 0 12 13 4 2
11 7 9 13 13 4 9 0 10 13 4 2
18 2 9 9 12 13 4 2 7 2 7 2 9 9 13 13 4 2 2
13 3 3 13 11 9 12 9 9 11 7 11 11 2
4 9 13 4 2
4 2 3 13 2
14 11 9 0 13 2 7 10 9 10 0 13 9 13 2
9 2 12 9 9 12 13 13 2 2
17 9 0 9 12 13 4 2 9 9 7 9 12 12 9 0 13 2
4 9 13 4 2
8 11 0 9 13 4 11 9 2
8 7 3 13 15 12 9 4 2
7 9 9 7 3 13 4 2
12 9 7 9 0 3 13 9 10 10 9 13 2
9 9 2 9 2 7 13 13 4 2
12 11 9 13 9 9 10 13 4 13 13 4 2
12 11 12 9 13 2 7 0 13 9 13 4 2
10 9 9 11 7 11 0 9 13 4 2
23 3 0 13 4 9 2 7 9 13 4 2 7 9 0 7 9 7 9 13 4 9 13 2
17 3 2 9 13 4 11 2 2 0 9 0 13 9 0 13 2 2
17 3 13 4 12 9 2 7 9 0 14 4 13 12 12 9 10 2
16 11 14 4 3 13 2 7 0 9 12 13 4 11 11 9 2
11 9 2 7 2 9 13 9 0 13 11 2
21 9 12 5 9 13 7 9 13 4 12 9 13 13 2 7 9 9 13 8 4 2
9 7 9 13 2 9 9 13 4 2
15 9 0 13 3 13 4 2 9 10 3 13 15 0 13 2
6 14 13 9 2 11 2
13 2 9 11 13 4 2 9 2 9 7 9 2 2
6 0 9 14 13 9 2
9 0 13 7 9 7 9 3 13 2
13 10 13 9 13 9 0 13 4 9 11 13 9 2
5 14 4 13 13 2
4 11 13 4 2
12 9 9 0 7 0 0 13 4 11 9 0 2
17 9 7 13 13 4 9 2 14 4 9 10 15 9 13 2 13 2
21 9 9 9 13 4 7 14 4 13 2 13 4 9 13 9 0 9 13 4 13 2
7 11 7 9 9 9 13 2
8 11 11 13 9 13 9 13 2
11 3 9 13 4 11 2 10 9 10 12 2
13 9 12 9 13 9 9 12 9 13 11 9 0 2
9 6 6 11 0 13 13 2 10 2
29 14 4 9 0 13 9 2 7 3 9 13 9 12 9 12 2 7 13 4 9 0 13 0 13 14 13 10 13 2
20 12 9 15 9 9 13 7 13 4 9 0 13 4 2 3 13 4 9 13 2
13 7 2 0 11 7 2 11 2 13 9 2 12 2
8 2 13 9 9 13 4 9 2
14 9 11 9 13 7 9 12 9 13 4 2 9 9 2
9 11 9 9 14 4 13 3 7 2
13 12 9 12 9 13 4 11 2 3 9 13 4 2
8 14 4 9 0 13 9 10 2
8 3 7 11 9 13 13 4 2
24 11 11 7 11 11 9 7 13 4 3 13 4 15 9 9 7 9 10 15 9 9 13 13 2
6 12 9 13 4 9 2
13 13 9 2 11 2 9 9 13 4 12 9 0 2
14 12 7 12 13 4 11 2 7 11 13 4 11 9 2
14 11 3 13 4 12 9 13 2 9 0 2 13 4 2
17 11 13 3 9 2 7 3 9 13 9 13 2 14 4 9 13 2
10 11 13 4 9 10 2 9 13 3 2
13 13 13 4 9 2 7 13 9 14 13 15 9 2
14 2 11 9 9 0 11 13 4 9 9 9 13 2 2
6 3 12 9 13 9 2
9 13 4 9 10 14 4 13 11 2
9 13 11 9 13 4 9 2 3 2
11 3 13 2 11 7 0 9 10 13 4 2
22 3 2 11 9 13 13 4 9 0 2 11 9 2 9 13 4 13 0 13 4 9 2
12 3 9 13 9 0 2 0 7 9 9 13 2
7 7 11 3 13 4 11 2
12 3 2 11 7 11 9 13 9 13 13 4 2
9 9 9 0 3 9 0 13 4 2
13 7 2 2 9 9 9 0 14 4 3 13 2 2
13 9 9 3 13 4 11 13 9 0 11 9 13 2
13 11 12 9 13 4 3 2 7 3 13 9 13 2
8 3 9 10 13 4 12 9 2
8 11 12 9 13 4 13 9 2
6 2 14 13 2 9 2
17 9 10 2 3 9 13 4 9 0 2 3 13 4 3 12 9 2
3 3 13 2
16 9 0 3 9 13 4 2 11 9 9 9 13 4 11 9 2
7 9 0 13 13 9 13 2
7 7 10 9 10 13 4 2
16 12 9 9 13 4 9 9 9 7 9 10 9 0 13 4 2
4 9 9 13 2
14 11 13 13 7 9 9 9 13 9 13 13 4 11 2
5 15 12 13 13 2
4 3 9 13 2
14 10 9 3 9 10 13 4 9 7 9 13 9 13 2
8 0 9 12 9 0 13 13 2
16 12 9 14 4 13 13 9 2 7 9 9 13 9 13 4 2
19 11 2 7 2 11 9 14 4 13 13 2 7 9 10 9 9 13 4 2
5 9 3 13 13 2
8 11 11 0 13 4 9 0 2
12 3 2 11 2 11 7 11 13 13 13 13 2
15 9 10 9 13 13 4 2 7 14 4 13 9 9 13 2
13 9 7 0 12 9 2 7 2 12 9 13 4 2
8 3 2 11 9 13 4 13 2
4 9 13 4 2
7 11 11 9 9 9 13 2
10 11 11 11 12 3 9 12 13 4 2
8 9 9 13 4 9 13 4 2
12 11 13 13 4 2 9 13 7 13 13 4 2
6 11 12 9 13 4 2
11 13 9 9 3 12 9 13 4 13 4 2
6 13 11 9 11 13 2
7 3 13 4 3 11 9 2
28 9 13 9 7 11 2 0 9 2 13 9 14 13 13 4 11 11 11 11 2 2 3 3 3 13 4 2 2
7 13 13 7 9 9 13 2
6 2 0 13 4 9 2
9 9 9 2 11 14 4 13 3 2
9 9 12 13 4 9 2 9 11 2
9 3 2 7 2 14 13 9 0 2
14 9 13 2 13 7 13 9 2 15 9 9 13 4 2
10 2 13 9 2 11 9 13 4 11 2
13 9 9 12 9 10 13 4 9 0 9 13 4 2
13 9 0 3 13 4 9 2 7 9 13 4 9 2
15 9 0 13 4 9 2 13 4 9 13 7 10 3 13 2
14 2 15 9 9 13 9 0 13 7 0 13 13 4 2
23 7 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 7 11 13 4 9 2
6 9 3 13 4 12 2
7 11 11 13 4 10 12 2
5 9 0 13 11 2
10 15 14 13 0 13 2 3 13 7 2
6 3 2 12 9 13 2
27 2 9 9 9 13 4 9 7 9 10 13 9 13 4 2 7 10 3 13 4 3 13 13 9 13 2 2
10 11 11 9 9 0 13 4 3 9 2
14 15 3 13 4 2 0 13 4 9 10 13 9 13 2
4 12 9 13 2
5 2 3 13 4 2
9 11 11 9 14 4 9 10 13 2
18 9 9 2 9 7 9 2 9 4 9 10 3 13 13 4 9 11 2
6 2 9 11 13 4 2
7 0 9 13 11 7 11 2
20 3 2 11 9 11 11 9 0 13 13 2 9 11 9 0 12 13 13 4 2
11 11 2 9 13 2 14 4 13 13 4 2
7 3 13 4 2 9 13 2
10 9 13 13 4 2 9 9 3 13 2
8 3 14 13 3 3 13 4 2
13 11 9 12 13 4 2 9 9 9 10 13 9 2
9 7 2 3 13 4 11 13 9 2
5 11 12 9 13 2
20 9 9 7 9 9 9 9 13 2 7 7 0 9 12 2 0 9 10 13 2
7 2 11 3 13 4 7 2
17 3 2 11 11 8 11 7 11 11 9 9 13 4 3 9 10 2
10 0 9 10 9 3 13 4 2 3 2
9 2 10 13 2 11 3 13 4 2
5 11 9 0 13 2
10 11 9 12 9 13 4 11 11 9 2
5 3 13 9 0 2
15 9 9 0 11 13 9 9 9 12 13 4 12 12 9 2
16 9 7 9 0 13 4 9 13 13 4 9 9 0 13 4 2
24 9 10 2 9 2 2 9 13 7 2 9 2 0 12 13 4 9 13 2 7 9 2 14 2
7 9 0 10 13 13 4 2
13 9 9 9 0 0 9 13 2 9 12 9 13 2
13 10 9 9 9 13 9 13 2 14 13 0 2 2
7 13 4 14 4 9 13 2
9 12 12 9 3 13 4 9 13 2
10 2 9 14 13 0 2 2 13 4 2
18 7 2 14 4 3 0 13 2 7 10 13 9 13 9 9 12 13 2
15 2 13 4 2 7 9 12 9 13 2 13 13 13 4 2
8 7 11 14 13 11 13 9 2
5 11 13 13 4 2
16 13 13 4 11 13 13 4 12 10 12 11 9 13 13 4 2
9 3 9 13 7 9 12 13 4 2
12 13 14 13 9 10 13 4 9 0 13 4 2
8 2 9 13 4 9 13 4 2
5 7 3 13 4 2
5 10 13 4 3 2
16 9 12 12 9 9 9 13 0 4 11 11 9 0 12 9 2
8 0 13 0 9 13 9 13 2
20 0 9 9 13 4 2 7 2 11 9 9 2 9 7 9 2 13 9 4 2
14 2 9 3 13 4 7 3 2 9 9 13 13 2 2
19 3 13 4 11 11 12 9 2 7 3 9 9 13 4 12 9 9 0 2
19 9 2 7 2 14 13 2 9 9 9 2 9 9 10 13 4 3 9 2
5 10 9 13 4 2
13 10 9 13 9 2 7 13 9 0 9 13 4 2
13 11 9 9 9 10 13 4 11 9 9 13 9 2
14 15 13 13 9 13 2 7 0 13 9 7 9 13 2
7 3 2 12 9 13 11 2
12 10 2 9 14 13 9 2 7 13 13 13 2
17 9 0 9 9 12 13 4 2 7 9 9 10 13 4 13 4 2
5 9 13 13 4 2
25 9 10 13 2 2 9 10 10 10 9 9 13 2 3 7 9 9 2 9 13 0 13 4 2 2
12 11 9 13 4 9 13 9 2 11 7 3 2
5 7 14 4 13 2
10 10 0 13 7 9 0 9 13 4 2
8 2 0 13 7 9 13 4 2
6 7 9 13 10 9 2
12 9 13 13 4 7 3 10 12 9 13 4 2
8 10 13 4 9 9 9 9 2
10 11 7 11 3 9 0 13 4 13 2
9 11 11 9 0 7 13 4 13 2
7 9 13 4 9 3 13 2
7 14 4 15 9 9 13 2
12 3 2 7 2 9 9 13 4 2 9 9 2
6 3 9 0 13 4 2
6 9 0 13 4 11 2
15 9 2 7 2 3 9 0 13 11 2 7 9 13 4 2
8 11 9 0 13 4 3 11 2
10 9 0 7 0 13 4 3 9 0 2
7 2 3 3 13 13 4 2
16 7 3 9 0 13 4 11 12 9 2 7 11 9 12 2 2
7 11 0 9 13 4 9 2
9 2 9 13 9 11 9 13 4 2
10 9 13 2 9 10 2 9 0 0 2
25 3 11 13 9 13 4 3 2 11 9 9 13 9 9 9 13 9 13 7 9 14 4 9 13 2
18 9 10 3 12 9 9 2 12 9 2 13 4 11 10 9 12 9 2
7 11 0 13 4 9 0 2
7 9 13 13 4 10 10 2
4 3 13 10 2
13 2 9 10 13 4 11 13 7 3 9 13 4 2
28 11 9 9 13 4 11 11 9 9 2 12 2 2 11 9 2 12 2 7 11 7 9 13 11 2 12 2 2
6 9 12 13 4 9 2
12 11 13 9 12 9 13 11 13 9 13 9 2
24 11 11 9 9 10 9 13 9 13 2 3 2 7 2 13 7 13 4 2 12 9 13 4 2
14 0 13 3 2 9 13 4 9 7 9 10 10 13 2
28 11 11 9 9 9 2 11 9 13 2 13 13 4 7 11 9 13 4 9 14 13 11 2 9 2 13 4 2
5 9 3 13 4 2
14 9 2 14 4 0 13 9 10 13 4 9 0 9 2
14 3 9 12 12 9 13 4 12 2 7 9 13 4 2
6 13 3 9 0 10 2
11 2 9 9 9 9 13 7 13 13 4 2
7 2 3 13 13 4 2 2
13 0 9 13 13 4 3 11 12 9 2 12 2 2
13 9 9 13 7 0 9 0 13 13 4 9 10 2
7 0 13 9 7 9 13 2
11 11 9 9 9 0 3 13 4 9 10 2
17 11 9 2 7 2 9 9 0 13 4 9 9 13 2 12 9 2
20 11 2 10 9 2 0 9 0 13 4 2 7 2 3 2 3 9 0 13 2
7 3 13 11 9 9 9 2
19 11 14 4 9 13 2 7 9 14 4 13 2 7 9 9 0 13 4 2
4 9 9 13 2
12 7 9 10 13 4 11 11 9 0 13 2 2
7 3 2 12 13 4 9 2
11 12 9 9 9 13 4 12 9 9 13 2
11 7 15 9 13 4 9 13 13 0 4 2
25 13 9 13 9 9 0 13 3 2 9 0 9 0 13 4 7 2 9 2 9 2 12 9 2 2
14 9 0 3 13 4 11 9 11 9 14 13 13 9 2
10 2 3 10 11 11 3 13 13 2 2
9 9 9 2 12 2 9 9 13 2
8 2 9 13 13 9 13 2 2
15 2 14 4 9 13 9 2 9 2 9 7 9 13 7 2
9 9 10 7 9 0 9 13 4 2
15 9 7 9 0 3 13 13 9 13 2 9 9 0 13 2
9 11 9 13 4 9 9 13 4 2
10 9 0 13 7 11 13 13 9 9 2
9 11 2 12 9 9 9 13 4 2
10 13 11 11 13 11 9 11 11 9 2
13 7 11 14 4 9 2 9 0 13 9 12 8 2
6 14 4 9 13 2 2
5 14 4 10 13 2
9 9 9 0 9 13 2 9 2 2
7 2 14 4 9 0 13 2
10 0 10 11 9 7 9 9 9 13 2
9 9 13 2 9 13 14 4 13 2
10 3 13 3 2 9 9 9 13 4 2
9 11 9 13 4 2 9 13 13 2
18 9 14 4 13 2 9 12 13 4 11 9 7 9 9 9 14 13 2
8 9 9 9 9 0 13 4 2
8 3 9 13 4 9 13 9 2
17 7 12 9 9 9 13 4 2 11 11 11 14 4 2 7 13 2
20 9 11 13 15 9 13 9 0 2 3 14 4 13 10 13 10 9 11 9 2
6 2 10 13 4 3 2
14 13 4 0 9 0 7 0 7 13 4 0 9 12 2
5 3 13 13 15 2
15 9 10 2 15 0 13 13 4 9 2 13 2 0 13 2
10 12 9 13 4 0 9 13 9 9 2
7 0 9 9 0 13 4 2
11 9 0 9 13 4 7 9 12 13 4 2
9 13 4 3 9 13 4 12 9 2
6 10 7 15 13 4 2
12 9 0 9 12 13 4 9 12 13 13 4 2
7 2 3 3 13 2 14 2
9 11 9 12 13 9 13 4 9 2
5 3 13 4 9 2
5 9 9 12 13 2
8 11 9 9 14 4 3 13 2
9 10 9 13 9 13 4 9 9 2
17 2 9 7 9 2 9 3 13 4 2 3 0 13 10 13 2 2
3 9 13 2
9 7 9 2 9 7 9 13 4 2
12 12 10 2 9 9 9 0 13 4 11 9 2
8 2 9 13 4 9 13 2 2
14 9 10 2 12 9 11 13 4 9 11 13 13 4 2
10 11 9 10 7 9 13 4 9 13 2
14 12 9 13 4 9 0 12 2 3 12 9 13 4 2
31 3 2 11 9 7 9 10 7 12 13 4 9 2 13 4 12 9 9 12 15 9 13 3 2 2 7 9 13 13 4 2
6 9 9 0 13 4 2
9 11 2 11 2 9 0 13 15 2
20 12 9 12 9 9 13 7 10 13 4 9 2 7 9 0 9 10 13 4 2
15 9 3 13 4 3 2 7 3 3 0 13 0 9 13 2
19 9 13 7 2 7 2 11 9 13 4 9 9 13 4 9 7 11 9 2
17 12 9 9 0 9 9 7 9 9 2 0 9 2 13 9 13 2
13 9 0 7 0 13 7 3 9 9 12 13 4 2
15 11 9 13 13 4 11 14 13 3 2 7 3 3 13 2
5 9 13 13 9 2
10 3 12 9 13 4 2 12 9 2 2
17 11 9 9 10 13 4 2 7 9 7 9 10 0 9 13 4 2
13 9 10 13 4 2 7 2 11 9 0 12 9 2
24 11 9 9 12 9 13 4 12 9 9 13 4 2 7 0 11 13 4 9 2 9 7 9 2
8 11 11 9 13 4 3 11 2
7 12 9 0 13 4 11 2
18 9 0 9 13 7 2 10 0 13 9 0 10 9 13 4 12 9 2
26 9 9 9 13 13 9 10 11 2 7 15 9 9 12 9 13 3 2 9 9 0 13 4 13 4 2
14 2 9 3 13 4 13 4 7 10 3 13 4 2 2
21 11 9 9 12 9 9 12 13 4 2 11 11 12 9 9 13 7 13 0 13 2
13 7 2 9 9 9 9 13 14 13 13 4 9 2
11 9 9 9 9 9 9 9 9 13 4 2
8 9 12 13 4 11 2 9 2
10 9 12 7 13 4 2 9 9 9 2
7 7 2 13 9 10 13 2
10 9 10 2 11 9 13 4 11 9 2
11 7 11 13 13 4 11 9 10 13 4 2
10 9 13 4 2 9 3 13 13 4 2
6 2 13 4 9 2 2
8 11 7 9 10 13 4 3 2
11 11 14 4 13 11 11 13 4 9 0 2
12 3 9 13 7 13 13 9 10 9 13 4 2
9 9 0 10 9 10 13 13 3 2
14 11 13 2 9 9 9 13 4 9 12 9 13 2 2
9 9 10 7 12 9 13 4 9 2
6 3 9 13 13 4 2
7 9 3 12 9 13 4 2
10 9 2 11 9 0 13 4 10 9 2
17 11 9 0 9 0 13 3 2 7 10 9 10 9 0 13 4 2
5 13 13 4 10 2
6 2 0 9 13 2 2
31 9 13 9 2 9 9 13 3 2 9 13 13 4 2 10 2 9 12 2 12 7 10 13 4 2 13 4 9 9 13 2
18 9 11 9 13 4 2 7 2 9 3 13 2 3 9 9 13 4 2
16 11 9 9 7 9 9 2 9 0 9 2 13 13 4 11 2
8 9 13 9 13 7 9 13 2
13 9 2 9 2 9 7 9 9 13 4 9 10 2
15 2 11 9 10 9 13 4 9 0 9 12 13 13 4 2
21 12 9 9 13 4 11 9 10 9 2 7 9 0 10 9 9 13 13 4 9 2
15 11 2 11 7 11 9 7 9 9 9 13 4 3 11 2
10 9 7 9 11 9 0 0 13 4 2
23 9 7 9 13 9 13 4 9 12 9 7 13 8 10 13 7 13 4 3 13 4 9 2
14 9 13 3 2 13 13 4 2 9 9 13 14 4 2
13 2 9 0 13 7 2 15 9 9 13 10 2 2
6 15 13 3 2 9 2
12 11 9 3 13 4 9 9 9 13 9 0 2
11 13 4 9 0 7 0 9 0 13 4 2
9 3 7 3 13 4 13 9 13 2
11 9 0 9 13 13 4 9 9 0 0 2
8 9 0 2 9 9 13 4 2
12 9 13 14 4 13 2 7 14 4 9 13 2
12 9 9 9 12 13 4 2 14 4 3 13 2
6 9 10 3 9 13 2
11 12 9 13 4 9 11 8 11 9 0 2
8 3 7 9 3 13 4 9 2
9 11 7 11 9 0 13 4 12 2
4 10 13 4 2
21 3 12 9 13 2 7 0 9 13 9 13 9 13 2 9 13 9 13 2 7 2
8 2 0 13 3 0 13 11 2
15 3 2 9 9 0 12 13 4 2 7 14 4 9 13 2
5 9 0 13 4 2
9 10 13 4 9 9 9 0 12 2
11 11 2 7 2 12 13 4 7 11 12 2
7 9 9 14 4 0 13 2
5 9 13 13 4 2
9 9 13 7 7 9 13 9 13 2
27 0 13 9 13 14 4 9 10 3 13 2 7 2 3 13 4 13 7 13 4 9 0 13 13 13 13 2
11 10 13 2 7 2 9 2 9 9 9 2
6 15 9 9 0 13 2
24 10 2 9 10 9 9 2 13 9 13 4 2 7 9 2 9 7 9 0 9 13 13 4 2
6 9 0 12 13 4 2
14 6 2 9 13 9 13 10 13 2 7 13 9 13 2
15 9 2 11 2 11 0 13 9 13 2 2 13 4 11 2
6 0 9 0 13 9 2
6 12 12 9 13 4 2
13 9 13 13 7 2 11 11 13 9 3 13 9 2
6 10 12 11 13 4 2
14 11 9 13 9 9 11 11 13 4 13 4 13 4 2
4 2 9 13 2
11 9 9 2 11 10 9 12 13 4 9 2
9 9 3 9 9 13 4 9 9 2
10 2 9 13 7 9 9 13 13 4 2
7 9 9 9 13 13 9 2
9 11 11 13 9 9 9 13 9 2
7 11 14 4 9 11 13 2
8 11 9 9 0 13 4 11 2
7 0 12 13 4 9 9 2
11 9 10 13 7 2 14 4 0 13 11 2
17 11 11 7 11 11 9 9 0 13 4 7 11 11 9 13 4 2
4 15 14 13 2
23 9 0 9 13 2 9 13 4 7 9 13 2 3 9 0 13 4 3 9 0 13 13 2
14 9 13 9 13 9 0 10 2 3 0 13 0 9 2
9 7 2 13 13 9 12 9 0 2
10 9 9 9 14 4 2 7 2 13 2
11 9 10 9 13 3 12 9 9 13 4 2
12 13 0 13 9 13 2 7 9 12 13 9 2
11 12 12 9 9 10 13 4 11 7 9 2
14 9 0 13 4 9 2 7 13 9 0 9 7 13 2
11 12 9 13 4 2 11 13 9 13 13 2
13 11 9 13 4 9 13 13 4 9 9 10 9 2
10 12 9 2 7 2 3 13 9 0 2
15 11 13 4 3 2 9 14 4 9 0 9 13 10 9 2
14 2 15 9 0 11 9 13 2 7 12 9 13 2 2
9 12 9 13 4 9 12 13 13 2
9 10 12 9 9 9 13 9 9 2
6 7 3 14 13 9 2
11 14 13 7 2 11 9 0 13 4 9 2
20 9 2 9 2 9 2 9 7 9 9 9 9 13 13 7 13 13 9 9 2
7 11 9 11 9 13 4 2
5 9 9 0 13 2
29 11 9 2 11 2 12 9 9 9 11 2 11 2 11 2 13 4 3 7 3 2 9 9 9 9 13 9 13 2
10 3 2 9 12 9 12 13 9 9 2
9 13 3 12 9 9 9 13 4 2
17 9 9 13 4 12 9 13 4 3 7 11 3 14 4 9 13 2
20 11 2 11 2 11 7 11 7 14 4 13 2 11 7 11 14 4 13 3 2
6 11 9 0 13 10 2
25 11 9 13 9 13 4 2 7 11 8 11 13 14 4 2 13 4 3 13 9 2 9 10 13 2
9 11 9 0 9 0 12 13 3 2
5 9 14 13 4 2
14 11 12 9 9 9 13 4 11 9 9 9 9 13 2
11 2 11 9 11 9 0 13 13 4 9 2
10 0 12 2 12 7 12 9 13 4 2
6 13 13 9 13 2 2
24 11 13 9 9 13 4 13 11 2 7 9 13 7 9 13 4 9 9 9 0 13 13 4 2
6 12 9 13 4 0 2
7 2 10 13 4 2 11 2
14 9 0 7 0 13 13 4 9 2 13 9 9 2 2
4 9 0 13 2
12 9 0 13 4 11 9 2 9 3 13 4 2
10 3 10 9 13 4 9 9 2 3 2
20 11 11 9 0 7 11 11 0 0 9 9 0 13 0 13 13 9 13 4 2
6 9 14 13 9 9 2
12 12 9 9 13 3 2 9 13 4 9 10 2
8 2 3 9 9 14 13 9 2
7 9 12 12 13 4 3 2
11 11 9 13 13 4 12 9 9 2 11 2
17 9 9 9 7 9 7 9 13 7 9 2 13 13 4 9 13 2
17 13 9 12 9 2 13 13 4 2 7 9 13 7 13 13 4 2
19 13 9 3 13 4 9 13 2 7 9 10 13 9 13 4 2 0 13 2
5 11 12 13 4 2
11 9 10 11 13 4 7 15 13 4 9 2
4 0 13 10 2
10 9 11 9 9 13 7 9 13 4 2
15 0 2 12 9 0 9 13 3 2 9 13 4 2 9 2
12 7 9 10 9 13 2 9 3 13 13 4 2
14 11 11 13 4 9 0 2 7 14 4 9 13 13 2
17 9 0 13 2 9 9 7 9 0 0 2 9 0 7 3 13 2
14 9 9 9 13 7 14 13 13 4 9 10 9 0 2
4 12 13 4 2
6 15 13 3 2 11 2
6 9 13 13 4 9 2
15 11 11 3 13 4 12 9 9 2 7 9 0 13 3 2
5 9 0 13 4 2
7 2 9 9 0 14 13 2
16 9 9 2 0 10 9 7 9 10 2 3 13 4 0 9 2
15 2 7 2 3 14 13 2 3 13 4 9 9 3 13 2
8 11 9 11 7 11 13 13 2
14 11 11 0 12 9 13 4 9 2 7 12 9 9 2
13 9 0 11 9 13 2 7 3 13 4 12 9 2
17 3 9 13 4 7 12 9 13 4 9 9 2 9 7 13 13 2
4 9 13 4 2
4 3 3 13 2
16 15 14 13 9 9 13 7 9 15 14 4 13 7 13 2 2
6 12 9 13 4 9 2
30 9 9 12 13 4 2 9 9 13 4 7 3 13 12 9 7 10 9 9 12 2 9 12 7 9 12 9 13 4 2
7 12 9 9 13 9 9 2
7 10 2 7 2 13 13 2
9 9 13 12 2 13 7 13 0 2
23 11 9 2 3 2 13 4 11 14 4 9 13 7 2 10 9 13 2 9 13 13 4 2
8 10 13 2 13 13 4 3 2
10 9 3 13 4 2 7 3 13 2 2
6 2 9 14 13 0 2
13 9 9 9 2 9 2 9 7 9 9 13 4 2
16 11 0 13 9 0 2 7 9 13 4 10 13 4 11 9 2
18 12 9 11 9 0 13 4 11 0 2 7 9 9 9 13 4 10 2
11 9 12 9 13 7 3 13 4 9 0 2
9 2 9 9 13 13 15 9 2 2
14 11 11 13 0 4 2 10 9 14 4 0 3 13 2
8 0 2 14 4 0 9 13 2
11 9 0 13 2 9 7 0 13 9 13 2
11 11 13 9 0 9 0 13 4 11 9 2
14 9 9 2 7 2 12 9 9 13 4 3 9 9 2
7 3 2 12 13 4 11 2
9 9 9 9 12 13 4 2 3 2
17 12 11 2 9 9 0 13 2 3 13 4 9 9 2 12 5 2
6 13 3 9 12 13 2
22 11 9 13 13 4 11 11 11 2 7 10 13 4 9 14 13 2 9 13 2 4 2
8 3 13 4 11 11 9 11 2
7 9 2 11 13 4 0 2
6 9 12 9 13 4 2
17 0 9 9 2 11 2 11 2 11 2 11 7 11 13 4 0 2
11 9 0 13 4 3 7 3 14 13 9 2
3 9 13 2
12 9 0 13 7 2 12 9 13 9 13 4 2
8 9 0 10 13 4 3 9 2
7 9 12 9 13 4 11 2
16 12 9 11 2 9 8 11 2 0 10 13 4 9 13 9 2
4 9 10 13 2
14 3 2 0 9 13 4 9 9 13 2 13 7 13 2
9 9 9 7 14 9 3 13 4 2
14 10 9 13 4 11 9 13 2 11 11 11 9 13 2
8 7 10 10 9 13 4 2 2
5 2 9 13 4 2
7 2 15 13 13 4 3 2
11 11 9 12 9 9 0 13 4 3 9 2
12 3 13 13 2 7 15 9 9 0 13 13 2
10 7 2 14 4 13 3 0 9 13 2
8 3 2 3 9 13 4 11 2
13 9 13 0 13 11 2 9 0 7 9 3 13 2
12 13 4 13 4 2 7 3 2 0 13 4 2
5 14 13 10 13 2
6 12 9 12 13 4 2
27 10 3 3 13 3 13 4 2 7 13 9 10 3 13 9 13 2 10 13 4 2 7 13 13 4 2 2
8 2 9 9 13 9 13 2 2
11 9 0 13 9 13 2 9 7 9 13 2
10 9 0 13 2 3 14 13 3 0 2
9 9 9 0 2 7 2 10 13 2
9 3 13 9 13 2 3 13 4 2
11 10 13 4 10 9 15 13 7 13 4 2
7 14 4 13 9 13 4 2
8 11 9 10 12 9 13 4 2
18 12 9 10 9 0 0 3 13 4 2 0 0 9 13 9 13 4 2
4 13 9 9 2
6 3 10 10 13 4 2
9 3 2 9 12 11 13 9 13 2
19 7 2 9 13 13 4 2 14 4 3 13 2 10 14 13 10 3 0 2
21 9 9 13 0 9 12 13 4 2 9 10 12 7 11 12 9 13 4 13 4 2
5 14 13 9 11 2
9 2 9 0 3 13 4 2 9 2
4 0 13 9 2
7 13 13 9 9 14 13 2
19 7 9 10 2 10 9 2 3 13 4 11 7 11 2 9 9 2 13 2
11 7 3 13 9 7 13 13 4 7 13 2
4 13 13 4 2
11 11 14 4 13 2 7 3 9 13 4 2
23 9 0 13 4 2 7 11 8 11 9 7 11 11 9 9 13 14 7 2 13 13 4 2
6 2 10 9 13 4 2
3 9 13 2
9 9 12 9 12 9 13 4 3 2
12 9 9 2 12 9 12 9 13 4 13 4 2
15 11 9 7 2 9 9 11 11 0 13 4 0 12 9 2
8 3 0 13 4 2 9 13 2
7 3 13 4 9 0 9 2
5 13 9 13 0 2
10 12 9 11 13 4 2 9 0 12 2
31 0 9 14 13 13 3 2 11 9 9 14 4 0 13 13 4 9 0 9 2 2 9 0 12 0 9 9 13 4 2 2
26 9 13 9 9 10 13 9 13 4 2 9 2 9 0 2 9 9 2 10 9 13 9 9 9 13 2
10 9 13 9 9 0 7 0 13 4 2
7 0 7 10 9 13 3 2
7 15 14 13 10 9 9 2
19 11 11 3 13 4 11 2 7 9 0 13 4 2 13 2 13 4 11 2
8 0 9 2 9 0 13 4 2
11 11 13 9 13 4 9 7 3 13 4 2
7 10 9 13 7 13 4 2
11 7 9 9 13 14 4 2 13 13 4 2
17 3 2 12 9 10 13 4 2 9 13 7 9 9 13 4 9 2
5 9 9 13 0 2
9 7 10 14 4 3 0 13 9 2
18 11 0 2 11 2 11 9 9 13 4 9 2 9 3 13 14 13 2
8 15 9 9 10 9 13 4 2
12 11 9 7 9 9 9 13 4 12 12 9 2
13 15 2 7 2 13 10 10 7 3 13 4 9 2
5 9 13 4 7 2
13 2 9 9 10 13 4 7 2 9 13 9 2 2
10 9 13 13 13 2 11 9 13 4 2
4 10 13 9 2
7 9 12 9 0 13 4 2
12 11 7 10 13 13 13 4 9 9 13 4 2
15 0 9 0 13 4 9 9 9 2 7 3 13 4 9 2
13 13 4 9 13 4 11 2 9 13 4 12 9 2
20 3 13 4 2 10 2 9 2 11 9 13 4 2 9 13 10 9 13 4 2
6 10 9 13 3 13 2
7 11 11 0 7 9 13 2
6 11 9 7 9 13 2
10 9 7 9 2 9 0 2 13 4 2
10 9 9 13 9 13 4 0 9 9 2
6 9 13 4 13 3 2
11 9 9 13 4 11 2 9 13 0 13 2
16 3 7 11 13 4 2 7 12 9 7 12 9 9 13 4 2
8 9 12 13 4 11 9 9 2
15 11 11 0 9 9 7 11 11 0 13 4 11 9 0 2
7 12 0 12 13 4 9 2
16 9 10 2 9 0 13 4 9 2 9 11 7 11 10 13 2
9 11 13 13 2 11 7 11 3 2
8 11 3 13 4 9 9 13 2
18 9 10 2 13 9 13 9 9 13 2 9 9 10 9 12 13 4 2
23 3 2 9 2 9 9 7 9 9 15 9 13 2 10 9 0 13 4 9 12 13 4 2
19 10 2 11 12 13 4 3 11 2 12 9 13 2 7 9 12 13 4 2
17 11 2 9 2 9 7 9 2 13 4 11 7 11 13 13 4 2
8 2 9 9 13 11 9 2 2
13 0 13 2 7 9 13 9 3 13 13 9 13 2
14 3 2 7 2 9 13 0 11 7 14 13 0 9 2
10 11 9 0 0 13 4 11 9 9 2
14 9 9 13 10 2 9 9 13 0 13 9 14 13 2
8 2 13 9 13 9 13 2 2
11 15 9 13 9 12 9 10 3 13 4 2
22 12 9 13 13 4 9 7 9 12 9 9 2 12 9 11 8 11 9 13 13 4 2
16 9 3 13 2 3 0 2 0 2 14 3 0 7 9 0 2
4 10 13 4 2
6 2 13 4 11 2 2
8 9 12 9 11 13 9 0 2
6 9 10 3 13 4 2
25 9 7 9 9 13 9 2 9 0 2 13 13 4 2 7 9 7 9 9 3 13 4 13 4 2
14 11 11 13 12 9 9 0 2 7 3 13 4 9 2
11 13 3 9 2 10 3 9 0 13 7 2
17 0 9 13 9 13 13 4 11 9 9 2 7 10 9 9 13 2
12 11 11 0 7 11 11 0 13 4 12 9 2
6 2 13 4 11 2 2
4 9 0 13 2
5 9 13 13 4 2
13 9 13 2 11 13 4 0 9 7 11 9 13 2
11 9 13 3 2 3 13 4 9 13 4 2
7 0 13 4 9 13 9 2
10 11 9 11 12 9 13 4 3 9 2
4 9 13 13 2
11 9 0 13 9 9 13 9 0 13 4 2
12 2 9 10 3 13 4 2 9 10 13 3 2
7 10 10 14 4 9 13 2
9 3 2 9 13 3 9 0 9 2
6 9 0 10 0 13 2
7 0 9 9 13 8 4 2
13 9 13 7 10 11 9 11 0 11 9 13 4 2
6 2 13 3 13 13 2
5 9 12 13 4 2
15 3 9 13 9 0 2 7 9 0 13 4 12 13 13 2
9 3 13 9 11 11 9 0 13 2
9 11 13 9 0 11 13 9 13 2
4 2 9 13 2
5 3 0 13 4 2
12 11 3 13 4 11 2 7 10 9 13 4 2
7 3 2 12 9 13 4 2
6 2 0 13 9 2 2
4 9 0 13 2
12 3 9 2 3 2 12 12 9 13 4 9 2
14 11 11 9 11 9 13 9 13 4 3 2 11 2 2
10 3 2 9 13 4 9 9 0 13 2
27 9 13 9 12 2 13 7 13 13 7 2 9 7 9 9 13 9 2 9 12 13 7 3 13 14 4 2
17 13 9 2 13 4 9 7 9 9 9 12 9 13 4 9 9 2
19 11 0 13 4 9 2 7 9 11 13 3 11 0 13 4 9 13 9 2
14 11 9 9 2 9 13 7 9 13 2 13 4 0 2
10 11 11 11 0 13 4 3 9 0 2
13 12 9 13 7 13 4 3 2 7 12 9 13 2
18 2 15 9 2 11 2 3 13 4 7 2 0 2 13 9 13 2 2
12 9 10 10 7 10 9 0 13 11 9 9 2
14 9 10 2 9 2 9 0 12 13 4 7 9 13 2
10 9 10 13 13 4 9 12 13 9 2
13 10 9 3 13 13 4 7 10 9 10 13 4 2
4 13 13 4 2
16 12 9 9 2 11 9 9 12 13 4 7 12 13 4 9 2
11 10 2 11 9 9 13 4 3 9 0 2
15 11 2 0 13 2 13 15 9 2 13 9 2 13 9 2
12 7 3 11 11 9 9 13 13 13 4 15 2
7 7 9 13 7 13 4 2
3 13 9 2
13 13 4 9 3 13 4 13 2 7 9 13 4 2
7 12 9 13 13 4 0 2
14 11 9 2 9 2 9 13 4 9 0 13 13 2 2
14 3 2 9 0 9 9 0 9 13 0 13 4 11 2
10 11 2 14 13 0 2 11 10 13 2
4 3 9 13 2
18 2 13 4 9 11 2 11 2 13 4 2 7 9 13 9 13 2 2
19 2 15 13 4 7 15 9 9 13 13 2 9 13 12 13 9 13 3 2
13 10 9 12 9 13 4 2 7 14 13 10 3 2
9 11 9 11 13 9 7 9 11 2
16 2 9 9 9 12 10 9 13 4 9 7 0 9 13 4 2
12 9 9 13 4 9 10 2 9 2 13 4 2
9 11 13 4 9 11 2 12 2 2
7 2 0 9 13 13 4 2
7 2 2 13 4 9 2 2
10 15 9 13 4 2 7 9 9 13 2
9 9 9 9 7 9 13 9 0 2
13 7 14 13 9 0 13 2 0 13 7 0 13 2
8 11 9 3 9 10 13 4 2
17 11 9 2 7 2 11 14 4 9 13 13 4 7 14 13 9 2
4 2 13 13 2
9 13 4 2 7 3 13 13 4 2
24 3 13 2 9 13 9 2 7 13 9 13 2 15 9 13 9 2 9 13 4 9 9 10 2
10 2 9 12 9 9 7 9 9 13 2
15 11 2 11 9 3 13 4 11 2 11 9 2 12 2 2
11 7 2 13 4 11 13 9 11 13 4 2
10 9 13 7 15 9 9 9 13 4 2
6 3 9 0 13 4 2
9 9 9 13 9 3 0 13 4 2
5 2 7 13 13 2
13 9 10 9 9 0 13 4 9 9 13 9 13 2
9 9 0 9 7 9 13 13 4 2
8 14 4 15 15 9 13 13 2
11 9 9 9 9 9 7 0 13 9 13 2
11 2 11 11 13 4 10 9 0 13 7 2
35 9 2 11 13 4 2 7 10 7 3 13 4 9 13 2 3 14 13 9 2 7 9 2 9 7 9 9 7 13 4 9 9 13 4 2
22 9 13 9 12 9 13 2 7 2 9 0 3 13 4 2 13 9 9 0 13 4 2
16 3 9 10 9 7 9 13 4 7 13 4 13 4 9 12 2
18 9 9 2 9 7 9 13 4 3 9 9 12 13 4 7 13 9 2
10 11 9 12 9 13 4 3 11 9 2
12 9 9 13 3 2 9 13 7 13 13 4 2
7 7 13 4 13 4 9 2
12 3 2 9 9 13 4 9 10 7 9 13 2
11 9 13 7 9 13 7 14 4 3 13 2
10 3 13 4 9 13 12 9 13 4 2
9 11 9 9 0 3 13 4 9 2
12 11 11 9 0 13 4 9 13 4 9 13 2
22 9 13 2 3 9 2 3 13 4 2 2 7 9 9 2 3 2 13 4 13 4 2
8 12 9 13 4 9 9 9 2
16 9 13 7 9 2 9 12 13 3 2 13 9 0 13 4 2
14 11 11 9 4 9 0 2 11 11 9 13 13 4 2
6 11 9 9 13 11 2
10 9 9 0 9 10 13 9 13 4 2
13 9 13 4 9 7 3 9 9 13 4 15 9 2
19 15 13 4 3 13 4 7 2 7 11 9 13 4 3 9 3 13 9 2
14 9 0 14 13 9 7 11 11 0 13 4 12 9 2
5 9 13 4 10 2
27 11 2 9 0 2 13 9 13 7 2 10 2 9 9 13 2 13 9 13 13 4 3 11 11 11 9 2
6 0 9 9 13 13 2
8 2 9 12 13 4 9 2 2
15 12 9 13 13 4 2 11 2 12 2 2 12 9 13 2
20 9 9 13 4 3 13 11 9 0 9 7 10 13 9 9 13 4 13 9 2
23 7 2 10 9 0 12 13 4 9 10 9 13 4 9 0 2 7 10 9 7 13 4 2
23 11 0 9 13 2 13 9 13 13 9 13 13 2 2 11 13 4 7 9 13 4 2 2
19 9 13 4 7 9 0 10 2 11 2 11 2 2 15 0 9 13 4 2
8 11 0 9 13 4 3 11 2
15 11 9 13 4 11 9 12 13 4 2 9 2 9 0 2
10 9 9 13 2 7 9 10 13 4 2
7 2 15 14 13 9 2 2
13 11 9 9 10 2 9 7 9 9 13 10 9 2
8 2 3 11 9 13 13 13 2
11 11 7 11 9 10 12 9 13 4 3 2
19 12 10 2 9 0 13 4 11 2 11 7 11 7 3 4 2 12 9 2
22 9 9 13 4 9 2 9 7 9 13 4 2 7 9 2 7 9 9 7 9 7 2
7 9 9 10 9 13 4 2
10 10 9 0 13 2 7 11 9 13 2
8 14 2 3 3 0 13 4 2
15 11 13 4 10 9 9 0 13 12 2 3 13 4 9 2
16 9 13 10 9 11 8 11 13 4 7 0 9 9 13 4 2
8 9 0 13 13 4 2 7 2
12 3 2 3 13 4 11 9 9 13 4 9 2
21 9 13 13 9 2 9 10 7 9 10 13 2 13 7 13 3 2 9 13 4 2
21 10 13 9 13 4 3 2 3 2 3 13 4 3 2 10 9 9 13 4 3 2
12 9 12 9 13 9 13 0 13 9 13 0 2
9 7 0 9 9 7 13 13 4 2
12 3 12 9 13 4 7 10 12 12 9 13 2
10 11 12 9 13 2 7 12 9 9 2
11 10 9 2 10 9 0 13 9 9 13 2
13 12 12 9 3 13 4 9 9 13 13 9 10 2
6 10 13 9 13 10 2
8 9 9 10 3 13 4 9 2
11 11 9 13 4 9 9 0 13 2 8 2
4 11 9 13 2
18 10 9 3 13 7 0 13 7 2 14 13 11 13 9 10 9 10 2
11 11 11 13 7 9 0 2 3 0 13 2
17 11 11 9 0 13 4 9 2 7 11 11 9 3 13 9 13 2
14 12 13 13 9 2 11 7 11 13 4 12 12 9 2
21 11 2 7 2 11 11 13 13 9 13 9 10 2 7 3 9 13 9 13 4 2
6 11 12 13 4 9 2
7 11 7 11 9 13 4 2
5 3 13 4 10 2
6 9 10 9 9 13 2
13 11 9 7 0 3 13 4 9 0 9 9 13 2
16 11 2 11 7 11 3 0 13 4 3 9 7 9 9 9 2
5 11 13 4 12 2
5 11 13 10 13 2
5 14 13 10 9 2
15 9 2 7 2 9 9 9 13 2 9 9 13 13 4 2
14 11 13 4 9 0 9 9 10 9 9 13 13 4 2
6 3 13 4 9 10 2
6 3 9 10 13 4 2
11 3 3 9 0 13 2 7 7 11 13 2
15 9 0 13 4 9 2 7 3 9 14 4 0 13 10 2
9 2 9 7 0 9 3 0 13 2
15 11 7 11 3 2 12 9 12 13 4 9 3 13 13 2
12 9 7 3 14 13 9 7 9 2 9 7 2
9 11 7 11 13 4 11 12 9 2
26 9 13 9 13 4 2 7 10 13 2 7 11 13 9 13 4 12 9 0 2 11 12 9 13 3 2
9 9 0 13 9 0 9 0 10 2
9 12 9 7 9 12 13 4 9 2
21 9 13 4 2 7 2 9 12 12 9 9 13 7 9 10 13 13 4 9 9 2
7 3 14 4 9 0 13 2
11 9 9 13 4 7 12 9 13 9 10 2
19 11 9 9 14 4 13 2 7 9 14 13 3 13 4 13 13 13 4 2
5 7 9 10 13 2
21 9 9 9 13 4 11 9 10 2 7 13 13 4 11 9 3 13 4 0 9 2
8 10 13 7 11 9 13 4 2
25 7 2 12 9 13 4 9 9 2 13 11 13 2 9 9 7 9 9 2 13 9 9 13 4 2
7 9 13 13 9 13 3 2
6 10 0 13 9 13 2
8 15 14 4 9 13 9 13 2
8 9 10 11 9 13 4 13 2
6 2 13 9 7 13 2
22 9 9 9 13 11 14 4 13 2 9 7 9 0 9 9 2 2 11 9 9 13 2
13 9 11 9 0 13 11 9 13 9 12 13 4 2
30 11 10 3 13 4 2 11 2 9 9 9 0 7 9 2 13 4 2 7 11 9 2 9 13 9 2 7 13 4 2
15 3 2 12 9 9 13 3 2 9 9 9 13 4 9 2
9 11 11 13 4 3 2 9 9 2
7 3 13 4 3 13 4 2
8 11 11 11 14 4 9 13 2
7 2 12 13 4 10 9 2
12 9 9 14 13 13 4 3 13 4 9 13 2
5 3 13 4 3 2
9 12 9 13 4 2 12 9 0 2
8 9 9 13 4 9 9 0 2
9 0 9 13 13 2 7 3 13 2
11 11 9 2 9 12 9 2 13 13 4 2
7 12 9 13 4 11 0 2
18 12 13 4 3 9 9 7 9 0 0 13 11 11 0 2 12 9 2
8 9 0 13 0 9 13 9 2
7 0 13 9 0 13 4 2
14 11 11 11 9 11 11 11 9 13 13 4 9 9 2
13 3 9 7 9 9 10 13 4 7 13 9 13 2
15 12 9 0 13 4 9 7 9 10 3 13 9 0 13 2
10 3 13 4 9 2 7 9 13 4 2
12 9 9 9 13 4 9 13 4 9 9 13 2
44 12 9 13 4 2 12 2 11 2 11 2 11 2 11 7 11 13 4 2 12 2 11 2 11 2 11 2 11 11 7 11 2 12 2 11 2 11 2 11 2 11 7 11 2
10 11 9 9 10 9 9 13 4 9 2
17 3 11 9 13 4 12 9 10 13 4 9 0 2 7 9 13 2
3 9 13 2
14 15 9 13 11 9 2 7 9 9 13 13 9 13 2
11 7 2 3 3 13 4 9 12 13 4 2
6 10 11 13 4 3 2
13 9 9 10 10 9 9 9 7 13 4 9 9 2
13 2 10 7 9 13 2 7 9 0 13 4 12 2
17 9 13 4 2 7 11 9 9 12 7 11 11 9 12 13 4 2
10 11 2 11 2 2 0 3 13 4 2
8 2 9 13 2 9 9 13 2
8 3 11 12 9 13 13 4 2
20 11 9 13 4 12 9 9 13 10 2 7 13 9 10 9 10 13 9 13 2
10 3 9 13 2 8 9 13 13 2 2
17 2 3 11 11 13 4 10 9 12 2 9 10 13 4 10 15 2
9 9 13 4 3 11 9 2 9 2
11 9 13 2 11 7 11 0 13 9 0 2
15 11 9 0 13 2 7 3 13 4 11 9 13 9 9 2
12 11 9 13 9 13 3 9 0 9 13 9 2
6 3 13 4 3 11 2
24 11 9 9 13 9 2 11 13 4 9 0 9 0 9 12 13 4 9 10 13 4 9 13 2
7 11 9 13 4 12 9 2
12 9 13 4 2 11 9 9 13 11 7 9 2
19 11 9 9 9 2 9 10 9 13 9 12 13 4 2 9 9 9 13 2
10 9 12 13 4 2 11 11 9 9 2
7 11 9 13 9 13 4 2
14 9 10 2 11 10 9 13 4 9 12 13 11 13 2
12 9 0 13 4 2 12 9 9 9 13 12 2
7 9 13 9 7 13 14 2
15 9 12 9 13 4 9 7 9 10 13 4 9 12 9 2
8 12 9 7 9 9 13 9 2
6 9 14 4 13 9 2
20 11 2 7 2 11 13 2 9 9 13 4 7 10 11 13 2 0 2 13 2
20 11 13 7 3 13 13 4 2 9 0 9 2 13 2 13 7 13 13 4 2
9 13 9 9 9 13 4 13 4 2
17 2 11 7 11 9 0 13 13 7 11 13 9 13 13 4 2 2
12 11 14 4 13 10 9 13 4 11 11 13 2
14 11 11 11 13 11 11 9 9 9 2 11 11 13 2
21 11 12 9 13 13 4 7 3 13 2 9 13 4 2 3 14 4 13 7 13 2
8 9 9 9 0 13 4 11 2
26 10 9 13 4 2 13 13 9 13 9 7 9 14 13 2 7 9 11 9 13 4 13 9 13 4 2
16 3 9 13 2 11 9 0 13 4 7 9 13 7 13 4 2
17 10 2 3 13 2 9 0 9 0 13 2 13 4 11 9 9 2
9 2 3 3 13 12 9 13 4 2
5 2 14 4 13 2
15 2 15 9 0 9 9 13 13 2 15 9 13 4 2 2
5 9 0 13 4 2
25 10 9 2 12 9 13 4 9 10 2 0 13 13 4 2 9 3 9 13 7 9 14 13 2 2
9 9 12 13 4 9 7 10 9 2
13 11 9 2 9 0 2 2 12 2 13 13 4 2
16 12 9 12 12 9 13 4 9 2 7 14 4 10 9 13 2
10 11 11 9 0 9 13 4 9 0 2
12 9 9 9 13 4 2 9 12 9 13 4 2
11 11 9 9 0 13 7 3 13 4 9 2
5 0 13 0 10 2
6 10 13 3 9 9 2
16 7 2 12 9 11 9 13 4 11 12 9 3 13 4 3 2
13 9 10 13 4 9 2 7 9 7 9 10 13 2
21 9 9 2 7 2 9 0 12 13 4 2 7 9 0 0 10 13 9 13 4 2
13 7 9 13 9 13 4 13 4 12 9 10 13 2
11 15 9 12 9 13 13 4 2 3 9 2
13 9 9 9 11 11 9 7 9 9 13 4 9 2
15 9 2 9 9 12 13 3 2 14 13 2 14 4 13 2
14 0 12 9 13 3 2 7 11 13 9 13 9 13 2
21 11 9 13 0 13 7 13 4 12 9 9 13 4 9 2 9 0 0 9 2 2
6 2 9 13 4 2 2
7 9 2 11 9 9 13 2
15 3 11 11 9 13 4 9 2 7 10 13 4 9 9 2
4 11 13 13 2
16 11 2 11 2 11 7 11 9 0 13 4 11 11 9 9 2
11 9 13 12 9 0 11 7 9 9 13 2
8 13 4 3 11 13 13 4 2
8 9 13 9 3 13 4 9 2
11 10 13 4 2 7 11 9 10 9 13 2
9 11 9 9 13 4 2 12 2 2
13 3 9 13 7 10 3 13 13 2 3 7 3 2
11 9 10 9 7 13 2 0 9 13 4 2
4 13 4 3 2
12 9 9 14 4 15 13 9 2 7 9 0 2
13 9 12 9 7 9 13 7 9 9 12 13 4 2
11 12 10 2 7 2 9 7 0 13 4 2
18 9 9 2 12 9 9 13 2 3 7 3 11 9 13 9 13 4 2
9 2 9 7 0 9 0 13 3 2
5 11 13 4 3 2
20 11 2 7 2 9 13 4 11 13 4 13 4 7 14 4 9 13 9 13 2
7 10 0 13 9 13 10 2
19 9 10 9 9 13 9 9 13 4 9 2 9 9 13 9 13 4 3 2
5 9 14 4 13 2
14 3 2 13 9 9 12 9 13 4 7 12 9 9 2
26 9 0 12 9 13 2 9 0 12 9 2 14 12 2 2 7 9 9 9 13 4 2 9 9 0 2
15 7 13 7 13 4 11 9 9 3 0 13 4 9 10 2
10 0 13 4 9 7 0 13 4 9 2
7 2 9 13 4 11 2 2
12 9 0 13 13 4 11 13 13 4 9 13 2
10 13 9 12 9 2 13 4 9 9 2
16 9 0 9 9 10 13 4 2 7 9 9 13 4 9 13 2
5 9 14 4 13 2
8 9 13 4 9 0 13 4 2
4 3 13 4 2
14 11 7 2 9 10 13 9 9 2 9 0 13 4 2
13 9 2 11 2 11 2 13 4 9 9 13 4 2
16 2 9 15 13 9 13 4 2 9 0 10 0 13 4 2 2
7 11 13 3 9 13 4 2
6 11 7 0 13 4 2
6 3 2 13 9 13 2
15 9 0 7 13 4 9 9 13 4 9 13 4 13 13 2
9 9 2 7 2 9 9 9 13 2
4 13 4 7 2
10 11 9 2 11 2 9 10 9 13 2
10 2 11 15 9 13 4 13 9 13 2
13 11 11 9 0 0 9 13 4 3 2 11 9 2
4 9 13 4 2
9 10 7 0 13 2 3 13 4 2
10 9 13 4 11 11 9 13 12 9 2
11 11 10 13 4 9 2 11 9 3 13 2
5 7 3 0 13 2
13 11 9 11 9 13 12 9 13 4 13 4 9 2
5 0 13 2 9 2
7 9 9 3 13 13 9 2
11 15 9 13 2 7 15 7 13 13 4 2
11 15 13 4 12 12 9 0 9 10 13 2
12 11 7 2 12 9 9 9 13 13 4 9 2
5 0 15 13 13 2
11 9 10 9 9 7 9 0 9 13 4 2
7 2 10 9 13 4 9 2
17 9 9 13 14 7 2 9 0 13 9 13 9 13 4 11 9 2
6 7 2 9 13 4 2
6 0 13 2 7 3 2
16 9 9 9 9 13 13 7 10 9 13 9 14 4 13 11 2
14 11 9 11 13 9 13 4 2 13 13 9 13 7 2
20 12 12 9 10 7 10 9 11 9 9 13 4 3 2 9 9 0 13 9 2
6 11 9 9 9 13 2
12 12 11 13 4 7 12 9 12 9 13 4 2
6 14 13 10 13 4 2
10 10 9 9 13 4 11 11 13 4 2
15 15 9 13 13 9 2 11 2 11 11 7 11 9 2 2
13 9 0 9 10 12 9 9 7 9 10 13 4 2
17 11 2 11 11 2 11 11 2 11 7 10 11 13 13 4 3 2
17 9 9 12 13 2 7 2 3 2 11 9 13 4 2 9 13 2
13 3 3 11 13 4 9 12 13 2 9 2 11 2
14 9 3 13 4 9 9 9 13 2 3 9 13 4 2
13 9 12 9 13 4 12 12 9 2 15 13 4 2
13 9 11 13 11 9 9 13 2 7 9 13 4 2
8 11 11 7 11 11 13 4 2
6 9 13 3 13 4 2
18 9 9 9 13 4 2 7 10 9 9 13 7 15 9 9 13 4 2
13 7 2 9 7 9 0 13 0 9 10 12 9 2
7 12 13 4 9 3 12 2
23 9 10 10 12 9 0 13 4 11 9 2 7 3 2 0 9 2 13 4 11 9 10 2
11 11 7 11 11 14 4 13 13 4 11 2
9 9 13 7 13 10 13 4 11 2
8 9 0 12 9 13 4 9 2
14 2 9 10 13 4 9 0 7 9 9 13 13 4 2
9 2 9 7 0 9 0 13 3 2
4 10 13 10 2
7 11 9 13 4 9 9 2
5 9 3 13 13 2
7 9 3 9 0 13 4 2
8 15 2 7 2 14 4 13 2
9 9 10 9 2 9 2 13 4 2
11 2 9 13 4 9 13 9 14 13 2 2
6 0 0 9 13 4 2
9 9 9 2 7 2 9 13 4 2
11 2 11 9 0 13 7 9 0 9 13 2
12 11 13 9 2 9 2 13 4 9 13 4 2
8 9 13 4 9 13 7 13 2
10 7 2 11 9 0 13 4 11 9 2
5 13 10 13 2 2
13 9 0 13 9 13 2 9 13 13 4 13 11 2
22 11 13 9 10 13 4 9 10 2 11 2 7 2 13 4 12 9 0 12 9 13 2
7 9 9 0 10 9 13 2
7 15 9 12 9 0 13 2
10 9 13 7 2 9 0 13 9 13 2
8 12 13 4 9 7 12 13 2
6 2 3 13 3 13 2
11 2 9 4 7 2 14 4 3 13 2 2
8 2 13 3 13 4 2 9 2
3 9 13 2
13 11 7 11 9 13 2 12 9 11 15 13 4 2
16 12 13 4 9 2 7 3 13 4 11 9 2 11 11 9 2
16 11 9 10 9 9 13 13 4 2 12 9 14 4 9 13 2
12 11 9 0 13 2 7 3 9 9 13 4 2
18 3 13 4 15 7 11 9 13 13 2 11 9 13 2 15 13 4 2
9 14 4 9 13 9 2 14 9 2
5 11 3 13 4 2
6 3 13 4 9 0 2
5 9 9 13 4 2
30 14 9 9 2 14 11 0 13 4 9 9 12 9 13 9 0 12 3 3 13 2 7 10 9 2 9 9 0 13 2
31 3 2 3 2 9 13 9 7 9 9 13 4 9 12 13 2 7 9 15 13 14 4 3 13 4 2 14 9 14 9 2
10 9 9 2 3 2 14 4 9 13 2
7 3 2 14 13 9 0 2
14 2 9 0 13 3 2 9 7 9 2 7 2 14 2
19 3 13 4 11 2 11 12 2 11 12 2 11 12 2 11 12 7 11 2
25 12 9 10 2 9 9 13 9 13 4 2 9 9 0 12 9 7 9 9 0 9 13 13 4 2
5 10 13 4 9 2
9 2 0 13 13 7 13 4 2 2
15 0 13 2 3 12 9 12 9 13 9 0 11 9 13 2
17 9 0 13 11 9 13 4 2 10 9 13 7 9 9 12 13 2
5 9 3 13 4 2
11 11 9 9 2 9 3 2 3 13 4 2
13 9 7 9 9 12 0 13 2 9 0 3 13 2
14 9 10 9 10 9 13 4 2 9 9 0 13 4 2
4 3 13 9 2
8 9 7 13 4 9 0 10 2
6 15 9 13 4 3 2
16 9 9 10 13 7 9 12 9 13 4 2 10 12 9 13 2
16 9 12 9 9 13 4 12 9 2 11 9 12 9 0 13 2
17 9 13 9 9 13 9 0 9 9 13 7 10 11 7 13 4 2
7 9 13 9 10 13 9 2
6 13 2 13 2 9 2
23 9 2 7 2 14 4 13 9 13 2 7 9 9 9 10 9 13 7 3 3 13 4 2
10 9 10 13 3 13 4 9 13 4 2
8 2 9 9 0 13 4 2 2
18 7 9 0 12 3 13 9 13 9 2 7 12 9 9 12 13 13 2
10 9 10 13 13 2 3 13 4 9 2
10 2 9 10 9 10 13 13 4 2 2
10 3 2 12 9 0 9 7 13 4 2
6 3 9 0 13 4 2
19 13 9 13 7 9 9 13 2 9 0 13 9 13 13 4 11 9 0 2
5 12 9 13 4 2
5 9 13 0 10 2
8 11 13 9 13 4 9 0 2
7 11 9 0 13 13 4 2
12 11 9 7 10 9 9 14 4 3 3 13 2
6 11 7 11 13 4 2
5 2 9 13 4 2
21 11 7 11 14 4 3 10 9 9 13 2 7 12 7 12 3 13 4 10 11 2
6 7 10 7 13 4 2
7 9 0 13 4 3 9 2
5 9 13 13 13 2
12 9 7 9 9 0 10 9 7 9 13 4 2
15 9 0 9 13 2 7 9 10 2 9 2 0 13 2 2
7 2 9 3 13 4 9 2
7 2 9 13 13 4 2 2
11 7 13 4 9 9 13 14 4 15 13 2
9 2 9 13 4 9 13 4 0 2
12 2 9 13 10 10 9 9 13 14 4 2 2
7 11 7 11 0 13 4 2
24 7 2 11 9 2 9 0 14 2 4 13 13 4 2 2 9 9 3 13 2 4 13 3 2
3 9 13 2
7 11 11 13 9 13 4 2
13 7 9 0 9 14 13 9 13 2 14 4 13 2
8 14 4 3 13 2 13 13 2
17 13 9 12 11 13 11 9 0 9 3 13 4 3 2 11 9 2
15 11 12 13 9 11 0 3 13 4 9 2 9 3 13 2
4 9 9 13 2
27 9 9 0 14 13 7 2 9 9 9 0 13 7 9 3 13 4 13 4 2 9 13 9 0 13 7 2
13 7 9 13 9 13 2 7 9 3 13 4 11 2
13 12 9 11 13 9 2 13 2 13 13 4 11 2
13 9 9 13 7 9 13 4 2 10 13 7 13 2
8 9 9 13 4 11 9 9 2
11 2 9 3 13 13 2 9 0 12 13 2
8 2 11 13 13 9 10 13 2
21 9 7 9 13 9 13 4 9 2 7 9 9 13 13 4 9 9 2 12 9 2
10 2 13 9 9 10 9 0 13 2 2
29 9 13 4 9 11 11 9 11 12 12 13 2 7 12 9 13 9 2 11 9 2 11 11 11 9 13 9 13 2
8 3 13 4 9 13 12 9 2
15 11 7 11 9 12 13 4 9 2 7 14 4 10 13 2
11 9 9 13 4 3 2 7 12 13 4 2
16 9 9 0 13 2 9 0 13 7 9 0 13 9 3 13 2
10 9 2 9 13 2 9 9 13 4 2
6 9 9 12 13 4 2
6 3 13 4 0 9 2
23 3 7 3 13 13 4 9 2 10 7 13 13 4 7 2 10 13 3 2 3 13 4 2
4 9 12 13 2
8 9 2 7 2 9 13 4 2
11 9 12 13 4 9 11 9 2 0 2 2
17 10 9 4 3 13 2 7 7 2 9 0 10 7 13 9 13 2
11 3 2 11 13 13 4 11 11 9 13 2
14 12 9 2 11 13 4 2 3 9 0 13 4 9 2
15 9 9 13 13 9 9 13 7 9 9 0 13 9 13 2
6 2 0 13 7 13 2
6 13 15 2 14 13 2
14 9 9 12 11 9 9 13 4 7 9 12 13 3 2
16 9 7 9 12 13 4 12 9 13 4 9 2 12 9 2 2
11 9 11 9 13 4 12 2 11 12 13 2
12 9 12 13 4 2 7 12 9 13 4 3 2
12 11 7 2 9 9 13 4 2 3 13 4 2
8 11 9 10 14 13 10 9 2
3 10 13 2
5 9 13 11 11 2
5 3 13 4 10 2
21 9 9 9 13 4 7 11 7 11 9 13 4 2 3 7 14 4 9 13 11 2
7 9 9 9 13 4 11 2
6 14 13 0 0 13 2
20 7 9 10 9 10 7 13 4 2 12 9 13 9 9 13 9 13 4 9 2
7 12 9 3 13 4 0 2
18 9 7 9 3 13 2 7 9 10 13 9 2 13 13 4 15 9 2
5 10 13 4 10 2
16 14 4 10 9 3 13 7 2 9 3 9 13 14 4 9 2
9 13 4 2 3 13 13 10 9 2
19 11 9 13 4 2 11 9 13 3 9 9 13 7 14 4 3 13 9 2
7 3 13 4 9 9 9 2
14 11 9 9 3 13 3 2 11 9 13 4 2 7 2
20 9 9 13 9 9 10 3 13 2 11 10 13 4 3 2 10 9 3 13 2
19 11 9 13 10 9 2 7 3 13 9 13 4 2 2 13 4 3 11 2
12 2 13 15 9 9 0 13 4 15 9 13 2
8 14 13 3 13 9 0 12 2
20 11 2 3 11 9 2 12 9 13 4 2 12 13 4 11 2 7 12 11 2
6 9 0 12 9 13 2
12 10 9 0 13 2 9 0 7 13 9 10 2
13 3 2 9 13 13 4 2 7 12 9 13 4 2
10 14 13 11 12 9 3 3 13 4 2
19 11 0 13 11 0 9 0 2 9 7 9 9 7 9 13 11 13 4 2
22 10 3 2 7 2 9 9 13 4 2 13 12 3 2 7 9 7 9 13 10 3 2
21 3 2 9 0 2 13 4 10 13 7 13 4 9 11 2 3 9 7 9 13 2
18 9 9 2 10 9 3 13 9 13 4 9 13 4 13 4 3 2 2
17 3 2 9 7 9 9 9 13 7 9 0 13 4 13 4 0 2
4 11 13 4 2
24 10 2 9 0 11 7 9 0 9 13 13 4 11 2 7 11 9 7 13 9 13 13 4 2
12 7 2 12 9 2 10 12 9 13 4 0 2
16 3 13 4 10 13 4 2 7 15 14 13 9 9 9 0 2
9 3 11 7 11 9 10 13 13 2
5 9 0 10 13 2
7 9 0 9 13 4 9 2
6 13 9 0 9 12 2
19 9 13 2 9 9 9 13 4 2 12 2 12 2 12 7 12 9 9 2
5 10 9 13 4 2
8 3 13 14 4 9 13 4 2
5 9 13 4 13 2
10 7 9 0 9 9 9 0 13 4 2
16 0 13 2 15 3 13 13 4 2 7 3 9 3 13 4 2
8 2 9 9 9 13 13 3 2
7 7 13 4 13 4 3 2
12 11 3 13 4 9 11 9 9 7 9 13 2
11 9 9 9 9 13 7 9 9 13 4 2
12 11 13 4 2 10 13 4 9 2 0 4 2
11 9 13 4 7 3 13 4 9 9 13 2
7 3 2 3 13 4 13 2
14 9 0 13 4 2 7 9 9 13 9 10 13 4 2
15 7 11 11 8 9 0 13 3 7 12 9 13 4 9 2
11 9 0 13 9 13 4 9 0 13 3 2
14 9 2 9 2 2 9 13 4 7 3 13 9 13 2
10 9 13 13 4 9 14 13 3 0 2
14 11 9 2 7 2 9 12 8 15 10 7 13 4 2
7 15 9 13 4 3 9 2
12 9 10 13 9 13 4 11 2 9 9 9 2
4 11 9 13 2
19 12 2 13 4 0 10 12 9 12 13 4 10 3 13 4 9 14 13 2
6 0 9 9 13 2 2
11 9 12 2 3 13 4 3 13 13 9 2
18 11 11 9 0 9 13 9 13 4 11 9 9 9 9 12 13 9 2
28 2 15 9 0 13 4 2 9 0 13 4 9 0 2 9 9 13 4 7 0 9 9 13 9 13 4 2 2
10 11 9 12 9 3 13 4 9 10 2
6 14 13 3 2 7 2
13 9 14 13 2 10 13 4 9 2 7 9 9 2
14 9 0 14 13 7 2 11 13 9 3 13 4 9 2
29 14 4 13 11 9 11 11 2 11 2 11 8 11 2 7 11 11 0 2 11 2 2 3 13 7 9 13 13 2
30 9 9 13 9 13 7 2 2 3 13 2 13 9 2 7 9 10 13 4 9 13 4 3 13 7 9 9 9 13 2
16 10 7 11 13 4 2 11 13 2 7 9 9 0 13 4 2
9 9 12 11 9 13 13 4 9 2
14 9 10 2 11 13 4 2 3 9 0 2 13 9 2
11 9 0 13 9 0 13 11 9 9 0 2
18 9 0 9 9 9 9 13 4 3 9 11 11 13 9 9 12 9 2
11 11 9 13 9 11 11 13 9 13 13 2
18 9 9 9 7 9 13 2 9 10 13 4 2 7 9 0 13 2 2
16 3 9 9 13 2 11 9 3 9 0 13 4 13 9 13 2
7 12 9 9 13 4 9 2
5 3 11 13 0 2
17 11 11 2 12 9 0 9 13 9 4 2 7 3 9 0 13 2
12 9 0 13 3 9 13 7 9 13 13 4 2
7 14 2 3 0 13 10 2
10 2 11 13 2 0 2 13 9 0 2
20 7 2 9 13 0 13 2 12 9 12 9 7 12 9 13 14 13 9 0 2
6 9 13 7 12 13 2
15 12 9 2 9 2 9 7 9 2 13 9 9 13 4 2
9 9 10 9 9 9 9 13 4 2
6 3 13 4 9 9 2
10 9 0 13 4 2 7 10 3 13 2
6 2 15 9 13 4 2
8 9 13 9 13 2 14 9 2
11 9 12 13 7 3 12 13 4 9 10 2
15 11 9 0 10 13 4 12 9 2 7 14 4 15 13 2
16 3 2 11 9 9 13 7 9 12 9 13 9 13 4 9 2
19 9 9 13 11 9 0 7 11 13 9 11 13 13 12 9 11 9 9 2
19 11 9 13 4 9 2 7 12 9 13 13 4 9 2 9 0 13 4 2
6 12 9 0 13 4 2
9 9 10 9 13 4 3 11 9 2
7 3 9 0 13 13 9 2
6 12 9 13 11 13 2
5 11 13 13 4 2
12 6 2 15 11 13 7 15 9 9 13 4 2
3 9 13 2
10 9 13 9 2 14 13 2 14 13 2
12 3 9 9 0 13 9 2 7 9 13 4 2
5 10 13 4 15 2
30 11 13 4 0 9 0 12 13 4 9 13 4 12 9 2 7 13 4 2 7 2 12 9 13 4 11 13 9 12 2
17 10 9 0 13 11 7 9 13 9 13 10 13 9 13 9 13 2
10 11 9 9 13 13 4 11 7 11 2
16 11 11 11 11 11 9 11 13 4 3 2 11 9 9 13 2
9 15 9 2 9 13 4 13 4 2
10 9 9 10 13 2 15 9 9 13 2
9 2 9 3 13 4 15 9 2 2
15 11 9 9 10 13 9 13 4 11 9 9 11 13 9 2
17 7 2 10 13 9 9 13 2 9 9 13 9 0 0 12 13 2
12 9 0 2 0 2 3 0 7 9 0 13 2
18 9 0 9 2 9 2 9 2 12 7 12 2 2 9 7 9 13 2
10 9 0 13 13 4 7 14 4 13 2
11 12 9 7 2 12 9 13 10 9 0 2
11 9 0 2 7 2 10 9 13 13 4 2
6 3 0 13 9 9 2
8 7 9 3 14 13 13 4 2
14 9 9 9 13 4 13 3 2 9 9 13 13 4 2
7 13 3 2 9 13 4 2
5 3 10 13 4 2
32 9 9 2 3 2 10 9 9 7 9 3 13 4 2 9 0 9 0 12 13 9 13 4 2 3 2 3 9 9 13 4 2
24 7 2 9 13 4 9 9 12 13 3 11 9 14 13 2 7 10 13 4 10 13 9 9 2
12 9 12 9 13 4 2 7 10 3 13 3 2
26 9 9 9 2 12 10 12 13 4 9 0 13 4 9 7 9 9 13 7 12 9 7 9 9 13 2
4 9 13 4 2
5 13 0 4 7 2
11 3 12 13 2 7 12 13 7 13 4 2
8 7 2 11 3 13 9 10 2
7 2 14 2 3 13 4 2
16 7 2 12 12 9 14 4 9 13 7 10 13 9 7 13 2
12 11 11 7 11 11 9 9 13 4 11 9 2
12 11 9 9 13 2 7 9 13 9 13 4 2
9 13 4 9 13 4 12 9 0 2
6 2 9 9 9 13 2
3 9 13 2
10 11 7 11 2 7 2 9 0 13 2
5 9 9 14 13 2
9 9 0 13 4 2 13 4 9 2
11 9 13 4 9 0 3 13 4 13 4 2
8 9 0 12 9 7 14 13 2
14 3 2 9 0 9 13 4 2 7 12 9 13 4 2
18 11 2 7 2 12 9 12 9 9 13 13 4 2 9 10 13 4 2
10 0 13 2 12 9 13 4 10 9 2
18 9 9 7 3 9 10 13 2 11 9 0 13 9 13 9 13 4 2
4 9 0 13 2
3 13 4 2
11 7 2 0 9 13 9 9 9 9 10 2
6 9 9 13 9 12 2
10 11 11 13 4 2 11 12 9 0 2
8 2 14 13 2 11 14 13 2
11 2 9 9 10 13 4 9 14 13 2 2
17 7 2 14 4 13 2 14 4 11 13 7 11 9 13 13 4 2
9 3 9 0 13 9 9 13 4 2
8 9 11 9 13 4 2 12 2
22 10 9 10 11 11 11 2 11 11 11 2 11 11 2 11 11 7 9 11 13 13 2
13 11 9 9 13 7 2 9 13 9 2 13 4 2
10 9 13 4 9 12 9 9 13 4 2
8 12 9 0 9 0 13 4 2
7 11 9 9 13 9 13 2
12 0 9 13 13 9 9 13 4 9 13 9 2
12 9 10 0 12 9 10 13 4 11 0 12 2
11 9 9 2 11 7 11 9 15 13 4 2
13 9 10 9 0 12 7 13 4 2 10 13 3 2
7 15 9 7 9 0 13 2
14 11 13 4 9 9 11 7 13 13 4 11 9 0 2
10 9 9 13 4 9 13 4 9 10 2
15 9 9 13 13 4 3 9 2 7 9 13 9 13 4 2
9 9 9 13 2 9 12 13 11 2
10 2 0 2 13 7 9 0 13 4 2
9 9 10 3 13 4 9 9 9 2
16 9 13 14 7 2 9 0 13 2 7 9 9 0 13 13 2
9 9 13 13 9 2 2 13 0 2
13 15 9 10 13 9 0 7 3 9 9 13 4 2
6 9 9 9 13 4 2
18 12 9 9 13 4 11 9 12 9 9 13 2 7 0 13 9 13 2
11 9 7 9 9 7 13 4 3 0 13 2
6 2 13 10 13 4 2
9 14 3 15 13 2 3 2 3 2
16 9 13 4 9 9 12 13 4 9 13 2 9 10 9 13 2
14 9 13 9 9 10 13 4 2 9 9 12 13 4 2
14 9 13 2 9 0 13 2 7 0 7 13 9 0 2
30 11 2 11 2 11 7 11 13 4 12 9 2 11 2 11 2 11 7 11 9 7 11 2 11 2 11 7 11 9 2
7 11 9 12 13 13 4 2
10 13 4 9 2 12 9 13 4 9 2
10 9 10 9 13 9 0 10 15 13 2
19 9 9 13 9 13 9 9 13 9 13 4 2 7 10 9 13 4 3 2
29 2 11 9 13 13 4 7 2 7 2 10 14 4 0 9 13 2 11 0 9 13 11 2 2 13 4 11 9 2
22 11 11 11 7 11 11 9 13 4 11 14 13 2 9 0 2 9 13 7 9 13 2
15 2 9 9 13 4 2 9 0 13 7 12 9 9 13 2
7 9 9 3 13 0 13 2
11 0 9 2 11 0 9 12 9 13 9 2
13 14 13 0 2 9 7 9 13 2 3 10 13 2
10 11 13 4 2 7 2 12 13 4 2
9 2 2 9 13 11 12 9 13 2
7 9 13 9 13 4 10 2
7 2 10 15 9 13 2 2
7 10 13 9 12 13 4 2
8 9 0 13 9 9 13 4 2
11 2 3 2 11 9 15 9 13 13 4 2
4 9 0 13 2
9 11 2 9 0 2 13 4 9 2
12 2 9 10 9 13 3 9 0 13 4 11 2
21 11 11 12 9 9 0 13 4 2 7 11 9 9 13 9 13 4 9 9 10 2
16 11 7 11 13 13 2 7 12 9 10 9 13 4 9 0 2
24 2 11 9 13 7 12 9 9 13 4 2 9 9 13 13 4 2 9 9 12 9 13 4 2
6 3 13 10 13 9 2
19 9 10 12 9 13 11 7 11 11 9 9 13 9 9 12 9 13 4 2
16 3 14 4 9 2 9 7 9 0 0 13 13 9 9 13 2
15 3 7 9 0 9 13 4 9 14 4 9 0 9 13 2
15 9 9 13 2 7 14 13 0 2 9 14 4 13 2 2
9 3 14 4 10 9 13 9 10 2
18 7 2 9 9 14 4 0 9 13 13 13 2 3 9 9 13 4 2
12 9 10 9 11 13 2 13 4 7 13 4 2
28 11 12 9 9 9 9 0 13 7 2 14 4 9 13 9 0 2 7 13 13 13 9 10 13 11 9 9 2
4 9 13 4 2
12 9 2 9 2 13 9 13 13 4 11 9 2
5 9 9 0 13 2
20 2 3 12 9 13 4 9 13 4 2 7 9 10 9 13 9 13 9 13 2
13 11 9 12 9 11 11 0 13 4 2 11 9 2
5 10 13 9 10 2
4 3 13 4 2
18 2 0 13 4 2 7 14 4 13 9 13 4 2 2 13 4 11 2
5 11 13 4 11 2
13 11 9 11 7 11 11 7 11 9 13 4 3 2
6 3 13 4 15 9 2
22 11 9 3 9 13 4 2 12 2 2 7 11 0 0 13 7 2 3 13 13 4 2
5 9 9 13 4 2
5 7 14 4 13 2
16 10 4 7 2 11 13 9 9 10 2 13 2 13 13 4 2
6 9 14 13 3 11 2
7 9 12 13 4 2 3 2
3 13 3 2
8 9 12 9 12 13 4 3 2
8 11 9 12 9 13 3 13 2
9 11 12 13 4 12 9 7 9 2
6 9 3 3 13 4 2
8 11 9 0 9 13 4 3 2
8 2 9 9 13 13 9 13 2
14 11 9 11 0 9 13 4 11 9 13 9 0 13 2
12 2 9 9 7 13 2 13 13 4 10 9 2
9 3 13 9 9 12 13 4 9 2
7 9 13 13 13 9 13 2
10 10 9 13 3 2 11 9 13 4 2
11 7 2 3 2 9 0 12 13 4 3 2
9 14 14 4 0 9 13 9 0 2
6 9 9 0 13 4 2
19 0 13 9 0 7 0 13 4 9 13 4 2 7 11 9 13 13 4 2
11 10 2 9 9 13 4 9 10 13 4 2
21 11 11 2 11 11 7 11 11 9 9 9 12 13 4 2 7 9 9 12 13 2
12 9 13 9 2 9 0 10 0 7 13 7 2
17 9 0 9 2 9 2 9 2 9 2 2 13 9 10 9 13 2
7 9 9 2 10 0 13 2
6 9 14 13 13 13 2
10 9 10 8 0 13 2 14 2 11 2
7 3 2 11 9 13 4 2
11 2 9 0 2 13 4 9 4 9 9 2
7 9 0 9 13 2 9 2
10 11 7 11 9 0 13 4 9 9 2
30 2 9 0 2 9 13 13 11 2 7 3 13 4 14 11 2 14 9 9 14 13 11 0 2 2 9 0 7 2 2
8 9 14 4 13 13 9 0 2
9 13 13 13 4 2 11 9 13 2
9 9 10 14 4 3 3 13 9 2
20 9 0 10 13 4 11 12 9 7 9 9 7 10 9 13 4 9 10 13 2
8 7 15 9 13 3 0 13 2
13 3 14 13 11 13 0 2 7 9 12 13 4 2
15 9 9 9 13 7 2 9 0 9 3 0 13 13 4 2
9 2 10 9 13 2 10 13 4 2
11 9 13 8 4 9 10 9 9 13 4 2
7 0 9 2 11 13 4 2
14 9 13 10 7 9 13 13 11 3 9 0 9 13 2
16 9 0 0 10 13 4 9 2 13 4 15 2 14 9 9 2
10 9 12 9 13 4 9 13 9 13 2
14 2 12 9 12 9 13 4 2 7 9 13 4 13 2
5 15 9 0 13 2
8 11 9 9 13 13 4 9 2
11 13 9 13 4 3 11 11 9 13 9 2
15 9 14 4 13 11 3 0 13 2 7 14 4 15 13 2
20 2 9 13 14 4 2 7 9 9 13 2 9 9 12 13 4 13 9 2 2
12 3 0 13 0 9 13 9 12 9 12 13 2
4 13 4 11 2
11 9 9 12 13 4 0 2 12 9 13 2
15 11 11 9 12 13 4 7 2 3 2 11 11 10 12 2
26 9 9 9 12 13 4 7 2 9 14 4 9 13 13 4 3 2 7 11 13 4 2 11 12 9 2
10 11 11 9 0 9 13 13 4 3 2
18 9 10 3 3 13 4 13 4 9 9 9 0 2 13 12 9 2 2
13 11 9 8 0 13 4 2 7 2 11 11 9 2
19 11 13 4 9 10 13 4 2 7 14 4 9 13 2 3 14 13 3 2
6 14 4 3 0 13 2
5 9 3 13 4 2
18 11 9 13 4 2 11 7 11 9 2 11 9 9 13 13 4 2 2
6 2 3 13 13 4 2
10 12 9 11 9 11 11 11 13 4 2
12 9 0 2 7 2 12 9 13 4 13 4 2
11 9 2 11 7 11 7 3 13 4 9 2
14 11 13 10 2 7 9 0 13 10 7 9 13 4 2
15 11 9 13 13 4 2 7 12 9 7 0 13 9 4 2
11 9 3 13 2 7 10 10 9 3 13 2
12 9 13 4 10 15 9 7 13 13 9 13 2
7 2 3 7 13 4 3 2
30 9 14 4 0 13 2 7 11 13 0 9 9 13 2 9 13 2 10 13 7 11 13 4 9 2 0 11 13 4 2
13 2 7 9 9 13 13 4 9 13 13 9 2 2
11 0 9 0 13 4 3 11 2 7 13 2
12 9 13 9 13 4 2 9 7 9 0 2 2
7 3 0 12 9 13 4 2
13 9 9 7 9 12 0 13 9 9 13 0 13 2
20 9 10 9 12 13 4 2 9 13 9 13 2 9 9 13 4 9 10 2 2
8 2 11 9 0 13 4 2 2
8 2 3 11 14 13 9 0 2
8 3 12 9 9 9 13 4 2
24 12 9 7 9 12 3 13 15 13 2 14 4 9 0 12 13 7 9 0 3 0 14 13 2
6 13 9 7 13 4 2
19 11 11 7 11 9 13 13 9 13 4 2 7 9 0 13 4 9 9 2
13 9 9 13 2 9 9 2 0 2 9 13 13 2
7 9 13 9 13 9 9 2
17 9 9 13 9 13 4 11 2 2 3 13 9 3 0 13 2 2
8 13 9 10 15 9 13 4 2
15 3 13 4 11 0 12 2 7 10 10 13 9 13 4 2
8 11 3 13 4 11 9 9 2
9 11 9 9 10 7 0 13 4 2
7 12 9 9 13 4 9 2
9 9 12 12 9 9 0 13 4 2
8 7 2 9 9 13 9 13 2
4 9 3 13 2
7 7 9 10 9 13 4 2
9 9 0 13 4 9 9 9 9 2
17 2 12 0 9 10 13 4 7 2 10 9 13 9 10 13 2 2
7 12 9 9 9 13 9 2
12 13 2 14 4 13 3 9 7 10 0 13 2
11 15 9 11 14 4 9 13 9 13 2 2
10 10 9 11 9 9 9 9 13 4 2
8 3 9 3 13 13 4 9 2
8 9 13 9 9 0 13 4 2
5 9 13 4 9 2
22 9 0 13 4 0 9 0 9 13 4 9 9 2 7 3 13 4 9 13 9 10 2
8 2 9 14 4 11 9 13 2
10 11 11 9 9 9 9 13 4 0 2
5 2 9 12 13 2
21 9 9 0 13 13 13 9 13 3 2 7 10 7 13 4 0 13 11 9 9 2
20 3 2 9 0 13 4 2 0 11 13 12 9 0 9 13 9 13 13 4 2
11 0 13 14 4 2 11 13 4 9 0 2
14 9 10 0 9 9 13 2 9 13 4 13 9 2 2
24 12 2 9 0 2 9 13 4 9 9 12 2 13 2 7 10 9 0 13 4 9 9 13 2
9 7 15 10 10 13 13 9 13 2
4 14 13 9 2
4 13 4 3 2
13 11 2 9 2 13 11 4 9 0 13 12 9 2
10 11 11 9 9 13 7 9 13 4 2
5 12 9 13 4 2
10 9 10 14 13 7 3 3 13 9 2
15 3 9 0 9 3 13 4 7 13 7 9 14 4 13 2
10 9 13 9 13 2 7 13 13 4 2
7 9 9 13 13 13 4 2
21 10 12 9 13 9 0 9 3 13 9 12 2 12 9 9 12 13 4 10 9 2
5 9 13 4 9 2
10 9 0 12 9 13 4 9 13 9 2
17 12 2 10 13 2 10 10 13 13 2 3 13 4 11 9 9 2
11 2 13 9 2 6 10 13 4 12 9 2
11 11 12 9 13 4 9 9 10 0 13 2
11 11 11 3 11 13 9 9 13 4 9 2
10 11 8 11 13 9 7 13 4 9 2
9 2 10 13 9 7 15 13 9 2
18 9 9 11 9 0 9 2 2 9 9 2 7 10 9 13 13 4 2
12 0 7 0 13 2 7 9 3 0 13 4 2
5 0 9 0 13 2
10 3 12 9 13 4 9 12 9 10 2
16 9 10 9 13 9 9 13 4 2 7 10 13 4 11 9 2
17 2 15 9 9 9 0 13 11 2 7 3 3 13 10 9 2 2
13 9 7 13 13 2 15 9 13 4 9 13 4 2
9 9 9 11 9 13 4 2 9 2
18 0 9 11 9 9 13 4 2 7 10 13 7 12 9 9 13 4 2
6 3 9 0 13 4 2
21 3 13 4 11 11 11 0 11 12 9 9 13 2 12 9 0 9 13 13 4 2
10 11 2 7 2 3 3 13 4 9 2
11 11 11 11 9 9 13 4 11 9 9 2
8 7 2 9 9 13 13 4 2
12 11 11 13 4 7 13 13 10 13 4 11 2
5 2 9 9 13 2
7 7 10 9 13 2 3 2
9 15 9 13 9 0 15 15 13 2
18 11 9 0 12 13 4 3 9 3 7 2 10 2 14 13 9 0 2
22 11 13 9 12 2 12 13 12 13 11 13 9 13 7 3 13 2 9 9 13 4 2
9 9 0 10 13 13 4 9 13 2
29 11 9 12 9 0 2 0 2 0 7 0 13 4 9 2 7 9 0 0 13 4 3 2 14 4 9 0 13 2
8 12 9 9 9 10 13 4 2
15 15 9 9 12 13 4 7 9 10 9 9 2 13 4 2
13 7 2 3 13 4 9 13 9 0 7 13 4 2
23 11 9 14 4 3 13 9 0 2 3 11 9 13 3 9 0 11 13 9 0 14 4 2
12 9 13 9 9 0 13 4 2 9 9 0 2
4 15 13 3 2
5 2 3 0 13 2
19 12 9 0 10 12 9 13 9 11 2 7 2 9 13 4 2 9 13 2
9 9 10 2 11 3 13 11 9 2
12 9 0 10 9 13 12 9 13 4 11 9 2
4 2 11 13 2
12 11 0 2 2 14 4 3 10 9 9 13 2
7 11 10 9 13 13 4 2
5 11 13 0 9 2
25 11 9 0 13 3 13 2 7 14 13 0 2 9 12 10 13 4 2 7 10 13 9 13 11 2
13 7 10 13 4 9 11 7 11 14 4 9 13 2
11 9 13 9 13 4 11 11 11 7 11 2
8 13 4 11 7 9 12 3 2
8 9 13 7 9 13 4 11 2
9 3 2 11 9 0 13 4 11 2
6 9 0 13 4 9 2
21 12 9 4 2 12 9 13 2 9 10 13 4 13 2 7 9 12 13 9 13 2
10 7 2 0 9 7 9 13 9 9 2
8 9 9 13 3 3 13 4 2
20 3 2 13 13 4 9 0 7 14 4 0 13 2 14 4 13 9 10 9 2
7 9 0 9 13 9 13 2
4 10 13 4 2
9 10 13 7 13 4 9 9 13 2
5 9 13 4 9 2
9 9 9 11 9 13 7 11 9 2
12 9 10 9 9 13 2 7 9 13 13 13 2
11 2 3 12 9 13 4 11 9 13 2 2
6 9 0 13 4 9 2
4 7 3 13 2
9 7 13 13 9 0 11 13 9 2
15 9 13 3 12 9 13 13 4 3 2 7 9 13 4 2
14 9 0 9 13 2 12 9 2 9 13 9 0 13 2
8 15 9 0 12 9 13 13 2
10 11 9 10 12 9 13 4 3 11 2
16 11 13 4 2 13 2 11 9 0 0 2 10 15 8 3 2
8 9 13 10 9 13 4 9 2
18 11 13 3 9 13 7 9 13 7 11 9 9 9 3 0 13 4 2
13 13 4 2 7 2 9 13 9 13 7 9 13 2
16 9 13 9 13 4 9 7 2 0 2 13 13 4 12 9 2
19 9 9 9 9 13 4 9 2 7 15 9 3 13 9 13 2 11 3 2
11 11 8 11 3 13 2 9 9 13 4 2
6 9 0 13 4 9 2
12 2 11 2 3 9 13 4 3 13 4 9 2
6 2 9 9 13 2 2
5 9 13 4 9 2
14 11 9 2 11 9 0 13 4 2 7 9 11 9 2
12 11 9 11 9 12 13 2 3 9 13 4 2
14 11 9 13 9 13 2 13 13 4 11 7 11 9 2
4 9 0 13 2
8 9 13 4 2 9 7 9 2
11 9 0 9 3 13 2 13 2 13 4 2
9 3 14 13 3 13 4 9 13 2
15 9 13 14 13 0 13 2 7 11 9 9 0 13 4 2
15 9 0 12 13 4 9 9 2 7 10 9 9 13 4 2
17 7 2 3 2 9 9 0 13 4 9 2 7 12 13 13 4 2
16 11 11 0 7 11 11 0 11 11 11 9 13 4 0 9 2
10 9 10 2 0 9 10 13 4 9 2
12 3 11 13 4 11 9 10 9 12 13 4 2
6 9 14 4 13 3 2
8 14 13 2 15 9 4 13 2
9 3 13 4 11 11 11 9 7 2
8 7 2 9 13 11 9 13 2
6 11 14 4 9 13 2
8 11 13 14 4 13 9 10 2
11 9 2 12 9 13 9 13 4 2 11 2
16 9 9 9 9 11 9 13 4 2 7 10 0 13 4 11 2
16 9 9 0 13 4 12 9 2 7 10 11 9 13 13 4 2
12 9 9 0 2 12 9 12 11 9 13 4 2
12 3 13 4 10 9 2 10 9 2 10 9 2
6 2 0 9 13 15 2
15 10 13 4 11 9 9 2 3 11 9 9 9 13 4 2
10 9 10 13 4 2 3 2 9 9 2
12 9 13 2 0 9 0 12 9 13 4 11 2
17 15 13 4 2 7 2 9 9 0 13 2 9 9 0 9 13 2
6 12 9 13 4 9 2
11 9 10 9 13 9 13 9 14 4 13 2
7 11 9 13 9 13 4 2
5 14 4 13 13 2
14 14 4 9 13 9 12 12 9 7 9 0 13 4 2
18 9 3 0 13 2 9 7 9 13 2 7 10 14 4 9 13 11 2
9 11 9 13 9 0 12 13 4 2
9 9 9 12 13 4 11 10 13 2
10 9 2 9 7 9 13 4 9 10 2
12 11 9 7 9 0 0 9 13 13 4 3 2
4 10 13 4 2
4 13 9 9 2
13 9 9 13 4 9 9 2 7 14 4 15 13 2
14 9 10 3 13 2 9 14 13 9 12 9 13 4 2
4 3 13 7 2
8 9 13 4 9 0 9 0 2
9 2 13 9 0 12 2 3 13 2
9 3 9 9 0 13 11 7 11 2
22 12 7 12 9 9 2 9 10 13 4 9 2 9 9 9 0 13 4 7 14 13 2
7 9 10 9 13 9 13 2
7 11 14 4 3 13 11 2
10 12 10 12 9 3 13 4 9 9 2
13 9 9 7 9 13 4 2 7 9 9 9 9 2
13 0 2 7 2 0 9 9 9 13 2 11 9 2
5 3 13 4 11 2
17 12 9 0 9 10 13 4 9 9 7 9 9 10 13 13 4 2
6 9 13 13 13 9 2
13 11 11 9 9 2 9 7 9 13 13 13 4 2
21 0 2 7 2 3 9 13 4 13 4 2 7 8 3 13 4 2 9 2 10 2
15 2 3 14 4 10 13 2 7 13 4 13 4 9 2 2
14 9 13 13 3 2 7 9 10 14 0 13 4 11 2
12 9 2 9 2 7 9 2 9 2 13 4 2
9 9 9 9 0 13 14 13 0 2
7 11 7 11 13 4 9 2
19 9 10 13 4 2 13 4 2 9 2 3 2 12 9 13 4 9 9 2
19 10 13 13 4 13 4 2 10 10 13 7 13 2 7 9 0 13 4 2
11 9 13 4 12 9 12 9 0 13 13 2
12 3 9 10 13 4 2 3 9 13 13 2 2
16 11 11 9 0 13 4 10 13 2 7 0 9 0 13 4 2
16 2 0 9 13 4 2 7 2 9 13 12 9 15 9 13 2
5 11 13 10 9 2
6 15 14 13 9 0 2
12 13 9 13 9 12 9 13 4 9 2 11 2
17 9 10 2 9 9 13 9 3 3 13 13 4 11 7 11 9 2
9 2 11 9 13 4 9 13 2 2
7 11 11 9 13 4 3 2
6 2 9 0 13 2 2
5 9 12 9 13 2
19 11 11 11 0 13 9 13 4 3 2 9 11 9 12 9 13 4 7 2
11 13 13 9 13 10 13 4 7 3 13 2
23 3 13 7 9 13 4 2 13 2 7 3 13 4 12 9 9 2 7 9 9 13 4 2
11 12 9 13 2 3 13 4 9 13 9 2
30 11 3 13 4 9 2 3 13 4 11 13 9 2 7 11 3 13 4 9 9 2 7 11 0 12 9 13 4 9 2
13 11 9 2 12 9 9 2 14 13 3 0 9 2
8 13 4 9 11 13 4 9 2
17 9 0 12 9 10 2 11 9 9 9 0 9 13 13 13 4 2
8 11 13 7 12 9 13 4 2
14 9 9 13 9 9 9 9 13 13 13 4 11 9 2
24 15 9 13 3 2 9 13 4 9 0 13 2 7 3 13 4 3 11 11 9 9 7 9 2
8 12 3 14 4 11 15 13 2
11 9 0 11 13 3 2 13 9 13 11 2
5 14 13 10 9 2
9 12 9 10 13 13 4 11 7 2
5 11 11 9 13 2
8 9 10 9 13 9 0 13 2
14 11 2 12 9 10 9 13 2 10 9 10 13 4 2
13 2 9 13 9 13 13 8 0 13 2 3 2 2
8 14 13 3 0 2 13 4 2
12 11 13 4 2 15 0 2 9 3 13 4 2
21 10 13 7 2 9 9 9 12 3 13 4 7 9 13 4 9 13 9 12 13 2
16 9 3 13 4 2 0 7 13 2 9 7 9 3 13 13 2
10 9 9 13 13 15 2 9 0 13 2
11 11 9 13 4 12 9 2 11 13 9 2
17 9 2 3 2 3 13 7 9 2 13 4 2 9 13 4 2 2
8 7 2 9 9 13 13 4 2
7 0 9 13 4 11 9 2
17 11 9 11 11 9 9 13 4 2 7 3 13 4 9 10 11 2
13 10 9 9 13 13 4 2 7 11 9 13 4 2
10 9 0 9 13 2 7 2 9 12 2
11 11 9 9 13 13 4 3 11 2 12 2
22 11 9 11 11 13 4 2 9 10 13 13 4 11 11 11 13 4 9 2 9 2 2
3 9 13 2
8 11 3 13 4 13 4 11 2
22 10 9 2 12 7 12 9 12 9 13 4 3 9 0 9 13 9 9 13 9 9 2
8 11 12 9 12 9 13 9 2
9 3 11 7 11 9 9 13 4 2
21 11 2 11 2 11 7 11 2 7 2 9 12 9 9 9 12 9 13 4 13 2
15 9 0 2 7 2 9 13 4 10 10 9 15 9 13 2
16 15 10 9 13 4 9 13 2 7 9 13 13 9 13 3 2
9 2 9 13 4 9 13 4 2 2
8 11 9 9 0 13 9 13 2
10 11 11 9 7 9 13 13 2 3 2
5 11 3 13 4 2
9 11 0 9 13 7 13 13 4 2
13 3 3 2 12 9 13 4 9 0 13 4 9 2
5 2 15 9 13 2
11 9 12 9 13 4 3 9 9 12 13 2
25 12 9 10 9 9 0 10 13 4 2 7 9 9 13 9 13 4 2 10 13 4 10 13 13 2
4 3 13 4 2
14 11 9 9 7 9 13 4 7 0 13 4 11 9 2
13 11 13 4 2 10 9 13 9 13 13 4 3 2
12 11 8 11 9 9 0 13 13 4 12 9 2
6 12 9 9 13 4 2
32 9 10 2 7 2 7 9 13 9 9 0 9 2 9 0 0 13 4 9 9 10 7 10 10 9 0 13 4 9 9 7 2
24 12 9 7 9 10 13 4 13 2 7 12 9 9 0 13 4 11 2 7 9 13 4 9 2
15 0 9 9 14 13 7 2 9 13 4 9 9 0 13 2
8 7 14 4 0 13 13 4 2
9 11 11 13 4 9 2 12 13 2
13 12 9 0 9 13 4 9 0 9 3 13 9 2
5 9 13 4 3 2
15 9 10 9 10 2 10 9 13 4 10 9 13 0 9 2
8 9 12 9 13 9 13 4 2
10 7 2 10 11 13 4 9 0 2 2
17 11 12 9 13 4 2 7 0 9 0 13 10 9 2 12 2 2
16 11 14 4 13 2 11 9 10 13 7 11 13 4 9 10 2
10 7 2 9 9 9 7 9 13 4 2
16 13 9 13 7 13 2 9 13 3 9 7 9 0 13 13 2
5 10 13 9 15 2
8 3 12 9 13 13 4 9 2
13 11 13 9 3 13 4 11 11 9 9 10 13 2
8 12 9 13 9 0 13 10 2
7 9 12 13 4 12 9 2
9 9 9 12 13 7 12 13 4 2
12 11 9 13 2 9 2 13 13 4 11 11 2
8 9 13 9 14 13 0 10 2
7 2 9 3 13 4 3 2
7 13 4 10 13 4 9 2
16 11 11 8 11 2 12 2 12 13 4 9 0 2 11 9 2
11 9 12 13 2 13 13 11 9 12 13 2
9 7 2 9 0 12 9 13 4 2
19 7 2 10 9 13 4 7 9 13 4 2 9 13 11 9 9 13 4 2
7 12 9 13 4 9 3 2
15 9 13 4 9 9 0 2 7 9 0 13 4 9 10 2
7 11 9 9 13 9 10 2
23 11 9 12 13 4 11 9 11 13 4 2 11 13 4 9 11 13 4 9 13 4 7 2
19 7 9 0 13 9 13 7 13 9 13 3 14 13 9 2 13 3 13 2
17 3 10 9 13 4 2 7 2 9 13 4 2 14 13 9 0 2
24 9 9 12 9 9 2 9 0 2 13 9 2 9 0 10 9 7 9 9 0 2 13 4 2
17 9 0 7 9 0 13 9 13 4 7 2 9 0 13 4 11 2
11 11 9 13 4 11 9 12 12 9 9 2
16 9 9 12 13 4 3 2 7 12 9 9 9 13 4 9 2
27 0 13 4 0 9 0 13 2 7 14 13 3 0 2 3 7 9 0 13 11 9 9 9 12 9 9 2
8 9 0 14 13 11 10 2 2
11 0 9 13 4 2 9 0 0 13 4 2
6 13 9 0 13 4 2
8 10 9 9 10 13 7 11 2
5 2 9 0 13 2
20 7 2 9 13 13 9 2 9 10 9 9 13 4 2 7 9 9 13 4 2
13 11 12 9 9 7 9 10 13 4 3 9 0 2
8 2 11 9 13 4 11 2 2
19 3 13 2 7 9 9 0 9 13 2 9 10 7 12 9 13 13 4 2
4 9 13 13 2
16 9 9 9 0 3 13 2 7 13 3 9 13 3 13 4 2
11 9 10 13 9 13 9 13 9 9 12 2
11 2 13 4 7 13 4 9 12 0 2 2
10 9 13 4 2 9 9 7 3 13 2
7 11 9 13 13 4 11 2
24 3 2 9 9 9 9 3 13 4 9 9 9 13 9 2 7 3 0 13 4 11 7 11 2
17 0 9 9 3 13 4 2 7 3 9 12 9 13 4 9 0 2
12 9 9 2 9 0 13 9 2 13 4 11 2
15 9 10 2 9 0 12 13 9 13 2 10 9 13 4 2
6 0 13 4 11 9 2
8 13 4 12 9 7 10 9 2
7 9 13 9 3 0 13 2
9 9 9 7 9 12 13 13 4 2
7 14 13 15 9 10 13 2
20 9 12 9 9 13 4 11 9 13 2 7 2 12 9 9 7 12 9 9 2
10 11 7 11 9 0 9 13 4 11 2
12 9 13 14 4 2 9 9 10 9 13 4 2
7 9 3 3 13 13 9 2
13 12 12 9 13 13 3 13 11 7 11 3 13 2
16 9 12 13 4 11 2 11 13 0 4 12 9 7 12 9 2
15 9 0 9 12 9 12 13 4 3 11 9 2 11 9 2
10 2 15 9 9 9 13 13 4 2 2
20 7 9 3 13 4 2 7 13 4 2 9 9 2 9 0 9 12 13 2 2
6 15 13 4 9 9 2
21 11 9 9 9 13 0 12 13 4 2 9 10 13 4 9 13 9 12 9 9 2
9 9 2 13 9 12 9 2 3 2
20 2 3 14 4 0 15 9 10 13 7 9 7 9 9 10 12 9 13 2 2
19 9 2 3 2 9 0 2 7 9 9 13 4 13 4 7 9 13 9 2
19 0 13 2 7 2 11 13 4 9 0 9 0 9 9 0 13 13 4 2
19 11 9 9 10 9 11 9 9 12 13 4 2 7 11 9 13 13 4 2
20 9 12 9 0 13 13 7 13 9 13 9 9 9 13 13 4 12 9 9 2
10 2 7 0 9 13 2 15 2 3 2
9 11 0 13 13 4 11 9 12 2
6 2 9 9 14 13 2
10 3 13 4 9 0 9 0 0 13 2
12 2 3 9 9 13 4 9 9 0 13 2 2
11 9 13 11 14 4 15 13 13 4 11 2
17 9 9 13 2 11 11 11 9 13 2 3 13 11 9 0 13 2
12 9 7 2 13 9 0 13 4 13 9 0 2
6 10 13 10 9 12 2
22 9 9 2 12 2 13 4 9 13 9 13 2 7 14 13 12 13 2 10 13 4 2
16 7 9 14 4 0 9 13 2 9 9 11 13 13 4 9 2
19 9 10 9 7 9 13 4 2 9 0 7 9 9 0 7 0 13 4 2
18 9 0 10 9 0 12 9 12 13 4 2 9 10 4 13 9 0 2
9 11 9 13 7 9 9 13 4 2
7 11 13 0 13 4 9 2
12 2 13 4 3 2 9 9 9 9 13 2 2
7 2 15 3 3 13 4 2
9 12 9 13 9 0 13 13 4 2
7 7 3 13 4 9 9 2
7 7 2 9 13 4 9 2
9 3 13 4 15 9 0 13 4 2
17 3 2 11 9 10 13 4 11 2 11 9 7 11 13 9 13 2
11 7 9 9 13 9 13 2 9 13 4 2
10 7 2 12 9 13 7 0 13 4 2
6 2 9 13 13 4 2
10 3 15 9 3 13 13 9 13 4 2
6 6 2 15 11 13 2
6 9 13 4 3 11 2
5 12 9 13 4 2
4 14 4 13 2
10 9 10 14 13 9 9 13 4 9 2
7 9 9 9 13 4 13 2
4 9 13 4 2
4 9 13 4 2
25 12 9 13 4 9 2 7 11 9 0 7 9 13 13 4 9 9 13 13 4 9 13 13 9 2
7 11 9 9 7 13 9 2
19 3 14 4 3 13 9 0 12 2 14 11 14 11 2 7 10 0 13 2
7 2 9 13 13 13 2 2
9 11 7 9 13 11 9 13 13 2
10 13 15 13 13 4 2 15 13 11 2
10 9 9 13 9 13 2 13 3 10 2
15 9 9 13 9 9 13 13 2 7 10 9 12 13 4 2
22 9 14 13 13 2 7 9 10 9 13 4 11 7 9 10 13 4 2 3 2 11 2
8 2 9 10 13 3 13 4 2
3 9 13 2
18 9 0 0 9 10 11 9 13 4 2 9 9 2 13 4 11 9 2
18 11 11 9 9 13 13 4 2 9 12 2 11 8 11 2 11 2 2
6 11 12 9 13 4 2
8 2 0 13 9 13 2 11 2
7 0 13 2 9 0 3 2
7 12 9 9 12 9 13 2
20 12 9 9 13 11 9 2 7 2 10 13 3 2 9 13 10 9 9 0 2
25 10 2 13 4 2 9 2 9 2 13 9 13 2 9 11 13 14 4 9 0 2 10 9 13 2
5 11 0 3 13 2
22 9 14 4 14 9 0 9 2 14 9 13 13 4 9 9 0 13 14 4 9 0 2
7 3 14 4 11 9 13 2
16 11 9 9 2 13 2 11 7 11 11 13 4 11 7 11 2
15 0 9 10 13 4 9 9 7 9 0 0 13 4 13 2
15 9 9 0 7 9 0 13 13 7 9 9 7 13 4 2
13 9 10 2 11 2 11 7 11 13 4 9 2 2
8 9 0 13 9 14 13 9 2
9 9 7 9 9 10 13 9 13 2
6 3 12 9 13 11 2
14 3 2 11 9 2 11 9 7 9 0 9 13 13 2
16 11 9 9 0 13 4 2 7 12 9 9 13 9 13 4 2
17 2 3 13 13 9 13 2 3 14 4 9 3 10 9 13 13 2
12 11 2 13 2 2 9 9 13 2 11 10 2
11 9 13 13 9 2 9 13 7 9 13 2
8 11 2 7 2 9 0 13 2
10 9 14 13 2 7 3 13 4 2 2
9 7 2 9 9 9 0 9 13 2
13 9 13 4 10 12 9 2 7 12 9 13 4 2
5 10 9 13 4 2
10 9 10 9 0 0 9 13 4 11 2
10 9 13 2 9 10 13 4 9 9 2
22 3 14 13 2 9 15 3 9 0 7 0 13 4 2 3 9 13 4 9 13 4 2
6 11 14 13 9 10 2
5 15 13 9 13 2
36 3 13 13 2 13 2 3 13 4 9 9 2 9 0 14 4 10 3 13 2 2 7 14 13 2 9 9 9 0 2 10 10 13 9 15 2
17 0 12 9 13 13 4 12 2 7 9 10 12 9 13 4 11 2
14 10 9 2 11 2 9 0 2 9 13 13 13 4 2
13 9 7 13 13 4 2 7 11 13 4 0 9 2
8 11 9 13 9 13 9 13 2
13 11 11 9 0 12 9 13 4 11 9 4 9 2
10 0 14 4 9 7 9 0 13 9 2
4 15 9 13 2
12 11 7 9 13 13 2 7 3 9 13 4 2
14 9 0 13 4 2 7 2 9 12 13 3 13 0 2
13 7 9 9 7 13 2 11 13 2 9 11 9 2
15 2 11 3 9 0 13 2 7 9 7 3 13 9 13 2
28 11 11 9 9 9 0 13 2 7 0 13 7 2 9 2 9 7 9 2 7 9 9 0 7 9 13 4 2
10 7 3 2 10 9 13 9 13 15 2
23 0 2 0 2 0 11 11 9 13 4 11 0 9 9 2 12 9 13 0 13 4 7 2
7 2 15 9 13 13 4 2
8 11 9 10 9 8 0 13 2
6 9 9 7 9 13 2
12 11 7 11 9 2 9 9 12 12 9 13 2
19 9 0 9 9 2 12 9 9 9 13 4 2 10 9 13 9 13 4 2
9 11 9 12 9 13 4 9 10 2
8 3 2 13 9 13 4 3 2
10 11 9 13 9 10 9 2 12 9 2
13 9 13 13 9 13 4 2 7 9 14 13 13 2
15 11 13 4 2 7 9 10 9 11 7 9 0 13 4 2
9 9 10 12 9 11 11 0 13 2
12 12 9 13 4 12 3 11 9 13 4 9 2
12 11 10 2 7 9 13 4 9 9 13 4 2
7 11 9 12 9 13 4 2
13 9 9 12 13 2 9 7 2 7 13 13 4 2
8 3 9 3 13 13 9 13 2
14 13 13 4 10 9 13 2 9 2 9 2 9 2 2
6 10 13 4 9 10 2
8 9 9 9 13 13 4 0 2
7 11 9 9 0 13 4 2
15 7 2 11 11 9 14 4 13 9 9 9 13 4 0 2
12 9 9 0 12 9 0 13 4 9 0 3 2
6 9 0 13 15 9 2
5 9 9 13 4 2
14 3 13 4 13 3 2 9 9 13 2 9 9 13 2
4 15 13 4 2
20 9 9 9 10 13 4 9 13 2 10 9 13 13 9 13 10 9 0 13 2
8 9 9 0 13 9 13 11 2
17 11 9 9 9 13 13 4 7 11 0 9 14 4 13 13 4 2
21 11 9 0 13 2 9 9 10 10 13 4 2 7 3 7 13 13 4 10 9 2
8 2 0 10 9 13 9 12 2
14 9 9 12 13 4 9 0 7 9 13 4 10 9 2
4 10 13 9 2
7 9 13 13 4 15 9 2
9 3 13 9 2 7 13 13 4 2
13 3 13 4 9 10 10 7 9 10 13 4 9 2
10 9 9 2 9 13 13 4 12 9 2
13 3 12 13 4 2 12 9 13 2 12 9 2 2
3 3 13 2
12 9 10 3 13 4 7 9 9 10 13 4 2
23 11 0 9 9 2 2 11 9 0 7 0 13 2 7 11 7 11 9 0 13 4 2 2
6 2 11 13 13 2 2
6 7 13 4 9 12 2
6 9 10 13 9 13 2
5 9 10 9 13 2
9 9 7 9 13 9 9 9 0 2
8 11 9 13 3 9 13 4 2
26 9 13 9 11 11 2 11 9 2 9 13 12 9 10 9 13 4 9 2 3 13 9 12 13 4 2
11 9 9 12 9 13 4 2 9 7 9 2
15 9 0 9 2 9 12 2 7 2 9 9 0 13 13 2
7 9 13 7 9 9 13 2
9 14 13 9 2 3 9 9 13 2
8 9 13 7 9 13 13 4 2
7 9 9 0 13 13 3 2
33 10 13 13 2 9 0 7 9 9 9 13 11 11 12 9 9 12 13 13 4 2 3 13 12 9 2 11 9 11 9 9 9 2
14 15 9 2 14 13 10 7 9 9 9 13 9 13 2
13 9 9 13 9 9 13 4 2 11 13 4 9 2
12 9 0 2 7 2 14 4 3 9 0 13 2
12 9 13 0 13 2 7 9 14 4 13 2 2
8 11 13 4 2 11 9 13 2
15 9 13 3 2 10 9 3 13 4 9 2 9 9 9 2
13 9 13 4 13 7 3 13 9 9 3 13 13 2
19 2 6 2 9 13 4 7 15 9 15 13 4 2 14 2 10 13 4 2
28 7 10 2 13 9 13 9 14 13 11 7 11 9 13 4 9 2 9 13 13 4 9 7 13 4 9 7 2
15 7 3 3 13 13 3 14 4 10 13 13 13 9 13 2
6 3 13 4 2 7 2
11 12 9 2 9 12 7 9 13 10 12 2
5 10 13 4 9 2
17 9 2 7 2 3 13 4 14 4 0 13 2 11 9 13 10 2
7 12 9 13 3 13 4 2
10 9 13 13 4 7 9 12 13 4 2
7 13 4 0 9 9 13 2
6 9 10 9 0 13 2
23 9 9 13 4 2 7 9 2 3 0 2 13 4 2 7 9 9 14 4 13 9 13 2
8 11 14 4 11 11 11 13 2
9 13 14 4 14 4 15 13 2 2
13 9 13 9 13 11 9 10 9 0 10 0 13 2
14 11 2 7 2 12 9 13 4 9 2 9 13 12 2
7 11 9 9 9 13 4 2
11 3 10 9 7 9 13 13 4 9 13 2
5 2 12 9 13 2
11 7 2 9 2 9 7 9 3 9 13 2
12 3 12 13 4 12 9 13 2 12 9 2 2
18 9 13 0 13 2 7 9 0 2 3 9 15 9 9 0 13 13 2
9 3 9 2 9 9 13 4 3 2
15 0 13 7 2 15 13 4 11 9 10 13 4 9 13 2
9 11 9 12 13 4 2 9 0 2
10 10 4 7 2 9 0 13 11 14 2
16 0 13 4 9 9 10 7 3 13 4 2 15 9 9 13 2
10 2 13 9 13 10 13 4 2 7 2
17 9 10 11 9 13 4 3 10 13 3 0 13 13 4 11 11 2
14 9 13 4 9 0 2 15 9 9 9 12 13 4 2
8 2 14 13 3 9 0 9 2
21 3 13 9 9 13 4 2 7 12 9 3 13 4 9 12 2 9 9 13 4 2
13 9 9 9 13 4 9 2 7 10 9 12 9 2
5 9 12 13 13 2
21 0 13 4 12 9 2 7 2 9 8 10 2 9 12 7 10 9 13 4 9 2
15 9 13 12 9 0 9 2 12 9 9 7 12 9 9 2
26 12 12 9 9 0 13 7 2 11 11 11 0 14 4 9 0 13 9 0 11 9 9 12 13 11 2
14 9 9 13 4 9 13 9 13 4 9 9 13 9 2
9 2 14 4 9 0 13 0 9 2
17 7 11 9 13 9 0 13 4 11 9 2 7 9 0 13 4 2
5 9 13 13 4 2
8 3 11 10 3 0 13 4 2
10 7 9 13 4 9 3 13 9 10 2
4 11 13 4 2
15 0 9 9 0 12 13 4 2 7 14 13 9 0 2 2
14 9 9 9 13 7 9 9 13 4 2 10 12 13 2
16 9 13 2 9 9 9 13 4 2 7 3 0 13 9 13 2
5 9 0 13 4 2
11 12 9 9 13 11 7 12 9 0 13 2
9 12 9 13 4 7 9 13 4 2
10 11 11 9 13 9 9 0 0 13 2
7 2 14 13 15 13 4 2
12 9 7 9 13 4 2 9 10 9 13 4 2
12 2 7 3 14 4 13 2 3 13 9 13 2
10 3 9 10 13 7 11 13 9 13 2
9 11 11 13 9 13 13 4 11 2
18 11 9 3 13 4 2 14 13 3 13 9 9 14 13 9 12 9 2
14 9 12 9 13 4 2 7 0 13 4 3 9 10 2
13 11 3 13 9 2 2 3 9 0 13 4 2 2
5 9 9 13 4 2
6 10 7 9 13 13 2
14 15 3 13 4 2 7 13 4 10 3 13 4 15 2
11 9 13 13 4 2 7 13 3 13 4 2
7 7 9 10 3 13 4 2
12 9 9 13 15 9 0 2 3 13 10 13 2
12 15 9 13 2 3 13 4 15 9 9 12 2
5 2 13 4 2 2
6 0 13 15 13 13 2
21 10 2 9 9 9 2 0 2 13 4 2 7 2 9 9 9 12 2 13 4 2
7 9 13 2 0 9 13 2
15 12 9 13 9 13 9 7 9 0 13 2 13 9 9 2
14 2 9 9 13 4 2 10 13 4 7 3 13 2 2
22 2 9 9 10 13 7 2 0 13 13 4 9 13 9 13 2 10 13 14 4 2 2
10 0 13 4 2 7 12 9 13 4 2
4 13 4 9 2
11 3 2 12 9 9 11 9 10 13 4 2
7 9 9 12 9 13 4 2
15 9 0 13 4 9 12 9 2 7 9 10 13 4 9 2
10 10 2 9 0 9 13 13 9 13 2
25 10 2 9 0 13 4 9 0 9 13 4 9 9 13 4 2 7 12 9 0 3 13 4 9 2
7 9 0 7 13 13 4 2
18 2 9 0 14 4 13 9 2 7 9 7 9 14 4 9 13 2 2
11 11 11 9 2 7 2 12 9 13 4 2
13 2 13 9 2 3 2 9 7 9 9 13 2 2
11 13 13 4 7 3 10 12 13 13 4 2
6 14 4 9 9 13 2
10 2 11 2 9 2 13 9 13 2 2
19 9 0 7 0 13 4 11 12 9 13 9 2 7 3 13 9 13 4 2
10 15 13 9 13 7 3 13 4 11 2
26 9 2 9 0 11 2 13 13 4 9 10 11 2 7 9 10 13 3 2 9 9 13 13 13 4 2
7 9 9 9 3 13 4 2
13 9 10 13 9 13 4 2 3 13 4 9 13 2
16 13 9 13 12 10 9 0 10 13 13 3 2 9 13 12 2
14 2 11 11 9 13 4 2 14 4 15 9 13 2 2
5 2 9 0 13 2
12 9 0 9 9 13 4 2 9 7 9 14 2
3 3 13 2
10 3 13 4 0 9 2 9 13 3 2
10 3 13 9 7 9 0 9 13 4 2
7 10 9 13 9 13 10 2
22 11 13 4 9 0 11 9 12 9 2 3 2 12 9 2 12 9 7 12 9 2 2
6 11 9 13 2 13 2
12 3 2 9 12 13 4 9 9 9 13 4 2
3 13 4 2
9 12 12 13 4 3 9 11 9 2
8 9 9 13 2 14 13 9 2
19 10 9 0 13 4 9 7 2 7 2 9 10 9 7 9 0 9 13 2
25 14 2 9 0 9 13 2 7 2 9 0 0 12 13 9 13 2 7 9 13 3 3 13 3 2
15 3 12 9 13 4 7 12 13 2 9 9 12 13 9 2
5 12 9 13 4 2
8 9 12 9 7 12 9 13 2
5 14 13 0 0 2
9 9 7 13 13 9 13 9 13 2
7 11 11 9 3 13 4 2
16 11 2 7 2 9 10 9 12 13 4 9 9 9 9 13 2
10 9 10 13 4 3 2 9 0 13 2
6 9 13 13 13 4 2
6 10 7 10 0 13 2
19 11 9 9 9 12 9 13 7 3 12 9 13 7 10 10 13 4 3 2
10 3 2 9 0 13 9 0 13 4 2
16 12 9 13 2 7 13 13 9 9 13 9 13 4 9 13 2
19 9 2 9 13 13 9 9 12 9 8 0 13 9 9 9 14 4 13 2
8 7 15 10 9 13 15 13 2
10 9 13 7 2 9 13 9 0 13 2
15 7 3 2 11 9 13 13 4 2 11 10 13 13 4 2
6 2 14 13 13 9 2
12 15 14 4 9 12 10 13 0 9 12 13 2
10 9 0 9 0 13 8 0 13 10 2
13 7 9 14 13 4 13 2 0 9 3 4 13 2
3 14 13 2
5 9 2 0 13 2
5 2 9 13 4 2
32 2 15 13 4 9 12 9 12 9 13 2 0 9 12 13 7 9 12 9 13 3 13 4 2 7 14 4 9 10 13 2 2
17 14 13 2 7 15 9 3 13 2 13 9 7 3 13 4 2 2
9 2 11 9 9 0 9 13 4 2
6 2 13 4 9 2 2
7 11 9 7 9 9 13 2
9 14 4 3 13 11 9 13 13 2
14 13 4 11 12 9 0 13 4 2 13 2 13 4 2
18 9 13 2 11 13 4 9 2 9 0 11 13 9 9 9 12 13 2
14 11 9 2 7 2 11 9 13 9 0 13 9 13 2
7 11 14 4 9 9 13 2
6 3 9 13 10 13 2
10 11 9 9 9 12 9 9 13 4 2
5 2 9 13 4 2
10 14 13 9 0 15 2 0 13 4 2
5 15 9 12 13 2
16 11 9 9 9 13 4 3 7 9 13 4 12 9 9 9 2
12 9 2 11 2 11 11 9 9 13 4 9 2
9 9 12 9 9 3 13 13 4 2
5 9 0 9 13 2
10 9 12 11 13 10 9 9 13 9 2
3 10 13 2
13 3 13 4 9 2 7 11 12 9 9 13 11 2
13 3 13 4 9 2 12 10 13 9 7 9 13 2
11 11 11 13 4 2 7 9 9 13 4 2
16 3 13 4 3 11 11 9 11 11 7 9 0 11 11 11 2
10 10 10 0 2 7 2 9 13 4 2
5 2 13 7 13 2
8 2 9 7 9 0 14 13 2
6 9 14 4 3 13 2
9 9 0 12 13 9 13 0 13 2
20 11 14 13 9 13 4 11 2 7 9 9 9 13 14 4 9 13 13 4 2
5 7 9 10 13 2
11 2 9 3 0 13 2 7 14 13 13 2
13 3 2 9 9 13 9 9 12 9 13 13 4 2
11 10 9 2 11 11 13 4 10 13 4 2
6 3 13 4 9 13 2
4 9 13 9 2
5 12 9 13 9 2
8 3 3 9 0 13 4 11 2
11 2 9 13 4 2 10 13 4 13 2 2
18 2 11 13 2 3 2 9 3 13 2 9 7 11 13 7 11 2 2
15 11 2 11 7 11 3 13 4 10 9 9 13 0 9 2
16 9 9 0 13 13 4 7 2 14 4 9 10 13 9 0 2
14 9 15 13 13 13 7 9 14 4 9 0 13 13 2
5 3 13 4 9 2
28 9 13 9 9 10 13 9 13 4 2 9 2 9 0 2 9 9 2 7 3 10 9 0 7 0 13 4 2
8 9 13 4 9 13 4 11 2
14 2 3 13 4 0 9 9 2 9 0 12 13 7 2
6 11 9 13 13 4 2
10 15 3 13 12 9 13 4 9 13 2
10 10 13 9 13 3 3 12 9 0 2
17 11 9 2 2 11 9 9 13 4 13 13 9 13 11 11 2 2
11 11 13 9 12 9 2 7 10 0 13 2
14 11 11 9 13 0 13 2 7 11 0 13 4 9 2
12 9 0 3 11 13 4 2 12 2 9 13 2
5 10 0 13 2 2
16 9 9 3 13 13 3 11 9 0 2 2 3 2 13 9 2
22 11 9 13 4 9 3 2 11 11 9 2 7 2 9 2 9 13 13 4 12 9 2
5 9 9 13 4 2
8 9 0 13 9 0 13 4 2
10 7 0 10 13 4 9 9 7 9 2
7 9 9 7 9 13 4 2
21 9 0 9 13 2 9 2 13 7 11 2 9 10 2 9 13 4 13 4 11 2
17 12 9 11 9 13 11 9 13 2 7 10 12 11 9 13 11 2
8 12 9 13 4 11 2 11 2
10 9 0 2 11 9 7 9 13 4 2
21 11 2 12 5 2 2 11 2 12 5 2 7 11 2 12 5 2 9 13 4 2
8 11 11 13 2 9 12 13 2
9 10 9 13 11 13 4 13 9 2
15 7 11 9 9 1 2 9 13 9 9 13 13 13 4 2
8 9 10 3 4 13 9 13 2
19 3 2 7 2 13 13 4 10 13 13 7 9 1 13 4 9 9 10 2
12 9 2 9 1 13 2 9 7 9 1 13 2
10 9 11 9 0 7 0 13 4 9 2
27 9 3 13 13 4 2 12 9 3 2 7 3 9 0 13 14 4 2 13 7 0 9 13 4 12 9 2
14 9 13 9 13 2 7 10 10 13 4 11 1 2 2
14 2 9 1 9 13 4 2 9 0 2 11 7 2 2
21 9 1 13 4 9 7 9 13 13 7 9 9 2 10 13 4 9 1 13 4 2
15 11 9 9 0 3 13 9 0 13 3 2 9 7 2 2
14 15 15 1 0 13 4 2 3 9 2 9 2 3 2
6 9 3 9 13 9 2
17 9 9 0 12 2 7 2 10 9 3 9 13 4 12 9 3 2
20 11 2 7 2 3 13 4 9 2 7 11 9 13 9 13 2 9 13 4 2
14 11 13 13 3 3 13 4 12 9 2 12 7 11 2
15 11 13 2 9 1 2 9 2 13 4 12 9 12 12 2
24 11 13 4 12 9 10 9 9 11 9 13 4 9 12 9 7 9 13 4 9 1 9 13 2
19 10 1 2 7 2 11 11 9 13 4 9 2 10 10 2 8 11 11 2
20 9 9 7 11 9 13 13 4 9 12 2 7 2 9 2 3 2 11 11 2
9 11 11 11 9 14 4 0 13 2
14 3 7 11 9 13 2 7 11 7 11 13 4 13 2
16 11 9 2 7 2 10 9 12 13 4 9 9 9 9 13 2
21 2 2 11 11 2 9 9 9 13 9 9 2 3 3 9 0 13 13 13 4 2
22 11 9 13 10 9 12 11 11 9 12 9 9 13 13 4 11 11 9 9 13 9 2
12 11 11 3 12 9 9 9 9 9 13 4 2
16 12 9 0 13 13 13 7 2 14 13 10 1 13 4 0 2
21 9 9 2 9 9 12 2 13 13 4 2 7 9 10 2 0 2 13 13 4 2
8 2 0 11 9 13 4 13 2
17 11 9 11 9 13 0 13 9 13 9 13 2 11 3 13 4 2
19 12 9 9 12 13 4 9 9 11 2 9 11 9 2 7 9 13 4 2
10 7 2 12 1 13 12 9 9 9 2
24 13 9 1 2 9 9 2 13 13 4 10 9 13 4 11 11 11 12 9 12 7 12 9 2
21 11 0 2 2 9 10 14 13 11 15 13 9 2 7 9 1 10 13 0 2 2
14 12 9 14 4 0 13 2 7 13 9 10 13 4 2
20 0 9 10 13 4 9 1 9 7 11 13 12 9 1 9 12 13 3 13 2
11 11 1 13 13 12 9 9 13 4 11 2
13 11 9 11 9 11 13 9 10 9 13 4 11 2
20 11 11 9 2 7 11 11 9 13 4 9 11 13 4 11 9 9 9 9 2
19 11 11 9 13 4 12 9 13 2 11 9 13 4 11 11 11 9 13 2
15 11 9 9 13 4 9 12 2 7 11 7 13 4 13 2
24 2 9 1 2 9 0 12 13 9 13 10 10 2 7 10 0 13 0 9 10 13 13 2 2
19 9 13 13 4 12 9 9 12 13 2 9 11 9 11 1 13 9 13 2
22 11 9 13 4 11 9 13 2 7 9 14 4 9 13 7 9 9 13 9 13 4 2
18 10 10 9 1 2 11 13 9 2 11 13 3 2 11 11 13 4 2
19 3 3 3 13 13 9 2 7 13 4 15 9 9 12 3 13 13 4 2
19 11 12 9 13 9 10 9 13 7 3 13 2 9 10 13 9 13 7 2
23 12 9 3 7 3 13 4 2 3 7 3 2 9 9 13 2 9 15 8 3 13 9 2
28 10 1 9 13 4 11 2 11 9 9 7 9 0 2 0 9 11 9 7 11 9 10 7 9 13 4 13 2
20 9 12 9 9 13 13 4 2 7 9 12 9 2 12 12 9 7 12 9 2
7 2 7 11 9 3 13 2
12 11 7 9 9 10 4 13 9 9 13 13 2
17 9 13 9 13 2 9 11 11 7 11 11 9 9 9 13 4 2
12 15 13 2 3 2 9 1 9 9 13 4 2
17 11 11 12 9 9 9 12 9 13 4 11 0 9 3 9 1 2
12 13 3 13 2 7 9 3 14 13 3 3 2
13 9 3 13 4 9 9 9 13 2 7 3 14 2
15 3 9 12 9 1 9 13 13 4 2 9 0 14 13 2
16 13 2 3 14 13 9 15 10 9 9 12 9 9 13 4 2
11 9 9 9 4 7 12 1 9 13 4 2
21 14 4 11 9 9 0 13 2 11 11 9 1 11 11 7 11 13 4 2 7 2
17 11 9 9 9 9 11 11 9 13 4 2 11 9 14 13 0 2
9 12 13 4 9 11 7 11 1 2
7 2 11 1 13 4 2 2
13 11 9 9 4 13 9 13 9 2 9 13 9 2
21 11 9 7 9 2 3 13 7 2 3 13 4 9 0 9 13 7 9 9 0 2
13 11 2 11 7 10 9 1 9 2 13 13 4 2
20 11 11 7 11 11 4 13 13 9 9 10 2 7 9 1 13 12 12 9 2
11 7 10 9 13 9 7 9 2 9 1 2
8 7 2 12 1 13 3 13 2
13 9 0 9 13 4 11 2 11 1 7 11 1 2
21 13 12 9 9 13 13 11 11 9 9 12 2 7 10 1 9 13 13 4 3 2
19 11 10 9 13 4 12 9 10 10 9 2 9 0 3 14 13 0 13 2
13 9 9 1 2 7 2 11 13 3 13 4 11 2
30 9 9 1 2 9 0 2 13 9 10 2 9 9 9 3 2 7 11 11 11 9 13 13 4 2 9 12 13 3 2
19 11 10 9 13 9 0 13 3 11 9 2 11 9 0 13 4 3 9 2
23 9 1 13 9 2 11 11 9 1 13 4 9 7 7 2 9 9 3 1 13 4 3 2
14 10 9 1 13 13 7 2 3 1 14 4 9 13 2
19 12 9 0 13 3 2 0 9 13 4 12 9 2 7 3 13 4 11 2
10 2 14 4 3 0 13 2 11 11 2
16 12 9 10 13 4 9 9 12 9 2 15 0 13 14 4 2
14 0 13 10 3 9 0 13 7 13 13 12 12 13 2
23 11 11 9 11 13 4 11 9 2 7 10 9 13 11 11 11 0 9 13 11 9 9 2
19 9 2 11 1 9 9 9 2 11 9 10 0 9 13 7 0 13 4 2
11 11 3 13 4 3 11 1 9 13 9 2
25 11 9 11 11 12 9 11 9 0 0 9 13 13 2 7 9 10 2 0 9 9 0 0 13 2
15 10 9 13 4 2 7 9 1 9 10 9 13 13 4 2
21 11 11 13 4 11 13 2 7 11 3 0 13 11 2 7 14 4 9 0 13 2
15 3 10 13 9 13 9 14 13 10 0 9 13 4 9 2
8 10 9 2 3 13 9 13 2
26 10 2 0 9 9 13 13 4 2 10 10 9 7 9 1 13 2 10 9 0 7 9 9 13 4 2
13 9 7 9 11 9 13 13 4 9 13 4 13 2
19 9 10 9 9 9 9 1 9 13 4 7 15 1 9 13 4 13 4 2
10 10 13 4 2 14 4 11 11 13 2
9 2 11 11 13 15 9 0 2 2
25 7 2 13 9 10 1 9 7 9 0 0 9 7 9 10 9 13 4 2 9 2 0 2 13 2
24 7 2 3 11 13 9 9 9 9 13 4 12 12 11 7 14 4 13 3 0 9 13 4 2
31 2 12 9 1 9 9 12 13 2 13 13 9 13 13 9 10 9 13 4 2 9 3 13 4 13 10 9 7 9 2 2
10 15 7 0 13 13 2 7 14 10 2
13 2 9 9 0 13 4 7 9 3 0 13 4 2
20 9 9 9 9 8 9 0 13 4 9 2 14 4 3 8 9 7 9 13 2
30 3 13 4 11 9 10 13 9 2 7 2 10 1 2 12 9 9 13 4 9 2 11 9 1 13 4 11 12 9 2
16 9 10 1 2 11 13 13 7 9 1 9 12 13 4 13 2
25 2 9 9 9 13 13 4 2 7 9 13 9 1 9 9 10 15 9 9 13 4 13 4 2 2
15 7 2 9 9 13 9 12 13 4 13 4 3 11 9 2
9 11 11 11 11 12 12 9 13 2
15 3 2 15 9 13 11 11 2 7 0 13 4 10 9 2
22 2 9 2 9 2 0 7 9 2 9 13 4 3 11 11 11 3 11 13 9 13 2
19 10 2 9 13 2 9 0 9 1 9 13 9 2 9 2 13 13 4 2
14 9 2 9 2 13 12 9 1 9 13 12 9 0 2
16 2 11 7 11 13 13 4 2 9 11 13 4 9 0 12 2
23 7 2 11 7 11 1 3 9 13 13 4 9 2 9 9 13 4 13 4 2 9 0 2
18 9 10 13 13 9 10 2 15 0 13 2 7 3 3 2 3 0 2
17 11 11 9 9 0 1 13 4 13 4 9 0 1 13 9 9 2
20 9 9 2 11 11 3 13 9 13 11 11 2 7 14 13 9 9 9 0 2
13 9 13 7 3 3 13 13 9 10 13 4 3 2
5 9 13 2 13 2
23 12 7 12 9 13 3 11 9 13 12 9 2 12 9 9 13 4 2 11 2 12 2 2
13 9 9 9 7 9 9 9 9 9 13 9 13 2
21 9 9 12 13 4 3 9 2 7 10 3 13 4 11 0 7 11 2 11 2 2
31 9 13 12 9 0 12 13 4 3 11 11 9 2 11 11 7 11 9 1 2 7 13 12 9 13 4 2 10 12 9 2
19 9 13 3 2 14 13 11 0 2 7 12 13 2 7 12 9 10 3 2
11 11 11 9 11 13 4 7 11 13 4 2
26 12 9 9 13 11 1 2 11 2 12 2 2 7 9 12 9 13 4 2 13 4 9 9 13 4 2
14 11 9 3 13 4 7 2 11 11 9 3 13 4 2
10 12 10 2 14 13 10 9 13 9 2
17 0 9 1 11 13 4 9 3 3 13 4 3 11 11 0 9 2
11 9 0 13 13 9 7 15 9 9 13 2
10 7 2 9 12 13 4 11 9 9 2
21 9 9 9 13 13 9 2 9 9 7 9 7 9 13 9 0 13 13 13 9 2
41 9 12 13 3 9 0 2 13 2 13 4 11 11 9 9 2 7 3 2 9 9 11 13 13 2 7 9 9 1 13 4 13 4 2 2 9 9 1 13 2 2
20 11 11 2 12 2 13 13 4 11 11 11 1 2 12 2 12 7 12 2 2
24 11 11 11 13 9 11 11 13 4 13 4 10 2 7 9 10 11 9 3 13 4 11 9 2
12 9 0 13 9 11 2 9 9 3 13 4 2
13 14 4 15 13 9 0 13 0 9 7 9 1 2
9 11 13 4 12 12 9 7 3 2
15 9 1 9 9 13 11 9 2 3 3 14 13 7 2 2
7 10 9 14 13 13 13 2
14 9 13 2 9 7 9 2 13 4 11 11 11 9 2
11 11 9 13 9 13 9 13 11 9 0 2
16 9 13 2 10 9 1 2 13 13 4 9 3 7 9 13 2
11 11 11 11 10 9 13 4 2 11 0 2
19 9 9 1 13 4 11 11 9 2 7 9 9 12 9 10 9 13 4 2
9 11 11 13 4 12 9 11 1 2
10 11 7 10 12 9 1 9 13 4 2
23 11 9 2 9 9 9 1 13 3 2 9 0 12 9 13 4 9 9 10 13 13 4 2
19 11 9 1 2 3 0 13 9 10 12 1 3 13 9 9 9 13 4 2
18 11 2 7 2 11 0 13 9 13 11 9 2 9 9 2 13 4 2
22 11 11 9 9 13 4 3 2 9 9 2 7 13 4 10 9 11 11 3 13 13 2
10 9 12 9 12 13 4 11 11 9 2
20 7 9 10 3 13 4 2 9 13 4 9 2 9 3 13 4 9 9 13 2
13 2 3 9 13 2 12 7 3 13 0 13 4 2
9 7 10 1 2 10 10 13 4 2
11 3 12 9 13 4 2 7 10 10 3 2
9 2 15 12 9 13 9 2 11 2
15 10 10 1 2 9 9 11 9 9 13 4 2 11 11 2
10 9 0 9 1 12 9 13 4 11 2
18 7 9 11 12 9 11 11 13 4 13 13 3 12 9 13 4 9 2
14 13 9 0 13 4 9 12 13 13 4 9 0 12 2
10 9 9 1 2 11 9 9 13 4 2
27 2 0 9 9 9 10 13 9 13 13 4 2 7 9 13 9 9 9 0 10 13 10 14 4 13 2 2
8 11 13 4 12 12 11 11 2
11 9 0 11 13 4 11 11 7 9 9 2
30 9 9 13 9 7 9 3 13 4 2 7 3 7 3 13 4 9 0 13 4 9 9 9 0 13 4 9 9 8 2
28 9 0 9 14 13 9 10 2 11 11 9 9 12 13 4 3 14 4 13 9 9 1 13 0 4 9 13 2
21 9 10 13 2 7 2 11 9 1 9 0 13 9 0 2 12 9 0 13 4 2
10 9 13 7 12 9 3 13 9 13 2
18 11 10 0 13 4 3 2 7 3 3 2 7 14 3 9 9 0 2
17 11 13 4 14 13 9 10 10 9 11 11 2 0 13 13 3 2
10 9 9 12 11 13 9 13 4 13 2
31 3 7 9 13 7 0 10 1 10 0 14 4 13 2 14 13 10 2 0 9 13 9 3 13 4 13 9 7 13 9 2
8 11 9 10 13 4 11 1 2
11 10 1 2 9 9 13 9 13 13 4 2
30 9 11 9 9 11 11 3 13 4 9 9 13 2 9 0 2 2 7 11 9 9 11 11 2 0 2 13 4 9 2
13 11 9 9 0 9 9 13 9 13 9 13 11 2
7 10 9 1 13 13 4 2
5 10 13 8 13 2
18 9 0 13 4 11 2 7 2 10 9 13 4 2 9 13 13 4 2
17 11 2 13 9 11 11 1 13 9 13 9 0 13 4 2 7 2
17 13 4 2 0 13 4 10 9 9 9 9 1 2 7 9 0 2
18 11 11 11 11 9 9 13 4 9 0 11 9 2 13 2 4 13 2
7 9 1 9 9 9 13 2
17 2 13 4 10 9 13 2 9 10 13 3 9 0 13 9 13 2
14 9 0 13 4 11 11 2 7 3 3 13 4 9 2
17 9 9 12 9 0 7 9 12 13 2 9 1 9 7 9 13 2
28 7 2 9 7 9 9 0 13 7 2 9 0 10 0 13 2 3 3 2 9 2 9 0 9 7 9 9 2
15 9 12 13 9 13 2 7 3 13 13 12 1 13 4 2
26 7 2 14 4 9 0 13 11 2 11 11 9 9 13 13 4 12 9 12 9 11 13 9 12 1 2
14 3 3 13 4 9 2 3 3 13 13 9 13 4 2
12 9 10 13 4 9 0 7 0 9 0 13 2
6 11 11 0 13 4 2
18 2 9 9 13 4 2 7 3 9 12 3 9 13 2 7 11 1 2
19 10 2 11 9 3 13 4 3 10 13 11 11 7 11 11 13 13 4 2
13 9 12 1 2 9 12 9 13 7 9 13 13 2
22 11 7 12 1 13 4 9 7 2 9 2 11 9 9 0 13 4 2 9 9 13 2
17 9 12 9 13 11 9 10 3 13 13 4 15 10 13 3 13 2
15 11 9 13 13 4 0 10 2 3 2 7 13 3 13 2
7 3 12 13 13 4 13 2
13 9 14 4 0 13 2 15 9 1 13 4 9 2
13 9 3 13 4 13 13 2 9 13 0 15 2 2
8 3 1 12 12 9 13 4 2
18 11 11 13 4 2 7 9 13 9 11 13 4 2 11 11 3 0 2
28 10 9 13 4 9 0 0 13 4 9 13 4 10 9 13 2 7 14 9 13 2 3 1 13 4 9 2 2
8 3 11 13 4 7 3 11 2
24 0 9 9 9 9 12 13 2 7 2 9 1 13 12 9 9 9 12 13 4 13 4 11 2
26 9 1 9 9 7 9 1 13 4 9 13 4 11 11 11 9 3 9 10 9 2 11 13 9 0 2
30 2 9 9 1 0 13 7 9 13 13 9 2 9 2 9 2 9 2 9 2 9 7 10 9 7 9 0 7 0 2
12 2 9 0 9 9 1 15 9 13 13 4 2
15 12 9 1 13 13 4 2 9 13 4 9 13 9 1 2
12 15 9 2 11 11 7 11 13 4 0 9 2
27 11 11 11 9 9 2 11 12 9 11 11 7 11 9 0 9 9 11 11 9 2 9 9 2 13 4 2
16 11 11 13 4 9 1 11 9 0 13 2 0 9 0 13 2
8 2 9 13 4 11 1 9 2
18 9 13 9 10 13 2 10 3 13 13 4 2 7 0 13 13 4 2
19 7 2 9 10 2 9 13 9 3 1 13 4 2 7 10 7 0 13 2
9 7 9 0 13 4 2 0 9 2
32 11 11 11 11 9 13 9 13 4 13 11 14 4 3 13 9 13 4 2 7 7 11 2 9 7 9 9 3 13 13 4 2
17 9 3 2 12 9 9 12 13 4 7 9 0 13 4 9 13 2
15 3 13 4 11 9 9 12 11 11 9 11 2 11 2 2
20 11 9 9 9 12 13 4 2 11 14 13 9 7 9 9 13 9 13 4 2
16 9 0 10 9 13 4 2 3 2 3 9 0 0 13 13 2
19 11 11 13 4 14 4 11 11 13 9 13 7 9 7 14 4 13 13 2
27 9 10 11 9 11 11 13 4 0 9 2 12 9 2 9 0 2 9 9 13 7 13 9 13 13 4 2
24 15 9 1 10 13 9 12 10 13 13 2 12 9 9 0 13 9 0 13 2 3 7 3 2
12 9 10 9 7 13 4 2 9 12 9 2 2
18 10 9 2 2 9 0 12 13 15 9 9 9 0 13 4 13 2 2
30 3 2 7 2 12 12 9 11 11 7 11 1 9 3 0 13 2 7 2 9 1 2 12 10 13 4 9 9 10 2
9 9 9 0 12 13 4 9 1 2
15 2 9 1 9 13 4 2 7 13 13 13 4 9 2 2
13 12 9 12 9 9 13 4 9 9 7 9 13 2
15 11 11 7 3 13 4 9 9 9 14 4 9 13 13 2
18 9 9 2 9 7 9 2 13 3 2 9 9 1 2 9 9 0 2
15 11 13 3 3 11 9 9 14 13 9 3 13 12 9 2
14 12 9 9 1 12 9 13 4 3 9 11 9 0 2
21 9 13 4 9 1 2 3 14 4 13 9 0 7 0 2 7 13 13 0 13 2
21 9 12 3 9 0 13 2 9 13 13 0 9 1 2 9 0 13 4 10 1 2
18 9 9 9 0 13 9 13 9 2 11 11 9 9 13 4 12 9 2
17 3 9 13 4 12 9 13 4 2 7 9 14 4 3 3 13 2
21 3 9 2 13 9 9 7 9 1 9 0 13 4 12 2 3 12 9 13 4 2
13 9 10 2 7 3 9 2 13 13 4 9 10 2
14 11 13 9 11 9 13 9 1 11 10 9 13 4 2
14 11 11 14 13 9 2 7 11 11 13 4 10 9 2
24 2 13 4 2 9 10 11 13 4 7 9 12 9 13 2 3 13 9 13 2 11 1 2 2
17 9 0 12 1 2 10 9 8 0 13 9 3 13 4 3 13 2
17 9 11 9 10 13 4 12 9 2 7 10 13 4 11 9 0 2
23 11 11 11 9 9 13 4 9 2 2 11 13 9 13 4 3 2 7 14 4 13 2 2
16 12 9 1 13 4 9 3 9 2 9 2 7 9 0 13 2
5 13 3 3 13 2
11 9 10 10 2 3 12 10 10 13 4 2
18 9 2 11 11 0 13 2 7 13 11 9 7 9 0 13 11 13 2
12 3 2 12 9 2 11 7 0 1 13 4 2
7 9 0 1 9 13 4 2
17 11 11 13 4 12 9 12 13 4 3 9 9 2 12 9 13 2
11 12 1 2 3 2 12 9 9 13 4 2
14 11 7 11 13 13 4 9 3 3 9 0 12 9 2
7 9 7 9 1 9 13 2
25 11 7 11 10 9 13 10 2 9 7 9 9 13 13 9 13 13 9 13 13 9 7 9 10 2
31 3 2 13 9 13 4 7 2 12 9 11 11 9 9 9 13 11 11 2 11 1 3 7 2 12 9 9 12 13 13 2
30 11 11 9 0 11 11 13 7 11 11 13 11 9 12 9 13 4 2 14 9 7 9 2 3 7 3 11 11 9 2
10 3 1 2 9 0 13 4 9 1 2
17 11 11 3 13 9 13 9 13 7 13 9 13 2 0 9 13 2
18 9 10 9 2 11 9 3 9 13 7 3 1 9 13 4 9 1 2
15 11 0 9 2 11 11 2 7 2 9 0 13 3 13 2
39 9 9 13 2 9 13 4 9 9 13 4 9 2 11 13 4 9 10 2 9 0 2 13 4 11 7 11 1 9 7 2 9 2 9 9 13 4 11 2
7 9 0 10 1 13 4 2
18 3 2 11 11 9 13 4 11 13 2 13 4 9 11 9 13 9 2
23 9 9 7 9 0 13 7 13 4 2 0 9 0 7 0 2 9 9 7 15 9 1 2
22 9 9 0 11 9 13 9 13 9 13 2 7 9 14 4 9 13 9 9 13 9 2
13 9 0 9 0 1 2 12 9 13 4 10 13 2
21 11 11 9 13 9 1 9 13 0 13 4 11 2 7 3 13 4 11 7 11 2
16 9 1 2 9 0 13 4 12 9 1 2 9 13 9 13 2
17 3 2 10 12 9 13 4 9 3 9 7 9 0 13 9 13 2
7 7 11 7 11 9 13 2
14 11 9 7 9 3 13 9 13 11 9 9 9 1 2
17 12 9 9 9 13 4 2 7 11 2 7 2 9 7 9 2 2
27 2 9 13 13 9 0 13 13 4 11 9 2 7 2 7 2 13 4 11 0 7 0 13 9 13 2 2
24 3 13 13 9 2 7 2 13 4 9 2 7 9 14 13 3 3 2 14 7 9 9 9 2
13 9 12 13 4 3 3 13 2 7 9 13 4 2
21 9 0 9 9 3 0 13 2 7 0 13 4 9 9 12 13 7 9 9 13 2
18 9 13 4 2 9 9 10 13 9 1 7 13 9 7 3 13 4 2
20 3 11 11 7 11 11 9 13 4 2 7 9 9 9 1 9 0 13 4 2
9 2 7 2 14 4 3 7 13 2
16 11 9 11 9 12 9 9 13 4 9 0 13 9 12 13 2
24 11 2 7 2 3 1 12 7 9 13 4 9 13 14 4 13 13 4 2 7 3 13 4 2
25 11 13 4 9 0 11 2 11 7 11 9 9 13 0 13 9 1 9 9 13 2 9 0 2 2
27 11 13 11 9 9 1 0 9 10 2 7 3 11 7 11 9 13 14 4 2 9 10 13 4 3 7 2
22 10 1 2 11 2 11 2 11 2 11 2 11 0 7 10 10 9 9 13 9 13 2
11 3 3 13 4 2 9 2 9 13 10 2
14 12 7 10 2 9 10 13 4 9 10 2 9 1 2
7 9 11 9 7 0 13 2
14 9 9 0 9 9 13 4 2 3 3 13 7 9 2
13 9 10 13 9 10 7 3 3 13 4 13 4 2
20 10 13 13 2 3 9 10 12 13 4 9 2 7 12 13 4 10 9 13 2
10 11 9 0 9 13 2 11 9 1 2
14 11 9 7 9 0 9 9 1 9 13 4 12 9 2
17 2 9 1 13 9 9 0 7 0 2 3 13 4 3 9 9 2
20 11 11 11 9 9 7 11 9 9 11 11 11 11 1 9 13 13 4 3 2
21 9 12 13 4 10 1 2 9 2 9 0 2 7 9 9 9 12 13 4 9 2
12 7 10 13 3 9 0 13 4 9 10 1 2
11 11 11 9 11 13 9 2 11 0 13 2
12 11 11 9 13 4 11 9 13 4 12 9 2
9 11 11 10 9 13 4 9 12 2
8 12 9 13 2 7 9 3 2
22 12 12 9 10 11 9 13 9 0 7 0 1 11 9 11 13 13 4 9 10 3 2
19 9 14 4 3 10 9 9 10 13 2 9 9 3 9 9 0 13 4 2
18 7 2 11 9 10 9 9 9 13 13 13 7 0 13 4 11 9 2
17 11 1 9 12 9 7 11 9 9 10 12 9 13 13 4 11 2
12 3 9 9 0 13 4 2 9 9 9 1 2
7 12 11 11 13 4 9 2
12 0 10 2 11 9 1 9 0 9 12 13 2
11 10 10 13 4 9 2 9 1 13 4 2
21 9 0 13 13 4 3 9 9 9 9 13 2 7 9 7 13 13 4 11 9 2
13 11 9 9 9 0 13 4 11 11 11 9 0 2
15 7 2 9 10 9 13 9 0 13 4 13 13 4 11 2
18 9 13 4 11 11 9 9 2 7 11 9 13 4 9 13 4 13 2
24 3 13 9 13 2 9 13 4 2 9 14 13 7 2 3 13 11 12 9 9 13 4 13 2
11 9 7 9 9 13 4 9 0 9 13 2
20 9 13 3 3 1 2 9 1 7 9 13 3 13 9 12 1 13 4 13 2
19 11 13 13 4 11 9 2 7 0 12 9 14 4 14 9 7 3 13 2
12 9 3 12 10 11 9 9 12 13 4 9 2
13 10 11 13 9 12 1 7 9 13 9 13 11 2
9 11 11 13 4 3 1 10 9 2
10 13 7 2 15 10 9 13 15 13 2
13 9 13 13 4 7 9 12 1 10 9 13 4 2
9 3 3 2 6 2 0 13 4 2
22 9 0 13 4 2 3 0 13 7 14 4 3 7 13 9 10 12 9 13 4 3 2
11 9 10 12 9 11 11 13 2 12 9 2
10 11 2 9 1 13 2 9 13 4 2
19 11 1 2 9 0 1 9 13 0 9 11 7 11 11 9 0 3 13 2
19 9 3 1 0 13 13 4 2 7 3 7 2 3 2 13 13 4 13 2
21 10 9 13 4 2 9 10 9 2 9 13 13 9 13 11 9 0 13 4 9 2
27 9 9 10 2 0 7 0 2 3 0 2 11 9 13 4 9 13 2 14 4 2 7 2 15 9 13 2
29 3 9 12 10 9 10 9 13 4 13 9 9 13 4 9 9 13 9 12 2 7 9 10 7 11 9 13 4 2
16 12 11 9 9 11 9 12 9 9 13 4 11 2 9 0 2
17 9 12 13 13 4 3 11 11 9 2 11 9 11 9 13 4 2
13 11 13 4 9 13 4 11 11 9 11 11 9 2
10 3 9 13 2 9 9 13 7 9 2
20 9 1 11 13 4 9 13 4 11 2 7 10 1 15 13 4 13 9 0 2
15 7 2 3 7 2 13 4 9 9 13 3 9 13 4 2
16 9 9 9 9 7 9 9 9 13 9 7 9 13 9 13 2
24 11 9 2 11 2 9 9 11 1 9 9 10 13 4 11 9 3 11 2 11 2 13 9 2
15 11 9 9 12 13 4 2 7 11 7 11 11 12 9 2
19 9 0 9 9 13 0 1 13 4 2 7 11 7 11 9 0 13 4 2
14 3 9 10 13 13 2 9 14 13 2 7 9 1 2
13 11 9 11 9 12 11 9 11 9 13 4 9 2
23 2 9 9 7 9 13 4 9 7 13 4 7 10 1 9 7 9 9 13 0 13 2 2
12 12 9 13 4 9 9 0 2 12 9 0 2
15 7 2 3 9 13 14 4 10 9 13 0 9 13 4 2
11 9 0 13 4 13 2 9 2 9 13 2
25 11 1 2 2 9 8 0 2 13 13 4 9 2 7 3 13 2 9 2 9 2 0 13 2 2
32 11 9 11 9 0 13 4 2 7 2 13 4 9 11 11 13 3 2 9 0 13 13 4 3 11 11 11 9 9 0 13 2
16 11 9 0 0 9 13 9 13 7 9 1 13 13 4 9 2
20 9 13 2 9 3 9 13 4 9 2 7 11 9 1 13 4 3 12 9 2
20 2 9 13 9 2 9 13 4 9 13 13 4 2 3 2 11 9 9 13 2
11 2 9 0 12 13 15 9 0 1 9 2
18 7 2 3 3 13 4 3 13 4 9 0 3 0 13 9 10 13 2
14 11 11 7 11 11 7 2 9 9 1 13 4 13 2
31 9 9 13 2 3 2 9 9 9 0 1 2 9 12 9 9 13 13 13 4 7 9 10 4 11 9 9 12 13 13 2
26 11 11 9 11 11 11 7 9 13 4 2 7 0 9 2 9 0 7 0 9 2 13 4 13 4 2
11 2 9 0 13 9 11 1 9 9 13 2
12 3 7 2 9 11 13 4 11 9 9 13 2
21 11 9 2 9 0 2 12 9 13 4 2 7 9 9 9 13 9 12 13 4 2
12 9 10 1 13 4 11 7 13 13 4 13 2
12 9 10 3 13 4 9 9 9 13 13 4 2
10 11 12 9 1 9 0 13 4 9 2
17 9 7 9 9 7 9 1 9 9 13 9 13 4 10 9 10 2
11 11 11 9 11 9 13 4 9 9 1 2
26 3 12 9 10 1 9 12 13 4 3 11 11 11 9 11 9 0 9 12 9 13 4 9 12 9 2
23 9 9 13 4 2 9 12 2 11 2 7 9 2 7 2 9 12 13 4 2 11 11 2
23 3 2 13 4 9 0 13 4 9 10 9 13 13 14 13 9 7 10 14 4 9 13 2
19 7 2 12 9 9 7 13 4 11 2 7 11 11 11 13 9 13 4 2
9 9 10 9 9 1 13 4 13 2
18 3 1 2 12 9 9 13 4 11 2 7 3 13 4 9 13 9 2
35 9 0 9 9 13 9 13 2 7 11 9 9 1 3 13 13 4 2 7 9 10 14 4 2 3 2 11 11 11 9 13 13 11 11 2
14 9 12 2 9 1 9 13 9 7 9 13 4 9 2
27 3 3 2 9 7 9 9 0 2 9 0 13 4 3 9 2 7 15 0 9 0 10 14 13 9 0 2
12 3 13 4 3 11 11 11 2 11 13 9 2
12 12 9 1 2 11 11 9 3 0 13 4 2
13 3 2 11 0 7 9 7 10 13 13 4 3 2
23 11 11 9 0 11 11 11 11 9 0 13 4 3 2 12 7 12 9 1 3 13 9 2
11 2 12 9 1 13 4 9 14 4 13 2
22 11 2 11 2 11 11 2 11 2 11 11 2 11 2 11 7 11 13 4 9 1 2
14 9 11 9 0 12 9 13 4 2 13 14 4 9 2
11 9 0 13 4 9 0 9 13 9 1 2
26 12 9 13 4 9 11 2 12 9 9 1 2 7 9 12 9 13 4 2 12 9 2 2 12 2 2
28 3 9 13 13 4 9 10 2 11 10 9 1 2 7 10 13 2 3 0 2 0 9 9 0 9 13 4 2
32 13 9 9 10 9 7 9 2 13 9 13 4 13 4 7 9 10 13 9 2 15 9 13 9 13 2 9 9 9 13 13 2
9 12 9 9 9 13 4 11 11 2
14 11 11 13 11 9 2 7 13 13 4 9 11 13 2
13 9 0 9 9 13 9 9 10 9 13 4 9 2
13 3 9 9 1 13 9 12 13 4 2 13 13 2
22 3 2 11 11 11 2 11 11 2 11 11 2 11 11 7 11 11 13 4 13 12 2
17 7 2 9 3 13 2 13 13 4 9 1 9 7 0 9 9 2
18 11 13 9 9 13 4 2 11 14 4 9 0 9 13 12 12 9 2
21 9 9 12 7 13 4 9 9 7 9 13 2 9 9 2 9 9 0 2 9 2
9 11 9 13 4 9 1 9 13 2
18 12 9 14 4 11 13 9 2 7 10 3 9 0 13 4 9 13 2
25 11 9 0 7 2 12 9 13 4 2 11 9 10 9 9 13 13 4 9 0 12 13 13 4 2
14 11 9 13 4 9 11 7 9 9 0 9 9 11 2
13 9 0 9 10 3 13 0 13 4 13 11 1 2
10 11 11 0 13 2 12 13 2 11 2
8 9 1 2 9 13 4 9 2
16 11 9 13 9 0 1 11 9 9 13 9 1 9 13 4 2
22 7 2 12 7 12 9 13 9 13 4 13 0 9 2 7 14 15 10 9 13 9 2
26 11 2 9 13 9 10 13 13 4 2 7 11 11 11 1 11 13 4 9 14 4 3 9 13 2 2
64 9 13 9 0 9 13 4 15 1 13 2 7 3 9 0 13 4 2 9 13 13 4 2 9 7 3 13 2 7 2 3 2 9 10 7 13 4 2 2 13 4 3 11 11 9 2 11 9 2 11 9 2 11 2 2 9 9 13 9 0 10 9 3 2
12 7 2 11 13 4 13 10 13 13 9 9 2
8 9 9 11 9 1 13 4 2
17 9 10 12 9 9 7 12 9 9 13 2 9 3 13 9 1 2
19 11 11 9 0 1 9 1 12 9 12 9 9 0 13 4 9 13 3 2
9 10 9 12 13 11 9 1 9 2
16 11 9 9 9 9 10 13 4 2 9 0 9 0 13 7 2
19 3 13 4 2 11 9 9 13 9 13 4 9 9 7 9 3 9 13 2
17 12 9 2 7 2 3 13 4 2 9 0 13 4 10 10 1 2
20 9 13 2 9 13 9 0 13 14 4 2 3 3 9 10 13 4 9 0 2
14 9 0 13 0 9 13 2 7 11 9 3 13 4 2
19 9 0 13 9 11 9 13 4 3 2 7 9 14 4 3 1 15 13 2
9 0 9 1 3 13 4 9 9 2
13 10 1 2 9 2 9 9 7 9 13 4 2 2
19 11 3 12 9 13 4 9 2 7 11 9 11 13 4 9 3 13 3 2
23 11 9 0 13 4 9 12 13 4 2 7 9 3 9 10 11 9 13 13 13 9 13 2
12 11 9 9 13 12 9 1 13 7 12 9 2
24 3 2 9 10 1 2 9 10 9 13 3 9 10 9 13 2 10 9 9 13 4 2 13 2
10 2 11 0 9 9 13 13 12 9 2
8 13 9 9 0 13 4 11 2
14 14 4 13 10 9 9 12 9 9 13 12 13 4 2
13 3 3 13 2 3 3 13 4 9 1 9 12 2
24 9 9 0 7 9 9 11 7 11 9 9 13 3 13 4 2 3 9 13 9 0 9 13 2
34 14 4 3 13 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 7 2 10 10 2 11 11 9 2
9 2 12 9 13 7 13 13 2 2
19 9 1 9 14 4 13 11 3 9 2 7 9 1 9 9 13 4 9 2
16 9 10 13 4 11 9 0 7 0 9 7 11 9 11 11 2
10 13 2 10 3 2 11 9 13 4 2
11 3 9 11 9 9 13 4 11 11 11 2
9 7 3 7 9 0 1 13 4 2
14 11 9 0 9 13 4 9 2 7 10 1 11 9 2
28 9 9 1 2 2 9 9 10 9 9 13 4 2 7 9 9 1 9 9 3 13 4 2 2 9 12 13 2
14 12 7 12 9 13 4 3 2 9 13 13 8 3 2
21 10 9 2 9 13 11 13 9 13 13 13 4 2 7 3 9 11 9 13 13 2
16 9 13 4 3 10 9 2 3 3 3 9 0 9 13 7 2
16 11 9 9 11 11 11 11 13 9 2 9 0 2 13 4 2
17 11 11 9 13 12 9 13 4 2 7 9 0 13 4 9 0 2
15 11 11 11 13 4 9 2 11 11 7 11 11 0 1 2
28 12 9 12 12 9 13 13 2 7 10 12 2 11 11 2 11 7 11 2 11 9 9 13 4 15 9 0 2
7 10 9 0 9 1 13 2
14 10 0 3 13 4 2 3 2 11 14 4 9 13 2
13 11 13 13 4 15 14 13 2 11 2 10 10 2
16 9 9 13 4 3 11 11 2 9 2 7 0 13 4 9 2
9 9 9 11 11 13 9 13 11 2
14 11 11 13 4 11 11 11 9 13 9 4 13 9 2
15 2 12 9 1 9 13 2 7 9 10 3 4 13 13 2
12 9 0 7 9 1 2 9 7 10 1 13 2
24 11 9 11 11 9 9 9 0 2 11 11 9 9 7 11 9 9 13 4 3 9 12 1 2
10 11 9 11 13 2 11 9 9 12 2
12 11 9 13 9 13 4 9 11 9 13 4 2
11 0 9 11 9 9 13 13 4 11 11 2
7 11 11 9 9 9 13 2
8 3 9 11 9 9 13 4 2
31 11 11 2 9 0 13 9 13 2 7 13 4 9 1 14 4 9 0 1 3 13 2 7 11 12 9 13 13 4 9 2
29 7 2 12 9 9 3 13 4 2 9 0 13 14 7 2 2 7 2 12 9 13 9 14 2 4 13 13 4 2
9 10 13 4 2 7 2 3 9 2
16 7 12 12 9 9 9 10 13 4 9 0 11 11 13 4 2
19 11 11 11 9 11 9 13 4 13 3 12 9 9 9 9 12 13 13 2
34 11 2 9 10 2 2 9 2 13 4 2 9 9 2 9 0 10 2 7 2 9 9 13 4 9 7 11 9 2 9 9 13 13 2
23 11 11 11 9 0 9 9 12 13 7 13 4 13 4 9 2 11 11 9 0 0 9 2
12 9 10 9 9 0 1 9 13 4 9 0 2
20 11 9 9 9 12 1 2 2 9 0 13 11 7 11 1 9 3 13 2 2
27 9 13 13 9 13 7 2 11 11 11 11 9 13 9 12 11 13 4 9 0 11 8 0 13 13 4 2
16 11 7 11 1 2 9 9 2 13 9 13 11 11 9 0 2
10 11 12 1 9 13 4 11 2 11 2
14 12 2 11 11 11 11 13 9 13 4 9 9 13 2
18 3 2 13 9 0 9 0 12 7 9 2 9 7 9 13 4 9 2
30 11 2 11 7 11 3 13 4 3 11 9 0 9 0 9 11 2 11 2 11 7 11 13 4 9 9 13 0 9 2
12 11 9 9 0 13 4 2 9 9 2 13 2
40 10 9 2 11 12 9 0 2 11 9 0 9 12 13 9 2 13 2 7 2 11 10 7 9 10 10 9 2 13 4 2 2 11 9 0 9 13 3 2 2
54 11 11 2 11 2 2 11 11 2 11 2 2 11 11 2 11 7 11 2 2 11 11 2 11 2 7 11 11 11 2 11 2 9 13 9 13 4 2 2 9 10 9 11 9 14 13 9 13 13 2 4 13 3 2
27 11 11 13 0 4 9 2 0 2 13 7 10 13 4 9 14 4 2 0 2 13 4 3 11 11 0 2
20 9 10 13 3 11 12 9 9 1 2 7 9 9 7 12 9 9 13 4 2
15 11 9 9 12 3 13 4 2 9 12 9 4 13 9 2
12 13 13 4 11 9 9 13 2 7 3 3 2
19 9 0 7 13 9 9 13 13 4 9 9 2 12 7 11 13 4 9 2
17 15 9 0 13 7 9 0 14 13 0 9 2 13 13 2 3 2
11 9 13 4 11 11 12 9 9 13 4 2
19 11 12 9 9 1 13 9 13 2 9 0 13 0 9 10 0 9 13 2
16 9 0 10 15 14 4 13 9 2 15 7 14 4 15 13 2
18 11 9 11 13 4 9 11 11 0 12 9 13 2 10 9 13 9 2
22 13 4 2 9 0 2 9 13 4 13 9 13 3 7 3 2 2 10 9 13 0 2
19 9 10 9 13 4 11 11 11 9 7 11 11 9 10 9 13 13 4 2
22 7 2 11 12 12 9 13 4 12 9 9 9 12 2 7 11 9 13 4 2 11 2
22 3 2 11 11 0 9 9 13 13 13 2 10 13 2 3 7 3 2 9 0 9 2
17 9 10 2 13 9 13 11 11 11 9 3 13 4 11 11 9 2
30 0 9 13 9 2 13 4 13 7 9 13 4 11 11 11 7 2 9 13 2 4 13 2 11 2 9 2 13 4 2
22 11 1 9 13 13 4 11 13 3 2 11 11 0 9 9 12 13 7 9 13 4 2
23 9 12 9 1 11 9 7 9 10 9 9 13 9 11 9 3 13 4 11 9 9 13 2
15 11 2 3 7 3 2 9 9 9 12 9 13 9 13 2
12 3 2 11 2 10 3 3 13 4 3 7 2
17 11 9 10 9 13 4 9 0 2 7 3 2 10 13 9 13 2
11 9 14 4 3 13 9 9 13 4 11 2
13 9 9 9 13 7 14 4 9 13 11 9 1 2
14 11 11 13 4 2 2 9 9 1 9 13 4 10 2
18 3 11 9 0 11 13 4 2 7 11 13 4 9 9 13 4 9 2
16 3 2 9 13 9 7 13 13 9 13 4 15 9 13 7 2
28 3 0 13 12 9 10 1 11 2 11 9 0 13 9 2 0 2 3 2 11 9 11 2 9 0 2 13 2
17 3 9 13 4 9 13 4 2 7 9 0 9 9 1 13 4 2
15 7 2 10 9 12 9 13 4 9 2 11 12 9 1 2
16 11 9 13 4 13 9 11 11 2 7 12 9 9 13 4 2
12 2 14 2 7 2 9 3 3 13 4 2 2
25 3 9 0 13 4 11 9 1 13 9 1 7 9 10 3 13 0 9 9 13 4 2 0 3 2
20 13 10 10 7 2 13 0 9 7 2 9 0 11 14 4 0 1 13 3 2
11 11 9 13 2 10 9 12 2 13 13 2
13 2 9 1 13 4 9 12 10 13 13 4 2 2
13 11 11 3 12 9 13 4 2 7 9 10 13 2
11 12 9 9 0 13 4 9 13 4 3 2
11 10 3 13 7 9 13 4 9 12 1 2
12 11 11 11 12 13 4 2 11 2 11 2 2
17 11 9 12 11 9 13 4 2 9 1 9 0 11 11 13 4 2
9 11 13 4 9 9 9 1 13 2
16 9 0 12 1 9 12 13 2 9 10 9 1 9 13 4 2
18 9 2 9 0 0 13 4 7 14 2 12 11 1 2 9 7 9 2
15 2 14 13 10 13 4 2 7 9 13 4 13 13 4 2
9 3 2 11 11 0 13 4 9 2
10 0 12 9 9 12 13 4 11 11 2
15 10 9 2 3 9 2 11 9 10 13 2 3 13 4 2
23 7 2 11 7 11 12 12 2 15 9 0 13 0 13 9 13 4 7 11 9 13 4 2
14 9 2 9 7 9 9 13 4 9 9 13 9 13 2
11 11 11 9 13 2 7 13 3 9 3 2
15 0 9 13 9 1 2 7 9 0 13 4 9 10 9 2
20 11 2 7 2 0 9 9 13 4 9 12 2 10 12 2 9 1 13 4 2
13 13 14 13 2 10 9 3 9 13 4 13 4 2
14 10 9 13 9 13 4 9 10 1 2 3 13 4 2
9 12 9 1 14 4 13 9 13 2
12 13 13 9 0 2 7 3 13 10 4 13 2
18 7 0 9 13 3 7 2 11 3 13 9 10 13 2 9 12 12 2
20 11 11 11 2 11 2 11 2 11 2 0 9 2 7 11 11 13 4 9 2
18 7 10 10 4 13 13 3 11 2 3 2 9 2 13 4 9 10 2
19 9 0 13 4 3 9 2 11 11 2 3 9 11 3 9 9 9 9 2
13 11 11 11 9 3 9 11 13 9 9 13 4 2
28 9 10 2 10 9 12 1 13 4 2 15 2 12 9 8 9 4 13 2 7 9 13 3 2 13 13 4 2
16 11 11 7 11 11 13 10 3 2 7 9 9 13 11 9 2
13 11 11 9 0 11 9 11 11 13 4 3 11 2
35 10 9 0 13 4 15 7 15 9 2 7 2 12 1 9 3 13 7 2 9 9 10 13 4 9 13 14 4 10 2 10 13 9 13 2
13 9 10 9 1 13 13 2 7 14 13 9 9 2
7 0 0 13 2 9 1 2
13 9 0 9 4 13 9 0 9 14 4 13 2 2
17 7 2 11 9 11 11 3 13 4 3 10 9 13 9 7 9 2
9 9 4 15 13 9 9 3 13 2
9 10 9 2 9 13 4 9 9 2
10 11 9 9 3 13 4 2 12 9 2
22 3 0 13 2 9 10 2 9 12 9 9 1 13 12 7 9 9 9 9 13 4 2
17 11 7 11 9 12 13 4 9 2 7 9 13 4 12 9 13 2
24 10 9 2 9 0 1 13 2 9 9 7 9 9 2 13 2 7 3 13 10 14 4 13 2
15 13 9 13 4 11 11 9 10 9 13 4 11 9 13 2
24 11 7 13 3 13 2 7 10 1 11 10 9 13 0 13 4 2 12 7 11 13 4 9 2
19 11 13 2 11 9 3 13 4 13 7 9 10 13 4 9 13 9 9 2
10 7 2 10 9 9 1 13 4 9 2
21 13 4 9 8 9 12 10 13 4 11 9 0 9 13 2 11 14 4 13 3 2
12 9 1 9 9 2 9 13 4 3 11 9 2
16 7 12 9 12 9 13 9 2 11 2 3 9 0 13 4 2
13 11 9 0 0 0 14 13 3 10 9 0 13 2
14 9 0 3 13 11 9 13 7 11 9 10 13 7 2
17 11 11 9 3 13 4 9 9 13 4 7 9 9 1 13 4 2
18 9 1 2 7 2 9 13 9 0 12 13 4 2 9 13 13 4 2
5 9 1 9 13 2
21 11 13 4 14 13 7 2 9 13 4 9 13 0 9 14 13 13 4 11 11 2
21 11 11 2 7 2 9 13 4 2 7 2 9 2 9 9 12 14 4 9 13 2
13 9 9 9 7 11 9 13 3 2 9 9 13 2
9 11 9 9 0 12 9 12 13 2
14 11 9 10 13 4 12 9 7 3 13 4 9 13 2
17 11 13 9 0 13 13 3 11 7 11 9 13 9 13 13 4 2
12 10 14 4 3 13 9 1 9 13 9 10 2
24 7 2 13 4 7 2 11 14 4 9 13 2 3 3 9 11 11 9 13 4 9 13 4 2
11 7 2 14 4 9 13 11 13 9 10 2
12 11 11 11 2 11 11 12 13 4 9 11 2
32 9 9 10 2 13 9 1 9 13 3 2 13 9 13 4 2 12 9 9 7 12 9 9 13 9 9 12 0 13 9 1 2
18 9 0 9 13 3 0 13 2 9 10 9 13 9 13 13 12 12 2
19 11 11 11 9 14 4 11 13 2 9 10 9 0 10 13 9 10 13 2
18 10 13 11 9 9 11 3 13 4 3 9 7 3 13 4 9 9 2
9 15 9 9 1 9 0 12 13 2
24 9 0 10 11 9 9 1 0 9 13 14 7 2 10 9 13 4 0 0 9 7 13 4 2
23 11 9 9 9 1 13 9 9 13 13 9 0 13 4 2 9 10 11 12 9 0 1 2
20 2 9 1 9 13 4 10 9 2 2 2 9 13 2 13 4 9 7 9 2
17 11 9 11 1 13 14 4 13 13 4 11 9 9 11 11 11 2
18 11 7 11 11 11 13 4 9 2 9 0 2 13 4 11 9 9 2
8 2 15 9 13 9 3 13 2
16 0 9 13 13 4 2 9 13 4 13 9 9 11 9 13 2
17 9 12 9 9 1 9 0 13 4 7 9 3 13 13 4 9 2
10 11 2 10 1 2 9 13 9 13 2
10 9 0 1 0 9 13 4 9 0 2
13 7 11 11 11 2 7 13 4 0 1 13 4 2
8 2 9 9 1 13 4 9 2
15 11 11 9 12 9 13 11 11 13 4 11 7 11 1 2
13 11 13 9 11 9 9 0 13 4 12 9 3 2
14 7 2 9 13 4 9 0 12 13 4 12 9 1 2
13 11 9 10 13 4 13 9 7 9 0 13 13 2
14 11 9 9 1 2 11 13 4 2 11 1 2 9 2
14 9 9 10 1 2 9 7 9 0 9 13 4 11 2
24 9 11 13 2 7 11 9 0 13 4 9 11 9 9 13 4 2 7 14 11 2 13 3 2
20 9 13 4 9 1 9 0 13 4 11 11 11 9 9 0 9 7 11 11 2
7 2 10 0 9 13 4 2
8 9 0 9 13 9 13 9 2
7 9 13 7 0 13 4 2
15 3 7 9 1 10 9 13 4 9 9 11 11 13 3 2
25 3 2 11 2 11 7 11 1 9 0 9 10 13 4 11 9 2 3 7 3 9 9 0 13 2
16 12 9 9 9 0 13 3 11 1 13 4 12 9 9 13 2
22 11 9 13 13 9 10 10 13 4 2 7 3 11 1 13 9 9 10 3 13 4 2
12 12 9 9 9 9 13 4 11 9 9 13 2
21 3 2 9 9 1 9 13 9 9 13 4 9 10 9 7 3 9 0 13 4 2
14 3 2 7 2 12 9 7 10 9 13 9 13 4 2
23 15 3 13 2 7 2 9 9 13 9 9 1 3 13 3 2 12 9 13 4 9 9 2
28 15 9 0 12 9 13 13 3 2 7 2 10 2 15 9 0 7 0 13 13 4 2 2 13 4 9 0 2
9 0 1 13 4 9 1 10 13 2
15 11 9 11 11 11 9 9 9 9 3 9 12 13 4 2
8 9 0 1 11 11 13 4 2
15 10 10 2 3 3 2 15 9 0 13 12 9 13 4 2
18 12 9 9 13 3 2 11 11 9 9 9 9 12 13 4 11 9 2
18 9 9 0 9 13 4 2 9 7 9 9 7 9 1 9 10 1 2
20 11 11 9 1 13 4 9 13 2 10 13 4 13 2 9 2 9 7 9 2
7 11 3 9 13 11 9 2
24 12 9 2 11 2 9 1 2 3 13 4 11 9 2 7 11 9 13 9 13 13 4 3 2
12 3 13 9 13 9 0 12 1 13 4 10 2
14 2 9 7 9 1 13 9 13 9 0 13 9 9 2
18 10 13 7 2 11 11 0 7 11 11 14 4 11 0 9 9 13 2
21 2 11 11 13 13 4 2 9 13 4 2 7 9 13 9 0 13 13 4 2 2
17 11 9 0 9 13 4 11 11 9 11 9 9 11 13 9 13 2
25 10 13 7 2 0 11 9 1 2 13 10 11 12 11 9 2 9 0 0 2 9 9 9 1 2
20 7 10 3 9 13 4 9 9 13 13 2 9 9 10 3 13 9 14 13 2
19 9 9 13 4 9 11 13 4 2 11 9 2 7 11 3 13 9 13 2
12 13 12 9 1 9 0 12 13 4 13 11 2
19 9 7 9 9 1 2 9 7 9 1 13 4 11 9 7 10 9 9 2
8 2 9 13 13 9 13 2 2
11 13 13 9 9 12 13 13 9 12 10 2
14 13 3 2 9 10 13 13 13 11 11 13 9 9 2
11 9 1 9 9 13 13 4 13 11 9 2
17 3 9 0 13 4 9 0 12 1 2 3 9 0 12 1 13 2
12 12 9 0 1 2 12 9 13 4 9 9 2
22 3 1 9 0 2 13 12 9 2 9 12 3 0 2 13 4 11 9 9 9 13 2
10 9 13 2 9 13 7 13 13 4 2
5 9 3 13 4 2
11 9 9 3 0 13 2 7 9 9 14 2
8 0 9 9 13 4 12 9 2
18 13 13 7 9 10 2 9 9 9 9 7 9 9 9 13 13 4 2
19 7 2 10 9 3 0 13 4 2 3 3 11 0 9 7 11 0 9 2
10 12 9 9 0 13 4 12 9 1 2
10 13 7 2 15 10 9 13 15 13 2
17 9 11 7 9 11 9 0 9 9 13 4 9 13 9 3 13 2
17 9 2 11 9 11 11 13 4 9 0 7 10 12 9 9 13 2
19 9 10 2 3 3 9 12 13 9 13 12 9 2 3 11 13 9 13 2
10 11 9 9 9 9 12 13 13 4 2
6 11 9 13 10 13 2
8 9 1 14 13 3 9 0 2
19 3 2 11 11 9 13 7 12 12 9 2 12 12 9 2 13 4 11 2
4 3 0 13 2
19 9 9 9 13 3 2 3 7 11 11 2 11 11 2 0 13 4 0 2
11 11 3 13 4 11 11 2 11 9 0 2
10 11 1 9 10 11 9 1 13 4 2
18 9 12 9 13 4 3 11 9 2 7 9 9 9 11 11 13 4 2
17 9 9 1 7 2 9 11 9 11 13 4 11 9 9 13 4 2
10 12 9 1 2 7 2 3 13 4 2
20 11 9 13 2 2 9 3 13 2 13 13 9 11 2 3 9 6 12 13 2
9 7 14 4 9 13 9 10 1 2
26 7 2 11 10 9 13 4 7 11 11 2 11 11 2 7 11 2 11 2 9 13 4 2 10 10 2
22 11 11 11 9 9 13 13 4 11 13 9 2 7 3 13 9 12 13 4 13 4 2
16 11 12 9 1 13 4 7 3 7 0 9 9 13 4 13 2
9 3 9 13 4 9 13 4 9 2
12 10 13 4 11 9 11 11 13 9 13 9 2
11 11 11 11 1 13 4 3 2 12 2 2
7 9 13 9 7 9 0 2
9 11 9 11 11 13 4 12 9 2
11 11 9 12 9 9 0 13 4 9 0 2
9 9 10 13 4 3 9 9 9 2
5 2 13 2 13 2
16 11 3 13 4 2 7 11 7 14 2 3 10 13 4 7 2
11 9 10 13 13 13 4 3 11 9 9 2
6 11 9 9 13 13 2
7 15 9 10 0 13 9 2
13 9 0 7 9 9 9 11 11 13 13 4 9 2
24 9 11 11 11 9 9 13 4 9 2 9 11 11 11 9 9 9 7 9 11 11 11 9 2
13 2 14 2 9 14 13 2 9 9 1 2 7 2
15 11 9 9 13 4 11 9 13 7 0 9 13 4 13 2
27 11 9 13 4 9 13 4 9 10 13 12 9 13 9 13 9 12 8 3 2 9 10 13 4 9 9 2
22 9 11 3 13 2 9 2 13 4 13 4 2 7 9 10 9 0 1 13 13 4 2
7 11 9 12 9 13 4 2
17 11 1 2 11 9 13 9 14 4 13 2 10 10 2 0 9 2
9 12 11 11 13 4 2 12 9 2
10 11 11 9 13 4 9 0 9 9 2
21 9 14 4 13 11 0 2 9 2 13 3 13 13 11 11 2 11 2 9 9 2
16 3 15 14 4 13 10 9 2 7 10 9 13 11 9 13 2
9 3 9 2 9 9 9 13 4 2
8 11 11 9 9 9 13 4 2
18 9 1 13 4 11 11 11 0 0 9 11 11 2 12 9 13 4 2
9 9 12 9 9 1 13 4 9 2
24 3 9 9 3 13 9 13 9 13 2 3 7 11 11 11 9 9 9 9 13 13 4 11 2
33 11 9 11 9 12 9 2 11 11 7 11 11 7 9 9 12 9 2 11 11 2 11 11 2 11 11 7 11 11 13 4 9 2
9 13 9 9 0 13 7 3 13 2
11 11 11 3 13 4 10 9 14 13 9 2
18 11 11 11 9 9 9 13 4 11 11 2 2 9 0 12 13 2 2
8 13 7 0 13 4 9 1 2
16 9 7 9 13 2 11 13 4 3 9 9 1 2 9 13 2
15 9 1 13 4 2 14 9 9 14 9 2 7 0 1 2
13 0 15 13 4 3 9 2 3 9 13 13 4 2
6 11 9 13 2 13 2
8 11 11 9 0 13 4 11 2
23 9 9 13 7 13 13 4 2 0 9 13 4 9 9 12 13 7 10 13 4 9 13 2
15 9 13 4 7 9 1 9 9 0 13 13 4 9 9 2
21 11 2 11 2 11 2 13 10 7 0 9 10 13 4 11 2 12 9 2 3 2
15 11 9 14 7 2 11 9 0 7 13 4 9 7 9 2
21 9 9 13 4 10 9 1 9 12 9 9 9 9 13 2 9 13 9 9 2 2
12 9 9 10 9 1 9 0 13 4 9 9 2
7 9 0 13 9 12 1 2
13 9 9 11 11 13 4 3 2 9 12 9 13 2
13 10 9 2 9 13 7 2 9 10 10 13 4 2
19 3 2 11 9 9 14 13 9 3 13 9 2 7 9 13 9 13 4 2
7 9 13 10 13 4 9 2
14 9 9 9 2 7 2 12 9 9 7 14 13 9 2
7 9 1 14 4 9 13 2
20 14 4 3 3 3 13 2 7 9 13 0 13 4 3 1 13 7 10 13 2
32 13 11 2 11 2 11 7 11 2 10 1 2 3 3 9 0 13 2 7 10 1 2 13 10 9 1 10 9 9 13 4 2
13 10 0 9 12 3 13 13 4 13 11 7 11 2
28 11 11 11 12 9 7 9 9 9 9 9 13 4 2 10 9 9 12 13 4 9 11 9 11 11 9 13 2
19 9 10 13 13 13 4 9 9 11 9 2 9 12 1 10 9 13 3 2
24 11 2 11 2 2 11 2 11 2 2 11 2 11 11 2 7 11 2 11 2 13 4 11 2
9 11 9 14 13 10 1 9 0 2
21 2 9 11 2 9 9 13 9 13 2 7 9 13 9 2 10 13 15 9 0 2
18 12 9 1 9 13 4 10 9 2 12 12 11 12 9 0 13 3 2
18 11 11 9 0 13 4 11 2 7 2 11 1 2 9 1 13 4 2
22 11 9 0 13 4 11 1 9 13 2 12 7 11 7 11 2 3 0 9 13 4 2
17 11 11 12 9 9 13 3 2 11 11 13 4 13 4 3 9 2
22 9 0 13 9 13 9 13 4 9 12 9 10 1 9 13 9 0 12 13 13 4 2
11 9 13 4 11 11 13 2 3 13 7 2
11 11 11 9 0 13 4 9 11 9 9 2
27 3 0 4 13 13 11 11 11 11 2 7 12 9 13 4 9 0 2 11 11 11 0 12 7 12 13 2
11 7 2 9 9 0 9 1 13 13 4 2
10 11 11 11 11 9 13 4 9 0 2
10 0 9 3 13 4 10 9 9 1 2
17 9 0 13 2 3 0 2 9 9 10 1 13 9 9 11 1 2
15 9 1 13 4 9 12 7 12 13 9 9 1 13 4 2
23 9 0 9 11 13 12 9 7 10 12 9 13 9 3 9 13 4 13 4 3 9 0 2
19 11 13 9 2 12 7 12 9 2 0 13 4 11 2 12 7 12 2 2
16 9 9 9 7 9 13 4 11 9 9 7 9 3 7 3 2
10 11 11 7 3 3 13 4 9 10 2
19 11 11 7 11 9 13 9 1 2 2 9 7 9 9 0 13 4 2 2
24 11 2 7 2 11 9 0 11 11 13 9 13 9 9 13 2 7 15 13 9 13 0 13 2
20 11 9 1 2 2 11 10 13 9 13 11 9 2 7 14 4 15 13 2 2
9 0 7 0 2 9 13 11 0 2
11 3 2 9 9 13 0 10 9 10 1 2
11 12 9 9 13 4 9 7 9 11 9 2
12 9 3 2 11 11 11 0 1 13 4 11 2
24 12 9 11 11 11 9 1 13 4 11 7 0 9 1 13 4 12 9 2 12 7 12 2 2
25 9 9 1 9 13 13 13 4 13 4 11 2 7 9 10 11 11 11 9 13 13 9 13 4 2
13 11 9 13 4 11 2 2 9 13 2 9 1 2
14 2 15 9 3 13 4 2 9 7 9 12 7 2 2
12 15 3 1 13 4 2 9 0 13 4 7 2
19 11 13 4 2 11 12 9 13 4 9 11 2 9 10 13 9 13 9 2
24 9 12 9 12 1 13 4 2 7 12 9 13 2 12 9 9 13 4 2 7 13 7 13 2
25 9 9 2 3 2 14 4 13 9 12 13 3 13 9 13 4 11 9 1 13 13 9 9 12 2
12 11 13 0 3 7 13 13 4 11 9 9 2
18 3 11 13 13 4 11 2 7 11 1 13 2 7 15 9 13 9 2
10 13 7 9 9 13 9 12 13 4 2
24 9 9 1 10 9 13 4 2 9 0 12 7 2 7 12 9 11 0 7 10 10 9 7 2
21 7 2 9 1 13 9 9 13 9 3 13 13 7 13 4 9 13 4 10 9 2
18 11 7 11 2 9 7 9 2 9 4 13 9 15 13 9 13 13 2
13 11 13 11 2 11 7 11 9 13 4 10 10 2
19 9 12 9 1 2 9 9 7 9 9 9 13 4 13 9 12 8 3 2
13 11 11 11 9 2 7 2 0 9 9 13 4 2
14 9 13 3 2 3 13 0 13 9 11 9 9 3 2
13 11 9 2 9 10 2 11 0 7 0 8 13 2
27 11 11 11 9 9 0 13 4 9 11 12 9 2 12 9 7 12 9 2 7 10 9 12 13 4 11 2
14 11 11 9 13 4 2 9 15 13 4 13 13 4 2
19 9 10 0 9 10 1 13 4 7 9 7 9 13 4 9 9 0 1 2
21 0 9 9 9 12 10 13 4 2 7 11 3 9 0 13 4 7 9 13 4 2
19 11 11 4 9 2 11 13 13 2 7 3 13 13 4 2 11 13 4 2
26 11 9 2 3 2 0 11 9 3 13 11 9 9 0 13 4 13 7 9 9 7 0 13 13 4 2
10 13 8 11 0 9 13 3 9 11 2
27 3 9 2 0 13 2 3 13 13 4 9 9 9 13 4 13 4 2 12 9 9 13 9 3 7 13 2
8 10 13 9 3 7 15 9 2
19 9 0 9 15 1 13 4 2 7 9 2 7 2 9 0 0 13 4 2
15 9 3 3 13 4 11 2 11 13 12 9 9 13 9 2
16 3 1 9 0 9 13 4 9 2 7 9 13 4 10 9 2
9 9 9 7 9 13 13 4 11 2
21 12 9 9 13 9 13 4 9 7 13 4 9 13 2 9 12 9 13 4 13 2
22 14 2 0 13 2 15 10 9 12 2 9 12 13 2 7 7 3 15 9 7 13 2
25 11 11 2 11 2 9 9 1 9 13 13 4 3 11 9 9 1 2 13 4 13 0 9 2 2
24 3 11 9 7 11 11 13 4 2 7 3 9 2 7 3 13 4 10 9 13 9 0 2 2
9 9 1 13 7 11 9 13 4 2
25 11 13 9 1 13 4 11 11 9 13 9 2 9 9 2 7 9 9 0 13 9 9 13 4 2
15 12 9 2 12 9 13 4 9 9 1 2 9 9 9 2
11 3 2 9 11 9 13 4 12 9 13 2
27 9 13 13 4 11 11 13 7 10 13 2 11 8 11 7 11 11 0 9 13 9 12 13 4 13 4 2
9 11 9 3 13 4 9 13 9 2
10 7 2 3 7 2 13 13 4 9 2
10 11 9 12 9 13 4 3 11 9 2
17 7 2 9 13 9 6 12 13 2 9 9 7 13 4 13 4 2
21 11 11 11 9 13 4 9 2 9 9 2 13 4 2 12 9 9 14 13 13 2
12 11 9 9 13 3 13 13 4 12 9 0 2
14 9 13 2 0 13 13 4 2 9 1 9 13 4 2
19 3 11 14 13 7 2 3 3 13 7 2 11 3 13 9 13 10 9 2
15 9 13 3 12 9 0 7 9 0 9 2 9 13 4 2
21 2 11 11 12 9 9 0 9 12 13 13 4 2 7 11 9 13 4 13 2 2
23 9 10 9 13 13 11 13 2 7 3 11 13 13 4 0 9 3 11 11 13 9 13 2
21 9 12 9 9 13 4 3 9 13 2 12 9 1 2 7 12 9 13 4 9 2
22 9 9 0 1 13 7 9 9 9 3 0 13 4 2 9 9 2 9 2 0 13 2
18 12 12 13 13 4 11 9 11 11 0 2 10 0 9 2 11 1 2
9 10 7 3 13 4 2 15 1 2
23 9 11 13 4 2 10 11 11 9 13 4 7 9 3 2 9 13 4 9 11 9 13 2
7 10 1 11 11 13 4 2
12 10 1 2 7 2 11 9 13 4 11 9 2
14 11 11 9 13 4 9 9 3 13 4 9 12 9 2
12 9 13 10 7 13 11 7 10 9 1 9 2
13 11 0 9 13 2 3 13 4 11 12 11 9 2
16 12 9 12 9 9 12 9 0 7 9 0 13 9 13 13 2
11 9 13 9 0 13 13 4 2 11 1 2
10 9 13 4 0 9 1 13 9 13 2
14 10 9 9 10 1 13 4 2 0 9 9 1 2 2
14 9 10 2 3 7 2 14 4 9 9 9 9 13 2
27 10 13 4 11 2 11 7 11 9 9 2 11 2 7 9 10 9 10 9 9 0 1 9 13 13 4 2
17 11 9 1 2 10 12 13 4 11 2 11 2 11 12 9 9 2
15 12 12 9 9 2 9 1 9 9 2 13 13 4 9 2
15 2 9 0 9 0 13 4 13 4 9 11 15 12 9 2
22 11 2 9 13 13 7 3 3 13 4 2 7 11 2 7 2 9 1 9 13 4 2
12 12 9 9 0 13 7 11 3 0 13 4 2
17 11 11 11 9 13 11 9 0 0 9 0 3 13 13 4 9 2
30 12 9 2 11 11 11 11 9 0 0 9 13 4 9 1 2 7 2 10 9 2 13 4 12 9 13 4 13 9 2
31 9 9 9 0 13 4 2 14 13 10 9 12 9 9 2 2 9 0 13 7 2 9 1 9 10 13 13 4 9 13 2
21 13 4 2 14 13 3 0 2 7 3 13 2 13 7 9 9 9 10 13 9 2
11 11 9 1 2 13 0 13 13 4 9 2
26 0 9 0 9 0 13 2 0 13 9 7 9 1 13 4 9 11 11 9 2 7 9 14 4 13 2
10 11 14 4 11 9 13 2 9 9 2
26 12 9 9 0 13 9 2 11 11 7 11 11 13 4 3 7 9 2 9 11 1 13 9 13 12 2
18 11 7 11 9 1 2 11 11 7 11 13 9 13 4 12 9 12 2
21 7 2 11 7 0 9 1 9 3 13 4 2 11 10 9 13 4 3 7 3 2
18 9 9 3 13 13 4 13 4 9 2 7 3 13 4 3 9 10 2
22 3 3 2 3 2 11 3 13 9 7 9 13 4 7 2 9 13 12 9 9 0 2
21 11 9 9 14 4 9 13 13 12 9 2 11 9 9 10 13 4 3 9 13 2
15 9 1 2 7 2 13 4 2 7 0 9 13 4 9 2
10 9 9 14 4 9 13 9 1 13 2
13 11 9 3 13 13 4 2 7 10 3 13 13 2
24 9 12 9 12 7 12 9 9 9 0 13 4 2 3 7 2 9 7 9 0 0 13 9 2
20 15 8 9 0 13 4 11 11 9 9 2 10 9 9 9 13 4 11 1 2
7 9 12 9 13 13 4 2
21 11 9 0 9 0 3 12 9 13 4 12 9 13 4 11 9 9 0 13 11 2
11 11 11 2 12 2 13 4 12 10 10 2
18 11 9 12 13 4 2 11 2 7 9 13 2 11 9 0 3 13 2
13 9 11 11 9 9 13 4 9 13 4 11 11 2
15 9 10 13 4 3 0 7 11 9 9 13 4 9 0 2
16 11 9 9 9 2 10 3 2 0 13 4 2 9 7 9 2
11 11 9 10 9 10 1 13 11 3 13 2
6 9 9 12 13 4 2
17 9 10 9 14 13 9 9 12 1 2 9 10 13 4 11 9 2
14 10 2 9 10 1 2 9 13 4 11 13 9 1 2
21 3 12 9 2 12 9 9 1 2 12 9 1 2 13 4 13 3 9 11 11 2
16 9 12 9 1 9 7 10 1 13 4 9 9 3 0 13 2
11 7 9 15 9 13 13 4 7 3 13 2
20 11 13 2 12 9 1 2 12 9 13 4 13 4 2 3 3 12 9 13 2
18 0 0 9 13 9 10 13 9 13 11 9 2 10 9 11 13 13 2
13 7 2 0 11 9 13 4 10 9 9 13 4 2
13 12 9 0 10 9 13 13 4 13 4 11 9 2
9 11 11 0 7 9 10 13 4 2
6 9 13 13 4 9 2
18 9 1 2 11 9 13 4 2 7 10 9 13 4 14 4 3 13 2
20 9 9 3 2 11 9 10 13 4 9 0 9 12 2 11 15 9 13 9 2
13 2 9 9 10 13 4 7 3 9 7 14 2 2
14 9 1 13 7 2 0 11 0 13 4 3 9 11 2
20 11 9 9 0 9 10 13 4 2 7 13 13 4 9 9 0 14 13 9 2
11 7 3 11 2 13 3 2 13 4 13 2
16 3 12 12 9 1 13 13 4 0 2 7 3 13 9 10 2
13 9 3 13 2 11 11 9 13 4 9 9 1 2
17 11 11 2 7 2 9 9 9 13 4 2 7 0 9 9 9 2
8 3 9 13 4 12 9 11 2
6 0 3 1 13 4 2
19 11 3 13 13 4 9 9 7 14 11 14 11 14 4 13 13 4 11 2
20 9 11 9 10 13 4 3 2 11 9 9 2 7 3 13 4 9 1 9 2
20 11 9 9 0 13 4 12 9 11 11 11 9 9 7 11 11 9 9 1 2
14 13 13 10 0 13 2 9 9 13 9 9 13 4 2
11 3 9 0 13 13 9 13 4 11 1 2
10 9 0 11 11 13 13 3 13 4 2
8 2 13 2 13 4 9 0 2
17 3 2 10 9 13 13 4 15 13 7 2 3 7 2 9 13 2
14 9 1 9 13 4 11 9 3 13 4 12 9 9 2
9 2 9 13 9 13 4 13 2 2
12 9 1 11 9 11 9 13 4 3 13 3 2
8 11 11 11 9 1 13 4 2
13 11 11 13 4 12 9 13 4 11 11 13 9 2
45 9 9 9 9 1 12 12 2 9 9 10 9 13 4 9 9 13 7 2 11 9 11 11 2 11 2 13 4 13 9 12 9 2 0 9 2 9 13 4 9 0 13 13 4 2
14 9 10 14 13 9 0 0 3 0 7 9 1 4 2
23 3 7 11 11 13 4 9 11 13 4 9 2 9 9 11 13 7 11 9 13 4 2 2
8 12 12 1 0 9 13 4 2
7 15 13 4 9 7 3 2
24 9 3 7 3 13 4 3 11 9 2 7 12 9 3 9 13 4 9 0 13 7 3 13 2
11 15 2 11 0 12 7 12 9 13 4 2
22 10 13 7 2 9 13 2 3 13 4 11 9 9 0 13 4 11 9 9 2 12 2
13 11 11 12 9 13 7 11 0 13 2 11 9 2
31 11 9 9 11 7 9 9 1 13 4 9 9 9 13 9 9 13 13 4 3 2 11 2 11 7 9 0 13 9 13 2
24 11 0 9 9 11 11 13 4 11 9 2 7 13 13 4 11 11 0 2 11 12 9 13 2
10 10 2 11 9 3 13 4 13 4 2
17 2 3 3 2 9 10 9 12 13 2 9 0 9 13 4 2 2
11 9 1 2 3 13 9 0 0 0 0 2
27 12 3 2 11 2 9 9 0 13 9 2 9 0 13 7 12 9 13 4 2 11 1 7 11 12 9 2
24 9 0 3 3 1 14 4 13 3 2 7 9 13 0 13 4 2 0 13 7 0 13 4 2
13 11 9 0 9 11 0 13 13 4 3 11 9 2
21 7 9 7 9 13 10 9 13 2 9 10 9 0 12 13 7 13 9 13 13 2
17 13 9 12 13 9 13 2 13 12 9 12 13 9 13 4 9 2
20 3 2 7 2 9 9 1 9 7 9 9 13 4 2 9 13 9 13 4 2
13 9 9 13 2 7 3 2 13 13 2 0 13 2
15 10 13 13 4 11 9 2 13 9 10 9 13 9 13 2
9 9 13 2 12 7 9 13 4 2
22 11 11 11 11 0 13 4 3 12 1 11 7 11 11 9 9 13 4 9 9 0 2
14 11 1 9 7 13 4 14 13 9 10 0 9 13 2
10 0 12 1 11 12 13 4 13 4 2
10 11 9 13 4 11 9 13 13 9 2
18 7 9 2 11 9 2 15 13 4 3 2 9 0 12 1 13 4 2
16 9 9 0 12 2 9 0 2 3 9 13 9 13 4 3 2
13 2 11 9 14 4 3 13 9 13 13 4 13 2
13 7 2 11 11 9 12 9 7 12 9 13 4 2
30 9 13 9 3 9 0 13 4 7 3 9 9 9 13 10 2 10 9 4 9 2 3 2 3 13 4 9 13 4 2
10 3 13 4 3 12 11 9 13 12 2
21 12 9 3 13 4 9 13 12 9 1 2 7 9 9 13 2 11 11 0 1 2
14 11 2 11 9 13 9 1 13 4 9 3 9 10 2
14 10 11 2 9 13 2 7 2 9 0 0 13 4 2
10 11 7 9 13 9 13 9 13 4 2
8 3 13 4 3 9 12 1 2
10 11 11 10 12 9 9 13 4 9 2
9 9 9 13 11 11 11 11 9 2
15 11 10 7 2 9 13 4 9 13 9 9 10 13 4 2
18 11 0 9 9 3 9 11 13 9 13 4 2 9 13 9 0 13 2
18 7 2 9 9 12 1 2 13 13 3 2 9 7 9 2 9 10 2
10 11 9 1 0 9 9 0 13 4 2
28 2 11 9 0 0 13 4 12 9 9 9 0 9 13 2 9 9 0 10 1 2 10 9 7 9 9 9 2
22 10 13 2 7 2 11 9 2 10 9 13 2 9 13 4 12 7 2 3 2 0 2
7 9 1 11 13 9 13 2
14 9 12 9 13 4 9 1 11 13 4 12 9 0 2
14 11 9 11 14 4 3 9 1 3 9 1 9 13 2
24 8 14 3 2 9 13 4 9 2 9 11 13 9 13 2 7 10 13 2 3 13 9 13 2
15 11 11 9 13 4 11 9 0 2 0 9 11 9 13 2
9 7 0 9 4 13 13 2 7 2
11 10 15 9 13 4 13 9 11 13 4 2
10 2 3 13 4 2 10 9 8 0 2
11 9 1 9 12 1 13 0 7 13 4 2
16 13 13 4 9 12 13 10 1 2 7 9 13 10 9 9 2
19 9 13 4 9 11 9 11 9 13 2 7 2 7 2 9 11 9 9 2
16 11 2 11 7 11 2 11 11 9 9 0 7 13 4 3 2
28 9 3 13 4 13 9 13 4 2 7 3 13 2 7 2 3 7 3 7 13 14 4 2 14 4 15 13 2
15 9 0 13 4 11 11 3 9 9 2 9 9 9 13 2
11 2 11 1 13 9 13 9 13 11 13 2
14 11 9 0 13 4 2 2 9 9 1 0 2 13 2
17 11 11 3 13 9 13 9 13 7 13 9 13 2 0 9 13 2
26 11 11 11 9 9 12 3 13 9 1 2 11 8 11 9 9 9 9 13 4 9 12 7 9 12 2
12 9 7 9 13 4 9 9 0 9 13 4 2
20 11 1 13 0 9 13 4 11 2 9 9 9 7 11 9 9 9 13 4 2
23 13 12 9 11 9 0 13 4 11 11 9 9 2 7 3 1 9 10 9 12 13 4 2
23 11 11 11 2 11 11 9 7 11 11 13 4 9 13 4 0 2 12 7 12 9 2 2
14 9 9 1 2 9 13 13 4 11 11 2 12 9 2
13 7 2 11 9 13 9 0 9 0 13 13 4 2
14 9 0 9 1 12 9 13 4 3 11 2 11 9 2
22 9 11 13 13 11 13 13 4 9 2 7 10 2 3 13 0 9 12 2 11 3 2
17 0 10 9 0 9 9 13 4 2 2 9 9 2 13 4 9 2
8 7 14 13 9 9 13 4 2
11 9 3 13 7 15 0 13 4 15 9 2
21 11 11 11 9 0 9 9 10 1 13 9 0 2 0 2 13 4 0 9 9 2
21 10 9 2 9 9 13 3 7 3 9 1 9 0 7 0 13 3 13 9 13 2
10 11 9 10 9 9 9 13 11 1 2
10 11 9 9 1 9 9 13 9 13 2
18 11 11 9 0 12 9 13 4 14 4 9 13 0 13 4 12 9 2
37 9 0 13 9 9 2 9 2 9 0 12 9 2 12 9 9 2 12 9 2 12 9 7 12 9 0 7 11 9 12 9 7 0 12 13 4 2
13 9 13 4 2 11 1 9 9 13 4 9 13 2
11 9 12 13 4 13 4 11 9 13 0 2
28 11 11 11 13 4 9 13 4 7 9 12 13 4 12 9 2 3 3 9 9 13 4 2 9 2 9 9 2
17 2 11 9 3 13 4 9 2 7 3 9 10 13 9 13 2 2
20 9 9 13 13 4 3 9 1 2 11 9 0 13 4 13 13 4 9 13 2
22 11 11 9 13 2 11 13 4 12 15 9 2 9 9 0 1 10 9 9 0 13 2
14 12 9 2 11 3 13 4 11 2 7 12 13 4 2
18 10 9 2 11 9 13 13 7 2 9 13 2 13 9 13 13 4 2
9 11 11 2 7 2 9 13 4 2
34 9 10 1 2 9 14 4 9 9 0 13 2 10 9 12 13 10 9 10 9 13 4 3 1 2 9 2 9 2 9 7 9 2 2
13 11 9 0 13 4 13 9 9 13 7 3 13 2
17 13 9 0 13 9 9 3 9 12 13 4 10 9 13 0 9 2
13 9 2 9 1 2 13 9 13 13 4 9 9 2
21 2 9 10 9 14 13 0 2 9 0 13 9 1 2 7 9 10 9 13 4 2
10 9 9 2 9 12 1 13 4 9 2
19 9 13 9 13 11 9 2 10 3 2 12 13 7 9 12 9 9 13 2
15 14 4 9 3 0 13 2 7 11 0 13 4 9 10 2
15 9 10 9 9 13 9 13 4 11 2 3 9 9 1 2
4 3 9 10 2
15 9 10 9 13 13 4 7 9 2 10 1 2 0 9 2
21 2 0 14 13 14 13 15 9 13 7 14 2 9 9 0 13 9 9 0 13 2
13 3 13 4 0 2 9 1 3 13 3 13 4 2
19 9 9 9 9 9 13 4 2 7 9 3 13 3 13 13 4 9 1 2
9 11 11 13 4 14 4 13 13 2
12 10 13 4 3 1 2 3 7 3 9 13 2
15 11 9 13 4 9 9 7 3 9 13 4 0 9 13 2
13 11 9 13 13 9 13 9 12 13 4 9 0 2
11 9 1 2 9 2 13 13 13 4 11 2
17 13 13 2 9 0 1 2 9 0 9 13 4 13 11 9 9 2
11 7 9 9 2 9 1 2 9 0 13 2
19 9 0 1 9 9 13 4 9 2 0 9 0 2 7 10 14 13 13 2
14 10 2 11 12 13 4 11 11 9 9 2 11 1 2
28 11 9 9 9 13 9 14 13 13 4 11 7 3 11 11 1 10 9 2 13 7 9 9 13 2 9 13 2
5 7 13 9 13 2
14 11 11 11 13 4 9 12 2 11 1 2 9 13 2
18 9 11 13 4 9 10 2 7 9 9 1 2 11 13 4 12 9 2
21 11 9 3 10 13 9 1 2 12 9 9 9 13 4 9 9 13 4 9 0 2
16 10 9 2 3 11 7 11 11 11 13 4 11 9 13 4 2
14 9 9 1 11 1 9 0 14 4 13 11 9 12 2
13 11 11 11 9 2 7 2 9 13 4 2 3 2
22 0 2 9 7 9 10 13 9 9 13 4 9 7 9 1 9 12 9 2 9 9 2
17 13 4 9 9 10 1 12 13 9 0 7 0 9 12 13 3 2
27 11 9 9 12 9 11 9 9 13 4 9 13 13 2 7 11 11 12 9 9 3 9 13 4 9 9 2
13 11 7 11 9 12 13 4 7 11 7 11 10 2
25 9 0 7 13 13 13 2 13 2 13 13 4 11 8 11 2 7 10 1 7 13 4 9 9 2
9 11 14 4 15 13 11 9 1 2
8 9 10 13 4 12 9 10 2
22 9 0 13 13 4 11 7 9 9 10 9 13 3 2 9 13 4 9 11 12 9 2
25 7 2 9 13 3 11 13 4 2 9 0 7 9 1 13 4 2 7 3 9 7 9 0 13 2
16 11 11 9 9 13 13 13 2 13 4 2 13 2 13 11 2
11 11 12 9 9 9 13 2 13 9 9 2
10 2 9 9 7 9 13 9 13 2 2
11 9 1 9 13 9 13 4 11 7 11 2
15 3 2 9 9 9 10 15 9 9 13 12 9 1 9 2
20 11 11 11 9 7 11 9 13 4 9 9 1 2 3 13 4 12 13 9 2
10 10 1 13 11 2 11 11 9 13 2
18 9 12 9 1 2 11 9 9 0 0 13 4 2 12 7 11 9 2
13 9 9 13 14 4 2 3 13 4 9 1 13 2
24 11 11 9 3 13 9 13 13 9 11 11 13 9 7 10 9 0 11 13 13 0 9 1 2
11 3 2 12 9 2 11 11 9 13 4 2
14 11 11 11 12 7 11 11 11 11 13 4 3 9 2
10 9 13 9 12 9 13 4 9 11 2
17 10 13 4 11 9 0 0 9 9 13 9 10 1 9 9 13 2
14 15 11 9 12 3 13 2 11 9 9 2 13 4 2
20 11 1 9 10 13 4 11 9 2 7 3 13 4 9 10 11 11 9 9 2
18 15 9 2 7 2 3 1 13 4 2 9 1 13 2 7 10 13 2
22 11 11 9 2 11 9 2 9 0 13 2 7 11 7 11 11 9 3 13 13 2 2
11 11 11 2 3 13 3 9 9 13 9 2
10 2 6 6 2 15 13 4 9 10 2
26 11 9 11 9 9 13 9 12 9 13 9 1 2 9 0 12 9 9 9 7 9 9 9 9 13 2
16 9 9 13 4 9 12 8 9 13 2 3 3 9 1 13 2
12 3 13 7 9 1 2 12 9 13 4 11 2
13 9 7 9 9 12 9 13 7 9 7 12 9 2
13 11 11 9 13 4 13 2 9 0 9 13 9 2
14 11 9 2 11 11 13 12 9 9 1 13 12 9 2
11 11 11 11 11 0 13 4 13 4 3 2
7 11 11 13 4 11 9 2
24 9 12 13 4 0 9 2 7 3 3 9 13 9 13 2 12 7 11 12 13 4 9 11 2
18 11 0 0 9 9 9 13 13 2 9 9 2 7 13 9 13 13 2
9 0 11 11 9 7 0 13 4 2
19 9 13 9 11 11 11 9 2 3 2 13 4 9 13 2 7 2 11 2
13 11 7 11 2 13 9 2 13 4 11 1 9 2
20 11 11 9 13 13 4 9 13 4 2 3 2 11 9 13 13 4 9 13 2
15 11 11 11 9 13 9 3 9 13 4 11 7 11 1 2
14 3 1 9 13 14 4 9 13 13 10 13 4 9 2
12 11 9 9 13 4 9 9 1 9 13 9 2
12 11 11 9 11 1 13 12 9 9 13 11 2
10 9 2 9 1 13 4 9 10 9 2
9 12 9 3 9 10 9 13 4 2
24 11 9 9 0 9 13 13 2 7 2 9 10 1 2 12 9 10 12 9 13 9 13 4 2
8 13 4 9 0 12 9 1 2
14 2 11 9 9 13 7 9 10 9 10 13 4 2 2
10 9 2 3 3 2 9 0 13 9 2
9 3 9 12 9 13 4 11 11 2
21 11 13 4 2 2 3 9 11 1 13 4 2 7 9 12 14 4 10 13 2 2
18 7 2 9 7 9 9 4 9 0 9 12 7 10 13 7 13 13 2
13 9 12 13 4 3 3 13 2 7 9 13 4 2
25 11 11 2 9 9 13 13 2 12 9 13 4 2 7 10 10 9 9 13 4 9 0 10 1 2
18 0 9 3 13 14 7 2 9 9 9 9 10 13 4 11 12 9 2
13 11 9 2 9 7 2 13 4 13 4 11 9 2
24 0 9 9 3 3 13 13 9 10 2 3 0 13 4 9 11 2 11 7 9 9 9 9 2
17 11 13 4 9 13 9 9 2 7 3 14 13 9 2 0 7 2
10 3 13 4 9 10 11 2 11 11 2
14 9 9 0 7 10 9 3 13 13 3 13 9 9 2
15 2 12 7 9 9 13 4 2 11 3 0 13 9 10 2
15 11 11 11 2 11 2 13 4 12 9 2 12 9 0 2
20 11 11 9 9 2 9 0 13 2 12 5 2 9 9 13 7 13 9 13 2
17 11 11 3 13 4 11 9 9 13 2 7 9 13 4 13 4 2
22 11 11 9 13 4 11 11 9 13 11 7 10 9 12 9 14 13 11 13 13 4 2
13 9 0 13 2 7 2 14 4 0 13 12 9 2
25 9 0 2 9 0 2 13 2 9 10 9 13 4 13 2 15 1 3 2 10 9 9 3 13 2
30 10 9 2 9 0 2 12 7 2 14 4 13 9 9 13 2 11 2 11 7 11 2 7 2 9 0 13 9 13 2
12 9 10 1 3 13 4 11 11 11 9 9 2
15 0 9 11 11 13 4 9 14 13 3 13 9 13 9 2
20 9 0 0 10 9 9 7 13 4 9 2 7 3 3 13 13 9 10 3 2
35 9 9 9 0 1 13 9 13 13 4 2 7 3 13 4 9 0 1 13 4 9 2 9 10 2 10 9 0 9 9 13 13 4 2 2
27 7 2 11 11 9 11 2 11 7 11 11 14 4 13 3 13 7 2 9 2 9 10 9 12 13 4 2
28 3 0 13 2 7 12 1 11 9 13 11 11 12 9 9 2 9 12 10 1 13 7 11 13 9 13 4 2
11 9 13 12 13 4 9 2 0 7 9 2
10 13 4 9 10 12 9 1 13 4 2
8 3 2 11 9 9 13 4 2
11 9 11 11 11 9 9 7 13 4 9 2
15 11 1 2 11 9 7 9 0 13 4 13 9 0 13 2
7 11 9 14 13 3 0 2
14 12 9 12 9 13 13 4 9 11 11 2 11 2 2
13 11 11 11 2 11 9 9 9 11 13 4 3 2
9 9 1 13 4 9 9 13 4 2
15 11 9 9 10 9 0 13 2 9 9 0 1 9 13 2
18 2 13 9 13 4 2 14 13 10 9 13 2 7 10 0 13 4 2
17 3 1 12 9 9 13 9 3 13 4 2 9 9 9 13 9 2
18 12 9 9 13 9 2 9 9 15 1 13 4 13 13 4 11 0 2
14 9 9 13 9 11 2 7 12 9 1 11 13 4 2
19 13 4 7 9 0 13 2 7 12 1 13 13 15 7 13 9 13 4 2
21 15 13 4 9 13 9 11 11 9 13 13 4 3 7 3 11 11 9 11 9 2
16 9 10 9 12 13 2 9 2 9 2 9 7 9 14 13 2
24 2 9 9 12 8 9 10 13 15 7 9 10 9 0 7 13 2 15 10 9 13 7 2 2
16 11 9 9 9 0 13 13 9 4 13 11 0 9 9 9 2
17 9 0 1 0 13 4 11 7 11 12 9 13 4 9 9 1 2
14 9 1 13 4 9 3 13 4 11 11 11 9 11 2
24 9 2 9 13 11 9 9 9 9 13 14 7 2 10 9 13 9 9 10 9 13 4 13 2
10 3 9 1 13 4 2 10 9 10 2
6 9 13 3 13 4 2
20 11 11 11 11 9 13 4 2 2 15 9 13 9 13 4 13 9 13 2 2
11 3 9 2 11 11 7 11 11 13 4 2
12 9 0 1 13 4 9 13 7 13 7 13 2
25 11 11 9 7 11 9 13 12 9 13 4 2 9 9 13 9 13 4 11 2 11 1 9 13 2
9 3 9 10 9 13 4 9 10 2
19 9 0 10 11 11 13 4 2 11 9 0 3 2 7 9 9 0 9 2
13 11 11 12 13 4 2 7 11 0 13 4 12 2
12 11 9 9 11 11 9 13 4 12 9 9 2
8 9 1 9 13 9 10 13 2
30 3 2 10 9 2 2 0 10 13 4 13 4 2 15 9 13 4 9 7 9 13 9 13 9 10 9 13 4 2 2
11 9 13 9 9 1 13 7 9 13 4 2
13 9 9 13 9 9 2 0 9 10 1 13 4 2
11 2 3 9 7 9 13 4 9 1 2 2
11 10 13 4 11 3 13 0 4 0 9 2
13 12 9 2 11 9 9 7 11 9 13 9 9 2
9 9 12 13 4 9 12 9 9 2
10 9 9 3 0 13 4 9 9 9 2
22 11 11 12 9 11 7 11 2 3 12 9 2 3 13 13 4 0 0 9 1 9 2
23 3 1 13 9 0 7 0 13 9 0 0 7 2 10 1 2 9 9 10 13 4 2 2
17 9 3 13 4 9 13 4 2 7 11 9 13 13 4 9 1 2
8 9 9 13 4 9 0 3 2
10 12 9 7 12 9 13 4 12 10 2
17 11 11 9 12 7 9 1 13 4 9 2 9 13 3 9 13 2
7 10 9 12 11 11 13 2
18 11 11 11 11 9 0 13 0 13 4 10 9 9 11 0 9 0 2
22 11 1 2 11 3 13 4 9 2 7 3 9 2 3 13 2 13 4 13 11 9 2
25 9 10 2 12 9 12 13 3 2 12 9 13 4 9 10 2 3 0 0 9 13 0 9 13 2
23 9 12 12 9 2 12 12 9 2 13 4 11 2 11 7 11 11 0 9 13 4 3 2
15 7 2 9 10 9 0 9 1 11 13 13 4 11 11 2
16 11 3 9 13 13 4 11 9 2 9 10 9 13 9 13 2
13 2 9 13 11 1 13 2 11 3 9 0 13 2
10 11 11 9 9 13 4 3 9 9 2
17 13 4 9 12 9 13 4 9 10 2 11 2 11 12 9 9 2
35 3 2 9 9 2 12 9 12 9 2 9 9 12 7 9 12 13 2 7 11 13 9 10 13 2 11 11 13 9 13 9 0 13 4 2
12 11 9 13 9 9 11 9 9 13 4 3 2
33 7 9 13 4 2 2 11 9 9 13 9 9 13 13 4 2 9 0 13 11 9 9 1 7 10 9 9 13 9 13 4 2 2
20 11 11 11 14 4 12 9 13 2 7 0 9 9 12 9 0 13 2 9 2
17 12 9 11 11 13 4 2 12 2 7 12 11 11 2 12 2 2
10 3 2 7 2 0 9 3 13 4 2
20 11 12 9 13 4 12 9 13 2 12 9 2 12 12 9 7 9 12 2 2
18 7 2 14 13 15 0 9 2 9 10 13 2 7 10 14 13 0 2
18 0 9 0 2 11 0 13 4 7 9 1 2 11 12 9 13 4 2
14 3 13 4 9 7 3 13 13 4 9 10 9 13 2
35 9 0 9 13 13 13 13 4 11 2 7 9 12 9 13 4 12 9 13 2 11 11 12 9 9 13 0 13 4 2 12 9 12 13 2
13 3 2 11 9 1 9 12 3 13 4 13 4 2
10 11 9 12 9 9 13 4 11 9 2
25 11 11 11 9 12 2 11 11 2 13 4 9 11 11 2 9 9 7 11 9 9 9 10 2 2
20 9 9 9 9 3 7 3 11 9 9 9 13 13 4 2 11 2 11 2 2
14 11 0 11 11 13 9 13 4 3 9 12 11 9 2
17 11 9 9 9 13 2 7 3 9 0 9 1 9 10 13 4 2
13 11 9 13 4 2 7 2 7 11 9 13 4 2
19 7 9 10 13 4 13 3 13 12 9 2 11 11 11 9 9 13 4 2
13 9 9 9 9 12 9 13 4 11 7 11 1 2
23 9 3 13 9 13 4 11 9 0 7 10 13 9 2 9 0 12 9 13 4 9 1 2
7 11 11 13 4 11 9 2
6 3 9 9 9 13 2
7 13 13 4 2 14 9 2
16 7 11 13 9 13 4 2 11 11 1 2 11 9 0 7 2
16 10 13 4 3 9 11 9 9 7 9 0 1 13 9 13 2
7 3 2 3 8 3 13 2
27 9 12 11 9 10 9 12 13 4 2 10 12 2 7 2 9 12 3 12 9 10 1 0 13 9 13 2
10 13 9 13 9 9 1 7 13 9 2
37 9 1 13 2 0 13 2 3 9 0 2 0 2 9 9 9 7 15 0 2 9 0 7 0 13 2 3 9 9 13 7 0 13 9 13 4 2
8 12 12 9 12 13 4 10 2
17 11 9 0 13 9 1 2 9 0 12 9 13 4 12 9 1 2
17 9 10 9 1 2 12 13 4 3 13 11 2 11 2 9 0 2
10 9 9 13 11 9 9 0 13 4 2
18 9 10 13 4 14 4 13 13 2 7 7 9 13 4 9 13 13 2
11 9 14 13 3 2 7 14 3 13 9 2
21 11 11 11 9 9 0 9 0 9 9 13 4 11 9 9 2 9 1 9 13 2
23 9 9 13 4 2 9 9 14 13 9 12 13 4 2 3 2 10 10 2 9 9 13 2
15 11 11 12 13 4 9 12 9 7 3 0 9 7 13 2
19 7 11 12 9 2 11 11 7 11 11 2 9 9 9 13 9 13 4 2
11 9 9 13 13 2 7 14 13 11 11 2
20 7 2 3 2 9 14 4 3 13 2 9 9 1 9 9 9 0 13 4 2
13 9 9 11 11 9 13 7 9 9 12 9 13 2
34 10 1 2 11 13 4 11 3 13 9 2 3 3 2 13 2 11 2 9 9 0 2 13 2 7 12 1 2 9 9 0 2 13 2
22 11 9 12 7 12 3 9 13 4 7 10 10 9 7 9 9 13 9 13 9 13 2
16 11 0 13 9 9 2 12 7 9 13 9 9 3 0 13 2
15 3 13 9 12 1 13 13 7 9 11 11 9 9 13 2
19 11 9 0 13 13 4 9 13 4 2 7 3 1 9 1 13 4 11 2
21 7 12 9 1 11 2 11 7 11 9 13 13 4 2 7 11 2 7 2 13 2
14 11 12 9 13 9 11 2 7 12 9 13 12 9 2
12 11 11 13 9 13 9 1 2 13 2 13 2
12 10 2 10 9 9 1 0 9 13 13 4 2
13 3 2 12 9 9 13 4 2 7 3 9 0 2
17 11 13 9 13 11 9 9 10 13 2 7 3 13 4 9 0 2
13 9 1 2 9 13 2 9 2 13 4 13 4 2
23 9 10 2 2 9 1 7 9 1 9 2 9 1 9 7 9 0 9 2 13 4 11 2
12 11 11 7 11 11 3 13 4 9 10 9 2
38 7 9 13 3 2 10 0 9 13 4 13 4 11 2 3 2 9 9 13 9 9 9 13 11 11 7 2 9 10 13 2 9 0 9 13 2 12 2
18 9 0 11 11 13 4 2 7 3 1 12 9 9 9 0 13 4 2
16 9 7 9 9 11 9 1 13 9 13 4 3 11 9 0 2
12 3 2 9 9 2 3 13 14 4 9 1 2
21 9 9 9 9 9 13 4 11 2 12 7 9 12 9 7 9 9 13 4 9 2
29 11 9 13 9 2 11 9 3 9 13 9 0 11 13 4 9 1 2 7 9 9 0 13 9 0 13 4 9 2
21 9 2 12 9 9 7 9 13 4 2 7 9 9 13 4 9 9 7 9 9 2
9 7 2 12 1 9 10 13 4 2
16 11 13 7 9 13 4 3 3 9 7 10 9 13 13 3 2
13 9 9 13 12 7 12 9 9 3 0 13 4 2
22 12 9 9 13 9 14 4 13 2 7 2 9 9 13 2 7 11 13 4 10 1 2
12 3 2 11 11 12 12 9 9 13 4 11 2
20 11 1 9 10 11 11 9 3 13 4 9 2 0 9 13 0 9 11 9 2
23 12 11 8 11 7 11 11 11 13 4 12 12 9 9 13 9 10 2 7 12 9 11 2
5 11 12 13 13 2
19 7 2 11 9 14 4 13 10 3 9 13 11 9 12 2 9 9 13 2
17 9 0 9 9 2 9 9 7 9 9 13 13 4 13 4 11 2
22 11 9 11 12 0 9 13 4 12 9 2 7 10 12 3 3 13 4 2 9 1 2
9 3 2 15 9 1 13 9 10 2
19 9 9 9 9 1 13 4 11 2 3 9 9 13 2 3 14 15 9 2
9 9 0 10 1 9 9 13 4 2
13 2 9 0 1 9 13 7 9 9 13 4 2 2
22 11 11 11 0 1 2 2 11 9 9 13 4 13 13 9 13 11 11 11 9 2 2
18 11 11 2 11 7 9 0 9 9 7 9 0 13 4 11 9 1 2
20 11 8 11 9 9 0 14 4 13 13 11 9 2 7 9 4 11 11 9 2
18 2 9 9 13 4 7 3 9 2 3 2 9 9 12 13 4 9 2
17 10 1 9 0 7 9 0 13 4 9 0 13 4 10 13 13 2
25 2 15 10 9 9 0 13 4 11 11 13 4 2 9 9 0 12 13 4 2 2 13 4 11 2
14 11 9 13 4 9 9 3 0 13 11 11 9 0 2
17 10 13 7 9 13 9 9 7 9 1 13 4 9 0 0 13 2
19 12 12 1 12 9 13 4 7 12 9 3 13 4 11 9 9 13 13 2
15 9 3 13 4 11 9 1 2 7 14 4 3 7 13 2
13 11 11 12 13 4 2 7 11 13 7 13 4 2
18 11 9 10 2 7 2 3 0 13 15 2 3 3 9 7 9 0 2
12 9 9 7 0 9 9 13 7 13 4 9 2
16 12 2 11 11 9 9 13 4 2 9 9 9 9 13 4 2
25 11 9 11 13 4 3 2 9 9 9 2 7 13 4 11 9 13 11 13 4 9 1 14 13 2
8 10 1 15 13 9 13 11 2
12 11 4 13 9 12 2 3 12 12 13 4 2
8 11 11 11 9 13 9 13 2
19 9 0 9 2 7 2 9 13 4 9 2 7 10 13 9 13 9 0 2
24 9 7 9 9 13 2 13 7 2 9 2 9 7 9 9 0 3 13 4 2 9 13 7 2
17 9 10 9 9 0 7 9 9 13 9 9 9 9 13 4 9 2
5 11 11 13 13 2
13 0 12 0 13 2 7 2 9 13 4 11 9 2
7 7 3 13 10 9 13 2
16 2 11 9 13 13 13 2 7 9 1 8 14 4 13 2 2
14 10 3 2 11 9 0 13 4 2 7 9 0 0 2
34 11 11 11 13 4 2 2 11 7 11 9 9 13 4 9 0 9 13 7 9 9 7 9 13 4 9 9 0 9 13 13 4 2 2
7 13 11 9 1 11 12 2
15 11 2 12 9 9 13 4 11 11 2 3 11 9 13 2
20 9 2 9 9 9 9 3 10 9 10 13 4 2 11 9 14 13 3 13 2
17 9 11 13 9 12 9 9 3 2 11 9 9 13 4 12 9 2
14 7 2 3 3 2 2 9 13 2 13 4 9 0 2
8 10 10 14 13 9 9 10 2
19 9 7 9 14 13 10 9 10 2 11 2 9 9 13 12 0 9 13 2
17 9 2 9 9 7 0 9 9 14 7 9 9 10 13 13 4 2
8 9 9 9 14 4 0 13 2
25 11 11 11 9 11 9 12 0 13 13 4 3 2 7 11 12 7 11 13 9 10 13 13 4 2
16 0 9 2 9 2 9 7 9 13 2 9 10 9 1 13 2
9 10 1 14 13 10 9 9 13 2
10 9 13 12 13 4 9 13 4 9 2
12 12 9 0 7 12 9 13 4 9 0 9 2
13 13 0 13 4 2 7 0 13 2 11 13 9 2
20 11 9 9 11 13 0 13 13 4 9 2 7 11 11 11 9 14 13 4 2
24 3 7 3 9 13 9 13 13 4 7 2 12 9 7 9 12 9 3 13 4 12 12 9 2
17 11 9 10 13 4 9 3 2 7 11 1 9 13 4 13 4 2
30 12 12 9 11 13 4 9 0 7 0 13 4 3 2 9 10 10 12 9 9 13 9 13 9 0 0 2 11 2 2
19 2 3 9 0 1 9 13 4 9 7 3 2 7 2 3 0 13 2 2
12 9 9 10 12 9 13 9 13 4 10 1 2
25 10 9 2 2 11 3 0 13 4 11 11 2 2 7 7 2 0 9 14 2 4 13 9 0 2
24 11 9 0 13 4 0 11 7 10 12 13 13 4 2 11 10 9 13 4 9 13 13 4 2
15 3 3 3 13 7 13 4 9 9 9 9 13 4 13 2
21 2 11 13 9 13 4 9 0 9 12 9 13 7 10 9 13 4 9 9 2 2
23 0 0 11 13 7 9 0 9 9 13 13 9 1 2 3 3 9 9 9 13 4 3 2
16 3 3 13 2 7 12 7 3 13 3 2 9 3 0 13 2
16 2 15 13 4 13 9 9 2 13 4 9 10 13 13 4 2
6 9 1 13 4 9 2
18 9 12 9 9 13 7 9 0 13 4 3 2 12 9 1 13 9 2
6 3 7 3 13 4 2
20 11 11 12 13 4 2 11 13 4 12 9 9 2 11 12 9 13 13 4 2
11 9 7 9 1 2 9 9 0 13 4 2
21 3 9 14 4 13 11 9 0 15 13 2 3 9 9 15 14 4 9 0 13 2
8 9 13 4 11 11 13 9 2
12 11 11 11 7 13 4 2 7 13 13 4 2
12 9 9 9 13 13 4 11 9 9 13 9 2
19 9 9 9 7 9 9 13 4 9 9 2 9 0 12 13 4 10 1 2
15 7 2 3 9 12 1 2 11 0 13 13 9 13 4 2
18 11 9 0 13 4 11 9 2 7 2 9 1 2 13 4 13 4 2
8 9 0 12 13 10 1 9 2
28 9 9 0 9 13 4 3 13 9 13 9 9 1 9 3 11 9 2 0 0 7 12 9 13 4 9 0 2
16 9 12 13 4 2 3 2 9 11 12 9 9 2 11 2 2
13 9 9 2 11 9 0 13 4 9 0 9 1 2
23 3 2 0 9 11 3 0 9 0 13 9 13 4 11 2 7 9 0 9 0 13 4 2
14 11 11 2 11 2 13 4 3 1 9 9 9 9 2
10 9 1 2 9 12 3 13 9 12 2
8 11 11 8 12 9 0 13 2
24 15 9 13 9 9 10 9 13 13 13 7 0 9 10 13 2 10 9 9 9 0 13 2 2
7 12 9 3 9 13 10 2
18 11 13 9 13 3 2 0 15 13 2 7 14 2 8 3 2 11 2
30 9 9 9 12 13 4 9 9 14 13 9 12 13 4 9 1 2 7 13 3 13 4 9 7 9 12 13 4 9 2
10 7 11 9 14 4 9 9 1 13 2
8 12 12 13 11 9 13 4 2
13 9 10 0 13 2 7 3 12 2 11 9 9 2
28 11 9 11 13 9 0 12 9 13 13 2 7 13 9 9 9 14 13 2 0 9 3 13 4 2 11 3 2
23 10 9 2 0 13 9 9 9 3 9 12 9 13 7 14 12 9 3 3 13 4 3 2
23 9 1 9 13 9 13 9 0 9 13 9 1 13 2 7 7 9 0 7 9 13 4 2
9 12 9 9 13 4 9 12 1 2
7 7 11 9 9 13 4 2
9 2 10 7 10 13 4 9 1 2
11 11 11 9 2 9 0 13 9 13 4 2
26 9 9 9 0 9 9 12 13 4 2 11 2 11 2 2 7 11 11 11 12 10 1 13 13 3 2
19 9 12 1 13 4 7 11 8 11 7 11 9 11 9 13 4 10 10 2
15 9 9 9 3 13 2 9 1 13 4 12 9 11 11 2
19 11 9 0 0 9 0 13 8 4 2 3 9 0 2 11 7 11 3 2
18 11 11 13 13 4 11 2 11 11 1 2 12 2 12 7 12 2 2
17 9 1 2 9 9 11 9 9 13 4 2 3 13 4 9 9 2
28 11 2 9 1 2 13 4 9 2 9 1 2 9 9 9 2 13 4 2 7 9 1 9 9 9 13 13 2
36 11 11 2 12 5 2 2 11 11 11 2 9 2 2 11 11 2 9 2 7 11 11 2 9 9 2 3 13 11 11 9 13 15 12 9 2
12 11 2 11 7 11 9 9 12 1 13 4 2
9 9 12 9 1 2 9 9 13 2
9 9 1 13 7 9 0 13 4 2
20 9 9 7 9 13 2 12 9 10 9 13 9 13 4 2 9 13 13 9 2
5 9 1 13 4 2
12 11 12 7 11 2 11 7 11 12 13 4 2
11 3 2 11 7 0 1 13 4 3 1 2
14 9 0 9 13 9 9 13 2 12 7 9 2 8 2
11 9 9 1 13 4 7 9 13 13 4 2
13 11 11 9 11 12 7 11 12 13 13 4 11 2
18 9 1 2 9 0 12 13 7 9 10 1 9 9 0 12 13 15 2
15 10 1 11 9 11 11 7 9 0 10 12 9 13 4 2
11 11 9 1 2 2 9 9 9 13 4 2
17 11 11 11 9 0 9 9 13 4 7 14 13 4 3 9 0 2
20 9 3 2 3 13 13 13 2 7 13 4 9 0 2 9 3 13 2 13 2
19 3 13 2 7 2 9 3 0 13 7 9 0 2 13 4 9 9 13 2
18 9 0 9 12 9 9 13 4 2 7 11 7 11 13 4 3 9 2
23 9 9 13 9 11 13 4 9 3 12 9 13 4 11 2 12 13 4 11 9 9 9 2
22 3 7 2 9 0 12 1 9 12 13 9 12 4 9 13 9 0 12 9 13 4 2
18 0 10 3 13 4 9 12 9 7 9 1 2 7 10 13 4 7 2
15 11 9 13 4 13 4 2 9 10 0 13 9 1 2 2
16 11 7 11 1 9 13 9 12 9 13 4 3 11 2 11 2
15 9 10 13 4 2 11 12 9 1 9 9 13 9 13 2
10 9 2 0 14 4 9 1 13 9 2
20 7 2 11 11 11 9 2 9 9 12 13 4 2 11 11 0 9 0 13 2
10 15 7 2 3 1 9 13 13 9 2
20 3 13 4 3 11 11 11 9 9 0 7 9 11 9 9 11 9 9 9 2
23 11 11 0 2 11 2 13 4 0 2 11 11 2 11 2 7 11 11 2 11 2 9 2
7 14 13 3 2 7 3 2
15 9 9 13 4 13 13 4 9 2 13 7 2 13 13 2
21 9 2 9 2 9 2 9 0 7 0 2 9 2 9 2 9 10 13 9 1 2
18 11 11 2 9 0 2 7 2 9 3 13 2 13 4 13 4 11 2
31 9 9 2 7 2 11 11 9 9 14 13 13 3 2 11 11 9 13 9 13 4 11 9 10 9 2 9 13 4 7 2
14 9 10 1 9 13 11 11 9 10 9 13 13 4 2
11 3 2 7 2 11 11 7 11 11 13 2
8 9 0 12 13 3 10 1 2
13 11 11 11 13 4 9 9 9 9 2 12 2 2
23 11 9 9 15 9 7 9 13 4 3 11 11 9 9 13 9 13 15 9 13 4 9 2
23 0 9 9 3 9 13 7 9 13 13 4 2 7 9 12 2 12 7 12 7 13 4 2
24 11 9 13 13 4 3 9 0 13 4 13 4 2 7 3 9 9 12 11 10 13 13 4 2
16 7 11 1 2 9 10 14 13 0 2 13 4 9 3 13 2
21 10 13 7 2 11 11 9 12 13 7 9 0 12 13 9 2 14 4 3 13 2
22 9 10 2 9 1 13 9 10 9 0 0 9 7 9 13 4 2 13 9 13 9 2
10 2 9 1 9 0 13 9 13 2 2
12 9 3 0 13 4 3 11 1 9 13 9 2
16 9 9 13 7 13 4 2 3 13 4 3 9 0 7 0 2
20 10 9 0 3 0 13 7 9 9 0 1 13 4 7 3 0 13 9 13 2
17 9 2 11 12 9 12 13 9 9 7 3 11 9 13 13 4 2
24 3 13 4 12 9 12 0 9 13 9 9 13 9 10 2 13 7 2 9 10 3 13 4 2
19 2 9 1 9 13 2 9 13 13 4 9 12 7 12 9 13 4 9 2
14 9 3 7 3 13 4 2 7 12 7 9 0 12 2
16 10 2 3 7 3 13 4 3 9 13 4 9 11 13 4 2
13 11 9 0 12 13 13 4 9 2 11 9 1 2
7 11 7 11 15 1 13 2
13 12 9 12 13 4 11 1 2 7 12 11 1 2
19 3 2 3 3 2 9 14 13 3 13 9 13 7 2 15 9 13 4 2
10 11 11 12 12 9 13 4 11 9 2
7 0 2 9 1 13 4 2
14 9 9 15 13 13 4 2 7 9 12 1 13 4 2
14 15 13 4 9 0 13 4 2 10 0 13 7 9 2
7 10 10 10 13 13 4 2
17 9 12 9 13 4 9 3 9 13 4 11 11 7 11 11 3 2
30 3 3 2 11 9 9 13 4 11 2 13 13 4 9 9 11 9 10 10 9 13 2 7 9 14 4 13 10 9 2
29 3 13 4 2 10 10 2 11 11 7 11 11 11 9 2 11 11 11 7 11 11 9 7 11 11 11 9 0 2
10 11 9 9 9 14 4 15 3 13 2
12 9 1 13 4 3 7 9 10 13 9 1 2
10 11 7 2 12 9 9 9 13 4 2
17 12 2 9 9 12 13 2 9 10 9 12 13 7 13 13 4 2
17 9 13 13 9 9 0 13 13 2 3 7 2 9 9 13 9 2
19 9 2 3 13 13 9 13 2 7 9 0 0 3 3 13 13 3 13 2
20 9 9 9 9 7 11 11 7 11 3 3 7 0 13 4 9 9 9 3 2
15 9 10 2 12 9 9 11 9 9 9 13 4 13 4 2
24 3 13 4 11 9 10 1 9 2 7 2 3 15 13 14 4 7 2 10 9 13 4 13 2
18 9 11 11 13 9 7 9 13 9 2 9 13 9 13 7 13 4 2
25 11 9 11 2 9 2 11 11 2 9 7 11 11 2 9 2 13 4 9 1 9 9 13 9 2
16 10 10 9 13 13 9 2 0 9 9 1 9 13 13 4 2
32 12 9 13 13 4 2 7 11 1 13 14 4 7 2 9 1 9 9 13 13 13 4 2 7 10 3 13 4 9 13 4 2
9 11 0 1 13 9 9 13 4 2
6 13 10 13 4 13 2
20 11 9 1 11 8 11 13 4 13 4 12 2 7 10 1 11 0 13 4 2
30 11 10 13 4 9 2 7 10 9 0 13 4 2 7 13 4 10 9 11 11 13 9 2 0 2 10 13 4 9 2
10 11 1 2 9 9 10 13 4 9 2
9 2 11 11 1 13 9 13 4 2
8 11 11 2 11 13 4 13 2
18 11 11 9 13 13 9 11 2 11 9 0 13 2 13 4 13 4 2
9 10 2 10 9 13 4 9 1 2
20 12 9 12 9 12 11 13 4 2 12 2 2 3 9 9 13 4 9 1 2
12 9 13 4 9 0 10 1 10 0 13 9 2
15 9 13 4 13 9 12 9 12 13 4 11 11 9 0 2
11 11 9 3 0 13 10 1 9 12 13 2
9 11 9 9 13 11 11 11 9 2
34 11 9 14 4 3 9 0 9 2 11 2 13 9 13 9 13 9 2 7 11 11 9 11 11 9 0 13 4 11 12 9 13 4 2
21 9 13 3 13 4 2 9 2 3 2 7 9 2 11 9 0 1 13 13 4 2
10 12 8 3 9 0 13 4 9 11 2
11 11 11 0 13 9 9 0 2 11 1 2
13 9 3 13 7 2 10 1 9 0 13 15 13 2
25 11 9 9 10 2 9 13 4 7 9 9 7 2 7 9 9 13 15 9 7 9 9 13 2 2
32 9 0 2 0 7 0 13 7 3 9 7 9 13 0 13 2 7 3 11 9 14 4 13 2 3 9 9 9 13 4 2 2
14 2 9 0 13 11 2 7 11 9 13 13 9 13 2
10 12 10 12 1 13 9 13 4 3 2
12 0 12 9 13 2 9 13 13 4 9 1 2
17 12 9 9 9 0 1 2 11 3 13 4 10 9 1 12 9 2
19 11 9 11 11 3 13 4 2 7 2 10 9 9 12 9 9 13 11 2
12 0 13 9 11 11 7 11 9 1 9 9 2
31 9 4 9 9 10 2 7 9 0 2 9 12 13 4 9 0 2 7 9 13 4 13 2 3 3 0 2 3 3 0 2
9 9 12 1 13 4 13 9 10 2
13 11 9 9 11 9 13 4 7 9 10 13 4 2
23 11 9 9 2 12 9 9 14 4 9 13 0 2 7 10 9 13 4 12 9 9 9 2
23 3 2 11 11 7 11 11 9 13 2 12 9 9 13 9 13 4 9 12 9 0 10 2
18 9 7 11 13 9 14 7 2 9 9 7 12 9 13 4 13 4 2
8 11 11 9 12 9 13 4 2
13 11 11 1 10 9 2 13 2 9 13 11 9 2
13 7 3 7 9 0 13 9 9 8 9 13 9 2
11 7 2 13 2 3 1 0 9 13 4 2
17 9 3 9 0 13 2 9 0 2 9 2 7 9 1 9 10 2
7 15 1 13 4 13 4 2
9 9 13 4 2 9 3 13 4 2
24 9 10 2 14 4 3 0 13 11 9 9 13 2 9 9 9 13 4 9 7 13 4 13 2
23 10 2 9 11 9 9 13 4 2 9 9 11 9 13 4 9 7 9 1 9 13 4 2
20 12 9 13 4 2 9 10 10 2 11 1 10 12 9 2 7 13 13 4 2
13 11 9 12 9 9 13 9 13 3 11 2 11 2
16 9 13 4 9 2 11 9 2 9 7 9 1 9 9 13 2
7 2 9 13 9 13 4 2
17 9 9 2 11 11 13 4 12 9 10 9 3 7 3 13 4 2
17 0 13 4 10 9 2 11 11 2 13 12 9 11 11 9 9 2
14 11 10 2 12 9 9 13 4 2 9 10 13 4 2
7 11 11 11 13 10 9 2
11 11 12 13 2 12 2 11 7 11 1 2
30 9 9 2 11 13 7 13 9 13 4 2 2 7 11 13 9 13 4 2 9 0 9 9 13 4 12 9 9 1 2
33 2 9 9 10 1 9 9 13 4 9 9 2 9 10 13 9 7 9 7 9 9 12 4 13 2 9 10 13 4 9 13 9 2
9 9 9 9 15 13 4 13 11 2
5 13 13 9 12 2
18 11 9 12 13 4 9 0 1 7 11 11 9 9 13 4 9 13 2
10 11 13 13 9 11 10 2 15 9 2
29 9 9 9 9 13 4 2 9 0 9 7 11 9 2 2 9 1 2 7 9 3 1 0 13 4 9 13 4 2
10 9 0 13 4 9 9 12 13 4 2
12 7 2 3 9 1 2 3 9 13 13 4 2
14 9 13 13 4 3 11 9 7 11 13 9 13 9 2
11 12 11 11 12 11 9 11 11 13 4 2
23 9 9 2 12 7 12 9 1 9 9 12 0 9 12 13 4 2 11 9 2 9 2 2
14 9 9 9 12 9 13 4 11 9 1 2 9 12 2
8 9 1 9 13 4 11 9 2
25 3 7 9 0 13 4 0 9 2 7 3 13 9 13 9 9 9 0 9 2 12 9 13 3 2
14 9 10 2 9 0 12 13 4 2 9 12 13 3 2
16 12 7 12 9 13 4 12 9 13 7 2 11 11 13 4 2
9 3 3 13 4 2 12 9 0 2
33 9 2 7 12 12 9 13 13 4 2 13 7 2 11 9 3 9 13 4 2 7 7 2 9 1 2 9 9 13 0 9 13 2
12 7 2 0 13 11 14 13 9 10 0 9 2
9 9 9 0 7 9 10 13 4 2
23 13 13 11 11 9 0 9 13 4 2 7 3 12 9 13 9 2 9 7 9 13 3 2
19 9 1 2 11 12 9 13 4 2 7 3 7 11 9 0 13 13 4 2
28 3 2 9 9 12 13 9 2 12 11 9 13 13 4 3 11 2 12 11 9 0 9 2 7 12 9 9 2
17 11 11 13 7 2 3 2 9 1 13 4 2 3 13 4 9 2
12 2 14 4 3 0 13 2 11 11 2 2 2
26 11 9 2 9 13 13 9 2 3 9 0 2 13 4 9 0 2 7 11 11 0 13 4 15 13 2
9 10 13 4 13 15 9 9 12 2
14 11 9 1 10 9 9 0 13 4 9 12 13 4 2
13 3 12 9 13 11 9 0 2 7 12 9 11 2
11 3 2 11 12 9 9 13 4 9 1 2
10 12 9 1 3 13 4 11 13 4 2
18 12 7 12 9 1 9 10 13 4 11 11 2 7 14 4 9 13 2
25 9 1 9 9 0 13 9 13 9 13 2 9 0 13 4 9 0 13 7 9 10 9 0 13 2
35 2 9 0 13 2 7 10 9 13 9 13 2 7 2 9 13 9 3 0 13 4 9 13 2 13 4 2 7 2 11 11 10 9 12 2
19 7 0 13 9 13 4 0 9 1 2 7 7 3 9 14 4 0 13 2
14 9 10 0 9 13 9 10 13 4 2 9 13 7 2
18 9 9 1 13 11 3 9 7 3 13 4 9 9 10 9 13 4 2
16 9 2 9 1 2 9 13 13 4 9 1 2 9 9 12 2
9 11 11 7 9 0 13 4 3 2
23 10 1 2 11 13 4 2 0 2 13 11 1 9 13 2 2 11 11 9 13 8 2 2
11 11 9 0 13 4 3 9 9 0 13 2
18 12 11 9 13 4 11 0 13 4 3 11 11 11 9 2 12 13 2
10 12 3 9 0 13 4 7 12 13 2
22 9 14 13 7 9 12 9 9 0 13 13 4 2 15 0 9 13 9 7 9 1 2
21 3 2 11 11 11 9 12 9 13 4 2 3 15 9 7 11 9 13 4 2 2
18 3 1 11 9 3 13 7 2 11 14 13 9 0 13 4 9 0 2
7 11 11 9 0 13 4 2
24 9 13 4 2 7 13 13 9 9 13 4 2 10 11 9 13 13 4 2 7 0 13 4 2
22 11 2 3 2 3 12 9 15 1 13 9 10 1 9 0 13 7 9 13 9 13 2
18 12 9 9 0 2 7 9 2 12 9 2 0 13 9 9 0 13 2
10 9 1 2 9 9 0 13 4 11 2
13 11 11 9 0 13 4 9 0 10 9 10 13 2
30 2 3 3 2 13 4 11 9 2 12 7 10 9 10 9 13 4 11 11 9 2 7 10 9 13 13 13 13 4 2
11 9 3 1 13 4 2 7 12 13 4 2
24 11 11 13 4 2 9 12 2 9 13 9 13 13 2 7 12 9 13 13 3 11 13 4 2
21 11 1 2 12 9 9 13 4 11 7 11 9 7 11 2 11 7 11 11 9 2
14 3 2 3 2 13 15 9 2 14 4 9 0 13 2
10 9 9 1 13 7 2 14 4 13 2
11 11 7 12 9 1 13 4 9 1 13 2
23 3 13 4 9 13 2 7 2 10 3 7 2 9 13 4 3 9 12 9 13 4 10 2
12 9 0 13 4 14 4 9 13 11 9 9 2
11 9 1 2 9 10 9 10 7 13 4 2
22 11 9 2 9 9 0 0 13 2 9 1 2 9 12 9 1 13 4 9 13 4 2
20 11 11 11 9 12 3 13 9 13 4 2 11 9 9 9 9 9 13 4 2
15 11 11 3 1 12 9 9 13 4 7 12 9 13 4 2
15 11 9 13 13 13 4 12 9 7 9 9 0 13 4 2
25 12 9 9 2 11 9 13 4 9 1 12 9 13 2 12 7 2 11 9 9 13 4 12 9 2
7 2 0 9 1 13 10 2
10 11 12 7 11 13 0 9 3 9 2
16 9 13 4 2 9 9 9 2 11 11 2 2 3 9 9 2
23 10 2 11 13 4 13 9 7 11 0 1 11 13 4 9 2 7 0 10 13 9 13 2
9 10 13 13 4 0 9 11 11 2
16 10 2 11 3 1 0 13 4 9 7 9 13 13 4 11 2
11 9 9 9 9 13 4 2 3 3 1 2
23 11 11 11 2 11 11 7 11 11 13 14 4 7 2 9 0 12 13 4 3 9 9 2
11 11 11 9 13 4 11 12 9 13 3 2
11 3 2 11 1 2 11 13 4 11 9 2
19 2 3 9 2 9 13 4 11 9 2 7 11 10 2 12 9 1 9 2
15 11 9 13 13 9 13 9 12 9 12 13 4 9 0 2
6 3 0 13 13 4 2
9 0 11 13 4 9 2 11 11 2
16 9 9 3 9 9 9 12 9 13 4 3 2 11 11 9 2
14 11 1 2 11 7 11 9 0 13 4 9 1 9 2
31 10 1 4 9 13 4 13 2 11 11 11 2 11 9 9 13 7 9 13 4 2 9 12 12 9 9 3 13 13 4 2
23 3 9 9 14 13 9 2 7 9 3 13 9 9 13 2 2 13 13 4 9 12 2 2
13 11 13 9 12 13 4 9 0 2 12 9 9 2
14 9 10 9 9 0 11 11 11 9 9 9 13 4 2
21 11 11 0 13 4 11 9 11 9 13 4 9 2 3 11 11 9 0 13 4 2
18 7 2 3 1 13 4 11 2 7 10 9 10 13 3 13 4 9 2
17 11 7 11 13 4 2 7 9 13 15 7 3 9 0 13 4 2
12 9 3 13 2 9 1 10 9 13 9 13 2
22 11 11 13 4 9 9 0 13 2 7 9 13 13 11 9 0 13 4 9 12 11 2
10 2 3 7 15 1 13 9 13 10 2
14 9 3 9 13 4 9 7 9 0 10 9 1 13 2
14 11 9 3 7 11 9 3 2 9 0 13 4 9 2
18 11 11 9 11 9 7 11 11 9 11 9 13 9 9 9 13 9 2
8 11 11 13 4 9 9 9 2
7 9 10 9 1 13 4 2
12 11 9 11 11 2 9 0 13 9 9 13 2
19 9 9 10 13 2 11 9 9 13 4 3 2 7 10 9 11 9 3 2
18 10 9 0 9 13 13 4 13 9 13 9 3 13 4 11 11 11 2
13 2 9 9 1 11 9 9 10 13 4 9 12 2
18 3 3 2 9 9 0 13 9 9 9 9 7 10 1 4 9 9 2
17 10 1 2 11 9 9 13 4 9 0 9 13 4 9 0 9 2
24 9 0 9 7 9 0 10 9 0 9 7 9 9 9 0 7 0 13 4 9 9 9 1 2
24 11 13 12 9 1 2 11 11 9 7 11 9 13 13 4 2 7 9 10 12 9 13 9 2
24 11 11 2 9 0 12 2 2 9 2 13 4 9 2 9 9 7 10 9 10 7 13 4 2
15 3 2 11 1 13 4 9 2 9 11 7 9 11 13 2
12 3 11 11 13 4 9 2 7 3 11 9 2
22 11 11 11 12 9 0 7 3 3 9 9 9 11 13 4 3 2 9 11 11 13 2
12 11 11 13 4 9 2 13 4 2 13 4 2
9 9 13 12 13 4 9 13 4 2
15 3 9 3 9 13 4 12 9 13 4 11 11 11 12 2
13 13 9 9 1 14 0 9 13 4 13 4 11 2
30 9 9 9 13 9 3 11 2 13 2 13 4 13 4 2 7 3 9 9 13 2 11 9 9 9 13 12 13 9 2
8 7 9 12 13 4 9 1 2
18 11 9 9 13 4 11 11 1 9 9 1 13 7 12 9 13 3 2
18 11 12 9 0 15 1 13 4 13 9 10 9 9 1 13 13 4 2
14 9 10 1 11 12 9 13 4 11 3 13 12 9 2
8 3 9 11 9 13 9 10 2
17 11 2 11 7 11 3 3 13 4 15 13 4 2 9 12 7 2
14 11 1 12 9 0 13 4 2 7 9 13 13 4 2
13 9 13 11 9 2 7 10 1 15 3 13 4 2
26 7 2 9 13 11 11 3 9 13 9 2 9 0 13 4 7 2 13 13 4 9 7 9 1 9 2
11 2 11 9 13 9 7 9 0 13 2 2
10 9 3 2 11 9 13 4 11 13 2
25 9 0 1 9 9 10 13 4 2 7 9 9 2 11 2 3 13 4 10 11 8 11 13 9 2
12 12 9 1 11 13 11 9 9 9 0 12 2
18 3 2 9 9 13 13 4 11 11 2 7 11 11 13 4 10 1 2
19 13 2 11 9 10 13 4 3 11 2 7 10 13 4 11 9 7 9 2
26 3 2 9 2 9 9 2 9 9 2 9 0 9 2 9 7 9 2 9 10 9 13 13 13 4 2
12 9 9 2 7 2 9 13 4 10 9 13 2
17 10 9 2 11 7 11 9 13 4 2 12 0 13 9 9 1 2
25 9 13 2 9 1 9 13 13 4 2 7 9 9 10 13 4 12 13 4 11 2 11 2 9 2
6 2 9 9 1 13 2
15 12 9 11 11 13 4 9 12 2 7 12 11 11 12 2
22 11 9 2 7 2 11 11 13 12 13 4 13 4 7 9 13 13 9 13 13 4 2
9 3 8 3 13 13 4 3 10 2
12 9 13 13 4 0 9 0 13 9 13 4 2
19 9 11 11 11 13 9 0 9 13 4 9 9 2 11 9 12 13 9 2
8 3 1 13 4 2 9 3 2
28 9 10 1 2 9 0 3 7 3 3 13 13 14 4 9 0 13 4 2 12 7 9 13 7 3 13 4 2
17 9 3 11 9 13 4 13 9 2 10 9 3 9 13 4 9 2
13 9 0 13 4 11 2 11 1 7 9 9 1 2
10 10 13 4 15 9 9 0 9 1 2
25 13 9 11 11 11 9 9 13 9 11 11 13 9 13 13 2 7 12 7 12 9 1 9 13 2
10 10 9 1 9 9 9 13 10 9 2
10 11 8 8 11 11 13 4 13 3 2
16 10 9 14 7 2 9 12 9 14 0 7 9 9 13 4 2
15 3 3 12 9 0 13 9 11 2 9 0 12 12 9 2
29 7 2 3 0 13 7 9 13 13 4 9 13 13 4 2 7 10 9 9 13 3 0 9 13 9 13 11 9 2
15 13 13 2 7 2 9 0 13 4 11 2 11 7 11 2
14 12 12 9 9 11 12 9 13 7 12 1 13 4 2
8 11 11 9 13 4 9 0 2
9 9 9 11 11 9 13 4 11 2
9 10 13 11 9 1 13 9 9 2
14 11 1 9 14 13 13 7 9 13 7 13 13 4 2
12 11 11 13 14 4 11 11 13 4 9 0 2
12 7 9 9 1 13 4 2 7 15 9 13 2
13 10 1 2 9 9 13 4 9 1 13 4 9 2
15 9 10 2 9 0 2 11 13 13 13 4 11 11 9 2
5 3 13 4 13 2
17 2 3 14 4 11 11 13 2 3 0 13 9 12 13 4 3 2
22 9 0 4 2 9 7 9 0 0 13 2 7 9 1 2 9 13 12 2 9 9 2
9 11 9 0 13 4 9 9 1 2
9 3 7 2 9 0 13 4 2 2
18 11 7 11 1 2 9 0 12 2 13 4 11 12 9 9 11 9 2
9 11 7 11 13 4 11 1 9 2
9 11 9 9 9 13 4 11 13 2
13 12 13 4 9 11 7 13 4 10 1 13 9 2
8 13 13 4 9 10 1 13 2
25 2 3 7 9 10 13 4 9 10 2 9 0 12 9 13 7 2 9 9 1 9 13 14 4 2
8 3 8 9 10 13 4 11 2
28 9 9 3 13 13 4 2 9 10 9 13 7 3 7 9 1 13 2 9 13 7 3 13 2 13 13 4 2
27 11 9 13 4 11 9 11 11 13 13 4 13 9 10 2 7 3 13 9 2 0 2 13 4 9 0 2
36 11 9 0 11 2 11 2 11 9 9 9 0 9 13 9 13 13 12 9 1 13 4 3 2 2 9 9 13 9 0 7 9 0 2 13 2
21 10 9 13 4 13 13 4 0 2 7 3 2 13 9 13 4 9 4 13 13 2
9 2 9 0 7 0 13 4 13 2
21 3 1 10 13 4 9 0 2 15 3 2 11 7 11 9 9 13 4 9 7 2
18 7 2 13 10 3 7 11 9 0 9 9 13 9 13 11 7 11 2
17 10 13 7 2 11 9 9 0 13 9 9 13 9 13 4 9 2
10 12 9 9 2 13 9 2 0 13 2
9 10 9 13 4 11 11 9 11 2
14 9 1 2 11 2 11 2 11 7 11 13 4 13 2
25 11 2 9 12 2 9 12 9 13 4 9 9 9 2 7 9 7 12 9 2 9 2 12 2 2
7 9 13 14 13 15 1 2
11 11 2 11 7 11 7 9 1 13 4 2
25 11 2 7 2 3 7 0 9 1 13 9 13 9 10 13 2 11 2 11 7 11 9 9 1 2
11 7 2 12 9 13 4 11 7 11 1 2
8 12 9 13 7 13 13 9 2
22 10 2 3 9 12 13 4 9 12 9 13 9 2 7 11 12 13 4 12 9 13 2
10 11 9 0 12 1 13 4 9 0 2
26 7 2 9 12 9 12 9 7 9 0 12 2 9 11 1 2 13 9 2 11 9 12 13 4 9 2
8 2 11 11 13 9 13 4 2
10 10 13 7 2 9 9 10 13 4 2
23 9 2 0 2 7 2 9 13 2 13 13 4 3 7 3 2 9 9 7 9 9 13 2
28 9 0 0 7 9 0 11 11 9 2 11 2 11 11 11 9 0 9 13 12 9 0 13 9 13 13 4 2
7 2 11 11 11 13 4 2
6 3 1 3 13 4 2
12 9 7 9 1 2 9 13 4 11 11 9 2
12 12 9 0 9 0 0 1 9 12 13 4 2
21 15 3 3 13 4 2 12 7 11 11 9 13 2 7 10 1 9 0 13 4 2
22 9 13 2 9 9 12 13 4 2 9 14 4 3 9 1 13 9 9 0 9 13 2
9 9 1 2 9 13 9 13 4 2
18 7 3 2 3 13 4 9 10 9 9 9 1 2 9 3 3 13 2
9 10 12 11 11 11 9 0 13 2
14 11 11 12 9 13 4 12 13 2 7 13 4 9 2
6 3 9 13 11 11 2
20 9 13 9 0 0 9 12 11 13 7 0 9 9 9 1 9 13 13 4 2
21 11 2 7 2 13 4 3 3 13 9 9 2 11 9 7 9 1 9 0 13 2
17 3 0 9 13 4 2 9 9 1 13 7 2 9 9 13 4 2
17 3 9 0 7 9 0 11 13 2 9 10 9 9 1 13 4 2
12 11 13 9 13 9 1 9 9 12 13 4 2
12 9 13 2 15 3 2 9 9 0 7 0 2
13 9 10 9 2 7 2 11 11 11 9 13 4 2
7 13 4 2 7 9 3 2
17 3 2 11 9 11 9 11 11 11 7 11 9 13 9 13 4 2
12 9 13 2 11 3 7 3 13 4 10 9 2
14 9 0 12 9 1 13 4 2 7 0 9 9 13 2
11 3 13 2 9 12 10 9 12 13 4 2
18 11 2 11 7 11 11 7 2 11 9 3 0 13 4 13 4 9 2
16 7 2 0 9 1 13 9 13 4 9 12 9 13 4 9 2
14 11 11 11 11 9 9 9 9 1 13 4 3 9 2
18 12 9 0 13 9 9 1 13 4 0 9 9 13 9 13 13 9 2
15 3 11 13 4 11 11 7 10 9 2 9 3 0 3 2
13 9 11 13 4 9 13 2 11 11 9 13 0 2
18 11 11 11 0 13 4 11 9 10 11 1 2 9 3 0 2 13 2
10 2 9 10 1 9 13 11 9 0 2
23 15 9 0 13 4 2 7 3 7 3 9 13 7 9 1 13 13 9 2 13 13 4 2
23 3 13 11 11 11 11 9 1 2 13 7 9 2 13 7 13 2 12 9 7 9 14 2
16 12 9 13 2 13 12 10 1 2 11 9 7 9 13 4 2
22 11 11 11 9 13 4 10 9 2 7 10 13 13 9 9 3 9 13 4 13 4 2
16 10 9 0 13 13 9 9 14 13 7 9 10 9 13 4 2
18 9 0 9 13 13 11 9 15 9 13 9 14 4 13 11 9 2 2
25 12 9 2 11 9 9 9 3 3 13 4 13 9 1 2 7 10 9 10 10 9 0 13 4 2
18 3 9 0 13 2 7 0 13 9 13 2 9 12 2 9 0 9 2
14 11 11 1 13 13 4 2 7 11 11 13 4 9 2
17 7 13 3 2 11 12 7 11 9 3 13 13 4 2 12 2 2
24 9 9 9 9 13 4 2 2 11 9 9 13 13 9 2 11 1 13 3 13 13 4 11 2
11 3 2 9 9 0 13 9 13 9 1 2
12 9 13 9 9 12 9 13 4 12 9 1 2
8 11 11 7 9 13 10 9 2
28 11 2 11 11 11 9 9 2 11 11 11 9 9 2 11 11 11 7 11 11 11 9 13 4 2 10 10 2
18 9 12 9 9 9 10 9 12 13 4 11 2 11 7 11 1 9 2
10 9 9 3 13 13 9 13 4 13 2
17 9 7 9 13 9 2 9 0 9 7 9 1 13 9 13 4 2
24 13 4 10 7 7 10 9 0 1 2 9 2 13 13 4 3 2 9 2 10 2 13 4 2
17 3 9 13 4 11 11 7 2 7 11 9 1 13 4 9 0 2
7 9 13 9 9 8 3 2
18 2 11 13 4 9 2 10 10 9 1 2 9 13 13 4 3 9 2
13 9 9 2 3 8 9 10 13 4 11 12 9 2
15 13 9 12 9 13 4 3 2 7 9 12 9 0 13 2
20 9 13 11 9 13 4 15 13 2 7 14 4 13 9 9 3 0 7 0 2
16 10 0 13 9 9 9 2 10 9 3 7 3 13 13 4 2
11 9 9 13 4 7 12 9 13 9 10 2
17 11 11 9 10 13 11 12 9 9 13 2 11 13 14 4 7 2
15 12 9 1 9 0 9 2 14 9 9 1 9 9 13 2
13 9 1 2 0 9 1 15 13 9 13 13 4 2
14 11 9 9 0 13 4 9 2 11 11 9 13 4 2
15 9 10 9 13 9 2 7 11 1 13 4 9 13 4 2
13 11 9 2 7 2 11 9 11 11 13 4 9 2
23 3 2 12 9 2 10 12 9 13 4 9 9 13 9 9 0 13 9 13 4 9 0 2
12 9 13 4 13 9 9 13 9 0 9 9 2
9 0 9 7 9 13 9 13 4 2
12 9 2 9 10 2 11 7 11 13 13 9 2
30 11 9 11 12 9 13 2 11 12 7 11 2 11 7 11 12 2 7 3 1 9 9 11 2 11 7 11 13 4 2
5 9 9 13 13 2
10 11 11 9 0 12 13 2 9 1 2
9 2 15 1 13 4 9 10 2 2
23 11 2 10 1 2 2 11 9 9 0 2 13 13 4 2 7 11 13 2 9 2 13 2
20 9 13 11 3 13 4 14 13 9 0 2 7 11 9 11 11 9 13 4 2
25 7 9 10 9 9 13 11 11 9 9 2 12 9 2 9 0 7 0 2 13 4 9 13 3 2
7 10 1 12 9 13 4 2
21 10 2 12 9 9 13 4 9 1 2 7 10 3 2 3 13 4 2 13 13 2
9 10 1 2 9 7 13 13 4 2
25 9 0 2 7 2 0 13 8 4 9 2 3 7 11 13 4 9 9 7 10 13 4 9 9 2
13 11 9 13 4 13 2 13 13 7 9 13 9 2
19 9 2 7 2 9 0 13 4 9 2 12 12 10 9 13 3 13 9 2
10 2 9 14 4 0 9 13 9 1 2
17 2 3 1 9 0 10 8 9 13 2 7 9 9 13 4 3 2
21 11 11 9 0 12 9 0 3 9 1 9 13 4 13 4 3 2 0 13 13 2
23 9 10 2 9 9 13 9 13 4 2 7 10 13 4 9 13 2 9 13 4 10 1 2
27 12 9 9 9 11 2 9 0 2 11 7 9 9 7 12 11 9 9 9 12 13 4 12 8 12 9 2
6 9 13 4 9 1 2
19 2 10 9 13 9 13 4 2 7 11 3 13 7 3 14 13 4 9 2
14 2 11 11 9 12 13 4 3 13 9 2 10 3 2
29 12 9 2 11 9 13 13 11 11 2 7 9 9 13 9 13 13 4 9 11 9 11 11 2 9 11 13 4 2
14 9 2 9 9 9 1 7 3 13 4 11 9 9 2
15 9 9 3 9 13 4 2 7 3 12 9 1 13 4 2
17 9 11 13 4 9 9 7 9 9 13 9 13 9 13 11 9 2
26 9 10 13 9 2 11 13 4 10 9 2 9 1 2 13 4 2 7 10 9 0 13 4 9 9 2
29 9 1 2 2 9 14 13 9 9 13 9 9 13 9 7 2 10 1 2 9 12 9 9 13 9 13 3 2 2
8 3 2 11 11 9 1 13 2
19 2 15 3 9 0 13 4 13 4 2 10 1 2 9 13 9 13 4 2
6 11 11 14 4 13 2
20 13 3 13 9 13 2 0 9 13 7 7 2 9 3 4 13 9 9 1 2
17 7 2 9 9 11 7 11 9 0 9 13 9 1 9 13 13 2
14 3 13 11 11 2 9 9 9 2 9 0 13 9 2
15 3 9 9 0 13 3 13 3 2 9 10 1 13 4 2
10 9 10 1 2 15 13 4 9 13 2
23 11 0 13 9 7 11 9 9 14 13 9 2 11 12 7 11 11 9 9 0 13 7 2
15 3 2 11 9 1 9 0 13 4 2 9 1 13 13 2
23 13 4 9 1 2 9 9 11 11 9 12 12 7 12 9 9 13 4 0 2 13 4 2
16 9 9 7 9 2 9 1 13 9 13 4 9 7 9 1 2
26 3 2 9 2 9 1 9 0 2 11 9 13 9 0 7 9 0 0 2 13 4 11 13 9 1 2
29 9 10 9 13 7 2 7 2 10 0 3 13 2 13 13 4 2 3 2 2 9 9 9 13 7 9 0 13 2
14 9 9 9 9 9 0 1 13 9 13 9 13 4 2
7 9 13 4 9 7 13 2
11 9 1 2 9 9 9 13 9 13 9 2
9 11 11 13 13 4 9 13 4 2
27 7 2 3 13 9 13 13 4 7 11 9 12 9 9 13 13 2 12 9 2 11 11 11 9 9 1 2
24 9 9 10 2 7 11 1 13 4 9 0 14 4 13 9 1 7 9 10 13 13 4 9 2
11 11 9 13 2 7 3 12 13 4 9 2
16 7 13 2 11 12 9 12 12 9 1 13 13 4 9 13 2
25 11 0 9 9 9 10 13 4 13 2 3 7 2 3 12 9 1 13 4 3 13 4 9 13 2
11 13 9 1 13 9 2 7 2 0 13 2
19 3 2 7 2 12 13 4 9 2 7 9 9 13 9 9 14 4 13 2
12 9 9 12 13 4 2 7 9 13 9 13 2
16 11 11 11 12 9 11 11 11 12 9 7 13 4 9 3 2
11 9 12 9 1 9 12 13 9 13 4 2
13 11 9 9 11 11 9 13 13 4 13 4 3 2
29 2 9 0 13 3 9 2 7 9 13 4 15 3 13 2 2 13 4 9 9 9 11 2 11 2 9 11 9 2
14 11 9 12 9 13 4 3 9 2 11 2 11 1 2
20 11 2 11 9 3 2 9 9 0 13 4 9 11 13 4 12 9 9 0 2
7 12 9 13 4 12 10 2
13 10 1 13 4 3 9 2 7 9 9 13 13 2
23 9 0 13 14 13 3 9 0 13 2 7 12 9 1 10 9 12 13 4 13 4 11 2
23 7 2 0 9 9 7 13 4 2 3 9 13 14 4 9 13 2 12 7 9 9 9 2
15 9 3 13 4 2 7 3 2 9 4 9 13 4 11 2
19 12 7 12 9 3 9 9 9 3 13 4 3 11 11 9 2 12 2 2
21 3 2 9 10 9 0 13 4 2 7 13 4 3 9 10 11 0 9 13 9 2
9 11 7 10 1 13 9 7 9 2
10 9 1 9 13 11 11 9 9 0 2
24 11 9 0 0 13 4 9 2 7 13 4 12 9 9 1 9 13 2 12 9 9 14 13 2
10 9 9 9 13 4 11 13 9 12 2
6 12 11 11 13 0 2
15 7 2 13 9 9 0 7 9 13 4 2 9 13 9 2
18 9 10 2 11 9 0 3 0 13 7 9 9 14 13 13 4 11 2
9 9 9 13 4 3 2 12 1 2
23 9 2 9 0 2 13 4 13 2 9 9 12 13 4 13 7 10 9 3 10 13 4 2
15 11 9 0 13 4 11 11 9 2 7 9 12 9 13 2
15 11 9 12 9 13 9 13 3 11 1 9 2 12 2 2
14 7 2 3 11 11 9 13 4 2 11 2 9 9 2
12 12 9 9 12 13 4 9 11 3 9 11 2
8 7 0 3 9 4 9 13 2
9 3 3 14 4 13 15 1 9 2
17 11 11 11 9 9 12 9 0 13 4 11 11 9 2 11 2 2
14 0 9 13 2 9 13 13 4 9 2 0 10 9 2
10 11 11 3 13 4 10 12 9 9 2
25 9 9 9 11 2 9 9 9 2 9 0 11 11 13 4 2 7 3 9 0 13 4 9 1 2
8 9 1 2 0 13 4 2 2
13 11 9 13 2 11 9 0 7 0 13 4 13 2
9 9 13 4 13 15 9 13 4 2
17 9 9 0 13 4 9 2 11 3 9 13 2 7 11 9 0 2
22 11 9 1 13 9 9 13 4 9 2 7 9 9 2 9 9 9 9 2 13 4 2
11 9 10 2 9 13 9 13 9 11 9 2
17 2 9 9 12 9 13 9 13 2 7 9 0 13 7 14 2 2
17 9 9 0 11 11 13 4 12 9 2 7 9 9 9 13 4 2
14 2 3 13 12 9 9 11 14 13 0 9 9 1 2
12 9 2 3 12 9 13 4 7 12 1 13 2
7 11 11 0 9 13 4 2
11 11 3 13 4 9 7 9 13 13 4 2
21 11 9 0 9 1 9 0 12 9 13 4 9 9 2 10 9 9 7 13 4 2
13 11 9 2 11 9 9 9 9 13 10 9 9 2
12 3 2 13 4 2 13 7 9 13 9 3 2
20 7 13 4 9 0 12 13 2 11 1 9 13 4 9 0 2 2 0 2 2
11 11 7 11 9 12 1 9 13 4 11 2
14 11 11 13 4 3 11 0 9 9 9 2 12 2 2
19 11 11 13 4 9 10 13 4 7 9 13 4 2 7 2 9 9 13 2
8 9 13 12 9 13 4 11 2
12 9 11 9 13 4 7 11 8 11 13 4 2
19 3 13 9 9 2 11 12 2 11 13 4 11 2 11 1 2 12 2 2
13 9 9 10 2 9 13 2 9 12 9 0 13 2
19 7 3 7 2 9 13 3 2 11 2 11 7 11 1 9 9 13 4 2
12 9 0 13 2 7 9 7 9 9 1 13 2
19 11 9 9 9 9 0 13 4 9 9 0 0 13 4 3 7 9 0 2
27 11 9 9 12 7 12 9 1 13 4 9 9 2 9 9 9 12 9 9 2 12 9 9 2 13 4 2
13 3 2 3 1 13 10 9 10 13 13 4 2 2
17 11 11 9 9 9 12 9 13 4 3 2 10 1 11 11 9 2
16 2 11 13 14 13 3 7 3 7 13 13 4 9 13 2 2
17 3 2 11 9 9 9 13 4 2 7 10 1 10 9 13 4 2
9 15 3 9 0 9 13 9 13 2
41 11 11 11 9 9 7 12 9 0 13 4 3 2 11 9 9 12 9 2 11 7 10 13 11 11 2 11 11 7 11 11 13 12 9 13 9 9 13 2 7 2
12 13 9 13 2 7 2 9 13 4 9 9 2
17 9 0 10 1 2 3 13 4 9 9 13 12 9 11 1 9 2
20 13 7 3 9 0 9 0 9 13 4 9 9 2 3 9 10 9 13 4 2
17 11 11 11 9 9 9 13 4 2 2 9 12 9 1 13 2 2
7 0 13 12 9 1 9 2
9 9 13 9 12 7 9 12 10 2
18 3 2 9 0 13 2 9 9 1 9 13 4 2 9 13 9 13 2
13 0 9 11 11 3 13 4 9 2 9 2 9 2
21 9 9 0 1 13 4 7 13 9 0 7 0 13 2 12 10 0 9 13 4 2
15 11 9 9 13 13 4 9 13 4 3 11 9 11 11 2
15 11 11 7 11 13 4 9 2 7 11 13 4 9 0 2
12 9 9 2 9 14 13 10 9 3 0 9 2
8 9 10 9 1 9 13 4 2
17 2 10 9 13 4 9 7 3 12 12 13 4 9 1 9 13 2
23 7 2 9 13 3 9 0 13 4 2 11 2 11 2 11 11 7 11 1 13 4 3 2
9 11 9 3 13 13 4 9 0 2
12 9 11 9 13 4 2 7 11 9 13 4 2
28 9 11 9 9 13 4 2 11 9 9 11 9 9 13 4 2 7 9 11 9 0 2 11 11 2 13 4 2
16 9 9 1 11 9 13 4 7 9 11 7 11 9 13 4 2
34 11 11 2 11 2 11 11 2 11 11 2 11 13 13 4 3 2 11 2 11 2 11 7 11 11 13 4 3 2 7 3 13 4 2
11 9 9 9 13 4 9 7 9 0 1 2
15 3 13 4 9 11 2 7 9 12 9 9 1 13 4 2
13 9 10 2 9 9 1 9 9 13 13 4 11 2
7 10 13 7 13 9 9 2
27 10 13 13 4 2 3 9 9 1 2 7 9 0 9 13 2 9 7 9 2 2 3 9 0 12 13 2
14 9 10 2 3 2 11 9 9 11 9 13 4 13 2
14 10 9 13 4 9 10 11 9 9 13 11 11 11 2
26 11 0 12 13 4 2 9 12 9 2 7 11 0 12 2 11 2 11 7 11 1 2 9 12 9 2
12 11 11 2 11 11 12 9 0 9 9 13 2
15 11 9 13 9 13 2 9 13 9 1 13 9 0 2 2
11 14 4 3 13 11 9 9 1 13 9 2
23 9 1 2 11 11 9 9 9 13 13 4 2 7 12 9 1 2 9 0 2 13 4 2
8 9 9 13 4 2 10 1 2
21 9 2 11 9 0 13 4 9 2 9 13 4 7 10 1 9 9 12 13 4 2
11 9 10 1 13 9 9 13 3 7 13 2
26 13 4 9 12 13 12 9 9 9 9 0 9 2 9 9 9 7 9 10 1 10 9 10 13 4 2
13 7 2 9 13 9 2 3 2 11 11 9 12 2
15 7 2 12 9 9 13 4 9 3 3 9 10 13 3 2
10 9 9 3 9 12 13 4 0 9 2
38 9 13 4 2 9 0 9 13 13 4 2 9 0 12 2 9 10 9 9 13 4 2 7 12 9 2 9 9 2 13 2 2 3 3 9 13 4 2
16 7 2 9 15 13 4 13 7 10 7 9 0 13 4 2 2
18 2 3 1 13 4 9 0 13 2 9 1 2 9 0 12 13 4 2
12 9 1 9 0 0 1 9 9 13 4 9 2
15 10 9 7 9 13 4 13 7 9 9 13 3 2 3 2
19 9 2 9 7 10 9 0 12 0 13 9 2 9 13 9 1 13 4 2
12 9 12 9 13 7 12 9 0 7 9 9 2
24 11 11 11 9 11 11 9 13 11 9 12 9 2 11 13 7 13 4 12 9 9 13 3 2
7 10 13 4 11 9 1 2
18 10 10 1 2 9 0 1 12 9 9 0 13 4 13 11 13 9 2
8 11 12 13 4 11 11 9 2
11 11 7 11 9 9 13 11 7 11 1 2
24 3 0 9 13 4 11 9 0 0 11 11 2 7 13 4 11 2 9 2 3 14 4 13 2
13 9 9 13 4 9 3 13 7 9 3 13 4 2
7 9 0 9 0 13 4 2
15 11 11 2 11 11 9 0 13 4 11 3 9 9 13 2
19 11 9 9 13 13 14 4 3 13 11 11 9 2 7 9 13 4 11 2
24 12 9 9 0 13 4 9 2 7 9 9 0 12 13 4 2 11 11 9 2 11 11 2 2
31 9 9 0 13 4 9 2 12 9 3 2 11 13 4 2 11 13 0 2 7 9 10 9 9 9 3 9 0 13 4 2
26 11 9 9 9 7 11 11 2 9 7 0 9 2 9 13 4 7 14 3 13 4 9 9 9 13 2
10 11 11 9 2 7 2 9 0 13 2
15 9 9 0 1 2 11 7 11 12 7 12 9 13 4 2
14 2 9 0 9 13 4 2 7 15 12 1 13 4 2
13 9 7 9 9 0 13 4 9 13 4 9 11 2
20 3 0 9 13 10 2 7 3 9 13 13 4 13 4 10 9 1 13 9 2
45 15 0 13 4 0 9 9 13 2 7 3 13 4 2 7 2 7 9 0 11 2 11 11 7 11 11 13 9 13 4 9 2 10 9 1 2 7 9 10 14 4 9 3 13 2
18 11 9 0 2 0 2 13 4 11 11 0 7 11 11 13 4 3 2
19 9 13 4 9 0 12 2 7 3 2 9 10 1 13 2 7 3 14 2
35 9 9 9 2 12 2 2 9 0 11 7 9 9 2 12 7 12 2 13 4 2 10 10 2 11 12 9 2 7 9 10 3 13 3 2
28 10 1 2 11 13 12 9 12 9 9 13 4 2 12 12 9 2 0 9 13 7 9 10 9 9 13 4 2
13 11 9 9 13 9 2 7 3 13 4 13 9 2
24 9 13 12 9 9 13 4 11 2 3 2 11 2 11 2 2 11 3 0 7 2 12 2 2
16 9 12 12 9 9 3 13 4 2 9 9 9 1 13 4 2
11 2 9 9 0 13 7 9 13 9 13 2
15 12 9 9 0 13 4 2 9 13 4 9 7 9 1 2
17 11 9 14 7 2 12 12 9 9 10 10 9 13 13 4 11 2
14 11 11 12 9 9 13 13 4 9 7 10 12 13 2
19 11 9 12 9 9 13 4 11 9 9 9 9 13 2 12 9 9 2 2
15 7 2 9 1 2 10 4 11 9 9 13 7 13 9 2
25 11 13 11 13 9 13 4 11 11 2 9 0 2 13 2 7 11 10 9 13 4 9 13 4 2
15 2 12 2 9 13 13 2 10 2 9 1 13 4 9 2
14 9 10 3 9 7 10 12 9 13 4 11 9 12 2
18 3 2 12 9 0 13 4 7 9 3 12 9 2 12 10 10 0 2
7 9 1 13 4 2 3 2
22 9 0 1 2 9 9 13 4 9 0 13 9 9 2 9 0 7 9 0 9 13 2
17 12 9 7 12 9 2 11 9 9 10 13 4 9 13 11 11 2
14 10 2 11 12 9 9 12 13 13 4 11 9 0 2
10 3 2 14 13 9 9 3 13 4 2
14 9 3 9 9 13 4 11 11 2 7 9 13 9 2
20 3 3 9 9 9 13 13 2 9 1 2 9 12 9 13 9 12 10 9 2
13 10 9 1 13 13 4 2 11 13 4 9 9 2
8 7 9 9 13 4 13 4 2
21 9 1 11 9 12 9 13 4 9 0 9 2 10 9 9 13 2 13 13 4 2
12 10 1 2 9 13 3 10 9 13 9 13 2
14 9 10 13 9 13 9 9 9 13 4 2 9 1 2
16 9 3 8 2 9 3 9 13 10 9 2 3 9 9 10 2
25 2 3 2 9 0 13 4 3 7 12 9 13 7 2 9 14 4 10 9 10 3 0 13 2 2
16 11 12 2 11 12 2 11 9 7 11 12 13 4 9 9 2
13 9 1 2 9 13 4 9 0 10 13 13 4 2
14 2 13 9 13 11 14 4 3 13 15 13 10 9 2
8 10 1 2 9 9 13 4 2
22 9 9 12 9 13 4 9 7 13 4 13 3 13 4 9 7 3 13 4 10 12 2
17 9 9 13 9 9 13 4 13 13 9 13 13 7 9 13 4 2
19 9 0 13 9 1 9 0 0 2 7 13 11 7 11 7 9 1 13 2
13 10 12 2 11 2 11 0 7 11 13 4 9 2
14 11 9 0 7 9 0 11 9 9 13 4 11 9 2
10 9 13 4 13 2 7 0 7 10 2
7 9 9 12 1 13 4 2
21 9 0 2 9 9 10 2 7 9 13 9 11 9 0 13 9 13 4 9 0 2
19 3 9 10 1 2 7 2 11 11 9 9 9 9 9 12 9 13 4 2
16 11 9 11 11 13 4 9 11 2 9 2 13 4 9 9 2
14 10 13 9 10 13 4 2 3 8 12 9 9 10 2
8 2 3 3 9 0 13 9 2
14 11 9 3 13 4 11 9 12 9 9 13 13 9 2
15 9 2 9 13 9 7 9 0 13 9 13 4 13 9 2
10 9 12 9 7 10 9 13 13 9 2
25 2 0 9 9 2 9 0 2 9 13 9 13 2 9 10 9 0 0 13 9 13 9 13 4 2
17 11 11 3 13 4 14 4 0 13 2 9 10 0 13 14 4 2
15 11 12 9 9 0 13 9 13 4 3 11 11 2 11 2
24 9 9 2 11 2 9 0 9 2 7 11 11 2 11 9 9 2 13 4 2 9 0 9 2
15 11 11 7 11 11 11 0 13 11 12 9 13 10 13 2
18 9 0 13 4 11 9 9 0 12 13 9 0 9 13 9 13 4 2
10 11 11 9 12 9 12 13 4 11 2
16 9 10 13 13 2 10 10 2 9 13 4 9 0 9 12 2
9 9 9 9 13 4 3 11 9 2
14 13 11 11 9 13 4 11 11 2 7 11 11 11 2
9 0 9 0 13 11 9 0 1 2
6 7 9 13 3 1 2
25 11 3 3 12 9 2 12 3 13 4 7 10 9 13 9 0 7 13 0 9 2 11 13 4 2
13 11 3 13 9 14 4 13 9 9 1 13 4 2
11 7 2 12 7 2 10 9 12 13 4 2
30 9 1 13 4 13 9 13 9 11 9 3 9 0 13 4 7 2 7 2 14 4 0 9 13 9 9 0 1 13 2
35 11 11 0 2 9 9 0 9 2 4 13 13 4 7 9 9 9 13 9 9 7 2 11 9 9 13 14 4 13 4 9 2 13 4 2
7 13 9 3 9 7 9 2
27 11 11 9 2 9 3 3 2 2 7 2 9 8 9 0 13 13 4 2 7 3 9 9 10 13 13 2
26 11 11 9 12 9 13 11 11 13 4 2 11 11 9 9 0 9 9 13 0 13 9 13 13 4 2
18 11 1 2 2 9 0 2 13 4 2 7 11 2 13 2 13 4 2
12 7 2 11 9 1 13 4 9 0 13 4 2
12 9 10 14 13 3 7 9 10 13 4 13 2
14 9 9 7 13 4 2 9 1 9 10 9 13 4 2
17 11 11 9 0 12 9 13 4 9 11 2 12 9 9 12 1 2
19 11 9 9 10 13 13 4 11 2 7 9 0 1 9 3 0 13 13 2
23 9 0 13 4 9 10 2 7 2 9 8 14 3 2 14 4 13 12 9 2 12 2 2
18 3 13 3 2 11 0 9 13 11 11 2 7 0 13 3 9 1 2
20 2 11 9 9 13 4 3 2 9 13 10 9 1 13 13 4 12 2 2 2
11 7 9 2 9 10 13 4 9 7 9 2
11 12 1 9 3 0 13 13 4 11 9 2
19 9 3 0 13 9 11 9 9 13 9 0 7 0 1 9 0 13 4 2
8 9 13 9 9 7 9 3 2
22 9 7 14 4 9 9 10 13 7 11 11 12 9 13 9 12 0 12 9 13 4 2
14 3 2 9 12 7 2 9 9 9 9 9 13 4 2
5 9 9 9 13 2
16 3 1 13 12 9 3 13 4 14 13 3 0 11 9 13 2
30 9 9 13 4 14 4 2 13 2 11 9 2 9 9 13 13 13 4 2 11 9 13 7 9 2 13 4 13 2 2
24 9 10 2 9 9 3 0 13 9 0 10 2 10 1 9 9 9 7 9 9 9 13 4 2
8 15 3 13 4 7 11 9 2
16 7 2 11 11 11 12 9 0 9 0 9 1 13 4 3 2
13 3 13 2 7 2 13 2 10 3 13 4 9 2
7 9 9 13 4 11 1 2
19 11 11 11 9 9 9 0 13 4 0 11 9 2 2 11 9 1 2 2
9 0 14 4 3 9 15 1 13 2
25 7 3 2 9 12 9 10 9 13 13 10 13 9 13 2 7 7 2 9 9 10 13 13 9 2
16 11 9 12 9 13 4 3 9 11 9 11 9 9 11 1 2
27 2 9 9 13 2 13 9 13 2 11 13 4 7 9 12 13 4 2 13 4 13 2 10 9 2 2 2
17 3 7 3 13 4 0 9 2 7 9 12 2 12 7 12 10 2
19 9 10 9 9 9 13 9 13 13 4 13 4 11 11 7 11 11 0 2
18 3 13 9 3 2 11 9 0 7 10 13 4 11 13 12 9 10 2
11 7 0 14 13 3 10 9 11 13 13 2
8 9 11 9 1 9 13 4 2
13 10 2 12 9 13 9 9 13 4 9 13 4 2
14 9 0 7 9 0 1 9 9 0 13 7 3 13 2
14 11 12 2 11 7 11 12 2 11 13 4 9 0 2
17 9 13 2 9 2 13 4 2 11 13 4 2 13 9 9 13 2
22 11 9 0 13 4 0 9 9 13 11 9 9 10 1 2 11 7 11 1 2 3 2
20 11 7 11 9 2 0 1 9 7 9 0 13 4 15 1 13 9 7 9 2
16 9 12 13 13 4 2 10 9 13 2 7 9 9 13 4 2
22 9 13 4 11 9 9 1 7 9 9 13 4 2 9 0 9 9 13 4 13 2 2
15 11 11 9 7 3 13 4 2 13 9 11 13 4 11 2
22 11 1 2 11 9 9 13 4 13 11 9 12 9 2 7 13 9 9 13 9 10 2
10 9 1 12 9 0 13 4 9 10 2
27 2 9 3 0 13 2 2 13 4 11 9 9 2 7 3 7 11 13 4 3 10 9 2 9 13 9 2
25 13 11 9 2 13 11 9 2 13 11 9 13 10 2 7 2 12 12 2 13 11 11 11 12 2
21 11 9 9 13 13 12 9 9 2 9 9 2 7 13 4 13 13 4 13 9 2
18 2 11 9 9 1 13 9 13 7 9 10 10 9 13 4 2 11 2
9 12 0 1 9 13 4 9 9 2
18 9 9 13 7 2 12 9 13 4 9 2 12 11 7 10 2 11 2
18 0 9 3 13 4 7 9 9 13 7 9 1 0 9 7 13 4 2
28 11 13 9 13 7 2 11 11 9 0 13 13 7 2 9 10 9 9 0 9 1 13 13 4 13 4 11 2
15 9 9 9 13 7 2 9 10 1 13 4 2 12 9 2
8 11 9 12 9 13 4 3 2
16 9 1 13 4 9 10 9 1 13 10 9 7 9 13 13 2
14 3 2 7 2 3 13 4 9 2 9 12 9 10 2
13 3 9 13 4 9 7 9 13 13 3 13 9 2
25 11 11 11 9 11 13 4 13 9 13 7 2 12 9 9 1 9 13 4 11 7 11 9 9 2
12 10 9 13 3 9 10 9 7 9 10 1 2
7 11 3 13 3 13 4 2
21 3 2 9 13 9 9 9 0 13 9 13 2 7 10 0 9 12 13 9 13 2
14 2 9 9 2 9 10 9 13 4 9 9 4 7 2
25 7 9 0 12 13 9 13 2 7 3 3 13 4 3 7 9 9 12 13 2 9 13 9 13 2
34 12 9 7 2 9 0 13 4 9 2 11 11 3 1 9 9 3 13 9 13 7 11 2 7 2 9 1 13 9 0 13 9 13 2
19 13 4 15 1 0 13 4 9 0 9 12 13 7 13 0 9 9 12 2
27 11 11 9 11 9 0 9 13 9 13 13 7 2 9 14 7 2 11 9 7 9 13 9 9 13 4 2
20 11 9 9 13 4 11 11 11 3 9 7 11 11 2 12 2 11 12 2 2
12 11 9 9 0 0 9 12 13 9 11 9 2
20 12 9 9 13 3 2 15 9 13 13 4 7 2 11 9 13 9 13 4 2
17 3 13 3 2 9 3 13 4 7 9 1 13 9 3 13 13 2
11 7 9 13 2 9 9 1 9 13 4 2
12 11 1 13 9 13 4 9 13 9 13 4 2
14 3 3 2 3 13 12 9 13 4 11 12 9 11 2
19 9 10 11 11 0 13 4 2 3 12 9 2 7 11 12 9 13 4 2
16 11 11 9 9 9 0 9 13 4 13 9 2 9 13 7 2
24 11 9 13 4 9 13 4 11 7 10 9 10 1 9 13 4 2 9 13 7 9 13 13 2
15 3 2 12 9 1 13 4 13 4 9 12 9 13 4 2
15 3 9 0 9 13 9 13 2 7 10 1 10 13 4 2
12 9 9 12 1 13 2 0 2 13 4 11 2
19 9 13 13 4 13 4 2 9 1 2 9 9 13 11 7 11 9 11 2
21 11 11 13 9 11 11 2 11 9 9 9 2 11 9 13 13 4 11 9 2 2
21 9 2 9 9 9 2 13 13 4 2 7 2 0 2 2 9 1 2 13 4 2
7 9 12 9 1 13 4 2
19 9 9 2 2 12 2 9 9 11 11 9 9 13 4 2 12 9 9 2
22 3 2 9 1 12 9 13 4 2 7 3 13 2 12 9 13 4 11 11 9 0 2
10 10 2 11 11 13 4 7 0 13 2
15 15 9 2 9 13 9 13 2 9 1 13 7 3 13 2
17 9 1 2 9 2 9 2 7 9 7 9 9 13 10 10 9 2
15 2 11 9 7 9 13 13 4 9 2 7 9 9 2 2
15 12 12 9 10 12 9 13 4 11 2 0 1 9 9 2
12 3 9 2 10 9 9 9 1 13 4 7 2
22 9 3 14 13 3 3 0 2 7 9 3 13 4 2 7 3 9 7 0 13 4 2
28 11 11 11 9 9 13 4 2 9 9 12 9 13 4 9 9 11 9 9 12 1 2 9 9 11 9 1 2
15 15 9 13 4 2 7 9 0 12 13 4 15 9 1 2
15 9 10 1 2 11 9 9 9 0 9 13 4 12 9 2
15 10 9 2 11 9 9 7 9 7 9 9 9 13 4 2
15 11 9 11 11 0 13 4 2 13 2 10 9 9 13 2
20 11 9 0 13 2 9 9 9 13 4 3 12 9 2 9 9 12 9 1 2
11 11 2 11 11 7 11 11 9 13 4 2
23 10 2 11 9 11 9 12 3 13 4 9 12 9 9 12 1 9 13 9 12 13 9 2
22 0 9 9 13 4 9 9 13 2 11 2 11 2 11 2 11 7 11 1 9 13 2
7 9 9 12 9 13 4 2
12 11 11 13 4 2 9 7 9 13 14 4 2
12 9 1 2 12 9 9 0 13 4 12 9 2
16 9 9 0 12 1 13 7 9 9 7 9 9 0 13 13 2
15 7 2 12 9 3 13 3 2 10 9 12 13 4 9 2
30 11 7 11 1 13 9 2 10 12 9 9 13 4 9 11 11 7 9 2 3 3 13 10 0 9 13 4 0 9 2
12 9 13 9 1 2 7 2 15 10 13 4 2
8 3 3 13 11 9 13 4 2
15 2 3 3 13 4 2 14 2 9 10 9 2 0 6 2
15 9 9 1 13 9 2 7 9 13 3 13 9 10 13 2
22 11 9 13 10 2 7 3 11 13 4 2 7 11 9 4 13 2 13 9 0 9 2
10 9 1 9 13 9 1 7 9 13 2
41 9 4 13 13 11 9 11 9 0 9 7 3 11 11 9 13 4 2 2 11 13 13 4 9 9 7 0 9 10 13 7 11 9 0 13 9 0 7 0 13 2
15 9 9 2 7 2 10 9 13 4 12 9 13 9 0 2
24 11 11 9 1 0 13 4 9 2 10 12 9 1 2 9 9 12 13 4 9 13 4 13 2
16 9 3 12 9 13 4 2 7 3 9 9 13 9 13 4 2
13 11 11 2 3 2 0 9 1 13 4 9 9 2
10 9 12 2 12 9 12 9 13 4 2
15 9 7 9 2 9 10 13 4 0 9 13 9 12 1 2
20 9 2 9 7 9 1 9 0 9 13 4 7 9 0 12 10 9 13 4 2
7 12 9 12 9 13 4 2
15 9 9 12 1 2 9 7 9 9 12 1 13 13 4 2
20 9 0 13 4 9 10 11 9 9 1 2 0 7 2 3 1 13 4 0 2
7 12 9 1 9 13 4 2
17 10 9 2 9 12 2 10 9 13 13 4 13 8 0 13 13 2
15 11 7 11 12 0 13 4 9 12 1 2 9 9 9 2
25 9 10 2 12 9 12 13 3 2 12 9 13 4 9 10 2 3 0 0 9 13 9 9 13 2
22 11 2 7 2 11 12 9 9 9 1 13 4 12 9 2 7 11 13 4 10 9 2
11 9 3 2 9 12 13 9 13 9 2 2
19 9 9 10 9 13 2 9 7 9 1 13 9 13 9 9 9 9 13 2
15 11 7 11 13 3 2 11 4 13 2 9 13 4 3 2
13 3 0 7 2 9 10 13 4 11 11 9 0 2
9 11 9 9 12 13 13 11 9 2
21 3 11 9 0 13 4 9 2 7 2 9 13 12 9 9 2 12 0 11 11 2
18 11 9 0 13 4 11 9 2 0 9 7 9 9 10 3 9 13 2
12 9 9 9 9 9 13 13 9 13 4 9 2
10 12 9 13 7 12 13 12 9 9 2
22 9 0 9 9 2 2 14 13 0 11 11 9 11 9 13 14 4 11 9 0 13 2
16 9 13 4 9 9 9 2 3 13 9 9 1 12 13 3 2
12 0 9 9 13 9 13 2 7 15 13 4 2
14 9 9 9 12 13 4 9 12 9 9 12 9 11 2
24 11 9 13 11 12 9 13 9 9 9 13 4 2 9 9 9 10 1 9 9 13 9 13 2
12 12 9 9 13 9 9 11 11 11 12 9 2
21 11 2 7 2 12 13 7 12 9 0 11 9 2 11 2 9 12 1 13 4 2
10 13 4 9 9 1 2 3 13 3 2
15 7 2 3 12 9 13 4 2 12 9 8 12 9 10 2
17 12 9 9 13 4 11 15 13 4 2 9 1 13 9 13 4 2
7 0 13 4 11 1 9 2
12 2 11 9 13 4 13 9 10 9 0 13 2
20 11 11 11 11 9 9 9 13 3 2 2 9 12 12 9 1 13 13 2 2
11 9 7 9 11 3 13 4 13 9 13 2
14 0 13 2 3 13 9 10 0 9 13 4 9 0 2
17 11 11 13 11 12 9 0 3 13 9 13 4 9 9 12 9 2
15 11 11 9 13 2 3 9 9 0 13 4 11 11 0 2
10 7 2 3 9 9 0 4 13 13 2
36 11 2 11 2 11 7 11 7 11 9 9 7 9 9 13 4 3 11 9 7 9 9 0 13 4 9 13 9 13 7 10 1 10 13 13 2
13 9 1 2 11 13 11 13 9 13 11 9 0 2
22 11 9 0 13 4 2 12 9 13 4 9 9 2 9 1 2 9 2 7 9 12 2
21 9 10 2 3 0 2 9 0 9 10 9 13 4 15 9 0 13 9 13 13 2
35 11 11 2 3 2 9 13 11 9 0 2 7 14 9 2 2 7 9 10 9 2 10 9 11 2 9 0 9 2 2 13 4 2 3 2
14 9 11 2 11 7 11 9 13 4 12 7 12 9 2
9 11 9 9 9 1 9 13 4 2
23 11 9 13 7 11 11 13 2 14 4 13 13 2 7 2 10 9 3 13 7 13 4 2
15 11 11 11 0 13 4 3 9 11 2 9 1 13 9 2
23 11 9 2 11 2 2 9 11 9 9 12 13 9 12 13 4 9 0 12 13 4 13 2
12 9 11 3 13 2 3 9 0 13 4 9 2
11 9 6 12 13 2 9 9 9 13 4 2
14 11 9 9 11 11 11 2 9 2 13 14 4 9 2
17 11 7 11 1 12 9 9 12 13 4 2 9 9 3 13 4 2
8 9 10 9 12 13 9 1 2
13 11 11 9 13 4 2 7 12 9 1 11 13 2
16 11 1 13 4 9 13 2 12 9 13 4 3 9 13 4 2
16 12 13 4 3 11 2 7 3 13 4 9 11 9 0 9 2
20 9 9 0 9 9 9 0 9 11 11 13 4 3 2 11 9 9 13 9 2
22 0 13 4 2 7 2 9 0 13 4 9 9 1 13 14 4 11 9 10 12 9 2
28 9 10 1 2 11 11 9 11 2 11 9 0 2 13 4 2 7 3 13 2 11 11 13 4 11 12 9 2
15 9 13 3 2 11 11 9 13 3 9 13 4 12 9 2
29 11 14 4 13 7 13 9 11 9 9 11 9 13 9 13 4 2 7 3 10 10 10 9 0 13 9 13 4 2
11 2 9 9 0 13 7 9 13 9 13 2
15 11 9 0 10 13 4 9 2 10 10 13 4 11 1 2
24 9 9 12 1 2 11 11 9 13 4 13 13 4 9 9 13 9 0 12 9 9 1 13 2
14 9 0 10 1 2 9 9 3 13 9 13 13 4 2
25 11 14 4 12 1 9 0 13 2 7 3 9 0 13 9 13 2 12 7 13 4 9 11 13 2
24 11 7 11 9 2 7 2 9 9 1 9 9 12 9 13 4 9 0 1 9 13 12 13 2
14 11 11 9 0 9 0 13 13 4 3 13 9 9 2
20 9 0 13 9 0 10 13 4 2 10 9 0 1 9 9 0 9 0 13 2
21 10 9 2 2 9 9 9 12 13 13 3 2 7 13 4 0 9 9 1 2 2
26 9 9 2 11 3 13 13 4 9 2 2 11 9 9 14 13 0 9 10 13 4 11 11 9 2 2
20 3 2 9 7 9 13 2 9 3 7 3 13 13 4 2 2 9 13 2 2
21 2 3 1 9 10 13 4 7 10 10 14 7 10 10 9 13 13 4 9 0 2
25 11 9 9 0 13 7 13 4 2 9 0 13 12 9 9 2 9 9 2 9 7 9 2 13 2
13 9 9 1 13 2 9 0 12 13 4 11 9 2
10 11 11 11 11 9 13 4 3 1 2
8 11 11 9 13 4 9 0 2
25 10 9 13 4 9 0 10 13 2 9 13 2 3 2 9 13 3 2 9 3 9 1 13 4 2
17 11 2 10 9 12 1 2 9 9 13 7 13 9 13 4 9 2
10 11 9 9 0 13 13 13 9 1 2
39 10 13 7 9 0 13 14 13 9 13 11 11 9 9 0 12 13 4 9 0 7 13 9 13 4 7 15 13 4 13 4 9 12 13 4 11 9 1 2
20 9 10 13 9 13 9 3 0 13 2 11 11 9 7 11 9 11 0 1 2
8 3 9 9 12 9 13 4 2
11 11 11 11 9 9 13 2 7 9 9 2
15 9 13 2 9 13 13 4 11 11 11 9 9 12 9 2
20 0 9 0 13 4 9 13 4 7 11 11 11 0 9 9 9 1 13 4 2
22 9 10 9 9 9 0 13 9 9 12 13 13 2 3 1 9 0 9 13 9 13 2
17 10 13 13 4 11 9 13 2 7 10 1 9 10 14 4 13 2
13 9 13 9 9 0 13 13 4 9 9 9 9 2
21 11 13 9 9 10 13 9 13 4 2 7 2 9 9 13 2 9 1 13 4 2
15 10 9 2 9 2 7 14 9 2 13 4 13 9 10 2
18 3 2 9 9 3 9 13 7 9 0 9 13 4 13 4 11 9 2
16 7 2 12 12 9 0 11 9 13 11 9 9 3 13 4 2
15 9 9 13 4 2 7 9 10 9 1 9 12 13 4 2
20 11 11 11 9 9 13 4 11 7 11 9 9 13 4 2 11 6 12 13 2
27 9 13 4 12 9 11 7 11 9 0 2 11 9 7 11 11 12 9 9 11 3 13 9 13 4 7 2
24 10 9 9 13 2 9 1 2 7 10 1 9 9 9 2 9 0 7 13 13 11 9 13 2
17 10 10 9 2 9 9 13 9 7 13 9 9 9 13 4 9 2
12 10 3 2 12 9 0 9 13 4 9 9 2
12 3 9 13 4 9 1 13 4 9 10 13 2
13 2 9 3 9 13 4 12 9 9 13 4 2 2
11 3 9 1 13 4 11 9 9 7 9 2
19 10 9 0 13 2 7 9 14 7 9 7 13 4 2 9 1 9 13 2
19 11 11 13 9 7 10 13 4 12 9 11 7 11 11 9 0 13 4 2
7 12 9 13 13 11 11 2
12 11 2 11 7 11 11 13 4 3 9 10 2
18 12 9 13 9 9 1 2 9 9 13 4 9 13 4 13 0 1 2
9 11 11 11 7 11 11 13 4 2
13 11 9 10 9 7 9 10 1 9 13 13 4 2
22 9 10 1 0 13 2 9 1 13 4 9 12 9 1 2 9 7 9 9 9 1 2
22 11 13 9 2 7 2 9 9 13 7 11 10 9 13 2 11 11 9 9 13 4 2
22 10 1 2 9 13 13 4 9 9 2 9 0 9 13 4 12 9 9 9 13 3 2
15 0 9 0 13 9 7 9 13 4 2 9 7 13 9 2
20 11 7 11 13 9 9 13 0 0 2 3 1 14 4 9 12 10 7 13 2
9 2 0 13 9 12 13 4 13 2
34 13 2 7 2 9 0 9 9 9 0 13 9 9 7 9 12 13 4 2 7 9 13 2 9 0 9 12 9 13 9 12 9 13 2
8 9 10 9 13 4 9 13 2
14 9 9 13 4 7 9 0 13 9 9 9 0 1 2
31 0 2 9 9 13 9 2 15 9 13 4 11 7 11 11 13 4 9 10 2 11 13 4 2 9 10 9 13 13 4 2
22 9 3 13 4 2 3 9 10 13 3 2 9 1 9 2 9 10 9 9 13 3 2
8 11 0 9 9 13 9 13 2
22 9 1 10 9 9 13 4 9 0 13 4 13 9 1 2 7 14 4 9 0 13 2
10 11 3 13 4 7 14 3 3 11 2
23 11 11 9 0 9 1 2 9 9 0 12 13 7 9 10 9 13 4 13 4 13 9 2
13 7 2 12 9 3 13 4 9 0 2 11 11 2
19 11 9 13 0 13 2 2 7 12 9 13 10 9 13 0 2 2 13 2
25 11 13 4 3 2 7 3 11 7 12 9 4 13 2 3 7 3 2 10 9 13 7 9 13 2
12 9 12 9 13 12 9 7 0 12 12 9 2
14 11 12 9 13 4 13 9 0 13 4 9 9 0 2
38 10 9 12 13 4 9 2 7 9 3 3 9 13 7 2 3 13 13 4 9 2 7 12 9 11 11 12 9 13 4 11 2 11 9 12 9 13 2
17 2 9 14 13 9 2 9 13 9 9 9 13 4 13 13 2 2
15 9 9 9 9 13 4 13 11 2 7 3 13 13 9 2
34 9 11 9 13 13 4 2 7 2 9 9 9 2 12 9 9 9 2 9 9 9 0 2 9 13 9 10 9 7 9 0 2 13 2
7 0 13 9 1 9 13 2
10 9 12 13 13 9 9 10 13 4 2
26 2 13 4 9 0 14 13 9 2 13 4 9 14 13 2 7 3 7 9 13 9 13 2 11 13 2
19 11 9 9 9 9 9 13 11 9 13 9 9 9 13 13 4 11 9 2
20 11 2 11 2 2 11 2 11 11 2 7 11 2 11 2 9 13 4 0 2
16 3 0 4 13 13 2 7 9 2 9 7 9 13 9 13 2
14 2 11 7 9 15 3 9 13 4 3 13 13 9 2
13 9 10 13 4 11 9 11 1 9 13 4 13 2
18 3 1 2 11 11 0 13 4 12 9 0 12 9 13 9 10 13 2
19 9 9 13 9 1 2 11 9 9 11 11 9 0 13 9 13 9 13 2
16 7 11 11 9 13 2 9 10 9 13 4 9 13 13 9 2
8 2 13 9 13 4 13 2 2
16 9 9 13 11 11 2 10 11 11 12 9 9 13 4 9 2
8 9 0 13 3 2 3 7 2
19 11 9 9 2 9 0 13 2 12 5 2 9 9 13 7 13 9 13 2
10 9 9 3 0 13 4 9 9 9 2
25 3 2 7 2 13 13 13 4 9 0 9 12 11 11 13 4 9 12 9 3 13 4 7 14 2
14 9 10 1 13 4 9 9 7 9 9 14 13 0 2
18 12 9 10 11 11 13 9 13 2 12 9 10 9 9 0 13 4 2
22 3 9 13 0 9 14 13 7 9 13 9 9 14 13 2 13 4 13 7 9 1 2
17 12 9 0 13 4 2 7 2 11 11 2 11 11 7 11 11 2
