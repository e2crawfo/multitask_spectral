76 11
20 1 9 9 9 15 4 13 12 1 9 0 2 1 15 12 0 7 12 0 2
25 3 10 9 0 0 15 4 13 1 9 0 14 13 9 1 9 13 7 11 7 14 15 13 9 2
14 9 4 13 14 13 1 9 1 9 2 9 2 9 2
14 7 14 15 13 1 10 11 11 14 15 13 10 9 2
14 4 13 1 9 3 10 9 1 9 0 10 9 9 2
25 1 10 9 2 15 3 13 1 9 11 9 2 9 7 9 1 9 0 1 9 13 1 9 0 2
22 9 1 9 2 9 0 2 9 2 2 9 11 2 9 2 4 4 13 1 9 0 2
23 12 9 1 11 11 2 9 9 7 9 9 2 13 1 15 2 4 4 13 1 9 12 2
23 9 13 10 9 2 16 13 14 13 10 2 9 0 2 2 9 2 1 9 0 10 9 2
24 10 12 9 2 11 9 2 9 10 11 2 9 2 2 4 13 9 1 9 10 11 2 11 2
26 11 15 13 9 1 12 9 7 12 9 2 9 1 15 4 13 14 13 2 10 9 7 10 9 2 2
19 9 9 15 13 2 15 13 3 3 9 2 3 7 1 9 1 9 0 2
18 11 13 1 9 9 9 1 10 9 7 13 9 1 9 13 1 9 2
27 12 12 7 12 7 12 9 4 4 13 1 9 2 12 11 2 12 11 5 5 11 7 12 11 9 2 2
13 11 13 7 14 13 2 7 14 13 9 9 0 2
30 9 0 1 3 14 13 3 1 9 9 0 0 1 9 2 3 1 9 9 0 10 9 2 11 2 0 3 1 9 2
20 9 1 9 13 1 12 9 12 3 2 7 15 9 13 13 1 9 3 0 2
27 15 13 14 13 16 14 13 13 11 1 0 9 2 16 15 9 15 2 3 7 9 9 13 9 0 0 2
24 2 12 2 9 1 9 4 13 1 15 1 9 9 0 15 15 4 13 7 15 15 13 0 2
29 9 13 2 3 2 9 1 9 10 10 10 9 1 11 0 1 9 7 9 2 15 15 13 9 1 9 9 10 2
23 12 2 11 10 11 15 13 13 1 9 0 0 1 9 11 2 9 2 13 1 9 12 2
27 15 13 2 9 11 5 12 8 2 12 2 13 1 9 1 12 9 12 1 9 0 1 9 0 7 9 2
19 2 9 15 13 9 1 9 2 9 1 12 11 5 9 2 1 9 0 2
23 15 13 9 9 0 2 11 2 11 2 0 2 2 1 9 1 15 4 13 1 15 0 2
18 7 15 4 13 7 1 10 12 2 13 1 11 11 2 1 9 15 2
15 1 15 7 13 9 14 15 13 1 9 2 13 1 9 2
29 3 13 16 4 13 1 9 7 16 15 4 13 7 16 15 4 13 9 1 15 15 15 13 15 2 9 7 9 2
20 3 13 9 7 15 1 15 2 15 1 9 0 2 4 13 3 10 9 0 2
12 7 13 2 13 2 7 14 3 13 1 9 2
16 4 4 13 3 3 1 9 9 10 2 2 9 1 9 2 2
15 15 4 13 1 9 7 14 4 13 13 14 14 15 13 2
14 9 2 9 2 3 13 15 1 9 3 13 1 9 2
12 16 9 16 4 13 3 1 15 15 4 13 2
13 15 13 2 9 13 2 15 14 2 3 9 0 2
8 3 14 13 15 15 13 9 2
17 3 9 14 3 13 1 0 2 15 9 3 3 13 9 1 9 2
8 10 9 14 3 13 1 9 2
14 9 9 14 3 13 1 9 3 13 1 9 10 0 2
13 15 15 13 16 10 9 14 3 13 1 9 0 2
14 15 13 3 13 14 13 3 3 9 7 3 3 9 2
9 13 3 15 13 1 9 1 9 2
8 13 2 13 3 15 13 9 2
10 15 13 3 13 1 9 7 1 9 2
16 7 2 15 13 2 1 9 11 14 13 3 4 13 15 13 2
10 4 13 14 13 1 9 3 4 13 2
6 15 4 13 13 3 2
15 15 2 3 9 1 10 9 2 13 14 15 13 1 9 2
7 13 13 1 9 1 9 2
11 15 13 14 13 3 0 7 3 0 9 2
14 15 13 13 2 3 3 1 9 2 9 10 9 0 2
6 3 13 13 3 13 2
14 1 9 10 2 13 15 11 13 7 14 13 1 9 2
42 1 9 1 12 9 12 2 9 0 13 3 1 11 1 9 3 1 9 9 2 9 11 15 13 9 1 9 1 9 10 9 11 16 15 4 13 9 9 1 9 0 2
23 10 9 0 0 1 0 9 0 4 13 9 9 2 3 11 11 4 13 9 0 10 9 2
17 0 9 4 13 15 1 9 0 7 4 13 10 1 9 9 0 2
14 1 3 12 15 4 13 9 10 9 1 9 7 9 2
19 11 4 4 13 9 2 3 9 10 2 9 9 0 2 4 13 9 0 2
7 11 11 4 13 12 9 2
9 9 7 14 4 13 9 9 0 2
12 9 9 4 13 1 9 9 11 1 9 12 2
25 1 9 2 0 9 1 9 2 11 11 15 4 13 10 11 3 12 9 15 4 13 10 0 9 2
33 11 11 1 9 0 9 0 0 2 9 2 15 4 13 1 12 1 9 11 2 1 10 10 12 9 7 15 4 13 1 9 9 2
8 11 11 4 4 13 12 9 2
9 11 13 1 10 9 1 9 0 2
11 9 0 4 13 1 10 9 10 10 9 2
12 3 2 1 9 9 7 9 13 0 0 9 2
33 15 1 9 0 1 9 13 1 9 11 13 9 0 2 9 0 2 9 2 9 1 9 0 7 9 0 2 7 3 9 1 9 2
13 10 9 13 9 10 9 0 0 1 9 1 9 2
32 1 9 0 7 15 0 10 9 0 2 9 0 15 13 1 12 9 9 2 12 9 9 1 9 2 12 9 9 1 9 2 2
13 9 9 13 10 9 0 1 9 9 7 9 0 2
44 1 9 2 9 11 13 15 1 9 0 2 1 12 9 7 4 13 1 9 10 9 0 1 9 2 0 1 9 2 0 1 9 7 9 2 13 15 3 9 9 9 2 0 2
29 1 12 13 9 10 9 10 9 1 9 0 2 13 3 0 9 0 1 9 0 10 9 0 2 9 2 0 2 3
26 1 9 1 12 2 11 13 10 9 1 12 12 12 1 9 7 1 9 1 12 4 4 13 12 12 2
10 9 0 0 13 0 9 0 1 11 2
17 15 13 10 9 0 15 15 13 1 9 1 10 9 13 9 0 2
30 9 13 9 9 0 13 1 9 9 2 10 9 0 2 1 9 0 2 0 7 13 1 9 9 0 1 9 9 0 2
