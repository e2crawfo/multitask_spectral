5077 17
20 13 3 9 15 1 9 7 13 3 13 15 1 9 15 7 3 13 13 9 15
28 13 13 15 1 9 15 3 16 13 1 9 1 15 16 3 13 15 9 7 9 15 13 9 7 1 9 13 15
3 6 13 15
7 3 13 3 16 13 0 9
5 13 16 13 13 0
3 3 9 13
20 15 3 13 15 16 0 15 13 1 9 1 9 3 9 13 1 15 1 9 15
13 16 3 9 15 0 13 15 13 15 7 13 1 15
17 0 3 15 13 16 13 12 9 15 7 3 15 9 15 13 1 9
3 13 3 13
10 15 3 13 9 15 3 13 15 9 0
22 15 3 13 15 16 0 13 9 15 1 9 0 13 15 9 13 7 15 9 13 9 13
6 3 13 16 13 13 0
5 3 1 9 13 15
5 13 3 9 9 15
14 7 9 15 13 15 16 3 13 9 12 0 7 0 13
6 0 3 0 1 9 13
4 13 16 13 13
7 9 1 9 7 9 1 9
8 15 3 13 15 3 13 15 0
12 7 16 15 15 13 1 0 9 13 15 3 0
15 7 13 9 13 1 15 7 9 15 13 13 15 3 9 15
11 13 1 15 13 7 13 1 15 13 3 13
4 13 16 13 13
4 15 3 13 15
3 13 9 15
3 13 13 15
4 0 13 13 15
33 7 13 1 13 15 9 7 13 15 16 13 9 9 15 15 13 1 9 16 9 15 13 1 0 7 0 7 13 1 0 7 1 0
6 3 3 9 3 0 13
9 7 16 13 9 15 3 15 0 13
6 3 3 9 3 3 13
11 13 9 15 3 13 1 9 16 13 13 15
14 16 3 3 3 9 3 13 1 9 15 15 13 1 9
21 3 3 13 9 3 13 1 15 3 9 13 1 9 7 1 9 16 13 15 1 9
3 6 13 15
28 15 3 13 9 3 3 13 9 15 15 13 9 15 16 13 9 15 1 9 7 9 15 13 1 9 13 15 3
9 7 3 13 15 3 13 3 3 9
17 3 13 1 9 7 1 9 7 1 9 13 13 15 16 13 15 9
7 6 13 15 16 13 9 15
15 13 15 9 15 1 9 7 9 15 13 1 9 13 15 3
9 13 3 15 3 0 13 3 3 9
10 13 3 15 16 1 0 9 15 13 13
9 13 3 9 15 15 13 1 9 15
5 3 3 13 15 15
11 9 15 15 13 1 9 3 13 15 9 15
4 3 13 9 15
10 3 13 9 15 3 1 9 3 1 9
11 7 13 15 9 15 3 3 15 13 9 15
22 7 3 13 15 1 9 7 13 15 1 9 16 15 13 9 7 9 7 9 1 9 6
13 16 3 3 13 9 9 15 3 9 15 13 9 15
9 3 3 13 15 3 13 3 3 9
10 13 3 9 15 16 13 15 13 9 13
7 6 13 15 16 13 9 15
25 15 3 13 15 13 9 15 7 9 15 13 16 3 13 15 9 13 15 7 9 15 15 13 1 9
9 7 9 15 13 1 9 13 15 3
17 13 3 15 9 9 3 7 9 7 9 13 3 9 3 13 7 13
4 9 9 13 9
11 16 3 13 9 15 0 15 9 15 0 13
11 16 3 9 15 0 13 15 9 15 0 13
11 16 3 9 15 1 15 9 13 3 9 3
6 15 9 13 12 9 13
16 7 3 12 13 7 0 13 7 12 13 15 7 1 0 13 13
6 3 13 9 13 7 9
9 3 9 3 0 13 9 7 9 9
19 13 1 9 0 16 3 13 7 13 7 13 1 9 7 9 15 0 13 15
7 3 15 3 3 15 0 13
12 15 3 1 15 13 15 13 13 9 15 9 12
6 7 1 9 15 15 13
5 13 9 0 3 13
5 3 13 15 7 13
16 13 3 15 16 3 11 1 15 9 15 13 15 3 12 1 0
5 3 13 15 3 13
5 15 13 7 15 13
4 7 15 13 15
5 15 3 0 9 13
9 13 3 9 15 0 16 13 0 15
14 13 3 3 9 0 7 9 15 7 0 15 13 15 15
6 3 13 15 3 1 0
6 0 3 9 15 13 15
14 15 3 9 13 13 15 7 1 15 9 13 13 15 15
22 15 3 13 9 1 9 9 15 7 9 15 13 1 9 15 3 13 7 3 13 9 15
7 13 7 13 9 1 9 15
6 7 6 9 1 9 15
16 9 13 3 9 1 9 15 7 3 13 13 9 1 9 9 15
21 3 13 0 9 7 13 9 15 1 9 16 3 13 15 9 15 7 13 15 13 15
5 13 7 13 15 15
5 13 7 13 15 15
16 3 15 13 1 15 9 15 16 13 9 15 9 3 9 13 15
8 7 16 9 13 3 9 13 15
23 16 3 15 0 13 13 9 0 13 9 15 3 3 9 15 15 13 1 9 13 0 13 15
14 15 3 15 3 13 16 13 15 9 3 3 15 13 15
6 0 3 13 9 7 9
3 13 0 9
5 7 0 13 13 15
9 3 0 9 7 0 9 13 1 9
11 13 1 0 9 15 13 1 15 1 9 0
5 3 3 13 9 9
5 1 9 15 13 15
9 3 13 1 9 9 7 1 9 9
13 3 0 9 0 9 0 13 7 0 9 9 0 13
12 0 9 15 3 13 9 0 13 7 1 9 13
8 0 3 3 1 9 15 13 15
19 3 0 13 15 9 9 13 1 9 0 7 13 9 9 15 15 13 1 9
19 9 9 3 1 15 3 9 13 7 15 9 9 13 7 15 9 9 0 13
5 7 3 13 15 16
3 3 13 15
5 13 1 15 13 9
14 7 13 9 7 13 9 7 13 9 7 13 1 9 0
4 7 3 13 15
5 13 3 13 1 9
20 7 0 13 9 15 0 7 3 13 15 13 15 9 0 15 13 15 9 1 9
9 7 13 15 7 13 9 15 0 3
14 7 13 3 13 11 15 9 0 13 15 9 1 9 15
13 13 3 13 3 9 13 7 3 3 9 15 7 9
8 7 6 0 13 13 15 15 13
6 9 16 13 13 15 13
7 7 13 9 11 13 15 13
1 13
2 13 15
4 7 13 15 11
1 13
13 13 3 15 11 1 11 13 1 15 9 13 15 13
10 9 9 15 13 1 9 13 3 3 13
4 7 13 15 11
4 15 13 13 15
5 7 13 9 13 15
8 9 13 0 16 1 9 15 13
10 3 15 9 13 1 9 13 1 15 9
5 7 0 13 7 13
7 7 9 15 13 0 7 13
11 13 3 11 13 15 15 7 13 13 1 15
3 6 13 15
7 3 1 11 0 9 3 13
21 13 3 15 16 0 1 9 7 9 13 7 13 1 11 7 11 7 11 1 9 0
8 7 9 9 13 13 1 9 0
1 13
4 3 13 13 15
7 7 13 9 15 1 0 9
13 7 13 15 9 1 9 15 1 0 9 13 15 0
12 7 13 11 1 9 0 13 9 15 13 9 13
5 7 13 15 9 15
4 7 13 15 9
5 7 13 7 13 15
7 0 9 15 13 7 9 13
7 13 3 11 0 9 1 15
5 13 13 1 0 9
6 7 13 15 9 13 15
7 9 13 1 15 3 3 13
3 13 15 11
15 9 9 13 7 9 0 9 7 9 0 3 13 3 9 13
6 0 3 1 9 13 15
9 13 1 15 7 13 0 13 15 9
10 7 13 15 1 9 1 15 13 9 15
12 7 6 9 0 13 1 9 16 13 15 9 9
3 7 0 13
7 7 13 9 15 13 15 13
3 9 13 15
1 13
4 15 0 13 0
5 9 3 13 15 13
9 15 0 13 16 9 7 9 13 15
26 7 13 15 11 1 0 9 1 9 0 13 15 12 0 1 9 13 3 3 16 3 13 15 13 9 0
4 7 6 13 13
8 15 13 15 7 15 11 9 0
7 13 13 3 1 9 13 15
5 9 3 13 15 13
9 16 13 15 13 15 13 1 9 0
1 13
6 0 3 13 13 1 9
14 7 3 13 15 9 15 1 9 1 9 7 13 1 9
12 7 13 13 7 13 1 9 13 15 3 1 0
17 7 6 15 9 13 1 11 7 13 15 13 16 13 13 1 9 15
9 7 6 13 15 13 9 1 9 13
7 7 13 11 9 15 13 13
1 13
8 7 6 15 1 9 13 1 15
2 0 13
6 7 13 11 9 15 13
7 3 15 13 0 1 9 15
2 13 13
12 7 16 13 16 9 13 9 0 1 9 13 9
3 3 13 13
9 13 13 9 15 7 13 1 9 15
14 7 13 11 3 13 9 1 9 13 9 11 7 13 15
3 1 15 13
5 7 13 1 15 13
6 7 13 9 13 9 15
9 1 15 1 9 7 9 9 15 13
5 11 3 13 13 15
6 3 13 0 9 7 13
6 13 3 13 15 15 13
9 3 13 3 9 13 7 9 1 9
7 3 13 1 15 9 0 13
3 13 15 11
11 3 13 9 0 13 15 16 1 15 13 9
13 13 3 9 3 13 15 1 15 9 7 3 13 15
10 15 3 3 13 9 9 3 13 9 0
10 13 3 9 15 1 9 7 0 9 13
7 7 13 9 0 1 9 0
11 7 9 0 1 9 0 13 7 12 13 15
14 9 15 3 13 7 13 3 13 1 15 9 15 7 13
9 7 13 11 1 15 13 7 9 15
17 7 6 9 0 12 1 12 9 13 13 1 3 13 15 9 9 15
4 13 3 1 15
8 16 3 13 15 9 15 13 13
8 11 3 13 15 7 13 15 13
1 13
14 7 13 11 1 9 0 7 13 9 7 9 13 13 15
1 13
6 3 13 3 9 7 13
4 7 13 15 15
13 3 3 13 13 9 13 13 15 1 9 7 13 9
8 7 13 9 0 1 15 9 0
12 7 13 3 11 1 15 13 12 9 13 7 13
4 13 15 9 0
6 13 3 16 13 0 13
4 13 15 6 9
6 3 13 15 1 9 13
5 1 9 15 13 15
5 7 13 15 15 9
5 7 13 15 11 13
5 13 16 15 3 13
9 0 3 13 13 15 1 15 9 0
5 7 13 15 9 13
6 3 13 15 3 1 11
3 7 9 13
5 1 9 9 13 9
24 7 13 11 9 15 7 9 13 1 9 15 7 13 9 9 7 13 0 9 7 0 9 1 9
17 13 3 9 11 13 1 15 16 13 13 7 13 3 9 3 13 9
4 3 13 9 15
11 13 15 3 9 9 16 13 9 1 9 15
16 13 15 9 1 9 0 16 13 15 7 13 0 9 7 0 9
8 12 3 1 12 9 9 13 0
30 0 11 15 13 15 11 7 11 9 15 11 7 11 11 7 11 9 11 0 7 11 13 11 11 9 11 0 15 15 13
9 0 12 1 12 13 11 13 15 13
11 1 9 9 3 13 7 1 9 9 3 13
8 13 3 3 1 9 13 9 0
2 13 13
2 0 13
2 9 13
2 3 13
2 3 13
21 3 13 9 7 9 7 9 1 9 15 7 9 1 9 7 12 9 7 9 7 9
6 0 3 13 9 9 15
5 7 3 13 16 13
6 13 3 1 9 13 15
11 7 16 3 13 9 0 13 9 15 1 15
22 7 15 3 3 13 15 7 13 9 15 13 1 9 7 1 9 0 13 9 1 9 15
3 6 13 15
11 3 13 9 0 0 1 9 0 3 9 0
9 6 15 13 15 3 9 1 9 9
11 13 3 15 1 9 7 1 9 15 13 15
15 7 1 9 3 7 9 13 13 15 1 1 9 15 7 9
11 3 3 13 15 3 13 15 3 7 15 13
9 13 3 15 15 1 0 9 15 13
17 13 3 9 9 1 9 7 9 9 7 13 9 1 9 7 13 15
7 7 13 13 15 9 15 1
7 13 3 1 9 0 13 13
14 6 3 13 15 16 3 13 13 9 0 16 13 9 0
9 13 9 1 9 7 9 1 9 15
12 13 9 16 13 3 9 15 7 9 3 9 15
10 7 16 9 9 11 13 3 3 0 15
5 3 13 15 3 15
8 15 13 15 1 9 13 1 9
8 7 15 1 9 13 13 1 9
12 13 3 15 3 13 7 9 7 9 13 1 9
8 3 12 3 9 1 9 13 13
13 7 3 15 3 1 15 3 13 1 9 1 9 15
8 15 3 3 9 9 15 13 13
4 3 13 15 3
5 0 9 0 15 13
17 15 13 15 15 1 9 13 15 15 3 15 1 9 15 13 1 9
6 3 13 13 9 7 9
17 13 3 13 9 1 9 15 7 9 1 9 15 7 9 1 9 15
5 7 9 9 0 15
35 15 13 9 7 9 3 15 13 15 0 7 15 13 9 7 9 3 15 13 15 0 7 15 3 13 9 15 7 1 9 15 13 13 15 0
14 13 9 15 13 15 7 15 13 9 15 15 1 13 15
12 15 15 13 15 13 7 15 13 15 13 13 15
17 13 9 1 9 0 9 0 13 7 13 9 1 9 0 9 0 13
8 13 3 13 7 13 1 9 15
12 11 3 13 1 9 9 0 13 9 15 13 15
7 15 3 13 13 7 15 13
5 7 13 11 13 15
3 13 13 11
16 0 13 7 0 13 0 13 15 7 0 13 0 13 7 0 13
9 7 0 13 15 3 13 15 1 15
9 0 3 13 13 11 13 9 1 11
4 9 3 9 13
4 7 15 13 13
6 9 3 1 0 9 13
8 6 15 0 13 1 9 0 13
4 7 15 13 13
2 9 3
2 13 15
3 7 0 9
3 6 13 15
8 3 13 1 13 9 0 11 9
8 0 3 1 9 0 0 13 15
14 1 9 3 11 9 3 9 0 13 15 7 9 13 15
17 15 3 9 7 9 1 11 13 7 16 13 13 0 13 11 13 13
5 13 9 13 3 13
4 15 13 9 0
5 13 15 7 3 13
9 13 3 11 3 13 7 13 7 13
2 9 13
8 13 9 0 13 7 13 7 13
10 6 0 9 9 7 9 9 9 7 9
7 7 13 15 9 1 9 15
14 3 13 13 9 1 15 13 0 9 15 16 3 13 15
21 3 16 1 11 7 11 13 9 13 13 1 15 3 3 1 9 7 9 13 15 13
3 3 13 15
10 7 15 11 13 15 1 9 1 9 13
14 3 16 1 11 13 9 13 1 15 13 13 1 0 9
13 3 13 15 16 9 0 3 13 1 9 0 3 15
6 1 0 9 13 11 13
21 13 15 15 9 9 9 7 9 16 13 13 0 1 0 7 0 7 13 15 13 9
24 15 15 13 13 9 15 7 15 3 13 9 3 9 7 9 15 13 3 9 7 15 13 9 13
8 13 1 15 15 13 15 7 13
4 7 15 13 15
9 9 3 15 0 7 9 15 0 13
7 1 0 9 13 11 1 9
11 9 3 15 13 15 7 13 13 9 7 13
5 9 3 13 13 15
4 0 3 13 15
13 13 3 13 15 13 11 3 13 0 7 13 1 15
22 3 13 1 9 0 7 9 9 13 15 3 0 15 13 13 7 13 1 15 3 9 12
16 7 13 13 1 9 16 1 9 9 1 9 9 13 7 0 13
16 16 3 13 13 15 13 9 13 7 3 9 3 3 13 13 0
6 9 3 13 9 9 0
8 7 13 3 11 13 1 9 15
13 7 13 15 13 16 13 1 9 13 16 1 15 13
4 0 3 13 15
21 15 13 1 15 9 15 13 9 12 7 16 13 15 1 9 1 9 3 13 3 15
6 3 3 0 13 9 9
7 0 3 13 1 9 0 13
2 13 9
2 7 13
10 9 3 13 9 13 1 15 3 15 13
5 11 3 13 13 3
10 7 1 15 13 9 0 7 13 15 15
8 7 13 15 16 3 3 15 13
7 16 13 15 13 9 11 13
12 6 9 15 15 13 13 15 1 15 13 9 15
11 3 13 7 13 3 13 15 1 9 9 15
6 7 1 9 15 9 13
19 3 13 1 15 13 15 0 7 0 7 13 15 16 0 7 0 13 7 13
6 7 13 15 15 9 13
5 3 0 13 9 0
4 9 3 13 13
9 0 3 13 9 3 1 11 9 9
6 13 3 9 15 13 15
5 3 3 13 9 15
12 7 16 15 1 11 13 9 9 15 1 15 13
6 0 1 0 15 13 9
14 16 3 1 9 0 15 13 9 3 13 1 15 9 0
22 7 3 13 15 13 1 9 0 7 9 15 13 16 3 3 13 0 7 3 9 15 13
14 15 13 1 15 1 15 13 7 15 3 13 1 15 13
4 0 1 13 15
16 0 9 7 9 13 15 9 7 15 1 9 9 3 13 15 9
17 7 15 13 1 9 0 3 13 15 15 7 1 0 9 7 1 13
16 7 13 9 0 7 9 15 0 7 13 9 0 7 9 15 0
6 1 9 3 9 13 13
8 9 0 3 13 0 13 0 13
6 1 9 3 9 9 13
15 0 9 1 0 9 13 0 7 0 9 1 0 9 13 0
18 13 3 15 16 0 9 0 15 3 13 9 13 1 15 9 1 9 0
11 1 9 3 15 13 15 7 9 15 13 15
5 0 3 13 13 15
16 9 0 7 0 9 13 7 9 3 13 15 15 3 9 11 9
24 3 3 13 11 1 9 0 12 9 7 12 9 3 13 9 0 1 9 9 12 9 7 12 9
21 9 0 13 1 9 1 9 0 7 13 15 16 13 15 9 0 7 6 0 11 3
16 3 3 0 9 13 1 9 13 1 0 9 13 9 7 3 13
2 3 13
7 13 15 1 9 15 3 13
22 3 13 7 13 1 15 12 15 9 0 15 7 13 13 3 7 13 0 9 0 0 0
15 3 15 13 1 9 6 9 7 9 15 13 3 13 13 15
5 13 3 1 15 15
12 6 9 15 7 9 15 3 13 13 13 1 15
6 0 3 13 13 1 13
9 15 13 9 15 7 15 13 9 15
7 7 13 9 1 9 15 13
19 15 3 3 13 9 9 15 15 13 1 9 0 9 15 7 9 7 9 13
11 1 0 3 9 13 11 1 9 13 1 9
6 7 13 15 3 9 13
5 6 13 13 16 13
14 7 13 0 3 13 1 9 7 13 9 0 7 13 15
18 0 3 13 1 9 15 3 13 9 0 7 3 13 16 3 13 9 9
10 9 3 13 13 7 16 3 13 9 13
17 0 3 13 1 9 0 7 13 9 0 12 0 12 12 0 12 12
5 13 9 13 3 13
5 7 13 9 13 15
4 0 3 13 13
8 3 15 13 13 13 0 9 0
5 0 3 3 13 13
7 13 3 13 15 7 13 15
15 0 1 9 15 13 16 13 3 13 7 13 3 13 7 13
7 7 13 15 15 9 0 13
6 9 13 7 3 13 13
7 7 13 13 7 3 13 13
11 15 3 0 9 16 13 7 9 15 16 13
23 6 3 13 15 16 0 9 7 9 13 13 15 13 7 3 13 7 13 15 13 7 3 13
5 15 3 13 9 13
5 0 13 13 1 9
14 7 13 1 9 0 13 13 9 7 3 1 9 13 15
9 3 13 3 9 1 15 7 3 13
10 13 3 9 7 9 9 1 3 13 15
21 7 13 1 9 0 13 13 9 7 9 9 0 7 9 9 13 15 7 1 9 13
5 15 9 13 15 13
11 13 15 9 0 9 13 0 9 1 9 15
12 3 3 13 9 7 9 13 3 13 15 3 9
6 13 3 9 9 13 15
10 9 3 0 3 9 13 13 1 9 15
4 3 3 13 9
4 0 3 13 15
4 9 9 0 13
7 13 3 3 16 13 13 15
10 3 16 13 9 13 3 1 15 3 9
13 13 15 3 13 3 1 9 7 1 9 9 13 9
17 13 3 9 7 13 15 1 9 16 13 15 7 9 13 1 9 15
5 15 9 13 15 13
13 0 13 9 0 9 0 15 13 9 13 1 9 15
5 15 0 13 15 9
18 3 3 13 0 9 13 7 13 9 16 13 9 0 7 13 1 9 15
19 15 13 11 9 1 9 7 1 9 15 13 1 15 16 13 15 13 9 13
5 13 1 9 9 15
6 13 13 1 9 15 9
7 3 13 9 13 1 9 11
7 7 13 1 15 9 15 13
5 13 15 9 9 0
5 0 3 13 13 15
6 13 13 0 9 9 0
7 0 3 9 0 13 9 9
5 7 9 13 9 0
6 7 9 13 13 15 9
9 7 9 13 9 9 7 9 13 9
14 3 3 3 13 9 7 9 13 3 13 1 9 9 0
21 13 9 0 9 15 7 13 1 9 15 15 9 7 13 9 7 13 15 1 9 0
6 3 13 9 7 9 9
5 13 9 13 3 13
24 3 0 13 9 0 9 9 13 0 9 15 13 12 0 9 13 13 15 9 15 13 7 13 15
14 3 0 13 9 0 9 13 1 9 7 1 0 9 13
18 15 3 13 15 13 15 1 9 7 13 13 0 1 9 7 0 13 3
5 3 13 1 9 9
8 13 9 7 13 0 1 9 0
6 7 13 15 1 9 0
6 3 13 9 7 9 9
4 13 3 15 0
4 11 3 13 15
20 0 1 0 9 13 15 9 0 0 13 9 0 15 13 1 9 15 0 7 0
7 7 13 3 13 11 9 0
2 13 3
16 7 13 1 9 15 13 15 1 9 15 16 13 15 15 7 13
7 3 0 13 9 0 7 9
7 3 9 3 15 13 15 11
9 7 9 15 11 7 11 7 11 11
6 3 3 0 15 0 13
5 7 13 15 1 15
4 11 3 13 15
11 13 9 0 3 1 15 9 7 1 9 15
9 7 3 13 3 9 0 1 9 15
4 0 13 11 9
12 0 13 1 0 7 0 1 9 13 15 1 15
17 11 3 13 11 13 15 7 13 15 1 9 11 1 9 11 9 15
5 3 13 15 13 15
12 7 13 15 13 13 15 9 16 3 9 13 15
13 9 3 13 9 0 13 9 0 1 9 7 13 11
10 0 3 1 9 13 15 13 15 3 13
4 7 0 13 9
16 9 3 1 7 13 1 15 13 13 15 7 13 13 11 1 9
13 7 13 9 15 1 9 7 13 9 7 13 9 15
14 7 13 9 15 13 9 15 7 13 15 7 13 13 11
9 7 13 9 1 15 13 0 1 9
14 7 13 11 13 9 0 7 13 1 15 7 13 0 15
9 3 3 13 13 1 15 9 15 13
4 7 9 13 3
10 13 9 16 13 1 0 9 13 9 15
4 11 3 13 15
3 3 13 13
4 13 15 15 13
9 3 13 3 3 12 9 7 12 9
3 0 3 13
25 7 13 9 13 1 9 7 13 12 9 7 12 9 13 1 9 13 7 13 9 13 9 9 3 9
15 7 13 15 7 13 15 7 13 9 9 12 1 12 9 0
11 13 3 13 9 3 12 12 1 9 7 9
17 7 3 13 11 9 13 1 9 7 13 15 1 0 9 16 13 9
9 7 13 9 13 1 9 12 13 15
6 3 3 13 12 13 3
4 13 3 0 9
13 7 13 15 9 13 1 9 13 15 13 16 9 13
4 7 1 9 13
6 3 3 13 15 11 13
1 13
2 15 13
3 3 13 15
5 13 3 11 13 15
1 13
8 7 13 1 9 11 13 1 9
4 7 13 1 11
11 13 3 9 0 13 15 7 13 13 13 13
3 9 13 15
7 3 3 11 13 9 13 15
3 7 13 15
5 0 1 15 15 13
9 13 3 1 9 13 13 15 15 13
5 1 9 9 0 13
6 7 13 13 1 9 0
27 7 13 15 9 9 0 13 1 15 9 0 7 13 1 15 15 13 7 13 15 16 3 13 15 9 9 15
7 7 15 13 15 15 13 13
12 3 13 1 11 15 13 1 11 9 7 9 13
7 1 15 9 15 13 9 9
8 3 13 3 9 15 3 9 13
4 9 3 13 13
4 13 9 7 9
8 7 15 13 9 7 9 9 13
3 15 3 13
21 15 3 13 9 7 9 9 15 3 1 15 13 15 13 15 3 13 9 7 9 15
7 7 13 9 0 1 9 15
7 9 3 13 1 15 11 13
8 3 3 13 15 13 9 9 0
3 13 7 13
13 3 13 1 9 13 9 7 13 1 9 0 13 9
6 3 13 9 15 13 15
8 13 3 16 9 13 9 13 15
4 0 3 13 13
10 0 9 15 3 13 9 15 0 13 15
4 9 13 0 9
10 9 3 9 16 13 12 1 9 13 15
4 13 15 9 0
4 11 3 13 15
7 3 3 3 15 1 9 13
17 3 3 3 13 16 0 15 13 1 9 1 9 13 15 7 9 13
11 7 13 1 9 1 9 13 7 0 13 9
4 0 13 13 9
9 7 10 3 13 9 13 3 13 9
10 7 13 3 11 13 1 9 0 7 0
5 13 15 9 9 0
5 9 15 3 13 15
6 0 3 3 13 15 9
7 7 13 9 15 13 15 13
4 0 3 13 13
8 13 13 3 1 9 13 9 0
7 0 3 13 13 15 15 13
3 9 13 15
8 13 0 13 9 9 7 13 9
3 0 3 13
13 6 9 3 3 9 13 1 9 13 1 9 9 15
6 6 9 0 13 9 15
4 13 15 3 13
7 7 13 9 15 1 0 9
14 7 13 3 11 13 1 9 0 7 13 1 9 13 3
24 7 13 1 15 9 0 13 1 15 0 0 7 0 7 0 7 15 0 7 13 15 1 9 0
4 7 13 9 0
7 11 3 13 9 15 13 15
13 7 13 15 3 13 3 13 16 3 3 13 1 9
4 7 13 15 9
9 3 13 1 0 9 9 13 3 9
4 7 13 15 11
3 3 9 13
3 0 3 13
22 7 13 9 13 1 9 7 13 12 9 7 9 9 13 13 7 13 9 15 9 3 9
10 7 13 13 12 12 9 1 9 7 9
11 7 13 9 13 1 9 7 13 1 9 0
13 7 13 9 7 9 13 15 13 9 1 9 13 15
5 0 3 13 13 15
3 3 13 13
1 9
3 13 15 9
5 13 3 15 13 9
10 9 3 9 13 13 7 9 9 3 13
6 9 0 7 0 9 13
10 7 9 3 13 15 15 3 9 11 9
4 7 13 15 13
10 7 13 9 15 1 0 9 13 9 13
4 11 3 13 15
9 13 7 13 15 1 9 0 7 0
4 3 9 3 13
4 13 3 11 13
9 15 13 1 15 0 16 9 3 13
14 3 3 3 13 7 13 12 9 12 12 7 3 9 13
10 3 3 12 9 12 12 7 3 9 13
10 3 3 13 16 3 1 9 15 13 13
8 13 3 15 1 9 0 7 0
4 3 13 16 13
7 15 13 15 9 13 9 0
4 0 3 13 15
3 0 11 9
3 15 3 11
7 0 3 11 7 12 1 9
3 13 15 11
6 15 3 15 15 13 13
6 15 13 11 9 9 0
18 0 13 11 11 16 9 7 9 3 13 15 7 9 15 15 13 1 9
22 7 15 3 15 13 16 15 13 11 7 1 0 9 13 9 15 7 9 0 3 13 15
26 7 13 15 9 9 0 7 15 3 13 1 9 13 13 1 9 7 15 3 13 1 9 13 13 1 9
9 3 13 9 15 16 15 3 13 16
4 0 13 11 11
28 3 13 11 13 9 15 16 13 15 13 1 11 7 3 13 1 9 7 9 7 9 7 13 13 7 0 9 13
3 0 15 9
5 3 13 15 13 0
3 13 1 15
12 9 9 15 13 16 3 13 15 13 0 7 0
5 3 11 13 9 15
19 16 15 13 1 15 13 3 13 15 15 7 13 9 15 7 1 9 15 13
8 15 3 13 9 15 13 13 15
12 15 9 13 9 16 15 9 13 7 9 15 13
8 7 15 13 9 9 1 9 15
19 13 3 13 9 0 1 9 9 15 1 9 0 7 3 13 15 1 9 15
21 7 13 1 12 9 13 11 11 7 11 7 11 9 15 7 13 15 1 9 0 12
19 7 13 15 1 15 7 13 15 9 15 3 9 7 9 15 13 0 3 9
11 7 6 13 15 15 11 7 11 1 15 13
6 13 3 11 1 11 13
15 16 13 3 13 3 12 9 15 12 7 11 12 7 11 12
15 3 3 15 13 6 9 0 13 15 7 6 9 1 9 13
8 0 13 9 15 13 1 15 13
2 0 13
6 7 13 11 13 15 15
2 7 13
5 13 7 3 13 15
9 7 13 15 1 9 13 15 11 13
10 15 3 13 9 16 9 0 1 0 13
6 7 13 15 9 15 13
9 15 3 13 9 16 11 13 13 3
5 11 3 13 13 15
18 13 3 15 16 11 3 13 7 3 13 15 7 13 1 15 15 15 13
8 3 3 9 0 13 13 1 15
14 7 13 15 1 9 13 1 15 9 13 15 15 7 13
13 9 13 9 15 16 1 0 9 13 15 7 3 13
9 3 3 13 1 9 7 3 1 9
11 7 13 15 1 9 15 7 3 13 15 13
4 13 3 11 13
9 6 9 0 7 13 3 1 15 13
4 13 15 15 3
6 3 13 9 11 12 13
7 1 15 15 3 13 13 15
4 11 3 13 15
3 1 9 15
4 6 3 13 15
9 16 13 9 3 9 0 13 9 0
3 13 3 3
9 9 3 0 3 13 3 9 7 9
8 13 3 15 1 11 13 15 11
15 13 13 13 9 0 1 9 9 7 13 15 7 0 9 13
4 7 0 13 3
12 13 3 15 1 11 13 13 9 1 11 7 13
6 9 15 3 13 3 9
2 13 6
8 7 3 13 1 9 13 11 13
8 9 0 1 15 13 9 7 9
7 1 15 3 9 7 1 0
4 7 13 15 11
2 1 0
3 13 15 11
4 3 0 13 9
23 7 16 3 13 15 13 1 9 13 9 7 15 13 3 9 13 7 13 9 15 7 13 9
9 0 13 13 15 1 15 7 1 15
11 7 13 11 9 13 15 1 9 15 7 13
3 6 13 15
14 16 3 13 15 7 13 3 9 3 13 13 1 9 0
13 15 3 15 13 3 9 0 0 13 0 1 9 0
12 7 15 3 13 9 0 12 1 9 15 15 13
27 7 15 3 13 12 1 0 0 13 1 15 0 15 13 16 13 9 1 9 15 0 7 13 15 1 9 0
5 6 15 9 1 9
7 3 6 9 0 15 9 13
21 0 15 13 13 1 9 0 7 0 3 12 9 7 12 9 13 13 13 1 9 0
12 7 16 9 15 13 15 13 15 7 13 1 15
18 0 15 13 1 12 9 1 9 13 3 12 9 13 13 13 1 9 0
10 13 15 7 3 13 1 12 1 0 0
14 13 3 15 16 9 15 1 9 3 13 9 9 15 0
8 13 3 9 0 13 7 13 13
24 16 13 15 9 12 9 7 13 12 1 15 3 13 3 12 12 7 12 1 9 7 13 13 13
21 7 16 13 15 6 13 15 16 13 15 1 15 3 3 1 12 12 7 12 3 13
15 16 3 13 1 15 9 15 13 13 15 1 15 7 0 12
6 16 15 13 13 9 15
22 16 3 15 3 13 13 3 1 15 12 7 12 16 1 9 12 7 12 9 13 0 9
7 16 3 3 13 15 13 9
15 16 3 3 1 9 3 13 13 3 13 15 3 9 7 9
19 15 3 13 1 9 13 13 1 9 7 15 3 13 1 9 13 13 1 9
27 3 6 13 15 16 16 12 1 15 13 1 9 1 0 9 15 3 13 13 15 1 9 15 15 13 1 9
15 3 3 13 12 7 12 13 1 9 15 3 13 1 9 15
11 9 3 9 13 9 15 1 15 7 13 15
4 1 12 9 3
3 13 15 11
12 3 13 15 1 12 9 7 1 12 12 9 3
13 13 3 15 13 15 1 9 13 15 9 15 9 9
23 3 13 3 15 13 13 9 15 16 13 15 7 9 15 7 9 7 15 15 13 7 13 15
8 13 3 9 0 13 15 15 13
8 9 13 1 15 7 15 13 15
20 13 3 9 0 13 12 1 9 15 15 13 0 15 12 9 7 13 13 15 13
5 13 15 15 13 0
6 13 3 9 13 15 13
15 0 3 3 13 7 13 13 15 1 9 16 13 15 15 9
15 13 3 3 9 13 13 15 3 7 13 13 9 15 15 13
7 3 13 15 9 15 13 15
10 9 0 15 9 15 13 15 16 13 15
13 3 13 3 3 15 13 9 15 3 3 15 15 13
16 3 3 9 15 0 13 15 16 3 13 15 9 15 1 9 15
19 7 13 3 13 11 9 0 13 1 11 7 13 1 9 0 1 0 9 11
8 7 13 1 15 9 13 15 13
9 3 13 9 13 9 15 1 0 9
5 0 3 13 13 15
12 13 3 13 16 13 3 0 9 7 0 13 13
2 7 13
9 0 1 13 9 9 15 7 9 15
8 0 3 3 13 12 7 12 9
2 13 15
10 15 3 11 13 13 9 0 7 13 15
3 13 15 16
9 11 1 9 15 13 15 13 9 15
5 3 3 3 13 3
22 13 3 15 16 15 3 13 9 15 1 9 0 13 15 9 13 7 13 15 9 9 13
5 7 13 15 9 15
9 3 15 13 9 0 7 15 13 13
26 13 3 9 15 1 9 0 13 15 3 7 13 9 15 13 9 7 13 9 15 13 15 0 9 1 0
4 13 13 3 13
13 3 13 1 15 9 16 9 13 1 15 7 13 15
4 9 3 13 15
4 11 3 13 15
9 13 9 7 3 13 15 13 1 15
5 0 3 13 9 0
6 7 6 15 13 13 15
9 9 0 15 0 13 16 13 9 0
4 0 3 13 15
4 15 15 13 0
5 15 0 3 12 9
8 16 3 13 1 9 13 13 9
2 13 15
1 15
3 13 15 9
6 15 0 13 1 9 15
5 15 13 3 3 13
3 13 15 11
22 16 13 13 13 13 13 9 15 7 13 0 7 13 13 9 1 9 7 13 1 9 15
6 13 3 9 9 13 13
5 13 3 13 9 0
10 6 13 15 16 3 13 0 1 9 0
7 13 3 9 13 15 3 13
5 15 3 13 13 13
5 13 3 11 13 15
10 1 9 0 0 13 7 1 9 15 0
5 3 13 11 13 15
10 9 6 15 13 15 7 1 9 15 13
3 11 13 15
4 6 13 15 16
28 7 0 15 13 9 7 9 7 9 7 9 7 9 7 9 7 9 7 9 9 15 1 3 13 7 9 0 13
8 0 3 13 0 0 7 0 0
14 0 13 9 0 9 0 15 13 3 3 13 9 9 15
13 13 3 1 9 1 9 1 9 13 15 1 9 15
14 7 13 1 0 9 13 15 1 9 13 0 7 0 13
6 7 15 13 9 13 15
3 0 3 13
11 3 3 13 1 0 7 1 0 9 13 3
3 7 13 15
6 15 13 3 15 9 0
4 7 13 15 16
4 15 15 3 13
6 13 3 15 1 9 15
5 7 15 13 9 13
9 9 3 13 13 9 9 1 9 15
2 13 9
11 13 3 15 1 12 1 12 9 13 1 9
7 7 13 0 13 15 3 13
4 7 13 1 9
17 3 0 0 12 9 13 7 0 15 13 15 13 13 9 9 7 9
6 0 3 13 13 15 15
4 9 3 13 15
7 3 1 9 3 13 1 15
4 13 15 7 13
10 16 13 15 9 13 1 15 15 15 13
9 3 9 15 0 13 16 15 0 13
7 0 3 13 13 3 3 13
16 7 13 11 1 11 13 12 1 12 9 12 1 9 7 13 15
17 6 13 1 11 7 9 0 13 13 9 7 9 7 13 15 1 9
15 7 13 15 1 9 9 7 9 7 9 7 1 0 9 13
17 3 13 1 15 9 9 0 1 9 15 13 15 7 13 15 1 15
4 0 3 13 15
2 13 15
4 13 3 11 13
5 3 13 15 15 13
16 13 3 13 9 15 15 13 13 7 9 15 15 13 15 13 15
2 13 15
1 13
3 7 13 15
3 9 15 13
7 7 15 13 13 1 9 15
7 7 13 9 13 1 12 9
5 11 3 13 15 13
10 13 16 9 9 13 15 7 0 13 0
6 3 3 3 13 1 15
12 7 15 3 13 0 13 1 15 3 13 15 9
12 7 15 3 13 1 15 13 0 3 13 15 9
18 3 9 0 3 13 3 16 13 15 7 13 7 13 9 15 9 1 0
14 7 6 12 9 13 1 9 7 13 16 11 13 13 13
5 13 15 9 9 0
6 9 3 13 15 16 13
5 0 3 3 13 13
5 13 15 9 9 0
7 7 13 11 13 15 7 13
5 15 13 16 13 15
2 13 15
19 7 3 13 15 1 11 7 13 1 11 1 9 0 3 11 13 12 9 15
3 7 13 15
16 13 1 9 15 13 1 15 7 3 13 9 13 7 9 1 15
5 7 13 13 15 15
11 7 16 13 15 15 15 13 16 9 13 15
5 7 3 3 13 15
10 0 3 15 13 16 13 15 13 9 13
14 6 9 15 13 15 0 7 13 1 9 7 9 9 0
8 0 3 9 13 9 15 1 9
10 0 3 13 9 1 9 7 13 1 9
10 9 3 13 1 15 7 1 9 13 13
11 6 9 0 0 13 1 9 0 6 1 0
10 7 13 15 1 11 13 15 15 9 13
3 15 0 13
8 0 13 11 9 15 1 11 0
25 7 13 11 1 9 0 7 13 15 13 7 13 1 9 7 9 9 13 7 9 13 9 7 13 15
6 9 15 9 9 13 15
6 15 3 13 15 9 9
12 7 13 1 15 0 7 0 1 9 7 13 15
22 13 3 9 7 9 9 15 13 7 9 13 1 9 7 13 6 9 0 13 7 13 15
5 13 3 15 0 13
1 6
13 13 3 13 3 16 1 9 0 7 13 13 13 9
13 7 13 15 13 3 1 9 1 11 7 13 15 3
21 7 13 9 12 1 9 13 1 15 7 15 3 13 1 15 3 9 12 7 13 15
9 3 3 9 1 15 3 13 1 9
4 7 3 13 9
6 7 13 9 13 15 13
5 13 3 11 13 15
3 6 13 15
25 16 13 9 7 3 13 15 3 3 0 13 7 16 3 9 0 13 13 15 7 13 15 1 9 13
8 7 15 15 13 1 9 13 13
10 15 9 0 13 7 15 15 13 9 0
5 13 3 11 13 15
18 13 15 3 15 12 9 15 16 13 15 3 15 15 13 15 9 0 13
6 0 3 13 1 15 13
11 16 13 1 9 1 15 3 3 13 15 9
8 16 3 13 1 9 13 15 9
6 15 3 3 9 13 11
4 13 3 11 13
4 13 15 7 0
8 3 15 13 15 15 9 0 13
5 9 15 13 12 9
5 7 13 1 0 13
3 9 13 3
4 13 1 9 15
4 0 3 13 13
2 3 13
6 7 13 1 0 13 3
3 15 13 9
3 7 3 13
6 15 1 12 13 9 0
2 13 15
1 0
3 13 15 11
12 6 13 15 16 9 7 9 13 15 1 9 0
11 15 3 13 15 3 13 15 3 13 15 9
3 15 9 13
26 9 13 0 15 13 9 7 9 15 13 7 13 1 15 9 7 13 1 15 9 7 13 15 9 7 13
14 3 3 13 15 9 9 13 9 15 1 9 13 9 15
14 13 3 9 9 15 0 13 0 3 13 0 3 9 13
10 3 13 15 9 0 0 7 13 15 3
8 3 3 13 1 15 9 15 13
4 13 15 9 15
3 0 13 9
1 13
6 13 15 7 13 9 15
10 7 13 15 13 3 1 9 7 13 15
10 3 3 3 13 9 9 15 13 9 0
4 0 3 13 15
12 7 9 13 15 9 15 13 15 9 1 9 15
3 13 15 11
10 1 9 13 0 7 13 0 1 9 15
31 0 1 13 15 16 13 15 1 15 9 0 7 13 15 9 13 9 15 7 13 1 9 0 13 15 7 1 15 13 13 15
12 7 13 9 7 9 9 15 13 16 1 15 13
12 7 13 13 15 13 15 9 16 3 9 13 15
8 7 13 11 13 15 1 9 13
11 13 15 9 0 9 9 15 13 9 9 15
12 7 13 9 15 13 13 1 9 7 3 13 13
2 13 13
8 9 15 7 0 13 7 15 13
3 13 1 9
13 0 3 3 13 13 0 1 9 15 0 1 9 15
10 7 0 13 9 15 13 15 7 13 15
17 7 13 9 0 13 15 7 13 9 15 13 9 0 7 9 15 13
4 3 13 9 15
5 7 13 3 13 0
12 13 3 1 9 9 7 15 3 13 13 1 9
13 13 3 9 13 13 13 3 9 3 13 1 9 0
3 7 13 15
8 9 3 13 3 3 13 9 0
3 0 3 13
4 3 13 9 9
6 3 13 9 7 9 9
7 0 3 13 13 3 3 13
11 3 13 9 9 13 1 15 16 13 15 9
5 9 13 16 0 13
10 9 0 1 9 13 7 15 1 3 13
6 3 13 3 1 9 9
7 13 3 15 15 15 15 13
6 13 3 11 9 15 13
4 15 15 13 9
4 13 15 9 0
5 0 3 13 15 9
6 15 13 9 0 7 9
2 13 15
1 0
7 13 3 0 9 7 0 9
8 7 13 13 15 7 13 15 13
15 1 0 9 13 1 15 13 9 3 13 9 7 13 15 13
3 9 11 13
16 16 15 13 3 13 9 16 13 9 9 15 7 13 9 9 15
7 3 7 0 7 0 1 0
7 1 3 15 15 13 3 9
4 15 3 13 15
5 13 3 11 13 15
7 13 3 13 9 7 9 0
15 1 9 3 7 13 15 7 13 7 3 9 0 1 9 13
11 1 9 3 0 13 3 13 13 15 9 13
10 15 13 9 0 7 9 0 7 9 0
8 7 13 9 13 15 1 9 15
7 9 15 9 13 0 1 9
4 11 3 13 15
15 13 9 9 15 15 9 15 7 15 9 15 7 15 9 15
6 0 13 0 7 0 9
4 0 3 0 15
6 13 0 15 3 0 15
9 1 0 12 9 15 9 7 9 13
3 15 13 9
2 13 15
1 0
2 13 15
8 3 3 11 9 13 15 9 13
4 13 9 9 15
11 13 1 0 15 16 13 9 15 9 9 15
11 16 3 11 9 9 13 15 3 15 13 9
10 3 13 15 1 9 0 13 15 1 0
9 3 11 13 1 9 7 9 15 13
7 1 0 9 13 9 7 9
10 15 3 15 3 13 15 13 13 7 13
6 1 9 3 15 3 13
5 13 3 7 3 13
12 13 3 9 0 7 3 13 7 13 1 9 0
7 7 9 15 3 13 13 15
6 7 13 9 9 9 15
19 13 3 9 1 9 7 9 1 9 7 9 1 9 7 13 15 1 9 9
6 15 3 3 13 15 9
6 12 3 13 15 9 11
5 15 3 15 9 13
7 7 9 3 13 15 1 9
9 12 3 13 9 15 15 13 1 9
7 7 0 15 3 13 15 9
11 6 15 9 7 9 7 9 16 13 9 9
10 7 9 3 9 13 0 1 13 0 9
12 6 15 9 7 9 9 16 13 9 0 1 9
4 15 3 3 13
4 7 13 13 13
23 6 15 9 7 9 9 16 13 9 7 9 13 12 9 7 3 13 13 15 9 9 0 15
7 15 3 13 15 9 15 13
8 7 15 13 15 9 0 0 13
6 9 3 7 9 13 9
8 7 15 3 13 15 9 15 13
11 7 15 13 15 9 15 13 1 15 0 13
7 0 7 0 15 3 13 0
6 9 3 7 9 13 9
11 7 13 15 9 13 15 15 7 13 1 15
12 7 13 15 9 13 15 9 0 7 13 1 15
22 6 15 9 7 9 9 16 13 9 7 9 7 9 7 13 0 9 9 7 9 7 9
7 9 0 13 9 7 9 13
19 6 15 9 7 9 9 16 13 0 9 7 9 3 3 13 0 9 7 9
14 9 0 13 3 0 9 7 9 16 13 3 0 15 3
25 6 15 9 7 9 9 16 13 15 9 13 15 3 3 13 0 3 3 0 13 9 0 7 0 9
7 3 3 13 0 9 7 9
17 6 15 9 7 9 7 9 16 13 9 0 7 13 9 0 7 13
16 16 13 13 1 9 9 15 3 13 3 9 15 13 1 9 9
10 0 3 0 13 15 16 9 13 13 9
8 9 9 0 3 13 1 9 0
12 0 1 6 15 13 1 15 9 7 0 7 9
19 7 1 15 13 7 13 7 1 15 13 1 9 15 7 13 1 9 1 9
3 6 13 15
6 13 15 0 1 9 0
25 11 13 9 7 9 13 13 1 15 3 9 13 13 9 15 3 13 9 9 15 1 9 7 3 13
7 6 13 15 15 9 15 0
3 13 3 15
5 0 13 1 9 0
16 7 13 11 1 9 13 7 13 1 15 9 15 13 15 9 0
5 3 13 3 15 0
3 6 13 15
11 3 13 3 13 9 1 9 15 3 13 15
13 13 3 15 1 9 0 13 1 15 9 15 12 13
14 13 15 3 0 13 7 15 13 9 15 9 7 9 9
5 7 13 11 13 15
5 15 15 3 3 13
3 15 13 11
3 7 0 13
7 13 3 13 9 7 9 9
1 13
3 3 13 15
4 13 3 15 13
5 7 3 3 13 9
16 3 13 15 1 9 7 13 15 7 13 13 15 9 9 15 1
13 7 3 13 15 0 7 15 15 13 7 13 15 15
8 7 0 0 9 13 7 13 0
7 7 1 9 9 13 9 0
7 13 3 1 9 0 13 15
16 7 13 15 9 9 1 15 9 1 9 15 9 7 3 13 9
49 3 3 13 9 9 13 11 9 13 1 9 15 13 16 13 3 13 1 11 3 13 1 9 7 15 1 9 3 3 13 13 15 13 1 9 15 7 15 1 9 3 3 3 13 15 3 13 9 15
8 6 3 0 7 13 1 0 9
16 13 3 3 9 0 15 13 13 1 9 15 9 3 7 13 13
15 7 16 3 13 13 15 9 0 3 13 3 13 15 0 9
7 1 13 3 13 15 9 0
13 3 16 15 15 13 6 3 11 7 3 3 13 9
19 13 3 0 11 7 0 9 7 13 9 0 7 9 16 13 16 13 0 13
4 6 3 13 15
10 16 3 13 15 6 1 9 13 3 13
3 6 1 9
9 3 3 3 13 9 3 13 15 9
24 3 3 1 9 9 0 9 13 7 9 3 13 9 15 7 9 13 1 9 7 9 0 13 15
29 7 3 13 15 9 9 0 1 9 7 3 13 15 15 9 0 7 13 9 0 13 1 9 0 1 9 7 9 0
20 7 13 9 1 9 0 0 7 13 13 15 1 12 9 1 9 9 1 9 15
6 1 9 3 13 15 9
14 3 3 9 15 13 0 7 9 13 13 16 1 13 9
13 3 3 15 3 13 15 0 13 16 1 13 1 9
9 9 7 9 13 7 9 15 3 13
12 3 3 1 9 0 3 13 3 1 9 9 0
36 3 3 13 1 9 1 9 13 7 13 13 15 7 13 1 15 9 13 11 1 9 7 3 13 16 13 9 7 13 15 3 13 3 9 9 0
5 3 12 13 1 9
2 12 13
4 7 0 13 15
4 12 13 1 9
11 13 3 16 3 13 1 15 9 9 15 13
24 0 3 13 16 16 13 13 9 9 1 15 9 9 13 13 3 13 7 3 13 13 13 9 15
20 15 3 13 0 9 7 0 15 13 9 1 9 15 16 13 15 1 9 9 15
10 0 9 0 15 13 9 15 13 3 13
9 6 13 15 16 1 15 9 13 15
50 16 3 13 0 9 1 9 15 13 15 9 13 7 13 13 9 15 13 3 7 13 1 9 13 9 9 0 1 9 1 15 3 13 7 1 9 1 15 3 13 7 13 15 9 7 9 15 1 9 13
6 3 13 9 7 9 9
9 12 3 13 1 15 0 7 12 0
10 0 3 13 9 15 3 13 1 15 9
9 7 0 13 9 1 9 1 9 15
5 9 9 3 9 13
3 6 9 13
4 13 1 9 15
9 3 13 9 15 15 7 13 9 15
9 13 15 1 9 15 16 9 15 13
4 13 3 0 13
6 3 3 13 15 7 15
8 13 3 3 1 13 7 13 15
7 3 3 13 3 0 9 13
4 9 9 13 15
4 0 3 13 13
3 3 13 15
8 13 3 16 3 13 9 7 9
31 3 3 9 13 13 15 9 7 13 15 9 15 7 0 3 13 12 9 0 3 12 0 3 12 15 3 9 15 7 13 3
13 13 3 13 12 9 13 1 15 7 13 0 12 9
7 3 3 15 12 13 0 12
15 1 0 3 9 13 9 9 0 7 13 15 1 15 1 9
10 7 13 13 12 9 13 0 12 9 13
6 6 0 12 9 13 15
4 13 15 9 15
10 0 9 7 0 7 0 1 0 13 0
4 1 0 15 13
5 13 1 9 9 15
7 13 3 3 13 12 9 13
5 6 0 12 13 15
9 0 9 0 7 0 1 0 13 0
4 1 0 15 13
5 13 1 9 9 15
8 13 3 3 13 12 9 13 9
15 13 15 16 0 13 9 13 3 13 13 7 13 3 3 13
9 7 13 15 13 13 9 15 1 9
3 6 13 15
16 13 15 3 13 9 15 9 7 13 15 13 3 13 15 1 9
10 13 3 1 15 9 7 13 13 12 9
7 13 3 3 13 13 7 13
14 7 1 3 13 3 15 3 13 15 13 13 13 1 15
7 7 0 9 13 1 9 0
6 3 13 9 7 9 9
18 3 13 9 0 1 9 15 7 15 9 1 15 3 13 1 9 9 15
29 7 13 15 1 15 15 9 7 13 15 15 1 15 3 9 13 9 1 9 7 13 9 1 0 15 7 9 1 0
4 13 0 9 15
8 13 13 15 9 1 9 15 9
7 13 3 15 7 13 15 13
5 13 15 7 13 15
5 0 13 7 13 15
4 0 7 13 15
4 13 7 13 15
7 1 9 13 7 13 1 15
4 7 13 7 13
7 3 3 15 13 0 7 13
4 7 0 7 13
12 3 3 15 13 13 7 1 9 7 13 1 15
5 7 13 9 13 15
3 6 13 15
11 16 13 12 1 0 0 9 15 0 15 13
12 13 1 15 13 1 9 0 13 9 7 9 15
6 13 15 7 3 13 15
6 0 13 7 3 13 15
5 0 7 3 13 15
8 0 7 1 9 7 3 13 15
5 3 13 3 0 13
20 9 3 15 13 13 7 13 7 0 7 0 7 0 7 1 9 7 3 13 15
3 6 13 15
10 16 3 13 12 1 0 0 3 15 13
11 7 13 3 13 11 15 9 0 13 9 15
14 13 16 1 12 9 9 13 7 9 0 13 13 1 9
23 3 13 15 9 7 9 7 9 0 1 9 0 13 11 7 9 13 16 11 9 13 7 13
2 13 3
10 7 3 1 9 16 3 9 13 1 9
6 13 3 9 15 13 13
4 15 1 9 0
12 13 3 0 9 13 13 1 0 7 13 13 0
3 15 13 9
6 9 3 0 13 1 15
6 3 3 0 13 1 15
5 15 3 3 3 13
3 6 13 15
18 3 3 13 13 9 0 1 15 9 13 15 3 15 13 0 1 9 15
12 3 13 1 12 1 12 13 11 0 1 9 13
9 15 13 15 13 7 15 15 13 15
8 7 3 13 0 9 16 15 13
12 1 0 3 9 9 13 9 1 11 13 1 15
6 3 13 13 15 9 13
5 13 1 9 1 15
3 7 13 15
2 9 13
7 1 15 13 9 1 9 15
10 7 13 9 3 13 15 11 7 13 9
4 7 13 15 13
9 6 13 15 16 12 1 15 13 15
4 3 15 13 9
4 0 3 13 13
9 13 1 15 9 1 9 0 15 13
9 9 3 0 13 3 13 13 1 15
9 6 3 9 0 15 9 0 13 15
11 0 13 13 15 16 15 13 3 13 9 0
4 3 15 13 9
2 15 13
9 13 3 15 13 11 9 7 13 13
4 7 13 9 15
2 7 13
1 13
1 13
4 0 13 9 15
12 0 13 9 15 0 9 13 1 0 1 9 9
24 13 3 15 16 3 13 13 3 1 0 9 0 1 0 9 3 13 1 15 0 1 9 9 15
6 7 13 13 1 9 0
4 3 13 15 11
9 15 15 13 15 1 15 1 0 9
3 13 3 13
7 13 9 7 13 15 9 9
8 1 9 3 15 13 15 1 11
12 16 3 15 13 15 1 15 15 3 3 13 15
3 13 15 11
4 6 13 15 16
13 1 0 9 3 16 9 3 13 12 9 13 15 15
3 13 15 11
11 16 15 15 13 1 15 13 3 13 15 15
5 3 7 15 9 13
10 3 13 11 1 9 13 11 7 13 9
4 3 13 15 11
6 0 13 9 15 1 9
6 13 3 7 13 1 15
9 7 13 3 13 0 13 15 7 13
11 9 15 16 0 13 3 13 1 15 9 0
8 3 3 3 15 13 7 3 15
11 7 13 1 9 7 13 15 13 7 13 11
9 13 7 13 15 16 3 13 1 9
6 3 3 13 13 15 13
17 9 15 16 3 13 9 0 13 1 15 16 3 13 15 13 9 15
6 7 13 3 13 15 13
5 13 3 9 15 0
11 7 13 15 3 13 13 15 3 0 9 13
4 3 13 1 9
4 13 3 7 13
12 6 13 15 9 7 9 0 13 15 1 9 9
1 13
5 6 13 15 13 15
26 7 3 13 15 6 11 12 1 12 1 12 13 7 1 15 9 0 1 9 7 9 1 9 7 9 0
7 13 3 15 13 15 9 13
5 15 3 13 0 13
7 7 3 13 1 11 13 15
3 13 15 9
3 7 13 15
5 9 1 15 13 13
9 3 13 13 9 1 11 7 13 15
19 7 6 12 1 13 1 11 13 9 13 9 15 7 13 9 0 13 15 9
4 3 13 15 11
6 15 3 13 9 9 13
21 7 13 15 15 16 3 13 3 13 9 15 7 13 15 3 3 12 1 12 9 9
10 3 3 3 13 15 9 16 3 13 13
6 1 0 9 13 11 9
12 1 15 9 13 1 15 1 9 7 3 13 15
9 0 3 15 13 16 13 15 9 0
6 3 9 9 13 15 13
17 11 3 13 1 15 3 1 9 0 7 13 3 13 1 9 13 9
23 9 3 7 9 7 9 15 13 0 9 1 11 16 3 13 15 7 3 13 0 0 9 13
7 3 3 13 12 0 9 13
2 0 13
9 13 13 9 0 7 12 9 13 15
4 15 3 3 13
5 15 0 1 15 13
5 7 13 9 13 15
13 13 15 9 0 16 13 15 16 15 13 11 9 0
3 13 15 11
2 15 13
3 3 13 15
13 3 13 9 0 13 1 0 9 7 13 1 9 0
2 9 13
5 6 3 13 9 15
4 15 15 15 13
4 0 3 13 13
3 0 13 9
8 3 13 9 15 7 9 15 13
6 0 3 1 9 13 13
2 13 15
7 7 13 1 15 15 9 13
6 3 15 13 1 11 0
7 0 3 13 15 1 15 13
4 3 13 15 13
11 13 3 15 1 9 13 15 0 7 13 15
8 3 3 0 13 9 1 11 9
7 7 3 13 15 1 9 16
3 3 13 9
7 1 9 3 15 1 15 13
7 3 3 9 15 3 15 13
8 3 13 13 15 7 13 15 16
3 3 13 9
4 7 3 9 13
9 7 13 11 9 0 15 13 15 16
10 3 16 9 3 13 12 9 13 15 15
6 7 13 3 13 15 3
18 3 13 11 13 15 16 13 15 13 15 13 12 12 9 9 7 9 13
4 13 13 9 0
3 0 3 13
3 15 13 15
2 15 13
10 7 13 9 1 9 13 7 13 13 15
5 9 3 13 9 13
10 9 3 13 13 15 9 0 1 9 0
6 3 13 15 13 9 13
12 7 13 12 12 9 9 13 15 13 1 9 0
10 7 13 15 1 9 0 3 13 15 9
5 11 3 13 1 9
5 7 13 15 9 13
5 15 3 13 9 0
2 15 13
10 7 3 1 15 13 9 7 9 15 13
7 3 13 3 3 1 15 13
13 7 3 13 15 3 1 12 9 16 13 15 9 3
13 1 0 3 9 0 9 13 9 13 9 9 15 13
7 13 3 3 9 0 13 11
7 13 3 15 15 13 15 11
7 13 3 16 9 1 13 15
11 13 3 15 1 9 13 1 15 9 15 13
5 15 15 7 9 0
12 9 3 7 9 13 9 16 13 11 11 3 13
5 13 3 9 13 15
6 15 13 1 12 13 15
3 0 3 13
3 13 15 11
6 15 3 13 11 13 11
3 13 15 15
3 3 13 13
4 15 3 0 13
5 0 3 3 13 13
3 3 13 13
6 0 13 1 9 0 0
2 15 13
5 7 13 15 9 13
8 9 15 1 15 7 1 9 15
4 3 13 15 11
12 3 9 0 13 11 1 9 13 1 15 15 9
32 7 13 15 9 0 13 15 7 13 9 1 9 13 1 9 15 7 9 1 9 15 7 13 15 1 9 1 15 13 15 15 13
11 7 13 1 15 13 9 7 13 15 1 9
20 7 3 13 15 15 13 1 15 9 7 13 15 1 9 15 7 13 15 1 9
7 13 3 13 9 0 9 11
5 0 13 13 9 15
18 7 13 1 9 13 11 15 13 13 0 9 13 15 9 13 1 9 13
5 7 13 3 13 13
7 7 13 1 9 15 9 13
13 3 13 1 15 12 9 12 1 0 7 12 1 0
9 13 3 13 15 13 9 15 7 13
9 6 13 9 7 12 9 13 13 15
7 16 9 0 13 13 1 9
13 3 3 3 9 13 15 1 9 7 9 7 9 13
2 15 13
9 15 3 3 13 13 16 9 0 13
7 3 13 15 3 16 13 15
3 13 3 16
3 0 9 13
9 3 3 3 9 13 1 15 13 15
12 1 0 3 9 9 13 1 15 9 1 0 9
9 1 0 3 9 13 11 9 0 13
4 8 8 8 8
2 15 13
10 15 3 1 13 3 13 13 16 11 13
17 7 3 13 12 1 15 7 13 9 13 9 7 13 1 9 13 15
3 7 0 13
8 13 16 13 16 13 11 13 15
12 0 3 13 9 13 15 9 7 13 9 7 9
7 11 3 13 9 0 13 9
31 7 6 9 0 13 15 1 0 9 1 0 1 12 7 9 13 15 7 9 13 15 7 9 13 15 7 0 9 13 0 13
15 7 13 1 9 1 9 15 13 1 0 9 7 13 15 0
15 13 3 3 9 0 3 13 15 13 1 11 1 11 13 15
16 1 15 3 13 11 9 7 11 0 7 11 9 7 9 9 0
16 3 3 13 13 9 0 1 11 9 11 15 7 13 15 1 11
7 0 13 1 11 13 9 0
6 11 3 13 13 9 0
28 7 13 9 11 13 15 9 0 7 13 15 1 0 15 9 15 13 1 9 7 13 9 0 1 9 9 7 13
11 13 3 3 11 9 7 0 11 13 1 9
9 9 13 16 9 0 13 3 13 0
18 13 3 13 9 1 0 9 16 3 13 9 15 9 13 15 7 13 9
3 13 1 0
6 7 13 0 9 0 0
3 13 15 11
2 13 9
1 13
9 0 3 13 13 9 13 9 1 9
16 1 9 3 0 13 1 0 9 13 11 9 7 0 11 13 9
17 9 3 0 13 1 9 7 13 13 9 1 9 9 7 13 1 15
12 13 3 9 15 3 9 7 9 15 0 3 9
11 1 9 3 15 13 15 13 7 13 3 0
5 13 3 9 13 9
4 3 13 15 15
2 13 3
4 13 3 3 13
1 13
7 7 3 13 13 9 15 16
9 13 1 0 7 6 13 15 1 11
3 3 15 13
3 6 13 15
6 7 6 11 13 15 13
2 13 15
8 0 3 13 13 15 1 9 15
4 7 13 15 15
3 3 13 15
13 13 7 13 9 15 16 13 1 11 7 3 15 13
14 13 3 15 6 15 1 9 13 1 9 13 9 15 13
8 9 3 13 9 0 13 9 13
2 13 16
8 9 15 9 13 13 15 15 13
15 7 16 0 13 13 1 9 15 13 15 7 15 1 9 13
8 0 3 13 9 13 3 13 13
20 12 3 1 12 9 13 1 11 1 9 3 13 15 11 7 13 15 13 15 15
4 0 3 13 15
10 13 15 13 0 9 1 9 7 1 9
22 13 3 13 15 9 13 15 1 9 9 7 9 7 0 9 13 15 13 15 15 13 15
12 7 6 15 1 15 13 15 9 1 9 9 6
10 9 9 0 9 0 3 13 13 1 9
12 6 15 13 9 15 1 9 15 15 13 9 15
4 9 13 1 9
4 0 13 9 15
21 7 13 1 15 15 0 9 7 9 7 13 15 15 1 0 9 1 15 13 9 15
18 13 3 11 13 9 0 7 9 0 1 9 15 7 9 9 7 9 0
3 7 13 13
15 13 0 15 1 9 15 15 13 0 13 15 13 9 9 15
11 15 3 13 15 9 7 0 13 15 9 0
5 7 13 1 9 0
12 13 11 1 11 0 7 13 15 1 11 1 11
5 15 13 9 15 13
3 1 15 13
7 7 3 9 13 15 1 9
17 7 13 3 1 9 12 9 13 9 7 13 1 9 7 9 13 15
22 1 9 3 0 13 11 1 11 13 9 9 0 13 16 13 15 9 7 13 15 9 0
6 13 15 7 13 1 9
16 13 3 1 9 0 13 11 7 11 9 0 11 13 9 1 9
3 13 3 9
10 13 1 9 15 7 13 15 13 9 9
8 7 3 13 9 15 1 15 13
20 7 13 3 13 11 0 7 11 9 15 7 0 1 9 13 9 7 3 13 15
12 7 13 9 15 11 1 9 1 9 1 15 13
4 7 13 1 11
8 7 3 1 9 1 9 13 15
6 7 13 15 1 9 15
11 13 3 13 3 9 13 7 3 3 9 15
5 15 13 15 7 15
6 11 9 13 13 13 15
4 13 15 15 13
2 0 0
5 7 13 15 11 13
1 13
3 13 1 15
10 7 13 15 15 7 13 15 1 15 13
13 15 9 0 0 16 1 9 9 0 13 7 13 15
9 7 13 9 15 3 1 15 9 0
15 7 3 13 1 9 13 1 9 0 7 0 1 11 7 11
12 9 3 0 13 9 13 7 3 13 15 1 15
7 7 13 13 15 13 1 9
8 7 13 15 3 9 7 13 15
8 7 13 15 9 13 15 1 9
19 7 13 0 0 13 0 9 7 9 0 13 7 3 13 13 9 16 13 15
15 7 13 15 11 7 15 13 1 15 7 13 15 13 15 16
3 15 13 15
3 7 13 15
10 13 1 0 9 7 9 16 3 3 13
4 1 0 3 13
15 7 13 1 15 0 13 15 7 1 9 13 7 13 15 16
5 16 13 13 15 13
10 11 3 13 13 9 13 15 7 13 15
2 13 15
11 7 13 15 3 13 9 1 15 7 0 13
9 7 13 15 3 13 15 7 13 15
2 13 15
16 7 13 13 15 9 7 13 1 9 15 15 13 11 1 9 15
29 0 3 13 13 13 3 7 13 9 16 1 0 3 13 3 1 9 13 7 3 1 0 9 13 7 13 1 15 3
15 7 13 3 11 1 11 1 9 7 9 13 16 1 9 13
18 7 3 13 15 0 16 1 0 3 13 15 3 1 9 7 13 15 9
20 7 3 13 13 1 15 1 9 13 9 3 13 7 13 13 9 1 15 13 13
7 13 3 11 9 15 13 13
6 9 13 15 15 9 15
5 15 0 3 13 9
7 15 13 13 9 3 12 9
14 7 3 13 11 9 15 16 3 0 13 1 15 13 15
6 15 3 13 1 9 15
18 15 13 0 13 13 13 15 15 9 7 13 13 7 13 9 15 7 13
10 13 7 13 9 15 7 13 1 9 15
6 7 13 3 7 13 9
3 3 0 13
5 7 13 3 1 9
9 7 15 9 13 1 15 7 13 15
9 7 13 11 13 11 0 13 1 9
3 7 13 15
3 1 15 13
19 7 13 13 15 1 9 15 7 0 9 7 9 13 1 11 7 1 9 15
17 7 1 15 13 7 9 9 13 15 13 1 9 7 9 13 9 15
7 15 3 1 9 13 7 13
5 7 13 11 13 15
6 3 13 0 9 7 13
8 3 13 13 9 7 9 1 9
8 7 13 9 0 7 9 13 15
5 7 13 7 13 15
11 3 13 9 0 13 15 16 1 15 13 9
10 15 9 1 15 13 9 3 13 13 15
16 13 3 9 3 13 15 1 15 9 7 3 13 15 1 0 9
10 7 15 9 9 3 13 3 13 9 0
15 16 3 3 3 13 9 1 15 0 1 0 7 0 9 13
9 7 15 3 13 9 0 1 9 0
14 16 3 3 3 13 9 0 7 9 13 15 7 9 13
7 7 9 0 1 9 0 13
4 7 9 13 15
1 13
7 15 13 1 9 15 3 13
4 7 0 13 15
41 13 3 3 13 15 13 11 3 13 7 13 15 7 15 13 1 15 3 13 1 9 0 1 11 9 7 9 9 13 15 3 13 13 3 9 7 13 3 13 1 15
3 7 13 15
9 9 9 1 13 7 3 9 9 1
7 0 3 9 13 9 0 9
6 7 13 9 13 0 9
3 13 1 9
3 7 13 15
13 13 3 1 9 0 13 7 0 13 9 13 7 13
3 0 3 13
13 7 13 1 15 1 9 13 1 9 9 15 13 9
3 13 9 15
9 7 13 15 9 15 0 3 3 0
44 11 3 13 1 9 15 1 9 7 0 9 1 11 1 15 13 7 1 11 7 1 11 7 1 11 7 1 0 9 11 7 13 1 11 7 11 0 9 13 15 13 13 1 15
15 7 13 9 15 16 13 1 15 9 9 1 16 3 13 15
13 0 3 13 16 13 15 13 13 15 15 15 13 9
13 7 3 13 15 9 0 13 1 15 7 13 13 16
5 15 13 11 9 0
9 7 3 13 15 16 3 3 13 15
22 7 13 12 1 12 16 13 1 15 7 16 13 15 13 7 13 9 13 9 7 13 9
5 7 13 9 11 11
25 7 11 7 11 7 11 7 11 7 11 7 11 0 7 11 7 11 9 7 11 0 15 3 13 15
4 7 13 1 9
12 7 13 15 3 9 16 3 13 15 3 9 13
9 7 13 15 13 1 15 13 13 15
5 13 3 16 0 13
8 7 13 15 1 9 13 1 15
5 3 13 9 9 13
12 7 16 9 1 15 13 15 3 13 13 9 0
16 7 16 9 13 0 1 15 7 13 15 3 13 13 7 9 13
20 15 3 13 9 0 13 1 9 15 13 16 3 3 0 13 7 3 9 15 13
15 6 13 15 16 15 13 15 9 0 9 7 9 15 3 13
16 7 15 13 1 0 9 3 13 9 1 9 7 0 13 0 9
14 13 3 9 15 7 9 7 3 13 13 1 15 13 15
5 7 13 1 15 9
3 13 3 15
12 6 9 15 7 9 15 7 9 15 3 13 15
7 15 13 9 15 7 9 15
6 7 13 13 3 15 13
6 6 9 15 7 9 15
6 7 3 13 1 9 13
23 7 13 15 1 15 9 0 16 15 13 1 9 13 1 9 7 15 9 13 1 9 1 9
11 7 13 15 9 3 7 13 15 1 9 15
1 13
4 6 13 13 13
10 0 13 1 9 7 13 9 7 13 15
18 7 0 13 1 0 3 3 13 9 0 7 3 13 16 3 13 9 0
15 7 0 13 1 9 7 13 9 7 13 15 7 9 3 13
21 7 0 13 1 9 0 7 13 9 13 7 13 7 13 0 12 12 0 12 0 12
2 7 13
5 13 9 13 3 13
15 3 3 13 12 13 15 15 13 1 15 1 12 1 12 9
3 7 13 15
28 0 3 0 1 9 15 13 16 13 13 7 3 13 7 13 13 7 3 13 16 3 13 15 7 13 15 15 9
5 3 13 3 9 0
5 7 3 15 9 13
3 13 9 13
23 0 3 13 15 1 9 3 13 15 9 7 3 13 3 13 9 7 13 9 13 1 9 15
26 7 0 3 13 15 1 0 13 15 3 13 9 3 1 9 13 15 7 3 13 9 1 15 7 0 13
12 1 0 3 13 9 7 9 9 1 3 13 15
8 7 0 13 13 1 9 13 9
3 7 13 15
18 3 13 9 16 1 9 13 13 7 1 9 3 16 3 1 9 13 15
8 13 3 15 0 15 3 13 15
8 7 13 13 7 16 13 1 9
6 15 13 9 13 3 13
3 7 13 15
4 13 15 15 13
12 1 15 9 13 13 15 15 7 13 15 15 13
11 7 15 3 13 3 15 13 13 15 1 15
2 7 13
26 0 13 9 0 3 9 13 9 1 9 7 13 7 13 9 7 9 7 9 13 7 13 3 3 13 0
19 1 15 3 9 13 15 3 9 1 0 3 9 1 0 3 3 9 1 9
10 3 3 13 9 3 13 9 16 13 9
2 7 13
4 15 13 9 0
5 7 15 9 13 15
6 1 9 3 3 13 15
6 12 3 13 9 15 15
8 7 13 15 1 0 9 9 13
4 13 1 0 9
16 7 13 9 13 15 3 13 1 9 7 15 3 9 13 1 15
5 7 13 9 0 0
10 9 3 13 15 1 9 16 3 13 13
3 7 13 15
6 9 3 13 3 16 13
4 7 13 13 9
3 7 13 9
3 13 7 13
7 7 13 9 7 13 9 0
3 7 13 15
4 3 3 13 9
10 7 13 15 9 0 7 13 15 1 15
9 7 13 1 0 9 9 1 9 0
68 7 13 15 1 9 3 13 15 1 9 9 0 9 15 9 13 1 9 7 3 0 9 15 15 3 13 13 16 0 9 9 7 9 0 13 13 13 15 1 15 9 0 7 9 13 15 7 15 15 3 13 13 7 3 9 7 9 1 9 7 1 9 13 13 7 13 15 9
14 13 3 11 3 13 7 13 15 15 7 13 9 0 13
8 15 15 7 15 11 9 9 0
3 13 15 9
2 13 15
5 13 9 0 1 9
3 7 13 15
3 7 13 15
7 9 15 13 9 16 0 13
10 7 13 15 3 16 3 13 15 1 9
9 13 3 3 9 0 13 0 1 9
8 13 15 1 9 16 1 15 13
5 7 3 13 15 11
25 7 13 9 0 13 1 9 7 13 15 9 1 9 1 9 13 3 15 3 12 12 7 13 1 9
11 7 13 9 13 7 13 1 9 7 1 9
26 13 1 11 7 13 13 15 13 13 7 13 13 9 7 13 15 7 13 15 13 3 13 0 7 1 9
8 7 13 13 15 13 1 9 15
14 7 13 15 1 9 13 15 13 15 16 13 1 15 13
6 13 1 9 15 1 15
10 7 13 15 15 15 9 13 7 13 15
15 7 13 7 13 13 1 11 15 13 15 11 7 15 13 15
19 7 13 11 1 9 3 1 0 9 13 15 9 0 1 15 7 13 1 9
21 7 6 13 12 1 9 9 11 7 13 15 13 1 9 15 7 13 15 3 13 16
11 3 13 13 1 15 9 16 13 13 7 13
13 7 13 1 15 7 1 15 13 9 0 7 13 15
3 13 3 16
8 16 13 15 3 9 15 13 13
13 7 3 13 9 9 15 7 13 9 16 13 1 9
15 7 3 11 13 1 15 9 13 1 15 13 15 1 9 13
5 15 13 15 9 15
5 7 13 15 9 15
5 15 15 13 15 15
20 9 3 13 15 7 13 13 15 13 15 13 7 13 1 15 7 13 15 15 9
4 11 3 13 15
5 9 9 15 13 15
3 13 1 9
6 7 13 0 1 9 15
9 7 3 13 15 13 1 9 13 16
3 9 15 13
3 3 13 15
2 3 13
17 7 3 13 13 1 15 3 12 3 3 11 7 11 7 11 9 0
18 7 13 1 9 0 7 13 9 7 13 15 7 13 3 7 13 13 15
5 15 13 7 13 15
5 9 13 13 7 13
4 7 13 15 15
20 0 3 13 15 13 9 9 7 9 7 15 13 1 15 7 13 3 13 9 13
4 8 15 13 13
3 9 15 13
1 13
6 7 3 13 9 7 13
6 13 3 9 12 1 12
5 7 13 15 9 0
14 7 13 15 3 16 15 3 13 0 7 13 13 15 13
14 7 13 3 7 13 1 9 15 7 1 15 13 9 15
6 7 9 0 9 15 13
16 3 0 3 13 9 9 0 9 3 11 7 11 7 11 7 11
9 3 7 3 9 15 13 1 15 3
5 7 13 15 1 15
20 13 3 15 11 16 13 9 1 9 3 1 15 9 7 1 9 7 1 9 15
7 3 13 3 3 12 9 13
7 3 1 3 9 9 13 13
4 7 13 9 13
3 7 13 15
10 3 3 13 1 9 3 13 16 13 3
21 7 15 3 3 13 15 7 13 15 13 3 13 9 15 13 1 9 15 1 9 15
3 6 13 15
11 3 13 9 7 11 1 9 0 3 9 0
17 7 13 13 16 13 15 7 9 0 13 7 13 9 0 0 7 13
10 15 3 13 16 11 13 16 12 1 9
5 13 3 11 13 16
4 0 13 1 0
21 0 3 11 13 13 11 7 13 15 1 9 11 1 9 11 9 15 16 13 15 15
4 13 3 11 11
8 3 13 15 13 9 11 9 15
13 11 3 13 15 1 15 7 13 15 13 7 3 13
35 7 13 15 9 0 3 11 9 15 9 13 9 15 7 9 7 9 0 7 13 9 15 11 7 13 7 13 11 7 13 1 15 13 9 9
9 13 1 15 15 3 13 7 13 15
5 7 13 15 15 16
7 0 3 13 13 1 9 15
2 15 13
3 0 3 13
3 9 11 9
11 13 16 13 15 1 15 1 9 9 11 9
4 7 0 13 9
11 1 9 7 13 1 15 3 13 13 15 15
9 7 3 13 9 9 13 13 9 15
12 7 13 9 15 13 9 15 7 13 15 1 9
15 7 13 15 9 1 11 7 13 15 15 15 13 7 15 13
3 7 13 15
6 13 3 13 7 13 0
7 7 3 13 15 3 3 13
7 7 13 1 0 9 9 12
18 7 13 15 13 7 13 15 0 7 0 1 15 9 13 3 7 13 15
22 7 13 11 13 9 0 7 0 15 13 16 13 3 9 3 13 9 7 13 13 15 3
12 13 15 16 13 1 0 9 7 9 13 15 9
5 3 13 3 15 13
4 13 15 15 13
4 7 13 15 16
10 13 13 12 12 9 9 7 13 15 13
4 0 3 13 15
3 3 13 9
3 13 7 13
5 12 9 7 12 9
12 7 13 1 9 1 9 1 12 7 1 12 12
27 7 13 12 9 7 12 9 13 1 9 13 7 13 9 7 13 9 15 16 13 1 15 7 12 9 13 15
6 7 13 15 7 13 15
11 7 13 9 12 1 12 9 0 7 1 9
7 13 3 13 9 12 12 9
20 7 3 13 9 15 13 1 9 7 13 15 1 0 9 1 11 16 0 13 9
9 7 13 15 15 13 1 9 13 15
4 7 13 15 13
10 0 3 13 15 1 9 13 13 9 13
2 7 13
7 15 3 13 15 7 13 15
9 0 3 3 13 1 15 7 13 15
1 13
2 15 13
3 3 13 15
10 7 3 3 1 15 13 15 7 13 15
10 3 13 3 1 9 7 13 9 15 13
8 7 13 13 1 9 0 7 13
25 13 3 15 1 9 3 13 15 7 13 15 9 0 7 13 13 1 9 13 3 13 15 16 3 13
26 7 3 3 13 1 9 7 1 9 7 1 9 1 9 13 0 7 13 15 16 3 9 9 15 13 15
8 7 15 3 13 15 15 13 13
13 7 13 15 1 15 9 7 15 1 9 13 1 11
14 7 13 15 1 9 15 0 9 3 3 13 13 9 13
15 1 15 3 13 9 15 1 9 9 7 3 13 9 13 9
6 0 3 13 13 15 16
9 3 13 11 1 15 9 3 13 13
12 0 9 9 15 13 7 9 15 3 13 1 15
8 3 3 13 15 13 9 9 0
17 13 3 9 0 13 9 0 9 9 7 9 7 15 0 0 0 13
3 7 13 15
3 11 3 13
9 7 15 13 9 7 9 9 3 13
3 15 3 13
37 16 13 9 9 7 9 9 15 13 9 7 15 3 1 15 13 13 3 1 0 3 13 15 15 13 9 15 7 9 15 13 9 0 9 15 15 13
5 7 0 0 0 13
6 7 13 15 9 13 15
5 13 15 15 7 13
8 7 13 1 15 0 13 13 9
7 16 15 13 9 13 3 13
3 7 13 15
6 3 3 3 15 0 13
30 3 13 3 16 0 15 3 13 1 9 3 13 15 13 16 3 13 15 1 9 7 1 9 7 1 9 13 13 15 9
9 13 3 16 13 1 9 0 13 9
20 3 3 1 9 0 9 13 9 9 9 9 9 9 9 9 9 0 9 9 9
25 7 3 13 13 1 9 0 7 0 7 1 9 13 3 13 16 13 15 15 13 7 3 13 13 15
15 13 3 9 1 15 15 9 13 9 0 13 13 1 9 15
6 9 3 13 9 9 9
4 11 3 13 15
6 13 16 3 13 15 9
9 13 3 0 13 9 9 7 9 13
7 0 3 13 13 15 6 9
3 7 13 15
4 1 9 0 13
5 13 9 1 9 15
11 7 13 3 13 9 13 1 9 7 9 13
14 7 13 1 15 0 0 7 13 15 16 13 1 15 9
26 7 13 15 12 1 9 13 9 15 1 9 15 7 13 13 15 1 9 7 13 1 9 13 7 13 15
5 8 15 13 13 15
7 7 13 15 16 15 3 13
8 3 15 0 13 0 3 3 13
5 7 3 13 15 13
3 3 15 13
6 0 13 13 7 0 13
16 0 15 13 9 0 16 3 12 9 13 15 7 3 13 15 13
12 7 16 13 15 3 13 1 9 15 13 1 9
5 7 13 15 9 15
9 3 0 13 15 3 13 9 1 9
3 7 13 15
3 3 13 9
3 0 3 13
1 12
4 7 13 1 9
4 7 0 13 13
3 13 3 0
11 13 3 7 13 15 7 13 9 9 12 9
6 13 3 13 3 12 12
3 7 13 15
12 7 3 13 1 9 1 9 15 13 1 9 0
17 7 13 9 7 13 13 15 1 15 13 1 15 9 1 9 13 15
3 6 13 15
6 3 13 15 9 0 9
11 7 13 15 13 3 1 9 13 1 0 9
14 7 13 13 9 7 1 12 9 3 13 1 15 1 9
4 7 13 15 13
1 13
9 13 15 1 9 0 7 1 9 0
7 7 13 15 1 15 13 16
5 7 13 11 13 15
6 15 13 16 9 3 13
7 3 3 3 13 7 13 3
5 13 3 13 9 15
25 9 13 3 13 7 9 13 3 13 7 3 13 3 3 12 9 13 1 12 12 7 3 9 9 13
2 13 15
3 12 1 12
11 7 3 12 1 12 12 3 9 9 9 13
3 7 13 15
3 3 3 13
4 7 13 1 11
11 7 13 1 15 0 7 13 15 16 15 13
25 7 13 1 9 0 13 15 3 1 9 7 13 1 9 15 7 13 9 1 15 13 15 16 15 13
3 7 13 13
1 13
20 1 0 3 3 13 9 1 9 15 7 13 15 13 7 13 15 7 13 15 3
9 7 1 9 13 7 13 15 1 9
10 13 3 11 7 9 15 1 9 11 0
8 7 1 9 13 9 15 13 15
5 15 15 13 9 13
3 0 3 13
11 0 11 9 7 15 11 7 0 12 1 9
6 15 3 15 15 13 13
5 13 3 11 13 15
9 7 13 15 16 15 3 13 1 15
26 7 13 13 15 16 13 9 0 3 13 7 13 13 1 9 7 9 7 9 7 13 13 7 0 9 13
6 7 3 13 15 9 13
7 7 13 15 11 13 13 15
12 0 3 13 15 7 13 1 9 15 13 11 13
8 7 13 9 1 9 15 13 15
17 15 13 1 15 13 3 13 15 15 7 13 9 15 7 13 1 15
9 15 3 3 13 9 15 13 13 15
13 15 3 9 13 9 16 13 15 9 7 13 9 15
8 15 3 13 9 9 1 9 15
30 15 3 3 13 15 15 7 15 9 1 9 0 0 7 0 3 9 0 13 15 15 3 13 1 9 9 15 1 9 0
21 6 13 15 16 13 15 1 3 13 15 3 13 13 9 16 13 9 0 13 1 9
12 7 13 15 15 11 1 11 7 13 13 1 11
5 7 13 11 13 11
18 9 0 13 15 3 13 7 13 12 9 15 12 7 11 12 7 11 12
5 3 13 3 15 13
11 7 13 3 9 13 15 7 13 9 1 9
5 0 13 9 15 13
2 13 15
20 13 3 15 1 9 13 15 16 15 3 13 15 13 3 3 9 0 13 1 0
13 7 13 9 1 15 13 15 15 13 10 1 0 13
8 7 13 15 13 3 13 9 16
4 11 13 3 13
5 0 3 13 13 15
7 7 3 13 13 1 9 0
6 16 3 13 7 13 15
15 7 13 1 9 13 9 0 1 15 7 9 13 15 1 15
12 7 3 15 9 13 15 13 15 7 13 13 15
3 7 13 9
5 15 13 15 1 15
6 7 13 12 1 9 13
17 9 13 9 15 1 15 13 9 0 7 15 3 3 13 15 13 15
10 7 13 9 15 16 13 15 7 3 13
7 6 9 0 3 1 15 13
3 3 13 15
4 13 15 1 15
5 7 13 15 1 15
15 7 13 15 9 3 13 15 7 13 1 9 13 15 9 13
5 7 13 11 9 15
7 3 9 13 3 0 13 15
13 7 3 7 1 9 13 7 1 9 16 15 13 13
9 7 16 15 13 13 15 13 1 15
8 11 3 13 15 10 16 13 13
3 15 0 13
8 7 3 13 9 9 1 9 13
1 13
4 9 13 15 9
12 13 3 11 16 13 15 9 13 9 0 13 15
7 7 13 7 3 13 15 13
9 7 13 3 0 16 0 13 16 13
9 11 3 13 15 1 9 13 7 13
11 7 13 15 1 9 9 15 13 15 12 16
5 15 3 13 13 15
3 7 13 15
10 0 9 15 3 13 13 3 9 7 9
12 7 3 13 13 1 11 7 3 13 16 15 13
10 7 13 1 11 7 1 9 13 13 15
6 15 1 9 1 15 13
3 0 3 13
10 15 1 15 3 13 1 9 15 13 0
9 7 13 13 12 1 12 7 13 15
12 16 15 13 0 13 3 13 15 0 7 15 9
13 7 13 9 13 15 1 9 15 7 13 15 13 15
11 7 15 3 15 13 3 15 13 7 13 15
19 9 13 15 9 15 13 9 15 3 13 1 15 7 13 15 16 3 13 15
3 11 3 13
3 3 13 15
14 15 3 13 15 13 9 1 9 15 7 13 3 13 15
8 15 3 13 1 15 1 15 13
19 15 3 3 13 15 9 9 1 9 16 0 13 6 13 15 3 13 9 15
8 7 16 13 15 9 15 13 15
26 0 15 13 9 1 9 13 3 12 9 13 13 1 9 1 9 0 3 9 15 3 13 7 9 3 13
27 0 15 13 13 1 9 0 3 12 9 13 13 13 1 9 1 9 0 3 9 15 3 13 7 9 3 13
8 7 16 9 15 13 15 13 15
27 0 15 13 1 12 9 13 1 9 0 3 12 9 13 13 1 9 0 3 9 15 3 13 7 9 3 13
11 0 3 9 13 15 7 0 9 9 13 15
3 0 13 9
9 13 9 1 15 7 9 13 1 15
24 7 3 13 13 1 9 0 1 0 9 11 7 13 3 9 1 15 7 3 13 9 3 13 15
12 7 13 9 13 15 16 13 9 9 13 13 15
4 15 15 13 11
7 13 11 9 0 13 7 13
5 7 13 11 13 15
7 1 9 15 13 15 9 0
20 0 1 13 9 9 15 7 9 7 13 15 1 9 15 7 13 12 1 9 12
8 0 3 3 13 12 7 9 12
9 15 3 9 13 13 9 3 3 13
10 7 1 9 3 9 15 1 0 13 15
13 15 3 13 9 15 7 13 15 15 9 13 1 15
10 7 16 9 13 9 13 1 15 9 13
8 7 13 1 15 9 16 15 13
4 13 3 11 13
3 7 13 15
10 3 13 9 13 1 15 7 3 13 15
5 0 3 13 9 0
3 6 13 15
8 7 13 15 13 13 9 1 15
15 7 13 15 1 9 13 15 7 13 15 15 1 9 13 15
4 11 3 13 15
4 15 15 13 0
5 15 0 3 12 9
2 9 13
3 3 9 13
2 3 13
3 3 13 13
5 13 9 15 7 9
5 0 3 13 13 15
7 9 15 0 13 1 9 15
10 11 3 13 1 15 13 15 7 13 15
3 12 13 13
25 16 13 13 13 13 15 13 13 7 13 0 7 13 13 9 1 9 7 13 13 1 9 15 13 9
8 0 3 0 13 1 9 13 13
8 3 3 13 9 1 9 0 13
7 9 3 13 15 1 9 15
6 11 3 3 13 13 15
11 9 3 3 13 13 1 9 1 9 0 13
13 0 13 9 1 0 9 13 3 0 1 9 0 13
8 0 3 3 13 15 13 1 15
4 15 13 13 13
6 7 13 1 15 11 13
6 15 3 0 1 9 13
5 13 3 11 13 15
9 6 15 13 15 7 1 9 15 13
4 13 3 11 13
3 6 13 15
53 15 13 15 13 9 7 9 7 9 7 9 7 9 7 9 7 9 7 9 15 1 7 9 16 3 13 13 3 1 9 0 3 9 7 9 7 9 7 9 7 9 7 9 7 9 1 9 7 1 9 13 9 0
8 0 3 13 0 0 7 0 0
34 13 3 1 9 13 1 11 7 13 13 11 7 13 15 7 3 13 13 15 7 13 11 3 12 1 12 13 15 13 15 13 13 15 16
8 9 13 16 15 3 13 13 15
4 11 3 13 15
5 15 13 16 13 15
4 0 3 13 15
16 13 15 16 12 1 0 15 7 12 1 0 15 13 1 9 15
4 11 3 13 15
5 3 13 15 15 13
4 0 3 13 15
4 11 3 13 15
6 9 3 15 15 13 13
8 7 9 15 15 13 15 13 15
16 7 10 13 1 0 15 7 1 0 13 15 13 7 15 13 13
9 7 13 12 13 13 1 11 7 11
6 11 3 13 15 13 15
6 3 3 3 13 1 15
24 7 15 3 13 0 13 1 15 3 13 15 9 7 15 3 13 1 15 13 0 3 13 15 9
4 7 13 1 11
18 13 15 1 11 7 9 15 7 9 0 9 0 11 0 13 1 9 13
10 7 13 16 11 9 13 13 13 7 13
5 9 0 11 13 15
6 7 13 15 0 16 13
4 9 0 13 15
6 7 13 11 13 13 15
5 7 13 9 13 15
1 13
2 13 15
9 0 3 13 9 15 13 13 1 11
5 7 13 13 15 11
4 9 3 13 15
3 9 3 13
4 11 3 13 15
1 13
9 7 3 13 7 1 11 13 1 9
21 7 3 13 15 1 11 1 11 7 11 1 9 0 13 12 1 9 15 7 13 15
24 13 1 9 15 13 1 15 7 3 13 1 15 13 9 13 1 15 13 3 3 15 1 9 13
18 7 16 15 15 13 15 0 13 13 16 9 15 13 7 3 13 15 3
14 13 3 7 13 9 13 1 9 3 1 9 7 13 15
7 7 15 1 13 3 13 15
4 15 13 13 9
7 0 3 13 15 3 13 11
15 7 13 9 1 11 7 13 1 15 9 15 7 13 1 15
17 0 3 9 15 13 1 9 7 0 9 13 1 9 7 13 1 9
6 6 0 13 1 9 0
12 0 13 9 1 9 9 9 15 11 6 1 0
8 7 13 1 11 11 7 1 9
3 7 13 15
11 3 3 13 9 13 1 11 1 12 1 12
8 7 1 0 13 15 1 11 13
5 3 13 3 9 9
10 1 0 1 15 1 9 15 9 3 13
4 13 3 9 15
24 7 13 1 11 7 13 11 1 9 13 13 13 7 13 1 9 7 9 9 7 9 13 9 13
12 7 3 13 15 13 9 1 9 7 13 13 15
4 13 3 13 16
8 9 15 9 9 13 15 15 9
6 15 3 13 15 9 9
8 7 16 3 13 13 3 1 9
8 7 13 3 13 9 13 1 9
5 7 13 11 13 15
2 9 13
4 9 15 13 13
5 7 13 11 13 15
3 13 9 0
34 6 13 15 16 15 13 9 0 13 15 7 13 15 1 9 7 3 13 15 1 9 15 7 9 13 16 15 13 13 13 15 15 3 13
11 15 15 13 15 13 13 16 13 7 13 15
20 7 3 13 13 15 13 16 15 13 1 15 16 3 9 15 0 13 15 9 15
14 16 3 15 3 13 3 9 15 15 1 9 13 9 15
5 7 13 3 1 11
13 7 1 9 13 15 13 1 15 9 7 9 7 9
3 7 13 15
13 15 9 0 13 7 15 15 13 9 0 16 0 13
5 11 3 13 13 15
2 13 15
5 7 13 1 15 13
11 16 13 1 9 13 1 15 3 3 13 15
4 16 13 1 9
3 13 15 9
6 15 3 13 11 3 9
4 7 13 13 11
8 3 15 13 15 15 9 0 13
19 9 9 13 7 13 15 9 7 13 9 7 13 9 7 13 15 9 7 13
14 7 13 1 9 9 1 9 16 1 9 13 1 9 9
8 0 3 13 15 13 7 13 0
7 7 3 13 1 15 0 9
10 7 0 9 13 13 9 15 7 13 0
7 7 3 15 13 7 0 13
7 3 3 13 12 9 13 15
8 13 3 0 1 15 3 13 16
10 0 3 9 1 15 13 16 0 13 9
1 13
2 13 15
4 7 15 13 9
10 7 13 13 15 7 13 15 3 1 9
4 13 7 13 9
4 7 13 9 15
6 3 3 0 13 9 13
10 1 9 13 0 7 13 0 1 9 15
8 7 13 13 15 7 13 15 9
7 13 3 16 1 15 13 9
4 7 13 15 13
6 0 3 13 13 15 9
10 13 16 0 13 7 3 13 3 1 15
12 3 13 3 1 9 9 7 1 9 9 0 13
7 13 3 13 9 9 7 3
7 0 3 13 15 9 13 15
3 15 15 13
5 13 15 9 16 13
6 15 13 9 0 7 9
4 0 3 13 15
1 0
5 7 13 11 13 15
6 0 13 9 7 0 9
14 7 13 9 1 15 15 13 3 13 9 7 13 15 13
26 9 11 13 15 16 16 15 9 13 7 13 9 7 9 3 13 3 13 9 9 15 7 13 9 9 15
9 7 0 13 9 7 13 3 13 9
11 7 0 13 15 7 13 7 0 3 13 9
3 7 0 3
8 7 13 15 12 7 3 13 9
6 1 3 15 13 3 9
9 1 9 3 3 13 15 15 13 9
5 7 13 11 13 15
16 3 3 1 0 13 7 13 15 7 13 7 13 3 9 1 9
18 7 1 0 16 13 13 3 13 1 9 0 1 9 3 13 15 9 13
9 15 9 0 7 9 0 7 9 0
6 13 9 0 7 9 0
4 15 3 3 13
16 7 13 15 1 9 13 15 13 15 13 16 3 13 15 13 15
5 15 13 9 0 15
2 13 11
6 9 9 15 9 12 13
20 7 13 9 9 15 15 9 15 7 15 9 15 7 15 9 15 7 15 9 15
4 0 0 15 9
4 7 0 0 15
6 13 0 15 3 0 15
5 0 0 15 9 13
4 7 13 15 9
27 7 10 13 15 15 9 7 15 9 7 15 9 7 15 9 7 15 13 0 3 15 0 13 15 9 7 9
9 11 3 13 15 16 3 13 13 15
6 3 3 13 1 9 0
8 7 15 3 13 15 1 0 13
7 7 13 11 13 13 1 9
8 3 13 9 16 11 9 0 13
6 0 3 13 11 9 0
4 13 9 9 15
5 7 3 15 13 9
7 7 0 9 13 15 1 9
6 7 13 15 1 9 15
32 13 15 1 9 13 1 9 13 7 9 1 9 7 9 1 9 7 9 1 9 13 9 9 7 9 3 13 15 0 13 0 9
12 7 13 11 1 9 13 3 9 13 9 1 9
5 7 0 0 13 0
11 7 13 15 9 0 13 12 9 15 13 9
13 6 13 15 16 9 0 0 3 15 13 13 1 9
11 7 13 15 1 9 13 15 15 1 9 15
7 9 13 0 9 7 0 9
5 11 3 13 13 15
5 13 3 0 0 9
12 3 13 13 3 9 1 9 15 3 13 13 15
18 7 13 15 1 9 0 1 9 13 15 12 11 7 11 7 11 7 11
6 11 3 13 13 13 15
7 13 15 16 3 15 13 15
10 3 3 13 9 7 9 9 3 13 15
7 13 3 13 7 3 3 9
19 13 3 9 1 9 7 9 1 9 7 13 9 1 9 7 13 9 7 9
3 9 9 0
5 13 3 15 15 0
17 7 1 9 13 13 7 1 9 7 1 9 13 15 1 1 9 15
9 7 1 15 9 13 3 13 15 9
25 3 3 13 15 13 3 13 15 3 15 13 7 13 15 7 15 3 13 15 15 1 0 9 0 13
17 13 3 9 9 1 9 7 9 9 7 13 9 1 9 7 13 15
7 7 13 13 15 9 15 1
7 13 3 1 9 0 13 13
53 3 3 9 13 9 13 11 9 13 3 3 13 13 3 13 3 15 13 1 11 3 13 1 9 7 15 1 9 3 3 13 1 9 7 3 13 13 15 1 9 15 7 13 1 9 3 3 13 15 3 13 9 15
9 13 3 15 16 3 13 9 15 9
20 13 3 9 0 0 3 3 13 0 1 9 9 15 13 9 1 3 7 3 13
13 7 16 3 13 9 13 9 3 13 13 13 0 9
7 7 13 1 15 13 13 9
17 13 3 0 11 7 0 9 7 13 9 7 9 16 13 16 0 13
4 15 3 13 15
5 6 3 13 15 15
13 7 3 13 9 0 13 1 9 1 9 0 7 9
18 7 3 13 9 15 7 13 13 15 1 12 9 1 9 9 1 9 9
5 1 9 3 13 9
14 3 3 9 15 13 0 7 13 9 13 16 1 13 9
13 3 3 15 3 13 0 13 13 16 1 13 1 9
9 9 7 9 13 7 15 9 3 13
20 7 1 9 0 7 1 9 15 3 13 7 9 15 13 1 9 7 9 3 9
6 3 13 3 3 9 13
22 3 9 13 13 9 15 7 13 9 15 9 7 15 9 15 7 9 13 16 13 13 3
17 3 13 3 3 9 9 13 3 3 1 9 9 3 1 9 3 3
7 16 3 13 3 13 15 13
6 7 15 15 13 15 13
1 13
10 7 13 9 7 9 3 15 9 13 13
4 7 3 1 9
5 3 3 13 9 9
19 7 13 15 1 11 1 9 11 0 13 15 13 9 13 9 9 0 9 0
7 7 13 9 13 15 1 9
8 13 3 15 13 1 15 7 13
6 1 15 9 0 0 13
14 13 3 0 9 13 13 3 12 12 9 7 13 15 0
2 13 15
4 1 15 15 13
6 0 3 9 13 1 15
18 3 3 0 13 1 15 7 3 13 13 15 0 13 7 15 3 3 13
4 15 13 0 13
7 13 13 13 9 15 1 9
3 6 13 15
18 3 3 13 13 9 0 1 15 9 3 15 13 0 13 13 1 9 15
10 0 3 13 13 15 7 13 15 9 13
8 7 13 3 15 1 0 9 13
12 7 1 0 9 9 3 9 13 13 15 9 15
7 3 13 13 13 16 13 9
6 7 13 12 1 9 15
3 7 13 15
11 13 1 9 7 13 15 9 1 9 9 13
3 1 15 13
9 3 13 9 3 9 1 9 15 13
8 7 0 15 13 9 0 13 0
3 3 13 15
16 7 13 9 15 7 13 1 9 7 13 3 13 15 7 13 9
8 7 9 13 13 1 12 1 12
7 7 13 15 7 13 13 11
12 6 13 15 16 15 1 15 13 15 13 1 15
2 3 15
2 3 15
5 0 3 13 13 15
10 12 1 12 1 12 13 1 15 1 9
10 9 3 3 0 13 3 13 13 1 15
9 6 3 9 0 15 9 0 13 15
11 0 13 15 13 16 3 13 13 15 9 0
5 7 13 15 7 13
1 13
12 7 13 9 9 13 13 15 7 13 1 15 15
3 7 13 15
9 0 13 9 15 0 9 13 1 0
21 6 3 13 15 16 3 3 13 13 1 9 0 1 0 9 3 13 15 1 9 0
6 7 13 13 1 9 0
8 15 13 15 1 15 1 0 9
3 13 3 13
6 13 9 7 9 13 15
4 11 3 13 15
8 3 16 15 13 15 7 3 15
4 7 13 15 11
4 6 13 15 16
5 0 3 3 13 3
11 16 15 15 13 1 15 13 3 13 15 15
4 3 3 15 13
10 13 1 9 15 9 11 7 13 9 15
18 7 13 11 7 11 7 11 1 15 7 13 13 15 7 13 7 13 15
6 0 13 9 15 1 9
4 13 3 7 13
6 9 9 15 0 15 13
5 13 9 0 1 15
8 7 3 3 15 13 7 15 0
9 7 13 7 13 15 13 7 13 11
3 11 13 3
9 13 7 13 15 16 3 13 1 9
7 9 3 13 0 7 9 0
7 7 13 15 13 15 3 13
12 13 3 15 9 0 7 3 13 15 13 13 15
3 7 13 3
3 7 13 15
4 13 3 7 13
2 13 9
8 6 13 15 9 0 1 9 9
1 13
5 6 13 15 13 15
27 7 3 3 15 13 13 11 12 1 12 1 12 7 1 15 9 0 1 9 7 9 1 9 7 9 7 9
7 13 3 13 15 9 15 13
7 15 3 13 13 7 0 13
3 7 13 3
7 7 13 3 13 1 15 13
9 0 3 13 9 1 15 7 13 15
13 12 3 1 13 13 9 13 9 0 7 13 15 9
5 7 13 11 13 15
11 3 1 9 3 13 1 9 7 9 13 15
13 1 15 9 13 1 15 13 1 9 7 3 13 15
5 7 3 13 15 9
5 7 13 15 15 13
15 7 12 9 15 1 15 13 13 1 9 0 7 13 3 9
16 7 13 11 1 9 7 13 15 1 15 15 9 7 9 7 9
22 7 11 3 1 9 15 13 1 3 1 9 0 7 13 13 1 9 7 13 15 1 9
15 9 3 7 15 9 13 1 11 9 16 15 13 7 3 13
19 0 3 13 1 15 7 3 13 0 9 7 15 13 9 13 1 15 13 16
5 15 13 15 13 16
11 15 13 9 0 0 7 12 9 15 0 13
8 7 3 3 3 13 0 9 15
8 7 13 9 1 9 13 11 13
7 0 3 13 7 15 3 13
7 3 9 13 15 7 13 15
6 15 3 13 11 9 0
3 11 3 13
2 15 13
13 7 13 9 0 1 0 13 9 7 13 1 9 0
6 9 3 13 9 15 13
3 13 9 15
8 0 3 15 13 15 0 13 9
16 7 13 15 13 1 15 7 13 9 15 7 13 15 7 13 15
7 13 15 11 15 13 13 15
7 7 9 13 1 9 13 15
20 7 13 11 3 1 9 13 12 1 9 0 7 13 11 13 15 13 1 15 13
6 3 15 1 9 11 13
7 3 13 7 13 15 15 13
8 7 13 3 1 9 7 9 13
4 0 13 1 15
5 0 3 3 13 15
8 7 3 1 0 3 13 13 11
5 1 9 1 15 13
3 3 9 13
9 0 3 13 13 15 7 13 15 16
6 3 13 9 0 15 13
12 7 3 9 13 7 13 11 9 15 13 15 11
4 7 13 13 15
21 7 3 1 0 9 13 9 7 9 7 9 7 15 9 13 11 13 7 13 15 11
4 7 13 15 11
5 15 3 13 9 0
2 15 13
6 7 13 1 15 9 3
5 0 3 15 3 13
6 11 3 3 13 15 13
5 13 3 1 15 13
11 11 3 1 0 15 3 13 16 13 15 11
10 1 0 3 9 13 15 12 9 15 13
8 7 13 13 13 3 3 13 15
5 11 3 13 15 13
7 13 3 16 13 15 9 0
8 13 3 16 9 1 13 15 9
9 9 3 13 9 16 3 11 13 15
8 15 3 13 13 15 13 9 0
4 0 3 3 13
4 11 3 13 15
4 15 3 0 13
4 0 3 3 13
2 13 15
16 11 3 13 9 9 13 13 15 11 7 13 11 13 16 15 13
14 9 3 13 11 3 1 9 15 13 9 7 13 15 9
4 7 13 13 15
16 7 13 15 9 1 9 7 13 1 15 7 13 9 13 15 15
15 7 3 13 15 15 13 1 15 9 7 13 15 1 9 15
6 7 13 15 16 13 15
17 7 13 13 15 11 11 13 1 9 9 0 7 0 16 13 9 15
11 7 13 15 1 9 11 15 13 13 0 9
6 7 13 15 13 0 9
4 0 3 3 13
8 7 13 9 9 15 13 9 0
20 7 1 15 13 12 9 12 1 0 7 0 1 0 15 7 13 15 13 15 13
5 7 1 9 13 13
10 7 13 13 15 7 13 9 15 7 13
14 6 13 9 7 12 9 13 13 15 0 7 13 1 9
11 3 3 9 13 15 1 9 15 1 15 13
7 15 13 7 15 3 13 13
13 11 9 0 3 13 3 1 9 16 13 7 9 13
12 13 3 9 0 9 13 1 15 9 1 0 9
9 7 1 0 9 13 11 9 0 13
4 8 8 8 8
3 15 13 13
6 9 9 15 3 15 13
6 7 15 1 13 13 13
1 13
2 11 13
6 11 3 13 9 0 13
11 7 9 0 13 15 1 12 1 3 1 3
11 13 3 9 13 1 15 16 3 13 13 13
7 1 9 9 0 9 0 13
40 13 3 7 9 3 13 1 15 13 7 11 9 7 11 11 0 7 9 0 7 11 15 3 13 1 11 1 15 13 7 13 15 7 15 0 13 1 15 1 11
34 7 3 3 13 16 13 9 9 15 13 1 9 13 11 1 11 0 9 15 3 0 13 13 9 0 7 13 13 1 11 7 13 9 0
7 11 3 13 15 16 3 13
7 7 13 1 9 13 9 11
10 11 3 9 7 11 0 13 3 15 13
16 7 13 9 11 9 7 11 0 7 11 13 9 16 13 13 15
11 7 3 3 1 12 9 13 1 9 13 9
4 7 13 1 15
7 15 13 15 9 1 9 9
7 7 13 13 16 13 13 9
16 7 13 1 9 13 9 13 1 0 13 1 9 0 7 13 15
4 0 3 13 15
4 11 13 9 13
1 13
2 13 3
5 6 9 3 13 13
2 7 13
6 3 15 13 3 13 15
5 7 13 13 1 9
15 7 13 3 15 9 7 9 7 15 15 3 13 13 3 15
10 0 13 13 13 1 15 13 15 7 13
13 0 3 13 16 0 13 7 13 13 15 3 13 9
14 1 0 3 12 1 15 13 13 15 15 9 13 1 9
5 7 0 13 13 0
24 3 3 13 15 12 1 12 13 15 7 13 9 15 7 9 16 13 15 13 1 0 3 13 9
3 7 13 15
8 13 1 15 9 13 9 15 9
16 7 15 9 13 7 13 15 13 13 7 15 3 13 9 13 13
28 9 15 9 13 9 13 0 7 1 9 9 13 16 3 0 15 13 15 15 3 13 1 9 9 13 7 0 13
17 9 3 11 1 9 15 1 15 13 15 1 9 7 13 1 0 9
12 0 3 13 13 3 9 13 7 9 13 13 9
45 16 3 0 13 13 9 1 13 1 15 9 3 13 15 13 3 9 7 9 9 13 15 3 15 13 3 1 15 1 9 1 9 13 15 0 11 16 13 1 15 13 15 13 9 9
23 13 1 9 11 9 0 9 15 9 11 1 9 0 7 9 15 1 9 0 7 9 15 11
15 13 3 12 0 1 9 13 1 9 15 7 9 0 1 9
16 7 3 13 15 9 16 13 11 9 7 12 13 1 9 15 13
32 13 3 13 15 1 9 9 15 1 9 1 9 0 13 15 15 13 13 1 9 0 7 15 9 9 13 9 13 3 1 9 9
10 7 13 15 11 13 7 9 13 1 15
5 13 3 1 15 9
13 7 13 15 9 7 9 7 0 1 9 15 13 15
31 13 3 0 1 9 7 9 7 9 3 13 13 7 9 0 13 15 3 1 9 9 15 7 0 9 0 13 1 9 9 15
23 7 0 13 1 15 9 7 9 0 13 9 9 1 9 7 0 1 9 0 13 9 9 0
5 7 13 11 1 9
4 1 15 13 0
11 15 3 13 0 7 9 15 13 1 9 15
15 15 13 11 13 1 9 7 13 13 13 1 15 7 13 15
13 7 13 9 13 11 7 13 15 16 13 0 1 9
14 13 3 3 13 13 1 9 7 13 16 9 13 1 9
8 7 0 13 13 15 7 13 0
12 7 13 16 13 15 9 9 15 13 1 9 15
8 1 0 3 9 13 11 9 15
7 7 13 15 12 9 13 16
14 3 13 15 9 1 9 1 15 13 13 9 15 1 9
2 13 15
4 0 9 1 15
4 0 15 1 9
12 0 3 13 13 15 1 9 15 7 13 1 15
4 15 0 13 9
4 7 13 15 9
4 3 13 15 11
5 13 3 9 1 9
31 0 13 0 7 9 0 13 15 7 13 15 9 9 9 11 9 15 7 13 15 1 9 0 1 9 7 9 15 3 13 9
5 13 3 11 1 9
3 3 13 0
4 3 9 3 13
5 7 13 9 13 15
10 9 0 13 1 15 7 9 0 13 15
10 0 3 15 13 15 0 13 15 9 0
27 7 6 11 9 15 3 0 13 9 1 9 15 7 0 9 0 13 15 13 9 16 3 13 1 9 0 9
5 13 15 1 9 15
5 7 13 1 15 9
22 13 3 11 1 0 9 13 1 9 1 9 1 9 0 7 13 1 9 0 7 13 11
13 7 13 16 13 11 9 0 13 15 9 1 9 15
6 7 13 15 9 0 11
6 7 13 9 0 7 13
9 0 15 1 9 7 0 9 9 15
17 6 3 16 13 9 9 15 1 9 15 13 15 9 9 1 9 15
3 7 13 11
4 13 9 15 9
15 7 13 15 9 15 1 9 9 15 16 13 1 9 9 15
12 6 3 3 13 15 15 9 16 13 15 9 0
4 7 0 9 15
10 7 9 15 1 9 7 9 13 15 15
5 13 0 9 9 15
7 13 0 1 9 7 13 0
17 13 11 9 15 13 9 3 13 1 9 15 11 7 9 15 1 9
15 13 3 11 1 15 3 3 12 9 7 13 15 1 9 15
10 11 3 13 15 9 13 15 7 13 9
20 7 13 3 13 7 9 15 16 13 13 9 9 15 1 15 7 13 15 1 15
15 7 13 1 0 9 13 13 9 7 13 15 9 9 15 11
6 6 7 3 13 15 11
4 7 13 15 16
10 15 13 1 9 15 15 13 15 9 0
5 7 13 9 13 13
4 11 13 9 15
4 7 13 15 15
13 13 3 15 9 15 3 7 9 15 7 13 13 9
5 15 3 9 0 13
6 7 9 0 13 1 15
11 7 11 9 15 13 15 9 0 7 13 13
78 0 9 9 0 16 13 7 13 9 9 15 7 13 9 9 15 1 9 11 9 15 3 13 9 0 13 1 9 9 9 1 9 15 7 1 9 15 13 15 13 9 1 9 15 7 13 9 0 15 9 15 13 15 1 11 9 15 13 15 1 9 1 9 9 15 13 15 13 15 9 7 9 1 15 15 9 9 15
42 13 3 1 9 0 13 9 15 13 9 9 9 15 1 9 9 15 9 1 9 15 1 15 13 13 15 9 1 3 13 13 1 9 7 9 0 13 9 15 1 9 0
17 9 3 13 7 13 15 9 7 13 1 9 1 9 9 15 1 11
13 13 3 1 9 0 13 9 1 9 11 13 15 9
9 7 13 15 15 13 15 1 15 9
33 13 3 11 1 11 1 9 0 1 11 1 9 0 15 13 15 11 16 13 1 9 7 9 0 13 15 1 11 13 15 9 13 0
30 13 3 3 13 3 13 15 9 13 15 7 13 9 15 9 7 13 15 7 13 15 1 9 16 3 13 15 9 1 9
14 7 13 9 1 0 9 13 7 13 9 0 1 9 15
17 7 6 9 0 13 1 15 7 9 0 13 15 7 13 15 9 0
3 3 13 15
23 6 3 13 15 9 0 15 13 15 9 16 13 15 15 3 9 15 13 11 9 1 9 0
6 13 9 13 13 1 9
12 7 3 13 1 9 9 9 0 13 9 7 13
11 9 1 0 9 7 1 9 9 1 9 9
16 7 13 16 13 1 15 9 1 9 7 9 9 13 15 1 15
13 13 3 1 11 7 13 9 0 13 15 13 15 9
15 7 13 13 15 7 13 11 3 7 11 7 9 13 1 9
11 7 15 13 13 15 1 13 1 9 1 15
19 7 13 15 9 13 7 13 9 1 15 15 13 7 13 3 13 13 1 15
23 7 3 13 15 12 9 16 15 13 7 13 9 15 11 13 9 3 16 3 13 15 1 9
48 7 3 13 15 9 9 15 1 9 0 13 15 1 11 13 1 9 3 13 13 1 9 0 16 0 9 0 9 13 9 0 9 13 15 7 13 9 1 13 1 9 0 12 9 7 12 9 0
24 7 6 13 9 1 11 15 9 11 7 9 0 0 7 0 13 9 0 7 9 13 0 1 15
14 7 13 15 13 9 0 3 13 9 3 16 13 11 0
5 7 13 9 1 9
25 7 3 13 9 9 11 13 15 1 9 0 1 15 7 0 13 15 1 9 15 7 13 9 7 13
10 7 13 15 11 7 13 1 11 9 15
15 6 13 0 1 9 7 1 9 0 1 11 7 1 9 0
14 7 15 3 0 9 13 9 16 13 15 1 0 9 9
9 7 13 11 9 9 0 1 9 0
13 0 13 1 9 0 13 1 9 12 9 1 9 15
19 7 0 9 1 12 12 7 12 9 15 3 13 9 7 9 13 9 7 9
18 7 0 1 0 9 13 13 15 9 7 13 1 15 15 13 9 1 11
15 16 13 15 15 1 9 9 13 15 1 11 1 9 15 11
12 7 13 9 15 1 15 9 1 11 1 9 9
32 7 3 13 12 1 12 9 13 15 1 11 1 9 9 7 13 9 13 15 15 13 9 11 1 11 7 3 13 11 7 9 15
27 13 3 15 1 9 13 13 12 9 7 13 15 1 9 7 1 9 7 3 13 15 13 15 1 11 13 15
19 7 13 1 12 9 13 15 1 9 13 1 9 9 7 13 15 7 13 15
12 13 3 15 15 13 15 1 9 7 1 9 15
11 7 13 15 13 15 7 13 1 15 9 15
5 9 15 13 15 3
8 6 9 15 7 15 13 13 15
13 3 13 3 16 15 13 9 15 1 0 13 15 13
8 7 0 3 13 9 15 13 15
13 7 13 1 15 7 13 1 11 7 13 13 15 15
10 7 9 15 13 15 9 0 1 9 15
12 11 3 13 9 7 9 7 9 1 9 7 9
43 1 0 1 12 9 9 11 9 13 0 11 11 7 13 11 11 11 3 9 15 13 11 7 0 9 7 11 13 11 1 9 11 7 11 13 9 0 1 11 0 9 1 9
21 7 13 1 15 9 0 13 9 9 1 9 9 3 13 13 1 9 9 11 9 13
3 13 9 0
21 0 9 13 15 7 0 9 7 9 13 15 7 13 0 1 0 7 0 1 9 0
6 7 13 0 9 9 0
8 13 3 13 9 13 15 1 15
9 9 0 15 13 15 13 1 13 9
5 13 3 9 0 9
6 7 3 13 13 1 15
4 13 3 15 16
8 13 9 1 9 0 13 9 11
12 0 3 9 3 13 9 0 13 7 1 9 13
5 7 13 15 9 13
3 15 3 13
4 13 3 13 15
13 13 12 9 3 13 3 13 7 13 9 3 3 13
4 7 13 1 15
3 9 15 13
5 0 3 13 1 15
6 13 3 15 3 9 13
4 3 15 15 13
4 7 13 1 15
9 15 13 7 13 7 0 13 9 15
5 15 3 9 13 15
11 13 3 0 15 15 13 0 13 9 9 15
27 0 15 13 9 0 7 9 15 9 1 9 15 7 13 9 15 7 13 9 1 9 15 7 9 13 9 0
8 0 3 3 15 13 13 1 9
32 13 3 3 13 15 15 9 11 13 15 7 13 15 13 15 9 7 13 9 0 0 9 3 9 1 15 7 9 1 9 13 13
5 15 13 9 15 13
3 1 15 13
32 11 3 0 9 0 13 15 1 11 7 13 15 9 1 9 12 9 13 9 7 3 13 15 1 0 9 7 13 15 15 3 13
4 7 13 15 9
10 16 9 13 0 13 9 0 16 13 9
6 7 13 11 1 15 13
15 13 13 16 3 1 9 12 0 13 9 7 1 0 9 0
8 13 15 0 9 9 1 9 0
4 7 13 15 9
10 15 3 16 13 15 1 15 13 15 15
5 7 13 11 13 15
4 13 1 15 9
2 13 13
9 9 9 15 13 15 7 0 12 13
14 7 13 15 1 11 7 13 15 1 9 0 7 13 15
23 13 3 13 16 9 15 13 1 15 13 15 7 1 9 13 15 16 3 1 9 13 9 15
5 3 13 9 9 15
10 7 13 0 9 9 13 1 15 1 9
9 7 13 15 11 1 9 0 1 11
8 7 9 13 1 15 9 1 15
8 7 3 13 1 9 15 13 15
21 7 13 1 11 1 15 13 13 7 13 1 9 15 1 9 0 1 9 7 13 13
14 7 13 15 9 11 9 7 13 9 13 9 3 13 13
15 7 13 9 13 9 13 7 15 1 9 9 13 13 1 15
6 13 3 13 1 15 16
8 3 13 15 9 0 1 9 15
14 7 15 13 15 7 13 15 1 9 9 13 1 9 15
2 7 13
6 3 0 3 13 9 0
4 7 13 1 15
5 3 13 15 9 0
11 15 13 13 1 11 13 3 3 1 9 15
2 13 3
11 6 13 15 16 15 9 0 13 1 9 15
5 1 9 3 13 15
39 0 9 13 1 9 0 1 11 3 13 15 9 12 9 7 12 9 16 13 9 1 15 9 7 3 1 12 3 15 13 13 11 3 1 11 0 1 9 9
20 7 0 13 0 1 11 1 11 9 7 3 12 3 1 15 13 15 3 11 0
31 7 13 15 9 15 1 9 13 7 13 13 15 3 1 9 7 13 15 1 9 9 1 15 9 15 13 13 16 13 15 13
7 0 3 13 1 9 15 13
14 7 1 9 13 9 13 9 9 0 7 13 9 0 13
1 13
7 15 13 15 7 15 11 9
4 13 13 13 15
4 13 15 15 13
2 0 0
5 7 13 15 11 13
3 13 1 15
12 7 13 9 1 15 7 13 15 15 1 15 13
13 15 13 9 0 16 9 7 9 13 0 9 7 13
10 7 13 9 1 15 1 0 9 7 9
8 13 3 1 9 13 1 9 0
12 9 3 0 13 13 9 0 7 13 15 1 15
9 7 13 1 15 13 9 7 13 15
13 13 3 9 15 15 13 13 9 0 13 15 1 15
9 0 3 1 15 15 9 13 13 15
5 15 13 11 9 0
11 7 13 3 13 15 13 16 13 11 15 13
12 13 3 9 13 13 1 0 9 7 9 13 15
13 7 13 1 15 7 13 15 16 3 13 13 1 15
6 0 3 13 1 15 16
6 7 13 13 1 9 0
25 13 3 13 15 9 16 13 13 9 0 7 0 13 13 11 1 9 0 7 13 12 9 13 1 9
7 9 3 13 1 15 13 9
7 16 3 13 13 13 1 11
9 13 1 9 7 13 9 15 1 9
5 7 13 11 13 15
9 9 1 9 15 13 15 3 13 15
7 7 0 13 13 9 9 0
5 13 3 15 9 15
22 7 13 9 15 13 1 0 9 16 13 13 15 7 13 7 13 12 9 16 13 15 15
9 13 3 11 11 13 1 9 0 13
26 9 3 13 15 7 15 13 1 15 1 9 9 15 13 3 3 3 11 7 11 9 0 15 13 9 11
5 7 13 1 11 11
3 3 13 15
12 7 13 9 1 9 7 13 15 1 9 15 13
13 7 13 3 13 1 12 1 9 7 6 9 0 9
9 7 13 11 13 0 13 15 15 13
6 9 16 13 13 15 13
6 7 13 9 13 15 13
2 13 15
6 7 3 9 13 1 15
16 7 13 13 15 9 7 13 1 9 15 3 13 11 1 9 15
20 13 3 3 9 1 15 7 13 15 9 0 13 7 13 15 1 15 1 9 15
9 0 3 13 13 1 9 7 13 15
34 7 13 1 12 1 9 7 0 13 13 7 13 13 9 7 9 15 13 13 1 0 9 0 7 0 7 1 11 7 9 0 13 13 15
19 7 6 9 1 9 13 9 15 13 13 7 13 13 15 7 13 15 1 15
18 7 3 13 3 13 15 9 13 1 9 1 9 13 15 1 9 1 11
6 9 13 15 15 9 15
6 15 13 0 15 13 9
7 15 13 13 9 3 12 9
9 13 3 11 9 15 13 13 1 15
5 15 13 1 9 15
14 15 13 0 13 13 15 15 9 15 7 13 13 7 13
12 7 16 13 16 9 13 9 0 1 9 13 9
2 13 13
15 7 3 13 1 15 13 1 15 13 13 1 9 15 13 9
6 7 13 15 9 13 16
3 13 0 3
12 7 1 0 13 7 13 9 9 11 13 1 9
3 7 13 15
3 13 1 15
7 7 13 15 1 9 15 13
9 7 13 9 0 11 15 1 9 15
10 7 13 9 15 7 9 1 9 15 13
9 1 15 1 9 7 9 13 7 13
6 7 13 11 13 1 15
6 3 13 0 9 7 13
8 3 13 13 9 7 9 1 9
5 0 3 13 1 15
18 1 15 9 0 13 15 3 7 9 13 3 3 0 7 15 13 7 13
5 0 3 13 1 15
6 3 13 15 1 0 9
16 13 3 3 9 1 15 16 15 9 9 0 3 13 1 9 0
16 16 3 3 3 7 0 13 7 0 3 13 15 9 15 1 0
9 7 15 3 13 9 0 1 9 0
15 16 3 3 3 13 9 0 9 7 0 13 15 7 9 13
11 7 9 0 1 9 0 13 7 12 13 15
7 7 15 13 0 3 13 0
3 0 0 13
6 15 3 1 9 13 15
8 15 13 15 3 13 13 1 9
6 7 13 11 13 1 15
41 3 3 0 13 13 15 13 11 3 13 15 15 7 15 1 15 13 3 13 1 9 0 7 9 9 13 7 13 7 13 3 13 1 15 15 3 13 13 3 9 12
9 7 13 15 16 9 13 9 0 9
12 13 3 7 1 0 9 13 15 1 9 7 13
16 7 13 15 9 7 9 16 1 9 13 15 16 13 9 1 15
5 0 3 13 9 15
5 13 7 13 1 9
3 0 3 13
5 13 3 11 1 15
2 13 15
14 15 13 1 9 0 3 13 7 0 13 9 13 7 13
3 13 9 15
3 0 3 13
8 7 13 15 9 15 3 3 0
17 13 3 1 9 0 13 1 9 13 15 7 13 1 9 1 9 0
51 7 3 13 9 13 9 15 7 13 1 15 12 1 12 15 7 9 13 11 15 13 11 7 11 9 15 7 11 7 11 11 7 11 11 7 11 11 0 7 11 13 11 11 0 7 11 0 15 13 3 9
43 7 13 1 15 13 1 9 0 7 9 9 15 7 9 0 9 1 15 11 7 1 11 7 9 0 7 0 15 13 13 15 7 13 15 1 9 7 13 1 9 0 13 15
15 7 15 9 13 13 15 15 16 9 1 15 13 7 13 15
7 0 0 16 15 13 9 0
6 0 13 3 16 13 15
6 0 13 3 16 13 15
21 0 13 3 13 15 9 7 3 13 15 7 13 7 13 9 15 3 0 9 0 1
7 6 3 9 15 0 1 9
7 1 0 3 13 9 9 15
8 3 6 15 0 16 13 9 15
10 6 15 13 15 3 16 13 7 13 15
8 6 3 13 3 1 15 15 9
8 1 0 3 13 0 9 9 15
4 7 15 13 13
3 13 9 15
3 13 13 15
6 13 15 1 13 15 9
12 0 3 13 1 15 13 7 1 13 15 3 13
12 7 3 13 16 13 15 9 3 15 13 15 3
9 7 16 13 13 15 15 15 9 13
6 3 3 9 13 15 13
9 7 16 13 13 15 15 15 9 13
5 3 3 9 0 13
10 3 3 9 9 1 9 13 16 13 0
17 7 13 9 15 0 7 13 9 0 16 0 0 13 1 0 7 0
9 13 3 0 3 3 9 15 0 13
7 7 3 13 16 3 13 15
6 3 13 16 3 13 15
4 13 7 13 15
5 13 7 13 15 15
12 9 0 13 7 0 7 13 15 13 1 9 15
5 3 13 9 9 13
7 3 12 7 1 9 13 15
5 13 9 1 9 15
7 13 3 0 13 3 9 15
19 15 3 13 9 15 13 1 9 9 15 7 9 15 13 1 9 15 3 13
23 7 3 13 13 9 15 9 13 16 13 9 15 13 1 9 15 0 9 1 9 15 3 13
18 9 13 3 9 1 9 15 7 3 13 13 9 15 13 1 9 9 15
13 13 3 9 0 13 9 0 7 9 0 13 9 0
11 3 1 9 3 13 9 7 1 9 9 13
19 0 9 1 0 9 9 15 13 0 7 0 9 1 0 9 9 15 13 0
7 1 9 3 9 13 9 15
11 15 3 15 13 9 9 7 3 13 15 13
16 0 13 1 15 7 13 9 15 7 13 15 13 15 15 13 0
14 0 13 9 13 9 15 13 7 13 7 13 9 1 9
12 9 3 13 13 9 9 0 7 3 13 13 15
5 13 3 13 1 9
6 7 13 9 9 0 0
11 3 13 15 9 0 1 9 9 13 1 11
11 9 3 15 9 13 3 13 15 13 15 0
16 13 3 1 11 13 1 15 9 0 13 15 16 13 13 9 15
10 0 3 13 1 11 13 15 3 13 16
6 0 13 15 3 13 15
9 13 3 9 15 7 9 0 13 15
14 3 3 15 3 13 1 9 13 1 15 9 9 13 15
8 13 3 0 16 1 9 15 13
9 0 3 3 15 0 13 13 1 15
7 7 13 9 7 13 9 15
11 3 15 9 13 1 9 13 13 1 15 9
6 7 13 0 13 7 13
5 7 0 13 7 13
13 13 3 0 11 13 15 15 7 13 15 13 9 13
2 13 15
10 7 13 15 1 9 13 13 13 9 13
19 7 13 1 0 13 11 1 9 13 11 7 1 15 13 9 15 7 9 0
27 16 3 13 15 1 9 9 7 6 13 13 9 0 9 15 7 0 13 9 7 9 1 9 0 13 1 15
6 7 13 15 9 13 15
3 7 13 15
5 7 13 13 1 9
3 13 3 13
2 7 13
1 13
11 7 13 0 7 13 13 7 13 15 9 15
21 13 3 9 15 7 13 9 13 16 9 0 13 1 15 7 16 13 9 9 9 15
13 7 13 9 0 1 15 11 1 15 7 1 15 9
12 7 13 12 15 1 9 15 11 13 1 11 13
7 15 3 13 13 7 15 13
6 13 3 1 15 9 13
7 11 9 13 15 1 15 13
17 1 0 9 13 0 1 9 7 9 7 9 0 7 0 0 13 9
5 7 13 11 13 15
21 13 13 11 15 13 7 13 16 0 13 0 13 0 13 15 0 13 0 13 0 13
10 13 3 9 0 13 13 1 9 1 11
5 15 13 1 9 13
4 9 3 9 13
4 7 15 13 13
5 9 3 0 9 13
4 7 15 13 13
2 9 3
3 3 0 9
6 0 13 1 15 13 13
14 6 15 13 9 15 1 9 15 15 13 9 15 1 15
3 13 3 15
8 0 13 9 9 11 9 15 13
8 0 3 1 9 0 0 15 13
14 9 3 7 9 9 0 13 1 15 3 13 15 1 15
12 0 13 9 13 1 9 7 13 15 15 7 13
5 13 15 7 3 13
6 13 15 7 3 13 15
10 13 3 11 9 7 9 13 7 9 13
2 7 13
2 9 13
8 13 9 0 13 7 13 7 13
11 13 3 15 12 1 9 16 13 13 1 15
6 7 13 1 9 0 13
43 7 6 9 1 9 15 13 9 7 13 16 13 1 9 0 13 9 9 7 13 3 1 9 15 13 15 13 13 9 15 9 7 9 9 15 13 7 13 9 15 7 13 9
9 13 3 9 13 15 13 1 15 13
18 0 16 13 13 9 13 13 3 15 7 0 9 13 15 15 16 9 13
6 13 3 11 13 1 15
5 11 13 15 15 13
4 0 3 13 13
5 12 9 13 9 15
10 12 13 0 12 12 9 7 0 12 12
8 3 13 3 15 13 12 15 13
6 15 3 15 3 13 15
4 13 3 11 13
5 13 16 15 0 13
4 0 3 13 15
3 3 13 13
4 13 1 9 15
6 9 1 9 15 3 13
10 0 3 9 13 9 15 7 9 15 13
4 9 15 3 13
9 0 3 16 13 3 13 13 9 15
5 9 9 15 3 13
10 0 3 9 15 9 13 15 1 13 15
7 7 15 0 13 15 3 13
4 13 15 15 9
8 7 13 13 1 15 13 1 15
7 15 0 13 15 3 9 13
4 13 3 1 9
4 9 15 13 15
3 13 1 9
17 13 3 9 0 7 13 1 15 9 1 15 13 9 9 0 1 15
5 13 13 13 9 15
12 7 0 13 1 9 7 13 13 16 3 13 9
12 7 0 13 1 9 9 7 13 9 7 13 15
11 7 0 13 1 9 0 7 13 13 9 3
3 6 13 13
5 13 9 13 3 13
4 15 13 9 0
3 0 3 13
19 15 13 13 13 9 9 0 7 0 1 9 16 13 3 13 7 13 3 13
4 9 13 9 0
6 7 15 1 9 13 13
17 1 0 3 13 9 7 13 9 1 9 15 16 3 9 13 13 13
26 7 15 1 9 15 3 13 1 9 13 9 7 0 9 3 13 15 1 9 9 13 7 1 9 9 13
20 7 15 1 0 9 0 13 15 0 9 7 0 13 9 13 7 9 13 1 9
19 15 3 9 13 13 15 9 7 1 9 13 7 1 9 13 16 13 13 9
17 13 3 0 15 3 13 15 7 13 15 3 13 13 7 1 9 13
5 13 15 3 3 13
15 13 3 1 15 9 7 9 15 7 3 13 13 1 15 9
5 7 13 15 13 16
10 9 15 7 9 15 3 13 13 15 13
13 9 15 7 9 15 0 13 13 9 0 7 13 15
14 13 3 1 12 1 9 7 0 13 1 9 7 9 15
4 7 13 1 15
5 13 1 0 9 9
2 7 13
12 7 13 9 0 1 9 7 13 15 7 13 15
5 13 3 13 15 13
8 0 3 13 13 9 7 9 0
2 7 13
3 7 13 9
4 7 13 1 15
4 3 13 9 15
8 13 3 15 13 15 13 1 15
11 7 13 1 9 0 15 13 1 0 9 11
8 13 3 11 7 13 13 1 15
4 7 9 0 13
9 15 13 15 7 15 11 9 9 0
3 13 15 15
3 3 13 15
7 13 3 9 0 13 1 9
22 1 0 3 9 13 15 7 13 15 9 0 7 9 13 7 13 9 13 13 9 1 9
10 0 3 13 9 16 9 0 13 1 15
10 7 13 15 16 3 13 15 1 9 13
9 13 3 3 9 9 0 13 1 9
9 7 13 15 16 13 15 1 0 13
3 7 13 15
18 13 3 9 1 9 13 1 9 7 13 15 9 1 9 1 9 7 13
12 13 3 13 13 13 7 13 1 9 7 1 9
25 13 3 13 13 7 13 1 11 7 13 13 9 1 15 9 13 13 7 13 1 9 0 7 13 15
15 7 13 15 15 9 9 0 13 1 15 16 9 0 13 13
7 0 3 13 1 9 13 15
14 13 3 15 15 9 1 15 13 9 16 13 1 15 13
5 11 3 13 15 13
11 13 15 1 9 15 7 13 15 15 13 9
10 7 13 1 15 9 13 15 13 15 11
9 13 3 3 13 15 11 13 15 9
5 13 3 15 13 15
3 7 0 13
5 3 13 9 13 15
37 7 9 13 1 9 9 1 12 1 12 9 15 9 13 15 9 3 1 12 3 3 13 13 13 1 9 13 15 9 9 15 7 3 13 9 9 15
3 7 13 11
5 15 13 13 15 15
11 13 3 15 15 13 11 7 15 1 15 13
8 9 9 13 15 7 13 7 13
3 11 3 13
7 15 3 13 9 13 1 15
28 13 3 9 16 3 13 15 13 13 7 13 1 15 1 15 9 13 15 15 13 15 1 15 9 7 16 13 3
4 0 3 13 15
1 13
5 9 9 15 13 15
3 13 1 9
3 13 9 15
3 3 13 9
3 3 13 15
5 3 13 7 13 13
19 13 3 1 9 3 13 15 13 3 11 7 11 7 11 7 9 9 7 9
3 13 3 15
4 7 13 15 15
4 3 13 15 15
4 13 13 7 13
7 7 13 15 15 13 16 13
2 9 13
13 7 13 15 9 15 7 13 3 7 13 13 15 13
5 7 13 15 9 15
8 0 3 13 15 3 13 15 13
13 15 3 13 1 9 7 9 7 9 7 9 7 9
4 3 12 9 13
10 7 1 15 9 13 3 13 7 3 13
19 7 15 3 13 15 13 1 9 0 7 9 1 9 15 13 1 9 1 15
37 13 3 11 9 13 1 15 15 7 13 15 16 9 13 1 15 16 11 13 1 0 1 15 3 16 11 13 15 1 0 3 16 9 15 1 0 13
3 7 13 11
3 11 15 13
4 7 13 13 15
8 7 13 15 9 13 15 15 13
11 7 13 15 13 12 1 9 0 9 13 11
18 9 3 13 1 15 13 7 13 15 13 15 1 9 0 7 13 9 13
5 9 3 13 13 15
19 13 9 16 13 1 0 9 7 9 13 7 13 9 16 3 1 0 9 13
4 13 3 1 15
3 0 3 13
20 3 13 3 3 12 9 7 9 12 16 3 3 15 13 1 15 9 0 13 9
6 13 3 9 3 12 12
5 13 3 1 9 15
7 13 15 1 9 1 12 12
6 7 13 3 7 13 15
12 7 13 7 13 15 15 7 13 13 15 9 12
5 15 15 13 9 13
4 0 3 13 13
13 11 9 7 15 3 11 0 3 16 9 12 0 13
3 13 3 15
6 15 3 15 15 13 13
4 13 3 11 13
2 11 0
22 16 15 13 1 15 13 3 13 15 15 7 3 13 9 15 1 15 9 7 13 1 15
9 15 3 3 13 9 15 13 13 15
10 7 15 3 13 9 15 15 1 13 15
14 15 3 9 13 9 16 13 15 9 7 15 13 7 13
24 15 3 3 13 15 15 7 15 9 0 9 0 13 15 3 13 1 9 15 7 0 7 0 9
5 13 3 15 1 9
14 13 15 1 13 3 15 3 13 13 9 16 13 9 0
20 13 3 1 9 0 3 9 12 7 13 11 7 11 7 11 13 1 9 13 15
25 7 6 9 12 1 15 13 15 13 11 7 11 15 13 15 1 9 13 9 15 15 13 13 1 11
9 11 3 7 13 1 15 13 13 9
12 13 3 15 13 9 15 7 12 9 13 1 15
33 7 13 3 13 15 1 15 13 11 1 11 9 0 13 15 3 13 7 13 9 12 12 15 7 12 11 7 12 11 3 13 15 13
9 0 3 15 13 13 9 7 13 15
9 7 13 3 15 13 15 0 1 9
6 7 9 13 1 9 13
5 0 13 9 15 13
12 7 15 3 13 1 0 9 15 1 0 15 13
13 13 3 1 0 9 13 15 1 9 13 15 9 0
7 7 6 9 1 9 13 13
4 9 13 15 15
8 13 1 9 15 16 0 15 13
20 7 6 9 13 15 7 3 13 7 13 15 1 9 7 3 13 1 15 13 15
11 7 13 15 9 15 16 13 15 7 3 13
12 6 9 0 7 13 3 13 1 15 7 13 15
10 3 3 13 15 13 15 9 7 13 15
13 13 3 11 9 0 7 13 9 7 13 15 9 15
7 13 3 15 15 1 9 0
13 15 3 13 15 1 15 15 13 11 13 1 9 15
6 13 1 9 15 9 0
9 9 3 0 13 13 15 1 9 0
17 13 3 13 1 15 16 3 13 15 7 13 15 13 15 1 9 0
10 13 3 9 1 15 15 15 0 13 13
18 15 3 13 9 0 1 9 15 15 13 7 15 3 13 15 13 13 15
10 15 3 0 13 1 15 15 0 13 0
4 13 3 11 13
18 9 13 15 1 9 15 13 9 7 13 15 16 1 9 3 13 1 15
5 7 13 1 15 11
4 13 3 1 15
8 15 3 13 1 15 1 15 13
22 13 3 3 13 15 9 9 15 7 0 13 9 15 1 11 13 7 13 9 1 9 15
11 7 3 13 15 16 9 15 13 13 1 11
8 13 3 9 15 11 7 11 13
17 9 13 3 7 13 16 9 13 1 9 7 13 15 3 3 11 13
5 13 3 15 13 15
9 13 3 13 1 9 13 15 1 15
7 13 1 15 3 3 13 9
4 7 13 15 11
15 9 9 13 7 9 0 9 7 9 0 3 13 3 13 9
4 13 1 9 15
3 0 3 13
8 9 13 15 3 13 13 9 15
5 13 0 13 15 9
6 15 3 13 13 9 0
4 13 3 7 0
4 13 1 15 9
11 3 3 13 13 15 15 15 13 1 9 15
14 15 13 9 15 1 9 7 13 3 13 13 1 9 0
27 7 1 0 3 13 9 3 15 12 12 7 13 15 1 12 1 9 15 1 0 9 7 9 3 13 0 13
6 9 3 0 7 9 3
11 13 15 3 9 9 16 13 9 1 9 15
1 13
9 6 15 13 15 3 9 1 9 9
13 3 13 9 7 9 7 9 7 15 1 9 3 13
7 1 15 9 13 3 3 13
11 7 16 13 3 9 9 13 1 15 9 15
12 1 0 3 9 13 13 7 13 15 13 1 15
6 0 3 13 9 9 15
6 3 13 1 9 1 9
22 7 1 15 9 3 13 7 13 15 13 13 15 7 13 0 15 13 1 15 7 13 15
6 13 15 1 15 9 0
14 1 15 3 9 13 7 3 13 15 13 1 9 15 13
9 3 9 13 15 1 9 15 13 15
6 6 15 11 6 15 11
22 3 16 1 11 7 11 13 9 13 13 1 15 3 3 1 9 7 9 13 13 15 13
10 3 11 7 11 3 13 1 9 3 15
11 7 15 11 1 9 13 15 1 9 13 15
11 13 15 15 13 7 13 15 15 15 15 13
8 7 13 15 15 13 15 13 15
8 13 3 15 12 12 1 9 13
9 9 3 9 13 15 15 1 9 15
7 13 9 3 9 1 9 13
19 6 13 15 9 13 1 9 7 9 7 1 15 9 9 7 15 15 3 13
11 3 1 0 3 13 15 16 9 15 13 15
9 13 3 15 16 9 15 13 13 9
9 1 0 9 13 15 9 11 7 13
20 13 15 15 9 9 9 7 9 16 13 13 0 1 0 7 0 7 13 0 9
8 6 9 3 0 13 9 1 15
6 7 13 15 1 9 13
5 0 9 13 15 13
23 13 3 15 16 0 9 7 9 13 13 15 15 13 7 3 13 7 13 15 13 7 3 13
11 7 6 9 15 13 1 11 13 15 7 13
6 9 15 13 9 0 13
5 0 3 13 1 15
5 1 9 15 13 13
2 3 13
26 13 9 9 15 1 15 9 15 7 15 9 15 7 15 9 15 7 15 9 15 7 0 15 3 0 15
2 3 13
5 0 13 7 0 13
9 0 3 13 13 15 0 13 1 11
5 7 15 13 0 15
4 13 3 11 13
23 9 15 13 1 11 1 11 7 1 9 13 15 7 13 15 7 9 13 13 13 3 0 13
13 3 3 3 9 13 1 0 9 13 7 13 15 13
20 9 3 15 13 13 1 15 7 13 15 13 7 13 13 9 15 13 9 7 9
9 7 1 0 13 13 12 9 13 9
3 7 13 15
12 13 15 7 15 3 13 15 3 13 15 13 15
11 15 3 0 12 0 13 15 13 13 1 9
3 0 3 13
3 13 15 11
5 13 7 15 13 3
11 13 3 13 15 7 0 13 11 1 9 15
15 7 0 13 9 9 11 15 3 13 1 9 0 13 9 15
6 7 11 13 1 0 9
3 13 3 13
11 9 3 13 3 16 9 15 12 15 13 13
5 13 3 13 15 11
8 11 11 13 15 7 13 1 0
5 12 3 13 1 9
11 11 3 0 9 13 15 3 13 15 1 15
10 9 13 15 13 15 3 11 13 9 15
3 13 3 15
10 3 13 15 13 9 15 15 13 1 9
4 3 13 9 15
10 3 13 9 15 3 1 9 3 1 9
8 9 15 0 13 15 1 0 9
5 7 13 15 9 15
7 3 3 0 13 0 9 15
4 7 13 1 15
14 15 1 15 13 9 7 13 1 15 9 9 7 13 15
15 3 9 15 13 1 9 1 15 7 3 13 15 13 1 15
5 7 1 3 13 13
4 3 13 15 9
12 3 9 13 13 7 9 15 1 15 1 9 13
5 3 13 13 13 15
2 13 15
4 7 15 13 15
3 13 7 13
5 13 7 13 15 15
11 0 3 13 13 7 13 13 7 13 13 15
12 15 3 1 15 9 13 9 9 3 9 13 15
9 7 9 3 1 9 9 9 13 15
8 7 16 13 9 3 13 15 9
22 16 3 15 0 13 13 9 0 13 9 15 3 3 9 1 9 13 9 0 13 1 15
4 7 13 15 9
5 15 3 1 15 13
6 1 11 9 9 13 9
9 0 3 13 9 1 15 13 1 9
7 0 3 13 15 9 13 15
13 0 9 13 15 0 1 15 13 7 9 1 9 13
13 16 3 3 9 0 1 15 13 15 3 13 9 15
7 3 13 1 11 13 15 9
6 0 1 0 13 15 9
15 16 3 3 1 9 0 15 13 9 3 13 1 15 9 0
12 3 0 13 15 13 15 9 1 9 13 9 15
19 7 16 0 15 13 13 15 7 15 9 15 13 1 15 13 7 9 15 13
14 15 13 1 15 1 15 13 7 15 3 13 1 15 13
17 3 3 0 9 13 1 9 13 1 0 9 13 9 7 3 13 13
8 13 15 1 9 15 1 3 13
6 7 13 13 13 7 13
9 0 9 13 15 7 9 15 13 13
3 0 3 13
9 0 3 3 0 13 9 0 7 13
6 9 3 13 15 13 13
4 9 0 0 13
12 9 13 7 9 3 13 15 15 3 9 11 9
13 3 3 13 11 9 9 3 13 7 9 0 9 0
13 3 13 1 9 9 13 9 0 7 6 3 11 3
14 7 13 15 16 13 15 1 9 0 7 6 3 11 3
17 15 3 9 13 1 9 13 7 1 9 7 1 9 16 13 13 9
4 9 9 13 9
12 3 3 9 15 0 13 3 15 9 15 0 13
9 7 16 0 13 3 9 15 0 13
10 13 3 16 9 15 13 1 15 9 13
11 3 3 13 13 15 9 15 16 13 1 15
3 13 3 13
4 13 9 1 15
16 3 15 9 0 9 7 9 13 7 0 15 0 13 9 7 9
10 0 3 15 3 13 13 0 3 0 13
10 3 13 13 9 7 6 15 0 15 13
20 7 6 15 9 16 9 13 1 9 7 9 7 0 9 7 13 9 7 9 0
12 6 15 9 16 13 9 1 9 7 9 1 9
19 6 15 9 7 9 7 9 3 13 3 9 3 13 7 9 13 1 3 13
7 13 3 15 1 9 13 15
7 0 3 13 3 15 9 6
17 16 13 1 9 9 3 13 7 0 3 12 3 9 15 13 15 9
11 6 15 16 13 9 9 9 3 15 13 15
18 3 13 7 9 13 9 9 15 16 0 3 13 15 15 3 13 15 9
38 13 1 15 9 7 9 7 1 15 13 7 13 16 13 15 9 15 9 13 1 9 15 9 1 9 0 1 9 11 0 1 9 11 13 1 9 7 9
3 6 13 15
5 13 15 1 9 0
7 6 15 9 16 13 9 9
30 13 3 15 1 15 3 13 9 7 9 3 3 13 15 7 13 15 1 0 13 15 13 15 1 9 15 16 1 15 13
16 1 15 13 15 9 9 16 13 15 15 13 13 1 9 15 3
8 13 15 1 9 0 15 13 9
20 3 15 1 9 13 1 9 13 15 7 15 1 9 13 1 9 13 15 1 9
5 13 3 15 9 15
14 3 13 15 1 13 9 7 1 0 3 13 0 15 13
6 13 3 15 15 15 13
9 13 15 13 9 1 9 13 1 9
3 0 13 15
8 3 12 3 9 13 15 9 12
8 7 3 9 9 15 15 13 13
3 3 13 15
5 3 0 9 0 13
3 13 3 15
15 0 15 3 13 15 1 9 3 9 0 13 15 1 9 0
11 7 13 15 15 1 9 13 13 1 9 0
10 7 15 13 1 9 0 3 13 15 15
11 0 3 9 13 15 1 0 9 15 13 13
6 13 3 15 15 1 9
9 9 13 9 15 16 13 1 15 9
4 0 3 13 15
9 9 15 15 13 9 7 9 1 15
4 13 3 1 15
18 13 15 7 13 15 1 0 9 16 1 9 15 9 15 13 1 9 15
5 7 13 1 15 13
9 15 13 16 3 13 3 13 9 15
2 7 13
2 0 13
6 13 9 15 7 0 13
13 7 13 3 15 9 15 7 0 15 7 13 9 15
8 9 13 0 0 13 1 9 0
1 13
1 13
2 13 15
4 13 3 15 9
9 0 1 0 9 9 15 13 1 15
5 7 15 13 15 13
8 3 13 15 7 3 1 9 13
3 0 13 13
5 13 9 13 3 13
13 3 13 15 9 15 15 13 7 9 1 15 13 15
8 9 3 0 13 9 7 9 9
16 13 9 16 3 13 7 13 15 13 9 7 9 7 9 13 15
6 3 3 15 13 0 9
12 15 3 1 15 13 15 13 13 9 15 9 12
11 16 3 3 0 15 13 15 1 0 13 15
4 13 9 3 13
16 13 3 15 16 3 11 1 15 9 15 13 15 3 12 1 0
14 7 15 3 13 15 13 13 7 15 13 7 3 13 15
7 15 3 0 9 9 0 13
7 15 3 9 13 16 13 0
10 3 13 9 0 7 0 15 13 15 15
12 3 13 15 0 9 16 13 9 15 13 15 9
6 13 9 15 7 13 9
10 3 3 13 9 15 3 3 9 15 13
7 13 9 15 13 7 9 13
8 0 9 0 15 9 13 13 13
4 6 13 15 16
9 13 15 7 13 15 7 13 13 15
15 7 1 0 7 1 0 9 13 7 13 3 0 13 9 0
24 0 3 13 16 16 13 13 9 9 1 15 9 9 13 13 3 13 7 3 13 13 13 9 15
4 13 3 15 11
10 9 1 15 3 9 0 13 7 1 15
3 13 3 9
10 0 9 0 15 13 9 15 13 13 3
11 1 9 13 15 16 1 15 9 15 13 15
51 16 3 3 13 9 0 1 9 15 13 9 15 13 7 13 13 9 7 9 13 3 7 13 7 13 15 13 9 9 0 1 15 9 3 13 7 1 9 1 15 3 13 7 13 15 7 9 15 1 0 13
19 0 3 9 13 9 9 15 7 3 13 7 3 13 1 9 15 13 13 3
18 0 3 15 13 13 0 13 15 1 15 7 15 13 0 0 13 1 15
5 9 13 13 1 9
7 15 13 16 3 3 13 15
12 9 3 13 13 15 7 3 13 15 16 13 15
3 6 13 15
2 7 9
41 13 3 3 12 1 12 9 13 12 1 12 7 12 1 12 7 13 15 9 1 9 7 9 1 9 9 1 9 7 9 1 9 9 1 9 15 7 9 1 9 15
14 3 13 9 13 1 9 3 13 16 9 13 7 13 3
10 7 3 9 13 13 16 9 13 7 13
12 9 9 9 7 9 13 13 7 9 0 3 13
8 15 3 7 1 15 3 13 9
32 3 3 13 1 9 15 1 9 1 9 13 9 13 1 15 16 3 13 15 1 9 7 9 15 13 9 7 9 15 13 1 9
9 3 13 13 3 16 3 0 9 13
18 13 3 15 15 1 0 9 13 15 1 9 15 9 11 13 1 9 15
13 13 3 16 9 0 0 3 15 9 13 16 3 13
3 6 13 15
8 7 16 3 13 15 15 3 13
25 7 0 12 1 12 1 15 13 9 0 7 13 15 13 3 16 0 0 13 3 15 9 13 1 11
3 6 13 15
8 7 16 3 13 15 15 3 13
7 9 13 15 1 9 15 13
4 13 3 1 9
12 6 0 9 13 13 9 1 9 0 7 3 13
2 13 15
4 3 7 9 13
5 0 3 13 13 15
13 9 13 15 3 0 9 16 15 13 3 7 13 9
5 7 16 3 13 9
21 7 6 9 13 9 13 0 12 12 1 12 9 7 13 0 7 3 13 15 13 3
8 13 3 15 11 13 7 13 15
6 9 13 13 1 9 15
5 7 13 1 15 9
7 7 3 13 15 7 13 9
12 13 3 9 13 16 1 9 13 15 11 13 9
7 12 9 13 1 15 13 13
11 1 0 3 13 13 15 7 3 1 9 0
17 9 15 15 1 9 3 13 3 15 9 7 9 1 9 7 13 13
23 0 3 9 0 13 15 13 9 6 0 1 12 9 3 13 3 13 15 1 9 1 9 0
21 7 6 15 13 13 15 15 13 15 15 7 15 9 13 15 1 15 0 13 1 15
2 13 3
5 15 0 13 9 0
4 7 15 13 15
13 0 13 9 0 9 0 15 13 9 13 1 9 15
15 7 13 7 13 1 9 0 7 9 0 13 15 1 9 15
14 0 13 9 15 13 9 13 1 9 12 9 16 13 15
12 7 13 1 9 7 9 13 7 9 13 1 11
5 13 3 15 1 15
6 9 3 3 13 13 15
5 0 3 13 1 15
6 13 15 13 1 0 9
8 3 0 13 13 13 7 3 13
4 9 9 13 15
5 3 13 15 3 13
3 3 13 13
11 13 1 15 7 13 7 1 9 15 13 13
2 7 13
2 13 15
5 3 13 15 3 13
23 3 13 9 7 9 9 3 13 11 7 11 7 11 7 15 9 1 9 0 15 3 13 3
15 7 13 1 9 7 9 7 9 7 9 7 13 1 9 0
8 1 0 9 13 15 9 13 15
9 13 7 13 3 16 11 13 15 13
3 7 13 15
4 13 13 9 0
11 6 13 9 7 9 13 3 7 1 0 13
25 11 11 13 9 7 9 13 13 1 15 3 9 13 13 9 15 3 9 9 15 1 9 7 3 13
6 6 13 15 15 9 15
12 13 3 15 16 3 13 13 15 16 13 3 13
19 7 13 3 13 11 1 9 15 9 0 1 9 9 13 7 0 13 13 15
10 7 6 9 15 13 0 9 13 1 15
10 7 13 13 11 13 1 9 7 9 13
5 3 13 1 9 13
8 7 13 15 13 15 7 13 15
5 7 13 1 15 13
16 15 15 9 7 9 1 9 13 7 3 3 13 15 1 9 0
7 7 3 13 13 15 1 0
25 3 13 13 15 1 9 3 13 1 0 9 16 15 0 15 13 13 7 13 13 15 7 0 13 15
3 13 0 9
8 7 3 13 1 9 0 9 13
3 9 13 3
8 3 13 15 9 1 13 1 15
11 3 0 13 15 13 15 7 13 15 13 15
5 13 3 1 13 15
29 3 13 9 7 9 3 13 15 15 7 9 15 7 9 15 7 9 0 16 3 3 0 15 3 13 7 13 15 9
7 13 3 15 15 1 9 0
10 13 3 12 1 13 1 15 0 13 15
4 0 3 13 15
17 9 15 13 9 0 7 13 0 7 13 9 15 1 9 9 13 13
6 13 16 3 0 13 15
6 7 13 3 13 15 15
3 0 13 15
9 9 13 7 13 9 13 7 13 15
3 13 15 0
4 9 0 13 12
4 7 13 13 15
2 13 15
3 13 15 0
3 7 0 13
8 9 13 7 0 1 3 13 13
8 7 13 9 0 13 0 9 15
3 7 13 9
8 9 13 3 13 7 3 9 13
4 7 13 9 9
13 13 1 9 7 9 7 13 13 16 13 15 9 15
14 13 3 15 16 3 12 3 9 0 13 3 13 15 9
7 0 3 13 13 3 3 13
12 13 3 1 15 9 0 7 13 15 13 1 15
30 16 15 13 1 15 7 3 13 9 15 7 9 7 9 7 9 7 9 7 9 3 3 3 9 15 3 13 15 9 13
36 15 3 1 15 13 9 13 3 3 3 13 13 9 16 13 15 13 1 9 16 3 3 13 9 7 3 13 13 15 13 13 13 15 15 13 16
8 0 9 13 13 7 3 13 13
30 7 15 9 13 1 15 9 13 15 1 9 3 13 3 3 13 16 0 13 1 12 12 13 13 1 12 12 12 1 15
14 16 3 3 3 3 3 15 13 9 13 13 15 1 9
17 3 3 0 1 15 15 3 13 15 15 15 9 3 13 15 13 9
3 0 13 9
8 16 3 9 13 1 15 13 15
8 7 1 9 7 1 9 9 13
12 13 3 1 15 13 15 15 9 7 9 13 15
14 7 13 9 7 9 13 16 0 9 13 7 1 15 13
7 13 3 1 15 9 0 13
29 15 9 1 15 13 12 9 7 13 12 1 15 3 13 3 12 12 7 12 1 9 7 13 1 9 13 16 13 15
18 7 13 13 1 9 15 13 15 7 13 1 9 13 9 7 9 13 15
9 13 15 1 15 16 13 9 15 13
24 13 15 16 3 9 13 1 9 1 12 9 13 15 3 1 12 12 7 12 9 15 3 13 9
7 7 13 13 9 7 9 13
13 3 13 15 9 13 1 9 0 1 12 9 13 15
3 13 3 9
5 9 15 13 12 9
5 7 13 0 15 9
6 9 13 15 0 9 9
4 7 13 15 9
15 13 3 15 15 13 9 0 1 9 0 7 0 13 13 15
17 7 13 13 15 15 1 9 0 9 7 13 15 1 9 15 13 9
5 1 15 3 13 13
6 3 9 9 15 13 9
4 15 3 9 13
5 13 13 1 9 15
3 7 13 15
7 3 13 0 13 15 9 15
7 13 15 3 12 1 9 15
6 7 13 13 1 9 15
4 13 3 15 9
7 9 13 1 9 7 1 15
7 3 13 0 13 15 9 15
6 13 3 9 1 9 15
23 7 13 9 0 13 7 13 3 13 15 16 9 15 0 0 13 7 13 13 13 7 13 15
4 7 13 13 15
7 13 3 9 15 0 1 9
11 7 16 13 13 15 1 9 13 9 7 9
4 15 3 0 13
5 0 3 13 15 16
13 9 15 13 7 13 9 15 9 0 16 0 15 13
6 9 3 15 13 13 15
6 0 3 13 13 9 15
25 6 3 9 13 15 7 3 9 15 3 13 7 15 3 3 13 13 9 16 1 9 15 13 15 13
15 3 3 9 15 0 13 15 9 1 9 13 13 15 9 0
4 0 3 13 15
19 13 3 15 7 13 13 16 9 15 0 0 13 7 13 13 13 7 13 15
6 13 3 7 1 9 15
5 7 13 15 13 15
5 15 0 13 1 15
5 13 9 1 9 0
7 3 13 3 1 0 9 13
6 13 3 1 15 9 9
10 15 13 16 9 15 13 9 9 1 15
3 13 13 15
9 7 13 12 15 9 9 15 13 0
5 15 0 13 9 15
3 0 3 13
4 12 9 1 9
3 7 13 15
3 13 9 15
6 7 13 3 13 12 12
3 0 3 13
3 12 9 9
3 7 13 15
7 13 9 15 7 13 12 12
9 7 13 9 9 0 16 3 3 13
12 3 9 9 0 0 3 9 9 1 9 15 13
4 3 15 15 13
14 13 15 9 1 0 9 16 3 13 13 15 1 0 9
14 16 3 1 0 9 3 13 0 1 0 15 15 9 13
11 7 16 1 0 0 3 13 15 15 15 13
7 15 9 3 13 12 9 13
16 7 3 12 13 7 0 13 7 12 13 15 7 1 0 13 13
6 3 13 9 13 7 9
11 13 3 0 15 3 9 9 13 7 13 15
3 7 13 15
6 15 13 13 15 1 9
5 9 7 9 1 11
5 3 9 0 13 15
13 0 3 13 9 7 9 13 3 1 9 12 9 13
17 0 13 9 15 7 13 15 9 13 7 13 15 13 1 9 9 13
18 9 3 15 13 0 7 13 15 1 9 7 9 13 15 1 0 9 3
22 0 3 13 15 9 11 15 13 1 9 15 0 7 13 13 15 1 9 13 1 9 0
7 7 3 9 13 13 9 15
7 13 3 3 0 7 13 15
4 7 0 13 13
4 9 11 13 15
19 7 13 11 16 13 9 9 15 1 9 7 13 9 15 16 13 1 9 0
3 13 3 11
15 9 13 16 13 13 15 0 15 1 9 15 7 11 3 0
8 3 3 3 13 15 7 15 13
2 13 3
28 13 15 3 9 16 15 13 1 9 9 15 13 3 12 9 16 3 13 15 16 3 3 0 13 1 9 0 0
4 13 11 7 9
3 3 13 15
6 0 3 13 6 9 11
10 7 16 15 1 0 13 1 15 13 15
3 13 3 15
4 13 3 1 9
6 0 13 16 3 13 9
5 6 3 0 15 13
2 13 15
14 16 3 13 15 9 15 13 15 7 16 13 15 13 15
17 7 16 3 9 13 1 15 7 3 9 13 15 13 13 15 13 15
4 7 13 9 9
3 13 3 9
12 16 13 13 9 3 9 0 13 13 3 9 0
7 13 15 7 13 15 1 9
4 7 13 13 15
3 3 13 13
5 7 3 13 3 15
19 13 15 13 7 13 15 13 15 16 13 7 13 7 1 0 13 7 13 15
2 3 13
10 3 3 15 3 13 15 13 15 13 16
9 9 0 13 16 15 0 13 13 13
12 7 13 13 15 1 11 7 0 13 1 11 11
19 7 13 15 1 15 9 13 15 12 0 9 15 13 3 7 0 13 9 13
5 7 13 15 13 15
4 13 13 15 9
23 12 3 1 15 13 16 13 13 15 1 9 0 13 9 7 13 0 1 9 15 9 15 13
4 7 0 13 9
4 13 3 11 13
5 3 12 3 13 15
14 7 12 3 3 13 15 13 15 13 9 9 3 9 10
3 7 13 15
4 9 15 13 15
6 3 13 9 0 1 9
6 7 13 6 3 7 3
8 6 3 9 0 3 1 15 13
4 13 3 1 9
9 13 9 3 13 12 9 9 0 13
3 7 3 13
3 7 13 15
4 3 13 7 13
18 3 3 9 13 15 1 0 1 0 13 15 3 13 9 0 1 9 15
12 3 3 13 15 3 13 7 13 13 1 9 0
13 7 3 13 1 9 0 3 13 3 1 9 9 0
18 13 13 13 15 13 1 15 9 13 11 1 9 7 13 9 7 13 15
7 3 7 3 13 1 9 0
3 13 7 13
3 13 7 13
1 13
16 1 15 9 13 11 1 9 13 9 7 9 1 9 7 13 15
11 1 0 13 3 9 1 15 9 0 13 15
27 1 0 9 15 13 1 9 7 9 15 1 9 3 3 13 13 15 7 15 1 9 3 3 3 13 15 3
3 13 9 0
16 7 15 3 13 9 15 15 13 13 15 7 15 13 15 13 15
2 13 15
8 1 0 9 13 12 1 9 12
5 12 13 7 0 13
4 12 13 1 9
5 12 13 7 0 13
4 7 13 13 15
2 3 9
4 0 3 13 15
6 3 9 3 9 13 15
15 9 13 15 1 15 9 9 3 13 15 7 9 3 13 15
5 13 15 1 9 15
6 7 3 13 1 0 9
5 3 3 13 1 15
27 16 7 9 3 13 15 7 9 3 13 15 16 13 15 9 9 0 3 13 15 16 3 1 9 13 13 15
3 13 3 9
5 13 15 9 0 13
8 13 15 16 13 9 15 1 0
10 3 9 0 13 3 13 3 9 1 9
7 9 12 13 1 9 13 15
5 12 9 7 0 9
6 9 13 1 15 13 15
17 9 9 15 13 16 13 3 3 0 9 9 9 9 7 3 0 9
6 13 15 12 9 1 9
11 7 9 3 13 3 13 3 9 13 1 9
5 7 13 9 15 13
5 9 0 13 15 9
8 13 0 13 1 9 15 3 0
11 3 0 13 15 13 15 7 13 15 13 15
11 13 3 1 15 3 9 16 13 15 15 13
5 13 3 9 13 15
10 3 13 9 13 1 15 7 3 13 15
5 0 3 13 9 0
3 6 13 15
13 15 3 3 13 9 0 3 9 3 13 13 1 15
7 9 0 15 13 9 0 13
4 13 3 15 11
4 15 15 13 0
2 9 13
2 3 13
3 3 9 13
2 3 13
4 3 0 9 13
3 0 3 13
6 15 0 13 1 9 15
4 3 12 13 13
17 15 15 13 13 7 13 0 7 13 13 9 1 9 7 13 1 15
6 0 3 13 0 0 13
4 13 3 0 3
6 13 3 11 0 13 13
8 3 3 13 9 1 9 0 13
3 13 3 13
3 0 3 13
7 0 1 9 0 1 9 13
3 13 3 11
4 6 15 13 15
4 7 1 15 13
4 0 3 13 15
33 6 13 15 16 15 13 15 13 9 7 9 7 9 7 9 7 9 9 0 1 15 3 13 3 1 9 0 7 1 9 13 9 0
22 13 3 15 9 7 13 15 15 7 13 15 7 13 15 7 13 13 15 7 0 9 13
18 7 0 15 1 0 3 13 7 13 9 0 13 1 15 7 3 13 13
14 13 3 3 13 15 11 1 11 9 15 13 1 9 13
5 13 3 9 13 13
4 15 3 13 0
7 13 3 15 16 11 9 13
3 7 13 13
5 11 9 0 13 15
6 0 3 3 3 13 13
4 9 0 13 15
8 13 3 11 13 13 15 1 15
9 13 3 15 15 1 15 13 15 13
5 15 13 16 15 13
3 0 3 13
3 9 16 13
4 11 3 13 15
10 7 3 13 7 1 9 15 13 13 9
7 7 15 9 13 13 9 9
6 7 13 13 11 1 11
15 7 6 9 9 13 11 7 0 13 0 9 7 0 13 0
14 7 13 13 11 15 13 7 3 13 9 16 9 0 13
13 7 3 13 13 1 9 16 13 15 16 3 13 13
9 7 16 13 1 9 13 11 13 15
4 11 13 15 13
9 7 13 15 13 7 13 15 13 15
11 7 13 15 13 13 16 1 0 9 13 13
6 13 3 11 13 1 9
15 6 9 9 15 9 13 0 7 16 13 15 15 13 13 9
6 13 3 1 15 11 16
11 3 9 9 15 13 16 3 0 9 0 13
21 13 3 15 0 13 9 13 16 0 13 1 11 7 13 16 3 13 9 0 13 15
2 13 3
15 13 3 7 12 9 15 7 13 15 12 9 7 13 1 15
4 9 13 16 13
5 9 3 15 13 15
6 13 9 1 9 15 13
7 3 13 0 16 13 1 15
4 13 3 0 13
6 9 9 15 13 12 9
7 7 13 15 0 9 7 0
4 7 13 0 13
6 9 15 9 13 12 9
4 13 3 3 0
6 7 15 13 1 12 9
9 9 6 9 15 15 13 13 1 9
8 13 3 15 15 16 9 0 13
9 13 15 3 13 7 13 15 3 13
2 13 15
15 13 16 15 9 0 13 13 15 3 13 7 13 15 3 13
8 7 1 15 3 13 15 9 9
8 7 15 13 1 9 13 15 13
4 13 1 15 9
5 7 13 13 12 9
3 7 13 15
4 9 13 12 9
17 13 3 15 16 0 13 13 7 1 3 13 3 15 13 13 1 15
8 7 0 13 13 3 13 1 11
18 7 13 16 13 15 1 11 7 11 1 9 13 11 13 12 9 15 13
3 13 15 13
8 7 16 15 15 13 3 13 15
4 16 9 13 15
7 13 3 13 13 3 13 15
9 13 3 15 9 13 9 15 1 15
3 15 13 9
13 7 13 15 1 11 7 13 9 15 1 9 13 11
25 13 3 15 15 3 1 9 9 0 13 15 9 9 13 15 13 9 9 0 1 15 9 15 13 13
5 0 13 1 9 0
7 9 1 9 7 9 1 0
8 7 15 9 1 9 13 1 15
4 9 13 9 15
4 7 13 13 15
10 13 15 16 16 3 0 13 9 13 13
7 3 3 13 15 1 9 15
41 3 13 9 1 15 7 13 9 15 9 1 15 7 13 15 7 13 15 3 7 13 15 7 9 15 1 15 7 3 13 1 15 9 1 9 16 3 13 9 9 15
13 7 13 1 9 13 13 13 1 15 7 13 13 15
2 13 13
5 9 15 9 9 13
6 15 3 13 15 9 9
8 7 13 13 1 9 1 15 9
10 9 3 7 9 13 15 13 7 9 9
7 9 3 15 13 15 15 13
26 7 13 1 15 1 9 0 13 15 9 1 9 7 13 13 15 9 7 9 1 9 7 13 13 1 15
13 13 15 15 9 0 13 7 15 13 13 15 9 0
5 13 3 13 1 15
9 13 15 3 15 12 9 7 13 15
9 9 0 1 9 3 13 7 1 9
7 0 3 13 1 15 13 16
5 16 13 1 9 13
8 0 3 13 9 16 11 9 13
2 7 13
3 3 13 3
4 11 3 13 15
8 3 15 13 15 15 9 0 13
7 13 3 1 9 13 9 0
12 9 13 9 7 13 15 9 7 13 1 9 0
5 9 3 13 13 0
10 0 3 3 0 13 7 13 15 13 0
4 7 13 0 13
6 0 3 3 0 13 13
4 13 3 9 9
2 15 13
4 13 9 15 13
9 13 3 15 9 13 15 1 15 13
3 0 13 9
6 13 15 16 15 13 9
7 7 13 15 3 1 9 13
6 15 3 13 15 9 9
9 13 7 13 9 0 7 13 9 15
3 13 3 13
6 0 3 13 1 15 13
5 15 3 13 13 0
10 9 15 9 13 13 0 13 1 9 9
6 7 1 15 13 13 15
16 7 13 9 7 9 13 1 15 9 1 0 9 7 13 15 9
8 13 3 16 1 15 13 9 0
21 7 13 13 9 13 15 9 13 16 13 15 1 9 16 13 15 13 9 7 9 9
18 9 13 16 3 13 7 13 7 3 1 9 13 7 1 9 9 0 13
8 13 3 15 9 9 13 7 3
7 13 3 9 15 13 1 15
3 15 15 13
5 15 13 9 7 9
2 13 13
1 0
11 13 3 15 13 0 9 7 15 13 0 9
15 7 3 13 13 9 15 1 9 7 13 15 1 9 15 13
12 13 3 15 1 9 13 9 3 13 13 15 13
26 9 11 13 13 15 16 15 9 13 13 9 7 0 1 9 13 16 13 9 15 9 7 13 9 9 15
4 12 3 9 13
21 7 13 0 9 7 0 13 0 7 0 13 15 3 3 3 15 12 13 3 13 9
6 1 3 15 3 9 13
5 12 3 13 15 9
5 7 13 11 13 15
7 9 9 0 13 15 7 13
16 7 13 15 9 0 13 7 9 15 1 0 7 13 15 7 13
6 7 13 3 1 0 13
11 0 3 13 9 7 9 13 0 9 9 13
6 9 3 13 0 7 0
5 13 3 15 9 13
3 9 3 13
8 1 0 3 3 13 15 13 15
4 13 3 1 15
7 3 13 15 11 13 9 0
7 7 0 11 13 1 9 0
4 13 9 9 15
8 13 3 15 9 13 1 9 15
32 13 1 9 13 1 9 13 7 13 9 1 9 7 9 1 9 7 9 1 9 7 1 9 15 13 9 9 7 9 3 13 15
4 0 13 9 0
9 13 3 13 13 1 9 9 15 0
12 13 3 3 15 9 0 13 3 12 9 7 13
11 1 9 13 15 16 9 0 0 3 15 13
3 0 13 13
5 13 9 13 3 13
13 7 15 13 1 9 16 9 0 7 9 13 13 13
16 0 15 13 13 9 1 15 3 13 9 1 9 15 3 13 15
4 13 3 15 13
5 9 3 3 0 13
8 7 15 13 9 3 13 0 13
3 0 3 13
6 13 15 16 3 13 13
8 0 3 13 1 9 15 13 16
9 3 3 13 9 7 9 3 13 15
10 13 3 0 3 13 7 3 3 3 9
3 3 13 15
8 13 9 1 9 7 9 1 9
10 9 3 0 1 9 7 9 7 9 13
8 9 3 7 9 1 9 0 13
24 1 3 0 15 13 1 15 9 15 7 13 13 1 9 7 9 13 1 9 7 9 9 15 1
10 13 3 1 9 15 3 3 13 15 13
22 13 3 13 9 7 9 7 9 7 9 7 13 1 15 7 13 13 1 15 9 15 1
6 7 9 9 15 3 13
6 1 9 15 13 9 15
13 3 3 13 13 9 11 3 13 16 13 15 9 15
34 3 13 1 11 3 13 1 9 7 15 1 9 15 3 13 7 15 1 9 3 3 13 1 15 16 9 9 0 13 16 13 15 15 13
8 6 3 0 7 13 1 0 9
20 7 13 9 1 9 7 9 7 9 7 1 9 9 9 1 9 9 0 7 9
14 13 9 1 9 7 9 13 1 9 9 3 0 13 15
15 13 3 0 13 13 15 7 13 9 15 16 13 15 9 15
4 7 13 15 9
5 13 9 7 15 9
13 3 13 15 3 13 1 15 13 16 3 1 9 13
13 3 3 15 3 13 0 13 13 16 1 13 9 0
9 9 7 9 13 7 9 15 3 13
21 13 3 15 16 3 13 9 15 9 7 9 7 9 0 7 13 1 15 3 9 0
11 3 9 3 13 1 15 13 1 9 15 9
16 13 3 1 9 13 1 9 7 9 13 15 13 1 9 13 11
12 7 15 9 1 9 13 1 15 1 9 13 15
16 13 3 15 9 9 13 9 7 13 9 7 9 3 15 13 13
4 13 3 15 9
10 7 13 13 9 7 9 3 15 13 15
10 7 13 15 7 13 15 13 9 7 13
10 7 13 0 9 16 15 13 15 1 9
16 13 3 9 9 1 15 0 13 13 9 7 13 11 7 11 13
4 0 3 13 15
4 3 13 16 13
4 0 3 13 15
8 1 15 13 1 9 1 15 13
4 7 13 9 9
3 13 15 9
9 3 13 9 3 9 1 9 15 13
7 7 0 15 13 9 0 13
9 13 3 13 3 13 15 7 13 9
12 7 3 13 9 13 7 12 1 12 9 1 15
12 9 0 13 9 13 1 15 3 16 3 13 9
16 13 3 15 16 3 3 13 13 1 15 16 13 15 1 9 0
6 7 13 9 9 13 13
5 13 0 7 13 15
3 13 3 15
11 3 3 13 13 1 9 0 16 9 0 13
7 0 13 9 15 13 1 15
6 7 9 3 1 9 13
11 0 9 0 9 15 9 15 1 15 13 15
10 3 6 9 13 15 1 15 13 1 9
14 7 9 3 0 1 13 13 3 6 9 0 15 13 13
14 7 0 13 13 1 15 15 3 13 1 15 13 13 0
12 13 3 3 9 1 15 15 13 15 15 13 0
4 0 3 13 15
7 15 3 0 13 3 7 13
3 3 13 3
8 15 3 1 9 15 13 3 13
9 15 3 13 13 1 15 1 9 15
30 7 15 13 15 3 13 15 9 15 9 16 13 7 13 1 9 15 1 9 15 7 13 1 9 13 12 1 12 9 0
3 13 3 9
11 11 11 6 9 13 15 16 13 13 3 9
11 15 3 13 15 1 15 16 3 13 9 15
4 0 3 13 15
12 9 1 15 0 13 7 1 9 7 1 9 13
3 0 3 13
3 13 15 11
12 3 13 9 3 16 12 9 13 15 15 3 13
3 7 13 15
15 3 13 15 1 9 7 1 9 7 1 9 3 15 13 13
3 0 3 13
10 7 3 15 13 9 3 13 3 7 9
11 7 15 3 13 3 13 9 15 7 13 9
14 13 3 15 16 3 13 0 13 16 13 15 1 15 0
5 7 1 9 13 15
6 3 15 1 15 9 13
3 0 3 13
5 9 6 9 3 12
2 3 13
5 1 15 13 9 15
6 13 3 1 9 13 15
7 13 15 16 3 13 1 9
8 7 15 13 1 15 3 9 9
6 7 13 9 13 15 13
8 9 16 13 13 9 0 1 15
9 13 3 15 15 9 1 9 13 15
7 7 13 1 9 3 13 15
12 7 13 1 9 13 1 9 13 15 13 1 9
3 7 13 15
2 15 13
8 13 13 15 16 3 13 1 9
23 3 3 15 13 6 9 7 13 11 12 1 12 1 12 1 15 13 7 13 1 11 13 15
4 15 13 0 13
4 11 3 13 15
6 11 9 3 9 0 13
4 9 3 13 9
13 7 13 12 15 1 15 0 9 7 13 15 9 0
4 13 3 11 13
3 13 1 0
13 13 3 11 1 13 1 15 9 7 9 0 7 9
9 3 1 9 3 13 1 9 7 9
14 1 15 9 13 15 1 15 1 9 3 13 9 1 15
8 7 0 13 15 9 7 9 0
6 11 3 13 1 9 3
15 13 3 9 1 9 9 7 3 13 15 13 11 1 9 15
13 13 3 15 9 15 13 1 9 7 13 1 15 13
6 0 3 13 15 15 13
4 3 13 15 9
8 7 3 1 0 0 13 15 13
5 3 15 1 15 13
3 11 3 13
10 7 13 3 9 12 15 15 13 15 13
7 1 9 3 0 13 1 15
3 13 3 11
5 9 3 13 15 13
7 7 3 3 15 13 13 9
16 7 13 15 9 13 1 11 7 13 11 9 0 3 13 15 16
10 3 16 3 13 9 12 9 13 15 15
7 7 13 3 11 13 15 3
6 7 13 15 13 1 9
4 13 15 15 13
7 7 15 0 13 13 1 15
19 7 16 13 9 13 15 9 0 7 9 7 9 7 13 15 1 9 15 13
6 16 15 13 11 13 15
3 13 3 15
6 16 15 13 3 13 9
10 16 3 7 13 15 3 13 15 7 13
6 15 3 13 3 9 0
5 0 3 1 15 13
5 15 13 16 15 13
3 0 3 13
4 15 3 13 9
6 0 3 13 1 9 15
9 7 13 15 9 15 13 15 1 11
6 13 3 1 15 13 13
5 11 3 13 15 13
5 15 3 13 9 9
5 0 3 13 13 15
2 15 13
8 11 3 13 1 9 7 1 9
7 15 9 3 13 1 9 0
17 0 3 13 15 13 16 13 9 13 1 15 11 13 1 11 1 3
29 11 3 13 11 13 15 16 9 0 13 7 13 16 1 9 0 13 13 15 1 11 13 3 0 1 11 1 9 0
5 13 3 15 9 0
6 0 3 15 3 13 15
9 13 3 9 7 9 3 13 1 15
19 13 3 15 11 1 9 15 7 13 15 13 15 1 9 0 13 15 1 11
13 13 3 0 9 11 3 7 11 1 0 9 1 15
7 3 3 13 9 13 1 15
11 11 3 13 9 7 9 7 9 13 1 15
19 7 6 15 13 1 15 3 13 3 12 3 1 9 0 9 15 1 15 13
14 13 3 15 1 15 7 6 15 0 9 13 13 1 15
4 13 3 13 15
9 9 3 13 1 15 9 13 15 12
5 13 3 15 9 13
2 13 0
4 13 3 15 11
7 3 3 11 13 13 13 11
4 0 3 13 13
1 13
6 0 3 3 13 1 15
4 15 3 13 0
6 15 0 9 13 1 15
4 13 15 3 13
6 11 3 13 13 9 15
17 13 3 15 13 1 9 1 9 7 9 15 13 7 11 13 9 15
17 7 16 15 13 13 11 15 9 13 1 9 13 15 9 13 1 11
7 13 3 15 11 1 15 13
7 9 0 3 13 15 1 15
14 3 15 13 15 7 9 15 16 6 9 13 1 15 13
12 0 9 7 9 15 3 13 7 9 15 3 13
3 13 1 15
2 7 9
2 13 15
11 3 16 1 0 9 0 13 1 0 15 13
20 7 3 13 1 9 13 0 3 13 15 7 9 0 3 1 0 7 0 1 0
3 11 3 13
3 9 13 15
6 13 3 9 15 13 9
4 7 13 9 13
8 13 3 15 3 9 13 1 15
3 15 13 13
11 3 13 3 15 16 0 13 11 9 0 13
8 16 15 13 9 0 13 15 0
13 13 3 3 9 13 1 15 9 0 7 0 7 0
8 12 3 1 13 9 13 15 13
9 16 15 13 11 13 15 0 7 15
6 13 3 0 13 15 13
11 3 3 15 13 15 9 16 1 0 9 13
5 7 15 3 1 9
5 0 3 9 15 13
3 7 13 11
4 7 13 15 11
3 6 13 15
6 3 1 15 13 1 9
17 13 3 3 9 0 7 9 13 1 15 9 1 9 0 7 13 9
7 7 9 0 13 15 1 12
6 7 13 9 0 11 13
7 9 1 9 15 13 9 15
6 1 9 9 0 0 13
14 7 15 13 9 1 9 0 13 13 13 9 15 13 15
15 13 3 15 13 15 3 7 9 13 1 15 1 11 13 0
11 7 6 9 9 11 9 13 9 0 7 0
18 0 3 13 13 9 7 9 15 1 11 9 0 15 13 3 0 9 0
26 0 13 1 11 13 9 0 7 13 15 13 15 9 7 13 15 1 9 13 1 15 3 13 15 3 13
7 7 9 13 9 7 9 13
20 1 9 3 13 9 15 13 13 1 15 1 11 13 9 7 16 13 13 9 15
7 7 1 9 3 13 1 9
17 1 15 3 9 3 3 13 1 9 13 15 13 9 7 0 1 15
13 13 3 9 13 1 9 7 13 3 13 9 9 11
18 7 13 13 15 15 1 0 7 6 9 12 13 1 15 1 9 13 15
12 0 3 13 15 7 13 9 1 9 13 1 15
5 15 13 0 1 0
4 13 3 7 13
10 13 3 13 15 3 13 1 11 13 16
19 13 3 11 9 7 11 7 11 0 7 0 1 15 15 3 13 1 9 0
14 7 13 15 1 15 3 9 9 15 7 3 13 15 9
19 11 3 13 13 1 9 7 13 13 9 12 13 7 13 1 15 13 15 13
31 7 6 12 1 15 13 13 1 0 9 1 9 13 9 12 12 1 11 15 9 11 7 0 13 1 15 1 15 0 13 15
15 7 13 13 15 7 13 15 7 0 11 13 15 13 1 15
9 9 3 15 13 15 16 15 3 13
4 13 3 1 15
3 7 13 0
14 15 3 12 9 13 1 11 7 3 13 13 1 9 0
3 7 13 15
1 15
4 0 3 13 15
31 15 1 11 9 15 13 9 9 0 9 7 9 1 9 7 15 9 7 3 15 13 9 7 9 15 1 9 9 7 13 15
10 15 3 13 15 16 0 13 13 11 13
8 7 7 9 15 1 15 13 15
19 13 3 1 9 7 3 13 9 15 13 13 3 9 9 13 15 13 15 0
5 7 0 13 1 15
11 6 0 7 0 9 13 1 15 15 13 9
11 3 3 3 13 13 11 7 13 1 9 15
15 7 13 1 11 7 1 15 9 13 15 9 15 13 1 15
14 7 13 15 1 9 1 15 13 7 0 13 15 3 13
13 13 1 15 16 1 9 13 7 13 15 13 3 9
5 7 13 1 15 13
13 7 13 16 13 1 15 13 9 13 7 13 13 15
5 7 0 13 1 15
4 7 13 1 15
19 3 9 3 15 13 13 1 15 3 13 1 15 1 9 7 16 13 15 9
31 7 13 1 0 9 13 15 1 11 7 13 13 15 12 1 12 7 15 13 1 15 13 1 9 16 13 11 7 13 15 11
10 0 3 15 13 0 11 13 1 9 15
9 13 11 1 0 13 1 9 9 15
3 7 13 15
2 9 15
3 3 13 15
9 13 3 15 7 0 13 13 9 13
3 7 13 15
8 7 1 15 9 13 1 9 15
10 13 9 15 7 9 15 16 0 15 13
15 13 15 7 13 16 9 9 7 9 3 13 3 15 13 13
8 7 0 13 13 15 9 7 9
12 3 3 3 13 15 1 9 7 13 15 13 15
11 0 3 13 15 9 13 9 7 1 9 9
5 7 13 1 15 13
3 13 3 15
26 0 13 9 15 13 1 15 3 13 1 15 16 13 13 15 15 13 1 9 0 7 9 7 9 1 15
7 3 13 15 9 16 13 9
34 7 13 15 16 3 13 13 7 3 13 13 11 7 13 1 0 0 9 7 13 15 1 9 15 9 7 9 9 1 15 9 13 1 11
5 15 3 13 9 0
9 7 6 15 13 9 9 15 1 15
12 13 3 15 3 1 11 7 13 9 15 13 15
21 7 0 13 15 15 13 15 1 11 1 9 0 7 13 3 1 9 13 7 13 9
1 6
7 13 9 0 3 13 11 9
5 7 13 13 1 9
6 7 13 15 7 13 15
11 15 3 13 16 15 13 11 7 11 7 9
4 13 15 11 13
18 0 13 13 1 15 15 1 15 13 15 15 13 0 16 13 9 9 15
12 0 1 11 13 1 0 9 11 3 13 11 13
10 1 0 9 13 11 13 1 15 7 13
7 6 9 0 13 9 9 15
6 0 13 1 15 15 13
12 1 15 13 9 15 1 15 13 16 0 15 13
17 7 15 3 13 15 7 16 13 15 11 0 1 15 13 1 9 13
5 7 13 11 13 16
4 7 13 1 15
14 7 15 3 13 15 7 13 15 13 1 9 0 15 13
14 1 15 13 9 13 7 13 1 15 0 13 13 9 0
10 7 15 13 7 13 16 0 13 9 0
16 1 0 3 9 3 13 11 7 1 9 15 12 7 13 11 13
1 13
3 6 9 0
10 7 13 15 12 9 13 7 1 11 13
4 0 3 13 15
8 9 15 13 15 13 9 3 13
2 13 15
3 13 7 13
12 13 3 7 13 3 13 7 13 1 15 9 0
4 9 13 3 0
16 13 3 11 9 11 11 12 1 12 13 1 11 7 1 15 13
3 7 13 15
5 7 13 15 1 11
6 13 3 1 15 11 13
5 15 13 11 9 0
8 15 13 15 11 15 13 15 11
12 1 0 3 9 13 11 13 1 11 7 13 11
4 7 13 15 11
10 13 3 11 1 11 1 9 0 7 0
6 13 11 11 7 13 15
4 7 13 15 11
7 1 11 13 3 15 0 13
4 7 13 15 11
3 13 7 13
7 13 3 11 11 13 1 15
8 6 1 9 9 1 15 9 13
3 13 15 11
3 3 15 13
11 3 16 3 13 15 11 13 1 9 13 15
5 13 11 7 13 15
6 9 7 15 13 9 0
4 15 13 9 0
9 16 13 15 16 13 15 1 9 13
3 0 0 13
3 7 13 15
4 6 6 13 15
14 7 1 0 9 9 13 1 11 0 7 13 9 0 3
10 13 3 13 7 11 7 9 15 1 9
8 7 13 9 13 9 0 1 15
3 13 15 11
6 15 13 15 7 15 9
5 3 3 13 9 15
4 13 9 15 9
5 15 3 13 15 13
3 13 15 11
3 13 9 9
3 7 13 15
5 13 3 7 13 9
2 7 13
24 16 3 13 9 9 13 1 9 7 3 13 3 13 7 9 13 13 9 13 9 9 7 13 15
12 0 9 3 0 9 13 7 3 13 15 3 0
6 15 3 13 0 9 3
22 1 0 13 11 1 11 0 7 9 15 7 9 15 7 9 15 7 3 3 0 9 13
37 7 13 1 9 13 9 7 9 7 9 7 9 13 7 13 9 1 9 15 13 1 9 9 3 7 9 7 9 13 9 7 9 13 7 13 9 13
3 13 0 3
7 3 13 9 9 15 9 0
7 13 3 9 15 16 13 13
5 9 9 15 13 15
6 13 3 9 7 13 15
7 15 9 13 15 16 0 13
3 13 3 9
16 12 12 7 12 9 13 13 9 0 7 15 3 12 9 13 15
7 0 3 13 1 9 9 15
20 3 3 13 1 0 13 9 15 16 0 13 7 9 13 9 7 9 15 13 11
19 3 3 13 1 11 1 9 1 9 0 13 1 9 15 13 9 15 15 13
22 0 3 11 3 13 15 1 9 15 16 0 13 15 7 16 3 13 16 15 13 1 9
7 0 3 13 15 13 1 9
10 13 3 9 1 9 11 9 15 9 0
3 7 13 15
8 9 13 16 1 9 13 13 9
16 15 3 3 13 9 0 13 15 15 13 16 3 13 9 1 15
5 13 11 7 13 15
4 6 6 13 15
11 16 15 3 13 15 3 3 13 13 9 0
4 13 1 15 11
7 3 13 9 13 15 0 13
3 6 13 15
14 16 15 3 13 15 9 7 9 3 13 13 1 9 0
11 13 1 9 9 13 7 13 1 9 9 13
6 3 13 15 16 13 15
5 13 15 13 15 3
16 9 3 13 13 7 9 15 13 7 3 13 3 13 7 3 13
6 3 13 0 13 1 9
4 3 13 0 13
4 15 13 9 0
5 7 0 3 3 13
17 6 6 13 15 16 15 13 13 7 15 13 13 7 9 15 3 13
13 16 0 13 15 7 3 13 3 16 13 15 0 13
14 7 15 13 1 9 3 13 1 9 9 0 13 1 9
24 7 3 11 13 9 1 9 3 13 15 13 9 0 16 0 13 1 15 3 13 7 13 9 0
17 3 13 3 9 9 15 1 9 16 13 9 7 16 13 15 9 15
6 13 1 15 3 13 13
3 0 13 9
12 13 3 9 1 9 7 13 9 3 9 3 9
5 13 3 15 9 0
20 0 3 13 0 13 9 7 3 13 1 9 16 3 13 15 9 15 16 0 13
16 7 13 9 13 1 9 16 13 15 9 15 16 1 9 13 13
18 13 3 11 13 1 11 1 11 16 9 0 13 3 7 13 7 13 15
8 3 3 3 13 13 1 9 11
10 13 3 9 1 9 0 1 9 1 9
20 9 15 13 1 15 1 0 9 11 15 15 13 6 0 13 7 15 13 1 15
4 13 11 7 13
12 3 13 9 13 15 16 3 13 15 13 1 9
6 15 0 15 13 16 13
4 13 9 9 13
13 7 9 0 13 7 13 15 9 13 15 1 9 0
6 0 3 9 15 13 15
7 0 13 13 7 15 13 15
10 13 1 9 1 9 13 7 1 9 13
19 13 1 9 1 15 13 7 15 13 7 13 0 13 7 9 15 15 3 13
8 13 15 9 13 16 9 0 13
7 3 1 9 3 9 13 9
9 9 13 9 7 15 13 1 9 15
6 13 1 9 13 9 0
15 7 15 3 13 1 9 3 13 9 7 9 0 13 1 15
31 3 3 13 9 16 13 9 16 11 0 9 13 7 13 3 11 7 11 0 3 13 7 9 15 13 11 7 13 3 1 11
16 13 3 11 1 9 0 13 11 1 9 15 13 11 11 9 15
5 13 3 3 9 0
4 9 13 3 0
6 13 9 1 11 13 9
2 13 11
3 13 15 13
10 9 3 15 13 13 1 9 16 9 13
5 13 3 15 9 9
6 3 13 3 15 9 9
24 16 13 13 9 0 7 15 13 13 15 13 15 13 15 13 13 1 15 7 13 15 13 9 0
3 13 15 9
4 9 3 9 13
4 7 9 13 0
5 3 3 13 9 0
12 3 15 0 13 9 15 11 15 13 15 9 0
11 7 0 1 15 13 7 9 15 7 9 15
29 7 15 13 1 9 15 15 13 15 3 13 15 1 9 7 9 15 15 13 15 13 1 15 9 9 13 1 9 0
4 13 1 15 9
12 9 13 15 0 9 16 7 13 7 13 3 13
3 13 15 11
1 13
6 13 9 15 7 13 3
5 13 9 7 13 15
3 3 13 9
3 3 13 16
3 9 3 13
12 12 3 9 13 13 7 3 15 13 13 15 9
4 0 1 9 13
3 13 15 9
6 9 13 16 9 13 15
7 9 15 1 9 0 13 15
12 7 15 13 16 1 11 13 9 3 13 15 13
6 15 13 15 15 3 13
11 15 3 13 15 15 13 16 9 1 9 13
15 7 13 9 7 3 13 3 0 9 13 15 9 9 7 9
7 3 9 0 13 13 15 15
14 9 13 9 7 15 13 15 15 9 7 9 13 13 15
3 13 15 9
6 13 16 11 13 13 11
3 13 15 11
12 7 3 13 9 15 7 13 15 16 1 9 13
7 7 15 3 13 15 13 7
4 15 13 1 15
12 13 3 9 15 9 7 13 1 9 7 13 9
10 13 7 13 9 15 13 15 15 15 13
4 3 0 13 11
8 1 3 0 13 15 9 15 13
2 9 13
8 15 9 13 13 15 15 3 13
5 13 3 9 1 15
5 3 15 13 15 13
3 13 15 11
12 15 9 13 16 13 9 13 15 7 13 9 15
3 6 13 15
12 13 9 15 7 13 9 16 0 13 1 9 3
18 7 13 9 13 7 13 9 1 9 0 16 7 13 3 13 15 7 13
9 15 13 15 13 3 15 3 13 15
9 15 13 15 7 15 1 9 15 13
15 1 9 3 0 0 13 1 15 1 9 1 9 9 13 16
5 13 15 15 15 13
5 7 13 3 12 9
7 7 3 3 13 1 9 15
4 9 3 13 16
6 3 3 1 15 9 13
10 1 12 3 9 13 3 7 13 1 11
12 0 3 11 13 16 9 1 15 9 3 13 9
16 3 3 13 1 11 13 15 9 15 13 15 13 1 11 1 9
12 13 3 3 11 1 11 11 3 13 1 9 9
10 13 3 15 0 9 15 9 13 1 11
21 0 13 16 11 13 1 11 1 11 13 1 15 7 13 15 16 13 7 13 9 15
3 13 3 13
5 13 3 1 15 11
5 13 1 15 0 9
8 9 13 3 16 3 13 9 15
1 13
4 9 15 0 13
10 7 9 13 9 9 15 13 15 11 13
15 3 3 13 15 6 9 15 13 15 13 16 9 15 0 13
10 13 3 9 1 15 1 15 3 15 13
4 13 3 15 16
13 13 3 9 16 0 13 9 1 15 13 15 11 16
7 7 13 0 7 15 9 15
11 6 3 0 9 13 11 13 1 11 1 11
11 1 0 3 13 9 0 7 13 11 1 11
15 13 3 1 11 1 0 9 15 13 15 3 11 12 9 13
11 1 0 13 9 13 0 0 0 13 9 9
26 9 3 0 1 15 9 13 1 9 7 13 9 7 15 3 13 1 9 9 0 13 15 3 9 13 13
13 13 3 3 15 9 12 7 12 9 13 1 9 15
3 13 15 0
15 6 9 9 3 3 13 16 3 13 15 9 13 15 1 9
8 3 3 13 15 15 1 15 13
3 13 15 11
1 13
8 13 9 15 7 13 1 9 15
11 7 3 0 13 9 7 13 9 15 7 13
6 13 3 9 1 0 9
9 9 13 7 3 13 15 13 9 15
4 0 3 13 15
7 15 15 13 0 0 15 13
5 13 9 15 7 13
3 13 3 15
5 15 13 9 13 15
5 13 9 15 7 13
6 13 3 3 13 15 13
3 7 13 15
3 6 0 13
9 1 0 3 13 16 3 0 15 13
13 13 3 9 7 13 9 16 11 13 15 15 13 0
15 7 0 1 13 9 11 7 13 15 13 16 0 13 1 9
4 11 3 13 15
7 9 15 3 13 7 15 13
6 13 3 11 7 13 15
13 3 13 9 1 15 13 15 3 3 15 13 9 13
9 15 3 0 13 0 3 9 3 13
21 9 3 13 9 7 15 13 15 15 0 13 7 0 0 13 15 9 16 15 13 15
13 3 3 9 13 0 7 13 3 3 9 15 13 13
17 9 3 3 13 15 7 9 15 13 9 16 15 13 9 3 13 9
10 7 15 3 13 9 3 13 9 13 15
19 6 6 13 15 16 13 9 7 3 13 3 0 13 9 9 0 7 13 13
15 3 3 9 9 13 1 15 3 13 3 9 9 13 1 15
30 3 13 15 0 16 13 9 1 15 15 13 1 9 13 9 9 0 7 13 13 0 1 9 9 7 13 0 1 9 9
7 3 13 15 1 15 13 15
18 3 13 13 7 9 15 0 13 16 3 13 9 15 7 9 13 15 9
9 16 15 13 1 15 9 15 13 0
15 15 13 13 1 15 7 13 16 0 13 9 15 13 1 15
14 15 3 3 1 9 9 13 7 0 13 16 15 13 13
6 0 13 9 13 7 13
9 15 3 13 13 15 1 9 9 15
20 9 3 15 13 15 9 16 13 15 0 9 15 13 13 1 15 16 9 15 13
8 7 13 15 9 0 13 1 15
9 7 9 15 3 13 7 9 15 13
17 7 9 15 3 13 13 1 15 16 15 0 13 0 15 9 3 13
6 7 0 13 13 1 15
9 7 3 13 13 1 15 16 9 13
15 9 1 9 3 13 7 13 15 16 9 0 3 13 1 15
10 15 13 1 9 9 15 7 3 13 15
17 3 15 13 13 9 15 1 15 13 7 9 15 1 12 9 3 13
9 3 13 16 15 1 15 13 1 9
10 13 15 1 15 13 11 1 15 15 13
5 1 15 3 0 13
12 16 3 0 9 9 3 13 3 15 9 9 13
10 1 0 13 11 1 0 9 9 11 0
13 7 1 15 13 9 0 16 13 9 15 13 1 0
11 13 3 1 9 11 7 3 13 1 9 15
14 13 3 9 11 13 16 0 9 13 1 15 13 1 11
6 15 13 9 16 13 0
6 0 3 13 15 13 13
3 13 15 11
13 12 12 9 9 3 13 15 16 15 15 0 15 13
10 13 15 15 1 9 15 11 9 11 11
12 13 9 3 15 15 13 12 9 0 7 12 9
6 7 0 15 13 1 0
3 13 9 13
7 13 3 9 9 3 12 12
18 13 3 9 11 7 9 13 13 9 7 9 13 3 7 1 9 15 13
7 7 16 13 15 13 9 15
7 13 9 9 16 3 13 15
16 13 3 7 13 12 1 12 9 9 1 12 9 0 15 13 13
9 9 3 13 9 15 13 11 13 16
9 0 13 1 9 9 13 1 15 9
12 7 9 3 13 7 3 3 13 13 1 15 11
6 9 3 9 0 13 13
23 13 3 3 12 12 7 12 9 7 12 0 13 11 13 1 9 7 1 9 13 7 13 15
4 0 3 13 15
2 15 13
3 3 13 15
15 13 3 15 13 1 9 7 3 13 9 1 9 1 15 13
40 1 0 9 9 15 13 1 0 9 9 13 16 9 15 3 13 3 3 12 0 1 15 13 9 15 7 16 3 13 1 9 15 11 1 9 7 12 9 15 13
22 3 3 13 9 16 11 3 13 3 7 9 15 13 0 1 9 7 13 1 11 13 11
9 7 13 15 1 0 9 9 13 15
4 9 3 3 13
5 13 15 11 7 13
4 6 6 13 15
14 13 15 3 16 13 9 7 16 13 13 9 7 13 15
15 13 3 9 13 7 9 13 1 9 0 15 9 0 15 13
5 0 3 9 13 9
5 13 11 7 13 15
11 0 13 9 0 16 13 1 0 15 13 0
3 13 3 15
11 15 3 15 13 9 16 13 7 9 13 15
2 15 13
9 9 15 13 9 1 9 3 13 13
6 9 1 9 13 15 13
4 6 6 13 15
11 9 3 0 13 13 1 9 7 13 9 9
4 13 3 1 15
6 9 3 13 15 9 0
4 13 3 15 11
4 15 13 9 0
16 13 1 15 3 13 13 15 7 13 1 15 3 13 13 15 3
28 15 15 13 15 9 1 15 13 7 13 1 15 3 13 3 16 13 1 9 16 3 13 9 15 7 9 13 15
22 0 3 13 9 13 15 9 16 0 15 13 15 3 13 1 15 7 13 15 1 0 9
7 13 3 9 1 15 16 13
6 15 13 9 13 1 9
2 7 13
13 3 0 3 13 11 9 0 15 15 13 9 7 9
5 3 3 0 13 16
5 13 11 7 13 15
4 3 13 1 15
20 15 3 13 13 1 15 16 3 9 13 15 13 15 7 15 13 15 1 0 9
5 7 13 15 13 9
8 0 13 9 7 13 13 1 15
6 3 3 9 13 13 3
4 3 13 1 9
4 6 6 13 15
6 13 1 15 13 9 0
4 15 13 9 0
8 9 15 13 9 1 9 7 13
7 15 13 9 0 13 1 9
10 16 15 13 1 9 0 0 13 1 9
14 9 3 15 15 13 9 15 13 15 15 13 1 9 9
8 3 13 0 13 9 15 13 15
4 13 3 15 11
4 6 6 13 15
15 16 3 13 9 9 0 7 13 9 15 9 3 13 1 15
17 13 15 9 7 13 15 9 13 9 0 7 15 13 15 1 0 9
14 13 15 9 7 13 15 9 1 15 13 7 15 1 15
10 3 13 15 13 9 3 15 13 9 1
7 13 9 0 0 13 1 9
7 0 13 1 9 13 1 11
7 0 3 13 1 9 15 13
4 0 13 9 0
4 15 13 15 13
13 13 3 11 1 15 16 13 1 0 9 15 13 15
9 16 3 13 9 0 13 3 13 3
5 1 9 13 9 15
10 9 15 15 13 15 9 13 7 9 13
8 7 13 1 15 15 15 3 13
14 13 3 3 11 15 13 3 13 7 15 13 13 13 15
2 7 13
19 0 1 13 15 16 15 3 13 13 1 15 16 3 13 13 15 1 9 15
15 1 0 0 1 9 15 13 3 7 1 0 3 13 1 15
4 13 15 11 11
4 9 1 15 13
4 9 9 0 13
12 7 15 13 7 13 16 15 13 11 9 9 0
3 13 15 11
8 3 15 3 15 12 1 12 13
6 7 1 15 12 9 13
5 13 3 11 0 11
7 7 13 1 0 11 1 11
11 3 13 3 1 11 13 16 13 15 9 13
6 13 3 1 9 0 9
6 13 3 1 15 9 15
15 13 3 7 13 1 11 16 3 9 15 13 9 15 15 13
11 15 3 1 9 15 13 7 13 0 3 13
7 16 0 13 13 15 15 9
7 3 9 3 15 13 1 15
5 3 13 9 13 15
13 15 3 13 16 15 13 1 15 16 9 15 0 13
5 15 13 1 9 0
13 15 3 13 1 9 0 16 9 15 3 3 13 15
6 0 13 0 13 1 11
16 3 3 13 9 15 1 9 3 3 0 13 3 3 7 3 3
6 9 3 13 15 1 9
3 3 13 0
5 0 13 16 0 13
3 15 3 13
4 3 7 13 9
9 15 3 3 13 1 15 9 1 0
11 3 3 1 9 9 13 11 1 9 7 13
5 7 13 15 9 13
6 13 3 11 7 13 15
7 15 9 13 15 7 13 15
6 13 1 15 9 15 13
13 7 13 9 13 15 0 0 13 7 13 9 1 15
6 3 11 3 13 15 9
6 7 15 1 15 13 9
4 15 15 13 13
3 9 3 13
4 15 15 13 13
5 13 11 7 13 15
19 0 1 11 13 15 9 3 16 1 11 13 7 1 9 7 1 9 13 9
24 16 9 13 9 1 9 16 3 13 15 9 0 1 15 3 13 15 16 15 9 0 13 1 9
8 3 13 1 9 7 0 9 13
5 13 3 15 1 9
11 7 6 3 13 15 13 7 15 15 3 13
8 3 3 13 9 16 0 13 11
5 7 0 13 3 13
9 7 11 3 13 15 3 13 3 13
7 7 15 13 7 13 3 13
14 7 1 15 3 13 7 13 0 13 15 15 15 3 13
11 15 15 13 16 1 15 13 7 0 15 13
10 1 9 3 0 13 1 15 7 13 16
11 11 3 13 3 0 9 13 15 0 13 13
17 13 3 9 9 13 1 15 0 7 13 9 7 9 9 16 13 15
3 13 3 11
11 3 0 9 1 15 13 7 13 1 13 15
6 13 3 9 1 15 0
8 3 13 13 16 15 3 13 15
4 15 13 9 0
13 13 15 7 3 13 7 3 13 15 15 3 13 13
11 1 0 3 9 0 9 13 11 7 13 13
9 16 15 13 3 13 1 15 7 13
13 13 1 15 3 9 13 9 1 9 15 13 9 0
11 0 3 13 1 9 15 13 13 13 1 15
8 0 3 1 9 13 9 0 13
2 0 13
3 0 13 11
2 0 13
5 3 1 11 11 13
10 3 9 3 13 16 1 9 0 13 11
7 9 3 13 1 9 15 1
14 15 3 1 15 13 15 13 7 15 3 13 1 15 9
2 13 9
8 3 3 13 13 9 3 0 9
3 13 15 9
5 3 3 15 13 13
10 3 15 1 9 13 1 15 7 1 9
9 7 9 0 15 3 13 9 13 13
12 13 1 15 11 13 1 15 9 12 13 1 15
15 3 9 15 13 9 16 3 13 1 15 3 7 13 15 13
6 3 3 15 1 11 13
9 13 7 13 16 1 11 9 3 13
6 11 3 13 1 9 0
6 3 3 3 13 1 9
10 7 15 9 13 1 15 7 13 13 15
9 13 3 9 7 9 9 1 9 13
7 7 13 15 1 9 13 15
8 9 0 9 13 13 3 1 9
12 0 3 13 13 15 16 13 13 1 15 15 13
9 11 3 3 13 15 9 13 1 9
10 16 3 13 13 15 13 15 7 13 15
10 15 15 1 9 13 3 13 9 1 15
7 7 3 13 15 13 1 9
12 0 3 13 13 12 1 12 13 1 9 1 0
9 7 13 11 12 7 9 13 1 9
7 9 3 13 15 1 15 13
3 0 3 13
2 15 9
3 13 15 11
4 3 15 15 13
7 13 7 3 3 13 1 0
6 3 3 15 13 11 13
12 13 1 15 3 13 13 1 9 7 13 9 0
4 13 3 15 9
4 9 15 13 0
5 13 11 7 13 15
17 16 15 13 1 15 0 9 15 0 13 16 13 3 13 7 3 13
9 15 3 3 13 3 13 7 3 13
4 15 1 9 13
17 16 3 13 15 9 15 0 13 16 12 13 7 15 7 13 15 9
13 7 1 9 3 15 13 13 16 12 9 9 0 13
13 15 13 13 1 15 0 7 13 1 15 13 15 9
4 3 13 9 15
2 13 11
6 7 15 13 7 9 15
9 16 15 13 13 3 9 15 13 13
12 7 15 3 13 15 16 3 3 13 13 9 15
5 13 3 15 3 11
10 15 13 7 13 15 7 1 9 15 13
7 3 15 13 15 3 13 13
6 3 15 0 13 16 13
7 3 15 13 15 3 13 13
3 7 13 15
4 15 1 0 13
5 15 1 0 9 13
5 15 13 1 0 9
8 13 3 15 16 13 1 9 15
12 16 3 9 3 13 16 15 13 13 1 9 15
3 15 15 13
4 7 13 15 11
7 0 13 1 15 13 7 13
15 7 13 15 0 13 7 15 15 13 1 15 0 13 1 9
7 7 3 13 16 9 15 13
4 13 3 15 11
23 3 13 9 0 3 13 16 15 13 7 1 15 15 3 13 7 3 13 15 9 15 0 13
6 7 13 15 1 15 13
7 0 13 15 0 13 1 15
11 16 15 13 1 9 15 1 9 9 15 13
7 7 13 9 7 9 13 15
3 13 15 9
8 9 0 13 7 15 3 13 3
4 3 15 13 16
2 0 13
3 13 15 11
8 7 9 3 13 1 9 1 9
5 9 3 13 1 9
9 16 3 9 15 13 1 9 0 13
5 13 16 9 0 13
7 15 15 13 1 9 15 13
9 7 15 3 15 13 1 9 15 13
4 13 7 13 15
4 9 15 11 13
9 16 9 0 13 13 9 0 13 13
14 3 3 13 15 13 9 15 9 15 13 15 13 1 9
4 0 11 13 13
5 15 13 9 9 15
3 13 3 15
5 15 1 9 13 13
4 12 9 13 9
4 13 3 15 11
9 3 1 15 3 13 7 0 15 13
6 1 15 9 15 3 13
6 3 3 13 13 9 15
5 15 1 9 9 13
6 7 9 9 15 13 13
14 0 9 13 3 7 1 9 3 13 16 13 9 1 15
12 3 13 9 1 15 13 16 0 13 7 9 15
7 15 1 15 13 15 1 9
7 15 13 1 9 9 0 13
8 0 15 3 13 16 13 1 9
5 13 9 7 13 15
12 3 3 3 13 15 16 9 13 15 7 9 13
2 13 11
4 15 9 3 13
6 15 3 3 13 9 15
4 13 13 7 13
11 16 15 9 15 13 9 3 13 13 1 9
4 13 3 15 9
5 3 13 16 9 13
8 11 13 7 9 7 15 13 16
11 16 15 9 15 13 3 13 13 9 1 9
3 7 9 13
5 15 15 0 15 13
2 13 11
12 13 9 15 13 15 15 15 13 16 9 15 13
4 7 3 13 15
4 15 3 13 15
11 7 16 13 16 3 13 15 13 0 15 0
16 11 9 15 0 13 13 16 13 13 9 15 7 13 7 13 15
5 13 3 9 1 15
11 12 12 9 3 3 13 7 11 3 13 13
3 13 15 11
7 3 16 3 13 11 15 13
7 13 3 9 16 13 1 15
16 11 3 13 15 7 13 1 9 7 13 1 9 15 13 7 13
6 7 13 15 9 15 13
12 9 15 13 0 3 7 9 15 16 0 13 15
2 13 11
14 7 0 13 7 9 15 7 16 13 15 9 0 1 15
9 15 13 13 9 13 15 16 9 13
7 3 1 9 13 9 13 9
18 0 13 13 1 9 7 13 9 1 9 7 13 15 9 9 7 13 15
9 13 15 1 9 0 15 13 15 13
8 13 3 7 13 15 7 13 13
12 9 3 7 15 15 13 13 3 16 0 13 13
7 3 0 3 13 13 7 13
5 0 13 16 0 13
4 0 3 13 16
3 13 3 15
4 13 0 7 13
5 9 13 11 9 13
7 7 13 9 15 7 13 15
7 13 1 9 0 7 13 15
6 13 3 7 13 15 13
3 13 3 15
3 3 0 13
8 13 15 1 9 15 13 3 0
11 13 3 9 3 13 9 11 7 13 15 9
7 3 3 13 15 9 3 13
4 0 3 13 15
10 9 13 15 1 9 7 13 15 7 13
5 13 3 1 9 15
9 13 0 1 9 9 16 9 3 13
2 0 13
5 7 9 13 1 15
3 13 9 3
9 15 15 13 1 15 16 13 9 15
6 0 3 13 16 9 13
21 3 13 3 9 9 1 15 16 13 0 7 13 16 13 9 0 13 7 13 15 13
12 0 3 13 9 15 15 15 13 16 0 15 13
4 3 3 3 13
7 13 3 15 9 15 7 13
2 0 13
2 9 13
5 0 1 15 3 13
8 3 13 9 15 16 13 15 9
14 3 3 15 13 13 9 16 16 15 13 11 13 9 13
6 0 1 9 15 13 16
2 9 13
10 13 3 3 9 15 13 0 7 13 15
7 15 13 16 9 0 0 13
5 13 3 0 7 13
5 16 9 13 3 13
8 12 13 16 0 13 3 3 13
4 13 3 15 3
3 15 13 15
6 13 15 3 7 3 13
4 15 13 3 13
6 0 3 13 15 7 13
4 15 9 13 0
5 15 3 0 13 9
6 15 13 16 11 13 9
6 0 3 3 13 3 13
15 1 0 3 0 13 16 15 3 13 3 13 7 13 9 15
18 13 3 16 9 9 3 13 7 16 15 9 13 7 9 15 13 0 13
10 1 9 13 13 16 15 13 9 0 13
4 13 7 13 15
12 1 9 15 13 15 13 15 7 15 3 15 13
4 7 13 15 3
11 13 11 16 13 15 3 7 13 15 13 15
4 13 0 7 13
8 15 13 9 16 9 13 1 15
4 13 3 15 11
9 13 15 13 7 13 1 15 0 13
2 13 9
4 7 13 15 15
3 7 13 11
11 7 13 0 1 9 13 1 15 7 13 15
5 3 3 15 0 13
4 13 3 15 11
8 16 13 0 13 3 13 13 9
4 3 3 13 16
4 7 9 15 13
4 6 6 13 15
6 7 13 9 9 13 9
17 0 9 13 7 9 9 15 13 7 15 9 13 1 9 7 13 15
17 7 3 15 9 13 1 15 13 7 9 1 15 13 16 13 9 15
14 1 0 3 3 13 7 13 1 15 16 3 13 0 9
5 0 9 13 15 11
9 0 3 3 13 15 13 15 13 15
4 6 6 13 15
15 15 3 15 13 1 15 9 13 7 9 7 3 13 15 9
3 15 13 9
13 15 16 15 13 13 15 7 13 7 13 7 9 13
10 9 3 13 7 16 13 7 13 7 13
8 15 13 16 9 13 7 0 13
4 15 13 9 0
7 9 0 9 15 13 1 9
25 15 13 9 0 7 13 15 7 13 15 15 3 13 15 9 7 15 13 9 7 9 15 13 1 9
10 7 15 9 13 15 3 13 1 9 0
16 3 0 15 13 13 7 9 15 13 7 13 12 9 7 12 9
14 0 1 15 9 13 16 15 13 9 15 16 3 13 15
11 15 13 15 1 15 7 15 13 15 1 15
10 9 13 13 15 7 9 13 3 13 15
6 0 9 13 1 9 15
9 9 3 13 3 1 9 1 9 0
5 9 13 7 0 13
3 15 15 13
2 15 13
6 0 9 3 13 13 15
6 3 9 13 0 9 13
6 13 3 3 9 1 11
3 7 9 13
8 7 13 11 1 9 1 9 0
9 16 15 13 11 13 15 3 13 15
3 13 15 11
5 13 15 7 3 13
12 9 15 15 13 1 9 9 15 0 13 1 15
4 7 15 3 13
8 13 3 1 9 15 3 13 15
32 9 15 9 15 13 7 15 13 15 7 1 15 13 7 15 9 0 13 15 7 3 13 1 9 7 3 13 15 15 1 9 15
5 15 7 9 12 13
3 13 15 11
9 0 9 0 13 1 15 1 9 15
8 1 15 15 9 9 1 15 13
4 13 15 9 13
20 1 0 9 3 13 9 1 15 7 1 9 7 16 15 9 13 13 15 0 9
3 13 15 11
2 15 13
2 9 13
10 16 3 13 9 9 15 3 13 15 9
25 16 3 13 16 3 15 9 3 13 9 15 9 13 16 13 7 13 16 1 15 9 7 15 1 9
11 7 13 3 15 3 13 7 13 1 9 15
17 7 13 3 1 0 9 11 1 9 3 13 11 3 13 7 13 3
8 7 0 13 1 15 7 13 16
9 15 3 15 13 11 1 0 9 13
6 7 0 13 1 15 3
13 13 3 15 13 11 1 11 9 0 7 11 9 15
7 13 3 9 15 1 15 13
5 9 6 15 13 13
4 13 3 11 13
15 0 9 13 1 9 7 1 9 0 16 13 15 9 0 15
14 3 3 13 16 13 3 3 13 1 15 13 9 12 9
5 1 0 3 13 9
4 13 1 11 3
4 13 15 9 15
2 13 11
9 3 12 3 1 12 9 13 1 9
13 16 15 13 1 9 3 13 15 16 9 9 0 13
7 0 13 7 1 0 13 15
4 11 9 15 13
5 7 13 16 13 15
4 13 3 9 15
5 9 16 13 13 13
8 0 3 13 16 1 9 9 13
7 3 13 15 11 3 13 15
4 7 13 1 15
7 13 3 11 13 11 1 9
7 13 3 15 16 13 1 15
13 13 3 11 1 11 13 15 12 9 3 13 1 9
10 13 3 11 1 11 3 12 1 12 9
16 7 0 1 9 13 13 1 11 7 11 16 13 15 1 9 15
4 7 11 3 13
10 9 16 13 3 13 3 13 9 15 13
13 7 3 3 13 16 15 3 13 1 9 13 15 9
3 13 15 11
3 13 9 15
3 13 15 11
8 13 16 13 1 9 1 0 9
3 13 15 11
11 7 0 0 7 13 1 15 3 13 1 9
4 13 3 9 0
4 13 15 6 9
12 15 13 16 15 13 11 9 0 13 1 15 9
11 7 0 13 13 7 13 11 9 15 3 13
6 9 6 13 7 13 15
10 0 3 16 13 13 3 7 13 1 15
18 3 13 3 3 3 11 13 1 9 7 13 1 9 3 3 13 15 11
15 11 3 16 13 3 13 11 13 15 13 15 1 9 13 15
10 9 16 13 13 3 3 13 15 9 13
16 11 3 16 13 15 13 15 7 13 1 15 9 13 15 13 9
6 7 13 15 0 7 13
3 3 13 15
2 13 15
2 9 13
1 13
4 13 3 13 15
5 15 3 1 15 13
13 3 13 3 0 13 9 0 13 16 3 0 3 13
9 11 3 3 13 1 15 13 1 9
8 13 3 9 7 9 13 1 15
2 13 11
2 13 9
3 9 3 13
3 13 15 11
10 3 13 3 15 16 16 13 13 9 0
7 13 3 9 3 13 13 13
7 11 3 13 3 9 7 13
7 9 9 15 13 16 13 15
7 15 3 13 16 3 15 13
6 7 0 13 9 0 13
3 11 13 3
5 7 9 15 9 13
3 13 15 11
7 13 15 7 3 13 15 13
15 0 3 1 9 13 1 11 7 13 15 13 11 13 1 15
13 15 3 1 15 13 1 9 7 13 15 15 13 11
8 15 13 16 9 0 9 0 13
19 16 13 15 3 15 9 13 1 15 7 13 9 7 13 7 9 7 9 15
12 15 3 15 1 15 11 9 13 9 0 13 15
32 0 3 1 15 3 13 7 9 13 9 0 13 16 13 11 13 1 9 7 3 3 1 9 7 3 16 9 0 13 13 1 12
9 1 0 3 9 13 16 15 13 13
26 11 3 1 0 3 3 13 1 9 7 13 3 1 9 1 9 1 11 13 9 7 3 13 1 9 15
17 13 3 1 9 0 7 13 0 1 11 1 9 1 9 16 13 15
11 15 15 13 15 16 3 13 3 13 1 9
17 13 3 9 7 9 9 16 16 15 13 15 3 13 13 16 13 15
17 11 3 1 12 9 9 13 1 11 3 13 11 13 15 13 1 0
8 13 3 15 9 3 7 11 13
11 11 3 13 9 9 9 9 0 13 9 0
6 7 13 9 15 9 15
7 9 3 13 15 1 9 0
13 15 1 9 0 3 13 13 1 12 9 7 13 0
18 0 13 3 16 1 0 13 15 7 16 9 13 7 9 13 7 13 13
3 13 3 11
3 3 13 15
6 1 9 9 15 13 15
24 13 3 9 0 1 9 16 3 13 7 13 3 11 1 3 7 16 3 11 13 15 13 1 0
17 13 3 9 16 3 11 13 16 0 15 1 13 9 7 13 1 11
3 7 13 13
8 6 0 13 1 9 0 9 0
10 13 3 11 9 13 1 15 3 13 13
5 3 13 15 9 0
8 6 9 15 13 13 1 9 0
24 0 3 3 13 9 15 3 7 3 13 15 11 3 13 16 0 13 1 15 13 7 0 13 15
13 0 1 3 3 15 13 9 16 13 15 13 0 9
5 13 16 3 9 13
6 6 15 9 1 15 13
11 13 3 9 15 1 13 16 13 15 1 9
10 0 3 13 1 11 15 13 1 11 0
4 7 13 15 13
4 9 13 11 13
5 13 11 7 13 11
7 13 9 16 13 15 9 0
4 6 6 13 15
11 16 9 0 3 13 13 1 9 0 12 13
6 16 3 13 0 9 13
17 13 9 15 13 15 7 13 9 15 1 9 0 1 9 0 13 15
17 16 15 15 13 1 15 3 13 7 3 13 15 3 3 9 15 13
8 7 16 15 15 13 13 15 9
8 3 9 15 13 15 7 15 13
7 7 0 1 13 1 9 0
4 9 13 9 15
5 13 3 9 1 9
5 7 13 7 3 13
6 9 3 13 7 13 13
2 9 13
2 15 13
3 9 13 15
5 3 9 13 9 0
7 3 9 9 0 13 13 3
11 7 15 16 13 13 1 9 15 13 1 15
8 0 3 13 13 15 9 13 13
3 13 15 9
13 15 13 1 9 16 11 13 1 9 7 3 15 13
5 13 15 13 9 0
4 13 3 15 11
9 13 16 9 13 16 9 15 3 13
8 7 13 1 9 3 13 3 13
10 16 9 13 13 1 9 16 9 9 13
9 0 13 11 7 13 13 15 1 15
19 0 3 9 13 15 1 15 3 13 1 15 16 13 15 9 11 9 15 13
6 9 15 9 13 9 15
9 0 1 3 13 13 16 3 13 11
21 13 9 15 7 13 13 9 15 16 3 13 9 7 13 9 7 13 15 7 13 15
20 3 3 3 1 9 0 13 1 15 7 9 1 3 13 16 3 1 9 13 13
8 13 3 3 9 0 3 9 0
5 11 3 13 7 13
11 13 1 15 3 13 1 15 7 1 13 15
6 7 13 15 13 13 15
14 7 16 15 13 9 15 7 3 13 15 15 3 13 15
10 3 13 3 16 13 9 7 16 13 9
11 13 15 15 7 3 13 9 15 13 13 15
19 3 15 1 15 3 13 7 13 15 9 0 15 9 13 15 13 7 15 13
8 7 13 16 9 15 9 0 13
10 15 3 15 13 3 13 15 9 3 13
27 1 3 9 9 13 11 16 13 15 9 16 13 1 9 0 1 9 13 15 13 1 15 9 1 9 13 15
18 1 0 3 13 9 1 9 7 13 13 9 9 7 13 9 15 13 13
5 13 3 1 11 11
4 7 13 15 0
6 9 15 3 15 13 9
7 15 15 13 15 3 13 3
4 13 3 1 0
3 13 15 11
3 13 15 11
9 16 3 13 15 3 13 9 1 15
4 13 15 11 11
10 9 3 9 15 3 7 3 9 7 9
3 13 15 11
4 13 3 15 0
7 7 15 0 13 7 3 15
4 0 1 13 16
4 3 15 13 0
14 3 3 13 9 15 13 9 15 7 13 3 7 13 15
5 13 3 15 13 15
9 15 13 15 9 7 9 7 3 13
2 13 3
12 9 3 13 15 16 3 15 13 15 3 15 13
10 13 9 0 9 15 7 9 0 13 15
8 16 0 13 0 13 16 13 15
5 3 1 15 15 13
5 15 3 13 15 13
5 7 16 9 13 15
9 13 1 15 9 13 1 15 9 15
15 3 13 15 3 16 3 13 16 3 13 9 13 16 15 13
10 0 13 11 13 15 9 7 13 7 13
10 6 6 13 15 16 12 1 15 13 15
10 13 3 15 1 15 9 13 1 15 13
13 13 3 12 13 1 9 15 1 9 0 15 13 11
6 13 3 0 11 11 13
6 15 3 13 1 15 13
9 13 3 0 3 1 9 0 13 15
3 9 15 13
7 0 13 15 15 13 9 13
7 7 13 9 13 11 0 0
8 7 1 9 3 13 1 15 9
3 13 15 11
4 15 13 13 3
10 0 3 15 3 13 13 1 15 13 15
20 15 13 16 9 13 11 16 13 15 11 13 15 13 1 9 7 0 16 15 13
6 13 3 0 9 13 3
11 3 13 15 9 0 7 9 13 15 1 15
16 16 9 13 15 1 15 3 9 13 15 1 15 7 3 13 15
6 9 3 3 1 15 13
2 13 15
16 7 3 13 9 16 3 15 13 15 3 13 13 3 15 13 3
10 9 13 15 16 13 15 15 3 13 15
6 16 3 15 13 15 15
4 13 15 11 11
2 13 11
9 3 15 13 3 13 3 1 15 13
5 3 3 1 15 13
9 9 1 15 3 13 3 1 15 13
6 3 9 15 1 15 13
3 13 15 11
4 6 6 13 15
9 3 13 9 16 13 15 15 12 9
7 13 1 9 7 1 15 13
7 1 9 9 15 9 0 13
12 16 3 3 3 13 13 15 16 13 13 9 15
20 7 16 13 13 9 15 3 13 7 13 15 1 15 16 3 13 15 3 15 13
8 7 3 15 13 13 7 9 13
5 9 3 13 3 13
5 7 3 9 13 13
3 13 15 11
6 15 13 1 9 3 15
10 16 15 13 13 3 9 15 13 13 3
7 7 3 13 15 7 13 15
3 13 15 11
3 13 15 11
11 0 7 9 1 15 13 7 3 13 3 15
5 11 13 15 13 9
4 7 3 15 13
12 3 13 3 16 15 1 9 7 9 1 15 13
9 9 15 15 13 15 1 15 3 13
8 9 3 13 1 15 0 13 9
10 16 3 3 3 1 0 9 9 13 15
4 6 6 13 15
14 13 1 15 9 15 15 13 3 0 13 7 0 13 0
5 3 15 1 9 13
15 7 15 3 13 1 9 15 0 13 16 13 15 9 1 9
6 16 13 15 9 15 13
29 7 15 13 9 7 15 9 13 15 16 13 1 15 1 9 9 0 15 9 3 13 13 16 3 13 15 7 13 15
4 7 1 15 13
4 3 13 15 0
3 13 1 15
9 3 3 7 9 1 0 3 13 15
11 15 3 13 15 16 15 13 7 15 0 13
17 1 0 9 13 16 15 1 9 15 7 15 1 15 7 15 1 15
16 7 13 15 13 13 9 15 7 15 13 15 7 13 15 15 0
13 9 7 15 13 16 15 13 15 13 7 3 15 9
5 13 11 7 13 15
21 16 15 13 15 9 15 13 7 9 15 13 15 7 1 15 13 7 9 1 15 13
7 3 13 15 9 15 3 13
10 7 9 15 13 13 15 7 13 15 9
6 0 13 15 1 15 13
21 9 3 9 0 15 13 9 1 9 15 0 15 13 15 7 13 15 15 3 13 15
8 3 3 15 9 13 15 13 15
8 3 3 13 15 15 9 7 13
5 13 16 15 13 15
5 13 7 13 1 15
19 16 13 13 15 13 15 13 3 16 13 13 1 9 16 9 15 0 15 13
13 7 3 13 15 3 16 3 13 16 3 13 9 13
6 3 3 3 13 1 15
11 13 3 0 9 9 7 1 15 3 13 15
1 13
2 13 3
9 15 13 9 0 7 9 15 9 13
17 0 9 3 13 9 13 15 7 0 13 9 13 15 16 9 0 13
9 3 15 0 13 1 9 15 13 15
7 13 1 15 7 15 1 15
21 3 9 3 13 9 13 1 15 16 3 13 1 9 3 3 15 16 1 15 3 13
3 15 13 9
22 16 15 1 15 3 13 13 15 3 3 9 7 13 7 13 15 7 1 9 13 7 13
17 16 13 1 15 7 9 15 1 15 13 15 3 13 13 7 13 15
14 1 0 13 15 9 15 16 9 0 13 7 13 15 9
8 3 13 15 9 3 15 13 15
4 13 1 9 15
19 16 9 15 13 13 1 9 15 3 15 9 9 15 13 7 13 1 15 9
14 0 13 15 16 9 15 1 15 13 7 9 15 13 15
14 0 0 9 15 3 13 16 15 9 15 13 1 9 15
5 3 3 13 15 9
8 9 3 3 13 15 13 9 15
13 15 3 13 9 16 15 15 13 1 9 15 13 15
32 3 15 15 13 7 15 13 15 7 13 15 16 15 13 7 9 13 7 9 15 13 16 15 3 13 1 9 1 9 15 13 15
7 0 13 15 16 13 15 15
10 16 9 15 13 13 16 15 1 15 13
16 16 3 1 9 13 7 15 13 15 1 9 0 1 13 15 9
6 13 9 15 15 13 15
6 16 15 13 3 15 13
7 16 9 15 13 3 15 13
13 7 0 15 13 15 1 9 15 16 3 13 13 15
11 16 3 13 13 7 13 15 9 3 13 13
9 3 3 3 9 3 13 1 9 15
15 16 9 3 13 13 1 15 15 15 15 13 9 3 13 13
11 3 3 7 13 7 13 7 15 7 9 15
10 7 16 13 15 9 13 1 9 15 16
20 3 3 13 9 15 15 13 15 1 9 9 0 15 1 9 13 0 13 1 15
9 3 15 3 13 16 3 1 15 13
7 0 13 15 16 3 13 15
4 1 9 13 15
10 7 0 13 15 16 3 13 9 7 15
14 7 0 13 15 16 3 13 9 13 0 16 15 13 15
10 0 3 15 3 3 13 16 1 15 13
13 3 3 13 1 13 15 7 15 1 15 3 13 15
9 7 16 0 13 15 9 0 9 15
5 7 15 9 15 13
6 0 13 15 16 15 13
8 16 3 3 13 13 15 1 15
13 7 13 0 13 9 1 9 7 1 9 7 1 9
8 1 9 3 16 3 13 1 15
13 1 9 3 16 1 9 13 7 1 0 3 13 15
9 1 9 3 16 9 9 0 13 13
11 3 3 13 0 9 0 13 15 1 0 9
16 3 1 15 3 13 13 7 15 3 13 13 13 7 13 13 15
6 15 15 13 9 15 13
11 0 1 13 15 16 1 15 13 7 13 15
20 1 0 7 1 0 3 13 15 7 3 1 0 7 13 15 7 16 13 1 9
7 13 3 1 9 15 1 15
20 15 13 0 15 13 15 1 0 7 3 13 15 7 3 1 0 7 13 15 7
4 16 13 1 9
5 15 13 0 15 13
4 3 13 15 13
10 13 3 11 16 13 15 13 7 13 15
9 1 0 3 13 15 1 15 16 13
13 1 0 7 3 13 15 7 3 1 0 7 13 15
14 6 6 13 15 16 13 15 7 13 15 7 9 13 15
10 15 3 0 13 7 9 15 1 9 13
9 9 3 13 9 13 16 13 9 15
17 3 3 13 15 7 13 15 9 15 7 9 15 15 3 13 1 15
8 7 1 0 9 15 3 13 15
15 6 6 13 15 16 16 15 13 1 9 1 9 15 13 15
7 3 3 13 15 1 9 15
8 13 7 13 16 9 15 13 13
5 0 1 9 13 15
19 7 13 9 3 1 0 1 9 3 13 15 7 3 13 15 1 9 13 15
17 1 0 9 1 9 15 13 7 3 13 15 16 15 13 9 1 15
7 13 1 9 7 13 1 9
7 3 13 9 7 13 1 9
4 13 15 9 15
11 6 3 3 13 15 13 7 9 15 3 13
12 3 13 16 13 15 7 3 13 16 15 15 13
8 1 0 13 16 1 9 13 13
3 13 15 11
3 3 3 13
8 0 13 15 16 1 15 9 13
6 1 9 0 13 7 13
3 15 13 9
12 0 13 11 7 13 11 9 15 1 9 7 13
3 9 13 9
26 13 9 15 16 3 9 15 13 15 3 13 15 13 9 0 9 16 0 15 13 15 13 13 15 9 0
16 6 3 13 0 9 16 13 15 12 0 9 7 15 13 11 11
8 9 13 15 13 13 15 16 13
10 13 9 15 9 15 13 13 15 1 9
11 15 13 7 15 15 13 13 7 9 15 13
11 3 13 16 15 15 13 13 15 1 15 13
25 3 9 15 13 13 15 13 15 7 0 13 7 13 1 9 16 1 15 13 7 13 16 15 15 13
4 15 1 0 13
15 3 1 15 9 13 7 1 0 15 13 13 15 16 15 13
16 7 1 0 13 1 9 7 0 1 9 13 7 15 1 15 13
17 9 0 13 15 1 9 15 15 13 13 15 16 13 12 3 3 15
16 3 1 15 13 7 0 13 1 9 16 13 9 15 13 1 15
20 15 13 15 9 15 7 9 13 15 16 3 13 1 9 3 3 15 1 9 13
13 3 13 16 13 15 1 9 7 16 13 15 1 9
10 1 9 3 13 3 3 15 1 9 13
5 13 15 1 9 15
12 3 15 15 13 1 9 3 15 13 15 1 9
14 7 1 15 15 13 15 0 16 13 3 0 13 1 9
42 3 1 0 3 13 3 7 3 13 9 15 1 15 16 15 12 13 3 15 9 1 15 7 15 1 15 16 3 0 1 15 12 13 16 3 9 9 13 16 15 15 13
29 15 1 15 7 15 1 15 16 13 0 1 12 7 16 13 9 16 15 15 13 7 13 15 13 3 3 15 13 13
30 9 15 13 13 15 13 16 3 13 15 3 0 13 1 15 16 13 9 15 15 13 13 15 16 13 15 13 1 9 9
6 9 0 9 15 3 13
11 15 3 15 13 7 0 13 16 15 15 13
22 0 13 11 13 1 9 15 1 0 9 9 0 3 13 9 1 15 13 0 7 9 15
16 13 3 11 15 15 13 9 16 3 13 15 11 3 1 9 15
18 11 3 13 9 7 1 9 7 9 9 13 3 1 9 7 9 7 9
10 11 3 13 15 13 1 15 13 13 15
2 13 15
2 11 9
3 13 15 11
8 13 3 11 15 15 13 1 15
12 7 16 13 15 15 13 13 3 7 13 1 9
5 3 3 15 13 11
2 15 13
3 0 3 13
2 13 11
5 13 15 16 15 13
7 16 13 15 9 15 13 16
9 15 13 13 15 3 13 15 1 15
11 11 3 11 13 9 13 15 7 13 0 9
5 7 13 15 9 0
5 13 3 9 9 11
4 13 3 11 11
10 9 15 13 15 9 3 13 3 13 15
3 7 13 15
6 7 13 15 1 11 3
4 13 3 9 11
6 15 9 13 1 9 0
5 13 3 7 13 15
11 16 3 13 13 0 9 3 13 13 15 15
4 13 3 15 11
5 3 13 15 13 15
12 16 9 0 13 15 15 13 13 15 9 13 13
12 13 3 3 11 1 9 7 13 11 7 13 15
5 15 3 13 9 0
3 13 15 11
12 1 15 3 15 13 0 7 15 15 13 1 15
2 13 11
4 3 15 9 13
3 15 13 13
2 13 11
6 9 15 13 1 0 9
19 16 1 0 9 13 13 9 15 9 3 15 13 15 13 16 3 13 13 9
6 3 3 9 15 13 3
4 13 3 15 11
5 3 9 3 13 15
2 13 11
8 0 15 13 1 9 13 9 15
3 13 15 11
3 15 13 9
10 7 0 13 3 13 1 9 7 13 15
7 15 3 12 9 13 1 15
10 13 3 9 15 16 12 15 13 1 9
8 13 3 3 16 13 15 9 0
4 3 0 7 11
7 3 3 11 13 11 7 13
18 7 9 13 9 1 9 13 1 9 15 7 1 9 0 13 15 7 13
4 13 15 9 0
5 7 13 15 1 9
5 13 3 3 11 3
3 7 13 15
10 13 3 11 3 13 0 9 7 0 9
3 7 13 15
9 3 3 15 13 9 7 9 13 13
2 13 15
2 13 15
3 13 15 11
4 13 15 7 13
3 13 15 9
15 15 9 13 7 1 9 15 0 13 13 16 9 0 13 15
17 3 3 13 11 0 9 3 13 15 7 13 1 9 3 7 13 11
6 11 3 9 3 13 15
3 13 15 11
4 15 3 3 13
13 3 13 3 16 9 13 13 15 7 9 13 13 15
12 3 13 9 1 15 15 16 3 13 15 13 3
8 0 1 13 15 15 0 9 13
6 1 0 11 13 13 15
4 9 3 13 13
8 0 15 15 13 9 13 15 9
19 11 3 13 0 9 13 3 11 7 13 1 9 1 9 13 11 3 3 11
4 13 3 9 9
3 7 13 9
3 6 9 15
3 0 3 13
1 13
1 13
3 13 15 11
4 9 3 15 13
5 3 13 9 3 9
7 3 3 13 15 16 15 13
5 0 3 13 11 13
30 7 0 15 13 9 13 1 13 0 9 15 13 15 3 11 3 15 13 7 1 15 15 12 3 7 3 1 9 3 11
5 13 3 7 9 11
4 7 13 1 9
4 11 9 9 0
7 7 13 13 3 3 7 3
5 13 3 11 9 0
8 3 13 9 0 7 16 0 13
3 9 13 0
2 13 11
3 15 13 13
17 9 3 3 13 11 13 9 15 7 13 12 9 15 9 9 7 9
3 3 13 15
5 7 13 9 15 13
5 16 13 15 9 13
4 13 15 9 15
6 7 1 9 15 13 9
5 9 3 3 0 13
16 13 3 1 9 0 9 15 7 9 9 15 11 0 7 11 9
12 11 3 13 9 7 9 13 15 13 13 9 15
5 1 0 3 13 9
3 6 9 15
10 7 1 0 9 13 15 9 1 15 15
16 1 0 13 11 16 15 3 13 15 1 15 16 13 15 9 13
1 13
5 9 3 13 0 9
12 0 3 13 9 9 1 9 13 13 1 9 15
6 3 3 13 9 11 13
28 9 3 16 9 13 16 3 13 1 9 9 1 9 13 3 0 9 0 9 13 11 16 13 9 15 7 13 15
12 13 3 9 7 0 13 9 7 0 13 1 15
27 1 11 3 13 16 13 15 3 13 3 13 15 9 7 12 1 9 9 15 9 13 7 13 3 9 7 9
19 7 13 15 13 7 0 13 9 15 7 0 13 16 9 13 16 15 9 13
7 13 3 0 16 13 15 9
5 9 3 13 15 15
5 7 3 0 9 13
22 1 0 3 13 11 11 15 13 1 11 13 9 0 0 3 1 9 0 16 13 9 0
6 13 3 7 13 9 0
18 13 3 3 11 13 1 11 9 3 13 9 0 7 0 3 3 9 12
15 13 3 9 0 7 13 15 9 1 9 3 9 13 9 13
20 13 3 1 9 3 15 13 9 7 1 9 9 0 1 15 3 15 3 13 13
11 3 3 1 9 0 16 1 13 9 13 11
19 1 12 3 9 11 9 13 3 3 13 9 1 9 7 13 9 13 1 9
3 7 13 15
10 13 9 1 9 7 3 13 3 13 15
4 13 3 12 3
11 7 0 9 13 3 11 7 13 3 1 9
5 7 13 13 9 13
3 3 3 13
34 13 3 3 11 11 1 9 15 7 13 3 1 9 7 13 9 13 7 9 15 13 1 9 15 3 1 9 13 7 3 13 1 12 9
11 3 3 3 13 9 16 13 15 1 0 13
6 13 3 3 1 15 9
8 11 3 13 1 9 3 13 15
19 7 13 12 9 1 0 13 12 1 9 7 12 1 9 3 13 13 9 0
4 7 13 15 0
4 9 15 13 15
3 13 15 16
15 0 13 13 15 3 7 13 11 13 7 3 13 16 11 13
3 13 15 11
4 9 15 15 13
2 15 13
15 9 16 15 13 13 13 15 3 15 13 13 7 15 15 13
4 13 15 11 11
7 13 3 15 0 13 15 3
4 15 13 15 9
3 13 15 11
4 3 13 15 15
7 3 3 3 13 1 9 15
8 13 3 1 9 15 7 13 15
12 13 11 9 13 9 16 13 9 7 0 13 15
22 13 3 3 1 0 9 1 12 9 7 9 13 3 13 9 15 13 1 9 0 13 11
2 9 15
11 7 0 13 13 15 9 7 9 7 9 15
6 13 3 15 9 13 9
4 13 15 11 3
2 9 15
8 3 13 15 9 3 15 13 15
3 13 9 0
17 11 3 12 1 12 1 12 13 9 3 13 3 1 15 3 13 11
5 13 3 15 0 9
2 13 9
4 0 3 13 15
25 16 3 13 1 9 15 9 0 7 13 9 15 1 9 15 7 13 9 15 1 9 0 3 13 9
13 7 1 12 9 3 13 3 9 15 7 11 1 15
10 13 11 9 13 7 13 1 9 7 13
23 13 9 15 3 7 13 9 15 7 13 9 15 7 13 1 9 15 7 3 13 0 7 0
6 7 13 11 7 13 15
2 9 15
2 9 15
4 13 15 11 16
3 13 15 13
5 0 3 13 7 13
16 0 3 15 9 13 11 1 9 15 15 3 13 13 1 9 0
11 1 0 13 15 3 11 9 15 1 9 0
4 13 3 15 3
24 13 3 11 11 7 11 13 11 7 11 15 13 1 11 0 7 9 0 7 15 12 1 9 15
4 13 15 11 11
3 13 9 13
2 13 15
5 13 3 15 1 15
14 7 13 7 13 1 9 3 7 1 0 9 3 13 15
4 13 3 15 11
5 9 3 15 0 13
3 13 3 15
1 3
4 0 3 13 15
8 13 1 0 9 9 9 7 13
12 13 3 7 1 0 3 13 13 15 1 9 9
2 9 13
5 7 0 9 9 13
14 3 13 3 3 1 9 7 3 12 12 9 13 9 9
15 16 3 13 1 9 13 9 13 7 9 1 15 13 7 9
3 13 15 11
6 13 1 9 15 13 3
18 13 3 11 11 7 13 9 1 9 0 0 9 12 7 12 12 7 12
3 13 15 11
1 13
15 7 15 3 13 1 9 13 15 15 15 13 13 16 9 13
12 13 3 11 7 13 9 7 13 15 7 9 3
11 6 3 3 13 15 11 9 15 13 1 0
7 3 3 13 13 11 11 11
7 11 0 13 3 15 3 0
7 6 9 15 13 16 13 15
2 13 15
3 13 9 15
5 11 0 13 3 15
4 13 15 6 9
5 15 13 16 13 15
2 13 15
3 13 15 3
