6471 11
24 2 10 9 4 3 13 2 13 15 4 9 9 1 15 2 16 4 13 2 16 15 9 13 2
8 9 1 11 4 13 0 9 2
17 9 4 1 0 9 13 13 2 16 4 15 13 2 4 13 9 2
8 13 4 1 9 7 13 4 2
6 15 15 14 4 13 2
24 15 15 4 13 2 4 13 14 0 9 1 9 2 2 4 1 9 1 11 1 11 13 9 2
15 9 1 0 9 4 13 2 16 4 15 9 13 3 3 2
20 9 1 0 9 7 4 13 2 3 4 9 1 11 3 13 13 0 0 9 2
21 1 9 4 13 14 1 9 1 9 2 16 13 0 9 7 9 9 7 10 9 2
20 1 9 4 14 1 9 13 15 0 1 9 9 2 1 15 4 13 9 0 2
26 9 9 9 13 0 1 9 9 1 0 9 1 0 9 2 1 9 7 4 15 14 15 13 0 9 2
18 7 4 3 13 9 2 1 15 4 13 2 3 4 13 1 0 9 2
10 15 13 9 2 13 9 3 3 0 2
29 3 13 9 9 9 2 16 13 0 1 9 2 16 13 1 9 2 3 13 9 9 9 2 9 2 9 2 9 2
12 3 13 3 13 9 2 1 15 4 15 13 2
8 3 13 9 14 9 0 9 2
13 2 13 0 9 9 2 15 13 9 7 3 13 2
18 0 9 1 9 2 16 4 15 13 10 9 2 13 14 9 1 15 2
24 1 10 9 4 11 11 13 2 16 13 2 9 0 9 1 9 9 2 7 13 3 0 2 2
13 0 9 13 1 9 3 0 0 9 7 0 9 2
10 1 10 9 7 13 3 0 0 9 2
18 13 4 14 1 0 9 1 10 0 9 2 16 13 1 9 10 9 2
24 11 11 2 9 2 9 0 9 7 9 2 7 4 9 13 9 1 9 2 9 7 0 9 2
27 1 0 9 1 0 0 9 13 9 1 0 9 7 10 9 1 0 9 13 1 9 2 16 3 13 9 2
25 3 0 9 9 1 0 9 13 1 9 2 16 13 3 0 1 0 9 3 2 16 1 15 13 2
13 9 13 2 9 2 7 13 1 9 1 0 9 2
54 9 11 13 3 10 9 9 2 0 1 0 9 2 16 13 9 7 9 0 9 1 9 2 7 1 9 13 3 1 9 2 16 13 1 9 2 7 1 10 9 0 2 3 4 3 13 9 7 13 0 9 1 9 2
23 9 9 13 9 9 2 0 9 2 16 13 7 13 10 9 2 7 4 13 13 3 0 2
15 3 3 14 4 10 9 13 9 2 9 7 9 10 9 2
22 13 13 3 9 2 16 15 13 7 13 10 0 9 2 16 13 9 2 9 7 9 2
16 1 9 13 3 2 16 13 2 3 10 9 13 1 0 9 2
11 13 15 1 10 9 7 13 10 0 9 2
17 13 10 9 2 16 15 13 3 7 16 4 1 15 3 13 9 2
19 0 9 13 0 9 7 0 9 7 3 0 9 2 16 15 13 1 9 2
10 1 10 9 15 3 0 9 14 13 2
11 9 1 0 0 9 13 0 0 0 9 2
17 1 9 0 13 0 7 3 0 9 2 16 13 9 3 0 9 2
17 0 0 9 11 12 1 9 11 4 14 3 13 1 10 0 9 2
11 1 9 4 13 3 9 0 13 10 9 2
14 0 9 0 0 9 4 13 1 9 9 9 11 11 12
23 9 9 15 4 13 14 1 9 0 0 9 2 16 4 13 9 9 11 7 11 11 11 2
9 3 4 13 9 7 9 10 9 2
20 0 9 4 13 9 1 9 11 2 16 4 14 1 9 13 9 10 0 9 2
22 9 0 9 13 7 1 11 14 3 3 7 1 0 9 9 11 11 15 4 13 13 2
16 9 4 13 1 9 1 9 2 9 7 4 13 1 12 9 2
20 9 9 9 11 13 1 9 9 2 9 2 9 9 2 9 2 9 2 9 2
25 0 9 4 9 3 13 2 16 4 15 13 2 16 11 8 2 16 13 9 2 13 7 13 9 2
10 1 10 9 14 4 4 13 14 9 2
14 3 4 15 13 7 13 11 8 13 2 4 13 9 2
2 11 11
21 0 9 4 9 9 13 1 0 9 2 16 13 1 10 9 1 2 0 9 2 2
11 0 0 9 13 1 15 0 1 0 9 2
10 1 0 9 15 0 9 13 16 9 2
5 3 15 15 13 2
20 13 4 1 9 2 16 4 15 3 13 14 3 7 15 1 9 3 13 15 2
29 13 4 3 2 16 4 13 15 14 0 9 1 9 2 7 10 9 4 15 13 10 0 9 7 15 4 14 13 2
18 13 4 10 0 0 9 2 16 4 3 13 2 3 3 15 15 13 2
18 1 9 14 4 13 3 9 9 2 12 9 9 2 3 16 1 12 9
29 1 0 9 1 11 1 11 4 1 9 2 12 2 7 9 2 12 9 2 13 12 0 9 9 2 9 7 9 2
21 13 15 4 12 9 1 12 9 2 16 4 13 7 13 0 7 0 9 0 9 2
19 9 4 1 9 2 12 9 2 1 12 9 13 11 11 2 9 0 9 2
19 3 4 13 3 0 0 0 9 11 1 11 2 16 4 13 11 11 11 2
26 16 4 14 13 2 4 13 9 11 12 1 9 2 16 4 1 9 13 0 9 11 11 2 11 2 2
16 1 9 9 11 11 4 1 9 1 9 0 9 13 11 11 2
3 2 8 2
20 13 1 9 2 16 13 9 1 9 1 10 9 2 3 7 13 0 1 9 2
21 15 0 13 14 9 9 2 0 13 1 9 7 15 1 9 3 13 1 0 9 2
22 9 15 13 0 14 1 0 9 2 9 7 9 2 13 7 15 1 12 9 9 3 2
9 1 9 15 14 13 13 9 9 2
6 14 9 9 13 0 2
31 1 3 0 9 4 13 2 16 14 4 9 13 0 1 9 2 15 13 2 16 4 11 1 10 0 9 9 13 9 9 2
26 1 15 14 4 13 9 1 9 9 1 0 9 2 3 7 4 3 1 9 13 0 9 1 10 9 2
22 14 1 11 13 9 7 9 1 3 0 9 9 2 7 4 13 13 10 9 9 9 2
27 16 9 1 9 9 13 14 1 10 9 7 0 9 2 13 3 14 1 0 3 13 1 9 7 9 9 2
24 13 4 2 16 4 13 15 2 16 4 1 12 9 13 0 9 2 3 0 9 1 0 9 2
35 1 0 9 4 13 9 1 0 9 7 15 13 13 2 16 13 1 15 0 7 16 13 7 13 10 9 2 10 9 1 0 7 0 9 2
13 3 15 15 10 9 13 2 4 13 0 0 9 2
43 1 9 11 1 11 4 9 13 2 16 15 15 13 2 7 15 1 0 9 1 11 13 13 2 16 4 0 9 11 13 14 9 2 16 4 15 14 1 10 9 13 9 2
26 4 7 13 14 1 9 2 16 15 13 10 9 13 2 3 4 13 14 1 11 2 11 7 11 2 2
30 0 9 13 9 0 9 2 15 13 2 16 13 1 0 9 11 0 9 10 9 13 14 12 7 12 9 0 0 9 2
20 1 0 9 1 11 4 7 1 11 13 0 0 9 7 0 9 4 13 9 2
6 3 4 13 1 9 2
14 3 4 14 13 1 9 2 14 2 15 4 14 13 2
15 3 13 2 10 9 3 13 10 9 7 15 3 13 2 2
6 14 2 7 3 13 2
2 9 2
2 9 2
6 4 13 1 0 9 2
8 13 10 9 0 1 10 9 2
11 14 2 13 2 16 4 15 0 9 13 2
6 3 4 15 3 13 2
4 13 10 9 2
34 16 4 13 9 2 4 13 2 3 15 4 0 9 2 0 1 0 9 2 13 9 7 9 15 4 15 13 2 3 4 15 15 13 2
6 13 4 9 1 15 2
5 13 4 16 0 2
19 3 4 13 12 2 12 9 2 9 15 4 3 13 2 16 4 13 9 2
9 1 10 0 9 4 13 3 0 2
18 15 4 3 13 10 12 9 2 3 2 16 4 9 13 9 9 0 2
12 13 4 1 9 7 13 2 16 15 4 13 2
15 13 2 3 10 0 9 13 1 10 9 1 15 2 2 2
11 3 13 9 2 16 14 14 13 1 15 2
8 7 14 13 2 4 3 13 2
16 16 7 4 13 2 4 9 11 2 16 4 13 2 13 13 2
16 9 4 13 3 2 16 4 10 9 13 1 0 9 1 11 2
7 10 9 4 14 13 9 2
4 13 4 0 2
10 3 4 13 1 10 9 14 0 9 2
10 10 0 9 9 13 0 1 10 9 2
3 0 9 2
2 0 2
4 9 0 9 2
3 13 15 2
6 0 9 13 1 9 2
12 13 9 2 3 4 13 1 9 10 9 2 2
3 13 15 2
3 13 9 2
10 9 15 13 9 7 9 13 13 9 2
4 3 13 13 2
8 1 9 13 2 3 15 13 2
7 15 13 12 10 0 9 2
9 13 4 0 15 12 2 12 9 2
33 14 16 4 13 2 4 13 1 12 1 9 2 1 9 13 1 0 0 9 9 2 16 4 3 13 2 16 4 13 1 0 9 2
18 13 4 2 16 4 9 13 7 13 2 16 13 1 10 9 3 0 2
8 13 4 7 15 3 13 3 2
9 1 10 9 4 13 15 13 9 2
8 15 7 15 14 4 13 15 2
9 13 15 15 2 16 4 13 15 2
5 13 4 0 15 2
7 13 4 1 9 15 0 2
16 1 9 4 13 9 7 15 13 2 16 16 13 15 3 0 2
10 3 15 4 13 1 9 7 13 15 2
2 9 2
5 15 15 7 13 2
4 9 13 0 2
36 16 4 13 0 9 2 4 3 2 16 16 15 13 1 9 1 9 2 13 1 10 9 2 14 3 13 1 9 7 15 14 3 13 1 9 2
33 3 4 9 3 13 7 15 13 1 9 9 1 15 2 16 15 4 3 13 2 3 15 4 13 1 9 2 16 4 15 13 0 2
28 16 4 9 13 1 9 9 2 4 15 13 2 16 13 15 3 0 2 16 15 13 3 2 16 13 1 9 2
34 16 4 9 13 2 16 15 1 0 9 14 13 2 15 4 14 15 3 13 7 15 3 13 3 1 0 7 1 10 9 0 0 9 2
7 14 10 0 9 4 13 2
24 14 13 4 2 16 13 9 2 16 3 13 1 9 7 15 13 2 16 14 4 13 3 0 2
7 3 13 9 13 2 2 2
1 2
8 9 4 3 13 13 1 3 2
28 0 9 11 11 1 9 0 9 11 11 15 4 3 7 13 2 16 15 4 13 9 1 9 8 9 8 11 2
11 11 4 13 9 1 9 7 13 0 9 2
28 10 0 9 11 11 4 13 0 1 9 0 9 1 0 9 2 13 7 4 1 12 0 7 3 0 0 9 2
36 9 4 1 0 9 11 7 10 9 13 14 1 9 2 16 15 4 1 12 0 9 1 0 9 1 11 13 9 0 9 0 9 11 1 11 2
8 14 13 2 3 14 13 3 2
7 15 14 13 2 15 13 2
51 3 13 14 3 0 2 16 1 9 9 1 9 14 13 14 11 2 16 13 15 1 9 2 15 4 13 11 2 16 3 13 1 11 2 7 9 9 11 2 3 16 15 1 11 13 11 7 3 14 11 2
18 14 7 3 13 2 3 13 8 8 2 16 3 14 2 13 9 2 2
25 1 11 4 13 2 16 3 13 10 16 12 9 0 0 9 2 15 13 3 1 3 3 16 3 2
8 0 9 0 9 7 14 13 2
20 3 4 13 7 3 14 3 13 2 7 13 14 10 0 9 0 1 0 9 2
10 9 13 12 2 15 13 0 1 9 2
8 0 1 9 13 9 7 9 2
6 0 9 11 11 12 2
15 1 12 13 9 2 16 15 0 9 0 9 14 14 13 2
14 11 12 13 1 9 9 2 16 13 0 14 10 9 2
11 15 13 1 9 12 9 0 14 0 9 2
23 10 9 4 3 13 3 2 16 4 13 2 3 14 13 2 16 13 12 0 14 1 15 2
12 3 13 12 15 0 2 9 9 13 14 0 2
21 0 14 13 2 7 13 1 10 0 9 0 9 1 9 9 1 0 9 2 9 2
11 2 11 9 2 7 13 1 9 1 9 2
21 13 9 9 7 0 9 7 13 15 9 1 11 2 1 11 2 0 11 2 11 2
14 3 13 1 15 11 12 2 7 3 14 13 1 9 2
22 0 13 14 15 2 16 4 11 1 9 13 9 2 16 15 1 10 0 9 4 13 2
15 11 4 14 13 2 16 9 10 9 11 13 14 10 9 2
23 14 2 16 4 13 10 9 9 11 0 1 9 14 0 9 2 4 13 10 9 3 0 2
31 0 9 2 16 13 1 9 0 9 0 9 9 2 13 3 3 0 1 9 2 16 4 9 13 0 9 1 11 2 11 2
34 9 13 0 2 7 4 13 1 9 0 0 9 1 9 9 2 16 15 13 1 10 9 1 9 9 9 7 14 14 0 9 0 9 2
18 9 4 3 13 1 9 0 9 7 1 9 14 3 13 9 10 9 2
7 3 15 13 1 0 9 2
18 14 14 16 9 2 9 9 13 1 10 0 9 10 16 12 0 9 2
4 11 13 0 2
32 14 13 15 2 3 4 13 10 16 10 9 1 9 9 9 2 16 15 4 13 10 0 9 2 15 15 7 14 3 4 13 2
36 14 7 1 0 9 7 9 7 9 13 9 7 9 0 9 4 13 3 2 16 15 4 3 1 9 13 1 0 9 1 9 2 9 7 9 2
25 10 9 4 13 2 16 10 9 10 9 14 13 1 9 2 3 7 15 4 13 1 9 7 9 2
11 3 13 9 10 9 1 3 0 0 9 2
32 11 11 4 13 1 0 2 7 0 9 2 16 4 13 1 9 10 9 3 3 2 16 7 15 15 4 3 13 1 9 13 2
23 0 9 4 13 13 0 7 9 7 0 9 15 3 3 13 9 1 9 2 9 2 2 2
30 9 0 9 9 13 12 9 9 2 0 7 13 12 9 9 9 0 0 9 2 4 13 1 9 9 1 9 0 9 2
35 2 7 4 14 9 3 1 0 9 11 13 9 10 0 0 9 2 16 4 1 15 1 10 9 13 0 0 9 3 12 9 9 1 9 2
17 2 7 4 9 0 9 9 11 13 2 16 13 9 0 9 11 2
41 1 0 9 7 9 4 0 0 9 13 9 1 9 1 9 11 2 0 0 0 9 7 0 9 11 11 2 16 4 13 9 10 0 9 7 1 9 14 0 9 2
22 1 0 9 4 13 2 15 4 13 2 7 15 15 4 3 13 1 9 10 0 9 2
10 15 13 14 3 3 2 13 9 9 2
13 3 7 1 3 13 0 0 9 1 9 7 11 2
9 1 10 9 13 3 14 15 13 2
24 1 9 0 0 9 4 1 11 13 14 9 9 7 3 9 12 15 4 9 13 1 0 9 2
36 11 4 13 1 9 14 9 0 9 11 11 11 2 16 10 9 13 2 16 4 13 9 9 3 0 2 16 7 15 4 13 1 0 9 9 2
22 11 7 4 14 13 2 16 13 0 9 0 1 0 9 9 0 9 7 10 0 9 2
20 0 11 11 4 1 11 13 12 9 16 9 1 0 9 1 9 7 0 9 2
21 1 0 9 9 4 13 13 12 9 2 4 13 13 0 7 13 4 13 0 9 2
14 1 9 4 15 13 12 9 2 9 4 13 1 9 2
10 14 3 4 13 9 0 1 9 9 2
23 14 1 9 3 1 9 13 10 9 16 1 9 2 14 7 13 3 14 10 9 16 9 2
43 14 0 9 13 1 0 9 0 9 0 9 2 10 12 9 13 3 10 9 2 16 15 15 14 3 13 3 2 3 15 13 2 15 4 13 1 0 7 0 9 0 9 2
14 7 13 10 9 2 9 7 9 9 1 9 1 9 2
19 14 10 9 2 9 4 1 9 1 9 2 16 4 13 9 2 13 0 2
35 0 13 14 9 9 0 9 2 16 15 13 1 0 9 9 2 1 9 2 16 13 0 2 15 13 1 9 7 3 13 1 9 0 9 2
27 9 9 2 9 2 9 9 2 9 9 7 9 13 9 9 7 9 2 16 13 0 1 0 9 0 9 2
6 3 13 14 12 9 2
14 0 9 1 11 2 1 9 2 12 9 2 3 13 2
19 11 15 4 1 0 9 3 13 2 15 13 15 2 16 15 13 1 9 2
6 3 15 4 15 13 2
10 0 9 7 9 1 9 0 9 1 11
12 0 9 4 13 0 9 11 11 1 0 9 2
28 1 15 13 0 2 3 4 13 3 13 1 9 0 0 9 2 7 1 15 13 0 9 0 9 0 1 9 2
18 7 13 3 1 9 0 9 11 13 0 0 9 1 0 9 0 9 2
13 1 11 1 15 13 0 10 9 1 2 9 2 2
9 11 3 13 9 9 0 9 11 2
9 11 14 13 9 0 9 1 11 2
17 1 9 7 14 1 9 4 3 3 13 14 2 16 13 3 0 2
18 3 0 13 1 11 9 0 9 2 3 3 15 4 11 13 1 9 2
11 0 9 15 13 13 2 16 4 13 9 2
7 1 9 13 11 7 9 2
25 11 2 1 9 4 1 0 9 9 9 2 0 9 0 9 2 14 3 13 12 2 0 11 11 2
48 0 9 11 11 2 16 4 1 9 1 9 9 10 9 13 2 3 14 13 0 0 9 0 9 7 7 14 15 3 13 0 9 1 0 9 2 4 9 11 11 1 9 13 9 9 1 9 2
38 9 10 0 9 7 0 9 13 1 10 9 2 16 3 14 14 13 0 0 9 10 9 2 14 3 7 15 3 1 9 4 13 13 0 9 10 9 2
15 7 13 9 0 9 1 9 0 9 0 9 9 0 9 2
35 7 16 13 2 16 9 3 13 14 1 0 9 2 13 3 14 0 9 10 9 2 16 15 0 9 14 13 0 9 7 14 13 10 9 2
14 0 9 7 9 0 0 9 15 13 1 9 1 9 9
16 11 1 11 2 0 9 2 9 0 9 2 13 12 2 9 2
17 11 2 9 0 9 4 13 3 0 9 0 0 9 1 10 9 2
27 11 4 2 3 16 1 11 2 11 7 11 4 13 0 9 1 9 2 1 9 1 11 13 3 1 9 2
16 13 15 2 16 4 15 9 0 9 0 9 3 14 3 13 2
22 1 12 9 4 15 3 13 1 0 0 9 2 3 15 4 11 3 13 1 0 9 2
15 11 15 4 14 3 14 1 3 10 9 13 1 0 9 2
25 3 16 4 0 9 1 11 3 13 2 4 13 16 0 3 3 0 7 1 15 0 9 3 13 2
33 11 11 2 0 9 1 9 2 4 1 9 13 2 16 4 15 13 1 10 9 2 7 9 11 11 1 0 9 14 13 3 0 2
14 2 9 13 2 16 15 1 12 9 12 3 13 9 2
17 0 9 1 9 0 9 1 9 12 4 1 9 0 9 14 13 2
28 9 1 11 2 12 0 9 1 11 2 4 15 3 3 13 1 9 9 9 7 1 10 9 13 0 9 9 2
20 9 7 14 4 13 14 13 9 1 9 2 16 15 4 15 7 10 9 13 2
25 16 4 1 9 13 1 9 7 15 13 1 0 9 7 1 9 2 4 13 13 0 9 0 9 2
20 12 1 9 2 16 15 4 13 14 13 2 13 0 9 2 16 13 9 0 2
48 1 12 2 9 9 13 0 0 9 0 9 1 9 9 7 9 9 1 9 0 9 9 9 12 1 0 9 9 2 16 4 9 9 13 1 9 1 9 0 0 9 1 9 11 1 9 11 2
30 9 4 3 13 9 0 11 1 9 11 2 9 0 2 0 7 0 9 0 9 2 7 0 11 2 16 13 0 11 2
28 3 4 15 10 9 13 1 0 9 7 9 1 0 9 2 1 15 4 9 3 13 14 1 0 7 0 9 2
16 9 4 13 0 0 7 0 9 1 0 9 1 0 9 9 2
48 3 15 4 13 1 0 9 0 0 9 1 0 9 12 2 16 13 14 3 9 9 2 1 9 0 9 7 0 9 2 7 4 1 9 12 2 12 13 14 0 9 0 9 1 0 9 12 2
21 14 1 9 9 13 9 1 10 9 0 9 0 9 1 11 7 0 9 1 11 2
36 9 12 4 13 9 1 9 9 1 0 1 0 0 9 2 16 14 4 13 1 9 0 0 9 2 10 9 7 4 13 9 9 9 9 12 2
32 3 13 9 1 10 0 9 14 1 9 12 0 9 1 9 8 11 1 11 7 9 12 0 9 1 0 9 1 9 1 11 2
36 1 0 9 4 13 14 0 9 1 9 11 11 7 0 9 1 9 9 11 1 11 2 0 9 1 11 7 0 7 0 9 1 11 1 11 2
49 1 9 9 11 11 7 10 9 13 0 9 1 12 2 0 9 9 9 2 9 0 9 1 9 9 11 2 9 2 16 4 13 1 9 7 1 9 2 9 9 1 0 9 7 13 0 1 9 2
2 8 8
5 3 15 15 13 2
18 3 3 13 9 1 9 2 16 15 15 13 1 0 2 3 0 9 2
14 13 2 16 13 1 9 2 3 2 10 16 12 9 2
10 14 3 0 9 1 9 15 13 9 2
13 0 9 1 0 9 9 15 13 1 0 0 9 2
4 13 1 9 2
14 1 9 13 14 0 9 2 16 15 15 3 13 9 2
16 15 13 0 9 1 9 2 16 15 13 0 7 3 0 9 2
8 10 0 9 13 14 10 9 2
14 3 7 15 15 4 0 9 9 1 10 9 3 13 2
13 9 15 13 1 9 2 16 13 3 0 9 9 2
7 13 15 1 0 0 9 2
9 15 13 1 0 0 9 1 9 2
9 9 4 13 0 9 1 0 9 2
8 15 13 9 2 0 0 9 2
24 3 14 13 2 16 4 13 3 0 9 2 16 15 4 11 1 12 9 9 3 13 1 9 2
14 9 13 9 9 2 0 0 9 13 3 1 11 11 2
13 1 0 9 0 9 13 0 9 8 11 3 3 2
11 3 13 2 16 13 10 0 9 9 11 2
15 9 14 13 3 15 9 2 7 15 1 0 9 13 3 2
20 3 15 0 9 9 1 9 1 10 9 13 2 16 15 15 3 13 14 3 2
13 1 3 13 14 10 9 2 9 7 0 0 9 2
18 0 9 13 9 2 16 13 1 0 9 7 1 9 13 0 0 9 2
7 9 4 13 9 1 9 2
8 3 15 15 13 9 7 9 2
4 13 15 3 2
17 1 9 3 3 15 13 10 9 2 16 15 13 13 1 0 9 2
27 0 0 9 10 0 9 15 4 14 1 0 9 13 2 1 0 7 13 3 15 3 1 0 1 0 9 2
12 9 2 16 4 13 9 9 2 13 13 3 2
22 1 9 13 13 10 3 3 0 9 2 16 15 13 1 10 9 13 1 9 7 9 2
16 3 14 13 3 1 9 0 9 2 16 15 13 3 1 9 2
6 0 9 15 14 13 2
24 13 0 2 7 9 13 2 16 4 10 9 9 13 1 9 2 16 15 4 10 9 13 3 2
8 14 7 2 3 15 3 13 2
18 13 0 9 7 1 15 13 9 2 3 16 4 3 13 0 9 9 2
12 15 13 9 9 7 9 2 3 15 13 3 2
9 0 3 0 9 13 14 1 9 2
20 11 4 13 3 2 11 7 3 15 2 13 2 0 10 9 2 16 3 13 2
17 15 4 15 13 2 16 4 14 1 10 9 2 13 1 9 2 2
8 1 9 1 15 13 15 14 2
14 3 15 4 13 9 7 13 4 15 9 1 0 9 2
16 9 4 13 3 7 1 9 4 13 10 9 14 1 0 9 2
8 1 9 4 13 0 9 3 2
8 15 7 4 13 9 1 12 2
28 16 4 13 13 2 4 13 1 15 12 9 9 2 3 7 15 4 13 14 1 10 9 0 9 9 7 9 2
33 16 4 15 3 3 3 13 2 13 0 9 10 12 9 3 1 9 1 0 9 7 1 0 9 13 9 2 16 13 9 1 0 2
13 11 15 13 1 15 2 16 4 15 13 1 9 2
11 14 9 14 13 13 7 14 13 1 15 2
15 3 15 13 2 9 2 2 16 4 13 1 9 10 9 2
9 1 15 15 13 9 1 0 9 2
16 16 3 13 0 9 2 3 3 13 2 16 13 3 14 0 2
11 3 13 2 16 4 15 3 14 13 9 2
15 3 4 13 0 9 2 16 4 13 3 13 1 10 9 2
7 7 15 15 15 14 13 2
12 1 15 15 13 13 9 2 3 13 1 9 2
13 1 0 9 4 15 13 1 9 1 9 16 0 2
9 0 9 9 15 4 13 1 9 2
6 3 4 9 13 0 2
22 3 13 1 0 9 1 9 1 0 2 16 0 9 1 9 13 9 7 13 0 9 2
9 3 14 3 3 15 13 1 9 2
18 1 15 7 13 14 3 0 9 1 9 14 10 12 9 1 9 9 2
22 9 13 3 1 0 7 1 9 0 9 2 16 15 1 0 3 13 1 0 9 9 2
41 16 13 9 14 0 2 9 14 13 0 16 15 2 16 4 14 3 3 13 1 9 7 13 2 3 4 15 13 1 0 9 2 16 4 15 9 1 0 9 13 2
20 9 11 4 1 0 0 9 13 2 2 6 2 0 1 15 15 4 13 13 2
4 13 4 13 2
16 3 15 4 13 9 1 9 2 1 15 4 13 9 1 9 2
10 0 4 13 1 0 9 7 0 9 2
7 1 9 4 13 0 9 2
15 9 4 13 14 3 0 2 0 1 9 7 9 1 9 2
25 4 15 13 13 2 16 4 13 1 9 7 13 1 9 2 16 4 13 9 2 7 15 4 13 2
27 13 4 9 2 16 15 14 4 0 13 3 2 7 15 13 2 16 15 4 9 13 7 13 0 0 9 2
9 2 15 14 13 2 2 4 13 2
5 15 13 0 9 2
3 1 9 2
7 15 13 3 10 0 9 2
13 2 1 9 1 11 11 4 15 13 13 1 9 2
14 9 4 13 2 16 4 15 13 9 2 16 13 9 2
19 1 9 4 15 7 13 9 2 3 16 4 13 2 16 4 13 10 9 2
10 13 4 1 9 7 15 13 0 9 2
7 2 16 4 15 3 13 2
11 7 13 4 2 16 15 10 9 4 13 2
11 4 13 2 16 4 15 13 1 10 9 2
16 7 16 4 13 10 9 2 4 13 2 16 13 14 1 9 2
7 16 14 4 13 1 9 2
11 16 4 13 3 0 7 16 4 13 9 2
5 11 4 3 13 2
4 7 13 0 2
15 13 4 0 9 2 16 15 0 9 14 4 13 1 9 2
10 2 1 0 9 13 2 2 4 13 2
7 3 7 3 15 13 13 2
5 9 4 13 0 2
10 1 9 9 4 13 1 9 0 9 2
19 9 4 1 9 13 10 0 9 2 1 9 1 15 4 3 13 0 9 2
9 15 15 15 4 13 1 0 9 2
32 11 4 13 1 9 9 7 13 1 0 9 9 2 16 15 4 13 2 11 15 4 13 1 11 11 7 11 15 4 13 9 2
19 4 15 13 2 3 15 4 3 13 3 3 2 3 0 9 7 3 3 2
3 13 4 2
4 3 4 13 2
21 1 0 9 4 11 13 2 2 16 13 15 0 2 14 13 1 15 7 14 13 2
16 3 13 11 11 1 10 9 7 9 15 9 2 9 7 9 2
22 14 15 13 1 0 9 7 13 1 0 9 2 16 4 13 10 9 7 3 13 9 2
10 0 9 15 13 1 9 10 0 9 2
17 13 15 1 10 9 7 15 1 0 0 9 3 13 1 0 9 2
2 9 2
14 9 4 9 13 0 9 7 13 9 1 9 0 9 2
25 7 0 9 14 3 13 2 1 0 9 7 4 13 9 2 3 4 7 13 9 7 0 9 13 2
26 1 10 9 13 14 0 9 2 16 13 0 1 0 7 1 15 14 4 13 0 0 9 13 14 3 2
39 14 7 15 15 13 2 16 4 9 7 9 1 9 1 10 9 13 2 16 15 9 0 2 0 9 14 13 7 16 15 13 1 9 15 14 14 15 13 2
23 1 12 1 9 15 4 9 1 9 8 11 11 13 2 16 3 0 13 9 1 0 9 2
27 1 16 4 9 13 14 0 9 7 13 9 2 3 4 3 13 9 7 9 2 4 9 14 1 9 13 2
35 9 11 4 0 9 13 1 12 9 2 1 12 9 9 2 9 9 7 4 1 0 9 13 3 12 9 9 2 15 13 0 9 1 9 2
10 2 1 0 9 15 9 14 13 15 2
27 9 11 4 13 1 0 11 2 16 4 13 0 7 0 9 2 3 7 13 10 9 1 0 7 0 9 2
34 9 4 13 1 9 0 9 1 9 12 9 1 9 9 2 7 4 9 7 15 0 9 13 7 15 1 9 0 11 13 1 0 9 2
36 1 15 9 9 2 3 2 14 13 3 0 2 16 4 1 15 1 9 14 13 1 15 2 16 4 9 9 0 7 0 9 13 1 10 9 2
21 16 13 9 1 9 0 9 10 9 2 7 1 9 9 1 0 9 15 13 3 2
23 0 9 2 9 9 2 4 13 7 3 0 1 9 2 9 7 1 15 0 9 10 9 2
25 1 9 9 0 9 11 11 11 13 11 1 12 9 14 1 0 9 2 16 13 0 9 0 9 2
34 9 9 11 7 9 0 0 9 11 11 7 4 13 2 16 0 9 3 14 13 1 9 1 0 9 2 16 15 1 3 14 13 0 2
37 2 0 9 0 0 9 1 0 7 3 0 9 4 13 9 9 2 16 15 4 13 0 0 9 2 2 4 13 9 9 0 9 1 11 11 11 2
20 1 10 9 4 8 11 13 1 9 2 16 9 7 9 13 14 0 0 9 2
26 3 0 13 9 10 9 2 16 15 13 9 2 15 4 13 0 9 1 9 2 10 0 9 4 13 2
7 3 15 4 9 14 13 2
14 3 7 4 14 13 13 9 2 7 15 13 1 9 2
21 2 16 13 10 9 9 2 13 3 0 2 9 9 7 9 1 0 7 13 0 2
33 9 11 4 13 2 16 0 9 1 9 9 13 14 0 0 9 2 7 4 13 13 10 9 3 7 13 0 9 1 9 0 9 2
16 1 0 0 9 3 4 7 3 13 1 9 2 2 13 11 2
9 9 13 0 14 1 9 1 9 2
10 9 13 0 2 9 13 1 0 9 2
6 9 3 13 1 9 2
9 9 13 0 9 1 0 0 9 2
6 9 13 9 0 9 2
10 3 13 0 2 0 2 0 7 0 2
8 0 13 0 2 7 3 0 2
6 1 9 15 3 13 2
11 3 15 3 13 0 7 0 9 0 9 2
21 1 9 15 13 9 2 7 13 13 10 9 0 7 3 0 2 16 13 0 9 2
9 9 9 13 0 1 0 9 9 2
9 1 0 9 13 9 7 0 9 2
18 9 1 9 9 11 13 3 0 9 2 0 1 9 0 7 0 9 2
13 16 4 9 13 2 13 13 10 9 9 7 9 2
13 3 13 9 7 9 2 13 0 9 7 9 9 2
7 9 13 1 9 1 9 2
23 3 2 16 4 13 9 2 3 1 9 1 9 13 0 9 2 9 7 10 9 1 9 2
11 1 9 1 9 13 14 9 7 0 9 2
13 1 0 9 13 13 2 16 9 7 9 13 0 2
22 9 2 0 13 1 0 11 1 0 11 2 0 9 7 9 11 1 9 1 0 9 2
5 9 13 3 0 2
8 1 9 13 12 2 12 9 2
15 9 2 0 13 1 0 9 0 11 7 0 9 9 11 2
9 0 13 14 1 0 7 0 9 2
16 13 1 0 9 1 9 8 9 2 16 13 0 1 0 11 2
25 9 2 0 13 1 9 11 7 1 0 9 1 0 11 1 11 2 3 15 13 1 9 0 9 2
6 13 1 10 0 9 2
6 3 13 14 9 9 2
13 9 13 3 0 2 0 7 0 7 13 3 0 2
9 9 15 1 9 13 7 13 0 2
18 9 2 13 0 2 0 9 2 0 0 9 7 0 9 1 0 9 2
16 9 2 1 9 7 9 13 0 9 2 1 9 15 9 13 2
10 1 9 13 12 2 12 0 0 9 2
9 1 9 0 9 13 0 0 9 2
5 9 13 0 9 2
22 9 2 13 0 2 0 9 2 0 9 7 9 1 0 0 9 7 3 0 0 9 2
6 9 13 1 0 9 2
6 0 9 13 3 0 2
14 1 0 7 0 9 9 13 9 12 2 12 0 9 2
17 0 7 0 9 13 0 2 0 13 1 9 0 3 1 9 9 2
21 9 2 13 0 2 1 9 0 9 2 0 9 1 0 0 9 7 0 0 9 2
8 1 9 13 12 2 12 9 2
30 9 2 13 0 2 0 2 0 9 2 3 0 0 9 2 0 9 1 12 2 12 9 7 0 1 12 2 12 9 2
16 0 9 13 3 0 7 0 2 0 9 13 3 0 0 9 2
7 10 0 9 13 3 0 2
9 1 0 0 9 13 0 0 9 2
19 9 13 0 0 9 2 16 15 1 0 13 1 10 0 9 2 0 9 2
8 1 9 13 12 2 12 9 2
9 3 4 15 3 13 1 10 9 2
19 9 2 13 0 9 9 11 2 16 3 1 0 9 13 9 2 0 9 2
17 13 15 1 9 2 9 2 9 2 16 15 1 0 0 9 13 2
7 13 15 1 0 0 9 2
38 9 2 13 0 2 0 2 1 0 9 0 9 2 0 9 2 1 9 0 0 9 1 0 9 2 14 0 0 9 7 1 10 9 9 0 0 9 2
7 0 9 0 9 13 0 2
16 9 2 1 9 13 0 9 2 0 9 9 7 9 13 0 2
11 1 0 9 1 9 13 12 0 0 9 2
15 1 9 13 0 2 0 0 0 9 2 9 13 0 9 2
9 9 2 9 13 0 2 0 9 2
8 1 0 9 9 13 0 9 2
9 9 2 13 0 0 2 0 9 2
10 0 13 1 0 9 2 9 13 0 2
9 0 9 13 12 2 12 0 9 2
4 13 0 9 2
5 0 9 13 3 2
7 13 12 2 12 0 9 2
4 9 13 0 2
8 1 9 13 12 2 12 9 2
19 9 2 13 0 2 0 7 3 0 9 2 0 1 9 1 9 0 9 2
6 9 7 9 13 0 2
4 13 1 9 2
16 13 0 2 0 7 0 0 9 2 16 1 9 13 16 9 2
10 9 13 3 0 7 13 0 0 9 2
6 0 9 13 3 0 2
10 0 9 13 1 9 9 3 0 9 2
14 1 9 13 0 2 9 7 13 0 7 3 0 9 2
18 1 0 9 13 0 0 9 7 3 0 2 1 0 9 0 0 9 2
8 1 9 13 12 2 12 9 2
20 16 3 9 9 13 7 15 0 9 13 2 15 14 9 13 1 0 9 9 2
19 3 14 13 1 9 2 9 1 0 9 13 9 9 7 14 13 0 9 2
9 3 13 13 3 3 7 3 3 2
20 16 9 14 13 9 1 9 7 9 2 15 1 9 1 9 13 9 7 9 2
56 14 13 1 0 9 2 9 2 2 0 7 0 9 2 9 2 2 9 13 1 9 13 2 3 15 0 9 13 7 15 3 13 1 15 1 9 2 16 13 0 9 2 9 2 9 9 2 2 1 15 13 7 0 0 9 2
19 14 13 0 9 1 9 0 9 2 7 9 1 9 2 16 9 3 13 2
7 9 3 13 1 9 3 2
21 9 1 9 1 9 13 13 3 0 1 15 2 16 15 13 1 9 1 0 9 2
11 13 13 0 2 1 0 2 7 0 9 2
26 1 0 9 9 13 14 1 9 7 9 9 1 9 2 7 1 10 9 3 13 3 0 7 0 9 2
22 10 9 9 13 1 9 12 2 0 7 1 12 9 9 13 9 1 12 1 12 9 2
10 9 1 10 0 9 13 0 9 9 2
22 9 7 9 1 10 9 13 0 9 1 0 0 9 2 16 15 3 13 1 0 9 2
20 15 13 0 1 9 1 0 0 9 2 0 7 13 0 1 9 1 0 9 2
9 0 9 1 9 13 1 0 9 2
16 9 0 9 13 9 9 7 9 0 9 9 2 0 1 9 2
18 0 7 0 9 13 13 1 9 2 0 7 13 1 0 7 0 9 2
19 9 0 9 9 13 13 1 9 7 15 13 2 16 0 13 1 0 9 2
20 9 13 1 9 9 2 16 15 13 10 9 2 16 15 13 7 13 1 9 2
6 9 13 0 1 15 2
23 9 1 9 9 1 9 9 1 9 9 13 10 9 2 12 2 2 16 1 15 13 9 2
9 1 9 0 9 13 1 0 9 2
11 10 0 9 1 0 11 7 11 13 15 2
10 1 15 13 0 7 15 0 0 9 2
27 10 0 9 2 16 15 13 1 0 9 2 13 3 0 9 2 9 13 1 0 9 9 7 13 0 3 2
29 9 2 9 7 9 2 16 15 13 1 9 2 7 13 3 0 9 2 9 13 1 0 9 9 7 13 0 3 2
13 9 13 0 7 0 9 2 16 13 1 9 9 2
33 9 2 16 13 1 9 9 7 1 0 9 2 13 3 3 0 7 3 0 9 2 15 1 9 2 1 15 13 2 13 0 9 2
15 1 9 4 3 13 0 0 9 11 11 1 11 1 11 2
22 1 9 11 1 11 4 9 3 13 2 13 4 15 0 9 7 0 9 15 4 13 2
19 13 15 0 9 9 2 7 13 9 2 9 7 9 2 16 13 9 9 2
8 13 15 1 9 7 13 9 2
21 10 9 1 9 9 2 12 1 12 2 13 0 9 9 9 14 1 9 0 9 2
11 1 0 9 15 13 0 9 7 13 0 2
14 10 9 13 9 9 7 15 13 9 1 9 7 9 2
16 1 9 0 9 14 13 1 0 0 9 7 15 13 3 13 2
10 1 9 15 13 9 3 16 1 9 2
6 9 15 13 9 9 2
20 1 9 15 9 13 1 0 9 2 1 15 13 0 3 0 9 16 1 9 2
27 9 1 3 0 9 1 0 0 9 4 13 1 0 9 0 9 2 7 15 0 9 13 1 0 9 9 2
20 1 15 10 9 13 1 10 9 9 7 1 9 10 9 1 9 7 1 15 2
16 10 9 0 9 13 0 9 1 9 2 9 7 0 0 9 2
14 3 13 2 16 0 3 13 1 0 9 1 0 9 2
15 0 9 4 15 13 14 8 11 11 7 9 11 11 11 2
8 15 4 13 9 9 7 9 2
21 11 11 4 13 2 16 13 9 12 1 9 1 0 9 7 9 1 9 7 9 2
23 1 10 9 13 9 1 0 11 0 9 1 0 9 2 0 9 9 7 9 1 9 0 2
19 9 4 13 10 9 2 9 9 9 11 1 11 2 9 2 9 7 9 2
39 8 11 11 2 9 0 9 2 16 4 3 1 0 9 11 11 1 11 7 1 9 13 0 9 2 13 3 0 1 0 9 9 2 9 7 1 10 9 2
17 13 15 2 16 13 0 9 0 9 1 9 0 9 1 9 9 2
26 9 2 1 15 15 13 2 4 15 3 13 2 16 4 13 3 0 9 7 13 10 9 14 1 0 2
17 1 10 9 4 13 15 2 15 13 14 3 3 2 7 13 0 2
12 14 13 7 1 9 2 1 9 3 13 9 2
23 0 9 0 9 13 0 2 3 0 9 2 9 2 1 0 9 1 0 9 13 0 9 2
14 1 15 13 1 0 9 0 0 9 2 15 13 9 2
11 1 15 13 0 7 0 9 2 9 2 2
8 1 15 13 9 1 9 0 2
16 15 3 13 2 1 15 13 9 2 16 15 9 13 1 9 2
10 10 9 13 9 0 7 3 0 0 9
9 3 7 15 13 14 12 0 9 2
32 1 0 9 12 14 4 0 11 13 9 9 1 9 1 0 9 2 1 15 7 15 4 13 0 0 9 9 11 1 0 9 2
24 14 3 1 9 1 9 7 9 13 14 0 9 2 16 4 13 0 9 0 9 7 0 9 2
24 9 1 0 9 13 3 1 0 9 2 4 13 11 11 11 1 9 1 9 1 9 1 9 2
8 1 11 7 15 9 14 13 2
18 15 15 13 9 13 1 15 2 16 15 2 16 3 13 2 14 13 2
17 14 13 2 14 2 3 15 11 13 0 2 3 13 3 10 9 2
42 3 0 13 14 2 16 4 11 1 9 1 0 9 10 9 13 7 13 0 9 7 16 15 4 9 14 15 14 0 13 7 0 13 3 0 2 16 9 13 0 9 2
33 15 7 4 13 2 16 4 1 9 10 9 2 16 4 13 0 2 14 13 9 2 16 14 4 13 0 7 16 4 15 9 13 2
7 9 4 13 14 1 9 2
22 16 4 3 1 9 13 0 9 2 4 0 13 2 7 15 4 3 13 1 10 9 2
19 0 9 1 0 9 4 1 12 9 1 9 0 9 11 11 3 13 9 2
31 9 0 9 1 9 1 9 11 13 2 16 4 13 9 0 7 4 13 1 15 2 16 15 4 9 13 13 1 0 9 2
26 0 9 9 13 9 1 9 0 9 1 0 9 2 1 15 13 1 9 14 0 9 1 0 9 11 2
5 14 0 9 13 2
19 15 13 9 0 9 0 2 0 9 2 10 13 9 2 0 9 7 0 2
19 9 2 9 7 0 0 9 13 0 9 2 16 15 0 9 13 0 9 2
14 3 15 14 3 13 1 0 9 7 1 15 13 9 2
5 14 13 15 13 2
22 16 4 9 13 2 16 15 14 13 1 0 9 2 16 13 3 0 2 0 2 0 2
14 2 14 3 15 3 13 2 3 4 3 13 0 9 2
5 14 13 14 3 2
9 9 13 0 2 14 13 13 0 2
17 13 9 1 10 9 7 13 15 2 16 4 3 13 2 15 13 2
23 15 15 9 14 13 7 14 13 13 2 16 4 15 13 0 9 14 0 9 9 7 9 2
10 15 9 13 1 15 2 3 14 13 2
9 14 15 4 14 13 1 0 9 2
36 16 15 9 9 14 4 13 13 2 13 14 10 9 3 2 16 4 13 1 9 2 16 15 13 2 7 14 9 1 9 1 15 13 3 0 2
22 10 9 4 13 10 9 2 16 4 14 13 1 9 2 9 9 7 9 2 13 15 2
7 7 1 9 16 1 9 2
17 9 13 3 0 7 0 2 16 4 13 9 9 13 0 0 9 2
34 3 2 16 4 1 15 1 0 13 9 2 16 13 14 13 1 9 2 15 3 13 3 3 2 1 10 9 2 0 1 9 7 12 2
19 1 9 9 9 0 9 4 3 15 13 9 11 2 16 13 1 0 9 2
21 3 3 4 15 13 2 16 10 9 14 13 3 13 2 16 15 14 14 13 9 2
27 10 9 2 16 4 15 15 13 1 9 2 14 13 10 9 2 7 13 2 16 15 9 9 14 4 13 2
31 1 9 4 13 15 2 7 16 14 13 13 2 3 13 15 9 2 14 13 9 2 16 4 13 2 15 13 9 0 9 2
13 16 15 1 0 9 13 2 4 13 9 3 0 2
7 9 9 4 13 1 15 2
10 1 9 0 9 4 9 13 1 15 2
10 10 9 1 11 4 1 15 3 13 2
12 1 0 11 4 13 9 7 15 13 12 9 2
11 9 4 13 7 15 13 1 9 1 11 2
16 9 4 13 9 2 16 15 4 13 1 9 7 15 13 9 2
22 11 11 2 1 9 2 13 2 16 4 15 1 9 3 13 2 16 4 13 0 9 2
14 16 13 0 9 7 16 4 13 0 9 0 1 0 2
12 7 14 0 4 13 3 16 0 9 2 13 2
12 12 9 13 2 12 7 13 7 13 1 9 2
17 1 9 13 9 2 9 2 0 9 2 13 7 13 13 10 9 2
7 13 9 2 9 7 9 2
9 9 13 1 9 7 9 7 13 2
26 16 16 13 15 9 7 15 2 13 14 0 0 9 1 12 9 2 1 0 9 0 9 14 13 2 2
20 0 9 1 0 9 4 13 16 9 2 15 9 4 1 9 13 14 0 9 2
40 10 9 4 13 3 0 2 3 0 1 9 2 16 4 15 3 13 2 7 4 9 13 3 0 15 11 11 2 16 4 13 0 13 1 9 0 9 1 11 2
31 14 10 10 0 9 4 13 9 9 2 0 15 14 4 13 2 16 7 4 9 11 11 13 13 3 3 1 3 0 9 2
14 9 13 3 2 3 7 13 2 15 4 13 0 9 2
4 12 15 13 2
9 0 9 15 4 13 14 1 9 2
21 10 9 1 0 0 0 4 13 0 1 0 7 0 9 7 0 1 0 0 9 2
28 9 12 4 13 0 1 9 1 0 9 0 9 11 2 1 0 9 9 3 7 4 13 0 1 0 0 9 2
25 1 0 9 4 16 0 7 0 9 13 9 9 9 0 9 7 13 0 9 1 12 9 9 9 2
21 9 15 13 3 13 1 10 9 2 16 13 10 9 7 0 9 0 16 1 9 2
21 14 3 13 10 0 9 9 2 1 15 13 15 0 2 7 9 13 1 15 0 2
12 9 9 9 15 13 0 2 0 7 3 0 2
14 13 9 9 7 9 9 2 16 13 1 9 9 0 2
16 1 9 9 13 14 9 2 16 13 1 0 9 1 0 9 2
11 9 9 7 0 9 13 1 0 9 7 9
38 14 1 0 9 10 9 13 0 2 16 9 1 9 11 1 9 14 13 3 3 0 2 16 4 13 3 1 15 2 7 16 13 9 9 14 3 0 2
18 9 9 7 13 2 16 11 1 9 1 10 9 3 3 13 1 9 2
51 11 11 2 12 0 9 4 13 9 0 9 11 11 2 16 4 1 0 9 13 9 9 7 9 0 9 2 16 4 15 13 9 3 1 9 1 9 9 0 9 9 7 9 0 9 1 9 12 7 12 2
21 9 2 16 13 1 10 9 2 3 3 13 2 16 15 0 9 13 1 10 9 2
20 1 9 2 9 13 7 0 0 9 1 0 9 2 16 15 13 3 1 9 2
13 1 15 13 0 9 9 0 9 14 1 0 9 2
17 1 9 13 2 16 15 4 13 14 0 9 9 0 9 0 11 2
11 0 9 9 11 7 13 1 0 9 9 2
15 3 7 13 2 16 13 1 9 9 12 14 3 0 9 2
10 7 12 1 9 4 13 1 15 0 2
13 12 0 9 4 1 9 9 11 11 13 0 9 2
22 9 1 9 2 9 7 9 4 14 13 0 9 2 0 1 9 1 9 1 0 9 2
24 9 4 13 9 12 2 0 9 0 0 9 2 16 15 4 12 9 1 12 9 13 14 11 2
16 0 9 4 13 0 14 3 2 1 9 0 9 0 0 9 2
23 16 9 9 0 9 13 15 9 0 0 9 2 9 10 9 13 1 0 9 9 9 9 2
10 7 14 1 10 9 13 0 0 9 2
19 9 0 9 1 9 0 7 0 9 7 10 0 9 15 4 7 13 3 2
30 2 14 13 3 2 16 4 13 1 9 7 3 1 9 7 3 0 0 9 2 7 1 10 9 4 13 9 3 3 2
27 13 2 16 4 13 0 9 1 9 9 12 0 3 2 13 7 4 9 1 0 9 1 9 7 1 9 2
20 3 10 0 9 14 14 13 2 15 13 9 12 2 2 13 11 11 1 11 2
12 7 9 9 13 7 0 7 0 9 0 9 2
17 11 4 1 9 13 10 9 2 16 3 13 0 1 0 0 9 2
14 3 7 4 14 3 13 9 9 7 3 13 0 9 2
7 9 1 15 14 13 9 2
26 16 4 9 13 2 7 16 4 1 9 13 0 9 3 7 3 2 4 1 10 9 9 13 1 9 2
4 8 8 8 2
38 16 13 9 2 16 4 13 0 1 9 2 9 0 9 2 2 15 1 10 9 2 9 2 9 2 9 7 9 2 16 4 15 13 2 14 3 13 2
4 7 3 3 2
3 3 3 2
11 16 4 13 2 15 4 13 0 0 9 2
11 16 4 13 2 15 4 3 13 0 9 2
9 16 4 13 2 15 4 13 9 2
9 14 2 9 4 1 15 13 9 2
23 0 9 13 3 3 0 2 7 0 1 3 0 9 2 7 15 13 3 1 10 9 13 2
14 9 13 0 2 7 13 14 9 9 9 7 9 9 2
25 9 13 0 1 0 9 1 0 9 7 0 9 7 1 0 9 0 9 2 16 13 9 1 9 2
22 0 9 13 0 9 1 0 9 2 16 3 1 9 13 9 7 9 9 1 0 9 2
13 9 13 9 2 0 0 0 2 0 7 0 9 2
18 10 0 2 0 9 15 13 9 1 9 2 16 13 3 0 1 9 2
29 16 9 9 13 7 13 1 9 2 15 9 13 1 0 9 2 1 15 13 9 2 7 9 13 14 0 0 9 2
41 1 9 7 9 9 13 1 11 3 0 9 11 1 11 2 7 1 10 0 9 9 1 9 7 10 9 4 3 13 1 11 14 12 2 16 15 1 15 14 13 2
8 3 4 13 14 0 2 2 2
11 9 13 12 3 7 1 9 15 13 13 2
5 1 9 13 0 2
6 11 13 14 3 0 2
12 1 0 12 9 4 15 13 1 0 10 9 2
27 1 9 13 1 9 1 12 2 9 1 9 2 2 16 3 13 3 3 2 7 10 9 4 15 3 13 2
5 9 13 3 15 2
2 8 2
2 8 2
3 0 9 2
6 13 7 14 1 9 2
12 1 0 9 13 0 9 2 15 9 4 13 2
42 16 15 13 2 16 4 13 14 0 9 2 9 7 9 2 13 0 9 1 9 7 9 7 9 2 1 15 1 0 9 2 16 4 13 9 2 13 1 12 9 9 2
31 9 2 16 15 13 2 16 9 13 3 2 7 0 9 13 2 16 9 13 1 9 7 16 9 3 13 1 15 7 13 2
15 1 15 9 13 2 16 15 14 13 1 15 1 9 9 2
14 3 16 1 9 1 9 7 9 1 9 7 1 9 2
13 9 1 9 13 15 3 0 7 0 1 10 9 2
16 14 4 13 13 2 16 13 9 3 2 7 13 15 13 0 2
16 15 9 2 16 15 4 13 7 13 2 15 4 13 10 9 2
40 2 11 11 2 0 9 2 16 13 1 0 9 0 1 10 9 2 3 14 13 1 9 2 7 1 9 13 2 16 13 10 9 0 7 16 13 9 1 9 2
17 7 1 15 13 0 2 7 13 0 9 9 2 16 15 13 3 2
9 9 4 3 13 10 9 1 9 2
17 2 14 13 2 3 4 13 2 2 15 4 13 1 3 0 9 2
16 3 15 4 13 1 0 9 2 16 15 4 13 1 0 9 2
30 11 4 14 3 13 1 9 1 3 12 2 15 4 13 13 3 1 12 1 0 9 2 16 4 13 9 1 0 9 2
6 3 4 15 3 13 2
16 11 4 13 1 9 7 13 9 11 2 16 4 13 1 9 2
17 0 4 13 2 16 4 13 2 16 13 1 9 10 9 7 9 2
33 2 9 11 4 13 2 16 4 10 9 11 2 0 1 0 9 11 11 2 3 13 1 9 1 9 11 12 2 2 4 13 11 2
24 9 2 16 15 11 12 14 13 14 3 1 9 2 15 4 13 0 2 14 0 9 1 9 2
35 11 2 16 4 13 9 1 9 2 16 4 13 0 2 16 15 4 13 2 15 4 13 3 2 13 9 1 9 7 13 0 9 1 9 2
29 14 13 2 15 4 13 15 2 7 3 13 2 16 4 13 13 0 1 15 2 15 4 14 13 11 7 10 9 2
16 11 4 1 9 13 2 3 7 4 13 2 16 4 9 13 2
8 3 4 13 13 0 1 9 2
44 16 15 4 1 9 13 3 2 4 13 2 16 4 15 14 3 13 9 7 13 0 0 9 2 7 16 15 4 13 1 15 2 4 3 13 2 16 3 13 0 9 1 15 2
11 14 3 15 15 4 13 0 9 3 0 2
14 1 9 3 4 11 11 1 9 13 0 9 9 11 2
12 2 3 13 1 9 2 2 15 4 13 0 2
16 3 4 3 11 13 1 10 9 13 10 9 2 15 4 13 2
24 14 0 4 13 14 3 2 16 4 1 9 9 0 9 14 13 7 14 3 13 9 0 9 2
7 9 1 9 4 13 0 2
16 11 4 3 13 7 3 13 9 2 16 15 4 13 1 9 2
21 2 14 13 15 3 3 1 9 2 13 7 2 16 15 1 9 14 13 1 9 2
12 16 13 3 0 2 15 3 14 4 3 13 2
16 14 16 4 15 13 2 4 13 11 1 9 7 13 1 9 2
9 13 15 4 0 9 7 15 13 2
7 1 9 4 13 9 11 2
15 1 0 9 4 13 1 0 9 9 9 7 9 0 9 2
21 2 7 4 13 0 9 7 7 4 15 1 9 1 0 9 15 13 1 9 9 2
26 13 4 9 15 15 2 9 1 0 9 2 16 15 4 13 3 13 2 16 15 15 4 13 0 13 2
20 1 0 0 9 7 1 0 9 4 13 2 16 13 15 2 15 13 2 9 2
24 1 10 9 4 13 0 9 9 9 2 16 15 11 3 13 1 0 9 1 9 7 9 9 2
16 11 2 12 2 3 14 4 1 0 9 13 0 9 9 9 2
3 2 9 2
27 0 9 13 1 9 3 2 16 4 9 1 0 9 12 0 9 13 9 0 9 0 9 1 11 7 11 2
5 13 4 14 9 2
3 2 8 2
15 15 15 7 4 13 0 1 9 0 9 7 9 0 9 2
6 7 7 13 1 11 2
13 11 2 12 2 0 0 9 13 14 1 10 9 2
26 0 9 7 9 0 9 14 3 13 10 9 9 0 9 2 16 13 3 1 0 9 3 14 14 0 2
16 3 9 13 1 0 9 16 1 9 1 10 0 0 9 11 2
28 1 10 9 4 13 10 9 1 9 9 9 2 16 13 14 0 2 13 0 9 1 9 10 9 9 0 9 2
35 3 13 14 0 0 9 2 9 2 2 16 4 0 0 9 1 3 3 7 3 13 3 10 0 9 7 0 0 9 13 1 10 0 9 2
32 11 2 12 2 0 2 0 9 11 2 11 4 1 9 1 0 9 1 11 7 9 11 8 8 8 13 9 1 9 0 9 2
19 11 2 12 2 1 9 4 1 9 0 9 3 13 9 11 11 11 11 2
25 9 7 4 15 3 1 9 13 1 0 9 2 7 4 1 9 13 1 9 9 0 9 11 0 2
25 1 0 9 4 3 1 9 13 11 0 2 16 4 1 10 9 14 13 14 1 10 0 0 9 2
31 1 9 4 11 3 1 9 11 1 0 11 1 11 13 0 9 1 0 9 2 16 4 13 0 0 12 2 9 3 0 2
25 1 9 4 13 9 1 11 2 11 7 11 7 1 15 3 13 1 9 10 9 1 0 0 9 2
13 11 11 2 3 15 9 13 11 12 7 11 12 2
9 0 13 3 0 9 9 1 9 2
12 15 0 13 2 16 15 1 9 13 0 9 2
7 15 13 14 1 0 9 2
14 14 7 13 1 9 0 9 1 0 0 7 0 9 2
11 0 9 13 3 0 9 2 16 13 9 2
12 11 15 4 13 1 11 7 3 13 10 9 2
25 9 12 4 13 14 1 11 2 16 15 4 9 8 11 13 2 16 15 4 13 13 1 0 9 2
28 14 16 15 4 13 1 0 9 11 11 2 12 2 2 15 4 13 9 2 16 4 13 10 9 3 14 0 2
12 9 4 15 13 1 9 2 16 4 14 13 2
14 10 9 4 13 10 9 2 16 4 13 10 0 9 2
39 1 0 9 9 2 1 12 9 2 4 11 11 2 11 11 7 11 11 13 1 0 9 0 9 2 16 4 13 1 0 9 0 9 7 0 9 10 9 2
14 15 4 13 1 0 9 7 9 4 3 13 1 9 2
12 1 9 0 9 13 0 3 12 9 9 9 2
21 1 11 13 14 3 1 12 9 9 1 0 9 1 9 1 9 0 9 1 9 2
18 14 9 9 13 9 1 9 2 16 4 13 1 0 9 1 9 9 2
13 1 11 10 9 14 13 2 3 13 14 1 11 2
20 16 13 1 0 9 2 15 0 9 13 1 0 9 2 16 13 14 0 9 2
17 2 1 15 4 15 14 13 1 9 2 16 13 9 0 7 0 2
11 9 9 4 13 11 11 1 0 9 11 2
10 10 0 9 15 13 1 3 12 3 2
16 2 10 9 13 9 7 9 2 13 7 14 1 0 0 9 2
20 1 9 13 2 16 13 9 0 9 2 7 1 9 13 2 16 13 0 9 2
51 9 2 0 9 13 2 16 13 9 9 9 13 7 15 13 9 0 9 2 16 13 1 0 9 10 9 2 7 9 2 16 13 1 10 9 2 16 15 13 7 16 15 1 10 9 14 13 9 0 9 2
20 1 15 13 0 14 9 0 9 2 9 2 0 9 2 2 16 13 10 9 2
3 2 8 2
14 0 9 1 11 13 1 0 9 3 3 0 0 9 2
26 14 3 7 13 10 12 9 0 9 0 12 1 9 1 9 9 2 16 3 13 0 9 9 1 9 2
14 1 10 9 4 13 9 1 9 9 9 1 9 9 2
15 0 4 13 9 2 3 13 9 1 9 1 9 0 9 2
19 13 15 2 16 13 1 9 3 0 2 15 15 7 3 13 1 0 9 2
12 3 13 1 0 9 0 0 1 0 7 0 2
36 14 0 13 2 16 0 9 2 0 1 0 9 2 13 0 9 7 16 1 15 3 13 15 15 7 15 0 2 7 4 15 13 1 0 9 2
5 13 7 0 9 2
13 3 13 14 15 2 16 4 3 13 9 0 9 2
2 3 2
21 14 15 3 1 9 9 13 0 9 7 3 13 1 9 9 7 14 14 0 9 2
24 13 15 13 2 7 1 9 10 9 7 0 15 9 15 3 14 13 13 2 1 10 9 13 2
27 0 13 2 16 13 10 0 9 2 16 15 13 1 0 9 3 2 16 13 0 13 9 7 9 10 9 2
8 14 3 13 0 9 14 13 2
13 10 0 9 4 13 0 9 7 4 13 10 0 9
17 11 1 0 9 0 9 0 9 9 1 9 9 4 13 3 3 2
12 0 9 4 7 14 3 13 14 3 10 9 2
17 1 15 15 15 4 13 9 7 9 4 3 13 1 9 7 9 2
22 11 7 11 4 14 9 12 13 9 2 1 15 13 9 0 9 7 9 1 0 9 2
29 0 0 9 11 11 11 1 0 9 13 11 2 16 14 13 1 0 0 9 2 16 13 1 9 0 9 0 9 2
10 13 1 0 9 2 16 13 10 11 2
15 7 12 9 3 14 13 13 15 2 15 15 4 3 13 2
20 9 4 13 1 0 14 1 12 1 9 0 9 1 9 11 11 11 1 11 2
21 0 9 13 3 0 2 7 15 4 1 1 9 1 0 9 13 1 0 9 9 2
43 1 0 9 2 16 15 4 13 1 12 9 2 4 1 0 9 13 0 9 1 9 9 2 1 0 9 7 13 1 9 9 11 0 9 2 16 15 4 1 9 13 9 2
13 9 11 15 4 3 1 10 9 13 1 9 9 2
3 2 8 2
11 9 13 0 1 9 11 1 0 9 12 2
39 3 1 0 9 13 9 9 1 9 2 1 15 4 13 11 11 2 11 11 2 11 11 2 11 11 2 11 11 7 0 9 9 0 9 0 9 0 9 2
19 1 9 2 12 9 2 1 12 9 13 0 9 0 9 7 0 9 9 2
6 9 9 13 11 11 2
14 7 1 12 9 1 9 1 11 15 3 13 14 15 2
45 11 11 4 13 0 0 9 2 7 3 15 13 9 2 15 4 13 11 2 16 11 1 9 9 2 16 13 14 12 9 0 9 2 13 14 1 12 9 7 13 9 1 0 9 2
14 9 13 15 0 2 7 13 0 1 9 0 9 11 2
13 0 9 13 11 11 2 13 9 0 9 11 11 2
9 9 13 1 0 9 0 1 9 2
12 15 0 13 3 0 2 7 15 9 14 13 2
14 16 13 3 1 9 7 15 13 2 15 13 0 13 2
10 9 13 9 0 9 1 0 9 7 9
17 1 0 0 9 1 0 9 15 4 11 11 13 1 11 11 11 2
28 9 1 0 9 1 11 4 13 0 1 9 0 9 2 16 4 3 13 0 9 9 2 16 4 13 0 9 2
14 16 2 9 2 13 1 10 9 12 0 14 11 11 2
11 15 4 1 10 9 13 14 1 0 9 2
17 14 12 9 3 11 11 3 13 12 9 9 2 15 9 4 13 2
26 3 15 13 1 10 9 7 0 9 2 16 4 15 3 1 0 9 9 13 2 16 15 4 9 13 2
10 9 9 4 3 13 10 9 1 9 2
24 9 13 2 16 14 13 0 2 16 4 9 1 10 9 13 14 3 2 7 13 9 0 9 2
17 9 9 2 0 9 16 9 9 2 15 13 3 1 9 0 9 2
44 3 0 1 10 9 0 9 13 2 16 13 9 15 2 16 13 9 1 9 9 7 14 13 9 9 2 3 7 9 14 13 2 3 16 13 10 9 1 0 9 0 9 9 2
19 9 9 2 16 13 9 0 1 0 9 2 1 9 7 1 9 13 9 2
31 1 0 9 11 11 9 11 13 13 0 9 9 14 1 9 0 9 2 16 4 13 9 13 9 2 16 4 13 13 0 2
36 14 0 9 13 13 1 0 9 2 16 13 9 9 9 2 16 15 4 9 12 13 9 11 11 1 9 9 1 9 9 2 9 7 0 9 2
26 10 9 4 13 14 1 9 2 16 4 14 9 9 13 1 9 2 16 7 14 4 13 1 10 9 2
39 0 9 4 1 3 10 9 13 9 1 11 2 14 16 4 13 1 9 2 16 4 14 10 0 9 13 16 9 7 4 10 9 14 3 13 14 1 9 2
19 13 4 1 0 9 2 7 16 4 13 0 9 2 15 15 4 9 13 2
31 13 15 4 1 9 7 3 13 2 16 16 0 2 0 9 14 4 13 13 2 7 4 15 3 3 13 7 3 14 13 2
10 13 15 4 13 7 15 13 0 9 2
25 9 15 4 13 1 0 7 15 13 14 1 0 9 1 0 9 2 16 4 15 13 1 0 9 2
19 16 4 1 9 13 11 2 4 15 13 10 9 7 14 3 13 10 9 2
11 11 4 13 10 9 2 7 4 3 13 2
18 16 4 13 14 15 2 4 0 9 13 10 0 9 0 9 1 9 2
15 9 4 13 9 2 16 4 13 9 1 10 9 1 11 2
11 9 4 13 0 1 9 9 1 0 11 2
19 11 11 4 13 3 0 1 11 2 16 15 4 3 13 9 1 10 9 2
19 3 1 9 1 10 0 9 13 0 9 2 1 15 13 0 9 0 9 2
10 9 4 11 13 2 9 1 9 2 2
7 8 8 8 8 8 8 2
9 8 8 8 8 2 12 2 12 2
4 8 8 8 2
4 8 8 8 2
7 8 8 8 8 8 8 2
4 8 8 8 2
29 13 9 0 9 2 12 9 2 12 9 0 9 2 10 9 2 12 9 9 2 12 9 0 9 2 12 9 9 2
11 0 9 14 13 2 3 15 4 3 13 2
23 1 9 0 9 7 4 13 10 9 0 2 7 13 14 15 14 9 1 0 7 0 9 2
33 1 9 7 1 11 3 14 13 15 2 16 13 9 1 11 0 1 0 9 7 16 4 3 14 15 3 13 10 10 2 9 2 2
15 10 16 12 0 9 4 1 12 9 3 13 1 0 9 2
28 9 13 2 16 4 15 3 13 0 9 2 16 4 13 1 0 9 2 13 2 9 7 13 10 2 9 2 2
44 1 11 7 4 13 9 14 14 1 9 2 7 14 1 0 9 16 4 9 2 16 4 15 1 9 13 9 7 9 2 3 13 12 9 3 7 15 3 13 1 0 0 9 2
24 3 13 13 2 16 13 1 9 10 0 9 2 16 15 3 7 3 13 2 3 3 13 9 2
8 15 7 10 9 13 15 0 2
11 1 0 12 9 4 15 10 9 3 13 2
24 15 13 2 16 10 9 13 2 16 13 3 13 13 1 9 14 1 0 9 9 9 1 9 2
37 0 9 1 9 9 1 0 9 9 1 9 15 14 10 9 13 2 7 16 4 13 0 13 9 3 2 16 13 9 3 3 3 2 16 13 0 2
7 0 9 15 3 3 13 2
33 0 0 9 4 7 13 2 16 3 3 3 3 13 9 2 16 4 13 9 2 16 4 15 13 7 16 13 1 9 3 14 0 2
7 9 9 3 4 13 0 2
21 1 9 1 9 3 0 13 9 2 16 4 13 9 15 9 7 9 0 7 0 2
14 3 15 13 1 9 2 9 2 9 2 16 14 13 2
19 9 9 14 13 0 16 1 9 1 9 2 7 3 3 13 10 9 9 2
7 3 4 1 10 9 13 2
15 3 15 4 15 1 0 9 13 2 16 4 9 9 13 2
12 2 14 15 4 13 2 16 4 14 13 9 2
32 3 7 4 10 9 7 15 13 14 3 13 2 16 13 1 9 1 9 7 16 13 0 2 16 13 3 0 2 3 13 2 2
15 7 4 3 13 2 15 15 15 14 15 1 10 9 13 2
3 7 13 2
4 16 14 13 2
7 9 13 1 0 9 9 2
7 1 9 9 13 0 9 2
27 16 9 13 9 2 9 7 9 2 15 3 13 1 9 0 9 2 16 13 0 9 2 9 2 0 9 2
16 16 10 9 14 13 0 0 0 9 2 13 3 0 9 0 2
14 16 13 9 7 9 2 13 3 2 16 15 13 9 2
11 9 3 13 2 16 4 13 1 10 9 2
11 1 9 13 14 0 2 7 14 13 13 2
29 0 13 2 16 9 13 9 7 13 3 13 10 10 9 7 9 2 7 13 14 3 0 2 16 13 1 10 9 2
10 3 4 13 10 3 0 9 16 3 2
13 13 13 3 1 2 0 2 7 2 0 2 9 2
16 1 0 9 13 13 1 0 9 9 2 0 1 9 0 9 2
35 11 11 2 16 4 1 12 9 13 1 0 9 2 15 4 13 0 9 2 0 9 0 9 2 0 0 2 9 2 7 9 9 1 9 2
34 9 3 4 1 9 13 9 2 9 7 4 13 3 0 1 0 11 2 16 4 9 11 12 13 13 14 9 2 16 14 13 0 9 2
24 9 0 9 13 1 10 9 0 9 2 9 7 13 14 0 9 7 13 14 3 0 0 9 2
11 2 3 13 1 9 2 2 4 13 9 2
17 2 13 4 9 1 9 2 16 13 9 2 3 7 15 13 9 2
14 2 1 9 4 15 13 1 11 2 2 4 13 11 2
17 2 7 4 13 9 2 11 7 1 9 14 4 13 13 0 9 2
23 13 4 10 10 9 7 16 9 4 13 14 2 15 4 11 13 2 16 4 13 0 9 2
12 14 15 15 4 13 3 2 7 4 13 13 2
10 15 7 14 4 13 9 10 0 9 2
13 9 8 11 11 4 3 13 1 11 11 1 11 2
25 0 9 4 1 15 13 9 0 9 7 14 0 9 2 15 3 4 13 1 9 9 1 10 11 2
6 0 4 13 0 9 2
17 10 9 13 16 0 9 2 7 4 1 9 3 13 0 12 9 2
21 14 3 13 0 1 0 2 3 0 9 2 16 13 1 9 9 2 1 12 9 2
6 3 4 15 13 0 2
14 15 2 15 15 15 4 13 2 4 13 13 1 0 2
11 14 9 15 14 4 13 13 14 1 9 2
17 3 13 1 9 2 16 13 0 2 0 7 15 4 13 1 9 2
10 1 9 13 0 7 13 13 3 3 2
31 15 13 1 0 9 7 0 9 2 0 0 9 0 9 1 9 0 9 2 10 0 9 2 16 14 4 13 9 0 9 2
6 10 0 9 13 9 2
7 15 7 13 0 9 11 2
2 9 2
19 13 3 1 9 9 0 2 14 15 14 14 13 0 15 9 7 0 9 2
7 0 9 4 3 14 13 2
24 1 3 14 3 3 0 0 9 11 2 1 15 15 14 13 9 3 0 9 2 13 15 0 2
10 9 1 9 1 9 13 14 0 9 2
25 2 13 4 14 9 2 3 3 7 4 13 9 7 13 2 16 13 7 16 13 13 1 12 9 2
15 3 15 4 13 0 2 16 16 4 13 0 9 7 13 2
12 14 2 16 15 13 13 2 15 4 13 3 2
22 1 0 9 15 9 10 9 9 14 13 13 2 14 16 4 15 13 1 0 9 9 2
19 7 15 4 14 13 1 9 1 0 9 1 11 2 16 13 1 0 9 2
14 9 1 0 11 4 13 15 3 0 2 16 13 0 2
15 2 3 4 13 15 13 3 2 7 4 13 13 0 9 2
14 3 4 13 0 10 9 2 1 15 4 15 13 0 2
9 0 9 4 13 15 9 1 9 2
6 2 15 4 13 13 2
13 3 13 2 16 15 9 3 3 13 1 10 9 2
9 2 14 13 0 15 13 1 9 2
12 13 3 3 2 14 1 9 15 13 1 9 2
14 3 15 13 1 0 9 7 13 1 0 9 1 15 2
2 9 2
7 3 14 13 2 13 9 2
10 3 15 13 2 13 7 13 1 9 2
5 9 7 14 13 2
14 15 13 2 16 13 15 10 9 9 2 16 15 13 2
8 13 15 7 15 13 1 9 2
14 12 9 13 14 2 16 4 15 13 1 9 1 11 2
17 9 0 9 1 9 9 9 4 13 9 1 0 0 9 1 11 2
13 13 1 9 1 9 2 1 9 7 1 0 9 2
14 11 15 1 15 13 1 0 9 1 0 9 0 9 2
14 0 9 15 13 9 1 9 7 1 9 7 0 9 2
45 0 13 9 2 16 4 15 13 9 1 9 0 0 9 1 0 9 7 0 9 1 0 0 2 9 1 0 9 1 0 9 13 2 16 4 1 10 9 13 3 13 1 0 9 2
16 0 7 4 13 14 3 9 1 9 9 2 1 12 9 9 2
15 1 9 9 7 1 9 7 9 10 9 11 15 4 13 2
4 0 7 0 2
13 11 2 15 13 2 16 14 4 3 15 3 13 2
21 11 4 3 13 9 2 13 15 4 1 0 0 9 2 16 13 0 9 7 9 2
26 0 4 13 1 0 9 2 9 1 9 1 10 9 2 1 9 4 3 13 7 1 11 16 1 9 2
18 1 0 9 3 13 0 9 0 9 1 0 0 7 0 9 11 11 2
16 11 4 3 1 11 13 1 11 1 9 9 0 9 11 11 2
24 9 15 3 3 13 1 9 0 9 2 14 3 16 13 2 16 1 0 9 3 13 14 11 2
27 1 0 9 4 0 9 13 14 10 9 2 16 4 1 9 13 0 9 7 13 10 0 9 9 0 9 2
19 11 11 7 4 0 0 9 13 1 0 9 2 1 9 0 11 11 11 2
17 11 4 9 13 9 1 12 9 2 7 4 13 1 0 12 9 2
16 11 2 16 4 13 1 9 12 9 2 7 4 13 0 13 2
19 0 11 4 1 0 9 13 14 12 9 7 13 0 9 13 9 11 11 2
18 6 2 3 4 13 3 1 15 2 3 1 10 0 9 14 3 13 2
24 7 4 13 14 13 2 11 13 14 1 11 7 15 14 3 13 2 15 15 13 1 10 9 2
4 15 13 3 2
9 1 9 9 13 9 2 16 13 2
10 10 9 13 3 0 1 9 1 9 2
17 16 13 9 0 2 13 3 3 2 1 9 9 7 1 0 9 2
17 9 7 9 13 1 9 9 2 9 9 7 14 13 1 9 9 2
6 1 15 13 0 9 2
5 13 1 9 9 2
5 9 14 13 0 2
10 14 3 2 13 0 9 9 7 9 2
3 9 9 2
3 9 9 2
8 1 11 4 15 13 7 13 2
31 1 11 9 2 9 9 2 15 4 13 0 9 2 16 4 15 13 1 9 2 15 13 1 9 7 15 13 1 0 9 2
26 13 7 4 14 1 9 2 9 9 0 9 4 13 9 2 0 1 10 9 2 16 4 3 13 9 2
9 1 0 0 9 4 13 0 9 2
15 1 10 9 9 4 13 1 9 11 10 9 1 0 9 2
19 1 0 9 15 4 13 9 2 16 15 4 14 1 0 9 13 0 9 2
14 0 9 15 4 13 1 9 2 16 15 4 13 9 2
7 7 15 11 4 13 0 2
19 14 16 15 15 4 13 1 9 7 9 10 9 2 15 4 13 0 9 2
16 12 15 4 13 2 16 15 4 13 3 3 2 1 2 2 2
37 0 9 2 3 13 12 3 2 0 2 0 9 2 14 1 12 1 12 9 7 4 15 1 9 9 0 9 8 11 11 3 13 14 1 0 9 2
39 11 2 1 9 2 16 4 15 13 1 0 9 9 7 9 2 4 1 0 9 1 9 2 16 15 13 2 13 12 9 2 0 14 4 13 10 9 3 2
21 1 0 9 4 10 9 14 13 9 2 9 7 14 4 13 14 1 9 10 9 2
13 9 13 0 1 9 11 7 11 2 9 13 0 9
33 1 9 1 9 9 7 9 0 9 1 0 9 9 13 0 9 9 2 16 13 1 10 9 7 15 14 1 0 9 13 1 9 2
19 9 9 9 7 0 9 11 4 13 1 12 9 1 10 9 1 10 9 2
12 9 9 1 9 15 13 1 0 7 0 9 2
13 1 10 9 9 9 7 13 13 0 9 1 9 2
24 13 4 14 2 16 4 13 0 9 14 9 9 2 1 0 9 7 13 0 7 1 9 9 2
46 3 16 9 1 0 9 4 0 9 3 13 14 9 0 9 1 9 2 7 4 13 0 2 16 4 1 9 1 9 13 1 10 9 9 2 16 13 9 7 9 9 1 9 1 9 2
13 3 4 0 9 10 9 13 1 9 9 9 9 2
10 9 4 0 9 10 9 13 0 9 2
12 9 1 9 14 3 13 1 9 9 1 0 9
12 1 9 1 0 9 4 11 3 13 9 11 2
20 11 4 13 3 0 7 13 2 16 9 13 9 0 9 2 7 9 1 0 9
9 1 11 13 10 9 1 0 9 2
19 13 15 4 2 16 13 0 9 3 0 2 16 4 3 13 1 10 9 2
18 11 3 13 2 15 15 4 13 2 16 13 1 11 3 0 0 9 2
19 11 4 3 1 11 13 0 0 9 1 9 0 9 1 9 12 1 12 2
12 1 11 7 1 0 9 13 3 0 1 9 2
33 9 0 9 4 13 2 16 13 0 9 13 1 0 9 2 3 4 14 13 2 16 13 0 9 3 3 0 16 9 1 10 11 2
16 11 4 1 9 14 13 2 16 13 1 9 9 3 0 9 2
36 0 9 4 13 14 1 12 9 2 0 9 7 4 1 9 13 13 10 1 12 9 2 16 4 15 1 10 9 9 14 13 13 14 0 9 2
10 0 13 2 16 15 4 13 3 0 2
4 3 3 13 2
19 3 2 16 4 1 0 9 13 9 3 2 13 15 9 7 9 10 9 2
14 13 7 4 1 0 9 2 15 7 9 15 13 3 2
16 3 1 12 9 4 9 13 9 2 16 4 14 3 13 13 2
10 1 10 9 15 4 11 13 0 9 2
14 3 9 4 15 13 1 9 2 4 13 0 11 11 2
18 13 9 9 11 2 11 2 16 15 1 11 13 3 1 11 7 3 2
7 3 0 9 9 1 11 2
28 15 13 9 1 9 0 9 2 14 7 13 9 1 9 0 9 7 9 0 9 2 16 15 13 1 10 9 2
42 13 15 15 2 16 9 9 2 16 15 9 13 1 9 1 0 9 2 13 3 1 9 7 16 2 16 13 9 9 0 2 13 13 10 9 2 16 13 1 0 9 2
11 1 9 1 11 4 13 10 16 12 9 2
16 9 4 15 13 2 13 4 12 0 7 12 0 7 0 9 2
18 0 9 4 15 13 14 9 12 9 2 0 4 13 0 10 0 9 2
15 9 9 4 15 13 14 3 7 4 13 12 1 12 9 2
18 13 4 15 1 0 9 2 1 0 9 1 0 9 1 11 7 3 2
51 16 4 1 0 9 10 0 9 1 11 13 2 16 15 13 13 1 11 2 4 15 13 1 10 9 2 16 16 13 1 9 9 2 7 15 13 2 16 15 1 10 0 11 9 13 7 13 1 0 9 2
13 1 9 4 11 11 13 0 7 0 9 1 9 2
14 10 9 4 13 7 13 1 9 2 16 15 4 13 2
12 9 4 13 3 0 7 4 15 13 1 9 2
47 9 11 1 9 1 0 9 1 9 1 9 2 12 9 2 1 12 9 1 9 9 12 0 9 13 1 9 9 11 11 1 9 9 1 9 2 1 15 13 13 9 1 9 9 11 11 2
26 1 9 4 13 14 11 11 2 9 9 2 11 8 11 2 11 11 7 11 11 2 9 7 13 0 2
56 9 11 4 13 15 2 16 15 4 1 11 13 0 9 9 7 16 13 0 9 14 3 3 0 2 4 1 0 9 1 0 9 13 9 9 11 8 11 11 2 16 1 0 0 9 13 9 9 7 9 9 1 0 0 9 2
15 16 4 14 13 2 4 1 9 11 1 0 9 9 13 2
25 0 9 15 4 13 0 0 0 9 2 16 4 13 1 9 0 9 7 0 0 7 0 9 9 2
27 9 11 11 11 13 0 9 0 7 0 9 2 0 1 0 9 0 9 2 16 15 9 13 3 9 9 2
3 2 8 2
26 3 15 15 3 13 1 15 2 15 15 4 13 1 0 0 9 7 14 1 0 9 1 11 2 2 2
3 15 0 2
29 9 13 14 1 15 2 16 1 0 9 11 7 11 4 13 9 1 11 2 7 4 15 3 3 13 14 1 15 2
19 9 1 9 0 11 13 14 0 2 1 15 14 4 0 0 9 13 1 9
28 2 1 9 0 9 13 10 9 1 9 12 2 3 0 4 13 14 9 1 10 9 1 9 1 11 7 11 2
13 13 4 9 9 1 9 2 13 3 3 7 13 2
34 3 15 4 3 13 0 9 0 9 11 2 16 14 4 13 1 9 0 9 1 9 0 9 2 3 16 4 1 9 13 9 11 11 2
20 7 1 9 1 0 9 4 9 11 11 11 11 3 13 9 1 9 10 9 2
24 1 10 9 13 0 9 2 16 3 9 1 9 14 14 4 13 7 16 4 3 13 13 9 2
22 2 3 10 9 4 13 10 0 9 2 1 15 15 4 13 2 2 4 13 11 11 2
10 2 3 13 1 0 9 1 11 11 2
12 2 11 4 1 10 9 13 3 14 1 9 2
28 11 11 4 13 1 9 1 0 9 2 1 0 9 1 9 4 13 2 16 2 4 3 13 0 1 15 2 2
10 10 9 4 1 0 9 13 9 0 9
24 1 2 0 9 2 4 13 14 11 11 1 0 0 9 2 16 4 13 12 0 7 0 9 2
21 9 1 9 11 11 13 2 16 1 9 1 0 0 9 9 0 9 9 13 0 2
15 1 0 9 15 9 13 14 1 9 1 9 9 0 9 2
37 1 9 1 9 9 9 13 1 10 9 0 2 16 9 11 13 2 16 1 11 13 10 0 9 2 11 2 2 16 4 13 2 16 4 13 0 2
25 10 9 13 9 9 9 2 9 0 9 2 16 13 0 1 9 9 2 7 9 9 15 1 11 2
17 0 9 11 4 10 9 13 9 11 2 10 9 7 4 13 9 2
24 0 0 9 15 4 3 13 1 11 2 1 0 9 2 16 4 13 14 1 0 9 1 9 2
27 3 13 1 9 9 0 2 16 15 4 1 11 1 9 13 14 0 0 9 2 15 9 4 13 0 9 2
9 10 9 13 9 0 9 0 9 2
3 2 8 2
36 9 0 13 14 0 9 9 9 11 2 7 13 0 9 0 0 9 7 15 13 1 0 9 1 9 9 7 9 1 9 1 9 1 12 9 2
25 1 11 13 9 2 9 2 16 4 15 11 13 1 0 12 12 0 9 2 4 3 13 0 9 2
16 3 4 9 1 9 13 10 9 9 9 2 7 14 13 0 2
30 9 9 15 3 13 1 0 9 2 1 15 4 9 2 16 4 1 10 9 13 9 1 12 9 9 2 13 10 11 2
45 1 9 4 15 1 0 9 13 2 16 4 11 2 16 4 13 12 9 9 2 13 12 9 0 9 2 11 2 16 1 10 9 4 13 2 7 4 1 12 9 9 13 1 9 2
31 9 11 8 11 11 4 3 2 16 4 13 1 11 2 0 9 13 2 16 13 11 11 1 9 14 1 9 0 12 9 2
2 8 8
14 2 0 9 13 12 9 7 13 0 9 7 12 9 2
2 11 2
9 2 1 9 15 15 13 0 9 2
11 15 15 14 4 13 2 16 13 1 9 2
9 13 15 15 2 16 15 15 13 2
11 15 14 13 0 2 7 15 9 13 3 2
9 13 9 2 16 15 13 2 2 2
15 13 15 2 10 9 13 1 9 7 15 4 1 15 13 2
6 13 10 9 2 2 2
12 14 15 1 9 13 0 9 2 3 15 13 2
19 7 14 16 14 13 2 15 13 2 16 16 13 2 7 3 13 10 9 2
12 3 15 4 13 2 16 1 9 13 10 9 2
13 0 9 9 4 13 9 14 3 1 9 2 2 2
20 0 0 9 1 9 11 4 13 0 16 9 2 16 4 1 9 13 1 11 2
19 9 15 4 1 9 13 7 13 4 13 0 15 2 7 4 13 1 9 2
22 16 15 4 13 13 1 9 2 16 4 15 13 2 15 4 13 13 2 16 13 9 2
13 11 4 10 9 13 1 9 1 0 0 9 11 12
10 13 7 15 4 2 16 13 11 0 2
13 13 4 11 7 13 2 16 13 0 1 9 9 2
19 11 2 16 4 13 3 10 9 2 4 13 1 11 1 9 13 1 9 2
19 11 4 13 2 10 13 10 9 2 7 15 4 13 1 9 11 1 11 2
30 16 4 13 11 2 3 0 2 15 4 1 0 9 0 9 13 13 12 9 1 0 9 2 16 4 13 14 0 9 2
22 11 2 16 15 4 3 13 2 4 3 13 2 16 4 13 11 2 3 13 1 9 2
31 14 16 15 4 9 11 13 2 16 4 11 13 2 16 15 13 1 9 14 14 9 2 15 4 11 13 2 16 15 13 2
20 1 0 2 0 11 1 0 9 4 13 0 11 1 0 9 13 14 3 0 2
18 7 7 4 11 11 13 2 16 15 4 1 9 1 9 13 0 9 2
10 1 3 0 9 4 13 9 1 9 2
12 9 4 13 9 1 9 7 15 13 1 9 2
49 10 9 4 13 9 9 1 9 2 2 16 4 3 13 10 0 7 0 9 2 16 15 4 13 3 2 7 13 4 15 15 3 2 16 4 13 0 7 3 0 2 16 4 15 15 3 13 2 2
16 1 10 0 9 15 4 11 13 2 16 4 13 9 1 9 2
31 1 10 9 4 13 2 16 13 0 9 0 9 9 2 9 2 9 0 9 2 9 2 9 2 9 2 9 7 0 9 2
8 9 1 11 4 13 10 9 2
24 9 12 4 13 2 16 13 9 1 9 14 15 3 0 2 16 1 15 15 14 14 13 9 2
47 11 12 4 2 16 4 13 0 9 2 13 10 16 12 9 9 11 11 2 16 4 13 9 9 2 16 4 15 13 16 2 3 0 9 2 16 15 4 3 13 0 9 7 0 9 2 2
19 7 11 4 13 10 9 3 2 11 4 3 13 7 15 13 1 0 9 2
14 1 15 4 13 12 9 2 16 4 13 1 10 9 2
16 13 4 2 16 4 13 9 7 15 4 1 9 13 0 9 2
17 16 4 9 13 10 0 9 2 4 13 0 1 12 9 0 9 2
23 9 13 7 13 0 1 9 0 9 2 9 0 9 13 9 10 9 2 16 13 0 9 2
27 7 4 9 11 13 10 9 2 16 2 4 1 0 9 14 3 13 10 9 9 2 16 4 15 13 2 2
7 3 15 4 13 10 9 2
11 3 1 9 4 14 13 2 15 4 13 2
12 7 15 4 10 0 9 3 13 1 9 11 2
15 14 9 11 0 3 4 13 9 2 16 13 1 0 9 2
41 11 11 2 0 9 9 2 4 9 11 13 2 2 1 9 2 16 15 13 1 9 2 15 13 1 9 2 1 0 7 0 9 2 16 13 2 16 13 0 9 2
7 9 15 13 1 0 9 2
13 9 3 13 9 2 9 9 7 15 13 1 15 2
18 7 15 15 14 13 3 13 7 15 3 13 2 7 0 13 1 15 2
9 1 10 9 13 3 16 10 9 2
15 13 4 13 2 7 11 15 4 13 2 16 13 1 9 2
8 13 4 7 13 9 1 9 2
29 13 2 16 10 9 14 3 15 3 13 3 14 4 13 0 7 16 4 9 11 13 0 14 9 2 16 4 13 2
4 13 9 11 2
7 2 3 15 4 9 13 2
27 9 2 16 4 13 9 1 0 9 2 4 13 9 11 2 13 9 2 16 15 13 1 10 9 16 11 2
5 14 2 4 13 2
11 16 14 13 2 16 13 9 2 7 13 2
7 14 13 15 2 4 13 2
2 13 2
14 15 13 14 9 2 1 15 15 4 13 10 0 9 2
7 15 4 15 13 1 15 2
11 16 15 4 9 13 2 4 13 1 15 2
11 13 4 10 9 7 13 10 9 1 15 2
20 1 15 4 10 9 2 16 4 14 13 9 2 13 1 9 7 15 15 13 2
25 10 9 0 9 4 13 1 15 7 1 15 2 7 15 4 13 13 2 16 4 13 0 1 9 2
14 16 15 4 13 2 15 4 3 7 14 3 13 3 2
21 3 4 15 3 13 10 9 1 9 9 7 13 1 15 9 2 0 1 0 9 2
22 3 13 0 2 16 13 1 10 9 2 16 13 10 9 2 15 2 16 13 1 9 2
6 7 3 13 1 9 2
15 14 16 4 15 13 2 15 14 13 3 3 13 1 9 2
14 15 4 13 15 2 16 4 13 2 7 4 15 13 2
7 13 15 4 3 16 0 2
11 9 11 4 13 10 9 7 15 15 13 2
11 3 14 4 13 2 16 4 13 10 9 2
18 9 11 2 11 2 11 7 11 4 1 9 13 2 16 15 13 9 2
14 16 4 13 10 9 2 15 4 1 9 13 0 9 2
12 3 4 13 2 16 4 13 9 1 11 11 2
29 0 9 11 15 1 0 12 9 2 1 0 9 9 9 2 1 15 4 1 0 9 13 0 9 2 4 3 13 2
27 1 9 4 0 9 11 11 11 2 11 2 13 9 13 1 9 10 9 2 16 4 3 13 9 9 9 2
34 16 4 13 9 1 0 9 2 4 15 7 13 2 16 9 1 11 2 11 2 11 1 11 7 0 0 9 9 14 4 13 14 13 2
37 1 11 4 13 14 1 9 2 16 4 13 13 0 9 14 9 3 0 9 1 9 2 3 16 4 13 1 10 9 1 9 9 11 13 0 9 2
16 1 11 4 9 1 0 9 1 0 13 14 0 12 0 9 2
13 11 11 2 9 2 9 4 1 0 13 3 3 2
19 13 4 2 16 4 3 3 13 1 9 7 15 4 3 13 9 7 9 2
8 3 4 13 14 13 1 11 2
12 9 13 3 0 2 7 0 9 3 14 13 2
23 11 13 16 0 9 3 0 7 13 3 9 2 16 15 14 4 1 15 13 1 0 9 2
26 3 13 14 3 0 9 11 14 0 2 7 15 15 9 1 0 9 1 9 1 11 3 3 3 13 2
21 11 14 13 13 2 16 4 1 9 13 2 16 13 1 0 7 3 3 0 9 2
20 14 15 15 4 14 13 2 16 15 4 11 3 13 1 10 9 1 0 9 2
3 2 8 2
50 1 9 0 9 4 13 3 0 13 1 9 9 2 1 0 9 2 1 10 0 0 9 2 16 15 4 13 0 9 2 0 9 2 9 2 9 0 9 2 14 1 0 15 9 4 15 13 15 13 2
27 1 10 10 9 7 9 10 0 9 1 9 1 0 9 13 1 9 13 2 16 15 4 13 3 15 15 2
27 9 12 4 1 9 9 2 16 9 9 13 2 10 0 0 9 13 0 0 9 2 15 13 14 0 9 2
11 9 1 11 13 1 12 1 12 9 9 9
8 9 1 9 13 12 1 11 2
10 0 9 7 9 0 9 13 1 11 2
9 9 12 15 1 9 13 1 11 2
7 3 13 9 2 11 2 2
27 1 9 12 2 12 13 1 9 1 0 9 1 11 1 8 11 11 2 9 2 7 11 11 2 9 2 2
6 13 7 13 1 11 2
7 9 12 13 9 0 9 2
22 13 4 1 12 0 7 0 9 0 9 1 9 2 1 0 0 9 7 0 0 9 2
37 3 4 13 1 9 2 16 15 4 11 13 9 12 2 16 4 13 0 9 1 9 12 1 12 2 3 4 13 9 10 9 1 9 12 1 12 2
10 1 9 9 4 13 0 9 12 9 2
39 13 15 1 0 0 9 11 11 11 2 13 14 4 9 0 9 12 9 2 16 13 1 9 1 10 9 2 16 4 1 10 9 10 9 13 1 0 9 2
17 2 3 13 1 9 9 2 9 2 9 7 9 2 1 0 9 2
4 9 0 9 2
14 13 15 0 0 0 9 0 9 7 1 0 0 9 2
11 14 1 0 9 15 15 9 14 4 13 2
4 13 0 9 2
25 1 9 1 9 9 15 4 0 9 13 2 16 4 3 13 1 0 9 1 9 1 9 0 9 2
21 9 13 1 9 0 9 9 7 0 9 2 16 15 4 13 9 1 9 0 9 2
52 0 0 9 0 9 13 0 9 1 9 1 9 9 2 0 9 9 1 0 9 2 9 0 9 0 9 1 0 7 0 9 2 1 0 9 7 14 13 1 9 9 0 9 9 0 9 1 0 7 0 9 2
10 1 0 9 13 10 0 7 0 9 2
13 3 13 0 2 9 2 3 9 4 13 10 11 2
8 1 9 4 13 14 9 9 2
10 3 15 13 2 16 15 14 13 14 2
9 1 9 9 13 14 10 0 9 2
23 12 1 9 13 0 9 2 16 13 1 9 1 11 2 3 13 3 14 0 9 1 9 2
12 1 11 11 4 1 9 13 0 0 0 9 2
11 13 4 12 9 7 12 9 1 12 9 2
20 1 9 4 13 0 9 7 9 0 11 2 16 4 13 3 12 9 0 9 2
3 2 8 2
36 0 9 11 11 4 1 9 13 0 9 2 1 15 4 0 9 0 0 9 1 11 1 9 9 12 2 12 2 12 9 2 13 12 9 9 2
25 9 4 14 13 1 10 9 2 1 15 13 0 9 9 2 7 13 0 9 9 1 0 9 0 2
8 0 9 4 13 1 9 0 2
10 0 9 7 4 13 13 10 0 9 2
24 1 9 15 4 1 9 13 14 9 0 0 9 11 11 2 16 4 9 1 11 13 1 9 2
9 0 9 1 11 4 13 3 0 2
25 1 9 4 13 14 0 9 7 14 0 0 9 4 13 13 9 2 16 13 13 0 0 9 0 2
11 2 1 9 1 0 9 3 13 3 0 2
45 0 13 13 14 0 7 13 2 16 4 1 15 14 0 13 0 9 2 2 13 11 2 16 15 4 0 9 13 1 9 2 16 4 11 1 9 9 11 11 13 9 1 0 9 2
14 11 3 13 0 9 9 2 0 9 11 7 13 9 9
20 16 9 1 0 9 14 13 1 0 9 2 15 13 1 9 9 9 7 9 2
8 3 13 10 9 1 0 9 2
21 9 3 13 13 0 9 2 16 13 13 0 9 2 7 7 0 1 0 9 13 2
28 2 4 1 11 14 1 0 12 2 0 0 9 1 9 12 0 9 0 9 13 1 0 12 1 12 12 9 2
25 1 10 16 12 2 0 9 2 15 4 13 3 7 1 0 12 9 3 2 4 13 14 3 0 2
24 2 16 4 13 13 0 9 2 13 1 3 3 13 0 9 7 13 0 9 2 2 13 11 2
82 1 10 9 1 9 2 3 15 4 0 9 13 1 0 9 3 7 3 2 4 1 0 9 0 9 13 9 2 16 4 13 1 0 9 0 9 7 9 1 11 11 2 16 4 15 9 0 9 13 1 11 12 9 12 7 16 15 4 3 13 1 2 9 9 7 9 2 7 1 0 9 2 0 9 1 9 2 9 2 9 2 2
46 13 15 3 2 16 4 0 9 13 14 9 1 11 11 2 16 13 2 9 9 2 9 7 9 0 9 1 9 9 2 7 13 9 7 9 1 9 10 9 13 9 10 0 9 2 2
11 3 13 1 11 0 9 1 9 0 9 2
32 1 9 0 9 7 9 13 3 13 1 9 1 11 2 1 15 7 13 0 7 0 3 7 3 13 14 1 15 1 0 9 2
22 16 4 13 14 10 9 2 4 1 0 0 13 10 0 9 9 1 3 12 0 9 2
15 10 9 13 3 3 14 3 13 0 9 2 13 1 11 2
36 16 4 9 13 2 16 13 3 3 2 13 9 3 0 11 2 8 8 8 2 2 16 13 10 9 9 2 16 9 13 2 16 9 3 13 2
31 16 13 9 2 0 2 1 0 2 0 9 0 9 16 10 9 2 13 1 9 1 9 3 12 9 2 9 9 12 2 2
18 1 9 1 12 9 4 13 11 11 2 11 11 2 2 0 9 12 2
20 9 1 9 4 13 1 0 9 1 0 9 9 2 11 11 11 2 9 12 2
19 0 4 1 0 9 14 3 13 0 9 7 15 1 9 13 0 9 3 2
28 11 11 2 11 11 2 4 3 1 0 9 13 3 2 7 1 9 4 13 3 7 3 13 1 11 11 11 2
13 1 9 9 7 9 1 12 9 11 4 13 9 2
9 13 4 10 9 2 9 7 9 2
20 1 10 9 4 3 14 13 2 9 15 13 2 16 15 4 9 13 1 9 2
28 0 9 1 15 13 9 11 2 16 1 9 12 0 0 9 13 3 3 14 3 12 0 9 1 10 9 9 2
15 9 4 1 0 0 9 13 13 14 9 0 0 9 11 2
9 10 9 7 15 14 13 15 0 2
36 3 15 1 10 9 2 16 4 15 1 11 3 13 1 0 0 9 2 11 3 3 13 0 0 9 2 2 13 14 9 1 0 9 0 11 2
12 1 0 11 4 13 10 9 3 0 0 9 2
44 9 4 0 9 1 9 11 11 13 1 0 9 2 1 15 4 13 2 16 4 1 9 12 7 12 1 9 9 1 0 9 14 12 9 13 9 7 15 13 9 7 0 9 2
6 1 9 13 3 9 2
36 0 4 15 14 0 9 13 0 9 2 7 4 10 0 9 1 10 9 13 9 1 0 0 9 7 13 1 9 1 15 2 15 15 4 13 2
36 3 7 15 13 2 3 15 2 16 14 13 3 3 2 15 2 16 14 13 3 3 2 13 2 3 4 1 11 0 9 1 9 13 0 9 2
24 16 4 14 13 1 0 3 1 0 2 4 13 0 9 0 9 2 16 13 0 9 0 9 2
3 10 9 2
8 14 10 9 15 4 3 13 2
11 9 13 14 0 2 16 13 9 0 9 2
13 3 13 11 14 3 16 12 2 0 9 11 11 2
19 11 4 13 0 0 9 9 11 11 2 13 7 4 14 10 9 11 11 2
8 0 9 3 13 1 0 9 2
17 1 0 9 13 7 0 0 9 2 16 4 15 13 1 8 9 2
8 14 3 4 3 13 1 15 2
17 3 2 16 13 1 9 2 15 3 13 7 15 13 10 0 9 2
34 13 15 1 0 9 7 15 15 3 2 1 9 2 1 9 0 9 2 16 13 1 9 9 7 1 0 9 1 9 2 13 0 9 2
5 7 3 13 0 2
15 13 15 3 7 13 9 2 16 4 13 9 9 1 9 2
13 2 3 13 2 16 4 10 9 13 0 9 9 2
5 3 14 13 9 2
9 13 9 9 7 9 1 10 9 2
4 2 13 9 2
22 13 9 10 9 2 13 15 2 3 7 3 4 15 13 2 16 4 13 3 1 9 2
12 14 3 15 13 13 0 9 0 9 1 9 2
12 0 9 14 4 13 0 9 7 13 0 9 2
34 10 9 13 1 0 9 2 0 0 9 2 1 9 9 2 2 9 2 3 0 0 9 2 0 9 2 9 2 0 9 7 0 9 2
17 2 13 9 1 9 2 1 9 7 9 2 15 13 3 3 13 2
14 14 13 9 2 16 7 15 7 13 2 15 9 13 2
11 13 9 1 9 2 16 4 15 13 3 2
13 2 16 13 0 9 2 15 3 3 13 7 13 2
15 2 13 0 2 3 4 9 13 2 7 15 13 9 9 2
18 2 13 2 16 4 13 1 9 7 14 10 9 1 15 9 3 0 2
6 1 9 15 3 13 2
32 16 15 13 9 2 13 2 16 15 9 14 13 1 9 2 7 1 10 9 13 9 9 2 0 1 9 2 16 15 3 13 2
9 14 13 2 16 15 9 14 13 2
19 2 13 9 2 9 7 9 1 9 7 9 2 16 4 13 7 13 9 2
43 7 0 9 0 9 11 11 4 13 2 16 4 9 13 10 9 1 9 1 0 9 2 16 4 15 13 2 14 3 1 15 2 3 4 9 13 14 14 9 9 7 3 2
12 9 4 13 3 12 3 0 9 1 0 9 2
8 15 7 15 9 14 13 0 2
11 14 4 13 9 13 1 9 9 7 9 2
8 9 9 15 13 0 0 9 2
19 7 1 11 4 11 1 0 9 13 2 1 11 7 14 14 4 13 9 2
24 1 9 0 0 9 13 3 9 2 3 4 11 7 13 9 1 9 1 11 1 9 1 11 2
24 16 7 0 9 1 15 14 4 13 13 1 11 2 4 0 9 14 13 1 9 1 0 9 2
50 1 0 9 2 1 15 13 1 11 1 0 9 14 4 11 11 13 9 1 0 9 1 0 9 14 13 15 13 7 13 2 16 15 15 9 9 1 11 14 3 14 13 14 7 4 15 13 0 9 2
26 14 7 13 11 7 11 14 0 0 0 9 2 16 15 4 11 13 1 9 2 16 15 4 9 13 2
3 2 8 2
14 3 4 13 10 9 1 12 9 3 14 0 12 9 2
14 1 0 9 4 13 2 16 13 9 3 3 0 9 2
27 3 13 10 9 0 9 2 7 9 2 4 1 9 11 13 13 0 9 2 1 15 4 9 7 9 13 2
28 11 11 2 3 2 4 13 9 2 11 11 7 4 13 1 9 2 16 4 13 9 1 0 9 0 1 9 2
18 3 15 13 2 16 9 1 0 9 13 14 9 7 12 9 1 9 2
21 1 15 14 13 0 0 9 2 0 9 2 10 9 7 9 9 2 16 15 13 2
23 9 1 9 0 9 9 13 14 15 2 9 1 9 13 0 1 9 2 16 13 10 9 2
23 9 1 15 3 13 9 2 9 2 0 9 7 13 12 1 9 2 16 13 9 1 9 2
8 1 9 13 3 0 0 9 2
31 1 0 0 9 10 9 4 0 9 11 11 13 9 9 7 10 9 2 11 2 2 16 13 10 9 14 1 9 1 9 2
29 1 9 7 0 9 1 9 2 16 15 1 10 9 14 13 2 4 15 13 2 16 15 13 14 9 9 1 9 2
15 0 9 13 3 0 1 9 2 0 13 3 7 3 0 2
28 13 4 15 0 9 2 9 1 9 2 16 4 13 1 0 9 2 3 3 0 13 9 2 16 13 1 9 2
17 1 9 7 4 13 0 9 1 9 2 7 4 1 15 13 9 2
10 9 9 11 13 1 9 1 0 9 2
13 9 11 13 1 9 1 12 0 0 9 1 11 2
5 15 0 8 9 2
17 4 15 15 7 13 2 16 13 1 11 0 7 11 3 10 9 2
25 13 15 4 1 11 2 16 15 4 14 3 13 1 11 0 7 15 13 2 16 16 15 14 13 2
6 14 10 9 4 13 2
9 2 13 3 2 2 4 13 11 2
10 2 1 0 9 4 13 0 10 9 2
23 11 4 13 9 7 13 9 1 12 9 2 16 4 13 9 2 3 13 1 10 9 0 2
11 0 9 4 13 1 9 1 0 0 9 2
8 3 9 10 9 4 13 0 2
12 7 4 1 9 9 13 10 9 1 0 9 2
16 0 9 1 9 9 11 4 13 15 2 16 4 3 15 13 2
24 7 16 4 14 3 13 13 2 7 3 7 3 4 13 9 2 16 4 4 3 13 0 15 2
8 9 11 11 4 13 10 9 2
7 1 9 4 15 13 9 2
4 13 4 9 2
5 13 4 0 3 2
26 16 15 4 13 9 11 11 2 4 15 9 13 2 3 4 0 13 9 1 9 7 15 13 1 15 2
5 13 7 4 0 2
8 14 15 4 13 1 9 9 2
12 16 4 13 1 9 2 4 13 9 1 11 2
19 13 4 9 2 16 15 4 11 11 13 1 10 9 2 16 4 13 15 2
7 3 15 4 13 1 9 2
15 7 4 13 7 15 13 2 16 4 13 9 0 0 9 2
6 7 11 4 13 9 2
14 14 3 9 15 4 3 13 0 2 0 9 11 11 2
9 10 9 4 3 13 9 0 9 2
22 7 16 15 4 2 16 4 13 2 13 9 9 7 9 4 15 13 1 9 16 9 2
38 16 4 11 13 1 9 1 9 2 15 15 4 13 2 16 4 3 13 2 3 4 13 3 9 2 1 0 9 2 1 15 4 13 9 1 10 9 2
14 1 9 4 13 2 3 9 13 7 13 1 0 9 2
11 9 4 13 7 3 0 1 9 7 9 2
27 13 4 0 9 2 16 4 15 4 3 13 2 16 4 13 0 2 7 4 13 10 9 3 0 16 9 2
22 2 7 15 14 4 13 1 9 9 2 16 4 13 1 9 2 2 4 13 11 11 2
12 13 4 9 2 16 4 13 15 0 7 0 2
11 9 4 13 14 3 2 16 16 15 13 2
17 3 16 4 9 13 1 9 2 4 13 15 2 16 4 13 9 2
13 13 4 0 1 0 9 2 16 4 13 0 9 2
28 1 10 9 4 15 3 13 1 10 9 2 1 0 9 7 9 2 16 14 4 15 13 2 3 15 13 9 2
24 11 4 13 3 14 3 0 2 3 0 2 16 7 4 15 14 3 13 2 16 4 15 13 2
11 11 15 4 13 2 16 4 13 9 9 2
6 10 9 4 13 3 2
6 13 15 4 1 9 2
11 13 4 0 9 1 0 9 2 16 9 2
12 13 7 4 9 14 0 9 9 1 0 9 2
8 16 13 15 3 2 14 13 2
5 9 13 9 9 2
15 2 13 2 16 14 4 13 14 3 2 2 4 3 13 2
33 0 9 2 9 11 11 2 16 15 4 13 0 9 2 13 3 2 16 13 2 1 9 9 2 16 15 13 13 1 9 1 9 2
17 0 9 15 4 13 13 9 2 16 15 15 4 13 16 0 9 2
32 9 2 16 4 15 9 13 14 0 9 2 1 3 14 13 0 2 7 0 9 4 13 2 16 4 13 9 1 0 0 9 2
10 9 0 9 4 3 13 10 10 9 2
9 11 4 13 3 2 15 4 13 2
25 1 10 9 4 1 10 9 3 13 11 11 2 0 9 0 9 2 14 16 4 13 13 0 9 2
8 3 7 13 0 9 0 9 2
34 3 4 0 0 9 13 11 1 9 7 13 2 16 4 1 9 2 1 15 4 13 0 2 2 13 2 1 12 9 9 10 0 9 2
19 0 9 1 9 0 0 0 9 4 14 13 2 9 15 4 13 1 0 9
14 1 9 3 4 1 9 0 9 3 13 0 0 0 9
11 9 0 9 11 12 13 1 9 0 9 2
14 9 4 13 12 9 2 16 4 13 9 7 0 9 2
24 9 4 15 13 1 9 0 9 9 2 9 1 9 12 9 2 16 4 13 11 7 11 11 2
17 3 4 13 15 0 9 1 9 2 7 4 9 13 1 12 9 2
28 0 9 11 12 4 13 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 7 11 2
9 9 4 1 9 13 14 12 9 2
8 1 9 9 4 13 0 9 2
18 2 9 2 16 15 4 1 10 9 13 9 2 13 0 9 9 9 2
12 13 15 9 2 9 7 9 9 9 1 9 2
18 16 4 1 9 13 2 4 13 9 13 10 0 9 1 0 0 9 2
19 0 13 2 16 4 14 15 13 7 13 2 14 4 13 13 10 0 9 2
25 1 0 2 16 13 10 12 9 2 13 2 16 15 4 0 0 9 1 10 0 9 13 3 3 2
19 1 10 9 4 3 13 1 0 9 2 16 4 13 9 0 9 1 11 2
29 9 13 0 1 9 2 16 15 13 2 7 13 14 0 9 1 9 7 9 2 16 15 9 14 4 13 7 13 2
37 10 9 1 11 2 16 3 13 1 9 0 9 2 4 14 3 13 9 2 16 4 13 10 9 2 1 15 14 1 3 14 4 13 13 0 9 2
12 13 15 9 12 2 9 13 0 1 0 11 2
2 13 2
7 0 9 0 9 15 13 2
11 11 11 1 9 0 11 3 13 1 9 2
17 1 9 4 13 2 16 4 15 13 1 9 2 16 15 4 13 2
26 1 9 15 13 0 9 11 11 2 16 14 13 2 16 15 15 4 10 0 9 1 0 13 1 9 2
30 1 15 4 13 11 7 10 0 9 2 0 9 11 2 16 15 13 13 9 2 1 15 4 11 13 1 9 2 2 2
14 0 9 0 9 13 11 11 2 11 11 7 11 11 2
10 0 9 0 9 11 11 7 11 11 2
11 1 0 9 9 1 0 9 4 13 11 2
21 9 2 3 15 4 0 13 2 13 0 7 13 9 0 9 0 9 2 4 13 2
9 9 3 13 1 12 1 12 9 2
12 10 9 13 3 9 9 2 16 15 14 13 2
9 1 10 9 3 14 13 0 9 2
22 9 3 13 14 9 1 9 9 2 14 10 9 13 3 3 0 2 16 13 15 0 2
10 3 4 13 3 2 16 15 13 0 2
22 0 11 13 9 2 16 15 14 1 3 4 13 11 7 4 13 10 0 9 0 9 2
30 3 13 10 9 2 7 14 15 13 1 9 0 11 2 16 15 13 1 0 9 1 0 9 7 1 3 13 9 3 2
27 1 9 15 4 13 10 16 12 0 9 7 7 3 0 9 9 9 2 1 9 15 13 14 14 3 12 2
26 1 3 12 3 2 1 12 0 9 7 1 9 4 13 0 9 2 16 4 15 3 13 3 1 3 2
19 15 0 7 0 2 0 7 0 9 4 13 1 9 1 9 3 0 9 2
18 4 15 13 14 9 0 9 2 7 10 10 9 9 2 9 7 9 2
14 0 12 9 1 9 13 16 3 0 1 10 10 9 2
29 3 1 9 2 16 4 15 0 13 1 10 9 2 4 13 7 13 9 2 16 15 4 10 10 9 13 1 9 2
30 9 7 9 2 16 13 9 11 2 4 1 9 11 2 0 9 11 2 16 4 13 1 9 0 9 2 13 11 11 2
25 3 4 13 9 0 9 3 1 9 2 7 1 10 14 12 9 1 15 4 13 0 9 7 9 2
5 14 9 4 13 2
27 9 15 4 1 15 15 13 2 3 7 13 9 2 16 15 4 13 1 9 0 9 2 9 0 0 9 2
27 1 12 9 2 16 14 4 15 1 9 13 9 11 2 1 9 1 0 9 13 9 2 16 3 13 9 2
7 16 9 15 13 3 3 2
11 3 1 9 15 13 1 10 9 3 13 2
19 1 15 15 13 1 9 2 10 12 9 13 1 9 9 7 13 15 0 2
17 1 9 2 16 13 0 0 9 2 0 9 1 9 2 13 9 2
19 15 4 13 10 9 1 9 2 3 13 0 3 2 16 13 1 15 9 2
12 0 9 7 4 13 1 10 9 14 9 3 2
11 1 9 1 0 9 13 7 0 7 0 2
31 10 9 13 0 9 16 9 0 9 7 16 12 1 9 9 2 16 15 13 3 0 1 9 7 9 9 2 1 15 13 2
36 0 9 1 15 2 7 14 12 0 9 1 0 9 7 13 2 16 3 9 1 0 13 1 9 10 14 9 2 16 13 3 1 9 10 9 2
17 3 3 1 10 9 13 1 9 0 2 0 2 0 7 0 9 2
22 1 0 9 9 0 9 15 1 15 13 14 9 7 9 2 16 13 1 3 0 9 2
17 16 13 0 9 0 7 0 2 14 14 13 2 16 13 3 0 2
13 16 7 15 15 3 13 2 4 13 13 10 9 2
13 3 14 13 9 1 0 9 16 4 15 13 9 2
10 15 13 14 14 0 2 7 14 0 2
29 7 13 1 11 10 0 9 2 7 14 1 9 13 3 13 10 9 2 16 14 4 13 3 2 16 15 4 13 2
22 3 7 4 3 13 2 16 14 13 13 2 16 13 9 7 13 0 13 10 0 9 2
26 15 13 14 3 0 2 7 1 9 9 3 3 13 1 9 7 15 13 0 9 1 9 1 0 9 2
12 11 4 0 3 0 9 13 1 0 7 0 2
13 7 13 9 1 9 10 9 7 15 1 15 13 2
21 9 1 15 13 0 9 1 0 9 2 9 7 0 9 2 16 15 13 10 9 2
34 0 0 9 11 11 4 1 0 9 9 9 9 9 13 1 9 2 16 13 3 13 16 13 2 7 9 13 3 3 13 16 7 13 2
13 3 13 11 12 9 1 9 1 11 3 0 9 2
12 3 9 13 3 1 9 7 15 13 1 9 9
17 1 15 4 13 1 0 9 2 7 14 3 1 15 9 13 9 2
6 2 9 15 13 9 2
10 13 4 3 3 7 0 13 13 11 2
13 0 13 2 16 14 4 13 2 2 13 11 11 2
14 10 9 2 15 15 13 9 7 9 2 13 11 11 2
19 9 11 4 13 1 9 3 9 1 9 2 3 7 13 12 9 10 9 2
7 2 15 13 15 0 9 2
11 13 4 1 10 9 7 15 3 14 13 2
15 0 9 13 15 0 7 10 9 3 13 2 16 15 13 2
25 11 13 0 9 2 7 3 1 10 9 1 9 7 0 9 1 9 13 1 15 0 14 10 9 2
35 16 4 13 3 16 13 2 4 9 13 0 1 15 2 2 13 12 2 0 11 11 2 16 15 0 1 10 9 1 9 13 9 1 9 2
8 15 4 1 15 13 0 9 2
12 12 4 13 1 9 7 15 13 9 1 9 2
35 9 4 0 9 13 1 9 7 15 13 13 9 2 1 9 7 15 4 8 8 1 9 9 13 1 9 7 13 1 0 9 9 7 9 2
30 1 11 11 4 1 12 1 12 9 1 9 0 9 11 13 9 11 11 11 2 1 15 15 4 13 12 9 9 11 2
24 9 9 11 11 2 16 4 1 0 12 9 9 13 3 3 2 4 13 0 0 7 0 9 2
19 15 14 4 3 13 9 9 14 1 9 0 9 1 3 1 9 7 9 2
19 2 9 2 16 4 15 9 9 8 11 11 13 1 9 2 13 10 9 2
17 13 2 16 13 9 9 0 9 7 16 13 1 0 9 0 9 2
33 1 9 9 9 0 0 9 1 0 9 13 14 14 10 9 2 7 14 9 11 11 1 15 2 16 4 13 11 13 0 9 11 2
33 2 16 13 10 9 2 13 0 2 16 4 10 9 2 16 4 13 9 2 13 13 10 9 7 13 0 9 2 2 4 13 11 2
23 9 9 13 14 1 0 9 0 9 7 9 9 2 0 9 13 0 7 0 2 0 9 2
39 9 14 4 3 10 9 13 7 13 1 1 15 0 0 9 2 1 9 2 1 15 13 0 14 0 9 2 7 13 14 13 0 2 3 0 13 0 9 2
25 9 2 16 1 0 9 7 9 0 0 9 13 1 9 10 9 2 1 10 9 13 3 12 9 2
28 16 4 3 14 1 10 9 2 10 9 15 13 1 0 0 9 2 13 0 9 2 15 4 13 14 12 9 2
2 3 2
23 1 11 7 13 9 2 16 4 13 0 9 2 9 13 14 0 11 2 16 13 0 9 2
29 3 13 0 0 9 13 0 0 9 2 16 10 9 3 13 2 0 9 7 13 13 3 12 9 1 9 10 9 2
30 3 15 3 13 2 16 13 9 14 0 2 16 9 14 13 3 10 10 9 2 7 4 14 9 3 3 13 0 9 2
32 9 11 11 4 1 9 12 13 0 0 9 11 2 1 15 4 9 3 16 9 13 9 11 1 11 2 11 2 11 7 11 2
36 0 9 13 0 16 9 8 8 0 9 2 16 0 0 9 13 9 0 9 7 9 1 9 2 16 1 0 9 13 7 13 9 1 0 9 2
39 0 13 2 16 4 15 1 0 9 13 15 2 16 13 0 2 0 9 2 16 13 9 2 9 2 9 7 9 2 7 3 3 13 9 2 9 7 9 2
31 9 9 11 11 13 0 9 11 11 2 9 2 2 11 11 2 9 2 2 11 11 2 9 2 7 11 11 2 9 2 2
20 1 9 0 9 0 13 13 0 4 13 3 12 9 1 11 2 11 2 11 2
22 11 11 2 12 1 9 9 0 9 11 2 13 2 16 13 0 9 9 0 0 0 9
14 0 9 13 2 16 15 13 2 15 4 13 10 9 2
12 3 14 4 14 13 13 1 9 12 9 3 2
6 13 2 15 15 13 2
29 9 4 13 9 9 2 16 13 1 0 0 9 0 1 9 1 9 2 1 9 7 2 15 13 2 14 10 9 2
47 13 0 13 2 16 4 1 10 0 9 9 2 16 14 13 9 1 10 0 9 2 13 15 10 9 2 16 4 15 10 9 9 2 16 1 9 14 4 13 0 2 13 14 10 0 9 2
23 7 13 15 2 14 13 2 16 1 0 9 0 9 14 13 3 0 9 9 7 0 9 2
29 9 0 9 1 0 7 0 9 13 14 9 0 9 1 9 2 7 1 0 0 0 9 16 1 9 1 0 9 2
18 15 4 13 14 0 9 1 0 2 0 9 2 0 9 1 10 9 2
4 4 15 13 2
24 4 13 9 2 16 4 13 3 1 9 1 9 7 4 3 13 2 15 15 13 2 15 13 2
17 3 7 13 14 9 2 16 15 9 13 7 15 14 13 0 13 2
11 16 13 15 3 0 2 13 0 7 0 2
1 2
11 9 1 0 9 13 2 16 13 3 0 2
23 14 3 3 13 0 1 9 0 9 12 7 12 9 2 16 13 0 9 9 0 1 11 2
34 3 7 13 10 9 0 9 3 0 1 10 9 2 16 13 0 9 1 0 1 9 1 0 2 7 3 3 13 13 1 12 1 0 2
17 9 1 9 1 9 4 1 1 0 13 9 2 16 4 15 13 2
15 9 9 4 13 1 0 9 2 16 4 13 1 0 9 2
14 3 3 4 13 10 0 9 2 16 4 13 9 9 2
7 3 7 15 4 15 13 2
23 3 13 0 9 0 9 2 1 15 4 11 11 7 11 8 13 9 1 9 1 0 9 2
22 3 15 11 11 2 11 11 7 11 11 13 0 9 1 2 0 9 2 7 0 9 2
17 1 10 9 13 9 3 3 13 16 9 9 9 1 9 7 9 2
19 1 10 9 4 13 0 2 16 4 13 9 14 3 0 3 13 7 13 2
21 13 4 13 2 16 9 2 16 13 2 13 2 16 13 0 9 2 9 7 9 2
8 9 13 0 7 3 13 9 2
11 16 13 9 0 2 3 13 12 0 9 2
12 0 13 13 7 9 16 9 2 16 13 9 2
19 9 0 9 13 9 9 2 16 4 1 12 9 13 0 9 7 0 11 2
10 7 9 16 9 4 13 1 0 9 2
23 0 9 0 13 2 3 4 15 3 13 9 2 16 13 14 10 9 1 9 10 0 9 2
34 16 13 10 10 9 1 9 2 0 9 0 9 2 10 9 1 15 2 15 13 1 9 2 13 9 1 9 0 9 0 1 10 9 2
18 9 13 13 10 10 9 7 13 9 1 0 2 0 2 0 2 0 2
8 11 11 10 9 13 9 9 2
14 13 15 4 0 9 2 1 15 13 9 16 0 9 2
48 12 9 13 1 11 11 9 0 0 9 2 9 0 9 1 0 9 2 15 13 9 2 16 9 13 0 1 15 7 3 9 7 9 2 16 13 1 9 2 3 13 7 1 0 9 13 9 2
8 9 7 14 13 7 15 13 2
15 9 13 3 0 1 9 2 16 7 13 7 7 13 9 2
8 13 1 10 9 1 0 9 2
25 12 9 2 16 13 1 11 1 10 9 0 9 2 13 3 14 9 1 9 2 1 9 7 9 2
17 1 0 7 0 9 4 15 9 13 14 1 15 2 16 13 9 2
33 16 4 15 2 16 4 13 11 1 0 9 14 3 13 2 16 13 9 0 1 9 2 7 9 7 9 1 0 13 7 13 9 2
26 0 9 9 1 0 11 13 1 2 0 9 2 7 1 9 16 9 2 16 15 13 9 7 10 9 2
19 3 14 13 9 1 15 4 13 2 16 4 13 1 9 14 1 0 9 2
32 1 0 9 14 13 0 0 9 7 1 9 13 14 2 9 2 0 9 2 16 13 15 14 1 12 9 7 15 13 16 9 9
24 11 2 1 9 0 9 0 9 4 3 13 9 1 12 9 11 11 2 9 2 9 7 9 2
34 9 1 9 2 16 13 1 0 0 9 1 9 0 9 1 0 9 2 4 13 1 9 10 9 2 9 7 4 13 9 0 9 11 2
3 2 8 2
47 1 0 0 9 11 1 11 4 0 9 9 13 7 13 9 2 16 15 4 3 13 13 1 9 12 9 2 7 15 4 13 3 12 9 1 9 2 15 3 13 9 9 1 9 7 9 2
9 1 0 9 15 9 4 3 13 2
24 0 9 1 9 4 13 1 12 2 0 9 0 9 2 7 4 15 9 13 14 3 12 9 2
23 14 7 15 4 3 13 2 7 4 14 0 9 9 0 9 13 14 15 10 9 1 3 2
22 9 1 12 1 12 9 13 1 11 14 0 2 0 9 7 14 13 1 0 12 9 2
27 13 15 4 9 2 1 10 0 9 4 15 3 0 9 13 1 9 2 7 15 15 3 0 14 13 13 2
32 9 2 16 4 13 0 1 9 2 4 13 0 2 16 15 4 9 9 1 9 9 13 14 12 9 1 9 1 0 0 9 2
17 9 9 1 9 1 0 9 4 13 1 9 1 0 9 3 0 2
22 14 7 14 4 13 1 9 9 1 0 9 1 9 9 1 9 3 0 3 12 9 2
28 9 14 14 13 3 13 14 1 9 9 7 9 2 9 7 14 4 0 9 13 0 9 3 1 9 12 9 2
33 14 7 14 4 14 1 9 11 13 3 0 9 1 9 12 1 12 9 2 7 14 13 9 2 16 4 15 9 2 3 13 2 2
27 16 4 13 0 9 1 9 1 9 11 11 2 1 9 1 9 0 9 3 13 1 12 1 12 9 9 2
13 1 9 9 7 14 12 9 10 9 13 0 13 2
26 2 1 0 13 1 9 9 14 9 1 9 2 1 10 0 9 7 15 13 12 9 9 1 0 9 2
27 1 15 13 3 0 2 16 16 13 0 9 2 16 4 13 0 9 2 3 0 9 13 9 9 1 9 2
25 9 0 14 13 9 2 1 15 13 0 9 13 9 9 2 13 7 14 13 2 16 9 14 13 2
7 0 9 14 3 15 13 2
11 1 9 15 13 11 8 8 7 9 9 2
17 11 11 8 13 2 16 1 0 9 13 0 14 9 2 7 14 9
13 2 0 13 2 16 0 9 12 9 4 13 9 2
25 16 15 4 13 11 11 2 7 4 13 0 9 11 11 1 10 9 1 0 9 13 3 12 9 2
24 16 13 9 2 13 2 16 15 15 14 13 13 2 7 16 0 9 13 10 0 7 0 9 2
20 2 1 0 11 9 1 0 9 4 13 2 14 0 4 15 3 13 1 11 2
6 1 11 15 14 13 2
10 1 11 3 4 13 10 0 0 9 2
11 11 4 13 9 0 9 1 11 7 9 2
4 2 14 13 2
6 11 15 14 4 13 2
7 3 13 2 15 13 9 2
5 15 4 13 9 2
5 3 15 4 13 2
35 9 4 13 2 3 13 1 9 1 11 2 15 15 13 7 3 13 9 12 14 3 15 2 16 14 4 11 13 0 9 1 0 0 9 2
13 13 2 16 13 15 0 0 9 7 0 0 9 2
10 3 13 9 9 1 9 10 0 9 2
10 13 2 16 13 15 0 9 0 9 2
32 10 9 13 1 10 9 0 1 15 0 2 10 0 9 2 9 9 0 9 2 16 13 1 15 7 1 15 1 10 9 13 2
12 0 13 2 16 4 0 0 9 13 0 9 2
24 9 14 13 14 3 9 2 1 15 15 9 1 10 9 13 2 16 13 7 13 9 0 9 2
14 1 9 13 9 1 9 1 0 9 1 9 12 2 12
18 13 1 9 11 1 11 2 11 1 9 9 7 0 11 1 0 9 2
29 9 9 1 0 9 7 13 1 9 0 9 0 11 7 11 1 11 2 11 1 11 7 0 9 1 11 1 11 2
11 1 0 9 0 0 9 1 9 0 0 9
7 0 9 7 13 0 9 2
26 11 8 13 10 12 0 9 1 10 9 2 16 15 13 0 9 2 7 13 15 0 9 1 0 9 2
17 9 11 4 1 10 9 1 11 13 14 12 0 9 1 0 9 2
20 9 13 0 13 1 12 7 12 0 9 7 13 0 7 1 9 16 0 9 2
22 0 13 14 12 2 0 9 12 1 12 9 1 0 9 7 0 9 2 12 9 2 2
2 14 2
16 3 0 4 13 2 16 4 1 9 1 9 13 15 0 13 2
21 3 7 13 2 16 15 4 15 3 13 9 9 0 0 9 1 9 1 9 9 2
31 13 2 16 4 1 0 12 9 0 9 2 16 15 4 15 3 13 2 13 1 10 16 12 9 9 0 9 1 0 9 2
11 3 4 15 1 0 0 9 9 3 13 2
27 1 9 9 4 13 3 14 3 10 16 12 9 0 9 7 4 15 14 1 10 9 13 1 3 9 9 2
9 1 0 9 13 3 9 11 0 2
25 0 7 1 15 14 0 9 13 3 9 7 9 7 9 0 9 2 16 13 9 2 9 7 0 2
21 0 0 9 13 1 9 2 16 13 3 0 2 7 1 0 9 1 3 0 9 2
34 9 13 0 3 2 16 9 1 9 9 7 9 13 1 0 9 14 9 0 9 7 14 9 1 9 0 9 7 9 7 9 10 9 2
21 13 9 2 16 13 0 9 0 9 7 9 2 15 4 13 9 13 16 10 9 2
12 15 15 13 15 0 2 0 9 9 7 9 2
7 10 9 13 15 1 9 2
7 10 0 9 13 0 9 2
17 3 13 2 16 4 15 13 10 1 9 7 16 4 15 3 13 2
6 15 13 9 15 0 2
22 13 1 0 9 7 13 15 15 3 2 16 13 15 10 9 2 7 15 13 10 9 2
9 13 9 7 14 13 1 0 9 2
24 1 11 13 15 12 3 0 9 2 16 13 0 9 9 2 15 4 13 3 13 1 9 9 2
23 11 2 0 9 11 2 16 15 13 1 9 7 9 0 9 2 3 14 13 1 9 9 2
47 1 9 7 0 15 0 9 1 0 9 15 4 9 11 13 1 9 0 9 9 0 9 2 16 4 1 9 13 1 9 0 9 11 7 10 9 9 11 2 16 4 14 3 13 1 9 2
22 9 0 9 0 9 4 11 13 1 11 9 11 2 16 15 15 4 13 1 9 9 2
25 3 9 13 1 9 0 9 2 1 0 9 7 14 4 15 0 13 1 0 7 1 9 0 9 2
3 2 8 2
11 3 3 15 10 9 4 14 13 14 13 2
12 11 13 3 0 2 3 7 13 0 1 0 9
25 1 9 11 15 3 13 1 9 1 12 7 12 9 2 16 13 14 0 7 0 0 9 0 9 2
17 1 0 9 4 3 1 0 9 13 9 0 0 9 1 3 3 2
18 9 15 3 1 0 9 4 3 13 2 15 13 0 9 1 12 9 2
17 1 10 9 15 13 14 0 9 2 16 7 4 13 0 0 9 2
18 16 13 9 9 1 9 9 2 3 13 2 16 9 3 13 9 9 2
22 16 9 14 13 3 0 1 12 9 2 3 13 9 9 1 9 1 12 7 12 9 2
16 16 7 15 9 3 13 1 12 9 2 3 13 14 0 9 2
21 9 0 9 15 3 13 3 12 0 9 2 1 0 9 7 4 13 9 12 9 2
18 3 1 0 9 9 3 13 2 16 4 9 14 3 13 1 12 9 2
20 1 3 0 9 7 15 4 9 9 3 13 1 12 9 2 16 9 13 3 2
16 15 4 3 13 1 9 2 16 4 9 13 1 14 12 9 2
15 1 9 0 9 13 3 10 0 9 2 16 4 13 9 2
21 9 1 0 9 9 1 0 9 4 1 0 9 0 9 9 0 13 1 0 9 2
3 2 8 2
8 1 3 15 4 13 14 9 2
22 13 4 1 9 9 2 7 4 15 3 13 2 16 4 13 2 16 15 4 13 0 2
12 2 14 15 15 14 13 2 2 4 3 13 2
5 2 13 10 9 2
9 2 13 4 1 11 7 1 9 2
31 1 9 4 15 13 0 2 7 0 9 2 1 9 9 14 14 13 9 2 16 15 4 13 0 1 9 7 4 13 0 2
40 0 7 0 9 2 12 9 7 12 9 2 11 11 11 4 7 13 0 9 11 11 1 12 9 9 2 15 13 3 3 3 2 16 4 0 9 13 1 9 2
12 9 1 0 0 9 7 4 13 0 0 9 2
24 11 4 13 9 1 9 14 3 1 0 9 2 1 9 7 4 13 10 10 0 9 7 9 2
39 1 10 0 9 4 11 3 12 13 14 10 9 1 9 0 9 8 8 8 8 8 8 8 8 8 2 16 4 13 14 12 1 9 1 0 9 1 11 2
19 13 0 9 10 9 7 13 0 9 1 9 0 9 1 0 0 0 9 2
19 10 9 4 14 3 3 13 9 1 9 0 9 1 9 1 0 0 9 2
13 0 9 9 1 9 13 9 2 16 13 10 9 2
19 9 1 9 13 13 0 3 2 14 16 4 13 9 15 13 2 7 3 2
16 0 13 13 14 1 9 0 9 7 14 12 1 0 0 9 2
19 2 13 0 9 1 9 7 16 13 15 0 14 1 9 0 9 0 9 2
9 8 8 8 8 8 2 8 8 2
34 0 9 4 13 9 11 2 9 13 7 15 13 2 16 4 1 9 13 0 9 1 12 9 1 11 2 16 13 3 1 9 9 12 2
39 0 2 0 9 1 9 2 16 13 9 9 2 9 7 9 2 13 12 9 12 1 9 0 9 9 1 11 2 16 15 13 9 12 1 0 9 1 11 2
9 15 15 13 0 7 15 0 9 2
27 7 4 3 0 9 9 9 13 0 9 3 1 0 9 1 11 2 16 4 13 0 9 7 0 9 9 2
18 9 1 9 13 3 0 0 9 2 3 0 1 0 9 7 0 9 2
38 7 0 13 14 1 9 1 0 9 2 9 2 2 3 16 15 4 0 9 2 0 9 2 1 9 13 1 0 0 9 2 16 14 13 9 7 9 2
10 1 0 9 15 15 14 13 0 9 2
6 13 15 4 9 0 2
8 3 4 13 9 1 0 9 2
20 14 4 15 15 13 0 13 2 16 15 4 15 13 1 9 13 1 9 9 2
9 10 9 13 0 9 14 1 0 2
10 13 15 2 16 4 13 10 0 9 2
14 13 15 4 1 9 2 16 4 13 0 9 10 9 2
18 9 13 0 9 2 16 15 1 0 9 9 3 13 1 0 9 9 2
10 13 4 1 10 9 7 3 13 0 2
13 13 15 4 2 16 4 1 11 13 1 0 11 2
25 1 9 12 15 4 1 11 13 1 9 9 11 2 7 15 14 3 0 9 1 15 0 4 13 2
19 0 9 1 11 1 11 4 13 1 0 9 2 1 0 9 7 1 9 2
22 13 4 1 0 9 2 3 16 4 9 1 0 9 1 10 9 13 2 15 4 13 2
9 1 15 11 0 9 4 3 13 2
32 0 9 2 16 14 4 15 9 13 3 2 4 2 16 13 14 0 2 1 0 13 14 2 15 7 3 4 13 1 0 9 2
20 9 14 13 14 0 2 3 13 3 1 9 7 9 13 1 12 9 1 9 2
16 11 13 2 16 9 14 3 13 9 9 1 0 7 0 9 2
18 9 1 9 7 9 4 2 16 13 9 0 2 13 3 16 0 9 2
14 9 4 13 0 9 2 1 15 14 4 13 0 9 2
7 2 9 13 1 9 9 2
24 9 13 1 9 7 13 2 16 4 9 3 13 2 2 13 0 9 1 9 7 0 9 11 2
24 2 0 2 9 4 14 3 13 0 12 9 9 0 9 2 3 7 13 9 14 14 9 0 2
16 11 13 2 16 13 3 13 1 0 0 9 7 9 0 9 2
8 13 2 15 13 0 9 8 2
15 14 2 15 4 15 3 13 14 1 9 1 10 0 9 2
11 16 4 13 3 13 14 2 4 13 3 2
12 3 15 4 7 11 13 2 16 3 14 13 2
17 3 7 15 4 10 9 13 2 16 1 0 9 13 3 0 9 2
15 15 13 3 2 16 3 14 3 13 1 3 7 3 13 2
12 14 2 14 1 11 4 13 10 9 10 9 2
8 9 1 10 9 13 3 0 2
14 3 1 9 9 13 15 3 3 16 1 9 0 9 2
6 1 3 9 3 13 2
16 16 13 9 0 2 13 10 9 12 2 3 0 16 1 11 2
9 0 0 9 7 14 13 14 9 2
17 1 9 11 1 0 9 1 11 0 9 13 12 2 0 9 9 2
9 1 11 4 9 13 9 1 9 2
15 1 11 0 9 13 9 2 16 4 15 1 9 13 9 2
13 0 9 2 16 15 13 0 9 2 13 9 9 2
22 1 11 2 15 13 0 14 15 2 16 13 2 7 16 4 13 9 14 1 0 9 2
16 3 16 0 9 14 0 9 13 9 2 16 13 3 0 15 2
9 12 9 3 13 7 13 10 9 2
8 15 13 3 0 2 0 9 2
20 3 7 13 1 10 9 14 0 9 2 16 15 13 9 7 14 3 10 9 2
10 9 13 3 3 2 11 4 3 13 2
14 9 13 9 7 13 9 2 13 7 14 9 7 9 2
21 9 0 1 15 13 7 9 7 9 2 12 7 0 13 14 1 9 1 0 9 2
24 15 13 3 1 9 7 1 9 9 2 16 15 13 9 1 10 0 9 2 0 9 7 9 2
9 1 9 3 13 2 0 9 2 2
24 13 4 14 2 16 13 9 1 0 9 3 0 2 15 1 0 9 4 3 13 14 9 15 2
19 1 11 13 10 9 14 3 0 14 1 9 2 16 13 3 0 7 0 2
13 3 7 13 14 2 16 10 9 4 13 1 9 2
20 11 15 4 13 2 13 15 4 13 7 14 4 13 1 10 0 9 3 0 2
21 11 7 15 4 13 13 9 2 11 2 7 15 13 10 9 2 16 13 10 9 2
12 9 1 9 7 14 4 13 3 2 0 2 2
28 0 9 0 9 15 14 13 1 9 7 0 9 2 9 4 14 3 13 7 13 9 7 4 13 14 0 9 2
16 2 3 13 9 0 9 2 16 3 13 10 0 9 10 9 2
29 13 14 2 15 4 13 2 15 13 2 16 4 3 2 16 4 13 15 1 9 2 13 15 3 0 9 1 9 2
24 1 9 2 16 13 1 9 0 9 2 15 4 3 13 9 9 2 4 9 3 13 1 9 2
31 9 1 10 9 13 9 11 2 16 1 9 0 9 14 13 9 0 9 11 11 7 13 0 9 1 0 9 0 0 9 2
31 1 0 0 9 2 1 3 0 9 7 0 9 7 9 0 9 2 2 4 0 0 9 13 0 0 9 0 1 12 9 2
30 10 0 9 4 1 0 9 1 9 13 11 2 16 4 1 0 9 13 9 1 12 9 7 1 15 3 13 9 9 2
16 0 9 9 4 13 9 9 9 1 0 9 1 0 0 9 2
19 14 0 9 9 11 11 13 0 1 0 2 15 4 13 9 0 9 9 2
27 0 0 9 4 3 13 9 9 1 9 2 16 13 0 1 0 9 7 13 15 3 0 1 0 9 9 2
11 14 2 14 15 13 0 1 0 9 9 2
18 13 15 2 16 4 13 1 9 9 1 9 0 1 10 9 0 9 2
13 1 15 4 13 0 9 14 1 0 9 7 9 2
18 9 0 9 1 0 9 13 9 0 9 9 1 0 9 1 0 9 2
29 13 2 16 4 1 10 3 0 0 9 14 12 7 12 9 1 9 1 9 13 9 2 16 13 9 0 0 9 2
16 13 7 2 16 4 9 11 1 0 9 10 9 13 0 9 2
14 9 4 3 13 1 9 7 0 13 1 12 0 9 2
15 1 15 4 13 1 9 2 16 7 4 13 1 0 9 2
25 13 4 0 2 16 14 4 13 13 9 2 3 4 13 9 2 16 15 13 9 1 12 0 9 2
6 9 1 9 7 9 2
22 1 0 9 13 0 9 0 7 0 9 2 9 2 9 7 9 7 9 1 0 9 2
15 9 13 9 9 7 9 2 9 0 9 7 9 10 9 2
8 9 1 9 13 9 1 9 2
11 9 13 10 16 0 9 2 9 7 9 2
5 9 13 9 9 2
1 9
17 13 0 0 7 13 0 0 2 16 15 13 15 3 13 1 15 2
11 16 4 9 13 15 2 3 14 15 13 2
16 14 13 9 1 9 2 16 4 13 9 1 0 7 0 9 2
14 7 13 10 9 1 14 3 0 9 14 9 0 9 2
35 0 9 13 3 14 15 2 16 13 0 2 16 13 0 9 2 16 15 13 13 1 9 1 10 9 7 10 9 7 15 10 9 3 13 2
30 14 1 15 13 0 9 7 15 13 9 9 2 16 1 15 1 0 9 13 9 2 16 15 13 2 2 15 7 0 2
19 1 0 9 15 13 9 2 0 13 10 9 7 1 9 15 13 1 9 2
13 0 13 10 9 7 15 3 1 15 13 7 13 2
32 1 10 0 9 3 13 2 2 9 2 16 13 10 9 1 14 0 9 2 16 4 15 13 1 9 2 13 1 15 0 9 2
10 3 14 4 10 9 13 13 1 9 2
9 13 15 4 1 9 1 0 9 2
14 3 4 14 11 13 10 0 11 1 0 9 10 9 2
9 13 4 2 3 13 0 7 0 2
17 3 15 4 13 1 15 7 15 1 0 9 13 1 9 10 9 2
17 1 0 9 13 3 1 10 9 7 10 9 3 13 1 9 9 2
21 14 15 13 13 2 16 13 15 0 1 0 9 1 15 0 7 13 1 15 0 2
13 1 0 9 14 13 14 15 2 7 14 1 0 2
9 1 0 9 9 13 1 10 9 2
18 9 9 13 1 15 9 7 0 9 2 16 13 9 7 15 3 13 2
3 9 13 2
9 13 15 3 9 2 7 13 13 2
7 1 9 15 15 13 3 2
4 15 3 13 2
4 3 14 13 2
7 13 15 2 16 13 0 2
2 13 2
4 4 13 9 2
2 13 2
8 11 13 7 15 3 13 9 2
12 13 0 0 9 7 15 13 1 15 14 0 2
4 0 9 13 2
10 3 16 13 9 7 9 1 0 9 2
6 15 13 14 0 13 2
16 3 15 13 2 16 15 4 0 9 11 1 9 13 10 9 2
4 13 4 0 2
15 7 4 3 13 13 9 3 2 16 15 4 13 7 13 2
10 7 7 15 13 2 13 14 0 9 2
16 13 9 2 16 15 13 0 9 3 0 2 3 4 13 0 2
15 13 15 3 2 3 4 15 13 9 2 1 15 4 13 2
2 14 2
16 1 0 9 9 3 13 2 3 13 12 9 2 16 13 0 2
33 13 7 3 2 16 13 14 1 9 0 9 1 9 7 9 2 16 15 1 9 13 9 7 7 3 13 2 16 4 9 3 13 2
7 1 9 15 13 3 3 2
25 12 1 0 0 9 1 9 13 2 16 9 0 1 15 13 14 0 9 2 0 9 7 15 0 2
6 9 13 14 0 9 2
24 16 1 15 14 13 13 2 3 15 7 0 13 10 9 2 1 9 2 16 15 3 3 13 2
8 9 2 9 13 7 3 13 2
6 3 15 13 7 13 2
6 13 15 1 0 9 2
5 13 9 1 9 2
8 13 9 7 15 13 1 9 2
5 13 15 1 9 2
8 13 7 1 9 3 13 9 2
9 13 14 9 7 13 9 1 9 2
9 13 15 3 3 1 10 0 9 2
16 13 15 2 16 15 4 9 0 0 9 1 10 9 3 13 2
13 16 13 3 0 13 9 0 0 9 2 13 0 2
26 14 2 16 15 13 2 16 9 3 13 2 16 14 13 1 9 2 16 13 3 0 13 1 15 15 2
25 13 2 16 0 9 13 9 2 7 16 15 13 1 0 9 7 9 1 0 9 2 3 13 9 2
17 9 1 9 7 13 3 0 2 16 13 9 3 3 0 13 3 2
16 9 7 9 7 14 13 10 0 9 7 7 15 3 3 13 2
37 0 7 1 0 9 0 9 11 11 4 1 10 0 0 9 2 12 0 9 11 2 13 14 0 0 9 7 9 7 3 9 13 14 0 0 9 2
23 1 0 9 2 16 4 13 1 10 9 7 1 15 9 0 9 2 4 13 16 1 9 2
12 9 13 3 2 7 14 1 11 4 3 13 2
5 9 9 13 0 2
4 13 0 9 2
20 1 15 13 0 13 2 16 3 3 13 2 16 15 14 14 4 13 3 13 2
22 0 0 9 2 16 15 13 1 9 0 9 2 4 13 3 0 7 3 0 0 9 2
15 0 9 4 13 14 1 9 3 15 2 15 13 14 3 2
3 0 9 2
19 1 9 2 16 4 13 1 0 0 9 2 4 9 13 0 2 0 9 2
2 3 2
28 16 9 14 4 13 13 1 9 1 9 2 16 9 14 4 13 1 9 13 9 2 1 15 4 3 13 9 2
2 14 2
3 4 13 2
7 9 15 4 13 13 9 2
14 9 0 9 15 14 1 9 14 13 13 9 2 2 2
13 9 15 14 13 13 14 9 2 16 13 1 9 2
16 3 13 9 0 2 9 7 9 4 15 1 9 3 3 13 2
2 0 2
37 13 4 2 16 4 13 11 1 9 11 2 16 4 3 1 0 9 13 9 2 13 0 0 9 1 0 9 3 2 16 4 10 11 13 1 9 2
8 1 15 4 13 9 1 11 2
18 10 9 4 11 11 13 13 1 9 10 9 1 9 16 10 0 9 2
15 3 15 15 4 13 2 16 15 10 9 14 13 1 15 2
14 10 9 4 13 2 3 4 13 15 0 13 10 9 2
5 15 4 14 13 2
15 3 4 14 1 10 9 13 13 9 2 16 13 3 0 2
12 15 13 9 1 15 2 0 9 13 1 9 2
12 9 1 15 15 13 9 2 7 15 13 13 2
20 10 9 15 13 14 1 0 9 1 15 2 16 14 4 1 9 13 1 9 2
31 14 4 9 14 13 1 0 9 7 15 1 15 14 13 14 2 7 13 14 1 0 9 15 2 16 4 3 13 1 9 2
26 16 4 13 11 0 0 9 2 16 4 13 0 9 12 2 4 1 15 0 7 0 9 13 0 9 2
30 7 3 15 4 13 2 16 4 1 0 9 1 0 2 0 9 13 12 0 9 2 16 15 4 3 1 10 9 13 2
39 16 4 0 0 9 7 2 0 0 0 9 2 11 11 1 9 9 1 10 9 3 13 0 9 2 4 15 0 9 13 2 9 1 9 7 13 0 9 2
16 11 11 4 14 3 1 0 0 9 12 9 13 1 0 0 2
13 0 9 13 14 9 1 9 2 16 15 13 9 2
13 0 9 13 7 13 0 9 2 7 15 9 13 2
15 14 9 1 0 9 7 0 9 13 0 9 7 13 9 2
20 10 9 14 4 13 9 2 16 15 4 1 9 1 9 13 9 1 0 9 2
8 9 13 0 7 14 3 13 2
14 2 3 13 1 11 12 0 2 16 14 13 0 9 2
11 4 1 9 13 0 9 2 0 1 9 2
18 12 1 9 1 9 13 15 2 16 13 9 0 9 9 9 1 9 2
29 1 0 9 1 9 2 16 13 9 2 13 14 3 9 0 9 1 9 2 15 13 1 12 9 0 9 12 9 2
16 0 9 2 1 9 2 12 9 2 15 3 13 9 7 9 2
7 3 4 13 14 1 9 2
22 1 9 7 9 1 10 9 4 13 12 9 7 14 10 9 13 1 12 9 1 9 2
4 14 13 0 2
7 15 3 13 1 0 9 2
27 10 9 15 4 13 2 16 13 13 14 15 7 1 10 9 2 9 7 13 3 13 2 16 15 14 13 2
18 7 3 14 13 13 0 0 9 1 15 2 10 9 3 13 1 15 2
27 1 0 9 13 13 3 0 9 9 1 11 2 0 9 1 9 7 0 0 9 2 16 13 9 7 9 2
21 9 15 1 9 13 1 9 7 9 2 13 15 13 0 9 7 3 0 9 11 2
19 9 9 13 11 11 2 9 1 0 9 2 16 15 4 3 13 0 9 2
22 9 4 13 9 11 2 11 2 11 2 11 7 9 0 0 9 7 9 0 0 9 2
26 11 2 16 15 11 13 2 3 10 9 2 2 13 13 2 9 2 9 2 7 15 0 9 14 13 2
22 9 11 2 11 11 2 9 2 9 7 9 9 1 0 11 7 15 13 14 1 9 2
38 11 2 12 2 16 4 13 9 1 11 1 9 3 1 12 9 1 0 9 0 9 1 0 9 2 4 13 9 2 16 4 13 1 9 1 9 9 2
15 14 7 4 13 9 2 4 3 13 0 9 2 0 3 2
31 16 4 1 0 9 13 1 0 0 9 10 0 0 9 2 16 4 13 3 0 1 0 0 9 2 7 1 3 13 13 2
20 7 13 3 0 2 16 4 13 1 11 3 3 2 16 16 15 4 15 13 2
28 11 2 9 1 0 9 8 11 1 0 9 11 11 13 2 16 14 4 13 3 0 7 0 9 9 16 3 2
7 11 10 9 3 13 9 2
5 9 9 3 13 2
24 11 13 2 16 13 9 0 2 13 15 14 14 1 0 9 2 16 14 4 13 1 0 9 2
28 11 4 3 7 13 9 1 0 9 2 3 16 4 11 14 3 13 1 9 2 16 7 13 0 1 9 9 2
23 9 0 9 4 1 0 0 9 1 11 1 9 13 1 0 9 11 1 12 2 12 2 2
11 10 9 1 9 4 13 0 9 11 11 2
39 1 0 9 11 1 9 1 11 2 16 4 13 0 7 0 9 11 1 15 0 2 4 13 1 0 9 2 0 4 1 9 7 9 9 13 14 9 9 2
25 14 1 0 9 1 9 7 4 10 9 3 3 1 0 9 13 1 0 0 2 0 7 0 9 2
15 0 9 11 4 3 3 13 7 14 13 13 1 9 9 2
9 2 3 4 14 13 7 4 13 2
19 1 9 0 9 15 13 13 0 9 9 7 1 15 3 13 1 0 9 2
29 1 0 1 11 13 1 9 2 12 9 2 3 0 2 7 4 9 1 0 9 1 12 9 3 13 1 0 9 2
18 0 9 13 0 7 14 1 9 15 4 9 7 9 13 1 12 9 2
9 1 15 0 4 13 10 0 9 2
24 9 1 3 1 11 4 13 9 7 9 11 11 2 1 9 7 9 7 4 3 13 9 11 2
5 2 14 2 13 2
9 1 0 9 0 9 13 1 12 2
17 1 11 14 1 9 0 9 14 13 3 2 7 13 1 0 9 2
37 10 0 9 3 4 13 1 9 9 11 0 0 9 2 16 15 1 9 1 0 9 9 1 0 0 9 1 9 13 1 12 0 9 2 9 2 2
31 7 13 4 1 9 1 9 14 1 9 11 0 9 2 16 15 9 13 14 9 1 11 7 16 15 1 9 13 0 9 2
9 15 15 4 13 0 9 1 9 2
17 7 13 2 14 15 2 16 4 13 0 9 2 15 14 4 13 2
21 14 15 1 12 9 11 2 16 4 15 13 1 0 9 2 15 0 9 4 13 2
14 3 12 9 13 1 0 0 9 11 11 14 12 9 2
15 13 7 3 2 1 9 2 7 3 11 3 14 4 13 2
5 13 3 1 11 2
8 1 3 3 4 13 12 9 2
4 14 13 0 2
7 13 2 13 4 0 9 2
26 16 4 15 15 13 1 9 2 4 13 2 16 13 1 9 2 3 7 4 13 14 10 9 1 15 2
11 13 4 15 3 2 3 7 3 4 13 2
18 16 13 0 7 14 0 9 2 13 9 16 9 7 13 10 10 9 2
10 3 13 2 13 7 15 3 3 13 2
9 3 7 1 9 9 14 3 13 2
21 16 0 13 9 3 3 0 2 0 2 0 2 0 9 2 3 13 0 1 9 2
17 15 13 14 1 9 2 16 4 13 0 13 1 0 9 7 9 2
13 16 9 13 9 2 15 15 3 13 1 9 9 2
15 16 7 15 9 13 15 10 2 9 2 2 3 13 9 2
19 3 15 9 16 9 13 3 2 16 16 4 13 12 1 15 9 7 9 2
15 9 13 1 11 1 0 0 9 2 16 13 9 7 9 2
12 9 4 3 13 10 0 9 2 16 4 13 15
4 13 4 11 2
8 1 10 9 4 13 10 11 2
2 3 13
9 11 11 13 1 11 1 0 11 2
12 3 0 9 9 0 9 7 13 1 0 9 2
21 15 13 1 0 9 2 1 9 2 9 2 9 7 13 3 0 9 9 1 9 2
10 7 3 13 14 1 9 9 1 9 2
16 15 4 0 9 13 9 7 15 13 9 7 1 15 13 9 2
23 2 3 9 1 0 9 7 9 13 7 1 3 0 9 13 9 9 2 16 15 15 13 2
16 2 13 15 4 14 1 11 2 16 4 13 1 9 9 9 2
34 11 2 0 9 1 12 9 2 16 14 4 15 16 0 9 1 11 13 13 1 9 7 3 2 13 0 3 13 2 13 11 11 11 2
9 9 9 14 4 13 12 9 9 2
18 1 9 4 13 13 2 15 13 0 7 0 9 9 1 3 0 9 2
15 12 1 12 0 9 0 9 4 1 9 14 13 0 9 2
1 11
9 1 0 9 3 3 4 13 3 2
20 0 9 4 14 13 10 9 2 9 9 2 4 7 15 13 1 9 7 9 2
25 11 0 8 8 1 9 11 7 12 2 0 8 8 1 11 4 13 1 9 1 0 9 13 9 2
20 8 8 4 13 1 9 2 1 0 9 13 9 1 9 7 15 13 1 9 2
40 16 1 9 4 13 9 2 4 9 13 1 9 1 9 2 16 4 13 8 8 9 4 3 13 0 7 8 8 13 1 9 9 2 16 4 0 9 3 13 2
3 2 8 2
14 12 1 15 13 14 0 7 13 14 14 1 0 9 2
17 14 3 4 9 9 1 9 1 9 13 9 12 9 9 1 9 2
17 13 7 2 16 9 1 9 1 2 0 7 0 2 14 13 13 2
26 9 9 11 13 1 9 1 9 13 0 9 1 9 10 9 10 9 1 9 1 9 0 7 0 9 2
19 1 9 9 14 4 0 9 2 16 15 13 2 1 12 9 13 0 9 2
17 1 9 14 4 13 10 0 9 2 16 4 13 9 7 13 9 2
27 3 4 13 14 0 2 7 13 0 9 14 3 2 16 3 3 15 0 1 9 3 0 13 1 0 9 2
10 0 9 7 3 13 0 14 1 9 2
38 2 6 2 3 4 13 10 0 9 2 2 4 3 1 9 1 9 13 9 2 16 15 4 1 0 0 9 13 1 9 0 9 1 9 12 2 12 2
19 3 4 13 1 9 0 0 9 1 9 1 0 9 2 13 4 15 9 2
23 0 9 2 3 7 3 2 7 0 9 13 9 2 9 3 13 0 7 0 9 1 9 2
11 0 13 13 2 16 13 10 9 10 9 2
15 3 4 13 9 7 15 1 0 9 13 1 10 0 9 2
11 3 3 15 9 13 2 3 13 14 3 2
7 13 15 3 12 9 9 2
25 0 9 15 3 13 16 14 1 9 2 3 7 15 13 0 9 1 0 12 9 9 7 1 9 2
4 3 15 13 2
4 3 4 13 2
9 9 13 1 9 2 9 13 7 13
29 1 0 0 9 15 4 13 2 16 0 9 14 13 9 0 7 0 9 2 15 4 13 14 3 0 1 0 9 2
21 7 4 15 9 12 13 1 12 0 9 2 1 15 4 15 13 14 9 0 9 2
9 9 7 11 7 0 11 4 13 2
6 13 3 1 0 9 2
30 3 13 9 0 9 7 9 9 1 9 9 7 14 9 1 0 9 2 4 13 9 9 2 16 4 15 13 9 12 2
3 2 8 2
16 0 15 4 10 9 13 14 1 12 2 0 8 8 1 11 2
29 16 4 13 0 7 1 0 0 9 2 14 3 7 13 0 9 0 9 2 4 15 1 12 0 9 13 1 9 2
9 14 15 4 13 13 9 1 9 2
3 2 8 2
8 0 9 15 13 1 12 9 2
24 10 9 4 3 13 10 12 9 2 15 15 14 4 13 14 9 9 2 16 4 13 3 0 2
13 0 9 1 9 9 13 0 1 12 1 12 9 2
25 13 15 4 1 12 7 1 12 9 7 16 13 9 0 2 15 4 3 13 1 9 1 12 9 2
13 13 4 14 10 9 2 14 3 13 9 2 2 2
14 9 13 13 16 9 7 9 2 16 13 13 16 9 2
13 0 9 15 13 2 9 13 1 9 9 1 9 2
19 9 11 1 0 9 1 9 1 12 9 13 9 2 0 0 9 7 9 2
8 9 13 9 0 14 1 9 2
41 15 13 3 0 9 0 0 9 11 1 0 9 2 14 4 1 0 9 13 1 0 0 2 0 9 9 1 0 11 1 9 9 2 16 15 1 9 13 1 9 2
35 3 4 2 16 4 13 2 1 15 7 1 9 9 9 1 15 2 9 12 2 12 7 12 2 13 14 0 9 1 9 2 9 7 9 2
23 1 12 9 9 12 2 16 4 11 13 0 9 11 2 7 4 13 0 9 14 3 13 2
17 9 4 3 13 9 9 1 9 1 9 9 9 1 9 0 9 2
9 9 4 13 1 12 9 0 9 2
15 0 9 13 14 0 9 1 9 9 1 9 9 0 9 2
29 3 4 0 0 9 2 11 2 3 13 0 9 2 3 12 9 9 2 2 16 4 13 10 16 12 9 7 9 2
25 9 0 9 4 7 1 0 9 13 10 9 2 7 4 1 9 1 9 0 9 13 10 0 9 2
40 9 2 1 15 13 14 2 9 2 1 12 9 9 9 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 7 11 2 2 13 1 0 9 2
38 3 4 15 13 0 1 9 2 16 4 13 12 9 12 9 2 16 4 13 0 9 9 2 7 4 15 13 1 14 0 9 2 12 9 12 9 2 2
8 1 15 13 10 9 0 9 2
27 1 0 9 13 1 9 12 9 3 2 1 9 2 2 1 9 7 15 13 0 3 1 12 9 1 9 2
9 9 13 1 0 9 7 0 9 2
14 1 0 9 4 1 11 3 13 14 3 12 9 9 2
47 11 11 2 11 2 4 10 9 1 10 9 13 1 9 2 14 3 4 13 0 9 2 16 4 15 10 9 3 13 1 10 9 7 1 10 9 2 1 15 3 1 11 13 10 12 9 2
18 9 15 13 0 2 9 4 15 1 11 7 11 3 13 1 0 9 2
16 1 0 9 4 13 9 1 9 7 9 2 3 3 15 13 2
10 1 12 9 1 11 14 13 3 15 2
13 0 9 13 1 0 9 2 16 4 15 3 13 2
47 1 0 9 11 2 16 4 13 12 0 9 1 0 9 2 4 1 0 2 15 9 4 13 0 9 2 1 12 9 1 10 9 0 9 13 11 11 11 2 11 11 7 4 13 0 9 2
17 9 4 3 13 14 1 11 2 11 2 11 2 11 7 0 11 2
19 1 11 4 15 1 9 9 13 1 10 9 2 16 7 4 15 3 13 2
47 7 14 13 2 16 0 1 0 9 13 3 0 2 16 15 13 2 1 0 0 9 2 0 12 0 9 7 0 1 12 9 2 4 13 9 12 1 12 9 13 12 9 2 3 9 2 2
47 16 15 1 15 13 9 9 1 0 9 1 9 2 13 15 3 0 1 3 2 3 0 9 2 16 9 13 1 3 0 0 9 2 16 3 13 0 9 7 15 3 13 3 3 0 9 2
27 1 15 7 14 13 15 0 1 9 0 9 2 16 15 13 1 9 7 16 4 1 0 9 13 1 9 2
18 9 0 9 13 2 16 15 13 2 7 14 0 9 13 9 1 15 2
22 1 0 0 0 9 2 16 1 9 12 0 9 13 0 9 2 13 3 1 12 9 9
22 0 9 11 11 4 1 11 13 2 16 4 13 3 1 0 9 9 10 9 3 0 2
19 14 3 0 13 1 0 9 2 7 4 13 15 0 10 9 1 10 9 2
31 0 9 4 7 3 1 0 9 13 1 9 12 0 9 2 16 13 0 9 3 0 9 2 16 13 0 1 9 1 9 2
15 3 1 9 1 0 12 14 13 0 9 1 3 0 9 2
21 11 15 4 3 13 10 0 9 1 9 1 0 9 2 16 13 1 9 0 9 2
10 13 2 16 15 3 13 14 1 9 2
7 15 13 10 9 2 13 2
41 9 2 0 1 11 2 16 4 1 10 0 9 13 14 9 9 0 9 2 4 13 1 9 1 10 0 9 2 16 7 4 13 13 15 2 15 4 13 14 15 2
8 3 3 15 13 2 4 13 2
5 7 3 13 9 2
3 2 8 2
39 14 3 0 13 3 0 9 9 2 16 4 13 15 9 10 9 2 3 0 7 0 1 0 9 13 14 0 9 2 16 13 0 1 9 10 9 1 9 2
19 1 11 4 1 10 9 13 9 9 12 9 2 16 15 13 16 9 9 2
33 0 9 1 9 7 9 13 1 0 0 9 0 1 0 0 9 1 9 2 1 15 0 9 13 1 0 9 3 0 9 9 11 2
7 3 13 1 0 9 8 2
18 1 9 7 0 9 9 1 9 9 14 0 9 3 13 14 9 9 2
9 10 9 7 13 14 0 0 9 2
8 10 9 4 13 8 11 11 2
12 10 9 13 14 9 12 0 9 1 0 9 2
4 9 9 13 2
19 15 15 13 14 1 0 9 1 9 2 1 0 9 7 13 15 14 9 2
19 9 14 13 9 9 0 0 9 2 7 13 15 1 10 9 9 1 9 2
30 9 1 9 0 9 1 9 4 14 1 9 13 0 9 1 9 0 2 0 7 0 9 1 12 7 9 1 0 9 2
12 15 4 15 3 13 2 16 4 9 3 13 2
8 1 9 14 13 1 0 9 2
26 1 0 9 15 9 13 1 0 7 14 0 0 9 2 16 9 9 7 0 9 15 3 14 4 13 2
31 1 10 9 13 3 3 3 0 9 2 16 4 9 9 13 1 10 0 9 1 9 2 3 7 4 15 13 9 9 9 2
26 9 9 1 9 9 8 11 11 7 4 13 2 3 13 9 2 16 15 13 9 9 2 0 1 9 2
12 1 15 7 13 9 2 16 13 9 1 9 2
25 11 11 2 0 9 1 0 0 9 2 4 1 11 13 12 9 2 1 10 9 7 13 12 9 2
18 11 2 12 1 9 3 4 1 9 11 13 1 9 1 0 0 9 2
22 1 9 13 0 0 9 1 0 7 0 9 2 16 1 15 13 9 14 1 0 9 2
21 0 9 13 14 3 0 1 0 9 2 15 13 2 16 13 13 2 13 0 9 2
18 9 9 1 0 9 2 0 9 7 0 9 7 13 1 10 9 15 2
16 14 15 13 0 2 16 9 14 13 0 9 1 0 0 9 2
7 15 13 10 9 1 15 2
9 11 4 10 9 1 9 3 13 2
9 3 15 4 13 7 13 10 9 2
10 3 4 15 3 13 0 9 2 2 2
7 14 13 0 13 10 9 2
13 2 1 9 1 11 15 4 0 9 13 0 9 2
12 3 13 0 9 2 16 13 1 9 0 9 2
11 1 0 9 4 0 9 13 9 7 9 2
13 10 12 9 15 4 1 10 9 13 13 0 9 2
17 0 4 13 9 7 0 9 2 0 9 7 0 7 0 9 9 2
10 10 9 4 13 0 2 0 2 0 2
6 9 4 13 1 9 2
8 9 11 11 4 13 13 9 2
12 9 15 4 13 1 11 1 9 7 1 9 2
13 3 4 13 14 14 13 1 0 9 9 11 11 2
8 15 4 13 1 9 1 9 2
7 1 9 15 4 13 9 2
12 9 2 16 4 13 2 4 3 13 1 9 2
18 9 4 13 9 2 7 4 13 1 15 0 1 15 13 14 0 9 2
21 3 4 13 12 9 2 3 7 4 9 13 0 9 9 2 16 16 13 0 9 2
4 13 15 4 2
16 1 9 2 9 9 7 9 2 4 13 0 0 7 0 9 2
21 9 4 3 13 7 13 15 1 10 9 2 1 9 7 15 4 13 14 0 9 2
4 9 4 13 2
22 2 16 15 4 13 2 7 15 13 9 2 16 13 1 9 2 2 4 13 11 11 2
12 13 15 4 7 15 1 0 9 13 1 9 2
16 13 4 13 0 3 12 9 2 7 4 14 13 13 9 9 2
14 9 4 3 13 1 9 2 9 7 4 3 13 9 2
6 13 4 9 7 9 2
7 9 4 13 1 0 9 2
8 11 4 1 10 9 13 9 2
8 1 15 4 13 14 0 9 2
17 1 9 4 9 13 1 3 0 9 2 16 4 15 9 3 13 2
14 9 1 11 4 13 9 2 13 15 4 9 1 9 2
18 0 9 4 15 3 13 1 9 2 16 15 4 1 10 9 13 15 2
16 1 9 4 9 3 13 7 13 2 16 4 9 3 13 9 2
19 0 4 13 13 1 12 1 0 9 0 9 2 16 4 15 13 10 9 2
6 13 15 4 1 11 2
13 0 9 4 13 7 15 1 0 9 3 13 9 2
13 13 4 13 9 2 16 15 4 4 3 3 13 2
15 2 10 9 13 0 9 7 0 9 2 0 9 0 9 2
5 13 7 0 9 2
17 9 15 4 13 3 1 15 2 13 15 4 2 16 16 15 13 2
7 9 4 13 3 3 0 2
13 11 15 4 13 1 9 7 15 1 9 13 3 2
5 9 4 15 13 2
14 9 15 4 13 1 9 2 9 4 15 13 1 9 2
8 1 9 15 15 4 13 9 2
13 0 9 9 15 4 13 16 9 1 0 0 9 2
13 13 15 15 4 2 16 4 1 15 13 2 2 2
20 13 4 13 2 15 13 7 3 13 1 9 2 7 1 10 9 4 13 9 2
14 3 4 13 14 3 3 2 16 15 3 14 4 13 2
12 9 7 15 4 14 3 13 3 2 1 9 2
36 2 16 3 13 2 15 14 14 14 13 2 15 3 10 9 13 2 16 0 9 13 2 16 3 13 0 9 2 16 13 3 0 1 10 9 2
6 15 4 13 0 9 2
14 3 16 15 13 1 9 10 9 2 3 15 4 13 2
21 2 3 1 10 9 0 9 14 13 14 2 2 4 13 11 2 16 4 13 9 2
7 2 9 13 0 1 9 2
19 11 15 4 14 13 13 2 16 15 4 9 3 13 7 15 4 9 13 2
13 11 4 13 13 14 14 2 3 4 13 1 9 2
14 13 4 3 2 16 4 15 13 1 9 0 0 9 2
16 13 4 14 3 0 2 16 16 4 13 9 1 9 0 9 2
20 11 4 3 13 2 16 13 9 1 9 0 2 9 4 13 0 3 12 9 2
12 13 15 4 2 16 13 0 1 9 7 9 2
12 3 4 13 13 14 0 9 2 9 2 9 2
15 1 0 9 2 1 9 2 7 4 1 0 9 13 9 2
10 10 9 1 11 1 11 4 13 0 9
22 11 15 4 13 7 13 3 2 1 11 2 16 4 13 15 12 9 1 15 1 9 2
21 13 4 0 1 9 2 1 15 4 13 10 10 9 2 7 13 4 0 7 0 2
11 11 4 13 9 2 16 4 13 0 9 2
12 13 4 9 2 9 4 13 7 9 4 13 2
9 3 4 13 7 15 3 13 3 2
8 1 9 7 9 4 3 13 2
16 3 4 11 13 0 0 9 7 9 7 15 15 13 1 9 2
11 3 4 13 0 9 7 13 9 1 9 2
12 3 4 13 7 13 11 2 16 13 1 15 2
12 11 4 13 9 1 9 7 15 15 3 13 2
4 11 4 13 2
7 14 3 14 13 13 9 2
4 1 0 9 2
2 9 2
3 0 9 2
14 14 15 14 13 3 2 7 4 15 0 3 14 13 2
13 3 15 4 13 1 0 9 7 13 1 0 9 2
17 11 15 15 4 0 13 1 9 7 15 13 1 9 1 0 9 2
17 13 15 4 14 1 9 0 9 1 9 2 1 15 4 13 9 2
15 15 13 2 16 16 4 13 9 2 2 15 4 13 11 2
6 13 15 4 0 9 2
10 2 14 0 13 2 16 14 13 15 2
13 1 9 4 13 0 9 13 2 3 13 9 9 2
21 3 15 14 1 0 9 13 1 9 0 9 2 3 16 4 9 13 1 0 9 2
9 13 2 7 4 15 14 13 2 2
8 3 4 13 7 15 13 9 2
11 2 3 3 13 0 9 2 2 4 13 2
6 11 4 14 3 13 2
9 11 15 4 13 7 13 1 9 2
8 1 9 4 14 3 13 9 2
12 16 4 11 13 9 2 4 11 14 14 13 2
7 11 4 14 3 13 9 2
10 2 13 4 13 9 2 2 4 13 2
7 2 9 15 4 3 13 2
17 16 16 15 14 13 1 9 7 9 2 16 15 13 13 2 2 2
2 14 2
6 1 15 15 15 13 2
7 11 4 13 1 0 9 2
15 14 4 15 13 1 9 2 7 15 3 4 13 3 0 2
8 0 7 0 1 9 0 9 2
4 9 9 9 2
30 9 9 11 15 4 14 3 3 13 9 2 16 0 9 4 13 13 2 16 3 1 9 1 0 9 13 0 0 9 2
21 2 4 13 2 16 13 9 9 0 9 2 2 15 4 13 7 15 13 1 9 2
10 11 15 4 0 13 1 9 1 9 2
25 11 4 3 3 13 2 16 4 15 14 13 14 11 7 11 2 16 4 15 3 13 10 9 3 2
23 0 9 15 4 13 1 9 2 16 4 15 13 1 0 9 7 0 9 1 9 1 9 2
10 11 7 11 4 15 14 13 0 9 2
17 11 15 1 9 14 4 13 2 11 7 15 4 13 9 16 11 2
14 11 15 4 0 13 1 0 9 2 16 4 13 11 2
5 11 4 13 9 2
7 1 9 13 3 4 13 2
8 11 4 3 13 9 1 9 2
7 2 13 2 13 14 3 2
9 13 15 1 9 1 9 3 3 2
10 2 13 4 3 1 9 1 10 9 2
6 13 4 15 1 9 2
9 9 2 16 15 13 2 13 0 2
5 9 4 14 13 2
16 11 4 13 2 14 16 15 1 10 0 9 13 9 7 9 2
10 3 15 13 13 1 10 0 9 2 2
10 2 15 13 11 2 2 4 13 11 2
19 11 4 11 7 11 13 1 9 1 0 9 2 1 15 4 13 0 9 2
14 9 4 13 1 9 2 16 4 15 0 14 3 13 2
24 0 9 1 9 4 15 3 13 1 14 0 9 2 7 7 4 11 1 0 9 13 10 9 2
9 14 3 4 1 0 13 7 13 2
9 2 16 13 2 2 4 13 11 2
20 2 1 11 4 13 14 3 0 2 16 4 10 9 13 1 0 1 0 9 2
18 9 4 15 13 7 13 4 1 0 9 2 7 15 4 3 13 15 2
7 14 3 4 13 1 9 2
17 3 4 15 13 3 7 13 0 9 2 16 4 15 13 1 15 2
26 1 11 4 13 1 9 7 13 2 16 4 15 3 14 3 13 2 16 15 4 13 7 13 3 13 2
18 0 4 13 10 9 7 13 9 7 1 9 4 15 13 9 1 9 2
10 10 9 4 13 9 1 9 9 9 2
13 3 4 13 2 16 13 15 3 14 9 1 9 2
15 3 15 15 4 13 2 3 4 0 1 15 13 10 9 2
31 9 15 4 7 13 13 1 9 7 13 4 2 16 4 13 0 9 2 1 15 13 9 9 7 15 1 9 13 1 15 2
19 11 15 15 4 13 2 7 15 4 13 2 16 4 15 13 13 1 9 2
15 9 4 14 13 3 7 13 4 15 2 16 4 9 13 2
10 13 4 1 9 7 15 13 1 9 2
15 2 7 15 4 13 2 2 4 13 7 15 13 1 9 2
19 13 15 4 1 11 7 15 13 2 2 15 13 14 3 2 9 2 14 2
20 2 14 2 15 13 2 2 4 13 11 7 11 3 13 1 9 1 0 9 2
7 11 4 13 10 0 9 2
3 0 9 2
25 1 9 4 15 13 14 1 9 0 9 12 9 12 1 0 9 2 16 4 13 0 0 0 9 2
13 1 0 9 0 9 4 1 11 13 14 9 11 2
9 15 4 13 0 0 9 1 9 2
13 1 12 0 9 13 0 3 13 9 7 15 13 2
23 9 13 0 1 9 2 16 1 9 13 1 0 9 1 9 2 8 8 0 0 9 2 2
10 0 9 1 9 15 3 4 13 13 2
16 2 1 0 9 13 12 9 9 1 9 2 12 9 13 9 2
10 1 11 3 12 9 9 13 10 9 2
20 3 15 16 11 13 9 0 9 9 2 1 15 4 15 1 0 9 13 11 2
20 0 9 0 9 8 11 11 1 0 0 9 1 9 13 2 16 13 3 3 2
54 3 0 2 3 7 3 0 9 9 7 9 1 9 1 11 4 13 1 0 9 9 2 16 4 0 9 2 16 4 13 0 9 3 12 9 9 13 9 2 0 1 0 9 1 11 1 0 9 11 1 0 0 9 2
3 3 0 2
12 0 9 9 7 9 7 13 7 14 13 13 2
5 13 4 3 9 2
32 1 15 2 16 13 0 9 0 9 1 0 2 0 2 0 2 0 7 0 9 2 15 9 14 4 9 7 9 13 1 9 2
16 3 7 4 9 14 14 0 9 10 9 13 1 0 0 9 2
34 10 0 9 4 7 9 10 9 13 1 3 0 9 1 9 7 10 9 2 1 9 9 2 13 1 10 0 9 2 1 10 0 9 2
22 9 9 4 13 9 9 1 9 0 9 1 9 7 1 3 15 13 14 1 9 9 2
27 16 13 2 13 9 9 0 0 9 1 11 2 16 15 3 0 9 13 1 10 0 9 0 9 0 9 2
19 1 0 9 13 3 3 9 2 9 1 0 9 15 13 1 3 0 9 2
22 16 4 1 9 9 9 3 13 3 1 9 9 2 4 13 0 9 0 1 10 9 2
15 10 0 9 4 13 9 2 16 13 9 9 14 3 9 2
23 0 9 2 16 13 2 13 14 15 2 16 15 1 9 9 3 13 0 0 7 0 9 2
24 16 0 13 0 9 7 9 2 4 13 3 3 0 2 7 4 13 14 1 0 9 3 0 2
13 9 9 4 3 13 0 0 9 1 0 9 9 2
35 16 13 3 16 0 2 16 4 0 9 14 13 10 9 2 15 13 7 13 1 0 2 4 13 0 10 0 9 13 14 1 0 9 9 2
14 7 15 1 9 9 13 10 9 2 16 13 9 9 2
15 15 13 2 16 0 0 9 9 3 3 13 1 9 9 2
12 1 15 2 16 4 13 2 16 13 14 13 2
17 3 9 7 3 1 0 0 9 4 13 2 16 4 13 0 9 2
5 13 4 3 0 2
13 10 9 15 4 3 1 0 13 13 1 10 9 2
11 13 4 13 7 15 1 15 14 3 13 2
13 13 4 15 13 1 9 7 9 7 13 4 0 2
10 1 12 9 15 4 13 10 10 9 2
5 13 4 13 9 2
31 3 14 4 13 3 3 13 14 10 0 9 16 9 1 0 9 2 10 9 9 2 16 15 3 13 7 3 10 9 13 2
19 1 12 9 15 9 2 1 12 9 2 13 1 9 2 1 12 9 2 2
20 1 0 9 2 16 13 0 9 13 1 9 2 4 13 13 1 9 10 0 9
29 15 4 1 11 13 14 1 0 0 9 2 3 0 4 13 15 2 16 4 15 1 9 12 13 1 0 0 9 2
28 3 4 13 9 12 2 0 11 11 11 2 16 4 1 9 11 13 0 0 9 0 0 9 1 10 0 9 2
13 0 11 4 13 14 1 10 9 9 0 0 9 2
26 1 11 4 15 13 16 0 0 9 1 9 2 15 14 13 9 11 7 16 0 9 4 13 1 9 2
10 16 0 4 1 10 9 13 14 9 2
23 7 14 3 9 4 13 2 16 4 1 9 1 9 13 15 2 15 3 13 16 0 9 2
6 9 4 13 3 0 2
32 9 9 4 13 9 2 0 1 0 0 9 7 0 9 2 1 9 7 1 9 7 4 13 9 2 9 7 9 2 0 9 2
11 11 11 13 10 9 1 9 1 0 9 2
19 13 7 13 15 15 0 2 15 15 3 13 3 7 1 0 16 0 9 2
8 2 3 3 13 1 0 9 2
15 1 15 15 3 3 13 10 9 2 3 15 13 0 9 2
9 10 12 10 9 13 3 0 9 2
23 14 11 13 0 9 9 2 14 10 9 1 10 9 4 13 1 0 0 9 7 0 9 2
48 14 1 9 15 4 1 0 9 0 9 13 9 11 11 2 1 15 4 3 9 13 1 9 2 1 9 1 9 8 8 2 0 9 2 16 13 3 0 0 9 9 1 9 0 9 1 11 2
17 2 9 1 9 8 8 4 3 13 14 1 9 2 1 0 9 2
13 9 4 15 13 3 1 11 7 13 9 1 15 2
32 3 3 15 4 13 1 11 11 1 10 0 9 7 13 4 2 16 13 15 10 10 9 1 9 2 16 15 14 13 1 9 2
12 1 9 4 13 2 16 15 4 13 1 11 2
15 13 4 15 2 15 13 1 15 7 3 4 13 10 9 2
19 3 0 13 2 16 1 9 0 9 1 9 9 13 0 9 7 0 9 2
21 0 13 9 2 16 4 14 9 9 1 0 9 13 0 2 9 2 1 0 9 2
19 13 15 0 9 0 0 9 2 16 15 1 9 13 3 0 9 0 9 2
8 9 1 15 15 13 1 3 2
4 9 0 9 2
8 9 1 9 13 9 1 9 2
12 1 10 9 9 1 9 13 1 9 0 9 2
20 10 9 3 9 1 9 1 9 13 10 9 11 2 16 13 9 1 11 11 2
17 10 9 4 13 3 10 12 9 9 1 9 9 3 13 1 9 2
23 7 10 0 9 4 3 3 2 10 9 9 1 9 2 0 1 0 13 7 13 4 9 2
16 7 14 10 0 9 9 9 13 3 0 1 0 9 0 9 2
20 10 0 9 9 15 4 13 12 3 3 0 1 0 9 2 0 1 0 9 2
24 1 0 9 14 14 13 0 7 1 15 4 13 9 0 9 2 16 16 4 1 0 9 13 2
20 16 4 1 10 9 13 1 9 12 9 2 15 4 9 13 13 14 12 9 2
17 10 9 13 10 9 2 9 7 9 2 16 13 0 9 1 9 2
27 14 13 10 9 10 9 2 13 1 0 9 9 7 13 9 2 0 9 1 9 2 3 13 1 10 9 2
12 1 0 9 9 2 1 0 9 1 0 9 2
18 13 4 15 1 9 2 9 4 13 9 7 13 1 9 0 9 9 2
40 14 2 15 4 13 11 7 13 1 9 1 9 9 1 0 9 7 9 2 16 4 15 13 1 0 9 1 9 2 7 9 13 14 3 1 9 0 9 0 2
13 7 14 16 10 9 13 2 13 3 13 1 15 2
3 0 9 2
16 9 1 9 0 9 3 13 2 13 15 9 7 13 0 9 2
11 13 2 9 13 1 9 0 9 1 9 2
13 7 11 1 0 9 9 13 2 16 4 3 13 2
2 13 2
12 9 4 13 14 9 9 2 10 0 0 9 2
43 1 9 1 9 7 0 1 9 4 13 2 16 15 4 13 9 10 9 2 10 9 2 9 0 9 2 9 11 2 16 4 13 9 7 9 7 1 10 9 13 1 9 2
6 13 15 4 7 13 2
28 1 9 4 15 14 13 0 9 2 7 4 15 0 3 13 13 2 15 13 9 0 9 2 16 13 1 9 2
5 7 3 13 9 2
20 13 4 1 9 2 1 9 9 2 16 4 1 9 1 9 7 9 13 3 2
20 13 15 4 10 9 7 13 4 0 9 1 9 2 3 4 13 13 1 15 2
4 15 13 3 2
4 13 15 13 2
14 9 11 4 13 3 2 13 4 15 2 16 13 0 2
5 16 13 0 9 2
30 11 4 1 0 9 2 16 4 13 1 0 9 9 1 10 9 2 13 9 1 9 2 13 7 15 3 13 1 9 2
20 1 10 9 4 13 0 9 7 9 2 0 9 3 0 9 4 13 0 9 2
21 1 9 4 3 13 14 16 0 2 9 1 9 7 3 7 4 13 3 0 9 2
7 13 4 14 3 0 15 2
9 13 15 4 1 9 1 0 9 2
17 13 15 4 1 0 9 10 9 2 1 9 4 9 13 10 9 2
20 13 15 4 1 3 0 0 9 2 13 15 4 7 13 2 16 15 9 13 2
4 3 4 13 2
5 13 13 10 9 2
14 10 9 15 4 13 2 3 13 0 13 2 15 13 2
27 14 13 14 10 0 7 3 3 0 9 2 16 4 15 15 13 0 2 0 7 4 15 1 0 9 13 2
22 10 3 0 9 0 9 4 1 0 0 9 1 0 11 13 9 7 9 10 0 9 2
26 1 14 12 0 9 15 4 13 13 3 12 9 12 9 12 9 12 9 1 12 9 1 3 0 11 2
23 1 0 9 9 9 1 9 1 11 11 11 4 13 3 1 0 9 3 0 9 12 9 2
16 15 13 0 9 1 0 2 0 7 0 9 7 0 0 9 2
13 1 9 13 9 2 13 9 7 0 7 0 9 2
8 1 0 13 2 16 15 13 2
32 1 9 9 13 3 0 15 2 15 3 13 1 9 0 9 9 2 8 8 0 9 2 1 15 13 9 7 13 9 1 15 2
9 1 10 0 0 9 13 1 9 2
8 9 13 3 2 9 13 3 2
3 4 13 2
18 16 0 9 0 9 4 13 11 0 1 9 9 11 1 9 11 11 2
22 11 4 1 9 13 1 0 9 7 15 1 9 1 0 9 15 4 13 3 1 9 2
3 13 15 2
8 15 13 9 2 13 7 0 2
7 13 2 16 10 9 13 2
8 0 9 4 13 3 1 9 2
17 9 15 4 13 0 9 0 9 2 7 15 4 13 1 9 9 2
21 9 2 16 4 13 1 11 2 4 13 12 0 0 9 2 7 15 4 13 0 2
5 9 4 13 9 2
4 3 7 3 2
10 10 9 13 14 2 13 14 0 9 2
11 0 9 4 13 1 0 9 1 0 9 2
8 0 9 4 13 0 9 15 2
9 3 13 2 16 13 1 15 9 2
13 3 4 15 3 13 9 2 16 4 13 9 3 2
15 7 13 10 9 2 7 9 7 9 2 0 9 1 11 2
18 3 7 13 3 10 3 0 0 9 9 2 16 13 1 9 1 9 2
18 9 4 13 9 9 2 14 13 15 2 16 15 4 13 14 3 12 2
19 0 9 13 0 13 14 1 9 7 9 1 0 9 7 9 1 0 9 2
20 9 13 2 7 13 3 0 13 11 2 16 13 2 16 4 1 15 11 13 2
14 14 0 9 1 9 7 0 9 9 13 1 0 9 2
12 13 15 1 9 9 7 16 13 9 14 0 2
5 14 4 3 13 2
35 3 4 15 1 9 10 9 1 0 9 13 14 1 0 9 2 16 4 15 13 2 16 4 13 10 12 2 0 9 10 9 13 1 9 2
29 10 2 9 2 1 9 7 9 4 2 13 2 2 16 4 15 14 1 15 2 13 9 2 7 2 13 9 2 2
19 0 4 13 9 9 1 10 9 2 3 13 1 10 9 2 3 14 13 2
15 14 14 3 4 13 3 7 10 9 4 14 13 1 9 2
6 3 4 13 15 0 2
15 10 9 13 3 10 9 7 9 2 16 15 13 14 0 2
21 3 13 2 16 9 2 16 15 4 3 15 13 10 9 1 9 2 13 1 15 2
24 13 4 14 10 9 2 16 4 13 2 15 15 15 4 13 2 7 3 15 4 3 13 9 2
7 1 10 9 9 4 13 2
6 13 4 15 0 9 2
9 15 14 15 13 1 9 10 9 2
5 13 4 10 9 2
8 15 15 4 9 13 1 15 2
6 7 4 15 13 13 2
9 1 9 4 1 15 13 1 15 2
13 3 4 9 1 9 13 15 2 15 4 3 13 2
9 7 16 4 13 2 13 1 9 2
5 3 4 13 3 2
8 15 15 4 1 15 14 13 2
2 15 2
6 15 15 13 0 13 2
7 15 15 4 7 13 13 2
8 7 13 3 13 1 10 9 2
10 3 4 13 0 7 13 1 10 9 2
5 10 9 4 13 2
5 10 9 4 13 2
12 16 15 4 13 9 1 9 1 9 1 9 2
10 3 4 13 2 16 15 3 13 9 2
10 3 4 9 13 3 16 11 1 9 2
8 7 3 9 1 15 4 13 2
2 6 2
2 9 2
4 3 13 9 2
31 13 9 2 16 3 13 9 7 15 13 1 9 2 16 1 0 9 13 1 9 7 1 15 15 13 3 9 9 14 13 2
7 7 3 13 14 10 9 2
6 7 15 4 15 13 2
13 4 13 1 9 14 1 9 2 7 14 1 9 2
4 15 14 13 2
7 7 1 9 13 3 0 2
23 16 3 15 15 14 13 13 2 3 13 15 1 9 2 16 13 2 16 4 13 1 9 2
20 9 15 2 15 14 4 13 9 2 15 13 3 2 16 4 15 0 3 13 2
8 1 15 4 11 13 1 9 2
6 1 15 4 13 9 2
8 2 13 2 2 4 13 11 2
8 2 13 15 2 3 15 13 2
12 3 15 4 13 2 1 15 4 15 3 13 2
2 3 2
3 10 9 2
22 10 10 0 9 15 13 1 9 2 16 4 15 2 16 4 13 9 2 13 0 9 2
7 2 14 2 2 4 13 2
6 2 3 14 13 9 2
3 1 9 2
7 7 3 9 13 0 9 2
11 3 3 13 1 15 2 7 13 0 9 2
24 7 16 4 13 10 9 2 16 4 15 13 2 14 13 15 13 2 14 16 4 13 0 2 2
5 2 9 13 0 2
9 2 7 15 13 2 2 4 13 2
8 2 6 2 2 4 13 11 2
4 2 14 13 2
12 2 13 4 13 9 2 7 4 15 3 13 2
7 2 6 2 2 4 13 2
11 9 4 13 9 2 13 15 4 2 2 2
8 15 13 2 13 1 10 9 2
35 16 4 13 9 7 2 16 4 15 13 2 9 1 15 13 1 10 10 9 2 16 16 4 13 15 2 4 9 9 14 3 13 1 9 2
9 13 4 9 9 7 15 13 9 2
8 14 9 15 4 13 14 13 2
18 14 15 4 13 0 2 16 4 3 13 15 2 16 4 9 13 13 2
12 1 9 9 9 4 13 9 11 3 10 9 2
23 1 0 7 4 1 9 0 9 13 9 0 9 9 2 1 15 9 4 13 0 9 9 2
10 0 9 13 1 9 2 3 14 13 2
9 9 1 9 4 13 0 0 9 2
16 11 2 11 2 11 7 10 0 9 4 13 13 9 0 9 2
15 13 7 0 9 2 1 15 15 3 7 3 13 0 9 2
22 15 13 0 0 9 1 11 2 3 7 13 9 2 1 15 4 13 9 11 1 11 2
10 10 9 13 1 9 7 9 0 9 2
25 0 9 0 9 13 2 16 1 9 10 0 9 14 4 13 13 9 0 0 9 14 3 0 9 2
14 7 1 9 4 3 13 2 16 4 9 13 0 9 2
16 9 9 4 13 0 9 7 1 0 9 4 13 14 1 12 2
17 9 1 9 4 13 1 0 12 9 2 16 4 0 11 13 13 2
6 2 11 13 2 9 2
35 16 4 9 0 9 11 11 3 1 9 9 11 11 1 9 13 0 9 8 11 2 14 4 13 13 2 16 13 10 9 7 9 3 0 2
11 2 12 0 9 4 3 13 1 0 9 2
21 3 4 15 11 13 7 16 4 13 15 14 1 9 9 2 4 13 10 9 9 2
8 13 15 4 13 1 0 9 2
10 14 10 9 4 13 2 15 4 13 2
24 11 2 12 2 9 0 0 9 11 11 11 11 1 9 9 0 12 9 14 4 13 13 9 2
15 13 1 0 9 1 9 2 16 15 4 13 0 0 9 2
19 11 4 13 2 16 4 9 13 14 3 7 16 15 14 13 1 10 9 2
22 11 4 2 13 2 12 9 3 1 9 1 11 2 9 7 4 13 14 9 1 11 2
29 16 9 4 13 9 1 9 2 3 7 4 13 9 2 16 4 13 13 1 0 9 7 13 4 1 9 1 11 2
17 13 4 1 12 2 12 9 7 3 4 13 1 9 1 10 9 2
5 2 9 13 0 2
7 14 7 13 10 9 0 2
36 9 1 11 4 1 9 0 9 13 14 0 9 11 7 11 11 2 1 9 9 7 4 11 13 2 16 15 4 13 1 9 9 9 1 11 2
51 0 9 4 3 1 9 13 2 16 13 9 1 0 9 2 0 7 0 2 2 14 3 7 15 4 13 1 9 13 2 16 15 3 3 16 9 1 3 0 11 13 9 1 3 0 9 2 15 15 13 2
18 1 0 12 9 4 11 13 7 3 10 9 1 9 0 9 1 9 2
46 9 4 13 7 9 4 1 9 12 7 12 13 9 9 2 3 0 0 9 2 3 16 4 1 9 9 1 9 1 9 11 13 10 9 2 16 4 13 12 9 9 9 1 0 9 2
40 7 14 3 0 9 1 0 9 1 10 9 4 13 3 0 2 7 4 1 9 9 9 13 1 11 2 3 16 4 1 0 9 13 14 0 0 9 11 11 2
14 2 8 2 13 0 0 9 2 10 9 2 9 7 9
28 3 16 4 11 3 13 9 2 4 13 1 0 9 11 3 0 2 7 4 3 13 1 0 9 1 0 9 2
14 2 13 13 2 16 4 13 1 9 1 3 0 9 2
20 1 9 1 10 9 4 15 13 3 3 2 7 14 4 13 9 1 0 9 2
17 0 9 4 13 14 3 0 2 15 7 4 13 1 15 10 9 2
15 1 11 4 14 13 3 3 2 3 7 9 1 9 13 2
29 3 14 4 13 10 0 9 2 2 4 1 9 13 11 2 16 4 13 3 0 14 1 0 0 9 1 10 9 2
38 3 4 13 0 9 0 9 7 1 15 13 2 16 4 15 9 0 1 0 1 9 13 7 3 14 13 2 14 16 13 0 0 7 0 9 0 9 2
18 1 0 9 9 1 11 4 9 0 9 13 13 1 15 1 9 9 2
25 10 0 9 4 0 9 1 9 13 2 0 0 9 7 15 4 1 9 13 1 9 1 0 9 2
20 0 9 11 11 4 13 9 9 0 9 7 15 13 2 16 13 1 10 9 2
20 14 11 4 15 3 16 1 0 9 13 1 0 9 2 2 3 13 0 9 2
8 0 4 13 14 1 9 12 2
21 1 9 15 4 7 3 13 2 9 1 10 0 0 9 7 4 13 14 11 11 2
34 0 9 4 13 11 14 1 12 9 2 16 4 1 9 3 3 13 2 16 4 10 3 0 9 11 11 13 14 10 9 1 10 9 2
17 11 15 4 7 1 0 12 9 3 13 2 7 4 3 13 9 2
27 16 4 13 0 11 11 0 1 0 1 9 12 2 13 2 16 4 14 0 2 3 2 13 1 0 9 2
18 9 2 3 15 3 9 13 2 16 13 2 16 4 13 9 0 3 2
13 11 2 0 3 13 7 3 1 9 11 13 9 2
26 0 9 4 13 3 1 10 9 7 7 4 13 1 0 1 11 2 16 4 3 13 10 9 1 9 2
30 16 4 15 0 9 13 2 16 13 9 2 7 4 13 1 9 10 9 2 4 10 9 13 12 1 12 7 13 3 2
19 9 11 11 11 13 3 10 9 1 9 1 9 9 9 1 10 0 9 2
9 1 0 9 9 3 13 0 9 2
40 1 0 9 7 9 4 9 1 0 9 0 9 11 11 3 13 1 10 9 2 16 4 3 14 0 9 13 3 3 1 15 2 7 7 0 9 14 3 13 2
23 11 13 2 16 13 15 0 9 9 9 2 7 14 13 3 0 1 9 9 0 9 11 2
10 11 2 2 1 9 13 3 16 0 2
7 3 4 10 9 13 9 2
12 3 15 13 2 16 15 3 14 13 13 9 2
28 11 4 0 9 13 9 1 9 1 0 9 2 7 15 14 13 13 2 16 4 13 1 10 9 0 1 9 2
13 15 4 13 15 1 9 1 9 7 1 0 9 2
24 11 2 16 13 9 3 0 2 4 1 0 9 13 2 16 11 11 9 14 4 13 1 11 2
33 16 15 15 4 13 13 2 4 13 2 3 4 13 1 0 9 1 0 9 1 9 2 16 4 15 13 9 11 2 3 3 0 2
27 7 1 9 1 11 11 4 13 0 2 16 1 15 14 13 15 2 7 14 4 15 0 11 13 3 3 2
31 16 13 0 2 14 4 0 9 9 1 9 1 0 9 13 12 9 2 15 13 3 3 3 3 2 16 4 13 3 0 2
43 10 9 1 9 1 0 9 1 0 12 2 16 4 13 2 16 4 1 0 9 14 3 13 2 4 13 3 14 9 9 1 9 2 7 14 4 13 14 3 0 13 11 2
17 1 15 13 14 15 2 16 4 10 9 1 11 13 14 11 11 2
10 14 3 4 13 14 10 9 3 0 2
17 16 4 0 1 15 13 2 16 14 13 2 4 13 9 3 0 2
2 14 2
19 14 15 13 13 1 9 1 10 9 2 3 13 1 0 9 7 0 9 2
14 1 9 1 9 15 13 13 9 1 9 7 13 9 2
19 11 11 11 7 11 11 11 4 3 3 3 13 9 0 9 1 0 9 2
19 9 2 1 15 4 1 10 9 13 3 2 4 1 9 13 14 0 9 2
14 2 8 2 13 0 0 9 2 10 9 2 9 7 9
2 13 2
28 3 15 4 3 13 2 16 4 11 13 1 9 7 15 13 9 1 9 2 3 1 9 7 4 13 10 9 2
15 3 13 0 1 15 2 15 9 15 14 1 9 13 9 2
35 14 3 1 9 14 14 13 13 10 0 9 2 7 15 15 3 13 2 16 14 1 9 13 0 9 2 16 3 13 7 13 14 0 9 2
15 15 13 14 3 9 2 16 14 4 1 11 13 3 0 2
36 3 13 9 2 16 4 15 1 15 2 16 4 3 13 1 11 7 11 2 13 3 3 7 3 3 3 3 1 0 9 1 11 1 10 9 2
43 9 4 13 2 16 0 9 9 13 1 11 2 1 0 11 7 15 13 3 2 16 13 0 0 9 7 0 9 2 16 4 13 0 1 9 9 2 16 13 9 1 15 2
30 3 7 15 4 0 9 3 3 13 7 0 9 4 1 0 9 13 14 12 0 2 16 13 0 3 1 9 0 9 2
28 12 0 9 1 9 9 4 13 1 0 9 11 3 0 9 1 11 2 7 15 15 9 1 9 9 14 13 2
31 14 14 13 9 3 13 2 16 13 1 11 1 14 1 10 9 10 0 0 9 2 1 15 4 0 9 3 13 10 9 2
11 1 0 9 14 0 0 9 14 13 14 2
43 7 9 0 9 1 11 13 2 16 10 0 0 9 14 13 1 11 2 1 16 9 9 3 13 1 0 9 2 16 15 14 13 7 15 1 0 9 13 14 1 9 9 2
38 16 4 1 10 0 0 9 3 13 3 3 2 4 9 13 14 10 0 9 2 15 14 14 13 1 10 0 0 9 2 16 15 3 13 3 1 9 2
33 15 0 4 13 3 14 9 9 2 16 13 2 16 15 10 9 2 16 15 13 1 9 2 3 13 9 7 7 13 3 1 9 2
25 0 9 13 0 1 11 3 0 9 0 9 2 1 11 7 1 15 13 14 14 8 8 0 9 2
20 12 7 0 13 9 12 9 10 9 2 16 15 13 1 3 0 0 0 9 2
30 1 9 10 7 0 0 9 13 0 11 0 1 0 9 1 9 7 9 0 9 1 9 9 9 0 9 11 9 11 2
17 3 0 9 4 11 13 3 1 9 7 9 15 4 3 3 13 2
18 9 13 3 9 2 1 15 9 13 9 3 2 16 3 13 1 9 2
25 10 9 15 13 2 16 14 1 9 9 7 0 9 3 13 2 1 10 9 4 9 13 1 9 2
33 9 2 1 15 9 3 13 2 13 14 0 9 2 7 7 9 13 0 0 9 7 1 9 13 9 2 16 15 13 9 1 9 2
20 1 9 9 3 13 0 2 1 0 9 7 15 13 13 2 15 13 2 13 2
23 16 0 9 7 9 15 9 13 14 1 0 11 11 2 0 1 0 9 2 0 1 9 2
7 15 7 3 3 15 13 2
23 9 15 13 9 2 16 13 9 2 16 15 13 1 15 2 0 7 0 2 13 3 3 2
32 3 15 9 13 0 9 2 16 1 10 0 9 13 0 2 13 2 16 4 15 13 9 7 16 1 9 13 13 10 9 14 2
24 11 2 1 9 2 12 9 2 1 12 9 3 15 4 9 9 1 11 13 1 0 0 9 2
32 0 9 0 9 1 9 4 1 9 1 0 9 11 2 16 15 13 11 7 11 11 2 13 9 0 9 0 9 1 9 11 2
18 1 9 4 13 12 9 1 11 2 0 9 2 11 2 11 7 11 2
25 9 13 0 2 16 4 0 9 2 16 4 14 13 0 9 11 2 13 1 0 9 14 0 11 2
12 0 9 1 9 4 13 0 9 11 7 11 2
18 9 13 3 3 0 2 13 7 13 15 2 16 15 15 15 13 13 2
17 10 9 12 0 0 9 4 13 11 11 1 9 1 9 7 9 2
27 14 7 4 15 14 13 1 9 1 9 13 9 2 9 2 16 15 4 7 13 0 9 1 0 0 9 2
11 9 15 14 13 0 2 7 13 10 9 2
18 13 1 9 0 15 9 7 1 9 0 9 2 0 1 9 0 9 2
7 1 9 15 9 14 13 2
21 0 0 0 9 2 9 2 4 1 0 9 13 0 9 2 16 4 13 9 9 2
20 14 13 1 0 9 16 1 9 0 9 2 7 14 13 1 0 9 10 11 2
28 13 2 16 0 0 9 2 3 16 4 13 11 2 14 4 13 1 15 2 16 4 9 14 3 13 0 9 2
22 1 11 15 3 13 0 0 11 2 9 7 10 9 1 0 2 3 13 1 9 11 2
9 10 3 14 0 9 13 3 14 8
9 2 3 15 13 14 3 1 9 2
37 9 11 1 11 2 16 4 13 0 1 9 10 9 2 15 4 1 15 13 2 16 4 9 1 11 13 12 0 9 1 0 2 0 7 0 9 2
45 9 9 0 9 7 9 1 0 9 13 1 15 2 16 15 9 1 15 3 13 3 3 2 16 13 1 9 1 0 9 2 14 7 16 13 10 9 2 0 2 3 1 0 9 2
28 9 9 2 16 15 13 1 0 9 2 15 13 2 16 1 9 0 9 13 3 2 16 13 15 3 3 0 2
30 9 1 9 1 9 1 9 9 14 4 9 13 1 9 0 2 9 2 0 9 2 3 7 13 9 9 1 9 9 2
12 9 7 9 2 0 9 13 1 9 0 9 2
12 0 9 7 9 13 14 15 2 15 9 13 2
24 9 14 13 0 0 9 2 9 7 14 15 13 2 16 1 9 14 4 13 0 9 1 9 2
4 9 1 9 2
14 9 0 9 7 9 0 9 1 9 3 13 10 9 2
19 9 13 1 0 9 2 13 15 2 16 13 9 7 9 7 13 1 9 2
20 13 15 1 0 9 1 0 9 7 0 9 2 7 10 9 13 1 0 9 2
13 9 7 9 14 13 10 2 9 2 14 1 9 2
14 9 3 13 0 9 7 0 0 9 1 0 9 9 2
6 9 15 4 3 13 2
30 16 4 15 15 13 7 16 4 15 13 2 16 15 13 10 9 2 4 14 13 15 3 0 1 15 2 15 4 13 2
16 9 13 7 0 9 1 9 0 9 2 16 15 13 1 0 2
19 10 0 2 0 9 13 13 14 3 0 9 2 7 13 3 13 1 9 2
13 7 7 15 13 14 0 2 0 7 0 9 9 2
4 9 13 15 2
7 13 15 2 16 13 9 2
5 9 15 13 3 2
13 9 9 13 13 14 3 0 2 16 13 1 9 2
6 13 1 9 1 9 2
3 9 15 2
8 9 0 9 7 3 0 9 2
18 10 9 13 0 9 7 0 15 13 1 9 2 16 4 13 10 9 2
8 13 15 4 14 1 0 9 2
13 9 7 9 13 3 3 7 1 15 15 3 13 2
5 9 3 14 13 2
13 13 15 1 9 2 16 13 14 9 3 1 9 2
21 0 13 15 9 2 16 15 3 13 2 13 0 9 7 3 0 2 3 0 9 2
22 9 2 16 10 9 13 9 2 16 15 13 0 13 2 15 13 15 3 3 1 9 2
6 13 15 1 10 9 2
14 13 15 2 16 4 1 10 0 9 3 13 10 11 2
10 9 7 9 2 10 9 15 3 13 2
15 1 9 13 9 2 7 16 10 9 13 2 13 9 13 2
11 15 15 3 13 0 2 7 13 1 9 2
7 10 9 13 9 7 9 2
12 0 9 15 3 13 1 0 2 3 0 9 2
23 9 0 9 15 14 13 2 7 13 10 0 9 15 2 16 13 0 2 0 9 10 9 2
10 1 9 13 0 2 14 16 15 13 2
9 14 15 13 9 2 3 9 13 2
14 14 4 14 13 1 9 2 14 16 4 13 1 15 2
22 10 9 15 4 13 9 1 9 16 2 9 1 0 9 2 16 15 13 1 15 2 2
14 16 15 13 1 0 9 2 13 10 9 3 1 9 2
32 13 12 2 16 15 4 1 9 3 13 1 9 2 16 4 13 0 9 7 15 13 1 9 9 2 1 9 4 13 0 2 2
18 10 3 0 9 15 13 0 9 9 2 16 13 13 9 2 9 2 2
20 9 13 1 9 2 9 7 9 15 13 1 0 9 7 15 1 15 3 13 2
15 1 9 1 0 9 13 13 0 9 1 0 9 7 9 2
19 16 7 10 9 3 2 13 2 2 13 9 0 2 0 7 3 0 9 2
11 13 15 3 2 16 15 4 13 1 9 2
23 14 13 3 10 9 2 16 4 15 1 10 9 13 2 16 16 4 13 13 9 0 9 2
22 9 7 9 2 1 9 15 13 10 9 0 7 0 2 3 7 3 13 1 0 9 2
14 1 15 9 9 13 0 13 3 2 16 4 15 13 2
10 15 13 0 2 9 0 9 3 13 2
11 3 15 13 2 7 10 9 13 0 9 2
12 13 0 2 3 15 13 7 3 13 0 9 2
11 14 13 15 9 2 16 4 13 10 9 2
23 10 9 4 13 0 7 0 2 3 0 7 14 4 13 0 9 2 16 16 13 9 3 2
5 0 9 7 9 2
25 9 4 3 13 0 9 9 7 3 13 2 16 15 10 9 9 13 1 0 9 10 9 0 9 2
49 9 4 14 13 0 9 1 9 7 0 0 9 2 16 0 9 1 9 9 1 9 1 9 9 2 16 13 0 9 0 0 9 2 13 7 13 0 9 9 11 9 1 0 9 10 12 9 9 2
5 13 4 1 12 2
23 16 15 14 13 14 9 2 13 9 1 9 9 1 9 7 13 10 9 0 9 1 9 2
7 9 0 4 13 12 9 2
7 9 13 13 0 7 0 2
3 0 9 2
2 0 2
28 16 4 11 13 2 16 0 3 13 0 9 1 9 2 15 14 4 13 0 9 7 1 15 15 4 9 13 2
19 13 2 16 9 0 13 9 2 9 9 1 10 9 14 15 13 1 9 2
2 9 2
16 9 15 1 15 13 2 0 9 7 3 13 3 1 0 9 2
14 9 2 0 9 14 13 13 0 2 7 3 0 9 2
20 10 9 13 2 16 4 0 9 13 9 2 10 4 3 3 13 9 1 11 2
24 3 13 7 13 9 2 16 1 0 9 9 15 3 13 7 14 13 2 16 10 9 14 13 2
22 16 13 9 1 9 2 0 13 2 16 13 0 2 0 2 15 4 0 9 14 13 2
22 13 7 1 0 9 1 10 0 9 2 7 1 9 2 1 0 9 7 1 0 9 2
17 14 10 10 9 3 4 13 0 0 9 1 3 3 0 0 9 2
12 3 1 10 9 14 13 13 1 9 0 9 2
14 3 4 15 14 15 13 2 16 4 13 14 1 0 2
10 1 15 13 7 9 3 14 3 0 2
21 2 13 7 2 16 15 1 0 9 0 9 10 9 13 9 2 1 9 9 2 2
3 1 9 2
26 9 1 0 9 13 0 1 9 7 9 1 0 9 2 16 15 13 1 9 2 9 7 9 0 9 2
39 14 1 0 9 4 1 0 9 7 0 9 13 9 9 7 9 9 9 10 9 9 2 1 15 4 13 14 0 9 11 2 16 4 10 9 8 9 13 2
13 1 0 9 0 9 7 9 9 4 13 0 9 2
2 9 2
3 9 0 2
5 13 14 15 9 2
11 9 9 4 1 9 13 9 1 0 9 2
7 9 4 13 1 9 9 2
15 13 4 14 9 9 9 11 7 9 1 9 7 0 9 2
5 13 9 9 9 2
2 13 2
3 9 0 2
6 13 4 14 12 9 2
44 9 2 16 4 3 13 2 4 13 0 9 9 2 15 9 13 0 2 16 13 1 10 9 13 2 7 7 4 13 15 2 16 13 1 15 2 16 15 9 13 1 0 9 2
5 15 3 14 13 2
5 9 13 3 0 2
8 15 3 13 10 9 1 9 2
19 0 9 1 9 2 1 16 13 2 13 1 0 0 12 9 1 12 9 2
3 9 0 2
15 13 2 16 15 15 13 2 16 16 15 9 13 2 13 2
8 4 7 13 2 3 13 3 2
31 15 13 2 16 13 1 9 1 9 2 16 13 15 14 9 1 9 2 16 4 15 13 2 16 13 0 1 0 0 9 2
26 16 15 13 2 3 13 2 16 14 13 13 10 9 3 2 16 15 14 13 2 16 13 14 15 0 2
24 13 2 16 1 0 9 13 14 3 7 3 0 10 12 9 2 16 4 15 14 13 1 9 2
3 9 0 2
19 12 1 10 0 9 13 3 0 0 7 13 16 13 1 9 9 3 0 2
3 9 0 2
18 3 4 3 15 13 10 9 1 9 9 2 7 15 4 15 3 13 2
3 13 9 2
4 2 12 0 2
4 15 13 3 2
4 13 15 3 2
17 1 9 12 1 0 9 1 12 9 13 9 1 0 9 10 9 2
9 9 13 9 11 11 2 13 9 2
4 15 13 3 2
4 13 15 3 2
16 13 4 1 10 9 2 16 13 2 16 13 0 13 0 9 2
15 14 2 16 13 2 16 13 10 9 1 0 9 9 0 2
44 1 9 15 15 13 0 2 16 4 3 13 1 9 0 9 1 9 1 0 9 2 16 0 9 13 16 9 1 9 0 9 2 1 9 2 16 4 3 3 13 9 1 15 2
16 9 10 9 2 16 15 13 0 9 12 9 2 13 0 9 2
7 7 14 3 4 13 3 2
4 15 13 3 2
4 13 15 3 2
5 13 1 0 9 2
17 13 1 9 9 0 2 0 9 1 9 9 8 11 11 15 13 2
20 13 2 16 4 9 9 11 11 13 1 9 0 9 0 0 9 1 0 9 2
4 15 13 3 2
4 13 15 3 2
4 15 13 3 2
4 13 15 3 2
8 13 1 9 9 1 12 9 2
10 14 3 13 9 9 11 11 2 11 2
4 9 14 13 2
6 9 13 1 12 9 2
4 15 13 3 2
4 13 15 3 2
15 13 2 16 13 9 1 12 9 2 1 9 12 2 0 2
11 13 1 9 1 12 9 2 1 9 12 2
12 9 13 9 1 9 7 9 0 9 0 9 2
3 9 13 2
3 13 9 2
3 9 0 2
7 13 14 15 13 10 9 2
3 1 9 2
12 13 1 9 1 9 1 12 9 9 11 11 2
9 9 9 13 2 9 9 14 13 2
3 13 9 2
7 13 1 9 1 12 9 2
17 1 12 9 3 13 9 1 12 9 9 8 11 11 7 11 11 2
13 9 9 14 13 2 16 13 9 9 1 10 9 2
12 9 3 13 2 7 1 0 9 13 10 9 2
4 9 13 0 2
4 15 13 3 2
4 13 15 3 2
3 9 0 2
3 9 0 2
3 9 0 2
14 16 3 2 16 9 4 9 13 2 13 1 15 13 2
3 13 9 2
40 15 13 16 9 10 9 1 0 9 1 3 0 9 2 16 13 10 9 1 9 10 9 3 7 4 15 14 3 13 1 9 1 15 2 16 4 15 15 13 2
48 3 4 13 1 9 9 2 9 11 11 2 16 15 13 2 0 9 14 13 9 1 9 2 16 0 9 9 11 13 9 9 11 2 16 13 9 7 9 0 9 12 9 9 1 9 0 9 2
3 13 9 2
13 15 4 14 13 3 2 7 4 1 15 13 3 2
11 16 4 3 13 1 11 2 16 13 9 2
5 15 3 3 13 2
13 13 15 4 13 2 16 4 13 9 1 10 9 2
19 1 9 1 15 13 15 0 9 13 4 15 15 1 0 9 1 0 9 2
12 13 15 1 10 9 2 9 2 9 7 9 2
14 15 4 0 9 13 16 0 9 7 15 13 9 9 2
9 1 0 9 3 13 14 1 9 2
11 3 15 13 2 15 4 13 1 0 9 2
4 9 13 0 2
25 1 9 9 0 11 7 0 9 1 0 9 9 13 15 3 0 2 16 4 3 13 1 10 9 2
17 10 9 13 0 9 7 9 1 15 3 13 0 2 14 0 9 2
12 10 9 13 0 14 1 0 9 7 0 9 2
20 9 0 9 13 14 0 9 7 0 9 1 0 0 9 13 7 13 10 9 2
21 1 10 9 13 3 13 14 0 9 2 1 15 9 3 13 0 9 7 0 9 2
6 13 15 4 1 9 2
7 11 4 13 9 1 9 2
24 3 16 13 0 9 1 0 9 0 1 9 9 1 9 2 13 1 15 0 14 9 1 9 2
13 9 1 9 12 9 7 9 0 13 0 9 9 2
13 9 0 9 15 3 13 1 9 7 1 9 0 2
11 9 1 15 13 10 9 0 9 1 9 2
12 2 10 9 13 1 9 9 0 7 0 9 2
21 3 4 15 13 0 9 0 2 0 7 14 0 9 2 16 15 15 15 3 13 2
28 14 9 15 7 13 2 16 13 0 7 0 9 0 7 15 13 3 13 16 0 7 1 0 0 2 0 9 2
31 7 13 0 7 0 9 1 9 7 0 9 14 12 1 0 9 2 16 15 13 13 1 0 9 2 16 14 13 0 9 2
21 9 1 9 3 2 3 7 3 2 13 0 9 2 13 0 9 7 13 9 9 2
17 1 9 1 9 7 9 0 9 15 15 13 14 10 9 7 9 2
22 1 9 0 9 9 13 1 0 9 2 9 2 9 2 16 15 14 13 7 14 13 2
24 15 13 9 2 16 13 1 0 9 3 0 2 1 9 1 0 0 9 7 13 3 0 9 2
11 7 13 9 10 0 9 1 10 0 9 2
21 11 14 13 10 0 7 0 9 1 10 3 0 9 9 2 7 14 13 1 9 2
13 9 14 13 2 10 9 13 1 10 9 3 9 2
8 3 9 13 7 13 10 9 2
16 11 2 4 3 13 2 3 4 13 2 16 4 1 15 13 2
8 9 7 15 13 14 3 3 2
5 11 15 3 13 2
4 2 13 2 2
16 7 15 4 13 1 9 0 9 2 16 15 13 13 1 9 2
17 13 4 2 16 15 13 10 9 2 1 15 15 14 13 3 13 2
11 2 3 7 14 13 1 9 2 15 13 2
8 1 11 2 11 7 1 11 2
9 3 15 13 1 11 7 1 11 2
41 13 15 1 15 2 16 15 14 4 14 13 0 7 0 2 16 15 4 9 1 0 9 13 1 10 9 7 15 13 2 15 13 2 16 4 15 13 0 9 2 2
13 2 13 2 16 4 13 0 9 7 0 9 3 2
10 15 13 1 9 2 0 1 9 9 2
20 13 9 7 1 9 13 14 1 0 0 2 9 2 2 0 1 0 0 9 2
25 11 11 4 1 9 9 0 9 13 2 16 1 0 9 13 10 9 2 16 15 3 13 0 9 2
15 0 13 9 2 0 0 9 2 2 7 13 10 9 0 2
11 1 10 9 15 13 3 0 7 0 9 2
13 3 3 0 9 0 9 7 15 13 1 0 11 2
11 13 16 9 0 9 2 16 15 14 13 2
12 13 16 9 2 16 1 10 11 13 0 9 2
30 0 9 13 3 0 2 3 0 2 0 0 9 7 9 2 16 15 9 3 14 13 2 3 3 13 7 15 14 13 2
16 7 13 10 9 2 10 9 2 10 9 1 3 1 0 9 2
10 2 14 13 15 15 2 2 4 13 2
22 9 4 3 13 2 13 4 2 16 4 13 3 1 9 14 15 7 16 15 14 13 2
38 11 11 2 0 9 1 9 11 11 8 11 2 16 13 0 9 1 9 11 8 11 2 16 13 0 9 1 9 11 8 11 2 13 1 9 0 9 2
27 1 0 0 9 2 1 15 13 9 0 9 2 13 1 0 0 9 2 16 13 1 9 2 0 0 9 2
8 1 12 1 15 13 11 11 2
9 16 10 0 9 1 9 13 3 2
29 10 9 1 12 3 15 0 9 2 16 15 4 9 9 12 0 13 1 11 2 13 1 9 1 12 9 0 11 2
16 11 11 2 12 2 15 4 13 14 16 9 0 9 1 11 2
17 1 10 9 13 0 0 9 9 7 0 9 7 9 2 9 2 2
44 1 0 9 13 9 10 9 14 0 2 0 9 7 9 7 9 2 16 14 3 14 13 9 2 10 15 1 9 3 13 2 7 9 13 2 16 1 0 13 0 9 1 11 2
24 1 9 1 9 1 0 9 2 16 4 13 9 1 0 9 2 4 13 0 0 9 7 9 2
6 9 4 13 0 9 2
17 3 4 15 13 1 9 7 15 3 13 2 16 16 13 9 3 2
6 15 15 15 3 13 2
3 13 15 2
5 14 15 15 13 2
3 13 9 2
8 13 2 3 15 4 3 13 2
9 3 4 3 13 2 15 15 13 2
4 3 13 3 2
37 13 15 1 9 2 16 13 0 14 1 3 2 3 16 13 0 7 0 14 0 9 2 3 15 3 13 1 9 1 9 2 1 0 9 1 9 2
28 9 4 13 1 9 2 9 9 2 16 15 4 13 2 4 13 1 0 9 1 0 9 1 9 1 0 9 2
12 9 7 0 9 3 4 13 10 9 2 11 2
4 9 15 13 2
8 13 15 1 9 7 13 9 2
7 3 3 15 0 9 13 2
14 1 9 13 14 12 9 9 2 3 13 1 9 9 2
7 1 9 13 9 1 9 2
6 13 15 12 1 9 2
14 9 15 13 1 9 2 0 9 7 13 1 10 9 2
9 3 15 4 11 3 13 1 9 2
25 16 4 9 13 9 1 0 9 2 15 4 13 2 16 13 9 11 2 16 4 3 13 1 15 2
24 10 9 15 4 13 9 11 2 0 9 2 16 4 1 9 13 1 11 13 9 1 0 9 2
8 2 3 13 2 2 4 13 2
47 11 2 12 0 9 1 9 0 9 2 3 1 11 11 2 4 13 11 2 16 1 0 9 9 1 0 9 11 1 11 13 9 2 1 15 4 13 11 11 1 9 0 9 7 0 9 2
32 16 9 9 9 1 10 9 13 0 9 0 9 11 9 2 15 12 12 9 4 13 7 13 1 12 0 9 14 1 0 9 2
21 9 4 3 13 2 16 9 13 1 9 2 7 0 9 11 11 4 3 14 13 2
22 3 4 3 10 16 12 9 3 0 9 1 11 1 0 12 9 13 12 9 1 9 2
21 14 0 12 1 12 9 13 9 3 10 0 9 2 7 15 9 1 15 14 13 2
16 1 0 9 10 0 9 4 13 2 16 9 11 11 13 9 2
7 3 13 14 10 0 9 2
19 16 15 2 16 13 1 9 2 15 14 1 15 3 13 10 9 7 9 2
9 14 9 11 15 3 13 3 3 2
16 13 15 10 0 9 2 9 3 2 13 9 1 9 7 9 2
16 10 9 13 0 9 1 9 9 7 15 4 13 13 1 9 2
22 14 7 15 1 10 9 9 14 13 13 1 0 9 7 14 9 13 0 1 0 9 2
35 13 15 0 9 1 0 9 2 16 4 3 3 13 9 1 9 7 9 2 15 13 7 1 0 9 13 1 9 0 9 1 0 9 9 2
14 1 10 9 13 9 2 7 14 4 15 3 13 9 2
41 1 0 9 0 9 2 1 15 4 14 13 14 9 11 11 2 4 13 1 9 2 3 16 13 1 0 9 2 13 14 2 16 13 1 9 14 2 0 2 9 2
19 1 15 13 10 9 3 1 0 9 7 0 9 2 16 15 3 13 0 2
20 1 9 9 7 13 14 1 0 2 0 2 0 7 0 9 2 4 14 13 2
27 0 9 13 1 9 9 0 0 9 3 0 2 0 9 13 1 12 9 1 9 0 9 7 13 0 9 2
31 16 4 15 13 1 12 9 13 0 9 1 10 0 9 16 9 10 0 9 7 10 9 2 4 15 3 13 1 0 9 2
12 11 15 13 3 3 3 2 16 13 3 3 2
12 11 15 4 13 1 9 1 0 9 1 9 2
5 2 3 14 13 2
38 13 7 14 9 3 10 9 1 12 2 16 4 13 1 9 2 15 7 13 1 15 2 16 9 9 14 4 13 9 7 4 1 9 13 13 1 9 2
15 14 3 15 15 4 13 2 16 4 13 9 14 3 12 2
5 13 4 9 9 2
8 13 14 9 2 16 15 13 2
17 10 9 14 3 3 13 10 0 9 2 3 16 1 15 13 9 2
3 13 9 2
27 0 13 2 16 13 13 10 9 2 1 9 7 4 15 13 15 2 7 16 4 15 13 2 16 4 13 2
27 9 4 15 15 13 13 1 9 2 16 16 4 13 15 1 0 2 7 13 2 16 4 15 15 13 13 2
13 3 13 0 2 16 15 15 0 14 4 13 3 2
8 9 11 15 15 13 1 9 2
13 16 4 13 0 12 9 2 4 13 11 11 11 2
8 9 15 4 13 9 9 12 2
8 1 9 4 15 13 1 9 2
15 9 4 13 9 2 16 4 15 13 1 9 1 9 9 2
11 4 13 1 9 2 13 4 1 9 9 2
12 9 4 13 9 3 2 16 4 13 9 3 2
15 13 4 3 0 2 7 0 16 1 9 9 1 0 9 2
23 16 4 13 1 9 2 4 13 10 0 0 9 2 16 4 13 12 1 9 1 0 9 2
11 1 3 4 13 9 13 16 9 1 9 2
18 10 0 9 4 13 0 9 2 16 15 9 14 13 13 1 10 9 2
23 1 10 10 0 0 9 15 15 4 13 2 14 4 15 13 2 16 4 15 3 13 3 2
32 15 4 13 3 2 16 4 13 2 16 15 13 3 14 3 9 2 16 1 3 13 3 3 2 16 16 1 3 13 3 3 2
22 0 9 10 12 9 4 13 10 0 9 1 9 9 9 1 9 11 4 13 3 0 2
16 4 15 14 3 13 2 14 7 4 15 0 9 14 3 13 2
9 13 4 14 15 0 1 15 0 2
16 9 2 16 15 4 13 10 12 9 2 4 13 3 16 0 2
14 7 7 4 9 13 9 1 9 3 1 9 0 9 2
11 1 10 9 4 13 9 1 15 15 0 2
11 15 15 0 1 15 4 13 3 15 0 2
19 0 0 9 15 4 13 1 9 7 1 15 13 0 9 9 1 0 9 2
38 14 15 4 15 13 1 9 2 13 4 9 2 16 4 13 1 0 9 2 10 9 11 2 10 9 2 16 4 15 13 2 9 2 16 4 13 9 2
23 7 4 15 13 15 2 16 15 14 4 13 1 9 2 9 4 15 3 13 10 0 9 2
24 3 3 15 4 13 2 16 16 15 9 13 1 12 2 15 13 1 9 9 16 1 0 9 2
9 14 0 9 9 15 4 3 13 2
18 16 4 13 10 9 2 4 13 13 7 3 0 7 7 13 0 9 2
3 7 15 2
28 13 4 15 9 2 16 4 14 3 3 13 1 10 9 2 14 16 4 15 13 2 16 15 13 1 9 9 2
28 11 2 12 1 9 4 11 2 16 15 13 1 9 0 0 0 9 2 1 0 9 1 9 13 10 12 9 2
39 1 9 4 3 13 2 16 4 9 1 0 9 13 0 9 11 11 2 0 9 9 11 2 16 15 4 0 9 14 13 2 7 15 4 0 13 1 9 2
19 0 9 4 13 1 0 9 9 2 16 4 1 9 1 9 13 0 9 2
26 1 9 1 9 1 11 1 0 9 13 14 12 9 1 0 9 2 0 9 7 13 9 12 1 15 2
25 9 9 0 9 9 4 13 9 1 9 10 0 9 2 16 4 15 13 1 9 0 9 1 9 2
20 9 4 3 13 9 1 9 9 2 4 13 9 9 0 0 9 9 11 11 2
41 0 9 4 3 1 9 0 0 9 13 2 16 15 1 0 9 3 14 13 13 1 9 0 0 9 2 16 15 14 4 13 0 9 7 15 13 1 9 0 9 2
10 0 0 0 9 4 13 0 0 0 9
9 0 11 11 4 0 9 13 9 2
13 9 4 1 9 0 9 13 0 0 9 11 11 2
18 16 4 1 9 13 9 1 0 9 9 2 4 1 9 13 0 9 2
24 7 16 4 2 11 2 1 0 9 3 13 9 0 9 2 4 13 0 2 16 4 11 13 2
16 10 9 4 10 9 3 13 14 11 2 16 4 13 9 9 2
15 9 9 11 11 13 0 1 0 9 9 9 1 10 9 2
18 16 15 4 13 9 1 9 2 4 3 13 14 1 9 1 0 11 2
33 15 3 13 9 2 15 4 15 9 13 1 9 0 9 2 11 11 11 2 9 2 9 7 9 2 3 14 14 13 3 0 9 2
12 9 13 0 14 1 0 9 2 9 11 11 2
24 2 13 3 0 2 16 14 13 9 1 10 9 2 2 4 11 13 9 7 3 13 1 9 2
8 2 9 15 4 13 10 9 2
19 13 1 9 7 13 1 9 2 15 7 4 3 13 13 10 0 9 2 2
11 1 0 11 10 9 1 9 13 12 9 2
21 11 4 0 9 11 13 1 9 1 0 9 2 16 15 4 1 15 13 0 9 2
6 3 3 15 4 13 2
22 10 9 2 11 7 11 2 4 15 3 13 2 3 16 4 15 1 15 14 3 13 2
27 16 4 13 13 2 15 1 15 15 4 13 0 9 2 4 15 13 1 14 12 9 9 1 9 1 9 2
12 9 13 15 3 7 14 0 4 3 13 15 2
10 15 1 9 9 14 13 13 1 9 9
20 0 9 13 2 16 9 11 3 13 3 13 0 0 7 3 3 13 1 11 2
26 3 1 11 11 4 13 10 9 13 11 2 16 3 13 14 7 9 7 9 1 0 9 1 0 0 2
37 14 4 13 0 13 2 16 11 14 3 13 12 0 9 2 1 9 7 4 13 11 7 11 13 13 2 16 13 10 9 14 3 3 0 1 15 2
20 9 0 13 2 16 15 3 1 9 0 9 7 1 9 0 9 9 14 13 2
28 11 4 15 13 14 1 0 9 2 16 15 4 13 1 9 1 10 9 2 0 3 1 0 9 3 2 3 2
10 0 9 10 9 4 13 1 10 9 2
9 1 15 4 13 11 3 9 9 2
14 10 9 1 9 0 9 1 9 1 9 13 14 11 2
41 3 9 4 13 2 3 4 13 9 2 1 15 4 13 10 9 2 7 7 4 15 13 2 16 9 7 9 13 3 0 2 16 4 13 0 9 9 7 0 9 2
16 13 15 7 14 13 0 9 9 1 9 7 9 7 10 9 2
23 1 9 3 13 9 1 0 9 7 14 13 1 15 2 16 14 4 14 15 13 10 9 2
20 11 2 9 9 1 9 11 13 0 2 16 9 1 9 14 13 10 9 9 2
25 7 4 1 9 13 9 2 16 15 4 13 12 9 7 9 2 16 1 0 9 13 0 0 9 2
39 1 9 4 13 2 16 4 15 1 10 9 9 7 9 3 13 10 9 2 16 13 1 9 9 2 7 3 3 13 15 2 16 10 9 0 9 14 13 2
20 1 9 1 0 0 9 7 9 13 2 16 4 10 9 14 3 13 0 9 2
43 10 9 9 2 16 13 9 9 9 9 9 1 9 2 13 9 11 11 2 16 4 0 0 9 2 11 2 13 1 9 2 16 1 9 10 0 9 3 13 9 1 11 2
32 16 4 13 9 1 9 11 11 1 9 0 2 7 4 9 10 9 13 1 12 1 12 2 15 4 3 13 0 9 1 9 2
26 1 9 0 9 11 2 11 1 12 9 13 11 1 11 0 0 0 9 2 1 15 3 13 13 9 2
21 14 7 13 0 13 1 0 9 7 2 16 4 15 13 1 0 2 13 0 9 2
26 9 11 4 15 14 1 9 13 2 16 14 13 13 10 9 9 2 9 11 1 11 13 0 0 9 2
6 3 4 13 9 11 2
17 2 0 0 9 2 11 2 4 13 9 9 1 0 9 0 9 2
14 0 9 15 4 3 13 1 0 11 2 12 9 2 2
39 3 4 13 1 10 9 0 11 11 11 2 16 4 1 0 9 1 9 1 12 9 13 9 0 9 9 7 16 0 9 1 9 0 13 0 0 9 9 2
13 1 10 0 0 9 4 3 13 9 1 0 9 2
17 1 0 9 15 4 9 7 9 13 1 0 9 2 1 0 9 2
9 15 4 15 13 1 10 0 9 2
9 3 4 13 9 1 9 7 9 2
23 7 3 4 3 13 7 4 13 13 1 9 1 9 2 3 16 15 4 15 13 1 9 2
6 9 13 1 9 9 2
10 9 9 1 0 9 13 9 9 9 2
17 7 3 15 13 2 16 4 9 13 9 2 16 15 3 14 13 2
19 14 13 14 3 2 16 13 9 3 13 9 1 0 9 2 9 3 13 2
20 15 0 15 4 13 0 9 2 16 4 9 13 10 9 1 3 12 0 9 2
17 2 1 9 7 4 13 0 9 2 7 15 0 0 9 4 13 2
3 3 13 2
15 9 4 13 13 0 9 1 10 0 9 1 9 0 9 2
15 1 10 9 13 1 9 1 0 9 0 9 9 0 9 2
19 2 16 13 12 9 9 2 13 1 11 15 0 10 0 9 7 0 9 2
45 1 10 9 2 1 9 0 9 14 4 13 14 1 0 9 2 14 4 13 10 9 2 16 1 10 9 13 0 9 0 9 2 16 13 9 9 2 9 1 9 9 7 9 9 2
27 9 14 4 15 13 1 9 2 16 15 10 9 3 3 13 1 9 0 9 7 7 16 9 13 0 9 2
34 16 15 4 13 9 9 11 2 4 15 1 10 0 9 13 2 16 4 3 12 9 9 0 0 9 1 0 12 9 13 1 0 9 2
26 13 4 14 9 0 0 9 2 16 4 13 11 2 16 13 3 3 2 2 16 4 13 1 10 9 2
13 11 11 2 9 0 9 2 1 10 9 13 3 2
23 0 0 2 0 2 0 2 0 7 0 9 13 0 2 0 2 0 2 0 7 0 9 2
21 9 13 3 0 13 7 10 16 12 0 9 7 0 9 2 16 15 14 3 13 2
27 9 13 0 1 9 12 0 0 9 11 11 11 2 10 9 13 1 0 14 9 0 9 9 7 0 9 2
21 9 4 0 9 13 0 9 2 16 13 1 9 3 15 2 16 15 13 1 9 2
8 9 4 13 14 11 11 11 2
21 11 2 11 2 16 4 11 11 13 1 9 1 0 11 2 4 13 9 1 11 2
17 7 3 1 9 4 13 2 6 2 15 0 15 4 13 1 9 2
9 13 15 4 2 16 4 13 9 2
14 13 4 2 16 4 13 0 2 16 15 4 0 13 2
20 16 4 13 3 7 14 15 9 2 14 14 4 13 15 3 2 15 4 13 2
10 11 2 13 3 1 9 11 1 9 2
19 16 13 13 9 3 0 2 13 13 0 2 0 7 3 13 13 1 9 2
11 16 7 13 15 2 13 11 3 1 15 2
10 10 9 7 10 9 4 13 1 15 2
4 15 0 9 2
16 11 2 3 13 2 15 4 13 1 10 9 1 10 0 9 2
4 4 15 13 2
4 4 13 15 2
13 13 15 4 1 15 16 1 10 9 1 0 9 2
17 11 2 11 2 14 10 9 4 15 3 13 1 9 1 0 9 2
10 11 11 4 1 10 9 13 3 0 2
23 9 4 13 2 16 15 13 13 3 1 15 7 16 13 3 13 9 2 16 4 15 13 2
37 10 9 4 3 13 2 16 13 10 9 7 9 1 0 9 1 9 0 9 3 0 10 9 2 9 7 4 13 13 0 1 0 9 14 1 9 2
29 9 4 3 13 2 16 0 9 14 13 13 2 15 3 13 9 1 0 0 9 7 15 13 1 0 9 0 9 2
10 9 4 13 14 9 0 0 0 9 2
15 10 9 0 9 4 13 0 1 0 9 2 0 1 9 2
23 9 4 13 0 1 12 9 2 1 15 16 4 13 0 12 9 3 1 12 1 12 9 2
25 9 4 13 0 9 1 10 9 1 0 9 1 9 9 2 9 10 9 7 9 0 2 0 9 2
20 9 13 14 0 9 1 9 9 7 9 2 3 3 7 13 0 14 0 9 2
17 0 9 0 7 0 9 13 9 2 9 2 7 9 2 9 2 2
13 15 13 9 0 7 0 16 0 9 0 0 9 2
16 1 0 9 13 7 0 7 0 9 0 9 1 0 0 9 2
17 11 15 4 13 1 9 9 2 16 13 10 9 7 15 3 13 2
39 14 4 13 11 0 1 9 2 16 9 1 9 1 0 9 7 1 0 9 1 10 9 13 0 9 1 9 7 3 13 0 9 7 9 1 10 0 9 2
3 1 12 2
21 9 11 13 2 16 9 7 9 9 1 9 0 9 7 1 9 0 9 13 9 2
24 1 0 0 9 9 7 9 9 13 9 2 16 9 2 0 9 7 0 9 9 14 13 3 2
12 11 13 14 1 9 7 9 1 9 9 11 2
21 1 0 9 7 13 14 2 16 0 9 2 16 15 13 2 13 1 9 3 0 2
6 9 9 13 14 12 2
39 9 2 1 15 4 13 1 9 9 0 7 0 9 0 0 0 9 1 9 0 9 2 13 9 1 9 1 0 0 0 9 1 12 9 1 9 9 9 2
20 16 9 13 1 9 2 9 1 15 14 13 13 10 9 2 16 14 13 9 2
26 0 9 1 9 1 10 9 15 3 14 13 13 16 0 7 1 15 14 13 13 0 0 9 9 0 9
24 16 9 0 0 9 4 9 1 9 13 14 1 3 0 9 2 7 15 1 0 9 4 13 2
20 0 9 1 9 9 1 9 15 3 13 1 9 3 0 9 9 1 0 9 2
24 16 9 1 9 15 13 9 9 1 9 9 7 1 9 1 10 9 2 7 1 0 9 9 2
41 2 1 9 2 16 13 12 9 0 9 2 16 0 9 9 7 9 1 9 1 9 2 16 15 13 0 9 2 7 1 0 9 14 13 2 16 3 13 0 9 2
3 1 12 2
10 9 11 3 13 14 9 9 1 9 2
19 13 2 16 9 1 9 11 3 9 0 9 3 13 9 1 9 1 9 2
15 0 9 13 0 3 2 16 9 13 9 7 16 13 9 2
14 16 9 1 9 13 9 2 13 0 0 9 12 9 2
26 2 1 9 9 9 0 9 9 1 9 2 16 15 13 9 7 9 1 9 2 13 13 1 0 9 2
15 9 9 0 9 13 3 13 2 16 13 14 12 9 9 2
35 16 4 15 13 9 9 11 2 9 9 7 9 9 2 0 9 2 2 13 0 9 7 9 2 16 15 0 9 13 13 1 9 9 9 2
15 9 1 9 9 13 0 9 7 9 0 0 9 1 11 2
29 0 2 3 0 9 9 1 0 9 4 13 9 7 9 9 9 2 15 3 1 0 9 15 9 13 1 9 9 2
21 9 0 9 7 9 13 1 11 0 1 0 9 2 9 9 1 0 9 7 9 2
27 1 12 9 11 15 9 0 9 1 0 0 9 2 16 13 0 1 9 12 11 2 13 3 1 9 12 2
10 0 7 0 9 9 13 0 3 3 2
7 9 15 13 1 0 9 2
16 1 9 9 13 0 9 1 9 2 16 15 9 13 1 9 2
36 9 13 9 0 9 13 1 0 9 2 3 14 3 2 1 10 9 15 0 9 13 9 3 2 7 3 1 9 0 9 1 0 0 9 2 2
34 0 9 9 1 9 13 9 1 9 9 9 7 9 1 10 0 9 3 1 9 7 9 9 1 9 2 16 13 0 1 0 0 9 2
30 11 13 0 2 0 0 9 0 0 9 9 7 9 1 9 2 16 4 13 3 0 9 1 9 1 9 1 9 12 2
25 11 13 9 7 9 9 7 9 1 9 1 0 7 0 9 7 9 1 9 9 7 9 1 9 2
13 11 13 14 9 2 0 1 9 7 9 1 9 2
33 11 13 9 1 9 16 0 9 10 0 9 2 16 13 1 9 1 9 7 9 1 0 9 0 9 7 1 9 9 1 0 9 2
20 9 13 9 9 1 9 7 9 1 0 9 0 9 2 16 9 14 13 3 2
27 1 9 1 9 7 9 1 0 9 13 0 0 9 1 0 9 1 9 2 16 4 0 9 13 9 9 2
24 10 0 9 1 9 0 9 4 15 13 2 15 4 1 9 13 14 0 9 7 0 0 9 2
56 1 15 3 3 13 1 0 10 9 0 9 9 2 16 9 14 14 4 13 2 7 4 15 3 14 13 2 16 4 13 1 0 9 3 9 0 7 0 0 2 0 9 1 3 0 7 0 9 1 9 2 15 13 3 12 2
22 11 2 9 15 10 9 13 2 9 9 7 9 7 13 2 3 3 13 15 0 13 2
27 0 9 9 13 10 9 2 9 7 13 2 3 15 13 13 0 9 7 3 13 9 12 9 1 15 0 2
18 1 11 13 1 12 9 0 7 0 9 2 16 15 15 1 0 13 2
11 13 13 3 14 9 12 9 9 7 9 2
26 1 10 9 13 1 0 9 2 3 15 13 3 13 1 12 9 7 15 1 12 9 13 1 10 9 2
16 1 0 9 14 13 13 14 2 16 13 1 9 1 0 9 2
28 1 9 1 9 13 9 3 13 1 9 7 9 2 14 7 1 9 2 16 13 9 0 9 7 7 14 9 2
12 1 9 0 9 7 14 14 13 0 13 9 2
21 3 4 13 1 9 2 16 15 4 14 3 13 7 15 4 3 13 1 0 9 2
24 1 0 9 4 13 1 9 0 9 0 14 1 10 9 2 16 15 4 0 9 13 1 9 2
17 1 9 4 15 0 2 0 13 1 10 9 7 11 13 9 9 2
29 3 0 9 0 1 9 4 9 13 1 0 9 2 14 1 12 9 4 0 11 11 13 1 9 1 9 0 9 2
23 0 9 9 4 11 1 9 11 1 0 9 7 0 9 1 9 11 13 1 9 1 12 2
11 4 13 0 13 0 9 14 3 0 9 2
20 3 4 13 0 0 9 11 11 2 16 4 13 0 9 11 14 1 0 9 2
14 13 4 1 0 9 9 9 2 16 15 4 3 13 2
8 1 9 9 4 13 1 9 2
13 9 1 9 0 9 4 0 9 13 1 9 9 2
13 1 10 9 4 9 1 0 9 13 10 9 3 2
18 3 4 1 9 13 0 0 9 1 0 9 9 7 0 9 1 9 2
9 10 9 4 13 1 9 0 9 2
16 1 10 0 9 4 0 9 13 9 1 0 0 9 1 0 2
6 9 11 4 13 9 2
19 9 13 0 1 0 9 9 11 2 16 15 4 9 1 0 9 14 13 2
17 1 0 9 7 1 0 9 4 0 9 1 11 3 13 14 15 2
7 9 15 13 1 12 9 2
6 1 9 13 0 9 2
10 1 9 9 15 13 9 9 1 9 2
12 1 11 4 15 3 0 2 13 2 14 0 9
21 1 11 13 14 1 0 0 9 0 2 16 4 14 3 3 13 0 9 11 11 2
36 13 7 13 14 2 16 15 4 11 1 11 14 13 2 16 14 4 1 0 0 9 13 11 11 2 16 15 4 15 2 13 2 1 0 9 2
36 11 2 12 2 3 4 13 0 0 9 0 9 0 0 7 9 9 9 0 9 7 1 0 9 11 2 14 0 9 4 13 14 0 0 9 2
14 16 14 9 13 1 0 9 2 15 4 13 3 13 2
25 9 4 1 0 9 3 13 10 9 2 2 3 7 4 13 2 16 13 0 1 3 0 9 2 2
33 11 2 12 2 0 9 11 11 2 4 7 13 2 16 14 4 13 13 9 9 2 7 13 9 1 9 11 11 1 9 0 9 2
34 9 15 4 13 13 3 11 0 2 16 4 13 1 9 2 16 14 13 13 2 9 2 9 1 0 9 2 16 10 9 13 1 11 2
31 10 0 9 1 9 1 9 7 15 4 13 1 0 9 2 7 4 13 9 1 9 7 9 9 1 0 0 9 0 9 2
21 0 9 13 10 9 1 9 2 16 4 13 0 9 1 9 9 7 10 0 9 2
21 0 9 2 16 13 10 0 9 2 7 13 2 3 13 0 2 0 9 1 9 2
30 1 10 14 0 9 1 9 0 9 1 9 3 13 1 9 7 9 9 7 13 14 10 0 9 1 9 9 7 9 2
13 3 3 7 15 4 9 13 11 11 11 1 11 2
25 13 15 2 16 13 0 9 3 0 1 9 2 9 2 2 16 15 4 13 11 11 2 12 2 2
21 0 7 0 0 2 0 9 9 1 9 7 0 0 9 13 1 12 9 10 9 2
41 0 9 13 1 0 9 1 15 2 0 2 1 3 0 2 0 2 3 0 15 7 0 2 9 2 9 7 9 2 3 1 9 2 9 2 9 2 9 7 9 2
20 2 9 1 0 9 14 13 13 1 0 9 2 13 13 1 0 9 7 9 2
40 9 2 16 1 9 13 1 9 0 9 2 3 13 9 2 16 4 13 0 7 0 0 0 2 2 13 9 9 0 9 9 2 16 4 13 0 9 7 9 2
23 15 2 1 15 13 1 9 1 9 7 9 2 13 9 9 1 9 7 9 7 1 15 2
33 13 0 9 2 1 15 15 13 9 9 2 7 7 13 0 9 1 3 0 7 3 0 9 2 16 15 13 9 9 7 0 9 2
16 13 2 16 13 9 7 9 10 9 0 9 0 16 10 9 2
45 15 13 0 9 1 9 1 9 7 9 1 15 1 15 2 16 4 1 9 14 3 3 13 1 10 9 2 16 7 13 9 0 9 1 0 0 9 7 10 9 1 0 9 9 2
41 1 9 10 9 0 9 4 13 0 0 9 1 0 9 1 9 0 0 9 1 0 0 7 3 1 9 0 0 1 9 1 9 2 0 2 0 9 0 9 2 2
46 10 2 0 2 9 1 11 7 0 0 9 4 13 9 0 9 1 9 0 9 2 16 4 15 13 3 3 1 9 9 0 9 1 10 9 0 9 1 0 9 1 0 9 1 9 2
28 0 9 0 9 4 1 9 7 15 0 13 10 9 2 16 7 15 4 0 9 0 0 7 0 3 3 13 2
24 0 9 2 16 4 3 13 1 0 9 11 3 14 1 10 9 2 4 1 10 9 13 9 2
34 9 0 9 11 11 13 2 16 13 3 9 1 10 9 7 9 1 15 2 15 4 3 10 9 13 7 10 9 4 13 1 0 9 2
45 3 4 13 0 2 16 13 1 9 2 7 4 9 13 1 0 0 9 2 16 4 13 0 9 2 16 4 13 2 16 4 8 8 13 12 9 9 2 12 9 9 7 10 9 2
39 1 9 4 13 2 16 4 9 7 9 13 14 1 9 0 9 1 12 2 0 8 8 1 11 2 16 15 4 1 10 9 13 1 9 3 12 9 9 2
23 14 10 9 4 15 9 13 1 9 9 2 16 4 15 13 2 16 4 14 13 1 9 2
13 9 0 4 13 2 16 4 13 0 1 0 9 2
9 3 0 9 7 13 1 9 11 2
16 11 11 13 2 16 4 11 11 13 13 2 16 13 14 0 9
25 9 1 9 1 11 4 1 0 9 13 1 0 9 2 9 7 15 4 3 13 3 12 0 9 2
19 1 0 9 9 15 4 13 9 9 7 9 1 0 2 0 7 0 9 2
32 0 9 0 9 1 0 9 13 1 12 2 16 15 4 13 9 9 11 7 9 9 2 16 15 0 9 13 1 0 9 11 2
34 3 4 1 9 7 9 1 0 9 13 0 9 7 0 9 2 1 2 9 2 0 9 9 7 4 13 9 14 9 9 7 0 9 2
14 3 4 13 2 16 4 1 0 9 0 13 1 9 2
9 7 15 4 14 13 15 1 15 2
13 3 15 4 1 9 13 9 2 7 4 13 9 2
18 11 2 12 2 0 9 11 11 4 3 13 1 0 0 9 1 11 2
17 1 0 9 15 4 1 0 9 13 9 2 9 0 9 11 11 2
31 9 4 13 1 9 0 9 2 3 7 15 4 13 3 2 16 4 11 13 14 9 9 11 11 7 9 0 9 11 11 2
25 13 1 0 0 9 0 9 1 11 7 3 0 0 0 0 9 1 9 1 9 0 9 0 9 2
10 0 9 4 3 13 14 9 0 9 2
13 13 4 15 11 11 1 11 7 11 11 1 11 2
7 15 15 15 13 1 9 2
10 13 2 16 15 15 13 10 9 9 2
18 7 9 15 3 13 15 2 15 15 15 13 2 16 1 9 3 13 2
28 1 0 9 13 3 16 1 9 2 10 9 2 9 7 0 9 13 0 13 15 2 14 16 3 14 13 9 2
19 11 11 1 10 9 8 8 8 8 8 2 10 9 3 13 0 2 13 2
14 13 15 9 1 0 9 9 2 16 15 13 1 9 2
8 16 15 15 13 2 15 13 2
29 3 13 14 1 10 9 16 9 1 9 0 9 9 2 16 13 0 7 0 9 16 0 9 1 0 7 0 9 2
35 1 9 11 4 14 13 0 9 2 1 15 4 9 13 9 0 9 2 13 7 15 4 0 9 1 9 9 1 0 9 2 9 7 9 2
17 0 9 13 9 9 1 9 7 9 1 0 0 9 4 13 0 9
31 11 2 1 0 0 9 7 9 4 3 13 12 2 9 11 7 12 2 9 9 0 9 1 11 2 15 9 13 14 0 2
36 0 9 0 7 0 9 7 9 4 13 2 16 13 9 10 9 9 2 14 3 1 9 2 1 15 4 15 13 9 9 7 0 9 0 9 2
2 8 8
4 9 13 0 2
53 3 16 4 0 9 11 11 1 10 9 1 11 3 3 13 9 12 9 11 2 15 4 13 13 2 16 10 9 9 2 16 15 15 4 13 1 9 9 7 9 9 9 11 2 14 13 3 1 9 0 0 9 2
37 10 9 3 4 13 9 0 9 1 11 7 16 15 1 10 9 1 15 13 0 9 1 0 9 2 4 9 1 0 9 9 1 9 3 13 9 2
32 11 4 13 2 16 13 14 0 0 13 9 10 9 7 13 9 1 12 9 9 2 14 16 14 4 14 3 13 1 0 9 2
20 14 0 9 10 9 13 1 9 2 0 9 7 13 1 15 13 3 0 9 2
18 9 0 13 1 0 9 2 1 0 9 2 0 2 0 7 3 0 2
4 9 0 9 2
8 0 0 9 7 9 11 9 2
3 0 9 2
29 3 4 9 0 9 11 13 2 16 4 11 13 10 16 12 9 9 0 9 2 16 4 10 0 9 13 12 9 2
28 10 9 4 3 13 2 16 15 4 0 9 13 9 2 16 4 13 0 1 9 7 1 15 4 13 9 9 2
38 11 2 12 0 0 9 11 11 4 3 1 9 1 11 13 0 9 1 0 0 9 0 0 9 1 9 11 2 16 15 3 13 1 9 11 7 11 2
14 7 15 15 13 1 0 2 16 14 13 9 0 9 2
18 9 7 15 3 13 1 9 2 10 11 11 13 14 14 1 9 2 2
24 9 7 9 9 11 4 7 3 13 9 9 1 0 7 0 11 1 9 11 9 1 0 11 2
35 1 9 2 16 13 14 9 0 9 2 0 1 9 2 0 9 2 9 9 7 9 2 4 3 13 14 1 11 2 11 2 11 7 11 2
14 14 14 13 10 9 2 9 11 2 15 4 13 11 2
6 3 12 9 3 13 2
13 11 4 13 1 9 9 2 16 15 4 15 13 2
12 2 13 0 7 0 9 2 16 13 13 9 2
15 9 1 9 13 3 3 2 16 15 13 0 9 1 9 2
7 13 7 3 15 3 13 2
13 7 13 3 0 2 16 13 9 1 0 9 0 2
12 13 2 16 1 9 9 1 9 14 13 3 2
14 14 7 15 4 1 9 1 9 1 9 14 3 13 2
10 0 13 2 16 4 10 9 14 13 2
28 3 7 3 3 1 9 2 0 0 0 9 13 9 9 0 0 9 2 7 13 10 0 9 1 0 0 9 2
16 13 4 1 15 1 9 7 15 13 3 1 0 9 1 9 2
10 13 15 4 7 13 1 15 1 9 2
24 1 9 15 9 3 13 2 16 3 14 13 14 13 9 2 16 15 13 0 9 1 10 9 2
18 9 11 11 13 3 0 9 2 7 4 15 13 3 13 9 0 9 2
22 14 14 2 16 14 13 14 1 0 0 9 13 14 12 9 2 10 9 13 3 0 2
15 1 9 13 3 0 11 11 2 16 1 9 13 0 11 2
29 14 7 2 16 13 0 9 9 2 16 16 13 0 0 9 1 9 2 1 15 3 11 1 9 1 11 13 9 2
30 7 9 2 16 15 13 0 9 2 16 1 9 1 0 9 13 0 9 0 9 2 16 15 13 1 0 9 2 13 2
19 1 0 0 9 15 1 0 9 1 11 1 9 1 11 3 13 12 9 2
8 9 0 9 7 10 9 13 2
30 0 9 13 0 2 3 0 9 2 9 2 9 2 1 9 0 9 1 9 7 9 7 0 9 7 15 3 3 13 2
26 13 0 9 2 15 13 1 9 7 9 7 13 1 9 1 0 9 2 1 15 9 13 14 1 9 2
13 13 1 9 0 0 9 7 13 1 9 3 9 2
31 0 9 13 1 9 7 13 1 9 2 16 15 13 1 0 9 2 0 0 0 9 2 9 7 10 9 7 13 1 0 9
31 9 4 3 13 1 11 9 2 15 13 1 0 9 9 7 14 3 1 15 1 0 9 13 12 2 0 8 8 1 11 2
13 11 4 3 13 7 1 15 13 9 1 9 9 2
17 14 4 15 13 9 2 1 0 9 7 15 4 13 1 0 9 2
3 2 8 2
28 11 11 4 13 1 12 1 0 9 11 11 1 11 2 12 2 2 0 7 4 13 11 11 11 2 12 2 2
20 0 9 7 9 11 11 4 1 9 13 12 2 7 4 13 10 9 1 12 2
15 1 12 9 4 13 0 0 9 11 11 2 11 1 12 2
15 0 9 1 12 9 1 9 4 13 11 11 1 0 12 2
22 11 2 12 14 1 9 4 12 9 1 11 1 0 11 1 9 13 9 7 15 13 2
27 12 2 7 0 9 4 12 2 0 0 9 1 9 1 12 12 9 13 1 9 7 15 1 9 13 9 2
39 10 9 2 0 9 7 9 1 0 0 9 9 7 9 9 2 16 15 13 14 0 9 11 11 2 15 3 13 1 14 3 0 7 0 0 9 8 11 2
10 0 9 13 1 3 3 3 16 8 8
9 3 15 4 13 1 9 1 9 2
29 15 1 9 1 9 14 13 9 13 3 2 3 2 2 7 1 10 9 7 9 9 3 4 3 3 13 7 13 2
22 14 4 9 1 10 9 13 7 15 3 1 0 9 14 1 2 13 3 0 0 9 2
14 3 3 1 15 13 14 9 1 9 10 3 0 9 2
35 1 0 9 9 9 13 14 1 0 9 2 16 13 2 2 0 2 9 2 9 1 2 9 2 2 7 4 14 9 10 9 13 0 9 2
7 0 13 0 9 10 9 2
12 9 2 9 13 8 13 1 10 9 1 9 9
28 1 9 0 9 2 16 15 13 9 2 13 1 0 9 11 1 11 2 16 4 3 13 12 9 9 1 9 2
56 1 15 13 1 9 0 12 14 12 9 1 9 2 3 16 13 1 0 9 2 16 13 9 1 3 0 2 1 9 3 12 9 1 9 2 1 0 7 13 11 2 11 2 1 0 11 2 16 13 3 0 14 12 9 9 2
21 1 0 9 12 9 15 13 9 2 1 9 2 1 15 4 13 1 0 9 2 2
9 13 1 9 1 9 0 9 9 2
18 13 0 2 3 0 9 1 9 9 1 9 11 11 11 11 11 11 2
42 10 0 9 2 16 13 9 9 2 3 13 0 7 0 9 7 13 0 9 1 9 2 13 0 14 0 9 2 16 3 1 9 13 9 1 9 7 13 9 1 15 2
26 9 11 11 11 11 2 16 15 13 1 9 2 13 0 1 10 9 9 2 16 15 13 1 9 9 2
45 16 13 13 9 11 11 2 13 1 12 1 12 9 1 12 7 12 9 0 1 9 11 1 9 11 7 1 11 2 1 0 9 2 0 11 2 11 7 11 7 1 0 9 11 2
6 1 10 9 13 0 2
12 3 13 2 16 13 0 2 7 15 13 15 2
21 13 7 1 9 7 3 13 2 7 16 1 9 3 14 14 13 2 15 4 13 2
7 14 10 9 7 13 0 2
25 1 12 9 15 14 3 15 9 13 1 10 9 2 9 15 9 14 1 10 9 13 3 3 13 2
18 9 13 1 9 10 9 14 1 12 9 7 3 13 3 1 0 9 2
16 1 9 0 9 13 1 10 0 9 12 9 9 2 16 13 2
19 3 0 9 2 9 2 2 16 13 9 2 13 3 0 7 3 13 9 2
26 1 10 9 13 14 0 9 2 16 13 10 0 9 2 16 3 13 1 9 2 1 9 9 0 9 2
24 16 13 10 9 0 2 13 14 3 0 2 16 13 9 2 7 4 15 0 9 13 13 13 2
14 16 13 13 9 2 13 3 13 7 13 9 1 9 2
20 16 13 9 2 15 1 15 13 1 9 2 14 7 13 13 7 13 0 9 2
13 9 15 14 13 2 7 15 15 3 14 14 13 2
15 3 13 2 1 9 7 4 13 14 10 9 1 0 9 2
9 2 14 4 15 3 13 1 9 2
21 16 4 3 9 13 7 13 9 1 9 2 14 13 2 3 4 13 3 15 3 2
38 16 15 13 2 16 4 15 1 9 3 13 2 15 13 0 15 7 1 9 2 3 13 9 7 13 9 2 1 15 15 13 14 9 1 9 1 9 2
19 13 13 1 0 9 1 9 9 2 16 13 2 16 9 13 9 7 9 2
9 15 13 10 0 0 7 0 9 2
12 9 4 13 3 2 1 9 4 14 3 13 2
22 2 14 13 2 3 15 4 13 3 3 13 9 1 9 2 7 4 1 9 13 9 2
25 1 9 2 16 15 13 10 0 9 2 4 13 3 0 2 3 7 4 13 15 1 9 3 0 2
11 1 9 12 14 4 13 10 9 9 1 9
18 9 9 0 9 4 13 2 16 4 15 9 0 13 1 3 12 9 2
24 1 15 4 13 0 12 9 2 9 9 9 7 14 14 4 13 12 9 0 9 1 0 9 2
17 3 1 0 9 7 13 9 0 2 4 13 1 11 7 0 9 2
18 0 9 1 9 1 10 9 4 10 9 13 14 9 1 9 11 11 2
18 1 0 9 11 11 15 4 13 10 16 12 0 9 1 9 7 9 2
7 1 9 4 13 3 0 2
15 14 0 9 4 13 15 2 16 15 15 14 14 13 13 2
9 1 9 4 13 10 16 12 9 2
17 3 4 13 10 9 7 10 9 7 13 3 3 10 9 1 9 2
13 11 4 13 2 16 13 11 10 9 14 1 15 2
16 11 4 13 1 15 7 13 2 16 13 1 0 9 15 3 2
27 11 11 2 3 2 4 1 0 9 13 9 9 1 11 7 3 13 1 0 0 9 1 9 12 1 11 2
9 2 9 2 11 11 11 15 4 13
34 9 4 13 1 15 2 16 4 1 12 9 1 9 11 9 1 0 9 11 11 13 2 11 7 15 4 13 1 0 9 10 9 11 2
19 1 12 9 4 0 9 13 9 2 16 4 1 9 1 9 13 1 12 2
33 1 12 9 7 4 11 13 0 9 1 0 9 9 11 2 13 9 1 0 9 2 16 4 13 1 9 0 11 7 13 0 9 2
25 11 2 12 2 3 16 1 15 1 9 4 13 14 1 11 3 0 9 1 0 9 1 0 9 2
10 11 4 13 9 0 9 11 1 9 11
15 14 15 4 9 13 1 0 2 0 9 7 1 0 9 2
19 15 4 13 3 14 3 0 9 9 1 0 9 2 7 0 9 4 13 2
13 0 9 4 3 13 11 2 0 7 4 3 13 2
16 2 3 15 13 14 1 9 2 7 13 1 0 9 14 0 2
24 15 4 13 0 9 7 13 2 16 15 14 1 0 14 4 13 2 2 4 13 1 9 11 2
31 3 15 13 14 9 2 13 7 16 0 9 9 2 16 15 3 13 3 7 1 9 1 0 9 9 2 9 7 1 9 2
13 0 13 2 16 9 3 13 1 9 9 16 9 2
24 1 15 13 9 2 9 9 2 16 9 1 9 3 13 2 7 13 1 12 7 12 9 9 2
29 9 0 9 4 13 3 3 0 2 7 4 15 0 7 1 9 0 9 7 0 9 3 1 9 13 1 9 9 2
27 14 0 9 1 9 4 11 13 0 9 2 1 15 4 13 9 7 9 2 15 4 3 13 1 0 9 2
23 0 0 9 2 16 13 3 0 1 0 0 9 1 11 2 7 13 1 12 0 1 11 2
20 14 1 0 9 4 13 0 9 2 16 4 13 3 12 1 12 9 0 9 2
24 1 9 4 15 13 1 0 9 2 7 16 9 12 2 16 4 13 9 2 4 13 1 9 2
48 9 7 0 9 11 14 10 9 13 0 9 7 14 9 1 9 0 7 0 9 2 16 13 0 9 2 16 4 13 10 12 2 0 9 9 14 3 2 16 4 13 0 1 12 7 3 9 2
17 7 14 0 9 3 3 15 13 2 7 13 9 0 13 1 15 2
42 14 4 7 13 0 2 16 4 1 9 13 1 9 10 0 9 7 4 13 14 10 10 0 9 7 3 1 11 14 4 13 14 0 9 2 16 13 0 1 9 9 2
2 8 11
9 7 15 4 13 1 3 0 9 2
3 0 9 2
18 9 1 9 9 7 13 2 16 0 0 9 14 13 9 1 9 9 2
28 1 11 4 13 13 14 9 2 16 4 11 2 16 11 14 13 0 9 2 11 13 2 16 16 13 1 9 2
21 1 15 13 0 9 0 7 4 13 1 9 9 1 11 9 1 9 9 10 9 2
15 11 11 2 1 0 9 3 0 9 13 12 0 0 9 2
17 9 13 2 16 0 9 2 9 7 0 9 14 13 1 0 0 9
17 11 11 2 9 15 0 2 13 9 2 16 14 13 9 1 0 9
5 9 4 13 0 2
9 7 10 9 4 13 13 10 9 2
6 9 4 13 10 9 2
10 0 9 0 9 4 13 13 1 12 9
43 1 10 9 2 3 16 4 13 1 9 0 9 2 7 15 13 13 2 16 4 13 9 1 9 11 7 0 11 2 1 15 13 0 2 16 13 3 2 16 13 3 0 2
19 11 2 12 16 4 14 13 2 4 0 9 13 9 0 9 11 7 11 2
23 9 4 9 1 9 9 13 1 9 2 16 1 9 9 9 0 9 13 0 13 0 9 2
18 3 7 15 4 13 14 0 9 2 16 4 9 3 13 1 0 9 2
35 9 4 13 13 9 9 2 3 7 13 14 0 2 16 4 3 3 13 9 1 0 9 7 9 9 11 1 11 2 1 15 13 0 9 2
24 3 4 13 9 0 9 9 1 0 9 9 8 11 1 11 2 9 4 13 9 0 11 2 2
30 0 4 13 9 9 1 9 2 1 9 0 9 2 3 7 4 14 13 0 0 9 8 11 1 9 1 11 1 11 2
25 16 13 11 11 2 14 4 3 13 1 10 9 0 0 9 7 9 1 9 9 7 3 13 9 2
27 9 12 4 15 13 9 7 9 10 9 1 11 2 3 7 13 1 0 9 2 16 14 4 10 9 13 2
25 13 15 2 16 9 1 3 0 9 7 1 10 9 14 13 14 0 2 7 13 14 3 14 0 2
33 13 7 13 2 16 15 9 13 2 4 13 10 9 1 0 9 12 1 9 11 11 11 2 16 4 15 13 14 0 9 10 9 2
26 15 1 15 9 13 0 9 1 9 2 16 14 4 15 15 0 13 2 3 7 15 1 15 14 13 2
30 9 4 13 9 0 9 8 11 8 11 2 16 4 0 13 2 16 1 12 9 1 9 14 13 12 9 1 0 9 2
25 1 9 4 3 1 9 13 12 9 9 0 9 2 0 9 9 7 13 1 9 12 9 0 9 2
19 0 9 2 16 4 13 1 9 9 2 0 9 2 4 13 1 0 9 2
28 1 0 9 1 11 4 13 1 9 2 12 9 3 2 0 1 12 0 9 2 16 13 9 11 8 7 11 8
7 10 9 13 15 10 9 2
9 1 9 4 13 12 0 9 13 2
49 16 1 10 9 13 14 12 9 2 16 4 9 1 9 13 2 13 9 2 16 4 13 1 0 0 9 1 9 10 16 12 9 15 2 16 4 3 7 3 2 7 14 3 13 14 0 9 9 2
23 9 9 13 3 0 9 7 7 15 14 13 2 10 4 13 9 9 1 0 9 1 15 2
13 7 0 16 0 7 0 9 4 15 13 1 9 2
9 1 15 9 14 13 13 10 9 2
9 10 9 4 13 14 3 2 13 2
21 3 4 13 1 9 2 16 4 15 13 13 1 9 9 2 4 1 9 9 13 2
15 1 11 15 14 13 7 1 9 12 7 1 9 0 9 2
8 7 3 15 13 0 9 9 2
7 3 4 15 13 9 9 2
19 3 16 4 3 1 11 9 0 9 1 0 13 2 7 1 11 13 3 2
24 15 13 14 3 1 9 1 12 0 9 2 7 1 9 9 9 9 4 15 13 1 9 9 2
3 11 11 2
17 2 13 4 10 0 9 2 7 16 15 13 14 1 12 0 13 2
8 13 7 1 9 0 0 9 2
13 13 4 14 12 9 9 1 12 9 0 0 9 2
25 0 9 4 13 1 0 9 0 9 11 7 3 1 9 1 9 13 0 9 2 10 9 7 9 2
53 3 4 3 0 0 9 0 0 9 2 16 10 9 0 0 9 13 14 14 1 9 9 7 9 2 14 14 9 2 9 2 13 3 0 9 2 14 3 13 0 15 2 13 7 4 13 3 3 0 1 10 9 2
8 16 16 9 13 9 10 9 2
19 0 9 11 1 0 9 1 0 9 4 3 14 13 16 9 9 1 0 2
12 0 9 2 9 10 9 2 15 0 4 13 2
17 10 9 1 4 0 9 1 9 0 9 1 9 3 13 9 9 2
30 0 9 13 13 2 16 3 0 9 12 1 12 2 16 4 1 9 13 3 2 4 13 1 9 14 1 0 9 9 2
32 15 4 3 16 4 9 1 0 9 9 13 13 14 11 2 16 13 14 1 9 2 16 13 9 15 1 9 13 2 3 13 2
10 14 2 14 0 9 4 13 3 0 2
8 14 15 4 15 3 3 13 2
11 1 15 1 0 9 1 11 4 13 9 2
26 3 13 11 0 13 0 9 2 16 13 1 0 0 9 2 3 16 13 0 7 0 9 1 10 9 2
14 15 13 2 16 3 13 0 9 1 9 1 0 9 2
12 9 13 13 1 9 2 16 13 0 9 9 2
7 14 9 9 3 13 9 2
18 9 4 13 3 0 2 16 4 14 13 13 15 0 2 0 2 0 2
19 14 16 4 3 3 13 2 4 13 9 2 16 15 4 13 3 1 9 2
13 13 15 4 14 3 2 7 15 4 13 3 3 2
23 13 4 3 3 2 3 2 3 2 3 7 4 13 3 3 0 7 0 16 10 0 9 2
13 0 9 4 1 11 13 9 2 0 1 0 9 2
13 13 4 15 9 1 0 9 2 1 3 0 9 2
13 3 4 15 13 1 9 7 15 13 1 0 9 2
8 15 12 4 3 13 15 9 2
17 16 15 4 13 3 1 9 2 15 4 11 13 0 9 0 9 2
15 11 4 13 3 3 3 1 9 2 16 15 4 3 13 2
5 7 13 15 4 2
5 16 0 0 9 2
13 9 4 13 3 0 2 16 4 1 15 13 9 2
10 2 13 2 15 4 13 0 9 2 2
16 2 6 2 15 13 7 0 9 2 2 15 4 3 13 11 2
20 2 15 13 14 0 9 2 16 15 9 3 13 3 1 15 7 13 1 9 2
11 1 9 14 13 0 2 0 2 0 9 2
21 1 15 15 3 13 1 0 9 9 0 0 9 2 1 9 12 2 1 0 9 2
16 2 1 11 4 13 0 12 0 9 7 9 11 11 2 2 2
22 10 9 7 14 1 9 15 3 13 0 0 9 2 16 13 3 0 1 0 0 9 2
9 2 1 0 9 13 10 9 9 2
4 13 3 3 2
9 15 7 3 13 0 1 11 2 2
7 3 4 13 14 3 3 2
10 3 15 4 13 1 9 0 0 9 2
7 3 4 0 9 14 13 2
12 13 4 2 16 13 14 3 1 0 1 9 2
27 3 13 4 2 3 15 13 9 7 3 1 9 13 2 16 13 15 14 10 9 2 1 15 4 11 13 2
28 11 13 7 14 3 1 0 1 9 1 9 7 9 7 15 15 3 13 2 16 4 13 1 9 0 0 9 2
61 10 9 13 10 0 9 2 16 15 3 14 13 7 9 1 0 9 9 7 9 1 0 0 9 2 9 0 0 9 1 0 9 1 9 12 9 12 7 13 14 3 13 3 2 16 4 15 13 13 1 10 9 2 16 4 13 1 9 0 9 2
17 0 9 4 15 3 13 1 0 0 9 7 1 9 13 0 9 2
19 9 11 8 13 0 1 10 12 9 9 2 0 9 7 9 9 14 13 2
3 2 8 2
21 0 8 8 7 4 9 13 1 0 9 2 16 4 1 9 13 1 0 0 9 2
32 0 11 2 12 2 1 9 1 12 9 15 4 1 9 11 1 11 1 11 13 0 0 9 2 1 15 4 13 9 0 9 2
21 1 10 3 0 9 7 4 1 9 13 3 3 0 1 3 0 2 11 9 2 2
31 3 0 1 2 11 9 2 14 14 13 0 9 7 0 9 2 7 7 3 13 0 9 7 13 15 0 13 1 0 9 2
19 10 0 9 1 9 9 3 2 13 2 1 12 9 2 1 12 9 2 2
27 3 0 0 9 4 9 0 9 1 9 1 11 3 13 1 0 12 9 9 2 12 9 9 2 1 9 2
42 11 2 12 2 0 9 1 9 1 0 9 4 1 0 9 2 15 4 15 14 13 2 1 9 2 2 13 14 0 9 1 9 2 16 13 1 10 9 0 0 9 2
37 1 14 0 9 14 14 13 0 0 9 2 1 15 13 13 10 9 1 0 9 2 1 15 2 16 13 1 10 9 2 7 13 0 9 14 0 2
26 9 4 9 13 1 9 9 1 9 7 9 2 16 4 14 13 0 9 1 9 1 9 1 9 0 2
12 9 1 12 9 15 4 13 1 0 0 9 2
23 1 0 9 4 15 11 11 2 3 2 7 10 9 11 11 13 1 9 0 9 1 11 2
12 1 0 0 9 1 11 11 4 13 14 0 9
13 1 16 13 9 1 9 2 15 13 10 0 9 2
23 7 13 2 16 13 9 14 0 9 2 0 7 13 15 2 15 15 4 13 1 3 9 2
22 11 11 2 3 4 13 2 3 9 3 3 13 2 16 13 9 1 9 9 7 9 2
18 9 8 11 11 1 0 9 11 11 1 11 11 4 13 9 1 15 2
13 3 4 11 11 1 3 0 6 13 1 11 11 2
8 15 0 15 4 13 1 9 2
15 14 16 4 13 1 9 2 4 11 13 2 3 4 13 2
12 15 4 13 0 9 2 16 4 13 16 6 2
13 13 4 9 7 13 11 11 1 0 2 0 9 2
24 1 11 11 4 13 0 9 14 1 9 2 16 4 15 16 9 13 1 10 9 1 9 11 2
11 3 4 13 2 14 16 4 15 13 9 2
16 15 4 15 13 3 3 1 9 7 4 3 13 1 11 11 2
6 11 4 13 1 9 2
15 1 10 0 7 0 9 4 15 3 15 13 1 0 9 2
23 3 4 13 2 16 4 1 11 11 13 9 2 16 4 15 3 3 13 7 3 3 13 2
15 11 4 13 0 12 9 2 13 4 9 9 7 14 0 2
10 10 9 4 13 0 2 16 4 13 2
6 14 9 4 14 13 2
16 1 9 1 12 4 13 0 1 9 2 0 1 9 1 11 2
16 13 4 1 9 11 11 2 16 4 13 3 1 9 11 11 2
13 3 4 13 1 0 7 0 9 9 10 0 9 2
30 1 10 9 4 13 2 16 13 1 9 2 1 15 7 15 4 13 1 15 1 9 13 2 16 4 15 1 15 13 2
6 7 15 4 13 0 2
5 14 0 4 13 2
35 3 15 4 13 2 3 4 13 0 9 3 0 1 10 9 7 4 14 14 13 15 13 1 9 2 16 15 4 3 13 1 1 0 11 2
10 11 11 15 4 13 1 9 7 13 2
8 0 4 13 2 16 13 0 2
32 0 9 2 16 15 4 13 0 9 1 9 2 15 4 13 1 0 9 2 16 15 4 13 13 2 16 15 4 14 3 13 2
8 11 4 13 14 14 12 9 2
22 3 4 13 7 14 13 2 7 15 4 13 2 1 15 4 13 2 16 13 0 9 2
8 11 15 15 4 3 13 0 2
12 13 4 1 9 1 9 7 15 3 13 9 2
8 16 3 4 13 0 1 9 2
6 0 0 0 0 9 2
6 0 9 1 0 9 2
9 2 3 4 13 0 2 0 9 2
5 13 4 1 9 2
5 13 4 12 3 2
3 13 4 2
4 3 4 13 2
19 13 4 2 16 4 13 1 11 7 1 0 9 2 16 4 13 0 9 2
10 13 15 4 2 16 4 15 3 13 2
17 2 0 9 3 13 1 0 9 9 0 9 2 2 4 13 11 2
8 13 4 15 16 9 1 9 2
8 11 4 13 0 1 0 9 2
18 9 2 16 15 4 13 9 2 9 2 0 0 9 2 0 0 9 2
6 13 15 4 3 0 2
5 3 4 3 13 2
5 15 4 15 13 2
13 2 13 15 4 9 2 2 4 11 13 1 15 2
15 9 14 4 13 0 2 16 14 4 13 12 1 10 9 2
8 9 1 9 15 15 4 13 2
14 2 0 13 3 13 10 0 9 2 2 4 13 11 2
5 3 4 15 13 2
8 3 7 4 13 1 0 9 2
4 3 0 9 2
3 3 0 2
16 13 10 9 2 2 4 13 11 2 16 4 15 13 1 15 2
6 3 4 13 3 3 2
9 2 10 9 13 2 2 4 13 2
5 11 4 15 13 2
10 1 0 9 9 4 1 9 13 9 2
13 2 14 2 15 13 15 2 16 4 13 13 3 2
9 14 4 15 13 13 3 3 15 2
2 13 2
12 1 0 2 0 9 4 13 13 1 0 9 2
21 14 4 13 13 16 3 0 9 3 3 2 7 10 9 4 13 0 7 3 0 2
5 3 13 15 11 2
6 3 13 3 15 11 2
10 16 13 3 2 15 9 15 13 3 2
11 11 4 13 13 9 9 2 7 4 13 2
15 1 9 9 4 13 13 2 3 4 3 13 0 0 9 2
14 13 4 15 14 13 1 9 2 16 4 13 15 0 2
11 2 15 4 13 3 0 9 1 12 9 2
7 11 4 15 3 14 13 2
19 13 15 0 1 10 9 9 2 2 4 13 2 16 4 13 1 0 9 2
15 13 1 0 0 9 4 13 2 16 16 4 13 1 9 2
25 0 9 4 13 0 1 9 7 9 2 16 15 4 3 2 16 4 13 1 11 2 13 1 9 2
15 9 4 13 0 1 0 9 9 7 1 0 9 0 9 2
24 9 2 16 4 15 13 2 7 15 14 2 16 4 15 13 1 9 2 4 15 14 3 13 2
10 1 9 15 15 4 13 9 0 9 2
7 2 3 13 0 10 9 2
21 13 4 1 9 2 7 14 16 4 13 1 9 2 4 14 13 12 9 1 9 2
18 1 0 9 4 3 13 9 1 9 2 3 4 14 3 13 1 15 2
13 1 15 0 4 3 13 7 9 4 13 1 9 2
5 9 4 13 13 2
7 9 4 15 13 1 9 2
5 10 9 4 13 2
12 14 4 3 13 2 16 13 15 14 3 0 2
7 2 11 13 14 1 9 2
7 3 4 13 1 10 9 2
10 1 0 9 1 11 4 13 12 9 2
3 10 9 2
3 10 9 2
3 10 9 2
8 3 4 13 3 0 16 15 2
15 2 15 15 13 16 0 0 15 9 2 2 4 13 11 2
15 11 15 4 13 2 16 3 16 15 0 13 10 0 9 2
12 15 4 13 3 9 2 16 13 1 0 9 2
17 1 9 4 13 2 16 4 11 11 13 11 11 1 9 11 11 2
13 11 4 13 0 12 11 11 7 3 4 13 0 2
8 13 0 9 2 11 7 11 2
12 7 14 11 4 13 0 13 10 9 10 9 2
15 13 15 4 10 0 9 7 15 3 4 13 13 9 15 2
18 15 4 13 10 0 9 16 4 13 3 0 2 3 3 0 4 13 2
21 0 2 0 9 1 15 2 16 13 0 9 9 7 13 0 9 2 4 13 0 2
7 10 9 4 13 14 0 2
14 9 9 4 1 9 9 9 11 11 11 1 9 13 2
21 1 15 13 1 9 9 1 11 2 16 15 4 1 0 13 9 1 0 9 11 2
48 10 9 11 1 0 9 7 1 0 9 4 13 1 0 9 1 9 9 9 1 0 9 9 2 0 1 9 2 16 4 13 0 1 0 9 9 1 10 0 9 1 9 1 12 1 12 9 2
23 0 9 1 10 9 13 1 9 2 1 9 1 9 12 2 1 9 12 0 9 1 9 2
19 11 2 1 9 4 9 1 11 13 2 15 4 13 13 9 1 0 9 2
17 13 4 7 1 0 9 1 9 2 13 2 12 9 7 14 9 2
26 16 15 4 13 13 2 15 4 13 9 7 9 4 3 1 0 13 12 2 0 8 8 7 9 13 2
3 9 13 2
2 8 8
26 11 2 1 11 4 1 0 9 9 1 0 13 10 9 2 1 15 7 15 9 4 15 13 3 13 2
15 9 4 3 13 15 1 10 9 2 16 4 14 14 13 2
36 9 2 16 4 13 1 9 1 0 11 2 4 13 10 9 2 16 15 4 13 1 9 2 7 16 15 4 3 13 2 13 14 12 9 0 2
7 9 4 13 1 12 9 2
20 0 9 13 0 9 1 9 7 9 7 13 1 9 0 7 0 9 1 9 2
22 16 13 3 1 9 13 0 0 9 2 13 15 14 3 3 0 2 13 11 7 11 2
12 2 0 9 4 13 0 9 7 13 0 9 2
16 11 7 11 4 13 12 15 2 16 4 13 0 1 9 9 2
16 1 15 4 13 0 1 10 0 2 0 2 0 7 0 9 2
12 8 8 8 8 8 2 0 9 1 0 9 2
25 9 0 9 2 1 12 1 12 9 11 2 12 2 13 9 2 16 13 0 0 9 10 9 9 2
34 0 9 13 9 2 0 1 9 2 1 15 9 13 0 1 0 7 0 0 7 0 9 2 13 7 15 1 0 9 1 9 9 9 2
11 0 9 13 0 13 14 1 9 0 9 2
39 1 0 9 13 3 0 2 16 13 9 0 9 0 1 9 0 9 2 15 3 13 2 16 13 9 0 9 1 9 0 9 1 9 11 2 12 3 0 2
12 1 0 9 13 0 9 1 0 9 10 9 2
26 15 13 1 9 2 16 1 10 14 9 2 0 9 7 15 1 9 1 0 9 2 14 13 10 9 2
24 16 7 11 2 12 14 13 14 9 9 2 12 9 2 2 13 9 1 0 7 0 9 0 2
23 9 10 9 1 9 13 2 16 9 9 13 2 9 1 12 0 9 7 13 9 9 9 2
19 13 9 2 16 4 9 13 9 2 1 15 15 1 9 14 13 0 9 2
34 0 4 13 2 16 13 1 0 11 0 9 1 9 9 1 9 1 0 9 2 1 9 9 9 7 1 9 1 0 9 1 9 12 2
13 15 4 13 9 1 9 9 1 9 1 0 9 2
22 7 4 13 0 9 13 0 9 1 9 2 16 4 13 0 1 9 9 9 0 9 2
39 9 4 13 13 1 0 2 16 15 4 0 9 3 13 9 1 9 7 16 0 9 2 16 15 9 13 1 0 9 1 9 2 14 13 10 0 0 9 2
51 9 4 13 1 9 9 1 9 0 1 9 0 9 2 16 13 0 9 2 1 15 15 4 9 13 0 9 1 9 2 0 3 1 10 0 9 2 9 7 15 4 14 3 3 13 1 9 0 0 9 2
30 1 10 9 9 9 4 13 0 13 9 2 7 4 13 9 2 1 15 4 13 1 9 0 13 2 16 9 15 13 2
33 10 9 13 0 9 0 9 12 9 11 2 1 0 9 2 16 11 13 2 16 13 9 3 13 0 9 1 9 2 9 7 9 2
28 0 9 2 0 9 0 9 13 9 1 0 9 1 0 11 2 12 9 2 2 16 13 1 9 2 12 9 2
6 9 9 13 12 9 2
14 13 7 15 3 1 9 12 2 12 7 12 2 12 2
10 9 4 13 9 11 11 7 11 11 2
16 9 1 0 9 9 7 13 1 9 0 9 3 14 3 0 2
16 10 9 0 9 4 13 13 9 2 3 4 14 13 13 9 2
17 3 14 4 13 2 16 4 13 1 9 2 15 13 10 0 9 2
24 10 10 9 4 15 7 13 2 16 13 10 0 9 9 2 16 15 15 4 13 1 0 9 2
19 0 13 2 16 4 15 9 9 2 15 9 13 2 13 14 1 9 9 2
31 11 11 2 12 1 9 0 9 1 0 11 2 4 13 14 2 16 13 11 14 3 3 2 16 15 3 14 13 13 11 2
39 16 13 9 10 0 9 10 14 0 2 0 7 0 9 2 3 3 13 2 16 4 13 9 12 10 11 3 2 16 15 4 3 1 10 9 13 13 11 2
17 7 15 14 3 14 13 2 16 4 1 11 1 0 9 13 11 2
9 3 13 14 9 7 13 14 9 2
12 9 13 14 2 1 10 9 1 9 13 3 2
4 14 4 13 2
14 13 4 2 16 15 4 1 9 13 13 14 16 9 2
5 7 0 9 13 2
18 11 7 0 0 9 0 9 10 9 13 0 9 2 9 7 9 9 2
6 0 13 10 12 9 2
7 9 14 13 1 0 9 2
24 1 10 9 4 1 9 11 13 10 12 9 2 9 9 13 0 3 7 12 9 13 3 0 2
18 13 10 9 1 9 7 9 13 2 16 13 10 9 2 13 9 2 2
7 15 15 7 11 3 13 2
11 15 4 13 0 9 9 7 0 0 9 2
7 13 2 16 13 1 9 2
18 9 15 13 1 9 2 16 3 13 0 9 1 0 0 9 7 9 2
24 9 1 0 7 0 9 13 1 11 10 0 9 1 14 3 0 2 7 13 1 3 0 9 2
8 13 4 9 11 11 1 11 2
14 13 2 16 4 13 10 9 2 16 4 13 1 11 2
20 11 4 3 13 2 16 4 13 11 11 14 3 0 7 0 1 10 0 9 2
4 4 15 13 2
6 15 13 9 2 14 2
5 3 4 15 13 2
8 13 15 2 9 1 9 2 2
15 0 9 13 2 16 0 9 14 14 13 2 16 15 13 2
12 1 0 9 4 15 13 0 2 16 0 9 2
13 14 7 15 1 10 10 9 13 2 16 13 0 2
13 11 7 4 1 10 9 1 15 13 1 0 9 2
17 14 1 0 9 10 9 13 11 0 9 0 9 2 9 7 9 2
18 9 9 2 16 13 15 2 3 13 9 2 16 15 1 0 14 13 2
10 3 10 0 9 9 13 1 9 9 2
20 2 11 3 3 13 3 2 16 15 3 13 2 15 13 2 2 4 13 11 2
11 2 13 1 15 7 13 15 4 15 15 2
13 11 4 13 1 11 2 15 7 4 13 1 9 2
6 2 1 9 4 13 2
5 15 4 13 15 2
17 13 4 2 16 4 15 13 1 11 7 3 13 10 9 1 0 2
7 2 6 2 3 15 13 2
10 14 3 4 3 13 10 9 1 15 2
8 2 15 15 4 13 3 0 2
17 1 0 9 15 14 3 13 0 9 2 7 10 9 13 9 9 2
21 9 13 9 0 9 7 9 2 7 14 13 15 2 16 13 0 0 9 7 9 2
16 9 14 13 1 15 2 16 13 3 0 9 7 9 1 9 2
18 14 7 13 9 2 16 12 2 12 9 9 1 9 14 14 13 13 2
20 2 11 4 13 3 0 9 2 1 15 13 3 0 2 3 4 13 0 9 2
13 1 9 11 15 9 4 13 13 1 0 0 9 2
10 3 15 14 1 9 14 13 3 13 2
21 9 0 9 11 13 1 0 9 3 0 2 7 7 0 9 1 15 13 0 9 2
15 13 7 9 7 7 0 9 7 0 0 9 1 0 11 2
13 2 1 9 13 0 14 9 2 7 3 13 9 2
6 15 13 10 0 9 2
19 0 9 2 11 7 11 13 9 7 16 13 1 9 9 2 13 9 0 9
18 3 13 1 15 15 2 3 13 0 1 15 2 16 13 15 0 9 2
7 7 15 13 14 0 9 2
9 3 2 16 13 0 2 13 9 2
16 15 3 14 13 13 2 9 13 2 16 1 10 9 13 0 2
6 14 3 4 3 13 2
3 3 13 2
13 0 9 14 4 13 9 9 1 10 11 7 9 2
9 1 0 11 4 15 13 9 9 2
21 10 9 4 1 15 13 1 11 2 16 15 0 4 13 13 1 10 0 0 9 2
37 9 13 0 14 1 9 2 16 16 3 13 9 7 16 15 13 3 3 2 3 16 16 3 15 15 13 1 0 9 2 16 15 15 10 9 13 2
6 7 1 9 13 3 2
23 14 16 13 9 1 9 9 1 9 0 9 0 2 15 13 2 16 15 7 14 4 13 2
19 13 15 4 7 9 2 16 4 13 2 16 4 13 9 9 1 9 0 2
13 1 9 13 9 2 10 13 9 1 9 0 9 2
13 9 13 0 2 16 15 9 13 0 1 10 9 2
14 0 13 0 2 0 9 1 9 9 7 0 0 9 2
23 3 15 4 1 9 9 2 0 9 11 11 7 9 0 0 9 11 11 2 13 1 9 2
22 2 15 4 3 13 2 4 13 3 0 2 16 4 1 9 13 1 10 9 0 9 2
13 2 13 4 15 9 1 9 7 15 13 0 9 2
15 2 1 15 4 3 13 1 0 9 7 13 0 0 9 2
20 10 12 9 3 4 1 15 13 9 2 16 4 15 9 13 14 1 12 9 2
15 15 4 13 1 9 2 16 4 13 15 0 1 0 9 2
27 0 9 4 13 0 10 12 9 2 3 7 15 4 13 1 3 10 16 12 9 0 7 12 9 0 9 2
43 9 4 15 13 2 16 4 10 9 13 1 9 1 9 14 3 12 9 2 16 4 1 15 13 10 9 7 9 2 1 15 4 13 7 16 4 15 9 0 9 13 15 2
6 4 13 13 10 9 2
17 14 13 1 0 0 9 0 10 9 2 16 7 13 1 9 0 2
20 0 9 14 9 13 3 2 16 14 13 14 13 2 9 7 1 15 13 0 2
16 14 2 14 11 4 3 1 9 0 9 3 3 13 10 9 2
43 0 11 2 16 4 13 3 9 9 11 1 0 2 0 9 2 4 13 1 15 11 2 7 14 13 4 1 0 9 1 9 2 16 15 13 1 11 2 14 13 9 3 2
9 11 7 13 14 0 9 1 15 2
8 7 14 15 4 3 13 11 2
16 14 0 13 1 15 2 16 15 9 7 0 9 15 14 13 2
12 13 14 10 9 2 16 1 9 13 15 0 2
34 1 9 10 9 4 1 9 0 0 9 7 0 9 9 1 0 0 9 13 0 9 9 9 7 9 1 9 0 9 1 9 0 9 2
18 13 2 16 4 11 10 9 7 9 3 13 7 15 1 10 9 13 2
29 1 9 13 2 16 0 9 9 13 0 9 1 9 2 1 15 4 15 13 0 9 1 9 9 9 1 0 9 2
38 15 4 13 1 15 0 9 2 7 13 4 4 2 16 15 0 9 14 13 15 13 2 16 1 0 14 13 1 15 2 15 15 15 4 13 3 0 2
21 0 13 2 16 4 15 13 2 16 4 14 3 13 1 15 2 1 15 13 15 2
25 3 7 13 10 9 10 9 2 16 13 15 0 16 0 9 2 15 7 15 14 13 13 1 0 2
19 2 7 4 13 3 0 2 16 4 13 2 16 3 13 1 3 0 9 2
15 1 10 9 4 1 10 9 9 13 2 1 10 9 13 2
30 13 9 9 7 13 2 3 4 15 13 9 2 3 4 13 1 9 7 3 15 3 13 2 16 4 13 15 1 9 2
30 13 2 16 15 13 15 0 7 16 13 14 15 2 16 4 14 15 13 13 0 9 2 16 15 4 0 13 1 9 2
14 13 15 13 2 16 13 0 13 9 0 1 10 9 2
27 14 15 13 0 2 16 15 14 13 15 2 16 15 13 3 2 16 4 15 14 3 13 2 16 14 13 2
23 14 13 13 0 2 16 4 15 13 1 15 2 7 13 15 4 3 2 16 13 15 15 2
18 16 4 13 1 9 2 3 7 1 0 9 2 4 15 14 13 9 2
13 3 4 15 13 2 15 15 13 9 1 10 9 2
5 14 15 4 13 2
7 3 4 3 13 10 9 2
14 13 2 16 3 14 13 9 7 9 1 9 9 3 2
12 9 15 4 13 2 16 0 9 15 14 13 2
25 10 9 13 1 15 0 9 2 7 16 1 9 2 16 15 14 13 9 1 9 2 13 0 9 2
22 9 9 4 3 13 9 2 16 4 15 2 16 14 4 13 0 9 2 3 13 9 2
35 10 9 14 4 13 1 9 14 0 9 2 7 1 12 9 14 4 13 14 12 2 16 4 15 13 3 2 16 15 1 9 13 9 9 2
21 3 13 9 2 16 15 14 13 3 13 2 15 16 13 13 1 9 1 10 9 2
14 10 9 15 13 14 9 2 16 15 4 14 3 13 2
9 13 15 4 2 16 15 14 13 2
31 14 10 9 4 13 3 2 7 4 14 13 2 16 13 3 1 10 9 10 9 1 0 9 16 1 10 0 9 1 9 2
6 9 4 13 3 0 2
21 9 4 13 1 9 1 0 9 2 16 4 13 10 9 1 9 1 0 9 9 2
26 13 15 4 2 16 13 9 14 14 0 2 7 14 3 0 13 10 0 9 2 16 4 13 3 9 2
11 7 4 13 2 15 15 13 13 10 9 2
19 13 4 7 15 13 13 1 9 2 16 4 13 3 0 1 9 0 9 2
17 1 10 9 15 15 4 13 2 16 4 13 1 15 15 14 15 2
5 13 4 0 9 2
38 1 9 2 16 4 15 0 13 2 4 15 1 0 9 13 2 7 16 4 15 13 13 1 0 9 2 16 4 15 13 1 9 1 0 9 10 9 2
7 13 4 13 9 1 9 2
11 3 4 15 13 1 10 9 7 1 9 2
24 3 2 16 4 15 13 1 0 9 2 4 15 1 0 9 1 0 15 13 2 16 4 13 2
4 3 13 0 2
21 11 4 3 13 9 1 0 9 2 1 9 7 13 3 13 14 9 1 0 9 2
20 11 4 14 13 2 16 4 13 0 9 1 9 11 7 1 0 7 0 9 2
22 11 13 1 0 9 9 9 2 7 15 13 9 2 10 13 9 11 1 10 0 9 2
14 11 13 13 9 2 16 4 15 13 2 7 4 13 2
3 2 9 2
14 0 9 4 13 1 9 1 0 9 1 0 2 0 9
10 10 9 1 9 0 9 1 11 1 11
10 10 9 4 13 1 0 9 1 9 2
9 4 15 13 10 9 1 10 9 2
7 11 4 3 13 1 9 2
10 9 1 9 4 13 9 16 11 11 2
12 1 9 0 0 9 11 4 13 12 0 9 2
13 1 0 9 13 0 11 11 14 10 9 1 9 2
24 11 4 13 1 11 3 1 0 11 2 11 11 1 11 2 0 11 1 11 7 0 11 11 2
22 10 9 1 9 13 11 2 7 13 9 1 9 11 2 11 2 7 11 2 11 2 2
16 1 15 4 1 11 13 14 0 11 7 11 11 2 11 2 2
46 1 0 9 4 1 9 0 9 3 13 11 2 16 1 9 1 10 9 4 13 14 11 2 13 15 4 1 11 2 7 0 11 2 16 15 4 1 9 1 9 3 13 14 1 9 2
21 1 0 9 4 7 14 0 1 9 13 1 15 2 16 14 14 4 13 10 9 2
18 7 1 3 0 9 4 15 3 13 7 1 9 14 13 1 0 9 2
16 1 0 9 0 0 9 4 1 11 10 12 9 13 2 0 2
16 9 13 16 9 9 7 9 9 0 7 1 0 16 1 9 2
22 0 13 3 14 2 16 13 10 9 1 9 2 16 13 1 10 9 7 9 0 9 2
10 1 15 15 4 13 10 0 0 9 2
11 3 13 2 7 13 1 9 7 1 15 2
8 13 9 2 7 13 1 9 2
7 0 9 1 9 13 3 2
12 1 9 9 13 9 7 1 10 9 13 9 2
16 9 2 16 15 13 1 11 2 13 0 2 13 9 7 9 2
9 13 15 1 9 1 0 0 9 2
10 0 11 2 9 2 13 0 0 9 2
14 0 4 13 1 12 9 1 11 2 0 11 1 11 2
6 13 9 9 7 9 2
14 13 0 2 13 1 9 7 9 7 13 9 1 9 2
23 10 0 9 15 4 14 13 2 14 9 9 7 4 13 0 9 0 9 1 9 1 9 2
15 9 13 7 14 12 0 9 2 1 10 9 13 0 9 2
14 9 13 0 9 2 10 9 7 13 3 0 0 9 2
16 9 2 16 15 3 13 9 2 1 0 0 9 13 1 15 2
27 11 11 7 11 11 4 9 12 13 0 0 0 9 1 9 0 9 2 16 15 15 4 3 13 9 9 2
18 9 4 13 13 1 9 1 0 9 2 16 4 13 14 1 9 0 2
31 1 9 12 2 12 2 16 4 13 11 0 9 9 11 11 1 11 7 1 11 2 15 4 10 9 3 13 1 0 9 2
27 10 9 4 13 1 3 0 9 9 1 0 7 0 9 7 3 4 12 13 0 2 9 2 1 12 9 2
19 11 1 3 13 0 9 1 0 9 2 3 16 0 11 13 14 1 9 2
20 9 1 9 13 14 0 7 0 2 7 11 4 9 1 11 15 13 7 13 2
20 14 14 13 9 2 11 11 2 0 1 9 2 16 3 7 3 13 1 9 2
22 1 9 11 2 16 4 13 9 9 2 9 0 9 7 9 9 2 4 15 3 13 2
33 16 4 0 9 13 1 9 11 0 9 3 13 2 15 4 1 9 12 13 1 0 9 11 2 7 1 9 4 13 1 0 9 2
29 0 9 13 3 3 7 15 1 15 13 2 16 4 13 14 1 0 9 0 9 2 1 9 2 9 7 9 9 2
11 0 9 1 9 10 9 1 11 13 0 2
38 9 9 11 13 0 1 9 9 0 9 2 10 9 7 9 1 9 1 11 1 0 9 1 10 9 1 9 9 7 9 1 9 1 3 0 9 9 2
28 1 9 1 15 4 9 13 3 3 9 2 16 4 3 13 1 15 2 16 4 13 9 10 9 7 15 13 2
35 9 0 9 4 15 7 3 3 13 9 2 16 4 15 13 1 10 0 9 7 15 2 16 4 15 13 13 2 13 2 16 14 13 9 2
10 9 4 13 1 9 9 9 7 9 2
11 0 9 1 15 4 15 13 0 12 9 2
33 1 15 4 0 0 3 3 3 13 2 16 15 9 13 1 9 2 0 7 4 13 3 0 9 2 16 13 2 15 1 15 13 2
26 1 10 9 4 14 13 2 16 13 2 16 0 1 0 9 9 13 0 7 16 15 15 13 10 9 2
32 7 4 1 15 1 9 1 9 13 3 0 7 4 1 9 13 14 15 2 16 14 4 13 2 16 4 11 13 1 10 9 2
21 3 4 1 9 14 13 2 2 3 13 7 15 13 2 15 13 7 15 13 13 2
9 15 15 4 13 2 16 13 0 2
9 14 4 13 2 16 4 15 13 2
10 7 12 9 12 3 4 15 14 13 2
23 14 3 0 9 12 4 9 11 13 9 2 16 15 4 13 3 3 0 0 9 1 9 2
14 9 4 15 13 9 2 13 7 14 4 9 0 9 2
16 3 15 4 10 9 13 1 9 1 10 0 9 2 0 9 2
14 13 4 15 13 14 1 0 9 2 3 4 9 13 2
32 16 13 0 2 16 13 9 9 0 9 2 4 3 10 9 3 13 2 16 13 2 7 14 1 10 9 15 15 14 3 13 2
45 0 11 2 0 9 11 4 1 0 0 9 1 9 1 11 2 1 15 3 13 12 12 9 2 13 13 0 9 1 9 9 2 15 9 4 1 0 9 13 1 12 1 12 9 2
40 1 9 2 16 13 14 0 9 9 0 0 9 2 16 15 4 13 1 11 7 4 14 1 0 9 13 12 9 9 2 4 11 11 13 12 9 9 0 9 2
23 1 9 0 9 1 9 0 9 7 9 4 1 0 3 7 1 3 13 0 0 0 9 2
11 10 9 13 9 0 9 0 7 0 9 2
14 13 7 14 3 0 9 1 0 9 9 1 0 9 2
35 9 1 9 1 9 1 11 2 9 0 9 11 7 9 0 9 11 11 2 13 2 16 13 10 9 9 1 0 0 9 3 0 1 9 2
2 3 2
6 2 16 13 14 9 2
12 11 15 4 3 13 2 9 13 1 0 0 2
13 9 4 13 3 13 2 16 4 15 3 13 9 2
17 3 13 0 9 12 0 9 2 1 15 7 9 11 13 1 9 2
17 1 9 1 12 9 1 3 12 12 0 9 13 9 1 9 9 2
7 7 13 0 9 1 15 2
20 1 0 9 7 4 15 14 9 13 7 14 13 14 15 2 15 15 13 0 2
7 0 9 1 9 13 0 2
12 1 11 13 9 3 3 0 1 15 1 11 2
24 3 16 13 1 9 0 9 1 3 12 12 9 1 0 9 2 13 1 0 9 3 12 9 2
20 0 9 2 16 4 13 1 11 3 12 9 2 13 1 11 12 1 12 9 2
25 0 9 2 16 4 13 2 4 13 14 9 1 9 1 0 9 2 0 1 9 9 1 0 9 2
19 9 4 13 10 9 2 16 15 4 13 1 0 9 9 9 7 0 9 2
21 1 0 9 13 13 0 7 0 15 8 11 2 16 13 7 15 13 1 9 9 2
18 1 9 0 9 4 13 0 9 2 13 7 4 15 1 9 1 11 2
24 0 7 0 9 1 9 4 1 9 0 9 10 9 13 8 0 9 9 1 11 11 7 11 2
24 0 9 4 10 9 1 9 13 2 16 13 1 15 1 9 0 8 11 7 10 9 11 11 2
28 11 2 12 0 0 9 11 1 9 0 9 9 1 11 13 3 1 12 9 1 9 11 1 11 0 0 9 2
9 9 7 13 14 9 9 7 9 2
19 7 14 10 9 15 9 0 0 9 13 1 0 0 9 0 9 9 11 2
32 16 9 13 2 16 13 0 9 0 7 0 2 13 3 10 9 9 7 0 9 1 9 7 9 1 9 1 9 7 0 9 2
31 11 2 12 1 9 1 0 9 4 10 9 11 11 1 0 9 13 14 3 3 7 13 14 3 0 1 9 11 7 11 2
21 9 9 9 15 13 14 11 11 2 3 16 4 11 11 1 11 13 14 3 3 2
16 11 11 4 14 0 9 13 0 9 1 12 3 1 0 9 2
17 1 3 4 1 9 1 11 10 9 1 12 9 13 14 11 11 2
30 1 12 9 1 0 9 9 0 9 4 1 9 1 9 1 3 13 14 11 11 2 3 16 15 11 11 14 3 13 2
12 9 9 14 4 1 0 9 13 13 0 9 2
12 9 4 9 13 9 3 2 16 15 4 13 2
20 9 4 3 13 0 9 7 13 10 9 2 16 4 15 3 13 1 0 9 2
20 1 0 4 13 14 9 1 9 2 7 4 9 13 2 16 4 15 3 13 2
29 13 4 0 9 2 0 9 9 0 9 7 4 13 2 16 1 0 9 14 4 13 2 16 15 14 4 13 9 2
11 3 4 15 1 9 13 1 9 1 11 2
7 11 13 3 12 0 9 2
13 9 1 0 9 2 11 2 4 13 0 9 12 2
11 13 14 9 7 13 3 1 9 0 9 2
5 13 9 0 9 2
21 10 0 9 7 13 0 1 9 0 9 2 11 2 2 16 4 13 0 9 12 2
16 1 9 1 0 13 9 0 9 7 9 0 9 1 0 9 2
10 13 2 16 13 0 9 3 0 9 2
26 1 11 7 14 3 3 13 9 1 9 11 11 2 1 15 9 1 15 13 2 16 13 9 0 9 2
10 1 15 13 9 9 1 10 0 9 2
24 3 15 4 1 9 13 0 0 9 1 9 2 13 7 15 15 4 14 9 0 9 1 11 2
23 7 10 9 8 11 4 1 0 9 1 0 11 13 2 16 15 1 9 11 13 0 13 2
13 1 15 4 3 13 9 1 9 0 9 1 9 2
19 11 2 12 2 0 0 9 4 15 13 1 9 1 9 0 9 0 11 2
19 13 15 4 1 0 11 2 0 9 7 0 9 10 9 2 9 11 11 2
22 3 9 9 14 4 13 0 2 7 3 1 0 9 0 0 9 1 15 13 0 13 2
7 7 14 14 13 9 15 2
8 0 0 9 15 13 1 0 2
20 3 13 1 15 0 14 10 9 2 7 4 0 9 1 15 13 3 0 11 2
17 1 9 7 1 15 13 14 2 16 13 1 0 0 9 9 11 2
36 11 2 1 9 0 9 1 9 8 11 1 0 9 1 9 11 4 10 16 12 9 2 3 1 9 12 0 9 2 13 0 0 9 1 11 2
18 12 2 0 9 4 10 16 12 9 13 2 15 7 4 15 14 13 2
18 9 4 0 9 3 13 2 7 13 12 0 9 0 0 9 1 11 2
7 3 4 13 13 0 9 2
25 9 11 11 4 13 2 16 4 3 13 9 2 9 1 9 7 14 13 1 10 9 1 0 9 2
3 2 8 2
16 11 2 12 2 9 12 13 1 15 3 14 9 0 9 9 2
25 16 4 13 0 0 9 8 8 2 14 4 3 1 9 1 12 9 9 9 13 2 10 9 2 2
30 1 12 4 9 1 11 13 0 9 2 16 4 13 1 0 9 7 9 1 9 0 9 12 1 9 12 9 1 11 2
17 1 9 4 13 0 9 2 9 2 9 2 9 2 9 7 9 2
5 9 13 12 9 2
21 1 10 9 1 9 7 4 1 11 10 9 1 12 9 13 1 9 1 0 9 2
24 3 4 15 13 14 9 2 7 16 1 9 2 16 4 15 13 12 9 2 4 13 0 9 2
3 2 8 2
12 9 4 13 12 9 12 1 9 9 9 11 2
25 0 0 9 1 11 13 2 16 4 9 14 13 2 7 3 15 13 12 9 0 9 12 9 9 2
40 14 3 4 13 1 15 9 11 11 0 9 2 16 4 0 9 13 2 16 4 1 9 1 0 9 13 0 9 10 9 2 16 15 4 13 10 9 11 11 2
18 15 7 13 9 0 9 1 9 7 1 15 0 9 11 1 0 9 2
34 9 1 0 9 9 13 1 9 2 16 13 9 1 9 9 1 9 0 9 7 1 9 10 9 9 0 9 7 9 0 9 7 9 2
37 9 7 9 1 9 9 13 2 16 13 0 7 0 9 1 0 9 0 9 2 16 13 1 9 1 9 7 16 13 0 2 16 13 0 10 9 2
42 9 0 9 13 9 1 9 1 9 2 3 4 9 9 13 2 13 7 13 3 2 16 13 10 9 1 9 0 9 1 0 9 9 2 16 13 1 9 1 0 9 2
13 15 15 13 1 9 1 9 1 9 9 10 9 2
32 0 9 13 9 1 9 7 13 2 16 4 0 9 2 9 2 9 7 9 13 2 16 4 15 15 13 1 9 9 1 9 2
16 9 15 13 1 9 1 3 2 16 13 3 9 1 0 9 2
16 11 2 9 9 13 2 16 13 14 1 9 2 7 9 13 2
10 1 11 4 15 3 13 1 9 9 2
9 13 15 4 2 16 3 13 9 2
15 3 4 13 13 9 2 13 15 4 9 7 9 1 15 2
9 11 2 14 2 3 13 3 0 2
6 1 9 15 4 13 2
14 11 2 9 4 13 13 15 2 16 4 13 15 3 2
23 2 3 2 7 3 13 9 9 1 9 7 9 10 9 15 13 0 2 13 3 1 9 2
22 9 15 13 13 1 0 9 1 9 7 14 14 13 0 9 9 1 0 0 9 3 2
2 11 2
26 3 13 1 9 12 9 2 16 3 16 10 10 9 13 2 16 4 9 9 13 0 9 7 0 9 2
36 16 7 4 0 9 13 14 1 0 13 1 0 9 0 9 2 4 13 2 16 13 0 9 9 11 11 2 3 13 1 0 9 7 0 9 2
17 1 9 14 13 13 9 2 16 3 1 9 13 14 9 0 9 2
21 3 16 13 14 8 8 0 9 2 3 0 9 7 13 9 1 0 9 10 9 2
32 16 13 0 9 3 3 2 13 1 0 0 0 9 9 13 9 10 9 1 9 9 0 9 2 16 15 13 9 1 0 9 2
13 16 13 9 15 0 13 2 0 9 1 15 13 2
42 16 4 15 1 9 2 16 4 1 9 0 9 0 9 13 3 2 13 1 0 0 0 9 2 1 10 9 9 1 9 9 7 0 9 9 13 2 16 9 13 3 2
37 1 9 15 4 13 2 16 4 13 2 16 14 4 0 9 1 9 13 1 12 9 0 9 2 1 15 14 4 2 1 0 9 13 2 12 9 2
15 9 4 15 1 15 13 2 16 4 9 13 1 0 9 2
3 2 8 2
7 13 15 4 1 0 9 2
10 1 9 4 14 13 9 7 15 13 2
6 15 4 13 1 9 2
22 9 9 1 0 11 1 9 11 1 9 12 9 2 9 1 0 9 3 13 0 9 2
18 9 13 0 0 9 11 11 1 9 0 11 2 16 14 3 14 13 2
18 0 9 0 9 0 9 13 3 0 1 9 2 16 13 9 14 3 2
21 16 13 9 9 1 9 1 9 0 2 3 9 1 9 13 2 1 15 9 13 2
17 11 11 13 1 0 9 2 16 0 9 13 14 9 1 0 9 2
3 2 9 2
20 1 0 9 4 0 9 1 9 7 9 13 0 0 9 0 9 1 12 0 9
26 12 0 0 9 4 1 9 13 9 9 3 1 12 9 9 7 12 9 7 3 13 12 9 9 9 2
24 1 12 9 13 0 9 0 13 9 1 9 1 0 12 9 2 9 9 7 1 0 12 9 2
6 3 15 13 0 9 2
17 15 13 2 1 15 13 2 15 1 15 3 14 13 9 1 9 2
14 0 13 9 7 9 15 2 16 15 1 0 9 13 2
9 7 14 0 0 9 3 13 9 2
16 14 0 7 0 9 13 0 9 2 16 4 13 15 1 9 2
49 3 4 1 9 1 9 1 9 1 9 13 0 9 2 0 12 0 9 2 1 15 4 11 13 12 9 9 7 16 4 14 0 9 13 1 2 9 2 3 3 16 12 12 9 1 11 7 11 2
31 1 15 4 13 14 0 0 0 9 11 11 2 16 4 13 3 3 1 11 7 15 13 1 9 0 0 2 0 0 9 2
7 9 13 15 3 0 9 2
23 9 9 4 11 11 13 1 12 9 2 16 15 4 13 0 9 7 15 3 13 14 15 2
34 7 14 12 0 9 4 13 3 2 16 4 0 0 7 0 9 11 13 2 1 9 7 4 3 1 15 13 14 10 0 9 7 9 2
34 9 0 9 2 1 15 15 4 3 1 10 9 13 9 1 9 2 16 4 13 0 14 12 0 9 2 7 15 4 0 9 7 13 2
18 1 10 9 1 0 9 11 4 12 2 0 11 13 1 9 1 9 2
22 0 9 4 3 3 13 2 9 1 9 12 9 0 9 7 14 4 3 13 10 9 2
40 11 9 0 9 11 11 4 13 9 0 9 1 0 9 2 16 13 3 0 9 2 0 9 2 1 9 0 9 2 16 4 13 15 3 3 3 9 0 9 2
31 3 13 9 0 3 2 16 4 3 11 3 3 13 9 2 16 15 13 1 3 0 9 0 9 2 13 9 11 11 11 2
17 9 4 0 9 3 13 2 11 11 7 4 13 1 9 1 9 2
21 1 10 9 4 13 0 9 1 9 13 9 9 0 7 13 9 10 3 0 9 2
11 9 4 15 13 13 1 9 12 2 3 2
15 0 9 4 13 12 9 2 12 15 4 13 1 0 9 2
7 9 4 13 9 1 9 2
23 0 9 15 7 13 1 9 2 1 9 7 4 9 10 9 3 13 1 0 9 0 9 2
33 1 15 14 1 0 9 0 9 13 0 9 9 3 0 9 2 1 15 4 1 12 9 11 2 11 3 13 1 12 9 9 9 2
3 2 8 2
42 11 2 12 9 8 11 11 4 3 3 1 0 9 13 12 0 0 9 2 1 15 15 4 1 12 9 13 12 9 1 12 9 2 13 7 15 4 3 12 0 9 2
30 1 10 9 4 13 2 16 13 9 13 9 1 9 9 7 9 1 9 7 3 13 1 15 2 3 13 0 0 9 2
16 3 0 9 2 3 0 9 7 0 9 13 13 1 0 9 2
19 3 3 0 15 13 0 9 12 11 2 16 14 3 13 3 10 0 9 2
32 0 13 1 3 0 9 1 12 3 0 9 2 3 0 0 9 7 0 9 2 16 15 13 9 1 9 7 9 1 0 9 2
9 0 9 4 13 1 9 1 9 2
14 13 4 1 11 7 10 9 2 16 4 13 0 9 2
4 13 15 0 2
3 14 0 2
16 3 13 0 9 2 7 13 10 9 9 7 15 3 14 13 2
11 0 0 9 3 0 0 9 13 1 9 2
18 3 15 13 2 3 4 2 16 4 13 2 15 15 13 2 13 13 2
17 14 4 13 15 0 2 7 4 13 9 3 14 3 3 0 15 2
10 7 15 13 0 0 9 1 11 11 2
8 10 9 13 3 13 7 13 2
19 15 13 0 7 1 0 9 2 16 13 9 1 9 9 2 16 1 0 2
15 16 13 9 1 15 15 7 0 2 14 4 13 13 9 2
15 13 2 16 13 1 0 9 3 0 9 2 9 0 9 2
9 14 3 0 13 9 9 1 9 2
12 1 10 9 15 13 14 9 13 9 10 9 2
8 7 14 13 13 1 9 9 2
21 3 14 4 12 9 0 9 3 1 9 13 12 9 9 7 15 3 13 0 9 2
25 1 12 1 9 4 9 1 0 0 9 13 0 9 2 9 7 4 3 9 13 1 0 0 9 2
27 10 9 4 3 13 2 3 13 9 9 1 9 1 0 9 1 0 9 2 10 9 13 0 1 0 9 2
16 15 13 0 9 2 16 13 0 1 0 9 2 0 13 9 2
16 1 9 0 9 11 13 0 9 0 1 0 9 2 1 9 2
9 15 3 13 0 9 9 1 9 2
12 0 9 9 2 8 2 13 1 9 9 11 2
17 0 9 8 2 9 2 13 0 0 9 7 13 1 9 9 11 2
11 0 9 8 2 11 2 13 1 9 11 2
12 0 9 8 2 0 9 2 13 1 9 11 2
13 0 2 0 9 9 2 9 2 13 1 9 11 2
17 9 13 9 11 1 9 2 13 0 0 9 2 9 7 9 9 2
11 13 0 9 2 9 7 0 9 0 9 2
21 0 9 1 0 9 15 4 13 12 9 2 15 12 9 1 9 4 13 0 11 2
21 0 9 1 9 4 13 0 9 2 1 15 4 15 13 9 3 2 3 7 3 2
13 9 4 13 1 9 2 16 4 13 7 13 11 2
21 1 0 9 4 13 0 2 9 2 1 9 9 7 9 2 16 4 13 0 9 2
12 7 14 1 9 3 10 9 13 1 0 9 2
13 9 7 3 13 14 3 2 3 13 9 3 0 2
12 11 11 2 12 2 1 9 3 13 10 9 2
14 3 13 15 0 2 0 2 0 2 0 7 0 9 2
5 9 15 13 9 2
18 1 9 1 9 2 16 13 0 9 2 13 0 0 9 1 0 9 2
31 14 3 1 9 9 1 9 3 13 0 7 0 0 9 1 0 0 7 0 0 9 2 16 4 13 1 9 9 9 2 2
15 1 15 4 13 3 13 9 7 9 9 1 10 0 9 2
24 9 0 9 13 1 12 9 7 13 7 1 0 9 13 9 2 1 15 13 14 1 12 9 2
7 9 1 9 13 14 0 2
13 9 15 13 1 9 2 16 15 9 13 1 15 2
20 9 15 13 1 0 9 9 2 3 7 15 14 3 13 1 0 9 1 9 2
25 9 1 9 2 9 7 9 0 0 9 13 1 9 1 11 1 0 9 2 16 13 14 0 9 2
12 0 9 13 0 0 9 7 0 9 0 9 2
28 16 13 9 1 9 3 0 2 15 13 9 1 10 9 0 13 1 0 0 9 1 0 9 1 9 0 9 2
9 3 13 3 0 10 9 9 9 2
19 1 9 13 14 0 0 9 2 16 9 1 9 13 1 0 9 7 9 2
18 1 9 14 4 15 13 12 9 1 9 2 1 15 14 13 13 9 2
18 9 7 9 2 16 4 13 1 9 9 10 0 9 2 13 9 0 2
27 1 0 9 15 3 1 12 9 13 1 9 2 16 13 1 12 2 0 9 7 13 0 14 1 9 9 2
18 0 9 1 0 13 3 12 9 2 1 9 7 4 13 13 14 9 2
23 1 0 9 13 3 13 3 12 9 9 2 9 1 0 9 7 13 1 12 1 12 9 2
26 16 9 14 13 13 2 15 13 1 9 9 9 1 9 1 9 9 7 13 9 1 9 1 0 9 2
10 13 14 9 2 16 13 3 3 0 2
11 0 9 7 9 2 16 13 0 2 13 2
24 1 9 11 7 11 15 13 10 0 9 2 16 1 10 9 7 9 13 10 14 3 0 9 2
19 9 11 13 1 3 0 9 7 14 10 9 4 13 13 10 3 0 9 2
19 1 0 9 1 9 14 3 13 1 9 1 9 1 9 2 2 13 11 2
16 0 9 0 9 11 10 9 13 9 1 9 1 12 9 9 2
16 1 9 2 12 9 2 15 4 1 9 11 13 3 12 9 2
32 13 4 9 9 7 0 9 11 7 0 9 11 2 9 1 9 7 13 14 0 9 11 2 9 11 1 0 11 7 9 11 2
4 13 4 0 2
23 1 9 1 9 7 1 9 9 1 10 9 11 13 0 1 9 9 13 1 0 0 9 2
36 0 9 11 12 2 16 11 13 0 9 11 2 13 0 2 7 1 10 9 4 13 9 2 16 4 1 0 9 0 0 9 3 13 10 9 2
14 3 7 15 13 2 16 9 3 7 4 13 14 0 2
40 3 11 2 12 2 13 2 16 4 0 2 0 9 1 9 9 3 13 10 9 2 3 3 7 15 4 13 2 16 11 1 9 7 0 9 4 13 3 0 2
32 7 4 13 0 3 2 16 15 9 0 11 7 0 0 9 11 3 13 7 4 0 9 1 15 13 3 1 9 9 9 11 2
19 0 4 13 1 3 3 0 9 7 4 13 13 10 0 9 3 0 9 2
30 16 4 9 13 1 9 7 1 15 14 0 9 0 9 7 0 9 1 0 9 2 15 4 10 9 14 3 3 13 2
23 7 1 9 9 4 13 9 14 0 0 9 2 7 14 0 2 1 15 13 9 1 9 2
17 1 10 9 10 12 9 13 0 9 15 2 16 4 13 0 9 2
25 1 10 9 4 13 14 9 9 7 9 1 9 2 16 15 13 1 9 7 1 10 9 1 15 2
17 1 9 15 3 13 7 14 3 13 9 9 7 13 1 0 9 2
54 9 9 7 9 2 9 11 1 11 7 0 9 11 4 1 9 2 12 9 2 1 0 9 11 13 2 9 9 7 9 2 2 1 15 4 16 9 13 14 9 0 9 11 7 0 9 9 0 9 1 0 0 9 2
37 11 11 7 9 9 11 4 0 13 10 9 2 3 16 4 15 9 0 9 9 11 1 9 9 11 11 13 1 0 9 0 0 11 7 0 11 2
21 16 4 9 3 13 2 4 13 14 0 9 9 9 7 11 11 1 11 1 9 2
41 11 4 14 1 12 9 1 10 9 13 0 9 1 0 9 2 3 7 15 4 0 9 3 1 0 11 7 1 11 13 14 0 9 1 3 0 9 1 0 9 2
17 3 15 4 1 9 13 1 9 9 2 3 7 15 4 13 9 2
8 1 9 4 13 12 9 9 2
9 9 0 9 1 10 9 9 11 2
19 9 11 13 0 13 0 9 1 9 0 9 9 2 9 7 0 0 9 2
28 1 0 0 9 4 13 0 9 1 11 7 15 3 13 1 9 0 9 11 11 2 16 4 13 3 1 9 2
35 1 9 12 2 16 15 4 13 1 10 9 2 15 4 1 0 9 13 1 9 0 0 9 0 9 2 16 4 10 9 3 13 9 9 2
27 1 0 9 4 13 9 1 10 9 1 0 9 9 2 16 13 3 7 3 0 1 10 0 9 0 9 2
11 3 4 1 0 13 9 9 7 0 9 2
15 0 9 11 11 4 13 9 2 16 4 13 0 7 0 2
32 3 4 13 9 10 9 2 16 13 9 1 9 9 1 0 9 7 15 1 10 9 13 1 9 9 2 7 13 15 10 9 2
30 1 9 4 9 13 1 9 1 9 1 9 9 1 0 9 1 9 0 9 9 2 16 4 13 9 1 9 0 9 2
30 9 15 4 1 0 9 13 1 9 1 0 9 2 16 4 13 9 9 2 13 0 0 9 7 13 1 0 9 9 2
18 1 11 2 1 11 7 1 11 4 14 1 0 9 13 9 0 9 2
12 0 9 1 0 9 4 13 9 11 11 11 2
33 11 2 1 9 1 12 9 4 15 1 9 11 13 1 0 9 7 1 9 2 3 16 4 9 8 8 13 2 1 9 13 9 2
19 3 4 13 14 1 9 2 16 4 1 0 9 13 9 7 15 14 13 2
10 9 4 3 13 1 0 12 12 9 2
33 9 1 10 9 4 1 11 13 12 9 3 7 13 9 2 16 4 13 0 9 7 9 0 9 2 16 3 13 12 2 9 9 2
5 2 14 2 13 2
8 13 2 1 9 15 9 13 2
9 1 0 9 13 0 9 2 9 2
39 1 0 9 4 13 9 0 9 11 11 2 1 15 13 11 11 2 11 11 7 11 11 2 16 9 7 4 13 14 9 11 11 7 11 11 1 9 9 2
23 1 10 0 9 15 0 9 13 3 2 16 15 1 10 12 9 9 13 12 9 0 9 2
22 1 9 1 0 9 12 2 12 13 9 14 1 9 2 12 2 1 12 1 12 9 2
14 9 1 0 9 12 1 12 13 0 2 0 1 9 2
13 1 9 13 0 7 0 2 0 13 3 14 9 2
9 2 14 13 2 2 13 9 9 2
14 0 9 13 13 2 16 9 13 7 16 14 13 9 2
4 1 9 13 2
13 14 3 3 13 2 16 4 13 10 0 9 3 2
22 1 0 9 4 13 9 3 0 2 7 4 1 9 9 13 9 12 0 9 0 9 2
16 1 15 4 9 0 9 13 9 1 12 9 2 11 7 11 2
21 9 4 1 15 0 0 13 0 9 2 1 15 13 0 9 7 12 13 0 9 2
13 1 15 4 13 0 9 0 0 9 1 0 9 2
36 1 12 9 3 2 16 4 13 0 0 9 1 9 0 9 2 1 12 9 4 13 12 9 2 15 13 1 0 9 3 16 1 10 9 3 2
11 11 1 11 13 9 1 11 1 0 9 2
36 2 3 11 13 2 3 1 11 14 12 9 13 14 9 2 16 15 4 3 13 0 0 9 2 15 7 4 13 0 9 11 2 11 7 11 2
14 7 14 15 13 11 2 16 0 9 1 11 13 0 2
4 13 7 13 2
13 3 13 10 9 2 16 13 0 0 2 0 9 2
8 13 1 9 2 0 9 2 2
6 3 15 15 13 9 2
13 13 0 2 16 9 14 13 13 9 2 16 13 2
10 14 13 7 13 1 0 9 1 9 2
15 0 9 3 14 13 1 9 2 16 1 15 13 0 9 2
22 1 9 15 3 13 7 13 2 15 13 3 0 9 7 10 9 2 0 9 7 9 2
13 10 9 3 13 7 13 1 9 7 9 1 9 2
17 15 12 4 1 0 13 3 1 9 0 0 9 9 12 1 11 2
21 14 1 9 2 16 4 13 13 9 2 4 1 9 0 0 9 1 9 13 9 2
24 16 7 15 15 9 4 13 13 2 4 15 13 2 16 15 4 13 16 9 0 2 0 9 2
4 9 4 13 2
16 2 1 9 9 7 11 4 13 14 9 2 9 1 9 2 2
21 0 4 13 2 16 4 13 9 1 9 2 1 0 9 7 15 4 13 14 12 2
19 9 4 13 3 0 1 9 9 2 16 4 13 9 13 14 0 11 11 2
22 9 2 10 0 9 4 1 9 13 10 10 9 2 16 4 1 9 9 13 1 11 2
20 15 0 9 14 4 13 2 16 4 13 13 14 9 1 0 12 0 0 9 2
25 14 7 13 0 2 16 11 14 4 13 9 2 7 1 9 3 9 11 13 2 3 13 12 9 2
12 0 0 9 4 0 9 9 3 13 14 12 9
15 0 9 4 1 0 9 13 2 0 9 4 13 11 11 2
19 16 15 4 13 1 0 9 2 4 3 13 3 12 9 1 9 0 9 2
18 3 4 10 9 3 3 13 2 16 13 9 10 10 9 1 0 9 2
23 7 15 4 3 13 7 1 15 15 4 3 13 13 9 1 3 0 0 9 2 11 9 2
35 11 2 12 9 1 0 9 9 1 0 9 4 1 0 9 1 0 9 7 0 9 13 0 9 2 16 4 15 3 7 3 13 0 9 2
25 13 4 1 9 9 0 9 2 16 4 13 9 7 1 15 13 14 0 9 2 16 4 15 13 2
17 9 2 16 4 3 0 13 7 13 0 9 2 4 13 0 9 2
5 3 13 7 13 2
3 13 15 2
7 1 0 9 13 0 9 2
21 14 7 13 3 0 9 14 14 1 12 9 2 1 11 2 1 11 7 1 11 2
22 14 2 15 13 1 0 9 1 9 11 1 0 11 2 9 7 15 13 1 0 9 2
9 14 12 9 1 9 13 9 9 2
23 0 9 8 11 11 4 1 15 13 2 2 9 1 9 0 9 1 9 0 9 13 0 2
15 3 15 13 13 9 2 3 7 15 4 13 1 9 9 2
15 1 9 13 3 0 0 9 2 14 3 15 13 0 9 2
18 3 13 9 9 9 10 9 2 16 7 3 13 14 0 9 1 9 2
19 12 9 1 15 2 16 13 0 1 9 9 2 4 15 13 10 9 1 9
31 10 9 2 16 4 13 11 1 11 2 4 14 0 0 9 13 9 0 0 9 1 11 2 15 7 4 13 0 9 8 2
7 11 4 3 13 0 9 2
31 12 0 0 9 4 13 1 0 9 9 2 0 7 4 3 13 1 0 9 0 9 2 16 15 9 9 4 1 9 13 2
19 11 4 3 3 13 10 9 7 1 10 0 9 15 4 9 1 9 13 2
34 11 4 13 11 2 3 0 9 13 9 2 1 15 15 4 13 2 16 4 11 3 13 10 9 1 9 7 3 13 14 10 0 9 2
14 2 0 13 2 2 4 13 7 0 4 15 15 13 2
5 11 15 4 13 2
14 2 0 9 1 9 13 12 9 2 2 4 13 11 2
12 2 14 2 13 15 2 2 4 3 13 11 2
5 11 4 13 9 2
16 3 3 15 4 13 13 1 0 9 2 16 15 4 0 13 2
7 4 14 13 1 0 9 2
15 3 4 13 0 10 9 1 11 7 9 4 15 13 0 2
16 9 4 15 9 3 13 2 3 7 4 10 9 13 1 9 2
22 9 4 13 1 10 9 0 2 7 11 14 4 13 9 2 16 15 14 4 13 13 2
21 7 1 9 1 9 2 16 15 4 3 3 13 1 10 0 9 2 4 9 13 2
12 16 4 11 13 0 9 2 14 4 13 9 2
8 13 4 0 9 1 0 9 2
16 0 9 2 16 15 4 13 1 9 2 15 4 13 1 9 2
12 3 4 15 13 9 2 3 15 13 1 9 2
19 7 9 4 13 9 1 9 9 9 2 7 15 4 13 13 1 10 9 2
8 2 13 4 9 1 10 9 2
16 13 4 1 0 9 9 7 15 3 13 1 10 9 7 9 2
9 1 9 15 4 13 0 0 9 2
10 9 4 13 13 0 1 9 15 9 2
7 9 4 13 3 3 0 2
5 8 8 8 8 2
2 9 2
24 9 9 12 4 13 3 0 0 9 2 1 9 4 13 13 10 9 2 16 4 13 0 9 2
33 13 15 2 16 4 15 3 1 0 9 13 1 9 2 16 4 1 0 9 13 1 0 9 2 16 4 15 13 1 0 0 9 2
22 13 4 15 14 1 10 9 1 0 9 2 13 4 0 2 0 1 0 2 0 9 2
29 1 0 9 1 0 0 9 3 4 13 9 2 16 4 13 11 1 9 7 3 14 1 9 2 3 3 3 0 2
13 1 9 12 2 12 4 3 13 9 1 9 9 2
18 9 4 13 2 16 4 9 13 11 11 2 0 0 9 1 0 9 2
9 15 4 13 2 16 13 1 15 2
6 11 4 10 9 13 2
17 16 15 3 13 2 4 16 9 13 2 16 13 0 1 0 9 2
16 14 3 7 15 13 16 9 2 16 15 4 13 2 4 13 2
19 13 4 2 16 4 13 13 1 9 12 2 16 4 13 3 3 0 9 2
18 3 15 9 1 0 9 2 16 4 15 15 13 15 2 4 3 13 2
15 16 4 1 10 9 13 9 13 2 4 15 0 13 9 2
22 1 0 9 4 13 0 9 2 11 11 2 11 11 2 11 11 7 3 0 11 11 2
37 1 9 2 16 4 13 9 1 9 12 2 4 15 13 1 9 11 2 16 4 13 0 0 9 11 11 2 16 4 13 3 9 1 0 0 9 2
32 3 12 9 3 2 12 9 12 2 4 11 11 13 9 9 9 2 1 15 4 10 0 9 13 10 3 0 7 0 0 9 2
26 1 0 0 9 1 0 9 4 13 14 9 2 1 15 4 11 3 3 13 10 9 1 9 7 9 2
11 1 9 13 1 9 11 2 0 0 9 2
28 1 10 0 9 4 13 9 2 16 4 14 3 13 2 3 4 13 14 10 0 9 1 10 0 9 10 9 2
25 16 4 13 14 12 9 0 9 2 15 4 9 9 13 2 14 16 4 1 15 13 12 0 9 2
44 1 0 9 4 13 9 1 9 9 10 9 7 1 12 9 15 4 0 9 1 9 13 1 9 0 9 0 9 7 9 2 9 9 7 13 9 2 16 15 14 4 14 13 2
12 14 1 10 9 15 4 13 0 9 1 15 2
26 3 4 13 9 2 16 4 13 2 16 4 13 10 9 1 9 2 9 7 0 9 2 13 1 9 2
20 15 14 4 15 13 1 9 12 2 16 4 10 9 13 14 1 9 12 9 2
26 13 4 3 0 2 16 15 4 15 3 13 2 7 4 14 10 9 1 15 13 13 10 9 1 9 2
24 11 11 2 9 0 9 2 15 4 13 9 0 9 11 2 16 15 4 13 0 11 11 11 2
31 1 9 14 4 13 0 9 9 0 9 2 16 4 15 1 0 9 1 0 9 13 1 9 7 15 10 9 14 3 13 2
24 13 0 9 2 7 13 1 9 3 0 9 10 9 13 9 0 2 14 3 0 9 1 9 2
22 1 11 4 3 13 14 1 9 0 9 2 16 4 13 16 9 1 9 1 0 9 2
3 0 0 9
13 15 14 4 0 9 13 9 2 4 3 13 9 2
22 0 13 2 16 13 11 7 11 3 0 2 16 15 13 1 9 2 0 9 7 9 2
36 7 14 3 4 13 0 0 9 1 9 9 2 16 15 15 13 7 0 13 7 15 1 15 3 13 9 9 7 14 13 9 9 1 10 9 2
41 9 7 10 9 4 3 13 14 9 9 0 9 0 9 2 15 0 9 13 3 13 7 13 11 2 16 4 13 12 3 0 7 0 0 9 1 0 2 0 11 2
12 2 13 1 10 9 2 13 4 15 0 9 2
16 9 15 4 1 9 0 9 13 1 10 9 2 2 4 13 2
29 11 15 4 1 9 9 1 15 13 13 9 2 16 15 4 1 9 9 14 0 13 2 7 13 3 1 9 11 2
22 15 7 13 3 11 2 16 13 2 16 13 9 0 9 0 9 1 0 9 3 0 2
26 7 13 1 11 0 13 9 2 16 13 1 0 9 12 9 7 0 2 16 0 9 13 1 12 9 2
31 1 15 13 0 11 2 16 13 2 16 13 16 9 11 11 9 13 9 1 9 2 16 0 1 0 9 12 9 13 0 2
18 3 4 15 9 13 0 12 1 0 2 9 7 1 15 13 0 0 2
21 14 10 9 4 1 0 9 3 13 9 2 16 4 1 9 9 3 13 3 3 2
44 1 0 9 2 16 15 4 13 1 0 9 1 0 9 2 1 15 13 0 12 9 2 4 9 1 9 0 9 13 14 1 9 2 3 7 13 9 1 9 0 9 1 9 2
24 16 7 15 4 3 13 9 2 13 1 0 0 0 9 2 16 15 4 13 2 13 0 9 2
35 1 0 9 2 9 2 9 7 9 2 1 0 7 0 9 7 1 0 9 9 1 9 11 11 3 13 16 3 0 2 0 7 0 9 11
16 0 9 13 0 2 7 15 2 1 15 15 3 13 1 9 2
18 15 13 9 2 16 13 1 0 11 2 0 9 11 7 0 9 11 2
32 13 4 2 16 3 4 13 13 1 0 9 0 9 2 7 4 13 13 10 0 9 2 16 14 4 13 9 1 0 0 9 2
26 1 9 9 11 11 13 11 0 9 0 0 9 1 0 9 1 12 2 12 1 12 2 12 2 12 2
27 11 2 9 12 2 1 15 4 11 1 0 13 10 9 2 13 9 2 0 9 7 0 9 1 9 3 2
20 1 9 7 13 14 10 0 9 0 9 7 9 2 16 15 14 13 10 9 2
12 1 0 9 1 9 13 14 10 9 0 9 2
32 1 9 4 13 9 12 0 2 3 16 0 7 0 9 13 1 0 9 2 0 0 9 2 16 4 3 13 2 9 9 2 2
32 10 0 9 13 14 1 0 9 9 2 16 13 1 9 9 9 9 9 11 2 11 2 16 13 1 9 0 0 9 1 9 2
14 16 15 13 14 3 3 2 9 13 1 9 7 9 2
12 9 1 9 13 1 9 7 13 1 0 9 2
14 1 0 9 3 14 0 9 2 13 2 8 0 9 2
13 9 10 9 13 14 1 9 0 9 2 9 9 2
24 16 15 9 13 7 15 13 9 7 13 0 9 2 3 9 13 9 2 16 13 15 15 0 2
17 1 0 9 9 15 13 13 2 16 1 10 9 14 4 15 13 2
15 13 4 10 9 2 16 14 4 13 0 9 1 10 9 2
19 3 0 0 9 4 13 0 1 10 9 2 16 1 9 7 9 13 9 2
10 15 4 13 0 1 9 3 1 9 2
13 9 9 13 9 9 2 16 13 16 0 9 9 2
18 16 15 13 2 13 9 1 10 9 7 0 9 13 10 9 1 9 2
11 1 10 9 15 13 0 9 9 1 9 2
48 0 4 13 2 16 4 1 9 0 9 2 16 15 3 13 1 9 9 7 1 0 9 2 13 9 1 9 2 15 7 4 1 0 9 13 1 9 1 9 2 16 4 13 10 9 3 0 2
19 12 10 3 0 9 1 11 11 13 9 11 2 16 13 1 9 3 0 2
20 16 13 0 14 12 9 2 15 9 13 13 1 9 2 7 3 13 3 0 2
25 3 4 9 13 1 9 2 16 14 15 3 13 10 0 9 7 16 14 10 9 13 14 10 9 2
13 16 15 4 13 2 15 4 13 9 13 1 9 2
11 9 4 14 13 1 9 7 13 1 9 2
7 10 9 7 3 3 13 2
26 11 13 11 2 16 14 13 10 9 1 0 9 2 7 16 10 9 13 1 15 2 16 13 14 0 2
27 11 13 9 0 2 16 15 4 13 1 10 9 2 15 7 15 13 2 16 13 1 9 1 10 9 11 2
12 11 13 11 11 2 16 1 0 9 13 9 2
16 11 13 11 1 0 0 9 2 16 13 11 2 16 13 9 2
22 11 13 2 16 4 11 13 11 9 2 1 15 4 13 3 3 0 0 0 9 11 2
12 1 9 14 4 13 9 14 1 0 9 11 2
27 1 11 2 3 12 9 3 1 0 0 9 2 4 13 14 12 2 1 15 13 3 10 9 16 1 0 2
19 9 14 13 1 9 2 7 16 13 1 3 0 9 0 1 9 0 9 2
17 14 3 4 1 11 13 0 9 2 16 15 4 13 14 0 9 2
28 15 2 16 4 15 0 9 13 14 1 0 9 2 7 15 4 3 1 9 13 1 0 2 4 13 11 11 2
20 3 16 15 4 11 11 13 2 4 13 1 9 16 0 0 9 7 0 9 2
17 9 9 13 9 11 11 2 12 0 7 15 13 1 0 9 9 2
18 7 0 9 11 7 11 1 9 7 11 1 9 10 0 9 13 3 2
17 0 9 4 14 13 2 16 4 13 0 0 9 1 0 0 9 2
16 9 14 13 2 16 1 9 14 13 9 1 9 0 0 9 2
11 9 4 9 13 1 12 9 1 0 0 9
5 11 13 10 9 2
5 13 1 0 9 2
60 9 10 9 2 16 15 3 13 1 9 2 15 4 13 1 9 2 9 7 9 2 16 13 10 0 9 7 13 10 0 9 2 4 13 11 11 2 16 15 4 3 1 11 11 7 11 11 1 12 9 13 1 0 9 1 0 7 0 9 2
10 0 13 1 0 0 0 9 1 15 2
7 7 15 13 1 9 11 2
14 13 4 3 1 15 2 16 15 0 9 11 3 13 2
30 7 16 4 1 10 0 2 0 0 9 1 3 0 0 9 14 3 13 3 2 4 13 9 10 9 1 9 13 3 2
17 3 13 11 0 2 1 0 9 7 1 9 13 14 11 7 11 2
14 9 0 11 4 13 2 11 7 4 13 14 14 3 2
11 1 9 9 15 3 13 2 1 9 13 2
10 7 0 15 1 9 3 14 13 14 2
13 1 12 9 9 9 13 0 13 1 12 9 9 2
16 11 4 14 9 10 9 13 13 9 1 9 9 11 1 11 2
12 9 1 9 0 9 1 0 9 4 13 0 2
19 9 1 0 9 12 9 10 9 15 13 1 9 12 9 1 9 0 9 2
14 9 13 0 0 9 1 9 9 7 0 9 0 9 2
19 1 9 1 9 9 15 0 9 1 0 9 12 9 10 9 14 13 13 2
30 9 1 9 13 0 9 1 15 2 10 0 9 0 9 13 1 0 9 0 2 0 7 13 14 9 9 9 1 9 2
22 13 9 9 2 16 15 4 9 13 1 0 11 1 9 11 2 11 2 11 7 11 2
30 9 11 11 15 4 1 0 9 3 13 9 0 9 7 15 3 13 9 1 0 9 2 16 4 15 13 1 10 9 2
14 14 1 0 9 4 13 2 16 13 11 0 9 15 2
24 3 0 13 7 3 13 13 2 15 13 7 10 13 10 9 2 7 15 13 1 9 1 15 2
14 9 13 0 7 15 15 14 10 9 1 9 3 13 2
35 1 10 9 3 13 0 9 2 14 14 1 9 1 15 2 7 14 1 15 2 16 15 13 1 9 2 9 2 9 7 0 9 1 9 2
7 14 13 15 1 10 9 2
28 10 10 9 1 11 13 15 0 9 2 16 15 13 0 13 2 16 13 15 3 13 7 0 15 13 3 3 2
16 15 2 16 15 1 15 13 2 13 2 3 15 10 9 13 2
18 11 15 4 13 1 9 7 1 15 13 1 10 0 9 3 7 3 2
19 13 15 14 3 13 1 15 7 10 9 7 3 1 15 13 3 3 0 2
17 15 15 4 13 7 15 3 13 9 1 9 0 9 7 0 9 2
26 12 9 0 9 0 9 11 1 11 4 1 0 9 13 2 3 13 1 10 9 14 10 9 7 9 2
25 1 12 9 1 9 9 13 0 9 4 9 1 9 9 11 11 7 11 11 2 11 13 0 9 2
16 7 3 4 15 13 1 10 0 9 2 16 4 3 3 13 2
22 13 4 0 9 7 9 9 2 13 9 1 9 9 7 13 9 0 0 7 0 9 2
8 10 9 4 13 1 0 9 2
39 16 15 4 13 2 15 4 13 7 15 1 9 13 3 3 1 9 2 16 4 14 3 13 2 11 7 4 13 16 4 13 0 7 0 7 13 0 9 2
17 16 4 9 3 13 1 15 2 15 4 13 1 9 7 3 13 2
47 16 4 1 9 14 13 2 16 13 3 13 9 2 4 13 1 9 3 1 9 7 4 14 13 2 16 4 13 1 9 1 9 2 16 4 3 13 10 9 7 13 1 9 1 10 9 2
46 1 10 9 7 15 4 13 2 16 15 9 7 9 9 14 4 14 13 2 7 15 4 1 10 9 9 2 16 4 13 1 9 2 3 13 1 0 9 7 13 1 0 9 0 9 2
11 13 15 4 14 2 16 4 15 0 13 2
14 14 2 14 10 9 4 13 7 9 15 4 13 13 2
22 1 10 9 7 9 15 4 9 13 9 2 16 4 14 1 9 13 3 7 1 9 2
11 13 4 2 16 4 0 1 0 3 13 2
34 0 9 13 11 11 1 9 0 9 2 9 7 13 3 16 11 0 1 9 7 9 2 16 3 13 1 9 9 2 9 2 9 12 2
32 1 15 2 16 13 3 10 9 2 7 7 13 1 0 9 2 16 4 13 1 9 1 0 9 13 9 1 9 2 13 9 2
20 15 14 13 1 9 7 14 0 9 9 2 7 1 0 9 15 3 13 9 2
37 15 7 13 2 16 4 3 10 9 13 1 9 2 9 2 16 15 15 13 9 2 7 1 0 9 4 14 15 13 1 9 10 0 9 2 2 2
23 15 2 15 13 3 13 2 13 13 9 11 2 16 15 3 1 0 9 13 1 9 8 2
32 9 9 2 9 1 9 9 13 14 14 0 1 10 3 0 0 9 7 1 10 10 9 2 16 1 0 0 9 13 10 9 2
18 9 9 2 9 3 14 13 2 16 13 1 0 9 13 9 2 9 2
13 9 9 0 9 13 1 10 9 7 9 0 9 2
10 9 9 4 13 14 9 2 11 2 2
15 3 15 13 2 16 13 1 9 10 1 10 9 0 9 2
14 7 15 15 14 13 1 9 2 16 4 15 13 9 2
29 13 3 1 15 15 1 0 9 2 13 9 7 1 9 13 9 2 16 4 15 15 3 13 7 13 1 15 0 2
33 3 16 4 11 1 0 9 0 9 11 12 13 11 2 7 4 11 13 9 1 3 0 9 1 9 0 9 0 0 9 11 12 2
13 10 9 1 9 7 9 0 0 9 14 13 0 2
15 16 14 13 1 9 2 1 10 9 14 3 13 9 11 2
15 0 9 9 4 1 9 9 1 9 2 9 13 0 9 2
25 16 13 3 0 2 15 4 1 9 13 9 2 16 13 15 3 2 7 13 3 0 9 3 0 2
14 3 13 14 9 1 9 2 0 1 12 9 0 11 2
19 14 13 0 14 9 1 0 9 2 16 13 14 3 0 16 0 0 9 2
9 3 13 0 13 1 9 9 9 2
17 1 9 9 13 0 3 2 9 7 13 1 9 2 9 3 0 2
18 1 9 1 9 9 15 4 13 0 9 2 1 15 3 13 10 9 2
23 3 13 13 1 3 0 2 16 13 3 13 10 9 7 9 9 2 9 7 9 2 9 2
22 9 9 7 9 13 9 1 9 2 0 9 0 9 2 9 9 11 2 11 2 2 2
9 9 13 10 0 9 1 10 9 2
18 10 9 13 3 14 10 9 3 7 14 0 9 9 15 15 3 13 2
15 9 9 15 4 3 13 1 0 9 0 9 7 0 9 2
17 1 0 11 7 1 11 13 3 0 2 1 0 9 7 13 0 2
10 12 0 9 4 13 9 1 0 9 2
13 9 11 11 1 9 4 13 2 14 15 4 13 2
12 13 7 4 2 16 13 1 0 9 1 11 2
29 9 11 11 2 16 15 4 0 13 1 9 7 13 3 14 0 0 2 4 13 2 3 4 3 13 14 12 9 2
11 9 4 1 9 0 9 13 1 0 9 2
19 3 3 4 13 14 11 8 1 0 9 2 1 15 14 4 11 13 9 2
27 13 4 1 0 9 2 13 4 2 16 4 15 7 10 9 13 9 7 16 15 15 15 14 4 14 13 2
13 14 10 9 11 8 14 13 13 14 9 1 11 2
27 15 15 4 14 3 13 2 1 9 7 4 13 2 16 4 0 13 2 2 16 4 15 1 9 13 2 2
20 1 0 9 4 13 2 16 13 14 9 1 10 9 7 14 13 9 1 9 2
16 15 15 13 2 16 15 11 11 1 9 3 13 1 11 11 2
42 1 9 4 13 11 11 2 1 15 15 4 13 2 16 14 4 13 9 9 3 7 15 13 2 16 4 0 11 14 13 9 9 7 15 1 9 10 9 13 0 9 2
6 11 11 15 13 13 2
14 2 13 11 7 15 13 0 13 2 2 4 13 9 2
18 2 1 10 0 9 15 4 13 1 9 2 13 7 15 4 14 11 2
16 11 2 2 11 13 2 16 15 10 9 13 2 16 13 15 2
8 0 9 9 15 13 0 13 2
24 2 9 14 0 11 13 16 9 2 3 7 13 14 10 12 0 9 1 0 9 1 9 11 2
19 7 10 3 0 9 2 16 15 3 3 13 2 13 2 16 4 13 9 2
9 3 15 4 11 3 13 10 9 2
5 14 2 13 9 2
18 1 9 1 11 4 13 14 3 2 16 4 9 1 0 9 13 9 11
36 9 1 0 9 2 9 9 1 15 2 15 4 1 0 13 1 11 7 10 13 9 2 16 15 14 13 1 9 0 2 4 13 9 0 9 2
27 1 0 0 9 4 13 3 10 9 2 11 4 13 9 2 3 10 10 9 9 1 9 13 1 9 9 2
30 10 0 9 4 13 0 1 9 11 2 10 12 9 1 11 2 16 4 0 9 7 9 9 9 1 9 9 14 13 2
28 13 14 2 16 13 0 9 1 9 0 13 9 0 9 9 2 14 7 13 2 16 13 9 9 7 9 0 2
22 11 15 4 1 9 0 9 13 1 10 9 7 13 2 16 13 0 9 0 1 9 2
10 0 9 9 7 15 4 13 14 15 2
19 15 4 13 0 2 16 16 4 15 10 0 9 9 13 13 1 9 11 2
64 3 16 4 9 1 11 13 1 10 9 1 9 0 9 7 13 10 0 9 2 0 1 9 10 0 9 1 9 11 2 11 7 11 7 11 7 11 1 0 9 7 9 2 0 1 0 7 0 9 2 4 13 11 1 11 7 0 9 1 11 14 4 13 2
19 9 1 11 15 4 13 0 9 1 14 12 9 9 10 2 0 2 9 2
7 3 4 13 12 9 12 2
8 9 15 4 13 1 0 9 2
18 0 9 4 13 3 1 15 7 3 4 15 13 9 1 11 7 11 2
18 3 4 15 13 1 9 7 13 2 16 4 1 11 9 13 1 9 2
5 13 4 0 9 2
3 10 9 2
8 7 3 14 4 13 10 9 2
12 9 12 4 13 0 1 0 9 1 9 9 2
21 0 9 1 0 9 12 9 13 0 1 11 11 2 12 2 12 2 7 10 9 2
14 1 10 9 4 0 9 1 10 9 3 13 0 9 2
26 0 9 1 9 9 15 4 13 2 16 4 13 1 9 12 7 12 0 1 11 0 9 11 2 11 2
15 3 4 13 3 13 7 13 9 1 0 9 7 0 9 2
10 11 13 3 12 9 0 9 7 9 2
16 9 2 11 7 11 13 14 12 1 12 9 1 9 7 9 2
31 11 13 9 2 16 13 9 7 1 15 0 0 9 2 0 9 1 9 9 1 0 9 9 7 0 9 7 9 9 9 2
25 1 0 0 9 13 15 1 9 1 9 9 1 9 1 0 0 9 0 1 9 7 9 10 9 2
20 2 13 2 16 13 10 9 9 0 13 0 9 7 9 9 9 2 16 15 13
12 2 13 9 9 7 13 1 9 1 0 9 2
7 9 9 9 13 3 0 2
9 1 0 15 13 1 0 7 0 2
13 2 13 9 7 9 9 3 0 2 0 7 0 2
16 9 2 9 2 9 2 7 2 9 2 13 3 0 3 3 2
11 9 7 9 15 3 13 1 9 7 9 2
39 9 0 9 1 9 9 15 13 2 1 15 7 13 14 9 9 1 9 3 3 0 2 16 1 0 9 13 1 9 7 9 9 9 2 16 13 0 9 2
8 13 9 9 1 10 0 9 2
13 13 0 0 9 9 2 16 13 0 0 9 9 2
16 16 13 0 9 2 15 13 1 10 9 16 15 13 9 11 2
35 9 9 13 3 2 16 13 10 0 0 9 9 7 9 2 0 9 1 9 11 2 7 13 9 9 2 16 15 13 7 3 13 9 9 2
12 1 10 9 13 13 0 9 1 0 9 9 2
28 9 9 15 1 10 9 13 1 9 0 9 2 16 13 1 9 9 7 9 9 2 16 13 0 1 9 11 2
14 9 9 12 13 3 0 9 9 7 3 13 9 9 2
14 16 13 0 0 9 9 2 15 3 13 14 0 9 2
32 9 1 9 2 16 15 4 9 0 9 13 1 0 9 2 7 13 0 9 9 9 1 11 2 16 13 3 12 9 0 9 2
27 1 9 9 4 16 9 10 9 13 9 1 9 9 2 9 4 15 7 13 9 7 4 13 3 0 9 2
20 13 7 4 14 9 2 16 4 15 0 13 9 9 7 16 13 14 13 9 2
30 7 4 15 3 3 13 2 16 0 9 2 16 15 3 13 1 10 0 9 2 13 9 2 16 4 15 3 3 13 2
26 1 0 9 4 13 9 9 7 3 9 9 13 2 16 13 9 0 7 16 15 13 1 15 3 13 2
17 11 2 9 2 16 4 13 0 9 2 4 3 13 9 11 11 2
20 15 4 14 13 1 11 11 7 11 11 2 11 11 7 4 9 13 1 9 2
13 3 15 1 0 9 1 11 13 0 9 2 2 2
10 1 9 4 15 0 9 13 3 13 2
10 13 4 2 16 15 13 13 0 9 2
13 15 15 4 13 10 9 1 9 9 7 0 9 2
31 2 15 13 11 11 2 2 4 13 1 10 9 7 3 15 15 4 13 9 9 2 16 4 1 9 13 0 2 0 9 2
18 7 16 4 13 14 9 3 2 4 3 13 2 16 9 13 10 9 2
9 7 9 1 15 14 4 13 9 2
4 14 4 13 2
35 1 9 9 2 16 13 7 9 9 16 9 9 1 10 9 2 13 9 9 7 9 2 3 7 15 3 13 1 9 2 16 15 13 9 2
12 0 9 15 9 7 0 9 13 9 0 9 2
23 0 7 0 9 4 15 1 0 9 13 3 16 3 2 7 14 3 4 13 9 3 0 2
18 0 9 0 9 15 3 13 2 7 15 0 0 9 14 4 13 13 2
14 13 4 15 1 0 9 1 11 10 9 1 0 9 2
8 13 4 3 0 7 0 9 2
30 13 15 4 2 16 13 9 3 0 7 15 3 3 16 9 1 9 1 9 13 2 16 1 10 9 13 0 0 9 2
18 13 4 0 2 16 13 0 9 2 7 4 13 2 16 13 0 9 2
23 13 15 4 2 16 4 2 10 10 9 2 1 0 0 9 13 13 0 9 1 12 9 2
27 13 4 14 2 16 4 1 0 9 1 10 0 9 11 13 12 9 7 16 1 15 4 13 14 0 9 2
10 16 4 15 13 2 4 13 1 9 2
8 0 4 13 7 13 0 9 2
29 1 9 4 13 10 9 7 15 13 2 16 4 13 0 7 16 15 15 14 4 13 13 7 13 2 16 15 13 2
9 13 4 0 2 16 4 4 13 2
16 11 3 4 13 15 13 3 2 16 4 0 9 13 1 9 2
17 1 9 15 3 13 1 9 7 13 2 16 15 9 10 9 13 2
8 16 15 3 12 1 0 13 2
28 0 13 2 16 15 4 10 9 13 14 15 1 9 2 16 13 1 9 14 15 2 15 15 15 3 13 2 2
25 1 9 4 13 3 0 9 11 2 16 4 15 3 13 7 13 1 11 7 11 7 14 1 11 2
14 11 7 13 1 3 0 9 9 2 16 13 3 3 2
12 11 13 7 0 9 12 1 0 9 1 9 2
24 13 2 16 13 9 14 0 2 7 0 9 13 2 16 15 9 9 13 1 9 2 9 2 2
30 1 0 9 2 16 13 9 2 0 9 2 7 0 0 9 2 0 9 0 9 14 13 2 7 13 7 15 14 13 2
19 9 13 3 1 9 0 14 1 0 9 2 9 7 0 9 9 7 9 2
27 14 3 7 13 14 0 2 16 4 1 0 9 2 16 4 15 9 13 3 1 9 2 13 1 0 9 2
16 2 1 9 1 0 1 0 9 9 13 0 9 7 13 9 2
9 9 13 3 0 1 9 16 9 2
23 2 0 9 14 13 1 9 9 2 7 15 14 2 15 3 13 3 7 13 1 9 3 2
25 1 9 2 16 15 3 13 1 1 15 0 9 2 10 0 9 13 1 9 7 1 9 1 9 2
56 1 9 7 4 13 14 14 10 9 2 16 14 13 3 0 2 3 13 2 16 13 0 15 2 16 13 3 1 15 9 2 16 15 1 10 9 7 9 13 2 1 9 7 9 13 9 7 15 3 13 2 16 13 15 0 2
19 15 9 13 2 16 15 3 13 7 15 1 9 13 9 9 7 9 9 2
9 1 15 14 4 11 3 3 13 2
26 1 9 4 3 13 11 7 13 2 16 15 13 1 11 2 16 13 10 9 3 2 12 12 0 9 2
15 11 4 13 14 0 13 2 7 15 4 13 9 1 11 2
14 14 7 15 4 13 14 0 9 2 9 14 13 11 2
21 13 15 4 14 1 0 9 2 16 9 14 4 13 2 16 4 13 15 1 11 2
28 1 0 9 0 9 4 15 3 13 2 16 15 9 1 3 0 0 9 3 13 1 9 9 1 9 0 9 2
27 7 14 16 13 1 0 9 2 13 0 13 10 0 9 10 9 2 14 3 7 13 2 16 13 10 9 2
5 3 13 1 9 2
13 9 4 13 14 9 9 2 7 14 9 0 15 2
14 15 4 13 1 9 9 11 0 2 16 15 4 13 2
20 13 2 16 4 13 11 2 16 4 13 1 0 9 7 13 3 1 0 9 2
7 9 15 3 13 1 9 2
16 16 15 15 7 15 13 2 3 13 10 9 7 10 9 13 2
15 15 15 13 2 16 3 13 9 2 9 7 0 9 9 2
23 0 0 9 1 9 9 2 9 7 13 15 2 14 3 13 9 7 15 13 1 10 9 2
13 0 0 9 1 9 13 14 3 13 1 10 9 2
11 11 4 13 1 10 12 9 0 7 0 2
14 7 4 1 9 0 9 7 0 9 10 9 13 9 2
29 1 15 4 13 9 2 16 1 9 9 13 14 14 15 2 7 14 9 2 16 4 13 1 9 2 9 7 9 2
9 13 4 9 2 16 4 13 9 2
19 10 9 4 13 1 9 2 16 15 4 14 0 14 3 13 1 0 9 2
8 10 9 1 9 13 3 0 2
27 14 13 13 2 3 4 11 1 11 13 15 2 7 13 9 2 16 15 4 13 0 9 1 0 9 0 2
9 14 4 1 9 11 3 13 15 2
23 0 0 9 2 16 13 0 2 0 9 1 9 2 4 11 3 3 13 1 0 9 11 2
26 0 9 10 9 2 11 2 0 0 9 2 16 13 1 9 2 13 1 0 9 1 9 7 9 11 2
11 1 15 4 9 13 7 13 10 10 9 2
16 13 9 2 16 15 4 13 1 9 7 9 2 16 14 13 2
24 7 13 9 2 3 4 9 2 3 9 10 9 2 3 13 15 2 13 1 9 0 0 9 2
18 14 13 4 15 13 10 0 9 1 0 9 2 1 0 9 2 2 2
20 14 1 0 0 9 4 15 4 13 13 10 9 10 0 2 0 9 2 2 2
14 7 0 9 1 0 9 1 11 13 0 1 10 9 2
15 7 13 10 9 7 10 9 1 15 2 16 15 13 13 2
26 10 9 1 9 13 14 9 1 15 7 1 10 9 2 16 4 13 10 9 7 15 13 1 10 9 2
12 1 15 15 13 2 16 4 3 13 1 9 2
22 1 9 15 13 1 15 1 11 7 10 9 7 15 13 13 2 16 13 10 9 0 2
12 1 0 0 9 4 11 13 9 9 1 9 2
26 0 9 2 9 2 16 13 2 15 2 1 0 9 1 0 9 2 13 1 9 1 9 7 15 13 2
5 3 0 9 13 2
9 14 3 4 13 3 13 0 9 2
26 15 15 4 14 3 13 2 7 0 9 2 1 9 1 0 2 13 7 13 1 0 9 9 0 9 2
20 0 9 2 16 13 0 2 14 13 9 2 0 9 7 13 0 9 10 9 2
32 13 2 16 15 10 9 13 0 9 2 16 13 9 9 0 9 9 2 16 15 14 3 3 13 1 0 9 2 1 10 9 2
14 7 13 0 13 0 9 2 15 13 9 1 0 9 2
30 11 2 9 0 9 1 0 9 11 2 16 4 9 1 9 9 13 12 0 9 2 4 1 9 0 9 11 11 13 2
20 9 4 9 13 2 16 15 13 9 7 15 4 3 1 0 9 13 16 9 2
20 10 9 4 7 1 9 0 9 3 13 2 16 4 0 9 13 3 7 3 2
15 2 15 4 14 13 13 1 0 2 2 4 3 13 11 2
24 7 16 4 11 13 1 9 7 15 13 1 9 2 15 4 13 2 3 15 4 15 14 13 2
36 1 15 2 16 15 4 13 9 7 9 2 4 14 3 13 2 3 13 1 15 2 7 4 13 3 0 1 10 0 9 7 7 1 0 9 2
25 1 0 9 4 1 15 13 14 9 7 16 3 15 4 13 2 3 4 14 3 3 13 0 9 2
17 13 4 1 9 2 15 13 1 0 9 7 15 1 11 13 9 2
7 0 9 4 13 3 0 2
14 11 4 11 13 1 9 2 16 15 4 3 13 15 2
7 3 4 13 1 10 9 2
12 1 9 15 4 13 0 2 0 7 3 0 2
16 11 15 4 13 9 1 9 2 11 7 15 4 13 1 9 2
7 9 4 13 3 1 9 2
15 11 15 4 1 9 0 9 3 13 3 7 15 3 13 2
14 11 4 13 13 0 2 11 11 7 4 3 13 9 2
14 0 9 4 15 3 13 2 7 4 13 1 0 9 2
11 14 16 15 1 9 9 13 1 10 9 2
13 14 13 0 1 1 15 3 3 0 0 0 9 2
23 15 7 13 14 1 9 9 3 0 1 9 2 0 3 13 3 0 0 9 1 3 0 2
21 9 15 14 13 2 16 13 9 1 9 2 16 15 13 0 9 2 13 0 9 2
15 14 7 4 13 0 9 2 15 4 3 3 9 3 13 2
26 7 7 16 4 9 14 3 13 2 16 13 14 1 9 0 2 13 9 2 3 15 4 13 1 9 2
31 9 7 0 0 9 13 3 3 0 1 9 9 2 16 15 13 1 9 2 16 13 1 9 2 7 13 14 1 9 9 2
16 14 13 7 13 2 16 13 9 14 9 2 16 13 10 9 2
17 14 13 3 2 16 15 13 1 0 9 2 16 4 13 1 9 2
15 1 9 15 13 1 9 3 2 16 4 13 1 0 9 2
28 9 1 0 9 2 16 13 1 9 14 12 9 2 4 13 13 1 9 9 12 2 10 9 4 13 1 0 9
28 14 9 14 13 9 9 7 9 10 9 2 16 15 13 1 15 2 13 14 1 10 9 2 16 4 13 9 2
9 1 10 9 13 0 7 0 9 2
3 13 15 2
12 13 15 4 14 14 9 2 9 7 0 9 2
10 0 9 15 13 1 9 9 7 9 2
13 1 10 9 4 13 3 0 0 9 1 9 9 2
15 0 9 13 9 9 2 16 15 14 13 1 9 0 9 2
12 3 13 0 9 2 16 13 9 9 7 9 2
11 16 10 9 13 9 2 13 16 13 0 2
12 0 0 9 7 9 15 13 1 0 0 9 2
14 9 1 12 9 11 13 0 9 2 0 9 7 9 2
12 15 13 1 0 9 7 15 13 1 0 9 2
14 9 1 12 9 11 13 9 1 0 9 1 0 9 2
56 0 9 11 4 13 0 9 2 16 9 2 16 4 1 9 0 9 2 1 15 4 13 9 2 13 9 1 0 9 7 0 9 2 3 1 9 2 16 15 4 13 9 0 9 1 0 9 0 2 3 13 9 3 0 9 2
4 14 15 13 2
17 7 9 0 9 14 13 1 9 2 16 15 9 13 1 10 9 2
7 16 14 13 8 8 9 2
23 9 10 9 1 9 13 1 15 7 10 9 13 8 8 0 9 2 16 15 10 9 13 2
5 15 13 0 9 2
10 15 7 4 13 2 15 15 3 13 2
4 2 13 15 2
9 13 4 15 2 13 15 10 9 2
7 1 9 4 13 15 0 2
19 13 4 7 15 13 7 13 15 15 4 2 16 15 4 1 9 13 9 2
5 13 4 0 9 2
21 13 4 2 16 15 10 9 13 2 15 7 16 4 3 13 10 9 1 9 9 2
14 15 4 13 0 1 10 9 2 16 4 13 0 3 2
25 0 13 14 9 9 7 7 9 9 1 9 1 9 1 10 9 2 16 9 9 14 13 14 0 2
4 15 3 13 2
9 1 15 13 9 10 9 1 9 2
8 3 13 3 2 13 0 13 2
14 16 13 1 12 9 0 2 13 7 3 10 0 9 2
24 1 9 9 1 9 7 9 9 13 0 9 1 9 1 9 0 9 2 16 3 13 0 9 2
12 0 9 4 13 14 3 0 16 9 1 9 2
12 0 0 9 13 9 1 9 7 9 1 9 2
24 9 4 13 0 9 0 0 9 7 0 9 2 3 16 4 15 9 0 9 13 1 9 9 2
18 0 9 4 15 3 13 2 0 1 9 2 16 4 15 13 1 9 2
20 15 4 14 13 2 16 4 3 13 9 2 16 4 13 9 9 1 0 9 2
28 9 9 7 9 15 1 9 4 13 13 14 8 8 1 9 4 12 2 0 11 10 9 13 1 0 9 11 2
19 1 9 15 13 2 16 4 15 1 10 0 9 3 13 10 0 0 9 2
15 1 12 9 9 12 9 12 9 12 4 13 0 0 9 2
21 1 0 9 4 13 0 2 16 4 13 0 9 3 0 7 13 4 9 0 9 2
18 0 9 0 0 9 7 4 13 9 7 3 4 1 9 13 0 9 2
36 9 9 9 12 13 0 1 12 9 2 13 4 7 14 0 2 16 4 13 0 9 9 9 9 11 2 16 15 4 13 1 2 0 9 2 2
21 0 9 4 1 9 0 9 1 0 9 13 9 9 2 7 13 0 9 1 9 2
24 9 13 14 10 9 1 9 7 1 9 0 9 13 2 16 4 9 1 9 11 11 13 3 2
35 15 3 7 4 13 0 9 2 16 4 13 13 15 2 16 4 13 2 16 4 13 1 11 7 3 2 16 15 13 1 9 1 0 9 2
12 9 1 11 11 1 0 1 11 13 14 0 2
32 0 9 7 4 0 9 1 11 11 13 16 0 9 1 9 2 7 14 4 13 0 9 1 0 9 7 15 13 0 1 9 2
39 1 9 2 3 4 11 1 9 11 9 1 11 13 9 1 9 2 4 3 13 0 12 9 2 16 11 14 13 0 1 11 2 7 4 13 12 9 9 2
5 0 15 4 13 2
17 1 12 1 12 9 4 1 9 0 9 1 0 9 13 12 9 2
18 2 15 15 4 13 2 16 15 4 11 13 1 0 11 1 9 12 2
24 0 13 2 16 13 1 10 9 0 3 10 9 2 9 2 9 2 16 13 1 9 7 1 9
23 1 9 4 13 2 16 13 1 9 13 9 11 12 2 15 13 9 1 10 9 7 9 2
20 9 2 3 14 13 10 0 9 2 16 4 9 13 9 9 1 9 0 9 2
19 13 7 3 1 0 0 9 9 1 0 9 2 10 9 13 9 10 9 2
26 1 10 9 7 3 13 0 2 15 4 13 10 9 2 7 9 2 16 13 14 0 9 1 0 9 2
18 0 9 15 13 3 3 1 0 9 7 15 13 0 9 0 3 13 2
3 2 8 2
20 10 9 1 9 13 1 0 9 7 1 15 3 1 0 3 13 1 9 9 2
10 1 9 1 9 15 13 10 0 9 2
14 13 10 9 2 3 7 14 1 9 1 9 13 9 2
12 13 1 9 2 15 1 9 13 7 13 9 2
12 3 3 13 15 2 3 13 0 0 1 15 2
10 13 15 4 13 12 9 1 12 9 2
11 13 4 10 12 9 2 16 4 15 13 2
13 16 4 0 0 0 9 13 0 2 15 3 13 2
8 9 15 4 1 9 12 13 2
13 1 9 1 10 0 9 13 3 13 14 12 9 2
22 13 4 0 1 0 9 1 0 9 2 1 15 15 4 3 7 3 13 9 0 9 2
9 10 0 9 4 13 14 12 9 2
5 15 14 4 13 2
16 15 2 16 13 7 7 15 13 1 10 9 2 4 13 15 2
9 0 4 7 9 13 1 0 9 2
12 10 9 7 9 3 9 13 2 3 2 3 2
11 13 2 16 13 3 0 9 13 10 9 2
15 14 1 0 9 4 10 9 13 13 10 0 9 1 9 2
8 13 4 1 9 1 0 9 2
15 10 9 4 1 10 9 13 2 16 4 14 15 13 0 2
7 13 15 9 1 12 9 2
16 3 4 13 3 0 7 9 4 13 1 10 9 1 0 9 2
25 13 15 15 4 0 2 16 15 4 13 1 10 9 2 16 13 14 3 0 1 9 7 0 9 2
25 1 15 7 15 4 1 9 13 1 3 0 9 7 4 13 1 0 9 13 16 10 7 15 9 2
9 3 15 4 13 0 14 12 9 2
15 3 13 13 9 7 9 14 13 13 3 3 1 10 9 2
13 14 15 13 3 9 13 2 16 13 0 1 9 2
10 1 9 13 3 0 14 9 0 9 2
11 10 9 3 15 13 2 3 7 14 13 2
10 7 13 9 9 14 1 0 9 0 2
42 16 8 15 1 10 9 13 2 16 15 4 1 10 9 13 9 13 9 1 12 2 12 7 12 9 2 15 14 15 14 13 1 15 2 3 4 9 1 10 9 13 2
20 7 4 10 9 13 2 3 15 4 13 1 0 2 7 7 4 13 3 3 2
18 7 4 10 9 13 13 3 1 9 7 7 4 3 13 1 10 9 2
26 0 0 9 1 0 9 0 9 7 4 13 0 11 11 11 2 16 4 1 9 1 12 9 13 11 2
12 14 1 11 7 10 9 14 13 1 9 12 2
20 15 13 9 0 9 2 12 9 2 2 1 15 14 1 9 13 14 0 9 2
11 1 0 11 15 4 13 1 9 0 9 2
14 1 9 13 13 12 12 9 7 15 3 12 9 13 2
7 2 15 7 15 13 9 2
14 1 15 13 15 3 0 9 2 16 14 13 14 3 2
15 15 15 10 9 13 1 15 2 15 7 15 14 13 3 2
12 7 13 2 16 13 0 9 9 15 3 0 2
27 16 4 14 1 12 9 13 1 11 2 15 14 3 3 13 0 7 0 9 2 16 4 15 15 3 13 2
16 3 16 15 3 13 9 2 16 4 15 15 13 1 12 9 2
30 13 14 9 2 16 4 15 15 10 9 3 13 3 0 2 16 7 15 15 3 13 2 13 1 15 10 9 2 9 2
9 15 13 1 0 9 15 3 0 2
82 7 13 0 2 16 9 2 16 4 15 15 13 14 1 0 11 7 16 13 0 1 0 9 2 3 3 13 9 9 2 16 13 1 3 0 9 2 2 4 13 11 11 2 9 9 9 13 2 16 13 0 1 15 2 16 13 1 0 9 7 16 1 10 9 3 13 10 9 2 0 2 0 9 2 10 13 1 9 13 1 15 2
28 14 3 4 13 1 9 0 11 11 2 16 4 15 13 14 0 9 7 15 4 1 0 9 1 9 13 3 2
3 1 9 2
4 15 13 13 2
16 2 13 15 0 2 3 15 13 13 15 2 2 4 13 9 2
7 15 4 14 13 1 9 2
6 11 11 4 13 0 2
33 1 9 9 9 15 4 13 0 2 3 13 1 9 3 0 7 7 13 3 3 0 2 16 15 14 13 15 13 2 4 15 13 2
9 9 1 10 9 4 13 9 15 2
8 13 4 2 16 15 4 13 2
13 13 4 15 3 13 1 10 9 2 3 4 13 2
6 4 15 13 3 0 2
3 16 3 2
28 1 15 13 3 9 1 15 2 16 4 9 3 13 3 1 9 2 7 13 2 16 15 4 0 9 3 13 2
5 15 13 2 13 2
14 9 15 4 13 2 9 15 4 13 16 14 3 14 2
17 13 9 16 9 0 9 2 16 1 15 13 0 2 14 16 13 2
8 13 4 3 2 13 10 9 2
43 7 15 15 13 0 13 9 0 9 14 1 9 2 16 13 2 0 9 2 2 2 0 9 2 2 16 13 0 2 16 13 0 2 9 2 7 2 9 2 1 10 9 2
14 10 10 9 1 10 9 14 4 13 2 16 13 0 2
24 13 15 14 15 2 16 4 10 9 13 7 13 7 16 4 3 13 3 0 0 9 7 13 2
13 7 1 9 9 9 1 0 12 0 9 13 3 2
7 10 9 13 0 1 15 2
10 10 9 13 11 11 2 11 13 9 2
12 13 14 9 2 16 3 13 0 9 7 9 2
11 0 9 1 9 9 7 13 15 3 0 2
17 13 13 2 16 15 10 0 9 1 9 4 13 3 3 16 15 2
13 10 16 9 11 7 11 4 14 13 10 0 9 2
21 1 9 2 16 13 0 1 12 9 2 1 0 9 13 14 9 7 9 0 9 2
23 0 9 9 1 14 12 9 1 10 9 13 13 0 9 1 9 7 1 15 13 0 9 2
18 9 15 4 1 9 0 9 13 9 2 16 15 13 7 15 3 13 2
42 1 9 0 9 1 9 9 0 9 15 3 13 9 12 0 9 2 16 15 15 0 9 3 13 0 13 7 15 13 2 7 13 1 15 1 0 9 2 9 7 9 2
17 13 13 4 15 9 13 3 7 9 4 1 9 13 1 10 9 2
8 15 0 4 11 13 1 9 2
20 7 14 3 2 13 4 2 16 4 15 13 9 2 16 4 13 11 7 9 2
22 11 11 2 16 15 1 9 1 11 3 13 1 0 9 2 13 1 9 9 3 0 2
25 1 15 3 9 9 13 14 3 3 0 16 14 0 9 2 16 4 15 13 1 9 1 0 9 2
20 11 13 0 2 16 13 0 9 2 14 13 7 13 1 15 2 16 13 0 2
16 16 4 13 2 4 1 9 13 13 14 1 9 2 13 0 2
17 3 15 13 13 2 14 13 2 16 1 11 15 14 4 13 0 2
25 1 15 15 15 13 0 2 16 13 1 9 9 2 16 15 4 13 9 2 14 9 9 3 0 2
18 0 9 0 9 1 10 9 14 13 0 1 9 0 9 16 0 9 2
22 0 9 4 13 9 9 1 0 9 9 9 2 15 4 13 11 11 7 11 11 11 2
23 9 14 4 13 3 1 9 0 9 2 0 9 13 3 3 3 1 9 1 9 0 9 2
36 11 2 1 0 9 2 16 4 1 9 13 0 2 0 9 2 2 4 15 13 9 0 0 9 2 16 15 4 3 14 3 3 13 9 11 2
26 9 4 3 0 9 9 1 9 13 1 0 9 0 9 2 1 9 11 7 4 15 15 3 3 13 2
37 0 11 2 0 0 9 1 9 9 1 9 0 11 2 9 2 4 13 9 1 9 2 16 4 15 1 9 1 9 13 9 2 9 7 0 9 2
19 13 2 16 13 9 3 0 2 16 14 13 1 9 2 7 3 3 13 2
25 9 4 13 1 9 2 16 4 15 13 1 9 0 9 2 0 9 11 11 7 0 9 0 11 2
16 0 13 2 16 4 0 9 13 9 10 9 1 9 12 9 2
24 13 4 1 0 0 9 7 1 9 13 9 7 9 2 0 9 7 4 3 13 1 10 9 2
14 3 4 13 12 9 3 2 16 15 4 9 13 9 2
13 1 15 4 13 14 11 2 7 15 4 9 13 2
21 16 4 13 2 4 11 13 1 9 2 3 7 15 4 1 9 13 14 1 15 2
15 3 15 4 13 1 9 2 9 7 15 4 13 1 9 2
30 11 2 1 9 9 0 9 4 15 1 9 1 12 3 1 12 2 0 11 2 16 4 13 1 0 9 2 13 9 2
20 13 4 2 15 13 13 7 15 2 3 2 13 12 0 9 2 9 7 9 2
9 13 4 15 1 3 12 12 9 2
4 13 15 15 2
20 1 9 13 3 0 14 9 9 7 9 9 2 16 15 3 13 1 0 9 2
3 4 13 2
4 15 4 13 2
18 3 15 13 3 13 1 0 9 7 15 3 13 14 1 9 0 9 2
7 14 2 16 13 0 9 2
8 11 7 13 0 2 0 9 2
37 1 9 1 3 0 9 2 16 13 11 7 11 2 13 9 0 9 2 16 15 3 13 1 0 9 7 0 9 2 1 0 9 7 13 3 0 2
14 9 0 9 7 0 0 9 13 1 0 9 0 9 2
7 0 0 9 15 14 13 2
9 9 11 1 15 13 16 0 9 2
20 13 15 2 16 13 1 0 9 2 9 2 9 2 7 1 15 13 15 3 2
14 3 3 13 2 16 9 9 13 16 9 7 0 9 2
18 14 14 13 9 2 7 13 1 10 9 0 1 9 7 1 0 9 2
12 2 13 4 9 2 16 4 3 13 1 0 2
17 1 9 4 13 10 9 16 9 7 14 9 15 4 3 3 13 2
14 0 4 13 2 16 4 1 9 1 9 13 1 9 2
22 0 11 2 9 13 0 2 4 13 14 1 12 9 3 0 2 16 13 0 16 9 2
45 16 15 14 4 9 1 9 9 13 0 9 1 9 9 2 14 14 3 14 4 13 2 16 13 0 2 0 9 2 0 9 11 2 11 2 11 2 16 15 13 14 1 9 11 2
12 11 15 4 13 1 11 1 10 0 9 1 11
9 9 9 9 4 13 0 0 9 2
11 3 7 3 4 9 13 2 9 14 13 2
3 2 8 2
3 2 8 2
13 3 9 0 0 9 1 0 9 13 9 9 1 9
18 3 13 14 12 9 9 2 16 4 15 1 10 9 14 13 1 15 2
33 1 10 9 9 1 9 8 9 14 13 14 9 2 7 15 7 1 0 16 0 9 7 9 9 13 14 0 9 7 9 10 9 2
32 0 0 9 1 12 9 4 3 13 9 1 9 7 9 9 0 2 3 7 4 9 14 1 10 9 13 9 1 0 9 9 2
26 3 4 3 1 10 9 13 9 7 15 14 13 1 10 9 9 2 1 15 4 15 3 13 10 9 2
10 0 9 15 15 13 3 0 7 0 2
23 3 4 13 0 9 2 16 13 11 13 1 10 9 1 9 7 15 15 3 14 3 13 2
15 13 15 2 16 15 4 13 3 3 2 15 13 7 13 2
31 9 7 4 1 9 13 13 9 7 0 9 2 7 15 4 3 13 2 16 4 13 9 7 0 9 4 15 1 9 13 2
28 7 7 15 4 3 13 2 16 13 3 0 7 4 13 2 16 13 11 0 7 4 1 15 13 7 15 13 2
10 14 3 9 4 15 3 13 1 9 2
25 9 4 13 3 2 16 15 15 3 13 1 0 9 7 3 4 13 0 9 7 15 3 14 13 2
7 3 15 13 14 12 9 2
16 1 0 11 4 13 0 0 9 2 9 1 9 7 9 9 2
25 16 9 1 0 9 14 4 13 0 2 4 15 9 1 15 14 3 13 1 0 0 9 7 9 2
38 13 15 2 16 1 9 0 9 13 14 0 9 2 14 16 4 13 14 14 0 2 7 4 15 13 3 0 13 10 0 9 1 10 12 7 15 9 2
12 0 13 14 2 3 15 13 2 13 7 13 2
28 11 15 4 1 9 13 1 0 9 7 1 0 2 3 0 9 4 13 9 13 9 7 15 13 1 0 9 2
11 14 1 12 9 4 13 9 12 0 9 2
10 3 4 13 7 9 15 15 4 13 2
21 9 4 13 13 0 9 2 16 14 4 13 9 7 9 2 16 4 13 15 0 2
14 9 2 16 15 15 4 3 13 2 15 4 13 15 2
10 2 1 9 7 9 13 9 9 9 2
11 13 2 3 13 10 9 0 1 9 9 2
9 1 10 0 9 9 13 0 9 2
10 1 0 9 13 1 0 0 9 1 9
13 1 0 9 13 0 10 9 14 1 9 7 9 2
10 1 9 13 9 3 0 16 1 11 2
11 16 15 13 1 11 2 15 3 13 9 2
9 11 13 10 10 9 3 1 9 2
19 16 14 15 15 13 2 13 15 1 9 2 15 13 1 15 7 15 13 2
15 11 15 1 10 9 13 2 16 4 13 0 1 0 9 2
18 10 9 13 7 13 9 2 16 9 13 2 13 7 0 1 0 13 2
24 9 7 13 7 15 13 2 14 16 4 15 13 2 15 15 13 2 7 4 15 3 14 13 2
25 16 13 9 1 9 0 2 16 13 15 0 2 3 14 13 2 3 4 15 13 2 16 15 13 2
13 0 4 15 13 0 9 2 0 9 7 0 9 2
9 4 13 13 2 15 4 13 13 2
6 15 0 13 0 9 2
24 3 13 2 16 13 1 10 9 3 3 16 9 2 7 14 3 3 13 2 3 10 9 13 2
10 3 3 13 2 3 15 13 1 9 2
9 1 9 13 14 14 1 0 9 2
17 10 1 9 0 9 1 10 9 11 11 3 3 13 9 10 9 2
22 10 0 9 13 10 9 2 7 15 13 14 3 2 16 15 14 13 13 1 10 9 2
17 1 9 4 13 2 16 13 2 15 9 1 9 13 0 9 9 2
26 16 13 9 2 16 13 9 1 9 2 9 2 15 13 3 3 1 9 2 10 4 13 7 13 14 2
29 16 4 9 3 13 2 16 13 2 15 2 16 13 2 2 4 15 3 9 3 13 16 2 15 2 16 13 2 2
24 7 14 10 9 2 10 9 9 2 16 4 1 9 13 10 9 2 15 13 1 9 7 9 2
14 9 9 13 2 1 10 9 15 3 13 14 10 9 2
23 16 3 13 10 9 16 1 15 2 15 13 9 2 16 4 13 0 9 7 15 13 9 2
30 16 13 3 2 16 15 4 13 9 2 15 7 4 13 13 1 9 2 16 13 1 10 9 2 16 4 13 1 15 2
22 15 7 13 2 16 4 13 1 9 0 14 3 2 16 4 1 15 13 9 10 9 2
13 9 1 0 15 13 1 9 2 16 15 15 13 2
14 14 13 9 7 9 2 3 1 12 12 9 4 13 2
25 0 9 15 4 13 9 2 16 4 1 10 9 13 3 0 9 2 16 15 13 0 0 0 9 2
46 10 0 0 9 4 13 0 9 11 11 2 16 4 13 1 0 9 14 14 3 0 1 15 2 16 15 4 9 12 2 14 13 2 1 9 7 4 13 1 15 7 15 4 13 9 2
18 0 9 2 15 15 4 13 1 15 2 13 3 3 9 0 0 9 2
16 1 9 13 9 10 9 2 7 13 13 9 3 2 0 2 2
11 1 15 13 0 13 2 16 9 14 13 2
16 1 10 9 4 1 0 0 9 8 11 9 12 13 0 9 2
14 0 9 1 11 0 9 13 12 0 9 9 11 11 2
4 15 13 9 2
11 13 4 2 16 13 3 0 16 3 3 2
47 9 4 13 0 14 9 1 10 2 0 2 0 9 2 1 15 4 15 13 0 0 9 2 1 9 0 1 0 9 2 15 4 15 0 9 1 9 14 13 7 13 2 3 15 9 13 2
22 1 0 4 13 10 0 9 0 9 2 9 7 0 9 1 9 0 9 11 0 9 2
24 9 2 16 13 1 9 0 9 2 15 13 3 1 15 13 2 13 1 9 15 7 9 9 2
22 14 7 14 10 9 1 10 9 14 13 9 9 9 2 16 13 3 0 1 0 9 2
31 14 13 13 2 16 13 9 9 1 0 9 1 9 0 2 14 16 15 13 16 9 0 9 2 1 15 15 13 0 9 2
31 12 1 10 9 13 14 9 2 16 13 0 14 16 10 9 0 9 2 1 15 15 13 9 0 9 1 9 0 9 9 2
34 14 1 0 9 4 10 12 9 13 14 0 9 1 9 9 0 9 7 10 9 2 7 15 4 1 15 1 15 13 0 9 0 9 2
24 10 10 7 0 9 9 7 9 0 9 4 3 1 0 9 3 13 0 9 7 10 0 9 2
9 0 9 1 15 13 3 0 9 2
42 1 15 15 3 0 9 13 14 14 16 0 9 2 7 14 16 9 2 16 1 2 9 9 2 13 16 3 0 9 10 0 9 2 16 4 15 13 1 0 0 9 2
48 1 9 9 2 16 15 3 13 2 13 14 13 2 16 13 9 10 9 1 9 0 9 3 0 7 16 10 9 3 13 3 0 9 2 16 3 13 3 1 0 7 0 9 9 1 0 9 2
46 0 9 0 9 1 0 9 13 0 1 9 2 15 13 0 9 0 7 0 9 2 16 13 1 0 2 0 2 9 7 9 1 0 9 7 10 10 9 0 9 13 0 9 0 9 2
12 10 9 13 3 13 9 1 9 2 9 9 2
51 11 11 2 0 13 10 9 2 16 4 1 10 12 0 0 9 1 9 2 3 0 9 2 15 1 9 13 10 9 2 7 0 9 9 11 11 11 4 13 15 2 16 0 9 1 11 11 13 10 9 2
31 16 4 11 11 2 11 11 7 11 11 3 14 13 1 0 9 2 13 14 11 13 10 9 12 9 1 9 1 10 9 2
21 2 16 15 15 13 13 12 9 2 4 13 0 9 2 2 13 0 9 1 9 2
30 1 9 4 15 14 3 3 13 9 9 9 2 16 7 15 13 2 15 13 13 2 16 15 9 14 4 13 0 9 2
52 14 13 3 0 1 0 9 2 16 4 1 9 1 11 0 13 9 0 9 1 0 9 1 0 9 1 11 11 11 7 0 9 1 9 1 11 11 11 2 10 9 4 13 9 11 11 1 11 11 11 2 2
13 7 15 13 1 9 0 9 1 9 11 11 11 2
20 13 4 1 9 0 9 2 11 2 9 0 9 7 0 9 1 11 11 11 2
4 1 11 13 2
13 0 0 9 13 0 7 0 9 13 10 9 3 2
7 1 11 4 3 14 13 2
39 3 4 13 1 0 2 0 9 10 0 9 1 9 1 0 7 0 9 2 3 15 13 1 9 2 16 15 9 3 3 13 7 1 9 13 1 0 9 2
25 9 9 13 1 0 11 2 7 16 1 3 13 9 2 15 13 2 16 15 1 9 13 1 9 2
14 7 13 3 2 16 13 1 0 9 1 9 1 9 2
12 3 15 14 4 14 9 13 1 10 0 9 2
8 13 1 9 9 7 9 13 2
24 1 0 9 2 16 4 12 9 12 3 13 0 9 11 11 1 11 2 4 1 9 14 13 2
16 3 4 13 10 9 7 0 2 16 13 9 11 1 0 9 2
9 13 4 15 14 10 0 0 9 2
30 3 3 15 4 9 9 13 0 9 11 2 16 4 13 14 12 10 9 2 16 4 1 10 9 13 1 9 0 9 2
26 1 10 9 4 13 2 3 0 13 0 9 7 9 0 7 14 0 9 2 16 9 13 13 0 9 2
30 1 12 9 4 13 13 3 0 0 9 2 16 1 10 9 11 13 0 9 9 2 9 7 0 9 9 7 9 9 2
12 1 11 4 9 13 3 3 7 15 14 13 2
45 9 1 9 2 9 7 9 8 11 11 4 9 13 0 9 1 0 9 7 9 0 9 2 16 11 3 13 0 9 2 16 13 0 9 9 2 3 7 13 0 9 0 0 9 2
17 9 9 7 9 2 9 7 9 2 13 0 9 1 0 0 9 2
24 14 10 9 13 9 9 0 9 2 16 13 9 0 9 2 9 2 9 0 9 7 9 9 2
52 9 11 4 13 2 16 14 3 1 15 2 3 4 3 13 0 9 0 9 9 2 1 15 4 0 9 14 13 10 9 2 4 9 13 1 15 2 16 4 0 9 9 7 9 13 9 9 14 1 0 9 2
26 0 9 7 9 7 0 9 13 9 2 16 13 0 9 2 9 7 13 14 9 9 1 0 0 9 2
11 13 15 10 12 9 1 9 9 0 9 2
42 14 4 13 9 7 9 1 9 0 9 1 0 9 9 2 7 4 14 3 13 9 2 16 13 1 9 0 9 2 16 13 9 1 9 14 0 0 9 13 14 9 2
29 15 7 13 2 16 9 2 16 13 9 2 14 13 13 10 0 9 2 16 15 13 1 9 0 9 1 0 9 2
36 1 9 1 0 9 7 9 2 16 13 9 0 9 1 0 0 9 2 13 2 16 15 4 3 13 1 9 1 9 0 9 7 13 14 9 2
17 16 13 2 4 10 0 9 14 13 0 9 1 9 0 0 9 2
31 13 14 0 9 1 0 0 9 0 9 2 16 13 10 9 2 9 9 2 0 9 1 9 7 9 1 0 9 2 9 2
13 3 13 9 9 14 13 9 0 9 1 0 9 2
14 1 15 4 13 3 3 0 2 15 13 14 0 9 2
32 14 12 0 9 7 10 12 9 7 12 0 0 9 1 12 9 13 9 0 9 0 9 11 2 9 11 7 9 11 1 11 2
21 16 4 13 9 9 2 16 15 13 0 9 2 4 13 0 9 0 9 0 9 2
20 3 3 3 7 15 0 9 13 14 1 9 9 7 14 3 13 13 0 9 2
39 15 3 13 2 16 13 1 9 12 9 3 2 13 2 9 7 9 1 0 9 2 3 3 3 10 9 7 9 13 10 0 9 2 14 13 9 9 2 2
20 1 9 4 13 0 9 9 0 9 2 16 13 1 9 2 16 13 9 0 2
18 9 4 13 10 0 9 1 9 2 9 7 9 9 2 0 1 9 2
8 3 7 10 9 13 1 9 2
7 10 0 9 13 14 9 2
25 13 3 9 9 7 9 7 15 13 1 9 1 9 9 2 16 15 13 10 16 12 9 10 9 2
13 3 13 0 9 7 9 2 16 15 13 0 9 2
15 3 13 9 2 16 15 13 1 0 9 1 9 0 9 2
17 3 13 15 3 9 1 0 9 2 1 9 1 10 16 12 9 2
20 1 9 9 13 9 3 0 0 9 9 2 16 13 14 3 0 1 12 9 2
30 0 9 2 16 4 15 15 13 1 12 1 9 2 13 3 2 3 13 9 14 1 9 2 16 15 9 14 13 14 2
12 0 9 13 1 9 2 1 15 0 9 13 2
28 0 9 9 13 3 2 16 15 13 9 2 9 9 2 9 7 0 9 2 16 15 13 0 13 1 0 9 2
21 2 13 2 16 13 0 1 10 0 9 2 1 15 10 9 3 13 1 0 9 2
16 0 9 1 9 9 7 9 1 9 9 13 9 9 0 9 2
4 0 9 13 2
15 3 13 3 14 9 2 16 13 13 0 9 9 2 13 2
21 0 9 9 1 9 1 9 9 13 2 16 9 13 1 9 7 9 13 16 9 2
21 16 13 9 2 13 9 7 9 13 2 14 16 4 13 1 15 13 0 0 9 2
15 1 0 11 3 13 1 9 1 0 0 9 1 0 9 2
18 9 9 4 13 3 0 1 9 1 10 0 9 1 0 9 12 9 2
12 3 13 14 0 9 0 9 1 0 0 9 2
27 16 13 14 9 7 9 2 3 1 9 9 13 0 9 2 16 13 2 16 15 4 0 9 13 1 9 2
14 1 0 9 1 0 0 9 13 1 9 3 1 11 2
19 13 0 0 9 2 14 12 10 9 13 0 9 9 1 9 1 0 9 2
13 1 0 9 0 11 13 0 7 15 0 0 9 2
21 1 9 11 13 0 0 0 9 2 1 15 15 3 13 1 10 9 0 0 9 2
17 0 9 15 13 3 1 9 2 13 0 9 7 15 13 1 11 2
11 1 9 4 13 7 9 0 9 9 9 2
21 1 10 9 4 1 11 14 13 0 9 2 16 7 4 13 14 1 9 3 0 2
15 3 13 10 9 9 9 14 14 9 1 3 3 0 9 2
41 9 0 0 9 4 1 9 9 0 9 1 0 7 0 9 9 7 1 9 0 9 1 10 9 9 12 3 13 9 2 1 15 14 10 9 13 9 7 13 9 2
9 13 15 9 10 9 1 9 11 2
15 1 9 15 13 14 0 9 1 0 9 7 9 0 9 2
17 1 3 15 13 1 9 1 0 11 2 16 0 9 13 10 9 2
11 15 1 0 9 3 13 0 9 0 9 2
15 0 9 9 2 9 2 15 1 0 9 3 13 7 13 2
4 15 15 13 2
19 1 15 1 3 0 9 13 0 9 7 9 1 9 3 2 16 13 0 2
12 1 9 15 1 9 9 13 9 2 9 2 2
14 14 2 13 10 0 9 2 3 13 3 13 0 9 2
25 0 13 14 2 16 15 2 16 13 2 13 1 9 14 3 16 3 7 13 0 9 1 0 9 2
27 9 14 3 13 7 3 14 4 1 9 13 2 14 16 15 14 13 13 1 3 15 2 15 15 9 13 2
26 0 9 1 9 9 9 1 9 4 13 1 9 11 2 1 9 11 11 11 11 7 10 9 11 11 2
20 1 0 9 9 9 7 1 0 0 9 3 13 10 16 12 9 10 0 9 2
25 3 13 14 9 9 1 9 2 0 9 2 11 2 2 16 13 1 9 9 7 0 9 0 9 2
24 11 11 1 9 11 4 1 10 0 9 13 2 16 13 9 9 3 0 1 9 7 0 9 2
20 1 9 9 3 13 2 15 13 0 9 2 16 13 9 0 7 14 0 9 2
21 0 13 2 16 13 9 1 0 9 1 9 10 9 3 0 2 13 7 0 11 2
15 10 9 3 13 14 16 0 9 1 9 7 9 1 9 2
14 9 13 1 0 9 2 16 15 13 2 3 15 13 2
7 2 1 0 14 4 13 2
15 3 0 9 2 16 15 13 11 3 2 14 3 4 13 2
24 16 13 3 10 9 3 13 1 9 2 4 15 3 1 9 11 13 2 16 4 13 3 3 2
23 0 9 4 14 3 3 13 9 9 1 10 9 2 7 15 3 4 13 9 1 0 9 2
22 0 0 9 4 3 7 3 13 3 3 0 9 2 16 3 3 13 9 1 0 9 2
15 9 1 9 7 0 9 4 13 0 9 0 2 9 2 2
10 14 3 15 15 13 10 0 9 9 2
11 11 13 3 3 0 9 1 0 0 9 2
17 3 0 9 13 3 12 9 2 16 4 15 13 1 9 7 9 2
24 9 0 9 13 3 14 1 9 2 9 1 10 9 2 0 1 0 9 2 7 3 13 9 2
20 1 15 2 16 13 10 9 2 4 1 9 13 12 9 2 16 15 3 13 2
23 1 10 9 15 3 15 13 2 9 2 1 9 2 16 15 13 0 13 14 1 10 9 2
38 3 15 9 3 13 13 2 1 10 9 14 13 0 2 0 13 14 2 16 9 2 16 13 1 9 2 13 2 16 4 13 0 9 10 7 15 9 2
27 11 3 15 4 13 1 15 2 16 13 1 9 0 2 16 13 2 3 2 7 16 14 13 1 9 9 2
12 0 3 0 0 9 15 4 13 9 1 9 2
18 9 13 2 16 13 1 9 2 1 15 7 10 9 13 9 10 9 2
13 3 13 2 16 15 13 9 7 0 9 1 12 2
19 14 13 1 9 2 16 15 13 1 9 2 16 4 14 13 1 15 9 2
6 0 9 13 9 9 2
18 0 9 13 1 9 2 13 0 9 7 15 3 13 2 16 14 13 2
20 13 9 9 2 16 4 15 3 13 1 9 2 7 15 13 2 16 14 13 2
14 13 0 9 9 2 9 2 9 2 0 9 7 9 2
15 13 2 16 13 2 3 7 13 1 9 2 0 1 9 2
17 1 9 13 9 2 13 0 9 7 9 7 9 13 1 0 9 2
14 9 1 9 7 1 9 3 4 13 9 14 0 9 2
14 16 4 13 9 2 4 1 9 1 15 13 0 9 2
17 9 1 11 4 11 3 13 2 3 3 0 11 13 1 9 7 9
19 0 9 0 9 4 9 14 0 9 3 13 0 9 9 1 9 7 9 2
13 1 9 9 1 9 11 4 11 3 13 0 9 2
23 1 12 0 9 15 4 3 3 13 1 12 9 2 0 7 13 14 9 0 9 7 9 2
33 1 12 1 12 9 1 9 2 7 9 2 13 10 9 9 2 16 4 15 13 1 12 9 0 9 2 16 4 3 13 10 9 2
23 0 9 7 13 9 9 2 9 1 9 7 0 9 2 16 9 13 2 16 15 9 13 2
17 10 9 15 4 13 2 16 4 13 3 7 15 1 9 13 9 2
6 15 15 4 13 13 2
20 9 4 15 3 13 2 16 13 9 10 0 9 14 0 9 2 16 13 9 2
13 13 4 16 9 2 16 1 9 13 15 1 15 2
6 3 7 4 13 9 2
14 4 15 13 1 0 2 0 9 2 16 13 1 9 2
11 1 0 4 14 3 13 7 13 1 9 2
18 13 4 9 1 15 2 7 3 4 3 13 2 16 9 4 13 0 2
12 7 15 4 13 0 9 2 16 4 15 13 2
25 13 4 9 2 16 3 4 13 10 9 2 7 15 4 13 2 16 16 13 10 9 1 10 9 2
11 4 13 0 2 0 9 2 3 13 0 2
24 13 4 0 2 0 2 0 9 2 16 4 13 2 16 15 3 13 9 2 16 13 0 9 2
10 1 0 12 9 4 13 1 12 9 2
16 3 4 13 3 0 2 3 4 1 12 0 9 13 12 9 2
9 9 4 13 13 10 2 9 2 2
27 0 9 13 0 9 2 16 13 0 13 10 9 3 2 16 4 14 1 9 9 1 9 13 2 16 13 2
16 9 14 4 13 10 9 7 13 1 0 9 0 9 7 9 2
13 1 15 14 4 15 13 14 9 1 9 0 9 2
6 2 13 0 16 9 2
5 13 3 7 3 2
12 3 15 14 13 2 16 16 4 13 1 9 2
8 1 9 13 1 9 7 9 2
10 9 15 13 0 1 0 9 7 9 2
10 9 15 1 9 14 4 13 0 9 2
8 1 9 13 15 0 7 0 2
4 15 13 9 2
24 15 13 14 10 9 7 3 13 9 1 9 2 9 13 14 3 0 1 15 7 15 3 13 2
14 16 13 9 0 2 15 1 12 9 14 13 10 9 2
9 9 9 1 10 9 14 14 13 2
17 16 7 13 10 9 3 13 14 9 2 16 13 9 0 7 0 2
25 13 7 13 2 16 9 3 3 13 0 9 7 16 15 13 3 0 0 9 9 16 7 0 9 2
4 9 13 0 2
15 15 13 9 9 2 9 2 9 2 9 1 9 2 2 2
12 3 4 15 13 2 16 15 13 1 0 9 2
13 1 9 4 15 13 16 0 7 15 13 0 9 2
12 7 14 14 15 13 2 16 10 9 13 0 2
19 9 9 9 11 2 11 11 2 7 15 4 13 2 16 14 13 0 9 2
15 11 11 15 4 13 9 12 1 9 0 9 1 0 11 2
22 9 1 15 4 13 4 14 13 10 9 1 0 2 0 2 0 2 0 7 0 9 2
17 1 15 15 4 13 1 9 1 0 9 1 9 2 9 7 9 2
21 1 0 9 4 14 9 12 13 9 0 9 9 2 0 9 4 13 9 9 11 2
13 9 12 4 13 9 9 9 7 9 1 0 11 2
21 1 9 9 12 7 4 13 0 9 9 0 2 0 7 0 9 0 9 0 11 2
13 2 9 13 9 9 10 9 2 9 9 0 9 2
11 7 16 13 0 2 3 14 15 0 13 2
19 15 14 4 13 13 1 15 2 15 13 0 1 0 9 2 2 13 11 2
14 12 9 1 11 13 3 0 9 9 11 7 9 11 2
21 2 0 9 10 0 9 13 12 9 0 9 2 1 15 4 1 9 13 12 9 2
28 9 13 0 3 2 16 15 4 13 1 0 9 3 12 2 0 9 7 4 3 3 3 10 9 3 13 0 2
50 16 15 3 13 2 16 13 10 0 9 2 1 9 15 15 9 3 1 9 13 1 9 2 0 1 11 2 15 4 13 2 16 9 9 7 13 15 2 16 15 1 15 14 4 13 14 9 1 9 2
29 3 3 0 13 14 0 9 2 7 4 10 9 13 9 10 9 2 1 15 1 7 1 9 13 10 3 0 9 2
26 0 9 9 2 16 4 15 1 3 9 7 3 10 0 9 13 0 9 2 13 14 0 9 1 9 2
24 1 9 4 13 14 12 9 0 0 9 2 1 15 15 3 10 9 1 9 3 13 0 9 2
15 12 9 9 12 15 4 1 9 0 9 9 13 3 3 2
35 9 9 13 2 16 9 9 14 13 1 0 9 1 9 2 14 7 1 9 13 15 2 15 14 4 13 10 0 9 7 15 13 0 9 2
32 1 15 13 9 0 7 0 1 15 3 0 7 1 10 9 13 0 9 3 10 9 7 3 3 0 0 9 2 9 7 9 2
30 9 9 2 9 2 13 1 12 9 0 9 7 0 9 2 1 0 9 14 10 9 0 15 13 1 0 9 7 9 2
10 6 2 16 13 0 1 10 0 9 2
4 9 1 9 2
8 13 4 15 0 9 9 12 2
12 1 11 11 4 13 1 9 12 1 9 12 2
17 9 4 13 0 1 9 11 2 15 7 4 13 1 9 9 11 2
21 9 11 15 4 13 9 1 9 1 11 2 3 4 13 13 9 1 9 11 11 2
14 13 4 0 2 0 9 2 9 2 9 7 10 9 2
10 0 9 1 9 7 9 13 14 0 2
36 1 0 0 9 0 9 11 4 15 13 9 9 2 16 14 4 15 4 12 9 1 9 11 3 3 13 2 16 4 1 9 13 1 0 9 2
5 0 9 4 13 2
12 1 9 13 9 0 9 7 1 9 0 9 2
27 3 4 15 13 14 9 1 9 1 9 9 1 0 9 2 1 15 4 13 0 13 14 10 9 1 9 2
9 7 1 9 13 7 9 7 9 2
6 15 13 3 0 9 2
24 1 9 11 11 2 9 9 0 9 2 4 15 3 13 11 2 16 15 4 13 1 0 9 2
39 2 9 9 13 3 13 2 2 4 13 11 7 13 2 16 13 9 1 9 3 0 14 3 2 16 15 1 9 13 0 9 2 16 13 9 1 0 9 2
11 11 14 4 4 12 1 9 13 1 9 2
22 13 4 14 14 0 9 9 7 9 1 9 13 2 15 13 7 13 2 16 11 13 2
17 12 1 9 15 4 7 13 13 1 9 7 11 4 13 13 3 2
21 3 14 4 15 4 1 15 13 11 7 15 13 1 9 13 0 9 7 15 13 2
9 9 4 15 13 7 13 1 9 2
4 13 4 9 2
31 0 4 15 13 1 9 7 1 0 9 14 4 4 9 13 2 3 7 15 3 13 7 13 2 16 4 9 13 0 9 2
17 1 9 4 13 11 7 11 2 16 14 4 4 1 15 13 9 2
11 10 12 9 4 13 9 1 9 1 9 2
5 9 9 14 13 2
21 13 7 2 16 4 9 13 1 10 9 7 15 1 10 9 13 14 9 1 9 2
19 11 14 13 2 16 14 4 15 4 9 1 9 0 13 1 9 7 9 2
23 13 10 9 2 14 16 14 4 4 9 13 14 2 16 4 13 9 14 0 1 0 9 2
17 2 8 8 4 1 9 3 13 2 16 4 13 1 0 9 2 2
8 1 3 15 13 0 0 9 2
30 16 14 4 13 15 1 0 9 12 0 0 9 1 9 1 0 9 2 13 14 0 2 16 9 9 9 14 4 13 2
9 14 3 16 13 1 11 9 9 2
29 7 16 4 1 0 13 0 9 2 3 16 4 9 10 9 3 13 9 2 4 3 0 9 11 3 13 1 9 2
44 16 15 0 0 9 1 9 14 4 13 10 9 7 13 1 9 10 9 2 14 16 4 11 13 13 1 9 1 9 2 3 13 11 11 0 2 16 4 13 10 9 1 11 2
12 7 4 1 10 0 7 0 9 13 1 9 2
38 0 11 7 11 4 15 13 1 9 1 0 7 0 9 1 9 1 11 2 16 4 3 13 10 9 1 0 9 2 7 1 0 0 9 0 0 9 2
22 3 13 0 9 0 9 9 1 9 2 0 11 7 4 3 3 13 9 0 9 9 2
34 11 2 9 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 2 11 7 11 2 13 9 0 9 1 9 11 11 2
8 0 9 15 13 9 0 9 2
17 1 0 9 12 9 15 9 2 9 9 2 9 2 9 2 13 2
10 9 14 3 13 0 9 1 9 9 2
28 14 15 7 13 2 16 1 10 9 13 3 0 0 9 2 7 15 4 14 14 3 15 13 1 9 0 9 2
7 13 1 10 9 9 9 2
11 1 9 13 3 2 16 13 9 1 15 2
9 1 9 13 3 7 13 1 9 2
24 15 13 12 2 16 9 13 1 9 7 16 15 13 2 16 15 13 13 2 13 3 1 3 2
6 15 15 13 1 9 2
11 3 13 14 12 9 13 10 9 14 0 2
17 0 9 9 13 0 13 3 2 16 4 13 10 9 3 12 9 2
9 13 4 10 9 1 11 7 11 2
4 3 3 13 2
13 9 13 0 3 3 16 0 9 1 9 10 9 2
20 9 9 7 9 1 9 4 13 3 14 0 1 0 9 2 7 9 7 9 2
34 16 9 2 16 15 4 1 9 13 11 11 2 13 1 3 2 3 14 13 13 2 3 15 4 13 9 7 0 9 1 9 9 9 2
20 1 11 4 14 13 1 9 10 0 0 9 13 2 16 13 10 9 13 0 2
26 11 4 13 0 9 1 10 0 9 2 16 13 9 9 0 9 1 9 1 9 9 7 0 9 9 2
22 9 13 14 1 0 9 2 7 13 15 3 0 7 3 0 1 0 9 1 0 9 2
7 13 7 3 3 0 9 2
21 9 15 0 0 9 13 9 11 2 7 15 1 9 9 1 9 3 3 14 13 2
8 9 15 13 3 7 3 3 2
31 1 9 15 13 2 16 14 1 12 9 14 13 3 3 13 9 16 1 10 9 2 15 13 1 9 14 1 9 7 9 2
8 1 0 9 9 3 14 13 2
26 0 7 13 14 9 9 2 7 14 3 0 9 2 16 13 13 9 1 0 9 9 9 7 0 9 2
15 1 9 1 0 9 1 9 15 9 3 9 13 3 3 2
17 1 9 13 15 3 0 9 0 9 2 16 4 13 0 0 9 2
16 15 4 13 0 2 4 14 13 10 9 7 9 13 1 15 2
11 3 3 13 1 9 2 16 13 1 9 2
14 15 15 1 10 9 7 9 14 14 14 13 10 9 2
35 14 3 0 13 2 16 15 9 0 9 3 13 2 3 7 15 14 0 9 1 10 9 7 9 13 7 1 15 14 13 9 9 7 9 2
46 0 0 9 2 16 4 3 13 11 13 3 1 9 7 9 11 11 11 14 10 0 9 2 16 4 13 10 0 9 0 9 2 10 0 2 0 7 0 9 7 4 13 1 15 0 2
13 1 15 13 14 0 9 2 10 13 0 0 9 2
8 15 13 3 0 2 3 2 2
12 15 13 1 10 0 9 2 13 1 0 9 2
14 9 11 4 13 2 16 1 9 4 15 14 13 13 2
11 13 4 2 16 13 10 0 9 7 9 2
33 11 2 9 1 0 9 7 0 9 4 1 9 9 8 7 1 9 0 9 3 1 0 9 11 13 9 1 9 0 9 7 11 2
21 9 4 13 1 15 3 3 0 1 11 2 11 2 11 2 1 0 11 7 11 2
9 13 4 15 1 3 12 9 9 2
25 1 0 9 12 9 4 15 9 3 13 2 1 0 0 9 7 4 15 9 1 9 9 3 13 2
29 1 9 4 15 13 0 9 0 9 2 3 7 4 1 9 0 9 13 0 9 2 16 13 0 9 2 9 2 2
18 1 11 15 9 3 13 1 9 2 9 2 0 9 7 10 0 9 2
20 0 13 1 0 9 2 9 2 0 9 1 9 2 9 2 9 2 0 9 2
18 16 4 14 13 11 11 2 0 9 1 0 9 13 1 9 10 9 2
36 2 13 2 16 13 3 2 16 3 13 9 0 9 2 16 4 14 9 12 13 10 9 9 1 9 2 16 13 0 9 2 0 1 9 9 2
27 1 9 9 7 9 9 1 9 4 9 13 14 3 2 16 4 13 15 9 0 9 1 0 9 0 9 2
21 1 10 9 13 9 0 9 1 9 9 0 2 7 4 0 0 9 13 0 9 2
33 9 1 9 4 3 1 9 9 2 9 7 0 0 9 1 0 9 7 1 0 9 1 9 0 9 7 0 9 13 12 9 9 2
10 9 10 9 4 13 0 9 7 9 2
29 11 11 13 2 16 0 1 9 3 13 9 1 10 9 2 7 15 13 13 1 0 0 2 0 7 0 0 9 2
9 9 15 13 9 2 0 1 9 2
11 3 9 9 13 3 2 16 15 3 13 2
16 9 9 3 3 4 1 9 1 0 9 13 1 9 3 3 2
23 11 2 16 13 1 9 0 9 8 2 13 7 0 3 13 14 1 9 3 3 1 11 2
29 16 1 9 10 9 4 13 1 9 0 9 0 9 2 4 15 1 9 3 0 9 3 3 13 1 9 1 9 2
15 1 0 9 0 9 13 10 9 2 16 15 13 1 9 2
13 1 9 9 9 13 3 0 9 1 0 9 9 2
31 3 7 11 7 11 11 14 13 13 16 0 9 1 9 0 9 2 7 0 9 1 0 7 0 9 13 3 9 0 9 2
32 9 0 9 1 11 13 3 13 0 9 9 2 16 15 14 3 13 1 0 9 9 11 7 13 1 0 9 14 1 0 9 2
23 1 15 4 13 9 14 9 0 0 9 2 16 4 1 15 3 13 9 1 9 1 9 2
26 14 9 1 9 1 9 9 9 0 11 7 9 0 9 1 9 9 0 9 9 4 9 1 9 13 2
25 9 9 9 14 4 13 1 11 2 7 13 0 9 9 2 16 15 0 9 1 15 14 4 13 2
14 0 9 1 9 11 0 1 11 13 0 9 0 9 2
11 1 15 7 13 9 14 3 0 16 9 2
8 7 3 4 13 3 0 9 2
14 1 0 0 4 13 0 2 3 1 9 0 7 0 2
8 9 13 1 14 0 0 9 2
18 0 9 1 9 9 1 9 9 4 13 11 11 1 0 11 1 11 2
24 9 1 9 4 7 1 10 9 1 9 13 0 12 9 0 9 2 16 15 4 13 1 11 2
17 13 1 0 9 1 9 9 9 2 16 15 9 14 3 14 13 2
15 0 9 1 0 11 13 3 0 12 9 7 13 0 9 2
9 3 13 1 0 9 12 0 9 2
15 1 9 15 13 9 13 0 0 9 7 0 7 0 9 2
8 13 14 0 9 1 9 12 2
21 13 1 0 0 0 9 1 11 2 16 13 1 9 9 1 9 7 0 9 11 2
12 9 7 9 1 0 9 0 0 9 1 0 11
18 1 9 9 2 16 13 3 14 9 9 2 4 13 1 11 1 9 2
14 3 4 13 1 9 3 2 16 13 0 9 1 11 2
14 3 4 9 11 13 2 16 13 9 11 1 0 9 2
5 3 13 1 9 2
13 1 0 9 1 9 11 4 13 0 9 1 9 2
8 0 9 15 4 15 13 3 2
16 13 13 2 16 4 1 9 9 11 10 9 13 1 0 9 2
6 3 15 13 15 13 2
12 1 9 13 9 2 1 15 15 13 9 9 2
12 3 7 1 15 4 9 11 13 0 0 9 2
18 9 0 9 7 13 2 16 13 9 2 15 13 1 9 11 2 0 2
40 0 11 2 0 0 9 4 1 9 11 1 0 11 3 13 9 9 9 11 1 10 9 2 1 15 4 13 0 9 9 1 0 9 1 11 2 11 7 11 2
20 3 4 13 3 1 0 9 1 0 9 9 9 11 11 7 14 12 9 9 2
14 2 13 15 1 9 2 2 15 4 13 15 1 9 2
7 1 9 4 13 1 9 2
12 3 3 4 13 14 9 2 1 15 4 13 2
26 9 1 9 1 10 9 13 1 0 9 2 1 15 7 4 13 0 2 15 3 15 4 13 1 9 2
25 3 13 7 9 13 0 9 2 7 14 13 3 2 3 9 15 4 1 12 9 13 1 0 9 2
46 9 11 4 13 0 9 1 3 2 16 4 13 1 0 9 2 1 0 9 12 12 12 3 1 9 12 12 9 2 16 15 4 1 9 9 0 9 9 13 2 0 0 9 11 2 2
42 16 4 11 13 2 16 4 1 0 9 1 9 12 12 9 13 13 1 11 2 16 4 13 10 1 11 0 9 2 4 9 13 2 16 15 4 11 15 14 0 13 2
16 13 15 15 1 9 2 1 16 4 15 3 13 1 0 9 2
25 16 13 9 0 9 3 0 2 7 13 1 9 0 9 14 0 2 7 13 0 9 1 0 9 2
14 16 13 2 13 14 1 15 2 16 4 13 10 9 2
7 1 15 15 13 1 9 2
18 2 14 9 9 7 9 1 9 15 13 1 9 9 13 9 0 9 2
11 1 9 14 2 15 15 3 13 1 9 2
10 2 9 0 9 13 9 9 7 9 2
12 3 13 1 9 0 9 7 13 1 9 9 2
11 14 13 0 9 2 16 13 0 0 9 2
6 9 13 0 9 9 2
10 1 9 13 14 1 9 9 7 9 2
26 2 0 0 9 16 13 9 2 9 1 9 2 9 7 0 9 1 12 1 12 9 13 0 9 9 2
17 9 1 9 13 3 0 2 1 15 13 0 9 14 1 0 9 2
8 1 9 9 13 3 3 0 2
21 2 13 0 9 7 9 1 9 3 13 7 13 2 14 16 4 1 15 13 9 2
7 9 13 3 1 10 9 2
6 2 13 3 1 9 2
11 1 9 2 16 0 13 3 2 13 9 2
7 9 13 0 0 1 0 2
63 0 12 9 1 9 9 1 9 7 9 2 16 13 9 9 0 9 1 9 9 11 2 11 2 7 9 9 1 9 11 2 16 9 13 2 4 15 0 9 1 9 12 9 9 13 14 9 0 9 11 1 0 11 2 1 15 4 9 11 2 11 13 2
44 9 4 1 9 13 2 16 4 1 0 9 9 3 1 0 9 13 9 2 16 14 13 1 9 2 1 15 4 13 1 0 9 1 0 0 9 7 1 1 9 0 0 9 2
15 0 9 13 9 13 1 9 9 1 9 9 1 0 9 2
40 9 9 1 0 9 11 13 10 9 9 9 2 1 15 4 13 9 9 7 9 1 0 9 2 9 7 4 13 14 1 15 2 3 13 1 7 1 0 9 2
16 9 9 13 9 1 11 7 11 2 1 11 7 13 1 9 2
48 11 2 1 9 0 0 9 2 0 9 2 9 7 11 11 4 1 9 2 12 9 2 3 1 9 1 0 9 7 3 1 0 0 9 3 13 0 0 9 9 9 9 11 11 1 0 9 2
28 13 15 4 1 9 0 0 9 11 11 2 16 4 1 10 9 14 13 0 0 9 1 9 1 9 11 9 2
11 0 9 13 13 1 9 9 1 9 9 2
31 1 9 10 9 2 16 13 0 1 9 9 2 3 13 0 9 9 9 2 9 8 1 0 9 9 7 0 9 0 9 2
28 14 3 13 1 9 0 9 2 9 2 9 2 9 2 2 16 4 15 13 1 0 9 1 0 7 0 9 2
11 1 9 13 3 9 2 9 7 0 9 2
24 1 9 9 1 9 13 14 13 14 9 2 7 13 0 3 16 0 9 7 15 13 3 3 2
42 9 1 0 7 0 9 4 13 9 9 11 11 7 13 1 9 9 2 16 13 12 9 2 7 10 9 1 0 7 0 9 2 9 11 11 7 4 13 0 9 9 2
28 0 9 4 1 10 9 1 9 13 9 2 9 7 4 13 14 9 1 9 0 9 2 16 13 14 10 9 2
17 13 14 0 9 7 10 9 3 13 1 0 9 2 0 9 2 2
23 0 4 15 13 1 10 9 7 13 1 0 9 2 1 0 9 7 4 13 0 9 9 2
24 9 9 11 11 4 13 2 16 13 1 9 9 11 1 12 9 14 10 16 12 9 7 9 2
5 0 9 13 9 2
7 0 9 13 14 0 9 2
11 3 4 1 0 9 13 15 12 0 9 2
14 3 4 1 0 2 0 7 0 9 13 3 12 9 2
24 7 15 14 13 2 7 11 4 1 9 13 2 16 15 1 9 9 1 11 14 13 0 9 2
39 1 0 9 2 15 9 13 0 1 12 9 2 16 13 14 1 3 0 9 1 12 9 2 15 4 13 9 7 14 4 13 9 1 0 0 9 1 11 2
14 9 4 13 14 1 0 9 2 14 9 4 14 13 2
26 11 1 9 0 9 4 1 0 9 11 13 14 12 9 0 9 0 0 0 9 2 16 13 0 9 2
30 9 9 9 11 11 13 2 16 4 15 0 13 12 0 9 2 0 9 9 9 7 4 12 9 13 3 1 9 11 2
9 7 10 9 13 9 11 9 9 2
29 15 4 13 3 2 16 15 4 11 13 1 9 9 7 4 9 1 0 9 13 14 0 9 2 0 1 0 9 2
30 1 0 9 0 9 4 3 13 1 0 9 2 16 4 1 9 9 9 7 0 9 11 11 13 9 1 9 9 9 2
22 1 9 4 13 15 11 11 2 11 1 9 9 9 7 11 11 2 11 1 9 11 2
5 1 9 15 13 2
12 1 0 9 4 13 0 0 9 1 0 9 2
13 1 15 4 13 0 9 2 3 7 13 1 11 2
5 13 15 1 9 2
14 3 13 0 2 7 15 9 0 0 9 9 3 13 2
19 3 15 13 2 16 15 4 3 9 13 7 16 15 13 10 14 0 9 2
15 3 15 1 0 13 0 0 9 8 11 1 9 12 9 2
19 9 13 0 0 9 2 7 1 10 9 11 4 13 13 3 0 0 9 2
9 0 9 9 13 1 9 12 9 2
20 9 12 4 13 0 9 7 0 9 2 16 13 0 12 9 7 0 12 9 2
8 0 9 13 0 9 1 11 2
9 9 13 12 9 7 9 0 9 2
11 0 9 0 9 13 0 1 9 8 11 2
8 15 13 14 9 7 0 9 2
14 9 13 9 2 9 1 0 9 13 16 0 0 9 2
24 9 2 16 13 1 9 0 9 2 14 13 9 1 9 1 12 9 1 9 9 1 9 9 2
21 1 9 15 4 1 12 9 1 0 9 13 9 9 0 9 1 0 9 7 11 2
29 1 12 9 13 9 0 9 11 1 11 7 0 9 1 9 2 1 12 9 7 4 0 9 13 0 9 11 11 2
24 13 4 9 0 9 1 11 2 11 2 11 7 11 2 9 7 0 0 9 1 11 7 11 2
21 9 13 1 9 16 4 15 15 3 13 2 4 3 13 0 9 1 10 0 9 2
34 15 7 4 1 0 11 1 0 9 13 9 9 2 16 15 4 13 3 1 9 7 4 13 9 1 9 2 16 4 3 13 1 9 2
42 7 4 13 0 9 11 2 16 13 0 9 7 15 13 11 2 13 12 9 9 9 2 16 4 9 3 13 1 2 9 2 2 16 15 3 1 10 0 9 4 13 2
31 13 9 0 9 9 1 0 9 2 16 4 13 1 9 0 2 13 3 10 9 2 12 9 2 1 12 9 1 9 11 2
19 9 9 13 1 12 9 1 9 11 2 16 4 9 13 9 7 13 9 2
10 2 0 9 13 1 9 12 2 12 2
10 13 2 16 10 9 14 4 13 9 2
14 16 13 1 0 9 2 13 1 0 9 1 0 9 2
14 3 15 13 13 2 16 14 13 15 0 9 1 9 2
9 1 15 15 13 10 9 3 0 2
12 14 13 13 1 0 9 7 13 14 10 9 2
15 9 0 9 4 13 14 3 2 16 4 13 1 0 9 2
23 10 0 9 7 13 2 16 0 9 3 13 14 1 15 2 16 15 4 9 1 9 13 2
24 16 4 13 3 0 9 2 4 10 9 14 14 13 2 7 9 9 13 1 9 0 1 9 2
37 15 13 1 9 0 9 1 0 9 1 9 0 9 1 0 9 2 16 4 13 14 0 9 1 9 2 16 15 4 9 14 13 2 7 3 13 2
15 3 15 4 1 9 13 1 9 9 11 1 10 9 11 2
24 11 4 14 1 11 13 0 9 1 9 11 11 2 16 13 14 0 9 2 12 2 0 9 2
21 16 15 9 1 0 9 3 13 1 0 9 2 7 1 9 7 9 9 3 13 2
21 0 9 1 15 13 9 9 2 16 1 9 7 0 9 0 9 13 3 0 9 2
18 16 15 14 3 15 13 2 4 3 13 0 9 1 9 0 9 9 2
16 9 11 8 11 7 4 13 12 2 0 9 7 0 9 11 2
10 11 13 1 9 9 0 14 0 9 2
17 1 9 13 9 9 9 2 16 13 0 9 9 2 1 9 9 2
10 9 9 11 13 1 0 9 12 9 2
15 11 11 4 13 9 11 11 2 0 1 9 14 0 9 2
45 9 13 12 9 9 11 2 12 9 9 2 12 9 9 2 9 9 2 9 2 0 9 2 9 7 0 9 9 12 2 11 2 9 11 12 2 11 11 2 11 11 9 7 11 2
21 11 11 4 13 14 10 9 2 16 13 9 1 9 7 9 1 9 7 0 9 2
42 1 3 0 9 13 3 13 12 9 2 0 1 11 11 7 13 2 16 4 1 9 13 14 9 2 16 15 13 1 12 9 13 10 9 1 9 7 9 0 0 9 2
21 13 14 2 16 1 11 10 9 14 4 13 1 9 7 13 0 1 9 7 9 2
31 1 0 2 0 9 9 7 4 3 13 12 2 3 13 0 14 0 9 1 0 9 7 3 13 3 3 14 0 0 9 2
21 1 9 13 7 3 13 2 16 4 1 11 14 14 13 2 16 13 14 11 11 2
9 0 0 9 13 12 9 7 9 2
16 13 15 2 16 13 0 9 2 16 15 14 13 13 9 0 2
8 13 15 0 9 2 9 2 2
20 10 9 9 1 0 9 2 9 2 7 9 8 13 1 0 9 2 9 2 2
12 16 13 0 9 0 2 15 15 14 4 13 2
8 9 4 14 3 13 10 9 2
13 14 13 1 15 10 9 0 9 7 0 9 11 2
25 9 9 2 16 3 7 3 3 13 0 9 0 9 2 3 13 1 10 9 2 16 4 13 9 2
42 9 0 9 2 9 2 9 1 9 9 7 9 2 9 0 9 7 0 9 2 9 2 1 15 4 13 9 1 10 9 2 13 9 2 16 15 3 13 9 0 9 2
6 7 13 15 14 0 2
5 13 15 14 3 2
8 13 13 3 9 1 9 9 2
45 15 13 3 1 9 3 13 0 9 1 0 9 9 7 0 0 9 2 16 13 9 9 9 2 9 1 0 9 2 9 1 9 9 9 2 9 2 9 9 1 9 9 7 0 2
35 9 1 10 9 2 16 4 14 13 9 9 2 13 2 16 13 9 9 9 0 2 16 15 13 9 2 16 13 1 9 3 9 16 9 2
27 0 9 1 9 1 11 7 0 9 0 9 4 13 1 10 9 0 16 0 0 9 1 9 9 0 9 2
33 0 0 9 4 7 9 9 0 9 0 9 9 13 7 1 9 10 9 13 2 16 11 13 9 2 16 13 0 1 9 0 9 2
24 0 9 1 0 9 9 1 11 11 13 3 2 16 13 9 2 16 15 9 7 9 4 13 2
28 13 1 0 9 2 16 14 14 13 10 0 9 7 0 9 0 9 2 7 1 15 13 0 9 1 0 9 2
26 0 9 15 13 3 1 9 0 9 7 13 10 3 0 9 2 16 3 9 1 9 13 1 0 9 2
33 13 14 1 0 9 7 9 0 9 2 10 0 9 2 16 13 0 9 7 9 1 0 9 2 7 13 0 9 1 9 1 9 2
10 9 0 9 1 9 4 13 14 0 9
38 1 9 13 13 0 9 1 12 9 2 16 4 1 0 0 9 9 2 16 15 4 13 1 9 11 11 2 1 9 13 1 10 9 3 10 0 9 2
24 9 11 11 4 3 9 13 1 11 7 3 13 2 16 13 0 1 9 7 14 1 9 9 2
36 2 11 11 4 3 13 0 9 2 13 9 2 16 15 4 13 0 11 11 2 16 4 1 0 9 1 0 9 13 9 9 1 9 9 9 2
16 16 15 4 11 13 0 9 1 9 9 2 4 14 15 13 2
17 1 9 11 4 13 9 1 9 9 2 3 7 4 13 9 9 2
9 14 1 9 4 13 9 7 9 2
6 9 4 13 1 9 2
14 15 4 13 1 9 10 9 2 16 4 15 13 9 2
14 9 2 16 15 13 4 15 2 14 13 1 9 3 2
18 1 11 7 13 0 14 9 0 7 0 9 1 9 7 9 0 9 2
24 1 0 9 9 11 11 11 2 16 4 9 13 1 9 7 9 2 4 3 1 10 9 13 2
44 1 0 9 4 13 1 0 0 9 1 0 0 9 2 1 9 7 0 9 1 0 11 1 9 0 0 9 2 1 0 0 9 2 0 9 1 9 7 0 9 1 9 11 2
25 0 9 4 13 0 0 0 9 1 11 2 3 7 13 13 9 1 0 2 0 9 1 9 11 2
11 9 11 11 15 4 13 1 0 9 1 9
11 3 13 9 9 1 0 9 3 0 9 2
13 0 9 9 7 14 9 13 3 0 9 0 9 2
16 3 4 7 13 0 9 7 13 10 9 7 3 13 9 9 2
16 9 1 9 13 14 1 9 2 15 7 4 13 14 0 9 2
22 1 9 4 13 0 0 9 2 16 4 13 0 1 0 9 0 9 0 0 9 9 2
15 11 13 2 16 13 3 0 9 2 16 4 13 1 9 2
20 1 9 9 7 9 3 13 9 1 9 2 15 3 3 13 1 9 1 9 2
25 1 9 12 9 10 9 1 10 9 15 15 13 9 2 9 7 9 2 16 13 0 1 0 9 2
20 1 10 9 9 13 3 13 1 0 9 1 9 9 1 9 7 9 7 9 2
12 0 9 13 1 9 2 16 15 14 3 13 2
32 3 9 3 1 9 13 1 0 9 2 16 15 14 14 13 13 1 9 2 1 15 13 2 0 0 9 2 2 0 9 11 2
24 16 13 13 2 13 9 1 11 11 11 2 16 13 0 9 7 14 0 11 10 9 1 9 2
11 1 9 13 0 12 2 12 0 0 9 2
34 3 1 9 13 9 2 1 9 7 9 2 2 16 13 10 10 9 7 9 1 9 1 11 2 16 15 3 13 1 9 10 0 9 2
21 15 13 0 14 15 2 16 15 14 13 1 9 2 10 9 7 13 15 3 0 2
8 1 9 4 13 14 1 9 2
20 1 15 4 3 13 11 2 16 13 0 9 2 1 15 4 3 13 0 9 2
22 3 3 15 3 13 1 0 9 7 0 9 2 16 13 9 7 15 3 13 1 9 2
25 10 9 2 16 4 3 13 3 0 9 2 13 2 16 1 9 0 9 9 13 3 0 7 0 2
11 9 15 3 14 13 13 1 9 10 9 2
32 9 2 16 13 0 2 15 15 13 0 2 0 2 0 2 13 7 2 10 4 15 15 0 9 13 2 16 4 13 0 0 2
31 1 9 2 16 15 14 13 13 2 1 15 14 13 13 9 7 9 2 1 15 15 13 0 9 2 15 10 9 13 0 2
4 7 14 13 2
17 2 15 13 3 13 2 16 4 13 9 7 3 13 9 1 15 2
26 1 9 13 0 10 0 9 2 16 4 13 1 9 9 0 9 2 8 1 12 9 7 12 9 12 2
31 1 0 9 4 0 9 12 9 13 0 9 1 11 7 9 0 9 1 11 12 2 9 9 13 9 2 7 12 9 11 2
11 9 9 13 0 7 15 15 13 0 13 2
8 9 4 1 9 13 1 9 2
14 9 13 0 7 15 13 0 13 1 9 7 0 9 2
10 9 9 13 9 1 9 1 0 9 2
14 1 0 9 0 13 2 16 13 0 1 9 0 9 2
33 1 9 14 13 13 9 2 16 13 1 9 2 9 7 9 0 9 2 7 0 1 9 11 2 8 8 8 2 7 10 0 9 2
14 13 4 2 16 4 15 13 13 1 9 0 0 9 2
6 1 3 4 13 9 2
11 2 13 4 0 2 9 4 3 13 0 2
11 9 1 9 1 9 1 9 15 13 3 2
3 2 11 2
16 1 0 12 9 15 13 1 0 9 9 9 7 9 0 9 2
48 1 0 9 7 1 0 16 1 0 0 9 2 16 1 0 7 0 9 13 0 9 1 0 9 9 0 9 2 3 13 9 15 2 16 13 2 16 3 9 13 1 9 0 2 3 0 9 2
31 1 0 9 13 14 0 2 7 10 0 9 13 2 16 13 0 0 9 9 13 3 2 16 13 9 0 9 0 0 9 2
14 11 13 9 0 9 0 0 9 7 0 9 7 9 2
17 1 0 9 13 0 9 2 0 13 3 1 9 2 16 15 13 2
10 1 15 7 4 13 1 9 0 9 2
10 0 9 13 14 9 9 1 0 9 2
26 9 9 2 0 9 7 0 9 1 9 7 9 1 0 9 4 1 0 0 9 13 0 9 0 9 2
19 15 7 13 14 9 2 16 15 9 14 3 13 1 9 1 9 1 9 2
13 7 0 9 0 9 1 11 13 1 0 9 9 2
28 1 0 9 9 1 0 11 9 1 11 15 4 10 0 0 9 16 0 3 1 10 9 13 1 0 0 9 2
26 9 13 3 1 9 16 9 2 7 13 1 15 9 10 9 2 1 10 0 9 7 1 10 9 9 2
11 12 1 0 9 13 9 9 1 0 9 2
32 3 1 9 12 9 0 13 2 16 13 9 1 10 9 9 2 7 12 9 2 16 14 13 13 1 15 2 3 3 4 13 2
4 9 0 9 2
11 9 11 11 1 0 9 11 11 1 11 2
14 0 9 2 9 2 9 2 9 4 13 13 10 9 2
20 12 3 0 9 1 15 4 1 9 9 13 0 9 11 11 1 9 9 9 2
18 13 4 2 16 0 9 13 14 0 7 16 15 3 13 14 0 9 2
25 16 4 1 9 13 3 12 9 9 0 1 12 9 2 4 13 13 2 16 4 13 0 0 9 2
32 1 0 9 1 0 9 2 16 4 15 15 0 9 3 13 1 9 7 9 0 9 2 4 13 1 10 9 0 14 0 9 2
18 9 15 4 13 16 9 1 0 9 2 7 4 13 0 9 0 0 2
10 9 4 3 9 12 13 10 0 9 2
23 1 0 9 4 13 9 1 9 1 0 3 7 3 0 9 1 3 0 2 0 9 2 2
18 0 9 4 13 9 2 16 4 15 9 3 1 9 0 9 3 13 2
20 0 9 1 9 11 4 13 1 11 9 12 7 3 3 13 0 9 1 11 2
30 0 0 9 4 1 9 13 1 0 9 1 11 7 11 2 3 7 4 15 13 1 9 2 16 4 15 13 0 13 2
8 3 15 15 4 13 1 11 2
11 14 1 0 9 15 4 13 9 0 9 2
22 1 0 9 4 13 0 9 1 9 2 1 0 9 7 4 9 13 9 1 0 9 2
14 1 0 9 14 0 11 4 13 0 9 7 0 9 2
25 3 0 0 9 4 13 1 9 0 9 2 16 4 13 9 1 9 1 0 9 0 13 0 9 2
24 1 9 0 9 4 13 0 9 1 0 9 2 1 0 9 7 4 0 9 13 14 0 9 2
8 3 4 11 3 13 16 13 2
13 13 15 1 0 9 2 11 7 0 9 0 9 2
28 1 9 1 11 4 13 11 0 2 16 15 4 3 13 1 0 0 0 2 0 2 0 2 0 7 0 9 2
17 0 0 9 13 9 9 2 16 9 0 11 4 13 3 7 3 2
16 11 15 4 13 13 1 0 9 1 3 0 9 16 0 9 2
13 9 7 13 9 9 1 11 7 9 9 0 11 2
17 1 9 11 13 9 9 2 1 0 4 13 9 12 0 11 11 2
15 0 9 13 12 2 0 0 9 2 16 13 9 9 11 2
44 8 11 4 13 9 1 9 9 2 16 13 1 3 0 9 9 0 9 2 16 15 13 0 1 9 13 14 1 9 1 11 2 16 13 15 3 0 1 9 1 0 0 9 2
10 14 7 14 13 10 9 1 10 9 2
11 3 4 13 3 16 0 9 1 11 11 2
21 3 15 4 13 1 0 9 2 1 9 9 2 1 9 2 13 4 10 0 9 2
26 1 10 9 15 4 13 7 4 13 2 16 13 0 0 0 9 7 0 9 2 9 7 13 13 3 2
29 13 4 2 16 13 9 2 16 4 15 13 3 14 0 0 9 7 4 1 0 9 13 14 1 0 9 0 9 2
17 15 4 15 13 7 15 0 9 1 11 13 1 9 0 0 9 2
17 0 11 15 4 3 3 13 1 0 9 10 9 7 13 10 9 2
17 14 10 9 3 4 13 10 9 1 0 11 11 1 0 0 9 2
11 1 9 9 4 15 13 9 1 10 9 2
20 16 9 9 15 14 13 13 2 13 15 3 9 2 16 13 0 1 0 9 2
28 7 15 15 13 14 1 9 9 9 2 16 4 13 1 0 9 3 0 2 9 7 15 3 13 14 1 0 2
19 14 10 0 9 7 9 9 13 9 2 16 15 9 9 9 3 3 13 2
19 0 13 1 9 14 3 9 12 2 16 13 1 9 14 9 1 12 9 2
43 3 12 15 1 0 9 14 13 0 0 7 0 9 2 14 3 7 13 0 11 1 9 1 11 11 16 0 0 9 2 11 11 16 0 0 9 7 11 11 16 10 9 2
16 11 2 0 9 9 0 9 11 13 1 9 14 14 12 9 2
23 0 4 7 1 0 9 13 0 9 2 1 15 4 13 9 12 0 9 7 9 0 9 2
16 9 3 14 4 13 0 9 1 9 3 10 16 12 9 9 2
3 2 8 2
9 7 3 13 11 0 1 10 9 2
20 0 9 4 13 2 16 10 0 9 15 3 13 2 13 7 10 9 0 13 2
11 14 1 9 7 9 9 13 1 0 9 2
23 9 1 9 9 7 13 14 1 15 1 9 2 16 0 9 1 0 9 13 14 0 9 2
18 9 4 14 13 0 7 0 9 9 9 2 0 13 0 12 9 2 2
23 9 9 15 4 1 0 9 13 1 12 9 2 9 7 4 13 1 10 9 12 2 0 2
33 3 4 15 13 1 9 12 1 12 9 1 9 11 1 9 2 16 13 0 3 12 12 9 2 7 1 12 0 7 12 0 9 2
23 0 12 12 9 9 4 14 3 3 13 0 11 2 16 15 4 13 1 10 9 1 11 2
47 0 9 1 9 0 9 0 0 9 7 9 1 9 2 9 9 2 2 16 4 15 1 12 9 9 13 1 9 2 13 14 9 9 2 1 15 13 14 11 11 2 11 11 7 11 11 2
20 2 1 9 1 3 12 3 15 4 1 0 9 1 11 13 12 2 0 9 2
4 15 13 11 2
30 9 4 13 0 7 4 13 3 13 2 7 16 4 9 13 7 13 2 3 7 14 0 13 9 7 3 1 9 13 2
18 15 4 13 3 0 2 0 9 7 4 3 0 13 1 0 0 9 2
25 9 14 13 2 16 0 9 9 2 16 15 13 1 11 2 3 13 16 9 1 9 7 1 9 2
46 3 10 0 9 4 15 1 9 1 11 13 11 7 1 0 9 1 0 9 9 13 3 14 9 1 0 9 2 1 15 14 4 13 0 1 11 12 2 11 11 11 7 11 11 11 2
12 0 9 13 1 9 7 13 0 7 0 9 2
21 16 13 2 3 13 10 9 9 2 1 9 12 13 2 15 13 0 13 1 9 2
21 16 13 9 0 14 1 9 9 11 2 15 4 10 9 1 0 9 9 3 13 2
20 0 9 1 10 9 15 3 3 13 1 0 9 7 9 0 9 1 9 11 2
28 11 2 1 0 9 1 11 1 11 4 13 9 2 9 12 9 9 1 9 2 11 11 7 11 11 0 9 2
11 13 4 9 11 2 11 2 11 7 11 2
15 0 0 9 11 15 4 1 12 9 3 13 1 0 9 2
24 15 4 13 0 9 10 9 9 1 9 2 13 7 4 14 2 3 0 9 13 1 0 9 2
25 16 13 10 0 9 0 9 2 16 13 14 3 3 0 0 0 9 1 11 2 4 3 3 13 2
25 12 9 0 9 2 16 13 1 10 9 2 4 1 0 13 10 9 2 16 4 14 13 0 9 2
19 1 10 9 15 4 13 3 0 0 9 9 9 1 9 1 0 12 9 2
10 1 9 7 3 4 9 14 13 13 2
16 1 3 3 4 3 0 2 0 9 2 13 13 12 0 9 2
24 9 1 10 9 1 0 9 15 4 3 3 3 13 2 7 4 0 0 9 13 14 9 12 2
6 10 9 13 0 9 2
19 16 4 1 10 9 13 3 9 2 15 0 7 3 0 9 14 13 13 2
4 13 15 14 2
16 9 1 9 11 3 3 13 9 2 3 3 7 15 15 13 2
15 3 1 9 13 14 9 2 16 15 3 13 7 3 13 2
5 11 4 13 0 2
8 15 15 3 9 14 14 13 2
5 9 13 1 9 2
18 13 3 0 9 2 0 9 2 0 9 7 9 2 16 13 0 9 2
4 13 0 9 2
15 1 9 13 0 9 1 9 9 2 9 2 9 7 9 2
10 10 9 14 1 9 13 3 12 9 2
12 13 0 9 7 0 9 2 16 13 0 9 2
10 0 9 13 7 15 13 1 0 9 2
9 3 7 16 9 13 14 0 9 2
7 2 3 1 9 13 9 2
26 1 9 13 0 0 9 1 9 7 9 0 9 1 12 1 12 9 2 16 13 9 1 9 1 9 2
12 9 1 9 13 9 7 9 9 1 10 9 2
9 9 9 9 13 0 1 9 9 2
14 3 13 0 9 0 1 0 9 7 9 1 0 9 2
10 1 0 9 4 13 9 1 0 9 2
13 9 4 13 9 1 9 2 13 7 13 0 9 2
17 1 0 9 4 13 0 9 7 15 13 14 10 0 9 7 9 2
22 0 9 9 9 9 14 13 1 0 9 2 7 15 13 1 9 1 0 9 7 9 2
16 9 0 9 9 13 9 7 9 9 1 0 9 7 0 9 2
25 9 0 9 3 13 1 0 0 9 7 7 15 13 9 3 1 9 3 1 9 9 1 0 9 2
42 1 9 4 0 9 13 7 0 9 4 1 0 9 13 3 2 16 4 13 0 9 1 9 1 9 7 1 15 13 0 7 0 9 9 7 3 7 3 13 0 9 2
17 14 4 13 14 9 9 7 15 13 14 1 0 9 1 9 9 2
14 2 3 13 9 1 9 1 9 7 15 1 15 13 2
4 13 9 9 2
8 13 9 1 9 7 13 9 2
19 1 0 9 4 15 13 1 9 9 7 13 9 1 9 1 9 7 9 2
16 2 13 9 10 0 9 3 7 15 1 15 13 1 9 9 2
22 9 9 0 9 9 7 9 11 13 1 11 0 2 0 9 2 11 7 11 14 13 3
18 0 9 1 9 12 13 12 9 9 2 13 7 15 13 1 12 9 9
22 11 2 12 9 1 0 9 11 15 4 1 9 13 0 9 1 9 11 1 9 11 2
15 1 11 4 13 14 0 1 11 2 11 2 11 7 11 2
25 1 15 4 15 13 0 9 1 9 9 0 9 11 2 11 2 1 9 11 2 12 9 1 11 2
27 2 3 15 4 3 9 9 2 16 4 3 13 1 0 9 1 11 2 13 1 11 2 2 13 0 9 2
41 10 9 14 4 15 1 10 9 14 3 13 3 12 9 2 12 9 9 2 14 7 0 9 9 7 4 13 14 9 1 11 2 16 4 15 3 13 1 0 9 2
25 11 2 0 0 9 0 0 9 15 4 3 13 1 0 9 2 9 7 4 15 13 9 7 9 2
31 14 4 15 3 13 14 1 9 2 7 4 9 3 13 2 15 4 1 9 7 9 9 13 9 2 16 9 13 1 9 2
37 0 9 9 2 16 4 15 3 13 1 0 9 2 4 1 0 9 13 9 1 9 1 0 0 9 2 16 4 15 10 9 3 3 13 1 11 2
29 9 4 13 9 7 13 0 9 2 16 1 9 0 2 0 9 9 12 13 9 2 3 13 9 0 0 9 9 2
9 1 11 4 12 9 13 0 9 2
16 16 4 13 1 0 9 9 2 4 9 3 13 0 9 11 2
34 16 4 10 9 13 10 9 1 9 2 4 1 9 9 9 1 12 9 1 12 9 1 12 9 13 0 9 1 11 1 0 0 9 2
19 3 1 10 9 15 4 13 14 15 2 16 4 1 9 13 3 0 9 2
21 0 9 11 4 7 13 13 12 9 9 2 1 15 4 13 10 9 1 10 9 2
16 9 3 0 9 4 3 13 10 9 2 16 4 13 0 9 2
33 1 15 4 3 13 2 16 13 11 0 0 9 7 0 9 1 0 2 16 13 14 10 9 16 0 11 2 1 15 15 13 9 2
15 0 13 14 1 0 9 2 16 14 4 14 13 9 9 2
32 9 9 1 11 3 13 0 9 2 9 1 0 9 7 0 0 9 7 9 1 9 12 2 0 9 2 1 0 9 2 9 2
18 1 0 9 0 9 9 13 3 3 0 2 7 1 11 13 0 9 2
56 1 9 10 0 9 4 9 13 14 0 0 9 2 16 4 15 13 0 9 2 9 0 9 9 7 15 1 0 9 9 13 1 3 0 2 7 3 3 0 9 0 9 2 16 13 1 9 1 3 9 9 2 9 7 9 2
13 1 0 9 0 9 3 13 0 9 1 9 11 2
15 9 4 13 0 9 7 15 13 2 16 4 13 1 15 2
24 3 4 13 2 16 4 13 10 0 9 2 7 13 4 1 3 0 1 9 1 9 0 9 2
12 13 4 9 0 0 9 7 15 3 13 11 2
14 7 0 9 7 0 9 11 15 4 13 13 0 9 2
28 16 0 9 11 1 9 3 13 1 0 9 9 2 4 13 0 9 1 9 14 9 9 2 0 9 7 9 2
25 1 0 9 0 11 7 11 4 13 9 3 0 7 0 9 13 1 15 3 0 16 9 9 11 2
27 2 1 9 0 9 15 1 9 13 9 1 9 2 1 9 3 13 7 1 9 1 9 7 9 13 9 2
17 13 13 2 16 13 0 9 0 2 7 14 13 13 0 9 9 2
12 15 2 16 15 13 2 7 13 13 9 0 2
12 12 9 9 13 1 0 9 13 1 0 9 2
32 7 9 2 0 1 9 7 1 0 9 9 2 16 15 1 9 0 0 9 13 0 2 13 0 1 9 2 0 1 12 9 2
22 0 9 13 3 13 9 1 9 9 2 16 1 10 9 3 13 1 9 7 9 9 2
22 10 9 13 1 14 3 0 9 1 0 9 9 2 1 15 13 10 9 0 7 0 2
21 9 7 9 14 3 13 0 9 9 2 16 13 0 1 0 9 1 9 7 9 2
25 0 0 9 9 4 1 0 9 7 0 9 13 1 3 0 9 7 3 14 4 13 0 0 9 2
7 3 15 4 7 13 9 2
14 9 9 4 13 0 7 10 9 0 9 4 13 13 2
18 9 15 4 13 1 9 1 0 9 7 15 13 13 1 9 0 9 2
16 3 13 2 16 4 15 13 1 9 1 0 9 0 9 11 2
4 15 4 13 2
11 3 15 15 13 2 16 4 13 3 0 2
16 15 13 14 10 9 2 7 15 13 9 14 3 3 16 3 2
12 14 15 14 3 13 2 7 13 15 3 0 2
14 13 15 4 2 13 2 3 16 13 7 9 4 13 2
10 14 3 15 4 13 1 9 1 9 2
6 15 4 13 9 9 2
6 14 13 4 1 9 2
6 14 9 15 4 13 2
13 10 9 0 11 2 9 1 9 9 2 13 9 2
11 7 10 9 11 1 0 9 13 0 9 2
10 0 9 1 9 12 9 0 9 1 11
8 9 13 0 9 9 0 9 2
35 9 0 9 13 0 7 13 0 1 0 9 9 1 9 9 7 9 9 1 9 13 1 9 9 9 2 16 9 7 9 13 10 0 9 2
15 3 3 15 13 1 15 2 16 13 9 0 9 14 0 2
10 3 0 13 9 7 9 1 10 9 2
23 10 0 9 13 1 9 1 0 9 1 9 0 2 7 15 1 10 9 13 3 1 9 2
21 3 0 0 9 13 3 3 3 0 1 0 7 3 12 9 9 13 1 0 9 2
23 9 0 0 0 9 11 13 12 9 7 9 1 9 0 9 12 9 1 0 9 0 9 2
12 9 4 1 11 11 0 9 13 1 11 11 2
22 7 9 16 9 13 1 9 9 2 7 16 3 13 9 1 12 7 1 0 0 9 2
28 13 3 2 16 13 9 10 0 3 0 9 10 0 9 0 9 2 1 15 3 13 1 9 10 3 0 9 2
8 9 9 13 0 1 0 9 2
12 1 9 13 1 10 9 1 9 12 0 9 2
11 1 0 9 9 14 13 3 13 1 9 2
12 9 13 9 1 9 1 9 12 9 0 9 2
10 0 9 9 15 13 1 0 0 9 2
11 9 13 1 0 9 9 7 15 13 9 2
10 0 9 15 3 13 1 9 7 9 2
11 13 3 2 9 9 13 1 9 1 9 2
9 0 9 13 3 3 1 12 9 2
16 9 13 3 0 7 16 9 3 0 14 1 9 1 9 11 2
14 9 13 0 9 0 9 2 1 9 13 0 0 9 2
11 13 0 7 3 15 1 9 13 1 9 2
6 3 15 13 1 9 2
13 10 0 9 13 9 9 7 9 2 13 14 9 2
11 13 3 0 9 1 0 0 9 7 9 2
20 0 9 13 9 0 9 2 16 15 1 0 9 14 3 13 1 0 0 9 2
14 13 0 3 0 9 0 15 0 9 2 3 13 0 2
37 13 15 3 1 9 7 3 13 15 1 3 0 9 2 16 15 13 3 1 9 2 16 13 9 9 7 9 2 14 7 13 15 1 9 1 9 2
11 0 13 3 10 9 13 1 10 0 9 2
13 1 10 9 13 12 0 9 1 12 3 0 9 2
14 10 9 13 0 9 2 0 9 7 1 9 10 9 2
9 13 15 13 3 3 7 1 9 2
8 9 15 3 13 1 0 9 2
13 9 13 0 0 9 2 1 15 15 13 1 9 2
7 0 9 13 0 12 9 2
8 11 4 14 3 13 9 9 2
28 16 13 9 7 13 13 2 16 15 4 1 0 9 13 9 2 15 14 4 15 13 2 16 4 15 13 3 2
24 11 2 3 15 3 14 4 15 13 2 16 1 3 0 9 1 9 3 14 4 15 14 13 2
28 7 15 4 13 1 9 9 2 15 13 1 9 2 16 4 14 10 9 13 1 0 0 9 2 3 0 9 2
33 13 7 3 13 2 16 11 3 13 0 9 2 15 3 13 7 1 9 0 0 9 13 1 0 9 1 9 9 2 9 7 9 2
26 10 9 14 14 13 3 1 9 2 16 4 13 13 14 9 11 2 15 13 15 0 16 0 9 9 2
30 9 9 0 9 2 16 15 4 9 13 13 1 9 9 1 0 9 0 9 2 7 4 13 0 0 9 1 0 9 2
3 2 8 2
18 1 12 9 15 13 9 9 11 11 14 3 3 13 1 10 0 9 2
28 0 9 11 11 13 10 9 2 0 1 9 2 8 8 2 7 9 2 8 8 2 13 3 0 9 1 9 2
13 3 4 13 0 9 2 9 7 13 1 0 9 2
18 1 15 11 3 13 9 1 9 7 9 1 9 9 2 0 11 11 2
12 1 11 4 14 1 9 9 9 13 10 0 9
18 0 9 13 13 0 2 0 1 9 7 14 3 4 3 13 0 9 2
11 0 9 13 0 2 1 9 13 0 9 2
21 15 2 15 4 3 13 2 4 13 3 3 0 1 15 2 15 4 13 1 0 2
20 1 9 1 0 9 7 9 4 7 13 9 1 0 9 2 13 4 10 9 2
27 0 9 15 4 13 0 9 9 2 10 9 7 15 7 4 13 15 15 13 7 1 0 9 13 1 9 2
28 1 0 9 7 3 13 2 16 13 9 0 9 3 7 16 13 3 3 0 2 7 15 4 15 13 10 9 2
20 13 3 0 2 16 4 1 15 13 10 9 2 16 15 14 1 15 14 13 2
20 15 13 2 16 13 9 9 1 10 9 0 7 16 4 15 13 1 10 9 2
13 3 7 9 13 0 9 2 16 15 3 3 13 2
25 13 15 7 15 13 1 0 9 2 7 13 9 1 9 2 1 15 13 9 1 0 9 1 9 2
14 9 7 0 9 2 16 13 1 9 2 13 3 3 2
21 3 15 9 13 2 7 3 13 13 0 9 2 16 7 3 13 1 10 0 9 2
13 3 2 16 15 9 13 2 9 1 15 3 13 2
27 3 15 13 3 13 1 14 0 2 7 0 9 1 9 7 0 13 2 16 15 10 0 9 13 0 9 2
22 9 2 16 13 1 9 2 14 13 2 14 4 15 15 7 14 15 0 13 14 3 2
20 9 2 16 1 9 9 13 1 0 9 2 7 15 3 14 13 1 0 9 2
25 15 15 0 0 9 13 1 9 2 9 12 4 13 1 11 0 12 9 9 1 0 7 0 9 2
18 0 9 4 3 13 12 9 9 9 2 12 9 3 16 1 12 9 2
19 3 13 1 9 1 9 2 9 12 4 9 13 1 9 3 16 9 12 2
17 2 1 9 3 13 15 2 15 3 3 14 13 1 10 0 9 2
14 1 9 13 15 2 15 13 2 0 9 9 1 9 2
8 1 9 15 13 3 3 0 2
32 9 2 16 13 0 9 1 9 2 14 9 0 9 4 13 3 10 9 1 9 10 0 9 2 2 15 1 15 3 13 3 2
18 16 13 3 14 1 15 2 4 9 13 2 16 15 4 13 1 9 2
14 13 4 7 10 9 7 15 1 10 9 14 14 13 2
15 16 13 3 0 1 15 7 10 9 2 13 3 9 0 2
16 4 14 14 13 1 9 2 3 16 13 10 9 3 3 0 2
29 9 7 3 3 0 1 9 13 2 16 14 14 13 9 1 9 1 9 2 9 2 16 15 0 3 2 13 2 2
14 3 4 14 15 0 13 2 16 13 0 9 0 9 2
22 9 13 2 16 15 3 13 0 9 14 1 0 10 9 1 9 2 7 13 3 3 2
18 9 13 2 13 15 15 2 16 14 13 9 7 16 13 0 1 9 2
15 14 15 13 2 16 15 15 4 1 0 9 9 15 13 2
15 16 15 3 13 1 10 9 2 15 13 3 13 1 15 2
32 0 1 15 3 13 3 9 10 9 7 16 15 15 4 1 10 9 14 13 2 4 3 13 12 1 0 7 0 9 1 9 2
26 0 13 2 16 9 13 9 2 14 3 7 13 14 9 0 9 2 7 1 9 16 1 0 0 9 2
6 15 7 3 3 13 2
28 13 2 16 4 13 7 13 9 2 7 16 13 10 9 0 1 9 10 9 2 15 13 2 16 13 9 15 2
22 7 7 3 13 9 2 3 15 3 13 2 16 15 4 1 10 9 13 3 14 15 2
9 9 3 13 2 3 3 13 9 2
34 10 9 4 13 14 1 0 0 9 2 3 7 4 3 1 9 13 7 15 1 10 9 13 1 15 2 13 2 1 0 9 7 9 2
21 9 9 13 12 0 0 9 7 10 9 13 0 2 16 15 15 4 13 1 15 2
22 14 2 16 13 9 14 0 7 2 14 13 2 2 15 14 3 13 10 2 9 2 2
24 1 0 0 9 7 0 0 9 15 13 1 10 9 2 16 4 13 2 10 13 10 9 9 2
10 3 15 14 13 13 1 9 7 9 2
29 13 9 2 16 15 4 15 13 12 1 10 9 2 1 0 7 13 0 13 9 1 0 0 9 2 16 13 3 2
31 15 7 13 3 3 0 7 1 9 16 1 10 9 2 7 9 1 0 9 13 2 3 10 9 1 15 13 13 0 9 2
39 16 7 13 0 9 3 2 15 9 14 3 13 1 15 2 16 13 2 0 2 2 9 7 13 10 9 9 2 16 15 10 9 1 0 13 1 10 9 2
26 16 13 14 0 0 0 9 2 13 1 10 10 2 9 2 1 0 9 7 13 4 13 9 1 9 2
18 10 9 15 13 1 9 7 15 4 15 3 3 3 13 1 9 15 2
11 7 15 14 3 13 9 1 9 1 9 2
22 16 13 9 3 0 9 2 13 3 9 1 10 9 0 9 7 14 9 9 1 9 2
19 3 4 13 2 16 4 14 15 13 10 0 9 2 16 15 13 2 14 2
13 1 9 4 1 3 1 0 13 14 10 0 9 2
24 13 4 9 2 13 0 9 1 9 9 7 14 1 0 9 0 9 7 13 9 1 0 9 2
27 1 10 9 14 4 9 11 9 13 14 9 0 7 0 9 7 13 9 1 9 1 0 9 7 1 11 2
8 0 13 14 1 9 7 9 2
11 2 15 15 13 2 16 1 9 13 9 2
18 9 1 0 7 0 9 13 1 9 15 2 1 9 1 10 0 9 2
34 11 11 11 13 2 16 4 13 0 9 13 9 1 10 9 2 16 13 0 9 0 0 9 2 7 9 2 0 9 2 1 9 9 2
16 9 0 9 1 9 9 4 1 11 13 10 16 12 0 9 2
8 0 9 4 13 9 9 9 2
3 2 8 2
18 14 13 9 10 9 9 2 16 4 15 14 1 0 9 14 3 13 2
40 3 4 15 13 14 1 0 9 9 7 9 9 7 9 9 2 16 4 2 16 4 3 13 2 10 9 3 14 13 9 9 1 0 0 9 1 11 0 9 2
35 16 0 9 1 0 2 0 9 13 1 9 14 0 3 0 9 10 9 2 15 13 13 2 16 4 13 1 9 10 9 7 9 0 9 2
19 1 0 9 13 0 9 2 16 14 3 13 10 9 2 0 14 10 9 2
33 3 0 4 13 9 1 10 0 9 0 9 1 15 2 16 4 15 13 1 9 0 7 15 3 13 14 1 9 0 9 1 11 2
10 3 3 1 11 4 13 9 0 9 2
27 10 0 9 4 13 13 14 0 9 2 4 7 13 3 3 2 16 10 0 9 1 0 9 3 14 13 2
7 1 9 9 4 13 0 2
9 14 0 9 4 3 13 9 9 2
24 3 13 7 7 9 1 9 0 9 7 0 9 1 9 9 7 14 9 9 1 9 0 9 2
11 10 9 15 1 9 13 14 0 9 9 2
19 9 2 16 13 1 15 2 3 3 4 0 9 13 9 2 14 13 9 2
28 3 16 15 1 10 9 10 9 13 0 9 2 7 7 13 13 2 16 1 9 14 13 3 13 1 0 9 2
10 14 3 0 4 13 9 13 0 9 2
10 14 3 4 13 10 9 9 0 9 2
11 14 7 4 9 13 10 9 9 10 9 2
19 3 13 14 0 9 10 9 2 16 4 15 1 0 9 13 1 10 9 2
15 1 15 7 4 13 9 0 9 7 9 1 9 3 0 2
20 1 15 4 13 0 9 2 7 15 4 13 1 0 9 14 3 0 0 9 2
11 9 9 4 9 13 14 1 10 0 9 2
8 14 11 7 11 4 13 3 2
6 11 4 3 13 9 2
5 13 4 3 0 2
6 11 4 13 10 9 2
5 13 15 1 15 2
6 16 13 11 0 15 2
19 1 9 2 16 15 4 13 1 9 2 15 4 13 13 1 9 9 9 2
14 2 14 2 13 13 3 0 2 14 3 7 3 13 2
12 16 15 15 13 0 13 2 15 15 14 13 2
9 13 4 2 10 9 3 13 9 2
31 9 2 0 9 13 1 0 3 0 2 8 13 10 9 2 16 7 15 4 15 3 3 13 2 4 13 2 16 14 13 2
12 2 14 13 2 16 13 0 13 10 9 3 2
8 14 15 13 2 4 13 11 2
6 3 15 4 13 11 2
8 2 13 2 14 13 3 3 2
14 15 9 13 9 1 10 0 9 2 6 2 7 13 2
21 11 15 13 2 16 1 9 13 11 7 13 2 10 9 15 13 3 13 1 9 2
8 2 7 14 9 13 10 9 2
10 9 4 13 11 1 9 7 1 9 2
8 11 15 4 15 0 3 13 2
31 4 14 15 13 2 3 4 10 9 3 9 13 3 16 15 2 15 4 13 14 3 0 2 16 4 1 15 0 9 13 2
8 15 15 3 10 9 14 13 2
16 9 7 9 8 14 3 3 13 2 15 13 1 10 9 13 2
7 12 0 0 9 15 13 2
40 0 0 9 2 0 9 7 0 9 15 3 13 7 13 3 13 10 9 7 15 13 2 7 13 15 3 1 9 2 0 7 7 15 3 13 9 1 15 3 2
18 3 15 13 1 11 7 15 3 3 13 2 10 9 9 0 16 13 2
31 9 14 13 2 8 13 13 9 1 9 2 14 15 4 13 3 2 16 8 13 11 7 7 11 2 16 3 13 11 11 2
14 13 2 16 4 15 3 13 2 16 4 13 14 0 2
12 13 2 9 15 4 3 3 13 1 10 9 2
16 1 15 4 15 7 10 0 9 2 11 2 10 0 9 13 2
14 8 11 2 4 15 1 10 9 14 3 1 15 13 2
6 10 0 9 7 9 2
13 13 15 10 9 2 3 4 13 7 3 9 13 2
11 1 3 3 2 9 2 4 13 1 15 2
9 8 13 2 16 15 13 1 9 2
7 9 4 15 13 1 9 2
3 9 13 2
3 13 15 2
6 3 7 15 13 3 2
12 14 9 7 3 13 0 2 0 2 0 9 2
36 3 15 13 2 16 14 13 1 9 7 15 13 9 1 9 3 1 9 2 14 15 15 13 2 16 16 8 15 0 13 2 16 15 13 13 2
12 1 15 15 14 0 9 1 9 13 16 9 2
10 10 9 15 13 2 16 13 1 9 2
9 16 15 13 2 15 13 1 9 2
5 3 13 14 0 2
10 3 15 13 2 1 10 9 13 9 2
14 0 13 2 16 4 13 10 9 2 4 3 13 11 2
38 16 14 13 10 9 1 0 10 9 2 3 3 14 13 2 16 15 9 0 3 13 7 15 1 11 13 2 16 15 15 1 9 13 2 4 15 13 2
17 3 15 13 9 2 14 4 13 3 3 0 2 15 15 9 13 2
18 4 13 12 10 9 2 8 4 1 15 13 2 7 4 13 1 9 2
10 11 13 1 9 7 1 15 13 9 2
7 1 9 0 9 13 9 2
16 14 13 15 9 2 14 9 9 1 0 9 4 15 3 13 2
13 7 3 4 1 10 9 1 9 14 13 12 9 2
17 0 9 13 0 9 9 2 16 15 13 1 9 1 9 0 9 2
8 3 0 13 1 9 1 9 2
7 15 13 2 16 13 0 2
13 11 11 3 13 10 9 2 16 13 3 0 9 2
8 16 4 15 3 13 15 15 2
15 14 1 9 13 7 13 9 7 15 13 13 2 7 13 2
6 1 9 4 15 13 2
19 11 15 4 13 1 11 2 10 9 2 7 15 4 13 2 16 13 3 2
25 16 4 15 13 2 4 11 14 3 13 1 9 1 11 7 14 15 9 7 15 13 12 1 0 2
10 11 4 13 10 9 1 10 0 9 2
15 13 4 2 3 4 15 13 1 9 2 3 7 3 13 2
8 3 4 13 15 9 7 9 2
14 3 4 13 0 9 7 13 9 3 2 16 4 13 2
13 10 9 7 9 4 13 2 7 15 15 4 13 2
19 13 4 2 16 4 15 15 13 2 7 4 13 9 10 9 14 15 0 2
9 15 13 1 12 9 2 1 9 2
5 11 13 13 3 2
7 2 15 13 3 0 9 2
6 13 8 2 13 9 2
4 15 13 0 2
11 2 14 2 15 13 12 0 9 1 11 2
5 14 13 15 13 2
11 9 2 7 4 15 13 2 16 13 0 2
8 15 13 3 3 0 2 13 2
9 9 3 3 13 13 0 0 9 2
13 2 0 9 8 3 13 9 1 9 2 15 13 2
19 13 1 9 1 9 2 16 13 11 2 16 13 3 1 11 2 10 9 2
11 11 4 9 13 16 0 1 12 0 9 2
11 1 9 9 13 3 13 12 9 0 9 2
21 9 13 1 0 9 2 7 13 9 7 9 3 1 0 9 1 10 9 1 9 2
12 9 13 2 16 4 9 14 13 9 12 9 2
23 0 9 9 2 16 4 15 13 1 9 2 4 15 13 14 0 9 10 0 9 1 11 2
13 0 9 7 13 7 14 9 1 9 1 10 9 2
19 16 0 0 9 3 0 1 15 13 14 3 0 1 10 9 1 0 9 2
19 1 15 14 14 13 13 2 16 13 14 1 9 7 9 9 1 0 9 2
32 0 9 10 9 13 0 9 1 9 10 9 1 9 1 11 2 1 15 13 9 1 9 7 9 9 2 0 1 9 1 9 2
24 3 1 9 4 1 0 9 13 9 11 11 1 9 2 2 16 4 13 15 2 15 4 13 2
41 16 4 15 1 9 9 2 3 14 15 13 1 9 2 13 14 10 9 2 15 4 13 0 2 16 4 13 0 2 16 4 3 13 3 2 16 4 13 1 9 2
17 15 13 15 2 15 3 13 2 3 1 15 2 16 13 9 0 2
13 9 15 4 14 13 2 16 4 13 0 9 0 2
26 13 15 0 9 0 0 9 2 0 9 0 9 7 9 2 0 0 0 9 4 3 13 1 10 0 9
7 11 11 13 1 9 9 2
27 0 9 15 14 13 3 3 2 3 15 13 0 9 2 16 13 9 0 9 2 0 9 7 9 1 11 2
23 16 9 9 2 16 13 9 11 2 15 14 13 9 11 2 3 16 4 9 13 11 11 2
27 0 0 9 2 11 2 4 13 2 16 13 9 1 9 0 0 9 12 0 12 9 1 12 9 1 11 2
12 1 9 0 9 15 4 13 9 11 11 11 2
37 0 9 7 9 13 0 7 14 0 9 2 13 12 1 9 2 16 15 4 13 9 9 9 9 0 9 1 9 9 0 9 7 9 1 0 9 2
22 16 9 9 3 13 0 9 11 2 1 15 4 13 14 9 11 11 11 7 11 11 2
17 0 9 2 1 15 4 15 9 13 2 13 1 9 10 0 9 2
17 3 13 9 7 10 10 9 3 0 1 9 9 2 8 8 2 2
9 15 13 1 0 9 7 9 0 2
18 1 9 13 9 9 2 16 13 7 13 9 2 9 7 13 9 0 2
26 1 9 9 3 9 13 0 9 1 9 0 9 7 9 9 2 16 7 13 1 9 10 9 0 9 2
24 1 9 0 9 15 13 7 13 9 2 9 2 9 7 9 0 9 2 16 15 13 0 9 2
22 10 9 4 13 0 15 2 0 4 13 0 1 9 7 7 4 13 0 12 1 0 2
21 0 4 13 10 0 9 7 0 7 0 9 2 9 7 9 4 13 14 3 0 2
12 13 4 14 12 9 2 7 10 9 3 13 2
8 9 1 10 9 14 14 13 2
8 13 3 9 2 9 14 13 2
21 0 7 3 0 9 13 7 15 13 0 1 9 7 1 15 2 10 4 13 9 2
6 3 13 0 9 9 2
9 13 15 14 0 2 7 13 3 2
20 16 13 12 9 2 15 9 0 9 14 13 14 15 2 16 4 13 0 9 2
21 1 15 13 14 9 2 9 2 16 3 13 7 13 0 9 2 15 1 15 13 2
19 15 13 0 7 3 14 13 14 9 2 16 15 13 13 14 1 12 9 2
20 13 3 1 11 9 9 1 0 9 2 9 1 0 9 7 9 1 0 9 2
6 14 4 3 13 9 2
6 9 4 13 3 0 2
6 9 9 15 3 13 2
12 16 13 1 9 2 13 9 2 16 15 13 2
19 0 9 13 2 16 13 0 9 9 2 7 9 2 1 15 13 3 13 2
16 13 15 3 3 2 7 15 4 3 13 13 1 10 9 3 2
13 13 0 9 9 7 13 15 2 16 13 1 15 2
13 9 1 0 9 9 15 13 2 15 9 9 13 2
33 9 14 13 0 9 3 16 1 9 15 13 1 0 9 7 0 9 9 2 16 15 0 9 14 13 13 1 14 10 10 0 9 2
14 2 10 9 13 0 9 7 9 2 16 15 13 13 2
14 1 11 1 0 9 0 9 1 11 4 13 0 9 2
6 14 1 11 13 0 2
25 11 11 13 2 16 4 1 11 13 1 12 7 12 9 2 16 4 11 3 13 0 7 0 9 2
28 1 9 1 9 9 1 11 15 14 13 13 2 16 13 1 0 9 2 16 13 1 0 9 2 4 13 11 2
21 0 9 11 11 15 4 1 0 9 13 2 16 13 3 13 9 9 16 15 13 2
33 3 4 1 9 9 11 11 11 7 11 11 11 13 3 3 2 16 4 3 3 1 0 9 11 11 7 9 11 11 13 0 9 2
11 7 0 9 11 11 4 9 13 1 9 2
32 11 2 16 13 9 1 0 9 1 11 14 0 9 2 15 9 1 9 0 9 11 11 1 9 4 3 13 1 9 1 9 2
16 0 9 9 9 4 9 14 3 13 1 9 7 9 9 9 2
24 9 9 4 10 0 9 13 14 9 1 0 9 2 16 3 14 1 0 9 1 9 13 9 2
14 0 9 1 11 3 3 13 2 13 7 15 14 0 9
23 9 2 0 4 13 12 12 12 7 4 15 13 12 12 12 2 15 13 1 12 9 9 2
17 13 14 12 9 2 12 9 7 12 9 9 2 0 1 0 9 2
4 13 12 9 2
7 3 4 13 3 1 9 2
32 16 13 3 3 2 13 14 0 2 16 15 3 13 10 9 9 2 16 15 4 13 2 16 4 1 10 9 13 14 10 9 2
22 16 13 3 0 2 15 4 3 3 13 1 9 7 9 9 7 9 0 9 1 15 2
18 13 9 1 9 2 15 15 9 13 7 3 4 13 2 16 13 0 2
5 13 1 9 9 2
29 13 15 3 2 16 9 1 10 9 13 7 16 15 1 0 9 1 10 0 9 13 2 3 13 10 0 9 0 2
24 9 1 11 2 16 4 13 1 9 3 0 4 13 13 1 0 9 2 7 4 9 3 13 2
21 9 14 13 0 9 1 0 9 2 16 15 4 13 11 11 2 0 9 0 9 2
22 0 9 9 4 13 14 3 0 14 1 9 0 9 2 9 11 11 2 0 0 9 2
38 9 9 11 11 7 9 11 11 4 13 9 7 9 11 1 10 0 9 7 0 9 7 15 15 13 1 9 9 2 16 15 4 13 14 1 9 9 2
26 11 11 4 13 2 16 15 4 13 3 0 2 16 4 9 9 13 1 9 2 16 13 1 10 9 2
12 1 9 7 4 13 9 0 11 0 7 0 2
5 2 16 13 0 2
5 1 15 1 9 2
7 7 3 13 9 1 9 2
22 0 11 14 15 4 9 3 13 9 1 9 1 9 7 7 4 13 14 2 9 2 2
16 9 4 1 9 13 0 12 12 12 9 0 9 9 0 9 2
8 3 13 10 0 9 1 9 2
15 3 13 2 16 15 9 1 10 9 14 4 13 7 13 2
9 3 13 0 9 1 10 0 9 2
13 15 13 15 2 15 4 1 10 9 13 10 9 2
21 0 9 9 13 14 9 2 16 1 9 13 13 1 0 2 0 7 3 0 9 2
23 9 2 0 9 2 1 9 12 9 12 1 9 1 11 2 11 7 11 7 1 9 1 11
26 16 15 4 11 8 1 11 1 9 13 1 0 9 11 2 4 13 2 16 4 1 11 13 1 9 2
22 11 4 9 1 0 9 13 1 9 7 9 1 9 2 16 15 4 10 0 9 13 2
3 2 8 2
5 9 13 1 9 2
12 1 0 4 0 9 10 9 13 12 9 9 2
11 1 9 0 9 13 9 0 9 1 0 9
3 2 8 2
12 1 9 9 13 0 1 9 11 13 14 10 9
24 9 13 1 9 2 16 13 0 1 9 2 4 13 9 9 9 1 9 1 0 9 11 11 2
29 0 9 13 1 9 9 0 9 1 9 7 9 2 1 15 7 13 0 9 9 2 9 7 0 9 9 7 9 2
13 10 9 15 13 2 9 15 13 15 2 15 13 2
22 0 9 9 2 16 15 3 13 7 13 1 10 9 2 13 3 1 12 9 0 9 2
8 10 9 15 3 13 1 9 2
12 13 0 2 3 15 13 13 7 13 3 0 2
13 9 13 3 7 15 13 1 15 2 13 11 11 2
17 3 0 13 7 1 15 16 14 1 0 2 1 9 13 3 3 2
4 9 13 3 2
32 11 14 4 16 9 9 11 8 8 8 13 9 9 1 9 1 0 9 2 1 15 7 13 2 16 11 13 9 1 9 9 2
14 9 11 11 4 3 1 11 13 0 9 1 0 9 2
19 1 15 4 15 13 11 11 11 2 0 11 2 7 11 11 2 0 11 2
7 3 4 13 9 3 3 2
13 3 4 13 2 16 13 9 0 0 9 14 3 2
23 15 7 14 13 1 9 14 0 0 9 2 7 14 9 1 0 9 2 0 9 7 9 2
18 9 0 9 13 0 14 0 9 1 9 0 9 9 7 0 9 9 2
8 1 0 9 4 13 12 9 2
24 0 13 0 16 0 9 0 9 0 9 3 1 12 0 9 2 16 4 15 13 0 9 9 2
22 0 9 13 0 1 9 9 1 9 1 0 9 3 1 0 0 9 7 9 10 9 2
38 0 9 7 13 0 1 9 9 2 16 4 1 0 9 13 1 9 1 15 4 13 9 2 16 13 1 9 2 7 9 2 16 4 13 1 15 0 2
20 9 9 4 13 14 9 7 0 9 1 0 9 2 3 7 3 13 0 9 2
8 10 9 9 3 13 1 9 2
14 14 13 10 9 9 2 16 13 3 1 9 3 0 2
14 16 9 15 13 2 3 15 1 9 9 13 13 9 2
22 9 9 13 0 9 2 0 1 10 9 2 16 15 13 13 3 1 3 0 0 9 2
9 10 9 9 13 9 1 9 9 2
11 1 10 9 15 9 13 1 0 9 9 2
14 10 9 9 9 14 13 7 1 9 0 9 13 9 2
31 1 9 7 10 0 9 2 9 2 0 9 13 3 14 0 13 2 15 4 9 13 7 1 15 13 1 9 1 0 9 2
26 1 0 9 13 14 10 0 9 9 9 2 16 13 0 9 1 15 2 3 3 13 9 0 1 9 2
17 0 9 1 10 0 9 3 13 9 1 10 9 7 1 9 9 2
21 16 13 10 9 0 2 15 3 13 1 10 9 7 13 0 9 14 1 10 9 2
9 0 9 3 13 1 9 1 9 2
21 0 9 2 9 13 0 9 2 1 15 13 0 9 1 9 0 1 0 0 9 2
14 3 4 13 13 0 1 9 1 9 2 1 15 13 2
17 3 2 16 13 10 9 2 9 7 9 2 3 13 0 0 9 2
9 9 11 9 0 0 9 13 0 2
12 1 10 9 4 15 13 10 0 9 13 9 2
21 3 4 13 13 9 1 0 7 0 9 7 13 2 10 13 1 9 1 15 9 2
20 13 4 15 14 13 9 7 9 2 16 15 13 7 13 0 9 1 0 9 2
8 9 9 13 0 3 7 3 2
14 16 4 13 9 7 9 9 2 13 14 9 9 9 2
19 9 3 13 12 7 3 9 2 10 9 7 3 13 12 7 3 9 9 2
18 3 13 0 7 15 13 2 3 15 15 13 7 3 4 15 3 13 2
13 13 15 4 9 2 16 13 2 3 13 15 0 2
9 10 9 15 13 9 7 13 9 2
8 9 9 12 13 0 9 9 2
16 9 9 12 13 3 0 7 13 13 0 1 0 9 9 9 2
18 0 9 4 13 9 9 1 12 9 1 9 2 9 9 7 9 9 2
23 1 9 9 2 16 13 2 15 9 13 9 2 3 1 9 13 0 13 0 9 9 9 2
8 9 12 13 9 1 9 9 2
22 1 10 9 15 4 13 1 10 0 9 9 7 0 9 2 16 15 3 13 1 9 2
7 13 15 4 0 0 9 2
30 1 0 9 9 2 7 9 9 9 2 3 13 9 2 16 1 0 9 13 9 1 9 9 7 13 3 0 9 9 2
27 16 4 15 3 1 0 9 13 0 9 2 4 13 3 0 9 2 16 13 3 0 2 16 13 9 9 2
27 13 14 9 9 7 0 0 9 2 16 13 11 2 11 2 9 2 9 2 9 9 2 7 15 0 9 2
13 1 9 13 10 9 3 0 7 13 9 10 9 2
18 0 10 9 15 4 13 10 9 2 16 14 13 0 16 9 1 9 2
13 13 14 0 9 0 9 2 16 13 0 9 9 2
7 9 1 9 13 12 9 2
13 0 13 13 10 9 3 15 13 13 0 9 9 2
26 13 2 16 15 4 0 9 9 14 15 13 2 7 16 10 9 3 13 13 2 13 14 15 0 9 2
11 0 9 13 9 0 9 1 0 9 9 2
19 15 13 3 3 0 1 9 1 9 7 13 14 10 9 1 0 0 9 2
10 15 1 10 9 4 13 1 0 9 2
3 0 9 2
4 4 14 13 2
30 9 9 2 16 13 9 2 9 7 9 3 13 1 10 9 2 7 9 9 12 13 2 16 1 15 3 13 0 9 2
13 9 13 9 9 9 7 3 9 13 0 0 9 2
13 1 9 1 9 15 9 3 13 14 1 9 1 9
26 1 9 2 3 4 15 15 3 13 2 4 3 13 1 10 9 2 16 13 1 0 9 1 9 9 2
17 9 4 0 9 13 1 0 10 12 0 9 2 12 9 13 13 9
13 11 4 7 1 0 9 13 9 10 0 0 9 2
30 13 4 15 14 10 9 1 10 9 1 0 9 0 9 1 11 2 3 7 4 13 11 14 0 1 9 0 9 11 2
17 13 7 15 4 14 1 0 9 2 16 13 1 9 14 3 0 2
7 0 9 15 4 3 13 2
10 14 13 3 0 1 0 9 9 9 2
7 9 13 3 3 16 3 2
17 1 9 7 13 1 9 2 16 15 4 1 0 9 13 1 9 2
13 9 15 13 1 9 9 2 16 4 13 3 0 2
8 3 4 9 13 1 0 9 2
10 9 3 4 15 13 14 14 0 9 2
11 1 9 1 9 4 13 9 1 0 9 2
28 9 15 4 13 1 9 0 9 1 10 0 9 1 0 9 9 2 16 14 4 15 1 9 9 13 9 0 2
11 0 9 9 4 0 9 13 1 0 9 2
23 15 2 16 15 4 13 1 9 2 4 1 9 13 9 9 2 16 4 0 9 3 13 2
17 3 0 4 2 16 4 15 15 13 1 9 2 13 9 7 9 2
10 16 16 4 13 9 1 9 15 0 2
20 1 10 9 15 11 13 1 0 7 0 9 11 1 9 1 9 1 0 9 2
21 10 9 13 0 7 0 2 3 7 13 11 16 12 1 0 9 1 9 1 11 2
12 0 9 3 13 0 2 7 3 13 14 0 2
24 14 9 4 1 11 11 3 13 3 1 9 2 3 7 4 15 9 7 9 13 7 13 9 2
19 0 9 0 9 2 0 9 7 0 9 13 14 3 0 1 0 9 9 2
9 14 2 15 4 7 13 1 15 2
15 1 9 13 3 0 2 15 7 15 3 14 13 10 9 2
12 0 9 14 4 1 0 9 13 14 0 9 2
12 1 9 14 4 15 13 9 10 12 0 9 2
12 1 0 9 9 13 9 1 11 12 0 9 2
7 1 9 7 13 14 9 2
21 14 0 9 4 1 0 9 13 2 16 4 15 13 3 1 9 9 9 3 13 2
33 1 0 9 9 9 9 1 11 12 3 3 14 4 13 2 7 15 4 13 14 16 9 2 16 4 3 0 9 12 3 13 9 2
24 0 9 0 9 4 13 3 3 2 16 4 13 1 11 12 1 9 7 2 13 2 12 9 2
18 0 9 15 9 3 13 1 9 9 9 1 0 9 9 1 0 9 2
15 3 16 10 9 9 11 11 11 11 4 13 14 1 9 2
10 13 4 2 16 15 4 13 13 9 2
18 2 0 9 1 9 2 4 13 3 0 9 1 9 9 1 0 11 2
31 2 16 4 9 12 13 9 2 4 13 1 15 10 9 16 0 9 2 2 15 13 11 2 16 13 9 1 10 0 9 2
14 2 16 4 11 9 3 13 2 4 13 3 3 0 2
3 14 0 2
6 7 4 3 13 9 2
39 0 11 2 8 2 2 15 12 0 2 1 15 15 4 1 0 0 9 1 9 13 9 1 0 9 9 9 2 4 15 13 2 16 15 4 13 1 9 2
35 0 4 13 8 8 1 9 1 0 9 2 16 4 13 9 1 9 2 16 4 1 9 2 1 9 9 2 13 12 0 9 1 12 9 2
14 1 9 1 0 9 11 7 4 15 12 9 13 12 2
11 1 9 11 13 2 16 15 3 3 13 2
36 0 9 3 0 9 0 9 9 11 2 16 4 13 1 9 11 2 15 0 9 3 13 1 9 0 9 2 16 15 3 13 0 9 7 9 2
16 11 13 0 9 1 10 10 9 2 1 9 13 9 0 9 2
23 1 0 9 13 1 9 0 0 9 2 16 13 3 0 7 0 1 0 0 7 0 9 2
17 1 0 9 15 13 0 7 0 0 9 9 2 9 7 0 9 2
12 10 9 13 9 9 7 13 9 1 0 9 2
20 1 9 9 15 13 0 7 0 0 9 2 7 15 14 13 3 3 1 11 2
8 0 9 9 13 0 9 11 2
13 0 9 13 0 0 9 2 3 15 13 7 13 2
20 1 0 11 15 3 1 11 7 0 9 13 0 9 2 0 1 9 0 9 2
14 13 12 0 7 0 0 9 10 0 9 1 0 11 2
15 9 13 0 1 12 9 2 10 9 13 9 1 12 9 2
6 9 13 3 0 9 2
25 1 0 9 13 0 2 16 13 0 2 3 0 9 7 15 1 0 9 1 10 9 13 3 3 2
9 1 0 9 15 13 0 0 9 2
21 9 2 16 15 4 13 2 3 9 13 1 9 0 9 2 0 9 0 0 9 2
11 9 0 9 14 13 0 3 2 14 3 2
12 3 13 9 0 2 3 2 13 1 0 9 2
20 3 14 15 13 1 9 9 2 16 13 1 9 0 9 7 1 9 10 9 2
10 9 14 9 1 0 9 13 10 9 2
10 9 3 13 3 2 1 9 0 9 2
10 0 9 9 7 12 3 0 9 1 9
10 10 9 13 3 14 1 9 1 9 2
21 15 14 3 3 13 9 2 16 4 13 14 1 9 7 15 9 3 13 1 15 2
17 13 10 9 2 16 4 3 13 9 2 16 4 14 14 9 13 2
7 13 10 9 2 4 13 2
3 9 9 2
15 16 13 13 1 9 1 0 9 2 13 13 13 14 9 2
4 9 14 13 2
11 1 15 7 13 14 1 9 0 9 9 2
5 9 11 2 9 2
15 15 13 0 2 3 7 13 9 9 2 16 13 3 12 2
24 15 4 3 13 2 16 4 13 1 9 9 2 16 13 9 2 16 15 4 15 1 9 13 2
3 9 0 2
19 1 9 9 1 10 9 1 0 9 13 0 0 9 9 7 0 0 9 2
14 0 9 0 9 2 0 9 2 0 0 9 2 0 9
11 14 11 4 10 0 0 9 13 9 12 2
37 10 9 2 16 15 4 3 13 7 4 15 13 14 1 12 9 2 4 13 9 12 7 14 3 0 2 1 15 4 13 3 0 9 11 2 11 2
3 0 9 2
11 9 1 0 9 2 0 9 2 12 9 2
16 10 0 9 13 9 9 2 0 9 2 0 9 9 7 0 2
11 7 14 1 9 1 0 9 14 13 13 2
21 1 0 9 0 9 2 16 13 1 10 9 13 9 2 13 1 10 9 0 9 2
16 13 4 7 2 16 4 0 9 3 1 10 9 13 3 3 2
27 16 9 9 1 9 4 13 13 9 1 9 10 9 2 1 15 4 15 3 13 9 1 0 9 13 9 2
31 1 0 9 1 0 11 15 11 13 9 2 16 3 1 11 1 11 13 1 0 9 14 1 9 2 1 15 13 10 9 2
12 0 9 1 9 9 14 14 13 1 9 1 9
10 4 3 11 7 13 10 0 9 9 9
19 1 0 9 15 4 9 13 14 1 0 9 2 0 9 7 15 4 13 2
20 11 15 9 4 13 2 1 0 9 7 0 9 15 4 13 3 13 0 9 2
42 3 13 9 0 2 15 3 7 3 13 9 0 9 9 11 11 2 16 13 1 10 9 14 9 9 2 3 16 4 13 1 9 2 16 4 1 0 9 13 0 9 2
28 15 13 2 16 4 9 11 2 9 1 9 9 2 3 13 9 7 9 7 13 15 2 16 14 13 0 9 2
32 14 3 15 13 2 16 4 1 15 15 3 13 9 1 0 9 2 16 4 1 0 9 13 9 2 3 7 4 10 9 13 2
15 7 7 4 13 3 0 1 0 9 2 16 13 1 9 2
28 3 4 13 0 9 1 0 9 2 16 13 9 1 9 2 13 0 9 2 1 15 7 0 9 4 13 0 2
23 9 1 11 4 13 14 9 0 9 1 3 3 0 0 9 1 0 9 1 9 0 9 2
22 11 11 2 16 13 9 14 0 7 0 9 2 13 1 0 9 1 9 13 0 9 2
28 1 10 9 13 14 3 14 9 9 0 9 1 0 9 2 16 13 1 0 9 1 9 9 11 11 0 9 2
18 16 0 9 1 3 0 9 15 3 13 1 10 16 12 2 0 9 2
68 11 11 2 0 0 9 2 4 1 12 1 0 9 13 0 9 1 9 0 9 7 1 0 13 2 16 13 3 0 2 3 13 0 2 16 9 0 9 2 12 9 9 2 13 1 9 2 16 13 1 0 9 7 1 0 9 13 2 16 9 13 3 13 1 0 0 9 2
20 1 10 9 4 15 13 9 13 0 7 1 9 9 2 14 7 1 9 9 2
38 16 15 4 11 11 1 10 9 13 1 9 10 9 2 13 9 2 16 13 1 0 9 1 9 7 9 2 16 4 10 9 13 1 9 0 0 9 2
22 11 4 2 16 15 9 14 4 3 13 2 3 3 13 9 2 16 4 3 14 13 2
22 9 2 16 13 11 2 11 2 11 2 11 2 11 2 7 4 1 11 14 14 13 2
20 3 15 15 13 2 3 16 15 4 11 11 13 10 9 2 16 4 3 13 2
7 10 0 9 14 15 13 2
14 3 15 13 15 2 16 13 16 15 0 1 9 9 2
21 0 9 10 9 7 9 2 16 15 13 1 9 1 15 2 13 13 10 0 9 2
19 16 4 1 10 0 9 13 9 11 11 2 4 3 13 0 9 1 15 2
16 1 9 2 16 13 0 9 2 1 9 10 9 4 13 13 2
15 9 15 4 13 0 2 16 13 13 2 15 13 13 9 2
11 1 9 1 9 4 13 1 9 0 9 2
20 1 9 9 4 13 0 1 15 12 9 0 9 2 16 13 1 15 0 9 2
15 10 9 10 9 4 13 7 13 1 15 7 13 1 15 2
6 1 9 4 3 13 2
18 9 2 1 15 4 13 2 3 13 14 15 2 16 4 13 15 15 2
13 1 9 13 15 0 9 1 9 1 0 9 9 2
15 3 4 1 0 9 13 14 12 0 9 7 9 1 9 2
19 9 4 13 9 9 11 2 16 13 10 9 1 9 1 9 0 0 9 2
26 1 12 1 0 9 0 0 9 14 4 1 0 9 13 11 11 11 2 11 11 2 11 11 7 11 11
16 9 1 0 4 13 10 9 2 16 4 13 1 9 9 9 2
17 9 14 1 15 14 13 9 0 9 1 9 9 1 12 0 9 2
31 16 4 3 3 13 9 7 16 9 1 9 13 1 10 9 1 9 9 7 10 9 2 4 11 13 9 1 0 9 9 2
3 2 8 2
22 11 4 14 1 0 0 9 1 0 9 13 9 2 15 1 10 9 14 4 13 9 2
31 7 10 9 4 13 0 2 0 7 0 11 7 4 13 14 1 0 9 2 16 4 13 1 15 0 0 9 11 2 11 2
33 11 1 0 0 9 2 16 4 9 13 1 11 11 2 4 13 1 9 2 11 7 4 1 0 9 13 1 0 9 1 0 9 2
11 0 1 9 0 0 9 9 0 9 1 9
18 16 10 0 9 13 2 13 13 2 16 15 9 7 9 2 13 2 2
21 14 7 9 14 13 13 2 16 10 9 3 14 4 13 3 0 9 1 10 9 2
16 1 9 1 9 13 7 9 1 9 3 3 0 1 0 9 2
16 9 15 3 3 13 1 0 0 9 2 1 9 7 1 9 2
9 1 15 15 13 14 0 9 9 2
5 0 9 7 9 2
15 9 10 0 9 7 9 1 15 13 3 0 16 10 9 2
9 10 9 15 14 13 1 0 9 2
15 1 0 15 1 9 3 13 2 16 14 13 14 10 9 2
18 3 14 13 3 9 1 9 2 7 16 3 1 9 9 1 9 13 2
10 3 15 14 13 7 1 15 3 13 2
34 13 15 10 9 2 9 4 13 1 9 0 7 0 9 13 14 1 9 1 9 1 9 9 2 16 4 15 3 13 0 9 1 9 2
5 7 3 13 3 2
6 15 13 14 3 0 2
15 9 1 0 0 9 13 0 7 0 7 3 14 13 3 2
9 0 9 13 2 16 13 3 0 2
14 9 9 7 0 9 1 0 0 9 13 14 10 9 2
23 1 10 9 13 1 0 9 0 9 10 0 9 2 9 15 13 7 3 15 13 0 9 2
13 9 3 13 3 9 1 9 2 13 9 7 9 2
11 1 0 9 13 9 1 0 9 1 9 2
22 11 13 0 12 9 7 15 14 12 9 10 9 13 0 9 2 16 15 13 1 9 2
16 3 3 13 14 3 2 16 15 9 13 1 9 0 9 3 2
27 3 15 7 10 9 1 0 9 13 1 0 9 7 3 0 0 9 15 1 10 9 13 1 10 0 9 2
13 7 13 9 1 0 9 9 14 12 1 12 9 2
19 0 7 0 9 0 9 4 13 0 9 2 13 4 15 1 0 7 0 2
22 9 14 4 15 13 7 9 14 4 15 13 2 16 4 15 15 13 9 1 0 9 2
8 3 13 3 14 9 1 9 2
18 16 13 10 9 2 13 3 1 9 9 9 2 16 13 10 0 9 2
13 3 10 9 13 2 16 15 9 13 7 13 13 2
14 10 0 9 13 2 16 4 15 3 9 13 1 9 2
17 0 9 13 2 16 9 14 14 13 1 9 9 16 14 13 3 2
13 10 9 13 2 16 15 13 1 7 1 0 9 2
32 16 9 14 13 9 1 0 9 2 16 9 13 0 9 2 13 15 14 3 0 12 2 0 0 9 2 16 15 9 13 9 2
13 14 13 15 14 9 2 16 3 14 13 1 9 2
21 0 0 9 2 1 15 9 13 2 13 0 3 3 7 13 3 14 14 3 3 2
21 0 7 13 1 14 3 0 0 9 1 9 7 9 2 1 15 13 9 0 9 2
22 3 15 15 4 9 13 3 2 16 15 4 13 1 10 0 9 7 15 13 1 9 2
7 15 4 13 9 0 9 2
28 9 4 13 2 16 4 14 3 13 2 3 0 9 13 3 2 7 0 7 0 9 4 14 9 3 13 3 2
17 14 4 13 14 3 13 15 3 3 1 0 7 14 15 4 13 2
21 13 4 9 1 3 10 9 2 15 4 13 1 9 9 2 16 4 14 13 9 2
16 13 4 9 3 3 2 12 1 12 2 7 15 13 7 13 2
7 3 4 15 13 1 9 2
5 3 4 13 9 2
24 7 13 14 3 0 2 16 13 2 14 16 4 15 13 3 14 3 13 2 16 4 13 15 2
38 3 15 13 9 2 10 13 10 9 2 16 15 1 3 0 9 9 2 16 15 3 13 2 16 4 13 0 2 1 3 0 9 13 1 9 7 13 2
7 14 15 15 13 2 13 2
8 7 0 13 2 16 15 13 2
9 1 9 13 15 13 2 7 13 2
5 15 4 3 13 2
44 1 15 4 14 3 13 7 14 3 4 13 3 13 10 9 2 9 7 4 13 3 7 3 0 7 0 2 16 4 15 13 15 0 9 7 4 13 15 3 3 0 7 0 2
7 1 15 14 4 4 13 2
13 1 9 4 13 0 2 3 7 4 13 0 9 2
12 16 4 13 9 2 4 13 1 9 0 9 2
6 3 4 13 10 9 2
9 9 15 15 4 13 0 7 0 2
9 13 4 1 0 9 9 7 13 2
40 3 4 15 7 13 1 0 9 7 3 2 16 4 11 13 1 9 9 9 9 7 15 13 1 9 9 2 3 15 15 4 13 2 16 13 1 15 0 13 2
22 1 10 9 1 9 3 4 13 7 13 2 7 1 10 9 4 1 11 13 0 9 2
25 11 4 13 9 2 11 7 15 4 13 9 2 1 9 2 16 15 11 1 0 9 13 9 9 2
14 11 13 2 16 15 15 1 15 1 15 13 3 13 2
35 13 15 15 2 16 15 14 1 10 0 9 13 2 16 13 10 16 10 0 9 2 7 16 1 9 13 14 3 3 2 16 4 13 13 2
12 7 3 14 13 14 3 2 16 4 15 13 2
41 10 9 4 13 1 9 1 0 9 2 16 7 15 4 13 7 4 0 9 13 1 9 0 9 2 4 13 9 1 0 9 2 16 4 13 1 10 9 7 9 2
22 7 9 9 15 4 13 1 10 0 9 2 15 13 10 0 9 1 9 7 13 9 2
16 4 15 13 13 7 13 2 15 13 3 7 1 10 9 13 2
8 3 4 15 13 1 0 9 2
20 1 15 4 13 15 1 9 14 15 15 4 13 3 2 15 4 13 0 13 2
20 13 4 3 1 10 9 7 14 15 15 15 4 13 15 2 16 4 3 13 2
9 7 11 7 15 15 4 13 13 2
13 9 4 13 9 1 9 7 4 3 10 9 13 2
4 3 13 15 2
7 15 13 3 1 10 9 2
8 14 3 14 4 15 13 3 2
9 1 11 4 9 1 0 9 13 2
8 9 13 14 1 12 9 9 2
20 0 9 4 3 13 9 2 16 15 4 13 2 16 4 13 10 9 1 9 2
16 3 15 4 13 2 15 13 15 7 13 0 9 1 10 9 2
9 9 15 4 3 3 13 1 9 2
13 1 9 2 1 15 4 13 2 4 13 0 9 2
17 0 9 4 13 2 16 15 3 13 9 7 15 4 13 14 0 2
10 13 15 4 1 9 7 1 15 13 2
6 13 15 4 10 9 2
10 9 15 4 13 1 9 1 9 9 2
11 3 4 13 2 16 4 13 15 14 0 2
9 1 0 9 4 13 14 1 9 2
19 9 4 13 2 16 13 15 3 2 16 9 14 13 3 3 1 10 9 2
29 9 4 13 2 3 14 13 2 16 4 13 10 9 9 0 9 2 7 9 0 4 13 13 2 15 15 4 13 2
22 13 4 15 2 16 4 13 1 9 2 16 4 3 13 2 15 4 9 1 15 13 2
24 9 15 4 3 13 2 13 15 9 7 1 15 13 0 9 2 16 15 4 1 15 13 9 2
16 13 4 15 1 9 7 3 13 9 2 3 4 13 0 9 2
21 1 12 9 4 13 2 2 3 2 16 4 13 14 3 0 2 4 13 15 0 2
6 7 9 15 4 13 2
11 3 4 13 2 16 15 13 3 2 2 2
9 2 13 15 4 13 1 0 9 2
11 2 14 13 15 13 2 2 4 13 3 2
11 1 0 9 15 4 11 13 0 7 0 2
7 10 9 4 13 1 9 2
13 2 15 0 4 13 1 9 2 16 4 13 3 2
17 2 9 4 13 10 9 7 15 13 2 3 4 13 9 15 0 2
18 9 11 2 9 9 11 2 9 13 2 1 3 13 0 9 7 3 2
11 3 13 1 9 9 9 9 1 10 9 2
25 9 9 13 0 9 2 1 9 0 9 7 13 9 9 2 0 1 0 9 2 16 13 0 9 2
14 2 13 15 9 2 1 15 15 13 13 3 7 3 2
19 1 9 1 9 13 3 0 7 0 7 3 13 0 9 13 2 9 2 2
45 7 11 16 3 0 13 9 0 9 2 16 4 3 3 0 9 0 9 2 13 2 1 0 9 2 7 15 13 16 0 9 2 1 15 13 9 3 14 9 2 9 1 9 2 2
62 11 2 1 9 0 9 0 0 9 1 9 0 9 1 9 0 9 11 11 1 9 0 0 9 1 9 11 2 11 2 11 7 11 2 11 4 12 9 0 0 9 1 0 9 11 1 11 13 1 0 0 9 9 1 9 0 0 2 0 0 9 2
37 11 2 0 0 0 0 9 2 16 4 13 1 9 9 9 1 0 9 7 9 2 11 2 1 10 0 9 2 15 4 3 13 1 9 0 9 2
30 3 13 3 14 14 0 0 9 9 9 0 9 7 9 2 1 15 14 4 13 0 0 9 9 9 1 9 1 9 2
13 3 4 1 11 2 1 0 9 2 13 0 9 2
22 1 9 0 0 9 11 2 9 0 0 11 2 7 9 1 11 4 13 9 9 11 2
18 10 0 9 13 0 0 9 9 2 16 1 11 3 3 13 0 9 2
33 9 9 11 13 0 14 14 1 15 2 16 4 13 9 0 9 7 14 10 0 9 2 7 4 13 13 9 1 3 0 0 9 2
32 9 1 0 9 13 0 2 16 13 9 1 9 14 0 2 3 3 7 13 0 14 9 2 16 1 0 9 9 13 0 9 2
40 1 0 7 0 13 0 9 2 16 4 1 0 9 13 14 1 9 0 9 2 0 9 7 9 2 1 9 7 14 13 0 11 1 9 1 2 0 2 11 2
31 9 4 13 14 3 2 16 13 2 16 13 13 2 0 2 9 2 0 9 2 3 0 7 0 9 16 3 0 0 9 2
26 11 4 13 9 11 11 2 9 11 11 2 9 11 11 7 11 11 2 9 11 11 7 9 11 11 2
6 13 4 0 0 9 2
7 14 2 9 15 14 13 2
10 13 9 2 9 2 14 13 0 9 2
24 9 13 3 0 1 12 1 12 9 2 16 15 4 9 7 1 15 14 9 9 3 3 13 2
9 13 4 1 9 9 1 0 9 2
8 0 0 9 13 0 2 2 2
25 11 2 11 13 14 1 12 9 0 1 10 0 0 0 9 2 16 13 13 11 2 11 7 11 2
18 1 9 7 9 13 0 9 3 0 9 2 1 15 13 15 0 9 2
29 0 9 13 1 9 9 14 0 0 9 2 1 15 13 0 9 2 3 7 3 7 15 13 0 2 7 0 9 2
34 0 9 1 10 9 13 1 0 9 2 3 16 15 13 1 9 0 13 1 0 9 2 16 13 1 9 15 0 7 0 1 10 9 2
21 0 9 1 9 13 2 7 7 13 0 13 1 0 9 2 16 13 1 10 9 2
20 3 4 3 13 14 1 9 0 2 1 15 4 13 2 16 4 14 3 13 2
14 7 1 9 4 15 3 13 1 0 0 9 1 9 2
21 16 4 13 9 2 16 4 13 9 9 7 9 2 4 15 13 1 0 0 9 2
15 3 3 13 2 16 14 4 13 2 7 13 14 1 11 2
11 3 3 4 1 0 9 13 9 0 9 2
16 1 3 9 13 3 0 2 7 9 13 14 1 10 10 9 2
14 13 7 14 12 9 2 3 13 14 0 9 7 9 2
14 13 1 0 9 1 9 7 13 0 1 0 9 9 2
45 1 11 4 13 9 3 0 2 7 15 4 10 0 9 11 2 1 15 4 1 9 12 7 12 13 0 0 9 2 2 13 2 2 16 15 4 1 12 9 13 1 9 1 0 2
29 1 9 0 9 4 11 11 2 11 11 7 11 11 14 13 0 9 2 3 7 15 4 2 13 2 10 0 11 2
14 0 11 4 15 13 2 16 4 13 3 1 10 9 2
19 9 1 9 4 9 1 9 9 13 9 9 1 9 12 9 1 0 9 2
22 9 0 9 14 13 14 0 2 3 7 13 2 16 13 0 9 1 0 9 0 3 2
23 14 7 4 9 9 1 9 1 0 9 13 14 1 9 2 0 9 2 9 7 9 9 2
36 13 4 14 1 9 2 16 13 1 9 2 7 1 14 3 0 9 0 9 7 1 9 9 2 16 1 10 9 13 9 2 15 9 13 9 2
13 11 9 9 11 11 15 4 14 3 13 11 11 2
14 2 13 15 4 2 16 4 1 9 13 0 9 8 2
53 1 11 4 15 3 3 3 13 9 0 9 11 2 11 2 2 16 4 13 9 1 3 12 9 7 12 7 12 9 1 9 1 0 9 2 1 15 4 13 9 7 0 9 2 14 3 2 13 2 9 9 11 2
20 9 1 11 7 11 11 4 13 14 3 2 1 9 0 9 2 1 0 9 2
23 11 13 1 9 0 9 1 0 9 14 3 0 0 9 2 1 15 11 4 13 0 9 2
15 13 4 9 0 9 7 9 1 0 7 10 0 0 9 2
11 3 1 0 9 4 13 0 13 0 9 2
26 9 1 0 9 2 0 9 7 0 9 4 13 1 11 10 9 2 16 4 15 13 13 14 0 9 2
6 11 4 13 9 11 2
11 13 4 12 9 2 16 4 15 13 9 2
4 9 15 4 13
11 13 15 4 0 0 9 9 1 9 9 2
11 13 4 1 9 2 16 15 4 13 9 2
16 13 4 3 2 7 15 4 13 9 2 16 4 13 1 9 2
5 15 4 13 9 2
6 9 4 13 1 9 2
9 1 9 4 13 13 3 7 3 2
15 7 2 16 15 9 14 13 1 9 2 16 13 1 9 2
14 7 2 16 15 14 13 1 9 2 16 13 1 9 2
8 15 7 3 13 1 0 9 2
3 10 9 2
12 3 4 15 12 13 2 16 15 13 2 2 2
22 3 7 13 14 0 2 7 15 4 13 9 2 16 4 10 0 9 15 13 1 9 2
11 11 13 0 2 9 1 0 9 3 13 2
29 16 13 11 1 9 14 3 0 2 7 4 1 12 9 3 3 13 1 9 2 1 15 4 14 13 0 0 9 2
17 9 12 4 7 9 1 9 1 11 13 2 16 13 1 9 9 2
32 1 9 15 4 15 13 3 2 7 16 15 4 9 13 9 0 9 2 16 15 4 13 16 9 1 0 9 13 0 0 9 2
12 13 7 15 4 14 1 0 9 10 9 11 2
33 1 0 9 0 9 11 2 1 9 2 14 4 13 9 1 0 9 7 13 1 10 9 16 9 2 7 4 10 9 13 1 9 2
12 14 2 16 15 4 9 13 1 10 0 9 2
14 16 15 4 15 3 13 2 13 1 10 9 3 0 2
20 7 0 9 13 0 9 2 1 15 9 1 0 7 3 13 10 0 9 9 2
19 12 1 10 0 9 14 4 13 15 2 16 4 10 9 13 1 10 9 2
18 7 11 9 0 9 1 9 13 2 15 2 15 13 2 13 0 9 2
16 7 13 2 16 15 15 4 13 2 7 4 9 13 1 9 2
17 0 13 2 16 9 3 13 2 9 7 4 13 13 1 10 9 2
19 12 9 13 0 0 9 1 0 9 2 16 15 13 1 0 9 1 9 2
11 0 9 1 9 1 9 13 0 0 9 2
17 0 9 4 9 14 1 3 13 1 0 9 2 16 4 13 1 11
14 9 13 0 2 16 9 9 1 9 1 0 9 3 13
17 12 0 9 2 10 9 7 9 7 4 1 9 3 13 0 9 2
25 10 12 9 7 4 13 1 0 9 2 16 1 9 3 2 16 13 0 9 2 4 13 13 9 2
16 15 13 0 9 1 11 7 9 2 4 13 0 11 1 11 2
12 0 9 11 11 4 3 1 9 13 0 9 2
12 13 4 1 9 7 3 13 15 2 15 13 2
14 9 2 16 13 1 9 11 11 1 11 2 13 0 2
11 11 15 1 10 9 13 1 0 0 9 2
26 10 9 13 2 16 9 13 1 9 3 0 9 2 15 11 14 3 13 2 16 13 1 0 9 9 2
4 7 13 9 2
7 3 3 9 14 3 13 2
7 0 9 3 1 9 13 2
13 7 13 3 0 7 9 13 1 9 3 4 13 2
24 11 4 13 2 16 14 13 13 0 9 2 16 15 13 9 2 10 9 7 1 9 14 13 2
17 13 15 2 3 13 9 9 11 3 0 2 7 14 14 13 15 2
34 9 1 9 9 13 9 0 9 11 11 0 9 1 11 2 16 4 11 13 2 16 13 0 9 1 11 3 1 0 0 9 9 12 2
19 11 4 14 13 2 16 13 14 0 3 13 9 2 1 9 7 15 13 2
21 0 9 4 13 13 12 9 9 2 7 4 15 3 13 14 3 10 16 12 9 2
15 0 12 9 7 1 9 11 0 9 14 4 13 0 13 2
20 9 9 4 3 13 13 9 11 2 9 9 2 16 1 9 13 0 0 9 2
18 3 4 15 13 2 16 13 1 12 9 14 9 1 10 0 0 9 2
19 1 3 12 9 9 4 1 9 13 12 0 2 12 0 7 12 0 9 2
17 12 9 4 13 9 7 15 15 3 14 13 7 13 9 1 9 2
19 7 13 3 0 14 12 1 10 9 2 7 4 13 9 1 9 0 12 2
15 16 14 13 9 0 9 0 11 2 15 4 13 0 9 2
22 9 9 4 13 1 9 1 1 11 0 0 9 11 11 2 16 4 13 0 9 9 2
46 3 4 15 1 0 9 1 9 13 0 7 0 9 2 9 15 2 9 2 16 4 15 1 0 9 13 0 1 0 2 9 7 4 13 10 9 2 16 4 13 7 3 13 1 9 2
18 3 15 15 4 3 13 1 9 9 1 0 0 9 0 0 9 11 2
15 9 1 12 9 3 2 16 4 13 0 9 2 4 13 15
12 3 3 13 1 0 0 9 0 0 9 9 2
24 0 9 1 0 9 9 16 0 9 7 0 9 9 1 0 9 15 13 14 1 9 0 9 2
13 3 0 9 1 9 1 0 9 7 13 0 9 2
10 1 10 9 13 1 15 9 0 9 2
34 9 0 9 14 13 14 9 0 9 2 9 0 9 2 0 9 9 9 7 9 2 14 14 9 1 0 9 2 7 14 9 0 9 2
17 9 13 2 16 13 1 9 0 9 0 9 0 9 7 9 9 2
20 15 13 0 13 0 9 2 16 13 9 0 9 9 9 9 7 9 9 9 2
28 10 9 13 0 7 1 15 4 13 10 9 7 9 16 7 0 9 2 7 7 3 14 13 9 9 7 9 2
32 14 1 9 15 4 13 9 1 9 14 1 0 9 2 7 1 9 2 1 9 2 16 4 0 9 14 3 13 10 0 9 2
23 3 7 13 3 2 16 3 2 16 9 13 3 0 9 2 13 1 0 9 9 0 9 2
16 1 10 9 13 14 12 9 2 16 13 3 0 1 0 9 2
25 9 1 9 13 13 1 0 9 2 2 13 9 13 3 2 16 14 4 13 1 9 7 9 2 2
8 9 14 13 13 9 0 9 2
21 0 9 1 9 10 9 13 9 9 7 9 9 2 15 15 13 1 9 8 9 2
18 7 7 13 14 10 9 0 9 7 9 2 16 4 13 1 9 9 2
25 1 0 9 14 4 13 0 2 16 4 12 13 1 9 9 0 7 15 1 9 7 9 13 9 2
17 9 0 9 7 1 0 9 16 1 9 15 3 13 1 0 9 2
12 3 0 9 4 13 0 1 9 1 0 9 2
32 14 7 4 9 9 3 13 2 16 9 1 0 0 9 2 1 0 9 2 1 11 7 1 0 9 1 9 3 7 3 13 2
14 2 7 13 10 9 2 16 15 4 13 7 13 3 2
15 7 1 9 0 0 9 11 1 9 4 13 14 0 9 2
11 1 0 9 4 15 9 13 0 0 9 2
34 3 16 4 1 9 1 12 2 12 13 0 9 11 2 11 2 4 13 1 9 1 12 2 12 2 12 0 1 0 9 11 2 11 2
26 2 13 4 3 3 2 14 1 9 4 13 0 2 3 16 1 10 9 9 4 13 14 1 12 9 2
11 1 12 2 12 15 4 13 11 11 11 2
25 10 9 4 13 0 9 11 11 11 11 2 16 4 15 13 3 3 1 9 11 11 1 0 11 2
15 1 10 3 0 0 9 4 13 0 9 9 12 12 9 2
43 1 0 9 9 2 2 13 14 4 15 15 3 1 12 9 2 2 2 15 4 9 13 9 1 9 9 7 13 0 9 9 2 16 14 4 13 3 1 9 14 1 9 2
16 1 9 1 0 9 9 4 9 3 13 0 9 9 0 9 2
13 1 11 13 0 9 2 0 0 9 2 0 9 2
15 3 4 1 9 11 11 1 9 0 9 10 9 13 9 2
18 1 9 4 3 13 2 16 15 4 1 9 9 13 13 0 9 9 2
11 9 4 13 1 9 1 0 9 0 9 2
27 7 15 13 1 10 9 2 1 0 9 2 3 1 9 7 9 2 7 14 9 14 13 10 9 3 0 2
25 1 9 7 9 0 9 4 10 9 7 9 13 11 11 1 11 2 16 13 9 9 14 0 9 2
20 1 0 0 9 4 13 14 9 9 2 7 13 3 1 2 9 2 0 9 2
18 13 14 4 14 0 0 9 1 9 8 11 2 16 13 1 9 9 2
19 9 2 0 15 13 9 2 16 1 9 14 13 3 2 13 1 9 2 2
7 3 13 13 1 0 9 2
13 9 12 4 9 13 0 9 7 9 1 0 9 2
9 1 9 4 1 9 13 0 9 2
28 9 4 13 14 9 2 7 4 15 0 9 7 0 9 1 9 7 9 2 16 4 13 1 9 2 13 13 2
17 1 0 9 12 9 4 9 13 10 9 2 16 15 13 14 3 2
17 1 15 4 13 9 9 11 2 9 11 7 9 1 10 0 9 2
21 10 0 9 4 13 14 11 11 2 16 4 1 10 9 13 10 0 9 1 9 2
18 9 0 9 4 14 13 1 15 2 16 0 14 3 13 1 10 9 2
14 0 4 13 14 0 9 2 16 15 13 3 12 9 2
14 3 4 1 9 13 9 0 9 11 0 9 11 11 2
15 0 4 13 9 12 2 12 2 16 4 13 0 0 9 2
28 3 15 15 4 9 3 13 1 0 9 1 9 2 13 4 15 9 1 9 2 1 0 9 2 9 1 9 2
23 16 4 13 2 4 1 9 1 9 7 9 13 9 9 2 16 4 13 9 1 0 9 2
19 1 3 13 0 9 1 9 1 9 2 3 0 9 14 4 9 13 9 2
10 1 10 9 4 13 13 1 12 9 2
44 0 9 7 13 1 9 14 0 0 9 0 2 0 9 11 1 9 7 0 9 1 0 9 2 16 13 14 2 3 14 13 9 2 1 15 9 9 1 11 14 4 13 0 2
22 0 9 13 3 1 9 9 1 9 9 1 9 7 15 3 13 1 9 9 0 9 2
12 9 11 11 13 3 3 0 0 9 0 9 2
32 1 10 2 9 2 0 9 3 3 14 4 13 2 7 3 1 0 9 15 4 14 14 3 7 3 15 13 14 1 10 9 2
15 14 4 13 0 9 3 0 16 2 3 0 2 1 9 2
17 1 15 11 11 13 9 2 16 15 15 13 1 9 3 0 9 2
11 3 7 9 1 0 9 13 14 1 9 2
16 15 15 4 13 1 14 0 2 14 0 9 0 2 11 2 2
20 16 0 9 0 9 13 10 9 2 15 13 1 9 10 9 16 9 1 9 2
14 2 1 10 9 4 9 13 9 1 9 9 1 9 2
15 13 7 4 2 16 15 3 14 13 2 16 13 1 9 2
14 1 9 9 15 4 13 13 14 9 1 0 0 9 2
15 3 12 15 4 13 0 9 2 12 9 7 4 9 13 2
21 1 11 11 4 9 13 12 9 12 0 9 2 16 4 15 13 1 0 0 9 2
22 0 9 15 4 13 14 1 9 3 2 0 9 9 2 7 4 9 13 14 1 9 2
16 9 4 14 13 2 16 4 1 9 13 10 0 9 7 9 2
20 9 13 3 1 9 9 7 9 2 9 15 0 7 3 2 16 13 9 0 2
22 16 13 9 1 9 2 13 9 1 9 1 9 1 12 1 12 9 1 9 12 9 2
25 9 13 1 0 9 1 12 1 12 9 7 15 1 10 9 13 1 9 2 16 15 13 1 9 2
26 1 12 1 12 9 13 9 1 9 7 9 7 15 13 1 0 9 2 3 7 14 1 15 13 9 2
12 13 14 9 2 16 0 9 14 13 1 9 2
5 13 15 16 9 2
16 0 9 13 0 2 7 15 13 9 2 16 15 13 2 13 2
30 10 9 13 1 15 2 3 4 9 13 1 10 9 2 1 15 7 13 2 16 15 3 13 7 13 10 9 0 9 2
10 1 9 3 4 15 13 13 1 9 2
14 16 14 4 13 9 10 9 2 13 9 0 14 15 2
8 15 15 4 3 13 11 11 2
24 10 0 9 4 13 1 9 7 3 4 13 11 0 9 2 14 16 4 4 13 12 0 9 2
17 13 15 0 2 1 15 9 13 2 16 13 1 2 0 11 2 2
26 11 13 7 0 7 0 2 13 0 9 2 16 14 14 9 1 0 9 13 9 2 1 15 13 0 2
15 1 10 9 13 9 1 0 9 9 14 14 1 9 0 2
26 7 7 13 3 2 16 15 4 13 1 11 2 7 14 13 3 2 16 15 4 13 15 1 10 9 2
17 11 11 4 3 13 2 16 13 10 9 13 3 2 16 3 13 2
8 3 13 2 16 13 1 11 2
11 3 14 4 13 7 0 0 9 16 11 2
11 3 15 13 13 2 16 13 10 9 0 2
40 13 3 2 16 4 1 0 9 1 11 7 11 13 0 11 2 7 16 10 16 9 1 12 9 2 16 15 1 11 14 13 7 7 13 1 9 2 13 11 2
21 3 7 4 15 13 2 16 4 3 13 14 0 11 2 16 4 1 11 13 11 2
26 13 7 4 14 13 2 16 12 9 1 10 9 2 1 15 13 14 11 7 11 2 13 9 0 9 2
32 16 14 4 13 0 0 9 2 4 1 9 1 12 9 0 9 2 11 2 1 0 11 3 13 10 16 12 9 1 10 11 2
51 9 4 13 13 2 7 4 1 9 1 9 1 11 13 2 16 4 9 13 2 16 9 14 4 13 9 9 1 9 9 12 7 9 0 9 2 16 4 9 9 12 13 2 16 13 13 0 9 9 9 2
41 1 9 4 1 0 9 9 1 9 9 13 2 16 4 9 14 3 13 1 3 0 0 9 2 16 7 4 15 3 13 2 9 9 9 13 3 1 9 0 9 2
33 9 9 4 1 0 9 13 9 2 16 15 1 3 0 9 13 9 7 13 1 9 2 16 4 3 13 9 1 0 0 9 9 2
28 9 2 16 4 9 13 1 0 0 9 2 15 4 13 2 1 0 9 13 1 9 1 9 0 0 9 13 2
13 1 9 0 0 9 4 1 10 9 13 0 9 2
13 0 9 1 0 9 7 9 9 13 0 7 0 2
20 0 9 4 1 12 1 12 9 13 12 9 2 16 4 13 3 13 1 11 2
13 1 15 4 13 3 11 2 11 2 11 7 11 2
3 2 8 2
11 9 4 1 11 14 13 9 1 0 9 2
42 0 0 0 9 4 13 2 16 4 9 7 9 9 13 1 12 0 9 0 9 2 0 9 11 2 16 13 10 9 1 0 11 2 7 4 14 13 0 9 1 9 2
32 0 9 1 0 9 4 13 1 9 1 12 9 1 9 9 2 1 15 4 13 0 2 16 13 9 9 0 9 9 0 9 2
32 9 2 16 4 3 13 9 1 9 0 9 2 1 15 13 9 1 9 13 9 9 2 4 1 0 9 0 9 13 12 9 2
28 9 1 9 13 0 13 14 1 9 0 9 9 2 1 15 15 9 13 2 16 15 15 13 1 9 10 9 2
14 13 13 2 3 13 9 2 9 7 13 1 0 9 2
3 2 8 2
12 9 1 11 1 11 13 3 0 1 12 0 9
12 3 4 13 9 2 16 15 4 3 3 13 2
11 3 7 3 4 1 9 10 9 13 9 2
5 13 4 1 9 2
5 12 9 1 12 2
13 3 4 13 9 1 9 2 13 9 7 13 13 2
4 13 14 3 2
17 9 2 16 15 12 7 13 14 10 0 9 2 1 15 13 0 2
20 11 4 13 13 0 0 9 11 7 15 2 16 9 0 14 13 10 0 9 2
27 11 4 13 3 0 2 4 14 13 0 9 1 0 9 2 1 15 4 3 13 2 16 4 13 0 9 2
21 13 4 2 16 15 11 15 14 4 13 13 2 15 14 4 1 15 13 0 9 2
19 11 4 13 2 16 9 13 10 9 2 16 13 0 0 0 9 13 0 2
14 2 15 14 13 9 2 16 9 1 9 13 1 9 2
3 13 3 2
10 13 15 15 14 3 13 0 9 9 2
18 0 9 8 11 11 1 11 4 1 10 9 1 0 0 9 13 0 2
40 1 0 0 9 7 9 14 10 9 13 0 9 0 9 2 14 14 1 9 1 11 2 7 14 1 11 2 11 2 11 7 0 9 1 9 11 7 1 11 2
25 0 9 14 13 9 11 1 3 0 2 0 2 0 9 7 0 9 2 16 13 3 9 0 9 2
13 10 9 4 1 9 9 1 10 9 13 1 9 2
24 11 8 11 1 9 11 4 1 9 1 9 12 3 13 1 9 0 9 1 0 9 7 3 2
11 9 4 14 3 3 13 2 3 15 13 15
7 13 4 3 1 0 9 2
7 15 4 13 12 9 12 2
37 9 2 0 7 0 1 10 0 9 7 0 0 9 2 16 13 14 0 9 7 16 15 13 0 0 9 1 0 9 7 3 2 4 9 3 13 2
36 13 15 4 9 2 16 13 1 9 10 9 10 9 2 16 4 15 15 13 1 0 2 7 9 2 16 13 10 9 15 1 9 1 0 9 2
29 1 10 0 9 4 13 9 9 2 16 15 4 13 1 0 9 2 9 7 9 7 15 3 1 9 13 15 0 2
32 10 0 9 13 14 1 9 9 2 16 15 4 1 12 9 9 3 13 13 9 9 16 9 9 2 14 16 4 3 13 0 2
42 16 4 13 9 2 16 15 4 13 2 7 13 9 10 0 9 2 4 13 3 13 1 10 9 2 0 16 0 9 0 9 11 7 0 1 10 9 16 9 0 9 2
7 13 4 1 0 0 9 2
8 0 9 4 13 1 11 11 2
10 9 9 4 13 13 1 9 1 9 2
9 0 4 13 10 9 2 12 2 2
6 9 7 9 11 11 2
14 1 9 1 11 4 1 11 11 7 11 13 0 9 2
12 11 4 14 13 9 2 13 7 4 0 9 2
16 1 0 0 9 4 13 9 7 9 7 13 9 7 9 11 2
31 11 4 13 13 0 9 1 9 2 16 4 13 0 9 2 7 4 13 3 1 9 13 9 11 2 16 15 4 13 3 2
25 10 0 9 4 13 9 8 8 2 12 2 2 16 15 4 13 14 10 16 12 9 7 0 9 2
24 11 4 10 9 13 1 0 0 9 2 0 16 0 9 0 9 2 16 15 4 13 0 9 2
18 1 10 3 0 9 13 11 11 2 12 2 7 9 11 2 12 2 2
19 11 4 13 0 9 8 12 2 16 4 0 9 13 1 9 1 12 9 2
12 0 4 13 7 13 0 0 9 1 0 9 2
14 10 0 7 0 9 4 13 1 0 9 1 0 9 2
8 11 4 13 14 3 0 9 2
11 1 0 13 12 0 9 7 12 0 9 2
5 13 4 1 9 2
12 0 9 15 4 13 1 9 12 7 12 9 2
31 1 9 1 0 9 4 13 0 9 2 7 4 1 9 2 16 4 13 9 2 16 4 15 13 13 9 2 13 0 9 2
16 0 4 13 1 9 11 12 0 7 0 9 15 4 13 13 2
12 13 15 4 9 11 12 2 0 0 0 9 2
10 1 12 0 9 4 13 1 0 9 2
30 1 9 2 16 15 4 1 0 0 9 13 1 9 2 4 10 3 0 7 0 9 13 1 9 10 9 2 12 2 2
22 1 0 9 7 9 1 0 9 4 1 9 13 0 9 2 16 4 13 9 1 9 2
7 11 4 13 9 9 12 2
19 13 15 4 1 9 0 9 2 1 15 4 10 9 3 13 11 7 9 2
17 11 4 13 0 9 2 16 4 13 9 2 0 9 11 7 0 2
14 0 0 9 4 13 0 2 7 4 13 13 0 9 2
19 9 1 11 4 0 11 7 11 3 13 2 16 4 9 12 11 13 9 2
10 1 12 0 9 4 9 3 13 11 2
13 9 12 4 2 16 4 13 11 0 2 13 9 2
9 13 15 4 1 9 0 0 9 2
31 1 0 4 13 9 0 9 1 0 9 1 9 2 12 2 2 9 0 9 9 2 12 2 7 9 7 9 2 12 2 2
8 13 1 0 9 0 0 9 2
14 10 3 0 9 11 13 1 9 9 11 1 9 11 2
21 10 9 4 13 0 0 9 9 2 16 4 13 1 0 0 0 9 1 0 9 2
17 1 12 9 4 15 11 13 2 16 4 15 13 1 0 9 11 2
4 9 9 11 2
19 12 0 9 11 13 11 7 13 11 7 11 0 9 13 0 1 10 9 2
13 12 11 12 2 12 2 1 11 13 9 1 11 2
21 12 11 8 11 2 16 13 1 11 2 15 1 9 1 11 13 1 0 9 11 2
18 12 0 9 11 11 2 8 12 2 13 2 16 4 0 9 13 11 2
17 12 0 9 11 11 2 12 2 13 2 16 9 13 1 0 9 2
15 9 9 13 9 2 16 15 13 9 3 13 7 13 9 2
32 7 15 2 16 13 1 9 9 9 2 16 15 2 16 13 2 15 13 1 0 9 13 1 10 9 7 15 10 9 3 13 2
13 1 9 9 3 13 10 9 9 7 15 3 13 2
21 9 10 9 13 1 15 2 16 13 1 15 9 3 3 0 1 10 3 0 9 2
9 3 7 3 13 10 9 11 11 2
9 1 3 13 1 9 3 1 9 2
17 0 9 7 3 4 13 3 7 3 3 3 2 3 7 13 3 2
17 10 9 15 13 13 1 9 2 7 3 13 9 2 16 3 13 2
19 9 9 0 4 13 9 2 7 1 15 11 13 3 3 0 13 0 0 9
21 11 4 13 1 9 1 11 2 7 1 14 3 0 9 13 0 3 13 1 9 2
12 0 9 15 4 11 1 9 13 1 0 9 2
16 11 4 13 9 2 1 15 15 4 3 3 9 13 1 9 2
17 3 4 3 13 1 9 2 13 4 13 2 16 16 15 13 0 2
7 9 4 15 13 7 13 2
4 12 4 13 2
10 3 15 4 13 2 16 4 13 9 2
22 3 4 13 14 3 0 2 16 4 15 3 13 1 9 2 16 4 15 15 3 13 2
8 9 15 4 3 13 1 9 2
7 1 9 4 13 10 9 2
5 13 4 13 9 2
4 9 4 13 2
32 13 4 3 0 1 0 9 1 9 2 3 7 4 13 13 14 9 1 0 9 9 2 16 4 13 1 9 10 9 1 9 2
17 1 9 4 11 13 11 9 2 1 15 4 3 13 14 9 9 2
19 3 4 13 0 9 2 9 2 9 2 9 2 0 9 2 9 2 9 2
26 11 4 13 0 0 9 7 9 2 1 15 4 13 2 16 0 4 13 10 9 16 9 1 9 9 2
29 16 15 4 13 1 9 1 0 9 2 4 13 1 9 0 0 9 14 0 9 7 15 1 15 14 13 1 9 2
19 16 4 13 0 0 9 2 7 15 4 13 14 1 9 2 4 13 11 2
13 9 1 9 15 4 3 13 2 13 7 4 15 2
18 9 1 9 2 9 2 16 4 13 1 11 2 15 4 1 3 13 2
8 11 15 4 13 1 9 9 2
14 9 4 13 1 9 9 2 7 15 14 13 4 13 2
9 13 4 0 2 0 9 0 9 2
12 11 15 4 13 1 9 2 13 4 10 9 2
5 9 4 13 0 2
11 15 4 9 13 9 2 4 13 1 9 2
8 3 4 13 9 7 13 3 2
5 13 4 1 9 2
14 9 4 13 14 2 14 9 4 13 1 9 7 9 2
6 11 15 4 3 13 2
16 15 4 13 2 16 11 14 3 10 9 13 9 1 0 9 2
12 3 4 15 13 1 9 7 13 1 0 9 2
15 9 10 9 2 16 4 13 3 1 15 2 4 13 0 2
7 15 15 4 13 1 15 2
7 14 2 9 4 14 13 2
16 13 4 2 16 4 15 13 2 16 4 15 13 1 10 9 2
17 16 4 13 1 9 2 16 14 4 13 9 2 4 15 13 9 2
19 3 4 15 15 13 1 9 7 0 9 2 16 14 4 13 1 10 9 2
14 15 15 4 14 13 7 7 4 15 15 14 3 13 2
10 13 4 9 1 9 7 15 15 13 2
18 11 4 3 13 1 9 7 15 13 1 9 1 0 1 9 0 9 2
8 1 9 15 15 4 13 9 2
5 9 4 13 0 2
10 1 12 1 15 4 13 3 0 9 2
12 3 4 13 14 0 9 7 0 9 7 9 2
6 3 9 15 4 13 2
6 14 3 4 13 9 2
13 3 15 4 13 2 7 16 4 15 13 14 11 2
8 3 1 9 4 15 3 13 2
11 4 13 2 16 4 11 1 9 3 13 2
12 16 4 15 13 2 4 13 1 10 0 9 2
9 1 9 4 13 9 7 13 15 2
11 9 4 13 0 2 7 15 4 3 13 2
7 3 4 15 13 1 9 2
13 3 4 13 11 2 13 9 7 15 1 9 13 2
6 13 4 9 10 9 2
11 9 15 4 3 13 7 13 13 1 9 2
11 13 4 10 9 2 16 15 4 3 13 2
10 13 4 15 1 9 7 15 13 3 2
8 3 1 9 4 13 9 9 2
6 15 4 15 3 13 2
14 0 9 4 13 9 1 0 0 9 2 0 1 9 2
14 13 15 4 2 16 16 4 13 2 16 15 15 13 2
6 10 9 4 15 13 2
5 13 4 15 15 2
13 13 15 4 1 9 1 9 7 15 14 15 13 2
4 13 15 4 2
9 3 4 13 9 0 9 1 9 2
13 16 4 15 13 10 9 2 13 13 15 1 9 2
15 16 4 13 1 15 2 4 13 13 1 9 7 0 9 2
8 15 4 11 1 9 3 13 2
17 13 4 15 1 11 2 3 0 9 13 7 15 15 4 15 13 2
23 13 4 2 16 13 9 7 16 13 14 9 2 7 15 4 13 2 16 4 15 13 13 2
9 13 4 0 0 7 3 0 9 2
10 13 4 1 9 7 13 9 1 9 2
17 1 10 0 9 4 11 13 15 2 7 4 3 13 9 1 9 2
4 13 4 15 2
10 4 15 13 13 2 13 4 1 11 2
6 11 1 9 4 13 2
12 13 4 2 16 15 0 9 3 13 1 15 2
18 14 16 4 13 1 11 7 0 2 15 15 4 13 2 16 15 13 2
8 16 16 14 4 13 13 9 2
13 13 4 2 3 13 15 10 9 1 9 1 9 2
6 15 7 14 13 4 2
11 14 2 1 0 9 4 15 13 14 15 2
14 11 4 3 1 9 13 10 9 7 15 15 14 13 2
8 13 4 7 15 1 9 13 2
4 15 4 13 2
7 3 15 4 13 1 15 2
9 3 4 15 12 13 1 9 9 2
5 13 4 3 0 2
13 1 10 14 9 4 13 2 3 4 13 14 9 2
8 0 9 4 13 1 10 9 2
14 16 4 3 13 3 9 2 4 14 13 14 10 9 2
9 1 9 4 13 7 14 0 9 2
17 0 9 2 16 15 4 13 11 0 1 15 2 4 13 10 9 2
10 13 4 3 0 2 0 7 3 0 2
7 13 4 15 1 9 9 2
7 14 2 14 15 13 0 2
14 16 4 15 15 13 13 2 4 13 3 0 16 15 2
17 7 15 13 3 0 9 2 9 15 13 1 9 7 13 0 3 2
9 3 4 1 11 3 13 1 9 2
12 13 4 14 2 16 4 13 9 7 15 13 2
15 11 4 14 13 1 9 2 14 2 9 13 10 1 9 2
8 13 4 15 3 1 0 9 2
10 4 15 13 0 2 16 16 15 13 2
7 2 13 4 15 13 0 2
5 9 15 4 13 2
6 3 4 13 10 9 2
13 7 15 1 10 9 15 4 13 13 2 16 13 2
16 13 15 4 3 3 2 16 3 13 2 7 15 4 13 13 2
14 3 4 13 1 9 2 16 4 15 13 1 3 0 2
7 3 15 4 13 1 15 2
10 3 15 4 13 2 16 4 13 0 2
5 1 11 4 13 2
8 0 15 4 3 13 1 9 2
8 3 15 4 11 13 1 9 2
9 3 4 13 1 9 7 15 13 2
16 9 4 13 7 13 13 9 2 16 15 4 13 1 9 9 2
7 3 15 4 13 13 11 2
4 13 4 0 2
5 9 9 2 9 2
9 9 4 1 0 9 13 1 9 2
11 1 0 9 4 13 14 9 7 0 9 2
17 13 4 15 12 9 12 16 0 7 3 0 9 11 7 11 11 2
24 1 9 4 13 1 0 9 2 7 1 10 0 9 13 11 1 11 2 16 13 15 12 9 2
18 10 9 4 13 1 10 9 0 2 7 4 13 0 9 1 0 9 2
7 9 4 15 13 9 11 2
17 0 13 2 16 4 15 3 13 2 16 13 3 0 7 0 9 2
17 1 0 9 15 3 13 1 9 7 13 1 15 16 10 0 9 2
13 9 4 13 1 9 3 7 13 4 15 0 9 2
12 3 4 1 9 3 13 9 1 9 0 9 2
10 14 15 4 13 2 16 15 4 13 2
13 3 4 15 13 2 16 4 14 0 13 15 0 2
18 9 4 13 1 11 2 16 13 9 1 9 7 9 0 16 1 15 2
11 0 9 1 9 9 13 9 9 1 9 2
11 13 4 15 14 9 1 0 7 0 9 2
18 13 4 13 14 10 9 2 7 4 15 1 9 13 14 1 10 9 2
9 3 15 4 13 11 7 0 9 2
23 3 16 9 14 9 13 1 9 2 16 15 9 13 1 0 0 9 2 15 13 3 12 2
27 9 0 9 1 10 9 3 13 1 9 1 0 9 2 0 9 2 1 15 13 7 13 9 1 0 9 2
9 13 1 0 9 2 9 7 9 2
6 13 9 1 12 9 2
8 12 9 9 13 7 13 9 2
3 13 9 2
3 13 9 2
10 9 1 9 13 1 12 9 0 9 2
15 3 13 9 2 13 9 9 7 1 0 9 13 12 9 2
9 13 0 9 7 0 9 7 13 2
6 13 1 0 9 9 2
5 13 9 0 9 2
13 16 13 9 1 9 2 3 13 1 9 0 9 2
27 9 13 1 9 9 9 1 12 0 9 2 14 16 4 15 13 13 7 13 7 14 16 4 13 1 9 2
19 14 13 15 3 1 9 0 9 2 16 15 13 1 9 7 13 1 9 2
21 9 2 16 13 1 9 2 0 9 2 0 9 7 0 9 13 0 9 0 9 2
8 9 13 2 16 15 13 9 2
17 1 12 9 4 1 9 13 2 1 0 9 7 4 13 9 9 2
23 0 15 4 13 1 0 9 2 14 16 4 13 1 9 7 14 16 4 3 15 13 9 2
7 10 9 15 13 3 13 2
5 15 13 0 9 2
32 9 0 9 2 0 9 9 7 9 2 4 13 14 3 0 0 2 14 16 13 3 0 9 9 9 7 9 7 14 9 9 2
17 1 10 16 12 9 10 9 4 15 13 1 9 13 14 15 0 2
23 9 9 9 13 12 2 0 11 2 16 13 1 0 0 9 7 16 15 3 13 1 9 2
23 3 7 15 13 1 0 9 2 16 9 3 13 7 13 16 0 9 13 1 9 7 9 2
24 3 15 13 2 16 13 3 10 9 2 7 14 15 13 14 9 2 16 15 13 9 7 9 2
27 1 15 13 13 2 16 4 13 15 1 10 9 9 2 7 7 13 0 2 16 13 10 9 1 10 9 2
18 14 7 4 13 10 9 0 2 7 13 4 1 0 2 3 0 9 2
6 1 15 15 4 13 2
9 7 3 15 4 13 14 1 11 2
27 1 0 9 15 4 14 13 10 9 2 1 0 9 2 1 11 2 4 15 0 7 0 9 13 0 9 2
11 11 13 1 9 2 1 9 0 0 9 2
6 0 9 13 3 3 2
16 13 10 9 1 11 2 16 4 11 13 13 10 9 1 11 2
15 13 15 3 13 10 0 9 7 9 2 10 9 7 9 2
22 3 13 2 16 13 2 16 13 9 0 2 16 4 9 13 1 10 10 9 7 9 2
4 11 13 0 2
5 3 13 1 11 2
12 15 15 13 1 9 0 2 0 2 14 0 2
14 7 10 9 13 11 3 2 16 16 4 15 3 13 2
5 0 13 0 9 2
21 13 14 0 2 0 9 1 2 0 9 2 0 9 2 16 13 3 1 3 0 2
30 3 7 13 0 9 9 0 2 7 10 9 0 9 15 13 1 9 2 16 4 13 1 10 9 13 10 9 0 9 2
16 7 10 0 9 14 13 3 16 9 9 2 16 15 4 13 2
12 11 4 3 13 11 2 2 10 9 13 9 2
16 2 3 3 15 4 13 14 9 2 13 7 4 15 3 15 2
19 13 4 9 7 13 1 9 0 9 1 0 9 16 14 1 0 0 9 2
21 0 9 2 16 15 13 1 9 16 9 2 9 2 9 9 2 14 13 10 9 2
12 1 11 3 9 4 13 3 3 16 1 11 2
9 11 4 13 3 3 10 0 9 2
21 14 1 11 4 13 9 3 3 2 7 15 15 4 3 16 3 13 13 0 9 2
33 11 7 4 13 0 1 9 10 9 2 1 9 2 16 4 13 1 9 7 0 0 9 2 13 4 0 1 10 0 9 7 9 2
20 0 9 1 9 13 1 9 0 7 3 13 1 9 2 16 13 14 3 0 2
27 16 4 13 0 2 15 14 4 3 13 9 1 9 2 9 1 9 7 0 9 2 7 4 3 13 9 2
16 7 1 9 1 9 13 15 2 16 13 1 3 10 0 9 2
8 11 1 9 12 4 13 0 2
26 16 4 13 0 0 2 4 15 3 13 1 0 9 9 1 9 7 9 2 7 13 1 15 14 11 2
18 7 9 7 9 13 3 0 14 14 3 2 16 15 15 13 10 9 2
14 11 4 13 10 2 9 2 14 3 0 16 11 15 2
13 0 9 1 9 4 13 14 1 9 0 1 0 2
32 13 4 3 3 0 2 3 0 2 1 10 0 9 7 9 7 4 13 0 9 2 1 15 15 4 13 0 0 9 0 9 2
25 15 4 13 13 10 9 2 13 10 9 7 13 10 0 9 1 9 2 16 4 3 14 3 13 2
17 11 13 2 16 9 2 13 14 3 13 14 1 3 0 9 2 2
11 7 13 2 16 4 13 0 0 0 9 2
19 11 4 13 2 16 0 9 14 13 9 2 16 4 15 15 1 15 13 2
18 9 2 9 2 0 9 15 2 15 13 15 3 2 13 14 10 9 2
9 11 13 0 9 2 0 9 2 2
3 0 9 2
24 0 0 9 4 3 2 13 2 1 9 2 7 16 15 4 3 13 2 4 3 13 1 9 2
23 3 4 15 9 13 13 3 15 13 3 2 1 15 7 14 2 13 2 15 14 1 9 2
36 3 3 15 4 13 13 2 7 1 9 1 0 9 4 13 3 0 2 0 9 2 2 1 15 4 1 9 13 14 9 3 0 0 0 9 2
22 0 9 4 13 0 0 9 2 16 15 15 13 14 1 9 12 2 0 9 11 11 2
28 13 4 9 0 9 2 0 9 7 0 9 2 16 9 0 9 9 15 4 4 1 10 9 13 9 0 9 2
13 9 8 11 16 13 14 1 0 9 7 9 9 2
30 15 15 4 3 3 13 1 9 2 16 15 4 14 10 9 3 13 14 11 2 14 16 15 1 11 4 13 0 13 2
17 3 7 15 4 15 13 14 1 9 15 2 3 3 1 0 9 2
28 0 9 13 0 9 2 16 4 13 13 1 9 2 14 16 4 13 3 3 7 1 15 0 1 15 2 2 2
10 10 9 4 13 8 3 3 1 9 2
13 10 9 4 14 13 2 16 16 15 4 13 15 2
13 1 11 7 11 4 0 9 14 13 0 9 9 2
14 13 15 2 16 10 0 9 4 13 13 14 0 9 2
5 11 4 15 13 2
20 16 0 9 1 9 12 4 13 3 13 9 2 16 4 3 13 9 0 9 2
17 14 0 11 4 13 1 9 2 16 4 9 13 1 10 9 9 2
29 15 1 15 4 14 13 2 15 15 13 2 13 4 0 7 0 2 16 4 15 1 9 11 13 0 9 13 11 2
20 1 9 7 10 9 3 4 13 2 16 15 4 13 0 9 2 9 9 2 2
18 1 9 0 9 4 3 1 2 0 11 2 13 3 14 14 9 11 2
26 3 16 4 9 1 0 9 13 11 7 13 0 9 1 0 0 9 2 15 4 9 3 14 3 13 2
5 11 4 13 0 2
18 3 4 13 1 0 9 7 4 13 0 16 13 0 0 9 1 9 2
22 2 15 2 16 13 9 2 2 4 13 10 0 9 2 2 15 3 13 0 1 0 2
31 9 13 0 9 2 9 2 9 2 9 2 0 9 9 2 0 9 2 0 9 2 0 9 7 0 1 0 9 0 9 2
37 3 13 3 0 9 9 2 0 1 0 7 0 9 2 0 0 9 2 1 9 9 2 16 15 16 0 9 13 1 9 2 9 7 0 0 9 2
45 10 9 1 0 9 11 13 1 3 0 9 14 0 9 1 9 11 2 16 4 13 14 1 9 9 2 12 2 1 3 0 9 1 11 2 7 4 13 1 9 12 9 9 9 2
24 1 15 4 0 0 9 12 9 12 13 0 9 1 9 9 7 15 1 15 13 1 0 9 2
6 9 15 13 3 0 2
18 13 7 2 16 15 9 14 13 7 16 13 0 9 1 9 0 9 2
7 3 10 9 14 13 9 2
29 15 3 15 13 1 9 1 9 0 0 9 1 9 9 2 16 15 15 9 3 13 1 15 2 16 15 14 13 2
12 9 1 0 9 15 4 1 10 9 14 13 2
23 11 13 2 16 15 3 13 9 1 9 0 9 2 7 13 9 14 1 0 9 0 9 2
19 0 9 13 3 0 2 7 13 1 0 9 2 1 15 4 15 3 13 2
13 1 0 11 10 9 13 14 1 9 9 7 9 2
12 3 3 0 13 1 9 9 0 9 1 9 2
6 13 7 10 0 9 2
26 11 13 14 12 9 2 1 9 2 16 15 13 0 2 15 14 13 13 9 1 10 16 12 9 9 2
38 13 15 2 3 4 9 13 14 1 9 1 9 9 7 4 3 14 13 0 9 2 4 13 9 11 11 7 13 2 16 4 13 1 0 9 10 9 2
20 9 9 7 10 9 4 13 14 0 0 9 1 9 0 0 9 9 11 11 2
25 0 13 16 0 9 1 0 9 1 9 0 9 12 0 0 9 2 4 13 10 9 8 11 11 2
35 1 0 9 13 1 10 0 9 2 16 15 14 13 1 0 9 7 15 13 2 7 14 3 13 7 3 7 3 0 1 9 1 10 9 2
36 0 13 2 16 0 9 11 2 16 15 4 0 0 9 9 12 13 1 10 9 1 0 9 2 13 9 1 10 9 2 4 13 9 11 11 2
12 14 12 9 9 9 7 9 14 4 13 9 2
25 12 0 13 3 12 9 0 7 0 9 2 1 15 13 12 9 1 9 0 9 7 12 0 9 2
36 0 9 15 13 1 9 9 0 9 1 9 2 4 14 13 7 13 9 11 2 16 14 10 16 12 9 13 0 9 1 0 9 10 0 9 2
32 9 9 8 11 11 2 14 16 1 9 13 9 9 2 1 15 4 14 13 0 9 7 15 9 2 4 13 10 16 1 9 2
8 3 3 0 9 13 0 9 2
18 9 11 11 13 1 10 9 11 3 1 0 0 9 1 9 0 9 2
24 11 2 16 4 13 1 9 14 10 0 11 0 9 2 13 1 10 9 14 10 9 16 0 2
26 10 0 9 2 0 9 11 11 2 0 9 1 11 11 11 7 11 11 2 4 9 3 1 9 13 2
17 0 13 14 9 11 2 16 4 13 13 14 10 9 1 0 9 2
11 0 9 1 12 9 13 14 3 12 9 2
9 13 4 14 9 7 9 1 9 2
14 9 9 13 0 9 2 16 13 13 10 9 1 9 2
11 1 10 9 14 4 13 10 16 12 9 2
15 10 9 1 9 13 0 9 9 2 16 13 1 15 0 2
20 16 15 13 0 2 1 10 9 4 13 10 9 9 2 15 13 9 1 9 2
11 13 1 9 2 15 13 1 9 0 15 2
12 13 10 9 1 9 12 9 9 1 0 9 2
22 14 13 9 2 1 15 13 9 2 7 9 2 16 13 9 2 9 2 9 2 2 2
18 9 1 0 9 1 0 9 15 4 3 13 1 9 2 12 9 12 2
15 1 9 9 0 9 13 0 9 12 9 1 9 10 9 2
12 10 0 9 15 14 13 2 16 15 9 13 2
20 13 1 10 9 2 7 1 9 15 13 9 1 15 15 15 3 13 9 11 2
20 16 15 4 9 1 9 13 0 7 0 2 4 1 9 13 9 1 10 9 2
12 13 15 4 1 15 7 15 1 15 13 3 2
15 16 15 4 13 1 10 9 2 14 0 0 9 13 0 2
21 14 3 14 15 13 2 13 14 10 9 7 14 13 15 0 2 16 15 4 13 2
13 13 13 10 9 1 10 9 7 10 9 1 9 2
19 1 3 0 9 13 9 1 9 3 12 2 12 9 2 16 9 14 13 2
10 3 13 9 7 15 13 9 7 9 2
19 1 9 16 9 3 13 3 0 7 7 15 14 13 2 3 15 13 15 2
18 7 7 15 15 13 14 1 15 2 15 13 0 10 9 1 9 9 2
19 3 15 4 15 13 2 13 0 1 15 2 3 13 0 7 3 13 9 2
17 9 1 0 9 13 9 9 2 13 7 0 2 16 13 3 3 2
23 7 3 3 13 3 2 13 3 0 1 9 0 0 9 2 10 9 7 10 0 0 9 2
26 0 9 9 0 9 1 9 1 11 1 9 0 9 11 13 0 2 7 13 1 12 10 0 0 9 2
28 0 9 1 10 0 9 1 9 13 14 9 1 9 0 11 2 13 3 0 9 0 9 2 7 10 9 2 2
9 13 2 16 4 13 15 12 0 2
9 1 10 9 4 13 14 12 9 2
32 10 9 1 9 9 4 13 14 3 3 7 13 4 15 1 9 2 1 15 4 13 10 9 13 9 1 9 2 0 12 9 2
9 9 4 13 3 2 16 4 13 2
12 11 2 14 13 15 2 3 15 4 15 13 2
21 0 13 2 16 4 13 13 9 2 16 4 13 3 9 2 7 15 4 13 3 2
29 1 15 4 10 9 1 9 2 3 13 9 2 16 4 0 11 3 13 11 2 13 2 16 9 3 13 2 2 2
7 2 9 13 16 0 9 2
2 9 11
8 13 15 2 3 9 13 11 2
15 10 9 13 10 9 2 16 15 3 14 3 14 14 13 2
12 14 0 15 14 13 13 10 9 1 9 11 2
12 2 9 7 1 15 14 13 2 2 13 0 2
15 9 4 3 1 0 9 11 11 13 9 9 7 0 9 2
17 16 4 13 0 2 4 11 1 12 9 13 9 3 12 9 9 2
23 1 15 4 0 9 13 9 10 9 1 0 0 9 7 13 3 13 1 0 9 7 9 2
30 1 10 9 2 15 4 13 0 9 2 4 13 2 16 13 11 2 15 0 9 13 0 9 11 2 10 9 1 15 2
31 0 0 0 9 4 15 13 1 9 11 11 7 0 9 10 0 9 9 1 0 9 0 9 11 11 1 0 9 8 11 2
15 13 4 14 9 11 0 7 9 11 11 7 9 11 11 2
31 3 0 0 9 1 0 0 9 2 0 9 1 12 9 7 12 9 2 13 9 2 9 7 9 9 9 7 9 9 11 2
12 1 9 1 0 9 13 14 0 9 0 9 2
9 1 10 9 15 3 13 10 9 2
6 1 0 7 0 9 2
30 1 15 15 4 13 1 9 9 11 3 3 2 16 4 13 9 9 2 15 9 13 0 9 2 7 4 3 13 0 2
29 15 13 9 2 16 15 13 3 13 1 9 9 9 2 16 3 3 14 13 2 3 4 0 9 14 3 13 0 2
22 2 0 9 2 16 13 1 9 0 7 0 1 9 2 3 14 13 13 0 1 0 2
38 3 1 15 2 16 13 14 9 9 1 9 0 9 0 9 7 9 2 15 3 14 13 2 3 4 9 13 2 16 4 9 13 13 1 0 7 9 2
6 14 13 0 0 9 2
28 9 16 4 0 9 13 0 9 2 16 15 4 13 1 9 1 11 2 15 4 3 13 7 1 3 13 9 2
26 1 9 2 7 9 9 0 1 0 13 14 9 2 16 4 15 10 0 9 13 1 0 9 1 9 2
10 15 7 1 15 15 13 0 1 9 2
30 0 9 1 9 1 9 15 1 9 4 13 2 14 16 4 14 15 13 1 9 2 16 7 9 1 9 14 4 13 2
19 3 4 15 13 1 9 2 16 1 9 14 13 1 9 1 9 1 9 2
28 7 1 12 3 2 16 15 1 0 1 9 13 0 7 0 9 2 4 13 1 0 7 0 9 13 0 9 2
12 15 9 13 1 9 2 0 4 1 15 13 2
19 3 4 13 2 16 14 13 9 2 15 13 3 1 15 2 7 14 13 2
11 13 2 16 4 14 9 15 13 1 15 2
6 7 9 13 15 13 2
14 16 13 9 1 15 0 2 15 13 13 14 1 15 2
25 2 10 0 9 1 0 9 2 16 4 1 0 9 1 9 13 1 9 2 4 13 13 3 0 2
11 2 14 14 4 13 2 15 13 1 15 2
9 14 13 2 15 0 4 15 13 2
15 2 10 9 7 4 14 13 2 1 10 9 15 4 13 2
22 0 4 1 0 3 13 0 9 2 1 15 13 9 2 16 4 13 0 9 2 0 2
18 2 7 10 9 2 16 13 0 12 2 12 2 15 4 14 3 13 2
34 1 0 7 13 3 9 2 2 15 4 13 12 1 9 2 16 13 14 10 9 2 16 13 0 1 9 7 15 9 13 14 1 9 2
7 9 9 0 9 13 9 2
18 1 15 13 0 9 14 0 9 9 2 1 9 1 9 7 1 15 2
15 7 14 9 13 0 2 7 0 11 13 14 3 12 9 2
26 1 9 1 0 9 9 4 11 14 11 13 1 0 0 9 1 0 9 2 16 13 0 0 9 9 2
14 10 10 9 15 3 13 1 9 2 16 13 3 13 2
18 11 13 10 9 2 16 13 1 9 9 0 9 1 9 2 0 9 2
26 1 9 9 7 0 9 1 9 9 4 11 13 1 9 2 16 4 3 14 10 9 13 9 1 9 2
9 7 9 0 9 1 9 13 0 2
23 3 0 9 2 16 15 13 7 9 0 9 16 0 9 1 0 9 2 10 9 13 3 2
9 0 0 9 13 1 9 14 3 2
17 9 13 2 3 9 4 11 14 3 1 0 9 11 13 10 9 2
11 0 9 0 9 13 14 14 0 0 9 2
21 3 3 0 4 13 0 0 9 2 7 14 11 0 14 4 13 13 9 9 9 2
12 1 15 13 3 10 9 0 14 1 0 9 2
17 11 11 4 1 0 0 9 0 9 9 12 13 1 9 11 12 2
20 13 1 9 11 1 9 12 9 1 9 2 16 13 1 12 9 8 1 9 2
9 9 13 1 9 1 0 9 9 2
19 13 15 3 1 9 9 2 1 9 0 9 7 13 1 9 14 0 9 2
6 0 9 13 9 9 2
21 0 13 10 9 2 1 0 13 13 9 2 11 2 9 2 9 2 9 7 9 2
15 16 13 0 9 0 1 9 2 13 15 0 14 0 9 2
13 9 3 14 13 0 9 2 1 15 13 0 9 2
17 3 13 9 1 15 9 2 9 7 13 9 7 9 1 0 9 2
13 9 13 3 12 0 9 9 7 15 13 10 9 2
6 9 13 3 3 3 2
21 9 4 10 9 13 9 0 9 1 11 2 13 4 9 7 9 9 9 1 9 2
11 0 13 9 9 1 0 9 7 0 9 2
6 3 14 9 13 15 2
19 15 13 2 16 13 9 0 7 0 2 15 13 14 1 0 2 0 9 2
9 14 0 9 13 3 0 7 0 2
13 1 0 9 13 3 0 9 1 9 7 9 15 2
18 15 13 2 16 15 13 9 3 13 2 15 9 4 1 9 9 13 2
17 16 13 1 0 7 0 9 7 0 9 2 9 14 13 0 9 2
16 3 15 9 3 3 13 2 16 13 1 9 0 10 0 9 2
14 16 13 2 13 0 0 9 3 15 2 15 13 9 2
30 0 13 2 16 1 9 14 13 2 15 10 9 13 2 3 15 4 3 13 2 16 4 9 7 15 1 10 9 13 2
35 14 1 9 7 3 4 13 2 16 13 9 1 9 1 12 9 7 9 2 13 14 1 9 9 11 7 9 11 2 1 3 12 9 9 2
16 15 13 10 9 2 16 13 14 1 9 0 9 1 0 9 2
7 7 9 9 13 3 0 2
9 1 9 9 13 15 0 0 9 2
17 15 7 13 13 3 0 0 9 2 16 13 1 10 9 0 9 2
21 0 9 13 7 0 1 9 9 7 14 9 9 2 16 13 9 1 9 9 9 2
14 14 16 13 0 9 2 13 9 9 2 7 15 13 2
9 13 14 9 2 16 13 9 0 2
12 16 13 0 2 13 0 13 2 16 13 9 2
26 9 0 9 15 4 1 0 9 13 2 16 13 0 9 0 0 9 7 10 9 1 11 15 0 9 2
33 16 13 1 15 12 9 1 12 9 9 0 9 1 3 14 0 9 0 9 2 13 1 15 3 1 10 9 3 1 9 1 9 2
26 9 13 9 9 2 16 4 15 1 11 13 1 0 9 1 9 0 9 12 1 0 9 12 2 12 2
17 10 0 9 4 13 0 9 2 16 4 1 11 1 11 13 9 2
9 14 10 9 4 13 0 0 9 2
24 11 11 4 3 13 2 16 4 10 9 13 1 9 2 16 4 13 14 3 0 1 9 9 2
30 9 9 4 1 0 13 14 9 0 0 9 11 11 2 16 4 13 2 16 13 11 13 0 9 2 0 1 0 9 2
24 16 4 15 11 3 13 1 10 9 2 15 14 3 14 4 13 3 2 7 4 9 3 13 2
16 1 9 13 12 3 0 2 1 9 7 15 10 9 14 13 2
34 0 0 9 13 2 16 13 1 9 0 9 7 16 13 0 9 1 0 9 1 10 9 2 13 11 2 16 13 1 9 14 0 9 2
8 3 4 13 12 9 9 9 2
16 9 9 13 2 9 2 2 16 15 13 9 2 9 7 9 2
8 3 12 9 10 9 13 9 2
26 9 1 9 2 9 7 9 4 13 9 1 9 0 9 9 9 1 9 9 9 7 9 7 9 9 2
38 9 9 2 0 9 7 0 0 9 2 4 9 9 2 1 15 4 13 13 10 9 9 9 7 15 13 0 9 9 2 1 0 9 13 1 0 9 2
16 9 4 13 0 12 9 9 2 9 9 4 13 9 1 9 2
14 1 15 4 9 7 9 13 9 2 9 7 0 9 2
16 1 12 9 3 4 3 13 0 0 7 0 9 1 0 9 2
14 1 0 9 11 7 9 9 9 12 7 4 3 13 2
6 10 9 14 13 9 2
30 9 9 9 7 13 2 16 4 13 9 1 9 1 9 0 3 2 16 4 1 10 11 13 10 9 2 14 3 2 2
25 7 4 9 9 13 3 0 0 9 2 1 15 14 4 0 9 9 1 12 9 13 1 0 9 2
19 0 13 2 16 10 9 1 10 9 13 3 2 3 7 15 13 1 0 2
21 0 13 14 2 16 13 0 9 10 2 3 2 9 2 16 13 0 1 12 9 2
26 16 4 10 10 9 13 2 4 13 1 9 2 0 9 1 9 2 9 1 0 9 2 13 9 11 2
4 15 15 13 2
11 15 13 1 10 9 16 3 3 0 11 2
21 1 0 0 7 0 9 11 13 14 9 2 0 1 11 2 15 15 13 1 9 2
14 15 4 13 3 3 1 0 9 2 16 4 15 13 2
25 1 0 9 9 13 0 9 9 7 9 2 16 1 0 9 1 0 9 13 9 9 2 9 2 2
12 3 13 0 1 11 11 12 7 13 11 12 2
6 9 13 0 9 9 2
22 9 4 7 13 1 9 1 9 11 1 12 9 2 0 4 13 1 12 9 11 9 2
28 1 0 9 9 7 0 0 9 4 13 9 3 0 2 16 1 9 9 7 9 9 9 7 9 9 14 13 2
25 9 1 11 12 13 3 3 0 2 16 1 15 4 13 3 3 0 16 1 15 9 11 7 11 2
33 10 0 9 2 16 13 14 0 9 2 15 13 1 0 9 1 9 9 2 10 0 9 7 13 10 9 7 15 13 1 9 9 2
20 1 15 3 13 0 9 7 2 7 9 9 2 13 7 3 14 0 9 9 2
13 10 9 1 10 9 14 0 13 9 0 9 11 2
22 0 9 1 9 0 9 13 15 9 2 16 4 13 0 9 9 1 0 9 7 3 2
10 1 3 0 9 4 14 13 3 9 2
26 1 15 3 4 3 13 14 15 2 16 4 0 9 13 9 1 9 2 7 16 4 10 9 13 9 2
32 11 4 1 9 13 0 12 2 0 9 11 2 16 4 13 9 0 9 11 9 12 9 1 9 1 10 16 12 9 1 9 2
12 9 12 13 0 0 9 1 3 12 0 9 2
17 0 14 4 13 1 9 0 9 2 16 13 0 1 0 0 9 2
16 1 10 9 13 9 9 0 9 2 0 1 9 9 2 9 2
28 1 15 1 9 13 3 13 1 10 0 9 2 16 13 0 1 9 0 9 7 13 0 0 9 1 9 9 2
37 16 7 13 1 9 14 0 9 9 2 9 1 0 0 9 2 13 3 0 2 16 13 1 10 0 9 7 1 14 3 10 0 9 16 9 9 2
31 1 10 9 13 3 13 0 9 0 9 7 9 9 0 9 1 0 9 0 9 7 0 9 9 2 16 15 13 1 9 2
22 3 13 3 13 9 0 9 1 9 2 16 14 4 3 13 9 9 0 0 0 9 2
12 13 4 15 9 2 13 9 1 9 7 13 9
29 11 11 2 12 2 16 15 4 1 0 13 1 11 11 2 13 3 1 15 9 9 14 3 2 16 13 3 0 2
12 11 15 4 1 9 11 11 14 13 1 15 2
6 6 2 15 13 11 2
3 13 0 2
9 7 13 0 9 2 15 4 13 2
23 16 4 13 10 9 1 9 2 11 11 7 11 11 2 4 13 14 0 11 11 2 11 2
10 0 15 4 13 1 9 2 3 13 2
5 11 2 3 13 2
15 7 11 4 13 0 2 16 15 4 13 2 14 3 13 2
6 3 4 13 1 3 2
9 9 12 4 13 1 11 0 9 2
14 13 15 15 4 7 15 16 0 11 13 1 0 9 2
14 13 7 4 0 9 1 9 2 7 4 13 3 3 2
11 10 9 4 13 14 1 12 2 12 9 2
20 9 4 3 1 15 1 0 3 13 2 7 1 12 2 12 9 4 3 13 2
19 1 15 15 4 3 13 1 0 9 0 9 2 16 15 4 13 9 9 2
7 13 4 0 9 1 11 2
17 14 1 9 15 4 13 2 7 9 9 4 3 13 1 0 9 2
7 10 9 4 13 9 12 2
13 15 13 0 9 9 2 3 7 13 14 12 9 2
21 3 1 3 1 9 13 1 9 0 9 11 2 11 2 16 13 9 0 9 9 2
4 3 13 0 2
10 16 4 14 13 2 4 15 3 13 2
20 13 0 1 9 2 7 1 0 9 4 0 9 13 3 2 16 13 10 9 2
16 15 13 13 3 0 2 13 1 9 15 1 9 2 7 13 2
20 0 9 4 9 11 3 13 2 7 4 3 13 2 3 4 15 13 10 9 2
26 13 15 4 1 9 8 8 11 2 16 4 13 14 10 9 2 7 15 4 13 13 14 9 11 11 2
15 4 14 3 15 13 1 9 7 13 10 0 9 1 9 2
9 9 8 8 11 15 1 9 13 2
40 9 1 9 0 7 0 0 9 11 11 4 15 1 0 9 3 13 1 9 2 16 13 9 2 1 15 13 0 9 2 9 7 0 9 1 0 9 1 0 2
25 16 13 3 11 1 9 2 16 4 3 13 2 16 15 4 13 13 0 9 2 13 10 9 0 2
25 1 0 12 9 9 4 13 11 8 11 2 15 12 9 13 3 2 15 10 9 7 3 3 9 2
37 1 9 10 12 12 9 2 1 15 4 13 0 10 9 2 9 7 9 2 13 2 16 15 3 3 13 9 2 16 4 15 3 13 0 7 0 2
33 10 0 9 13 1 9 1 10 11 3 0 2 13 4 14 15 12 9 1 15 12 2 16 15 4 4 1 15 9 13 7 13 2
12 9 2 0 9 2 13 2 7 15 13 9 2
15 16 13 9 0 2 9 13 1 9 7 15 13 1 9 2
15 13 15 3 2 16 15 1 10 9 13 1 9 7 13 2
42 1 9 2 16 4 13 7 13 9 0 0 0 9 1 10 11 1 9 9 2 16 13 14 14 0 9 2 9 7 0 9 2 13 1 9 10 3 0 9 0 9 2
13 11 11 15 14 13 1 0 9 7 3 13 9 2
22 1 9 9 15 4 3 13 14 10 9 2 1 15 13 10 9 2 7 14 13 9 2
17 13 1 0 9 2 16 13 1 9 2 12 13 3 0 9 2 2
7 12 0 13 9 12 9 2
16 0 9 9 13 0 9 2 0 9 9 7 9 9 13 0 2
13 16 4 13 0 9 9 2 15 13 1 9 3 2
10 15 13 0 1 9 0 9 7 9 2
25 9 1 9 13 9 1 0 9 2 0 9 2 0 0 0 9 7 9 1 9 9 1 0 9 2
24 3 13 15 1 0 9 2 0 9 7 0 9 2 7 13 9 1 9 1 10 9 14 13 2
8 9 11 13 16 10 0 9 2
4 1 9 3 13
12 9 9 3 13 14 16 9 1 9 0 9 2
22 1 9 9 9 3 13 9 2 16 3 3 13 1 10 9 8 13 10 9 1 9 2
21 10 9 13 1 9 1 9 9 1 9 0 9 7 1 9 0 9 2 16 13 2
16 9 13 1 9 0 9 7 1 9 0 9 2 1 15 13 2
22 9 9 13 9 7 1 9 13 9 12 2 0 9 2 16 4 13 0 1 0 9 2
17 3 13 14 0 2 16 1 0 9 0 9 14 13 10 9 14 2
9 3 13 0 2 3 3 0 9 2
15 13 1 9 0 0 9 2 16 13 3 3 0 3 3 2
15 9 7 1 0 9 13 14 9 0 9 2 16 15 13 2
20 9 11 8 11 11 4 9 1 9 1 0 9 13 0 0 9 9 9 11 2
38 1 0 0 9 7 0 9 1 0 0 9 4 9 11 11 13 14 9 11 11 11 2 11 11 2 11 11 2 11 11 11 2 11 11 7 11 11 2
