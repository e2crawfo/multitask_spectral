322 11
5 3 13 9 1 2
21 9 13 3 1 9 7 9 2 15 15 4 13 3 1 10 9 1 10 13 9 2
12 11 9 4 13 12 9 2 2 13 11 11 2
21 11 13 1 9 7 13 10 0 0 9 2 1 15 3 3 4 13 15 13 1 2
9 11 11 4 10 0 7 0 9 2
38 7 3 4 15 3 1 0 9 4 13 10 0 9 7 10 10 9 1 9 1 15 2 15 4 13 1 11 9 2 7 1 9 13 13 15 0 9 2
13 9 13 15 0 1 10 9 1 15 15 13 15 2
6 15 13 3 1 15 2
7 9 3 13 3 0 9 2
9 2 15 13 15 10 9 1 9 2
18 2 11 11 11 4 3 0 2 16 10 9 4 4 13 1 0 9 2
29 15 4 3 0 1 10 9 1 9 9 2 7 3 4 9 3 1 10 0 4 13 1 9 7 13 9 1 9 2
31 13 15 0 0 9 2 4 15 13 10 9 1 9 1 9 9 7 9 9 2 16 0 9 3 13 0 9 7 13 9 2
33 9 11 7 9 11 2 15 1 10 9 13 3 1 11 2 3 15 4 13 1 9 1 10 9 9 11 2 13 3 3 1 9 2
27 6 1 11 1 15 13 13 10 0 9 2 7 6 1 11 2 15 13 10 9 2 7 3 13 10 9 2
5 2 13 3 3 2
15 2 15 4 13 10 9 1 0 10 9 2 15 4 13 2
9 15 4 4 13 1 9 1 15 2
8 2 15 4 15 2 15 13 2
10 1 10 9 2 9 4 0 1 9 2
28 14 4 10 0 4 0 2 11 1 8 8 2 7 14 4 0 9 4 3 15 1 10 0 2 15 4 13 2
30 0 2 15 4 3 13 13 10 9 1 10 9 2 7 16 15 10 9 13 10 9 2 3 4 15 4 13 15 3 2
27 9 4 13 2 16 10 9 2 2 3 9 2 15 13 3 2 2 3 13 2 16 15 3 13 0 9 2
16 15 13 9 3 7 13 1 9 7 3 14 13 9 1 9 2
35 7 3 16 10 9 4 13 1 9 9 2 4 15 3 13 10 9 1 15 2 15 13 10 13 9 1 10 0 9 1 14 13 1 9 2
4 11 11 13 2
4 2 9 9 2
25 13 15 3 1 11 2 1 10 13 9 1 9 2 4 15 3 3 13 15 1 9 1 0 9 2
19 10 9 1 10 9 2 3 4 4 0 1 9 2 7 1 9 0 9 2
3 2 3 2
58 3 13 10 9 1 9 9 1 14 13 9 2 3 1 0 7 0 9 2 16 15 3 4 9 7 9 13 10 9 2 3 3 16 3 4 13 9 1 9 2 7 3 9 2 15 13 9 2 13 2 4 9 3 13 15 0 9 2
21 0 0 13 1 9 14 13 9 1 14 2 13 9 7 9 0 1 15 13 2 2
1 9
34 10 9 3 13 2 16 10 9 3 1 0 9 13 9 1 9 2 7 10 9 2 15 3 3 3 4 13 1 14 13 9 1 9 2
27 9 1 11 4 3 3 4 13 2 16 9 4 13 9 2 7 15 13 3 9 1 9 1 14 13 9 2
33 15 4 13 1 9 2 7 15 4 3 13 15 3 7 13 1 14 13 3 1 10 9 2 15 4 13 3 3 1 9 1 11 2
8 7 15 4 3 3 13 15 2
11 3 10 9 1 10 9 4 13 1 9 2
13 9 2 9 7 9 1 11 13 3 10 0 9 2
17 2 3 13 15 9 2 15 4 3 0 14 4 9 1 10 9 2
16 1 0 9 13 1 15 9 2 9 7 9 2 9 7 9 2
19 7 1 2 16 9 4 13 1 0 9 2 3 4 15 3 0 1 11 2
4 1 9 1 11
9 7 15 13 15 1 9 14 13 2
14 2 15 4 3 0 2 16 9 13 12 9 1 9 2
35 3 4 15 3 3 9 2 7 15 13 3 2 15 15 13 3 1 15 2 16 15 13 0 9 1 0 2 7 1 9 4 15 0 9 2
19 15 13 3 9 1 14 13 15 1 9 2 7 15 13 3 10 9 1 2
24 15 13 9 1 10 3 0 7 0 9 2 7 1 10 9 13 15 3 7 13 15 10 9 2
5 11 4 13 1 11
37 7 3 15 3 3 13 11 11 2 11 11 2 11 2 13 15 3 2 15 15 13 9 1 1 9 2 2 13 11 11 2 9 1 9 9 11 2
20 9 4 13 9 9 2 7 3 13 9 1 9 9 7 9 7 1 9 9 2
39 15 4 9 1 9 1 9 1 9 7 1 9 2 7 3 1 9 13 15 0 15 2 15 1 9 13 1 10 0 9 13 1 15 1 10 0 0 9 2
16 15 13 15 15 2 16 11 9 3 4 4 13 1 10 9 2
28 10 12 9 13 1 9 13 11 0 9 2 11 1 9 7 10 0 9 1 9 1 10 0 2 11 11 2 2
7 2 3 4 15 13 9 2
42 10 0 9 1 9 13 11 11 1 9 1 10 0 11 11 2 15 3 4 4 13 1 9 1 12 9 2 7 13 3 1 10 0 9 2 15 13 1 10 0 9 2
24 16 15 1 9 4 13 2 16 2 15 15 4 3 3 0 2 2 4 15 3 4 13 15 2
34 7 11 13 9 3 7 15 4 13 2 16 15 4 15 1 9 1 10 0 9 2 15 0 9 9 13 1 9 1 9 1 9 12 2
26 16 15 1 9 13 13 9 1 10 0 9 2 13 15 3 10 9 1 9 3 1 9 1 0 9 2
10 2 10 0 0 9 2 13 15 13 2
7 15 4 13 15 2 9 2
19 7 0 13 2 16 15 13 1 9 2 16 10 0 9 3 4 13 3 2
10 3 4 15 13 1 10 9 3 2 2
3 11 0 9
23 15 4 13 15 15 14 13 2 7 15 4 3 0 2 16 15 3 13 1 10 9 2 2
16 10 0 9 1 9 13 15 3 2 15 4 13 15 1 14 13
26 15 4 3 3 9 2 1 12 9 4 15 13 0 9 1 9 7 3 1 10 9 2 3 1 9 2
11 7 1 10 0 12 9 4 15 13 3 2
21 1 3 4 15 1 11 13 15 1 10 0 9 2 16 9 4 0 1 10 9 2
2 0 9
24 9 3 13 15 9 1 2 0 9 2 2 7 1 12 13 15 10 0 9 2 2 9 2 2
10 9 1 9 13 14 13 12 9 9 2
8 9 1 9 13 3 1 9 2
13 2 1 9 13 3 9 9 7 13 3 1 9 2
20 16 15 13 3 1 11 2 4 3 13 10 9 9 2 7 15 4 3 9 2
18 4 15 15 2 16 9 3 4 0 2 3 4 15 3 13 1 15 2
2 4 9
29 0 11 11 2 15 13 1 10 3 0 9 7 9 1 9 1 10 0 2 13 9 13 3 1 9 1 10 9 2
18 9 4 3 3 2 15 13 3 1 9 1 10 13 9 1 10 9 2
17 15 4 13 11 0 0 9 7 3 13 10 0 9 1 0 9 2
32 10 9 13 13 7 13 3 2 15 4 11 2 15 13 9 7 9 1 15 7 4 3 14 13 2 16 15 1 15 4 13 2
2 0 9
8 10 0 13 3 1 9 12 2
11 13 9 3 1 9 2 7 3 1 9 2
19 2 15 4 3 13 11 3 0 2 15 13 10 9 1 9 3 1 9 2
29 15 4 3 3 13 2 16 9 9 2 11 11 2 3 13 1 11 9 1 9 1 3 11 11 11 1 11 11 2
10 2 15 13 3 10 1 9 1 9 2
17 16 15 13 10 9 1 9 1 14 13 9 1 9 1 9 2 2
10 11 13 15 1 2 16 9 4 0 2
31 15 13 15 2 16 10 9 13 14 13 2 16 0 11 2 15 15 13 1 10 0 9 0 9 2 4 4 13 1 15 2
22 9 4 3 13 3 10 0 9 2 7 10 0 9 13 3 3 1 11 1 0 9 2
8 11 13 12 9 3 1 10 9
52 9 2 9 8 11 11 11 2 15 15 4 13 10 0 9 1 14 13 9 7 9 1 9 2 3 9 2 13 3 3 2 16 2 9 2 15 13 10 0 9 2 4 13 15 1 2 16 10 9 4 13 2
38 7 10 0 9 13 1 2 16 15 15 4 13 1 10 0 9 2 10 0 7 3 0 11 11 2 1 11 11 1 10 9 9 1 3 4 0 1 2
34 7 0 13 3 2 16 16 11 13 10 9 1 12 9 1 12 9 2 3 4 15 1 0 9 9 15 2 15 13 1 10 0 9 2
18 1 9 1 14 13 13 15 3 1 9 7 13 1 9 1 10 9 2
13 2 6 2 2 13 15 7 13 15 3 1 9 2
24 11 11 7 11 11 4 9 2 7 11 11 11 7 11 11 4 4 9 1 0 1 12 9 2
21 11 11 11 13 1 10 0 9 2 15 4 13 1 3 14 4 13 15 1 11 2
59 2 16 3 12 9 1 9 3 13 9 2 7 9 9 1 0 9 13 9 1 9 2 3 4 10 0 9 4 0 1 2 16 3 13 3 9 1 10 9 2 2 13 11 11 7 13 1 9 1 9 7 13 9 1 0 0 0 9 2
24 16 10 9 4 13 2 13 9 1 10 9 1 11 12 9 1 9 1 9 1 9 7 9 2
26 15 13 15 1 11 11 11 0 9 1 11 2 3 11 13 9 11 11 2 15 4 13 9 1 9 2
15 7 15 13 11 1 10 0 7 0 11 8 12 1 12 2
23 4 15 4 9 12 9 2 3 13 13 2 3 3 1 15 3 3 13 2 15 4 13 2
28 9 7 9 13 15 3 14 4 10 13 9 2 7 10 9 13 15 1 14 13 9 1 9 1 10 0 9 2
30 2 7 3 13 15 3 10 9 2 2 13 11 11 2 15 3 13 2 16 15 3 4 4 3 7 2 13 2 9 2
7 0 9 13 3 0 9 2
48 2 13 3 1 9 10 0 9 1 2 16 15 4 4 10 9 2 16 10 9 4 0 7 0 1 9 2 13 15 2 15 4 4 0 14 13 2 16 15 3 13 10 0 7 10 0 9 2
12 15 4 15 3 3 3 13 14 13 15 1 2
15 8 11 13 10 0 9 1 15 7 13 15 3 1 9 2
4 12 0 9 2
23 10 9 9 2 15 9 4 13 1 9 11 2 4 3 1 9 3 13 1 9 7 9 2
17 3 4 15 13 0 9 1 9 2 7 13 0 9 1 0 9 2
22 15 13 1 10 9 3 1 10 0 9 2 3 9 13 2 16 15 4 13 1 9 2
13 9 1 10 0 9 13 3 1 9 1 11 9 2
17 1 9 4 11 11 13 3 2 7 3 1 11 11 4 3 11 2
26 11 13 3 3 3 9 1 2 16 9 1 9 0 9 7 3 1 9 1 9 4 4 3 3 0 2
17 2 10 9 1 2 15 9 13 3 1 2 13 1 10 10 9 2
23 1 10 9 13 10 0 9 2 15 3 13 1 9 1 9 7 3 13 0 7 0 9 2
24 2 15 4 9 2 15 13 1 14 13 1 9 2 7 10 0 15 3 13 2 15 4 13 2
18 10 10 9 2 9 2 4 13 1 11 9 7 3 1 9 1 11 2
13 7 15 13 15 3 13 2 3 0 10 9 13 2
23 11 11 13 3 3 9 1 9 2 7 15 4 15 3 13 15 14 13 10 0 9 1 2
10 10 9 4 13 1 11 0 9 9 2
15 3 4 3 3 3 13 9 1 11 2 10 9 4 13 2
19 15 4 3 9 2 16 11 4 13 10 3 3 0 9 14 4 4 13 2
27 15 4 13 10 0 9 1 9 2 15 13 3 1 2 16 10 0 9 1 0 9 13 1 9 1 9 2
24 7 15 4 15 13 15 1 14 13 2 13 10 0 11 2 15 3 13 14 4 9 1 10 9
14 15 3 4 13 3 1 9 2 4 3 4 10 9 2
10 3 3 13 15 3 7 13 15 13 2
27 9 1 11 11 13 13 7 13 1 10 0 9 2 15 3 13 1 9 0 2 0 9 7 9 1 9 2
73 9 11 11 2 15 4 13 9 2 9 9 2 7 3 13 1 11 2 13 13 1 2 3 0 9 3 13 3 2 2 13 15 1 9 2 16 10 0 9 13 15 1 14 4 10 9 2 3 0 0 9 4 1 9 2 3 13 15 9 1 9 1 9 1 9 1 10 3 0 9 1 11 2
20 2 15 13 1 10 9 7 13 10 9 1 10 9 2 16 15 13 9 13 2
3 2 6 2
7 15 4 0 9 3 2 2
13 9 0 9 13 1 9 9 1 14 13 1 9 2
14 13 3 3 7 3 3 1 10 3 0 9 7 9 2
20 9 4 13 12 9 2 7 15 4 0 2 16 9 13 3 0 9 7 9 2
26 9 1 0 9 4 9 2 7 10 9 1 9 13 3 0 9 1 10 13 9 2 3 3 3 9 2
29 3 13 9 10 0 9 3 3 1 3 1 10 0 9 1 10 0 9 7 1 10 0 9 1 10 3 13 9 2
16 9 1 9 2 10 9 7 9 9 2 4 3 0 7 0 2
15 0 1 9 4 15 13 3 10 9 1 12 9 7 12 2
20 9 4 3 4 13 2 7 3 13 0 9 1 2 16 11 11 13 15 3 2
15 15 13 1 15 2 16 10 9 1 15 4 0 1 9 2
14 15 13 15 3 1 10 0 9 7 13 3 1 9 2
36 13 9 1 9 3 2 16 10 9 7 9 4 13 1 9 2 7 16 10 9 7 9 4 4 13 1 9 2 13 9 10 9 1 10 9 2
26 2 6 2 3 13 15 7 13 2 7 11 13 3 13 2 16 15 13 10 9 9 3 2 13 11 2
23 11 4 13 9 11 11 1 10 13 9 2 7 15 13 3 14 13 9 7 13 1 9 2
22 16 0 9 4 0 7 0 1 9 2 15 13 3 10 9 1 2 13 11 11 11 2
51 15 4 15 2 15 13 3 1 14 2 13 2 9 2 7 1 11 11 1 9 13 9 14 13 9 1 10 9 2 10 9 15 3 4 0 1 1 9 2 3 15 13 14 13 9 7 9 1 0 9 2
16 11 11 13 2 1 0 10 0 9 2 10 0 9 1 9 2
14 0 9 4 13 1 9 2 9 7 9 7 1 9 2
10 9 4 3 13 1 10 0 9 2 2
9 11 11 2 0 9 1 11 11 2
16 9 4 2 9 2 2 7 9 4 13 1 11 11 2 11 2
14 9 13 2 16 15 13 12 9 1 15 13 12 9 2
11 9 13 1 9 2 15 4 13 1 9 2
27 4 3 10 0 9 7 11 9 9 10 9 13 3 1 9 2 16 15 13 15 1 9 1 10 0 9 2
15 7 15 4 3 3 13 15 1 0 9 14 13 1 15 2
16 9 4 13 14 13 9 1 11 7 11 7 13 3 3 12 8
18 15 4 13 2 16 10 0 4 13 1 9 7 13 1 9 3 3 2
42 0 13 3 1 2 9 2 1 9 2 7 1 10 9 2 15 3 4 1 9 1 9 0 9 2 4 11 11 3 3 7 3 13 10 11 1 3 0 9 1 0 11
21 3 13 15 1 9 2 15 13 2 16 11 3 4 13 0 9 1 11 1 11 2
38 2 15 13 1 9 2 7 16 15 13 3 2 4 10 0 3 0 2 7 15 13 0 9 3 3 1 9 1 0 9 2 2 13 11 11 1 11 2
1 2
24 2 16 15 4 13 14 13 10 0 9 2 11 11 2 2 13 15 3 1 10 3 0 9 2
8 11 4 3 13 1 10 9 2
19 15 13 2 3 1 3 3 13 10 9 2 15 3 4 3 1 7 13 2
8 15 4 3 13 10 9 9 2
20 15 13 8 9 1 15 2 7 15 13 3 1 2 16 15 4 13 1 9 2
7 7 4 15 3 3 15 2
19 15 13 3 2 16 15 13 1 14 13 15 2 7 16 15 3 4 0 2
9 10 9 13 3 1 3 10 0 2
21 1 9 1 9 9 4 15 4 13 9 9 1 8 15 15 1 0 9 1 9 2
34 1 9 13 3 0 12 9 2 15 3 3 4 13 3 1 9 7 3 1 0 9 3 13 1 9 2 1 9 7 9 1 9 9 2
14 1 9 9 4 15 13 9 2 15 13 9 1 9 2
32 15 13 15 3 3 1 15 2 7 1 10 0 9 4 15 13 0 9 1 14 13 1 9 1 10 10 9 2 2 13 15 2
20 10 0 9 4 9 2 16 10 0 9 4 9 2 7 15 13 3 1 15 2
36 15 13 13 2 16 15 1 9 1 10 1 0 9 0 9 1 14 13 10 0 9 1 11 2 13 3 3 13 3 1 3 10 9 1 11 2
18 12 9 9 7 9 1 9 13 3 2 16 9 4 13 1 12 9 2
37 15 4 0 3 2 16 10 0 13 9 1 9 9 2 7 3 1 9 4 10 0 9 13 14 13 9 1 0 9 9 2 7 15 4 0 9 2
8 0 9 13 3 1 0 9 2
27 7 3 9 1 2 1 15 9 9 4 13 3 4 13 1 13 1 9 2 13 9 3 14 13 1 9 2
12 3 13 10 0 9 1 10 0 9 1 9 2
7 15 4 10 0 0 9 2
19 11 2 6 2 6 2 3 2 6 2 7 15 4 0 2 13 15 2 2
28 10 9 7 15 4 13 2 16 15 4 13 1 11 1 10 12 9 2 16 15 4 13 9 14 13 9 9 2
13 15 13 3 0 2 3 15 4 13 10 0 9 2
9 2 15 13 14 13 1 0 9 2
8 10 0 9 13 10 0 9 2
6 3 13 15 9 2 2
30 10 0 9 1 3 10 0 9 1 14 13 9 7 9 3 1 10 3 13 9 2 4 13 9 2 2 13 11 11 2
26 9 13 1 9 3 9 12 1 14 13 0 1 9 12 2 13 15 1 9 2 9 11 11 2 11 2
36 7 3 1 9 4 15 3 0 1 2 16 10 0 9 9 4 13 10 0 9 1 9 9 2 3 1 0 9 2 16 9 13 1 9 3 2
11 2 13 15 2 13 10 9 1 10 9 2
3 2 3 2
8 9 13 10 9 1 0 9 2
17 15 13 10 9 3 1 10 0 9 2 16 9 11 11 13 9 2
2 11 9
1 2
20 15 4 3 10 9 16 15 1 9 1 11 13 14 13 9 1 4 3 0 2
9 11 13 15 1 15 1 10 9 2
9 7 13 10 9 1 12 9 9 2
19 15 13 10 9 1 2 16 15 1 11 4 13 10 9 1 10 9 9 2
32 7 15 4 13 0 9 2 15 15 1 15 4 13 13 9 1 10 9 1 10 9 2 15 4 13 2 7 3 1 15 0 2
22 3 1 12 9 1 11 9 4 15 13 2 15 3 13 9 10 0 9 2 7 3 2
10 15 4 3 1 14 13 9 1 15 2
8 9 13 3 3 10 0 9 2
10 11 11 9 1 10 0 9 4 0 2
5 15 4 3 0 2
20 10 0 9 1 11 4 3 13 1 10 0 9 2 7 3 13 11 3 3 2
43 9 13 9 12 1 9 1 12 8 2 7 15 4 13 2 16 15 4 13 1 12 9 2 7 1 9 1 10 0 9 4 9 1 12 2 16 15 13 1 9 1 9 2
18 1 9 2 3 4 10 0 9 3 3 13 9 1 10 0 2 9 2
33 3 4 15 13 10 9 2 11 11 2 1 14 13 15 1 9 2 2 13 11 11 2 15 13 0 1 14 13 15 3 1 11 2
17 10 9 13 3 1 10 0 1 11 2 16 11 9 4 3 0 2
10 10 13 0 9 13 15 1 9 9 2
19 15 13 10 9 1 9 3 1 9 1 14 13 15 9 1 14 13 3 2
6 13 9 2 11 9 2
29 1 0 9 9 4 9 13 2 16 10 3 12 9 3 4 13 3 2 13 9 7 9 3 7 13 1 0 9 2
15 15 4 15 13 1 0 9 2 3 0 1 9 1 9 2
19 10 9 13 1 10 9 3 1 9 9 11 2 11 2 11 7 11 11 2
16 15 4 3 4 13 1 10 0 9 2 2 13 9 11 11 2
8 7 1 10 9 13 0 9 2
33 9 1 9 1 9 1 9 7 10 9 2 15 13 1 9 1 9 2 4 4 13 1 12 9 1 2 16 9 7 9 4 13 2
50 1 0 11 3 3 1 13 2 7 11 1 0 9 2 4 15 4 3 0 1 14 13 10 0 9 2 3 3 1 9 1 11 1 11 2 3 15 3 13 10 2 0 2 9 16 15 13 1 9 2
15 9 12 13 12 10 9 1 10 0 9 9 2 11 11 2
26 11 11 11 13 3 1 9 2 16 11 11 2 11 2 7 9 11 11 2 11 2 13 9 1 9 2
9 15 13 10 9 13 3 1 9 2
10 3 13 3 0 9 1 9 10 9 2
35 1 10 0 12 9 4 10 9 13 10 3 0 2 3 0 9 2 15 4 4 2 13 1 15 1 9 7 9 2 7 13 13 9 3 2
9 13 16 10 9 4 13 12 9 2
10 9 2 9 2 9 9 7 3 3 2
33 9 9 4 0 7 13 1 10 0 9 2 15 15 13 13 1 12 9 3 2 7 1 3 13 15 1 9 1 12 9 13 9 2
8 15 4 10 0 9 1 9 2
37 9 4 1 10 9 3 4 13 9 4 13 9 1 10 0 9 1 12 9 2 1 0 9 2 1 3 12 9 2 7 1 3 12 9 3 3 2
14 9 13 1 10 9 1 9 1 11 9 2 11 11 2
5 15 4 9 9 2
10 10 0 9 1 10 0 9 1 9 2
16 15 13 11 11 1 11 9 1 14 13 0 9 1 9 3 2
7 12 9 4 13 1 9 2
11 15 4 3 3 13 1 10 9 0 9 2
14 1 11 11 2 12 9 2 4 9 13 10 3 0 2
11 7 9 4 13 10 9 2 15 3 13 2
53 10 0 1 10 0 9 2 15 1 0 4 13 9 1 0 7 0 1 10 0 12 9 2 13 2 16 10 9 3 13 1 10 0 9 2 3 10 13 9 2 10 0 9 2 10 13 2 10 13 7 10 13 2
25 10 0 0 9 2 3 10 13 9 11 11 2 13 10 3 0 9 1 10 0 9 9 11 11 2
31 15 4 3 3 13 9 1 14 13 10 0 9 1 10 0 9 2 15 11 11 4 13 1 9 7 9 1 10 0 9 2
16 15 13 9 1 9 7 9 2 15 13 10 9 9 1 9 2
15 2 15 4 0 0 13 1 14 13 9 2 2 13 15 2
21 3 0 4 3 13 1 9 1 9 1 9 1 12 9 7 12 9 12 9 3 2
5 15 13 1 9 2
19 2 15 3 13 15 3 2 13 9 2 16 11 4 13 1 9 1 11 2
24 10 0 9 1 11 4 13 9 1 14 13 1 9 2 7 15 13 10 0 9 4 4 9 2
8 9 9 4 13 1 0 9 2
7 9 4 3 13 1 11 2
25 15 13 3 1 14 13 7 13 1 3 14 13 9 2 15 3 4 13 2 1 9 1 15 15 2
7 15 4 9 9 1 9 2
8 15 4 0 14 13 1 9 2
5 0 9 1 9 2
1 9
22 7 9 3 13 9 7 10 9 3 9 1 11 9 2 7 3 4 15 4 3 0 2
2 9 11
28 11 1 9 11 2 2 11 4 10 3 0 9 2 3 9 13 3 3 2 15 4 10 9 2 15 4 13 2
14 2 3 10 0 2 15 13 2 15 4 3 13 15 2
7 2 3 4 15 10 9 2
5 11 13 15 9 2
12 3 4 15 13 9 7 9 7 13 1 9 2
10 15 13 10 9 1 9 7 0 9 2
7 3 4 15 3 1 9 2
26 15 4 2 1 3 11 7 11 2 4 13 3 1 9 2 15 4 13 15 1 10 9 1 11 9 2
24 10 0 9 11 13 1 9 2 16 9 3 4 13 9 1 9 1 9 1 1 13 1 9 2
21 15 4 13 2 16 0 9 13 1 9 2 2 13 9 11 2 15 13 1 9 2
4 12 13 1 9
6 2 9 2 11 11 2
12 3 13 15 12 9 7 10 0 9 0 0 2
13 7 1 10 9 4 15 0 9 1 1 12 9 2
10 9 4 1 9 13 1 9 1 11 2
17 9 13 1 12 9 1 10 0 1 12 1 10 9 1 11 12 2
11 9 13 14 13 2 16 9 13 1 9 2
1 9
13 7 1 9 13 15 2 16 15 4 13 9 3 2
23 3 13 10 0 11 11 2 9 2 9 1 9 2 1 12 9 9 1 9 2 0 9 2
17 1 0 9 9 1 9 13 9 9 1 11 1 9 9 3 13 2
16 1 9 1 11 11 4 15 3 4 9 1 9 1 11 11 2
12 11 4 3 1 10 10 9 13 1 0 9 2
21 11 11 11 4 9 1 12 9 7 13 15 3 13 1 11 11 1 11 8 11 2
28 9 1 9 0 9 4 3 0 2 3 12 13 9 2 1 16 15 4 13 9 1 2 16 3 0 4 13 2
6 12 9 7 12 9 2
10 11 13 12 0 9 2 9 7 9 2
6 9 1 10 0 9 2
36 11 11 11 13 2 16 9 4 3 0 2 16 15 4 13 1 12 9 1 12 9 1 9 1 14 13 15 1 9 7 1 14 13 10 9 2
8 2 4 15 3 3 10 9 2
18 1 10 0 9 2 0 0 9 2 4 10 0 9 13 3 1 9 2
12 15 13 0 7 3 13 11 1 10 0 9 2
25 1 10 0 9 4 15 4 3 0 1 10 9 2 15 13 1 9 2 1 0 9 2 9 2 2
6 2 6 15 13 3 2
14 3 13 10 0 9 1 9 7 10 9 9 1 9 2
18 2 15 4 0 1 2 16 15 13 12 9 7 12 9 1 10 9 2
10 9 0 9 4 13 3 1 0 9 2
31 1 10 9 2 3 3 3 13 9 1 9 2 16 3 13 3 0 2 16 15 13 0 9 1 9 2 13 15 1 9 2
9 2 9 1 9 4 13 3 3 2
6 7 11 13 10 9 2
6 0 9 13 1 11 2
5 11 2 15 13 15
10 16 9 13 9 2 13 15 10 9 2
2 0 9
22 2 15 13 9 1 9 13 3 2 0 9 3 7 0 9 3 3 1 10 0 9 2
38 7 1 12 9 9 4 15 13 3 2 7 16 10 0 9 1 9 13 13 3 15 7 9 9 1 14 13 3 1 10 0 9 9 2 13 15 3 2
9 12 9 1 9 1 10 0 9 2
24 1 10 9 1 12 9 13 11 12 12 8 13 1 9 2 15 9 1 9 4 12 9 0 2
33 9 11 4 3 13 10 0 9 2 16 11 1 0 9 13 15 1 10 3 0 9 1 9 1 14 13 1 12 1 10 0 9 2
39 2 1 9 1 9 0 9 1 9 13 9 3 2 16 3 4 13 3 1 9 2 7 9 13 3 3 2 16 3 13 9 1 10 9 1 9 3 2 2
2 9 13
22 10 0 9 1 10 0 9 7 9 1 10 0 9 1 11 4 13 10 0 0 9 2
33 1 9 1 9 4 10 9 1 14 13 10 13 9 13 1 1 10 2 9 2 2 16 9 9 4 13 1 3 13 9 1 9 2
11 7 1 13 2 10 9 4 3 10 9 2
10 13 14 13 15 1 9 7 9 9 2
11 15 4 3 13 15 15 1 14 13 15 2
36 16 15 13 1 10 9 2 3 15 4 10 9 2 16 15 13 13 9 1 9 2 4 15 3 13 2 16 15 3 13 3 0 9 1 9 2
7 2 15 4 3 13 11 2
42 1 10 3 0 7 0 9 1 9 4 9 2 9 11 11 11 2 13 10 9 1 2 3 15 13 3 2 2 9 4 4 3 0 2 16 15 3 13 10 0 9 2
25 3 13 10 13 11 14 13 11 1 9 7 13 14 13 1 9 7 13 3 1 9 1 0 9 2
11 7 9 13 3 10 12 9 3 1 9 2
