484 11
20 12 9 13 1 11 1 11 14 15 13 1 9 2 7 3 13 9 0 0 2
23 9 15 13 3 1 9 10 9 7 10 9 14 10 11 2 16 13 1 9 9 9 0 2
35 9 10 9 2 9 11 11 2 11 2 2 13 16 2 13 9 0 1 11 1 9 14 9 1 11 2 3 1 3 13 1 15 9 9 2
33 1 9 12 13 10 9 13 14 9 10 9 2 7 1 9 12 13 9 10 9 7 10 9 13 9 0 1 3 1 9 15 2 2
37 11 13 16 13 1 9 10 9 7 10 9 7 10 9 7 1 9 9 10 9 2 1 9 13 14 9 15 14 12 9 0 1 11 1 9 3 2
42 15 13 16 10 9 13 9 9 1 9 10 9 10 0 2 16 13 9 1 9 9 1 10 9 1 1 9 10 9 7 9 10 9 10 0 10 0 1 9 10 9 2
22 1 15 2 13 9 10 9 9 9 7 9 9 0 1 3 16 13 9 0 1 9 2
33 11 11 2 16 13 1 9 9 9 1 9 1 9 10 9 2 13 16 9 10 9 13 9 16 13 1 15 13 9 0 1 11 2
19 15 13 16 9 10 9 13 13 9 1 9 11 2 7 9 10 9 13 2
42 11 11 2 9 10 9 10 0 2 13 16 13 9 9 10 9 7 10 9 2 11 11 2 13 9 3 2 0 2 16 13 13 1 9 0 14 10 9 1 10 9 2
27 9 11 11 2 11 2 13 9 9 16 1 15 13 9 1 9 9 0 2 1 13 9 15 1 9 0 2
17 9 16 13 9 0 13 1 9 2 7 7 15 13 9 0 3 2
42 9 11 11 2 11 2 13 16 1 10 9 13 1 10 9 1 9 13 14 9 10 9 10 0 3 2 1 9 9 10 9 16 4 13 1 10 9 1 9 10 9 2
34 1 9 15 2 4 13 1 9 10 9 7 10 9 1 9 13 1 9 14 9 10 9 10 0 16 13 3 1 10 9 2 9 2 2
23 9 11 11 2 11 2 13 16 9 10 9 10 0 13 2 9 9 1 9 15 10 0 2
17 10 9 13 3 3 1 10 9 10 0 7 3 1 9 10 9 2
18 10 9 10 0 13 1 15 9 1 9 9 2 16 13 9 0 2 2
22 15 13 1 9 10 9 7 1 9 9 0 1 10 9 2 16 13 14 9 10 9 2
31 9 9 10 9 13 3 1 9 2 16 10 9 13 1 9 9 15 14 10 9 10 0 7 1 9 9 0 1 9 15 2
24 2 1 9 0 1 10 9 10 0 2 13 10 10 9 10 0 1 9 10 9 1 12 9 2
16 1 9 10 9 3 13 1 10 9 10 9 1 9 0 2 2
19 10 9 13 16 10 9 13 1 10 9 13 1 9 0 2 1 1 9 2
43 2 10 9 3 13 14 10 9 1 9 9 9 1 9 2 7 3 2 15 13 1 9 10 9 16 10 9 0 16 13 13 1 9 10 9 2 13 1 10 9 3 2 2
34 9 15 14 11 11 2 2 10 9 1 11 11 13 7 3 13 2 2 2 10 9 2 12 2 2 13 1 9 15 3 1 9 15 2
50 1 16 13 3 12 9 2 7 1 16 9 9 15 3 13 1 10 9 0 2 15 13 9 1 9 15 14 10 9 2 10 9 7 9 10 9 10 15 2 1 12 16 13 3 2 13 1 10 9 2
42 9 10 9 16 13 1 10 9 15 2 7 16 3 1 15 13 2 13 1 9 9 7 1 9 9 2 7 13 1 10 9 16 15 0 9 0 0 7 9 0 0 2
36 7 3 1 10 9 10 0 2 9 10 9 2 2 10 9 1 11 11 2 13 3 13 2 2 13 16 4 16 1 10 9 3 3 13 9 2
36 1 10 15 16 13 7 13 1 9 10 9 3 2 15 4 13 16 3 13 3 9 2 7 15 13 12 10 0 7 10 0 1 10 9 11 2
30 7 1 15 13 10 9 2 7 13 12 10 9 16 13 1 10 9 7 13 13 14 9 15 1 7 10 9 10 0 2
30 1 9 10 9 2 1 10 9 1 11 2 13 9 11 0 1 9 11 10 0 7 13 1 9 9 0 0 7 0 2
31 10 9 10 0 14 11 1 9 1 9 0 7 1 9 1 10 9 13 9 11 11 2 7 7 13 1 15 13 1 15 2
11 13 2 2 1 9 13 1 15 9 2 2
9 3 2 3 13 9 2 11 2 2
36 15 13 3 14 10 9 7 14 9 10 9 13 1 1 3 2 1 9 9 16 13 1 10 9 2 9 9 13 1 9 9 0 1 15 2 2
21 10 9 3 13 2 9 10 9 13 1 9 0 2 11 13 7 11 10 0 13 2
35 10 9 2 16 13 1 9 15 14 11 11 2 2 3 3 13 4 13 14 10 9 2 2 2 13 1 9 9 0 7 0 1 9 15 2
18 9 10 9 16 11 13 1 9 1 10 9 1 9 11 11 13 9 2
24 15 13 1 15 9 10 9 16 1 15 13 9 9 0 2 7 1 9 9 0 1 9 9 2
22 9 9 7 9 0 13 1 9 1 9 10 9 16 13 1 9 2 9 10 9 2 2
37 10 9 16 13 1 9 9 1 9 0 2 1 9 11 11 2 13 2 16 1 1 9 1 10 9 3 10 13 1 10 9 16 13 1 1 15 2
15 7 3 2 3 13 1 10 9 1 10 9 10 0 3 2
16 3 13 2 9 2 2 7 9 0 2 3 9 1 10 9 2
2 3 2
6 9 3 13 1 15 2
22 9 1 10 9 2 2 1 9 16 13 2 2 10 9 2 13 1 9 1 9 2 2
3 10 9 2
20 7 9 10 9 13 2 9 3 1 10 15 2 16 10 9 13 0 1 9 2
29 15 13 3 2 7 10 9 10 9 2 2 15 13 9 0 14 9 7 9 7 9 9 2 2 13 9 7 9 2
25 3 13 3 9 9 2 7 9 1 9 9 10 9 14 10 11 1 9 9 10 9 14 10 9 2
43 10 9 16 13 1 10 9 2 2 9 1 9 10 9 1 11 2 11 1 9 1 11 2 13 2 9 0 2 2 2 2 10 9 2 2 12 2 2 13 14 15 3 2
73 11 11 2 16 13 14 10 9 1 9 9 2 3 13 7 13 1 9 0 2 7 1 9 9 0 2 2 13 16 2 12 10 9 2 16 13 1 10 9 14 10 9 10 0 16 1 15 13 9 1 9 9 15 1 10 9 2 13 16 2 15 9 0 16 9 15 13 9 0 1 9 2 2
24 1 9 10 9 2 1 15 13 16 15 13 1 10 9 16 13 14 9 15 1 9 10 9 2
17 3 3 16 3 15 9 0 7 15 9 0 2 0 1 9 0 2
47 15 3 4 13 7 13 16 10 9 2 7 9 10 9 16 13 1 10 9 2 13 1 10 9 14 9 0 0 7 3 15 13 13 14 9 15 16 10 9 13 1 15 9 1 10 9 2
55 15 4 2 7 13 2 13 14 10 9 14 15 1 11 1 9 9 7 1 9 9 2 1 13 9 7 9 1 10 9 14 11 11 2 16 13 9 1 10 9 1 15 9 0 16 13 1 10 9 12 9 1 9 9 2
46 15 13 16 10 9 14 15 13 1 10 9 14 10 9 10 0 7 13 1 15 2 2 15 3 0 1 11 2 16 3 15 16 13 1 11 2 9 2 1 15 1 9 0 3 2 2
48 15 4 13 16 3 9 15 0 2 16 13 14 15 1 9 1 11 1 9 11 16 10 9 13 1 9 11 11 2 11 2 13 1 15 2 2 11 2 7 13 9 13 2 7 3 13 2 2
25 7 7 15 13 1 10 9 11 2 3 13 2 13 1 11 2 7 7 13 7 7 13 3 9 2
84 10 9 10 0 16 13 10 9 10 0 1 9 15 14 9 15 7 9 15 2 10 9 16 9 15 14 9 10 9 13 1 12 10 9 2 7 9 10 9 1 9 9 15 3 1 3 1 2 9 12 1 9 15 2 7 15 9 2 13 1 9 10 9 14 10 9 2 2 16 13 9 9 1 9 15 2 3 13 7 13 15 13 2 2
24 15 13 15 1 9 7 1 9 9 2 3 13 3 2 1 10 9 2 3 1 10 9 2 2
5 13 16 13 0 2
46 9 10 9 16 13 1 10 9 2 13 6 9 13 2 2 2 10 9 2 2 12 2 2 13 13 14 10 9 1 10 9 7 9 10 9 10 0 1 9 15 1 9 9 10 9 2
28 15 9 15 10 0 1 3 14 10 9 2 16 13 3 1 10 9 16 15 13 3 3 1 9 15 10 0 2
30 7 10 9 9 13 3 1 10 9 10 0 2 13 10 9 1 9 3 13 14 9 9 0 2 0 9 7 0 9 2
23 13 10 9 16 10 0 1 10 9 10 15 16 13 4 13 1 9 9 15 13 10 9 2
24 15 3 13 1 9 1 9 7 1 9 2 7 7 1 9 0 2 7 3 1 9 9 0 2
48 9 1 9 9 7 9 9 0 2 1 9 10 9 10 0 7 1 9 9 13 3 1 9 0 2 7 14 4 13 14 10 9 1 9 9 7 9 2 13 9 15 14 15 1 9 10 9 2
26 15 13 1 2 10 9 2 16 13 13 1 9 15 14 10 9 2 10 4 13 1 10 9 10 0 2
31 1 9 0 13 9 15 14 11 11 2 9 9 9 10 9 7 9 10 9 2 1 10 9 2 3 13 1 10 9 2 2
37 1 9 15 13 9 12 1 9 15 2 2 15 2 9 10 9 2 13 1 9 15 10 0 3 1 9 0 2 7 1 10 9 7 10 9 2 2
18 9 1 9 2 16 13 3 14 3 16 10 13 3 13 1 9 0 2
17 15 3 10 9 16 13 14 9 10 9 7 9 10 9 10 0 2
30 9 2 1 2 15 2 10 9 1 11 3 1 9 13 1 10 0 3 1 10 9 2 7 3 10 0 16 1 15 2
15 7 7 1 10 9 7 1 10 9 10 9 13 10 9 2
27 1 10 12 1 11 13 1 10 9 11 11 2 1 10 9 10 0 14 9 10 9 2 10 9 11 11 2
17 3 15 3 13 1 10 9 10 0 1 9 1 10 9 10 0 2
21 2 3 13 9 1 9 2 2 13 1 15 10 9 1 9 9 1 9 9 0 2
17 2 3 9 2 2 13 10 9 2 2 13 3 1 9 0 2 2
7 11 13 9 3 2 0 2
22 13 1 15 2 16 13 1 15 3 9 0 1 9 0 7 1 10 9 0 14 11 2
20 9 13 13 1 11 1 9 0 2 4 13 14 15 3 1 9 7 9 9 2
24 11 13 1 9 10 9 14 11 2 7 1 9 15 15 13 14 15 1 9 1 9 10 9 2
38 1 12 13 11 2 3 1 9 0 0 1 10 9 10 0 2 1 9 0 2 10 9 11 11 13 13 9 9 1 10 9 2 1 9 15 1 11 2
11 11 13 14 10 9 1 9 9 10 12 2
24 9 15 13 13 1 9 0 2 1 9 16 10 10 9 10 0 1 11 13 1 9 0 9 2
17 3 3 9 0 13 7 1 11 9 1 9 2 7 3 9 0 2
15 3 3 13 3 14 10 9 14 9 1 10 9 10 0 2
32 9 12 1 10 9 16 13 13 10 9 10 0 2 11 11 11 2 9 0 1 9 9 10 9 10 0 14 9 15 10 0 2
13 2 2 13 10 9 1 11 2 2 9 3 2 2
17 1 10 9 10 0 13 10 9 14 9 9 10 9 1 9 11 2
17 1 9 0 13 10 9 1 9 9 10 9 14 15 9 0 9 2
29 13 1 15 9 10 9 0 9 2 7 1 9 15 13 10 9 2 2 13 14 9 2 11 3 13 3 11 2 2
8 2 11 2 13 3 11 11 2
30 2 13 14 9 2 2 13 9 1 9 10 9 10 0 14 10 9 1 12 2 2 13 14 9 3 13 9 0 2 2
59 1 9 9 9 1 11 11 2 10 9 10 0 16 13 14 15 3 1 9 0 2 13 1 15 1 9 12 10 13 3 4 11 13 14 9 10 9 10 0 2 2 7 3 13 14 10 9 1 9 10 9 10 3 2 0 2 1 11 2
9 13 1 9 9 15 1 9 0 2
20 9 1 10 15 2 16 3 13 0 1 9 1 11 2 3 13 3 10 9 2
52 1 9 10 9 10 0 14 11 4 13 16 10 9 13 1 9 11 2 16 15 0 9 0 7 0 2 7 16 10 9 10 0 14 9 16 9 2 13 11 2 3 3 13 1 9 13 9 0 1 11 11 2
15 10 9 1 10 9 10 0 3 13 9 9 0 1 11 2
32 11 11 10 0 2 7 9 15 10 0 10 0 11 11 2 3 3 13 13 1 10 9 2 7 13 13 1 10 9 10 0 2
15 15 13 1 10 9 2 7 15 13 1 10 9 1 9 2
19 1 9 10 9 10 0 13 11 3 2 9 13 2 7 11 13 9 13 2
44 11 13 1 10 9 9 0 0 2 7 13 14 10 9 1 9 9 11 2 11 13 9 0 1 9 10 9 2 7 13 1 9 10 9 1 10 9 1 10 9 1 10 11 2
18 1 10 9 10 0 15 9 0 2 7 9 0 2 1 9 3 0 2
29 1 9 9 13 9 7 1 9 10 9 13 3 9 0 14 9 0 2 9 0 14 9 10 9 10 0 10 0 2
24 1 9 9 10 9 13 9 15 14 11 9 9 2 16 12 1 9 15 13 9 1 9 9 2
32 1 9 10 9 10 3 2 0 1 11 2 9 1 9 9 13 14 10 9 1 9 1 10 9 3 7 13 13 3 1 11 2
22 9 3 2 0 13 3 7 3 9 13 9 1 9 2 16 13 1 9 9 10 9 2
29 3 2 11 11 2 9 0 1 9 10 9 2 13 12 10 9 10 0 3 14 9 0 1 12 10 9 10 0 2
23 1 9 0 1 11 2 11 13 12 12 9 1 9 9 0 3 2 0 1 10 9 11 2
6 11 13 3 12 12 2
25 1 12 13 9 11 11 11 14 11 1 12 1 12 7 12 9 2 16 13 1 2 9 0 2 2
16 15 13 9 3 2 0 2 7 13 9 16 13 1 15 3 2
39 7 2 1 2 9 2 15 2 9 3 2 0 1 11 13 3 14 9 15 1 9 9 1 9 10 9 2 16 11 13 1 11 1 9 13 14 12 9 2
17 15 10 9 10 0 10 0 1 9 11 16 13 1 9 9 12 2
39 15 3 13 2 16 1 9 1 9 1 9 9 15 10 0 2 13 13 10 9 1 9 9 10 9 10 0 10 0 2 16 1 15 3 9 0 4 13 2
16 9 1 11 2 16 13 3 1 10 9 1 9 9 10 9 2
39 9 9 10 9 10 0 13 3 16 10 9 13 9 0 14 12 9 2 13 1 10 9 10 0 2 1 10 9 16 13 1 9 10 9 1 12 9 3 2
49 9 9 10 9 10 0 2 11 11 2 13 16 10 9 13 1 10 9 1 9 9 16 13 3 3 7 13 1 10 9 10 0 2 14 10 9 13 1 9 15 2 3 7 9 9 1 10 9 2
35 10 9 13 13 16 13 13 9 0 14 9 0 1 10 9 2 1 10 9 10 0 16 13 1 9 15 3 1 9 10 9 1 10 9 2
39 1 10 9 10 0 13 9 9 10 9 2 11 11 2 1 9 9 10 9 2 11 9 2 1 9 10 9 13 9 0 16 13 1 9 13 1 10 9 2
18 11 13 16 10 9 13 10 1 9 9 15 14 10 9 1 10 9 2
38 9 9 10 9 10 0 13 3 9 9 7 1 9 10 9 10 0 3 13 9 9 1 10 9 10 0 2 1 9 15 13 9 10 9 1 12 9 2
7 9 10 9 13 1 11 2
22 9 9 9 10 9 2 11 11 2 13 1 9 11 1 9 9 1 9 2 10 9 2
23 11 13 3 1 10 9 2 1 9 15 1 10 9 11 1 11 1 9 10 9 14 15 2
13 9 13 1 9 15 2 7 15 13 1 10 9 2
18 11 11 4 13 13 1 11 1 11 2 7 1 15 1 11 2 11 2
13 3 13 4 13 1 9 15 2 16 13 1 11 2
14 9 10 9 11 13 13 3 1 2 10 9 1 11 2
17 9 9 15 14 11 13 3 3 1 10 9 1 9 9 10 9 2
21 10 9 2 16 13 1 10 9 1 10 9 2 3 13 14 9 15 1 9 15 2
14 9 11 13 1 9 15 14 9 15 1 9 10 9 2
29 10 9 13 1 9 10 9 10 0 2 16 13 14 10 9 1 10 9 10 0 1 11 2 16 13 1 9 11 2
8 10 9 1 11 13 1 11 2
26 1 9 10 9 1 11 13 9 13 1 9 10 9 1 9 10 9 2 7 3 13 9 1 9 15 2
23 3 1 2 15 13 9 9 2 7 1 15 9 15 7 9 15 14 11 1 9 9 0 2
23 9 9 10 9 13 3 1 10 9 2 7 3 3 13 16 13 1 9 9 9 10 9 2
22 11 2 9 12 1 9 15 2 13 1 15 9 2 9 2 9 2 9 7 12 9 2
8 3 3 13 9 1 9 15 2
36 9 10 9 1 9 10 9 1 10 9 2 2 11 2 2 13 1 3 1 3 9 9 7 1 15 9 1 16 13 1 10 9 1 9 0 2
16 10 9 0 3 2 1 9 9 13 1 15 9 1 9 9 2
25 2 11 2 13 13 14 9 10 9 14 15 1 9 9 0 2 9 15 9 9 1 9 10 9 2
31 1 9 15 13 1 9 10 9 9 1 9 10 9 2 1 9 0 2 7 15 9 15 2 2 10 9 10 9 14 15 2
11 3 13 1 15 10 9 16 13 1 15 2
16 1 15 15 13 1 15 3 3 7 15 13 3 1 10 9 2
8 13 15 13 1 15 9 15 2
11 9 9 15 13 1 9 9 9 3 2 2
15 1 10 9 11 11 2 10 9 1 9 10 9 7 9 2
25 7 1 3 16 13 3 14 9 15 14 9 10 9 1 10 9 10 0 10 15 2 3 9 9 2
57 1 9 10 9 16 9 11 13 1 9 15 1 10 9 13 9 1 15 10 9 2 2 7 13 1 15 9 9 1 9 10 9 2 3 13 1 9 10 9 1 10 9 2 1 13 1 9 0 13 7 13 14 9 10 9 2 2
5 10 9 1 15 2
4 10 9 13 2
24 9 15 14 9 0 13 3 1 10 9 2 7 3 3 13 1 9 2 9 2 14 9 11 2
4 3 15 3 2
58 9 9 10 13 3 2 1 3 2 3 1 15 1 13 1 9 2 1 9 2 1 9 7 1 9 1 9 0 1 9 9 10 9 9 15 13 1 9 10 9 10 0 2 14 1 9 15 13 10 9 16 3 3 15 13 1 15 2
25 1 1 9 9 2 12 10 13 7 13 1 9 16 13 1 15 1 10 9 13 13 0 10 3 2
16 7 3 2 1 9 0 2 13 16 15 3 3 16 15 0 2
6 13 7 14 11 11 2
10 1 9 15 13 1 10 13 0 0 2
30 7 1 9 1 0 13 16 15 13 1 13 11 11 11 2 9 1 9 9 7 1 9 1 11 11 2 11 2 11 2
7 3 15 4 13 1 15 2
19 7 13 3 10 13 10 0 1 10 9 16 3 0 1 9 14 10 9 2
49 1 16 9 9 11 13 13 14 10 13 1 9 10 9 1 9 15 2 10 9 13 3 1 9 16 13 3 13 1 13 1 9 7 1 9 9 2 10 9 10 0 14 10 9 13 11 11 2 2
44 7 1 10 15 15 13 9 1 9 15 7 1 9 15 2 1 15 13 14 15 1 10 9 10 0 2 13 1 10 9 2 7 13 9 9 9 16 15 4 1 9 1 15 2
4 3 10 9 2
8 9 9 12 2 13 1 9 2
19 3 10 12 1 12 12 10 9 16 9 0 13 3 9 13 13 1 0 2
13 15 12 10 9 1 15 16 9 11 0 10 3 2
39 1 9 9 13 10 9 1 9 2 1 9 9 2 2 13 9 9 2 2 1 9 1 9 0 2 1 9 2 1 9 7 1 9 0 3 1 9 9 2
20 16 15 2 3 10 1 15 13 1 9 9 0 1 12 1 12 10 9 15 2
49 3 4 13 1 9 1 9 0 3 7 3 2 7 13 1 10 9 9 1 14 15 1 9 10 9 13 10 9 2 1 16 13 10 9 14 15 13 9 0 1 10 9 1 13 2 9 0 2 2
20 7 15 13 13 1 9 9 2 15 4 13 9 1 14 15 3 1 9 9 2
36 3 13 9 10 9 9 10 9 10 0 11 11 2 16 13 14 2 10 9 1 9 0 3 2 2 16 13 9 1 9 1 13 9 9 0 2
44 3 2 1 16 13 9 0 1 9 1 10 9 14 15 3 1 9 9 13 11 14 10 9 10 0 1 9 10 9 14 15 16 0 3 1 13 9 7 1 9 0 1 15 2
10 7 3 13 13 1 10 9 10 0 2
28 10 9 1 2 16 3 1 9 9 2 7 1 2 1 9 9 2 0 3 2 7 1 9 9 9 0 3 2
34 10 9 10 0 3 1 9 1 10 9 10 0 13 10 9 1 9 9 11 1 9 12 9 14 10 9 14 9 11 3 2 11 11 2
34 10 9 13 13 14 10 9 1 9 9 2 10 9 14 2 11 11 11 2 2 9 16 1 9 9 13 1 15 9 12 12 9 0 2
4 9 9 12 2
8 13 13 9 9 7 9 0 2
17 1 10 9 2 9 13 1 9 2 13 11 11 1 9 10 9 2
66 9 0 1 9 15 14 9 2 7 14 9 7 9 0 2 13 3 1 9 10 9 14 15 2 1 10 9 10 0 14 10 9 2 1 9 2 1 9 9 7 1 9 0 2 16 9 10 9 16 4 13 1 15 13 9 9 13 16 13 14 15 7 13 14 15 2
11 12 9 1 9 10 9 13 1 9 0 2
23 1 9 9 16 4 13 1 9 0 0 3 7 9 9 0 1 9 2 15 9 0 3 2
35 1 10 10 9 2 1 9 1 10 9 13 1 9 16 10 9 1 15 0 3 2 1 9 9 7 9 1 9 10 9 7 9 10 9 2
34 3 3 1 9 13 1 9 10 9 10 0 16 1 15 13 1 9 10 9 9 7 9 1 9 10 9 7 1 9 10 9 10 0 2
20 1 9 9 15 2 16 9 15 13 11 2 10 9 10 0 13 10 0 3 2
4 9 9 12 2
11 13 0 1 10 9 10 0 14 9 15 2
41 2 15 13 1 9 16 13 9 9 0 1 9 2 7 1 15 1 10 9 13 14 9 15 14 9 10 9 2 2 13 11 11 2 9 9 10 9 1 9 11 2
37 1 12 9 13 11 13 9 0 1 9 9 10 9 10 0 2 9 1 9 9 16 1 15 13 1 12 10 9 10 0 2 10 9 10 0 2 2
14 3 13 1 10 9 7 13 14 9 10 9 14 15 2
4 9 9 12 2
6 13 13 14 10 9 2
31 1 9 10 10 9 13 1 10 9 10 0 9 0 1 10 9 1 9 9 1 9 10 9 16 13 1 15 9 0 0 2
22 11 13 16 1 9 10 12 7 10 12 15 4 13 13 1 9 1 9 11 7 11 2
18 9 15 10 0 14 11 13 9 1 9 11 13 1 9 9 10 12 2
30 3 15 13 9 1 10 9 16 13 1 9 10 9 2 7 9 10 9 13 9 1 9 10 9 10 0 1 9 9 2
7 13 13 16 15 9 0 2
32 11 13 16 9 10 9 13 9 9 16 13 1 9 9 13 2 9 16 1 9 15 4 13 13 9 0 1 9 9 10 9 2
10 7 15 3 13 3 0 1 10 9 2
21 9 11 13 13 0 16 10 9 13 3 14 10 9 1 9 9 10 9 1 9 2
10 11 3 4 13 13 15 1 9 0 2
29 1 3 12 13 9 9 10 9 10 0 1 2 9 9 10 9 10 0 2 10 9 10 0 3 1 9 9 0 2
4 9 9 12 2
5 13 9 1 9 2
17 13 9 16 13 13 1 9 9 16 15 13 9 1 9 0 0 2
35 1 9 15 4 13 1 9 2 13 3 9 0 16 4 13 9 7 16 3 13 13 2 7 13 14 15 1 9 9 1 9 2 13 9 2
22 10 9 13 3 7 3 9 0 1 10 15 1 10 9 16 13 1 9 7 1 9 2
34 3 15 13 13 9 16 16 15 4 16 3 13 13 3 2 9 7 9 2 9 7 9 9 2 0 14 10 9 7 0 14 10 9 2
25 7 13 2 4 16 9 10 9 14 10 9 13 3 15 1 10 9 2 13 7 1 9 10 9 2
29 13 16 9 10 9 7 10 9 14 9 11 1 11 16 1 11 13 9 0 1 9 9 1 9 0 14 10 9 2
19 3 7 3 13 9 0 1 9 15 2 0 1 0 16 13 9 14 9 2
26 1 9 16 13 13 1 9 15 13 9 0 7 1 9 9 10 9 7 10 9 16 13 1 9 9 2
46 3 15 4 16 1 9 9 7 9 9 13 10 9 2 11 11 11 2 14 12 10 9 10 0 2 7 3 0 16 13 1 15 10 9 16 13 9 1 9 0 1 9 0 7 0 2
4 9 9 12 2
13 13 9 0 2 13 7 0 2 1 9 0 0 2
24 15 1 12 9 13 9 9 2 1 15 11 11 2 13 9 0 1 9 0 3 1 10 9 2
56 15 13 16 13 9 1 15 16 9 9 13 1 9 9 1 9 0 2 7 10 9 13 3 0 9 14 3 1 10 9 1 9 10 9 2 10 9 16 13 11 11 1 9 11 2 2 16 1 9 15 14 9 13 14 15 2
36 11 7 9 15 10 0 13 12 9 2 3 2 15 13 9 13 14 10 9 14 15 1 10 9 1 10 9 14 9 15 2 1 9 9 11 2
21 3 2 15 13 14 10 9 1 10 9 13 9 0 3 1 9 9 1 9 0 2
15 9 1 9 15 9 13 16 3 13 15 9 14 10 9 2
27 2 9 3 13 4 13 9 16 1 15 4 13 9 0 2 2 13 11 11 2 12 10 9 1 10 9 2
53 11 2 16 13 14 9 11 2 11 7 3 13 14 9 11 2 13 16 10 9 3 13 10 2 3 13 9 1 10 9 10 0 14 1 15 2 7 13 9 1 10 10 9 10 0 16 13 1 3 9 7 9 2
21 15 7 11 7 10 0 3 13 16 2 0 9 0 14 9 16 4 1 9 2 2
16 15 3 13 2 13 11 2 2 1 3 13 9 0 2 2 2
52 3 2 13 16 9 10 9 10 0 13 9 1 11 11 2 11 11 2 11 11 7 11 11 16 3 1 1 10 9 10 0 16 13 1 9 10 12 7 7 1 9 9 10 12 13 9 13 15 1 10 9 2
84 7 15 13 1 10 9 9 1 15 16 11 7 9 13 14 10 9 1 9 15 2 7 7 3 9 0 13 16 13 1 10 9 1 9 10 9 2 15 13 14 15 1 9 10 9 10 0 10 0 3 2 7 13 1 15 16 1 10 9 10 0 11 2 11 2 11 2 11 7 11 11 2 11 2 11 11 3 11 13 1 9 10 9 2
3 3 0 2
33 7 3 15 3 2 7 0 3 16 9 11 2 10 9 10 0 3 1 10 9 10 0 14 9 10 12 2 3 4 1 9 15 2
29 1 10 9 13 10 9 12 9 1 9 11 1 9 15 14 11 11 13 14 9 10 9 7 9 10 9 14 11 2
14 3 13 9 1 10 15 1 9 9 3 1 9 0 2
26 7 10 9 13 9 11 1 9 0 16 13 1 9 15 7 13 13 1 9 0 1 9 0 0 9 2
29 1 15 2 3 10 9 9 10 9 10 0 13 3 9 10 9 10 0 10 0 16 16 1 9 0 13 14 15 2
28 9 11 3 4 13 3 7 3 12 9 1 9 2 9 7 9 0 2 9 1 9 1 9 3 2 0 2 2
23 7 15 4 13 1 12 9 9 11 10 0 1 13 9 9 16 4 10 3 13 1 15 2
34 16 1 9 11 9 13 16 9 9 0 1 9 1 9 10 9 2 9 9 12 2 13 0 2 16 15 13 2 13 9 1 9 0 2
46 7 13 9 16 9 0 1 12 12 10 9 16 1 15 9 10 9 13 1 9 1 2 11 2 2 1 2 13 14 9 10 9 10 0 1 10 11 11 10 0 14 11 2 11 2 2
66 1 15 2 2 9 10 9 2 2 10 9 10 0 1 9 16 13 9 11 1 12 2 13 9 0 2 1 9 9 0 3 14 9 0 2 1 9 9 7 9 0 7 0 3 2 16 3 13 9 9 2 7 3 13 16 10 9 13 1 9 9 10 9 1 9 2
25 13 1 10 15 2 3 15 13 1 10 0 9 15 14 10 9 1 10 9 7 3 3 1 15 2
18 16 13 10 9 1 9 0 2 9 0 13 3 1 10 9 14 15 2
21 3 13 9 1 9 10 9 2 10 9 10 0 1 10 9 1 10 9 10 0 2
19 9 0 13 1 9 1 13 14 10 9 10 0 14 15 1 9 9 0 2
33 1 10 9 7 10 9 13 1 9 3 0 14 9 1 9 2 13 3 9 1 11 14 9 15 1 9 0 1 13 14 10 9 2
4 9 9 12 2
8 13 9 9 14 9 10 9 2
15 1 10 9 0 2 9 16 13 1 9 0 13 7 13 2
45 1 9 9 10 12 13 7 13 1 9 10 9 10 3 2 0 1 2 10 9 1 9 7 9 2 7 1 2 9 0 2 2 7 10 9 13 1 9 1 9 10 9 10 12 2
15 3 13 10 9 1 11 7 11 11 7 9 9 10 9 2
23 3 3 3 13 10 9 10 0 1 10 9 10 3 2 0 9 0 0 2 7 9 0 2
25 10 9 10 3 2 0 13 3 15 16 13 9 1 3 2 13 1 10 9 3 13 1 10 9 2
27 3 2 14 10 9 10 0 13 2 13 9 13 9 7 9 9 0 16 13 14 9 9 15 14 9 9 2
4 9 9 12 2
8 13 7 13 1 9 9 0 2
29 13 16 9 10 9 13 13 2 9 0 2 2 9 3 2 0 0 2 7 13 14 15 1 9 10 9 14 15 2
28 9 10 9 10 0 10 3 2 0 13 16 3 3 2 4 3 13 1 9 0 1 2 9 9 10 9 2 2
33 10 9 13 10 9 10 0 2 16 0 1 9 0 3 2 13 16 10 9 13 4 13 0 7 3 13 2 9 9 0 0 2 2
55 7 9 1 9 9 10 9 10 0 2 3 1 9 1 9 10 9 1 9 2 13 1 9 13 9 15 1 9 9 10 9 2 1 9 16 1 10 9 13 10 9 10 0 1 9 14 9 9 0 2 3 14 9 0 2
8 1 9 15 11 11 13 9 2
42 7 11 11 13 9 2 9 1 10 10 9 1 9 3 2 0 1 10 9 2 16 13 15 9 16 4 13 14 9 15 14 9 0 1 9 0 1 10 9 10 12 2
30 13 1 9 9 16 13 13 1 15 9 9 1 9 16 10 9 13 9 1 9 0 7 9 3 2 0 1 10 9 2
35 9 15 13 9 1 9 0 1 9 10 9 2 9 15 14 9 7 9 9 1 9 0 13 1 15 16 10 9 3 0 1 9 0 0 2
68 11 11 11 2 9 10 9 2 10 9 14 10 9 2 9 9 7 9 15 14 9 9 0 2 2 13 16 10 9 1 9 9 13 2 7 9 10 9 1 9 15 14 9 0 1 9 10 9 2 13 14 15 1 9 0 14 9 2 16 1 15 4 13 16 13 10 9 2
3 15 0 2
34 1 9 2 10 9 1 9 9 13 1 9 10 9 10 0 1 10 9 10 0 1 9 13 1 3 9 9 1 11 11 4 13 0 2
12 10 9 13 3 13 9 0 1 9 9 0 2
19 13 9 1 10 9 16 3 15 13 12 10 9 10 13 3 14 10 9 2
31 7 4 13 1 9 2 16 10 3 9 12 1 3 1 12 12 10 9 16 13 9 1 12 1 12 3 13 1 9 15 2
25 3 10 9 13 14 10 9 7 16 13 10 9 1 9 0 1 9 15 7 10 9 16 1 15 2
48 1 13 1 9 15 1 15 13 3 1 10 1 3 2 15 9 0 1 9 15 14 10 9 2 7 13 9 1 9 0 2 1 9 1 9 15 14 10 9 10 0 1 10 9 7 3 3 2
16 7 15 13 9 1 10 9 16 4 13 1 15 1 9 0 2
25 10 9 13 9 9 1 9 10 9 1 9 9 9 4 13 1 10 9 10 0 1 1 10 9 2
14 9 9 3 13 1 10 1 9 10 9 14 10 9 2
50 10 9 13 1 10 9 7 1 10 9 2 7 1 12 9 2 2 12 2 9 13 13 3 1 10 9 10 0 2 7 3 15 16 13 1 3 13 13 13 13 13 1 10 9 10 0 7 13 13 2
21 3 12 9 1 15 13 1 9 11 1 10 9 1 10 9 7 1 9 10 9 2
16 2 12 2 9 10 9 3 13 9 10 9 10 0 10 0 2
50 1 11 13 3 3 3 1 12 9 1 9 9 10 9 1 10 9 2 3 1 16 13 1 9 0 2 7 1 9 0 2 7 1 16 13 14 10 9 16 13 1 9 9 10 9 1 9 9 15 2
28 4 3 16 1 10 9 1 10 9 13 9 15 14 10 9 10 0 1 10 9 2 11 11 2 1 10 0 2
20 3 3 1 10 9 1 10 9 13 3 10 9 11 11 13 2 1 9 0 2
36 9 15 14 9 9 1 10 9 10 0 13 13 3 3 10 13 13 13 2 7 7 3 15 13 13 10 4 16 1 10 15 13 1 10 9 2
33 1 9 9 11 2 9 9 11 16 13 1 9 9 11 2 13 9 0 1 3 2 10 9 14 9 9 9 1 10 9 10 0 2
11 15 13 9 14 3 2 9 1 10 15 2
22 10 9 13 1 15 9 0 1 10 9 10 0 14 10 9 10 0 2 1 9 11 2
16 15 13 14 9 15 2 14 9 15 7 14 11 1 10 9 2
20 1 9 9 10 9 10 0 13 11 14 10 9 10 0 1 3 2 10 9 2
15 2 9 2 2 13 2 2 13 1 9 10 9 3 13 2
15 9 9 2 10 9 10 9 10 0 13 9 14 9 15 2
28 16 13 1 15 9 2 16 3 15 13 2 7 13 2 3 13 2 3 15 13 3 15 2 7 3 15 13 2
5 3 15 10 9 2
9 3 15 9 2 16 13 13 15 2
14 3 15 10 9 2 16 13 13 9 0 1 10 9 2
8 7 3 15 13 7 13 2 2
38 1 10 9 16 13 14 10 9 10 15 1 9 11 13 10 9 2 11 11 2 9 2 16 13 3 9 1 11 1 9 9 15 10 0 2 11 11 2
21 1 9 13 10 9 1 12 9 2 7 1 11 13 9 13 1 9 15 14 11 2
9 15 13 3 1 9 14 12 9 2
23 11 13 3 10 9 10 0 10 0 2 10 0 7 10 0 3 1 9 10 9 14 12 2
23 15 9 0 2 16 13 1 9 13 1 10 9 16 13 2 7 1 10 9 14 9 0 2
14 15 13 9 0 1 9 9 0 7 1 9 9 0 2
28 15 13 1 10 13 14 9 15 2 2 9 9 2 13 9 1 10 9 2 2 13 1 15 1 9 0 2 2
10 15 13 1 9 0 1 9 9 0 2
32 1 15 15 3 13 9 0 0 2 9 2 16 1 15 13 3 1 10 9 0 14 9 10 9 1 11 2 7 13 9 0 2
17 15 13 10 1 9 15 16 13 1 15 10 9 16 0 13 9 2
12 7 9 15 7 9 15 13 9 1 9 15 2
33 7 1 11 11 11 13 16 13 1 15 2 9 1 9 12 7 9 1 9 0 2 2 3 1 11 13 4 13 3 14 10 9 2
102 1 10 12 1 11 13 1 15 9 9 1 10 9 2 11 11 2 1 9 16 0 1 9 9 12 2 2 15 13 1 9 0 1 9 10 9 3 16 13 1 10 9 9 1 13 1 9 0 2 7 9 13 9 0 2 15 13 13 1 9 10 9 2 11 3 0 2 1 16 15 13 1 11 13 1 11 2 7 13 2 13 1 9 15 10 9 13 1 15 13 9 1 9 15 10 0 2 16 13 11 2 2
36 7 3 10 9 10 15 10 9 13 12 9 0 9 1 9 15 14 9 0 13 9 0 14 9 9 1 9 15 14 10 0 10 0 11 11 2
21 15 0 2 0 2 4 13 1 9 15 2 7 13 14 10 9 3 3 1 9 2
22 7 13 11 2 4 3 16 13 13 1 9 2 7 1 12 9 2 13 1 10 9 2
31 11 11 2 9 1 9 11 2 16 11 13 3 1 9 15 1 9 9 1 9 2 13 3 1 9 15 1 9 10 9 2
13 15 13 7 4 13 15 13 1 10 9 10 0 2
8 2 3 3 2 2 2 13 2
11 2 3 1 11 11 9 3 13 13 2 2
14 10 9 10 15 2 1 10 9 15 2 13 1 15 2
16 11 13 3 1 10 9 2 13 7 0 3 1 3 2 3 2
20 10 9 10 0 1 11 13 3 14 9 15 1 10 9 10 0 2 1 12 2
12 3 13 3 3 10 9 2 7 3 10 9 2
19 3 12 9 1 12 10 9 10 0 3 13 9 13 7 13 2 7 13 2
17 1 1 9 3 13 9 0 13 16 11 11 13 10 9 10 12 2
52 7 1 3 13 11 1 9 15 1 9 10 9 2 13 1 9 2 9 1 10 9 2 7 13 3 1 10 10 9 2 13 1 9 10 9 16 13 1 15 9 0 13 14 11 1 10 9 10 0 1 9 2
10 13 3 10 9 16 13 13 1 15 2
7 3 13 10 9 1 12 2
66 10 9 14 10 9 13 13 9 0 1 12 1 10 9 10 13 3 2 10 9 0 2 10 9 14 9 11 11 2 11 11 2 16 9 15 13 1 9 0 1 3 12 2 7 10 9 1 11 11 2 10 9 7 9 10 9 10 0 14 9 10 12 2 11 11 2
15 9 15 3 13 10 9 12 1 9 1 9 9 10 9 2
15 10 9 10 0 13 1 10 9 13 9 0 9 1 9 2
9 11 13 3 1 9 14 12 9 2
46 1 9 9 10 9 13 9 1 3 2 9 1 10 9 2 7 13 1 9 0 16 7 13 13 13 1 9 10 9 1 11 11 2 13 13 1 9 10 9 10 0 2 11 11 11 2
26 7 16 15 13 1 15 9 13 1 10 9 2 15 13 1 9 9 0 1 12 9 1 15 14 11 2
27 11 11 13 10 9 10 0 3 1 10 9 1 3 13 9 13 1 9 10 9 10 0 2 1 9 12 2
34 9 10 9 14 15 2 10 9 10 0 2 10 9 7 10 9 13 9 0 1 11 16 15 13 9 12 10 9 10 0 1 11 11 2
30 10 9 16 13 9 10 3 3 0 1 9 10 3 3 0 13 13 3 16 9 15 13 1 10 9 10 0 13 3 2
14 15 13 1 15 2 16 9 1 10 9 14 15 13 2
26 1 9 13 16 13 1 15 12 1 15 16 13 13 14 15 2 3 7 3 2 9 0 1 10 9 2
28 1 10 12 10 15 13 12 9 1 9 2 7 12 9 0 13 1 10 9 1 9 15 14 10 9 14 15 2
10 1 15 13 1 10 9 12 9 9 2
16 9 9 1 9 0 13 9 9 1 9 9 10 9 10 0 2
29 1 9 16 13 3 10 1 9 10 9 2 9 10 9 13 3 0 1 15 9 16 13 9 9 9 10 9 11 2
29 10 9 10 15 13 1 9 2 3 1 9 2 2 13 3 11 11 2 16 13 1 10 9 10 0 1 10 9 2
20 9 15 10 0 14 9 15 2 11 2 13 4 13 10 9 1 9 9 15 2
16 1 9 15 14 9 13 16 10 9 13 9 2 7 11 13 2
6 7 10 9 3 13 2
25 7 13 9 0 14 9 10 9 10 0 14 11 2 14 11 2 14 11 2 14 11 7 14 11 2
10 1 10 10 9 10 15 13 11 11 2
16 1 9 12 15 4 13 1 9 10 9 10 0 3 1 11 2
21 15 13 3 1 9 11 2 1 9 9 10 9 10 0 7 10 0 3 14 12 2
35 11 13 3 1 10 9 10 0 1 11 2 16 13 13 14 10 9 10 0 1 9 10 9 10 0 2 9 10 9 1 10 9 14 12 2
23 10 9 13 1 9 9 2 7 13 16 9 15 11 3 13 7 13 1 10 9 10 0 2
23 15 4 13 1 3 1 9 2 1 10 9 7 10 9 16 13 10 9 10 0 11 11 2
12 11 13 12 9 1 9 0 9 0 1 11 2
33 2 11 10 0 2 2 13 11 1 10 9 10 0 10 0 14 15 2 2 15 3 0 2 15 13 1 9 9 1 10 9 2 2
41 15 13 9 3 1 13 9 9 2 7 3 1 9 15 13 10 9 13 14 10 9 10 3 2 0 1 10 9 10 3 2 0 7 1 10 9 10 3 2 0 2
38 11 13 1 9 16 10 9 16 15 13 1 15 14 10 9 13 1 10 9 1 9 9 2 16 9 9 15 13 1 3 3 2 9 0 1 9 0 2
8 3 13 11 9 0 1 9 2
29 16 13 13 1 9 9 15 1 9 2 13 1 15 12 9 0 2 16 13 9 16 15 13 1 10 9 1 9 2
10 11 3 13 14 9 15 1 10 9 2
18 15 3 13 1 10 9 10 0 1 9 2 7 3 1 9 7 9 2
25 9 1 11 3 13 16 9 15 10 0 2 11 11 2 9 7 9 9 2 13 14 15 1 9 2
26 15 13 1 9 10 9 14 15 13 1 9 2 1 9 0 9 2 7 13 1 9 10 9 10 0 2
8 15 3 13 13 9 0 0 2
25 15 13 1 10 9 2 16 7 15 13 9 1 9 7 15 0 9 2 2 4 13 7 13 2 2
16 15 13 1 9 1 9 15 1 9 0 1 9 2 9 0 2
22 15 13 13 14 9 15 14 11 1 10 13 2 7 13 1 15 1 9 15 9 2 2
27 9 0 13 1 9 0 2 3 13 13 9 2 11 13 16 13 9 1 9 1 9 0 14 9 15 2 2
23 9 15 10 0 14 11 1 10 9 13 7 13 2 7 10 9 13 1 9 14 9 15 2
6 15 13 1 11 13 2
4 15 3 13 2
26 1 11 13 1 9 15 11 14 10 9 10 0 10 0 3 16 13 3 2 3 1 9 1 9 11 2
36 9 0 2 11 11 2 9 10 9 3 14 11 11 2 9 2 9 2 13 1 9 0 1 10 9 1 9 11 2 10 9 1 9 10 9 2
20 9 0 2 11 11 2 13 14 9 10 9 1 9 11 1 9 9 9 12 2
26 9 12 2 11 11 2 9 0 2 13 12 9 9 1 9 11 2 7 3 13 14 15 1 9 0 2
15 9 13 2 7 13 1 9 1 9 11 7 1 9 11 2
17 1 9 9 13 7 1 11 10 0 12 9 1 11 7 12 9 2
11 10 9 12 3 13 13 3 1 10 9 2
9 1 15 13 9 10 9 10 0 2
15 1 10 9 13 12 9 2 7 3 1 15 13 12 9 2
30 12 1 15 2 11 11 2 0 1 9 11 2 13 1 10 9 2 7 14 9 15 13 9 0 1 11 2 11 11 2
18 9 15 14 11 13 9 0 1 12 10 9 10 0 14 9 10 9 2
24 11 13 13 9 1 11 13 1 11 2 7 3 15 9 0 2 7 9 15 13 13 1 9 2
25 9 0 1 11 13 1 9 11 16 10 9 1 9 15 10 0 14 11 13 9 0 1 9 11 2
11 1 10 9 13 11 1 9 14 12 9 2
7 1 12 9 13 10 9 2
31 1 9 10 9 2 1 16 13 1 9 15 2 13 11 1 9 9 7 13 14 10 9 1 9 15 1 9 14 9 0 2
13 15 3 13 16 13 9 0 1 9 15 14 15 2
23 11 2 9 1 9 10 9 1 9 0 2 13 13 9 9 0 1 11 1 9 9 0 2
13 9 10 9 14 15 13 1 10 0 3 1 11 2
7 12 1 15 13 9 0 2
21 1 12 13 11 13 14 11 11 1 9 10 11 2 1 9 13 1 15 9 0 2
37 1 10 9 15 13 13 1 9 0 1 9 9 9 1 9 15 2 7 13 16 13 1 15 9 13 1 9 1 16 9 10 9 14 15 13 13 2
9 11 3 13 1 9 1 10 15 2
13 15 3 2 9 2 16 4 3 13 1 15 9 2
18 3 1 15 2 1 9 9 15 1 9 13 13 9 14 12 12 9 2
16 11 13 10 9 10 0 1 10 9 3 16 13 13 9 13 2
27 2 9 10 9 2 13 3 10 3 0 2 1 16 1 10 9 3 13 10 9 10 0 13 7 9 0 2
24 9 7 9 9 9 13 14 10 9 1 13 9 0 14 9 2 7 13 1 15 10 9 0 2
31 0 2 1 9 9 2 9 15 14 10 9 11 1 9 0 3 2 16 1 9 15 9 15 14 11 1 9 13 9 0 2
31 9 0 0 1 9 15 2 11 11 11 2 3 16 13 10 9 10 0 1 9 10 9 2 13 1 9 15 1 9 15 2
23 3 1 9 15 13 1 10 9 2 7 10 9 3 13 1 15 13 1 9 0 1 11 2
36 1 12 13 1 9 0 1 10 9 2 11 2 2 16 3 1 11 13 10 9 1 13 2 7 3 1 9 9 2 9 2 7 1 9 9 2
8 15 13 1 10 9 1 11 2
29 15 3 13 14 10 9 10 0 1 9 0 2 7 9 11 3 13 16 13 1 9 15 1 9 9 15 1 9 2
34 12 9 0 2 13 1 15 14 11 11 2 13 7 15 3 1 9 0 0 16 13 9 0 2 15 14 11 11 7 15 14 11 11 2
26 11 2 16 3 13 9 1 9 11 1 9 10 9 2 13 1 9 10 9 1 10 9 1 11 12 2
15 1 10 9 2 1 9 12 2 15 13 9 1 9 11 2
18 3 3 13 9 1 9 11 9 1 9 9 15 14 11 11 2 11 2
28 1 12 2 1 9 0 2 13 16 13 9 13 1 15 9 9 1 9 1 9 15 14 9 1 9 10 9 2
15 1 12 13 1 15 9 2 9 16 13 1 15 9 0 2
15 1 3 13 9 15 1 9 0 14 9 1 9 2 9 2
21 1 10 9 1 9 10 9 1 11 2 11 11 2 13 3 9 15 14 11 11 2
54 15 13 1 9 10 9 10 0 10 0 1 9 1 11 2 13 9 0 1 10 9 14 10 9 1 9 9 7 9 2 13 13 2 13 14 9 15 2 7 13 1 9 15 1 10 13 14 10 1 9 15 1 9 2
7 1 10 9 13 9 15 2
15 9 9 1 11 13 14 15 1 10 9 3 1 9 15 2
41 1 9 12 13 9 0 16 1 11 12 13 1 15 10 9 11 11 9 2 7 16 1 10 10 9 13 10 9 1 9 9 10 9 10 0 1 11 7 1 11 2
14 1 9 12 13 10 9 1 11 2 7 15 3 13 2
22 1 11 12 13 1 9 0 9 1 9 15 3 2 7 7 13 2 9 9 15 2 2
8 7 3 13 1 11 10 0 2
13 13 9 16 9 11 13 3 14 9 11 7 11 2
48 1 9 9 16 13 1 10 12 1 11 3 1 11 13 9 10 9 1 9 10 9 2 9 11 11 2 1 2 9 10 9 10 0 13 1 9 14 12 10 9 14 11 2 11 7 11 2 2
12 15 13 2 2 12 9 15 13 1 9 0 2
13 3 15 9 16 12 10 9 15 3 13 1 3 2
21 9 15 13 9 0 7 9 9 1 10 9 2 1 10 9 7 1 9 10 9 2
10 15 13 16 15 13 1 9 0 0 2
31 3 13 1 9 9 7 9 1 10 9 2 16 16 15 0 1 9 14 9 16 13 13 16 13 14 10 9 10 0 2 2
4 7 3 3 2
7 11 2 11 7 11 0 2
9 10 12 1 15 13 1 9 12 2
14 10 9 13 16 10 9 10 0 13 16 13 1 9 2
15 3 16 0 2 16 15 13 4 1 9 15 1 10 9 2
30 15 13 1 9 9 16 0 1 9 2 1 9 0 2 7 1 9 16 4 13 9 16 0 9 3 0 1 9 0 2
35 12 7 9 9 13 3 1 11 12 12 1 9 15 14 11 11 1 9 9 0 2 0 9 9 1 9 1 9 2 1 9 7 1 9 2
33 1 9 12 2 14 13 10 9 13 2 13 10 9 12 9 0 2 12 1 15 3 2 7 12 9 13 2 9 16 13 7 15 2
13 1 9 12 3 13 9 10 12 1 9 7 9 2
19 1 1 9 10 9 13 12 1 9 10 9 10 0 1 9 11 10 9 2
13 9 9 11 13 1 9 16 13 1 9 10 9 2
9 9 9 0 13 1 9 9 0 2
8 9 9 0 13 1 9 9 2
10 1 9 12 13 10 9 1 10 9 2
18 1 10 9 13 9 15 14 12 1 9 10 9 2 16 13 9 11 2
8 10 9 13 1 15 1 9 2
17 9 10 12 13 9 0 2 9 2 9 0 1 11 7 9 9 2
17 9 10 9 11 13 13 14 9 10 9 1 10 9 1 10 9 2
13 3 1 9 9 15 13 13 15 2 7 1 9 2
39 9 10 9 2 10 9 2 9 11 7 3 10 9 10 0 1 11 2 10 11 1 11 10 9 11 11 2 13 1 9 10 9 13 10 9 2 7 3 2
27 12 13 1 9 10 9 11 2 1 16 15 13 9 14 9 7 13 9 7 9 1 9 10 9 10 0 2
23 10 9 11 11 7 9 15 11 11 2 16 13 13 14 10 9 11 2 13 1 10 9 2
34 1 10 9 13 9 10 11 11 11 2 10 9 11 11 2 10 9 3 11 11 11 2 9 11 11 7 9 0 0 1 9 10 9 2
16 1 12 13 9 10 9 11 13 1 9 14 16 13 1 15 2
7 10 9 2 9 16 13 2
24 1 9 9 10 9 16 13 1 15 1 9 10 13 2 13 10 9 10 0 14 9 10 9 2
44 10 9 10 0 13 1 9 15 14 11 2 2 10 9 14 15 2 10 9 14 15 7 9 10 9 14 15 2 2 7 1 15 13 1 10 9 2 2 10 11 13 9 15 2
7 3 13 1 9 10 9 2
8 13 14 10 9 1 9 2 2
32 10 9 11 11 2 9 15 14 11 11 2 13 1 10 9 1 9 2 16 2 9 15 14 11 13 1 9 9 2 10 9 2
6 10 9 10 15 13 2
9 1 10 9 10 15 13 9 2 2
43 3 1 9 15 14 10 9 11 11 2 9 1 9 10 9 10 0 7 9 12 1 9 11 1 10 11 2 13 3 9 0 2 2 9 13 9 15 7 15 13 14 15 2
4 9 9 10 2
4 3 9 13 2
7 15 10 9 13 9 15 2
16 13 1 9 2 7 13 4 13 1 9 2 3 1 10 9 2
23 9 1 9 7 9 1 9 2 13 4 13 1 10 9 2 7 15 3 13 14 10 9 2
4 15 10 9 2
11 15 10 9 13 9 15 14 10 9 2 2
44 9 15 14 11 11 2 11 2 9 11 16 0 3 1 10 9 11 2 13 10 0 3 2 7 15 13 1 9 15 2 7 3 13 13 2 2 10 9 11 13 14 15 9 2
14 3 1 10 9 13 14 15 7 1 11 13 14 15 2
11 10 9 10 0 13 13 14 15 9 12 2
15 13 7 13 13 7 13 14 10 9 16 13 14 15 9 2
16 13 14 9 10 9 1 10 9 3 2 9 1 10 9 9 2
6 9 10 9 11 2 2
18 3 3 13 10 9 13 1 1 9 1 10 9 1 10 9 10 0 2
31 3 1 9 7 1 15 1 9 13 7 13 2 2 9 1 10 9 2 2 2 9 1 10 9 2 2 2 13 9 2 2
13 10 9 10 15 13 0 1 9 7 15 13 9 2
17 3 3 1 3 13 9 14 10 12 3 16 13 13 16 13 9 2
5 7 10 9 0 2
16 9 9 0 1 9 10 9 13 14 9 15 1 9 7 9 2
17 12 1 15 13 9 7 13 1 1 10 9 2 1 9 13 9 2
8 3 13 12 1 9 10 9 2
7 9 9 13 14 15 3 2
8 9 13 1 9 1 9 15 2
19 9 0 14 9 13 1 10 9 10 0 9 12 2 1 10 9 10 0 2
6 9 9 10 9 13 2
8 9 1 9 15 13 1 9 2
12 3 1 15 13 9 9 14 9 1 10 9 2
8 10 9 13 3 1 10 9 2
17 1 9 9 12 1 9 9 11 15 9 1 10 9 10 0 3 2
