2595 11
5 11 11 11 11 11
8 9 9 13 11 13 9 11 2
13 11 13 0 11 11 11 7 13 0 9 0 9 2
9 13 3 9 9 1 3 1 12 2
14 9 15 1 13 12 9 2 15 1 13 3 1 9 2
16 13 11 7 11 1 0 9 13 2 7 3 9 13 0 9 2
13 3 11 7 11 13 9 2 7 15 13 3 9 2
15 0 3 13 2 16 9 13 11 13 3 0 9 9 1 2
8 2 15 13 2 15 13 2 2
5 3 13 9 13 2
6 13 3 0 13 9 2
17 9 13 11 11 9 7 3 15 9 7 9 9 13 9 13 15 2
8 15 0 9 13 3 13 13 2
16 0 9 15 0 9 13 3 0 3 13 2 7 13 3 13 2
20 0 9 9 13 0 9 2 3 3 4 3 13 2 15 9 13 15 15 0 2
5 9 13 15 0 2
10 15 9 13 15 0 7 0 0 9 2
13 15 9 13 3 4 13 15 2 7 3 13 3 2
18 15 13 9 13 2 16 9 13 3 0 0 9 2 16 15 13 0 2
18 9 13 13 9 9 13 2 7 13 2 16 15 3 9 13 9 2 5
11 11 2 11 7 11 13 1 9 3 13 2
15 9 4 13 11 0 9 7 3 15 9 2 15 11 13 2
18 0 2 3 3 13 13 9 15 9 9 7 13 2 15 13 9 15 2
10 13 3 13 0 9 7 13 15 0 2
11 13 3 0 2 16 3 13 13 15 2 5
8 11 1 13 13 9 15 9 2
13 0 9 3 13 15 1 7 3 13 15 0 9 2
7 11 13 3 9 13 2 5
13 0 9 13 15 0 9 7 13 9 9 9 1 2
9 15 3 9 9 7 3 0 9 2
16 15 13 4 13 15 16 2 16 2 2 11 13 15 9 2 2
15 13 15 3 0 7 0 3 2 7 15 0 9 13 2 5
17 15 9 13 3 9 2 7 0 9 3 3 13 11 13 9 1 2
19 13 13 13 9 3 3 2 16 15 2 11 7 11 4 13 9 9 13 2
9 13 3 13 9 15 9 0 9 2
9 3 2 13 15 0 9 3 3 2
4 13 13 0 2
9 9 7 9 13 0 9 13 9 2
7 9 15 7 9 9 11 2
6 3 0 9 13 3 5
10 11 2 11 7 11 13 9 15 9 2
17 0 9 13 11 9 15 0 0 2 7 3 13 3 0 9 2 5
7 4 3 3 13 9 3 2
12 12 9 13 13 15 2 7 3 15 3 13 2
17 13 13 3 3 2 9 1 2 9 2 9 7 0 9 13 9 2
9 9 13 0 7 15 13 0 9 2
7 9 13 0 9 0 9 2
12 9 4 13 12 5 0 9 7 9 13 9 2
16 3 11 9 13 3 9 2 16 4 15 1 13 3 9 2 5
9 11 3 13 3 3 15 9 9 2
7 9 4 13 9 9 2 5
21 0 9 9 13 3 11 11 11 7 15 13 13 13 11 9 2 16 3 9 13 2
21 9 13 3 15 0 9 15 2 16 15 9 4 13 9 13 9 7 9 7 9 2
3 3 0 2
5 15 9 0 9 2
11 3 13 13 11 9 7 13 9 3 9 2
18 3 16 13 15 3 9 1 2 9 4 13 3 0 13 0 7 0 2
9 13 3 3 3 9 7 9 2 5
14 13 3 13 3 0 3 9 2 16 15 4 3 13 2
3 3 13 2
7 8 8 8 9 2 11 2
28 16 13 15 0 11 13 9 13 2 9 13 13 8 2 8 8 8 2 13 15 3 2 9 7 13 9 9 2
20 4 13 9 9 2 15 13 9 7 13 3 3 13 3 13 9 7 13 9 2
29 13 3 2 16 13 13 3 0 11 13 8 8 9 2 7 9 13 13 15 9 1 3 2 3 15 13 13 9 2
4 9 9 3 2
29 0 9 13 3 3 3 9 2 16 13 4 13 13 2 13 13 9 3 2 7 9 7 9 2 11 7 3 3 2
32 15 3 13 15 2 16 13 11 9 7 9 9 7 9 0 9 9 7 3 9 2 7 9 0 9 2 2 3 9 13 9 2
21 0 9 13 15 0 9 2 16 13 13 3 0 9 16 13 7 9 13 3 8 2
33 15 13 3 9 2 16 15 13 13 0 9 2 13 0 9 2 7 15 13 3 9 13 13 0 8 15 2 2 15 13 13 9 2
12 3 3 13 3 9 2 15 11 13 0 9 2
15 13 3 13 13 3 12 9 9 2 3 9 13 0 9 2
18 3 13 15 9 13 3 16 9 13 2 3 9 13 4 3 0 13 2
28 3 3 15 9 7 3 3 3 3 2 16 4 13 13 15 9 8 0 13 2 3 13 3 12 9 12 1 2
5 12 9 13 3 2
22 0 9 13 3 15 9 2 15 4 13 3 15 16 13 13 13 0 9 9 9 15 2
9 9 3 13 2 3 15 9 13 2
24 15 9 4 13 15 1 3 12 9 9 2 13 9 2 16 9 13 9 13 0 15 9 2 2
17 0 9 13 3 3 3 12 9 2 16 9 13 3 15 8 9 2
6 7 15 13 0 8 2
10 0 15 4 13 4 13 3 12 9 2
17 9 13 15 9 15 4 13 15 2 15 13 9 3 12 9 1 5
5 9 16 9 13 2
6 11 13 11 3 3 2
10 3 12 9 2 15 13 3 12 2 2
4 9 13 9 2
2 9 2
13 13 9 9 9 2 13 13 11 9 15 9 13 2
6 11 9 2 15 13 2
10 9 9 13 9 16 13 15 3 13 5
4 9 7 15 9
19 13 3 15 9 1 2 16 9 13 13 11 9 7 13 13 3 8 9 2
15 9 4 3 3 13 7 2 13 2 2 16 11 9 13 2
12 3 9 4 13 15 9 2 7 13 9 9 2
11 9 15 2 3 15 4 13 2 13 13 2
17 15 4 13 3 0 0 8 7 15 15 2 15 11 9 13 9 2
7 3 9 13 11 11 11 2
8 3 3 13 2 4 15 13 2
11 13 11 9 7 13 9 9 2 5 2 2
11 16 9 13 13 2 15 4 13 11 9 2
5 9 4 3 13 2
4 13 0 9 2
14 0 13 9 5 7 13 0 8 2 5 9 2 9 2
11 0 13 9 2 8 8 8 8 8 8 2
10 0 13 2 16 11 9 13 7 13 9
15 0 8 13 9 9 1 13 2 3 13 9 9 0 8 2
2 9 2
5 15 13 3 0 5
18 16 0 9 9 4 13 3 0 2 3 15 9 13 0 7 0 9 2
13 3 12 13 11 7 9 13 9 7 15 0 9 2
15 15 9 9 13 11 2 6 6 6 2 2 7 11 11 2
24 3 13 11 11 2 11 2 7 13 11 9 0 9 2 15 3 9 13 9 11 7 0 9 2
24 7 13 3 13 3 3 9 7 0 9 2 3 9 13 11 7 11 1 9 11 13 3 11 2
17 15 9 0 9 4 13 9 2 15 9 13 3 3 4 13 15 2
8 3 2 16 9 3 13 9 2
15 9 0 7 0 9 13 9 9 7 9 9 2 0 15 2
8 0 9 4 3 13 0 9 2
11 15 9 13 3 13 9 9 7 0 9 2
2 0 2
2 3 2
10 7 3 3 13 15 0 9 9 13 2
9 13 3 0 9 7 0 9 13 2
13 3 3 3 2 16 3 13 15 2 13 13 15 2
13 7 16 9 13 13 13 0 9 2 13 3 15 2
8 6 6 2 13 0 9 13 2
12 4 15 9 3 3 3 13 15 11 2 9 2
10 13 15 13 3 12 9 0 9 13 2
2 13 9
12 15 9 9 9 3 9 7 9 13 13 9 2
31 9 13 3 3 13 9 2 16 15 13 0 9 3 9 7 9 2 15 4 13 0 9 3 9 2 9 7 3 9 3 2
15 13 9 4 3 13 0 9 0 7 15 4 13 3 15 2
15 13 9 13 13 3 13 2 16 9 9 13 3 15 9 2
13 13 9 3 9 3 7 3 3 0 9 0 9 2
9 13 9 9 7 13 15 3 9 2
10 13 3 9 0 9 7 13 15 3 2
6 9 13 3 15 9 2
6 13 2 13 13 9 2
10 13 9 7 13 3 9 7 0 9 2
3 13 9 2
13 13 9 13 0 3 0 9 2 3 0 0 15 13
11 15 9 13 13 9 0 9 7 9 1 2
8 13 9 13 3 9 9 2 2
16 15 13 3 12 9 13 9 7 9 13 15 0 9 7 9 2
13 13 9 13 3 3 9 2 9 7 3 9 9 2
1 13
19 0 9 2 9 9 13 9 9 13 0 9 9 12 9 2 15 13 11 2
13 3 13 0 9 2 16 15 13 15 9 3 0 2
7 9 9 13 3 9 9 2
18 15 13 0 2 16 9 9 13 0 9 15 9 16 9 13 9 9 2
15 13 3 0 2 16 9 9 13 15 9 16 9 13 9 2
11 9 0 9 13 9 7 9 0 9 3 2
10 15 9 4 13 0 9 9 9 9 2
9 9 13 13 9 9 3 12 9 2
11 9 13 15 3 13 9 12 9 9 9 2
17 16 15 13 13 9 9 2 9 13 15 9 3 13 9 9 9 2
6 15 9 13 9 9 2
11 9 9 13 3 3 0 9 7 9 9 2
9 15 9 1 0 9 13 0 9 2
8 0 11 13 12 12 9 9 2
12 3 11 9 13 9 13 3 12 12 9 9 2
8 15 4 13 0 9 11 9 2
9 3 2 9 9 9 13 15 9 2
13 15 13 15 2 16 9 9 13 0 9 9 9 2
7 3 0 9 13 15 9 2
34 0 9 2 13 3 15 9 2 16 15 13 13 15 9 9 2 16 13 13 15 13 9 0 9 2 15 13 9 9 7 12 9 3 2
33 16 9 13 3 0 2 7 9 9 13 0 2 13 9 9 2 16 9 9 2 7 15 7 9 11 2 13 13 0 9 15 9 2
18 13 2 16 13 9 1 13 9 15 9 0 9 2 7 3 12 9 2
6 0 9 9 4 13 2
3 13 13 2
39 0 9 2 0 9 9 2 0 9 7 9 2 15 13 15 0 0 9 2 7 15 15 2 15 3 13 2 13 2 7 13 15 3 3 9 9 2 9 2
14 13 15 3 3 13 2 16 13 13 9 13 0 9 2
26 13 3 13 9 11 15 2 7 13 3 3 13 12 9 15 9 2 3 12 9 2 15 13 9 12 2
31 11 9 13 9 15 9 9 2 16 11 9 9 9 13 9 9 9 13 0 9 9 13 0 9 2 15 13 15 9 9 2
17 0 9 9 7 9 13 3 15 9 2 16 0 9 4 13 9 2
9 0 9 9 7 9 13 9 9 2
7 3 9 13 9 9 9 2
40 13 15 13 15 2 16 0 9 1 2 15 13 9 7 9 9 9 2 15 15 9 7 15 9 13 9 13 3 15 9 2 3 15 0 9 13 9 9 1 2
14 13 13 2 16 13 13 9 13 9 1 13 15 9 2
20 9 12 0 9 13 9 0 9 9 9 7 9 9 7 9 9 13 9 1 2
23 9 13 15 2 13 0 9 9 9 12 9 2 9 2 7 12 9 9 2 9 9 2 2
22 15 9 13 0 11 9 9 9 9 3 15 2 16 9 9 12 9 13 0 0 9 2
30 9 9 9 0 13 9 9 7 9 9 4 13 9 0 9 9 2 16 9 9 12 9 7 12 9 9 13 13 9 2
23 0 9 9 9 13 13 13 9 0 9 9 2 3 9 7 9 7 9 7 9 9 9 2
10 9 13 9 9 4 9 9 13 9 2
11 3 11 9 9 13 3 13 0 9 9 2
23 3 13 9 9 9 9 9 13 9 3 13 4 3 13 0 9 13 9 7 15 13 9 2
24 4 3 13 2 16 9 15 9 13 15 9 3 2 13 13 2 16 15 9 1 13 0 9 2
1 9
11 15 13 15 9 2 15 9 2 15 9 2
10 15 13 15 9 7 15 9 13 15 2
9 9 13 11 9 15 13 16 9 2
16 13 2 3 13 13 15 15 1 2 13 2 16 15 13 9 2
12 9 13 9 9 7 13 2 16 15 13 3 2
18 13 0 9 2 13 13 15 9 2 13 9 9 2 9 9 7 15 2
16 13 9 7 13 9 2 15 9 13 9 7 9 13 9 9 2
10 13 9 9 2 3 9 13 0 9 2
12 9 13 0 9 2 13 15 2 13 3 15 2
8 15 9 13 13 15 0 9 2
6 13 3 7 13 3 2
9 9 13 9 7 15 9 13 9 2
14 15 13 9 2 9 7 3 13 13 15 3 0 9 2
1 9
6 9 15 13 9 9 2
9 3 0 9 1 3 0 2 0 2
25 9 2 15 9 13 9 7 15 4 13 9 2 13 9 7 9 9 9 2 13 9 13 9 3 2
15 9 13 9 2 9 2 9 0 9 7 0 0 0 9 2
15 15 13 15 9 7 9 2 15 13 9 15 9 7 9 2
9 15 13 0 2 0 7 0 9 2
10 15 9 9 4 13 0 9 9 1 2
19 9 15 13 2 16 13 3 3 13 0 9 2 3 9 13 3 0 9 2
4 9 13 13 2
12 4 3 13 3 2 15 9 4 13 12 9 2
12 13 15 13 9 3 2 7 9 13 9 13 2
16 3 15 9 13 2 7 3 15 13 3 0 2 0 9 1 2
9 13 0 9 2 13 15 13 3 2
13 0 7 9 13 9 9 7 9 4 13 0 9 2
5 3 3 13 9 2
10 13 9 2 15 9 13 15 9 3 2
7 16 13 2 13 9 3 2
7 13 3 2 3 16 13 2
28 13 3 13 9 15 2 7 9 13 9 1 9 0 9 2 3 9 13 2 3 0 9 13 13 0 9 9 2
14 16 4 13 15 1 9 2 13 9 9 13 3 15 2
2 1 9
15 0 9 13 2 16 15 3 13 2 16 15 9 13 3 2
6 15 4 13 3 3 2
8 13 15 2 16 9 13 3 2
8 15 9 13 3 3 3 13 2
10 4 15 3 13 13 2 16 9 13 2
12 13 2 16 16 9 13 13 9 2 15 13 2
14 13 13 9 2 16 16 9 13 13 2 15 13 3 2
7 13 3 2 16 9 13 2
13 15 13 3 15 9 2 16 15 9 13 9 1 2
9 6 15 9 13 3 9 13 13 2
21 0 15 13 2 16 15 13 0 9 2 16 9 13 3 3 3 3 0 9 3 2
4 15 4 13 2
4 15 13 0 2
4 9 13 13 2
15 16 9 13 2 13 0 2 16 6 2 3 15 4 13 2
19 16 13 9 7 15 3 9 13 9 13 15 13 3 15 13 0 9 9 2
50 16 13 9 0 9 7 9 2 16 13 9 7 9 9 13 2 13 13 9 2 16 13 9 0 9 9 1 2 3 15 4 13 13 9 9 2 9 9 2 0 9 2 9 2 9 9 2 9 9 2
6 15 13 0 9 0 2
40 16 9 3 13 3 7 15 15 13 2 13 3 2 3 15 15 13 2 7 2 13 13 2 3 16 9 13 9 4 13 13 13 9 7 13 3 9 0 9 2
7 13 15 15 9 3 0 2
13 13 15 9 0 13 9 3 0 7 0 9 13 2
9 4 15 13 3 2 3 2 3 2
9 13 9 0 13 9 1 9 9 2
3 3 13 2
3 13 13 2
10 3 13 3 9 2 9 7 3 9 2
20 3 12 9 1 13 9 7 15 13 9 13 2 16 13 15 9 3 9 13 2
10 7 3 9 13 3 9 2 3 9 2
11 13 13 2 7 15 13 2 16 15 13 2
2 0 9
6 13 13 9 9 9 2
12 0 9 9 13 4 4 0 9 13 9 9 2
9 3 13 7 0 9 9 7 3 2
14 3 0 9 13 9 9 2 16 0 9 13 3 3 2
15 3 3 4 13 3 3 0 9 9 7 0 9 15 9 2
12 3 13 0 13 0 9 13 9 13 9 9 2
12 3 13 0 13 9 1 9 9 7 15 9 2
13 3 9 9 13 3 9 16 15 9 4 13 3 2
21 16 9 13 9 7 15 1 0 9 9 1 2 13 13 0 9 2 15 13 9 2
7 15 3 3 13 13 9 2
8 15 4 13 3 13 13 9 2
7 3 15 3 13 13 9 2
14 9 3 13 13 9 1 7 3 9 15 0 13 9 2
7 13 0 16 9 13 9 2
5 9 13 13 3 2
16 15 0 9 13 4 13 13 15 9 7 9 9 1 15 9 2
16 9 13 3 15 13 9 9 3 13 7 3 0 9 13 9 2
17 0 0 9 13 3 15 2 16 9 13 3 9 7 15 9 9 2
16 3 4 3 3 13 15 0 9 13 13 3 3 3 13 9 2
17 3 13 9 13 3 9 4 9 13 15 3 16 9 13 9 15 2
10 9 13 0 9 0 7 0 9 9 2
12 0 9 0 0 0 9 9 13 9 13 13 2
16 15 1 9 9 13 3 0 0 7 0 9 13 9 13 9 2
5 3 9 3 13 2
6 13 15 3 1 9 2
11 3 3 15 13 9 2 1 9 7 9 2
6 15 13 0 9 9 2
5 13 15 12 9 2
14 7 0 15 13 2 16 13 3 13 2 16 13 9 2
9 15 13 9 9 13 0 9 3 2
12 13 3 2 16 4 3 13 9 7 13 9 2
15 11 4 13 11 3 12 9 12 9 2 16 15 13 9 2
13 11 1 11 13 15 9 7 13 9 3 0 9 2
2 2 13
5 11 13 11 9 2
9 15 13 9 2 15 13 15 0 2
7 9 9 13 13 13 9 2
13 9 15 4 3 13 2 13 3 9 7 0 9 2
4 15 4 13 9
8 0 9 4 13 9 7 9 2
9 11 13 15 9 2 15 4 13 2
3 0 13 2
15 11 9 13 3 12 5 9 2 16 15 11 13 12 5 2
3 3 0 9
2 3 2
10 3 13 3 3 9 7 9 13 13 2
8 13 0 9 13 9 9 3 2
2 13 0
7 15 13 9 9 13 9 2
18 13 3 3 3 2 13 15 3 11 2 15 9 4 13 2 13 11 2
2 9 13
8 3 13 3 13 13 9 3 3
19 9 13 2 16 9 7 9 13 3 15 2 15 13 3 12 12 9 9 2
6 7 3 15 15 13 2
2 13 9
5 0 9 3 9 2
8 15 13 16 13 13 15 15 2
7 11 13 13 9 3 3 2
9 13 15 3 2 3 13 0 9 2
2 0 9
20 3 0 9 3 13 9 9 11 11 13 9 13 13 15 0 9 11 11 9 2
7 9 9 13 0 16 9 2
5 9 4 13 2 2
9 9 13 13 16 13 15 13 9 2
6 3 9 13 3 3 2
6 15 13 15 3 13 2
11 3 15 3 13 2 16 9 13 13 13 2
8 11 11 9 13 0 0 9 2
5 15 13 9 9 2
9 15 9 9 13 13 13 1 9 2
5 9 13 9 0 2
12 16 12 9 13 2 3 15 13 15 3 11 9
7 9 13 15 2 16 13 2
9 9 9 9 13 9 12 12 9 2
4 9 13 0 2
8 15 13 3 13 13 13 13 9
8 9 4 13 13 0 9 9 2
4 2 3 0 2
6 11 13 3 9 0 9
7 15 9 9 13 3 11 2
7 11 9 9 11 11 1 2
6 9 9 9 9 13 2
11 15 13 0 9 16 13 0 2 15 13 2
4 9 13 6 2
13 9 13 3 9 2 15 9 13 11 11 7 9 2
7 9 7 9 9 11 13 9
7 11 13 9 7 15 13 2
6 13 15 9 2 11 2
10 9 13 3 0 2 16 13 3 0 2
4 9 7 9 9
2 13 13
11 15 13 9 7 13 9 13 2 0 9 2
3 9 13 9
2 0 9
2 9 11
5 15 13 9 0 2
11 16 15 4 13 9 3 2 4 13 15 9
5 3 9 9 13 2
10 15 15 13 2 15 13 0 9 3 2
17 4 13 3 0 0 2 7 15 13 3 13 3 0 9 16 11 2
13 9 13 9 7 13 2 16 9 13 3 9 13 2
7 15 13 9 9 3 6 2
9 2 15 3 2 15 13 4 13 2
12 13 13 9 9 13 9 9 9 7 13 11 2
7 13 15 11 15 9 3 2
6 15 4 13 9 0 2
12 9 13 13 15 15 2 15 3 13 13 9 2
7 15 13 2 16 9 13 2
9 15 15 13 13 2 16 13 9 2
2 9 9
7 15 13 3 9 15 3 2
4 13 15 9 2
7 9 1 9 4 13 11 2
45 16 3 15 13 3 9 7 3 15 13 16 3 13 3 3 15 16 6 16 15 3 13 3 15 0 9 3 3 15 13 3 16 6 16 16 3 15 3 13 16 4 15 13 15 9
7 13 3 9 9 1 1 2
9 16 13 13 2 13 9 3 13 2
7 3 3 11 13 0 9 2
2 13 13
9 0 9 13 9 7 0 0 9 2
11 13 2 16 11 9 13 9 12 12 9 2
8 3 13 9 13 9 3 13 2
2 13 15
6 13 3 3 12 9 2
8 15 13 0 9 13 9 9 2
5 3 9 13 11 2
6 15 4 13 0 9 2
15 13 15 9 3 2 13 13 3 2 7 13 15 9 3 2
2 13 13
5 15 4 13 12 9
10 3 9 12 9 13 11 3 12 12 2
4 3 13 0 9
7 9 13 0 16 9 0 2
18 15 11 9 3 15 13 3 0 16 15 13 16 15 3 13 15 9 2
13 16 11 9 13 11 2 11 1 0 9 13 13 2
6 9 13 7 9 13 2
6 9 9 4 13 0 2
6 15 13 15 3 3 2
16 11 13 9 4 3 3 13 2 16 13 15 13 13 0 9 2
6 9 11 9 12 1 2
7 15 4 13 0 9 9 2
10 9 9 13 0 9 7 9 11 11 2
7 13 13 3 13 0 9 2
7 9 0 9 13 15 3 2
6 0 13 3 0 9 2
29 11 11 7 15 9 13 15 0 15 13 13 9 9 2 7 13 15 13 7 13 2 16 15 13 9 0 0 9 2
10 13 3 2 0 9 2 9 15 13 2
2 13 9
10 0 0 9 4 13 13 9 9 1 2
5 13 15 3 0 2
4 9 13 9 2
7 0 9 11 4 13 9 2
5 4 13 3 9 2
16 13 9 13 9 0 9 3 7 9 13 0 0 2 3 13 2
13 15 13 13 15 9 15 13 9 9 0 9 9 2
5 6 6 15 1 2
6 15 0 9 13 9 2
10 3 9 9 3 15 13 15 9 9 2
5 13 15 3 6 2
10 13 15 9 9 9 0 9 12 9 1
3 13 3 2
7 11 13 11 0 0 9 2
5 13 9 0 9 2
4 13 15 9 2
9 3 15 4 13 12 0 0 9 2
4 15 15 13 13
2 11 9
16 11 11 2 15 9 13 3 0 9 15 11 9 13 15 9 2
12 15 15 15 0 9 4 13 13 3 9 9 2
13 9 4 4 13 3 15 9 16 15 13 9 7 2
8 9 11 13 9 11 0 9 2
9 11 13 2 15 13 9 9 9 2
6 15 0 15 3 13 2
5 11 13 3 13 9
8 9 13 9 13 3 15 9 2
16 9 9 12 2 13 12 9 9 12 2 9 7 9 13 9 9
177 11 9 9 2 15 13 9 11 9 9 7 3 15 12 9 2 13 9 9 9 2 12 2 2 13 9 9 9 2 12 2 2 7 13 2 16 9 9 0 9 9 9 1 12 9 9 12 13 9 9 12 2 12 2 7 9 7 9 9 0 2 0 0 9 7 9 9 9 9 1 12 9 9 12 13 9 9 12 2 12 2 13 2 16 9 13 7 13 9 13 0 9 2 0 9 7 9 9 0 9 9 9 4 4 3 13 9 7 9 13 9 2 0 9 13 4 13 15 9 2 15 1 4 13 0 9 0 9 7 9 13 9 9 9 7 9 13 9 9 9 9 3 2 4 13 15 2 16 0 9 9 13 9 13 9 7 9 13 3 15 9 13 9 13 9 2 7 4 13 0 9 0 7 0 9 9 2
5 4 13 15 9 2
16 12 9 15 9 13 9 2 15 13 9 13 9 13 9 9 2
2 12 9
5 0 15 9 13 2
20 2 9 13 9 2 2 9 12 9 9 7 9 12 9 9 7 9 13 9 2
33 2 9 13 9 2 2 9 7 2 16 9 13 9 3 13 2 15 3 15 9 2 15 0 9 4 13 9 13 9 13 9 9 2
19 0 3 12 9 13 9 1 13 13 9 9 12 7 12 12 9 13 9 2
2 12 9
62 0 9 4 13 15 2 16 9 13 9 13 0 9 13 9 9 15 9 7 9 9 2 15 15 4 13 9 7 16 15 13 3 3 3 9 9 7 9 13 9 7 16 3 2 15 9 2 9 7 9 9 7 9 2 15 9 4 13 1 9 9 2
22 0 9 13 9 13 13 13 9 9 2 15 15 13 3 13 7 15 15 13 4 13 2
32 0 9 13 9 13 13 13 0 7 0 9 13 0 9 7 9 13 9 2 15 15 13 4 13 7 15 13 3 13 15 9 2
20 16 9 13 15 9 7 9 9 2 9 13 9 4 13 0 9 3 1 9 2
69 0 15 9 13 13 9 13 9 0 9 2 15 9 2 0 9 13 2 13 9 9 13 9 4 13 0 15 9 12 9 3 2 3 16 15 4 13 15 9 9 2 7 9 2 4 13 9 1 2 3 13 9 13 7 9 9 9 15 9 2 15 15 13 9 13 9 1 0 2
16 0 15 9 9 13 0 0 9 4 13 12 9 13 9 3 2
2 12 9
13 0 0 9 4 13 15 13 9 9 9 9 9 2
59 15 4 3 13 15 2 16 15 13 9 13 9 13 9 2 9 2 15 13 15 9 7 15 2 16 15 13 13 0 0 0 9 15 9 7 9 2 15 15 13 9 7 9 7 9 2 15 9 13 3 2 9 2 0 15 13 9 9 2
25 0 9 4 13 3 12 9 13 9 13 9 7 3 12 9 0 9 2 3 16 9 9 4 13 2
33 0 15 0 9 4 13 13 9 7 15 13 9 0 9 7 13 15 2 16 15 15 9 13 9 4 13 9 13 9 13 9 9 2
2 12 9
32 0 9 4 13 9 7 13 13 0 9 0 7 3 0 9 9 9 7 9 13 9 0 9 13 13 9 0 9 7 9 9 2
36 0 0 9 4 13 0 9 7 9 7 13 0 9 15 15 9 13 0 7 0 9 9 9 2 13 3 13 9 13 9 9 7 13 15 9 2
13 15 9 4 13 9 13 9 9 0 9 9 9 2
72 3 2 16 9 9 13 9 2 16 9 13 9 4 3 13 0 9 2 0 9 4 13 15 13 13 0 9 2 16 0 9 13 4 13 9 2 9 2 16 0 9 7 9 4 13 0 9 7 13 0 9 2 0 9 4 13 15 13 13 0 9 2 16 15 9 7 9 13 4 13 9 2
17 0 9 4 13 15 2 16 0 9 7 9 3 13 13 0 9 2
2 12 9
41 9 13 9 13 9 9 13 9 7 9 7 0 9 1 13 9 3 13 9 9 15 2 16 0 9 9 13 9 13 9 7 9 13 3 15 9 13 9 13 9 2
40 16 9 7 9 7 9 12 7 12 13 9 13 3 2 16 0 9 9 13 9 13 4 13 15 9 2 4 13 9 7 15 9 15 9 12 9 13 9 13 2
2 12 9
25 16 13 15 9 13 9 2 9 12 2 12 2 13 0 9 13 9 9 12 12 9 13 9 3 2
2 12 9
22 9 13 9 1 12 9 9 12 9 2 15 4 13 9 0 0 0 9 7 9 9 2
6 9 13 15 9 9 2
2 12 9
21 0 9 4 13 15 9 9 13 9 2 9 7 0 9 3 3 12 9 9 12 2
7 15 4 13 15 9 13 2
20 15 9 13 9 4 13 15 9 7 15 4 13 0 9 2 16 15 3 13 2
9 9 4 13 15 2 3 9 13 2
21 0 9 4 13 9 0 0 0 9 2 15 15 4 13 7 13 15 9 13 9 2
2 12 9
7 15 9 4 13 15 9 2
7 13 11 12 9 9 12 2
5 9 1 11 11 9
6 11 13 2 9 1 9
19 0 9 9 13 11 13 9 9 0 9 15 2 3 9 9 9 13 9 2
18 9 9 7 9 13 13 3 3 2 13 0 9 4 9 13 9 13 2
19 9 0 7 0 9 13 3 0 9 2 15 13 0 9 16 0 9 9 2
12 3 2 0 9 13 9 7 9 13 3 0 2
5 13 9 7 9 2
34 9 3 13 9 9 9 2 9 13 13 15 9 0 3 3 3 2 3 16 4 13 15 9 2 13 9 7 3 13 3 9 13 9 2
18 16 9 13 9 9 0 9 2 13 0 9 9 0 9 7 15 9 2
16 0 9 13 13 13 13 3 12 9 0 9 15 3 13 9 2
4 9 2 9 9
7 9 13 15 9 9 9 2
15 9 2 15 3 13 2 13 9 7 9 13 9 13 9 2
10 9 13 0 2 7 3 0 4 13 2
14 9 9 13 15 13 2 13 3 3 13 13 2 15 2
19 11 0 9 13 3 9 13 9 15 2 3 9 9 4 13 9 3 9 2
25 11 9 9 2 15 13 13 3 9 13 9 2 13 3 0 9 9 2 15 13 9 9 3 3 2
9 15 13 4 13 9 13 9 9 2
27 9 9 13 9 13 0 2 0 9 3 9 9 13 13 0 3 16 0 9 9 7 9 13 9 9 9 2
14 9 13 3 4 13 9 9 9 2 16 15 13 13 2
2 9 9
16 16 9 13 0 13 2 13 15 9 3 13 3 15 9 9 2
9 9 9 13 3 0 9 7 9 2
8 9 1 9 13 13 3 0 2
22 9 2 15 9 9 3 13 0 9 2 13 15 3 13 9 7 9 13 3 15 9 2
20 9 1 13 3 13 15 3 9 2 7 9 4 13 0 0 2 16 9 13 2
8 15 9 11 9 13 13 13 2
31 9 1 13 3 9 2 16 9 13 15 9 2 15 13 13 2 15 4 13 15 3 13 4 9 2 3 9 13 0 9 2
7 9 9 9 13 3 15 2
13 9 7 9 13 3 13 2 16 9 4 13 3 2
13 0 0 9 15 9 13 9 2 15 13 9 0 2
17 9 13 3 9 9 13 9 2 16 3 13 9 9 7 9 3 2
19 9 15 13 3 13 2 3 4 13 7 13 9 3 9 2 9 7 9 2
14 3 9 1 9 1 13 15 2 13 3 9 13 15 2
9 3 15 13 13 13 9 9 9 2
7 15 0 9 13 9 9 2
17 15 9 13 9 9 7 15 15 9 2 15 9 9 13 9 1 2
13 15 13 3 0 9 2 15 4 13 13 3 9 2
16 9 13 3 13 3 3 9 9 2 16 9 4 13 0 9 2
15 9 13 3 3 9 2 15 13 9 0 9 15 9 13 2
14 0 9 7 13 9 13 9 9 2 15 13 0 9 2
13 0 9 1 13 9 9 0 16 9 9 9 1 2
9 13 2 16 9 13 3 3 15 2
3 15 9 2
16 9 0 9 4 13 15 9 2 15 9 7 9 13 3 9 2
16 16 15 13 13 9 2 3 9 4 13 9 7 9 4 13 2
13 0 9 7 9 1 9 13 3 0 9 7 9 2
6 9 12 9 3 9 1
16 9 4 13 3 3 0 9 16 9 12 2 13 0 9 9 2
22 9 13 3 3 0 9 16 9 12 2 9 9 5 9 11 11 9 11 11 13 9 2
16 2 9 9 13 0 0 2 11 13 9 9 2 9 11 13 2
16 11 13 2 16 9 12 9 9 13 2 3 3 16 0 2 2
9 2 13 3 13 9 7 9 9 2
26 9 0 11 7 11 9 13 9 13 0 16 1 11 0 9 2 7 11 9 13 0 9 2 15 13 2
17 11 13 2 16 11 9 13 3 0 13 13 9 0 9 0 9 2
23 15 13 2 16 9 13 9 13 13 9 0 9 15 9 2 2 15 3 13 13 9 2 2
7 0 9 0 9 13 0 9
12 9 2 0 9 9 13 9 9 9 13 0 2
17 9 13 13 7 9 7 0 9 9 13 9 9 9 9 7 9 2
15 9 13 11 9 9 9 0 9 13 13 9 11 11 11 2
20 11 13 9 2 12 9 2 12 9 2 15 2 3 12 0 9 13 9 9 2
23 15 13 9 2 15 4 13 2 13 3 0 9 9 13 0 7 0 9 12 9 0 9 2
19 13 9 1 0 13 12 9 9 12 0 0 9 2 15 9 4 13 15 2
7 9 3 13 12 0 9 2
8 2 15 13 0 13 9 1 2
23 0 9 13 15 9 13 0 9 2 15 13 3 0 9 16 15 2 16 13 9 13 9 2
17 11 11 11 13 2 16 9 13 13 15 0 9 3 16 0 9 2
21 2 16 12 9 3 13 0 13 9 2 13 0 13 3 15 3 13 2 11 13 2
29 9 13 9 2 15 0 9 0 9 9 0 9 13 9 13 9 2 3 9 0 7 0 9 2 9 7 9 1 2
15 2 9 13 3 15 2 15 9 13 2 16 13 7 13 2
18 9 0 9 13 15 2 16 9 13 9 13 7 13 3 3 7 3 2
14 0 9 9 13 9 13 11 1 0 13 9 7 9 2
12 2 13 9 3 2 7 3 13 13 9 9 2
4 9 9 9 9
18 11 9 7 8 9 9 4 13 8 9 9 9 11 11 15 9 9 2
10 9 13 0 0 9 9 7 8 9 2
15 11 11 9 12 13 9 13 9 9 9 7 9 0 9 2
17 9 4 13 11 9 9 9 5 9 2 15 11 9 13 9 12 2
14 9 9 13 9 11 11 7 9 4 13 13 0 9 2
17 9 9 13 2 16 9 4 13 0 9 2 15 9 13 0 9 2
20 9 9 13 0 7 15 9 4 13 9 0 9 2 9 9 9 7 9 9 2
12 9 4 13 11 9 0 9 7 8 9 12 2
18 11 11 13 9 11 9 7 13 8 8 9 9 11 9 9 9 1 2
27 15 4 13 12 0 9 9 9 9 7 13 0 7 0 7 0 9 7 9 2 15 9 4 13 9 9 2
8 15 9 4 3 13 9 9 2
23 11 11 11 2 11 2 3 11 11 2 13 0 9 12 2 11 2 11 2 13 0 9 2
5 15 13 0 9 2
16 11 13 9 12 11 9 11 11 2 15 15 9 13 11 11 2
9 15 13 3 11 9 7 0 9 2
16 15 13 11 11 11 9 12 7 4 13 9 9 3 9 1 2
7 11 13 0 7 13 9 2
22 15 4 13 9 12 11 11 2 11 11 11 9 2 15 15 4 13 13 3 11 11 2
15 11 11 11 11 9 11 11 11 0 9 9 11 11 11 2
13 9 13 9 9 9 7 13 9 13 13 7 13 2
7 11 13 9 11 9 9 2
11 9 13 9 11 2 15 13 9 13 9 2
13 11 7 9 7 9 13 0 9 13 3 9 9 2
19 11 11 11 2 13 0 9 12 11 2 11 2 13 9 2 13 0 9 2
20 15 0 0 9 13 2 11 11 11 11 2 2 12 2 2 15 13 9 9 2
9 11 13 0 9 11 11 11 11 2
26 9 1 15 9 2 15 15 4 13 9 2 13 3 3 9 2 12 2 7 11 13 3 2 12 2 2
9 11 13 9 12 0 9 9 9 2
15 15 13 9 12 11 9 1 9 9 9 9 9 11 11 2
8 11 13 9 12 9 13 9 2
19 9 13 15 11 11 9 0 9 11 2 11 11 2 11 7 11 11 1 2
14 9 9 13 9 9 7 9 2 7 3 9 4 13 2
12 9 12 9 9 13 11 0 9 2 0 9 2
9 9 12 9 13 0 9 12 9 2
15 15 9 13 0 9 9 7 9 9 0 9 0 9 9 2
12 9 13 9 11 2 15 13 9 11 9 12 2
8 3 11 13 0 9 13 9 2
9 9 9 0 9 11 13 11 12 2
15 9 9 13 2 16 11 13 11 0 9 9 7 13 9 2
7 0 9 13 9 13 11 2
8 0 9 9 13 11 9 11 2
15 9 9 11 13 11 12 9 11 11 13 9 0 0 9 2
11 0 9 0 9 13 3 11 7 11 1 2
13 9 13 3 11 11 11 0 9 7 11 11 9 2
10 11 13 3 9 9 1 9 13 12 2
9 9 11 13 11 9 0 9 1 2
9 11 3 13 11 0 9 1 12 2
11 11 13 11 12 11 11 0 0 9 9 2
9 9 9 13 11 3 13 11 12 2
12 9 11 13 11 12 11 11 13 9 15 9 2
8 0 9 11 13 11 9 1 2
13 9 0 9 4 13 12 11 11 11 13 0 9 2
6 9 11 13 11 12 2
13 11 11 11 13 9 9 0 9 7 13 3 9 2
12 1 9 0 9 13 11 9 11 13 0 9 2
7 11 13 9 3 9 12 2
9 11 11 13 0 9 12 9 9 2
9 0 9 13 3 9 9 11 11 2
8 11 13 9 1 9 0 9 2
19 11 11 11 11 13 0 8 8 9 11 11 0 9 7 15 13 9 12 2
8 9 13 9 9 7 9 9 2
11 15 13 11 11 9 9 2 9 11 12 2
11 15 4 13 12 13 0 9 7 9 9 2
8 9 13 0 12 9 9 11 2
7 9 12 9 13 0 9 2
22 0 9 13 4 15 1 13 2 7 0 12 9 0 9 4 13 3 3 16 4 13 2
29 9 2 15 9 1 13 0 2 13 9 9 13 9 3 0 7 0 9 13 0 0 7 0 11 9 9 9 13 2
12 12 9 9 3 1 15 9 9 13 9 9 2
13 9 5 13 15 9 9 9 7 9 5 9 9 2
20 9 9 13 12 9 9 2 9 2 9 7 9 2 9 2 9 9 7 9 2
17 11 11 2 9 11 2 13 0 9 12 2 13 0 0 9 9 2
13 15 13 9 12 11 9 7 9 9 3 12 9 2
10 1 11 9 15 13 9 9 3 11 2
6 9 15 9 13 12 2
6 9 15 13 0 11 2
24 11 2 9 8 2 11 2 11 11 2 11 2 11 2 13 11 11 13 0 9 11 11 9 2
22 11 13 0 7 15 13 12 9 2 15 9 15 13 0 9 2 15 13 15 9 9 2
12 11 13 9 0 2 7 13 13 9 0 9 2
11 11 0 9 13 11 2 11 2 11 2 2
18 3 15 13 11 9 9 9 7 13 11 11 1 2 9 0 2 9 2
21 9 13 11 0 9 2 16 15 13 9 2 11 11 13 3 13 9 7 13 9 2
20 9 1 11 13 9 9 7 13 11 11 7 15 9 9 13 0 9 11 1 2
27 16 11 4 13 2 11 13 0 2 9 0 2 9 15 0 9 2 9 11 11 11 2 7 13 15 3 2
11 0 9 15 13 11 11 2 7 13 3 2
17 11 11 11 11 13 9 11 1 2 7 13 13 15 9 8 9 2
19 15 13 3 11 7 11 11 7 11 11 1 2 7 15 13 3 0 15 2
13 11 11 2 13 12 11 2 13 0 9 7 9 2
8 15 13 9 9 11 11 11 2
24 11 4 13 9 11 7 11 13 9 2 12 2 7 11 2 11 7 9 11 9 2 12 2 2
26 0 11 11 2 9 11 11 7 11 11 2 2 3 12 2 0 9 12 2 13 11 13 9 7 9 2
16 15 13 7 13 11 2 7 13 3 11 11 9 2 11 9 2
6 15 13 3 9 9 2
18 11 0 9 9 9 12 2 3 9 15 13 2 13 11 11 13 9 2
16 11 2 9 8 2 9 8 2 11 2 13 9 11 9 11 2
9 9 12 3 13 3 12 12 9 2
14 9 13 9 12 0 11 9 9 2 9 11 11 1 2
10 15 1 9 9 13 11 2 8 2 2
8 15 9 13 9 9 7 9 2
18 9 13 9 2 9 2 9 7 9 2 15 13 7 13 9 7 9 2
8 9 13 9 2 15 13 9 2
17 9 4 13 0 9 9 2 15 13 9 0 9 13 2 13 9 2
16 9 13 15 13 7 13 2 7 3 0 13 0 2 0 9 2
20 9 9 8 13 9 9 13 9 8 2 9 0 9 3 9 2 9 2 9 2
12 9 13 9 9 8 2 15 13 9 7 9 2
11 9 4 13 0 2 0 2 0 7 0 2
11 0 9 13 3 9 2 7 9 2 1 2
8 0 9 13 9 7 9 9 2
14 0 9 13 9 7 9 2 13 13 0 9 9 1 2
9 9 4 13 9 9 7 9 1 2
11 16 9 13 0 2 9 9 4 13 9 2
12 9 13 3 3 2 16 3 9 9 13 0 2
10 0 9 13 9 1 0 7 0 9 2
6 0 9 13 9 1 2
21 3 0 9 9 4 13 9 2 15 13 15 9 2 3 9 13 9 9 7 9 2
21 11 9 2 9 11 11 11 2 13 11 9 12 2 16 11 9 9 4 13 0 2
13 11 9 13 9 9 2 3 9 13 3 11 9 2
14 11 9 13 9 13 2 7 15 13 0 7 0 9 2
11 3 3 0 9 0 7 0 9 13 0 2
18 11 13 9 11 0 0 9 2 15 9 13 11 0 9 7 9 9 2
14 11 13 0 9 9 2 15 13 9 11 9 9 9 2
22 11 11 11 2 2 11 11 11 11 2 13 11 11 0 9 7 0 9 12 13 9 2
22 9 13 3 3 0 9 11 9 2 16 15 13 0 15 0 9 13 9 1 9 12 2
16 9 4 9 11 11 7 11 15 1 13 11 11 7 11 11 2
11 15 9 13 0 9 12 11 11 9 9 2
37 11 13 11 11 11 2 9 0 9 9 11 11 11 11 9 0 9 7 15 9 15 13 0 9 11 11 11 11 2 15 9 15 13 3 9 12 2
13 11 4 13 11 11 11 2 9 3 9 9 11 2
23 11 4 3 13 9 2 16 9 13 3 9 11 11 11 2 2 16 9 9 13 9 13 2
16 2 11 11 11 11 2 9 13 9 9 13 9 9 13 9 2
11 9 13 3 9 2 15 13 9 11 11 2
18 11 11 11 2 13 11 11 12 9 9 12 7 4 13 3 9 12 2
17 11 11 15 13 9 12 7 9 9 15 13 9 9 12 9 12 2
27 0 9 11 13 11 11 11 11 9 9 12 2 7 13 0 9 9 2 15 15 4 13 3 12 9 9 2
23 9 13 11 0 9 11 11 11 9 7 3 15 13 9 3 9 12 13 11 11 11 11 2
9 9 13 13 3 3 11 9 11 2
19 15 4 3 13 0 13 9 1 2 7 11 0 9 15 4 13 9 12 2
4 9 9 9 1
13 3 12 9 13 11 9 11 11 9 9 9 12 2
15 11 11 0 9 7 11 0 9 13 12 9 9 9 1 2
6 15 13 11 1 11 2
4 9 13 9 2
14 11 0 9 9 11 11 1 11 13 13 9 11 9 2
13 11 13 13 2 13 15 13 0 9 7 9 9 2
12 9 13 2 16 11 9 4 13 9 9 9 2
13 11 9 9 9 12 0 9 13 3 9 9 11 2
9 3 16 9 13 9 15 9 9 2
9 9 1 11 9 13 9 9 11 2
12 3 11 9 13 3 3 11 9 0 9 1 2
8 11 9 12 9 12 9 9 13
15 9 11 4 13 9 12 9 13 9 12 9 9 13 9 2
6 9 13 9 11 11 2
19 11 4 13 9 9 12 1 2 7 0 9 1 15 13 4 13 3 9 2
12 9 12 11 9 9 13 9 3 12 12 9 2
18 2 16 9 13 2 13 0 13 9 9 3 3 16 13 12 9 9 2
8 15 9 13 13 9 15 9 2
7 15 4 13 12 9 9 2
15 13 15 1 2 16 13 9 9 12 2 11 13 11 9 2
2 11 11
9 9 9 11 11 13 3 9 11 2
16 0 9 9 11 13 11 9 11 11 2 9 9 7 15 9 2
11 9 13 9 11 9 7 11 9 13 9 2
7 11 9 1 13 9 9 2
16 15 1 9 11 11 2 11 2 4 13 9 9 11 9 1 2
12 9 13 9 9 9 2 15 13 11 13 9 2
4 9 13 9 11
16 11 11 9 13 0 9 7 9 13 15 9 11 1 11 9 2
8 9 13 9 12 9 11 9 2
19 9 13 9 9 13 9 9 2 7 9 12 9 12 13 2 12 15 3 2
8 3 13 13 9 1 9 9 2
13 9 9 1 9 13 9 9 9 7 13 9 3 2
11 3 9 13 13 9 9 7 12 9 9 2
22 9 13 3 0 9 9 15 9 16 3 0 9 1 13 13 9 2 15 13 13 9 2
11 9 7 0 9 13 4 3 13 9 1 2
3 9 13 13
10 11 13 3 9 2 16 15 13 9 2
16 6 16 15 13 16 15 13 3 7 3 7 15 3 13 15 2
5 11 3 13 13 2
3 13 13 3
6 13 15 13 3 9 2
13 2 15 13 3 2 16 3 13 7 13 9 2 2
3 13 13 9
11 13 9 2 16 13 9 9 3 16 0 2
3 13 13 9
9 11 13 0 2 0 2 3 0 2
22 15 13 0 9 9 13 10 12 0 9 15 15 13 3 15 13 0 9 3 13 15 2
5 9 13 10 9 2
4 13 3 3 2
4 15 13 11 2
6 9 13 7 9 13 2
5 13 3 1 9 2
4 13 3 9 2
13 15 13 3 13 2 16 12 9 9 13 0 9 2
10 2 13 13 9 2 2 13 9 15 2
12 0 3 13 3 9 3 11 2 11 7 11 2
6 9 13 13 9 9 2
7 9 9 13 0 0 9 2
6 15 13 13 9 13 2
7 9 13 13 3 9 9 2
5 9 13 13 13 2
17 9 13 13 0 2 7 9 13 9 9 13 2 13 7 9 13 2
3 3 13 9
17 3 15 3 13 3 9 0 2 3 13 0 7 0 7 15 13 2
11 10 9 13 10 9 2 15 13 9 1 2
5 3 3 13 13 2
5 15 13 9 3 2
13 9 13 13 3 9 2 7 9 15 13 13 13 2
2 13 11
14 0 9 1 9 13 15 2 16 0 9 9 13 9 2
26 0 0 9 13 3 12 12 2 7 13 12 7 12 9 7 15 3 0 9 3 13 3 15 13 12 9
4 15 13 9 2
17 9 13 12 12 9 0 9 13 13 2 16 9 13 13 10 9 2
6 13 13 3 13 3 2
7 9 0 9 13 15 3 2
6 15 13 12 12 9 2
9 11 13 2 16 11 13 3 9 2
13 10 0 9 13 3 0 2 16 9 13 13 13 2
17 3 11 7 11 13 0 9 2 15 1 11 13 0 9 9 9 11
7 9 9 9 13 12 9 2
6 9 13 13 0 9 2
14 15 13 13 3 11 2 7 13 13 10 9 9 13 2
13 11 9 13 13 9 2 16 9 13 13 9 9 2
12 13 3 2 13 15 13 2 15 15 15 13 2
4 13 15 9 2
6 15 13 3 9 7 2
6 11 9 13 13 9 2
10 9 13 3 3 3 2 3 11 13 2
5 15 13 0 9 2
5 15 13 9 13 2
7 13 9 3 3 0 9 2
2 3 3
4 9 13 3 12
8 0 9 13 3 0 13 11 9
3 9 9 9
6 15 3 13 9 13 2
23 15 3 13 2 16 15 13 10 9 9 2 15 13 3 0 7 15 1 15 13 3 0 2
7 15 13 13 3 10 0 2
2 11 9
20 9 1 11 13 9 13 9 13 9 7 10 9 2 16 13 13 13 9 9 2
4 15 13 6 2
19 9 9 13 13 0 9 0 9 9 9 13 3 2 16 15 13 9 9 2
13 6 3 2 11 2 9 13 15 2 16 13 13 2
14 0 9 9 9 13 9 9 12 9 13 7 9 13 2
8 9 15 13 7 9 13 13 2
6 0 15 13 3 13 2
6 10 13 13 0 9 2
3 15 3 0
15 15 13 3 0 9 2 15 13 13 13 13 3 0 9 2
9 10 0 13 3 13 9 9 13 2
3 13 15 2
5 10 9 13 11 2
3 11 9 9
2 13 9
8 9 13 9 3 0 16 9 2
8 16 9 13 2 9 13 0 2
13 9 11 13 3 2 16 9 9 9 13 9 9 2
14 15 1 15 13 11 2 16 3 9 13 3 3 9 2
10 9 9 13 0 9 7 9 11 11 2
4 0 7 0 11
14 9 13 2 3 3 9 11 11 13 13 0 0 9 2
6 9 13 13 15 13 2
9 13 10 9 9 7 15 3 13 2
4 0 9 10 15
6 9 13 9 9 1 2
9 9 9 7 10 9 13 0 9 2
11 10 9 13 13 7 9 13 9 13 9 2
2 13 9
9 9 13 2 13 15 13 11 9 2
10 9 7 9 13 10 3 9 7 9 2
19 3 3 0 9 13 3 0 11 9 2 16 3 15 9 13 13 0 9 2
6 9 13 2 9 13 2
2 13 3
9 16 13 13 15 0 2 13 3 2
11 0 0 9 9 2 15 13 13 10 9 2
5 15 13 15 13 2
12 15 13 3 13 15 3 9 3 1 9 9 2
11 11 9 13 13 9 9 7 11 0 9 2
7 15 9 13 12 9 9 2
11 15 13 13 13 13 13 9 2 9 2 2
8 3 13 2 16 0 15 13 2
10 2 15 13 15 15 2 16 13 0 2
6 13 11 9 0 9 2
5 9 13 9 0 2
5 0 9 0 9 2
7 9 9 13 13 3 3 2
8 12 9 15 13 3 3 9 2
12 11 0 7 3 0 9 13 13 13 9 9 2
6 15 9 9 13 9 2
7 9 13 3 3 9 9 2
6 15 13 13 11 9 2
4 11 13 9 9
2 13 13
6 13 15 3 3 9 2
4 15 13 9 2
7 3 15 13 13 9 0 2
9 9 13 0 3 3 0 7 0 1
6 11 13 9 13 9 2
19 10 9 9 13 9 15 13 0 9 2 16 9 13 13 7 13 11 9 2
11 3 15 3 13 2 16 9 13 13 13 2
8 9 13 13 3 16 13 13 2
2 0 9
17 7 9 1 13 2 3 16 15 13 3 3 13 3 13 3 9 2
8 9 7 0 11 13 3 3 2
26 0 9 7 9 9 13 9 2 16 13 9 9 11 13 0 13 0 9 2 16 15 0 9 3 13 2
9 9 13 15 13 13 15 3 9 2
7 3 13 0 13 0 9 2
7 9 13 13 3 16 13 13
9 9 13 13 13 10 10 9 9 2
13 16 9 13 0 7 15 13 2 15 13 3 9 2
13 12 3 0 9 13 13 15 3 10 3 13 9 2
6 3 15 13 9 3 2
5 13 15 13 9 2
6 0 9 13 13 0 2
16 9 13 9 13 3 16 15 13 2 7 13 3 16 15 13 2
17 7 0 13 2 16 15 13 0 0 9 2 13 13 13 0 0 2
4 15 13 15 2
17 13 10 10 9 13 7 13 15 13 9 2 7 13 9 2 9 2
9 13 0 2 16 15 13 13 3 2
3 9 13 0
7 6 15 13 10 0 9 2
3 3 13 13
2 0 9
11 7 15 13 3 7 15 3 10 0 9 2
29 16 11 9 13 10 0 9 11 11 2 11 13 2 2 0 7 0 13 3 0 9 9 2 15 13 13 3 9 2
3 9 13 13
13 16 13 11 13 10 0 9 2 3 15 13 0 9
16 0 9 13 9 0 9 3 7 9 13 0 0 2 3 13 2
6 15 13 13 0 9 2
6 9 13 9 12 9 2
12 16 9 9 13 15 0 7 0 9 7 9 2
21 3 12 9 13 0 2 16 11 9 1 9 13 9 2 7 10 9 10 9 13 2
18 3 13 13 13 13 11 3 10 9 1 2 7 3 9 7 12 1 2
6 15 1 13 13 3 2
9 3 9 3 13 2 13 9 1 2
14 16 0 9 13 10 9 2 15 13 9 13 3 9 2
6 13 13 16 11 13 2
9 9 13 13 3 9 9 16 15 2
8 9 13 3 13 9 3 12 2
9 13 10 9 2 16 13 0 3 2
4 9 13 9 2
2 3 2
14 16 15 13 9 2 15 13 15 3 15 3 0 9 2
12 11 13 3 0 9 2 15 15 13 3 13 2
7 13 15 15 3 13 15 2
9 11 13 9 10 9 9 0 9 2
6 11 13 13 15 13 9
13 9 2 9 2 13 0 16 15 13 16 9 9 2
4 9 13 9 9
10 3 15 13 0 9 2 3 13 9 2
8 9 13 9 2 16 0 0 2
8 9 11 13 9 13 13 15 2
9 6 3 13 9 2 11 13 13 2
18 9 13 3 9 13 0 9 2 15 13 13 3 13 0 9 9 9 2
4 13 1 12 2
9 15 15 13 13 2 16 13 9 2
14 3 15 13 13 15 13 13 2 16 9 13 0 0 2
14 15 3 13 11 13 7 0 9 2 11 13 9 9 2
6 9 13 13 3 3 2
12 9 15 13 9 9 2 11 2 11 2 11 2
10 9 13 16 9 2 9 13 12 9 2
4 15 16 13 15
2 13 13
6 15 13 3 3 13 2
3 0 0 9
13 3 11 13 13 0 13 12 9 15 1 3 15 2
6 15 13 2 15 3 13
5 15 9 13 15 2
7 9 1 15 13 3 0 2
3 15 13 13
7 15 13 3 0 10 10 9
5 9 0 2 13 9
6 13 13 3 13 9 2
5 15 13 11 1 2
5 13 13 3 12 9
9 2 15 3 2 15 13 13 13 2
8 11 13 10 9 12 11 9 2
12 0 9 13 3 13 2 9 13 7 0 13 2
9 13 3 3 2 16 13 13 9 2
6 11 9 13 10 9 2
12 3 10 9 15 2 15 13 0 9 0 9 2
14 15 13 2 3 13 11 9 0 13 9 7 13 3 2
4 13 15 13 2
5 13 9 9 13 2
6 15 13 3 9 9 2
5 15 13 3 9 2
9 11 13 13 3 13 9 7 9 2
7 9 3 13 3 2 3 2
5 13 9 0 9 2
11 3 13 10 9 13 3 2 13 3 13 2
19 10 9 9 15 3 13 2 15 15 13 2 9 2 9 2 10 9 9 2
7 13 15 9 9 2 13 2
6 6 16 15 3 13 2
9 3 15 13 13 12 0 0 9 2
9 0 9 3 13 12 7 12 9 2
4 15 13 11 2
10 3 16 13 2 13 13 13 15 15 2
3 9 9 9
5 13 3 13 9 2
11 16 13 3 9 3 2 13 13 0 9 2
2 9 3
3 13 9 2
8 9 13 3 0 7 0 9 2
5 3 11 13 9 2
5 13 3 15 3 9
6 15 13 15 3 3 2
3 13 13 13
12 0 9 13 3 13 9 7 13 9 9 13 2
9 11 13 9 13 3 3 0 9 2
3 9 13 13
6 15 13 3 10 9 2
5 15 13 9 9 2
7 9 13 9 3 12 9 2
19 11 13 3 2 13 9 7 13 9 7 9 7 13 3 9 9 13 9 2
5 11 13 12 0 2
9 9 13 13 13 7 13 11 9 2
7 15 13 13 15 2 16 2
8 13 9 7 9 9 3 0 2
3 9 13 3
4 13 15 15 2
16 3 2 9 2 9 9 13 3 15 2 15 15 13 0 9 2
13 3 3 9 13 3 9 2 16 15 3 13 9 2
6 15 13 15 3 3 2
3 9 13 3
9 15 13 13 15 3 2 0 9 2
7 0 3 11 13 13 9 2
7 13 7 15 13 0 9 2
3 13 9 9
13 15 13 16 6 3 15 13 3 13 3 3 13 2
8 9 13 9 2 13 15 13 2
4 9 7 9 9
14 9 11 9 13 3 0 2 16 0 9 13 3 9 2
10 9 13 0 13 2 16 15 13 13 2
5 9 13 13 0 2
4 9 16 15 13
6 15 13 9 11 1 2
11 3 3 15 13 9 2 3 9 7 9 2
11 9 13 13 2 7 13 3 13 13 3 2
7 13 0 9 9 3 3 2
8 9 9 13 9 3 9 9 2
16 9 13 3 3 0 2 16 9 13 9 13 3 3 3 0 2
8 13 3 13 15 3 15 1 2
4 13 15 1 2
8 11 9 13 13 9 0 9 2
9 15 13 9 1 13 0 9 3 2
10 13 11 8 7 13 2 15 13 13 0
5 9 9 13 13 2
3 9 15 13
4 15 13 13 9
13 1 9 13 9 9 7 15 13 13 0 0 9 2
7 13 3 9 0 16 9 2
17 9 11 13 9 0 9 9 2 9 1 9 2 9 7 9 9 9
7 11 13 11 12 0 9 2
5 15 13 13 9 2
5 9 13 9 9 2
4 9 13 9 0
6 13 2 16 13 13 2
6 9 13 3 9 1 2
16 11 9 9 13 13 13 0 9 2 16 9 9 12 3 13 2
10 15 13 3 9 1 2 13 15 13 2
8 13 0 9 13 9 9 3 2
7 9 7 9 13 3 0 2
10 12 9 13 11 9 13 9 9 9 2
11 9 13 13 0 7 9 13 3 0 3 2
6 13 13 3 12 1 2
34 3 15 13 10 0 9 15 13 3 13 3 0 15 13 13 13 3 15 13 3 0 16 15 13 13 3 10 9 3 7 3 15 13 13
5 9 13 15 9 2
5 9 13 0 9 2
8 11 9 13 9 13 9 9 2
14 16 9 13 0 2 13 15 3 15 13 3 9 9 2
4 13 13 15 2
15 15 13 3 3 3 10 9 16 3 16 0 13 9 13 2
17 15 13 3 12 0 9 15 11 11 13 13 3 0 2 0 9 2
4 13 9 9 3
5 11 13 11 9 2
9 9 13 13 2 16 15 13 3 2
5 13 13 3 9 2
6 10 12 3 13 9 2
12 9 0 9 13 9 11 9 7 13 12 9 2
4 13 15 3 2
9 15 13 13 12 7 15 13 9 13
8 11 11 13 11 9 1 9 3
6 13 2 16 15 13 2
3 9 9 2
5 13 0 13 11 2
2 13 15
10 11 13 13 9 9 7 13 15 9 2
2 15 1
6 11 13 13 9 9 2
11 15 13 13 3 2 16 3 13 10 9 2
12 13 15 15 2 16 9 13 9 3 12 9 2
13 3 15 13 3 13 2 13 3 9 7 0 9 2
15 11 13 9 13 3 3 16 9 3 12 9 13 9 1 2
10 9 3 13 2 16 3 0 9 13 2
14 10 9 7 9 13 3 13 9 1 7 13 3 3 2
15 11 13 9 2 16 10 9 7 9 13 13 13 9 3 2
9 13 3 9 16 13 13 3 9 2
4 9 13 15 9
2 13 13
5 9 13 9 9 2
16 11 13 13 15 1 15 2 16 15 13 9 15 1 16 9 2
5 9 13 0 9 2
6 9 9 3 0 11 9
5 15 13 9 13 9
4 13 0 9 9
11 2 13 15 10 0 9 13 2 15 13 2
11 9 9 13 9 13 10 9 3 13 9 2
19 9 13 9 1 7 13 10 9 9 13 9 11 2 15 15 13 9 9 2
7 9 13 12 9 0 9 2
7 13 11 9 1 13 9 2
4 13 10 9 2
8 2 15 13 13 0 9 2 2
10 9 13 13 9 2 9 16 3 13 13
9 3 13 3 13 13 9 10 9 2
7 15 13 13 13 13 3 2
9 11 9 9 13 9 3 7 9 2
9 11 13 16 15 13 0 9 3 2
3 9 13 9
7 9 13 13 1 9 9 2
21 9 13 2 16 15 15 13 15 2 15 13 3 3 2 16 9 13 13 3 0 2
4 9 13 0 13
11 13 3 13 2 3 15 13 13 10 9 2
15 15 13 9 10 9 2 16 11 13 0 9 7 13 13 2
5 9 13 15 9 2
3 2 15 2
12 9 13 13 10 15 2 15 3 13 13 9 2
16 15 7 3 10 15 1 3 13 13 9 9 2 15 13 13 2
10 13 3 2 0 9 2 9 15 13 2
8 9 13 9 13 3 10 9 2
8 13 15 13 9 9 9 9 2
9 15 13 3 13 13 9 10 9 2
13 9 9 9 13 13 0 9 2 16 9 13 3 2
13 9 11 9 9 13 13 9 9 9 13 11 11 2
7 13 12 9 11 13 9 2
8 10 9 13 9 7 13 12 2
4 13 13 15 2
4 13 13 9 2
11 3 13 0 9 2 13 9 13 3 3 2
15 9 13 9 3 2 16 3 9 9 13 0 9 9 9 2
11 11 13 13 3 10 0 9 8 13 11 2
14 3 15 13 13 9 3 2 3 15 13 13 13 9 2
4 3 15 13 2
7 13 15 3 15 13 13 2
11 16 9 13 13 3 2 9 13 13 0 2
6 11 13 3 13 9 2
13 3 3 3 10 9 13 15 2 16 15 13 3 2
4 13 3 3 13
12 11 13 2 9 13 9 7 15 13 15 15 2
7 13 15 15 13 7 15 2
2 13 13
7 9 13 3 0 9 1 2
2 13 9
12 9 13 3 13 2 16 11 9 13 0 13 2
5 10 9 13 9 2
2 9 1
5 9 13 0 9 2
6 13 2 3 9 9 2
9 10 0 13 13 9 3 3 3 2
8 7 13 3 0 2 0 9 2
3 13 9 1
7 9 13 9 0 0 9 2
7 9 13 3 7 13 9 2
11 11 9 13 3 0 3 7 3 0 11 2
14 10 9 0 7 0 2 7 0 2 9 13 9 7 2
8 0 9 11 13 11 12 9 2
17 3 13 3 3 11 13 13 0 9 9 2 8 8 8 8 8 2
5 9 13 13 9 13
8 6 3 15 3 3 9 13 2
6 10 9 13 13 0 2
8 0 9 13 8 7 9 11 9
6 9 13 9 9 1 2
12 9 0 3 12 9 13 13 1 9 1 9 2
2 9 13
9 13 9 13 13 9 9 10 9 2
4 15 13 0 13
21 10 11 9 13 9 9 9 2 7 9 7 9 13 13 3 11 2 11 7 11 2
4 13 9 9 2
14 3 9 7 9 13 3 3 13 15 1 13 9 9 2
7 9 13 3 2 13 13 2
10 13 3 3 13 13 3 3 13 9 2
4 11 13 11 9
15 0 9 13 3 12 9 7 9 2 15 13 15 3 9 2
15 9 13 9 7 9 13 9 7 9 7 9 13 0 3 2
11 10 9 16 15 13 0 9 2 7 13 2
3 9 13 9
8 9 13 13 13 3 3 3 2
6 13 16 11 13 11 2
11 11 11 13 9 2 7 13 15 13 9 2
2 9 9
2 11 9
5 9 13 9 12 2
6 13 15 9 2 11 2
4 15 13 0 2
9 3 13 3 13 3 3 16 3 2
5 0 9 9 13 2
8 3 13 9 0 9 9 9 2
5 13 15 3 3 2
4 9 13 3 2
3 13 13 2
8 3 9 13 2 11 13 15 9
12 0 9 13 9 0 9 13 13 3 3 3 2
6 3 15 13 9 3 2
3 15 13 0
5 9 9 13 0 2
8 15 13 0 13 0 9 9 2
5 13 2 16 13 2
8 9 13 13 12 9 9 3 2
4 9 13 9 2
2 3 3
11 15 16 13 13 2 13 13 10 9 13 2
2 9 1
11 9 13 3 9 2 10 9 9 3 13 2
9 3 13 13 0 13 9 9 9 2
9 9 7 9 13 13 13 9 3 2
5 3 9 9 13 2
6 9 13 2 13 9 2
23 3 15 13 13 16 15 13 10 0 9 7 3 3 9 13 10 0 9 7 9 3 7 2
6 15 15 13 10 9 2
11 3 9 13 9 13 9 0 11 7 11 2
4 9 13 13 9
3 3 9 1
7 11 13 11 9 3 12 2
6 0 9 9 13 0 2
3 13 9 2
13 10 9 13 3 13 16 12 9 2 15 13 9 2
5 13 13 13 9 2
2 13 9
5 15 1 9 13 2
22 3 2 9 9 1 2 9 1 2 13 9 13 9 9 1 9 13 10 9 2 9 2
7 12 9 13 13 3 13 2
4 11 9 13 2
21 16 9 13 2 11 13 13 0 2 16 13 2 3 15 13 0 9 13 0 9 2
7 15 13 9 9 3 3 2
18 15 13 9 11 11 2 15 13 13 9 9 9 7 11 16 11 9 2
7 10 9 13 13 1 9 2
8 9 13 0 1 9 13 9 2
10 3 13 9 2 15 13 13 7 13 2
11 11 9 13 13 10 0 0 3 0 13 2
6 3 13 3 13 9 2
10 15 13 9 2 0 10 0 7 0 2
10 13 0 9 2 16 13 3 13 11 2
2 9 1
3 13 13 9
9 12 9 11 13 3 13 11 12 2
2 9 1
10 13 10 9 9 9 12 9 12 9 1
11 13 2 13 9 7 9 7 13 3 11 2
8 9 13 13 13 0 9 1 2
8 15 13 13 0 0 9 1 2
23 13 13 0 9 11 2 7 15 13 3 0 9 2 16 13 13 15 13 10 9 7 9 2
11 13 9 2 16 9 13 10 9 3 13 3
9 3 16 13 3 0 3 15 13 2
2 9 1
2 3 3
3 15 13 9
7 13 0 9 2 15 13 2
5 11 13 3 13 9
18 13 15 3 13 13 3 2 16 15 13 2 16 9 9 13 13 13 2
8 3 0 11 13 9 3 9 2
16 10 9 9 13 3 0 3 13 2 16 9 13 15 3 13 2
8 15 13 13 9 2 15 13 2
8 3 15 9 9 13 3 9 2
10 15 13 3 3 16 13 13 15 0 2
6 15 13 13 3 9 2
5 13 13 9 3 13
10 7 13 16 3 2 0 9 13 13 9
11 15 13 9 3 9 2 16 3 13 13 2
3 6 0 2
9 10 9 13 3 13 0 9 1 2
3 13 1 9
19 9 13 13 3 9 2 15 9 9 13 9 1 13 3 9 7 13 9 2
13 16 9 13 3 9 2 12 12 9 2 9 13 2
6 11 13 0 9 9 2
8 9 9 9 13 9 0 9 2
19 16 13 16 15 13 0 2 15 13 16 15 13 9 13 2 3 0 9 2
11 9 13 13 0 9 7 13 0 0 9 2
5 15 13 3 9 2
18 10 9 13 0 9 13 15 13 3 16 11 0 9 13 3 1 9 2
7 9 13 9 11 9 3 2
5 13 9 9 11 2
12 9 13 9 3 13 3 13 2 7 13 0 2
5 7 11 13 9 2
10 10 9 15 13 13 3 2 3 9 2
4 13 9 9 2
9 9 9 13 3 9 13 9 9 2
9 9 13 2 7 15 13 13 3 2
6 15 9 13 3 3 2
8 9 13 0 9 0 9 3 2
11 11 13 13 3 9 2 13 9 3 9 2
15 3 0 13 2 16 13 3 9 7 9 13 13 9 1 2
17 13 0 9 7 9 15 2 11 13 0 13 3 13 9 12 9 2
4 13 13 13 13
13 13 11 13 2 16 10 9 13 13 2 13 11 2
6 11 13 9 3 3 2
10 11 9 13 3 3 11 7 11 9 2
17 3 15 0 13 16 13 13 2 0 0 2 0 9 13 9 0 2
10 9 13 9 13 9 2 16 0 13 2
13 9 13 13 0 9 3 10 3 16 9 9 9 2
4 11 13 9 11
2 7 9
8 15 13 3 3 3 9 1 2
9 10 15 15 13 2 16 13 9 2
8 11 9 9 3 13 0 3 2
13 9 9 13 11 9 2 15 13 9 9 13 9 2
12 9 13 9 1 13 7 0 2 0 9 13 2
4 13 3 15 13
13 13 13 2 16 11 13 0 9 13 13 9 9 2
7 3 3 11 13 0 9 2
2 9 9
5 3 13 13 3 2
9 11 13 13 3 10 9 9 9 2
2 3 9
2 0 11
6 13 3 13 10 9 2
4 9 13 3 2
4 13 9 0 9
2 0 9
3 13 3 2
7 15 15 13 16 13 9 2
7 0 15 13 11 3 0 2
2 9 9
8 0 9 13 13 9 7 9 2
4 13 15 13 2
5 13 3 10 9 2
5 15 13 3 3 15
12 9 13 13 0 7 0 2 3 13 13 13 2
7 11 0 9 13 13 9 2
12 6 7 15 13 3 3 3 3 3 3 8 2
8 13 2 16 9 13 13 12 9
9 10 9 9 7 9 1 13 0 2
4 9 13 3 2
2 0 9
7 3 16 3 9 13 9 2
6 3 15 13 9 13 2
2 9 9
15 9 13 2 16 15 13 0 9 9 2 9 13 3 12 2
2 0 9
17 11 9 13 10 9 2 16 0 9 13 3 0 16 13 13 3 2
5 11 9 11 1 2
5 13 3 3 12 2
3 9 9 9
6 13 15 3 16 0 2
11 16 9 13 13 3 2 13 13 13 3 2
9 11 9 13 3 13 3 3 9 2
6 16 13 3 3 9 2
8 6 16 0 2 16 15 13 2
9 9 3 13 2 13 9 13 9 2
11 9 13 13 9 9 1 13 9 0 9 2
12 9 13 13 9 9 2 7 15 13 3 13 2
10 0 9 9 13 9 0 9 3 13 2
3 15 13 9
10 13 13 13 3 16 15 3 13 0 2
8 15 13 10 9 7 3 13 2
4 11 3 13 9
10 13 10 9 2 3 9 11 13 15 2
8 7 10 9 13 13 3 9 2
4 13 15 9 2
28 3 6 3 15 15 13 16 13 13 7 15 3 13 16 16 16 13 15 13 15 15 13 3 13 3 15 13 3
11 11 13 9 0 9 0 9 16 11 3 2
5 9 13 9 13 2
3 9 11 9
25 13 13 3 13 9 10 0 9 9 15 13 3 9 7 3 13 3 9 0 9 7 10 0 9 2
11 16 15 13 13 9 3 2 13 13 15 9
11 9 13 9 13 1 9 2 3 9 1 2
3 0 15 13
7 13 13 9 3 9 1 2
10 9 13 3 3 0 9 16 9 0 2
9 15 13 9 2 15 13 15 0 2
3 0 9 13
9 10 9 16 15 13 13 15 9 2
5 3 9 13 11 2
11 15 13 0 9 2 16 13 3 0 11 2
6 13 15 13 9 13 2
2 9 13
4 15 13 13 9
2 9 9
10 16 9 3 13 10 9 9 13 2 3
6 3 13 16 9 13 2
21 7 16 15 15 13 3 10 2 9 11 3 15 13 3 0 16 13 15 13 15 2
2 10 9
6 3 13 9 13 9 2
6 9 1 9 13 0 2
11 13 13 3 13 1 2 7 13 13 1 2
4 9 13 9 2
5 3 15 15 13 2
8 9 13 13 13 13 3 9 2
5 13 13 15 13 2
17 13 13 2 11 11 13 2 9 9 2 7 2 9 2 9 9 2
6 7 3 3 13 9 2
19 0 9 15 13 13 2 16 10 0 9 13 3 3 9 16 15 10 9 2
7 10 9 13 0 9 9 2
5 11 13 11 0 2
28 9 1 9 9 13 12 9 9 13 12 9 9 13 2 16 9 13 13 12 9 2 12 9 3 12 0 9 2
3 15 13 9
6 13 3 13 10 9 2
7 3 0 9 9 13 0 2
8 10 9 1 15 13 13 13 2
7 15 13 13 13 15 9 2
11 12 9 13 7 13 9 9 12 7 12 2
13 9 13 3 7 11 3 13 16 3 11 3 13 2
8 12 15 13 9 7 12 9 2
6 13 16 15 13 9 2
5 15 13 9 9 2
21 2 15 13 15 0 9 7 10 9 1 13 13 2 16 15 13 0 0 9 9 2
7 15 13 3 9 9 3 2
8 13 13 3 13 15 13 15 2
5 13 15 3 0 2
10 13 3 9 2 7 9 10 3 13 2
18 16 3 13 10 9 13 16 15 13 13 3 1 15 13 3 0 9 2
7 9 13 3 3 9 13 2
6 3 9 13 3 9 13
4 13 13 9 2
2 10 9
14 9 3 15 13 0 2 7 3 9 13 9 13 13 2
2 13 13
5 9 13 9 9 2
5 15 13 9 3 2
7 0 3 0 9 13 9 2
15 11 1 11 13 0 9 2 15 13 3 0 9 11 11 2
7 9 13 9 0 9 3 2
4 10 12 11 9
10 0 9 15 13 9 2 7 15 13 2
6 9 13 11 9 13 2
5 6 13 15 9 2
9 15 13 9 7 15 13 13 9 2
5 13 9 9 15 2
11 10 9 13 15 2 16 9 13 11 9 2
12 10 10 15 0 9 13 13 13 3 9 9 2
6 3 15 3 15 13 2
3 13 9 9
6 13 13 3 9 12 1
2 0 9
8 13 9 13 9 2 7 13 2
13 11 13 9 15 13 3 3 3 16 13 9 13 2
3 7 10 0
4 15 15 13 2
6 13 3 16 9 13 2
5 11 13 3 9 2
19 15 13 2 13 15 15 7 13 13 2 2 3 15 1 2 0 3 13 2
22 15 13 9 9 7 15 13 9 7 15 15 2 3 9 13 7 3 15 13 3 3 2
8 0 11 13 13 3 9 9 2
11 15 13 13 0 9 0 9 7 13 9 2
12 3 0 9 1 9 13 13 0 9 9 9 2
6 0 13 10 0 9 2
5 9 13 3 0 2
4 2 10 9 2
3 10 15 9
2 9 9
12 13 10 9 3 0 13 2 16 0 13 13 2
8 13 3 0 13 13 0 9 2
4 2 3 0 2
12 9 13 13 9 0 15 2 15 13 9 13 2
12 9 9 13 13 3 0 12 3 13 9 1 2
9 10 10 9 13 13 9 7 9 2
2 13 13
4 9 9 2 11
8 11 11 9 13 0 0 9 2
12 16 12 9 13 2 3 15 13 15 3 9 9
5 13 3 13 9 2
6 15 13 9 9 1 2
13 13 13 3 13 9 16 15 13 3 10 9 13 2
8 0 9 13 3 10 9 13 2
14 15 13 3 13 15 2 16 13 9 13 0 15 3 2
2 0 9
10 9 13 13 2 13 16 13 13 3 2
2 13 13
8 11 9 11 13 13 9 1 2
4 3 15 13 2
4 15 13 0 2
10 3 9 13 12 9 9 9 3 13 2
10 3 9 9 3 15 13 10 9 9 2
4 9 3 0 9
11 11 9 0 9 13 3 3 1 11 9 2
7 9 13 13 3 16 3 13
12 3 13 2 3 9 13 2 7 13 0 9 2
5 13 9 13 9 2
2 9 9
5 13 13 15 0 2
10 15 15 13 2 15 13 0 9 3 2
9 3 3 13 9 13 0 0 9 2
8 9 13 9 9 7 3 9 2
14 9 9 9 1 13 0 15 2 16 13 13 0 9 2
19 11 13 13 3 0 9 2 15 10 9 13 9 2 16 9 13 3 3 2
8 3 9 11 9 13 13 13 2
8 11 13 2 16 13 9 13 2
9 13 13 2 13 9 7 9 13 2
14 3 2 3 11 2 16 15 3 13 0 10 0 9 2
5 0 9 13 15 2
6 9 13 12 0 9 2
4 3 9 7 9
6 3 15 13 13 9 2
9 3 13 9 0 0 13 9 9 2
6 9 13 3 9 11 2
3 10 9 1
4 13 9 3 9
11 9 13 13 0 9 9 0 7 0 9 2
15 3 16 13 9 9 7 9 2 13 3 9 13 7 13 2
2 2 13
13 2 15 10 11 11 3 13 2 2 13 9 9 2
15 13 15 13 2 10 9 2 13 0 9 3 10 9 13 2
13 13 2 16 9 13 9 9 7 13 3 9 9 2
7 9 13 13 9 3 9 2
6 13 9 3 0 9 2
10 6 10 0 0 13 9 2 13 9 2
4 15 13 15 9
2 9 9
5 16 15 15 13 2
13 9 13 3 9 9 2 15 16 13 13 9 9 2
4 13 9 13 3
5 13 15 9 1 2
33 7 3 3 3 15 13 10 10 9 7 13 16 13 15 9 9 7 7 3 15 13 16 16 6 13 3 16 13 15 3 15 1 13
10 3 15 13 13 13 2 16 13 9 2
16 16 13 2 16 9 13 7 13 3 9 2 15 13 16 9 2
8 9 13 9 0 9 0 9 2
4 9 13 9 2
8 0 13 11 8 8 9 9 12
3 13 9 0
12 11 13 9 3 3 2 16 13 13 13 13 2
23 2 15 13 9 9 0 9 2 16 11 9 7 11 13 12 7 15 9 2 2 15 13 2
2 13 1
11 12 9 2 15 13 11 9 2 13 0 2
7 13 9 13 3 9 12 2
6 13 3 3 12 1 2
6 9 9 13 0 9 2
7 10 9 13 13 10 0 2
5 13 3 0 13 2
5 13 13 3 9 2
5 13 10 0 9 2
2 10 3
5 9 13 13 13 2
8 3 9 13 0 2 0 9 2
9 3 15 13 3 3 13 10 9 2
12 9 15 15 13 3 0 0 13 3 3 0 2
8 13 15 3 13 10 9 3 2
3 9 13 9
11 9 13 13 9 15 7 15 15 13 13 2
5 11 13 0 9 2
10 0 9 13 3 9 2 3 13 13 2
15 11 13 2 16 0 9 15 13 11 9 1 12 9 9 2
11 15 13 9 7 13 9 13 2 0 9 2
4 15 13 9 2
12 13 3 15 13 2 15 13 7 13 9 9 2
11 16 9 13 3 2 9 0 9 13 3 2
4 13 15 0 2
3 13 15 15
10 16 9 13 3 2 13 3 13 9 2
28 3 15 3 13 13 3 3 2 3 3 10 9 9 2 16 9 13 13 12 7 12 2 7 9 13 10 9 2
11 13 3 0 2 16 13 13 3 13 15 2
12 3 15 13 13 8 7 3 9 1 10 9 2
9 11 9 13 0 16 11 13 13 2
6 13 0 13 0 9 2
3 9 10 9
7 15 13 13 0 9 9 2
5 13 15 15 13 2
13 9 13 13 13 3 2 16 10 9 13 9 13 2
5 13 3 9 3 2
5 9 13 9 13 2
9 13 15 9 7 9 13 9 9 2
17 10 9 13 9 9 13 3 13 2 16 15 13 10 0 9 13 2
9 15 13 13 3 9 2 13 9 2
2 3 0
4 13 15 9 2
2 13 0
13 16 13 0 2 3 3 9 13 2 15 13 0 2
2 6 6
4 15 3 13 2
9 9 13 3 11 0 3 9 9 2
6 0 9 15 13 13 2
8 7 10 9 13 10 9 3 2
7 9 3 13 3 0 9 2
3 13 13 0
10 13 10 12 7 15 9 13 0 9 2
2 13 9
7 13 9 2 16 13 0 2
6 15 13 15 0 9 2
2 0 9
12 9 13 13 11 9 9 9 7 9 0 9 2
12 0 9 13 3 13 9 9 2 10 1 9 2
6 0 9 13 3 9 2
6 15 13 3 13 0 2
4 15 13 3 2
8 13 15 3 11 2 3 11 2
5 6 6 15 1 2
2 3 0
23 16 11 9 13 3 9 9 2 13 12 9 3 16 0 11 9 13 13 3 12 9 9 2
7 10 9 13 13 15 13 2
5 15 13 13 12 9
2 13 13
18 0 9 13 3 9 9 2 16 9 13 10 9 16 15 0 9 13 2
5 13 15 3 13 3
5 9 13 9 1 2
6 15 13 3 0 13 2
4 9 13 3 3
14 3 9 1 13 13 15 1 13 0 2 15 9 13 2
9 10 9 9 13 13 13 1 9 2
7 9 1 15 13 13 3 2
9 13 3 2 16 13 13 15 13 2
3 12 13 2
16 2 13 15 3 15 16 11 13 11 2 11 11 2 9 2 2
13 9 13 0 13 2 13 9 13 13 3 3 3 2
3 3 9 2
13 9 13 12 9 2 15 0 11 9 13 13 0 2
7 13 13 9 9 1 1 2
10 9 13 0 9 15 9 7 9 9 2
14 3 13 10 13 9 13 9 13 7 3 15 13 9 2
5 9 9 13 0 2
8 13 3 3 16 13 15 13 15
8 9 2 15 13 9 9 13 9
10 0 9 7 0 9 2 13 13 9 9
3 0 9 2
6 13 9 2 16 13 2
2 13 13
7 9 9 13 13 13 9 2
9 13 0 9 2 16 9 13 13 2
14 10 0 9 13 3 3 0 2 16 13 11 7 9 2
6 0 13 9 13 9 2
5 9 13 0 9 2
5 3 3 13 13 2
8 0 13 13 1 9 9 9 2
11 11 13 11 7 13 15 3 12 9 9 2
10 9 13 9 1 13 3 9 9 0 2
9 10 10 0 11 13 9 9 3 2
2 3 2
5 15 13 9 13 2
4 0 9 15 2
13 15 13 3 3 0 3 2 11 7 15 7 15 2
4 3 15 3 13
15 13 15 13 15 1 13 16 13 9 9 13 3 16 15 2
7 13 3 2 13 0 15 2
5 15 3 9 9 2
6 7 9 13 12 3 2
13 16 10 9 9 9 7 9 13 9 13 9 9 2
8 11 9 9 13 9 12 9 2
14 9 13 15 2 13 7 16 9 13 13 3 0 11 2
4 0 15 13 2
10 3 15 13 15 2 15 13 11 13 2
7 9 9 13 13 3 13 2
4 3 13 0 9
2 13 9
6 9 13 0 9 9 2
29 11 11 7 10 9 13 10 0 15 13 13 9 9 2 7 13 15 13 7 13 2 16 15 13 0 0 0 9 2
4 2 6 3 2
11 9 9 13 12 9 2 15 13 9 9 2
3 3 3 2
7 9 13 11 1 9 9 2
6 15 13 3 0 9 2
12 15 3 3 13 2 16 13 13 0 10 9 2
15 13 13 11 9 7 13 9 9 7 13 9 9 9 9 2
2 13 9
8 15 13 13 10 10 9 9 2
5 9 13 9 0 9
5 9 13 9 1 2
7 9 9 13 0 1 9 2
6 13 12 2 13 3 2
7 15 15 13 9 9 1 2
4 13 3 15 2
4 9 13 13 0
12 9 11 13 0 2 10 9 13 11 13 9 2
2 0 0
6 10 0 9 13 9 2
16 11 11 2 15 9 13 3 0 9 10 11 9 13 10 9 2
7 9 15 13 7 9 13 2
6 9 9 9 9 13 2
14 11 13 13 3 0 9 2 15 9 13 3 9 1 2
5 9 13 1 9 2
8 11 9 0 9 13 0 0 2
3 9 13 2
10 9 13 13 2 16 10 9 13 0 2
7 0 9 13 9 10 9 2
5 2 13 13 3 2
8 9 9 9 13 9 9 3 2
7 15 3 13 15 3 2 2
12 15 13 13 0 9 2 3 3 12 13 11 2
9 15 13 0 9 2 16 11 13 2
5 3 13 3 9 2
14 2 15 13 13 3 2 7 3 15 3 13 15 2 2
8 15 13 3 3 9 9 1 2
11 3 13 3 9 2 7 3 0 16 3 2
3 9 9 1
8 16 13 2 13 13 0 9 2
10 9 13 13 11 7 11 12 13 9 2
12 0 9 13 13 15 16 15 2 15 13 0 2
3 9 9 9
11 9 13 13 2 16 9 13 3 9 9 2
4 9 13 13 9
5 11 13 3 9 2
5 2 13 15 0 2
18 13 3 3 3 2 13 15 3 11 2 15 9 13 13 2 13 11 2
6 11 13 13 15 0 2
7 9 9 13 9 0 9 2
2 0 9
7 0 7 0 9 9 13 9
5 15 13 10 13 2
15 9 0 9 13 11 8 8 2 15 13 7 13 12 9 2
17 9 13 0 9 1 3 2 7 3 15 13 13 3 0 7 0 2
7 13 3 11 13 13 9 2
11 13 3 13 2 16 11 13 13 9 15 2
3 0 0 9
5 13 13 13 9 2
9 3 0 13 3 15 15 9 13 2
5 13 15 12 9 2
14 11 13 13 0 9 2 16 15 13 9 3 0 9 2
11 9 13 13 9 7 10 9 13 10 9 2
7 15 13 2 16 9 13 2
13 3 9 13 9 7 13 9 2 9 13 0 9 2
13 3 13 9 9 3 13 7 9 7 9 7 9 13
6 11 13 3 13 0 2
4 0 9 13 9
15 9 13 13 11 2 11 7 11 0 9 15 3 10 9 2
11 11 13 13 12 10 0 1 13 0 9 2
2 13 9
2 3 3
8 15 13 2 16 13 15 13 2
13 3 3 16 0 9 13 9 2 13 15 13 13 2
13 9 1 13 3 9 7 9 2 7 13 10 0 2
15 1 10 9 13 9 1 13 9 13 3 13 2 9 9 2
4 13 13 3 2
18 13 3 13 2 16 3 2 9 2 13 0 9 0 7 13 0 9 2
2 3 13
10 13 3 15 13 9 9 1 9 9 2
9 9 9 13 13 9 3 9 9 2
17 16 15 13 11 9 2 15 15 3 13 3 9 16 13 13 15 2
6 10 9 15 13 9 2
3 0 9 9
9 0 9 13 9 3 16 10 9 2
5 15 13 13 3 2
11 13 2 3 15 13 3 13 3 3 16 0
8 15 13 9 3 2 3 9 2
17 13 13 3 0 0 2 7 15 13 3 13 3 0 9 16 11 2
13 9 13 9 7 13 2 16 9 13 3 9 13 2
9 3 13 13 7 13 10 9 3 2
18 10 9 13 10 9 2 15 15 7 15 13 13 3 9 2 15 13 2
8 9 11 13 9 1 13 9 2
2 13 2
3 13 9 2
4 3 15 13 2
5 9 13 9 11 2
10 0 15 13 15 16 15 13 13 15 2
7 9 13 13 11 9 9 1
19 0 9 9 13 3 9 10 0 9 7 9 2 15 1 10 0 9 13 2
3 3 0 11
2 13 13
4 9 13 3 9
3 0 0 9
6 9 9 13 0 9 2
7 0 8 7 0 9 13 9
6 15 9 13 0 9 2
9 10 9 13 9 9 7 9 9 2
5 13 15 13 15 2
15 16 0 9 13 0 2 3 13 2 15 13 13 10 9 2
7 9 1 15 13 13 3 2
13 13 11 9 9 12 9 12 16 13 3 9 9 2
10 3 9 6 2 13 3 3 3 3 2
4 13 13 13 13
9 3 9 13 9 7 12 9 1 2
5 9 7 9 13 15
3 13 0 9
10 13 16 13 9 3 7 13 16 3 2
8 3 13 13 9 3 3 3 2
15 13 13 13 10 0 2 16 9 9 9 13 10 9 13 2
8 10 9 9 13 3 9 0 2
16 0 13 3 12 9 9 15 13 0 9 9 13 7 13 9 2
18 3 0 9 13 0 13 2 16 3 9 13 0 13 3 9 13 9 2
5 15 13 12 9 2
18 9 7 9 9 2 15 11 13 13 2 3 13 12 9 15 11 13 2
11 0 9 13 15 2 16 13 13 9 9 2
11 12 0 9 13 12 9 3 9 9 11 2
13 9 9 7 9 9 11 13 9 13 12 12 9 2
6 9 13 3 16 9 2
19 11 11 7 15 13 0 9 11 9 9 9 2 9 13 13 7 9 3 2
10 9 9 13 0 9 1 3 12 9 2
12 1 9 13 3 9 7 11 13 3 3 3 2
6 15 13 13 9 9 2
14 9 0 9 13 3 0 2 16 15 13 0 13 3 2
5 13 13 3 13 2
4 13 9 3 2
2 0 9
4 0 9 7 9
12 13 13 9 1 13 9 9 9 7 13 11 2
8 0 13 13 13 15 3 9 2
11 16 13 13 15 0 2 3 3 13 3 2
9 11 13 2 15 13 9 9 9 2
14 15 13 13 9 3 10 9 2 7 3 3 13 13 2
7 12 11 9 13 9 1 2
8 0 9 13 3 13 7 13 2
2 11 6
4 9 13 9 13
20 11 9 13 3 3 13 0 7 0 13 2 7 9 13 13 3 3 16 11 2
7 9 9 13 0 16 9 2
7 9 13 16 9 12 9 2
11 13 13 3 0 7 0 9 2 16 13 2
5 10 11 3 0 2
2 13 13
4 10 9 3 2
9 15 13 13 12 9 16 10 9 13
4 13 15 0 9
7 15 13 10 10 9 3 2
3 9 9 11
10 9 13 16 9 13 3 3 9 1 2
7 9 1 9 13 13 11 2
4 9 13 9 2
6 9 13 7 9 13 2
19 15 13 11 9 13 3 3 3 0 9 2 16 13 9 9 3 3 13 2
17 3 9 0 9 13 0 9 3 9 9 9 13 9 12 9 3 2
11 13 9 0 9 7 13 11 13 13 9 2
6 3 9 15 3 3 13
11 13 3 2 16 0 9 13 3 3 9 2
11 16 13 0 9 9 2 9 13 3 15 2
7 13 3 13 0 3 9 2
4 13 3 9 2
9 13 13 2 16 13 13 13 13 2
11 15 13 13 15 15 1 2 16 13 9 2
4 13 9 9 2
7 2 3 15 3 9 13 2
6 3 13 12 11 9 2
15 9 11 2 15 13 13 9 9 1 3 7 3 13 9 2
2 13 13
9 13 10 9 9 13 12 13 0 2
6 9 13 0 13 3 2
9 13 13 2 13 7 13 13 3 2
4 3 13 0 9
7 9 13 9 12 0 1 2
10 12 0 9 9 13 3 3 3 11 2
10 0 0 9 13 13 13 9 9 1 2
13 9 13 12 0 9 16 15 2 15 13 13 9 2
9 10 9 7 9 13 3 0 9 2
3 13 9 2
8 9 13 3 13 11 9 11 2
11 9 13 13 15 3 2 15 13 10 9 2
7 9 9 9 13 0 12 2
7 9 7 9 9 11 13 9
2 9 9
2 0 9
5 0 15 13 3 2
11 9 13 3 15 2 13 9 7 9 9 2
4 9 13 0 15
3 11 13 9
15 9 7 9 13 13 9 7 9 2 15 9 9 1 13 2
7 3 13 13 13 9 13 2
16 12 9 0 9 0 9 13 3 0 9 7 12 9 9 9 2
4 9 13 9 2
7 15 13 13 9 10 0 2
8 13 13 2 3 3 13 9 9
20 16 16 3 13 13 0 9 2 9 13 13 3 2 13 9 0 9 13 11 2
7 9 13 13 3 9 12 2
5 3 13 15 13 2
13 16 9 13 13 3 2 15 9 9 13 9 1 2
3 13 9 1
4 15 13 3 2
8 13 3 0 16 13 15 13 15
20 3 7 3 2 3 12 9 2 9 2 9 2 8 7 9 2 9 7 9 2
15 15 16 9 13 13 3 13 0 9 0 9 2 7 0 2
4 3 13 0 2
3 3 13 3
6 3 9 13 10 9 2
9 13 2 16 13 3 8 8 3 2
8 16 15 13 13 3 3 9 2
7 9 9 13 3 3 3 2
6 9 13 13 13 9 2
12 0 13 0 9 7 0 9 9 13 0 9 2
12 9 13 3 13 2 3 15 13 0 3 3 2
13 0 13 13 3 3 2 11 16 13 11 13 13 2
16 10 15 2 15 13 13 13 0 9 2 13 13 3 9 9 2
16 16 9 9 13 3 2 15 13 13 7 0 9 7 0 9 2
11 9 7 9 13 15 2 13 9 7 13 2
12 9 9 13 3 0 2 13 3 9 7 9 2
5 13 3 9 9 2
18 13 3 3 3 2 13 15 3 11 2 15 9 13 13 2 13 11 2
8 3 3 13 0 9 13 9 2
6 13 15 3 1 9 2
7 13 10 11 10 9 3 2
2 9 13
10 13 0 13 9 0 2 16 3 13 2
7 9 1 13 3 13 9 2
9 11 13 9 13 11 1 9 1 2
7 9 13 13 15 3 3 2
4 9 0 9 9
4 15 13 0 9
8 9 9 12 9 12 13 9 2
2 0 9
9 9 9 13 15 3 16 9 13 2
10 3 15 13 13 12 12 9 3 3 2
11 15 1 15 13 10 0 3 0 13 9 2
13 7 9 11 7 11 1 9 13 0 9 11 9 2
10 7 13 10 0 16 3 9 10 9 2
5 13 15 13 15 9
10 9 13 13 1 3 9 7 3 0 9
4 3 3 13 9
13 16 11 9 13 11 2 11 1 0 9 13 13 2
10 9 11 7 9 11 15 13 0 9 2
10 3 16 3 13 3 13 9 13 3 2
12 15 3 13 15 13 7 13 0 9 15 9 2
3 3 13 15
23 15 13 13 3 3 16 16 13 10 9 7 3 3 16 3 13 10 6 15 3 9 9 2
14 0 9 0 2 0 9 13 3 3 0 3 3 13 2
12 9 13 3 9 15 1 2 16 13 13 9 2
8 13 15 15 3 15 13 15 2
16 9 13 1 0 9 9 7 13 2 16 3 3 13 3 9 2
9 9 13 9 13 3 9 0 9 2
2 13 9
8 13 16 15 13 10 9 3 2
7 9 9 13 13 0 9 2
7 11 13 13 9 3 3 2
2 13 15
5 13 15 10 9 2
20 12 9 0 9 11 13 0 9 9 12 7 13 13 9 9 12 0 7 0 2
8 10 9 9 0 11 9 13 2
5 0 9 13 9 2
12 2 3 15 10 9 13 2 2 9 13 9 2
6 15 13 13 3 3 2
4 9 1 13 9
9 0 9 13 9 7 0 0 9 2
7 9 13 15 2 16 13 2
3 13 9 9
14 13 13 13 3 9 2 16 9 13 11 9 0 9 2
11 9 13 9 1 9 7 13 3 9 2 2
11 9 9 9 11 11 1 9 13 11 9 2
5 15 15 3 13 9
8 9 0 11 9 13 3 11 2
17 3 15 13 10 9 3 11 3 15 1 15 13 16 15 13 13 2
4 2 13 13 2
9 13 2 16 13 9 13 3 13 2
10 13 2 16 13 10 3 11 13 11 2
4 15 13 15 2
7 3 15 13 13 0 9 2
10 9 13 9 13 3 0 7 0 13 2
16 3 15 13 3 15 9 13 3 13 15 13 3 0 10 3 2
6 3 15 15 1 13 2
13 9 13 13 13 3 10 9 16 15 13 9 7 2
10 3 12 9 1 11 13 0 9 0 9
10 3 9 7 10 10 9 13 13 9 2
4 2 3 13 2
6 15 13 3 9 0 2
6 15 13 13 0 9 2
10 9 13 13 3 3 13 13 3 9 2
16 7 9 13 3 16 16 15 15 13 2 3 9 9 13 13 2
6 13 15 3 13 9 2
11 11 13 13 13 9 13 3 11 11 9 2
11 3 13 3 9 7 3 9 13 3 0 2
2 9 11
10 9 13 9 0 9 7 13 9 9 2
6 0 15 13 0 9 2
3 13 3 2
4 9 7 9 1
4 3 15 13 2
3 15 13 13
14 9 9 13 3 3 9 9 2 9 7 9 9 9 2
16 3 9 12 1 15 13 13 3 3 2 16 13 13 3 13 2
10 15 13 3 13 2 16 15 13 3 2
6 3 9 13 3 3 2
5 15 13 15 3 2
6 15 13 3 0 9 2
17 11 13 15 13 3 3 3 10 0 3 0 9 10 0 3 9 1
9 10 0 9 9 13 13 9 9 2
3 13 0 9
5 10 9 15 13 9
5 13 15 3 9 2
3 3 13 9
6 0 0 9 13 13 2
7 11 13 11 9 7 9 2
5 15 15 13 0 9
2 11 9
9 3 15 13 13 3 3 9 1 2
9 16 13 13 2 13 9 3 13 2
12 2 13 12 9 9 16 13 13 3 9 2 2
24 15 13 13 9 0 9 2 15 13 3 11 11 9 15 13 9 7 9 15 9 15 13 3 2
10 11 11 9 9 2 2 3 13 3 2
12 3 9 13 10 9 2 16 13 12 9 9 2
2 9 9
7 7 3 15 15 3 13 9
6 15 13 15 13 9 2
10 9 13 12 2 13 9 7 13 13 2
7 0 9 9 13 0 0 2
3 13 15 2
3 9 9 2
4 9 13 9 2
6 9 13 13 0 9 2
12 15 13 3 9 7 15 13 9 9 9 3 2
26 3 3 13 13 3 3 7 13 9 7 13 9 7 13 3 10 9 3 2 9 7 15 13 13 9 2
13 15 13 13 9 7 10 0 7 15 13 15 9 2
4 9 7 9 9
12 9 3 2 16 13 3 13 9 7 13 9 2
23 9 13 10 10 9 2 15 10 9 13 3 2 7 0 9 13 2 16 9 13 9 13 2
4 13 13 13 2
17 8 8 8 8 8 8 7 11 11 8 13 3 0 16 11 9 2
2 10 9
7 10 9 10 9 13 13 2
4 9 13 9 2
7 0 13 3 13 0 9 2
6 11 7 11 13 0 9
7 11 9 9 13 3 11 3
8 10 11 9 9 13 13 9 2
5 9 13 3 13 3
10 13 10 11 2 15 13 3 1 15 2
17 13 3 11 7 11 7 15 2 15 13 9 7 9 9 10 3 2
2 3 13
32 11 9 13 0 9 9 12 9 2 11 11 0 0 9 10 9 2 11 9 7 9 13 13 12 9 2 11 9 12 9 3 2
5 0 9 3 9 2
41 9 13 9 9 0 9 2 9 9 2 9 7 10 0 2 9 11 2 9 9 2 9 11 1 9 9 2 9 9 9 1 7 3 9 9 3 10 0 9 9 2
6 9 1 13 0 9 2
12 9 1 13 3 15 2 13 9 3 7 11 2
7 0 0 13 10 0 9 2
8 15 13 12 2 12 7 11 2
4 13 3 13 2
5 9 13 3 9 1
6 9 13 13 10 0 2
4 13 15 3 2
6 3 15 13 13 13 2
6 3 13 9 0 9 2
9 13 13 8 11 1 3 11 1 2
4 13 15 13 2
3 13 0 2
3 13 9 2
8 9 13 3 10 9 15 13 2
7 9 13 0 9 9 9 2
6 9 13 9 13 3 2
6 9 13 13 9 13 2
10 11 3 2 15 13 9 12 12 9 2
12 0 9 13 0 13 2 16 9 13 13 9 2
10 3 12 9 13 11 7 11 0 0 9
2 9 0
15 9 13 13 3 2 15 13 9 0 15 15 9 1 13 2
10 13 15 11 2 3 13 13 9 9 2
4 0 0 0 9
7 0 9 13 12 9 12 2
13 3 11 13 9 3 8 7 9 16 10 10 9 2
6 7 13 3 10 9 2
19 11 13 9 11 0 9 0 11 2 15 9 13 13 3 13 9 13 3 2
13 15 13 13 3 3 3 15 13 10 0 9 9 2
2 6 6
9 9 13 0 2 7 9 13 0 2
7 13 3 9 9 1 1 2
6 7 9 13 13 15 2
2 13 13
10 11 9 13 0 2 7 13 3 0 2
7 9 1 15 3 13 9 2
24 15 13 13 3 2 16 13 3 2 15 3 13 7 3 2 16 13 2 0 0 9 13 3 2
7 9 13 13 9 7 9 2
7 15 1 13 13 3 13 2
14 12 15 13 9 7 9 2 9 15 3 3 12 12 2
12 9 13 11 7 13 3 0 9 0 12 9 2
7 15 13 3 9 15 3 2
9 3 2 7 9 13 3 0 9 2
18 0 15 3 13 2 9 13 2 7 15 3 13 9 9 7 9 9 2
6 3 13 3 13 9 2
2 9 2
13 0 9 9 9 13 3 13 13 0 9 9 9 2
6 3 0 11 13 9 2
9 13 15 3 2 3 13 0 9 2
5 9 13 13 3 2
13 6 9 15 13 3 2 15 13 13 9 6 3 2
10 11 13 13 0 9 9 0 10 9 2
3 10 12 9
10 9 9 13 0 9 9 9 13 9 2
8 13 0 2 16 15 13 13 2
8 11 9 9 13 13 11 11 2
12 16 15 13 13 0 2 3 15 13 13 3 2
12 11 1 9 13 13 2 16 13 15 13 13 2
12 6 3 12 10 9 13 9 7 15 13 13 2
7 9 9 13 10 9 9 2
7 15 13 0 9 13 9 2
7 13 3 3 10 3 9 13
2 10 9
2 9 9
7 15 13 3 3 0 13 2
9 13 9 10 9 2 15 15 13 2
10 11 13 9 15 13 0 9 2 0 2
7 9 13 13 13 3 0 9
17 16 13 9 12 0 9 3 2 16 13 13 13 15 2 13 9 2
6 9 11 9 12 1 2
7 9 0 9 13 0 9 2
10 13 9 9 2 16 13 3 13 9 2
5 9 9 13 9 2
11 15 13 0 2 15 13 3 13 9 15 2
9 15 13 3 13 2 16 15 13 2
19 13 13 3 9 2 16 13 3 0 9 0 9 2 15 13 0 9 9 2
4 13 9 13 9
18 9 2 9 7 9 13 3 3 3 0 9 16 10 0 0 0 9 2
11 15 13 3 11 2 16 3 3 15 13 2
27 7 10 9 7 9 3 15 1 15 13 3 0 9 3 13 13 3 3 10 9 3 3 10 10 9 13 2
4 11 13 9 2
11 13 11 0 9 11 13 10 9 3 9 2
15 11 13 3 2 7 13 15 3 0 9 16 3 11 11 2
2 13 3
8 7 13 3 13 13 3 9 2
6 7 3 15 15 13 2
21 11 13 13 3 0 3 7 9 7 0 15 2 16 13 13 0 0 9 2 11 2
3 0 12 9
5 13 15 13 9 2
6 3 13 13 3 13 2
15 11 13 13 11 3 12 9 12 9 2 16 15 13 9 2
7 11 9 9 13 11 0 2
5 13 13 9 9 2
18 11 13 13 9 9 2 15 13 9 1 13 3 3 16 9 13 3 2
6 13 13 3 3 13 3
4 9 13 3 13
3 13 9 2
4 9 13 9 2
19 9 9 12 9 13 12 2 12 2 12 2 12 2 12 2 12 7 12 2
35 3 15 13 3 0 13 16 13 15 15 13 13 15 13 13 3 3 16 13 13 0 9 16 13 15 3 3 13 16 15 13 15 13 9 2
5 9 13 13 9 2
7 11 13 9 7 15 13 2
6 0 13 3 0 13 2
4 9 13 9 2
8 0 9 13 13 13 9 3 2
8 9 13 3 9 9 3 3 2
8 15 13 0 9 13 9 9 2
2 3 3
5 10 9 13 13 2
8 10 0 9 13 15 13 0 9
12 10 0 10 9 13 11 13 7 13 3 9 2
5 15 15 13 9 2
14 9 13 3 3 13 15 2 16 15 13 9 9 3 2
7 9 13 10 9 3 9 2
6 11 13 9 0 9 2
5 9 9 13 12 2
10 9 2 15 13 15 2 13 9 13 2
6 13 15 13 0 9 2
4 15 15 13 2
4 0 16 9 15
10 10 9 15 13 2 15 13 13 9 2
8 16 3 13 2 13 15 3 2
21 11 13 16 15 13 13 11 7 11 0 9 10 9 2 16 15 13 10 9 13 2
6 0 9 13 3 11 2
7 3 10 9 13 3 9 13
6 0 9 13 9 9 2
15 9 11 13 13 3 9 9 1 2 16 0 9 13 9 2
3 9 13 2
2 0 9
9 6 3 2 13 11 13 15 9 2
16 0 9 2 3 9 13 13 7 13 9 2 7 9 13 13 2
4 13 15 9 2
3 9 12 9
2 3 16
13 9 13 16 9 7 13 3 2 13 3 0 9 2
4 15 13 13 0
2 9 9
3 9 13 13
10 9 13 15 3 2 16 15 13 13 2
11 9 13 9 0 9 9 13 15 15 0 2
13 13 13 10 9 13 16 13 15 13 11 10 9 9
5 9 13 9 1 2
6 13 0 13 3 9 2
9 9 7 9 9 13 13 0 0 2
9 15 13 13 13 15 13 13 15 2
9 13 13 2 16 9 15 3 13 2
7 0 9 13 13 3 0 2
7 13 13 3 13 0 9 2
16 9 9 9 13 12 0 9 10 10 9 2 15 15 13 13 2
6 0 9 13 13 15 2
14 13 9 13 13 7 0 9 2 9 13 9 7 9 2
14 9 13 13 9 2 15 1 9 13 13 3 9 1 2
3 9 9 13
10 11 13 11 1 9 13 9 9 11 2
7 13 9 13 9 12 9 2
3 15 13 2
13 9 13 3 0 3 9 9 7 9 9 7 9 2
7 3 15 3 13 0 9 2
6 15 13 9 3 3 3
10 3 12 0 9 13 3 13 3 3 2
4 9 13 9 2
10 9 13 13 9 12 9 3 12 9 2
5 16 13 9 13 9
14 9 11 13 13 9 13 0 9 9 3 9 12 1 2
7 3 13 9 13 11 9 2
16 11 13 0 9 2 13 15 0 9 3 16 10 10 9 9 2
7 13 13 13 3 0 9 2
7 0 9 13 3 0 9 2
15 0 9 13 3 3 13 0 9 8 2 15 3 13 9 2
12 9 7 9 13 0 13 10 9 2 9 13 2
9 13 15 2 15 13 9 0 0 2
6 9 13 3 9 0 9
16 16 13 3 0 9 2 0 9 2 13 15 13 3 0 9 2
4 13 15 3 2
9 9 13 3 7 3 13 15 13 2
4 15 13 3 3
4 11 11 1 11
5 13 13 15 13 9
21 13 9 13 3 12 9 2 15 12 13 3 9 2 12 3 13 9 7 12 15 2
17 3 15 13 3 16 6 6 9 16 13 15 13 10 9 3 13 2
4 15 13 13 2
15 11 9 13 3 12 9 9 2 16 15 11 13 12 9 2
2 12 9
21 15 13 3 3 3 2 15 0 13 11 2 15 13 13 7 15 15 13 9 13 2
10 11 13 13 13 9 3 9 3 9 2
6 9 13 3 11 9 2
3 13 3 2
7 15 13 0 12 9 1 2
5 13 15 13 9 2
4 11 13 9 2
5 11 13 9 13 9
3 9 0 9
14 9 2 15 11 3 13 10 9 1 11 13 13 9 2
6 9 9 13 0 9 2
4 9 13 15 3
13 0 9 9 13 12 7 10 9 9 13 3 12 2
8 9 13 15 3 10 0 9 2
3 15 13 9
7 9 13 0 9 9 11 2
7 3 11 9 0 9 0 9
2 9 9
4 15 13 12 9
6 3 15 13 10 9 2
16 15 13 13 3 3 10 9 10 0 9 13 7 10 9 13 2
3 2 15 2
8 10 9 11 9 13 9 9 2
2 6 15
9 15 13 3 9 2 11 13 9 2
10 15 1 15 15 13 2 13 15 3 2
2 6 3
3 9 0 2
7 11 9 13 11 9 0 2
10 9 7 9 13 11 9 9 0 9 2
6 9 13 9 13 0 2
7 9 13 13 3 7 3 2
3 15 1 16
11 9 0 7 3 13 13 3 13 9 9 2
6 0 9 3 0 9 2
2 9 0
6 9 13 9 13 3 2
20 15 1 9 9 13 13 13 10 9 9 1 2 3 9 13 9 12 9 9 2
6 15 13 13 10 9 2
2 0 9
10 15 13 3 3 9 0 9 9 1 2
10 9 13 3 0 2 16 13 3 0 2
7 9 13 9 0 9 9 2
11 9 1 9 13 15 16 9 13 13 9 2
13 9 13 13 0 2 15 9 13 9 10 9 13 2
5 9 13 0 13 2
4 9 13 13 2
11 3 3 11 13 3 13 9 7 11 9 2
8 13 13 3 12 7 3 12 2
2 9 13
10 7 3 13 9 13 13 2 3 9 2
10 9 12 8 7 9 13 12 9 9 2
4 0 2 0 9
17 13 3 9 2 16 9 13 3 0 9 2 7 13 15 11 3 2
4 15 13 11 2
2 9 9
11 13 15 11 9 13 9 15 10 9 13 2
6 9 13 13 9 1 2
7 3 13 10 12 9 13 2
6 13 9 9 9 1 2
6 2 13 13 3 9 12
18 7 16 15 13 13 9 2 15 13 15 3 9 2 3 16 13 15 2
7 9 13 13 3 0 9 2
12 9 13 3 3 12 0 9 2 0 0 9 2
14 16 13 9 11 9 13 10 9 13 11 13 10 9 2
4 9 13 11 2
9 3 15 13 15 0 9 3 6 13
15 3 13 11 9 3 0 7 3 0 2 0 0 9 9 2
16 15 2 15 9 13 2 13 15 13 7 15 13 15 3 0 2
16 12 9 9 13 3 9 9 7 9 13 9 9 7 9 9 2
10 9 13 11 11 2 0 9 9 9 2
8 13 3 11 9 12 9 9 2
11 11 7 11 13 9 13 3 3 9 9 2
15 0 3 13 2 16 11 7 9 9 13 10 9 13 3 2
5 13 15 15 3 2
5 15 13 15 9 2
5 13 13 3 13 11
17 16 9 9 13 13 10 3 9 2 3 0 9 13 13 10 9 2
15 12 9 1 9 13 9 9 15 2 16 9 13 15 13 2
3 6 15 2
8 7 13 3 7 9 13 3 2
11 10 9 13 13 13 13 10 0 9 9 2
18 11 3 13 16 13 16 13 3 0 9 3 9 1 3 13 15 13 2
10 9 13 9 2 13 0 2 0 15 2
10 3 9 13 7 3 15 13 3 13 2
4 6 3 0 2
7 9 13 3 15 1 9 2
5 13 9 7 9 2
11 15 13 9 13 9 13 12 0 9 9 2
3 12 9 0
9 11 9 9 7 9 13 3 0 2
5 13 10 9 9 2
17 9 13 16 0 9 2 12 9 2 2 7 9 9 13 3 0 2
15 10 9 13 13 9 12 9 2 3 16 3 2 7 12 2
4 9 7 9 9
6 15 13 3 12 9 2
9 13 0 16 13 9 2 15 13 2
12 9 13 9 0 9 7 13 9 9 16 9 2
2 3 9
5 9 13 9 1 2
2 9 0
5 13 15 13 13 2
17 0 9 15 3 13 9 11 0 9 2 15 3 13 0 9 0 2
9 9 13 2 16 3 13 10 9 2
9 13 15 0 9 9 16 9 9 2
13 13 9 2 16 13 0 0 9 13 3 15 1 2
5 0 11 13 9 1
4 9 1 13 9
8 13 0 9 13 9 3 9 2
13 9 13 9 2 16 9 13 13 15 9 13 9 2
15 9 13 0 9 2 16 15 13 3 13 0 9 0 9 2
14 7 9 15 13 2 16 13 3 13 2 16 13 9 2
5 11 13 3 9 2
15 7 13 15 13 10 9 13 9 12 9 11 13 0 9 2
4 11 3 13 9
6 15 13 13 9 13 2
7 0 0 10 0 9 13 2
7 9 13 13 10 9 9 2
10 9 13 15 13 3 9 13 0 9 2
4 13 11 10 9
9 11 13 0 0 2 15 13 13 2
3 0 13 2
6 15 3 13 13 15 13
5 9 13 9 13 13
7 13 16 15 13 13 15 2
9 9 12 11 13 11 9 12 9 2
3 15 13 9
2 10 9
10 9 9 13 3 13 9 13 3 9 2
3 13 9 9
3 15 13 0
2 3 13
16 9 9 9 13 12 9 2 7 15 16 0 2 9 2 11 2
13 3 15 13 13 3 2 15 13 13 9 9 13 2
11 13 9 9 13 13 3 12 9 9 9 2
7 13 15 3 13 13 9 2
12 9 11 9 13 3 9 2 16 9 13 9 2
8 9 11 9 13 9 3 12 2
7 13 3 9 3 15 1 2
13 0 0 13 16 9 13 3 2 16 15 13 9 2
14 3 11 13 2 13 15 0 9 9 2 9 7 9 2
16 0 9 13 3 2 16 3 9 9 11 11 13 13 9 1 2
10 3 15 13 13 3 2 15 13 3 2
4 3 3 15 2
2 11 9
11 9 13 9 0 9 2 15 0 13 9 2
14 11 13 13 12 9 9 12 2 15 13 12 9 9 2
6 13 9 9 2 6 2
4 13 9 1 2
5 3 13 3 0 2
13 9 13 13 9 7 10 0 9 2 15 13 13 2
7 10 9 0 9 13 9 2
9 15 13 9 1 7 13 9 9 2
2 3 2
5 15 13 13 11 2
8 13 0 2 16 15 13 13 2
5 15 13 3 3 2
7 10 9 13 13 0 9 2
3 9 9 2
9 3 13 9 2 15 13 0 3 2
14 2 9 2 13 9 13 0 9 2 15 13 13 3 2
3 0 13 9
7 13 9 9 9 7 9 2
15 13 9 9 1 7 3 0 13 2 16 9 13 3 9 2
8 11 10 9 13 0 7 0 2
4 13 3 9 2
10 9 13 16 9 11 9 7 11 13 2
2 9 9
4 9 13 13 13
20 7 3 10 12 10 9 2 0 9 7 9 9 9 1 2 13 9 7 9 2
9 7 13 3 8 7 11 13 9 2
12 0 9 1 9 13 3 13 9 0 9 9 2
12 9 12 11 9 13 2 7 9 13 13 13 2
2 13 9
12 15 11 13 13 9 15 2 15 13 3 0 2
17 16 11 9 13 2 13 0 9 2 16 3 16 13 13 11 3 2
14 11 9 13 2 16 9 13 13 1 9 3 11 9 2
10 13 15 13 2 16 13 9 13 15 2
5 13 3 3 9 2
5 3 15 13 3 2
5 9 13 9 1 2
16 9 13 13 11 9 3 2 7 10 9 13 9 9 9 13 2
4 9 13 9 2
8 7 10 12 9 1 13 13 2
13 15 3 13 13 9 2 3 9 7 0 13 13 2
7 9 11 13 0 9 3 2
11 11 11 2 15 13 9 9 7 10 9 2
15 13 3 3 7 3 13 13 3 3 16 13 2 9 13 2
8 15 3 13 13 0 9 9 2
5 15 13 9 15 2
6 9 1 9 13 9 2
14 13 13 1 9 10 9 2 7 1 9 3 10 9 2
5 15 13 15 3 3
5 13 0 7 13 2
10 9 1 13 9 13 13 9 3 9 2
10 10 9 13 9 9 9 7 9 1 2
7 13 13 3 16 3 13 2
15 3 9 13 0 16 15 9 9 12 9 9 13 9 13 2
3 2 13 2
4 15 13 15 3
4 13 13 10 9
22 7 16 15 3 13 13 10 0 0 9 2 13 3 15 2 16 15 13 10 0 9 2
8 13 15 3 13 7 13 15 13
9 9 13 9 7 12 9 13 15 2
5 9 13 9 9 2
8 15 13 12 9 1 13 9 2
8 9 13 9 1 9 13 9 2
7 13 13 16 13 9 13 3
7 16 13 3 3 13 3 2
10 9 9 13 9 13 13 13 3 13 2
8 15 13 3 13 13 13 13 9
11 9 2 15 9 13 0 2 9 13 0 2
2 13 15
4 13 9 1 2
7 0 9 13 9 9 13 2
4 15 3 13 2
2 13 11
6 7 3 13 3 9 2
5 9 13 13 3 2
15 13 10 9 13 2 16 9 15 13 15 10 9 3 13 2
19 16 13 9 7 13 9 13 11 2 3 3 3 13 2 16 3 15 13 2
13 15 3 15 13 16 10 9 15 13 3 3 3 9
7 0 9 13 3 13 3 2
6 9 13 9 13 9 2
20 11 13 9 1 13 3 9 2 7 2 3 15 13 2 0 9 13 9 9 2
13 15 9 13 0 9 2 15 13 13 0 0 9 2
6 13 3 16 13 13 2
3 13 9 2
6 9 13 9 9 0 2
4 15 15 13 13
8 15 13 3 3 0 9 3 2
15 15 13 13 3 10 9 1 2 15 9 1 13 15 9 2
13 7 15 13 3 15 1 16 11 13 13 12 9 2
3 13 0 2
6 10 0 15 3 13 2
5 12 9 13 9 2
4 9 13 1 9
6 15 13 13 9 3 2
10 11 11 11 13 13 9 11 0 9 2
2 0 9
3 9 13 2
5 3 15 13 9 2
2 9 1
8 0 9 13 9 2 15 13 9
10 15 3 13 2 16 13 13 15 15 2
11 16 15 13 9 2 3 15 13 15 13 2
3 3 9 2
4 13 10 9 2
12 3 13 2 16 13 15 13 2 9 3 13 2
8 9 9 13 10 9 0 0 2
10 15 13 2 16 15 3 9 13 0 2
18 9 13 13 13 9 9 15 13 3 2 7 16 15 13 9 3 9 2
6 2 11 13 3 10 9
5 13 9 9 11 2
11 3 9 9 13 15 3 9 7 9 9 2
14 9 13 9 2 10 9 9 2 15 13 9 9 1 2
2 0 9
13 0 9 13 11 3 3 9 16 0 9 3 9 2
14 9 9 0 0 7 0 0 8 8 8 13 0 9 2
8 3 13 15 13 9 9 11 2
4 0 9 7 9
3 9 13 9
9 3 9 7 9 13 3 2 16 2
5 13 13 15 3 2
45 16 3 15 13 3 9 7 3 15 13 16 3 13 3 3 15 16 6 16 15 3 13 3 15 0 9 3 3 15 13 3 16 6 16 16 3 15 3 13 16 13 15 13 10 9
3 13 9 2
6 13 9 13 9 13 2
4 9 2 9 11
6 13 13 3 7 3 2
12 3 13 13 13 3 0 15 2 15 9 13 2
5 15 13 3 0 3
4 9 13 9 2
12 9 16 13 9 2 3 9 9 13 13 9 2
13 11 1 11 13 10 9 7 13 9 1 0 9 2
11 13 3 13 10 9 3 0 9 0 11 2
5 0 13 3 9 2
6 9 13 3 9 7 9
2 3 9
8 11 9 13 3 9 1 0 2
5 9 13 13 1 9
2 9 13
5 9 13 9 1 2
7 15 13 3 13 12 9 2
14 10 9 9 13 10 9 2 12 0 2 9 13 9 2
4 15 13 3 13
19 9 13 0 9 2 9 9 1 7 3 16 13 0 9 13 0 0 9 2
6 15 13 3 0 9 2
17 11 13 2 16 0 9 7 0 9 13 2 16 9 13 11 9 2
10 9 13 9 12 9 9 2 9 2 2
3 9 13 9
11 11 7 11 11 13 9 13 12 0 0 2
5 11 13 3 9 2
12 9 13 13 9 2 15 13 13 11 0 9 2
4 15 13 13 3
8 8 7 9 13 11 11 1 2
6 13 3 15 0 9 2
7 10 0 9 13 0 9 2
7 15 13 15 3 13 9 2
2 0 9
4 9 13 0 2
6 15 1 9 13 3 2
6 12 9 15 13 0 2
16 9 13 12 9 1 2 7 13 3 12 9 2 9 13 12 9
14 15 13 13 9 2 7 10 9 11 0 9 3 9 2
20 9 15 13 13 10 9 13 9 10 9 15 10 10 0 8 7 9 13 11 2
7 10 9 13 13 13 9 2
6 15 13 0 9 9 2
5 13 0 9 0 2
7 10 9 13 3 0 9 2
7 9 13 9 7 13 15 2
6 13 0 7 13 9 2
9 0 9 11 13 9 9 0 9 2
13 9 13 11 9 13 9 2 16 9 13 13 3 2
3 3 13 9
4 9 13 9 2
14 9 13 10 9 13 9 9 2 13 15 3 0 3 2
11 9 9 13 9 1 2 16 13 9 13 2
10 6 7 15 13 13 9 16 15 13 2
16 0 1 13 13 2 13 7 13 3 10 9 1 0 9 9 2
2 13 13
10 9 9 13 13 3 10 12 0 9 2
12 11 0 9 9 7 9 13 13 2 3 2 2
7 3 10 10 9 13 3 2
7 0 9 9 13 0 0 2
8 9 10 9 9 1 13 9 2
21 10 9 13 9 12 13 9 9 9 7 0 9 13 9 9 7 9 9 7 9 2
5 11 9 13 13 2
4 9 0 9 9
11 9 13 13 11 0 9 13 3 12 9 2
7 13 9 9 7 13 9 2
14 9 16 13 9 9 9 2 10 9 13 12 0 9 2
7 9 13 3 16 9 0 2
8 7 13 13 13 16 13 13 2
11 9 13 3 0 15 2 15 0 13 9 2
12 15 13 10 9 0 9 16 3 13 3 9 2
12 9 13 13 9 2 9 7 9 13 3 9 2
12 10 15 13 13 9 2 3 0 13 16 9 2
7 12 3 0 9 3 13 13
3 13 13 13
6 13 13 9 12 1 2
5 9 13 0 13 9
7 9 13 9 3 15 0 2
19 11 2 11 10 9 9 13 0 9 2 15 13 9 11 11 7 0 11 2
6 13 15 15 15 13 2
10 15 1 13 13 13 16 15 13 9 2
3 9 9 2
16 9 13 3 13 13 9 7 9 2 13 15 13 3 13 9 2
3 13 3 13
5 9 13 13 9 2
5 9 13 0 9 2
5 9 13 13 13 2
10 9 9 13 2 16 13 15 13 11 2
24 0 7 0 9 0 9 13 15 9 3 0 2 16 13 9 11 7 11 1 10 9 13 9 2
2 13 15
2 0 9
4 13 15 3 2
14 9 13 9 9 9 2 13 9 0 0 15 15 13 2
8 13 3 3 2 16 15 13 2
8 9 11 13 9 11 0 9 2
5 9 9 7 9 1
3 3 0 9
8 3 13 9 13 9 16 13 2
7 15 13 3 3 16 9 2
6 9 13 0 13 3 2
30 9 13 13 2 16 13 0 7 0 9 9 9 2 7 15 13 13 0 7 0 3 9 2 16 3 13 12 9 3 2
9 3 16 13 15 2 15 9 13 2
8 9 13 0 9 9 0 9 2
6 13 13 0 9 9 2
7 11 13 9 3 9 9 2
5 13 15 15 13 2
11 7 3 10 9 13 11 9 13 9 13 2
5 11 9 13 9 2
9 13 9 3 3 7 3 7 3 2
3 11 13 13
16 0 2 15 3 13 7 3 13 13 13 3 3 15 13 9 2
12 15 13 3 3 9 16 3 10 9 3 13 2
7 0 13 0 12 9 1 2
17 9 11 13 0 9 2 9 13 0 9 13 2 9 3 9 13 2
9 7 13 2 16 15 13 0 9 2
11 15 13 0 9 16 13 0 2 15 13 2
12 10 9 13 2 0 2 0 2 3 9 9 2
8 15 13 13 3 0 16 15 2
5 15 3 13 15 2
11 9 13 0 0 7 3 9 13 0 13 15
13 13 3 16 13 11 13 0 16 15 0 13 13 2
10 9 9 13 3 3 3 16 0 9 2
7 13 15 15 13 9 13 0
7 0 9 13 9 9 3 2
4 13 15 3 2
5 15 13 3 3 2
7 9 0 9 13 12 9 2
2 9 3
3 8 7 9
11 15 13 2 16 15 13 13 15 9 9 2
6 13 12 7 13 12 2
15 15 1 15 13 13 3 9 2 16 9 13 3 3 12 2
13 15 13 13 10 9 15 13 9 9 0 9 9 2
2 13 9
4 9 13 13 0
2 9 2
12 7 11 9 7 0 9 1 9 13 13 13 2
16 13 0 9 0 7 13 2 13 9 2 15 3 3 13 13 2
18 10 11 9 3 15 13 3 0 16 15 13 16 15 3 13 15 9 2
7 0 9 13 13 3 3 2
3 13 13 15
15 0 13 9 13 11 7 11 9 2 3 9 13 13 9 2
3 15 13 2
9 11 13 15 0 9 9 3 3 2
7 9 13 13 9 13 9 2
15 11 9 13 9 2 16 9 13 3 0 2 9 13 9 2
6 15 15 13 13 9 2
6 9 9 2 9 7 9
6 9 13 13 13 9 2
2 0 9
5 9 13 9 1 2
4 13 9 0 9
6 9 13 12 12 9 2
3 13 3 2
14 15 13 15 2 3 13 0 2 9 0 9 9 7 9
4 13 15 9 2
7 13 3 10 9 3 3 2
6 15 13 13 0 9 2
8 3 13 13 11 2 11 13 2
8 11 7 11 13 3 3 9 2
7 10 9 9 13 3 11 2
12 9 9 13 9 1 7 0 9 0 9 9 2
36 6 2 15 15 3 13 15 15 13 9 12 9 16 12 9 1 7 2 15 13 15 13 3 3 7 3 10 9 13 15 15 13 3 16 3 3
6 10 9 9 13 0 2
10 15 13 10 9 2 15 13 13 9 2
10 3 13 3 3 9 7 9 13 13 2
2 10 9
12 13 9 1 0 9 2 3 12 9 13 9 2
5 15 15 3 13 2
8 16 13 13 13 9 13 9 2
2 9 13
9 9 13 9 10 9 2 9 7 9
6 13 3 15 13 13 2
7 9 13 13 12 12 9 2
5 10 9 13 3 2
13 9 11 7 9 9 13 0 2 15 11 13 13 2
15 13 10 9 3 2 13 13 3 2 7 13 10 9 3 2
6 9 9 13 10 9 2
7 9 9 13 3 9 9 2
17 16 15 3 3 13 13 2 3 3 0 3 2 9 16 13 9 2
4 13 15 9 2
6 13 3 15 7 13 13
4 13 13 3 2
8 9 9 13 9 10 9 3 2
8 11 0 9 13 13 0 9 2
12 16 9 9 13 13 0 2 15 13 3 0 2
12 3 13 3 13 9 13 16 9 13 13 3 2
16 11 13 0 9 2 15 3 13 13 9 11 13 13 9 9 2
11 12 9 0 15 13 13 9 0 9 1 2
9 13 15 13 3 10 9 2 9 2
5 15 13 9 0 2
20 15 9 13 3 3 13 15 2 3 10 0 1 3 13 13 3 9 13 9 2
4 9 13 9 2
3 13 12 2
4 13 3 9 2
5 9 13 9 9 2
6 9 13 13 9 1 2
23 15 13 13 13 13 10 0 2 7 10 9 13 15 9 0 3 10 9 7 15 13 15 2
19 13 13 9 3 3 2 16 13 0 9 2 13 3 0 9 9 11 11 2
6 13 13 3 0 0 2
10 9 15 13 3 13 2 7 3 9 2
13 11 9 13 2 16 9 9 13 9 9 13 9 2
2 13 13
12 9 9 13 3 0 2 3 3 9 7 9 2
2 3 0
2 9 13
9 0 9 13 3 0 16 10 9 2
