241 11
35 15 10 9 10 9 14 13 3 14 13 15 10 9 10 0 9 1 9 3 10 9 9 1 9 0 9 13 7 14 13 1 10 0 9 2
10 10 9 9 13 10 9 9 1 9 12
42 10 0 9 2 1 15 13 10 9 10 9 2 9 9 2 7 10 3 9 10 0 9 2 9 9 2 13 10 9 1 9 1 9 9 10 9 9 9 9 1 9 2
4 0 0 9 2
9 0 1 15 13 14 13 0 2 2
18 13 14 13 10 0 9 2 7 10 9 2 13 1 10 9 2 13 2
21 3 2 10 9 10 1 3 9 2 10 9 7 10 9 15 13 10 3 0 9 2
45 3 2 3 13 10 9 10 2 9 2 14 13 14 13 10 9 15 3 1 15 3 7 1 0 10 9 10 9 1 10 9 15 13 1 9 7 9 3 1 10 3 0 15 9 2
15 10 9 13 10 0 9 10 9 7 13 1 3 10 9 2
39 10 9 12 9 14 13 14 13 1 10 9 9 9 2 3 1 10 15 10 9 13 1 12 2 12 2 12 1 1 12 2 12 2 12 2 12 2 12 2
42 13 10 0 9 0 1 10 3 9 7 13 7 3 14 13 7 10 9 1 10 9 9 2 7 1 10 9 15 3 10 0 9 14 13 10 0 9 1 10 9 9 2
14 0 9 2 10 9 13 14 13 9 1 10 9 1 9
22 13 0 7 15 0 9 14 14 13 14 13 7 13 10 9 7 10 0 9 10 9 2
30 0 2 7 14 3 0 2 10 0 9 14 13 9 15 13 0 9 1 9 10 9 1 14 13 10 9 1 10 9 2
23 3 2 14 14 13 9 14 13 15 7 10 9 9 15 13 3 14 13 0 9 1 9 2
55 1 10 9 15 14 13 3 10 9 10 9 2 3 1 9 10 9 10 9 10 9 1 0 10 9 10 9 7 10 9 10 0 9 2 7 13 3 10 9 7 10 9 1 9 2 10 9 2 10 9 7 10 0 9 2
33 3 7 12 9 13 0 10 3 0 9 15 13 15 10 12 0 1 15 2 13 10 9 10 9 14 13 9 7 14 13 9 9 2
29 7 10 9 9 14 13 10 9 2 10 0 15 13 14 13 13 7 0 10 9 15 1 9 9 14 13 15 9 2
69 10 9 15 10 0 9 13 3 0 2 7 13 2 1 9 2 1 9 1 10 9 10 9 10 9 7 10 0 9 1 10 9 9 1 9 2 7 1 9 1 10 9 1 9 1 10 9 10 9 2 10 9 7 10 9 2 7 13 7 13 10 9 15 10 9 1 9 15 2
20 1 10 9 10 9 3 10 9 13 7 13 3 1 10 0 9 15 13 13 2
18 13 7 7 10 15 9 9 14 13 3 10 9 10 9 1 0 9 2
8 12 9 10 9 9 1 0 9
1 9
35 1 9 15 1 0 9 2 10 9 9 13 7 10 9 13 0 9 2 1 10 9 7 10 0 10 9 13 13 14 13 10 0 10 0 2
4 2 2 1 2
74 10 0 9 9 13 10 12 1 9 7 10 0 1 9 7 10 9 2 10 15 13 10 0 9 9 2 9 10 9 15 13 1 10 0 9 2 3 10 9 13 10 12 2 7 15 0 9 9 7 9 3 10 9 2 10 9 2 10 0 9 7 7 10 9 10 9 2 10 9 12 2 10 9 2
16 0 7 10 9 10 9 2 14 13 14 15 13 0 1 9 2
33 10 0 9 10 9 15 13 10 9 10 9 1 10 9 9 13 13 7 2 14 13 10 9 1 10 0 0 9 1 10 9 9 2
10 13 3 0 7 10 9 13 0 9 2
17 1 10 0 9 13 10 9 9 10 0 9 2 15 7 13 3 2
38 1 10 9 10 0 9 1 9 2 10 0 9 2 1 14 13 10 9 15 2 13 1 9 7 13 9 10 9 2 1 10 9 7 10 9 13 9 2
20 1 12 9 2 10 9 13 0 7 13 14 13 1 9 10 9 1 12 9 2
34 3 13 2 2 10 9 13 1 9 9 2 7 10 0 13 9 13 1 9 7 13 0 9 1 9 9 3 1 9 10 9 9 2 2
15 1 0 9 2 13 12 1 15 10 9 1 0 15 9 2
19 10 9 10 9 14 13 10 9 1 9 1 10 0 9 13 0 9 2 2
17 10 9 13 9 9 7 10 9 15 1 10 9 13 12 0 9 2
10 13 0 9 14 13 9 1 9 15 2
15 10 9 1 10 0 9 13 0 7 10 9 13 13 0 2
33 7 2 10 9 9 13 7 2 7 3 13 1 9 2 2 3 1 10 9 10 15 9 2 10 0 9 9 10 9 13 9 2 2
18 3 2 7 2 13 0 7 0 10 9 15 1 10 9 9 7 9 2
10 3 2 10 12 9 14 13 1 9 2
1 9
20 3 10 12 13 1 9 10 9 2 10 15 3 13 9 15 13 13 0 9 2
37 3 3 10 9 10 9 1 10 9 9 2 10 9 0 9 10 9 9 13 10 0 9 10 9 10 0 0 9 15 13 3 15 10 12 0 9 2
31 7 10 12 9 9 13 7 2 10 0 9 14 13 14 13 7 14 13 0 9 7 13 10 0 9 15 1 0 9 2 2
14 3 2 10 9 9 15 14 13 10 9 1 13 9 2
18 3 2 1 9 10 9 10 2 9 13 14 13 10 9 7 10 9 2
21 15 13 10 0 9 3 1 10 9 10 12 9 9 10 0 15 9 1 10 9 2
22 10 9 13 1 9 10 9 0 9 9 2 10 15 13 3 9 1 10 9 10 9 2
46 12 0 9 13 1 10 9 10 9 10 9 2 10 0 0 9 2 2 2 2 15 13 1 12 9 0 0 9 7 10 0 9 0 9 2 2 2 1 9 1 9 9 10 0 9 2
5 1 15 9 13 2
15 7 2 10 9 10 9 10 9 13 9 9 3 9 9 2
24 1 0 9 2 10 9 13 0 0 9 1 10 9 9 2 10 15 13 10 9 1 10 9 2
24 10 9 13 7 13 1 9 10 2 2 13 3 10 0 0 9 2 2 13 7 3 10 9 2
32 10 9 12 13 0 9 9 2 7 13 15 9 14 13 1 9 7 14 13 1 0 9 2 7 13 9 1 9 7 1 9 2
26 13 3 10 2 1 9 10 9 9 15 13 9 9 10 0 0 9 2 10 0 2 3 7 15 9 2
15 13 10 9 3 1 10 9 9 9 2 13 10 0 9 2
11 10 9 15 13 1 10 14 13 9 9 2
14 2 10 9 13 14 13 3 1 9 7 13 1 9 2
27 1 9 15 2 10 9 13 7 13 0 9 1 9 10 0 9 1 10 9 10 9 10 9 10 0 9 2
11 3 15 13 0 0 9 1 10 0 9 2
27 3 9 1 10 9 13 3 1 2 1 9 9 7 2 1 12 9 1 3 14 14 13 13 7 9 2 2
6 13 3 13 0 9 2
15 0 9 2 10 9 2 10 3 0 9 13 1 0 9 2
6 10 9 13 14 13 2
34 13 3 0 7 13 14 13 10 0 9 1 10 9 15 13 14 13 2 3 10 9 9 2 1 15 15 13 14 13 2 3 10 9 2
12 10 9 13 9 7 3 1 9 7 1 9 2
14 13 14 13 1 0 9 10 0 9 1 0 9 15 2
48 10 0 9 10 9 2 3 15 13 3 2 3 13 3 10 0 9 10 9 2 3 10 9 7 9 1 0 10 9 0 9 9 7 9 1 10 9 15 14 13 1 9 7 10 9 10 9 2
23 10 9 15 13 0 7 13 3 1 10 9 2 10 9 15 7 10 9 10 9 15 2 2
14 10 9 13 14 13 7 14 13 3 1 10 0 9 2
1 9
31 1 9 2 10 9 10 0 9 13 14 13 0 9 2 9 9 2 9 9 2 9 2 9 2 3 7 14 13 9 9 2
31 10 2 13 14 13 10 9 1 9 10 9 10 9 10 9 9 2 7 14 1 9 10 9 14 13 7 14 9 1 9 2
17 10 9 1 9 13 3 2 3 13 10 2 9 2 0 7 0 2
55 13 10 0 9 9 1 10 9 1 10 9 10 9 7 13 14 13 15 10 9 2 15 13 3 0 1 10 0 9 2 7 2 1 14 13 10 9 15 13 3 2 14 14 13 15 10 9 2 3 13 13 3 0 9 2
21 0 2 9 7 9 13 13 2 7 1 9 13 10 0 9 0 9 7 0 9 2
56 10 9 9 13 7 2 10 9 10 9 10 9 2 3 10 9 15 1 0 2 0 7 10 9 15 1 9 9 7 9 7 1 0 9 1 9 7 10 9 2 13 14 3 0 0 9 2 7 7 10 0 9 10 9 2 2
33 7 2 15 14 13 14 13 1 14 13 10 9 10 9 7 3 10 0 0 9 15 14 13 1 14 13 10 9 10 0 0 9 2
19 10 9 0 9 1 10 9 10 9 10 0 9 13 10 9 9 9 9 2
28 10 0 9 10 9 13 10 9 10 9 7 13 7 10 9 13 13 3 3 1 9 10 9 15 1 0 9 2
35 14 14 13 7 10 9 7 10 9 10 0 0 9 9 1 10 9 9 1 9 10 9 14 13 3 0 1 10 0 9 1 10 9 9 2
24 15 13 2 13 2 10 9 1 10 15 13 13 1 9 10 9 12 3 1 10 9 1 9 2
18 10 9 9 13 10 12 10 9 2 12 0 9 0 1 10 9 9 2
17 10 0 9 2 3 12 2 2 14 13 14 15 13 1 10 9 2
55 2 3 14 13 0 14 14 13 15 2 3 14 13 15 9 9 2 15 14 13 3 0 2 2 7 2 3 13 3 2 7 10 9 13 9 1 9 2 13 14 13 15 9 1 0 9 7 14 13 0 9 1 15 9 2
22 13 3 9 10 9 13 10 9 14 13 9 1 10 0 0 0 9 2 9 2 9 2
16 13 3 14 13 10 9 15 13 10 9 10 0 7 10 2 2
13 1 9 10 13 0 9 13 10 9 1 0 9 2
20 10 9 13 2 3 2 10 0 9 14 13 3 9 7 14 13 10 0 9 2
16 9 10 9 13 10 9 12 9 2 3 7 10 9 12 9 2
36 10 9 2 12 13 10 0 2 0 0 9 15 13 1 14 13 0 9 2 3 0 9 2 9 7 9 2 9 2 3 7 9 9 7 9 2
15 7 13 9 1 12 15 9 2 14 13 3 13 3 0 2
24 3 2 10 9 13 13 10 0 9 1 10 9 10 9 7 14 13 0 10 9 10 0 9 2
13 3 2 10 9 9 1 10 0 9 13 3 9 2
49 10 12 9 15 13 10 3 2 14 13 10 9 15 10 9 2 1 9 1 10 9 10 9 15 2 14 13 1 9 9 1 9 9 1 0 0 9 7 14 13 0 9 10 15 13 3 14 13 2
28 10 9 13 0 9 10 0 9 15 2 10 15 13 3 1 9 2 7 10 0 9 10 0 9 13 1 2 2
12 13 1 10 9 0 9 2 7 13 1 9 2
43 10 9 14 13 2 3 2 10 9 10 9 7 14 13 10 9 15 1 10 9 10 9 2 7 14 13 2 14 13 10 9 9 10 9 15 3 1 10 9 10 0 9 2
24 10 9 9 2 12 2 2 2 9 2 12 2 2 7 9 2 12 2 2 13 0 1 9 2
19 13 0 1 10 9 9 7 9 1 10 9 10 9 2 1 10 0 9 2
12 3 9 2 10 0 9 14 13 1 10 9 2
16 10 9 9 13 10 9 13 10 9 9 1 9 10 9 9 2
27 3 13 10 9 1 10 2 2 14 13 14 13 7 2 1 9 10 0 9 2 10 9 14 13 3 0 2
20 13 7 14 15 13 3 10 9 7 10 9 10 9 15 1 15 13 1 3 2
23 2 0 3 13 0 7 15 14 13 15 13 14 13 2 2 13 10 9 2 9 10 9 2
15 1 9 10 9 15 2 1 9 2 13 10 9 10 9 2
1 9
37 1 9 10 2 2 10 9 9 9 15 13 1 10 9 13 1 10 0 9 2 7 14 13 3 9 1 10 9 15 9 15 3 13 10 0 9 2
57 10 9 2 9 9 2 13 1 10 9 0 9 9 9 2 13 10 9 7 13 12 0 9 10 9 1 9 9 1 10 9 10 9 9 12 2 2 15 13 7 10 9 9 7 1 9 9 1 9 9 2 9 1 9 9 12 2
20 10 9 13 10 0 9 1 0 9 10 9 9 13 1 10 0 2 0 9 2
17 13 7 10 9 7 13 0 10 9 10 9 15 13 10 9 9 2
37 13 3 0 9 1 0 9 10 9 2 1 9 10 12 3 13 9 1 10 3 9 9 9 2 10 15 15 13 1 9 1 10 0 9 15 13 2
14 14 13 1 12 9 2 10 9 10 15 13 9 9 2
17 10 9 13 10 9 14 1 15 7 1 9 10 9 9 10 9 2
10 13 1 10 0 9 10 9 9 9 2
19 14 13 14 13 9 1 9 2 7 15 13 1 9 10 0 9 1 0 2
45 10 9 15 13 10 9 15 2 3 10 9 0 9 3 1 10 9 9 2 7 3 14 13 3 3 1 10 9 9 2 7 3 1 10 9 9 2 13 9 1 9 1 10 9 2
55 3 2 10 9 10 9 10 9 1 10 9 1 0 10 0 0 9 7 9 1 9 10 9 13 10 3 0 0 9 2 10 15 14 13 14 13 1 9 10 9 9 7 9 2 7 1 9 10 0 9 10 9 1 9 2
22 10 9 9 1 9 13 13 0 9 1 2 1 10 9 0 9 7 10 9 1 9 2
13 13 7 10 9 9 13 9 0 9 1 9 15 2
31 1 9 13 1 9 10 0 9 1 10 9 2 1 10 9 9 10 12 0 9 10 0 9 2 9 2 9 2 9 2 2
15 0 9 13 7 1 0 9 2 10 15 13 13 1 9 2
26 10 9 10 9 13 14 13 3 1 10 0 15 9 14 13 7 14 13 3 9 10 15 14 13 13 2
72 3 2 13 14 13 14 13 3 10 0 9 1 0 9 10 9 15 1 10 0 9 15 13 1 10 9 2 3 10 9 2 10 9 2 10 9 7 10 0 9 2 9 15 2 3 13 15 1 15 1 9 15 2 13 7 1 10 0 15 9 2 1 15 1 9 15 13 1 10 0 9 2
87 13 0 9 10 9 7 13 2 3 1 10 9 9 7 1 9 1 10 9 10 0 9 2 7 2 10 9 14 13 0 2 7 0 2 7 10 9 10 9 13 7 9 10 9 2 2 7 7 2 10 9 14 13 0 15 14 13 10 9 10 9 7 14 15 13 1 0 9 7 0 9 1 10 0 9 7 10 15 9 2 9 10 9 10 9 2 2
51 13 2 3 2 7 10 9 15 2 15 13 14 13 1 10 9 2 13 10 12 9 1 9 1 15 13 0 10 9 9 2 1 9 1 10 9 9 15 13 10 9 2 10 9 7 10 9 9 10 9 2
17 10 9 10 9 13 13 1 9 10 9 3 1 10 9 10 9 2
52 3 10 0 15 13 13 14 13 10 9 15 1 10 12 9 2 3 2 7 13 14 13 10 0 15 9 14 15 13 7 3 2 7 10 0 9 14 13 1 9 10 9 15 13 3 1 10 9 9 7 9 2
31 13 10 9 10 9 3 10 9 14 13 10 9 1 0 9 1 10 9 15 14 13 9 1 10 9 3 1 10 0 9 2
9 13 9 1 10 9 10 0 9 2
36 10 12 0 14 13 1 12 9 1 9 2 9 9 2 2 1 10 9 14 13 9 7 9 7 1 10 0 9 14 13 9 1 9 12 9 2
29 1 9 10 9 2 13 10 9 9 3 1 10 9 15 3 7 1 10 9 15 14 13 9 7 14 13 0 9 2
11 10 0 9 15 14 13 14 13 10 9 2
23 1 10 9 3 13 10 9 10 9 2 1 10 9 10 0 0 9 2 13 1 9 15 2
39 0 1 12 9 9 13 1 9 3 1 10 9 10 9 2 3 1 9 1 10 9 3 13 10 2 9 10 9 2 2 3 1 12 9 3 2 1 3 2
6 7 12 1 10 12 2
12 10 9 10 12 9 9 13 1 10 0 9 2
19 13 0 3 9 2 0 9 9 1 10 9 9 2 10 15 13 14 13 2
17 10 9 13 7 7 10 9 13 15 9 10 9 15 13 9 9 2
31 12 1 10 9 10 9 2 10 9 9 2 13 7 10 9 15 13 1 10 9 10 0 9 1 9 13 10 9 10 9 2
16 9 2 10 0 9 14 13 1 9 10 9 1 10 9 9 2
8 10 9 13 1 9 0 9 2
33 13 9 1 0 15 2 10 9 2 10 9 7 10 9 2 14 13 15 10 0 2 7 13 0 14 13 14 13 7 14 15 13 2
39 1 9 15 2 10 9 13 2 1 15 2 7 3 14 13 13 9 1 9 10 9 1 9 10 9 2 7 7 10 9 13 13 10 9 9 15 10 9 2
15 10 9 10 9 9 1 9 14 13 10 9 1 10 2 2
23 3 1 10 9 9 2 9 1 9 10 9 13 0 9 1 10 9 10 0 9 10 9 2
33 1 10 9 15 15 10 0 9 13 10 9 9 15 13 1 10 9 14 13 10 9 2 13 7 13 9 1 10 9 1 2 9 2
10 15 13 7 13 9 9 3 7 9 2
59 1 3 2 10 0 9 9 10 9 13 10 9 7 2 10 0 0 9 10 9 13 0 9 1 9 9 10 9 15 13 1 9 2 3 7 14 13 14 13 1 9 1 14 13 1 0 9 15 13 10 9 9 9 1 9 10 9 2 2
3 2 9 2
37 9 10 9 7 9 13 7 2 0 9 1 0 9 7 0 10 9 9 1 9 10 9 13 3 9 14 13 10 9 15 12 9 7 12 0 2 2
23 10 9 9 13 13 3 12 9 2 0 9 2 2 1 14 13 9 15 13 10 9 15 2
3 2 9 2
23 1 10 0 15 9 13 3 7 10 9 1 9 7 9 13 0 15 10 9 9 0 9 2
32 13 7 15 10 9 14 13 3 1 9 1 9 7 1 10 15 15 9 9 10 2 2 7 10 9 13 10 9 15 1 9 2
18 3 2 10 9 13 10 9 0 9 1 9 12 7 13 1 0 9 2
30 10 9 13 1 10 2 2 12 9 2 2 2 9 9 2 2 2 9 9 2 2 2 9 2 7 2 9 9 2 2
30 13 10 0 9 10 2 7 14 13 10 0 0 9 7 14 13 15 0 0 0 9 2 10 15 13 3 0 7 0 2
44 1 12 9 2 13 1 10 12 9 9 2 10 0 1 9 9 7 10 9 10 0 0 9 2 3 1 9 10 0 9 10 9 13 12 9 2 12 9 7 0 1 12 9 2
9 3 2 12 9 1 9 13 3 2
26 7 13 9 1 10 9 2 10 0 14 13 3 1 15 7 7 13 0 9 2 3 2 14 15 13 2
13 13 1 0 9 1 9 10 9 1 10 9 15 2
47 10 12 0 0 0 9 13 0 10 0 9 9 12 9 1 10 0 9 15 13 12 1 15 1 9 15 13 1 9 1 0 15 9 7 10 9 13 1 10 9 7 13 3 14 13 15 2
21 10 12 15 13 1 9 13 7 3 15 10 9 10 9 15 13 9 1 9 2 2
11 10 9 9 13 1 10 9 9 1 9 12
29 3 13 3 0 10 0 9 1 10 9 15 10 9 1 10 9 7 15 10 9 14 13 1 9 10 9 10 9 2
20 15 14 13 10 12 9 10 9 2 10 15 13 15 9 1 9 7 10 12 2
22 1 10 0 9 10 9 13 10 9 10 0 15 9 2 3 15 13 3 15 10 9 2
14 10 9 9 10 2 7 10 9 10 9 13 1 15 2
14 1 0 9 15 2 10 9 9 10 9 13 3 0 2
9 13 7 13 9 1 15 15 9 2
19 12 9 13 7 1 10 12 9 7 1 15 10 9 10 0 13 14 13 2
16 13 3 10 9 10 9 2 9 2 7 3 10 9 10 9 2
26 10 9 10 9 13 10 9 10 9 1 0 9 10 9 10 0 9 2 10 15 13 1 12 0 9 2
30 10 9 13 10 0 9 1 10 9 10 9 9 10 9 7 13 3 3 0 10 9 15 13 1 10 9 3 10 9 2
34 14 13 10 9 0 10 0 9 2 10 9 10 9 10 9 2 10 9 2 10 9 9 10 9 10 9 2 10 9 0 9 7 9 2
18 1 0 9 10 9 10 9 13 9 1 14 13 10 9 0 0 9 2
14 1 9 1 10 0 9 15 13 2 13 14 13 9 2
29 13 14 13 10 9 0 9 2 15 13 3 13 2 1 15 2 10 9 2 9 15 14 13 14 13 1 0 9 2
24 10 0 10 9 13 1 12 0 9 15 3 13 3 14 13 15 10 9 1 14 13 0 9 2
41 1 10 3 9 10 9 13 7 14 13 14 13 13 3 10 9 14 13 10 9 9 10 9 3 1 10 9 0 9 3 13 10 9 7 10 9 15 13 1 9 2
39 1 0 0 9 13 9 9 1 9 7 10 9 10 9 10 9 1 9 13 9 9 1 9 10 9 15 13 1 0 9 14 13 3 0 9 1 10 9 2
49 10 9 9 10 9 2 9 9 9 9 2 13 7 2 12 9 1 10 9 13 1 9 2 7 13 7 2 10 9 13 14 13 1 7 12 9 2 10 15 14 13 3 1 3 13 10 9 2 2
17 10 9 13 10 9 15 1 12 1 10 9 15 2 10 9 9 2
12 9 9 2 10 9 13 14 13 1 0 9 2
10 13 10 9 9 10 15 1 15 13 2
40 3 3 13 7 0 7 0 9 2 3 7 9 10 9 2 9 9 7 9 9 2 2 1 10 15 13 14 13 3 3 10 9 1 0 9 9 1 12 9 2
23 3 2 3 13 10 0 9 13 1 0 9 10 0 9 2 10 0 9 7 10 9 9 2
23 9 9 13 10 9 2 7 1 9 12 9 13 13 10 9 15 7 12 13 13 1 9 2
11 1 10 9 13 0 9 1 10 0 9 2
52 13 7 7 2 3 1 12 9 9 3 1 10 9 9 9 1 10 0 9 9 2 13 13 1 9 2 7 0 14 13 14 13 1 9 9 2 1 10 15 14 13 14 13 7 14 13 10 9 1 0 9 2
12 9 15 13 10 9 1 9 10 9 10 9 2
24 7 3 2 1 9 15 2 14 13 10 0 9 9 7 10 14 0 9 1 9 10 0 9 2
23 10 0 9 9 10 2 2 9 9 2 13 1 12 9 3 1 9 7 0 9 0 9 2
27 3 3 10 0 9 2 3 7 15 15 2 13 14 13 2 13 3 0 9 7 14 13 10 9 15 3 2
19 7 10 9 13 3 9 2 14 14 13 14 15 13 3 1 15 10 9 2
42 10 9 13 12 1 10 3 0 9 10 0 9 7 13 10 0 2 0 0 1 9 2 2 0 9 10 12 9 2 10 9 2 10 9 7 10 0 9 10 0 9 2
25 14 13 9 1 14 13 7 13 14 13 10 0 9 3 7 3 1 14 13 10 13 7 13 9 2
33 13 14 15 13 15 2 7 3 13 10 9 15 1 10 9 2 7 1 15 10 9 2 9 7 9 2 10 12 9 15 15 13 2
8 13 7 10 15 9 10 9 2
17 9 9 2 14 13 14 13 1 9 10 9 10 9 1 0 9 2
29 14 13 9 10 9 3 7 7 10 9 15 13 1 9 15 13 3 0 3 13 10 9 15 13 1 15 10 9 2
28 3 2 13 10 9 14 13 7 0 9 1 0 9 2 7 14 13 0 9 1 9 7 9 15 13 3 9 2
6 13 10 9 0 1 9
27 3 2 10 9 13 10 9 1 14 13 0 9 2 7 14 13 10 9 10 9 1 0 9 1 0 9 2
40 10 0 9 14 13 1 10 9 10 9 2 10 9 10 0 9 2 10 15 13 1 9 15 10 9 9 2 7 10 15 13 1 9 10 0 9 10 12 9 2
11 10 9 13 9 12 0 7 0 9 9 2
13 9 10 9 13 9 7 14 13 14 13 0 3 2
45 10 0 9 15 13 7 2 10 0 9 13 14 13 10 9 10 0 9 9 2 10 15 14 13 7 14 13 10 9 9 7 9 15 13 1 10 9 2 10 9 7 10 9 2 2
37 1 9 10 0 9 7 13 3 10 9 10 9 1 10 0 0 9 2 13 7 0 9 10 0 9 14 13 14 13 10 9 10 9 10 9 9 2
28 10 15 2 3 1 10 0 9 9 7 10 9 9 1 10 9 9 7 10 15 3 1 10 0 9 10 9 2
31 10 9 15 13 1 10 9 10 0 9 14 13 10 0 9 10 9 7 10 9 7 14 13 10 9 1 3 3 0 9 2
31 7 10 9 10 9 10 9 1 0 9 13 1 9 9 1 10 9 2 10 0 9 10 15 14 13 1 9 10 0 9 2
32 1 10 9 10 9 3 0 9 2 10 9 13 0 7 1 10 9 2 14 13 10 9 1 0 9 9 3 13 2 10 9 2
25 15 13 3 1 9 10 0 9 2 3 10 0 2 10 0 7 10 9 15 13 10 9 1 9 2
54 3 2 1 0 9 15 13 10 2 7 10 9 10 12 2 1 14 13 10 9 10 9 1 10 15 9 1 15 2 14 13 3 14 13 13 9 9 1 10 9 15 7 14 13 0 9 15 14 15 13 1 0 9 2
12 7 10 9 13 10 9 2 10 0 9 13 2
16 1 9 2 1 10 0 9 10 9 13 9 7 13 10 9 2
57 1 10 9 3 14 13 13 2 10 9 14 13 10 0 9 1 9 10 9 7 10 9 10 9 2 10 9 10 15 13 1 0 9 7 1 9 1 15 10 0 9 15 14 13 10 9 7 14 13 10 9 15 1 3 0 9 2
39 10 9 9 10 9 2 9 9 2 13 10 9 9 15 14 13 1 2 7 15 9 10 2 14 13 9 1 0 9 3 9 9 10 9 15 13 1 9 2
54 1 9 2 14 13 3 0 15 15 13 10 9 1 9 1 10 0 9 7 10 9 2 3 2 1 15 2 3 1 10 9 15 13 1 0 9 2 13 7 1 10 0 10 9 2 3 1 14 13 10 9 10 9 2
23 7 2 7 10 9 15 13 1 10 0 12 9 2 3 14 13 3 3 1 10 9 15 2
12 3 14 13 10 9 10 9 1 10 0 15 2
32 10 0 9 1 10 0 9 10 0 9 0 0 7 0 9 3 9 13 14 13 10 0 9 7 14 13 10 9 10 0 9 2
36 7 7 10 9 9 9 1 9 2 12 13 13 1 0 10 0 9 1 10 9 2 13 7 10 9 15 13 10 9 13 3 1 15 10 9 2
12 3 1 10 9 13 7 10 9 15 2 9 2
16 10 12 9 13 10 9 10 9 1 9 1 10 9 10 9 2
4 10 9 9 2
41 9 7 9 2 14 13 10 9 3 10 9 1 9 7 3 13 14 13 7 10 2 9 2 1 2 9 9 2 10 9 2 13 7 15 13 1 10 9 10 0 2
1 9
31 3 10 9 9 13 1 9 9 10 9 15 13 7 14 13 14 13 1 9 2 1 3 13 14 13 1 9 1 0 9 2
38 10 9 13 0 9 3 13 10 0 9 7 10 9 2 15 13 10 9 0 10 0 9 10 2 7 13 10 12 10 9 9 7 10 12 10 9 9 2
14 10 9 10 12 9 13 1 0 9 15 13 10 9 2
11 10 9 10 9 13 1 9 10 0 9 2
25 3 2 10 12 0 9 15 13 14 13 13 7 10 9 13 10 9 10 0 9 1 10 9 9 2
30 3 1 10 9 2 10 9 10 0 9 7 10 9 10 9 13 10 0 9 10 9 15 13 10 9 10 9 1 9 2
23 1 9 10 0 0 9 2 10 0 9 10 0 13 13 10 9 0 7 0 9 7 9 2
29 10 9 14 13 14 13 10 9 10 9 15 2 14 13 14 13 7 7 14 13 0 1 9 14 13 13 15 0 2
31 10 9 15 13 7 10 0 9 13 0 2 7 1 10 9 15 13 1 0 9 10 0 9 10 9 3 1 15 10 9 2
29 13 3 0 2 14 13 1 9 15 1 15 9 2 14 13 14 13 3 9 12 9 10 15 13 0 1 0 9 2
