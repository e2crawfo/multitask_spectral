1115 11
6 16 15 13 2 13 2
5 9 14 15 13 2
7 1 9 15 13 14 13 2
5 0 9 3 13 2
10 1 9 4 13 11 2 0 15 9 2
6 1 9 13 1 11 2
7 3 13 9 1 15 14 2
9 13 0 9 3 7 3 1 9 2
9 12 9 13 14 15 13 3 3 2
5 14 15 13 3 2
7 1 9 13 1 9 12 2
12 1 0 9 15 13 0 7 0 9 1 9 2
7 3 1 0 9 4 13 2
13 7 15 2 0 2 6 13 2 16 15 4 13 2
7 0 1 9 13 9 15 2
8 7 13 3 0 9 1 9 2
9 9 11 4 13 1 9 1 11 2
7 9 15 14 13 1 11 2
10 9 11 15 13 1 9 2 9 13 2
7 15 0 9 15 13 3 2
5 9 13 1 0 2
15 0 9 15 15 13 1 0 15 9 2 7 13 9 15 2
13 9 14 13 2 0 14 13 2 7 13 3 0 2
8 9 1 11 13 14 13 0 2
6 13 14 6 15 13 2
8 6 13 14 4 13 1 15 2
17 9 15 13 1 0 9 7 3 1 15 13 14 13 9 1 9 2
7 1 14 15 13 2 13 2
11 15 15 13 0 2 3 4 13 9 3 2
11 1 3 16 13 0 2 14 13 1 9 2
11 16 13 14 13 9 2 13 14 13 9 2
15 14 13 0 2 13 14 13 1 9 14 15 13 10 9 2
10 13 15 2 14 6 13 14 15 13 2
10 15 13 3 2 16 13 14 13 9 2
9 16 9 13 9 2 14 15 13 2
9 13 3 1 9 2 16 13 0 2
14 1 14 13 3 1 9 15 2 14 13 1 10 9 2
10 14 3 14 13 9 2 15 13 9 2
14 3 0 9 2 15 13 3 2 15 13 14 15 13 2
13 0 13 2 16 15 4 13 3 1 9 1 9 2
9 0 9 13 2 16 9 15 13 2
7 0 9 15 13 3 3 2
10 1 10 9 7 9 3 15 13 9 2
16 9 13 0 2 1 15 15 13 2 7 3 14 13 6 13 2
11 13 15 15 13 2 16 3 14 15 13 2
6 6 13 14 13 9 2
15 12 9 13 4 14 13 7 16 16 13 0 9 1 9 2
6 11 13 0 7 0 2
7 9 11 15 13 1 0 2
5 9 13 1 9 2
8 10 9 13 3 1 0 9 2
9 13 0 0 9 2 0 7 0 2
5 11 13 0 9 2
7 15 6 13 2 15 13 2
6 13 15 1 0 9 2
11 7 6 13 15 2 9 2 1 0 9 2
16 7 1 9 2 3 4 13 1 0 9 7 9 2 9 13 2
7 1 9 13 14 15 13 2
20 3 1 10 9 15 13 9 15 2 16 10 0 9 13 14 13 1 10 9 2
12 16 13 2 16 9 13 3 2 11 15 13 2
5 15 15 15 13 2
8 7 3 15 13 9 1 9 2
7 1 0 0 9 13 9 2
11 3 3 6 13 10 9 7 10 0 9 2
12 1 9 13 3 12 2 9 15 13 1 9 2
16 1 9 15 13 10 9 3 2 7 9 13 1 9 1 9 2
10 9 2 9 2 9 4 13 1 9 2
14 13 2 16 3 2 1 10 9 2 13 9 1 11 2
11 9 6 15 13 2 7 15 13 9 15 2
12 9 13 14 15 13 1 0 0 9 1 9 2
15 7 16 9 13 14 15 13 2 15 15 13 1 9 15 2
12 13 15 2 1 14 13 11 14 15 13 9 2
8 7 14 13 9 1 10 9 2
3 15 13 2
6 6 13 3 15 13 2
9 13 15 15 14 15 4 3 13 2
7 14 15 13 15 14 13 2
6 0 10 9 13 0 2
5 14 15 13 15 2
8 13 14 13 14 13 1 15 2
5 13 3 14 13 2
9 3 14 13 2 15 13 1 15 2
5 1 9 15 13 2
6 13 14 11 9 15 2
9 9 4 13 2 1 14 4 13 2
5 10 0 9 13 2
9 10 1 10 9 13 1 12 9 2
8 3 13 9 1 9 1 9 2
11 3 13 3 3 9 2 16 15 15 13 2
6 15 4 13 1 15 2
8 9 13 9 1 15 1 15 2
4 2 13 15 2
14 13 14 13 14 15 13 14 15 13 14 13 14 13 2
6 15 15 13 1 0 2
9 3 13 2 16 15 6 13 3 2
6 9 13 14 15 13 2
6 15 13 14 15 13 2
6 13 2 16 4 13 2
5 13 15 14 13 2
6 13 15 14 13 3 2
6 13 15 14 13 15 2
5 13 2 15 13 2
11 9 1 10 2 16 4 13 2 13 0 2
12 10 9 15 15 13 2 10 9 15 15 13 2
10 15 13 9 2 1 15 14 15 13 2
8 13 9 2 3 14 13 9 2
10 3 13 1 15 2 3 14 15 13 2
7 14 15 13 2 16 13 2
7 14 13 2 13 14 13 2
7 14 13 2 3 15 13 2
8 13 15 2 1 14 6 13 2
5 13 14 13 9 2
9 15 13 9 2 3 15 13 9 2
3 11 13 2
5 13 15 14 13 2
6 14 3 15 13 9 2
7 13 15 2 16 14 13 2
8 9 2 0 1 9 2 13 2
8 6 2 9 1 9 4 13 2
8 6 13 3 1 15 14 13 2
9 13 1 9 2 1 14 13 15 2
6 2 15 13 0 13 2
9 15 13 2 16 9 14 13 0 2
13 1 3 15 13 9 2 3 15 6 15 15 13 2
7 15 15 15 15 4 13 2
5 15 15 15 13 2
5 13 15 16 13 2
6 13 0 2 0 9 2
13 13 4 9 1 9 15 1 11 2 11 2 11 2
21 0 13 9 1 0 9 1 9 1 10 9 1 10 9 1 3 0 9 1 11 2
26 9 13 2 16 9 2 1 15 13 0 9 2 13 0 9 2 3 15 4 13 1 9 1 0 9 2
32 9 1 9 1 0 11 2 0 1 9 1 9 1 9 1 11 1 0 9 1 11 2 3 13 0 9 1 9 1 10 9 2
12 6 13 3 3 14 15 13 10 9 1 11 2
24 2 1 10 0 2 0 9 11 13 3 3 0 9 1 3 11 1 9 2 11 2 14 11 2
20 15 6 13 2 7 9 15 13 1 0 9 2 7 10 9 13 1 15 0 2
17 3 15 13 2 16 1 15 4 13 0 9 1 0 9 1 9 2
10 1 10 6 3 0 9 15 13 3 2
26 0 1 9 13 9 2 15 0 9 6 4 15 13 1 9 1 11 2 3 9 6 13 9 1 15 2
13 10 13 0 9 1 11 14 13 1 9 1 11 2
9 13 2 9 15 13 0 1 15 2
11 14 3 11 15 13 7 1 10 0 9 2
13 13 14 9 1 10 9 15 13 0 9 0 9 2
8 9 15 9 15 4 3 13 2
39 16 15 13 3 9 1 9 1 9 1 12 0 9 1 9 2 15 13 1 3 0 9 1 0 9 2 1 0 7 0 9 1 0 15 9 7 0 9 2
14 9 1 9 1 0 9 13 0 1 9 1 12 9 2
21 9 1 0 9 13 0 9 7 9 2 0 7 0 1 0 7 0 9 1 9 2
35 16 16 14 6 13 14 3 3 9 1 9 2 15 13 0 9 7 16 16 14 9 1 9 15 13 3 1 9 1 9 1 9 1 9 2
11 13 15 7 15 13 1 10 15 13 9 2
20 13 15 9 2 9 7 1 3 1 0 9 13 0 7 0 9 1 0 9 2
22 2 14 13 0 7 3 3 0 1 0 15 9 2 0 1 9 7 9 1 9 15 2
8 3 7 9 14 13 14 13 2
16 9 2 15 3 13 9 2 13 0 9 1 0 9 1 11 2
15 10 9 7 0 15 9 3 15 13 1 0 9 7 9 2
11 2 6 2 13 0 9 14 13 10 9 2
43 0 0 9 15 13 1 0 9 1 9 7 1 0 9 1 3 0 9 1 9 1 9 2 9 7 9 1 9 2 0 9 2 1 15 9 7 9 1 0 9 13 0 2
14 3 15 13 1 0 15 2 1 15 15 4 13 3 2
18 13 4 3 9 2 13 15 9 7 13 14 15 13 1 9 3 3 2
11 15 13 1 3 0 15 0 9 1 9 2
14 15 15 13 1 3 0 9 1 9 7 1 0 9 2
8 13 7 3 3 6 15 13 2
8 9 3 15 13 1 9 15 2
16 7 9 13 7 15 13 1 9 3 7 9 13 1 1 9 2
20 3 2 9 9 2 3 3 3 13 14 4 13 2 1 14 13 10 10 9 2
29 13 2 16 9 1 10 9 14 15 13 1 9 1 0 9 13 0 7 15 13 9 1 9 1 9 1 10 9 2
18 11 13 14 13 9 1 10 9 2 3 15 14 13 7 9 1 9 2
9 13 4 9 1 9 1 0 9 2
21 1 9 4 13 7 9 1 9 7 9 1 9 1 0 9 1 9 1 0 9 2
18 0 13 7 9 1 0 0 9 1 0 0 9 1 9 1 0 9 2
33 1 9 1 0 13 0 9 2 1 15 13 9 1 0 1 7 1 9 0 9 0 9 7 0 9 1 9 1 9 7 0 9 2
4 10 9 13 2
7 15 13 14 13 9 15 2
7 3 14 15 13 1 9 2
4 15 6 13 2
7 14 4 14 13 10 9 2
7 3 13 0 9 1 9 2
7 9 15 13 1 3 9 2
9 2 13 0 9 1 9 1 9 2
8 13 1 9 7 3 3 9 2
10 0 9 2 13 15 2 13 1 3 2
8 9 1 0 9 13 9 11 2
8 15 13 1 9 1 0 9 2
10 3 2 7 9 11 15 13 3 9 2
9 7 1 10 9 9 13 1 9 2
3 9 13 2
5 0 9 15 13 2
10 2 13 9 7 9 1 9 1 9 2
10 11 13 3 3 9 13 1 9 15 2
11 2 10 9 14 13 3 7 14 13 9 2
10 1 10 9 13 0 1 0 9 9 2
10 9 15 13 1 0 9 1 0 9 2
6 13 15 3 7 3 2
11 15 13 1 10 0 0 9 1 0 9 2
11 3 13 9 1 9 1 0 9 1 9 2
13 3 13 14 1 9 14 15 13 2 3 15 13 2
5 15 13 0 9 2
12 13 14 10 0 9 14 13 9 1 0 9 2
13 9 15 13 3 9 7 13 9 3 1 0 9 2
14 2 13 9 1 9 1 9 1 9 7 9 1 9 2
13 15 13 3 9 7 13 1 9 7 1 0 9 2
13 3 13 9 1 9 1 9 1 0 9 1 9 2
15 9 3 13 9 7 16 13 14 13 9 15 2 13 9 2
4 7 1 15 2
13 12 9 13 1 0 9 14 15 13 7 12 9 2
17 7 15 13 1 9 15 3 1 14 15 13 14 13 3 10 9 2
14 14 15 13 14 13 14 13 7 14 15 13 1 9 2
15 9 13 1 0 9 1 9 9 1 0 9 1 0 9 2
19 7 15 2 9 2 15 13 1 9 15 2 13 15 9 7 15 13 3 2
10 15 13 11 14 13 7 13 3 9 2
42 15 13 14 13 3 14 4 13 9 2 0 1 9 1 9 1 0 9 2 3 16 15 13 9 3 1 9 1 10 3 0 9 1 11 2 7 15 13 0 15 9 2
16 7 15 15 13 2 13 15 7 15 13 2 16 15 6 13 2
25 1 9 1 0 2 0 1 0 9 9 2 9 2 9 9 3 13 14 13 9 1 9 1 9 2
7 11 13 14 6 15 13 2
21 9 13 9 1 0 15 9 7 14 1 3 15 13 2 14 6 15 15 13 15 2
16 7 6 13 14 13 10 0 9 2 3 6 15 13 3 3 2
15 13 15 3 14 13 3 1 15 2 1 14 13 9 15 2
25 3 3 13 14 15 13 2 16 3 3 10 9 4 13 7 1 0 0 9 1 0 9 1 9 2
9 15 6 13 14 9 1 0 9 2
19 13 0 2 0 2 1 0 9 2 7 11 13 14 15 15 13 3 3 2
6 6 13 14 13 9 2
20 9 9 2 13 14 9 14 13 0 9 1 9 1 9 7 9 1 0 9 2
8 13 15 3 1 0 15 9 2
6 0 14 13 0 9 2
28 12 9 7 12 9 13 9 2 9 13 2 9 13 7 0 9 2 0 7 1 3 2 13 1 9 7 9 2
6 2 3 15 15 13 2
16 9 1 0 9 13 9 1 9 1 9 7 9 1 0 9 2
17 10 0 9 14 13 9 1 9 1 0 7 0 9 1 0 9 2
18 0 9 15 13 7 1 9 1 9 1 0 9 7 9 1 0 9 2
18 1 0 9 4 13 0 9 1 9 1 0 9 7 9 1 10 9 2
20 14 15 13 9 1 9 1 9 1 0 9 1 0 7 0 9 1 0 9 2
20 1 9 1 10 9 10 9 2 3 1 0 9 2 4 13 0 9 1 9 2
17 1 9 1 0 9 13 1 9 7 0 9 1 0 9 1 9 2
13 10 9 3 6 13 2 7 13 14 13 1 9 2
7 9 4 13 2 9 13 2
5 10 15 13 3 2
9 7 3 15 13 14 13 0 9 2
6 15 3 6 15 13 2
31 7 3 15 1 0 9 2 0 13 2 16 3 4 13 9 2 0 9 6 4 13 10 9 1 9 2 1 15 15 13 2
6 15 13 10 9 9 2
17 9 1 9 1 0 9 1 11 7 0 11 2 13 9 1 11 2
11 3 13 9 1 9 2 1 14 13 3 2
9 9 15 13 1 0 9 1 9 2
19 0 2 15 13 14 15 13 13 14 9 13 14 15 13 1 9 1 11 2
19 13 15 2 1 14 15 13 10 0 9 1 9 1 0 9 7 10 9 2
8 7 15 13 0 9 1 9 2
8 7 10 9 13 3 12 9 2
22 3 3 4 13 0 9 1 0 9 1 9 1 0 9 1 11 7 1 0 0 9 2
5 13 15 3 9 2
22 7 15 13 2 16 1 9 1 0 9 3 14 13 3 9 2 1 14 15 13 3 2
5 14 14 13 0 2
10 9 1 0 9 14 15 13 1 9 2
13 1 0 9 2 3 13 2 9 6 13 1 11 2
10 16 15 13 2 14 15 13 3 2 2
13 16 15 13 9 2 13 15 7 15 13 1 9 2
4 15 15 13 2
11 15 3 13 0 9 2 3 15 13 3 2
14 3 7 14 13 0 9 3 2 15 13 14 4 13 2
27 10 2 1 15 3 3 13 0 9 1 9 1 9 1 0 0 9 2 7 13 1 9 1 9 1 9 2
6 0 9 13 1 9 2
22 10 9 2 10 9 2 15 13 1 15 7 13 1 9 1 9 15 13 10 0 9 2
22 15 13 1 0 9 2 3 9 7 9 3 13 14 13 9 2 6 3 1 0 9 2
11 9 1 9 1 0 9 13 2 13 15 2
16 1 12 9 1 9 7 9 13 2 16 13 9 6 15 13 2
33 3 13 2 13 7 16 15 13 2 16 13 1 9 15 2 13 15 2 13 15 9 9 2 7 15 13 7 13 3 3 1 3 2
13 9 15 13 1 0 2 0 7 0 9 1 9 2
18 15 6 13 6 15 13 3 2 9 9 2 3 13 15 6 13 9 2
9 0 9 1 15 3 13 0 9 2
7 1 9 1 0 9 14 2
21 15 6 15 13 2 7 13 9 15 14 13 3 1 9 1 0 9 1 0 9 2
10 4 13 1 9 2 16 6 13 9 2
13 10 10 9 1 0 9 15 15 13 0 7 0 2
16 9 2 13 2 13 1 9 2 13 15 2 7 6 15 13 2
4 15 13 9 2
11 15 13 9 2 13 4 14 13 3 9 2
10 9 13 14 13 3 7 1 3 9 2
8 9 2 13 2 13 1 9 2
8 3 15 2 9 13 0 9 2
5 3 9 15 13 2
3 7 12 2
8 6 15 13 2 7 3 13 2
13 13 15 7 15 13 1 9 15 2 3 4 13 2
14 13 15 1 9 1 9 15 2 15 13 14 15 13 2
5 2 13 15 2 2
6 2 13 2 13 15 2
5 7 9 1 15 2
26 4 13 9 1 9 15 2 4 15 13 14 15 13 2 6 15 4 13 1 9 7 9 15 15 13 2
6 2 3 15 13 11 2
3 1 15 2
3 2 7 15
7 9 13 14 15 13 0 2
12 11 2 15 13 9 1 9 2 13 0 9 2
8 9 15 13 3 10 0 9 2
13 6 4 13 2 16 14 13 3 2 7 15 13 2
34 6 16 4 15 15 13 2 3 14 13 14 13 1 15 2 7 13 1 9 1 9 2 1 9 2 15 3 7 3 13 14 15 13 2
38 9 15 13 2 6 15 13 14 15 13 1 9 2 3 1 0 9 7 15 15 13 1 9 2 13 13 6 3 7 6 3 14 15 13 1 15 14 2
5 14 2 14 13 2
13 2 15 13 9 1 9 7 10 9 13 10 9 2
10 13 0 15 0 9 2 13 9 15 2
3 1 9 2
13 2 1 14 13 3 12 9 2 15 13 9 15 2
7 15 14 13 1 9 15 2
8 9 13 0 0 9 1 11 2
12 15 13 3 3 0 9 2 9 13 3 9 2
15 3 13 0 9 2 13 15 10 2 15 4 13 1 15 2
39 1 10 9 2 0 1 9 1 9 1 9 2 9 1 0 9 2 9 2 9 1 9 7 9 1 9 15 2 15 13 9 1 9 2 0 1 0 9 2
1 9
9 1 15 6 15 13 0 0 9 2
19 15 13 1 9 12 9 1 9 15 2 1 3 1 15 4 13 0 9 2
20 9 1 9 7 9 1 0 9 2 3 7 9 1 10 9 15 13 1 9 2
5 0 9 13 0 2
17 9 13 0 0 9 2 15 15 13 1 0 9 1 9 7 9 2
6 0 9 7 9 1 9
10 9 1 0 9 15 13 1 0 9 2
18 6 15 13 1 9 0 9 7 9 1 9 1 9 1 9 7 9 2
26 9 2 1 15 0 9 6 13 0 2 13 9 3 1 0 9 1 0 9 14 13 7 13 10 9 2
14 9 1 9 7 9 1 9 7 9 15 13 1 9 2
21 9 7 9 1 9 1 9 15 13 9 7 9 1 10 9 7 15 13 1 9 2
2 0 9
20 9 7 9 1 0 9 15 13 1 9 1 11 7 1 9 2 0 1 15 2
19 9 13 0 7 3 2 1 3 11 13 7 0 9 13 15 14 13 3 2
11 0 9 1 0 9 15 13 1 12 9 2
10 9 15 13 1 9 7 1 0 9 2
12 0 9 15 13 1 9 2 9 9 7 9 2
10 1 9 0 9 13 7 9 7 9 2
15 0 0 9 15 13 1 12 0 9 2 0 1 0 9 2
9 9 2 9 2 9 2 9 2 9
10 7 9 1 9 1 0 9 13 0 2
13 3 3 13 9 1 9 2 0 9 7 0 9 2
11 11 13 14 13 14 15 13 9 1 9 2
20 9 14 13 1 10 0 9 1 0 9 2 1 15 13 13 6 1 0 9 2
17 3 15 13 14 15 13 1 10 0 9 1 9 1 0 0 9 2
22 7 9 1 10 0 1 0 9 9 1 11 11 11 15 13 1 2 9 1 9 2 2
23 6 13 3 10 9 14 13 1 10 9 1 9 2 1 15 4 13 0 9 1 10 9 2
6 7 10 9 1 9 2
19 15 13 9 1 9 2 15 13 0 9 7 13 14 13 9 1 10 9 2
10 9 13 3 7 13 9 1 0 9 2
14 3 3 0 15 14 13 14 15 13 1 9 7 9 2
5 3 15 15 13 2
12 13 15 12 7 12 9 2 15 13 3 0 2
5 15 13 0 9 2
16 16 15 13 2 13 15 9 7 13 9 2 9 14 13 3 2
3 13 11 2
23 16 13 3 9 1 0 9 1 9 2 13 14 15 13 14 12 9 2 1 15 13 9 2
4 13 7 13 2
5 0 13 1 9 2
5 13 9 7 9 2
14 6 13 3 0 9 2 1 14 13 15 1 12 9 2
9 13 9 2 16 15 13 1 15 2
11 9 13 14 15 13 2 16 13 3 0 2
7 7 15 13 9 1 9 2
3 13 9 2
20 2 3 9 13 9 2 15 3 15 13 3 1 9 2 1 15 13 14 13 2
10 1 15 15 13 1 9 1 10 9 2
13 9 1 11 11 2 2 11 2 2 9 0 9 2
14 0 9 13 3 1 10 0 0 9 2 15 3 13 2
2 15 2
7 1 10 9 14 13 0 2
12 7 9 13 1 9 1 9 7 15 13 9 2
26 1 0 9 15 13 9 9 7 12 0 9 2 15 14 15 13 1 0 9 2 0 9 7 0 9 2
5 3 14 13 10 9
5 15 13 0 9 2
11 13 0 9 2 3 7 9 1 0 9 2
5 15 13 0 9 2
14 0 3 4 13 1 9 1 9 7 9 1 0 9 2
28 10 12 9 1 9 4 13 1 9 1 12 9 2 11 2 7 11 2 0 2 11 2 7 11 2 0 2 2
32 0 9 1 9 13 9 1 9 1 0 9 1 9 2 3 4 13 1 9 2 9 7 9 2 11 2 7 11 2 0 2 2
12 9 1 0 9 13 0 1 0 7 0 9 2
35 13 15 1 9 2 9 2 9 2 0 0 9 2 9 1 9 1 0 2 9 2 9 2 0 9 2 0 9 7 9 1 9 1 9 2
11 2 13 15 1 9 2 9 7 9 2 2
8 2 3 6 13 1 9 2 2
9 2 3 15 13 1 9 15 2 2
13 0 9 1 10 9 13 2 16 15 13 3 0 2
7 9 1 9 7 9 1 9
24 1 10 9 9 13 9 1 9 2 15 13 1 9 1 0 9 1 0 1 9 1 0 9 2
11 15 13 1 9 1 9 15 1 0 9 2
22 10 9 4 13 1 9 1 0 9 2 11 11 11 2 2 11 7 0 2 0 2 2
16 10 9 3 6 13 3 0 7 13 14 15 13 1 9 15 2
33 3 13 2 16 9 1 9 1 9 14 13 0 9 1 9 1 0 9 1 9 1 10 2 15 4 13 0 0 9 2 16 13 2
15 1 0 9 14 13 3 1 9 2 1 15 10 9 13 2
9 2 13 13 1 9 1 12 9 2
11 11 11 2 12 9 2 2 9 2 11 2
19 10 9 4 13 0 9 7 1 11 3 1 0 9 2 7 3 12 9 2
5 13 9 1 0 9
10 11 3 6 13 10 9 2 13 1 11
21 1 9 15 13 0 9 1 9 7 9 7 15 13 9 1 12 9 2 13 15 2
11 3 15 13 0 9 2 3 3 13 9 2
11 9 1 9 4 15 13 7 1 0 9 2
16 15 13 9 11 11 1 9 1 2 9 12 2 1 0 9 2
13 13 9 1 9 1 9 1 9 2 13 1 11 2
11 0 13 0 9 1 9 7 9 1 0 9
7 9 13 3 1 0 9 2
17 9 13 14 15 13 9 7 1 9 1 11 1 0 9 1 11 2
8 1 15 1 0 9 1 9 2
6 9 13 12 9 9 9
17 9 1 0 0 9 13 0 9 1 0 0 9 2 13 0 9 2
28 1 9 1 15 11 14 15 13 1 9 1 0 9 1 9 2 13 9 2 11 11 11 2 2 0 1 11 2
19 0 9 2 11 2 1 9 12 14 4 13 1 0 0 9 1 0 9 2
17 1 0 9 1 0 9 14 15 13 9 1 0 0 9 11 11 2
8 0 13 1 0 9 1 9 2
8 0 9 13 1 3 0 9 2
5 9 13 12 0 9
18 10 0 9 1 9 1 2 11 11 2 13 1 9 2 0 9 2 2
17 9 15 13 1 10 2 16 1 9 9 1 9 15 13 9 12 2
8 0 9 13 14 13 7 9 2
13 0 13 1 9 1 2 9 2 11 11 7 11 2
17 9 13 14 6 15 13 9 15 1 0 2 0 1 15 0 9 2
12 1 10 9 15 13 11 2 9 7 9 11 2
18 3 9 1 11 13 9 1 9 1 0 9 2 10 9 6 4 13 2
25 9 1 9 1 2 11 2 11 11 4 13 1 9 1 9 1 11 2 13 0 9 11 11 3 2
7 0 15 13 3 1 9 2
11 11 11 2 12 9 2 2 9 2 11 2
5 2 6 2 13 2
13 13 14 6 13 3 9 2 1 14 6 13 3 2
22 13 10 2 0 9 1 9 2 2 15 13 9 7 9 1 9 1 9 1 0 9 2
18 2 0 2 7 2 9 2 13 0 12 9 1 9 1 9 1 9 2
10 2 0 9 13 11 2 2 11 2 2
18 2 9 13 14 13 9 6 3 1 0 9 2 7 7 1 0 9 2
21 6 15 13 2 16 9 15 13 1 9 2 3 15 13 7 3 13 0 15 9 2
22 0 1 9 9 14 4 13 1 9 1 9 1 11 2 3 16 15 14 15 13 14 13
19 1 15 13 9 2 9 2 1 14 15 13 0 9 7 14 13 0 9 2
37 15 13 2 16 9 4 13 14 4 13 10 9 7 4 13 3 1 9 15 2 13 0 9 1 9 11 11 2 15 3 13 9 1 2 11 2 2
13 15 13 14 13 9 3 1 9 2 7 0 9 2
11 1 0 9 0 9 4 13 9 12 9 2
10 9 13 14 13 7 9 12 9 9 2
13 15 13 2 16 9 1 9 10 9 14 4 13 2
8 1 0 9 13 1 9 1 9
5 0 11 3 15 13
10 9 15 13 1 0 9 1 12 9 2
11 13 0 2 3 16 9 13 1 0 9 2
21 12 9 3 13 0 9 1 10 9 1 9 1 0 9 2 13 0 9 11 11 2
17 1 15 9 3 13 2 9 2 15 14 6 15 13 1 0 9 2
12 7 15 13 1 0 9 2 0 3 1 11 2
21 10 9 1 10 7 14 13 9 1 0 9 1 9 13 1 9 1 3 0 9 2
10 2 13 2 16 13 0 9 1 9 2
14 1 9 13 7 9 1 0 9 7 9 1 0 9 2
11 11 11 2 12 9 2 2 9 2 11 2
11 11 11 2 12 9 2 2 9 2 11 2
13 1 9 15 4 4 13 1 9 1 9 1 9 2
15 13 15 0 9 2 9 7 9 2 9 1 9 1 11 2
24 1 9 1 9 4 13 7 9 2 0 9 2 0 9 1 9 7 1 10 9 1 11 2 2
7 0 9 14 13 0 9 2
20 2 0 15 9 13 2 16 2 1 10 9 9 3 15 4 13 12 9 2 2
5 13 1 12 9 2
15 9 11 11 13 9 1 9 1 9 1 9 1 0 9 2
10 9 13 1 3 1 0 9 1 11 2
17 15 14 15 13 1 9 1 9 7 0 9 1 11 1 0 9 2
5 9 13 9 1 11
33 1 9 15 13 9 1 9 9 12 12 2 0 1 0 9 2 14 13 0 0 9 1 9 1 2 11 2 1 9 1 0 9 2
4 13 9 1 11
2 11 11
8 15 13 1 0 9 7 9 2
16 9 1 9 1 9 7 9 1 9 7 9 1 9 1 9 2
6 0 9 1 9 1 9
14 15 13 9 1 9 1 9 2 15 0 9 13 3 2
9 0 9 13 1 1 12 9 9 2
10 3 9 14 4 13 1 0 0 9 2
12 3 9 1 9 13 14 13 9 15 1 9 2
12 3 9 2 15 13 9 2 4 13 1 9 2
11 1 9 1 11 14 13 1 12 9 9 2
8 2 11 2 13 3 1 0 9
5 0 9 13 0 2
18 15 13 0 9 2 7 0 13 2 16 15 13 1 9 1 0 9 2
21 0 9 4 13 1 0 9 1 0 0 9 2 11 2 11 11 2 13 11 3 2
5 12 0 9 15 13
4 9 13 0 9
32 1 9 1 11 2 9 4 4 13 7 13 1 12 9 1 12 9 9 2 1 1 9 15 15 13 1 9 1 0 9 11 2
5 1 15 13 9 2
7 9 11 11 13 1 9 2
16 3 0 9 11 11 15 4 13 1 0 9 14 13 12 9 2
11 11 11 2 12 9 2 2 9 2 11 2
14 3 3 15 13 14 13 0 2 3 10 6 15 13 2
9 16 15 13 3 2 4 13 0 2
13 9 1 12 9 1 11 11 13 9 1 12 9 2
20 9 15 15 13 1 9 1 9 7 13 9 2 15 13 1 9 1 0 9 2
34 11 11 13 9 15 1 9 2 0 11 2 2 1 14 13 0 9 1 0 9 2 15 9 1 2 11 2 13 1 9 1 0 9 2
7 2 6 2 14 15 13 2
4 2 3 6 2
14 11 11 13 1 9 3 1 0 9 2 7 11 13 2
19 2 11 2 15 13 1 0 9 11 11 2 15 13 14 13 3 1 9 2
23 1 14 13 1 15 2 9 7 0 9 15 13 1 2 11 11 2 12 3 9 1 0 2
15 3 13 9 7 3 6 15 13 1 0 0 9 1 9 11
14 1 10 9 1 0 9 9 13 7 1 12 12 9 2
16 9 1 9 4 13 1 9 1 0 9 2 13 1 0 9 2
7 13 11 1 9 12 9 2
6 13 9 1 0 9 3
7 9 13 11 0 1 9 2
20 0 9 1 11 13 0 0 9 2 13 3 9 1 0 0 9 9 11 11 2
18 9 1 9 13 0 9 1 9 1 0 9 2 13 9 1 0 9 2
4 9 1 0 9
11 9 13 12 9 2 12 9 7 12 9 2
7 13 7 9 2 13 15 2
39 0 9 4 13 1 0 9 1 0 9 2 7 1 0 9 4 15 13 1 12 9 7 9 2 1 9 1 15 1 12 9 2 9 2 13 1 12 9 2
21 10 1 9 6 15 13 2 16 13 9 1 9 2 10 9 13 1 12 9 9 2
40 0 1 9 7 9 0 9 14 13 1 9 1 9 7 9 2 1 9 1 9 7 1 0 9 2 3 7 1 9 1 9 1 10 9 7 9 1 0 9 2
7 9 13 9 1 2 11 2
10 13 12 9 9 9 1 11 9 2 12
3 13 9 12
17 1 9 1 0 9 15 13 12 9 3 9 1 9 1 0 9 2
3 13 9 9
5 13 11 1 0 9
29 1 9 2 9 7 9 2 14 13 14 13 1 11 2 1 14 15 13 14 13 1 9 1 9 1 9 1 11 2
13 11 11 2 12 9 2 2 9 1 11 2 11 2
8 13 13 14 13 7 9 15 2
17 13 14 4 13 10 9 1 9 15 1 0 9 7 0 15 9 2
14 11 11 14 15 13 1 9 1 11 11 1 0 9 2
14 9 13 9 1 0 9 7 13 9 14 13 0 9 2
11 11 13 9 1 9 2 9 1 9 9 2
30 11 13 9 15 1 9 0 15 9 7 15 13 1 0 9 2 9 15 13 9 1 0 15 9 2 13 2 9 2 2
20 9 2 15 14 13 9 1 9 2 14 13 3 0 2 16 13 9 1 9 2
14 12 9 1 11 4 13 10 9 7 9 2 13 11 2
11 0 9 14 13 1 0 9 3 1 9 2
5 12 9 15 13 2
6 9 4 13 1 9 2
7 0 9 13 9 1 0 9
15 16 11 13 1 9 2 12 14 13 9 1 0 9 3 2
37 3 1 12 9 13 9 1 0 9 2 1 15 13 0 9 2 9 2 9 2 2 0 2 9 1 9 7 9 7 3 0 9 2 9 7 9 2
14 11 7 11 14 13 0 9 1 11 1 9 1 9 2
5 12 9 15 13 2
21 14 11 6 13 9 2 0 1 12 9 2 16 1 15 13 10 9 1 10 9 2
22 11 14 13 3 9 1 11 2 16 11 6 15 13 14 13 9 1 9 1 0 9 2
16 3 12 9 1 9 1 11 15 13 1 0 9 2 13 9 2
6 9 4 13 1 11 2
6 9 15 13 1 9 15
17 9 15 13 2 1 14 15 13 9 1 9 2 9 7 0 9 2
15 3 4 13 2 3 9 13 1 9 7 15 13 1 12 9
12 12 9 3 13 9 15 1 9 1 10 9 2
19 14 15 13 14 15 13 12 9 1 9 2 13 0 9 7 9 11 11 2
21 1 9 15 9 15 13 9 1 0 9 2 11 11 2 2 1 15 4 13 9 2
38 1 12 9 2 0 1 0 9 1 9 1 0 9 11 11 2 4 13 12 9 2 0 1 0 0 9 2 0 1 9 2 1 0 9 12 9 9 2
20 0 9 2 11 11 2 13 1 11 1 12 9 1 0 15 9 1 0 9 2
18 1 3 1 0 9 1 9 1 11 13 12 0 9 2 0 1 9 2
26 0 9 1 9 13 9 1 9 2 15 13 1 9 2 7 9 1 0 9 1 9 1 9 1 9 2
17 15 13 2 16 9 1 11 11 13 14 14 15 13 1 0 9 2
12 2 15 13 14 14 15 13 1 10 0 9 2
6 9 15 13 1 9 2
25 1 9 1 0 9 14 4 13 7 9 1 9 1 9 7 0 9 2 13 3 9 2 11 2 2
22 12 9 13 1 10 0 0 9 2 13 9 1 11 11 11 2 7 13 14 15 13 2
15 9 1 11 2 9 1 0 9 7 9 13 9 7 9 2
12 11 11 2 12 9 2 2 0 9 2 11 2
8 14 9 1 9 14 13 0 2
18 1 9 1 0 9 11 1 9 1 9 4 13 12 9 1 0 9 2
19 1 9 1 9 0 15 9 13 1 0 9 1 9 9 1 9 1 9 2
23 13 4 9 2 2 0 2 9 2 0 9 2 9 1 0 9 2 0 9 7 0 9 2
6 9 14 13 11 11 2
6 13 0 9 1 11 11
12 15 13 0 9 1 10 9 1 12 9 1 11
14 0 9 1 9 4 13 3 1 0 9 1 0 9 2
10 11 11 15 13 1 15 1 0 9 2
15 11 2 11 13 0 9 1 9 7 9 1 12 9 9 2
21 1 11 15 14 13 1 9 2 3 1 9 1 9 15 13 9 1 9 1 9 2
6 0 9 13 9 1 11
12 13 1 9 2 0 9 2 1 0 0 9 2
18 2 3 13 9 1 0 15 9 2 13 15 15 1 9 1 12 9 2
13 9 13 2 16 1 0 9 0 13 9 1 9 2
4 3 14 13 2
14 9 1 11 11 4 13 10 9 7 0 9 1 9 2
16 3 0 1 0 9 1 10 9 2 3 0 2 0 7 0 2
23 13 14 15 1 15 14 2 13 14 0 15 9 2 15 14 15 13 1 9 14 15 13 2
12 11 14 13 11 1 9 2 11 2 1 11 2
25 1 9 1 9 14 4 13 9 1 9 1 9 1 11 2 11 2 2 13 3 0 9 11 11 2
19 9 15 13 1 9 1 0 11 2 15 13 10 9 7 13 1 1 9 2
22 9 3 1 0 9 1 15 14 15 13 1 9 11 2 9 12 1 9 9 1 9 2
5 11 11 13 1 9
8 9 13 14 15 13 1 9 2
11 11 11 2 12 9 2 2 0 2 11 2
9 14 3 9 14 15 15 13 9 2
9 1 16 10 9 6 13 3 0 2
8 2 11 2 13 1 9 1 9
18 9 13 3 12 9 3 1 11 2 1 14 13 0 9 1 0 9 2
32 1 9 13 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 2 11 11 7 0 2
21 11 11 7 11 11 13 1 9 1 0 0 9 1 2 11 2 1 0 0 9 2
6 11 15 13 1 0 9
13 13 15 1 9 9 2 9 2 9 7 0 9 2
7 14 6 15 13 1 9 2
31 1 0 9 9 1 9 9 1 0 11 7 11 13 1 0 9 1 12 9 1 11 2 11 2 11 2 0 9 7 0 2
19 9 13 1 0 9 1 10 9 14 4 13 9 1 9 1 9 1 9 2
18 9 1 11 3 13 3 0 2 15 1 0 9 13 14 13 1 9 2
24 1 12 9 1 9 9 13 9 1 9 1 3 1 12 9 2 0 1 0 9 1 0 9 2
17 0 9 1 9 2 11 11 2 13 0 9 7 11 1 0 9 2
14 1 15 3 15 13 7 9 7 11 13 0 1 9 2
9 13 0 2 15 6 13 14 13 2
16 1 9 1 11 13 2 16 9 6 13 14 13 9 1 9 2
6 10 9 14 13 15 2
8 11 4 13 1 0 0 9 2
10 2 6 13 3 14 15 13 0 9 2
17 2 1 0 9 13 9 1 9 1 9 2 15 15 13 1 9 2
12 14 13 14 9 1 9 1 0 14 12 9 2
5 2 13 3 9 2
15 2 13 13 14 15 13 2 16 14 13 9 7 1 0 2
4 13 11 1 11
15 10 2 16 15 13 0 2 13 9 3 13 14 13 3 2
21 3 13 2 16 3 0 9 13 14 13 1 2 0 9 2 2 13 1 0 9 2
11 3 13 3 2 15 13 14 13 1 11 2
15 3 4 13 0 9 1 9 2 11 7 9 2 11 2 2
13 16 13 2 16 13 0 2 15 15 13 10 9 2
12 13 1 0 15 9 2 15 3 13 1 9 15
12 0 9 13 1 3 9 2 13 9 1 9 2
19 16 15 6 15 13 2 10 13 1 0 9 2 13 15 9 1 9 11 2
10 15 13 9 1 0 9 9 1 9 2
18 9 15 3 13 0 9 2 15 15 13 9 1 9 2 3 13 9 2
6 13 9 1 12 9 2
17 1 10 9 15 13 14 13 12 9 2 7 0 15 13 1 12 2
8 13 3 2 16 13 14 13 2
11 11 11 2 12 9 2 2 9 2 11 2
5 2 3 13 0 2
20 9 1 0 9 11 11 13 2 16 1 9 6 15 13 1 10 9 1 11 2
18 3 9 4 13 1 9 1 0 9 1 11 11 2 11 2 1 11 2
7 0 9 13 9 1 9 2
11 3 0 9 1 9 13 1 9 1 9 2
11 0 9 13 0 0 9 1 12 9 3 2
15 3 1 9 3 15 13 7 9 1 10 0 7 0 9 2
13 9 1 9 13 1 0 9 2 9 1 9 2 2
20 9 7 0 9 1 11 11 11 4 13 1 9 11 1 9 9 2 13 11 2
8 9 15 13 1 9 1 11 2
15 9 13 9 1 11 2 16 3 4 4 13 1 9 9 2
11 15 1 0 7 0 9 3 3 15 13 2
10 13 10 0 9 1 1 12 12 9 2
15 13 15 2 16 9 13 9 2 15 6 13 14 13 9 2
21 3 1 0 9 4 13 3 12 9 2 16 9 13 1 12 9 3 1 0 9 2
9 13 9 1 0 9 9 1 0 9
17 12 9 13 7 9 1 9 2 15 13 0 9 14 13 9 15 2
25 9 1 9 3 13 3 2 16 3 9 9 2 12 9 2 13 1 9 1 9 12 2 13 11 2
35 13 9 1 9 1 0 0 9 2 0 9 2 0 9 1 0 9 2 3 7 1 9 2 0 1 0 9 2 1 1 0 9 1 9 2
6 9 13 9 1 0 9
9 9 9 2 9 7 9 13 9 2
8 1 9 1 9 13 0 9 2
13 1 0 9 13 7 9 1 9 1 9 11 11 2
7 0 9 13 9 1 9 2
12 0 9 1 0 9 13 0 9 1 0 9 2
11 0 9 1 11 13 9 2 0 11 2 2
10 1 9 1 0 9 13 1 12 9 2
24 9 1 9 4 13 1 9 2 3 9 3 9 2 1 9 1 0 9 2 15 15 13 3 2
24 1 0 9 1 11 1 9 9 13 0 9 1 9 2 1 3 14 13 9 1 2 11 2 2
20 1 10 9 2 1 9 3 2 3 13 9 1 9 2 15 14 15 13 9 2
24 1 15 13 7 0 9 2 16 1 10 9 15 13 0 9 1 9 1 10 9 1 0 9 2
38 9 2 0 1 9 1 0 9 2 10 9 1 9 15 1 9 1 0 9 1 11 2 11 11 2 1 0 9 1 9 13 14 4 13 1 0 9 2
12 3 13 9 1 10 0 0 9 1 0 9 2
7 9 1 9 13 3 0 2
17 2 3 10 9 11 11 13 2 16 9 14 13 1 12 9 3 2
12 2 13 3 9 2 9 7 9 1 10 9 2
11 11 11 2 12 9 2 2 9 2 11 2
16 0 0 9 13 1 0 1 9 9 1 0 9 11 11 11 2
60 9 2 1 9 1 9 2 2 9 1 2 0 9 2 2 9 1 0 0 9 2 9 1 2 9 1 0 9 2 1 0 0 2 0 2 0 9 1 9 2 1 9 2 1 9 7 9 15 13 0 1 0 9 9 1 2 0 9 2 2
32 1 9 12 1 0 9 15 13 12 9 2 7 9 1 9 11 11 2 11 11 2 11 11 7 11 11 14 13 1 0 9 2
20 9 1 11 14 13 0 9 1 0 9 2 11 2 2 13 9 11 11 3 2
27 9 1 0 9 4 13 2 7 9 15 13 1 0 9 7 13 14 15 13 1 0 9 1 2 11 2 2
19 11 11 2 11 15 13 1 0 9 1 9 9 1 11 2 11 11 2 2
17 15 13 7 9 1 9 1 0 9 1 9 14 13 9 1 9 2
21 3 12 9 4 13 9 14 13 1 9 2 0 1 12 9 9 7 12 9 9 2
6 0 9 13 9 7 9
15 3 13 3 2 16 0 9 9 15 13 3 1 0 9 2
19 3 13 9 1 0 9 1 0 9 2 0 1 0 9 11 2 13 9 2
25 1 0 9 1 11 9 1 11 13 14 13 0 9 1 0 9 7 1 0 0 9 2 13 11 2
21 1 9 6 15 13 1 10 14 13 0 9 1 9 2 0 15 1 3 0 9 2
11 7 9 0 9 3 14 13 14 15 13 2
9 1 15 3 0 9 4 3 13 2
6 11 13 14 13 9 11
11 9 4 13 1 9 3 1 3 0 9 2
24 9 1 11 1 0 9 4 13 1 9 1 10 9 2 15 15 4 13 14 15 13 1 9 2
17 1 9 0 9 15 13 12 9 1 9 7 15 13 1 0 9 2
5 3 9 15 13 2
10 9 3 6 13 2 7 9 15 13 2
10 15 13 2 16 11 3 13 14 13 2
10 9 1 0 9 13 1 1 12 9 2
13 0 9 4 13 1 9 2 15 13 1 0 9 2
21 1 9 9 9 4 13 1 9 1 11 7 9 15 11 1 9 2 0 9 2 2
8 9 15 4 13 1 0 9 2
4 3 13 9 2
10 9 1 9 2 11 2 15 13 1 9
20 1 0 9 9 2 11 2 2 1 15 12 13 0 9 2 15 13 1 15 2
10 9 1 0 9 1 0 9 13 0 9
17 16 15 13 1 9 1 9 2 9 13 9 14 13 0 7 0 2
15 10 9 3 13 0 2 3 16 13 9 1 10 0 9 2
22 2 13 9 1 9 1 2 11 2 2 9 2 15 13 0 9 14 13 1 0 9 2
11 7 13 9 1 9 1 9 2 1 9 2
7 14 13 1 11 1 0 9
10 0 9 13 1 9 15 1 9 1 9
5 11 13 9 1 11
15 1 0 9 1 11 11 7 11 11 3 14 13 0 9 2
12 11 11 15 13 1 9 0 9 1 11 12 2
24 1 0 9 1 0 9 14 15 13 10 0 9 2 0 1 9 2 2 9 1 2 11 2 2
10 11 13 2 1 14 15 4 13 3 2
4 2 3 14 2
11 13 15 1 0 3 9 1 9 1 9 2
5 10 14 6 13 2
23 9 3 13 0 9 2 9 15 13 7 15 13 1 9 2 9 7 9 15 13 1 9 2
16 9 13 9 1 11 1 9 15 1 9 1 2 0 9 2 2
13 1 9 1 9 15 15 15 13 7 13 0 9 2
15 1 9 1 9 14 15 13 2 14 11 14 13 1 15 2
31 11 7 11 2 9 2 15 13 1 9 2 11 13 1 9 1 9 2 7 9 1 2 11 2 11 13 0 9 1 9 2
23 1 9 1 11 11 15 13 10 0 9 7 9 2 15 3 13 14 4 13 1 0 9 2
16 1 0 9 3 13 9 2 15 6 13 14 13 9 1 9 2
10 1 15 14 13 9 2 9 7 9 2
10 9 15 3 13 9 7 6 15 13 2
11 2 7 13 14 13 0 9 1 0 9 2
17 9 13 0 9 2 0 9 2 9 2 0 9 7 0 9 2 2
23 1 0 9 13 12 9 1 11 1 12 9 7 12 9 1 0 9 1 0 9 1 11 2
73 3 1 9 13 11 11 2 11 11 2 11 11 2 11 11 2 11 2 11 11 2 7 3 7 9 2 0 9 2 2 2 11 2 2 2 11 2 2 2 11 11 11 2 2 2 11 2 2 11 11 2 11 2 11 2 11 11 2 11 11 7 11 11 7 0 9 1 9 2 9 7 9 2
22 1 0 9 2 1 9 1 0 9 2 13 9 0 15 9 14 15 13 1 0 0 9
35 1 15 15 13 6 3 1 9 1 0 0 9 2 6 3 1 9 1 9 2 7 7 1 9 1 0 1 15 9 1 0 9 7 11 2
11 9 1 0 9 13 9 1 0 9 11 11
13 11 14 13 1 10 9 1 12 1 0 0 9 2
31 15 13 9 1 11 7 1 9 15 13 1 9 1 10 0 9 7 9 2 15 13 2 16 14 13 1 9 1 9 15 2
14 10 9 13 2 3 13 9 1 0 9 2 13 15 2
20 1 11 11 3 3 0 9 13 14 13 0 0 9 1 9 1 0 15 9 2
15 9 1 9 1 9 1 0 9 13 1 9 1 0 9 2
21 0 9 11 11 13 2 16 9 13 4 13 3 7 13 9 1 9 1 0 9 2
14 9 13 10 9 2 16 9 15 11 13 9 1 9 2
20 11 11 2 11 11 2 11 11 2 11 11 7 11 11 13 1 9 1 9 2
19 0 9 11 11 2 9 1 9 11 11 2 13 0 9 1 9 1 9 2
34 1 0 9 1 12 9 1 9 1 0 9 1 11 7 1 9 2 16 0 9 11 11 3 6 4 4 13 13 9 15 9 1 11 2
14 1 9 2 1 15 9 1 0 9 4 13 11 11 2
20 1 15 13 3 14 13 9 1 9 11 11 2 15 3 13 12 9 1 9 2
6 13 4 9 1 11 2
12 11 3 14 13 0 9 2 1 14 13 9 2
21 9 4 13 1 12 9 7 4 13 1 12 1 12 9 1 12 9 1 12 9 2
35 11 3 6 13 9 15 1 9 1 9 1 9 1 0 9 2 11 7 11 7 6 15 13 1 14 12 1 9 1 9 1 9 7 9 2
15 13 3 14 15 13 0 9 1 10 9 1 9 1 9 2
12 2 13 1 11 7 9 11 6 13 14 13 2
10 15 13 0 9 2 15 4 15 13 2
6 2 10 13 3 3 2
8 1 3 3 4 13 1 9 2
6 2 15 13 10 9 2
8 11 11 13 9 1 9 1 11
11 7 11 13 2 9 13 0 9 1 9 2
20 15 6 4 13 1 9 2 7 0 9 13 0 9 1 0 9 1 10 9 2
10 1 15 0 9 1 0 9 13 9 2
20 0 9 1 9 4 15 13 3 1 11 2 11 2 7 11 11 2 11 2 2
27 0 9 11 11 13 3 1 9 1 0 9 1 2 11 11 11 11 2 1 11 7 11 2 13 9 11 2
9 1 10 9 1 9 2 11 3 13
10 4 13 3 7 9 1 9 1 9 2
14 9 15 13 1 0 9 2 3 15 13 3 12 9 2
24 15 14 6 4 13 1 9 1 9 1 2 11 2 10 9 1 0 9 1 9 2 11 2 2
3 9 2 11
21 3 3 13 9 1 9 2 9 2 2 3 3 14 4 13 9 1 2 11 2 2
16 1 15 1 0 9 1 9 13 9 11 11 7 9 11 11 2
25 13 14 4 13 0 0 9 2 15 14 15 13 1 9 1 9 1 0 11 1 9 2 11 2 2
22 9 14 13 1 0 9 1 0 9 1 0 9 2 13 9 1 9 7 9 11 11 2
8 11 13 3 9 1 12 9 9
12 6 15 13 3 3 4 4 13 2 11 2 2
13 3 12 9 14 13 9 1 9 7 9 1 9 2
25 0 9 15 13 1 9 1 9 15 2 11 2 0 9 2 1 1 13 14 13 1 9 1 11 2
8 15 13 0 15 9 1 11 2
8 10 9 13 10 0 0 9 2
4 9 2 11 11
22 3 13 2 16 13 14 13 14 13 9 1 3 1 9 2 7 1 9 13 1 9 2
10 7 3 6 4 13 9 1 0 9 2
20 1 9 2 0 1 11 2 11 2 2 13 9 7 0 9 1 0 15 9 2
7 13 1 9 0 0 9 2
18 11 11 13 2 16 1 9 15 2 9 1 9 2 13 3 0 9 2
14 0 9 2 15 15 13 2 13 9 1 10 0 9 2
13 9 4 13 9 1 9 1 9 1 9 12 9 2
22 1 9 9 1 9 1 0 0 9 2 0 1 0 9 2 13 0 9 1 10 9 2
8 9 1 9 11 13 3 0 2
10 1 9 15 13 12 9 9 1 9 2
16 9 7 9 15 14 13 9 15 1 9 11 2 3 1 11 2
8 12 9 13 9 1 0 9 2
5 9 13 9 1 0
10 12 9 3 13 2 16 6 13 0 2
24 0 9 1 2 0 9 2 1 0 9 2 0 11 2 2 3 13 12 9 2 13 12 9 2
6 11 13 11 1 9 3
21 15 13 2 3 0 2 0 7 3 0 0 9 2 2 1 14 13 9 1 9 2
6 13 4 9 7 9 2
11 0 15 13 1 9 7 6 13 1 9 2
12 3 15 13 3 14 15 13 7 9 1 9 2
13 3 11 14 13 0 9 1 11 1 10 0 9 2
28 1 9 1 9 1 11 2 15 13 9 15 1 0 9 2 1 14 15 13 0 9 2 11 13 0 1 9 2
16 3 7 2 0 2 9 1 9 1 10 9 7 9 1 0 2
11 9 13 12 0 9 2 0 9 1 11 2
6 9 15 13 1 0 2
7 3 13 14 13 1 9 2
11 11 3 15 13 2 14 13 14 13 0 2
8 3 13 9 1 9 1 9 2
4 13 0 9 2
13 1 9 1 0 9 7 0 9 0 9 13 0 2
9 1 0 9 15 13 3 0 9 2
8 0 9 13 7 1 0 9 2
18 10 10 0 9 3 13 14 13 1 9 2 11 11 2 1 12 9 2
13 9 15 13 2 16 1 9 13 0 2 11 2 2
10 1 11 12 4 13 1 3 0 9 2
4 3 13 9 2
11 1 0 9 15 13 14 13 9 0 9 2
15 9 13 9 1 9 1 9 2 11 2 1 9 1 9 2
9 1 0 9 13 7 9 1 9 2
22 0 9 4 13 1 9 1 0 9 2 1 16 9 4 13 3 1 0 9 0 9 2
6 11 13 9 2 11 2
11 3 0 9 1 9 1 9 13 0 9 2
9 9 14 15 13 3 1 0 9 2
4 9 1 0 9
16 0 9 2 0 9 2 9 1 0 9 2 9 1 9 1 11
15 0 1 9 7 9 15 13 1 9 2 9 7 0 9 2
14 3 6 13 3 0 15 14 15 13 1 0 0 9 2
28 1 9 2 0 9 1 9 15 1 9 2 9 15 13 1 9 2 11 2 2 3 13 7 15 13 1 9 2
27 0 9 1 2 11 11 11 2 11 4 13 1 9 1 0 9 1 0 9 1 0 9 2 11 11 2 2
25 12 9 1 15 15 4 13 9 14 15 13 1 2 11 2 2 1 14 15 13 0 9 1 9 2
26 1 0 9 15 13 9 2 11 11 2 7 2 11 11 11 2 7 2 11 11 2 7 2 11 2 2
6 13 0 9 1 11 11
11 1 9 13 7 9 2 0 1 0 9 2
11 1 0 1 12 9 9 1 9 13 11 2
5 13 9 1 0 9
27 0 7 0 9 13 0 1 15 0 9 2 0 9 2 0 9 2 0 9 2 0 9 2 9 2 9 2
21 1 0 9 4 13 9 1 9 2 11 2 11 2 1 0 9 1 0 9 3 2
12 15 13 1 12 9 1 9 15 1 0 9 2
14 12 9 15 13 1 0 9 1 0 9 1 0 9 2
15 9 4 13 1 9 1 9 1 0 7 0 9 1 11 2
22 1 11 12 9 4 13 7 1 12 4 13 1 9 2 0 1 0 9 2 13 11 2
18 1 9 1 15 9 14 13 0 9 3 1 9 1 9 2 13 9 2
6 9 2 9 2 11 2
11 2 0 0 9 14 15 13 1 0 9 2
17 7 16 13 2 16 10 9 13 0 2 1 10 0 9 15 13 2
15 3 2 3 1 0 9 1 0 9 9 6 13 1 9 2
29 0 9 1 11 7 2 11 2 11 11 2 1 9 2 13 9 2 0 1 10 9 1 9 11 1 0 9 9 2
21 1 9 9 13 11 11 2 0 1 11 11 2 11 11 2 11 11 7 11 11 2
8 9 13 1 9 2 13 11 2
6 11 11 13 9 1 9
8 9 15 13 1 12 9 9 2
9 9 1 11 4 13 0 15 9 2
7 13 14 3 0 0 9 2
14 15 13 2 16 15 13 0 9 7 3 14 13 9 2
14 7 6 3 16 13 14 13 1 9 2 7 14 13 2
15 15 11 13 1 0 0 9 2 3 15 13 9 1 9 2
10 1 0 9 0 9 13 0 1 9 2
4 3 13 15 2
11 16 9 15 13 2 14 13 9 1 12 9
4 3 6 13 9
7 2 15 13 9 1 9 2
24 1 9 2 11 2 12 9 13 2 16 15 13 0 0 9 1 9 1 9 1 9 7 9 2
7 9 6 13 0 7 0 2
19 3 1 0 9 13 7 0 9 1 9 1 9 1 11 1 9 1 9 2
24 1 9 2 1 0 9 0 9 11 3 13 9 1 2 11 2 1 0 9 1 12 9 9 2
11 11 11 2 9 1 0 9 1 9 1 9
30 1 9 1 9 15 14 4 13 7 0 0 9 1 9 1 9 1 0 0 9 1 11 2 11 7 11 1 0 9 2
23 1 15 15 13 0 9 2 0 9 2 7 10 9 2 0 9 7 9 2 2 13 11 2
20 9 1 9 6 13 0 7 6 13 9 2 13 9 11 2 0 9 1 11 2
16 9 2 9 1 9 2 13 7 9 1 9 15 1 0 9 2
18 0 9 13 9 1 0 9 7 9 1 9 1 9 1 9 7 9 2
21 9 14 13 14 13 9 1 10 9 1 0 9 2 3 7 1 9 1 0 9 2
18 13 4 7 0 9 1 9 2 15 13 1 9 1 9 2 13 9 2
22 2 0 0 9 1 9 2 0 9 2 13 9 1 0 9 1 9 2 2 13 11 2
19 1 10 0 9 15 13 14 13 0 9 1 11 2 13 9 1 12 9 2
2 11 11
24 9 13 1 9 1 9 2 16 13 0 9 1 11 1 9 1 9 12 9 2 13 1 11 2
17 1 9 1 9 1 11 9 1 9 15 13 1 0 9 1 11 2
22 0 9 11 11 14 13 11 1 0 9 1 9 12 9 1 11 7 9 11 2 11 2
12 1 12 4 13 0 9 2 1 14 13 9 2
15 6 4 13 9 1 9 1 11 11 2 3 15 13 9 2
8 15 13 1 0 0 9 1 11
19 11 13 12 9 1 9 1 9 2 11 11 11 2 7 2 11 2 11 2
21 9 1 9 13 9 1 9 1 9 2 1 9 1 9 1 0 15 9 1 3 2
16 1 9 2 9 1 2 11 2 12 4 4 13 1 0 9 2
17 2 15 13 14 2 16 13 14 15 13 3 9 1 11 7 11 2
7 2 15 15 13 10 9 2
26 3 1 9 1 10 9 9 4 4 13 7 1 9 1 0 9 1 0 9 2 15 3 13 11 11 2
8 3 13 9 2 15 15 13 2
15 13 14 13 0 15 9 1 0 9 1 11 2 13 15 2
7 9 1 11 13 3 9 15
27 15 3 4 13 9 1 0 9 2 1 10 2 16 1 9 15 1 9 15 4 13 0 9 7 0 9 2
15 3 9 13 2 16 1 0 15 9 13 9 1 0 9 2
13 3 9 1 9 13 1 9 1 9 15 1 9 2
23 10 0 0 9 13 9 1 11 1 9 1 9 11 11 1 9 1 0 9 2 13 11 2
8 9 1 0 13 1 10 9 2
13 15 13 1 11 1 11 7 13 1 9 1 11 2
10 0 9 1 9 1 9 3 13 0 2
8 11 14 13 1 11 1 0 9
31 3 9 11 15 13 1 9 1 11 11 11 2 1 9 1 0 9 1 11 11 11 7 1 11 11 2 9 1 0 9 2
7 9 15 13 10 0 9 2
24 3 10 9 14 4 13 0 0 9 2 13 9 11 11 1 0 15 9 1 0 9 1 9 2
2 11 2
24 11 11 4 13 1 0 9 1 9 1 11 1 9 1 9 9 1 9 1 0 9 11 11 2
11 1 9 1 9 13 7 2 11 11 2 2
10 7 13 15 14 15 13 1 0 9 2
25 3 3 2 16 3 6 13 3 14 11 14 13 15 14 15 4 13 7 3 11 14 13 1 15 2
5 9 7 9 13 11
14 1 0 9 3 15 13 2 16 0 9 13 0 9 2
21 1 12 9 0 9 1 9 2 11 2 1 9 9 15 13 1 0 9 1 11 2
22 12 15 0 9 9 7 11 11 11 11 11 4 13 1 9 2 0 1 12 12 9 2
13 0 9 3 4 13 3 9 7 1 9 11 11 2
15 3 15 4 13 1 11 1 0 15 9 7 0 15 9 2
13 9 2 0 9 2 15 13 3 9 1 0 9 2
20 0 11 7 9 3 13 0 9 7 15 13 1 9 2 0 1 9 10 9 2
23 7 15 13 1 10 9 3 1 9 2 15 15 13 0 9 2 15 3 15 13 3 3 2
24 7 3 16 15 13 2 16 13 0 2 13 3 14 4 13 1 15 1 1 2 0 9 2 2
9 9 1 11 11 13 9 1 0 9
24 13 4 9 1 9 2 15 13 9 1 0 9 1 9 2 9 1 0 9 2 0 1 9 2
8 0 9 15 13 1 11 7 11
18 15 14 15 13 1 11 7 14 4 13 1 9 1 9 1 10 9 2
10 3 1 15 15 13 9 1 0 9 2
19 3 15 13 2 3 15 6 15 13 3 1 9 2 1 14 4 13 9 2
5 15 13 12 9 2
24 3 2 16 13 1 9 7 15 13 2 16 13 1 9 2 15 13 1 9 14 15 13 3 2
12 0 0 9 1 9 4 13 3 1 10 9 2
15 13 2 16 9 1 0 9 11 11 2 11 14 13 9 2
13 2 3 14 13 10 9 14 15 13 1 0 9 2
5 2 16 13 9 2
19 2 16 15 13 1 9 7 1 0 9 1 10 9 1 9 1 0 9 2
9 3 15 4 13 1 0 0 9 2
24 2 9 1 0 9 1 9 16 16 13 0 9 1 15 7 13 0 9 1 10 9 1 11 2
5 2 3 2 6 2
12 3 15 13 10 3 0 9 1 0 15 9 2
29 3 11 3 15 13 1 0 0 9 2 7 9 15 1 0 9 4 13 1 9 3 1 11 11 1 0 0 9 2
9 0 9 1 0 9 13 0 9 2
14 3 1 9 1 0 9 1 11 13 14 13 3 3 2
15 1 0 1 0 9 9 9 1 0 9 13 0 0 9 2
30 1 9 1 0 0 9 7 9 1 9 1 11 11 7 11 11 1 0 9 13 9 1 9 1 0 9 1 0 9 2
13 1 9 1 9 9 1 0 0 9 13 12 9 2
17 0 9 13 15 14 13 2 16 6 13 9 1 10 9 7 9 2
17 3 1 9 11 13 1 12 0 9 2 1 15 4 13 9 9 2
18 9 3 15 13 1 11 2 11 2 11 7 11 2 16 9 13 0 2
15 0 13 0 9 1 9 2 1 14 15 13 3 0 9 2
8 1 1 9 15 13 1 9 2
12 1 12 9 1 9 13 2 7 6 13 0 2
14 11 4 13 9 2 15 13 1 0 9 1 0 9 2
17 9 1 9 11 1 11 11 11 14 13 3 9 15 1 0 9 2
17 1 9 1 9 15 13 14 15 13 7 9 1 10 9 11 11 2
18 9 13 2 16 9 1 11 11 7 11 11 1 9 1 11 15 13 2
14 1 9 1 0 0 9 1 11 9 1 9 13 0 2
9 0 9 1 11 13 9 1 9 2
11 13 14 13 12 11 7 12 9 1 11 2
29 0 9 13 9 15 1 10 9 7 1 9 15 13 9 2 1 15 4 15 13 1 0 9 2 13 0 0 9 2
16 9 7 9 3 6 13 14 15 13 0 14 13 9 1 11 2
6 14 9 6 13 1 9
7 15 13 9 1 10 9 2
25 2 9 1 9 9 11 13 2 16 1 10 9 11 6 4 13 10 0 0 9 1 9 1 9 2
28 7 14 14 15 13 3 14 15 13 15 1 9 2 1 10 0 9 2 16 13 14 13 9 7 14 13 9 2
22 0 9 1 11 6 4 13 1 0 9 7 3 13 2 6 4 13 7 1 0 9 2
6 6 13 14 15 13 2
25 16 13 0 9 1 9 1 9 1 9 7 15 13 10 0 9 2 9 15 4 13 10 0 9 2
21 9 1 9 1 9 7 9 1 9 1 9 1 9 7 9 13 0 0 9 3 2
26 13 4 7 9 1 0 9 2 10 9 15 13 1 0 9 1 0 0 9 2 0 9 6 4 13 2
9 9 13 7 0 9 1 0 11 2
27 1 9 1 9 9 1 0 9 1 0 9 7 1 9 11 4 13 3 1 0 9 7 9 1 11 11 2
18 3 1 9 1 9 9 13 9 1 0 0 9 11 2 9 11 11 2
21 9 11 13 14 13 9 1 0 9 2 3 2 1 14 6 13 9 1 11 11 2
15 3 6 15 13 2 13 2 16 9 6 15 13 1 15 2
33 11 15 13 1 9 11 2 3 3 13 0 9 1 0 15 9 1 9 1 9 1 12 9 2 9 1 0 0 9 2 13 11 2
23 3 11 15 13 1 9 1 0 9 1 11 2 1 14 13 9 1 0 9 2 13 11 2
9 11 13 14 4 13 3 1 11 2
11 9 15 13 1 9 1 0 9 1 11 2
18 1 9 9 4 4 13 1 0 9 2 16 4 13 1 9 11 11 2
22 12 9 4 13 1 2 0 9 2 2 13 9 1 9 7 9 11 11 1 9 11 2
13 9 1 9 7 9 1 9 3 13 10 0 9 2
13 15 13 1 9 15 9 1 9 7 13 1 9 2
6 9 1 0 9 13 2
19 13 14 13 2 16 15 4 15 13 1 10 9 2 15 6 13 1 15 2
7 0 13 2 16 13 10 2
14 3 13 0 7 0 9 2 10 0 9 14 4 13 2
11 10 9 15 13 12 1 0 9 1 9 2
28 6 2 10 9 2 15 1 10 9 15 13 2 16 13 1 15 7 13 2 16 10 9 6 15 13 1 15 2
11 9 2 3 0 2 1 9 13 1 13 2
10 15 13 0 9 2 3 6 13 10 2
6 9 13 9 1 9 2
8 1 10 9 13 2 13 3 2
10 13 4 3 3 10 0 9 7 9 2
29 0 9 13 9 15 1 9 1 9 7 13 2 16 11 14 13 0 9 1 11 1 9 1 9 1 9 1 11 2
8 13 1 0 9 14 15 13 2
5 10 13 10 9 2
19 1 10 9 13 9 1 9 1 0 9 2 9 7 9 15 13 1 9 2
10 3 16 3 3 13 10 2 15 13 2
24 1 9 7 9 1 15 4 13 3 9 2 1 15 13 14 13 0 9 7 9 1 0 9 2
8 10 13 9 15 1 10 9 2
18 13 15 1 0 9 2 16 10 9 1 9 13 0 2 0 7 0 2
61 10 9 4 15 13 14 6 15 13 1 9 1 10 9 2 3 7 1 3 0 9 14 13 2 3 14 15 13 1 0 9 2 7 1 9 2 1 9 15 1 9 2 15 1 9 13 14 15 13 3 1 9 2 1 14 13 1 9 1 15 2
7 14 9 7 1 0 9 2
9 15 3 15 13 1 9 1 9 2
9 10 13 9 1 9 1 0 9 2
11 10 13 9 1 9 1 9 1 0 9 2
12 10 13 10 9 1 9 7 9 1 10 9 2
14 0 9 13 14 1 9 15 3 9 1 9 1 9 2
17 2 10 13 9 15 1 9 1 0 9 7 1 9 1 0 9 2
29 1 0 9 1 9 4 13 2 16 11 2 15 1 9 13 11 2 4 13 11 14 13 1 9 1 9 1 9 2
28 13 15 14 13 2 16 1 9 1 10 0 7 0 9 1 11 7 11 0 3 13 14 15 13 1 0 9 2
46 14 13 3 3 2 16 1 0 12 9 9 4 13 3 0 0 9 2 7 1 9 1 0 9 15 13 9 1 9 1 0 9 1 9 1 9 7 15 13 1 9 1 9 1 9 2
20 15 6 13 10 9 13 15 2 10 13 10 9 2 10 9 7 10 9 13 2
24 2 3 13 14 15 13 2 16 6 4 13 14 13 3 9 2 1 9 14 4 13 1 9 2
11 10 13 9 1 9 1 9 1 10 9 2
19 13 15 14 6 13 3 0 0 9 1 9 2 15 4 15 13 1 9 2
21 0 13 2 16 12 7 0 0 9 13 3 0 7 13 1 9 15 10 0 9 2
14 9 3 3 15 13 7 9 13 1 0 9 1 9 2
23 16 13 0 9 2 11 11 15 13 2 16 6 13 2 13 2 13 7 6 13 14 13 2
20 15 13 14 13 1 9 1 9 2 1 15 15 13 3 2 1 9 7 9 2
8 13 9 1 9 1 0 9 2
25 10 2 15 1 9 1 9 1 0 12 9 3 13 9 1 9 1 9 1 9 1 9 1 9 2
19 10 9 7 9 1 9 13 9 1 9 7 9 1 9 2 1 15 13 2
30 0 9 15 13 1 0 9 1 0 9 1 9 1 0 9 1 0 9 7 0 9 1 9 7 9 2 13 3 9 2
13 2 3 0 9 14 13 9 1 10 1 9 3 2
20 13 15 10 9 7 15 15 13 2 16 13 10 2 7 1 3 10 15 13 2
17 7 15 1 10 9 3 13 7 6 1 3 15 13 1 9 15 2
16 2 13 15 11 2 13 9 7 13 9 1 9 1 9 15 2
13 13 15 14 13 1 9 15 7 15 14 15 13 2
17 7 15 3 1 10 9 13 0 9 2 13 15 9 7 9 15 2
11 0 9 13 1 10 9 0 7 0 9 2
22 9 1 0 0 9 15 13 2 1 1 15 15 13 3 1 9 2 1 15 4 13 2
22 13 2 16 9 1 0 9 3 4 13 2 7 9 1 0 0 9 3 3 13 0 2
11 3 13 14 13 1 9 2 15 4 13 2
14 6 13 2 3 2 16 13 10 2 15 13 14 13 2
12 13 3 14 13 9 1 9 2 9 7 9 2
15 2 9 1 0 2 15 13 10 9 2 6 13 1 3 2
55 15 13 2 16 1 0 9 10 9 9 13 1 9 1 11 9 1 9 2 1 14 15 13 1 0 9 1 0 9 2 13 14 13 10 0 9 1 0 9 7 3 13 0 9 2 15 13 12 9 7 3 6 4 13 2
25 3 3 2 7 6 1 0 9 2 3 1 0 9 2 15 13 14 13 9 15 14 13 1 9 2
14 0 9 13 9 1 10 2 15 4 13 9 7 9 2
8 14 12 9 1 9 1 9 2
9 2 13 14 15 13 1 0 2 2
17 0 13 14 15 13 14 13 10 9 2 15 3 13 14 15 13 2
8 2 15 13 12 1 0 9 2
22 2 11 11 2 3 13 14 13 1 9 9 2 13 0 9 1 9 1 15 11 11 2
23 1 0 0 9 4 13 12 9 1 11 1 10 9 2 1 9 16 13 1 0 15 9 2
25 9 2 15 13 14 13 0 15 9 7 14 13 9 1 9 15 2 4 13 0 0 9 11 11 2
26 13 14 13 0 9 10 9 7 9 4 13 10 9 14 13 2 16 14 13 9 1 9 1 9 1 9
28 15 15 13 1 9 1 0 9 1 11 2 7 13 14 13 15 13 9 7 15 4 13 2 9 2 1 9 2
18 9 1 0 9 1 9 14 4 13 2 13 1 9 1 9 1 11 2
14 9 1 11 13 9 1 9 1 9 1 2 11 2 2
24 10 9 13 14 13 12 9 9 2 16 9 6 4 13 1 9 12 9 9 0 9 10 9 2
18 3 10 12 9 2 7 14 3 1 0 9 13 14 13 9 1 9 2
25 1 0 9 1 0 9 15 13 0 9 2 11 2 2 15 1 0 9 13 9 1 9 0 9 2
15 0 1 9 9 6 13 1 9 1 9 10 9 1 9 2
26 1 9 1 0 9 11 4 13 9 15 14 13 1 9 0 9 9 1 10 9 7 9 1 0 9 2
10 9 13 1 9 9 1 12 9 9 2
11 13 0 9 1 2 11 2 1 9 1 9
11 2 9 13 14 13 10 9 1 0 9 2
15 9 11 13 9 2 7 11 13 0 9 1 12 1 12 2
13 9 4 13 1 11 12 9 9 1 9 7 9 2
13 15 13 1 9 1 11 3 9 1 9 11 11 2
18 12 13 3 0 9 1 11 1 9 2 13 3 1 0 2 9 2 2
12 14 15 13 9 7 14 15 13 14 15 13 2
20 2 11 2 13 9 1 9 1 0 9 11 11 1 9 1 9 2 11 2 2
23 2 3 13 2 13 1 0 9 1 0 15 12 9 1 11 2 13 9 15 3 11 11 2
30 16 13 14 13 1 9 2 15 13 14 13 3 2 16 6 4 13 2 6 13 1 9 7 6 4 13 9 1 11 2
17 0 9 13 1 9 0 9 1 12 9 1 9 2 15 13 3 2
8 14 13 9 1 11 1 0 9
6 2 13 0 0 9 2
5 2 13 11 11 2
27 14 15 13 2 16 3 13 0 2 14 13 2 14 13 12 9 2 14 15 13 10 9 7 3 14 13 2
12 1 9 9 13 1 9 1 0 9 1 11 2
15 3 1 15 9 1 11 11 11 13 9 1 9 1 9 2
22 3 13 3 0 9 14 15 13 9 1 9 1 0 11 1 15 2 13 9 12 2 2
5 14 0 15 9 2
16 0 12 1 12 1 9 13 1 9 1 9 2 13 1 9 2
5 14 13 7 15 2
23 9 13 1 0 9 1 9 15 14 13 1 9 9 1 0 1 11 9 1 0 0 9 2
24 9 1 9 1 11 4 13 1 9 1 2 0 11 2 9 1 9 1 9 1 12 12 9 2
8 2 13 9 1 9 11 11 2
6 2 13 3 11 2 2
26 15 9 3 13 1 3 0 9 2 15 14 3 13 2 3 15 13 0 9 1 9 1 9 7 9 2
16 1 9 15 13 14 13 0 15 9 1 9 2 0 9 2 2
25 1 9 9 1 11 9 11 13 14 15 13 9 1 9 2 15 4 15 13 6 1 9 1 9 2
17 2 9 11 2 3 13 1 0 0 9 9 1 9 1 0 9 2
8 12 1 0 13 1 0 9 2
29 3 13 2 16 15 13 9 15 1 9 2 3 14 13 9 15 1 9 1 0 15 9 1 0 9 7 9 15 2
12 9 13 2 16 9 10 9 14 13 3 0 2
19 6 13 1 9 7 9 2 16 10 9 13 12 1 0 9 1 0 9 2
7 9 7 9 13 9 1 11
20 3 0 11 13 1 9 1 0 9 0 9 11 7 13 9 1 0 9 11 2
13 14 14 13 9 7 14 13 9 1 11 7 11 2
30 1 0 9 1 9 9 1 9 1 11 11 11 13 3 14 4 13 1 0 9 10 0 9 2 15 4 13 1 11 2
29 9 13 7 13 2 1 9 15 13 0 9 9 2 9 13 2 14 15 9 2 0 0 9 1 11 2 9 13 2
21 9 4 13 1 0 9 1 11 7 13 9 12 1 0 9 2 0 1 9 15 2
60 14 6 13 2 16 3 13 14 15 13 1 0 9 7 0 9 2 0 9 13 14 15 13 0 2 0 9 2 15 13 0 9 1 9 7 15 13 3 1 10 9 7 3 2 1 10 0 0 9 2 15 13 1 9 15 2 13 9 11 2
46 16 3 1 0 9 1 9 1 0 9 15 13 10 9 1 9 2 14 9 1 10 9 13 0 9 2 13 10 9 9 11 11 2 15 13 0 9 1 9 2 11 11 2 1 11 2
37 3 15 13 1 9 1 10 9 2 13 3 14 15 13 2 16 12 1 9 2 15 13 9 1 10 9 2 13 11 2 13 0 9 1 9 15 2
40 3 16 9 1 9 13 1 11 7 9 1 9 1 9 15 13 1 11 2 16 15 13 7 15 13 2 14 13 14 13 0 9 2 0 1 11 2 13 11 2
51 1 9 1 0 11 4 13 2 16 2 4 13 9 1 11 1 0 9 2 2 13 1 0 9 1 9 1 9 1 0 9 2 2 13 15 4 1 9 2 2 7 9 15 6 13 1 9 1 9 2 2
4 2 13 11 2
25 3 13 14 13 1 11 2 1 15 3 14 15 13 1 15 2 15 3 1 9 6 4 13 0 2
22 14 15 15 13 14 15 13 0 9 1 15 2 1 14 15 13 10 13 0 15 9 2
8 15 1 10 9 13 1 11 2
18 6 13 14 13 10 9 2 3 9 14 13 2 3 1 11 13 1 15
4 2 13 11 2
19 1 11 13 14 15 13 7 0 9 1 10 9 2 1 15 4 13 9 2
12 9 4 13 1 0 9 1 0 9 1 11 2
4 2 13 9 2
22 9 13 14 15 13 9 1 9 2 15 1 9 4 13 0 9 1 9 1 0 9 2
9 10 9 1 9 13 9 1 9 2
35 15 13 2 16 9 1 11 1 9 13 9 1 9 2 0 0 9 7 0 9 4 13 7 15 13 1 9 2 15 14 15 13 0 9 2
20 2 13 14 15 13 9 10 1 0 15 13 1 0 9 2 2 13 3 11 2
7 0 0 9 13 11 1 9
21 0 9 1 9 2 0 15 1 0 9 1 0 9 2 1 9 13 0 0 9 2
22 7 16 13 9 2 7 1 0 9 3 10 13 0 0 9 13 14 15 13 1 10 2
16 14 10 2 14 15 13 7 14 13 1 9 1 0 9 14 2
21 15 15 13 2 3 13 2 7 7 15 1 9 13 14 13 1 0 9 1 9 2
17 9 13 1 9 9 7 15 13 1 9 2 15 4 15 13 3 2
4 2 13 11 2
36 9 2 11 2 13 0 9 1 0 15 9 7 9 2 15 15 13 1 9 15 2 3 16 3 1 9 14 13 14 15 13 7 9 1 9 2
13 1 0 12 9 14 13 14 13 9 1 0 9 2
13 11 1 9 11 7 11 13 11 1 12 1 12 2
14 9 13 1 15 0 9 1 9 1 9 1 0 9 2
32 0 9 2 16 9 1 0 3 9 14 13 7 9 1 0 9 2 13 1 0 9 1 0 9 0 9 11 11 2 13 11 2
17 3 13 14 15 13 7 1 9 9 14 13 9 1 3 0 9 2
26 3 13 9 14 4 13 12 9 1 0 9 2 1 14 13 9 14 15 13 1 15 7 14 15 13 2
16 10 2 16 15 13 10 9 2 6 15 13 3 9 2 14 2
11 12 1 12 1 15 13 0 9 1 9 2
7 0 13 10 1 9 1 11
24 7 13 1 9 9 1 9 1 9 15 11 11 2 15 1 10 9 13 9 1 9 1 9 2
6 11 13 0 9 1 9
20 9 1 9 1 9 14 13 3 9 1 9 14 13 1 9 1 9 1 9 2
16 13 9 15 1 10 3 13 9 1 11 1 9 1 0 9 2
25 15 13 0 15 0 9 1 0 2 3 15 13 1 10 9 2 1 9 1 9 1 9 1 11 2
15 0 9 15 13 7 13 12 1 11 2 13 1 11 3 2
9 7 15 3 3 13 1 10 9 2
14 1 10 0 9 1 11 4 13 3 0 9 11 11 2
7 0 0 9 13 11 1 11
39 9 13 1 10 2 16 9 1 9 1 0 9 13 3 2 13 15 2 9 13 14 13 15 7 1 0 0 9 2 14 15 13 0 9 1 9 1 9 2
15 6 13 2 16 11 14 15 13 1 12 9 1 0 9 2
26 1 0 9 1 9 0 9 4 13 1 1 12 9 9 1 11 2 7 3 15 13 1 12 9 9 2
6 13 14 9 1 15 2
23 7 7 9 7 3 10 2 15 13 0 9 7 0 9 1 9 2 3 6 13 3 0 2
24 3 3 9 1 0 9 1 0 9 1 11 2 9 11 11 2 13 0 9 1 2 9 2 2
6 2 13 15 0 9 2
14 0 9 11 11 3 13 2 16 15 13 9 1 11 2
26 15 13 2 16 14 13 9 1 9 1 9 1 0 9 2 9 1 9 7 10 9 2 1 15 13 2
22 15 6 13 14 6 13 9 7 14 6 13 9 1 0 9 2 1 9 7 1 9 2
12 0 9 14 13 1 0 9 9 1 0 9 2
38 0 9 1 0 9 13 1 10 2 16 9 0 2 15 13 9 1 9 2 11 2 2 1 0 9 6 13 14 15 13 3 2 3 16 13 3 9 2
26 11 2 15 3 10 6 4 13 1 0 9 2 13 0 9 14 15 13 1 9 2 15 14 13 15 2
20 9 6 13 9 1 9 7 2 1 0 9 1 9 13 14 13 10 9 2 2
39 0 9 13 9 1 9 1 11 1 0 9 2 3 0 1 9 2 15 14 15 13 1 11 2 16 0 9 1 9 1 0 0 9 14 13 1 0 11 2
36 12 0 9 1 11 13 9 2 0 9 7 0 9 1 11 2 0 11 2 1 0 9 2 1 1 14 12 1 15 6 15 13 1 0 9 2
